
`ifndef GUARD_SVT_AXI_SLAVE_TRANSACTION_SV
`define GUARD_SVT_AXI_SLAVE_TRANSACTION_SV

`include "svt_axi_defines.svi"
/**
    The slave transaction class extends from the AXI transaction base class
    svt_axi_transaction. The slave transaction class contains the constraints
    for slave specific members in the base transaction class.
    svt_axi_slave_transaction is used for specifying slave response to the
    slave component. In addition to this, at the end of each transaction on the
    AXI port, the slave VIP component provides object of type
    svt_axi_slave_transaction from its analysis ports, in active and passive
    mode.
 */

typedef class svt_axi_port_configuration;

class svt_axi_slave_transaction extends svt_axi_transaction;
 
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  `ifdef SVT_VMM_TECHNOLOGY
    local static vmm_log shared_log = new("svt_axi_slave_transaction", "class" );
  `endif

  rand coherent_resp_type_enum coh_rresp_tmp;

  `ifdef INCA
  local rand svt_axi_port_configuration::axi_interface_type_enum slave_interface_type;
  local rand coherent_xact_type_enum slave_coherent_xact_type;
  local rand xact_type_enum slave_xact_type;
  `endif
 
  // ****************************************************************************
  // Constraints
  // ****************************************************************************
    
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
hVoGPG+ya6YnfRjaTeEA6LUf2azA6QnxP+9XeYqCo/zbskLTZSVgRMI3p4BAXNO5
9rz6WOCMGCFv9w1MYAXGlyx8cepqEDmdJPQ0nmXUwUXQgBwVAcA5S5KnGSPVBLET
4bVRd1Jvg2UoEf9kinma5WcdGigxqKJxk0NSXJmf7Yo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 328       )
FMczhrS3Eq5FfVMFLOkB5FcnO26e96AYkUQWNvMc98Dcf/MtXrZbT6VNlSn4+m3p
xN6vX6rqPHc6pAdjEAkLAd06/Apw/+rOoS1QhcUr55yOy09a3IRM3mrqDve4V41H
pWPxj08bPP7/AyUTop/2Rem8xNpBOIFI60cGADn0mrEA3FvrpUJOjuk3HC/OG7fG
VIx1d2UMXLVgJIOuFQQLDF91N/Id6PwzjmPdtBM7VLVFX6KtgfhWEoAgAbKvifxF
RCBhjQtrSh9WfrW2SkL9KzlXt8SCzXR0Gl05EnelR1LHIjgpfeuUXn70w9lm5Jr/
tDZPCfOCNYy3Alvo237nPnhlHe8LJ7T3xv8a3j9qQdiwBEtRYnoCp6Vhg47rh+P7
Gp8hwMNSPJvkeK/4ekq3dB9vakMZfBUY5QF4PFB0VXqGG2NIaTEuyTtx9Ep+a2dO
`pragma protect end_protected
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
D2+AwW3mdXjz8+aPyLyObIEns1LGGpHGby6gw/XeE2YqJNt6C8TuXLIF7p32EGaB
xkIauOpkJ34l3wEJQi1cUeb+dB0PHLcITOqYgVwNSlLjxh71TE9MBH8b+w9U1xZo
GRfBuGQi9PRq+sVz54pJtjMhkp4u/6E1YO52JRXHrXM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 29215     )
7PPUgVlYjXvwUtx//u/ddQ+2RTd6cf902+1tWnbO9htIuS5MEqay/A6Rik2q3RhD
rZvu+zlyQbBVEc0xhlQ7jbsYuCccpYZYvl0t5p2i19l7X5hGfCDczO+zVo5E0BsX
j6lv/x5h1hcand3z8603zQdtCuDs3NXPGTKzX3rJsKr4pq2SVhrqjZKA8Tu40fCh
xLWRVKTiGQK481EUHUgcPp1HPZA1QwJNPx0DexlwD7HktJlE2pLixmyikzyfdTc6
fnDrgyZXuGURGJBbSKInKMX036HaZacq2qhRqIKaxzOOBDvrPudRza2U+qPX+SdQ
WMD9kW0ZlG7SwEHX0LWMWah5OOGD50Z9LlwRCWtToYYTdC4ZMLbqZd1yTFNYFjmj
2LyQJXDBPUil0pBGn75Lp0C93d0JCnA7xAfPyTI22S6/kyKNIhQE5sZIGS6NBd54
E2A+UffH+W20MylZpGWcqr3wDRrnhBrNjhgJC5xX93QaK7WR8fol1Psa55wJCwb9
dT4ddiOQDc+lVvEwnAmdNCWg4tRcx/Vj4d8vDES7jbKPocjhh0+ziJStNvTxLj6l
Pr8z7iHRMaIfsuORvp9wSKMSAb2HOOscN48+9zrB3P86BQsF5b3+kvtfB8n6qIYT
6p9axXhjJ8LCo0JkwZdqgNsDJvw+Tw1L9PIcMs3or7Zz2z2fxE33TZYaTzduXbIR
TIfRosIIRGU9E7F0638c48QujCarfyOdcaNoKyUZ7CIWBSKNiAc0/SHjfddeB2GL
dR5WX2cOH5FrZ6InL5u/IKcFNuvEaECqiDnMMiLLLG0xLFW2oViirDBJz0H2idfy
+tMegPpEQejxH5J/tjS2HaQXlNU9HSFtExZoExjSr9A9OPx8wqW+zxmi1B0Cihjx
eIYBKBQ8rkFvauiwWPl0E2awTHKl1mOaShzP2pZozdHZjCxeCzzEUBQDJPAkL9oD
yqxM3PJuChWoV/nYzLvbG+zE8Ka6VkrmxzoDFjXCuLKqvGxTaUB9m1HafU+xHVIh
OLEiOkzqkr5iwmg5i8XQ0X8AtU8QG/7/M9U/rjfK+AB+SWwjSI4w59Tecptgwmcv
jcIzDc1b6DKcxJ0cMjfJnsYRMaEQgkObfZoMsZj813z2qKgOaOw0VD37vvG6HxdT
oxv7XhRCMZeFJMdTiUomqt7XrCEh66MVxnKw8Enou8cRcgKr1bOlVxO/oOP/kaQJ
fZQjhbUPNi4LgdnLJV9RZHGWPDBrsWPJ95sK0uWNYFFReWZARyPh8xZO5gH7HX+A
moH8r9EPjzhyS57/Dua5dr4ZPsiTFWB4xhQelzF8DyC5412wmJAD9wc7rxlzjW9W
ZK/X4DrA2gLkcOnZUhnJHUsfyi+yiOlAJI4bTAGuTF/TKPV5b+4W9M5yvFvpgWkv
AocWr+S0vvenIonKethcrKbs93pE0C2ZdE3MigUZGB/8h1TuedmAAopv7rIVWVbb
+T/L7yEwA/S1I7eFPN/pQFGtWDzMbM2MJWrFUfothRWtdII7b11qn1mLEGKhq92b
37a3XeCDE1vlvXMnoGmVzY+gyHRXtT4MQnjnVllH+9Mlp/jLcZuQy2YhPMvECpo5
Do6JTN/ZwglkaeQ6mylDLpxXTDvyeew+TiEfzaLqxKK98L4TKJ0ZFw7iVbDHfvUz
ecdEhwNQEgyPFgu2vf09mUsVgoZzilBvfHvO/p37sBGEGe6XRefHnkiCmrAUyFa0
XgGKdrvw98tMqBf7bg+guvX1PPtJ5dqv3Ij3JJ9BEf7HYxe/Swy66aYiqEIuf8s5
345xsve+O0XDogPTFhOHIw1sY9z/BYdbzHlwypJ4Q4UK53o6fFejJyJzqaFXVbD3
GWskKadv6oCmBIyG07fMyAicRMgtvuyIFGjpF2r+CxJ0+oOmjsbvHvzik6ZXae75
NIzRjSCRYtDuz6Pwdc+wjRJ+anhgtmmb1W+SypWbzA2+WRUeqssp257vUq7iilNr
LrwFSSuS9Bu0cLLhO76+ukseKTnxsExUCq5pId7AIR6Dn3mW2L/ydQjgIKbAXcfR
qpZyXlt2GHLdLSf2z7CRg/aZoxEHfHRJqVxHYCH2sJBAFqfWci6gqi/aKPRBbVSG
ZwRSqxpjDMF579icYvrUuGWQrRgh96Cykx+JiNViX0keXFkD7dhwB0WIghjDAxjK
N5HFJw+zUaBauKIeAskTy4S07d60y6AwO5Nrf1U2URQtO5HAon14Zg2rjxHTEJ7q
rS+XNRpNcja5FE6Lf2EkeCQjYtxfasJppiPUxeotNzd7DI1sCk722yUNoo/YBOCm
zTLLUMJjZcGuLBihezv7k/nVy+EZf3r+RytwmvgJPo/jpwOLYb6UUpy13ccRHXGW
HTpMhDyMGomHCNcRSJtOrazr00puot1Rb7S1IKh5wFFmu2+SNf6eiM7OqecdRlT0
vk6m6vZvI31xMvO/62ISGhv4u5XkwaOm43v9buS+OMkNyQRCa2MNA9hUx+dbxpT+
1XJPiZSVf7NHcRB82wfPFSf/7SIQy1nPZnE79XJyGW2Koul3PFyTiQ8kUeWHk5ZG
WqRm7rsxvsLCWcXhFHtfuF28CukKy4YhOa4cc0Wwag3BA8455OJ9iQaxin+hVroX
7wlYK9lk5lz4L8N4jGnYtvGFuJ41gz9mMUj66Pof/UKSHqhYzqbGBkS6Stn3ppIc
wB74/qLF5n9f/HWHKsdgq2DFhebYJPY3xVXxkFaUdR60URjZHb0OtcN6lQjeMTaq
9Ej6FHRlicfskbvkX2XLPzZzsT9Foxk58eSigf+69DtqGUxt+bb9sPdAdvEnWm5n
MJAmQg1E+YQYt4Vd2V/H0MX+i+SwpwIFHH1QtUD2XHxJ6nthSLuf47eDpYoWLEWQ
f10BR/xS0GtKTW8kswHSN9TUq9Kmo8EQUgay3K/tvrloHQaNEJVzwFZwMupuZEmU
7cOCvk/SHqPGX4+kAiH8tSoJt7gPLQgJ+J6lgPt+SWBVgJ2Vr2PAA8NERCNIendo
kWsdCQOo6lmpjocJq5wKW2GxVThxSTKsmNF92kTZAumZLLm1U4VXqPGnPan6kqwA
3gprSIeFLPWBwb4tZp5DNxhySwJqrhllhRGclXrImx6V76K27rFzWN7Q4v7BTdYE
sSp9MyltJ25DBluUR4ETmnQQ9abvv/04iopihLJ48fwYy3cIuZ6wo1f72d5kiAJI
VcQkh5hjQDIZwSYiQZlofkia2vWRZkxmdxDck2ZF8XjcqVBL94CZUxcA6i9eX8Ng
x3vswWpmSU2gvpUzVAkt68xpq5T5IagTQGrRsFqtC3l2ib2a/dePz8zVtar2t8jq
A83i3qftODiHsaV+0T3l6cIMhxRk9J2CUoEGj8E+Geg0PFu8hiNDopaDnsuDjslv
ZbKOC2+v0ssGLpZoAxqDaRII4lCzy31QFr9Jcw0Nx+O9ZF286F5LQqctCfr07MQs
dlsuyl9KgdW/Ho7RkNkNK/ex6ny3TOGkM6cT0IISFkroN8Io42hXwevXJmeO7zl9
6l9rbgfVRqYchxDIB1lFcDubkt7Ctbz0S+ZkdWHqu7/fnpB+uqE45b2jmLXvY+lu
6dPLR+c1OdDSWvN5jAgJk1Gqc/cK0n0m8XfNTYDGpZYfs4qVBpyvr1S8+U7pYcqD
OFhA0LDGX2R+WP7W2CeFvfDV170q7iQB/WbYt1xuNIXXok/uxqxN0fdnhXdRi2tN
iPBIxuvjBfj81N+3LiEbDE0athPlUjydawX+HO43CURN0P+H9sKSfKYB732RtNV9
cZV+6kOJkhNgVGybralNRtNSpOPZkwWnJV11v6K7jxSnGTdjCbDKZPusIGPggNpZ
uHC5wskDP3t+9z7SoKExU/Au0WwBquEkh8F4lvZA7eT4w419+xQvzOkykP0du85z
6WUmyOJpwyp0C/FvY7FeMO7MB6q+aBpx3b8iNOM4UBPHiqWHTuuo/cCyQDlmFBKb
HqfbWt13OPLqr8fzGSRh+9ZtNozbiMh7CVR52afrgQeALjlRaq3eRNlZy9S4y0M3
jwloGe/Tiu4SGQkfD5c5JJXUmr/1RGqmOdOB7Cwr4bwf+MgohbbdlK0Oq0EU9szn
QNBErPZX9YY9SQGnTQLcbvQvBq9iy675ZTpOMbURvXNqLNAS2OPUga0aK9eMmWbb
evLglvxuQyoBZ006KVUs2c6qoDXGQpjejHadjj5BA3KBUIX1usjuDJE+eEc07IYd
rdW2+GeB9Uu8UVcCRAT/KLJ2UWkn4V1NAwCQ5HCccETh3OaGrqM/Z/9oW3sWyzU0
k5CGGMEXvYV5GJpiN32mfqndCAlFg+wDjYN2ILJpl/Vn5n5Drwur8wF6rk9Eu35i
WbhQZ6b6lNgTZlMpo3NO8CSlh+r7oR24XEC12z/q30kK1JTF10gU9CbXLmJPVW5X
N0GlzaCTZs5PcJZ5yxxDSUOxkQVDroWjliHj6TesT6byXj1sigAqWPvj5DAMrVWI
2YgazYDuKGjY2Zcius9SG4clCyXkequLKPWDoavwJwdVvk8TAE6KJ3Kq3cWHvfdY
BI1IIZtzzSvvu2378C1FlAAgefxHVZFHghxNKK/Oz+VehTjV29UQoJti9bdZEYoO
/HDiseRL8/0ANBHS+FGNGPxDJdR+HBlNS9OrZiwtTXmPsLA31Td5c3FhJfnsEEVJ
p3zcNCZ7oQ4CEej2lFTpQLLUug66npk/OmBbX1v6QH8BG0wwtBg3ZdldO243pFja
rNCJ3CB0OwR29Y6AxZMCf2TW2jG1TOwsFd6/k4/YJ0rutT4zFtqa92n1WryS1gIB
bqckAs77QYYUqNxKLcexB89ujkzG5wAdqFFX6bclWJo5K+ANLyvuUymOpW4j3zaE
fhWhRTfnHcdIo//0pIbXtP4pWVgk/woj942ZvPLoKk6mHnNAdxz2ab1d3mRU/Qp5
rPip9bA6nh4AZBLElUMD0um2N5To5KhANIldxdY2KAILfL3n1AUOf+zX6ehe9iVQ
dU+STsBUmbq/aVt61wa2HJC2URejqeSQ6J+KVpRHSp5v4gDdb6E5HD6pT31W64/c
dOpg/fvNoAMMahlrbCMaYwXsFmMyHrUUbi2f5bQGcJevwUG/PEWgn8vjgryY7euY
vuM+A+lIZHjNjC/sWIbYElKn8F29zMVJOq7vJewuyeuNYgpsY9t7jNQgQTCoK20Q
nsRdD15flvaVCqaDaKchWsb8zxxcdByynewRVQycqAULHuA/fi8LvsVV3Ybn0Ve7
hO5HXJo/El1+2i6M6Xia5GKQeYHcJgjJpzJA5NXaNuE0txnu95QS/dH4XEx6kBps
tqE4dGvEx5orHLjEM4BfbsdHgSlTIrvVov5GyCbKTXJ3HmWwu161ojRlqUswl/kL
5sUQvm/TixPMdegB63eWqJsNLyqiyyz/XixYsGEqvcAFcz1aHVdufV3nfkTNM6Vr
07mQ+Xg2A1p9g7G27pPNLFTKg0qvSSlCM8NdnGwD7yHCS9jXW0Ex1k0Owg265blJ
5jamR8wWbaBmLbNIJcpfA8l3Mkrlq77SlAdLRIfwJqqFdW3UmSMUcVSKCBqexX2v
7zsCvLRdqXI8NUlFQqzBBH9JviZrnGAfmA16L0U8N3LEBY1Us04hE+GK23spcZQ5
Btjd0gwEfOxvI7rmafsqpbJfpaK6PvVTp6JleW3bZmgr3EqcufT6HUnpUwBZ2RT4
5lSrebMrqrob1HhQLPt+FrJE+gnzazU1gksWOF7kp76sZ/kjTTlGqCOm6lgrki7S
4FcYvA/jw/ZbAMiOkZo7FAWOSb9aZA49JdiyiZRbP7lC74GSVeHgKVbHLGU/mEgx
O32uXTESFzDm/tioEGxgG6S9JrFKGZrW8u0PVa8hk/6FtfvgvAZ3wlbTe5H3bCEw
C4tyJ0GbbYDHiU5YDnsWPV9sbdQ+aBxM5JHgK4/mmiFJg66j8zmuiJqh+R5q7XbQ
7xdIl3n6CwOR6SaY0Q9loSI0gb5hRKJ1x9HxZElSKhRBFI+OATUfsk5YP7NKTYsT
fQs6WRC9iAe3PbZHEXAwO60Fyn8UlGwwmiCtr8cSU9JyEOjCiDkzlyLl5G/tqV6g
cVhYVPQFQhaRFnZ7XRL8a1iolacOsc0CptWQInhcUZRRIpNzETVnpn7D/jsyLRLt
ciCEdXEwW+C37PCBa8AcM1kOaO4ebuNAQLWp3wixWgDHZS1j93TNWsDKjGsCCpjW
0u2ZL7/NQTfWst5QHeYOdKXUbOHBX+zWgWnzM7zSIdfJLMm5Jdal/IP2FdyE47yb
eVA3gvOeNiSIHup7BkTWiQdSkKCcTznw+YSRvDYCFwVU14eDjfI2XKORlj7HdEOC
pWYJd+VYqBKLODjzUjrr/OdvcBxZ59fthp7tlYBgFUQpjmdpyFUqSBPfrMLcaojc
1kwcMkjpgYbThMZ3uiXIP2Y+73uuo4TQp7zP9I6+DHfh6RbEKm1PXCo04RspEPr4
89FxqKnOrVHGKMAWdCj/jTxE/bZFKSPAbAPDZOuwXAWIFN2eVl0KB8Cql1Yr0UOA
UOP9L3ppfedvF0PbbkDeH7ArVPwNZYs/tksiLBfnYVBoe+Du6TLTjU79h2J7TDOv
6dHWGIhF7zsDUvXDxl0CiWP9TrUFgt0PpSPkHWr9WBGl/6jtenEG6yRq0ADQ36jg
KUuYy113K8bRRhvw5SP6IOqqn3JXQIZEABHXq9y32Ssbp0nct20ZX4DxkiwVdHfy
h9dzQr4lAsDmnEgT39kOjZE4c3Ys/JX6z7CEbX97f/TNQSccFxHOVNieSh1mck+1
v+9yqi/Awb4Bzz4jgYlICA58ogR4q+zJnP6paGLmR2AuJpApd+bDr64GwUYWosTQ
Lj6tZOnl5YjhzLmWUo3Wi5vKGYfLO6UC1RP3Z0+/MqwZk0XIudRH8eHmbe1VVhBI
AKDdeTUv7b7sDxlTqdEgL5Z/GCcGI6+gF+gFa0snYgpzqqrXM1NEmckNME9kk4lb
YrWdWhWhVdmrPjWt0IU+HR1Mi0IAC4+LHsENZx9I29NCddfeqUaPDwE4XBxgYHek
aDR1PVMh1VNRxThM4CE0zst9xPXLXp/HaqNavQUN4l9xqnt3PBtvb6WbEFvZcXh6
nEHSRTnbDy4P+RLiDqZHdX0LUOQrqPUYTVKunxmGGviAW+U9ta+a34jsRS55VkCH
9KR8dtJZnU+5wqWC6MmRFgFDPshIfYAiTK42aO3+BsGvfuqLXghNuOFDT3G2R0nY
0VQENh5IteJZfDJl7MRP/2wXWLHJ1hm8AsyxVPpOTHR8GnvmZ+HRc8H11eTpV+Z0
o9tWaUU3pkEv/77YEMEn56oY8poWLeyeel5bdGrP7XVNDD3g1fL5zQVLAdn01i+Y
VfiSWRsP5SMBy2c7h+Ok3OgO95B+eDfoq54MKMURMeSkuKqiC8D1rHY4GWLmTo2l
XBZIRExdE1jFwmMgnmefxdo4t0OCUojeRTGQR2hTfjSip+mF5m+pYTKGaPrV7TBN
Rgz/PGPRtpft1wwY7Z/qYWLZ87J0Pu7TwxHVelxvKh93rjZpB16QvasJ0l8KJrpa
KopV3M4xseOc/UxVVz3qfmegMBMIcMudsGX5k2C55HvrNWlqVdFU7p1KP2GuH6St
X2CHVZy/XiiB1jlo4x+G0k6KRqoNIpwA1kaJTlqfNsCTAjWfkVfZGtn9MgsWa8TQ
RNRCziRi9/yyQhwGHesEoPtnBaAvSyAJImecuYmFI6LA2eQbluYhVN6cwzUxsLlO
XnnUSkKnE8+jf4/rx13yFkEJ4bycQFjj5XSj22RBpe8Ki/EuzmXjChchK5DrvFCu
BUQn7cKnFlSE6XjHoMsXIJxwUSwRwT3RPrjSQQJKqxy/qh0oy5/4R6SAOpYwPLlj
CZv+V8E43hMwlKWPjuVXj70bKWbQfkrP28P2ds24RY2G3yKaYwa114bMqIIKFKB3
0HGamroRBWhoPj6ejFenDujUTMNH1C9w74hvFr0VuyYe1jghYY6qmkQxqf7yAalS
vF3uDEkqRx0QjsO+1RGnGyxsye9M+jg7O2tdFmR2ahWOMVlQNDf5AvRtRtfGE7Jf
2Em5FDmhTh/QpEYDCWiMmsLHO2WMMWkX/hDAEEuth+OfrKLoB3HBHlk17kRPcKNz
UV1b9GbQJKnJMpxtY1nKUaN3DAJYogVT3Gb1958fvyM4mRbUs4rqlPHgle4D24sA
0EHD4mfRvFgEKPRnpn6WkcVgs0nqSaSSVCnzIiBPuZz3itE/MPWVft2ij0WauNzb
kLCa64wBXtfeNXN42pq/vByzUP7IOsj6GmZgOu/uFC7TQzcO3dReerSvW3Jg4blE
5+pc4Hi3lBoGZPTaRnxUeFzapWnFfbMnAB3TzXiLgvdfbVOPmC8A3lwW5oCo45bq
bznaLB0wzv8utqUg3V3yh+UNvoTtuRYrhZ/qCZegtLqBhiDR3q2yM+0lEx4Z9szx
Igw9Y/nJExneCjOw3GDkUkM9U/ah09S55f5EXxSsUSYiMZ7D4OPOCJCi5Y9KvFHN
PZyoXNV/d0mbi/D+7vyvWWIYOoHABzzQJu1u4ionty6j9zm/9Bk1UrM8eI4uxGHE
DywWP4iTC1VdDUyMHo5YmwkbzeV+RV1xYxVH0c5DsixXl+XBzby6r0nPEU+y8jWa
OeA0IKqit32lyHjYcbAvrqysqmnHMGxnIk7P08hOFuctX8U1lEV8V+gW/fKUVPMR
XKUlcEWpM4CfxVMAj9nE4j1JW76ThKJJrCOSYgKwyIIVqA+CUB6RbLEWer3TDdXM
zQydquXkWZGs0Pp6uRTeOoINIvS8MEl5Ayv+9WgVOdW5QxgJc2idw/cbauFdP744
3DupP+p81rHfzGHR8iMQFsdy4TuJb3PJqa4teGCfxSEjVmJorNVErnLFOjdz5X0C
jntdQQoRJ/AdcLndEoTj9OwkTb88FoP9Y48INuziYV7Vqq3GC9SNsh6WGzgipfbd
jKbnbUeObLFxj3ZgaHp8hlc4fPeca9ORnAdNRaHQMfykGo6PpCAflTdmi8afDbn+
M7+YoQOt6a+bXNcI9qXSkzveW1EnrUj4KyE1Tj/zj09qB+2IAwemCPPS/ilSB1qN
D3NM+H6GpOxJS8al96vGzvzqfHslRzKb1vXVuy4xDYPY7dPHYM3PM0XTZnHor2Tq
g0oHQHWsJ7vhO9PZ0EXrr1WA156NuKGazxMvg8bcuQ0eNcGNsriJt9tTbDmKJrVY
taliJHG0NUVZjds5ezu0LYvc7sNxxqEjaroE3cIi59+q3ZvcFDamHlJkFTj/C8OV
sw7KCnJzZOSrs2MfFRHMgoIZxkD5d2IOkg3NoEyO+uo/j4MniZlQId5ImL1EAVTG
aDPyc2ncERG3k6+qZT4l4j271K99/umGCoYgREaJCY0RlCoZZcxKtdR/q9azLEHp
rawWoUZt0cPmaM7DNcOHj5bdOwjYOEz66/QQT8JbcPuq4h/l9DftIbgDA2DluuET
kqXCj3y00jO3aEz5Yr0oo7CC9Ak/sbpYX9ZRF5XqBX/VQaQPfkmgicH+V7hNnuTi
5ukpGd4xsszHWPN9AA2Q0TiEAmr/WQQrl4Zk+d5P4kNtw5xczZgNL3ycJ2L+AYnU
s95mewF4+0faD6Kz3kQUC1ovzzcF+cMtapRZs4CuUG0yYWubWs/oubuG/5Uaocpu
sDr5rYMM1kbaDotSuTe29W5G0UXuz48eIcPERlsJEsxZI7DpBphHjgKenCPWEzxE
aECCK8tx2Vhm1PDwtiI3b8AzRqYt5Lm9Pu7TwU3m118G8t4Q0+bGQxkLEZu19NiU
O73ySsH3KDeNV+pT8/4FgwSrN3KAX1sNCFd28GVntHuKYbwX7CkyXdEV59NGpukd
sxGOFF9mh0Tsfcm6NGJjrNm2239rReKgZ9D20JbqsNv8JtQGiwCtFbdS2X4mNpek
gZMv+UTi4f+dlr8jfxL50hDVYrTP4E9XPMDIH7onyIQnxStTTzr7I9FRi0ksm7AB
biitIU7Xz2+HqxkPtEuQy3NBIlm40rpHU1LmZmH14b45aCY+E7WDTbS6jvzcIgBB
8+V+sctpKi/AS/OAA/GQf/DWyPJWEvgSDdnHJL0lVd6caBjGQCmSbdfjPx1Wxf7X
ANBJAR0eqArj93DX+1WIoY8C8v03iMJ9x5RyMQPwYDJ+zfUpK61KPtMaSQRxNfIw
GZGFitFZdmIT5uMH7QYOvT7Jqvssi8bwKMe61e2MVKCjf6M14kq18Jsn3Ey3NhNC
qbWFRoMUwznPWEAQwEQsrjy4Y9HUZTLROVEWGaQ9vAYHIJeo9nZ+bfrr8ai3cA7y
W3hJD+yAcnVs91b72uojWzzH5QBlG16D72thB3tB+iMD4OFXYhaG5vq4zl3QiCsI
zgqlvuSQYFEhlIetlrBWfRF+Q1x3Nk4yy8Dg109+uk4iW406pYdKqfnPj7RtBdXZ
js3773jjmuKBC2kzq4/kp+PG8gHM3GIlu5OSUhX7BUO5POcYfTlnhaibnxTxeuz3
m72+EJ5s1otiYMIajrqOF+QWTmDC5XlxzMYvcldYWhgD37fDBcI7WM+xmivDEjVV
GY3ZT4mVLjSbfM7JH32obOLQJfgzVNlXHmC/X7ArBrWZzDn1d2Sb1HlU7TW/KLbq
ImH7LwLUelJ7EQ6iPBveBaX2NNbM6vdUwoWG1WG4M/Hz1kt0KubxTTr6LvpDsb6t
VLPip6rgCGlHgr1g8y/MLLcoZhEb57E0LEgTIkrM3MIulYcvn/a9DUaAYN+mvHIP
CV7fRN6kVAXMy3xL3HwvKbO9YA4Pv+lkZmM1NGgpiqcvhUitrO++PdI7hVWwMYW2
h53O3zFuBocgX0uiSxC40jiw16/Gw/YKfCDyTXsKYEQpuFiq4ibrqSNUoqiQOdCa
u7YMTaIUPgq6L5p6E+63UYXCnarOdnNLYQd79nw0kuLdraLBz+7YYKZPASWzr1aG
0kh15FSyD4jWYio7locR18n+ZVZFBZubsAW3y1DAJtc1dFYX1NYo1+gmxogCPaz1
57NjaiB3/JpM4oRYCXXnGbSdoBBgNBiM39QkJomGDHnLcHV3aH+1+71d+kP4vkcA
5eL6qzO4tlm4UMXsxF3PgHQDNRDPCJBQlh1JF7CzF2UG6lhL0uvlch98tqT1Rj4/
ngW13y+rJEnyJF09uppC0RSeB6TnEN1sUcOmeJneydRWZcWdxWJ14pYNgWeLOTet
n7BD5lC5Rw81P2yoPcLduFmqEUpaaj6oMPcm1yuMizGHqMO9o49VopLb8oTqAZfc
g+gkQAERkCqNtRKwdi9A9AYOwNOVZ2jFqoh8hrTDZnz95VItwqXPJscGZxThCNaU
2yzCUV6npsM6oUDdhdcl9g1Ajz4qRS95WS2esgCwdDCW39ZeIdsNXYLH0o4U+PGl
XlO3sG8PeuOnNXfLFPv7+ePL3tOm7abclZzyfBP0ZMAFUeOtFHSYkT68HcvQE57e
NJHF9e53oLYxrJm3hwwOWO9xv0pbP3l2wK7rlGhEbxhO0stH35uKF8exctRM8bDg
mK2zk1k6HrPxXddc7i3p2V4osVxe9DoSqTxd/x6IttTYIwE5nAG1NIfp4zcZzTAk
r8sq/saKmSr0FIaf6EWxfXLd8laRzVlDE4+DMOyK7JtQ2MvjPE21QEc0g/VxnbsT
TjKWzdxu6CjGjdwcTlJMSNBKNMksAeG03yKgsFZzGONKvD2BuvtLgHNfXln9bjM+
wMy1XsyFOfIsOl6+Hw78d6wozvjHRUFSD2hlnXBH/uIenGJeWF6spA3sdrXD/bDF
zBbJggmYwibMsr2LSbqoO0vpxaha4+Cptq3nc+1q+UvEhrD9Orky8VnaHCvNHVl2
T1+mxVbxTolCe6MfHtPMxC1J9icRyB38gdHpr/+NUTpvMXz2S1ObY3IITeTqNgyg
O/yQuxJ/0kQH1kzod4bukCFpeFpjiNLBm4LXTG9RJ3hnRGoYAB/STa/Ys5KsmGKq
ShYAHBQmfcvrvkfPkshAybOOtkh/L21TwwXTUQUQDE1auu86w10j1Y+jotIQY2R6
KiM7kBV5yis9b/qAS2yn0mWNsS7y9zQwzPJqbIO8M+ANJwBDwHtCu20UxydbZ2tO
9JopR/evsaBYsaODruy5Mqf0o4h8o2ZhLznkvxExTQ8JquEBX4eoI1I3YzOijL1H
OLvqZzti4W/xHLrSK106iMw+qMK8taJl7szIdhZ0iPhWX79Brwl4QXQqOtmIN07u
ylEnUvUVeR0vsbLnggXU/ks7zqdk2nUUkEIYHYcQ8IwQ3YTrnm4w+OxvKrfxVfTC
GwSjJO99BvQxRkNJ6fWHoHFjsr3043pePSpWvYT2H84Ekoryc7dUbmGAHq5ceppZ
2XZ/iIYR29mvIT7FKxiCaGq4kZ1AXwY0UWt0yCKa6EbWxEONMYefRtvc36vk7ajD
suz4hJ/u0zO1YuGtrpZawYUT2egnYILQQKxAK+b77SDzzTw08gcQw5JdyYr43feP
6zi54ZlJmtxfYaKJwixlFYO8RTNWrpdxEmHa6VN8KCyThCj6kcQcpfdpJqBRR7Gh
22Jn+4KWD81zLllgDAlRvHDKwpdc/J090UCrVwFA3t5W9AFDsv+ufJLUoNGI29NI
B3qovhfjoRTQKlagPfbbjsbTO3Llg0aWPF5m1hssts6bLfc8+ZY+wEt4ETQKzNVk
esQf0mWUeUe28f5vcfuUupJlXqrYRppPkuWj5aZXRKP9+Pi/MOb3N+OY0BKOQs+r
eqKeBTIwQ3vyBfxUREX34x4C74UJlpKUflXzQuOjilz66h94xShWKRhJ3HSLL9a4
7tfyvNKjYCiEmcOTFT8lAyByBZrTy3wwJaTnoP70xa2UbSW0wbtdanPPqe8qsdyW
hmK9kpehEJXilQNB061zGiaiYoqSV4Laic6MwH4cdtNOc9SZf4PjZ/2OCrM4jRmc
1LKUXBjj1kHq2/cpNMXwhbtGqL/mwot64AJWSarY99cCBX0o5pZ+QGSM1r+A89A8
+M5bFIFatTNV8a0Ws0WwulluTNSc4yaTGch356hHBCRUIoqDU9rLyEHlB4q8CICZ
AsQUL2ySQqs/XgIxdNeOYi8+D6bN0G0R+dHUqmXgslA0/lcq1uPg25OnOQGybbH/
0kEftJr/ISu1t67FEhxdgtnWoIMDoFJFrWtCS894zdi53JPjgpWPqNtQYesq79Vx
VlRovkCkawVc9tk9NMDSYylS5VT6c1v36cGinO23gMxsKck/prPhjuT15lnz3jCK
Fp4jV5crmtMJrUnRJsc4k42dc8ks16V89M8g2mK0vK5EX0emO+2WqKB8/2GJCcuw
/R6lX6yfDkZePT2bYjH53QSyuAw+nzfn5D+Z4drC2ILpU24KHB3xJVrh3A8ygL73
hUbIzryzwOUnGo5w3Cm/IzGlL7dFhUT2vK/ryOoHqPHmwmD7pqHmfPfrdw6M17FB
y7rEJHceqXKRoVregst+yimobvkA+rkIrUPqLLFoXlUaxK8MGZC9cyO8Dg4Q7rpe
JYTv/0KJZg4dNhMetz2HWywgs57OIlGQU87crQzSfgJijWtjKSFPx/YhEoLVtVP8
6VlLx6mfOi0KS41bjEYgel6wHzpU8NV1Y+h7Vsc6AzetVcakDG/RKlvWOnvsR6vH
uc6yzVf4gTnemxs4u2f/0n6W//N04lZ0FfKp3ef2NqadQpxNlKwyty4FwyexGa4M
6/n8x5Fltpu/YQHUIUIXyora+tIOC0DIEWtjxbHXU7XEhO7KuVq16ZWgLSbbniC7
nq8iS6pH0GTsply5YJTFJkd0WwDJt1oTdXLQIaxYXWD4z0sfwAgPAKL46DZ9EMVm
OoyAGffNInIMemrWr/Ur4jeHwVhNAsCGL9t1FCNUHvCP3EHCxCxKduGDgJl2y1OR
+lSOLa6gVMQJ5ws12m51WW0u04Mx/cbcrQ5Smjtbt281UQiV6N20dbtnrntNuXlC
qeCnyrkc5PYOZKOcBKZd7zABZiYf0/t3Cy4JRT/gYBiKTsxhkX87LAq+g9RPHlfP
XDyF5tbIU6xhU+VON/kXapXjsLQrlniWSp+hLudsebszoB5FxHr0h6Xm/KgBI3bB
AwAR7eFXrNYQD3inNtuHWc0sxZn6TSyrEFarkRFfkTDpNJ2CZAszn3E+SbhdAKHO
gQd9s/kIY9HqdwZAMZWvvOptJAtU5UWHwjJA87JSc1iPcqiMkbPoIWAISppBQINE
NQbEn88A1nvbEuXZQeH1hr7ZMfsltoYoccGK6mMd5M8EHia44rRUv6KpRBq3TRce
OHSb6cCUDeKSkctgTRfca6MZOsmttTb5F6N9a6bbV1rywpVexAuV8USs3K2zkaNm
hpwPkNgbyRifqT03D33C7vyL4Ga1zQb9YlvzM7guyy46m46ppsjKOLaOAdi89v0k
j3ZmJ9Sioh1m4Tn0vY5rgitfIsHXKpUwdvuatXpIbMimI3Fhjroyg7lkwjvpoqDa
Pfc159nHQ3rKDDHCVYzrR2UtX71TfsxxPbfvzlHBTBLsG5xkfLX7wG1H0pvEv7RA
LlcnEL+edy+gq3QYV17TksVA5+U2rC5mhGmtH4g28tZ0t1ovYsm9cQZkzmhd85gB
TK+mgwlwfKk0kzL8Lqwx2WU3r79rGWM/5CXhFDOmScEZjn3wwhlswtq65ur3WhjX
WNvVjquCdWbP1m03WlTWCl/DqDoGYkk5jCCaMIuiG/WlXBS1oW0wXofYV6x0r8PW
XdBnzitl5PpQV82g2WZDwDJVTvfKK4K8U4/4EC3JCaI8Zd2ExMrL19Vec9kz2P7U
2T7w79wzseP8lvUy+qX88NlWxfQV6cQJGtyvTFg6UUwJw/tXzbmDGWP07D2Xb7JQ
Opz5bk1Bapqwmj6LZcd+JnLAwhkBuse6hUyzKIcSRDfWcYG8dHSL7RYi0owCI7/Z
9YH9GvMIvUPdSmeVCNvvioV/5NUvZcP4BL1KThWd2ipIVaNcrrAEk4IlICeJiClJ
9fUUUt3n3ufssEl1idl7bwgl2v6CM7nd0XTAWJJ0Kbhtxd5pK5u/NW08imvr1k7Y
oxd3j/BkPpxd1p9sR2nkdN3mLkVzbDaMmITdcM4A3HigbIWTqh2jTKxgnZA26rcu
S+E3KPLcCqHLQ3aTmLpaUJYwu0mmWgIuijStmShEm8cNbLlHohlA5LdGkumzjNIq
oljbf+Qds10/2G+XGpx69c9GFA8FMORt1x6IkXrqNN0b/SOX5FaQzeflmulmEMir
QDoklp1YWtdkpLBuyB2eH6GAavAr/rel1woSHgeRXNpzNebyxjdHDmt3iV1KOw8G
h89DF3/IPIcmAf7qMZvMnwcOMZfT+yXFOoawXNE0TkLn25Ml3h3QBMIRSOzgvOoj
BbOdk0NVAYR5keNuBvNJuZmRHwYQwx/lYzwIJpT3tmVIAcsV7d2MKC9G+M654Fd5
d7ocD9ykkiE7qty6owsqJdb8X80kRPq2fgjlQQp1O4tUfpWrKXcBeELlMSWA+Ut5
CJ479RAMWw0uFcGp+BA2RVQZqr2M6dAMEq23cDhF8Gaqm8Bc0UoZLWrN0k23D793
j5q2kfC8OtxZ+BBt95bltFXZNxkCnLRIF7I0yXNeUUrnA0Og5E62+wCnDYw7eQkP
qufsAHKoHsUmJEmIA9zMQiUE6DexFA8lcb1tgdp5HQBiNkQH1GJyLfl5BDsGJW/Q
UrXu05YlOPVyfFKmZfSX1bxBu294s6WDMpZnUldJcLYdN5aNSdBCNDQa+EtAR4Ju
+whkbQapimkCdtUB50ulZn5PWH9wptylOCU7RJe2yppk3liZ72ycjmy0u7VXWao1
sASCS9g77S4daaeCX7EVnfNZ8nCkouG0hsYEmXzMUlNi1rwZ0dFS+EGQsDkwI8Zf
GFEJq6p1w8QCO/fOXH4+SyVP5w7NxgA8fqnQ3KUt+dxsceW8X15BIWmxSXCVvzAJ
r8RgFW9WZigX1ANROZu1e0cr+y3ktXWZd1naM19dSBLTXQjbwr1zFLjF2mcF1s5h
dMVQIWzzXRY02qU69G0uxf6/kbzfuFj3HWHTTWZINR68bELePs6wSQDYTRT1sFV+
GtREZWNzl82UfiOZFG6rDN7Dr8H9iP4wt+Vumx3IegQLO5ixgNuN5fPJXEWqP+Xj
QazISA5lucJ82vNzg/zvp5EA52re5t+dsL5AniPUsJI4deT7aAjQTHebZlNXDDYB
ufSzZ3+pH8CnBVtPLacq0PxLBdZFpcGPUKAjKTbqbjEWJ9UuQvlScwW/QTfw4ZEy
R8QsaPYcEzZ9qciqjWWJZ/u94lXUR5DLe2jzc0bdEx1GMVupg1Wcy6GAveKt4hhY
qsiOcVK2nj1fp8q/u5R4VrRgDWgK0P1LKWZkRhbD0IuAUk3rtiJ5Aj5ajoaOmUs4
EnFswKmX1IsYjl4QvTLJ2XVVpS9XLnOB3J3+7pQQlhYbmzN2d9oSdd03TQ+wXF+7
2aAqCWSChBlcrw3rnjaaIKIZYvQAKQ3p16J0cULM0ga8TIwrb6NdZM5DwE0zFFnQ
BgUprroyzoVNVuFpbXCEsBlwTXEC5lRjzQA1Ys3I+Eee5r6O0+IQ9eq2FXLAIv90
b4N9yBVnjLVjPTVqVm6YUrI26zj7k2U+vbhxC3y65F5rA3S/6PiuAD4RytnPyHy6
p1YK7r/tXhK46f7Yz6t7KP3zTfd1h97HZAYVw5i8DCFTRA8++OKG0brovnei7yyi
KhLALz8TRF7YPCAUPJbEGbF2Q+oauYMYxuLy3Vu71wOWAsCji8U6PzuEMuvmDHlq
wpTQVGb9mlJM0U+61Pl+shi9DkuuOA0h1gHltR7jGfFWZ4MbFTzBUTJQJs0sjS3T
llBuFUdgxzLfHAVyFDwFwcqBykBt+4BQd+4F1JtZVt6iWAepASfI9G6PECVE7y7m
pPFUUHiC70HjP9/Z3KhrOX7tdSoKACVqurCY3KPIKnI39XRg7pPc+QaOT7am+HrF
aYyY3yi4il971to+LaBUdBe6vmEJhJy7mKCYlQBH2AZeQ6OqUt+HkOjZUEDeI5FM
PAP/M9yf3jZMp+m+A8UpNvqJg46C0qPOuCsm5fWeSiDqoiwXzDA1TVi3qdfueoEE
rM7lOU7QK7S9LUmTEcBkNYlBAG5FZ1YIL6GWJjpKn5a20/pa6tnuOtl8BcoCVEKD
y7vcgUwSAuF9jKHaREk3HLYQwCB9VgeidBN9vZSDpr8xYzL0P52L7ali35YfM2rZ
N0EFoxCP4hstcy57/o54WY+a/IWW1RPeWy5QvH/56OeB1OvAhFK/50oqwtH/U2Ek
5XSAT7o/P+VjNiRhiHI7conEnGnLkxxHN3Kkv7tKaPfrEhl5+PB4qkCMR3D8VfXM
JBq6h06ZrPnknuJArD6V4iOy0O6/y5K/Tuc5rXBRMjR+RdMbyJyvpLWLSQICJS0n
cSNsCeGYOQn1fTfna2UDttlMSV5861FpYJzgpjqC8hLsoQ2El8tQD4suvxCm8xwG
5Exv3wc5XwcBu9+p1wwJQpK2fy+rzjIz63mdfXQG23ehyYso7l3l5AIZ0zW6xw3D
oLa9hwTY2kfbE6DrKuPQUDajyQSBeGp1U3Skz5CgJ4wBcPZZdfH87iKPROkz6BWj
gV2lt4AJyAHKuMvAQ38khGThkqo8kSC4Nf+PfzkE4Av2KhtKWn+CK7Nt4tkbwHvd
mphK0AP7z5ovsjGEWF/SVsTcrQ2I8Zdz1yVGOgzHPmFsq7/b2Pum7om16fSK++uw
xb0Jwjd6L1QHIsrt/aOkWU3VVRys5FZaf2acVJg6pUgp43BWjrNKBmai81+xd1zl
sPeWBth5Lvm0ysTJIfYXBQIrP2dz8P+SHh8Bi1hC9gmEYYIQ404EYP+0yrir2tqg
q/RxVyN1I6OHk4EoGuqvLIGItxaBnYDAX6m0xU50OARyR1y27AtROkWXCYnvJv5i
p+ZMp1pqVtOVy8IbFeuThZo8oYLfXsbLPlhTGpOQxaGALYNzTN+ke2gEHwVMyuTV
KM2kdz9tUEAztdQrskgRZ1pmDDK4VEsPBaUXtZPq1j49DyadTMM8JDbhwyo9eRfs
CfcgKQ7aZ+p/w10QSFs61Vmd35YDiGPFh+wtsQpjUXamqTQipelN5BjNbiy3arqg
b43xnzwjcbEx9MBaqhTVeJUPNiSIKqalv1dDfjJyy8C1U1E6g983CdAuD1qpwZGI
2Pe0gH8P/04vEB88yDpZzT+HjiPo5mTSwNODJC4NKRTdyj49a+TPvZNDwblUDs0G
rtPfWeTND/F4ZSRsgOfd7VbuoHiXuNBR84kqeQoKpvnNKYdtokYJNKpDQdNTL3zO
PJ4NF1ujfJvwNUAHykm0fwgBM5w4cHyZUmqRlh3sDmpdAld66l9948fBq+m67pzU
CmG1aQM+xFSdyClS6uxDcWtfjcXw4nI3ZMStbO9iM63XTAankUr5pd0Ymu45Ca88
VZqcHMldGQ/HMPiMVJ7Zj2vhmXgzY+PoXhk/fgrP7DCNrqlGCzRPxZFLNF4Auq1C
81jKIT37AzVnTgb+rvKDPEdBB7Jfu6RGrhFWi2veqsOt7IKc0o/wz5vdBAjS9bI0
xy7YuSm4v/FTWqokl8G/zgLixRbceIOWNEOjfDERXLrtnpQzREV75+nR4SvDx3dp
FrW/8NPE3CLPBXVQzPsDxGD3gQQXHVDJISCXykZF1+ok7+dMgfLM6tYoX0LbR/fi
n0HhG7RwVqLDhzE3xZLq60f7Q9umP8TE1hlGamJzNOmvmRNIlSrzoSUvninAcMXM
12MSdIm4orL0zXIlQVJSayT5sriu/F5Zcq8HIgmHzjE4JFf+YXbcUyUz9sVsh/BN
KbcWVifL+QJNohdjxHww4kxeOZiQnVDqDIWprC4f4+dLqS8m9chKs7O0wTiEAbrS
zR8BYvg746jFNx2/FxREhgnECSvZTStL88W9tfV6aJloyPEYec42U0i7w7dhZPAD
ME0Ef/ZMJ2FuodPBfvQalu0gV+oSinIPJcZx9WpbHGTsjkdsT0NoOhaFtSjQp3Vp
0x3uxu8mYAsAO1y5fsk9oxLh8lIcbPAC3wQ1ygBrlRRvszHHbik1bAQDJPqe/S6I
DdOqbaLTHie8seM6nBlYx6ldeh2QUF3bwfew3NF3nSwOlbbrXnjO+12oe8SGu/ln
QxsTOpZloKrqNNnGZoIxYr6NcJlolwbxKa+CDoVVHjaMFywbN9OmooEXYZ70/2o6
G7ZATyhiEa8OHRlWcW7Bc+LpwNTD62IbKDdgyi1YWZgftVK706SloKVnkTcxkKGV
HC+aPtPQs9zERtcCkAtY8zf/k/uJwgMiXnrunlGU3C8SHJmMpBVXZ2Rsr4YfW11v
oHUje0uTb3z3/apT8quaZ+S7epdLtBur+4JynsNLzXFQj1m0D1lLlNyRzsj+8nvX
3ay6Pcfm9JiWwjQGHiBqdFAk30KHg0Od0N7wflD7XuYjcR6Qt0lZ6FwvjBlcBidY
l+97JBP3tLi00qhX/SVsveTbwhufYC1MoZ5bzUG9HSdfC4grdHPDaxjh48nt6qS/
x6eaaLiz34vOL03tDBqTtdKoh8K1w0JKiIEbcCwn9cn9vIN52qAdlah1UB2fQWFK
+6gD33HlAQjMkv2qg0npjyZHeyeJdK+WVO8cdNJtphQEF0M+fn6to8LzIPBbNaT7
1OZ94WJRAX4v/Mh3t+pwQvlip/f72KJdenZmzSGxJ7zCvBPPL/40TlGIAA8q9LsA
Xj/49NjCRJEuBhTPWjeFAhfT+AmCV593FsWpo1F2v8aUapU++CgXYQg0orKvpPdw
1FDhPUJjmOLEKml6/IBwj3kxNUgQ/qFgW6cP6qynEx+pl46pis3AeUyhrN+H2ejn
nHqsSFZ2N4l7F8NgznhIy2XyZJOKzahq1Ic8i5T4DxmSRXcW7tnAh3LWhmE15On2
Pr/t2JURRM7Y0C0RGcoi7i5rHRvhUwPTEFiM1vk0H1smN6/6M/natR/medzoE5x2
CaxEnUwtMCSYKrmtOj8QURpMkf/EqeBl/cTS6vYF/jA7EG3ezQdR14kG+rS8JJlp
/Bh7R/qw2vyBgY3S+rGr0IRKgN48d0AENa1NAoTJSEu7YhV3wotWtyOQSz+ASg9Y
wlacGlPMu5tDcH0U1bBgfbsMav+vePwx1Mmchl/ccqLZl8YMq5CEAPGxJQa7HFkW
VKlwkBHoAjARQn5iNM/29t4ol795Onw+gBv+RIDRg3B1VCJ3aLFpCfGwNC9hTPFv
MYXxxwSrEr5x/svbHHpR2tryK57+0hNeDmzi5a4iUtvOWRq0Onj1yMdQmn5+WGgw
aR1esEM46q4pvKPPxKC16vIxNzlZR0CCHZWCK3mPl9YTsv0fJPR0Nw7UxZemm1gQ
IJgZzChtJgsbFmN95DhIxrgBkyA32/CKv9MeQ0xXhXv2MiclKF5aZgaW3doXehpM
JtzkI25MW/MN7v1lQfSVFJ7gwnKjfiALbzJ5C7itCvMhcFqgQAPAiUXXi/uwlM5g
zcc/DfjzdC1V+Oqp4re/HWT0eEctpVGcOR1AmlM8+idCgBAb0TFQJUHywEjbj4qK
abg68PpwdQV9Ly3e+5P+GvPRiB3lIu9wqTMOMtG7Xvrfggm0m5IBFn2J2uM8ba7v
MPWPYrUQMYiJ12z/wZb5x64oq0tatkDLNhFF3AKD/eaYuLYMjgCXYrKpnW5HOCZi
tvrLOeccZLZrBW3S/idhrZqtw/kxpN4A7pLH86Fnxy3FVzbjiDd04UoNcfQEoR/9
TjwDuJf6XKz80tPJcpHLQ6FqSfTF3zALy+MPpDjIbdrThtwyrOFHXsatNLb22hvl
IE79GNdQaeBCHxRTfq+LoWX++Qp6Was8yR/4AMckDyCiKtOW0FjEFRewQ2CNcq/M
XhzDQhXIo/74ImUDGjrkA/+ydf4t5ze8/KH+UBZq1CWCRiPqJAH8ZCkLOD2UEVnY
IhaXHruTRW804qdwZO1uf6stMWbewFEL2caS4rZ8Op6UpXgaeo1CwqnBl1tjMTHm
uBDDl1TI/QtW2jQVZAZ9USaLSuwQRIQnmUlTK8Z0ihd+2GnlWuCHYRFgOIHD89Ph
83DRWBez6ErNKR06QOC3S0wsP9Qy4qgvpy274z4saoWcl6fSJdeQ08lvuzGRc2YY
4OkzhqQGKYDSfdwIFHKXNxJk4tmB9xxqaZ33U+hZffyRYQpHsr+pcC4f68xzurcA
fd+w6cHn9tUmxHBhZgl0G22oyItRijiUsIDzCtW5cCGieh1OdMMJo9Sww9aGKamH
oPBnyVYfBVYZiLV2+bicEOu7jnz/xrFElpmka2x6+OR66asxeib8zqfktIfVfOqE
ssTvzOadp5eTyOOHXIka4lvGVVxxhdbzbe1vkT9VrRUN9NxswtGBto3FZDJXx1CD
ebbr8s+QZBywb/CUnUfztfHOR5GZN0Ov44GEcC6IPZNAyCJr04oSPThWZ3U9Z8vj
PU6NboEM6W8rPmUQH1JDy4k8sBjsrji+ZWLchn1k9Z1vspkfJB3IKcNPgxSlE/PZ
VBNW18flYhsZuFSfOD/e3rmXGJ0laBsaxHUNnxRPPOKlTRwliZ+Km4SdRhyFHhuE
BLCyL9dC70RLx/InHkgV2zuYr/+IOb56SSiUDjyvHgSqM9UfWBRUObv/AvaMlqNg
sqXy46geMcusWIzPoIFVx05EvIQrJrThq4iMlCXn9rwBL+55o7HeROvuFbOtJOcj
ElGnzVAWIbfDwAo7y/IXDwmBwKxDYn14Q7cCMufJBwwOr9Ek6ApSY2Z2LbY2kgTd
SV4PSfwJAqrrFvAAGNyzU642Q9dneHdFxy4/N0e0dILIxklQ1Jw2qZUvKmu5vkEB
TlsSHutugCUrBgB9k4TqHS8C8B3rv+0syeVXpR4q09rzoRww/1kR6QTTv9uqxTIE
G97MOUuENgn9Z0M/F1w6MYdSOMQ7yvQvC3s+hraIPOZDVAERcI5ah9TIwfgaOwUl
ZPR0bSI5eQYGebZiMOly1oj7X3P9UoIAslFxzjK/xIcE/migTrnQXAWsG7BwAkQB
XvIFvusKdmAesLvvtKNsQeo8wEE6/2NE63ZoKYcNFqIhuLqZsVCHahxZ1YMOpCdr
6ODu7zuYDcXGd4HGeddM1k13RVFfujIcpVowUbylL5iPckZjG6AX70U2sKrt+hzM
OPqEsWO4xOok1tLJb6e4z2UYCiyv/NTw6vr4LrKp1FZZ2Xlo3r8adg13oMo9R1gf
IrxgsxDaPuflS1pcu6McXNKihO/OAoTZRDh3B0szYrKdzNdHiJwiofcu5ODHXQsA
6ojXK2rNazF4N4Fsun4JUgnKZOSpZPunfJLs348Af+VDJfwiLxjBR86Q1h1DhDRH
skg0DJpYrIhRptoEIjmgE0+Cb+o8jFYNIBP6htQMGzutw3gfu5045o0i1TNDwFBz
jUL5OPCtHpOC9OECBVmuFSBbfej/qRJ8OW+KLgzYtT/PSHn3Nr1u26B9Ahv5k7zT
psNSZIgdZMQ7lI8WUUj0edVjwgg6rQ1BHONl+cIgu6mBpgU2mD+nG7XjUJuL5Rpu
julQl28WDvOuw33FMa3QJfZbpsSj416gWUWlDSFM3nHlKwE8wg6YBx2vaKrsOofL
srKlcpFgPqBw0gPFnu2HIri1IndZFx8CQvH/wOgTaMbkIVIMfo5Nhr6T4xM8enzB
czW89hTn4renVw532/l3xTODGO6/ESayuwjnejHJHoMsOozoNGahKulJ6bEgf85D
/vti0K66uhtiS6dYukgS0rsjx7Tj9M/meHVdhe5MUjrDSsIgfxEKDoVpZjshIj9z
1ba9/p+mq6jm58BSREkNu057ZRHIxBIsHp5C6OR+2ZnwYDWMuTmUHjXVBildSUz8
3/VAi1eC8SQLHE+gRF4p/w4CfSKefuOr6zRuassrPFu0u+RyVMT/1SJka/IHYS4z
KYUvLkLdBHMvnItSUlE1m97BY2bcaHjYgTeA6OkKPvYwJZxcJ86B+vWjYXcSUYC/
oKCkMbwtAqd0qljrh76PMYvUgqT0VFVyD581de5M5xpMn0dtqfKzC//p1oFX3SYV
hfMUq6hUEPFu8rnw9uiTATTC1+zWrWiLc77I35Ccxr1havLfQbW0WrQc5NHPdiU1
JHb0AegYnQUIX56yX05LpdVBJCfkvhbciNhmBIx9ArY2k63sxPChcYce5Ln3+dal
2utTV0Ri4aIPsDUW6vF9sYqsE8Lja+8Ow4Ye2x0lr4O2LjzivCPekPJmr4Do3Q2d
Le0CHuqYS4gw26SncYbCCFmv7kQxBocoto7OhM3kKQ3Zwndw3eTklQ9t8Wt4CPMo
qwCBgsUplMor2i4YKx3DVrVE3EgIYVjBQYwlsjCfgU5u8tinBdDdN+uIU/x7PBeN
Zsf/a1Ev1vyRjdZjYMHjGnhgKd7A2oyZJW0k46eh2dVic8DCvBzlhb/yqhmVvtaW
308i9V0CAO18kTBSv8UofMjb4VXu8LbJl7TN/ERNNqw1YF3hWFFCQxlyKhBb1/2U
mnjWoh/Xn0qdyO1DYzCaqR6dSlRrdTuME9WNbpU79XSsY7BwiHSmLfv4dSJit/h+
BOMMM/2UH8NMjwQmlllGEAiGiAcK3nfGNDohy3oG9r8c6XHAceGAoOrPIplKcHX2
ntipYuUVhmbBvok5Q83rbaaHSkIstS8NHf2iasTvU8WRfRApetW77LQLkxxQdE27
7qEqL2/xAPJblszHqlXhmZ9kTy/BX/oBml6UxpZAz44x7F3AS2SK5K3lLlwm2s//
jPsRUlGaprnxYFGC6EiFNMvSRJeFBfv2hsbYs6cVlhD7hHJVl9vzdPxz6s2+IgC4
DjHA5K137JTDcNP7WykkTmzj9Y+HVBzJ6yRtzR7WxNNyi8+mzFt5cnCBt4lD+qne
zHX9SCkjFb8kRKt28opAfLlFq1ESD+/5W80SM2spXPz2wCAW7QvfjfE87Xxpl1iU
vWLXuZfOflGdRnqmjy7G1uY9c9o2LBn2LHVh3zy4Sjif/UYtiJvu60GnnT5AAU18
8t34vNDgdPaBVOBq+pHAoEkxSrxXU/cTsJ1BNaght0960S3cVfKiLRZRyiJ/EvCT
eSdr7Vp+atFY/UwRdUvl7Hg1ZBEYB3xpQW5tl3tkDvq+wzJM2+6mpio0qUwpQehh
UCGLHnEw/1VxOVt6lnNOfETXH60966UVBbjxK/ziHMV4b1mY4AYHaeUFG2mBXUHX
0PtrIRoKU09Rh7e8y6dEKJvzeiBpN0BC6syXDrS1dsLV6hQgqaJvKMO6zKVtnTaH
wPZ1Hgxh1WLmiI9DWnpvaEJOojapPv0JfcnJ76XHmbGgkGww48RQt0N/nFnirNmX
PrTW1i1HiXN5K3hAx1VM6YSrIiWrOH8CIq6+q1+1rlyBBNbyBrAkuKu7z7e8N6Ai
1EW3bIiICB0UzUu7Ly5LcR9hbzCsumvcghSQ7/In08HmE1al9Pv6olkUtTaOnSpV
AO1hcok7GUs4rMeJo/Mcb9U1AZhPfjj+bh97ZnXy4H1UvYpEBLoIzVNIz5Uc8Z0b
CwaFLPJty8XBvXrB0gfpeKRtgRkME0Ctb1H7zdT45CFnqZBRD+iy8A8uua0S88IX
y8IusjZfjBtnxRF13zJntZeBQD8ZIusSKyI3GblZ3M3kL9z4xcFc6GpNc45ux3Hu
YODeo4arLLTxl+tPtzDeBUHMvA5LY6OG5Jn5XH6MM9QRsb09ffQPq8ILF6nE7WyE
s3fR8RBUgCiF80GmbodCKQ+JrOMb1tDtJNVmcT9t2H5J3vy7ajrWHtUx5v23PgoL
AnQMXdQNKMsJbChEElbM87FGpFoTnEgaCu2zpE0SMW97wv7AGCCwoJowuYva7Szw
jcIzWhvlrU4YovRpxF1lEdHPkJpCQ/cVdtJPtzQqm6l9WC1wNYg+bbWYZ/9RB6xy
XQFQwBBNYymo2Yd9S2OreXAqo8mKi4PisxgtFILqnCWt7MEU9TyrX2jmUIO0xS+b
sYyxLBKkgDgV+wXrgrAMg4ZRubHPt4TVXrCttHcCkB6P/wgz7yeC1CYVSvEWnVqU
ENmwWTuUoWpze3SuArN2JfAuWBanqlzqUyc0YrkXpB3PXCAU/AIvKjueCYnML6Yq
GVPYkfE+j424K/HykUPaA78AlBEIaXTatxoU8k//wGf8iMg9IE+AxYFIRD1ms5lT
awck1gXXwVLVXT6wiukvb4KYWcThtYEAhBBi8xloc1qLZkSEZlwZPh5dI6ITvPyR
myi/HXLKmdJlCc6tBe4yWFvibpznZq3ffAeCu1C6ZdAOueh3t5COJQhXmAHD0Nd7
wr737TgP6YChNcyPp+OUx6edWd3CWybywfAbnE53WMaQIxPwkrXbazk9y7qmluX6
u3tO8nYo8n4Lfw4VBP2tYPMXRC5ln3J3kgBdv7/hz8IglmoBD8rhKGIWIbVrs7Jk
FR5/LhvUfciqLL9bcrDZ58/RsD7X8ioSatfGAvk6zPhQ/s5TLdmfH/PEMOyeKGll
GEdtUCH63RhCwFBYSZnRKYWt7HwD8k00zIuhUPnpI326UVMEph9Be63Np6l1oMd0
AbEU0CLryNrRwnd0W4JfO3AWxoQt5AYXs4VkLtoTRzx5+azsYF7HH9JDyrezC/Fk
Yxo2bnBb3gvajoFDNjY+/p1yResMjUtGf7t6CcpN/kDrXkRO2bgFN2JOBMbGbthM
Ys9cekEPkp0uc2NmnJZYgaOc7yoeX8stvxCr6gPD1onB6WrApJVxhN+llq4s7UI9
4TFSz6gJyf3QSWvnJoEncpy2r9rPaLQxm2dhGcR394b/2OcqYgnTw06IpmzMysEK
EsKKLSLj6YjgB/aHLiYBDR72zVjwwIU9vO8ZOLYYFtIPhjwdJcp5wnk4iGpq3l8x
pQPpcPlCAkCKiMVn0tCpsgqVUpaA4ubJeBxaVrJME4rTtSeZvWVuSx67RCcX/Q3y
QVHAm0HQGPDXBQ7fZ/want5Q0KyY6kTNDe0jEtMdpBbeZu49mZEi0Ww+N3Wwh+Ce
I09CLzZO5QzAnwrPhqdsFmpqJfDcrDq4uKN7K3z0gNwCW7UbZ4T0yxLXS0XSvBk0
4QUo58CNEGlu71H7HiZdls6iSwN5hEY7Syg3ZrdoqN6tmrtPhcSfg4v7xTow4bLw
RSVEgBPLMxQFW8+ZsWF4M0Fr8tgn9Pwizs+8y1Zk8YCXq6fL2b1dbYQkGpYpx8i5
j9p3lhenY+USl5HY3EMCphRYNDbnRpv1NTSjskZhPWsU8gQc4ZuNHn1QqGuBIR/r
I6ZeDlk16Wkv6e8fL9ojQ+BQsS7DaRh7OtpsLXrpf0L4RF/YUry87BAU8ZpXOHWn
dyyXefwfYVMqYPmKOjGgevObrGReGDqwWW0n3sh7RInLDg8k60w9RqZhXXdniyZR
VDmMiplEPZCA4bIV5rgA048kxooPk78lWY/ArsIUaFcz2psOXnqA5BTET5XR1Mhl
8FHgLYgawDPwSj73eAcuIVdYa/20UeGqtnLwS1R7in9t4qenfP+R92JnXsu/OSVC
w+EjPK3hEpTcNgY2bovduPnqIAefjk/wMOdZDYQ83omqeWfEmHmx96ue9AT/jkQu
1fE8bHPuKNISOwYutrnUipa5fMA/rKsJVcDnqtI5Yt0DNsYMdk3OJ/8s9NxN2enZ
9ofd7Z9SAdh6V1zSgv/zcGJlTrOM27ALheIGMCA4D4MReFx8VY9e05YOr1spnhZm
BKYVMW/QphQbcqfxPj2tHA/ZxNtp7ErWIRRsd3hTT+y0KwaTTOqQgUWQnetUVG1M
W2VnDhIi2BOCqx35+ZKMmOpNdxeZPHSZ2PYlNbJlptj+GjdwB9QbxQt0bbfjucUY
yODzO0Oxu8/VV+lU/lyZbLGaRv79dvVDXj48dyBpraTAh2oHBAgWBVYgsVIZhtgI
rNXvqIxBElbpqUA6FJEPe6fNHYVK50bt17JGMOixj64ktHE7OH1AHc+7KYbnAXT8
ZMqS1jEzNsjcSi6fbUP+Dt7DpCNrrzyynGuxW8Yt97+b4mxQFgMTEMQ4Q5z+W12g
b3N6i6QdwO1hyGRfeZkzRCuAo8lD9Hbl20dQi/Th7afBPDyAtHnXQUUSN0sEsvui
zzA2KWNmAIrbRl8uGjn1urIX5yvrLkxEZ3dB/1T69CQu3YpaXYtCov96qWMTzOQw
FWnAN0FjQyJKr6cYXLei6vJXUQ+jtz+clePfxMwzKN9DrzIurpCmO1QtQPXLdfRL
YyKqaUR2kDnbYdim6/RG7ZUoNG+Ks24ObqpwKK8H3cs7Wp/kreBUf4ECsBoss/vd
CxcmLUBKZT0+w7GI23nz/eGHMDFX9fE3nNGKstxgAYgFwxcGYN+zCkat/+tqQMgk
MnEwpxv9Zae+q/0kvSfi5GyUMRXrORjz8hdwaqffq0+CxYFuSRweSgC8Wb7B3e23
PDafGCgzzMhZJlXb+C9DbXiYyPUNHZ1HaNCc0ZnNqaBRvw7WJp0RuYOCfBkkcXiZ
z/wTCksXpl1u8C0NwDHvgc5TyO5FrqzCym9buVuOQuoBhhhFG/3JcZVFFmcixqdf
1jERRXjqUA/XbnHQKwgW7GlYeNmasxb8df2gTShvFOsCILjwT5edEpxIB9Ca7dOg
Fh3OBwyrJ083neGhDhxlSV+NeGlUVX0MksGhyzXky/274amu0/YEoL8b+2rgGtBW
VHgghUQGY5QrggIXBU96Cf5ZU02RRuS2KV2/wKeDqWbaD+T+fKIykXjWpN7psITM
G49hYRzliCInyOcjzEkAWjZP+Y7oNsVoSCpi5JbRWKrx2rG3fIaKvUrlzVv3eOt4
MUwhXDQkHOdXD7cPl30tTPEjQnBFkCInshyhe7inkjB5hDg7GJ8N01BrF2ZfP1DN
USSKS2Q76e3Cq2G8DE3TO/yDJFe1KPGCnASScuG/c5eTQrpz1/6gzBv/2dE85nxs
AN/Ar/Jee2WEUCKAy+J+Eob1DFY4W1EgEXDWvwj/Mgb1piWNDCV8Nw6RWIbqjLWI
cBFhCXr+EYhuMkagqZs708peXZoFc0lBRx1TGZ9s21nkgg3QEcuXLV1vr6QqcP8i
F2/wmJvETaRXpXo1S2jmcr59927Eke/xwvfADGOestbqtGzztd6dkHy9gHhynFS+
w732HVYtfL7KrwucMgVV1a7bGYcwlHjQh4JbHMyr1AYBp/W69tEyuhoy5i6mRPVv
IEEwa9KFem7iE5zIeihVYlrkOCt9vPJMhgh2cZ5Xvi+j1X02J0jXMp/b/9skwiOD
9jjU6mNi2kv4vdHl4IzIPXPpr1h7O5uOcZXMw32W+rW9dJ3s0fSRrurLlY4xm7AE
hE0BqI9/cinwMClD44Vf7RUV5PCrYbPtPuUZ1OZjbjzY6NNgq5/+wPIGSbTYjN3J
DDjDeTQ4cm2wdfC/3lROKT49+zz7TCWvnqZmcJlke15KL0x1n3rKht4hCpqRSPz5
/yesGhR850VznfT4VqXG42+QAFpUp3BzUshNgiDAESPzt29Wo+6cYMNoBP9whWji
6lLOe+9YxwbLQQOWfNgrVTtmJS01LCTEb1aBNN4wxm+acsYS8qFd9EZgMgRcmkzK
ogdy7JMr7/MaNIAjC2zM+RO5wNNK89kBgWc6SazPXNYf/TxQHadf6HKy1sXKwBxP
NUvcnO1MzeF+LlyOrE00L6aj+d71Hzpd2o4alv/+wQceYVKWEDCARkAskl3ZVxhb
Y5V5vTJWLubcvUaZ0Hw4TBe+berXhE0NiUBflFHqfaKalXekLIjZp5M1g8cIbhYl
Xo7P3B0Y48AlXfDPmvn+TSltH3A8q7jrOw58qnWBzD/oGqlTTmPPz0xrB/mFdX5m
bU9uAZLTMvoTWu7Bkk7J8uih9ee95bOU+sStsC3CvkBk5zpC5pi4CvyQ/QlrmsTD
C3+2ylgZxmzwzlszqTc2uBVp931uFIkf2blIG67RVdFMSXcysSiOIq56IzO6fZNq
Xf4V4JfH+QQvOchp1iIhXQTOah9Fqml1/SOqHez9muYZmkQMkxJU/flZ27etEimf
M376IyUuanyn/dWxGhtHJcfsH8w/Ir226B1siY3kVN2h4sfr0gzeNTbgUZ52nBgW
oLkCik2V5oWJeg48EFAS+w7b4uQmnBIMLAeB+cKcb8jM1P+6dMmjc8jtZWOFkyCN
ex6UiQZSBn6dgNwcwtQFubx6HWr8wW1fZiwCT5vymaG5EO19yPBTnB5Lw0gMj5UV
B59BKSUxystr4CAZ98HSqLgZKUVrO5N3oayFkkFLCpZ8HhsOjnV3y3eYKxR+dRR9
KkPIZhTfokCnH1yHo76J5W/U1kZxkj2G7J0ZLl7Exk8Vj79BOH2ETBHGINLSZH7a
YERf2cYYu7O+KV5baLp366lul2Aj+5fnXUUXiJJG9NxhpnqludO56gFEOE4q4L4e
D2kS3upI3jN0GNCuAuGNXO6K/lQz0+PhsP0wryPrf9Mw/v7eOC3XFA43/e46+L2x
2SRxOmqaChcL+Uwpefy8dTvyuXC0hIVAGuQKlwV1MhFJNBGQ6bm8xao5apo/6cZG
BA6m7qm0R9+J8N4Fy2PubezNakIVcTYhACQ0P1G4oH1f9ymek6j0khRJQzq+tCh0
H6Y3nbeyL+eoLgqgWvu05DLzMRTUZG5dL3Y9FsoJZtIWbELzSth0SKCMD5PfUxye
B6Tn4pL5CLNMLx8ibua39pcEHpOq8LsCAq5w2LIfmKvmJhryFzvU3ExZhF1Wl+7L
kds3CkkQsQvbe/XDxusmIfS3ToRlbFzp+98q5x2JCuToU2T2dN9skLnRi4wfG8bU
iTM/vDhOBR9+H6FLI960dQw+3ewjj086ZqsJNnIr553763jMNj1BJnvuRqCNNSVd
hAXICiSCrzodSU8mwuFnzzkpxBHmUP9bq+Oh6GwQ+pGq8IylMXgMdGxz4bHXTTqq
wdN3Jzo5qrgjY50now4HcpUhicWrSpOY2VioJKEW3DoadvSg8nYUfw7lQcvZVWgy
jAjVjKlYR0eyRWxfSaMh1CpM+w0PxVYiNW1v+IUb2LUbmyTU3DmLYkoOA6igNdKx
FE96bGgoJuWLiJuy7TKhWRC7EwtacoC9GEAm72FCXpJsx68aMUwGJRN6EA1JlMRF
1ggF2mReSe663FZhtI72aYXhittVI5hA+PDKTC84f6wLXpw6khsn04c49oKq06+3
gbez7AcD68afifhbULhj3G0JsXDiweNVIpLRjtzhESPzv6R11XtnI+avl4Mj0TaU
bTSWoJhzoa/BQqyKfzbeqx20p+9maBf9Fv9lsMt41m2SjT3OclpMmCf9BRc0IrGC
BT8nQjX9NNNpz8GhTpY9GE+4sVWN4wMeZC5mYvo030h5AqldpsIQCQCRZeUMkz3B
034SRKj846M/y1Na6U27d1e3KBHa6H92l59V0/v6YWZUOfDt6B6v2AoLAseJnnTA
Q/XfbRBZTJLJ9UNvpM8AbKkq08zYxQzrXiZW77Lx72unTbHbLSbRj1VQzwdUGABL
CQdWvJdeygc2PsFG7hHAIIpPxtT2A8bQ6vQfpwRsIJrIATkNikg0f8hDfjTOWM/X
bNmkul1zpx2oaGtdHCxuxe6gbohXOwYyKUXvZIX3xFa3opzZ6rdmZvyDfGmZksnQ
5Xc3HdVwrFL6CvreA+NKtPLa00WeGc6FVuFP0CtPZea8LdOSmsKQO4I0+VMmEb7t
QJ1Yapbwi8ziSRmKEDzFETGxloGv6QWLLfErvmo91vZf28wMP1s1MWO83ubtUNVr
lEvCFPfSYDCpWQORH+nOacbRFfezGZkHpz30kH7LFaLIo4PF/ueD6VXhc9iLK1YD
8vCjal0TFJkS9KN2egzdFK1xCwWNWVo2Y/E2coPOgcTW8rusQ6AlLGGsZoSFyEQv
FMvBLKoXrq+JAdKC9+gwJ1VQfAM14riwxrTD3roj+HlFsi4NftS9WH6NzyNNUKRG
qCyNaLT2Aef81IiczZvhTNpwwzYHMUKiCccb9AcWjfjoH7oGIqAEp3+Hq9whXgJT
0lcZSRjdGqKCb7dgQFWUT0B+A957gIb9IF6NGYAJeqFufY4T6QJGWiCcgw11+or2
/NUq+TYx54v1xAsukeTlbXvqTAhIBps2dgRo9iQrNwtS9iqaRfzSVHM3xkfH4cgM
vPM+QvGttchPqHhxFWDAzk8XVH5K75qS5sfF48IBLdxGcUhlsPs6mDXiNr2kkfws
MPwidUruA6uwrKBJzT6CJDG3dJxNQEUavLUJMe2vG9YRYX4QWwQ0m/fkk3n+mIT9
KFfy+MAZkiKj+EhvlKXM3UsnaveSOIBqTtubuBMnxkipOdWSQXLJlQkaXqj0aSe5
6SbJmBs8NHymaCs8r2SVJZDz4LVIsIQKCQWfKW+sYOwgg9ypNsUKDNKeYZsVlsxm
yIBoia+n2+V8osuAujZ7Ca8Rh/oLpNGUeqWa/jJ0p7WweELdHHPSj8HV3qHzSuih
3gu5HCTuNOGuQJbqvf09pCcnv94I93pMXx4x2yn+EWX4LlmX2hASif6QW0QJIqmV
sEzqtZmRhajntmU5EMA328alGeQVOjV0EYUxOfVRyFoztNCqZQm/sUX8r6wC0JLi
f3FzsDykly0aotpeGXDoEDOhgIhgM773+udC6gyKnrHrbcc3IMDexBxUktMDHPGj
AwQnJXWelmAiVviJv4Fla6eyHsbFP09sBoeHmezyNGhXTPRzixtbBwgxAilcBxHO
4Q8h0JVwZAa2BEIW1XsdxLByn8WVjbK+BiV5bwci9xDDhghvyNZY7AoAbgwKufaG
BtjwK8pWuHzLPrZ2zPeU3af4D77+5fZ6RGBH2pQGm13Wo2WbcI4HjQ8jbQLtw+ey
zm3kL08WRues++APK1moF8gfEkceC9ZnSIe4VNT7glnIzSl77I6wPrBKNrOeLQ3I
fh93y0FNCIOT+pFNepaJ0hjHbzPXmIuCjhgCuC5xwnpLWDEv8FKfBw/P9p+cLLmt
HWT4HkYLAtA9znuXciXT9rWHqCp1NrxAO+E+S/r6iTFJtsv+LLTKMPYyyV4Ekb1C
+WWvrglYnqmuz4Sz1zpww5NozBQ5gCJbOvq213PbHy8v4IsQ+PV42SX5Z76oygej
mdbUEo2YpGqX3hLo7hh31KkAH49dd6HxePnvc+PkrJuJBucgy5SM1qRV9EsFUxCX
ePyEIhIY8YhY8rQKLj/ZZ0bc/Vwb3GOMEOZCJlVVb6antcsgywrktLY5RzrpNRZs
b77nCinFpbba7u/fx0DeDGP91VlqZwAXyEP7BvhIcqIJS8I4vSXAx3zx64rme1sd
BGhbgQlOWKSojru8hAvh3AsfjmNXWcU+UEknCDjV5TMGAdPk/jG9tIjLdrGexW61
lRf8U59jZm9ZGVIYBgNbKcd8NUrimOx2wMsV5rqt+Scv2292ioA0TxCgX1v7vqZF
XrVsh53PLp1IEmGmaFLyKO8t82tSOx9xII6ceH6Ht685ABboB0C5RPW5a7I+83ek
o1b/WI3hO+umu09x0OvepWtcNu6mhm+kfXwyGYjN8IveVvWc3kjBx6lUL+xnIgKn
DhQFMQn0+k9bBOAwleAYuZg+UzZvejjT/Tre5wpiwqqoCveiPggT32hFcGzjGMM0
8T0aYRnsl/3K78pI/R5riPEbmpv1uAo3qVXNGujw6gKVqkh+Twg/AMteF4wr5Hbe
kvwCr0BK7SyQPZwt6GigXfqmrjN/+bE3fdcY2iA/uRUS9nj+1Vg4uADnLLdvlpIz
b6XTBSIgQ14kDKx2d+wC7G3mmFuZ+9chQXtmt4Zl5RxFwpxS0EcEjL9IUAhUP/Mu
ARsUNlZmatxiFcenfA628uvf+DYtHaglOFnygl1j5OHLsyzbroamv7vqVf/FjC/R
sNQuhH+9on04f0OjUtLosFTgj4wJUZut058AiBl20+AYtLZhhUxRhKz2lp5CNSRc
GtXytWQzg+acwz0W7xstL1BhElZVZKLi83wsXf1rIQ6/FKnbYOIqQBiLeu/Irsvv
KV+B6pTFExLL3e2vkj5pfAeAw+9keASVQpkz1vg0X5gNWyCUUkFJ3ejtrSasE00d
Lu1IHjwLcd6YEyHgxHjlspSy0QJ+bxjM0YBtru3MQE51TURiT+TsQy59qo6yWhM1
nFVA5PEty7v7YVsq5tpupbMrryZMpcOvJ1tIOWlXfLo/+4s2wzrHYzbpxjTKD9p5
2/+skK6af3rcjAx21POlT1ndUrKTZsD9BbtRKKvbw7rI3N/NgIxsv6PygX72wmer
1XjpXu8I4Eg/kh1xe7nO8mLRzAZ56k/YjsS6UmFYxZWgWWi3ZNpApRASZOx79Opz
0CFfPb6d1ZBEDgzFIZEY6nzQqL4YKsNO03SGoaWMim8Ee/WOmQxadj6iR2sFx8j/
8Gezz4FW5ktmYTK2+saqqfse2Ji/w9rgbtrbNQ226046ZDaOYJJ3d2vOZN0Eq8mM
GVxxi3oSHdeuGbkPRqT50OLz8TCPLYdH2iTMDHaywFo4TqDQZDRM1ACezILbV7uT
OVRwv0mCNQDbkq8jdqHId1BtrxkxN+/WU0QjF0kHmjEUrBQgWwKBVC7ZB9ARY2cc
2KH2hutwuUvNpN96iHwA/n00C2tPatMhBB+lgMlwl+4R3egrejjhN/7DDsuS4ouM
sriE7DGevRfmPIhwCqEcoYkr6FxYIWhAHJq94igKf8ne+OKc3xbxomsfj+MG0Pjw
6OiULJWnR5GicCoDjI1H2SgKj1lZQ6kadpHUlUUNciFvBqq6c6o/94LbmRTw4Jsf
YuNiZOFrdaK/Jcntvq5sQCNWwzhyUhjWQGDoiahl7N0qNA+WwR7rHzgQ49kUK7lQ
GmBQNfc2FMa1aXwW6USQ0IA5CAv9UPGQid3kj68AwZxxPLyGe1MCn5nQlJwTHW/a
ozn9REpo8a7Y4oLPEKZcRChgIqBbFn/GoCsPAxEZ92r8KbC9yEKepmMTIy2npsJq
+Yry3/dNh+l2JkvtB7y5zDPPvRGY5LSpThnCkGkV/ulzy1HT2FY5ts0OO3/AfGxi
D0VCEGmf+/kYJnbHwBld8K4PTvThWH2BluU1eDRlz/dcWzERBSZxXDZmxyZ7oOhm
9+JYSmoPYDVh4gN0I0iDhUQjJbbb7+0Vvd+GvvHEbrD6qrNQP6AYII6vIpAEpJlI
GtVxilqX7r5uim3afa5sKNZo0xBNKoOcG8gzXhQaTYlezMNCvYxjTovVVF1k6bde
y5s2ypya9J65rwE7ZcC4C8xTuwnMWRhGeKwYa4oGKC7TiUZk5f2RCl7p+cHilnj1
Lbp/8nK6pPggTSVaUOcLAL8aB67VpwLV7Rg6lkduOv0PY/LPqEeaubtXlptXX4r5
vewxpABQ9ovCLrmx8p75vpPuJzJ56Yf2gNClpUYNu4K8VwYl3ODDL32OliPThFIi
C70yqNQeBIOvuk5cawimtZDq6GSZZX/e0e2BNHTATLeO0pqKpbtGokaCVPyCZ/hN
gt5n/OjgbRLEC8KhtOaeooGL9yWCR0ZDdwLfVU/7BsnH/KMHVcWi4KjwMIM802FJ
FHZEfzAVK4OeGZZaG8+8epb8eR/o8n6gRa2sGt4uwcsKxfMe55m/Zw7V2TH29Qt9
XJds0QbURoHYdYzCOAUqM5iCko36ERA2ZC5YHZD19KuklTwunTQMUC45jr/KZYlR
q5zIUA6Q5LnLDGYKiLtQHA+JshNLMlyZeE2BtyjpY3RF4MY8UC5WKMW5sJmvxsU/
fL8knDXxNTD5fL+DnKLRf6tjVM0qiMD4X6K52nnhE4u7eMIf1AnCDcTyu8GRFYu9
TJQcg8Paa1Dby+DH5Us/HefkOr4xqI14NJlbB/nZrGq85xGMMQK3eQFbUv+hhz10
3W3xFxaKwU0xsBZsOTG0/q6jLSCrj03NCd193NdtNYHJ5z9YKgytAqeFpDXXjq7O
x+J7B3WjqG1v1KNHjw30Cytlsbv6fe/+T4jRWK3x/EGBrhBUOm1t0fVSRMkLOHjQ
pCKflT11sV2z7dsW0TyqQkhxe6Zf2yI3q3wE/ZHmopC8pg4Xb8/PZ1qFA8H1a/hT
MEH4pW9gYrYzeI8/kLu6trRgQ7uss6CMsR6zEOcpnzOdn+tjQgijkdhAZ3zEfPyE
8pcQwhAy9kOeSUCORWMaB8T3gNkCYpPcxfgCx85eqBHq3c3jWfyox+aZ7gX56u1Z
yEUvZN/qUAiqxx9IrhPjADxy2l0iCEaanIFMnypD9/YKxgjPPplNtMN6Je+2x8Ei
pU1g/LjLJ/7PSX2rSp3A9Ble4ePDIMe5L4OICKB15hpjHMMA+0Yev/syT/X4AJx5
bnml02YgUOM2i5qOZz9+2JeqzU/FeewKfHW4yyRr+PwLGEhNKjY7QzjhZK4MNyJb
7yc+EApR1UuEEeHQCT+5/K47AWx7j4y1sUDyap2n5SZNqvxJtmGsg4E45ySyrCh4
s/wjne8eAbwfoc5ya180Jykb6Mrer0EtUVUA0ImuxxciY8QBUJotz7zoGr+0c1KS
WeI17NSUfWbz1gqlHtXgUAiWeKV8L6QD3NAMVkchGvYLpLygMJQhYbzChviVk5Zh
fgPG6noMAMtCj5MlNIayAWt0HxveGkV26taYJbv8FkX53teoxX7tP7wgJn+FXwDA
Op1Qjh843A8nQIJ8w4wol7Iyx0P5KE8uy+h50yDvkuAnhL5QwC7bvXldchkGbelJ
1SvzmyKSTRz0w6eMISG2U6lhlkTOynylzgWbf/b0dUR+llKpixY5vYVfVtbPshfe
JJz+cctTP9A2on7z/23Y7a6zkwSetTmggA4xaUaD8UiI8i8nMnSi4dmOc6xO1eMA
B7zwimBWBa1ixvz3kC/uQJ25p0etTEHUzVeRDqxIzH8785pwlItLmUb/5apjEe5X
HP15MMDYjaHwvs67+vEQk+r6IZwjVmjI0qRRyxmqy2N9GhycsSk0aG4kicLXcua1
0Wp82QSP2njCYHASkHkl5EdAMZK3Cal2ttPPvCffEGcMh7d2/D0XUD1zh9qR6V5T
V2adrZ9sGA/0kzInLpmoS24SZBh2qFGInlEcW0J4XwZpkQ+Fe34Q9hGE9RB4hAbH
WvRIorW8T7p8uzmIPKA7xR69bJC6pgElDnUPu5nIbBqqN5NuLEx1U4rqsYSkH11F
XxlYv9vAERc3jQmRrK9efLh++KAGu4ZbmQfV291zYZMPNwAaZp7Mpn07HSr4+Opf
sasQtuj26/bk8O+8uxj0/2KYshn+y4CXKT8d8NMZMFdlNsXbXKtsUxf3NVCFA/7o
jyq2sGFh6owmNOwBtlBTI+TeTpZo1ZpDT4qEg3YG+PHQtFxraXzgicYi/+8bsr3M
dDdqwHtQxO9oShvDAt8kzLNmt78v1rISB/cfYLBPfOvQ2XGYVZftzif9yxcPE50w
j1w3PsIYK0I3RPh99aqg7HlX3A3kclBw68WHf/GLl62K1O4UY+PdAxjODe3lFhwp
uXbQx5t0ZZPHBssUEWnqyhlsr9MwpD4Q8O/4TR6gxRb+KOIpyfPG7vkpxohP43By
JwgitcmPrhkv4c9ujxf7O+jF7yFffpVHxpGv9tM7Q2WPdlUOSO7MmrN316I/2bCr
BQiWJxCPm1lRMhllzdlF0vYryYyPT/rZf8gjXkcego4l+1nxE5PZUTm9CUMQ3Whe
J9XBki6LF0WCzHdmWDikTd1i+XGg5IWnoCKDePbVWsTL+B7i18LX4YpEgZ9H+UFy
BPb32WMWDmHn/pXwR6Cd6U5QZECVsXszRpGIyuLAMHm/m4PdMj4oESfX/wArKmZK
MPzUkYctLerWsw7BgovhSAuQTp9ctG1E6rVDAAj+RHrn0QR/vIXp1J9x4l8mPBZq
GJfsDYAQYGWIHNjNWrpCgV1re4cogARo8HTAmy3LWRxDdDsqu1uQBAGeya/+wSlt
0TTjz3UH04YfCvWUAV0xryjhwlG/HkcMurP0M+wXPTurmXNHpPEDutSjh6qJ+MdH
I2vXJxQ8Amp1mQg8gaIpOLkJxiKkqBIaFuwd0cytjES4quz+30T/v8yN73vWiLeT
+M7ITuF5pWPjnugVgZv9D1/GRh1pNn3m2GIYpdp8TBa9ZnrV+aWyBYP8tkDv5q/G
7vkc+7wdpSr2qRjLZArqJ/PInvI9MS/HOTmp4Fk+XZtqhsHtZHmtrdi2gtwHQYRW
pR3q9ZlVN3DKjKuOxBiroycQ5OZKWZPItstHG4y7ESNNfRwyuTiy8TNs77IqYZVR
/YNyDfUrGEbBS/PlGcEH5yJh10+kEkJ1syn1zakUP1GbETGerwzoyNmua3Fd9Nt5
+98geNLZ5dFD5RLFUPk/cMB7gv351paW7DTYLqCC9k945uA3eQKvjfrnCfa9F0qg
CwUPmedLHL8jPYnpsdoIWkF29JbkslQ+p9/KPDH31joJAL1w72rqDsN5EewKEEfQ
yQGOZSErOwIUHYEAhgaNoyBfVCFrE9fHlFxSK7vsc21Q7sdF4DSw07NQC33Js54O
J1TkCuvyEOVhHAdqE62HnCj1ZU/+Z7l/9EEhGpYyxAbF/O8v+BRrVZK0w+z2Rh3X
/leaYEnfspH20gVb9EiFIcIvUvCDUUJw37RHM5fQlz9AYPaMq+en7WRJoKb7+Y+7
Fk6XeP5YQj/50GHURb/vjHkd+oO8KqKgDtilAc6XmNa73TqV4MiScXR6Opv2Sb4F
ffQHsWiEKu+zWP7lcF7Vem4kLHjYABwYRp1k/riUTvXIxKaMW25hAcGo1lPUUP81
/jNHg5uyu1re0z1QzjEyaUateUQzYuP42hYHc1grlDgkzAAKIxl0mPAEYfjVaEU6
F0C2dg83EQHzlDAgZD951RwwTfW+96BCQtEgMNKOe52115/+U9mp6dT2KS0z7rjP
ZOVyFkjwII4W1Vhskm4Qy/ubhapvDf9Kyrac/pP4yyFRd5nfFFDaJgQYyZAUCr2C
WNim4Pn9Uh1eJ8dC8leqo6+N0ZDTnEKB37UgyT51kZxBH/OQ/Kg8Yqrn7Z1UMgyw
nwhskJSlRQ2uSC2ul4BBgvQEb1lQOG0/st00FtPWYi9A+6GEKv0x9pT5/506N8sv
L1WipsuaoBlqlJbpt1kgQzITaG/C3FhFPnkJ1gDQt6qMzOdI390wjEuzxwTziYv0
FTzeDZ92Hl8kbvDrtAyVhNVRy3h8J76YudWtJgja328KOtEslXTMbtiS2nos/feI
TV6ouPJTmA34lZBbIWRSsbufsEsm4gQeYppZ71UU1QhsKcQuiNI/y6dYVwnX3qbv
45IkBIcWWQegPWBo3Q69Dvi1/fqapGr5OpszGCqK11pPWL1ipJ/X2yYH9BaP5FK9
fsg9xscQdf/9HLAG9paJN5/eA/oP5gl3Bk1pTgLbGK+t7MDQQPZes1VJBxemmkXx
DlDQmQLYWA1Cr7GGg7cSevHNb78uI6WkEaRMzmRBQ1rIjCMNKJ07l5HBhPJDch2s
MbT/TmubDH0dwgdeq3L7GcPkG4S+HefLM6pBkgY1O7y5eRrrUFir2FNh4J4SqsXn
JIyUnTK9AvgiPO1l3kW5hYNZ5OETc2kNMv98dnw/yy8+x519iLQWdjmTJeGWZ/4G
`pragma protect end_protected


`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_slave_transaction", svt_axi_port_configuration port_cfg_handle = null);

`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_slave_transaction", svt_axi_port_configuration port_cfg_handle = null);

`else
 `svt_vmm_data_new(svt_axi_slave_transaction)
  extern function new (vmm_log log = null, svt_axi_port_configuration port_cfg_handle = null);
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
  `svt_data_member_begin(svt_axi_slave_transaction)
  `svt_data_member_end(svt_axi_slave_transaction)


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) Tests the validity of the configuration
   */
  extern function void pre_randomize ();

  //----------------------------------------------------------------------------
  /**
   * post_randomize. 
   * Calls super.
   */
  extern function void post_randomize ();

  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode (bit on_off);

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();

`ifdef SVT_UVM_TECHNOLOGY
  extern function bit do_compare(uvm_object rhs, uvm_comparer comparer);
`elsif SVT_OVM_TECHNOLOGY
  extern function bit do_compare(ovm_object rhs, ovm_comparer comparer);
`else

  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_axi_slave_transaction.
   */
  extern virtual function vmm_data do_allocate ();

  // ---------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare (vmm_data to, output string diff, input int kind = -1);

  //----------------------------------------------------------------------------
  /**                         
   * Returns the size (in bytes) required by the byte_pack operation.
   *
   * @param kind This int indicates the type of byte_size being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in a size calculation based on the
   * non-static fields. All other kind values result in a return value of 0.
   */
  extern virtual function int unsigned byte_size (int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset, based on the
   * requested byte_pack kind.
   *
   * @param bytes Buffer that will contain the packed bytes at the end of the operation.
   * @param offset Offset into bytes where the packing is to begin.
   * @param kind This int indicates the type of byte_pack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being packed and the return of an integer indicating the number of
   * packed bytes. All other kind values result in no change to the buffer contents, and a
   * return value of 0.
   */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset, based on
   * the requested byte_unpack kind.
   *
   * @param bytes Buffer containing the bytes to be unpacked.
   * @param offset Offset into bytes where the unpacking is to begin.
   * @param len Number of bytes to be unpacked.
   * @param kind This int indicates the type of byte_unpack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being unpacked and the return of an integer indicating the number of
   * unpacked bytes. All other kind values result in no change to the exception contents,
   * and a return value of 0.
   */
  extern virtual function int unsigned do_byte_unpack (const ref logic [7:0]
  bytes[], input int unsigned offset = 0, input int len = -1, input int kind = -1);

`endif // SVT_UVM_TECHNOLOGY

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>read</i> access to public data members of this class.
   */
  extern virtual function bit get_prop_val (string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val (string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
   * Does basic validation of the object contents.
   */
  extern virtual function bit do_is_valid (bit silent = 1, int kind = RELEVANT);
 
// ---------------------------------------------------------------------------
  /**
   * This method returns PA object which contains the PA header information for XML or FSDB.
   *
   * @param uid Optional string indicating the unique identification value for object. If not 
   * provided uses the 'get_uid()' method  to retrieve the value. 
   * @param typ Optional string indicating the 'type' of the object. If not provided
   * uses the type name for the class.
   * @param parent_uid Optional string indicating the UID of the object's parent. If not provided
   * the method assumes there is no parent.
   * @param channel Optional string indicating an object channel. If not provided
   * the method assumes there is no channel.
   *
   * @return The requested object block description.
   */
 extern virtual function svt_pa_object_data get_pa_obj_data(string uid = "", string typ = "", string parent_uid = "", string channel = "" );

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB.  The pattern is customized to contain only the fields necessary for
   * the application and tranaction type.
   * 
   * Note:
   * As a performance enhancement, property values in the pattern are pre-populated when
   * the pattern is created.  This allows the FSDB writer infrastructure to skip the
   * get_prop_val_via_pattern step.
   *
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
  extern virtual function svt_pattern allocate_xml_pattern();

 //---------------------------------------------------------------------------------
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
e3MpcpVsHiYlJ0Xw6IUjDolzreckis63pd9Zx0jYQ+O5cJfdDd3ManzSP9Nfe5RS
Jn1B9UzbDq0ZS9DKFEitfKqKmwubrLjj58PjdPIxeLUsjRMG9B+TkS8LkOqRVocg
HDdJVWbfvNJhotFXDePhRCAybfdnMvNKTSVkzUICHE8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 29335     )
YybehXSA56rnFejabKKd3K4a3RyyjqYB8gnUURkphxHssr8+HOx7mgKHaBym9MhO
DQrDuW53tvuS+NAmf1Xgez6CLfptESq7bGAJULoHI0BU6tNTwMCV3xOPAvaDZ0dt
zvdvAR201TwuApN0nmlRUs4+Ie55sJnza4IWoUQV86A=
`pragma protect end_protected
  `ifdef SVT_VMM_TECHNOLOGY
    `vmm_class_factory(svt_axi_slave_transaction)      
  `endif  

endclass

`ifdef SVT_UVM_TECHNOLOGY
// Declare a sequence library for this transaction
// -----------------------------------------------------------------------------
`SVT_SEQUENCE_LIBRARY_DECL(svt_axi_slave_transaction)
`elsif SVT_OVM_TECHNOLOGY
// Declare a sequence library for this transaction
// -----------------------------------------------------------------------------
`SVT_SEQUENCE_LIBRARY_DECL(svt_axi_slave_transaction)
`endif

// =============================================================================
/**

Unitlity Methods for the svt_axi_slave_transaction class
*/

//vcs_vip_protect

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
m1eEJEAdn6NVdlQQDLknqcaIJjN/F1I0r+BlkeVCqnEQ2L6NEydtQfIrRj0LTOZZ
LWMCGMUfn3GCooV3PDeDFJHsm8NvxN3nhShCwhJsTRZBvToTSjInJtVK7mQs9TUP
RNuZ16KrUUqlmE04XuP+fYE1zj4EmtEHq2UkO/ZJ1Wk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 29868     )
HEvYE+23txDkej6AtL2dgHl7EgKDxGNYcLEDXyu1NEqHwjO8obMfWhK5NYIVCaN3
8u84AMTgvNoKirSyFi9I5GZZxcGc6uFoZnGz1qVu34d0yC7FXm0zGWhCGBlPXch0
ZVZnBeMAF6qAkgquzphdxKzsaZLtakkoqsh7s/PA75f75XY+o4qSDQRCGS0ahRq8
ocKJk+Blw3nU1vRI75tXa19x/kAYL3jcguDMuhrzXN35EpGQA7EDJmgfOIRQU1LV
70zHvgXDLUWwAnZUbjXSRgDzmnOy/7APhboEmSD2Rq+ALEAh8vfG1cWve0rStlT6
p0BB8t36kzDdcYapt0zj8TGofCE8Ny3qZrd5Hc1vd3PgN/0XY5TK4uINmTeuthfQ
bnrHXAYDqhiFcgHXBSd75u1ytK9TGw9VQ3uitioY0lUeG52S9L2Ovxd53+75891S
a/x8lLTc5fP5aja0OzAazy68prvsCXwDCRemjTDDu3WtzRuoILRBdvgVf+e7vW9i
sQxcp8d/o1slGHcxT/PHvHlE/yN6YNgFd/FnyVbKDOP6AvE2bJza9iYEV1esig0I
1hQqnlKMP9rG0QBGq4pFlCjXi5cXbHxWXhUyPIUjwsJ2Tq3qTEdwWCq10cP6lmGO
0ZDDGXMPcfhg/A0HzmhOu8ValsdixfFa4zffnx1kggQlE0/WA1XHzkjIVpa/qssJ
p/+t0P83YuemSbRdfxJoUQ==
`pragma protect end_protected

// -----------------------------------------------------------------------------
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
AmevlKD9Im+QkVnVpucQExTN58XxF+ZcGl3/eOEFfQQnNi/6E1iT47zppXxF0jZ4
s33g5gMw4QcegYu2PC1jpyWtJgVpYgSujnVqUXgZciZLVNIWKGdJ49+yuiEU+JOj
FQvafhd0eWNVjnjotp9GGfDE9f1isUFaNk7mG2+u6Fo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 32419     )
peGtK2jK5BcrG3Zg2DrMR5AjbUzXly/BY+PJiyc3WczO9t0HUqbbsATuiq5tREfl
1/YNR2oPWVLvCHZG+ANxWPHt1EMpwXfyLLaMnu4rtsRapDlQ3UIiFFUGdO0dMg9M
ONfhzHBitVwBYhx+iirlZR58YSZ3YufWobQXaIa3ZrxvbRIXJ0zgS0r9J9OYbbvL
8HjsPlZWy1XQbWyp5s7wW61n0gFtwev6J1LZd+5588TGHeUz6RdGPAt10n1qTLl6
DValb1toS4BRRrwWcQ0yFmnOA507wn1Q5Xvac6FTLBKx+6MqgmMZa6oWVNZIGzq7
JQj6pyu4oqBR0P9L1sRhDW/hLPN1WBUQW1HtX6rAdvqa/io2ejIkh+EQabpc3cVc
siMXu/0/9vhvPgumu82a2kgqm49+BCISsFCaH4Nupg308TxGac0IHGxyuz08aMMa
zDKB17E0RlBZVXGsaIvaSVTf7iftsTfiUXxEm8x3jY1LDkkLron7qhEQo+FNHlca
v4qrvNtXdpcsyDQgH5mXc6MD8WA99dEmArF3Bm4v4r685azxeMHyaLexMWLGYzG6
LBajOrdUn7D2cyZ9pry+wr1Ht85VU5dVsNy5P6QIYQC5EwA+7fpTYYALC3F2Kn04
1b862/y8eOf3qSmYdTLcz27ae39NpYyxnGaEz0jo3XyRGQc4IAzuU+wC3akR8ple
PLKsgztQjxWVKoYbrKUa9a92495TJGwtFGawwshDyDZwvfcbe7qEMCr0bOGPU5QE
oGebi6mtZYXYiOEbYacQY075o17JBqWGRqYJsHydnXJrGyerLnfjj4Q+m2G5Xrxr
2uig28TP+vvISySCv9qOBYFVt+/hQDvAnxNCnIhPjud7RxPVns3SF53OPtyFHO8B
TR6nft/B+4iJZWAUe8WSk1Jo6z7icbGzqT6Eq0n5tFnyan7a/Q2jNvWvC+xcKdOg
3PTw0mbaxLMoZCgh70n9utsjX2jbhhiGZFZxynieYQOT5QtfBogjOm6/1V04U9w5
DZLTu4VkYvWmnvFSY4WJ1m8jyyDyoc6J3eIMyY4ermXjfAUy6Cc6Ap5nFuMzM49a
wbhNM7PgHOAFP9pxHicUG1P1C/9IZxAjGWVDl/yRQIl3tyH81sBxw+mUhg6ik97V
M4nh9psNWgSTwCL/hR5wJ0AHMGczAn+4rFlI9MAPEL1iGEUkm5v9LJIhRUI2iJ1o
ZqcwzqqpTueA7RGZR+AytHW1g4Vjda5adtF8L3yhbiqDrVux4eduE+qxTlzzfw6u
AzhD6oAeuyRnY3IY43DR4UcYkaniiqchgn/jRgD63KqrEHWo3++7U9jCULEjI84c
Vdp3vqXf7ZIiQCFNnpjB7ChW0jvVJFYPEEYO7FBacIOxKs8IZ7Fe4IQ1FJLydOxb
3MEosF+pDjv4HCKhSVUh2y/bTQJwc7euV6l68ceme1Yft07gutp77fEDtyomAuKc
PlUD0YzIfxwi/JkGIvkQUIRxv9wEVD9FYRKJgdD1S6WkYx7RKd8MOHFzYS+BBT/d
lHNF66TtWP+KhqmZdKNOcecf+t5ugo+oEmyQYCd0kAq0x9Hzuaa3u3v5bk3t2Lip
q5CUzKgdTIWFacdLLAsSEJXrs39g5prBhM9PjKTOd0xxT+wm9BLmRjXPchF6eS8g
opox/Wii21sSSRerLGubz9ar1jxrfyiPG/FXrQbSnRkh84lTFHyZ0+P6LXfEWN5G
5p2zmC2Hd1RRGUEjwjlb95jRiz++Vww/E4lMAqOzN4g0JfDFaJCaFWblHpqhNa8d
UsFIDliPaJ8kza7mkridASiB98JIIYa+5s9snyHjHh98lYD4Ystzr1bQAkerstw1
mYwy/Z32bwW3A216tvV4YZYhcBQog/Q2y6Vjx/FLn9+GB5B24dC5urWRQXdqUR7l
IAoZMmWywNRp/yqwdmuujO932CgcsLioUxVF20YEbYF+Kaabd+9WilavB4lgv0MU
Hnl/1eR+ZtOo2z7rfNUa3pRKlIBkYXNu39QEZ6t6CmgGU12Fi/gHDWH8Up0/sWnt
wff9vV1ZoNnYCJZThDqcRY+k9UI8RGBig4pulS86wNS2EkSVy9IyD4dWIWNOJtAI
+Zdb+TtMDf+p+OZWxiwTvwq7oM3oyHizGV0PEOFSVNdkC1/gwyOR4ZLpOhb9OMQ2
KuLWFlan7mGmKQJh4TnevhT3hQvjnQ3j5PrVpt9lh+A6kdsdhsc0qqPmyVX5U9uL
JKhjVRzbvTZ22GLlsbeRdSv6aaTP/VhbXLQ0vbnCYJJ61wwTUQC19VFZMGwwd6VN
Fbx+c8KMecQ8KP9X5G7x8zxfrxd7kNcPCcYYcpUT1ngS4ZZOoSPXE12i9NMu71vg
MTeZ8uzeE6ZAiH6+kC171CVO40QsZsxZ/eLlh7uE0jmNTVmj535JaVpJP//ckLeD
dhRvikm0w+mhTAYt2vMjA+xO0KX20aRdZHxG022JwVQvrZdhymbtf9UfOO3KfASP
1VD06ru3pTr0bMtKK/1BCnlYqpK8fvecejLx+kKThR4d1SnavbJ3Sju1J1ZSKp4+
uyQmlT4TkoRmjtoEfRokY/mk4QXM6CerQCK3WW5QeiF/xZAYoGvybLchMtbeFC5Y
b92uG9FCHgzCRBbo1VL4sA7PezeI8x864Jt8mRwp0xK9+Kx2IdFR1SqM2CjjXbC2
mcWaBAhWdNBmsW6RApR7AZUT4iLwKGqsDbaVNAKIr/1ZqlL9FL96s8+DAW8E4jE9
EJcXPLJv+V44bu6nwTPvirlEsQZItMnyn/Sez4xc/+OqvBwU50SJ50/TWp2b84/P
NCty3xOULqtSFrwoEGBxSxgheAe3b1yX6clp43BY/871CJ/xGrhbQ3a/M4yBlN+O
x+vIffBRjVXKSd2X/J4mawINfs1A5ZKN1BIhv27kveEakFjlr7yURxpZASf7zsZ1
uKrxqijaZs7BMMj3sNqMHO6oOeMbdZGwAC5nVP8AoV+XQA6ivJ3VQ+Trb6UPWVK8
SUw6/hUMP0uKDWDMjDTYIjIodzgthzm3LCsGC7Hluc4M4ZpRX2YVYwSXj+lG8ABo
oBEAJ+CSElKSoJ1Q+NuELB0URD4q2OyVsT9Y0CIVdH9QmoZG2bYvEY/4SPq9eHYs
7l4WSbQtV+YjnuXLka86WfPIS76gL5+5mlJa8iM3C6tAMTx69dgbBF05JVR92U7K
6ETmI/9Xc+o325rkjBkPNLlhM+ov4Fn1UGN/4DZYJo1liVUcB8zzYKbUU1koneXE
wBN9OwOZP4vxi0AcNGcQrwzil6wjG+2CEKW4N1gu8r36izwV4TYyN7ONLtj4jMCe
jH2yM7XJethcDLskISakm41WX/NB6Ghf0mkLoQKEoGC5WYOJVD1lXx1YMyBU0IUR
E3Wkim3CXpwpe5AyFG9m8A==
`pragma protect end_protected  
// -----------------------------------------------------------------------------
function void svt_axi_slave_transaction::pre_randomize ();
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ZVB+Pgp3T9nFUTZmBlIJPSSr71an/LsUA0QldHI2KDdkS7fjr8qYTABZhrYY1E8l
UTvTNKnLLuusN553mHNwnS/8AoMKqqb+Bj1w3mN4Wvk9mo0xYS+lExvSfJI/fqgM
XOY2Y6iKfJcye9DLTUmqd/6Q0eG5rJpFrI4ap9n5+nY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 33584     )
I6Iu9COFgwiaIvZMBf5uOXLFDOwrMU5WQEpuHO9lRFZMnQEnJkSIBfp/5EVjfp9q
A+zAZTvKKP8895ItWUJ0Y9dkXbvJUYKxEgecrZ8hW9/RtypCTJIOcpoSp1ODriyw
GV5kL6wPMRBHQTF5vlub8gFUFti5YiJ/c3aTjyB9s3t9MGgwEkWxzzPNOHvCOwcx
AgWGWUlMNHxl+J8BjMRNR+TtwV5UGq+8DeyHsvJKTEauicgWTWckOCmEuovfZGpT
wD/mpSg9rJWtGy6D+FBzu+aU3LlVOmMsIwNoKZNS1e7WEZQPR28c1ayBgEj6ebSX
Emh5IU9nAjPPfD20VUkGEDwlrlI9l6uBpKfzl5gr/Id4BvSk2VsjRLL5AhjwQOHb
Nw7+c6cNx/phAWMd3TVvh3ttSNbuCY6sQvr6Dszh+cpFq7NJZR0NFgyF1kuBaKGQ
1da1GvZIsCp7EbCyA6GkGPSjcKOxF1SkxeAclZ0wfNNma6ZiTUMJbwvvFBr9PmWz
w19Z/13oer1UIOaUlRBPtwhE060vc8MpmyLUf4a2/QgjSMrdPiwJRgeV74UyLPRp
WrKHAID9njfb5E+zM29xzTzxbI+/2sHyfjxCTFqBo/7PvMBqDglvNmi0xWO05erD
XOVBzUbok11WXnwYHOrPtFxn24rQG3t5mHJ0HlRdGVZ19/ZXhgpumQg68Hx2A4mK
7REErmaxCOyTRu8xMEgtHAM5y5sQ/zoD1X8szL233UUkwhAQXmYxx7CYLfI0KHCZ
0uTNLkJ2ULhgBS+bxThgcEfAkb/jZDnbGKtME11XpxtKgmJ8lQlZeGfrQDByS2jf
HxWrAPh1HFkoZ1YAzHq4rUupuJMOMg0h78HsU3ChkKV4fpMhM6pYARjWqiTSkvd8
sytwx0C6Th75KLRT5kWaM/uytzCDAYwWXN/fjPxlR8VWDPotlIriRD/ObumfM4Jh
k1tTdpds+9Ve8y+pQakSRN3arG327KNHbRnxmipAH+PWXJeSPlW9l9SRba41ZON7
Na9g6zDpTwN0QV8gr04G4HXdBWK+pM92sgasq4kQ0SJ6bx09yaGq6eakCSwsV62+
G6TTC71Xkzyd7u0qkJMl2jU4Cgn3jxRoCul2Ap2Uyug30EV5VHq8QFcXyyNHN70n
DScJzPbNDhK4xjGBBUm17TGfRdsw+6Q5fnijYBjgRKxYIcM+WfTUIt57PbLd2ETu
RIc59FhRezIVgO+8u1sDkuiDY7x3r4+mIWSkYWdfzq7blx9H/ToAHi+AOJ0AGVQo
WvUXKsMVB3AasdgbHwR+h+VJibBxGp2zJBnABDSPkH6g0hDqNLZ2GrQGVQ2SCZ4/
Tof0+LqVXeLQDYLoCODPsX2gmgUSAcKjvXwrm5k3mabep1ovBJhgwgc7JvTI6WMp
ZDZhbiKTZZX+1tfkLdeCIrXEk8oKS0flnKI8JJ95mxNAtqojvJCqFt9aJDdsOFl2
F7i5QmU61lkE64qB6xC1HcmClr+yFxIMYRLTiOKn3Re0scA9V7UXZA4OLVbVv4Fb
VOPsxw/OlSUclNYsE7LWpw==
`pragma protect end_protected
endfunction: pre_randomize


  // -----------------------------------------------------------------------------
function void svt_axi_slave_transaction :: post_randomize();
  bit data_only = 1;
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
SW+2ywANWzHlvxjgnA+gx2ExKOLbGhOg1PzmOH/Csebb9flWvAYnFhxfFbRRuANl
A8/GUyc2KhBx7pUuJEOcVq2EH7k6zrx1AIknWs4UX669Gt125VNsGQl2A9U6oinL
ajjfPQeusxKZwV3LJq0v1+knqM+zcylpbFD5086Tm3U=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 33693     )
ALg19XXQx3uzUaYNz1h7GQsA+rdH22EY+fDFeBVj+9T62226uI4JlAmTrYMQC6dA
glMHo3PjmibhC/R0OK9sbglnyGH0gjmLuD01gyztAkNZXs6UpWDO8tmsDD9hIbHJ
YOvStVbVIF73lnAoZxbN9A==
`pragma protect end_protected
endfunction

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ekEdZ7yM+EzXBRT1oCeBq9gdhG7luzCrZLPHdFSUTcweDXfnMCKrHCW8SrpfHFfh
vSKKzdMlFEEPW6o+CLkIHoHFGpoTE4C3jLE9dyEPxxUmMxYYiySfv25t3twW7Xi1
AvNRg9fXutTx2EwtGqreWZ+acion9ZPmgwc5lmhtN1U=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 64299     )
1DdvoFAgxdos7iEaOp96tNtbiHJl6pqusbJ2vS+tNSaQ9TGG8xj5dg6xUEUPUXzp
XWuoIDJUByDwmWRyUPq88aaCYF7hO1cVFyvJtgsXwZGzsBMECWSM70JpMhC2Rtpf
60BitCg6TQlJuFvu4PuayaKX4IRsWUkn1Twlirg9fIwWIL/dWcwiOtQlYlY3qWYX
KNbjwcRcF+6o8V2OmSIA6jhxrL/Fw+BnibOAXo2kMLYKhf2vB3KVdSL9MMoPOK8e
hWLP16VvBL4X5j6AljUQjKSqiXx8EIrg0zIjp1Ww+w6ZOWo2LeK1pk0V54oHAbBY
j+pxJQ6lxAPxwn2a7fAJoxCTIB/9xOq8tNsNdi4dWh/hSmbvAlkRKdovpBFFHP/K
rRZcPwVCFRZvfNNbmlCKjagHYsOQzRVTlCpOu1tlDZ09pFP70B9rFnOl0KdRxTep
G1ySVp4F1cQg4uywmOM+5ZFdNAUMv6cx++6d/gzVLzCtphtD1O4DlaKSD+gPkDnJ
o9SLqdIP2QvkKSkGJyZ5XS1R0dj+LpvI49Q0zTdI6wjYLsAbkWtcinlrL8sDx8xR
qOrhxRrQICPzvJ6bGWL+6X8grroWITBe//PZmQBZRfFFcwZ0n5Qk+zTCbdVE9zzp
g6xaNyXg04N1RAIPDt/jbj5rVTj9uy3aufFdro/LH6rvq2lGxHoYiSQIEOSvrbdo
c2vymf3brZAr3bvbhr/rnIU+H7mp/umfhV6iQIEiXCyIA9iPg99eyaQOQh2Dyt4H
VI2xxIa+9Ex8hBZFmdtcF1jkMS+dgkeIbLRK8gC25IPVEqZltRksNvxvCNbGVc7F
SKAU+h7i0OAkdiVDAbdoG4qj770m0O7lJAbsr26vyn5RsP4knCUoaGNAl5Kv+GJp
wd6BwLzw9s2VtsgoYmxta+ZqLav21UY4+TijzHRWwVwRclI0DU5frg9D45Ls3KGP
Xz3+lA6thcRNU5QM2R/sFpnmanNPY+Dc3Ff0rzfdHkBV+dlN/Q3frlaklCQHwEAB
20AU4uINZKXLKOheqjSYrKjKiDWxEWyXTiNdM0vxRy+gVw/T0hOjlHwozEyrZcbb
O2sIxWj9jCFJusb9zEX+CCpkLtntZw0n2vGv8bolIiVtEIZDX+5GhP87F0PWR1ou
es5x98XxTZ6yRf+TPyZhnLacwN7NcJajHNB6DW7O4hb/4sOse9ziO6AJDivx9B2j
PD91G1hJMGE10tKRKt0ymAPwyWrqxpHNYZZ+gI9WScrETBmIeXqT3b9KoH0EzwTK
0VY1/X1RRJ0R795E+OAUQ05S6qQtfmR97hQW+ArYoxxAbyDzl5+ngxudS/mdOh67
8fsuXTKHIC6CfuRJvqKDKQ5+5RziGQ80kJUUv6KzBI77EKqXUsbFuylo7a0MbUTg
jHh/wrWadCR0BYlbS/q4vRkghS6yO3VAw9FMumrWl7hFhiGp2JoemOCur019etoI
aRW4pGX8fmrpJPZprGumRLFa5BZjY4zrlFHbJ8CiI93YwSk/xxoNyYnWjVfqYrrN
RDOg8xKYrxB5wSxiLs0NI7/VRgJicFDn4/jpg6r9TT3wTVot1bB/Jpid+qyC1gfe
zticlX6wnx88PhAWEJeUdT52L7vosApJGYPuZ42DKcFg2JKVc2fXCN8cWHHYdkYB
Icxes1gh4HBkMtJNvkcybh21DkZSM5v2nWFKQogURcIa02XZWyGGOfE/ytPu37PT
dyukhd8iwKvRUi2wAAIoMXj2n73w6MEic1G/2XRi5s2n/RVFV3/KtDNcopiAVSuR
5kE2mz7uhxRAcrYZPtGAdnBf85B/nuulZlW50DadQmi/XXSTT5ZeDhmUKu1p4FRY
HV45jlUQ84I1kaK5kki1upZL0ooNXUdSjuKBg4Tcfq3W4wRgcqz0YahLoszA+zE4
0uGMoLkS+/6EngSJPqzeWvZwJNxrNoyhDSxWZk9Khz0+rpXwokiTPJVQOqQ6kmpI
cJO7s1giGNUdcb0UAKQOMTWAaDUN+NW8nnJ042b1zS1sTf8FOHE50GaIVWNtA2yU
xeZNswrhpCKrS+FB6KIEWDTEGoZnP438m4A1kU4sqNZgEyYhhlvbCr4EWJoHERZ5
DtxMczzXNEfN9wZiIvkH6X0GoTJ4bRDuc3XUhitgqwydu6PwEX9iTOjeButZgN6e
wGl4oPmJZytJK9KvRsAYWz79B1l+xys2yhgg5vGmNB9wPBjUGnVqHrSRk9ecDCFu
OtzrfdoZrsfi9DJfsCmF/yQ91GBlWzpBFh3uYLQ+1vipLtDQguFHD/HriGwvS9O7
RrjsH+zQlYwJntJ3uNciqasG7sh3KIsXhgJJFvS7AVqL3qXZIlQzPtzYuhzy+DVu
ke2jiBiQ5pthrJ/FO/LFWS+YybZeHBw690dnIJ87q0BPxBM1THRWcP42S8BJO2vl
r0izs2KkA7/FXoduWV2AP3oRFIdkr/yk+O8gXXAeZLCi2acz+kn8r+SQ+EU0Pf4s
YtlMFprrI0wlu7vcqyDXU8A3KmezOs0YpvPvSw5ZEAZ2Z40k92jXT02puj0oTTmr
aegb0Q8lMjFhSHHOCFrRM6+zyGON+4ODUXaZuE/bqLp41kMN+HjEi23Z78nMRiwH
WC7q+JMDoyyeDhmx7HMmFqbWfUT4Obopu2qKv3cyIKgBFNdfBrfU0gWdlQHB5iPV
AghckVVOHv63MHtx81BFUgHeo95l7mnjGXexssEnkmKG+yVF3PH4XjuPMswB2dlg
3DzJh9SCtkVeHbGjHM6TJ1DQ9jB1CyConMyIxw0OMwwJcN7twD80JMhmggWeweKq
AyOzmANYL2wN0LlIH5ZZ/OsJhpnd6HWo42eoEMXaaln/c1f3JzDeKffG2jenNv78
LfuRYeV7zhmX8pmz9XaPt9IBh9BVyrXuRW+3GkvsQY226lMkbN1ENAKumFjQk9Xm
1A7Zw+sYirQM2PiIopD/axcLIp09Zd3iN7B1y4GW2wUxwR6kaaLvbIyiFYqy/I9f
K4J3UTBYRf1uCGLn3XYy+B4OpLR/6mGG+rwP2gmCzOzHdvtizSLlbYkGfOYOFwuV
X4XmDcfMVfghauE0P+iLnb3hO1+RMFHgCZcQ2RNFt+VWrA0x+y2p3Ix+0oYKJIS6
8Iz1vmyKYsuC/0brmToaCvjucgQA0u3Nf9Ye2sgrphpU6x3pXzEYawNjznRxA2NV
mhsohH/NbZODBjosj5BmTXJiw3enpC9CBhWSgtrSpDJ0yOQM6aVh2t1JSu9JQNSs
+ocI+JEwGc9OGPTUzlNSjrcgGO02WeR6UTZdrVm4Fz1LWy2koqbw7DxnufgLPqO1
BRw6RCYe/SrRz+p/hwOCuLOm/S4Q7RefihL0wAYK+cJNlhq8ki1JNGLVsgjXHdIn
8dhFqMwKBa0B59fWO5HmcpKtCJKJ+OTUXy9gtKSvSFy2/hXaDPoh0lii7jeCqtX6
0SxzVr7dsLjOY/cXEBCmMIRncW80wRQA/rW0JvgZW3sRW/Wf7RZ0SX5eGiEbU6ZF
FEGmo4LUNhEebCf2S6t3Wp7+6RXxQpYwjN30AGG9bKL5ClUGojrIvdNUBFylui/O
ePgJAcoAQX3Kqg/6k3uf5DTytyBEbbMS0+l0XloeyfOaIb72JB77QYR1nOvN5SvF
mTS50qH8IbB+8niLR/SpjUpta0vXYTte6f7WcuqfFqRMljE+Rww2RTa2YKoiDVFU
jrVfHSABHCOY74CLYfzYTflmV6llshSQMJnazf02AbLN6JeoeSjLxeoZeCg05t9b
y7b8IpQFtrPPsvrGSujLUcbeMdC1TQPfW4TQhIvoXVafowr5/8y+OFIvMQ9owmjK
DnoXzqc0CB3gbAL+BYVvDEMqxzhSEkkITXOlrUD3AcVnXST/tmRjzPnTx0Bwn50u
whmxrYdHvJDezWytMwZ0ChC/f/vuxkKx++cxFIxVVz9fgMU8MfSg2KEi2X5VOIff
ezuUNCyPlOAqImZaoEGaMlKWQRhR+XT0hlogJsl4XfYzi1F7NVTWK7b4YNQomawn
wswAowgzSNLq3r6L3onuc9iBOQxX4eUZyi1XQLuZIfrt+XXRRg81J5soMuLd49F/
Da7Dr00eLp8b63SXWmNGWsrGWb28/0e5gwDfgzFwC9bXZ/F8XtI2cVeltOgWSuHf
ctPj2AF/4DjYZ8cL2pwQ6w3cS1qmGUBbqFN23i2oFRFuLao6s7WORKDPrhcT57KI
bo4bc1Ma7WccqDOPhA+Yhb9UxuG6gQcf4S9EUeCjBTRzpGlgYz0WD0s/lcUMXeT6
xKJKoraprDJmgi/FYoa6BiHpD4HzkgDWRSMpV0x3DE3nUpDxAfJgTNgcUo9xSg1p
ZgviHaqRH3ehGBzQO8g9xyIdZrd5+VNVkblYdKq/4V+W9aVMa7vMDP+b1AwCO9HG
1ShZSnrtd0Ds7pM0XsfIabbCxdUtCALWGnyE5d1LZPIFqwVZswmyNA/+7i5NHzZ5
tzLiu+kWhyBkXJBLwpCSJjw96MDmd66bSYKGBM043Xu0uNcPSL4OkIVkJ2xuVRZE
DnesFGrSq9CtzKS9srCYed4ptg1xLRNpYnhxQecKAnIjEdV7zsEdpqloHO57EBV3
ab6JTH2lfmeRJ+5PiOgGx5KuR9AIOtkT3wgFJnydD2AoyX2UleoumQJIpdj2HBFr
vM486FXMD8ykJpjzEssv+tHy4dGkPotVnNCAg4riGxV4I58mT12JMlMPuLNMxcES
nxGa5+pnXCzRHe/kdzaWXIrrYFnDKC9AY9rS+CSJciN4QQPhBcLi00DkTUIb8KiM
QnKAu1F5Vrnqs6I3b7wkULNXF3ZLXdU6eZ9qRoMDvLaJLp5lBKFDzTqtaIkyK5Ic
nVFnMI+nKHr6WMsIImi/5gyRRBytBZpRxh2ZPkOgOrm4kA/JGRDwWSmCLneWM0G8
ztDDjGLEFiwbHpnn/wWDE3MdVHxrRFYunSCpFVoEcH/nWSR18vf3eLYnbXmFnIkA
0TTbmKECnQo9fdtff3kC2floW/ErMcRTKevgwXyrTB/aFMZw8jGTayQ9AmRgG+cC
x7N2KzYpwICPtkp1djNaSylwWgmDOskBu7DNNtrlmL2vaVxEXOiY1nMb3jqeyqeI
OzzOsdMvtui1jA1HL5YUnCDCGW8/oXg2X0bQTVZ/1JpdzJWXrnNElvHQfGa3DvfK
j7ldTm+CDjpVmkCSIl9+u0ronWtEWc+EqDi7nIR/Kinl/nRss/epvWiqxRHc+3e1
IRZJYuivWo9gKCW7ufRNXsYrUuqsO/7Noj3j+bCd6kKkDC0aQomJAQOTDsqdxhNN
OIaAfQM1DqzgpqDysfH9JbjphupQOEStivUygEqzzKX5P7tjg1gddB73acupXOnJ
IL43XSJAwgU3LJANd5iKl8X3Htp9Vd8VcRLyF0LONg3X/atUMerm9jiyryZR8iHc
5vl94Df1Mj/MM3PxWs6ZCXkkpcCwi9Jj2m7KqCuLsHPZR1HOLNobFQZjXVfz+w0D
e+VL/q35XGuT3swxf9ur1PsfS6iq66OKOQ0ka4xpHJjOn/BnwBlESP5QCV/GlO5G
TupgIFHvIG5IK/YAKgDVxixTp79ZhF6zSvWxxsMiR6A54AwhjrklFl7a7IBzLVx6
w7baVSUwgf7hao1GTRKYIIN+dJLC9cnManRLz0ejUrAKiKnETgefPRwbIQwCttPu
FqKuBffcYQbc9Fn3p27sNoQMatjhUZZRXWd8z8qYcmO4ctUsQ1xVrXYRCKVYG1GR
gLE/l9WuXEZzFwgsiK8YwCHOiQe2viv/FdsFH9JMHABjV4lsWxmq5iXKp2tkPUwu
2zf4YsOGIQOChz4lJ6FSnJrZnpLD+eG4FT1oADHfml6XXbIR2w/56iykUD0H91dm
PJA3mdZ0DEUov/OpTmdhf6L9FltiY0KfPL33ktlNacRg9Mf2LJPXdwWjhCLApLwc
YRWhB//vmdl50jiFdAOMlrEnv+CIrj15Pm6l5LIXALT9ZtWr4DP5HKBnaOCJHkMs
z5pnPXqNxTdcMdetf9xrzDd2wzUfA3N6M3uJQQT/NTOXCSky7ecINDjHUiua2ppw
hPkrn85jbLxM2SPYcjb8sd5YIqRi4i13U+gLRmBMuXV2Dw35cN0lGJTmMttCe898
gxv6yKm7GfGkt4B0Ii0LC2KvQf4czCu1Tm7ygjkbsVYfhaJH1VDvvM2b6oMOMCIJ
ALMbLC/OMSX9jXzVIRo1s632libfS2nfgWn7009k3/NTJ13AUv8cQ6+gl1AoIJw6
R/T02JnSyRDJ1c7MhKklxlKbh/GvQrVfokDOfwX95vFfhQ1bPlxvvgUrK6ef0vv6
j1Xexa6hIESfi1YhDntCCpIHqObC9F0akbJtHCqsHiOFOIgQDTJ7j9ZxWUDd+L11
x8Lu2cDvT2ycfwYnlwlTc2fnHnW7b+9+wjViYYh+oLcKkmhhXDKkaBhunvdLR+qY
oAKjxfl0SnTO+FzanbI7baZyABDe0iX80CZmUDZDHPZR/palk7Vx43KZoomQxWPT
DmISrW2UBS9GM7ozeRra//f+IiD6DIKuvUUPLO22cxRtK24MFkkxYwLpBicERKy9
kXEkO7aEeneyeUWnjAfX5uE3Egd1blKO9mvx2R16jKUct+e+dUSQ722u8Fv3jkUF
6tSVkJfq0NcrEDXNxerKrZVgCar+2yGc5ftSi8SaDV+O9DyXfzxVmn3RgAI2k7pQ
NMMZ1owK2B/siI0JjJ2Q730V0zP+lyHzpniGizrioTqPWi80XOXCR0kvbFhIztOY
j5JJ+1silS30gx15Z/qTNUC4aKu17HL7Zkh9q/mIuvnJmuyjjEqsB2wzEINh1hGW
TyLG/DeljU+zMCzwJ2VnHKchxAjKhgbCDNhN7nXLjl7b/DlvTa0WiTO6x2SoLNk7
Gm4oynkoxTjfAhJUDt9ExxJDdmT3skgQ3/N9YowjC3Ygb6Kr/T6vv0W34qSQ9Zhp
yiQjCRuAjOLKHFzVNsXP9+qZqo52J+VCa2eraRxiCcbD3TWnfzby1Qh7cEyWW0kG
w/HKpuRpMQGtIhHoYY4O7kpTDswKpGtluchC94bdTev8+YuPWx0mvQ526UAA9h0v
qMHmafyLVpolE9KTEnSFajsCydretgYn+8vwfFowcpEi0ACNpDnru06h/6Qx3QhV
dyU/LO2IxjWzOIQZBkZTHc3W4OP9PDTdzldVql/lGzQ8M1VEP0bfcAvSLfTNgt+2
mmteTN8G/qBvvhix2qX7HziYsr7JacY0nNrRKQdG3IydzjLfRhfJ+pPDHlH8vw/M
seAyAHaqVdcTbtkuNN/Ht7uyjqyCZfAJ+uS0bMaqO1g4KFDvgRpqrl8u6sjrZyV6
yGY4x4YDsxRCTagI5B63SK/Y+ICMAO2iGyKjpsPwD+btbTn2oo8Wbj8/83nsFi6K
7QjcCHMiO/P7YZR8KmdX6FFOqPKPtaOTdy5m9ooQ6057vLSqxTuY5cpTBohP4/x9
+2iQkeYABMrVCg74IuFUKlDuUop7MnjaaiSJ63AKFQtB5LG1GhulKvkqttqIOzTl
CX9yDiT+Tru0wGLV5OeEtHU1Btbd14ZsZBvZSABHy7ihbO8WopYXJIte2SQDIv8j
Er1g7oJtQb8OLizM4g+6RqxfSZzoADPyQyjZkGlZR3WgicCtbgPM+Xpx+ySov7UK
Pujy4RUGdBAeA3x5MLJ9crn9gNHFDvez5R7oF3Lxr/E73AHQuW8/ddjz6/8/ccmi
QxAb3g3+89FoAr/wJ5itDlra6p6hAFC9siUalzk5I+yzGWNNNYwNENz0dA5mDMEd
kbhsCeyHH5PaZTxZsW4Q+ObC1ew6qUEXgJi8xdOGltxkU3au2TBY3CPCvWwbBgmW
kATnIpTTEU7wLscF/kcSkxshyaH29TUfeEY43LfY6oa7QjcGsu776P9ReR3MZdmV
eRj2mSp7Ls8MgcZ0tGuu9eIw16+9u+UB5g2k+ZGiTiVUAiBKhzVPDZ7DgL54Q4lQ
BRt4T4c127CxLWCCMxgY8VyvFsWdEsLKIrNtT+yucwUojHs0czVyR8+l5Gwrz7KO
0OxBNiAREBXdQ7Feb7sFF6SRkWbZt1ixPrhCF7fMFpUBM5mGslhWOs11JthMoJ/V
GU3cHS49npTAp81+//BGOeGehiBLxz5ny4hQPQPHyL7y9Zz6p0If8iOSZroz7n59
TdJ3XXa50DkZ/prGHE1+LC/RyFjJ9xkI/iM5kHy9fpyCrmNFAWCBkgeJSZkrMtrZ
RGu7Ui61HNEguZqaDFzUuXz9S0gcGBZrt1S3u4iLCS/MY/6AhFQnU9hX2FW2pJmO
0dDxPX4mjXJcgBZUTSWtll9czV7Ol5Eh7Hk0XcPDq6Aiz4hnA5d64R6vXmh7DNPe
i0b0MG3wYYEpclF/iUESjV1xZy7UyHrRBtAUkrBcTVrplMYa4iQQgX8jCuimu4dv
CK+OjoNbSYPV13iMczXnFQ5wpvnJLeJGZtcjZEkJQQRgwpRnMsvSUdWyqxjJ36Gp
S7CWaMUogpOJ35mmRk3mV+vyP0Lkt4cZRGD96KCsxkC5TfNOF1Duj4DtLT2mXvPF
+qJ2pv9vj+FQTdosXeLUE7Om2e50X5ImJ6UD61ZS5x4kX/5OKoL8ElRCybgHCb6V
EPkdy9gdrC0R7/YKZVKG3KDyrvL5D+zm1gHhQyfauC7d4K5jjPHxx4x8Yo0ahpaP
1zr9BLF9+UE3uQiX56lDw9HzQF9NhUJQqtq6uOo0Qvi5me6YT1baudZTxKPxw+Wq
6p/LueEB55E0N0SrXy0NYq2lhwLAO6iF5HWt6pcNuCBBx1YO+D191bGV5tV/R253
zI+ioLD57A66JX0+3ZrroyHFQ+LsFjh4A3DXCDCNTVMpQRsXAAREU/CtHjn25CvR
lF2DBv8pRWBn+zOqjNl35L9Gv4LPRKfhgsXYDOFEG2v1pxJ58250OzG7YpLaGGkf
uesdd68l29fbjFQXBtTd9bLVFdw14lAO//pN+QqQ+1dazlLo/a6t5ENVnpKRByhe
fbhnCXd0lXv5ndn4YxOT/0nNYNzXDTMiK8Zrmt5OD6UPkH5qA6ejzlrJX5wsRbTu
tFoi2RrX1EQTH0xksHFNVnS0S8QbrXRpVMckUuC0P/r+8MYicssnLUIP+BAJhIyk
rvgZ38uHleJ1fwU008mJtfZx1PhORpXEGqo/UoF33SASi62oHAI/p31sEMfyYbZJ
JMYGvj3nZ/h06FS17qo+8PdnEmW0r9YJ1MBbWKQGBcyee8jiK5LCo09DDkeZzINk
3wRk8B+kVi5dvAbeqT8IdiZab44vzgcxcPIHtOKG9Fe/O0njI1p3HIb+fr/9AtK5
JyiNWJ4J0CpA/Uc75MvDfmJcdzqL8AtMPLfhAFNSFDJe5nTLWS9QXM4+JZ+7qnwf
MvtIDWcEhCDKoYA3CkcNUHYhvB20lBOjw9K9SIpGtf7pucxxw+stHcmfVQaQUJ3T
uBTQs4qZ9KVoLvne/k+bWWqoTFK6P1S5GRd2vSY2/jmS/e2s48+2qECZ7VtxdUbe
6xtCkNvHPin1taNyHAr4XhHuDKmwtEa1mpN4zSRyldn+KXN+ZVyFjb/dcz9DxRkf
V3RyJOF+y/KddRu73Mn5ZB3y05icINDcFUKAqncp9DDFqgLlmEW5tYsh/bL6zc4z
BrTzv1kBpDhtF06yh7d/5pZ1pHYRY92LVLd1ryXSdpcWSOB9XoCOwx4Bszi9r+WM
R4x1YVm+3LLvrMGSS3C9yn3Wu+K8LSuVemWpsV92/AM+G8NGUR/msK07PqM7ioyM
PfmrV0pODaF+BJpZQmQFKkEl8p4Gq0AFnLRNcmkqP1ywawDTS2C6/TCNkcJH59DF
cthimIOKsJDNd4XsjSMoESfDyo1auqAc07bkFEcC4sQ0rT22SzCn6VHwrzmcDApK
AxjtRrIAxPXoQgRz3d3nnVMSk5dlDxv4/DsLzYn+GN1hINkZmGEeOI5RB5rNaOy0
rYzrwXKF5O7A07qVpVxZ4H9i9TdVoyNbBkLzJr48+sIPIbg854R6rN79Aw0dqvL0
Gqw+5A8YQATuZs7Js+z8VdODmBpMm0GC60AFy74PtBTTj8v2EbWbOpVSbsjBJWoe
Juo1OqplXyc8/0A7cKpvNuYMSiwe7pyvP1t2vu0ps4GMgQ1hLCiRBKLSLBYSfeZ8
w7QtoGL5SqWpQPsajkMkDt8YZQNNyr+ax9HCX3glEGxsZe0iJhkQQ2wmBuJU8Fyv
JjlqaiGKVcQGotySlqNtzVyeNkFnIUkt588c5DgSQPo2D2252VjSfIsvQrVSb7zH
anYzIsu+U/qGBxeSHVI5Cnx9gRzcCTJKEebF0TPOth13nGyQZzTTcKtFp7tw3v+R
0nDYTViPWtFoBKW8cd4d/BOg5N7w0T4/k9f7NyOSpLhi+UdiGns8FMY1wDPQIpC5
SBCWG5P+rseirGZlkBX1DxIWn3q3qR6G0E5thpNPsIzz9GECD8+oGs6h2MbL5oCT
bkV3sEh3x9hun61m/ii5D5e5hTP4CbegM57PM4iTqj9yZQs66aMpajAlh3GR/tee
fgA24BKRxT5YzgumRIAYdfyCbzn1EMWEhxSAHD9Ep3UDh81S/mTRKDbX75N8p03n
ILedt1H6TAw3LOg4TpzgRuO0db5oMtCcZpMu4oVMEwITWhu6nbLt20u00IsGUbdp
vap7esQw+eT2wsYWdOzs4DPGSwAOSWH0VdBoTEJnBn9mwp8mwdc6iYOyQEaOTTyK
8XMyBfh1yJa0XkSXyTBsq4yPqRN6T/tIS5drb7rsgXtXhaONOXOxy9lHfCiMiO7a
8Izoukgmnd52/k8Y0ZgFzmgYaA4sF6Ty9fCUkhiKYyXofEe9RDWYmMvdoh+JYRJi
Pvzq/ESHcTOdfiaK9srQ5s3PRdwpmXEGXeuwqaui2s993eBOCilCa/iBsGW0UPdv
kRN9z7/Z4bvUq3lY3wTK+kGZ1ciIB+EG06iV4scwAjqp60/fZU+05nvYZngOwXs6
KDZp+n8x8bN/T7ynFpdX1sHrVkIp3crZ+tS3FfXGkwohAe5Q+PpTfLCAG3bGSuAT
OiLs0tr9X4AgcjXCVQBiV9KDmOGMr865SylzYPynGvjaBWFKk/YqmYVXprEkQtYO
ii0jcUKtlVlrQHO//pTR2yyk924EfV8ccgskrlkyl6KgAILBjBBj9FVeDK6l/WUx
RZa/2PCmFSsAHR2oShxWJWl4liqkerbR+cKI71cevDqwKNUxwGB0kcsu97deUICU
A8m8z9ZW2Z+7Jxa/52OStubFLlVewTE++jveG9ja1+ufZzGHwlPgJgfLfAWmrPxF
HgchURNyl+7e1BnmTszdxqi570aQob0WxdzaJxnf/eN3sxXTUzsE/EcWbM3FBSx4
7XTniQmTljgfFbY5sR69u/3v92EwSCwTrxVK7MSruiTkaOkGGG0RMyeSC8a/iC2y
CrGpT03h0ZZ0kyXs/5s/qVFnUIzUcF0Jm3hs7JPXv6DUEO6JAxvowjAXvDfDQOcr
wrPDyIwGpL7HIRh1/hqd0QGbxq1TRbrhpz72HE+IXnx54+P1t23fp3xApgmbLB+W
kOg95UVhtuW4OJoesnp1ezpENM+bl+2QimYrGa+W9yNUElh9TFCi5hQh9PB+jTRA
NRFJYaHLLcqCfapwecMTKq/P41VnaDCXHxTL9XqcNKz9pCk5jYGSOyEeMCcrLIO4
XhXL3IOIkFt1KtkYC5ZLzrWa5ip4iQzPT6sx7ySaYvCE4A9BOy5Qx775/MTq2KkP
tFjakcAkdbK7T043Rr8/54TMZg2W6PF+TlzLOnluXKV175l4t7kmpu1VtD31Bxt5
Na7JsTmVhDL86xfp6sy0pfSOCRCyvtQDwEyaZ7GqyM38u9YCtVOyYFXQN0vzEH/4
Dbcz+dag9ZSfg5maUNloeyMTGlnl54Hp/tU3NFM6s+ok4TLhwek8mPM0MYWtxrmU
oF5yHyalzNx5drPVWDEKOqxYuXrRPqG981YYlGFS9PiS5CWrg65MRk2OkQPYgqsc
3KWbMEmeBhAzRbe+wlLmYY/ycSYTpENsmYcHe5YlnA7lo4IJ+mWoIjzQHDLCYpWo
bpkJwkBrM8dzUlHNmw3g1ti674+9Sq9lgZB501XA3AtmK8HnErplMDZovB/4LkUl
7xIBKQURKlRrwEbbJO2gJb2jWDiTiZx0sZBbrRKxgJqYTuQpuXG1my7SXZQnnjE9
TEmmwEfHBSEfKEWKoPsVZFbGCOHmqyWk+NRvmqx+VJOtrtlnJr8zXrwCM9rv3T9a
9Lh7ju0s6GzBa1uhd+i/zT5ERvgyopZNGNjLMgVUoUnHcN8gOgILbZ77DdUpChNS
Z9z2TIozaU1hnjPJGCEwY4BsG91Ls5NvOw3fQmjg6JxEMjqX/91xR9HEqNubKEXO
kU7U3QDnj7fT9EaPtUdRShhEqx8VR7TKBKKcGE9nb1GbZiJYW/C+klagxyIR5eYo
myYi/mrF+nucIpKBGrVvMUA67QRr8uv7LFiFfv3XhgSKZAbM/ZAjW689f/Ih7QF/
Ke/i1ODDUopzGe+7JBK+E7+sWGFgjB+9TcfIptcj6rEkt0egdhSAaPwfYnK6P5Cw
AvzNdHinrH0u+zQLTjAFrqrea1ljZEqHlenqYsu+gXCfiFLQR9MEciC9Weyi7G9T
5FuwrDPOgVGxLtpseLcYY99G3yNY7j3PGbAScFzxQMVy9OCrNINktJ2mKfq5N5Hh
m2JnaYqnQU+KLcktDYp1vsuSQHLupePWPUktTP2EZWWktJTRUrTiNuRIcPK3uV3v
DzI71onznnseW1ubV2Nl4wCc/2IMo8Si+IYRnW9S7p+r87tGXYqGv2bdY3qqGUTq
/qTj4mgcjX6Zakn3Pe4aQj2IjqJ1+mW15fGDzP9GGIiIVRS7Afo6S6tzJ95nXiW3
WDyGcX7EeDU5DwSc7hvmqMi3pYjw7sGfV1/cR+iD4Ib1cTTMEGOgtMXwKH6sopd5
oycD2A5LuNZsmLIivr6cVteEpahb1V6CEbTxT8eVLS0GA/o7SoRHcpLMxMPbWrql
IHO/nCrPubrPAKGa5hqMtd4IBGoNXQpYHymrd1JcHJhwIbKSJWju4b/ZfwmoAGPA
7YZWqG4iW0L0ln7tvGRirllrC5V7+9lLSFHl0Hg+NPySTq8wqcu09RB68aMDe9Hh
p5Bg80IFb2kLL2C6iL5hhlO1ybM3ESaZJsiNvK2t5EcpHzElEFDjWL67Hj5mWiVu
lQjXzPIVRZDz2kS9l5NrJLQq+PJ0m7vw6HjWbfUpcpHcZJAdryn9mwY6Yr3ESDEn
TZ7mQsp7tuY8exO7Ym174NwYvQV69Lxz4KKQkmpvS/hiKQREJ3K5Ej3ILHxt2o0h
IygYoBSEzXXQ5g9NS0UvgIL9k2Hx1zz+eV9Y49O1CfGM5ueAyNXjrJ+VElKOpWqI
D2bPKp59sQeM2lKZp9eR2Uf3JzFC/UhfXwW0YaPR2yNUg9NoYsitowvLPb8KZu3/
EC1yat1i8KHYnbcHJjN9JwIspDYNQAN4RtrdFSJ13Kuafv7Nsu9xEXdIGX7BJcKj
gk50fY4qMyOrZHemeZ+k9xggcJ8KOli3dG424iDi0OOoMVSlZvFmH5GPa6dPzj5h
EqwEmQjokDqyVUDf2CiTNkJyJroK2tU7Bn/BhiotjZCCrBfj6gvmetBnWwKmnRve
xkcIrWGKxotG7TnDbGMGcuA4TZMgj2rNoz+0Jl9DeI5HeD9az+2KMRPJU8U+BfRh
2t0AwkJDAB8Utgt7rb7y9IiTn7dGnPk0rk9bzCvZlV4jcIPUmAy8C3IHvAiFC3fc
x95hSyM2yJKiCki4QjGyDN9JfSXJlF0kwLW5qwgd3XzNL6tlu95nhV/ymmGh3Qvu
t4+n1j7nqSI7yXCcgmu7KFNtI69MxZlQ00yMAsuNnISxiVLv0yvHrhiyATtqJw7W
vavTd57dUx0y9RKc8sfmW3DxKB0TT/0uNVpJN3DKv3HPk+R/g0ColUORcmrMp1Qx
f2QyvSZXIhUIA2Sik18OFPNcr+d8g473ksVuJth4Jf2GH3vspfjSjD2cF2bQn1Tl
DShYTxHvWP3tofQlBHXGNrNA9TmEfsX4GQv41bY9P/1sH+iu25xhdFXwuiL46P9t
RN8pTAuRX4GOB4rEekGSVCu9LjyLsS5s9inXfRFLtedxmDvZEX46DCg1GN33iiIm
X8m9ck+6ciiX22runoenRuQeZJVXSLWBOgxXm580lAHo6coMnkxW/N9hEPIIYUkT
A9IItWEUpV+S7mh77iAZDv4hGaVXRMfXGQ+a9bACyTIGy4BxEYW6uN0urrHi4Xxs
JqTWynDHz/B2M3Uad1qMwkI9Q0IRS4bG61qBvciMcuZr8p8a56NnR02Z8KPXWtYH
OniW3pgXnaLwFC9SwzJdWWcKRxX9H34MmFKKysrShtE8ZeE/fVROfhzHFtDFOxWo
GOH47zqOGCyiTNK1liZSOENrXqSVxPgJ1bfqYUaeHUZsS7ahXxwZKO2DpCw0JYZs
I6yEGTbi8Q5/K18IHmiZ73uCSAMMChWQ4bvbRZ11gBYqcAAk6wdvPU4ynzjG4Ked
vyYqTVnlDZUwp9lXdaSXPYPMcyAWkOnghuC4UgHH1RFnqcAz3nyd3ltyWw20mvVF
GAIgND6DYRyupNIQiU4aIXblnIo82m90GvsRNwc8ui0nURSrbXtktnBBV9YzWNpx
gr9/NSYbJTAWIrw/sJ0oaV95MFZhvh5QH8UGPkT6PwXV4V9OXUc1IUQb+44oHNzQ
EyNyt5lnv7bGEZDg7uM+Ccj+17b2xuEUVYCtUrZdIduN7vIMlJSfs5/Jh2yJRvKC
gsqO+Xzzdb5ML0PTW32F2DUs9MEpD2GM5NmnCD1TsAgDAarIlwMVDgF3OClEAUQH
snG6k2Bj6b3rEOcHHfq6nEiVygYkXL20KP8qtyDfKZg2Y8lxDclMbjh+1lcqvyui
Jk8uVH8FNW4qeQkK4tQzg0sRQDC68a7wP4s2ouALKWtMJ+PL0WMdG7g7T8hkUGrf
qNi6VPhehrw5Cy4oLG9hLePVJN2oRBVb/xmmUMSpLpbPwmAq1/vzYDueeL4pqfFm
ocoSM4m5ILxvHOmE7j6CbGR5uvlDX9hR60mUpLkuv50fLZ8zHlyC8Nvnx6NDFgc4
mX5X1wwoVLTOTelt+dpYbGKgsJL2MxXJGcPXj8f47q6VymuOWYJ5CtezNdGjtI0B
QRdi7TLVASWvtNIcFFJokEPQUjigHTDtEKYjR1t7WGb/BUl/Tr+0n+5y5DcuF/n+
g+i64Yq8AxfuMF20tqEQ++U0K+BDDuIJoPCoX+0L/6Uto+ujAo3lDNDdb1JlGREa
T+KWjPzDiu7sjwQgjy4LikoccYrc2h/H+3jXlOryRGc2eoEn7bTkvME96OP86Af6
Fs4W2Znm8owyO5grQ4T/wsL6keH2koCgGHqD/Pvpj4nYx7phodzCLIFhx8BXMew2
l7KAKDpBBL5KhH9UIsrwQdnCHRA0zttfH24Z5KShNyl0KSQACVbVjdprOzoTTGb7
9UHY1kJ2gtiDRtmcwiq48BPDmV9xo+KMv6rh4sr7rhACuxmYKip80GhuaCobaVs0
NGZWrQokMw7YcX3v6bc/ihkxtELrMFfR/kL3CpmkZg9UfL3t61bGQYzy8XKjuhV7
uxWuVmjSD2/nNZrg9wc3oo0ImPTiWr3rsnaG1SCh3vS4iqukLAuSy0KBvtW/mR8f
qWEc6sxhaUpqiIYt38Rjfszr+ixWr1nnD7PL3X/alwrDHgGTmG3O0bexGvYNeeSn
XTCUT3Lq2mw5/mxGubZxIS7EG9/eZTLaa/155SHhPAZUjP6zGka0o28ZU3MPPehP
9CfB0tLsWBV//G24el3kkYjZ2vcyhuSpKavub40sjW/2Pxb4zhRIale3UuGNRBes
DXPSrLyi3tnWFF1VhDri/zvD1WGF27SjwZaL9kffpKq8NwUSQhqHAbz9zatrXYaJ
gcACi0VDsXKbTqlXgjcdfDg7SG7UFgEjQed38BbIAhqD3xsMQkcM6XlM1bwqrM4W
MhJ91KCBMOOLkbAq3czHBaHCS3B8dnxZzmdZxusorJnABuV8Fv4bp/8+M3uMjn9H
eTFEB3rBRWHQblBDIl7R+z3Wej7EuIuSKJDXint9QN17gp3Hcz1uw3cAjvh8xUFf
Z4fki3EJrmibmdOY0iGT5czPREk9tPYWH9khEKZrX7LNVn5/6OgN8Fu515IcVZ2E
dfgeXBayAXrQseM5isu9Q4EezE6NT7OtHA80Q6IfiqnT1ZFDgZNhi3KxjDMuHabm
cduld49ig3+/2PNv7gl+MEzvzeZj6RkRtLXT39RZSG2TlBi0e8TiIcftJi6LTzpc
yk2beOoRlEtTM3bU5Ay8YwFHcwyql3Unyq3M3pj04LKQ7rUC+iLXwFxvzyhZdXvs
fYpPLddMHWELJoTr2GY5NC2selb6FNjHlf60oX3fG+PdDCunyotJ1ctVwPpco3SA
Zbj06av6bDDH+JgSiaEZ4Z94xvLQ80L9UN4LvItls4a0dtG5LV1qtYs+KMQhTOBE
Lh4hSwl6OU76tt9GhgWuKAYS/yvZAW9naquzE+AiTWrGfPqxg/KOgW39YZ89QjLh
WhW51/pqQCVNCtSfXEAOSH527H8L18AEjIjWgR+/Upw87UNJn6dDl7jpQwlp+aOm
+ayi6iPN2fuppxjzWRSCTosRVXQu/p7p9ie+y5R1Z8vogFeNkWs5a7W/vM35cUJU
pt58skfC3lQMcFYja3vqAF4i6R4jSuy5rqdDB79e26SxX3AlZf00aMPgXogN32kn
UCzZfhNvaN3mLR4gy5CCZet85DRMRFW/05E40KyNVHtI5pCSvh77CAckjIpP9fmN
9m+/xP6vj/uc0mUxo47/W/TtNiG5SPAACYpeQ0HPEGfUcAPgJ22jPKQE76HBjkEJ
itkDE6a4V1ZmCHjMPEgHV+ETA1dAHlP5x51K2pscm94tKMsGTWq2g18YoTHDWveN
xCVx17X9bc8bbF809M/V2ss0LOmopqD6R6q9jNkWpxT/QJZuwK7EcUa/dkTtlM3r
i9hnGRxF9B5huqcYczrFLcGq5yymhmiDWJ4ElKbc20DzNdhtda2VEJeUHaqgTrwy
qnxf2Y8/2HUTFlTZ1RdiuPISli3gTVAWpvlxgaBidb4FeRvSXmC8MNJ4hLJcyxeB
iL9JQ3caUgTDy8pIDrMzD7aaEtmbtL12ggWWPtSl3L4k5lPWqhg+OVhAzpPwQ1LV
M2lzmZkYKwKq1coq7/MXNem2U5ozDa0mvrBD63ZNI50zeJJcvW3dMwU0fU+gvGtu
Y271cMPb5tgEefguJbYUmhUr24VunFSQxu4IA/Jpoz1cnTN5GBKH/UnBh/AMIurU
DK3dQZ1+veYFscHOVSaEY3lHacsPG9Yyn25emNWoCH2xRbYw2n1ajAfhtd10u+Vf
xfefkAFMkqFIGPYsuk2WR+AjuO3awYlFQCO1QQHe9+7SmKOjkhXbK1lpJ/A3TA9+
CHuO+UvUZKhytwZnqykckauwNj4GcMWpPEg2aCb7wj1OIpmnlSATI/CIcbot3L5+
ie6xpLtAEoEMzl0pRhyPHE/4lhAb0JMGpDc6RTOLUOzb7OGJMJ32RvxHm7DYmbiP
yUoV++5WzGxQm7KiwCc6BHd9/OdzUfofqa4XavljEstD81Grw9EcieLOOEfoZ7Nz
KxbrHdWyh2CprjV2scfD85QbneSK2xqDakpgGczBO6XTzvxtyL424kXh4mTPxhe3
zbTv5TF16SdO1Okt3whUFPOQf5tO0wGl7PIHBKi4oZYixG672ptfx4aLvUL5qUjp
sNxWDoGPSBL2Yv7HMGwXpiRZHDtLXw4UpEuSxPtErdFacNJQIRBiI4Hw4ylYokKb
b4l/PhxF1xHj3uEv31xKeMtcaeZm3uxjiUEuv//smSLwPQm1Y1M2JiHgc+sJm9Um
MH9fZIVJPUs6nwmdTrgH7KpIUfMLye4KdEpaR1OiosxFV1n9aUVKQdEPVMjkIKqx
mbaoAUmMKzHUWEoVd077ac/+mPCAp712CDcBKept3nWXbn4BduHrrIESnQ8N8zk2
FJCWhBN3azx2ytJH7zV+7kqmzd6dSwkHZ1Pu9RoYnkryg0Wl/qCKdDR9D625nHuJ
0twU5Gzizb9dCmA407xHxOW58EJK+dAQy7xBAnaxD9Dxkb2ed8APbn8Nw6GeNt3s
ZqgnbP8QMjD2Fz2QXDn3a3Un97c4RmfoNSFrnuBxEzvjP7KfYDh21oYnaeaJZS+U
AYr1rSJHxv1OytHe0gs4DbGl3sZqUxXJkCJGY9VmuOv3LLbxSRUoEbQLxPjQSCNg
5s9hRjkShs0MeRsiLpDZGH+SzBS+6ZVNubF+elqWezqeNjYzvKb44vT3bdNfSsqG
mbHDdvb1f67gYPgiT+2VPjNxDIUOIhgd88N2qjVILnhPuldzjhcMrDIEbYcfGY6z
musibv2tlZCiTe1dB1MEF7NRdDO48F03JbRggcAbtJoXl/h7rncVo8QpQs8Kd6Nv
v6HHvk49OT5coreqGL5aUr6zwI3xXKDkMy8xb5zamTFNV/XrXs6D6RWnONiAA410
zhghADfTBv3zoBS7UASPe5mBHU2+VVJc3a21hmlT6rQf2lO3/85ECZTdJn2OkVnt
/BHneSb0R+ziV9H+wXsQvMpbckHRn2f2m8eCWNfkih/PIKree6qcKnm3T2yqVV4M
ksh5mYsVnYWjj+jNNqv3pUGtK0r3bJ6oJ3ze7nGs386DoKnqy1rPLRiVr9OfyHCw
FnoESkcOcKpONUT95a7+G3x6YbL+ju5/RdoxIJyyhtHD5VdZ282CHpYUuMwGfzlx
OI5RQxZXgxF0Zc2/1ybOekeXwwV4PWqwOt6I+1VisWEP2uud8x8IV6FKzfHb1ELZ
Aklf0Joc+ntQ6TJrTW6QxMXqDaa29RwCkjcxYcLBR2Ws4S89UZe/gfI1gAG4ZijI
M4WFNAc/oppWtrIVrOT1c5ZoCPl7IS1vqzTlUqVUppCYpJB90XOkXH7i3fHNEGFq
8MbpcKrZG7Ptz2EDwYuITkWK7RQipHWP4a9HzO0Ryie0pHI4kRnhIIuxCPDuw/zY
6Jrf4v33nAgxTq1sZRP93wHDCpLGMNSLBSTIlnk7lf9248xK3rtqAvE6g61wXEjl
DB0ASEXCkm10Fsy3ITdZbdshcXhXtTUnJUfzzJWpLzQh5eRjvFCr+JU8ASQqqi9h
gtwYspuwTsvn/o+Fo02SW1DWJvWP6SApmqoywRioW05lcrTi575ycAZiMl3eQbL5
J8qi0j6AI8HHpT+B3SSgoWfr8nenWr0Z646xr9FdS/8hS+Q7RnaKtqz2JpFpRfqW
vpDjJ4WoRZCvztXvdTmkthLF5+RCsuQfj+J/p7B6VXi0QkVx9KTg1vPre+5FS7rI
Ts5014w8GG8FR2pPzwz797pLEiVDnL08/36IEK5bXvd1V8WdoPM1zw+5dGSgYPv7
L8EDOY0M2zymWLLx/CGeasDNUiA5ZxqthWVkJtgVA78LikYuG3Bz4VoKRjL+vAwc
elPecI3De6CBCU4fxkyKOMFa21/lQJV3uPTJRCwxPrzgzIZNlxiW5aQkEWzabztD
cbVrxjsRW+cO/+9ysDYSsU/fpQKtIIcmcaiYBMvqetZLEmIKdRLlVcpiC525dv81
VZtx7Wjaq6wos6BAMzLIObF/wLUNcxOejop8FGYga75R/9K+Jl0iYaZJ5E78Wsoi
h0t7qhr/TpATQvJGVngjjJbnvjGK/BxKhhEb7lpZGInXgW1eFlxbu0B3PXLNU5vw
x2lqRRU8w4ZmWfpjcSf9FAKGI2rNL/bZ/Udpm4dsdipLQC5eroBrIRCT0iQKvojo
cWN9phulVN1gLs6god8v3rCrHXcl9inQujjJpAkdD/Ekg11ltFDJ+xyQXvTqWelo
5LCZdgLRz4qTCEjf0tueLObeMOUDM+Fb1x8FDJ3n8xUClxKgR1uLPYS0AmMTwQwp
WS5nqNm899Njw9VXXYkD85Zv0qE3uPeeiXroXPe0DkuHQFZ+mNWyIGBVRKs4qu9X
J3mSFTYJgjM3bBnItcNk0v6f26vN4WgJACYq9O+cOfl0YxWXCvVIMQmOdFLdZ/4+
vAl+xcmjjGMa294Qmnf5PEKxK5b+OJEGUAu1RlRrQ8I23xb22Onps0EX0629qXsG
AE6x738aJ6WIzd1vIlPIvUwiZpxg0OuZJ9Zigd8TXXF0io6X5YF0aRIPeNIUm/IS
nJ3bYYZoe71jjlHHHa14Wurib8yW8P+vQV+EkF8tpSTRZVM6P7tWxKyh/E/FQGvC
fspJjBbsPDLi43msKg33/XAIw5xEMHFWqjJ4sHmBFf6iApdFTS6Y70qFyUEPIuGq
xJgjbHsFNqIFA1JRvnahtFphrbpolij6IMI/mlXu/Hu4gfFoJEWrV1+HVO2e7UjS
MzvfmJQA1SphFvLT2xNzYUHUiV24D3F3Pnq3qXyjECKSBWsPLSjeAa5avVn5AtcS
OUGmm10fPQ7FdPk+79Lb3EYGFRqfbUZLoQfHa+murEHENxQtkjUF0YayhZf2aGN6
QG6VeKXmQcQatq2uy65q1kuOtKpmWJmHbDFnI7gN96PCPNYFSLOWVUG9hvmj9jF6
PJxKV+ETmrH1ZQasP8K0O2TxbEjL7GEwAqcdamIWIFBTLlwxPdYB+hYezXrbUYdw
7HFuXCKEflvq1G1YetvsNorwqlqYPz4KjmgsuWfNbRs9vu/BcdzAAY0lxsFtwMaF
I7u7LjHQdVXpG/jOdgd6bxV/qTGCgSTlclcF7IYftpgpkOYxh7wgRiiyEagJJ54k
Rj126UqTETca7aFXKqOjNipTsEaupsOJvetpAaKwxcCgRLio5NQXm2FODq/4lPwO
QF8zSR1v7LB7d09jvGRtJZ4JSqKB6Meq5DOoPu282QUYQNm/V97+UlO2WHfeh10M
wiSAIX6f484mPh4skSn8q8POBSPmBik4Ub4aPsdBGP1wewJPyidWELVaUSxEz3mk
D9Vd+GfcwjiyXafYWTeVsqAgtLJX5ts70jq0IDn9pBxaXn0Qtfs82/JdBQbjcEBX
RQbigIJgI5k4xl+WREnXNuhpFFYoqX7fSOT1Vo9tq25L5W1pPrCUcs+gwBXP9Wu3
a30iDsQns2N59xKuscH2jL7N2X6jZgqcUEPZ9cVu5THi6/I8sT3+KGKiiF6eyS1i
u/l35efw6yDxTtPPHoCEpVmt6YQBxkLae/UhJ7hh4/wCeOIkBSqU3fjdHbkylDUr
H2i3qohWFxza8IpGIVsJ8+7pikQfuJ1kJmFJYkI5hwDIhMuYdHkqkfHCM4MSlFXy
hK1WvP3hhqIsCq/dFQnvG1rj4Iw78LpAtJ+jfcltZnaIh8vWynuyMhBn3QxLTFCN
f/cs8MtdqI72ZkcNj9BwuGxAVTpMSI8V3pr7mXKTdAGC7HeyMgVJvk8yrg85Jg5P
8bYzQYReiKZ44+P3eDJGw3rTkJxSXouA4QdBomeqmCgvmwAlz2EBWjHf8j9cjPVs
K+fLF8ChUniv3he8uHTGGGhuiEyrNsrg9T+g9AWm5Ccjw9bqiV3hR/cuMeM6w8v/
Syp82tIlEOqE6zSp5/2xh2oAyzbm5ImvDxih8Mi0kOONoglGm7677WTE1NDYCHo8
o/uUFIxfe+Nt2qNcfPgvarrLxJPaO5AKjXJSKKbVisS/R5B/ofOJVyb6JD9DnTRd
3SdhVf/ZW2atumXp8f5CkeMa5ytDfPUCM7rTnRcHyCVOEoyH/Axji4wkepc9jkS4
i5Glach8f5NTJRth8jDo/DistFsOdJpsErMfL5cWsdDesINuGAxWOhzNR+RAmQiq
L4q/lfycHwz+XvIEa2nKauqxMr7oZNX3E9HW3QLW+Occ2QLN5vJONw14Dq5UPn/V
s6ozUWVuCqQ9a7aUDjFy+VGx0Tn5sqRh0SU6W1mLC0WjDJPIDbTB8HSr06RJC+dU
zY2u4l9JEszOZ4SrgAPZnPyJjp2GsX728QyugPdVO7BtuiMY4ABEZ8YVrsrHFMqh
2oFo4jqtE7zf5QtNEmjJrs/rH9FpfdPMgM/Z3LJzL1aAnZr+ZMUjX0CfRqTZDuk9
SJTd9lXYBY78NNkKYyhQ4eC1JOjecxaWNdG38FiC2t7Oy79rG+Axl9GISlEm9ZeX
M4eWasxAeUim82vlqGWmuddsYZhTvwN7hX5OeOH4ktLWQf7WBD48wsSpdAf+YDiz
He6b8ru6KJYeN4NMY+6ZZ8dHbguZnoCbHcw4Q8FcaVHRBP/5RxskgWXsSbZPnarb
b7rGRGGJHd9Ik2eG6hPdX03agb5Y64T7WF6eDV9rX9r++K+p3cdaQmsRgxRtnyiS
pxol8pCymn4F53kAM1UE3ei1r2/5FAvzJVnCmF315Jwv/cFeUd3ak8gfbN2K08l2
WqdZixpDoJxSxTVH1Q6ynJkLkjKsEn3kz3JlMi1tGpOAx22wrPyrcOkIdV3grd4B
mmOay/j1Xmg4pdBlr52L/ZxoIMTc7dP3vRz4WldUTMVQPvsTfqmxoYV4L7hAhLeB
lYBoaY420cmRJj4hPCIdQPAtNlHEdmczcYEGiJ+YF+MmE+c/nBRQ8ij0NgSjiP9b
viws0tHNZxewrs5VW9yMq0CsEvFSqyuHRSnyCdDl1z1SX1LOXdSWz6AmPGb2VpEN
eTQtBoNQjbmdYfEwU5FoOTQAYtLzKKHN3fupcCOm4ks96D9jxt8XZeb3ZA1W5su4
v9yjLhxOcKXfWd8ZpYo9oCft1WxSr2h3CSvAmG9wtf6o780138aZlyZLeKzzUrTz
E1WzV490dj5bS+l+LB2i431UraDfxdLxAUdDD64RexzHpZXqgcTliqt8QZFLIt5j
6AqvuchNWUGjPeTomovPswSAeyXn1N62BbPssaHsCoShgLxJ3X9bGTzbQNsUH78f
vR7iiN1RAaWhVpimrykaZ52LMbRAIiPV+2MqcsKkQdrO1hkIfEYWdSjLgXogvVbv
h0Bz0PrH3Sv54pH7hns7ME5u4NWNsRkP2aLb/TSWI4SNKlv5PU4IF1/y7aKCaIa9
XTe1VOWPFlG8zu6fp7ibRN0y8KtsekpIZO1zL3aE/IDfqu9b/DTG1TEHnxpQhJt9
+9e0CKHdSZ4q0DnGYho3M9mzTFYOnryEX3QKUyyvLYT69cWga+cw1RQNhgXugo8y
TCjUXw0Mk/pyAebNqieAm2aCxOO6mz3Gmgmc/GjQ67O9G2u1hp6s8u47EHYDvU4t
L5KQvFJJtATCG4GxP4j2FwtdMyiEGzTyCVSJlefU39RzAn3fdNn1DGG88TQ5faNr
1QwfeJL8FObVrRbDMfu/vcqsFfxF1D1rpGgZKfGZekvSln4itYPViXIhbaii7hDE
JSAlvn8BdRTk7qhqB9ROM8aVI5pqMUoAM21KaqrfB6X9SDwwHWiBbvkwLFfj74mw
cCgU1AM9bl/poqyau31bVSF5505GAAZJCyIr2gQyyabzwyTgjtZKFwLHNa9liTPi
9BpxsIuugsAAuF5GjpICMaqZEEp0/e8lAb1/86tuo5tRlrBwmATNFP1iNfhd5vma
JeAUJdUddEanWyoPFNCbnnhfsQAkzjYKkHL8b0dI8vpUl6L3pM6UECgl7VrBIARx
3AipuREhtNOQIpjc481m/45etHy1lLTq9IXLsILebaBMtzXjlZU1ScA1JBiaz/vD
8C2v2hZ79G4uoro24jQZKA6C3Qv98GkiPCsFQE2p0tAt1GJrTkvjj5A6Dd0m0e5J
mBsDRlyu+m7IEPkyOud5R8wkuBHENTSdAUsIiEdtjdhvh4LfOYgiuEvukz/xNX9C
/VXRubIXnn61LZ/9YG1257BXhz/fF7G+xXPI+o5gL7koDqfSC/XEi8MZa2t4URcd
aBRYCQAlkWDeQ3ICy4kCILca/wXEvBj5ZdHMXyVGppNh+Sbrg+jZs74sRM7pSsX/
J/KLmWcK+q6cDaPKLVBjyCKS1DuG8yIuFtwp5DV7gAqPPsoxHiPIRGfSsZFgyloB
zjOwZOS+HOmyiUFKlP2Re3OP7TG4oYs+QxOVGOtjIVgJuR9N0U2pD3/cyJ/VKazG
C+sjeh5T3IZU76iCvbMhOZaXwS4UJOp54QB/zBI3VsT4IM4rMzw6BjgjjUMQC3Ms
win6dI5hE5N4JG0rv0pSScB1wENHCzqIcKYt+CFUvHuZ1eb1vCDBOMILYCjymIcc
jgn2R86hKDHPEHTlgYhHcYhmN/6YV8t32b8nNFGcXl6om6ctObL8UoWp5cq+cSuB
Kxq7Jvpbxb8pX3lrwYtzBppqhIIEkIeEr9TwdCyU/xXck38mSN7eZgFTkHfSrQLa
76a+D4f4WvIz5ZNcDz+rQodycmGhHnGt2RVGHs7Fw7m4fsWjSAKdnjrdCPHVGnvg
x9XYczz+nyqim8BFTCm6A8lAIYLbiFDxnFaIeleIHgmZ+qn+I9KyqXLw4PubSDPC
N3SktJa9SuPcjzpioI86vPsAUlxWGeRlzjZ+6dosMySB9vCAJqHeSNHVJ0xyFXyQ
zqob6HTA6ts4VT+IZZmdN48Dr63q2ip24ag7Upb/1s7ya9iHbCuXWJi0YrP8rg1Y
I6shRvlvejWdCnVykJlJK7eOtfbcrDtzBuJr/x152fz8FlTfCjGePyrEU3ZLZ9s7
rH4nW1r/4GLZa23B1RbUhGFALY8qnmx3C0AiNBR8+74bMArXITpGeZ2t1CTtzMI+
R7hqt1PAVtUYVS1t5I8ybXQNF7TazVcL/9oEcS4e/SKrP+YcYcQlSmTjliJ+afrf
MxI40GzoUc0/4AMsJriNYB9vYesvO605qkCDgnA2LfcF7rPO98IIT610MiMftCf1
wKOcLdyflm9UGASfmNbQEXgALBQc39uFd29PlGw6tUgFEXuVRzpb3bgjcEZOcekl
Dd5brz1OO9kPhEH72fL7DEpGIvY6TAhSLFNJpXfsZJlzNB8umXwdC0j0s0YqTHVo
ofkr7VbA8g1cUQXPEHylMauV9HgdM8m/wcNNWDk+FNqCEojSCz4vmB0g2k8yA4Lt
HK8dRqe8DCRRK5OiyvB/jsmBe4N8ioWnNwbwFOqX1WgdX3NubgHbxs//c3sThSYS
/n9AFqQkMm5g/iNqpdQ+4Rs3gl9fccoo3bkoob4LAgtofdm+MR/6HYNAOk/gr8Rp
REznnQyrf/pPK7qXUtLxpPVK36bnIiKzx6h8qzU3PTB8S9MyGPs5vsVk0qnJfIy3
vCFwCgrEIGMoYKjBXabXhcn/hfD6eQ8aSdLjYrtz0hEDlX9SMX785nnOWbOIDGp1
qWXsD1SLu8OW5JJBmIOaiR0ycvBZln4nbJ5Y+TFbgb51f9mhZtDx8Fxh4A10obsi
2pOyX6di0siktx9p2H8pW+Y0s8lA7yERQURDFxYXeuBV6SxSsutLFWKyALiEHe7B
FiUWSk7AUr64jL0736HcShxTEdIg59MNJtAGd1YfvmvhIncFInHhK56fmwsGFasZ
yE69CVHNpJNcpF9DHRY1t3eWWanrJkrWeAKctipydmesS7/PrZlErCZCI72oazdQ
DRT+VdJgnZpTEWnLkhPXrbtIJUR4twZC9GRVy3kd8HYEChXbzSbVMPEwLA5MBBsu
HUysZELJMrtFlqkvmgThRPjK3Cg9d+x90Jvzm5pU898j3I4mwvUJFoWQUwh1Ry6v
wCIfDJsRWJ0kW6TGxtdVrh58W1vpn45Iqi9uotH8Ew9CqPTT1xPaTmc9Eoz3eDBk
depfvasGsl9peCLjGNv4xJuhmbqPPVcDQW3GHVJ/mLr2QrDX3NjeYOJeAsf8I5ub
NBC7k13KrbQdfLod4oxJjcU6AA6SzMjjaQ//XBh1DwGyHFwyVgwzAxTNOikqUgBB
yV7Em6vF2oh2hlwneQ7fFo/hcmVzAp2WzDmOin9A3Vyunt1fq8JLM8IGO8Mw3fwD
VOV4B1xfDmKiUO3cYeVGt3Cit9lRxHYTZCv7vpq1mdafjDTQnqfXPxTuaq4yn0JX
V6u5kslreFVW19BXMEF93Et82ATkEJbCSDmsjXXfAQGVzVGrKfzvfBaCXvfZmNIx
edvmihovmwG5XYKZ/Gun61R5tgXRZC4cOQvN9MXgCHgRtWsotnYI66waOZ2L2by5
EFoQIybsHZHfvL7phrSVxE52vWm8c8jvdi8U6wrD9AoslImGlONHXSnMsOtUuXqU
wSulf3Z7av3SIz8u0EgLvrWpp4iDTR/hU1Pp9J5c4bQEYgL3q+dywFdx3FeHY7iX
PINfrErLI5fevQUOwoKoArgKXIDuUnGcNFwOs0R1C2GFZW++ruPmS96ST74/YfiX
sfIyYtVOpR5an0Pxd097KqEC+eIjPECFY2dtoT6dK780siAeiDIQWJRucYjI4iFy
UzT7K6/cNFhSEUbKzSk3wy0mUnguEgUSCIzROfnGzylnd4Y1oq9GEOyvaK4TrmjQ
xwrMiDCemB/fkagaBh0buW88tpYZumPdStQfRvNhgKASxQRA916OK3J7T+TbWBea
0ocg1D3oBeRfr6qKiqiyMREISOaMwjR/0WCKT5UG8yen6WesroKCxNV/g3Guc93d
8apuEiWhGnl2O6Ru6DrkHZhvqCeXlHXGnEYCuRt+DD0+U8uoapfHpUWcs8X6U9it
HYxCNbEQjlhFzh0zfplECoN/A9elT3Fm8aK4G5kmR3+b7Sbgz8NtLHtXQ5CtoLfZ
3u/sP+7bDv3XS89GwDs5G/snactXHN1WkxAQTGRuuJlMLf8xoJz4OflW9orWarIc
oXklQeVi/C4wCkZ+09YEeUQssLqj4APPkrCCPRX2zzee37b4IbYk68ia+AYWvjvz
+vsV9zA0vn60otftZZ5iBw9EgWD1resxdHDjlyRgQEplqsAqLHGlpfUvhSaXw+aO
5jW2N1IhyQjliHqZ9sC99aOz/PS5NzvS+//OoNsrONlrXHbIufXi07i3m8Kb5lGz
mhEUBhWmMAB3pEIqtoQJ6gK/5mm6nWkg4VZbRDntGYD+0y3BhyYQbw6v5bjxsbby
AIulb4dPq9hNfd64ANZOdrAlLT35UmKdI4NTvJOaPFyjLVf+Yjxh6xufABZzOxdn
34m6UTmYmiXQcs6wWzAaCui4PFDo6Vmo3GfTSkCHocwoHu6cgGqsg9VzciNTjh2F
WiWKTVtZzh0bo/rpykyNXix1yE0PXjd5oTox+jcUVGExdyH0LdaZViSRD4utMqDs
2pkd4SJRRZr0uRxWWjBIFceSClz1Olt/5RUE1zOoj3APLU0qd2kcwNwBu3RFBSdc
fWiPiWOqXlFHZ5h+fv2N6rqSdDCRiF52JqzfYhybbDmgGv5z3j5MPOXg3PHzJwv2
WkH1ASgnFhJXwMaQRYC0PVToAQP+wL/LGse3bvzojZVRJiZoyOgtcl9ZIqOG7kye
SPY49bCDSkFMbOFZAuVwOiKJXYOKhG3jVxKlNEZW2+zqCMFo52jsLbbwODdb3zlk
BoRtMt0Y7w933ACufbRTKThoPjdk67kKmLQryHfIR5wqFldUYrxfaK78bkPMsYv8
2FAdYpEudDACw/iUqzYkqaRQlxLpGaybrgr3InL5ZcXALYQA2gnaGXA2811Ki5OJ
C102dHOdB9Ckp70krDBLoac+HMw7uJrEksqgfVU4SxEPQk8oq/sWNakPKnPsmIR2
QGr6zoUXAoNz1SL/jNMamPKRH7qcjmwPGiEmxzH3ygJnoE30DgBj4+2VmXG88KlS
UxjKqpkPmnwzptZ2jCD+MbzkJjjY/EmWW2EUXOB7Yj7pI6rTo+FQGmPIDySwN0Jd
KMTYCRSiKpSGI1Rqx+dp73/49pR8yHoBp/zelpsQ1a2H7kcZVmTnDhIJsNV/g7Wb
dICau9uN0MvR8r+6mip8+8Jba1hPIPYSy8khueOxjOr+pgNyGFBX3s1QkVW6iFyX
X3hf2JsBaX9sJdsAsN1+NsqSvhUOtT0lGw5Z+eHAdSlIqR6phFaeapZKZrLBKoIm
nd/c3c5LKy+xYzMrI2Q8/MblF8+2Z1w932sGTv0K/GXaJTE6XSCJDQPu9z1p5efU
qCkCkj43dtnweTi/EyfWHY9VtwSDPwG3aolx52jsdwy7oAs++kqnb2+PDl1MR8sh
7zrObWX2K8pMLnZcNXifSQX6m5hjOQWfIs3qbu0+2OIdINS3o06QKsD+02fvpeXg
K3u6ERtkP9ZB47Cx0IdSwbGtLXxmr4p1t+qyFWSrLRTnDQXgO4oTcY6aV/4KxrEQ
nEx67YIgUF6ITAjIZKJ+n3KEDetcw4qGKEuZp+UQpPuEsp7zTfDnLNWsEr2FHkdp
2kdDM3/sfPMPy5A4QkT8/dkvtME623qXlynKqB8erF49TQnhe/DLNBfVlwn0yxEv
6gzQSUyB5qr55OslcazeB9dtTXlKYNH338bj4f8E5/U9L4GRtKDOy4ZRstwgUEOQ
JyUp8UlPZvc5A95TFL9yNSxHQkvxNfmGeXx1gfoKlEjFeBwJWNAhIlDXi1EkAt/9
WN+XpzAzbvwSv4yLcOEDv+ZuF+52ngCoFE1D6bSv2lcWmIerkP2XaIpklfMQoMMp
v9mqGc4wCytUQJWCRNptpTzjq9xZ3r9wAkyvAd9YIKz7qsH8s6+75Sgx9dtOcF8N
iGD6Ls2WkrC5QBe5Td7zvgTiWEt39TlPJZSOl3fK94pHSGdKIEahc9hM3aLX8slm
yvw5jwDvf5DwrhNI1Z8f0sO0smRmZgHPRq8qfkdusDQFFgCHvGq1/5i9YMvVFPP4
ZDYaLPsmu2LYlB/jRvdXB3SpD2JYC9/Gui+/RFKHvo5emUomjiYr6dbdCwfUlKzc
MVVt75zwrL6OFoG1/P0hQu6UTSoiu6Di8HJQgAemVlyLHLk+qiwLHir5Y+exYYje
yxpIFBPuYcNDiT+RFHHBY/hq+AUpcYkr4ehxJt2yzXupIQ0Os9vVbYDxDzM7ijsJ
cD5406PcshhW/XdlydtbMo07l3DEOQNdFSPh2dsXcalIhMNDHl60kna2Dy6CoccM
BV8TJH3F/LkTAjrQp+cs/8aCBhnnRTKc+10bzsaFIa6BDJ2Jyc8+dm63ft6+MisF
/uToFJ0qBFVrxvwaet5a53cLrF6ZrTrwIFNZ39cWoOTEhOF3FWJ8K43v5bnwT+xd
pGMnbpedoMpA/9WV6GYA+z4kdmy7rM0I198c48zN4ASoHouGi12NjGIDSnSEpCIL
cEbLy3ICQ0aO+cD6p5uhXcaQZoXB9NIaboW8d3HKfi5Mha4PcHg7vVnrXdpT3o3o
GfA2kivva5ks8RNHvjG7nQye9hxO506PLJic1w1wsmfAPQofvcwZBZXhqCER3lIY
g5t6Q/6ujCtbfb2bBUN0f8I87RA+MX+MwwVM7fb7iNyRTEVI7dptMgAR1LZRSpLX
6ofTlSS79QClg0qZSAiKngynJU/8oIpwBCfNnFHdmrKGtiyFlVRWqVghetrfq4An
CzTdVKT8h9nRdpN0cWrY2zXKYEZPvnJpDzSpt/tOe0hPLpdN6/CvRoeVrZ3+A4Xf
KL2F7j7Nf8ULrXO0w4VX3CXIlJaBVkwyst5vj66Lr10JbVomIdMsFJe9tEn56+yE
7ZpOzVqMltwgdwvpUx+SrrH4N5n2wzyfVlgAdg3ULec1o+9bPw8Ln9GgG8Tc/TvF
3i0cVXOR/ovyU1Mo7WycjbftXWndz+RewH7Y6FUqg1eXxoqOhkVx1Rb+HkKPTBqj
3hlBb7SUCNoHsZaqMzFz1kuAKW6jNbqU/LeAH89RendgH0bOqz3bh6ub29JxQHT1
HdvJLI9BfBP3i1C862emMwD33v9Elh7ULuKQCF8ZTdtgaW+vFGOF9bbuhO2Qdun3
TcOOPLFCPqP8wcdfdVEjsk0EsgxZqhfTYAP+smHi9rgbBwPbW6i7++tG5Z/3exe5
x0YiMj4b0B+hNxT3Fpld5vyTr6UMwwBfAcinxBRcm7ALg5L8mFtWDLcUHSw7SEOa
WfbXicRI59xytGkDLZc26wC2g5C3KeETIE985jaNfyJoOOMlDNXoH32ANkIjIMl1
W3gg4ocMs/VssLTIbW4d3CDW9EICBr901zcyA3OBxjLo3vUDgwT0WQEsywTdXKxt
slAoNlublPWnRTy9yWL28vL9rvWhIVx+YMpM659mLpPBuO7kN+ApPBmded3XusK1
WMbFXThKbU3h7ucWWIUcJMRj5eGa+ePN+IGgqzIO7jV3hm48jXs+Zn3/bcrlGwBH
GgaeUYFDGsFNB2s1IMKlvQXaBG5lhtnbB8uYDxz2JJJFSL3hHEr6DhHNF2zmJ9Zs
ydlRa3Q00MLOsV70zG4/hqfMFvBzEEbaAcDEDt9m0r53IDC7fhXeo4Dps8lOQfi+
rlFJIaz9jOSVcDjCguPvDD8pru08LB7lBVgb2ZQ3aVfVYUTEu/YQcRiSbnVaHN5x
yIDIyzPBJwId6ezKK7isLoWAijkhvCYXwH/PlmW2nrx0AFHJT1yQ+7nrcMxSJjQ8
FxcPmdmRqWbAcTo+GitNDeBN2jewTCMux0iHwBq/myrOrB+/mCjncRcfbhmTFZZN
dtuU27EmH0e/R0tOuqPgAkCMPPfewun780EI/BA9sS9uDWGgxyNLh6VFBawDu0cU
q00ZjbzNoDScBEscLoMZ/7Q51m9DSSU8JV9V8eUokUILUJfxJd7uA8Ms5B3E6hvI
TnVLYxFJF6cMGuOkJr0IKSBPss1hJXKXB8PaPITawvRtO1Nj4fZ4edNHMbH56MkS
71jZGojycnqHBeSlfs2XALno1X9ofm2pWKPulLjDU5qrj4I5YreXHkJinN+4IgoR
/6zXEU0vpXdJQpaLziSOPJkzcqvZITWITMO+dIVWYNrm9/H6WYAQl//yvKpseVzo
tTwVwQP4A47MGxR5IGKufCU/Y/QePHe0tpjTKevhAIAn/s5ltN5XFWEmL/1ohakL
FTgk9U1mCQsCnHu4smDN3SFi5rAAmS7sTUs1w1apjTbhsznF9KK/w0dptga2EwzN
uBP4QPFWqeRVOnr5nTQhyJFCvqw8qPVg7vM+e0CfJlyG1vZus+d8k5VykGyV2B4C
+9/Zgw8d9cDWVu4UywKfTpHli46/CPsfiAVqbxrUjMhaA9POMgsfRY93M7jE49JB
717AEICcLw790HcKgBWdX+ToByHLrai5bbrpnjPFMzdu0fDGBLMchtLjiVAObe08
4JM82xe0NtyX94qMy2wrLCIa1s3ikpOqe3L12ZnwFAEMvl9+ngEwL/MVS6xwLPyM
cRYL3S2Aj9eKmVBE4vfQ8JDuM5VwROryS3c6569hYrWxjck+Ukk6rKCmawFKiyyV
cHpnTwfrxbAhLSNgP0VCSWLK6r3YCZEiyRDhJDmofvZUtKDXoVZhBF4vS6VkKrwp
XzaRN3DM6ik/42JYl0rzqVJ7FJMFueN0T+qfuK6uLweX6XxZyVxq63AnBItiWL2F
6hLfkLs5muxzMW9MqEsbXanZQVMr4rAy6Bi6k1seYn5jfO72OnJRghVgpTjy3YdN
tuVNtExKLipn3ivZt0Mt9gI91dBvvTyRF3PrlAKXgnJae0mQD7dXcvIHt8K4k1Zb
mFGrHB4Sj2A+hohwP1wpyEq2+Jt1mN6v3Z+QW39+56djS6vjkoVx6GtmU7wNBER9
GCWdZDpdtKYt5lID9tFHuvFOctMGXe/ryp+KNcNX7KdCkomggPFnxAfs1iNfAKkA
Vau3GZlr/vrgBj+AXOejJqAIQx2xoxd2NvJum86zf2iAdOz26j/Dxs8R53DJ3B1+
eH2vrnJsaY9vL/B+QQaSkrG0RrB8Mq5G7ZQ2eWvFJkSLsSGFSLVPp8pjBZEuPHjP
pIoogZeHQNGb2Q+3FaDAit694RbHnpac5bSqB1Osi5gwdMsL96vJ6xR3PxZ+D2O6
WGSfDjPd1cBR4BghdDNuDzm5W816jH9Al6b0htCuxe4y88CReVjYbtvZa8ymhKy9
wBE2bKmpSzSKoHLqko9KDaWnyOhXa3zDIqET0E5pB2OXbTYQ+F8PoeTOsMzs9DNX
QBq2Khy3/bbUFO2xKCtR+y2mHCBIOgP9APvWq0awY8JwiI4ZaKQHokMij5+rq6On
wlgNgMJ0tvhPHkt1jHpCbQobVaDm6J4FXtIS8ASzvy7nMaRKgpbak4v5dW5Wyy7u
pnuS5AEi1w8J4au7K91UEwgtQ6hBsgdkXv3krrt6BJBjqefzegAbVS/FyxjJZ8RJ
uaB54KQXXqiLM/RFAlNJnxEOLFHW/nRtQ8C71QWGQS8GQkr51sbZT3P3kbzAdQIn
dvGEkl5TCej7jnd8PAZb1juHu+jyb1ALLWk1Qerj93/Tfj8mp1cbJ2t3loW7FWA1
ipd0opFkM9SpelD2BlWVqEheqK/HzXqNv2wq63HxXpMStvfdWyrVpizAjGwpklYL
K9NcHowT5hGgcJCfxG3Wnqy5Gj2uDHhnTz83RQh2F73OpQednhF/N8C+AK7EF8X4
uPxCImHwUszMVtIvGu0GTq6FifI4u40PWbWX9r/LgixVmo692K54UKobw45B4Lqs
QAPIchLMKHCvRSE3o0GpTxXLcI09xQP+Sp2MODmFRtfmf67KTQBvi7aI9S0Y7jaq
oeqnaEFSNFgtc6VRa5dJz7NnWdb6pcJ+4rggwvovHZsAQsaIGIGNY27jkyvjjFWT
3C52KrWcfxNHQbP09KSyLN5PJxBwU2xZfDFCvY6JoSI/lZN0R1YOBy9nPyScceXO
21ile2DKCr5qpZd0kchdcBkZshneB7gimx0qVVxclr9YmTTjqR8Z5j2h87oNtHek
im8PlgKD4KrlIbDeapny1l4xX6QfPDxzjF1nyiJdPiU4MmX1RuGdxA2FMnSFzYDy
QQTo7JVE7Dy/ZILvCHmAJXwugYyq8RmKleMzt59Sz8UvfZZMpr2NYl/55EGksl2D
q0IG8/lI1vWZSt4N0JDQd7Yk2/W/yXm3GqG5SSDNKuU/TYQCoTxB0OWv/Rp4jTVv
hAk7R3gNlNs+WVuYZys4vBiT8hgIbgdnzlumig6AW9/s/V4XQc2FpGQuzN+ZRLGS
Am/YbmDrPzbJLtS6VdTsnw+TdhhxG3rlwotmNuzZYoiRLhp2jwS/SrlCE55Z9Wgz
E2p1JsPkDo8ocinvQVwMUKH0JX50hRzKsbBJI2YyWiDruCepTbJsSX8A+mUzstIP
IwH011ADNRyH2T0iktrhjBnn0ysi15hkX1tuxGoFtq1lexXPkrLmuL4ESHH2yeyR
fA309/JRB0subPYds5LW3RT4E+cTivy6BXv/IiecjvIzKsqWOXnXYPdrATKuklun
V8m75mGxlVgbNTl4hvWTp3m5qVi9Z2aO008GBNcI1ZYfDjsZSX4YTIPpiCSlHZCp
tJbdq83FhYnpir+Wo7/ykoc+ggTnOoRVwLEzX3WQdubUNqkiduXk8kaFKpjs4KvL
+3OWQhVqUc2Y7Y33dcOb6WofR81op8EN0CZGAB6k+s6SW/4OyEOJOTXa14dwwaL+
kyDFPYnPkidnaUWfHPoJ/ozgI5IGEZs2RR+fVQ9gaWiOj2IsqwHq2TaXeMGpt3RV
WCFGdqBL+lt2z1hZwxhc7xeL42CSedAzlNZ1ZrD/vcYeZuWUq/GQP4de/vP5AwCh
WgOz1nZxB5b0R3b5f6x6gZZ5x80ZS+m8DFzE7HrPTQ7IcLsnWOmTW6P8xwD4wRDZ
g7ps96/03jMCNun1Iucri1yea93CJo82KCjcyZ2Vu/7CIEVxk0wq9biNlbxEpwm1
JcqoFRj64cIKWF8hFPyPYBQqz+8OJQABckHI232yb/VsRsZDq/nj82E1sFV74r/m
WxHmg0UnEv3Lnhz/U33PIifSjrR6VM0ve8G/zzU1yxQtjylgHVeQyJKk5p72RJM1
sbqpnz4gIJGj/1c0nzo8Ywt498y5SUJ3lVBMxHqXQMfSx0HPGWOIsZsraw6X5sLu
PPILVHRlsKu3vm61N6ZZpNKoRaLzy/hqjYkpcjc4risn4l+jkxGik7W7nVA4p8zO
X0qADx1Gye6Ovk1C1aVXFDfqetOZgX1JSNDXSxG9pEKO0eXar4ku2bGgFz2O1vKh
r7yFQHXvDWixM55+ggjYoYWvaDcnYlwJs4CRatJCy1YptTDSLIw9PKoP9kTn/l6b
fCQgiIGvoS4wyVlnUgPj4bvRRSPuYEL8qOPkRX/tqyx4pXgkfiFUXYHAHAB+F/a+
4RMiu1ppVGo5xzsUnrc0jjoB/srUpl4+0mqgGuC1DKgtYiZYgPLpuw/joPbq0l1E
u/QVoHWdqsVqkBwi3fZGAbgwyBOejjIChoAZLMr0O69nalqTLdf0Bksy5WHW0MAS
N+KBNULVIIjyJq9aIIcbg7GzlzCbo1JHuZ0L+Esoqd48detpAp7TCrPU5scpH7Db
exEYK6yTC2YwCQlVjDowZfxzFqHWMnIpyl88o+vK3WTxoKRXQzYyhOofZ77mKCBI
66sJzpx8V1SMYWfT93i3RlnFiswNVw+xwnhVqyePuL/0t3h1RU6UXjFoK/0Pwx+3
CyI02SDJFrWmi0ewdenswSwvq0MVhMEc5qcZvpqFq5MybU8KywerLU/aFFo97hO4
iutpIaa8GhhTQsgJ6n0XQokB3SljH7OpZwxOz/tgEHZHPf8WciBa/C98pI+egsSv
QW21dQT0nNleWsq/CIUwL4zHjQe/LImCin09hVsc+SQ4DFRcEa4ax00U3cre0VV6
BBunoNPHbgdhPhjzDyD3GpUgeDT0RkMi3DhG4NdXcNkP4YryBbsX+C3JDqmZM7nB
JhV9RlFzl9RHzzz+UMxvkOmVm+Hdf/QmlaeeiKacjG94/3O9zK1/Bx5VMc2vzz0E
zBWxEtx/nSTB94O3PvMAODVN9atA4cKideI9Z63yuFYr6cCPqi9lccimpw/NhduW
aHuybHb798WHjF2sTP1GtxT2Ud8vCRV98RZTiATtmIT9/iudyytP6UUIfKp/zXa7
ycAvVYwXPP53/xJB9OoDvpGTPs3oseKEx40RTSrRwotxJRjGLj6M77HZZYhvrJ9J
vKetJrkDi9Z8t7mvDt+/4h4ViCZcBwxTL6aF5NJ9DWRBViHeQyg+l8rpvC8XCXyC
KNvq8Ah+9MifahNYmjYOOuIycxE+AY1UlnYEReS4wui8qQXCpANIRafvSRXUyjLd
/q7zM7BnLRlhIVmcWDm6ciNOLMH7Dl4IT2e1cvbgazhwmY2op+YkVMwpmwIBKPZ/
H5f/ROZBjxfQ3+IESoUZxzFFYmGoKptkCDd7o+ZHnDH41c5Cah/l8Ho+0IPMoEoS
auJLP9AeNHCxIpEK+7+QenGR+FlgweZHHpXrcXBrZGdQRHoGK6uqw7srPXa2rwHb
Ci7LwnTfMROoDFrTA9sLakaiCeYaM84f9/tPvTJMAEVTra5gUmsHqzgljgkPeQBk
j27qP3kXvUm3hRq3EiOWuAz5xQsNkb/uWLcnY6V3XnzWpmGVNmyqSXTKpmgw8DDO
OfoU7ZclEyQaZlL3Hy4lCfsw15NZxSxPBZBButUGGJrfyBVftjYIMHpzMHkc2NXR
XcGLdrupTFjyVfJF4KDSXtE9w6fK8t1afNPlRDPaEmApgaPVvdazZwORNlbCSGP/
3B9ZLbUQUuDUIupgoXw2WpVJUa42uWvS7s/Y6aEeVCxLpWupoF0G9AXC3ZGe09ru
TANWt5EIj5BEzMdWi9YAEa49lVkl+6sYkZXrE2AcrpTioxVvtJ3bg06gUqPGOuWU
FffrPg5hvs/93D3T4nuvKl0bJEdel2s5f9jN3aeTQwz3BZpFRwW9h0uz9YYsI/IG
9yUIrgti7K0r3fHJA9EYoGAiaq3Gye5HIafsGsoJ2yp9CLliMAfrf4Ljc5NzutsA
j6q/hdmwNvex+TKAhQ9UizJTLaXqOh01FArGebzwrYDKkiUKXBGOmtVdJvdu0ulx
AFMEFToyOlqyYWv15SYCEQ10XWZgiwyl/7ITyHA6BxdA+O3EhmKuGgFmiGmGF1i5
2YGMLvNzhsFWHIzcfd6JK82csKNy/7Xal/LfKjLZ/ieyv0+w6k++k+17t97Xotf/
2dC1e9GepIKsUkEeGBP9jlFGOOtqafH6UHdAhTSOCrk6bDY5GSXJDrpRU42pQJ6j
Pt2Z+tVVjh8REWSD0VWlPqEv0VoXQUGK/bG1W3JD6X/6FQjyJKdTTP9PPSTLq1Jh
PG892mnPhz0PEKvRP/emKYitAXR8fOMpVH+3PpjnE0VScyY7sbqNBBP75hxxliBy
fv7a2iPDaZlBU3n40ZBNxEOCl/xDcviI2uh5y1QHS3ogydPF7tOfe5Qvb9elnEao
6WNZhyWhebTrNLfFEYmgIK9OvxrflHbm5s9i1rdTH7yA8QKToL7mFGOjBLZX9Yd1
47by1gnkhk/s9cyveimr4XaPzAw4pnGx1mQNdP97jADAp1n3Twp+TXeldtw2JFGN
12pd4hZa36ETsJbUNrvZ6DaFQrsQkGp3z0Evn4pHyeWk0ZCF50GdUWaIPqRex4gA
lkNfwO/vK1OMPVQBXXluKhJ1A5ac09F8O+p3pI0D/6LIa/3gUufJnAcj6yoFxUd2
y+8KkHGf3QoafHznxJr3UvH07JDb+nGtgBPnSYwH/QRWEi1+Ge8x0ZJxJJO47Wo7
aXIcYwTyjmpUpEHQ2p8pKdYAzkITkd66Acb5vAGCx57X1LGK8XZKxbLeXHevOagP
FF61DyWnrq2ih0tdO8yjTXBqLp9AYsqzMIrU+5tyA2H0cBO357r589L782ZMneuj
mv896HUGa58f7rQmklTEObz63c7vfrCOa9wMrzwDVPbEb+ladFn+KiWpT9q8Lo/T
WhEEN/CQiopf3ekkfkmVEeisOms3VVyfhsD8Chqw91Lsytulfy4k+c3t007RCejO
cNcpCqbIETjHGZq4XQhwqme9QkJZlsLhxe0nyvN9ayqq7btI16MT5C08VSmmKcKm
b01Z/oN2jmUN4A9UzSOFaPCXptBXN2NP5qKvzCBGNQjEf0jxDGJM/M9g8o/3PJxw
lJ+IHwfTHUHDGam24zw7wqActnJGIRfr/8EhcRJNSlOhRXHouMMb701tmjEpK3uM
ERGf2vc728rTkPBHQpHaBujZswEiOAEq1/or2J++Wrejh0ktVFj01d7q41RaRs5u
YjhtWqOUucJCgZCX044lvRf90LY0w+liOE6Q/czuApN4tJmgM/bv2KFaWA1RpeCi
5Cqt8lY5m+M413bZ/esVO8GC3axxQmC73yjLV4CRciWDpuwfRmyU5WtN4fxA7MOh
s/HmXwdKrOiqD6Omd79ImqoQuGHCj704L4xrWcroXxSRJJg5T5nPScb7uCpcaqze
Uj2+yhZTZsWfyIRuVHYBrA7Q/IZCgYgj4V/JUX9GL2E9ScSJfLc83ydAlpmS1+lx
Y1DPPuutjgH0zGLFNY7gtzdm9vO6BB0VmbKP0Za8tjpTdiy57eqxJXlEhk7MyejR
/QRTiuyScQ99Icg4meuJfaIs4iDIuDWxlI8gGPbemze719BK0bWCkSrbyDNf+YKV
O1tdf179h7PmLKekU1aXBiX7NFf0bgcKCzvrY+4/ARrBZdKQsLaUUAPy+H+I5u+O
kpqsOJtyNGIi9qtjXjFBZllTeqAV6wvLkMOcXD1lxKBJpzNJtqQEMGRHaVaqSJva
9+s3lVMRFSUZf6Mwjcs3z450LkH4tcEPYMH9pb3LUJb2p0huCmuuqao5+WjmZoOc
+pWFoTALjwyVxrk639Y+C7e5OLBimwCvcA9BsWX0kHop2bxVIKEGZt89Vh7i5IHv
mAYxJvwbPy7lY0LpAJ8tkl9W9eyTRaTDZAzW7sumL2dMuXdaTNgPw7A7eWnocBhH
tT+VeVpffBrviyCgPpLK7hFgJFeIR94x4zP9oHwmYwHxiP42L5GYJHEKr4/v3Udy
yxhtRJv0tidXK41B/gBWJ8Kk1//WOqOXrMqxhC1yb2i1/sCpCc3U5LUBpzikR9sf
DNID9mZNGqLiD7WmTGmbmShCmHmHrNhVRSh+UvJ/FuYXhgYGpxGibHRUTNWRikLK
UXx6RsnCXxGk+btB+mtAY1zd59peMrX4qJR4LV0uYhZplkMGoLVP16qgPfPSMP8W
5/ywE5/jCC1VbQhqywQUGR6KL9EINuof9KKtTrbCOr32uKrmnTtSsKPKmat7vNCl
JL4qWcegaM+PBbuAd8kIEhiTxf34PiFLMBi/PCGNAmokDjxG+cDpzxD6cqmwkfuq
Kx/17PN+QDA5MoMS6akvEVQBaUoqKUgNgeFTFdWkGRfLjwv/2boAdxBRWnuA356Y
u7eXwHP9D1cAioFc/mO9jixfpD/WTaxmEEMbE/G2UcKBO2w8RQEnIzwXPjJ6wr28
toodoGll8UU5wCXa7S0xXgWiEU7ONoVwsC9nXpUGmjG+PuSsfc7axNtD3w6wNS9U
4CskcFkpUrrmyjKG+aAnvi4DUJNHAIenaNwsr/vmzES3kLKSqrdPAtLg4VTfJ5k7
/Nmf4cLPYksSfleIl6oC9GyaYYcyCSEaKIPZ3dsjfAXll/Lp+L+NuCYhRRLQpu02
ovjiGdN1ULaJjWPzVjvMdSjg+Coh1fceyHwzQEcQXkuKfT2CIzZ2YMmE84eheDKi
PrBwiEboSHCUUjXjZHqpCNkxBZpCqvCVnUdSomkYmQHWOGKkVRKH0gmyvK7T9rWm
Ho9La35dLb/ih3CW2F8eTaE7hVVZDYqeZk93OeIKKW5+pwIm0HQ2nbqeb587U/pk
dPi6NGUiWUzuAvEAAE7xZq2PMdpXXL8UH+JZ67Y1q4z5l5jUi4Ndwitd1Du/UCeb
f8eM0nFGawm8fARKEHqSIpkiq/5CWEyBZqHqycuCfRVtHtXUYFDkbQru2QvdNqbq
xBkib3Oip7csCr0G6IfLebCglBzlZW7Aha8bvCJ4cD9v+zHljdepTAfcZfygudjg
1DodryM4AlAI7dXMvDQoVSP1YXNjpUvTeT5B9cpLkZ7Ws78XWBt1zjMEqY972es8
1qBwwGrMfTR7SlcJVHs5TokMHUMKK33eJtsn9uO309yNyqy/hWN11Hr8cnOvDifo
gWz73maQTp+NjluGG9pg1tTzbdi0N1pazWaSZoiyNGwfvfOXv8MUeMp6MlvHaAmv
UETDGE1QPjclSrVu8mKE0fGYDT+cwF+fX9TjhNBPLWX9f/3Zc8hEdu8ASD1GgieP
/vf/BtyqHQlZw4fI+/AFxvybGhsy55KOpWfreIan1dOJ+xsa/PpGW9DEUrZccDU4
NN1lC5qs/fbFzn+cbpanShb2PyKvijyb8slSsdY040CTRKZsEGT+JLzXwXRtW8bN
dz+a6pxRpdzJizqcjHtE7VHUOFibFvvBS3ew+H51N3GZALXCx+zJk7Rt7/WAucEb
NU6c8r1Z57jf/bHRrWnc2X23EAmcaZy5QscmHAAwRKF1qyDTvnukgqJdQj3HQZve
72NoHbVFZCvMnlJ7jxLCuw8hJ3KYhpBNHYoWhgdsmYYULlMtswVANbl0Q878P7vD
5I/UodyMPxtFNMREGj2br20nY7sS70nF+GP2tVxWeiHYtAtzWrRAHWMn0oabvQSY
/wU6aLe6gr8n/PjFcOgHL6ZGOJ0ZrsGpck7MLCtfv+PBqDpyw80M0f/7M9pRd7og
mjzo6zJ0gbDqiQz4KZa86h0aEHtvCz2l3N+rVtUdfZ/iwtvU9nKHe7TqJLF9/JIk
Ww36Yw8VqiSLn+hy0j6cnLnnnGcZzR0G/tt1zN3BTSsbhTnQHfTrR8h9FgISaKzM
fdJx63GdAKMYnVQ7Suc1s/Xc1awMq7LCNYgwjGnyzJX88KS/UK/rlm/sKAbOOOg+
iTPxp2H7T/hfs26yDlABvhHJ7eih49sLRMZI7Ml7KktrpTCdLgwVjK8YpmenFMbU
Ir+gZd1VwwEAXRHCVhjQ1/hVUfJgNor1qzEXMLha7kMWU/dDFauscwZN/evs/vWy
BqDAdNp7Gyd0UN57rt6WhwZSifCXZJgeDdqR+C4DmZKdceE8fff28LO8Q0GiBzCX
E5uBCF3C01dm7lvSZNfcBhnDSP73x1AXb43mhwq71lKrpI4fgblFoBafNRcV05AM
t/wS++1ySewTf5H4ZTZWeJculk6BDYJNgwL2AmUi9MNwXOgbjBkKoePNMfOkEKNb
uBG6JM3xQjnjCSebBELQQp9w+AyyuISmx7QlnjVPNJ10JiJQxtbehpvecHXaR/hT
4wrQeHwNfQOLWLs9uij7+9J+R3fPqOUgqe7F6/NnlpAVIemiFObp5Q+SHgs2T3Fu
3PWIHwTxSjuYrV1reQeN2TxBiaVq1s28eNuAGZN4lTvP+M4ZVREzdg5wwvWUJnVU
/v0EhotW3kyiptadIj6tqJ6ltScFOWyaUCX/933jLnlnYR++/hlYPDq4fVvOCfmc
m3l1JEdtMu0ECnQ3AFzOm28HlPVtCgPp8pxVgOakwDrK7BDswLHVWbi+pFE3V9Vh
jU+YCJnZPD30rq+oVBrmek3lC33i6o5ocFuQ5Fvr7REAunMd5X6NpfCvincbjfsU
TQrqUKDLODQ3EoHTP/3IR1mION+RnEntuqSTih51qaxfnsYHGQYsc6+qNWacWXc8
O5MvKWEd5m0bOTwUIbgJsZlMdr/2RsF7TTXgB9ktcq5DFD9nTpHqAD/sUDEtyzM4
fVYHkNOAxmXHxmxgVUMPEdOYWMKd5ZSkdzmtFiQ4RMCE2kkm4aWWK/Nh6jAQ0E2b
TuY8FXrIgxe7FDLnQMXjvdngu8NwIRzJ29zcXI3aicA=
`pragma protect end_protected


`ifdef SVT_VMM_TECHNOLOGY
  typedef vmm_channel_typed#(svt_axi_slave_transaction) svt_axi_slave_transaction_channel;
  typedef vmm_channel_typed#(svt_axi_slave_transaction) svt_axi_slave_input_port_type;
  `vmm_atomic_gen(svt_axi_slave_transaction, "VMM (Atomic) Generator for svt_axi_slave_transaction data objects")
  `vmm_scenario_gen(svt_axi_slave_transaction, "VMM (Scenario) Generator for svt_axi_slave_transaction data objects")
`endif 


`endif // GUARD_SVT_AXI_SLAVE_TRANSACTION_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
XE7RYfbmfSUClOj/Gsza3jeMpmlgNk2nPJCWi/RZkK7vTBzT5TiU4sgeUUtyO0ro
qdEW6tMLW9NIRmtaxHQYyLxfopGzOSgmyprbF2HCS65kplguGbMWY63555TgQ6CA
5kIsi/OrlrfyqZuqdOk+6dtYEU6/c7HFSN5fbIq/Cxc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 64382     )
JAbGRtntQWmMGyQxRwUxjPWuiVea5Bjenq/NHnYuWw1vvtI6r9Bt5a20Q1zeYTG7
jPMal0DrvUxoqIUCkN1KmYZnmkB8edCfcrda3eTAPSgY9rBvC4Po9l6FERZztnGw
`pragma protect end_protected
