
`ifndef GUARD_SVT_AXI_SLAVE_AGENT_CMD_SV
`define GUARD_SVT_AXI_SLAVE_AGENT_CMD_SV


/** @cond PRIVATE */

/**
 * Special command assistant handle container used for objects returned by
 * the NOTIFY_CB_PRE_RESPONSE_REQUEST_PORT_PUT callback.  These objects are
 * first provided by the monitor, but they are then transfered to the driver
 * so that the response object can be handled by the driver.
 */
class svt_slave_cmd_assistant_driver_handle_cont extends svt_cmd_assistant_handle_cont;

  /** Handle to the driver data object */
  int driver_data_handle;

`protected
.e=CL)0Re31CDJ&)Xb7Y5Q#b<V;3VDHg)=/FYD1^+.91CQ93CEbG6)G:T0BIRa&@
c?M.KB@R.,J\69,e?aKVBV^R@#DFE[=.BP(&X,=JV184LJZ(\\D[--/N]K3S6f=?
;]TN8(C8<.g.aH?IJ#JN.X\a<V+)/IJ9d:JHXWQ]dOf0<fBJS-ZNYMWd/2L+Lg_f
F8-OaHV\2ad#K6/YUcF_/N.S8ZMO5WNMV[2bN.#EM_7cUP&@+>L&4ScBUbJZXg(^
Y7W?ZQIVRVM8CfOEC+-^UKa9f+&]F1N=g#([c4c1W8/)\\HUS>AOYYc#6&eQ/)81
N9F]D<3X=Cg_B6C,CT8W+1cf)^<A;O_J6cfHE;7+5=fROTd,&>E>-A.?d3AG&F49
I)P_9H[A2WT^&S3/7.1A0UfJNE/_b:6QB8>T8(IG]d[OUa)^V&U#OJ+OaT<Z5-H#
7bI5D:gV86cWJ\#Og&-),?KX>L\+AR+)RKf3<C16Sb+0<0<0+8UI5cdK<F\E0eN_
BdA##]N+1N0PLQ=C^@dC?)UXU(CGH>.8(fS<f5d.6/7(O+ggbHX6&GEHOP=:X:K<
Z>6LT<cS1L3(/W9O/3QI)aH\P?bQOUe;OUa0>59Pba9TZ>+RN3fBegJ/)<8a6)Kf
Q)APL7fLQ434]P-+=f&JVA&JQETZ,\358Dg,5P4fb]Y8FI/3.LKRN95g9BU<2AQN
b9]-?62U)L;@BJDbX.Y<B_\dEQ^ZD_JcJ^RJQgONW8G0\W7)6/JbL5OaHagUVHeL
cM[Jf(K=,Xd_bTPcVO/0A_aL83R@Nf+3P:D=Y988A95W6,5=;#fG4_92[e6a17V3
EL:aNPRTS0b&d8A(\8VKWI5;3+YGX_a:0))^#;U&]#c2PDP5c^L37DD5SF1AK,#M
L,^1)Y69W>g/SHXfbPEcDE9\H>AfggR996X0.dYEV>6;7?:MF^#0-;2[/bgP_P<f
>DX^6I,Cg?f//$
`endprotected
  

`ifdef SVT_UVM_TECHNOLOGY
  function void do_copy(uvm_object rhs);
`elsif SVT_OVM_TECHNOLOGY
  function void do_copy(ovm_object rhs);
`endif
    svt_slave_cmd_assistant_driver_handle_cont rhs_;

    super.do_copy(rhs);

    $cast(rhs_,rhs);
    rhs_.driver_data_handle = driver_data_handle;
  endfunction

endclass: svt_slave_cmd_assistant_driver_handle_cont

// =============================================================================
/**
 * <h1>AXI Slave Agent Component with Command Interface Support</h1>
 * <hr width="75%" align="left">
 * <h2>General Description</h2>
 * <p>
 * This class implements an extension of the AXI Slave Agent component that implements
 * the Command Interface support methods, as declared in the <b>svt_agent</b> class.
 * Apart from the constructor (the <b><i>new()</i></b> method), each of the methods
 * implemented in this extension will be <i>export</i>ed as command accessible tasks.
 * These tasks will be declared in the shell file that implements the AXI Slave Agent's
 * <i>module</i> definition (which is instantiated in the command testbench).
 * </p>
 * <p>
 * In addition to the methods described below, the following methods are
 * available in the model, as command accessible tasks:
 * </p>
 */
class svt_axi_slave_agent_cmd extends svt_axi_slave_agent;

  // ---------------------------------------------------------------------------
  // TYPE DEFINITIONS FOR THIS ENVIRONMENT
  // ---------------------------------------------------------------------------

  // ****************************************************************************
  // Public Data Properties
  svt_axi_slave_vlog_cmd_sequence     vlog_cmd_seq;
  bit                                  is_cmd_cfg_applied = 1;
  // ****************************************************************************

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * Indicates the last verbosity setting requested by the user via the
   * log_set_verbosity method. Used to enforce this verbosity on the subenv
   * if the subenv is reconfigured. A value of -1 indicates that this method
   * has not been called, and that the verbosity should therefore not be forced.
   */
  local int last_verbosity = -1;

  /** 
   * Status flag to indicate VLOG CMD user to provide default slave response
   * debug information. 
   */
  bit default_slave_response = 1;
  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  `uvm_component_utils(svt_axi_slave_agent_cmd)
`elsif SVT_OVM_TECHNOLOGY
  `ovm_component_utils(svt_axi_slave_agent_cmd)
`endif


  //----------------------------------------------------------------------------
  /**
   * The Constructor simply calls the parent class' constructor.
   * Note that the parent class' name and inst parameters are
   * not included in the parameter list, as they aren't really known
   * at the time of model construction. These values must be set at
   * runtime via set_data_prop commands. 
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new (string name, uvm_component parent);
`elsif SVT_OVM_TECHNOLOGY
  extern function new (string name, ovm_component parent);
`endif
  
  // ---------------------------------------------------------------------------
  /**
   * Run phase used here to raise an objection for hdl testcase, it will be dropped
   * in hdl testcase.
   * 
   * @param phase instance of uvm_phase, which is utlized by the base class and 
   * helps in phasing.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs overrides the driver implementation with the VLOG CMD extension.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   * Connects the #driver and #sequencer TLM ports if configured as a UVM_ACTIVE
   * component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  //----------------------------------------------------------------------------
  /**
   * Updates the subenv configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for the agents.
   * This extended method insures that if the user has used log_set_verbosity
   * to force a specific verbosity that the this new verbosity is enforced
   * after the reconfiguration. This is only applicable if the agent has
   * not been started. 
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ****************************************************************************
  // Command Interface Methods Implemented in this class.
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * Command Support:
   * Instructs the component to create a new data object of one of the types
   * that it supports, and store that object in a command owned reference object
   * so the command code can get/set applicable properties of that data object.
   *
   * @param is_valid Functions as a <i>return</i> value ('0' only if the
   * <b>data_class</b> argument does not specify a supported data object type).
   * 
   * @param handle Functions as a <i>return</i> value that <i>points to</i>
   * the command owned data object.
   * 
   * @param data_class Specifies the type (class name) of the new data object
   * to be created by the transactor (must be a <i>supported</i> type.
   */
  extern virtual task new_data(output bit is_valid, output int handle, input string data_class);

  //----------------------------------------------------------------------------
  /**
   * Command Support:
   * Instructs the component that the command code is done modifying the data object
   * (config or transaction data), and that it may now be checked and utilized.
   * The result of a call to this method depends heavily on what procedures are
   * active.
   *
   * @param is_valid Functions as a <i>return</i> value ('0' if the <b>handle</b>
   * argument does not point to a command owned data object that is currently active).
   * 
   * @param handle Identifies the command owned data object that is ready for use.
   * 
   * @param delete_handle Indicates whether the handle should be deleted.
   */
  extern virtual task apply_data(output bit is_valid, input int handle, bit delete_handle = 1);

  //----------------------------------------------------------------------------
  /**
   * Command Support:
   * When called from the command, does not return until the specified notification
   * event occurs within the model.
   *
   * @param is_valid Functions as a <i>return</i> value ('0' if the
   * <b>notify_name</b> argument does not specify a notification that is
   * available for the command to use).
   * 
   * @param notify_name The name of an <i>vmm_notify</i> notification event
   * configured in the transactor, and intended to be command accessible. The
   * name should be of the form "EVENT_...".
   */
  extern virtual task notify_wait_for(output bit is_valid, input string notify_name);

  //----------------------------------------------------------------------------
  /**
   * Command Support: 
   * Retrieves the value (into the <b>prop_val</b> <i>var</i> argument) of a
   * specified public property, in the command owned data object pointed to by the
   * <b>handle</b> argument.
   *
   * <b>Note:</b> If the <i>prop_name</i> represents a sub-object, this task
   * stores a reference to that sub-object as an command owned data object, and assigns
   * the <b>prop_val</b> argument with an int that is a <i>handle</i> to that
   * sub-object. It is the user's responsibility to manage references to such
   * sub-objects.
   *
   * @param is_valid Functions as a <i>return</i> value ('0' if the <b>handle</b>
   * argument does not point to a command owned data object that is currently active,
   * or if the property specified by the <b>prop_name</b> argument does
   * not exist in that object, or if the property is an array but the
   * index specified by the <b>array_ix</b> argument is out of bounds).
   * 
   * @param handle Identifies the command owned data object whose property is to be
   * accessed.
   * 
   * @param prop_name Identifies the property name whose value is to be retrieved.
   * 
   * @param prop_val Functions as the <i>return</i> value (the value of the specified
   * property). <b>Note:</b> Regardless of its actual type in the data object, the
   * property value is converted to a 1Kb bit-vector. This return value must be
   * dealt with in a manner applicable to the actual property type by the command code.
   * For instance, the command code must understand the int equivalents of enumerated
   * type values in the data object.
   * 
   * @param array_ix Specifies the array element to be accessed if the property is
   * an array. This argument is <i>required</i>, but is ignored if the property is
   * not an array. If this argument is out of the array bounds in the object, an
   * error is reported.
   */
  extern virtual task get_data_prop(output bit is_valid, input int handle, string prop_name, output bit [1023:0] prop_val, input int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Command Support: 
   * Assigns the value given in the <b>prop_val</b> <i>var</i> argument, to a
   * specified public property in the command owned data object pointed to by the
   * <b>handle</b> argument.
   *
   * @param is_valid Functions as a <i>return</i> value ('0' if the <b>handle</b>
   * argument does not point to an command owned data object that is currently active,
   * or if the property specified by the <b>prop_name</b> argument does
   * not exist in that object, or if the property is an array but the
   * index specified by the <b>array_ix</b> argument is out of bounds).
   * 
   * @param handle Identifies the command owned data object whose property is to be
   * accessed.
   * 
   * @param prop_name Identifies the property name whose value is to be set.
   * 
   * @param prop_val The value to assign to the specified property.
   * <b>Note:</b> Regardless of its actual type in the data object, the
   * property value is sent as a 1Kb bit-vector. This return value must be
   * specified by the command code, based on an understanding of the data object
   * property's type. For instance, the command code should supply a string for this
   * argument if the property is of type <i>string</i>. Similarly, the command should
   * supply the int equivalent of the applicable enumerated value if the
   * property type is an enum.
   * 
   * @param array_ix Specifies the array element to be accessed if the property is
   * an array. This argument is <i>required</i>, but is ignored if the property is
   * not an array. If this argument is out of the array bounds in the object, an
   * error is reported.
   */
  extern virtual task set_data_prop(output bit is_valid, input int handle, string prop_name, bit [1023:0] prop_val, int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Command Support:
   * When called from the command, does not return until the specified
   * <i>Command Callback</i> event occurs within the model. This happens when a specified
   * command accessible callback point has been reached. At that time, the model copies
   * the data object of interest (at that callback point) to a command owned data object,
   * and assigns the <b>handle</b> <i>ref</i> argument with a pointer to that command
   * owned object. The command code may then access the properties of that object using
   * the handle. <b>Note:</b> The Command code must complete all accesses to the object,
   * and then call in zero simulation time either the 
   * <b><i>cmd_callback_proceed()</i></b> method or this method again, otherwise the model 
   * will report a <b><i>fatal error</i></b>!  If this method is called instead of
   * <b><i>cmd_callback_proceed()</i></b>, it will instruct the model to proceed 
   * with processing after the specified callback point (potentially using the data 
   * object modified by the Command code), and then return when the specified
   * <i>Command Callback</i> event occurs within the model again.
   *
   * @param is_valid Functions as a <i>return</i> value ('0' if the
   * <b>cb_event_name</b> argument does not specify a command callback event
   * that is available for the command to use).
   * 
   * @param handle Functions as a <i>return</i> value that <i>points to</i> 
   * the command owned data object for the specified callback. Additionaly,
   * the input value may identify a handle that was returned by a previous call 
   * to cmd_callback_wait_for for which to automatically issue a call to
   * cmd_callback_proceed before blocking until the specified event occurs within the
   * model.
   * 
   * @param cb_event_name The name of an <i>uvm_event</i> event configured in the
   * component, and intended to be command accessible. The name should be of the
   * form "EVENT_CB_...".
   */
  extern virtual task cmd_callback_wait_for(output bit is_valid, inout int handle, input string cb_event_name);

  //----------------------------------------------------------------------------
  /**
   * Command Support: 
   * When called from the command, instructs the model to proceed with processing
   * after the specified callback point (potentially using the data object modified
   * by the command code).
   *
   * @param is_valid Functions as a <i>return</i> value ('0' if the
   * <b>cb_event_name</b> argument does not specify a command callback event
   * marking a callback at which the model is currently halted, pending this method).
   * @param handle Identifies the handle that was in use by the command for this
   * callback, so the transactor can now get rid of the corresponding command owned
   * data object.
   * @param cb_event_name The name of an <i>uvm_event</i> event configured in the
   * component, and intended to be command accessible. The name should be of the form
   * "EVENT_CB_...".
   */
  extern virtual task cmd_callback_proceed(output bit is_valid, input int handle, string cb_event_name);

  //----------------------------------------------------------------------------
  /**
   * Command Support: 
   * Start any sub-components
   */
  extern virtual task start_agent();

  //----------------------------------------------------------------------------
  /**
   * Command Support: 
   * Stop any sub-components
   */
  extern virtual task stop_agent();

  // ---------------------------------------------------------------------------
endclass
/** @endcond */

// -----------------------------------------------------------------------------
`protected
GVPDQ+0D9T/:GBbB97)D+?Y>M\E<T-L\.@U5R_M6?8(NSV#9YH.R6)SHHZcI5699
^#,3<>Yf5?=OY4=USLgT,EaNCY1YS]MO5AXH@=:9QJ;WKeEe53)H>#MXNDgTb;<B
^8.(f;+;JVbP@8Gb0GUO&#;d62I6Qb?#F+.\Q4>/77AD1Yd=G^MaF;Nf1<6PJ;@3
WbTgH#1R;XZc:+OVJ7].J,E-TcK,;ZD;4]K-gP_60OEK7YS/)FWJEWZMM56b_5VO
47C8>6V;8-GL/.cNIHY\9\/\dU><V)>P=[X5-4(GCMK-&^gY[Z,#,8A)P?KE^:ff
Sg\\X:Hb5+FS=1M<4<N?0B_d8b9Yf[#e,00Z=G2>PP/+>TeP9LTZ00BfG9N)Y4BN
[\D[4J[FP(Y1JGHLO_^<QMBTd1_W]DTRA6c9I(@R4;EaE9QZ,S04B/G&2;U?J)f?
=OUOB,_(Y\.H^(9FDa@82e22O]N,g(((UWTc0BBTfScFC3VW2;;G1GD:fdD&_VD_
>3LKSF8<7S8EZE@/ECe@1?81,<<[f<EQRSVF>ea5SJ=76F#Ec?\Yg_8Bdg.+fa85
G9@40^#^@cK3#A83#(93NJPUY-)1BC_TT;WF]I5RfX&d#\);84)@=]2abYT,9MKe
@LVBCbVAA)(-M?+D\OW/LQ_6/06W)KGFCY]\#_\9GMJ@:6ZG4b^#;?_YGH]_4,C+
XBYWR/^EIHX8B#BeV0PW9g6=X&@59E9.ce.KL-UgKNRNe;=:,QJ6bQE;THH5fCD5
.0XDI3Y8DY:3ScXOG)fKG-,J720=P]#Q>0X#aM;8X90.7a13WRgacY=YC@#[I<Ga
)U3AL88PRH:9SQYTNN83Q(IL)f#;]DL9.ZD(;^b&XRX495&0K@[LPFPD[ae853/(
ZSN3M<?0G<BL[]G.6+4Af>:<?3)/LEFS]=_-Z,(dXVfJc;.b+[f,HDF=<@TJF9<@
/dUA=d.0F8F<9/SBUZD&CaQUe+2S@B(afF8Y/-3BP#>>Zd7^P6;N975Na3.E/2c6
),M?5>>38IbM<M4^.Sf19,I>f.-;;6GX>-K^;g#8NHA+]daS<A<RJ>(WMJROVNX;
^(T?(]DD9QACZ3_<_(QP)FZST.EZ_CO=D+I1/,?g2?(TV784(O0eQ&3^>6FI91W<
_HW?DXe>+#]6&KWR;7]^:/,PBE^]<T^+A_BY7S-?dP)S@YWOW\(((LdB;[GHH-7?
eDeXg4GfLWW7Lg&0#W047U)]<BHY05H:Sf5@eU5bX51+dadEI&^d;J)S((143E97Q$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
dc^7&^K0A,;gD_?M1.NeL)I;L0OM&Vf7E6W1\UeB4gRGaJY,)5ZH6(#H-Ke/6GfO
E_cEGbd4L(A-81]HKb8MUJTEc8X-;QXA#Z2ZAg#AW2]:ZFJ1J-f#F(OR^J(JDSd#
5=KI>.;PH&4e?c-8MMITUQ<5<=4HIgg4f1EUa4J?E276)ag1XG)TEP0DWBTI)=Ke
TO=5.7CN>O+73;7J)R/_Q(aL:>X.H2\TUbbSfN6I+V^KNK^]]EeVcK+VcIcR2)PG
MEeO4dZ(RHCBA)9-WM]YAT):ZV3T?V)9[eGG400eDZZ2_dE?^-4+(G42@GHA.bIB
&TESV[<Z+E2]VP9cc:U7c=_eAgJ>^BM>2OHAZGG3],P3N9>1&Y4dbbXUeLKE)G6R
X</+cV7_a/\Ug[_\QDNV1_?<>F940#LW3g-V2:>MZ0g]3.HZ;+V2aYW]3<-RQH1_
1SR5@59)g931D\SNSZdNK.X745cRM;S64>SG^65J0^.^4CN=>?6_48M9)E)G0GcH
fEW:QW@NDXK&/Z4O]@H+V;CKITY9-]#fL.caYU]=SF>+RUa_/<0/_^6/;?g?c#,Z
=/R)K(1G9MW==U=<W?1.0R-8U@S@0CVA.;CCB#LMQI?X1C=_T/:gQ=>ET+^>H6U7
16C9M8S_9(]cP23M<G=.FdV>KDR9N,MP(6cH7MWO&=C,M/f_0_<1H<K-XZ7-K=A+
g^g/PHJS#cBQWMLRXg[\<<OX3+?X8JFQ]dOM51QS1Ogd)2Y+BUM,DDXF]LK6A#58
DaVZ74[H6+T>^09Eb;V_WaPB8f,YY;<3-f?4aaW2]07=42Og@+7^dI>2I-#R.f\E
[[B3@BQ9+SW6>DULK[H6c7^NgF)5QA+R9@30e&]FSaU?8O4:,GB[MF40AdOH,Q;,
\@eUB<GIOF\-=7G\R6<J.5cBRMb?;TSK<c-TaKZaN/,GOfWJTJ+7CJY768M5^/7S
GF:DYdK<RLKDN2>NK(Bf(XCOF[d.@H//c?BHT#0L.V0V(6KTVUC=#O5Q#A=_7:[I
(SVC9a<55]9-4d9X@^5P3W,EbeOcC;aHd8.[?&G0QV:SaU2S#1DG^#\JL;O75L)5
JN0UL@A=GQ-\)FH[[AXTC@9G6&YEL/+VG)QM4E5:K@,.T]]Gg;(,H6^U2\QZD>@\
&WX1^9>NB?d8eT>YVX>O:NBC8b<GY@PKaJ-+<8]X;ZD:N_ZaHDN8;fBWS5S7W,1,
e],Q88&c[RGT)+WHY9eYH[BV\B_+=cBQJM)1T+(aW(?CaE4H?=?(LI@=V7H&L#dK
#KW-:8]O1[(EY+HQ/#4e8aW:7>_/4#]\CF9DK^=c7eUQSa]WLX;RgbVR[MQ4@_gf
bL(2fN[KSL[?#gLN+&+;a1eG?.2B?QU^0&/O6_U2SeYePe&==7SV#2SHO65XVK>1
bN9&g=4(([]e>PG7KAbQ/3d9?07-UTQ]S?FS-C]>BK\]a,5WMfX7N5;C[.U:@7.c
RQ+VKeZ:J):MQ#J):9CN^ID@T(MZ/KfD64[K&&0NdT-_.)^-8M]GbD6GGd=]^=D/
MKaIM3K<4[ZXf3H^dRJ&#UTF8-1YYDddXc]>)Z;Q()dH=QUUa5\acOa_e84IYXM3
@[P4cB(c0QU?eKbegX&IV3BW63-b/16NZ.]#ZN6bFBOXG_ED1+DX>3C83=;O=A2^
c;N5S=&\,+G0eP87H;GOC6N\2SKegf.U1TR?1M7;3HEFcVA-@9HcJLKY\1U<[dP7
f)dOCK.],3[;E[=G]>_F(MeGGEgAf1/a4Ye8,4Y3BU7J(@-32#A/-Q)6MJ,FX1)[
AF6b&L-(8TIE;\M_6eZA2B9X#ODSZ3[aR0+EJ]GfUcN@Tf)ESKQ)V(6aebLSWJ^:
C7E5bWJNA+K/YNXI>/DZI@.Rd?@-.Fa<:])7H7.cD1?c&CV.F9+;GFNCV32<20;6
65UQ-4C2(K8GXY0^P,[J<:Q(N;F,O9PQCa9YL^M[Q1W-K(&[BY&fC_AN0PSY9>-9
K>[XR<G;]B9DGZb[+QES.MT<<T;gTNN3#6aQUV0+;,?NA+Ja01^VGO_>+L]Y@;Mg
Q^X.OTdM)U+.3XJS&VK1M&9ZYMS[7<ZPc-1U#MaTPW3KedVa0T5@(-dHeH<=5ePg
ZSGEUBD<aQI355aSJD5@&8:EOQO37:/ea+U9E-[1^2XZP]2PK/FSN],<6eC,TV^<
d;,:;T[)6-73_a\gJ/_H+Q>:-9gJ.<A@7E3(:?JTc-JTC/DA/+C[])_C(bR\85?&
L8,L@?E:Xf9D+Z][\O:798,Q6@89g?F]<[Wb.C.KG5\&67&^2I,ME2fUa3_AG,+5
198ZSS0#KZL=bgGKI:_0_^;R[DF,<F4-2;,@RdfH<L#N]&ZJQ;60=#MP8B]8^7(D
b8X1>6TSA-8M\KRL_YJ-7U@H14aB-4<()7R,FLQ\;7-)aQFcK@\8-K6;XP1QO#3G
1,O9e9d/]8(76\?HE1d25>/@eQU(XQ7Bbg@P)?U34Y0\)?g?d(&[CB1fOTQ(d7M;
&S+2&0^_\X-5>M+0<B94LE6c8@Y=-X.-:@7JQ(D411IU/AHc/aIRc]#J]eOAUabg
;3(E]?agX:fga9_^gM\HG:>f=1(9@I=94B_,#5(1JR)(X)GB/,[&TTKNTIfQ1XeD
bSR:F[0M(>T6Wg/:KH]]J8J0RW2eDgL7^4.2_/97cJa-(IAGPMe[ca:4+@DLSJSa
V(Kf=;9IWCNd:EcSe@=;cdH&bGU/B5[35]\HcGO5>+\c[8>^+F8KcdbaaNdAV;#N
]+>T=&OX,&8SPM79-8N17=[NRJ>]^Y,L3R:7:RB@/SM9U]PD58F\74Sa792_XG[J
74Rd(+,dG+b4Rc;V:];W&/@@66[FF8B0/QOb0Q)OP@\=&S,&DP6@45_BOQS0?8ML
HbXH8/d(?:=5K#;aUO;G(1JRVU26U0#bA9?b=gS;[INZ^Eb]#3e/H3&E2>+TFXH2
HT;cg+WcX#)67>)[NT^IMgVM^R=_gHT0,]6^,=OGI()[HG]AQY0RFN23]7?M,GOO
<J^9D\Y0/48Y1<UL(8IHJEPWAK/\c),\0.=aYAP0A=^\(FM8U#N=B?A>[E>SK,H[
AS(V714_RgF,[Q8&d#CFH(Q\-GO-MJ5.,M,BCbC5#LYDEg7A#,E/eYgL4;((Og.d
a)X28F>?IfFDf&\>7_>5A()UFR[O&Ud>?8:EBY\S0:K]OgSEBG?J^R^c;#f=;f/7
T?WVE@ef:C+=EF4LFC(2Zg)7DT8MIRGdBeX2H6McDL\eHM2bQc-:,E96/W2FaGeY
_&MSXf=69EHfKD\J0#6&82[OKOPOB:>H^.M<<GKNVe@Fg+S&_@aNV7FU5B#fEX8P
b^,7&+DU.bY8,W?1>,<U<;dB;D?^NS0DZ4KE9a-D[G<E5Z3VA_[_0g_WaT-T+CdW
HMdH6-B>gC_Q-<]>R0d7>J&E:de^PWe[::(@I9K-D)6V)QfGV/O(P6>ICU-(VFaB
/-J27;&bU:/&O&7;b+3ZJUY^VA7V(<:dS20=[E1)LKd212e(9K6\2Wc7&8N,:LD)
#(3<MZ&J.+SQD0@Z,3UESf<-5#?V>#a;M-e=W9c1F]A,A6F(3GG089A:8.+-d^C:
MX>-FE9CK^VZJMRWPWH4Ta@#>@2.;4M7;H^OV)DF_PW7,5GXR=RNR,C\dY#,8GW7
S,JS]9&K<.-OA7.D(GM7/<JbFL0O(:OXI/_U[8RMNFG(^XJEV]7G&M5D&]90E&@P
JgF]RYH9,<fYP42WI7Y+1Qf(8?IB#@:1A&4T-?9,a0>a=GeSNLF[VPRD3O?Z8fZT
_(RD+E3#[HNU8NeI\d4Q[0HQ<LZT,:WS.7^=O)J#PX0K-@IF#DPLF]DV:0C-d<)6
];<)(_F\WJ?2O3(BK4&NMDJ0P3aH;.-=D^XWI6fc&bC(a(7^cUC(-:(ZY?N5@K_G
CV;dFV-1d_^?-KQ.#^W[22JXaePA]1<3]b[aSPHO<Rg:KbKJ])R44E3XT3:cGL6=
F8[Z/+HBU\,c;2g[bCJ(O6MO<592a/2J\-<PEN.-MNU^ZKD[\Bd8:?X\\9f:@,V:
T?KJ=CF]/f/HIcV(IdU5W<91]98.RMVX1<<025&d^I[<TB=fL)M&cfF7?^+RE/#.
@)[O+cF#2T2Z7FF6U[f=NQBB6TOTMLOGEGV,C&NXXK0fI/9W36@/:b<gQKAeH5.9
dR\a?cMKW&aR3<+bXd-D(cNF9BJ;-dI<H]]H8@?_B0V5K+8X8g.XcJB87K9eYR_R
@<IO/(,bc_dE3fXc[)7b61Vg()P=BFP;8@W<8TE,6>R1+D?-X>6T2I&8P?8X.M@@
A#.\GRH)d@XU1ZNMW6^^;S@Q01YXB?62@)/:.<)Nde+@.e>2Y=M1#26VBTIL_Z0@
?L2?U-)8F=56.X.ZAZ+dECKO<a27IP3dX,E7OK>gLTQ^&:=K8JKG,3R<I>OIZ+,[
9F5SHJN7G2aW12cXZe7c2HC-\c.U590_H1(f,2+b[6MFPB)-b^PLL(2MT)e@:abH
ZDO\.4)Yb]XEL[e8WGBG[;&QeB#(S[fbA]5&E^b+f-Mg3+J&.UW)6c,?^DR_[ea4
7f9V#T5:_))8c9eG[19Wf3,378&dXR,462Bc\=KJg@e3D.(46-?U&)O_<(OBg:?V
0?/@/[99@Va.PgY2a0^XV0R747[F@8LWIW<(Udc#[AEWe,R-]?:H-B)DIM/N33/1
27@bUG#I3\FPB]>CVYM45(DYJMLOZSE_B-IUM]1ZEUXffBg0A92;@LOJU)Ncadg6
H),[Z6>)FGL?E36IH75Kb>?.^a94dIXV_44GOQ].d+gNV2.7&,D)fUf.[bH,@,I^
(X3c4CF1_YKL?1gBQ9gRCYVRXRDOe2OEc4V61;]H]J^?QV=/f<=gf<T=KKK;CB(5
8EL&1,Ze2@F=dZITXUZLNX]&-S)4Q>b8=@__&3S+WgU<^Ub,V/EOI;;]+7[Gg2dR
(-D;?/G;2,7OSNKCVagYU,AL:6H+1#<PGK]DNb-SZcKX7VK/7d4DKSYV@B/,f1b;
]2T>O9<O7TOS):TV6+8(4I>1X3<LVOR1G@DBYK>1.-H6?[N_c58O\d9>.<=MfBZ8
?TQbM(dbbH;>9gF275#gVTGf<PQZ:B>93,.UI4[N-/F.e90Ke2-7-7fKL?ZSRE,e
V,b2PRF=fZ3ODHV9L(FI>G&W05-<6ZS+^M^>TGRGZT@9D:^-JV_O(\Y_=[+_ATY5
?.PL2.P_L#+-.=+M91DP]A^.?@TPU_?PSILU,ZBTPR9Y)(BIZLc3@B/HdRL__4g@
cY;5+;PYS[@/W8/.EH1,U1RMD<O/b>e.dS92Za/A?DNbDYMN,Of7<75/>0MbPR(g
db#8&6N(EKM_R\U/YgW>a<Q#G+eG99=FM::gBF1XJ,K[OK_+eK>#\^2.6P#&QFY(
-J16/e=])[ZS<\^)KXV9;F7f-H[bdf6dgWFe7U)IeA+e&6.4,O0K#O7:=,U\YfT4
#Y7Y_g^V04JgQf,?-R&\^00H@^YPS/N5fFg984VC,C)[I.XHTAA_\&3I\/8)+Ef3
^/R_#M?34T4^dC)G\I.R\&^=/MY]FP;gQ/<NLU2=?G8gL^W8_]EW/4)KW7)<gG+8
]3&HWf^QP]e4c?68DW-_PKZ#gPKM)gED7DUYJ?E>G?/bQF^.+4#SVM=,dHA)@a\U
ae\)NW-[7(gE#>U9b?<.14\EZ;e8WfaKfAL6e6;(RLRD+1M^F5&R=YORg1O[I#C0
3cER,ceTE:-\G.UAKgaJS^?f]g/Z/T7]7-QI_=?KKGU9Y_::1(@J2G=d@aO_:JbC
5UaIN)DXY(07&]F/LNF>>MGbD34=[NX5I9P<2+M0GG/)]Q^V3?F;H1^0RJCU&N7_
M/,94ZP^c^B(MZ#5NS-4Y_O8V:/(Q\5_[Q5UcLC5fTaWK)SbfDQNXWa0K@AVK1:-
F63IMMMCKX4FK1&JH^Sa:&2Z;9=Y(^NS)gZCH5.+A:DAS,+\PW4(Hg)-E)BKK;TI
T?1f4WC+W&_Z9FLWfM[5)GH@^T/38F]25?9EX=DeH)6]0FC1<gD+=??)^>)3K6#S
.e@Da#(I,WT_)P1LV4:9E(K_eIGe\gVJ=+\LI,0S4=:JU]Gb7_^AdG:e1GaDaHc?
5b65LTLfYCXHg2IFYP\_@H[AS#fVW<6aL4AB/@_d0CE0?VT6gPGV+FB5X5<J5@H(
H4:J+;9)Y4J<dS0JFE\-gPC7&1Jg5cYI<LUAQ9G[@[8AUc3gR8e&d8MMVIT++Q]T
;dB4PW3UWc+5(@S]0V1cQf;L7][\9G@J,\=(VG407[LTf(EAY-bY-7O;3YCTb&?A
^L/EbZS6T+KP1T52+S]-I8)1U/TMAZVNAYd?B)ODHK)eSYR#C?DXZUU7##=&1;?)
D:HT4R&.a8HcC-4?9NM;]d<Ra0O/QPCWP2M<&VZ;7H6W6FDdHY@?DER6,K3)_J6,
@C\\.#NOaf9Fc[AE2V22=a:IbVd3A2f+9Bed9KG0.?W0[ac,2Y7M)8fRBWD>F+[4
W2)?KND2563R33OV?,L=#L&4[TVP9D^J42.VARII(cYEZId2BJF(X6E1fEY5(.\U
6bW.A#fa8(Pf\,.-2-U1S/<I22U)5^@V/L(K1XO^5:BMOf/3I04NE<P@,D(NI&#c
b=LSTS7N?D2U,a<F):f=R;UQ=4@S^051=WGBIM>1,9:KWXXdc+a^>INS(AOgIQ))
,O6LaI5gUIACS_#Cd>(<.(Y@NTgU8=D3.F/6=BVO(Zb=CXUM#-7E_S9;e<73,U4^
N:RRB-H?=MG=N@W8A7LR&9ZK\_SaS3U)1.4^;[E=:W/[;L8\U>CA>((CTJMFEX&c
TB;Y\F?1?HF-U3HZQIbI?9R]=LTDTUEU/6.2Le.Ee#;GFPEfYVbHH4g@0>63:Z@8
Cc;g-89\g>P9W7XYQK8Z#50>;>feQ@&T]Qc.f#1DTd2:24:U#gL#F;7?dD6O]OC@
#+M>2:+][?[K@f=cEOF.Jb,UUA&(/LMI3W60@1QUK8d?>]+/1PS:5_Vg8HWVT>f0
Q]^9U0SK\X(R8^>?O_D;>f(<[QB[Q5Y:W1F4@-=4f+=)c+I+I^=MKAKORLI0=aP3
>IM]O?H[RP9P^bDIg6,:MaDCC64WP?XGKUbB6GHXR](d,J_ST?Lf7(IO&V^XQ5Z6
IYI_&?L3&DN,SH2:R:/Cb1=IYVIe.2=5UD\&^P#XDC+YZUOf)FdH0NW^#ag952?b
XP&2@.7e\1>3BB6?T[=a#FZa36V0(LJF]YYD#f+Y7=W2II2OEIN+[<e+-T_XMJP\
.EO:V)D5],H#DOR+T.d.(88GSXI-L&b-&adY3>2@A2ECc6#>FL5#KERc6#/FS_-_
ZY7fH:f_Y&U^/_ZWGGPE+3^WQa?WgA]U28IK4)<>U55#N=gX&I1^efLgZC=I?\C;
RdDT<=Q7360:G2Eg5^?PD<T:=W?06XJD:ADf(fDVO&d_=Y9fbEW86[1/d1-4WC?<
DSSERC3]1GBTP#\4cAYeb<#;/NK+N]fC/;:CJ\AN2IC7E/D@=Wa&Xg=]K7a8?P;W
YP6#LV/>Ab+?8:FF&TERa-3-V8(Ha9,d6fXE8]<G(0.[\_UT+IZ.e2,[@d)Y(\N6
Z&W>NR4.MGDgR2UY:76Q8EOdXU8:a=3SE&QES18G48/KMI1MV+G1#I/IcI2@e]2:
4_+FI.=dAYMCb<AdA?GP>&Ha5d<?,A>aY9d7(@f_K9b@^7KJ1[aJ<&4\JcP@CWd=
;fU/dJQgg,8c0IRFE1JC55:3e:62+<;7_D9/;eVO<@aN)\:Q8,Ub-^=b-E2(J&OT
RDT;9M.P<dRT0J,_L&6=N](?<^.YHJX&P>EaYN<KAeQ=/RbA?WfMVUJ/bYe>.,a_
eYFJLHR?C:<G8b_EDe9TWfE7c]<RO;)?4#7:DPVU3&B&[MCcR^RFM646=A([U.VH
S]LRSM_K\9@3OaFK(^L16F;8dW4#VJIfA13R,]ed,_f\1RHW]R3+4_e()dNR;f1+
ZZcZ]b^/9D_9?[<T/G<E)+,-AbW]g=0^JTB^K8K#^OG7E/,K8DU&@?=HaFGf5MaJ
GO;+?+]JaePK@W3#,S#SBM@fVcE8F\.4R73feS00ROR=IP1,2I\W.],MY5fB],YN
(N91NB29K_\5L<RL870MYdX\;E>I1E,,&+(VH7?;?49>)O+,1L\>feJ9EML@4Z]4
D.^UaXLg8WSfI:G(T&7E35Z#e]>:HM,G#Q7cY:gQcXH-GP&/+P)-T9DFP]3HXb6Y
.7V5-.NKML.60[Ye7P;]UHTN^.M8g(SbS97ACGS9>QaCM4I@\3T:6&bZ7EUgS6J,
X/,,[CE&]Of>DJB@T39,Z.JR<U9K?\@-X(NQ;1-)E0f.[>Z@.7RG-YSI->J:A1S6
_2+<cC7;^V+cLI3X@]a&_E1)1;T.fC.P+U_+=V9PKT]PQ.H/?/NV<5(BcF]X^APE
Y9.&:)Ma)d1&LLX/UM:WK)bZE2Zf:e5CfOT/5L2K?NFI+BN]gNC4f7GdLZL4:VEK
L1V]fFb6.b09/C85<+A5?/Jd/YQT_1>A:<\b:\-c&)UPYEgT1MN;8;,A&C(],8JZ
g0eUIX0#HbRG809C>9K<T-X22E1Pd7>J#_IgL7@U_@M39>;,RSUe_H+J&b\I?+T+
/]CTB/eLadDNR=12>A+S=O_6)8[H96Ne,5#dd_e(Hae)LB:L;&>3Z88E?BW=/\Bc
c-?E.WDaW]54RK)VHfTTJSPEAHA#2b:Y1BJ^>ecHPG6c0Le=0YW^c[b/UPI.f15N
+O=I.#^AU6K7K8FT#C<aIdAFW84+RGCfO;^;@OQ9Y033_4O,@U@5>e0D0X-LRKAd
<+^Y9];2R<.9.=4J09dEGCYdQWT-cQ,b>6c,PF.Y?FPE/_K<QIYY:+L.-W7&;6GV
H&BJ?;+eXP/&<BZ6:4OGKH7RO,Vd>24&KdA0C.=-)dM4>Z)[eg8;T>=:T/@;,7P=
X2B6>Lb5+Z/TI9I3H^5QcH;K9Hb[9OZNVDXZGC&c_V5XG)GO45g)6&=LHW:^Td;-
5#HA)LHH+QVLMJac<9S_FFI]b2&HC\FVdPVbe7:>(;.H;S55[<G2#.OZSfRQ_U)^
6WW#8(gg8&ag1]gO205=6ZEP#>gL&(:(9aAOTD7_,N4bECVfXd8?6TL\g7b4WeS6
SLQ[1aMW329OcC-fSN;MeWTK#L?^TIg@JT8#14/>H&3OL^KWfBUZ^_3B.S1D=5I\
EaPPG=/CU;5A@O<G0X]>/O8VQ1HOZ->((P3LDAaK^E-F(3I-X.8fL@CbO\AU@H,(
C\<M8g)__TV)^QUE\_.^QgdBT^cH6N5O4.5+E3B?3C1S\K6;/9d/E+G]4E=7BY]O
&aGRR=C<DfSF@d.6U3Ydf,6+W]&_+Z[/BSWdGNQ?_Wg#]3AE&P^@N8<@[R)RD0KO
0)U/cZL].c?RBTTI3+20DYGd934B+G4@<)HJ(LMR\3e]CO^S2g?)RS[\NKEL83/^
=DOF3J05VS.8Q&,;I7b-?7G=:3GHXQ0_?#>L&,YIX;0_+-X5RS1>HMU6:\_fO\BV
ANXSIUJI?4^I8cKX(VZ;UMgdWXMeR6\9-687)?68ZH6K9]H[(UI-:3N#,<37?@04
CL8<[@JG(NcE5K>A(+ND(a8^dZPF/6^7GNCO/=31G3IO@e\3TLW+f@]bPU8XKA(C
[-=ZB/XL=A<gF?QK5eG@b3P0;7H>)<gPb[_<0Z_B3=Q#Z7g]S\+[<?D&cH-f#E1\
,bQUd:+d>EVK-?PR@^@M<:^7ZJQ7HV_gJ3-J9Ef7VU=&)Q1KLW]3&X]?;L;J.d[8
WV9^DGcc\DW5^-0c+IPL-F/)MOV2#XFa,8-d,LZ0HFF+]U2>eC_OO:9^D:0bVFON
L(._E]_e7ebO4>aPX-CSIb@)@-b3B,T]B.9Q:P5DVN_Z^ICQ3P46a0e1,\>-c@Y0
VQa2]C7_1e4Kg?KAD><.e5Z5c:]^bfF<#\(W>;e-[WYH35P95NUJ((537Og0d.g)
08[6)edZd\\>-.>I-_;KQ)b2<e^\SL&-8NSdK+[9[])3,I8QVC,Of@\:/ZCPIPPI
Y6G@)Pd+\NA-6#,EUH3gXMOS-4DSU=;;6g7K(RI^a2D]9;>f[L-6R#_UJ-(;(dM.
SE)?NOBeXREPcOATf^[S]7NJf,RfMG@C9DBagHGXFN9TW+<9V,8[J2:]6_3gC+b@
&?:@W5<#G=9fN+L<(,H;63X<[Cdd:8C7KYP,8>WAIgM1f4;:Q?GG?4>D+U;&XbN7
0;LM;E<^NKJ59PX,P)_Q&_AS0W)XL^:GS&=<RTH]:KTQ53G@([(\bE[2?:a(H2b5
eRM-R1T[;FO>WR7\2f+NNX]HR_0(+NNOF^/8HD:#YX@S5^fE_eZSP6JN7Y9HdZ#L
1>GRP&3^Z2EP[RCL9#:&FIB#=U)^ME&a[P2-gS</2?)8ZZLT@OE)Q9^>>gWI^B[=
aR)BIIdJ+_^^MFTeTDWAEQ0P]e4U=03)13ARa>a=HX4/YbZ13]ROfNdfQLP]MaPF
PR2X(#/d)dXWVS3gKK5P_6e(RRR)BafE5AZSd3_-^UOVT/,?VK)T=@2bWF41JLKe
EMQeA1@^FFZ#2C)KL?/)OD5\^,2eF?;LMfF1gZ;_GLA9RMa^@ID9HM@=-S#+[:)E
IfW1YJA9]QW0A.U<ERH=M.f=4-]YW9+a^fQW;,(GZZ,S,S&AUR^)eBC>JM8Z1P3(
d&2OMcf9O+gFM@NU&P_4fdH@.D8=SV0NZ5+HW5:;34b-SgF5++,bN#3&.14S]8bX
P&7]e8ZDC2<56>c_e=#T(M>XPb6=)^)8T=JcVe>V2dfa?O^0@GZ.0A:UZ3X>ea4)
9U7LbAb[I</,G&BJ?EgPHCb,>\B:XV[fX@D3OK&W;DY=e)==1d(<L@8J]4037_BN
VA5P,IB_>XKU3a09gM;YD.bHAd67V,6/M-Sg0M8e,U_TdHf9^>7[J8>G68IJd,dR
)X](4?GDE^f#H;DUR]dND9U@]^+,NDDN;R2]//e)S[R=;2I-ZTE@NM[SfB)5#HF6
9C(_+W6E7]K5IZZT.]4eb2?Z(-T\fV=+UUFK3[FG+a90&eMA2J8^-\YR&ca+^8:0
L2KXA9-A3Y?V(4_Lb6@TAG+[>bTNB+]g)>^U4J&;N3ZUNG:RX\KSH,/4^,8S&,Wb
0;C)b=E[A)E&@eb[R#BH_A/[^A^79DRXgK1LD)=eYQTNL^cS,gb@H:a?5a-R;Df8
d:W<e([R:&A&MPLW8I/eTIXb2GGdZFK3XQ7aC=^3E0ZdbHg)W8I&I2Jb68AOFMAJ
>N/agG@&JD+3_=-.):^NF6K@PEO62_WYO,f#(]E>e54O[M;W\?\Qa]a?),Z=AgQO
3J\[6ZR6_Q@MJNS9;FQF&>Y;-S<?PDB&#5eJ:LW,LQc91JY9b\Be(N8\-.1<Y]R5
FIE@e.0]V6\H=OC,R4a.g+b^b(30H?,AaRY?I@3ge;Z4OTI@dL7e19@SCP-Q(7\V
2#^/SV<9d-CRME6W.9?JD]L#_Mg?<:G@^MQ1gO2LGDIXF9CS[9b+1cC(QdO9(BSN
D\D)ATJNF2Q[,bO>e6ASKQCV71[f?]M^d39BQNb-Q.gJG^([eJ9IF0,YKUK@S7=(
/DXB:FHDSWeL<.O;402CYD&;/S<]7&&)TcT,JI=9R,,E)a#acMTfE<D?ag_SIUVJ
\D&WF]K^X;UPZ8KGJ?.P6C]&JeBb_988?/(G[1[eg8:;W8G/a;0LD@+AZ]EFXT._
J,\PT_Sd47].5VNU][1EYTLO/c8?P\VE,bO:]8,-=dO8O8#&SRN^9.196#fO\U[A
YKL]H+)ZYc8(FJd/N\g(;I>(YS?_N]Hc>9T]G^97E/^7NA<+.N)DZ>7+I\JR.F9K
SV.+)<X2+D;@6e5F[L=O;M)O&;bTI5]c]03)bY<PRAfe,6(TIg(GT8dU0,MQc412
X0^IX1f\^LVHHc]]&Oe<#L37\V1OPR&IHGMa=MT@Y<1cYbJ6QgZ(9^YO(AH,M?(D
.^_R,DY]V<Fd6BSOEH]V-Q@2\7E&09fd&fB6-+f8-P/B.+X&W81JJ?bIM#/gdIOG
P8S+Tc^^=XQ>8(XTb+8>VJJaH6E[+abGT\J+K8VG^Pf5J.,]D;c))P>JBUg)5TVb
aINT53b?8#J2;EPZRUOGWVNHY4M@F[HdEd,aX4[3#77]448BggM?dCY3[2e-M^+O
[IU[cL<<d/-3O5(^QH>.7IYM1(\4<c]aA<YU]^A^TPS2?\,Z9^IP\VZ):=]PA<L^
L4Jf<4]@GQ43:._[/SSODM8M&AP5/R\JTD[^)9:\<>&C9HR:SU7NDe91&L][2W9]
KIf^R,9Vf,O,EA7EC(QLMDT1X2Wb@=B3f[9VN)=E@:^S[^WEK]@GY;2b5Y84[<)d
-X9NOZIf?IY4[:SCCG]c43A-SUIQ_0(f#:e5Ue/gH?<\VI222E6+K):):d/5dBY/
STd[463/fKcYP\^#?c-/\UULI9(#/AZDB=b;cV&e[8X;3&+W53-C7T9(R:_UK#<3
E<R9X,C5OdAUGeaa&gV+6b>;FdE;D:_YaK]-PK,/CGf9\/B4NdKE=DMK(bG>L839
f6KY_XP.>JO0#eJ038/AFa-gOZcdbA0)=NUO<XSc22V(-5V^A@@+T-KHcdYe/a+_
#I3Ee(JYQ_.#dY6.)^K<==CW:A;>F[]JMX?Q_RK,6J>a-fJ,OaIfV7aEY-):]U70
Ga.923d_=Y6H1SEXPCB8+(9CI&+J(W\[BbDA]9:3c#_,;MQO5=L/EHJUT.S3Zege
8(4Re>PR/Z.c#\K8eMHYdQX9g/PaCI>B#9QOIcK@UMbc_:[G>;<X2UB1;,V.:IK:
U4+-QVVc33Q0(fNd;_XZE,Ra-]IeEe4d534ELUY-B\>]4M#eMa4YQP1>6&3]]_AH
66S7]VdU3:D_B4F527e1<VPa9+/8/Q)1AgBe9\fQ):,HcDNLe?]0Q);EGaKV(<;@
4?c@4:CUNAI)A5=6[:G&DV,<-70b7XPOE)[-?5?-_(S-PG#7P.E<?78UW\RK;^3E
7Pc2Leg5A1NXgTEdJKGRV&MSc9SL.eH([aARBWP7<aEF@+2+D1-;&;\#;cE@^#=/
&(/cNEQLGWV;DM]d7A5,fZ:MK+DQPH&]6WK(H7S9M^,T3\2547f0[&fT,->B<JX&
NXcaKV]+1D7O96L&GeE;fe=URIF2_--bB,)U[d7Z6Ue0ISYE):\8=MS@PKO/<-<H
F.O3G;UL&9WS_g&B;8PQ&(aJGdZA.A?#LB&[W0^)HOVE-/CfX7N6/@a)R3aMOBD7
[^^dZM;8fFO7(,CN=-_C>XP;BgZ#P_\;3D_PYO19TA:V,Le51c)&VY&YO-4]2NUW
6c4]R[Ke;0ABP6eB,dXg[#2Of0g6/HMCSW>#G<@g1f?(R9/Y8Bc[,8LcZ&;,e5TG
_B:_>W:7>D(H09=@0,=e=G?4[NE<_A?:V@JR1A>D0124<E([b[#O&TFON<B2T5eC
]1)1eHE0/_X[fa/T15I?a+4(6-CJ5&B-bG76:3D((9/cA#BA9GBI^]9;#1MBB][]
^1Z_fRE4=33-A/;b0=;eLN4D]X3(<7eT4&CcgB8/C;5Eg<3TY;/#HJ@^-4T7042#
D0]VKgg/T0((2XC?H(FJb5B/-5Lb2JEX7b11U.=(<E9JM:R449aRY\B[:EU=gC>2
2TODY-OaFb)YV=W+K+8Sg^#7)IYIRJ+3DYN(<\RLA6O<[X5.9+cK_T]_.<KL8#N-
:5eAEg+NcH(5e9GR_/4K5g[c^@&X0O4Je1E^c9#gW7_Z,4Za:9,S1;9.X5:cf3=P
MW&:F^a45aCVWCXZP0cE7ZeaUM2gNf]@2T1)TVg2YRN1D@CG&#U:4)NH^KQ@+5:S
WCNS0a7dLG>.cAT[S(0S97BCISd>^Ceg&>#>)Z.Z\=YT>WZDaDgcW98([YEM8](&
+L()_L7Ig)-..2X^dZ3V;71X+RT)=2:<=/@30?HX=U.2<\>TY)\0&f_?c))R]_AU
cKN+_\=7Eg,G?8dU;W#b+X&=W)(Efa2Z)U?=7c::JH(L?FF7a?ZL3];cV?a397_=
&(;TW8UU\gG75A/HaNH@SR4eQ7L0g0_=ca8S?&I;:gA)AfUaW>=7B.UK3R]:I:]_
\b:_UA#NTbG;9g(J+@D@;F.@+Jd)UY<(HIC.+-&Q7+H&bO861aV\Q#+A.CTcL:cK
[XBU(#&XL:A((b0ML.IeB,NVR?@-Z@=S\ReYbA>[4>3^?<KKPGM^71^[D_Z4JC=_
W,>RU90KVL41UV=RV)PSV<LZA@UXIUKI@W_7Ab_cd4>NY=@Y]F1J3H+U2d]]^9J/
0K<;<\J>F;8&>1HdX;Q\Z<_JW7<eId)H]VVcdP]SFC84=@AWg=4b-UZ:V9NRZ@0c
&J-M47LO4;1Hf76F#)_:OAW5E=+9aO(;;Q,a>b1[?[Z1=<N-c2fB&W_(EEH+\Z)a
V1M_1/L>+>WOR8,ILN2fV+C6K=[-DFNb4E1d.5>W18>CFG=/8SLOG+;b\,H</LRT
Va9bV7OA<F0g1-M#(LO)9O(10=MGPRc@P[_>F6,=RO&6ePTI1B98C>gV_J[ZeP5V
6/DPO@._]+#07S@Pe-]&-UE4H=FRRaECJVe<[aeRB(P>7e[PQD[]B<N1UT5a:Ye+
7>=(&KgC9;V#fSb^g8_JM_G-0-/0_)(ZeVAM<-e+._J,QL/0<Be4+5S<ZN\7LBKA
#8<PW57eR=NACRd96A1(&>EVg.DC6H35-(--)OQ4&/DV\X7a-3GBec13P0RUZ0Uf
[(&dJ>(c22QG@.9RSBVK&aS1=.3X(;SA-,:A9Z/\\N+5P0Ee^8OW=>)MJ#@PG;;V
8dBSWWAT8[NbNYc+GUN3NDDQH?HV&H]=<TU.+9+b68B7d7EOP-&be4(JV;&fG>Q_
4J<Rb(-(LNO3/>I5[5L)/TT8-D.6E9K7_I^42K0O@S?1(5>LPMD_3GU\Q&7A6TM/
D5B<WGN1GDX)g/c-KMOJNOQ&=[0QNC(\[6/2bJf3<87KV]a6[gXPAgg<\U9g>(5T
Pa.V;<74dTSM-:@+7V\g0#V43\e#a:fa4C=TeDK5cQb+50A^-FIK>9S#@a6K)=YF
YBAIF.0<TC/:FF(CRROL:[B2NP9C98XVS\[=4\E\490=YXY[;Q#)Ofa#UbUJ;P00
DHgX(@1#@:1/:6@V,(I,(P<AIEY9]=14EL2.Og7-8WL,_He&e;>B@DeQ:ddZ]<Td
-]>7I]E9^\-A8ZU<^A.\0#M\D+KN3M47I>CBd&(Z8#gbGU(/??3.@fYY.LeE1@aM
0CX+[CI[8?5M6T331V\]HPeLa0P,C>XG]/=//<D+0FUgPA+/[9&P=NCB20K,eR;_
Z>QcQHZ:<&01.IC4Q01T@eNB]CEU]#a2,76cZ6W/-KF3WIf#bSJ3]b6be5F-6]])
438d7\&_0<HJ-g[5?KKVgDX1HeR:+>07@D3L@6)IZ&Xgadg,Zg\aCW3Q0PUR1.U4
[NR)L[8I4Y^FEUPY-:5JEf1]T8HY_DFQ02C[AJL1_EOVUa6aW6[L@,cfU[^^75X:
d3&7JDRC0B660WS5)VZ26P<?+Vf/N=e8Ef?0f51VP6dB,.XG+O[0aOPJ,4A[Z9bB
d&e)PB_@:cBNSB.fD^XORGM21OG1=,6FgI.gCKFD(^gJ_G<<M<Z7)K[WOdG9bY)X
48=(WJdP@7/801HHQ:Q[WGIe1e1gGLPC/2QA-V)\1>LA8X=Vd]d<2;9/c[;7UM[-
MFR[J@D#D>#<3GIIcccd^6e9TOZ<0>_DOUd2=1_ZA>abFYUEC35MR55dI-W258UW
5[2_KZB\?LOZ+9(IfC#8/M[#P;_[UZ<9b658aWBeVD5H[NVH+TY)@(Q:cg#Z6]+L
(H:gf./AW/Nc.,W\>[:_&:T>6)):(Zg0MYJ[V/dPETZf#<6G(:J&F>CU.DZS;)J;
JPX@/&RX9Z4JbTA.(gV[f#7PL<.&(UL8fWG(6eIO:,D84F>;A>6[>=f>A4^(V8fc
D:P_V856^F#fG,aM8K/D/@4FfQIO:[?[9:X2<_S@VF,A3EBTSge#W.e>4<>;<+R,
a]&+?7DBQU;KD_PCPET/05A]AYTY_B?7XDQTWdOSb]BRB[aF?E_2ZW&R]PDAG+:@
A9HGcW+WPZ7EY^2fcO8J:3F+JH@6K8LEWBT2:]I9DcO6GC.+O.[.4)93T6Q2\bd?
ggb^_F(_)O-c3?J<;HO9LD)#_gCU1A[<fA(?Q#U/9DD9K[g0#U.C&Z\2;Q(aG^N7
US:,7e_Q?RdNJJ0S\^M^,)9^RJ7PM=UOb<_I]I3ePNgP1ZT;W)9CCV1JTA;/1OV0
R7P7]_\9C@Hf58QS?X=JWCe515)+eeeQL?:TBGO_J_4SQQ@A9AMOZS7GV=<LPgW1
,(,]b)/9;BL-1,@?F959b;CP.VKO/<Z<[&R)JDT5+U9?5[-TH@V:5.<aO@R51,U#
]fC+)=B[aBcBd<_ccbC:-,a?V)aaccEB1_^06M,dSTBQ)LV4Dga@&7A=A9K]H,0a
,\S]Tg>f)0CDTYa2WcR^A&8GILPB_g11JDE^2f>TeL;W\#SJEf_d,GNPSN2C3D20
>#N.JYb+G06b]c;/b+WYI6P1PSf-a.cVP+L.dFC&RH:SQ)Ia)/-U5.9_@4fRO(1V
KJLLM7851(g1;9Pd]/dWFUeOA(;S3g&2a2-dTfDT62#+EV:N?]LZE7=eZ[IQ:bdc
F;2C5QG5f\gL2Y^L7Gg[XYFZS^KI;Se5+?<X#-CO9T)E?)<ZL0Y:M4->W,45fJ=J
#J3.XE.PGXPd_YY\OU05NXaKEE61UH.H\LEY38c^]LaOP@P;B4FJ5KK&gXE_096c
V-POK#M=]@Z3W9e8D@5Q>[8C_g^6&5)\90bZ>[/c.Y&efBgJT68SALb/P-_/XW0P
MSAg1&_FG0OXCQCS-ZU0eEEIDKIACX)G9f1&^KW_8Hc\XK.9,73Hc0##9&BC.9J8
\413:(0R_Z[gN/F\K9:6&/SSg#V5WHI;]UE=UCUTH)[P=+=1M0Zga@MG<)3aVeDX
LM-RF.(fLEGF1b?4W3\b+-G,.F8N0CV?[WX;<:A[V(g;;#1W.4C?\PFKL?4WK[BH
F36f:QO9_>QbAd5830XJR5-NQS#&FD6U/TB:.K25[fBFR-<P3=U,_WCDa2+X[cNd
0[-]KA[Rg-cMP<G>R_RYS\?;2T[RQP@3O@8R8Z>N-\RASg8@:b3<G\XW9&?TX=;1
F_,(A<_R#Z.f[>&]T<R[#HWbN3IfJ6SCN,c8D\94PYI1^gd&Q,(S-eP)[S=f_1;]
>Q_Mf(,Y[?(gV(Ba.-:=)<P0:J8C&#;BJbOf/MH[&2KTc56V9>>Hf=EZY#b2[1B>
513YF60TQ[6)A[Y(UHfe4;?\QY2TS78HUR<K?HDD)[HA]MfIecGT^C6F_8GW,[I>
;5Y?]a[^]g((K(NXT/cC@P)a?b7,99E.g/Rb1BY&LV3ba<E4R0Ub4(_WT#D[<T@=
d98L3D/#Ud;S?ABV+:Zc-/3X699=IC0>?8fX\CTcGN,+^P8cWTbfX&cSbYI8>WXK
,Q[Yf0.4SG?>gP@D9.3NRAI6>2QMC=\=?S9KfL5dUX)BZ&>?gWH+b8),We:4G-C&
c[]dIYSWG)CQ[_Lb_B8XeIE6<OU6I\>Z\.M=7[//:X.[Mb>P]5Z_TQ:)Y-AW>XF&
6+D-Ne=M,:S>9,(B?dZ\[K.gSNF8Y=^R2@Q@B(#EAU2[b(=H>G\dE[c>;N\=eLXY
D<T+\<eI[OA<V/@bXd?7J.dY&BKZ93W;8c-UD0-KNCg,PX8cGC6FfWg@\G_\9dgb
^,<?1B.2,-a#.2(],&Xf<YV7_1LB80--_c,KBVU8e2-<7[M2GDT\DbVTQQcK\Y13
C21?JJcLg:f-4;5)]5QOYcbOP/,J&Df92J3@@V:JW?3Q_N-R1ORMA&+YARKI\TMd
LeVV#F+10TLYg+Se@0#XCEBXOU[B#Fb4\D]5TdD8MP</[WaRdd[D3UPOUCJRbG+@
/@=]9F14]A81]@MZY7@4)>dS]DL3R[]IE=-OMR3-@&PVN8?^6J[e@K;KaZWT-F@6
@EA+83[W4RJB+Yf.(D.)]NY+bOO\MY&\Y^OX)@SR+60#/3-P3YHaFE<=fb)@?X#&
ZTR-1YW&N^2J82&VB(^Z;@Q3VC8ZbSD.L4X.8F@YN(_D(+ceJbgSFM2JQR-B2JUD
CbMD4\dWFHbX:c(J2PS9OAT/DHb4G^#87&4>:4?<CEcHJQKHTA._[Ha?05@T-\/a
@.^;4[&2]<4OX8J\<C5IaX8Ra^e=:@@MFcPKZ@:X_4G6c7.O[(HP,IfIS&2M4fgK
Y0:&OE8FC#e03;?3#OL>cAU0XOfH/5OK@gA4eICT(H:Zd[TKbH69,WI[35L4MPOG
5eQKX:Oa3dO2.C])(TASd9;8O/MJD)_^9F2-13;Lf:HVf]4EA3>89<ADBbg<+C\=
J>8I)X9#M><dIEJ9-]H11;I^VgYAGV@6Z/WL7-Bc^N6-EZ6&Y1YD;V8OCSf0?F/D
7dZ6\SP21eX/dI#@\(I92g<LS+C=;B_FE603]?)(:#\Fe8fB#I<8OS(4)4PE\5CI
bQ-@)>]2058<ddC^V+]SdHfDGSb9dUH62;.VS;])#7XJX,UY1[^]PgQQVKK2FeV>
W;;U<;4P9(50K-a,e+RX19-G#cfB((<:E=9BWAWIAb4@&Ng)OE<7H>Q;OHV+TbW=
_UUf8XOdW@G=_D&]6VO4Cb/T<R:6#e7U3a@W6f&6E(;1[KBVBSCB/#&f4?VCRMe=
XA,gO9RW7CfPQGAH:AYY&OJgeC<aa<J[?aCEV05Ac]91DX1caKg>Ad5E,^J;O.#M
&23YHdFZLdW83X>/HbJc4QT5]ICJ1FcSe,d=9QW&#_T7BR(\A9D;S_P.,F-05CZ2
e#;c9GfQE2.+,7[=,UHfL79#fMUT,A[S]]1Q3BU1=_I.5:(7-YM5g+)D25Q;/R)2
XP/edMGIZ9Nf,+Y.R\aG3]S0[(1/0_?;ZMCZbT_V9cGJ=b<e6)<^bUO;I463@[33
DLPJ\F+,V<-4:PLU(LQUe(0H-1,=(51G0F2dJ_Vf#\:G;0089<XKT?&dYC2@Dd@(
BZ[Xc2P]R#>A##82J7P<L::GKDeNSTWI<XWJXX]<[@](:^7Y9F<,Jf@46_)1?BM(
]3(1=+1HM8YS>J8DVB:;d.S2>-X#7CA1FA8PJ9X/TTD[(Gg)(<JdF-PA0U(UG@E2
WdNAH/YC@_,7MCeV8S2&VCEH]<KN(d96)\?/YMS9c:<aO8:Xg<7a^EO9^-S?Z_<O
4(Y-+K=UM-_H4?W@3aae#4Ea06DcgV([/<X,>I]gGN>ZR;8.HX(-BeaCg.<gGg2F
b8[S,-A3V^L)e@5]gHWQHODM1UN4aQI6AX^d7g.@?;5#GZ=eU,]e>S>7]U3d3<5_
WU0Dd6P3])7Y;]6O\H,Y]WR<?N8c:IA8BDdO))=45_/9AN8B(8F0gX2Td;#_Q-6<
@Z:TDW1998fZ4&g#@WYV9X]X-,\AHaQ<2-HbLWMgD[YOQMUgGD[R5&MJ@@LP_\5R
7R9ac1BAA2Qe>&Z:XG)Q/,HUc78(O+fB9LWT]A7-PT(Qe81\0gJ^W7.4OK]9;#\[
[5dL,Z\#B39]V(01S6_FKECKMU@eR6V<0Rgf889>C_IFU[3#EVM-1VW0(d^V<,V(
IIeLNd+)^87VG]UML[A>Td8/B0N86dKa6S=LPCQNDK4e23aH.P>?J4\Rg@HfK/HM
[M=ZQ84_OEZaMI=WQFSb.]ES&CbC/SZG/-@ZCC+#\^7YEHC(S6Re@D..AJ\=F.1c
W[bG.?a+c,[SN;;9/UTF+g3@YTR[b<Fb.DJNHdBa<_L?X(]=G[1^:Y0fK:2WZGI,
3L<aN)-dO@Z;GbB;55#BZGGD\&[8c.;aT,EgI:CB8X2,96VBde=_dHN)7X+.e(C.
6>QbBdUG6DfL&6-2De27gM@dLb?fL84I1/=B[>@fOM8;>.@MY,__:96gYCE]_cSG
HLYadbK7#<DGcdeS@f9C_6Gd(K1O)1EPgB_ZSK5&Z7XW\@&>4K8(;5d&C1O4L=]T
PZBe/]/@&_b1DQXWR((^[-@1LP&ZI#W#;e\<7AE,G/FKJ.H^1TA)B=8E205IG&5N
^C+&Zb8@[JE@Db[Z.-V02&+-+1OR5\N7;;GCRc#H3[J]_YbD@SRcC\7N4,_QfHYG
g[Qd8))8W8#e3_J3Y^3&\Y77]D,W3GJLCY)40MN<=J4GCV[TVQ9R^e@_[<:(N<JL
#>5]X+==&2a?94H.>N)/FY+C+T9f:V?efe4306KH[\#/A+:&NVYU(R[.QWE-.S@#
ba:4NbeGfH9V7Z:FM:^RP3>T@\3(:dS=+CdFVT8Yb.>\<.8@CX&J<cDAQaa6^5Qg
OV9A6-N\&;e#8DE93b\HJ?:#^Z[S8J:YaFM3<f.Ob>dcb<JFCUfVH0)\WO5e8e0&
G@SIMO7AV]KL&VC\3[]\C@BX<TD390\\35CI>,UIN4L50[_NOe(T:fb/Ja;-PF71
1WWa(]50GbA<U+W6(aZeSVR9FbGDWM9PF_7^-@600V>ASICI^W0XAd^eaU<5@Ae@
K:-X_&:B8dAYcH3f7&O#-RL6F>IYJABM\36THHaOc);#3=AfV:eD+fe1X-DKT@=K
NIYNaZeH/]TAQcQ)T^J5f+RF>#<4P6A,GPJ1R;cM=XCDHM&5-_@SY/c--_6.<QCH
]XVQQ,B9F:RcVS@CK)VMg7B8b-CYI;dR_VD;]M=-:\VgZf9K2eA7Z[=Z^#CD,V1+
MOKD1dM9<E&4+1EKTVN4IBe^>@C]DQ[HW5OcWRYA_<L1U;PR,I8c];)MYO2<e./6
\eVa_[_N15<;3+AKO1dMNe+_)VXNP.I46(>>?3+6^9>J#f2PY82V#\g@5^I:E)]O
O>^]Rg],=U0BJ&KdC9&CV;9;Ge53ED[6/2eKedH@0UAgCM<8FXP7OL<]7T?#NKM?
e6XbZXVe]b)<dYWZ:aZ\FSQC]X#/Y;2&W-;.U_T/&e^2ID72^X0aOHgH5W[92V>e
10-WE\ONLLAOV5?#2PbZDC9bQ)dYP[a=18K>0BU-VXV@3W[(A,a1ET8_MJH9E04S
f484B9C,TJ@+5,:S&NH@L-C:ZQL#J?F:0.(--S>#D<9+<_QP^P6eP(H#-O+PBU#f
O(._0RRE1ab+))PVV6?<LIWN#IA0dBVX86H<CWS?Jb3JO.Zc84cTD4[.3FVECWFG
3^d2,U+4dX??C(E&+F0T-&dR7#3:,eGL:4X8[;MS,A_+:<2=Ra071V5N?Y)4#@QE
VJEb89+B#KYH][3_Ed0/,J+fU(1gW7M_2LHXX^U3f#85SQK#/+D=B+C\e0)_J;4E
<><2.O+(R=;XGZ@=0V8HB(X(G&73VK[Vc(H=;0J+D4/B,U^E5+:P-;2dW[IZS9@G
S[\Q3Ed@/2GCFQ7FgdNWg>\U-4B43=4Pe>5F_Rg]2J9YbN^:;08PJ3/X_W<PgUJA
0TF[W3.2&W+:#50Se7,#?8/K>^aAL#_R;aWJ4(L7Y+[VdB[-Eg<36XFJ#gTHNg)9
YKAG&0#UG.ECG=V];G#4@UFda)F8X8?ca_5QHYEJ&LR_E;@[\GC/;6e>&IM_,NgZ
-=<e8O>)@M6K_&4>J_6X8ZNDgJXK;=f8ZOgF(CcDKEd^P=K+FMG_:R-\b1.e/JDa
XR8PDWa+=6EYL#fTcVGB#d?K]cF6@4<EVNPI#B1DeH8)_ZN+U5<5Qa8@YOX3\LO=
>.Sc88SUYT/OVdP7S(SW<D>V.76:C#+F<@c?J6QaW_bdJE#(TY_0;:=;7S3JgFX]
XReA7<HPgdV77@T]4aJL_2cSd#:a2]8cJLQAD==V0Ob:a,I/@f-[XZUYMIF<1bH;
E5_8)0g\bbMc825/QNbILY=J[.OgZB=&&#B056K.<3>MJ^Ggc8&IgEWdC4Q.Z/4H
V<_?[EU=EBR)7P/OgN)GBf8E,T5GVG>7-)<,/CLZ3[QRC]_>NeU@W8cF;3fRKLVJ
>ZT[L9?g&.X\^&-6?@N_V,bM1U++^YTU7CAX1L3GeEAXR+YG=36P),83@gY7:3MB
QCCb+ZSW\9a[Ib([46&;cJLW)R+YO.>#&&YgF>78aP.#c32GFSO3P1T\LC+T_;fT
61g7f3,M3J&C?&L^.ZNRHZW&IE;DT<628_Y<aPL::Rc=f^d?C2)]7HC8W,1>N.\<
7(;&Z(RbW=cIf(8YE40LFDdF.7./)0Rg[2ID\,2[#AKaX^U0S=/2c)04X5/.VVR#
-A;f35bQX]2DZU+C5G+O[Zg^g^NVDT2FC3]90X)+?@)ZV^>?@EZN0e5XAV#GgEE^
cLeUL[\@[TF;c.5@Md8KLAT5H91<5/@DHfX\Z(_?9a,&?I4@3a[B28=0\0@#</3d
&@U1VF:3XK4(3(4;;9\b2a,&3GZ:3YW0S1&Ae8UYB,Sed0E2T#WY2F/UedO3e<.)
/\5_]UG;a=3e-7+/C.eMO.VQVK1EZ1Gb8a(9C8^M@9:F\J7<JDCEU4T#=EG6a=4>
E@=@HA3c.5=ARaP#+[P=;.c3ac)0AeB)-?N:K).\b2L>&9Kgg-3:8=VNC2^:_:?d
O4GD+48@KgPL>(,]W7F#Y5NZZUGAZc_,RbK71;d_35J.=@.b_2YNFOB0LEb^0:d&
KT1_=2QX0).a3N3[IJ-T7fgLb].]\1_UVT97a)U.^bQ3EQ6.WK>TS9?1BLZ4[NV<
dUCK\G1840HQN2bO+?RJ?Lg>IT2#.J73,_9-4&>-Db\#<<=BU\JDSICSJC[&1G(R
V:2[c^;ce=9aI+ff6Rg1#UfH.<SIfe.I9-#=M?WUO6Z>_37WJH<@bM:Z\^EWXZB<
=B#;AZ-KYBa-QO3JB;3g]PYA)XU2[;1T2S?O2FMab9>:#FXe?T4&\?+Bb]@/-cPB
>/g@4,8NF_.U;2.[VOe^9I0Xc.J^P<,H3C,2M)V9LI+FG>1[+aS>57W-,:Ic0?[?
(]:J8F+T7aTTIZZVCgKLFEHP<Q9-H7,9;7&3OM,1>4GL^7_GQM?F#+N;aP19FdX7
0++ME1:bR+]d,OHE.fJ(UO+IWg<^/S\6/UE2)INWEJN(G[gR9RZ9f[-+617)?@aO
aUV>,&CAH>J]<b#>++dV@fMC@[95b@&W8H5<UKdY4#WTf_.]7ee8Dd/:8P+1R^C&
Xa>RT]R,I@Q-aId-3dI1,Z8:N_\5&.:cRTIPd-c>:5;=a\eUKDS,INJc;]77/XBA
RL1YF.)+D1,d?_,a]B>becHH:dLc&HF9Vc<:]3W@[AfCB66067?9>G3\A?<OEJMQ
0J^B8K^WVRYEI?2+I;SM]97;Y/e8gT-c)3E0f5B3MI6P_7_#G)6SJ=4^DK4WNNGP
=N2R&D>Z4=5:V+6GB44O2M?Z]X7;OXd?92.T=Y#Y\0]fALeaC3(NF)J#7eWR@)P1
B.?I5Q?]=<fDDQS/_&J_2JG=;&Z]f^bIbF:^M4:3?9,1K1Z6++]54P8I\)c24E4<
+7ba9A?741UW?9TI1E,:CBBdS_]Q6JSD](M/4.>0c2-d1<\:b,)-I2OWSB3CEDNM
&.J+]XQJ1bDD/JQWMW+aWDJETRZKY+^+6E&Y+I3IJ8C@J?MA@deFd@9YSRf9#?U4
Ba6>C?RAY&K_2=<KN\LLU1WI?f8O](D.WdNB/><b\T[7HW=0JScHP#cc(-9d:3W7
JGdA@@;]7gOMV6<e9<[RcKPcUVDKcO=OW1Q1:/Z9ME-RcFXX<D_9/_6I&9<Kd>#E
D>8,()WaYGDgEP,F7+3#BcL9@@5S5d4IW:U-B.3^OIGB\&1b1@[)5XS+CRE?Cc<)
G@;-08#=>,\,<X64,C[R6_&VMG/;-DOT?\3WO3M8QQ\5J&MI_N6&<BP-P1c_][);
-PR5N#E:GYE+T/KOC/b5#JVKK?c?/ZD#OLM1[77A6S>E6GQS.dd:-9c0LSEU5>1T
OWQPd)c;,;LcP:(T7\aA,Zg7L?DP[=a_4BD:TAOc[?^J0D<I/9Z6#3U6,fQ#_U:+
09>(#Q35/,[]5):KOA.1aG+U>GJX?@HKM1Sa,fSVRY^VB[IVI]#JN^5QdS)7:)T_
?1D_/>OaX10NbEg(6_.0f..V,FK4KC<_]@O@6].JZJ&K30M0WY?K-Qd:HdR9(44/
bUIAX/e(;R_20P5<c4WdSb^+]Od&=Z9,R]+,QPVWZT:b.A2M]6RP)79?)g&W\<89
[X0WVf&_;\6E8#(=40cc#b=FW0E72XOCcTWfZG(1W_O8V7cIA8_2f=NXSK=&WbB1
4DUIaLB8/8c)]LbVRZHKGgY)3:)AYQ+Z5#Y4X0(\cfQ[27J4527ZJ_I.Yb4UCYU<
_8dJ[K8K:XdfB(S@P?B7/NHJGc@=PW2L<W(b>.5f+;O(AO0Xc&L-gfH=E)O&(?W+
_H9fKFNa@/.]H?]A44]-;b>)H@T(/eUd^9MACY^fYdV7:A0TP_L.O#3gYXUZM/\L
O^Y5K9M=fd0]XP1c9HgB4H)3R9Ba[5G5_U60T[#AK50M^\I2]R<^V@\=@b)7a42d
+D4MI@3b,CP<M[+\gIBEU8L\YH1[IS37(e#^C&,fE&a6P3I1g\FZW4FOQ:_?+g:a
#EMeCBPF4GW(A8Pb60P<8;.<Ya8(59^b&.OL>gDdY4IC/]XBbA#d+RdT+BU_449H
Z&Qe;P___U9>:-V&FegJWAQ<RU7>g=-;D[2DKOCG67197\afd:[015eGSG2GgA^H
N=b[\V4^/73OXO1-5;0aQ]PSDT^YaCc0R^gWV^&/G1dW6]MK/M#aW<Na#[O/79O/
Oa6JTCEEAbYCP8OXTEY,T]8:\A9X=6;56-Bd,SM[a2OEHOd>&5:SSJ0Y0>6W7;W1
^,34[EX9>dNL:9AE(c@K]WC([JR,,MZF6Nf5QTB8M#BA=1I,[1P5+V:fB[.<(J2e
S74_JH-f5=H-MUI0&-c_]N^0MF]<T>G6U4&_Z\&M(RP(?bLX:c873HM7@A<.BaIE
\>,cKGE4R?.<?>Z4SA)I&S-+,T&?7-VAQJO:fHeP\8.M5/:#S&CW&M5-QO1(BOg.
J,?E7T^bRHQ)07@Yg6JgS=],SK&EBU+_/FJ3A\;BQ]1-DTY6X\-9W#CZH?Z)aPSJ
P&[fA3dQ@&+<]Y,1BZ]#V#?0E.LEI]WW@)=9#M?.IcR;<8DU==Qgc9?=FKXL_^HD
,5Vb=dY6La(5Z&b3<FU_>KH\?-dE4]94;#BB/T&66UI\G19E5c4N5Fe+cR^PJHR\
.GC_81F?6U;N(;=-2XA[?UFa&P\5?8:Z^7M63(/V[)5Y+PH^+g44Y+?aR:gc#].C
S3#aVc1(<O?f4Y>d]R:[GPR)GP&MU0C;CT:b;cWHLgJ]\f=+9W2Db?)4^YWaaWGK
JEH_3OaG@+67S)cDJR1^[X2NZE5A;6X&-Y<LeR^7gS8U;ac^7\=2b+aV]51:URL3
PD,+NWEQc:TSC_OZ+6=C+&-D.K&,-@dBVQba7KD8A032f)4IfP:[TD5aQJ\^d,S,
T\38.KFP[aX^GKOM:c3M,I_L2N8JIF^O_3Cg2&G2-L@\+VQS;^,M@+>TK[VNLbSD
(S+;X^)E@O+;WYBeaUaT#eF6\8+G]abY;g0\F^K9N,UcH7b7QFKFL)C.N6^0Df#:
58aB+<YL>46XMKQZQK2SK-\@0g];>YA8YR4\T&2.-.3SSYWdA>Pa&I\\^BZY7@&B
Hb^(cNeH&&Z<8/d=J(^<,7[?1Sc]U:RF35C-eA#+fV+].VMV4DF?HC:7]#04\+8C
,HGdOM?((e4>GGS@Pb]f(,6FR?-\GcFf)aW7\C#O2IZUXcY)/58,?aL_KRDWa#GV
YCEfY5)La\[g;E#(3dgZgY55WI2@+D:Z9+0KDITcSG9cTV1XY<_,KH7&FA7O.CH+
O0Y.5KVVOb@b(YWFAT05G@2Re#1>Q2G]bO#A8(;b[g0+ZQ520dN6R<3.N)gM=B9>
7</-5LM5GS^SZH/GO&#V>e9>RO96E@^5,GWN67,fVTKQ/ZGd,HMeCLg(^B(.HV&S
;-1Y6cSSY.S;6YU1c8^fY(Z_Fbe@\4Z-ZXg/KGZFG](;=\0AXfe39Q<+^KO,FD/P
4R90_+gC6af/^Q>f#-c?5cUJeDg89U#O,E:+Qb&#[5RgcZ:PK4b<15(g/49E=G6-
1<(TDbZ:P+5=]PW+^W;)3.PO_.9B;0JfZ&2)L)CLY/C79fF(C\c:JX91d2B[4^DJ
M.f99-+IL,HfOg-;97;-#(D:-D/_6)SI#V:(O,Fb7V/SbQ4N/J^7M\U&,#&)&=6R
H0#RP)Y_G7g9gLGKgP>=Jb[#Y.&>.d3BQ4NWebUQ#>Ja-?Pd5RLgeVN+DZ9:FWcN
aFD17U2J>UWL&STTG:HZ5AEHO/J96D?2c8bB-66]#cR1P77:a1=T]KD\7^LQDK5U
\ZacG=CX.?f0>#&U?cS.Q/8baMF507A./G(F>=;NBG.bJQcA#49L9H60Y3E7Jd(Z
/>)eZR1T=O\AcS6U#V1^8G=]/K+g+.@\_e;7-^]AVWA\[HQ8cK9\JTDZD5M&9>f#
6aN6^c<]e7OJ)a4N1\:E56(K/TbC8/W&2?>L;X:Fce()I2B0EUBB==WT&JI6@DO5
(3\IBIM2^L_/,7eDb\gH3RL1b>KA4K1-DQeBW>K:Uc=3OVL3?FDMTaC4gb3eSO(V
82gFV2Hb4caHUgCV,,UG<cE@5C1ZE6Hb-TB7VD9[_-TdJI4>XW:OPD_-U->c-8aD
B>TfJ>,?[\T_^5UNA//V7#71NY+.OPU2N(#[UV+BY^d08_]Ce.8=EW93\,FF)-0F
X5U@,F914eB7M+WI_QHWJ>8T:\f6Rf(OC,.2Q/WRI0O?Gg4++;:_2E\&M:R\,=M;
d\)/.aO@X-J#I><CG97T6#AOfeG?[,c4:(.\c]C6>PKS_9A4=Yc2P;=):,&+/7;c
YXT8<TBJ5a>;Q#=b\JV,)ffBQ/a(0TSL,b8fB,80JG:dA-fb#1R<QFQ<]U;HX@d2
N3eUb+09CVKD.D]bL?^?;3U@8GOB,>R3_VXRU^7//7a)^,<75g,cc11)ZB4E<OKU
bQ@6ZL?c2785UM-D.>ZPd,J;(<X30>.;3#/7#TXW>^b<>=W&U4b=M@:SD2cUNYC^
)]J(WFH5@1Sc@/&]+aTOOX3SJ+@G#K>E^Kd&f>D?e-d1>TR>&PY.X6D\7-=L=cAH
_MZG[CZ+d[@;=P+@<82&[bRO];]O4;-9)Z[WN?D<^P_;X]d;#I0(c0K.[Pc7WVe-
=WF@]/F/>cLBD.L99c<8[37I[fW)8J6H@0/b[-.8.@WF;?<Z46b+0Ca&=ZJK/4&Z
-Q8Y-,(?0E0MP.b[<&HIZ[FEEd>B;W]Wf_Ca^]I]WeXGg<R@_e.JYKd7@4^aNaGZ
GWb_,>0f=)-4-fW::YZ.&L]?>5?U/L&g4Gd^>_6)<<E@B:3PPGEYFc,S,Y8e7a])
GXbg^b3AGaF,8fF_P;L_Pd6\_^EFf?#8Z=4cOJ0SGJ(@LLQQYXbG1)NL&-YYe_TY
V[SSMWB8aZ2<Z:35>+dB7R_,U(4<+H-C6K2HC<<e^KGZ,/f.)cS\#d7X#K/)#2UI
[XBQa8#Bf<-@^7C3NL_Ad5<,=O<,g_Y=&@E&\7GTUA3QdI)SY,K=Hd\4OR1fPfHg
^NA)K++CA^3cW];b;)9&PCZ?E^56bG>A-e8:IYHLQR)J[[c4LHEV#/+eEdX(E3De
15?@-Fd4EXQc_fQ^2NQbZDL+8a0/;HF??+B)7Zcd30<fK@5FV-T(DKbHHT_3KVdG
FU)&Q<^ISbbd8\bKX/T\=]&3V?VAEC,OMRU/>ScOL.)7R??.2c0_=X&(\V3LW4>[
f>dBRZJ]J.UTd4T8O6:\RUQFADQM0BFged<(1?EGNE[U6]VXD7ATE0;N,6QN;2VM
;4814b\>5\7K&X(-^X;D2VN=&Q&[UB77e6LEf#G#BUT)X9gL;^4VE(KHJHe694If
A(.f(\(FF((ee^_._d<&S_+GdI^J_;d1f25I.3LE-#bHT7ATa_X3#RA6eEF\dE[H
aC&W:CI^V:dYaH1U4RM3#(R?Db:ZNTS46[MMSH[8GAG3-6SAH(6J(Eg01_><;PTG
@F=:OO6X0])JB_7HCJ=J,daBTe+(QLcI0@#T:gIYdg)#@XE?8PWd0,>9[/dJ3;KX
d(2NFGKZ.ITa[[P_:W)5(O2]+,8;5^bGb1;A&^2)c;=K#F>0A9g:,=XMSc_.A&B\
+\VA[[E@AF<UJ1E/@<L&.;70[UF4D7]1NI[J=)Z#)^OCS>[L/^7;a>VF^NGM.UfR
YK_D<Le2Z,MH:QD=-f?;7C;I<S3dC[@;3?/Mg..O3?RcgOJM7gAdCQ=e<76.)4WQ
9E;,BM\I=dVXe4bCge3HV4?=0@Z2cC]4\+OF8/2?.(<#6)\1&ETR8;a;B^HF.2WO
c?=)DYUccXEQF2.cV3CP5W&(2CXUdR_U>/Z.NU^D6g5aK)TZVU[Z@JY+Q4S?cW0/
WO@-MZg0f-EHa0\L.S-e(\F18SYI\WZ_:+#cOP6VKWX_C2;;,[F8T7MPL-/NJ/^X
f5C<G7D26B+5SU912a_IXbA@_e=F[(#J.g;GbD;HcN#HR17fLU8-NfQAgZP;eQA8
5?OPb),QR-UPc;>4Y)A/G/Fb.T+J]/eZ(;/HLcXORcIY\/-8IGXIJ-5a@^M1]ED_
\DB>3T>(-3;3c#4ab:gIDMc24D?C?4#A5BQY)#MGR9]-J(4N//^F,H&^[5XZ.H&e
NWWbGP2H9gE&eT4:BP;:BO8[9Qg>6g7VDO]gE;0bb+,5J@V(CXB7\<>aL7XHd1fZ
fL0fQX,HEJ(0aFZHgH\B]^2CUMUJAecPCNR:D<gQU1_dfGCOCS\bQ;bdYdNNNR>^
^5(NEOFR(cd;MB[,P)-0(8F6LKEOaPAXHWdWP\2Y+YeD<5P6&0b5N1gQ:L_b3Ng+
A.67UM<O8>Og?&c#-aA\5H_1ETcFSL7CTabO9b(CLX&1eeBG8W<H9Gf#D/AOP^ME
JK4c;GPd<L8<<X/(5]8ZKV>]_ZKE/G/#a-/NLbINJ5G-1C&N,O.2OCaO(Pc(4=SL
_fQ+_IQ-J5VdL.,IUZ^3/B0F?B73]Dg=(dKNP(((.;T?a[B,O7d/S)JYV_S/Q(E3
-;Cd87&FK<:=@QOfe-K_?Q0ACXQd-J0@4H92)#1RN]1J54S40^T3@_Q>N<5Q#0Z-
-0D_M7WcO)OMge+P8OfS<W/G?Z&;AdQ@+,JNc9;GS[PaN]_XVERG/@MbaPaWMALg
UD)Y=[&R;Pc.c,]&RGZSE07:HE2f_0YU;3EBJ#\2;g>bcC/\e<IceY+[NI>Kd;KF
F&:TQ#CASV/21<UXE:e5H\CJZR=6Z/@6<X>1[)]I\^WG7.LOI97MIS+gJQID:3_&
.4E@A>-P#9Q2&FK3L/e(/).]H2d6K+G)XK@&f/?gB,044C\cXX96@0#L7C@=D-8<
M3#\a^?EJXUQ#dR&MGFYN@U/3K8=VIg=E.ECN4C+MR^V-a5g;ABZ8EL(I04U5[0b
<T?.=8aSJ^[_HT&-M=(J8#N&0+g,6V16,&9bNF50&X5FI2aQP((/JQ;HBdJ>0aMD
FaR-Ca)Fa<;IJ^AAA7Lg,W_^8(8ON[09V>@9D6CB=aLB)=Y.C^6/CId95KR6baBD
Af6Fg2@J21U8BbbRO7+9(SUd__KOO]/OOZ9X5fJI)]L[g06:/8V6/aY&4X0cgY#?
4e-Vf,2T-7#&ZEc/Ega-YbK,AOX6S@PFY<N&E@]5.D6M0R:UYR),8LTe2W>,PQPV
T)--Yb0fKH\BWOS-^A#-&,8#S)(L^H<ZC1T0#E(X,UQ?D+eb8>W/5UR]:1B>Y?CB
eVQ;_OVZU@Z2f#U\S,EG>=V0._@aa&F?gWe?BT)JMR1UXK0S6(?2\S\W#WPT,P^X
VPd_&O^]b#=K3_7)<\4/F#GDJ;FCec;#3<XFX&f3,gGR&;\RHV^7XKFO=_a_-_fQ
H6X(gTQN<BTP0Sb8(ZNCWSd/=-[0e[]^1L_.6aEM-&[N>JN@PL_(:#HCW:b8QW))
TTBW;VJ99F,BgM0-^:<2eM5<_JD=68c._><#P:DJF@Z\7fE^b^MQdBbPe6I&3]B8
-JY19#P;-K5B]YR2Vc1eTDYG]IaE0/>aZ/=#3A/_cQbUBMXE#L,@=FQg(N#ecB(6
9ZI5JN:g=(QcZN\c>?EKY6CE>6V<RNd8[@T,51?_[Fa^:<AJ@V<(V@If/KbW<(d8
.WVJ.fVUdgSRXV.NU]Bcb]Ha?;POEA:_\J@RTCEM/V:ZC^&9bD8)FeONHZ3YHMO,
R6TEMDL;XS7,IC<WaeR,)dZJ6:7F=1^-[/GJ<6Ng4(92c4f2U[+.JJdTZ6AeIN3\
JP#8e;[\&G.Y=\)EZ0#(fTeEL3PbVX7I&7A,XCEM^:88^GYEg1)EOW)_0X(WMHa/
5G^&G1&L]C[-0]/(_V8.>@aIb>H\EYCFWJO/4G-#Y+f1LU3&6MbNLB9/gWa_IZdE
)FF;D;]088RXTQOVgSY[V#RCNC>FeGSHWbFIR\&B]8FCUfKM-^dNa^N7I19X[UWc
(M9D]Q892cB80/(/^=M..,2UEeDY>>-I=A@ZZJ\D01JGWJd-c0YX-0Q;FdQ[YX.0
;b:2R2>RMFfMM6@[/\ED:GBK-X5)AC.:DQ1,1T:SN:Qa_3)=;f8HJId=J99[YABU
]0)WN22SJPWcP?g#=bRGK1c&U-(BARWT=]IgbT9Fed+HE/0a,^]&^g],?FRcNE1Z
,_F=.LFH9D,cG;M\/cN,2FD)H#FB##NcR&[5N(H;bM^P)MZK=aU1]T?fFcg>>403
;]ZbZ#U9,I?7=@2N#H(JY.J[O:^7?XH^d:1]XZPN)P<_PNRUgM4B(cf.eI_H_:\K
S0\cPV4Q@O5N\dH?X72(VD@8)API5aK.N^Q1086=AS=dDMK>RU\-a9aeN9LQZY#g
Y)8b?EcWT(+UcDH/La-Bd0^c;+(LWaLIa^Y>AUVV+#G,47VA\a2<_.[,=AH(_a;=
@Mb/HTeB4b/8E8aU;b0DECXF32>[.cP(,#e/PZP:,KN>673]7<RH+#T6QDGEDe=8
8\C#c#cR_4ERd[]0.#Y[2_bR8L.GC_+UAVaCZE>0IeDdR&TW-(J<d7K91\7\)HT2
W\RJBEU8WMX\gB[De[#=X_V-(CUcK](UZ(^,Fd55U)MEJ^_64<5GJQ7NUK3&00\8
P7.b8c\c+=60B?CX?(=[5L1aY?6JK1]Y=^/D:^7Z6C5MBIXZJ4eZ/GG.Y2g;/=,N
V03T-T-BF:e2;(b8C4LfLFaFMb7AG-fdEX8=Ig\gK_J@PXH@Ud8Jd<b;,+9S\,=)
]8H22+(9B&6WFJ;G07De466:gc<F4RP#M6BUAA36=OI=7F>b-9C\BMFc:cEF>[G,
P.a:Ob87bbS(?@+NI1:-&UDN?3IP<CZ,KgX\=PV8,O\5/GK?Z43)8OYW8Z2]\5Db
1C[0O:@4bXF26E]Q^[dCY3GH.,,I16X>VGYR@)Z61MP=B7L9eJ3cL7D14^g4X72e
8^2A1P6WX2#,@Ifg+DB\UV;BZW;@KNNSdO#(Wc[K@(L1;:E+A</eCHffVK[T9@G:
:+=9C0[-7&&LTN::9LA]=M)@81G7L]U?OU:4=/)UQD^MAbM:>\=;FP3]UMe(M0+M
\We>/FS/6&WRS6=b+-RHJV6B[^4Y<&fWN3PS3W7((_DZ).VAW=2LbfS+0aa^G?@8
A/9.@(@<,XE:1)ZQ@M9+;=[UA#NeZ\SW(LKG&a5BT0cVaDX8QcSQ9UX=&5dCQ@W4
SOaHWIcJPH4Z3\3C)KL+XUG=X3a.]T+/9\&K5BAR5=bF^AU.0@N6T3B<D44g\CG4
1?TMN-R76\VW>5H=]aMAcOS#f8bXQ;<MaREIaV0^eE&#E[3T(cU:cA86S(>HM7BC
>a;3ef4.EdPNS9(CU0bL8D96gK+LQSWd6&72SZMV,/&QNO4\IHJ=?/9d-f,?M+;7
gWb2f@T^E4+F3)Ge/BE15Sf12eS75<C5bcZ[;6RQ_g2Eg(-@5;DA^Ydag)6APd5.
LX)Q7cH(g>C7gE@^<Q2WSR-+G=IQOb5_OC.P7Z;.cEf1G_gR\+61O3Q0>KFJZC,J
a&cL9E:+F[(V_B8c<#HeO06A5+D,?)?WXE#?&,HIHQ.a.SW(5aWZTBIdLH\K^+N>
\IA4SEV_[cXA&2)AEg2Q)F,PGeMe4DJa3)30\ZS;(HS1UC4;5Y5V<614D8W=:=QH
R_FRUL(;egB3PQPF0X8(TS1]9U<f@NN)3IeM_HdR3Wb]KFJ39XE^KK+(76C\L[)E
T5S>DQ:(I^>fRG<^3&P\Z[FH=Z2SQZ\EN;O7.Te7SEL:ONa^&3MIK.M6(;5KX]0R
#WUg,-MD1:N4PIM5.AMea75TKY/+GCLRG,WXI-W[Z;(O(\b8DQPI4g&V41]M+@gW
BTOF-:)](+g@)KT,fX:^RE&<H35dNFFM=?ZX10gc@#KI;F4B6SI@fSc(W@<P^9g3
C:C[P.WOWdJM)Cf<O.LY=);T9M/&Q=WU^URT?(c8/BVBZ2g(3EEeKHXOR_+cRH@S
689W&+)(^/7f4PMfGRT/_T,?XbEU/I-e[[)GSTL])bHB9I08-96OJ?K@1UHY6.F@
QL23C)UL?\H6G,T,97991,M(7NCMSaWUS8BVd]TaW3@07KIA5#H,202?@d;>KP.U
G)I7KfD4KXGM1)9E],<aPXIG_,7Z)_<#W8[Nb(,^W^R8E>4>aAg#?Y\2P@3gg<8B
ZfY&TLC=,XU<C_e)8bZ,R--NB8#K&6gf=-Pd:/BN29F)9X)FC)D_;P@8?/bQ+;VG
+>K[(RNMdXc[)D_5cO[;0-53eL12H3.WB>bM<BE4,;:A1#B(FcgO4>/.2&U9\#fT
AY<W(/If;P:b2aT<R-R&5P4C+Ka:],RcX8JfL]d^M+A2W1RKbA/+?YE^>fV<NQ?K
X2H+J;)K/<U8BW3g+fe[fQ3FP=.TgA(fDXRg7Y]ZGW8A,^W7)QR9SO)VAaJb;(g+
,2WK5M0H&[[F<OeUfaY(2)FV>2Wg>D)C.9DV.bE]+S8I5Q,\46Z=@DLA9Y+U26Q;
DB&gX9?5\+c?AeLcDG-&MfN8cM7(.dKSC^a-(&_R>=+I92N:(3Q9fQ7-6NGSHB:O
Z3-e:_df;#b=N0-RgG):^W/OBYB+A2#P1S>BU+B8+RX8DCeK6<_L[O@fK[[S2f8U
IM::#7MFS3?(O>V(4DA.Q)5MN:2&K6Aa_Ja,C4K5eda42[YC:M?<Q2(/.SV4QT#N
@gO-_NJ1<]3))#Q>#cY7V:?VA>]c+R]4.&Q03E](2+N1PfL&.2O3-R=g+6Z0d0J:
5\?D3H,?UHeF1f6+B7W:Pbfb@R9_U_CTA>3AL-NdRDD;N+d-3Y_CF830?M53YYC<
=[BB3TY_g&8IXNO1+K59Q82fOZQQY?#Y4MEBNRd;TgBQ\,5Z3[e\UgJK^L+[Kg)9
)?SA\?3S11.&8&FZ95X5YPbYfXDAK/T\W](N/@-7aU+R^H@7gA?)g:?,NE0>QR>S
(D=D;S4g56,I0G]DV;[DT+3NVXU<g<7+0CI6.:bZOAbW?D-PR>7g4eZ4GMK]VDM0
_DVB491J)dES#Y+/GQ6?\A/39ICU,(\f-:>GAD45X^/]I;_9781?MPd7_QM/<2;7
+./[)JFR>5c40(.19daD[9?)9J\UCBag@AKYH4A-7])AUeGX=A\1K:f\-fb;S\K@
LCBOC6fR>Da[4PS#DQ+<c;>R0[EKZ_9CN]UA)I5TQ3B,4595U3g&)(9EB9<GGZ)&
28P/YFFOgeG\=XWdf23cMXEW_ACdK)+32XM<:+cYg6KC-\NPX:F@3XXI?4Sb<7_P
UVH\A9eNMQH.;/4Q&<5a;b)WgIc&+fAfUO1<L/0c&EZJe/WEG1TUA.@?Ne&ZXJ)R
HO[UC(@OJL,934VdB4FLgfU=GaBa>S61F6K<M#7-2a8AU@T?0^afC<?/8cB)[5;@
0c19(CI:@8QeEfb\).IfK;9>]WZ113V+3)/:,G6OKB,,LT3/ggJf89B(,;a>&-C<
8L44PVJHAOE@I>\D#806Z3OV\[4abd#>0UYCWg4,:NeRJ8SQ0EBM^0I<1e1OY^,2
c/2#c<g#REVRf=K_J(+<>/P0[B1H7_O(7^HYZ&fDRA:^_FfZf5P,]=_SF5&b<T[Z
d+JUFDZS/[CSVULQ1B-e9H]OGgL5=[1AWUSR(b:]cMA?U8P<@=93<)5-W/5GfE?E
,aZP2B;2>J9g;-G<05HPe+bY1f1L66;gfQ@?a8OALc<O..H7DY>VOF.S\O^e2Ze)
:Z^>,]WGYHe28O=0X)TaO8K\?:W,E#?4aT:XVe9eR1H>^<WQ06@deYJ6WHR8:3LY
IcWOgD_A6HLOd0d>C]?P9BDX:^C(H5Zd<)Eb2Z18?dfed:FV+7C/FJ;Q=6DDE4X,
/)-CN?7NT+M\/M3G/e3X;@KNSA,bS)dE9.cIFX7bOYd6];:5J7TOB@caT0MAC8>C
Z3J05SQ92_#Q:<8\>aB>&/SK<V\9BA(.EA<,ST@6M^ZC,R-PXM7&Ef@RH./N\6.E
c<-+>H?2&4FD3OdY)F+T-_^<&L5aK)EQP,2cT_C-B,)bO+Sb[X/eZ8>(WeBf;?>H
4\&AC1/H00P7CTT5I@)D;J.VIB2f:J5F@c64N,-[fSBK.e-F9CRX0Y#EZHRF:XMB
X?&9QXXFJc9ZHC>0D]55[V,,HKD7^Q:U_98ZF0EP0=Z+FV2Nc3D;K[;P2;=6=baR
TaEZA<3^dBC1RMZb8W4ZO7E[6<^&CH32DGEOPe]::ITfcZXe8J:1,K.E@1a^[1e0
+LHgGg4H[P19<S#/EWfXV6HKe6&;)2[U9R5O6ZN5aD__V^XZMf0Rg1D\L1:T^(QQ
/Z.XZ&B?:Y<?[C1Q>1g@H<8K:J3_BFaK=LCa^&K:,9TN#2c/@)<MCEae@)IHZaKL
--SJ3#EG5N1#UO,YT=Q/_.S7E9Lf?d7cYF,,&;T[DK/ffR5+[8,>/UT]>8[d6I88
;C?\bXH0I7SG/U_f=F.a-<A3+Y3#K+YSH94BF\PLT[R76D=J3W<7,T/:;O_f2(=Q
V3^U09<[Y.#A:9_7C^dVf0QH1PC@N0V-e2b&gA<NO:b0&2L=&BK6^/\6c2P;5:aG
USfI<A)YG^5N13TVO:1)>=G:WM3(,WF9Ed1()UP8UMRLR&,1/(#c>^I&-/Y1<9S.
A+RBTMV^:b<0(FNE5V,PO=R=8C8X&:FZN:+g-AQ0DEUKf.f7d=S.IJ[Y6LC<dXc(
?Zd4SF-)5a1ZBTY[QQ(?8&TJ62Jb4[ZLX5>2R:@f\KRYZ+K3;\NM0DKYJ][864D4
d?UJU)?JbN38)]:<C7Q@BQSag(YY,4ZR-&1M)^GK,<A<#<f50_Y<>=b6C2A9\Y6S
:R?-,E8/83@31C/6<Y>>00;+PTL#F,&MRCgTGK-S^>.RE4\-8cI:C7;37PY\697P
.#bCE^C7GP]:Z@D)R.g4[LbS#YGW73Xf/:5Ffa0POLT/8VV;O611J,&48371#UL7
.bQW]OgD-O7A7[AJ<eN3MP[=#ASB3&c_>afTWIbA4)NBA#L(W(M=B]MGQIDQ6CAL
>2SX@MbI]L^(P[g/5YE8aB^1Sa6]-N0d5ag4[;gAg6NE/)Q;CRJQKY#4KgU#U<+R
OI)(>g[A+<a7O4b+df/62Q+e.64LRO88HW&JQ1LT0\>?G65d]gXd,f4LE0G:,PD1
;9/Sc3/,XYZAa/=Y>Hf@F\\?MU3M9,K+1<g(B;WLOS/66K986-cNCcgg>G(J>9-/
Q-PJ>V^.0M+<^G1EDa\-3Q;BR^DgR=VYJ9IZ_YUQ))V93S):U1Gc0YVJ;19(-DGF
M<S2-(PLFJ0S?+(@&:,\?^YeR=:\Y[BKK5G3/N<=)#,Q&,FRYU&/)^US^4[g?51f
YMM16P?b3@UU2+2@,.WP/K4QZbIFCSc4#Be[>2CUVV[_<F3LM>0WI/4_A4Z+1A0/
)S\)-44Z]@IBB5])+T@3\0P\\S2QG:GEP2?I0Ie1E&M\JO:T:/d>W\=NYXc^0@NW
Ua@LIeK[2PEO[D/B54Z1C#OO5c:3Ha3#<M<AY@>WZWbT+UMe5;04SKT/eY,BO:0B
:caIF\QB5QW[4_O2[\4dVK=[J.gHWH6cY,_eN:W<DW.&_R19FE#U-;712,4JL\D8
<M:.1@4)Q<1W5IMR.37K@cUS20I<)#2gc,c2P(V8>T6J=,01N)(I3cVO&0Y^)CS-
.(f8,8a<T./-0XGSIYc+7I-]WT#OHMC5[dVCB-E@ZP0d\:bNE^,(cR.?6;^=;L;G
4X\bSOY@-^c(<^[UeWT6:Dg:5^G:4/aBKL^C:HfY&ZPL?H;.=Cdb>#eA2I^BZ+Sf
&V3=B9fIJ+SU;SP/+8eW/3AD,GWG@]LAA?DB-@9aF5<>^Q.608,dR5G/I\U\J7C]
DZH9N]N[@26FMd6C^e5<9QQ9&IbC6U-3A];XV_3B8V;,7F_9;U#-S8]#Y^@:V4+/
KZFNIZLLJL9U,NN-2b6H_TbE6;8&##B]?O<bB0d4:E741FY<3CSJED_TA<Ha.+f7
eT90ET1[H_97-Fg\?2DBF/B^S-/UO;eT9=IXU56+_^>5U==a)V_)7[PZ)]ZUN776
FO3O[QI<819]OB<:O=3KJZ46;(-;P^;O_/S[WG?\c;)2[6MDFeU^B,N21/@:CI2g
)4.^:.GRgC?6D3;N;[L,+)b8]R7=G9=2&YPDYb9ca<3GPF\bNWD:<0_D>f.f&YRa
TQXXQ&R\<X(T&N19ZaDVDL7e_/X)-EJZY8bA:G\1<H@6@_&+,0ZdIH,GBB0@E[Q.
EZXM/;R]/Ue(N[7\_K1I:.[F.C>&VNaP,OXB&L+_OB\5EGKeM.AZ_d5[Ade(M^Cc
F3fW,;?GR821JW/AO,QQ<JPJD3;7@^eUU,Y-4.g8G7fIX\g\GfXE-_-ZQ_LR7AVA
W5\gXF^_I/KFRAOXFDd\9fb\bf0-TACO?C9^M48;8.a1+39MHb,UO://@[=8]=cC
G=JDAH0H?Jb>4@(AR6N2gZRPBCf)\;\0/c]FI]DRHd25IaL,NM[N6=HE_+7b_WgT
35[U,+PT<RDFCM)#=?2,MT2AM&CS7]a@PTD1Z_&eK0E&070P:D6/;P_HE^ZI76N8
G-+HVV>43[^8R4c(UTNN;P07^@@9,Wa-DBX<C#Y1cQcL.I6eV3MZC-&I[XaBGc7V
(BB.I2U/[2DWRC0CIGIP)[a;7DZ1F=fd;fAA\UdE_fe^/^.ONP;FSg=L[EPDJ[DB
EXA>UfE5WA2W&S.7AJ(GeZcLX5ZH[,&G#7g[HfTDM+OCY/6g?&R^a]A&&)N=:gf;
YI98,-2,J2=R(XQd[Q:Yc;gLWPJJ)_Z6/NPH&G20VK77V^b^1>:R4B&@S5M\JUF^
Q[bHHH&2&L#_J1C95/-4cG<8\b(9gV<7]Z_XCM<I/Z?Bb@&)Bec64R&43e?4eB?)
ZTZS1RQSR[;F#4GfUUXgA]0&L:(5BKNF:[2bX1c4#M2+c^P&&^]FZY1>J_;?_[?1
G#/1;cQKHfU4Bg7^CM[;)?XcfP]V3EM.1Z39MRe0:DPG,GYE4SIRLa@2]?Y(e7Q]
fG7W0fbX?HK@G9JgT:T@-L-f@/,8aZZ8WKGMO@O+W<Y[(HG;<@(C0XdKg6]7@a6a
($
`endprotected


`endif // GUARD_SVT_AXI_SLAVE_AGENT_CMD_SV
