
`ifndef GUARD_SVT_AXI_MASTER_SV
`define GUARD_SVT_AXI_MASTER_SV

typedef class svt_axi_master_callback;
typedef uvm_callbacks#(svt_axi_master,svt_axi_master_callback) svt_axi_master_callback_pool;
// =============================================================================
/**
 * This class is UVM Driver that implements an AXI Master component.
 */
class svt_axi_master extends svt_driver #(`SVT_AXI_MASTER_TRANSACTION_TYPE);

  /** @cond PRIVATE */
  `uvm_register_cb(svt_axi_master, svt_axi_master_callback)
  uvm_blocking_put_port #(`SVT_AXI_MASTER_TRANSACTION_TYPE) vlog_cmd_put_port;
  /** @endcond */

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  /* indicates if user configuration has been applied from the command layer */
  bit is_cmd_cfg_applied = 1;

  /**
   * Request port provided to get the snoop requests
   */
  uvm_seq_item_pull_port #(svt_axi_master_snoop_transaction, svt_axi_master_snoop_transaction) snoop_seq_item_port;

  /** @cond PRIVATE */
  /**
    * A reference to the cache of the master
    */
  svt_axi_cache axi_cache;

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  /** Common features of AXI Master components */
  protected svt_axi_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_axi_port_configuration cfg_snapshot;

  //vcs_lic_vip_protect
    `protected
(0&KXDJ6HO[&-g?O_3_7.\VcG@_1Zd-SPNc8VSBD</#4?a/d5T/,+(+-,@6e8O)S
==B8-TIL]XFKC)Zd]I)a9H(/)95&;4fWI@AF@6>/.Q:NAODKWW42Tf6_30_]\>4Z
R/@9DHa^b9Xe+f/;>D/0^/C3<DbOF-5/#3A0(CUYfU)d&:c<R+][:3ALN4O)L\;b
\c6a5.NeI._U\AJCPJN,;9BDM:SWBAfV5QDJO[2:R;DUU3Oa&TH:H5Se_JR5gT>T
W&/B\0,-5#Z&TU-3P,/M6)5?#ZJ@c6LB97aFdZP7Qg+LD@a1C-,0B7eNQO[][(Q@
B(L5BL,4f<8A?10YA@4[(R)SI-(<8LQJ@+8Y&#GeeE^3BSE2M)?9K.b&Weg.dg8E
M4Y:])E#fZ&FH=#M6U;SX;]B7?I#)P21]C?Y5D2D)GCd.<Q/PR>^)-GQWOPH>U_E
FY.6A7I>\ggFBSggQ0O,8d4X9J0+?P/PIF/PO72D33B-3F/8.5J@G,Aa[eRe+JLO
_]U0e(e@e5>dagag.X.IOYY2S9A2bYYO:QC92VV6I@L-G=N4a=/1BO2eGc;e_fY]
0@V^G)>1T3ac98HF.Vb?3Uf:4RT[V@@5aJLKE(K0(XEIY:S\)+S)gRL2c1WIP(/8
SgYa_I+LgIWC8#Y[GJD3NcP(]O6[aZ:>##)bU9b([<XHMT9@b2G:^_Tb>B2KRF7F
D<+6=:8->G6e==9W9fI/&4g7^@a9XR>E6FJbU>3C9)T=Gdbb?&bE?N80=^E?ZeU]
+g.b^B=SU/:Q=&SEPV:AH@[DVNOF2--2^3.Q8I:]:1O,P4-Z,]0RM:K^g@>I0:()
)FIa/FLEU6#O8;AJKO;I0DeO?Z@F=>]S&S_>Dg],;AE?Q20C6&;,[Gef#^f#eeHA
-MN8(J#P2[C?+Jd[[T(K6UN+<63gd;XBecNN4U?#8>)O2<eMY]A\9XI[0IV5TP:)
H1[S<_&F\1_N\\+OT)VfD,QC#fafCH/T=L[XObSFPBDJQ8/F0F_APd]=X(;VOF?2
00U>:C2[,.O-5BK0aN_+:\UZf1:aWO=NPTAZ&QOfa;@WII=f5Q8/XB]LG1\5FEa[
CREH1M+e/UG\+Ha+2R&53.ce2ZS-;e7<9JK5L6JT:4->DTeJ\-c2F/<1VJdB/@.,
e=6WD1c#g58ZC.Q9N#]03Gce4$
`endprotected

  /** @endcond */

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_axi_port_configuration cfg;

  /** A semaphore that helps to determine if add_to_active is currently blocked */ 
  local semaphore add_to_active_sema = new(1);

  /** A semaphore that helps to determine if add_to_snoop_active is currently blocked */ 
  local semaphore add_to_snoop_active_sema = new(1);

  /** The process that runs consume_from_seq_item_port */ 
  local process consume_from_seq_item_port_process;  

  /** Variable to indicate if the consume_from_seq_item_port is blocked waiting
   * for a transaction from sequencer */
  local bit is_waiting_on_seq_item_port = 0;

  /** The process that runs consume_from_seq_item_port */ 
  local process consume_from_snoop_seq_item_port_process;  

  /** Event that is triggered when snoop is added to queue */
  local event ev_add_to_master_snoop_active;

  /** Event that is triggered when snoop is added to queue */
  /** Variable that keeps count of number of DVM Syncs which are accepted and DVMCOMPLETEs
    * are yet to be added to the queue */
  //local int num_active_dvm_sync_xacts = 0;

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `uvm_component_utils(svt_axi_master)

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new driver instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, uvm_component parent);

  // ---------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
  extern virtual function void build_phase (uvm_phase phase);

  /**
   * End of Elaboration Phase
   * Disables automatic item recording if the feature is available
   */
  extern virtual function void end_of_elaboration_phase (uvm_phase phase);

  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads like consume_from_seq_item_port()
   */
  extern virtual task run_phase(uvm_phase phase);
  
  /** Report phase execution of the UVM component*/
  extern virtual function void report_phase (uvm_phase phase);

/** @cond PRIVATE */
  /** Gets the active semaphore */
  extern task get_active_semaphore();

  /** Puts the active semaphore */
  extern task put_active_semaphore();

  /** Uses try_get to get the active semaphore */
  extern function int try_get_active_semaphore();
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** 
   * Method which manages seq_item_port. Sequence items are taken
   * from the port and added to an internal queue.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_from_seq_item_port(uvm_phase phase);

  /** 
   * Method which manages snoop_seq_item_port. Sequence items are taken
   * from the port and added to an internal queue.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_from_snoop_seq_item_port(uvm_phase phase);
  
  // ---------------------------------------------------------------------------
  /**
   * Task to drop al objections if there is a bus inactivity timeout
   * 
   * @param phase Phase reference from the phase that this method is started from
   */ 
  extern local task manage_objections(uvm_phase phase);

  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_axi_common common);

   //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void post_input_port_get(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param device_id_queue A reference to the ID's of device type
   * transactions which are currently beeing processed by the master.
   * 
   * @param non_device_id_queue A reference to the ID's of non device type
   * transactions which are currently beeing processed by the master.
   */
  extern virtual protected function void post_vip_randomized_xact_id_update(ref int device_id_queue[$], ref int non_device_id_queue[$]);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving the address phase of a transaction.
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void pre_address_phase_started(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving a data beat of a write transaction.
   *  
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void pre_write_data_phase_started(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving the first transfer of a data stream transaction.
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void pre_data_stream_started(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after randomizing memory update transaction.
   *  
   * @param xact A reference to the memory update descriptor object of interest.
   */
  extern virtual protected function void post_memory_update_xact_gen(svt_axi_transaction xact);

  /**
   * Called after pulling a snoop transaction descriptor out of the input channel which
   * is connected to the generator, but before acting on the transaction descriptor
   * in any way.  
   *
   * @param xact A reference to the transaction descriptor object of interest.
   * 
   * @param drop A <i>ref</i> argument, which if set by the user's callback
   * implementation causes the transactor to discard the transaction descriptor
   * without further action.
   */
  extern virtual protected function void post_snoop_input_port_get(svt_axi_master_snoop_transaction xact, ref bit drop);

  /** 
   * Called before driving the snoop data phase of a transaction
   * 
   * @param xact A reference to the data descriptor object of interest.
   */

  extern virtual protected function void pre_snoop_data_phase_started(svt_axi_master_snoop_transaction xact);

  /**
   * Called before driving a response to a snoop transaction. 
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void pre_snoop_resp_phase_started(svt_axi_master_snoop_transaction xact);

  /** 
   * Called before writing into the cache. 
   * 
   * @param xact A reference to the data descriptor object of interest.
   */

  extern virtual protected function void pre_cache_update(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
   * Called when there is change in the state of the cache. 
   * 
   * @param xact A reference to the data descriptor object of interest.
   */

  extern virtual protected function void post_cache_update(`SVT_TRANSACTION_BASE_TYPE xact);

  /**
   * Called when barrier_enable is set to 1 in svt_axi_port_configuration and
   * associate_barrier_xact bit is set in svt_axi_master_transaction class.
   * 
   * @param xact reference to the data descriptor object of interest.
   * 
   * @param barrier_pair_xact Barrier pair associated with this transaction
   */
  extern virtual protected function void associate_xact_to_barrier_pair(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, svt_axi_barrier_pair_transaction barrier_pair_xact[$]);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_input_port_get</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task post_input_port_get_cb_exec(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_vip_randomized_xact_id_update</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param device_id_queue A reference to the ID's of device type
   * transactions which are currently beeing processed by the master.
   * 
   * @param non_device_id_queue A reference to the ID's of non device type
   * transactions which are currently beeing processed by the master.
   */
  extern virtual task post_vip_randomized_xact_id_update_cb_exec(ref int device_id_queue[$], ref int non_device_id_queue[$]);

  /**
   * Internal method used only for logging and playback.  This method is called by
   * the consume_from_seq_item_port() method after detecting that the value of 
   * suspend_master_xact is reset, but only if the overlap_addr_access_control_enable
   * feature is enabled.
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task after_suspend_master_xact_cb_exec(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving the address phase of a transaction.
   * 
   * This method issues the <i>pre_address_phase_started</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_address_phase_started_cb_exec(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving a data beat of a write transaction.
   *  
   * This method issues the <i>pre_write_data_phase_started</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_write_data_phase_started_cb_exec(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving the first transfer of a data stream transaction.
   * 
   * This method issues the <i>pre_data_stream_started</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_data_stream_started_cb_exec(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after randomizing memory update transaction.
   *  
   * This method issues the <i>post_memory_update_xact_gen</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the memory update descriptor object of interest.
   */
  extern virtual task post_memory_update_xact_gen_cb_exec(svt_axi_transaction xact);

  /**
   * Called after pulling a snoop transaction descriptor out of the input channel which
   * is connected to the generator, but before acting on the transaction descriptor
   * in any way.  
   *
   * This method issues the <i>post_snoop_input_port_get</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must call the super version of
   * this method.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   * 
   * @param drop A <i>ref</i> argument, which if set by the user's callback
   * implementation causes the transactor to discard the transaction descriptor
   * without further action.
   */
  extern virtual protected task post_snoop_input_port_get_cb_exec(svt_axi_master_snoop_transaction xact, ref bit drop);

  /** 
   * Called before driving the snoop data phase of a transaction
   * 
   * This method issues the <i>pre_snoop_data_phase_started</i> callback
   * using the `uvm_do_callbacks macro.
   *
   * @param xact A reference to the data descriptor object of interest.
   */

  extern virtual task pre_snoop_data_phase_started_cb_exec(svt_axi_master_snoop_transaction xact);

  /**
   * Called before driving a response to a snoop transaction. 
   * 
   * This method issues the <i>pre_snoop_resp_phase_started</i> callback using the
   * `uvm_do_callbacks macro.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_snoop_resp_phase_started_cb_exec(svt_axi_master_snoop_transaction xact);

  /** 
   * Called before writing into the cache. 
   * 
   * This method issues the <i>pre_cache_update</i> callback using the
   * `uvm_do_callbacks macro.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_cache_update_cb_exec(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
   * Called when there is change in the state of the cache. 
   * 
   * This method issues the <i>post_cache_update</i> callback using the
   * `uvm_do_callbacks macro.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task post_cache_update_cb_exec(`SVT_TRANSACTION_BASE_TYPE xact);

  /**
   * Called when barrier_enable is set to 1 in svt_axi_port_configuration and
   * associate_barrier_xact bit is set in svt_axi_master_transaction class.
   * 
   * This method issues the <i>associate_xact_to_barrier_pair</i> callback using
   * the `uvm_do_callbacks macro.
   * 
   * @param xact reference to the data descriptor object of interest.
   * 
   * @param barrier_pair_xact Barrier pair associated with this transaction
   */
  extern virtual task associate_xact_to_barrier_pair_cb_exec(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, svt_axi_barrier_pair_transaction barrier_pair_xact[$]);

  /** Gets the time at which an address was invalidated due to a MAKEINVALID coherent transaction */
  extern virtual function real get_makeinvalid_invalidate_time(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
    
/** @endcond */

  /**
   * Returns the number of outstanding transactions
   */
  extern virtual function int get_number_of_outstanding_master_transactions(bit silent = 1);

  /**
    * This method is used to get list of all IDs which are currently under use by outstanding transactions. However, user
    * can choose the type of outstanding transactions this method should consider while extracting ID of active transactions.
    * "mode" and "rw_type" arguments should be used for this purpose.
    *
    * It returns '1' if total number of unique IDs currently used by active transactions, is less than all possible ID that can
    * be used by an AXI transaction. This helps in determining whether randomizing ID field of a new transaction which should
    * not be part of the all the IDs currently in use, is possible or not.
    * 
    * @param mode Type of outstanding transactions this method should consider while extracting ID of active transactions.
    *             Currently it supports following modes (defined as string) ::
    *               - "non_dvm_non_barrier" => all transactions which are neither DVM nor Barrier  (default)
    *               - "non_dvm"             => all transactions which are not DVM 
    *               - "non_barrier"         => all transactions which are not Barrier 
    *               - "dvm"                 => all transactions which are of DVM type 
    *               - "barrier"             => all transactions which are of Barrier type
    *               - "dvm_barrier"         => all transactions which are either DVM or Barrier type
    *               - Note: if "rw_type" is set to '0' then only read channel transactions will be considered for non-dvm
    *                       and non-barrier type
    *               .
    * 
    * @param rw_type Indicates which channel id width should be considered.
    *               - ' 0 ' => only read channel id width and transactions should be used
    *               - ' 1 ' => only write channel id width and transactions should be used
    *               - '-1 ' => common or either of read or write channel id width and transactions are used
    *               .
    * 
    * @param use_min_width If set to '1', minimum of read and write channel id width should be used otherwise maximum.
    *               This is applicable only if "rw_type == -1" i.e. no particular channel id width is specified.
    * 
    * @param silent Suppresses debug messages from this method if set to '1'
    */
  extern virtual function bit get_ids_used_by_active_master_transactions(output bit[`SVT_AXI_MAX_ID_WIDTH-1:0] id_list[$], input string mode="non_dvm_non_barrier", input int rw_type=-1, input bit use_min_width=1, input bit silent=1);

  /** waits until master is out of reset state 
      @param mode if set to '1' then it waits for 1 clock cycle after reset is detected deasserted.
                  otherwise,         it waits for reset to be sampled as deasserted and comes out of reset
                  after waiting for the negedge of the same sampling clock that detected reset de-assertion
                  to avoid any race condition.
    */
  extern virtual task wait_for_out_of_reset(int mode = 0);

  /**
    * This method returns list of transactions which are currently active and pending inside master agent.
    * 
    * @param silent Suppresses debug messages from this method if set to '1'. Default value is '1'.
    */
  extern virtual function int get_outstanding_master_transactions(bit silent=1, output `SVT_AXI_MASTER_TRANSACTION_TYPE actvQ[$]);

//vcs_lic_vip_protect
  `protected
.I.IOVH_W]1HHMNc])U_3bR/fKA3@;36)AJCc<1Bff&T-TH2J5LM6(7N8H8;\?2e
<SA@M)@=.-AW245SZ,IK;#bH.fY:[,LIYNZ[GH5b)K?X,838_g_1?4K==OD6DES3
e9W@8302Q3AYJKK&/<f#a5gZ<)2e4Cde3/M9g?E\CF/(.#D>SFE7Z>+A[f5_b36L
HV1^=f_4]>>FCK8<=<:eO8@#f:J61c^]P1;Q&P7J6OJQb4.3)=^(E\QES@OaQ(QR
;^YSIUL#bVZ=@GCCdbO\?+@#6$
`endprotected


endclass

`protected
)LeMPba\a?F&M9S2=SR\2F116L5[6MZ+\3:;9FQDRB8=e68O52_Y()^3;CI[97fd
+.7<Q1P#@_UI?1(,M^;W@f&gRH0W9FX([&HMWZN+[aZ:b+C/-\,VIO-_0<R\DOTM
[(GIXGNJA0MU85Q.cID4_N=R^9&:98PS:;<(I43;1_,PBeQ9VX+bb;[e5,DfT@80
ELE6>N9<^PIUGI(CFP-3WKKa5e-ZT6;LL>fBc/=J^,WJ^S81;HS;#L2VX\(CH.KJ
U(3C/Ld:&#BRT:VEI7GQ+=2d(Q<<W[FGbF7T@Z8(SX[_gF\>\#W6]:W&9102fX@M
^K1EM@D.\8b?McFe6TX;JcX)SB@QSB&7Z#3Ld=^Y]R[\S,bZ;O&2b[MJ&FMM64d)
U[CMg[aF7e7V\/V+#5]]CKF.+)aM5AIA)DIHICIK&^ZO;b;/SLSMTT4D.;W=&XDU
U<D&DQ68_:1-Ff6J=8U2..JD6>&SQGT;OZ3R\NGOT]NZ[cbK2L]I3f6(YFA3NJ9U
LI&c?FV,U8)N2.9RDY@>N-A6W#ELK?-25U&[&[0dQ>G>Ia5@eOLA-XfL&_KU(4)?
JIESOd@QYBYN/$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
,^66MaCB@Z560HV_gc/d/-^S.5-8OS=.K]XN.QgKIL,-c:@1JOSe&(6/[S25aP6+
#28CK[1/\5RAbc8OSe4_QeC#)#W?P3JDBH>R=9IIC0>DND_#@VNX^#eZM+eTTDa8
YXD(K7Z0@C(6[0.])WT&+HA?X2JXMZKK;PB/Db]]56XOGd3N3.4>/7?L#8R_g?gV
1^dcG-?]^>a9&LA]FWDT3,LTWG2C)7]1U4I39-U2D5TFVSNSJ@2X)&?\E:_MF=0g
BZ-c2+#QQVCgUE6)>D:OdJSUPC7YIC.2_D/<W^aB[GA25F0>LPJ;J)4/\]348TBg
gf0)&W],ZQMP++1V[bJR@Q05/R0G6VO\f4FX?LDFgd.:XQ4TIN7AVRbcRG:J_UEE
aVdOJA8)YgA?Z9\gNFU.ZP2U^G,;QVY9&R8Vc4M5S_JYLf/G0FN0eEbgIE+P?^NC
[d[M5;W\(;KaHK4JIE>)0D[9\<@70SDGb>.@cT:XEJ6V6aHTfe?#fZDE4Fe12+)D
,8R:F[cXN)W(KN,Q#_aOb+#4)EE8STe<UJ9_EeKRb/W[\DEeS\+QZDJ+>6=CeIUL
J+&c>=PR3RYP@M8L6D@CD&=2FC0J/3-S;F9YZe])W^1=dHQQ?_V/+c/CD.6V_45Q
(WK<GY_F/PX?B_(>=MKfXDF_:0>d0..)cW[?dEI\[E3G5dX2I0K@\f^9<+/fc4Gf
JdV_2d+IY7-e<B7_AB9WPQPOP[@(I1G4A[Mb2\@Z;R6\.JXEKc/_HK9_L))T.18I
4LE&BETYE9P2@4A4LZU9EZA4M]f3G429V=ET>K8W_Z2FMU_/]UW3TJV_7MaAN-/?
5Q:2.A+KP;;3O\.]H7T7H/4U+NRQ4K#,^0H.(XWVM[fJ6<]dD\f7T[gf^.]e:Z4O
b?a+<aR?TOJ^-dP>,X44GNY+_)]]g[<\]+AJYe0A&)&-d-a#D(Z>0I9N;4/T2J:5
X85I.D#D+<C6F&I,Q?eg2bg89V,Mb:_c-FV3-Xe1U=ZEMfK\&C(Y)>;^:(g,+95P
E(dZ7ETDaTEL^(VK&YT87)P.ZJGV9a<.d0+SBQT2EWc2#.R<H^LU1E]e;ZggU:WX
6X7C]4NV<03eEf/Y5g/a?8U<P&beL;@:<+,dE]5\HZ<Og#_F.Pg>3D\]NP2@Y.)2
><_;\K#^0&6KMd\J:=8Z=),&dZ_@/L:BHAbJ,N>ITf8;QZXFB?[8D,dEM9>g(HO[
>GQ[&-@d?HZR@L<@e8@B>:8g_\TNNT.+<V2=TCD&A]]PQC,Ib&gYK:?g96c@N\-9
E3</L,:LaROE_Cg)dII5ER[eBg9JM[VVX@XSNKLaLcEJOG-6FZ_-a,B(DI5<G9TY
:SR@P\S[S?1\3TSg]RD0Q),Z-_aI?FdAI@b>,&-,V=e4@52N&<KK40TK//1^0_74
ZL;7g5dXg28;J/0_ONKaN^^@-E=D#5G.&9[:aN.P;]TCAV6SQ>1fKa3_(3a^2^2S
c3D#&:gVVUdP3_N58<ZZ3I@1X@P1b?#S>OLX3\/VKZA4USde5&FN7D+e&O95?7d6
=PMS(dV4J)<?ZfgX[Bg)D_86V.N-F5.K#^>CPV6S(=B#KAE2EWGcFa/c<+_=NJc0
.d]@YELOWG9e,A@)FL#8g4gQE@#ACd)X-.45aFd__>QON[LWIGADW<g^SEAWf,Z\
b2+F?2;OSI<JfSH;T^HB6K6B=<CYM;,E<B-^\X+K7]bGc644JJD;WgI.0W]OcL?^
,,>Rb0eYZfcEc;^):L=efX.LS.M3,H5]Q9eC+HYL2W;,9c_BGBd-SDZ11LZf3WZ^
<?##DVVfEFC;MPe4M&3@<;-PUQ/?V(TM/+#g(,.;O/1EM\agS4)S8.)_U?Me7Q9L
dF(&21,.V)D4MD3[d8(#+<]U4gU5J5(@BW_a):]M<6^]LPI@Q>-&M?AX5?[L/;A-
PL3Ha.OJG#;O[dY?E/Y?Jg)=+5Xf&85XL&]bOPgHe>&4.:>X,?HgVHd8Y@&c5T(F
1WFL)1[XS7Q2=[>-39;5QQCPPZYE/P^[)<W_gf&/ZN[a6]#VC6#01YVLB4KBC)<[
:ca_HSH2DI70(HZXfL>O]H=K,fP?gb29+EQ3P3R=:R9[6IUJR&H##R&8QA?Og>CP
0.@]<\(;Y8C[6N<#I,P:[eWP)&H^1]-]_8(B-#\WF6-&[];<.LZM1@O[MB_3=].b
YDH.V0A\JC,G6#I5H9e_5I-aRNUA_S@>4<F-,7>U;TcQ3QG10XS1_0A9LE\U7PT;
e2;L=eNf;ZAaD;(OHC3?1Y0^<&NMOD><CMfX=TWI0V#;3-YG;92V/?N)0I3g[M>_
I]?J&MM7F7]C4EV?dQ()\VH4c?<A?OE<UXLJ=BIZP?D<GIIE-8DVA;0C^)gMI4Za
cJUDbA9AJEf2X?Z5&YLB)PJ.VP\gOVdXB:RW9)bf)/?PX19X^6EH769T?]ZL?LTX
(WeU#36XEQN3JXLgYIP1B\B_X-Z^@MHV6HaL_C-PFK66R6O?I>,\I,]0&QVb:H&-
_>T;^TBXSc,KK-X)-?F@)#Z;BCcLXU]5d)@d>T^,O0LEY\=,3/WNgf[AXEZ8=@7T
fMBGe=UBP0d_#I9Y\I;^-6462]-H=f^^34&R/@F,4\@?XMU_M@42YYZf(QINL-M6
6(_fB<K[>Q>ZWM2+J5JWbVTVMKJ/V@)^cI\A&1D9Ec<0DJdWJ&I6cL8;7J0N1JYG
[Z+JAXYJ/M^dS0,4ObAc^6&F79bE9KXH37E2Z^_BO5;+-d,2R@3[WLJO&XQ^-D_f
=:#R<BD0FNW,F875.L,c4bR89L78E@BH+#c-.JX#/aUI3EgHQD7^7;K:N5]eWc:)
:BH-5G=RS^9D?c>gC5I])4A)V<=WZ&>dV-GgIGR3.6LeRdJd_/>722VFg&d?F6S2
W7(7K;a_BQ^e?5W\BAe&/@3QN[F=&]R@:bLbBf^2+Z60JfAM^+E>XVcZC_MdS(#8
/2b5@)^:(EfSDM1b)R<+O4<^5WfM]H:#S?:Lag^fRH^H<-Jf.(^)B#Q[R:#^>LLK
.U_C074/[A0bX]R4E5P\7b)>#f=W3L(JX6#+W;?HN(0940ZLD;@1&Y8(M;.3CG6O
f28CgLDR_(F_JPI)/d(?M^NRRD9)HCMfM[?PCEF&\MDI>-GePd@=4KM3IK;(E_J6
0-G)6KBF>7@J4LPVg0:<S\CKA?LPO?-aJWZWE@dMgB):@9C7\M)X^/LT&,g>78JD
Ec+BJU]M@L;cSbSU.D2_a:F->B?1O_f>5,TO^31<\YMA_LHeRZg#V/?Q/4D+IKf[
<gH;JAR[QB4#T0Tc&SfTZP,F@.MX6\A#ZF5Y+9.KDHcLPQGdHfZ=/GL>=gA?2b6A
W,e>5C@c0P]2</7=>O4Z?FA+HQGGX6,gD(<OUKIg(8A8(M&IT::;d5c(+Y[WbH-V
Y9_:A3#dJ:aT90NP+PTf.[_fPMCbA\Fg#0W:1WNP7,fY]8Kd\K+N]M-./agTU.51
W;41#Vb^KASF2JeaVZ[7fO38C3JbdBB<10,ZD,U^0N(NB-\DFGMVg-T5&@K]O(<Q
3,_9(\KMM<\b<@06X)eCe2L+BOB5)Z2_9RX1<We8aPfe,dg>@<@=A^#?8[W-a-;E
KbY5R[J:I0YE[HE;X]MRK+N->Nc&BY66bK]^,<KFS[AM9fZY#7c=-:TG^+cF)>95
^K\b+>#)bS^Y\,SB:U5e3/NWLbMfQe\2M/dGV6,?@?A/#=SbWU5#/f.:LT]\WL(+
\[HIGeF.49+cZ[7]6+5B,B/7)[\E/[51-eLgW\#gP2DIYIbH76>;&EQL,IFN,S4.
WTZ2V)G[Mf6#e1J+HGd49HR-B0Z,=;_Ag44:f7?-LdD3HR-,54Xc]Og>R:cO35U5
H6c287E.\+=-9?8XePWY6bC7<:Z[A,)1U]77UL\1e[.g0G>IZgSI)ZbIJa^bbgLd
W3J80T4I4QZ3)XX;g]^HO>A0f#?AC\?KF(/G?4:E0@bdge+B\5=2<@2(Tba?V1B>
RS;Z)&fBYG(028fHb&GP^-5@,DYQN4LZ_Fd@+ZPSKDeI?8SQCaG)(P&K3_HSPN;Q
TJEF=>^4=:1C-<+D1T9gJ1PdF;+;>J-7&ce[OMVNT>>]Y<R4YS.fJ=MZF#:SB:IK
C6]C1cCTER;8<fb5_f4_ZN))4O@SCb\WI)/4;D?JGP3f=eU?4b]G/f]/FB[L\?A.
N0>=H#28<_Q>+d^V7d5c&X4_+\^&04;0Q@4U?d76CD#GI89ebHHXMKcc3(Rf0,GE
VfcaOeC5bd=/CPQY05),CHfZ3H;<_XLb,P83LHgR:53X:ef,5;7RT&Xc_/gOf6FF
^^SBX&1U<^Z\E.f6&b8]]YYBc2L&J+W+)E^^D-(30^?XD+2GLcAEF;:B1LdTK(M>
>@82&b2J\>:@=5]@MVbeDZ&;TKY(VKSN>eaPYL>+b:b,UK,aeH7,\_RCT<JE]LGP
,Q:@B>C6UE^U922cgaA=]cGRS<VM.)9X^b4,\<Q,29#(AP3<MAVZ0SB3Tc23MgU>
[(K;#YKK<YQ.=<;7&TAdAQ]C\]d/G&?f5<RL#a12Q_O<_6M5&LN288GG,><><N[Q
-T7Ke7L2a7ZdR7Ufg3<Y#Ee1GMT(/8G:QC05b0;G#5JbB1VGL-]=#@TN]O5(MYRT
)4.K?f6^R6]eLSGZJK+090FC@/3=A<&g<A,6C@]S:]Fedg:dX:HD6gM2Dd@If/c4
<A-.&C0L:;e@6^CX[(5FRe.EP2DFL8?:UVEc>/O.@KMH5F.N-Nb;_OSO632C0e+2
GZP34KgM]ZNQAJ;0^L6L-,;657ca0\3cC(S6_SV61&=ICO5EI))UXVeBY;:;T-H>
P/=VN<@1WV::0KUO>C_/A8:URFLVR<]eg5K07DG?e,:fPISf<9>3ULYEgTP(<(8_
\4M,Hb)[QMI(525.R-8[eVZG+E=DNT<R=Y.eL?.V@I7)9KV&FYV8S814N5f_,O_)
L)<.I8^5P/BJEa1f+WM+aL;&PG:bb1\IX\>fW6YZbbbETP-J3[02KMMDbIGO7+G&
:_W2S9@gdLPOE69(fHTD<f6W.>9OVC&66X5S/5OKL=7X)/,WBB?c&Sd[-Xe3<^[K
]FXePHUUTR)4I8([(\G_Y<:58<4&X]VdNQFL-V?a6)SR,C29KAdU==gS?]a+\Z=\
=+F<KHKF=675eJdY/^UXGT6>-N:-e6^I6H:ZVcd+19_\GdISXg4&\IK)g/_Ed5X;
\\eR.P.?#]KQE1<K\g]bE,Wdg#>B:U6;7AJSVfUI8Ia[?5gXX)ZZ?U4A4\A2]@SP
#BQVM<]B/\fI<@)<0.(LF=XN]@3)LZPe-fXDVPCX6S?[7C/dB>GC=>?Q-(U-F5YA
Fc003_;07X<17<b/eA:b5E/&,/.Rcbd8daLZK9deU6(TSO&g#9K4P=O>A<OEb(8W
J5L+CBDUed)028dZ=WOa-X+Dc3a2g7=:TU\b8@Nf(\2Z40H:VN4PEN2SfP3M-e->
aa7WZ&^d1.HEH+AdM15KcBW,(=/=bGd@c>2=+N,<&Td#+>=B0gcSG3g]UNa@e\?5
N4U\SAFcD^cB/;Q0fg3^CTd+^dE?VYXacX=9_J:+;/&_(bRY5d=T?OZ-1&4YEM0f
G_S9[B&UW<T@IC0E,\--;g&c=C#g1eaeLHD^:GM>3FOU^D1IUJ=2S:^AB@4NM9U;
]N,MB8;\/GP+3AS^?_dGgX=2PGO+S4d--IVL.XSG5UEC9f;&>Uc640W8U@=-3PSb
a(aT#@]-9+S7+I=(CKaD=099_b?I0:T^H)]TfI:R[0\#c5b9TI2cGJMW_Bg:]1KU
#M[.?JP5OE2^d_#&&A11Hg+I7cB^N,B?B.I<XTOV\_<=;)eLS._b7ZAM0SR3a1D_
XG9)]A0PD6Q<[<FAC@/&X91&^93=Z4M6#WW1[PWVLD_H:[9@2gbH?/5^O\-dXZG[
J3OXPb++<1=9T76c>g,F_:2>G##VL7F\AVR5XHbG=]ZD37)b-d_9QGad.D[g@3>N
J?NIFA@4MXB=&K\#(I-:W?\?_\YEYT;^S_2P]a_bOU^WSA,0bO#,E<2WYW68(-L.
/fGP=IADgeU7@HQ9V[6dc+UeZXb_B5dP#YUC@WY+)QFJ]BARBWIUa?GZg.66K9b/
FN[X^N])9g-_1&#R33189]\E2>R.;+7;G)BYPW--+L,eD=#2QVC]g&JK;:c#0)JQ
T?^,R<fV:LB:VdNe+eccf<_[fVf2<eaJ.HWF?dZ]PBY723<6G22ZNBPdE05OR3Wd
NdbLS+F.F^L1K:MZ84Z,E;DUc,8?E3NZ&1DPaVLFWdEHA33bK23g<ggcF^O(811O
+GOI=5U)]4aB>^C:=>0\,<^fDBW^G-M;S?YEF^,Df3(NTQ,97,>TFAHbEf=K1AP[
7S;1,U<c791<MWE4gKSE,D0:-/\)5CId4M(2.:4cP-Q--_CQ\C<8E-0=I(fZ-P>_
XM@Z(1fF#E;-f4>T9(3[]-O1UYSW/:<-81Y@35F,]KYM-Z?PfFC4c-L+0HI9;@D/
2)M?Bd8T?]8I,\UY9Y2UOZJ.,f6[CGE]^X:PYG/D;E3a_4d,:ZG@-.M]YX_U=D)g
g1R1SE/XKb[@WeJ3E.827OZ5c+840#7^IaW6b>LY>JT:Y9-#=T,H21O&;^dPc.X<
_,#0P.d4.)S9<cL-[Ed71;>HHTEH[:^4L5g,Z3E^b9RCJ2NZ/8RceA_Nf@E/4\)N
S=f+&?-MId6J+8&?AW(-C;b7\U;-D.6^RS+N-V:EB@RWceBDMe3DG,&54^F,MO,>
7,CPZD1PC)6O+.S37A4K@;a.a>b<3C(_<)ffb+N403?41:-YgDHa0Zg9f/VaWR?K
;(L8VH^Q0.dKdegSdBGE]fXdPNP+9fGTH=2#&Y3Edde)NTd.W#34f+Eg@4@0,M?b
DQ-N7:bRRQ8Q9<._Rg;Y[9aeXFE:@83)#)(UBL6cU)gQ,JGc><)Q(.U@c:[Y9-c^
^(Q:U/G420FS=MR((](?&R9[#d^7DRUeW)T&.;LDQYQ&9?33c8SI<]7A53&4D7U)
5bf1/M_U<WYI]RU/G6<9T(5HgUae@f#aE/F>SUI2IA&Eb\87?G)+M,ETTd0+Cb)/
5)PH65>HMe_dG0P)1g]8;<JcTSG+cF]3[g5P.aQ+@<I_+eG>Z3.(VF]ZK:.[5e(g
PIH5;<2\HJ4KTM=>GMBH7RTaA0Q=@=ae:D07.]XgUBK6+2=XX@MBFW1AQHGBV/EP
O@c6^OOCY4-308efG2cTQ>-Sc,7:_;c9Y,^HFJ&D#(J6O-9(bJAb<=-J]HSHSJIX
XSY9T/Ng9R[^I/Z@QYa^DS?SJ_,E>RWR0J?B2NeS^+8X(/F\U<FZ9JML_R1(Q3QR
](L&Q][(gIX]Q@KTG<XG&>]B[(32O^G(.,Se_+>4]Y8=,8XdW((gGH3\HBgYg\7a
EM=]Xg7=]#-d0(W9?HK.AC+C>>b19[I&V<)X25/]DI<ENW9d#d^U:]ZG^S?KB06e
CW7e/-5JRW[2N>_(FW59CfXZG,I55K.]7^c[7NYZ0Qc7e)OaX+)FC=Y),-WRdEW1
dAJUL7J_SG0^g(0GGg;CdCD4B^\,TQY[X[Y3[MGLAAdgERML:.VSR>/4FcD0/@,/
#\5ISK]@&D[UM[dZ=TNUcKGA[2^QV#URP>8M=]8U14Yg\9gRWC[dOb3eTI-,Sd6#
#X&c<39<P[1P\>J,I4O.]g.8C;bSe>\^:DVAA+Vfce=H\-N[IKKBZ1ME@bHC>a4G
Fb?OR+>;QeI-XYJLK=a0G<QYUgQ@M4-];DHKOC?ZM(VS^^[O<0YgMG/F:7e=87?.
UQ43dfPa3+V1IQMGf9bK:Rf&?8NfFDV-ba42_KaVQd7,QR0F6].;L70O39BSP]WP
6AHWC=@>AOR?9X6VX0dggKfQI7Z^>SF6X2I^5LPZV&eK58Q.W?cODO&LffMF<S>R
CJOE)X,1ZMCdd,[W65(4.bRWB5&QX@M=/ERFSOeZ&_CS07[J9ed0<C[g#;YCA:.E
]44_\CHYJD\bD/7TZfYa^IX>_19]8)P)\A1PB[KgH&6:?#=+O[Ea,cGV\(;M=RYg
L+44fa[2OQR3J)=<EL?.QZ,P;7GU9<64YK[gaPP8f0fE7X&bDA,Z<W?TU-?(OfN7
/&Cg7_\[I@,7^;#d:2B\:QR0J^NTAC+=X=K2,40=@8,-4P_E5TRFg7GR.1BR3cHL
XL[_.J=UBRFXdfdf-CNeR;SYNe=LC+ANYDC+B<]U2^:2ggRVFUEPN@2?EO-_Qf@>
d+]d)ef1L0+AP^84S4ebg1&.5a/B[#TEM>OAL->0=O;>IT1d=FP3#7C>VPLFJJ^0
HJP\I(24H/b9Y,R8MIPB)Td:/Z4X-@IL@.eSF/ZIRAT&/e?0Ld71OMS.Wfd0B;:T
(90W>T96\0H?A<OP,5Bc=Q@CeHdE3[TcQL^gHWW-0e&bI?[DA)2LD/cHELcUWg_(
b[G\8_F:&9\B)N#Jga4<&&0AOE1[6IG=E(Y\SK_A>@_.2E:G7,<F#A^L[,:6,=:5
C.FDD36X[IRBXB_P-V=<-S#O\K)V[ZL6@gJ-d(XK:DT0P8,,DT4YFTD1990;<DgQ
2AYaI_YT[dZ0Qc6bPS[>TRBg.EGQ94:f;]9^KgULd)^YBbI?FA+VfaAYVC#E<&O[
4&IM>.6@@=e/4,a=^G:D:R9/&(Ra^W@7Y\K=/L9PcJ@66&Nf3-+--OFf:;MK)=5?
+Q3ga+X[L/WES^YdK>;3S3ZZQ,g(Cf9.5/WZI>Q+(.9]bPC.:5J3LUc]@[\:IP,J
.APV1cff9KR2A\#f\.74\EY3a;Xb&)=[DQb_M3.dZVQ+:B=]VH_B9U&SSQ5)W1&C
5?0UQ</^\P.[F_=1T^[dO&HPI:P;@(::g1<H<\/1(O?:5f[?&9e5\=Z\40^0Y(UF
f:.A0g=IE1?=4:\<\]1@gWNAgXRa8=2B=)=bPA7D&00Xcg=4SEVGbFf3.874,4GM
\]P<+NF5SH(>5(3SA,7A_AL]I>_=Z[Z2X9D&McE7Y#7U)@PgE]c(\L=I?T#)HYfc
HbP?SXIK(Kf&gd5?M7IS]_@7)gN_+V]XKYQ0X8JRU[YfbS_CT;bVYX#207[[UW)f
@B5A(f#K_1Y^8W@#DUQ0<;b<W1K)gb(\>8YLN(@>EPNHM_0R6(X&<4\+/F49+@-T
I&2Pb;4LVE)=b=]I@UYEXP,2-1/<TO_b+>_=Q#TWIWa0/)?FbG6.7IWX8Ee>:>f_
RQNBI7USKJH#O,1W-c>52<F.R/7Uf.FZg0F8e2D+B)T##e8@]OF/a2/_6_1CRAN8
4KI7C:Tc_#\&ZFLK2?=W0@)c1H7_5B/>3-P)H.fOIJfT<Z#I@c8;/1gbRfB)]OV0
W,:-5@>bQdaAJ@W>01)&T:b+DG_W\e5Lf#cceffLQ+J806LeN>7RYLJF@g)=7@dQ
L&A^bSAWFf2,,)2RRO8FNNBefHC])NQE+a4T),gNK<e<ZYQ7F2>9XB\b@Rd7]L#>
-<8.XT].:B8&Gc.FEP5@9627a.A87@=Y+X#BQe/2.DC):IN7c;aEJ8Z_V&_^9LQH
(RggXg;9Mc5:FG(+B=4GYUEG1N>O]MLfW,4)?]5&SW?=M8Y59JFES3Z;a7JN07M#
3#FB[^-Ug.b>E@-235P>8SO2348;,EYa\0.cDV3>Lf7B6:(NdEF:MR&_?@bfV2Vd
#&6N:V>@H]ZY..2;aWd4McZ@GDHJR],7R6^A8Ng\2EN;D0gbK&N_+&3MEWJf]KUE
GN?egfSHQ5BLLcQbJD>e,E[QEQCN^_C]E11R7c53-FSAS20UX6>bBGGF>72@X3fc
CV@CFHHWFTA@7KQ_JD[80=VT<>RYH0\8.6Zf.T/OQI^gA:d8)=?QS<Mf]L6K6Q3,
6M3Ie-RJPP+@fYSLEe2&&gR+)47:A.MS<0//DAZ>(QAaCO5>Z<^fJ^@TPf5E1Nc2
GJOU\0FQKB1,NN:^R9(+Da21,K]0+d1T@E+CM)7+M;XLTWU;EaaJL]LZ9]<AR>L3
)1_T:>+Q-&b/_EKd-fb>-5O0&]U?=[\ce0#T0IGELEHXR3^JPQ&_?WY?N<J?9(Dc
P<Q_a7BO0H[,W-B57+FT3EdF?EQ8K&VEJA-f_7_7]-PaJfB2O_f\T74]/B5f0:7<
IEHV#NJ3=\2H3?H14)JAd9EW[P]&5>IB&&a#N,<46dW-5AY4T1<@<ee;5df;8<d>
f7IDZ>J,\&PYV-(0-=8\Y^c?;=<]0P:X7e?T@U4d_<R#G97B&=KT4.aQPGA\69]+
K<+[f[/@Z\^6XQ0,]C#C]G.OJ_Y[PA:U&L:9SVZZfc28Z(/T&,X:DO[4Z<Y1gKS#
-@ALP0J]0c@eceT.MWKLIg0bBJ&b_4&f?LB#=MJ48556U\:-Jd9DSY>.S]H48df2
DX903CY(Z4QPKF.0YZ]>0U9)&:APga&9VGIWc<HeGdc2AQ]8/962&L?:S[IG#)YI
KAD)+BA7+H8f(d13GH@S]c/-10Y0_+>[9CXe?R&O3RU5L7)ZB=a1,G<_b57?H)FL
/#WW_Y7Zg3HG5UcLV\[>._<6^NR/7]#G+M6gG_\&YS3//LSSE/30A-g&:/Bfgd>V
UHFe-4;\Dd0&]+^3:cf.+?fTD_06g(]MC7d.8+9[/,M9[,4/;)R-^d/cE7#,Bc=;
H@N8JAVWfG0=D\aD3cJ\aVH44R?D/9YSXQXe4,K\bSW+8(/J\H?R7L//].g4^.Kc
M[6M(ZU5L=1WNA<U=([5FaO/0g]Y0g8a[N,E[g8#ZA,_]ae1^g_(&eL:1YOFeYIA
PM0Q<>==OJR7,U9We<c(XX6.KT;KQcQ7+f_WQPNX#(4=VJMFgZIH?fR3(.[0Y=&\
a030@C^B:S3TF+?:<OEMIT^_\#;\8Gba][LLI,N>7R@V#f^/UPOI@:2MdIB2MU/\
L=TX1.\;B)ba&@&YK.Z@BTQ>4:c^XDd4gMFKR(a]70C/>7bGYZ4ZZ,V^S=cg]c_R
SXTX0?LW_3P?]P:+V\AWEeFTO2.&ZAfOf@8Y,POI:M6=&AO;+cE\PWf-\_5aCK7_
/VM;&((>QRG,Y9HT-<)V>6234D>ab1P(AL68Q09YIU0d\],&>X@#._[2RGZAfY,a
4;f[H<d(SP&ROMY@SO1.LN^4RP28Q3O58VAgc_Y)==<Q\PH.f,S3@dF)5d9#bF2L
4-a\1H3H+b[J?WVgDK;05#>2D11Ldc(/W&#[?BQXgDaARS-D44H/1#T7L&&:,:.7
N(SdbS(aM,;Z@L.?JA(5[_8VefMg,FSSS>DeA2C4M@[S:9>7-(L[ATJ+BQ2:a2a(
.@A8?NU[IGQc-TcU(1-20&:]KfT&=Y?WcLT_YRNb[R#MAH)aC1P1SC#f[OYQdK:g
ERRN.T,VM4D.<Q>IZ0)LN@(WBU0bAB@8XMI,W_:6GcV:MO7HQZA;,S/T6@)?M4=L
gWTTgCWgLQc0e\AeYB1..<0,R57^8IU/.BONBCTGSMB+5CNU.=YBDUL8bNIMEXV_
:P448M:77cL4<]55_a;33NNRE=/)M)YXE;D;L^a0g:9edCWdd,M(9=IEF=,G67#f
KFP[JJOJT4QOHAZ;H1^UIW:Iag@A3e0]@6;?ZUOI--^.[8;:SSY;KH/bgJYfc=,D
;/-Y\V(W#>,I[,?HU;BO1@c4c5Yg/(DA#-;2A7ZgS4K#6(]W)\N(NXE4W]\VSA):
P8R<RB0H]A4LIK&3XE0()#>9b^E&M15WWOPOfL==_C)J6RN079\A]2Je;G7W3]0B
R<V2FebL66ZR8:1gV7D/L2QRIJ#\?dN,P5\XQLMAK?^9@N+P?.d37:a:V&ATbIbH
1YR-eO]:JV2a/HFM5X6A\a:;d6=SHSEU,/.8##JNf.M]ZJSKWL#0>gQ-;>-@ID[M
9e1GTOL&e^Yd5J9AA(@(TbL0ZS(+.R#=A@[63N)#_0:I@.]VYS-Hg85>2D&>W]=7
2ACUe-4@1#8P^9&^,#^8Y9AHABLcV>MW([HQD:5XSS[L)ATU.Be.0#]^?]Q]8XZK
;Y9.Y8bM77_B;4EEbT;^29^:2Ogg:cKLa_CO)K^>4&MWCM^P9O/)W]g5MaAV\CAM
>C?M<@^A-Q38X;[ff_.gd<W3fR4O^6&VN[[TA31/HA<..;NN67D+^1PZ[15AMZ]#
g>B]-KB(Q,VS:5-,dTHS/-8M5;462<Q<U-(>Q(0Y5K&R<\]ced:dB5[[4+29SL<[
f0\TZ_EYZ4fOS[G2D,IV9XTc.Yd,FEY^[ePBEK\_cK9I+F7BA]f0N),S^F7)_McE
[Q]147\SEA80#Fc1VM4T43XcFR2DZ_\gFHT&NCg[dN98<YCdP-LTaQN=e]cf]M(X
)6776VQ>]eONe]8O8g[,@IV[TQOc@-ED=+JgGX,/VQJYX:PDQUC+P+2eR;W>B([F
VH]P2OaJ^.^Ub7a12(CT^]4MP+cc-b6.X&455>A9-AYc+_8R-[_bR.LSQ=S1WHba
?T=2-DUQfD4V(TRO#+C-2D5]_V7@N(\C8WHJD6SA8(ELc:S?..7YfHS\LU0B:_BK
ZD@;@2J71ED^H:QN+V4V&2<Q-F7D/PA\bTTF(d\92+fad7.O9S^e2I].^FL4?<(J
cL&K)aLAMXB&.PW7\<<X+9(d8D.[a/PG\(F<[X1ZAUGZI?^aS4W,/WEf3#KF:T^Z
a0<L9cHB4E#1T2Ug6L45^>[,&cO\G2F95:921;9):[K(-)5;+?B@CB\GR7PNDZFD
7NfQR=J,O406IUSHK_Bd74VaH;(-bgTY[Z<#gSWI)N_T4+Sf-CaFE3Oac-PMO(&R
--450Z7;68QQ,9[Y]d42VDT&\UDH-dUF9M)eYC+H94XF>=6Ie4b_U^\UGO#Tb)JU
cC/NaI23??)fa._7@S&@0\=5T,EA6YXU]=bSCF0#2Yc9GM0F:WT/Xfd-6&gUQ.M>
IW2.6E5+/(7=(R#Hed,.NTc<<7.aVKN;?6b+PcSdH_+ZDc[eW-&X:L(Ve&5+@9))
2Q:P,SCJ:V>Z=T3=c;_HCf@V,P;C<^AN#\Y@HcJK=8@_3E,;Ja-X[SU(V>AH-e0=
1T)\/[D72.aD7@G:A7c7G\.d6IT)E8>BBW>Dd?\bBfc+32fANeMXNG(fc:=-[48O
4S(aYK#D+L<Z\gd[MFb590L#)dBD9g]]@(+>6W_5+&2SYD2_B1QFN6^9ARW)_N3/
E?;+(aE/;+F^(C9@:@+[KRK52SB-ZD[)KG3#G@C9gEOAc=(\N,ZGT9W:W@[F[V<=
:)7E;WWE[a_7HT78C6C=,CIHM0Kf16>^O_fZ/L7\8^VJ:#f>>.XP95-U1=W9GPag
ZC0GaYE2:ZO=f,RA[/REJTf?XEL,5f@<LE<8U(Qe5S4c-[]#G,]VU>U?eV7O7b\3
J(?[MA#Yb@8N-VTbIL=EJS?>3F1S8:=2N_MNC^][[SRKCZG916ENCGeV/Z85\aKA
2AUT<@,&Z+;(P:B?#D3MbXV2eggEL@(I_AON>/#Gb>^DDWeEc+cfG3+?SSc&LST,
C+EP[O#fXJ3X(.#=>DdW-;d<ad_D8INR1fGJIEgO\1(gOC?Cd^6MIC4eB84O=:U\
ff-D(W@59IXSf.6?68ae(b](1^RRYDL7ADWP0;f>B1[DX?eMc((fVXCaQeS#_PR<
dJMFFP.&[)XW9KV?3Y;cg]TJ3Mb([S-;U<^Y+eG(3gB:MYYfKI4Q>.[F+ZF2N3,:
/76;+b?ZC9\#02T7JP/SO(^<,f:9MGWDcS3HYT]VSA.,OG:/d]2dU1O7c<Sd:Jb3
>>(TgZ?,MF,ZW=8c.+7D&SOD0O#^6d?W06>S+]UA#8VD6;D1f0HD5b=B8g&3#Wb,
A7CV1>>1KgN99OV#I\2Z+a2d1f#[OBfVC[cf]\BU=](,/1@CP#e+.eR?1PW5PI/]
I2_f@1Z6N@3.G.O[@R+^fV\8Z3aUG&FL<>WD?fK.+,QR.+=8^@S]BeV:1C(CNJHa
#\7g<8Ydf[G::<15]8R3]CF9;=.Q8&F?[MSZ>g;;@/JQg7,0W4]S5b>=D-ZZ4B=f
bcU_0;ND\:[Ka>GK\Q>^GX1:Y<HFTAegAb((.&e#P,EBAFJ?OGOB=Y+]9OJ<(@8@
;Q]g_\YB9V(@N1SLCS1Q(HH+9&+ACKHEB\d4g?1UJ6b(R4HM&I6P>?TdXa[\#P:/
=#GS?1gdR4I\d](JF_J+OIJ9Ab7]<Y;N1dH:.3d:>,KbFR=3WNN8.L\aFP5(HbbW
-##b9NK;OGZcIaZ5LM^c-S6&1f=XZ=f7e.YRQDcW&,8BgL;PRG@_#U[GFI06<H((
J<;Bc9BV.Dag7VfQ_E\B@.4d,cL2;\Q0ffE^fJ1VFGb<3_8#3:&6.)PR#HQ?PTMO
?NS#S0;I@W/XP/)fc9ag^8HXg4-FeDGb/O<:FJRW1U6VVZW:C5aG4RQ4OYg.3T#G
X21690(T+HEP]]BZCDTCQSO:FR]>Zc?]3Q5(LPE34^D5c8AJaS5UQ)_JFAPF,9#I
O1M^5MAQ1(8M4I<^G3C^,?ID1.V50PW#0^F8=b7(,;&(26IK0fbcP7/:A]TPE@d]
PO>MeRQQ;<2SXDFL+-PgPf^a\NX:].SN(@/SXSLK\1M=A<8T)W5G0HVH:.L=C@SN
@MH2;Dc^c@J1O5,O]^=&?L-K=eHdHYDRZ;-E^>>@NE/77M&R@_]12:,J&\@e:[9Y
ZS,Ac:&?;,I(/B)T@c78O;U+^e0=Ib5-7AFI4>A6EHEg#:Y\1>C9/Jb)c)7dN?(?
JT+6)^E046dE;<L5#@U#BOQF@A;]II<f#&(]8LCBK._0V\]9U1FTT>a&0fCL:P3\
5eV,a-L)G[2Z.P#D/O&^+OGUPO)WR5M<;1U9E]YOAKMALHVSf=5E7CE(J\-,XUZY
H80#<f&WK9]J04;3Va_d(6V6:eVd1DP]-eJ0NW^^+I06V3+==O8\B.,b#_a<JFLM
1PJ#bJOJ#QP:V)<e46^)Y@N8U?7CJAHV2ecH@,)@[HCgGLGW#F)K34G>-&K_9[Mc
HYJ.96c](OEX2Gd_N):_?@OJ3aROe@4&:QODBefVZS,@?XCb;+-\HZV&&^A:+(CH
N)N3GY?[7A[M,+WH3I^A71H.^Y-ST:BI-fcXIDA1G)B)0BK>&YfU@C@?_3f<CK-E
S,e^Yd.@];ce9P##R?6ZY7Y7PU[NFd.X]M[&Ye@I&7g>fVDcEDCH48eIH^.+/0#P
^^EW?bK9[3&S9F5RdV2Pc+&K:L=>54gMM8M^X7=a43&XWL<L:0#5/T&e_-<#@<\&
3N3(Va:bSJ4bR;X=ba?+6W@]C_Z8ZTH7g/;aEE,aPQFeUbT<Q@MDOPP(A0@[HF,&
.#A]R&5@eb/T.-ZHd#aC,CF2QTX/>EPCOPa7VH63^ZE)M?faFDcZ;1O\&g;=\)c^
FEfD>QL;?T0UYC/LSM7aACPA]UGXNOEF@1X)^]-;&G5)Aa-75b\,5gEP6YM6GK@Z
1AC(B5UaN[>;>1@4C=)Z8H<?Y>.^WT+^fHdAH>cIM2f\T[cPf/DIQE@I6)F7Qe.W
6ad1TCUN;W/Y;eU,^):>92?7R##-g3NSN4DeDd,b6QDQ]5VE&M<[23V9TBCQggN/
I=V:D,)><a1>R=JA&(JK&(-)fLeAcG@Dg\L&Sg#\_2LL6#M/JB?=6))A0).T^79^
/;;G(LNUAT=CSa>>:DCg.YOCbR(WJGgL+,_S,A_09R.bgf,6VbbYMLIP?:1C5ZKM
:aO79L:I?&8MQ9A=2)4&3[>7Q=G#K>bJ-XDL^\+E6Y3K#S?>-RI2ULBQ?5L9\NC/
QY&4?#6_PXN^NW>;06]:E5\#[S71\&=S])[MC&KFM/(;HDPUPM9b#+G)4_U8/7(f
.He5fcD2a0SgO(0Jf>70L@9Y7Ob11?dRF3bV)YMN_]bR\^Kc;Pf_:=VY&Nc&[?\&
Xe65Z/MBLM[&YA5g0cP>7>a+GL[^dbHC<3NK_c:fa2T;TF.:]G?e8#@eBHc0KUNN
bZ7)0)L87;5[dCa&0PD#b<3cAWO6Gg>C_2/@]H6,F8>Q:(R1g,daWL^VCLYL+B^<
09W2]aDQ@0\af^.Yca:+G_)Xg</8/EA;7=M^#EO5>I[9B-MeQ1=UbedXA3gfKM,P
^RV0^#2aEb\12_43F\,N4J.2[@R/6]7\OT_R9N\YEcA&7ME@E#Ga<7M1>1GJZ=<0
Q->d]6#V^W5df@f#TQ1824gUZ8WON.69HY4X=TE@T)^(;<KYbXTN23ZV9X5V/;2L
f:YB+@]0UQ/Z_e^LC^=+9#?KW0C+D]Q5=PSb[Hf,PLHU#-\VaRZM,K:\:R\#9bf2
8D+e3+=M?d[LUCS&-RT=+N;.,)_QeEL4K6.Z+2=05;LF4P6@(8#JJQ<>D&]Ma@KC
ZUT&Z[9[BT_G=B3+>PRQf^1<2b5EPQ1OU63gOTY&K:.]#05?Fb[dOCc=&A6JN=5]
<0?_N^1Y1.BZ)g7PJTP8/SXD2J+,Kc.S/P6[ORZgN7S#=]UCe\4OD/LR(6BQYSa3
?Q+#(TC]D1N-cKM?g+2[ge6Ub;.\8\g[]f3V0LX\K@[3XG7gXTY<&M]NFg/e>2X_
_1DQJSMH(Db.@44@IcBf)F#&,>GW6EQb;_5&53YXNa0JdH?8cWT@;R0E^=HN#_4g
M;:3Q+f+?T<-TT>;G(,BWb\8a:D<39HY(U=A0eeE]MfeX]fG-gZF/V2&+Qf,0YG;
<3g5AZZgd50e2/]c_<.a,[N6EK]GKD4.Z]612KIS?Nb/?VQa\c#]U4OZa2JH2D7P
111@G7ZQ3^/W=VU;IM;8f8M]J;I@4>>J@<P(>T9ENX85WL>TX7\@2SYGNW==YaD<
-(bbV>XWO5WO+3CDBB[?;bO?OI-3K4Rg);0_>92&Y,e8fE^H?a,T429Ve(7]/2(E
PYLH)DA\#R)GO+.f<VYdB=&:KbT/c3cM75V[LO/O-]60ScKd<NIL-C[<0#_TD1BB
AGcUM@8?OJGdARgFR:3J(:U8XR=Vc0B1>#]9NL3M,=LO12+U\WHYCUMB[]R5?=:;
M0N9XTI_gJ9DTMK6QQ0L=/-69_W3YF+,gYN<V=/]VYgc\AN\C0U\R(a7X=Rf>DJQ
bGI;b=SBO8L:0K,U;dG=d-9P3+^bURb0[CHfWg>2LT226J-d0P^F_+O=/@DUN=g3
<Fg)B()aVD@00&][R<]cFTA@X,;AfV=BUOa&a\#40I1FbOGH3+D)JC?K_HF<8U.>
F,9#:&G-J9M5);^b0[,:RS_S=CVa?\+8V-32#K1M4:aVM4_g24K?S#b#T^80_WGS
3CH8KXPQ?.dMXXBDadVIFZcd@S>#GG\_P:b</Y9d=GC+UZORCc&fc+faX9.eZBOG
b7.7Fa_6AbF2(K.(9Aa(2E6#YV8PA)&0_04cATfSf@)@(e<)INE]QUTTSY)<Nb5a
9Sdf<LKK/PA/:-Y]W0:bZdHf:V:,1U_:ZSe2dGNHaf@8bM@O.&;P<\WHA^,NVVS<
F,4dZ,a2bTCUEc,L,OV6dZ/;2-98+\+Z6_GT<<BKBOI]_M@<6faW)0,YdURf3^9B
M/;fQ&8T>\6;DTcF]dV:EedaUeJX;+E>TAQ+DWIIU1R,g0YBOg2NBL5IVR=P\+@2
.?(;938A^Ie)1C;QdM3N+)f@.VPgY0<V(D(5/6F>G7_V11ON2.:-&I1XMT(Oc6>V
+;?eaTTb)B-50+U9:FW_1A?a8aZ8D,Td?8L<J=G]gW[#b55#eO7:>d\39eIR-=CT
>CU&]^&V)4BEc))+1#<J,]Y^eBHX+&VZ=7)=RN>-@6Ve84-;=H<H@&f;YIVAIDL)
I_XWE(;.F)^F9@c\M\QW^XJQ,OVM()3.(+AH>_HS35[_>21M1/DaOeWKDJOb,J4b
4[WC6R\SfGCS]V[VF-2LM5:Y4,Z5c?3(_LdN+Z.3?(=^]c7cYL;WE0+@QDI;cf=C
2@U9ZgAAAgFP/XHUG[22H[ec.K0g:Z4QgWY:YFJV&fAYbR>E9\Pd9ECb9N;1c6</
W7AF8=-^J_YI:S.TU+&QX[CAZ^T2b[//BE2g)F/W464N&FbP2-gAMH+cYU8@W+GZ
2gO6BUBa;VV4EMPf=D:f22VM[,@,DNMAK6d+1>#N+1/fB(&K3X(8L(1A@PLF[MaL
fN0)@3XFIAf]4A+0@MYL:9_f@?W@I1+OI8G7W@X:M-MdaTGSFNH55@A<75X/87eM
T2F)0]>=TL,1>,BU],7N79Yg2eO;.OWb3?57SEW(Dd/QFSMZb4YX6,WU42:4B=(@
c<W1?>=@Td]4;d;193.e,D6Q8E_YY[1-g6bDD8>:a8\7QU,DG/9N+e#XbV)WC\N2
g.e<g>fb41DIN-U/(f_YgS3M]Tg0RPYT5BQ6O61A>^65X_OS_c8\I53.2GCQVM.K
a9^KS1e6W7JAU1OVHOa+E9,=71bP:NKPJ8=)TdB;5e;g[I/PRT820&3MGAP\cOLB
Z?J^O>>aL1N7Oa-VQ>..GI,Dec3KGa<P>6<C4Cf58B--C3DT#HZD2c)_TEfV__=&
ACU&RBPRY]f/4,\^#dQc<:LT_=YXYg3]@@DRM?5HH+^@<X,>K:DE949@+R>:T.EC
g.ENSH.=A=V7V(([MbI,VM@:C/aAY4:1+A<[-JXedSeLgLL3XPGCF63<//X?a0c:
8abCMPA4,2[F;=gH/_H;N0bGN\aQ>;C1e&7.Ja2T#5FGSb0FYN0Ad-Q7YYgacZ8N
@T74>>=dU+[FQ>5K/cb>>/23@;cBW9&U:fX^S1B>OA[(QJ#K=\;F1Ya4I+(T31Jf
5[NF?H2>C&-eBdP39@A?@N>FYD20Z,R\/WSJSR?;,?P\WWDD@M1<R(A,.Q2bLSa<
<1f8VUb5#b7I[:F<4+,-#E+K//#Y>f[#PPd0/.BY#H?P;Zf+)2@_aBC8),HP=V/f
>8Hf^Zc+,2^A(-CafLT0COPQNA6VLFOObVA5\IZW5NAY<29#G1AFb41>/>KgLWdQ
)\E_cf[4B,AB[16&g,f^1K4+([Je,c:?/#7.b\_J3CYARKXYaOf.#M[(66:CL\L?
S0U=c.+Z60aL@cADZIa;;a=^PH))2Gg+YSH[T_PM)a\)G<J[J)MXTF=\a;TF#R1]
)O+9A7M0a/7:H1^0.Caa4D1SX-ADMb/\PEV602CN[>0,Q5,dF0PC+DVO:\3>E(7#
9/7(_[P096@Y=5W2XW7\?g0FS_Q\;7FS^=bDb^=X/M7(I3?^TRS-:I85=AK_26II
H0Y8X3,?HNA6#NC>C\<N,LREJ[1L3bB]S:R?3NFKOEQ.BIE7XG3gb@[K35-4Q[B(
/#-,[@,^4MV^.AOEV?eK#(,5]R<3E>80L2\E[9[g^.ZSbSKfLIP2OOBM#Qc:=CVN
P^^<H[)HAG9/M-bc/b)JMEL)7NA5Wb_)#\#74H3TUD<C7ID9PNfZSefIT7<c=E64
W.]SJEVHd+S)F(RS:f]0[S=^JJ_[QLZe_Q)6PDf2KAJ,A9V])<HQe0&BIOFaXM[:
QTE:KHgUZA6?:XFFIKIYcbTWUB#]9)_1;@W8R[I/Z5@:[Nf;fYb+d7g])+^/<7.1
(07Ce1.U^@I0Y>LdcGKBSUBJB)))@4NNNcgFM/TYDgY+T970dRca8(8F=79VZK.f
Z^B/(>A.Y^7[M([Z0^D)/58SC_V0<-R0&aJ.^bXK03=&9;BF82)).9X+_SW_6F^c
Wf:<R52Zd5MV[)I5@fO6<#a[6aH[AV;T1d-fHHQNCfPMER&0@_9P22R@eVN8ILaB
=@VSKe3;X:0NH3RCS1;NO@[Q<]7:3/AS17&HD_eLfK)OVdAJd)^7)<AJ0-B=E)UL
EZ)RSDNGVWYcN(;^a.+)VWfa9MadP]Eb:]IeK9+D3C;0I_(ZQOF]3EQ#?^,((N7Y
[+5N#,)J&S\;;BR+JP<OS3/P:6EdQa/MP(]R7_g\C-)1?QdV;75U)7VIFPYUe1CB
XDS(a5?AdELea8=-8g+U5)W+E60?N>D=8)-d[/<>fAH;WWg7BUggb6SMgTM:>e@=
B&F<<g\(aNgK]@>fHE3[(MZaG/[>:.QT1)0HDLQY[FZ<WfbTWX^6/QQ#D)acJ?>K
NEM>IA/Z)-4NI>-2C<\E5VVL1g^@7CI2KY3M^4,X-cXHa:SYX4?[4:Bg4#/^(Y:J
&Q+8dPCe-=aAV)U,G-]CeIcDXV#40PfB5[YA<eD(D7T84/(O-C;R4[Ig(CH2O5#X
GM4&0_)2--</3@FO&WZDTb#+E,a5GEHB18#)8OS._f-\#=/d@[V+#O_#+4P<RU?e
8GFKUCFb+G#H>R,,dNaN>PfKQAaSRX1ZU1ZG+RdO^e@#4V,R[_Y#d>5WT#?.8=)M
aZ<P<>5H^_f=L8B&f:)#==YID3)^b)dfE?#@D?8B)AESfc6.,&aJ8LC9-_G:+W<B
&:YOMg4_bN.76LYGLF^=O<>O1U0?=2F8.@Z[Ye)]GMYC\KIL7T)C]945_Xc126KQ
FR=(1?A#4N0(+fb7]gU0Sc6C4<>;9D<(ba8JC2.(aQK8RLI&@MQD<_XZ0R016031
(T,a1d^2(?AQ@K)YUYYHFO/\=3>[F<B?BLQ[b;T;c-<)(BK\>?62ZC+TK(OJN+08
_:@CX76#&C@R;KEbZ>B\3&42AZEH5+H5NBEd,eQ7;T66[T_6.DKJI>1\[MJ:]Od?
+N7QNR?N@>=4^d0ML\YA:AO5[dP926K;W@\;<)[NO0(JO8fN>5SU?4OZ4@Y4N7))
PNX3HFWVGTKXf3U\V;(3^MEZ&,TZf/VG.21gVL5W\:29@b)8:Y9,a2X87SM#<>80
#<XWIP)^LF_Z8c(AKG-95A/W0^G1=PDN780CN7c:>,)P3a(5OJX()?KCCSR0c@S0
)Ne^<5.^G]&dWSPU):\N+--aXJ_APbPZW18D9>JJTIdg/268IfXQI\A5=&@U7B6E
V/f3WI3:Ed+#F)AHgFb+3TN1HGcPU0/=JLB]9AJ&A2fKJ-e?4RBcD4TYM:J0YD2V
)D8M)7/G@)5:)d];8ZHSK8[f7#f^FLO>.(/Xg<D6,RaEWD1]Na\AMb+CBcIE-:aL
]1C-NW)=AA02D>A83&H<D?F)H6ERX0aVGDdUT0JK8/73&Ue39LXZFLS_KO<+.SA9
6B&GIUJ\OPQYd#ABS;^,)Da;GQ)eOGKVN6?A+R0FYde,G4^O/>7=(WKJ1/.)eeO8
(BJI59E-c3TA;\4(./)cR1(L]8Y)#dXdC^?Y/CFdHLQ+TJ<9?;cRQL7g&+&eMX9<
.GRbK8:O^YHBMG:-_-dBM_GMba/MT(.ZK1GV.7>+f@]e[Cd1C9>68DKFWd<KV(ET
XV=IFRY>0AL6OB5,gL\dACPZF;^N=59[GHFa01-BE>;<N94gT&\QL;D(C3bP3BY1
ZddQ/2,,F//P#J2E9Xb4e<HDgTH3;b=UA>#.gDf+?e([R6X.EV&2:b?0cLbA4BDI
YFJEDPeQ,4TeL&/;R-+M)TXdSfbaREJ.-CHf]]SF,,)J#J5)P&=bI4QE06;:[K\A
TKSV-:::QMHe6>M>>]\2/]&^DdafSRF;8<;N[D:D,L(;@c[Y4P&ePN\\I-)RW7-<
HZPI?dEE)/B/2Bc8g+L8?Tcc#gNF=A&@^&MDES&O6:89R5_ee+//Y?Uc#=f&Q)/G
THJ9GXV]8BKAY(HGNJ2\,.(HG&D5efJC3)HC<R@^GIQ6BO63BQ84\91&e/9CPPe,
?TTWe(7f?CPReZ9O>##OKWd43dYf@/>T0OJ#?933?J=JdM-e(8PQBXdYe<(P^.7^
D2S-?KCT44SEK#__aRc0-JAFY)DY>[N;UK.9N(-1M,W.66,=6D)UgX80(L_NRZb;
N(GG1cA2[e?cQLOEU9&7(33eGd3I3fXWT>HP\>dQC1?4RgIcI(5RQHE+\&cVe4g[
]^JdD?Te+^d_I,Z6+IG.UY-CG^BOH/R:&_BV5:9bd;&UPKT-bI9O0A9Ba2Ea37\S
1K7<ICT/ba]RQDIfXGM56+#?e9DM&,J;MH_fN_13XTE0;Y[(_G4D=VZeGZHaT,dA
I.:X02?\410f@WKMUfLBaBP^9L[JG>R7Q,cZ@COR1De+aWa;,#bG3d/Ue4ebbJ?W
9M7\>,(VV,FBQE#[L/\aAKKPX?2IYcMQF1N58<SCM1=M3YPBe9@],CDQ^.QBX^[A
&\f;]BVMUK.IF#6ZS3OG]OA5G\DNg#]Hf0OS5#f8LHdT,7AKag8OK;J7U44)aLH0
bCUAS&X-<a9_>?)6H;<C6P_O9NJeYY>F_)T(5Yb#&..:d,7bJJ)T)^eZFPS/LD7.
(LVB^3Oe41f,L0/T\8RF,]WIX,-BX?5RV04YE-VRX?;AZB9_NST\1c;V74FZ,gJW
>-T9>7+QbJg?F@IQKLO4#G<0?MDEGVZ&73+:bO6fW1^3=D>DJ;#APUg.cT9FUYW3
3]->?]6]W=82#f\Jf\T8fA\(g>2CPdJF^W\0QSYdDdM2gODg;\RD&YG_]N2J8@G2
dW9==_VPbU<]4,K^N4d.a/VCIf.R;cQNDIc7\g0P+WZe/5)g.X9?A;O17(&Uc=,Q
DaGKM.3F=Wc>::HGgAeZM=5KEJ)BK(Ia,C;LAc.D.25Eb<_D6fR(8PL&5[#[3SWS
,V4(c#9M_I?W90]OP9L8Q:#]A_RD5GdCg=1/7RBUYe=5d.OKQL5STe5[ceHMe^65
D42U?@1gXb#@c9@89H3]Le5-&5KfCI+4]O@;MU0J11NZPAc-gEd8:ZKYE3,C936Q
PM&HB2(-)deOf@)ZL;fSg)AbU7YE[^Od(f18-:W+:D:IZR5]5^\]-,PQ0ZB+0DC1
Nc-9=U4bCGY\gWCPF1)#)2=&<]2A.:RFc&Gb[VXU+]UcMBb:[CIH/V1U:I=gFZDG
_D>C=UM_Y35\dSWeV#CHL+CNbE+BFcfA5d3DTcf<F\S,5HDd+1@A1,FI9@1=[P:O
SF<c^QXX-<?,V;fN8C>.RF,QLGeef-+Aa.9:GB.CPb]5;>0J&gO<(R@BbT/Sg6_K
(+1OB5HYRN84;#;dN:O>S8Q=3b[V6GYX8;E?ReR/5\(e5/W7KeS2O@T,,)d@IK8R
2f.9&5Ya,e,#)-CKL(aMggU;89J#WdWG3=2FgTN7YBP80NBOLPXc>M,_A6W0+2Z6
>_DGb]Z9_N(<BX3dL-IQ-H=^Y?<OX^aV+fB>OXN?@e[:1A_,;R:(I_.+5Cd,:4_<
NP2#0Ed_#H^KKYSPdSFF6>b&J<K,L2R_-YgK_GO/ZQ;<.2I?S^;U[C]#YC7W5S3U
B)<0S,4EHb3R3I7KVN6d7Uf+dC[ca^P&Fb[E_I,eHfNfFU/b@TaEN>/-?Y+agf=#
Zd[:ZDP(U68fG9dS]2E3CG#XbYM1(?[<AH#c]c1DU);.O(,_M?S1:#/5?Z/.]6/W
P7#R<JaW@2(TU<]P@PGNS:@P15S/9(MBR-b,B/F6KZVI@J)PYafL(288AM[<<:/(
_\4^4XK.U;P+MC8W[dV_;24UB<>f9BRH=4N1WHaZTM@Lf97A\@.-c(Ugd<=0.P9e
4aPDUQg(\dMYBCG:E2N9X(dL-W[[/3ZK[Y/FSgLRT^Df#TPG:;]K<d\+19I/PD47
E,:4CcObVd6>U8c9>>GCfgT(J+N.CCEg]>1EbQGO)GJS7?=Mb;PgNUN.GfG1_(TZ
aPYI5PGEHUHA,YD>ZR,H:=<F7(\bY+HS#XL&A-bC-@)6WbZ0(+#-4I@L/=4e]8A<
.,CO@2/Y2T^6B#d&0aF=<22C_g2&#4DW,8;+[HJYc6:F7K+>201&\6=effgWRC/f
QE50be.^EVI;XUaY952D<7B[aCB7[Od;>.TY+JeV6a]&1XWZ1INg55IO4e>e=5KP
b;&G]CD0^&)TOOP\U,Ug_3N/LSf@#B?ADPaQfU^#@Y^DLUC?BGIdTZM_IW&BBT_c
<-gY:d;)Vc]?Af<dN,)?I/=Y43YGaIEfTO2&=42+9:-Z#(07PG0_8@+69+H.MRU&
M;:T+,PL9@7K+G_2&c)1#7e@=T48.:DR8:(7>+XXg12H(ZKMAP[]CD1d[b-_)]1R
[f>N1ZPf[]D4S/8aES5F4KEe9E0ZgWAPc1QT>0D\4I.#TcC,DY-9,AW4^5;;fP0E
V]C:CRMU:0HUY,1bU+VI+cDOdc1)GSP2Bfc7P?L+#.,edE4KYe&D7^TI8?<:CSI:
Le<VA-JCC3UO.5,B\^GSNQOO:L/>\Df2a=)XO)#1\ZOYd>I-)-42A]:3(D3@S+Y7
(&YU3_+4F#71DW74]2:F3],cU(e)U(),F.I7PJ?KOB]X<6c+<VN92RN+?7B;Q@7-
gNY_TbW[ge,O<6,\UUcRU)BGI/,JOcVQAQ+)a4cEJ(BHbXbdDGaX-1=Qe2+K9J.9
9VGbHEb<-#05\?&HXdV#=L;Iaa;_01eRUf5#/G37c[MO[?1S3_#F/#a#fFN44@Q.
32#Y-ESNK_PS,EBad=+g4)G<H/C-U50.3=K.HQ<a+KB3>;3Q;<aeTDU8fJ1YSg>V
,MEAMQ-_4_+69(M&V:V=N1@db/J2R/R&UJ^6d7(F#=/[&RD]1Cf3H(FcMRE)X2M0
2Xf,@;3)<.(H]K_4T+^^g=V\a5T-Te6H2?1bU07c_1HbVPd,A;^>+I[OK^SV6_TV
U?L_0+U51:]RScF1Ub,dIFR#3BNQb=c;=c7@#X\M,:ZJ+JLf38[L\HR)_U]XCOWA
JCYMe4d0>UA:cg6W4N(B(7R-;>_,gLT5@3/6e\aY5C(N+YI<P]WU0/I743.Y<[WU
7c/=M4VE4:BbXa-+Q<T)dCJ^Z(Q@.gZU_;6JAEaVXCE]0S+DeA/-M+_KXdd8+@[Z
AD(;CFf3)#K_REKK+bXXNVP<6_2I(dgW;SdQF1b#K6bBf(ETWY@dP#CZ#J,^)Y&H
Gd2SLEGX0VGJP1QA)X<AaKS^F6-,O:^B36:M_L6c0gOAXIX\&VOQXURK\<b1DQg+
\?6f/+VQ6)LP=]YE35g=V25G5OJcF4ZZ[+gVR28JcISb9b^GaJR26ZRC3V9@f^G(
TF3T1E4I>A9e#gAN6_R-3[,26dE;-\UdQA#5>gA[3TdH\,UHXeE7aK#CaEW:8^]H
_:=GU?>_E\2bFV3#\;C0.AaN)WQd4[g]A(8g&HZPZ:eR0O;;fC:Fb?b/MWL_4-F/
3I):aWW;?B_IZ=XQQ2[Rc/Z<L=[OT4BE6[GV]5JY9HZQ>SDeNF>SXI).1^Y2adUI
M\F/OYDNR7H7[KG8N22/Db/S&Z0TWdW-M:#QaBROO#^JR3IVP+2H-]ET+XLO@UB&
:T6+1;:M@LYSW;WKB8N&b2KaU8_/67)&aY]7VPg,AdP:e&)Q+E)9&X(=/&.?>Y#Z
gdaI+1L)#2G[&Y3Q>KN3g#KHf#b0BIAKEX[H/RE?@)#0gg]G2DZf4=LE&WYPdd,G
ggAHXIHK7,67dP6:7ggM+>0KD+;:;T4^)/.43Q^>R&?7-ZU4^]0<2RA@FF#V\]^D
^J8g4f5e=Re-5c9&1P\+&5U=V5PJ..Z\;ZcT5.EL/I#5cF(aUBPRBLO+S.E_+)[#
88fbT+WgULAZb;c:NE&Z[2,=I-^.BC-2@G-:.T)gZ5aLN5EOUTe?@BNFA#;Jd9)?
6(0a)AE-MIX&e[R/#A#Q5WJa8Ygf)]J^TIC.6ZM(ROgeUIXUQ^/0X[<bbO=H_EA:
1X<>6\L5[1?_>6+I1\[]GX2E,HWE+1[_Na]IPINL:TH]YDV_EK\404/#bYNGF;.>
J7/^a,cTUV#3(B,8HKc?RG]G.OJ_bHNXLNX1#7f^0H5gMPB(QVe;fBS@H,YN[+1[
bDgadC-GF=#aYSe<_(C>EX8.BI:O/[8#)0=O5?C7Rg0U43V&9MYFS0D3Y:.AXJMD
?XJ3R@]M#=C@Q1^^?)>bZE)UGRcgaUd1##T=Y\ed4?gdP_H9A^5AeZb>AS>R9)6N
ed:Re^\Y+2X:M+)VJ3eegQ/aTW;8d)ZW1]N#?&?P\PID/00GR\T@Cd0IAe?XF0MA
-NeV0=@XVR0IKg,R5MIIP?L,g?]=4PV5M,?#5]eM;ZNMSE/.e,8@9M.(-#7dNS/J
<[F)WRGQ-+#[AMW]^5_HA/B_VaNB^#=D#Bg&^T0V8?g^VVbEgAOG];#TR.3M<]5?
Na+:(:Kcg?+cUg#)+;07BgG&OKb343/HC>BePB]#]3,1B<5]<U_JQ@(.R?PMP1G_
?T=-Y[<@]WE-#EK=;7-:#NHe1ZD9f\BZ?IW/&XJ7bRFFR_R\6MU/.N4.MX:7+/C@
<A6@@/UL[6La=:L^6??2>;51C#Ue]gEaR9_)?)0T+_#MeDUCg-HB2Je<N3[M=)]X
Pdd#c6cWfdd,[VTL;Z&<)@0>dBgA1]MTQJKgGUTF+:>+.)9b:FMNF(E^B?-O@GUH
/;.OQd[Y<+,^&NDX:6[)(-IQ92+_&X[<PdGK&fDC;WZ106^AC-44U,?:.K&(DZYa
]Z2cUY]#21YaQ+8X;.0XB6:T.^dNc@ed:7@H1LLdfPCCHSc6T96Z2=&>HI8SU&RS
IS(;#\eQ4)#PP3]=?9bKF.BV^f24?f..c<fGII<T.CSPX.QJN<FS[P/GgAbgT:c?
RW;;b9;ZN=Z#8+BDA@b;DC/&a6cUcEK1F0ZJc9TeNC<<73,:T1C3NeMZ1>T>0a#G
]9c]+.VD5VdLNT<WIOWZcU,XYSGC-S>PF/gCg1Y)ZHI4O@XaU]+TJf?ge48SVb@C
L>)48:\.F.WN^_Qb+P(?=a<F9C=N<_KGG_)XT<4Fg\^KJF)5EMPTL::&&c7US,&N
f4f1^U1>R5Ne8KCd]M9]Q)VLA;dI:fIG00&R&Y/U<+D[L=SJG\W_PUB#1<FO#aV3
J_^3]H\Q^0@8?2N(5,\3Aa5e14O8XT<;)9DD2P;:TVGKT:)XDOC3X\5XEEH-#>\:
=-@JD<5\K<\RPTJ0<L+&]<2(2TDGGcD04MM]EE56EfINGGPM[1&H+0A)HC9+_@E?
(-EM3)AW;8YcN]d+2ZG&S]S?0-VZCJ#bQM9/_WMF=C5g5)C80E0_Q>(N:LA./:T-
B&=5R,,31DP^U@)CY5>K4N343UWdB.,\KVJR,Kc\\H<CE2XcHNeWBg@_08I1)J=g
59AJ6O[./dMP(YC(gVKb[4R#GM+TWe+;B2IC;G@IXOBHMI/5f(bLV.H0?eeJ1V-B
JaEKSIN8C#CM-O;>PZ5UO^R39=<9ad<,L);PNF#9^d/T>_@eL:O::[NREHg(31T9
HUK;Df,CI3KT[FESeH(T/0JJ?IeQ4F<.0#>82-fF\QB9Ab#&H-?N^?]@#AB86,UQ
\X1Hg7=YHfD+#X+>3PAX+S(FH5XQ)&3XD85=b02V)1PD.LX+<>_Vb]>5<ME3K@ED
I?354bP[E^3@B]YNS0/gNE5=0P=7>-5>-C-\<9#HfAQL@\).NFZ<@7K+XES@^<,a
\e&&-CBVM&<0AEP-,(ab&8_[\3aEQPD4E6eV;9:JRX6<C,SRJ3-K@=B<3G_C?0MM
N2;J?eBQC(a<1G_2NF)W01TR_IXA,848>(S]P9LB+CB<MGHU&]9RQSC+Uc#-fPc:
Cg.W4ORCYgW:T3&:5g/DM)8H.Qa]-X6D&W;>\G.>Xb]P7J>A:,NH:dWbZT/]VU>J
DaN67QO9@;dJU7,1Y05Q6ReVE&:g8==U7JLL-NDI\I2::+TI@f8#QD3D/3@<YXXO
J5+QU3^@_dDG(+.@21#WKdbf,^JIQ],JN[:R(O)/TK5A.AdXbVcQdX\R+M\2_NF\
4<F-L@674YcX3gBQ3L-U1c>DY&V/.b;dBSQ6]\KSAV66T7.B9HB<+a>;W6W>4>f_
Q4#[gW\(X6#5UF/C@&Z0,b7V0W?6&J+=(TbgI.&C?_[>3B)37aG.1),_KaBPNST.
fbJC9V+#YId><&A^996c)9-BT^#/?</-XG0RMG6K232dAWK87#VH#H9^E3(ea5F/
>==Zf<,N[<&AL/Mcea,N:OO14<f)0PZfS-CPDW]REH5LS@9>cMKG^>a:_=LMca1R
?)3:eG4WL6_:RX.Q+2=^OHM5Y1&S2+N6,H0ebe-A>CCA&;-LR:^G@0f@\=ZW2?Qe
.=)^#_AS>==8<BD5EKYfKf3b7_U@HMQ/:HaWLGEd/JE?&+IAb@3.Y)(cfW9b^?F&
2=1DfS3+P38X451C-[4P72]XJ01KB(<gQ-QHZV.Q^#J26.G2FH>@.9<WQS98b/5_
#K/.Q-&\DG@JC]#;<_^ON1:Ad:O4UAM[MM2.ZZ22R<e#)M<H1&GHfB6C.Y(TIc3J
HPdR@H3]3@<D[^(=KJ-D).X\_H\:K,)3N-W#4Q+&baLY0DOZ5J-9>e@ca;3YPD)b
[-<7\R2;./M\R?P30T,@M53,Tb)LXY_A,^U-Z7:E<+8.]V5MK@ddCY@5#bJKbb&Y
W8]/A.Z;a.Fd+4HZMTZOG+;IH_gMP2+O@OP.Z@]bDS_eJf3:dPLJ4UEEFHTg?5dD
J+P-LR+VBcHW5<HO42Y?9/G9_->G-;gG^VC]^)(D(:GSO@c4c]MXY43O@/LCWAG&
cWHJPHT3(5-TB#)Sf[TE[S/C]IP].A\DXT7L8f]E8Tf&8V4=NH_IU6?\.I;gbeMY
YIQZ,6H3^,>U3g(ZJPM-WX23:,&VG4,9K68INE&8L-1Y]7EI,GX8MF+Z8_I>D5-J
6Pa57RbTFBGc@=bWc:JAVbCbKQZ=.=DL0>Ga+3XSD+-5e[JHI+^eB)aF814=NB-.
[(gT<Ca20K74D=dL&RI/.MGAMe6C2\@6&>@3b6Y#XDQ7V?C^#0)81#U4.Y^7>L/L
OYeFZ[b8C2+>M,6L13][ZgQZ(2,cN]?5ACK.cJ4;S\#YHX;TXS=]C8.JWL(;B(bK
\SdUEJ8ZeX;Y>Zb/Q6a3Z48W2&KUC@2UCfeMQecMf9WA@S.M-d(6,fd:+FZDN\1=
(WF3VZAM[-,\;Q_:Gf9c5[&Mb;,YcE=F\4\6?/S&_d2V^OcI9de7/J(.(O6S.9Mg
8BbY,;OZS^W#>R:d<ERX=e57XgIdga\6V+eUMZ1<W^S?O/&ZOe(2;17Z\I,H/PD0
0R6:LU7.&7)M^3(,-JSgdN:BOV2/4UHCV@?K&RQ:I+LAbW]/_6&2ba1(D:-WX(/J
9Z[[L6YY^<;6JK?3_OITEDG[b;6<0?IUfS;#3IJRf(KP13LHJ=5X?e3ZV:F:N7W8
7LK]C2;2P;c@)R^RY/NX\3#2^0X++]dSX35R,;C^A@VZ.=(G-fe<XZ-.ATMTE6@e
)gJ&H7:\A10A9gU>a?H9QKfgRHBHVMFKLWa]8ZY9d[g:c(1K[^S)a\b@#fP?:XHM
>1H3ZA.]W1-;(BY8.FWb)E[FaM]5HG;SgCR2eUX(a5QT/_FE<,O;^ZQ2N0.9+.TD
1(O6VYHD-@+:&ObFKLe\SQQQL[gL,/]ZG4YN2+gLA/AR8(d9a8QfI25MSd&.HbW2
X1.0=<6+8(Ec60M.^(8T64./]b?;UB9D)I==3Q-^C#.B,d(^LIFV,SN+T)FN<FPU
=O.8E^S#KNVf>X]c]SL1V6G&B@@cOSGYC(FbESH&8:>J/eOFSaEF4+A3JT-6=>9U
0F_LddG=_:Z7EZA#VMU,APZ]M.d4[AN17T+d8\TQQeH(VA@ESEBIB3P]7^2J?T0g
Rc?3/]43g^K7;W_<g)Y&N?<2ALZ;++3:BUDaW7U3;#EXbVNcIPefGe,bIPW[(VND
;DPXT)0_Tf?5QE_DH0DTa]MK_bZ9ZT_;8e^S)ed+)EU@V1,Q5Xf,<]C]Ie7A;?T?
b:TX-?8F90[P>L4dR_]T.GJ64O5P#.GZ3-+b4:B.--.?1.:R.cba:M1/5)fgXL+D
P2g#3FDQ:;;[/CS5d61:,]4U6F\V,8+H-cd^[Q[<^K>Q5Odb46J4.?XAYKS@d:;A
4+3-.,/X8HZ62GI_.<K65)\I0E=XQ9(1@X-1bb>U6&?g).#TVN9>FFT+G<)J:V2\
OJJ5ce#AB];bERV6e&bS&ST#6EU\&2LFXA38d_0A6_e:<?=U3e8?fg(UX2NG)UK^
L)Z4=&F286BX)5R(;BIW7GPEI&\\Zf>fD&f+b<GV(?;>0UFUTLWE)Z[eeZ,&5c2W
cK<ce;L,1T#\CJ;eCI]R]9Ud_:T(T<&E7VQOE]a>#;L>A::=fPA2T(0]G\Zg#A>+
^0XN>>,(6+7gT2I7TdNgY2,ZH&]YS\8-_(/gUF#7fJdL?WQd3#=3;7F+M(Y7::HV
/F;U5C6S<[D/0g^4RIAe5>Ra>HL&C;0(M?,3NR>.774Nc#+B7XV9D<VVEaGTY\fV
>XECUgH2a539HH^FW]d7>eOeZ&T^d2+[].7+5E/N7(VXR?5-()[./BLPUJIA@,bK
^G_O96SGMZ_MC2_#ZL:XN84MX1:(A0cf\?6_<NcHWab@4:BSYYC5Ec3W/M:,S@Z[
NaCYYfWC)G<>,H]>74\5R149(@K>7^U]\_D6;,-0e]PD?cB]O_LIM:(K/ORU,]@=
?:IcaG>P0aJF^V4G:XE\>RLW.9B@A8^I?,6WVU_Z^)g_E,[+V7YUG0V9B6,-UTEV
FK[Vf7aNNW<AB>S[.-EfKP4[BP;edHA&X+1)?cRVA=H:QR0;SF.-1N\FgC[&6bQC
2WJ0W_F7KXU8c^2)+?bC4:B2fa)F#)WN-.[Y(-VTX(6AZdW51]3[=,AdE>\N]<Rc
,:5Y/89[H3LPB0ZW,7Y<aReeG#FB9KQP]?SA7JHPQZ[3V-(=X)G[dF23aaI;KM]?
Y:V/][>C63WOA3V;97PR6+7&CVTCW]HV]8IVX[D9aD2RLdXeP+RCHZP1g7fYb3R[
3e>OagP]0Q)9,NMRE[JM;_L)?>d?M8=d1B#-4:eH@2O@RA7?4,H1N+6WecY3C7EI
d8_/<=:<>:Ie#H,/AeS6YI>Sa]:G2+fc-Cb01Y@<]AF\EXWf2Ude<F:SaMNZH#12
4X31DQ\X(A[MGXZ(.Cd,f-D68c6bYCc0f]:#f/0b2f@65A=3L47E;\f3ZQ+>4HUY
c\_/YT[ZD5.O7b@F80=Ba9G2(2Z.PQX?NA.CBSA8F13OB,;J2O4@W_&E.);X^MKB
8S1Y]6_?=:2e04HDZ4_2ES?#+f66W,Q]AWA[f&06;IcJO?2We;DGMcH7U+PBW&eP
#.@8UE5F[M32=TGOJ2>Pf2MV_N9+d?c;O[1EQ.#]Y877I(,VS8<C-V[.BHB:#7G)
]LQJZ6GAW-_f<)?aX0ZABF9SN7&<ILY]QT8./gDY]b.V8\bc(e+IF8^74VX.Df2(
\4Q>-_UG?Ad72\G:Me>9)FD0ONL]WdN]]?b8>^Q(]2dSJL4b4:b-1Y6Fd7IK4P7^
#>(e4,=(-I_MT?dQf+3AK]8^E-gc,\@255B>+#be7,[fbN3bC;1fFZYHc>ANbM9W
E2?9bX(d7QR;NP5WD5WVUOfJ^0<d7J:N#9[H^4ab/;W,IVVF/6.g\&N9,-Yb28A#
9Od&D?+KY2E>f?;(;+](6,E6G=VXBY;3<+Y26[S:0#[45.(=06c4bMZ@ADCT@Q(&
WXX?e],:V5[Ba8I.?>^^[0+fegaV1V2]e1069D:MK=Tb;OR,0XPX5HET0\FUL58+
OH</HD184DLW(V9-,7?AXGYQPODN=N:5V,0AI1LXPQIc4[MBAb3HR<DbIGU2bO:]
26=,gH][VcIQE:=:cdM=-TR70PEA#=fB:&D=30:Yd)3T\[U5]#Ag2#WBa_YNfF/b
_&dcIgY8O=X#M1V;Q(f6@D^K-Z@NbR,73NE(cZa@f,DbWY=:W^MDR(D<__\ZU5MD
)VfB[&+)W]d2H@N;Wf1D3JV0+2T)Q5<US:>G[^V5)21-SA:Te3EJ=:O,YPYeS,6G
GB(,A6T[NNLa#+GN)UP=46G4#[4CbFBgEVM.[]Z?;8597bMb/M3HNF6e?Cec+,9C
C&NS[)IPE\-/4I(U)Hb69S@Ub:SM4FQge,K\RAGS+<JL32?&J:>)&Z],fLT&,(K8
UE?F[UI1N0a0#KS9=bRRVH[^@_Q.aGIXFeQeaTEVSE1Y-#LO1-Od=g^N:;,d;+R&
#L7f)Z8-cf]N?^WSL-AAN5f373Zfg-?A\bOeQ1bGJC([cU]7]]EJ#,)?Lb7cMM]g
Z)54.DeHNCdJ7b.]U+#OI-TI8(+R=2KAZR76b4N2O,5B@e;JZ]#CP_M<60)cM^I:
_B-39(CQ2XWWEPFe03f;H7e_FZAdP4A&PXVO@_H,0,97MHB?__,&;VG+]SA4\ZE<
B.e6>4Q)LA&)X(35H)&GASY/T6:X3,SGQN/,&=VZ>[>^N)6RN8<ESfW[/c&bHV-#
LLH98)++1EU]BJ>Y?R49SFFdU<;B/X8ON73,_XOQ?HbMG7#0546A=_]LS&F=1e2,
Z_Pg=F>\@bX0)fO>?[WPc_WdYKgO\f_6?C2).\fGS@NS&f?WI\4>f^0g\6AUFgL]
4aM5(bc-e/U,(?5/\<=.G(a=V&\)Bb#;[R.>@]Y,^98W.X#;Y[d9=C,T##@4c>\B
HND;VTg&Lc0FdON3Xf@MLK[]25U&NO=PaKa]ggO4Yd-3)RcGW7D(M0Ie]QJdT^-4
B_58OH>eOMR(cO+WLcQU=_;/-=5-6Y</@-T1,6]=HYVR/9bP>ePd6GL+c@[B#g0S
c3-TDG:[@Zb#)XG[@?\#DWFFeW.0SAd?Z-@A?D,R-T&7.Z/b&PdGP;a/;EFfLA).
2OPY[;K:]1^_;B]cA1gOD48b@=Q0S,M:7.>;/KHB;Z2\c+8P_c?;ZgTA+fS6=8?d
a_=<UI36]7_)V26+e@7cP<=B4D0aGXQfKREJ395TC5#N1Yb?86D89(XXQ5&OZ>/F
M?]@E(3d_:;0H7cH]RG>,(D.LJ:MN/QH04b?RIce@#F?_2AN0QR10_1P^<b.8Uf8
S7RTKg(FHb2W:A-&HGL1dPFYKegG.>A]e05XN()<@F43d);CQ&(.?>PFO??L/MT6
@TK\<AIN;ENZ;S#\J9f[e<bS+)+5S\U?S71?#bOC<4.5XH0@gK0f.NF0NIY&g[A<
fcHZf0RNI4IBQNbUD5H1Wf+.4aDW#^T0<eA9:LZS[QSA@JRZMB_=+?)Q_432S3M+
OGDYM=,Z\HEM7D]27@>.M:\,[97\.4PbT.L=MJa9(PP-U;LCfS:^.KNC<]QC0b#B
(O+,9J=H_7OT=_T_1F3?aa1X>ZZDd5eFS&5MH^?9QNUA4CQc.2VOW9FAZ]/\CUF4
W/T/5Q>^YI1MY(ERH99SHTKY+c?a+?YZL>YdKJa)]A;#NG5KdLOW#A&+4gLK):8/
<aZ;gPZ5JJU&#d<+4O7+BbeB]F8>WV9-a,>(&c@P6?XGV8S;^X+Bff6>-DWC<R6[
I\f\]c0__D,XFP[F+K?87C1PcBfLbg-K;+]&^6I&?,A)>Ca6,c9C,f08^<XZACW3
OUWPD\L?deV)(.;ga&E\D?QCZ(9D:SJQ&&_.HY5bZ.4A)I_I(_QZ7fa-BO&B^13P
&eeg6MaA@_g:g/PE4fBDg#6=L<U0_5G;_C-?_IN,1\bWR4fWG5L.W?ZSHU8W]V;a
VQ)LS9I:@I@;R8gIeKABG1D&J[/Y32Db=.eC@7+(B.fQZe+^b=AP2@(D><X4c]=c
8#Da=6BZ.<26K(D\/d#\63LNBV@\<;.#Mf.7+-.Z9X/<?D?:Xd[1/f,=IL4IOZ=D
c+&.BH(C]AOD7b52#\#^AW76E>^[D^d(S3,<W/dD6DZ_9X7CCe2:K9cd;LW([VC7
d?7IFf9,LOQL[Z+60V_.cCc?A;:<\Y(IE_OSUIbb#9>R2^,@Ce<#MY+4bb1_]7RE
51TVZELHRaRS=SOa:#1@/Ab)@N_9VR;=Yb4I7\DAOP3T]aV]4GFG[9c[5(_:9CMD
G>\X5@]JTNE6_L:f1#.VX]-A@&gFY926BaC+/M7M]63=Z=)AeNXSUTa;?[eFW3Bc
F(HGDJE_c^E?Jc8IPe[I^g2RVd4EK&QR-)Q&S6<c6S>8X(F4J/f#T:IYF(cD8g=&
&[fT<Id]^S+[FSJ3^b:c+_8ITKLe#ZXH1O1dDQ_#aY&V(PRgPA2G6>15\E&ee>Tg
KXHD=XB(P]A;LPCA5:;=^,;(MMB2ZPQP[1C-AWd]&@SAUd]2d807Kbd2VFVLL;\(
Z_S[2;\e<Oe[-D&5FGJAYF)K6e,\YA4HO6M2XAU=fU:5RXGN[;E/<3^gT+CXPR3f
R^GK9KJ17c[A1>T/2?VSaM2+c@g0EWBda3S.d@MR&UGMeDO,e,N1B8GE(]fKL^,6
9.b+U@W@@ONK:2./=\M;S?-^J#?AMUfZH26H+G3:\c\&@@BMV-UOb[02\bCY]&E6
8W7W&e&M9]Y:6)OJN9AIS(W3,?&eC=-/:ASLMURG5VX9W/f+<[^#0.#)ROeEbZ:S
_^S1LKX^\M)0GWWY221F\,<2f6]UTa]2L4]Q_,RI[VK_2IO9+>cF74RRc8VLK@>X
7D;cSfRBIGJNE5&943,A.0g7+L.BJG?E6e[?LTM;XE6c@[P;f#&E0.=6R^3c;#<5
G5Q87Ee^[4JbK8BcIGYfECbD7V&:a_86LAYH+M\7_M1:gg@]C<dKNR944@_#2>7I
b(XL,a(fNM#4:aaKFZ(_EA2:;I;#5-HHf6bb)@QPE-Y:PHF./aIHPUY@ZTS8,Va3
4DeDfYF=\CE6O[^S25+MIDUAI>eF9e64_=HEAW(-I3EH8@aDD[)6L9bJc?O=fHX/
XQ[,00,6QS8XbO\?@86?<AR.(B)#3]/^aU/UKQRJC[b+T0/OKacWJC;3e=;M#;I\
-0SX3R3]B2d6Yb<)@EQ\>2]LGcR=[DK\GY1GBM-AQNY\Z_e:O0<RFKZEQc]Zb37:
PV_OT]cS6,8/Gf;=++gW5a]9dQI6B(W[?(YZO4DfJA;d09S=M5IW<KP1CU4agI^W
3a:2ZX?ZO2P]DXCN6S/KV<c7JQOBJYL);8P6MaHA:Ta]T.<L93\7\.8Y9Ye5ERV3
4gB?5N:O8QW-HOSTH3W/b#^D2UfA0J#FC+1[7;N:\ZUP[<;&a-ID^aCKbg#[_[]G
;;^LfN:2U9>T1=)dg90K?FT^;BURgT3T57;,@K(@bUBECb-.J#.+4NFfVPAYD;ES
A,dX1J_8ga927Z);I=XD.F]+c^G[Za#GNQ&AUPfORFTL0e>_.HUaE+<Y&[BfAOLI
g.PD,@2?)E3@A&gcT<[ULdOe0M3:N<R:,A[&BG>c[.QA]\&]@RA\X=#1Q[NY)dU?
5Z/7L/2?B>]Df3--=eI(+[PA;NH:9/8#DP(:71:5<11TPLQD14TAE)&LOEZI#=58
6@ZbNEH^SL-6FR3:[EIY<=QWF(Tgf7I\9N6_)Q]#98)@+LOO9SaTe\dPgMWI,?R+
&Q0Y8PUK#:6E/+0FcFF1((/0-U1cFSJ5/L+A@>+FB:-HI=bF[#M=H9LVIe>4[-XC
#Ma&C84MUd5:?C<7B2-^8/B[NeD,+0&gU@32Jfdc.=/S>Yc\8.5^V2]82\BBHc-<
4WRY0#J2)V5d\-E.O^X+GaY8SX[d](f[NA2Yc[9E6V)<&J[+#F+DCGZDL5M;2#/:
FVBK9VHOSMA_ZU(:]N(J1=c@EM?&aa^UIcF:748&-/QD^M0,XUEB(>_.0(CODBQB
42?aDJS=VGfc#9ED>>C;LF4f1LQ5dgSIB#LY5)?_DBN:L?5ba/0/F#9c5\X@CffB
&_IR.2XT5(70c4a4(#OA@bP<:ON,GN;D?/c)->N7HQ7],3UfOeKTR+b(,QJ5Va#c
^8a(->d,fK[+A-KG,gV[TTUC/cWP?\TWdQA(MXCAI6]YHC[@=G@cIZ)f&a^QRfbQ
4Dcaf&e;#VP>:7,<)/M<[X>0BeEM]SRDVLN?f?P-9e]0+926\@)ZK3>-10Oaf3AD
eP_Y<d#N97O<]F[EJKHG6fg#T87[EXBN\1:cPLMR3\/6:IH@DNPF(_@7,8U]/WK-
4?LGV4,7@+>3<YW7,&>/#d-<V/5,A08aK3Y=>cf8AS2Ue7.Jg(+(#d8F_WU]_4(+
VPY.)&=+1F08MLE1X#_L>#:Wd>N#EB&=Y<f:[MY_,+8KgC-Y+KXEMb)+1/ME3U,;
KK2<5/0^/QNPDf+2GJ1ULQ\,;1TI9,33HYcL8#@=0d2e]I3GNKH1aSN94)_T_bLB
V8Hb&BNWe;S#7TN0QEJC>WG3O#]Q4H0;/;2-Qe,aXbOJ(0;#V8d(7;UTJ7]&Gg9g
KLU]/#M=9.&9ZQ73X<8f)aHMOMR3#FW^2:dO(C(,-MJAf-AL?LRC0_R?Q<:FL(7_
Og/;2C,5[NE.(<YCgLXVgILZB<O>C.F^A9>@g-Z74&V[+LbTA\9ELTMY^@_R.d]M
[32RI(f]U:c&F6UYf&YdcAe391EI>L@DU0a>L;+]G2;,Q]6KYDQJ:Ee2eAO@P(gJ
IOP<)fPV2,^5\CRV_e\HRKI<)ERY&+DET<[f+[eg)#JH@TI&U.1<OgBY-2JfeUD9
\ZdV85Y?D9Z1d:Fb@Wf?HO6)QF#1ZLR2U/(56<b^)W0JaF:&(gd8+MH4K;;5@6:C
daI#7ed3#3\M.0fX_Jc(YN?=:.9YH,G>+Pd@Pe+:bINgLYOP=^NO@I.BF2BD=3DO
eBI.L\8XID.J<e9\cPV\U#57/C[dXbF)>Q;J-GScB1g5,.TYc1XbV@NO>#f@-_&(
VB@L0S8cTUG>1a2JK[dL]Z97Z^S,#gXJL&BK.&:C-\]Ke&?Z4V#O7//K2^E>?H?Y
8G?FXJPSd9^FIIT>Q5-4E@R();K2YCW7ZNWeNcL-(M+MS2A(^Cf9BJ7\]7cDIUV[
^C^?B(OCQ9fIZ;7VO,6a;\\JN8-g]+4:I;0+D^_9dTCUQgNdBF4@9C[]+O8Pe)_T
7eYXEbC=aeQVgB+T-IHLcd?7[Q>9G,7[FKY=.0=#8<XN<[OH2;O1PU,\N64V)daN
J>>ND&W@H5I:::V5K?A^<V</P<PBQcS21&7U=c&\.@6AHIGd:)_V6dM<aK4]8UN=
-)N<Fd61F/:XIGZSEGTbeG-O/<?E+fMSC@0bHBAMU(,0?JA06fd&UKRV2SXWU=+@
F:C>(@Ge1;f>C)<\(cJeVa:EM,[SN)X8F#e<?3;0&/M3S_^a+V_FC]a+eQA]g9]D
A[AaUSCIJQNQg>BOL8AP:D+)9UCK@S)US:R1b2DLE6EbFU9P(9:,YZ\O,<6GQ=Zg
d:Ng[F3P2]?IaXWT];>E<JC.A_J0QI<S.I;Vf)cQJFH4?<+/?_/J9</3OM&-LRP7
BSK7gM(b7[6]-S4Y;TJ3@#IYER]L<(VE2M+P^^<-S7I:D6/^V:VLHK3e@7(H\NED
58#W<YYVH&GO^CeDPU1R^7>>5#,X<TI8+U_8Q/14G6gN\\S\R]B3BXT;WGZ\ES]V
DT#]C)I[)GB:89W4A;T:D3B]+Eg&>EI8g0N@3MBA@#V#2I,0IXbKLH/39=9>QX]^
=SE^N?>47bV-M2>2#-+4b_]RJ7FPEITLT.8/2eI2@F.U5#:W@-/0\a9Z.-YIGNg]
@W43/>_gOf1d_JcIJ[5BCVP>MJ5#Sdf6GE/N(.^c8Q?2M9@<:GeR+=f6[5e4>_#b
e2G,0VF_Z]<PELce,0--@Ae#b,F-MZJ(_eW^&</bD1)<D)Z4:6cOI9E0A#LJ74UV
S^;O9]RLLA&:I^OD.ZR@TOZ2CLRBMNI93G+7@[dE+N])fX[0Q1^N60\0Y]RF#>&>
,_4BA/U?AQX)?QfcL4[@G#4=c>83(RXCD=G93:WO4#+N>AeD(>Y5ORT_B885/3a0
4_-,9;)BFDH_-S,.:,0^.@6T(X\SK.LBCKfJ35I,Mb6Ud(&90Kfb4<7@/b-4]OPU
gPC5XWTSEBK,HfCJCg4cYb</M)GP,WM_gfg#d7f>(CB@?3XHb9\B8PP=+8a;R4BJ
W+Q(3SM]aeC/WP2#)<;Q&1FdI4Yf,JZ#GD-Q:_bK-T/BXfPD_?R&&/U.,A],EA;J
898a6B@RAbPM09FZGEdHMaFM8HNYQ](T;I#::YgcZR_N(WUD-e-&6I)e6;H>1YH&
Y=P48?S1P0W=?MQ<T?a?S>GW2a@]1]^2HFLb@=e./9d/[^[=53&2g@[#JaHB/@A7
eBO7ZY_7ca;A;R1LAa=Z#73UMS?W_d\;bGR#C4F;?e2(Q3/2@,D3MSfQaHK<g:-:
2RBgR=,-T0U1^E1(c2);/:7MR<_+4=OAU<20Kc,=#AB?aX?eGP+3T:&L:=8fV(-C
Y/TJbQb:_0WI\Ae/5A1NS>,@4CT8D#O,>458?]e@R\S6HBEC5e]5A2=b(0[;Sdg_
MeDU/::L?=>Z9D=:5Y=BR0#G)gY+447B;17:2Y3eG@CfU(EZNc6Ha)<8HgI@LMLN
B)3A;aTKILfP7+Se?:;V\-[Zb_cB-7&S].+da2=3Tg.a^(S@R_a5C6GdJ_;cC04E
G5_4_?^,CB,ZWM(\>2=gH1>Y,bV[&F1:9MgGN-0RJK_abPcZZHOF^2Q<?IEWbRWK
)Dd>Q><@a(bQ1==O0N-GA.7dB.(IC,Y9d\##1dM#N]H368N;VRP9G-UL[1S5e:T4
PH\73[02NId9J&0CgFac[[7gZJD3=1babI\ggB;:<:F>M:QHXgQaBXd#H1/KMDQ;
/,RaeMbQ>M:SJUb-4)eQ1OTDY&Fc_V55;DWd;CG]2ff@4,3PYH8:[^)7#52)+0\2
:Nb,].5XLP?gbVN&>2FFd(^P2649JbZWZ<c,TS49_b.9YD+=]7/?X8)L5QdW\)^B
IeYAY7b5,ES\:6Pa81Ba_YVOP^LZ\,1OK]>Pe>IX^e3K<0+XPbN-C#&F453MWc-D
6X:_&&0KA5[^]eA<XPge6N<?JH30]#YDHTZb?DA,OU3/7&9>MZO/f4ENce,7._9?
:LR/fHge7(T+(]G[9ONS7MY:PTN7[NQEe41DO39G60fTHL@c2_.g9F[HJWde-NC&
UEdTSM@[:CA;S8<&Vf>?F666Z?0UAfCZf&8.A&Q_bMR^N)/fIA\TID3_X,gE)>W>
eBX5P[(;5X.RY)^bL<=M#g43:7+>d0NB0\@U84W>KQc1W>T&&8K75#;>F>DG;OgA
8/T>c<.eID53]&:^^+Y2(3]Ub>26L9CW>O<_dF=YGY)e[MA8H[fM4=<+QD5df7:/
&Y6Mf?b0K\eUH/(fMYKAPcKR-I(+9,INS[A<))EZ>F6[A(/SFSZXB/DgJA&8;b^2
@dK6XL4+?6/gE[YP\Y=A?-[VXE^);5E(^L1dVG70NAZaR/]6Ed_e2MJ,^#D52]8Q
9:g^WT?;HPRb7,@-d@8X-)fBa2=-dd>DBGI#PHE0;9S4F2M<^#T[SG-FCR<#7b/C
^dC&:R:67NF_KNL+cLAH.HE6;8.86EE[6M0Z#IV9VZI:/_,@ZWWdDVR)>4BMVO_f
X=?B;b&VeDYa]/a.+C<NdM_bI+:4XG43HB0?5\H4O:V--H,4PMCf@)D.gaQ2c=[A
Y+Lf9]S+]DKR?4/F>/8S8Z_YT6MYJA,J^,HN>b74(2<&I\@f#^gH#^G4dXRe1Ic-
If99?3@GEgMW@c7UPO3K99bP3GQ5?Y7O]X+<0/P?79K4+>PD(Y,\Z1XTc]V>g-c]
B6_5<.^b?QAC=.J;8aKMQ]&.?e=2^GG;:)9d8905O<>L.L.TKDJ-:OUA=2E2EcPZ
OR<X+S)<WW9PW1VV9O7P/a8ZP(J6>_>8B0N:GddA<6Q56KVX0VWA]G+f=.I<0T,a
N4PK_<-UR]5c>RTGGg9N[(FbP<QK]^@2\1:YF;eE7CAL_ZDK3+0LgQ(]:gOL&[dR
6KXfQFV+FXD?D.H2,2XFe+?ZA(f)#=_=V1/<\\cEA)2fXQB?AWV750cIc0DN?E;H
I\-c1eI&Sf0WCQ\Ke^&(#/]g/.TUOKEGfMFGCSfKd<(SOJL><TM+_:ZPD=N,)>a]
]_F<eUQc/5(d)Z.)K1EIb9^cX6<Dd=2B9ZGNS.dd^ML,RMB,W4\gX>+/=EJbcWBC
dW3\GSC7:=cDP\D+C]=JgY/DD]@?+1Pg-9T8Y2>Z6a>7I=W:VB9S@##MZM.\EeIO
-a66P91XA<6=/V/7e+N7b=NGV[=9KcA)&4U;L=;6GRGS>[]RNK_c;DH,IC0ITf3-
+S@FbP,7f?)Q]TS/RAJ.G8ITe,0Z7_c^A7\W:cf6.B;0e8T@=eBfDcJMM/+?fdIH
(SV4NT=c3(<<G;ZW6BO5<L=/MEIS;CVW&c>#@4de\+LE(U,bX7MDc93X2Q4I&MXe
7Z[XM1ZV3>aF]?0_ee_I50GbF?RQ_^d)XM<ceJbN=<C?I;JXQ:-PYU.BL:2aPU;A
XQCH@a^aR(7bWGH(RG2&53M1=gQ&D)G?>?_f.fa/g0E@f5M?1^\,/9B7?Z+(CS]R
:f>/AHO62G?4_cU^.3U3W2c7+;Z#(B.CMeC48?Dba0bUWW&E?0Ea(aI+[WeM>>9<
LLa\5]TLHU,<4g+@/)32WJ-,2DA)\UNS-LQMEbgMAG\IHF]A:<DYd\,QS7Q5+8I7
<PCVN/W4GeZN0<dJV_gI_QQaCO&Q;-=_;<<g-L9APFFD=QU;GRK\44_;7_49Dfa_
4-5C:::MN<gXYR98()63VQW7(STO<SOQB\<K/^GEb+bJ_5[+SR1]O=<TOd6D5^a,
Q5__R867>V/Y=H#B(C#OaTWN/;>+?#6FaSZD[8KTDQ\9:<.D,&=-/BE.[U:1;&#F
:bf8;LJg&:FA0@Gb&Uf@HAY([EKNQ<)?f90MM7259I<cV_CRRSHbK6=+1(7-e.=I
?#33adRM2,K(=Jd+[VfVIG\bV04]:<WSIL7)O<^P](>bYA@Q_-(5ZB?-.P;MY2E]
X25_/IQ<:6bUc?V]g4e[0b=(>YU:,f+#6=VJID^HSC\9:]EX(,QDXCVNV;9^XX)5
AWN=Gb;&<>P894O]2@,#N28+Y>a[<L5EY=Sf))OA-#8.eMUaUN7W8>X@baBCI.=&
#P)W:I)3aMY=gZJY7P.,[3EOfa#H5&0TS0bFa7YgBO+K0A[V&J-3B=^N8R#?I9E+
bO[g2GC@?9?A8-e?2I_Y1B?^4BEPR?T(CSEI2G]D5^=<d5CbQV:S&QL/;#7/NG]E
>(KCa_)]VNgfYMfS6QJ7N&T465_]D[3JF_Y]b)O?K6gDXD5e,A,DC\-fB?YE0B^^
#M/I7dgAT/6Y3WVB,Z:@XDIW&?/Y8.FSfb=:eV:5KU#Af2N?b5-F&X1BL)_E_57d
6b@b]O1AE=,@V]cM+6GN?/7N(d39Q(Y>KK4D2W#Fa:KWAED=Q+Zb05:H4CZ.=CHC
:B,4<?BIPCXA[6aH#DZKU1IN1[7II(;[26U=G4(Q0#M9MZE7(CO(F,bI#/b:TCIb
._#ECfaVW:A4W6?FI/QH\BW4EBU(aE#>Gd1I9b(cSOF6Wd;2R/LUZ(F1L-T?]fG;
(W6D7N_.PU(-#OPH_D#Y9)_AAc0O?N[JU1,W&a5#[dH-HW,THgQ79(CV/=2^H;LP
;(]_LKC7&Y)7V+Tg2]0(g_IXQ_GEC=9UTILN)/4H:WNAFCQF]>A:0f?/Y<DF3][3
M[6a1Bg(dTe;2(,B<3C?C55,Ie;8#M[GSDR80]=C:<XE?FcL[((@M0?fJL_W;7?_
4/5&CMCSM</JE\>.++K&L=?H8I@b-L5V[Od7(KaWCE=6;A=AgcUA&:X\eHc:aCdK
&G7I(F>G#],dEMf5bUO;:[2&]O8af(,-<VLWU#8P4Fc@Q^D6Ff^@gGG5?EWGE7FY
7EOLQNG>#=2I<Wc>g0AYIY28G;Ra+?C_3]D;?_?D+OUPY]A[@<g(BAE/fcTDf[H7
\2I7NM3VdZeg5NE:<[3:=N:O,U(2P4LQHH]Nb7KA8Z>5U@O:UI)-NSN0,WB:M&5T
RaYX3Pg2_LD0(-@?YHBKBIDa&=O75]BFD=2IVY#,J@4If?J.OES\A3(:OIe/WbY#
A-KeA@[5B</9@KM?](/E>PFf=2HM3Y43ZSKQGJcd<U1;QU734H]5;AED[M.MO#aO
gPVKGRVWMgEJJbX2Lf<?I93Q[b\d([cQ.1=+4(>aL19@+UMC)37ZX]gWMV@C/;9<
:_O4T<939X0O@cgNFP>A>E^2\a@>KbL2LC)dH4H:O.61,(A4HRHe7IOafdaM]:4_
(\1R+E^ZgC:,4FJJ.)bea6P&ZQ6N#-\6:M\ba\Zf1?Q7YQA8SPa=Q2d3-(<cL/f/
PI#_geX-6U-)6(V[8=7-]K(.:.6S4H#8]f/0aBU_^&5+DaDT8:=VLe\8ZF:Y3FM_
Zg&aM>F,OO[1JNe.d<S@L163+R<A<Z+1Y;S4APC#\Z,0E(Tc^dX:W4MWYf?=LCO.
Jd0>eCd@I4>CGaT[C<-^J,EY@0e>VK]LEXaaSb[PSf/MRNK0QL6=G8RU+9JDId[=
3b3^MUeVY7Q&g2=bZ/9dY[;1aA[JHC/NOYF&1(FWF.&FEH>e:O4A<[NL&Nb+6&[<
?:P>7Y+GX#aeOAU8I836gU2VX)cfQ/.d);TB6cV_?e:T)gQ[Z:VHHU0.LY4H-CRY
;,MBKK8>L1IbW)Hb?U-#<I6@8NFKDg75>:_4<fg(LR?+4][6RbM-X_aeb;>P66K-
8CaK7KCF6P:BZLUSb@2C&2O1R3JPfUI]6UecSa]48BDBM_37B2bb]G,#39>&HQA&
cC9f^6]MP_)QAaJX>5T\9Y<;STKSACGK[9S(GDA.F/<e_YeCU4AbVP_R.\5#>8\c
J6Q+L_PRX4Ta6AS#XWT1^\8d4G==XWg;g6]Eg(EBQ#MU+>GG5JZ:R)a;e0a]@1g\
A,P;X-LB[/,=0.G,J#H)71M_ZZ7+XWEX\5g>:E+If)NT7+Cb+ZI=;eP::(^6@]N\
aDX]aKW(Tfc(gNM(SGRVVcNG8T>DVD\_<8T[Y23(7FM7Cbf0/P?5#AD^B,VC^ddZ
KDO/9A42\IL18L&3YI@T\UV4=-Y6KU;^[^<K07:WQ-.U\IF9FX?:],JOT8<(4c;7
Gg<Rc,\?L<Ie7MGW3.?U&?OVeHBU=V^<Ug.J+7IH8b+-UU(JW75^ZQeFHH0:??)\
#dPV@NDFa(DKNEH:FeY;@f)fSCTe:YJAQR=SYM)f0GBO3XRW)+W>T)@73AU5+_L.
&aL?SWQf].0(eO;T(L1b6^_BTV:65YU9/UCeO0c2e\cLGJ6,VaFP]8[4cQIOFS],
B8K[SE6fT?#R]0ABSHUeY,>PBW+&ZO4..B>[F.HbGd2LLG.78b<9?)4[8WM5D,9-
9KT^MKKL,EO4K0Je])a1FEP,fWIB]OL/#C-@LK^V,2>TF=e5OdXgPLbTEfRTV5N+
(O\H/^8E.9eMYM9.;/</9QIg+5I5SZA;fMC;1@51?Z+8O(:V]b-9&V8/U[+0c3;d
P.bBR6Eb,c)GMF\;eSQ_FVVTB2KYgf._Tgc=^;4CBO@V,+aBHA->b@PH;[[F5;3(
<a=eBM:TTWb4-9GW<fe.SM,TC&O@;#.;;fR1IZf[2bF(B.617_W.eMFTTMR:8]1U
,/DUVNG4B->@f6\^BS68A1Y73R\EBOga6&VN+d/9\SP&#E]QNPV#UTKV0(XCUfNU
2OX,ZA;BV?B.EdJEKa2G[<6_S.dF)>?Ob-/7=:FOa/B#1#UT5]2WeDSf3J1SZ,c(
J(PC2Y)\OBZSa00/X2?#d7Uc@G7GQdQDA1V/2+<&:RX891Adg09[I</Z^\)TeF-@
:,dZ0PZG74ES;_&0\3U\G-4QfP3X/J8#I@YSH;@[+&1>;CH^L+YG5SPY):H02^5\
\AG&&2OH?7NL,L3b24WKR+b;ACS3Yc#XQ;E4UJ3B(UOAORAB\d2NRa3A@XGa+N-P
HI)/Fb)>38AS<=W&g[87_=EQX)=G:0[,IgJ8>#H#4=WYD#/Ig4JDX:Z/3K#Ee_>4
Q0[e,?bN&E[gc#H+,TAD\BE841D=>SBFTMIM8++TO-0RPA1H4=F_UV6V#M@dGY]C
KZ.S#NR+/GDZ</O^]TO[#Udd<Aga,e3HW6aP?fECLQJGK/5O.?4ZYQQYFH^#D;X^
YG)P4FcbVVC7R^C2V9>/?&DfAS\;GNCcP31^I<[]-77\@NGW-fX#Og^\(]2LTD?J
_2_&@0]f[NXE^AIK6<WT@,<9C/E0(IK_?aF85<fG/+_9DaQ,O]RG6R#bOg5G)#H(
8S/&Z@[.J272GM5O?A5<3-ZPR9B+&e\3J=GgVBU[^PO4@\WWLL(UNWOMWEb77(5e
QR\+e_f0f^X4=T(2Wb8a]XMe:EVLWO12S@^H+,\VXX4U])C.CH:f,a\K6XW?79(_
e[(,8;#-K)_AdS>/8ELQ_<e2d](/B1Haf]=XD.ZLX2,9Yf[0B0)AQ?^J7;7&f:c3
\eV,4>-F<XdFD&;=R++VCA>::5?Fdd&+W-0Z0HUHdTOLN>(J,>@P)CI3W=?FSF>O
?bF5-WG]B.)?-/g::aRfE\MXg3]3(W/RZKGb6Ic]5-5IF]RdBC9\Lg0e:7I[TMND
dgS^L0Q)>1c0[M>JA(ZAUdP)Z@F@G4<=DWRe3KdH.)5CQB2\f:9Wf[KLV(N&;f/P
=#bH7>,AUVC:8=A+2NT;@W@F4d1XCf08PO4+c[V<41c7_M9&R]G@LV,5#MccQe3C
\HcTK0#<UZCBQF0MdaP@.GF]\7-]A-\#f\V8H510+/Y#,:)44=LQbK4I8/d1BdZN
+C_WNTSaF.J[+?7)M_YT/K9eVc=D:9KO^.,ebf,d0(N12MGBGE:I5UaWaUfJb@U>
FeR36\1\0F/.3aM,+E:V_@FEHW&)GA@6A-<J?IX(#<(7JV4ced0aC2P.ff@<VObS
@W8G;_VHKCT49fG+QQc_+,DCe)77]g#-^K4.bMGc_=\3NTF3&FbAae?,J;SdfFdP
a42SL59HaPb1P8Wd>3eGX^]TK)4SNb3)#0g5_VWWS7d72#HN:;.-QJ^H>LQ_DW49
HP]&M0M&(RJ610E:Q:^+ZWTXF.IGHcNC+=d>&2#YNSZ#C@PR8J&TVPPOI7#Rb#\H
Q#VLJKFc[43-K]5;Ld<K>,GbdWc;VV1c#GR,-OQX_c;Q40HW_>EUX\SV?\W,?UD0
@7P:IQ3NC)C1[2QS&)SJc,IZ4]NQ2f(@:We:a:BI7?5K]cQXMQGR(O+2GeG3eC-8
a81+9I@[CIgT?g48FfdUb]e:6/#NY;_.2=/-\VCKQ4)Y);>&,A2_-^JbO_B9<B55
1+1W=WSM.?#[W1GQ<9/J,LTG.b.L5a/1_aO^Jb)LOT<K2<??2gd9g5<[=S9IQ5e^
1.0N;OVCeDC2A@PN>8O^1&>eSa79C2;N8c6[K=H,@KIF)E.(Xd(#84[@YYNf@\/X
7O[W>@,SdL=EcTMO=291aASEa&T-P;B?+U?cXA8I))FgP/]J@G:]c7:;?-Q,X7RU
.WUAMbB@[&C3(B@gbJ,8AB0ULKRJ2ZN.Ya_3#0V[=\6A2(R7bLG8):2gG:C5S<]W
f]P@F,T1(I>-X)c=Z6C5T[U]cN+W]CUODbVY-7Z9:=R-2]O17cCGaCgK^&cS7gU2
(3R\Q8TTZ&,>B3MP0Y(#a-+LcY?)O;LFN6fYW+0Ze#DAZ^b,MNd>[91dLA>H>B8W
4UX(H0AB<fSa]X82JF1g]GP<a1?S\MW>6O)6CA7<:)d)27aLRg>;71CNZMNYWM+=
1L0c5\LYQQT^A3C(TS[AT^0]T^;(AR1:;,&DDD2NM&Z45Z@Y>V-+WULcK&aQ>96E
#a+S3C7C-BWI,e(8,3_OfCA8.+^&]EUG.<4OCXEDA(MC5H=4/?d?Q\7b8;(62>dB
ON?_bDGL6_1O2B@(ePDU@;3MGFIKBWZ&@D&bg?&W_2Db:Z8\&ea]7,ScDa542Kb-
JT1L5HL#D[HP-,E7dB?W+e/Q&YeUAA4X;MfeC]3;L>DM<:3/D=XPS_PB#.9H0b6,
=5&71:J8B;;:C^_Hc41#-XcXTZV_VgZ,I??ENd^AMBCZ]RKf#6bU[fETM4cW6WLE
]e.:cY_U68Xe5+V,2L\^&3QaJZ^3R9K/-fID(EN&d-NO5S4c8UWV69<3c#1KU3BW
)Q-D0RQMH;CX_B[ba6CAbf)AX<?W+8:TI>)-J\[V1ec8b#8Y71_U#?L:J3Ub5@9Q
WIWA9R)W#0>Q6QbHZ3a^YZ6W+dHTH5+LUX.(eV>V:\+N8,@2Z,2N)WF,=&OYP#B6
5R]8a-eMRG\8XJca^\_UO-#T:E3,D4U5#[a8b5NN[R]N8KY[T.>fa1PZN#CAG:Z#
XRQ1f\D<OW2,,;E-XKB=@>0T92X;:3M4R;RC]f^;Qg1OV#68+OAKeM/Rg)H9RZ:[
RZ,S>2aZ_b_4GJN(]+MF1\G3B^)K:f2UA>+7&K1M]3A)d.T;XNe^XD0=M_GB&\[Z
DWbS3L4-(_8H9G[W-(X_dfaF45?3,FWANPD<24,/P)&;GI:4?>EGI-_](33.>DaK
+UgA3OA7_+3T,5_V40D@ZPb90;(FXB.M,<Y:;(2>08H/C_W<2AN#2JAEC&)1:)dL
/:UJ(C,OH@REUC//K:MHR1d<@5,aF[6&3>1EW=,Xf[.RT4M<1#G_gBgEcf,V3)<;
X8/H;U8BIf.)Agd#]efT<<#=]Rf+W=Wdb0BC.<ZKBI;@,QTB:D6\@_c[e:c0\Y]P
_LF>M:/bT=a.bM<@<ZODFS7L8PHN1ad@R<--4gW0.?=C+A9XZ1+A@OY50+Y8^6+:
GF+c&\?-@,3gH_+GBO1&&,0RbSdU,JU\BS9;]Z(5_G@8SBPD4K9U()_aNZKKGCH5
IVMZVPCZ[a9B6gS+)IZUK7C=(R=D3Ga1A0\EGbU5Q+^Ng>]d9M4Y+Z;3B(D3T&F7
<H\N)XTdfRH]N+4d0bUICTWO<[-f].\]&A&bJAFE,(\L]F4GD\]^BeLZ:CEADYT?
+6-e<3Q:F;?,?IKFLfMXG2;1bd8@=JKcS&=cEa/KYW4[[T;&Z1VZV:Y0:VfbX00U
#E01R_YZEJ5UXA<C\PE-M,0dY>J#]GAX.FNLZ]N,7eGEG&?7VE)#F:f8OS1+g63W
F<EP>>Ye\^33g44gCUVa36JB_Wf:^;ZMAfCaY@c@W2)3b^;\EQfXM?5LX&D7Pd;b
9UdaF]g/e+HN<C?SGRHM:8g3Q,=,)J,3;4+ZRN0,)/5I3ZV@-),?LW.-6A^LE3)V
_<_387F>=cPe+K<_L^6YITBaE1,GccE?+]Cd@R:FN)EeQX1#6LV64NeTND@XG;X.
e1fA-+e3+HM3&BG9.eG#<1B@P:KDR?9</E6@]P3/J_<5L/Y:C+(++;[AcRegLXcI
,J^1^Y1&35]dQH1<dL>ZE;&G??&4bee?L3^&63-N(BG(7#OgB<\DA(.QD5D#GI5a
/&U3V45+_,MM<1+F5,6RA74aXNa^42.5NWL;P)CHFO/?](CfTU1@Q39Y^0IDPZ/T
?.e845f[26/fX)H#3/5<&2.,&H7PDG&)5BV7;-586RLf@WT,,>G;Qe=MQ#++(VB[
&ARQC?B5)?Z-\_2c:Wa0OSXf,]<-b3\P4)e;[L43e#HGQBe>@HJ<2Q7^\#+BN+/=
/<CY8^ZZEbV.&+5&_8,6P,SGAQ7S(-TX2baX(#+0d<2WT45K)&825dLRbKOeU5GW
SCDJ6?,cbJ<0dRBf_S9.M=,&Y:)DS?J+]NNb[BOMRe;KbQ)3GLA1;Y\D8d4W\7ZT
gOSOaI0Ydc4@OIU10=@XIGd-Wg3-:7\fTc<O1]U[LIK8Q#^Z[[4f/]ZXI-)55eUQ
b)?_V6E=G5+=V&]MD75M:eVM[708G(X;3a[aW5OKHgT4BBJI+1]S4211LGeS3>=(
A?MD71bQ)5,YedfM^I0R7D97KUD6Le>TU<L4FYedA@S:(_[FbAZe+8_EFE;B&7dH
JVEbXYXB0UGJ&Q?DL5c,g3;>>9,3+E((6PU+#EU6W0&a_Y,L(<87((XYQYCM\9D]
RLE+5@8&YQ1dI1EZUI>e_PK6UXGSTg3eV=.NfAFJWI](IJ[6Q@9)Z^[7VOeXLYcQ
Sab(JN,\8&gYc[g-L@IA5R38?H:YRAEKCJ)WXU+U&,eaVJ;(XOK0A.B;=OIgEb.X
)OD@W8eFTT/He-GB3K29,IUd?Z&S-W>X@.K3PXY?B47A\/Y]/:\ZTS&)#BC27,H[
:4ICT#@BY31TTH^1V)NQ&3/FFQPbF6be.ca+&ODN(cgMVR\dR+/aXKVZ9c[:Z>Xc
-.,5Y>D.7B67g1c&SM4V?NL;H3U+^(Ma(=+a3(0]32@4K@:_D5;0_eCVRS/eg;cZ
SM4D>]5>0V&Ff4>A]DH5F)]+f]GBaA#TDTaTH,D8<SZ4Y2_DJ)5aM]?I/79A?JBW
(]2ZSQWTKR^J:Ta\8#D;/E.;EZAFHF4Qa4/E./L,K7OMcK&8CE=:._==T>AM-fWB
CQ6EQ^BTBS_Y6H,MbcK?>DHA50GeH9]c;)#=K.#UCBa@&LVO4=23e4N1.0U;+4,_
_+NQ8.7@gXW.-HT.S@BLYH0BD9KEb:g;MHf:@9FIHDfEN(+U;,)(HcDHK_&fg2+b
H],]BDB[UX94IULX\C0Jg:#S_U#B(=[a,MZ(CBT/YP?6(09I1Y6c8[6OL-WIQM>,
35>ZW]J9TBaJ>geSTHNR\\QL:f?BH6VKG9X7bY@0a=bH4RY44ScWZ#8BOfVHJ5,G
BLBa>V>\T(T8gdWIA(\3M6@=-SQ#O8g58F4,I\@4_a[Q2K:(RZ[>U:HYCVgP6&OB
G06IKXGW2-@[#.Y694Q7N7_C#SfF,>H2DFM6&S2DUC]&304eVANI#>M2Y-A.^AHX
D:#B097OW#E7XU2@f,>Z5[+0S[5/XBV)V2[0-g^H;C9&5H)gQ82^MgVV3V6<Q[F>
]6S>L.G\Y,)VSb(27a8<a,&bf_H7O&P(9<J/WMbFPTB^<GQR./@dM9#cf-#5.#W1
K7J\PUX41J+^<EE0\b?((cVXQ.H8^-9;eWDKfWAfW;bR^9Me;DY1M6#cP$
`endprotected


`endif // GUARD_SVT_AXI_MASTER_SV
