
`ifndef GUARD_SVT_AXI_CHECKER_SV
`define GUARD_SVT_AXI_CHECKER_SV

/**
 * Class declaration of each of the error check stats instances using the 
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 * 
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */
`ifndef SVT_VMM_TECHNOLOGY

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
JVExvbQdRcxnQs6fMjsqt+Mbm020vn3lfPrh8uVm6Xfg99haFZnma1E1ygLfur+j
35zBV49Hk/VWnYUjz5hERnKIDBWF+xatu/v91vfmYC/NTwKOWg+IQnYprwZSW9FE
IOvLnAjS46+MBmIBwSCG3kpRaULNkA5V+eWKxeVI4Co=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 41456     )
vQIokPnjjKTs/4mSSMKioiOWccw48PESMwPzLEp1aJ+awPcmiWr41tmmoWW/sz+I
nwX5PEl+HI8hEVE1hXJ15rIBrQtK99IJL/z4/C/wyMhzVO+6ehQArVQPc9uj7ruw
TzKRrhtQdFc0BMb7JbtA7B4CLrgrkMMT6jSBfexj82gGJCzJTlcZM8MtZDHHqRWN
WuE3Nhn9JYEPf/o14aIGMIHJM+/CUOlsadHjKCGWVX0mURKRpd+tGjdOnHLQRIdJ
4ucChjN9Z2ugwLKQ3/BAk8BEOMDASGStXxX/T0LPnE3e7/RrA3ajF2ItC6Y38tZs
r7gi9FUf9uZH8ccy89/mFpipcY5NcArQhukX1NW1QbifMimO96LuNZZe7DQ51F+R
KEKrKGXuDyTVfBp6pb3tgcSHLRORnFrHgyAE/E7X/1zSPN3E0xyf4+tv3h0wk00b
wefKwncKbPHzue9A+IP57ws1wxboEfmOoJ150erwDwdDxs8c56nN1dcpNfz13KhQ
jq9DjZaswJAIwnbJgFWPHZ3dk4MTN6Z0dRyLaCR4i3yg4HprxreWV/W00u9TBckm
yM5xTheYBO9Bpj4Uk7a0uUg9gbokNN9xdVkV0nKuhrS+AFQmdMImDU0daUS6tVKV
A1TF9UlgBIQZq6U5UPDQTBJKQWKjD7lK+CK8Zg8fHeQb6XNXjqIFlus3fsr/gTU6
MTcF06h8+RJl1axGGLMemzeX92yF4vxnJXdjTEbJIUAVPQHPgBwUY2IzKKHz+o9U
i7HAG8oPDAQzeZTpUrdgVlLsNEct6bu9d7dfqLZ3e5qbaPjq0hs3KbtDO+tkY7+y
TUYYtv639Pt/ElGxN2l0fvMsbfciOdRPma9L6AM749spUKNshhzv/873CqfWnaiK
kGSYCPKJUNGfyz6ysoMOyN9WWSN0QSyuoBo6KpSZ2pRPT9qXXmSiMJuIgUqCKsoL
9uqwBuQo8FI8OgcGZQ0nSSxIo/dZzzyQ6c8WVV57lwENbZSYS8ePY+Nk9i8GC797
OJAPXQ6LfaLlXxbQztrFjyiP1su2mbVIviMfsjGmwOG6BdgWdarTtlG0e0bmtn8f
A2OhjyCI++5xKEFnqtYAUmTtTs7UPZ2Mm+QcHS++RfSK7/ZgOXBRyS+dkXG3u35H
2qSwKmw4uodrZz7zu0S5tkigU073NqoIRlH4oIgmsZJyqy1vFR120vXiYxNn8OVF
4Tjf+sDu1N1pMA4ozZu8mcQzE7T/1cMJH3Wrl81Kx7iM3YPnJgLMcBcaF1aPR767
fwlSlV5yI61u8s284IE0H3CNo5+cn6/Iv11g6q7GdrZGraMqlXuHL83Rmf+04mTZ
56go6y74kyRTEs3fOqBupMz0u3GSmJEXUIdUWMHEZ8MIcW+qGC1n4rrVFXlUz2NN
8jEg0+mKYpkbWN7F0WLkXP1+oXxnyAqMxKNK1EeG5a3j718In76wBn78wamSrzOo
mr0GzFdPZs1u/uh89Vg8r3LForOCKhmweq/cq8qSrNJlBlCsRolh9MH0uCCGNAEP
k5S+R2AnOaxEDcdoNoqCII0eBkmlCGfEz+OxzbClXqRl/0ik0AIz/YAGHWbk2s+Z
I9OyNNvWFZtDR1GoaCSpFD/7iUge03mZMOS69YvziDvo55re0N6CSHGm5oxqyqmH
nItmM/CPulxdOuhfAS0/Ea6KY6UIVtLHazgKkHXHX8uB5J7P5GOfvMjo1tjRMxoW
Pz3p5EWRQLKmftWjTSZMX7Dpaq6+LD4LMohUXUrZIb4MSvlQOsV1QX5L/C/M4xgG
WFwYItudHwV4x4njOa6uUGjNMnvL6jL5CmLLRdc5VPbOXK4ZmCVXcC80SKfd51Ys
aKMZAyFPNGFAiTiZLlo39TuJ8nsWVBmVos20NV4Qh+1gD+GVm7w8xi+Pjxgvls5U
QMitD3+A5o1v3v3I3qXGA5HdTH9O5iVV6H6dy9yr5PVZcnFrcfR0Rs8grAk+5gb5
qp0h2pGxM+U8DSmWAGPuiDYdg4yZXfvu/8oMJy+ZI1yfU9h98BOdgoiUFqQosiWs
Adhq8UlF/93Un0YN81sOleITmGA3Dmf+YB7gq1Qkep2cdDXHfLlALBFT7jp/IhTC
cScgL/cwh5BW6Aws5qn8s5JDCAnF0WnfdA0D10mfIhCnzoXLIPUY0zYK/l6vX0cz
4Y3x4WpxSeIeLGK7UPZjGUemPbmhSsaWQvHzqBDGWlwUWvN2lGt/wxJRa2iQVKSu
QzCGiLwYZn2sf7MgTLjvamZ05e0NbW8M6MimgU3XrsPm096BtEIGQdFg6IPUDnjE
sggM27v36zLhps1VBNhzUiLSK0Vtn7YIFHep73E+p2Xi15H0UnXOd3yGhHqDjMti
jXM8NNTJBO52de+qlIUwnpV7FUe0og3APSGYB+b5XbOBMhiVKAyopm0mR5D/9QAG
M9s9f7618CXOpk+fmNZyt+xx6P93K2S3ofmV248084Kb2df2MsSfRMXjN6005Xwh
1lu2nllo7546yMr4UD6OehdujIcca/Qfzop9f4+DG17upN7d3/pmR6VBS5cIy9RT
iLeSg1K8nTH610VUU1uBBZVnSh/SqUgmGTyD4hXUspjWqdKL/F806xguUKua7zUS
JnOAsXUe2n0p90yWrZD6/vTKGfw7f/kpdxRD8uu4+hQzONGAKyaVcoMX9bJBVH0j
PyGo1WdOPlkUFXeLdgx/TW4V+LQt3nK3Vh1WLFQ2Szvi/flQ1BuhC9sNSZ6C2X+a
tUyQykhAZh0xHm/b9NK7sGC6LE4NIJIJ2ijsrB5VAEzA2zv4nKw9yHQx3R6yT7gT
pwmaj3pSU5Hi68QgCNqEo1Cko+QI9bHan38MaWk3DJTKszBdK3ArHsJw4gTM4tRW
LNs23KmY9PgVNQPNNCqB/QcIZ8zSLqctRLISp92mXPy5v3R+T4HCX8IlzW/UkkjU
TRcqgn14PvkfJA6ASeOgJLh+pfPTF+DAA2LHmlKefyayQE2bH3GSzRsbuCgYWLWD
2sxUH6xLb8fhBp3DvbbfjukfLIkg8ezRbOweS/xakuWjB+b7T2ffiyX4I2dzj25d
OUT5YRQMhAVZF5YDImwP7cfFrjg8gdMoDWhRMiEu6IpAXRMDuEPnZYnmJ5eJi6pN
7xf2QYxlQyb8v3wYBspUsL5x8hmQHqb+/JqSX0AyVP4p7FX8Gdz3DgirgSJipEGp
tXpSWthRnZh1BF2FVxHj1Vsw28622V9lNMzVe/kPLfcqi/6VCJzpdoZ7AtF3Q5fm
18ynwhCK7Abj5iw8aJhx6T425Lz50/K2iKRmk0DBCHXIDWFq3uIcQha1Lx0hYoGZ
NuwWzx3ysEawmqzDLfcYC7ZtfWs2YqxCdwJXt124NDjBJmAubRWhgpSZftj4DDk7
Eczv9m0hejwZ6g5K2B+G4PhZzJXt/XwRbe2pvbI5z3y02jWGVOMVDFskZLjre03g
uz1duxip4YVhK1kR94Q/BGPhwjokls+uhXHIDI5K4sNWCBJVx5lYxcyb50lf5EFD
MzrTLf4flwO9J+GrHlhdat4Cf7qqJDdnIWDSxUDxDQixj3g5QOKk5wXQrb2fRm4I
WPTrIsEuKFOueMqyOWdmUxqajmyEhH28I5yo6UiR2sQ1j0kiSrYBRGZac6B3L8sx
WrzBlXjbnFvoB52s5O51DOxfVQ+DEVlHAC4GB9vtqblPfRJffbRXLbZAUSDzrkc0
bm7bSCIClMiZ6YgbDOzsIXv58Xd8GxzzXdjE//dk/h+kLiV0zffGiPwCA0ADlLh6
n9Oj42fPoqKdTm/Gwfwcfk+puk4fmJvaNWNowlFLrLuyfxT8UWsPXQ+T8G5uK7GF
hGzEk8F6/YKXLSmogzEolnYrumxAjy/qesKeBFJunTMI4WeN2vfQllwKWsMCdudD
UoZKcSUS5wEqiNiVk4xE2j/Pluz0MZWN73ggjWuH+3GYCPcALrc9tTjgXYWX50cQ
GjypZGMjN+vTT111VuzBJwomDiF1Fh0hs7ssFloG8sfHFoUUowtPNW0MwPhQHDKY
kNhcafhhCRL6PLWGLv7grU09aUFTwNbWhTQ/Ayq6OTO50buYFKH5+khutjfrztOQ
SVHM/a5qHfcMw8mU1DIjXafV97AdB91v3mGZpx5U0bCdbJwaVzY+No+1QPMTx7ZD
1OpTxPPLewngyB/Fr2Pr1fk8BDhoA4p6br6xBSUJVJd8gkum9gc+uHqNAO+HmyOG
5Bzq0VwdTiV4Pnf4TS5YZS38Tuqi/6lgiVtOAeXpwjCfnXP4D94JqHQZuV/ke9Gq
k4xRyRPOwB3YYt0yvoai1J3x6xQ53EPbKApu/nalw/LabUK58OKSkEEPqpnwmQTd
lGCjN6NVARz9qxUjMMLUJfR0IUwpq92SrwU0a+bw7tcOkQR0iQ61/MRYVn7zmLlW
TwVO2qV1JovydTfQVuLAalddBC5UXPp3hd1uSEq8FGag2/pMSuJzKUs0SLgd7FwD
tkWtuM/iqLiFYwKqLbPxZggccDUs76AsURkspjjC+rKzydzZYLgZ5maX8Xi2puwj
YOCnsteiUKoWsPqxnJ1ySWjSQZMBa4YIg8kE3HM+3fHxPXH/TAVK065xqnBeMHHw
SmfCm7X9h+O5zXU6rblUufV5swWOeSg2LPgIDAUejvWmrJQLeJEuT0Oj5vMDr08r
4OUCs8bTiL9BW/aIALGYsEDpSXjMXIfXAwynOB9IzqgtdDqfA9So9wBOOm780Th8
Ti1GtzkyNviGW3/Nx2t1WDhhH6hQS66RN3OmPWCob3KiCTD3HWjM3nakMjl2tcxq
nDz6UpcoOSfK1Yu4BbesMqPMFzwX3JeRHrqvz5Sg2JGjUlLdHuCchftxSTiEx4+y
P63lRcesyLUHR5rGB4xCzfISs3jm+xbp34f5l02cbAhmwRxbWDEMyfH7PqSBhhJD
SSratoimTuiDkiUMChtHXoR2Q2/MmVQ+aPyKLyw3O0PFI0TSjt22ics7kqbVLZhP
yukLySFnKcDwqWds+3immwS1YlPzZZ0dby/A9rAdLJTGv/MCcfD501JYGUow2z2v
neiy4BpO5BhfsMQQ+yx9bmhVKhsxWB/fi/loXty9O5ItA/W/sV3gQ2Rrexb8XGpN
kIixD52L6MgRwClBoIgPQCiMcFATFYdJplpxUl0HeUDneyyo6l5gMnQllU8qU0S7
UuRCU7VG6BjBhcR3aLaEvXUz1iYkniD4wInzi51ylITyyQWyRDBi7DjAQ+/NvL56
TZvO5OORQJRqIMC8la1o5Ie5rLIBudUHp/dSrd5TwLACS+Fr0PFGQSXZNaKptwCY
8D0hfLxxv5Zip0Py0Unc1hEfa89/28Bt0vidyxEllsjymFtZ949Nyp8nJ/+T0iQ3
08Aq8uumpsCDmxKDMXJPSsqsGOTAUcIWebLsTa5ZP3sRRoJuREkdk3o9Izh9EzpA
fsRnrye2WwsYdVcR+LXKTQlOWL/BtAYPzWRM1hrG73dpamC63MZesKc+pOX0yrby
QZKr3zZQ8EWsSthTFYuU1BCDobZ1zcXZWtIqH1N7HpDoqdgBFb14UwyYQKVFptd9
iQ1VfqlSPt9voJCmSQJIdSAcLM/wFnRSQJoq5GbPcQPd+PeAXKIyM7ZUk0tmsyrt
Gd+eGGkIcB8NsJdILO5E3zdAiV3MpMVk3YeAGcwHQ6z6zdTvj/LgBGc/5nJKL1Ng
Q2vJlB4+kWNl4HWreTIsadWjcUuT5g0uYmRX+chdcLtszQhM/kj6DlZLKIfDBRA/
R6d/T1f61Kx2NdiSAt6exOwIQI5fweLnhMdkbFqnNxnj3i6M1LtoJQyrH5NMaA0S
CmwT6RfDGS81QftrtpD4IRJWdk6LDzlXOXPcJAx7Rf42mozKwP5r3E/fLumH0o6I
gr5mOT1grn5HnB79Jzm1p+sJAzYTG4JjrbEUn9ZJ6ApITcrBqBxUL6RFgb3F7sku
0zo7IynLlBEOX4b1RHe2oKq/zIKX2PjnIUUNpOs6iEtGT8IsP3WA5YyvEk7AHzaa
KK/CgCPRV7vaq43uvSXBjcqp3kvlyv8M85gN9nNXfjF7Nd9TxU74bgho3XlMj6JK
WR+xn0JsqiIhpISlHCU6xyIH/yb15osQkQNOLixZzEy9mex/0y5LTzC0egSmDrG4
Jh8bo5nRxtOrxsY2I7HRbEKcuBpaeoSiT4R+jjYwfaZ821M6S6YJe7CCNZCrPQZt
KYZN7QdLKt39xAIPK5xpDnH496942816WGpFTNB/wf0H0cyXDhvYs/m/4Pvollxk
OZqgOr3VI5roegxHlcpRTm0z/8Lwkbgk7R7OCCisBna7701oOZZ3QsaV2tE7ReNK
jJ6wIEYX5PPGZ82532yWg80u3LzrEKwMDBocAZxt/SuwWY3uzJTtUgs0dTAQTDeH
6iTm1sFAxR3Rqm4J76x36lX6G/GLWhXvUglcURQJo4rQZLddNe9mUMnMKDePDhSy
s4vQ45iyJ5wf4He6alzgyK4YuOpYAdhWo4gPSfWC0YQEOkltbUhI/YgCg+TWH7X5
ggAIvo4dYwEZw+9DZAIYXASRVdGPkn06CZv1+hZmY6RhJK4CP7TvLN44iQGkflgM
5Eg3vSKBPA9mLx4KYV/ids3TeDLXn9l1ZXBDOiGOpr3DLt7QmY/solV5UM9YPsl/
sxV9ovm5wgr8beUquER8oWybxb0Sv1JBAUSnahre1176w4W6UW39/4w+DqkrAgzx
itsKVuYuz2R8Ybjpsw4Ec2fIPW2Xq9eTmGD+Jt2TWsIQGnG683Ud/68Gk8dCqZQ7
PZfh1/PVRw8d7czl6QRR4s9/KGd/xWP8eihjmaz5uFWf0BSdBH0g+bi4okb2vRWi
91PUIyxHoMpDt4ckuy2pdHkbfXR2k1wU8myzzWeYpcsirhamR7Z6mWQuMmbH2vZ9
yIb48Eukn6LB4QrolWJC4larAYMl0G3/39tZ2kAOgMZuXOHouvHzXXIJpq/KYFTh
oWRHkJuS/6m1kUSmjEtkwPK9ViS6z1uY1War5/QsEAuQ34WQVX5+D5Ck+M4tve+6
rRt5XI8KD56mKt6Z9Maa1MlZ7fEjT6k6g2Ir+r7YDuC2Ph9lBeKsJRlm0aIYSHfH
sDnvjpqSZSk3hLOFcoEEu0w04K+WO8Jcy/zBra9bOcEyLQGqrR40aG0tRCimH6Gy
g28yaa5NCxzPrXr+CSJRrYCtrSf6IioAiwIV+K1G1dl/38m4IR4Opqr1q0Wky4is
7Vc6XuhHEBejlkoooja0Y+8UFo56Da7mEQT2SNXf5i/77JsJJp/cYpUYqFT0Q+4P
CMRs8xyaCvJ7IPrmbgMhLxV4xHIYq2trYbZX8JKZ5VqoQsZnUJkb+UKHbzIFi38w
cesRdiA3iR+d5NaTRuop2JYvhdY8Bmxz/cQPCaWyiB2iXfkE5z4PE59whG0FluCl
wPDpykjfmnBjfA7prua2wngvdDS2PagfhdPdgA3yWOZmlEBTcaIQ1rwP+gFNcCoL
EfKAFLyxRuAccpm8KQ50Yg74fSeN/7/n8MVNQ8NjV5yNoKHvnzeMf3XOtoKCqzEZ
sx/+IvFnat/AAU9eH79N9kT2G2ZTegSDI3S2/oDoyaJL9tC5bzZ8VlZWUbPH0n2K
OKLvUqb9jasgJfRIHBsyz5Dq082T5YNagKNBkP0ZFVvL7gOH7HhjS7vUJ9/d38xp
gLD+I5CT7YYGsrSSECKxLtE1o9P2AMGAiTl/q6gXEKHvjPXbxhCTWNyn7s0Z2d/I
nov6Z8P2yAN39AgVl+ruulRQH0i6B+S42QQz+KdFrXOPcwT3Q4MrFdKZ0BPU56J3
4ZvDYehhDmFKgAJ41sjLNRscwRhzeMCYab2o2i6jJ+FovGHjC9RxerHlRXnydwpU
JoZ9Xie36fJU5zfL8QzAzrLklA/lahej1ph+QQcYj2VnKsRUpGP4y5VL9JbnWMZT
nHsh899b2s4a0T5ub7MZwD0Qf28dDBpuPmedpdCfkGKXKIUfS/0p3/yvSbqeuovE
XWidd0vuAPa5Xr7Gy5vjT/wwELgZIYyJejnrVjPfSvVGWdSQnJ82rWShYolLywD5
q0uRkvkgT7+v483u6tjRsQWn8g27+JKcOoIps6tD+s8qrFnOOm6R3/RYj+PbaEhX
rPtrEy/ucDpPtpQuZR/QOGpBbK4aX+HEm5xcZqkNUPZTyas4JN+yHg5ppJVMRpIQ
9EaVbASHUmllDEOf+e/y5i85VPgjIffQ92kv32iw+03IOiCxNL2798KNyZqFgpdc
Dh8HQIm8dUDn7zesmXzIuAVt+MrErBSLIqfkHTIQFBpBDTy41aQwmEpze/qAlcnf
0pdiy9S3IlgLEFLpZrneEHMHhhNmiii5Uky+5q2DoR3ZrHs1Aaw/6jR/sXdfYXXN
H/cpSOaH/NGdDtpbXhXpb8fJzIR+SANShX/i7IlaBYTHQLim12RSYM3MGv4lw7bl
y0DjAnhVipRf6A7UBrtXaSOmjDbR1/teF5nD7PkEtnNWjTf5UOkj52YOZzxMAIep
WB/TBL691QeJw8TcO95bNlWnhpirpEKPVYkw8SI8Ibt0MXQRjEhBJRU6bN6xX/OY
i8dppa9JNOsA5NKQa/PIaWvnr7IoeG9UHG5KpC6ru84Wzvf1rKmgXR2x/IKwIljK
T6nonQ8iSdPYfcXTxljh6I5m5fZcOwb1ctXoxl8Xt9Id7zdoqppGqHCJuShy5v1X
lbhzA3ByT2s/vtC5bWKfE9EV5KaZ4whXyMlqcHM3z67R25SdD4Cgv1WPL6O/hGrj
xuoo7TZmq/9l5ZlN9PYwcI1Bu3DnJYN9MxyURdp/g2eNAPwc272Y5V+0StRIiLp7
cTeR9rGsM7NFmYr6+5EUsp42MdQGwyRHlA99qbark1bfjd8CvzcuYG2QjvfqS4RR
+YG1JR8LrLO/IhzuMldrNQh81TA5cV7zp4sjaI4cJlo8K3Ee9ve0kQazg1Zjjwki
9prOjzVNk7iW+FanNWJwV1YAYEz2m7HktdmazmNwyxJdFrv3eAyn08ibMfsSo2ga
Tfs2q62IwnNWlW+5mtEZSzBdSe0hVgEviR/N+gYtTpSTNO16cmaMP3pinbmbo/Tv
lXCK+UIQaMePX8/1JNNH+kc1ypl7UME3iFbFmbz+ZKtiFRyM6ccyaAbRAXEV73Kp
v1LqshdJquc9spXR2xzSaSDauMwnhc/8zJ2UmKra7JZ5lRXe7v/j4/O8DZ7PFPWa
MAZpL1i7iY/mmJZxZqmSbSljgpf1s6hDC7EYu2J3DhXtYKMMNCb5HzpaUsmyvMyT
h+oenlWvVc7C3r74mlNfkNUdNdiqWbarMvfmddkcMws5WTL96YUTJG1V+om0go6V
PTcG9NuE47y8jJK9Soci8d3oDjtKmzSLMFwYYn2lkUpkhqslVCic5qhArMu4H6mb
pSszC8T8fULkkaxAnY/d+9Vyr+nl+nOIsIom90UHODWAjxfVnF8WB2jvrXVrARC1
mOHPPAWYvw5IzexyHTtpVGhOsQal+Z82hB0iGYW8gzOsjKx2EBUH6pFYRdk0aKd8
6VTt5erF6AOsZNyCjC69lCWwglLuiOgomI3uDvwI//33DuM5LqCcB/lSZMTKJ9y0
bItvt1/V2iFTf+iTGoot1vj2mN41AqfMgZ05RoGMCQXH020fOLQhWyA98q6xJ/9T
yBkN4pDKe+t521sUUFQGxmAe5PhWkagqrEgNjniU3jgYLrDMPaNXy2xKEah4T+hn
ZfoTwCQNR+Sjninps55M8iLhtVhH8s/O90dMpnAaEKvTLJrkO7CyYBUWHQGOTF9N
HUiTg95/IItqGb7BC/VYKT/IVjPskUDZOObXk2gxrrYQct3tAiuCPmhjL1zIZQWR
ThcJdukNDK9JvHiEsmyn64pgzyVR5wt4UMzZTHfvDcEztVJzTEwIcPTpxh2squgL
uSw22tNDmmV2KclsaonUEyFdGcI8qme/JFB+rOUB34Q6AIw13iZdMBRPcN209D8l
FmrPwdjqRNdRt4UsCcXgTiV8iHqO84TjyCCz2cbdBl3ukhh+MhNN6pPh844eFONK
0Pj7T/bvI2sivryCBrsbTa6HJpmc360sF/flUGnDZIQEtI4lt/JeNswcCRAYyHL6
/4uOICiIrrXOELRHOD9z0FYchAUV0m8D22C8mdTAHF5J2k+KhKdvsOe/j7DzxEry
Zl9NjAYGEMQJt4CZpGBroi63JlREjuaoSyYPfk3zuHELF+lxuF5l7jdVbGYnv5HV
b/wfmbxa3gewg27+Nw3XNQF1mHUD2AZr8sjyfk74P5NWPBG3lH3fvkrrSIAnt238
ds5ZqiQZxzLoeham24lpbBsSkFEv8vbREp2/kfztCr6MCdTdemf3kPS26j/bPxlP
zOqT8wEaim9VHgcM9wXv8HoR0zKyCqBEfHYGemICV/oWYnePPgE3TtYc/eHMJHHm
BjWNBCuS9fhA9EngaA0nu/eBjBdL1hDGiMXJgfojoiNfHAkN0prqDdw3ep0m3msy
yFwMHUIUIo+pwHfX/JaH56kZk3i0yg+yP9iXUs4/fVLrgqiSJSjr9pL1pJMJ2q+T
IA+NCntv4MYVEVD9sdNBP0vc29W8aGyoPeJ/j1zsnLjqHdLz7RK+WMhsgg9L5mvX
kRgVS9WGGe5ctr6FfDtnXAwK63Sn7gjPmh+gDXyWs+UE8w+N4ZsxDiHpyQl/toCy
yelUUIu8MUnDfyXQdhf7u0IWslydzagkxZbXGslUB0JPD5CQSOCdKpzU7JWFppWV
Hq0ETzVtKT6ARoz/fUQegK8nPAyggyv9q2IjjAQgtZIdQzv73ogrAAXl8QmhcqP0
q24LOIr1XPOd4/Cnbk9M4VJ7CLg4xugCcYqtgR3IZOpmXssESAMctpRHlOmbtVtV
vMtYtRrDcEmnt/+MXCxHnZmD74Y9XCrYaPfGOe+2ve7nIN8NJ+5j4sLODcYX9uoJ
zNDJUj+iFHFWWVBY/0VNaGIhayWgPDSvzKLkK7NtRGF+cNE22BdrwOqiBfIe4Fvo
6JoKsLtvHXq69PunZKxaQuXD4dT30DvqE1K5cHggacgtwbezrBlUC08FMREelN3o
kHJLzvTkfUQ7q19zhMQA2WF2ucnoppRJxFT5z6dPJbGcEu2uPdbtcHxuFREUMp2x
Yc3xTBm/Qm5bMeMzB6Qx0339PvzKZ2RqS+64duWBjTwBs08Evgphy3h0ktepnxHd
+7/YG9UkCZ8yC+VieS20vT7ZPTQbCecFhF6UjG5wM9L+TXrRxqXSd/QmVBkY0NO6
sfZTjw0wxHKmdh9PUfutpgwoJC1sH7pK0XGNok9esVzUty+MR7WbJ2RrwlO6/g37
8jfo397S7wnfouwgtOkHNbHjStGajY9MOG6MsJmEOeBfXnu6GAd4vzDG5vyb9ROG
EiOFlHB2FalwNgZgrjA6cXtZhjbsPF1ZZC855on78Mggp07RBaUTdi2PzeAa7BvD
h70w7NnpCW+9IwvEEKjWySJzEo0O7nOAoJcgw2LHLnHlzBP9po2bPmLGeFsUemMe
RjzvADf/5K0uSOW0YwJWxKpbs422exk4IENJvdPdmU112EzhKEoWRtDD1XNmn19T
kaAsSEH4fUM1OuDCjL+bORnmcZtF9TY7WWdrCOWhs9/Ku+bhYNopd3ZEJFI3k7dr
miBl2CJxhKGVTCA9iRn5WsV/X9VjyVXJ6uFs3GugYc9HKF3GBNEZCkxe9JW/bbg5
cDGF3+TBWsKURyz8Mr5a22AZUkpbAUCvojtfNcbZjfpA9VQIOsJJLO9GqFbfM6U+
d4aOhdFdK6eXlBRtquhZUWiufscrOhkIItyYnIMg17Dvn40h7n99M2LwIV3RKhe+
H2A6zyYlw0jX/YecMePKinDYgLoFtT9/W4G2fpgIsqbzbXS1skH+s9VkKXd2Frao
qfyrHyf4Hbe6CalRQqwIA1weF78G6MENrXW/iklv021jKix3VcCrOo9xb33aATk+
mGZdIdP0wFviKsSb/aCwbK3QT5g6ZvHOR4Wcig49uTL/wxLeL2Zw3yfHivdVThIe
X0vGIvzdHLrrEuo4U2kdYBLiGxasfscoPGmDWdfuubhVi7MQ0WCg33rFU1X/qDIi
coRt6eCdPpiNVB0w1kdcxqBz3zn9rZy/I93A4GFTqV/5yNRCQGy2w/rKOcEoQslq
9gqt0hpzwvek64llIjyN2oqIq5nE9OKYBQZvLKps7A5Dc8PLXseWbeP68Df7dHuG
Lpx8RygEfELkqdA+HnNc2iyVu4K0OkAlkBxUM+7r5OrnY8cEXiKlN8CwZtE7AvoR
Ixbpc9Yv0ueaaWP3OGjRtQHh67TnLqQTyM3WaAGdDwMEgL0Vmc0IAJUUwAdfO2aq
iAhCn/0rvLszOZi/upCKJCmfR7VgUTHygT3Jj2lK6+rwPBEbKv51vNww9u/yTwZd
LhxTl/oqlHKennWoS+o0w01OHXXXw4uUYgZYT2Ws0FsLhrDb3h+F6muRNtOV+4OW
6QQm/i7FuGsTUSYeC6klHGaZH80s5ERSsrztReZqNpF8vuZucR1NfqUZBHoHbCzr
pc5WpA8Lq3RxHA7zv5xYyGoE8AxgT32aQM/c+c/1p6G3nahDQrxfx7e20F8DpAqp
GdRv7V2sSmqp0CvOux0k5Ghqw3rsAKtvi9SuAEIb5ZZH2Z9y9yRnUtpZPyoXa+WF
tHMp5GyaSo4Ere1KE2R/WRkxuzXKeVjRtHD05yRt8WYac0HAtsYzb+kQPKKwBTnQ
MpVX6qMyq4ANXrTXx46G56upAj8Ms4iJZGA7H7XaDPZamkAq7isyuk+vN9sTwH9f
KgYYHd+19L8CO7/5Rv2MXjIIyYVcxmZcmgQ0hkLS800X2PUNn2UEp2anHKn7Y3oo
eA/cVvVj+tEsBBRVWER/2p3OgZr8l4kVBfgWCnVE011g6fRvUZvmYr3jQ5yJvwtQ
dUSIhkKaSH5iRRiflg+Orwb4+9M8h+vfm+HjoIb1Pbgvunt/wHvU3kfzro1TsW7G
rjHDzL6B4CIU1w/LGTSgmz5iEeRVV2DeT4vBycuB3nWCgIG0AxEfERmktCpNfuxT
z9XqMJ4BENaqqFoVLmsdF+whnk+1dNUmrSdqsp8zb6Q6pwaDb5cjfGD7182FKb3n
ssR6CmH+GPm2nfATEDnUWJgZemX8TNrbp4fgtoEredZ0v8JgQRaP5MIAQbpIPA5b
3kLSBbU+LoB5eCzSrizwBoGTZ71KG+99pc10Pl+bltlkwOJZW1qgolC7UqXwin0c
rrIRXXIQ6ULXiv7dRhLr4hFAF9x/Xl/4M+qZgp/iYjVmzErOvXZRPBqlvK1BwgYT
pKana7g3xpjrc2UMf6P2MeAvHIGpipOe4Ck37by3JP9zmfmDIrM9ivEHCspnezsS
qVI5wWtqENtnG1EEQG5bh7+V8f5pSfC7gx/AflH8dObBUopNxkBMvajPiA8tQlX9
fTszOdKDne9TrOSzXP1VThfTLCe+RQnQDUZ+cfNJAIl6f/GNmeIhwUGJgJjkkrSL
AUxSihsgHKoGADPo9gxVteq2DFeTDg2XzvjX6sKj8zq0yU996nqQhM7Sd9yYmJVT
rHkxIBQkUIgXldHMWCJXz7J9TdGPal6tuLiQw2SAvtYvZKOtfPop6JxsOt6Cg7t0
T2hN7zVatA9KnqaBbRwo0+ZHKGPPFfsHvHYMAYEcY0I0oVI9kiZ/HF4m/p/WM6O9
QwgdIC1wuKKPJOsvvuow4hCIbmhC9gpxMyMomaKd+31p8AXzpGt3YQLOZoBHsY+K
pBmA79S4kFT04k4OiIKKB9dAzyZudJ/IikMR4XZTnQaEW2ZE8bBUJX10SI/zFZml
CM4tQmC45vIBRsXLAUS7+3i/+3egQceVVzoTFX8PdvExuCUdO/UI2Eo7v+xCA3ws
a4Q6o3Se4mDrpgHQXxbip5Z/042RdHqrFYaoz6yeelb6gWH78PLFGhJVuLaeSic8
ZMM8PFND20qFQTT/DHl0Um2MIqbY/71SlXWLC5NhyUpiqgFrFVhvTvKoy9OXT1zV
BLDzA0M+O8jYMQXsioySTEeLfWmaACWSq0HEMWOXxl2rY/4G4c2lmAw0TSzTz/h7
DptZ9O3Rkbb02Fd/szCPIkraJCD4JKWsomPxUtLv1fAKJ8aJUSOBoH2oT7nYvOQN
+/7xAeId5052kNYyiM23syya/v7AEPdH8vY6jQhMjORIXBPK3LEQrE4s/OO77Zu5
0LcqWV1jFjvFo+Ffci+D4tM8fAPaCq3WlMhTfbQMutHj72+QciH/l8+trlBIP88F
3ETt1y3qBjIVo+dMu5KhmSTc6AhhlHm6tsBZ7Frl9nRmd8+bPP73GZANy/OHiqsk
0mZc910/dva20kmhxv3gtDfVS/StELP47RheQI5qVpax6m/kARHotASKDsX12Pfy
i4+gHhYHZ9Eiw+rMxGOFKZuPDpg3LC8pbxRx3hVVhsxu1cHsAQBbUbAPvLPCEwil
5yWiIVwnAcs7aycUoCAa5JjdphGK8lvfF/04vYblsNOkghlieX/nkg4RxSTs35M0
TQBieDkT8gMQLutvflHjXk5NQRxCMd6mtY6QFctsa4Ybj+VMG5gIURML2Y+qUcf1
tfRnHOTeGkUZG1NsCCksImN+eyzFqDLxec5TIXwnxNpEWfzZNNh5u/+TKG5UJNXh
Go6JR3kt+yENlfBj24XLo4vOjnryQMmWA6jcZCjeeD6WouOmZBCjpGnhSmNWcql4
f5tKWrBzwFTQbBqNzH6LjVgVhC1jr7xW7WyoGE9hLvMXuBBNPxfb3u7fIqvkiVRu
bnAEGB1ytRPycR/AwrXY+SGTMTprLmPxhOQVREQ4GtFaJVyxUztTM+Q/gmz/C/2S
19xi7u4R5jeDL23sAtjP9LXBEtx2vQkcyaGqaSpRvMIdD2hWrzQ9MOGggig2e2zF
4pQP5rVFBMuVJLAY00oagn50jzaWNq+dgqZxESMYFSCa+YpL3NHjoouGOWWosC3N
HmKyr9FNdJ7JbQlqD074zHVo7UgloR/hBkYvrRXaiRIm924JMfD+6l3qPALVFRQD
lkLsg8oV7dcogKVm4DYMwO8Nx86e3oJPRJ7boK03yA3VhvNznBw+PUavj0Rg8Sam
3PAtgzmthg7gT0Fooo8o8tZ8AiTM7i9VBfUe9+StcLFju5Ru7HOIxebQee/ZVPkZ
ViBd52o+9y+7eVFAVtcYueTSooDTx6Dy8i0DzN0yhsOTQU2NN2tHvgUagdyzOP16
K+oo2bewSyQyr5YORBMrz8EustbU4q18EYcYDsUYup/LRk2t5T3c6h4f5ZkAUb1E
wR6fXMv4tZlAmvjexs0JKWQXsZa7STrFh1YT/x5zp9xUQPWPyA/KXncehhtDIGpT
d4l4NcB15rpsajCnyvTSE41m6TFsFYLLYs5RTa9pa9vyFuWT/FkHbx8ne/SjP3cW
r9aquy7SzeduTLJbXWx60z/b3/EdmRJMtpLisAoX3g1bs3kQEFTevhl5mQQtBD/r
gEkO0Z+KDqI58hG5rx15qWsVRCs/AphDLGnGXTrrxIiqvd0uZM6SK9CpGtGqO3sp
L+9RQw6pBq5VuakGrV6P6CCUj4TqyD2ws3ByZhlblAdjplV9870yWhzCFzXuikd4
32LOt5psV1AwxjhCZGcrSLkXnc/bwkmfOif/CzXHpcglEv4B3BlzFS2K7eh5XkQD
2/iImB399rgsK81Zhl+nbwTVVndjEzecW3BaKSBX88CSX4jbrVRmcLp+d3uS6dx7
Nn/g4jHS887Z2vkjCNEK+ht7yn3L+hoizmZmXfgl89n7757PJ65UNXwCnE7QWR/b
wwBpIHHeaRZL/ZsP3kwafQQTxJ6rhXKhaKPBZLwhnoraSjqtNDSG02Jrk1kJu04s
xQSDRNPrVCdlyDRpmZYSH7Dx24x5ebWDN/JjH+dObcewueKsYQIWDJRV4kW6HPwi
EDM+nAm2VaZ6Qz62uT9SRiZhxdGQG7PcDSuaoS/N9OJqVlzreTf5WbAki/TI6inu
cdAU1vtTnXxnGSsj8RbayKJmB+xIRDiETWhWhOZm9cNjSgj/ouZBYbPWZdjhH8RM
koWty6t1BFisIekfzY3eeFGB/+K+dW47BfMd1r64MgiKH1m/xzVNBMxJh9+EAE86
MUdpm48f9Gy/+97qNJfA/EZVI+KDQgHf3oeqHkGTM88hAxMErVFjd5Hp/cGf9Van
8GdM/7iYOR3iFggiqg9Ke5Tk3g/WQ5wSf+j+HcRR87ZLKuNkVn85sNkGKoiA0Hfr
q4SdDejdM6aBZ0WwnGTgFK7K1WC6P77Fbdc5EjldE37YySmPKyEOtJZ7TBd6QHKg
qJM3m6lj9Qw9VDBsb4d/aSc8DBvYiiWDjULdTNLrfynb9mLHVeD+kkHre/P3uy/E
Fw9qPlEudvNzXFO+VzYx4PE3iOpWYTFk/a7xISBmAQLIm35J1L51tlR9pGwRsaVq
/Sx88OYcJCRbMiAkp4SQKSpJS210hidTOzm79ZRi2/N1ntysgncjY0TqVIcTBZS1
F3Q0R/Fd8I6IWc+YXb/MPfcMGAqpKjlptejkjqh1b0hDqofEppGz3TjwO86Z9122
DZc2ewLX4PYyp3DtpwRQ3AuKAG5JY2hbvA0/8Y7YMDHrMWbQ6V8NGhh8/o957Ww7
8Fn7WPv+hA7yBEk+y5n1OoGKs90WGCL3N5nShqb1sv3wiN/q5KrL6pM76H0Un8H8
Qunw2M4fyVT4mWks8bEsf3qqwWDW05cr+SbpjzIbM3zXe8rfsneAAreCvSAPxNhx
qn/s35lSCRQ3GHkZ+OABDcn5UaLfJJ/WZDM3RVXfXAB0sThwG21neCgLRndFCOBT
uPpzraDO38dIfM2mgZWvpKBt3dkRbvTP79RZ4dnXpJWrhAdb0fZYWBT0YtURPz0P
gXFI/QPhD2L9AiY0FmJ9A9AD1rQkgCIF/bIWRXnmDPoUjivcH1/WcER4DCui8zqt
oLKjUg6YbUQs9pa5zPlqTJ4I/hskkDWHkG8LHxaZBDrdzp4dHuLMx+a+Vsw1m3/f
wugs94laR3UcI25YDaXbJG1n05IVs+NiLVeYUT1iPVnGTuz4wUVCDnEybqmvjY3b
jD91N+CekpEmc5zP/nFW50M8Kq/Oq26k1tODUb45A9yyVo7nuSvkCqq6GWNwikkp
BbuItR2E3ApnmXft72qqabZf29N1Qo6l19ay5SbWI6Rn07svwRu8Ag1WcRB2XdcP
ySQPAijcey9sddcnsP59VDLZF3V1cxse7UGErWaI5dpiwqgpbdNGkUyj4UpMDU6J
46tPR4q9V7Gv/e6bO5x0b+JgxooxfpM/GaiASrh1E0P5M/8KXBF9g4y4b1o/oxl8
UcShtKH+ajdqnUAhVq/jQ9pltkf1EceMTt/gIfmLSuVk4x7050htGVe+TzoCEEiy
NRaOUIgZ3gyrm+URlk1uQ1gxNUF9+JRFTG4k2FZcbjMwymtRc2CxuTGynSdD4MhW
8d1LxOCm1Bb2twesGVYv42JG6gKALpX4M12IC94DB8sgpPpv9qBqnrusSHmIxYlC
hmc2Uqm62TolDVLiU/PD9upWByo4LH1248fsraKm+rvwz4vkjdWbIRcpmBk8Nl20
QP6lSY1stR1ZV/GpJ1dAS3e2FZJI0bojDuQlxwiE7lJqcZzcENt4gcZwqQnUo64G
4oVBLcjvkKHyeBDZAm3KBXw9j14vKgQG1W6XuRbZQeUO7FC/CQRuydeaCBlL0Npu
qzMrTRs+Wvdd09Tb4oTIzwiEFfxsjDLfFfwCjcHlCpqjBqtwSPklygmXcxM4zPiD
w7UPBUPIPemo3GFa8fTSDSysXahvpd9dpXr76j6xHisjGZCH5IUI4IvfmIdSRPap
3OqMvbJPeyTfTIfyLVgUTWIqHjv81ecucYPsc27X1r1G3n9Yd05pfpd12B5IFNPM
SYODcdf2rWn5wqDv+dgoO6lmN2nXlhj1BGaRv1CKzQtW12rVmFfPwhb9u9m3Mlph
AlejDtYBUHGHTioz74tpFFiDnUbqKJTVHu6oO/t8bhv2xV4bVlmK9dzON7UO9ujE
9FOGQSBGpuEr7Ke85ox+Qo7YN1+E0jBMSFiUF5AgT0Ox+KkEWITVZOawVwa2DGZq
+3i8WDewPoKIO5mEJx+GWmRuxBoB47zvkkINYqsBFDsbByQnilcxjcbIH7iMwmjn
1V1HPjq3gUAHCVB5ga8Gxx7hbe0Xnn43uBNty2jR5o4j/lVuMNWmA/2xxaSIGyFK
HtIMp6pa6D1uHhoNimVl41v2u3a2jnPv3fgJbRA3B86SunQV/kvISNz+wy/+kRGV
lHEQIA0+HqXQH2aglxx1+CCXUdtVW1oTNQbIOeQi3eEq4JIe1dJk5ZuWStJsQ9X9
IpaZWR8JMPgvq+oTcodKSVMepEVp43ELOmFCNn+8o5XDgSyfFa6/ktrsrol/nuSa
AN7ef2uyPYhAZgXUcm+IyZL55XIpd2POIe1eZAm239hau44lKlQONIuwOccjhvv4
i9ZyYC2T65lGGyznjUBAOqpBn2E+4PFaDlKfTO0GZOhOsiP2bXTm/jKVLyw+lR7o
4QYlONaM42YJ+a95Xhd5Gu1DZjtqncEt/5m7hF3l3e1QrSnob1a9FEklf64gpnHM
PorVcpMgdLuMr3l6XbOpcbkFwxdcWLN71HZJtbbV83ohar5WFclgliU7JUTeSoT2
kMvcNEGYJ6EyJ4+ysRZ/G4VzKNEDmWuZmGFkIc8nV6UkB2x54baY0bsAyfypUIJM
t0B+Uz/ES7uQop4Il0o/ECcJmyAFPX6uDR0TDH7AaTT1DsRWYEbfnxvvmAf530qB
c4f8Y3bgPcr3U0YIY+cAFeNRZcRETOsbFQuiV3sovKfB1cgpuap/bsEQUnQ3Gs26
Gg7edLM1ByraxOI0kj34Zs+thnnQzY/7Hh1QpDKlaSgCzNUUjNJWDUS+L3azG1Tc
EpmMfJ/jqd1BZBCV+lDTzYFalw0u+pnXhwgnEH4MWoV7HlO6mbc1COoTsPhNkiHf
YBQs0PC97w2f+KyZ2kO0wmK/lubMt7LatMw1O82C/fJx6S9+J/XLxPDEKjYb/Le/
dEagJJ6c+564GvUt0W8e4VJCIBBXat59AAcumE/i6v2zdAFerFGkuB2si9HO7lT+
qNEGsaOHd09y59yDhTAfyH3PjJ/4kToEgQ680FaZOWJfmeN7LyXM3bqlEK+JLGIG
yAEsWcZ73Hm/g4XFICOnJfH6Xs3QldmMUF6DbWA6s9Ls/qomQj0nVgD7bO56CE/c
ANAyoeFfXmkThrtkD9Iu9g6S9Pa27WNI4oqAkBDpR3AAEx7kWVeQEkex/O6e5uda
nZGdR14bYDb2N2elZAW087JZjUwFnlsED3q+/hyK067XmP5fq6t+NgUKqgBEDEQs
AFCINUQyvmAsSIuLgkcfVW1i1hNoPabv7He/ho0DEAKRyxJNhuWiEIyy+SWoOr4w
aRMa7G8uqjog252xidE4x8O+3fr0uiYAooJT7xUPpmjjJNxN6xmNufYKOe4mmzJ7
q7/NdZn3BtE9lWwBzDb62LZChCSzoj602a/LUT5R2R/heFmzr7Gsg6wqBDgTE2wh
YjgecpwyHkFIg7YauOu7v2Z0to+IyOPnZvIw7ruDvrVPJyzIjN6xxqqmWlItzuRi
bSxgBcZqrg06TQ0TcGGSRVMHuIXFRGtDtM4KXL5Vz/OqZLXOvzrUeuLWO6ieuc7j
rLswliuUaELTlYNwnibv3iOCYyLs+sqo+Qz4o/PXKeL36VYZvVeJ8yiY4aWqNvLH
R/YDESRKruAN+m/6aNCitzFLQAurto1sxcKHfVD8Yr5SyHldiBAQwDEXlLCjJ4Z5
yJ/38xQnmE8zxCopGOjv0jtie3CuHj+/SgKPbwX3SCLaM9eHv9lNJt5zfHVhltG2
giVIZt3lwMFJe9R6d3G5DCZS6t0f/uAtBh3dekTzLjIDz/kAQMpdjqwtIGxFsgd9
PcDIaxfmMbUsdv3e8nJY9hdDUK/C6Rz7qPaFc8+QY1pbgz3O8iHm4htjNJ0wmSwv
1BHw/IRpf4mHuoFKDxzVFxzWa2JQuzZt1uHBlUm1IDF6VhfKkcERmhLSOFFi4wnJ
jWqrDzJokT4rkLdyoNna1IEO5TORl9O9Bn1LJ3/enp9hOc4enwOVJTXRQc44CCRC
7LJLc8VHSUH7rQyfLOAvaDkxyiLhJwx9rZ+0Fi/pyLTGv3uUvTWnclzNsEjO8yXL
fO2q2iYsKdOxb+rJ1acQLXg29QF25lkJniX0P9JC+TwwdT5cjZLYAsTjUzgPwhB+
0rJSu3WRHlHquTnLcscwLneiWgpDToO25Y78RhJ3FuzU6c8MZqmjIig0AOLYRhi0
5IoCLPwEsPbSLO8eCvwCMkmzw48XoY6y8zRHKpDcIKP20Wg5ubBH4ATOQ3l8q9qf
xBxxPP7w/9sKQZpJ5eIISpO1xBds45Ad9Yy6LcGuWjOP4quPyxMJ8eHjwaaC/xlD
O8N8Ok5+9iSB9sbFkk2wLK0yjBj/3VtI019I36u9Cmy8gIGbGI02xxbumbJgxUe9
mk7YKvThKcaP40E/ivcRZYQNNn+HEUGonJRcsXUhXqeVnDsD8t76lJBGlY+sxWKr
bmIvUmPMpKlae/0YyisUdOE/l2K8y7yJMY5JqfQMdIQD8FtVPg4Vc4JlYc21mZux
EfmqpvjxQGdko8ppetwms3jTXvXLB5gGc3Feyx1polbE4gBAcr5MvxPGqsSMopYg
TzxJGgfzQ69ashf1DvnYW65h7GKuTpMe1ez2tjFPDKO1Y4R+MJsH5yMNGI4Vc7Hk
GETRSPS79WX5BYJO1kv4cQ70MrNfVo+q4vQcrdP1Hgp23wpIH/Glww7Nw0yaJI+L
tlTNznGbS7/KIlW3NLqcI5pdakOrr9runW/nvEXxwbsEOtigi12ctLIRNGBLgB0g
l4PiAnaEDfCb/2mXEVNptsI+6njMPwowgyK/ki9XKqp7CTGk49XixGFw1u/IKuEu
s14Su0gK/AadM0M7DGOuyjpFu04DuOpytd3b0YzNeJIBfC3ZGvote6BAdrlQqA2Q
kC9QBGKY+qhhkHO518r82wYxoibotA2S86hGZIgkh3W8y7u2UM8RdVZb8mVGjWV8
sllA1yzfXpx2GAY1u5FKRVeZxGKLxR3ueRkyVtnNlwq+VhOCRZkaMo2HFNoRMzLF
h7w03LmkYRqFPa8PXgR9Ktk80M4OlXDQ0fgU+B2sUxf/5SF7FTBaiYMl6keaCymp
IfkBsn1M0yucKgp+eDKA8PBMjWjA/deUm6ObczCs1Vra0/Ci/LmN6vvKkNOKyse2
tF3jcQAxS5Qtuk+VMfHkvl3knMwoNwX+UIR0+HDYhYP6o5w+GrXWTl6G4ZvH+LzP
rhFryV4+iFI0Ao6mIm37tfq57RYLkQYZjAdATnGNKnIc5NLwRYfPrKywk5HGzDo7
iSPPCjjfLMhFVLR5QCNN8Hqg6C7QDucnYz/M1acpjs/l+ox9c/F4qRn00iNejqwM
Po7Gzh1CgWcf3zyZbITMx16mJU8BtpNnPSeHkUbT+u2MPNogldJzMPRK/DDO1vhv
/+80uO2WN9NZWKeBevstGvwczh5VwUYqDWR5mgAtTxG97KnU/GF38j719bKS/glk
v3Wyali62gGam5KICsRgv6c9T2liYBmC9LgzOP2MsVr+R26M6q7L82Y55NXAQlqV
q13OueIvQdElDOdrGMo1THBTel7APAHMmF+o0D0oyn8MEaCR46TF1T6fFEUFSBsu
WgcmDh54lZcADSl2a/9K6UFLmBy2M5LIwhSJ9ALK1K2zT6IOVWn/DEpYx/54gBdy
7l6GS/1OqQlV8tLY1fso9vdlhQ5LW5erk2Zk63iLN5rW6j2AWMoiagwlnVEtn2yV
38X4Sy2VrPEX3qLa65zn331PtYzv7AE2JrWqDV03s02XwbGwZ/iK2ps3s1jG40AY
TrFrQ6QQz1YycRMJS29rUcjpst4XZ0SPFcxb3oOLM3WlkZj9dghyYFoMT4MzRp6k
f8mRAafyodNieZ5nfHjM/1fkN7TanKzmx4g+pJj14DgKLgCTzf8Ag3M6Zv0utPIF
PljbcqnzyEugaWzGyrQJfCt/dpC8JuGrUwQLP+Z4p5ayXO50/FgJvL6H0p+Vms8z
XNjA0TdXINkeMidxMozcrk7ogRNu8L1ygZ1HDKDQqIYjh3u4Z3m/0irVcieSN2Fy
xclOwFYxEG9ojPeSsi467ZJYbLsMOBsiEL0n7sntN8z0i16H/MUL2EqX8tWfcXTo
yp7EM+g9JO0QPVVZLUM8xPg+xsv+RgmCTQr8rNyCwjuJBoML427rYXebTWHeHb5k
vKW0nHulRdjaxHZiVDb9q+TrtAL+QxZrvJvUJ52genibOtO+UAsw907CSfM0bBRf
SP4+Qm7fDEVb0wGSozI7EwdWcygdqORxpvoF+n5xI4mMRmAKB+GzudoGx8idPXrY
AYw38seyHP3PkHmzEG2WEUuKnpnLm9pgcenxTO1k4TGd66IbPu25TaYn7rs8UVKz
dUyqKq6VzpFldNUeJt7FzPxSPuT94ute5NftaNB6GQ0Qkb43oad5sAv5dRb9tBlZ
H25W+VQfky4RSH++v8r2SsG147PT2aml7MfO9YeWtZqVcNTejAwHqtqjpCaI0MsY
MELay1EAduNhJCg52haj5qpTnTYNaluCE2peBrCtwFi9XINWlWNH9FLu1gf5FJrx
Z8gNg9Q+yXZ1ZoI1jW+DDcGuIXfv1LLhjkPPKIKzY7sPflDrR1lxG9ZfNuf2613W
Waq8FS4k+EuKq4oOS+UqO3CD+8GLB9/QwH/BXTLG4s3YrimC9RBw2tDIwwhF6oaj
NyW5GXuYoXmqK/aP+jqK2h48bDwD10KKW7zbGwuGu/2yvGywo4dRFce/37NmRbLH
DDrobxijtbrKXNRi380idckYTka01CLaCdnnMiFOH9tV+DQtQFhdNcDTa/dZS+om
1puwdj35nMsYSo+12UzHODqJhX59nqDEMY7ZicJSWpbK+b7XGTm1V5MBaHIvpEpj
iZ0B0CJ0YoL6rqGXQsayjfwriEKEtfuDiZhSZejhUciSx7vizZrN6yWNBwrdLIpB
tsDCvNZM5DBISfjp0X+gspYTZPDOPbUBoTgJHqjZUsW8IWg5KrhuWkYVZlwvUwRE
OVf8C94eSVc6980Bp6FM7ZVen5WRKJZBiRWFMw8dhkDmifFzjZXXVmjoVEvppFYU
/nvD5frKjcjkR6CFSvyV9kRXDKulZNtTqFiNy2VQZfmjzm4o7Uhog/9WshGqK8aO
UTsqKwPo1ky7r6nQy8Qwtg8uZ4KjF4cnHpIBgQOU5IV27DVhew+hw3XA6QqK/UzU
kPJWY3SW+0xAHzUWsI9haEJ4HfkgE5VixPOp39/32SEIEO7F2r0OI3KoysqwlAZX
yX0hPyahf41Vc1Rgi5bg3ppC16F+KnZn8Z5LoiSeO+XVoKwupIKYXtKCq4z1pKy9
UVapWHG+3eym3emCoR9wwShCANVNSXlLJrysmRx4hutGJz4bZQXmpPdOLBGJ9F8k
e4isGDYDJEyiqJFlcfTa3nKCcLwf4iP8iXq6xO7K+pFcCUC6anl1UD1N0SUjMOZS
ljszOgifOpVD6IB2p9u0WRtN/7qIy5AcN1bsqy5RdBlLviortHIHwNZIWKIyEz24
b+oGBmuZhz+T6wrUtW8DUQUQTZysERBNLcVoHs4Elml/SOPlLFFhnNd5CjT9VAyU
RkCLHxbxCiRPFMG5WudVxGgCIIkEmwZFOouCZ0UY2VsCqGXCPH5/FraapEjAGljx
j+e/hhUs0SNIU3e0l4FjHp8uJT90Kj771FagUJx6Rq+xclYfbsKNxXGL67cciqjr
oZMlzS84HtqnZxsF4ytAceKmpggoNTut6iZ7CdIC2mjT17hzEhwm+DoVqNtgqued
pN0Vws2e419E2FVA4Wl9GtF66FrQqRYsHqhIkmfE4X1xPZ7KP+PbFF8suMJVdQJr
lIyrfos+uAffIpZ+m2H3NPHBkl9r5XPOm0Ro5cADJ8sQtdV7LvoirkMpbLw0cXiy
UXh16mIJYq+X9y9SqGqiAKVoH3SpQHr0QZphdf4c6YcNwLaAqkLfPBWK0eEbsBNj
gZYFr49tBGyMvY/fSaJ/UxnsmsLaEl3HYmA2Gpgcx2lUyGj7tiXtQyiONUBoJKOZ
H0fhZ0fa+xjGR2Acp75EGpg6gLz6/ebO9Bi0zfFFd9eAVbaciNfL3fAkvWPrtzWE
u8n9Bq7BWwNuMQUpgdHHyxNbOxGMAqbvtQeKzO/gE49VYqWl4/01ZU1g9xWiTeO4
X3mcW+2Bvk0KrjQ64mJtNdmtYna3mDJNQp531f+Jct8AnshcYCEKp8mMch5wwWs8
iiaqAelJpYfgCXpaaPUFoEskJYixei3vlrxh93kyjOJXFKp4ioFegmcMF6SPw3zy
6/B3IRoyk3T1qt+ywMCBoytfbjUKR0kIhhdbE4SQLkF5/YLlsn2kPghCLAgSJbx8
rc3ttxGTKuolG5viWf8NKEAnvzn/7+NixTLgxuWbWNVHrCmObwZ+D1iDRA7zwxu7
/2GyVFw1QRvnPOUWHlPvnWm429QRgLOgAor0Duf0fX4Zp8E2r04UBwUOvtrs93b7
OPbgIjzgw5mfttYrQxvnPrMXzi+mp/whC/dcd+i+io6k33gYSLak4HkHKbefYj9o
jvlLc+Maoejkl0ZuwFJ7253S8K6EOOE/8ysG5cUwrKqaBCwsB+idI6MyERr90tYv
KWECxPlNlXLxMEFi9oCC++9jofxik0GTfWBoIzncZan1XHwr9NZO0CYmPQw1EutV
lzhUVX5Fw5NXfX2GiyQgV18RXlxyJpMqJubxrzznKuOeXTQYuitAgoZ1RsOMooRZ
nBjBx//jDTFos84s8LdAKxcjBm4lvp6zdYloT+4eyth9kZAaIy+ALw1CeQJI5omE
MckUEZF+w64vJ9x02uDnTsTNV7Dka9Q4WJAN4dzS287xdzGKeI7SayonwkpPaibN
gJnhWx6rnNv3otTC3hOtZDcaHbyzE2ft1YKNm1Pg7D66UgQi2jt+4XF5CPMGVTvW
KiaWTbPKpVHGbYqE4Bw1wyL7ESGS9/egyS+km/FV+K/KUd+5L6TI7d1ewSP5bdO5
AnqmMJsLLQgMqLcWfj9h6NHujoeTrzwABUSdd6d1alQzhiMc1VqL29LDcThmQO7N
TIYBHZm4bqnMD95tx/W9TtYGixhJ/m0FPrX9Q8O1vCqBz7BgCjA/ZLOb+/YPpSSR
yaHe3xRuNwjS6k6h8eYXigIexCLzhN8pCMepj/nEXQdZ/eKlbEEKsZl/bhzLwbKT
leqcq5srKhUP1Yth6jLzPUd+qZet/LTkTAZIQ7OzrHr3MJCCVFQE2GQ/Nw1xd+Fb
S3B2BJvVCih9tBr/0TIbPtqdZZqWJsO9eTFEGOFQvKIAsI8FnXEi56TFHMAwSh9R
Xd43eORrNFCSqR+Bs6gXwmzskoknjj5hKZGVShUqxRc7Yp8KR7NPZOhQgzXVGFon
q2p54PqazvqUkC8XUgeXfcOJuZmLSJ1pJZT/iRihpN4UwGMP1RuvhNsl0SkgqBhF
tqGBM2EpkEYz76eBi6G+AcNyjyeudiEOshJA1gTkkMHkFyX/sI459oUTxqu6amiR
BiqQugRlpIL0V0kU3SXDeHQuQzomcOF8rDrMEK4PTpyAneYgNbJhZOp8U8ue89Dh
riyVM+kSuyWunFFM15CcF59f9d/9wj4ATCSwTH7/HOdmpmzsAqUplEZH7CB+ANOE
CCTp6wQSWanW96KbndMImdPBjXtxFXcr3FRxPWuHJwq0dfbGlnMepQQ6AO16hSo7
FA8SSDvXNFoGJlBjEeK8Q36eBY/44yWQdnuLzqUiLyzY0r5fQjjnyTzJGN/hQ5no
mNm4++VGecGLWTh7P5ehLO367OAMUK8eNs94/mzSXH3ZfLj+8Xg1lMTXp/wYop2i
IsOlMPUqclEy+2gFc859zXOYLhb+CtGOyS0H20weaH9pWmwdWSDhnTzt+PamFwlY
jxfvWmS3F8t7ekJHghcBZtFRrmQj+DNigDVGntrHk35oSbg+NuCcjSFM3fxQMIhF
strwjgfufIMmXxnRyASXjf7VLn8b3k4ymG6k/Bj4AtGf47hHm6u7+A3LdqaAevrP
qJchF2WbfHIar/ewoMSeEHlCkqtPFn+oaP5JiaasLbuMg6kQmphBG21tzUHPjzZ+
4SuOjJlbzWp2D6lmEh9cyWmq1kAuBZWNDfZLLi/Mj4jW63DUyfrKRmxSTS4VSpky
Ij1VHk/q8hjd9itBND+P9x8xc9M8h7ly8p+bn253llOhi2Z8HxDfWi17ZHjOpEp5
04XkQeWsY1e4d+6KN36gParcOgjbwFADgt86gJfa3qqbglYQxmd9AGLsli5zT4av
hZjo/y2k+ooMZVDXhTapEOxUtgHQOIdLb05j0VQy0+7ouWazYL6z4LVRbsjonY2n
Wrc2RIpNnbXUEacyhV3WzchgDwh9fyfFacnZNdvyEss0fEOAhyTeCtEfTa40MYAP
bQdCUqL8Vd73V+ZJeTo5AlOQhpSVTQ6927VEYkiKRHhXNp742DaFDlOJfc2k4hJc
ywu3fxc9lMe6HKH/VANsWgfmUf4AV+BW5qFbRJLNqt6J0l97VyFd3sz3Zo6ZOwJe
XOM5O4/K+VOa/vxxrRrWiEsQCqOr1yAF/MgKEE1JwbEHtWkl2lHuQ+W2EZCrGLrh
NDD/LX6gSsrh6JX9V7MR+1Lz01nZhV0S+Eq/Msgjr1Xvhgkv4F7l2PzpXQTJjsWs
tFr4yQ1X0QqUCzPOxKeCndY4uXw+ierACbALvFKdOuvuuu8RiM4+u6jad+Xu4/7q
DQQYkVdBzoegyIvR7sy2mONZemXzFgt4iGZcFPLALokzX32lQ4L4daQSXRw41wLG
6rqdnD8Y2Nw/rcKhCHRDvqLuol94qIq2odptEDPUvx/oV3Q3KiwdZnRhQsJhtq5V
94r9DBbcqP8jobR6ncTAbS/47TitImEW0TWE8vHjda9fluaoPXjTPDnNbEiTg9Y9
nie5t+jTjZEvtGllW5jiHbiRis/VriCQTguva2wnKEk9Or0fm1pSXfeQr5S2ZxxI
NOtoyyLXByMxMT6YyP1SNsIy1mqRNYDfVUcnfcADnBicB27+61wVQ8xQKoEVO+6O
zsTmY32H3OrF9Sqn6prPVrO/9VGuvQvBKpt5Zkgr6jb3Z4oFTJYkMbXtsLwRkGzs
z9IxBHe4jhUnu1CdzR4+2McKcSww7H8AlFJcmfuH4AGcO+tKKVjZiRD5XrFMUHm7
5boR/IeMqg11o1M2iF5aFPiVbjOuXsEAbrYEqczSCloeJJhlOmDOvcyndS3fzKis
PVKYAlsLWA7M0EyvioQ5pydFMqu8UWbk8erST/+vlOHcXEkDI2URNgMohylip57G
4CQsqfIUgAbZ8Wfxya1cRGTmAcIn2IZNpOvs7v/OZ9GUZ9CW3UPJlhLQspkqFMUB
mbM0ZQUNXluVA5KSTRi8FZiMjOYQ9a2NTmOYcGh/nJEPw0TT6we0PUNgQo8p1IfQ
y53BvbBSG2Xs4Kl6QC8iwNlHHhEEwqn1W5aTWhNJu5QaxYQosL6kvvJy5ztwEIB4
nR+x4rt0RDwXeDE2Fg0SvHUmVlBgfRiRHR4roSKMglZVymDE2bShsrKsAW/LNHrh
eXT2W4AA/cJ8Eb22CahvEfflMDgyaBAM4E1KVcdUmWvLHiKlTNsuWpVyKMRp5qq0
9PLO2G04rr8W4d4fxeJ+xhBf33NLrRD8CPxxXM/zJITYIr7ecfAQntJffbjYqlJJ
PZSH4Dc7lySvcy069yMICcQvynCURUvjlV38RPsan1DoAMT67DlINeLV175axVmd
LRd966pv69s4OFZI0NQlHa4i2NLj3dCK0J5wltoEI12/dyZ5XGRmePWGbuXeJUAl
PkJrdrcpNbqj0eVgbwGYCg5ZD6AWrlGTe1NzsRQTR41E9C0YPycBe3TjxjoBIa/q
eq/YvKK75qgsmoVgDOB5vRkt9ZnNBCkobFGY89PwJyhzTjLu6dZTtk4Hkazo9WMI
OquvHVvBI+YdMRvjxrkTuRlN8WNEvYw7O9SLCb2Lx6CebRFkQZOalw5WhyCQkcxz
bPnhtmjE3Y0OiyOSW/k3RAE7SoYlYtG1G8ndTVRgZMrOS9Hpkqj6ArphqRYlPLCw
Jnwfl7SP+WPJBxNXmK1mx0S30v4dxhEO0/CleJGANLmXtY2naSecLGljb0fIYPN6
zJZb3SgtDAlrdyV8FasXX+u8co+O9O0dnbxsvBA17bYZmEt/2l9ZCEaLfZ9zIyoA
fZckinpR6IocjjFGASI/bk/HubMtAxC0ZNMS7cM2j9OrMlSS8e4BTQw5roCLxY2z
0tu10jowTrZXcC+B8eMRtyWITyPOS40gvf86P+8es2L32PM0njVsXrC4FISiVcCA
1+SOPXvwAOz98QghIgs6A8eBAzz726M8LZs7+bOPUFPU4QyJ9c6jXYW9P0jjEHyA
m+eWSYOWweELoW9XsV58tKgAfxe39xa1UYD18bxTLUVw+CI2/7BbkrDCbdHvw17/
MTfdZHiBzqO5lAD35AWyOwhEnHxY0ylU8ihsM7DWj5ywAhVpsnXXP7JcImAZHcM9
bSmc3H6YirAlhpSCmnt3QuP688S3qjwYZGHcpfwc8qvc/E1UOUekXmVLhVhq+2aa
8o2kFinfTwSIiDEcWzprin06UYMgcuj2L3CyGIhDl2Le721zCkRd+aVAnUKVNEOa
Cb5IB3iK4K0ZmRbvpnJlXcKar1l3N4n1h+sNvyc6d0BqiJ8ZnHCYD2gO3cJKam+u
A892bf4RuBbgPNpqeDkaWuyvKOQ5mQSTxOkzzZvOgwQf8+mnfqXC1yRvJS3HLS18
krejRx/zQmitICNoX4wasKwF0x1+tI8TqaN1S0TF0S0aSy6wyViYVIaipWKqGc8R
97tmp8cg+FraMAI5zniMOhzs7rfu3Xc52JVvZVrgr3pvsIYaaD22h6ltomd/NIFL
Ru2wZoHoQXhD3lKsIzfm+0iFmC44gYab8OxE6SWJRJAkA8Y+LNmhXMsvn7tcajCx
yCBua+c3o+Dp4idrGhh5iJz+cw8BOfoUgKH4SNwGcWtwwiM3njCO1wh5aJc8f8Bf
KPOuXNG/MHGb6RAC766XxpyWrv6GCx/U54yttcqwIRIc40D+wpSVVDi/bGvWp0QW
h90b8juTaY4nmWKOavA5yOQ//mT05rlyqegSWN1x50UxOby2fK12p1t8pTbFHHh8
8cdyDsgKe+OLchDE3ZkuPAX5/bgu/MR2/sSGRlJrLO+pK6iUcPPSIP84nwtmDAq6
Wh3vhU8u3VeCVTmKyRECclp0OekTZXZXNfjCBZADaDIV/uBmyEdcZ8rbQJ88u620
ikcXk2PwRxbHLM2j04QPPU979W5wk1uzPk0I6uRNP/qzezkhoO51m1rDYN3g+v/H
OPkaZxrpvIPHHVK17J1KMwBFN2cH+Q1p8PWZQgDS79gk1uZWDhBELYxeWa92gOkp
Va0Ksa4jwamAkaiArY7EyZh+eUiPym7XOh3MdqqUOe1zEbn9f8sOuYOIgz0Gobpy
V52GsCFrpE/uEGLM/RI1NOJRW1/fvoWFMkBy5wIs+Szq3f9ncAZx0sQCfbB63P2C
1RT52xltPs8RMOQ7AHVum4EJcuwx9k/D4LclDM/rXTnV5sqTo13jSAfm78FwlQBL
8AdCZunDtiFm3R2f4HQiglkZkDpvdKr545mhCNvjlcojaeQRiqm5ub2WnRZlOSCP
TRBz6PCoUsqvZYwdAeNZZLTi86XXPZnrKCDyY4wKB+Zt9zeIpF1zFGKGJ9kzuVSo
rLCgIEZ8MWR/lmUxqNI9Su/GTDniv5KWVlFXIUUb7zmXPOWCK3z3ikxotdi6sdK/
HQUc9A+IPMVyhiLJR2yz8DteO3Iwz8eVTkNLhIAiI2lAtNahBwaJjVFFlsVxJqdC
Vbw/tC0/9s8S+J064H5NXFz8YvZq8d5qkzSVbIy+7vle4NEztJuSoCoaLaWokPfG
qXoyfgUPjExadX9O4/9yW5exe9SAgD/EkCqf8Dil1NU/a0awVyFL6FVxp0noIkpy
mcE/fXw7g0ma+v+3z+8G4zuaxNxsjyixBpRjzx/eS5RexdxhHU7nC45RUgT7eqaA
8C9bNfH+yjrWfvYkQj3S8+nBjmCUC4klmMObz2RgQYZpmd5UnLeyrXhqaaAwvXFp
yISbtS75W5wCw+HwmNVsLjXaH2EcV39XGt2k22wG9kifm5e/KVKnVORJ2fe3g3Lh
CDvElIPIEqNzrT6X77GLWyzFpgqTW0CdjIrp3KitbGd+XgTI5ihitNWFy0xe8G4Y
EZZmcqGRnES4uDDzw7SaDT0B2lBIecXmbZ5d9vvzCBnpJ6eUBPYldWymcWdT8U1L
ajaSO5yuSNHgTvGC3K8Dj9mhL6RZCbjotLnkM0OR8gb8Va5VL+OvbExY8VyaSxPT
BSAMnnUJLV/xt4TiL7VX+WrMcMis7Vwyr94En2YLKGOsPxHsZrSvjCVICRRKVD5z
l1xOWctWBUYvbWk6JgIUN6Kkt55QihGlM5Hcayx1UF2nuXYHxxAR9jRh4x7Ix7Vg
2NtTb6MjVsBhUS7Wjp/DlkTot1favlWrRaKhAEkBKrxdSpIpeP0XdqGdqcPhn5oI
xHQLSV4S552byTJxylH47/qxBmEHSbsy9sn7j8r0X71xA/CWVGZMHMyUBJOncGZp
PvEoYJFE+lITS7KD+CoPrdbZQAXrW9gk1ymKAMY4O8YfX8Uz+/VLk4kdTfzXLx74
l9nenW0xKQ5d9dPSWxJITrvZrgu/iM4yQEA5UvsfbltmlOU47MVnuty0UFDSg67B
zQqv0qTZhaKxrozkJ6kjgqbvCsreyBPliApMazNHlHuHuEntuDEjkr6GCWyr4nC8
wPKKkXDsKaSwOGYhhJCYeBd00Fk9hSy443mHdV3VnlxDFcF2m54WdLr3DrYMsJSF
ZIwyd5iMVdudvX3EUMo9HAU9VnsAu1rpyZwUud3rnaN6stUrGftvfv77kP3zU2pf
mBYJz14daSFVcEN/9OYpm1TaqFYucTu6UcamyHiqD0QkKtPxVQJpeduji0cFjOa+
0wtwKmBwuzNjAnP/85+4aYygOCUO7rXwLVTs+IJi1n7D4uxpVp+3dfnP5p3ngvJZ
yTiLm6D9hUCKIab6FGztbakzadRQg6MTg08Aewnalk/vVKj95Mg76G0LvYEBGF4Y
wOsXB7OXJXDnCqYCwd9NEJqGpxtB0eqON8qzDI/bphyqVhOFa4Oe5eOQZyZHJDc8
bn/2t73UdovVY2OroEaaqDyAHIGmSc2kXCdbDAki1XFlJ733e8ijWnANZ03R8kcd
y53SEUPd7fpDZAqzGA1Lm5kdU74/zPlZtBnw+nUU/Fp3L0DjRWzE0nkBCoG+yMHz
FiVeKPjDJpEwZYXCgNZOqOx25PKYY8s63Pl19CJgiy4o7FiX/z4i1UlBckhn6SPt
ajX7S2nVlGLdCV1zNLtr4Pnpvae7gGX70b508iq5Wb+Pndd8smICgZM1KRLP+2y4
qY2FHaAfR3MNtKQYSZr2zgOiyjwDIYKrqvMn39IoQKkMg6FJoMqzpVcObujrIO4E
uVC5XbkWwxGIJSctdbs3XKJJVVaWOSgNujpFA5IQAm47EBljDp/k0soOmMdfZ6Ka
iae9WtpQJ5/9qp+qL9vNQPPziwxzyyi53wj7PUj5mY6YosF2Y+PtKriJSSK7Z7Jt
NWBHSlXL9dD6C8Z+6+bqKgPHYs2VuHeYFiBBu+WHJbHnd/JvUq3Om2E8MAjfFfSv
QHjeV/9t3+2rzW7KicNGnciGx3Y6y/4RUFCxbJmNwa2LcLVwsk0M9dk7Kr2J6auF
x+vZH8eyYNv92vUhawBtj3laYU+XN5T1UAIusFZqPdibBvhqNeSp1TlgY2meqD/S
KOom+0RFPc5CxnVe6bIew6FQ1t4lUfYOyspl4NMOCByENfu4u5FSUsKzVyTFL+8e
1M90qlRksesdMcgOXo2sBYUDIAWAMlLdJYs8E+1z9RwBN3NKzvqx241N+JDpGVgQ
TmxVyGK953MaRYa85wh75kKlc0yd6ZlD9paZUx4F+QDeikTqE/u2Pzj7IExUe0rT
6V3CjfW2LWmiYO10taVvPgmdCqhORgPoMdXShlO3pKZNE4q9nQgi+xseGS84AlCr
/xjuHbj4e3YBL0H6o5HSgafLjxjEKLelzW5udKhLSy0ghl6OxxVaWGKnO6AVWeCV
RUaRPGRU2kiPMgI70OvPkP7JHVWEOdc2YFm+6yqv5fU7HMxvaK5kN9uUyarsXnMN
fPkLFP/JD+5XsdBhBipKy8gO5h0xBLUGVSMRP+uJHXZGF3GsJ3kMFXKLVnxFqXuj
Q+D/yhfBZRP/4hBNCE0bXeXj1CpE4+Qu4v0NL0tqoG57jlO81us51Nu2SfI10KJH
4cd/gWTGAuvMEibbmky9PE0pwt6qXZFEmJ7NAFRYgRkPBwLc2txcjxKHT7qYG5yp
YbPGfCZDT0uFA+27MycokFzZzMCuc2usv8AZuKZtClYR2/Ik8ki3i5NUOJi+3Lmg
oY8NFOeX/MOuA0LYO2P72aPct9RElH1Q661LFdVpvHGhz7hF/YOMQYzF2Pr8vFN/
8Up/9hWSE/jThNoWWlyEnWFPcwzFplXoJ1q1lMxUXnoru3jKQdDMbIMpsu7Q6sOz
A6e91Reu8tpI1HVXs6rJMv5GDrXKHlohTZDFBCoF5k8rBlL/Lbn9/CzV0bfNYENV
7IpkkgyAKTR1C32Rzp+dwyfDyWDTGMKxJn8RedmfYV1vXoXl/6co3EzrFGQbwteW
Ym/mLAbiyNZMg/l7z/W4+ex2J+cGju4nViD9HAmK8IdevazUiKPYdllg/hVXrGjT
nTVFWe950ULOsdh8b1G9e9/rbCG8CN0eFCrvPD0s/VR+NPJ69mBllbJNyurwEjrQ
Qg/LMcvwb0g+4n7gHu9qsm58xRibbMD/OpdxhbZIX0EX2Wt+lCMOCDkgAYqXSiwg
Hz1MKNSpH0IZfL0C9bUV8A0FLdkXNYIyx9Ca8FmhQj1qQlCfqwMyvUoHHS6NuWNO
6JCwnuu0DnfOZpFU7L5Bjg0J5NKbZXGobN2IWcck2CHNWqlRz6BLi45TvkkMAJOK
VOgGluBKqcxm7kOHlAE9gD/xkElHcAchC61BIwrU1Ftu/AiprXdj8nhkbruCKKzl
brZ20CeYr9FOEHy1Y31fRVRveGTUF9mIcUhpuzP2K3UpFhCX/V1Gpp11nXImRjB7
iKBfSnsGar8FZLSIMX1tBHirNQmMHCE1MqitXaly3PVTAQ2eMQ9W63++o0C4lCa/
8yksJP/JsnnVAjzM8xp3rrwGogcTRysyYXZjRLU9M6Pkbk1zq/xK5ApRQDHTpGea
Z0fWHviwnGfhuw1TC3JbQiR0j8wbyj491Vb/veAUbsdGod1xhgOMOtROt3PAspRZ
iMIcRT+xZuV3qejMtyNJOEzUYAplPewHCyNe2Qfy7nAB/8e54Rt1ENndTAl+RGVR
8pEP5UZOtrTgCFqnDRdogn1qNR5s8wCTJI7pzKCNKC1EVuRaL/0EGCYHS+DsvTXS
MyUeJLdbJbSeDpzrOqgPpiiP4E658TG+IZny7XCWdHp3DcljQAZDTxchwUftDjiU
FT04UII8Mosf+BB2r+oslvv5DvLgtwhiK1MvccQD0n+A86wdyhRfuMZBZqjxyvTU
GziBaOTYTqdDbP4x9PwbxEwkNKsvMsYPULeCeb/LMNugs/1qsJeB00lOgebjpy6p
LqyDpKZIM//vnoSrxoz0QEuSciDeLk8fBME4DhoEslk6tKJSWwAltvd1QhYlYBbY
rxGEAzNVwHGpooMNss8U+ZaWgQxIUVUhdFh+nMs+XofoTIre0xo7olUS/UP9FtYg
+riBIUNtAsb6t9cV2QCXUewRNB/oP2xqdqwAT0iS4ca0/hTos4jAUPmR9sCMahsm
xvWcG9y2etbiWORwgfCuOn9M0MnE6HWhr5wNbemFEqsOwmqqpuCuZwOgjFv6BuNv
oGyC0S2OLwBBR+K9U4lI5ghdtdRchOrvO/tO0lypql86eRxh1lMOcPzAxtq8n1Jb
U0VNUCzcwJNMuY2DaknK+y0E8gimMftwwzUGE2/H205bR5h1DbUSp405OXUXFAIN
XDH+JhJlg2srZzTwZ84Xw3bCv7t6O2ZnLB2F34Q/YNWvhWYxdnMbG+FSlzGkv61c
+HGHbefdyEPBHiRoU1LPsdCIcFyxDVRL01KH/0FINR1j2qY/SfqPiQozx0vjuTOI
Z13hxTCyRl/gk9WPV3+bV2VlEEW8p++QnzD7g5M7SYIqL+j0qHQ2+Mi35wPy5V1J
mHBiLdOlZNsP5Fz3E9fmLuA66rqaMFkkkd84Z+KSnXC0Vlen/nVSboQsqXp8k+NO
moungcR3KsUePbZaBOCred6spUoA3YUudnIS6QdOSBLWUXyh6U0D9sq444XYZOBu
R4oPcFCgsrY0Yae7dBYOFHge7cRH0JE0N7RLRH7poju7905Hg+0Zkt7OfBeZs9V4
Y9hEhTaqucjzl6gxc3KqLJg/xwmoRumLWisNU10uT7DpJyIzAUw1EKvGUxbFtM3K
uRuj0I1M0T5AIsuCoCFnE4rTcXDFFIweyiMG02VjGh5wNg825EZW+RRVP/4RehOt
r+NhbwfEXpXktZXNjwX6Ybyp/QF1Rr9RLZNSwQaa7d5v1f7vs9CLUActHuV69vw3
CT+tJDxOUb0sGGNyCvlJNjWf8BkVLxBzk2ZNld0QGRJ2yFSAMm/BO86gK8TgfWW/
azOKNBfdq7ol2Ay9tFOsDyD0PgS/cTKy4qQYYkuQbKSSFNgA1J6oBCT1EOx39WjA
VTmpyoHObWMjthns7fYGasFM8wJyPrVlYByYCuEEwke9qJ9/s0HQw2ah9ZCdSx3C
5qTVbgTCVwf87JuG8SiVEfSVYhudaZZXMbfaoFmfVmTT7VrzGPwSeo/yYfqfjiF8
pXyc7D/WkSjlNaBSXtOXBWzGxU/R8dvyi8Jmu6F9XWUWlcM9IOwV0jbUzqrrsk1x
EdQLxP7vjdgLWfILjeYAQbRr+ksGdcUQacJ+HbPZwj4BtFTDdr/7kLMbfn/hOYF9
aiFszVHZVKKnBhTARwpEvnyibMIlYKYs2eNmWwN9A1CV2vBZhgRsE4mzfZFYsTGc
8a/J6SdXnTm2LcyVVMQJbhR0/ravVtu1rroTpCvmenB7ZzY5VMrM8D70FyLmLU6R
Z4nAcdb4fgyjcBRD0op+lPcT+nV9rCkiqHBtZLY+f2V5iEht66IgQ4A7hYIFbWzB
vXM3Bh3v38+KShgUzGBSIwU8JmBIKUOOBnOSdjCvVdLfJ5TjSdr6WekQigFW88Px
SV7OKVpn3QRn2zYsx2+T3384BRPzJpKOSaYWRsDDJ14V4Qw4yO3Kp2vNhBZ2rB5j
BrtDWgqJZNdPapVc31LNjHmcZJamFA0/+zJt38MM+6ejyBAxsiGQXpb98GoG1jQh
AhAVGvF0ySuqI+q6nWsnIZX0IllCRTUkGJab96nY7uB4krtAhvyckbqezsbMGeEh
MuA6ReQv4jzYGDBITKHmDUyr7zj/etvd9SthK0K83iHAd5co6LSsIeaBmwtCL5VX
J915AzuJLrEphn0zzsmrRy8YlVtP/wTXu7YcVdLX4q+3xE+w6TPvhXyo+WbsMD1i
ROPLI+F5hSWSu2sQSTYF2BEeKzwqwKcHLTqLjJv6TpzKU7NYEIFLclRoFKiyWWWA
mEa9GUjG8NUTQyEKmowsCbaWRI5Jyw8Zc2pTkxK1J1p9ZxVNMK4tFRE21PzM+59j
uQnquxOhheXmgMaaB4wpwjTZAOfLoTcsvkgQoJbPjcz4meTFJ06+EbKkza5yVxUS
SrgzLNeRMisViAXhjNDrJEMznqsmvAM16fFzrB16d5uzeG1ZETsHFw+lmMBSjPku
nB79YBLPTf3eCV/jNFYR6H+vi+1gRIOANucwB/1zk+91/6KXyMQSoF/+ChUsNH5f
kNzWwy7XAa+9SODDZZKgO4MKt7n/KSbvo7ZbtpeNyZX5VfEK4IQHOnOM8ZwSdxRh
YlSN0kdRbG8mVPQi0Z6JnP6f73HC3aeEIq631Gh1DpxlU4Btbh0hgBcSrtNGWBbP
aMTW99DlkE0Vze0beaWCkMEQeXkjju1n75ueJcStxiabhxLIkotE1On3cEgfpo5U
IlDJSGYVKeFS7Y0pWWNRITkQN5v2OEYCBy5jn4ySuzotOIW2QYYNIbytT0g1An2e
9Ubj1Nk4V0hICyR7KdfZNvh6GzKWH5KOrDYcM4yOutGF00+MowZ5DPVrIaSRc03b
HC5y6JFnGkBxBHKLKNFYCGqKyKxtdhXZGQykuVrD8WuT/Sntwa2Msxhdp5U5CCBV
nSNDAiWxsbhITrziJZDDHgyT68sSdx8WU7IgzrBQaDPtLJrBbqg//9XtiXiNWXnc
pMDTzpn4YIeAhNjnT7Ul8VTYLxSfKcQEkLdgiZDg7ZLWYOGNybcM+VT85rZ/RqgW
yao+uaRQvb3rtsrAUXUlxf78TzpTlXhLHvNl45+dea5fo9aw9mqB4BTFyaWls3nk
WBVVwAg0w4k0nHkzJ7gqB/gFArqOlOFnRyXEl8VCtQ0VdXMq1MsQACDAblvQumIh
Ploql3YVgfNReQ32pJv/sXsTNTkBrHcgUlUYjy99YhOsKgIgLb5X3uiKbk32fg9X
FunKlsgS2yczBvsGWuCF2c8VP77KI/hzoPYbGmn2ocgxXsdDpVIsDR4wZxuHZFMA
qnXQKRN2zObU0PPPrUOF5sfo3aQXX8eHQUtVb2wQNKVXgkOm0jR6OkCK6rXo3wCY
3dahf5RYJQPV/M1eI29ly10tQJ9pta47vl2i8ybGQ7gz3ejtpbYDmqpYIGSmKbU+
ANpvjwTNfmO8bQfDxCvDxPx3mc2Qq0TSMVulaUdYBVQljN1pTHLlr2uAqcFQlN94
DvtCkx5o5A8fP+8k+DVRQ4qY6YvvN3I6SFc72NimdZ2EQGECKExWaNnkBaXDR2Qe
R3SsnYp0CVPrZ/gpNu7Xtlz+KNM5a+O1Urmzf65eg52IF1LtRSR8CWSKc+3ucoSV
IbhU7TQEjSGvxOsapV37cQtkYiMqQB21IAsYW5j9hmHiNK/6yuUtyQhAUWQFxkvb
oL4jKhCJ3hQFLxn4oF/zKk95ECr6oz1Qb6FNHBa08VofkLbTLWnJO2bwj8WA17zF
kZzzuNVf+gR6aR+JfcNteVhuXe8qzGm2ZQvUYlUEXaKVz+/ZURKZfDYMwYgJQB8j
vIN0rhMOLwkyD8xSIvp+HZ6Bwz+WZ0kvqzpOBp6Tn341W8/KKUTZgPbIJ9R2fYa4
sWgDwTuxWbdc6sZzqVP4XVLkoydeE+24CpkaSBxzB3zM2EY8SYdFIrMk67HVcjqH
HlJwH09FfPCKR43iv5HtV7N8oZJCcD4CGZgwo4GmVxWgUHwgzb91xEkXEPLA7byV
x4K6Vmc/66lnUlG3i09NXHZQdML9TwpTI3dzQBfDAWPaC9xsPdH4cLuqf3GVvFYF
Bf5GXarNmcx3ASVcoRJ3/G/AREPa40r33cxpr5IHxxTO4Coc/Q733UulvmDr4o4p
PfIMPhX1iiWEEC2WQr39XJS1ATFT6Tyrg62wthhy0yq+Or6yoSnApUWu10e9PvbX
KjlKvfUcFvccu4mS1WhARwcA+qe0DbpB0S0TZgCQKc45n8CdSsnuBGohPR5RJZ68
9KMMP23XmS3jQ1qQQtDHp5wGp9X4cC7L5ycxOY41Ev5ZSTG0azfum1np7p66vmgj
SYeN9ICHcUr9PySHUfkY2NtaemksTMLOenWPAZsZrSsmDX5QKTe5VdMlWGUdQaUP
TV5bSFJSpAsgjt7XBJerU4GvLnemOEyZrnYfB9cCKX6D9xob7XE8Mii0aREHDhXE
nEEzMERR/epqxNss/EqbfmdLDmfkEWTiC/jTiumlkHDQ7jevzvHYXeRVC3GZayfe
etz+oIxkX9n7Aih1rjCHFeQ52ZvMPov4/e+G+omlGnmWFUuhhyEJ8gorpbVa7mrK
YPJQzgWF3HzsBtyB6GnRdtcMBzhovMQUQmR0xtQhFHFE48zfc98jXRZoLca//orZ
OOa3kXFRcguBZ/SKikZz3oP0WglC5Wr4Sj1ZeAP88J7kgfhyHR7QuY6sYlZXcvVN
KKnKXgB8ZME5FwNDiSDvUhK7oaSzI2/oKmSOZoZcbtzB+OR+Ip/k1Br1y5hta5+7
yqwd+NH/wa6H3rNWT7g9fDEffBm7cw9k1RSd6RtYfdqRUtd2KI9RulNKKdWZ/kGN
U5VUAo3rGUqSX2brv1zWoehfsCzu7qOn1kS9GbnuNjw4R2zJ8he2d31rpZLmm+J8
K2g3TgAqsNx56HirICLQcsJPXne9QhuUH5rl2+/x5tFpkYz1mJrfoJsO5EVhVHcN
Oq07/3m01s9wb+zsOXQirY1I9aCgcwSUNM2NInkRd5Ju8dkIq81vXSVAL30BpII1
3NOgnRv803H+TitcIvVwc3epMtWMtWDDvqxUQMjPVEXnDIfDWZsrORky7iX5kI0a
jQTxSnXton0jhxDYWzqZPPJ6V1U7XPGyGqjMpHNgUnW8L+ZrdD6Hhc/sCWGnD4Nj
KizhlQg/vnJswp7mXGmaFELu0S8neVi1CO4On/jEQdDYaYvTthkVIxd8aN9/kXhA
tYnCYTu/AaMFx18pC5WaX5WBZn5IUJgX8ZM2tWH5ET7a4BnEckeYWAlJPj5toLYe
0w354dRawfABLA1bt9T8J7np5mlgkNd1m3KGykKL6s0NCR7EWxFJFW+T2YVefSYd
4iXANg895TtcuN+od7yZghxmbY9g8/XQxUTUr47QTIBNdJHMyZXZd/1y9MQAW450
THsAvviM+YhbShRz7yhPUZ6TCVDjXmH0oa/+bkW3J0LpAaBaK3ZI2sYXSwRtOgwN
o/0rQo8lr3E4JRSlsYiNKHJ0k4BRTGOpRhhNNqHese+Rz6YZVL9ZIhnQHZngnOcn
TNQ+n1bMMoatWCuICRu7pGJfz4FvVisuoT75BRtOOL99unKZRbjvTr0HVu/PBAhj
vXZmD1cWMM1kLCnWlWtxF6quyIMkoNI1EtJyxB8/BQ/q5WmXjEXT+iMBOyh553dL
tawpYsnMKVZ3iZB94KsztLJeE0oSWZqlsVGyefJUCYQ6/UdzSSg4SiqPkpmu0GDR
JG0k1ZwYoH0Pgx9o9HOWbtWJhr+fMQ/UW570FsRzEoegCpf2cxrxqMjJUGWY7cOt
MyZqPogpRmWJwsUVXqZR+piuKRHyXnuG8tksXIQ2OKOttRNCH2GuOYvRuBwzCcAT
9VtRMPt/31cKeem8lS56IzsMTJ7Ih0RyP12uiw3NoSSEYsO4zF3SOgCVsxqN/B1J
q8T3HYevB/lJI2H9P/F+DqaaDwhQiXOnXqC/JzPs/gmoD2Fc9Xerpchk5bO1EeAW
mcUUIWtbnTSYgv81KUfvM9Z/ntsSXPrrD65jg5w3WgYiu681JHXazIVZOHmk5RRB
zlWpjwV44LL30DRFIUFR91AvIqnFTfVCRHSb3200fOhcntg0bqnnQz8QI2CysvxS
919XlZhV6DlguVSKiYaNt1OWx8KILw7NtZiCAdcxyreOy2L1pnHsk4e5MYr2w7f6
P3TMk9z49Zf5PHDs5WsXBesC8L9jq2AJSgInjcyZN1cH73PGT8MZPkcqCQ2Lddwq
46gkDQtirFRKg67nVDqh9zkbNTfbzjhepX/ibuZyIK1yBZP+5NmOTKdF51GazBCm
masGcQAG3mz2HRqzgyORCaJCagxdX8iwVsV3JQ60ErRb/cQycQDp0DAc5ng6ap6v
7N64SobDvUAJb/QGmenBZVYQ6DHG11dqYi6AmmYka0bm8E5zDzpRS55s8VtUJ/U/
9jKAqHl6+uij3iA+KTkB8/SZHdzI5Vx/fHNWFK3Tgj2Spxe3u1W1OO0Crym7zBWh
E/4KRFrzBKQ8kN04WrbhuhArU/SWjF2zNwENdA+uX1qUiyZua+mL+u93eGtz19cN
5nzxbZTE6WHJrHVQR/JAm57mJ3SEh/BAAd8/I7UIlCH8HUNIYi95xCdmrhLIwPAq
BYIE0eCxDecbZSkRGoVSyT5PfwlvTU3Kars0fSBxoNF4GreHez99aAidLdl7VVMg
jXBJakm9Z8ElsGF6oA4Xgxn8KFQgXYI4jra3SFJV5+jDVTWFIBmjHCUlRk8lMLB7
0f1/H1cY+k83NTcPsiBu3iKDtwrRBKe/ab8611wmDCTJgT6972DdXYqeP8cmH0VT
dFxn0KRouxq66Ii7cvNW2ew0PBRiWtQ74ZFv2G1tNETtFBJUod0EMmFC9tjtb6Wi
z21wBTprwXhlAwcUZADaUnxFi8goGigiIm0PircPGZ3jrYuMh9Ge3ijw6i1a28MG
Qlfl3Nkg8v6RiSkCeedTkGHU2/2qMd8DPr69UAs8uAOUIrKJGcKEFqHqGd8OsZ7d
1+I3vLRxa9w7QOuQlP9Kc57s3x+fPBF91KO0HEOOyXIRGpEFnpMg9MFj7aAbsVy7
0u2WIbzQKnB/5/G56ACqrNEqQrR8ZXm2M7zLjJ+yZLHIylcmVk9rVFTA7TAMWxpI
5QciNikD56zZSC61MXOQsXMUz9epFDVwxBtyuAn2rftQv10Bwzgqbu6oZTvTqGWT
Irm8IxKNbEg08u3IzbCgUZTmeBm5xjrDLhFX3Jlzd0oV4xIX4aMxQ7PgzlGZ31Ku
VfjbHBXiDqt1gw0xpkkd82f2QLsLF4DtZWuqd/BE37gEg8FZxZBmIaECsxk5qI0T
rB0J0/UPVCH8cxExDlG6j8LguipupoRpZL7WBWxHrp4sjLvBhBfqOxy2AUHzAlZ+
bc9bQjKVREoHQS0WHrin8DGs1q5bbn3nCfc/1eYccoW2+3X70zhdcLyydrGpGgii
AmVvGC5Zz805QJV4RSRljX1gGJGmsiqK9/Wg9Lr5AqbKvc637BxELhK2BaRoVmPG
3FO7FM5kFeJftZlfFAFOiCCZCP6BHXTeZ1KAETitaw4hJfjlq3GrP+cw/UjhWx9U
xLUSUjhsw6HJJG9+rcw+sC1G9PpszrBJXUax7ZjtGSfyAnHTrn/oPTz4B/jU8PL9
nYmWN8gRqsf3AQmdxGtmy4AI0KrXsDXgCDkJgYXESGye3Y+VBibvhwBK+HlthVx6
spvUOoowfMe4SCLkaNAU3fSq8g+OFVyFFRRST5nXjmXzw2o8Z8DyC1p1lr20KpjZ
I6BFuU2940/1pTbmICzQ9TsanQCcZ0RVr1K3IXQfGwubnRJfQhFh8RKr2lrYuaIY
2bhQ35z1fOpCYNb8cnDaXDenl+C0ojJD15VyIoEkhodd+2Wn3Qg5khsIYO4dnOWb
Uawl2Wpt0//OC4zqKen4IQL+7bcqbEsQLfx+s4NKNUFW5QfTLV7bXfgX9TIPxLu/
/pelQxwNKItSCNs9oGvkywekCbI3jXTBStF4MoAwXqk64hI+NwgzANniKaTmhMiK
R+vZXEfJ+Ac5qFYIIed45/2IDJFPuEH+bhtj5FaHiM3Wy7VSE5FxDhKKz3vZNRXr
zC+U9O7sgb1Zum4gtxarf4vnTMMGdv5IEyJkfCJ0vCvJ7ZocR2gm1BFyQemapNYK
87sgBLNt8HpKVVPLs4ER09ABcn2/S6iaFUg/NLPOOWWnoW3odcBA0GLMoGv5nckx
m3m7wQeVWB9pCFtnnLlj20z3SjZdPHjQT5y1rhyRBc+oECsI070/baVu+NH2wdv6
9DzilskXygDR7xAEsPkk6ZyJspikVhujvW6hhiXoZfJVs9haYKPLlRLcrR+dumlX
QxE3kbAQLOpPbzxdJicD95BJfB4PONZEfIBdUyF2Kpy6f6qU+LkKuoqpMNQQRI7T
JI+CdMtUBbQp0XTEVSzvsJaJw1GnB/wzEBiwnmpBrsMijcO9t1uTuhDwko1pxAS6
mb1BOhYT2dyY1WMxvjh+qCN/mhLMv5Q5SZwGNQK45FiFe/veLHicIrbqyDzXC6jy
QB0TgBZRAfUpZ+4sKrVyTB+zpCJ5RkW09fPyqyFMXvIqkAU868cf8l+MyH8EhIEd
fiX5C7ejAbosh8Tt/OZCgmOYCsRisRe2EMCKfHWjAH3PW201a6ukUFmmVeOlUpzg
UAM2hmbSAC+ZTJ3n/mqkLPzJtHMQ274OstA5Jn6S62hJBrKPN1/c3kChCDxFMJ6e
mUfbBP/62fEO/McfpVuh7xp3Yr1IoseTCiR1AmMbxCXqCFE1bPQ5vFCv0CBcPUdS
DS98xkwhJyqVMrMv9eLmOZLa/SFzq9s+Rapsr6d5hOLCupi4BSbggVOxxdMDtwtY
lBr6tyCOtklJzYtguq7GVcYnUjehjw57nVDaCliqIenthBp1etPCUG50Oo4vPBl3
TvszQsyGJ6X43U7BsTaZsmDQOFM2BP5aNkbLsDjG9sNN9NETwalB5epaGAokGtiC
d8ZO/XRzuq9zPzeIBQOwOecU9Rm0HdZ1n/3bczaVWcrauVcSfYxXQJRPXyqorEte
chN+gkhCG9VWHGTBnQaRuXR8GBACh68mTlpJMFAM7G83QOta41/+qVV/7WDcZhMQ
lRprWe7apUAoAl2QJUyyPpyQu0Gh+MZ+5JmE3l7m5Z1eDbwz8PE2JGKzTU2o6oMV
xmPuet0bvTda1g4gEp44hdW4fK/jfpVn7+aZGZDidNFYkj+BnCEsIMxOyeQ9sYXo
k/NRKpRm06bATpPHjNV+HPcX4/zpaS8H1J5rvqLUTbEXKkkUwc3jt1RlyD9I96Oc
TZ4u8tbuPtdxg37rz9LB6X9B6XqvgZyzleqPACEVyFkpExsYTG997L3+qroPuf+3
ijHJwhoT0s8MHdjJEH0MEZLQIk2o4Dz6Be/zcr8pDbSV62RDCV8MXmMspwyzc5BY
Il3e3xVgJ+gNZ8AZVXg6+ADWl/HNa+TVgTTpAp+sQBTUErhPSukmjuSoBeYcAMzZ
JREQDT0MdRQMaHNsin4WyrC7U8rjkU9YnXd382B2w9IUtH78MIlzQ382WMtRc8UI
m/MuVPaSE+6z1MdBCPE81SFnvPgZ6MbPsOecB+rTkUD3Xp4HRnucMSq+8a9HIMZq
lM34wz3UqykSaxVt9EdorQ9g4LTUsWXTrk5L4Vq1b5rNsOViuwnfDMEYWDzDC2Z9
2nhdNItOsI07qsB15NAX9P8CZu1pskAjxlp9LH0dYjYPDQAAuraFnSNwWdYyJeSa
JnphR8s79MgX36r0cfxLtBcGwRv00tuC9OSLxaFlio2qKlCfQ4gc+RXG1EBwWaQL
BcsOMyUqcQg4czHSD41hxVUPsr181dVrdqk8NiaUy4FcysXrS3Q7SZi2m+WwhG9V
axZORLQbLtlqMJ7/HcIy5qK8440qCZSPusrDuU2XLZZOkQFPJ4W3xHiZYPdkJyHl
UTW09koN84dzH4gOkw5OhxrLE+oywsCV3YTjO+DsmzKPvsOboCtRKvOPaLNLUPP4
4viE/8gRitX8ru6e8iXG/QakQH4ClwL07SPLO286gsyYHUf7/Q423LLpicvLBmXD
9dobI8ibzZY6K6ypTCmU/S66qgoyFmXBAaucaOWxZ70mykrdE/GbGqBVP8ndVw0f
X66La1Dyv64N2g08sLZdWLrMHGLMvo5ORKocYzqH23qZ+EOj160qOAqTatlm2+2n
g0ENY0H03pzUVGnKP5QNAW0o8tVAdDnmxiS6u0H7JSMjSEoDqw58rKjhuQ4NCesv
UTfDabMo9Pz77Z1h9/zocdB6xYey6Y/KgfvJ7vKQC0d0GADNU1ZVfeKdLDQDtWOB
+oQ8zXfZRDnvEvAt3hiyRAaJtnNHiHbqzZ8E1T9MBf+Po5G8nFXiWzWk1/fRY4hR
OqNuznvSC4sQY7MAqD2U8wOr4n0/G0vvtk20KjAF1ZO72TpxUZuUz3kiokUuii/N
gSAZn465IpkrsEjpYrkxzO+UurnSVDPwcEfmvGZqkmRt9WKGF2u7BC0TJtRzkGQK
vlCRiJkoYIbPksBiJF6aXyr8/WUQRO2Kufgjt4mCLYbo6ktfQm50KDPfCvPfYgDR
ndS+fu1WBrmm/3NSVAcYUmioKLWHL8AMs+zkfbqiMJekZJWf2C9S+beUVBY+sgsT
tJT/QLAVCX0Nr3j+tbpx7pVVJp9QWdqF3kN7RrfIAXUUhtKnY9w7EVZTcPSmdRmB
2k9a4bWBRWVnr7Yd28bh/5vBiqMufUYiPk/YhpDFgPFD/xECQK9Av68vivIWHb5G
A1KxT8p/xLINS+31viEJDmPSv5XyBB+s0kBPX1tZCsgGJ1enZnM8eakvNVB3kb0a
czPaeyCbNrNWZxLPNbVOUdsfvFFDsZjX1//bh2JOsToO08qxncOmjex71AiRCsic
JjebteXrVxO4VJeqCoKdyj+GWXanzqOgEDrSp78Fo+UEVilOKQJKxbfiRREnEVjT
X4xM7+EmQnrnWbu+4BGKwNix9M+YeoCh4B8sa6wW64vNV+s4P4eymdINxm+8hoNC
/915drACR9PKehQg1qtf24ysOzINecCbzUB7Tq2SKH2pZbVyQb1+sI9j/jn2BqBX
fRvW9OGRZk9uSQVsy5hSd07edNfPAW+AI8XPjqPwjgYnI8KQM86yKbzZUTzVf9Es
fv0mnPPbvRmt99wj2/WrZZlONgr6WQgtp0n9i/2fi7+D+naK/h8UuQcbhNoaVZYj
g0veFjSj1gzTeT3swr4kPVUp7zH29GXKegzrUKUoE9O3XKeP2S0ztXFMKfk7kCAM
mwpwl+kLvBi1Nz26cmrwJJs5W75OzIciI0syc4JwV/NawY6+wh3NrZwQI3pwqsZw
+IhbDcjyjCbm1c1JZk52urlxhQnYmO4Nqu3Rl+EPY6MrmqpszWD4Zx8Jn+ULIZOV
eSRTWosX619oVIM7CFw7G2uuRw7zfI8hxo2FJavjnVL4+mgf+ala5OwNW14mTReS
qFm5mdw0dWM+RkcbSz/J0qgZhn3j5UCuiKLEpeKD2vuvhAwLXcStT7YjznSKlJ4G
gRtPTiN7cSM/se9V1Y5JBwJfGJc99jWdGoLATV5XNkmTloMz5+LJ93kcL8w1Cguo
X6oCGfVned+4PhpgxI9RQ4k4vDCez1ZfXp+eUYqmvoIDR7H4rqgMBkEm98ZQoQQh
JqghFrVL4KT8D72YGNCQw1e0ceqNfM5Reo5qiUNvopPHvIoBRCZZ11/7LA1MzB62
YqOsT/VWFMgkaB9rUaAlQbalYlylOu6Gnvg1PZD7UU31LXpjR5XAZ1/LISqxJ02b
HEq2QXfQ3emK0h8jqUkFDAU/dgBonvvBkiIQTqVj8z1vgcZ3knPeIUn4s5KFR3QY
oxTf3YHFlyhLuOzm/6TvrqJm2321sxVRURlgrgVzUkdYhxeWu+NIIDf0we9HkiCU
TiKu5Tb2Y1zHn9D/IxhzSKip93706h6V0Y1h1iVZxQBb5W1BRfk2iTlBP+eyKHy2
LpB0rLswGMU/xL0FOa34pptBqu1TPkJUKbP4CtmFncrbx6eUQw665xBoeX+3leUT
5AKL9Asfc5fjAb5whZWxWUo7a0GxPPEd0H3ZqqIqp1ZTl4HDjsYDvSzIqsJFAKYB
3C54BQyWVw/IrhBy1RJ9sQze/VRIRKarzKCV+ZIz5UY7auwy+cXvR5TAbCYHcDoi
obzW4gzvIJSdaVvK43Ha/3LEBtEY1uZjSyggOHEG2NO//A6ll0EE8bISkzkNjjbU
CYaUHqkuDC6QTzcQG8dacNqJrXQyXpx6WDbvCBjPtIcQnZ+ZhPYeSsxyJBUhuxXR
TIr9RoOausgMoE9V7iItJ9Fu3SB1PFzyI3pJXpw/KA+CJ2jYk1Alv/SL+xor9n8X
OyVcX1HZG81qjvhlH9Xx0CB1P0KhNJungaLD5OCAi7T1cYJrMl1n4z08JT4EUyCk
XrA0oZmETtflNSq4IvKIixRMQDlAXsAVTclGwVIWWeWER1FnBnnGCMl19YCtOfCV
wLY7EryRafIykYtuOYC1u6UUSLicNYMjhOB93PxvC60VW5jbHoykICN6JT3OdlKK
t8PR/VrxhbdeoYSqmQfyeYetrqQqlsO5nK54eocrajwQGvnzePja4g7fA0Gf9QHg
VnYGVYnEkOMP8yJyikp4KxfDuWgkfRBSGbBUuBHda5gWThwpm7KMBjyukdO61kmG
NFG+BQmFCFXASwgjCPyn4zIwXTeBkNZsoAheCFErgJVioOmvQpY2ynV/5hh4S+DH
dcB2hrez4+jhJ1TWw6G8RrwlKdlK2RdWO/t+IIDBDAzAVyVwIXr6uq66JVHv5qbY
m38LK1Ss58n0OYMHiufFDglHI8awcl4WbVBOGxaiQPYq8gmWUyztlP1moC8WmPNW
xDiHOL/LO7jPCpV8gSd1n9I1olSmPSKsMiNT3qPcppPfA+51KeDEN0gizlxSR+ia
U/d2UTgU9WUeXjgyGi4sSAs0ggcxloS5yu00YV1rfqg8zGOF6KFRc5v/KdIZRubk
MwdHiWT1gxhpWYlurAlAcpTuEkibt1/Df1bbJt0zJ0YTtMr45Y24vQWBmwhpG2uu
JVK3OQ2HgUC6VQV1ib9CYfbP1EzhWanc8GX3G6f0+8QJQL5b55wk9BgXnMgOVpN6
2y0efUm0QbosoKvu7QRlXJF8lh7XGheN4+R/8FdQERhYiQDoIyEYGhifL8P/+FLF
A2NbOcS+SeVafVXOmMO8ydYsr2BQ0GNKBvz/nHcs62LzZuy7z/WYMcu0FLyMfy8r
HmJjOlF7Md50aget2qsmwNYfQcqVGtnWPhEJPGCAwnuBp5J8dnm/rnAqq/qjogrL
sLQD3svZ+EqkQq5xb+NLc03DlHB1J47FuP3cWBeDi+VFUEDBpDstQ8X53Z5zG6CZ
tGYE6XKTzOfwT1C6AT0QqbBIFPknb1ormOI7CKw/befJCmSzSCys0SXzcSOHmxo0
gRyaEtUvI9dz/zQcJE1QfLXxK7iK81Xi3uzRbWKRKSj6vlf34fuoIbvb6h1+oA2u
Sq2FZUczwJbpumQR4NL3XA1Sc297wPeKNJWeh1mQ0h3IkVqrVziI3I6/eb2iQ8+a
9WQ7FBfIN1sTXaYRcW6VHPViM4XtXVrdB3Vb/tdOHLQ9ZtWOefoMYabcO1MpTGxa
AX1lBOiUAyrFLqt8Re6yqb4ANT6dpYzKl6KCRINi01PqaXDGZreh/Kt/NGqGlutZ
E8i2ccxP5Wenvy/82g0ylbmZq84Ya6HuJFUafZoLCqK+16OP1SKMs5nK9yqNYVtb
TX8yx4SqRxaKFtgInZxn1wo81R+RikrgMKl/eEvHCeWUMwploG4DhvRFRGSH5mPP
jmfpLMjnUVD6VddItGRn/VjqH42m6Col3Od7Ds6Ylg35Nxuq2hH0T/r48Nmp1Pdk
l62myjuEGqBqGjPt0Tj34OeQhLuCgwJ1gWJm8s2YlrFfoFrZGW7XihRhtwfyX0O6
BvYAvYV689+zyhijpgAtypBL2CNtOHwqzibPd4RLUe3ob9J2eg9ui7ySscPWZba7
p8/Z96QOmwFflc4S4o7CpFQMmSCegX3W+8vuf38VMNjaYFbYqECnL3JZsS8oHf8B
KX47oY+am9UL6HIZV5JLqR8Us5kTfmSNt7Bf+iBPU+bHjWuUt4fjHrEVxH4DbURx
HzgQgbs3q0d8e6Qw6vTl9DLAst4ZqofeAQT7sqffbjkpemgTxx9DA2LRznvugm2z
lWlXEzcjBMj2H4uCJmOR7h6D7F6h/kkDbZ9xVBzQfLTpj0d/xmVvwC0SS+meoDaa
di08YP3jftUv3f1TWK7xMjE7wVdjTOBlDQd8EiwS8VzIgKMhblYpy7EuKA8dfRqz
+lKGk2OPJ96yPmEOY5bufkyd78Die4Goe1IjFOUK+xu9rzKFkYhUrsNeWkGZGKcu
Z9ZmH5n6X0L9lN3JO9lYDHZ7K66dO3h179ffUVnM7MAR2I/VUgyQN2I2ghwjJdIm
OLkjfkmM84UpW/IRbxAN9vPC29bId5NJjl92DQxzaONAVdyXYO7s5TU9lZuoP8Es
PdgsV6Qe39UU6LJX6wN9ldslg/lM1RcGSp+fTZ3yTORMtRF91eXs1tKM6uZHdlRW
a40hWqUgrKXgUMjNdqpTUyG4WQmWA3nahuTmadXuR4l2XYkCDRHy9tkJ6QuusCkw
/x9NROYs62MnHvmwjH5rBHpyAPZ4th6VFuzVcrJ6eHXQ+DTSxpDmsfdplBjFxGXe
JGvvcnhf5nv8Y2eDogq4pLXTKb9BK/9wKZVCXwCdI9y7SxTX4zvENid29VmMZ2hF
aRC4sXJxRwliTwns02S7YmglBYDFQabaKiosEuXN+WEpwlPYEMKd0H5zAJkYTiHF
N6yXcwm820xlc6+iVp0f/SsX9nOPeP7Vf9h4Ga67l+2EWXmCYy9AmOrgR9djniSS
imMX1ZdaGXbplIMZRICudbrFEpmuCYDIS1zWFXtRKh4m9WEju8omDjivyd6nWdfA
mawyNlDEMiurcVpLBeYwm2wNxDe0dIPHrntNC9YC5ZQ0NBPsZfpvsCKYMNyO81I1
bR8We3nfr/L2F/vRx9rgeQYnHMuriRTPF7IPi8icyXETLpEFjXE7YR74vvNOqMo+
jgIMRwg8r/OHuLquLugqJKER1ycGqD6ZHN3yxK3UguVdqfQ7fDeZuZcaC/0FMeyt
YIwu81qlIpM6uH9b4Xo1FT8L9foEey3ywXy3nTTDXn/VKsgqfOORUdap0tbnHkay
tFUTmML8iS98J573hmAUm5Skszzm2/m1egaEOI3M5TuM5TSh2uuknpPBN5RUWCTa
CDl+6oJnUk3174B+ebSPCJwvb+BrsMITYkJKbGWtz9qnM7K0nrjA0J2VvskrACXF
U+GXcBP0Z7ax3ftx7jEREBB+uLOtM02ZaflDxUuntZ4i0ACpJyHjz6EwrH1IajHO
GwCuXEnQoBd8wW2U1JzBh+3oJRkeN0vQ59G/IfQybbxnC9MnFTU+9Osu5/hjLiq4
tE6J6p6/ed2cR/orXpJFoKJn1GjUgavSY+3x8UfIrm4dWyI6KoK0hOZ0BxmGSyir
Ffygg7LhyR+i0fzAX2qHecjGL6QOONsely1FSyHoIfvdJCoRcNIQAee37YDZUXgn
A9iI2EFN+JhvfWWulQPP6xAAut3AwXipLnmC3IPkh/ydiPPXDRysEBEtQKXHpZUG
2S7RN1G741hGQcV/FBanlWCg8k/jFV9WtpnG8eEoj42JTPMIhS76OaMdx9X4h9+h
BLWUPr2PpePhu7XUrceTJxd6bNYSABKLdRnI8MDVANuMMWexh2U1Ul9wXqXjx2OT
bzqyt9oZmxQnDQT/FH1+995qJw4oznqn6nsr88eg3IDmjMxPciJLCdwWzzT+9aF6
J4I80bC9CHENv94x+hS63KObWS0laVvrbl65VQWikq22oB6IvsrzoyA96Fb8Cgd9
GjM2sNBirdafEsiopVH8chOUKYouAtl33Z7oHZXqjFn7fRybPTESwfhNml/vjdKY
2buROBJWlv8HF9DqiRgS/Zs7oVn6uSyfus8qCPXiS55nJb8oa333Sw2esQyYeJzP
qtYumP0eb6j1qOf2xg9n5ZXoueEN3+2hkOpk/sCjcxmSwC9XX3egezetc66flVId
DBvUcEaEF9vtjXYe/c2qtVDTna6TzEeofjuh0XX5WqGhYNBuIUUvsukQPaiEfRGT
W0PXtvDqtDwBc2sKuTejsLAv4acdTKd0QRMDTxDZCzu0MUcaJYSz0gQW67/rIrX8
EAgnNQgdVckZJJz/UFcXkTDrUN2M65FJrieAsdJtKVVcih6hdDEkrloX1+Turnxr
atnCP7oA1FvmV8b0j74kgSqR9OsI11JhuinBO1bTxf/DfSY8KuW19K0wkCHpi7Dm
0QRwlayrvWFXoe9bWhMDMuW1nKuvPf+nZT4cKRbD70EnSrelBYlrRtL8g3GWUXRP
/TWz8ncRLXFXQDu4ekxxe40c6gSCb7fETFy42HJZbhCNHceT7LhF/cZhqMQka/XQ
vOK6KF5l2E0sjG785njEMjxsnZ0sxvD0NSnagn2KUBF3y2IZh+U4uQzQ7jCZMAIO
nDGwxAKW2Nw3AdkrQugTnKDpioqnbLNhV72Vy0QCMkX8HdUYGSdNQg6eF6GB0PJa
9kjASmPpH1iHzhVnvNhMgyIZ/+JFQxjE8LlDC71nB3iY2uaLEYnGDSKCnbp3cU/c
CW2StH/ayU5iLmAedQtcQghmaa0aQoRfBLynObiH5ANniGKquxmRsoKWOXWtY3Wu
qeyOcQfW1tLR9kzI/oGEipxnLVnzQjLt9PwDFeHMQwJJ36QipMUr7DfM6OYpYZ4T
J4mFMDg+YuytV4oj9H7MV+0PLTx8uDVXAmF8IpNMbaNo56hMtOrjM3+pDKESuNb9
VQJeRZ7tGrhWRK3AYSl7cNw7Ap9gpx4P7I8gSk7uYF6TjulCU6NyS3ucKBRJA7y9
p32/LYa5+9omt7GVky69prlTnBw9w54yT8L4GkBK4UUoFjrKwSULwMwQEM73iAwx
DsLKhh45T2g2VnxftWOIcI/NIMIfdz0BA8ZCHwOMeYvorSYe7blztXdJ3faKLn3T
4CrcYO9mGSRGviq6508ElepqKZha6/enaDRI/TynZxL0Ti7xxfAF46Ozvkn+6vap
/Q5yaE2d5TtxJ8++B7HkRPnGHS5YKRrlvm3kmeAtfkY+K33ghwIqoKHLTt3qwI4n
pTnp4xephCDO4hxV8QzE3srlZYnGBICWNvFmLf+cKDrtUB7MJgYszcdxewz4ZkWa
RYjyO26b4Oep1l6x5vhDUF/gu729Symb+DXPOUoHGSt/u1mypsMLXlphAK3R9oS1
aMC02IvxMgWhfNQIKwbmqRpx9d5so8/ojqHFRE+yKqwrngRQa3VHjJJWuDwqsMKa
t2FDOKOuQ3tbG65edHbqE3iBXY5iWhinatQPa8jPWcz0EpDSeQZdAl4GV1NDxZyG
H5CYoE3+fOBb4Xca/Xnf/I0HhSYXoOLoKcwOMx8et41UhtYFDrLoQenbapZ0s1l2
QxLwpCPKjcXHDxrwJmiIeoy2FxesZ4ovnl4hVUqdjjmnaqdW7fT9sKzMAe5/k5jz
zzQ9T3c2L9LdmTZSswMONMUVjenOu1wpScgZrlgeaZhXR9U0WBTEJieghWziqHhz
MPS3kmynatLEkbPblyDmpqUfPwkZ0YmOSSdgu3socKRrzz6qMs2jO6Ka1USHXRDX
NwHhxeYvCxMu5Teu7z8yQgyZdhT49QZIXigzL+aEEu9xRy9M2qlzZZLd43bSIuLK
IX2BpDYHd4XVti4/8301c/n+PHZDtg3Kt/9ygJsrHzfc4xnnKgDX2bKXpYH3Wd4y
xkFel7pqgswYNke40Zq5hT4e6kqUwMwL9xUPrAMSOFAfn4lSYMVbQUXJYrGiD0pU
QlKumyYBwx9llvZAeZYEQKWLCbXn5gcaL4X4oGNhLSBxtur63SAx8cnTU8aCN/gH
uXenJnwqjbn7ExTMzDcuV91+RJLI/BBXqUPYMLTBzyu0PDi0JzMiAWL8QlyYe8ab
PWcq19UOD42/57pSSstRgbu+HQH+vr080jVG9hQfDCwXbK17/N0LX+MyqwfHzH4f
eIjGVeCyUy0hHShTcxvz29mUrVlp3Wte9duWEefiLtLxT8YWD97Ko5EXc0+TxEIC
l7eDeCUsdBzrdX5afkfHcvTe+gWgPROg38O2GKPJcidUxmsuR/PIjlA3+VJaaZjB
I3DRxlE3NiDG8FO6zJVs05VexsWvYw+wGebRDtu3UJ8+xMbpT85aCu+8UaF3JYSy
eO5tJoBiqz2A4J3z0fsr9NBo/J+2rAxOPFjumiWXZAD+suXoN3S4EAZKRYaQh0tK
UBTrzEz9w0XtS9sWVw6NRtcbfCrc6un+TgyoppNmj55iO9zd9VDqCmPBP19J5ig7
ksyXMI6TaFV1HR+6HjJBLXKsSuW8RlBU6XP5/2kZePT9Gesv5cliU5LySwgH9nU8
W6CYccLgR3tnerrcJHzw4GpwPzRGsKmQdG8F2tceVbN4YSIVJEVyCVM1BsQzjXQ+
A90w1aEtycmKQaQNUMowkMu95A+IUx32icTzBhK7lkqf5HxsOY7WqbL4NKK7ZLs7
eXXGMC9cUo6aDDp3DZr8Xi7LJPgXkxKlNIXnca5LfsPjyQlDCmp/bFSZy7qjD9ZR
HhlbymJxVBPKJcntdniyXXGJHy7JiGdmU8meR0guB77R6YNb6zcw9MyPkJBgfpdo
7ta2x5nmSN5lypHY83iqJjjRzaVbZ6etLoCXMkjBfpzYmG0K0V2luLuN0AMMMQ/C
4gARAPH6mVhXq1EwgO+yQWOpoh5XvgPSfSgdOJ8K3TL34HRSWB3iyqfAncNVWcLF
6d+9nq/ts46WOwJYmtaAuCMZuMuxHGZy1h/lZo4jzmuDLXbOUyIgueUE1fEofKdF
X8dki84WNTp2q6x1s4S0/Sgodr6N2kzJbTSo+ULtT5/xN35RJkReFPOyI1W6UD7L
pa3HyiZJ7o79JqwxCQvSwOoyDBzHd0FEILDpnP0p6fC1YfRJcmsJvB8GwJrNgImh
YjCYmssjbg6smLs+utihx/5+/ZN0sflk4HUMgkw+y4o5zaGO047ZdeB3Cw0Stf7w
bS+SKnvq2QUJOL/51twaD+u57sCbAUUb+drtMDExUQa3I4U2v5k0ofB6HpqAUcBY
h1QtFWVV70gCs4zUgucd2zkMBBqSu9UuxEy45EjO41Kr5b7SkuWSMd6j2tfRJbaM
GGd6HQTmp9fGpgRnIQ5rKwMxBVFq9SXGemD9ek4skt7xbtH98SD+jL3VqRvgJDOt
PcnIie3Lwce12GmWfRWsik23cfo6oSqielWbmOoo+gPl5veFfD7mRC8n8nZS+HZ4
ArcxvBULI64jlQdk1S/zUUiBx54bLUpHCRS3gONf8KqSNwFS4TDTvNPBmOIKjDjt
N5L4C5mirT6QYnqmf6WsUCagJgj1h653D8f8XyXIDuS9I8ocduMcKM6DeKytsm86
IK3//3CW0SQff0nKlFxKyTJk/T+AQZegC3KRlpqxF5hBNxJ67v3c5Juqr8dA5txM
m3FgJAFS9pkQou5x1sKXklO+Mg3lV7EcrxoguaEWJcRXcCg80rlHX/opZ6rbVdVT
XBcrb1yK9f8oB+IIs9gV6ssrHsDJZyL55vsIxv+RGmYitw3GFjbgrWMpCpchs1mb
5wZ0zQZovIW4EvXsn9rEZP9ezkywBfaXFKtVFnkrkEQdys9dr9Iggphb6rPydS/k
rMwdzMieZrbl2WDlMIbhVoXZltMugvufrQKgrmXe/3Th/jHoP88XaMmEMFjG30ap
8uhk1RMiewbhEC8hnerZQNhZF7HqMqix69HYMgdeOM5XB8U6M/vlf5/1uJJIqwQE
skjbBRcvpjF61WHLvJmNJaKzNBC8BtWjFqe4L28EDPQvRvs9vAPnnp/YNEWZp7or
DtIRmZ9qosRxUFSIsLb3VsQrmuDfe2GDYLffassytitI5d+5Xm1MdHjUyYOUT6BQ
NrrAQUGkUlFxrQbxFvxdcXXRfscEehBgur6j5JWuIkho1EvMbsGdI+2RPbdh1nNf
h5hmxdP9sVYuqHeGE4gWHCOvz9BG0KSjk1neNInpdxhSwuDUH/FQ6aZI9+P3mMf/
TNOkXRiYB+xKzkfWe8ehaulkUjGSUxNdeLVNJAGBxjR7o+uVRguP71K8iD2Zi9nk
C0dlyqQNs5RdjGcU74Z7I1MiS9gMbsPjyfdN3EsQzhkA4XkeyGLOkVoeEYVkY8Bn
p5hSkvPOVAgF2d3homP78YUcScvjoR5qsGTrUSsHbHFn/yJaN0B8GmVNICfeJ060
9VqyPmQFQjVp11gVvRrCk6PkDbtezK81klAyJar2TRnJn2jT1yarZ5diIS1ovhCs
CDEngtlAaa8b37dcI1Rd0Pg5NsPhz+kC1qBOaecTrW/0PiH7XwrL1zBtZAsQJmMt
69rnKe1k44qhWhmCtkSvcyBqpzxB7znfQ1jyJOk+gF+bfBOS0gdQKodecT76W0ip
w+CnNr0r667BsOBbEzUOKKg7+fua6TuDFK0/LILU5FARjNzKbYn0T2ckGkwF0ROR
cx3zJ2UlBmc7LwvbgEDxW8Zb17Uf9vd4cMhtyhVMshTlOhF5CaKqPeQ6rGE8XyUe
eudsYnqsZlSGg75OXEAY7zBkpbV5yC9UWPGsvcdTK9eZdcdCUvSsYGAkEvKVidkc
wIfXR6pgeNnWKXDNUvoxMHHBhL0sdUaGNeHpAax7F7iqn+70C3NG8zZsRxPXmc0b
SH2CqxICAZpsV3zN6M0d94CUF1JKqEq85A8I7JNboIj2xaZPeKZTgDMZGZwdwTey
z+rKcZSbK4R7ZttLCn9iBzkSWUU45d12xDRM7RHe/8EKhJOVZ8rKz7GW06M1EVyM
r3L4WrCwjAdglweova2FTPd1CdQestB6PGuC1RE/+0FuuGcTUIWVzoj5uxe3jPc7
ZDX9o6DtOv/fT2UXa0C8YrBcl953vun5tQmI4q+NdDEcT/rrvgV8qyRvs93p93cb
rpSOkWcIPjZipLi5rSI0M9hTm2fnJHvGHUne3veKqC0VfauyBgepFUTdnV7tn7hf
RFNJ95HTN/ldyVQDdt7clifA3E1ojT6o1tip7fH0HCmtnIc98uPaKXRDbnT6JtFq
qTks6j7fA0JPpOILzJUwsKn7LiPx1WfCx0XJxwAYUU4ibq9v9jcqj8dh0xKjLcFC
QayPuwJCoiclyel7YzRw6uTB2WdrM0n3HkIgQ+xaC+pV5oPoYqA8OXN2kh6bHGXf
+bkNjBXJeW+aRxZIH5HVTLubWnGOhXI/FO/yhxg99kcY3+cm9vsxizKxaVbN6MHE
Dj6E584mM/BGkUEeRRqxnhKe1wsxR3bMPvqSIEYk0AjXNb1DAYJqtug8Ocv9R0sm
npOzVVUQp040QzkuqIpjexNhEhU2/KcEqAm1xpd/eZnOIFo63e/ZNABKHCMmCHP+
zRCasPBMbtIsVmU+OQiycrxX6DxYUigduqY+WZgdz7i+412tvgMIQJllMUm+d0RT
LJrKJygI9QU5jikQ30MMGk3/+KCPIRGBd+vRah6YIeyuPAc2IVkalpdf1FtCKGpf
AYWQRRIJIiiNf3z0UpCGa9ltOYZ4CEgJbZb6ULM5bqVWGGQ6xnhYs6G6KNcRjdw8
`pragma protect end_protected


`ifdef SVT_AXI_QVN_ENABLE

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
GKeqfb7OdtdzGRg/VaX9hhcoeoFUGXiQBkra0LOGUXnY2b4DhzRRxeveLujs4vsg
mwcnrHSMucoFQFXvOS3otg3aEY1PdF7G6BCviNUCfmNORUN/zse+w3Gl5j/fGxNo
5eVg7+6zSbJxp+ybujzU+nirdFJnrjVMgGz1XdeROPk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 43498     )
i59I81hb6jVmO5HkrglO26l4Kb/sJM1VcOlO3nTmL1brsc4Dv9oBfg+rgRDvB9eg
Ha/zLJqsk57/PIK+uY6FA+K/XUIrWLAgp3R/Efs0uQEebyuClGR8NxRzVvSmpob5
im1OxRYxw0ZpWoZlazbYysIE9LcSgu6DMDqh91qNVWBU61kfn+5/z2ndkoRcd+Rd
Q/bcnuHYq91+JS+4xHq8OGoxRffIEaoRKrBbndcqcLXIEFS7emIKX2iUa2MK6bXN
hC/eblSgbmkzVppdsdEJIvLKdhTAe3yG7gmdN4lvhfF9IsZn91pe4lz08PJw+4DQ
IJPp2eaTUJZ8VhtMAv/vbxMTMVd2MEWQ8zqQxQZTIrHmvNj2dvq03NlzfpfXfDvn
V7njdj9mqapCZV8Th5SBLjPUfveRvUWzlfM/CoUmC7JFrBA/roMDAnBF+95kuh7q
JtyhJ/Q/i1E/nwfWUoFfAyFcpbom4yT7TxAIHvIbf+tEVoAoDdb0DHB8a/oLSuH6
J/FeQ+Z9xfDPD6mLy8gHp2ZII+HvFWXAgSBbO4gEYSabRkrJfvfADhF94fh/qlFT
mEUF8XNDd9fK6P/5/s/2SNx98F+P711/oXsWBimbowKMF17Mqtdn0/dlJcPA7R5G
qFZgtBatCeMBKIMtRkS/6feJYy5k07VnONvmERjuyIC1fec4BjD/A3bOkFMo2NV7
CW9X48rSM9UhXtifQr3XN8N75S53bQ47goa8dE3RXWI9DYbwXU74pTnsJV1k6h4b
ZhUtt7nPpq+K8WJ8RajovvkFlEAdqFGfFFxEOvN3xpLz8jXM7O72yFKZr9B3o7v1
/bEvwvUMmRE34ap2hJ5ZY6LeIdwKHI+Nv1S3RhOiQPyjjp/eOrBaeK70whQmgBDR
q2gsohC3MrRqagwBbcZsV417pIY5j4PRXADusmeZfIPRibQlWvvmLI4Cxv7K2D0u
UqMfdBtBpDEPh39dfW2bso8F4umSF7tN9pkhmaukG8mpvrv2QDBeGV37LKKZUYrs
HqMmjZ0QWfB8CiZCz3WX4+8fNopKo+b/ORqL4SX/0VncSOkJPM3S/4rt4NZuUjjM
x0MSpcvf+MvaFF6ik+YJhZaAeCUgTUwvClEgQ6IOEuE729SLAEb3TiSdyFd+o3xj
AWUUmvQhcLwOKuniKF7+h1tnzi6x8VfswHAUbM9VSXoYTxmxSlRwWgvjwIHjzJ4r
A+dhLI6PQLLIaEKOsfuLgUwALk2QnOb26l67wXoO8lM4/pxSnv3kjcw4K0hQkxW2
b6NELU4qzoFqkb44uoCSnropsom7FUaPk33AUPa7JVU+icrwuEYrN3Wc7GKJb0u8
RfMqYiTo0ysGNJEyWyebcec7dq5iVeW6H+kaoWJhDtzh2oU5n5DNgXH7PZ31KhYn
OUuv5G1Vf5HjUoM2giNGb94GGffeSJP5R9RXfUy/mkRA9svuvq7zwZMMcdr2PXZq
u22EELJ1colkiwonFYzFu40XyJGHRkhFRAzD9mLcKp8dBF7wvX92bVCBYIdG/E0z
eMhzodwvOR7eYtaT3cHWB1ihe2uSEdL3XHBaoeMYSdK78ZIVz1PymXbpoR+PWB8S
t+hgooSCWR+m3AFWYYwbWv0hB50jkc4ePiBTYXmJn/wjtCg09U7OpTW+Z67c4b0v
tqsi1BCQydpKV28RZ6XGhPr9Hwu5Kxes1umt+udGUaeNJtT0B7zY4EjyYV174qa4
LbYqV6p5OzKDKhyCG3mN5TD5ppGu0CO34NKWHVTxZDXQY3bpgJHG4CJjfDF3pgyL
jsmtMa049x5QNPdsxAjOm6klnDX52W9ZQCdIT8GJvt47ckJTivMYZjFbrKenX/AH
S2I1mRe5E5fv/OZFZbiASQ5hc2sJcn01rVryP++eYxMWKTCosHZEz+exctVaHQNY
4U9XwwSXS/Kf7GDmQpQcEoP087PUXOe+9h4c+4AxcRPlIh9SMa+fhf3VYWaJlzjj
blYeoflimHXUui3W6FpoeDDFvunUZGjNE07yKpUNU3911jjqNam7jpxy2HbDkIDX
YYz773cB761/+hSMpDc2pIgUZCwb1F1NowvvyuR847Axa7nV5i80XmymWL6Vkmnp
qlWnChCw+c39qDsGDrJzi9UQ4pFlTIFGEseudwrSvSwSj0R9M4zms1qehqmQcWOw
+xcJO0E85ns/m3Fh6WDZheSQbqgOyTTWbDDrzKdSDViTEA3sT40a3o3PD5ahwhvd
j6/xMeZNMbQZGmjM7bkHI/+sON4l1ZdEYU+S+1luLN5v6Sa2bqFBHT0+vqlZrLGM
3HW7RuTxtLabMev+gqVvT5d8faRBGjUlO5I+PB96SBGXkxToyRH6e1bFw/0xPuQt
doQVv+fBx/sxe34nzmaU+OFywK9FA0pnKLyPoTYHTJEwPWX2i2BX28Fx5Rox2QJ6
hoZE2c+/CL1vtlUXMLlJqj1Ufmcj73AW3nR0hgrVkAnMm/w8oyEZ7OENIpCeJ2+v
Ntgzg2dZR2uFBRK0nx8yEFpQHBP4osm26sI4wVhhrcURX/CtggcwDAz5ADiwLp5r
vpw9Tf0o4d+6hkfYPAJepimkUf63rbjBpAuBGdXxNHwJAvSJ4izhRtQ5ADyTDMVE
lfDobpoIj2KnRwcuua8WSUTEmCuYLm6Y6G41q8nNcG7JkrDt0qlK7ZhWEnNls7CD
qlUSxGKiqkBGxKT1DR7rFjuRawJpb+epHjDMfL0Phfg=
`pragma protect end_protected

`endif
`endif

class svt_axi_checker extends svt_err_check;

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
YxbfNg6F8JsmFBZTBuO59rrJPUSzhGqdIkdP3N3X0jDb0kWv4fvJfZF8emI2iJal
HgZ+/9RIM1TUGd8KMoMlQ6l6mIleLXEdHvPSPE/q/SBpLkVxpYbLWJ+tvAAydiy3
wAn6SiXNqcTweEWQyZepREu0I6/0h7zLQVsaSK/DyOc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 43698     )
Q0zadrpobcYAYv9GVnUZNxkvURFeoC0UYMLgyoi94X9TXriK7FXUytIQZhjPvN05
Umvy8p1u6i2j7hEe6H4SohCQp/D0/er6ziwQYylhyOoOzManZ8xwZmphx3tGfzbZ
8lFsXdcLoiOaYNXLophQv5e1I/96JnI4JetnHrLNwP0Na+1HBs2GCP9KItgFApnW
4thIM1DLT5XctyO8+lryT0+4lvaB/HeXWJoQ9xvBe0hze8ZtqIrzueY9fN5Jh6up
m+/1NAIGIis+eaKZc081RQ==
`pragma protect end_protected

  /**
    @grouphdr port_interleaving_check Port interleaving checks
    This group contains checks for port interleaving. 
    */

/**
    @grouphdr trace_tag_validity_check trace_tag related checks
    This group contains checks for trace_tag feature. 
    */


  typedef enum {LEGAL_TRANSITION,
                ILLEGAL_TRANSACTION_START_STATE,
                ILLEGAL_COHERENT_RESPONSE, 
                ILLEGAL_COHERENT_TRANSACTION,
                ILLEGAL_SNOOP_RESP_FOR_INITIAL_STATE,
                ILLEGAL_SNOOP_RESPONSE, 
                ILLEGAL_SNOOP_TRANSACTION
               } coherency_error_type_enum ;


  local svt_axi_port_configuration cfg;

  local svt_axi_transaction barrier_xact_queue[$];

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
enY8hsSH0In0zpnTPOKHArfZgKdb4+9jP6I1EyYvvRoQjdEFZ3dYtZPojbV7bd2N
UHEN3XbClSJvTMfJRXnYWAjUlSgjth1c/TKAdSTYzs6kO4FMhj87ZIBPacbax2sC
WnnXYFgGcPPIlRdNg/43dGEJOjCQ7Q4iZL49hG04hhQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 43821     )
bb8HobQKmfPfx5W+8Nxn6cuaiNZkl6rBiAlRW3wDBlD7Eh7Bx32EMXhfJokVVKEP
8Dd0dp8aQZCaSldBgwrhl1OXgpibTAAt8PZdvWXJTN4MA4OP5iZtVcjbxqTV+aAj
sqAU7mutABzKoOmUoDjaGhAzvXYiVDrPsWCNTehJCF4=
`pragma protect end_protected
  local string group_name = "";

  local string sub_group_name = "";

  /** String used in macros */
  local string macro_str = "";
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
JPf3Fkz+bv2GbS1q+x/ESJUHx4X/qqOxNxnQZP32RHp4XT99lq0QFJvcma1Y+c4d
WOfBDXUapmVNKBwfYiyO8E/4vGYVqVuN/LkUZrbkj82g81DbjYXXa/lL6a3xSVDC
ZgjKsGOX4DhOmoByapxFMqUo75/xEwjNY1/+dQW0sSw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 44152     )
Q+IV+KDSoy6QTDZCqBqbzzNf2GD4rKBvWFvP5FHXPW+sFqVCe0KFXLjR4B3FwJD6
ZWvEHH8/qniID4bJNn1b2XKqtuCD6J6nYENIbP2cT3W+k676DIahq3ymPLqQaWUU
vqWIFXeB/k19JjxsG82/aBdZLpfmOtNMm79gzhnEbs3D76xh3DnwCFbHEei32qub
Xw8+4XItbmSdOySGqO1t4S0IdJf41xlzoeClS1Dqgx/bgnM0LKG4QkhljQuueeHK
SctPsXCuyiQmV0X99lIai74dlZHJa3Lkq1leEOa4Hpp+6n1yuwFhAbYySKgqbm/7
oPIIYwcbb7NZm6rqhMqDbgjho26Psak20g5w57rjdWyE9uzkFmBZNsmS0r0LGTB2
VcaOUG3APeqmOrwJuKJpHx5IpqNlHRDeAeTyipsd2+bOMnGMMieLxHYA7BHvGnGq
`pragma protect end_protected
  logic previous_reset = 1;

  /** Delay from ARVALID assertion to ARREADY assertion */
  local int arvalid_arready_delay = 0;
  
  /** Delay from ACVALID assertion to ACREADY assertion */
  local int acvalid_acready_delay = 0;
  
  /** Delay from ACVALID assertion to ACREADY assertion */
  local int cdvalid_cdready_delay = 0;
  
  /** Delay from CRVALID assertion to CRREADY assertion */
  local int crvalid_crready_delay = 0;

  /** Delay from TVALID assertion to TREADY assertion */
  local int tvalid_tready_delay = 0;

  /** Last sampled values in read address channel */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_arid;
  local logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] previous_araddr;
  local logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] previous_arlen;
  local logic[`SVT_AXI_SIZE_WIDTH-1:0] previous_arsize;
  local logic[`SVT_AXI_BURST_WIDTH-1:0] previous_arburst;
  local logic[`SVT_AXI_LOCK_WIDTH-1:0] previous_arlock;
  local logic[`SVT_AXI_CACHE_WIDTH-1:0] previous_arcache;
  local logic[`SVT_AXI_PROT_WIDTH-1:0] previous_arprot;
  local logic[`SVT_AXI_QOS_WIDTH-1:0] previous_arqos;
  local logic[`SVT_AXI_REGION_WIDTH-1:0] previous_arregion;
  local logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] previous_aruser;
  local logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] previous_ardomain;
  local logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] previous_arsnoop;
  local logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] previous_arbar;
`ifdef SVT_ACE5_ENABLE
  local logic  previous_archunken;
  local logic[`SVT_AXI_MAX_MPAM_WIDTH-1:0] previous_armpam;
`endif
  
  local logic[`SVT_AXI_ACE_SNOOP_RESP_WIDTH-1:0] previous_crresp;
  local logic[`SVT_AXI_ACE_SNOOP_DATA_WIDTH-1:0] previous_cddata;
  local logic[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1:0] previous_acaddr;
  local logic[`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] previous_acsnoop; 
  local logic[`SVT_AXI_ACE_SNOOP_PROT_WIDTH-1:0] previous_acprot;
  local logic previous_aridunq;
  local logic previous_cdlast;

  /** holds number of databeat transferred over snoop data channel for current snoop request */
  local int unsigned cddata_beat_count = 0;

  /** Delay from RVALID assertion to RREADY assertion */
  local int rvalid_rready_delay = 0;

  /** Last sampled value of RID */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_rid;

  /** Last sampled value of RIDUNQ */
  local logic previous_ridunq;

  /** Last sampled value of RRESP */
  local logic[`SVT_AXI_RESP_WIDTH-1:0] previous_rresp;

  /** Last sampled value of RDATA */
  local logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] previous_rdata;

  /** Last sampled value of RLAST */
  local logic previous_rlast;

  /** Last sampled value of RUSER */
  local logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] previous_ruser;

`ifdef SVT_ACE5_ENABLE
  /** Last sampled value of RCHUNKV */
  local logic  previous_rchunkv;

  /** Last sampled value of RCHUNKNUM */
  local logic [`SVT_AXI_MAX_CHUNK_NUM_WIDTH-1:0] previous_rchunknum;

  /** Last sampled value of RCHUNKSTRB */
  local logic [`SVT_AXI_MAX_CHUNK_STROBE_WIDTH-1:0] previous_rchunkstrb;
`endif 

  /** Delay from AWVALID assertion to AWREADY assertion */
  local int awvalid_awready_delay = 0;

  /** Last sampled values in write address channel */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_awid;
  local logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] previous_awaddr;
  local logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] previous_awlen;
  local logic[`SVT_AXI_SIZE_WIDTH-1:0] previous_awsize;
  local logic[`SVT_AXI_BURST_WIDTH-1:0] previous_awburst;
  local logic[`SVT_AXI_LOCK_WIDTH-1:0] previous_awlock;
  local logic[`SVT_AXI_CACHE_WIDTH-1:0] previous_awcache;
  local logic[`SVT_AXI_PROT_WIDTH-1:0] previous_awprot;
  local logic[`SVT_AXI_QOS_WIDTH-1:0] previous_awqos;
  local logic[`SVT_AXI_REGION_WIDTH-1:0] previous_awregion;
  local logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] previous_awuser;
  local logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] previous_awdomain;
  local logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] previous_awsnoop;
  local logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] previous_awbar;
  local logic[`SVT_AXI_MAX_MPAM_WIDTH-1:0] previous_awmpam;
  local logic previous_awunique;
  local logic previous_awidunq;

  /** Delay from WVALID assertion to WREADY assertion */
  local int wvalid_wready_delay = 0;

  /** Last sampled value of WID */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_wid;

  /** Last sampled value of WDATA */
  local logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] previous_wdata;

  /** Last sampled value of WSTRB */
  local logic[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] previous_wstrb;

  /** Last sampled value of WUSER */
  local logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] previous_wuser;

  /** Last sampled value of WLAST */
  local logic previous_wlast;

  /** Delay from BVALID assertion to BREADY assertion */
  local int bvalid_bready_delay = 0;

  /** Last sampled value of BID */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_bid;

  /** Last sampled value of BIDUNQ */
  local logic previous_bidunq;

  /** Last sampled value of BRESP */
  local logic[`SVT_AXI_RESP_WIDTH-1:0] previous_bresp;

  /** Last sampled value of BUSER */
  local logic[`SVT_AXI_MAX_BRESP_USER_WIDTH-1:0] previous_buser;

  local logic[`SVT_AXI_MAX_TDATA_WIDTH-1:0] previous_tdata;
  local logic[`SVT_AXI_TSTRB_WIDTH-1:0] previous_tstrb;
  local logic[`SVT_AXI_TKEEP_WIDTH-1:0] previous_tkeep;
  local logic previous_tlast;
  local logic[`SVT_AXI_MAX_TID_WIDTH-1:0] previous_tid;
  local logic[`SVT_AXI_MAX_TDEST_WIDTH-1:0] previous_tdest;
  local logic[`SVT_AXI_MAX_TUSER_WIDTH-1:0] previous_tuser;

  `ifdef SVT_AXI_QVN_ENABLE
  /** Variables used in QVN token handshake signal checks */  
  local bit is_varvalidvn_deassertion_check_en [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local bit is_varqosvn_valid_change_check_en  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  local bit is_vawvalidvn_deassertion_check_en [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local bit is_vawqosvn_valid_change_check_en  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  local bit is_vwvalidvn_deassertion_check_en  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  local int unsigned qvn_ar_token_request_ready_timeout_counter_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];
  local int unsigned qvn_aw_token_request_ready_timeout_counter_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];
  local int unsigned qvn_w_token_request_ready_timeout_counter_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];
 
  local logic previous_varvalidvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic [3:0] previous_varqosvnx [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic previous_varreadyvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0]; 
   
  local logic previous_vawvalidvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic [3:0] previous_vawqosvnx [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic previous_vawreadyvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0]; 
  
  local logic previous_vwvalidvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic previous_vwreadyvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0]; 

  `endif

  local svt_axi_snoop_transaction  multipart_dvm_snoop_xact;
  svt_axi_transaction multipart_dvm_coherent_xact;
  local svt_axi_transaction        active_multipart_dvm_coherent_q[svt_axi_transaction];
  local svt_axi_snoop_transaction  active_multipart_dvm_snoop_q[svt_axi_snoop_transaction];

  //local svt_axi_snoop_transaction  multipart_dvm_snoop_check_guard_xact;
  //local svt_axi_master_transaction multipart_dvm_coherent_check_guard_xact;
  local svt_axi_transaction        active_multipart_dvm_coherent_check_guard_q[svt_axi_transaction];
  local svt_axi_snoop_transaction  active_multipart_dvm_snoop_check_guard_q[svt_axi_snoop_transaction];

  /** Enables protocol check coverage provided it protocol_checks_coverage_enable is set
    * in the port configuration as well. If enable_pc_cov is 0, then protocol checks coverage
    * will not be enabled, even if it is set in configuration
    */
  local bit enable_pc_cov = 1;

  /** indicates if only partial ID bits are considered for exclusive transaction */
  local bit partial_exclusive_id = 0;
  

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Uu11ooNgIuvpKigHmtAuf/kh+nteq63ZRYzxHb1oN+DYSmNRdu9eN+fhaH7RwlHz
Jo+okXiIYjmI8EkcEj2H+P7Lbr3kEmhxi54yP+SuPAXDsYhsVC0wYaeGt5lWTGA5
Ip+IjV2LIbeB3uhLSxn3XwDCK0MwBYzIaeAxdqVQHTA=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 44354     )
OqvMue0doqVEw0fo4/VvnKjAZHYrjs0srdl69EbQHloBTfzljgXgMGxbiy4UQSyP
SWqB837JsQs/BwmAZVj8lBivKnst+w7TZcCdMKOU4cSqO3BbEQ/hZTNhEbthsPjh
9VF8Lx98M14DxyySTCRDfMnBAoXPNpYgSO/Pg+LXre5YajKI3JHZihmr2ubXbw87
HOHGor7RoievnDNJnSIxu+V9DXFBzMNMHmqlNm8L44E9gxEZ61uWRfQ2cSj4GGw1
FKOWCpJhpwZhgpVnltxpJw==
`pragma protect end_protected


  //--------------------------------------------------------------
  /** Checks that ARID is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arid_when_arvalid_high_check;

  /** Checks that ARADDR is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_araddr_when_arvalid_high_check;

  /** Checks that ARLEN is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arlen_when_arvalid_high_check;
  
  /** Checks that ARSIZE is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arsize_when_arvalid_high_check;
  
  /** Checks that ARLEN and ARSIZE are valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_arlen_arsize_check;
  
  /** Checks that ARCACHE is valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_arcache_check;
  
  /** Checks that address is aligned for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_read_addr_aligned_check;
  
  /** Checks that AWLEN and AWSIZE are valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_awlen_awsize_check;
  
  /** Checks that AWCACHE is valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_awcache_check;
  
  /** Checks that address is aligned for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_write_addr_aligned_check;

  /** Checks that address is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_addr_check;
  
  /** Checks that received write data is not interleaved beyond write_data_interleave_depth value
    * An error is issued if write data is interleaved beyond this value for Write data interleaving */
  svt_err_check_stats write_data_interleave_depth_check;
 
  /** Checks that the order in which a slave receives the first data item of each transaction must be the
    * same as the order in which it receives the addresses for the transactions for Write Data Interleaving 
    * transactions */
  svt_err_check_stats write_data_interleave_order_check;

 /** Checks that id is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_id_check;

  /** Checks that response generated for exclusive load accesss is correct */
  svt_err_check_stats exclusive_load_response_check;

  /** Checks that response generated for exclusive store accesss is correct */
  svt_err_check_stats exclusive_store_response_check;

  /** Checks that master does not permit an Exclusive Store transaction to be
    * in progress at the same time as any transaction that registers that it
    * is performing an Exclusive sequence
    */
  svt_err_check_stats exclusive_store_overlap_with_another_exclusive_sequence_check;

  /** Checks that, once a master receives successful exclusive store response EXOKAY
    * from interconnect, then no other master should be provided with EXOKAY response,
    * until current master acknowledges completing successful exclusive store by asserting RACK
    */
   svt_err_check_stats exokay_not_sent_until_successful_exclusive_store_rack_observed_check;
  
    /** Checks that READ_ONLY_INTERFACE supports only read transactions 
     * Applicable only for AXI4 VIP
     * Passive Master,Passive Slave and Active slave will perform this
     * check
     */
     svt_err_check_stats read_xact_on_read_only_interface_check;
   
    /** Checks that WRITE_ONLY_INTERFACE supports only write transactions 
     * Applicable only for AXI4 VIP
     * Passive Master,Passive Slave and Active slave will perform this
     * check
     */
     svt_err_check_stats write_xact_on_write_only_interface_check;
     
     /** Checks that READ_ONLY_INTERFACE does not support exclusive access  
     * Applicable only for AXI4 VIP
     * Passive Master,Passive Slave and Active slave will perform this 
     * check
     */
     svt_err_check_stats excl_access_on_read_only_interface_check;

      /** Checks that WRITE_ONLY_INTERFACE does not support exclusive access  
      * Applicable only for AXI4 VIP
      * Passive Master,Passive Slave and Active slave will perform this 
      * check
      */
      svt_err_check_stats excl_access_on_write_only_interface_check;
     
     /** Checks that burst length is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_burst_length_check;
  
  /** Checks that burst size is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_burst_size_check;
  
  /** Checks that burst type is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_burst_type_check;
  
  /** Checks that cache type is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_cache_type_check;
  
  /** Checks that protection type is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_prot_type_check;
  
  /** Checks that exclusive transaction sent on AXI_ACE interface are
   * only of WRITENOSNOOP, READNOSNOOP, READCLEAN, READSHARED and CLEANUNIQUE type */
  svt_err_check_stats exclusive_ace_transaction_type_check;

  /** Checks that ARADDR[2:0] for multipart dvm xact is not other than SBZ */
  svt_err_check_stats signal_araddr_multipart_dvm_xact_check;

  /** Checks that ARBURST is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arburst_when_arvalid_high_check;

  /** Checks that ARLOCK is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arlock_when_arvalid_high_check;

  /** Checks that ARCACHE is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arcache_when_arvalid_high_check;

  /** Checks that ARPROT is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arprot_when_arvalid_high_check;

  /** Checks that ARQOS is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arqos_when_arvalid_high_check;

  /** Checks that ARREGION is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arregion_when_arvalid_high_check;

  /** Checks that ARUSER is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_aruser_when_arvalid_high_check;
  
    /** Checks that ARDOMAIN is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_ardomain_when_arvalid_high_check;
  
  /** Checks that ARSNOOP is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arsnoop_when_arvalid_high_check;
  
  /** Checks that ARBAR is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arbar_when_arvalid_high_check;

  /** Checks that ARREADY is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arready_when_arvalid_high_check;

  /** Checks that AWDOMAIN is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awdomain_when_awvalid_high_check;
  
  /** Checks that AWSNOOP is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awsnoop_when_awvalid_high_check;
  
  /** Checks that AWBAR is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awbar_when_awvalid_high_check;
  //--------------------------------------------------------------
  /** Checks that ARID is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arid_when_arvalid_high_check;

  /** Checks that ARADDR is stable when ARVALID is high */
  svt_err_check_stats signal_stable_araddr_when_arvalid_high_check;

  /** Checks that RACK is asserted for a single cycle */
  svt_err_check_stats signal_rack_single_cycle_high_check;

  /** Checks that RACK signal must be asserted the cycle after the associated handshake or later */
  svt_err_check_stats signal_rack_after_handshake_check;

  /** Checks that WACK is asserted for a single cycle */
  svt_err_check_stats signal_wack_single_cycle_high_check;

  /** Checks that WACK signal must be asserted the cycle after the associated handshake or later */
  svt_err_check_stats signal_wack_after_handshake_check;

  /** Checks that ARLEN is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arlen_when_arvalid_high_check;
  
  /** Checks that ARSIZE is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arsize_when_arvalid_high_check;

  /** Checks that ARBURST is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arburst_when_arvalid_high_check;

  /** Checks that ARLOCK is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arlock_when_arvalid_high_check;

  /** Checks that ARCACHE is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arcache_when_arvalid_high_check;

  /** Checks that ARPROT is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arprot_when_arvalid_high_check;

  /** Checks that ARQOS is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arqos_when_arvalid_high_check;

  /** Checks that ARREGION is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arregion_when_arvalid_high_check;

  /** Checks that ARUSER is stable when ARVALID is high */
  svt_err_check_stats signal_stable_aruser_when_arvalid_high_check;
  
  /** Checks that ARDOMAIN is stable when ARVALID is high */
  svt_err_check_stats signal_stable_ardomain_when_arvalid_high_check;
  
  /** Checks that ARSNOOP is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arsnoop_when_arvalid_high_check;
  
  /** Checks that ARBAR is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arbar_when_arvalid_high_check;

  /** Checks that AWDOMAIN is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awdomain_when_awvalid_high_check;
  
  /** Checks that AWSNOOP is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awsnoop_when_awvalid_high_check;
  
  /** Checks that AWBAR is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awbar_when_awvalid_high_check;
  //--------------------------------------------------------------
  /** Checks that RID is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rid_when_rvalid_high_check;

  /** Checks that RDATA is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rdata_when_rvalid_high_check;

  /** Checks that RDATACHK is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rdatachk_when_rvalid_high_check;
 
  /** Checks that rpoison is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rpoison_when_rvalid_high_check;
 
  /** Checks that RUSER is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_ruser_when_rvalid_high_check;

  /** Checks that RRESP is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rresp_when_rvalid_high_check;

  /** Checks that RLAST is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rlast_when_rvalid_high_check;

  /** Checks that RREADY is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rready_when_rvalid_high_check;

  /** Checks that RID is stable when RVALID is high */
  svt_err_check_stats signal_stable_rid_when_rvalid_high_check;

  /** Checks that RUSER is stable when RVALID is high */
  svt_err_check_stats signal_stable_ruser_when_rvalid_high_check;

  /** Checks that RDATA is stable when RVALID is high */
  svt_err_check_stats signal_stable_rdata_when_rvalid_high_check;

  /** Checks that RRESP is stable when RVALID is high */
  svt_err_check_stats signal_stable_rresp_when_rvalid_high_check;

  /** Checks that RLAST is stable when RVALID is high */
  svt_err_check_stats signal_stable_rlast_when_rvalid_high_check;

  /** Checks that sample read data has associated address */
  svt_err_check_stats read_data_follows_addr_check;
  //--------------------------------------------------------------
  /** Checks that AWID is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awid_when_awvalid_high_check;

  /** Checks that valid write strobes are driven */
  svt_err_check_stats valid_write_strobe_check;

`ifdef SVT_ACE5_ENABLE 
  //--------------------------------------------------------------
 /** Checks that stash_nid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_nid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that stash_lpid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_lpid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that stash_nid_valid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_nid_valid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that stash_lpid_valid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_lpid_valid_when_awvalid_high_check;

  //--------------------------------------------------------------
 /** Checks that awmmusid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmusid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that awmmussid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmussid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that  is awmmusecsid not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmusecsid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that awmmussidv is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmussidv_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that awmmuatst is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmuatst_when_awvalid_high_check;

  //--------------------------------------------------------------
 /** Checks that armmusid is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmusid_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that armmussid is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmussid_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that  is armmusecsid not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmusecsid_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that armmussidv is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmussidv_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that armmuatst is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmuatst_when_arvalid_high_check;

 /** Checks that awatop is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awatop_when_awvalid_high_check;

 /** Checks that armpam is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armpam_when_arvalid_high_check;

 /** Checks that awmpam is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmpam_when_awvalid_high_check;

   /** Checks that AWMPAM is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awmpam_when_awvalid_high_check;

  /** Checks that ARMPAM is stable when ARVALID is high */
  svt_err_check_stats signal_stable_armpam_when_arvalid_high_check;
`endif

`ifdef SVT_ACE5_ENABLE 
//--------------------------------------------------------------
 /** Checks that ARIDUNQ is not X or Z when ARVALID is high*/
   svt_err_check_stats signal_valid_aridunq_when_arvalid_high_check;

 /** Checks that RIDUNQ is not X or Z when RVALID is high*/
   svt_err_check_stats signal_valid_ridunq_when_rvalid_high_check;

 /** Checks that AWIDUNQ is not X or Z when AWVALID is high*/
   svt_err_check_stats signal_valid_awidunq_when_awvalid_high_check;

 /** Checks that BIDUNQ is not X or Z when BVALID is high*/
   svt_err_check_stats signal_valid_bidunq_when_bvalid_high_check;
   
//--------------------------------------------------------------
/** Checks that ARIDUNQ is stable when ARVALID is high */
  svt_err_check_stats signal_stable_aridunq_when_arvalid_high_check;

/** Checks that RIDUNQ is stable when RVALID is high */
  svt_err_check_stats signal_stable_ridunq_when_rvalid_high_check;

/** Checks that AWIDUNQ is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awidunq_when_awvalid_high_check;

/** Checks that BIDUNQ is stable when BVALID is high */
  svt_err_check_stats signal_stable_bidunq_when_bvalid_high_check;

//--------------------------------------------------------------
  /** Checks that RIDUNQ asserted or deasserted when ARIDUNQ asserted or deasserted */
  //svt_err_check_stats ridunq_asserted_deasserted_check;

  /** Checks that BIDUNQ asserted or deasserted when AWIDUNQ asserted or deasserted*/
  //svt_err_check_stats bidunq_asserted_deasserted_check;
 
  /** Checks that there is no outstanding transaction with same arid */
  svt_err_check_stats no_outstanding_read_unique_transaction_with_same_arid;

  /** Checks that there is no outstanding transaction with same awid */
  svt_err_check_stats no_outstanding_write_unique_transaction_with_same_awid;
`endif

  /** Checks that AWADDR is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awaddr_when_awvalid_high_check;

  /** Checks that AWLEN is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awlen_when_awvalid_high_check;
  
  /** Checks that AWSIZE is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awsize_when_awvalid_high_check;

  /** Checks that AWBURST is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awburst_when_awvalid_high_check;

  /** Checks that AWLOCK is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awlock_when_awvalid_high_check;

  /** Checks that AWCACHE is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awcache_when_awvalid_high_check;

  /** Checks that AWPROT is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awprot_when_awvalid_high_check;

  /** Checks that AWREADY is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awready_when_awvalid_high_check;

  /** Checks that AWQOS is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awqos_when_awvalid_high_check;

  /** Checks that AWREGION is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awregion_when_awvalid_high_check;

  /** Checks that AWUNIQUE is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awunique_when_awvalid_high_check;

  /** Checks that AWUSER is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awuser_when_awvalid_high_check;
  //--------------------------------------------------------------
  /** Checks that AWID is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awid_when_awvalid_high_check;

  /** Checks that AWADDR is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awaddr_when_awvalid_high_check;

  /** Checks that AWLEN is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awlen_when_awvalid_high_check;
  
  /** Checks that AWSIZE is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awsize_when_awvalid_high_check;

  /** Checks that AWBURST is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awburst_when_awvalid_high_check;

  /** Checks that AWLOCK is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awlock_when_awvalid_high_check;

  /** Checks that AWCACHE is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awcache_when_awvalid_high_check;

  /** Checks that AWPROT is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awprot_when_awvalid_high_check;

  /** Checks that AWQOS is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awqos_when_awvalid_high_check;

  /** Checks that AWREGION is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awregion_when_awvalid_high_check;

  /** Checks that AWUNIQUE is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awunique_when_awvalid_high_check;

  /** Checks that AWUSER is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awuser_when_awvalid_high_check;

  //--------------------------------------------------------------

  /** Checks that WID is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wid_when_wvalid_high_check;

  /** Checks that WUSER is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wuser_when_wvalid_high_check;

  /** Checks that WDATA is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wdata_when_wvalid_high_check;

  /** Checks that WDATACHK is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wdatachk_when_wvalid_high_check;

 /** Checks that WPOISON is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wpoison_when_wvalid_high_check;

  /** Checks that WSTRB is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wstrb_when_wvalid_high_check;

  /** Checks that WLAST is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wlast_when_wvalid_high_check;

  /** Checks that WREADY is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wready_when_wvalid_high_check;

  /** Checks that WID is stable when WVALID is high */
  svt_err_check_stats signal_stable_wid_when_wvalid_high_check;

  /** Checks that WUSER is stable when WVALID is high */
  svt_err_check_stats signal_stable_wuser_when_wvalid_high_check;

  /** 
   * Checks that WDATA is stable when WVALID is high 
   * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=1 ,
   * it considers only valid byte lanes of wdata based on wstrb. 
   * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=0 ,
   * whole wdata as seen on the bus will be considered.
   */
  svt_err_check_stats signal_stable_wdata_when_wvalid_high_check;

  /** Checks that WSTRB is stable when WVALID is high */
  svt_err_check_stats signal_stable_wstrb_when_wvalid_high_check;

  /** Checks that WLAST is stable when WVALID is high */
  svt_err_check_stats signal_stable_wlast_when_wvalid_high_check;

  //--------------------------------------------------------------
  /** Checks that BID is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_bid_when_bvalid_high_check;

  /** Checks that BUSER is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_buser_when_bvalid_high_check;

  /** Checks that BRESP is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_bresp_when_bvalid_high_check;

  /** Checks that BREADY is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_bready_when_bvalid_high_check;

  /** Checks that BID is stable when BVALID is high */
  svt_err_check_stats signal_stable_bid_when_bvalid_high_check;

  /** Checks that BUSER is stable when BVALID is high */
  svt_err_check_stats signal_stable_buser_when_bvalid_high_check;

  /** Checks that BRESP is stable when BVALID is high */
  svt_err_check_stats signal_stable_bresp_when_bvalid_high_check;

  /** 
    * When a write response is sampled, checks that there is a 
    * transaction with corresponding ID whose data phase is complete 
    */
  svt_err_check_stats write_resp_follows_last_write_xfer_check;

  /** 
    * Checks that WLAST is asserted for the last beat of write data. 
    */
  svt_err_check_stats wlast_asserted_for_last_write_data_beat;

  //--------------------------------------------------------------
  // Checks that need to be executed externally (by monitor).
  /** Checks that ARVALID is not X or Z */
  svt_err_check_stats signal_valid_arvalid_check;

  /** Checks that RVALID is not X or Z */
  svt_err_check_stats signal_valid_rvalid_check;

  /** Checks that AWVALID is not X or Z */
  svt_err_check_stats signal_valid_awvalid_check;

  /** Checks that WVALID is not X or Z */
  svt_err_check_stats signal_valid_wvalid_check;

  /** Checks that BVALID is not X or Z */
  svt_err_check_stats signal_valid_bvalid_check;
  
  /** Checks that ACVALID is not X or Z */
  svt_err_check_stats signal_valid_acvalid_check;
  
  /** Checks that CDVALID is not X or Z */
  svt_err_check_stats signal_valid_cdvalid_check;
  
  /** Checks that CDVALID is not X or Z */
  svt_err_check_stats signal_valid_crvalid_check;

  /** Checks that ARVALID is not X or Z During Reset */
  svt_err_check_stats signal_valid_arvalid_check_during_reset;

  /** Checks that RVALID is not X or Z During Reset*/
  svt_err_check_stats signal_valid_rvalid_check_during_reset;

  /** Checks that AWVALID is not X or Z During Reset*/
  svt_err_check_stats signal_valid_awvalid_check_during_reset;

  /** Checks that WVALID is not X or Z During Reset*/
  svt_err_check_stats signal_valid_wvalid_check_during_reset;

  /** Checks that BVALID is not X or Z During Reset */
  svt_err_check_stats signal_valid_bvalid_check_during_reset;

  /** Checks if arvalid was interrupted before arready got asserted */
  svt_err_check_stats arvalid_interrupted_check;
  
  /** Checks if acvalid was interrupted before acready got asserted */
  svt_err_check_stats acvalid_interrupted_check;
  
  /** Checks if cdvalid was interrupted before cdrready got asserted */
  svt_err_check_stats cdvalid_interrupted_check;
  
  /** Checks if crvalid was interrupted before crready got asserted */
  svt_err_check_stats crvalid_interrupted_check;

  /** Checks if rvalid was interrupted before rready got asserted */
  svt_err_check_stats rvalid_interrupted_check;

  /** Checks if awvalid was interrupted before awready got asserted */
  svt_err_check_stats awvalid_interrupted_check;

  /** Checks if wvalid was interrupted before wready got asserted */
  svt_err_check_stats wvalid_interrupted_check;

  /** Checks if bvalid was interrupted before bready got asserted */
  svt_err_check_stats bvalid_interrupted_check;
  //--------------------------------------------------------------
  /** Checks if rvalid is low when reset is active */
  svt_err_check_stats rvalid_low_when_reset_is_active_check;

  /** Checks if bvalid is low when reset is active */
  svt_err_check_stats bvalid_low_when_reset_is_active_check;

  /** Checks if arvalid is low when reset is active */
  svt_err_check_stats arvalid_low_when_reset_is_active_check;

  /** Checks if acvalid is low when reset is active */
  svt_err_check_stats acvalid_low_when_reset_is_active_check;
  
  /** Checks if crvalid is low when reset is active */
  svt_err_check_stats crvalid_low_when_reset_is_active_check;
  
  /** Checks if cdvalid is low when reset is active */
  svt_err_check_stats cdvalid_low_when_reset_is_active_check;

  /** Checks if awvalid is low when reset is active */
  svt_err_check_stats awvalid_low_when_reset_is_active_check;

  /** Checks if wvalid is low when reset is active */
  svt_err_check_stats wvalid_low_when_reset_is_active_check;
  //--------------------------------------------------------------
  
  /** Checks if write burst cross a 4KB boundary */
  svt_err_check_stats awaddr_4k_boundary_cross_active_check;
  //--------------------------------------------------------------

  /** Checks if write burst of WRAP type has an aligned address*/
  svt_err_check_stats awaddr_wrap_aligned_active_check ;
  //--------------------------------------------------------------
  
  /** Checks if write burst of WRAP type has a valid length*/
  svt_err_check_stats awlen_wrap_active_check;
  //--------------------------------------------------------------

  /** Checks if size of write transfer exceeds the width of the data bus*/
  svt_err_check_stats awsize_data_width_active_check;
  //--------------------------------------------------------------
        
  /** Checks if the value of awburst=2'b11 when awvalid is high*/
  svt_err_check_stats awburst_reserved_val_check;
  //--------------------------------------------------------------
  
  /** Checks if the value of awcache[3:2]=2'b00 when awvalid is high and awcache[1] is also low*/
  svt_err_check_stats awvalid_awcache_active_check;
  //--------------------------------------------------------------

  
  /** Checks if read burst cross a 4KB boundary */
  svt_err_check_stats araddr_4k_boundary_cross_active_check;
  //--------------------------------------------------------------

  /** Checks if read  burst of WRAP type has an aligned address*/
  svt_err_check_stats araddr_wrap_aligned_active_check ;
  //--------------------------------------------------------------

  /** Checks if snoop address is aligned with snoop data width */
  svt_err_check_stats acaddr_aligned_to_cddata_width_valid_check ;
  //--------------------------------------------------------------

  /** Checks that a cached master does not initiate WriteUnique or WriteLineUnique
    * coherent write transaction while any WriteBack, WriteClean or WriteEvict transaction
    * is outstanding.
    */
  svt_err_check_stats complete_outstanding_memory_write_before_writeunique_writelineunique_check ;

  /** Checks that a cached master does not issue WriteBack, WriteClean or WriteEvict
    * transaction while any WriteUnique or WriteLineUnique coherent write transaction
    * is in progress.
    * It automatically checks second rule which says, Complete any incoming snoop 
    * transactions without the use of WriteBack, WriteClean, or WriteEvict
    * transactions while a WriteUnique or WriteLineUnique transaction is in progress.
    */
  svt_err_check_stats complete_outstanding_writeunique_writelineunique_before_memory_write_check ;


  /** Checks that CleanInvalid and MakeInvalid cache maintenance transactions are not 
    * initiated while any memory update or shareable transactions are outstanding. It
    * also checks that CleanShared cache maintenance transactions are not initiated 
    * while any memory update or any shareable transactions that can make the cacheline
    * dirty, are outstanding.
    */
  svt_err_check_stats cache_maintenance_outstanding_transaction_check ;

  /** Checks that WriteBack, WriteClean or any shareable transactions are not issued 
    * while cache maintenance transaction is in progress.
    */
  svt_err_check_stats no_memory_update_or_shareable_txn_during_cache_maintenance_check ;

  /** Monitor checks that when master initiates a CleanShared cache maintenance transaction, 
    * and receives any snoop transaction to the same cacheline, the initiating master must not
    * assert PassDirty snoop response. It also checks that when master initiates CleanInvalid
    * or MakeInvalid cache maintenance transactions, and receives any snoop transaction to the
    * same cacheline, the initiating master must not assert PassDirty, IsShared and DataTransfer
    * snoop responses.
    */
  svt_err_check_stats valid_snoop_response_during_cache_maintenance_check ;
  //--------------------------------------------------------------

  /** Checks if number of databeat transferred over snoop data channel is valid */
  svt_err_check_stats snoop_transaction_burst_length_check ;
  //--------------------------------------------------------------
  
  /** Checks if read burst of WRAP type has a valid length*/
  svt_err_check_stats arlen_wrap_active_check;
  //--------------------------------------------------------------

  /** Checks if size of read transfer exceeds the width of the data bus*/
  svt_err_check_stats arsize_data_width_active_check;
  //--------------------------------------------------------------
        
  /** Checks if the value of arburst=2'b11 when arvalid is high*/
  svt_err_check_stats arburst_reserved_val_check;
  //--------------------------------------------------------------
  
  /** Checks if the value of arcache[3:2]=2'b00 when arvalid is high and arcache[1] is also low*/
  svt_err_check_stats arvalid_arcache_active_check;
  //--------------------------------------------------------------
  
/** Checks if the number of write data items matches AWLEN for the corresponding address */
  svt_err_check_stats wdata_awlen_match_for_corresponding_awaddr_check;
  //--------------------------------------------------------------

/** Checks if the slave must only give a write response after the last write data item is transferred  */
  svt_err_check_stats write_resp_after_last_wdata_check;
  //--------------------------------------------------------------

/** Checks if  A slave must not give a write response before the write address */
  svt_err_check_stats write_resp_after_write_addr_check;
  //--------------------------------------------------------------

/** Checks if the number of read data items matches ARLEN for the corresponding address */
  svt_err_check_stats rdata_arlen_match_for_corresponding_araddr_check;
  //--------------------------------------------------------------

/** Checks if the number of read data items matches ARLEN for the corresponding address */
 svt_err_check_stats rlast_asserted_for_last_read_data_beat;
//ACE CHECKS//

  /** Checks that ACREADY is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acready_when_arvalid_high_check;
  
  /** Checks that ACADDR is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acaddr_when_acvalid_high_check;
  
  /** Checks that ACSNOOP is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acsnoop_when_acvalid_high_check;
  
  /** Checks that ACPROT is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acprot_when_acvalid_high_check;
  
  /** Checks that CDREADY is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cdready_when_cdvalid_high_check;
  
  /** Checks that CDDATA is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cddata_when_cdvalid_high_check;
  
  /** Checks that CDDATACHK is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cddatachk_when_cdvalid_high_check;
  
  /** Checks that CDPOISON is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cdpoison_when_cdvalid_high_check;

 /** Checks that ACREADY is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_cdlast_when_cdvalid_high_check;
  
  /** Checks that CRREADY is not X or Z when CRVALID is high */
  svt_err_check_stats signal_valid_crready_when_crvalid_high_check;
  
  /** Checks that CRRESP is not X or Z when CRVALID is high */
  svt_err_check_stats signal_valid_crresp_when_crvalid_high_check;

  /** Checks that ACADDR is stable when ARVALID is high */
  svt_err_check_stats signal_stable_acaddr_when_acvalid_high_check;
  
  /** Checks that ACSNOOP is stable when ARVALID is high */
  svt_err_check_stats signal_stable_acsnoop_when_acvalid_high_check;
  
  /** Checks that ACPROT is stable when ARVALID is high */
  svt_err_check_stats signal_stable_acprot_when_acvalid_high_check;

  /** Checks that CDDATA is stable when CDVALID is high */
  svt_err_check_stats signal_stable_cddata_when_cdvalid_high_check;
  
  /** Checks that ACREADY is stable when ARVALID is high */
  svt_err_check_stats signal_stable_cdlast_when_cdvalid_high_check;

  /** Checks that CRRESP is stable when CRVALID is high */
  svt_err_check_stats signal_stable_crresp_when_crvalid_high_check;
  
  
/**Checks if the Device transactions, as indicated by AxCACHE[1] = 0, must only use AxDOMAIN = 11.  */
 svt_err_check_stats axcache_axdomain_restriction_check;
  //--------------------------------------------------------------

/**Checks if the  AXCACHE and AXDOMAIN value are valid */
 svt_err_check_stats axcache_axdomain_invalid_value_check ;
  //--------------------------------------------------------------



/**Checks if the  AWSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awsize_valid_value_check;
  //--------------------------------------------------------------
/**Checks if the  ARSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arsize_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWLEN is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awlen_valid_value_check;
  //--------------------------------------------------------------
/**Checks if the  ARLEN is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awsize_valid_check;
  //--------------------------------------------------------------

/**Checks if the  AWBURST is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  ARBURST is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arburst_valid_value_check;
  //--------------------------------------------------------------

 /**Checks if the  ARSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arsize_valid_check;
  //--------------------------------------------------------------

/**Checks if the  address is aligned for AWBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_awburst_wrap_addr_aligned_valid_check;
  //--------------------------------------------------------------
/**Checks if the  address is aligned for ARBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_arburst_wrap_addr_aligned_valid_check;
  //--------------------------------------------------------------
/**Checks if the  address is aligned for AWBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_awburst_incr_addr_aligned_valid_check;
  //--------------------------------------------------------------
/**Checks if the  address is aligned for ARBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_arburst_incr_addr_aligned_valid_check;
  //--------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_awdomain_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  ARDOMAIN is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_ardomain_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_awcache_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  AWLOCK is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_awlock_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  ARLOCK is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_arlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_arcache_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  AxBAR is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_axbar_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  AxLEN is correctly indicated as per the Cache Line Size configured */
 svt_err_check_stats  cache_line_sz_eq_alen_asize_check ;
  //--------------------------------------------------------------

  /**Checks if CLEANSHARED transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats cleanshared_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if CLEANSHAREDPERSIST transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats cleansharedpersist_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if CLEANINVALID transaction starts only from INVALID state */
  svt_err_check_stats cleaninvalid_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if MAKEINVALID transaction starts only from INVALID state */
  svt_err_check_stats makeinvalid_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if WRITEUNIQUE transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats writeunique_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if WRITELINEUNIQUE transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats writelineunique_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if WRITEBACK transaction starts only from UNIQUEDIRTY or SHAREDDIRTY state */
  svt_err_check_stats writeback_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if WRITECLEAN transaction starts only from UNIQUEDIRTY or SHAREDDIRTY state */
  svt_err_check_stats writeclean_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if WRITEEVICT transaction starts only from UNIQUECLEAN state */
  svt_err_check_stats writeevict_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if EVICT transaction starts only from UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats evict_correct_start_state_check;         
  //--------------------------------------------------------------

  /**Checks if snoop response has data transfer bit set for cacheline in dirty state */
  svt_err_check_stats dirty_state_data_transfer_check;         
  //--------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for ReadOnce & WriteUnique Transactions */
 svt_err_check_stats  writeunique_awdomain_valid_value_check;
//------------------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for WriteUniquePtlstash Transactions */
 svt_err_check_stats  writeuniqueptlstash_awdomain_valid_value_check;

  //--------------------------------------------------------------
/**Checks if the  AWDOMAIN is valid for ReadOnce & WriteUnique Transactions */
 svt_err_check_stats  readonce_ardomain_valid_value_check;
  //--------------------------------------------------------------

 /**Checks if all transactions (other than ReadNoSnoop, ReadOnce, ReadOnceCleanInvalid, ReadOnceMakeInvalid, WriteNoSnoop, WriteUnique) are required to be a full cache line size */
 svt_err_check_stats  full_cache_line_size_check;

/**Checks if the  AWBURST is valid for ReadOnce & WriteUnique Transactions */
 svt_err_check_stats writeunique_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWBURST is valid for writeuniqueptlstash Transactions */
 svt_err_check_stats writeuniqueptlstash_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  ARBURST is valid for ReadOnce & WriteUnique  Transactions */
 svt_err_check_stats readonce_arburst_valid_value_check;


/**Checks if the  AWCACHE is valid for ReadOnce & WriteUnique  Transactions */
 svt_err_check_stats  writeunique_awcache_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWLOCK is valid for ReadOnce & WriteUnique  Transactions */
 svt_err_check_stats  writeunique_awlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for writeuniqueptlstash  Transactions */
 svt_err_check_stats  writeuniqueptlstash_awcache_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWLOCK is valid for writeuniqueptlstash  Transactions */
 svt_err_check_stats  writeuniqueptlstash_awlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  ARCACHE is valid for ReadOnce & WriteUnique   Transactions */
 svt_err_check_stats  readonce_arcache_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  ARLOCK is valid for ReadOnce & WriteUnique   Transactions */
 svt_err_check_stats  readonce_arlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWSIZE is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awsize_valid_value_check;
  //--------------------------------------------------------------


/**Checks if the  AWSIZE is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWLEN for INCR is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_awlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWLEN for INCR is valid for AXI Transactions */
 svt_err_check_stats awburst_awlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWBURST is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awdomain_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awcache_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  Address aligned for WRAP is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_incr_valid_check;
  //--------------------------------------------------------------

/**Checks if the AWSIZE x AWLEN  not exceed the cache line size  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_wrap_valid_check;
//--------------------------------------------------------------

/**Checks if the ALOCK is 0 for WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awlock_valid_value_check;
//--------------------------------------------------------------
/** If a snooped master receives a snoop transaction when it is has an
 * outstanding WriteEvict transaction, then it is the responsibility of the
 * snooped master to ensure that no other master can update the same area of
 * main memory at the same time. The snooped master achieves this by delaying
 * the snoop response until the snooped master has completed the WriteEvict
 * transaction */
 svt_err_check_stats snoop_response_to_same_cacheline_during_writeevict_check;
//--------------------------------------------------------------
/** While a transaction is in progress which has the AWUNIQUE signal asserted,
 * the master must not give a snoop response that would allow another copy of
 * the line to be created, or an agent to consider that it has another Unique
 * copy of the line
 */
 svt_err_check_stats snoop_response_to_same_cacheline_during_xact_with_awunique_check;
//--------------------------------------------------------------
/** AWUNIQUE must be deasserted for WRITECLEAN transactions */
svt_err_check_stats writeclean_awunique_valid_value_check;
//--------------------------------------------------------------
/** AWUNIQUE must be asserted for WRITEEVICT transactions */
svt_err_check_stats writeevict_awunique_valid_value_check;
//--------------------------------------------------------------
/** Monitor check that all byte strobes are asserted for a WRITEEVICT transaction */
svt_err_check_stats writeevict_wstrb_valid_value_check;

//--------------------------------------------------------------
/** Monitor check that all byte strobes are asserted for a WRITELINEUNIQUE transaction */
svt_err_check_stats writelineunique_wstrb_valid_value_check;
//--------------------------------------------------------------

/** Monitor check that all byte strobes are asserted for a writeuniquefullstash transaction */
svt_err_check_stats writeuniquefullstash_wstrb_valid_value_check;
//--------------------------------------------------------------

//--------------------------------------------------------------
/**Checks the valid response of EXOKAY response is only for readnosnoop Transactions */
svt_err_check_stats exokay_resp_observed_only_for_exclusive_transactions_check;
//--------------------------------------------------------------
/**Checks that if cacheline is in invalid state then exclusive load transaction is issued only as READCLEAN or READSHARED */
svt_err_check_stats exclusive_load_from_valid_state_check;
//--------------------------------------------------------------
/**Checks that if cacheline is in invalid state then exclusive store transaction is not issued */
svt_err_check_stats exclusive_store_from_valid_state_check;
//--------------------------------------------------------------
/**Checks that if cacheline is in shared state then exclusive transaction is issued only as CLEANUNIQUE, READCLEAN or READSHARED*/
svt_err_check_stats exclusive_transaction_from_shared_state_check;
//--------------------------------------------------------------
/**Checks for no data transfer occurs for a CleanShared,Cleansharedpersist, CleanInvalid, CleanUnique, MakeUnique, MakeInvalid and Evict Transactions */
svt_err_check_stats perform_no_datatransfer_check;
  //--------------------------------------------------------------
/**Checks the valid response of  cleanshared Transactions */
svt_err_check_stats read_data_chan_cleanshared_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  cleansharedPersist Transactions */
svt_err_check_stats read_data_chan_cleansharedpersist_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of makeinvalid  Transactions */
svt_err_check_stats read_data_chan_makeinvalid_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  makeunique Transactions */
svt_err_check_stats read_data_chan_makeunique_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of cleaninvalid  Transactions */
svt_err_check_stats read_data_chan_cleaninvalid_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  cleanunique Transactions */
svt_err_check_stats read_data_chan_cleanunique_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  readunique Transactions */
svt_err_check_stats read_data_chan_readunique_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  readnotshareddirty Transactions */
svt_err_check_stats read_data_chan_readnotshareddirty_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  readclean Transactions */
svt_err_check_stats read_data_chan_readclean_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of readonce  Transactions */
svt_err_check_stats read_data_chan_readonce_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of readnosnoop  Transactions */
svt_err_check_stats read_data_chan_readnosnoop_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the CLEANUNIQUE, MAKEUNIQUE, CLEANSHARED,
  * CLEANINVALID,CLEANSHAREDPERSIST,
  * MAKEINVALID, READBARRIER, DVMCOMPLETE, DVMMESSAGE transactions
  * have only single read data channel transfer */
svt_err_check_stats coherent_single_read_data_transfer_valid_check;
  //--------------------------------------------------------------

/**Checks the valid response of readbarrier  Transactions */
svt_err_check_stats read_data_chan_readbarrier_resp_valid_check;
  //--------------------------------------------------------------

/**Checks the valid response of DVM Message Transactions */
svt_err_check_stats read_data_chan_dvmmessage_resp_valid_check;
  //--------------------------------------------------------------

/**Checks the valid response of DVM Complete Transactions */
svt_err_check_stats read_data_chan_dvmcomplete_resp_valid_check;

//--------------------------------------------------------------
/**Checks the valid snoop response of DVM Message Transactions */
svt_err_check_stats snoop_chan_dvmsync_resp_valid_check;
  //--------------------------------------------------------------

/**Checks the valid snoop response of DVM Complete Transactions */
svt_err_check_stats snoop_chan_dvmcomplete_resp_valid_check;

//--------------------------------------------------------------
/**Checks the ACSNOOP reserved values */
svt_err_check_stats acsnoop_reserved_value_check ;
 //--------------------------------------------------------------


/**Checks that for MakeInvalid transactions a data transfer is never required */
svt_err_check_stats snoop_resp_passdirty_datatransfer_check;
//--------------------------------------------------------------

/**If DataTransfer is asserted, a full cache line of data must be provided on the snoop data channel */
svt_err_check_stats full_cache_line_datatransfer_check;
//

/**Checks for readunique cleaninvalid makeinvalid illegal response  */
svt_err_check_stats snoop_response_channel_isshared_check;
//--------------------------------------------------------------

/** Checks that CDLAST signal is asserted during the final data transfer.
  *
  * protocol checks : port level 
  */
svt_err_check_stats cdlast_asserted_for_last_snoopread_data_beat;
//--------------------------------------------------------------

/**Checks that the FIXED burst type is not supported for shareable transactions */
svt_err_check_stats fixed_burst_type_valid;
//--------------------------------------------------------------

/**Checks that ACVALID and ACREADY to be asserted before asserting CRVALID */
svt_err_check_stats snoop_addr_snoop_resp_check;
//--------------------------------------------------------------
/**Checks that ACVALID and ACREADY to be asserted before asserting CDVALID */
svt_err_check_stats snoop_addr_snoop_data_check;
//--------------------------------------------------------------

//--------------------------------------------------------------
/**Checks the combinations of ARDOMAIN,ARSNOOP and ARBAR are valid and unreserved */
svt_err_check_stats arsnoop_ardomain_arbar_reserve_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWDOMAIN,AWSNOOP and AWBAR are valid and unreserved */
svt_err_check_stats awsnoop_awdomain_awbar_reserve_value_check;
//--------------------------------------------------------------

//Barrier Checks //
/**Checks the AWADDR is valid for AWBAR  */
svt_err_check_stats write_barrier_awaddr_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations AWBURST and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awburst_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWLEN and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awlen_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWSIZE and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awsize_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWCACHE and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awcache_type_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWSNOOP and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awsnoop_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWLOCK and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awlock_type_valid_value_check;
//--------------------------------------------------------------
/**Checks the valid value of AxUSER for write barrier transactions */
svt_err_check_stats barrier_transaction_user_valid_value_check;
//--------------------------------------------------------------

/**Checks the ARADDR is valid for ARBAR  */
svt_err_check_stats read_barrier_araddr_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations ARBURST and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arburst_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARLEN and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arlen_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARSIZE and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arsize_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARCACHE and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arcache_type_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARSNOOP and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arsnoop_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARLOCK and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arlock_type_valid_value_check;
//--------------------------------------------------------------
/** Checks the Barrier Id valid and unreserved.  */
svt_err_check_stats barrier_id_valid_value_check;
//--------------------------------------------------------------
/**Checks the Read Barrier valid response  */
svt_err_check_stats barrier_read_response_check ;
//--------------------------------------------------------------
/**Checks the Write Barrier valid response  */
svt_err_check_stats barrier_write_response_check ;
//--------------------------------------------------------------
/**Checks that both transactions in a barrier pair must have the same AxID, AxBAR, AxDOMAIN, and AxPROT values*/
svt_err_check_stats barrier_pair_cntrl_signals_check ;
//--------------------------------------------------------------
/**Checks that barrier pairs must be issued in the same sequence on the read address and write address channels*/
svt_err_check_stats barrier_pair_check ;
//--------------------------------------------------------------
/**Checks that ARADDR/AWADDR should always be aligned to Atomicity Size*/
svt_err_check_stats align_addr_atomicity_size_check ;

//--------------------------------------------------------------
/** Checks the RACK for valid response.  */
svt_err_check_stats rack_status_check;
//--------------------------------------------------------------
/** Checks the WACK for valid response.  */
svt_err_check_stats wack_status_check;
//-------------------------------------------------------------
/** Checks all snoop transactions are ordered. .
  */
svt_err_check_stats snoop_transaction_order_check;

//DVM CHECKS //
 /**Checks  For DVM ARBURST 'b01 Burst Type INCR. */
svt_err_check_stats dvm_message_arburst_valid_value_check;
//-------------------------------------------------------------
 /**Checks For DVM  ARLEN All zero */
svt_err_check_stats dvm_message_arlen_valid_value_check;
//-------------------------------------------------------------

 /**Checks for DVM ARSIZE Matches the data bus width */
svt_err_check_stats dvm_message_arsize_valid_value_check;
//-------------------------------------------------------------

 /**Checks for DVM ARCACHE 'b0010 Normal non-cacheable */
svt_err_check_stats dvm_message_arcache_type_valid_value_check;
//-------------------------------------------------------------

 /**Checks for DVM ARLOCK 'b0 Normal Access. */
svt_err_check_stats dvm_message_arlock_type_valid_value_check;
//-------------------------------------------------------------
 
/**Checks for DVM  ARDOMAIN  is Inner shareable or Outer shareable */ 
svt_err_check_stats dvm_message_ardomain_type_valid_value_check;
//-------------------------------------------------------------
/**Checks for DVM  ARBAR[0] is 1'b0 */ 
svt_err_check_stats dvm_message_arbar_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMCOMPLETE the valid value of  ARSNOOP */ 
svt_err_check_stats dvm_complete_arsnoop_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMSYNC, DVM Operation the valid value of  ARSNOOP */ 
svt_err_check_stats dvm_operation_dvm_sync_arsnoop_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMSYNC, DVM Operation the valid value of ARADDR[(n-1):32],[15],[11:0] bits */
svt_err_check_stats dvm_operation_dvm_sync_araddr_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMHINT, DVM Operation the valid value of ARADDR[15] */
svt_err_check_stats dvm_operation_dvm_hint_araddr_valid_value_check;
//-------------------------------------------------------------

/** Checks the value of  ACSNOOP for the DVM complete */ 
svt_err_check_stats dvm_complete_acsnoop_valid_value_check;
//-------------------------------------------------------------
/** Checks the value of  ACSNOOP for the DVM SYNC */ 
svt_err_check_stats dvm_operation_dvm_sync_acsnoop_valid_value_check;
//-------------------------------------------------------------

/** Checks For a DVM Complete message, ARADDR is defined to be all zeros */
svt_err_check_stats dvmcomplete_araddr_valid_value_check;
//-------------------------------------------------------------
/** Checks  For a DVM Complete message, ACADDR is defined to be all zeros */
svt_err_check_stats dvmcomplete_acaddr_valid_value_check;
//-------------------------------------------------------------


/** Checks  FOR DVM Message the value of reserve address bit should be zero  */
svt_err_check_stats dvmmessage_araddr_reserve_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[11:10] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_hypervisor_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[9:8] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[6] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[5] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type Branch Predictor Invalidate */
svt_err_check_stats dvmmessage_branch_predictor_invalidate_supported_message_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[9:8] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_secure_nonsecure_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[6:5] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_vid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[11:10] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_invalidate_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[9:8] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[6] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[5] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_addr_specified_value_check;
//-------------------------------------------------------------


//DVM snoop

/** Checks  FOR DVM Message the value of reserve address bit should be zero  */
svt_err_check_stats dvmmessage_snoop_araddr_reserve_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[11:10] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_hypervisor_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[9:8] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[6] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[5] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_snoop_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type Branch Predictor Invalidate */
svt_err_check_stats snoop_dvmmessage_branch_predictor_invalidate_supported_message_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[9:8] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_physical_inst_cache_secure_nonsecure_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[6:5] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_physical_inst_cache_vid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_snoop_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[11:10] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_invalidate_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[9:8] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[6] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[5] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_snoop_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks the overlapping AWID of Write Barrier transactions with any active Write transactions */
svt_err_check_stats writebarrier_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the overlapping ARID of Read Barrier transactions with any active Read transactions */
svt_err_check_stats readbarrier_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the overlapping ARID of DVM transactions with any active Read transactions */
svt_err_check_stats dvm_xact_id_overlap_check;

/** Checks the overlapping ARID of Non-DVM or Non-Device transactions with any active transactions */
svt_err_check_stats read_non_dvm_non_device_xact_id_overlap_check;

/** Checks the overlapping AWID of Non-DVM or Non-Device transactions with any active transactions*/
svt_err_check_stats write_non_dvm_non_device_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks that all transactions of multi-part DVM operation have same ID */
svt_err_check_stats multipart_dvm_coherent_same_id_check;
//-------------------------------------------------------------
/** Checks that all transactions of multi-part DVM operation have same coherent response */
svt_err_check_stats multipart_dvm_coherent_same_response_check;
//-------------------------------------------------------------
/** Checks that all coherent transactions of multi-part DVM operation are sent in successive manner 
    and no unrelated coherent transaction sent during multi-part DVM opearion over AR channel */
svt_err_check_stats multipart_dvm_coherent_successive_transaction_check;
//-------------------------------------------------------------
/** Checks that all transactions of multi-part DVM operation have same snoop response */
svt_err_check_stats multipart_dvm_snoop_same_response_check;
//-------------------------------------------------------------
/** Checks that all snoop transactions of multi-part DVM operation are sent in successive manner 
    and no unrelated snoop transaction sent during multi-part DVM opearion over AC channel */
svt_err_check_stats multipart_dvm_snoop_successive_transaction_check;
//-------------------------------------------------------------
/** Checks the overlapping ARID of Non-Barrier Non-DVM transactions with any active Barrier/DVM transactions */
svt_err_check_stats readbarrier_dvm_norm_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the overlapping AWID of Non-Barrier Non-DVM transactions with any active Barrier/DVM transactions */
svt_err_check_stats writebarrier_norm_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the receiverd RDATACHK is same as the parity calculated from RDATA in a read  transaction */
svt_err_check_stats rdatachk_parity_calculated_rdata_parity_check;
//-------------------------------------------------------------
/** Checks the receiverd parity is same as the parity calculated from respective signal in a transaction */
svt_err_check_stats received_parity_calculated_parity_check;
//-------------------------------------------------------------
/** Checks the receiverd WDATACHK is same as the parity calculated from WDATA in a write transaction */
svt_err_check_stats wdatachk_parity_calculated_wdata_parity_check;
//-------------------------------------------------------------
/** Checks the receiverd CDDATACHK is same as the parity calculated from CDDATA in a snoop transaction */
svt_err_check_stats cddatachk_parity_calculated_cddata_parity_check;
//-------------------------------------------------------------

// Checks on 'Sequencing Transactions'

/** Checks that Master does not receive a snoop transaction until 
  * any preceding transaction to the same cache line has completed
  */
svt_err_check_stats resp_to_same_cache_line_check;
//-------------------------------------------------------------
/** Checks that if received a snoop transaction, response to a transaction 
  * to the same cache line is not received , until snoop response is sent 
  */
svt_err_check_stats snoop_to_same_cache_line_check;
//-------------------------------------------------------------
/**
  * Checks that the if DataTransfer de-asserted then no data transfer will occur on the snoop data channel
  *  for this transaction DataTransfer, CRRESP[0]
  */
svt_err_check_stats cdvalid_high_no_data_transfer_check;
//-------------------------------------------------------------
// START OF LOCKED ACCESS CHECKS
/**
  * Checks that there are no pending transactions before a locked
  * sequence starts
  */
svt_err_check_stats no_pending_xacts_during_locked_xact_sequeunce_check;
//-------------------------------------------------------------

/**
  * Checks that all transactions of locked sequence have the same id
  */
svt_err_check_stats locked_sequeunce_id_check;
//-------------------------------------------------------------

/**
  * Checks that when a master does a lock transaction, it does not target subsequent transactions in the lock 
  * sequence to any slave other than the locked slave
  */

svt_err_check_stats locked_sequence_to_same_slave_check;
 //----------------------------------------------------------------
/**
  * Check that the master follows as per the recommendation from spec to  limit 2 transaction for the lock access
  */
   svt_err_check_stats locked_sequence_length_check;
//-------------------------------------------------------------

/**
  * Checks that there are no pending transactions of a locked sequeunce
  * when a normal transaction is received
  */
svt_err_check_stats no_pending_locked_xacts_before_normal_xacts_check;
// END OF LOCKED ACCESS CHECKS

/** 
  * Checks that AXI master and AXI slave are not exceeding the user 
  * configured maximum number of outstanding transactions (#num_outstanding_xact)
  * If #num_outstanding_xact = -1 then #num_outstanding_xact will not be considered , 
  * instead #num_read_outstanding_xact and #num_write_outstanding_xact will be considered for 
  * read and write transactions respectively.
  */
svt_err_check_stats max_num_outstanding_xacts_check ;

//-------------------------------------------------------------
// START OF PERFORMANCE CHECKS
/**
  * Checks that the latency of a write transaction is not greater than the
  * configured max value
  */
svt_err_check_stats perf_max_write_xact_latency_check;

/**
  * Checks that the latency of a write transaction is not lesser than the
  * configured min value
  */
svt_err_check_stats perf_min_write_xact_latency_check;

/**
  * Checks that the average latency of write transactions in a given interval
  * is not more than the configured max value
  */
svt_err_check_stats perf_avg_max_write_xact_latency_check;

/**
  * Checks that the average latency of write transactions in a given interval
  * is not less than the configured min value
  */
svt_err_check_stats perf_avg_min_write_xact_latency_check;

/**
  * Checks that the latency of a read transaction is not greater than the
  * configured max value
  */
svt_err_check_stats perf_max_read_xact_latency_check;

/**
  * Checks that the latency of a read transaction is not lesser than the
  * configured min value
  */
svt_err_check_stats perf_min_read_xact_latency_check;

/**
  * Checks that the average latency of read transactions in a given interval
  * is not more than the configured max value
  */
svt_err_check_stats perf_avg_max_read_xact_latency_check;

/**
  * Checks that the average latency of read transactions in a given interval
  * is not less than the configured min value
  */
svt_err_check_stats perf_avg_min_read_xact_latency_check;

/**
  * Checks that the throughput of read transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_read_throughput_check;

/**
  * Checks that the throughput of read transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_read_throughput_check;

/**
  * Checks that the throughput of write transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_write_throughput_check;

/**
  * Checks that the throughput of write transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_write_throughput_check;

/**
  * Checks that the bandwidth of read transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_read_bandwidth_check;

/**
  * Checks that the bandwidth of read transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_read_bandwidth_check;

/**
  * Checks that the bandwidth of write transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_write_bandwidth_check;

/**
  * Checks that the bandwidth of write transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_write_bandwidth_check;

// END OF PERFORMANCE CHECKS
//-------------------------------------------------------------
// START Of STREAM CHECKS

svt_err_check_stats signal_valid_tvalid_check;

/** Checks that TREADY is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tready_when_tvalid_high_check;

/** If tdata is enabled, checks that TDATA is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tdata_when_tvalid_high_check;

/** If tstrb is enabled, checks that TSTRB is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tstrb_when_tvalid_high_check;

/** If tkeep is enabled, checks that TKEEP is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tkeep_when_tvalid_high_check;

/** If tlast is enabled, checks that TLAST is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tlast_when_tvalid_high_check;

/** If tid is enabled, checks that TID is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tid_when_tvalid_high_check;

/** If tuser is enabled, checks that TUSER is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tuser_when_tvalid_high_check;

/** If tdest is enabled, checks that TDEST is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tdest_when_tvalid_high_check;

/** 
  * Checks that TDATA is stable when TVALID is high 
  * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=1 ,
  * it considers only valid byte lanes of tdata based on tstrb. 
  * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=0 ,
  * whole tdata as seen on the bus will be considered.
  */
svt_err_check_stats signal_stable_tdata_when_tvalid_high_check;

/** Checks that TSTRB is stable when TVALID is high */
svt_err_check_stats signal_stable_tstrb_when_tvalid_high_check;

/** Checks that TKEEP is stable when TVALID is high */
svt_err_check_stats signal_stable_tkeep_when_tvalid_high_check;

/** Checks that TLAST is stable when TVALID is high */
svt_err_check_stats signal_stable_tlast_when_tvalid_high_check;

/** Checks that TID is stable when TVALID is high */
svt_err_check_stats signal_stable_tid_when_tvalid_high_check;

/** Checks that TUSER is stable when TVALID is high */
svt_err_check_stats signal_stable_tuser_when_tvalid_high_check;

/** Checks that TDEST is stable when TVALID is high */
svt_err_check_stats signal_stable_tdest_when_tvalid_high_check;

/** Checks that TVALID is low when reset is active */
svt_err_check_stats tvalid_low_when_reset_is_active_check;

/** Checks if tvalid was interrupted before tready got asserted */
svt_err_check_stats tvalid_interrupted_check;

/** Checks that TSTRB is low if TKEEP is low */
svt_err_check_stats tstrb_low_when_tkeep_low_check;

/** Checks that received data stream is not interleaved beyond stream_interleave_depth
  * value. An error is issued if data stream is interleaved beyond this value. */
svt_err_check_stats stream_interleave_depth_check;

/** Checks that the burst length of received data stream is not exceeding the maximum
  * value allowed for stream_burst_length defined by `SVT_AXI_MAX_STREAM_BURST_LENGTH. */
svt_err_check_stats max_stream_burst_length_exceeded_check;

/** 
 * @groupname port_interleaving_check
 * @check_description   
 * - Checks if address does fall to correct interleaved port.
 * - Valid when port cfg port_interleaving_enable = 1.   
 * .
 * @end_check_description
 *
 * @check_pass
 * address does fall to correct interleaved port. 
 * @end_check_pass
 *
 * @check_fail
 * address does not fall to correct interleaved port. 
 * @end_check_fail
 *
 * @applicable_device_type
 * master & slave 
 * @end_applicable_device_type
 *
 * @check_additional_information
 * @end_check_additional_information   
 */
svt_err_check_stats port_interleaving_check;

/** 
 * @groupname trace_tag_validity_check
 * @check_description   
 * - Trace tag value on data channel or resposne channel should be valid as per the trace tag 
 * - value on the address channel. 
 * .
 * @end_check_description
 *
 * @check_pass
 * For Write transactions the check will pass if:
 * A slave that receives a write request with AWTRACE asserted should assert the BTRACE signal alongside
 * the write response.
 * For Read transactions the check will pass if:
 * A slave that receives a read request with the ARTRACE signal asserted should assert the RTRACE signal
 * alongside every beat of the read response.
 * For Snoop transactions the check will pass if:
 * A master that receives a snoop request with the ACTRACE signal asserted should assert the CRTRACE
 * signal alongside the snoop response.The master should also assert CDTRACE alongside every data beat of
 * the snoop data that is associated with the snoop transaction.
 * @end_check_pass
 * @check_fail
 * If trace_tag in the request packet is set to 1 and in the spawned response or data packet is set 
 * to 0.
 * @end_check_fail
 *
 * @applicable_device_type
 * @end_applicable_device_type
 *
 * @check_additional_information
 * @end_check_additional_information   
 */
svt_err_check_stats trace_tag_validity_check;


// END OF STREAM CHECKS
//-------------------------------------------------------------
  `ifdef SVT_AXI_QVN_ENABLE
// START OF QVN CHECKS    

/** Checks that VARVALIDVN* is not X or Z */
svt_err_check_stats signal_valid_varvalidvnx_check;

/** Checks the VARQOSVN* is valid when VARVALIDVN* is high */
svt_err_check_stats  signal_valid_varqosvnx_when_varvalidvnx_high_check;  
   
/** Checks that VARREADYVN* is not X or Z */
svt_err_check_stats signal_valid_varreadyvnx_check;

/** Checks that VAWVALIDVN* is not X or Z */
svt_err_check_stats signal_valid_vawvalidvnx_check;

/** Checks the VAWQOSVN* is valid when VAWVALIDVN* is high */
svt_err_check_stats  signal_valid_vawqosvnx_when_vawvalidvnx_high_check;  
   
/** Checks that VAWREADYVN* is not X or Z */
svt_err_check_stats signal_valid_vawreadyvnx_check;
   
/** Checks that VWVALIDVN* is not X or Z */
svt_err_check_stats signal_valid_vwvalidvnx_check;

/** Checks that VWREADYVN* is not X or Z */
svt_err_check_stats signal_valid_vwreadyvnx_check;
   
/** Checks that VARVALIDVN* when asserted, remains asserted till VARREADYVN* */   
svt_err_check_stats varvalidvn_deassertion_check;
   
/** When a master sets VARVALIDVNx high, it can change VARQOSVNx proir to the slave granting a token, but only if the value increase. */
svt_err_check_stats varqosvn_valid_change_check;

/** Checks that VAWVALIDVN* when asserted, remains asserted till VAWREADYVN* */   
svt_err_check_stats vawvalidvn_deassertion_check;
   
/** When a master sets VAWVALIDVNx high, it can change VAWQOSVNx proir to the slave granting a token, but only if the value increase. */
svt_err_check_stats vawqosvn_valid_change_check;
   
/** Checks that VWVALIDVN* when asserted, remains asserted till VWREADYVN* */   
svt_err_check_stats vwvalidvn_deassertion_check;

/** Check that master must only set ARVNET to values that correspond to a VN where the associated set of token request signals exist.*/
svt_err_check_stats arvnet_for_existing_vn_check;
   
/** Check that master must only set AWVNET to values that correspond to a VN where the associated set of token request signals exist.*/
svt_err_check_stats awvnet_for_existing_vn_check;

/** Check that master must only set WVNET to values that correspond to a VN where the associated set of token request signals exist.*/
svt_err_check_stats wvnet_for_existing_vn_check;

/** Check that master must have read address token for VN denote ARVNET, before it can send read address channel transfer (Except for a Barrier transaction).*/
svt_err_check_stats rd_addr_chan_vn_token_availability_check;
   
/** Check that master must have write address token for VN denote AWVNET, before it can send write address channel transfer (Except for a Barrier transaction).*/
svt_err_check_stats wr_addr_chan_vn_token_availability_check;
   
/** Check that master must have write data token for VN denote WVNET, before it can send a data beat. */
svt_err_check_stats wr_data_chan_vn_token_availability_check;

/** Check that transaction with the same AXI ID that are are sent on the same physical link must use the same VN.*/
svt_err_check_stats same_axi_id_over_single_vn_check;

/** Check Before entering a low-power or reset state, the component must have the same number of pre-allocated tokens that it had when it exited reset.*/
svt_err_check_stats pre_allocated_token_count_at_rst_check;

/** Check QVN token handshake signal are not asserted on unsupported VN.*/
svt_err_check_stats qvn_sig_asrt_on_unsupported_vn_check;

/** Check that slave component is not granting more outstanding token than its configured.*/
svt_err_check_stats slave_max_outstanding_token_check;
   
/** Check that token requested should be granted in a bounded time*/
svt_err_check_stats qvn_token_request_timeout_check;
   
//-------------------------------------------------------------
// END OF QVN CHECKS    
`endif

`ifdef SVT_ACE5_ENABLE

//--------------------------------------------------------------
/** Checks that ARCHUNKEN is not X or Z when ARVALID is high */
svt_err_check_stats signal_valid_archunken_when_arvalid_high_check;

//--------------------------------------------------------------
/** Checks that RCHUNKV is not X or Z when RVALID is high */
svt_err_check_stats signal_valid_rchunkv_when_rvalid_high_check;
  
/** Checks that RCHUNKNUM is not X or Z when RVALID and RCHUNKV are high */
svt_err_check_stats signal_valid_rchunknum_when_rvalid_rchunkv_high_check;

/** Checks that RCHUNKSTRB is not X or Z when RVALID and RCHUNKV are high */
svt_err_check_stats signal_valid_rchunkstrb_when_rvalid_rchunkv_high_check;


//--------------------------------------------------------------
/** Checks that ARCHUNKEN is stable when ARVALID is high */
svt_err_check_stats signal_stable_archunken_when_arvalid_high_check;

//--------------------------------------------------------------
/** Checks that RCHUNKV is stable when RVALID is high */
svt_err_check_stats signal_stable_rchunkv_when_rvalid_high_check;

/** Checks that RCHUNKNUM is stable when RVALID and RCHUNKV are high */
svt_err_check_stats signal_stable_rchunknum_when_rvalid_rchunkv_high_check;

/** Checks that RCHUNKSTRB is stable when RVALID and RCHUNKV are high */
svt_err_check_stats signal_stable_rchunkstrb_when_rvalid_rchunkv_high_check;


//--------------------------------------------------------------
/** Checks that ARSIZE is equal to the data bus width or ARLEN is one beat and
 * ARSIZE is 128 bits or larger for rdata chunking */
svt_err_check_stats rdata_chunking_arsize_valid_value_check;

/** Checks that ARADDR is aligned to 16 bytes for rdata chunking */
svt_err_check_stats rdata_chunking_araddr_aligned_check; 

/** Checks that ARBURST is INCR or WRAP for rdata chunking */
svt_err_check_stats rdata_chunking_arburst_type_check;

/**Checks that ARSNOOP is ReadNoSnoop, ReadOnce, ReadOnceCleanInvalid or 
 * ReadOnceMakeInvalid for rdata chunking */
svt_err_check_stats rdata_chunking_arsnoop_valid_value_check;

/** Checks that ARIDUNQ must be asserted for rdata chunking */
svt_err_check_stats rdata_chunking_aridunq_valid_value_check;

//--------------------------------------------------------------  
/**Checks that RCHUNKV is deasserted for all the transfers when ARCHUNKEN is
 * deasserted */
svt_err_check_stats rdata_chunking_rchunkv_zero_when_archunken_deasserted_check;

/**Checks that RCHUNKV must be the same for every response beat of a 
 * transaction */ 
svt_err_check_stats rdata_chunking_rchunkv_same_for_all_response_check;

/** Checks that RCHUNKNUM must be between zero and ARLEN when RVALID and
 * RCHUNKV are high*/
svt_err_check_stats rdata_chunking_rchunknum_valid_value_check;

/**Checks that RCHUNKSTRB must not be zero when RVALID and RCHUNKV are high */
svt_err_check_stats rdata_chunking_rchunkstrb_valid_value_check;

/**Checks that the number of bytes that are transferred through read data
 * chunking must be consistant with ARSIZE and ARLEN */
svt_err_check_stats rdata_chunking_num_bytes_transfer_check;

`endif

`ifdef SVT_UVM_TECHNOLOGY
  /** UVM report server passed in through the constructor */
  uvm_report_object reporter;
`elsif SVT_OVM_TECHNOLOGY
  /** OVM report server passed in through the constructor */
  ovm_report_object reporter;
`else
  /** VMM message service passed in through the constructor*/ 
  vmm_log  log;
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_port_configuration cfg, uvm_report_object reporter, bit register_enable=1, bit enable_pc_cov = 1);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_port_configuration cfg, ovm_report_object reporter, bit register_enable=1, bit enable_pc_cov = 1);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param log VMM log instance used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (string name, svt_axi_port_configuration cfg, vmm_log log = null, bit register_enable=1, bit enable_pc_cov = 1);
`endif
  /** @cond PRIVATE */
  extern function void perform_excl_write_addr_chan_signal_level_checks(svt_axi_transaction xact, 
                       svt_axi_transaction excl_xact, output bit is_excl_wr_error);
 
  extern function void perform_read_addr_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_arid,
                                                       ref logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] observed_araddr,
                                                       ref logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] observed_arlen,
                                                       ref logic[`SVT_AXI_SIZE_WIDTH-1:0] observed_arsize,
                                                       ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_arburst,
                                                       ref logic[`SVT_AXI_LOCK_WIDTH-1:0] observed_arlock,
                                                       ref logic[`SVT_AXI_CACHE_WIDTH-1:0] observed_arcache,
                                                       ref logic[`SVT_AXI_PROT_WIDTH-1:0] observed_arprot,
                                                       ref logic[`SVT_AXI_QOS_WIDTH-1:0] observed_arqos,
                                                       ref logic[`SVT_AXI_REGION_WIDTH-1:0] observed_arregion,
                                                       ref logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] observed_aruser,
                                                       ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain,
                                                       ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                                       ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
                                                       ref logic observed_arready,
`ifdef SVT_ACE5_ENABLE
                                                       ref logic[`SVT_AXI_MAX_MMUSID_WIDTH-1:0]observed_stream_id,
                                                       ref logic[`SVT_AXI_MAX_MMUSSID_WIDTH-1:0]observed_sub_stream_id,
                                                       ref logic observed_secure_or_non_secure_stream,
                                                       ref logic observed_sub_stream_id_valid,
                                                       ref logic observed_addr_translated_from_pcie,
                                                       ref logic observed_aridunq, 
                                                       ref logic observed_archunken,
                                                       ref logic [`SVT_AXI_MAX_MPAM_WIDTH-1:0] observed_armpam,
                                                       output bit is_aridunq_valid, 
                                                       output bit is_archunken_valid,
                                                       output bit is_stream_id_valid,                              
                                                       output bit is_sub_stream_id_valid,                          
                                                       output bit is_secure_or_non_secure_stream_valid,                              
                                                       output bit is_sub_streamid_valid,                          
                                                       output bit is_addr_translated_from_pcie_valid,
                                                       output bit is_armpam_valid,     
 `endif
                                                       output bit is_arid_valid,
                                                       output bit is_araddr_valid,
                                                       output bit is_arlen_valid,
                                                       output bit is_arsize_valid,
                                                       output bit is_arburst_valid,
                                                       output bit is_arlock_valid,
                                                       output bit is_arcache_valid,
                                                       output bit is_arprot_valid,
                                                       output bit is_arqos_valid,
                                                       output bit is_arregion_valid,
                                                       output bit is_aruser_valid,
                                                       output bit is_ardomain_valid,
                                                       output bit is_arsnoop_valid,
                                                       output bit is_arbar_valid,
                                                       output bit is_arready_valid,
                                                       output bit excl_read_error
                                                     );
  extern function void perform_read_data_chan_signal_level_checks(
                                                      ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_rid,
                                                      ref logic[`SVT_AXI_RESP_WIDTH-1:0] observed_rresp,
                                                      ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] observed_rdata,
                                                      ref logic[`SVT_AXI_MAX_POISON_WIDTH-1:0] observed_rpoison,
                                                      ref logic observed_rlast,
                                                      ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] observed_ruser,
                                                      ref logic observed_rready,
 `ifdef SVT_ACE5_ENABLE
                                                      ref logic observed_ridunq, 
                                                      ref logic observed_rchunkv,
                                                      ref logic [`SVT_AXI_MAX_CHUNK_NUM_WIDTH-1:0] observed_rchunknum,
                                                      ref logic [`SVT_AXI_MAX_CHUNK_STROBE_WIDTH-1:0] observed_rchunkstrb,
                                                      output bit is_ridunq_valid, 
                                                      output bit is_rchunkv_valid,
                                                      output bit is_rchunknum_valid,
                                                      output bit is_rchunkstrb_valid,
 `endif
                                                      output bit is_rid_valid,
                                                      output bit is_rresp_valid,
                                                      output bit is_rdata_valid,
                                                      output bit is_rpoison_valid,
                                                      output bit is_rlast_valid,
                                                      output bit is_ruser_valid,
                                                      output bit is_rready_valid
                                                    );
  extern function void perform_write_addr_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_awid,
                                                       ref logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] observed_awaddr,
                                                       ref logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] observed_awlen,
                                                       ref logic[`SVT_AXI_SIZE_WIDTH-1:0] observed_awsize,
                                                       ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_awburst,
                                                       ref logic[`SVT_AXI_LOCK_WIDTH-1:0] observed_awlock,
                                                       ref logic[`SVT_AXI_CACHE_WIDTH-1:0] observed_awcache,
                                                       ref logic[`SVT_AXI_PROT_WIDTH-1:0] observed_awprot,
                                                       ref logic[`SVT_AXI_QOS_WIDTH-1:0] observed_awqos,
                                                       ref logic[`SVT_AXI_REGION_WIDTH-1:0] observed_awregion,
                                                       ref logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] observed_awuser,
                                                       ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_awdomain,
                                                       ref logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop,
                                                       ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar,
`ifdef SVT_ACE5_ENABLE
                                                       ref logic[`SVT_AXI_STASH_NID_WIDTH-1:0]observed_stash_nid,
                                                       ref logic[`SVT_AXI_STASH_LPID_WIDTH-1:0]observed_stash_lpid,
                                                       ref logic observed_stash_nid_valid,
                                                       ref logic observed_stash_lpid_valid,
                                                       output bit is_stash_nid_valid,                              
                                                       output bit is_stash_lpid_valid,                          
                                                       output bit is_stashnid_valid,                              
                                                       output bit is_stashlpid_valid,                          
                                                       ref logic[`SVT_AXI_MAX_MMUSID_WIDTH-1:0]observed_stream_id,
                                                       ref logic[`SVT_AXI_MAX_MMUSSID_WIDTH-1:0]observed_sub_stream_id,
                                                       ref logic observed_secure_or_non_secure_stream,
                                                       ref logic observed_sub_stream_id_valid,
                                                       ref logic observed_addr_translated_from_pcie,
                                                       ref logic [`SVT_ACE5_ATOMIC_TYPE_WIDTH-1:0] observed_awatop,
                                                       ref logic [`SVT_AXI_MAX_MPAM_WIDTH-1:0] observed_awmpam,
                                                       output bit is_stream_id_valid,                              
                                                       output bit is_sub_stream_id_valid,                          
                                                       output bit is_secure_or_non_secure_stream_valid,                              
                                                       output bit is_sub_streamid_valid,                          
                                                       output bit is_addr_translated_from_pcie_valid,                          
                                                       output bit is_awatop_valid,
                                                       ref logic observed_awidunq,
                                                       output bit is_awidunq_valid,
                                                       output bit is_awmpam_valid,
`endif
                                                       ref logic observed_awready,
                                                       ref logic observed_awunique,
                                                       output bit is_awid_valid,
                                                       output bit is_awaddr_valid,
                                                       output bit is_awlen_valid,
                                                       output bit is_awsize_valid,
                                                       output bit is_awburst_valid,
                                                       output bit is_awlock_valid,
                                                       output bit is_awcache_valid,
                                                       output bit is_awprot_valid,
                                                       output bit is_awqos_valid,
                                                       output bit is_awregion_valid,
                                                       output bit is_awuser_valid,
                                                       output bit is_awdomain_valid,
                                                       output bit is_awsnoop_valid,
                                                       output bit is_awbar_valid,
                                                       output bit is_awready_valid,
                                                       output bit excl_write_error,
                                                       output bit is_awunique_valid
                                                     );
  extern function void perform_write_data_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_wid,
                                                       ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] observed_wdata,
                                                       ref logic[(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] observed_wdatachk,
                                                       ref logic[`SVT_AXI_MAX_POISON_WIDTH-1:0] observed_wpoison,
                                                       ref logic[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] observed_wstrb,
                                                       ref logic observed_wlast,
                                                       ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] observed_wuser,
                                                       ref logic observed_wready,
                                                       output bit is_wid_valid,
                                                       output bit is_wdata_valid,
                                                       output bit is_wdatachk_valid,
                                                       output bit is_wpoison_valid,
                                                       output bit is_wstrb_valid,
                                                       output bit is_wlast_valid,
                                                       output bit is_wuser_valid,
                                                       output bit is_wready_valid
                                                     );
  extern function void perform_write_resp_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_bid,
                                                       ref logic[`SVT_AXI_RESP_WIDTH-1:0] observed_bresp,
                                                       ref logic[`SVT_AXI_MAX_BRESP_USER_WIDTH-1:0] observed_buser,
                                                       ref logic observed_bready,
 `ifdef SVT_ACE5_ENABLE
                                                       ref logic observed_bidunq, 
                                                       output bit is_bidunq_valid, 
 `endif
                                                       output bit is_bid_valid,
                                                       output bit is_bresp_valid,
                                                       output bit is_buser_valid,
                                                       output bit is_bready_valid
                                                     );
  extern function void perform_data_stream_signal_level_checks(ref logic observed_tready,
                                                        logic[`SVT_AXI_MAX_TDATA_WIDTH-1:0] observed_tdata,
                                                        logic[`SVT_AXI_TSTRB_WIDTH-1:0] observed_tstrb,
                                                        logic[`SVT_AXI_TKEEP_WIDTH-1:0] observed_tkeep,
                                                        logic observed_tlast,
                                                        logic[`SVT_AXI_MAX_TID_WIDTH-1:0] observed_tid,
                                                        logic[`SVT_AXI_MAX_TDEST_WIDTH-1:0] observed_tdest,
                                                        logic[`SVT_AXI_MAX_TUSER_WIDTH-1:0] observed_tuser,
                                                        output bit is_tready_valid,
                                                        output bit is_tdata_valid,
                                                        output bit is_tstrb_valid,
                                                        output bit is_tkeep_valid,
                                                        output bit is_tlast_valid,
                                                        output bit is_tid_valid,
                                                        output bit is_tdest_valid,
                                                        output bit is_tuser_valid);

  extern function void perform_slave_reset_checks(logic observed_rvalid, logic observed_bvalid);
  extern function void perform_master_reset_checks(logic observed_arvalid, logic observed_awvalid, logic observed_wvalid);
  extern function void perform_master_reset_ace_checks(logic observed_crvalid, logic observed_cdvalid);
  extern function void perform_slave_reset_ace_checks(logic observed_acvalid);
  extern function void perform_master_reset_stream_checks(logic observed_tvalid);
  /** Performs checks on AWUNIQUE signal for WRITECLEAN and WRITEEVICT transactions */
  extern function void perform_awunique_checks(logic observed_awunique, svt_axi_transaction xact);
  /**
    * Performs check on WRITEEVICT transaction that all wstrb signals must be asserted
    * @param xact Transaction on which check is to be done
    * @param check_all_beats Indicates if check is to be done on current beat or on all beats
    */
  extern function void perform_coherent_xact_wstrb_check(svt_axi_transaction xact, bit check_all_beats);
  extern function void reset_internal_variables();

  extern function void perform_burst_4k_boundary_cross_check  (svt_axi_transaction xact);
  extern function void perform_burst_wrap_address_align_check (svt_axi_transaction xact);
  extern function void perform_burst_wrap_burst_length_check  (svt_axi_transaction xact);
  extern function void perform_burst_size_not_exceed_data_width_check(svt_axi_transaction xact);
  extern function void perform_write_burst_value_check  (ref logic observed_awvalid, ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_awburst);
  extern function void perform_write_valid_awcache_check(ref logic observed_awvalid,input svt_axi_transaction xact);
  extern function void perform_read_burst_value_check  (ref logic observed_arvalid, ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_arburwst);
  extern function void perform_read_valid_arcache_check(ref logic observed_arvalid, input svt_axi_transaction xact);
  extern function void perform_write_resp_write_data_check(svt_axi_transaction xact);
  extern function void perform_write_resp_write_address_check(svt_axi_transaction xact);

  extern function void perform_snoop_addr_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1:0] observed_acaddr,
                                                       ref logic[`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] observed_acsnoop,
                                                       ref logic[`SVT_AXI_ACE_SNOOP_PROT_WIDTH-1:0] observed_acprot,
                                                       ref logic observed_acready,
                                                       output bit is_acaddr_valid,
                                                       output bit is_acsnoop_valid,
                                                       output bit is_acprot_valid,
                                                       output bit is_acready_valid
                                                     );
  extern function void perform_snoop_data_chan_signal_level_checks(
                                                      ref logic[`SVT_AXI_ACE_SNOOP_DATA_WIDTH-1:0] observed_cddata,
                                                      ref logic[(`SVT_AXI_ACE_SNOOP_DATA_WIDTH/8)-1:0] observed_cddatachk,
                                                      ref logic[`SVT_AXI_ACE_SNOOP_POISON_WIDTH-1:0] observed_cdpoison,
                                                      ref logic observed_cdlast,
                                                      ref logic observed_cdready,
                                                      output bit is_cddata_valid,
                                                      output bit is_cddatachk_valid,
                                                      output bit is_cdpoison_valid,
                                                      output bit is_cdlast_valid,
                                                      output bit is_cdready_valid
                                                    );
  extern function void perform_snoop_resp_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_ACE_SNOOP_RESP_WIDTH-1:0] observed_crresp,
                                                       ref logic observed_crready,
                                                       output bit is_crresp_valid,
                                                       output bit is_crready_valid
                                                     );
  extern function void perform_axcache_axdomain_restriction_check(svt_axi_transaction xact);
  extern function void perform_axcache_axdomain_invalid_value_check(svt_axi_transaction xact);
  extern function void perform_cache_line_size_transaction_constraint_check(svt_axi_transaction xact);
  extern function void perform_readonce_writeunique_transaction_check(svt_axi_transaction xact);
  extern function void perform_writeback_writeclean_transaction_check(svt_axi_transaction xact);
  extern function void perform_axi_transaction_check(svt_axi_transaction xact);
  extern function void perform_read_data_channel_signal_value_check(svt_axi_transaction xact);
  extern function void perform_write_response_channel_signal_value_check(svt_axi_transaction xact,ref logic[`SVT_AXI_RESP_WIDTH-1:0] observed_bresp);
  extern function void perform_dvm_snoop_response_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_acsnoop_reserved_value_check(ref logic [`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] observed_acsnoop);
  extern function void perform_snoop_resp_passdirty_datatransfer_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_full_cache_line_datatransfer_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_cdvalid_high_no_data_transfer_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_snoop_response_channel_isshared_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_fixed_burst_type_valid_check(svt_axi_transaction xact);
  extern function void perform_snoop_addr_snoop_resp_check(svt_axi_snoop_transaction snoop_xact );
  extern function void perform_snoop_addr_snoop_data_check(svt_axi_snoop_transaction snoop_xact );

  extern function void perform_arsnoop_ardomain_arbar_reserve_value_check(ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop, 
  ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain, 
  ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar);

  extern function void perform_awsnoop_awdomain_awbar_reserve_value_check(ref logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop,
                                                                          ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_awdomain,
                                                                          ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar);

//--- Barrier Checks --//
  extern function void perform_write_barrier_transaction_check (svt_axi_transaction xact,ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar,
                                                                 ref logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop);
  extern function void  perform_read_barrier_transaction_check(svt_axi_transaction xact,ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop);
  extern function void perform_barrier_id_check(svt_axi_transaction xact);
  extern function void perform_barrier_read_response_check(svt_axi_transaction xact, ref logic[1:0]  observed_rresp ,ref logic observed_rlast);
  extern function void perform_barrier_write_response_check(svt_axi_transaction xact, ref logic[1:0] observed_bresp);
  extern function void perform_rack_status_check(svt_axi_transaction xact, logic observed_ack );
  extern function void perform_wack_status_check(svt_axi_transaction xact, logic observed_ack );


//--- DVM Checks --//

  extern function void  perform_dvm_read_address_channel_check(svt_axi_transaction xact,ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
                                                       ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                                       ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain);

  extern function void  perform_dvm_arsnoop_read_address_channel_valid_check(svt_axi_transaction xact,
                                                                     ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                                                     ref logic[`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0] observed_araddr);
  extern function void  perform_dvm_acsnoop_snoop_address_channel_valid_check(svt_axi_snoop_transaction xact,
                                                                      ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_acsnoop,
                                                                      ref logic[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1 : 0] observed_acaddr);
  extern function void perform_dvmcomplete_araddr_valid_value_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_araddr_reserve_value_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_tlb_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_branch_predictor_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_physical_inst_cache_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_virtual_inst_cache_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_snoop_araddr_reserve_value_check(svt_axi_snoop_transaction xact);
  extern function void perform_dvmcomplete_acaddr_valid_value_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_tlb_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_branch_predictor_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_physical_inst_cache_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_virtual_inst_cache_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function svt_axi_transaction perform_barrier_dvm_normal_xact_id_overlap_check(svt_axi_transaction xact, svt_axi_transaction active_queue[$], bit execute_check=1);
  extern function void perform_barrier_pair_check(svt_axi_transaction xact);
  extern function void perform_atomicity_size_alignment_check(svt_axi_transaction xact);

`ifdef SVT_ACE5_ENABLE
//--- UNIQUE_ID - OUTSTANDING Checks --//
  extern function svt_axi_transaction perform_no_unique_id_outstanding_transaction_with_same_id(svt_axi_transaction xact, svt_axi_transaction active_queue[$]);
`endif 

//--- NON - DVM Checks --//
  extern function svt_axi_transaction perform_non_dvm_non_device_with_overlap_id_check(svt_axi_transaction xact, svt_axi_transaction active_queue[$]);

  `ifdef SVT_AXI_QVN_ENABLE
//--- QVN Checks --//   
  extern function void perform_qvn_wr_addr_token_handshake_checks(logic       observed_vawvalidvnx,
                  logic       observed_vawreadyvnx,
                  logic [3:0] observed_vawqosvnx,
                  logic [3:0] vnet_id);
   
  extern function void perform_qvn_wr_data_token_handshake_checks(logic       observed_vwvalidvnx,
                  logic       observed_vwreadyvnx,
                  logic [3:0] vnet_id);

  extern function void perform_qvn_wr_addr_chan_sig_assertion_on_unsupported_vn_check(logic       observed_vawvalidvnx,
                          logic     observed_vawreadyvnx,
                          logic [3:0] vnet_id);

  extern function void perform_qvn_wr_data_chan_sig_assertion_on_unsupported_vn_check(logic     observed_vwvalidvnx,
                          logic     observed_vwreadyvnx,
                          logic [3:0] vnet_id);

   extern function void perform_qvn_rd_addr_token_handshake_checks(logic       observed_varvalidvnx,
                   logic       observed_varreadyvnx,
                   logic [3:0] observed_varqosvnx,
                   logic [3:0] vnet_id);
   
   extern function void perform_qvn_rd_addr_chan_sig_assertion_on_unsupported_vn_check(logic       observed_varvalidvnx,
                           logic     observed_varreadyvnx,
                           logic [3:0] vnet_id);
  `endif
  extern function void set_default_pass_effect(svt_err_check_stats::fail_effect_enum default_pass_effect);
  extern function void execute(svt_err_check_stats check_stats, bit test_pass, string fail_msg="",
                               svt_err_check_stats::fail_effect_enum fail_effect=svt_err_check_stats::ERROR);

  extern function void register_err_checks(bit en = 1'b1);

  extern function void passive_cache_check_post_coherent(coherency_error_type_enum err_status, svt_axi_transaction xact, svt_axi_passive_cache_line::passive_state_enum initial_state);

  extern virtual function void passive_cache_check_post_snoop(coherency_error_type_enum err_status, svt_axi_snoop_transaction xact, svt_axi_passive_cache_line::passive_state_enum initial_state);

  extern virtual function void perform_multipart_dvm_coherent_start_check(svt_axi_transaction xact, bit drop_xact_if_error=0);

  extern virtual function void perform_multipart_dvm_coherent_response_check(svt_axi_transaction xact);

  extern virtual function void perform_multipart_dvm_snoop_start_check(svt_axi_snoop_transaction xact);

  extern virtual function void perform_multipart_dvm_snoop_response_check(svt_axi_snoop_transaction xact);

  extern virtual function void update_checks_on_reset(svt_axi_transaction xact = null);

  extern virtual function bit is_current_xact_multipart_dvm(svt_axi_transaction xact);
  extern virtual function bit is_snoop_xact_multipart_dvm(svt_axi_snoop_transaction xact);

  /** 
    * This task waits for the last transaction of a multipart DVM. 
    */
  extern task check_and_wait_for_last_multipart_coherent_dvm_xact();

  /** Returns 1 if only the first part of a multi-part dvm is received */
  extern function bit is_second_part_of_multipart_pending();

  extern virtual function void disable_ace_checks();

  extern virtual function void reset_multipart_dvm();

  extern virtual function void reset_barrier_checks();

`ifdef SVT_ACE5_ENABLE
  // E1.11.1 (IHI0022H) Constraints for rdata chunking for AXI Transaction
  extern virtual function void perform_rdata_chunking_check(svt_axi_transaction xact);
  extern virtual function void perform_rdata_chunking_num_bytes_transfer_check(svt_axi_transaction xact, logic observed_rchunkv, logic observed_rlast);
`endif
/** @endcond */

endclass

//----------------------------------------------------------------
/**
AXI  port monitor check description
*/

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Ubc5UovD34LhQp8ABj7A9dyu1I///ViWv9apfJHvmTdZQghbNsg7Jehitdux8n+1
nb38dxppSGVLURWcaZjLLE0kuVfHjTPJBuaIfBD8cpP3QLfXutMcqsKM4aB2sg4r
hn7wHimZ/3NCO7M2O0vkoI5vN696ogUkHwt/1KgI11A=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 51003     )
TG4GzWtztCJ8XWDfqVIr8tCfgI5WcNJkHSyAlTKr3LlQZqEEs2jMc5Of3h4eGsFt
NVsgxT5CwsRkWEFN36gNVvXhCEBDkIghzGblP0aP2QHDgXAyU1ibul0MWCplQ0xv
hE/eXvmpb+yzVVPh2T8Xx8zcHiAcwv3oySd6ndyDoRYnVgFReCkA8sBI/hjm21Zy
jc1Fg0/oo/PItxojjVLRCaK6QJJAZuNzbfd+S0EIC/SqwoUnXfq4AUAk8M+iGlZ2
rM5c8/PAFXkEnbcykETgOhtcOrhVU8V/wjK8B6dj6EhhHMUHste9fxxf04nCgGmS
xs5uxBwnHZgf+S3Ir2qp1vOx6p26P++0rlu2fjzLo8mC3qZdbT0bYBZF9+nbxX8u
b6A9JoBP1cTgaFgwS42g36YiBBm9LzUThUr03JE15DzUjOoHCruXRLtizXeKkYkW
dvX5bT9rbjbuDABgq33d2kdWGBzFPWqKFeB/AeGQ7hAirU10exnK7cef9BuGeTZ0
nHfNrY2b2XUbRck/UABdvXsRe9dkRw4T4rymK0SpaITdF3pFl8tkph66iwa4L58C
rry8dSGCHM1+WK2boigDAXqXVotOVZGPcxMBV9KzDSPzIP87aC2qzDjnMtVNdrzM
aUCyPxIJz6m9T+q7CRGvGg6dBfOFMyRsc6vkxdARe9//fLecmNL9u8uMqnF/bvWo
cg4gdp1rQL154pgp53sv4p/d003GRTcGzArePjudTY7MKC/PW4BPwvrZbPMI9m5o
HBccgVsJdp4cVsCaJJ7AGXntUAFk9Aj3hAn0Ai4kghZVy6xeso8DuO7cNGpYSzDE
crjeENBtnot0rNE51JcdsfLAk4+JpJWe1P8eKfe/+9mN5/lLLy/FWqicHHoqvFt2
AoSBLYPpItLM+YQ68oHY2zk9/lThnQCAHoyGe0IjgrKby57AtAmBWl6TXnXeBRsP
rUr3ADJ5sa5R4HcbWOzbRsDNVOylzCeGIQFOlZFNBPQy6XlfWsNmbdJg7ZObra8S
GOM1SiDg16j+G7kQFYnBHRdDP2h6+OlFLn/ASWukRqx1jzuRIxRbZwEK2bNV9Fzi
KAvqrtkpKemIrFvoaDE/YkZxvGxcsfrVntw82G0NR6zzS4uNSfUG21aaovf+ebRC
zObJ6D8jfZgCQZOba9RD7Z1ZzBfV1qRM+ZOyWlL0KX8y9fr5vX3Hvu6VtX2ircCZ
1BitfjnZBti+Cr3vhhF9behdZvBRP1jjnwab6uhnllHwRMcsUA5Ubh8Skr/GLXxx
BSuRZUl78ino4Bc+ycpYmKuzvwL4tv+Y30Es5ZZnjG6DTeHbyFxknNQjgS2WUXpI
h4WiSGu/FBrXaz3T1sJdakrkhHTTFA7iZjxY2VsiyY77pxZNAWVKESGo72a3fI26
X10UExDZss50NLVrbzbbZuZ0hg4w4j4/p1tGcQqE99DEzY2vUdJkp1BXZozPoyZf
pY+YT7ebjy1yUBI+aTzPpExzC8D7ZpttCimh4CQGy5NZeRlO752OnOAU2LR/fJ3Z
RBkAeZlnMSziaJuIW5lbQzpnm6UNG8peMfTu+nQqy6AGy27maqJKAPrcB0Wg0iQk
flhWgKJ/xE7gk9wLgTqlnDTgw6vd6TRiu1QvIdMygM8adhAV0UGe3L7r7+3g4j+L
7HeSmm0GQ1XuZkkFkSmWT9RBLOr4+kom+ZWKwma6cgBeSVkt9z+J6o3Ww2iaBXR5
nL5bqSaT7NQx04KcZkWQskNiUcTNH7MRRMbOi0QQXRqCClvg97t3XIDAGZMNGcg8
wC8+DNcmuf3yj/ZsMWwxYjPiReFpaoOYlIV74r4Gi9WN5SC76Nt1Q2UnM1FIij7K
SGXyAizWiFfCC+w4VLpLsCNBz2lT/p8OxtNWY/F4Ef+Bj281qvPCQco9s848cyhB
jsZW8mZnC5k2QAsIEK6DUqcPtxIrhHY1GD7Bnc/hLONNXmj3+XoH9BRpgq5A9mPx
GmMs1Ww3j5MMupwlYWje98iGUMpy7EC2lpYlg35u+VnVaKiX15Sl0u+O36KmX0AT
+0qQ0RZwUrZLfZHmI5qu1qZmuE51KmQZhX9cAGEu9zp+5chlVZTkxK4W78AtbW/y
E3wK1dV3dE0Ss8TLlU83dQt/MLFDEgpXXAwzOG1iZ/fZ0FfhQGVPc1eh3ionKUvP
EZ779MpPAEJkGGRnO9CNQMBQM6gCFGLYrJN9zJHNHEOScQpM/mHLVMj9cbf27xGb
BQHnJZl9VQuctCmGv7Osxi90bc0AihLupj04iyETpOvCv3DsafKgyREyyaiK/QNv
Nxq7PBhhZeAOC5zD6gNa6pa+bB/VaQ/RQK/yMOzdGDnjos8cgLx4AKLvfGyUmcX1
xMY85jaoPyXkFgZ+Y5E+psBUtQYgAOro2uAIbeZR2CMpGeNzNO8JEw4ItZb6Rlwn
g2YWTuEMYUYRoKEjoKUODi+qDcUD1O+Z2c+QMCtTGgdtL21Y9ruV7ONF0aqZrFRl
KHxftnAak0PAJsLhnnFlojahTSwLo4k+xiIX/uVNTouL3x/KnhGJ0jgW3QqX1LEh
HkXYPJA7y7R06jUINja5VXpqwf9bylgNLyYRvFsH5YKyhIJ5E7bQ8k2sIuE0Fb1z
phowSo4YKv3coByDbN3StvSEzhQMckLjMSgYrbvvASkQHZNSWN25uQYThl2RGQcP
r9uRBT09R7hvktY99hFzCcnH+tF3DzC2ojWcUzfzLb21Qs8TBjH1BSCFT3Tw4H2U
lQZlJfUUpqFxvb8zqV/jM/VQEZL3hmRaOm1wODup7Yz1krW2xlENTMDelxPMW8nx
3xrMzz2NlQ5JFbWchLWBWLNJZ5cVOT7HT+MCZkCh6Dp2xFZT9qA5ZuYPdVN7z0jQ
53rKj5imwNvtgGWOn1w+LvVPkCGCCeqsREsKcRtaRd6uCHJV2IaRmqt7mtMUznDA
O7p67+1xgAulJGxTidg7LWzr45DF5+z/Vzi8k+aqK2APnUHS9JrC8FHe+gZXdpXj
yKQxTWxKPTCohFZsSYlRT1yMh9EfWJ/TFODN59jXbeCQDIvSdBOvm1YMCDSv3ZKm
pzSQqgUg7r2lNcMVueSk5Nn89q7WKzdva3boIV8Or36Ni2jy7yru6WK1BTMBt4Tk
vz3jC16qr6o1zfZrzypTr+197Bz6l5zeHqo7lKRIIhXdKlx18Mo/+js54rZVWmFo
IzBWJleb9T+HESx/kxxVtXugDBv8z7rChnf5yyMFX6hLb9SR0COYBaQpEaXV8OP1
aYQqcKSGsrzDgO10eiPy0UDrZW2QRrJE1lo0EILVw0sL/9h2nKV8OJhpAQan23cj
jJFPHJzvoSYB/M3RCTtuMNNnoqBbIg5uGHEU7n+3f+Njpr1obRrcm68MonmNBlBt
yzMf10Xd51HbzPP3OT1efcgksjsEmMlbzwgb4XsXbDH5ktyYlgPMpKGzu5sVuzWe
GzD9RJlmR9Bufm5NFzUaqOCI3pGhFE9H318NcNFAkNXANwLj37Cmr0UzbH3KgFXN
2ceVA7t6xIXS+sy4NGFLzmFzG9Rxq7JyP2i4Nfngd9wVit3hs8JZd6uz1KByC4Z+
xg4HK/ZiecfaljQSkVbBm2m/LO9i/YOrm3f7uTFsi8ZXv4zYOvL7/5PO722nZOsw
UeQQR9JZLi+pY0fWZ0Vje2asjn7f7Nti3o+04ekGERyZjAoBo/ZOyNWGZTP6wtwj
0eixqLSiDao2wSx84dhfVmaiihkOGKM+owThrCXFMAggr3ghGqLAee+YO1y8gMjO
nKP48CoUwhtF9gFSttbOTBbf2ORQUDhw69OjS/MT9EFnGm+qvIWRYVyFDqa4scfd
6rMAacfu0EOy8nhZqxlfFvgk1+tLq7rhpl8clBptvo6t1T1AtKmECLF5KJXvFzDa
liNnU+88mIcWLY4y79vy97MxLHkkIPQGGbSpNQuC2VO6MgCHq8S2oE8a/0jZB2Or
4sLQKpTIvq3Opk+JjVBisff47kHMLWx6T8n0n/GzZ2q6RBo4Ubs3eOOfgw2dt4aL
Sz/Hr3hVLqmjCtS1zKqgkeFt/C42NKXfJX3yDnxMHeSQKGFZHcgqQr5s9K+ymx+p
0xBb92roPtncibfKxrV/subk96ztWFpRTt0wpYwHX+DM0GveV+d92l2BcgPPFNrE
iCR1xT3jKBkFXTD27S47Xjr5EvPy2wM4mCA0ISMJOF4MwATLiFELNDD/i062DOma
QHvEtSWtEZy/Z4pxktzqKDOsS2ApBaiu8hGjJD+82XnMog3OGDKhJAc2MUkNBW5G
TPQ/dilk9l246gFp4QaVEu2N1hsz0oF1ybPPivhqPJzXjc24tVUbkzWu01op2WnT
9I3kb5PJ7gLGfrVqLLDobZe6t59bhl0YgXoq6+WSvvw1snnm9yceb1q9mnb8QPmY
9JNLccYe/tLApk+yYwFNvVLqAiqkMEw2/8uGPd514Dd0OBZ/KZq6XwVgh8eZVYmM
up2BOEOJbqB6ymdAPShc1VvpX3KOnkGwW2EsmWUFYlnTsGTuGKzP3/tZHSzwrPOY
a2S/yLhY9OvlImo8yNBQePrgLdJlLNsmZSW9aHXmF04RUo+d+BxCde1z3nWjULju
5yGXShiesxqIMgAxF9DyuOIvYDShdXoPzKpOXH08MZQHVcbaCJuyGVagrhZgDAzj
kZ0JaZRypAaZm+NdDF2N88GMIvxA/3bMJ08gfsjm6bW1YKYArAwrnmbKYMWOzlca
ghqmRyuyiYlFlPkBrr/EfcPMVynWVIcecIeE6j+eQ802VItsLWDqYRhwY2UXPvEU
h7O/raHX4eEHkw1hOxo5+NdFsjCMV2yewQbcEISpI05qp2EsQdy0ZL7sYB0EesHn
eIe/t6LmNYrHoi3lIlDEfNo8x89EynCYQclFInW/oaJ+wrsJZGDg3+XDix9KmV+P
Z9gK0WOZC/sMfIWVefWqsXfD5+aIK8MsMEkFlwUtRYUtfagcArphjGFCn+7Ar8rO
q//lC3/qHBOFgdZXB4uODKYZQfVZdqCIrdhonwkhG0eqzYqoACvnzaV/CnmHBUZz
694lAcOpMBmr/a9J6sQo6BUDlTkSovFvQfismzRQ0YIhq9KGr0zLPdyT/6Z+/aBz
Xdu1fWMn5PK3Yk1l4RaAjBsJM1jQJr4+r4o9AW9pqo/TooW5fzjPqN/K+Tq3D9A7
muG3xWZLukxhTa/svD1cl1I+abiouFJLY7Wo7xGy6LDDo6pYJwbLZoFkLC8o5eKg
1FLT3IUN10LEIKpjNAZKG299II2HZjDGPxmlDjDdkuNDMBKPhkYIjkk1PX6fjIRw
aj2CG2a9ZF33u8psJ2VJJ6N8ISZ9BkC9zS37aZK1jz4VRlSNKJso+eTiqAKOwzFV
awhkBiIhFanyNOW93zlS6g5eU0+2oLO9HT/CMOmZgIfgh2+KoBLtag15ZToxQznl
OxdGJlo00j9qj50akfe63IhG87kXv0qG3lTdIm1jbiVr4XyuQq7Jy6dRMM71WIbV
J1/zsGJJHBtCjCIS0rah7Kd73zWEBZT6c3lt6FJQPeL54Fc1XLKyrM6oXM67BUfk
ETo3KnhqgM/ecGDu300+cBDXxFDiDCE2tU2NAz1dsb5iCcFExO8E8ZgdGK7F3POR
/cg9YhfqU4+XLrRR1wf38IDc/Jfdkiivc1U88gZWkzrOI2pbRruK64+ToFgWtluQ
CNBoTTxGykW4ZXMIWD/weNJh+KaT8J9vOgaYD6pYrtL+squyQdnMj0yX0KQv4FYi
pHbAOpI57vPZ7CnQWFJWImEOOkR7/QOtybUa+Mf5i2vCI0xDcpjSad4xwCM/M5wr
ykPSrWvlRA/m1JjuTQ6lAhL3Af93P/EXwIoFK0KzaJvd/nMw2pz7FMCof4ruqQkU
fXhJsewGHGogHFmOKT3FYD02YCkrT5dGLicywY3yBUl+mOKRrOK2gk7gSTFz9CNi
69B11uvDwByOdkIteUY+LloK1VZ9DdgobAaNMX5U2awnOoGtV7h/6vTNkOSCeKST
sfRmZldqkWRpmjdJ1Xld1xeu/6dpXTV8tt7o+FShrICf+cALNc5p7jHYV0w9hyII
8rjZ5nd2KFArmSKFZPj+tY0W1+wDYhUkY42T+XQj52HjYM11G97Q1MJDVo7SxrVl
51V/oDRXBpqFTE9yvxU5MUgEgjJXqyx1sN8bqN7yJxmY1t4kj31paC+zDo0Uv4d8
iYj9dOUs1/X0qKvRJkOf+B93aVE37pkLDNaP9ldwmsIFjxFNw2xex22oGCGpT9wo
McCX/cGAqyoypA4p/4/mr4cAFLCKHL6VEwUC0IJWVVYQBLekd57EimV5G3ETMcCb
G4W8t1+tTs5YpIoRGeKBB4eXcXwXCl2/gwxfwUD31YBrjaTtybiCxEqfNb+X6ypS
vlXs9T62eFqx6r+U3EPeWipedsyaA69YQeSmjMoLF32ODH5JkEeT6994TD3dG93r
uPZNmYvIO8PnrRwMxNaMFF7J+xDV4zswtwWEWWNtaxJqJ3jtG7Xi427Fi1LEvZ3H
1d1F7FYaE01kMqCgK+hkziHpAiNcQxo3vRiLOadLYs3koNXRevtlGmUJqWfr1Kak
xXp/7sm0P09LBA0zLv6eIi1bFMUWXb401dwWqf5sEg5N+9kIXay/0SmlSotDjCqb
xDik5mpHdQmgcJVGkD3aIE7dmwzAtmY08csfYrcnWUllkI1YZ3iJ7AhvjuKe6Oty
147QxZ33oaxCjiWckju/6zVBnyS9213TT682yYPAriB2vM47Hix6RI7smxnHEGM0
m6TSVZmP8k379bHDAtSmTyXfhi+YiTsf2mmH1Hn/jVNxx9kU1wrwkVpqM9NNG245
kyWlYjceusAUHxWsIOfUtNxfq5CgvviWNRndgOZgrdNvh/y1MN8WICDNGSv8Mms0
jPRaSmS71WD4AoeRr9gEmER6jEXYuWoMmEAF1eXBNjj5qr0B46OqrPOfNIJuD18u
Sju1lh12/2CE7snsYWrd7hTOLIw0gMNpEulupZ/p7d8AABVC+3FMavLSZr3J05yK
rA7TLf+ui3R2neE/1Eno5SNs5RbwMBHlkKecj8MeHJ6ZXZGpiZEC0oF+l1q79oFL
/hUg/Hjmt3UgRPBOcc20GTtRLY7yaDLsqFmNbjHAL9fwVohhyjBrAh5XXgXoXaEY
E8TSj0eyZ5sP/iEKjrTv+NoBytniX7/GHeVm+VpS49hqeilBmh2o1MtsIH+TjWd/
U3ImG1H19dwcWEVrQHJzwywBhYcxBCUgQH1HHtOQ4gYNA4GgSun+IaGl0UZ25lS9
n0W6K11wkWJB1/upozzbjQXt4XrwBy7WpqVeKrk7v9Xnu/4R+6XiAVgyEFkzuRev
uKrYe/+DPVDRPeY8Yhf/AhlOndi7WjdssELXKdvl9YuybVgCyrTkIzafEuxRG4sG
pwCEqb04+Mhk2Iv6D5tRDMxWn3u5H+oTo5j1n5BMnhHOMyHz38nlpjVW49ZpnGs4
K6L4vUvdfdS3UKVjpGxWQoeLfvv7/6owurZBtpPUFV8KmzCb02ZOU5UIf8qoTwpb
mM7x+zH0UlPEVmpjKZ6sEB4s5Fdwti1YuAEosFLIJSLxFNLxQSVBDjuS+6KXQG6I
RDQfDH1eeISPKjhSQMS9fjuTlFX608TPLlA/XamOR/FyNAcDhKjQmqiVjjtTnbhw
lVy/1HYvkYlXezh94ZiSl9E63sNg/SFIaeAtx2/r4QH+fW5V2uuvlBSGXTitkm7h
uDCnigSLGYmvB0oavHGT2uwp4MV31M/6/DwZOpDgYo3UXTYdSv33650pFFGCZv0c
eruJvSllMSsIrw1MTT/U/uxNJExoF4/J/H+Xv0wyJCgJgaLNFCXy0MSK3bWo9KP2
xQAdXkjyYB2UELPzsF7Hp9Vz4ZbdkCZfYL64zLMacGRtmiOSvktmnLnO6CsnbvVr
JBvjoJIfzZ3cSBv6NWSWMYxzYJzvo9FPSdiGsSz6Per4n2YtNAdS17okVHFyGt8y
fPvRyOkx/iYt+aHwb3qZ3HGt/8xH7FCIOtZevNbp63RK2Q0kJpTsZN5PwaWZZtNX
EG2xQlo1CYgw0E5gZnQ22AVwns07+7pjZZcFQF/FTzSlJIkZxOO7HOoQIiGXlXVm
0F6APY+u/mdNVDcee0XN8ZAduL/3F7VBwHe6SXjFMbV/bzLXNJaYjMtIg6lcmvL0
GnIEVc4a8m6fj6HR6DiBJ1R6TFOMMu62IpGAX30VKhAei5DyAebGZAXIIyTdf3ES
vAT/SVsWjk3zKcjD7p/p3/RYl6I6u65Low0q8ok5C1E+ykKwFMjwRCXjLPmJgsIv
iZny7tusFK8dCVXov5gAcZieGfFMIlerSSVJYf5iFamQicpVOT6/SYpjcbbjNUsp
o81gxDIwJPe1LY5yMQiaDNsuP6vl0o9cmrdTDjENZ1p5y7ruvTm50QJBVT3QV1C3
DFdTXKzW7JpdB+kRRt68toIPsIQBYy5ZWY9PVa1OW32wii5/3+8NdyOIr1Y+skag
Kgn2/IU9c0xoHLa001Q+ElXvVFVAU7wUWG8nTYMFi0Uk+Xz52VmT2VitdZ3Fdn+Z
GUmeaI11LNWrz6MLwuOXm/WC+k6BMBZmyHeLz1X6CKMcJpI2WmjRQae8vBPp9KwR
VV7lPVZSw25oXxbs6a7Gk163fgaJlA5Ula9c+yJW2V4LaZUkjH7+BQrTwumiPf4i
2Q+cTP0EGtrqQK3GkeGiiiSe0esVhXCpKHIT4OMeLhrln+BZC5ZtF2VsyBISzMbp
S968jwULOKL5IMc4Vej33Jxt+hE79WR7bZyUi0gmwm7XNN4JmEYHB875kD7p1Buh
GNQWAz4FMSyC/Sj/VXK3zcTAwA1JJ/k2J9x6y15aMBo=
`pragma protect end_protected

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
kdVgbWmPuYCl5hJxGkIPZ9FzcYCC3W45xT0I2OQ/7Esp2tfi++l5fgRein/k37X7
lJAyOTtYx6cZVldKVlL17FA3Kmywd95Alryv1t9dvsqnmANnqwWdvyK7u1OC/Em7
XHMNS82Snk5lPjfEISN1amkBHMNofM9sDl2wuIaXXsI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 210837    )
Qz+Vid3EI70wL4BlWm4G1n5uJ+xyw+urWG4/Ml7sRR78AC/uF6uP4f6GBrVAcPru
4Bi7O9NPISh1b4PId+8M2uUpeS0r2XtqKx0BQNCo+SE7p/8ikzntaHgHB2mZTU7c
45d7357UOuH+znlxK0nGA+E6RY+V17auRe2j3kj2HZ7uEIXvCq7XHpnwSXuVIqhR
MjFHB1ZctuqL3hB9kmgT2r2E+pAu/kzfKAscvJBOx9WNV9mTCCwHqrH8i8/YAS9w
ayqNDGRiUbFiEeA/K4PjDGKFthqFa1l1C/Er+pe329ozMJQB5TFAKlY2PRhUic13
95YeLIV0CrP9oNkMA1g5i/QVXlRE1w80oIkn2nJrl6fhyJDp/bpL3TV2eYVdAZv3
4Np+yFuFXW/tsxlGOWt3hTmG8GXhRRO1xwfsT3gCBXIVGOrp3q2i1vdMltghO9Xz
gk9+9jpBgM461iVTZqs/i/zRBEmWwsps07Nki6U36Ml0dft3DV9r1CPBfj6uyN0m
zytF9hNxZ+2QUUgWx4BQ/j6XDpsxnYXWGO03m1DJAsXtPJWDRRKt06f2QKeBv5WP
ptuTuABZ0O6Jp1Rbshu0KM8KbabI3+kv8/yerSDh30wnYJ8piXRGUumz/OzRJOTO
l7g2FHsUrVr19G2VzO49zhiHcmSlopdMnwdexyBqOO7LGZaMMzdGT6rXaWeSHDYd
oujDSPESDf6RKJObcBZZ1SBIcz37NNrqrPZvBGJGLTPIZVLSxhN4tqPAU3axas4Y
p5x3JalPpd8gRDLJUZTqXtWGiGsdnASNrXbJbi+h3MDIo92dM8jWv8un2ZDAOiKe
fx/eY2wsdTfk70GzunG2K7fo5c/t/cAU8Rysj9o4UkgVjFeCl1tvCgPptBoFiRsc
6EX14pcwbrEyr73RaFgJszw/5ltLGIom4qmti+FMjbmTcVawQaNnJ6S8H4JgRBAK
UmFi080v4h2iRP3R1JHPcHO125MAIGnsY9LwrT9wxWi804bgD2xNuq0NkkM758vz
Kv34KCeuCzsh9YnXr9vA+0mgb3P3T3ofY83rvYY+AJRpF26jqlJskvSrbeUQl4J2
/9ACwDYN9RxUdl1w2MHYsyPw9ad/4qz8o2rF7WdpXAnp5CIxKI0Dg0N/q5BwKt1F
iotV2L2C55Hyf8Ygd9vcFKVSz4aH4D155QGud+yQ6adW3ITHqSPxMhRg0IkfslEQ
sjfbExDRlWAo8BrStFUr+6yxI7b6r4KfDG22PDqaUZqHW2x/tn5MqRgZrrm95j4m
jxUfjS6Jhb7q5JwanDsnXkFIMCbYoArWS0KlPpifaQ3LRu5ohQma9e2OCXpJwvFi
3MxJQI9f/BQL0uHqcNHUZCN+59f0OgIfjoJe1ShFsGUbCo5zTR/GM9231iWn18Zc
lpxNJyOvJJj23nnUV1sD1jMWATwkhVnu/AGHA025XZ+9SR84NSf/81pF5Ysi4Z3q
vpzWPTH0VQevL2+33mxAAAiAto8mUArCENpsUjEHcagC+xelenxCj/vUkdZf5Qzx
yWC/2uSShZ85CiiHbItxFXxTjPUH/jZLuCVt/JyHbyonHWEW0opQGLQp2ohpexqa
z4qItvcLFFFHnpnYRqu+W8946t0FE4tMU2+8qjgnydjUl97O9aCJfvAz46DLoJK1
G1wPeyZE0mVrjgBS8OQfYUnnq36ZLsCmu0NYlDv1nMv0LTB0eIkq655Rgah3HYxx
u8DdRcWoUvdDpP9aRyMB4hU3R+Aa3/xL/QBzNUUaSIBuNgEiarK7e3nsNn+KZK+A
7dikq47127t8cGkTcJVpBszPpVdYLD7eHqwo9ABSpDoufcRs8gQtomnx3L6qqVhY
P5LrRx0zvgaTLW74gaugAEKXwB394lZua8pTB+bvDOD/0YkrrYBeRVfPxE52iW/M
Ow0tLZ/DQSq+oqwfD4l81r1wRD+aGNVyL/+cLvFzh2rk7LqolbWqklTf8tsUR2fO
w8H3k+E9jrfi3BCK0inN41vHPB9rHNVCt8MMhfDMAx4FSObxoqXYpiXBrrA1mJBA
dti8T/TtPmHpKsLpxTPVF2xQ57yxDP5K6N9EvTxsxhjAiKW2S9VQYP4PjSYJy7k/
OqhWBfrnfWmT6RqyvC2meqI0eT64Bx8wqtulo0M0L/zvFucjtR2rwqGejWp2HTpB
e2+JFZnT9gxM0Z4wMvuRAKgL1lFxCAUNXurOsblEzARS/AlkyLvQe0/uu0e0wxm1
/qB/FwdauZ7ttY9LL9q2z/VhImo8JBECAmhc4ZImJyIjKuZYNKyXXJ+P1xPFb2zy
Cl6kTTWbdAXKyT1wvp56ogaWcbl4wX4ZFDm7Lht9xbAVZhfthKjDN07sOdWCOvnE
USPyUYJNSftZC2m9CgcEkmRqE2o+S8uvph3CckxFxyFF4D3fJ0Rn+gpAiJLICVHZ
s8MXeN8t/iDnTU87+klpho53sSm27BI2ryi4I6CaQ2DViBiLPKIrfT/NbM19HNWi
4vaFothm4HhMs2eaBtKPC1Iri+93MIWPCogRCMCR8DqaYRH0Dc2pRhgXEbUYIDLm
n85wnpcPPiX9XMkiFaPvO75u39MEkFZ4VygdsGS+LngffmhfbZeOR8+fBMSYdjA1
O8wEZxw4iPIJLEccgGhejzDr3Jtm3majtAUqkTkQUKgM+j5TU7uliACtNuC5TAI2
Tw5libNdc+MTqhJ7+JlJZJFv3cYf/5IooBXbNkvfCYDIZo1QC8jofiTwOYklLui7
B+/2tgBCEp7aw+c/TH7VFCsRcJSBS9w4Jn0S0uEqWcSgTNr65NYyxdaMGBXde+UY
nGkTIVhHWyAHVTzI1xEOjAjmXi0laefCViAtX9hYikP+jOM1WHITA5Ln9AtMlKbD
MkPpase6u3BLD1g3Pnv+n7QF3kRat+7AJLYj0OcxPsVgdzqS/x7HU1ETt1210uA5
Hh1CJRcgQqT3NU5EuWgX+qi/dwsEkKnOZzWr5F0GtlbAbUktuoe5Fm98vNl8kBbj
/R2F+8DwCqPAwhk0tdS4TJf4gNCcBKLA1xlFrqKkwDrLXtCtCOORC++b93BsvnW+
MfmZSAvNT5jvlwJ9CUmsoQAW7ADY6yfJTpq3RKpbyM8Uk3ddUR3GyslqvclwLpA1
c12i+zR78/0yCx3/DRwFnYGMq9PMIKQvneyEQy0BGqg8DM/ULvIXMqD4Ytinhjio
Y2CCe2YHFiDy0kWDS8XpshxhhYMdjYoLuKWrq5OLHMvw/RyrRNmS23bC1E7ioA5b
/gMTj+mANWyIVMTCs29ujRCxJetffSfy5KJIDoxmkCTuiOQVE7BV0nt/ceG5hPrC
vr1psRSyyaFhak8ph5NeS8HvSKbZbWFOhsH6i3ui24RX0OzTQCY8J9DZ3vHYipFF
YmLrJruTl6mE9PMeFoi88wcSCbFOCPA4plCSJUFZ3Wi1lXHKUWpebtma0uSHRbxv
6WchDQ6IPyUG3W+Y/laMB9wjJW6gV8zUlmSTYw5VHtJGopvvOntsxBhKA1N/H+53
uPXSxagZEHjnwT0dX9U/UszAvJFYM1ON1hBzem+Qm5COn02o2bbXvzkfO3bq0Mgk
oUa090iuB2B9AvAsvqccV4+1XyZ8b/kazWMVmRPoS2Ko4MKeWCjwsPZCfhZz2uPE
VFHZYqTmMGHHDuagWamRwEGXzoo8zKDP0DH6HfhfLUKiViczt343CX9M6QdpAxnk
/57EUUB2VCn0RTkSHZl/84D/x+uvsBd46Z8mnA43G588NjmYw6L52JGyzq9h0Qai
JiMTtX45B3/H5a+120ywuNECmzzOIAu1NR/HUg+iLn66DzUs7//FR0rG4yQBHf7O
k9OnSaBcBdjjabGk+JQ7OwGSUpTD0AlFQncKGn9Lu3AWq6pQM/qnNvKkaP8NcxV8
/0DvsV99JNRmOWBpvAsTf1AscREy+vn+2H78jiVh6Ikg1oPY1avsvTPgqIrtp+RK
MoAXL4EBNt2sF7M1ZDh4/LcOmSDYeFi5uvVIUmoVraq/FKQ8nRKMM90pO3K0xwsV
KIGiPcQRnil5dvBigNYE3T2mROfy9EH8Jl7pi4RUArbMLXtkMxqKrtKgShvI+oHR
eQSPWCXbEzmMDsfhvq8jsg6vjOXxjQPoO8JmviUV97T4jgKyoBJLlHCL8s7zfhxL
LwtOItMh4uv+4v134RCuWs85I0vXdzDmba3pNF7rALkss4jb9KrgwGBpndDkOy7i
XjIdCYoj8gOmez/5o7LPFdy9s6///V6GMritQGqqmRF1iTxfUiDj7o8eJf0xJzsk
40A2/wlFoTAHK1lzCSIX+swU86X6MoHJpPtbWK7PLxTZSkH3oH2hTKZGB7xK7FD2
UwqrENAEsWcBdOCnpbZMFWq1cMVQyWI14esqLR8IQiSFc1IhpkOZdxWoI9dd3HGQ
PapfXYz+9IOlytHD0Nk91bPLbBC/mbjuz6MDnWEHMSORjV561r0HeXvc8mDbbyDb
uiPVOZewrE/qOzg2uw8mmhiMGrH8vEyH9Ca6BOCChGL+fOiGndSFg6w7bni86d2i
x/t1pOn6I9T005QLhaxVX58s7f5LVnVFnB/eRsK835zCPXldCvVFAph+P0XiE7g7
Vg18UKvzUxH7NznLdW6BqA0mMCeLyAaGM7XHUHNhELcZVqu7jiaOc5aXHSFyVjh5
RlMvGdiVaR90VPNKEOstgmalXLBGdrwpPkrbpJIIqrInuiB5IKE7YjHsz16aJnk+
se9O5LcUdNF7ps4y9X7XWvmxAuvqQjPwmNDKWUGzN5CQXrR9g2/NgULbuYvknaLs
fXhGYBXNSVvSCLAc0ClMQtxkkhkVwtg/GHxWclM164oDmjha6c6zdRF6nmiRKJyW
vf1YtsHWFNQLmBAcDRdWPambYov8yXaFW4jBWFsbUaB3/IJaRt1qhQhnSJZ6UAWU
OVLFcje8HAO7VQDcx2xXpf+uzG5PiRcAuT4HCvyQGXIYDeBSAlMLZuQJ8xWob4pL
mgkXYszC1Mel0tEhPeBq0vUCOLllKnxEubbnenDJOpfKcWsHubbiDJR79PnZfQrc
3ENQs0p1uXxH/aSL8vrdhbVK/13hgxjaISA99iljsSTZkl8SP9zBArX8kzALLbm4
2aYuPB/QwBg420r6IROgGGeTPWPZZfgWVAvuZenkhl3/WNi4l25gkVlzO9va8Gac
m1wElZLqpdVe0xnz73pgpb9zvtw36a7wdpLLZpzwCQulg4q2t1GXPJVrt+syir+4
Pi3zUzKhUFAFZrvuqtvEBRn5U/X3X5Q7Wg9YsY8VD7j+4irEjN77Mjh9u8XOnjEw
Fbl+5ltfiaSdrz9LaeQnWDxc0ryJbk5L91c91RHgBdXO15Gy2dn0ds0zpGDpOfoQ
WP4bhDDxwnLXaztsiRcztcSUfkHto8z7Vf9K6Qb7pQjF5Ix/gQEHM3f1bqZrTewp
ngjKxmCCLcljqoCwGrlD2gz49BHv+YKQ6tLmbTfIqa6vlGEgUk4p6qcMqwaxsEoT
q8H5IUV6JIGnBmEFaCrnA1rqsE7aIy65vWkcBuyyAbQ7JEXm8orwQPTX6/qnr4cC
YNvoZw1gOWFlwV92WlFohdQhGc8LGcgW1N2MmPIuET4pWw7dfN0rugcOqT0STZ8Z
Sh6AN/7C0lj+23NVkbkd8HXsrk5ccwQrlMJp2hRoqXUURGWJANg17NjNzWNKneUI
ei35pl7PFAuJQvsu8HdxpFqlR/daYt8U026jQH+PE3sPjFsKae5B4J0d5qq/KW89
GMGnQMSeB20gj0jVh0zZS+gcy8EdpMlVI5QJ75WU3kDni6vFYkvFo0cIhGBrXSO0
ILhzXKBYqQ5UiEtqRMVpw5gpf22vIKi7ZXNcHEg9dGtkGcgoe6q4NsR0nhDv9B/E
XYBrj3CoCLQdTUbyvGkcTxGqADfMfJJFM2ZUlAPYwcP91+K/jTN5UhqQAR4IixWz
PIkNrc7IeaYrpvfon0ZSAIT/a15T2nn9vrmjb+FDEXxNI5c0CvNFEXSYwHB9KXTg
EViVHAPhP5sebwxGaDNTUotnCnnQBzGoaNWespi7xTDKNYB0S7lMN5OeNrOzxzjX
WJJa5CdC+sqeUa6b6TXq8oXdNZDIvBtZqpxmk6I0NS3gUFMnVfPECx+9NFGQbv4+
2hzxmrLOqjhMbV0UZ9+AcINgQ1re4IdOHuKwRDuR8DzUH7vu94g/y1c49H84SFk3
7jnpJzh/FkvR5brRtcwsaZmIrgInhnSzP+0X1DJrxze1K8pRGGzXVXOWbaA+Ks5M
4JZuXRhWW/KO1NxETlHHAybZNE5BVNM8ndenaqb4M609cOGQ9wa1ekO1U9PYKaol
WsdDBsC4YnGvhdILOR4RkTHr0HIW+LgAErfUlIyXpQqzAmkgA8Wr1/2USmj0rtwX
qAHEVPkcEytBTUNcRudfPIYK/HH1hK6y9kOSa7KN92l5xbeDcxfUSaE8m/zIgCTc
7ONkXqp2ESlVgtI5wjOvY5mofddgNrSM+xcWwJsAnj2hFSmzfS9tvUHAqFZ9gohL
emMSbFnUWR2qrP1ZcBuGUl5bVgtTl/bO3X+8OORg+J1jRVJTuCjR2dWMXl4YCTU7
snAuSjQe75yQeQAU241pvSbt/rcKjQ1L0Wcql8+XwReg1UVWpjm4ceMSE+PM2ynD
3dnLJrsY2JZ6GF0O0Ckp5Hb2+vAdGdH1LdbiNpvC8rPznk0HtCq2UeipFsN6BXja
wZRX4pGRBNQb6rFNohWgWGVaYhLiMtK0yPgLyyQJTRWTMZJB/McfaQRu/fKHJvrS
0RSRNKPCm8Iqio2hAFO0jCvH6Eikt30Md339AQD8Cm6O8iQ+iziYwrB5zPcFvQA5
keGik1BB1e0VTX70nZYS7eFTjdbvrdSCr3S2sBqSCukGgJrCDlArZnPbFdnin0CU
wegooJQEpEsq7ScC3Pne4Dgkf0cSbLNJimkWVtHGzb82SIJ2TL3o83XwZL0waS9M
YZj49lxTuzeObu+Hm5d1pRUcKevkbUeyEANyUwaoWLmIT8k/JmHKNfoAJlF9dW/K
0X/p+PrCS/rezmPEzScT2sytEU+xyxuGKZ8LFqOvvx9gYk2s8c2oyBZUBGvEwakm
GGZW7qOy6pEA/5T8RhmGAt1ff1ma5rT2SrA6TK/nWELn0qhplQw/Ee57LvjlGIXr
XLFSljuff18WNuFxbr721L8v67z/Oa7XkL/mMaR8w70GU9/nXI6pJyMKSsiJcuPa
YXs8PzReDi55gtI3vmMH1GPRLRatKQgZq0FZBzY0lyX1vv/UrhCCQQ2OsEKIne3G
wEgCs4GGoqMH4jSs5XHrgdTfhKQeM2p1IdI2T/1ypXOKs191BWx3EUNg6pLSGvn/
P4eYK0f3MJ1dLrou4KztOBgGE40SUyZNtiC1Li9nKjgDjV+H8PfmsLYPj94aTHHY
NV3czcMFeZPbJQmWG4Hdnndi3ilFZPDoyHesQCbl0gQuePweA9J0nHjI57bn8Mil
ZZxvjHICbOwu4a+fLPknsF9turqzDgiJ7m8HQQw2NBMdaZAw62bR61ULj/2CZdAE
WlEtL/eBYizEJGOoZMJkcBSmf4dcJaI2m5zV1g8TY39Ze3c4Wup9oPpsKcCNPr/l
YLpvKRfNp38EYLOKI/7jJiAGTJVzwXAsd7f+w+QMpL8oJGtNBvDnqwHDacuaJntP
a5hMUE9haD2FdD9e2UgCjHEu5u3jmSUTzVvwjELsxlg+KC8IkgpsBxhtrmFCqr6x
3fyWYceHO10XcgQQPXugsBU5nUhqCRutclZZD3v0CKU8rRhsLl0iG4sspscltEND
pWP99r86+2QXMNYe2rfuqFttDxt0IG8MhGrUSU53fmgiNbo819/YvU73sByiL/aN
/9X4AHae+eMNDhW9cuk5rPNCMlGj6xk26Mx4kUYyRE20xjKSBfy7QAQ2Lo9qH3Iw
9Qy05xbnxIShCKWBbTQ3ZlNdDggpjwaVI25Pb8lv7CxSEtfz8NhKqiM704anhZ01
rL7ZYxu14ZJkAszU9rkIu2WTJ84Vi4Fgf1dLlse6d6AxiTxMHs2c984MJ36LOza+
IXiPB7MjMXQ/EYAlvtEQ/2FLcUdC+Xs+WEJyr1vdQCmyXfqMjhS5g7digZd1ZoI6
57DgpHLv/Hu+yJeQvYom6xSpSbfb8lgGc84NIUJhUFfRCUZx2oD36jvbYp83LnC3
Hz1lU3OlxvnKiW8aaAFR2EWox1sqZfy3n6VpYTo+A2V5Ph1RPf6ZZlFqKiqn/Ty6
TNWmlttTuUfhAcSWUNn0MLCeU3Dotvf/gK33c0jh2PZIdthbIixZXhHHSNbDDEw7
Iy4wivlXdcLWH3DeNMZ/aOM4yxhOQiNpO7VYXh0HxQPzsY0Np4pnemPTR8sq9xgp
/VsC3r3jLnt7AY0MTPEqFlLVf7DETHhVsb6W+BVMdgL2sEYYqBFirFZxZgB5smMS
jarguJ/cc/IjNDpOTeqJGd3XYN/S2f/f/EBRl7wYaCJJg8do+g5tsI12UbduQJbz
iCv+HG6SfXd+5AvrlB05KSzZI7cVpemA02FClYqUMtI+8Mfe3qSdsDty2W+MV2Eu
qtNAhKm/Aa1Syp11vwc+7c7X2Lc8Z3aOqOyjJmxgMKQccgU5EmheePb+MoE+cKYF
7+gg0YubWSUmQUl3zJ+eSChJUYTiPmkMpR5aIPxnyF6DCqFuz0HSn2ovm2BmQqeQ
bYnXsWf93Q2oSyh/smC6qm6cL3h1F1lTKPL0jviPld+MORfS4NLLVNZEaVdV2lE/
DL/fDySNfuQSzflvf/9bwTy/WAsAADaiDy2n7yysYlh3NlFsBMH4VpPI+fuizTny
68a0/jaY7UyOXfFZdbFTVrT2CpXEJnC0dLhVllXQjLIbZjJMERhiVLlp5Vt1jwG0
VEhwDa9Ve8o6XNTkP395/sLO8KsvrKiK70AJfmpFROriaLhyJN2GrwR86PxLT9CD
oAVnpKypPaaX9PVOOcEAQjnvddL+JeK+g6oeCots3JPa0Xp+fYviie2Ezyp2f8vT
+jhU7mnjWbmwWJTJ0Q2C+kaYzPnknKXVr+6RsbQjIpX8oR2afh3y2yYDuOVkdM8x
gYQvqrpmQm3rRVP684MJ/toHpiUFRQxWKf0rSA3Aum6DA/N+kb2V7HKL/JCQEhX8
Qx/9/De2bodXK/MRmWOUWg5DPe5VJ4OBXiEzXubTtAKrRqdsbV7JDWVudplr1RCH
37ET7ev+lxUXTk7HKu1Y8mupaf8D/hW6UFlUKbHgI7ozBatQRrWfTjDD6dQyKvTj
5Jbd2zmTrmtXv+HUtTu0R3eMdUoUzzJoYI8IUtRQ6BDcbV0et0uIN13cyneSvUr2
7VYaC/Oc1xfqxmmArk2CFld6hwIl9P5dZRpAFIzmEyAlHe4qRgX9tLTVZ+2DQx/N
GULtjZYVLNta8Bb+MwCRC4PXQHWFY35TrzkF9A68VjYaM2BmJoufI2zkaiMBmavo
cSdvkNp2NNb6GcWa7aOPAC784O+q3f38bakVXOihEbYYKGK0Lgce9qQFb0jvE2wF
KgKzfi9Z1rz15dC6FwwyuKEOysp5Q7cYEVYhY8gh5J6VkrbU6dznCFdYjeFa8ujG
KsRzFFKyJI07Bi5t28wVoZioPcl1izqFYCiviMQUpr1OtQg8jZU5kKGdlIW/1vrj
qSR98A81C9TQq60PHPTkZEPeUytZIrYfrlDfnG92Wi/j+UynY+WfqWOmFqHl3y90
PV87A0x2xYsHM3ysCGJg+A9DvL3uBNn74G/q80rl0LhAg7xRG6hflxqQpldeRt/Y
UKDdE1tTEWJYCBtCf6tZIIAYORZsKwPe6RLQQ4pY5Q8CRTauWEQaUqc9LWtquXSC
yX0swpDn5w9fXqknz3wmcRoRU8yKeL/6ZDtxBFjF5RtsPyfRKsRRbl7TawjXAGZ5
a8NXg5/sCh8ZMWNyJdUfze7GjF9TysH17kKYarZ5LIGP7rzAX98GJ4UGBh0DEqFX
bAEnR4+A4KyO32C6UtkNtiSzagknjrTXRcNlYHqOPhor0kNAi9pLgbhwkD2bzx6R
Uovnm20JA1nMCipWYI6AJiYjDeJNppBiaPtIG9ExyhDkcnp2Bkz9aPZj9dKmEgVn
OxBI2VDWcLkOMZPRA4yG19V0V3QvSZOaG9qjZDupeZQaFSkS4PznYdQ7GDLUkCP3
2KZLXfl11bOzqOnXplgtNzjisj/1eAJIbDgjHc8ggCcD6Yg3DYD4XuH5isv6Gneq
ANNKSlRfSjSGSOS0C/VRdde4zQS6GReUVKEznEVBFIEBx4LsH3p3sPLrQByoXZhh
WMUbq6sWsjwS9TTSQ8OBW1lRwCpS5bUhUCAOFPMLCTlZ2Kk3aO/SjZ4pc3a4ukul
V4cmFIkl4Qg7iGK0Pu+GoP/Nw19e9Y9ygLerGwe66gc/YEond3g0BDnuFMdO7me/
z16wakBdj7sT5ws/4/anwKJ7+qeBBb5xodEyRDk0FnCqVzQfggn51wFwElLb2IdN
e9AvoaB+zio2E28VkXGPsDPOj5mFfAElHKXN/ywtPL5HuPl8TgmDuvAHZQh0mGfI
zphLwltvKuc0CeSw6vDvjjfyySQeWlh/hUfRMZJ4S35nYfyhEOfji5RVfO6HkAbk
uPwSLgQOn6FQvQwqOWNOoFeeUwqcg0+XQEdEUJqUd+6oaHCGaa2WEMvMjkwl80Pj
SNqOHnO2bj3ojkLQTp27Bqy6hNlXgCGf/iIdE072FnSd0Wh5IT7R556HKtlAE3P+
PBSK+B5wMpxQIvlnYgWi4srax8l85NDJ6exOvnD2v96Uh9yKGjvdI3oe9Zdu/2uC
om/eWqEwuDFGAJWOTPT3kFcPJ0L5JjGZRbUStXS4rDhTu9jQxNL+Y88678j7D76Q
ma8MUSKJEAcOpT09/GqasiadNkLvtcegmaRnJJNKTd8AJCqdpq6HPrcjAEB7udCM
Mz5oi7CXD/d7oAzerqi7D098XHGmN13Sp2qVh6j3Q/yPWzMESy2SRnoRwruSmsgJ
vbehyQLNYQ4VI5ubZAeUtJdWnXLjZf35AFatwHUkS1YkRprUFnXQkmeNndZR3VqI
2ZQkuvI9ieDhYgffP8Bpocob9bEulG5rmsU0JOIzp18uunDK2sslbzFk4bhGED1l
MAJ4EzDVG82vQiFHNAkL7eNhWpGWO3TA1Cjm1kLq2pNtH0vUwc4s/Zqfv7bdCQn5
KhfyxahudAEIMVv6L0OvtR+O85+UJwOGewaWpoH5wMlnDsPNb8uP2vnpU0B3caXK
2j67qMh4omI5H7zwHK45jWthMx2BV/p+PCH1qhCFBv3llT356KYgSh6BkUF7QS1C
22xGwHRZ4rq0UxzlFu+9JKwyI+ukOl3n2S2lKargTFwqDBA4LPnzxfspOp+zRfka
6GDixZKurkyR3toKdTxWucVEcbrCQkpUfUTr7bZHTXGfNN55qu73pXJZbIPTjQbM
e/0WbSQUNWJAPAlmrCHRh2K1icWQkUECc6VBjf7iQZS84UOHPkTnm4vURFT+hwQ0
8B5o8+vMpFFm1KKBML+hV7qb/u5tEJIbrn+RtrDmBpaCj8Ppq9fpYK/kWKkUxnuM
BysRDOFhxh+A/5I0ymlcf+zxcRFaOi8NzSJZ/OvcxKhPCwfwUCxvRp6rC53et2h9
8C5A4BrXE+hRSyI1Wb+HRjjrVSUBa1C8hhoTVTLL4g6t7+pI6ltKoF7U4CTwdTO2
ofZBIEhp3Mb1R83lSJbpz0ZLjVIN9EvXrVkRSvMt60XsY7fx+AA4GknSsZW005JU
0/QhhNkOCD3nmNLsFmSj/y7bN+EKzeZPkysK/9fw/FvAL2SjLpWhVfyawS9gqwm1
9LUTWBArjvecGusglZUAyANeDRTXDn8LqXlVtV7NYv57R4HGmVdPh1ew2Yb1wJoU
WoNVcTH8brfoA1d4otigeq0ALiBF8ZAkyfXLQZnBHn29E7ZYi5o4qHi/DKeBOl3x
it7pV9bAv6JOs7TfPam7iJKw9T8JrTpqnHinQ1G7bwWb4nGKd8JhvPPOyIxPYKaJ
Ck4w+Ophd7cpz38hXPTYhi5SM+JuRATWJ3uVZ9WpDl0mz0s1uev7A8ookd/friFt
35lErYZ0ryX8Ba7dY25IdJir2nyN6f/lzNJ/qpBZRtYEXIAJAnqKceTmNJ9VdR+q
A+r91SGgxkoyEBjUtJDMsmdK9eTGixJcqI9aon5rAMGtF9ya5bVPdgSdUPHpukIP
B4GFNgptyUFgGgfmVYbJ5CBnrtcbJIMbIrOlMQAmW8kRsJyvoJ4T9eMQ6RUnwXRp
4lVVEZBeB3JWO8RbFerOtpLlVgjrl5MZ72FXdCs+0e42ZGEn1v/J/tgqTNEZqEEe
mOf4Dd2k7L3PPF7u59ZfJKrpvNRxTy6kzoMjxX74NaPAzW98EjLCnzbyHYBPt6dr
kRFQ90awpLfPn12bQiLt0GpsXBgiymFzAOwn0gT+5g1OYxRlbfllj2zVXE2ZA1Ix
9r+/CP64QLr+pZZH7G4zKO4nQaCKn4FbWgeu50wiGGu92kATRKPy3ABynOekiF+H
3rdxSpkusDUsxnG3Mo+Tb679RqWi5QhprJ+vBzhsQCspeqrQkHRTpOt/qBVOMb3A
TE7AIk4yZ3lTLd90vlrI9oC0+NiB+z2Kl80vBpFWWbG54yZg314qUEJf4zlI/xYX
UYNCxGHzpmesw7ZYOpSJrHcqdB4rVTdUqZiLjANTdCOcc+4uXmhVb0tVHZgmtAth
55oxh9bMh2bkwqoJYXlJAZcE3z54AyOkfsX2lkL3lsdAgXfnvAQRpZZKVzlg3g/c
pdjgTaJr+4Jq5X0uvOc95YG7PQV0cE+GodwlH+joa4yCAJer+0rgTKrpEDEck0sG
LhX4aP/k25isikZtZMNYXZ6Um3+tzrbBRw3brxXYCu+cHoCvwJhtKe520vOWsvnz
jPCwDJMcJUqMJdiBe9MgEDSSJHrHlKT8EEJAIYV0LKCQfp/5oUxuAXpSTSgrN+gE
67OWZWZRLkPBcbtybfPvq6NFOay8Pqb2C2pa5M0lUdUlbsoG4hJPmqHU2SkNB5U6
smYRcrhFZqev8EkfLIhG5oEa+DzY+KTZWTdV7e2t2PM3DY7VaM5DO4civ9qYW2vP
1Hwrzq1woSUoAQI4M86jC7bxZRlvgsKb+xZWrnD+kYMow9ayPKWY22+UiNCAkm7a
uqThPj/UuIEFb3WNMeLl0LuW+kMmyYHQDLiG0DK+2nkd+TaZbi008hv0Qr1C9VWc
kM6gWizv/WOD4rqLm6lQsiU3Fzd+2e2vgh5T1Elx/ySiTsWGmofi4q0JPjaV5bIc
34mashUrZAFZNc4yxYUmMeHAHv3LaUSlONrVQs7K0cD8TgKrk918GOVw8s+u/8S+
nC7MxvJBaUZtUL7LlHu2coN1TPStryoHn5jwXztDEpx0xivf1mWAlh+mMObhGglW
8CVkQF16LVu7u8er8oTnF6qFRXn47QKcWWiRAY/iu0uTLMubP5VJuTSMP67z/8Ic
/daRi3KatQOl9qqfz1ZOVc0FNuG1N17gq+w//6GnWNvvIZAub5HmhYI3R7R6+gWj
mUHZ2uP0M1rUF8ybLgpOC7QNbsAXhAHAsHSJyjRpncX6+tvj9zGJ5QOy3/7t8Xcm
Tj4GuklMEU9C/GHZHg4T+l+Q6c1kTXnIR2dj7pnfm/9wuu81M03KoIIGNWHykLHY
l1NPfhMZn4j9yjRZvo8fCH2u+oY/2LlNZvqHrAhdgvXudonR3N4JmI87xhUefGnM
Vq9uL+IqLw0EE7COmS/A6owgmbfETqpTZx8NCbPadwGw4JuI9tj5feQJNBUAmdkl
AUgiEj9shTrHntxMygYneNQe2imbB1RUgzTu/l78V7GfFbW2LdW5Xu0ScnOPC804
L+rkYyLTxxdYB7YwWR3kEMjVUt/QFHACJcLtOsLK81Znn02K8gQ3mKB0qbR1M6ZK
7zppuguGEnr/y/ZgjEwPbSK6EIG2p2tMFqkJviYY9NtZOHYMZ1gIIH1jI6OLrQhN
pf/Xp1fp6+mQV7IlYJfFNJ2dFgt9Fb/8PZW1cuHfNW/RdmzXoLZIDVEB3cC/jyaI
NVrsf0uUmHExWG1hxuWfHCbjhuNhrNh4FkdTJ0T8ZZAwREhi69JZgYgs6oZTalxc
h17EhSXXhM4L1M28vsQApjzDG8JWiyyS/0fCFzz2DYGKqOW1wwwfxwo0UtmfNtsh
M/5ob5YZlu6ZRhe5Z28hD8Soi9MBdl1c6yAeNXFDR7fuovP6hMvOR8hotveOP9IE
dv4x836ryy0En5N5eMXtOYyJHkBETklOoCuCoCXZ/bdA7iwwwkOiJEpcAmldM5Bu
b0qjWXGOm8Wrhbm6n/FpUKgKO9GA5PaCr299rkS9lelyrrtWNNNl8wm+xKJpTFLp
/Zxp7bx4yzlhQ6A7EsS4bBhh77UCxMhS36J/9CycXd6bfeALGknYWnh2TbovrNTq
V1Ets7wVj6mZ3P/CE/7sXvBQ/g5BWH49fO6mzNOEhMkNiahw2gk0WEajzjrKjw75
bRCEA0SkPaAgTal7dKhxuc7GsNoUG/455xEyL2fWs4u1yv1azL+wYsl/WSPMt771
GDOYLd1MmR9Kcw/I0ume+AzDavrOqDF0/hqqD93RYa6XM4q4s7lNJ8z4IO9OjoFv
HFEIchW8oL7t5/qnDlIAiYGF0WVtNwuPNxd0VsLoZnuwYukx+qEVcvOFxveedtCF
SdTutbrtazlQhC3hyI4EV3h4rdu+EyN/egZtvS8tfolgGgNqC6uEfFaneMygkCx9
fb5MHn8sqXsLQsvWEBhrSZvhzU3JtD3BTeZhmzYMYvpH5W7ljyTeuAvggXzTucCn
nnzqdODNmueT01Vsg/YNDs+H0m+9APaBw7zjn0Vnt5NWirVC5hrcEmmfiPle7p7d
/6JE2R9lRoT2HtjmJeh6p/RZBGjT/mOn1Dx/I5wX4ZDIOkcV3nP0qJCCgaIN5Q+2
hp5n0RIXQwnn0SmCaSy85si8k73tPmrEbB4nmb8gX1Ld/j3fFAnQMwA3Rnm2dhVd
OGirVjwXGgzt/bMKNMIU6Q4/EimkLm7PGNs0ZgqETTR40UxKmuMfIPR6p1bZ2QMZ
dZqLDzVgvuB+TZNRGn5Sawv6wAQ11W3AmcpWgr48+wZl8JqaxjG2DVNfSZzE2Knw
NQB61Pq3Y5+EoY+7kivDF00txaqvbcWtHdrFQEk9JWInzgdXLkGElKfwHY9VRUck
XV2jAPlPC0kdCQ1kdd0rojt3WcWeR9ysORebgeJ8kXpYnlJW3l5I+aKNHd3fNX2E
EYUFX5osuVwsZ736caGqXw0hM6GYk2Lu3fhZu1C2Xjc/TiBtQ46dG1juDGMB2ft8
1joQ/9Z63lT1WX1VaqXnOAZxQRzeKtrR6HZ4zioWMXyLhUmFuDs5ZRA7v5f9ISt1
2wMrQvYTS/YJTPnTgzTFZFQ6in2F3wI8YpK5OvmpUtw5VI2GuCOKWBWyEs0Wj8aU
DEB7JyNHEZFUFGJ270Et60FFoyr4DKyDJmsGhWlJJgzTiwaAmjJlKYr+NQuUkJJJ
VjvvwQemIpU+DYOHy16Ya1Rpag/A5I5rQginIIMvTzNexzoASbioDMUyqRCeJuUk
s1V+0zWehGpJBrtPYNo398BJJCHsTj1PI6+f1pttN2y5Z6I+xAwmgjAKd6B5itg+
TvWYKuyNJdubjYJ5qS1ROWkXEtmYQIkIxCy0NhMChq7U3MXZpqC7P/TqDznfbWhg
gHLYjcLHbA+0DMet5dd7q5s4zrrXcI4i1clx8zJCN2zeS4lce4YjP8gWZhmgGG2A
LihKxb2j2gLfS7OcULUWpZZeNEYKZmtGCdMzYtQJmmJUu0x+GCQRiLP1qSbJXLh5
nAzcDbsVB8rfHKXCVW88RTUO7G1OBNjdHHRyFnv21U+7HR3GxdBWpcLHT555wW4u
yqdvxE7KRu1bZ13dWjxQn+8mKlZuRf8xECE+SJTJrRt+OV3FvJe1T7B/xKya0f20
cSHQZEZnuL5vbE2ugK6OsVmugY6eNhQ4dp01wOxvULSPbyCZm3SS/IXpqvprCISW
Ayh50BIrATe+9qfqRbPu9e6X9TrXreNlgBbkBXtBGKnxu+gJtJsrKS751VIa+e+8
kwkZah20xBet7BcFxW6KY+WcBkGnYxIC7v2hSrvR0SS/6tfQ4u4XPD0I5pr4Mo+s
YnlswJTLQ07mXm8ddH5oKRLy27aSjjRA3niNR/7CArBHtuKlISI6xw6F6HbKwj9o
D7kZcjI77la2dbTLLbmRrRWZYXRC1uurFxXlsHKyQacIEEidBASbGyrSyxY6c8Vw
suVheQVHeeXo2xQDVXJKMsu4ZMMcwxeAeOBWRqvzeSLRsu934ppXs0ZdYH/zljRP
2ggmHzzeROxHNAXU0V5o05SvNURUEmwdsKIn8zoKCbNEZMo37TGSBG06uDWw7RFy
oHL1nRZRZsZYrvYDweCoc3UIF47y2jLJg2abzg7krUEy91KA+GJ7nlLZjPgqaxei
vCryM9k0KLT7j6s6SQksHmT7ssZlJVxOQ5nJBRjB0sFyfhrX1mPPAB4/PNt5ztq4
6K75jK49b/dlHHmTtj2nVkWMNLGKi+Ckg2tdG5zM2g9bAJwSeKMUtoQcvbe5hrD+
Byd/ih8BPxpC5EIhu0ppo6t6pBj4uHKHznsfu350FowSQ2D/Exr6WvcGVhs9eoK8
OrvaCVIgsOVYyJuxjHyJaeXCn4qoIA1PLcUZ/diYxj7vgQVB5ojMepq5YHVqcTDS
t2Mpm7Tobh325mPnoZotD+UrBcVsVcjtDmVfDe9tIvcewlzPWZEgto7LAuuVluHH
oLwoFIbUcqD8pqGgkkIa6yMzmbDpED+EMQH0GytGTY4YLsHJafBpRSawN7YiGhWU
H+uz2zcrgOV3J9XUJ2zJum7LJ1Wqwn9YyRbgUij2K9c4i1plCp3e+fmTSofj+497
iQYY98hT2MAuOAK6G7ed8YLxRwaO8yoDFEKBMDi3F3UMjj7n0I6Hf9WuwOBY/zOf
WY/pJdBKTYBqaOBQePsgYJxsit3zSRccdxofsypbrgy6k0JDVPOvnSIvAYeYc6jv
X00Xldot/69cWalteQR3Pzvm7Kmu2RPj+pUEbEmScxh0Se4scXRWzBLKsAkVRaRZ
PhSAyDhAYJRPNgEtr2RnIqjG/46nrz6MSRSfst/XZG2plUImKZVJzXGcncNSOgVm
9RnexZHdCYMaT1NKp4b6Q81DnoReWL9+UZur2RgBp3Mk6qK1PsflCN52JHWbfYsS
gJZoljEAZkdE5eREU6uLQyUWnAo9IaN+G2nlGiL3KFsLeRlctoJO7YIAfMyp1Tqe
FazI8RttSlb94DazC41bf1ahS2d5+7HoROGsPMH4Dugh8pyHv1WuwE/iwTOWnXtE
snrfXvjHtJo3vW8f9oMDi+gF2XG6lBwb0MWBRHWkam087tEzAtLJV+GdgGDfokI1
/1I9Nh4BbG/5pGkb6knFts/rkdE35I3L+PLtGn4QzFAQx6hJqgYjbW6GT1Xul7qt
OcT+bFgGTvlFcq3IqXMhOCI8/VJr6rG/9TZ6n+WtpQTf6rqE0D7Ck2ixlaeI32HC
ZoaE4pxHP/AJCNjOBGvdKlcmI4nZEC1kmy8gwi+omNw3HDAcsCBMqvy6tyaCDh9n
NWI7CC10BeTSrA8RhrkgxQkItewARvR3bPIyt2ulnpdaJ84H56M4KjI9OjrQVJZ9
SfLjCtspfbywcSN3E6qqY//inC8Qm4rfRm7yUSfV70Z5WlB1OOn5p4z4ZEDXQwbC
AK5MTNHlDzMWd2/IACYLeOBdPXefd9B0RnnG7/5YVy3oW5/KcTrWLTYiRAiXY2sx
Gue/gqEYbFbeMrrhLf5Xi7hnWCg06THJfFgwlyPzxDKCDItfrhtKLZ7Oksds+9J3
J1XraZGi1ab9TcExIZ7YIz147qYWACH3w/OFCaJGQAuVsd5Uhe8E5+RnbyeN9WXG
kcEUqqn3GWa1PpZ/6zS40OykCvwtfqstW00mQIJeKJCKibDz55ofgkdYiTaVaxK9
9bfULaKRAbQ56dYlACGAIpueM3GalHAmqdO/K9x9WgeCHbGysqHCeL0Mh32Qdf7T
uiySXXRXb28Whj84y+iYNcyPl5EsA05ad9TwGhY4nCBY40DcRzlOhB8LUcg8z29Y
taboLwCzpNSu6LhPk8XhE61L4qojc4PifwO0fHJ1KCvUloEEFgV6IjsGfr3UcyvG
i+UU8OdO1tbztbgUBE3zHoKYbRc+S2TpcYSaVBp1B88iCbAxs0bPTj00RQxCkE7L
PaS8Cxdtl/QVT1icWYq+3j0jx6ZuE5Yv7cmQQQ53WRExMgjUhSskYVxU1c+/punM
3bEYec7tw8rM9SWfbMxe0zb6/oMOQDbHl1oVnBtMxo/UR5RjPtu+I3PfHunTJlKP
6ATc+2vaVvJ2/IpwZIbUXnWQUs2LAHnMGnrdbBCpMFsp55CZ+inANqvCoI4HsAU0
FgChvZdX8yk4NtfSMqHrHMexIDI1ep01KNzMjp9xZRRiL9SQ5//rYtB4xUBLUclk
EFFb6qodJYINI0koze9OqMCmEPqhofXC6bztgoS2VvczfPUvuFb4ymVzdtN6mypo
B3XpmY2lzrCfmQGSttZjvsg9QY3RoIwQtFGbV5j1kQpPT3N0eicvbbf9LT+ZjKfx
0FQ9sMGvx6sPyubgtKfESqZEIrEbwqhwdb9xQApbQ4UlIE8kQcfQIXwv7FvJDupX
pXcTvfqVjn+ge7X/Hj+k6IrW3TtAI5HbpHebGayf0wFMksKlN1WLzuSMIJ7m2mYv
Sa/FKQeG20hlUz+FUVZXi9wLfFcpm/xxayMcEksMbu81oKJWpRfNbnTasQ8WaNaV
tL/TE3RGVu9U4kP9DuqTzIF2zX5zlTV9Pm+y+LK8ZTNs3qeTCnYVZfYD8FaO3JSK
irQmWxs9gMTYM617dayttrJ9cZFvc9AF9KEtpNqEHXolHC4ug2BZ1BW6sU8MV49H
u8eu6eg6SJsZi3mMPmjgmRrlRpV1Kp27xJUDQYFeT0st7Z6CjGbpMcrdJOExPPqR
cZZnoUBZqTG9SdCSp2zqBsg5pvXIi+2wGMgq79fWhRvtNiPH0kfcBeJh/yFFutbh
zp0sahXZHi9zLwZOUQQk40VP35cHnqwrENboyZbGZ+o0zng/icQSsqhuRI+NOBp2
o3kjEQeKZg051R0RwFRyZDuVdoZSQ4RI7+10f/srYSRcyudn5cpHOM5cwFKLdvFo
72UjeUeom+8Sm1r10+2Wawss6X703sEKI8Q8PxcHNCyw5FBdDVJ9cWmY46ryzEV9
2AcXITjsTCE6bR+Ig6G/UQnh0SVxAa4xj4ZQUZDCH/pppj9/qLb73EWO6BcgunRM
VnkIPTNNFuHMApczyefHdE3rzjTnQg7EZ+wc3u3bFD2lyRJS5Zllknw74rRtkKIY
CkUA6euhPXZlw3F8eKYubEAvDr9qprv0nfKrTwteqnQBnJMTshxmjpVu8aVJlHV2
vRiSRHNGcftdB5IRtK3wFt6ZLa6jd+fbNiyoy6KZ0zRrA+OUpHltWHBcmA2jgaXH
SLXFURhfKhq0WqM4YN7STyZnUCplkPQfnJPAJq0TW7vRhDHndnFcjKie1U8L0jz1
33wVn53DB1ztljjWoCMupf8RPAhkN7Nr6LSvz172JZIFIlsFPlsAh+h2Vksar8rT
tJ54of9yAocd2QMSYIuUIaOTLnp5OK2TQjngY0X588fuzzNAJVAUBJPR3/MlwB0h
JLziloJDRLrm+y6k0N3G2d9WU6uZ4CRxk+DaroqdMhyaWDBtSugzhb8wZ72krfMz
bfHTy0L3OLSWIlJR49lSSSv0GXtAePrEoixnXMIrsMuOkXB8Co+gK4x9XNjIj67e
cF8XH1txMunlqdpbCgMt3OiHkZIqAmtjfSO/ZdlevNuW9esDdoG8THty3SNWbCvO
64nV38akTeYPxo60g1xW7HO6g3xlLlkhfJ5Kh7SQrGGJdu27OUxNesDwBVGz4qpI
H/hEzxKlKN2sZSLfdjernHdx7xjDpjp6iXx8C16Xauxgycz+tufNgfqUDH0ndmr8
2vltJ/MKjgkjfY7PiIreO7KCAlPleO6x5sM6aoW7AG6/3e7DU106c5QXZrroI68+
5iWptkRxhdEAZtKsD+axaXE9mVhEHtB8jEpHG3OYDLm6khJmfATtqC2myOILzRKI
5SlP/RGraPOwla1LjbR5s3afvOyo9mLile9kOHSYjX6/QKYc7j5tEmWHDAucJA0N
ZURA+bkn/cOFd62MigjTf3270hvrNtom3vln/hr8M0vo3jyEK9ZNMlanKAxmhgk5
fzQgX4Zfgr7u2fHrqTM75KZcNYTJd2I4IT7ueCV0IAVx8RC4L8qhLgn7HLDGtfVV
KZgGaeVIVuTVKuo5C0n4QnC1Z6KJi1OEcy4mQdFA93BRGUpIOALU9j0jC44j2dYL
fRyOs3vDHKWB4OK6MdVCaaQ7Nb9Oa300gcKxVktmGppEOwGdE9Px5fTcQ/0zACc2
BAzcW6rXq964PG05tKBuYWVc8JczU9FVUjtJIU1kM7Qo+azKHVZgGg3POzwGKl2W
+h+jCeGFbyc53vEw8HFAmpXj4Qu4dat+m1fkzDWwsEmAaUOXq4r4gkTYW2gwnEbO
XbS51lqdNKI0ml4g4Taoootq4RgY2cmxLBhgvy/54Y4MWMLnO9DpvnQy7VDjz7ld
i9nBpUIsZgSmhiUEnqFtXORj8TtOCB5SU56Z2PQPxxd9/F0NjPahtoMGkVWiaNXP
fZB2WEGJLdrHwZMcHCxYQ4ZHnpZTutQi9cnebbzggkOFF3Lci7VuiHIMe10WjoxU
1BWFWrVshb50utM4i85bHMjbWHkhmKAk+IoMGXKB6Xa2otUGDR/Zabkj3LQeIEIW
PdLqiILjfLKsDYuRzWXyTPSlxZK9/wZ0l+3RBOo0dwsVlHJphZd8QS9DZC+Fu/Lg
nysBJ9yUGK5ZXW0PqHg0DRzYxl4VYifprj5utA1k4y8Qt6ePtbJoTUwvAkVBk3AC
avtTszM761GTh1R08HQnSJihH/xcaZ86TuhlRLdyNNm8YU6GhTchTxAGG9nCSblk
9MZSkKMR1rOErMbgQzFBdDJycS6N3hSfgJC07rWu6H3CcoaekEEyLyeLASWcJua5
Xp1lVqRhjsKl18Qom+fgJCxDn78V6xJKNE+g/r+omkKayjbMKXUcNziZn6Ove/ke
sH6MKtAfWRUs4+182dxJ6llGZbWzMSwC+jGNg+UROI+Kcb6czGAaXiyskRran7Sm
d+MLq72WAuocIRebvtkiSFvMPXYOTH1nBFJFTPi+G0KhG87DBGEh2/IfrSOjY+1t
ERH3WAFO6hN+GeTGkADOhxSNzJKKpRDzX8RASZAttveV1bY5jud4Q4SOLdNxlvpN
k0iWivLLCO9M105SQlb1ZH22WUfu/CeIm5nRuGXVdoH6TKUYh7rmC7pdtqOIJ6sW
VNGBzMtN1uB5HQPd6MWYu2TC/gyX4wOo9XOG3pTeVNytGsXILxy7X6FGdQm4+XgZ
rENDPp4docsPlNFZiOn62g/llx+iai5QR1bhoUeRfSkkTN2JvGeY4kFr3VZBh7BV
VvbhJy21IfKYKGLT47Serfd4J/RbMmbZDsf1qm8J3nXbra2vxKUizvCq65aM87Ru
BYPSmHXSw6bCV20b7ASOyH59hPZaHivmqt3CwV8cxJTgoAqnR3e3kyxwuHnFY8l1
faZqarcE2C7Dbef2dtETQvuHMPkoFF5da8gv6Ege+L03Xoktjcy4MgARgPKXEtDN
d8cwl0Uu2J6LLFN/mZqUsHXSSiNlSIWAH1XgSt6MB2fVlGcEKrYEXeNKFi5Ws/yO
+DBUtx8ci6HT0S532W0NZP3BgmuHw3ih8ujh5t4/zS/zlkIqdigTXyL5c0HfELRV
9xQfq14DB+LaTHyn+lFrZrg1s7d/ZFBjfhNSS5QGnnHaVOSMJHuzVdyCgGAPo97r
TtEIdcbx2BLbEQODPZdnEDlvT1saf1Ar84q5y2YtNCumTzTbIM/FE0uKaG1z65n3
vVJBRUmEla15FJaeVx/LetL5hDQ5uObLsLojnTyKqb4l1Yvr2dN/gdcjx0e9bp+h
CKdcpTrgMc5KsIxBx+xMMwuQpKgiHCJIMmGStp0skgzY0lq4RmCWQf9pcEhJorPJ
t3aPp7qEq5qqh4xCurV4isdsAY1lCW1QUtH/4EwqJtrJF6XX2Ohg2jgkYa+NgN46
lcyEONyD9/yGGgDwkfoGOxkXYLzMgTkRAWh+v9wpdCZv2AiCHa9xFAb/8J5Tdb0h
2BsBwi3/E8UfrNBuymrhBmq/SJthrGbTD07BpszIpO4vlHTPXC8DKzkllJ+MNUX9
LMRm4zD9aNAFQNDBFJHaY5LhKosmE86RcnEeJ7J0ixTAtjS0RNDew1i/macQClwA
0Q4Ng2XEqb+/OY3wyNR0j44lOzXiQtVfvvxWAVhjhxNoPzvTbzqGvKKSkz6IChAd
qCbj5L2C6M+95Ol9L7LtAe2mnjYRx50y0/Srltj0ACRtVWEhz0oaOcJG87Bd4bvZ
1GQbBj+Ua/+msThumYhK057Q0SJ++wguuhMdG999rF3LfJLYTjWF/+r71urZbHgF
rcWl39R/6ZiZeEYIOpomoXAz5Y1baJ0iw/DInEKgNprWb/QN8TlNGsU1P+YR4M/6
FVzffQbsFo+hwWCul1R34+M6HfWEZZ5waZd5fVcexElzaBXyTGluiPxUXaLYh3oq
14aTZsdgpTDEG7RMzUehtvUvVLz+w3yHgPpLn3bVlPCM1g++ePPaDp0nOaFGEzqf
v53ruIZb5WNuYsx/jVq9E6p0Xpk3dlz/BKR1iXdYzQzUpygVxC1n/z7bSn7rCH0d
T/ND8G95HuPymIheaIrVfzao2bU3gMauQU0xkR6IufUOdl8dBFMCCz/jOLuTrPw9
gOMpce/VilRVjeRR45qvSjOg95p8B8e47MT3AAELdltr1Bqw/3wdxaWk2pwF3DP3
ZCT+LbSGP8YkL5dveHhtRD/5h81FgUhLFns4hSJ2gi5qQtzsbbE2D3WeVGe9txM2
mBzzJy45knJ7f2YpCNR/2EbkuPuU10PQpxu26WUdHBXJ+MIcDoJKw42X6rmYe4TJ
yiiIKsIiAbXbbXYpF9lp6WxtBjA918CYh+9KSNUT0hZbreFaGOfo8lybk1G12r2N
yjw7CQvDhXdDbsjo6QrPFr/QMB7Lg5zkkv4JXxVybkYIa/ITU5aZNFSf9mLjubhP
rpBIXzxZJr/U8KgvhOseAWkWThdHKPMRGPmK6co1viazP4YrRS343CElnphT9d+0
jzjyv9uepZoJT2SZTE3Hczt+IeqQFnkYfZkYY6svbbxn9w7zqv9kuVi+HeS7GnRc
Ws2gz3rvGbYXs17HQYB6Gd44l1uvRDjaXHzosrw7f8GqouXrfsdFdPzDETgB8TjD
lFLcesuQplNmOdNEG/GnKzx1RY+05gh9vHdFJiuXr/gqdXJhiSuAI4DXUpic2x5S
ra/T+UTRxDHnWUUaYqIZPTkBg/om6Ekp0YIfuR8E8N5a20EtZD6oX5CaAzLUE/ye
z6+KNEYW1oDB4rJb8+lOS7WkDcdFk3ybR1gJ0X8PJ9EjFdIcaycGDeceJulDaYBu
Fsd2wh/nXq14+xaRp0r/CgomDYJ0p7VbMrHxXRzQIEtlSMv8hCA28+hTdU9jQc1a
hvIcWUKwjRhR7ddMjAsIATdMS9zckJM1RphfzMfzH4E83lnKpD8raGYwQ8kOIiNa
H//pusr98w3MVJYcMEOtQSfnlD9ZCzNgqMJ213pHhExgXP0dfsPwVdygSHSE75di
4hIBn13PB2DATqzffB0CEe4yWnad55gT2TrNKhqjgR4i/mL6dmxwzqFjSZW7zZMn
AR0N+KX/JgttQeJHYH+NrvfcwOu692e2/7JJD/CzlTkOS3751jZcvvgVuDINZaiA
vAA6XXso6FhLYqvBsh4IGiPWm7itLXP3X79ozWNnP4zSDcnmQ7mTm2AlrtU346MT
P+Ot4xmpmTcaacpC/XBfKVXeQTFY+TtDDqkTAS71B4Q/o1yISG6LiqPU5PnAOe/d
Jz8Vx0s2Txpr2lYDcIM1lUkZdoWgQ4QgvstEvqCpL3u7etnWZVp24UHKX8Bp8HCl
b6DVqdTeJx4yFvp1s7zNXfXG/tNzg8gAqLhmAbUsXAyI9zKhgG8s0ZmhCC3aL/OZ
oJ/jdF44Nil3LSRRATylKRGTykqH3IHDupF2LDG4U0KIXppIRJAD25KqcC8qD3Ae
fo0g/Zzhs71qLzOEfzKv+sZktjwckoTMLaci7pnOySyLlDRxrEZUS02FxEHjKX9r
yGv/fHjtuu38a5I7hDlcChUUSJHMDake1eayoWJh8DO7NcVB3ZxZWc2bWa/udXdj
YVrDMcdsXoTTqY4syDZMoS0/Its0sCLGJTo4Fbn01246MXG97Wl17JbqeWiZg0Dl
DCuclfMEw+/5E9fm9TiLU9yjzRx7Xkr5rHtcU9NFM7+dDqNhBz1Fe5a7gfeQ0pUm
iUEKHH8hKyLtfoR4hfSSCHKTYBJae8hCYJuO3xsjgDdbZmNSt5DQwKyqhuiouLiY
vr2mkydP/W6z9brKR5sd2zxKq+/72tH+nmtL1q2trTK4JQEXolCXQPW0T1OMiI78
fI6v7SUAShz8wny8M687+G88jAw9iRNgx17wHA3KISHP2tsZpDD/W3vrxPPRJE0N
uTPfLXxyNmGq+Ady7s8FBLsy4luGlAeJHto4APNofL2P6UL18hXf7piFSTOZIxy6
JpZWmvxaLBC2IvLZJM0zydAZu9FSjltcolF6zPSHtytVmTZz41CZUnqQyhNTYcu6
aEX8GJFTq+tNsP2025J4FftYl/PCwryQlnFSNEp2iszc0xLtbBiZ7ZSwkoZOJPk2
4w1zv+bpo9CijQY6Xa+7seGqBBkIh3ub/dOam7zoY4lol5qPrsxYPWaMNj6XnpKZ
+RDqSNIPW1myU4rFIjgxAN9QgZ+E+MXqvwhNSvNIkeX3n4BIpeuiOQEEWl8etWn/
xhr85mjuy0+NYktnmoazxYP33HEpOkLJ7v6HC6xolN2Vmdor7L4mfmkbtSqMrX2Q
WSxBkBzXIJ5oHA4byGnF0JbUlBSp0w11080o63vHMDZxDmZgD0/DoHKUR6zUSybR
g62ulnVe3T7hFrxzlw9y2nio7BO9Thx973rxZiwN37JJ2+vgMT4WNEw4mORQ4ZYc
H2QrS6uFuc8KQx+NJOIf5re1YuEaNh0xfJO7ntoQT0vc7fzsjTy6wXjxoxemQQYL
mFs+27HSDTK1/DRV8QL9+6ett4J/kHUsdnrjqIMFqMjHbEF4Sa2pGDIDz/rCRn7o
W7kdQKrVghEe9ErOFNKmxU5d31RnyH8kX/0UrvqRfasBBP8FXjGl4sYjd84eTMSp
/7YbmSLGy+17NKHTE9fNrXwnM+UGqdeM4Fr0sA8ROTgN7XT/ESWRSzU7458nxgni
O6PXNUM9v2RMR+z/9t5ZZTpXVzsz5w/AJf+2mpKGs+zsvZfFk4BPHCbb/OqenM6W
ALxcX4vKAcaQOpi+qqLIotbRLtRwNrzIOOfgBjBJfxn1ICQ6VM47VX3TPNAw5R3s
PoJ5/p0gyRHFd3J/bgfl1Q+EDpqqBtrKA8mlf/SM/s6pwGJitLhShqvuDqXRLxzq
8pLxF/bjVw4dCixoyw7dCNR50MAbULcpwVUJ4Wh97hPJlaB+uC9ouTcgC6ypqIlZ
sgPy0MJLAnRsDVHZ6S8s1adEujaDSx0U/+rMGjLNcNpwllwzzQmFQ19MKpWNdM7d
QWzLKCbMzMxL77mExJ22mbOhOD6tNOrakXD6v5O6mKX9HYTsW9AjwJ0vYUJrBDqb
GV/L3I09M4qi6Y4nAmNQSoMLrotOwQqnVZaehdKiE5ZV/GwiIAx+oXHH2wqoZ/R3
ZO6gKmCg73SW8uD0H/qKLttYvq8y70cMBdqL/DJM7Y7Z5X0Sn+L0CZgmsvjYO52N
2E++cFYWUwdd3H9mmYv9xUplFxnpASv6ZdmGIqC1Lx6If7mLxrchsYIknsGM3lFQ
bR3z9fSyScy5NMW8ypWMX6EkaaEuiB7rc+BR3rA4R/WqRfGlE2I8CD6NtHil8Zea
qjGLPLFnJUD9ZB4ouXddSMrEKpTf1CAJAQqpLI8sSHrUZKb5/9QDzHZTagKXGWRI
LJb0mhZacS0CZiwRe4/oNywfwzkdQOwjNSGWHg4E4At5JuF9sRr9R/0fd6wIbwDy
DE55aQjfcTghhzbnzutwwhZi+Lrxbe270uUgJ5pdrP+uCZ03O0cJfWOnryq2Kt88
YA2FMlaQpcAB3YuNuC96WrqziJZ1fytB4Pj2IEN7ILC6QOHCjBq4BfMW/6zEYXb/
Fi+JII1jcH/vs+qBWH8DRrLpvucZHYG6RsYUlAgRKoxXraJIF2bRFQ5vrtSZRKN5
icC6U0Z9XWBlZsgqyBX6bst1DK0H650j1urJ/SHK+Vq7AaYTfsltRwfEAHl2D8dB
uudv+YpQ3rxVb7RShQDIwfw9xz1XWQ4wEKUUehauwzGcpFZzmwLwKowIJyPFPE46
Dm4xd210jfKROgEl0g+fr3OsdlrxNCBh75kNNsy5tNceYjVtmVs0ZG1xpxH8syDZ
MiUH3J5MdccJ5g43UxLb6Hg2q9a4LwIONTESx1neCYv/1e2PCgSwgbFnnAfA5EbI
dYlHlmsRyb3u+ccMZhJItAgieNQ84v+/ntL4rd0KWTCuQFe4NErAyDERfj2mRPfK
7J+clZwZqYBQkuVCZEbXJZJMuw1rRvlyEK60zM0zTN7CWfyoWqZljhIhX3yvfLtA
7hXeNQI5sglBU+2ceAiZrONLWnJ7YGfJ+O6tYBHdxHSodvimc0tEd3SEFK18JFSR
lnGgCuLuQN2GOrDEabZleNJKb13aQHkqciGBSz2kFPVbtXI0f0heGHMdD/d3E+8t
EuRp/dG35ZkBtEq5axGTMZz4YBVycVOs/5LzQoBZydNxr+d/wIV1Pa2TgP4yUR2I
R12RpWYUwLZn2A/qwFObgDL/mNCFQE0sKPIo9772ueyXO1kSz6euOc3gTEJ8B4xx
R0ISOgWvUj36DuU4zj2+KT7prBy/sfWLVA3pNRaYTqu9o0FozbCtktkIs3ABr+rB
CsUblhJZ2MfYkG5lkY+HRiNLsT9uYYsUo888kpUW0BwpHw19M7Fxz9RSfy/W+ymv
IVzbriLxCOpWEsfLB0Iw0MbXocru7eRshBs2A+s4lLIhuxe9XFb2ml/s10M+Dsd3
4BIoZ6mgILF7INTxj7NCp2QoQ6gHmuqNJiJicFDaXTlOxBOUuS5bWHzqR0Ru0wUr
AFCu6v8d6stj7nuFv9wOfVUcoaBNVrEucMGlRF46XMy6CC4zXX4KgyEodR40Gxif
nvNrkntLMAqZQuDLXQOZ6zDv18Cdnej4KZwW5rimWshtMVO7y6e42yZMUH27Wu1+
5fWQ7zAF4AEGH6rjNYq2UVMBCPMlJgVRszg3ajWcacKTWBu55vCyMlCAiUb6Zwt5
O9G7VypNv41v9p0gYn16AP6bGiSRDkHWg4JwxxrQZNJD4YdfKRvSETVhArQNc3b2
KtutwCxhfXttTM+WtARIDgmba1fnXHhHLiIiiyUh8HkrCeIIg2pHyegXVf1kblBT
MdwDSD1alhas7eJnwgnyo2qfg6DM0yKUT8ld+mHdh4a2aTJQSUA4VL2CbmklM8uE
sjUujucqtU11BlJocKys1EuVga3QX1nS7HdoVs26n3oMYP3ysGAeDzWRPqSNDGEL
2StJttWF1hDAxVm/83VhtLRtt8KUxzx7FGYCS21FwhCK9Qg8Qh23R7prDrbEQbtK
riTwyuYpjjM/Ucu0fwTBNY+V1zItg0g0yJoNEUFSDUZMlafJ09a5RMYdenCdh1R1
Z7Nh135cbv/qSMZBznBKjlXX9DwMoGBC6WRXWYgUkHn2hiXFpHM2W9vNYbcB0k6t
SGJOXMaw8pT4LxfYUGC0W4I1IPT/Cpsq43EhyBRIDhr+WMj40w8jUeUVRqioYD/Z
Q7Fv4YmqYeSdlhivEeGv/43Tf/pvBztQv9K/4QU7BJSQG4HUhfgzhNGtlI+xfXtF
HIjFXGGLYBr1jySZp1/+5Rabd0FV66izMVbT5ds3Mn4S2NldJJ8/9aWKqo+u0kLy
DsF/7RbPArA+Tox2/BtmfKrbtEk9JS+6k5vIjUgJHqeglzwRaAG4VGbHnexXq3Cr
UPbnU26BSxUhe/Iw+HsEQokkrFb7t7vKNcSYTPIrYKFPgKOoMUtMbNYrxQGuJF9i
2z+gZHcrv59j/HqT9dyh2f6AhtBvP8ZrUIFuBGRUDQlzkcumEALGSQPe7Xc+7xqJ
SbXcSXyrsQCgsTJ8zpmmJxgeNgxJi2or11glYOuI+rL26Miw7f38JMjGezWAw8bw
CkYex/MZVukwtr0fS3KKsdwzgWq2mIeXsYMTNERXK30P/UviBppotQtfTCBU0ZOi
B3H50P3IUTLwINiFKi4jo0BsSnZi/wYRABQkm8eiWFuPIukI1AEpDAJGfD9IcG72
kvOT3osHJi4n10teLcLXFRXPqftFXAZFtn/kxp/IDRvgA46zDDS6O04XRR9jj5la
e5oQEIl16S9Q2Wcw6G/eUDZKB11pSjTo+TxHJUrKABGT70oLizaCAjMBVkU85yKL
j+ZoiEfVP4Az5mQfKvP40+38d4MLQ0Q9+059V+bQE3GleSEzDjs24YCaB0UjrqAJ
GLR0hK7xdm3xj9FyO0X4RZhTwkP5XDLNPK9N8mqa7pR3XIcXJGNoCWsH7d3i2WL2
PEZPDRAHybxaTFfTczAyJftK97C88CGDQPn4b8gmUrPGftugxUvMlwaHpEAtLtOy
XOIqax+bR9/WuxVfm/iR9aYqHfvGqYoAP5ZqD9fd+zmKC5QzTGr7XQkau/GMfvu4
EOXAf8/XvME/W6v9y/2P8QxVWenAujZCJ17ML6S3v4PXeGOrrEtzbZg7YAeeexgI
VMj7P2PgLVNJi7j8W7MXtz+AliQMxp7nOJkrp8j+SzwyhnV12BfQAPtmp6gdvvIt
0nuA31nAVG4RoTqy05JbjDnHEBzYD2xmQzAeP21HTgfFLS5R8gOdFs+dUaIDgej4
ZcouxktxjVc8rR4VkLiOzUA6iv4WN0VbSATDZq2BDTaMdejtDFPNQcr6e7Si7g+9
MVV69lzv26YLoeOJgl8GmFC4I8hStEykQpRG8HxTqPtwy7FAbRWMoCXxKRn3gZb/
CVmi1gqya0iWOjvW5HtFRfplleR6WxxvvGJX7pZP5TsQFS473W3syPWBs4iLDdPH
8T5ieq8ah8oJaCRCC+QTvOS/OHfqc2WKIdH5/RVe5V9xq8EgHMoAYcD8rKMVGq+U
up2oKU+6tFpqAGG+tzyLIrNsmeQ6xT4h8ZQS6jcjzVEqEDyTbfntraliJkQCkRSz
eU3i3qbesByKPcJbz2vm1vcnWAYcE2m34Uyg8glmHiYg6JFrUPrUDGMi3Mber0A3
LsOqdGReC03VpLBPWRxz3pXwXwlLEIeqg+4jJ/Glbgicv/C/NIBWvMknliUh/H+W
vsc7zoLOlxt8Om32hgLdPNjWi2sSmH921i/wpjNIxoUugwOehpYNZZpA8gB+GBIK
Al877f34xG8LphbifOY0xR/jrcXXIbyQvMHMWeiGvd/OvvTU794TUsPtKOf0IMpw
fZ78N8QNHE8Zp4MnPX0bdkDrV36n6nxRl4NByCkFta6hsVJKIgKpp8GCeCPtXgFZ
Hk+37gvzh9YuufNvYPaOtS3fQiTVDOIHDWOV0btQQHApZNoV50BkxPgvGkR03cWg
Ulpxd6bIfu86Mt13AcF3QP4XocReVxUSd1gO+oWX3lVs/i59B0f6z7V10Husdh3q
z5VuLnU9/0pynRLXjy4YBlw01DQSFxko1+SwDjYXdPFn9h8iNwfD/p0H2ree2dqr
GIPU01DwVuNsXhkxQU18ivrfWn/PhxBFAw1+TZupwrjDj7Srl7kLVW+5quckqk7e
DMEmVAHWyts2nNQbLRlidYHPetQ/xtxpJOSrVwC6CraSj1R8vu3N033gf8k+Cgj4
ulzwJwmaySkA7QCfIijT2/dXtDXRXiub4Zf2pCFSiv1qaf+TxaPppKyH7ERwGHaj
4x17Xp3BYsxtxf5YWX2BaDGwsxHsASUvWtc+ebXtkEVx5NMzr1YrL0vWFSQgwdt1
BM/YQwH7D7hbtFXjhhkIvhYlPVj2xAMal7drcPZ2sSF5PDy10PauqjWPchcKs8KN
Ajt6XMo3mrl7UlZazs6pVOCDv17HAp9Di8yZyUXIexKIxjm8z44B2eiNtKXPJevW
k4SmiwNwVT7Y3RA4rmfjOB57X8OmIxRv0YhaJ1NQOsxk4KYuzUrq/R5IsD2TnHvq
dpq9KrDAFmEgaPyJ50640QjM4UXeOIxIx8ccd7zbCMb7OmxNMoEfDXopTqCKJ+9l
9Q3fkk+mRIC0B5gxJC66iE1MWTW9ctnaMilJAJJKCzLpm7KroC/VmJ3iV3/tH12/
0nVA73ZzA5II7t6MK1sYtkSgZG4xqqNSJxGeC/N6bP80kU6KCOXF+np+9mliXjAn
yMSBNnWip8VV67xMDjDzEnfEBelNljMQGcQ5PtfKalH/OzyOBj6CXa3Xd+PI3qzF
0BSuOYqjWpN6203JMVN7Sll9Aapj/+uit0fsHvqtV4NJZj6z8PE8OYtWOS09Vgum
72UMxonJgDMDf3H8OemtKqFHrOQhy68JLZHgN8geS87c4qgBFfWT/rLeOX1mMQWk
fCT2CZD/5ikJiogmWsXC8p1NEKwBCaDqQcCVTyIIGpBUMGEeUVPehBNsGtQdciWP
Np/sF112xU8gkgEdkSY18ndUw+2L15uleh8R/TtvNVFmd1BTLaLQ+CBLHJtJ93QA
yUUw9qaaY66G1Lt1G7oYmnYHKi3vq+W7fFv69ENL7sl25/cRuOrsRRfw5HuCQ2Dr
GnAMv+7MZuDvPilTGqKfV2FZpK591JhcYmnKLjpj/1FK3wOP7KkUZlMHnbprusvb
NBK+gf/ogUPB/MtRDUzb0pMY4Ccv0Y6+y1I4jciUmIcZU6X+jMsBaKhxIRMC5Uxd
oQ3UzQC/nIVpCbchypEVmbcIlixDVHufsP//ebzYmaPP8ZsFPCFzgkrc931mewAE
DEYK36How8dDezD8g5WNyYgnsiC6H77peaXyZBxDt4KLW23nUXw1Kb+H2wXZfmop
U0aXjeAM+fKY/fyTpmjaWrprbr/q7eNIhypgW5WCEsKeaBuQulgrzFNJ/s3Na0Su
GMFRVqEDEKw0UdsNfTM1cLsbTuI8YZHU/8AnIuhy1kep84m6zvRr0sJtHAXEE4yL
rcHtBmOXg9HmhDmyb91rl/ZxAdIP2HpkL689X0PlvVnMBDtxyoouJiTPqWJNl0uZ
fjOA2Da44IoYgrVhfsW/QAySbO0NY53FpWitHuVtIXsOWQ5ebQAEPDPJC5HUZIGs
K3Qssq6LJCr9/NWxh5vY5v4A0Lr2mjdgVx+LcRIskvgxyTXejT3mciLVGNRCJJYm
r+J4ksSuMQCK7sVVFRtS/aT+D+OfkdQUJVoOoDq0XZs/WVwkU4TxiqYbmubpjrU4
rNQErRtOrLproLUcTzT+hO1IfM6OHYXNASY+NvPdLLFQ6VTCt8I7E8LBlzNUUkhj
Va9cYQ51QifH74aoO92Z0taZnlUbERJRV9RJETZNwvaoFxHmCLNQ8A70YUT4kibk
zn1KXlFQ8nqMJyCaEmTNHHBkAqq6TJl/rVCyXKTmxFDvqejik3nKPUGRSwuVonGy
ALRudiy+p/7fjYv+4Feaw0r9c5jEvBnc/gcubvtAIqjA7D4gETAYePq8gEu7bNjE
vX+L5hKkXSRQH6zv+zRd44FIzVdKcBEDj6e9Ob174/FtatkDbEDGDVfhuIC1VD6w
y2AVxaJbXczM/OofKZ7BJSlhYO6S9Tfyqv6FIiFOioIUGHvG5TwpUAAlxDDNIlP7
Vm22WZQ/WUxHfGEYXWgvFFJZcR77gnBwG2Hm4+vRLG2DwmX0vPJkOeZqdvC+Ry4W
gBKvD0qNC4r4DscoAY0UlRYR0uoFQrO6TT/L69Y6x5Y5zmEDLVm4zeP7q+qreiXy
S2+7B4wuviGXy23xTNBzfFFPxi+8b+UN9OWnDdRaTwG/KBWKzUbNDzJ4TW2fksQt
E/jvJbV6xjWd7EjJn1r/8QjznPATuiLCkk/3NvqqLcRR3azERGbMZ2hpuHQGLLCD
aVayg06uU03gy8MkViy+nnmg5UgmIHDhWWz0X8aQGA1tB9AV6Q9oKXOv4HSXYc0T
y4o4n3yljs0XslZ4TPLtjNQlwDu1SStsNHWL4MD3FBB12fzY5j8i2sJF1190ZFnr
Ciaifr76w05flFvM/eaIxCpOjo3Lrc+Ha4O7JgloLkF2CWd/nqRAc+b799JiNj9T
IIGe1Je/vnl889ObeR/R2ZI/+MK4YOOzOfrU2zqkgnpB8S3AJbreiwLHu2dB/MJr
9VYEhaQcY6nFUmA7IVFmT8a9+sFZr3FsfbaKLQDC0q0QkNhOHPyeoN7eVYC2oZ9Z
z/p58NAzYW8fdUP0md8aCQJJc7neYajhcIWbO1kfDnyjG0T6s254IgQtX98NJ3bM
Lhp/koO7boUW9UaCihaZT6Dw575rwQ7I+Mjh9AEmeLg2a32UJWNEwQPNw/9qXqpJ
sgmLy8CJmdoVZE9+HDR7ykXskSGfv1B31sb6HSav3VywvbCN0+veUwnH0ZM3ZsPP
XYb5LCqa1bXWlEW8ZtF96rlQNgLZYcBjidl51EvSUJHZ/VQLVV6K6ntcXZnPPbi+
r6j5JQWpeIExvjaz7A2msytzIFXvof7xeGz4yg+KP52Hl2ZaA0SLQzU5+mpUkZOc
MkKeUa661GNgOxTncB9+6ErZEFjb9ShjxMMuOEpYthiFKFymGh/SMrVAOKhXUbhz
d34BmahGDR7J23VBEY3my2KfgC1NYz65b2R167rHxHG1T/JwCPMEFQ7+AEVsEpjN
3ey1/knkAS5Tt86zXWzYot51lchKeAH2TrV8olbT/BaPRTnFZ3+3APbHEAyQHv6x
yMZ/bKaEx/+vPWY+M78xLKqgYfMg7XSiZDX6FcjJTd76ehJhv0twaGjOK/9ML6q4
cjExAJ3z6RNL12Wo4+xk94eo2umz4CjjT5wCs1SLwvXaXisVqEv2nqIaYVyiJ0wa
KG4wqZ/BQ7qHN3oNr8m+E1xRZXKLkBdiM4f+KqU6NGhJrzDk4oq28lEbL8YURGfV
Q+DCp5GQEAfZCb+WhQM1hf8ss3yMw8K4bzVtgpyThdss7c8LAf6AmXIe/Mx484xB
kARYZ2nXSvMxcHXwqjWDU1Q//CP3h0oPJsEQG6BSaatu8mAyXBRMu8rBU++5lE3j
UGFJx4oYIgDR5bv2XzabuqdwsZtByp8DzQ1ZZxf5X3GM7bUP5O8VRL+nLsC0bdlC
bDS5+lLDwtxTb76jSfZFzlToQfwYB8OjsqJJ1XyrnzY1QMFnNwu0P9Qz0753WA9q
/4N08uUFQ+5+qKMQFnPS8lowiEVsRLsSSVl2DkWKJCUcONFNct07fW7qzIQlYm3L
XSONZmO97jx92NYOf+aCi9sv3/gDF+FENM1c+0Z3qv1D3fwF7UeuRduW+uDDPTEN
/SgF1y9H2sax4gK8TToc0n80Z/yshXT4LZSpmtCFGF3IQEaHW9JYBn47X8YWdOyG
W46N2YqJMwzzeHjDzYyNPrcsjFwSuHHuHLMu0s+ehGkl5NzlYsm4QQX+RYvpgMKL
UjWBmToF8Qp3eJoY/qfudJjOCwalpK2HHOaawNHaH1/mMSPJT8wZ8fS9zkJJhTxT
3SP2YZbvkwidBeP4cKOXxHKlQRU1wlFVIoU7rkwwh6bUr1ngHpKqTJb0pNYNmaU8
6gkFDu05bLr6jDNDU6etX7oDnBX/6CoypsFF39KGtoUO1qejar3CaKJgILDz65mH
CEC9zfdQ6Hi0eKxP3IW4tgpaITZzeLIa0nFwoFe7e/GY1yi6QfY/HFCT7YBMCYlv
JSAuzdPMVhZXykGLhi09E2DdLH+B3ubqWVcu6pkiRL2d4Uum7JrH6+q93sOK/yXY
dtld6eG4kNfLWiEAJgvl6UqkrgvpHLC22PNCnVMOwocQkVSOjVFd48xYDgpx86AV
X84nCof0KeGSijy+PcbI/eiGVTYui56GmZYWrPrx/ql/jUQYhzaTld2xNIp91e5N
aJlhNOAaRe4C4biTFfu8A16WtcpF8s53FKmnzFzHsnE+OiH9ovcoYASuk+EK9xKP
zZ1YCFyS38s9AL3zf/716/eUEITte38aJ1kSv8fcN2vkgM4SuvKQmdQ07C1OZxL2
vVVNYLF3snCXgsnssv0Zd0ddGHPG5t1mtc+7J93hmFk9v0PIunHzMBgwzxfKqWfu
AcG+9FxYlg2WazqTubeozWGXf6XHpa3L99N8A270PevKY0bHk/Z7xH1gclkDo6Gt
jcbXTQ6jOJ9RG7iDmsbWiciXoLI+DEVfLrBka49ow2Mfyjxc8SGyN70UXv+KxBMd
CdS7Ss1gwiQEkn0eP7Z9xV/BHQLeFs25digE4+9jC8SIyI0cY56cldt2HVAHV4RQ
aNU4RZOS21Ui5HW7/TCZvkoRiR4egWKuflVOC9ZBnO21nB+ap3v+ybPtJopACxPI
elM5ZIX7bFyLOUkGVBOWaDVACguk394nGoQG45L0uyoIzCxo5D556+zf8issHXQT
JthzSsbgKgiykdrESPziTmVnIVM+zXYHgdB5z/LAu42ru51xXKeCbTVn0oQOVf8w
w82qPOcTsORu8w/MTIiiUXhBuhZuMRqFBpP3ducbpnmtSQbEZTVI1V68uTr6bOYs
CA9VCuRRRPxR31j5ktBbApPvVjQFWTnggaBX/ZqaZA76NPURnYXzBhlVUPSkyGbG
m7+SQ3ttv2sbm/S2GnjZ+rNq9nPJ8hOBp26iuE2fErk3TCp4qGAMsUeqkcdWtSLP
xFM1vNwCLXXdfFESISuW+tETgMJaELJ5BbCHh367GXQRG2hlVKEXKfC07ztYP/O0
1cJXZcFt4uiKH4j3bqlbp5OVJns1mzUTAyUBchP6Dwg+0IEWCio76UewIMNzY19A
HgNswzXsfwBr1ag6Yotz2uGHIQjn3BBPavQcdNoR3ePP/Lby4LjSdeU+Zj726g0n
PmKfAgs9NueKaPmZnbC7cWI3fSxgqok6uWzVnwm20qTPQxh+Ct5aVFVtltDJQCnq
4cHOYqY0X1GZZOruuJknGDKnl1OdvNjQj9V/E7jRAHeDqsINVaLFOrVt4swSavYU
UqnKqn56VamaKisb/7LkSo/YMWuNVuS2kS0Tzk+KK1i3kByICWi0k+8zuXw7cjYw
yyeSnzNErPIqKrrGaBX2++XXFGRfjvPslpphXKpgGjcT23ljh3F0llWrTDewvh2S
wFGqtNWM3uKXry1rzM6JOPjLIa6ZG2IgPZ7k5k2W/OygAtD+HV2jfH5bubMcygpL
v/3cyazD8H3UrOC9YV16P3GSKXNQeAeBMcSfcmUrZjEGQgonJTO1/Ckw4DNESGT5
s9pO+0m8hxt8EuenVFDvOJenD8a8szQ/5Zn6Bk/iKrnk7Dwo04/xyozGI/88hjfG
1zP10tU8x7Oq553ylC3TQV3xNe3z000iOGPvIFvx2nuTfa9wa1/JH+Kd/iRi4Myy
aAsm4vneGjoq/xQieyEptPAY5LWghVMHHfcOQ3oWoF+Kl4atfZtKg1DfjFuLq2CL
ez1DhDJdExNkKvylIkUyQ39ZPbjiZPkLag2NcxW21qCY3odQNAeQTR4eboYbKX0r
uJveywiWW63ch7pVpboY5egu3lRSkR+yTQGnMlaIr6B3lWoq/zu0We5+eaX4KB/W
rlbiWlLoZFk9fXGTNfiiyfNGEakrbSwCluBKe9T8EOtrZMkAl/ZphmikAM7KJL9h
DNsMIPSrcz0BAHAnJqsl5FZINXMjw2CThdCuzCcY7jECEgUeGreioV6cb19xYKR3
DsXwTwGxZSrV5e2bk3r9Du4lrsckH394N3jLLgYmxDCRAtClZAg2g8zmHOrJSl57
QgYnM61XYMRX6vABLNrxMvrgGj1t/4l3hcFv0D/8JbHJf/HQaxjnjNMmX2rA+I+S
17pr+qfk7HiUZ1Vyykxecm7TJZQmDOf96BQLgf1XDhuEjF4GcB9cfFXodqBmANyI
Ja02aRKbzMI2wu0A/kKELSjvOoS7z728SpONgbChog2gGh+3thISnfo+rlZKb9i5
sWKlsG+PgFOcB8c0ylIUSvKP7OCesZy4sH7X1bipL70qKz/bOnZ6ZZVwykuYGAi/
n19tUREhkzAv1Dv6gXXMyz0qSuqkTioh4RCokfCOwpvTExc+tQOzrR0nn3HzVCKm
Q/3iFBxQ933cXeiZnX0sREEFToNY/4ma2ZDzGWAdk6U7BLqUY/S5qXi4YDTFbuWZ
jJFQyip6ZNO6S5AZ6DC+amFrhuE0PZWcQAOzvdf9//AzUO7WJpytF6m0cYzn2C2G
JYWK6AAD8h2+vEXKKDiW95TUzn9/Nf9MptSJICc8Jga96a2nLAfz8jhcCgyPhnsi
Nj5G04npqNIZxDDzlxJyo+Nv3I5g1bErigZHBAhotTkzqoonraacKOvmlSTevTQ7
Zb68VeY5DyX1cpk4Rk50F5YrbT0A+GbRSQD1tNskhbS5Zxjc83ssJ5SykA20K69B
N+4ODVSfWbPPLPapeBwWSrR6KDZHJYyg6JkRiJlOfv1H8gia1yP8qUhRosYfOUTu
MQC0/XDosH5fXCo3lroN21ledAQOzdmUrKxllh3ZShIHzxSP58Sj3a+oeJefIbqo
cJVCalk+a76/jEKRVagR+U6liTklFg/RaLxx+DPM7XKUEgX/e1KdXOAD2Qp6Oc78
Sk9OI/I91n3eozVuKdu/n4rzS2hC2P2FxeecvDFZn1OR3Z+od3sO7GfX4BE+Wng8
OxoI0IrycoEglqAqR1kQck9W9EQrrH8jQLws2IpBmClBbnQtNQH2+dKnBfUTeXVN
zlkCfxnXtlPnlB4U1C/KrQz8gnWJWl/j4JKPIpNFR8dgq9vEsxmfv8IBEYiPEGPs
7Sig5awMycn6QDWV/6+x5sdZBnyVeO4IQD6Otcn4N5TyKDygQRTjtf+WVlWdd3Ie
nbOc1xipquFDxC0Rgr5/E16JPd7z6X4jjuccS4UyQ90F47gTUqTwykYKvZ9sQ7zM
fw1ThZyRQeugAL3j6uTd2o+ugb0ZFXcanO/7DwprmccbM4rBV8HzhmudF1FRiQsh
pYE6O1notR2cOVYVQYpetJgLgw6Ou2YjSj6ujmjRACtWsY2quDtRV3RAPiVAm6kQ
0amyCTI4+oAtqEy3nG0B/f7TOCiQkTMJieZYAMCzru6XIRWoU1PhDpOcMNVV2csj
0+ZOkDXkQ6euZrDqh9pf0HZOtsiCsNMwjv7wiZEe2qovZ/vGRJNqINNmSM3ZeNog
ISHdsuVOo2GFML6b1HnsF+99VlaCEWlhaHKyBHa4TE6IRKqfbp2pPFVAczTwhLaD
3tLyi8ukMn8KGCwzqxMMDKXhu5W90++wHoLJ/SsGM/tl8+y4fGnrkpNcXN+OiBtl
ybt1HHCB2ufhfKUMSyvgg05JS0LTg0ccEo/df8n37OOUouatdDP87I1T8BdLqMym
g3I6hoYb26THQS19CINeyJlSp3u2OaLuEexFkw+qHMX4+T8G35F1eDHlU+FYUepy
DxrbeEDEbLVRTZKX850f1XRBn+xt+GO7O7AKzu+DQz/9pcBFkzDrAhchW0y7n30Q
c983sX9bgc1IHVScbHUmsWfVeHqgyZunrh8QLcPFCiNGRCGyMb+wyIm1CBErxEx9
E+GTjZw0QL5OBLjDiQzhcN/J160WGt+IslGaXFT+Ipe9UowqbtOgeN5hUtNKAqz6
gAK2JULrPuQsjzQysry2p02t/TlHVfyzxAhfZOez6d231xG7Zxh2pHzwmsEGRj6q
q2MIGaCdUYgCEvuFVT3Scq6DiVUWUFWASKt6Jkf0MVrNFyu566gJSbk5P5bMOyLQ
d1a3qJgE+2C9hgFKVJOJ/g0dLO33hr8YSk1fdKuW11j/CiwKRN9S3dpFukjWwV2N
iyhvUo83wIuU4kKyMm9kU2qN+1WhZkW+kLvGxnXTyQP1I9k6o2mk9S8wnGP2nXeC
qKDLBzmTJdz2E5kqZzXZ9u915vEZVxkvs6qWxzqzIWU4ole/LjdMZuCLgDqB+gp9
QGYafhGQiiLLsBJjaQuvRSejxeGSMjufv1l+Hzb34+ADcgc1j4mg6Ez52Aklt/Bj
4Olh1bGH2Lz49ugzgqx523G6PjrvRE6cldMJzMQLgpiYjikzy2xzL8gxrs+/2SVn
Ert6RvHsryzxn2C2ocNcQSB29oC2D+dkfEOTYTDQfDa86769WQYYdKAZJq2VjdlE
59jZsSM/uPailD+1pbRq3cmciozTo1bowBJZXBkooDNCdKVYBHRtnTUWgYp/2Q3G
p306p3PNMCbg0+36ZePn8ga8RMlyFVe7snhnwqIeXx551dY02PPG2BaoxXezsLXj
zfjR4UVclEXHpireOqDjePGtqmRBt0PrDVIo7NKJurzKhSlL3L2NzyzTVczvANzN
8bT6KkqyASe/RviIueytgqpdqLAFSLL9n/ExktGmhi9MC3/9x0L5Kbx6UYqeRMXs
8ivCStSS5bPvDMpiMtNX2RfmsJBtNpvFn7Tpa61s7StJ4BaWKNOEHGnXix0UVb+n
tsWYb1s/LbPXzE7LUgUtdFdpQWbSFSUskEsX5Ge/9ScbJjwOIhwi6q2IJBXgGoJS
s2WorvSUWeWOybXuWROU4Gz8i8tYBlencTFgXEKo8l9wUnrAlhjpKBWdGqipT+Z+
KP6u6ZwRcrY+ViTL2XYPwT5R/NOazRjvdovFgJF3w70mK6ChGSW4noghJuJEPWBF
h7JVzj73sE18JjDuZxTOCbr8kF8350uc4qIKWamif7txSyEn07Zipl9y4B9s+7lr
GxUS05jpjE0sel29yvNhmVJSOCNnJ96RG9L8Cve/XPzD0/Evw3yrOPV1JQIi2ZlZ
qJwjD/sMIRIpDTon+iq5B6M/Dy6Tyk9Z4eALJ7txPCtWUwdhM3RSVLOa1KkgA4/8
hLe+nipfRbRZzaP5A1XMsOotdUqQh/LB7CzGFmL0zLGaQF2IQ5PRGB4eqQAgW2I9
4y4kv1gB66kyIMl9c4Cn+i5W2dGPbR9cfK+gSBBBfjeaJwW3bo5sLaeoLiKTMZ/7
O6W3KItVW2E21fmBFmSxYU15RgF31ha9Vy7l0IQsWnBOlGQXW5oRBWX6oYUhXERw
f1Jav5cSe77QPVR1/rMWfYzJCesGYKRDAEIEmhZ2+HQOTebg2qfUgvLPNMZjRtGz
07zcpY2nulFxXKBmZW8L2PSpL1dUmE7DeO04WWdLHQNHoaBfJkEjO136IU2IzTlU
wuRnhSV731B1MWVf1oqskXRY6RE9dsCijy+3C/O6h0nRZ0aOwsnYX24YeZEdvPZn
JmcEaoa5mNacA9KKyN863QvdibpKIOiMvgI8QX1bvAXAkGmLoii2GT9u5btk9BYx
54wlmcUY3LIPr7GlV9s7Wszqwc53d07Pu3tlcQTeukjyThPL9/urThpyXRPKDvvP
r32s8FtxmKpFKabNh0+NZmAM6gaaMcyzhrQ7kdAOXzg4NeAu4DpsooecMgyYekm1
SXlICOSXu6Vx6L3ldZnU9/fFu5yBZqGhziQViTauzanXpPdZIFeXpEtC8d/Gbd90
XVkppCKNskPk6eDMCYve8DFxKXUl1lQfRgPUagl2fx84ygRX4Ywcn5PsATLcwbog
CJ5W0+0n9vsXCd8JAtw95cykkR067ixV865U2Ae4VlqHZdpSb9n0ZkFsxMr473ui
1YHs/8hpHcUbV43P/SjBwF+NfyM2yWBYVTaiN/aP+gnrnL2YPZOAq+ylGplDTwHV
Z/x7Kz7Y3rI8RrdTtNVrZ5Pd7N+zE3T0cs+3atod3zW82co68gTvoEnyYjlJA/yV
zxyxdjy4stiXHYSh+Y3wNSb3vEfZLKpwguBbYzhm6icYoqVbiu2RYNOSPOjzQ2XM
z5kOFR/vKo6R6xiQmtMgwmAV/d0bgh60UOE2qg07L+QjPaKUphgfUaztseLjTS78
o0yUUsJTYIMgMdUyI9t59zy0B0kI1YgnYu4DMOgtgd0QlXIX72Vj9k8FHd5NxRy9
NwtNfYfzbmvfNCE5KVVHQq6NzUsBbcII1A4dTL/yZFAJXT9u2kA7lMXjyswNOYGV
1PE6RHJWZR3Los4XbV0vinK2L1U60sbyYqYEhxgrmfsw8I7HwyqBbQA1LSJNuoZi
BBDp9olalmgiR0XtDwlhFyLRul8YYU8OqW18ciDxGYBwohjrhJB+rV4u0rceEq98
Ahmcfx8CN87xfUfl9UP5gZA6sRTm7k5HuNq/zxkXGNk5MsCC/F1xbcavGKdgG3sB
LxP8vx1TINRq9NFwySwYBgMdocnGgxTj/qGHKoZNxn5WhxcOtmdOMXsIOfl4lwEC
GHOtH2dpVNSJeHW45fAGRwPCVeqEBzLB1PBgO4C/ptAZKiQzQEZIC/veDRUZjYe2
z5/5gLtblPIcis3CCrrjvBF7LsaCDMWxp4MpH/T9XwER0lg4Om8MbXAAWoYqFLj7
n22Zr6R8BtaWCV+lqQoK5/4EJQtvHn7sHuYUPPTgGmq8k+QOGhlRDowTjRvCoKn0
hRIiIXdlZY7DpvnIf05O1d6rR8Mw/TaR0D/Tlmj43OfW6l++0ql5BZGcyE8WyJOZ
O6he5pIjN3PZ7QJYx3Q831SvRsFrFbDwkmBGvM3uKO6NV7rafjTw19X5wVgrqU83
H7iG33AwMt/gd8bsxc+l5enCI8+Il2DBL+D9I8rjfqo2CDEu153Sk2IthfkA3WWV
1CKXEB+EO87Pae41qGhVaQ6mGmEEpTx9TVEJdeWlHbGcY1USXkYfVoxYKN3KRPAD
Ekx86/vCIjpIA06+l8zn3Pw/MOTNzl5pjvO/uO66FOYBFIQCggp/4ziSJwuvnvH4
r6hwso3lEyORz15cs7frdz0h8FX9qcwJW2Y+xcE8yRuYKv51sjJTdV4UYD0JXT86
CdB4ND8xNrNMULjPEAdvFoWBgZv59g0oLBIfVp/ySCdV2wG28CbLOz4EOpyHkBzl
/vVn0b6ez3XBXD3RCYh0+kqoMAoFpLgVBL3rYcFKwfEJA2JKAhBbReDq9XoIfDe8
46sD+UaeLhX0pBg4IKN+6fTc6cYgsytYQBuM8GSOpwrDJ1ob/47/oP62IcSRdSqY
Gs+YUpIqADsQz9goih5NHJWrYDIR+sgXkwhCEyYCXrUnAvopX0iCPw58C7r4xHAx
YeDAcj3YCzUyXb14WSFgjsY5V0k1gflOUEQogJFGjUvYxbmnsZ4v9cZytSilMq45
QiPHr7L6ucb32UmIEYW/SXmHtosL6ZDTxZpsWPbLmcXQ5BbI2MSZLp6aDz1BHw6u
8XS9K9tRTRonjH6zPGpLf55nXPjPIWTHuVDFzWGYXzcFJHLjwLT5ToJIp2H02zsG
kQfcRMgcYInWT5Nw6jKgViQPQcltRlSyIp/PmqqVyTOkURgHXSqPRE9GDLKrgjSc
Qm8CStxzPDz9z3kab2L8NmjHClpkxIlFT0kJF/p+2Qj3pd7m2+Njx7Qf6VSiBtSG
aX11AUjeMMZz8BwbKuc6ZYHj6qy7rSrB7ZRTHO0nwDbVZscFRt2Hbm7BHdPk1OSV
csLPh7472aLldXhm3Jrh0J+VnnZ71OkMB/dXemvy5GksBKUfjS8n3ukeZDw+1QZz
9wv3L9JrMpVo3pBLnQ+9xcafXcJ12U/JrX0M9Bjhtc8bMbFyfu1fnjxqupW314BB
3Ob5aOazz/iPki5yr1shiqs/NsOSaLdSV9D/FubTM6enly2NQxKV/PqGHzErz1t8
9oiHVmspY5b9Lu7KLiQHkqv/frDpu4Z4eWTbST3aIB/LrIEUJESRGU5guFd+YSI9
5/+l71j1qUY/pf6kFvXqLVjGkMC+oMLRYpi0S7Sfbd1rdwpzNHuHrRvv/F/PAOx9
Mu+l4C/lhZzpJ/bTehPJqXa6z2JvM8MBDJlu2uRMfi6boeY7fi1YFzJXBIyps/Rf
We33XT9CV9yC//69kAkUV0s8tJZte0xC52xVYD5PZ3XUKDEwrcaDHhRwPk/KfHcF
ZiWVawWubUzOezbpYo8L/A+rQp9hLtktol7o9pNdRS5yIsBMEXz8KlQkX9tLjGQs
zNgvbQm26Hd+GDASUpvtffK4jtb0d5C3gejkOFJizCR+s9siDhPJ338O5nQwGuPI
QcJmFPD8CyINMV/ALOtAmiOZuoRp3EYBzMfZDZNEXXUPt65psvgmkzsSciVTscgn
XLpXZ9/vUe1JxVWRVBp9e7It+SIhsyFV7HXEr/p7WH/l00ahkMPwGZie6p7HXORj
4lZ1FMrtL403u3RWoJS69rKk+kjNk/At2HbmFN6KHNtF+Ko/Q29vgDCKxSAWLTPC
GQSBNL1sQAUDBd2W67copMlmPtESVrTua2sVdeAe46W9Di3cpbrCkT2jYjus35Aa
yZPqDnqa4adMudqHknD3Q2kNCHUNsxvZ6k4tjdAgb7uvozu+9BGdNdiYtuWzl4gD
Xc2W0EgLAv57kyS7pUEQ3EqzOlSY+D2B0UlByd55knkncu+bCTsCqEwNOESOgMiR
pF8r/36n2bz87ZAKl9Mt0ELCC1O5YWuhpRpCadzLivyxwN2lIcpjBXVIrxK9fS1g
jYlGDnv6rWNBbihD9fszoVATW+mPAaIC8sd6GCoS609SXrulWvSJMbMQ+q9l/jwQ
dy/jOyXZd4sg7vzfoKqggdA77DsfEf0WbLMEnw3LMiqrp/dxZZ9H9HYWv+1OJH2e
38sF91hsfxuLQmTCpMZ1ntl1zsSXqJl5oKy5oVF7qJ9g4gOjY8GzPPcfmNbnAK+C
CE4WjNSfzmIOIRYiMrMqBkiiivXplVhVJrxzBbPscDqAq3V7sPfHcBWjwi8yLaQP
kwJiakN9hIJ6tghfly8wKj95KUuOy0xIVsstvUHwKekWGnluRkrUk9b7mLgbZSaN
GBYOfAikUXOBWTfI2dRM34fcr+tbrdOBikydUEWDK+V2qOBHrc6KwXoKqwiWipnl
CGtIFlAyKel1o14oukWtnW/LWywfeXytJ2N50bKbNMSraPCov7Mgr4wveLL+I+XP
utuft6rWKHoTgcDxAfPj65pjjYfX+d7SzTBiuLjNcs6IRO9bHo10elKObyf5v7a3
pl2TeeU+zizKzVz7STF45jajRYNMfVX/03C0BtrT1LcZymnEPxrKxeHT3JytMFnS
OdDQDtpTvI1plAt9veotbM2jqVcakQ9qm4v5TIKfDheeA0hgXwsE+Hon1koi994w
4I1O8kf7gk3Y2Hv/YNsxP5xNFndY6m0GO0tQbYhdySR32ITKb8P+XJmj7BNwtgDn
tsFUZkitQlVo1P2eVoMa+rMCbHE5BJOskHW/3XaUPsOXFSmvdTIezVUDxh/gAAID
WZ+X1dr/zRVTTsoqk2Y2GblSne9X45ZP4Uw/jWPGpIeZeF89xJnlFIWfod/lbm/U
gvbCBqfcNvxVyPaGa8d5iqI+fDJ9SfauSrHT52HoxurGqTU46uumlnVw/O78zi+r
9vT2b0X6sowjN5FUXPscDEBn8EJz9LX3tiiLEt8MN2kJ+cjP7uyb4xUb2t7KcZls
QoQq1SyrPZsfBkChyyZ7y35jSDSLQ+ljiALkR2Nq0ltFrQnFxEj37ozEhblYburT
yxmKIQ8wFuE8mvuh8C2SVZ3MmwpoDYIRyHockN2rGiYywoMgGJmhLlpbqjFS955m
LFUAM6v3P4pl8GJkaxxzmH8AgRpHHtJTnTLRpF/ip9Ryi1/Sg3rZBPxA9BLoIxdj
hUorTdoYLwY2agv1G3AcfnYwyHDW/WxcBJRGwT55cr6bUZJ/w9jmcPaFaZJYmIeM
1qDhqQqJlY7GGidSQeH6CLQx/KiprKleE9O4UN2l717NnFIbIWGgcsj5iAM7J4Hg
8AstTG55IF5TN3GV3dVtoWsviN9y04NJ0Aw52p2FnXy2zn+2Tb1bLX+Noqmwgg+x
yMxXrVKSDQuyIgBpY7hh62Yp5UOxtu3TZzyZSj5FJ7OPrn+38bxLnHuk3uFl4VND
dEVRTE0BeJLFhTZKyUo6fv/iOzhf/CJLmpsSTYOR/LBexxgMpRSnoH0cFD+asnqK
L8aUqPIM88xIipCy9qYTMVZjKrrMenkmvxwonuOn/DYiSUQoGioKCmOPSgM7lcBA
v3p6ioAFzN1MdMvnZsnHwg4S/bfxL6L3655zdR4eKiro2H2qZM7tMgcOAJDFVnfv
ogIo5a6EnsvH4LBgFVkGLKud/V2Jk00KW9/Tgrra/SEvGqz8VL9SCUDEkB5J4Onj
ctKK5EYrtowDcjX8xkj2dc7FA3aRY8MvLYoGS2y2IYvInAYLlhF+jPfUyCZOgBpA
OTaGOaQkdv83WywSkZhfHW4VvjPIdAQ1WeXHqb9TF2Q11nLV9Pf6aiaMvKKsXCW/
1N6dTXcHU+tAFHgqWmZ74H2PUVccWpqzj0Fp6e7xG8aMan9quAoNTyy6U7MUpNmq
AKWHMNzL4cZyUYkp/PEFSayIIicHp20+MuMdr5HcaDrs8FGhUd/KOe3BaQO9NCY1
12BwK1w4c/1dzCsY0NLSD5rkYYFloP+Saa6Rgb8XX3/C3TLSrZiXGN/rTW8djZek
k4yTtKDko/nduk/cVsXUnFIha3VewjAg/IAOMGCj0o2u06vPV5WHP5iV9DMS9E3Q
CI/i6QI2JXUbAkfNT4/AR9y3tXL9r7fPUw628ZNsDCRmzwLgYS/rf6jhSf6tf32V
I9iD7TWiiBHEYbS5q3W1knFVw3yvZkydUsoZ+wCZGnRQ0Qq/v3nUuzGi5oO8T8OV
GSdWBPTWhOx7IQRx+oFBQlGXTxvSfFLJvxYji40YGf/Rn47rzbjEm5NckIwYyOpx
Alpr6ptZysuPl52j+6lJU1IBEBtfCTEh4UL7ILLSYfzb3YpO8y+j8PsCbMJPVt4F
mQoXfTk8+717wL4Xn2L6k86AyWLEZxYH5KzDwEc0sKEm/4jfllUXwCsJbVKMKuEm
zSAq9JAkAtMzeHOsVIz3pQNLpkI4veFamoElIv6dYGt5Yz1Boa45GlkMkyzPwloy
Gb8ozH0qYJey6stH6wjTVeVqLKC+SN2zHwTkhfzhhUs1ob/W3WQuRjCzSoJ7n8l8
bTuSfIn37Mvcsa+SEHmhLtKHqmn9LaGY/O1Zi9TFP8pw/4qBsEsjWtl/PrLkTowJ
mMzUGqdZlGbcaf+4q8mXeqfmRYMg9NodKi0sWaUyg+Fqv++dftUgnIVQZvpKCKYT
ONNp2Q27bEGrxtQHhI8R/a8HwmXZ16ZPMF7XQVT8qUjHXznJIQRNwEP51+jT7CXh
6qXKHPO0CNfvSBfUjLG09xi7mSk7d3yZ4OCQa6DMGhzB0eWIu/hcI9DpFDutLOaM
chQ3zSiHf04Bg0uqPXA+5ZSZBjeIxyfwoj3UY+GX5vY9sCDiMGIQ+5pZ7Reh4kxW
SES+N26kMuWPipJrV42QZP3FFt0rOXLuYAprRgfbWJ0yoG2mR9gukkXa8/Gnn6wY
B8AQr1mo3Vm+CkoQrsiEmTyIlxFFyUpUDE9d8wIucM/xdNmvVnitd42HcoRU/lmt
7q4wI0t6eEOn764WKnskwE3ZQSNf2Qszu9tzGxkPVCaKKjYMcZ6KXh9wGQ1frYvm
L45QmLzgaSiDsJp/KFA1avDbZKdIYmJQ95VKkAmICtzPp1Xh6olZb3d5632UNJhI
GBgnnNKY6VJrrSDf4ojLDjs2B2A/dABw9a9PtqCrsmU4bE+GZz3AQqBWKNwjn3LH
AEysCttyEX3b5LXh/tRljGB+eb0mskOLPgsNoK6P4bHRNCMqTM9b8TLKK9C/MaVH
Ykv7CWzrKYf55+WCDfozzspUYQMmYX+hheWXJz7TWub6uCLz4pMcvHWzSMo44MnN
LG8vdjF44J5X1SYUi5ntN+MNEl33fq4FsogOmZFdb6Z1NU2ctF3NQkSXewjAVc2z
OF3Qt+b//7VNSS4AXQ2Go6gWxweFK6JReHuzDbEsGUhfKXEXV5Q3pJii4xX9OR9c
ICLRvd8EHQGIEEbZAqau6OyrsVJNiqDf6l1p6Z2zxcZk8RXCMVcq3OEdsCoTPfwT
oQWUyF7FJEpBMuCViieQD/wb4w4tCm9eWoASxR2lBWbzpChEUI3/2oMSm8RlUfKe
wAwZ+bFvhJlUOz+O7SuXZzOg/YaJJXPj3BXy7BqBoNFFpzNNQnpqbiZaz4n4WsS2
2gsGe6/h+e+xGCYoSTR0w4BV31Aq9GpGC9/up8MA7IStukvuj+xZPLHeNEYQYlTk
vnIRO8L1jCj+An63xM9IIgnfWIhUcC6GwzekO9Oyy1La1f9TqNTDphPr+cgdGOMs
wcDTcfIOSXZUxB7qVLA1+9+pj/Ts1frml1c0Bf82JmfxMBK0FGlFasnw4uujAGfc
60N72SYJCuChdVWmh8X3ggsdEtqDiS6iAaDHAgVBjf5cl7cHLvha7J9WCNN9opEr
My/qvzukz6YWMOx2GAkG+EtA0Zf5QRkJUdCpnvamB6N1tKJEBjAMALucj5Lv3nzo
h/lg7YzhV+x8LNFV0dV6fWR3g1v/17h5IgxOPdo7uDl2JDBpf9P3blJttTmpxL0P
mRpkrCzJeUHqnQqYfBiXcFgTx1qncY9GHsFRRhFqpnpCLXHreFxbFX6+weO58NsN
XpYr3Rfs3isquwZdemZXWQdzAshTnsKL7PpbtXE2EUaEnJL1vj9LiFYmjdML1Sue
S/kMjb4ujCOKA4XjE/2laPJq7y+tsmf8fjdpFfaDj2gfj7Dx/U5ozJFGDnqeV9W4
D1D9OdhmPeJiCyK5t7CXHbKqJJn7ALuj+zJdIFSRd7XVizrMlNP6OEKVF+e8OtBR
/PDOmT2HSzJgrHUGcTsmbyzjQusiGvcJy8LpPP6r+yVt/QVGhg/KsfSqGZAkuQIx
xHM+U5wlEQvOhzcoS1ngKkkJoRbAjwBso90H84o2kAN1oiP2SBItx2NsiPu18v3M
tfidlPdbuYULjljG7qwh2gALjxgiGqSJ4txlHEz/KxR+eTJjF+1yxYdVswZBjlY+
dzl1vXV8cMBkIl2oaxkXYSZYJjDRovRwxU6BHGaMdy9eNsPRE8lrg9PaQMGWCK6Q
6IqlT+ll0vjJIlUdtR1xsWWjdMFdu40o2o6XnjoY48lng3vrVNrnXimICrW7IbhF
tktKWcnZjNYqNCSR5QOTu+6zSU3r6intbo2JJ2n6ean2laFQaZvF1YN3FxbyINnC
PPWY6NvG9o5ukuObjt2ciIFo4xs6Za7miQWusbiho9yyIry4mSuOhAl/O3brR1sK
yjeZxjy+Lz/PDuroKwPwO5RoUL1iHfBsoDYOYGBGaSzFnZ7as0YS2pvRZsO48R6J
0WFRuWJONB3TRhhbAHQusV2uySuLppyO0Dsn820tbREebt7O1nRUL2pbEqdk0THp
8iK3/ZvJApM62M9L6CKRzjLw0FabWjEZQAw8gDjzYbFhet4viOZc99dYHaahJLrG
O6tjvA83Sdm9TZe0a/AwpmcVRVBSRb4Hv74dbTAP6zV+4gPYAc2n/qTF2bTCKNab
hO0Wig48A9Uel23Dt+MMbzGQfq7CFhpcoDCMn4X93KgyCRnVzLWJqzdfRkz5rvCX
07BcpwiKCMBQiNjEakbHsQrOJDqfdLHD1IOyiU9lxCTrhFEyPFw7/8ivVlufZZ1H
jRxHfRvvpBzo/syj4EMp7pIL3RZuOoyBfUisA9h3NiwwxQ3mwQqzsMukgzYz5prA
vl5QupRzl/FPwtR3fnkV6URO6cE5MXrZJEo9PGYZNk4D+WEzlmAH6yn5N7v3c2KX
24U4RMgMdn34FhhCoF8qFxahHAGrzOhdQAI2gGPMYKaHkcsP9ZbdvyWZZU2PRtxd
wkq9RvxQjnKy3E5LxK7zwyWrm8JHtkoTdz8ugZhwA6cLJ01zXd5asp8LFug2Y8tH
sdJ3ujiZ+HVFPo5sI5CweJfYq03z2mB8mh6SRFQTQngD9cQI8Z2XJbmQOaLoDguG
CDwm70o27c4HkngW0VNM8K8UEjBktDGAzunLjpeg6V+hqV4MRNXesBpR4vtupCLx
X1EgKm6wBQNLU+Js+MYE2HFQDH4UQ3g08jvF5L/on+10t8Cm5V5YkdPHIdztWjkn
O4pTyKSKtwvMRjKi3KJg5AxeG/00x/NFZL8JMyPQ6cdWeite7CEWc79E4aSvGnYf
mIZPmqr48v2wCrEPfmsh8mxiGYrqy0o5HbPDzfgUCvdURKkA5ztSrP8uqqkgQS/f
DQcj2wObBiUidY5+X5uFhBL3Qgj3LFQUzmOUSBaMrf9dD7omytY3O8TP5LR4GGZF
aRfxDe/cjyFaOaYmUQGEUJwUKhL5bGKimshaLlMpSAtqNmzE8veU+NX7X5dDSnif
VuQ497j6d4oD0JUN3ISYWfU9Rc+YHMHRbpLdzq1WnM7rPglQt3bCQnnUDo/q60Cl
seCGEiqfoSvdlOnAErcfUb1DRvg67aC4jOi9dKpdLJ/RhwWbp8BJLpJ9iGK9kWfk
T/ng9QRIz+8FNCAI5MBmlbU0YSRxEK+H7gvuAfac0XS20M6MvptbPpqHncXk6khi
rMwyZ4sujizYKg6T6rXOYluqQggCpbpmwnUbAg/YnorBEi/27NGU85l8ThpEMAGp
QGSPOSXS81ZZjLVKEL47rJ7f+ToKLciUIv9dMrdoPEgk5iSSJwL/+KGKpIncPijU
YRw+w0Aoyw+CFOMkwWBJIUf77o0Ob8cwUpqLztfIV87DoYFIi8RbEAbAw9wlZgkD
vJj4x1cFAWjW9Idb9pATxwqX/LNGoLbhJBtJyvWpHh3m3pOsn7v847daQRf4WR6V
tcVG+pn3PHff7+lKaalaQZ1TXUpKtGVZSMV8N0c7099DuegDuAo2xDdWSRieh1hn
BPdtPDjouqpa/bWbicZrfDU6/7e12/J3nPDWXPUqMG7LT8DdI8hlV8bF2IgNVnl9
H+aRgNioshaKEsXhYwDGXzXneTLQZTh5oTpJU/VQsHiBtMBOFPTSmYAUyUbF9Te/
fXdiG+w6dWTcpbbu6BCkCN21dEbwJn62Ngl6cSC/su6taGVq+Ufo3CP44rA0aLQy
7i8v5aq1VvUywGefVq6G1KRaXCSoaCVl2hPxoT+vgNiMmkAHkPu1/ZsGA5e/r6ny
jkSG+CHzUpgSEnxUS9ocI1d0umBd6d/TTEOgUIU7GxCVHP0YGMYZtB7NXYIcNHSZ
qlWyO82gy2DYbUYFYvDZs8Kys4a/U+UDlohH3C0qY/xJvaTS3sGfJd7g6406Bzea
qSBH0A6OTLEwqQeU1PsIy8eQubr/F2XhCh20YEc90Q5oCT4jvt1TcAkEmlRWkcfA
/utJlzWBfJO5pt0ZKfGYOjYCi/7UXzq0Xx5W9ShCrf6twmyeKv5hlpyqVKALixqd
ArIHjbf2oNs0whTZwCiWlTd+P2cyWUkXJVu4Bx9k7jv51oi3qX8CCULTnadYmJqt
0cJjB+wmuEnNyF2u3wShsiifYOUtz+4Fctt9pJKB7Z2BJaPkH6tgT86Iqz5Rhu2L
7qoGL26VVWUkC9JjviesW0LNTlsdzHcprb9+ItPtHDVytum1c3rwfrH5tciFGENe
m6QrH2ydhBh6219EArJoK9n0ql0UFaMs5DY41PVI/vXIoV/m1ghIctm1c/EVrqZO
bfVqjnjDOr3m8DgLsOKf6ik1YwbAYFF5+IFfmAQcdOpUGqT7PvjSAxXqqO0iLTRh
nNvAjdNoR6Y51C1/m7vk3PVDRE4dRFtkhqvOBOa4CxSHiFR6YTkEWA0TCTlOySML
gpm08Gfu/Mw5WD9jOzHKxZ3q5lrO8s+owWwP8q/7V8J+I6008+nyY6wseJOQvNvb
Z2zSG0WIEEZbtfgcbWAvxV5M7XyS6KgIpbBVUbAIeLbK+PUQbnL570MvtzorO7+b
HKIC4xgYPpypkrjWw9JW26GU5HWrnMDkgoMo1zGb9dwnAyF9U0cyRjRRPbssSprg
tEEA5n6a8wXjPoeHJ+LR7fgL5GgE/iPXFxGErQIdffcUf3QpwzCyRSUNj8LN8uFh
GGO5D9qNVkzXtLoyo13q5rHxEvCmgo/94F6XPGVvL/ZKfocEyFejBoR0EBBlN7/U
Br4vXcGeQBn1KwIjLWfEiyK5cTkCZIYrP0Y4oTZ61QIaL4bu95G+4chvgjBu/Rwl
MCBN6i/Y/jv8TkbeZ/99a6SBZH0Q2tL6QpdJ5klM70kcYEWqtjip8pCneAmhRVwY
U5CMO1XaF9xsUz0KoyKb+VP4Swga4c+OME/DPEwjj6qtfPc0diXV1rMw2Hr+u8rw
KEriwXLNT/mMzI/W1BvFG/wAFLDfItjgNTpM2sLGNNbwUSZ4epLjH47nJUSnH77N
q1bjyCv6y/0n1lAKNDI0MHVRkaV5E7qmU3v50MBh4z9qlI/zMcVIoMc7wxu1vOS6
XB9vK6qTHKBwMlQjT4s1y6Nc5Cv4vRwm5uBouKEiWz9XXT+v/v2IJDgrai0STx9q
vQciFv+bkyMaB0h2bcf40lNdyAWNSPWYqlqSRNNqHs/MI1CXjJlxObJL8uDBuGRw
OKarIIjcdKxRoFV7bWpMcZfVFpm6/iq4UcSTcMLdcBRGcLva+r2hS+KtCIFvCPGg
4/IgGXLARC/39MC0tPzeAZixt1nhNoKnWjFhnZwnaTEqFi06lrpUXEC3oVhuASj+
6436Ueo31ZoP6TseveGAyFPlrX6OVb9T+KKdh01kt3Gmbw++L3LehQHbgj6QgHZy
2xXWcICD3vOmvVyXsBBWlNpZ42BbrqICNF5JJkvVbuYL/4F7mT4rfgLsUq+oPuhG
Dk9S0qKb9MP+xFRIR8I2XPqk3w4VzOWgZZtoopMa03t+5BL3eW8BW2wENIWmX6BN
BVF6HCPeLuXgDsJVWZy227856bBRwwo+5GCUb309KwH4BZEWfMN1GcAh/COX1sg9
GhI9DP3XnHbC/oEgvN9AlrjlZ4E0QpN+Q+qZuoBUc/Pk3G25Y44QPkbnPkXXVqOh
Xa5hiijbmN+WgL4JyVvpCz0RGhl/3RMxa2GKhjRtRtURIHFj6PNm72Oqowwo/xlo
Wol+5PxIQ3petJl2TKOrvon/dyqitQdKjlPKJbEsgJHSYZwDxN6WZoAMiST/gSyL
5sjtlEsOezcGZhwoXfa3UdPt9av8Hc731PG3+041RordL+P59dqvW2zPLN9VGvFy
jMPj7IBTyH87zgRaDnnM6l4Nq25KbB2P/KMZWsuco2foXHwFHIkD4irx0lE1cH1t
2PM1h6i1OUQSZVqV6oISl9HJNu5+PpR792E+DUkMG5ajTRGV5w0Blx/TwwyRxZJv
kJKbvbwNE0gD/xVNOwBD2vD94uDXlmyZSk8y5TX6Ho+X5ZNn2Twhl7eztuT9KsnZ
NCRaM5LsY/U1IdLoFq6bkLNTCynU0c92EgNUeCD72xBjIhii86g3dGYCjPVZO2No
GQXkTae7xTW2EYGjPlymUujn2DsgwmdeOZUKNa2Ik+b6VbPR7wmowr0WmWLP2M5J
u9vBxNCIA9qg3H7xg0ViL7KHbd/f4qAF11Rx/MSzYgPfyIjesWxUfLzXz0Af6Y6O
qGUh7+oE9Y+Hf35GIIhB0MUYkF+xKqapUORqdKkK8511LmbNyQ9P2w2RSxki3Sco
TjrJP5waS2yOoJtarH5a3JTqk6dwKaYj5y+mGyw4qPhEFlRg2+tABJXCqQ3RS7kP
th405zPn1nB+cQ82qoEzZ8UYeIb/XwKPwJ06Fd2rRRNhZ2dl/pm1lW0M/Fl2ppcD
Xdcr3Cj4SCbe1QOdSvx1CfyVOGtvV1O7G0BI2iUJcZD2ex4FrkV8uHFj2slN5vy9
fLhuc71fPMOhYgUPElLMYl+xqQlEH+T5SBOM0wiHS/Z8uPyyG5Y+bkSgxQIlIeXU
1VEH6zZdqYDNGVOJvweU0v0adX/kAmkMK6KWm2JufnDLXXO1BGS6sHp7uBORZ8iD
xUHDFEeXhyirBT0XI8in2X1QWb/p0xtxK/USKxUeypvYwpFGMcPm+LExmMJGNizF
IIY6KTzMksrwjgAVVX7N18CTpin10pnpp3Ia3mJU+ozlt1RaiUZYo6DpWbYz0uvQ
gvTkVJMxuz/OezlqljtTZYOOYglvzhSDSsRfjnBtBvvy/nV7KS3nE+aisN3x0KXe
vfK5RxHk8OqP0/acm5fcLLGdcc3h7jjPGOcQVvfVisP4W3h+I3e8HinC9VO66vkL
+k0ztIZcNI8Rn5iJWKUHNxaon/3lK/UAsMO604HNN1gBi59rSr+mgjXK8xUff3Jq
570o6vQ5lX6LwbkeFlnrhTla/PTHgJvkoJKmZzW9+V0ZPr31nHQOM15l8r9ke3RB
msJqpg+RCrStBou08e8db72uFHGDFj0ztMB7FjRDpZ8bJAMLC+I0v0gfeZC56r0p
rx32e8tQ8DbuOrXEIpF2PQfdxAI3rXGgjRP90W+As31ojj4hJtn+A238xx8i5oLr
AwHBqshezVv4q+PdeRKxp1lI+Vy3CvcJZKShE8+iL89jDUq+5gJeRi3oylfQIJtR
BSn5Vmh5pyot7BirMSN9eZr411V45sMX9eKQTHTSczUy6m7lnHQoAFKJoY3VX0yv
E509Hxt0esSGaQ4rky+6tVYd9H2lB73ojPEHDGB6lu505MHdZGDQ7tMi71MHV4wq
0kauYErXoJ/9sDe8PITlGQT5ZquWBw6YRq/ujYqj3DyT0I93vJkCg4sMPdVE9JF9
Z9F29/levkpfVIE9Y5Uiv0ND2fhDhbzKnwF0/70zYUrrZNpHI1Zbn+wFkILziXec
UlAUxDFzEGC88m3hhaMoP+l+VY/Q72wf2hQTXozyjX28CCXsK7Ut6KPgPixKT9I9
tF/GAj4aZYjGvu6zbDkKfYx4nThxwbrkWZV10i0wDG8P2bhjI5ub5tXJbqdjyDZ1
j57qWt5JrIAS/jwssHjMigH9lQrjsap0XHyp3kNlWn3p2IM+WMPrMpGbcoCg5dNF
Q9fn2n9d6/xQLv5b6+kljwPhcxGDECGUO2Dto9jNNJfe4kOU3MzZqcnXUVYPS2Th
05i04Vu3ff7F+yYL9Zq8YAD1s7EFL7pIS0AwGjPmvin1aTzTbjQ7cgFXcPRm171P
VQKKUIdJIzTOrYMWuvcT7+O7wR4/4taZTLQ3Kwmov0p3UC2/8StLdT1j8CUsfUzk
RIS3DrC8zYheWKBheyfRSO29bnedoI4vGUStMCSZ6h7vOKN8hTNaZRGW+Gle/0SV
AARpwbhusNOTauQIVxdrQpVAE+EEanjZIGMyyhuJS8ha3IQFT70lZP8EtdbMjOQk
UANbXl5YJ+KoE1etHuST4m6wqErqFMv7ONOeYKlM6QZ3l/GjBmd2pHdqGbq2BmYx
27AyZ4IVELto5v7pplUUt7/IMVBhGg5Xi4sirNPkt17GDKYMfz/AO3//VZEPYHPg
BjwEvDVut8Md++2OOzj/QCGG6nK9gOweSY0kzlejzXOcjm9vuoXbP1Yyl89/Yq8g
hvwT1fGgUMWqy7At3MUOby/okRBtALQvcVeQKM20QIxRIK0I5Uc65+Epwi9sFW8i
iQ5Mo+Yjdm5sIum4nprHE7fg5WrWiAMBJI2Slc+p7ir09YKU922uIECtKr01145p
wNicMawyAiwxaaCfL/phl1L15+GmzH+SYb2sR88zda2LCBrLcUwWR2+SDqP9+ukX
nuQxcypgckFeaDNtHzTg+FLktJc7x8btbxgS8LfmGabZeqZNc/bOYFkt4o6vyP+M
cYXCXsm+dAuv7Eg7IpXPk43EpFJ/7Y1GXnxWZ/YLTxmsbp+76qPTlv2BoG0jxzAd
E6pmpq7vuDplYNBOKMbsAU4hvO0TRLObQik0zmkkHPupAYlGDVjX7CEFKCa56tUE
slK6Kh4Za6+y1k01LgZG1D4X4HvReETJm7LK2r+jRz1WtQMpSb++SBuBtH55Mm2+
DnDFJNJ+kxRKl7ULd9NO4Cj6PSiEdgWL0wxRcoUN8gPTin3Ko2zvDdh8Fpm8U5N9
10JsNqSw/lzqd/4RKa/zL6wxqy2dvL1henTuchdRiR+c8PcZE2DkbR1cyt2NWF8r
leBbz8pDeaNqUZkELYucf9F4GNZMsK6/biFSjwCsrIZd0eZehQXvsMOmTs1mzri5
1pV8ZcwMTZdM5wF7TFCKDW1fIS0zJmx9QfLc2ACXvArbrfNdVVxpXNjSApzqu62U
dt3TrS1BKln1IkOQYvT5HHDeqmnbve8my/ayksA/0gkJpcd3EU50Iorzb8LMiBUi
xFfL5kaLRlxG78USjLMQifKOdKIDkahB0ov1Z2F8iaL+sIuUymtLl8eS1HJgbSLe
JOWyHwvNLyxjV6KMBkMVc1ARdpg31cPC9gKAUR/BsMuBPWyBcHxCSNJLFhaXkSJb
Z5uRxbQQEn/huaDjMv9IeV4TQ4VAXWT9KMM1NM+yEsE29P5Re3Lu1HvOG8Mhm8gJ
SW2zfVTLtIaUuBLh6bhjAQKaHojHQHTZJ00SJBMT9fBoUEE5yAQ6x++iFoJSdasV
YAxuog+f4ZMKPc4R/fHAURnEMU1NyVjSHhvFQwSCwY+nHvViROOi/sLPyVLla33o
Li2YtkljOg4nIlZ3n7+aSeYqJuG6KTMWcD8kki9W1l9Rz5T+5iTp5iLTEIKUCpoq
mXpF30B4WJJXs40vFCQk4p803VTzwQIBwg8lsBuqbfksGyo62XAFugI+MhUgvYDd
Ik9GTSv5Y7NeNaaMfHIqoNS7eGvmFHZ//ekfE3jmGc3YZe2y/U38uNgy79WNKqO4
lEf6fxI/JO2u2XXO8vIQy0RE/SxSIqnvlLYDfong3cSK7vreibBbyT+jiYKK5dR+
hNSzMAyOHdOLgFYFoNDqi98hd1Xpgwz6tB9T+o8F+TbE3p2SvxCWjXH/xSHiCX1j
DjBVUkKcJamrq71OMUVoX6mMgPsaIJb5U26zRrKPA0v4na0hJLow5nG/BMawXRyh
s7QW0N/9qegLFzuLBISb5lDqlmNtD8z2pDb7TgoWHg2VIx44Vgkfx4QquW5StEsk
tmRIEm8vDTL7+Vw1qu32AsqXmtSiywgycwGJtOJPPV5WFJwxxEhMvVhbiGmho+HK
UGkDU+Z/uGhu9oOrBHuHWFz2oXp3OMPVJDXZ6nmTkBpEiH8LzwnZ4cL2znLfr3S3
S79McK/sSMaAtk6LhdZa1eBGXAsUxbGrPRK/uIfGRgSzUum1qJ0XlJ+6Wg5siJXu
DeWVkshWjux1RbY14dQDD1ZkYRXPAIum/681lsXZrX2p06ZXRdJTaz5tZqF3QgpZ
KlLjnrnraLXusl+9rryfU75zd3paXsuMby9i68fYuTEmoL76P79qJ92RAKi5tGJS
CH+a1C7g+yR2iM6IxrPPFKTDpIzHj38nAFTlSpsQAN/VQY3IRPF5UgmIISRCx7eN
HBOLckomVrWtaYRBN7zYED+gsfXZPqpsj9w5CW/+XdlX3K3IZIoF4JajE7VvPAor
RhPaKKAUD7ZPgBFPWB84cVxs5kGFxLO/s3g73uUi9VEYBjvNBmjdNwKmZzscmAC4
ineyhrCXM8E6LQSxtmWMhyavfHbxLCQ/wn+9yuX4lQmX2siwWB8dSDEE98NaAJUT
VusuTTv7NzBau0e7vZ2tR5ghIYk3iKWRVo81z1cfVDrtsiKuM2zvarapDtEoNOn4
QJaiA/XwTF5Mn2CbgOk7BpT7MfNB0cOwDP50Kvv0YwKBS59ut5DiVYV8cvfIrqRN
lWXHfTFeBDKGTq/g4fACRnP0qwDarvXaxhJ+ePEtVyt8FBNvJzevTsLnLSyYI6tY
kMo3RRsRYWBZn6SFOfPe+H+Oyx5TpjPiZG32JRC4PPg0lw4E3vlsl4mXtpE3tCiV
9gIV3LPWVZqnJr6JgAUgTOXFV+7RtplBoBv/GP7qDmVMXrBpLRgyV2EfqQcokWwO
b2/UOl65KKJ+2YHXxbq/j3NieTEGFlSAC01wR6M6l9uI+hW3f+2iJUYW9tAAf4eS
/cF6slcV+UF60hvtmPTzF6rRqfiYgImJRAeoe8UzN6e4BFWBLQQG1IfNL6NEl8aR
PklvzkXr0qGGQr6Ssz4JsCvFccEfWfTrzDbfpEI5YImDCotDzKZgaL5UNjyQsYR6
70UHhEai8b8rkvqDg5xITemXpFapdBlLUNjKD7Hm48ngGczwhn61f0C7yjaKlNmT
YRhosqPuJBGLr2pLuEQzCO51IzzLojv+7o0y+2+sFYjA9tVxjUPjkKbONRTD6tdX
3FI2yA+YydSxJ7qckttM5JT7StXNBbSuwWOdusCtGQQ3d1PLWv5QhdoWcZ1rQlgP
WAhyqjT3fOBC1nfBGy5QOihbLgt1P8GzIDS4UNQQe7PeIUDJP/zCK3tPxkm8pLA8
b/a2PZbNi5MlM4kymX0dGKPUky4O9SfWRNsckdR3iomq1fbfrPH7bH6Ca/MhBuEh
j8mNVBUGKPB8zfcZTBKhN/eK0NTsxzQwsKckfc3g8glmXIxT7H+VOtZajQ44MKce
sJUdWKUk05POBhAaz3XvTe8zeybNPzc1+mV+b9WMpX2FdoqCUgQJioP9jZtN5CrT
xtvwxXS/0P5dYoLfq7dc//cUn1Q7MfgWSD/QuqZ3LSuAWnBUSr4vhJn+3o6bFcXO
bzLoXAsQOV15G5ZKtVw/q+onfpsUsdggMBXmas/SQpXk4L2onvYASyWxL3NGA1ZS
I0Gqw7DDG/CabapqlwldCCsgU4ki2IsXfddl0+rvNWjlJIwrGkQavbMWY8WMD/PG
SopFzNDlbgNJzP5Pv8lEg7Uo/6by+pIbpG2MxO7lhI1w68EpVRevgdkghrLjzJNl
JQrl35B+mcwm3h+fbR9LgvW+DhimHXY2yGfNyWBVKMPJ+1u47AQjDzmGg6zK00iS
aO4S6SdB7qoFmjV8HwMnzXWkn8qORip1t6RQieajgofxS49n9eBilw3x5GWooF65
AxRjaGMBraHQNnJnoAFjHIZsNrz+QddGsiOff+UGOOjTyvFQVuzMRRMZR3P3cC3k
qvWoJV3fAyIaitQQ5FsCm5ALF/Xa2yo5wxvjuES+d42Yb81drCaocUOJi4Vqp3QS
KsUP4mDIyQ/BYRSzRVBM3PsznghxxsOkrvBj7GDICU5ymVvfgNnSzFEwj5kc3Hm4
lOTPnQJMxF95zfuJ3GvjsbukoFc74YDOVa+Cj+LVGTnLEHhsLQ2Fcguzpb63H9e/
ufdlxLmUWfp1H2ZxHciwU1hBFqexJsb+JofLVx4E/MMhe9H5morMXZpep2wuYnZR
lR+2+p4d/JZd1w0+CFkDcU+JehxSgpiw95SsdYSxETh3QKQJajoacVSnBVTZaMF3
FEeiWaGh3mcXAENDj1BgmJKgCLEIgpGPBxCw/YR+ythjI0bVNwhiI/q5xxL6xuNt
9PaVt5qIfAlNWqITMy0LUUz934FxT5vU2bE1XM28FeKcMmVhpnw2kIOIqF8kbYIP
zGeIoShOmogBrzD4nw3xi73JnTXJ9AJ/TQJE45nWkEfQFifCEuxePsFzxD6exJ2E
S+hkwryHJFwbmNvvUKnybDCej1SZjskjcCWr+g5t4+ilCZdo/7rg2lek6JqYDwK6
qXWS+AB5GGcxfF/Y7LI2qGAAHasQOVk7V7WTHaFErwwTHxZg2mpMTzhxQgLrF8nu
0Iu0NcSwqpytylK6sCpoC8v3/tLXzHPCXGMZyg1AhO80LeoCT/PIq+FNBQtoZen3
Wylzi1W1ash7EJQqEV7ey2Wj2xC47XmU9PtMiuGYfGd/JAWkKPRMhOlSxqEwt4M0
kfamew6nmCLn4pgZr+EtNcUdjWpG4nfKwbE6odpBPTU+1WH3du/nAcDLn6rWOUq0
SwOHU7+wRCkS+Z6oB3kzkuVmcVEFbfukALAR9TVxVw7SP583z8gC7rKchFXqVFTN
nlSMPfOqnjkjFQZ7gQ+B0wHDYgqgdqv07AXji38mK/sppqmIyvEgwvr5bNDJAIYe
CBu6wU8KvEjj2VAfn9hwQoVHUFxw2dtpXtcYgrb7VVT/z8hwBAhdZjUtwEj5PT9t
UBgMGiAsKSWp32UyOo2DuigZzgoiH2rkXMNGzcWYoURI+Gjd0Gr8xQfbpscmRkzR
GQuWCZC3ifDhVq7wBzqBB2bG4EcvTAeMKi3jU4vhvety1vhifNcPGaOCsQhYQ4DH
ehaLrywWYDorYTblZCstnFG89adZlf0n1JDcyKWcb89mLfAGd7i+3V9bZYtFbh7Q
/zrk0GpJqZE9/Yfl4A7ptF0KS303lsP7bUUzEh9xoLXXUPEOb17IhFg0uGvPShsb
xQoyqiYi9X3X+T5d+OD5poHr5sq5Yc4kT660j9rEVFRvFCHdrt5PN74gnzm2ETOI
morRsfPLr1GDZJza83GYwEL4Y43I+VifvvNP1bERkkF7GWmWDXQXBT9LziP1t9e9
dkY9AN9yIrVP3LHsOHe3rMKpTH5i2rmY5UXG9ESiE1UP+rigi6KvM3EM0UG7Emd3
vB+e3XBb63/RCumcwTZhKNGFWQeoFhMWjrb3+ac8jJ9rmyKP3MMlWrBxUr5dKiXY
Af12nQ4wuYmJZRz04hCGkCYCHRg4gdmS9ls0XdVUDQFZYL2QpARnlUPiOKluZDfD
utPFlhfdYuDvydrSoHn/d/l7wGm3qTuWWCQqh3WTGmQWb5fiI/R/irImN9DMbtt1
dmnNzyyBcUMyj6JXboi3I7iJ8oXRFhr+FCa3bpGVmronJPfrGkdfsTen6qcOuVm5
fZqUN0CaL9Zms/LAP4wLeUi2XNg9NjW/LPkGfVTKhpk024wPFWY0ni3Qo30AixWR
KSAT0Gm0sdnBJJeQqtH+VoW2c95qyuE21zIrZOBeNUc1SPnHY0p9qd4GktgOhlu9
lc5FkOrUpmm/ImUBRHsrenOQqGJqWun72yI5JMdAHJ2KgxNEi4v3Q0qeMTOpJLsC
eiRW60xW4fPV2JjTcS+KvmrJWrlhKyW+U/T7WrM8qi6nKwQXZ3JcyjosUPBi+pw7
UwxpqHjdKiIfIAYH2tbGxWiLyJn/gGIQ/xns7LNHo4iRw+zQnW5vzf7Q/91/0uWV
uRGrukysjjWsB2JbmauJBrohpA2fsCGchWIQTEJG4mQPc4g/ropM5O1yrU6ezl3m
H0saYwGNOZnJ3Vr+ksRWBI5t/ZuO2bQ4Djc1CRktAr6ANLpIms14kqGpGbApZYa0
q4mgujhx8H/mUeYPUbrjBKF5IV8PCLG/Xsv9GnEOpGt4G3yC/fHLYv2L0PZVZf+Q
+PM4fz0SmRMCRuYUfke4RYYRPreuzhnXMGiNALp8dqoB/pjM2QnWS4o3tdqm6+Tp
THGrzdjrYrIA4unt3hcVrL4k4s0Fd8tmO1YLKXxRRKgNwlXY1Ax56xX7OBWpfeTp
uVXEeuTKgXe9nx/goF0oS6vLDXP/CI9jENdTlauRA2jbnVXDZ8HU3xO4ISFbtRTA
3UpepBA13BXD/axdydi8WMR6taiILSkYyFcyHhYMjekBH3/iFNdzefFvOYZRHuMR
c196dwzIjBgggZct3XLG/AEkIJ5udG3kUJZwqqmXjEGvUgl0iu+L3UvL/4Xm+rZh
verutyRihPf0tiKW3KFm50SRyrQVsGClzbn+zz+n8a/YolNm0cQNdipfi+VeXOqg
yvjk0e9dGMds6vS9yuX5jK3azna6EVrcXXbdvSiynCa778TMmfTvbHW+TqmmDkvD
/3GXwYIfP9bRjP0AKrlnoOH8cFly5zvOScG5bYkmnj/SCzlqwcVh5JMMzHAwExKm
yD4nJf+m2vQpQ1vc0dYj7CS80PuW6wH45VAdBumqUBvqE6VoYFoAtgV80fjDPECy
D7Ptyocw/YmS8ZZu1iIirNySOrXxrXHQC6AWHWa5Fkcv0vN5oYDGRVzYJinAKRTo
ue4xnypZ7yeW4++9wQj7AizCWYqRW82rr433V0XSBokno73ko8JI7WerGcxlULGd
N4GRWA5TyhOtyJ/CYI5kn5RpfyZMKGrBjkci4J9DtZ5F8P5H+FMpLAtTqIfCC7Rr
G04agKBkAVB1yo40o+AGhuQlsJZXxT0w3lZ9I6m+4GrnIX450oED+SaCok31s672
Lxs43DKO6EF+nAuSv0EGMDlq8ijT16hs4cxmYlQjBvvL13dDo5c3JzL1c1TVGUhj
S7lgO1DVEzQMXzIDG0Xjv1Qk7vr9vXOysBIQcH+JwnRI3f+6W1BIIA+GDI544gNW
c8DP22rKqR3pXTB8wsFyZ8wms0TtPkPlQm2Frf9WgWEnF4YL6Mc4rPJDorCpuqB9
QIE3Ye4lSPp8BAwtPh7NxnbimbyWoK0igIIrcKMWyj8kpGLxa9AV4qWIb4XNMmAV
Hema78SZUS8sjZTJmdhWQhwp0L/Gropd17mlbmQ69NxCWtu+5DEgM03XeFfEqL5O
ZS+LeOcBaN9Bl8qtULEHEhSak1XEQ6rOMxKoPnpOXBGYKnKDEVypMBhs+8PjfKvG
ngCYJkiqiBsGsPqDZUt/iN0aB654cc2TwYFGZgIQmK+amp/LYkgH7LbXoPIjuV2J
eLsHqLYo7mYJVeZ7qN0r9PrZYIop3N7ZP0bqVFnygLaiX0zk9IRK4zXLQvjI/jOS
b957tJQigWRnLihlX7LNwKbMyb+02RdkLHipYlUlOBYanhL4yGAzzQLJ38/vX0g4
I7qZ9HpI7FJuGZESBq7W+cfVTYxUoFrY1ZN1W3Gy3zD65DbamhVNNnkVZbxUd1aH
bIqmcgbSI2N1OW9fNuCPBnEhaGyJit9WKHzDj2MFmr3WWZUWVGLCckWwB9ZTJi1d
gHmokxB3UMTIwD6WNqd186HzGzwVuncLBtVn30IICQguxexKg1wVnr738y+ESJUq
7PZhNLNSTf3bsFsd+2AGI++Gb1Tj2Qwjm+W8VVM1vTisfnrrahTiCXPWj178mGI7
05hmU6V8QufS7ZdF3zRLa562SBsOMfB3Sg/ehxjdEM5nJnFDgKzsJE4Qwa2yIzI9
MUMR0CrWAnC1ynWe9ksM/b7iH0G1WEB9U36zzT7zQN2Yykhu9H+rmlvAdCRGvPxd
Me0eKJhx1MJyxPzyB+3KKF6yu5C0hAnLJ+RgHypeWbH8uIqWnWyHXhcWU/IiU7p3
seNALt0paTx35xXpHMgzXxedB4jS+haTl6ENKZpGgogmKjoD+B2BAwTxGxQLUATG
YyKNuHSve3mu7k3VqztYUYT+l8TOYBSIaiUszdDc1Q+CCD2a5AXTw64RRa9eu+PU
i1wW6ejyrmMrFs2ishLrem8JuiNXjxq5JmBoffX/FlOIYnUnh36eIJjdN6p3jNpT
z/mhqr+oRAVHPZ6/nl64XXCINbQI21sM0x5MuTikj8sUorK1gdeHZoMOwOxZ82k2
hSuwx0okWKmRwNMVpdJ9rjwINRjVNnZe9zQ7gqyXNMGB3Qi+LxJ/z7tYJNAZSbWR
TY7eWlht/qKVg8L8uNnmZp3Tj6LXGgZCF1yrRh8aJ3kbveKphbHLO2naD3BltLQJ
RXHNdJLO5dveXkw2B3XQe+o7miGmzVkU2dGShz7auJQ4r2e5cXaDO8HvGtgrQQqj
yQjFWKOvfpylKThlodf6UoT6aHoHyRpFgCZ0wH1714+ZJ/xd4neNcWUYWx8B1P4T
MiMMymRxCzW4IXoPQLD+o8DDuFPACwStLe4TvMqWVTMpVaey5RaKnbrUlgU2ZbE7
mZlrP+z7S1YEX/KZs+5MXLpX16MLoyeHFKKx6ybcI/XqGH7r7t1t/OCFm4tHHGps
YUAU1DE3ll46Ykpv9wR3W4WeRDZSsk7gmr8pF4npm2uYo1jfhydRXWxRZ8OFqMRB
+t5vFD3QhYBPQ0Se99+XcaxTMvQACZesr/4Bdnjg6cDqGc3Pgy5S6nIRzL5Dtx7P
hajjUUc9LF+rI5S+LTKgMNMsT6734MjczbEnrMPpwkFT4UnzejFdm362vqaixjPa
eKEhkCaHhbi/Jnrgwl4sX8eXRnU07LndTRScGKbw4ezZB3heL5f/S/it1nwFD2uZ
/DnhhS9sVFk3oRwBdNgg9DN1yJ1bRHxIpOU8+6sMJSZmrlFxwHw2YEe9b2kykM+Y
B29zzCpLDV4OkML/tCXINQuwFcW5fk+GRPmh9964Mg6rJf2K5RNwYc5jnyd3IcSR
tl9fMCT9ss22/53A93dZOxRjKuHy2pq+wx9kjkAroxkHhGNr9q4owGHsj2OHzPTP
+vcsPiF9H+pclz91LKyTVQ88KRYL/BSQRj9481a3v/4k8hPPCoOdxMulnbMpheuE
uarhldWPKY9/clhSfxP6kH/VQEJ8wCl5Gl0mwUIlSRwFtZI/FEzVHZyh2wT2AwfQ
njLJI2NMXNHWN0s9CaaNnWUb7SjeKbz4sX0leFljWbqRoWYSZK0zXl79x70oJtYp
V0eGSf4FYOZZDSn/kR9i+GjXlA1PO+heS4o8+2u1Kcq54/o8YQbtCINTDB7+AW3U
fJi18JlULzk1oujgN6i6NUdtoD+EOIoZGYFa1G5s9QMZZ7X8YldcMDVJbogBYaHG
+csHVLX3OXdAGb0mA40XNoAh7Tn1WkSQWFtleLuCW10q86rVuD4rrGn0Rzd6sWLp
/VKqB6BDQaCBDngkktmtRPDC0olyqkaj4Gk2e/TKFjKFAxHKAZiATHbCVfb2e7K2
RQ1wwxa1xv74xT0afACkgCt0JHgDoO2pmPGQH63GFiOo5D/0Ug+TTIRNFxu3nDKU
fxr2jr7Gs5UIHh8ws8qensnw6CjlcIyz/LXofKuyAz7cTIl7hOZyIHai1Xev5cjA
j9Vvi83J8b077umTQZ1n/fouGwCEfTuSjFkKLupnxeTkCIXvFSrclORX41/7NLL8
raK+wjMzi7kkdnVvM4Vl2euIxppbhZF6PYT5Y6XgBQHdpUO5IpM26R+huDlijKF/
9VvwP4cscXbQsklUF7xCFQp8tx4AOVdrQxAaC5WCgRPvWpk3BpAp+25/VzkIIqun
6/kUpFb0fUX4Vc77uupWnXXmo+soq2jQpNdvtYjlGV/roQBafqkUG+oZ7/CyZa46
EuQBIDA/heT+oXFBflFXHExKSIhR9cvRig3DYQk5YUQRKT6RPi7gBz+f93EUa4YC
UL5uvgg2z7qvYk1N6yntCj3VIrD6gatGZLRLz7s8CtuTwD6cK+yywYR4c2ANamQp
n7hDkTcrVPzE1eTolqdU5Io4rq2XhzQySTOo0kUZ/c0uTnf9wF3tJWzNl2SqzO+D
qXFAQSfhcqg34ltEXdcL0/sA6fFQrqO2KfHcXqTwzTOdsqCOaUL0BsQ37+Av8II4
b65LjKgjCiJtGJXIAUBNS3UulPl4q9PoEBuZfSZ79AEaD6bpztbQvf/IctnOPY4b
673iNPBHaJekZhHh7XJGPyrFL0ZWsGXsWEbxNG+iyfsXLnkTY0XHV950BcwNEDO9
BKvzL4ZWX7cVROT3u12SuY/tjXp3yrHg+Cq62em7u13k8es75Q7Vl2+gUaxLv11j
DLb+mjh9J6VoidP1IKirbMTnZfb+dA671a7dO7ESg5lUIaMcvT+X9MF/tEfROHPe
7XB6J+13/3PAwE3DDgGkYRMOpwm5m5+lnh6OC/FMUsK5Ua0KELX2TdGNeQmRrezJ
V+20cPiWfBbBQ6POSOY8ltvYMne+RyViqgZjQ7Gtu/4zhkwRlHe4molvsaIndYA/
VTaWLOD1sjgc4Lkj27XI7w+VAAYHvEOvjbzsaZX4zz02GXSzcd5R7ygVbVUi3VUT
Ek6dYDSUypP30/auKTN8Oxo6quTyNwNNxI8xyf4tGRFdD1gK1J9C0J6oFibXQG4d
WAWWLsYjwsA72R6X51EWlj4y5QuBDpToNmXJp4A6q2LvjORTf//fRwiwlnXl0iI+
pmkgsGsuL1m/p0MGZI7ue3kt4bSaaOqmskxBfMjsxFzdj4N1LM4wniNtVQvQAn20
53eDxnGnAkibq4pDJJV7Plh6T8Jgoh/VnxWPllRELjDR5H8btGAHXfPdu53OacsH
oWafjVnMkssJ3i32RaREG31LgfX2QOAYe2HCrc7Gm/n694ALv5UEBzYcYM0a34aB
1s+0Y3Gm/BHrgogDbspCFnxyChaUq5yBwivp24LRY9Zc8UHIj2u+SuMbClK741Y9
CK4HrcN/U+8VB7tT8+C6+0WUsesBLwZfz5b64NwTSLM5Xt/oYfok79IaexXRNmwa
YCn4A7S/Sy9XDV9JES8NvqrfAvBjqVQB2+z2niePSqkeOIhpL1pmSDs01I4zOpvD
WZyDjlIad1qFKqw6p/fUyl1iv2iR3UsYXs/zBERQ8ao3Np4nG0rJZUMV+jo87B32
sXIEIpUj71Cm7HO+VYrrajxnYcUKtc226cw1WmKYtd3IBc8O18WVIUB4pfauYK33
OS8C07/N59cTxMJVMn0HBhFtWS3YfMwj4H+yS5ZZURMXl9jWBhQT5x6S+jjcRAWc
1Fbw0SykQ3pjwR3/cj9x6Nrn4PsLrXNbZRzWmq+60j0tKcxHvarZkf1Tc6A4OhT6
31Sq6uPf0vSxkXAnn1GDuwlISsz4uoSDKrOwvGcZxHL1xihcnWCWGHG/ICYu3jrL
id9mnM80obLH7FqkcshrcaQaYrrHPS8CVi6q4qB4aE3l4L2S4lHH7ngLyoqbr1xL
kgbGRI1YBEIhwxjvTcfHZLjLjtcp85ZDr0s5qWzPxRE+ySMg3xV7oI6X63fMZkal
dMX9Exjsso4bcbss5QozmB1sMUljd588waUT2HGm2R4d3V4PU5S2urAoFVAoyaiB
D2/yquNBNAI2eRAzNqOT13h2qGqk3ZOsweX8z5/0wdI3BW3sm39gzzbvbwQ0xYFO
h4oYabPi89KbRiBM4K8ypUgobmigOTf20Qh2jotlDPR097mYJDuaw8OT3b/40Yg1
t8t7qGdne9UNvWPxKeQHJmN2mIAVJCOHSPJ4bVIDj9rACCcrmu/rK8HGYr7ba++p
e1/4OXGsLkl9gYkci7kBhTUMeb8jtrnhfatjDLm7T5WrkMfLZ2umF8JRvkljkdug
woepA2myblQ2hztKZlkMIWPEi4mYBUSPFdVfa5YMGTN7SHasMAjh44NZLsbObwAW
XBCgHNTI7wcjH+KPbVc7TDLvse+3cyuZ5gGfsssarFgixj7PqODGtFDZ1bNtttUN
zo7iLjdDN1rKA2KjqRQvi95yGyjQRh04Dcapxr+PEf2zePXJt0XbcbCI6m3XFldj
tJtP/JSLLcmLUBV0hSS06DXyecPhERRpM0Qdmfo7vgwkXAia3BIzh7iK/hKSfWAV
D+P9a6yDqqgMpff4XnBOVayY7efFmfbgWGldwORM/xKty7Y1IkDXXO+sXkpFxv6J
6aZWCiDJnefzT10JmCuDvdWuFO5ikbYvUNkU2vI5lvMIiTcsNhaqsNUZx8NkhxDN
y5QPyhXIiXwaSYoPhPGiav3tdM1k7vAE/MFji/qDaByBEa3D1zcT6bZ9/JjFkdHQ
GJRw88BcK8MZ/SF59d2WJXXzB/8XY1Tx8aHTiySqnxRSqMcM7O0Yp8dmycgZ6XtR
OgqowXRzM3BpF/nnFg5VjDfqTEkQez+lkIlbBw3Aca/po0UZOTqE+6rYnxRsjU9m
IikgGLKSiLRJOUO6jPUZiMjzceo4vPGQgUq+mPIMZpq4a3rxJTnhY7dgiJSOMR7+
XT7/z+3JAQ6ahrXHUtY3fCiDmcXTl1GAXhMISJniEDgwX+EvQKBsjlOnzFN0HF2I
x5TVqwr0k9NbmQjgz/lL0lh9nt5VlaIyKwlvyqee5vX9mWpZRuWYfLe8mHweXbBz
24lfv1Dmi57gJoIw1M6u7pyf0O1MK0yVzRT+DzhKzH6qBjjysVusEP5jIwB9G2TM
RN3xBWyjWHfCtSEYvRcOMatPR/eKP4OLJdbXmt4wmwH8KYyvL9p35YNJNaocu1tf
EfD6KUvWgS/InlRauCfC0UdZVGB4UrYSUlpX8ShqwD6ckMW/mluGOW8e6bmLoSUv
xLjSaarx3kmatkfy17Hb/1I5S2AmzeOj1S8zXgqLEOGRUHkGBW5C95wXawSp81qf
KWAF/3icU1koclAOgz3Rh3/uumHo4KG2MvDmO/c0sQzEo3lyeXfuDADar+09hU1Z
UN+9FNf4LmneYhEoqnzvz5tWyPjnO+ygQdoG6XOoSj1/H8DMaUdQ6P8fiRZ6b7t0
mdw5GwSCPsJRVu88i5ZxkHEOehMsQBZkI0rMV6xf3E6lmhb8BCrrkPuOzn4SagGu
lSG0mzHTb6NY8S12CPENp7VBpXMXvhpKy2Zd9WMGvhVt17eZNuX0k2xaIpmmwf4o
Q2DeZiUPZGDxoelI6Bca+GlvY9cj9iYmDlldgc9xdf7hSrz1AHGccMwrt4TScoN9
XAiYd+Sbw4w6lYYNhLSsFO2BpVbJpQlEjIn8OltxjIA9UxckKJ2SD9N5gGWq6Hhy
GevahSoofL5dkCvudFz5UYQNU1qBxCygnbQkDp1PcQ1T7J767j3t0tSvywOUnXFI
8y+GtAmFkaRqrwc5FIBkTpBiUhvSVt/PEI081LBVEWR96h0tKg8yCwjiZptAJXdc
hz+zcD1jJ2bUqDK/aIsDUqPEPu5hMOGZiSSjZ2jB0+qlCwgbHLYXclU/UPAkJ5jT
3muiZACgYT/0vvUfBlf1QMGtH7azek4hwit1xlMyyW2zBH74KWHJ2etpGb36lysz
Q26H4xYpAhv/NS190A4LJifA5alQjYzuj9dg/1/kGQDFdrNuegTUe3nSmenYVmLB
OqrYXWd6QC87keOVAmnBVL6fFg/ii6pyQpr1VA1UOoNbQ9M6NyUlIHL/5WtDEJSE
U4kHfGee4y4xkDG/+xXqGVK86FfaRe0ZufGqj85etXQo2hn9l1fD/gVO0a2EnZGh
RPP8oBqc9d3NcYe4lSnTyILJ1hUDU9EA+WvBq39hyVYjqoXIlSkT2lwz3qRYLpCn
OSo7qgBygix69Lug1jnieVF1B/+1BT2Pmz9jq3eMQ4QJUoIP9DLfDcfjxjwX5xE3
XxVBvdPZFa2lhfojd4q7ecXrCQovvAfBQH9zNvl/JStzPShxiqq7/dMW80BO/zM4
bdLgsa0H5Se+wd98ItZ7L/gFGzHK4fl5P50yexYH+18BiMRT1IBH95bggawF0uv2
m6axTt0DpTLtWJZNl7M6s9XjE1CEbtNG/JJJjeZcJw7kLirnusDw9p2pj8HkldCO
fVHpFToO5y8BIuJr0g1qXrpS3OFQ6e4PIweMXObyr23garX2NSqhR7lLv0eB2yzS
3UhIy/xreW8s5yqI866OrrLfPbd1sUkKQFYfCAvVoAlKEAtx/gklXDmilJeSO28C
PuJxQWDX3O3id0QYMPF6rETQB2br7kLUt3a8SWClxctsCHPXm79kOdYP0ENb2vf9
XXl7sfZqsjznuZawQyJznMi+njMMmxY8eUZ1uiI8u0Kfj++n6Ed9yYTOeXP3XjQO
FvDCi+TnBlfPDy6yW6US2grGQo8T7DgympoVHYN6CXWXAiscA+EpbxV2fAZi3coP
GGD/vS6ySTGY/tW7vN+lAR09ZlHgq0BObMnJR+C9gOVA7fI0rclZ7XPRA4fsY6vo
R3ULJaLkvqo+4tGKQCIq1+pu3LeIANloJsQ3VnlIdOgRORq1OuVBwK/2XHkjHGoM
axoU/mT79A5BOMYQdJfKBLEF5rf2hBrHOH4Kqi2M7V2+gSslLkmJWHsCOGU1wZPF
ezIdH0UF77rI7nqYD/5Dpr90pXMaitHKHZPCDm403t70wOFz7u1OLO6j2sLIhLw6
DqL1HR9LwOgCMQTvoNK2qLbTqQS7+wc8T2IsSAw0Dg+ZC9uWp/AnVw1WUDDl9BA1
XkSF/uFKBm0BcD25JPCexOZjf+XR5SnRooQcXr1ucyOyD065VN7ASd054CU3TtcO
mWgplj0ONOqAsAX3u6lTpo0dkPOEGHp/TMwrpIJ0/HnFBnokk0yDUpUhzS4kzCzp
bQmZRKfz/odXmIf2oWOkBVss88ND1MI9O0kABeAidBKL/yR2GplIRQd+0imRj2JV
cY1sNWknIKXVk2CMuxXorsgki2KvHcazDj+M5od6ier7Hh/ofU5vv/xSIHSE9ER1
HutTtMC6hXCM//8idrX37n6lZpAi+q2xxYRcMkAIzkHep+zMgY4nLiYiE3x3ggys
D7K1pYq9vapsiSPfHku5FS5yPwwVxEIEgflj9XoI/S65mUtmEUTvYmvXFVudKpZk
zXDHsM0uXIUQdlOb7WGXldAtTbXkH7M8c4UluMq9HzfWqj6NI0eL4ZYaXF+QfBpI
ZGI1213SoJMblmq1uLBtlBI+66lkMnicuvjnQ8px+9RXD5oyfx9ETMMQTHBjbQMO
uFxtrHxexl/xFWVKxDHpl8mJVEenr6tTTlnOwT6PwURtnVT8WxG/j7PaXCAaUQlk
OaNqC8wwnhc5pnwkTfC+r63yMOJJ4+WzkFIH/nO+xrihZ/j9OAyiabvPMymKUUuA
9JPnM7h1Y86oOMD5vLIGm01plHKDsuZDw2QhX8Pn8dq1uzbYkUx/1ZH31DoOTEHi
CpyHz3w2jO4akvexnY988CG9Eqawr8Ck0VPF3Su4vx7xKxgGqOS7EocjdrYWU+pi
UrmxQcoKZDK9JDb2OWsO8x+cJa8nUf3Zp10Er1dMMfkGQDUWfD/HX6YKPC6UYJng
w4Vh+j8x37Wuy4WKZPju47DUO5FM0nG6uh36HYHj88v2rGrl0kpU9pqyR6LlI2ER
CjQOD0JAqjrjFZSQSH0FWeQq9P7qcsKdd9DFRvSeTqAgyCq7lNUGDTOx9rrl+9Hi
1i1m6gKXKgXjw2p4fRD8yZJpFMM3YJ5F96XokU8Zc25uLDp8Mg7+1d8ySIKzSmCw
wyFPb8GSHAqo9TtifnV6zIm33fx+GDGgE1/70QcJtwhcbFSZwqDN9jb1cLpSKgMo
5HzHEjnr5gDrLsg2eUW039lRpvq3i8NI4M5b3YOj4vB/qikPiTCLsj4AND3kiO07
exohbq4V5XFqsThSSoe92D3HqQ3OH6i+zi2oFglcAh4QFiGqepKwqqcBMIoQmYSj
w9iszZbCFWCld7ykTD/pbmks7rxFsvdvBQT21sm3LFdqE3Dw1DwOdjlrk/ZQc+Fa
modSNefUdUcDPRT0bGSDuBG1Tsm40jAekg6R6XFgBKKAbVyUVJaPv8t6F+mOtqgp
fFHPv1amnzV1VFdnJdzOIMvEElcFDWLWnYwqbAVVoprSrYsr/mmMD+9jJMwRL7uY
cY28QWRFfiOIxu8fMHCPAJ/Mzo6LSgwcTJLcI7hvoftoqydbKo+po86enJ/vycl3
Spq4OkRNSTjolFkI5o7s4RetUq/gbWG0RcatnhRgxTsQ2tQyK6NCFvzEU+X1WBS5
fnfGQXwnS0sNewKte4kBKmu31nJm4VEr/VP+tG0WA9ZPjlxGnBQikx0qgJagvzXr
NhGRudfBA9DwRs/GxYIWpmChebBHiaOrizPQDKeZ7TsWpUU3cip+kvFnkC7eJY94
GN+CVxt8Rqzu9rU1AUvomyxsXveANnSWk0jdTINU5YytCnkHUWR1DDltVpzHa0vn
y2no0JIiQjKXFV6K5xiS/0+DzS43KnL4dxsiPvJqPRW33jo4VVnrvBCeCcHH1x0r
Yw6NquI2oThsQ5JcH/QIpMDCH9OriEXCCDCrk5NQvfLilTLxaxDTNom/LKNqIDNH
1qal24oBRTG7/aqbLurnePevsBQIuXSdiw51gNbdzc2X1lpHe2Bt4X/HBWov9qYs
B+k+jITVtGWNxzOIizspydQpqpfUCS6kOMMbFZkeKKMuC1AZGgm/9xR8ERQZHG2h
lqiRO9qzlRRfn8hQja5yLrquRyn3ncaHlQlzg1V0Gk6Dh8YyTxr5pexw0/vWjvHo
EvaRsAizjuyE3pUijdt0I+4+9t1Dp3sg7/8dLww336u94CCDUuad6c1XkP3OTiF/
9ngSFJH2e4CJmJUjMNy7eyxCx2T0ywI+Pjtnr01jDnNFuRMkTyS0ypayW32kTsjO
iF6GL4r4xZqOW+Pdc/rliz8Am7AqhYecAK6HME9JbSL/Ces4gbRdkOqhLLTFM6mn
sdp/1Vn6BILmps7SS4R/UAUq8A2EYfNoLRYA2mu5dWwV2N/Y5tU5BrfVN/fDYmE3
SxUM3tciTYY8e5NrxvA3ctqlxBLVNabwr1zMCyZzwsf93L75tHeQs0K4alQuQkPe
9t9xoNKsuDv0Bga03NEtwon/tdLySPayKG2ipEhPLNYAPBso8ilGwQ6aMwuTm1WV
HQALec9+0EhAKVQN/S8mpguMFi5MnlrzIA6cdj+lOsVOEOR+jh8bvd+wl3hdnNbY
Tov1MZRTcfr7NdmG1PfmgXp4vNjZYmOxVxq7kiGaUIMIgLjwhc7kQt179fWfYjKv
2u2cFk+Xie+uyr4k6MKBUfHZ+7ppBD/zDYrQxsONqso9SxKoE5XKXg7k1PDsi3KY
2e1oz72uxWFSg3FRPIdui2oG+cgkNdxlMyesmD4kIvdxU3R7EFrht7VfyumydBpH
wcTp4pkIFG/+gwZBFtP8zI+wxH67LzdCb7tx6K1SCXblRHQPYSX+KWbSbccdZ2Ds
/9GbLC9qWdZvksMkZuZU3lNqmEXRGt0gAA/Y2K254LJ2Yb9qxR7+euaPfXUmoMPf
I4MgQgP51/MabSZj2CC0MljGsmtdOY85eV9vech7ZEGL67b1/7aeBPEZDVDA1onU
uA2xQT+MoFCttPRVCT4J/ik+hEHbPnFOm1fwj1AenklWFINVOHiPADu81FZ0mEhb
EuCxvTSQs1z8efrKfIRHD8OM3kGx/q3CVicX7+d3aqfQmR/T4eDnc7MwrwGPVX4d
C7J8dosVSS5pOmJO3uCplTXENCBBrz942MMFS6aeP/xfZ0OoEoMMhJiMtGCxWZS0
mUpZ0spJBsQyjxUKLleY/7mgRYpQ72VAz1mnEYELYiRX8vJuyVT7sHHv13pHJlfc
miqrI395xnoN02o2NryE//ic22d400lEC91BFCA9WAsfP2ngb+y2CQbQ2CRVRCcE
1liu383P28zTMgk4g9ZNRHIA6RyVO0agRJGGJtRJiBVLei+Wx46IF6mpa/b3ggsU
r5p4Mkm5W35BQFPbuBM+HWzAfAbYXLfz+j68w6SycJN4rCgd2Vfi22PpU5SSTxx2
KoYcN9vBcrERSKjvTYjrbTI/+q3RfUnnc6xLbt5ni0x6xbtRtK+pZRa/BOMBKuZ5
B2TgQIqLvo2wIlHiqDUUMAbjOUNG5Er3bqzXz96uWsLe1aLgxjtRabhroGMcyTte
V0qcmHkWZ8em6qAgvfI9j93FeYs0I1WUkleMKTPwZQctiMs5y4BkNbmmJDb2eHEC
GRB1C371AjkBHE6X3rNv78BuIyF6qK/a8ijRBNMk9ER0aHfycfp3teZpvLUhXk3B
M1y0XmGzARw3RRyfjulaISkp/XbPNu0s4z1MJd7ET3RGoXJELvBAVcBbGrBS0lQH
eRha/fYLO6GQl8F+QNzSncY8IfzDwBQfgimhrzs/4XZqd0MAndr55ICWgS+oaxEP
PgYMnff1mrhwHxNI5MvTVJN+XRb0IPFzepfYAw1Kw793qxKJnEtU74fBonnaLVft
m36/GULrUXjqDV4k9IvbhLvwvd9lQ47s47g8DmJ/yVDnzKvdeCR/SBqZFMGgNNTm
A/cipEE5FNilDKfRiPxL8pdqldEgyYzh7NYZ3cwsD7UvhKITNGKv4LihQu05FsOb
OTZOcONcVFPqWg5lGXX27YCn3syk550Vcx9CoxisciaXpcTzCh4L7WOYTB5d3a5q
3qE34lUn5ECO+DKccK/e5/KCVWHGHsd2aCC30tV6rirJ2oMQrSF/LlEEKn3524QJ
It5ZzgSCio6ec3BweaiFIB/KTGBIyB+fd1MB9q9snsQJQ8+fUekPLwWvwSOBfZTZ
Q46JcU4YtNdQ8McfyRpHXWbzytEESupZS4EddCsiKPpTuWY0IxmrSHRvRKOyVxob
7zoC9GbPui7PD7AB3mFA6YXuc/pAeUboSfUrrdX6XEugEOytrqZX0couT/Ntxdlv
R25fwF1InVRSDzKG5xEzZYlwPR6tPttchVEGzkzViCtpDGi12GJtxipmgQ50bRsi
D4Xh2tZ6XqAF7lQEqr4AkRwuWX719QRoZY9cSDWX49qbRmCLZJG3ffCvRaTeYvXY
QI/2ioAzvcJLGnGX5j+nom9LR+git4OEMmN3xbniwblIwvW2AQl8YnLSRKPmfonc
lc83fZj1amf59FD7OItITv1GCCNuau26F/w3zJEqL3/NmG8o9h+ZjfLbwkpRtlln
OHuVetaCUg0z85/9BCoAdAA7MD+kgt9THsXzItxMY9a9Gd14hyLkASGV6rA0njKR
OFZyluqkdvQNEmPjy9cYR2ki/SA7ycfi0pzChsbbQr6JElIb9eGlhSDe/pxUqrCC
4j1/0WUb8jSuN40eCaTdwQ7KCXXfoZyn8SexemujG2qXQOMOAyq3sT2HlD2rnLpK
vs65YG988fNV4GmJXSm9wUM8blWABqVzL+ARPa7fOG4M4NNixPmZoDdwWeuGLOID
6/JyBfDb2x72OvWj/7+NF82ymGH7LSIi5udFZJIB0STvYEIuquV/Xx+4oI3+rLu/
7gdV1LhG8t+8kpmbDiSuCfVRU3Vn6M2vR7D8isEzTj+bArpuXuLP2uQSqc6lrzDV
p9PwvxKqi+z1p9skM3JhRui2XNWsyuLFZgHbS9KvsbudeaKE+cyLYd519CSw5cWH
JLflM0TLL9NZu3S6rCEp7QA6Y9H3Y4QZrH+ly5kJ8Vh/pE20rDRXP+eHw/j1+TKw
S+EA85GUcxtEdyxmyd7UoUZCyE0JKQJwZSJCi8FreFKhpiC53SdWcAaD81brcCjT
jYRyqpwMuY5Hv2amO2oK1G9BhjliVdNjxnFsMC0smN1jv4Bi/N/mX7588S4xq06m
1c+o4+oHzM6+ZR4gghpMtlcIJts3ETNmrmerFIMPt5MApPpvY+WskLd6HzWomEiN
9dRI8iTsBsRO+T7YtnL02kS4s0zHboj6tZSNQqACzmwy6j/rBFiAkpB4Ya0EpxS6
X55hMngpdoJMA4VGFCMX2PW1r1UQVR0MQ9SSQwbMwLIDGBi9wP9sApgRErbutK30
wFWmghF7noTEl+uPyY+xQRQ6qhGe9Kydl690ZJTanK6aX36ss4kavTnG6cvXzRAE
/iyB/k48AlHbdxtGsey8hlMl4USbXM6CdHPQo7kfJgUsgids/hnlPmQ7rZskOhi4
+fkshUK1ztdC2FHTdbDjHwQfdx5DuVUwLW1TIgiFCH6Upr8xbE2CapI/GgVNOVeN
amcYONILr2AeXxxe36XF9csQqurDEhVK6Ue1kGRvjqxlFzx7KLd73kxZZsvciR/v
7KStJ5poW8ZFbvfSKmMtlJslwFj/RAEaDNMQFZHcD1sb2XTRDQLIbz8IqyjtiTCU
Gl2cSSaDnvVK0xvX+H4oTZ45ZAMPy3Y/3W0POcfCq8KK6fBfVfUI2hgf5E9A/8qB
1s1GwAbeZ4fM+f9qYqVCH4NcCAyaZHihm4bLIafsaEQzLMHsbfdvSLlLDcexCBx+
TevR2fhMv26wUsevxAIeI7OCZYb/lk81zZgIC9ib/Jme5f5BrrDq9kFAadkM832/
jOjUH/oGzBoGPrA7X4gDGRrE9sHZpvOoiM6vA/WxZlPcQTMu6xq04FzLdJ5gPB+q
yYuzauC1Hk4bae7hznPTE2gTiWNfjvfYS/5VEvmMevgHsvNrfwyO/6qrDSFi/88Q
9+GuWnw2OTsrZjWTmfxjKDkx0TBRKZqp/qxxCJXbwS8hZDAfFWDiEbu7n4JkZMV2
PhxM+HHpzieit58agEUFnNid/EuE7j0CMN1aO7AilsSbv6Tgb1Dyc2M9ROP5AHpd
Gt82Nv/eFEP98mzU36NRCmSxfhFVM7x5kM35Utmi8cyrv2mGArmWW0+AgfXvhM70
wSRaLjacS7iEp6GhdkawJymRKpccnycWPRIIuXwWdJX5WtVVM3no6bQA4kksPna5
eAF5l3iwNWLflCRaRFeVDCjlu2vqyjz8vBGPRF80EWplBlzlbdMulGoIP0jWenNE
GuRVrnitw+RUoZaSoF+km7awOmb20N7Q+fiSdnE2gVriRVm4JeN5zIXscQ2FCy8g
t2Ks0H5ZCuV9sAEQPZ5FusRqu+CFmz+WaO8/s6pf7sDptrCFcyw+AdmwigvdcONs
Msop5vE5Q4X8yY9GqzYTEg8/479ahE3WBo9xy2j74Hxoahz4eB/Sg8FI0sw3y/gj
Ac3WlWOaJxUxb+jNjxsb0JN0B+BKlqzPYLcBLVf9rpx7EZy/lreStbR8sU1/K5BU
kAc/16KTnPzpFkYX7q0FBMmJE0k6/DRUcp52RXXc8uGURkspkQzVAHI4Yxtio14m
2S0Q7cxRkFUSUP/uvcEzN1ZVFBZPcys0cejiQKEpzbKeKoQUl3WL+y+rr/VslSrp
dr/XzQrP+nWw+3xnV8GF4Escs05zVx68tCJPoksusA21iE1cbW8PfGtgAbl7wtWh
A/wFebwqozC9cann6zIoRGQCzWDajG0ZxZP63Q0GS1PeukexwGYy8oISfMmmUGw/
6n6B4J25IKA5QWGKtFla3y9H59He9hCawmXNzOrCaB3koYjnO7j2vNFY0tS/iDE6
HJty5l39Ch9iLeMGFBabsrLhHEYVw068O7NBUwuPsqGqSNmhSLN6mrVMcBqqXAiM
qEKbkRVuXuTzp+dmfZPy3YuJSayXMuqMjiqu8FH1HX7Srl1a2ArbM14WKZKGiOdT
1QPbWW9LSLbhYj9FQ7iqav75C0sTKBnm0KS/jYQoHIq0urTSeOUUL/rGbAv/bG4Q
1t4XUtfhf8MOLhUcO63IwvxyAKkcrqWEAlYE7SuJhWkOcCANED/U5OI5/BZshoeE
dFEFMmvD29DK3Obf7KoRk+j/v2O3ibRKBd7bi+c61ONM2dDPVjMbIXUNJB6PgPq1
Szwt6SoG6LhrG25iXNv8lcWzNcOdfzTGvbEYwnieEtWv50zm6sS/x+ggGdrjihNG
vffAgzXsMvX5ZMOLiLDQNP295pn5o/TU4ZQc+gEyHpu2FV44xc2W6k+KqV5p2yH9
SqVQNVquxjULejHSxyrczwnQ+jWP0mJZUTFqa/p6SSzp0JbtLj5NPN4lbFOwlSPq
3oiFZ6ssz3R1/+I++jBWVsu9MMqChzHfw5njGKLzRx6uHlH8sl4WMOLQYPR2lffk
v7cuzr4nWjZAH1WAe//MUjnsFOPXfuI2eFnJrZIsPU99542sBDXsIzx1ZiJqkGU5
Qf3TaySOq/VWW7Jvu3s0cRLjYIlOFZNnXB1QXcX+mcWsLfK+PhGHhh3l9ZQz42kf
s2GF4/h/U/jDWjSU6aiWccGlFhzWN+Q7RUrkc1efih3eGIFYKj1k+RfyGj9OCzLY
2SQJWLv0iSAW40S4jFPcBcenD2kumAMN7mwCA0Vs2J95xft82m4WwXU4pjSf8oIC
eTgj4tLppXkgFmGLNE4bX5oTQfdUNMC9ubKz5QsK6/BnhjV57UT7nHOqWrBW4gPi
p7etjKg62yj/li9AjxCYfXQhwr+mkCedi95H6PtrsTyCzO91gEVqALVKRqU+0Utp
xmHtbDlLvv+oN/grLqOVVlnU0zVFTFmNM8eeHBVUCsEYT95lLyVyCA1nR4z0B39E
LOs97T99gfk2Pv9t82ZDyE16gAMGa73YzOaR7kAT58EPVuQ11K23OGuqWy8yVJn6
jj+b0aAd1FSDm7UQcv1/HWfI0jpBzGtqHPTTLaLdBFTx50kZTcvT1dME2QQDuSSb
K/cuTQuPyCUnaJFZvnQPRTJLBB9ragT0M9HCFt/tGZ7FoijNXDudleS+BxahB6Y0
aKuBYAe027tm9vA7jP40+AKe4jPQeIxoLDxhvioUrNpt1aho793tCb+3jE5nNMvq
7xrYYwki0GbwLdRF2P8IamwHFch8RDDfT64lqK92IkviILa0DoejwCvYo0+8USDJ
8FdXd14Q7FHZBObKooc01yD8JBykk/RiZcNY3axhMMzRiueYErq4bldPWyh7sZ97
nJlmzgnyGuktbMU6KbkaCKuLhhGSm+OERFKHUXYFNVFiZK7c9jKPwn+A0lZvLVOb
cgazea09ZeXypfmOhNvnYkOMUoqxfOhtog4L5sLJptLJiiHIzqfxeauqIWOrlZIz
CmhpCQCajSz3fxp+QvXFedF84pQr10ldxD2JqfXQDKvbhC1AXdAHT5952jjJIbDv
tdim8unlDkWZaGjiXx+jV8TEor/nkKliQfydJ9TDcaxIEsUMP5fDGwBvF/SmNmPi
0tjkQ7S/ilQTgSVoUJ0OSuV80axb1SPLgu8AA9Mhu/cJ3ezo0xAgp9E5PaZH80dC
lHl27+xv3bbpvzXV3VAO14a2bEZCE4ulB/Gpih0ZB1JcOe5897YPHtEgtvSvDXo2
95VdlT8FCs7xTnazA24zRkRouZ3q+YLahnslQQw5Mq88UGnTBccC/nTvmdpBhFrQ
g2jgZAJQWzeKxDCE69FDOzYJ3sSVAPNeTrGmRTITJlg1hyUi2RgVDK2flRoeR7SW
P1rp6Viv8cOuvCyaDEjzhp18Pxviuq4OQXcEyCZFyLR/Mi3Hotq6MzIVtb0T7iBA
Oz3Zj1WNtYX4COfCsUF59gY/kBehzV9B6DcrumE+IE3r/FyKunedDkMjG04Vskom
RZb2wkAIEL5EkQ6MyXhXlvWrJCVq8VaA5oun77MZS3+piUdmXtcDz9SOWTi2OctM
rnN5uY31/ys8q+oYa5AhIu6pGQx1TIV7VZVKRtqug48k+N3Z2bjGRI4l10/UGgJX
rcUF8Jhb5ci0VOaL9cbwatfp7NYDNzI1AWoDuXj3MmKglK+mAOBlZSUSB7umYMPY
3QRiitYFlN3V55CKh9B8j/PX6tgjCzJDo0dJJ9JZQueSAIAx0cXI7GEZCjUSQGHA
mI3GOkQsgpvPxnibBtp+Gj0xmQD82g2a1ZWlvy9NOzOtN+9PZi3Av+pPOVhxOa0R
pvYBhYKLEcoY6Cky+eKQH0sAHoeLMqrq2Rfde790kwKvSekmwNCX5JEnt9saCZmN
3ClmCJ7lgkjLFc1qb9OatF/FTC0JPZo3N9blGscFLKFtAt6iLS4mENzoAhd/7tXS
/mKHSFnpV/DI/We1dt0GJgg8jRDiZPIYS32sr87dNGJezy+PQ1vfWI3YKH24AB1f
wR7WTAqd2T2PTyHezzo9NFfjUql1H7WQOnQAvWwsPJtxriLDKVHPkEpHB1PnmzrY
alEeLSn7IuTKpcZaEOETEA5KN48zPBpahFnkcWe9cmp5B6mhlK1that4/7agzXi8
TIsvEbQKzele7+0lecdE2ZA7UeCft7DFxgcbKKk3tKpuDYp+7jRVBEJFXGXnWW4b
u4fBQS0YFhW0rI1TKjUWCmWKQ3zZt8HrBmmchodt/BdNYnpwS+1gTtNwHb+534VT
FW7y3jrG4Y09o/HVIGNEM1DswhHFVGej/Bb3kiUt9+F2Vdszgr3RJCjp4poX178+
qGCFNdsHcf8C9VQb57slX4fVjtn6mcgYfEHYnODWjxO/43hhlhVKO97J9ftmQEfM
VnVySYMHVblKcanh0WXEG362BYrjEdpiTEMaaNHCDfTqM8HKsR5+C4JoaYaWoJbC
oPbb8r6LSrnYs2He7eG7vqQ9NIyvh+TXAPrbEuczcM+MecsFuXNtCnNX6jZk3IAf
JqG2OqnGfSMsIwy5uDKrfcSwunsAq1eAakj9Qh7B/tG2WQ9pCegzAcWjVGExPOiK
I2565F7qEqZqtnegFXdZ5vaJ1MQSw9NL5WzIB/3IqLdFJ1PHnexGZjdFgowFwnMD
52N6Ip8EAdihJgJdVuEhi1LvEGV/id0m1F71k/7w7uG0+joRsHdJi8jWbgpSUAnh
+v5W7v0LYomThI6pqmddCChm32xyJ0dybQbQF7SCi+6NNIIvf5lC87FGVa6qVvUK
y285kPCyYMXnEtcKUUvquBoTWgkf/RLdSZ6j0piRZL8hrMUXUMFBPEg2n7hyrFcy
dl1bgbExzfZVZ+40sETBHtVf1jdBC+ixAOiZ6jDTl+jKtsAirSnIfC8X05XZ0Gph
xvMtdIIIpYAMO8rWU+g554se1PMWChKev0lJqCpeGR8DMAfHOe3IcLswYYr26Cr7
NyRfmhocHUkzi4gJVvKYyTgwglxQrb8glJAlD1rcloqB1JMj+n30FTZz5hZ5FY7E
eoPryfA90Ck/uwjN46RcicKFNayjFiTWMXHxl0e9rAaMI34RVUlG6SFjAAykGiqP
q51UOjn1rpZAIVrwSeu0XNvHxApHQ1kjMLbwFJghXIskPf73fuHZ1hndI6iZdxU/
zhppntoX9veX1YflFx2GxjSKBAl2e9LFVUESG7bqcZc6ibtWePhauifWjqIP9jat
wtp6nlimzA47rfhGYdUnRHUUexAVmPypg2DfqVq2YOZIHwbUt0xfSWmi/5/9Iov0
wH/q2zueEMYSxLgiuTKoaOi4trJaEtNWUoAlgF6FsbcC9dx2GDlYwykZePicpEKK
TwN/mjxuVAmwVxWYZwjb2sT/1wMXSJiOWsx+AZMIWYO9CAsD7MzGO6hSQgkPFnaN
+lum27TFtsZ3VYetVL5/ThTPocEC+4n9wCX/KuoygD8SX9frTlj63Q/LYYu7MgPL
D7362HTJiynCo/NWMRWruO9ptJRNiNfxTdkch9ZfzoO1gxSAE0ZJVVxFt4rYOKFl
v+zhJraWKxN9AovKAokzC2xw1m26G/5QbBw4fDo7psLSc2NB2Or6Bis8Wb5r55Tl
XXpiuIm9CMyM2OsVtZU/zxgI8FIyUQ8A9tT8fsd6IalrDNRRw/gS2YH5P7P9mgF/
rsifJjZ7Gxv0xwxdBC21ASLOdDfyMY8+imNP+FTzcFYGlNmAdJHF+mDbCPJAUTTW
ziFZT2QYYHGTznNk7bitL2kDzMrOJ5/ovmpnGZDzvPWaz4Aq4rNXhNjUY4Q6+y2y
aGFWS7Us5RxXbH3gOkzjVdWkQo0aY1ct+XwPN70yOENRodtsIg2DaLXgXC+5zW1r
Ghxqc7w39xp+zpeK2usDZSgCdzWqJmfpQ6+AOiLX6SO5xweu5RH95DaLJmEc+sm/
RrN91Z0Yd+CkXa7cJMLQdZQ9oOvHNU4x94wnd3adXjqGEZwpZ0PwXXgZ3FtZ/Swn
TTWJ7GHi386Zvd+3mGlXQG1j2ZAjSfE9FA++6E+UBSwS+jxfVw/ms4nqb2Ll9Sg9
qiXmfCP8kOIBscNq4BUjp/rsBcTvuNlUXxhWKymIyMr97FvgnxPOsmpaSmZO0xkQ
QaRMR24LvDPJnWniYPchnixr/umdlu14xRfNm3jOlZpt89mvqqMXHEwAlbFN2fRF
Ohy7UNKRXpEJCjlXKBbNaOWa9VPTl5PY6gf9JDHMw486J5s5t94fu7LZ4KYPxHKS
9ZgidgvjowEoe6fw43sUwQLABVRuyHUMSUcDVIHEBVUkCpR2/xAeo0i2RlGaabzr
AqJR43jhDxf1SQ4ziwbSB02+tmINr4s578dt1h/221DdD2VSkFQ1olUtJdAutKDn
/hiHbn8yoZH/KJCtiNEc6sH5FpK6NOf/OP2zl0eHkhtgx5slWdosx9CihC3aBqfi
HkcxRUFa7VTG8oWuM+v6a/ho9B2hojoGebv/Hjp6ZOCG/gNq99hvGNyHz+PkQlrN
8KZqGjrmUWXNiW8hzW/44kxB5dROlYKzCI3Q2ky6XnWI6lON2fGg9UPuE2umnaAQ
CvxpWb1Kz6jeeu5Wo6PWkJL2spp3M6cBlFgWSvMvhkntAA88nyS3HfnIWr4k7Qat
xTV4ypjC+3usKC62k3aa70yCkvQI4ibN71dcLHhUwpne9v7WLb84qGBXI+H+wgiy
ClTDywPHDqOK1u/g1sOF6Pn0eWhyj7jkDK7zZIuLWyInzQXRk7CiNWPCaukPFgVt
UYdTORWLuGmtFF2yeNDViP/jWPAi+8xx4NVnwOfcbDFDjPBB61BI9k3pa7N3RrLI
R260cf16y59a80rFcbVV/NP48/InDqanILKto7956vgDKfZU8FNhSnyV2zrJP+iF
PraaKtoA6o7a7Xbb6DlowDCXxBZXhJQ3/m+aVInTEvYKZU2wlAVoMJkyUTFcHCCF
c75KHFsi7h5rkzgU65hdXDGeRb1ZT1/YNsOE5qJHWUAzHw1zZxM3WTNIvm5KHf5I
1BzagF4DtS7h0VE5HurYo9J8riUx7CUSLyJ88Ze2a1Vt0cP8b3+VkhPOE0kCPcaM
wgJB247GcrToJ8VBGW9fqH2da+Skv68tcQm+Y2ErePNQnFiBnSc5Dj1TMgq07sUZ
GXh1p3nH+my4LKZ8+6wkFMXwGbnCC1ByYGmSZKywzps03nrt356ZNLfzcRrHdHxQ
GHvEbvuPSld7JwqBMVtuSoCjSPfTSQwAzUSPgAA6wyJ4NP3+wTPeJMxT/X8PZqaZ
v+0Xf+eBGaOqgihTIBJTt9yTWKtMRKgkeMR5+DrVV+daSwOlLH3/vVxKWRBGAzO6
Y1POAFaqwv9BkYWmav0D4I65ygrPvAibUap/cuVYSv4hWCIyiO8V0gHovaW9Nbv4
ef+Cpa2/2g/0qJawrMS1r5vsg8bMVR1aA1/1eOw7bBifc4GQE2c7/+W4t5F+Xnk6
8kNUgJEP/OJFOyd9mE3V9tB910nquxeSw+qnOmEB4rGDAdkKl/D0RR69vXwHc14W
RcSBDPOA6At5y5JacvJ/UjCc3n8xrE0oV7MYcFI25w6iV348AeIDym2yG5KApas6
18YfThkuz22m55BrkXLLhiZ7xiiLb9EVzoS61xxrQuP+DZJaINP3hHK7R14R3NMp
KBVjJtn3jTLc0aKKcPMh3h/9ImOfLDlTqvVQre+CrKV6TCjAWb7TlwNwdHr4j5Ag
X9eCDC9vroUe5FzA1tlgcDaSjMO1gy9VAD0dsf6u1eIB6+vyucoGkouHaxEetjMg
zmJ7px49nDeloFK8I4ELFz9iGl/bO+vX+4vleXOLx7LLSvGESdyN6Wk186dMu6gh
eB+4/W6ihCAQ4W4d5JP9etVEhf7lxVgg7KAuYmkwGNWAXGoc534aD5U/dyThgY7S
/uVDEe+sHwDUU5hAW1jO0CBI8yjpnvTJKGVpQ1uTqNsX8HJtGYaku1/gu+B7QZBT
ALUy4U61uN42xyQ8H+sxvLoSydKNGn1H8tbCqE+lkl+GS9wlRGzEfNV2R/dfFy7Q
RUeoRRFC06kr5YDkwcvA2r9bto9CaLkjP4jTsv1pz2Hb0OkXRQw3scK8vhdjeJG0
zucpiu8B328rjBDGFJiN1+nm34HV1zoweOaNHLLpeJFyZ0lHBIu1BixMDrffgEtL
C1WbaslQ7nkCwdzNU3S0070SOGwJkscvHuf8Ys2jOmnIzXZEbCk+JgyIgoib26ZV
JEm6z/TW3euv9XHhNTw+k1Yn5c187Eb2wKarG6PDr/eioywucxzYNs5GcCCxsUQ1
M06rxESiq+CnEX/DsqyZB5isoZH1n+lDx62PzhF78FKYnesV7jgpquxh9BRKfyzO
yQ9EtvlWZnQ64NZqTLwebV4gGHhY5GoAqKQCSGSskvSgbHEePnl/LIqjWZwm1xcd
dwUVvSs/zr8kBcGXdMZ5ZDVfUSXtLVIkpAkaK/FtUS1QFp8fUrzcYkasdtSjtepm
R0rINPhPJXrgZJb5r6PZsOpoFY+mmXEWfr4OWZ0vWdNUD0dQdEnNd8mHHBIwLXho
uoHULtTVpsoM5EJy6rSZAol9NpRvnEiOQbQfdTFAKppCM+4haRnFQA9Yzeeg9eLs
Z0d8BEzXnJi95Vak9QX4rTBGJLiSvxiAVL6Z484a0WPYjoVltwW/GIN1YZTVFrQ/
UZqBeeot7gSkW/1PhmftATqZyRAk0jD7QWcHOCmykbAeucYCfDamouLyMYqru+Mt
M4QGH4N+EsWe2oidxYMpDD01gNeTzU6dmgpRsHZcFD2ueBwYVRhmXgtQHYzZC9AO
8Ylne+iHCgljuddajxsoONBxYllbuG0DRIOKMeoAwqnPTKNfWAf+exz5ICqNqvdX
lYfh0f9kEIzgxSy5bjV6PfV2YS4K+lqoO9j/KMrkaNMSENe2n2a7aun2DNzfZhRx
2fCACjTyELq1IHiY0Z2QJ1Rx2rKQG2CfvCrbLji0nDo7RUqkA/DobHldskNrqW7X
Xx7v/rluVMLp5MgkOr8UhBZSKMzmAImOC50fweygFyRLMy9joLwg9PyZiS5vWzYo
z+LdL98IREWLsxW+tTM/8LTaYTtFiPTve23RNNIMOU+vbJ28L/A6fE9pJqI7OMIM
p72cubevx6PKMxdbqg0ldoxREYZ93Ib3/zAJaWdwZzSSH7EuV/J5KG5seNAsP/IZ
fZ6MGfg2x+ehfM2/I0bQRWQHncc4JjLSN100dmBminjqigQwYfbsItl4ONv8Wf/i
mxEvi7isw8ZbuZtcc7SrK+53rVX6TcB/PQLn3NA8WolkLCrxBFexWJkKRTfsuQUS
MtJysY+envhMlxlxg3LpQK3F8FKpUpqO3V54g9ogEYhkEuZ4kubjIPxE2Qh6LAg5
Zrq9m6iv85+Kcadl+w3ptU1eal12eBKXwWkCbqx4B6jbDGb2cAu7dgrnKrHMtao5
EeQQlMXb1O2yC720aXpwLKI1j/3AT+6IhBgAH4tv8VQ6rtyiLb0RvRWimm1WaZWw
AEdnfwe3fpRhPyUCuobgkjGvptB/AFa7iK5dg5mtkqAQYEJ1e7G9qMgZc2vF/zyy
za3jrJyI5rr8gV6WPp0Y9MGozQKEwWwGJCpZllaCqtx0eGpX9scQdkfZ8VuEJO23
50YETewi+kbF1MIkwK2WhpXXHIRzb/AzAl0TIIW/VM6qcdbhuY4b5qyjaeo9Vn+c
yUMPvvF1eUNYhk0lzNAzzh+fCpmMX+/055DxVGrFX65wKJSkZIWU2ESP5gzS7EAj
JYs9Ts21Tcw9DzT773VNlTJkaK9QfROUWbZ5Xb/6Jts5n3d8DQnY9eUnokpPyBKB
HPiAIF+pLsCv7w6an3D2Y+KD/Yoy9eaTydy8XNjA/xrTN0KsO1C4qaUk/DBAALOB
ERACZ2USa2vsNJ46KPmsZJzfrDgtCvMPQ6/FNwVxS967ZVTcMQOvz+VZAeOmAZHr
o2xptcr658IQEDnRgKKNYNbZCYJ/OjiX0+sJHFDrb6h57Ne4MqBS7qx1Sr22s4HU
lnL0rCO4lLljurG69RxUAMzZdSMYyw6py4q+vt9SBrXnuIuHZGVbVO2wamAGBJLr
S8Rw0a2liTmXw8uuSANMUP60BCQGCKROpaXodWxoClcEl8gPAZzU2YylMkgMeIY9
r9Tka+/hXHpqyqX+06m70ZLZwXde6t9oa58G4n1dYLi7k8LIrfmgGEf3aFBKjsW/
H+L3ZTv8dvzlWrDVtgTacb5fMZKuFTX/iTqFmo83CgxIyuoMVrJM80k5LDd4bXB4
UVxolE32C26XQZN25ET53YHpou+A7YrKGL/36GdI6CY2QhqBWE1qV+jvAltdCTmt
RD29jtYzDLiQphcwvWeI6WmtDOBpYQycQz/OM0e+uVvIHXibklbJd/QYA8UGf1kU
/5FVSz1taHL7YVeT+fo2ehFlc5QUaW6Zuqlw8VFHcCSLUZX3dR5uTI5mtnU+E3By
WtbaWnVxCZ3ocSQbydguL3ABgh4LUU9Nz6z30OENylKKj3Tq4eMgCpE28AbwyA9c
Htelib/gpcWx0W9/Fqq7NgebYwqBn50c3x6jzsLVbvnvb5xXaUyeVA/dQkOgwsAz
+WeDWO929JUg9MVfdCo3UTlk+V6iJU0+REBziKdVEDmGHfC5SeDlpgWRZvs06aAG
Lq1k794qqWtTqOYdssUbQNWSclUTm/KFPadQTgnQEj/4X8ZOTrzDSYOdA85QOOBz
HSA8Tqwy6vQy83R15/StSeC4YeZlUGCR324ES2P6l+DSgpJXthxpw/SyCpcNS9LE
UR2H2lY0og2SVHdTOeOuAuLE5ZvS7pmuqr8QkupvrTOTm7NoKz7g9KZLFZR2QhMV
D9ABHcWEBw/FpQIfNQgxz8fNB5oi7jNwnzT8r7MR08ePlxLhGp8lY5MVdcNe0Q41
iNZze1DzmcObnqEUC0kmoD/NBcq6kWEm6wTATXW+LDdQ8nf/RzvqsMNJCwpSk6IU
p7ZigumfB6LD9VTRnXsQbuS8t092aDEg0IviNtcMdve9kfNJkx+Gaz8TZAnJvfya
iGEbtGwQprtHCHLy1dqomWCtcFj7jCdX9sSRxtxBiLG6HskIAjspriY3tpFpkf6L
KBFTpdexdgqR99EKxxZmQBsXk3FbBO9uZhQGtkrUl9B4xHg6MGLuMT3Ga0H0IEvr
Fw/4HYUUp9i+CSu2m+BwwkDkCy1xOTuLj9F9MNHFdVoEzUacbGjo1svGO4d5rWR3
PtBr8k+Za81FkQ6CGVOT2RtCyiI6e3jkgY1gpsEHiS91r2H9Ypu4aYxRGuJoSqli
IJY6gcDPklmLkDua9xGCztL85Tn5SnN1MVuwsKy09hL0+84lyX4DMaHaJNgghRbz
+R6vPkRgKxYu70dLT/7vzBCmEF0iea75wJwka7yAM7Ze8MSugM5PA2Namp4M3v8t
HPbiPlt1VGGCYHda6EoY/gOuVttItUwhc6TajLc1LQwDWPV8p1I4S1i/u0xMg0l8
5aZsqhfnC/CFGOC+ty7AMLpxi+Pevi8RgTKpmQW1WVH9HOhrtXMBxS5ZfGSDW12e
ssehEzBsIwOSSh02lPR5OQFfkf8ubGuztv6Pi0WywBigorEk2zbwy8KYo5zan6ta
hniLkEtExfmWUCRK+IwKx8zBJCxmXifGGkhLFfPx7260nt2QUwZ2H9O5j4+aWVUI
FzUbwXyFfCtlmUL5+bJXzd5FtIsLAAye7MsolXMoLha5eWXloObVg6O/CVdkvz+M
fQzahhfD+br1DiV59+lUQDx+pOccfdJhkQEcxbLkQ8BPyTIETMrb3qOXgyZ4ZdxJ
hmQPKb23XDXXy82F1XTCGdao+axSVXbUiOcpm6MxkMD+vCM6TYQw82o9EoriTiCX
/xgZMEl11jG5ygSINCM0HLrwTNsRTw/9qPy3OWfva5HenOOT/P9Lz3vGeHhvSf//
ASoESXijOZyIktFmC0hLyU+kCpewnZ8CTEIFEfO42cRTvGosP729kDR26DTltAwc
vVQVkhte2+RnLwBhyWbaAHBxRnl8yIeUKy1X4lM1sUl26MD4LGNm9biqZAwReE46
zbfQWskpbMTdOyVez9rPfZJM3ni/ImPzxd6KFBqh2YVfKgkB3xZGkP1FSTZKmOtd
BJ61SiQxGcRF0zcqdJSyZydjaAU9/W2HdNVBBdhQnuTgKd0f75P1/hBjTKAKt2Ai
ROTtNSAG1i5DL2GNQ7BTuyoKrMdiat8ZsSincy5ZW7T/4X8qec656snNUdxsX9BX
zFeR1XNKLSl/PyOvX5LFldVaKW38YCBVDxDjwyIh8MLRJCjP158ztnkwfCXr2r5M
7Qs9Vo5PS44S2ztVmU06/PvAqjPm3zhoqyLo6eSXgBGi1VQ8YsrrQV/FFXDZ5KAs
OqerilqZW24f5RoAmCZxtmQRJcDFklvwFc6htXd5wmD6sJVAwsJtHtVU1W9MYdU6
E6WDqyeCWHQNuK/uqhUUeFs0A8mIup7X/oCYPFifacrhwMpz1Svh8rUUYVrGI/fr
hkbpr2WMD0LPpr8vqIfAMdC62JY0a/PLS4vj1Au09JaOTNu5yZJCslLNnWxTJGw9
3xkDpmUYEVcuwiH6O8ShV5rDT1eBCcrgnBbnyxLhdoJou6f5I51jE2ini2uphDi0
M+GnpgPioF3ucKHMkUhHmrZNoIDBKjtJHUR7tVECFZ5TZSqkCiXCOIngJL4i3OY+
L2orkC7lk4s9JSijAfkxj4LvOlQQW05WuLhozuqXIDr00aVgSc+1GrYqcFl9CKUr
bAMPmMqcG/rWgos1HLjSGx2lWnqAqhTu6alRompR4Yu6YyR/2uyx8KQ8pubHYyh6
AJy7BEnifxcsfWZMI23OSoCW89nmokQmsiGyoZzqhrHZgTZtqCrNuaYwfXHmPcSK
M7nct6s4hK3/4trznqUcJ5u3q22aDcIdECc8tZjU2izkrDKz0JauF7yGJIpQ7gYD
xbaJjhrFSo4RL2WgwA9n2WgJ6Am+gLYQKHWUsvbakSqjn9wstDkzTjIu8JRShiXX
t5nxDBe6f4s3ZHiiAbDKk7oa4TefsWFu4vqfvZeqvLX/Pt0U8wQgTEp7HeeXk7gL
4vTN6lNdcNvJLCvVYvW3hfv/TdchuB1qWog2+lqIk5qNzkf4aI1ksSIy1jlk2pyw
LUWaJxu5/zwv1MeHdkDJ24SPnPIsagDwXyZGVEFiUGLyvM8Tv/BYBO7yCvbfQoaD
yVqryjgQI2SPD5ORQ8PBHhxN5QM5jUCjZyzewqcNF+OctdioiPo3ThseUcf+g+hm
ODrbWRwfL0Qdwbak8T417vicSwLZ7P9ED/36fklOAbBSnJx+PtEUrCAF9Jb4fM39
sHio+Ol7PIuzySjub8IldjOxn6eC407JlMwo6kLC5QEjF5jWRPeyZBfh1IQ3Np/C
Fm5g4/HRze69tzxJtURVKTeLStuDO/073hi6J9fIbtxIqLERkH+wTng+2WcZi1Nd
GN0rC/EZqcqiw442hshNmMI8wgQawwfrQk2WmB7frxiywBsF/PtXqHUJR26YvAJo
Bokk1G/M4ukd/sL1suZmf9BiZk+5Jl1kEXPafvs68mf9Hx4eFTuYaLKWCasy12NA
hO5k2tJjrkj6xFNBd1lfastLRSlSn3QTZ3QFQpDuecJUw5HHP9QqZsJaRdQj8urC
kPsFNJxs++ytizb90WOGnZZAkqsVuX+HrPepEO6viqrJJARypkt//tYvSuAQVyDQ
2IuNIPYCLRNKiAizxMs+60uTaiV7gwgU5FtC2T4YJhZO+ZSRx5X/cSmzLLvaKwng
b7BUPLX/bWNPuC5P6OCrPpOAKwWbinpvTjKPR9nVqMdxvlE3XUl3iStVpP/nQVtB
U36qaXvamZqSYD+bBx6YrLqVXoQSLcuNaCT7YLAakQO9YVqsevBupwUnPlKsKbQ7
IzXqyXigEM0PmcprJeVW5N6fPbJoiPAkFnA0YN5Ysych2a4HDvAlTsMtvvWMUPtF
p5ZavWwOkjjIbLW/x7Xk/nrTpllZpHcI2ZlKJAQJYke9PknvHGcgvQ+tTBYt11g7
2oYYDYQYh+swnJZcWwC13DBTXqlcK5b2DPZrEXYf6YtpInr/MKmAp0N93Hf12C6F
MM3PNv2IjdQDDkhQKVDD2VoGj8nVr+vPtrFmqAjqmcmjGf0K8aRlntJCUgExHCd+
51L6zr0A+vuyyTE++owhUi+U7fNqWUfu4XqVTTwEjV962BJCtr8qstgBF6/j5SMc
0k74kvZ4eqGLwg3MOAmd1SD015+C6AQJN52u2+IJ7FpRysh4YSP0mACaZbpjzi6Z
lHfRq/3RdxtlMhEd7OH4ipWhSFHoZNKH/z8x6/u99K+/o97b/n73KJa3pO9jZ7vO
AkJzZeq8J8raFhGnCZUytC9HsdnvUAymokhD95fnpLPZDMFLmoVtY6JCIHN+kwhX
qOHOQqXUwwkl8G1XiUR9JDbENVv3GherOEMxvBSt+G2JUTSObcUKOt/xkoiLgcNj
n+SNnwnDw16LJuc+31dueUHUv8Pnap8PLP1TfOwnOSI6RsPsibaGkFJGTKZNgIFv
kl17mu30Mytf7yfte1qk8S522Sc/HZ6hQkc1q+5JxPaycTZjPzNzFGr+v4rS0ECh
aaLiuRqavgHiNJbFpMitr1FCuG3lHeEZuImBsWMA8ihCRmQgD5l2RzWw4hRyY7/z
edge+EZ+/WOyghB2KP9OOzEByfm+jy1/H0xyBJNEfR+kl0z881IxbPtHR8jEUXvA
+TImchNH7hkzBYc+2Aslfya4HlyWBPxRDn/Y5hhAzw0ym50pOKXO3HA6MujhRhjz
RCMFDdtDOOOp3THhvmt02YmBGLVB6PQpBEjTVmBaQU2kBuOGvGQQiFf79alZGKO5
kZEJitgkS0GFyNsMKS/vsY0LTb/if9+6xFs97GChIPZrqZ1fXkIyhlPYKlq+xqed
TzIQSS2fG1hGsSuZ9VBEeb0Z6qXDSQai7motQR5gyOu/k89zybhQX/CXUZuH8BZ+
o7eebut4Gwgv9GlWtwQMFLwqoWuBwtmDYVLTjrRyikSfpRNd4wcMghYgE7U9bg8G
MPfZYcBjq3pj2n2NWjas7/kF5kpwKJnF47tk1k4fIa48jTz+fuwbzH6RuJ2qmLCk
TNCP9+atU0LNcjYIxDFZm1qv7tLHtog0fssHh1jDoIOifbtoRk15QZCRRO1kFRpA
qreAXACJ2oq7WheqP1JqPOUlDWx9fQo9YbK8JxasKH+wOfGiOtFBSyDVjMaA3sIB
PfZifYlMKcbsKDMtv7YuVwP5Ay+HmRmPqex16zal39OZKrFZhlbotxgYlNwJaU6s
by5dTU/txCuav0/RwAnNlnFnOhwKN6j4G/0A+v+CoJK/akq7O9ZO53fAGhmS08Wd
rE39PdSsF63AeIpnyJALgeBSNNS2z0kzdfZwe+XoiqUV6mkdR174Ljh4NK+sBNoc
ITX/Kge5l1GInWXbWo3p7MY8tHa5wh+21N2TK+v5iUNzhpHIN4Lm5WMOJ9HYkc5H
efqZjdamwcMln6LfSRpZKC1Y8LuMRJbh5L+BdBhGo0DXWYZDQm6hqHy3GknN/TCs
1zEPyt8DJcuLWfw0sqSBeEkDkcWBozbzAelBic/bcG9yeWvxPM6KM0I+R8KwZY9z
twWo1AErh+Wu3QeJS0TzmI+dnL+8URCvxEeJz2yzfXpXUeRXIRYvB7eehom3UFWH
6gjlduPOlzDQCsHGI5kfODn8nlOTf42kMj/tdeacDg7xssiM9vKT+DJxThfYk5+C
AY7NxEwXRg2zquP6N233ptD18dBC/LriphbhXEcSYyJ+f18F26nZ4R1WVNRsadgm
NkjyiKB5EQEYUHjuY6W4zIMoAr6lUPEYeYCom/Xx4EgM3EkCKtKWe1y/mLrNq5zv
uqspBxA5YMRksBHosalSxEGa94SLgBWJ9w3YR4yO+gyVJK+aTHmmI/ClK0j/KIrO
mypEb/LTlp1eAobywZhl0zzGbvbEWsiW20oxmZTcAo8QptLV1VCDVr4PRrNYg4iV
Gqole+3GV7MI5SYu6nOtxDsi0/L9dAsanUvaiEpVMFu8QG+Nc1vAoLFC5FGFLGUA
GgelcW3Lzc/Yhkhe8NPyyYb8wPoxt1cuvTqHtT3OuBd6cGYwhfAco2LK1loZs8OY
paxPiFsSLypw2eOTKX4oaCrKV6R6pEbdN5fohlDAC5eoXWxJ9MmLh/WnCKRPsXO+
0u7fSVaNhGBtHIQRqpXXeIExG6KNNcQ1uQl5CkXyfxyPeghggfymhYn5A+A3u8uu
u9OTfbunyqdosx4jaJTuZ2bpVJBUi7j7sUjk0q1iy4UYqQR7OCGh+ieYE43SYla7
mg6R8SX/dbgAJTX/Cm5fGoNyGMsRoSTzf3PDLAjrgAQeVmptC6ZEDt39BBFlosE9
y1fTsVDG6vKyUpF8g3vaCpufIYcMBvUdQETW0Pa37ubUdAvGN578XQmLTzT2EJJD
5v1IpZRssjBxMyIn6YtGXRIDZl/8wcq/S8Dy+4xdEAMd0njnGEgMmE6LynXS1Div
GhnTt+qv21KhdLBDtmxfxZrCBdtMrjSnXljE1EC7WCegJW1YSGK/hkURmi5kgHhK
LUQTRr2r2pY0N97QzuJ+jHbbypCblURCOYRF8EtV1/Q02U2fUCL8pipjf7zPuyMT
GujygBghieo+4CLKtSliyQdcxqJpdPuJRy+kvTnQ5s9ob8Z+Z3OkEW9xKqPayLTm
mNOyK0TH3YM7B2HLjDzAJPpdZ+66ev8edeVckG3HEoy//ER+bH9yj40XsENDxL79
t/sed9oLIbrKGxhRz9QgEvl/gDao6Qv7fCYG1d0RVwhBpev2E33nRD9DYsJYQfU8
QWjm4FvArv0HrM4JqOigvoVJzx+b4tF24tq3wmC5jfBiGpdBBr222ID2prishzP7
yJOnZfN7O7kMP+F7r+MpN1QgPzrOiJohkrfOdIlF3HLoykIMmyt0pZEYw8qRnGHz
P08xCp9X8+ZI2Rrjhy5ZN4NjoWKvTfJ9FkyqvMPair4L6KDKH1XdaGhmmgxqYKdt
8lGggFtgooJxVbSc3WAjQDawaqysgjn+Gog7Oxk4yLZcGRYWznKY1Yh+KDpJ0o0D
SynbK9PKn41II5U75GBN3E9RwRN8Yoe20/RH2x575crlvXs2ygoTFwC9p0NfDWli
39vWcFrMvd7mB0TWbKG+wJ0SuqBuMbq15QXeXz1iE12N4txmO0k7L/2GJS4SVHie
oWHw0qEyGyfI5lYabrhCI4FAsA+EvXwYO75Rw5Su4Aj0RM2A/gsjMBR/X3LKp8nz
Mv4sKkqOuW6qq9CnEtto+UA8C0/fvhoMtJ+7TFL6hCM7fVR45JpkFKual5oTxiKh
6wo5OkYOlogLmNKxvhA8G8c2dSjRfisR3Uawd7PSjHRnNlUEwCEmE50irsPsYWCG
ksLRfWNyeDsPNrpuEda617wFkyr872gEsbGMc1LogsE/5oGi3NvPDXNxZOiYAqNa
SmiH/s2POtwGefTq9h4EDrTFj1aRAz9cNO8MKitscokJjJ485ENirKUH5jVxGzRA
hnpU878Tny4HIQpfbHL9Wfw0V+vwuttC7VFVjHgRwWRp5yy6IwkL6A55RrpQvM/t
hvN4Cc0pYg6dmCmbU6WywUsAawvNa6OYyJn/O9kBJs/uXu5dmcu5P/IZzH01toWq
54k7PhJBrJIrrahJ96dkRzHVhnIy2enF7Br4CvcWDdmePnEx6nBuxdHL5vNBq0je
+Nb+H/8ky5JiQUvf76GtHQswqMQUCevdv9LLMTongcU47ada69j1gjJTt8E2aD0I
JbPBVAY6wgKXI/BDtKAqNL0K9mF69bJb/Ba0a3nisTmCZL7Kev7Rt2dRMLzW3q3z
WLDzmVtc9T+2DZQT2wIMXb6DUFQTEafsgy1O7rEMdHBrJnf8IABJqllbvdMollcI
sUfXdYzonq1uVCcDyi+1lo2398u9d8OVql3p3lNiIc2QBy25t3ChdmGZbvpjZm0K
G0Zpa48UxKntztXtce+pTNRiYeAYgxtHokv+CXRrSXdi1L3v+VgMzwgu8SLiAQTh
pxilN7o6NPs65kpeQf5wkCBdJtwLG8GtpoJoOGamXI4OAo2J8Ua/GyauZUfIJZTx
6JLtdNKXCrJjaw6gbd4g4QQ5Xy3w7D+t0HcWPGmSqTsMIcIa4fzlsBbUVujPMywV
gXRIaVEiS4QFbdKoZyw/QE8vTB+6Q/5ciy6j8uI0fV+fRBicaZIJTEQ6AyZcNVD/
yG9jR9gyl0DwbadTjmelRUVJUgdKHczuULwV2Ont+i1EwNJbpSlZsgY4v+lyGZpp
//rZuUIKhtuHDgOyBY40YTS3ULZl5GTdxrRaM5KFJIP2O8IUGw4J3nZYdtarBT3G
rQB0h1mCIx2mSHHI7lS1d2T2l0nrG/Worye0WZy0clIlRsjb4zOEmicB+exxkA6/
WsbiXoUXz3yYQQwjR8eVKCRCxgmBvpHUPTLaN50d/xOPVzGJNtN15l+nSn9mHWDa
Que90ju4LJNiT7jsJvAXavwMOjvh5BdOEz7n8cVveCkD0+p/yrJ1Xfc7aFgrTmsf
jDPjmqdKkWfUuiFTAZHuVGN1HIkYvHKHqUmOMRi+v4NiG3nXg2FgnxUq4FEh+iIk
5acEGdj7hbvHsbrlh5qbJXjYA47bvbX6NMrATelvtS9G07DhEf+7CEKFdjtiNfYR
j68LmBREfucuIhWG8EpnreJ7ouibQQBqWpJzZ9AP/SKMdlsRiEixY34AJifdMgTF
38AiHt84qbn1rQYyAVeN8owUAarsfHdhY2CV0BHGejw34Qxras9kx1efGuyu+T9Y
gktvGXZClVPJWtaBPggDYl5IEXXL5Q9SSM/HnMDWR94zKIQF3PrIK7Amj4iBXArP
ugkuK1vJiBdwXlQaD9Fet6xPiRZX9NlujA082MckpNZNULWtoC5hBwL1TRZm2++h
45sJ6tPwbFblJlyGD1nRQy+F0ivqkmehavydyI2l8bc6neYIf8jJyLaRH1tvBLFa
pKKawGUebT7ySJ3QPagnjbHHoGqTJ78D46f/5nK7ATFfzGDjOFQNYR+9ZbVrq7oT
NL2NtGerdjpWkFfniTLAwsggBBwFkolF8TMSNEF8vwyDlo7bk0bBK1fdUHHZXccs
GpEfQbxwP7dGcX7Ba0MBoO4DGM4PM3zB4SkWaCXpyPvXk4bwUIeOZerKwGhecF4x
kk2/2Hyo5LeW307RcaPMXk3ivauh/kk9P9cEYd9V+WvY+rG9QhCHy3+iv3opVxXS
5wH2DHzewGHxgB3mNh4JKSYII+BWtz78yzyI4iePmvmLUA5J7ZSCXNv2pcLe7SL7
fhWuxoFLd1hSlHiJ/eGY/KUB7jp11xPynDUmZ4/wUwHXYIqjQfZ/ifBplA1TzsUN
8ku5f2ymqyuUmfMWBPbamUi3rzWM/TcR3dTWrO06I7u802CQmOd213shuryixGli
UlVhrHEjJJrU0Hvbiy3fijD2qQxhRWJJHVdPj1XV8ldeM0hN5hvlPVSBRZANVMjw
CbIHf2SmMbgfuHZyUqqS/liSlWd/0a0bmuKdjnkzS/1nLEmAllFWab4V/DpZ/4/J
95fC9MDQuv/Xx82VAgj5MFtNFhFNtdCmCcPh9lWVOJ0DL/rclD4A6Kx+oyLmBkis
IHZjB71zcejDmj4l24drBFdtzTtdaNZWPA9IlcaCNtxoZuPDS1YTB78p1zDsGlUm
SiRJ7nwnJj0fM3KBrcw9ddLm5HIkVaAFYA7Lo349Db8DpbAysPbDni1ODioMmh3v
d9dMx22z/QOG6b2IlYq6lt0YKdvpZdLfH1nvypOuR1fxe0Y1qhsWDyd4c5wffKZn
O1toXh2wZyfd1oNl3DMadLosMn124oHgBhgSdN+nP6VjAK4TGvC3MfkB8Te2jo1K
1roIFP40utr6tJTf1h072CwpVn/ne1S04r4g/lCd3opdlB3DTnrGrS2BKAsw1WVH
0ZTMcZMYmXNptnpPCYFFYMPBaiE/OBlkTIkq0Zf2MVVOXhB34S1UBkYB1ln2Vc2Q
NZcBLr6Ww2hJTENSmpYbj7jRweA81zFSXKMgvrpg3rRVY3+8kRZEqphoa3qwoNki
FFBqnQHJtrjWCxgHTBLSqet7awhatgyQLUSUdb2UdBvAt9uZUDrF8dAorcuaHlYF
SpF2HIgJHYSz0n6WJv6jNmHTsq525Bc92cGd1gdKy1pCNmlT6CTA44+N4LS6HTKB
IVHlhO9EQfyRYjshZz43SApmoj3EjKNnZia5/v9HbIYSro0OXLgis8ZHq6QOQMPA
Rfjx85rjV3N9RJoMoo1296kxkaQU0qgXaSJYzTHOeaFjUt2PLni8342lK4/Tlti1
BcY7FHod9B6EBAo9Axo730hjIM0oJD01FZPdXB4bBTZ3tCwOfR/uA3fZ8cdGHbes
JHqicWEnx0yHhYEw3NYOkU0gY3a/mNvXXbbLhjJnp8vEX86KutGcWOBB7dpM1PnV
NKm3TLVERvZLSYsmC+vbSFRW4JABvtl9Hk2Ij66zQ6aXh5ftbol1GY+OojwURmxu
hgQsNv7RCUGI4X8kFi2qCbdByl3sb8HrxEykeb/sjEz0xuJfDjgNXCLFTJnXZzuv
ZQJwipE8lAfLQmDCM9B7077ha/SB0gzQRtdnm75CVB7oZmKIAtHSKUdPZ3ZuFgs+
G99GRS2ziFk6dGKgk63dRs+L81SJ8sl06EevL9Ggn804AEB4EVA2bwkj01SAs+o+
6okc0Co/5ESaM6WLMAqlq2VTw0ejT64G6lDl1mWWsuTZUg0Vu9zCl6KviPJ9/ral
CGOrXRNUEFTTs1h++h71nKhnMcZEWYRGlDNCLm/mE6GeyrMs0LLyYem5ewN0YWHC
JPbY4/tEj6eGV0f6i4cHovWJPc5RzxyvmPYijP1MbaavyFII3CCaxS7juTwqtb6y
b6GelevPOnBl5fEQYj/prbWAJimAVETHnS44DAtdF43KtHnDmOD+PBG+/laU5JJW
L5eVuiB5KuwiX6L/M6rhUo54YbhNo2HEoD3KGcXCQAye1efsF6ROeMj7SGK3uq6C
7skbLH7K0igkDmpIe2emd0TWUZE6eoiKCP7jXzmNi9mJStnw+yT0/uCXxxMcX55s
Z9SSN+1dBtJkAptuOzNRTNKc/e15amZyjiL4Yy/vquavGRLVLzgP8yIQ2/m01MPK
Ih/aB0Syh0qAoQgj1ebUGVRL6oCTRCR+V6H6ime/vb5JIzs7+/EjxFpKsL00s45V
ikegBVRZHfDLHpPo+za2l7EOcokBGlzlOzCwVbSq9FeYhxM94XaZN6E+FaDwGOe2
T4XbD2rKJzeZNknetoD1OYPwCJpNGsUYA7sMhodDuAvUmbTSOYXRyiG85cVvi+Pk
L+eDJb+1shYsTte4pitIp26iqZ7cdqNqQLogrPx7fy5H/PhKEg9gksdXdRMIliXu
JkjYScjru7rh7tZeKyFeXBJu4F5VIRWcprOzrffS0+K5se1DeKBunVAvZ2cv0bpZ
Tzaxa5ADTfhDpX8OgEH4TXoH8GEB8sH3GZa5Cygx7WC/PFIovcLez4QKYFpCaR6O
DTRnQBIGTn2FO7GKmFqkdF/kCLU21lI0mSMwqbcUJSNccQ3kO5dqnd9+/j5bSt1F
JHrY9cpfDQBKatv82r5q4FdnEUASUe1IKqgdpmhmN7rPzy8y2JtlBMExyag+ll1C
xxsqLZi6Tgb5T2GWbGpOJCZt/O6EYHY5Tp2lxihRw1WpOYauMFmdUVvy72sBrceY
nVTICW8VLg8i6aVILtsJns7D3kozvJ437cskNYNFBiPwhSAfwSKZclb+IXccUbR+
v+uEXm+kt3htpnFtgbUW1HPJLeJCnViz8SROST0zlkjvuYzHLqXA0xYvBMknfL37
q4T+J9Rw+GIb1LGmdk0y0Gp9u38WVp1i0ZqhWaWCDltE/82JPWsSIIi4+iYnFgeI
amSIOLkOENrXe7z21pAbZ2LLPFj0bSJRLnRjfz5gUtxNyc3JW6Ttxf74vYMY6Oze
utQdPq8efg/zKcWd03Zcz8RWX5nWEfx8bCBhJJK5rOzQiGiyjA+D82qGGPZ9yx9o
T//Qe5wF4uYLYyccb8LF95VlvfPM/fRnADmmussGtKuDBuxXWUfcaerzyxF06fNt
DU6uF68QtQUtODfJ9ssw38Llm7IEkteV4rGCySmASGTz1vs8OBdBSniwnLqW+9qP
9UmA2t7aatLqK4wQU/mphn8RXFFCBd5S51uwURNdIQCsSINVOR1lKQcdoPIpro19
Eef8Md8mZwpeiDYzewZ6K6GsQHNvGPDFSV9USWD8Pgo14ITKVe/ssynLNvjDw+kP
LMQ21UXitEv+gWKKV96G05J7BFm/hLn2HU7xrcyvSmmbi4xicl2RWGaOU/0fOq1Q
yKNsJLyUK+N9e0Vn/HLK80QG4FLOsnMPweQu4QaBbnNT3RN9/0b5P2Rj4ZI7Ef2G
WVoru8fGHhUFrkfgkG9AyKfrLa/2y7LBLhssE1Sg3PZJSy+Apy2vEtDgvyl03XZu
7LPtcri4M1KKE+tx8lR+SCkIMSSrjT5xud1lIKjPxA2FYgW/+wnRFslAuenN6aG4
bF1GtQpV3P5FEvMUUgYSfgBMrzCj0yKw1f8rANAECddBzcq9KNBycl1cOj7BB1HZ
3anBk/YR/pyWUmI1OkOBm4GltJCPzDQN6thhsfbgH9SzWGFb/5IQULPaPABGlJ3s
Kmk0n+yP3DRoIMnTj+AmOdwrPD+cm28thkB4p7P4LH3pgCH2w9+BlbZojqAKEnV4
gAmY55AD6325pQ2M5YQUYh2YzVnCIROYth47AWGuJAQ5Klk1++349Yff5DbAXFkl
Nm99SS7Ez70sehcDLWMbi4l6PuGiFF1/soxuo+3bH5+FiiFRxYBUXzuqbubqbKby
0BAnCJdNHM1JrksClDQhRaYOEjOQ5PpzRscK56oPT5scX89tAbzR7LjeHvYftdZV
gX06dCEg5CuILPICUKY0LsK9Ln7cXHNOnVAiUypf4t7dDpZpRzeWDIqoXUPNvLK/
JMdNFDsAuE5xEKUGaTLJa/RLzKrWMu/NTLuZvUEFIDXkuCWyI9QB4liZCKucWvPP
S2hTVy/fTl/2F3SeNXcb3bGkCCKpS8j0r6ns4pcKTVtvzdnPHuNAkCT4l/zWpRah
vcvRqHXigsAWsdHMgjSdRzR5+onqMc7TkgUdtPuKppMEvuBYejQVpgcAMje5WwRr
PXRVzll3volQmpTMbbu6lXuiSz3zheXQB0Tt4ExdEKoFznYMkPhmzxoWr/MyHo7A
TXbMUpUfeEIjnfV3KN07xscWYrH+e11R6GLoLYNca0AF7KnPKshPkBf+1GXiHW49
/XfCHPWIkibiONBqIv5cxnNSF9Sshg781iQ0ca9RPBkgVU1BRoFl6xn5TQxfDguS
eFeeGXPrmGT+CO8tYN4yeoKcY2g9jRau9qScsFxtbyTHO5M+CT3RDeEgY2g47Nvi
Ff6bp0Y2Ed7H41ok8yfAEFr2fIPrT8lZgXxFzoDu9lIHXZ+Iq7GeP/FnkQGsurat
vo239s2zOplHtGRCM+oIPqrIbLpAs0NSPikjGqH8JwFS0nFYOsIF3gYUviaCVrfS
n+5v9e5SSvLDbCSoAntWDaeYNj/ndUwU30O1UhJ0Im38dQqOv1YNv1NrSzr7+hcT
ZzR5g7xP4g9JQcnJnMlq0zdXQ/ldbSBNKY99TWmRUGeBHGO8akve/T1VX9dLoGKO
KCXVFVoBCPqs+wobrCYuZm2mC/icQlFKN6hDpdYL/A46jXD/uazJK67xwjxk28M+
O9KUCxZkixOwTg+httEjM/FARApjQDtITwQ8G75BHfLvOZuVyKrnr/ZmO5nFEtf9
w17Rp/QOuVFYjN6e2ghG6NtKz6IuJlTkuRu1O46D289y8/hRJJhF4u5kiOoItLm+
MXi9C/XeERIvkeDqtRVUWFf8s0taEQg4YVxSS/RH4N2Pnc5pXYw4z6jTA7fbJgkb
+7V4yR7sQpv338msJHgg0M6JNG7/ZqZ9MujcJX9fzvc9y/jSJMj4md1H3zJAwc4V
LuGplx81kal2mfL6crG9+8cURSwyi/siY2ZiwixUxUGnLqV2pZIIGR4nPzjBvB4o
n60BIqEREfKPhPotOrWGMfJVFlU3+83uPxelu7hCuVq+iQI4NS033m1wh8UyLViW
b1wj2YCFtnG+PZfMK9vgd1162GGR9EKNObusFYRLLEvnafZKdX2VxT8czLMnjKie
oIzNVauQ5JXvxK3FCA4NIRr5/XLMlKWAvUxmsbOBFw6BR1dAkT4WsmC79yjqpuT7
xes0664Anv9TVSuMDsFpU4qKzWlmAuBb9FMkPCt4ubFhDlenDHq9/JgWr9K0pMF+
xMiAhkFZLc1g6+mgF3tBGxG5c15FjNTgy5gZAj8APedR1A28GwoktiRUPvIxcZ4F
AB3Pp7P9FM9n6sxY6GmzAI4gnvzP+P9OdK1n1elWZDWvGMpfbphcKrRhezt4eiz2
JN3mXlmg46LR8cN2bCKievpeUVnPZ50DBVwtpZ4AdLn7fQtnLljaagT++zq0xjNh
q6HICkcdD31siUjPfYAVOQ+m7zM8udPEdpEZyaVYK/r20C5AHXLG9FMNNzpwERl6
lF9ddjX+DQ8Ws6AaJVLaieXSqhdab00bLivfpzyUFNHI8BUPqun4yuFJs5j1NjIu
BMOa+QLzfTNt6NH4LvX8r0AsROjmGKr3udvxm8B8dUCwkL84XTFZdD1MVT9IcHLr
jMGvZe5mw4Ier4UrO8ipIzYyqNAGQ9r9ptvrrRx7VrkHLHoGn4i4NaDyUU2ExyNl
gSTiVLXJCwpUK0Ap2HOgpKQPtBpPHRb472t2Z21DhC90LO3eUVQRPMdGUR+L/e6b
wPI6NlB5CCh+k0Rspay7req3Nl8QhQa9eH24/RVN1Ep/0z7zOz0PvDb+YjgpcOiC
TzMJcorw7VMkDG90mtB2XR8jqjs/oCZageZrn7HWRkrtjT4FqFnbcAeyhLxwUtCR
uIqSrH7qIWtxXgvSjhl5rOmuBJQcAmmKIVP3/LO+S7rodrBsnMNt5r+0j/u/XQAV
jAvjqCI5TpeT1PnCfb4sPevK55WTxHxZtMkM1tPf50GiaXaEalOzEQn1bVBWsCcw
dBI8ajdNn/DnYVB0W/NezREs1W4uuoO4nzE2pfBNT292BRuNX0i27EUSZo3FuhS2
GeoMNPpsxAdUm7K3h2E41+Q9Dl53Lry8LwDX2QrucE02ok7O7pe7EdbWcFnrMIbP
jeeTPZThI+Cs16IozPtNMl9Sv+xoF/qtUc5nrhr3vqpwnw/CjKKRZezifeIyvb8Z
fdEHS0h9T6gn2OFg1J7kAmN9UAEhFmh9aGZIX2CF+Nyp8FATuUypEziuRHV/kuup
sI1ygEvHd4MhWDijhkI8AFH98ZQYS2y9VRnR3nUeY6KIuoIbd/nuYDqdD1Vy05fV
/Y68Pz+S2wmNLW6/gX9ueUj7MB2LC2lz0uH/hvQtj20j51R8E4Z9/rrVBQb1JfVu
Xv1815A8fNzQBCvZHPw5ztvA6zjLIyuS0lHzybYGPkOsqcbz2frVwJ+gXkyXDjpE
60+nUhPULlgzT9+j7pIYlLvwfLD++V1iGQz5omU97Bm5T1UFzPVak+qfAN8Eq58K
C6QxiJaG06KXXmpNGH6fuBMi8eLhVq6D/iwc9ICH2EZlwl+3ca1oBWLOQ6jcWcNI
GgKqp6G/nQX2ET69TKdIt5xXFwZTAffDyruvTR4hFlNumpapolZw6FhjsEgbpEqq
jFm6kXvRCu5BaZF2SCAIckIcl9gr8lZFhhzyouwbgoYVNq2FWFTpoua+LQyPUvjq
YglO76gvkkeT2iJRh5N6ESU2uZJCOGYF0dX2bEN0vLOiTgOhiN33XJA6jgr59iPA
IbtZgWD1PPGzFFYSOEQ24ANGzC5bkEFQBnpKZT8Dd42YcxUQB5W/iABie/qNawVE
vlDsL8J6c5QQN+I1XgbxKJKMzPITQnzJH0HcZJ6f5+zSweN37JG1lS/+41vtEClw
mNpQ0tsT8eu/Ls56DzJArsDU8sSj4h1HOzORxPb+hcm8dxzQYVmgduu7MooA8vA5
K/qOOu4uvfqiX3xTjBDJD2LAT6ViCLCBR5IHVdgH9T6KiAzfhco4gS0w18JtCm81
n59Yzu8I7z0ATu18KHlYn51QTE5zUvR4SMnrB8WdNLDObs54Y8BGqEg0zoVslktQ
aV8fyrEnp5fxkCf0SWOqYV+8lxlRezEXpOGES8kzPOquzoRrgdSrc1pokiReD69q
68U8HDuY1wNooAdYjkhnVmaZhn0Vg+yesJhDOs76o5Z9JasfdjNYEl5CWgQI97Nm
M/cVD94dkBU4K/FwBDFjwvf09W2f9WSwDHWdd0M43L2RkVGFXz4w1bg8lDZCmIfl
TMuu7b9KMO6siuwhw0TV0+Wdoiw3JCCH4hPDR7tOb8lUMq2XxczWe6oFAAd9h/cG
ZmfVIwXIqfj2tgWfu6syjaiCbS5egmQCsmca3JisdIjBbJn5JX5RrW3aHnZotFSl
Sca4+a0uPEYwnvbXYFoujiKwa391DhELrnsqpekF4xNUB9vDnmcUYqdX9hof/kr6
7KGVMI2HbdMciDYr3uZlebHZqGun6tdUwmtCEa/ZRB52UhG8w+/4Fyrd5djcxI0u
eDDbyAKtroOGzcR8aDMQEZIl7Fv6OEzXr86CmhmFDzqmAUrgkhDcPvwr7c6BZoxs
PdujeVBKT3hryGimLwNDuiIV5M/8mhfgPmzBp0pTY96IIpwegqBeMNV+Jaop2R+W
Ux/o+lpPFBGScZ68M/ZqBWy0usiZc6qOv2YtIjXYnQtZR+qEJjIwPe02yJo6g+hB
0DaD/xRFPTxN2TCP7bdZ9fp2uCWGy5mrwZJyZkKiCN3x7gVcpBL8E3pM4OtCCQtK
GIok/rx4iGTRxYYulN9i2fOwJmhAGhLvdwAX5sv30zYBVy2w5nLTrRad/0XkSPI3
kr/Gmjd0YXDXjLWgAawuQiUfl3GPZ+7Li4s2YHb1fzjxWuQQhq/w26/COGEhSdX1
pdd5SGBqXJaMB8l7msV9IS0JmHKso37cWYLgqT46OU3Peh1a3zcdtWsVeWG/Jczi
7rz4QsHRXClVEv9JIzT1itEWY/3vff4KCyXEbt9BzTfFf3/gopQDhA0e1GqRq4cV
CzV3X8NQ5vXznt+vmZCbGyve4JUIPI8wT7YTaKXpYgnfc2AMdi/TOTkwLuMW8Ndo
FiQBLXj5Dvupn0SdVRl9jUtcJEaOLDfQk39fXGTBwW9SlcR2GpGeazWWX3NUwEY3
DexXhd6wECX75AjX6G2QSqAYE3U74MFRJba9qJlautWcJ8yul46B02kzb/FAA2Wx
iKKUERvR4Zoy9iDdOsYt+5UY+mjuHAayVEuOZ21NYurpK4LTIJHGWBudPS2zzMDq
/t2KbFa7rMrcBsAYWebnWzFZr6mhMAMILqMGj/wwqXP3r2NLsHWdt2OtwRTdJ6zA
UuH+Y+z2vLA5dVGATpZonJZbIWlREpFiDJfYUWrOyVzpaznuiCST+OtX6+a4VnL+
FoOcP9V0M4FVKLtjDQHebZpIH48eKmyO3wVIcgtfYhObdqo9PVdXPnW2ymFKabZi
qSeZKlFeAhA1sgadzH5UUIbZrJ8pXC56kenuw07CYRNHskvKqRF2VP7HYhw+hL75
i2ET9E96cm+/rF/EAxWytZGNTbNWtYmOMONzJOttej1dPRl2YrfTlM4lYAUBgeNY
ums41jyk30fVmpUBuz0ZIloHnEw5MatbTvmrM0I/vBTSSgRCAGvdMPIbG7OFjU6f
47VOcwUd8uYra+Cfq6c14EfWRedOPU6aw0B+ilAxeCfBqDbtNw89zCXW7REJRVaB
lRuqIvBjM0cjPTDxSD9060OBuhZ0jCNye5qgQMb4WW9ZPSkymV0k4gdqquT2xz0L
q7aqqg6VAzA0PwijRGVFheZ3t11ze7zi5dwQkkrLA0KnjvVtL4mRdictYXlErfrJ
Y6BfOKGLjZY+x1lAmxveIiwEDlVr5t8rGxlrXzNARI7pO9wlMkfkFRtz/HZKfVX2
HWSKNWFJ9zVB0nHSVgzbDYEfw5O+U9XLBCH18lgZBdUonx9r6w7uvGOTNJ70eADy
mZGIytfgihb3A1294uLecq+3Mp0IJwB1VAbkh/uMt37ILGNuwoH2c2xSBYv/IW9P
qpb9wANfHbG7KckfO9oWvHGc69bXKC3yCR3OnBKWMR1AUQnS7Pcz6LqmHyR/PR7v
EHC0Et/EG8oEzja7z3rl6opGavDNxBMB2YBMDjGOPLsHTIaCgRTbClP/w7XWnCZ2
Z4hKXFejjTlStw4V6eKbg29TK82+bhpIdWbJasvsd+UDFoNNlT2OtIAcjrinW1Tt
2sx2TaL5BoAfBqRI/nE6+pxnxDrMNZPeLi2RoADgvDV365YfAPfNzgtNNl6Mi5+5
IWMYYGazGXjfIrWgUF3r2AwRI0vWlQmr4vNM1c6SeRli3lJ9lmagodCCSfN1Tajo
tsx0bMFfRBehKhl/w9K77Afm3jIP3/ewgE0PXN52rlQe5Nb8ENZWqIOplMPM6/6/
IBPDGb/uJXg4blL11Ww1ZsIZ4bnfaDkyXMU3R8Nc9Xltc2t0MTrHH5/D266vCJCp
Vb2XH+YT/tpnUA5LqCRvt2tD64zVMKXBHDa8qR5yPfIkioBXSLM/Ey3U05KQQNj0
0UsPGLYwfdKbQNT/hqtdiZvFCd7LMA2g6f7A11iNZAxG1q3nZrD/+G8eUIIcBgEL
dtwM9n+9yB+B9B7zxd9PyYEKgze0FDaTuXrzqku/LNaibRnyQ8GuuBAm9YLiL/Mt
FD744eQ35XYyHGv+1vCu/gM+h+ugwNKjBRCtXkon/vIfo/L00SZGbBpEUSEQLlXI
2qUkUthnfxG7L2ROlh+7zq6ZOmT/q/LF8Z3AlPAIEeYcDAzViEDM2SkJMh3XoW0X
Pfus1/luQ80tEx8ZvH9ypEVL+fhE3oMdeytEpn3NEjuS8tqjkdYhRtTep9hOwSAi
e3QIwnoVDGWQW3jmT+0uFuT+Sjj/TgZDaJqbIt4CcgS/5glGeAOTb4Jg9J6Kwf/S
6yHmz153N9AyWP5KJebHl7gOdjHub46hxrX2+oIAMJd8e/mClqwcPwgAPBpReVPD
roNggceyvk9jiNfE8dtAQcF97l8mSdnug8A49kmMVRHIRcRQZ/U+sVBJtHqcGcNv
lKLLjf/3k6CCrCq3L9upLFX+0ezD9nUS+iWm955PkPma0ni16c5JKPzyY7bWxPsA
KUb8IZUpXsQec58496YsPsHuj1+VJE6Zy4wJzI870B3f6r2dHSGoHXLEw5mybIBf
M8VB0lLufpLbWA+VlvNka7iiD/nWaVbsAc88VBfFzqPcaNEALrVTHpHli6ZZxQ3A
sEYFwyHmfNrouWDiUfEmCukHqObS0qVzsWUXiDhOo7egXtRww18ODI3ylhT+6LvH
LDGgsfpQbs23FSyzGtVLydwR8f5o6bswPxo/QW+bKZfIzS8wJnZZlssxqW+qkgkZ
DFG0YnGmt4SXttebHFywgkWYbfH+yp4mu2bT7wShx+P+PW0nwpUA+J7eqNWNlVTi
J0Cm2XotXA7QdY83u1BEc8aQe6L5+31zUCwSMOrS3+k6LMNDhIbdYG8bc0GI+sIv
5hUBc8+xXZp/BqMwCCyD5Nr1KQrQMxQzAf4HOFLqJQGeKopLuSYlyQw+X8eKJKSj
pIy1Jh1BlqpHWgAHIM1IA5QwYqVAKAaQN/os0rbTT+1fJI6o/fM788UV69ely9qP
5QJVLBGQT6VZDWKkF9f6zD1yPIgjMoFYYR+IZ4GdiO5p2932sc7PN2X6uKB4fmPF
YeCOpepzavUnn9WO4HpS3l0W02TKHO3kHLCLqE7yVqT9p7/sS4MeXPnGTkxK9Se0
bjkttNPGS/CRjnItuR7/PsKeN61RDZxpp1AqtVlo+dSlqyvtnnKfTLSIr1xtSCoT
AokEEcYsoYEZWbRyy1GLFfFzjjNZ4A7kPdUGicrYJNmsAo2bk4Zf88NLsAkOXPSb
ZYrMNwc9a4xYgpnhkWqLWltZmITYrdNtxMdNTwTeSJ5DvFHxb/EG2gdCmRzuJGU8
+cubLNbzLXYKIpFpI/DNqPdzUtgP2FlZlGpvw6Jr+zTjhs/fe79xrNd/WDRz5oBJ
M8qo19O8BWCAPZ6TvcqA8Ryop2tQM4t9jvpOSjd7g/Qq2LX1y5la6d0Lp6S/lO76
Bn34hI80jCxRBJSgOzJe6GLc5Y+KBKS18MafqO4KI7lkbE2sBrXdKGqSwBqQmvrO
UPQXJJa5WTww75IDFZZPy2te9FhOHcOInoDs0vMSnbioBVHRuA9ksjHYmZv5PzUt
E3bhI7qBVgsWVCCtr0DYXY7sPp6/luW2NWRLa/WhJE9BMs+6zuByf+2upkcTvFSg
fMwV3EP2/la1rLe2a/9qXt84UvVKLy6+20t1VogLKezogJLooITkIp5yh4jfwNgi
zGUAi2NKoP1Lt8VCHsZHC5OVMJxvYkhoOcO1uAGI4kNIo4SIYXBKcdxMRzN4cNEI
j4ZlphTPTnWVzVBtavPzVXke4S/z/8s8pd+lmp/iuYWmFE58vF7PlaB9vYTOQrZQ
Dq+hByKoevpBNB1okHKGwli9rXmSG42eHw955GGpHHd+jHCOEiP7kTYdJoVHc6Hg
mNdyJy5i58dPKkTcp6d15ef3j5RNySbpxHlodecZnMiCJXPf49diw/ouP8vBNpks
aIEN4nL0LETc2o8BcgMDIW62aNe8cpExE+4CRqqcvs+fgr47kCXF17ZjkP0ONOWe
BQAaYvwfxt+rQaDu8MUhQOJk8UeRki/9hgHvAGyGze394O0CHZJBEqX603U7hpMb
a71dWdpHMV74V+bQbyuvdeSs51Fa8sCfQV3sOtoHpqytL99ER/tOSONgzJH9EbBx
KbTGPSjqhhb7UcQk1rZy15rWRPBjTVXRSh1XB4I/vWmcF5ajd2LX+CI4bt2gW0mw
z+3tF62iHfFqUQk3gz00lqzwj2CfoOC7brO/qpKTJmS1FOjKgvZ5losey6ntpnEn
a/EeRbX+WZXJCZpuCHa49q4RraA4EoooZUeJFloDi/XVmcJ1udx6SY8wxjQISj4k
/ZjfjFbBmof7cp2OWbM950YfxWByR9dJLLqzOWkCAG3udfH94vI3vTp3fOOBk+3u
6iYJ+ih9XONItzXgf2GWk0Zvv7nLwi4RSz8nSrcgGZ9lsMthIbnRKd15oz6ANrzN
qecf36w6Qq3ctF0N0LqVEI+aKqGwdBfvdkkCiCJdsYc4PM++4zGVWwwv3yV+Ola+
4Y6v6lm89VffghbOVWCW0cU5bBdT8wT60pAIVaIjvcVG1Bw1rz62XVfQOVFs7emp
weEXwF+DTpI7IlRBDSEJYtils51EYWeY8f9JBRZGwViQ43o7580nXJv9d5dktP/w
BdE8sl9ozkiUBwzEkjm00VJ1DVTJ+FPi0RGJurVxEMgYYE1x/lC6HprrHwFqFB2Z
zqEK5QRGAlXrhVAoO/fC+5CLyXoU1TonSYneQSI1FlFfNM/1C8BCKlpzceek1Z4U
QAF4VLkXkifoPh0QHmpxI3pXvOsqB09wx6dNeQy2oxiv+nc5gGzv2KgNUnlD8W8D
Frbio0iplR4U0c80PGiM6/lsd6SFuEoz7Z5DU6FRX4y1Ax4VI7CrTkXvaKrJPH34
4MwsOTzpo62+f4MOC2y/SMHloTglH7O90u09JJ7AzwaLP8jfmtHL8paqD5YVwhJ/
UTQvEmwS4huveedwWpU+/tMUl53rocnrD04hfRTwZEVFuRwYqjfuNayy0D17m49E
ULVAltW421Dy41NmjHDO76Hw2hH/hUlLA4bzZlzTx1azG5sCjejoHUbqrmScbL2x
Nvbv6SPGY/L/O4dfRBrDxcXWkQjVYZyYe6MBgWXOjHjfcGlmLAodGwXUkHDtG7E8
BGoCNjHb6Ls23Brc/hXbS5ZCv+KNOC5hvOnZ5BV5T1LDHn08Lh+GhW0bdVNBpcyZ
WdMw+IkmE1vjmBJGqxwwmROw+kWFfEAz6iIk0SpHFBTZhuk5qVJ/9UCC/TMrRf2B
+I1fZbhUknH19sjG4VzmU9uK75h9vVX9T9fmovlaRN/fBpOeLK9TYCBvQ8vhmAyQ
gpTyz2Wrx+dwvBB+YkCXYXp0YMCuV+yD/jMj4bdi/82tTcZbgiB8a3Qum10i9GVQ
F69posEoGNcwJqJXaqBW+P/TqjyQU52TrpfrVpUt+IPGSN+bQuCEYiv48TOUiptJ
OtLlUfARABiuo1sWvsgVdbpSoOLyZvQurDpjlPC24z1gZ6fcwrJmXfeZ1cvZbPln
yQWJyecs45yMkAqyeTaR8tN31tUuQ4TX5Uk/BLJbI+8qYgHMOosUPxkr+bHmjS+J
IyppZNEU6U99rTPCeXYaCMzNawfHTdSKeOtmosY4T+T4gqTPNop20VzD+0QxdWhQ
OgoS+yL0ZWgNMdX3+glZGwA8YNKEVoM9xBhdaJtX+a7M9esPWtEkEvaFp4hlRVZv
0v1XGVh0va5CqpEAkoQczXgNBaQmrObcepbz6cUZcvewB8ZY/fQGlpNNJhlXoC6H
mkk9AU0stHSsHYPBSd4XoTHRYYqrSJr1YL7c0OuhXhygk9CF6YZi/lTur7zyJHK8
8HrDch+KBl4cMfsqwF8ODaV6g2eThqcB1B2Nrd6EfN14Nfu+Am/g3SabLDj67OvE
IHVCtK3BVvjTx6aybNSfOc/90mGjl3MU72Q7tSxxg67xrdMY/yk3BwVdIIDsVJrg
ZzEOxikTEhZzc6EPOT8OHIYghUifAChimjGV1CaCmqaFYVBUhmzijfjDK55zO6ny
nK7z+UVtjYvITTMoI6SmfRm0QWF5NOvZ4ol3ZRVjsrZiACGxvVqMZJzR/M7gF+mz
dO7EtVrXLT5L9nVyT6H8Nx7sCKIeF1/3q3vci4gnUOIAkl/EOIxm+zHPW7r2+ZCp
rH+WGPTuTgbYyIaUy5HqAzLZjk7u9Lr9XxGsNG0pTaiBlUSHU6/BwqhRKjWL8OTg
kck3Vwcc+m0L4X6kL841ZiTJJNV9JrxSQjz2qDrnK8OxZS9g0lcfSk/lwbpfOykg
XlZXhGhEtsgb+k+juZNjWa5u5hXWYPLjPfgGfd+e8H7LW+gHnc2mTezoWBKc2M/i
QlVjptExaEnFyVAiGSw+wwZuNreoUFr9D1XI0iklVdFf9J5jc5Krpo6sZcEKbabc
igqSB83kx1uSppafttlno7barXMjv2nvQC6cpz2XlYYulN0aJikC9Hn6QBiG3laM
B37K1HWr/qWpPi8sS4iRoR/Pi+YUdsuxL38fRv9DJlxjQyhoukT/sM+3iWkFjxp1
DcIJraz7vTpH5KD3XqIY1f1st6xjE5xbafZQ+C2K3bvREAr/afj8pTkI/9vy3jQj
tR35NGKaOE9hQvASgGLkYItwG+QznIgp1Gx8D6u7ABnnNlROds3lc2KaacH4K5wH
g/9Hpwl8rmB/YYh/QKPKPMsdCltVmLajHmWFEgOVEblP5ozkWMu54uXduSeQF9kt
++FJH8Rhr7JeWnzrNG4LmXeh80JG1GPpn4maAKzsUV9nyzC7Ixx/FCi962oCHxcN
baoVg4+MKIxaZW1pEUxqh0k+ubC8oUADXT9xHb+TrYNeiBxVUcXLvZ6Szh30y6fF
+cFmXzQUS7EBpAizZYFFaN1+epwfRL/hDjDDSXsmiR8lCSe3hjcLOCemGMnbBdgb
X7xmwTartK0WjgWIYUWz1ilOqURko23s+rfoWwuZGmtUtofx+mWK9Pod/R/+s1ms
sek0MpvWbYebQElhx6+dJyC/Z04xiAfVG3+2ArP7En3VbEn/G6Cm/Ee2gNM5OheT
/YFPqTBY7g0dyfvykGm38oOoECsL7QoeEI4q1mm4E4jik0mdRYjDS67ECNUIOmnz
zJN2JlHk6tPxjNvvALuX0A932nC9TXEAVe5ViEyL/dBYaDfF2+j3eeYRhqMC7YTv
u6Q0+z65h5QiLR9pMaoQEA91DVYnDgf50dnXqZJCpIAJCNEqCoBDsm53UdRSVKUR
/mb3DV+1Th5j0CyqtjzKnlYhUCN5tA3h7oC0uhqZV2SFnL40YwuMeH8FXdyR28pP
k0/8AUIriMfdpRxVYNotfcJEYpYVxhiv00tFi0gfHZptghGvaHUg0nE/w2d2VmFh
FbfegymzjWwzJOYiE2gvcZMqUM7pZwUBCx4r1ehUehYZHhYFZ9zyuHZz6WxUB8zv
IpkUfY9up6XnarCGcb4A4EM6BPepCKGgxVowp7md/L33OqZ9EhAb04Bu7xvDERZk
MFiyxYrH/eZZq6OPcoKECD/mr2RNYzSNvWEKOWH3bzZs/JocctrL29PUmTnZX2sY
mkZ/btruLeHPM5lj59uzDEUpi6eFJcfInj4HcgK36ertHSG82M26ESTXUXGhBOgE
KiJV2d9WXrNVmzreVgJqhMsdfld7/CfpNoLdYDwAt1bA+gQ8Fn95jvha6BFYRUaU
0FTXUscZmI9loK2eXOfEzEq9l55xdQZVr4hi0bUKAMBzMDWOTb9W0SOk3XFT2Yj5
VtGLRQewF85aJIkVXOajJvDvnVbMxtLHppIsLUXgoLisa7y+CVk5706uJB1jxmBM
aGRrloaGEf2TGTaoupweb238t79CxGRM1EdGCGKy0b8Vm4C4PppexSbpdY3lLjBN
qNLFhWUyeHk1l3vSLZ/DBL+l/8Sd71np1u3W/sNX8U8AWt+/HfmyxPXKfXXRVrpS
H1DvJl1X19zKiCqduIqw98wqZ7za21F+gOOO43ADckkWM8cRFXeADRWJ2SvyIPrz
D91kjVYnR+CvE0rak7F4IUVPPlVZjb8L6ei/EEBpEWT6/NpA5twZn0+fE3yz//i9
D4QpNfjj8OmWLnXrROf5IHck6X6L1ZjNWfwGSdzc8ERXfYwhVGv7I6XgYl46O9fx
LJEipK9WSTvlHi3leUeC+svuKZmuxl4XmkJlvNc0/YCjbvHdLVgY0w7SvtEkxwt9
FoA4ir+/I/8ySoHKsww/uUMWrhdnu3TDboL6wQrmkIEs/N9vYT4I3TqY5k5654/I
IG8hMD6NV/QJ9MG3usWGG+9R6ezi5ISolIk/f62HvKxTCWPGml3w7Q8y5uDQV4Zj
7FsQHiYlou9hVG5QieDzACDMXss29k3d8Qk46aF9jKy31KMaJakixysEVps+1qCc
wCgXKUwCDuoXNb2gIEM6umSUUAqc6DhhXxPGMVIJ+FR9F+1ac7lPsuK7uYxPkiOX
MAt42sRnoTEYEyNhezQ6V7uq5SCBCn79n6rM/c5Io/44LgpKaiew8cHcVabgUxOa
HXocpjJMa+8F0Z9Fe7jUuNScMiOSmjKYFpRfWPZQducxhVUwYA5kT+jEna/mR4wj
tj+D2iocZB2sJ6T4FSNP0qUAViVszhkAtZCaZTN0iHn30iNm9X/tJGDfufpKbTHI
4X4+QodFbRo8Xnk3qGdxMiw7gMaPGs0uKSp/1guZPEzpk44uTZuW9SiJeuyuKrrJ
qOTfzizRIMU01z7U0dL6K1Llz73ZlSvZAnDU5ys3iN0h4H7039vSrDL/1moyaeEY
IY0MRf0EIMIvQimRcQMSiJ+b1OYjara+4UF4j5Kc5/mpTrUjOWYHmPv9gRJRALKS
psMNboHaocboSCj9/dfcLmpGZM1IE8ei4iH0cGA0r7n+8WbqSgVKYpXRMFRwDIRG
mD1xuGKPM2bEjGHcPBNL7pXl8WtFHMNnCt6AD5SSH9kMTXNzNql3ab4V0WdDsmql
KtX5u7CrmdrPxrPRobQ2NHIvb0OFdDwxOnbOD1J/Jg37XI095ussehVNp/vAwEHh
U0wOk2uH1Su6zZpSnClFcBwopW2qGJPejhs5eIdQfpTBAg4/Km2cifihDfzp9YAn
Q0g1P9gmx5aaGihNDBflQHBcDN2EP8CxJszj5bzUoGV0ANr04ZNbICKNOud7qGbG
SUE6hXiF7700DPNWLJ6vOeByEZXNojwJ84tXu4chXDXZv8c0Z+gZu0aamrWrBQLg
swk3g7igd1wKmUngQ+LaVlzPhEwjjnaMS4gyCM7D1nLjuXBWXOK468niVr4xLIBU
b+vrIGggcgwTC6624dx6779udMLIatWpVIBE2XzVCFP4njNwCMEHJaGSG4dGvPCQ
2PSneXUY5Kaq8VeOifS8mN3vearBCLBmoV2skzty+ab4K0IfmVgKRfFY0luSrcWu
UTkk4Xk7E1VoYop6Bt1OcMlDI6QDiVZLTz7hOmYqTS5Jj6XZMf71RGOB/1Jb1t93
r3WcO//8V5BVnDV21mhZ4hMYcFsfLfk7MS/2ORYk6TB1V/uIjY7vWDP9NLcX+Uep
XpeL1AhLXele03dLbuXYlfdjyibrs9ExTH8hfg2CzekqvJDxU3/Y62+UfD1Rk+ee
3NxJ0hS4bzs43C9atuloUPhip+BSbZF1BY2pP5J+BN0Mmhz5Hfe8jTpgSrIokl6I
J1TiwFd6u5laKVNHx+VFhNi2/BmD3w7Vr4n9Sl43/bCFzJneFPgkNE043gvt2oC4
J6sxILV4dEug8Kw3jN2ZqB6nBgVElCoZMEZZZeWMgvSp0/ZcvXWjC+yTOp3+eTH2
iQbMQv76lmQFLMftTXSz0/YJds4rZXHRW66bj0+o/G1DGfUDJyaQE7ISsAyUZrVO
yKPn7thChSu972MtLBWLJep+PW9NAPLd0BR53Hmd27jLmouKOhL29147cNar7ph8
oZCYw8DKtHMcNMmFK3R5WnlcjYPwVjcYvD+pSwk0kdN2K+vuUY4gbfA7FcXKGRL8
/cptkpTc2auq4Yb5givfo3bn5NzVHBRYw2wWQ+iASoDduVIznZAdzKkRUonZZb6D
0qqKcuD5YQSbxG9fJ3XFPE84amgkh24s7Bsikw++V2ub9hBIsn78Ea7PoHBoUqtB
cykei78bQlVhvvKbAtiLC0abgAIl75z02p/hg76vGU45QB8R/FD7J2/dGH/oYvVO
DPfAbxT0+IfqWF5xWkHV8HA+G4wFMzRgrAdfAk2qzqs7Nrjr6Qgz9XRp0zDPslRB
8zgSPpC6T1X75qcJ9hUbvgF7uEyK2Qy5wSQZxMT/XiRICr079LHqFmleoTKxl7/i
Ht7yGXm96ritoIBygj0AhfCRwD3gCXUE3aBbbLarCHtbx79jjZ8lC++Bdeuiyxdz
5sIthfPttDNCYGd8ZR9NFS2pCU4Tx5E5tYvXsOeeIarJFz6Aqdv7mXz0z1xnXa4Q
Jox7cl4hwD3Nxv9io/6daSO84VtCOmfZgmda8H80RNPAX04wSbrpJS/XU9JhwlyG
kR8gohHxvhCjIKkKXqT57PgICvlVwTkIYjdp3Cajcx9gcSnJY8V+63ZEJ2IJ9Hqq
lhwxcCqDq1b4Wj35Xw7gmliRkYgQ8dy5qFLUArUgRgU0O5EpxEy0QxYQoQc3f2Oc
GNGa9igDtlaRt+G7tCZWjEtlYk0xqKbqsL+ANKclB63uoCZfg1KHkeS80lS3Phds
pr4kJ5RB844w0RCPYMBVkbjCnht1MfZN7LYXksT//w/6LrExCnocqcooCuLQWzRb
9kaBU+L36QGsXl2mIxBDdlpafIZwDxed7Ji7A3TBvOFh7nYqIagEbKeQ1x712Eaq
kttyAHlBknPfjKP8EYkRU30pRprzKoueVN9SJMkE0P8e2f8hac2XFLgU5Y5DXuHI
3l/Pz8ExegQuFNnIlgHzRHFzZ0g2cfKt7CK3W+IxuNXeDVxZGy0BYch0XEGKvPZa
JmRrfud9+xIHb3/qSEYJ4LyQ97UO9d5cTyaQGPfHGUa5LQaXLW7K/xU8DNGkkHtL
ZZ0zJNrBADvbztDRt0Cm2aAjUDBLWtnvXLGXCN2ZGmitBT3RsAXSyyz6BaSqbS8y
LW9MDmYcg6hr/6D1ftkQLfp34COc6aYOT0sHr5BfQyxf9JGE8qd3LZwVOnmjw+6L
MNLeNhsEDXQF+ephCEQXyeRr3j7isxqMNiHQVQSnyDW6r89unLDnhcwWAK0X91it
Eni+0ULKREMdF3IoS7f7pJbQFNU1ln+r3Xjr3JyrGTGCBkaNxvTeN66rHck77PHe
APaXzMuAuYjqJbLKyuDbTpLOrEZiBU40Ipsj0TqTSdjFRqD9UjsIzQes0TsskEOk
3z1uMc7ERBgzcBwfLxAAkvJReNu1rbACf0CRudbEPaSQ/6VbCGtMOUFcCf5fdB1u
9kRzjrH7tC2s2i5KCWYlVhxJjBVXIWQ10BF8Vuuqp/JaxxMSGnD2Ks97uHnnGaSs
Nb53XBQ9ScfpQd0Y4OlLMBnL3XJL1dCbzA4PsZIBb962Rd/H47U0LxlEndoLwQpV
lm2Aw0KMtNJ6z8bKysRR7VmogxHRv1c/PwCeBAS1yc+ZeBp7pvh0DAdgS6L3Iywk
52HVOCi62lDz1LKBsI50wfxIKAyYMzFDeZwQJlxZJEEdxjT5UCNr398B+mMC1m8L
9rJCkazmZZZWQQ7lExXZoILUTvarrnhRgOXSFRSU66L9kGWGCEVNWHZ1QCwOAkFS
vzqoT/WHo0AEOh7Eqjhr9R7GSbMkUJ8SVrMptgiL5MU3Y0TrIPetbovjwU8gwjS8
vEyZXUEYqqmavDeWgWVvb369JcedXC/rua4xBeBPRIBizSt6fDA4zPZom9ApsfHn
/Ro0vL8yHq9sO6HVUpuADt+Lz6dkuYCVOSFMgmhMrBr9/157p283gxUtLGg7SW+s
ztkdfQ2qTC2pIj30RGgRWiQDQRbaUQm9a83Qvjg/GesTbG/T5H9CdOdq9Y1cL7ok
YHSfPQeDKO1SpjrAZTXGnHf612xwwy7yMnaRScxZDRjmNbp06dZxFPlyzOP+7Rdz
EX1R/96bvRL/3w31MvjAS9i9y4hhll+45G2RaJ25FHvHx86Tvn9BrLakGzTmVbRi
nJPS5I/dhKEu65fiJLz2TJVfMkGZn97AftftPgeeSll5txlA1WSHS35I781rhomF
LqpuFvfp64/q3ZPod9ISGFcuGfN5MxRaK6z1e37YbzzWmI0pQsOPirGuBwo0Qmcx
lHgtFR1N0XyaHh+IJqsmlYeANHhWb7/vsw/TTjDuUFE5Eg53vOSiCDoSWrzR/S0w
Nlgr3NH4g+/WjlxPhlNKV+GmAnFjSFw40YUdjbfajkXF40tvig+omgKX2QxNOgiE
+QfAXQ/b1iwKSkkHsjBQSq5ZKwmcLkQ3gutIIHIH+WHX+W+cG5DFrt7iyAPKh00y
ahVZZM17Wrp55S3eOVwO6vafA9AoR3pHgmv9mMi6eZeK2xoLM7uJnhRGRLoeYQ6M
ushtyr++auytNVyr7SUWyk8GmOO3FgjdmMvqVE2lU5bdv+JAHT2EUSt0Hs7g6N8Z
pZWtFTbzEfpmuU4VhYpyymklbDxCBrqatv8dWQ7ZVQneplOxiOXUZS1CpnCkemNC
0F7xUuNZjyXz0qOYBF9/kU+qC/gzzE2N4FT98kVV0xP53P/y3UySRiL5oCKXjNaV
f1afilDjp0Roy3A7MkWe758vAZWgGklO92b3gF5Bn/Zoj/G4ivwOqbC3Jb5iNdd0
sGuTWEWgEZ7GwodiA0eE1FjJ4BZOc2ZWDsWgDmntZLXAaM8AEiiESrOQVqyhVtSH
MhlIuhIsP23Bi9fLeAmLt2ULTjoPebb+b1ViRUmwBMJqiYeMZj/fP80KoE2DgTSt
gGA56eybZnPiDbjNqSyCsU1q/rkAxBR+YFVrFLrHKkjwux0hYT1h7ZsllU7yvG9/
rM1OlSRZaUZcE5orbI8bJ3oy5n26KdejN2ih5boXmnSq40GTPQI5CerW+IpESZGc
TXCGIOWPn2xyXJVN6QIsGyMKB8nuO38EXxY5F7IqLpbRAJGSJbDj4MFYaIjr5rxe
nF4aT5obxuEE4G/2yyxm2OOFU8qK8lyFybidrIZ5pIZRFoQ3qntghDr5mSIOnN28
qtrbBdgGNyfIp2AQc6gkcqnpZapMYFBlsQASEF+/Sg5hl/BaKocmKl8ERgTJFavA
HAehhw1iQTm3f+b9LS7Wcn6TR6Vv6KFgdFCl51QGBZecVLWJu/DBn9n+f3z8JFiz
LZbUOe1DVl225Mnh/PiR7QEnWxz/mUwiVaUnaYbOC+x0yJMKX1XHYiZ9lmzREYSV
2LCmHBsFwlCHQvoNbfiPNct/TSJLNT0uSyz3fvrUDkRzzJB+Ijxr08NpXXsM/zD/
lqYnkVZ98ebKXj3RLKHLEwyBBYix4btgJYNbippDP+mqnFe29uQnTvdkfijRfXhc
3s5Gnj0I60qmDTRkfYrpKvfBw+hMgiDbqCFiuJILFH7UvoWU0wthL2UtCG3jk/wN
v5/9oxuq+Dinryk+GpcXK14bMFp5iF91y/IcOJg7BB1AHvYx/1qmMC7+l4Wn7fFz
hlar2FAQSMK2AMcQwCj1wTdMf3divtR8xSNOdgl6vgMrJLRo5s/LSJypiFxKF9Vq
jtWRKXDuLeC4LtjcFgs2daK5cLAZF3My5WiwkW0GhkkiIfuLJ0PhSLOwVUtWNFVz
IWJ5iY4bbyh8X4ZxHal7pAm6zpgNNDN7b0vQ7/Mu0FuEwI08W+9nnKIg2Z/KkHAz
RmUxHdoHDbPTtOBTjmafmA0CePakll5aJi/c3H4DlxcgUZM0lg8P1g7iEoYU8M4b
I1QQZlOw6l+V8+OhItvaharW1syTztL9967iyEuoKO5AFxjoINNI7N1MOZ49K2t4
u8S3xtuC0xVrOFPUZIown2oDyJl1B6SZ3cZ5eRMGrzSsABP/TGyNhhc9yw0v6BO9
BI0Xs8LH3m3/vCvv7BueX5YFL3hYvorUmnjNfJVsSPZQ5TYFEqwNSr6EikPU29/n
UCsyUbtEK5dzQ8S/NzmpTpJmfponSR3qQLlHbXeBWOmXwP2LbHzytNnWZ15hWsVs
yeR4l8z0+GZ3ZnhDOfwmdc9VX27zLphxxr5EysJJs3n7Gx2oxMrFpF2bjy1aTOJV
RTVmrLsYmqZI35bzqnItaZ9Q4rD8g2UqS8v7B0AwXuEaiEcv8UfYF7ycosWt2JzC
HU3BayAZybAbVYIzNFY6rpNmvaYMAh12jlPOtrC4eGZphobplvDfiFyXR45W1Kx2
ltCMjgzGuDBKlRpc5JiOt3+Q56g+AC2kXzRgj1Ga+2wwn3tFGJ/krPk1ZXHL3wcc
jnUKc3m+lE75sG63TEKJpfc8doLY/YmRWygF58HB9jhT8geR7yRAr55LiAIGbE0J
BwoFGeF9kh8+ngypKxBHqr0gL2d3D73SQH2LjWwFHZ2T7/3+xxMEz7QQs76bSNcq
8XgI9/HRLJoQbWePNypiO692neTpyVz41YlhIDKaP9Tlabn74PWjE9TzVLuyJe53
cmambssVqPgQ2cLsyC1794VC27h7nPFs1s5Je4ayrQmUwdJ+Zupsg0rsdLVSnFsP
Ho4U9MDwawwmDzlM9UCcacWuaZYsft3HZaQzeeGbfvhDrpHMBCOVwVsiXX4ug/Tm
6HK3i40fWci76BON3ns8PaFBEithChXhh2TuXEcMvCXxrYvVPyQ4FYOJ9ciskwuM
OUfMIbmuMog+QVI0ZQrp4Nb3VaeyWyDUd9Nd3a7TnVL6IXuvctiEI1XG0FTGgcVE
lZY7Q8wR79smJ2K5BKsYtC/PRH/5QbqRcjHIqxzMwk0PeS5zTILrBHfvxme09WXG
YdPj0BNwnVqW1yY3VLDA+zKYRJzT4Nf0JyKm3H1/0bPt+Jn5W7LLmDpfCyzuA5IQ
1AoqJWrnyXbd9aCzut070wO3K+fUfQF1p6xcqV99O9q6Z6PvKnBoxeBDgllyIjFO
gCQ4duftFv3JBPs3gd2gj0fgTfgUSjDZg7e0AKvt8H67D/zraJptx9u04sJ2exDb
n8Sij5JeEI7kYdp93skcaawEjlwL8S+j/u4QhAgU4YdXggjAG0grewNliKZg/+Se
RLqXCsM2A7oZBHNQnbc07chemagl/vjYjA6uWXDdkCS+Zk9KbnyKWwP6PCdrxWhR
+xzWE15PgJoLD3+PMrJluOFfo4NO+iRCZnT8TCo6YqlkHMqHXDDGnmLaV4BDEUXO
lK1hIas+3fzIwYkKEJDaL+YVFocGYYmE0JRRNAjGDW5HABjBf4Yciik8151aR7yH
sKp2ZNzdVt92rvRvuGK/SaqOHCtf2IAkdsw1kNleTARRvotA8652bhaFUKEUc0n7
EGS06cqNX8oFZ0eWWY0CCcLtE5V5zXP2HR0EBgwV6ajTZa0GcEEja6OAIjwaRv34
L2mJQHWmJBn2sSdVXhpwoOUOYUH/bm1bBID+DxtgIJzh7a8Ds/r2ZW66WHgiunp1
zIHfxPvQKzl+7U/OiBq45TmyUgPI485qzVv4JrsGXC4coOJlTslta0KhE3tPTM51
354IiB/tfTOxZ1Mk/qiZ5MLj5MGBcdcMct8B8Ffs52eqAx0URlFaaOAbLLAFHpSD
23/v2jeVv+dJCHpvXwPKtdGvkaAiwKvWhnu1gqBfH+R71Sa4yajjYO/KTUzllj+a
+1Zbrt48AEsD8qwY0AB3pcXBOJEm7QWijkose8bASWI+0iDUZiUYUa6RGm+CHteI
sF1JV6nujnQ0AGvmONRJrMKsgaLyUCMgWgCpzqpjpXVsZ3fe+sXK9UE1wCaJWjGI
Y9uSwX8MamwMcnrUwQdIbls7QCvWQMUEKyyNo96zfydejLH0ozUbf9EbVm8YNZ0G
rPmuNkldjuPI7yeEUE+UYL0A/AlvjJLhv5LYbMy6kCBMT2NGpU47bDncVNdaN9nB
xt4qCP7EBDdFW2oWZ7RrYdC6qqApdhhtC6p4MaeoyYagbobYxbFlSpTyY0+YTGX7
eitQkTA/UUa3Cj9FzLq7kr1Gne1m1GNEAy0G0YJs3pfDLWHBks0bbU2zC9IkjR65
8/x1SXG2l80ytoGxUbx93+EzZ7qddEwTNcaoXew3vlLvxiKHi9O+xIpGMOmRPAOX
0k68mbscymzl/dTeFK/zKqb765RhDH+PEjLYI2PLqMqLPDQpbf8P37X9ne+b2M1K
0Ww2FbhaUXHs7hHnlY+xllsrn1ry1QZeEPm0NJdm/te0vaSzGyNpG36JEXbPZunz
6pnogqrX901jVNXdVQ6GYK5vZYh4xGQAqESuU8gTV4fmjoN9ePARB3nup36Aqwzc
7SkawTMAkZI4A9ZFnYp+lDg4QKx0fUbLUuhn2IX3uxaihF9dyeFyKl1P1T1B6q78
aoxDDsyvShWx+DTg1LEMtsWg8dWP3DT14jva1s8UmaVonBH8fV0mzb2QppapxMfI
NnYyxzA052tZ0r6Bk4UvOM2E1AuDjgnNzO0dM7YMt5uVrsIEYQnkbFO7iTs1Ec9t
uoz2aJWNIEBS+3/bOrXRz5LGujn4rbdsoFYQEiWbgotKFnY7u/7xP4ydUZQJJ7uq
1SRlipQkA61kAkQeHqZKU10v5trENLyMhPM9mWN5T2hUy7oxBr8TlXEZljwsA8Jw
FoFJ0gfWmiDsHSoRxtIkGqgmpIe7CxKXxB7+CTOg5YyUx/nD90hHn4qwSmWWdiTM
//8ymnxNFLJlk2OeDqpQ1ld+hAQpGu2QqQzCQSliz6lbAkTy3nqDGbCYRfF+iWX+
rD3viRUA1xVYAY+teDu37PR29sAFRiqIT2LDmj1ycuqMuAVRkyMVGOg5WD8k6qqJ
t/dJ2ipiswzYF4jQM+kldccAl5Al3P24NddYZFF/pi+aWZPOEGEFcJgVNbj9NJ5W
88hENqKct8nmnffkpay3b+q1SddubhVU3nATTptR1btNgw0rdykf9y7+YftMLRVw
m03vER4eOvKB9rsE3Mj790wg3MRXpfYgwBOffuy3SHNT1hHMJGthJ8GaMwuzeyIU
fILFo2eEP2CYeZj5RcqYSuGTEKVsnMP1Pr3Dar/uQUj5DSuQipdQdZAXbRJtvuQW
ZP7KaFjXJ30jZGxkDyqUEN8ZGZgM73FunTpASOTwDYUd+B7pje7MBJo7wQUfctZH
N4i9g0F4+FwuINSTD7hl64qzcm5BzAgCUL52uU8x6WqLwGSUo905gcQRZ4XDfEoN
YpoIaJwuE5Q12e+SKnj+CfNt7ADjIutNbw8A2EOrCmgrKPaQdTjRzpCfMaSha1Vc
0TaKDlu+VSHLT8WVlzWtwojNEuYFutPsGK2BVdwCjYEgztehPVQpwnoOd1AYjndk
6SXUBUjhTPxsoqQOkXVPxPoYNIP8Jj+VsL3Qb6/kjgmt5/hqcWJmKdNC+3N2mOlx
4D7QkyUaItqi6NkPVrLyGNMDJNx6Ljq4G/wz8Ba/wtkDZet1xwN8205z68tTh7jp
9wLhPQXfZyKSM8YtENCdHIZJ6EYcx06QxQvOB4+wkeraCbUlUTwSGIt8D9R1cxpj
jUsw+PVS0ADzNlzkGclrZPhzxSbdcav4n1ekp7gPusYFbQ7iEyv2ZPM9vQT+wTzP
nCWLofv+r6we5G18isK3FppJok28413SpkEn9kYq+ZDRfRhDS0z4xjYpHhtI3Rpt
TrvtdXQN4ZxP686u0UTopVytM70ZFtcuDUXSffFVC+ah7hSZWGSUfDR4qTXXtigm
Dll/XhMUfR29z5DBVQSZuiMgSLObtw3Rh4ZGixeK/14YkEdUazjhsOYBcTzxxJIp
rRiZyK3xdZzrNn5/FolpJJz2K76MnSG1j2f1WbauV1doYQIl6wWFTgM7iqHHgt+V
Vp39g+dMY3EayGavJEkMv+1PWl9DcqET1pefpVGeJxoEL4R5tHL8NQ/ZT7ZYPnlm
tUVLad7Om81xpmAmryoq+XG5vyZ1rqlfSdrcdVHiffdnkWd0yOEXhGMV+mENBQOL
K+aVXxIEtTwXfr+GCp7n8C0NJUUvSFcc/mg1NyIGA2xYJvJmgoFzNyJSd33N0Hh1
3hGlIGDj/t8aqD1QmGF/DvlD/Yk5t3B52FxuIcHXaDC7ucasH51Tfc6WWnuDTTGi
+KmXzAirY/yqBCbUfUUp6eWmVMHjP3GPMtJu17T7vIYyZUG9tZ1phMnaVnzvd1Gu
h8wpP9CZ1wQ08FZ2SicODZGOqJZHZVtI53B8yH3j8rPuLW6wz/259aS5GFz0tGic
q/Mcv4UVNN1+H9xi8J2FzhYnJHNnIhneZkB117o+bo0DxI1O2/i6pBjZLiz/nvAb
ba4kfDsozcm0Sh5aFM8Q7dnIOw6oNiUKqa/PoO3Ph6uOzlWtcjGf3U08nMKwp8NI
eX9wVRR0d2BNaoTw8Sbh0iljJEgFXD6uzwAbZk505rKK7DCOBRBWVSTr+Iz6UpyL
LraVvsjzp4V61RbnNfX7QBRIts0CdEOlgjqZcGLGO/enUk+MECf6qRMLSR2y5OFY
hHSmjGt7D7Im26HSieUD3LyQHOBftKVzzKoaKxQ3fC1kn0xMQnGffGl8VAJb5QpL
+aQeyp+UtBnthbY3Ej6sBHqGLyMt33z1LOesJtF9cqtz9Rl6F43V9NQMl6KuNc6t
4pF7JZOlbfvc7J/QP3BCOD12ArkFdzgipYAAiFDVSfsuVw2PYHdPQr9qK1WdcJh1
nK2fqZdjSFJ/MhOkbcDYm3FOOyFwBMVu7B3oB1yQoHx2N0eY8q4qTGnepXxy9M0R
rhQ0/bcw8SUuS0Lpdvu/vRzs1FI+eQtcp1TmmlElCl9h5DxorZ6r/LArk0OmeIFg
ifc75DDi4DFslTzwDm5UUSM9KVCtVRRFDdsAE9CndbbRH193/lPBEktIgq+JjrMi
PnE9BCwVImq/CYu2lkjS0KiXSD/DK1RKKyKuGUDb0+H0X7cWlSmDbuY3zwYe9N3X
f6f0qkWFZ775ybDmdiFWhZvaUdITReZ93gZj1yymT8ynYAERRM9yGwwxadHskDew
D5xuxHmppjwhqs5f7ofAYUyG7qnrISMDCy/ixiTCQHokLCPDILwR2+7n2r84B+Aq
SaCOkWkRbj/6Xul+hold5bYIK64EZiIVI9Vn/tQICDeYPwg/gkMCj9VUwm00ViBO
M2R0vJGMWU3sx56XX436QmNM/aLwqvs+ruRGFKAhlc4H+9u+laXWYZZZeDsGONiC
vGAGxuZXeGCVtF/rs5unEl2Prm6LED4fPTMaBGQhsqeX/s6lp0nQovIiLapBAkTU
/2ipCyZHPlp6i8+5+9nRUapqczXV78GQYAtZrwoZwx0LvhIWq7kofHMSnxOGfYQd
MN/Z5rsnfHB++jPjs5XSalyQN3ytlALLGh1CP4Bhk5tWwR9N5ZDKyVC/lYpW23L5
QLeOq8TRWTzVy2/QEHhyLpLOQugwcDVn5JrBadYVNrFpSQnY/ixeP2qJ3GV6uI9i
gSlWjeZt5+vl49TSo/hcictv47tU5VoMF2swv10u998egfNUaOrea5i1QzFOvZ/f
F3JaLigR/NOqtFzMwELzo67nWx47TgRjM4x+uTBY5uwz/JnyyHPR/2jgzbu63xO4
Svz94cwn5XeKY2Y27gLuNkVXRI2az2cEVjSMEABDgmOvZXB47Ly6kQdzaRFFCbx7
lyAjCeXapAAq2ra1H/+jiS5Yyz5seMVuCrqH4qw1eIn4iwDcQVhBsOWUk+uZpPY0
Ff0+v1AQHf8ctKOABLqw9kP5VjlkXsIwfmL4NNqdiZ2TnVmPUO8dJXa3+mqZ2a2L
s/UqVTwjmVveKeCM0i6BgkGju4Gx+PsEZrLM4KMAtdGEhRf3ndM/6lDqvXqmFz23
VEXEQdqfyWEkqss3f/qcQMfM2Diiq05hZOdd146gtp/7ni10YYQ9KcE1P7EVedFQ
/gPTpFtOLlTx/s5e0t0bcBk6xll+Q7DxSle3jFypLh6faFAR2E3dOxnOiD5Avn04
5YnURYRQjoz09dddatSPLKKqdfCII4g1Mn5ixCuNrfg8LeK0m1mDNibygQkJZrAt
rfb00eD2CftNV/uOcWgqW6I35UAof5L/6DR1srIBWXtwmRg9Qi05WrClnRbq3LRf
BgLSthJEXG0gUbF9sV3CEc128X4WuvELzM4hmNRAL6bzSwc0Dajq8EA4gva8qpAJ
5lGFljpWt8Hplh4888Il/5ehscsHkUgVjCOWJcobbjnbkhOh4nQE+qcxyrnYZWJc
yfoDZPjWIP48kgebWgBapbqFStgrMu6BY1HAO9VmxrmwMEwWfGCDlWalMrhXaPzL
EsqxmPS9ynVGeeC1T1eHa7ytcrwFxzG1R0uQVuqXe5eD6dexIgh9Q6ABmbxa5z/N
bAizQvW73CNNZJHjOvM9ULHKQVdFLnlnz2fcTh2h+BSWKCOAo6lvZu6W8hGxaI4e
/buemZbyg4C4sBrA9t0PUELmRfTgsvap2N1l5zEFkjuF/DtclWt+NjgF7YarPV68
rVowfXOum5Cu5ZQ564Cv8cd2+zaxyq2uHc+4EMwx1sQ9f/65nX7v+h3b70chuby7
k4o5IQEoVXZ6I3756bYgej5ZxEEmbbzyHobaAg4IWl6727mrI+eanBBKQ5bA3liI
8hadLLMX7BgOvAOXdTC0Ew8PJRbMXx40+0yC6LXUUmb5T7VPy5CqPYQ8wZ4FdMQy
H5DwsVan+D5RO1P2o05A5TkitRhhK5Y3NgRWW5dosi5lFKdWc34QGSze2adBvAN/
u/yuTh+MfWHFns2gI42h3xSRKShPPFu98W+usALH/5gIMUOUqh+sMub0Y6DWDJBP
+djBJVuM6yYgHF+rufdztted99MdSVarGBnFrzFG8+4NM3plt/S8An84RpmruB0P
R9EsJeyH6yRppHDhRekMKz4gWUPyKTq9qMMGBpNJwFGpCfkPl/0yEYdQzKme93a8
GoaYg6NuHxF2ub1tleCmXu+sA1jIeMm4Hc9x35BkiTkJNIJ7TsFcd5+qamcfhayd
C04GrBHx/Xx/TUJ2BHdS98iZnd6D3G5gDOhbQrCur6qgmKnQcytJZ11AGpZUKvFg
MFBeE3RoAXy6LbxT+QaCXd4Hf3WMywZI0AI8jpDLuygLjE1DkwWx1CkSswmSGXgC
5IDTryZlrzsrHQVSJWcrhs2QnkbDrNTXFT+mcwYfGD8Zt51oU7UYGRSMkEAtF7kD
fncq6oZaL8gCFmN1j+AY2NbY2hxn/XSYHe6C5iv0Rs0IZz9PXBHGeZOPTn9F6mpB
gPH2PGblyM7gjf4yvCoRahrjIaNkNmSUiAR97WARQ3wx1MX76S5I0mum5rRGkX7b
rTQqRTdQWoB7huhoaw3riKG5+7lzGGmbgcqOLWAPamXN4rkfdgjMOHKqukNcpq9s
CS4OWtk0hFUnZbUFxrvHMzTDsqy9G9gzKoDHfdqjCqgCcoV1eL7Qs/bP9OzcORMb
Zcc/wdGuXXMTSoG2nUEqeJreegMC9lRXCcjdBu9SwIqVvlqHZR1cuyzC0XQzSV+d
BLjbebIe2ZvsfkU4G4N+KtMMrGJ2mWUye2+HpAGU4T831y+cRcEW86tdbgnCXKK5
VjYdWza17Bl3C1XqXdw+CWQqKPzzop7XA5C7q6q7UOiyTmbiKTdglh5X6tOD2CSq
DipyTzPBMUc/AG74TRT6AoBRSuYJo4iQPmcAVAzCVWUTs+n87l0P8DrG8hkiATYL
4VDLVPIKAW/690Z29AdFercYpKrbL/IbOaf8Oh53Yc0I2HwzDpEF7LXIZjb2je9T
MUNKpu6WXg/vuN8zPqUzEPb/ArhNuut2FGEUfEG9cMVb9d8mJhzYPKH7rXrwKAMy
v8pd5TwR7QkJER+yvMIshvazZ9g4JwxM044euNWGQZ253OR0Fs6cuF8E4xUpQjtF
JFo7E91ZWxeoJuNnt+LD4HTJsu2GSvBvKKIVpc4o5AXOt2m5+o50BIQsrOODGaTq
3e8QSzNo3vrNe2jEeKnF8WlVi6slH8pBIfN4zIW/7ZwU6jkNPCw28x5bVjuan062
HTiP58VIstNmtfza4oENoMbLlu0QOUuYGHrlBJSO50ThTfyFgURGR2PwQowp2P9F
07Im3I/7enVhl4FE7QCcbGupj+LtzzAujlxxUlC+z4igIX9IImY2VvwGGVtGXb4F
9WYR8Z7xJBopvjjp5LpRV+zQkDJWcVDsfCHstUM4XMYtw7AP0o7bir+hYWuYxHgc
qIUoNE4glai11W1GF4pQdIcljXroen+vJtqfQ7WQp/NWvD9Z/89c2NN7WjeGHrDt
ZfXEv5bNq7CXcgfHODkpecOTLjtNqd91NizuXROzBIxrg+Hks9uhkCA3hEUIsTmn
LZkKd4AxjxfN1rK66Qi9SjhtjK2qhIvW9ZohOiRFrjqndaWidKzwT0z5k6yHIOlh
nQqEn0YA9TJ9BkhUrnYa3sP6VWOaGKr9mzkgIVip5BXtrc1EBWgePKbL4QlbN5qr
Sw0AotyIdOqStZKnTqCWU3A27kr0SW0DubLAzuvXzoAYzRo5DsDnQv+KYbnSgTLT
Uj/GfbPCk67TUy8fQteoo4xwFY6IJwPKU4AYSlBEJdhlD6W9tn0u2r5FFXQLSRp2
xFdL+9h2DKBIuKwQBUiCECNxVu3IrYAIRTZrszglB+9SVBzgjp4WXKfUkH/6rd8w
TQ2v3JwDQo50w2fvk+6ksp44otRnaAZju+ySkpjQYHCtRxZve2/rEs9+SQLOVC/l
O6k0yj97hIW5F7sELQqxzdxM7/TFVHuRIaYvO24q2ICB0mSvkYiyyYE9HcezrkbG
Aj+P/ONeEGawdgpD+PrnoWRse45PMmJK+SWcufcP8AjC+9uIxuDRTvrhz6arCeDS
ZMx5obqSpgJ6l7dzAXD1v0fNbvF/m0wl7+8XNRwyZl3BND9eFyUc4de2m0esZk0I
lorwhiYCVYTlqVl4WK8dCLdyRcJCp28bBPrylDl410hHXPfaj90DdxvV+Z1NBBzO
c1E5JS9KSKwM6GJz+oWVD6Xb/SOXGuGHDDRVCT8O0j8kCmn662mxXXax9nU6+4AA
bx7aUH+XFh1kxaUpT3DOR8jjyQ3bx7FQQyr6heYSNsEOELmnvoujVimtKz/wjk6t
6ynT187552tBjTHlFHI6wlSat2OHTOpUEQRCzfxzLBmfLL2DII5vcrp37SSHLSe0
kNnPsN2jH876XQz00vH8V62/ztPx9IBjsgiEmwoODJvccNM+agxFjru1X1/8YwNy
vMQYa6Qvd49lnAF7GMrFU0D+z/7nY9FDi7EvoxQrMJw5qeNhWUJoBs/kmGJmdOA8
2pArsLj1e7xb339e36UB2FaYBNgZfPPvCj15VqkkgETZQk4l7OrQ39bqF8VhXf3w
pSCFvabaOHAOOXFezr5kZM6Xrh8h53AuqhWLcaDJWvbhGLdS2POjTWrGmlSAdToG
CW5AW5Glv32/I/iThbrRewI1c0zIlxbKgsRXZzQOoL/+tSumnL4z6Oz79r8o2Y/T
+xGRDyb2Iu4k+TwNDbraBE64hK+UlvUZbP5ody3Dmdf+C0AjXpaelGWyAyT3Dd0N
zTti2NsDsaWZceP4OT7+ut8ALzSllBpdLnJCkP+QI3GiqhrgHACXkwRyyBcUz5d8
uvDLXd9fkm+148iJ+GKaYQcAgwy3FH/GEFLwxHfOOmoZ41eJazS1xqX7MZibp9UL
Brdhf094crJDeLSaaqFlvMAvEUFFPqK/jvg27Ig7YmUBDqRDT78+5T1rdKmrX7Ov
vBFnJcl5pIfpRcTtRvdFRBaIUVZ+kzcqPgI4E892XwTp1X8Jkvf4JX4AXM2LJmc/
Eb9rD7lPQB/3bY7CgKYi4DtgFaeYeH5//vCg8iiIhEdJDmlMg7Dr8cofCTVNOH38
jakxhwhWVEEE9OPQ6wWdiQmZ7qRfeH3lmKGX1TEonUAsZ4flb2ygenOup2Dzx6Q9
yjIu/+KgSkivwgSLgO3PErlf5B7sx4Gx9ddxbJtZ0g1NVBGUGKRW1fZwn82QHqgR
posFCdo2D/MPu79n5etXKZCkbjmQFkYfd4ZqZbQzUETZCdJ8uHFkZA1jOlLqoWXU
rx+vbTNtVYTisrCgjK1yMtZGyT8f1FiK3Nw0U+yGH/pkrSHoDSR3rPz4RHSIfHBj
qX4tmgsjM/GLnlj9ofy0HNfstACnej4Gb6sxXtFh1STAecoG4bf5mwIDVfY5tpWW
+v+QzZnablUe1cViksy0KWK28bkyworgQ1T2unUjZ9WABRaGKd4bCU/QRKbnM6WG
brOQ5o48eWC7VRVTtvOuCuQb6OGCqPXuR+4KoLlPOLsbRvKSHzIjzBiifaULJL2D
FQCtYG9H8MtGi90KzPEWhQh+6JZZbN0XpluVGm0v5Fg5Ix81sTteGa0ooqVoQ0n+
JhUGzddCoXVp3J35O4caUTzhFJaMAlO5JchE9Cfr3vT/n7OLZZgmypHN3AAc3zsp
V9zkVTfnmKdkgRw8X0j2SQ6v+ECe9JgywkypHjZoZHbJf/X6TLrSxZ4kmIOxdBRv
uFcWsQ/vq3LRWI4GmPSSwGg4Gd6n8QzNTyiHrVFP8M9/lfYw2H+9uVU9crGnALba
29m+0ayNJB+Ky3DtCkI7bMlYmVpmNrHqILXrp6g/E1P9Vjwhs4XXR1xdsvXl3pNq
VuBeXvuoB428LQLt29hmftlRf0HtDM0HVdz7sltEBJbbUj27KAwIv5q2YqxIKd+J
PS3kEwRD3cY59gNGLKxGft6AUunxPWNIjDpCt5EhBwiHbize5WLim7d6MYtdCLke
LKRfQzrXG8zvaYLEhdmAhtv9n25Pqb+2UURjHIbLsECUyDlRbEJc3IZEmCsumjSx
M4AJ6G5iwNyie106wnLUY6u3R5pd5prvZz6cl3au/hGOvq4KuA0lUDD+GBNiFQw0
nunVT0hcSKQgHHiLU0qcfOCfbq4hv4tP6lbEKsjfXPJJC4jgBrhc+SIDdoUvM5X5
Qz2SBjnhfqXoNMHFgXxGqFqlByJnP+JHEWAguj9wIDjHIUm3EP4jJaozV8q2ODNb
jZZuxTik4yzKBpJl7nyrGoqdoDpX6N+XZle1x3MPP3eAfV/iIAMCq50SsAkPbOGo
bGs4v13bJSxYetGrPDdMLCg59KkSou1nUasjyp9a4VYThwt5zeFbefKSIra59kC7
TU+/5SCafk8WIpA8wm9h0U50kDaS4DMr8jmpP8lO1DHUhW5XkriyO4RsusrWtphN
dBqx5quayS3ZmyHvLKP8u0ZHulYcrNml/+6MCpEKA7TETaQiP2m1OQ/tDZy3MItB
njWsCPg56vS2qcc7TblQjzACQB+h+uYhdq7L2rlTE03qPZGxa3Ij+fjzjQsYXQ0d
aAoZUSGyCCp+9VZHQWW63n25AbfQUBFEQMDzeoMmr+YOPrmFlcwrFaQ//vAktu6K
NbV4iyJU825rRSXM7jTud3pcpMyk4OELAWUzc+DgeS21gEA/pZBNEyNDlTED6IAt
ReD/5tf/MpTB9+N9GKvgsxB1zpMcFDjIXPkzhFrjpzX6dyDbalANmoJYmRTPzllB
2Gc9kAbF1gisRlgXyR+Q/kWxME8I7ZwkMGOb55KzwHyF7yU7ufWbVjd0drEamZf6
pxbNAlQxACscS42f95ASHxOaVZE3TTFgLTuse+HA03drZzRlPEDVtMl48LY69h8E
u1rq2sg9hiRLRPECIF7Le6Upt9FzavLEYqSxQngMoKht5hccRz+x0DrtZ4hQuiJU
W7NUTiHba3UOzs99ccLCtXGd2KU+uC1J3M9cNXI+rMllHQbqv820NYwCUiEP4kf7
lD96UPj3l9VJm5u6/22APatDnv+8kYdYjvfW3Gk5sRbV+7LMm5rLe1xvxEO9ZfvX
adjnlcRMxkWzuGLjryy0wY493F7y1S/bKsut8Tnwp0RwJ/3g8HhP878uegVnT72Q
MmD1uTl6vN0MBTnbZDvFnFVqrQb4glar+jKDhjZYpbbWuqXE7B4nuN4I23F3Oyb7
8gg8igcgZx1V/wkhYNaqZxFxfWdEub5SaIVWxGvCgKiZTzuq9Lr5ucJax7nCx9rS
WZaamY/hh66iNDfkiyopO/W8+WA8jWFH9yidmdjh3KJ8vbRzqxVHEPBItmzgox07
oZrjUpfkVnK7D+lCrsG8GzjFi5GWohpKfmAxIjRTmha2KqOib0Z8gpUlxBI26wch
wGjWL986Jz1LXgL+uqanReMeqjLcAmWEFtOyMNJ2EUGATEepqrL7msYLT87efHGb
tsp7TAM1m58klEvliSatCqzh7K8wl2Cfo4dmOWkQXg1Jx7J0vz4fT+mW84zbpbbn
G7RUqUT3NvUmFgMd7YA/zHzKtFE6hlHesuOqqtBrHTVPZKwcUbzcsUJyTThYKm8g
nTUMiuDSaDtkiAenYhKARa9QlnkoB1MQdWQjBi4A2BpAruGyBJv5u5Mtuas8OYSU
FPLzbLOKQAPeQ9lpBUqVUGHePkDBDOilyZnVsUz34swTeFaZze0d8vS6gwwh/yME
AqDQIgFFOLhu1bsEyMhFeG+vCb2YGMHOxoATedLCoPubjZOANuEIORzsWBzZ9lxb
Ik0vkeJS8b/MhhXS/FOjLKpQI0zZLwS7kdQzDiomHgQ08rjYsHLRXPwsSylLGqZ0
GS+HZ/cTFMgTR8iwANBhGRSDJaxfavkhZ4VnICUM1bPOqlQqnW+LU7+cyUGDSCe3
sRFRvUNthZH4yGqQsoMa9cGLrmGw694fmXgGCyaYl1pFOd/p15ItGP4jRd00k2V+
CogSuOBuGOGQOxHNgesgZ+ZHCONca6mXFM9XxWuFdppxiXCksTajfQ7tcYUJW1LZ
KT3oIyJ6Z28j2Ixew2jY6TQaGffGpCTwsNWnKga4Tj3p4vPZm/q+0g/e2GD3S8MV
APJ6bkVi+mzbYtcd04utigubWEuwCka5wgjcQ7eMTzIfxG6yih+JG8EK+mJqfUQO
OSYwjkdDVgfyaEqb2DYWIsiwGeHbKaOzHK4xr3cnPQ/Q35Qh82isckH4gsa4xM+T
KwxjR5j/e64DIOwFw2Xd+4+oDgTL7EJhcZdXXkC56vUa/KzOsAq2gfKBHVu0AZqb
LS2zk4XlyK+RcTZXlbCK+7m83yybBj1RYTi8Ocs/AllIGBCbKl0vz8noJKhTLUS/
478YGhjssYGX51Tgfz6WnRZ8XOjErdA1pWlZUqgXqMFmJKLkNOZ8DY/u3mRbPPmv
pvONQ52gNBxHMiZbsUNvR6HH+mU7+crZ25VRGNSOjioq1QsNCQAt+GqE4sJsSuLY
JQ34kUyVSYjUh/58fkqg6m2bCQWeCA2u79PbjgouoznnA1MPySH0q/jt8DsS3Ktl
NkgVMabl7zsWNZI2K58If9SoU+MROgNskTL6W1CG5D+/Oubsv4gRIRRw5HO6zDUx
9q9iiCecL7xgfu0c2loTMXhCgZ6dkXuhTkIXdchXxFvPn6d3nS1l4s1LCXfizMbJ
AFQVRAb6AlsdDHsjeo44HjNiYM3ZjUU4wHeN6A1g2oNlWfQwHVItG16GqSEmZYMe
sH8idj6X4EJjtwWnDXRh/N7c+3kRkGUbRpsBoEMki24Jf1g/be+SwgDvryqie8F/
ugUaAmeqzCHBO1qlEHDuUh/LL2Cq3PTvcIkd5E3Tn3XayXXN5pN0zdXg1kJsgMEC
ucAWaabWHDtExA8CH+fYLWRTR8GOD+J5cHlPFNOpZavj9htWUwrMskmIp/k2xiOq
7Kc4Yg7OUXmTyEc85TX66kQ4rMuFD85eYZuHR9XYiwrNekEA+GVuuicn2O0a17al
aHtDq2AMWBxA2buC8MuJFHqNeJo5OXt771TbeN9soa/vXUCu5Bnc5TeIlvaZP1Y+
SYOUskYDVEdEKtRA+AX75wdtdRPk8VeVRVecOB+NE4yosF+3o6oaypabWRMstKaE
cujjYvLaP95Ml1tfw6oWirtommDGur7kdT23E5fj925roFeUnHkW5QO572aGfyg+
IlSIgg+dHRKTqjAsegQ4bCKEj14uSzlVh5/HuKvu4kiCjFBbBby8T09yrB5YBjQd
TGTuyncwytN8vEcL4n9sFA+DCgK3ZCUkvuuPzvA4JtzC7dYc+4XKWSzL6a2qsDZ6
25MtZ6rp7J4b6Zk3zguJWzfvopfp6nh8S8fA90lRtE77C/P9ANuREbZ7S1L0J9Jj
MZZLxk2Scl4k8v1crH763Fof4LlBPyyHUcygXTYYMljlJeUyHaR0da65d9pGp7EK
HCFrTczmCi3FjE+8qMGnr6fj2vgtaZvppRyojlDJhQm3u4IrvgYiv+Qb+flu/7oj
EoIK7jPExOXYYLo0zlppf1MH05/PAYbMOpYpNwukWldcThO69N3dL0WcmJPRr+m1
qhWJLX+SF4EqK9WKO9ocomO55OqYCW1I8ru/CsRpr+jPixYxeVbnpfxuRmmDN6Pk
1drkVm5r2pTXsU1k77C+R3LgtzdmJKcAv9oJlM6P8Ev4eELl+xZp+bZjIvUArwOr
RV5gcKGEBG8xZsu2S4bRhTU0JbPmreyZHHJMWWA+SryhUpEklT+D6cw4XHXQKgwE
0jVK0X+9Cssllv4KRASO0XnfNkx9d9fQvB3gmZ9o3BT4Fx0pGEHrc4ufL9Yk/LRb
wb7t5cI7sjorK9mwfp3Dr+aQGolBC3FGgaNJOEXU4HP/qgIXKNjlF9BgGVcOD+Nw
jA8h9+cslddYf5Wvf71ABCZkaXOg2eF8yhEIoNN1Goq/jUbSTMmBBHCILD3yE5vj
DL2/K4v8apbyYwPJZNslu/i6ZHcXBeyo1UMdpVv9g/imEo10gaDWf1mPuOAsQAmm
VoEylulAQx6bZMAYAhJ2zIpV1NKlVu0S3kbVhnHL4U93K50eUZZ4Grurs1n6Y4+G
59tkMbXzfj38lZ8uIUkIsRDhja0GPaAcEvCmbuPnUdJHOj3CchbC+5hVdyQv4DCm
+vUDcUWcv2WUzD/c0WxaMr0S6koAbCfYbIRcglVWcORBKjzOlB3HT8pml8MRLyQU
mJ1Sf16hpuHonHP+beQKBJGqYs+NwpL32s/rfk1FYapZhI4UPJ7EWZD5XDhq07Tj
fDTljNNbdwvOcZqNx1vJtCFeljX6eQFFa8V13zT3zKj1jho3FH+xqzUtJ7UC0vEY
Ws3W7jX6AOxd298ozO5GPFDmDa4uiJALCu7zSEPXasY7+lrt+7Y0yXiwnw2oL/rZ
5l6HbfPTXJD4Y7PEu7PEgqubSqQoLqDyUxrcMXGjSJ/csOirq9jHtPDqCmZMZ447
PQhkuZgib00tZw45cOKCDw4VgSxh8+9fKcnjWwOEetvE3b6HGR8WVbOvUkigjYMv
XSml75+5PHpNzOVhCu7W6ZK7h8qqp6WZmHh+ElQ8VipzF1dSNVWdXl0sJSR24HRU
1a8+4Kgy3KDYibThJ9Yuh69oPwaHXQ6QBrWngS2fvGk77rM3U1iheQ9vCgLmxhWe
GalpbIxKW6rwq/UdMBRSORRA77x/8BVjq3/0vKY+l2MTw37pToNlYWha9p/ttbdM
EQs7sB5Hl4UNixiLXCyEKnQ+30xvlYkL0hVx1Avj1Hqk/nUqtQur5vbbaqepqLor
/+UzdPbWm+3lLnt8wpIrZNn8jGTtg0XgFHbrnD8iZSZWmCNKgwAThE1pq4tNQ8Pa
U1Via4Kc2te1PzPKDtO3n4H0kB+5ybXtatU8D0bTCZc6AsL3N5aHEHlvcyxK+Vnf
WL3TvkYbM2StLf4FuMvJMp4vm745xh+V/6flcNqBC7Y/6rRVGejAsl6wDQQmY3jG
d53cNbBsHMHEGtHOw6IVcqa3APEL7z3bL6h3J3MoXPKVUQhGWA6LZxweAfEcEQcj
sn90WDn+vFSKPsCihYk6OetvBW9d0/cYCV71NUyO/Ee2h8SKCosekp/byLMP2No5
P060NV2hZiEKv4Q/0cfbSu2Ot2whKxb7XuKEsfVeQCc9EntZ96qxVFTXs3m13CDj
ySHbg40j7CKWY9zUUcApskOAHWb49Ti/KlRwNesTAAWCIg219lEAQKR5twh+Kgvo
rR+PFUlyLDLTOY+kjpXZEluBhUl8O4tGzi0ktfG1zjFbT4IF7RJnYsjkmkHYuIvs
oer0GMgnyopKeQ/xagrZPZGglWO9Iy9m7oi78T2WNqMo0dce8KyVG79zjeSVyQ2G
35IhQI55xYvEwXyJ1MIt4ifUk7HAGsyMuiP/tUnxi4OhfYYxvZknYe6G/maGVbsW
1pAmYzeEBd6rukgx+5QaxnIyBG1MCd495XuIDpGC0Miru4ci8AuNl9IF2QDyji2k
LJNUvyRIT/ZskQX9B6TByiIQnG6Smq+LhuFh11KzCX2iWECiPsR0/AYSgKepRF9q
7w7rfNdMeGY4/DaPmJ1D6OlAYJOOXZmtNl5xLYzSwq495XehIgwRXXvB3KxYpyo2
m9fbdbCQZVO+sLzfLdp2G6j4bOdRbhJUQPuI6+p1BkGLtGEZa8cBjoD/Js8S8M4e
jQKPfGdGMrwHEOoSlKkwCVI4tea7oxdTlaPE8H/OjXJEm4L/k348zmtE+f+qnzxM
brPr8VMCM3ds6Ilw+6rWrPSgjfRZDRwV2MoSUnMpEjcp+Uv5TcG+EhGU3EuIX7pj
/L5Ki2RXYY2zrvULFVsmLCaGJEFWMW6cOeSkHbm781URbMyMkEfxczHJs4Viwf2w
j0YtBP/xbnwjBwnCxfsxTX8mW0IsrYg5v+iDNgooIWn96oiKhxHlc5q3YQ6qehpA
FaVQs+DwEzBOoPTlU7EhULSl2c2XhA0JMMoW8Q37nO/1Sa1kooIyJjeCEYlS6tgp
wLcWmcU+q03MyhhfcPH/AADXTPeUrDxVGhQvxZ0KGu7HLb8rSV7cJQDSFa5S0czN
88Ieqt7mqceCcl1LGx2s3STqBYNN0r2Rc6jKwRWAhmOLcytB++IT0R1eGpBrkAQD
Zt6idrJrvZTF2iJVl/T8nE7ssXApR3fnMv3i/qXELh0Wp3a1WK2y8xMmDM06spJJ
Dmn21bSFh3U2tA7O9GmB2ODevRV3WkprDiSPrObU8EF4soyZhKmiZueP1APs1CXG
/QZR4viTLRKNmwbf0ghFx/O3LNjLu7iYsWehYXwXjMGPUVmW3Z9s6U1jo8uZLxS6
M7XKrFH4gTvD+xtNGGpx0uw+cD79Xhyv3gMTGoHcymsnHzAZJYlonCBr3TRS5MjT
ZIl4TzTsu2ixSTo+t0LSGUca1Xy1zqHvT1uxHxfTEuD8MzYK64o1C8RTzJHOFhEu
CaMN03r/65vGEVyGYncUSrH8zz2Y1/wnhSLLK9FikMa3kXk0CH1ab3Mxa4zgxOE7
RZ+z+NrQbzt/4au4lPw9sEIEoLmCYb6M7AQHdMekgXIQsckQOxgXbikuAMF/esxO
s8R8IoE0Y8MwxvbsvFkjozHMWMPv/ss8vUNxDEkMw1nO+p36nytoOEgd8ihR46Zy
36IDSm7BPRg0xUjWOXA4HGoCIsTmAmyEqaBv2KWWpdeyqfHLjGfdm3XrqxkW/LiV
5+jBB30ko+smoxE8PqNwSdZgNoAMdIpnKBYXhjnT8pjHR0cXlUsmePhQq+PhWqSR
MkMwUsTkuKscESitTWZXSsuwspoKK2CH7NYCBI+fVq30jQvf5wFdYVGdeAzW0OBn
9OBbjH4sFOX2ye3SfB9Ar/Oa//qs7ceLj6AyzJlzYnAF+mVTjT6WDFuYiuBaY/ek
M2lZB5PDVojSd8n5OQ5cJ+Gbdocbi8QjgApf2ivI03N/Z3hucSifQA7ovi91Fqns
polqMOe74An+aaRb3w+aZn/lwvkDQ/8bMR6MS9O/LbzVaFKhPIlGxfRmDKvtFF1A
50mgHBs4duqv1VaFPmqH9E/EvfswkBJMTDX70SBG7KiO8TnR9W321X+bzUWoNsze
N8PvLY+h5X7nM6o4KB1Wd5eed7rbpgLVtckTjJJJl+xwajZEhcJi3n9aivwhnK5B
zc2mUttlitjf6uKRMsL4xOE7aV5iEdkFBneND0hCHnoHBMpax4HGGOlcHD+PQf3T
Blxd72sEPmV+Lfk35h2x1gbBhW3Dr/JqQleIQ+YFKLQGxH0K30MhGL4V9nmJH5On
iNOIV8Whvr/k4LO1+CZPdHSr9vC2nzVH2oXJYS1tBsP7d7x1gAhDeQO6fQrfZt/z
jRAIZ4uihLPynQcE5FMvm4us4bWODc/FIGw82sSirggAvs1CYjzQAbo7uM9EeITx
kraQfdyjmYqppqKjxQ1uufBc9SXjBlSWekETAzUHrJYmwYVj37Exc4BDsAMq/G5W
2Ooeb17nZ0JPcrmjNIXTXewiNbUGIzNc+RkFs2oMx7GahKCXFyj98zjo0L1lGKwb
YuWiHyyaV1L67cP7PRTxURPHZdG23Zvvr54hoQJ8cfDzyZ05KBm/XHDngW5Y1sKx
ofHP7WvtcKY7i+gwCU1z2FAAkNGJlv0lJld9R8veGsXiiBy/Vck0MFdYwEHM0/HB
Lw605Qc29hz1FNcFiTr/oalqFhP5V2mX0UsLyfWUb+XRaZ2CSXD3awgiP3F0/4ES
u0wUM5mL+fVR5skVaZUqVVuCCCIdFE5FAP7BElPEmsWD7Gd98aR6klKrbGx21PAI
+lOKV2MSiwRbNkV3uSTWjq/xg0iq+na45CEwcRgt13ccPx0EKxSzqzl4m+0utgGc
349PjeFOLPnHNvLuuC/ygyaizzcbO7/NT+iBLjU8Gf7E0BqRpBEVDFAWqidJLyDP
MKbri87PugoHMWsuMKG1zwQ6rge3eTY1yodgMrO6Le3B4k0pU7JEDZjF6WB/T1/Z
UachOkHOwq/agkq3VaB73TEBYRVUfQuXf4hW+luCL1H6VQilsh2GmjWUp3tc180Z
VCoY0SjbWh27Us00NR1OaVsKM4QCVWZVToXmIqp86fwAHx7AhClDfYgmpc5L5n15
m2ED4mG1P/Yj2oo1/kX6ZdF0xG1Fw5X6jP4sdf/GbCWRQQ0IT6tMU8R5pmmexRbp
w2NJQ4ehqOysC6A/9kRPx0NNCmsNZolCBJoYHVqiy3jqVNQz3yeH8ZC4I4J8LIYd
wM8RfDReF56dVmUQkKbWyg1nL0c0UfV2bZQ20JpYN0coDx1pjGGtuvoVWN3nr1zF
/ThRq9qliF2Q6O0iq+1+KJsvrkopkVyifO3HbV1HMBqWMWX/ZW/jMEaMnMN6ee7H
hJ4UOLicUl4P4NeCfFQYtDTybH6uObjxjomhrZRPoyoHm08OPkwKnWKTaLUfo56U
ezYMOd05pRV8FFnm4l7a+sDJ3v3cgksSv1cZsxnUWkk1MUvu4gCiyk3CnX7UFC0W
2R7EghEZwi5xJGdGjV977VACc46D31WG+LdNLpYz8IQ4zmebHBKbADGzFXs+eRO1
dF/2KiL4AOMgXpsDp6Ow6oTKeotlE5S4ANrRFFGUJR8EaS12MmqkNZQHjiaIS/KZ
7kVY5r8E27Mw/jhju6Bm+01EDVSZvGWKjs4HPmPZpLIrr31BqWaUu0bP+bM1IIAC
czdlgc4qlYOsiPxivzSiciuNFFLRu8xsnst1A/a9PcHVMny5hSIkxGW8P+4Kt03u
X4flMjMIemgJjZQEXa1dGEYmnhjZVATSaK2XYYXJuDcUiYaluwS2YgNrDSEHxeXd
xl8P72rsfD3pmA4qiRSJcss5UE2boNDJM+IIv6Eeqp5NB6ysaNa9gLOab8ZFyKVy
hkljFN/HdILCKS3CTQ9MVV94LH6fMEeDQKqKlWEEUudX1AWuuPNV0iYHKTSEFOf6
ALFCbnacDvoZEpY/C1CvaImb68soojI0ctQrdf2XikMqYSf4KYn3NRZvc780CpRE
b/j3vXTuBVuBzPRu5gU1ZFYQNPAuWMClIdViSc6Ica+aFznLZ/F+lpqiovVV4pTo
VM/M7wIEkSd+SYD/DJKz7hiRe3QcDK5NGEhK49mcQnzUIoJL8iUSI4SLNRSUGfrr
lXmsyRtej5d+SiL9QSQHHKlDZVF2SXJGJ4qQBmPGkdrdHJNNeJdAoFTFi2BaFg6E
k0l8qfpWi3d9P0Vu9RRLj6snJPXWet/YzJbe+/7yBWAf1TUv0WVcmsyhgY6Bd9OG
YgTUFtz8+KMjHRprn3jmd6FmNbG/jYQeRmApDkb9CH3AXAbb3237uOybLKz+AguN
RPyiDBE5eE/niec+MDbtf4Hpj5K4wbchw9bvA6k5EphxpLSYp3mGfPOIZja/lHwT
sI2CnOoUw7H5vHuCSIKeO27CYDscVcPDDpkhJiTutIKXBlJcWipR8S0UphUUFXQR
+XuKbXKLabiYp05F3dJUoJNvrkXQkXmsSvE7KMgBsSokawPv5StgxA/jaKHWP8lE
wOzpeWfqfwR5Ss11+BgRHwSllAeflIcDAOBOfUnM1vnDkfQhNRwyZcCfBT+GPND6
BtOqLI5Ji9xb8H+x+EPMJChepsp5CQGss9G8uTjkhtD7EmDaazTYBFuKqQoZG9VH
1yWB7B+9sHXy57dQTRfVpOAjf5OUDi9oa/Pn+7UzTN85+KHSKzF3ynuKFmxGUj5A
OLNot41YSf8BqjzFLd0u9nYYsMhWJEoH9sCdPtf2yvmHsJ49pO79f1Cfvhuj0Saz
Ybe4+YFDFM6G/662Yb2rHHJCizF7NxzSJii1ZGUFuU8y+1mVPQJ86IaM9SGSy1I7
XoTry7C3PZpjn4fdxGjnVawNlEo6tt1yaulB+0iBHEhyeaOWEwQAXl9yAwvgy24C
glTyZ9NKgFAobya6DZ1RLrHFSbuGWiLN6egpP70RmaCVBOiMEK95fxcKjMb369n/
0aNmKTSPAsJwCACU8nP/0zumhK1VAn6A0GD6qadqNNgiWVfyLGwDz41/nVtuPlVh
xwbd/h1gRxXUBS3+dwK9wEdAol0HIEthvz0aPx4Pzf7P6NOtNT62NlzFhelEJ+YS
OdXc/nHUn4hVVyn/CQEhYs8mpSCgfgKW8WaHSn8GvzcvU4K8wCiBpQ/ktd1k4p0z
v3Kt9Dod+2XLyoS2rpTArVXqU6ywPxZ4D5i8OIkkIpHeR+IRfRvs/P1jaL+pv+eL
IcF+FY0zTJeXAi07wfgpXnZ1BNZ/5MHSisJR6Me6IwcZ455/JiKaaUD4iERGPIP7
trwoBAXdeFh57hu4RR6QR8EpvIV2GmKRr+nKmG0OgVKlVyqSmQdN4Vtq5XAvORrT
IpFDq8TeVY1KP3cK0gmADjGBm/1uzUBaJph+QGonLbAuttjWqGiXBKbBf2WpIgTo
oykDJJ6WAGPSoZclM5YVBiUXZkf8wSUlWG+FygpDW+l6rS80JrON0abLlqRuhoqj
cdsDshcrHLixlfrp6LYZ//I4E1HKc/VF5qsqYJ7p+ax0hwP7taWsrZxxwsMrPk1d
saBSel1YrMnDVBrY9TlJAsR15W9i+K/Ok6KZsvZ4C82ZfG7/oBOiaTozcwzFSAh/
NRRCwpHuAkyVtG1s8fmk3wZhv+aCkWJrt9kS5Do0zhqlD5xKQDMzicOuifkxvzLm
GbSAgZSoD0pnI56FJ0xjXvl1KtX+U9oaNWB8NFVS7Avg3MnK+TOKINrjUA4A6fuy
wKtkDF4wkDSQFsdKxLGrn/+EAKB/NObfdtzgMASezXnXXTNqQO0DdA3uXVNxyzJg
4JdY7zBvtv/mRiXsWT5GsJC8iIO1k+9EIGFS3hTIMINWh1soB+MbBfkPYnk+eugd
nWfEs/0sgZXFs/IvRynUrOUnIkcYQN+d24oyQhU8KIRR86R0EQcRevZ5+8QjQZFX
2k7ir7R0vI4f9n+kvKM9IiBuUm+tU5SzZuQrHTQ4FEMNUKsUqXsF9Og4p2zxFRwG
Gjx8tSEOlquvJ3cr0MppS85YlbnwMscIzTQ9Pv1OoUJ9Tq2V7o/Lb3VWH8rG9c6a
inGL1acp+QfiYUyIIiN5ralDRU0H6UMnSmMKfPFcS6KrdGizWTcKVAHMCk2ZX57o
rcZfSDJW9najS926DB+BvPq1bwoyAAfV/YN0/Hzd0TMmq9bqp6AYPQA9s6Jzds4F
ORO7QVB/8uGYtpyDNXo9vuFa/5X4aAgKV1baJqksWOqQEbk0QZ6YQRjeJdNmFTNi
FajJryMo51MDIKvpSEy84xj9u97iUeAzfZEh5C8SMS5lw6hvycqxtiDZdO53Mejy
rMr359I1hIhg4teQkLi4jAz9+j7Jtggygbnks7Wzn3oAughhGxqq47o5g7hh/4X8
WNcpL7RZT/3T7+mr5Q3ESZsDpsD7dP8f0xPwFm0qnj2k+QEEtErISvHLox3pe2Jc
i+mNI9JTMnvydXGXCLe8o8R37RhPr4zj4w2erzk/rF5OY7D6Xoie4qlVNafTXiNt
mtStdM/7X/SYxLjJF8uaQuQRO/rUivDeCmhnoM8VccSGCrMjToQPDYRz5JuLWLZQ
hW8B6EqEETF4bii6dG+oQwW9AAcn3D0/5AFkJpOHxWvFZgzS7NdK6G8W4ibFxUCx
Q2kfTAmr+G2QVQ54PWSqVpUF2ZJJ9XI/epaNwHwnrjrE+3G8UrK1XQemmB7Lyf+p
8d1bawIpSLmOO7Ns5T3K9KstvQiP3ipO4XAtKVSKOykpUDW0cVq09C9TVUBvYe/O
6FK8vsvXgAYVf+M7vCXyoCbztvz7Q6XBjBMpv62lnqMiEy2mGBRRTnnnNFedHXY7
NA0xNU/zdPJHwFYWHnLHEx6fHGuf1I4pxr6UzLZZehcxN1CBo0ELApfQ4zozdQvO
Fhg3t0LRGo0T/Yb2NvylFx/gR0wuqoKXdl4CVX8LzrVht8qI2OAs1NzjgAO71faB
BsVjiQxZ/KA63T5nIGr0wB7XZp6bTJrKiKkJzbUE9wqM7CO8K9OkWLCnqCJS8/tn
zpktwGbo4XSTszpT1aLp7ydHX8RipoWuXyStIAfGUDJnE8wIrmYoXwEyffMvyHxB
bm6a+aGHeRDoDpcUpGWpoX7boltOQhS8zReBTHSnVnMRY5sdjI+VdBMbEPXE05j1
6gxGUmhneWNb09l0tR+pG1V4NmiWPHXKSsc4l9PenFRm2ppi09ZwlX2mOZtuTTie
sAzQSGYDCOjBwZJkmPanji8V788pZMWKbRFE2WsSrkO1SuPGzlFU6YuNFkq2lVhm
Zeac/0ZoZLBVrjL63K73QOgCKOzmQgGDJ5b4ynpPFxwPib5kbpICuE4Dg0BrcYah
V4wqy7xt2FlGL0kD35rDhv3TnYutV+z42PO10Q3zXUbfGFc8z2jp4f8A0Lweg6oe
0cphQ/bOP6PgWwzTwXoCn/Qj4mN2zF+4EwLqKLffBWt8E3jpGxtuP6Of6Cc8Ol9M
F1pngOlMvYf4lYQP7euob6vAkkYH+M2+ewjE87HFk70RPU6WWuv6ubjwYIVEludL
skpVt9kQ+BCcTT9V1AMOZ8FPSqouj9LL7ll3PO1kBE+kipb7uAbiMsjCHAkXV/Qm
6kUVfBGSqiIBdqYUTgpOFMUq0D9sohhuTq0kv44loFkBLZ9gzZ4aZe2Za/+ETWy0
YNIoe8pDdqgfsxNduzukW/3gxeAjDwgnsuXl/StZ7rLKBmVyZnhYgYoaj80Zp4/i
5rHP/cgFy8GRKolN2UDbnUNzw1klNIiYCHutxVA7Ny48tKRdDRw2nP3tNVOf3F5l
g2RwCLyy7Z7IF4DlYdtG2AtEQ3qK95ZdG8PZubON0xCQ7XpSHTxmYL7OoD+Y6pFV
kMYIrTWqtKLFGjwC4SJgA8V/peVYfMnbNmHQAGjJq+LrxGBGAcgOwy2itDlhoe7R
KDS13P78smccZtp1ugnCKiQRAbsE2PtRF2LNR7WPcucfEguJWx/ijNpEOVGUQfn6
Nf5C5fBe3QAVt51psEuuCFAcvjtShZ/484pXqAPkd9hhbSQVyKgds3Br++GOXIEE
2ubs+yAVRZ4/s/qh/zncU6NMLmzZFgWkll/jGRGehrRkcWux3YjWlMYhJE18SZKJ
56mQrCiF0UbHV7+11vsuaOS2SE2ssFx+5BZXAxpD5X5/uiZRu8wobSUWHiYwvHrB
wPjprWHdAe+xZP6rsz3bdunOFNU7twg8mqvzLFnqrSzP+BNbTrh9qsQFlrDyrPI5
LNoVYjGRfLt4hWe0fqFsDorE/q7MXL49b9xOvciWbxSv4xCX2Fe2ezpmyRPbzFZc
5ustLfB0x5ZYD6jHG7jWLxIc/8HWdl/ACN2SZoOWTuYNzqaHBoW6eDtQfxC4faMg
Y6NSCJtf+gLCqhlZbKXjkHA3lSMqjNYvf4Vra6yGBKufBhsjFZ/pBgvC9ah1/qo6
IiyJ8jAgq2wBZXny5h3GzOVJaD5KZDdVwsdiOk6ZlLNBBRDFEWR07O9jmkJg5Jxp
9t/0lF1SeF/VO8Do7g0IrwZX5QWcy+g6kQJnAhqytOcQVj3TypUYUCxAKG50jJ4E
VRa/20Krz/jnsVWqO1mRLn7/kB1jcck/3/X7P4CdL9IdIiFw0oJWQ1VzDUyvwvXO
jLa3drRCrzCBaqibxSNnC7GCFhd+0YPZrxsfF4dyqdyGbptQ/UHQL5ZL55ia0djq
GlfSLxsDcksBgreNsp7/wNY2DJi9kPUApA0JUgakpvw4Dpij9laGo28pAPdk87AO
4cxKbCYFDJSOBjIDtFH8ziQtNh1LJ5zQ7cIh5BecDUUcx3orWlT8pW2UdCF7RHme
WN3q7EsMMDxAeEYIHO+LOjsZm32TT2Qp3MHPzfRHx4483ksU1CCu47B851TdLxCz
mufTPRIbrOWj0PnH+RcTDCSXwfNiH0SgBThqY62kUUkZqSLtju4CpMMeIluLceQL
JW7SDfvHn0GXSM/dSDhTm1M4RLV0y7vWD+d/yVbv1hDN7P5REYqtnO+dfUbacsca
9eivprmdWGPXR8CLvEMiNeDQUP/hwGTznFx3mtRR1QP+5AEvF42EssQn14ZZILy9
jYKd6ruu94FN+j6IK66p1PHOfj4e1iA1i7ngeP71hpRc3wa8YitORpYeM+oFPAO5
hL9HaZvyEuPpFTsdP6L7ialVWIlWkQW7dOJSmeEhbdOD5GuixC8MIEtXMYe4lfo6
dTBF4fFr81NxAXMEY/8fOgR76xppexKHHJo+UZh4Ucea0swbiM8zcGhABNoQ1mCt
XLaE9y3ch6cyOOGk8gLRs0W1XhoPss2dF+E9KmaUlyWQ67SZmKy73rgxfBGANcxj
WvYzIm4V0lxE3fsK2fvWExldB0ZB41cW/ZuWmow5sQ2jLTmNze5BAWLcih61Gugl
xfmyp0tTmei8Fg+KuTVz79/TcgAR/yaQzknneTvq8ImV3/9lIwaKXg5upbWHFDqg
lGlKWzgy037PZm8VHcw0/rp027JP5SLD2aolMCf/Q78k6jym42yIG+W4K88BECEq
sTIFEt/U0nj7O5OXOk068MyBO+CLbbEGETw4px9x6wm1V34aefFCOOp7btG4gVJZ
bGhYQoe0MM72P03YiKZCFze5qwvI/p047Lev9Wwj9vT6qXfqsS4TOgGYCUjhQxFC
FUKBGP/Dyf0HbKoGXGeV3h1KS1oRj2VTYle9AtxBNzH/KOh7RlYvknP0iG8qjPP1
BEdskkY/jC+pb/F5kTDgkAqLXbT40w81BYUupAFocvZ2meFTa4jexUrHW9r+EFq4
8QGmLOhAT7EQ7ptBkiiYlM5fVW0Vsd272jerbMoOMRawClG40nXCcBXX7jAxBedF
6SLJJyrnIlMzwozOPiFrCge4sVN+0+ZXe365skn5/qQlJ4VId3y9x9ws73CXjgFO
hdW+ThrpQu8gwrJnI+v+qP+VCufVGYN2BfOpiJxzfgN8htyYnxmQ7DfCRve8xmQh
LuzN0DBOpkvi3ZJ3HOA5GWXYYm0rJoLPbm0JSwe6AFUif1dn46baU7BH/DOauk4q
o4loA+4j//XcRda5CRAvr+qHUspmyWo1EsljzLKaXQls9aZayyAeNhcGPIJsoOGA
2f+su4eHOpXsrfCr+kFac3biIRtM2Pi4ARNqmH0tPDba0J6r77byzF11nJAZGPKc
jCoxHFN22jiaZShqViFOGw9+AxduqdqUDzNRGryc3qotwILymlpsmxj6UZ/S/M/y
KTIKomkF3kd6D6wX3uEwS5J31vy1lnafUmfZN5tNCHK2mia22BYgr8nXiIzZp720
XWhIWUgbj3HStOMNqWZN34EL5O61Ip1nuUR5fwPph8vNo/lTLDFVVgR7uZ/poAUJ
RcAsY52Ez6D6iBqbBz9c2zEqc//AWVg624UEdrNFNST1uqIlUBx0itMua1HAMtFI
ZmQOUhf1d5tUqalFFi+socxnZbxb/FfSqxoR3kC8IzEI9nBEV2cdrm1zhkzZr52e
Je89YdR95/UPWnBrNJLb/t10NFPqhHtsriejPiKmUiHEs4bpB5C/xXM/F4P2zzZy
MlgSwxqnFe++bZcUwv6FYkaccXESIw5FM7gJqxz1pIi8C4cgqNBbkewrgHWoGjjv
cwVUm55jsdiuJ4IfJe8RJI+ue3Sqp6DDv5tBtn1VQOFUEfit3rBQYZjO3Xt5+ESf
F7bo1XEJ1HVKQQ5LB15W/xr1JcU/k9zENp1ccLXLxqcvTdrnUP1ZbiSoYCR2udRT
r8m33ZO3hidtFXqGjrVxuL2tNis7qqE2Ohr9UkbyJm/kfgFhHvtzXcggKHB12W29
LprOv6odghbW4b6ViIHlICluyOPIU92nLMUEHH+bJv8+iFwRkbnTmp7nchBdLRzL
WwCo+1aPf3cY8g0SMX28MkNFf6/Uav6BN/BA4Un6Pruz7c4gUOONESZw/x9rCd8N
+NGW+CiP8r5IdJydzaOHa0kyDY0DErnueCxYoFNlXpRiEGciqOG89kyUCb8MwqiO
kHqxutGQY1SXOL34Avaz/KqFYKo17fprBJXmUDaQgOSj9W+ll4LTN/4Kzr4/wuRp
VYRJeL+VRRQudls9OCd0N91Cyk0RO7mN21IauLuD2lmQZGkJqcfoRg9EytZG1sOH
sf0rDP770/UsSAl0reczUV0H/byyOKLUqBC3dQtSufc5wu0oSyG8NgSyuuC9P+RQ
7sPWfs8pBjwfCKy0AQuP6uPjzh05q7qJJUDo/ezVhee/s4UYR4Qyy6/Av3JVwriJ
Fv9eOSGmm+hUbCZQLlo7L4wyYI1mEUtgPDkiF88q9sUWvq2Duj7rY0WFeIUGgOLU
X0FMUSsinVcpBRzVYVzxfP0GeOQaW5j0EogGL+wfzNXeZFvbx760AoLgADsJvp0b
gjPOHokk3xa2t9pOW3nR7ITOnTHN2NO9q5virX9WXjQ0rk0dYsQYpYQLI5EPFHiy
5okkzb3LeLn66a0Hb01//sOI8MG5a/GfYOmOHOQ1WQyq5woDM9B+/T1oDCTpowGq
7bFZ91Gzsj3IpsQD0wYm5MaW7rqiD4S/rCErZvifJdYojF6SE1lPnEAlSp7l1H3m
tCxJ5ViheVcCHCqaVaMSV5lTxNl7MDWv6NeXkMsxxejHATCdF0ytaYh6pLm8LfRN
iSTehLY2MiNxYEZUtgyR5sr+tttf8Ve26uhZrL25NKxIvku39pIelvBGF4Vrhyj2
v2LV85l9XF+kVipc2VsR7OtSss4fGRoHzGIx/JBo+SVQkPDLW6HmquLYwqjS1y9t
N7sl0dogNQCl5eUFvAXwblsIcswLN1zZMtfyAWLoaGoeNtZJbUFfaLZwbT2QXFOs
FKRH9EqbaP8V+ntAUX6ONE3hIdZ4bjBB6OfUJniYR9iBnE1Ej9y73Dg6UWOLkDdF
VtIptuXIidB7wivF+WlCX70HFDgduPq8/CNR88KWjpbMMW8aanFQxCljGnafGLyo
wjjYi5GPK5i1etAOLHu8j+Zh/lef3sum8DzTA5QNyuU7TFvnVm0NkGFyG4DsonMj
d/1ZMQKqc6SSGdG4ojfwOZmGiDzaLbJGYlAUTPy8TuvYTmn2Sj4r6enjK9h4WMIb
bpnQvjNCbwmRRKFNFrIolltoH52VN0y0fnWzBo+yY0+4uwayT29J/8VwSPUPbXz0
CVTQZzEqLpF8oY3Sw/wJtoLCcDTkrfq54cuDXlg3VNRZBuk/r6OsoDfmRLCqTKD4
MXYzy+/EAVnAeqHFpSSHC5Jjo58NizYa3943EjvMqMPb857m1urmbHx/RnjpC8X0
xwlCXCymyAPkFBXwLF4SgOgAeX7TzNteFFn1070Yk7qEDSv7RZ2tQDIaimYyCSBt
K6cB9Z6oiK1OivvAhu2Sf9CmQz/+qogvxRUp5tOQFgQx+eF95wCSB1MVLCE1ZdE9
rfvu9QU9Q/2xMJ9G4AjWqQsLrs8AwJkVbyXdteunFy8Z8mqFy4gdHF6ycWSoRULR
+TVhN9B1KJWyl7R07ZCeiBofHTZuf/8gKvq8FnQdNkbNOOO33VeDqjCgZlZ4UY3A
VyD600XLxlpS1ZemTt8tlhjkQTwmBzzmFQWgOVkKViG6CGR6jBSwg4Ah9/UHGo3p
ZWP9etTlzXOYj6DMTYygsHeteqv3hFG+LFX5t0bAoOq073U9c/HJ2jbfbbphg4An
Uz3m5+BQnUmKlm8kneeLPIrum1K5GgCCB0R22ru2x4m0PmARSaBZ1bxZ6f69EoM0
PY84tN2rs225RQVTQh7cy4t+H1CJ+1RW31wuGnn8Da+h9FzoVhSR5DWZxihrWe5o
6as2XZvbsRQbMQuXvra9Iw9H949emVCeV3juGqN3tV4ZowX8zt6oIX8onKPW52oO
3AGDwDTGRoINhm5oyJOX82Nx3Z+i20L82eAf2X8CxsVUOOeiIAwqxlnEQgNnsTvY
+Mk8t1LpEq8p3+WCHE1O3zUCQjDU5XItF5n3apXDsyD6rif6tyt6/W6ApX4AsAfC
uXljvQxhdHtJaf7NnOO55qHgwZeN/BL1nKLRuOAsM5t8Gq2PHx3XW37LM1T3SJda
BBeV+HnXOxnKnr2rGbPS9VlhwuR1q7TSPIBpI4aU7G9axKVeC2GcXl6J0i/JJDMw
XdPGwzeomp68kSEaQzPb2skwGxqyBBrbAM5fkC86TyzADPFSsqQXv3+InCvm9yiR
RdH1UlNlxFAyI5f9QhKFkuCdsbU5F9j2vrXdMF1p/uRgBDaGudsiVTquCCMZ8N7N
oTYUn2nP1IElUfXUk0HSWG78n1GoYT7d2Ajtf+01CMnmawhoQEb11twh6cyAXJoO
23MZvaFHCvBXuT5k4YFY0u0yx1iNW5+XgXn69WwfSDFuYz0HIghBxMjvOpw6CNFE
Gtr61zp+XskZQTGawjuti3utZGsYHPEeGsqN+s55bIeZ2Dbyfc1IZk2vauZqEbQw
4CxGIJhqfFP4jyP4UmfFrqCFso5SKVgmqaUKZK39HUpuYdY44BFzsR99sZucMLF0
qoP76fqqw9OLt5XHPRbB5bRSCO8EQoN6Qdqth2mbWNbEicL2g03NnpK2W3BjAz4Y
SYAuRmxISrBmrhgkvucUwvVdl1C6YJkN2A/DFwZG7hbLI8B+VHSuqI72APXwrRKs
HTXKChnbJ8qZLYay9PLMRCEShWhpk95364dERMYNENu/y4+lfyCjH7bz4lycsUYW
Rd08yby2runZwhTN6QWnya0a3h2lfRcDaF7AXrZS8+nohMIXj02ot9S6wEPcEckb
hibc43mgXZaYU2K3IKvLRghLZu7MXlV3x6aqkPTqGXfoobE8ci8SAUoiPyercijJ
2d+rZySWDGPIsP7y4rVCPzrSmJbk4F+OAp5yjTVKNRZQ9+XYC1xLnH4RdWPLmCQT
Jr1XoUt6wZNf0NbHqgt9R0DN/7h8XLLXWV5ymvZ6uESg+REXI/cpMjFNVjSgBbb7
Vuk+fM047WLU9Cpq17Xd1h1345/ORxWZxMFuQ9wU4fMeIohRB65zAk7lrogbYNbQ
LfIQXGy7eHnfjFmySDsOhL1Fg3/LUGSdhFlQMzIBDcw5SnPv/3PMDo8ncyNQ/CfO
EqEqoVuaWA+t4s6qezRRO4tych8HnNiDpD+PyEilCn8+QTe1fNH7BqJK6g6QGw/9
ysIhdXWnrBP+qVrJRmxvwa9v+TeYVpLS1iyKQ0EGjTrUkVv2usWXNatbmdjCYN/6
6o9uTp1DL9OBJT2lmv+mN7eiBdGB1JGCyjgoEh1tnW72karviA4ZGO0kET5sb7sg
Ax5w/HW04g4TJDZUbaG6HbwoeoDsb++Ha1n6i6Any5sy94FvyRgWViBO66UJGXfm
VKFJXLKYwliuMqKbwtgD89Mp0XbwDDC7JPY9Y4KIlgOhi2VXi2QpNNKKqwXbMva4
U55Upp5Ix1pJZRqiB8R3Uw9yf2fS/VvANG6j9LqBmyRzJW+OdmqCj9jE1asjVTUJ
Y85uJ61UxFjgrCVjKPSCj5xMlj2mQI21cKgKtPirk4uiwTXBhCcu1R8yO0NSSgkg
9VBwJPnZtquwHhDQDxAuR+Eje40GTTga2ACb4Wo4wg8VXl55H8KMMmSwJVH4bOQn
a2/9TVeVyZCwlu+mpbE9CqyWFVMefc3YfEFV5ipgjsfdgZ/OkCFHCwT4a9wlDJq9
M8IXna9tBhuqid8ChVJLsMY0cs2NwIA4sWh+DPnm3Fh2Bz793IbcNX6rxQqZIhvv
6s5mfbPMxEXO2plnOYa+R7NuQmX1dvto2VrfzJvIa46eJdl53gP6Pl57tOmBf1OO
wYzn9QjKFrJ6einqllLtgk8gBlIHQZeFec/TUMdHQwOszYNEad4fSRgFDYV3BYEm
PR9yBn0p2cB+ZyPBFTvBqaq8LRedBV9Tw6ToDRriRBazXjySSrcyVmracgdOlAjJ
9WO0DwS65m1gPxFAWSiW7R00KuskRyFC69KQ9UHADWcxETriPrhcUUktjiIaw2SG
KiwwYEYzQKEjrdrgu9pDsdAPl3nQ2tWIL5+Olw2dEmQqjlQVEPlm4H4U9hNe+FKN
rMP44cuTT3N35xAmy+4MJ5NruWm1CT+s6r3QFgd9NvSScEwW8fsKSjVjl3YUSZEm
Gpok3PR5IvBvL43qYTxGJoHh+RrqpUdV3vwaibdTr7rWQr6/qR91TgDvBq6WOdU3
201TmcwtBCy9NtYEjW0mvkWMAznlY8PsYtP1KO/i76kRP1sVxu2essKZlvsCT6BM
os03XkHhBHIR4QTy7xfjTJwr0P9FxamujqMrOK8nLd4GFbnTTrV+ebAugPq9ab/6
mG9lcoxzPIS2bodi20DwHLXyzIZR5U9HIHIgS1fDNRR/aDZLMpKPGBlwfiy+qcPN
HoGadf1C+3WBnZjHot19hV2ZR9pTJyLKgdFh6fGp9cO98nFFUfRpmp6NabLCNbcX
ubwDX1ohRTgZZlymUXI87HTCFffsv41f4qErRRQEAwa0kLAPlUdzwpuqfdVZG1Zt
UNghTXeTeStT1vAOpNOIU1foiVTV9m2oajofUNr3Kl/rqvBpU1ig+l/g8tpF1LCI
jQxE7vqkA8v7FZa+XBg62AP5ncXf4ixEMmxJICSdSJIjdqPftRX7zZrSGXIhMHbZ
KXR0IUJX2uywKnydtoYYMjEcBfNMPZSiuk7jzw4m+BeK+l7Fc2eIf760Vk3UxfKc
x6fwEOc8B1dhO0cA6fT1zwPfoi034+PZlc749PgAko7DpPNVeu6V117I3MxBrLy5
9VSx7OEJZUluECWiOeKNssDXX7dzNoQnuFUo2abA+aFcYujS1wrT/kwd+/APqYGD
UUIOtmeBrNk1ryVh9ld7mf4QUUWbXZEj/+krkPtde82CGchRcYj1w6Wg3+3z/NBT
aehq0aYX4bY+3MMFYxjiWYt4Wcuy81nW8uXiFwzrrmcnFtWD6tdu86lv9zeGYbxX
L6ehmc62rLQr2by0DS3xeuFDUSrYsHfLhviqSDvwPlfs3yuEVdKfpGPwKkMI/LPp
fy03eAvbuNqxSLSjmpQh7WA7rjsDbLk+HMMmVvVp7DJASHANGcLxGmvJa9n8sUvj
xsDdeQx0Hhb+UOKyuHoNVj30uZ4RG22r6Awf0g9ewqfEJRMmD7oImjp9F48UJ2qd
+WZCGGWncD5LIuewdWTYCVDV1KsbDudZlOYJbM2OMcIyQ26IyFR4K+AMT9EPvzcM
2KnaXp27fU3cQdV3kUI2/9hKmese4tYtiqfv1aXbmbYqNbpxCxi/9y2QCNd9DFg+
j5lzsDmbxtILBW7Yo0pUYsA6VwaYYB/mwC6jcyFg8LrJLslP+oI8MVA7+95jJ7wE
jPnfBpKuUPEwcnoc1jaXCRaBpcIq6ZuiF77bUzU7J8X4bkwp1mLbcXPiULTnocfp
DxVuRtja8MLOyPt0BDdqIMbt/IaNm6cn9JxEXUgW/csFHOFgS2KuXkH1AuyRUfak
+hFzXOgwWuJuctId0KM0zz6+rcvO8pz2qaWKepILpjq2i+LyHtVOxjgSkIT1Fs77
piV6VXFKkQ0wdJSmSG3PMCn1fLhc8PUdpwfnQRHdF92/iImUYXZLkSu+pnVXCj9n
CkJz/fTq4NMudFF3YfqKeYxRd6HeRIOwnlmUpE4Shr+4+/en3qBlE7q6E8reaCrW
V8fWdFsBW0NgLcFHkPQL5k+EJkG+sOBK8PMNSWrXT/h5I04CpqEA1vcMzHWBCNQ+
28dOg2tjxvfNstNhIK5Xc3SuagrUjaNo90/GNYv6rd/iT3WMXr5u+oMyX/s0nWkB
cJY1E1UhHQUOrtrfOAIu9xS0hNgYqmJsDQtF4s3GkZvEK/Eo6jAXWXP5wX5CJX5g
nTzZoim8ZE0kY+M1k7hlCk7jW4X8DC2lyu0z2PBVR0QQwjbzF82d2Sexm7J4dEt+
B4aUMrQeldrUmG63Kk3MIZXa3d9dRlwcYBBFIGIT2tBGduqH+g7FFLtSgKMFYRw5
+KAhAaRBzaqfgeDzEHio/O8Y/b3CipR6L+FM36ZacZeZ2yY263eGqHC56GGuY8uS
+JrLBq0Byt5lMtAsRWZaqTmSkkUGAqVgLRHS20g9knU3Hb57FrwmBtbe488NQmCg
jOut8WibR7arBlmFwTPylDe22gABFNHNz1FrRydSQ7jVho0tUMZ0w2hy/kI6pu8u
kbvhO+Cpl7aXYEw2QcCAvEhRv0btBivACDH4zBxbGfTtSLkOyb1yoZ2K+W5ORAuu
JLl07VSz+KAJyKCngmz6oOZ6ktl08PNwhsrhrIcNMary0aBtHXD5xeFfjNk0MqPa
XWXZC7J6D+sFwbKNPRNpdimWsZ/LdHIAkRfM3oB4uufB5Hw36425p5tttyAulzyD
j9Jzk6+hma2FHILT73CopHLzkl+gATSkChiZPhjQPckiXPJ24vgvRt8sfwoXSOE1
alOC/KVd720JbKBG1h6m9jewdrXHB71NUj6vkPkp1F3+GUSBr/4H7vqY0qccbYTF
3iXVO1Aw5wZO4BHbDfRRq/14K+fC3U+vSfrckKuXrabCLAPCidu3sgxT/AAdL9uB
8VV5tzX2rySSSZ1gum24Vcj09JFvJjqjx0668EFRMuc47Bxb3CeH6nvu5MfqWQih
LwVdycivfXhUDfdBA+6Idua4IzNQA4RzH2/H2s5fyciUjZj1eWtQU9U22U6/A4tM
3PVA7JSpdPyAVMQp6ivbAttA7egCm/RmhVeL83XvNXNzmvNiSzEy3M7tNVN3opwl
JH9OBhMZtXEAj38hrnT9sBBaQJ8fPTl8pBonkznTIfpxhq3yu2ocP1/qFX64C+o6
NClFeN4zeoyC7cR6yzxCjsaZR+ul9tS0Po6IC1pdsF/lLqRPMkf6b7sMeBeaRdYb
CG+HcI5EZw/Ad2NQd/P42gWcOFgHzMXiBL1HV+mZScMMlRalbh7uZL9T9xXtDhwL
Z4JUYlah0vMWAza1ncklttrsQ5QbXm01H+/Z2jJrEZnzlpYugavC3gc+tUKg9BzL
6mAKD2DtLCN+5w7qigfQdP0vb+fD6Tc7Ri2Mtu7GPQFGHKkaLS+nztBftsk9z3cv
ExHdNLWV6HFi0MLSOyp0BKl/Gz/uto5HOLSG/gGp03hVm8V5U6JBCRvyURCLlXak
v7H6CP1+X8+ex1Lb/vTWiCKc27shnow40vGj7oztLdksDSgDlr/TEZnVKYvfM7Hz
IbMOARzKrdEmmz0j6QUnNCbqGyGGCMPQPLS8mM27ZHiut+G14qRcqsa0PDsEwRvb
gr+D2ao5m/eDk+h2X9GGhczn7Qvos1fbagmiF8bdBr3fHswYkudplj59CnznluHT
lOGJYFmhuYHkGUH6ikDEKhZSseZhQx6E+jYzBbmHqIKLl70u4NqyqSuaXH8HRHgE
hTEztklNtQ6M9oqhSo1f8dOrjzL1YajPzXch4C9Fd9UKLScm5gKtTtKuE61aDgZI
GNLSn9ZTmcmqmguP9BUiYwg/Jn6qB6QXd5TiwPdMHZIunxdvpghvwotB9khvPK9Y
oV/yf4RMDkmyi6ezeVuB+k2aqfJeGg4mFEND9s2QV25wr05Dqvl5cW9KOxrsCChK
/DhYe+Z7zVUJVRIrGQFMpKieM9qnb02N7z+YV/jRVBb4KPaJaXUd9n/z+72i9b/k
0o+XFy9J03HPVhlf39gVsgU/wf3x21g2AO/KsnMsKFVH99uF8jcb5ycGbTKncEEi
xQLa/q0Wd5Hmd1mPjxta20u19mq3m2wD86gLS0I+x3CaLCADUnLSzXzunXzY81lU
RZaXQt5iAKwfU/wlXBvRzA86l8Ms0lXmNlCY58a1zruKCH87IU5kWhhMS3sJTPlt
dVdrJPgnDv7GzEzFjF5F75t5ahiEL+aKudz2VrsIMyUeXPlcS2FyZhIzZT84uC50
XgRMqrfWq9abHsmkG2g1ERDhLkUFfo2AQR37dAh0aE7cMxGjCip/U+dY0NTSuYlc
DduGP80C7ULRK7GV4qbstgQ93xbHormV9NamFgKz5mPC39o6xz6RAke91TwlrlOW
xoAnwdjaOKKCTcpkBWUPBSH1PBXTEka6EpR/li8KKgiOrQCehjYBWWytmoD9rGS8
S1VxlAsw9UE5YMwTpP5tCENATllm4QjfBNA5rEMyHHuXPgvHL4EIoh3G1eHzgJJb
TsbSzXByL5TTtFEmnZTK/WnKnn8Od3Ut4SycX9sbCBXR3gFp7AIvfqotUSClFrmY
NGxbuBw0QiJAjhyT8m5d1NWZ1nnj8yd/STxB2tK7JARWAPdW+7bLckP2SaIpy9J4
eFSavlGA7ccIZm07b7gwWhAw31kJB/Vxhtwm0hCqzQ1TK3kHDhnjumT/8S2wi0cC
3pgFtwSRytEUAiDJ0aAbjuuH3zIHS6cnmPYcWyteAOG3LKG7Gu6ifasUf3hX/0er
xn7I6sECAeBt811rhy9KmPU0EsYuqyR6dtY8mQRxEnx+8BMUeEjx/+CJu1xswcI2
XNYXsLCEbhb7smIIC3gTEfpUiKNAaM6ecSLCgj3UI6eyjW80GiGL8ajTYqRwNfpF
qyBJgLwTXP+KbTaB8LPU9tEtYY2pQ0aRkWAbXAZvtJpDUB2bBYpPHQuLt2kohNIA
D76t8Yr45tRmKwHUiW8K5HqjGGZkkOAcU1ejPXwF3iFjJmrKPxxZ29SNkArPOH6G
pKo+fl9pebH1+kxg42kwMCfzOCrZStSR1cHONU6k7jxiLRWu10w/cTHCH8p7sNNp
xxLOwW+QqcpDNsqWtR7HyQF6JJm9MEL4pitvOlhOeyhzoZN584yw6gSm97jlfoeq
BtGH+cIAxSyMqFW2XNaVu0aBtCEH+3czQ6RR2QWoC0xEXvHbesLb2wUbieLh2yX5
9xtjIPmuo0UDbz0wNhmeQWrl8BYEy0HDr8jGORyAroZu6e78uF3XzVdPbVbcOckm
ZkJqHFXZ6ixz6igbY6NbB8U3fb0bYTU2wrZABuBFccp+vX3VTfZqNodJQuS8HeSx
R+Axvqth+dDemTnxY792QKCvedOtqU3271G2e/+NbSPEIQ3rPpjVujZXGTWScztq
tBeLGdRHQskEuTYecrma3fHLiOxmDlUkHcAUWxvOYNRxaCzK9VXd6UdoRqL1xOJ1
My1aWzwNVmkSytkF780j+TQW/L1I3TpyGfzxQdLb/UZnbG/upZXPsttqR+4+olC7
sp/UlyhQc+tjFP6cUIZFB4TLqpx2apoQWSRja0XK3vW8kyf6bhHDOm8IEL7Wx8xT
Ig4FkgTgRrpngyJqi4eC7vxjZUZvL/sRhwG1MkCQfrdUuLnmadLzFthqMOfnLk4o
ZpGZMZZSKIIrWYBXAtDDPRP7kqNuh3tzWI/BEHR7hp0zAYS9mVheYxmK7jCBYS3R
vXeZHsLWg+U7s7vfcvDuP3rWju7f5+mZl3thGLzQtYLivxlUrxgIBbltKYQcOv5P
oK4LYpgQnVo1g4RsszVx0WsP2gfOT6MoKWwxT1YEMOiv8A1vRmaSrAjTmfM43U0a
qf8oiQD3+vQCfmKtcBvt5QXGBc2+JRXEpztJMf0yWsAwRzFFNpFuwoeoWI59ah9C
F0srQ6bdiTgxXZ9yuT3fNYlHbDDW8OMCgQcq0veOGxKZrfDHp1UoBXntNjnfMO+N
GVap0P30ug/xumnceLOqnIRNoBa1pAd3umpmQ4/SFjiTpJQKmZK7Xe48Fmv9do2+
4917VbVXEltv8EP8lO2Vh1qnRwngfyvCaYMuvzVhaxN7yAXPK9nmdOAcCH820WSj
PLFqBFoWnH5UUcNhH8A4I0B8suy0wcdqmgv553acVCnqVb4chwAmf7x2mfS3t8xm
CyN0Uo2gxnj2bZGXAudQV0N8uKHTTdBmRT3SD9jTDi81WmNrIByJluGYYaASWhX4
R/VvET9enFuXsQyvDB98FeN146XtH4SCQGHKSn0FVn8ci/vFum1jQprbwdT0bbxQ
Y13zj3Lzsrum7jmez1lhwfeZ5FP/lqNEuQeI626bOPyF1MaSa2/OOjMFR6ICU+PF
Hw5wkumC/1grpiBh1yr0bRGOG47lKuOAr2EF7oPQKZoJa/aatkM/YVx5su6Rh/l/
4M9ieUq8q6wdt6bE1jv57jHb2ceheVN3834oX7H7jQC9TTdaEKf/8Wg0ZcTzChf0
78BVRGTg8Qp3C87Rncf5MKE5yOLSc4Tt/BzvTVc3ma1xi3AdtaRiSpx7hi+1BJEB
ZXIjeEYl6Ldy7C0CSKfcGtmYxpAsWixP5h4uKGSW8mtbFtoXBoAC3MkxnLHO8yn3
ATqH3iZ+v3xzS8MTuCV/xsPmDzMQFZiDOZVEwmWIw8s474QmRYg970WVfKLfsTom
tbIbi9/yEQEeXyyfk0YC06b6iPkZuDOOwk41p18TfQQKysO6hUtQmqaXKqH21zZF
ZfjmKpSFfxqaOlojGgE5c0rU9mJxT/pgtuy69MVNi8nesCTSVWh7Ok2XvIzDRYfH
GALq0egMsgOn1NlVR2Gw73CyqASkOlB/8S/jKhPQZ0g/RJ43a/Ww59IpPnWGC5DR
LqkAY6m7EnZU28cwKRwm5g32lDScpi6uG6u72Z/4RDUhgVlJOipQ7NsZtImGzvvP
j58XjBd8/qk4askvLKsrhZWQX/CpENlSAVjB1r8ok2c1wS5SMFP4chrYxmtZxqNR
ctFt2ebxBmCBluJW1/ty9S9ExKI7tu1USgOLYqsfGxxOpmlKziiQosGv9tknhmjh
DuDEqv7l4FoEIOTsfdyjOwqgCs5sOlxACll0sOr7reTCXzm0ckaksJbphXZxpDtS
bC7w2DwRjRjOG9GnC4+yWQqiJVXVQ7CPDHUALgYln+e+qUvDmqp+6BcVYtwKvhrH
/++oaCecsNhhnKs0DfYvxSS6HdS4UsovSMb+O1HtO3wO72jn6oNsb4oH7lQ9uFzX
Yzx0agmRFGrxrvT/OhzZCZPa6jPc7DHcm4JiwSN5TGudVUYzB6lzjFLw1PA0lo80
2fnXjIBHr1lnTGQyivJ0pFE1P32q8mVcnb5Xv0d83qy88DskIGKjGdf+WuMWygqO
Ky2+zWjp0TWpAqhZXJ2NLToRQBK+gnNTOgY/JKJaL+SggciK1+2/Qpj4ofrDSG0/
vSXtPKRqM18Kve6KKJpby5LVTS8RqUTOVsDQhq0GMDBezphMBvojVQCszyi+dGoO
cIkwabTpMPJLYTf6NGtvWWwiSLWUor9ZkBBzwJB6DfGrmA3lPeGYPaM7WcLkQaIV
UcDo5A7PrayxqCmeLQISp949QJS1cTWPqoATYS9v1IaGihll4Zr5PtAymfeVAMMr
e7sn7Iac/fyVAiz9wb/xT9tnyKe2IBT/EzlVRJiTV1l3vXd6/223R+xbIJfW2GDQ
c0pmTFJjpBYjwL/kO61dTaiyU48ivzhdCPUMb3c/Nu/Qyp8rwmI4kPktqNBBb1yq
wVLVt4j1kMi43u7tnFGaMQyIaDQ5H0+9ZMAdpKgr+x/5P+qq+gsxWEMuUQZtWMiD
FxQApWHlwi2SHIcMAhgs43yvEqWHu69FPR9cIMyMtK1z3y6ay3xuhq0rLQUG7XHT
OyQ0T84Kmn68lO/T8fSo0eKHPbvSPzFODeZjOX7G0IULhTD+haN+wztrmkoETLtq
y/AhqkcrdFhUgIMRLclasFpnboHKV499LPmSAltkPhLYZ5BAeHXp7yxty/zlGA58
7TnzNy+9hBfEw8MZ877a5Iu0pGNvrCKULduUfJE/Fiukq68SyFUJQVuODsnNP3Vw
qximcavuDu3zcCQCO7xWilmTGgR+Ax801YzcSM2jTRYToCkjsSNg7yeM2Iqmxcp6
FOZMaVu8RuTnKA2maDLJX+mAP2mOsBZTzwHQU1QNl/swpr5FJfEGJfz4EXQoJW9p
V90QDaZFaNDyLA2Puq4RgZCK3u7OS3XHxhZhzvK12BaqrtX0/WlYKalrbx5klhdg
JoEU+hOy2IS/shuaMdz5oLJyJnYtqd8UXEiRxQT8cwkAy5tH+9SsVDerOjyZAVxQ
c0jaSuZ1YJyvdSKAiWKVQ+zPhUxhHM+/+MEjDic4UJgMlIcebFOLkxpsUBEpA0dt
jexJux1bsWWg/awZeqoWMMtcGal4Iw9vc5231FJAtsqRye4ERf+MMT4nhoTDe+TP
sxoTceEU6g/pCFu8/ch//TLwMO4inNnhgMEmyJaQBhzF8djo3KD1ZTABdMuWrLFu
mJYRCbNdfGx1fQastM0QZTnsKVraDk8AviE/dHQInmAkyl9LwOLZAWby7z4yHcoi
cYLbOChdPXojQB7uZ7cny7EneDl0vODrlLoMK13tsVTqE6hArYfBP/PtURJBBZsL
dL8IYMZNGqpflGXkRGGe2TBp7YHSDhBX3edP/9tQ8hIuEDRzq8+lOYyBMdYk1URL
QRggkOI8tS/sm2v3Pn1Hr6CA8c0rJX1uW6b0Wh2CnhxZ+Ywut74iNyelh79PYQZr
/5CNbocz4qRyjZ5MHknCJWzw2W6NWwMoGba4xii+nKKSurHdpuf9vLaYBlKqhn/j
qRnP0MnF1qeiH6Lo/lSMb+a5Ok/glln9sVcJRaBMrh98WtSI3Y9Zkx2B+OqGAPou
Y7eHwAs0UkhKnQAEvH5k1JuA/DcAwexdGdGsmaDka2EU0Rv6GmHEvX+XZ9YHUt06
ksv0GwT2wDAWrY25vYHKTe5GIQXK4c09S9db6F2FItWIx46TNf6oupKpqlToHE6m
28MBoEM0xK1Qfn9kd1JMmQQZ/zrXdfGQvkQzoL5bl9zbe9heB3Uhi6yh+DSeWh/6
ZeDXT7ALMxADiGBff3l6Yo7eo7WAqg3dyeNqahhsSpFK2XuDC04gY5HCjxF5tIl2
nDP+9KLP7srmDse5/WanXdKdMBJ+btdz8jIu6sc0Fa3JepbJjszieeSQWBDicu00
mLxYgF031PHPozdD1Lr64LSWNe/Q0gLQvuuTuWhcafpjw3rm/2M7+oKMFa2MDhCb
Igo/PSETGByTmU1cAfyCcYJVOxbsAIVr4rKuebsM4k+ZXE2CdzMv9GhfdGVn+1Q8
EhmOW0qF2/2KTAtxRHJODgrQSgcO39m2DZLiVxxOE94/29qrfGLGNbH3ouefhK4O
G6n9MhdNvjvXWlPXakgbrhHObMFhsZM60V2NeF/EHvzK4LRZol3nSxciFUj5ZLgO
mb/q3+t/LoEu+St0gY/17GVxQNS5uwbKlOag8c1iri+ws/iHloZZPsqVnNyYvAZF
2bGNJwTMTWw99MtDm80ZtZ5rihyBpK1W0n6UsNVDTQPqPtyPxrarveGzbAkZ2U2P
zE4JZ95DhHwQLPq175XJg+e84uX1Kgl4kRtb39lMjI2nNUwtGJfr5faArR2n1ziH
ZvyrFWynD4I0GEd/IKWGwAadfSmY8cyRgfpFssuQThSeTNcWxDaERQFfRz5VLrNo
p0MQ+DjXzg9BmfepUCgMQYWUmqcg1MiWh3JlcJ6L/l5J64k+BaIwyTHjYrJ2ACou
Oz4DKh+2i7s9faSfbKYMPIdCGyWHptHrKkprcQ/F9jbOUpLHTM30suEvGTCraRbW
3lC4cwnoWvjxYmyiMs8yWHd3eIlvxDUUftprPzcqWWFXWIAluY46/Kg0caMEhd5B
4z+iIdVfcwRSdL78nuiu028Ebh7GUDdoHvxMpNwHKramH+fALbFmiBUpjhovyHg3
O7qR18ePAS9odJTNuucWeXPNMeuo5tMEg1rvZTFci7m3FI61+ccsMuBmz9VW3QN3
3Fjlk3AkyW/5F+GHGUdteELz6eWaHRg0blYeBV2RmQhTCBWlOdOfsfsuXUWEFc4g
wCeGvs1zYdEGJOdiC655hRA5lPJQ1QhAslOYAQRwUcXizMambO0yvlnZCAdL8Xjs
nYxlj7noYBCFODzttp1+0Ph65hEpIznCS9DGMDpI2S+952iHmbCKW4BNXEsJPkK3
NMzRlJuCOpwbPCpfzKtbX1FjA/j1cn1jYrnOUkoVjhUz3nvWofg718JnftyskDv6
U6xDl7K2PpQp75t7ljVlKNdf6ME5UwX8zH8wMhTahee/zjz9/EkA0lIielIvJPAW
+xjRaMwppLU8pM4RSaBOqdM0+7VjqZ1wsxPJcZrF5cmobRiWTAufVzi98b50wTmU
LreZhqKj/OUIgnHuqMs8DqqYZ9nS0pe73CBsMLKYFLwF6MAQI38cLfW05X0XOKl+
3VQD5rkgC6Q4zdbgh/eSn1rW/mE/mAHNbTz26eYNDK2IzQYzbcXjYgisTw2nvz2r
ISKJ+YDKVeuQRtEBsCyegzDpxKeGT7CZY1wy8Xclr5AAYyQzDD25i3wfkQKGqvyD
DQ3bXr78Csrr+cbvr4kvjl0sl7q7kX4q/g9Mk6CVX+V9Ug4l7nlhakN8XM7ajeU5
nSzPsS781jWM3P3HOfkh8PLx5/Efdlqm8zZGJflT5hTmBKlyDKcdL3XU/4axlX8o
nX57CCf2FwuqM4Dhp+UOZPZ3lz6WYIueIqOdNFa01gVulMVMbNA8BnX7+oMq8Ry7
Y3OZ4LwGK6uqJX14o+DhZrwCvMm3cjOBr2Bo2HNQK0aFWzKIL7X1ChYI1yVUyQNz
6C4/84HWMv/HPgHzGWmyKH352ETZcpnqAr45c+usB7dauPxGF5ke/tECkuLnV7It
eR6mkvFUhJnMa/p4GHudXC/5yN7HDXJi/ECZmZScLC64f0MyFcKlLh95ggX2EWve
pAl0sV1g6hlI3w1s/VQ+xno5tSz+2vwkioyDhQ3KGtr0hJV76fwe73SbObku9kYx
oJzdxQEdJOH7W5Db2fXr+NTwLMeI3JxX7PVvwBOzx67Ee4AR3BmnELEcaYWtPgfD
xebsTAR9T1Y7FPKwpG4AQ6Xmop7JOkggU8g1w8K07CNUrzZ6MenVJkZrlOUBf/gA
cBYAVT2otvsmhpWihO98STPNj5HypeyNHppQprWnjyhCnCeQyp/HPbttm4OlcjRj
R9+C1fEMbLj92VGSwF7hbN+zl1SzKMfqoBZMVWDO8csciZ3g6CgpTrxpwpVP3/S9
tdmF3vWeET1awzZEpF1nzvItf5dmamrVDOKPLFS6wCzUKphQxXahkt5zLeyNqXin
G114Fj9NsvgYNlFA8GKOE0fHhIMD4X5s17eBwGj0U5jgb6bgkVCOAqF+jJAlpN12
14hXsSrMYphj4e2JzTI+uKk4QJYfFfrIfgW2B5PmW0nq7FZflgHQJHUzHb1vI9FI
nNvmkxaU/5X4Ih7sVtFb2MaXeXAgBMSlhCzOtZDdwDIzsN6aW2vx/dTjKJQcrrBe
Urop9NpPjXll7018+WbjLOpXubeGhH+dSX667pCdSjZaRCxiUKjd8QmB6kqm/053
B4DyMSivAo5X95l9s2RE9q95uigzFLpFcDXyLZpw5VFCBLyHYKYOtoZUeNdzvusO
vIZ4tf1ob0oRAGeDFNhGxSigo7NlLDjOHKQ8B+LSBKyhWYlv7O6S3zHhWKnaInPc
gYn+dtADkcrlo0w+KNaToZWxDCTGqUl2NNVCs+Pdr1n7Puyz0YGs3li77k+eCwYM
e1ymwXeudyx/6KADnPObE/fvCUYFyYHJgwbyotkmH5XBOuvwRxcpv7pi3F+alwBW
eBpGhSa84nflclS1yDxinhgGltWYbAynKQAwpBwbAZEiWS/pE7uZe8wWNeMhLspn
bz/I0JPnpfWU4RpBQZ7UVqC3T1R62u4wO/Z0V+Z1erQxGlIkqr/x4SAaN9Ltu9q2
D2znd6Hg6cDLlSeV5zMxZgP1MqC2W0Like0w2/tpLkko4il2tjzVdVtwPZEWDnRy
38cnZQUCWl8Tgmz6Ao7n96mUxP7W7YeVshqzymm//K5cyKlae7dSIP2zEOL4Skyp
/Y7A1hU62GtDRig2VkTU+v28PuIr4H6IrQVX89ujDE2zAHpdY2kx0L1OVRGFf439
DbclEAZQy9yRt4jJmmk4YiMXsF9yDp9Yfi6apevzgHnJLStT47IZfIijldVUC4/o
n7FtbRJQqHMZ1gwG1CZZGgEoDbns79SnWlC16Jw36Isxq9yVjZgOe77jE7U8WFMh
LlTaB8DqjoP0TU9tSk1E1bHj7hLqi1gw7eUZMzz+6jhvVtEdTDOzAueUmA5h9VaP
T4kofJCeiVN9vVhQx9nt09887ekn04fHt/OyZgy9YXoqwIndaVuWAcTd1YTwOema
NtHcRWTR+4MWHoozRdI3p5DDiMFZ2bVV8WY1OTnifIjX5dS5+IACHk9Oqgu79x4J
I0OQjW2g0gYNCRrLKZfqc37shjsxvcI8tUFjEe+W5aSiIk9j+98rq72jE/T4axcH
mGpF+ZBJ2RFBbdWVhzW8JMk4u8aWi3ZNA/gGwO/g2wNeQA7ehUhNDHgYbbhbV1K8
BFwa7qEA6b6N+VaCx2SwIx270AXwBtZ5VQ2LwpxmvhfDu+8EVxCn7V6pdF+vdVn1
otz74FyMqE//UyXtCcmRwO41OsJaaaaxBh4UOQ6jeHWN83YXECo/y4Cc2HzZgS02
o4y15vIgNwaZ94nAIRKGQLRZxnHf1PtQw8s5c9lYRi4MFnl/WaW1mQMLe1MBrfa8
vIWV4SbuI9BJXfwuWSEIe430v4uFLAP/zCfB1keYCROamIl6D4InaFR8gaPj4uzo
Chd1td/2HfG52CInT042ohRGXkreyfxjk+yT/7y6a6a5gofqoBYIpZgnKbmER4q9
SNb8GYgLg045q1eeWbSEN+YIx/YSdbzCFQyOjlars/sApLDhIwSCmmF6FaPGC4sx
jWyMIYLilMT7JFJO9LhnxNpLkF8o+RgMOINUatcm5RNJkZadzzdxBSpD6Rif8y4P
nrOyfNAms9J9mTwxRpK8SWp8MTUqWf1hVHgobpyfSl322OC9gowmV+kGv3ZcS5AS
Cfkb5T0Yl/Dn0mtnBG73hFM5Oe7m1vA/hmMn31JpWbUvqBltTZ6hTXR7LQ0LRc7X
gLeyAbQMxNL8RMZ1VKtLVqtDGBRXWUeKd3DGVjv+44Lo+TrN4uNCeSee5Y0f5f4j
Rba4apvx+AqOp+/x1iibAoiejVTtXlYmb8zL2L+1JFiKtxpOhAKcX2CsF4ojWFtt
ouIhw0OXG4OTRbUTzbSRg/MfVtawNEKNvkQmMOTMo6y5zxwZ9/GzXMnoeW5Vzw7J
FIIbniPizWZOrXJkEFzvcumiZH8ruwbDqJOYYgmQmpKL5YxJ2YK3oVnqEq1mtb+E
Cs3VfKgrqGuy8vnMFXNG3hwG5AZNCAALh/ytDmJipDAk8E3A3IuT1PQe99iAWr7s
itNGeuPR1Ma2WR9CaDNpCnszWkEZpL/Ke8Ji4IdFyfN98rLDBlhjxxbeDgIC+5/L
n/wKjzp/en+b1Kq9LseifVm0bGTL2b8wL/LSFWViu5t9IAdEyOjQbHbZ4xp9fFIp
8sX4a/zdxYX7Dn/mysi+Yb7iVpIQ/e7xXjrOWhA7oT4Ypvxm0NhJYiuX5UjQzs9E
B+ozKDk5CBNhFaAz2VK1J8Amub/Do1A5F3B/1aaY8pwMlZXCRTeFbHLtHHAkgGW1
7vYrKI6uXzc4dZndGZXhdZgaaqaqrL20xy7DohDP1Uhpy3CsqaKNFthNy5EWgy/9
eCFD042Tfezgf2hCeqi6YkH39Dq5mQ6IoUDU2pdvEOzVabKF6GL6fgebW0O/9THl
7phgmOGwbwkmpSBmn/m7VXLtkr1+p6BgF5C21tuvOYqd5vmWLQkTFdQ+sERgNFdf
42f88ln06mIXZ+iGBjzXU9i9j+zgbWqBlkGpfviRortt5Ug0AgpHpKYAwjUa9l37
eQh4jTEvwvZMTtdSV7uWFT4wMhuReqphiUtUPsL1xYne8WWdti8XvjrYCN1SuofK
SgYaTgDHJ6ZWg5w5j99der/Kp5sG6tG0ALyoN+kFwIJXRA2shmSxUFC+y7MXgx3/
HgYVg2ufAtrZNKojA4RFgsOUEpoh3AGGS74+irSG+PkWj8wDVAaWhBjp9yvaDu06
o+27E5/MgIqdow8p2h5DG4qkfPO3Gkpc8utS4CKoLfeRDFSLh69pPJ35oDCcQfIm
MMdHg2uVhLzguJUFRURfuvFp/I1NWnO/CdtDwf2cBBr4JrnuLcP28zVdwSDcA6S9
TZGYmjo8ZrrAStuhclU3BUBQEP8wrbgKLHe2vyRYo3lnct2VQJojBmeP58FtHYLj
ZJGUtA3y/0FT1qDcyU7VRb6kgsBDtaExzR8sB4H2etSJUzUKCr1dRyBwA08Dzx2y
mm2HZLsVKGSI6NCGZpbzarxQklRxZ0O6rlDMDmnZhPpTWUqElof5mVKo/bMqJd2j
kXlhZD+qPKucB4k3QKl4N/99JlcBQUFvgtcXeDCPOilbGYczv3KVSL7HpooMzdpx
1lEgr45jGRdYg6DBVP6NYOTyTN/1qZv2EI1WGHMSasoeSdo6LTMbTJMykEP31Uqj
+KXjtmIkBiruEfjMaMSs2E4zLhPLCAN7mgw1SDz1X8IH5Pr47/NGfdjSTTXsxJpT
bz5N4nKDvsFyVYJeffT3lwnNkOCLFltNNzvsKg34jelU/r8paYepFVC+1F43bFGN
wBWtRKKQlSAwLj5B7oYAQWkTGgVmuXz8XBUUV4sMlfXhePwd5Sz0uVZJuKa3WyKQ
ljHubkjLc5l6qzX5FYoY//NdD/UkXxDMdD17dGfwYVXlgSp+MMWg7W4p9CeYSsdj
/76gCEroOfkKUjOltLk2Phndf1DZmsXZcBVKE11V1d3mXc+CMzH8Gh+Co4DqKHoj
1lBzT/EeEW6vSuWb6Zz8TFPIhzN6Z0aOBFc7T/GvkHyJ9SNnNIr4Vzdt7v7HyS0l
gyu4V9oUZhT6rIKXzcdZ97VkijaPwoT1cz8RIsNr5WTUnIyGDmnFpTyOL0iODNCX
2oarEjZCBsUo2/XmzhA8h/j9xpJBNsOiMIjltNxf3XZIm5rMgeYYuklz2sfPdPpw
E1xeN8QmfEJuUhhiHuf7T12NLgJZirh4VKTq/rLJ0sPh7UDs3OiWo7+Snj/KuGP0
pGQ0OrCCMOl6hn4iCY5s2KX3FIBwrlWu21FTsbMpxCyyV6Pn3w/4ScUbv/q+ZitT
dhj80ZU0ReFY8WmIHrfl20noyRr45KnJoc8OdIgqnLgTbRip46/WRkdUrd5cPmb0
72U7C993ScRJHR21H3j3i65uqAF9MG4NQB76SjDpG1PY57ghO3T+jy4ThU1FFx2f
qF32d9Q+AyWAF5d/mPM/6Y/VLh/tQL0vl1QKT2sE4v41peUXv2En+to6czKJaplH
ebt5eU3XwG+Kjykto+SJPP2D+XHaLcr+Zp4EHnDvcgZsBg/fD7PDzC0co4N9ERZf
7Ym8p16LpLt1Y1bfNqYE+CnJR0X+f12+qmz4tHQcYqvQmogd0n0SkuI2hL02QnOl
AJyQONk6C3iogjntvCBRYKdmwq6dVYiRbBl3E4JdHCjAw51knBffWy0/WYQQ7GZi
G4rIALt1DhWG/X2Fzh0dYWtzTgnWUKiBCMfxQ6rUrygrxdjKr0Dip4cFh3JSUojD
SSZy1C8+HrLtY+k107GRMMtH8qWNNiZD//EnDfAZEhgybypJFQJ/+azInCoMayXT
zCEl4gRMvpaPgMRnuaZ5upOR+/Fn6imyA1LzcKB1eoLT9ShCn6yd4v/tHLcM/lR8
4s22bq5Kx3v+K5nO72yClXxNtXUAxAK2ZMe9MYEGwwN7mh3BRyEFqXj6zUpckdUP
kch0NMVSvR9n7r1/o+FHnIIqb78K5fhQGGPrO+agoStmut4q/ryjCfZ9+t1ChJ1q
Jz6yMI3pPsMH8MrUHhCciATuNZfZe6OAqygw/EnrK/udJ7QW3xkCPZuKFIOEzQKK
ZDBEgx1/KZSrcN9ygHfOkVxSYkXXBIBntWzdTXyopPllSuNjbG20aQigKEz3uJei
dZd/qpzVFfVodsgVYX769QYRGsbYpy+h4HzvPkFF96wW3jowVaH5C1LYpj6+NxJf
9/u4dmLbfEHVpUf28SF5gIgLEm/T4+jPlIr6OIRY+LxY7fiEXT3R5nn28k7kOb5w
GOV9aUuYQl6lxxd677DRZZZrdavrQ9pWRCxT9qb3Vrmm/l5E0I/1jrK0aQlJ7BQk
KX5zcoRt8LlpdnO7qQGjoY3fsL+yzCODQ7pzYUwFrdR2M2XspRtYsFqcWMcc8mGx
hD/Z6AGw8wL570LeCm8QLvhfODzK2KzuyDNlpX9Yzd1yPNt7y2FR02LQ6gZS6ga7
l4KyiTDpHv4lMRfCcvxjHIkFhgZllDePHVfVIHiJfJO/38q+qMJco0XM7xUS5pwM
N6VFQr/zks/ZFhWOrbIVss193Snh6AJnMxJpsINMiwuUPujKMA8nQNY6183PPr0n
CbllgYnFl3/i6twxQQQ2AcwREBHxIETGFef5qleLabsdCAqDoApK1ZrG8HzgMsL6
UD4wB/WqNl0VT5IBno3CFc+LEwxpsU6po5dItVZEetbLDnM6MYvPkoL1BUao4gEN
QqZareZANUz7Geabg9wzVCVXYtU69EIf3mVcsZ3kMuoKV2MHnZ2bnCZjFEzIe2a3
36V4ykgLHs0KqiqH9EBovl/6Hq6G4cYhcBEI1VK6zPGeQ774ZvTHcd/BdexoYlPR
T4mcjE0eMHzG6oUrUX665ozYbrHNRia2+VVj99vkl4zcKuNGdIIAKd7G6ySGPcs1
ukwTBr/wTSw4kstBBR4LkVMbPpfYiuo94rnJZBrZcLvH+FsqYPp5uB6ATw7aOFuq
YQq7wNZAJg4NXjCqjaloy0oMLeYktFqsDI4pcFuF85xRW/tCHIVmBdHuRf7kVSXe
vY7Z2BijcmEtknSsFylsCwzxkkeKE4jq6uSHPoDETRqsEcw5zaWIxILH39wQGVZV
IeKyIAPOPBSlAVGmbj1tFhHms2gDezpqYY5ofXZRgQL9QhdQgxYJX7F5MXdcHaQ4
bhfUv1A2iI6YQ6ta+YzHkov0Iu2ugy1uF1HP4QQI3fUDLs2pHIKjJeg6MLO3hsij
m+JOGz6H6dmO4GIMwgsO5IgEJGyu4LxZyW3ldXKYUaEcUFy5DenLn/XlPtXzWWmC
VJqv+k0DgEiRjFRPK/q/LPlTHhGrSmZmQ9R0AHXMhuLRBVl3Rh9ABM/OAi3O+0+D
pHMT+o/GvjFF85pxmZTmDiNMvNXe8uHZ50FU7uRA4IQTDxlmNVHSgjnwLh+HBbE0
A+JEsAsbay++CkyBMoJ51p1/RkHxgAEbpdzVw6jc/TYVr3ADEcFZv9yp3tUEJ03p
/FQDQ9td8dB+kzu/pNHVrFhWdWBOG84/q2BKwUevFeUoOHDrrl67XhEWwr4SUga8
3H7dlvUg0S1zH5M0Yb3HgTk4ATmYkt/AcaAJqvyUhcFeiKJzfteiHn7DFJOd/cWV
WriXGBcCnZHKI8RvLtlSdwDpSNgYquQjw5cy3ptF7+CgrDZx4+HcSpivUFA+PM/d
kx9bNPAAB7UPPWaI4u41TNSK/L4L2xXapiIWYKVBucL+BLwJZ4fDDo3C0C/gUDtC
FC1ZXoD/odV0TVZeJ+B4Eyp2ANenjHeC99mapvTSiZkwcwm+2nsXCeCDuZ7mFXcg
rJ/SyGjI4yCI1EOgExXyQTf8MZjkh7pOnpAfF5WxM0WzoiRDX3cZuw206baQX35Z
KdXPRy0k8vuqbr/G5ntIRiAl959oPEi1L46OxqPwhbhdC7uoYkyPR+nGuWHbkB5L
WN+AlFgJMgWDNzn7A/V+E1fyegV3ouDFPuMBDde7fNDNp4VZb5z2X6aJhpTwrogf
pbg9x4UEUfR6D8+9SJvOieSPzWpVbVCCJWSQoQRBhhbNgLYQLEk9UwW88mut4mWJ
X88iQu1dXoGl96Yft/RayhzBGGd3gIK/NafIgj0DXMHurGhWKwZ+vAkUkpLBfd4U
mEeswFw86NIWa03cb/crdixRrbPIc8It5i+NLgrgy5LepNtPtWm54QYp/oB7cdZX
4T6YhEnhOeXB+Ux1yhShXTCu8yI65hRVic5hHxQMjtMp507vtGvQVMOznU5CEV3N
l0asFPPmX0KUmI58Vfl+I7KRY+o9FZn8WXlgkZ0vUKTgZQtkXZAlmVrg+vM9sjA7
lDql808MyPTPvH2jlNm8T0fiK0mFw6+DkgKL1EJo4Zd8MH3T7jbUb6vmZFE8rtbN
aAGnDkfQBS1rbEjYTwlk0xfWGwaGbSSJYjrV09F7ma3+FcepYHNzpA5Y6tvCM3Vz
X74oinOeW/qpvR6iaDs4TiWx0Xr3Hkj62bNjayxUbRnot25h3Qjc+PBGa+XGfBVa
7wdGZybJo5lzUXEkslhC0a0J5nv9d7lq78oxhbCQdeaLNpi5Xgmk0sF3m1vRBAtr
11man4khKZfb1OsQ9I4YtB4suUbjsSPSr9OzvPRSYhYgCGqYueXHKbQ9rdS3C0NQ
d+elzlkNSB/uU7Bq76YujdF4h4usr3e47oju+MoXZuQzKByuMZV3Rczy5p+fGhmJ
bku6dWSMog5cF7H2Q1yLm59Aor6/cnK+7PqtHv9dEz67lzW4/qMWK+CpsmT6jB2Z
rwWhL715QoxQQmkKVm7BLAy75kEKBOrCNY5Vdqk0GpeVo1T0V9jBOc17W5yXoRNC
GZdhu4V56eGd9fnt46A6/usU0DHNgjY/wMI8okUvm7hyKzte2Bp5xyRe4GgxXN5y
nwyMcC/xaqvt+AwJcezOeZPAp6qe7764x3UkPNTcGO8HA2tdMztyooD8d0yxw0yh
PUHXzyevOCHS6pQ8MQw44vgxF6HWvpVO4I43NYs3wwKe/zEjW3hcF2bQx0B4vq0/
KWrsNlTfVyoMjgDgtNCywDO0rS3tUpu76DNSUc+2A218MezxdV0SGsig3oTSbN2O
IOM/LY5ma6mVq8ea3RSOlhZCBj7um3STY938PAVbCXe284SHYRcoeiNo9tNilIKG
lCbmsEd3kFQUFTmA0Y1icVM291HSeWpki/tV/QoPBla/tbWpJ80N5gasexHTWUbo
3F83fK7tN+oeOeQWebzp+zP+xUGg/0YQ+248QBPrCLfnE1Jh5SXOKK3hS1CMz2Rk
lyeOHtp84eGGCuqqS0BVK9v5zimd8cDMIkGlDjJwB9Oi9e5BIdebsL4HIJ+VZuYz
hzXaygFK1+lxbNi2gr6dfOpGvsOGN1zh/TgLTGIXF/szlDQ1CFabBYsHdV0hIhS8
wJ2Xg81SkxdiyLa5FVojlEb5mAYxa88MBkxeQk/P3kU4BWucsGV4MzWy8RbQAgBs
85jJQ/t0BHaUHSWL/LuCP8DNZdh1eNgV7cVw25X3BPkeXf5rOEauQ3mo8mQVCGts
jwEnSR3sqfyKNgfK4seqWoX7YCj5ZJBzUjy67G5ms1ra0xdYz0ETuVCVxT0XV39Z
Ec0wgAm3vURjsErGlJGaKh4YpqgrMfRB5KFfNX7w0r1vCketyRepmkzp4dXGBoYS
AppLfP5nPvBCOKLABJnzGHiTwGDu61+mnUe30E6rlsDTx2b7uCp7TbRNsIViw/+/
2ycE8tvCYPp1I7r0EHvreOVxZopvRQ5N5gpWLtJ3uGlOvNf1s8Yq0Skhs9ZILRo0
yOu7nsHTKUfqsQbTdN5ZifVtdgwCz7zPFbfNnkiVSkjd8eP1On9mg8VAcEP39euI
xQSuEI0T/VUP4mKBd0NpWulitzW+WwR1gT8qgz1yRcIG5HrpoyLSnTGsYGcgpZeu
ms9OZZHIpp6Fy9EOuDhIBU3iu9v5+WviiCtiJm1kLrk/oEcJkKGIGZ338hQosK8L
ZswqOwqN0Xfiz5txYTts66PES836j/wiDxc+cwM9UIop2tT1St6wDgm22TA1JxAI
u3zf4suwmMnVUi1m4MYcijrIswK+etPOx52wAacLqyPBrLeuLVPV9ZbV8btmO4bV
Tvl9XuHDG/pju8ZnC6jFQV5uuEokN9CtmCEh8Z9fxMfKiUPCctuVqqQkLKrl4aVd
U7PqzwByDqoOVtprE0Hxeloqh5HcvTcy6JAVdrCucRMTplYwm2xN74+9abVyBNMD
vrY5fZZ3gWmin25mPJX77P/ln207wxS0jY8Nqk4YLZPehZ4fjZiC4HevfqVfkm4d
2XAQ5017KVNZR//DUZPUIfpMmjhRMxDBn4iONp/pqBwfg46xBhOO/Y7omI2+1qGz
5OUvQAcDv2rLcG7IgzaZNCMZPlx/Hn+agpfOxp7W3Qpv7+Tq/SoIkTtzrhr9cWy/
TPojsgfxbkdrzJyuM2oNGicO0nvDhmKXLsIWTeGEtlSBLakcZsTrMC/WPGxFeCJW
ZlXA4E97fmjnxR1oU9aW83EJivI/g1YHUbwDCKeQTIBIiqHAFIWyJcRoAgJL73Gk
36XOhjNzzenl7sZ/YAbGMUPmzvrCwxrP6gsZMfMynEoaVC/lP36sF4VhhMmsiDcA
5DAFHPkIxpWcDXMVvaDf1Pn8TMl8yHAHUZGkjfMGhDLHpJFI7LYfXmc4merqMEkG
fqn6iXjevDBdbeYJKNQVgHu/Ykox299LbEE/xEJgaGb81V943c+QOjnesVoll80L
Ru6E8fV19xzhYgdmLMXFZdlrfyg3UYkjW4lDjkNbT5dOCXAE27lQRc7pZRfYVNyQ
I/eyZmSjOA2XAeMz5CnEO2ceNSGQybu8DrQo1nHImRigMBP/3FRL0FKMRBnFx1XB
Eqd2IApOBY4LiTw8FhbCwMOFBswEy9CSt0k2E4buHmhexe1aGAhgyFugObb9bMjk
Z9FNdXrxwLalfvV/1EVLCHoO904Kk31FBUIlDqyZZR48Lwc8o5+Vv4oqaNzngdRD
a1gThiKy8sMXh6BB7BnPdIj7K4NKIzs3e4vPzJhgN2m2Y1RKecM/g51pw9YiH0Ou
bAYiKBL46K3ODGla2QWJ7frE2R4nRJg/5NZu4jtgdtoi8K7KojZbUehElHs6YLDB
ymLWimDKPbuKjeillsZvuAWKOeZbtKS5bJXN0AC++KUw+b9hzVeqAsu+8skclv4b
PbDAeg1eJhTmAST7q8qwj99iq9qugUeaOokCf9dHwnYL7ZkLL0FhKCwD3uAYylLS
1rfy3sSB5L6uMCuAP6WNqoN0cMh1PrYODNSy73zP2hMxmFeNNRD1Mj9/nQeSydwI
sopTrm+3eZ4yUgUsbbdr7BCTZfOg03xcnk60oQTAGV1pYADo1cbGWIZgZnT9Wx9w
LqWFEHINQEFiuXzRn4H58hYGtOOBV4dsxMPaooZ6SgiqJhbL5VKHTxfx8EEYfDqb
WAYnDdBhyc4CLIooK6lcf/MEz1trB0oOi8j1NnHmBcMwU+Y7TLE2TrwqHOXG8LGP
QEjpaEbpAysQOTnVwN/Vna+ZPRyoqv+/1qQzg3zRkZiTUh+2w3K4UI5HO0+5Bv/O
Ckwteupff2FPLc0WUH8SCRZtWwBrcA6aO52JQr85rbJU27gt3iNA6pKydAuMX+KM
VBwY/YN6s7cOPSzSv07lcQDQmASF2+PJcERFk61FcocZFq1ytlAWY1ruGDz/Pl/l
LtcTqGAYR/v08bRzpCm2mDmsOxT2qMR8/VNSyDPRPo7S7FZ6wy7HPPSa4MLn2OxK
gfU8HVuWB5QB+f8+ZpjxZXb2d6UKBY3ZV/ee+ba6yCJDyXuwC/+IJvsDvQFdf/CE
sPgjzewfLXEXvKTFfwY3XW+KFRc02KdOdgCqgoRBMtG745zvBRWL1b5eO4G6UKF6
opC/QAQr/mBVhE0ygTrD8LCk2vVMB3GomrqROu8Tyj3uShCRPxBNbTsG4dlxZy7Q
SZ8tX7avU6jhUV8kJl9XiUt/obQbft+j9P7b0SRYDNwGstPqzEcRGKBWhlyBhLzo
AHSS1UoTpDfTJkpQIGPA0LYibWWGUXl+wjQS3s6C4vlUT2V8Z2mtCnzvGG5hbufN
L3Pau7yMCcNxvu3gHoIO8rGST2aQxwRb0xK4Zl2wi50ykQSsoCkoJN4/FY05AhSt
SzhuHed3JkWL8umqXMD870l4/RS81vVXu1ABlt568zEi7xlxJEacWA9MtoTrENRg
5JNs0EBFqp6cGx9cnzHhA1cIkrsSx9kZlxVzVIqQboqtUmgY+itHeAyPh5zpW5Z7
RO1rq4oeTjb42DDqr5/6CNztyqabG9nfp7Uq3nj2hNPboiBEVhI7jQ2AaOGYTvyz
VPWzT+SYDDF280HLloGrlV3hCMdSF+1E4liBVsTrEvcwz/ZbPSrjSbCh+jLbkxp1
2+plz9S2AQaY7nwFaEYQo2jQzaDVXCXzzL4M0B8hnLpCzFsP0OW+lNI7nMVkgRag
BkkNpCLmPQHECC+IF1N9YmYTIHvlunxpeY3nzMAunZqTbbk+zBnQPiPH28I+Lizh
Cm1SfPzJxvb13BpIZ10QSpKj8baKVp7bWM7htJvnqH3J2qIr4TUMagPU5Fk4b2xW
hKEGYlJveu1QUObgDIvPJ8kYcnqN/IVOpRx6mxNbXCSPpYAq9Y77Apjv8ASA3XJm
w2J2Hn33CHq6XGwtEBvkz4NKMWkIRAPb72P2sb0qW8wE8Oor2mGhkbKOWOvkIrNL
ZyxNe27Ifwah/dnY6DyxSQIbeZeCDj29tvHsiGv9GeAwd42DQgOZmzU4sQsUYrWy
d9mcss6N+3+adYVAJzg7I8q54u37s4cuLGQRuglBKJ0pMkKj+jPyjryxM5i4p3dg
G+4pDskbrggVnXqV3o2HgzbMWOU/UMgJttQ8zYIyJntBWaPzDE9l2VB6hD4MRz6z
nd1NZokWg9bNUD1NZIZRp9nZEVbIcwO531qHRNffu5p4VMOlHC/8NAATvZDB/5Zh
s3UsZkuKa95LxhbUgDINwG1Fe6ApFS5kiWxEOHffjYTz+9aPLEIzcx17z4NRHY2p
eo9isWfj1wqNmL6BkpBD2nQCG/OKcI0MPyT2iWrR6XJgzK+20P3GUUgNzBYPgOAP
9J4pZSQygWztRO2w2GyfDuz5mUNsOilV/+y7YIMtIIIDFEixfX/Nx6Xflr/XcAIA
wjpC76EA9zWPHqTssouMjsxvcxsrYZw6jHcV1flDDckw0Ffl+1ptgZ/mvsac6mmi
m9dntXUe+NHUzKGy8tA6OLpuzOjBs7nUZaqZYHdqYjrRLg962z6TR6dOVLCPo0T5
a3dWdwNLeyGaOSdbMFP/gOT7gupQ/HpZdK044/EICSuWPS5oyxRdsv4q98MaLIit
WhoSDxrJh+dJ6ycn0RxZEwN/lXP4OzUAQbqmqOg3oz/cJyY7oHABWavV0NwzScwH
wN7AAW+NYCuxsB85DF05jHVn7wHDkD7B9S4e3V3Fkd7qPLXPl03fIDRGFiprmxfk
4FDA3VeG//omKKEgfOBzfM2+kjohbEQRGWc1EqzQdn9bLnkgMCT9IU/OmFbJGexI
/Ow+GU83h1tOPoERvccwmLGHXc+LRiEWft4VQUKcoaeqD+l4hY5oZKXvGRS4Bokc
emUoEb3g3g2CgP8/mqNzHYWs1/xpKdRLU3xmiNENL5NAd7SRsasL3TwEH9tBnqiA
POKR3NTZeS1+Ukscn2yePjSmk/fCMWyqq7M78L8ynDvtLYpi0vppzFIRAHIbchhI
qWH9/Y9YhMTPl83VcBqX1wstcLq4wyCIZhMgCo/VsEQBTeqJQ5eTOnjivrambvny
HQXNJcASxMxjqMENwQ4uJJPaWZj/K7JbzURQdoNDucP+UZtTEDltB1H9jJhZHLsg
+6TxnwducOVQz4/IYQqoutf19nSkPGudLfcz+cJmEYmWxyxBTvngufzO9mMK1tDc
MMSYzJ4E6x+jut9wwVXcjvcNQL6zbNg1w41uSADCxydUQdX+pz5ZmeZAWYnh+rCo
CDrcfsS6XSiba8BqXekzw6webut70OAYb9LO3M4yFv7QQ+9llfcs6hWY6RHlx7FC
SlKdioNRyDKpMzdSOl1xLT/6jSGxvoOZWJ1vnnC+9GI2kgBACjvUy+2e5b0ykVLm
h8YAe50kYy4/kLTYz6Cveb1JdlNkWRo2Ju7D8lMSQQCNsKaCbUdwpKV4FPYTndwj
qu8wq81LmKnU/7+FmXoo/SfrK0pfO2ETQ8DlnsMpsk+0EG/pPiVELLfMkrcF14BM
UAsaPieoTp103Byrog1gGApDzQ2X9SMGGrLF3AgSsR/JqXDMk/Ip36Na85W8Iycg
49pBozrAHmJXdl7ueg8YJ2f0hF8MIGR2t84WBzZpPGB3nNPZd9COjsGaMYN2xgFk
enaYPioT5Qc4d2nPBUhBRlCEw6bOKSxwEWVQ9bAqXnB3KTOIe+Baj/l19ExfEXNF
CW+WEXlXh3vCRhbCc0L/l/P7TOkCHCWd3yfvSWNz8IArEUeNQxFDVtFxQrxNRodr
lO15We3a52X1779TYKLOXapZb+LdEoh/ApeYUlDT1nVEWPEfxtbObCdezwrGTaA+
IKLYDS9z/FbY0N/kjBRv+h/JXwOl5RehO4I5mHG7wsIzrPoia3PZ3wNvOV9uJmF8
TPmBNWK0c0Jd7BvnIeda4DVDmmrFCIbGafp4Iik5VVR/QZgugoqqpWL1jYGcNmrP
cXq+upw6eg3ZLEjtUnfmfx7wcsSyxsAb6iEPhholoPs2aY0gNattplLDZU7ZMEnm
v9IUsWKqlgriOF5JxQAIXFN9ezCelFQ+21bVE/knwr+3ut57lNHu49w0cQ8NZ+xs
Oshga9aH8xB2gh/ZNP5rBeESqN4gStYqN7U+XnI8PcOJhDdh62kNs9/rrjihlW3M
1Ec10Cxk5mPn2GYnj0BAUlG8aZbiBYyu/Qe/LTeFy6NCK6DTN/YGClUGSlZqmfni
AGP7aPppYPrSUtu++bfnL9wMMkAdfxSslOArhexPTwT0TJiirOd4mjD1evd1ABgy
v5fy4uHLXdJCo9BuuXjgv+pjPCWaFC0gzsKvScD2jaP3mvblLrrn0OJiUsmAZZD3
XtSz9aw+133EBl+VxL9Ewhbph+fX+7EloT2PuzN+douVuSoW1s+EaisbAFMhVlkH
Ehd/OWT4TTwhaJ3UPOwtGznjgfgTLz6T7Ir9rU/1Hm29R0ccyRtmWTKm+eU1/sDq
82sEM6GTSRH1Gq1InLzGZU3UmITNabn0liWVjTkr8WrLfmwyXXIX13OKjcK5hkFl
TFEcGUePId1ZhfZWjLORnLPo0Ynhzfm57SStGFL7xtup+gXVIjIckpEobb96nRyF
CI5y2nLPMWwAL6rD3WQ7zti2cW/4q1rfCvZJnLRS3fcfMUehgof0CIZCxMTknk8o
1JdP+EsNF/NCa5cR8rSew5j3gVnbantx3vB36tjWfwGdJ8qIZWaWCzmBRI3C6TWO
yEL5zr8I/tdnt5i2J+ZMIHVPUf9VS3OQ+Oe87Mfw7g7GL6JkolZROkztmXd1rkah
QmfpNM9ZK2Q4eP8osiUFgs5X0MO2ce2r8ErI8YzX2BJH34xDg5VJ2J6V75St96WO
hsKk9ftrqK5ef9QXh4zBVv6dBqfzWsTg2XAKN9OPEWSSQsbY36Rx9EKew+d2m9xV
7xrk82tvlI2SQdWt62KxLHSpPOgzCuZ4C56cmjbfa1eMuKxE7A7R0m6XR/emUPwa
HdhOwOedlyGHl/gwv7lXCMdms0AZ0Ow+nffhRB98juylqyW31/6zVIt2BnkqTJds
6ydeEbQoXCDb44sY1QhUPVFDkelwaPCcR8VdD9QaRKkZGAke6MSNQEeooSsIxLEp
M5BXu6OPqzPkIAYwB6LWawjTVktS2DZGe1V1pYwMwu7eOoiN58JV8SRvrVqGV4qv
OKJ4sTeTeDL1cQoxpZT61kQP2CB1VH/iC6t3vtXU8fYvC3KBBO4CtIY+JiveA7/T
Pktr4nyU8WcnwxspjHjRgQW7emp0PlzugzlffdLk5r36ax7c2+iGmJm9YQqzpkvH
1rTSssqmq7y7sxuzm7oCxut3tsbgfuNTdjMHcimK9a9E5WAUIc1ATfbDATN0XmPa
UAoXLraUV/JmX1/Wp/Cv6h2E3/+jd6CK6tZqJRCf3he3en8VxcXkQE4sh5dk2DiV
8SePoPlCZZiRMRsh6AvdPvsGKUcgYwAqQL9S23Vb54M1MHYJGH72RM3qYLAjLHOo
SMvEN22Be/GtZ4EGYsIJOV6BZ37E2oyISVaIdrPzS4EGS40I0zq4RdNwHocFHnmw
xXZDqMuffxVqQ10iOynC81hBlfCPUvuTZlJgb5rJxHeVlu7hs1MS54oXgCJ3uvxs
aOvCjebWJUYexCaec1PaVwrsZ4TeneeyWidPmu0crGDcvRgO2rF85nnAjoTFZFXF
NwFOwh1UTMezGTUEWMqtpfM3Fgb5e3llDS6G/8hWWXbf/21wRLlnGj31QNuAw6Mz
/tXVidtZRdYvV/njGcfc6Kw6iE3FrO5WBhtC4Qfb9lO6DJwd4cgt3/MMYQDrNTEn
WCYZY6LT/RqhgvDoVlxCwOOLV6dqmnEF9EKaMY8L0mEFLVv0KgwBwYxfrIgDSPOh
yCjpS8gb6jruCuKaLlI0nzhFLV1RmE9wXoxPjdCRGYRs4MX7l/zRMmKRoFeNTEw3
GGC0WOf3cALY7J/DOWgvqKzSQfoAi5Gh187k6bg4SeOMJsg620DxtqG8FiSlgNYR
WaJlPXtwpk5aekG8aD6K3pNuaGRbdlCluxiOKLLJdvfhVbUgyvVy/Nh/6HtShDgl
CQzTDfZbBndX/KFbo/stSHp8566iwEhatE6v2L+2TqltqM3Tn7xZfxbaJ7zrZSU+
UDE/8+QNMk0omcMSWcCqqZ3hKf5mC3ZbEjw8Er1J8e3/4UActaIoY6Zm98IMmwmp
fJCj4LOkJjKUeA3mMTBN/nag7xGPSYOF+h6i/rOoEHBA/U9r76JHAcNQzZ8DuBuM
QoN/z7aWWvpcPfDHvrORmHIMjuP1n7TWlUuQBVJ3yHhKfYNi58aM6Jpdw/w++52y
jEfmOCecuNsxp3rnQNA8nFSftow0an8Mt9+ohuGtmGG0DmB7NWwTIxEzHja4zUc2
5PnFeWLZrdPoLNwOV99ugo8pjNMzHifh5fQZoWHUYiSVCbE/oIjnvAcJVLfZfmH2
vxK21ztmItqllz2Ax8ifUlmQiiqF/1e/1wGnTfLuAqRAdWGqXeaqSohpRsK11U+j
XK/ubbWnx1af6j6zDtTmcU1hnWDb6VOzaJxFVZf8ReiqkkyQBxMCuyStIuECIVDC
jVx131YAHRBmAuD48DNqGgu56AoAlD7V3MXkp83/p9bbVf0f01XlPVpAF7IjuSpr
b7A3Dnw9LsH5OpkKnqGQJRdc5VHu0gsgZRrAclTCowOTvPb8BeRxzdbGEvrX5+ay
qAVNPppV8YhWnsEdES2//ufVm1CLdbSIvsU2i4EUv4eof1fKKlcUNlvArZqvr7Zg
Q87VlT4m/EwW41ZjCAQgXzqX0sSQjqc+Wf5VFNUM3ysNNWC+MxA18w5e1SBTTN/9
CKlysDkTyrR7DHJbxUI7EPTYXCFKnGOBKWe2mwL31zupBeverJlZabdJoRi6dLaA
WncT29+yaJpj5pta2INhLHY2p5t+hTFaOoE3HbMQs5NTRe+thEQ8it4GpZK9a00A
eOG0WLdQcT/CjAp0RgaMEBGZ8DUPtksR708wIDubXWPgSIC5ElMlIRLc4j6QDysu
k8PSs4BeYWigQd4RnAnJ0BwQHZ4nTTroLhcKQsRGxn089krhqhuHSv3VFh9fEwp7
T3HJzU0l0pfyHmYIl+z9TaYo8j2jcNIwjCHZ4SYaAlhLG6te4gZe+aDLdEu1bzbO
i4n1sNjVj3npk8s7XwmgFkqBRDkouNZcuzSvW+I2vUUJzDRqMAfzXXv2wmsWx+/V
UKXSKESwHcKhZiJ/wFBlzjlMHIVt1nuH0xiPeCu0aobeIbPj61cnfYkrHcimVFTH
fsydC8OOInoHicJkWCb81SMKBO6YKvZ9PAmHWfHcGgQU1PIMmkNQjx0apStdtLHR
J1/Px3/DLSGXgG7zSTs1tNURGtOGJursUDf9iK13QfWY/6aP1Ck1WmiTif+yx9hM
YGMk4LqOJ0I2Co9eO64K+CRJx9ByRQa1+5KU/g7nbSFL9RdVLTyxR8OKE71tViWC
b/nvrpOax3RhS5x+xlivRCUILoaBGO92N42MBe8S/QNur3spzf61Nq5svL+96iMB
942v+Ou75W+Mm4hkQonHrda/AOLaMCOxdIciSz31eniXiWLXZM6cn7381p+xFeJO
ibKprQ8Kzj7pPbD00YLRB/i2nhStrdOAzW+7ZOWRyKKZubZgqmcwciSHOPwGSf2g
NxlcUhMdlOUVtnqENjy6bOa+jm+ubHtcoDibGsXsMUHUdbCwPcWjst9+Ar6uh0Vp
RR5qcCja6GfsemYPE9oFf3SmVXSx+yZsBO9T4jVlW+YjlP574uSCc5MgBpy75YbK
5YltVfqhu35FWYpZBu/Oe5sZ8vcN2X11zIedzc8hJrQed5EntRUIVyPMAFX6EArU
Aa7qLAfYoSxwBWjVSKJUOUeUoyveRqC7XHa1zlDfIyaIb4rWcSmEHJeoyhOqYNpx
czlbBLmBR1ALDVUB9kvAXYlgAyqW5x6MfhmeUbJodEsattjDmD3ZrVzqzo/xubJd
E+UpocYgzE/D9P0YaMik+ejFXFa/LX1w21RNz4Ez/maEPSWTan5FpyJGIzmEOpQ+
5y6hghhX+dil/kcwsK5Y6YitdjLlodC3a06DdLf3sZ7qxn3mVVbhRgq+TITankx+
eLqtX1opKMKmsp9CiFmqlVw4e8GNgQavEcqxjwFaQC+yLE6PxmrqsMD2HnNX5fjR
cVlni8ctZD9umAe955WKIgwqmSffHfK3n26BRJHYLu5oT1W8406ieWAA9Ydp0kCN
H3qi3faFoIRaB2isg1bRAvUSQKuzIpnDPD8nk1SF+F9InZz+b/pKmdk7k9FGk2e3
xnXLr8eI+JkU+NfdqPj1KJn02qnLSm0jZzXQVCV9u/D3PdFzMzn0bqrqLh6wKlV8
snaBnDiGeBf7+bneledHQCq75Gna6Xwz2nrwO5+D2nmYnISSbBhn4SAcYgnPmwgZ
1ug7uAjbHc51s0n1ooSMCTn0kcfaITP9vCjrjDjNrm5OVIgfiQODZWfyg8HwrkDj
uglroDk13xOBDtkQMsYFfTJTqKuQ6RWt/6ELCl43FRrh644FJZ1Ssa9lKEwTycjW
dFDhwz+zqdx9mfYqsPUmfyw00QFZQPnlFmOOF7/UkehAXxdyo72ydvSOvoO4GUAi
2bPqfeNADsQ1kXWWyQkjRr1zBmPkjz4C4z/8RqWEt+gnobfxW5NwE3RqfkOzuvQm
0jyULxxjpU1U8g12P+9Ugt8k68N2U/2KKnSR75SQPhz9uAif5rC8UEM5gJ/XFpBL
Oua57u5RlMr27wLhyRCfzkcnCJ3WWYzSsbdl41uRAHPlaIxhoAiQIthSRP7dq07X
7iGv0UYqUbdNaDJloFEt3bzOBznmg8HZhqFtrQk+Mjwnf3lA0S+Rqx+jLibcNbel
e0o+aa4yrWqQP0IZUcl0ExyWFgUgxJm+khAXLLW4bPRPkurVyokNuLNbI+YZAJct
kNl68fn1/bIcdR1uU3iFoeJNZaDEqSGuJsPTTKnLqCcRBp28cwSgIfDt0x/J4/ZV
1gHMNpdKki002glWlapriTcV/IYi0jKURKAYSn2g9sCPURFNWjf+tQBaJVESnorq
d98MqEtJpHhUGKfUCRYx7kPthFIAbrzX7jZRfCNHp3at7NRXLSLiNcP6wpnXYZ1u
+Xo3CRuTfBS2sUkEGrSwCZyULopn3u0DV9wH9F90ORMtgVkTKsVrFeaZQ89JCqVM
Z8yW9AZdYIsdZC8Zfh7j3Iihp1CrAGvLbDEYY0HoejIASvr2f0A2Bh2KSosSfEHm
h60aJemdoCvUpQTnbrBTbk8S3/tAdpuxDsZZYrzfhOyLSNCIya8x/0kniTPQWjPU
DN7BONvqOC0NOIjoiw9ciwXo/wfz2wMuZ7RfI9VnawM17tgmsAQPou2WjC0VUOVo
2xox4dyOmS/AVz7yzHk46EB45bIWh5x73bwPQ0g6XevFY6nojtphglvTnzf4CvcN
CeJaf7rjcGesjr9n6Ozj0Sf3rlwSZYnPrs/um2Wzb50hpR41SBPeoD+tzubCAKM8
qOPFrQlZ/0HzBLRLvYV/zCuhS+bGiZXywEjTNsFDhDdWAI+Snpv+nmRmS0iQurK4
CTpZAvv6QIgp6lRQ7PjW+7Dt8oalMNUfFPClfmlOx8aUWNJv4UhfoE9yVnXAqKy+
M9Achu5tieOEljuHSrFT2yOccGt1wZB0lSTvgM1+0bjzkOGnycLXlUBwBtvEc6k0
oCaJN4chzfURT2OZb9mTA946I4IC7Kwnj2dWByLTIs2qAA/7kt2Q8VRNWlrlMz/9
FZPZGhHSEwQ3kk0bTJKzc0atf0we5dXCSLfSumTwTDwrY8sKSiYiSo3uzrpoHq7q
NJ3QUlJrdkdqInBWfopCFX713u8RJemFb4RZeuz36/H1KZQRPhPoflmqmFcdazgS
vv+VFLiEVwUxerGX1MqopTEQY8zTK/4IJpgwnCUCKWnaKAReT+yjuracW9rGhXqw
0FDCsmORpuZqjjgz13EEKHxhK37rLcmOKg97A9FxbHw1CODT6ctouat0qCNN/QIU
8jwGqTEk/hOA3hjNO6l/B/QMCQoOz22kSOLajM/WUQJycWjYeN1HtJAJ8vSvVEuk
HfbPQXSz6g7EZ54FhyuUMxRZw5Efk4YrIt9ZB45P2nJQE1eKt7YOlIuikxKVI8A+
GTFwy3Gb2Y7oKGe3SCyUvxVnKe5TCm8X5yIx+BpNeSbYaMYN3EvsqKegNPEVjuzN
GTSn9ceW+SUEqapgKCtUOOWA6cGGZm160zOBkf6yotaDu7Qhme5KcNYu/jHdgp91
cYDL1JTEWJ+CMqnsJaYOdqFL6CA75GKap8pM59QiFXj6lwB5b18K1OWxcKZtayca
alyuuSXPLQvlapQr5x64YBVgCW4GxQpjgDtEd3dsMbGswMzFWLDh9M4wBZkLpww8
FHy9tS9+bjiycDB9/oDMHBGdlmj9/Eo+OEpxUHcie0kipE+S8tPF/ZSVqzJeuxjJ
QTKFVx1Z5Y9feNDpqqA6+Rsvc3Lrq9qpRXGRW5iHwyTzAkT9SLggI8MN/aUomZNQ
qsNtvezh/jOI1+jrvUCnJOFBpugrjiAI64ZliB+BEN5I6clrxbTsm0nTqVu4Kust
zIPPxK1M2pz6Yhl9stj68gFC+q6DgMyIKd2dg8owZpBXEn1xvi/2v/tE1+c+zCo3
mLsJD90c0jRi2n1JhdDcfIwxLTTyWwV6DkfQihLCvoW7CuJnYAv5EbthD7xa9aQ1
XPz1JvCBwA8kZPoZVLQMmGyGlr1ndk57QQjhHW9HSb0PvM33JAZHxc2JkqOuLedt
UFb0nmqYFTnJURt2gAVjvD5VAkIVWRfKaVcl3OGds6BuI7qt9HUm3/F79IyyHZU9
hH7gSmATH5h6Bnpl1rfgjA61LZi2FlclVoDN3JH/OkdnX57GQ35Mmvq94kuOakg/
F5U66RVyMN6VhFu74TUKm78E/KHNyyNULLi3n/Z4K20aNJdlShzX/c9Lk1IJ/9D6
GmuJfZi8RClj5uHS59nj+uAYAYBmVe5c1F07epSWzJrXA1xQbztooa1372knmXPp
9RptNx7DOlWgqJOb094Op8Rd+2lpl20Ye4UYvsXJVm0w//YDffT1863sTf5m4Eaa
RR6d6syWvkruOOEg1Sv6zrp1dr0LV49EZnsvWKjAiw0pxEAG/jggTvBDYXu/viju
v95CmSPAPO5ZHtQoQosV1aNPlQ/j2bUMP5sYNqTds9GwJHNggXAkUwyErbo3jukf
Y992pwWJUdAukbYEiLvZeh1Nf/mdRgg9dK7mtbrGhln9fjDw+npNHzTx/QFuHYMi
oj+XU+t/hHxTsPmSUAnoactqnsXxA5j8+GE1F6woQ/InLLx+re1jIPWWQL3qXI6f
FNTGX+ysOTV7BLG6N0WMBwFXAmzOto6kZvFGkzuHZwznl4yH+/YPn3q/tg7Pb7Gf
jmYHe4lTK7SJSJZJOpEqma2ymzyKwK9uH9l5c7HYvrFjW2W+U3ZJdy2CvWRHL2Ki
l7TKPwk6wwI7kdS25kfs+xzc5A3MQ2otoNs55NoKRoMBFjh8HqnBL3w6S8U+gfSm
uk7DdjdJe08a5ASPcYmkGORVrAS5G3eCapyAzYzi1pakZJENy0JAvaoP/DXxhhfD
5g9qBHJLKQEP8sEuwmzmbxukU2QFtrXmuabC3MCG/mQGdwpTGEDVYQkIyGRhjgxJ
VEZreX68RKKt0BzoM7rnjwPtRHUPwLb7be2Xf3Z5+QaLG+o2tIVK26Ofi5VG6oS8
B7HI6Gkgj3A7YJheOKVCihrShKsJPpjf86p+hQuPASLwpy6KcEXLlnu58l4m1lqh
zXmsPQOS+p1u4FHa502iI2C71cdPRzOgv49bRrExPzfklwbl6CWPJLifMRAooPl0
XvzTKYuvovMDZB3/26z2jwgirgg46jj01hWirDeZ32M/y+1TRzvhAAPEnpAfqawi
I6QrfPjVzyVP7k0gCNnB5u+W2M/AKB/1Va/jRG71E314VGVE2d5iS9LahKqo6znN
Q73z09Hh63zKxmYUIz5RxJx60HmeZlBUVUvNgJhAoAUgEiVx9Vg7oKQjmkOliKgB
4I/+rSiAQHljX5Ph0tG2O/kr+Eq2iicGoZYqVUnjJFhXikyYl+Pp1l6/XLn551pQ
M6fwHTTE/2Kk+yIQ2G6AkjuduEHXyyYtMpcgXqSvrCJugrIZTFBLKPhhzGCFpmJ6
n690EEQf1UfGHoa70n8QicTFFyjLGDxJFr+N3iO0ivgJW3sPRmg8lwS4M8A1cIYw
Ahk89QUos3Nm21dR5uzucKwLE0zpUoWRtetpShnFL3Pa6kVASOB2Ykm+C08nGI1O
IQ7VJtGFYWgGTlN4hKSxoGpZcTb03mYHBTC7mLlz5MtKA34JrtsSUSAPVEer49RR
DRuQMQUuuma5vieY+YnOlo6kXhTUE15wyQCIlj0f6Iby76XAbIukOV0jppZ0dEdw
nNRum5fhjAWi10D3uZc2xzBMPNV+CzPseBh83N9CFwJXpwzbN9TFJJbSUnB66ZM0
QhO5e3VFxtZipjXa5hJUFFDyYlT6DLOnBSFAlMDYuc0h5flQLl/wR1jJu4chtnT/
ayKgwzpiR6pS6+gZpPnL08yr63S0ssIcOcI5dWn5l9i4kwbZ7Csv6jOLGrOL2HY9
eco94iWBEXbTSw5innbXXRQazeRqiWkoozhx5iNl7uQAMKAbEIJlEdfafSdtyBWc
aEiyOMRNDmKmJOVwtlIdQ8IUSAHbTvZI9HSmAM2wTe7VEQUXRgMMdrylANjhjbUQ
bPwsCin98KpzsQr42Rb615KxsVPIk0e5c5CRg85joK5pXQTriH5i9ow1jeA1nqE2
rwVIjiwnTdTBowVnpixfN76NJQnthYwxB2cV1TPpEcs1AIk0f6AuWlkPyRveqplj
CNs9yQF1VRElv19F3esC3N3tjNcQH108e+n7TdBBSwc11hJTMq2Wr4wVinnlVZAc
Psirj1F8jnxNs1baGFr+/jj5naRMemLPgfDbIpKnPpHamZytvJ/+5xYQgeMACvJi
fOu/6f+gUtm10d1qooW1olHL1tdSuIps2nxBp8b//+KRd5LM8Ou6qsjviciCnIdV
ci6+HOnewP8vJ6MQFoy/MZKHWnk4v1BpFrxdnrQMYNY9D2oQ6Cy4YhbZh32ai3cQ
wmBPOtuoRoqEUFP30T8OMsOlw6Y1umWSeGoVgHeeJ097iozjRC4KGLouPjcebume
fSBfcwUbMMPVfZOP8RPt/31PhPhoTMa7cLObBaYl36cVUf4WJ1k2/yyeGoCv22Q6
+CKsgCOOJPCKyYoGv3HBZp0nM38TolhtR7vAWkRHD9F4mtvLdFkAetgzIUCThy6f
Un9Z7DYUA5fWAeC8zJH+DYr4Su0AgjGbix8w6xqGajSQFdN502mrI4l4tIXlNinA
lbBKEMVuycMHiUFtXfWVy3M0qA0jAL51tMdyHbfM6DXhsbEkv/4iMUdiEn8//4F/
HlvU9rHQ6/y2TpgVczFHLRwHRqVXOq2gNyg8QxMnyAdstYM7OgVoV8sD1xMYyPeI
JsFSxdRdi59nevgLZ3cdw9V+hixw/T6kSJoK068eylHnGdbhhvzv3RDOTiIj+nP7
uGsogx+AREdBwm8mhGpCP2nE5XF4+mXjCeIZgTwX8ozSyGrhQTDKtpmn5Z8iEQ6R
VL1UD5k7miyKiMfVfzI3qb02+SJXhkf6xI4K/RnL0WXLusRuHtq4Nm/vcu2aD9cK
GL3GudPqgZaCuDCLIRoP+jGkb8yni9eay182V0qoSWm1V0pLtTRS+c0VQ+1L0ZQI
JYzHURLAxRtgSc+6xqabsYE2NIY7LiXjcQIVWys6fI4a2RE524b/5cXOSdn8TrOA
6gi7umSYSr2p0sp6LWQ7ktEfgQwRV1geb7tYgIFIZwJ1w9d7kAGJZK2B/biqrrdf
RbrpmwI4c2A9fBwmqVwEyEUKBdk0KGdTwfUBLa2gh8nxUAmwgEJlvejpF0WZQZS5
oiYULhb0//HJOk2r+6c5lOMaRlXgFjN4vKFe8o4CFN5/KmReMnc9d7JTGL17M+tc
MsaBK2SfilGBMJhK4y8CEkYmAY5IIEDOpc0bM5zAcafpkquLaVsakIh8tHav05Se
/QHeBijlrvZV8Vyrj+iOl3ecmL/biUvFbyXK4TAoGNP1KKnVlqMPg+EtxCT2Kag3
eQexld4eAS8tml/HJxhMugzd3qg5messGast0HNwlIjAtq8oVMK9qnNVOw+Z4V6y
MAggc4ZrT/2eJkNXJdLWMmYTFhJgLync5zGg63SmWYXa8KX7Kry7tXAtxebh4H9Y
ZpFS8lfej+kpwbcxs7I4kwv5I8mHvNeyqz6aeZH3Ka7hav7ZALRgUedLRFpc2qpm
3HVw3bWx/R0G47NMPB+iIlc5s3ABob6A+u44OyYiFUUZ65CbnGhx/arKazr29qhL
S6jz8MBGc8eQIxt1kq5qoDz6RgpyzD1F+ygMrFaDqiGMCo3VozNOuMBLpjjCK0jE
1szcIm18jetnxw5Q52Jn0HTda4vKfeqUOl44cr/QhzTiZCLFxf2j6j0jbx8RTIuD
UX4bt836LXyF0hcArUtNGxkbJ8CWlpfKlEMfzsMr4/lcbaF1fQabZLGSgnyMUSXV
t72fERW5AR3Lhs+qjGyGrjGXBgFge+ocnaQSZC455QQx4DdIY1AeKrlT7j4Gcy14
BUXV/oF4qSOLiSjDe/ASq4eoIvt3mHT+pNHoMFkWNwnzOdg5IDtBR9gUdTDvQlQT
tKs+JZpxDzO2CUGcgIlh45XluSoWN2rkAk6xd71Vm8BnWplU/obx5gBnGqsaC7bR
Yzd6jDKc38h1DiG1snZi0HsmTQrSGBtLpMTlK+Si+WDw67rht5uaXDWV6Ll37rgZ
aAMRPQ7WHCw8uWeamEcabShn5Oghohy77y8VgXCGczL2abt8/8c4Bz4aSQu1ZP31
O8RngQskegWPXegoO+7ijRxRRbFmjYQF/ZaN8unEAM04ClrwcCo2PggAUfvyqRYW
EpI7VSR85aL8LOr2WRIZu58pmYhSZGfPpkUPd3LtUjQzEOiGtmWewuKmW1LK2nYO
yuqoTqfDQEzbffhSaEX5WJbUvGaLmGw+az847Q0MedpwoTjXMJf+n7XKlBoOzeXq
rKP4qzf7LJQ7dIc7+m3jQXoWGz9Uk0CfhixLB6fM+AiRduIT1xbynMk02l78KURT
et5yeSxPR0ew8sccfOczzchI0Ys8lpWLlI3HtOf0xDqL37GKbmi8cbTJ+LYk0Wgj
8YEzFno2Fei4i9j5JVij4Pjhru12edXFyLNtzU64dLnrPkOPjltisHt6z8QXZZHH
0QLP0G4CuQPZzgeIisWiBgj6/zVVsAUxvT3OIMlZTLajWY4N39OwqW6tOR2/wxkf
tbNxIRhGPUDTzb79VXnuSCDenovkQXNsU0KjC0s3KRimO6+FWduAifO6H4HOkZOo
iikx284acLc0LVRuGhyT7Hh/iLMfpbMknyzPpAk9mYk3qD95fXJY7vZnsE/rmoAV
zTPR2HDJe64glYdnPaQaC0Da4EyAX0Lyfqz5gEtBEpezWSR8ycNpDhaQGlu/C2/t
UYXic11jaN2l3b3Xq2ha4JkcgEpCn8cy8AXYmkzwANYSySDrBHO0nKvKQweeTnw6
FIpmVRVNWqItfB/FSyRvG53il0DAAMAnNjtlhAalzsj8um0zxvmcvOejjCT1PHpL
4YocNMD1cgLHpl+iecyHOnry7FoUpW3wKjyWC5zXUUWqtP01CBFW+alvY20QKHPF
/sg95Oql7TVoEngf3b+c7m2iAq52rKfd/BO9sSKCqBaSSN6XLu+mhtMlRqMZWugy
GYCCyfDgNxY2mLJ9bmX5P9wZZPS872/xQTB4szEGbzpB1jNAAOdI+0Xq+PL9YuMK
PaGnhPvhZ2grL4soTRbFdqzhr4cMv69K7ZbpIvZqvfNonLiBP/q67U4Cx2omkRDa
o+1itN5VoOiKdn7adLMPAOEH6+ZAECqhzDei1YKAZ9tDDnyMpRJ8TalDEoRmsfB5
dhQMN7A29G/4Ark1sU6p7HDwpILyDtW/678Ywky9Wft/za5urCfMVkK/lb9f47xM
HfDPKPljFJR/ichRkYoiVAl18+l7Qk+rIYbZ+3cNWj3lO5kXxIDZM9OVJyAtGVCs
EB2ASvdKYphmkIJAic1mbDPJZ2idn0wOzPXgstqby4DNcblqAFeEGd3ubior4aX2
pyzVTNc/wKI7OurGMbJsNQTA6l7+YnZG0Xs3mwGC4n1cW3pco1AGJPbcIe8Nkcjx
1FuZV/rIjSL/fQvKlxVW+V/87sRQdSj4JbINPZmwtLXGW54YhwPymVE8W3FRMUpu
vs4rN8dthGsUgGgYzM0dmo2RBTjIWFiSfJbHYrnXkIcnBjGGIngdDZDuSOT1bAiW
OlMlkXdAvtzXhn9c/MR2Y7AphOm6yZWKOKJ1XrTt3wolsvhcqfxQvpI7wc62oeka
77JkXpHImeK9OvZmX+UpKSm60MnScX9y6LRMD/C5CpQsOQTihkDg5BosDzpcsYiB
4N3MNjN/Ji5KPKbgoa8OO8eXvG7rJ9XxaFEYmFmSoGI45sKyaWcfMo/SNzIiIgzn
2ReN5JQd9M4fPRlFWeyUwt/4hp5HYGsamPnBxVilxQIyzPVgPgT8Jn6vCeHZbXBa
aX/8uxgfsrwtvF9pHweZ8Q6j8cmaCRthezXocSB3NW/Yld1gHq4w54L14zz/j5+S
5DChwKCH8cwKZ4AxrpuI4NbNzcQUX3nid9nMW9fyoPIM7XIHGJFnrD4aIsLTiLYR
DzMFka60VmRGebBVQrADNMMnhRbpsMV8+T+hCu8rq20Bbna/suhmg7iPpE4Kmz16
moyUYahnNnyd/hgjMtS44hJybywJ4wDZ9P9thXrPoGPLmcl41a7y7tA5Wjb4DVGf
fRGm++r2oyAbgMMQuNlRoxNlfYaYMUPv0/xtQ4sYTZDjq1TqJ60HIxdcZqTC5qAO
om0Nzkbk/WvqL10oLsWOernRh1tXZAIgM89DARCk3ahwS/0ueW2krGqiigslO5Xx
S4WNFlM8OKwqqe2RNIn3yU1gBF49L6qxb32gTAnVOm8pvUw7BjCJIUUjx9hxvTOe
6Fr2O7qvS3nG+gOWL77h1O/+gQVBACRH56WyLGjFGhblikbzBTCsCzbgDMGL0J5D
fv6AIR7unwQ3Ch/PKShOwXcJWTRD3NtiFy69qG/xhLMp7Bn6vU9xkQbNSOJ7J1Wj
UD7qO41S//7W2dHyYaGAqhkJpC+MVMy++Z3VUm0GXw5OmxY+q50pAaGLA1991Ymy
2CthIbCQSTcRMnUBidUsVdhwDroEBuf7vCo+nKiwOSllAZ3xezASYyrJcbp+bQmY
JdcCbBi217evC4AF/aC0+U++HJoClAmw8yU08aPUhjQE/2HdhLx9DllpMO231WJ5
n95m/OXa6hAV9Rj8Rp3npeQLRtYt4xaMpetCW7wpHRfAUfqTQK/4Ok+7WgOrHGYj
yCkX4FajHFprYNu8PYD1ptQDMTks9/gWCjvuxEJL4cpl6vLy8ndjB7UkAUUUC9wp
zj5ahKPNQrwiLJzB6JSvqi6OKGsQS99+zz3xVwSmCmNUXqT2tNGNzg5e70N1+dyL
82FtvzBLMu4yIGNrqtQjM6e54fG91bEyL6DHk//hoBrmODXZBaAgPxHTVE0eVrP+
bxKe6xBciNzs29Hgw32zhT6chQZ5JO4L9u/zYcSDhEqp0H/35Lku6NquPthYm3N0
na5uHQXbr2GCiTis1vSDalh/wNDDUQRaMXiLXkoHPpfMXE8yWr4GzcRKOvDMg3Nn
EytwZOVe3vVy3sKhTy2cnM8xOerXEBOM1vfQx39hnQtyHs3BiSJLfxtBU3u2NaGL
O+mtD9Q24KKkoGs3c8kXs2Je+G0rCmFM4t7C25y1jaPtBk4qEdlovzJp1nKeSn1d
Jtar2ywkQ52d50dwRXEUhqAAiJcohiOd7FOfjmEv+3LGt39qVr6vJmhdncLvnSm3
RJx27/TIbRxp/+QFtrIqM8EV/p6kflknGvjhoemZWR5QlLVLXuoNbJIl1pHdLM5s
EGjrjoOZ18DSz5aMR/ztpdzNPNHJyaxbrbLuJHmTttftbRZkq7HFJnV02T7JWC63
ekOq2ssd4hDicgAHz90JzXhQgOQywLjMU0T7SJR7FwCRgAyNWlsgfljpIu/DYxah
pyk6TtN2zcrIxPpdlPTYcFjXo2rYSUIyvuxzsEET5B48ljjz6Sx2N8BaifI2c2aZ
N1CGd0aRlHvtfl2vVIrEVMMqKTDfM7xmDZo0m75mRSeWtjyzR9Eq14Bcvq0+qvaJ
VAdw9w7KjvdxGMO0/l8pirfD0Mx6wJkp719BpoN8W+wn63bFsN7ZguUwdHGNDWLY
Bnvfy5UJkbHnKI6J3Z8Ru2ZINLvqnpkoir6jPEsKvSrpKsSaEFv1RyDIzmmG0fN/
0wXRaiirbk7VMuTnmxdaX1hLb5Htw8hncAoYSclDtphscB/457gubzhHXC2CIU4m
w4wIZp6mQEhDqugmSnn33Mtd76tKMYUfrgUmwZzHrmy6YXRH0iTFjmxmVX9G3ujQ
sPO1msr+3xjOXon+TclRIExEekgBOUXfKbUOzWsn7JnkKb1mP6PZERqjumrPPVVz
eWbsIm0gJqmMxV8knljImn9ZEIzSoMWb3Zpxxnm//UBmsTRKEuntwm39AzDST/k4
wR5Qi3HqIFWvXgIUOTmg1cf5o5PguJix224Au2KQkYMYSPZupvxV1WSR63gn2EKm
Xo+AYdOk4TUzlwQ/tGXLL57Ypv6uYhIbQLgRju1pV8qnCIIS7UTUu4RGFRD8Om40
+z4R944t+rQE68bUoJ9sXq4+8W9LI6zPXB2+MX+sxNjXRX9qTnWl4Od0peZ2qN3t
TxU7gwBefQnL3LtAXPJgxDnT4YaNeJkhuc8Uhan9juUzuhBYwkQ5fAzWR/Kv/tKs
iz/pmA+/TdgY2eSNTVbRBDNIg+AU9qdLgxbJUhe1FQ2um3+yLf2LjzxOjFnUh/gJ
4GiL9bN/xJG75mBa/zU0X2+JbyxoxNYajuZgoVwizDKsqXFIi9x9XsqKMk/R2vV3
LhHYudu/3WdA1IPbwbnGbLhvQ2uzZ9XW6Pkgp7VqEipblXOP7bWMETbAJlzz0UBr
StRc7VLK9afBaEchCYK/mr8cD6wBtwzPdx+Ok4J6yHOlLcrwRUTRKOmlMqnCKKTM
KFelGgZna3VDZM2uzRjEpN1WnzhlRMzFXjQSXvDuV5cVBT/3TZ2KQs1aqW8+HV0n
uVUOEATGHuJ0awvyTrhaZrOvOMTR4PE5pC7q/ZU8oBqR5AcP7uhXlkTgof+4d1K8
4IvEo7T34pVwZOqyOZN7HXYY0oRduf0Yi0ltnF9Oj4dwOWf68QW37O/qP8VYAz0D
XCy4vA4L1RPFMZ8InSvomX5XaYGYNwA6vLAjw64yDvyBGZ8kdIAIH7jS2PI26I90
EfOW6Q22XohZ0qoNz9IQP7YOigygO+ttOiUDWqZGZQT+6IXku+OnJA2I3JGp6n2R
jtyehkwEbgQSS5SEmkELXGNHS3ELRSunjqlYwnvZcF67QUKKIGx9yliyCZIN6RV2
pDenOV2M2FOicEtZdLG9udCOjxvXxFyBeSKVlC4ip3eHuXpVrNF3/Daqjrqt03sk
7FkSzrj07qQsoOs+/FYuSzfHr0hcv0oLeTXj4ZpA+mfBcP+n5vRkoA6l75JKTfGA
hCf43cel+/2HfESJxO/oAbnXZp6NSmMfVWPcaEIcSc5APkwuSwTXjiAwerTokl01
XTvw1mUWfQtFaBo1D6tIXygeCrikdlEfmzTtMlvrhVjkbjVk3L8YYkNcQt+g/y54
mocCvTCKSzU1pJf2IkCvZHzA8eyz5vXMtOZdi+uINptBbQ5Br+CqgH/W2u+Cn1/x
mI/Eoi0gpC0nfOy0sq1AOjc0dhrU1RR48c3v7jqDbkoVPtbo3xa6zqd6r0jOGO6q
hOC6sVqBhN7HZSmh7q0tVl0WuC+eBDo4T77tXc09shnPW6x3fgTsbrfHdHXgdoqm
7IjrNH+mP9j/F24d3bf8Njm0EC2y4VkHYP/lWTrcYjUNnRBbJRkmVIyrQjvi+OI9
LQI/VtLQ6zogZpFwtgW0rQnjWU5enUsac6c3Fl9L74BDOcFNQzENhZ/A0X2JlRLj
i4Js2g6ndBed96rSvCPwnOjj+UfQvTTLBmTTPgxx2/tH5MNbMpGcGeVNOfV22GnY
iwir27QKkgmFAfntGkndVXlcYA+3RuKJhE6SXFcETBt6adeV6LK+fOJAlyiMHzHk
fhAYocrG8ObrQ+C1DdFVzjS2kfD9yEVwEWwbUwiMKESJa+M/uwRi6dyEVPyjq/dI
V8l9Nb9LZVniN5jyGa1quX6MwSgghSaRxDh8+bmCGEJm/e6a7FTSOoSxbFSpmNra
T6lKSY3AZ4TTpLBVGLmP8j1M8FYMFugILT9w7hfBMAY04HXu1D3Hbyqqh6bkwBBv
HXdaKaZUBXwkRceHIUnX9J5Xoz+jHqasU7lOoyoW/HGcafXl/yLCkLnjC3+BfKtp
0aROv1nUo/n8KKuFFliiw/nJitX866lV+n2WHm/NNh62ycY/WZap4LsaXKA2sRTC
zOclcbPGEdgvUmDVhVhGLvNKC70PCwBmeGlqIT8vZhw1uo7VDZMiX/gIY5vHFa+T
0E9eJ4aCPBxjcAM66m5rB1K+4AA8hG5N1wT/DEESE2OPcpsWNOCuvzlqHrvkK0sA
hGliZ59W+2/ACEXi1EpWuyBaxylj0Uk1TAkbj+w9zlZlh3CY8o8Y+GCsWpMfPqzm
M86YmeZf2FlgSRulJKjnqDG4H3Q1orWHddt6LzWPNUMFRwfaMu/2FWQ2mGbQ+vP4
CwZ70kcVeq97RU6P2X7v7FcBWR2X6yJarq7nkUEZQ5y1M728d3RnOxIFFz3/9wuu
aBHOzc3CDdqBIkn3wZPSVqve5c8WZzK3nutAQXK99/57/oYfdlpACoYFRQnOIRj1
9Gf+891Mc9JudUezbrWIN/Vrcw96fP+ZzIaSCVmXKen7a5FGwrC4a7FHPGo5ASv2
cdajr77QQxhMTpbWTf2JdX3vQBOXXbvsXQbD7FZTjdHAupjikmYmtRu66yZcz9+i
STWhSw9AerIlZgahvjgYl8mQisEGi0PhS4MPEIwOvMFjTTqCuctr9yxd1wzUArtH
sAwufhPLAi+JOOf1A+zxiveIUSutRWxRv39hBGMuXuZRQi6A3Riuz6K6O8wMeHYG
6UmDiYs7EK6zXPa6SS02H1DGORFQ0RUbctW+mgFaelcRgyjS5WQsHkCf82wOIoPU
gYnYZqRFlSy9fd44gsqy3gVOMwFO+ynhvJ58QOu7ACIhvAtuApAGs2isb20fDLcm
HkAz2GQ5sFl0WYFaIN9AS5YW4e8R++t/H+jBjfIZi2hrUSVpqVkqLJq/dIwIDctu
L5NJPS4ZRRviesxqPHzQmQ8HWCb4ldnjLugtbA5Cm5NiQh8S4HCk6jHOsFVF8FAe
3bo1n9pmUyVEmUkFvxu1K27YbMChlATvoka9y7vSB/pwoIIWhn9Be07S5tR1Ke/n
tLu2RFaATLMsrzZbccAXo9qi3iVxfCZNfrtd8ziILM+oRIfWS//905/1o0ZYGCMO
leEBmDf4jiYZUAqI/0XAcZtwWNBwZ985xRInEVgGIIB1ouZyAA96KWDhmwOe17la
2XieX6/trDFligvMEmlHLk0DD5vDu3FvvfbIytHYYVgRSgNuGjagDiNVGrWlCwO5
7NZNJJ1HUqDfE2+LdidU0xwRUCKB5YmPLvXnBXY9RE1j2abhOftaCcRh5wF3kRry
bTFS632RacNsWTTu28+C73lA6NQLk5k82iBq2RA9ov03wQDTQWxMFU8bwTysR9uo
rlKVJ97r44NpiL8Ig+YK7hOUxGJAft4SUe9knGRZ3VCvFDT+yHuV2DKqFAvk7Vn3
cnm+AkijZtmomQElpAjJceMdjM6j7LNNJna3PH8+zNCxv4q4H4aAtnbG1yyl+7ff
JnPrB4gXWPrOoIgy56s1O8xSH7VtVkJV/bNU33B4XEFDaT0IX3/0NA2F6VBd++JV
yQsjrjp5PC4KHf+Iv5RCXCgrGT9QJsSZ2LgB+Ud3G1WEIPP+G1xhLZF1UcsV3Wch
8JOE9W5dlbDDf0tQNZKFQx+2dBGapajKCemfnArrKPOCw6OsXp6suj8plN/KSE6c
Z1AuUuXXSVYZgXC0QkumfYSsjmpqTBGa2b/GRPJQikKAU+Rh8wHjxA4lozuVOhzR
GXss6EfS1zdgdLgAASoGUrLOFTFSc6Xia4nowT8u5d8V84k9xyGSkj/2MZS5YFpI
AEYCvEgR+JgAe/lbyrf4z7eqRoBIzKH70yIgRbDqBtGyta6Wlam1CCnv+ja9Zjd6
w7LIqdN+mDuDKRZhwl3yfUofUGzYjwLjSBYD9EziK1LWK2FCgoOLU2KsfJfkyMLw
edT0MXRos/NQdmIHwYeAraa8htf2QDQRn7JtQsnXsiDJzGJUfP701CgMZec5qfwJ
crFxLDuao1wzlKK4by+AEbrZpbcy9N/PmQzs6yQ3sgriSsDwvJ1hKusRV4dlB/ry
wzZW86ggzHMOQ0HVe+OonpAJUM/odJW/fmsC0JngP/vAGdCn3pe0yYWOSLU6Zt+2
kiuZUZAzjVB+kXreOXrI4N3d5WF+7j9muwlCSoISScohdLNKiRIqB33RnSKcR7ke
Xs6UbyZYKlOpr9m/NSssmeI+4EE3mTeGes4o4U0569KsK3ncu0I8qyWu7T5Rc0Ew
cE4Me6wwR8VhwD8s/Z8c8jxa0IeQ9XltIiBGZysTlROFr1rq+Zid+hET9SnOxZSu
Z+J2xu9QN5OIAKCgTOs4TaxAbH41+o+v8BaYZKPGJ2beos6vwyPpUJXwcO3Gk4jd
KFg9OyQC+aIeOdvBC0Z/ut+Upg7xGPM7fyfCMB1VQmtySKk5k0rmHX2ISZxgChgS
e7IZELuoKWpfTnpi1sOy+PfYPThAfMnksrrsqWcvrrBgKDAOy2G7Mcg0+6g3slUM
lWahuYLPNussUGo8Ih1UdJ0vFbl2AMIsscJmG+UV6RqNtx1/+fNjUQCwLv8a2By/
pHecy9YH0zuzLh9spWlmdzyazT30mUlWQGEp6R14UXK7laz22vVLdDWpIi7VLqO9
zw6CdnPmCUzMNfH8Dq2+6oRbjIAHA3X4gujj8CavOO2sJXSsYX4YHdeknQu67nuU
+J1Wab78SSXfXugY6bHgn+/TLPWBprDUNCwwsXIJVtqj3zFbhkVYCJS//e8Thvkr
RVoSdDAC9fLyyHLuuJcPvcm+J5ulMqT9om9n5ODgC5Z5CqJSuGQ3FwbDatIuZMVU
tg4JMa2DYccvwBWNCgNOwmXcPgD5APmNrDhDcau37dXyg51VOsSOyJSBbIBOo4G0
AMgZ7j1rF6Xt6w78SJzjn4Y+PlYGeMZxieSZCidGi7R0EN09ClTJGhFpoKaY6mxy
MK/yItz4HJaX3iTCJyau3cg0dwBbEruUlbCz8DbjgJg6GAZXJJTpZYCehMhf+jWm
vRLvfHyuhqXrqhuWxdOmX8QCcTuyo+ekLJBXLOukejBp7oEsOL2YX7Ygw8S2m6VR
fuJgX0GQREKC9uTM8DbZ9JNU9UFZ0Ar+5sqAhUYMk4cWzQtXYXLAj3jBNHDSWYp/
kr54JQaNyciESwsLSlK3XmHQGCYRkvpuex4K0SOTFxXIVgRVG9f2K0kawzgEyEBE
n0dOmYROZTnWPi7uj2plNeinjaTGdM3dN2scNT37kJknJlYSjJXKy5hhFXsERRRc
DHyB18stzXzx/0BdGVoyBUqXFfmL3JwsG1KF/V/wc+yXbrn3NF2hTtw6Wp5tzBsH
mcv0EW1iBkWcK++Dl1lYfbEDRACs6FojhfacF+CAu3BY5zUnCsTR2h2nLFoDJQox
CJcesOxi2H3n8cPUMTqeekVb67NQGG21K9L/Q+ZzFjhssdyHptwhN553aMx6Okxq
6lW9nkoBB02h+h9aIOPH82xUsRAEmnB3By07ll7bLyKKLpF2vpldWS6DaRS+imRQ
RFcKhrG2s/Pn51emZ7+HjJZepwEuxhPzaDXbGR2D0G9zTivXJ8FY5SpGsEKdlROS
Usm5ehZr5IjToaWPZ2atyAmzUNp4WDIlt1fvkUI1mP15FPPLVcXga3A4y1pKozDB
fYyITXdddLojcmtKDo945lGVeCB2B/iFXEjrEnPJv5+Y/NZnsdTRZEAqjqcVIdcy
kWjhr4FzaZI90N1pg6srUgNrpPyBBPgShDCqma3Wr+J/0kxsXCGaNA3AtTOkYVNb
XDr7XjC3Fg54/vB3Sxt6hvXc5QsnVijrhdogMBIHntMR6bd6sny9EWUY5zmg5cx3
zrPVYYjY+biu1L9s+KtbAAF1G08T5WXR8AMZvj5HFCqdhE3pXP2ns6ZBN1MQP+Iz
4xU9zJIRpLlKdmlrw15rRXi9t01J01IkqvLGgoHPimec/6bWe8rhzPqJRatsHwi2
4fr2M3FDyK26omhXg3t9mBWn8NF/1HW7Cyjv9E+S+SK1hhmWGWl7nKQFZJfQkrEu
icgRNedTSXIyhoGWeqJuHSG0PMqH1wt5qcde/c7JSYT5A20RMkR/uRXYwJmCm1mC
kFkOD34Bo2ZtTS5AuDRbYp2XDWi+q+HP/dH81fauu18CiBH+z3UWRxpzubheaByT
oH8wY+rV9e4K8xnlzDNwtBS0zTZdmqyddA/IYeXBTzyv2xVcvsfv3RLuNV7N9dif
cxH3mXOcXgJusLrNtgdNIuZhzimzmxPx78RCtsScOZbyw0VIPHlSnKftgHVRoxAh
aKLNiHdxuz1O4YPBFDOowgdMCNSXLJPWe5+kvQmw+j2wmIl0tyrTvE07PJs27LqO
mh3r1O3ShZlgrJC/UsXEcNdDbxSeSWGEexnFdbKThrHGCT/xnraUwvv1R+tj0YkW
15bhGm+Nshb1SoKzQrCL/08jb8UbWh87ExvbQ3aQDw+GugkeSBsoZ18ZwfEX2Esq
nS7yjzAdLlls8JkO3t3SNWdus/JzinVxh/DPV/K9uhMxhH5LTDKs0DHBIV6uat5p
aCaTNwMpMMq2rcT3bSD8TuXc64DFoXfB86rv8P1BLXqfj5h/VJksYEIsfoeknFeq
mvnPZqHuW+NFPygExoeo/aviqWanRuBDk752BRa0FstkL7QbtXW5+IH1nc5ri+Y5
nLecE8tx+68mnU5dsyXbdO7e6V1tXJ1Znw8AG3W2idzRkapO/Gye2ebwmuGl99gP
1Pw9btmVpGUhrrdg1JrSoCAD/IQvuLwApK/CmKr4NEUYPs0Y5+ZUiqGbXma4MJUQ
0D5QmWn9Pe/rf9fcfEK87TbFH4KTP3LhqUoZY8S88VYrF2n1miMpOoXAVZg59YKN
hMvUBWoLxSz0MZwY/or/8ktvaPZCRwZhT2SEPD1taiEw55IS44/mwMKHnREBe8Lf
lyBNPEw/7beW4bpjGic5rKMmIDekQxjvKU6v1hh4fiUuTk5Ry4CXiYbbnQHFSypX
UUUE69uWyfN2U6GBWV84GbmTsRg7U945yzKxZ+cblJueeF2W6qEGQucqPfjbZFrQ
7Fx62V4qfWVydCBo2tnV2o/XpmdbFw7cswutP33U4mm3Zgrf9EKTvut6hYFgOk0p
c+E6XQFVjhICeUeP3jsUXBDwNyNvI+vlb3R+VdgkP2CnrUY6VmDoB51Oob2+T+/U
04PBXIb1Xr1LOpa9Z/HheVR6diitBtqWzLRpgocqORdzBXZz28wIPJgYPhfVbl/C
4hBSkqe3UW/adq1hmrJWV51raDpl36PjW0tR9q3pySgr0VDmSTbLhj3LuWvNdfXb
s+m+BUrW43vgXpAxb5hZhhvk5ImiKkXD4k95m7PbhAheylpYYc+KQDsSuWJR1Cf4
RtIZXorChFRcggMvu0TYQlU586qys0XyzXIz1XdzBIhOzX86ya6lJkFSr7tPYPCJ
0a2GF8VJo89J/WNIvLDEd706YCzvznXz4FePtIszQh9UcPr7qnlY+o9HJf9sfU67
9lsBi11Du0VjbWLiyd5104re5gQ8F3l+iccz1jGhIEmtJYSRczLIqF0+nUvkVY2s
h2wsJFF3urUNo80ZW6hSEgmy9fNUni9WXq2/XGinf+FONNRJIN5NgbdHBjViRHKy
cTYGpvWwvQw5iNW3Tr8EwKXMqn7QROqyX3r+DrE0iA9bUVZ6v8jeTxrPMWeHbf7M
bA4JQL+mG0LZ1La0eYu9yDMhuK+9Hc7y+ofk8sUxg8c+htpLDsGo8HPnA2q3hQwI
ukyQu5iTxbFCqUBmWKjezIb+1B5Sqa3XjC6ptMqlcV/Ds56nYPxafhWhctntQ+P8
aERmebPryE4RuFbgzxdKDlQSn4320oXwc/HBEmfRlPixTeU/gVq1ja2Cb7kbvJuB
rlePFZBl4KLOrs4GlCA6HSIq5Rk5z5LX70EQOvTGiSTv+vxEQMrHf8HZN2gTW5Gp
OmwAUwp9cBBUGxQ2zo54+IPAzj/PIc2gGLTwq91gXxhDTpSgUBuqIII3vS6echsX
Z+2ZE5elHQTkXZClaMjcLGWtdddXyyngBtzLetvJYlkEIr2eUAAz3EwyJ47hg7kv
yIEd0rWMQ4/I0eM5+NdRriUNCpaDrCqa1HqgvbWceruI2E4oM+t1d89z4yjXMdz5
MGgoj3blqY3F43+besox8AvrNv5TZ3lUp7ZpDylYBupGiSHNVkY+8aQ5dPuUpJrH
3fRGbRuur1/qIL7vSidNB92lbvhrYECDF0pY/1QhXTR2CJ94/KogP25jo1mZqXY3
uXGcoRAIZId/99xvjoU+pGFuaoIBYIXRgGECjH+Lsf72Yu26BIhQwY+PpJmr9psJ
7TV2oZ1pIKkEMiwM6i9AmZvxiCEiQy/NRLDGWHhrhN0m1AzkV4GijxLGQVM7V/1J
PK7nn0eEhWi1BkEv8dOOMBpUxG8MGgiqwaNGnk15zvqIaMePaovjCrEHstSIvh2c
JSS3Dr40WOYZUNBX11tAn1iWAht6jt72vD53AmIRIr4Tmmyi22XNJTy2guXJnSRP
M+7xpr27CEUOPTT4NWk1Kdrkbp1eer9VbmKQeVXhQVGJkwYDn01iR2ReK1GeDwKz
P/N6AgXWKV1xZ8kBaqoTEcraY/JJHJxE1Nze3hk4FGbHKUSgnz+LUDsHsKehnUck
SasMxNWK1Q9VmxK0Fc0O11emHKyWRDGqtJY1uXuhJTgAzawoc7auaCpVIAKmjQO+
sFl5qmJKXC/MY3C/hlnTqdzvUj1yCXcq62tXejfsDZUEFVa3aDGiYpPdhqf5AtYR
xDa7wh1KtEyhjBts2IZgktpBEW6NV0pjlUCE0Zw2CFAsKh5CQ5kP6MjWwjEcz5hL
QCF39dreC/pqJyXhZkRi6xWFFdVq/LpLQd5Q13EE414T+qPN/txw5XVQpLpoby8R
hVM9LZ8eYAehoazqz0XwWdMr2MRSuiJT5t+KqlNrhXvv1Mt9l9xWA/pBHxXXVcaj
YGD4wGB10Pjt6Mkci3VrwxaTbZR1RAmMxgUF5S/2N8xyCOT5pRjwjNr8J5o+v0l8
LhuMUoXMctdNScBQUQJ+sVCcB9hN3NB9Ki51xY1JM8PR4XCdkxiGqT7Z5/b+1Kdj
wBCwXS4h7PQF/zRKL/PAV3ksTHCXwTi9zHN1JZfH3uHailX8xz4/9W2BH9gMBBMD
4DTJiUbX5/gN0DqU6aIc/jTibtXd63+TkW5I5FwumSNe84Ru7zpSYb7gkdLYFq72
wZ6M9X7nX0xoRGGa+NIhLOmXOgaSPuenXuJGHBu85lwgnE9kAG9u53pu24TzoWsY
l1p//lLuJspoOnQ+ADTV1UE+0J31BLCUK4mT1CwDwR1/2Z1Vd0xVfA6P/57/+ChS
Kg3lOdB5TMlfs0r6Qrkh4IQfQS5Bon17FKZBpvCNCXrh3YP1FWJmu4PiPee7X7HS
+fPuPBZU6csokdf5bLWBDlfl+lJ8Tm90Sh4icB7U0ys68YWvwW0twmnJjoRkYlwh
zp1Bf2SKpJBq+wby43Qe9SbR05pfWcl/VsK+4uWiOBWI2MMHRE7kTie3SdM5vsNO
p7O9M/cTZ2AQH1dMM6CSxfvaMC/bTUNzTNuKLDHMG/p+pEQ4ZaGfBSUzn4pWNGNI
NmxKTF8z+1WAPoGeFzH2wmxcq+LZvGCSqxCVNQs9iBMgZZ32D3ZyBqk1+Z41ULMV
qElB3TaoGk7+OmGWoidlQNYbw5IcjIoboi/oW71jXgiGMLwRN9bOpjc6Khd4/PA/
iwelrx5LRflkl45CmT3EtMX8fYdaclV6KnZJFPdwzrxYZH7iC/N0VIXKjrvIfceb
wnBSM7PhAs5NkXbL5zHntpilkx2FhKKF2Os4nqU5EB4DpAZ2boXahOjJugsuzNMC
Zn14KQLrg0jIAg+Kpp1b0taSQclFeefjYnU3ZqE9tNHlpKdo2+o+m5Uv1BhWMub9
Cm01DBx1FCrcA8WGNYF+uIHQFToL9gJyb3QVUOjItsxmCNA8zj5x6pDO/eCvTkn1
B9T3q2IYhKfLQg4rttR7Uv/1eV8lH/8hUR66vC2IH9F8Pqhsb//ohIpxv5E8U6vO
e+hGZX1pGHbduUkXHaX1b1HbX7iZO7UJ1uyR35g7u/0VV0nHtocJw0le4Xv0XpY5
ytOqKykFecaiV3C9giq8tay7wfjO1T7FOxUGVQggf9T4N4//Xz4aNeRxwnniAHjn
cU+DMqaCJlElqYmrbX/A6+HVCyJyQl4o30aeBhP52zf6J9YZCJSfbVtjR6+eARij
IFt9f/R80iZorvIsSTYe+bgg+Xle6nPcgEXg/5gF3tRPlt/UM8F8WENiXczwxKWK
6XCAVDbFVUnWUKSm27/y9UKrxHwt6SQQ6UmGCsiB4Q4/CEb80mGJlNXbtbNK2eR1
Tx7jXiJDyPcRyYMDOH9OR3u5rpTg82atJ1JIpqTZZ+vq8w7RjVikcB7l37LYkH0i
j3J1OkKVPZgMcNFlFXfdOScXmzSi9A7SOvUjkAdB/AnoR2h6w5dU23Z9gQlkjyND
PF/BgO0eveYp669GVprvcCHW7p0r5wB5hLy9hmc0aDQPTU1ibtuFVhZjY7q946CO
edgT/gkqTnYF4H6uDj+4Cv22mydIpE/KtCtKmzhIy46K+PNM2XtMVwR0y5RHlFjq
WCKGtQOqT7pi6t/Lay2hridh+lUoqqwiE6sg9XJjaVuEVUdUlUfCmDkLQB47MiBT
Fuz0DnMEQfhTyOVe/1t6JVekmYCkwjOwhuzihxppitN5UQ5W7LQ0R5pxkRZiFDzM
QkWhijuXH9X+2bS7s4/iUW+kXiyxdOSJqjaZCBrVP7sUd+SeZ8SHqT38f5WtMlPh
03d7LkSlj1BMM4Q/JDsL93cHc+Fxy7KKxvxw12JJb1ZMPfZq966m8r7HctrcyEBg
KY6nSOxr2LTmSJcH6QcEQJ6vBkHNTtvxok4oOX4ViewHYx9/JIphuc6yMeQ2grvR
3XoQONJ9147qUpWREwqpPTNAbGyEP3T8TtVcjjhM8gL41MNSQIdp7n8+eB3NuO4p
8mqjWv4TpZQTYqbah1PbCSJxCsQzFVMOLRRBYdo0IHenvD4HKZ2bP6FGNYYUI/Sy
CsJqLin+P69Zx2ZoyhtueXXTINtHENWDGA3u7ZcySKoJs8rusChFFZQIVzvV+LDO
jPWpKBY08Zr4sGrtdH7eOLox33k3rlrDq0U7v84ov/oVCZEv9hudctg0Jz6gY9Ek
vIABbpYTxew1s+gTAT+lP8XeAD8h0sLvO6MyKPqoNyXohyXbjljCEcO4E1xouzcz
5Cvs5wFlZyLk9srDMwhENH6oNP5LWIgn3qfKJ19WMRWgq4gm5HfwBZtA8OTg3PUu
YS/FYEQbZZ8Tgfgo55pe8nWVlbYrQ1mmw4fnPilo8IAVrbZPT9odabRWJjPCVqIU
bUBEczlLthFmupjBkRCT4kViH/0oFJ3Qmlk0eaoDS8pI3ofMmgqzauUGuXdchcWV
1Hr5cXJZwUN9c7xCdTtnLiBw2pvFzzZK7vMAVQZDYbwj9+JHSalFYG0G3eGuA7GM
+NWy9tr3RkmwOWwVXPrCQC4RNzjhmqPP2IkHZdj6rWWVJMS2jO+QpACfepj9kCcA
YXTbgnkilz2GM2dTYm7npOHHud748p0/irRXiZVdFB4vH/lCAR2qhG8FFZtuyUoy
WTcFdIZPVAeVqPX7x1OH/bo0mSmt4mMFyg9FLUKPovHSlrPfpDokoGz9lTTf/aXG
KN3TLHEE91TSRhcKipjQaHJPz6vmDvgkS2NTAMTDPZmgmHpM7YGxHASId3aGgnNN
Hede2id2HHNFO+xadDB3ma967SuryJPqlvfeWpH2CLSCgQO18E1f9xNVHXUFHiGK
oTIYGWNgek8q1OOCNmsrRFu/CiQp0c61T6qREJmQbRK7/3A6JUb4tmWh28QKDPdS
JgTpSH4VrPqwWQHmRTikiR82PQUG/y6aRINH9ma2Jb69jD8wL6T+9S/i6UgxyPst
CD3IbDKSM8gkpKbEpCKBRxw+wZxyi/Koa8Y1XBCA0y/ViOeW4XvqBnOGZzZNQPwW
y1G/RCoYcGfu5tEjVT//tcql5GBKd/H3WnUIIeKWLYxZ6Sdlt0p4GjLBWNNVwM9d
NHcDysuDaMq9WhvMxLrQWlz3jstOV6nDJIYQNoEV3BFYsuSKdCBtcXf3pDM7w4L8
61X1hJ8FNdcNkpaZzy5QkI7iMWi42uG5tbo5k6cQcQ+9wKifQFEB1uIvT8ISlhsR
KGCR/5ZgvJ//w9YOL7PUzUbCPBYSOoZaEyzTFa1uge24HLEbY5/FUEMBhHKQ2eYL
zNRkGAKpul6oHzSU7cLQu1uNDMXVwKQxZNDJneQJFNabCye8xgvp42zSnrEhbA/n
HA7x9BjwGvRXse2cFX2dUSNovRaUCIrDMizeYkcOYv1D7abnqHopObstjUEPrr7S
8wgqclPnCDBNF2N2T4SwAZgJr546cS8G1xo5zY71sIH/e0Z4DD0iXeAPNJ6Xv3Ze
C9UxRnfT6zbS4+pASk99exh4OxxgiJZvYwGDx+mhyBdpYI6JtnBdOdjTkfymJKVS
h4qPhghPO3uAn4gFjO0FOB0ONfpNXu1t3XHx5hSkzOESesu5HLigDqpMGvsf3+8k
tCWs/sqnMc0zd/8t9VKkbTntRSX12qhFADSM7KlgGKxlXrmPihWZYyW2I+gmWGqs
0qvL8rR9Ou171uCa2o3fExYnU92qXuNmVtxO4ohXsU0dFaUTZP7hj8oHvB4n5EZ/
H77+T2YvRswE+clSHm5XI7aNzO3QL561H3jk/Oq6xEw/tPM18yHsRCBt7Dy9y4JG
I+liRclfHqJSAKevqyibrflVbX6w4jtrBE6K1Pohn0NdiQVVOxdYbsguvJmcg3Uv
8bZd16rzl9RTCc7nF8nTfz1gHiEhq39fICtD2dkdIlY+owrk1hf8IwkqWohiZzpQ
WeZh+tg/jeGam58mM4ZsrPwPjpLFvqXPDYWxHuSJ5szyzuiydQP0KbbPnrE4ihVJ
0frq/uz5U2GVgsy7TW/R6/kqh0rzFIGPbcWb/LGTSRJPtDONVyalfG1gqzoGtDWS
+xbRVwzZejYyy6yMlSfK5jg3S7FCuCgpbYX8EAybG4veqlDTGAkCvjmq5+R4F0Ml
fBPFqCCkc9n33A6VskS03Otmqi2Pfe+wzGrdnf88kchhRy42fQxiKey/pvZuC67R
rWLFun1QHaIJGGBTU9gbddXXztxoNEBrBzbU+Nh7yDymGfa6daGs+FS14SaqobnI
4qij0ZKALzce3Rgw1hbYXkRShP5kGYfmVxNVyNnZ6vME5KjGbWcoiyhkbiWFrUhG
NDmMS1VQUUP3XG7S0GNIKBEm0XuNciEtvZnormrBYcJUr+rxPRNSEDzS+XYJIQVw
8r9zoF+O2TBYtPFFsQwykeTy/OVYwhpno00DDFpiK2LIKCGIgZBGL9yBHkN5jsCg
ZXcAQiD9X1tKb0k1aCNSNn/Efq9q5O9jyiTO+m0UgjglhaTB/Vuyg2B9FjnK6PzY
vBYriC4/VfkD44GQqx0fV4INEYqpGrl26w4KGNBty9Ioy0L1Q6MrOp7Jk0pmO7gS
01KO4rG5Aj71SyucRuCi6JBBMvADRUaAWQAZgIchGCSmp5/q7krZH+mhIowhrkpP
wXDI9O2M/JXzDP0aFiwXH0xw1zHxf5SyGQ5nBDtAGI6Hwm135eNFK0gcG+kUQJMr
U57dwAuzwD9CnBuryp/EAexk/odgwA7yxK+hA9aAdhLtRoLG6AjzGVYoT0PyQk8a
DwftK2UsFznQyKZPNB8kK5L4my9IWulE/3+8JIw7nLsp73uVzYYOlsJydctkB1u6
KMDt+tOiz/6jVV2wd5CUgR4ppufpMtD8TO+IGel5seAK8KYFA5FDKfgCcf3mRumY
bbyQjouMP+3ACOAuxH/REbR+R2mgLVJeousD5cHONL5KhwZ0aJb4yMCa5dss7bBG
HEb8Ud8ofXlxStHIqelXdOAIdg57Sz/tBlrWHlR1q19yY9Swyg8pJqAUp5kR3F2E
BnWWYf0dbI3rjI1pbq17QtHYI1i/9HcdzsTbb6RyseWEVvBktK3paWB2UZQBEwcB
3ZCs/7JWOCzuaUj6KbZfV4Dx5jraLt6WilFwYzMLzdLeebynRwXCuG8kiV5FYC2g
6eKy1m0Cfhc1l50iXqXOHWKDEytfH4L69WCHwBVmIwVs391yFhzifU31oizdFrmx
no36fgD5VrTaMczUzRVN8xzylhs/KnZExfdGi33FnroI42SHTWdoU+pJPYWs1X4y
85yzOSMCCMbbIFug2lYUEzpjXD59Nfe0x/PCoyM8cySb9HGLcWrgzKXE3OteAcOI
RWHXi04FkYxnO+aEZazQYW+h6FZspzYuRHw9VCi0yfD+Z+Pg+11JL0dJ5LMCdm+E
kjFkFq7bxHSwMISs5sLne5MB7YVF3FyZNABByjz0LCNKGinpnv5tVWja9o7gpl3+
0hgVW0qQJ1m5a4heRdQbvWDCN8YMj6zWodAi2EgNllWcMm5euuc+IMgwQeKAB33k
ojaATugrF9M3PEGb4b2Y06QWFixadHtfDl5C2hd1/5aDlMrFXvX84Px7DRsm8oQI
oG/FGwb+SbDQ2UAVrBbLO+SlQ/LNP/32C62tgSWfiqX6nFJcZI8hszu5OeDI+X1r
apioCxkantyca7Zer1a9Z1vmYq/LlJI6ndImmv8C/7Y45vBxBONAtB1I1udn3ITO
iRcspdBVdRhThdt26rKwrnG0HKLPoRhbKo0yRxfUsOTM1H0ur6MZoa9w2cikACgh
JY2AX/O1sWC62xZ0+LOHVs25N65htetod/afEUliwH2TDxd1/j7BW+LcL+5JSyHi
U4y7O/JNhd8GnI6AXPVoHqMyzWZtzaWp2YHQWudopRaL4519xq61Hk7kzoPpj3Jt
T+EaseTeL+3th7N/qmvWjAk4knWKCAt7zjPBgRo5nOzyMRhGabkX4Qv6oz3J+hKA
BKaOWOxI36kCUJWP++QgCY+lACmmpKeHQWkQd4vv7XmEI9jd+5aOoOSCoMfdtkRe
t0CrK560eRFzldfmnmLSZrObdWyosvQ8ejWNKHx0Yw4UzdrWxLNe+A5wLeoh/qpg
Q6vEvN4n1fbAda5es9eV9RuVg0pGNlhwYu4bFc+/aGey3TMa0P/6nzZ1jVF6nhOa
284C1kskvlTlFhteZvEnv19853fiZSMuUmK5AbrC67pw+XtXpXdKz73coGMvRlcS
jYyMM0S+CGFvVFgXiZGi2hNJhygtU4v/I21FBZ7KbCtmEIqC1lQw5p14O3AD7Wz0
2Y7di/w5AWMOAcHG6jel3ITjtfbE8CsaI9K29ru0ic5L22wcSWmulAMYvR4qtJ1U
XazZLxZ5uOIjP4LZxJe3+n4dcdJBBeJjht9PxFWrTCfEmvDzqaEG662oapB+Aj2i
6R2nAYT2bKvcykChcToqgh4MfY4viepjJ7ay7vE5LXIYDL8D2gl3Sr360zq26jNv
D91h75ULILldlGRk2dniHfm9zQbs86V85nNC1DotXfe9CUWwv8OJwWe4e5Jl14IZ
gfnP+ingdr5ZhGmsPPk08TGHsCTPnfUapiitTB1XZgw2hSemxC4AdVqKZ7UUhf7K
8ELJAlxvE7eWlGq4lKaISgNLNvXqgAqPGr2QjuD2mEACSx5x2jz+U7W9fYTDM8Jd
0RtTt6BuOidB/uQpQSpMG2cHWFt/j2P71obMTP7zydB9LGH3iheMNkEHqrX5IKje
ce5BwaADSxLgvikK0PTsmRR+Wyym21BbSlhyAHba2i9uC/CZdBDPpY7Z/RNYp8JG
TyI2jmD4Pb3M3hPg489ivbyqnFZ8fb6XzBdOVccqcj1hK274ZM5wE3AMXS5g5lCp
NFz8CV+UY/f3DS2X3z0Aer/ZFJeeFiXAEs6r08itU69N55aphwebVw3d726CEUOr
rCXNCknp42EwYdyP4fCewyC3GXTtcGWaaLmXvSPkT79bG2McAERVzeA1/Zfdfpdd
Nc9KC9dMU/ANfLTr708508Wh5XKAm3pb0sA7UGArLnk9jUyRRyBLDesRpw5JL+ux
EKWUxhoUvYz2cFE8FXzLLEdlavHXuE0R13ePaHT8bkPR3d9hjX8KUtsdL8s2E/KD
sQm7OphXic1ufM1ujts4Q+zRLFwB6gcQEvbt7lRUkW/QVXw7C4Q78IMTmokKyw93
vXZLTUtaN9FHOp7G/LbCCHr5ONgp3nQoqrBioducZT2IYEbrgGj4JrzhHJY7v/bZ
q8btxwumRXOeY+BWYCqUbvF1+HwbnqcFCfaGc4mwn52rcRBSnSsTcbzpc2mt4KaH
xNApcK5PwQ9gsyfXVnsKwi2lqdD4WeIy46Q9OcJWOWtE+hDq71wJTFFyvv6CttSD
yizv2SSVSXDMYKQK+SIsZUeOT90dCNz8TpF5bmAKBBoK201ZpamYdSF+TakHLgEm
UTjmNzWSEiCY/9wKVOzU00QJx5FDDMxddFBWOSq1WBN/wvwCJfcLWV6vGthkQzEM
QAhTsFhpxtJpNh8koW8ESbi75+KtoYdzyTUBaC6oiBeNFI0/oZOSO7DPQSoc597J
pTcoh/1MEWnyHjzpQyOjiQ2GJG1e/ONRmZt+ldN0bqbxe3fWQkaWFBDLO0AV1fKl
sZBRIBlxnYjRqZqWfxg5WGEPrqiUzvrqSTyTDMLde4J5sK/keT+YflcxKeggsO3R
VORAzb3LCYmwfqOKhbGAVRUAWbH1f8s+MOp+xTC75tbA0grsJT/Ty/bE895c+/pA
coq+r90Ibszg11FgZpAqqk0rG6vYOMSfAlF1jb/GWVgm0SRNWmTy6fmJpK+wB4kq
phDh0ur9SGiCEPIwpk155yFKDQicMffjwNPxzzaaKYnWtpFD3S6M83c345IQpfP6
pE4ECXZn9FmmCZZean1Hep/JYS1Fz9a2UYONapJo/OA3hjrL7V5XXiTN72DflSL7
jziXoJrwobvKvgdnmAPlU3F+K0pZ/htINybCJvbd+KAwVG74WGwJ2thfz6nAJXsq
xfMt6WEWE1YtyUc3UyQEpcxrUNFpEQfQkQdcgDFuSWwx4V7ySPRFQAXvGRHWErWu
iL1ubDyg7gj4yRoRZ5k38IbfmkLmmnuyQTksUXGflVZvgNE/OUEmJBPlLoFWmtZM
gYM8qeFpqiCA1ABgxoEdxLMCTLaHLO0mQM+xY856/VavoM/z94PNJ4Jq6DNVKXUw
hXdAdTr5fTDjYbCl6ofTdWyn15l0q1BzGhoHErbpRZJ6LiCysMZemBQKECXnewsx
y0dF1SgSJQuGskBPYsV67qi2nBUPV2ReM9UdfzL227rTXozBH922PBmHY8mu/g7k
nKKcG32z8+FIjqSaD7p4yN6GwBAlZ5AwaoIvtAUwDnuHaBZ7dadlgMoHAtYVm3qM
JMKLFTID87aBVhQuCFaVUcs9iJHWCBHB10xu9sUc1eQcgRWALmtDuMqbzMwOa4GF
zDvIbLhGLjGC4k4zgAKn31YvUdHp5qo/rJFY9t3bEOA7NxSEUvFT1Kx6l88Ck9JJ
Mp9N/46PHKf20N97oA+vZ7okaZijZ2Nu04jOug7JH7H/UaBJQOuNDVEfuuZgQRFY
g1K1xE+bhOmRGWZc319CABWqrU0clCYZ9EDAqISS+2eYOTob0JMLOYkWKFKnYlpg
198AvArBKmqRQiib//449fIKjNVCsxzR/XZz7g14ikQBa24zEDhexRrOgyzCObcw
ycn0CKS7TIkT+RAbe/csHMCynvMSduANPoNlDvkQs68l4nQBugOoRuHh2kcoba09
UVVpDMxt7YxY7lAPOPv0id+/HCAe6ER0s9gWZ0hwtngoDIFLW8Vq6P14b0V6ZeWF
5EIbt0RCM1v4UV6gwqhFFXchnFBEgwiNWPOL3sjAuOGaIMcnTLwABjem+0uZamhQ
F/coLnJmLpqKO82P2uq7NF+Ackyj+v47oSc3jtEinb4mmpVuswOT3mhvcWIHTzJN
nlpBm41qo1QQ5pxzi2MVOqVVYGBGi/99uByTPVDgXMLy+D3ZwCHtd79g6J98i4+D
jkHjf+CmqOx5BgSXHheOXgZ/QZUF/ajkU9LxdAwPzkCYI7jcTxW6e7CzWqyb91Y/
9xeqctPNvK0NTAH1L9qipI3RrUAM8SPmiSNHEigQ9yPXMuFUHY5XfRvsSK2ccwiR
Ru4fG5u+MLQ92y626slk+ENJUJ6MM/HoB3sQdOOH25gFWX+FreydH255AfG+/x81
Nojeh6bmWwwf8xIbz8akHzHPblBTJnwsHjVxfT30kntI93IPXTBhAQ3hkOESyNyy
LkoFGE8V9yOeeyhw544LuvmJ20UhGlgPpYP1f2JVqEtG4cw6DfjE+MEE9NqnP15R
cDHbD42oyCJ4TexbwpLrneOqj12Rxgy36bYDSFZLq+Oz4kc9Z03w4sx2hk0eNy9O
Obr6aphtRW8gI9fIoFJ8oDhfaUMwZ0H+P0ooBoOipcBf9nhOZh33/eMKK50oGHt7
zGjwpn94SskhmuLvd8fahOCdCP2DSICHTsbN3+Nw8+J7Y5dkmPH0Uc8WlNk1+PM8
n4jzNYAg7AVQjxMQ9krg8YM2s0Ho/3be6D55Px3fFDwiMN0o8KrqvCOYs+lqoE/U
LRyXjLfQXxyWpjjdrd9mObzFsahyLSUDMANYBGWJi4YoS16Lt5IY4wwTJapu8jlb
rBQep2C/f6xhvReI7LP3Qwp3+L/gWDatXdFLik5FLAQjGsThyNK/jXhLeyZVVWnO
a1DU2Ur0LEqjpVB0JPjKFYFpfbRM/RBsFbMI1/Fd1i2TITIEqgl+2iWEQ4lYA7lK
d5gpVbPJQnI3iX/wsXghfKe47+BpXZZf/noFsGqNIb8OtHzRGFGVc6aV9dVyXgRX
sU3k7JwSAeZnxSXO1YfIFnX+waqGxgAVA2eH05Pa99nwaX/V3bMnd5px8GsXafrz
fjEdb9SQRrmvS5RzicWWis0kTigq2DX4cV5yZOv0hVkUDbDYI03UZp3KpavwCbkV
vYgsYlfzUwldf/F7QgpqGAh1ut2VLtMUfNwGRlcBItslnSVXKaCEIVAg76bptL2/
aFjlxvJmRb7yWuFxcsGelT8qhpNZ+XYidmcf8FZz9TB9Wew7AhS+cdWc2t6x45R+
EWmIbhTJSTciIpV39gEU2ZA6DtWWXFm9q/yzlw+NYi3Ri1H7dC4wJw8c3aYr4hW1
Pj9wampwnxzK4V6QZ3o2gUhqXHYsgShraEqgvAMuPEwjyKdWH1nB47tA+N7v40jQ
n7er8aX8PhzkSfRTZBuf+We1QUVHxrSuuzfzBtgAYjRgwkfkAMWo+8+QYy2lHh4F
ewpAqQkPbN+Bz71g6LAxHllzpKV83zfD8waqzjcTeENPiyhCj+tb4WWBjRYXS7Q/
27tyY5BmDWbrfLWtKvxR547UzyPrf/GfshbDQWM1AsA8QGWO7iQaX/+5AE9nw2UM
3Jb78IW45LT+nymU+P350V+qHQt+LsvyRa331FwC68pCyAbIQN3aPoMdcceX/rWA
k0qTykewcPCRR2+HXStLcLqUR98kPIOYG7q9JU59bBxr8n0tD1h47r98yKqXFWfL
T3yw3EzJ2aJLY+N+jg/p1gpEEKGdapX73EtmzExLIGmhsbac4gLE4DG/wOPjEKyS
bSwjoeOt6Lfv6HwDrbAkJDARC1meUsEpIKiCHK5tD4u6JrS93eIVISms3FHiLJ1m
yePrb9ovRQUF4fmLh8lCNHf6wgWIxsllS5eJ5aSy0A0fv0lnZKPxuLuO7rZQeZ9j
WYHGKkvU7CdflYPm+ysc4c6xQ3DSneBOx+T8LEZHfPsmiS/1FJU9nOX6QxXmu0fD
JQ+RovlevzuijBqvnHhMM6pGz1liyFxNC5K6DIs0d57LrC3KI44g+bulBZbbfogb
aIMrPY94CrupMRbNvbxOJX6TvfmrxFr4YniRDWzNEpvjSu5VrHEXB5cqdrbcAJOS
aO5ddEoo1amjuk2UF2AvzA3+5VgleAVAY1/B4sV17FlCBvvqKyr9xf67k79R46/5
XTpClpzjsLED9tZOHmAReiq7BxRqXQ2mAJxk7N5xLELBtUHSaEbLvY4Mo07A3eOm
TS+FkV9kR+NnLyt36h4LwsEBB+66cJS+s+9j+z87FLevB3ZjZJOemFuJk60kBE/3
obzxktqKp8vVQ6HEn1o22JaSgu+Sd03+bv630hcRinS5PS1GnqHPrpWV3m2RyvM0
dOMZ6LkH6ZgOeMCMIuK9fdhU18fPNX79gLyhWh/Da0Ceka5phBXR7w+yHROJ67KZ
1K/Ad5Yt3svB5ThDpeU63n+nL0jiDhLfKOtWMINtLsPm9CBrzDPkbhzTQua2VjVk
fw+LbFt88iMdksS2CamyOqCTzdcY4TJeYhmNU1FTL61AYntjFVnjXp3b/e+ca1u5
/S/9Tfjkwum8GSHvEWKNs877MV48Yvdt8hsdy4ZRp0Lf12CJhnhu+ad1ctTi3aic
+sUf2MP5mmP5wZL2KRndWeMSCvYsyvSZhIm0X6A657eG4m0NYtmnVp8ZJm53iB0o
TzdhCgbtA6t4KzD/BB/96HKdwzzGCAlyEPxiHhYTwyP0xmsif8rrRXDoT4V1Q4Bj
Qk1bVaEjn8ijgUmrpBaG88ojTf+H5PpmXfBx8htQkC9lcwaDNMc69OY0yslX1zWI
6P5FrqdPluIX4xYwzmQKB1OpeD8QQPLHmJaz9RGc3gYVdUoeEDZlAtiIim0WsnGw
61fFo6Hfiv3WiYBq41oNyIBQZCdEhPCZLrAxiDkFa/ANPxJ1cdK1jM5wChdf9m5x
hlEMTxLyLmd4tCIzLAR2vCd422RkeIXaPwQhcSr2hZ4Ul0UAbiiLUVxW3IcqakT9
IquHPobStI318rZ8wUTJkKnKxy51pYOxpJwp3Pv9QJab3js20UfEzRbvkOk2/JuB
X+ihT80NPGjslGPz4E0EWbwhPrON7mEXVRDWHKjqzINe0xRVKKlEhkPbk0gVAjEU
yLAzrHDC3YS/tGx3cfv42Eaxg9S1vZEdh0KVHF6KRmK8yFhN/tmKEGVP2ub1JniA
WZno3rtBcoXPsvIGZs9SKzMwTfhgeN9CxKG8bj52Ij3VfxxKL7/TWqNm1PsH7fun
R0T3azlVEw4xb/4DzPW214EVgP2ZYyLCiGPVbgRmU11f0hBEDdEYt1+vtW9VKuic
xsDyO3evx5uC2ZnQ8dS2TLJdsfpHP37JWdFrms5IMYzucTOd+wHH/OhNm0aH3na4
l7vvHhStDp8b7hZ95aqyYxy2Jzj+OZ45zG44rpzHy7XRoNQobtqvX5vDCPBlYerp
Ca8Eazzwk7ezESbyV36RSK8O8jxwNXaor/Dm5/vPfGcMSThk7bDx48DlNFocgJXU
cm/DQO/NmRxUfFk5Bn6f1Ux3RfRCYnuJfF/TgENcHy5QA7uM65GH/f6kZ3i/IHCn
C2QYuc7NEbe4znVHaJ6TU8rpDp2bGyLEZfsw7InVzELtqzKmEDuC3qJwKWW0Bf+U
a9n1gvgNcoPyY3JlVMZD905uSoRQZPXhVXn+d5Fpc0uPF8USwKs/Nh3GyQOJnhNT
STEC15CXReBCv7de2lKwa4xKlrh/rUtrF94Ly59BOGcef7SxJAjdOYIadxb0MJXy
Ri//z6xtSObbzGIBwWEYOMsQhL1xSDl7hbEU9Wrc9Ab8dTWNO13OI3VDlWuYk4ky
Nqe/UnolvC/2RRYEyOwV8WXFUO0MYBWJpsYalD/qbNBQSrMLErl7etp/C8xTaZhH
C8riDi1bVTPIwGqGW1FmiH0pB2wHjudslZnl07NBUMPaDoUQCv0f85jXxl9oGY9K
tlc3IVGxNfqDaWyEkS7QN1sUJczh/nl4DyZGStzupcEZcBTZSD7C0RHTAVHuaVOR
5sjebcoc2oBcvZbJ7GEGh76OUSsdU0m20/f8p13yH0g5RccGxv8yl02U3v5rLrCT
bJjiSLixz0QmQHYDgK2ASk7QWC1hJIgpDEDqE/LhHw/Ufr1C7x4PTX1kJ3q1KOEd
DoOonGhtgC+USX4q+J1v8bMVDj/ootNKhJJJZDv9ViU6nX7w6rj7is/YsJTST60g
5UB2CeFHmLxtrjXy21NmIlRhYLg0PcOrqhly0T6dSfwhEStmtLMRQaMwTke640cW
C3FCMYtTkLGPs9Ky1OJM9gMyIuNqSjK+pxvp/OGdUJfKoKsVgzh8ZB7AW5ye6y18
GjlqHbJd66bC++Wks9/p9vkwzIieGMEo3gai846NnVx+r+cO/GbYsK2VVr+gAY0K
NV8mbcxzhDC0LjsKSh1a+Lvpv5i6HIP7bbJqE6NS4OnV1Msz97PHBm1fyC6p9HNk
t8zkojb4VsTdTynj7/bCTVFcaZnd17kFeD7MvW/oup0jf+7g4BJFnWfN4a223r3I
7doswYdj59f1vC7fxLKbZJz/dSu3S1XXL9mkBNWMI5e1+PHxNMgAgf/2qWMjO2Mv
7SFqOeKcLpwSISydBut+whjLSfYyse/8rl36hnCeSes6SzBwwyhBBjQdL8355uhx
DHMH+VxI7nsay9hclCyy23i+ducSWyTloXfNqEo7b/2mHezNQuh5Bdu2Wgl7NFwl
1xBgNLI8mBelZ8a+SRASNIP+HVe4UGXTXA+UpOpsVoYMJgP9H5ij+RNKFmpB+kVY
t5cf1Ne8Qcomq9oPyQ56/N0MbLiOgqAZc8ruIha8PuCfiLAVEcIOeBly0redzFOe
q4ghO7BEB3CWwjkgFbJg5uDqA6o2kcPpg/6Qnm3oed1SaD2xExVmCbeK//JtiEaR
droS6kxydtuG6vrLhF86ta/9StFaU7fLma2QAH+IBdvPeJ6q8eJKB2lbyToxCWBt
CDql1vmiOPwlV8Dzu+E1osb2ZAEoZtOFYO4PKrTYOgJj5XYTjTmzd8zgkJg7k2dI
E+fDP3B0u96404sWHEoZmgZAYPRPbO44vu/YhrCDMb2r4l3lHn0kd/v9XgLePYUh
yOtra1A0Ikhy4YeqKM88t/uJs6jMehgmTXf3ndVGjYzo21QQKiWv8WkT6y9Zodq4
kec9RQehFusHz5/j/By4VXy7uW1386E73TiCGEefM2C5JIwIwMezBRNWztCd2/vV
65N7a7/WWhuA0ShiIjuRxhf3VQBAfkUwuA6zk42r+VKRg5CUJrXrPoxUX3VYTfRx
jml+8aKf54wmWoLoncWuHoveFvs2UvTFYdyF7N49oxE/r8IwMI50yV9uw8sfcagA
+tMVd5IDj5jRxw3p5T8IPAB2UVLXZYhdL5PbeFDd2tY5F92UrMtx4i2jVGZ7UDd6
gpWs6Mi3noNca+T75LGUZUQcKn0Hs4Zfz3hQ1BXPPqTFhAe+eo4m/XTz6pvmRUnn
V8MF0u5EYIaHZrSZtDPO5uz60ZRwgW7kXqwZtAx6e2y5ojzDfyqiTCAaWJthwODh
v6CiMwiUByplidy6k1s5BzADpxokuFZpq+CBSHbwclBJZekzj2ERcXGwd7qJUwn2
PhO9u3K0nj76cO+jRb5JqMqWbWE0I6l4Xot+IE5h5d6XXSIK3GxZFgabjrTHjKXB
4xKDlL1Gqv5LArSRDSMqVvkw6vjIrMqGDC991D1H6Z/ZHz3exhNki+U/AMbo8j7c
yQYoKXnFGWicrML0XrY+RIJgRa2YG7DOb7MulQBaeh83TODZDBEXaiJQ87+CPcSJ
p1nmpr4qWRdpgNXqH3q1jUZK+nBmrFKMCfe/Rvc8pMITNfjoP6oPPbJHTf53lX5j
wU15AP3RZFx7KkTYNJ6uyrtnzfUg1HD53UFbQeOoa/7aimyUFCLloRUHMLeCQECL
7kB3Vi3iTcaG6PrwHChN+ukhED2pdyWYR9kJswDsvFemWHhfBmZW71ewTox+ZAX4
tsz7ZkEmKCmiXy93qwhn4+v0gzMyBenICql3yL4RYwIFZF/R2NydLl5CDNcYkyZU
9cvQ3mzLJ/Uq1OVfVbZIPWFLcA4gkOFcv2x2FOZdfJn/bPI4GhEv/NKfQAdmxoiu
XBesVKSU8bWifkK5Gg6Z24eN0lP0cBBObnZWJ30nJHLnmPEDStK+WVEYHFLS4ZCY
+W483bhet+Gaz2iUv4tr6FP0bJtZxAWcUFUjEOa6jf6Evcsg3b27cO/6zJyxUh9g
Ba+WuAyaZ4XhICJBQm8Fbuw7auop+LFa14vvhSfB/z9eUFhdVsycgguK0fZ+TDYf
iuMwb4ACMl0Fmm5U/MV/fzqYkNJKv/HIqFwFuGaTYMZ8j2MWrhl4flADxrFlf0wP
alRSK2uULoorLUNOS3JyviH2VoVsTsO1RXCfjaKCjBRd74KWUnVIVh+cU8zfACBH
J8LGgx6+E0vZSmI9elLQ+TVTIJvZBweOLYENiltZU+TvJf9PxiwY7xnSR8xTXt02
B0s4ZZwt1SnlqOirjGbbup5qaSquYngIzQzGSFXofcoG4t5hZGTc8h27DI6FCz/L
Gst5wZD24uIeFqZxfjCN/h0iNArkE7O9OAm5c6wRccm2At5aEXBqzs22or0AmCkP
BrZbyJ07+a5pysQnJ/T1GsAtBcZJOu4uzgthhs3oC3qrs0Whw0R2jaybVL37pHIY
vSL47A5161pSPLHbmebYHSQ4xkcka+8kO3TsPKauzjkxW6toLaBiddaRuCbXwZOV
AOthpedLdeM9pyQ58DHs/rce4hzybhkNe0f/U+9Ii8i841nW+hv5+i2EMPIScECe
sCNleqIy+1PDHwfHGJ5fZH7fn90zFzn5W0ZrqWcHbKTv/rKmC9UW8JkPzr6b9fqw
9vujqHkf8BJ2h7CWeG19TVAk36ehI6bofgNrmBNw3ZuYWOhTZUhflr+T5qfGWE2Y
AGfzz1r8P/lHsFV9wPl8bgydNo8Kqk+8ycX0FrqaNHib2sE6I1G/5elmShecRjGd
dz+fvEwPcZa0gOwivUkNrYUstTy9zo42+ZEVt8snZAIkYf2hZIjUd46tS0zR+rQ7
zzx70iyjm4hjWubMBODwdr5ixbDLL4uJjKHHpP5LAINQqG3bV7e3SVOd6N4Lp2rR
bb9eKi0TDM7vJJH4jfDX4scp0+CxaeeAFXkb/1sWzkebbwyu41Fc1NjkkvxfXRjY
bEO6lImUB5UoroFi2oJJ0TZ7fqOEmyzi15dJPfdyraLtdapG+SZ9+AIszY94VTXD
Uomc3QR0hYxjXYEdH0tZ62aNlTBh5CujB+rbZI2iJwK9MQ1u0CsDslRz34lUd2MP
jb73UCgcHdtuHYrOVzG0XsOJrC7o4WK3gspPnvjRDD+A/kK6SaK6YVDeav408qtX
710GMGvn7SNW2Hc8joR+gIWEs5uU3bixxIRZQ2Hr3P5N/ub8kJR792t2e5ei7Eg/
cQoLvabn/eD0bWRCvh3e8WvoJxkpSRFyzIP1Bh+vEXN+x/286p1T4XqcUXozK6lt
JAhnzNjSNpFYoSqdOj9jayj2D8buhw/svs1Gykj9o5Jiz0K5fd6719F8iYQfBpUE
Cl0fnIu8xJ4xQhC4mCMK5tSrZFYennhXovFKQY7EpZuL+KemJsNWsRE2PnkOWvjy
5xouk9pjwpEEpGS/YQrNtlh5yvMF9Asp8lDE2zS0bD42jHrS7hMhS1ZMRxkvO8Vr
kOe1PDgv+ym8G5GEh5GJHWqfTGjRB9jpSirCjQ6zMj89Zy2yATfp0XLPYF1bC8F3
S9mgHk+tQ7jRYd/9wBjHywCSh1L9/ZW7ziHuCPrO508dA4kMCjS421iBcDN5txli
0+AXsBm1Yayz+9r3Bml5kUFJlSPdg8JDn9E8lZHOliRtKYbSNE+QPZLBRDxDgCUv
lu2HzzNKZK+icLoH870UjeniiPQAaPCywZL0cP7mfZRmdNn1OWAccgv31/D9Q5dE
RAPzjMjTX9clbpeNzPverxdUyAN3v4WDaeCymirHlfySRCwNxZilB/W2Imr2LI+b
9Ad4jreSEwaSzhcyb20ElgTf64Yf2teJVn9sJOHhOpPQaKthhUoqVvMU0E3a4T2B
VY/Irlvvwth01NvKYuquLjIjKmOevrLhvD89pfzD+uXK/fjif6xQiL7BI2frtFyW
DkEyLQazSAmeBnIs+d9HxuXawme8ekep5tvuqT2AuO+XCBp5VdX1Z/jeDU1rlv4M
xUpi4dhGVvtfaIOUV7s1G8IflYE0wUBwhIkeJJhwfur2cYbtcmPIcirq9mrD62fe
DDZPm+kIxIflA+YhwBI8lsQkCEpXbR6hm/N8rMZXfRtp1eKLjT1XN5NE6Kr3lhtA
YrKp3xOXb71UAhpHdE1DVJgyZXEJ40gt6A7A6p+M/qLU3OD0Dv6jakvisDtQGueZ
ns2hTGHxmxAGREHopnWMAC8q4xxMw3XjSOwF82Du67RAl9RsCYjfdVC50clNKBNZ
1oibaISmxDw3Z1OVBXr0KiNyawcGmVXImpIciU23dId5smalXu1hH8ZdRL4PvI/M
sxls+AIT+/PzKmudNuZr+rB6AWJSAqEuBhO90nV0bsmcGGGEmX3uBSkQj+NOBUAs
Zs1fcQNafALxF5Nk5J1FvNVwPK/P+ATVOTDHIyIygU7FYV7AjbiQ2sS6DzlPo1bS
b1DNo04zyP3IWfnZPzG7iUUpLUL1AW5J/k4Q6g34VzrHhqTfJqt6jRUsPu7BrHn+
5i+FHFHnfduloIB2ZtfyK6mLFkjtPPPLnkBXAGiyuOGpfPlqzybB5BuUI4yy9O6Q
DRVyvbUrhZvusc/1EJ9FQSXM1HCeCSKxsTvNI8LlYu8wl+XDcTL7LpSD3CSb7FYh
8ZiDc00C9h5VVOxxZ2U3StnNi1MJsLSQdMVvSFJ01unOjiXl321cKmjhTdGhuYSd
7CoPUQdx3P6RTXs3Z5XHFfZBg/WCO0NY95RXPusrxIh5HPkq/reAxdxxWHBVgYRz
2HEEYXu1yi3WatU0cktO1Nl/rlSgyEgTXJWwFda1fUaExFkHKciwTeonZTikZ8M7
eifvCH9QigKi44RPOvpbFIBKR8OzDRklcLZ9N5Qy2q0hq/7uI18IGpx9n000mWAm
PUxXK1Vq7KB9tpnVKv3Qb1euGmjhEw0xphmEaLFcqukwtZ3JFZAiINT+HajesyVL
q7zj7JP5epLb14TalN8lQl8yq3C9ZM625Z4Cqiw4vq04muCESD0Hn5mpks8IDOG4
6im0pTmBYeDtkH79qBGf2za/Ll14huX1fZ6k3H+k7tFSMqE/j9tROtAJmt1NvlaQ
yA+4lcN7/UV6Xol4MdJvxUCdw9vTwaT/lUBzm4i/YOn4OWDMXcsJ8zkJPucYISch
nLcoeKoER8j5DMc5UJ230h8G4NdMYVBYaN1HBAToH9Dyaf5Ov4a9hOnLdYVR4ES1
bKy5LSiLX1bjaQ0ghWYV5AwV6pz7Sgpk5ITDteyfd1qf2VzJe6vDeWGF1R9TCYhA
E6RPs2evyDjhaO7DkksgfIs8nzXDuLICqIGxwXgwQ3kmfXJRlKlvFK7PJRjpdSKf
vBXVYcPW8edb6jK5JFiZie2FD8shO6RrkUTlcP0x5OtSNuoG4D7GmdITaLyq3gqc
Fl4NUNp+irFms7px57gbbTuAuAMZYU0tdSjWzC1/PA1hjWaS+iVz8iSQoonfF4Z7
BEggbmVLWgzTqJz8FkOPBKCmz1msq2Z+LTgRVjlbYg++TNfdvnFKpff/sguYAnor
rPBNBgfdxIQGug3DV8b6HgsFckXhMuRuOxdhHG8bpARMvcIJAMdxWl4GRTvfZh6J
QQ0dzpE5YczwGV8eetR2yEDZuqt2zeID1FIGN1TPH0wKgX95pDuBVFcPKGBtkxRh
x6T4AQtmi7EYvubqaoGZbZ5PK4o7h/4qf7G7HcYGss9ErWswyTnTNcnG7c7uhsKh
GWWiMz4bUwwssdRBUHbqdEua/x6XnYu6vI4vkhGNuYrkAu1GT38aI0nHfbeaog2K
RY6kQhbmquF+2pbDdeR3QaIC06YTgUrkgm5s30yM6PHvCaurefWDfbnUSMvW8cKT
kAlinPZ9xhz/o9b4On8zYrtSaWgNLOiz7XC0r69OSZzXhjR41m8dDahlv74Fyffa
gXqAYcDzRWlCcJiEKipRN9srzK5cMcAmh4GYlAcm3LKbJ2YPEHeUUGiwduNgLBkN
UoUsRN5xMWDoXieS5eSpKAMyDrbAdABphwyrER6u8216mdFVEcAqC45xpuTTE/tG
L62awMW/UFa4jNLjbQLxOGHoGUT0XemcQaF29sTlHuUB5yUTBEUPCJF7slTn7aTm
sOYvdEKXU9xNLPh9jMLoS2esSF8IGD2E4mkn+5pFUPQiaC9WSbt8A/YoGpHF8cKi
UygQc3iqLHqEjY3QN73/A9LtL50EzsX2Q84WD/DhtLAXgZwpuHvhCDiOrPrSaFeB
mhz4yoxyZi4nji+Ql2uvG6+6p8sw/j+jru7CVG/kagQ+nn/PI6uROkIq8eCWncVW
I4sGXxidJZ6qM1vhVoezqRCYzHzq8rq0XgCK96ASpNZ+9m/KMvl/OVPQPgf/oMnW
hQHVSFW00nUkt3gofqa3dS7DuVKejLkrw4sB5BBJ+ozBi8SNJp7Sw6jSG5eOWFgQ
SSccmQEd1/fzNRktQlfZC3yP3uQf2GAQujz5dzYjiHS3X2YscRKz2gwBmepRlWuv
aCebaTno0lm2TK1WJNjUjrK92O00xkT1pFm+ff2sBWvSz7zZz/gIvdCdw9pgigHG
xocNp0n/d0EWgJPG/QScfRZoAJWoR43e6v6vEBjiwmPGXZeDC0I56m/rdARiXqTm
zqEnbTlkHDFVRsV5PS1d3VmAF0qWqfQdedFho2rVRLvi9FbvbJfjnZLrgOENbD8s
CkbE1VdeJh6Dmh4q30oARBZk0FxWswu2djN1LgArWDToJciOBMsC+raD18ByX4pe
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
NcSurOYfAw+LeC+/S0WYt31GKV3yXMEXI3YP1Ovib5XtY2g1QP9zxJK/BW9tMM8S
cUz5PQWgOD5wP2BQJwBnf9i/84K6U6SGF4X6Zl8r+216BtkUKWymIAh+sUoKMBdp
F7cGS1/bRuYFYIZ8S2465FB1Wb5M9OjkMPFoXYZhCdk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 211028    )
NVF+nDvWfu7Q+a0Dp8w8+b6lrWN5iMZ2MkyiCTtAWBV354qF1jddI4+o4Aj/rN7E
GcBLV/+YtfuJCpe/12r27hr0iy9rBEJJlImFWJu9Awys7cLxrRS/GQRDCSSKMT8R
6zxwlycPvV2Pk++t8jcJ++DIdyt+0P4xJpeP1ruPx7zIRgTTgiVcyeKU9HrGJRS3
lNAct969TfS5q8Eh46ThTeNJNEzpeKG7O+fsTkKQKWp2LDkDxGTzrD7YK7Gu6kXe
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
eyNVKrKz8N9JKSX5Fcyis7hExhQCJipphXhL6qypCThomr8kKSX0DnSyJqEUpRmH
nTm5d7XugNlBR6hka6lXVUzVFyxgSqtLkD8AbuBe4wB2CGhSDmPjCb7x416GpZkn
da6PiMhxUBhDP1K4SJMXvqmZfLGE3fqFG9vAkx0Oevo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 226746    )
Qlmi4H3780HUIK7pIzHf8duMrFEhb9QJuskPi0DrBiTIjsvB7oURloJ6uR1Q9zPP
1fckGyaP1w8zXRG+KXMrRc7iIKV6oGvAbMUU6RsM6sdEXF9y/og+IaWlkrOLel5I
iUCDO6sDhR7A7O6tY/dgN+ww/mRtWbuAiAjwUDXQc/1qUJaV35d6gRiwWQOQ7ifN
AHw7wcsFTi98GjyrVs9aypQDH8Irz3Qi4CeLYZf4VgFYyq/9wW1sWmqUnvmn+APS
ydQ64EA3zrylif0RV9GBSoFH8W06V3PmSowsbtFRhnH9+tzu9yf82n08fIcg2dm5
dmni6+9mu/QEYun48OuonDzfrVairXGqgZzBdqhNqRME/aouJSd6qEgVK13OUKUW
lofsfSlQFNw6RHSJ+9FLXnQxoPUWGOBF8iy17nbdKzLlYwaSrFe81ugEh3pRknVk
f/waYQ3oGYrirHe+svrRo2yx8eYxBvk5St5MuY8odcRszsR6ZEZa2nr9vwnLRozR
5FjelkeD2eL3C6teNFhP8RjdsoY3L8WZfnaa/M7HUhIOMARbn7pYhmnmhUB/ucNo
Hees3s8np6apfE5+P34Cmx5m6s9O5KidPh6WwjHYKz/sobnO3JFe3AO09zj4fmoV
VP2rx1CIhZdqn4mYlooEHk2XaXCt0M60lnVgTzCR4FGVS4nWOqq73egAtHaRejmQ
L6MfpvMEUmUFuJ2CC0/NAX52ZDFwqWd5lMY+/EBXdK1chgvj4Xok3O19xksWwcZC
hmDshKFz4TfG/nhz15R+jYUogELSREXYjC6yhg9LCrDJCKIydqxh2Fc9fIV1JavB
kAtZwyh7uupEYQs7BOO8OCDTz18lsk3NiwHUm9QTefAac/ATvacwt5UTgPyL1Etd
HAl/wnnX3iyx2yjsmHe9BFnRGWgBsfNX0njT3CC7d7+5aBtR/y8Btee6lZbQhLl5
l3vKcg0AowxPDIj0dADxNYIcBcWDXVfSwbERM3eU2UqE2hEDN3vnbg4T+ZVGwWfJ
KbrnzTfoVaSiJsnTMaSP72Jlm1eGaQAM645RjAcyIIIRvZR/6Ebz2EGOYc6H6uUh
clxf/Jn/ADGzhzFdPgvbU/Ip51Mo9lxxOhfiKrg7c/7C8D4rhNsNH2cwgcMMLMEg
cDWLbqftmPaZAboSFpOIz1efyCpirHrgZbNp2FQLbAEWusSSUSCO9t188nl/iivo
019nTgn18bTVpUqLASxJ8q/kz8fuuw4Jn9ToqoWjhm9MDkEgbktIwAdwpBRMGRRv
JfqoxD8HgfAqtJXDEXzRuUAGKi6XDuAIjZk4GaBKVmd5tOTQcoDEjWPROGscupv5
hc4ZOIu6A+KuNj+zrKB2Bxgux/CtSl3Vcrrfse7djDtei12NZQtZoqPQR0h3Y8SD
kJ7tV7nML22rFEGL10pjvGFQ4ZWIx9z+gAkt/xw3c6sfXuykgB9y5OMcAOHHXZNO
adG2DhMVTxOKca959JK1kFyMkEImq0vCSpbKpugCLv2pdN6KbgQYhZG6DmzcC64x
9rMTv+F3lg6o/vvRTfa+/qvF+P5oyFo3bs9GaZ0l5RFP11Vp/Z4UDfwU+qP2+FJ9
nr27ZXZrcQ8wSKrLhcum2RGAZlKjYfLIWW2w9cD4M3h3OuvjEeP6k/otnIkSsvnF
rePmHks70d8XAVqfmttymQObG65Ii2Q7fQ3OdINyk4RL5TPNEC4UOuAReYpyskGq
V2y7Ew1sKDafgvt+ppLpGpvUJqE3bqVz5gPv6LQGaUNn7ejALEeGuBCv8PJhTyYC
PzDxxdVUVLtZqv5kT9qEPvqrf3JQn2IOwx+h8wzzwN+yugAkyb6up5yjbNA7sXL5
N7Jjt4Qz/W1uskCd/+NOFNlJHgTQX0np96BhmTfDs0a6pWBPf3A9ZXCchBuPUBC/
rXOAR/2Of+Tc+idcoHV+U0xg4h1NU3ZX6e6aZThCdfxUnHUy9dod+UriJ89vRf4A
Hd6PN3pX4SMXKGz9EKWgMaa9YjkuzQPlii7tyIGIxqQ5oU1CAzj0eQS61IJpqFdI
ZWiGldlsX7Vvrj51DbaXpzhnzhzk6ctGfVKDwqmFJAVcx8+CPokezfpoqmKjDKhD
Fw7p2niCcM5mT9U0L/gjIZ3w5HjrcGwqBS2I/hlBVvKkBF1q+bEmETLdQwhjua2D
sTaNmQ2TZz4gz1E6IhIKYtqD1silPFAAIpJmwroFJIuSWjECm1wTLlUlur2bH+9I
YDAhlF2SCo1963BDyZzYOeMGC4DicpFuG1t25RdMH1PXqaNT2e17raomFd+XI/c6
1FbvNoebWKjzZTcHcmNyZa+KiEwY2R/Ullm+PykrlDnDfexHQEjGeP+V2j6yIeWo
ciEOwkk+YqjIy4MTereFXvFe6dBKmA2cWKfZQBFufWLK645UwGU9yeTCQm8zCwJq
9z2N/W/SZ7WGGo7RRny6wgcWlKUwNtTI70epdFr5b+Roxweyku/WaxxpzNoj85zo
8X1LKFFo5pkvUJgY5D5+UrJCxaXb8jLE7Ht5poZIZl/7jOb9W9ruJ6ioBD3Ik9Ur
2LS6ZzmfL77oPBpCW6WwvXUpnPQqv+aqiYODhoX4dMZKKv0c1nNzCwgFAffKhDLd
mP3Bh5yzDQ4vxv/C3F2YKKuDg5GVxoYzMHwhKSX8Q+PJXQVDKSVxn+5biyEpvzl8
bt7fihpeKSI+u0++O6DnfrQSZ0RHgfpjIcpibMXr+1EJb2tIo9InsxE1GcQMAfc+
mT5bRBl46uoGY37IbTQlgv2b9h4aV/ehguXonSMJk2gt5vkrK/MgqWxr25qkztXm
dXb9LWaQU7W73ezA4f8dDSR+VU1TPLNSwd4Z3MwsqxoGywF/Yf8N24mUmTD5c32s
7ezHKCiLjm5rjoUn3gkoHogwyzHXdpWTNVA2Xumyw1ovVGrnsWKSP9mN7wFKN0cE
ak77Cl6QdYso07MpW8xrLipnR/DZOR+uP2U+agCMgYollMA4NOrZ5fjN0OCDyBHQ
acgKHrvsTZNwIlja5lMXzfscFw3b43BMHHmaM7ux/hY4gXIvT/BVeO/hxH2895j4
53PmruYxymPoMkXQeWZltS1jUGhtCijZ7U3KLPGqnr4wAZWINjqlIULhHKLGGn07
9OfuBd7bZTqUhWNBPqMRjf6IK0oAdR6SIv+SqQ9mLvN6ya6hK3/u3n8z2CgmD+7E
RYQ8qjxUhg5fKjDH5xbgVwoNSkhYnK/B/pGoRaBPo5zbsQkBkvb7z6L8bFQUFcJM
f0SD6iZiqtRxittRHmbwLhkKv08XIgUswKNXIC+wVNGKV1H3wowhvAIsaeswDdpi
fusCl51osN0mUfDA7SEUjg9ArzWNnidMtv3W/OI1Ruh1xWlTUQqkxI2VCZut4E8n
YaOY9hdXckAFTbym2voPpwHAuOg7COcTlNw0OMXrmUoCvwGS3/l8r4cfWN46wU44
sj7Tw30YZ3HPcha9YGqEd686ANhqWrqv38/wlZJTF7tzl5HveqDvZ771ufjawrXX
isJ/zyMOlAsW+CiSFPQMWV6+p17vIWow6u11mqZ4nSsTz5V0KfZwdPSog/iQzHWX
c6SZOv31gPkOkPMC3TT2cD8GUbGVy1GLXWDn8ZjuYT6csAdCoP/ExXcS0lIaT3qD
GJ1B+gxKSFtWv1MhOP34nXXSm+A/Dtubf9hEwgwgMe7iygkuCpfPdKwu8b85tvfC
wrxdK3LmbOExkmN2AeccvFH+iseld3NqNxUKYZL9jj1hjzkT/m7Uq03gMEOkGW3M
3WlvjhcMKmrisBqjvxKmvx9gV1YDMvPq026BcAziLsfzWzjlllIVlP2yVQ+tAv4O
qlPEXJHpMBpujUH0BiIQb+lr39S2iDGImIxQYYjCG6lYgIqJYcjht0IW/avs8GFb
YDa9GAbtAZOCQPQUugR2jW16X6lInoGd1ixvPn0U5O4Od7tPUnRtLKbkbQcFpTXo
7VjWgLLvcsE3CpECEaklVqj0K8K1kUjBvscReqdITXZnVg+SmmOJr6kUf4z4kdpr
c0Q5WvIfljawXQHwBL8lcRzeC+iwBD8KsUApyKBc+NsMHPdOqpmHn2FshaMegcRD
UiJMzWwenvQRilfZ8MXxPAXd/0UBXiTyx7FL+oVvhfzOzMDdbmyXSpz1/mF8cgf9
VhH8SZdS3sQW9bkk+Jc/HND0DpjbeSpcYTPEMA9nVUFt5MOfwxPIqHwzzaa2w26Z
uy/UgVJpL1J+5HX4HmKQEzKzNPbNsZZ8CvRJ6pKdsK6cqiWWrboiX2Ds0vsTtVJb
gPfy+AVNdYH68szxtAEp8P5oRZx45cRaqg5CdZLIM7SFeW44ymJbwf5Q37La74Au
e5jn413OZrfGMJEnY4CExHJxbfaBnxrwYK39DdwJ+BmUAenZipQJET+BNMH7h/2c
r6NVTpEE3J3xE0cqvwfUXYkc0qHAeCTgCtCgmZuvapFdbwFc292x9ULMqJcoJdL0
+aebstdb4OWELahtWRwKt+a0VFI5kTObOErOp3cJkxrw43NMYT5HSjQn2ZCYj4hw
A6jeZunfegwHQ5LLkjEY5h6WC8QdmgfyPitHVa7LdRpwOEX9ffnvsou5aciu2sjK
Q1LuGQddycdhuMRU493f9D/DDp9HY6puiWWnwE0BTcKo8OE36hd+bs054lt82JzH
IR8B8yCEtN+cf0B/UOZ6S1/QGz2AMG4+0HLXdBY6qyaJ+X0d255vMkzJrkeXSiNA
fTQX3q6h2UTJV408ss1y+4xlJupoyN39awkuBK8vKzXV1+ssm1fTQaFQWGP21YcF
BL+4f9u1tBUIybvDabLQG8uFAoCWAxnyF/bu+WgUPLFUMTzT5yQ6Q55m7hkIoykU
eMPsm+yZuODwcsVzsLZpZZH6fT4209CLwITjX/YmLH0cKy7xfeljQFzLnNWJVtop
bXHX5tQIbwAsv2Uv8C+mlB3SY+uYoQRxR4kTkAbkj7UPMLYiRjv0KKDTiF5ie41c
ZZhvDKEEV4AbyEAyeD6ZCYKn6lpBUiMvt2lZf5LtGUo1IOHLToF8Ra1MI5qBmqWA
oIC8dMcrv9ej0rwLRSpO+v2YUJqm0jseGYBJ7izifsWJeAaDu5FogFKZ3GXqZKgA
l96raRNabyZguVVtmDXsMK7ohjLZa1Pvx1yD+j+55x55S+raCae6vgD4tnj5ilw6
ji6tW0802dSEE9DSCIQMcLmSNMAJuwU2WSlvGrdbjjF6Zcxxiyqk0uwhjV95Z6bZ
pnMG/Dup5ertHvflF3620bHveLGA2Rv6vfhd4y4pjHSwQqnMqVEKFOw5y+5SxrNS
mk8Sj/x8yl5DviX69O1le2BUE6P1G/mjZ9cQ0g626Ug6ZZa2zLFCLnsQ1mgIS3Ho
uni3FBQDPiqtXwBCY84uJsL2b1lDNRt6dpLCZoZg22uCCD8l/pitxUL3MMESLzz9
fVVM9xrdGFhPs4r3nq+vjQfa3P/gDJj6drqywJsb4LMknEzOIPIgCyQ1oH6h5Q93
fUd/kO32Yhu+SbZBfp4MI9qTylKB01Q8gs/KHPUnwT+50t+FOBJmv5PHxZLt96ou
cI3fzzo4Lau7fvOINOrWLnw4Shbu+kPDqhg37m2Foc0CsN2TKlP8ngxIJ3eXgopN
tfNGfpWuY+CsIkEJICf6n5kz6euYbHd4mpwE2aC0/J1Nfqij9uXyUJE6pkR89CsQ
PHvM9+XHcH+P5biJihmLYtn/Mvzg8hm2W9wv0eBpX5iA9Bz7H2lM5fWrRTk8qkgA
+8yn807saN4O79bsFRXpL1kdX09EEmPAaUVqLpvIcu2YEUPeOtEtCgqorViSmO9+
LuKYuiJjc85nQhCCMF57GIlXe+D+HraBe09xTydC4o0bmafV2iQqnBqE7SoqA7iJ
Q9/i3nZaZh6I+4YPkOTiqd3DxFABprVYtN6MfLm1rdUeLr3k65Zen80GJHP4rM4G
J3h/pOkpew21yVlxfD2QIpadcbZqOnPXkAqs5kRZ3uRoirAA2C9nvxj6IaRBtwwX
DjjyxsDB2J+7vMpmegyZDgdB5ieIlMQk2BqUOFw/be7MlVUUlagwGICs0zyqR94M
hDHUSv3On1Ym7mn24DX2Y4jeBsd2Zj2TycdrNdsKJhPlyAr3NuXYXANpyX00x5oU
/0gLDu0+FQU9hwTipYTUABeUibGoQSHUc01XS4B1yeloHQfRfgouLqAvUFJ/rZjQ
eS4tHSAAZVbbix9iXvzAwrw4oULxwcpBP9xVwpPxvQf7VgmVbHxSEucrzJZ5iYxU
+83KpIlxd5LJf2kGbc3FOmumucpWgTdxuMJhj/xLZoMBYAYww2698bKpE14AqPZ9
HOA7OC9Vp3OIckO390CFvZxrnm4n+c0zXkTqXwOoufj7WPdAYrzuzyF/dr0BeWBM
IASVrHA1Tlg/F2Bu+L6nVQEdDwIpBPjV8isJ/SJFNqqlmW9pigpjtajQ1LCb/k9x
qmO9xgG6E00fQhuNqTamIz88EqYoJbzSN1+YsJXyHRRiJMmLCqjfF7xRg3M9Cggk
mcAmD/bV7SRittfh76CRsUXKw6OCY6Vcte86ASCu9nYFaNlLL62r6Qm73105WpQk
TkwBy13rI+fAH1t3uyMy2/mjSAcgJS9l0fIzPtcqrCZ+O3LBnr1ow/4ROmZhfsvN
yXOVALRDTadQpXxZZXG2ZOlQnj8ac0JhzsciqQVjlruUFER712oyZMLveA0GIMYc
lP0gQIx95KkM+jlC9YIokgIs/lx3NOOwvqzpWbXd+ihDjkBxBJgPp5tfcwMezy1P
sLNk1UERHOoahqtuYfH+fa0srHbp1JKJpTMRXo2XKtZuMuFX7f+IOY8xmbz0aPxW
XEtfFoqGOjg4wFRRTWLSNB9o/sUPfkqXbTaz4+p73U7KK2jDHzuIO56znUDZuw7q
hul3879/VmT1n5Ir+fYB9+4/YmpApSrGr/Mgu5anvOkdIm1LpGlmMUsyz8qqFunP
LHQ176DKNA2GQCtKF1REaYBGiFFub7raP4z6LllRupNLGdDIMPelQMD4rK10njfU
8sW6cBpzkJVBPfTA35hcXOFBf55rrrTJEd85nwiLr5K5ybv3jbyJ20dJZw0KhUN3
3ENIE5typ+vAnejC8AC70Mjdwv7ZuUvpRzVI9heugZMj/bGaodH9gnZ6S/GvmT+i
tHNy/Z/sSeQHqkzSY63EFjzLx8+dJPhcxUlRAsPmpjk7QCc9kOCfCs+ZmrHuzocA
TuEs3CWqREWrYfn+k+zDk6bYG1mZQqqLzW7GcyihSO3h42Yf2EZmbcAl3qDqxJVA
OJZgiSF7RpryFR+Tnn1tcodomZS0t/hH65BtsfnXGSI7mU/k7mKW9BsJA3viDHU4
vIgH5dnDkTIBY1JdrWq73V30YoBGmVjdGdlsMz6Ugxpz2ooTPGavM+FUf2+KJ62e
Mm61vEKLWTKhlkM/JeU2hLk3jOOGcTSHspmjHz1CezmQTebDN8p9odN78KOfiKbZ
h3a59T4d8UdtDYSruaLGHl6K3jKIr01uStpusJVAjZeHsX0WiO7Y8Xoz7xN8JnwR
GrR4zFAu/rdIhib7VzUDi7Xy9IqnfZRTuihQSnrGj54VWzLzVfOri5W0akQAx4gZ
XA+fAdTzO2vWsc8QW49BmTDGiAbuCB2+2N1Gu/UnBZ8DybZ4bawXJyG2Qmdd6Iva
qimLT1l3bi7qxyJ+k+3DrrsB1meBYIZsrBB3/hg6TvpJ2obyABRINIU45nDQ9qGE
0Lih957osx9T31WU674eMRkFtF1MU+Dt4mBUPCZOjm4BExuTyihogk/HlyW45y3M
2VIHEUMj8IQ30beWvcYIdMbHFLMOMbJoIOKjSbJXKS8j8quxvJ1yRNk8jJZGbIfO
X2BIrvF+Cybpf4b5q0lnv0WgCrVeibrZ5+tTDNdKIEOArAnXeNpLAgONVXPZ6kQl
2VS52eLUH6XVu/StC6lnACEVDO13U9FOMPmfF73qJacAKxVv2IsIKslbpPC4mHJp
TsimO6C0r93Bsnx+V0BkDmfCVmC1jk4CDfOsx3vpGsKGohGlYXy9xjKtsah0vPfM
B9CHbUIIcmkmvzXDK9jd3//axhwOWoC/Eqa9nkNvslL95sgqlgYWFYqsgpkvj2cL
25t2wHh3dFSTZdmvrnke5SnS6rphpVgWHs18tobWfhsmGQWljjdWmyBOtT7m6Z6W
Awr9uRH5rW9fLWFYOEU/ecGitKxBSb1q2fUEpCo/bNb1qogqqV5Aw/kErvNDZwEm
Lkjylweh1l61+k1gCTj7A9YSLrZZ4ugZ+58AQu3FgHSSnHG/QnB0HaaL7PN5Tb2A
XQVaN0gyaaQHutwNACI3Mpfxmv0VPuR5cjv5+XMwVX/kvH8E2pBYyMOrnhzeKJPd
1evbn9I86cGigFf7Xty1XJNjas87yHPtwSdWzHswqnidteQ+fkxt/cpuh10iLBYl
a1c7D7mlcutFobrfucN2WC8DZFAFpLrCbNeb6xyFKdBmN0qosgULRunkUvjljDCf
3wm4htSghyjJJX78FSuz7kWcApHl459G0N92UyCay/vQnP2b7CX+On5IuHf8brGR
w5xqeuf43zvOhu2mDQmqrb5FIOSnFsWk/lr+uFLFKxkOcF9VCfos1DbslH8zd6c6
E2vN4SJF+UQy2a/PdfRm/Mi+6OGMOKU3uSeAVVHcgfpysv1YNO7g+3JcmuvCLOhs
fy9gFY+kDisoPOR8VFZ8njByMA0t5owzfSfVSNSKsciblSbiuj9wIfZnZ8GSf+NR
YBkOABmkAfepepEewT0fRVOGlXfUqSDodyT+32FLXjNI2o4vSnsiuXBfWpHCda1A
ByQ3dad2PeVpF/BZ4az7pH7n40I+eG2rNi3BYr3lOk4LrSM7OkHPlySmaJnjKHT2
eqwWxSgPbF+N914iAMPctcUCqfley+TBkHwZdhYhJc3MgcXBm0X83VxEYpjlqbsZ
Z4Cr1g/rg5KqFf8Nq3ipBf2JRt3PRarwJFT09q6f/I/p5r8Xjc9CvJEP8w0UA4y9
5ZYB29oOS6HPGpc9aB7zJSuxUrQJGbsjUqJemoHX3XnVjE1I8bO4rN7AZ7cvpdgA
FUeKNgLS4Zdi0jupmwVkmKjgb8VYpWx7m5+gJ3f0b/jAN9PDhLq0UDOIjmGjpOCE
gg76U3Hr6VCXqDxqHbgwNyyJL+8bkwHy4uO24eN6eDrlLHIlkc4Fg9SZZSID1UMx
Ehpmef8sZKm4HHynNKBwpe01x/YANZ6OifK1PT+7qCpy0zBGiBieT1TslMp5Yq+/
kfn/GOTCi912nxk6G+DSbm7PiXX5crkhMPaCCQxEm7Xs0JEDPXu4pSsT6AaSq/u9
IT3Z0+mvLmQDc3vCbOAOElXcoodczT0u4b3zoN4DMUdx6zio/WSWZqBN8EN+bzL5
UCMJtIYohHE3v7o03klr4fA/K0Z/Q9v0b+ZVygamQBWOsBHrj8PStOKVFYGozGt/
w7Klrd+/mXKJTjSDpH6cDz34H+1Xas0Rq3ihNg/IPEyS5H/rz2lnJqsXj79y8hdN
ODS6VoFwnTbAMvaoL9LdtvpFzWqGyM15cDSjszJSheEsUa1ic5abOV60FzvzLpuP
+fIuetiuKD6vrmK2jFKMt1qlrq//lFbBaFTpk/tpr8DSWkLKC3QCIDIE2Ff/pcm9
On47v76lVDLZl2gumqGuTgh3/QPzOhr7T/3SvCSMxrPrgknacO1Pc1HopYzBRb6p
AVP4C3Wp2uZ7y47QZHLMArMd0zPzf96sW7vC1W0LqApr/9hkL6ZAI/CQzCgyH4Ag
vWNH23sGcrwPlEu+r6VhVTTZuanHv0IKZnArssDfsHV8srTwdeGf3r1UcTPxhWzz
1EMKh69j/DQeeZ25/DKA8bmtvYtnVUxZHiJ7lnEgifrEeRTbi1s70HuygNxHq1lU
AkoDgVbAcy+HIc3JtlMj2+Q8DETFh7UcHeCpq5PePFmyl+pdVZE1j+96AM7Y6/XO
rE4JaiMXW29c9UhKVSQjjTNjOW071cMvDSum/CUvxNNbddpuhF0HarttDkwT+LdE
j87BWThZiSJrkahJbVBEpQ5sOPzdNFsDZzClnGhqiGQj7/5F7SlqAmwFBx5F70RW
RMRzk/28iEU+Eu3ubiFHA4rz0Cxnod3rL6ZwW9NWSP9zB10JG1oVfMYQHeEUP02g
ysFPjX5Oe9Fkd+CmkafQvjqWICJEf1jt99E7R6E4DprQ5gQ6wxRMmAioKM2RoD8r
Oq5kBpkbWT0dvDKi5T6DxCeHs/4BbR1/IqKnBHAfRnztFv7ENq8dEAP13Mgfitbx
UVL045aw7e6/XjcwqAMio0EJ6TDI2cFwiWGaJeQDxrh+DJ5n3zNFlwVEDu3QCLQI
zOixM7dg0jw3mRkk3Fsd1cSKr3qATg50cEOZXpJMJ1avtfJdSSuKa72FJUAwx0Vz
KWytaAZ6+qZT2sjx1h2sNYp9plzsRRHIc4ws/Vj1m6b7FwS27yTFyY6jxl8KIX6X
P4HlJj5a3Hrrr3cSAj84cNUd8PstnkHz0PPHCtYjz+BnEJLX0+Uoe2NDYjCmiWCx
HhKP0tbVzGbd0+hpU0uObj5TAoJYv6mig0U2wCgYZs1HC9oKqEI1gQzrJIu8VRX4
/8Y0UQrFh6UncDrzJKgdFl8N++4Rb41SSt8r4TvJ0NPtLGdh8tEcr3aCrUxHlhS6
KyuCOiK4Ytx64GEF9THeaXZC1ELbbAXnGS9XHIceb+VNcMn2xz/GMfLbxwdPXH8O
/d/yNNDkZH5inE14zTMeX1N3fEg8ZdHXK6tCwDEan9ceQtG81f85jRDJFuCH7uYF
i7nTER3lZkZEoNzxAnkDYWCc4Q0HfmXIwDAKNiN4NtZD54515s3fg8HR55HeOZGB
oB++upxCp5OV6W8BsgdIgicZwT+657OXyBQMGRKTVdFOZQlZBWK7Ly4uYebvVNkZ
+o/SyjSoBhDgteE/KwmL9da6bBWlcEareGbb8fVRsclXXfBeDdgi+36CRqb0fduD
1lxmdEBF1sE/p13Q10yWB2c/KYSLGnAs8K9pGL9U/RasqlVi0QN1jyvPtPBwja2O
mh6poke7DvCTR6pcJW3ROdBgX5lZ3swqc0EkvsVUoUrM5m4MCGCltzMyFqHAPwtb
yl3OOq0Nh+HRBW5a2y57rMgMILqOEeA94z0t6yXysmVtn7ASC38g1hjcA95Zt9qU
HuF+9DJdmNrm9UT7yxlReHuKDjRws/vQk+3hMK8rPQURKsXJAOT50Nt9iUq0imag
GlaH267u0Pd1h53BoK5pmVLSDBL33W+QZWxpXqaWo9eP6CuRcq/0qZav34Pu1sqJ
a4s+b1mVBlkLgcZkA0rBPlvpLpEDlnq29wKDVvN/gQ5+++oH7kdMQUJak4yy3+Ez
YLJk697uWgf/1q96ehCNGdFDbTfOFInS77JaklT0Hmd/SdSxwoTDB1m0AR45pnKD
MqE7uzg89HOinGjFutAJK++QnjyghvSK0jbYmNM3/uA0XXZmXyKsq2iMSxjthyH2
K+xBs3QG06SZxuiG96s/9vesJDjdrJRJAPi7GgV+MPEUZtEZweJMtSLlDrc7nvDC
x2IOlxb6CQmNqXcVG9GbCv8HP0SSGq1v+3nAduaET8oyIK0oOiurWgIjY6j8Ujnx
GQpNlZtGks/B+jq2WgrJXOAWgYJ/PccSPNo6kFgmu3CpKnXPJ34fSqhTtMUZklOe
AkCsF677V+Vb7SvYCw5ShHwHLBJY7avHUrpGqjI8wlZbP8Rlz0HHmfzjte0dx7ew
2q2N9ZDtHzdzNsjMJG214rXio753g623SYCa3t7xUZSC5+1q1umT1WTlHezYVkh3
rJi+0yUjOmiEN71c+E2nM/EdbbU82CNTM7jhAdAOzPinjIbvQa3UUfiiFUz5Viw5
O1J5hdX0pL6nRDGh7r8xzCjqhTu05cPVul13hgLbencixUSzMH3d4XxAnTzAsUGd
ub55Qe9uGRhgogsD+PBqJf9lBjMHUxG5utyegtwxg3uQ0KwIQQFdOSC+7xGDuyZV
13hLmjKhWTR7twd1Go0WnSDa1t45UCnNvBGMDnBwhZkbqSM3ZqMw8NO0uxEPExMS
4nFBQv12gEjyJn+8RUhUkphHPudOvx5XmZSxmOD9ZVwYrKOTtbKEVt6aOi9zTWUa
aRjE7fiEkYXNx/kLFTTBRM+CDmhUavH46fZKnlEq81DS+oJvMPl07d4OXvgAD99F
sJQDqcEfSxNn6Xm8mmVs9IATk4sN5/nX8XmOFiEAX4QfBLqvcAwTJmpvRYTl9wPs
rKgtolvbeTEIPl+rPplmWNTZ8wa+dOPTR8FEhVYUBo9lwxiULzpobipRGCcFSn7d
tEW1Ejj0xt0GeP0uF+Km2YNygmqPZz5+06C1h+hRaKWi0szuQA3+SBolO0BHiD3r
UasdVjr85wr6SfP+YHYwhBBGp1tc1Ay3gOka42xmuZlbebckEkglmKHXv87h0k4V
NVoFVhqGsNFwwur5re2GzWpxYJDFGmHWIaXAN8gq5jiCxC+Cl+9IXJ0ZI4T6I/nt
66wXu+Yl3UTfaybpPsdflPg9hLGaQJSFGEuKDcK5q6o8MYzagxM39ntogTHydNDV
hvUiKFZ6F2cFm4Fwr6kI36al+SRNNxbTRLfxPK7o+LnlzMd/VB9quVrrk3NUZCgm
otfRZMqZcmVNTuuXt9shGJk4m8Xb2RjHvdvLDDKSABY3bG02aB8lCDPbKjLlOIOc
1nj41riuzIDCG2ICpQKc83jC/4yaQPxuwlojZUdXyxnBRXzydSD+IVEbunjFYPKc
R1bIICCEYeITbddQhYyv+dwCkoJQRNTs+PL/xMaIc2ts4x/X582JmSFFl/YMckIk
prBAdOkTNPIIjz/XHtJGuJFONCWczg8WHj4M8n5TbN8RJJn0JWq0zL05iaueLH/t
3s+ZCrtxXICq5x9pBforvF4o3JyEgb3bdY7D2i6HIst9B/JTjfdEVJfi1WZ5i3VR
qSYAJ8bv5LX0bqQRm+aJ1D3/8SskGpEduT9V2O34mppcl/+rzsw4zDE/0yvb84FI
nM0Oy40ga6wsMNPKBMmBEq2+8J7pyG+YOs3rcga4j77dqUPSQgfsVkYm2tNG/klF
hV+dM0QHu6aG1+d9u3JMzudSfTzL1Vb7kitNTyRVjAsqT0clGT7E2yRpHCPlhDHn
34ajK5MvQ/zM+hbr9h4LmnMmyNpkES/SVpa87put4lzIVyPtmp61PUQbIUiiQfHO
KsYDQ3Nr33DwCXr0yv6vO0e2GbQfP54v1Lnc4GhDAJURZjUrZ/tumHS0mAILexg4
tYTCMuawk2PBvuNRrZ2DR2XQbo6QkeAgxeGKOTWPlKPgG9JPxVQOi0EjNYZg1D1p
Ifrv2X0HwGjWvcx6TnyRVZviwADsvs6LokRc0g4qFsPaHhJ2HUDUjPiaQicF3uYp
EZHSL2PAb26GrPBEx8TMc/iXr2OkJt8NTY+Rd8+BEl7riKuL2RVCiC35VLaknbn7
v5uInBG5+g9ibEM2w0lOzCBukwpR6fEIFRmQIThPoXYXti7W1BB31LYUfp4mNTRW
j86mn2l5H8Dp7q/lisQO9hYxr67acAQcSfiGUTHsuHbHVnuSTmJvhUIHJwi9e6Iw
O+LLWf8RDO873plpVkrKL+dyY/uQSkvQmoB/+UOo9kyhDg843qZW/zcIMYapJ/kS
OqhdPoTsv12UB9yN19V2pJyPqvzWt5Orrq6Wyz0vTTshN1dh8lEw7NkqyzzUfPIc
cdjJqJePeFPjV4UOPBmBvSsOJEqg48X44e5Bm8Bole6vCdgJi7AO6ET0rKWUs0Uc
3VsAYHynawgXO/IJVix9y/eAI2kuexdVjRUMF8S93M/zdnarFEL8Y/wpmAzhvLue
7+13Mm/GFFSpXn71OgeKAl4CkuHwQQ80EEft22IZ7sMK3P3aHh2Oj2oURCoPM+Fe
OcR2ZrrmxSk2NUbFat+vzKeSrGZZ3vP6gqr9qZ8dLPZwns7ujlaYb0G4DHr8efVu
1awNdisBoRGt+ZykJG6BFZOlH6r8Jvge2CsngtVEOChNOMBSKIthNUAFA3KdM6Lj
dAWSRr9RHvoohroryTi/yDUZZAkVMnvudLMj7ndiae6maSoD02mIHlPVyxPwwU5g
c9U9DCjBNg2rXa/QrV95uURcxf6Wbuj9nTbsSDJG4A9e3yKUdHu/OJkas6gps0t8
r6e6uqnaLu0TnH5cTHloHyQNwGW8Wdlz69GDmjsglSi5E6OhDh0DnXNQow9gUPGy
jFbzsaZyxIaF0CXALSVPjkyerdaQZxmTQgIa77pcZ4uEWhT6bBa0KexFt31U5kCo
3DiUSKRahY0wvBGFaRxVNvcZQAayVjAn9F2Oy0Cd7AJCn1ICT+r7xtejslVF+fK2
cQpFgfytHk3OR0JkxjCwMgA1hAhKYvUj5XxrxkJXLBar1komh+qKLGpgXl2YG7f5
DO7cvxvEzjPLPmDkoXLqexc3iST+biJOOfPpQy+SlMh2GIjpN5nT3CnNWUZ01REI
7jOk8HrRKL5SVcFooJNRn/iCQIRXq55vG29jgBmsPU12OZlD+nxtve8uAeJEAudk
omqagNZtGA46+lj7UEWJ6ygMZozxxRWn/SVcK+lXzk/Ck9zQri/KQ3WZ9tZPsNWx
iLmUpNrOhfuoMu1xLbxzYGnnml7r0UjMk8LRlJw9YU1OOeitQPrponUaNZYmRQm3
fst7k+D+vVz966PJJ12Hpf7A6Qnqy+D+3n+llXobAm+BYeluyc7EeW+nyQKryNqm
oxQOtwXR/z2HbQzPaBchp6jm6LFAY/sfndchTSFaQ9yjdch0y7k0m8HZ0weprI89
+1cLLSuTRwEwaSvM/Je3fqsYv4GDXHyAhi6wz1r2B7hqLGFxVMO+AuiN+uMx9gkt
FPtVYlca5fdxtiCWYWCaKP3SpImh3jWbbtJy7w330zDZ7gX+BxpCb5MqgQ5N0Lwl
UbuNjK3SOjhMC+nAGpOaAwiK6cjNvldxGFMtP7ub7kVG7ald2oM5BXAOaFHIPij5
TrDlm1Y/CKKXtKIKSvaUxlMQCJ06opbYEieWZtgs1ER3gr3bugVbmew6Y8KbEVtv
ea7kngru3LNtP3JXHDaIs0ukwiPxSoxLpYCBTdMwLZEuYqk9fl8oChuaFOuwg+66
5XDjN4OvkzvlP35A++tRW5yA+DX5dF+TW+pV2yobk00imOnt2/FI32Khh491BcJC
TKeKBvqepml+iVQvMlA6KPoxkgd3I7X0BiWwctriad2aCce4bLJT2iFdJKwTUDUj
/Vq6fbpOWHQto4Zw84wzqA2HGEGfS9kPZPzbN/5HTXrOD5fOpk0qs5w3Z8s7CPda
OMXqzWF6rpLhv+JMkdN2X00rbUZBOqzSI5KswvmIVMkYprmnuaZq4UYrmipDs3j7
8PPMxj/SDC68ampp6K9KgL8wDiEhATV5hehLvcJyN12fDhNWN3XcPZpLgNGmWxDN
5lsrPvG32mT6t+JC9QobgEzUEy0kgRUeskU9tw27nuaTbfj367JjytN4yZ0J4KgI
unpIXzKbdlVGU+AXOntGVWszUlWxPYVmp/5Vg/D/a2okxF081jjZjRaP54UU/3g4
sSaixZFnnKUK3SWLAjIvJ4cqMXKTWdy29idqIAZGTmBS9+xhSoMVg4Na+ydrZWAH
/EEADWc1UXGYaxS7GM5x78+YgySiG5x3s4haIFzbvz9NZzRVpOSuqSDhHn4gLWI9
fOWAi+8a4H0fnRf44dFS3cc2h2OZMbSC6mVobtpXYYUNYr+DEUPgu3G7MtMgG0h3
uO3/VErCkOgKFRFGdBq8Wl0WmoskHyMsAMSIGBBmNU6pPuhfQ+TCRijasGMBv4nz
44ttcDB7oG9bnqvvVGjxclgILU4mD0vtHKalTjH9XHHSa3s/uoES0bkfH0XiHZ1g
Y16ekRO2/zfyA2nTyNyFJCX8lHGoKxgG0x66wdWbSdRbkbwnKj6bNt3aWHBo0pDJ
abqcUMQPZOAhu/EbiUSLmDN/1RlzdBKf72ZZEqFb2nVzmtovaHZzKYzlAYge2fgo
QeSjgoND9CQxgsHGJ99SNbxULxIDnRyguZFVDDVFYfVMyqu0vc7XcV+3NGh0Isgo
LiyhE1hTVaL8NPiPdkpPYWHg8ykLnpXSlIR9zeji+zO8CUV708sGTojvzsWktn1D
GLb+IxjQ5TBjSQSLaABztd0WMXlBWloARvgzj6ljeaRXCN855oRhwgiPDUMQekQw
GvVqpwiwN1ZvIUHPWxxDyqSLp2hrK3xNPdxjrp5terQDNFH6gbmKbWdjCX+mC67f
kUP16AWxzMs2lYKHmO3XL2/QbiQhkFGOy22QlgM69m+8r52gSxZRnCSAy8rnIMDz
7soUhmCuThc2G8D21ujyNxCDmi9zchH1pIalc4d5oQyiUlCi5DQ6WrUUyweRmtDY
pZb544/VANkrV2o31H/IslkZNq9unyf4xtWZZ2UgrGTbxqMAbHtMB5d5gST0ZlW7
qS3E4qsj7yDThpAM5RkSHbs84FdzfYrfch/EkLk0zR5eEAtoaEH80pEaySbnZABT
d8jmpLAKdW2OiG/GDWSVpwOHV3W9cJgZtWa3kPa2l8nmRmUlh/zoKUXCya2Irzlo
7DNBRkgH9m5XD57RS5Uw+IkMDG2XeSj+wzizyLWWQJ+FZyncK7UypqUqJLUksKpD
tsGXYr3RVOad0aN0Sap95m652v0Fj3fomUxeJy+XQkdFTLwZxLJw6zcipILtRQss
OIbtvuhZ9DDzRQ6GpgB5VTct351GCJ9Z5ORbZJKqWmUuRyRTnZcoBaT1aCMgcjBP
cZC9VUsW1kaa8kd6Py4Fd3f7Wv4I9RXz4xagToUSUlHeZtol61yxIvYgiOIzDi8A
mZoRnFg5CWCp0qW1GaTHNHKrUowajVRicFq86OWkCYEIiCWjcI9RC3oCzhDH72EC
AdbfD18YQg1JL8doVBUAcue30gqnN5BAdR3bMy1Q2twty6fvyyLXAxNPLtTx9JCb
aKot3TVEm2CgiE/3hUfyenBY6riI1kpD3A3UvPf8QfmwrqPQgSN2P1pJrfNvB4T1
yE3BzvdkdEcLgJTt0ZkjAzAK8KeHH/tu+YoTv8451M81NIDoaHBVEFdPLCZyGJj6
h5znlKGZIj5IMDlOyzVF2G25DOLz1AVFUfrpPwKcfG61I3w2R3lIujjo3j5EdVoU
8+JvPjHWAD4S7GGgSoyBzVH1jMuu/GQGcpJY2uKsNtwijSLni5lTWaxF/MGgAPTP
ipeKO4IjcBtmvJbmRR/KQSZX6NkI+jeZBuE3nERDaMKZtb3CuVK77xMomPFqgNYN
yXy7yEBE7F2OJt1d7wfsNxSkrugeTtphPmmY7dknwqgWr5Flk/2Zp3O0+ko59AKo
zfjm7w8iXyadz7uIIbS6IuSZ6JALfa8DPexaeMP+MANGEdnk4dIN0XskuXRAHzOd
nEcx/qYQqQ1vEEg+WwnDmW+tiePXyF4QWBXZ3Vsz8vCpJpU1t+njaINDRMlkDsrR
HLLpEleAd0Yp80CVbRySuhIan7EuXfq5ktf0iha6Na8+vQsYRooQYClPGsykaPSl
qs015MiXWRznrZ18iyaHfL0cHm6DflmP0N0hz6BoiADz+IU4p9vTu7iN1mBFcaes
vERS5WI/JGzZNZ8KGTYVqkHPeHuw+N0rUJyTbFJ6UlHUUacArNyYChH2hAbL/oGd
W3H5NUv4qIfUoXLbpRSkvEpyrPhHIOzoyfLmDg/XbLX/Kd/AUzfhRwE+jMZ9c0ur
QskmCoDMhj66/MkRmo0PjoO/L+KH5x9BgizFRszooaKUkyv+kJwH+3XqkS/gI4ob
fFGa1Gf/nk7Xu+rYeryJCnotlOBRzbL4plx8Wu1Mq2izL6B1OukGgfp6d9TiMbuH
7pZhuPgy02q3Q7XqhTLQnv1gu2YU02oQ1PZqzbE17hinangOUgLiuXh9WrLfTOtc
/6+YDPnA72tsJVH841QD5LJwZBJ8r65k6/qPmub2hroTAmShMUEQbii5JuCNb1ON
75EwvdWXhhiotMtyOLwGPBPqbzQd+Fwslvg9rhckw9+CZPk3P43oFVBEgNHHtpkD
Vs2jWkOr5rUfxnQZm8VWx2D27Xt693nQ/SJj9WN549lyas/ozVmOQ3y6Ys1AJpUr
XxntgkMlKNRUykjwxqkoJvwHOnPvNXq82iN/v2EDRQHB//x32WhG917Lpx/rt4O6
puKvDeUhyBK8VC+tiSu6Hz223WlvtfaaZYNtXm+uPGvj1wjqPc/c6TIkiAMX1zme
M/5GU+0gvB7+cEP/9vvxQGM5utUyIUs4Vb4niP/PTALc1Vhla4OSyod6Kn7I0hYC
DuLeqL9f5qk8jDiOZiuVUWVboHjt/hUhz9JLmVuEp4769rXnWUbEdq1b+ZD5iFer
rd56re+ezmWIrTvzOPQyqKKeDczcnfEXt0+gSPn0sK4cSh/+ug7mo6MjXh7oeXGn
TGboDTFDXDBS2SyhjFaAj1rRs0FkQXbXbKCvaFXJkhYakR1JugYWA11yJgSpEIMD
1ew6JfKn3YMkZkIv/yJ9nyryOjIEHXzO4/GKI/l8DACOKl56eKwHHq617kKx0I3q
IR3ojbEba/w++m4GPKcRoyKMVsmrDTUQ9ho9bJMCRO04Qyt/2oZrryRIk1C1i+sx
R4S6mAvWGagr0WR14Ym/ZxkXOauMm++COS51fgRN0DvfgJYI/HMlucR5LTHzAPCd
zr5WsRRV1XrEjtBmBNsNCRNNIwqceNa249eS+STg273Wh1u2CTroEzidBNWNhy1G
x5CvPw2cL5J/zUciWwrGTKZtMik+nmd/fGWFCYAvIvlMK0KZAEuvILW1hPNB2Jtt
MFU9f7WhjwYAoDlHuF3qZzkjeJrScn62E0nE55g7i6Zrrb7AV++WbIh8dVBOKvMx
xgmqFxzkz05jpRQ6Ya6WCO9ByPY5khssSHFXkciSG+rfbzk9JBm8AID83RygPq7K
fPgsI3LZ9sFnoQfwsd+jpAAjxHMA+mtgb3YKZOonjqeohBXID8OP5pUecj53lUBl
9cma2ixxw+uVt6JYKPkAwaL9eu7fBu8yvqWBJE65F6v95XjiMkQdUtllI6ZXN/+6
XRm6uuoUKasob7P8C/gCnDXUYn7Q+9egTCFbCYSklIEfivk3MU8DxD5WQx7dbjZP
41cUIlOGw8eyVBKwNXzwjP/Pd3e5qRZfp8Jsz0iU7u7+ZrNUrfHMKSb2ter95kWi
eZ4uafWQBtp7nKG7vM/u1THPvcplAlp1p4rf5yFr7SGLXy6CQG7CuwBqTVK9RK7T
rS+SEnAcbLPHY7/+DZwLhxPGXVdpIVpBR3l05pLEMvzTqx3Z0GbbmWnb9+9FfL8H
Od7QAnt9x9vDPY5UfqHtqAo/oFx2NSRM3g5Lxp2TVwAMMguYuFYfJ4UPa2LNIy7w
eh95tik04+SBPk+KgAy9cdfXldy3QllNxKbf/aPeiHhMpkIs3N2DrlGLPMqQ27pW
L/0Q1WLDpnAIEMsowW9MZ/6znPQebmwTGW27aSLoecxfHVUXVA6zQ/uj6+emhOoA
IynQjigeepzl/w3XjKUAHnC+zZlcvRjSDMARc6d8AToVAX5MlIFRd8J6eCZqRW4P
ZzIZcEMb3ASsMwzQM5kIae6nlaXj2geM9zVfzYMVKrdCTpS+btZbtV1mIZjQVW4Y
YEpDjaO/9DIXReornEOWNuhV+KIX75xMi80kZHWlqnrhAzeVtryLFXBNNONTox+q
Zr+xYCADnmSRVypd3P4RGaCy0aZfpmzaldofjXuhRBjgoXPVv6wlLu0cSxyIZyn2
7qn3FzCS+k3/aWHraJfxWd9SPCcUohKpbQ0vu//VtqdN7QspXEwlDVd50IuqgvSC
gMkNf1fi3O2dvpUBRX6LzuVdil+kTR4mJTx+Bbp6Zcwk3F/dYrI0QPFDmOOOo3io
qE81zsFdXMdHaAE0riSe3Y5mnW7prNtxDWUMbhS6uC4HaXwtG/4hCX8qo1cHxi55
akR2D0MHWw2f0a+jNZH9PQLNZsWygauMX8bZQE+o9VqaByK3eqcjBF73rsQHqMK3
/1m6+SeTVS1xUQOkLLWMa9O5eDhdJuxcmDNkFuFsM2JQF0E/8GtvSflXtweMkOTi
za5nE4UVaFVX/4SiW1m/2XJjruflyARBjQeEozDg51LQpGnu7yGJ9yJnOY3Sr8wb
g1vT7i0IF/9woxn/VoLMnFeq+Fa5l/o2PAOQh73kRKZT3YX6KBqLI17JyV3/T/vn
mf78kltwLZorMVsGJOPPY5qXT48zpYReDgK06mK4QvDJsKjsUwbnbcHwZSFi/nFl
FvFPtPAn1HtCwhnww1i387+XMLODhX3EbiUXpSnX3ZItqBzRg9XtaJeCLkUbctXq
kKAcS4YAL+YcaTnczRg0pwtPhvOnpTc8ozpFn9ydwja0/0SA/e3i0+bJ/JguHCUD
M39C5NxN11y063p9L2SphDasebS+5MQehha+oSgDpVHpdXSpRoI+i9wHQDesUozk
2vJdMleSZ2+TTgLFMoLOK6lkZRK2gqM6Eg/uuXDJQVGpGQcfUJMwQvC8rlHlHLQj
wRrTwgjUef92gH0bJ9ToE1tcI8T2/dt9plJiKN3s0ZPBnlWuYMDGVpnk3GPNcSnE
hVukHvxBGmZd/rDmE9uHo07pyeVUbk1nvtPApl+6X68gewRXNuDin09AwhEjSdL+
0elLELAIdlgSc4e3vAw8SwTbjNJW4CD+24w33WS3jqTM9n8BgJG6z+GgCPlcjY10
NkMi7XMxWli8De6U/aSEDETSQUZMw9BQHx0N2H0TwvHYVeK4wax4eNRevy/K75SW
opFNYqjSZzM2TptqoZn/ZexrbP0pf6sSqix9VWDA0YHT5+qzE5+2W70H6MRY90jD
8EXlzKA71izczgqPg9iXOPB8NDnLFtA0Cf+87V6zbiM=
`pragma protect end_protected          
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Y3K/BzUWjM6db9TE0vPN3+w4z+EZzT+pvUTSSN9iWkZ9h6YXSeNZ7zA272XVis7A
SZJxomWkoUSBnUp4X3lqy39OFCrA4n+nPGM9DHlUcI5U1wP9PzlHOxxwrSdNET6B
0TqgNr83jNZgu7v3Gv0/qPX81h6YTa8xzRuhpCIlYSs=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 227205    )
rmyR60NlboTMFqtqmnJ/l+L9HIw1YBQy+VCYCDg72N8/gPFux8hvOwLoTK6X9D9V
hg91f6Ce+WRYlZOtFVRGW2FZQgb57w1iBy6y73uGjN6rGf1Jrssaw5508pBSPlnW
76PN2C6ponFtzqTqDFWQfKeHlV4gujb7oAJ7gNn0b+yxU1Mb+Tx1bs4F/WVYNY/2
XHIqSfPJY60ucBUduKn24oWT4m5dW58o3CLcjAYSMbJWULT3zTtnEIpdTQFiM2BM
uaU+q43yenBx0kNErrbZ14rHMZCGQPGTiswArr2506kHb043cXF9g6ymHAs+/gNb
J9Do2Ph/9ZynJxqb0YAGmdRZjrxX+fVZLes2u3mPDoUrBqpEerQ7iKCwjq6I0W8Z
IWJcwDG8tj5YoaxyhnyusOqDqEtVKjr9Du366zEKXyquE6wCvTFqAzv+tQ97WK/T
TDCeOzEvTzUxY543EwQMAI7RebXOebMdeZyl0EYgK2i+FbPbRElWt/+YnACrB3WS
qaMdh/44XLDk8sf8HeFBiJk6/5WUIeKw4JEG1Z7LF2F9vs4tcCoDnCyDSui/uKWE
LVkbzpIBMjl15EhZGXnGFJ2ZW3afFLmNnTUalU4/S5g=
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
oe0jCnlxn/05AJMcASOBlemu98PT0HwxayZGh/16MlUY+Q6yvjBf7T1vBS8+ud00
+kJ2sGC+y9JmN7lNMFeDi/EqAjbMwjiEYJ2ePv12w0VgSjGwnN+0f1GUMeHPmEuI
pQ4WQ05xZ25E2arySHF444+Is/OnpXADM/7jYTpcryg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 235349    )
gcQgyX1i8rAZ4LWoaGVdVFw+59BqHxVCbJ0BCdRbRLjz0332LoDIXW85rO2h1oB/
0p6O0QNjEioYAFhVOAjJ61+agqYTTsQOsJbK+Ghl6XXwV/9Arpdw8TQ7Pk6Nmr5F
n8b66EXu+1hfBKnyrWX5MvtRwYPouoXimZf6sIZ5Dc+8tU4zJnLpHkg+oE4yX4Q+
QXtblJ/S20PoeV6niEjXBtSiqt8YrAmQTOX3UL2PwFGvo0ZBcsjQwKYDaRgvr/i6
zm3nIZn0RoYfnp2ogMGihiIASex0zdcH5OfrgwWctMC2PdYKI7xu6DuG1I+CMpAv
fRNh7aqrKmyJIL0D/JXMsEd+ePdppjS3R7bp6Q+Fk6bicrJelv7okOAImFwcSFgW
q68Sqmgw+U61oxUOLwO24iIuBaCGx9u2+BFwZEIldOMrJd0vJaxmN+m4AWKU6UcI
voJ1N68P9Q5tmjg8CQA6JmHv7xwrX88Z+dggP8oUDISvGnXqW0A7nnHTe83EuD/6
h8pJio8oBRE7lr2korrHYLunX/JVH5QumWcJetjEjJofHQXIFDqx4VLRoql6q7Vs
tf5b34p2X1Wubmhk5v87P7xV2eNmXsMEZEpZqUbUFsP6TeOtdgMrtHip76q8Jb/O
cZbUPGk8eqi24VN//mfH2RYstcaLWGLHgRVp8QCKxfSaNZtCMYiNrdt8kJyWsxQo
qZIcIkdEY/Ar3o310C/Fww4ZkKXSZRekooIQP9ahZLEcCNDoXrgb3vYTCr/ahuJh
amVr/9Lh1JypsfyU7GO4i/JD01TF1u/WNEocwvLUb0FUnLqpVTAlRh9h2gFj6K0l
88Vm7O3g+Ed/E02shWBdMA34UJl2Hx0tA5zbxv2pvOMAqGZYRQlEk+mRjA4v6mPP
0memblZtTUa3ZVA6AaYxRl/qmP35Eg9PrWn/0QI0q50Vg+qGHBg1WWJ/2u+LQ3WI
3uLOwEYBQlhGKmV3eTE0ny1q5ZbJdXLLaJyYFNnmrmK5i1K5lM6v8eX9PynsDF7J
5ZdbQ7fmzbmVNGgwdLlJKolpV9g4/u/du2CDhBKD4PRl+/yhHvI873ndJc7YX6dF
wCzXhvPGxqWjGgSqLFJvO31pwHpZHlVH8OZ9YQQviNKPZaR8RGemht83QM1TsN6r
JRtMa9UOvYbgaJRH/SewAz1C1oLzSDsna1L7tB4/lX8CAFOohXOLysYvovh+fbqU
7zRhyATavxg5hm53VwQ14EBXXWQwhbbS4FTX6SQAWiMNZ8uXHAn/R+YH1M1kQqUp
ANdWDO71rE8TE/vrB/X0rM2IslO2p/3+1VNnIUY3sPfe/o+iUnXozpJBAnTLuady
1y87T3PX2gbVcckkAWcsbhRPuS67S07wa8R1qSHJwHcmgxkpWIKuIfcouh5hNSbO
zrPkFPC6oVINOmypL0m76jX8mIoaZoOomFjPpW60E75/06jlRgfoHl5974KK6a6o
3AghCsFgynfwhWBCu/J7gn9l09M97YzC+zyFbC2iMPnhu25EuYXV4vTC0KoSH3dT
YMXK5tihzxmoF/5vRJOgoyG+KNf/23c26DxBvOzNqiGknswXbLLvcyU7hfMjsCSh
y2zqvlcAm1eq3GMR6phhybqNNAK5z1vf66MgPV1R3lX+gy/JYSyMk97+pb9ecMaL
Nsyt1FG08Ovf4l1eIwzNMD8EjsaO+6a3IHCK6kaTmtmOhTELmQAgSBHQBHv2EdUK
yOIirJOTLTejLIJ6uBnQk5MHylXSt/AYyBz0w4pIspCOaAYLKBuNHUXRHhKQyPCp
EJ+6+/XGF3HIiSci2NBz4FBOFd6h4XXajE17/7T4sR2k04RfNJ5PbuB62nT2WD6T
vhcTcWdGP4Bhxdy1OsJzRvlEziOAc+996zdDyDqLQOu5LSabLNXhSD4oBNk+Vrr3
j+yegfnJKuc7gtpbSFNShAIx/Be/M9tj1Xq+6mkZlnsgd+RH1Ni/CUVAv5Lcy5W1
BjX8dts/BCnYOEEeAXyPiX8BG/IHE3/SlLdYxuzsM6rIKANoXt9PKnRKOmsUhmEe
+10d4+c2S3vwYlbOfg9ewj06ogg9UpF5AmPCOSLlbpdZtwPpniDkiTU4sb+9/BeX
V/B3lWDcmXYWy8GEaX0WhaJO5UqJghvp4t28I9XU6CL/OITCogC4nLRLoDrOmYBB
lAvp4FlyCJ+Kc0WE7rbMHONJhy0IUHp9pg1q2N6BsL66QQGFxHt1vnxyAQTCgbAy
++wSTixsmqPQ1dsllqiiu7Zb47/z1wXGr9X1RP4brxsHXCP3XCtUInXCrXuPBWS6
zZHOVLqLftBWNmZchWt3FxzYYNyF5ydscv3hLQY1dubZow/hKmfqdradT/c32jqk
RtQrm7HYRyXGTqlCwbk9R6wxNcXARJMK2rj3dpPqOSNKCC6g1BoZ7xMomKGHuSpV
bnPrRXGfbudWPL4vyvMntM7EFmTXvWzrKgBiVWKtSFEdG0GDrWpAFS5tE/Tj+CVP
SVdtq2VklxOh4Z8AGw3sSMWOtE6RlwdQ8oYacBj7z8/OipvocO/EQ3sShmABIfoQ
IuQ8SWpfo+LKYBY0WiXEspv4P7DIcpArcnR+puyJgX697jVb7Nt5PdAwi6GyXEvj
mrYa/HRadsJxej88wkHffz1jQI72TlggsZ+JhDDBos+qos+TGkder+jjModiDust
rn2B0kh+otnN4jGlSvQmx62HIsltn6rhJxfHO+Iwtqw9PperGlyan+z8FM6yo+pM
8mwb7P92xI26c1FNfkgxmZrou2nk7lBHa89Tr4eBkEM89sI/eEQ9aLiInsTIpENL
LWmCN7TWyTeVAJD37HRsMg4Vx8fsueC27fzewnd3n1OI/qCbZPji9gbwffmC3vdR
wM4C9KzrS+o1dX6eV3FXhb5CAguVCSP561NHxi/hsG+pUFCA4KInztlCD1YDuNbT
xSV/ZqY7PNyuWOMudVXUYEIOvUQfR3H1gVv8+Y8aoinUEJNcWtzg4yVQ+DGTDzXy
FEu46oULVoYoSvkBcWCJvNJvkoYlDWPDN9zi1QCI2lnZrmyaRwfjnGXop6y7NtrP
iwn+OddwoLanPBd1a/SI7tos0DOql57m7B3TyQJ5JaFPVsLFEoaOHNRkQBkCUddz
BxChFiWNm6wNWp6dKJXbOkxBVmY+pGb9HASwGbuM8XDLb/vLw13x/k284NwyaqKc
lJ+Rj1cpKiNJ9KeyPC43V9ifPf7HvjwxhsLs3CEGBstfJsndmGF54NaQfvinoKSH
DvXs+8m0xcv8PSCi0vIquBO2jbo5RjLYwmtHuleNzPIYrMYAQdCJXbFXooRS7AQk
/3GSTfhFzGoiT2aVDsus9+cFI44bLOMeqj6P2b53P4WyIH9k6iQAZH9HniOrnn4Z
+5+NTxCGJOUbr3r2gXcVNa5aGPKfKSI7qO8btu/qf1P1Qej0dWgTKsEXe8Ld5vmq
W5fQb5ITmHCb9jN29S3lcQoUggXv4Vkr4zcrPZutrd4xv5+MebMdNJum1LMbRdPn
X99ZbUoFHi7jtSCKZixxxe8M/G0+6j60gZ6w/5D2gJEfQSMLnF6WcTtyf04cBnxy
RRuQR1U2B3K9Inw14ZxuYvS7JdIBOAzmMm7LQPMrxMTMHkthqzLMnrOreKcuQcqu
/vx/47GrHGGfu1t8S9jppO26gnvUScBmXYJSY4RNTDcu5oqf2nPxc/JCpvoX/CX8
awAAVc29H1BPAZH57LyoS2BrDhvz+73HPfe4xGZbNZ+2HMTz1hp0jIM8+D/fS/p1
YUDxGpqnGX6Ftr70ZGB/no7LGhh7/tEEgZNd923xqRFZ/wy12fPKZuY6/26MCu3B
3fl+RWygG9voK0wfn3001UAlSTShepI/DP20tkLEyS2sPy+LtoOUbhoylCMZE5iq
0LSvPlzdH8QtAoLUbw/oFFGh7TfsEP7t43+AbQn6PdV7AG4l+RWLDZwu6Kab4R8C
FJRMexp3rW607iC2l3Jvu7vTg/jLrwG7KVv7ixHFvLr3s1WI+mUMIB0qFlBW7TGC
EF8kEI3/wKqQ5s8IcqvqSlhzqUxBXsHjbp2qUMM/Zc+9zfvsOnzsfqbfG7YbOY+m
iIVrr2bVwUR1sWzcw+KpC40wiMSJPoq0L2zU2rhithI5WEnQRg83IhLN3AR1Hv5e
Ym8evbALQyuVZF3PBJq7BeHIy3OliBCBRI2hZhsMslCUhOoKQ/mnsEH1If0YEnct
PycWDhmRFjcF191qXO04Jzwf1T7OhG/L8E1RLALnrvckN+Jqxk9n95Oy+0+YUe8q
OvZNdYDh9Py+sulGpKabxOFO8Lnnk70E5mtCxzAkXC2B42R4LEQEmjus9wg3xSah
jt1kXKVd5msB5PxzTqoh7Al7p1WZewOfJcBCg7TmN1zgtAsuGPw2K/BaEtFoVuLp
CmRq2VMBFiaCQdly3/N6F7PXkbBK5ETyxHS6DouCfGCUA8FFArBTTB7QBcVgGSC7
DRLzp2wiOGXSVtYDPHaoyvYkmsKh8ZcMGrYUaDcILpTiZOnDbKlleA4Pp8k973A2
zd1P3++lLHjGKFTnPLB5nMYv7uxngiVJJkvqbFC/c/7Jmc4qXMs/DfYYzujMMkok
7qGf6/sfVJc9g6JgvDy+g7aiL0JwCIlgApnwfTgoJD+KbUBkByrGoSn5XFZHRLBH
QaSwWHQCDX0cXBRMoXtQCKePHtgv1UkAhJEiUnIyhzo6a2L9DGCj9OJsSMFlI1GA
U8bOY4V/cUOSYxNrAl6Fh3lNAOsPYfTfX8+cmGDLjT2givU6zulgWFKK9RYSs3ez
qukAObhjxmoZX5Z1nlYDK4cBworYw7eNKHojovKq7gyGCVvTq+fighGvQ05FGGBb
8+AkYVdNDfHrvCdd6JJhuhPKHEsUSm0kr/FXKKcTYiSky28DLQ0eJ9h9E1rm/bYz
4YLtSECj4Wu5JkzFl9wvIOLnSXeHhyUfIT9L/zfYO0FYhb7HG5dWr3QyAww+5XZj
5CJThEmTf6BHWQOSa6H51uFjecpTbDXmcN2nW1bh+NqZLncsaK6xGLqK+mU63xaZ
POfQ6BKDq8+ipnlNHauT4VejCR6kSIXZ6IEdURJCn3wypGNofnh1iVTYehvAf6z+
h3KwRfPSuUeDspwv7VksVFECGlixDnXrBblQFgx1G3bfUjZnHA2SB/uvldxkTsKL
GjmzbQvBtU6jO9OX9mWtZc1wB+M5U5IV5+M+d7K3/RwDT3psjsfLb0dHE1tXPYN4
FQHB6g75Pd8CFbRgLGohsrdpjterjwOwOGE6drzL4X5KqtNrFkOWtxVpMYOiEg4H
T1Zn8YHvTta4opx1kTN2qAnuoJAOSwiXYbpbJvVlVyyFmD2mkakACZOEsHC3GZPb
QdG2zpeOM6ERqg4Z5WS0cD13ijjU0drNeQ0mjGXqsgt/kKWv/ck6DQtI4OFn30b1
P85sGIeGqP+8qukp5Iq9geb0ZZc0Q91gecUqEjShqSDU+OHaMmpI6Wu5nhSpkcXB
r/6PI4KhdeuDsKGWfw3ovI6yfo5bpwDvy3yPW5zmp6Qbky0oLu25fo1vXdZTlEpp
3wpNEfQ0wI9AxiHxDsEizbBJYxYTrFoMY/cZ5NL1EeBf8s8FB1k20G8jMGZ539oL
Io3nBgDnYJuwM1AeRME4EhT817p4RNXjnBeTKU/WFhF8Z/9VaaHxWsB4tde78u4E
/J5qICAE0/DI6W/xzw44MzAtl8h1Hx7SL6EjzOW55H6CZdg3YxpLWNwRzdtXYdaP
aIRc5sMcIkL1cSFVIvv/JYXf7lRRD9Z7QlSXb3cHxjL4Q0tLmEyX/tMCZ5m61fEB
qwW5yS3QiYC+HPoGgTd0V/etfNy5ZHzFU+XeLlRTt/F/jEMK0+gkdzPOja8KvQM3
7ygvEz8ymYm+z+XjQaHXaBN+QjID7lzBEF7c1l8Ng3TrkEFrSaObW5u4mbSTMA6l
Efc4c0AuQ0J07ufOA+ibGbkXZeOBaCP8LEyoO+ysI/DwLO52gi1N9ca/9O0zL0/U
LbUZHjnYdNHvz0BujB66IQvjjY6ubaC95EzQrdd6mmKK6jCAmNT56GyEqseTWqtX
fA/IyUwLBnOmqQpcTZ8uKMhT5jR8pbPrd5q4VzUBUZ3ufouvvJz1rUIS900OOO3p
xo+fe9FcVvJvpr/BP0Vy2gGDwxuv3KttbcNMEUyD3S3k77MYhQTu3EZxZBnMhzN9
UEqzr1NlwYnP914CfqGfCDj5VM0cK/f+hTr9WfzAIpF6EidXW0s4g4O2tUgy//vQ
E/rtOHXdIosdQkKiORx72sj3HpLkImybehDs5YwvThdDOqcMqln2NWNwzVrsYHFo
ctA9GJKYe/hrNnF7lK1QcyTqCcKSFJxuSSMRAcH0Cv0oTl4Zd8hSZPaZttmgEhLV
xVJzqVaRRFzQPmzd2wFr1WXOKZ2JNr2Rf4b8oNdaCNbpzGl7kTD4A1k6yuugMXm4
9CxrOqOccl4eQjxBDs0O2JyOJeiLojnsW/xQxv/OjbivK/+chHvNDQXqGoT7QQFD
Lfb0+fAWWR8Lbu4JQ2lrnoj/ly65setYP0mGGpx6A5uFqoEckOATi0oe+Af+3r0g
JO6l5/o5y3wFK0X8+G8zGhzpIyBVRgkG//WEqw/ApsCQizGjJXTcaZlZGmr8VvKl
uIZGJ84yNL8jFYyYhQTv5zLSVpPmnV2nM5PnogOjr8KGCdfXJKh9AJ85RYhSmEAJ
FOtcyCQ/npFWWihfsgWy/Ap4FleWzEmVjD3+0IN6uneUwxYhzhoLoroacLzoM2/9
1B1fbicnDKEB83fSGIeEKmV6/yQsMEDGSa4jm/jReoFvTZi4jj3vmHuSedd/yzRC
jl93YIGJUI8cDN8dcTNSuKQAC2UAZXEKFjFqMItRlAhILFfCD7LwHcwTQa6TYVFq
LGoHiJetyyDzJ79Lgyf5uA75a3S4Mpwrwzrk1fKDbSDs8d00KFK9BAn5UqBFVO+o
6iKRdR2TSkET2iWQJoulxTDy6r7dqi938K2+HQgna8Cwh41KLRNz13abOJREN2lA
cY1lIdJ5sIJgNAF3/X27YtCSjfVe72ONFbUAvmSUQqmdbZKu1RxQb0YaE4fQVRWf
309F9BWtY1/Ajdv4zyqjc+R0CqlAb/hNkSLrGxnDdefazFhN0vp7/6JKrUV2uknI
D3wxcAMY56lY4vDMQhjPwBrPIpYNC5Lh1m2eZtPUC1/kJubKitfMu1AJbnjhP2CV
0oRTAkc2TFXRZEbTokNpt+jEwyeDan1moJz6FL1qSwB4SB2xmfQ4YMpj2+vw7twQ
+DAMu527d75UCcjJVLrtmBa2wSgaX4FVbh+g1z7yjUIJHeIyUoEXtSta7+IVQCLF
A4UP3tWJminrTt2im1AUsQeXkgKYXqUWo+r22zxBI+xWYkzfLZYC0MBvtahITQ78
3K05KOxdAcgMPjxzun2r86s8RCxw2LZWMzZZ4OGb9vJ5n8jBfhLju2C+hUFJdgap
8759e5l504s1jvWw/a+F5OP3h4KpqRXieXsjuCoDkJAT96FXr6gQ0eiKkQDP5M12
dx2TNQ21EvhqadwJI78CbYh19IOFBoVF9wMoz1vzB7vtTct3XH37n5iJkk1Y5LyI
dBtB+fOTuTKU1v6+L+Dr5/khBdGCU9wlqM9kgerBuMfNodS3uUvK9V5aZW1FtpLX
sWALh8tx26icrSFUKPQErFhoRjmYuN0Dc3+jOqCOR9eg3rouFdekVX7o3at0Fzbp
GgQhSvMIlMPWiJv2hs0hC5fekJ0Nj7wYwtlcEOedQrNQUCjzfMbv1UkpV12HXCdU
3aJ+q3OQXGBEBkgCixKpT4Di8ucS1b/sj/BkXPmpejnhezI9y2ILFHsCaSGnfwK7
I9Cz1qf3+bIEflGYMVhFXjzWOYEqKdHFLh3h8e0WVFs/ZfNqaabGLOgRb1xwJ17S
1YtvEBRM1vuib2Y83cwL/eeXuVGeGsarx4kyByk+7sJAKlo/skGlBwIFIplslF0Q
unAQTpwE0QNVjwBfZ2uI2cHYVTM3yI56YStx/swhD2E682FhfTs2WPNSD+dyjPvE
ORs/RrzcY/ZgCr3A58vfqkpfD+jYlBGBrNvv4ZjlyUyW512MuS+jtlJLZ3/TJC4l
61DLNJrbV2Us6pc/cgA8Qprkqja9skgeHxvlK2iukjOAk0tJDPKbkbeLuT4eV2LG
ip1kFlvuCx0UQ+scTkv2cE/njCdLcVPfw4uunGFZXBmzFvDBAKHL+hen1QtIrWC7
1Oz8CQ+fkyihLdHA6DLlAYN+/TJNrNZsebEkHVmALid0ptPSqEgpO88397dPBWMS
xkPA9/rToOw+zu82jbbduRCyYNxh14W4gbZF7bh2ujDJO+KSnyO47qIuKaDEakNH
e94FXU2qjrAevXpVrFMLDyvJa94ClCr0GIWDUnOCWRCXv4os9J1C8bI3uanaemjM
um9IK699k/GlX1XYbIxPVudXBQwFrUI4d4U+TdGLEdG/X7yJgm/NP1P6toJGVxiZ
YhPZzc8dPrckMMDoH5PPnHtKxAKzN9V+OnOG3H31p2yGTBk0mD/GKrm94rX+Uo2z
IqFlTH6GXpoP0Xpmorl0Fncx/fl5Bgfqt6TfxAI6ndog+erpyqUdveTaPWaU2ilm
KOd/KVlhiaNNpHxV4xipdeWksM2fJsuLftFa+K/J551wOrzYTXf3gHMJSigS8IUm
Vz7G4eSmDWRsUYpoVVsRwwekFGkQWRfPuH4VT+B4kkqmOP4gg/kkIH7ZoVdFPeWP
UUqDx1sFVeBvFnAbX3HYyHmJFuR2jmy4/uqKP6D6ZCKCxNIavQjDUYgpCrqhTAok
AXSQ9M6C5+RG8n/76wB8HR08SScaX2JqiHMiEQHvJxUgxaFmMnRgpPrM0W3s46U3
qzhkxxM97o+ArDAFu04NRqrI5BsnZZTMvcDbCj3iO4u1y2Xd/34cqnsj/oD/iwy0
KkecXPjKtnM6NieZA9WLPAlxBbWnIw155BC2fJR+6u40sb+hXXEnGktU3ZOPysJc
vryiqWiAU+KBWmu7begQqnoKvc+l/zAr6A4fgQoOwRbbwZ5LUpRGr2LTdmfFRNHF
6irhTXekac2jo4m88Q4yl6R/gSbelJOTrbsKOImJCK1nsZEmzxFJPJ9yMqIv/msu
v+GBLXrvwcItHCfmiZjJDemI2rEZEfDZjW/T27tRM9i5Z3I3sR/DnIQaRHTcx72L
UT2eddTYh+80fOxa71d5DjrmmmP7rGkYUZ2g2e5sFdQwhLfAx0KKy3iV2wutKEeD
/8rCNx9Qomai8TgYLV6+syMv4u0p1neQ1IQQY1ZCWLP7p+Ws6N93xiCMwfDXVwaj
0CQpStltAhEKAxC34bXh05Zf/S+1o1OM6+LTlzNn6+Rw9E0EEMm6X7fY+FrWEUY4
onhaWQRx5p/+hL4HafHkpC7FeyyikMjbl9a40O3PNmGVDvgDtVi7KOOQDv7I+rUF
A8V2WHVk2JTojTCHt/XkjkTg70XRqCXW37px0kk1cffG9A/hue7E+jQK8tKCdSjU
qmV9QhbA0N3rUJ65vMvyu5/9YEmXumYFRx4TuZjBQMu+WsBQSB1zPh3hRY5xtIjm
cQWbwP28Q4+5iD6hAlmgIpbdm21wK8klXNdVd8dPrx2FMV4MA0egNCeP0Jz3u+Vx
v5XfI0MJpmlYbdQFRQFG5lWE+soaHV1nh+NjPki7gbzeq8qASFjlgjBq+JZRBAG7
Z7k1zfni5vK+T1k2rUteGDBeTH9JOMkmdbVih7GlmnqmavjjUYQSikShQWnRTZXH
gfEvNe8R75ax1gr3VFeFuOxJBdcYzc7sT03vdYaTbTdrLVXeZsWk2L2kGO18Pjwz
sCUA+soVooLZ0WTFeEwwAD2ccYQyEwdDLGnfMUEXvYuJAqnYEDvfEbcteOez2U6Q
q6mtFrLyV7tMHcK1yojCq42ah66/0IbcTbDWccB5eozUNGrMnELqgiDBinDey3j0
SGmcDaSL7c4lwqAcXhHqrqa3Rp1Jtgfody/bagsqRLiMiCjU1lIcKocOdDY954PA
09gKyWtnVD7wPCm1c57EES1to2wa7LuAdGnP92H5Wg+kNfzHpABh0y5jEz/uxsqq
+XTBN1xRWRdwEA4KgnHtIIDOjGHDBcFqSSbfuqiT1jA/Lw/DqJ0GZnGXj9LbsUp5
AdtHV48I4yxnVmoIi0UAzezzMGVRJOpqsQZttTVUydmkaWnOZvqGabSMDIvIbYdv
WbO6lNNEMIYE8qfUNNkBIdBNhDh+n/w2EU6wWBZWUrWkXM7rVetK8phNft5cWoZ1
2fPqJWpu7ZBcD3Vl4gygaVq1rjlyeMsKTS1vbasvj/wc3CRp426X8/tGutVo82Og
0wjf0l4NwopUNEcDSQQCvVDU220kFNIqJQaGbxQAWJZSGmKerUUnbOTeWEG1t3tk
LBurzaAyusDiyAmWUW0T6ZcbrbwfDyRC3Krf+wzyzkG5MJT0Mn1/DwOIjqHMXw8D
nou1M0DmXF7D16kRXqniBSPB5hav2tdypqajQx74Hs/004KUweDxeuvdz6m20CI1
AdovNsS1p37ydX+STnZ4po5jL9IJyY8EKSKMbW6VWir/xEtUFnWkJN18ZutkHCOA
McSiO1ZlSYIQ4uinQ4w02y/2UNOxaPytY15ye0nbneh9VTvxaQjo5rcmF4YdWWak
ypNpSesKRzT2tPiT8l1iB4DhfKD/RCa613lC0WpVoJL7f8iLXuQBfhjx2EbTE4oo
S8m0y9dhAvKnJr10QGniI48bt4gNoy95mBWjJoqRsuExruIfG4BgH8PqIw8PhG2p
eiu8g7BelS19tnl1vHpH5WgeQBiQajnpPskqrsu61ATf1cnqOg4e85R914+fxdGb
`pragma protect end_protected        
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
c8QHULRuoUTBrG3pu2u8/OycVbxk8fPEMGlBCw3Zzlip+m1XGl99/dmmuI70xCQa
loA0NYdhpibreoQYvLASMvHdQYNpvanxH/FVi7BFyBUfjs0UYTzv9udrjE2/h+nl
lqppveY6NwTdIIvH8jAW8OOeSANoF1imScSUuT8VZlo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 235480    )
Poybhjo7pnXgwwa1Y6gnFGn6VWvYzPXAtRkGSuhvkPpR5u54b1Q/xSHm10Ms9KZJ
DNno4V1c2G05NIes1njZrMHQOUEO+M7erfFYPCj+3f2lHhY++JHNENIds8iI6yds
gvBU5w64ifPzdnm/SBs1GtiR5I2AOgF508+sYpBGBMRCaGOKVC3am4N8bGTzy25H
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
TD8VjQa50TFuZb52YIDfjpf6I02fdazGpe5bbKAAnsHjbYU/yYCaZNDvnFntb+oG
uVF6HKv9wVw87qzRDwnfMRDhx+lrReOsZeagnn5RgelTvMLqFUcg5yzWRGn6TwG6
rRWG8ZmYOIJiYWA+i8G/tPOXWB6W4hYV/BqgGsH1CQY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 269556    )
GO/+RwaI/xoqdgMD07rzVBbg5UJuuEM53EuR7vYMeTwZDRp8XpcUBhGHjDThiUdM
a7QS2kF1s4MCFYQQ/4ytMEVSYNmzq4k9n3FN/s8iuPq+WDNOaC8fuubJRRUpOjMO
XG+qf96T9n92o1eLK2dfllmzy/jtxzyKLQw2n1qcYTXCCHGv7F/jQpZIutPcw4al
YmARIBF5ZcnGp699Y1YdpLDyklYQt3kNqRW+xitS9IuHML9/yAL2buu0N/N7ngWD
725WoYOs7HKGjqKXX0wOrb+UHmiPo8s4lp4tB+qUyg1FlFVq32nVH+/xNZhk1mct
MvjOfyRXDpUcQnmENO6EmqCPYVLpIBimFxz6SupgqDvx4a4a1Cwah86eDeeB2FbQ
KntUL1vl16lviGyfwNwuAOQvdTUhWkVsHZwHH6/T46+zH8injoRKTxdMcrqey9jW
ewhNeoL2F4dYRu0ngkul3iyVbw5A/OpNaPdDETC5LIble+fiA+5mDw0Ed3nODttS
Cl3ga4/jVPM1OutnNM/qB5fwcxDvRQhxb8WK/OWURztN3p/PK/u7sjY+ncwDJf48
kMUXybrElvIH348cRX262fxiuMu5mQsRj7BrWIDlOD3RmMHg2ThpT259OMEKrY6O
EDJUvbrXbmZF8Om53o0T5KF0ioGdxl+JrUILYfp49+tCmtl2tbkYRpnVbYegvFIC
8ZMKbhqB7b+y7t8DH82aw2xbAwHRxuuV8R36oRYQkv5LBy3X6qKvmCo+IdZ/XJBk
ng13uF1UTU4qXg1+A1duxfpWKCHXiSTE1CpOCBpnxYvu43y8RAlwoL95j8n2KpMR
743Tglpk61BNewHto81/vHuwk7LhEXsigiLv8+iNAizLGNpVXjOMNB5tuWxgxTgd
GN0AypgU7glXE+aU25ffOVAFbboF8DbiTR5Hy0vt6TQ+euRVJ6qxaxDJZrr2y9wA
jhxo6KtUUi1NZegmdt2XNgM+eyFrsk0zX1JS4tgymWfH6Xbedq8n6ZAkc507pF8L
FPRUJOWas/DSrwSjLXxgnOUqPle2jpciBmsudPwpJDD53CzX+y0QPmtHyWwzVM9Y
kYBWLy8wePmz1APz7HoCwOZG6bBdtjoyt6AbFq3nhIsAj1JmqzXc/EVu5uDNbw9Z
LP2wbYhr6c1jnSwLqv/eUtGAMYMIwD4I7HeYhFiDXR8YsXvpW5TZSJX47u/xL31c
3eLLgbqKov3u6nrfgpauvLGOtmt/EZGQ4jqmutWJH2pocpbX1irzjuatILFVynDh
aSih5z3qRfmEzrjRfo7FurVkiuDl6Gi7Nbp1cVOpzuit7a6Ca460tjvF2ndrjTj3
J87AcCK3LAm/7Xk2hJAgajIQDa7I2Wr+fsS0XE1d5y4guK8oCpLAhjy2ZEzUnkUH
+4gR3psYTeRkyx3SQxHwVY1Owzu5w4rLiA/7SIvSPUC44sC4OmERatgMxR5snrvP
ZuOh+RAB4LUVvPW0qSZcdAhB5ICvpZpDq293Z5bXY3wkFT8P4QTujV/0XX26MjsJ
5xIyTiSYpvfo+LL6EMLpJAsCk8xubNeq6T0hwo04bnBwvAnjF6/uYBXqR0gVM8/5
w/MB/teBrCrhAUgWrLtyCrhqh5+45EG3kxWZZpy0BH+oEq4eoLqF0xlXQGYY1i0l
GC5iERrYYp77CouVCd2MHJR6bHSByjAUSU05g5nI3Rd8jfJVmfcRmQCoqWLI+qY3
GmeAIuGPvWSMnvX+z3K2/5QZE8Ngfyzi9FZbSw6yuD5k76RAk++QlfuMjgdpw6mz
clOUyulGOjwpQfLPFTBk6liy4/sboD/tw9iXHXXaaN2MWVQicHxdPB7M0F2bV2lY
a1gNWmsnm+gMNX785IJZw1ylRoah1loCMcZ6Y/ePO6dWmAbC+qcsY/IgZDb99MW9
SOjWHjDN7MQ/nCCQJqeKjQhlia44ZDj2apfSV2u2gxrzcYqDHP3mwzw7Hih/ivdj
Y/jUU87MGE3ebQ8vYl/7P00Qpf/UQZcYGcXKTqApcYo3r/SnQTNjUUTUBTkmzskn
8ojsmLwyPBIf0dYV+Fjj2HAzs2jUxFq4FzMg0x8L2CgtPciQrV03qL2wQ1nR1Hxy
5KD2yT1oNxRGqsmRB9V1D3LwNEdiw87uFXr7AWhP9lK2lIBSRj0rm+VsU5P7qCt6
0kpmMuJgU1WKySqr9ymuzXhJH6snbir22QEit2zhM4CKADR4eJgUsJquHxGEQQ5D
liTQWfNG3U7DscT8/pKQnEhG8vmCcHrPG8p27o1G63R51mTPqy/XyNXVX9/ei01e
O5zmv4PGIPeNshcZBjOoYTjzkaMB579E43Qb3qg6+GcxBWnFlXNPNCElJl1nL+hk
bfMPuJ0KmUbndWTTAs56emWH7mehrrMAJMNvUh3cyUDPSWHpWwmgq09wMVM05p6q
/y/m+tb/SUPpHk1wHsQP5oMRmphKhberbrwzzv38gfdOGSm4POlqXX6QKbIkK19o
/EK7BWlfU9UxBtGxaCSy3hejbQJwy/8ij6gw+l8d4rXbknvrwOBPfOwFRluhm09Y
h6vEoVOFLq6Jh/9rHKAqJbDCuHrx/r2sahQAtBfoVoT2z7omi4sZ7WfNbYJA28M1
qz9Ugy3mE6IHFfUOviRbsCLxJ5w0Ln5HioVkcTUAHbhUhTkca1t4VX2ekN7T5tbR
j2EEiEJfUa+UXwH3HqFCCUS8hPI5OQwjen4QNpPJTie87TACc6OsuNxWonTOx7yn
5iMSPkpZ0LUSGPgPI7MudPtpEpAbH9ByP2pDT6yg9PeoREbomO0ldI37SnAE93kc
hnNOyhyQidlExilYy8XSEDzbK4EeThvrEasVeTUhabKUBcTGOvqM7lIYHg2ry05c
QuAVgAL1zb1n+y1RiLtod/Tt5DOaoowZvwHc8KIvxw3y2foA25AcU3hBnnwWG7bj
QI2ry72gvV4gIqmRUWLnlO7KXdR5dfIFg02YsLd+nQ1KlkVZ8QSewkyQDtzJZ8TJ
6Jxhh5Sa+XuAnbb80XpnnQH+pj/p2CbJkgpAi6AxJSn+uV2aEZxBc0IaKOuTN0Pc
GLno2rkLSunuvhGczlU6ejHwSniQEgb4FAqvUwVUsRg0sn4TBUztRD7zBbSgclVv
pQWZ+cDeHT8wv//Vv/ojtkc6jxmyNsh5pa30Kg0BVJRSYzKfBkeN0mLPEYnrbxA+
6vyYciaVjOgBrsvsm2rA/flVXQySy+IJ+0JEAqu/VK5uj7NJ1W1fSyhgwqUa5YPL
vuTeXWQzlfFt1rp592iUrYXJcMMIMhY3LheJP0GS4A0Xz21e0tG2JnrTV6FES4hj
n4huBipX12zsit6TuzwAqJjOE+NWszanuau5zfhlu11Vaj4usiZ/i6gb5qg9+VzH
L6gmMNU13LvZHdHkhMxE7ZnOneGrZmr45dC4MrMluuUJOxaOc7nrQu9LXT7bB7Pg
syZjz14z8QCzDXlnsRUWWkRSfMq2wZMsWO774mvBhjDEGgSxuFmIlemTQUyBD23L
fQZxy2YYmFdEIf+yUPYKjVGCsdnrrwQ5oZi3CEXUcCIfivYN+f8lfF8jSu9L1AhO
2oWz7G2qzsnvYzXZX24I3uJeVAx6TLVF0yDpAz6vjgvnRL/kji87N6axzJUALhcu
ozxmcRwn4pIQYsLGAHqixLjx7G/vJJlRkI8clPk2SB0WQqP1oZTNd77u5D2THFyr
SnIgmxppHuQ6/hIS4EeTa7isGP3rRgO7hfBw26DnKFYSVDPbUyV/gpS42tG9qQAX
iSzViYwrNpObwKdC46oEhH93BEdpmPIKoYm3p3BNz4mkCYc0g954zDECX9hKKtdv
3PXGroLocTiH6ec80CZgSpf26RE1pNJ4cGbHA9bE58pJ3MTzLAjl+E86H5q5GXAr
6J/VwlrH9LM08dxn3IOmOEzBh5SfNWoS2AZwRgDyvPKcL7ni92VILwsAqrQgC2Bq
LUrZms1e8OG/1FyJc8JiDc7z0YP0lT7HT6Snly5uHpWb5YkLJ8coTfMi2F0+Wfm9
iERMMxvxqrKUGIuJAteaKniwgso1kaU19KvVZbiunfPuPtS+PlIaxjvL3dPkxDyL
/ZmpSDRVZS+zQRMz0eJPDglIk9CVDPwKh5aD/pxO7hw6plxwIx8t2OUDZ3IWt+Q+
TE9YYS/6iBtEvmHrfQ+hhdVzSQEaW4m9e7McOK2luxFzNpRlZqyAyGYozVwqwnqQ
0+CcEHoEhC0+/QS93ymbSODUHEljm82WEooHHx8EPqVpAtrSHz3vVh1o26thqsqA
BXCh8ErRSo0e2qp2Aq4lYEi4RR0tYIDa86Hzr2u2NFjRHBKQLWF434YUcqXNbqhj
70t62XyseT56UJ5C4pD7Jb85QVGraNpAhuAr9eWw+9E48XRcNpB9rBToKaimyrbt
dS/PTJyqlt2E+CHP16P5XhEGh6IoMPjEZvIGh+HdPcQ0imPvfXDsVqjj0vcXf0T4
w2cjlILH572w3bOLB8JkOPoGVcFhsPaFCNfBagWVa4wehH7rMsp4TqiSt7sAQyH/
iFD8THM4TRngyPAwN4rMIlo7r0NgG4t15pB3UHWKxmxJ5H5XmvfjYnGGF1LTL1AS
l892HtPc+fa9OpNeReNYsjakfpDw+fwGRQRKsUFHZkbjoyIZZ7YWo/wB/s3mHvAV
8Jvw5JadOTwT5xWPxdk7UwAcvQ+xYRJdMmyHSJobFlESo2kpSfR/c50UrnZLpSQf
eVuM7wxc6YswXXJPd3CHmuayz1yu9M/4IUOE1uCKPDLWDKx67m5GVHc8UqlpjDtO
6t5VX0HpxFwm3xjBPaAWhoB4tur1oWxCD2fMun12N9vdO4AbQS1cjoubkoPvz8UK
dPQGKeeJU2Puy+xdiOl6spVF/TCvt4HdLn/PmCe2bSTkPxEjxUZjqzZFcCeu3i1z
dQQ5chM48KwuGsh9VSGQD36WiP3JBGyo6fO4ddo5XHDRrX5FXf8OROKHGYwCo9dk
MZRfgEk/BxD6HpiFnmdrLN7yvM1MpfhF7OA3EB5QDWpDuMbDlhXgno9jqKNmH80v
ISAUSilVU7jmBfofndiDKe9QvJ0+FrbqytCiHCiydMdWK6w7dPJVFohMA960mc6D
QQKJ6KvLsWns4FDx7c+xa8reXYK2Rvl5d6GX0t4nTyoCp1fLCYktpXt4fDbVA4on
4VDhJcDNoyE7qQidi3SPLVSwcbk2TeeYDezO5R9sDr7MMqyDqu1r8lLtKSqWY5W5
gq4fTVxdJKRji8NkDWamnz9SoNEtqxlZmaKidjrnGlLiLCNuws7xIAREj2t8yhk3
9RDIGjs4n8HpwjdYFbji/oiOlug+nBf5v9UTwgQefYLvZ7aW4b4fNuTnzz2Ns53n
RbIZvh4GYn3yas3tUTGZv3lAPrSziu4eYx11+9eaJzhoIcpScfONCcR9Xb0VOGjP
lrF43+fZqRHQhzvn6wDN9V6mjNFOKP5xy7ISl0fklWdQ6EaKthamB4sG6o9awNAt
f/69EaR5oiZr6m4Xip0BP5+l9XoqpLKNsh9aAL76EjSBZP5wNNenZb6Gs0Hvk0Iv
BpzfoqH+0Gl2SaAZRe2h23NFloGZH9iMc7qwLTG1hKAMTbA+jJCm73/I2tW7LRXt
B2xEkE76T4nf92a5PZOkWMKeMhBYoW2Wqham/rDcKwVuCXFm6N2Qpw5psi0tpI+x
6AU+EbyGwnXtnNloziywbiL3mfqyZN5aClapa6GAzkyRU+tIhF/UrJdFUdXKVQq6
K7vpUgzfhs1725iOOiWkveJuk1v2noIAwM7O0ZKpAxbmIb6zzI0cHK6out//gVZz
wtaTZKTQ0MqTscTjKT1X24kyDc7N3NtQv/IqmR9DlxEX3GYVvUNkBIv99sgGxG4r
devgSkjWayUDYOgnZ4IB1bVKgHJ2jqt35RrmzL8cgQb7VKYDjGZ9j8faJfmOMsIG
h6GAFKfecPzVXYpvpI/rcNEKFV/hUjeqknPwKheiQDd1Cl2Ub2W1DudMISPFZkA2
bKNNKR8TrtKZAcM2ORNmURPnlX3ETayELnQmfJyQ/brzpFNcUUHlQwTjUJgxe/oe
s/hjvDOt8Tc9+t/Yt1voJTpVaJGNLcxxz6bi7RgrYgz1jOOtR2RQOoeKOCRIXgfH
5wr8tXK2+9mWhR21e9IOIB3dDfhci6XABoIE5RPZn49FhCuCMBLomO4U7PVxA81H
jq08f6+ocss0aal8z+qZN94ImmINvm4ip1+2YfrVbF/crKljmbfSWQ72R5e7QAyX
FvA7/1/Kalv8K1VeZHA5j1XMqBgV2qQl4ReGTvFmKgj0qe4IiLS4q3SaBwQLUmK8
rfGtc6vR7bHqfScnmKYHvY8WuiZ9VY/pN/uveoXzyfCBAKGobqJygKe3j6shyxod
b9OBNZ/abTpISFyPdg6lhPevEx177+aPmCxbYJ+7Fypd6cLC2DSxqXYjlyCTolUl
3h0rHPXgQgqD9ml0J/Rs12W4XxUIUt28e5HXdzRqkHWsmnTF616g/tCJWbxi1BQt
w+36fN1L2dp+6utK1SbEpO9qD7eJ4P8LQDMwkoox0x/dwF7UdK9LULpKp//QrVBo
4bBgG4sbY6QHnLun2asF8LLicOdvWa/SXvPd8eZBGCzD60Y6k82JFQn5SKP8aBXT
fvCiZnZzYxxeSRa8Pzgh9O/UOhYhSCkow/uRtLAcXh9hjhJiCcF9rMCDk0KY41TC
46FL3cF0n3C9r87NhcmkhjWlbA/001nAvb2imq95NCEf8ztowE+povVMG+CQERpv
Vp2Av7XnsPsar87hweGSCtuw1Ijrrvw1KG8+J2HV4WrwoMc7XMH2oHubTeoZLeFH
S0k8sPUqlKqwgb+5LHIK284uL1Kk7ESGTIEOYIwo4L+oXKseV5vdOkUPKlaJ9LAo
6SGFpK4jcZeANQMQ1DvToXD2MVo7xFGdluaAOgBmKu0wfFdALx8lprfzZxHh2kXh
rEWWlUlLkgEstuoRRsX/SDbQ9p74RaQkquvzYelveBvrmXcmMsB91hdtbtJt8WeH
Dz3I/4UI269hbW39xbXHOklqGYdeJC9xIgxEgeTpMN6Id1sEX6G6m96xAi8kmSbH
h0LDcScGZnAzBJMXfWn6yL8xgL+FF/j3G4ZWqZ/FEXgL7SQ0eGJ8WZuMPxDl092A
P/dN67nEcrdvoT7pcXJpbxS/GalTecAKiyZMgmFUnIlY/gdqG3Ue8AJrx58EcBmF
gwmRn4s0nbAht7tLS6F8ti9oPskblbXUecWzpPdBKuxSKIADYkomRsvX4vGIZ4Lt
zypy7aI/7J6JBdsuvVqiILrssEQ9KQwvH+DSQXLqydYfn38XG36qwGE7Iu9tUpYJ
q6g82xdD3LnMx/Edx0C1Ecgm7Iqyh7+6utDUhHXn94/VZM/Gp5I9lfzJmdUAZ5yo
DraLD4Ap6TC6raZc6LDhpClEwpYtoL43LcWTmBXHeJXuho8kc14T0J3tWBSGzO5P
XgO+5A6lnA7DBA+x9aY7LAMiWO66BoAeVL0cAOkgGBXuxDWn9o0C0eaXhKITBb04
FWPTYj9nPA+UMy+21Ir0j3gsoUBvvjwmWptzp3oIwit4u1n242SJigkFHZYsf3VE
S+ShcJbkgD68XbmAEvYIpUaJfTWmDrTYpUB1is+37Mgz/jjx2o/azDQb+QMwbqTx
tVcPDX8aXxE5Fnv7OdIrYqli+08vP2eNY6HpGwXXZi1/7RAbpABLg07rld4TZ4uB
8vILXuhs2zj/ITNgZr3zBWgPl/72a5mK3HcmXeUPSvP6STg8RZFu6CFnoPP1zjS7
YAAvMJc3voyZJV/dh6NqXNn0zbwCJ0UkWdU8VDAWPBYRv4MMwHxM9G6AGMm4T+dY
cZZQcHaoRamkOooKdxBXRs5SFF04HLXNqQvv1hc0Ffk7OoHrzdCQsL9a2QjtMQSg
XonkjUaKt3RqOsBT7+FWNmsWEhrbQQgPb4TVVBFhEIb+49S6lCCLkEV+VHpCYJeB
ljFw5SOo2AWExFHqAVqLIc4XwyyvTvaScXZwCUp49/zko2KCso+P4ldrKMuXZFMe
B/0XY28dNq1HMutgoUxBvqIgYuZN16uDfLKHoCm/Bw17gb0bXgId832+yt4Hx43q
l9NqLWK3taL6FPSRZjPMWqHdieUo42WOayPynmA2mby4aJAoRcfjyDH2lOguDnfl
0uFrRkURcV1KwgsKQZAZ9xgYY8+8ZKhcQcE322lp+jTx0jQ0ZL/RBEXp5xryWqhY
70itLtIRT73DbRgRaTXs3f25NL6SiolIx82Rye2c2wCsAWq8zs2ZyG4cLLmO0IHU
jIuB3eeobuYTD9/gs4X61Sm3uiek1uLrlBILxjjL9to1rAFHASs+O/+ocD0+i4Z2
67fRKZD6c66AZyRDL/wovDJ8MFRA52uDp5Q2IthzLVc6bXcQh8PcD0ly2aB4ZmfR
jPybYfvBSZ8Dh2/+fKgY7cHc+/FQ9GJfFIe5zTugHQHp60WMpPZw6XC4b9k+SjOq
PnQhQSk81fII5jL1/UlIZELt+o51GDh/7sxs6WI6BxE2J0oLlR5cUnxUo0Wx1oYP
JVKQRvvdewx1JPt+36hx2+vPHkQb20akjais7AMPxxxpR/0LqDJUn9ZM132GGZk/
zdO4uCtz1oS5gZXTLVg1af//pFADJA7PPlTo030bTuBbg60xIVt/XUXmnOAXFj8r
wKQtqm3Nbo2KmW54gyQeWxCXi5hdyHmG8CtBjIuV368XaIWwGrL57aeF719uhFio
bk7ndv8OgfrhFBbUrH4AZD5MFrPmJnFMbtKiDw+yUBQdxv3w5wFfrQipkl4gUzMU
b3HsvWtRsNSH1MOYuan6EHhaC1Cl8MNgK71iS6GQkB9oApgpLJhHAVweVVgFjTGf
wCXpEY1MWWESmYET1EAnl5UC3y3gxQJ/vOvd/mTPnVlg6hxO2OJKJdE7fMOfPxEU
VN19Nus5v0Bw0tWf9HTGPXrE5lbLKXI9jJmZ2h9WiK2iRDxkwoaC3JHdbllABUql
M5tD+eHzh7IRoDRwSN5p9Ur6LNXOgxpxt+W0m9AssxfyMun7ULDYxE3SlAGd8KW0
P39KIrmZqF/1ito/fYs0hop3L1eX7MQD0Xkhv+uD7evY/nbA47IJ1T7ABlqdWw/1
5/11ZvF07y8OphS5RaKK4RcO4Q/j8vPOHTGtrX9eIMmPuVEcrcWTlUJSf2FgqGHO
PThJKJKUZ+7ZNnGOo/F3O8hoSVJ26CFWslrtb3UiCv+3p11X1Sz7ZV915SOBxjdD
o2eMoogNmkhGvuFSZUgLP7/dxRmAiYhRHHMxCWDkXHT8Lt5c/7+mWtn4CkWh2Rbz
zymAV7NctEePId5rWILjitr30/Yk3iWXbkqSDU1NVJyPWkTmqRz/VEccoI2u70I2
mqmnHTjZik4uRwiDBjJdC0vLx4RatS0//thfmsRInUbAK3MNKg0s8vFM3rEv5WE5
INu8gDjYrMK09OoeylSVmuf7shTam7xo+mdZFJ7Ag3F1/oG1o7rxSH2NjgPy6wTD
TFLMtOUigV2NXgN0RnjoVB/zCQb89aca/cW0tuaGwcP+jcp6pvDtjO9qr32wVBZF
PevE00a/6Qw259d0mQ3sDP6G3gE7RZ2JBfJzEychi1f0WSuyBrz/hTmLXVmHO35P
Oc1SW5R8rcGdD/h7hyxtZoCpjscuMeR/O6QFAXpDvPNB3Vgllsq2rdav7Y7Mjuhv
YuEc1PhO/yNS+K1/F0uXehozGw01xCqNx3RV4hhMJ8pbYxWRRCQ3nGPnnyMPjFoR
lqWPsIj2y8JcXddB8x+Bop9XMCgqeomKsGL0Qd4sdXOwUqtdCzZ3KQxrxvtuEdoq
8hpnwo0dzU0u/oFP+OAgaiujRPdKgdX1QK57642dFe2Slx2msWLI3hfxxoYrfVbM
M9Mp/pa1LLDyt+BsH55L/l9RM5acDlqcURfze1UIpLevFv/1dN3ljGLwHkc1ojB3
PH0YiG3MyvISVRrFp0aBShhb4NktQSSmEnbvTtSnu1Uq2t1hA0zaDsvhdpedKt6g
nRQMAGbnHbfRMp18Si5w2n4ngiRd4uDiC2Ne+izhOMESPkPFPagDxflD1UzqbpYo
Yb5Ia/rc3lGZRxsOf0YV/rTZue8FMIeKYxKpF+I9RknHlBploPUyOcjYDIeqcMf3
z9oxe4uPs7JdBfMiHSAjeP0hR0t0j7VwmMi6S4iHAiwQhznYSfJrA9frMtTQiURW
P08h/nlPa3wWGDU5vKCEvY/9uXcsJaQHAKnt/F9c4t5snqU40rvTtQ4RPStVj1ML
F6f3AW2ZbA1ya25JyGbe8KaeQ9eFURTBYR+1xT528nFKk66EZS0MvIHPQUMNwGxC
Znwf1IoisKijr9uGeJ+r+mmRM4KqCi4NcXiLDwdLDJh9HVUJtxQI7bX7k8mRZGT7
ziCgj2W8cZNcHzDebrTvbpc8m7CqV6en1tDcORPx83NrXId836TdQwDcQrao6hF9
583Fm4zOlm9MK0zIlImHI0/bcHPO3qNj7kyzzQDXMGB3jBhQJV0TCV8o5kbiwpcr
s4OaKkVdFPcSV9hAGudBvupXMhFoVLK3tYuIfP84R0mfcTDWJWDymsDGSsOr744P
5mHP1VkUc3BZkaLOlT7+ivz7fd/U3Vd9NWo4TixMYbo3a5NQH186HX6SMfcPU3mt
rDddFTURKQg88EgCxBD7ogWh7iSgRGr2HfGqH1IclzkfBLtNBNWMp/YXXOVu64nY
vidVEZDRfJ04gVBBY+KR/3Xv7NdPGjWM1KaqGUx+rjRoSlF4c3SKHyKte3oLvEDY
879yjIlEpT021oHUovn7PIjGHWPT6UFXJq1mF/wLml+lcd67BCs+d6cYf7wUjr5V
ojjA+fnj1FhKCGzF8OlTPoZ2ne9ElXpPCbBT/KOA8Fb6feATgxaqTrFlFLXkl6V8
0m4sn8gOVSC5yNAv+kC3rZ8PPGb0wo6PWbBDdYXV6uuVsHBSMMJBZ3rRU0eiUr+B
p/8VW22U5rHVhnNSt8VLCG56nRx7tT9RU1mT3eIGdvR+x9nLFLcXmODP4QC2ruGt
9Dzq164VTV1dXo/rdqjYnzraOeOTDNUDAlg147GzqemWZp9uZ21250EIsRkcYwa5
RCKTXZHAAP8dNFeGCOGIozq8BgsbiiHoyGPsn3Rs8Q1lYyC4InbwM8en6ishauRy
pZhA/+d0mUYdEfRs4GxO2flNFBT6tPuoQEamkNNQ+AkDZ5FaAE+Q4IueHGGf+kTM
UyGCHf7yuzMm3xdrcxVPrEcu5mNfDJ81DkfxvP2YZ2nfMHh+i+6oMmKwZhl1QDQG
0Dx40ZW/XUTGakgqMoeT1e+I/zoY51hrqeLkwOu7EpIP/J1lz168Sll3n14W/ele
qgBVEQxtIb7u07NlowGUf5hUH9KlvuAHVyrrwchWM0x028w973kAV8EyxR0DO8SZ
eg2EQ5W1+qvQWlGEDJSHmN7xpmkiBQ8TDc3qG3GwKUHDjU0IRputxy1yiYJAFpQV
TLNpxfRVAKI9fw8dlgxgjxYRAeDS4FyNVMBMMzR3tbhy+gqFS/RqFoQ4U2ohejHP
kFDEetBZ9OrHMkGBtVfaBi3q77L9fCJCQ2Y0VM9lCDMwroUJZib3EqR0/LrHnsd/
JV8XmhKQQBtE8pcgsPN26S+FyNcsufSsDzjFjMuZ18tVizdvpwhIzYy7PaQK8v6X
KG7WlAg1ePxr2YmFVSHj7IXLXiQukjMUBIFooZfN9IzL/JQBCcizGYOWi1EZW//n
SDlpzym41slHKnXbEAK++uYLY17OUeb9V5Rt7KmlFtnObBQg9yYyQ/anCSe4YXS9
OThU2qwScj0m5UceUVSlwwkuXWjZcTmKkOAI6q7DzvGuvZKhoP7FF4TReTRu203G
gGmdq3IzMDQL2PWCaiEziUigSVHBa0CDqPXYoqId1q8Qjid+3V/ahUouql8rWK0F
W8mad07FgLGYJwVPOIGPLVKDaurbFzApxl03ul/DLVzvfL9dmYUIv1ZobYn6Nv9n
Ad0jEop0onGaINsNpy1Y9M3N959UTG360r2p0ucq9QNNdc5oEDrYFBGG1URjSVdJ
k9jxX8e03glQBl+NyR3PASs9WF7yextc9CT0c2XsfnlQFAxLlO+Hf1Nn65kEHRPf
jMrp3mdgq/0bgh7sooQFYUi3O8qAGeXT9TKLGMaptvoSk/ycvULMje4ccp5KZPXz
kOPPUc8pezK901g+qLpIyDw6UxKM+jjSomzcE8GTQbmEQ3kaHvTRNXaSP5MdAML7
Hw8JqILF6J6qRRgPgDRrx9DdWJDmmZczzAFIp62wdH+YGsf07nNlqTsUAP/t3xsw
dMH+dk9mOzkwXJemon++8N3u7aVCPLmULb7ksFjg513Quo0NyfjfcXfejcjxXSkJ
MWQ5umMAXjwxCVZcyab6SG0wOXwlIYL1rKMupM22oGl8TQ8ROcuYTjkJTW+Z5u8K
Lkavr2h3UU9SHicoMhItSoh5atnhOIN+j4mqNwhNn+b+0M9At2BYjbY41f2l904L
hI7aJCWNrxMtKImGxCh0URWP0c7RE9YktGUZMhwfz+6Gtcd+W+C4PFBJt/Tf8sOU
BXKXZ5ZRQuO1ATzonp4R4TnHr7+Asdsi2/vS9UCqZ8f5brKyNoZspsQ+3l9ycXbZ
bVBC9nfcWW5N8RxN/Nfi6xnik1GMluj7fzGQmcUZsPhjYiI5Pwmai0XwqPRCp08C
Eu4MYhoMGc6Knz3fpNwGSfUnbdLtRN/dQOZwmla6X+h97VUdDCFNMzBLL51Vhmzl
T3rQoQlo6vB8XCTe4X670VddHfVlxN2phXvxW920pF4XTSYSQgdDKopmGqBphYAJ
ln3Q5oF6hEs6ngX2xJW7yLhXFC/h6RP9AMVnrc6WYXkQYEyVPY5UIwTEe+dYH6fR
46MLwEYetGDLeuaxKclN8Yio3ieZKSzNSwPrn1zkAqMDI6m4Zy/WEZg5Fe4KdvIu
Jcej6FndzhdOrpSu8iEQawSgvr/iG3U5SkDds9APO4ap6V2iB4EdRBZJw/ea1Vij
4aqElJjxSrh/2C4tHdNH1UA1fP7TsZhQGfAe5VyJr+utfVXzZYT1jZ9BI+NtyJHT
8S7OvaDBVVHAYVf9OI0czwBupMbpdSzEJ728IhaMrEmqqFJD6Z5rNwFq2rxIReDQ
bf8jN0/o58Ujg1qXXWmuG7cvH4BFoOxi2qIOl2L9KQXGI2nKfHSxfQfZdJYXNkOS
9EijB2yA9ur1b0wIQMQp4wiu5N3t/eZBugj4Hreo5uBQPhkjyczhPKu8duDw5Rhs
aJfZLVf2dUyya9ntS74qHtFrz0hs7176xXIAMk9/rBUOX4YMciv/b7ooOG2wVUuW
jta2/IlA53r85pTc4VuiBTMQ+cpsBEglmlfQmJdrpshp4L5eK/XrOcssO5sxTsJl
Dm2CELhRFIOr/PYt2DV6KpPvYiwWsXcyqfBTc0q1BA3fnnR8Xy5qH6nxTDctDxSF
z6OoxooSyUDo8BCzIcOnh9gKCYBv6JJMuOl69sMY4CMbs7Prlu9IG/EIBxE+NiWp
U+dBp0zBXE66DFF9HVOaMlT90y2DVErCEnBaRY1LzxasK3kdy4D628fGOkV05fP5
txAnuhMrSog5h+4vN806MZh8lzBIwOo+YUA4CszQQtyb6f7ZRAMvTIw/5iGvOg9I
CebNNlP+TCSiRFTCtKNmpOS+lGMZWFvPiSVfi09G4Y/1pgUrQ9yz0z3sHfsFA/wY
gzsxdeD/9h7//MAHJDSQy6XL/LS6ECttsxGya6eWQODOKSuIAP79iLdtcbHvEgzF
JIAD8smaeNnFNlGF4IWDefGsk2ESfaUogkAd/OalBFt8/foJcOrbc90IgtLPkWvy
sG3m7T/FgGolohLHE6xsDZcr+Ir7AElMER696ZvyCIHO4SK7Joyeb85bpS/U75qA
U15j7Z5EIhLJJ7G3NAABBEO80uD3ygliBdruaVdoUMDjOoycBLY753WRQTrxZnRV
DxDIuVX3NEpL0M+0r7U+WU6j0PBRduBFHwmIhAZt/KvBKowqpSBNrgBALH3eD/ho
+VpCLAqEGzrO5RGQ+UUbPXjc65be4wqojrvaHkhRRaB6QE3m8tjPeuhBr9q8Fe5K
1q+CZWrWLShsH2cCannvzKEvwFDri8psgv1YNVUSSQOAiwS99QL4hMvfnpd4AU8L
WIDDAtWczhcMK4PGJ23uJ1oEqiAqQHGFjSQdt0dXmXMOgxfmJzBWnmXJ8aVqLFPr
Y+Fs7cbwDG/aH8NCNDo9KQwBjOYStSSWqT1/vFK6+dvMl30Oywvq0fmgN1mMXg8X
UvNRr7nt5BcoWVp++RbRZCOMViHtNJMo86QYIaSVSWIoGUGprQJUZ35yitLpVMvx
m12tT4HiihyLNnpH6RA0vORNPDNf2RR/JsYfYJ2TaDY2yemqPNX8pEC13keJ5Whh
MokhjzqjqIJpLP0PfGAQLLZDROdymYnvETRVaY4fZV6aN8VdDEuCzH7ceRzxYE1I
iUKKMzd5ZS5I5mmr0mr8CPKMgxITFy0OPPGAAduf0vTsO7d+V3PXWtxibi0Q69aD
KdIn3toXCXeoEE4OjDTi3Zbv6JAaALma2xA6CJKRGm++yeXP86Um/ILD0YjTjcY2
KvYxs9kfiqT/doYsjrnGn29tRfSutdHrOXS/8PwENaiGVc3j8hIy9afB/s9eKNPk
dG4BC+DvJ7cRFCDAmZtmc2mZ4Ev+niCtJLxyguxNn8TsRojwByRPXBdh7Sxwauwl
PfCfGVBvbklP4n8ZzqYfQSZgOnEMeISnJj8poF8URM0NyvJfyjAcCJ+jvvxwuFiK
r4uSdhWSaEGLlff5q9PN0jvx+rH0TNna/RDpZyoNsNgZVrZ6tjyPGOep2/Oo8N6q
viJ1zZq0PAFEUuJbMroIWJtwXiWVl6awWBkbXZX82QwpyZBkW9VDOKEVxUFPsmxK
jPpa6KqUAySdpr/iunVP++06sua6f4EQfDcuMencDO6Oes38G8Jg3hIyD0BCDy3z
ZcbxvgGMk1VfA26QV6Gsce4ay7c/qRm90WrEKTbUgpyavl8Z0rPrXEWCHz80bakq
Tw38IG/oqYvnEw+Pm/NIa/rbhxYKhtMw5QsEdCz++/mcJNKkZOdlr2y2F4Gr2r8g
hmMJmzOiOA2LwfJNEsw2/f1S/I3mQw6CKAQSz2LMbjwzzBqQWspaXqKVmDgeU6Vu
owWRHQ3GbfRRSVdIL1qZqyrESE3A63oZkDKu3GOrkNyw8AvFU5ZLpoc9y1vj3Zd5
aSnkvfg1/waXirU3nbh2nkgaxrqVdxroC0yZ8i2DVo2yFzc/6sfG6uzdUCyBglyn
bIbAGzYPUgDvlJ9uS6sEGYaagQJ1XDPnaXcyztr7c3epIK26vLyuQhJ9r7o1Vphe
T8FsViZwVYG0W0ErUXJfQf24Byx0YSxs4FEjriTaCIlZSVVW8lJVKfn1NvVnPTXi
EKRw1hS8b4ok0z8jgzSdcYt5RHCs4hC1XlSQfqOurRhO9JWp/hP+sfug1GVTonn2
uqsIqpSbyyu31fpzDyQ5gkQx6nyeWR6Ca6tVKgNmuM9qSCiiHwiw2JiiaSxwToqp
PQCaE7HPNPxVWKmBUK4dlsLbf1uXSoL0uuNe/lV9g85YkXkqVh0OJwOCRb3QBx9H
heQrTSWp2/4wM1MD2VB9sXQJy7JZZQI5yxKyF9FpeYzH71lxLwnODyHVhjDpTHdv
1tCtj5tooVr69JhgbHguMe8MqFXTNpGdT8pXqO1SHSc/X39NXzSItctQj0I1fzjq
qsp3tOY20maqCrGSRiWKw/WoRMP0IYrJoA5cCvKwwmpF9C0Ikjky3X7Hroh6oSs9
kS834SAElGuXzgSlWacHFhf+GWOYQwwJUJZq+2PR8iUgowL23MQe1a8hzDS75Ye1
MDnujLBc8GaDES3TzJjNTDlZj4AiG4+Nq7k5tsBRMsb5QzZOUXyQHmtRzky4w63F
gTKfnWhJNPghOIy7ykF/sZ8/ZbRORNoMAO7R3yGpWpWTYZgOhaz+5qz9B7kZqlK+
Ap/wDM3HUblisB3Vq8GxcdEAh9ktleV09TAwh1tk1NeziFnH8Z+/RV3jBhubwzNN
gn1mWHy3dU42X5fDAWTMiQERmesrlgldL1dQMG/9m1QE0YFpy5lf2jiPrE1P+uDk
L/D/7wkC5egeVSIxpk48xkodaISoiMOPH9Vfa9d4+MJqx1awP0tacvlCNue+FGA4
vB1moi4UoNlOFkUS7i4lI8CZ/X6bTpTzgo5k59C8++A42QZKwnG8TVZAIOmdVULF
YblKHFpE8rpM8ENtzd7wKffrvpTa7h0WELMVTUZm37S1dkEyUHxgv6tbIYGINXGo
169jbIJ5ofGXwyL0jK6Et85sKxz3fUH5Kf9QyegA5ejE4dFGXT2HoAYSZFDqBOEj
6i6NkrpJlm6mwWETLz1yAf12pfOyKSKEiV5IQU6smeJFcNGNr/UxHHrIzhvA3hwX
P3wRfARGxd+zwoiVJKW4Lip7APJ3+3Z1yXkw5/ZHap6izVBHwTCx6OGR99hdBdwy
8ZoRDHQHLcO1tr19EEvet9pnwzGnZL2EX5+bzB01trtuOdiQlV42RbfPbNVMnuiF
oJoug10ka1+zZ35n4mhTwwcSK/DyiqRjKwtbVHUq9BusrUu5dGI69nhGvaEIKTRc
GKGVAR6FzrJgNLjpFeYRKZ/WpY/vNoe/fclAvt+390xc/arFTLmZkeJCcLBpZssX
UE1F7Vlsn1ZldX0M0junMQGHqPvHHNKEwHi45+2a9goBL1KujIfDWVPTEcfSoK9z
Ru3o7YkBNTixtMnLWAhS9E8SdB2WEC38hAR73/dpwGgDxbLdHFb06/9eEr66ZklG
8j/NwEh7sn5Y3DwihX8A/XqQIeI79o0h9S4+fugxvafk3sOzKwUEPC2sy1j6Bpa3
AYPuvf0ChBMsGAEuGjEfwxFu7Jgcqg/ZGvpkfIpE26x/SD7EKMSskoefumfOfaKi
tx/35q1HuWPVeL6JEWXRnCo5KZl/q1CTEQiNgPNhYbWFCoxQPQ49bYMWokVAElnq
th0xB4bQmwKt6ANVaEpxxEVEqmGleVsyFh7h9Uz7svZiFvERvQK0E3m91bjvmjQb
+cjQ3esio7NfOyvEdaQ+zjl1BxVOcYESW7wfok6G3rN0h9EjpJPiKGbSQ8+7xsA4
rPmZE91zFtUVu9WYLw3OwDAKzp7NzMG+upC2gTGu/5LQ4AlaeblNJQE1QzEMB2qa
mgFgCyd8HuI5Ad8hwU/QdXm6RNRDyYzq9o8fxW5gQnK2ZPbAkRHLhC6hgKarlNKO
N8qsQ5vLV3stuIGZiCUnB1UqT+yi1wWU/5TtoBCWQiUzqCpdwn7dkVkAJfQ4OAYL
boInzu1Y3LaLPORPaZnNX5y7dVQtqMuB3vaeyouinmQNZzw7ipyhmn51HYBrC0gd
90uXDK5DPiEt5hMglnL8alXOmhuoU+CQChBrY2AYjrQeW0Ih+YV8gN6fTlms3OdY
lONwoRJzosNWutrAj2fw/oVKtnNrRj5V6gIv4mV/vzBMk0rjLngNxknvAButjU7A
rFjhFQbQT3eKUYwSsw6jC7giKQZOyaA4Mau5mMfUc+z38bR9VgodbJB03Wotn6p/
Nkh0yMO7AkH+/vMftowe8qMgJNH1wo0rpYdUm6P4DUZzE5vvGLsYOLhBmFSOBnkH
cF+pgfhxx5cwWZd1N/yuaViXXdEvSrOCSM7AY+2keGYPeisV4Xgsh7FcTwU2RU12
ZRje0gwcNFVRO8HmTDVb0ZXCb0AJKbZZ5QePajOHVJusJlt+KjM6a8pOmHKrWJmE
4AFAjZDvEtjNbErW7tKKHSb7gWfi+LHBqm1BwbKmQqbMVmiJIOrIjNE2o0A44em0
oOkTg6oF8m5pCEBewIJnN7r05/YXA77LR2d7LrWLcG+e0hMBA3BB2Xa63q4U8eQW
oav/Jelszt/noTMv4AwQa8fPlq4umcx88fhcvvZGc77uXTlD3tCzCv1RcmLHxWfF
nycGCwzX84FBwEFcgOO9w0HgeUt79H9ZbJO1FlXyXmR6xpUu33YbjJXUXdqDfQAR
5b7cO01Lw2ZI5z8pCRgqUqP17kxGnzsyQJGmsmQ0ZeZHGe2Tr+vyb8R13bWAfCiJ
UktxB04RUXw9/YxoMgT0MHkOXe2Fk/sYg+TaYUrEN1farkxJDoqUunsOkpBHzEhc
4S3wJ0qp/9nBtNQjlOTN8sULQBbncwv32MxkjNbwumHKJrG5VRxQryBgCBFg7Puu
4PXWZMS9uvblUH/TKfUOf3nMW9GkvFBEWywF+HJiw4JGjCU6YYoAXF7ZXgnOVhO3
3BOpUxY480GxmwfbgiWLz0ou8d45GNBYcge2JQ+lGzuM1vo/IvtSwVIFM3WqrPUr
eKEI7H4R15r28T12fdeO54d6KOfyeIi9QCS415B2m9s8Gst4aP4m1sMiHTwNPOSw
+lHQGn9QodylILIvzgOxDPt1INexOrskphfq/dSpMV1Hpy1+2rg16uSAuR5Nz8CF
7MfIUVFssjyITrOL9EWFSpFL/e1I9QpWntc11sNQCMe+T+DiXTnJ1haoDn3WSa22
ZMJUDvIDzD/1kvTC7sptiRfEWkdzLCk0yDuOZLXKRUA/wlStkPJgwN5roEY+LHkt
yzgetYGutkxha7vLvutpzppyhYsvGXZubjwwheMyHfc9fUeLZJmkURddZJYbiAhQ
rW5YaMgAYkpjPp+9B9ed2HQ0TF3AvjtWoeZ4+o8l1O2hiY5u82v1EfCeh8GjwJ2+
u0HSusPj4TKUsg/RCD9TTWcLOGTFFhRQ5CqMzplRg5dpCSxMN/5TYxJuNIaj2xaP
LfcYKYLOqLuEBbK6kcpLg8plVhGVFN+3nUAdMiokGyXthLq/jFyF37O1UqE6rqLB
CzIhOTF88aGBi2upGcG37OXVB95Lr+qVEeEonPYbwkMUTQF9xqW1Z6AVqVZZzBj7
l0ZZyCkVAJem58SIMDiHz+AgWm5WjW7dCl8dDVqSaJZQUqs4Xn33lHpzMC1L7SE+
V5KucKT8SQWVPdRoTfQXlqbxUPAC+nbBZ3UEWM5hWPGRFrt2DkX00iX4nhH+3PQ7
b8H0i1h5HXr0QCrh2jRQcxWrMOFyqHHefRJ+0nKRboF4nauH1OVLiZ/Qa/7nPaG6
1aercud8vmKyG9eDl4Xm/JZuDuW7JlFnOLDbUfDHCa4oOsw7MGDEB7euLpdS7vWj
zhY0BjS/O1RbsIEBiRRyzkgq0TaPflYPwctUKvtS8+Y12JWnc5O0ef1U6r36ttN1
JN/pL//ZxRsASCy2NCCryi0opp2I7RupWSPLbt7nKLZ6nw/wZUeVq/7JpEd2xo7z
N5InLWLWOIGLKP/73D780vReXCxL3+pICeATpwj5LL/SUNSW4FhYcNQbYuw4b122
OoaSXWEn0koWGST7NemXQ8PT5GP3InhiXYqnYyMVSo83urkGGqNy4Z36OdjAS+WG
5hlmh7xADRkn+zEbJ9Ts4irx5PV2NamErkjjVTKmTQH0lepQgO8E1Sa87GWubCKf
6g2WxUzmj+ExZPcWcEiq5gbJC4SB5M2dcAXiArH/mdnKmmfA9C1cLVvk82eyQx/d
Et7b/2aZuWKwOYeGcDoAA4+MkAXtg7iE5GxYEevI3ZmoNtYuweKRfJ3Aql9YDV3Z
PSL8vBafEeLtkCxyRENzdpL5VKQu9q78rvnNs+C9EN+hikZWyhYz2IvK+ss5LMtI
XkdrZCwn8MB1TS5fS4RGAOMwDcBQUWPkgpSbbZrnDLMe1/vBWbDYkNo3DUFJvjv3
X1V2pnSJ9zy4mwCBgl69mlNKqQRZqYuGoDike0GYA6EIYahfC8FMoUEchcq2qH9t
OnuaSwgiwqFLC5ES+SHptyv5l3qSiDff6zhJ63RO7AE5bHXfkXUXf5u7vOaViIkn
izrKsqpnkg1wAsYRSrHn0JlgiMRm4jmwhRBxBnohOvT8JyQq+9PnjfrA9CrEikyz
r7TpoYV02xESM7LKi4g419x0530Uh7sfDGzYynmuTWPllQlFvmkgVpkSGxH9gxj2
fEP4pSu6iMNH6MhP8VNBsWWLNGn4HC0sPVOTTExj7mxGz6Z/Awdyv9nNyrHdBNcI
NiILL/bvBiWlmysToWsXy6JuD4R26kenY0tfwnm3+GRQflVh8vg+hDN1zPwOKumY
ndXUlrOrSq/8NEoKNCwH/lvED8ASXIA7gVbPDqXhrRqLB1yCjLqY/DuxJSzqjYYZ
S3s2QRppza27n+O7swLk3ShFTZhjPEIEoEEqgHsLfxgTzHwWjX/bmXUH7xgLdbg/
entDoFwWWk51iFke5jNHOqOmshTvSD9Kcbv7effz5XqCw5rJxLMPwG8+rL0a7JmR
f9iLdKm3OReLC28jw9Qn9MTiEjlsmGix5v9gbkkVR9YNwx7RyAnvO05l3FqvKCRC
sHm7k8ynhC8tvirlvz7YsWWjYdoDO5QBqPMCkcL+AIg6+RlwB1tHGer2blFlEcNz
x4dEdbcEenysWCVeUfBlVbCehNvvI2YCGNhGgRvsa3mPv+Hhfbob2onr/HaPVXdS
wqXCKMOdbXIjFWxx+SUngkTsZN7azJy6N/nrSssMYD1ggB47VebBl2jFFfyFdNC9
INTkN25OgWVpvVtyUmKPHC0fqntOupPKC8JOYIUQ30S+bJVKIUy/MswVHEpNu1Ei
x0wD/9Jhyv3AnHlCpKZ/ZbrBViLFR4VaCWbzmfnVHXOHzRopyjRXilDBFV6DC8Tl
/92NXGSgYknEFecSttl6w56khk271EwIynTNcu7iQQiRxLFv5pmpFhgM/nDGASpN
/rZC8urN5qXv/oYPwcfYmSYF5AZxytvaT00qFaVDpmRI8kmEOQ5ESkYKAQmPcoD6
RY2z4amwySSD4t5dbhyCE24hJ9MPABnSMaHZfB+pfTEca4DIhqvEBGKA89HGYfvU
GxWTiVXFlagAsBNFUvk7SOLv61F62lwUXfZ0EUTz1BTxvoTEY7OMxfwtPqeJwtHB
kwih3ykjmwylNQ9BnMsGgLvs2T6wFsbpI/QTu/PKfi3VOuFmrYvpS+mmvHX8IHTY
Xp+JJaGMLzV9V0XmZn+lNSSyo2OGJwSoRhS3e5t4Xdfyq2xB6S1RFr0XcnRe4ptj
c+yF9rLF3+IJe3stBDeX8XrOtvy9CGnP5/mIQ5y6XaieEQuiAri9KNzXhksBMd/2
t+wwcMV52uDNRsmgd4QR21X29e2umrY6iwNh5G7HVC4NBmSW/z0ATte8MWxrAYCz
/mS8j/wz/fdOMPHPKn56HTomEZypmzR7DwKhhbhXq9vVfhx9462Ki4/y5UX6oeXL
ahdC3gfiA5h6iQeMxKDdUKJ3Z2aK6RMnXpnAskNyQSttQkQzMZTtZGpNuJNrt4r5
MPlCzBHnpfHLNWv6sSPb48NUziTQ4CaY+sQTfTI7KNVa2F6SU1aFUhNHH+YNfGgW
fLJ6dqyamUCErnFU03jm5J38vPIdPzs9pAaIU+s4fWMECYgZbrOWmqFKkbLgq6He
FOCixovzY8N4sj2FTeAH0Vzeynb9eHP2pbymg4qRPjZNNZ1oBPNTCAEcV4EXjm9f
2VHhdIdtGxr95tH4IGIf9wb+b6yVoGVUt4Oi1ZRO10J51lWtQXRMVmleMbAj7D+O
4O04FXqnK0BgkBg6N0q01i2SuG1+Q5eIC8oBcBG9LDuM+hGdnoN0dwuPz1e6m7z1
mP74ld23Zu2lklLTNYbn3lkLuyqEax6MOCpbgV7tYMPPNTPZMfS8JbRekC8EdA4r
NJRKq29B9IwvscHIT/9oquuOdDQ3FexbN3gaS291y7WhtB/6513qr2aoxtNukEBb
3rYwEHcbwWOAkdiiC+QNmXE/aQCgLeth6ZK3jNhE1V/5AepoaLWNoagxKAowzDUx
uF+MTBncbYqsCWHrH5iJG/x6cP5UKXXwA1kbeu+W7eBvGjbgsE9yfIVOY4NC4DAE
nOu3g90w7QM2Aewxg476GJYxXEVRSIPZ+CXt1/DeRbJBw2QPxmw59zr0CMmJItCJ
JglQ4t5qaS8x0I/rObNqwfl0kowYs8BozrnPaddY1XcqRv1kp6+Y8sufX4K4jjWP
oPi5fEqr62029ZJB0hlUjDFbgAcxolgmcAyoExMgFxiPpdYRpBuVGskkdjQXsQfG
SNiiJlLZKZXqMy48+sJySvLQwfqagBBsPiOcDI/5G+KURwSSx6O2c+Fu/dQIcxiv
amHTwtzAqQHktRhflVPuOk64hLeRLk3jM8msN5qQxlp7yc4O2EejOV+nhGcUh/oh
w3TT+dXvcBae5rvCGdSm1yK/pHy92DqDnTRHpc+vbFOLm8akYnfYyVVo+re0bW+q
deeN1QmHQYfloF5rruFdym8gfAn3BIiW3oplRkLSZUtRDAH3qev6ayOAzxTBuy2+
U4aLGPsCaaqhHlAiYoDfuBhTpwBflQ0YxWWDj3o3DGn2e6jCsvHAnI/103sXiNv1
Q9De/bZXE+PojmW9HhLvMWexkXcxaonTLAN8CaXrVfrUhcFSP2aUqprvoab03oSI
ILaZXuFewMAx1SCGpcMTR4PBANWs1cShUt3AYDgK/MCkOa+6/icOXo6F/kBEjOnO
KV1JFPHuhx0mlnp83uRfRgkGLY4pzzfdSEuHSkasQiBgl5beLmBKD6ODmvkihgqr
nevJro5bdtbOoACQpLHobVhzd7ubfvAnp7CloiPvLR2MQ7uZ8HMexsTGUXYPBpd8
s0L7Mt8A+Bek7ejQ7c+ba0gqfKsq9V6fWWDcdffEsRezBw3uSkAOyBdGrY6kRILR
Fg1wzNAtTki4dpWHRqgSD1vJ2fH/nbAI//hFyQaDoZXBCbYzkgoefzIbYuiXgyH7
Ljg7/CyRBYj/fGfyr1ueFAJLwbwNTGKxJiNXTeCI2c172Kk8h2ulRQS38M6wtSYE
h4ANrtMsuueZrEQ4ihCkaKRjiR5oz3+p3rqrQclJPqO3E9vYdIX5vT5EyJ4KhyJJ
Faw/q7q/ZHYmJHTDHSyzC5JgZcSx9VIqojGqbcY+yXPTvdEPvN5dx8cIBS2Lf8SE
AuyW69CnV4kfA9/wG4Ql5mc9YTdhkUZOH/sKzOh2VeGmqmaJe3aTTBrH8hjx+ASp
xL+rZIbCz6hinAmobx99GfEVxMXHYndvBSxrx9eo+DONYC0SYOyBTPOX6g0Mzs+R
TUk2/MieyEoRh4tIdkkKPKuSE5jQbBqlQKjrslJeBtEkHTmrtMyQpDBP94fjhBmQ
Tib4+zaFVElYd6+arrjRwbbf0DPhoENAMvfMs9O1Hg04HC1izoX9QqRiBp+lDguu
aT66jc+5Gmv6Sbzvn/Jv7G+fPAf3dk8imuU4y99ub299uVvfv+RlwzbPcnXAZ+qs
Us8FcFCBPj7KORAtw1cl5FlAgqPXWUlYw/2p4F1d8et0o31LGTv+9ouoUNHD/U2D
DjrnDYm+anNAl+QuD60ZLKv4U6rOEab08sWpU6c5m+ilJLpoe95X0ooMHD/IQpoc
kYpEEBgEef0GhxqHlLH9gYO5agKaojMzxM4UZfrRe2R5MG4LKo2vXQ1OBGQcgF+h
dMGq/6fOG2JAWV4W1ER1zAuMyxRb8kh8RVpAfwvbrr33CkCm0/y5a8g+k2Es24bG
7HCA59h2FMv+U4dvN5oKERwUhNsmHYbmy49yBcsBvS7xU2eLdnuFurodKsatn9o7
nMKzIxK65x7IS7UZW6D1TI2WMm8JemBwQgroxQla/1QDR10ShihISDqpTbOhFuYd
4p90LPNgtgL8uhlCK24rLtxjH0v8ztGLiRulKxdw8NgugnxspxMF6BQk9xwMHLsi
JnPzYHXVnJk34duFPfAKs3G8tWIkZnMYB3LtcYGi9j6/Y/PjfJ2LaBJOWh5XY4Sj
O6xGQlPvIesFhbTy7uwXhlpFSMdaJWK5t3aBjowea6vZ5B74IHNOnKskXJJGxERD
WvgKbnLpW31OJbkDR9QEPn+xs93ZmxzrwlJLK1VNMLv86J5RUg0l3553l7U21wn9
N9sCtbvrCKzHkCRmXXlZ43RZeLL2iAKEmwMZOXmFTQy3kgPlCtrVdwKL2fjuU5Ln
+akkXsNYpmqcNuiIPjjpIv7aR4ccnOsJtjC99a7BM+iRm1Qpdc5cG1B2ZgxUrqNV
dVI0i5qliOJobSCNVCB0bZusWdndmvN8f8Z6nTMeoKBSNsImXuziEGZpYnKR/pLY
8KKGoLquoA/sdBQxPxG/R/GAg8tntaJ4/P4Cc0JLwrx3WyxsNdR6a7okakvD0W+B
p2LtH7ktTEiLKofPNCas9DRyadMBGxGvctDGWqNgJ1C8ar82OoIgVnc/sMDpLdRC
B+pxbkuVneTYpZ11tegVgO9Vf4gRmnIXhLzKkgVLkmnh6lnuT4ynObcpGyJ+Teyv
gu9AczPrUWQCPVZxk2cSr0JzLPSK6B0PBZHvwZb8UdEDR5exnmyl25NDxTPF9xYa
bHO38lAgGA7rODq9aWtkvnVgotDuX8N+hNW9yBQW7Cc/tm2oqriJDwKDVOlxR2ZK
uw2QWZbcdDexpg+p3rbfBr1iyufBZdmvvJsTOILursXf7h1fm8gzTUl3x9dJaPPN
X/kUVt8WxK15IRxoWyP3G/8zLE4Um+/lWlH9dKDwbLTBq3u0RyTkDLnAm26UpNOW
Dus2ZFx4jJsmH6u7/OrQsviAOrM6TaiWIVoei4fCODP+XLt4jiMoHXXK8Gghko29
c1QKJvJJEzBxuI2Cik42u6BuQwb4uthLgJEEQANz7dmT34lYuoctQK1WPhKnX+5J
CuuiCaqSGqU/PJ4GhyD6LM2M/YSEq115h/H4rhwq/HpfpX4ilEiHcxhke33vVJWR
RlIn9Ete+JW37fgdhoUjmvfuoG43O1GeiHeh4IJn8LUtRhEmOaJoDw8tELHbLGxB
66sEQGdrnZslz44RMkV9TzWy9BmnQrmu0EJpH+1eHIuf/18nHcD1Fxf8ZpAAacTC
sbMTDLM5hTL3rMKxgYfQShjndLPKUadX8YKK9c8vWR51O94Z3g6XUOcx+6VlWHfM
Nu4Psn4nrOqeN6OvHdq4q/OMvCf7EyBeQowDscKWNzer1bbQHw1ef0n21LOVMD3x
QUY2v8YWINNZ4AB7c3J5445wl3yGq6x0Vl9Dqs3EVrR94SDGEz9HWN60NjF2SeIu
W2/vqgwCZfHN6xpwD3Y5kleB4p9V/cKMAx0wZ/7pTt/zXjwLZ1kHtIyloVRJMi/g
lMSVr+lA6BuNwLov+m9LHVhbOaPN7Lq5nT77VXnj3drC2JCtUKNv/fghl24AH3TK
WaO2DOf2yxHaYrXnnMGoLXeSjaLiToLWYZPlFRM+ToI0H5qhZd+kVafmqbAwK33u
h4DQd8Rcwmxnj+fPFwdl9+2vPbYap7PiTK9mNgn3C4fTuHPNRMGb89QB40H8+dF7
SUa2w55+AVUviqVrVNXNuqG71TDalrqxwEMJj/YINarZSSmXg7SiQaAmks6ru/QA
DRPrtfwaaulobbAufExhDJh7O4AYp8dYa0zWUYIVezUIMeSj/YZLXQ7PUE2uqX84
fP67WytHspxI6HYv58jdms+WKJVkgcKhW9yyQCCIwy4v6HIBNjrBoMRp30twyTMi
/j8To/xS5jo/UkVqeGQZkyHg/wwZQ+yT5E4dTqbZ4/eO7/UusuUw58ZMWyUagT/X
hF6jHL9xdbXau+iqX5hpByA+JStiytVBfpRBivrOEKKzBrfh9JieJvrumPwwx/YD
MVh0XNF5l3Q0XXuavt3d4AhtIuIkEZFdono0k+J1/bnh6daTgeQHIjTJjTJsX+VG
XKb/b7eTp6LzIElwtgT6ov5OXwKikT0KkQk/qax1gAb19uiqDl1UPkHebmlOCF9q
ZEiH/IuazdEOWISvam3XjawMrYda1t01sBMaFaZgMlDDKJPjB5XiH5GBrOw2aMpW
gGuwcsbaHVMJhVcu+MS9qw9BWxCtWF6J+1Y0REeyFQyScr8fGX3RHXGp0ikRNlgq
tzhgRHvfQzD8QoSb4rTKYeKEQEd8Dedzrmrb/LKznWOniqlZpj7CpVCnR7l833jM
WtpwjvtOLpuF8CAuagU/O8n74BVsTYmFznKpK4xVd4n27SeiVknECb8yLorUsbnB
htiwhK1qqFqCrbOeAD7t41LFrlzWo6vXGurp4owF6+vnYcSUx8VWy6TWSCJiPQQ/
l8Uz9pthc+J9vdMzhTmdW8tYSfHXB1l9SkS/WcU7ouu0dBWh745BVg2DvzDouGy6
89Hb9r8ywOKWMIIEssiSGqkW2lEhfcss/NzrNiWIMf5MMvc21+jjUNQcLhrXPs/u
3BGYz3KM3jOAybn3QklBcsntB/y8S3/4VLchqRo1GlpRq5KI/P8JcrnJhTlHvW7w
a+LA5DbXpiFuiZYWSH6TI+oORMbOAtp0E8Ulh5xYQZv0+lOv07JuSZ0Buza7Vibm
dQY91udNaZbBPOcdEFr+CtAZm/yulFc1t42VIw6ilexwN+J87GJP41UwYSWQd4vn
v4ttv7wZvcAqTS+4btegddL4Vw0NojNU3nVpiny5uAzzceieCpiLE8KRl0qwB6s5
9NeeYOP1sTRSe7PoB5mrAW5P1jzstlfAMarGRBhYvqsCLa+gR502/BTlCufCOy49
/vUhVeUR8DCblUZ/qcjokOjrn0DMjlA66zD/onRy9LIBAvaA033DFmYrEpXAtzGt
o6enhONEfUfqlfeRGz8TCooY/EfG5Uw5SycnL/8QgkpSn/lIbKLfmzUb6NtIt7YM
rjlI2cJTJjJdZhSBxIPS3q84cx+8nSrJ7Qhuiydm2Ups/hoLR65OW80QOJJ1p0e6
M+JAgIAJaVCS5bhkeBTyVS1tdaTu+GfjilHSfG0NRnn2HbUhzVr1eyYPUiaXXIoK
GnOGUPV1Wz8cGqauQNpQOhVCNE7IWi4yLX1a36s8voV2IgVqidn4MOwzYzND257H
rRdIrwys6//ZrSJesLNwyJ6fTWMK0hAFTe+37BhlMXAZrA8nKdLtsihg+8Hj1IVN
OFELquK7/mf3drautBGWK0b/n4w2zpwnPE8VefprWHvjVbd2eahELdnf6QVwyLx1
HJwoMJb+SsiPAgYJFczaUC+cIs4osgB41ZMVonXdh3o4JWe0H4uQpFv/sADpFFjI
nSttyXT4oHZtjiULL3lK0r7zM4dQDYsCkBeVE0AFJhhEqE3TvqGD4yKyQljK0oDN
BjgQtaoj18195kti6C3dftVxcu2/ebjnlDEUYdS+eQCVxAwCzRWhlF6DWIqosoSR
UxKutVo+VEDWGXC/wjttoBVuAlxkeJBcfgkhWpeJwp0UEPFzfKhMD68Ww7Xw1ygq
Y5FLu9bFfF4ziIt4iWJMxzrhsywxKWup09O57No7LwKE94qpHNjE0P2jKPPHm4wo
lESMhnYOLHx8+/glrUwm5GmHkFjCYbp2INjWwxFaLxwWeQEwoNj3AVMI6JqbohdM
brHLOeghqydNT846Ji7nWufmjyrb/UaqrdzlAjKWETvXt2iZiGqRzjIw0oKGR8S5
D7MYOukb2o8tLHEmUZj/2nUY8tDj5ecZnLGbVIrq8ClBdnUrfzQDCrRuUWl/MFxY
lU600z/qf6OBFWQECDJ1ndqFWEW36lUghrQSG1hc+J9JKbjsHznikdWnJCKdpUJW
tX3m3nsHGNzs5jJBKFZPERfor7iGihZUNK/+qG8qzJLSb+2VysZBhOVEki5HC/Wn
rmz5AOnuI1d98zdjOk4rtYwUYLNQPjEbwL8hv5t2/VbFVtN2q6/9zsR3CJntWRdT
geSAvYmdBCNOZ11SuI28rezOOh8GCsvIkWcRT1qfMURIo+LNQ3VxVwLaPWPQkkB6
MAV7h148AlzbVZxXWfNIz3oKeUiCdTHwiTmqf1sCu96w46pqJ6DBlHpfooOqm23c
2gI6y5ko13pQNKlmX2qJXxfyTPM7mFO+e+Siaiku5tvZTypCB9pn9MIprbU3CNjA
v4e0HkV/GKkjc5i0ZjUo45no+Vjj/nj3fBvHZd7McdSz4ysdbG0L4szAJuqcMGnL
DAc41aizPV+zg7/PLDGRCfLP3Hywl8o5d7v5O1YDc7UVQLxXbpdrtlKVK5sszVDf
pHHn4TBu4hKGUpoODja+Bf4Ee15cS+y51vMrrcUUSyJ2ZbHpPNyZBPxcvshf63Kx
9vzWiMqACjl0JfAUn8NiBjLpP1PNyAzA2MFPwySoMydqzxk3OpuKHZ36rByyCD0Q
yVPV+tI7C7jtu7wCNsir+6WTQUcEpkwDvqCxYuAdqqyycNVAAR4iFRGCyGg0MLs2
TCRYIFzBl61Gib5ofQnm7D0OTwCjY5RMvPbaAqDsJsR49WK3PwQLPad8iHbi82QP
K4uHi7kufSFNJlHQK0kanM/X3KAJFUB1Ju5Fu67eXSyMhui6yLhrFo+0h9Cjkl9X
KKWgqzq4uabm4sjDR4tz6A+BDOUbZ/vCLMYOcZhmvsn2VgA0nFy8w/N9j1HUxluu
TuCYosyBDeppMXHrE6fxETrgGzUOvdg3ezrW/HCVxh/8aeRBWZhl8oLXqxGBKHYS
tY2XX0Z6vruoGQEbKozf9qab5azuArQ7ds2P5oW9NPsAJcrMWrCqEOGnQtpEWGAt
HKAI49h6/SZ8pjbdwLGBNV53Sj0kMYuY7wNMzdRpRGXD49XA61WwtpmCrqi5rJia
W53AOVZmMJi5/fnE3rLpesh60D35hpnrSJT1JZWlBLqzJpVaIVx/DOW21Eb1iMB5
7+bf4cP3lWj0qEdjkM6BLV1yc4Fep7KrbjuKqQNw9ywThk/qtlwdaEwvQVPKSHQu
QB1oCIh/I0N+DoxEvIWTkyrKzSy+IUZrTN97xU4ApKv5J2w0c8NRO2rOl5qAa+TM
587PNcspgdv3azbfP6R+Z7ksnnnuAmZ7Z5Kp8ISVTUd2dFLY+cWW8ytEIY0LJWtF
mrONQoF7yMuXwxYY7lRS82jZYCVmw/gUsKxlbOutkt6EtfP+CIAz6vh5iHoH42RW
Jzq49OUSgv0bOHsTPYPKDKoPZf1nWZatH6QJFj/MaK4bjs5VtvTEoigW0bKqHoEp
fYQnQf/rEMwpw9s6e6CtCGMSoG2Yy+7vCzeZ50HGB0MvsY/VvSUfZwPR4lRSXR5l
lfrVVYoX3N+UKgOPQHKTA2GT4FaLm/Zk3OJ03MkIdcE7hNNLiyQJ2sN4XN64fN88
F2VuFWUhuey2q/VUPyQ+5AvLXO7PrL0o2pTPWC8Vy3roAbKdkVa/KDQ+B9RcNocF
Xus5Relqu3gLMRuYavNn/rnRihsJy/9wmmIg6607KurnZcbiY48ORGLh5eYVwdCo
0UbmamcV1sSrF1w6/nBfXpYTGt/Z3FE2G7LAzxHFXm3sIm+Z93fEVTyUNGarkn0U
lQakopnRI0MMHj9UYNwX4YLBojfSYaYIxWnpezf5mgODgfsVqym3dKri5Uzbt55x
aSDegI1p53WXZzLIBsJ9tJV5gLOZqUMd361kY1WPc6sSv4SHH0O3HgQ6c0pLwM8u
9dd8yBuphnDqJAorU00OVMu8zWwMa+Hk7Vio8Oy1CYclTN+N4z3pTOVwO2M+qrbk
66p/GTjk4Ro3Fqjq5jQKoC8Jls7i2dP/QUbJpAlzYWln4iKnj14DQCuTa4scWvyV
ZtV5UTsveLy/HMRmMls746VgfMgVcA0IG0+xhapPGDBzp6j2x6ZBI5WkPDgOd7p6
vQ29/13DnfI7qdpefVMjbzv0//Wo+awb8bKDU8vCjLliq4+EB/lKhAcDSlneMhXB
uCMzLUqBAmKwGk6rmN+9/M7zyGEuaQbSaU9MB8VRJvu9FSKgqDmN3LuX9l4vYB6X
EdIAQkwJy9XQavi99eBvEKUBEa94tzUvBZWXuplHJjj7bfw4UGAt7EDM8O4+GI/R
a+An5NsQGzI39pYJnUkrQRRTWA26gWRBHjKqQLIMB2bRrEm/xSnnn/Q192gWNCW/
y43UkjflnJiax6loIJZ/ho/Aeb+Q3MUBcPal3aJ66mOjqDgGxBYOfyeuw0rs3k/P
fFKbVIqAO7N9G8n3dyqyFUFPWv/7dKDMJ5+Wo/1jZc2QBPCS4ZAtFIASjwJIyKMr
Rr63VIzGErUitM5I9+X6TNEf9Uhk9CKw1AXHcfnfFhogXIahybGhQwdK4ORJjlrS
kIlKRRJ61m/N/+7z0Gj1LdQT810alrPWgiXoqofC2CsQBe4mlhQ1G6BcajV+ughF
OtrUVjja31Nyn/5sooBoSYDFMJ8RLgVhvjzc/zdhTvnob0RaRoAAsEajx+LpLLT1
+vzwVoiTYx8IKKdwkZkAokx2yxNzQ2M6qfKZE7Vbm+jHe1dPmxvq1KqaFowq9ezr
4P4uxz0AlROSIZhi0cwZ1xKw5xxrKwduKjUDtdJhP2KhM8cF0qkmhlNnJa80NNVt
q9jc9s8gDnLues8rm85H3GOAQceumL6Lnq7n/HCanJn54X7Ti/9+X2hgiQbMRdd0
lTNgiBh3iLjZ0zEmcF1aPfIipw0v0gVVzkKvzLn0qoKhr3A25P2qr4HBpjXLkqR8
ht3wWTQw+IQ4A9RMh57+bznxcm+SVm7qZdrQR12e8ysG5oi5WlhWMSiVwkZUhLkR
31SCKVyxDhMi9ZMo30P8ttM6611tDPeSo996hPsgDsQ/++tIAcAZXZb+pKxO5IKV
ByTtbVehO9S/cUq+tr6kWDuvWiMYLA9vx06zTkCPHtqRK6HSTwyL/s93NYpqxxWy
MqafcD2qI6+n8IlKz5mMLyAkvFY+jRmA1wd1XMxgZDhHsLUnXIj+gg6T530jEMBO
ePu9SQoSjgh2E5wqPe3LkYqtuRZ/PDxQQaC7KA2Thd7AN9oDjatn+u0a+BAOy9WE
pZvK0xziujDcFKMgihcXBuF/yuO93bZEjjWvfbS12loBjL2IWBvXKFhqnGQdxc6T
nrDM+4xXgLb95+aY4i6wN3lkS+8Oq1RWNeGUqXO6AkR9+UJHYjRrB6/ecZQMKaTx
vzzLBQsdWFTmini1/zNBsm4XaRmkDWEthxj3r2p8IV10ySb6HtC5v1i+T3mIvVHq
6A/UQ00+s6LaIiT+R+ZFkYrLBub954UsD5IkrRVwZsaRGKGlHwdntLjHzYObR4SL
VpRILIwwdUVGrtBb7qBT5+YuISk32ETtUVyK/ws8r3y2f8MvFPUguBjZT4rFNe34
erzXiXXedWKJx7OU2EBI9meWDO1rgNE95K5haK0vl7uxLGFUD5Oe2aYssX2kN5+8
qpe03FLDTEgCk099luUylXVdg907+D+SdcOF6R+6pwPX4C+GdrEvomwyepDTiEWV
uGKI7cdECRAyGHA8rGCpFpaFcP58epLnd7gMs8Q44RWoBDD4YbqOeCt/IOPkoT/m
RXiTAa9U77AldammRRWOSSeQX2cSvc+gBVV+9bTj7z5Qts8dv4ipI5ccE6DqL4PL
reovMC8zrJcrD4UrfpGzXA1PMftUwWnwtTmCJL0q29ByZZRXjRkz+D5t8Iuuu9/n
zQHsOuf30dM6g7lOl37UkiaHZgOhKTNDnJwPyiif01P9CaXcROs3dVDBoMDQvaLL
jAkgOjj2qEOUp8+yvoQVXtI5n5M7t846cETptzJnaC1se9KF2If6tWhVIQi8givG
0cSz9KcIvOB7lcYtxma6/J6KKWLO8j2ojJDXmoS3VF3sTCdbNB+N6sLG1ZcfKBOY
oUT8XxXBxXTNZ0f+aEvcRCtlnYxFPwNu+OGJ68YXO1ChoxL1j2vIjpAAjbpkrmxL
FEIx3fnlBg/C/VdOvkbJ4DKYHIl0bvVn1V0BwNOOm1DevNbD30zkwRoggMbrqaq8
RlZKGuNJTqjtrBZcF8tFYNtjQHAdqG3iwCbOba1S4prcAG1X5eGszbVpiv5tZPd5
d1KXTXg5xpsqDrvXjcDLDilqwsZDl7ARh+UfmoG/IxxZ90YtKBpUllFHfu4qf6ln
FAUi7B7qxZOxHTWwpoCOkI8wp9P7+suPBHTrKOmRxQudM06infykRX9FwR6o6JVc
hQjoGcZBRykq5HP6ZLJjeO46XWHdutCMFPE9yYL+EZWhteTDMXIAhbjAahZKTmoT
6IzWosBi9o06In+9dGB4CQ+8EiWTMOodOLuwKAbzpzN9eLNVarpOzvfkFjaSOaAJ
NIOeqZS7ppjexX5tHFJgah1EzFJCN6XLTCWUyzwSKH84V0evDMAyPoNbn60anOd+
cN+KRqYLyzXy1eNCPMqZVWn2qEGtiLfzuSerd+F9u+kl7LElnqYd9UGp/Y7RDsX0
32cMZTg1NiNNv6cV/WBwfhiC9b9/pC6F3/s9cCLKjJloCSIMsXLosYJx/gyLTSHK
Ep21irCMdQTXgT/uaCooeSlP8ch4qAlXhwfVNmkvfL3ar8Uxy5I79puMvmb7bxdb
4YNzQ2I+7IhP/qrbJ++5DqtWXEH95EdQ7F9gdoZsYPl8mnXNPHL4A1YmCCHJG6DY
9STxoesorwB65OTrhPMR+o/5iHwOL2ZSJivhCfBj4ZK+Kbm1ofNvOynJUkVOcjQw
b7P+ZIt3fFW8JgcbLe6m0fe39ZUXm3z2uKlp+ea8DXURJRNuwi3FGeNjrAX6EEWB
0Mcnc9pa+slh5y2EnSHiFQSOEdNeks5fElnHbG/dS7G/2QpLg1M/AgiS30EhRstP
smogLqoW8mlgrcL98OcKxXgzt4Yq3jK+Vx7PUMRPv5SweU99Cp0DqYZTNx+NFKRg
G4GvMHgMCbZIWkSt/XSTOeYPdqJbRowS7KsWv8YgLOSEbvmxOO6vdscLuzTeBzqs
Ot3NLHnZxye9dLqV6tj4wRENNx68uEs01CWbcQIYfS/08d2TKUIx5BsF8SOmXeaz
eEPzBHd/9SLjyLO4bp2Zq8QgHaaZad1gder2geYMyx5lSHvgg5Hh5AAcOu0t7i6g
sPmij/imyFw/0lCs1IDEdWe40ry2Q22moSn4YYonpMeAcTc9Qgal6UARLtvC3IuS
2u7SHEo+wqmVNAmx412fB1J1PV+2S/TjCdKWqFkbDWkkUmdwN0AzVy10duDacHaT
AYtdXzmZkHXeydKi6PNUYEfzzMYumzIlDP1FU5S838pWB2U7Cvkd0qTgZPy8ses0
4Bbkf9T2KZH02NA4edKjoj5MOqpRBqBYBc0c8F1Tg8WtNV72iS0a/eEJMuTQSMMt
uB5DT/kQ1O97CAdeckUe9G1sc4x3TqbH3xE0esaVFwPnyQwC5g5BOrUY2r67Acgy
A58dQT1S0k93t4K+MQXj3iACrKDYyw3hcLqF8GxzOBzaJM7ev+IeXkg/n5svxngA
S92F0zA0I3Z4kHIzqC6RYILe3yY04cluWOFKc838MSpuVRzytAw8RRyNjVY9l44F
BU2tZZqSHlhqfgbtzoA/+I9IvfTV/7G0NEz95lINzV6omJ0R+ZJGqfV305fGaqEm
4FPmdRKpvBKWcArgHrFsZOKGKBtpHrriSqpuU/naEsKo0S1iWwtFnpeRLmdCmpAd
KGMBUNVBV9jD8l/f5htfp2RPXW+0wdAOaq/S6S50R2Ij1fHwYdxLxlv+sFqE7xdq
Kg5d0opw3sOZObm7C610cNk9xwEdJUwwVUXlS7+PJQIKaMkLTJy8k50aFm7TBO+f
IBR8SbFls/0KPqRHGBEDZrXfPs+ogsgJ/N1nHaD08JAY0NAdAz1+YOP7v++qa3eR
U38F42YKHli1fkxIL4OtM85Pz+wlFBZzgGPFLwg0FBFdzHiONs6zTdBJnAQjHGqi
Cw+oHfNSE9iHWvXUpjNzCIomf/c0zzOJX+0dNlbHbPVQwiMOXkKbGZcvKIYXKxcz
HW99XipQJn1z1uRfSk2RAWbrZjRgcA6GXxPa1k6hdpMHHH5f/G3YF9jKSB5N7HOE
cp4fHNuVK8rLWH6IFzfyyEG2BDgrCQHRbg6lTTe2D5JGEnn9Nda3/zPBTG7IdgeB
doKxFNqUPTRywqhWT/QfXyxL7/R5RyglL+MFu8mF04TJX8B3BLpp+FSqt5TL7YoY
yI2aS8QLbK1EZbfC8uvQF5C2zac2PHUe2Z5J1fL1Unt74WnYOTaN9rLToIaC3xPo
rFWo+mJBkePRwrglb0um0EDkmargVpT8H9RINFgyRc6DQoajDd/L+/dpsmnmL4IH
q24XLxlIMt3g8xlnYnweol1u1AnI7GwWWnSyG/jS0XrqkkjJAc2MmQI9KsBBl8X0
K51YQ9291/UEhAfoZ3KOUUqdT6ewcJciHxnr4OKkOSIRk6tuh6BF6KZy2wWGhbK1
oJMBNCCC1Md5dJwcOXJwGDtPbBBdT7+sQcRL2yp5e0o4e0krL8vxucgRbdbGChbg
VWJdSveRFB1/wfzAiZJu/teRLbIJs+h54wvEMIkZWCiePzyNlVImG9hPLAII8w9v
L8NG+J/nbO9GzlNxvTcOEKmzVFE3xfmrbpbdiUzZnUcPnX7PEBTFxMClJ25Roa43
7PAKhrEkaPyOirBgig+Wax1ObC7+UYXhdxleEe4AxAhnrpez1iHIKwj7VcJjAteW
RngLP/QyMOKMOI4HDeeJxIo/mViC9bEerdyNjKQ03IbaU3Rp8tXetensTwNSr9ND
SJueo0uLOzYdaSxTlYOUHzCVKtJi7cN/Fmf/iqNP5u1X5qMCAHGhUwRaiZcsnmIj
PEGZBX5irxw4J7dU195Vrnh7Q3dneVFSw083aK999ZZiSLFnuurIJR9Gnx4gpZbP
aJUB4L26SWBKHPpew/ePL2H2ZO/y1o3bkvR3px5jISqeFlCgAMbkMIxMGvAENrfd
VWwQWznRTBru2USmJ3P7LlOslWPcpi6VAiVlTTiM99Ow997S0C2fDrypZGFzKK5N
ssh0y2Uc1Lyv3sCSUkfkLDUheBPXIIM8O7QzTUKxXACPyzOn27MsVLYD7SjMjXrx
Sc99N7i4HTbXyHT67NB8GZZotsnTwZbjJq7jH/IqAYaTf9OZChCyXSIhQ9CRuBfQ
uLyq5pqWhxkWdj2l/gYT19sv24yvU5sWg7lnLsjfmoJmg1z1mEA8MBUFQ/fBUR0z
raAEartNDXRtTbs1+DHDhZihxZ/5y1Om714pjQ8w/iOaW9BL8AP9OaGoe8eZPy0E
1/Lk1t8EhrBMuWdNS6NjQK5zWjIPeWb7aFc+X9jj132hY9OJgLbeVBZSt/crc4dU
XrN6hZoxMlDo5AgzN5JGIGq7N+vpGBIW6RMAYv0vGNsx7i+7uLCrl9qCTg/n50uw
wlZZTSDrwMRvo0FHuoQmmzxko5rXVyCG58bu3JOvf4weWcn8thkKHF8kNDz1FlGE
RgZcRFvDF1MkzVOYsExhKwCnPaC6FDl7vAS3tjLdHUuTE+lPgCtD2GSIbTNGzxuD
QRKhYdZF+A0ru+qVNmUi/Hi8EshXkO2oDKNXDWMXOgEQFbXbmdBI6RCj+DEDWvNe
m4kWk4H8pzvf6QPmtNE2K6Ia1w8aUT6swJXTsSavewcYFd/yLaRUhhXlN0KlXX2C
l6fsTYaxCVKyL1q1ew/kctAd1ebsMx8HWgbKriAuOgWVvdHV7g4Yo2qCLs0eLPkG
PO6fmTO7LooUHAJnFTL2pu2SaJxnMMkC705bBgkq/sPKihqoXpPrXzbV6cR1z9x0
8oj9QK+xCz/u63AqexKwZKBvpDI7vQy5w32Cj6R1DtRzarhQ5y3k96bicMZWDTjE
b9pHN6VwcNyYK6xaCqBNJ+/4ElYPp5V78XJR51sY6gRGD3IqIZXh4WS+3+OrYfTB
lNDn8JvVZKXPOQlgl0MIgMar+M9gTNs8Kcjlaj5j/gLaSM8M3mwW1Ssm1nYuSCjt
eMsc1ps7HWJvWC0Mlu3dlaGvpX+CBEUqbv9QuY2qkd7UFlpdkGzzWBKlCLMdUxb6
eb1RzUENuL7qTA6CTQkS6J7I2Wiji3hbor0NBlbsCPp49DD8ecBrYGufTJNnT5HV
iy2uoLr1iwjwKWemfVSbGjxA4ObFnGQ8XNOMhg10IlWMzXarWfqGd3e77S6dbd+X
IrfArPpcU7hqbq1cuAMV7iz8MHK+9Hi4rn4RY98nYFeesEsNiPhzLMbwuO7F0SFu
fLx5vPpZ5KE0FkgUu/2v8SLAU+FhUXDFsvfvY2pvJRFePEKRJo+76sAr8k/3sv62
rwO+qANx3uBTnK9qDfBxEAJ8D5WSu3/BNNoebNx7A//dA4JG1uYoq3z5PrUElXxG
82FimwYZqizKE7KI+ggLyE6kRMo5KHtEOO5UENu9FeFwbh2eMEl+yOgW0EhV2Tam
WSTpWu7gG2FuajpB73ADcqHZrMNhxPTWr50c0EmaxmYCNpstA3vXWKZCBnHEXHBB
TfKQCKXdVawimp8U1qH7IWh8iPGjhyzstsjDSsi373ueVdomxWxCFlvXrPUE+dTm
vqe+E5d+43unrknZ8KIcMsVF1n0ozB/NkxTJLlBXkSocb+6k/BV3zYNs0+B5+Lt8
ToTHQNv/vvB+ZH1tAITqZAYnyeOF7G6F8hrey8Rst2xGcvCAVsx/V9ktNHJu1McC
c+SJbMahePZWVIkTz023ebNLIgxuNjAtCxVu16XMVA7ikOqHfxQhn/5qkPHLeeXr
2DVeT/z2pa7/EHNztqbb+k4bybxp17cOOhhhx4okLMjQpmPTTskorZAJEOtgAJum
n7Mi+kje/30kWME2fHMCqET5HnH1TQwzpDB0TW89T0oDkycfAOiYuXPlRzeOcRj0
mi0+hYUcdqgpbUFbvmMarAxSmpH50B3G+vj+ZHYC2Hqa9P9snopyp/YDinxgSYtT
zwNumYNYfsbFfIwGv7zrT9hGGtiX21JE+n9i07xG/eAeWGSitNsKgWv+xAHwTVAK
4R8yaZKifYZRLv4A2D5bN9vBQRdsqBuchEWvU2zciPj/3OHTYYp4aPaYSpyapX94
eNU1i4qQlBUA4P/qJDHXYi9mg8gaYuXx4mjmf2kNfBgDHqSy5ebCBlNQzDH54TaX
Ki4c41ff232x7AhAztt1wJoKNjoP+tXl/FBnvFH1k8vSqZQ/MeZewaHANwu53XVG
RS1MOshhC2NSteec2rD2WxkKzp6vIirgqEZtfYkYTedyRDjcVcoz+b7ML50fIh3a
dNJJlLY3L/lms6yccdtknlXXNpDbCRn9cfhlW4lgNb05X6wXat0a/wrHv80OmzjS
kW2iVxHOmDxzQq3qw22J/5frSQPIJWaZXd0ZFn5gjLLi1LI79q/IPkSBqNV9ZGx9
hY+XhjPprpRWxmma0rkhp5w1M4tHdJpAlbJciDarvfkyo6HmSKBBtMKDcZyINRnU
oZ1DH70RPFTlLtTZwXFsMtZTZtMdTqx5cmbaYL3A/BU07XydvdA+ED1QXM0DeFmm
NA4YHTzckz1wL2eD3WUc8Ehpsc+tAk4Ic89hyTeaaWiacZ+uekjlJwrwkYTaZWah
d3hCHubkhDGD1Zyg12mqxAF1nJAoB292258yekTua9dDKCYFvYjH4CrndTmBxacJ
/qX1p+ZXHTT6+uQ5AJICve8zu/tdKC8A9ivtW5HJibBlnc+zVJXsbmGp9oIjG/Zc
VFnH0mFgJuwtnKid7jd/3tj5LZB1tmYwsHUvNhTzLr/uR/utVTkhv/x1iUg5t5A2
a9Jye/w2tKhnGezPgfNbHyj7YNq7i/1/Yw/Jwfi+enEr8Lzk3622Iz5JP37eWeXW
z7hSXqNTrxVMkVnYzQ9I0rSjxIcvogv9tLbKOIDOlGd3EUXpot+3m+aEZYChuucj
zvoSwDAxzgkCOAXJI3CyoeG4N2DNDhOm1FluAj4bzbInd7IDaasHpZ+oCh5Qi0rX
B4OF7tqw6XcL7J9iVsgsUG/69ygsvbcvhyhrj/LZ6uV2QBihDX4yujBYiJTdt9SA
oD7/ZfR0198zHqe+L6YYEXULQx5KlMCRkkLZIMUeRfylyEiq/3ktGnI+OibUDLsd
shAS1lFSq74TVyRjdWrhkUqSbgmVFzAplZmaajaIaDJXx3anA4cSq+kj35TOSHUx
6OxHgKlnqBUmOm3FWUjqAYhu3M52G2rSbJPKG8jhIz7D6wY2LfYddDk1YNYZ3Des
lLaD1G1Hbs6TxA0Kfx6qeoMNVXty4S3hWl4FALR+NkI7ppcckhzJ0GGiZnekE9So
US5Zsu0QSgdDn5JHl1U18yPo0JOEOQk+bW/uVcNonM1eSS7KMLrnd/V8KVWg1kT/
qC3dTSKOkTsG4GKwaUjqxxZK4kBKAZYKHfK7jrY8/zceJ+cy45jHco7FtIufLyeT
yyyMFR7Og4EaLNRJldXWrqAd5sh+H+H7sY9GYxgOZKJzzNU3yuISbmW/1Nl2vl63
CDXQKNrm0Ngaw8WpqgTLlILkPI7at40yK2i8gPkrcOv9CXfcOSpzqsYm34D2A7U8
3YhROIpNFkpti7cS49oDFYsxxYpeXWPAQzBiBT3O6sibmewKfNQf1Wlco6knvPH5
WXMM/lKw8ygik1cYRK/tMD46QOTzLLm9llvKDIxwoGQRPSklV+ZXYAiKDRBFCoDE
j0KnDEZHUW9bv+A3eVovvJO19cIhgL1+1WjrTOYqNXuYX7zd5vddf7zRXWOwU/gw
O0/eNEjsABR5q5qBPL/uOnNrxj+sNubBIe2d5/LqIhMCLi4p/g5OUoPhseR2a8WU
suf4gGbZ3b/h64+1dhAl7OJAFTWCJGHckFPGCfvyG+5Jvcj4YCQg8sQDsJjognei
5ZupUp8gMaaCSyOTpvWHmXpohnzQC6R5a1NnJU5ujC+t1N5YDaxiYvOx0giwR0hl
4sw0Zi1WIjSIg6cAwEVA0ut3YYDqrNKKTZk8NdCmWQqGfjsJPRqEqj0sRYGaiH3x
GAATxeoeLV4TJprqsEk9O1p5tQMluK+ShZ/cqlU2k8neygDSLtOQ+Ci/Fs3bXtoq
ZWkL8x+cCkhqAt4wXn7PUJ4Gfy9cBOYRjcMPAUpHUymItSEve2LghJhYdCgn+TUG
YLQ/xfm5hv48y35aN/DNX7jD/J5bb+CcCwv276V3sWGFixBwmmROUMN9yOFOJHxE
B09E6pbl+asamoL8+E6FHaHLVVr01dKolzCSaQ4XH5QlKlCaPVSlF+tc8AfGZliw
ml/mnlII4Vw/Nsa+UzOPu+4vvaxWaPhnep/6EiuofTbCGE1I6AU0e3KJ60m6ESM+
2/j4IZj2dcMPGaTOPgau3pUk+DrnRi06OgT1eqrhK2yYtlv7IZ0T4e8VdiDUnpT8
y67CjGsjOVrv4G8Qi0vnRl1gMu3+zXWe/75cET2g77vy/f9abjw4cy1uCi8eIck3
0AJEzYUn/IhxtI5LAoLsbJ4nNuz+ZkKyhuY4H4BP3ccK1nGYXtIEGNVzsTB2l4no
HgRPYaNnJALbjjUFLpmJjjts892YVEHI4qEMZvoxQOOBwqa1CEomrAmAFEWaLNgU
ev7cbXko4fV9KIKKTWXla5yfoqMRzks3AChFovOiE0+YujUYCRkU9ogvkI9tV578
oppWf018jcjA4wZa+bQODyXs/SxwWZnTVdGXhlMoLp2njz8h+BgDjn2PL4V9/rWt
qg6fy8SKlI7MGnCQc1GxQlGd6DtPUQSC75m/9JU6woHFCburbL18Hlj/ZI4ZB6f4
rJIr3t/1Fts2TXUUX8lZ8AbTVYB67J/mmNPJgMk0JIGxNy0CqH4ZCRV2DOB7yKYG
PJ7LRNwj86a3Pxo4nriM7liwk8LQke+2M+ArUYyRdo8rfNOerQX4uHRdXJEoimML
tf+aSWGVr+JMRKkM772aF45o9jKxuiPnLwFZy5xVF7gYlaU2D14wbvq7zshCu2ky
iF8G9rvI1C1t3ofWtPBEGhSkLzdx+8gBVygkCVvBJGnTs+kiO6jK5OtBCNQq8drZ
tpD/D+ozJSI0Oeh0VYwYGRR8iL8tIC2a5SEHpjbbtCzdS7ESOuHhXkeGOCmpTHWK
eP0v3Fu2MSVBniGJO6ls6vMM6VBCulvoQPsNnTKtPZXPdc8OH07No0Jfc1k8NW76
ODEFwbkFp8emAABfsjUDehGvVRsut5nEaZ0yR31pwSz1YmnfoLUt3GUUWSen15L3
g7djTCiPc3plwykmd2IS3xO907jJkwVXzqxQxt0pyHfLd+KpVwkBFsmGBcVn1mLO
QWNjjUvJvCF2DKGKhND8X+Or+a4b3i7lG5e8EFyOryJdB9QZGutgmjPxYXStTQuW
VPb0usNCLeSby9UGjMl3yN9wUOb38s35ZE6hAF4tBK5XITzT1Ez7Z90UT4i9p0Cq
/TfmF8oxm6VbJrBvo4DILIdTuZsWoTXH1ndIgzxljA7i3zUVv/bQODc5fX52BFb+
u17Wjtrhvrq/a8VsSr7v9u0+pfWk8qUgAP6PEilogiE2oddDHKBl33pxeQTRG+Ax
N8zEFjs9Th2DsT2vYSaqURcipdkPS0dWq5F9X+c90CYIEP4FSfXlsqs1OP5IUroj
TJyUwidH8FlplfAbZ5Xw3JhaoP18XIuqRtN2C7P3Eryx/CuK4VwNa3jcYpSG8+9j
U2vOBRYFVf8Nyq+aex/YgkBLb7L1hmTpjsjW/vcP6vJtLFdrB+oN+3qN7Qed2kNk
0X2OPGe1Stmwp8u6G/MQsqdEw/PV0wXsWwJFmZD4S9r+3oaJtE18utjMq4UUPACb
Ocmo/NYxhbgtysGc+daWP2u9yEVtcAHOFjsll5QW3asQrVzOSFcF7u8eMBuO9v7K
akeE/BPE9owimseWSiJn7Mn9doYZatvqfX+gTCui7vhxy9jo1CX0ebXO71kQvnqP
+yIEogMon357AkTvMy3VGMRz1nnE/G0GKaeWw0LdLEQVmSChcqP9gsnByGuYe/fE
jkaKeReALW/9ohTdbIXyJqHhiSL47vAUo77IuFdMhfmi5td4KoEPPqCJbRnqveGY
dNW4wKhlEu/BPrukrae74bbe2hOyuFeLuNsnyIzqMxfB1emw1BpXgYLU6SMpr5qO
QW+JzSsWnXDDvTTVInDi1SstZoeZwGcTos5drJJrHZwTT9VtSIa5GEYecrU3LxGb
2fplPn+7DIcp9O5lJTlWw5TvetWQtCCM1D4nVEOpJKveJE+sdUaON1oxpL1uiv+o
MJIUyXYo9w1mS6omlpnYzRRpv9iCMLNI03gg2cQNoy7ENzu3muXyzDMUtIUe/GBG
kED1jJ8vxqV590+RcZDbP0slig9UjwZ9IkIuc5xzVtEX+v4PRnPwjTCEL1PvFh/E
kiftxXUgsAbD8nFRt4KjA6uyLwqf1Pt2YQKL0/oNDQ/dt5QqN/yerpL0rpfUZ6NE
Tn2fpREtVT2rpTAcW4bWdf+KGdOkNI1ZHb4hTO66G/airylWTCJCsUgafH7hlCax
mMxCev0ucDEL5X47/OAZa4uQ5bqMBiElY8HruQghKECsgxMu+bHwFY71WvkCtVMo
0TAgPPpPeYDoOilkM5aETeH6rIN0dE5ZSjdB0/jxKC1ZkMXa1AWHeocFpVNFPZQz
5Fzpqpk3sn3HmbIGMNBAmSVkgChSy3pZVN1vkEIEly77rKoxPuisv54GSQm1JAMw
1h+drZbE7UyyLTU33g4CpPPvKUBaMKW2i58IsWkXZ6zxlq6HYFyKkpQIwhAR8BPx
xScEqOD4xNqNxREUON/qXj+OrsHOrHxqtV19RWiKfNZLDfjdbPMcHl+uKE3pmBUi
SbUBO3qUpWWTcjtP5zx2lhtNCE2EMAgh7QcFaz2oqseMARS3A8+oZ/SYjwrq74MF
1IbZpblo0puqcG74kwKGhEPaTP/1yK5gTA/FZWGEoSTAN7TCVtU3/L/8b6D5mew2
J1CHS+vzZL5rSPmdJ55mw6ZmyjYBI+M/Vnnu6/FHbBxZkXolCqxSX1eK2ppg6q5k
qr844E9tVeiQZ3LRgYFHBBhaW6zmdY0piYy+Akg5NUyGqaQAnBOTvA5HFVCGUoDR
Ht+PPN6LocDsDd0wqmudgSXCy5gUVRqGlObgpETEznAZS6B+GB5CK8xq0IRI643F
Dt0hwH9GK2j5drmSeBQ01ekmcgFhrUpA0/zFczaIp3LE71/6ZU4p+WOxg60u1xE/
1GwMdJt1pg8VncIMnUUhRi/qPgqkV02ZNYuUdDd6Nl4sKY0lZTpJYLWvM7ltmdZU
0GD7D/R3cKt2g2GYTcz57siItYrgZHowmJ+oDepsHCqOrODysXJNpGqzIRrzeOv9
S8DRoU6wzYygW5rU6XQb8J0DgTEcEkHSfccBEhD6hCoNLAfy1x+Y08zwRzL9zbnn
ov+9W+XVbRHtbYmARoJG/a7KuVENQ3By0/GSNvKWjl09ULYu26Qjj/06fL8MT4DO
theF0/0BdvmUHsJ6mRwkg2stBO75byc4XvCK524VPR4PwAVHm1R59KC9SlfdMsYP
QgjL+fRvKweq5NKgvG32lJEv3JtaFvGbip5C4FwqwNjHQ0pnaOwsSAC6XvIxEeu6
L9QPpEV4shzIrZjFGVYpeDxg2MBrAgwvfpNvzIT+GDpWeu1QpxsSTI1Yc4TbOVUp
MDPHBGGFYSsyOpws8w87TAXjTQZ4gpWeentTGWDtd9R/T4lWcwP/h79kqtFl26H6
1OIUese73ihjrixSp7H/dp8NtOI0uFyKtC52UTZQFsZWlIKu7KiMlIU4KVCv+BiV
VjGiKJ/TC2C12qSZHckyOfGA8jXvkhwV+YO1n52M3Q9n9axuMrBqfJZOdnKP1rx0
O52Y2e3Ns8VA+C+euqwKQ9enwKpQpWhVrL80haMxoH5gI41aY+UBgdYPMBqrPzXH
9WUJcnQFfkM3YHgFU2A39okPyobT1cSYeTN9EUE5yiYRxjyRaEOF3XZ4GcKM11F6
7k2wwgmXnQn6vxJr9pDz9vi0NVT+UIkfuci7PZW7T6BezlcEmNvLnKqvjZf29IYg
WFRGqxmHdqxRVGdKW9PLnNtiBYA3jcVubnAw9bjFd0QbDhWsFZSXu1tXMfqUJaHs
uwHmdhkrFSkbnlo+Dz6Ls0qLf+i90fm6WPyaw2QXGjV8HjThowGC99MudZ7tJSUM
6f1LakSoj9rkLWu3/7jEYrfreV8O2Co/7dqLWd0oGEdmN4o6hIpbcpUIbMg/u/JF
rsALBDK5tBkmXsL+ZaVgDHCqLCLeeaUbrv+B6CeW41sWQ7XDq+JgdriMfoanbh3n
BiPPioCRx/qmrYAoa8qHPBIPUH5q/OlbXFk77bSo+KMde8Tn+a8tAwcisDo+LbOm
Ah00/XNwepI7bVyInvIWEU7qCqbUrluo8VJAphTfsb6nHjgS/lJSlCATnd1lhHP9
PLZZXUDL51xJ+3jYMwB2M5WExISXK5dOo5o0Y0vDD8ETe4c73tU6oCcnSgmFbTcS
KrQKUT5WmOkSVGBaW8o5fzay5sT5N7TfVzyuoVDwy5Q1z6K/P+/zGvwj2doqiRbU
cypsXP4jPSGDBxnFvnhY/aDmCDN4e1NLjZ+uMFA0ck5ek6ohdX8clvwbai02Bm/S
YJ920mUNFRJzNu39hBIR0w2jgu/YUa93P47r2zQ760zzswZUtvc+sUIM7PO4DQ76
Zi5CWm3N9qVmKmr/zrNPMrz8gtkFM4whaZy8MbQvniBHF9LG25SvF+aWXC3OQPpZ
yVimyBK4PSiSoKMysSEqSRdi+J7SA9srtjONBU11J5DNTQ8+5kxJETuxP9NrVJH3
pYgB6aJf0Nnd6VDpf6+EqOtGr9M9GSfcN/GByxsLYlE9HuyOLWqKvIjgaHdKpuhR
dOt5cCl9zoqWmg8oJSjyQ3bnd6vDNDP6Romei3upLYpRY31+tk63fVTcSmpZoRgL
uj90iXU2gJaWqfpvDXzIzwurEv1ZlAXMAAI5iMw9Ote++Vb98OvpDoOFzHP7mExc
Q/ZRbyajb26dhKpxHZop5IgJiW/Ui6W8f10RybIhQ+DzRusuCh8QyO7DjN0TU3gs
qINftU+6DUBFFc8zQSQcKYAX1LSXe7XY0NtaHYgGcJrh4iRS7XUqwqzWQqFP8kyF
MUgXlC8oBf9AEfXdNVsBYGtsRBq22a6ZvuxZuHH4IDVppmBwY8QOR+JEme0lbJCg
SqrtcL7WvJq4J3n5DwS79tnMAXB1bcIdeRAo+M/RTEaxvpVJBDCH9qbja0prXTFP
cByBDts89IeOPDvrj86gd2X/+GHY1MG5aqtQJ3z05YqWM7+UQk+FaJpzHgI5xE2t
w5+/nX0YMZQiWrIHlIy8y9zR75KnJA9xy+vTlqTt5rV44zNT5g31mgxTcVisxdz7
bgIJZP35obWv9u2m1GiugPTDmjkmk+zjr24/KLk1NxGaDsEHwAdoabqYws6hFVk3
st2xox+lKGiKnjde/8P+wwno4EBTVc02KejmloRceTn17pIWNaPkwzSsH1DDsOo6
HCDzNco/74wInNH/OxWVuZA2DcWJ8lUeV6pAu6jX5K0cE0JC4mtqZ9eZPXqrNV+1
IXUUCMVnQZd9Y/uMpsu51Kt15bBqAVRLtU+Vzs/ZPUKvkcjPSAt4AiC7ZoCqdzF7
3Y6nXZGC5jSYEAiqcp0XwEpFoeNU9vYFRDWusqrb2HzT7RQxEuhZ0t8etv0Fi7Pu
Kn3f35Csr8iO9lPTov52R182gRr/gDKhecam3vdX8iXLLPJOduoLOhnROFTmriPx
CLOVnw5TTjPB6HZecIoNPNEbwdLLYwC/5S3vjddOKGaY4Cqol/mbsj7frhafR6tk
+53JoDuyUX1n9yrj266Jn/vACMM+ALY4b6euUGsBx7XgHX6o8+DYfXH7xO5uqRV/
gyTpZONtxW/2e8pn4VccYun+VefeKA+ismYpAPxTbTIwN3JYR3rLzbum0dYpgiW3
OnYZuvp2+IIL+wjjNMH4Pi5XxBX+oKi/RutYqKseoYoqxvSiRZG+O8d9GTgeSLfv
E1FqBu5Xo+aXTj32kMZov1LWFT4iAmwDfPvd8sf9eZeFSTi0tqFY4CavklTgJteu
s976gT+u5QWS2WJI1cIB4YgEX0U1E1tHl7cmoyGd07npThTgj+5c9uUZgwabvcnN
dJHBQkTrALX/2QFTuGfks1CPgUJWZ5RdjVuTlH6QLN8ACzmNh/OGcl//94nzChb8
ROI06IFdWFRreNM7E1hSNxLTBBN+Ucn9y3tp1cuyEuskTZP524I9fiqVgrqPSzIi
x+plVwVZBe9qHb7M2WJUJFuxBQCowBv4I3Re1JcXe/UuJMkz3I8Z3cSYr7fZYt44
fz43AouC44viRSW/zaMPWpMQsyvv6fFrTHHHQ8JCL6pi294TLy5I0nSruWzupsEQ
4kiWc/XTIoiGz2v1wCxcB6aayaj2xp8ldarUDWbeL+Cm5J+ttGErfd3lstb4NAoO
sCrf2sZr/Cr/VJm3ZRJVLX4xEn3kjaoeVKZfahZD5qM1u5juncZUCCAVLjvcbUZb
LwIN322/jcZoCXoVXKr2ARm/1juLD3trGTO+6vwJGYos5pfWu9wiXOyAI0PiYrmn
`pragma protect end_protected        
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
kAji1chAANL7ybQxu5Ph4rRZz5pKrH5BfyimVGHhs8p6Mv64SUuJ7halIMc5vUYm
AAc1epHsVTnNsK70TBIgQ+KyDr7xIBwAc2V/kajwXkqebeXujhAoytIR+75k/5yK
CPf0nXxcKecZzhdd03DdvP+MtMTAtKkzz5k7+DWJfxQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 269687    )
ND5FYYrioQ3kzMb7GdOL4y9do51J7TsZL3oX9nEj1QaCmm8kqq50NruvHGbamYpG
u3b0n3Qe/rQl4fYMEFU7if8qvBW2SfhEIkMb8Qq5d6H/kfuHgjzbOr7Mh6WW7Y2X
y/O3DvFP94kACi9e37IJSoCd7KZn2+NH7QEs/yE8oEXNK8pWcoRryjmUyNIVObx3
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Iq41b6QVJdZiFdLB2jZoJAFalO/M8DrBwFywtRh1IUlWA9IcC1dAcj0L5V2ut64B
JIGz1LWazdMZJrRYm2XUSjuTj31fpIyNMrVRUELsJkou1RsCoCKAsBAIZPsMSV/D
0vwM6luWZXdbUamIP/+BihYhHa42OtzuxYPcDusY/54=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 277579    )
kedpwBxfiOZ5y+qy1alw80ZgarcFuGfLymVYjX+DQI6mX8G9IafDs+CF+D6zdNZb
EbTXlUQGMCgREu8fzimc9uJIN1K6rFKFe4FoN5nZDpGjvJsJSmbmAsl3i1xStEwv
LZMHQe80Sm44oal1X9HrnlfftgQ/9p7j9c0T4tne+ZhgTcbyhC5FRJDqDRMbWfMn
5MpwU76rBrZWknyd9wvLVjxr1+qub4GOvuB4pGVrSkKL4QNvL8o/0NhjpKT12FxI
B+CUdveVpR6vMGRA9LhY/K+4Fz1XmCzAuAFOPhlKZbnsRQnKxMvtAhQf27+N1VNl
Bcsp4OuQSvbWBYCBU1l4ENeOt8IspA5Obke7fme5gKQkJgArlARtZgpAoDBayWCR
gwMtXJDsWioGz5sCHxmErus4ximth2Xy/GW8wLQvYM9mvG7Uz97xD97x0Na6xIle
WeK7I+s8mM2P6xbwId5jQMbZFB5mbp1ItEZ5n7C9ZBEg8hcHoCVG71pfdYa8Yh5f
AbJKkUgH0A8XH7G2LBHfkGO/ZBwr/Wt1bOrTGavAgEXGgDZHAJg7pwV8KFUEBxvW
tANoHZjuCLza1EY3gHM2VTRPqUlqaBHL1CB+N/xiizxgqlpfvBQdB0j8KSGeJOrD
4t+iGG9utZKL0smNt5eeyq1CQnIU88F92sHnzdDIswq1c+A3JPR+mArotUUNH1rB
YwIt6eK7+bAHgH/IeQ0ij4P4CuoNzCbajL0zkzTqHDG+cg6pVO19Jxt/TXNYY8SW
F2p/rZ6cEPAYipeoyKGz++J7/3xE0K7NZI20jKOKhlv4vBUBf73jEdIdDjDhPwEr
dzgoGpxfx5tbtJvYhQcfOPOtzy7RErVm/AGlGAftB73qRtg9W/3bXnay6toTYbwA
EcXedTrBJAdpUP2/KB1x03/+FveSGgteN59AV6j6rS3zQeIqgHU7zjpXDPcRwaUw
WO2ovBDoFaauKvhFBuABVDqVc3ZMj5oLpcEbf5SDhLSAoc1576TTxpyRgdq0JqP0
k0DxjjpDRb4x7i53fwFgVkQ9MsIiVVlI6cvck97Dj2WgS2sUHbifF3ZrkmshBRqk
wjNguExGWWsYETvz7T77u/FjNldfM9QgSuYRtnNILTNSgqLC5fUG8mmLBRX6yEbV
JOcKnj6C8AtfoQV7II3qwHcTePKVbQqb05M77awntgVPDcvGQRwopWdKbkSJYlBy
SZLg0cFXF/KPvMkpjj0hH5RehNhl+jdMSkjMX/+WXudCZW3kZNeRJKbpxrWVNHLl
SdiEfhz3nPxW8YyvyAT5rCpgvLXVzQ/1X0Xq3pxxbimhV+I4rn7Kg0T4/uSkmYcP
ypbEG0Us5nvfxVYk8Z79LkiWBeOW2XO9Zq79NLG//E22bWHrYAQ3+UyWGedD+mLo
cyHtjGlcXSpEABTGQtiIWnwMAR9NHC/xp6FSUVHPQNiRNhERnjwKytgjc/G/95mw
Ufl4Mxo6CkusDc0OmtRNvXcV7AtbsuiqB9cx/qbl8nYrgJHC0x3wueskT1xsvLLZ
MDQAe593iAg9birlnSGeserdayuq1t3IPLyX+0xysxkZKiCMk3KadGvdjvjzr8A0
3kWaLvGP+axqSPUz71GAKeqoXjBqNskuzrW1OffbLFf0Yq630AeywVRWpVEAL/xP
7QGWSvS71EIDecvvXX20MZ7N/OZ8DCMDxYjsmOu9UyRaSbeJ+hUF5dvKCmGHKcGT
Sts4pnYefPSTaIIZCxIxxH5KZR3PbQ/Ob7VDXzMNmbmSabqkbla9lzd1Q/hfDc1I
JYmlF5F85M/7KMYCgml6h4yabzdetjM9XM9ZFUh9wD2Aw1Uan6XBzpySTpN04lK3
+MMyLAM8Q2Gprdi35j0XI8BmPqsa8v4PEpzp3ddZ/ykmnExUTtoWAHDUkHbh4+R9
5FTptILNbMuApL9W0XDnEd3gKZqHESRGcaNqt+2/j752Ua7xTi3k0q7xrgm/XpZg
/G7ZhOIHbhzaXqKSCKurWxl4bxnwRL18dctZzhe8tmGeycAlLSosaOdIcoaZXcLC
nkdAyQgRE/NloN6Sj/tO7ufEBB+xXMIv1wh26fylBxLQCTds2OSMb/a79UiL1t+d
zkQ28f4y3lJgIHvE5Ke2MSGNIjM1j+/ZPCqy9ZQccnfAXMhg/91Km+FkFEcOACsQ
DLhJFaADLpvQUtcKgnGvrwdhc+qo3LJ2iM4uq/2e8y3fGbfESCXDvdtUMfirFoyk
Vnoud8UtUgDPGhwod8+C3eElEBd90290t3smk1L/+ptbb/c0y7Px9+XLAF9343+k
+KWLiIjki28jtUykQiV7H3u/awHm8zyTq+maWEoxPe1+x6/Zs5oA6tVAIBN3SR5s
vsMlj1aruN9LVqVKhUTcP5BLdOCLA88k6CoMtRgARajDgJiyQuEMcUfqsQ4nXZ54
mR8mNHAbe0Y54bnDSc2QR8xTeqN0lAB1Q/hPHeShiOhZm4oVgH1+gHPUBAL+kARj
l2Qo+MO9JB+y5QVR86/sDuu6pRQwcZVoOC2CIt5EyLZPyG4xHWm8BAYdqeCtqVI4
0/NmXLMzn+SqKHaFn/b5sjiubtErY5ci3RJ4Thm2AUI50PYLzSnZBb3hUqIzQXIc
1lVEQlkOCuchoh1hKugBPnbazKAEr4/KuO/ryQQ7r6Bnu+f+RhPwrykhsW+9H1Xk
JswrMPYWnq8XYQTbEURjnMoKjcmhs3JpyoZvZS64eteLQskCeLeCo+RU/pigtABQ
VRGqQs33XGzvekMznZbkZhGLykjI6oIrcisleIlWz+Jo/G3CSaAT9ExuTz3m1qwY
h2JmI8mWBYsuBWW1O26b5/Qa+f9SPWFEwJVdY2dybw7S3iniVlWHETyLB8lhCLmp
aSFLSIA1/X8gO0XQd4ZmoCjWb2ohqTPfyJ9OoAjiYuOfts7dv2hpzusPhDMc+5+g
24RZ43Q6YmJ2QsGuSUbCqQ26Xzh0xMO9Pt2Iky4aj3QBSPhtCMLiyYmbLREXVHlx
kl0CpMO/GkJpXNiJqU5iO7KK1sxEiKm2zca8nzdUfF99s0ePVwPK3vLW8gfOJY4i
uNHoDBb/dA6qB/7KnIdA03WbBq1RRJLdnByDR+dTMaPF5ihkfZx6Ds3WuY6dTBE3
TDXIYZtBZfblyln1gkZuVij00WkwmwK673emRVQQ/+Pio7aFTqTUiMblJNbgihsz
JaTrFL1kx1pme2OsbZVg3fAxHf/ArGUhvfqIZcfv7IsjvAXhKHVnCndwWXG2uyBo
HJRhgMiXmr3bIRdWt8hkvsIz0Af19sg7OgRLyZuva407T2bLcsMTMzsgONiN+3jC
tr7k8wbSDHfyxZRt8mrL3CwGKhfvSkB+kWTfCkunkgyUf9zEWnAfWTxhLa1U/0VM
yaWKP2Oj9+Gj9Byex1RWsIig5ULFSMbInSBStrv59+WbiPGQwKdZLa5JfwX0buWA
fNcMS6kE6D7b9FXOqH2Pqy/yrdwwemICSfDw6eOtCCRm2Ts7w2dyhCXo4FbYhs5C
VHRSyF8qEJ6UaYmh2z0XtDQMwuMtSqAP4fce9Rjlc1uPZY4IG6+k+Udh8Sjx/aws
ISM7jXJijrW0XBEfbKqeYDHsDUT1grVKJhMYSco3FVmnCa/6Mp19XJZUtAzOGOZI
R7PTGvmQrpKsZ7oeDaQ6Fg/Kw4KX13iBs6h9m2iwf7rhGz15dpZNLtWdmAMMNm6I
5dQy1zSle71CmuAhWYcQ68/BZUolQOzmgkzI82x04sPCRbRDj1OzvvE0tsrpVYUs
Lo2sxrl8THvdamrXBsOIE5IovwocDKnbBcJ4R2qwc9qEHyTdMkhsTdUXxOyodss2
i96ENvrBlA2MYY8BpbDysXgvmeCBDxWWA8Ab2rk+mKf5x5cRDsiFdso1U01A4Ku9
wYH2uYgEtDaRUXwCecrO4DlqDKsrnFUCpKvdk3qloA1UtqLvsmnMGWB0CFRLb2CH
JlW1//S3xkDGJTilIlEHeGvr+kJTv7ueSPnE0DM6xgJ6rgn0oiR/YEg5fDDFeAfx
3mABLfiVKM7zkm7jM+G4KwincY+UwlWrNSJ4gUP1Cm90TVWMZkmdO9BXh18EhrEc
Cz6W58qEQuSpNmQpPXO6z59Vt/qcWBhc5NkS2hBVRYaF49befelHSQnnHzCKvXRQ
GFsLypXUGIT6GPlJqrKPNSy1i/7JVXCdTi9lIXjbGkqoGJib28Q2NfGhDaSh6M64
MMdcdsMTXvaNJgQkrzdjuZzgee9+xvvD9HQZnP/YCFXRysrZg66sVMV0xyWdDmKb
qg/Rh2vI5sg34ymE0VkvoSjZGoDzMQW6L2wfjwBK0z/q+fkkTOyV6puq7ib73CL4
jYOXIbvH9E07K90dyniVrPo6UfJ5fg8LXzPiBFolv80FeJRqVOtRusThzCPrjVaC
+V3Ztz8dwentBGafaiLQWd2oRmICmkzGVo72IwKSokUiyoWfXQJArukgYuSWhfhs
wlz1tUCSFW4CLdqhlIC4Kl6GmONXyJALM6vxZQuzQN7OQsh5pLYRu1Kz1UDYCmId
Igh6q1LMejtmBaXDEFKkI1qjwdb1sCbxaNEa3G5HcafmpSYFY0e6c9Maq1anXJA+
JgSl9IfO5Yj6rGZBXlHfSX6kcROsWd9YWITHnNaQAS/R3UWJvZ9LHxje0Bh8YGjK
f5kzzGdQjCLwcBKYLVXP3ouokJxYCgXolzQ7qeAOsOPcxJjxFKtlKpr4tzvv/x7s
Za7/ZScl1cWl2G3p165sEAL/6IVXEhXOsd+1W3sQphDq+Ub/L+Gtsaxf7s34yz7X
wY4hlYcWB7uF9Uz7xcsblS1g5Ynm7InAGljwpfNgN5LltXD7Q99fT85jzjG/ICwA
w7QmC+bY0jW/rDb06wOtEUQNReUyzWSIkKgsC3gagmGJ8DqztMdKa5uYVULJcsos
dIp3zMxH6rAYD+efD+54/XTNrCbgxyRRH7i0LWiR6hmOb2ZmvXw6a9VoCYy+brWD
DkxqESzmSYiWHqbE+TiSmQibTgUiAp4TxmKhF8kAvAcuEWvYNkV+an+lxSQJikLI
BkgSk7/kPBOwmaC6jrRgvadvRNohVHKQ79ANV7jhOt2wWug9uxd+H6rWkszbpl+N
obszWKDhz2lFJ5Ly5twBTxFVK5VSJQ6enAGhAiRTUdCNiDAGdm7tf5qaX8zk3XVQ
3Uc5OwjNWAdSBF5Ghj8KvVFvsNnF0TLyjceu3fq5DrNxEQFMAIm0VThya7JUK6as
6kWxwyHRk/AeBp6ZsnVUkUiGLdBYYQ8S1gi9xI8+Wt7o7o38wu/HNujekiBbGD3B
yF2aRDisn6kfp2PIpEQ2H1gp4rUl3nGqeVX7nVamcLfcArkKdey03vouzPVtmXmI
gCqFIfiatYcEGjMKAri5yGEadtRHmVf8sY9S9MGnWhvdADhJF3ttYhPxjDD+/n98
RwAmqx2ILvN1k9razOk/cpOyb8a5MU89STUkAi6b+2rSOM2V5rn7L3wvKr9Ud7lB
KyhA9v8vnY4JO5atcN9dTTwlXzWEdbRGM5g764tg63M9ejWk4lMn/4Q9JB6r6RiD
A5nNtaxAplHQwLkaABgxMmEokX4ea2JqXePYtB3SfFKfSdKQv7SDOM7JUvWpRbE8
tns3T0SZjtgsG5PIsZ7AjRDvHLD/5izL3mfchFMnECBzru0YEEE2zmv7ETn2VXVi
heHYt8KBYCyzOqkiRZUp0v9gCQfOV9Jfh5CwapfUpSD4FTL27X/dHIz2PYqjZu87
9X99N0/BD4lQPaQvohgWly7JyLjV2LpPGZMKViVY5h4MAYW1js3bN8yQTZguzGk7
QZ40dR1+9KPu++zGijifLfqXUUIMK9fvZbhY1cOKzFhRH/vTdEyaqUYXU3yOzSmo
0wj6qqQYKchG9CPXci6/ByUTFbdQljqEG0z0F/6QL0oeyCuQYuvEXgfuYUrohXeg
Dc8Ccp4Ru7FaZoacuEA6sT1sScX/u9VJGth/oTULJiAVIFUlvnFbdgjj2QVGB1mF
l0ibDQ9Jc0reyPN7g6/bYZ52z+Zg8ClGe7ihu+VLZ3U7IAStikjf5TfR/sXiQu8c
Z3+Nk9GWvbbdirI140+ksuZm40Ey6QiWs76+0AzsPhPSiJAzbsA7y6sfpyeaJPEK
VVWeY0fzRXDNfBkfZA1r6ilvEZsx2ogXtfqDl76foh4LbYkkp+EMAA0hSfT0ljqi
MCmzcCLZ2ooQL1G305wQaxk5uQmPK3u4RBCFNuFdSG3y3Pl/MF1ElJQPbGoGi8Re
XrnLq1r5bUKqBZyQhGcUtHoKvvMoyZIDlkaMYcS2Gm4tqinOM00NSHvxD5CBrK+X
05Xykx0MEXrLIkYNOWthrxAinPwzuv88RCJ4OMynlndALmpfo1PV+jIVaBb/QTWx
VFaEGWYp344FgRNpJDFxKzf9qI1xV3uUY4bC62JkCf5igDUCWEL3yUBrX4JJiIXs
ND5z6Mg+sXkWoCog2hr+AYfQf9r9yexIm616oamMRXyucKBjP+i8S+8DydZwdL8h
AsQf05RCNrmGPy53XIQGN81Fpf57HOh7DG0Jh9C/U+lCMSdR83QJ1Dz05PB1hdi3
B2YIOnfaYTFa9/ikrAXHDSQjAkgZMhjnpSwUCgjXfiSpAI+nc5eCU1gHHmg6e7D3
dCL4a5Yg5dmGPcTF2+uOtZFy4qlRKdhys+2+Hy0EPKygpzObJeNQA+TlXpqotKI+
cwKF134WFYBIbihVcddXHVbbp7zz1C6Doifqq48LEDVF4tj8Td53CVIyJSGQRcLz
h84NNN3y4SWkgKMu0492UD1WgevU4/NqiexArrd8kcp0uOP0cwyIq6j/RzcnkauS
RaahZN3plidQb+3s4dR+Zob1Rlxui/86iXWAV5BlpSpbtLU7CRt5eXv/QCeDKCEK
vAijzmr8tv970xEZamghGWayR2AVRiS7rR08eSekWtwnIyelBXFJr4SbvZkPcdIX
EgzPjtWTBrstFE91s3oGfyxD7H/WF2vV91Oh6OqVRQD17ZUwEyhpDh7nZvUlo4gr
gF6C8rjD0ZRyJhVNd8VfuIgmdZMIWfeBRBNEOGo2anQauX5LY824NKWvxu9LIAfm
vPMzALF3wZqOoZpXjh2Mbs1eGNPV1OZ1FTUvhX5k+qThhd1rudLhuI+b68S2Ai/6
CPyNiBQFOgpTdaODGz57iZk2HlxTFyJ7gvj45CXjwcCz7nn1LaR95rFQ1GY6pRzU
/0s7Q2FjxuRjQN1HOErjJNbInXyu+ib1xab72WEkFRz3Jew/9KY2Pqqr9C+DjB0m
dM631Tzwa2N70ZVuR/RtZSIwECc4UNBZmFEnv0c0gxHPgT6Me+VVT6MmwUYIlVDL
LhEJLUD+8h2GC4f9hpD0AA4bxF+jRsm3FsgLMhhVN92GNVBLDaS1Hs37NDd1G/Bq
E/oNTJF8EHldIfsdSFZb0X+EqDm6JRmRPLO4DqbqcUhGoH87O4bKmR4JJ4FVsDCj
NG1SlrJd7ZSx12sxE9CkQUiJo1Q4x5Qvvd+r/jcGesbgUKTf7a6j4f0EF+dTXEqo
nIRcHkbiwX7fJKtNms40DU2D2oPdT47djGc8pXw2dneTE3Zq/tnqOj+jga7SG44A
s+BIfWqBLnJjI2RBBTCCghDwar+92pIb2j8NqqM2C/c0Rg204/Bse9AmqzpAIxCz
T0TlJGtuFADi1CYp6EqiOTBQ83s37aCAP0XzMVBlWbycSwLHlc4zAidyLK7wL38N
MPp8wUUF2aqlLq4o7qKYkBNvoAFO05fZK+M0ZAo67lU2v2vo1pCZO5KpKbZE4vng
0HPPktVqoFLfGFEfRgbigmMv/iTxZbUSXFwXtQ21URW72x5V6nrIPWU7S1q0N3Vc
4Lhpgghhscb/bggm3QHzpYZe2LeDOpZcEI92XhS4BZvYvXLqWoUcTjx7d3pwY9Sv
FSonGhqtienILIyveMS/M+gH25eH3Ol4OVR0XJzN4LGk+uLSnDiIqSNqF5EaN8/h
uH19H+/Dk2EEi4U6dA4tmKVoksC8ANGOHhN/MHQVdBQio6YeldzIzxYqmmQo7RKR
tLuvnA4Dn75mrEkG9E49JVucdKnsCWvk854kF1Zzsvnm15AeWUZEbvhgkZ4QMqHM
MSa1wcCb8Vhzt2EKA87jdNCvnKpGozsgehu4LSEK/dkeUokkNWKj/mqbvWIjUpJR
jllawgOJX2n7Cstyhz+kO/Xg6ZdJKJCxoYYiYB6YOSRIxwgKcYorD12SXz+q7nAm
lP9Qgn7zR36g+z5cnabkYS6/2CeXOtaK+dDbCaHHGNsS7MRX6c8kfp1G65WMQ7Ch
tDtR9JaLUGbLxC+SR9xmZH9HoIQe5qbiKdP9AU2BTnLyXQyEUf6yWIm9jWCHMoAh
hKkiAM6OFBrHNNHkqM97DR/w3v9PSAglv0pJYLTMaUv0MGZShlgYmEpu2dkdHBzM
0vPLigQuxCxIHzF/Dvo42BAeNc5hTSuuKoTnIW362TqFzFtaTSlIxxZSCTl1dlgQ
UAVy7pTGhGBcPfsLvtyXHeoMFYNOKs3zPBZakgBKTQvunRtmtph3qDZUiJhQCd5h
fKnmyFEqunRwhODzDVh+MZA2OvrmaC4VomBuxT0ESRG1oLg+Mn8vvTbbDp0u+8+J
zui+C3b5cKksHexI7OGP5MLXDgmz+aWjlcdo0MeJOIyyQdqfWvbprMhrPeYXmRJX
8x0laqVZjPuTrqTroS0z8AA8uVcoqzllk/fOtfMuOYf4BBFlw8WwykYfJ9Tp2JyT
MtHdjEJacLQTLs+67i70O+K1odDOsiW5QJhDNtLJTVwT0s+hOa3DYKyf8ZYpoAWA
42sP0X26lNXOC3zOyOSI6lGXj5SU3GggicuzDLUlpbwR09usQjHFzmPT5qRbf8Ic
Aqd4J6Xz7tn/bbWrCJF1oNqSXtXzVQKSFYGqPWBiCuZ+OCBjqa2X3BqD2AmvMLZm
5NaPMmvedyhxEV6I5dSrjE9JO8sGnWJajWAO1NN+j82aIrsRlqmQYb6iH+rlixQH
OeCjob9y2CMbTxpiu1XjoKok3wVckw7cVTHB9xIDiCCq669iHqDdHd0R1MPpYKTL
scVTLTwqXeR5Mi3FyQLI6TdmSeutvODfV7kSCHC6zFpyGslypKeM1y+P77Z8yCNG
3hcHL8/uWCYoHa11Upvq16N4JCRtKdpOBU8TVCTg9WLWqZBfWz1T+xCVmNsy8aE/
h+WYXVwtxzKEhJwX8JH10NhavdP2CLlowZgYK56K43P6+tAw4tkf/lPkW0g/8LBr
UjBMbjNWjXZMB9SG+Qa/nM7+kegrZPSA1HOMrq3IP5HuBGHjPnz5pCFtpwcprKEq
LF3dop7h6NeNmGeGLkr1iDaO4PllbV1CwFljxadyRQBGj2Oc+u3UQBNbY+oz6Cx5
umD+0bTgPXkYxiDR/KQO/CTtVcjaW4vQ5BPDikWiRiBhEie7ZLixJKu/5QM1BK7f
eIU6KKPhtXadnZTczQwNLCOzG9UeGxBqh9UaUV+cJsqnYcjt5dlhXzFH5yN6lJA0
Yo9pQvoXMhRsUQ1gndE+tQHUr+COC1N9dDLsUFbNMP5Ns3MZI+kddTWQJzET+p/l
XQe5oTKS1GGjlQexHPASDB6eKX+rsxJY/rGqmWsZFE9lPY9bgremM97rliqd9zQT
qR8d3w+e8CvIu+MYj6qzEumyamLDF9C/xkoTDm3T53vH1yLqKwMhP8KUI3jrcLyy
SsXoaTjbYK3LTkfJz+YFsEGDOFRKB7L/CS/dqxW1weOD7PSlVflB2owLQn06Y0/G
N3fyPrVXoKxU7RbrvV5ZAhtTT3KWTFnAWuGfwHb1/+YWCeQzPkX1A7TI3jOyGKGO
9SOa1CbM0C3vWyisvHexbGv3wyHcEqw4SyHW6Pn7v2lNboankDzoczljGgogsuOL
JXunnWlQT5T5vzY9LIZQ6/ArIftlJFLl5hP8iE7XuarHmG59GYrij+y/KmtGPPbz
3bjj4vP8v2dxYf4jZAOeUy84QbBZWtb1xasx9llvUIvNJ6B4GEjzbZXeX45VMBtG
Yskg2UC+7igrfTQ9DD/gS1Mvb7fXtKp5K6WHfXKvUbJS49YULjqwplj6ON+ZWAXG
6xt3enjV3Df7mPcHrQ6T4rhiu4wZL1OV26lavCDgvGGGFdZJcGjLNILIk+39x28X
gCNaCu6HoqOVMySAbi6DJkR6lR/kve0r4mbQN474oHTFLbZVICuBpDVPH3s5Xz3K
pEy8QgytKiSHZv1CI3odSX3nZrR+tOzLs9+c4It2R9cg05xJccZ9vaNCJk+VWf2o
VG8zQBZ8Z/11GgM6n4lfsLjvYX0xeKRG2le8jEZ0kWvghu8xczCI4yUe9JCjU+3m
lwFlv5soglxFKDWCejqovL5FgXKv5v8p1+SlbEgeOAAe+hKWwJtlluEx5zRmTukx
/6vdiHmDFkTHut/sw1RGOvGBhp1IRAXhE623MpAT783F/DtRkn9xuRNMIUdW0PUr
1iOmjNNHkxEVhiDgtYlbUcprSueRj0pqd9/AILd7N9w=
`pragma protect end_protected        
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
VTTwMWL1do9qBeFbeNnd2Ekb20MovVAunwdor/T8JE1KRHOMQSMCrevE2UaR1m8I
H05txGhMdicwFA5264rtjRQgLB8BXYvbZSdjdlT91aZ8ysYb5jzQIvT55q4lAsQo
0XzKHWqTXnq0rGz5XveymerNfayjWRODwAMaENxwf9s=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 277924    )
aTcNi2TFTzzuI4M9KGx1XoyNf0/ftoBXu3KXELZp6wY7cIpdHDkBJhb1lW2Mzrcm
EC9UsoahQsEVuhwjAPYiNExEc9AUvKYg9G4PAMdk31HNRRG63mfxVxE7nOncC1/b
TRSaxydrQzpXC5jBlHZ7/bD9JEfpynP7VcipcYGwFzudUk9hQNDpk2DlLvRn03EG
xxKiDWjVUWSC3kEhpPElVepNzaY5jbEhNBzN8EUVpefzzeRqDF6EKnCo3AZdVhj9
uKuHiSXT5usvr7KqgY2bl72YFUFDwNhygqSiP5T6K/BwVK9QGYwIYsKapRhteiUe
p2Vyt6NPW9YkPTGiuVhJRDg0zZ4KOkdlPlQ4MyJWdDFAVhhWVLH7nZRon7WZ3sBK
iR06O5MGKQppzZNvuddFX17LV4FcjnfD2J9VMFe003dAaUQOIS4oLf3i1gxlzCgM
fAJMjMoSdoWMwip/k/FRIA==
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
G2hiH4fRsIl9eFIsOKylKvyjgeCU3g58F68po5n3WcfY7iHYcLuJkOWRpYSH2RJe
GkOuMhKJf27xFRmA/dNuSYyi2nPbpVhIZ6aoQO/e9TbW5fYLZjwwXvKZ6DQAaJF8
JxPxa1WqGornHlZ6U3MZlpxcIo5UzeARLXAdTyieeZE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 289117    )
stKrGqTkPWMl0aQruedQxzduETqEQ2ClOShy7EaUPC2kzs36b+4BZ5e2x+qD8w8n
Pk3Fsyx2k9s2o+3ZWOJLPm1oosduS7/fINt4NOkjOJmoDu0+r30seTeVfrc8lFOx
YFnKanFw8Xz/rrSj1ArkqbhIfZHnUSqax0GHzjhHjWQ/8YTWEmk0Bfi9zmwEPmr8
e1pLFIdhoxLoK3MOithQ4o7xo1OLCFrUJaMz85dz7PZhm+tc4Yk90UxF5vRQQGuW
IcUCVgTOhr8nhKw16BfF/TmAxnrmq0ZCwv6NK+L3DXz/sJ9NKS6bVm0p3y+QHDJC
8PdMS1lhDKDH5lH8hnhTIDAVvno79KyTJGlDuXpJ33BbCZfqSfGLv7UU4w5zQUO3
AUdskMdTBGzh5XkB+SGheDPyTzuKqQXTs8Qp8X40/6ZHD3tp8TWWKjmA8pp/jdVg
1BJHnfZ8pFxlTINHFuJNVebJiN6J/8tdlXQg2WntGb5HyPChxm6bY4xXtXcXReF/
zH0p6ioWxqjZck7yvHFr5UgFBW4Tjrla2s4b6I6+3d7grSnW2pa4/2RYIPtoyeC1
w7GXNUlqXr+nYMtp+vsBK+SdtgyOpzraJXWSMnV2c4O5fFLVwdDNtN2KDmxlON62
gPM7jO+KaK03r4pZF7Lw2TDRe+C8zlSfUZvUzSRuEecT8/Aze9czindTDArcI6BR
oGeggLlBSV9+j5k1iGEzqHPqMfVhuhf9LvA0G5O20h7QLTJjArm4XQQ8CRyDyfEf
5QFSZ6QbqE9kjv/xvxGLLsp7PBrfHhCxR6xhDi7jwsRD5RJQtXVhG/vfK+csH3no
j3oGroQQN30SkctwYvxczeoWwoM4mDNm6VKEaKVy/IxDc/6jIFFsLkJZU8i9D27Z
e9BQveFKfDc62d/RJtM5NSckyEqJs5D+MqclP8+SPo+b0gXlI7Ra0HCdNAas84Jz
utVokeKQxpljfbGywTpTQKbN6/RdsJya3TPooc52HebKZKg0qUleZB6o0KLGOn/c
JR6PVP5CxmkBmB+DOcQJSwBfRdo3VyyZOBuookRot0YFsNd66ziCIeYVHyQhJ+mc
518q46wl71/jPVQG6WVdGNGq05snq7YH/TOpgc/LG9LZ1m/hT1Jl5kwLnA5yIoR9
0L2bT+j+lL4j8Z/9xPjj6e2CXfUvTIYOvO4Oxdvfzrx0MiWTt0dsrC5TVNxkRLkL
kvGUu3pzpMWMryDjj21TuKRbGHhCrDGbHIhxW0jy09XHX5swD5YIVTRhBYjqowyB
mFf9c1m4jq2tYE0aphJG5i7ISnYPW3CvlJzcrtU1HWTUaaX1/+VejtsFrAtEbjyS
haccJs9GiUKQ9XPWFwV4Hwlu1Neyf/rn7TbESK8ranJ0T8ZqH3Z00VdQvtWUMjM2
l8MNWDPd2OVwhfkp57OzPC63uDoiGURCYYoCpnoS6xDS4Srt7YLsdFVadvLdlF0x
0EOyBqbeoVTdwCnQ/yTlBq0m0vMsgGcQL9Legr1166sdR5HW/ENjKXdwo3IcmunM
4B+281B4qs3VOthfI9GI2eCEsc23GzaSNiOeyoYDcmA/R6nInUVujq7wTKgkQHBK
ha5ZA8ccK+xcIeM063ZzOWO/Lmidjg/FmBNJEOV7is0oTgEpuysa1UVU/fbIOyMK
ZaK5zipJ0DWdj6FZ159/lROvB7c55C01vdWU8Rr5HHazuqSL58sNWdRoYQ0tBIDg
nVpxH8N2WF4anwzc1ShMBDdw8Ppf+oT3CuJx33vcORgShjKP16KCHrQr3JDEcUqD
eOwvahCi5/fEaGdrZz4u9+qb4RlJgbxS28Ri6OMnqaVzaBwgriAFbk5HaU+YmZO4
txZFtjlyliZL8bhKlv7nFOh23LvGhjhiGF39ipqgiVeyE39LamORuuokLsUOTuB2
KUkntnZvuqbz+8Ao/IhOOlhvPg2sdaqYamyFcDb0AlHg9g4Z4UUWKu+Qtb9hE7Lc
ccZGXDyikHIA/XOrihdJhwqQWKyDh06SKFCIG2xHcLkV7ZQsbiy9u9o8ltfgm4T5
55aibbvTQ3WTmZ10r0YmwWoLrgyRZnAfC0yoQ3BjX/XVQbNUc/W1z/T21RuP8IDB
CaGY5j9SoHyrw5nviq1uDGu4+JpDI2FrA/ITlLgt686j/Bnhz9qxWYwvBJ2sJWZR
sfs3asr+mKzghQw5dmFzkU8MP9eDrb0ubM19gBRk/zCK2SBOr+NLRDtfJ+yAmxwn
7B5BkIjwYjCASCLgC0MyNIRvnENPtjFToq13F9+0DIzOWBsfmUCPAPPGQUfnNNAV
eUoTcASnSL14SACxHmu5U56GSTTJ9uW47kpz3TUoqoCo3LlFE6QKy8YPY4X8J2cr
R2m58a+hcmiqHNBTUeU7eLFrDhuCnhCwmQ6cPv03RqN+bDLF6mJXTukj7AQnF6no
8v3oIJB2y9bHkNLNH8yfw5JKiVaZYN09gxhRr1Rn1CStUVpNFDUHha5MYOAA8J3z
jo3WX3jZsTr5tW0P8v1uF6KRYPEDpBKv1RTek4JAOOBqGd7JT/NNGOy9+lW+y7On
GbOmyAxM1oY8FlrJLbcp5xrQsuSkNUPlwMHzhFMHrFn6ghzanGccYqj4DiuJNKs3
Wd3TT0R8jR6A2dRJeCCBWnyHUHbqKOgGk7cfgbIRR/xPfUxWlf2BztrwL7ZABg8X
lhwIXonXhMM/CO7ykITeIGtT42qSbbba6A6vco8nrQto64DUP8VKApN1rdgEHxrU
zQqLfRkdVZK4DiZa21GnWX+fwNZTBtJMvN43RP8ELmjgqhPRFmuiWBi7C5AcO0qH
bYnkAJh8ZoAj2ap/H8Tt/S45b/b2aK7VVzccYx9N6aomw+DDcY+at/dG54GfCe00
C3ihhBIbxo9N9obkpIZKmGzLz+u18VzeaYFO54AeizBt+eEwiFSIL8NdTCVcdFoA
4Ai+se35pWGvHcgWI+f/+TSO+uINWDouV8uexs7c4phDtnNTe510hM/ObGhKyu3E
AIdHG+2E4ogZEVNMPxLFfxvVMd/9AE1XgnargKp/gF+YXBbwIyFoB14WRBGtv6GD
sI2YdPhzt0A21ffhMNdqEvgXov18QRaegkdvDmIeb9/TulLc3pAuN0fnjgiG+blT
ZVWNQZa3A6M+/N/MYWpAQflysHwpXsI1GdGjrc07eWnqQBezYOa1dq0N69/EECUP
ftl9+iA48aj9tP6gFRSOgXSDTA+Ntf3eh2zo1L0bhXmOx0DHOmDo22q65r6lDQUS
KdXLBeUmEud8quDpdcW/nVmGAz0HiSThqK+K5suCZqT/e7l1tYqknIG4CO+mvdaO
nGO72a/u0XdeBr8TwgjA92zouFp3+qdnavLSotbe0ljyJBpCwe6CHMHL3E0Dn6BV
P7jueIMe9bIWg5fPdepOOQ9/6il8KjsJTI+5u2HWpuaBDTEoXnrk011Xy0lFsRdU
stHKcBiNWQub0SpeRtwtYCUsuNBgKGH2csorP7tEkC6UouAeLkvKJ/rPWKcJi3xy
PGBbg2watHk9IGh/v5hahDRXMdnVxDXsLT0hytTip2pg9ZeRMNStYgt4GRdrA6Qv
V6xhzKLFpI1LrS5lM4mQvbya8nGRUFsk3S8k3IQuSaB1dglJ84Xv912eIr7IWtUp
VvGA0fIW06bARSzFfo60T+gOuyY8viiCZ59vuDW4UymrZg4CZcjGuh7Jpe03cDL8
tVBCAFHHfGWLLIxgOaHT5Cr79dHaLwdT6Hx7CQQqOsTBSQHEzgZflbklK2Wud4Og
d8eRPYyxK2eUwknw8vOJN7mQv2jL/q0mYaWT3Wka9i/hikrWc3uG/kDwXsu0LeGn
hM8N4z0sHJpUFITZ3pQdZ2iq+TXQj1fBe0XUC4caSpl7/XcMS7bhtyrLGvbOlMfe
WjVNhN+C7DbOswIl/HUDGhX31r7cyPVpQrJNlPfjuBJAitFvABm8M/qjibEQza/T
c2Kz+45hf/sQMX3CmGbBX02btMGzmTuAySGChiQ7/lZoDBQjm0UKZZYwgASJjIe6
daQ3IQqEnfZFlq5qcI2FsUjlavN+sLz77Yv83K9OyNTN1+CTC99CrwojOBtkujmd
6TiGYQzL//SyD3/PUe90Rn957wtDpu5ie5GJ8Y68SymfXzcAPpWJgmKh0VUPKx+n
s++NZty3dJedlvio+XT8Ghlb4DCRTAnIL0l0zzFodCj1NKg7+BXwm6+wPY/LoRTk
FxceHMNQLLP2ogcid4dDIf6/xar/2cuq+ws5ByXPme4HOH0JPwYsxcyPSQi8M46g
eZjlosRmkY0202bHq5KJEIjoKFBENDQ+vsgrFiwTmxUEzuwwsKNNsBK0C8IPwxhn
fhZFv2IZcochGqTo25MZFq8qahBVUqF8PecwLniK29NlHTw1zfJzQsZD4vzMQV1l
82HJHtsrTJJy/VKgJEEBhQtVY/Ka78y43GdD6N/iQL8cAVQD41Y8lV4I14JpTVsN
d5DQ4TAoacxQxnuFCsPPkxSgDFY2iTu6sIw65Zh3qbOYOFb3PEs3AZmY8upa3N4n
VcRw/DUv2uMG0gWnJfv6VLrKC3QdwScn+4kLbqYVTN6sEy4MwpJzAMbICjbLipjB
7IxUhPmByDLJ3O6rdkp4IJ4goZIpkaLows6qdv62vid6og80omSOonb067h0HuYM
ipBTOCmwkAyo5RErl/IeZnspfN04KHnEyuqKqQ4P4Z1KgLeMnHRxJvoRvtJGWKG/
c/UhBznFaBuYENItVmAl2XlU5qXrdZbf347iYRwE4zSxuoBbOzR2PsEGanRvUZ28
nVaW8x+HBbXrgNZtNnHPzCWfR5M1aeYN9vDGgUmmy6iUIzaf0LJqXj3Qiqm9QDa6
esbGT4szgTpQJ08WbN8ol4ODHz0/OGUkaqel3XrVXQFfGcVk9B8WlepLovyA7q4u
azbMwTuNO0r2ujaMDf3ePZ8H+9TgavcB56iSDNiHNtbb/VCGTl88/Y1xQAcvCtVS
122eoG9vXwkQrtRHxBwu9YWDMRSsNyaDoyrkvum9n6Pi9Wd5rsqhCdC/fallxikk
gbf/ZTBTs6R/uJZxvs4zaAqqVnSVQUTgklgwhyBiq4kCs2kIyIl2JOtiyHulP8Ts
C0/TmV9vvSORVMxopyTCDsYgtDodKbGxkDfeUltRbP5eGpB5gx7gh7fL15Y+PhXu
Mc4JaYLmHvLJSjL3koRjpgO01IbNLa2XYc/lcfuMeG+/WSuVSYQr1zBkZG35UNel
GHw7EfEZM0XnIOWpe7pVfr/D/pfz1Rbc+YGQ3d2/hNHFYC4umDQmy/aIublA+igP
KBSbgIp+hd0ZzZRp/MwNJIVehB9YAWEetc3AvFIUvhobR+mFIgM9bKVoY+B1z3Qz
wzNd1bxebPlTktB23FDO1byfSt0tHUySBa8PkngYF67UKLmsvG4kuWJaqWYFMUdn
T1JNDS2XjAgRDyr0G1vGmAd+1N/boZw9FHqyEU11yW00pAM+b3rm4TGRArR/yM1p
GcV+0kQXlk+Ew7FBp7gJTr9HtCAQOCLO92qPwFsTX+q91lBESzB8EvZcK0iRAfDo
Lfw3yZpQNTvmK6Phe+WNtv9IFApxfb2Jkx8HjoZWyu4q1/eI6NZWsJa+5IEwMInH
8JD58DUMoiCZA/s+a3m/9l5bxzvjHuQgGACK5lpdeGzceb1xDBMu4njPM5+vwA1I
1WbcAAtyZblwtJI2tAcmoS5QfoXFuaAmjDNNBmwJf8IS32g5wuBJfHKkSds5ZIIG
4EgciGO1XbbE5kRzoGt9sLVybGBNiSlnyFRjEY9sEFsj3sDkWvfW0Axc3RI84OYa
VTeVMDJ4/X95b170wfyaa68Sw35y/caWvaDxwNxwttJKm9FSiQpT9naLxG+qvHAS
VvQoHX6V6kJjj143qVa/EpIs0axJDyarQ0IcQXIZaL7yW/TWFrVUWxzkwUlhO6Y5
rm9/yk8jnCktNBJTde577ZZri3exKhIjx7b0+k0YvFak6rBUEwSTR3tafvX0Y17d
n4TR/LmDs2dRbHXL19hA8OA6RVXRC9mvfP6pIwD1yizceh0ohusNILw0xFYC5d+e
48uvHLsli3IFmctmcqkulZQohUnTZVy4kOGsNg2JolFrnYb8ErjAiI+o3y+qJORa
NFVm9OKOiklk6rHfhBKYeCgRattKpGBlKIz/+IzgxAa/u9pHHnVzijZXfqw3eIha
HtA9UrkdKwiYrxpaqCoKaAzZYNRlZ+9TL7QTiGe1eeuhtsRYaBtC0z5rN2ntISjm
DeUCi7VGOM1MPir9BDZkyVoULm86vH2UnajtFfiNas3BRdioWfS2Ua0HR741YLqs
9qAuZGw3wyIcOKjeGYmUso+z/XABnFlLOe6cE7eEpt1g9l6piN6cmNF5G0Jnbhmf
Gq2q4H1UFEdapn7SWZOD7fOGkZrWJk1SpfspUHpDCE1UVr+bTClgUeufdGElcJbe
JRcKghltlbeymGqU3IyUYgPzG2GGyKIdl//vyykBp4XY9hyytg2IGzUNqJRw6MQv
1sxuVmzy4MdUxgjxSS39iGbT8ui9jERdp4IYXttS3SVGK8+AXM0XeV4iT/jazSyd
xPugKrBBR5QV6ogfoy2SjSQ+P43boZxIqYBpuUrUlw2XT3x8yVLLUR89kMi1zxlu
ggsdIL+eRWQKfaVpRbpM1o97DX+ILM01heKfQ+iYwezBLQWG7905GnEVFuzSN1h+
e6zGcCsfLwwOKBYzL0dStNc/1Iq3VcNEUXKmCHiyQcXfDnNbdHkfcMMyBy7EqlQV
r2tzWmOx6oA0L06isrFKoYiSLfi2Bu/SwwKA7w5dw1XrisJSzeO0Ojg2HIEgftXb
IlusxZjzOYP/N8tzsPJmvmuWIhVLHvkIw9ylOmd6PA3gDYTRTm1kctx/JLmRpx+Q
Hs4Yhw46uGqwPmijE+e1xK69grNvYz3d0TebvauK9Z9iEPY3maOE2LfUx7eX6WM1
cKlcG2+aO7RhugeRrc1rBFovs2z5AYRH5avp5n0OE1Jifqdy6U9NwjTdIcHVzp2n
zOzAzczulm7hCaEoiTmXFLqN7btdRm0HbTuTT/jtXb6BMhbCIV5gvkgj0OLT8Xfd
3YDUzLIPjFZK4eETRa0rZoOFGFdio8Ts70VdXVLYB1XrZPM8BEtH87Xpddt+JTbM
0o11hh0TZR+NAPW3qgrK2+LKjHX1dZp3qrV9fGfh1ll3I6IpDh1mMcKU17CelfLd
ZLhQdyxehNq8g+Czmbxmw/fgh7K8pqSi50DiElBaJAOEVyAnU13Uw+wQOH2AbjcG
/a/ElK8Bdl3jgWL9ChXnTh5jKqvjnbrUlGNf4BRiZNN+xLbOQYIhy5TIuaUhylr7
l7lG2zckUifBtjKUNmLYZGBJbywag/riZDQdKiLydNLanQNXmJ1cpiA61nyaoDe9
QrdFcrAuuRfi1EdBBrKE8avk29YuZjeHy/91fk5vBlMd1rYCqxyum3G7uFs0okAO
pBCzmuKZKEj/tGNuo59d414C+KqMsxpCtln1DAJa5bV1HEN/QoXxEZb1h25SXJiK
OJsIjmIUjgCWH7+B5bGZflZk3V1aniW3tskeZ3BAqodBDH1HJf59p5e6qSP4vD+c
4MNiqR2ovsXzHU1UFqlT38xa7Co0GKb3FQJj2RdoqeI5h/6Xv+bXJlhsO/ahCGe0
hghnGo+fL95qm5+UWwleryNpZQzUM4v/Q1ffcAVn1lXYKkagslg9PT/QN3TnlywC
dOTaSDeuB3D8wzQwuIVAx+M7DpBYF7ME7FKnGtN+R5GssakAQ6TJuvd/9D3exFOU
HbEoR2i6MoQWrnVuKtOlAPCAeaw+b20vQD5m8hUPth7ykM0eqmsvcsADRlscmENc
W283aqLofIVoxYdehAWETg2COackDtP9K7QDT+GrjGJUyuYAmY3Abn+gQjJCp0ia
YYkozEEkc43k01fsWlVltNkVTHhxelJyzRnrg/YnC2aTOwSVUljaz25SG/lJxLwB
H1bnggNDj8ebmQRe2SkGM2ovumkjDTzja16yl3BxB0/0pk2DxWUiqO1O/3DOefCc
Xtbq4Z/9JRdeSR6Jhi8mp8sk8BRnkSBSL2NtkTVvTZXYqnzrHcXTgzJiCKdPDg4W
O4iMpKm3JPYLS9wPcGNiWU6BtcuJuc9M3NzyEFxcQ5A+7lGRZ9sityunrR/aaTLy
SNeO5jymqH1jsS5j/dh0c8nfpUxTkdjuo8hQJEv1l7kvc7tiU8PnxIQ73eyRK0mF
bVXx0jjJTRY5AAaxeaNdTbncmO9z9NWZ+FtSUBF/9cyHnLUms7LyAES/RPDBLpIz
LBcSOflZlgqUe0xspKVSDS377aUYFvdFqNWUhGFmgWFknjuAyXd3GcZK5T32wGR8
B0wjeLGpigKfGpZXE0pr0WGdOKpJgDjRd5g3UERHEtpIgbxsHsKW077yzaWgwevS
2s4skFi8DtzSx2p9whvUH+acXSFQIJnLdHeEh0XaTQRj4uWfydGyrPg42ANTrfm4
f0OrL07EyojeAeC2p2l/TE34VCxvVx5zOnz9fitArIrajyQb5//41DCJgRySp1uT
6P8CHMKUb0X2GI9DOgjo/rS8D4TwXHlTadXjAKzsACWA/pEYvy6lmviZUCqjwKHc
uBOspBeKKTFWv9KbM8aQ1ZdnXlSGkPtJdp4deN4cn1BSuTu/NESBDIrHaC085W6y
7Gopcsiclx4TpilRrGQR4mPO3xhUlrQddFeFmTo6vRY1LQoLiQGl635P95gYiUB3
MZUQHVjUtmSIsoOGAxk3J4Dpcd72bJLzd4xg+r3WuGnsczac9bR7YdJtANsdSjJf
KRFGuAX7Acgc2CwaB2lFJhm9ENl55B+b7nHSjEGqqgugL3poFfwtEMX5zXYjoF3r
M4Pz10cqNtZpNiJZB0Uvu0SzWadOKWiUYXkKI/4l1ishstWySzkLBxCCzs/3S4hb
d9EHCCuIiaVk8ZoKyp9xTXiB7gzyWbLtnP5TMZyVqI3csoe84jnVdwwTtGJPgqtu
TiCe5NXdFl07t1KNBP2tVe4hMBmWi8zKPmYH/l00HsKDFJ3/TX5cmREd9nR3MZQg
W+flC+CbbWh5piodlN4J1yhz12HHafobHdRj4u5i+aPyxUkfkaASre1QNveee6hR
1EjxP+B0XdUaDLcZibeh/ut0+IAgLyg0laUITsaMD4R7RBIPU2EOW8eXZHPwsXSX
6B2S8feCj6+xK/5lPptjLwz6ozdYMjHx2InFhbRKboZgw7NIRhZANmVgb66cr6fJ
zpSunrSFJAauWZMOrsHCNa0W46WNzbWSoTYYhxk+hi4iKwFHbb2e6S0JQ9cepZf0
nsSWdRCfz+pPiHWuOWlBZbTIwv6ur55vJ9ZkPoVtK/2rpWF0CyfH4qWWKT+avD6f
i/eyR5DqLma4laCrEI7iiuK69OOJmX4IIsVKB1lAt7x0eZZTQkHYvSeq4XuIKQlc
ZS2uxMbx9U3Stoy0qtppX6O24ShZ4N5R/bCaoUICbdT2wWOVVQNFA7+VAaYbsJ+S
uXvmbq7YTydhAn22Vqm6f7nmYp1Lo88wo50yYiYK7Ucd7bjfhtFGUynDCf19dGQC
f43ij9bf7CeDfDR3AalaJnXjnkX6O84xKSGgav5KScs/I6Y4y16eLWYcWiQ9QNkm
TwDhwE+sLFM8d5xEqbv2ZQoqiziaJlHUfIyzgkVkl/pE+QUMiLCFmxcVatr2CtI5
f5pz5GEF5ZeE0Nguvd0Dt6VRBBKdXQRS2ItSE8lw82P+UrVlp7AvBoG5Rj1tZqnK
bLoa4vf12OpLPlmJRnQSMQtvLSguTSMSjJEVnG9ocoqhW47YiGCBZx6cJYX1SXSy
ESWHOyv6AAzg/obyCHVHQrMCtApedeArUHD5hhdIYgRybOLVz2mNn1fOKqDXZhsG
G39kqvqXzGh19zK3UiBxpRgRLVZ/XiR6tlxnocizwsFoq00rx/2HfT2vOGp72HRe
1dPrU0EGVwP5fObkd+ILHMH0ofhD/i+UPmmMJ0r7UqM3oLtRSjjNxcHhV2k9VcJL
OUr/wG5uKrGWASF8EbRGf4uEqw/1Z/vz66lXBG4G9Uz3Ddzk2TXtLlW2Ja3fNtQD
uGbfDa/pRknRabc4JNZwLytiA7lENsYymMdxI5/7bKjDEkANIX+hYREVEBa2ZB5U
J2fPO73mcRS5T6QEGXS3j79A+8h2IizQWYPKf3Ejv7MwSmbGmNaK/p+RZJ4E7Q/w
BrEzxLUMvTd05WPuUuG2FcGVnFGL3LF3ecptMv7wqyj2IZGD/LsIsdXAwlNHvCVM
JC1jLZBkbzwr8dNfcu8hrt+upGmHXKdNKOsSr6V57uIQJ2Sgi1tQMHb9EQwGa4cg
5LR07i+c4v5aygy1vOPRPidbXgcpGkXjybaDrud10nJYjH2guCeWzcuXP9Y4rek6
9RYogyz5DuaZfBgZcig6TQ2yLPt3yfuSNJ37sGW6n26ktH3OGvUbeO2sAh9ObCEE
KWmlBLZOv9W/O1iFr3QAL0x7xMUjfCciGxRv7uDRMtbDylcN3P/rWuRCZPGrTjv3
zIpIxVqIyPK+ln1zrWnot2AxRWwfXENxNfPJcSB1xj4uJeJD7xPurfEya1GcndgA
+RnH6uepmyo/e3Gbl0JOfIu8S2r6ibWoNgL9FYAVp8GmIDN/DMBMNo9a0VrSJN0a
TiGaoi51dhgIlQ7TNnEqKuh9KYSinYuctqIltXtSZ03ii32EdzFbJqq3Y+ty3RJS
NE2INEO9RrtKWMfn23VJdpT/Mv5Nt6LFWCMmhDFHQOBF1o1WCs3wRP/dRcuYtsEB
RjOPbKTxu7Zfn7qxkBvVzbU7AWYTkP4gVHJwhHRH3kXae7P5zti23WqM9F+qY7U2
j3bOuTReRwcWbmeH1QvjQNyPc77WN2t7OWMJVLgzGRcPEvZ5Ydim2zpqYwF61tq6
IeFOawmju0j/ZgAuBzzZ2rFeW7bg1SaxIqCvJsOpGztwfNnyDTxcPRhJOXmPsaxL
am1k64+dR6FWvrDAr+71ZQ4t00bd2PTrm58Y2BGuwlhFGOFAVpL3ls/luWJswQ7+
RAL8eFdTr8Vg5UR8DpLtUwnCw6Z5QvKMw9DU2gRKyJ3RhNd5YrBBNYTdheyBFR2R
BspehfC3UWp2G3kYpcW8wu+2RWaq4gfzGncu37W6ZtW+caYcoc0pKKc+YLCdcz/g
Tnye4U7vL5L85VL5eMhX6Q59075zMvnjkQOyXkitp0/0S6Lv/dJx4GqyRyd6gk8B
lVoTd/dvDu8l9mosfsB19vm6T/yNKFvsf56aqvKQARt6omQNZB1khrEDLaNzaYzT
EkQCh1Y81dFZlDmIwntWMvClaqf8iSLeEAIsWizh2P5liw9WIJn/GnfyFbilQ6p/
Ro2WrSM8dGn7Kzidxzm6zd8onN/g9p69n3l4UR24VQa228Xqt16aUxfTa1sBUEUc
Y589HBnMrfLP7Qc8w5HIUDcD98nGuTCsp2t+VCSoLrDghkIW8lJRjBWdKqWZfVC3
ximgBQG2dLesGE2t2GIwhDCvZUjDNUoFGQNNDeSy0N4hq2Gp/7uJCr+NH877eMm8
tF9U2KlzK97yCOf3Hup2ty74Eb5JceuqKkb0EI/Ub0TdZExJIi+d5lCGWZulbWwJ
nFzDx18Sgl2bQZGOcnSoBTz3Ok6ZqJtkBS3uBg9bSphNP23DLQlnCHLeUoqNnYny
6NGYfsGXkHTAWL9jK/uZXBTcl45pp+hp+NDQgOFGAAytVOxB8LHQdgptxTPfCQIb
ypbhRfnwzRc5vJ2P8kfKqX36jFd/YuFDwR2w2FLH7GtCFKodCBVKLWEwhMb0GsAZ
FUjqOYddp0A4I/LDSbpefvuFbeMhvuFwkDEkZDORSSQWLLSjPydtRNUbA4vmeBLL
Sd6Xn4S0ZN7cSEAIchIjOrKo7ml+PP9ej8z3uBt67Df5Fzx/yExRfVO5Z6ehNHRN
tvp5pHJbNTPNYE+xivmAsxgDfwaSkhhEWBRVH0VZ3shcovi6jnrztUGyWRBeO7ug
4jr+h0GzEYd1XEwmdvAMVoWY+wDOUAhMQxOCJge5B8OnmU6HVNclC9OBHXCH88/l
ZBGJjSQTilVFtJDPqaR5GB9zlq0oiHe9P4fd+1w2sNAl4zwq1b3WSuiZs+uj30a9
jSgNzGE881aTWV9zhugM8q2t8LbGj7ou3xUwHWWDNBcxBq54pndymZ1UF1ePyy2b
Ci/czOhJbjtzJRpC4aTWWN6d0tOEBC0OIngW5fhL+RUeNWFVbB2FbbpDjmQ01hGF
8Z6oP+qObHEtWxSnEi2BTut7U2UcxNXF45VyeWjUWRLS1GDZ7ap1M0t1xcTfvatX
I/vx5fo3DIk/xigVobBJ1wERGrOwCDrCQiwuE5/8/nstxs22AhcqsB33Vti+HjK8
gypXeIinmZHY6TITX2tVvohbPFKEX2O6mchdPxtc2N5Vq9uXFgeBeETKgvd3iYYd
j0tgIwqtfFn5Uiy/EuEMDCPhnTMqoOAwRMduAm3+Dmki/lKWplhXV0CBZBW4nwtI
EB8zSoD25crkET9aRqo2w24PpEaJw5x5SmCmtOXqUFWDbXQSG7QtiPhzqU3gkknD
/gar/JcmZtYovG4yGYSCmTkK4VmRMncFNweYLHlHL73rth2oVnlmBSJp0oBOaLJl
y9XV4Sy/16d6IMsRSn6rmGxjUeCz1d/pQbvgBGRASEmrvQgX9wif9LoSQiRsYpVJ
YAdf6azRCdk5m1wIDelui/68mI6cGcVbkNp4od5dfWSMIPg0Yfh/MJKeM6HqbQGh
yNPYhgun39Nu6JHztJiRrCi3K5F/YkzL/AOmeP3h2qKqLwsAG/ySgHTuO2/7Zf0J
7m35LprhhHVW8+XUqYGqEY+yScI5mAdGfapjTjwX3qr1CoYAO3S65hr308WHEq2z
Ip4Zvbdg8b35UPGYmJz1RkqZm/DsuGMc+Xi8t64Y5XKiuGnKMk9VBUU5hAoXWYUy
gpkP8ck/Sx6TElpEu4gF3fym0LDBFXsE1Qwy0Hpnf+DuCLa4mHvKBB1N2/qqgwZV
B2Cwb+k3rVWnEo7WVoVvHHMM3Hjm7o3REw1yG+xu9IDLeRhqRfa9jLRrNnWUmfsF
ge+qWRaZSEu9PSjpkhB0Cu+phD4zq1FyN4LWKw+XauzAwI+u0gisHEcN2dXUS2kw
mfB7pPOXy2b5gu0QcrzvxkvdEIItp4dtmF3JbKD92D+VLurbGyWFsCdJKCRnwX2h
c+c7dT962/YNVsnmDqS6ATNk1IjETHBW6PILhBYAy2l6+Y8LqsRN/qwCceLh17Ww
RrNxJ5NnRQ45F0G4r4RgeD8AkwOeCt097w5TTngziq4XK8sbHevN7yJJEctxdVcE
23kd0eVLALgj+ShsrqcL0HG7t4M+N+ZfmQ2jdd+XZrk44/7P+vLAf9NkznF7M3mB
MZNPS9D0K8jqkkDd+b7x+g+rbwtZbZ70DYkIL73fxKSubzpie0b+J+YFSO7KIXj8
BUoRJj1OQjfe2pLWCRFMNKE+acTYaQBNNJ3c2VhVGHP7fJ4y26AanJWHWCzRPE4Z
JQ78oys+wP9yMC/jCy/qpirVupyFLaFn6GGc4/gykYwuQO2UdG61hgUtqqZ53d/U
5K9SQ4SQxxBMn67g7De5ERsAodhq/xVlSq3urVZKlIRI+k0gXOMzJQsLlc7LG4Kd
C4pjs5fi+RdmdornfO2P26c8hsI0gZw/wfd78/9BX2V5L3Z0jcNM05h61hoM4IEN
UArDAlZa9JJUmyYbHTLxm6gNu4xh06ViKSjK6brvx4DGrTkre6ihFFpHQOvIAjeD
OS9rgL0U2sY/4KWI67DBzN0RJ2GUANDaTapg9mGQGijoNrkSTy0zfC2gEBBHJd0a
2tqR2NH86CLVkM0IV6wcTnBrCZxhw9G+Bj4YzM5Pi8H6L1kiZVfXOk5+SIWwoeNT
BbaKJAYYL5Fs9387SqF+Q1r8BRbxH9O3GX07f6tsES5u2A3BK0tjLR3mlxGFzmTl
pEchrgM7haB3v8z6jAsekwiqIUZXvFwozd9ipuqB59NKgPI1s/eYfwARGQjNl6n6
fid1yXeblSUTc2ZGxzH1OuOUeugQcg859n+UsTlxE1A9DoFmj1piHQgJVSr248sQ
JjVq2WRkfin9gZ2RrDXZgTniQtsNmraNq7UjrPgdxIO5CTxZj92k8N0dWpzI4Ag1
BPGZ6wPWWKuc5lGf1jvcMAXm01GB1FJ5a+OKRnle30shNDqcAL8PlLgKRASkAZcN
+zCA+tWxAQsSB7p41Z2DqOwson1l60f5t65+KTQAzyaXS1ks/3bPMrmZ6h13ZyLE
D5hxhAk/0EY7HJCLdmAFE6bS8k6Asl7FOrx4qmr45omO3c0c4R1UqG5NUZlv/dcn
vMK+bwJVT5mwYDITDUu2mVomSFLBiHWJoUYAoVAl9TR5mKrpyi8C/QVrZnkuo3nM
RDU2ub9Wgeis7yc+VWbBdvI2l4vvIps5JkUty3HwHj+APWDmlHFzj7ybYB7CfmcG
t4tZAtYAHl6Lia/Nb1nJKvGBgvz8XcHxhk3es4uy/Lk6C3B318XVw0fhViURagow
IeoNQnKSd4Zc1CyJ+nKrsYh8caaz+Tusctqqu1qIJz+qVaPjtAdBGCsNOFKHg6JQ
FChsU70P8acRRmAAYH5bP+ej8QNDaaG6zbmmTMGI1F7WXE29fZVaz/5GrkEv9RFX
D2gP69DGWhDE+3Qx6jn2NtpB2Q9WBYLzVpogOHq+XKRZDRN+sOVn4xqS1hNFedB9
2aN91KIJ/+b29cKtuFQaSbxpYBNveHlByMjpORmYyr4jRVFzz4clAjfcxG1vqvWD
rMcuyHdd6cO9p36lVaVMaIoM555YK8BAH3+6+uy3Qh+8NwPx3yGbBc9lGqiPKPiu
L5qwAm239+HXX8uZJi6B3Q==
`pragma protect end_protected      

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
PbON2WwUXFiIrx3lWjlDZDiTExj9pMKkGfvkN1oHr7cHrjUhNAtKG9vQDuSHXLnm
PbbA+/EXGNQxndyMxvKWvGxIhVnVpXhVvFoq1PfrrK9Dl7gRhpPKEI4VHy/MnWqz
2RUZC2WTguMC7HOWstSifG8HBSGageipFKlu7yn17J4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 289228    )
33iwUOoHDRY5RzBPFeeMPa0n3kUY29ct5klaoV2d578bjO5LcxBG6zW+k2ZrpnaE
7R3wZ026Mmc2talyLduhFe5BlfkdtXxChovK/p2fabhjV/szAuRW/bkjFo7C1yF3
y6PBByxiHEIgmd0Kbn9VnA==
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
dmX5xuFkGKEmAf49yzi60sZKmGmZx2ZeMG6cRYdnKHHHsCZMomSKopKgUinXeYE0
HIqZPD8Mkd+LVa7Y/GfRyd75mbriE70h/dG0MMCJZRWuKMAS/Wc9cZAucJfCmQJU
UeKl3KmlovE6tkQ2hQlqoCbkmr8/FVAYsAahEw4tp4k=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 294211    )
SqEHCo5YAn0gow4ELHsme3JveW42s/tcV1Tx959c1nlVBNjdzz2mKkifKnVxg50y
KW8sIJdj04LdKC6TQ8UsFNm+JhApBS017F9mjpea7xZ1+gAoX4sOjWhLaa/t/Kac
B9dJBW1R379LoWRDOiIgjfbS2bDG/eTVODwswA/wAO+q8XeSASztRMlca+Fcesx0
vUbSw1tjUnPkXYRCGxHuy8CsAAWZNTQw8pxFhWnL1dktkwArzXZ7Ia05xLa94kuF
Imq0lm66mlS9Q9+MwOn017FHOw4vmS2xUIH0dRCUk6RVMONY/x+dNMfOeWwq6TnA
gobfE6JHVzm6sp1wowK4i/Wk8ygnxBsEargAxjyLc264AvFtdtU4n4r+v0SxBag3
XgT1mmBs0e6YhnGTy9M7nAGdVUWp9l4+jfqkSW16uEbAVp3VAR9drAZ551o4tpzv
szmYdK3S8XMednKQYHhc0cOh7u9UvaLKLsQGDdZHe2V/7uf+GOBqCUhO6nAgOl9+
TIA/mVIBNAY2Vj7OxqvpUzEdE6A/JIK9Sr8w1p/RMrESoSISMV1hVNDJQMEPWah5
kaWSRrch/Ka1KrgNORSVnNh5oNADE9Q98JY4laBG1GkiHKq99O+QRnGd6EH5vP5B
gvBiCz5vXNvx8L6VZxSA7JzI8unUmp9ei3YrH/+J3bxJHAB+9v3VO2uvFPE3hg6k
HyQiL9dLzvTnK2aplCB/9AEc7/fNrvPp3VObmChrWhNo9xoTKYqpjuUBbhrJKa7v
Z1LIlQuT3sLCUyQG8X79zabtpnHDJ09ec4BeIHzFiRISoAuLs5GmF1/93GkQE8ne
TVh7LQujJXtpaiMUdZdNBuVdySdXyDZwyG+AW5ZFB8bupjBOnXxxoaryt7g9OvLr
vOKtLMiaGIHiw9jqveSaKtK/B4zRQwJGmtIV/b12qdkTp1kOHnh7Jvd7BN0Boesh
J1qMvGVvmd8kN4dbuY8f0f4R3nipwynet9URxdz+iOobi38/cdCuqs7ABvLq3LMR
K1FowObaGBlYUMMRKStzfKKAZnDi8of0w5Ev4fgCnNnAb+yf0Oz0489lEzLJn2Y4
rhQEBElHpTN4H4LizkHKHiX9QaIvmRkIqf+r0wUdIcrZBVudIMD1+XKw80CxTqq6
7Ex8vcZ2SLCDz9+xdVo4/hEiKxiSqY7TXB0i5x/rRWR7AseDFVRxEClCsP8IeYvY
YHOW7+0VwoYSXKVS+oGLhpBtnx61SjxNfYRsE95iLa6VgycR69IuSLrdBCKo2wLn
bjvfq4TfE7HLNR9nDyG80sMMITWC9Ji/Lrn9ig+81Z/4g/OTrQARgsL+8EeRSvqG
Az2IKElKxqPVtBmVXCkULCuF0UZtRsUuLNqYYuoJ0FtSJyNVrgzxkC4pyBiOW9RF
+qb1zlSsvNWWCwy7EH/LIyuF1gVdaMwdkaTN/qI2n7MtZTyL0REC6AtSUjiqduiC
GHz3EP15WjgsOIcV8l8cas84Ks5k7/deEbOtMwWUEBkCkSpBs2G4GpmmEO7q7F+j
UlSO77CoxjmrcFWAyvSlonz4hX0NaYnRjnbjyYeHi5G233mJlVekuzXLX83D2da+
pCw/Izd8eyTUUuQrD9QpbBjnojQkg2CbeiZF8TS2+ySdfe2WlGMoEMdAY5Ds/Cf8
/8vGLbVr38jGn+IH1myvuSuhRW4MepIYzZld2p4PIhP36J8XraqCMaB8I2Eour6l
wcoI/aLjxVD8VaAb/QdMgl3uMO1+kqFBgW3JOlvHu6U4Uk8xkdky4tuG1rn4dSqU
QCmcdyeYSmju4HCMYN7/uXpv8T/cZ/5lX6cjnKPs7n4utB0xWf98Rr8nQLzVhbeY
xNbyVrRK3lu3avCPpogI3DeZcfwazQQ4BWKDsbqY96Fx83oQFMplzdodFfIlf5rN
WmT1RfJkk2/qrtoL3M426Qq0Wob49IjcTH0WKWfdrmNiY4H7/7PZRHPaYcAWwLHC
lS1MKxcU4nsLYl20iVt3W6z/DVsxTUZTXhHAlPmwgmRDklERB/GayG6llQ9N/wWz
QlpO9Eh3k7D2Pf+Uqvntp7zPUM2eWwtgbImvKF3hbZshRpqRHALVTkqVEcW8JXMV
8CISZ9VRtux9VMpt8Q1bxhKV5JupSwAj9rIbR8ILM0S0vFu05PBlamtl2r3Qk721
TNbeqvBFZWMxnNitiimGMTUi0ZQsuQUBwlph7vL5OfFvdq4yWniugJXSE1nCfb22
bzqkvG1sORzEJWyoVEje3Yv0TRbDSH/UR+rsV1qRkdwhYl+USfwLsDw2+iCsJ6eT
a8owGoh3RMyZa2iWtTCU07t1pzvpM9dwP8diFUjUS4UynPd3Os7aMB2+COgwJ68D
BaEUtM5OokV5MknFpL/c6oMlKyXZ4izrCBhj6djIi7wHdVdSBc8yAfwaLfs/SBrQ
4DC0wnRP3zl+csifFnwe+zdjUvHssk4Oze2UhUpY4KV2Gm+LhH6tfI9Lrcx1nMER
AOUV82ddiMCN795711I6ibgaT5tReCo/mJdlUyGB+fk4ibeM0PjyaUrO99tyN/F1
JmXvT18jJSls6yCvWFZnRl7jtjUI6bjMC+MhTEBmJ4zSkkbbPT76U/X8IT81Ll1X
i6zLHA+SpYjiroEa6qsGIMpGZAJhZAzYsUOBBx/X83dkBZWlShfNcV7r80BndNsJ
181paZa+suWDXTJm014F8stZWIN85grmjGEJ89Rhed7bcq1CFZZio2TKISBARqpi
d+4Namki0chAm9pbvTlSSItDL9RYX6aYrBo0mES4B6Kw/wQxj5JMy2S3YOa2sMuF
vcFXy0Stp7KMGz+zJDVcM8zkWhl9MGoxQt9fb5iKpUNvqCZnY285n8BOKcizRju6
wEFMNh7vdxrDDTcfEkja5ZKl9F4Tt2GHBepG1/aV3SMfLLYifZH68viCTLXHrZV/
GNV3IQqsYUymBWj3+0RDB7vhPjEKOXe8dzpwg8gE70TsHfDNJCJd/Mguhw9Nc+Cs
tL81ohLP0fC8h9rPSEd3yZj/1j4H6Xv6jSDPHFMecIJI/E6HFHQrkY+Z6zbcg2nw
QEK98dTsqP7S7rE7n/oJu9e5kBqb+r7KfgtGX1UlAfHlQTvf2qmUILldaqRuYH9X
vXKjdZnGTfMkjFg0Y7zYr3KL9WEgkxl7XyqdhAA5/RJLcMUP7HcM1gcbxemxudQ6
LtZ2JVPB2x+6ZB4Dn1P13Cflf6HifRDra3nSXD4RoRfeSFW9zWlnfxM9k+FKTqNC
VWLJfcY+93R/Ml/8jmOFlJ16ApZIeA82oioUPIjCScGdYBtueco9ny/Wst1SOon0
vc9rEX6F2elB+NklfTvxHhRHHiNshtrzJZu0NlIDo3SBLVM4dATEARwCQf/DZ2sS
4PDHLucPnDP0xv0K2k6lmbU/rkZW7eT9J0zEeoWEnpbsLRhoUbZgsulLxCZD5+Ey
AVoNPeLBtgUn9uUgKSXjwR+xWBxBV+SmOMiSUwG0N7W/QyuuUFXYiJvhE3kqx743
MuZ+dIfStymFeKpqZV+pHoddsiEhQznT2nf/THuiFYBbDOD4e1g64ed+k4UQMfbI
zug9a0ZtZzccoPyUuwc6+vx3Mpy+KU9rbw4KC3C+N4TcEsnNdyoop8Wzz3PxiM3S
OlsD+hcoXAV7gLZtynI7Xx/NonDpVesR7DfLh1f/qJ6Y26NAkNQX/f2/08/v2CcW
7XQyXO5HTMIQVHSJOCWX9Ua7LPtj9vehf8R1aSOi3qxICrDgqD4+GqM2yvmuiGU7
jl2Eabx0ixQI2Rfwz2s5qLZrdkrZh7CXxMFdOirAhgvDoI9GwQyUgbHxLefso70e
fezwrIx66RuXbDaKJpY6UU+VBL2hEzsOc4HBfPx8mNtO0PV4XhmKxBg0Yim7umrK
1miprTGZbLtnkQlbObrNZm+FTNjd/KvrRAZjKO/n1m+oPMZkMJ0sHn7A1/p5MMzJ
2VzjnapQwsWK7QFimlHVLFzpV2i0Zyrf4/jTy1wgjD4K9bRADevHFIVn4NwNm0oS
LfVIwqmhhfvQ9KrwAp469RyXTBlUUyP2aLE+68+UguzPp0xXHINyvs0eOs/FQZoK
sbohcTMF4arMugk0f3oW0ahVj33CeuQ8gZmRR3Kk9M59q7tPBeg1bT2HrSKXYndj
Rn7xtGSyCOFApCqsm7CMvIBFuDtMbiTmd9cHQvlTkbzVMaLPJWxi2IJZQQfpJqIb
dquXRwdDshnnSAo/C2O2wgJ8uBQJXY3OMNW/qRfxbCTrO/TLKrDA2pTMg7tKcGHh
phC29w37ErJ0UV2ZrZluK8Bj9WID1Yjq53O9i8EUzLLnUYcoUFGzveCCmGeS5TEr
5Z9s6v8ghcCLzf94eGgsKM7wo02oVTWJdLAYzp8uLae6Tan29hq593s2ziG6r3J9
Hg9UAYkz00lAWijRRFTY71sg2g0pfnQoMV3HXxshQ2YRB1mTQZRX3LwE05WXAkvq
dE17I1cpvY6mTxThG6d6bVB0snvFl5ZhYfkigPBz3m576lTNsx+MycSvP6dU+NvY
YvvfuBam6++rgXVAMwsswzCibKhff87DWHrX7AJyKkLEKwrxblHCnKdtDlr5ydMy
dSoBufcGriksIJls8Fhq7Wj6TQFvME3fifEK/vFWnJSOLKfJ6/xtrWOVWPtJEMp8
sYIrDNQF42JEVzn0bMyN4kN449xdlO+XMfIyNtfAB2LP87tDPw2tMqejcFb5Wq6A
uLsS58VoYFgsPE7/0Pvx/eohx3q/+Dt9k0fkq16EUlLxmi327f5sEXhVJ1zIugpw
82rj1n8mhtTfLcrpf+KkVtUyUy0KYv0d2cFX05fbVnQIbxJ9CZ/EsNJj+6hkEYhB
SCw2m818NWG7gQo1imqIaHMWzWmWLQp0BiElP3/ArHNFjoym6lGrBNlfpAKkxtXW
+akATL2uuG3Qo/xhfbsMm51y8GJWe0L6U+XWb3h4eSAh0S6Dp51z5ctzoo8l9wmT
mq40vF2rj0IrDshtJglhye2D4QMLTAoMVpxqz/WpGgCr90zYYtr1UUy0uuIqfQ/B
QahNhKQ7GS6TBn0+SaVuUoRwt3ZcF/uWvw2FXvZVKa4ZdAOxBGmBWxy0hMpoxyxU
gazegjptAjIlwCNslpw3/KjfyvCSn408jcVmz5larDHDHwnVliCm48l+0PqMx2u3
s/BaZa29TuinmOptXa5uYd2e3qe4X/jASmLuotDHK74dOh7vX5k5Mq0CfaimUY54
F/dnzo4biMrnSX2cgOMQJVaKc7/ChDerktIFmOfTeMl9uIJYOp2SyQrCDS/9eVcU
9gllCJ/UW4oQB1zQlzhNZ7gsAlHdmMMX0GKdBZDOomIhN9DwOJqQNgTBK1Pw6mev
4TDmXTH0NNCGG8H2DP399HC7Ur0rLBbhHJFbM0Pk1lb/7XEKVsCmEitxEWDtnTlc
3BKtH91hcw+mx6BKq7z6vHfPIuLtSjpI614L09+b4CC3Wax0gs0N3V/YLgcOYQ5L
fNaTmdbQqu/c2TCbo9feVnfwrcOhXC3l0YGZjUfYxkDjr2zSKNw8Dhe5iujksKXH
TMwtOT548gbtgbtYykl1GF/fvt4EYLf3xYF9XYULQlvuN9TA8JADrAH5X6nvDpZ2
D0UExF0/Oc8XSWyviDm9+Bv+tDiMGqnJE+VT0WLitGNFsqHgHpsEM64FMa9Wk8mR
D8hXEhWEOgl4NinGL1KUkIvAIjP8g5GT2BQKdHoq1wpoy1osIfSQOuZnmwWx8ird
+4oqB3PejmSXvrd2TSCZL2+u6q3TvfoYR1zIdEXhSB8oJzdiejCMnb5pYB8W1Mlt
sgNPyZBVMMWMKpgB8smSFGWZEQNabMwWJHdzjZzrsFfI1SOdD1FDpKXDgE3q/OkF
dmsyji3Ac1h9FwkGuUOQMpjMo+4bbtL8lBwCAj+GNfeM9U4+Jz9hQvJAL/RP+hYF
91MlYZtp2D2wzwCBSEFmd1v2w4k/5GbXtyj/0EUqFcA7DPP2f9MVTw7a1RCmZblP
XXVr0UdT1tIjHa8Iele5k3bFPBR7MC/s0q6MaG/LANvE3DzrjMlrOTnDgRyEifu3
y6Hn0kS4qQYYiJ7LBipRt9+4J3xf5EWRz+u3g87Cy5F3XDupW+vH0SOgNu/R6TQQ
AAn9tZdMUQwg9MsmZuuCJpNQhHim5Krg5oQKqhnZkaNTVmN4/yC+7iOMqhqIDA3e
zFbAlwCg4pslsn7FXSFvn4B4K6XQhGZJDE75mMjpPxCkCtm6W3JrS62rX++qk1wX
cvi0SJxromqaWEW6C+iZpNFuDWRJWXHSP9CF/XtGrvlkgIcllUC8YE7EIduzUJJv
RN23WubbIduub3i8w8gfPu0Z6YXSKgmwb14WaqYk1Bh67cTHJEEq8zJBEDL9Hp+h
iPXDsuvevqVRh5vPLntkrz4shpkl0gk1jdx/3wlKicWtiOsi+Toepbd2HD43EBNK
vGOvzYg5yPUYAFuF9CyYSeSfMbYLQEpA25bz6gG3+oxSHTBwVXcHrMNKagogAw6u
GGD/iwLvZooG1HPW3KRb3frXW09YuU+emDwIFpSIGabxKkMJD3cBPAGOe8QTv0MX
9+SvSBQRfTBNE4duMZDgo/LxgpmsbAY46AEd2CLkbJfpOdKG8WlNidQYuCrd43uh
`pragma protect end_protected  
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
oq0UN1jpqC6iR7aiItjFsSS4k4moLNdqqjimocmEnBgLj9fEfZRo/vPYL4jmzik8
Isw5aemQ2/xFZdWTkM76OQOG6eoVzke12lpBlr7c18MVi2Dtnub8DqfUUtOU6OcS
PgpR56lxC5N3CMYVnCfpevtqRytInZyIixxy3Tp5S00=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 294350    )
W4/C758PAhhwV596KHGaBtzuCAf778KwltCwQuke9r9EUp/4zg+GHnHiumi7bTCz
5gdrethTht+k6wTa7gMQwaHGjbjAeFckuSGBLCtZlBvX5PakDHwvkAfueYp6yPJv
YBBxBQQGo/trsWrkXKtC//Lc5J7bkIcQSiFg8p7RFYJWmChU6xbd21bNI+8UaU0/
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
H0f2Oj+GkK9odU7HBOZvHfAbV/yj9hpUyrVUsm2dgIsWQciY0gYx9YoR7dLfoHyY
SS9iDBLzOM5AEh4KE5k78LxZU4GXRFEKX/ea2MkRTrvq7eqkqZw8QdNgT7ZwePSf
IMTwC1NRUaaGPkWdzB3hf8EfeKmYDyZQIQ0PqUYagB4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 295116    )
GLEwlZkQaXLudK89S5xanJtyQVbC8sArZotU8T0Iy/I+Jbqv75IKpMqCryoq4Xpk
UzoZbOHBUwjtKUXS7DePqthdQsK8QExEHf5XzsEqGD+QSJ29M6NH2JkX/xjE7EbC
qVruOJSLor+HtwK5LmsPNSz+h51W66D8azx1lUjqXBkMhkcLH8bqvl9KwI+OOeoF
KnMVGJwazveshqTvy6U+w9HYD7DS71a7si/azBEJ4wWLv8+nXiyRO4Aq3gKcPx1U
oF7mibETV9Aqgxq02+31KefqJtff8b+bEvx/sgZxnlCsEQEgcQu1bnv8jKn4Wtpf
0MMhFOjemt1mQ5XLrS8QTQ9SNSnj4XIVhTsEwvgIB9+RBSgXRnt0qBJ6ojvvKg1l
OIh+AI9iD8HplqjGTnIQO3XLWW3Wk5WZ4bVHc7a1J4I749QdxkI/W6Fgjz5Lt8CR
4MwVH/VdlRzQpC05HEKtZ6Ua8DUHQOyOTSZbDZTEOxc/hJczFGp6wzYfc/7XpcOY
Vbmjp3WQe3JA4fPGwrQCygxZesNhPiog/CrvUgbRiU6QeU5tnQxfxgcYEKtsWJJK
B09NBwO/FCqa2LFZkbSOB4W67ktrr0Cg+Y2foGnOUdsHIK8O1UH/DXhiR40eeut2
LybhuQUkFs9FCtk5AI7Z23A9fWPsQWiC6/u7KCSdna4ej1+JY20Xw2AkM40fdPvK
ItjsyDE7nRbXv4RPnU3KDJA795tFA0HhXdUIdrzrI0nkLmAbIcA7BDuWZE0Yvpol
q9wxA2C0teX676QDQXIdbGhTfreu8Gae+PtQzjsgNkrFo2dfpiTnZn8zUuQy2+IP
VTvspUX7u+qRW+tq6AddeedY0lL724CjMN5MUeX2FmsxsV8Ls9gCFXxgRLLICKfe
hADQLDdL+nyZ448TdUIo5uEdaBFm6GY0jRPf8LvddOJT1Q5EmhBuU/R7gxOI8yID
Kzsn7e6WPKSzu9kRi5t0ICeHwutLVu/fPzNqAPJymKf7ZchTOSKWPdPRRacuQ/by
`pragma protect end_protected  
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
nKvlyDKbNxEKgjzKOQsLv0wT5J8T9uqFqHm4vZIP1p8MhqjM+nd4is7pcT/HtMJ/
ABD2zJywxj/jtybao3FHv4Tt4s8OJjcm06kpzz+eTHMSWfxglowVbRy0Qz7vsKgK
v935c8/yCojKSohjqDb+fEiXuKS4VCsl6rTYINvnJu0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 295255    )
oL5NtoVr1La5bykK6rbZsF6Vi9wsRhLGBxLIelkXmpiNHRTmHD+5aOvkCxofem57
Pv1oxycTzku9on6V/a+ChC2LJ1gVmHNm2BSiMYSFpu0jPYKuLfe1zzeXMFiby102
GY9i/8h7P/QMY2Dh3TBzZ1Fa3umqdKbuqkGH2zTr680fEPXc+l3l9v9Tn8IUpgS2
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ht4eRSI4Rl7OJYpeXruxYAEAm8GImH+iNk+NmYkdQHGtGPrTz4mfDZjWlb17lBd2
l6497KxQXOwpAz9GyvPnUF1h24BqYpqBuv501RQ9UlBT1Q2B3dKOIvFqIGMHqxeP
MoHJt8AvHlxLV8d+yaU8kKl6TFLbbORfz/uW07WFWgI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 295937    )
j4ckOaZW7XntqGEMdYWtisEgVUBGYJtOTCkSojwUeUFMCaPZqz8FpMAoxUkGqb2T
X2ClVgqwDG1S5X4PjFLI2OoEwFmHtRmb75HJXwpdiU3Oh6J6c0BWVwdAUomcouVL
Veri+7rD8GwSl1VMXPsyByd3lrttCBeZJnyBtdEUH9NgyyhVxUe2LiuYCoPkhSSi
+wwDECTW1voCBJd34R6AS076FTtT8nWKLZGoxfUVTHRmcaYqZPwS+mpXko9axB20
2mqEiUgO8lbmsZMVgC3vte68KRO1mJ5KEs06J7vyjsRqm/FhHaymzU+7ZWG5mqPb
iVyKu70LwHkLTO9cHE535zmKFah4kdb0tWowZLqxgYolOwmkiV6s3iFiihK/gyJK
bVUBxMakAUJCoOSHx/HSieKFFOyfgtBV75ZV7HMf/OWAKFOE8b/WK8IhQ+D9P9e0
2mvfHzS84L2sEFZ24rL0ycxLDy2JoThXaVxO+sCM0DVFaF5yxpM6vpC2u167kAwz
pWnQzcd3NXcgvpBx4zTx1lQQfmUXeRSEB7fXdxco85rwhD1FKXAD1d14btlUxscD
BThPDc1o3G6tx7IS5p7VWRcEc//SMyCyJxaKhfevVXkQcNIlpLw9r6LQtZY07Al8
MNkbI1dF0RpOi4uNTK6PUhEqxOs0dr8BxoR5aUO7lvDjWgNEqDcvRipU0oMXljHX
g6gC0OG8d06Gz0LzXs8iV08cou484YlE5z9MvEtf27oJrZD3rQaSRV3jYhHh5d/K
RUb2a7qD/+l9w55uFsTrT4CaQA7FSPCipeBLJSm3aiL+nI5VEwnkFGtuiwSXiYFh
RN3vsVJFUnBeVgKzW6T2yjH+fDxocVRxvaGIoHf4fkUG32IM0g2VLKUt07VNpFzO
Ni4X+E5GWctVS5MBtGlJeA==
`pragma protect end_protected  
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
XOoailBQ+F7kjErAjjS6aTL5Yi13h3tXJDFyn7q4vrnMrad64gjdYHQgxMDjY+sZ
0xB7FbvJhnoJsQ0U+X/KtnBmImjxHEldjGy2hWe+JmimlCWmHAcseoSz28HZcOqz
gmZ+RT3tl0jQAnSlzUJkFTyEiuFwuQo0VqzatTFBwdU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 296076    )
nX+050lZNRi5V5THIeHvh/u4LJwX329aR1ruk5Mb54gRAXFzLAkMYWPdsce97A8d
HMxi3bwWsrRWU5B0HKgCVWpQfE3+mXF7Y1VpNiFcCq96BxPXxt5I9xgaAR5IOp9z
TrydcDDEo30MSvxxnVirYH2xkqLFDKnHafnxp3n2JO/fp/qT+Eu+Mo02UaDUhCs2
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
mg7k6gRE0bVjzGCtZqhV7C345JWP7E+gkkiCmxXfUFX5TL8IM0i9GJ8Z0HUk8mOs
guHyqAwX7MijBioyFBLZRLZS87zuX8Hh+I5OBTnm6albSVeTMxXygUyKS2JMkLZX
HzqNHKbMRCNExNeBxqGvC6IQyEGn9Uyh47osC+mBJHQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 308508    )
yhSwyy1haYXylJ6Jq7nxvp2pzbeZ26cvKFpxPk2BOHn6u2Z+4C1DxyT//F16ywRb
sfziMN4I98xM+7H45Ui9K8vHkfF26z+XqrVk7yNH7sXLPGnT654PTroEKbRyCi3Q
z5DePelYXywsj08jPhesohmtqYA+i/sDfvN4lHGfHNabK9kFm6w3zmBulK9IQ4Nw
a4pGvOLBAX7+65gwwD3fPbLBprDEbxoQ2LEDhGG6LhYE4F+/ws9UMyzymPwk0Z+h
OKIdi8MCKrpxlZoDfEBE7yxJq8ekc7OD6MPczFIYLNN8xI2nn1Gm+OuEjpMNrGEo
H7Ik5SE1HRwvs9keaC2PTJA6oTYS+9gJoQGMGgMHKEU7efHuLhYyfI0W+fUXXTVE
sEMyJP4b4O4K+QUmp9W2iRc0zYhbi18zDHU5LnNM2MZtFEv+s2UrFyP/5vgIcGJz
F318qya+XJfcNhpX+xUw1ZMV0N0dL1V+3nnkuxiFDJHkWZrnv2kcu6YcZVP7GFYN
l2gN+ZykNqBPJkjLNcchtypr4vCF+cWty19x6SUwyUv7ocn9kB5FpfB7VlXj19tD
q9i4G18Kh3QACd4yKvFINxiVHnJQLK/GabdJJcqyG8Evixhib94UfmNY8yOjJrRu
CjiLj5pDqjQIx4aMGoIsSVBptW8Irc3aLQ+pVr+z2lKUOiQmjCyTnIYQVi+E/glO
t6r9Tb8aMppclh1XIOafDh+7cchcgxcicF7NKCFDCYqZl1HKqKRQm1IxsJehcTU+
kkp/LfwsjWGy8E3MyYPhULdqPdGmHX58AtFmxkYbxWvhHdfWzEhZ0y9Ln/l98Cc4
cUF/FZxBZs99QNbvicWGAIxpPZ57vkKfwfnhlIxDxXANyekwx/frIKjlpVweFC22
MEvk+TpwW+kk3+VkIELuTIqGZZN6kkAoRF3rwLwanF1DbL+j8XHyo5/jvRVjoZMa
u9wHL8dTpPIM0ufIqfRreYQcaTOpnb7QmjTeq01nyIsjc2FxVEdlpEYRsF6bHd/r
6fLhA4IzuslEMaRJoaqcVwiFAnF+rP3I9xLWk1PvgLRP+LLoB/8NRkitFMrPl0YW
98RiY2wM2QlgLiITjuTg5inBR73aLIhu5OEKM0wtmQeRqAFVmHH1gGBbCVdD+be7
40K9eMcv8geplrjfOoMZDTLiBo35wiKUXxmuOklzsguJe4MM7F/k3qk+zjvzhidS
xhv6Vqku3Q1AeUeOk3YPWChzr9d/dhVVhQ2DyJP1giO4DICxTOnC/4dzFGiPFI79
auNa5lto154+XLjseW2wkOzimbugx02ue1FFk62Dqp0agf0Lz7u6wluSf9BU3V2u
/JpSfZw4/Fvik+PJq+DnS8X7+GnG0UJBNJ+UtpUnvUArC9L3xfIlh8Rt6uFvvH0v
IFOcOU4xlFFppSYVkTvX/g0bJ2Rz8NV8jFUSPiIfNjtWnT8DqKgY2J8Of39q77gq
fAzbaJStqVEhNvBcPNhcUdMa2TdM6hsidSbjulTLlU2PIbHCkouIpBxXKTj4iD1c
/K8RoNzdi9FSGgIcxv6TJyTgZYJ2io69ipNh/3pI9dt+HoGWtDMSh4vtrMoCmFTU
rk1D5SeNp0H4CqZ7vIim4NYF1wDsiAplZakvDk2Y+9/+jrPMd5CK6fpHbkPCboNn
2uS+CLJ/EZAos8X29ckGzZriL4QHQJjoEjMk7aGBbxr3txPtQT0KQB8O4zOXY+mg
YocwwauoL65sv9GHQZH8Uqr5+ZmwUKXiBbE5fCZOXpL/w3hd4rgV4m60BKGkzEsY
41V+7sEou4WWCbaiRGIqgaI2AlyeT6aPajLR0cI2upd1rKr25tt9f7lZO5gSgU/g
4OYoH8Slc0pJAe5b3XrSp0rwko2awKXzgGaQI1YFoDVQJbtn7cdG516xzZ1p2+YJ
dR8Fn/CJaLmIoGTjNlpU2wxDRWo6WlWLkKkYykbODn7y1aI1IzqC2gFAAjv0k8Mo
qC4LOHWsDo5Ednk2jCRb21gFdAxA8U+hAVDTOnt++6YQs6NQj3ipVw6hyMVv2bU5
e+RQJd19L2XXUVor3wCpv61ti4LoOKYGo2JLuoZwKmlk3/gPmKqc7R8hxSJaJfUC
9L8R4aWT8LqRET0AIcmSNoGvxTbK/juOYSasdzzUyxU7PfxpLMlWfloJ0rux5IA6
6FWkzTqJW7p9iK8lpfuHKFVzlPDNtj4FxjOmbTMJAks0SQ2TWaSjMXzTuoSyrTsQ
iqzqqFiWBy6kUj9KoRF6fVf8AIYWxIs25CKZuZsGlcvp50BZBX84zHKJ7JGeE8Mu
ZTAyOQK3DEEdagLs0vLXk1N7dtXqrabZ64uA4QvCiRpS8PeDCKXcLoIJ1NDQtS3K
kvccf/zvHAw+mKz3RhmuVzx/mghHSJVRXEXP64IK77vNLnA7D6DtlGKVXDzZgXfT
wuDcYZS1FL2RxmYrSXA5+eF9+Hz45wLPhXfiFCw2RhzXNsxVADyZRnwtHaPa+RlS
L2MJ87qZIVKe7xodtldHPhVLJ8O7z5+FLUXxGjsxcAb271VbSaC0qqTgiDtVABrl
XcQYMKkIubxy45T2BIpCrs9bdAwtyCFgvAVcSRZXCfEBfZ++fMrVYVs5We6TZBQu
dQYYEeKT32vjmNzj/Pc3MV2c8mPHcrwWn78UVS85b1yyaj+rk9KUVLfW2KV1p9q5
jKAvt79XZwRrUNZQehkPi57E0i0+QLb9Gx1rrRN86Oo4QJM0jxr1RmVPTCVB1pva
5WvHF2H2tLcFljiqZDl06dlAibkTm4lDYKzIF71rUFYhOo8dh+nTIgLw42RGoP4H
vye4NFR+glYi753cvc4+E41j2HJFpI19wBVZdHYjo1s7Wt4Zx3u6X2L0UlC7S4wf
1OC4cQx+z+9fn8Qy9piDI36026n1ToiPEKfB8k3LXvxj0jJpoUvfkT/4+6Agfizb
7784EeyM1viGIJKrZPm0oMx/rEXI8SxwVB0M9inRLELoNVv9lwj2xihZ2LLUnu7O
mtrQiHJ6gC5FjW0T+5fLZ+pi1PXccDD7qmOkyA9d3RaIazfMUT+nqpJNfHpZhdMp
FSphi6hq2Vr9uNes3tYjxw9F0NfPeuzXQn2CKF3txqihCIrgbOPLxo4rJvGxlien
jD3qmXYXH4BebgLEFaeFmS1aoKFUMsIKszR1PPvwS50uADK+7r58IMYLd9iwGiGv
T6v9nthwCZFSqgQo0NH8Vxd7Tx1xq4LH8O8vEyBSaX/8M+6IOnxpTnRYxFzGha11
xqPzJwf7eC+PVeMjDsMd8ZtIiUP2/wYN1M146XF/HfA5dE3CRiL50Kb87JXWiiBR
lHmr8LIykSE/XcD6FpsiomLMb3lZMKWByXhe/e3xOqPBuZU+LRMSyYCnvybFLkXo
3ZQqq+GLqS7yPmYhNlVZaq/zyxvoQx4ElrUtNBhn0GDZf9JH0BMS/uDYl/4XeFHf
vlNQldcMyl7OkAxg2dgKUTjE89H1tcD/Jh/v5JffyYl7WkEnLzvmTIVhbbJHZl0p
uXL04scHUVFrMvKLfMnMs6IszFzKtbaLBnmzssp4mGpDScviENJ7AZi7MDBIGqMi
cCfNtBj+1iBmQ/l/aQJmvG2ZHGXOOK6knojNvNx2OSueyNQbE7mJsPwowkg/5Qzq
cIg9us9g1KLSNgkq9ocut9aQ0uxNYQp9CJHwUayLyEbrVe8f02mt/eIYUvSlSui0
/FIxD6N79efb7woh1juKD6s+bnO5INmxakIChUD+1LTVzk89RCuFRqN92rFOw0ny
25WywuZAbv2rXECbI4r9sOF+j20LVm3MDcwsu+jS3VKpmLVbWKFM0NAF8Gvu+zQ+
RVMkNWy6HyGZLUne7vuMCLNcVV2sFws4zRjWZfX+iWxNgk/zfnLShP8aFHif3Mnf
Sz0I4E7zg9UP+osmhxLmCqH1sobAX3l76llsEPGYBNjMTC78rEupltURy7lcJkzD
GnXcNrroDviaostHS3/RaS0hxH/r0jCdKBu8NNHBM8BL9mme3/TJej6IGyfV9CRo
m40oYMWBFrkfca9c2NCT3gn79aBS7BIsg4nIJp2Re6cnRWCAJKjnT/P49+iG7Y6/
FebABa738MFDoJbhdXsX2NCbnPa4Jc6iahZsvuJjnD20Nq7v1FNuPxG3+4Q0L/3b
oYRtoKA3Elh1iTZMO9NEiMFLpP9MsqXKcJgcuKnmov0Z4cZtlGBNAbcBqdvkBcZt
feu3MXC5B2YBC10UOHtUtp6PbZh9QtCna+UBsLUxOgOB96S1B10xtil95REtrrE+
Fk+T09iP7S5z8lAQihKgc4xXq08JfAdNHeNGEz8pLsSy2GeJiHy17Tf27UpVd7n4
Cph7U0plrbv0sNV1HHZGsCPDZLKfZ3CeWxfQT1jfqpvyp8ekm13z1lRrh0tQyqI4
1ahhK6FsQeNgjnJIEmXk5QzucztGRYuW0OeblxE6uPbn/JQF81KfS5ruuEGlc7ET
Kwwcsb1tfTzMVydK/wqvzrT9Xwq3o7td6bzePjMmLSKq1CrCJTqe/QN+z7lIhYnL
XoY6FrVbEPzNIsaioCQ9RXdBJirkydswLoHQBMNkYMgjK9dfAnxp5opMNedD6w2g
AwIJYkDZOUzGM6VeMAdbRPOh/aLTBqIK5twygyftVkb/L0fq6KTp48HQdVHolv0Q
ntrekOADx0sfFlkMvpogW864NwFRPzQjRsJ9v9/Pr2ylisdXI6PkZEQFfA1VrvNT
HbRfnhMUadVwGobYHreOj2AJIjE/LQzK3RAbRiQt3Gu9PnTqM1PfM3m136rbp48k
Y2mcnxSl4zV7UvwXcdO2BV7KJTzbqqazet06U924+wZCfPjGYmy/K4Q2V2lh6WTg
00mB98/aPfzmMXarCj8S5te8crPrZP0FdaIyJHq27Aw8Yn04c3+pnf2AaBpLjcQX
nkd7HM22kXMcH6SAZav1H836OQ9I7yKVaFKnmalK3aTOsTHoC3JVwzmvmY2QfzqU
KXyitub5FmaZCs3TtBTRT84T3wWXNfTfwMWS5RHSi9D8vs5Ts4kCigkPjVnM7Jql
hkfnsZmCP2xX93V3SEe17w1zlq69UjtRuX+6iKy6A6EaxTVA9n48x6PKF0lpBKlX
Lryh2mp++QWmCcdntMlBFzMDLJGtQrS2dW0atR5N3KguMk9/ru5Re3v3vSc4mBBk
qgIbeXcgaiW8VlrOrzHL6iK2JH6XF8F1kKuXp46tOjx6sjg0LGbBPuDAfHg5RRyC
EhqYUjg2gDzKBUQUXH/n660T5BLLjtGxDYnXA4BbG/6aRgb+ctx0KjJWQs71ZZZL
D7w17ik8HA2ZbuOZiQoBoqcBx+NcqalgUhXhaVum/aKItsPSL94JQ/+q9nwSQAXl
b8Vb29ElswhsWeLJxKIQ8zIte4Al9HGm9wUu5XadSmwoiJ5L2om6nDRlQFk2B8Tk
8ES1a5tT7rmBP/BtPPyS3Y3QPLwTCi4kpY1sTFeH/3K02Qpt9tlUsuUpdhJn0Pdp
2kAOd5UNm9xzmWKbSwOTVVdMfDj18yYHY3aXmodZ67dHC/09LZ34hQgW05gQcgqb
wEQSGnZmBvG7lOgWVcn8yG5UXuIU7i72L+bp3H83mjDvk3uPlY89Yeqa1I40699A
2LGkk+Ax93BqAGgqqQG8U7lBw5P18Z2GTsrSvYUXhCOnED0gStz/JQlMXYZ6xlyc
49Sehhd9R1zaw9++kumt41JcFzBvnkRUf3iaCOkx7uRgyaKiEueaURvsfCL5+Ui0
iCU51DjkOu3wxKyMvTJElPD38RkvWCMa2KOPh0cpa5JLi/QTaeuCeAHcbn6W91u4
rokRcWtNrGtqtonA1itQmxgki0owB30tHJtpeqkZQrqcvc0hBLMuUXSiYp1WUSj3
kf+yjqWUjU0NFPm4V3WF56NzPv+kssrIE0V1+eNRFm0+eY1UWCGYZ7I8+Gu2hS0B
PVyuXXYjLbjNRftWeUGWcqyYtKJAFxRf4EY/3zM37sLhqo9qavxs3+6TAsL2tCKk
aj/HDYBR/uRmTrNetM8YOGd2CzXVyueW6vPQ9Y84KnN+QLopbhEWyOzPY+As5xbb
+0MLeSoslZYD/8nGwM5TaJMj9IE7PxsNw5VVusw1+1PpBAmhc18m6fRV+L+QsQ+t
QxkJepc5fEegLWz2z9Tc0xL+nxaytcjY4ok1nAAgf+E4ygb0uP3yQZToeU8fOFms
cP9++D6VKAeJZr9w+3y/Bd7eHUguiwEOX/XAfeslYQLO4GqbC6cHVes+Ddi9v9hM
jqTnQhNp6uX3K4DN/pcBDATLUjC9HOUDhIX7qudHGRt8LfAKDrWb7dOPaDtDCZ+R
Dy1Zt4pi7OtIQmP1j1SnI8EekO2O99JHcFxgzGANiI0VmHcd4IBZFswfVo1iocfi
ZuVSMLKJkz+XqEOOTNToK+zrTqtNiTpfnGzAFfVFqobSnvGnn+nVaKEvs7bdjvMw
nxOCDSVGPZKmT5vGZBnif8O0MAyJhIX6vxPoLQxh00EH8ykikmvutJ/lpGW3kbhm
enAx+eEhWrUTycEGxkwfZ2vmqUV6ETA0D60RRZQLsKaeiI1tobfMmLayDQDB4wK6
quLIEpvOgvUj6+7tome+L4gEXaYJNu25BIJcieOE2Lrboyuri9hGE1i23GmntMD7
kJeGjfsLYhBdZdb9tWOaBvEttFeajL8/8EjsZ7zrx1XTeSNWDI7PL91ulIPl2z8z
zr0esY8crOrqqfGuHCotlDhoVFzN/wch/Vh+h2CuBTZJDUZevvyijZgo7GcP9aKd
sDhrODnrbWsnRGcchvBm4PQ9S5bmc+wA9+Nov8U0T2/s8btoWSQQfd13Tw//5Qn4
DYnlG42cshdVTdGUYA+EXXF+o0duihXdqviOQCMcHVPYwtwWaXDgQevqvqewK1L4
v5hMQevn85fawyRgBDfcMq9cOZvgpH70/Yf0IfgLDhCkg43ve9kgvxxJqVRL86AR
dx1A+HNn+dft7jGdkmMXEFcjcl/+PgANuoapyfCcsk6JGf1bAhwUJ0ToWQUEqzQx
DF37k0wj5ZIDw1GTlcnMUVz177UeXpioZfyqlNunYax1LSE1XHf+7KzfcXww5i3I
Po9bhjXQErZF22NRJYp752yWyAevTERIA2fPU5ixxi9Zp88+IwFm6qVrWE7DjlpT
kVp2ORagpnIX37yuwWzaCmyTQw1p/fGJimfiHW2ypsOIsE2+WUsxNKxHEP5qPDZ/
CEkITSqMue+wiJQ767bQpU9au87Ohfz589qdKan7EFNnfEp3es3ZIcJ/c0jzM1Un
gP0uejGGXJbTqZMXLIt+xyWi9bhpH5larIUMbSypi5MAQt4tt6e5jj4BuMEtm6bE
eUdcBqUvq+8ahcOYaFVWu5kfbDcH8cD3OAGsto36TqNHRLe5cPGEGhlBHVUTjqOS
OfU1h7DAVWfEVNn86/+HybJeh+r+D8EjWsfOoVPBcSw/cogEKUe9fVJLeTX2G7no
f7tqEn3I/ivSQ1+WSmXJEbHlJ41DPL3H9+p8szs8wozClgNE0YVJBJ2Jvff4KYFY
vbMCIFv/Llwx3R9LM9Qa40ZFgzo/s08/YI1JPWCNdo5Yv2upXbNthW8tq/+hKF31
x68EYqkkUvPy0QbuW/HIBtOWSCIvw8gzbLuiQXOqTfe6G+iE5G5kk2ON09DcmaLo
Ni4ePQEFkXDhoxvDsLJtxQfk/3ElqNVj8wuauofgPmJZIN6T2A0tRcanehyYmhIA
x8Rs0vdsSWjgWs2e0lvb3Ne4CSvt/+yjhboY2wlXbKqmddkU0j/E9ldANL+zzvzq
1LTrF7NzE096hF0Tb1P9FmGxSW06HZFn90uneJ0Vel7aJuVD1zsYd6o2zQsc9bQA
w9y9BmTaxxGrZPia037aeXfUUYZc4TUHJ91P9vtbFmlfJPvf3WjTrqRMQkbNkjvt
51cHJP/rxaUzBOXfg15OoThshw6ZaSJehAOAjPPsx4uo3Rkf6Vvt9uKcpsBruNmR
KtDy6F9yyhDEFdYw67VkblNY0Hm+WrKj6imaH4j1PlpS4PqqWVuIWbZi+1AyDJkJ
83QujWWar5d6a5PtJP67rz4U73PgS6LEGl7r5LqWPvH8UMc7NtHNeIft7rX50K0d
+x00jhRJzwJpc4oJ+1VLcxbpigkNeN57ZK11nTsgD0R0YvLVRRCCQERbAPvXOrz/
cAxEmMwVWocCxl1Mmp5zpwlbo3n90bobzUm/BhLOKpnm6+uHxJ1uvwRZgvLLtE2l
7OijVbUH0U8lBRdYtAwDJq9EMND+pp8St0iWmckFney+rzcKa136BVojkYzRiJiH
7nqQZ7D1xtp4eL8WrppKl6gUvAjR0LpQuAR5G+oprmhkyM9zse2BBmjjJkBwMA1S
TqBGUNbGByjTGvnEGHpwv2rlB/jpD6iZeumtr9dEoB4yN+A1qvmJnrTGhEu1A3ov
Culyh6zKimHg8nc8AwBIWY4QBykMt2T756DWPPFIiZKJ3Gvw0jP8Cojr2vmFTWCh
L9kJ+0dKd6bIwD9/RHRaUENNyAty78sr3MdK6FMa5Vq12vylnX/Gu5sXuPho3jGf
E5itI66R/81HysEkQKVGGNDTjBL+U8wD9H1DTJyTcptsyoDE6ExooY80qHbiZbC7
+J2yOFkhdWBqW5eSomKyfg8ke5WF0c2uq/DbatGPy1teINxqKgf4ijfrR2ib9E4g
Q1e8pZIlI0QD0TvJoWVpi1AfSRevFEnTGU+DnYJf600uNnGYu0bdwyNFNAU66YwV
BeGIwcAV0vcagvjS9ONRQ0TZdkcpRmCSJoT9Pw95tYjlQr6KZZYbWe4HRCW0peML
BvqRqtLF97ZyGiRp6aUsMtmVez38fdGy7GbEY/0fkzc44J9pzoGQH3tWubv6k0yG
Jiy+2OUI3FgCfM+TCPSAtQ24NicRZ+DQUVjKaWKqDh63liqXjieOXpKo4qIIlzfw
kQFJatZjptPN4kgH6taZOq4x/E3XM+1A4LAu2t4znswgGOFuuFBZWlhTafJ8+rVn
zWymGFI4oDuAvwGhcs5GzXlkH7veoDnjf0wYyXVfz6GA7jW6nG9mM7rh/CrY/5km
XZ0XraK3BWKaCmR0tGXtrBeSVPMr/j9QzjZPqtKS+WQ7fP27hMHuGVoYAR+lnMfv
ICpFNffbngXCG/P4936eESsrAk1SrudQLp23TJnwtS7d1jChZAx84eKgt1qnhjE2
Mxj2k4Tc9pEhOd9lLzeDENZhnt+9s4CEl7uwWQBVL5+z+mBYTM5ywWa4xN/xG2iy
3FhcHHRp+dlV2RpXsIyyjDdvekX7kforFHgjREe3q0a6QSmjhGMo6UdMOryblC4j
MvNnRGrsdB3PTF8IdNNkbrYwVNEZi3o66maPwr1Jg2d9l1DAJjpLtk+653Dtkqz9
9Gw+L3x9Q8jJZ7msuYbRbzCGjw5dSxCvy823Z4PyOu67EAztx4YS6ybHVj4hc4hC
itY4X5+aWRNoTD28fqYY6ahRi1ULLBeZe2hIdqoX25hE4koU6EaBZFf0xbUsU5Dv
ZmGI2PVzvCF4Vq1v6qldCNBL+rJsD8V1db3yj3JTwa8o1INebkrS0PkZeKBCXevd
dh3MSpz8/jVExvby1dpjf5jGCO/zpDbnrHTx3gORFtvLIga8GsPTcovznPSPs7Sx
xS9Et7uCrYWjMobRBL45AveWXwWqGUEIJD0cAKIimhyfJbKiL3u3StWzAkO6iXFw
ia5RGtCH59iBeL28Z2PIVzP74izJQU0MCkK88VfU+S6OqdDaHFit/t3YSJ1MweNW
KLALJQ4of0kNB7dOyCTM0B5Q4rsNN3gTX4IwdjpOxXQFeIeEQmieWj4kdvqJXZ1E
6nn3RuZGEDE7wLAZe32hmcUBpyVXDAYFlTLWk4OCVR5wsSEN76sW9meU3aXq7FbX
gRnntzVLO5lDleTVITVOHaWGnRLFwizb+cxSIy53uiTVvxmq7VBiTsVdw0plHb4I
Ug5tIft4T5yLF+c7EhiyoOGoKnGY/DXbBDOkqm+r5PFU9SydauhbNhskQJ3ZsL1y
6EGM33AfQuhJUFDwW+IAJUwSnpvtbZ7XNncDsC0szt6yTV9ggzDRrcwDgJYWKKW0
ZlXQDvWU+je1VBsKgOgkWux7l4LgtWJfXb4Fsqkh9F8tNZq7cY8iSKbm5bRG/lDA
D3CtTcxkyh4b7SHqgm+XvSh6of5yh5i+wjmTqEAuC+ushu4/0Xd+n51poSsHppn3
zhXhXodAffwjv+7WaYGX09fxN888qKabLXaZOWq1QCTePgf5iC7370LZjufebmqy
AZEHB9EREVLTRwtiy2qAtfwTl4ah3joGtHZ0LMn/xUiD2NSSPz6h9ApwdtNe61md
lgKDDTsDll3sv1eQNQSFhCrssc7z0WIwEGmNgZTaT+NI0LDn+twB4R0v3UdYkcuZ
UFbuk8inr+yyJ+3sWRvBSOL0IFo5up52VJU9J/sYEllzsX27GyRP7FzE3qQVTgEj
6lj7e0fWDQoXk9eHwgb4anDIQAHwG5KiYFpzlS/lLC36nbR9aPLUNJ9n2f0Hrx+8
J4Co5ZIrVEotbqP2FiKNLVP0a3comY5K3d35OBbp+qWKrxcuk94/MBaubpgkCzXH
Z7DTYBLLBNMqZ1nKfqI17tPNipmXWLJcUbdU5jdq7j8Ihv/VqVU7f7bjt8/AGE40
s/hnOj/gd5+SC9DX+PdEtQdbvssOvOPlujbRsz4zocLJo+P3SBWFMZuMbas5ab5v
oeG9yStdQlGka0ZpOYuYbApSf/1Gq9HL7eWKnNXo5245oQ/2N1S/yOUe/8j5bt+R
nKnm/C0qQLaUNnUJ1o0Uss63rtsSzevoE72eSBf4j9wfmZbLa4oMLXZCzAnXBfee
wZCgo488e52ZX9pDvfv9vWliSqg+n5olsjaKyoW+H8czcy6rTOm2WDnk3wdzavvw
gFlHBij7jB0d6EOuDqXUxVYJdjLjzoZhn84P2axX3osM91fdtNbLDigziCPaBr6a
DhTv16waQyciy1bfGxTyA+eYkWL7NOQXQv9JkYPXCfx3cexNA6twfFnIMl0rUEzm
niAeFcHTeF4gaAakFg2nPIE2nWOeImkWhuuYgnwHiMcndGemvxuit5xHjNRZ3ZUW
Rti9XNctOfpmRW4MzgYtryPfY2tx5fEiDrg/BQhX0wjfFJXnV9JGIgTbnlMorVLj
4+ha3RlPUrmsZFlDMCX/x+B0SHqGELVdiDSn6OGDlzMRHFwLPHrJ9G0M/HEQzLFK
5lTlOr+ES7053ng2/GopZ6kcsaHCK9fFVTF3kFZ3xcl/B81oX1J5jlTGZUjfLCMm
LIdi/uinb87w7CPnFZeaX9fwFxJ6wL4ZjRqlnCAKryILK/mUW68f1V5Wtc/ll6CA
ErABztQGTXUujF4XavwViqe2zbYShF7E9YspC3yL9UR5QLpahC+D65NXAOAGT7bb
tTsqahMe5FlH9NKcLLe6zzwRmKgwzXrM1AhRvsTVzL0Y/EO8rIs4PuhQNmv9fThJ
VsMyFdfCy3H/SIrUlWMasVdZEPftWOwNWFOBI1jA62GS5ZAefklHwwSpEfG0rsef
oBF61oxXyveQtrpFUtTGGG5kZbJOh+tE6pnoHFePdp07KX1k4Vddw2PQeAP8YdfG
Y7L87y0oMWKdJy5DiVd+D7jXzVK2JvFTjY/zyoK/kYOj+Yy10CPA1m8alDBRok9x
TyXbjmA6nIrPNPYhwBwY540HGC21x93DDqIeq/9VVMm5fBe78PCd8rjUc4wtCxKc
tO5qOrjOSApyNO3VZFaKJZHoNXfPbi4H61ior/N9hGecBTgVuIDXVtORJ4hymJLU
aGDnVMFEBkFOFDvg3ScA+LsjMiytAhIFEBQH9KURExyrFCmzQjch3owHoNsqPXzj
IRotWbCC3wKlWNLo9nm2DF1iFO+Ltmr/Zbzil572hj4j/9iUcvYgs5VqpUMUDPLU
qlm+aGGbGwz6eFal8LZIDDQ+bAqJdd17ilsSkYudXC1eGuWyj9mGr+qwjiyXDEjV
u2YzITYKvhD5lqgISTsZd8i+EUurNjuezsmHd8ckMvrPIYkwXlv40ChK+M+whJoV
uG/sEdxnYuoy78lq4wza+1cz01x5k+KMfw7aWKRI9ILDJt/MNxG+iKP9mJpSNPHn
DNvR+lBK4GoPk+Gwya1MfBkErBGIxzqyEFnfH+ULTViTsePmB75RISH4gp/jbYjm
44A8SiLU7TA9RehBkAYgr9CTGBSVSXNYs4nQBCoyWpHm3WFtyUJueqnLRntFqKll
rHAlOIe0dWP43t3sgvcbOEYThb9BrH3rIbEq4zcuCF4X5x6eMoMg7o/dKhikpKpd
6acsX67BUybF09MKop1Szwjivp+jXH/uIIKlliHfIUUDkZcwYFXf3JEaVxcxe5NC
wzDDNSKPfvXPVvLycwicdpCUG13vsX3wm3/bxNVgeAwkD+vlJVriCCtHE21GSITA
LE0Ch6ckGZ2WNLUZkwZgQDoVTYX2U6cIyFRxDaFOY83Ucsb540vVodyinJOcsl3x
8kktqKgMADchYYwKEk8GQ1HEEjjMoQPl6TS5vtfOBB9rS3E0HLvBPpaASAuNkQA9
erKW3iRNMuNUfUqfCWHKsBgxyGLeW98QjV5pIfkk9jzUBo+jr4NkTWwlQQ7nnk1W
pKieNeY6gNOe2SdmfWcatqfFnU8YS/DlIifoxv3wbYJCi04/bFx79ZLgApjqNuVj
DDhaHNMRJtXpV/XHR0I4rOc+j4fqC7TU/OZXJyo1sGy2YzS7963UsDOqfPWaMI0u
om0IlBIjAGtegx1gBnjmi2Q2AVPx7Myv7C9ka5u4l6DDKt7SC0MWXhS0cbucYuoh
bh3puRj/ojo88DmXdwsyhLH1RH4DdmsrECfxV6W1LTzyLmoolbZyiAJe4O4BIcIX
eNTkzCq3mW1y/xnI0dUEYhvRHa+WOXmqovXqsQ5kKUa9cqp9/wmEfkm56DAKQNyy
Un6NGjC/3Nz8ezGKCZXCxJOaPMvku/HxgJjxT0IQ1lcjxCy3d2+Cog/X4f98R8dc
ueyOZXrqW34DaYR6eduHoom0Rzqtc8vPmAYoGPIDNFvLUgPvzjlvxf7EGM92i/CX
uZvPUovQJLXQpxEFzKyjW9e3qr1oLWvaU4htOVXQcoY/52xuq9KJBR0TRwbwIAkm
pzGEuYyV+JalxnTo3jMlHBqKk5IjcNV/fgG7gWId1zA3nRjZ8UnTfG5/O+iQ/6ia
u5L8xKOZRWnP0i9D6T1jSJofoTL7/GjSxkPT/uqc1AAXRMrsO0rnaQK8qhX7Posw
7Jo7iV9KHlfTHnDuVuc5Yvfimyr7ZkJ5i0xdxCo9b0he01k5dHsp9IbmCudzVmb1
wl/POIyHLhwL5TLdxRGVR1dxSMZloEhdHudfl7VY5477MRwloz35E4N6mjhNb4d9
BrXyuyiBLXvy7C9CeGYU4t1AW8TZbsY/1rxI0TDnxwkcfGi/OpLT/fVkpgUROY4i
Tt/5VWcG0DcO5OKKEFFlmmfV/wjCr9gtMu5ApyAl5OJM9UGI/uYbvPdoUmhdgsfP
b3dnIydsP0/mD8EpPcAZGqz4+/O9fKXkmDDJQlGwPYfSeju04Z6UoOj23hVsFGlI
AONOSrcjV7yQ1UhVSb7MiNzGKrZWBc/Kisdd9YxKMgT8qxeX00rYQCFANpY5Swar
VAJMcOOkhPj+VydwggkQ12ZXjbYPknauwezFESroGKjT6PilBXvHKotQYYCToS9j
2RVadNcoPZAjRBySYEdC/L1jQ8MCP93swiw+T9AnrgomslAhiBgiugKcqmEEeho+
7Rpjq6cWYRxI1f78HbPE+17GZ+avXtK0RtTndc0IdwdX0hJFOZ8++aGZ6OFG009S
R77F/YkVoJ8r5aVDufoVpmXg2pOUe/24pYkmdE4j3BIP/cANNHpl0/Ovef+ZCwmF
6VaOG1k34XQgq7PoEEXFpcWx81qacYh6Dn7/zQ9V1vBENvD02PKzj4otw55nLN72
RXzPHzb/jVRxssvXV17jGZYH/BsbBGRf//uE8zahVr09XeARDR1Dr7fYFc3NW0DJ
IIRaKMJ1ziyp4yIMp2b0Cj/hLlvjvhe5kX1phhusQUQSwstBodNX3DBJTF9F/kF6
VHfNWwjyZNcZ9Q9YdD+HJXWeJ2hebg1aoqpvFUYj6iGYMdNdxw1s3NX7D10J4eav
wz/m6I/uV0r/I8GLgpDboedtIugjorN4jmm1GGLA/UwsB989fl+1TwLCtlwdEO5Q
D0XEEHK6gUoR6fx05vKHhzTG/x803Qb1whZnc50jO1Pxr13BXST2K5jQjPgGUNC5
my4KMqRELLcsmcY/EyzkffO+L1fGLmgGzm/HUGMKZ4hHXNYWQIYAR2ZcBA97nutd
LtGMjgqx1jBwJC4miHw6dHvKQUqCAg0BhU9Yd28YZHvEq1okx+uOMdKeo3Eo4JXH
gTgVLMrEc6a3ocGp1zz6Mm5bOxSQGrqV4Yfj0nSr114GhXJB5Aw3OBsfaYKWkBJs
ro5FTClmIo/a0oUDbpRococNotUKiJsCzgJa72Y1ru3Coi/WG7+4kO74fiXgWdDB
ssgk7omYa6YiiH8VlnAonrBF2nU19v6qPiReDCbwQSukucEBVit0NWXxK76ul+CY
ZAF5zPUkOSNFEru/ZABTS49VISbItAcIZd89niLPWAt5YCNsT9qWwGmM7KrSBTPg
SW1t2QG3zSDwUeiVvDSenYD1QJdaTqIfNV6rxr5iOVfFSaSKgsIjXnbucdtezIJz
KmG0qUxFYqzNu/mNlD7SoMYcRa90j7Ykc5+80dfbLxZZlxIkcPZ/mGxu9dvy8vzj
xtTriU2LVXe+BVMlVt3fhjrnL+LYF156Di1zFF/5rhwVbgypXl1NR7bJVtRvZyKt
8FOhH2K/xIQappmh7lh8FAEerxswOkt9KzkTEHN067vhx/eKmTHXlBeuQ+PeOevi
BRf60Zat+k18Pfq/MsP22oUuMWuqd/LshkGGboXAC4lmzDgBHaZ73qwpN2L/SyIT
0Bfgxi2wgWvpZN7SX2XNM+gyj1Xn65Tn75QRNO58Os5VsjYW91gsLxTDqJaFpxeV
2L8Qfnn8/sYzh7QfYoHDLhbv9s/ZvEk4tiYHo6VlbE725he/+I90C07FliZ3CBVG
jqyzFQEFPHLCIenp1N4WFYy5ck8U5O1omAQS5mVfOO8OAoRsWBq6/aJ82UEM91Lc
/GgU34FK6yy837rkULe1Mt0kHkP56D+1Ts4ivB+FxV+rNKlSRQ9X2QjRg46+jBNE
bnuouBgO2ieOk9bLaI92pUtx/6MATKInTo3+ocNh0ntJYTEPCYX9+ERmX003LNAo
lLB+mExTKON8xPXaxc6e3s0SJMUvJiG96cxORHAegHG5wogHjdSTSfHBpf6ZX+SI
qy6GJ8wtcE44gAiKGFfuq1op2cQoRqRYaEG64jJi/VjAFL2aNIc+YVDmo7u9xJNa
rr7dLDjzZWClBMbnmzcpiXxVNSpf9lpOfyBPlJr2YktxJoOZzYrnqby6urI9F18q
s/FQzlUOO9w/qx63oNZW+CKAiK+f04TpzCzY3bLyzgfslHKj+ju1iw1P9jvRNW7W
g3jRqVkHOe0wwNv5Gnz9tXzzG0OA9YMr7OgiCdvexkFgHOPRO7rU+u2b9g23aWOb
T3UmpDitEl/xxfml08whzwNMyji4B5+zo/oU912hxj8qT4AkQmd9rroQYhmhO5U1
jQ9PqXkVf4iLvTqlpvmwUyJCnEQ9Yii8JpKMmmBZa7vPhvLC3q9M/e4+9b9tGcRO
Csx8Wf9XZ9xUv6srbiLTroiNMXQg9X//O7QYBP6h0htMH0e2kO+kZhC7+q0pca9T
+OSV6AxRGyVzEMIRG9Ao7n8Wn2nWHv39JjJFzkYKZMtTOBMRN7RMOM7sC/0DnkCH
G7FEPmzBOhT7O29+PIi4d+X2vUfWuTbxc33365J86xWA0UaGZdudQXAonp84+cxx
U1ylBD3C+mTLzIQJ4+WvP0zNykWYg1yx+KZ2jwaalULMj1CE0LYdR0A/mmHuxise
eOOTRnkxWa2DFXPshIqw/0kgHoWRuQVN7amDXyNvije0HlYpZTH/3AYJuZz5D5j4
A+0rHnv1tU7b69af3KGzaELh+0Pa4J5A92Gvg6i60R34p03pc+qXvBnGIcf/4zcz
tXJ89GlCLLspNLPkmEHyezaEPjsMbZtjOLTPsS9Za5rvOmE6eceasrpV6GcJDuQo
SaBXY9mywk/DxZCG7m6BAM+Jy8yU3XYDpKgfAtbvCXtug39O0maJdr8UwsnzHzrT
hmQzldc+BSb2PDWvU4+TGjHwIbKHJZ/7B/RZKN8wccp1z8nZxY/ek93r59mDofG0
QGXpL4YUcT7qBnqD3gecHVfbGEJoKOffIpwKYhn1rbEvyCqIbNREsZX1JyorI/oA
wa9Kbt6N2b0E7bDi76SlqlP5sGpovlBUW12kHqPGmtLrSUtGqpozopAcsAZ6I7o4
xmciK8h/VkwJbyI9LEQjUKZOnheH3VrkwnZEpC00towQNv4wzX1SiEPUDuVaO9Uf
kGFJi8mnrnew2K31Stg12g==
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
AQH9FXKy5EYAVA5MHCJ2DkxWMc5neyM3oYg8T0/cOMximtnxzu+y7xNHHO3bDdC+
s75QCannLsW6Mtm8i4eRSLn/BLYpc5dZtyb+H2uJHOyojiG+qk/3T4f/Lksjig12
co+DZzHS7FHMr3y+xx4pFUkMkc9cPBVt4a7nsSki4Fs=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 308857    )
8AgXpDP14m9B4z1iqyHs1Ne/TJe6VQozuC5Gw0RudhdiHG5w0C6OLs2f0x/AnVPs
NxGb6pyak1iEu3H6s23UIXPNq9PVl2w1x67t5TFIZNSpqOU14e2xTXHl5F2H8GKP
PpZdPCOEP3teyP/zm6SmSLndnOYBEImajUDtfjA+GWvKEkFMA1po0htAxkXa9qeP
oIcc0LXOV4qQqHQK48fze7uTOkUxMhHWR6HMCW4E1ROZ8k/IsQ0yFsYUBJJU6uVO
vksHk96J7Hp/TNjkJVS1Ld356nmpXIBLOQXvv7wiNakU1pnJoFrQsu0VcYu0dDmA
ExBiefpI0XRUGRsdmkkDHrUXpDIwIpyvq6lGiMS4MX8/JuhY13I9DJ1WtXSFpfGE
JmsEb4j05nuLCnrfjt+0baFCyLsZncGWsC9Q6eLkvkPWfsJX9tdR0iRY/zaItqjf
+xPokk7Rs8d4VnRKCC1BSQ==
`pragma protect end_protected

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
H4S/lfBc97nuWIawe3F+skd5koHnCkH69r16wnF8e9Wm7wijc+h3oieuZOTcAt9f
ipc7D5GTRW9Q7lgSzrBPINGjYzUZ8YVEZYIb3chfPxZzJUX+yXZy8ehoaOCQaEsq
NYkVAibw4xFUL2K0QzhQb9azHO8KggKvTZipH2rqI5A=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 365375    )
0ROhp32nUA0X/yp7jeAtk6Dl3gFnKxTbdWAlaFv6KxK/30DzogjdntojrYy8KDrc
gkOBnIFP08S2fai4j17WgZaPbulE1K532+nD2N0YhoJ5KDrpEmM2lo1pFaS6Ainr
QX0iDG/oiISg3FYeJ5Fc4q9xJMlIZN2TaV49HvVDx9zGTvygAlTT52f21cgSQLFW
lJcnUdzDwMZBiDPB031k8CeSiQjWXh7pA1vIbWziz+3jBwBz9i0gcwjwd98CqmCA
1Fnq0TJZtrXlMggsN0N3NrDBHG5NLBuvs/8RR94fZ2WEledMahS4cvFsYo7wuae9
IhSU26mYXo9Ca5QapFbAmM62yfohpoody5SpRp4pdximnNxzkX9eakEc+ffYgrVk
NklXSo4oEf0pWcZHcfhZ+qvKjzVa0IQO+w9/WINy+E66GEQf4uVFn7R5KSOJt/XU
AMuFIrT8pnyEuvGvdEhlRS9v+eQgkCKydoIgtvg1wMDfASyQR3eyq6VMw+v3XQMI
JF33pPFtrk1X9I+oHf2VZYQLlwLgPO93KX74IWZc4y9l8SSIjT7RRkLXofGCbnun
6iryBTRgIQyJatBAwZS6esR95ymfRMKCu9bdxY8X1RUv0BLxiS4Lcs+Q9m/0i/rt
XDd0y96JJwcn+hNWFuvUBKw6fN1/Wom5FSJawcCpMKnQdHpMV8oL7BwCLjA06CRQ
dAWcmf168PGp6zok3vKSMieDV/B4NNTjdbP6hUlCVe4lununugP2IAZyGvZ+75Vq
AkQrueglUyUlZUjtJseJXbMH1aymxhWSGridVw4l+gs+foSu7LI6sPVCRP+hu55O
ZPUzjs/dqg2e9YLfXuwzE9J4XBUSPGZwH2G8BYzqOHojr5z+42RnxbJvfJkP/rll
2UX61/8dFqxoRqUGJkH55cmtDa/gYnr5oMzPAOTQwiAuVViLGpjl9omD7h6APgwg
Qd8J7Ke/RWL1hdn/XHqZu+RXsswa2Q1SWdBJ5vrg4kzkZYB9+rUM5LHAn+YaWCsQ
FAyk3fwCcgi3tM0JqeRJ/22xJE2omPLL+XbaziOeN66qpl0keDNGfNaA/7u5CBIx
VxvBb6wz6rm64UrN/BYu+xI6xmJbkfmUTCTVxT/6k7botTw8WcGQoGV3IAXNh/bE
MJeXU7jiSvNJJvIVyzhvoZf7cAUouVlauzEEqw+zlfEDaLVbT3Row5VwvRg2/MaO
SA4OPoIxi5R1xGFtA4D+AJ8sSL4n8ZO9nfrSlctirvKOf5GYVEOq1cmBDpTF2poT
cp1O5PTKpAkXmbIKENZkjaL4YsIMTBpilisLFRdfT+lYgqiQ2MN+sIL5n8aF2hM5
A1vfqaEzeR0mxsHn3XkJZO1Zs4WL1iCvHHrBnfG/p6KFgSt1cDH0dKg949QHwHvF
wzGMUamUYIaptzEllYCxYIAb52ArUBgb8I+NrqHpj520doFEpCrMZkP9obKqKRoY
nYkZJ6GvPfNWHN/IM7O8rRwuAcaF6vlKsXimVLkkpHQEdcwIw38Hu0xGcAs/P4Gp
DgdvQjjl4MAwPKbuChF1YdqoEeJ3tec+C2aCZzhn6+a7L+GIuwXvNjh28VZKJzJn
tvrGTipyzB6GhSjYpp4/mZCSK6t59sxFgf9mD5Evyy2fQECya+x59KYcJ508Ht2j
cbvmHOzvasEVmbNKBrBL+uXtR082T+Zc+QJkOpDiYBUU4kZBFgQ/LxMoPMJX2EWs
Cst1m11LRR+nKg5w892WEQu79yi+r27HUttZO5dQJi4+83WME2WfOkedhk2OQdAe
bsjOTV/mHnORNnPq0L0SN55kkParBGpMTEhM3hNgS1mERsp+3EHGJAqgaicXX78m
LYFbmga4SBA41QEL/75wOa22Ah6ryDGTdZE+Mr8ngYEQyuXzsarEa+4xPZn7ZZax
SbUo34TrFja/uK6Zn/Z5CIUlNrON/kW6O7oEPVuMyqzpinWo42Rs+7aaEN9Nb5+S
1BWkGxDBJWRfl7eDRddjkwyMavaIeWu4B5H+osUsZFrf3htFQL+WBMkFtSu0Zwod
/P/fr0/B/Jc0aigxmVg9wC9exZoPCbteDBecr4lubzj+q/Y/eqewlAOmy/nPpGV5
Ehyl3uHsnhC2pdoh4jdoo+SaSMDtaEagcrlhAbzbaDkhD7ilWdYTZ89xLMML2jwD
IVMGXlRx1mImHBgyI0NBmsloQ+AMg58j0JRfkDphUPUM6W1Z6cjwtHxFeElJPQR+
yIqtLAH3icFPseJGaHI+qL3oaRqTcMyMMO3NgTQO33Eptsa/lxuGfz3KHAEKLAcq
DxAmAYaonTkHnaq4uyHTilG9sBUayQZQQNfYt6tGwat5nizE0YQdAkMW/1orY43U
BlVHPnZG+qyFI4bmvtK/tT6AFH+Fq5AOnmao14JZs5+dlUdkHu+HBcUrGguqo/AN
XThNjCtlczOOigik6qIQgmMvZY1dm4xLczEE7IL2TvYm8jMg4ocZWc98krm7tiyh
OLd7MdjcRb9k+saPV26tSsnQvP52gUbnHz1/ZDcpDDKpUMB3PdptE2/iXAvfKaui
EcFt2fYC25g/YqxSE+cM81ItwZYLLU7M/voRT1rPykry+o8S9bDgcJ3vDSouIw91
mhiDVQzWyyQ+K1S52dRIM+HVlZEAzrMHdh1oJnwDv5hVXY6pOcjYGNDeVTOIrJ1l
ZuZz0jzjKjlJ1IA75Jvml0PLKt6JrF9fC1ovwhNrJTmwdUUBSSKNvtY677aCZ/FL
HtQe+HbhEaRRiYAHewr4c6mDGx0BmtrhfLiHdrrrYUgFYPXPiwapsULFVkbCMYfk
FqUzBqIUnwIoHpdrStAVDZ05RQSV7MyRefcxiGjjpK/ofbGBSR35e9ReJMkX3P6R
qT8kG3iit5xzYYVsznOja5zno9MoqXL7q3gjzvADXZIrlIMnv2EKVb6ncmQo2suI
U2u0KpDw7G2S2+RAiJcMvYgHhwRUEJuDOLHakbGuPmFo20WMO8Kj93BYrz8TOrQI
T6qxFeRTWq8vhBxy3YzD3+GBPwJDwvBSy2GjdCd+tIT/M9E2jQURqzMXURI+QZ0t
OWeUtrJJLXb0aI81b8ASnDOqeWJ/fI4YKnp+tdCRXTN9WoTi5jAqWQfx76zLr4Mg
HDb/U7yvRtNwEWA47cYJDBKNHl6YDL/qzvlUCkyw0ov1cJAv9V2j/TPnQqkLKLBd
foNWpOJua3GcYU5oJJJ1zhcU0bb+f9m3fRX2LdeJejxDINzd7Nmd/RrDVO0jdD2t
et4R+mrQ7+w1M2btsZQE1uGpIQpVTz7UNgNsZ7W1PY4VP5Ck+REEi6lXCadO2MWu
Ju0WZAHgfEKOxMltLOz95NrrsBwerXdeiybK5EAiU3YeYp1yca/VZmgIej/sPrB+
fh1KRRnz5i+WamqcHtI2lM9drGDbY98VXZFPUpk4O7iQT+x69nfNNGbXM0EGj4bT
yS6G2BIlvnHpxFoAuGKoc5BZr/0VZAdIt8mW1g3UkTw6lODNiKC6zGtV3o7J6yiX
gAM6fwyX3WxAOzU9Z/Am8W6WJ6MWDY4vwHqy9vMW/fQlLedO/LJSsqWHPlz1CdUt
eASg8pm9NPBqDNOL1vSVa6BVeWGIJsUMkhhNCC9WlDIuhCdejFEUImQsh0tIYHau
i8pXCALJGKfKzKnA0IY8QQxuo6aI+pfnn6VPasXy7lVc0a8XHvyC+qLVjs3cUJ+5
2H7uJyMauv1vFRsgdCbZ/B+LnhXu0NRs+25ehkMSi0HRimcIQNwNWXNgMYYyZQAV
V5rc8gEOWewoK/dtlMhoeYKtXie2hCYKtQaeIZ6HbQJweaVV+Afk0D7VFKRlinJO
1j3lDWbRmZXIpBNfGwr+O/2wx+ifOXC4ZtKaHhi2bbTmWQHg3hGcZkDolYHuI447
0BGIJp6h5W44iVvBQVJamI2/u3wnNrjBSBkWiogKjfSmr+KYlyZk0xTF3a4QgAbQ
mFD0N/H6pCttxe/Op6WS03GrM9fruyq0N43T9bpK8df8o/xK+m/9I1zgYGNVSW18
bIK5nQ4KI3XeGaWvQUcRk65FDNm1Vcp2PnTr8iaQBjTdOyRulLJ8tnOnHMXz8P+U
gOmCsuoSCtXntETTaeaLGD7uiTReYii2mz0sS0pFDtcP5QSUqg9Ljzkva7ex3sgg
EGYwwgD/p9sWwKO7k/iiUYwnfbQEbKNjria1ThX5UJdyFe63QcRYfYz4M/1kmgz1
FUwAI8Exk5ImTaWKGcUu7lahcdyEfU4xRjm7f3QoKUOrOLp/69+V4szu92rgor6o
hD6O5P3bL44sMBeHadZtCLXMwS49jSl6dbR4KkxeilffkPQj0ESKTd2Di64JDSpK
gv5UXDATuVt1rQK9h93vPEQnWhE9XDmQWcgii5p2eJiGJqlLgzpXumOyB9xvVDka
klB8IGK8gTyssoi3qF7+oO6Zkq5r4BklAcX/45UQJ6RsfJAIAoAf600q19p86wXS
R87MJOxJgToGCx+m76OCXWCIH33AdQNfXuIIejCJVpdAMwh2ynsgt00hmfTIAWFw
Zm+y/THxrwWzD9TzhQTjBdpEwvEg3Xw653Vs2onSkEoSGSvrie+CfBQ9nPLkXW/q
hSqf8Ag2aca3/ZNVKE/RyurO3ce7fGzi+fntS6Z9TwcKtXx0EITaxKtVdvpV5X1E
ZeMAOa7cuN+3g34d/BggX+SsZ8YsqYkE3q5WDgMPqOcHtquQ4g4BnmuNthOttGMk
li41yhjKSrQGgmMgPzWm9xzgAl7JRpSRLaQfSw47a71wDSK5ztZqejhxyPTZkLXl
4GzXP/iDlY7BJ9tX2/U0KLoDf+LGEPxjBUoGqbiG1TynQMYIGwUNds6Rrrn0hKq4
SUZ2XRuLOVRhqgGyFiaGg+NQ8FftF2rNgTL3vjy8ZofvAq49KzHe/acbKeHAi4RO
i8/+I7BcDiDvCgHF/8kIdNEvbS9/5th4DPsNk0q5vSU9eLBsoSiwkTt9BQKqXFxk
Qh2gvafHBcA+N4rCYzR4pxgU8zYVbUS2ERb8tWxZv11gSBKA2dOJGmFs3Ppik8LW
W/3NDd/uhVRmYmifh2MlDJa+oIVoME6JcdvuMZdJiryih84nwPSt6GljZUUBK/rB
onfdqlm0dUh6NBeNQ4qoZW0bEaGtaIQC8rwmTOJGOwG/r2CmZl1v6EALtBSbIa16
PAIXJ0ryGknUjZPlv3prZtArSkw05vVoOQsK05kZHbD9k2gSJTec3mJiy1hute4I
WieWgdfinYVMUzcKDnofsuo7sq064NGVhktrWyDMseU30SwNGUyIK7PksexOQIH9
Y6UIhy7HE9cJYOk3Atfn/Uz5qGuoDfpjkf6xK5uSlbBZ00L9QuRJaSk0psRtpyb1
oL+t97AEdxEmaIvJphnVpbC6VkOTTUUd/66SLuWsy0WQVtpIgCeE/V6hCEHTR52R
gd+0kMF0J+180NpJJeOYubG45tEXhCBx6Tylu29TsAmKzcSaQFgrh6V5hPZIj0el
jw6Ww7V37r4GD5qOyIy+ftABonxHdn+HvhIOfppuEZZzJifrKAhgGCyxdJzNJ8Oz
O9kr1wZ15HryEvQ7wtP7oulgQTTnKlLM7/ZqmyExthCd2KCs8Aj+JDv2O09oIsWW
czuchVRMFOunV71GwZE3RUe5qWDhy96qkrj/pgF1nd2Oxd8WA55QQuA3D+GT+dkS
BdN9P9bTZ0PNI0ChyXhtE34B/nlrClNW4myi+k0DwH72jZI9EpEm9X3xzqTchY/G
83vEiGOojNpLxNbXX4D0EzEIZ5VrZXoQfAikRyZC1WJtrDpWP7fQFK5cn5+R7onK
B7r3PlchmmKNK970NZwA+z4ZxfiKlI7r5dNiCsXeJ7W+KzZZTQzEADh6m3aCNsF3
u+nhC0OzREmKPC0Z5jt2nMDu+0QRlclVCO5WNNa/ng/v0wBz+CVwQt9JOFIgMg3L
N6Awabv92lVt6YFVMWcXNLX1EIAAIIEnqWSqXBt1Np0gUBPCuBKiyfe0W9XYC+28
IxUMAMmttET7Q4F1+Evwvq/IrmIJqac1y+yOFTumkKGReUr660tdBcos02z+ZwC1
AraPjm35+o0Amijyg6bXjrpDGU+Hh0Pm46x9G35GL9t6UUrLf6baxJGj/1VGE+9V
JCErc7NO55dZpjwqarIkyqdAYOvpKaWHdVRTbA2Q0VeLUH9H2kqf8NICKAQwRLP4
P2ZrBeW1aEzZgEMfYHKhUQ0VUgmV+2TTeKA4O4cOK99OECBgwDZI17OvYyFrk4Lm
paz2LmdEnKPIJpOszKY0C5gpmvstQC8kPz7g43L7CHE8JAgd4xXCQ/3kCbFPaD3p
pVZiaIaes4lBgFc6E19xLzphJa4s+989KOi56HZxjiBmcgLY44TJGAm30PPxaxsz
k82u4k4eA2jOfoY1j75Ke4LvRcee67b8JThMIN0YcPPROAeuF9KSiFEAxsRURX9I
1jd8sNoWscCgGoUNoAWd5Wi1LdYykNvLKjWEoIo4A/YKJXefoxnZAQzVUdF4OHhq
ywHwSCF9qTUj9LDj08fyM2Eq8e2yFmbCnzC7dZMO3SxTkvbSw9FJXVKEAX9GLKkj
nG0vkB12CitgGvvcQ53D/BZOzZaLTfQbAzLZuC7PjTKXQjC2b7RGexhK7RiLB87p
SF2UVdU0kEQFfm+U2aodEmE4eqE5+5Lm09fSJrtPo9XUZV3+DKSF9mntMl8UGcnB
/Siw2Rkzm/HoSdXwHom9fKmRbWxpIQRbkAjvBixFlqLZwUI4muNWF06GSIMEff9m
dDvd6h8NdHaiUGkDkrEOzY0QWBrQEQticLCigZgZZpHb5NFRF8v/B+RsuE9iuk5Y
zMv3qZ2ODXD2++VhJLuYFtpjWoWGaMdDsH1H2vhdLwrcpYlu4uEJUL4fCh3yx2ar
2WS24pzeIUTgflnG59FJmNTCKkVHw4UxGA7rrylj6w9IzJasvYKmDGkjwCUAZA0m
XrMaemzMd6YvbcSO+pdbZvuhNIEiaPmKg1CqD7coDBnRkySuQd3O2soRYSPLNBCp
ckJB4cEI865/InAS/ishxv6t7eZ9djit5cOFBiWatTpiSu0v4ZXaoz5STaO+EG2l
kiU4FpgOoLYZkPJMTpghZ0KbpOkwfVPPJnRmWkUhh7rpxapWqAbDp3H6MBX3NsQ0
TfnHjl1/h2aYzAW53LZx4B/ml/zanvBl51iBcLIYsvih2BFDFCqawLElrztH0Hnx
DkKDU3dFhhlYyLvuZbqaRdSjs7J7qc4g1ksC4DTKWWpRky+oceLvLmdf9Zb7BzMA
DbEJaSHc6QSHvQxg9TgVEl8a4HtSh4RhRBeRrWlKruULj3DOaPu8jY3My1s7FmWE
HCXCtj+XnaTAaJUun+kUPM0nfPzSujpxzvUC7C2KU0i0munL5qXSsIILUdzutlim
OzKRr6JfI49bmywofrQlC3cG5Ffhf7Qeu6HOYdehfirWKdr/+aCvB1/HV+YC543N
Ac9x7YMTunws1eS7hdglm5OhJNhCkEZfn32kyhKavnIRYMzgXZCB3GwYRsWUQuZD
TAFrk5sna5RMn3VaL2l7iikDoBKeYlrvacY3l3V0K5qWpfMR3+jj+9KPpujB0Dsg
Bm9nB39wnJUMH7tVMd2GRHaN+JRVxaHXodi4Q0g3g4i/C9SHo2LptIfTxuNW664o
Rk5oq+/+9RR49bwidZQK9wSH0o9MhFMfwxFSEGPVP89HySF3Coz+cX9CziEam6+V
ZleAFPFR6mY3ZfSr89l0mYdF6grCTPMUbgxvHKOvN9YjIbLDq0BCplHjHT4FHGCM
qP/EGl11EBWrtLxBJXGpQPiRU0BXPgIdGIenbE7i/Kpy3gqHO1wlAWIBryvhP6jO
8ojeIj4DlDwegjFjDfbMSvGUl9yst9EsxgokIEq/7IDwOFuprroflHzeZ5C0a8vd
0UQNs3/bymFbt2JTFjLeJJDTPucj+OGWTHFzFoGsa6qpXntDl7TV1UQxrVacLcL0
BHoluMtYPyFBp1TPmUxSSI2oQuX2ZVi5S4Jkgy5o+4wVO+sXuO5P8K4QZNfE3C3r
4uHMgf1miRWNuxnmySeroHoW+KSaJEVu/YTvnr7OZCvgsiDcyS2OEBe344wOc5iH
lMmvNMhBkex+fNch+BstAEP4VbATepHawid+6B7q77+F38lwWTMDc8ZklHVk68al
mZDj7DwD8u7zmCfKvcWufsFEcgCMMjarJMy29vmCmEXxlsZJfI58kacw64CX+pD2
gBzCtnsADCghDVbePaRH91YX7pLfFANkTmTVL6peqy2nVjlRJ5V5aLg+fNKKxL6l
3GRc+PZvEEnkpRGEftBQbhom3V3cFvtsmWc+S9SA8tiwE2glQgCOs4ag2u0Svs4W
MrnM0c6O3q9EYsejTfCeDqSEkaXmT4e8QaCzA/ZWZsrhlQu0Sl2K74w74oCvGXJv
A+xmAJhW6DD09XN07ppSC2GhwDXd9rO6W8qTPQuISHXyM4Tsb0TbrFz/4WV/Gm10
DsydW5uvATes9X0pihNgF32Au2JyGsJObVYYj/QsvYNfW/JYXzC1Hu3viW321vzP
4bHi4YDNuxmCUJOBw/BsREj9Z0+I2aaxnZ9D9vS1j1W8kWZzi8G4WzcAqDd6ms5+
WVw5VwEI4UESbBq7/uHQLQ05Qz7gSI1Ve1DECbhgS1WhPaLzefAnZpm2VA+n6ldY
g6Fige0hnjqn2VwjKK4b5QNsKGAj8i8z9fALrcRgPJNeW3G7GwpUA0RlDvwAUOAT
3QpUmyYivVIOKdFTXxIu9YkY2PzZPtz6J8zT7FrCqIGsqhQn5lwHqUJUvqwXCQLY
Tqm9yTPOX1u/lWS02S/LJYoZms2MyeV2Ydwu4LZH0obJRRIHYouhRxyNSJTgsaGp
Nw8AmLHPhmWMwimQYNFmW0brvirits2D8ykrCBuR5vsfgenvxImnsPiuo7aI3gco
4JnQreumGiFPKOLc0U0XuGE/V3OWAYGucZ4PxGpp9NGtm6c4e3kCpDB+x9fP/BOR
3Zps4C2LrOjGnbp3lvuF1mef6v0/8W2e9+g9mNRPFM2sz3UwSWsBwbc1U8tXypcv
KcJsQbhdMha5onzZieJXF4w6cdRaY/hWmR+Ps7tfhPEjVoAhgWD5ijHw33Y1W/Ct
HBCRILT3C3kcbY0imYcUEG66lo2isksk0iFHo3ELzAHXzUhc1/C68/sK7mRexMMe
X3tjIkSNA/avBQ11EjUAcVnaFWnLVI/MczX9/ls1mr3EN1V3FlK7WoCiaWWFBM9l
N+AcF1g0u6hxc7MH7t6I0AFsMmRksApP6ZY0KlLKaiNuz/wgBtS0oygSx/TNrE5z
qlepI/EnzxnXqfo30EYmScCKPh1p3ZsQ4x8lhqVex7XCwazeL81EakiatBybRI9k
W6K9eGV3GTDcu6pHBGi98v429G5+47Oilrj+FAaO3jijhTYvHDtTtHHGqQ5HMsaM
BJj9ZsqNk7KrliV4Df9/nAnL3mkP56FuwIbybBXFisoeD6mtB4kYxMFHTVJ/wCCj
RybNKwSAOj6yZU0wW4twQRR2vhmU5jJg0aTcAQVCzPzzKcNJDSb78EHHdaFV+Jiz
KDuN4AwQNT+dwdFFzoXsJX93mtHuNGJF3F3PZ9ZdOLSYaoO5I8uPoxJ6wD2iM8L/
NNC8NPRoWADJIA5btf3u/MKYUIOOe5dQdVVsprkEgleI7SaOtrrBFRnBE/fFkTwT
80LGyV48tg0rUygqnO2PZf5vXZj+K9S3S5zyY14OCthGoEcQCIx+BbaHeSuK/sbI
NQBBfcy4pWB6qHcSKtJP959pI8doaYC3fjXiVX+m6XMrPQYnew+4Of44No2n88br
p5RjhJ+E/rFOuajq+w6d1c4SzCQW8ikaid1/pdeduCe3t7gvavudJlJ2SOSNFPD8
CVo8Pvwx0KWy+zS8jloP76kfoXh/eTD8iCpevS0HLrkbobdSzzLltqQeVECRjXH0
3onkVQskrTLevNRhtzKoHp54nHOlBKZgDacVuYh4mFIEvgDI8oQrcz30BeKA1xE+
v63ABoiJFLz15/qtrbEDTZek7rRTLp8d376b2kFCzIlEHsqZkgRc+vVCsY/CdTiI
sqhfkH4kn0d5EgLzVKWh/mwS5NoVf3d3e0fWfPVF0pNxL3OqtLs4m7K3RJJmzDC3
JdZDVYKu+lS1V40yVbnbJXldnGZtIdTdhBJHHExiHTkXmfeNnD4Rmo2/YOjBWqma
hkVz3AVMpci7/5HzLQLhOEVmM2WUarn+2u5oXr56YhvbGxF9ZN9wYMH175GL0xHl
xrqELx4OfBBABwplzCoyttfeuglwb8fuCKQKt7xKUTkl1fPl38DcNL62zuEpnwkH
M4HnmMa9sK6lOoDoEtQkwd4fB8BFPtwhY2ADGk1yeyCcoi56c7DrwIO6VvEuqqNr
sNxv4VIEk/Pbb4YXhid9U6LUM/AuehjxisZJQRCrXEXXqY0bn+mI7aMGWa4ARSFu
5BECh3KD+3IeArZgcl562ieBfIPGWcwR0JKk2NJnpxZCPjpgENvENXYpvu1WYAK+
LpahXx5OsTXD60C0dI4gXUnudTXfn4BtFhi+OmC2O7evhFBgx4f0eNvkoM6kb1SO
n9UBoCQfrq3QDHKY/TcUeZ0vJ38+PZ7c5WdqhT0oJKWjQHyljPWSiDbCsE0pJy1P
4yD9n4B78vwbWvx8OdsCByK1tt4lbb1c89JKLIeYf7S5xE+YyQXXSTI/TkkEIKyj
1BVoJ9iH1YVu6maVB1E6lOA2cvp4zTadn/BvLyNBkBV7sNZ+ML66vyX1rtGkW9b8
kEbpkORxAl78yOtoEDz02Jzj8wCJtPKlordyNDTUrNje4dJ5QCs3K4qBYYAJKSMi
IPQsqVDmIDMsBeu1PKwaVs3arpjnFWjfdXLMXMPj2zhgmo3W2BF6rkWSXjBRt150
8d0/XZ6avd2bFxdx2d9aEiiv0WhHKg0vLgQ9mQY5LsLGU6svH37Mk6d++UPQg/AU
1vb0EBma28jw94pT7YhiDWJs6Yob5V/Yhbtv9wZNEDuC2GC9c3D8og3HLa+hzVsd
EOhp4N7CkF7GOHMmmUAnZUylAFCwzQVvCsgtzQJqwygmecZpHeteCkIgJgOYymk/
vDS2nJUjh1xatOd8TRTYthCm0SGAVXLpMAusHN64r8b881fg8Hv65NIkEWbC4te5
ANiWRiw3mWTJhxamIhJXaXAQ30OJKl+FHB0bXE1U6ZQP7XgGIU8GKj3JDKywlwpm
5cOnpd23+SpVZPYV1ubfrx18qQzzft44PqeGMfOIsaLlzvCeKpJLVV85nIzRmsuw
2kVtB7fWboPkVFeNtJeFg+WvEM6NLuWN95YgxVqsgiEsyW7m4RMTB76U/sbv7aDP
Qukdc4YtgtCKHFQKozdY9GPOm4E8kbRlDiESYW5KxiGnULJLN1pKwnxUBYhdqaQ1
optwsRfobfB3TJBd1/JEozgifFOs2EWSxzRj8nNoAUFwcNQuD/aXFCKBU/PTMdHb
rZUcwBXfSGj57E7Xg3tu7MaJ0aHyO3zJ8/AA4zDEtT680kou09c9H1+dNw0/1vT0
GDS6IZ8K6biMNVoyj0gOVbySySPoTrlQzvyyCrtzWKV8eFPKDUmHClzgCifaaxOg
Wz13xVnlAWHetXx1ZpzwQ0mwPjF7x0AWfzP0ABBMlidiOP2GA7EUc9+9MNF2wCtp
25KZANV0MeQlCCmz2vpZWT6M7dlvkTTw/jIOIp6S8JuxVIRw5MGfTNtrw36vsh8/
UxTElmnBCjOlFPArGnfm1a7ZMels7AXUIhPbb6n7cRcABb5dAG45fClNI5TgJxQn
t8HyrrGvnCR4yK8XSqoWI/W6cnE0UsFHZa2kQzlei5gdmG4tfRgAFVYzXzEBIDsV
sR5f+3NTEoUvJSgi8otni2b3P4VYxgtFpoUyYQ5vPumlGtg2Q4jHDxiGkUbPhz9j
NM2DhuZWiI047SdW5LcQYpo7of7+Hvk+vGx+5dNdteshZu+TZgBZYhX7tX7kaq0D
XK2bd0NKtRSjOfkp26LqFWSPNq3iSr74SPRlntozEj7Zf0cnTsN52bU24dIWgrMT
tAgoA1zstNxObGIXHHRknA+H32o2emjIw9AcF34uCuUVVyNQOcbzZ7x6UnYwDdRc
4eCwuFhgdSr+Lth6Gtz/atPT71YOmj/Joqs2mYkXhd3Sxc635XYmk7ORs7Moccfh
su0Kjp3SG2wazywgy9+tXiKmxZAZ5G6p0QNXypRzyTO9Wir4RkssuuAgQB1lv5u8
3tGEW9VVdWi8weSuldcJBiAn90qOdRoAbVzdcXBYyACUBTCXQO1fORnUWUwaFflf
/gpsD805GUZQr3x9acKbt0V/z/d49UpFfEHSEqXJAfyKf0FqTzRKtlq6ATA1nJyz
UKYMJt+5BSe+q8OcnEanmHFinoXmwfb/ErKbzMpO9JlTBPjuXO8dPJD7qfbFScrj
oGIk9TtsJ1oWpArCKBlmodA9sR4rh2j5Vd6ZUOQ7fQzarBzXD6kE6UplNiWb9ZWg
ZLVv4NkV7SrvBzcKTvtcSy8HkPxO54QoY4S7q/jPbJWUCNaltYZcN1IwaMgR3DLW
ynZNXtvm/r9CtzD85GG0j0tQ1QMiJKUO5JVh+g7ZLkmaqfkdINGrHk2EhfpLASU4
BpoVq3+OMn1ukGwftKEUozvGtH8VY9gCR+ZuWMmiM6w4HY7dBFuETRzdDNnu/iRm
Oo09riBjJTKy1Dia39AtDj4ituvyMYnrw4Np/E57zh9+Ll6kB4+wdgzwd86u1TMO
RWuZNxR6SYIdLOTTkSxRsoKFo1hD9ii6P4OhcfyJUQ3Lj54ZX+QSf1JlkM3SOJSr
nBOvbTLKEfmk0qPGKoOcehey1oJ7NIZ0rYDsVc3Igcdil+CqKNCr08YXEsx5QWdp
iaWMw8O3y0Sj8M9d0KHK4LU4vrbKI8dPjfZAQ8gCj1SldZsBEWwEq4QgLX3VijOi
C9nmUexue8jUhV2A9QPq8IW0Dj0D1k04yMpBGPMYnm5/Yt9LfHCEWMh+gU+zoZKZ
rO42YH9Wr+8ovPLhyLV7Y/3ixiUlLtXtRC/LrXzaedi+5+pW484w1tg/rEOrnWU+
KrPZogFRHblmRGaCWHmYsTVJsRwznT2EOmlaMzUadC5i7IIxUn7oOKqsxwQ/HzxX
PZ7y/PIlgb0VOG+satRbIspnKat+ddKL19yewJ7bUH8ZkZNJDMxaxX7JykFnriOa
NnfmkBqsQpn+wzS2A1XUpwyn/WktXw5ivMdaqbTfb3Wxm3rECZwbGW2awZrAGafS
I99S3rGJjnjQ8SclZEYivmyA/6bDGfznHgOOviK/1GRlnhNR3V6Nnh0/kgUVlOr2
EQJyvuwhGwIgBMSMGMakY5j1DJwsgNxzauGrejxoUubBLb1HT/vNAFA3Cx9YTaMR
/8/ZOf5bOjTdaI6QX846kvwxlp7Ck8EUQto8fGHveS62/eQzO6gSmhfYDe0tbCnL
IfhSJzhWVa4IX1oG2yzNpChIJOKJtkDlZ4v4B1YsL7L2i1wL12PjTz7E5EMq5m49
D4twuJqFf4HB2PbYk4l4fkcELexYJDmNSP7wZGZJ4YB35ZB95XI9qkmINLxOPBs4
7DaqI1YN7eUfSN4JG0vdqzRQSlvb+n+4JIyioLSw1pY6SdJyv4s6wjdFG6cSOLU+
En1Vw/FyoAbgbszToUKPnpNg/b3BChuBvNq4hdsqyURe7SxV7O/sMvny9zCDGVDw
h99H+nQA1iXBf2f/iBvcIvRGJbcDfyEsoM8x/UiaiNzg6BqtA/wDV2qnth8ISKR0
N9kjA1Gma3ihgjrU/CzZyd0xD7TZnaF4gtIX+/tifzYbjwkJu47jwYdUMAB6qN35
/VlFiPIdwuIZewz9q7Jkftggq2XbPERYq4YTVyYbIxthGFYWLgnIQ2MhZjx/yMaB
5aOsq8V8Lu9p2OCmyxSLZ1zbeSAa9RtIA+yA5QwBN9BV1K0QS2pMmH0fRrboDwjO
vk8+igiVCmXyLtLDy6wfFi3VkTxmsIpIuyCffVt6W3D5sOiRPGfQQAFXDNH29UZT
fMxygFxHvYGWq9dlwIDXQAstW+T33yWR47At+g1EX0LA4DcgClybiCtkGx7OdtHY
QQnmnPGgSIoGnDEZmY0G3qUsbp13Tw6uD3rjVTgJsz+UpEbwb9EOUxs2DMUQrEwK
FvayCOJcPPTpgdj0iDxpT0wTpYPyNTHV0TrAfYXdPj5Q30JV/shgKisWgTc+4m3h
1vVBpBrxEjrMVgVCgRLOAQ6UltYEn6BwWInzFKmbgGl5hUs+4ZfD1K8C4njfrksx
HAMMPR10p83pH6BLL2WwuZcP05UnOvvUMzpcjgg3FMiHvCdQQfOtaWBlGuhMtYg+
Q05WTrlIFR4CzErlM37lvIKamLe/sN1Pjm1dSbBnQAkS/f/XBvSw+oZnlSnTyWCN
cg/s2jtnYGN4yq8CTOoAgmia9quVuStUSW8rQkDHXq332H3qW8hfl9xrcXGkgNVI
hpNv+/nDZms5yiyMYwVx//fjQvJhpH4SEmkXRzkC8l7JQaVmkalKie+AE3k8F+u6
wP7P8WilWa2dMCNinT7KfNftJOs5wDg4Nhl928QsUQjwWaeavMXd4xKk1ZhuyEo3
Xt1qhcJTD5H3qcj6TzWOzK2CF2W9wcCaoez7n85MJt76sYB6d9jm9Ddjpx8P1I8p
rs0a1mOxaUF0HZK+tX3BLixz0JH4sM/58a6VRlR/hsX2sTOHKE62POcpk8bAosZr
+pPpxBl0677DA1br219VSiZj+kro93Sj6Gb60p/6MBzWsrA+6SAKxW9T4Hr6x+vG
8nhp/2+IZfXoGDqyvNo7OPxBDotFDdsyReoV/KZV3nrsvVSPIuiSKzrQsM33zVc/
gcKpxW3QErf8SLkJMLyF19qykR4CSHD06oTqOMdHP0J8Ui0R6osvrR5Dfz2eJAvk
8OFe5pYCWpDhUsGAtFXjqnqthMKMAh540JNZCSn16Lpum3aKsPsT9I8RLxcC1dU3
YDx84p61zFN00RDSUg+2YuYxTWnYrwcksXbKKaHnJWQUQ5JhTUSQDrPvevtrPtII
rTp/YYMt2boNZFKHKa0zNM5GohDc5QaWArfickWgC6wE3o5YlQJO3SR5NLklYgdl
njIblIm4SWpKYAc+S4H1JJgmHS+iILBrRKZf157bUCRXK5L1gSFhbhHiCBYae+yO
1DI/jrvRnZ9/JcMRnDaGyJrCa0B0jjBbs4jKRdav0TKzmMgK5oLzd3EofsgQqxWt
4EmYkSU6AGb+vmLbbmwf4LPA+3FiiWHFvfY+tEhI9+ZiLHIUEEfbqsc3D97ra/mU
7SN8eswooMe1evP6prNATcoVJoBgWqVbW+ehcU8PrFYH9RzXA3RX7VIxARtL/qlM
nxCRdkcKGP8hTB6ddHACnFOYcCsD2rBjqzZ/wtEb1fBWweRw2+Hf256JAsis4e+A
f24TGZhYby9j145fRRS5B1dOcXUI6+h10U3AJjZ9PLuPiRGW6Bkt7xLILdf8brE9
XYilgF+eI8Wt42+5UCsnj6gLNKxnbRZFnPQYrieWaBw5UlXywcKzdJaa846MixAT
CM1qxxtQyXogbBTdBJLj3MbS6Uw7fhN0XbJyRPfkxfWNvbqUFpuCDgMoGSEXtae0
uNleIyjwYX3ZWWpeL/Je2xvx6ReolmOotRKdyTzQ+BAzdnBBVhuXaEzg+fETCu8C
2bPTBiMqueJcL3GHt+o/3wWqv18UCt5sC/d+aJrp0RL1ERnqG9qUpJM1zSBT0QKr
wh0y4+c8ltZKvwj51IhUoOAtiBYHKr957dViKoe89znWKht78OFR13JGAl612Phq
Qn1RCQqRg5/WSCFUCSR2t2dNspxlOQy3LGU43AejOGAMMl0ZRv2ibR9M0IZuoW43
OUhxkfM7O3uEmZTrIrESuFA16j8TzGzxHj7Un4W/LH6M8EHXXdXK23HV5WdRq78j
Lk+pbYYUpMSz2gt4BihpFRtsVUyu8bCJlkU6rK65Ij4rPM4iBagF8gPiMzQEtAHA
j5j+J5OP0bd3Due4KbDyCf+BtvX9ftXoCph2MSp6VG8j9SLgwiV5FwAViZx9ldgT
ZoVgMxGhNhuJYuwtatImOl1AU43kXKuBH5j6kWqRHzr2jC4lgiMnOykhrzoThqAl
V43+9ylNvnaIr8kDvIjuVAHPTuzlOok81eLYqTbdUoH1TUPH81oOci9mHHQ9fC5+
Z98jBvlf29DprqYpbcGJ0DgNRxr37bAD+UekCxZVjdi4HN+T1tbqPlv6UnKavrjV
809wb51mkapjrg28RLzYCcASo1CEHqsnAA1ItWZ9UnF/O6zZCI0mdMDQkHCUZiv3
rFN/FXKBN00tJ/17tWQeAVxMAATl3dz98barvqCDIJitPRl7ViuP+hjicYtkVXCK
sxaIjCZVhUxNpRMNPwR5v24Qx90dkbaaS1IEz71yLc+RrIkjK1isNV6PmHWKWju/
0zHcMXmZ0jXaB5ZJDjDuummIeWPmmdL86au/5YssYr5vkgPwJNQeObtyhe1O/dyw
8JBasO4JlZYjNqdW+ns1TDLtr5vaFUhS5e8x8rOTRLniTp6W1geYmfqQBSvJsOCo
6aReAwLJpLLyS/WhJJ1tlBUemvjX52F87Ddv2Dty2Q0QKKGdTR1KpzfFgkqiY1wl
A/qWo4aXQKMIHldcnQFovmBqgx5Ck4hBrg0rNBO1zqFByRY486Jlso2IZ3nhgaCm
bZa/VqHI0ri/8dtCOhNYZZcIQp8L4G+hwFE8csmBTB0E5fg1iqAokX3cGFeu68rf
hHU2q2xAfOzdFaZzVBavou2FipQc6bzv+L6ypmsDm4XH+8YTMDRSAGMBc78hn8QF
Hk1PR63J+in6u4OT47nd+5OBX9Gm+tphuF16dy1rqC5BO6UOCzOqgU1ELdHtbByj
TE10FO9AQYmBVWfvFYXSKhQB6H7oikJESz/l/9rpJ3MkGG2SUClvRgl9CJLoZ9m5
OcLIvXHXanHk2ugSEuqPvM3VXTXSo8VPu92s9aKz0+GLWb+jER7KkIEbZaA8no+j
Ww/3Nms/HHHXheuT6yIqbIvKQUZmBlHes1h7CnZXCebU12LhX+XwHXV97U+bnhIf
9iHHvSkb13YFbAbMwIbc14sopAtJJUqCN2hIhxqPCNnDKQ2spDmDtH4axI7EonCW
EyrBZICEpEeI+1ZOu/yQRRFlULvq+zwvTHmzUHaLwT4J3eZQMbojOVcTK9w+QNZf
Qz3gbZkwh77r24Pkc+1LkNAl4+n0EDQ395GhDqWYBS5YEx43W8ZRpcvpokXzW0Cn
cnU238su1s8agn/FN9oz2sspZ1q0RXjt/LtjseuM7Jg/zW7XJ8UsPnsTJQ8JF/n4
3V8eqI69lAoVqxPTHJIAz4wlwGGLFHaZrhl4/13qqeFjCQeCVzAmcc8O4vAgGZMw
uV+iXHVRtjHMUWVWrRq5/2E1ndeptwr5VERgjEjUuYiIO03/FAYFHZRLrFUmAbKW
4IGw7VEPVGMZIBBpNEY7+AVsKF6z7OweqZbvznQV+5WKBqazFkNAHswTPHX2Vj99
PA/ostD53DBBAzKDsf9CTmjuT4MlGKm0gv83sgX5PGYWzRTGyqdg0xYRO0JyEzDv
BY8YL3MwKRzXgxBa5ZbrKovHH9Q4c1ztckwzMx73eAE/kLldylRVNAUpa+fIJRIY
XAJGLnnGmZhUDhMyNabmb26tdeGU+HRTfljzE08gNrhCVB3H9mBD7x13EjdrpqOW
oQXcRfimvt00s7OtHZS3GJaqbhUgra7k4k5k9wP19YrdlA6/r4XOQQSaL/scgrJa
y1FvgBDwJo/oSAc1iFbVkiwR8fvdT94jMxUISR3FloN0tTcTQwmu+TL4JjH8cDsP
F3P9fMa+4srmZNDywCXp6eJ1PQTIUJwLUWMuSNxDqoBaV+/n0vlLwo991mLv+s0t
Td+RN5DXBlw7yK7lc1M0drrqyJR/hxpYO5KMCtTV2pLveozpzJKuc/X2tzdSc6Ol
f5D62akiwK9yjQtB9rUH4X1P4bGiXDYXHOs3G9eniavte0hVPkufBCSryhI352NP
0ZylG4Zfpreg7wTF6xQHgOKbj2Y3qrfIo1loyic7K6STLAV2Ob0VM8KyUZQutgbn
Qvew/bMldVYgWPooNUawTNeLHd3MXDbuhXH5arXi/WEHkeVRCAsifpXSsUnqARzj
4dpDBiBy60nGCohu7lDsd3QYzdmMhcC/Kh0/ptrBiqvk552TWxHIBJEX69AUU8IR
EGFx7jrBt0VreGKjZZOPzGenUtjh1K6RWsismovU0DcWn2t8iijZDQNLSgyHUWw/
okASNpGQquRsDad1sgdDuaLLGnXekgjGxXA08Ug+SQeGwJjozcwA95duRoXw5j00
wglzwNlgJYu85MW446yAXfewvOmVlau1cPWChe/aplPg2iZjnf+ruVWZgJ71q6NQ
pL55kkrLq4ohcwqFGGm98LcSRgfUcbbzjA0c07ooMaoRbNBFm3jcpNuoRYVQ7C5x
SPbZdlOwSaILSqqi3Lzr2STOjyrfl21n/zsfKzcWLv57xqC0ZWquMIb6QqlgTaRx
AeDVoIWbZ1FnRYbf7OK1jvJ+1LkKH7XTu35qX24Svf8BuP2FnXbBrujlVZk/vytl
lQK+7ugGDrtO3CnuF3zFopxpVXMoweDG9405dGBizZYJox2M3CpS2d3xfqb8fwcP
U8WUhZmiOeBHReR+vHLNeMbpy9sGJgjeUdiiMJ0yfE0oJyaY4SD7shy8xNRPDgAI
+yLJl0r4Sr7KHTxA9njrro/+DL1tEuFA/6gpNRGbWpK97tFz8svg9tYrvoAe/MiK
t7EYyIxWqIqdwBvQmsJ0o2iZF7+xy6qkBKHv7H0zlL8AhA/6LzbIVlU/G/6ok8rV
ABnKLf2JCvUmGK4MQuINu5MMF0VK+SnSnvoQ8lcIAgOcf6JxRK1HlFmkMdxC52Fd
PAJkBUpT9D0Gq66O+74m2M9R8GvlnQBxE0bM5y1EImcEdHUVR4Jd8txpekS3CW9v
BGEfufhfd83BWH3em2dojJ/gihFQZjcswfpjLHg223HtgH8zJFlHQqxATfCCcamT
H1I/vtF5zPhEnVwy/gDmI7tZIHTzpUlAYVI1o2PYqfRELdx9/IDunH3po+bXsbVQ
A0xprm0QuK8wyCtWd/se99Bc/VyQiZEtEwChJpJh3ojL8yEvnLTkKlMkcnwRc4SY
ai2osyKAZ33e+ByPv/xyWrhK9nCTWhRz6Sklymc+AR4r/zHHYXqQ/hD8BWB6luvl
e0Y+N6PpXWtlbwC2eoSQaogRsa3MDLy0+pg0QdZ2Q5UKyUMBWreVv8JveKHBdMMJ
SW8iPrC1jTqtzznr0fOTyR0kdKUoqWxPNNdskGXJKwKguOih2n/BJ/r4T/ffpvkH
rKThSHjJ0ST7LUu79SdPT0R+qSdPTgLegbqEEyg52W9BtLZMTkj0/csW4qREYysD
GNojWInOMAVc10l4cbzLdCjdMMsCR/eWuRQ/OgqX7y/s1fmc3UIZfwWRl3BZayjP
4MnaaqZNhifA/3NG9ZRT3lbwxPW3y7FSYM1Mn5ciQsMT1m51m4rGwSZkzdlxkh+O
/EAJq4OdZj6HQC/wkHUrwwumBr83rgOINVCQAwIttWfBvQQmjJ34Ax9aEMrMzV/o
U5r+cmYmWVjaeC8atkhkKGje8DJ0T/tb7csftUgRKSeqC9nNLamDWmh11HhmeAA3
q0HTd1ARNjUINjgKE10EPFFAQh91xwpnHA7YunEq3dTkP/KEfrK5Ge9gJDJgMpIZ
LHdsM3KZYcUN6y6Tzx0b0XgBvulsfpLskB2+slKXcXR99IHc3couZf7V/S+0xcV9
k58MUNbUiUCmTG5NSKc2jSCfIaZFUa7quUtw75Ac2pjqLll9oSCUTI6+0eUDFIui
8LQLPzX1Sc8OWFD5/ZD0qFf6HGlprlAiaH64fKN66z35OaKJ3kzyfRKYb1BXDAQE
JyPXz6+WQ0EegkfssbT6sb1WDP64htWsd6YI5618TQ9Ramzy4otslRIYEF9CB6vD
/MPhpZiEg/E9RIXruaSYiw/5xcqhYUTxzDX9m4tcT0KqFsjW5E/wNSUYUEYMZDHF
39iBAdMcJAkUbFttV9zBPka7vI7jj8y4Rl9QdMMm2blGF9V7vAJD+7ReuorC7A+9
7jYbnNMkWjTxHMzIIsnvGayyfCeE5OtSW9kYr//ScpwH3McFR9KCEH2s9zgaBQWF
HzUBNZ52ci4G8KSjGqhWMRpyCVyN4ZhUKADr1QYtjU9JDotkSGoWYIX3LByamNrX
fCKfhyd5vugeGo3jjUUTySo3UZp8snP+gHgoYUeE7bkQHYC+ne0vIlbHyx3ZpCCR
Sac9uYVF4gq0wTvyBJ1rCh/UKyzqStzTa49j9Dm7GPplHC4CjXAh5h76gJxBL+Ja
wLa/bqfbs8k33vCq7QOJRfbc6PTOJ/ClkO4KV6B14VouDIFrH33UpJBfVu7t2e3M
T2wfzWE1N9Ov4S2tefd7KMMhNqqLVcUheHWECXQP//aH4rX3Twe41JUCpJkHXcKy
OQLgpsnm0jU65I6PR8Ou2HywHxUxZy3KwYT5P1CoeGVLN0b2nktMwl57SyqOxbBT
h+ZXEBo0gtssdkOsEFlO/9ucY07H+st2lUD3dhovx4sAKmGOosCXfuREtcBSZ81U
IhfLghWtqxodOrRdNtW7CGQJf6lFMc7pDjCJTqegaXECve+TnTqwhBAaHt1ido/z
39eT4rQRfJlASJ671ly+v2UMsdEjITDwVYEMsazHjxMgKMEnQqSSHVriZKCmhyX/
LEgtJoPOvjlX2F4J6bvbdn5M+RGkdxvrzn9R7f7wFcC+zo3Zy7So4PCfB9W8RFA1
q/Du/jfBThIBVFpkBJFc9qLLwbenPvJgCHKDTF3ya+cTcgP/JAuWDOZ7c87D9Pif
/EFt93S4xOP4mu1//gk36aCOHBbnrk2Ol7KboFyxSmAaPWZGWclhA7c7jvchqL/X
EH8WULFFkVrY01yjMjsJDtnfVi6L4KJAgZ7CjWQH+vTQ2qH4Wsbz9TYEyWJOpvO4
w5tFCd2nm5628gSiRoM+/WDonwx2dILVewsSrgrdPJaFmHpMCQkioRDNDUQrG/Dr
L/KZMPAdn9Ukq+LRS+DqMLAM8gUfN1mZN0oKqPR2dsaaopILaSSjyZpSkOn0nids
iNikrPt2dTcVuHdTAamgDiB/RE7C+121qE4z5Imb01QPc3g5dILTmTADvSbq4od6
eqx5FV6lvHTnhXxCq38SFCYVfu3oJq2dUu+cM7mFuzoQmG/uQNCxJaJSu4lrOrtz
SP+8pmotoMkEspUX4fMZ0qKU6y2BC9OtBsYl9YcACR/+jl1t+cne2govEUaUsmw2
dJci6QV0aN0k+blDud2Hq9gle6bgY2yzWujtCoph0t3gjDYvfsfbiAYwZxzVjOu7
/e9oOdxDfPOeTJ0WjhKXdXsO4U55Thbv6E2jZ6lmAlaPytftSYGRwVdX9C7ZTTx4
0XJeYMhq1i2eZKQ4eMmY7oPA0LKIdR5Is1IazC5e3mFwmovvNP/KPndL9iNURtJi
ErUI6jbjUo8tP4++kpOsXQ4H2K+LCyjxQFvyD1FJ1z2b9su8SphruzAI54oROZXh
U5K4pWvIRgdY29Xbbpub7b8yg7DbOLFqTZSbvi+sgzrRWWL8pe9p2bVFULt3TgR1
oetHziWTXYYzZFbcHeGypZfwTRdbF1HW4fre+cbJsaUUqja0EqqajuP9dlOquU9T
7KIVvrlC9ni5JiqEfLib53xdqN8Am1hCDICf936/IYxbTLOjiYXY15CzZZ2m2iQe
zTEp4NHkFP1ZM+HsmHgcUa79dLQVnIQjEJXYjVxs35DkOkSai5IynbwRjV0/rz32
PuldjnIJ5cw0iF/fxZBiSoLC5n0m0cEE7Xwj1MZ2oi0sVVKG2pejjxi6LnvtPhy5
/WrE8t8XaufqkJ3vw576Id0feCP8TbnJWZ+YWk5w/E/ASCebeHWtLY5YBdcmMQq9
h1f1E9R0CYweltKy17aHIvGTWPlNBUPH3pi5+M7rAEbG3sXPj4dhhbBFajt9tFpU
7fXcNBxHjG1f6603GxE1xG7kBWgwlqzqBHObcURf/fVgUbwahUAgEavcY56jqWr/
IKLraJm4cc/Iww5VnMb3qDS/61RdsiZGtTLKOBXL4ccGxL9om8Ruv9lI6Pp96yGP
8aK03bRukcowEhvhFo2jW6I6qYpBo0cO6DN6mVpMiITt8CkOQf7NFqMjHSOGshD+
tK0tMl/jUil6j2/OgQHqIknANvKkAUYXnlzIrFyzKm+ChzfsoEks6DnS8PFFxqcH
xzJ47d+ZVabr9LkjZ2K+mAiO2xAnRu9C/KoQzj/xqpEsmQp28jTDDWDRyth7GT6s
sLEyl0VL0IdIhYLzzmRNR9b/kqNxMv/+Xug2c3aiHZ83sMxMQLwmHOogdkQ26/yG
UxUKVII7Ia4XZfjz2bb4gKwzIDZUXHu98BtWwraFhM7ZdqWvejN4qUdBykcMznuS
vMunsNVDQPoOE8Bpe6ocsJ60YCP+5KHGx4l3bJ2MQwSa5xJdjNvOwykNIpARTu1i
S2wSfQ0pHVWoV4poQoki+lWN7Usw4sPrGF79Ls2gpOmLdXHZg9Fdv56ctH4DPvK8
qoNofODlDifiNIOZyLfUKix1nrIHGHTbNwjjf8tz1zY1S1oRWSUHmIhx/6vGVWcU
nUvO5d/4i4jCpPLSNBoDphnY8CUEgmlmVgig9xyl7m1cGXbHRFfZAN2Ri/sEXs2a
jsKSKXyW6UiN4Q5FhCcqLLl2KkVyY6Q0spOSJskDpxWBZSh2xtmj+/sbFimNeAo7
WAuwIG00p8St40ckjbOmpoSA474aJRqZueCFGr9Z/RVCzDcpThC9gpGhgtSWZK13
F0y5VLjsaR6z0enkEKF1od/stmRmwwWvjAOjsHwnyiCs59FVtUDh8bDZabWYvI8Q
+LLS7iKVSUvu4dzAjtPKgLca5lmxvDxgLtS4WtPa3vNthKwxw+O+R8IqNE+Djx2k
IJmZZvcdwVwliJ2mYcrMkWZY98QZB0JV9dcIXIYfRmi3cljVojctmUDX1ckKc3Ka
pJvUadJGYUaOVtsQq+NDG5J0ESQGmKUhOxFQNyVklfx0okjAfL0jYIpRbv4gao6e
2x8dw4FSxoLEO+qH+LIRhmrY/qnSNTMufarxJFS2L2XCcroCRGshNWHEHRBucaKj
7EmPcapVDL4xUrmLT1RdZLmdUtiv+9pOumPH1KIW7MkXEW5vlYGBUEMzkXgCEfdU
0pBv5m7wBlqTkLFSllmhpC5DtIQ6Z6bLiOQyQmYM3aiCOVIlMRlVon8DE3g3huYu
9AuxipGzHzROlyzSvazOze8gEUzeN98rjg7HBRXCMVqGU/F34qEJCe+eBN215xjy
XAYV3V6mWgmQlowtkZht+UuM8bSAaS36oEzqMWK/Oa+vOCILiPCRgI3pp0EJ9RWX
nLqbIYkzcZ1wD41weTAAHpKz5Hvr9bSYNldc+1Lzx5uaeBKcvyCx3CW5nXNU9wPm
1s5P0pPrwgi7B0JLE+rDr8uTOsJQR/N7JkAFt3YXtIL3CvFbsAyf8FuMBtWVGDqZ
/mOo6IjDE+27OUtv9qT2A5+9QNbzi4EituRZrtwZpGrckrrOn7ZkCE49k6iXFzMr
P2v8LO51+NOH3GvF2kTS5vC0koLKHrkxd4ff0vHKJj9IAZQkvGqkMzW8IuuW1sFd
y7RsgqTh+ZfKUy3gpyrX9aDbN5AekhnIkhI8WETJKaXto+3fIWRrMBkmjI/OOgds
AKophrZg3EYNmXjPUCa2hLwA/p+1k09K0p6XPTBcs8sLKxSfghjOLg3ll2LGfHHW
i7h1N/nlGpelRNB1ML/tod2WmyWLxogiiLoDHNwgqWsg6AzJx7WStT5oALOuJhx2
8ri/NNVIMSG0BVu8GA72ykf9pqv+yPn4Ee1NDxdl9ASQbrZtzam37JAMIcEykNY/
QqPjcKXdFFvnjpJSSsBNqFJS1/zceXEC/6ROhXYHK3r75bQoNmYPUW09EhKlogxW
z4t6HdfE8mTqj9BUCyHGYp9U63cnOF88OuyCPr796GF7YpQDbsgqkBDb30iEMIwL
dQEgkeZ83XmwRq3UU9pqGHG0OwA9eQz9eDQ2xk6KWgis2pTVbtRd8N7sXLqhUjk2
DZh7ssrRDYtqndGdaMcCX0BZgwBTFuB3Flbh2XnG31hsaFD5FSoqP+7kzW1ufLUz
tlgiFd7Tw3GiRnc06J0iPwaS7DtpFwJyhFrwD71qfmvPKjYic9XoQdDincD/xCO9
lqg5Kp/3/8oEjPYVNn/xZNo4TqDqCyZGuHbrO9CjFg25W4wT2hEq+uYQh/zkHWLP
BgcR9nEnVd20IBeqZcxH7Qld1inQcxrSWPvmFuahKXeHUZu0RwkFn1xA4O1odhGX
s7fstj3JIfaz2ToQqOkL9eWnuaOi+i81Z5NxoN9W0gWJP3/xwYqtPBx2peOIUgMz
cWwaReL+5wBSq8rAALX5mYtWtvwJ/zmanFP3+v+iZR/ihFrq0kvecKfOZr+VRF1l
tVxyEki/pz+6nGL4qjg3X5t5NiycJs+J0yF6gp8Q4Ni3oyLFPMMwOQKdkmPSJcz2
RI9Ab/1BFX9D/0VScEF74vEi29L3h2E6lyXWmtvGvQktkm8QcJET5PNhn694oebu
/J5VagWDPF+9BGBLH5gOFdHmyJAdcAIUtEBK6EBLaoHqEn5Wx2ZAmZnFP+ARfdgo
yj3Jh1I41XLmKSth4fTEw7sJBP38RtbYEykVW9MpW617PzX7/eE9CI2nrtAJq10p
DxTbkdkRYjjQU5F0IaYyiWWRp/7dnDDC2pWGD2midcoYy4EqodG9UbKJpu/FNIDw
pUomO+DzRQZ/7l2oCntd+RduddlRavbM3p5kGamYNKuNVrVDGBGVDtBIdOsnsyRh
FaYzCvj+kobLTk5aaF3GhwbnvTM+k0/4jlk9D/pzhwZpCHLEVWaG757OAa5u38+4
asV9rWoVD8xhfJiZaXmZAFQJjyuozxm6YlEujLKlb4T5AtExomT1hreBNIo5bWKE
NNDBLItLrYJIyoHotcWTZ2vacO5y2/Chq6FSsY3tpCXIBVtAVBBr8CeD0+u89r7g
c9/7Ub2yqaw1tvQiouaYDnRicR/DAhsCp7OCehjKmvLud7ChFq5fJm+YMt9Q1wDv
/4b8Ob2WqRevYXzjDxYgbFaepcuf91BIEjQocNgGLuMGlPJrinQUTgy+wpVQ2VW5
tcvUisnVywRSus0nQRoIeSJSB1RiEVEJ7HkBwvtyWxQsU+0svSuLBazscyjhNGg3
dun7IeP+50RcOYCHW6EQzY5/dYZpV8d7607nN4wH66vGcYIRGFkXnAUkktOS4eNq
v47rmBJPO8CGO98nSuAh6cKW0H3Fr05BROnUoa3GGIr9uZDsRu1aoaY8Vxw62rPP
0lHouwu7uzi58cgtc7wRJKiJBDrZuoaTyUjaOu7wwaSmtFVSMjlQTirBR29bqnYu
cBMc27CWOkSMIJ/n7qrHe881QZfRCW0BTh92bXkuRoyHOR5OkR+ylI81FSyv0crR
WfAjrjiry2yGih88ZpaPY2SxYEJdpmRaSnBhUMKw/CX78kB2/5c6XtfwwIc1H2ix
wl59WRpzbY2IvzClygIMDEI3PiDrsa34k4DFa0mE1UXdNTNqzbl32fg4lJ+hHDtL
hxu7kCXUO8WDIX0I+2mQA2T7l8wpAtut4E6tOo912dk7LsXDeQ2cjTvVHxK1EA5L
c83QbQPq9VOWdnNbew0xhmTDcPtARE0ok7ro/epZU10ZVewb620gEbzQ4nvYHZvJ
xeu3AywFDxS15IFdYDJmqi0tkOXX06fakicPJW0s21aUkL0ni/TJDxVy9yQnMRN/
EoDt7n2qvf05W8woS2jqsgOSjLYzXFEQ6DSZ4SrGe1vyTM9UeTdfJLo/wEk11rC+
xnMpL2jTEZ4HCv1iYQzDpT8+9l6GGH6ZFiA+OQohT4dm0g3E89VWSL9n+/QO0crG
30mSUZWiUEnHNf6NtoxE5tjCVITc7MmUduIvBMYR1w9YhHFaUExVjxlWHdYzuDkV
gRqZi0u0vH9ZWEwjf+sLC5BfyrvFG/rVHGoA7KzJsXm6qrvESfMDUgCnVUeYtg2m
umyyX+UGPg6kk4dd87Tg23UmN6jk3a5wbuopu6XI4sHou60Poo/tLPkcoTtU5nSs
IvHobS3dXNYIPbADCfrShrD4jJtY4nkLPH8Elr86EcZVp3M+UoagOmX73QfUHsSX
uyLzhOSIbWrduHsVn13PSBEalKFnMPzVbnLFwq7Ok1awLOD8nK0HjJEl2Vr2eIG3
VkP2SRirYw4ErnfnVGicqApmCzSWZqMIJqzNpGRLs1+TugbacdnmiT/6g8EUARef
C5n/OuD65rTlfiIFgkTEwxfmOqHfKSBhUWJ4GoNYyr0QaDE9XYpOQhDSFE4l8N6V
2JUA+jGPulrvJaaVpvU74jy5r+sARBi8ZRt/QQZc8aOt/caG+gLR6KnT5I+4K2pQ
s2X1T2P98Q0dBvkoo7lT0uKwxJVqoyO0lIrXqRIAiyOyTBAuAdRNAvLTnN/InDxQ
5DItw5UJJGyAMQwg8G+5e0Yvbgl9U005+TZq1PXHL/AVY0eu8NkFKJr8cc0/MR3v
8zHbKmCgJjrP4BnQ9c/HzZtaYS0CLMfaXOznzihbuISyrBWQdBfUPivc/8HA5trN
5RZSxFXKYnmR+2jHXScihNkar4YEG5+tuOeupiXrDP4F8hglgfuf+OFVlLWeV0Xz
Sq0jnpRIB1865+g5hragA6nLfpxtHLVNblmpehaLz3beWm5s/iN6M+l+KZDNi2bh
cclZKHTi09fMZERtBKFMJ9JaxgDKcQYYbJAjFO2o4GPBu6qo+SroV43msph5fUgo
IQJZC+BcLY2pcJ3yZCdTpWXSdiJqxHUH9sAgFiKFbROW0gqVMwusS4N6fjhEJI20
IJc2muaxzbsDzY5wq1m0lcu0z89ZFvuIGw0lrCdnPUblDPQ7X/hrjmp4WvQNZTre
c60TZuGKUKxKYNUpxWzrjStmMPWQuRCZwmETG4xOv2ChCactPs75r6CVvqyPTKj4
VFYq5NuOeSq8SUdGsf9siDSLjyiI99uSPIXlV+AemL2ts/XMkPHOuUPuXZ40dP9I
/lDy5F6tC4loNSYt7FLwVGKhdwiX0L0fWCHR+nPEz2T/5SCVvJqhUoDsnkUvNfWZ
DnRAeRcGeZlgOVr6tcsB+qi07ZcemagB0OjSaTOOL8pfMfoDDLnUtYA4SNmORgjC
myrNyIpjIuD+JaxceJYtRpG3GNX/bvvg82Pn8xlRFZkoDkxMmnDrHU851jmNQYIc
jTMTwD7GAHEUBXRdReBNFLqUS5xbCP/AQIWwGpbvAzEVTVufM5g9zz21e5qH4MwN
I0WdKkMuI4ETX/nj4u0lmzzAyA6+m2ZBpOHCNbIKuawzhsATzOcoavjkwJ8F4ERA
1gV8EOza8kMsry2JLbzSEQWYTVTwcdgGIoeLFz2rCGxkd8Z/OALRz3ShA3qCJOCq
T8403bdIQaBUG21lZyFOmMVQv5AbE2uJdS1cRYe6qyOIT9jtf4iFld3sMtU4gRGu
Z+/O9uAXy5fW5W5CtBMy1Xp4v6z9D3GL+F+6VS1MFiq7EIc0rozQHENdDsqf6/CO
4CJmq8ZoHUBx55g+KK7gwrpFyrl5yQKddaYs99VKX6bxbZIBLYcS9BP+n/CWAN9S
HJUEKB9YMm1/uXiZNHURReUDncXdIt0qDncqLAiqmYc8OW22xD5kycKaxF6oAsZF
0y84PgnJBdL0d2wP8VrnOOJD04kdytdBklZqXlQTryUGt6VD6PWHw/FyTet51Isn
is8cFIVxYBc+WE2oQ7fFPM/vmXZXtjk5JhG0eVRTIXU9ur1Z2k0regrBpftiqoKf
tBw4Hjb6gmaEZodWcrpjFJPXgmwCJDPh3EQZbDkRBYgAJsXqKYTZ3JzgAUGr8PvC
kv3IXq2A9XxK2JIpDdPJPAosQlR3VxUPeI9FXhQr8o9x+k6pJJlFdRqpeVsIBrBB
BSOG23h7TFOcnrM/QGSKdsuJi5mR8Ddp/QeHDcsgL+uYWpjwkT0LxHjvHoZnlnSk
8+Gnyw+xJofdPDwkt9Awiw6p/+amnAUwRUC6JUOvRVQBJy4GW5dhoGo7RmYB54Jx
Ze0H0gANGh7aVm17+DwVyfIRIM/5noMUpbPgEnbkbvR7C8F9r7HZ3ev77b35XCOh
rkacpv1jQ1YyIclbbDKnjyDVTAeYvv2kra+jDYoy+Sr9JVmi0dKKuLuYZVUcxKod
/3oRdcbEhckzsZD1jycbYA9+AhzNkJyDh15G78F7bjm8s8coB/83cRTUXKPu3teX
I19oDTu01X842XbfcgenLNFcPBqmCBfRGq7W1MSxGYplyyI1k1cUeYx6xQm1QjhE
pQL7VYODPa8F5KJ1MYSK5rXJJMx06cgAnRrVoc6XCTSbzyHRE5FRpUBbzHUAMSAE
fcGAWGKQ629Se57uJQ/rXe88EYWBBv49wzCtnBIOi563nM7rXkuolLag0eIaTpSl
j3BB0pqsmWRNxe5cpz5Uz7Y5IQKh/o1y4Ll/9YMa76Z7mJkauv11mmxPECfgR+39
QPesvKCb+BKGDOZYWLNS0p1Rq4gFqcyk9GEXzSnA71b1DxOKXq3qvmK7XhMoO3pq
IDclZvlggY1fdkADOkgqPpoqHJTQ/9UWbog/ehu3O4tKqQqLvhCEsWn5VA9I0zKz
2FEMc6fwYmNJYyPDic0mx98gCVomQNQdwr2j6mKqWN41Z3bJ60U271qkMvpBk0IQ
VNAveTaOeLv7pH3XL1sRNjOFx8IdQL+qP0xMDBtupk5nLhk9AVKcnQImxhG0TM0y
zxXiR7NaKZpju7RLltGIGrqihF4DQTB5bAi51r4ezBMTEDH7UFnuZauw7sY6ytC5
TVMEhSMuEWnirKcjXKzWOAPutxjCpNdHaUfqjY0XbUxrBRtlS4XcZ92zYQYhlpHi
+mVtID6LNqrpYNZxk6R37Qvsz56i4wXvNGeKSsEdaWnzGP1kgpSwReIXUORDGuzW
M1B2ekLiRsAHhyMVEMiMevl655lQEUBos3TTUHScoYNOydaDpP+ub1ULFFp7ihWq
JbwTbRKXrVyx4Jc6m2meWrxSxkIKuVFquu1aWJwdL0sc9A0MOyEkqgHcW9CT3Mri
zR2TTTH1F00Jwm63350t8Sc+3txeUSMZIdGPijEWRahrFr7AimLcQR7JO4ZHj2tl
bJsOwgepBXbSIjsub7BvIbQWQubJWsjOBzkkeKD2R3Rm7jH+8z5SpzxrV+sDsE/W
YzKbth8gT88jW/TeKnDIPtb0KFuLCs04lSf7wuH/xaCzh5or7hAYo5ZnjoyhZIME
cc4Kco1yNFcJTaZMLkJmm5K5+gDfKD8NVi561mpJBz81Yw/IzmXpf7jfMfkJT624
ZwrjuVn6OsCcM3sn/iDCgL0mHekE6X08TGdDzkkYJtxf7RZwODkwwtxdQ6BG6zhv
pyi3vIKJ6pNFfzQ6ROPoasJ4ZSh9Fc98ybG85K+B69sTOfuxsX7VXM4gZElIb3ID
Qd8b8aD+O6aPmeH8InLbjTUIploNNH6B2XcmMkSitnLs8duzoqUzzr0GtzElP8o6
xSX/HViM9A81UU1vOeKWK/h/13+Jp4GaREpcJgV8Q1nLZaqFOnM28YObryrBU3N3
PHEgSin+vCHAhS4sW0xO+cYruQ8Hg8YGdRXiCtUr5aWfBWxzASeHJqsf9raf2hP4
E+57WImzD+d3Z3c5UrG4cAYZM2ISkv1ehst0MD28N/WS3hBF7Wvn0Cf69EHRwv+h
5C9ThqCnUchcihW5YAWTHd2quUETkNz9cmtFEjVHdpQ2YtXqeh+/yyJcXeRRcp1M
D3x9rZhUu/VjazgrEcqh6lGLvHjyrq370X7LBtJd+68GFPHK8x/56E5r+wzGSmEt
FW6MF7WHGpOfNoDkHXarJL8NUs6bTP3XkW9lozKKJkzZUWp16ZoND4SBGVLSjJ/O
LMNQW/vUksFSss7kBzXjyZh3++8EYGKboN7wCQNWuhkWLeu/XTNTd1ohfcKMmns6
O0RmYdf5KICs9KpGhWil+RmfA9SXdHFN2CYYgJxx0nWDgduSAmar5qn539v+81NL
I+hY13wRVLJD+nFPsxE5YcOmWrrpckXLEkREVqmim23FLwfE7ccM+qlh15X2oacv
5CYfMxdmFd4PCI0INxaZN0NpYd9T9zkFY8jCJ2KZ/0RHcY3RtZ1E9keOW/aiQ6yB
ZBq1jK1KvPPGtW1oXviK5XBTpIHjfc8hOT3XBdekJDvhfWucqtUFjT8Hg9RK9oMM
YcELt6y81HOXEmztZRFBVDgTWdEMBizMinOKVUm3YmW2gTpSwN6buOehawzIkben
Un94ZGokYyv/hTpVrc7fz88INOgYeJRsdfkBrlljanoWhiJc2rt2oGLOBbnS2IXL
wx+M22tNAbGlVeFGG/J25PV2rGKEYa8AjEvCblKbuF89uG3/czvBE6C52BkwDSuq
QX2lD8Abk+80B4UvuWE4jNY+STb5xWR2aGrP5TKCAp07oQs6ZNS8f5FtMB2dx20P
PGIe3SjYVrq8Xfy4Scug/e/0xrQyROsFjE9xtlC0F2EUPHV5zYzPOroUAW7o0e4x
qDIT/dyJwpiCJ/rwW9m8bn6UQmfKp0q1vgudg55QgYMuZgBslvM3DlCAJoVrvGjO
cLnyBCTA0UiEN9AcXEQ41ARtGEzu9SEF8uD/mwLOt+VMEYHaXdgfLT6pjgOwuxPi
snsXt1dSV6wW4ciZYae+Sy9sJJXAtKPdaLUtmG7/v0qWVWrzSGr6d5W1hFOwzg7f
84nf3IkpvQW3pk7o2gd8mMN88oys2ciN/HOFEn7SnamHN9IIDbs0/6qFvojJ+LGE
kRQ0HpszZWKA3zGJGRexG1yby2ozRyzHuJH5aflCj0qyH+MCIUq564JSGP5wToN6
fAkvqFIgIKe+ZT15ck5XywKT7oH/JgkLRJ/fsTm9NVoeN5Q+3zSDyqrYozRJWjYA
01WmZQ8OjwNtymWtihZamgr+6NKhSFFj/JHNcY2/bJY0RnY70rNyWSMTAZY+Rz+p
JhbQIJ3oBT/t/nZcS6m/YIrZI6T8pZ+/0Y/4HmiPrLySLY+rCN0/KWQqLqLZZc9h
nEF5P3KUjA1W91JaRV/i3p2u1n97ezQ7Wwe9626mV2Hn6UJsc0YPAeaLEnpohBPw
KJ6mrE3ACCWwZQhjjYTd2pT9LYbVvSdkH1vSC2yn8BTLvzgMxcquDV234tRw0phd
ZOrzWU2Z3ER4QYa/aRPNIGl9frUsIi7XgAPAIlQ68txnqeXhFj5Vt5gqs4qXBTkG
WsJXpUlwlbNkXTnQmIOgWUwk/vmlRO2nkTMs1C4PkiDyJgnqbRgGXkuJeiMy23HM
0jNn3tAmSecUt3oVZch/Z7x5UOggSYE2Rb2PoG1YtuZ0F2Qfny4uq3LaWy7yidh8
ctydiBJ7mSjj8/pLYUaqGzVmI7MlxP3qUryLNfBUcofnOqs0mPE8o+U7rcNev2AL
Qss2iod/82A6QAwBgjMcu0D/ly1Jid0Pv35uRuGj1BMtzJAQNgANWOOM98xJ2pGX
ZOWNUffWz//tNT1eNigEVImPWN1sWh0X8HeXSAtqD0s8hOiFWzugHfQiOfBi/52L
cHvUpC629+74NWELk1SCkQ2vk1TxzYEaSzjRObOCZ52fZiibCVDSVCtyM3HdGiOA
gNklIPoYEIlxOnPoYpRvW7Y6YJyTPAJKyg+gwcRob8OADIhBBARDFXjJAp69c7Zr
3Ix0QteNI28UY/joHVHedWBDPez90LBdl5m83FNa15j3FrpGOayOFCX5CR990VBA
whhuiv8OIfr5TkrZYy66zRXhhj/C0O6JOI419lCsEnofbICf6oFFjgZmOj9R6+z6
byh9AxfC3cd3RiSa2QOIe4IyznD2HC6b3M4BERugJd1zBhpDn4BBAxEqxOFlN5LS
zAvGN5s2Kshee6rUGHp+kW5qgqrAuw6j5o0pZTpqB7h54rz1tyj1N8AjJOeK/cWV
c0/XwgYU3vnzL3G9Dip2H/BBDlV2h3jfX3NF7V2IRigh12z46KPMwMhX/DN3SzIu
gW6PJWWQsCPT9zbLFJAd2d5KWoI03akXQ+5oK5J+y4fS7St+fW9hNDyU4uYT7TiY
t6T96ygDrIEAfCIzCeSpn9m7d2nJFEsrHjvblsVddeeobDz5Oft3YtM9cvOfClhJ
1CESyQ6kYq0jwj5I9LHkw4Cp3xVD3DiFKSZreggCltPWZQxx4KQBiSWs28rs4yxU
6OfXviNO89cH3iyp6c6LjHYr7mJ33Vh77RpiJejVrM8IVFa3Vrnvw174DqtmFPkn
sk8QH0+dszuC8p/ufmDKmyvl5MDBTZXn0RpDpFjlOt5kiIB4JeXV3uRo1buEApEV
4Ft5pa9fxlmGMuPtNPNNkV1j/tFOZyXevyaGFkRQtkTT/6dDJHnT9QQ6rRlpuIeR
Kww1DzTjOjApilVvhHIJcjVLNeWefM5VWP/1z3f1YhPp659w92YGljlZL44OpP/B
FCpaWMianE/HBnPmRRDyZKWmRvx1bkHFIlhgP7uzxME+TCUcV73NilGbXyQQXpSA
4aZwPZZDXdt3Xrub9ugbS+HaiEEEgPbpMMaN3HRquStSVgbeofM8xic/zBdyIous
hNKaZd1vFZn9h90KN/bWmXB9zvLMJ9gS94aELJtyUcRr0bMnC0fVr8yG2k0HQb6s
CBw6P3ZmjQMk1r9POfwdZmhSQKnioAdoxWuQ27meYkKsqkfMXiHW30dLcM+WyuEw
xJLtlUjtpTTCQRM4SeKa9Wzf+XSwwYrPfCbmo//VLgeMnenvzdBLvYfeWa3+yxHH
OmHPR/6FvvfbfjTxQgfqK0rPIW6x+whnS/J1ATMBNqPLR9x0i+Ys+KoW4gBN6Y96
eC2Hnr6tq0D+ctpdH5+gMPk8XHu15344Vn6NBaIsURemN7dYNNHaEDVP2jl1XsRp
n8FBjp+4bLvxUi0YiXPOt9KLAZD/14LJ8p2UW2N6dOzK6qQLuMECP9L75IKcSXPt
1UYJ9uxIP6aqnEytj0Gj3IYrIlXj2avy2w3z9IhWrKaS1keoWO4Yt24b9LmXAkrB
sTPSdfzZim3DbR3+YXgty7xvFOBMuit1tUgnRxjg4YEUPMpF440SYkCKhx/NKVA/
FJu6940d/fQQJACW1nrBwrDDB1M2Jdvi/wdUO/BIM0qaMKbtUxlNFj4XYRQwgwhQ
WwR1jwn28lw/ehTnGLcEBPwWA5XjyV8ciCS1l5INvR1wU1g4B9UrQ1iDL/M7YRDA
wQKhXTPDXMzA5QIBrxNZXg8pVzneY+f/KJlePyNsHu8QsdDHrxlNbl+GPKvbLNNx
cPv4fYhekDAxXoG3fmkK4U+/vmQmorRCz8tTdLk7SfdijhTlPPUfw5pz+Hf60O00
2RXrlukxBgI1ABwbNiZnKM7aHxr5AQwLQY4CXdQtkF5GA1PK8WuhK6F9SLhjn4Dx
5jnQIeE1WBx6a1/DqPKW4yLjDy4r2rhShe9rw/FcNYO/chdCZZJ3Y1kUA4oyHhBn
8CLPhYXs72ZMkjMSGjnJawta+U8qEIEf5w8DG2vGRaQbLWFG+H4gJhXPMPwpTKju
lvm5AcAUqLv96IfBZe46xM6U7JkMI2dbJ22Z7QL55H8VSaDHCCu/sFLYIDly2EQt
X9pfNooXGmq+WQtHQIX/wVOXGw1MGXFdZhnHmYyk/+IQ1jZZyssAyee1Jb7D8aX8
jCSrCR/OOTtMZWLQzyU8JTets2DQFzKn9i61M4EfuRuz5210JRo/YUqDDHpkdgzV
9XwqrF9IyRAcqUQBU0aIFMmiSxC6ob36XzAH6YnqKEvbXvp0kNounXbdkb6M+eVZ
DhzFucvw78OO7GrZ4NskmCZAEQjaD0Yzqaez1cGbabmes24SmWR+7f3pnnIpYu/5
NZZu+Npypjgcq25LFWg9sPVbJ4QRC5871+H9TbVNDlffyRt/fnU7/typykeusKrm
/FWR495HhEQKQvtdmdydN1m41D1IfHX2G01xLI2pRjW8YqKntz7Xe6CUaIk4bVM9
nAd6DpuGvM+xUvtrblC1jqChfALkxdbZReSSNCJVRT6du10f5LYUkxnS9h56HzlE
ahAIR3rhROHRttyVQqjlhoDrqZP4d0jSaJiIgqVd9oSFMH9QnEyT7rSzm/nzftLm
27jVu6oczpdXHmiLLr6LT0TA6zHVXs/dUat4Ra/icI/wpCJyBDLUA8Nx7OAVqsp4
whvV652ZxEm6cZFjJxORAtTvYcGSeSWS2+LJLI++hgTyAkU57nxZuInntLn+jTC0
NaSaqlan62M5FUj2W2jexOMqBDu6SiTWsSpjiFq04xQt/80UDT70CCug91uQBFh9
YPfInfb0JaIjqY2qZ6K31OGhFchhjuvAwNImcSHu62KujxIeEnVimoJH3EXjMEdn
eJHCvH/DtmZKpTgrBGQMrL0DcgYP0k7HDk4HSz83lp18MeEkluMRvV/y55uJ/cie
+KlajU4YabEMer+qdpizFK86IdRmbO/8Zhw3Awsa1ry9PuMW31hiaC8DLQxYGGxz
InUbeyGHGSJ8dYS0NGPETsLpDJ4WajXURsxxwyeL2v44k50I1lAcmrNg0TT/b/W5
Fq3eUTpB8OkSSB8q5aQhlH4h2Y12lnBevZmNZTsSv9BJSwPiKgQcpl+3WkkM237W
myeofPzxC/F8w4e+l/zjaSeWwAd8ypFQMIp57l9Y2UgQuG7lEPukG1LtrHL28RvO
HVTELyEd6WN4Kdc9tQaWNypsc7JII1D90AwSNgDle7G0PKqTWrah1kwzkeNeXEp1
e7bGTGhAIPDITzCk529ak/diEX8quuZW3Lni+ecITnTwPg0XRq2WG76LJazg+ffe
Kks5hlxE7J3FmUFH6uAL4lKE2+TsDc0UyuTYDVAXz9qCtegXZXSYg0JG0B7IriFu
3vNGvWfONpnoz8UgAupime7N3hqv4rcb/N2a2tKjH1eri1YzTej4K0anGkSICqgJ
WaG9BEM8KBOEFgbYOOrwWQ92zivvbDFXCKE4POvBwKvnG9fB1quLztOVNkLCOnww
x4gEWCnqbyryL0WUuLA6u92w9XhMBfbEoYWP8CS9Xmpf9e4UjPnohvlKmwLNUQwK
o+EOM2C0tE8nI+HTcSaEhTqHu84McthGWsidb+wh9OaN9DY1qyttwVKc7A1UHSYE
3/U/HwV+ew7jXict8WaAgDtp2P2cm9+HZCtHx34DI+EJen9x706XqsbRf0NiUbPk
3+iyd9RJY819EzbyTjfjUUlt7IbO+nPOAyBery+b9hPM3qAzOhdvnhymXoJ/U8Gh
r3ZKKv7a+0SomUzDD9f1Zw3w7x221CORlmV/DLh4T/7WkreJgFgqPst4dqWg72vA
mlOpHO00d2ArS3jDNrFVhfYp8GGK/XFAmeQeEhA9dk3cu9H3x5LYceURinU39OTO
nfZ7z6LITzWRhUxPqJgD4Wn7GNN450W4ToQb+jrTHOZmvKQ+9kKpH20xS40xJXoQ
eqNzZXRHdoXtOiZccl9h0K1V1D3H4vk3LB37b1FLsBAEhT7uyvlgdSm0gZp+Dpiw
b317EmWWpyb0ZJYEKQaOmy3kOj5biKizGwq+h6EQnv1qugNBgeoQH+OYG+YsThEt
AzX21PBtYvfe/lJ4t4nJ/Wdicmt+1zWZWwzX5QI97WL6BzFkqbrQIAPLxXb1XQf8
8ob84jKq4JoKmcf6GWq8qLxuz1VOKb+KSCPakDIgBOr18cdJg4ICNbtE2l2s1sc2
nyJLw+cFG6OP6TFfNMMF/ateDxo1aEI14NiT0p7bBvy3uaG/X8mykgFBarlwzF/s
+JVuOaePx96tB7yqvaxeBXfXsTvkUFC12FG9Wtb5biVsMpCWLElBKbgEU5iZF74P
JLZpB5nbz3/TtlsNZalgAPxecvZju2W9sTvLj9VQWaXr0HNYYw61fcgUBHXEjji/
iUtT3nJROHIToK9nU0fbFYjUYD5RQVFgugc8TQYP1m5rALKVeBgScGn4U+YSX5PS
q2TyaISngsmLpUopH5K0R8dVl+Xh7viaIHuZMiel3/Wvj9RnPLx+m5C5pkqnaA2M
JQPeHbqVQGJrqnB6Sg8m/TTOTzEJ+BBkVoAimsG4F1uONF4hvf3VuAWStX8FMvvQ
owwyJh/Xb1Rmxf8D7azzGfb11t1tAZVA8qEOKlOWBBf1hIhDUY+Z/aS8TEPFYFNb
o90cc7xa5pQt2+Fzz2wRVlSRD8PMFw600Z9/f9eYVaFdYgwxDVI1DHw6+6GNNe3a
gF8+qPaThCMHCfYWI10BzDb+up8+8SbZ+bQT5whpLBJeKBjbWFYmtTDqsX9drFQb
P1UaYtpHZmZgOfBVGxg6kCA1sgPYRCRrf1SOOAntMuYgz/JzZHnjADFdNcdaK7nv
i7mavmbNj9UQtRbViHAAbZZHn/KakmZ4jsrg4MctuRQVeBvR2Zt8w/BlFjD5M0Uh
mQM8a1gWJsk929P+NWv7pH8useRD9ZLjtBLULOJVbBX0jLm6hkhYEA4dfovFydaY
6Zi+5UD9Dts38U4yIvchN69e8dMeAYkZLikDDD4h1beDcB/WaAD619XHPLtrtAGI
4/wJNQtwkmhpjfGufZjMm2n+Q0G2KTgRFXRuZiTVn5UBBZHYpBF+yS/Vqi1y29Nb
l0+e95ORw6fZ+M6WYnnT2V3J5UYqV5xwFenxpJl16lQoEp0KO0OZS8Q3PJrzgm5P
rDNAJrycjb4O9DirEvYcfsjv//sllNx4zxlhpu6X1tdnyogyUxaJ2ycpcgRHlkeF
o7v0539HKD1VLzg4sEGEDyfMjsTnX+2/qPR6EGh1RJ4M9gg4XWcwRTA0Ha97vPcj
3uTJSpPhd38oEPVmGHqEot++xbZpvQZRpWZA4Eduv4xPCX6x9+mbALWQK1BkKp/t
PrHZ10o5kbr74UNsWfYqXmWZP2EERd/vwmKrahdKRfiwHVJRonJvWWSFf03+plbn
Dug2JiBvvBd/FFWUGexAmFe40FUfln+NQL98M2Mi2lx+bKkZ8IN0jm3OhOnX4xgi
9I4w1mTibZaEspvcsCP22M3xxa+DSAOjf5ykgyDvxw8MIinu80xh2wKUCqCS6ldn
PedDDB9aahFFABsCkcNhcjxHs59KdwSYf08S930J9+7Qbe5ljXXjiIkzU/xck/3v
r81q8hbt88jQdVp2pZKhOpyXLm/DgYVCWtv3H2VPjSofqcXq1ywECREKR0IJKGFB
Er0N+O4BzwO05kMFEserqqRh+ML1C2GP2N9zIc14zgTxRLZ5Njc+v70aJ/x4I/71
eLNkAKmaxlpPj6KeRF6wrZGkR+DAM91fR991+fv5cUdaA308vyUZVZg5/01SMKfS
hupDxCSKzYMiyAfSa6EzpZXK7Fo/s9nNj+nu7DJCr1kustbdOYuzR2cCGU+kaTAt
bUu6hx/wKUkff/I5Taenx82c9v5mlTYj8g5tw2GWg/O9bN57QrKJK/9eE7DXNvrB
xeKE09icqwJ0EJxdRVNKMibNYobUEpLfG7FPSiKlWzFxbsf+uxu05Wy9FwcBLgw8
nQfwX+aFBc0YaIg5lQGXxbQvh9dE9WGYEkF2xg/4UxCZ7w/sNPkf8wfxQo9VH7+D
7KCppCowBJCh2V9mRCsfRSHn+oEofwxAGrFasg7cLbbLmHkRWTVF1nVqHjTU4g3z
lD+/wWhC1tE3hr8zLlsSlmuxyxe1hp2e4csSgpWBtf2k5yUPOeyh8Yenu+hiq1p/
egBnq/mQLmma/jCtkkmry+lYHEeImfj6i3qrvaT1WfTQNBkBkjQr5Z0S6cxtCXVr
7P4Xo6T7Uf0wSEEtUgB9n2KK0yCohPTxFbQGamPeNIMToLZXWX6o8sV6gzNbMXmB
Ca/k9P4PKJH12aFs2za4jB+1bxPbPKnMn/BFExwMYa6inFsA2pBIlnFB7rwyWrkW
Do81zZL/WbICSGAvW0Te9had0w2PWLF8bc77xsZHY6Sv2tAN7iaGo7oQxGdU1oV3
LTTsotPutBsxoh1Rxr+VMoZai98+aWb4EXFLB+7dfblbSRX0j71eVvstfC/ky6Ip
9BkmN7cj9COrbefsGudssuohZm2ContDtsijlLCnvCvdOKFaRIrz+pxQZRvGR7EL
4LWkH8uqBCyr7vAPbhunD7OhDMTfX9Pcr/c8ayLPzZuIwWTk//X4KwxMqDFpEiDs
jzJn2LITT2GKmCNW6uC2q1nr6XV6dGYwWPLJxVNQVu9g4+E+aNdggxwutkNFUeRQ
q4VTUGYlpCCoy6k++vDSC+QiW074EX/8uozRbiz1xYe8Aeg2/PO68VqIeQ3b+Way
FD37ZlZ5I/XdeQJpsRH8nBU3Y9vy+DDfgF4aYHTsasHGkSNQPL+xowMIcSn+Y3Ip
GkuZIC3Ngx2tNeJBd3jJEBPOLlR4ja1Uoz9sDTtWTrMRzIaHyvyqb0dNDI9AaJ9e
KACiDYQne+Iyjnp0thdS3IDpMTH168R1PHzIBuWoFLvtylmXUSmcyMrmLUqPQ9GY
usLLBNxAxHulqoLX7oO7SphNauQAOb2K5kh4mIkwfW4fp1GA4lx99qntMsZ6U4BA
G4UvHCzmeIBZGwncXWXFP/BQ/VM0fl/U8VYDYgWu7InLGhVwQ7u7+S72EqpPANOc
GGc5xPAtJ0xI5hLmAjCCn4QQUmm48qUdb0LFm//99Fc3dy2FguPyx3zu7ko2HrHi
WeTdRqBff/5u84w0vgHIULgD0Sv2UGjdTxXY0tDbLSGmMQnH0m6pvrDJue+C9ORY
+V5r0IVHJZ30LEfCJMt6EPAC6mFO1k+R/bNQ0rhI3Dmhe0+GD60AHjNm2azn1p6j
0E9l3ThPAYfYLiqh2BX8f3cGVnk1l87mJZvoLfvlhE4TPsLJeqgwWWM6rZHNMwJK
UJ2BrP/unf/y7orBtZUoZ4cYiF+fx+kfLBXDBM89JAm+tbqL5fr76xjFnjm3OzXc
DQxgvaXQgHnYWRMP23ig4zC04Npv/kAbGadYa2YTySxmhvR77fDM4CYuxEqIWQFJ
d/ZFAiSWhWfKnQtNQKdtckd9MozrWFTmhmEFVfbXQn+tiPuMZH9eB9dOzEupBkp0
RkfSvqYtzSCDQImfI7TBTVYliMWnEKOir3zKGz8cMfSUpYMDMqCm+K7YBUWikzO8
KAmJA4O43VwwOl542K0pktj7NrAFC4hspYQIzF29VUFTqouFXftXos0z8yjWDDCG
mJajg/SDHzS28G1CUqZiRBSZnt5ruXiA79QteXjOFdsmBiQJm4OynIr/Tf/0a/1r
HKan1hsgu+0ibHsjauNXtbNk9qkWs8fyadKnWFQmz53kSk8wTqDiwmgSmpij2SSX
68RWtZMdq91gPA7eL3c7l/r1H4ELgS4HvGEYvUbfRqCwzYldGDQxQpHDDAlD4tyJ
jrfWF50VSmWONxTqMhrP384JptkD75a4XQRo3PczdokpiL3Lw0zSDadfvBpgDclF
OCEHFl7eEt6MpDCmQYAEb7WLoNj+9GGg3mbD7oVRHOzX2cobb5t42wtGoiVAHpc9
HlCTCFaESsQSjGjBVi6SSfX87s1eTUieV8R/2yKEwQ65uRZ+XjIwx0SEPTcAnfrr
FuA/YMCJ0ay42d32p55y8wzF/+UNobuImBx0RBDJKzj/HAiaEak8XvFKqiowK4hs
5DUp06tsyHXIe/kPn9up0L12TUU98LcQiyl6vpLYNx8Z+QO+JwoddQjtR4r+YuFt
H7RM04hmaqxhNW1sm+ysIqSltAEO3emwil1DDsFaS3dGK9iRr0cU8LC/MLYMDOEb
7XPft3xRiQUYeBTkBaUHJjtmHO0IPBN9enPoz9q3O+MW0FobsSjV/pRlaq5vn9PM
7SZAhILgvljPi3oP18EuC67wvkIUfJtL66+Ia7Aj++9uXoz3+Jejd7gPrENmvjx5
4MSf657gQmQvc8kfJgGW0wtBcBmtaZt4BVkxQDCnIA4e75CspG/HVWl5RBybn8Mb
XgXGQm1jQGCGzFwGFFJeAwoD3L+Hc/gEwDb9E/aOpe57ccqKl5IaDqI26kpp/IYS
ipnCA7VtyjTED5TgW6jFYsjCNczoHOA19CsH2z0GQBBVDjksMiPWpilKnXtOPAQb
xmz0puy4DSeNl/1Z5a4X3+DncY/DEAIaeDXd4nArIWSaABgdovee+ENGkI/cg3Ci
Rja6xheg2U1QrnWRwgthgJ9XeZPKpRRyOTDaEwOb+0T2UbWx0Sjhc0huvTzj8f+U
1qosuCQTYLbyz47+nlcaXaDXixefhyRThw6dhvwFJiDhCVvawt9PQdU/jxJia0aN
In+gJ52/tsSX5MvMfiyES8QITiFo4nB0rzqe9ey3Bv+YTVs41OtISrll4yOmbRoX
7ChIiRb6NUfCaz68gKOjnR58HVvW3LJimqJyMXYXOW3CKiRDMptFh5Sr4HNG03bL
87AICuBEsWnaDcLXRBQ5b7hvYwDb6/wZbcrX+POmVnI9AVvV8/UymcbxnisFaO8f
kfu+fRXw2UYSgpoK8omqpNvio6NwniAkL+oKm9B931Tg/ZUpnBgsS5JDdtrwwq8x
sSYZELhbQFzwht5wdgEW5qNNO8UOH14JaTP6R6H4LeJLFQwa40ttj9F+GXZky9mJ
vy6hwX+KNS4zC8uZUpfFE5IRT4KkU7gBTGFYXMoKKC8vIwFdWvfQw2MbGrfpW9mT
7IJ7aDDAYa6pdBu5uaF5dx2oIA7ydStraRc/xP4tJsPhXyK5kpRdf5lWnttQHtpz
kHwEufGvIvFGmF0ZPrH2T3APqsuFEMJhfwNxcyPulZfoxDK/cnWYyVqDskWM3EHH
MwEVzMw3ifH9q5zsf4yMRKSlId9S4UtwJ8VMBy/IeYbH8G9r95OJW3RgdB1UOLhv
M0BEGfwFc5n6KcqvunfnRuznrP/rBeY/IRy+glpCyDQCNIs+pEqtjS8E9FrUJ4nk
5mDuIJnNQF740Vh2SDF1CWX2q7h6473E/Fg9cfpXe6r2bhAYKHn0XBsD7o9tDrfj
msfqcU6jAEwfI597J03ezEgsk6HIad1RzCN02TxKN93hIOFLnl4K4NO67bgYjGXY
qamEF1qtlM8j1JMWopEu8YpInnZnMRnyBBrC4Pa9URUqc2cVQXn2gsUkwZe1BpPk
SqggZFUc2IOWDmQSQaQbufQkhgBcnGgCAUO33tjb7LT/b0wYw/qNummtHoB2E6nK
ICg+9fQk8wQ5pVrXBrSd59oGQD9oVuYXD9ViYWZcPXnm1WJc5zyivPqLUd+waGKv
qduj2+dHEbq/tQLPkXQeZrKGbYLoR0Gu8ppY28ZRCF15wLrqsixVE+2f7fI5Je5/
vRiWFVgfa2xyzYEynYUM6Cgfbl00gWeQRO8ouKwaVOCqBpPQeyqO64vfDHokRVVE
CiTqHMYcPlSDwWImylYqHe6NwySS5v/qR7X/QoYVi7GUnZbatbQFpm7DaReQkmTe
jxHj4wADqH0tQDunR5SWerAU/xkP5fwIFH4u811iDwzdIX4toL8T7R36Grx54mrJ
nl6DXD0lNi8D6kzYoBaWyiN4N8N2evFXS0kUZzwhaJktgD6POwQLNFK2BtJInBeh
lZYVmntR34NQxKNgIaOcr/v2ecKlu4cns53BHmqFPgH9SNkCwCTlhxD/Xz3hvHtF
o5nBauM/lpSzIavn5YyH1/vDJMuFaHDhbkLbFilZjvS7bwzEovP8zMTge4Z1WiJT
I4QksNBoZH9sUG0jj6lj+rrp4LgYVV4/KbpMmVbbhgzNVEX/HfNnXTRPMebdSzRH
JfMXCpKvpojE1AYXLpO0n9Hn0qdlkMjgZRMohX2tNcP5oHRaDL08MgKW4vLmYMBL
wn/GJjFYqhYuG1nVeHZPK9TRfU0g4wKJVDKJoI15G9X61nRLtDy9+I9hXug8v+bO
c03GgxAEZNrMPVtQlCsEBeKpbJ3NhoXQN4Lm4Rqo0MNF9LW83bHFFgMsyyoRyj+v
966Xk4NW0WIep1J7AHtTSlVZK93oXKIcJBlNfjavLkP8KXXUHuXofo3jp37U643G
3xFWD97y0EFFj48vEKbaARg2h6dNHevJF4Hs03Tedbz1KE2KwAywWjJtTRFFjdo5
4UT1qyK2tQep1nbK5SbSAS6jxsDEZWTftIFOWtYPX9PdVths6RVccVtJxD5+zG/c
wJDETeQ89PToFXtamnAIYtILyK0QJzvtW7UHk835zN07WbmPR7HNPj1tUVeFeIXy
VyRIQWn3Jx1vEN81bKOk/lv4/Ar1tBKPrA07xU9m86BrpiC6Gn/H2Az8nGZNwdfM
Udw+Exvldl14J+AnAL0J32pairJdQomf84ZfgVfK8LidAhRwxDw0ylk1c+hKme+R
f8xPcu7KNkU6WoijHYCe85mYPJ+lAvPQ9MGxQ+0t/7DajYPgaFUG0YTYYjC1JpEG
EPM29KQ4fLHTnEEwpKdafC8KV7aw48ZER8FZPJfemaUQLOxsJojdhBKAmKUhN0gu
L/5OK2MxwaWZP92brebavLcQQ3riUMgA26bqW6oiYANP8xzsELDkfPbbQdrUMAQN
txai3XJVB6f3/k10a8Jjhj9+3dHOZJXKu7MjvSgTxLD/NBeaFRgjWNfHouyvF2yJ
b8JNYDROsWkTmsaKo+zKt2Tff4JttxghXyLuMIFE4Txp9Tch6NS5WifsZ3LnwSdR
YV9L+lHCQpBFvsJrHu9iJsy2jR55CQJiGI8IpVzu+1qCwnOcXRzjNB5kxYg9afv+
tmKJddI4PuwMR2RYOnACDgTic9niFhExJxiizAhRMaZ8NxXZUBWFysu7772/4plK
NhR038p0yUa70KB/RRUn9uuqw9+tPEI65huVE4gVsJzudRAW2wjtgu+XkzSvweoC
/2h5Y9aLWWm7NhKoCBGXOiRjRN/I3LsMeZ54+LeVPmPtYwGfxzRjW0E6uRfkAFwf
WH/bINc01ZX+/45355KNwMZFPXBm+3qokOHojKIOKC/MRxYIa7Ax+6ah+vE+NVie
RfmHu/QtR3AoyfXQRqHv7W0RkQLJX1aRPSpYoEBi6Jzg3VUIFtvvnZNzW6w2JxNt
VKlGv3hjd+VFw37s6+fsd4pwi+5fuhI6L46nXCHWI6UDtU0U1U9GLTTGkjETZ2Np
4clzQ6Kt+bQL0g9u/HiP5VKZWvIoqNTqRmWSh0pVcaQR6qp8vzx5lqGgnGa+jP8F
qZQqMq6mdF6n0sdkNx0OkFIEn6VSLvo/lWQR+gLnLKXstVDG8yLyuEKjaFSNCQRN
BFmAscdHBzVVZk2+FHPEgJ5yuPXnFwmbIVU00LCS1xdchN77ymbl89KmWqQ78FIC
iMpyTdrP2GJMgVRg/HI0RwcE3BLLAjx6ElHemEOBsIyYIcpYJPkr3qReOnmi96Gp
7sjBwRwZBjMgv1WbrmzbOjrDxN1nL6nus4tXnw1ejt5BoyDWbmHwINYrEuNI9Vya
pQi0KLxTKSoz2+8Uw/f10ItFlPMLb+lxUYz369lDvomHTsFDv1JKnUgOG5SA48Ir
uv7KDLLvVAvPXZKUNrFWACq3ejT3k/VeNVE6DPsJR8MwW5OnUNpWvIW7nKQZXFf8
1WXjoe9CsQ/9A03qr5mF4jLznJS8duTjIpnk2pwMApWEQgFaghl+GrknZ84mUjA1
Rd2i5cZ6xkZvFcDsb658ip3gE1oD8lgn2mM8RTv7xqVA5BKTe088M0UvEjTb5sq7
gBbhBEhpwc+dtEp9RScXuuc4vyzYAfAG27gJTFVhn+vuyElOp78ldktr1F21frV6
YXAkzc7MbgTG2OqDB1jAfvCb5zmcIKeenLP3O1Lz31ck0zV+4e7shbIRDgR7h4As
vWQ/eP8qYJ8q57235dHewZWu80514+mfQqM4iek0r0Di3PCptYmgRZ1rYY8ezRpj
4eH6yzUwvViCi66chtlAlTCx5it1vjsmxx99S9rPCajUKTQwUB+emp2xk/tvLI2y
c/s5vwr3gA8l6RiBTuaL8v0cBtC+ivJusV1kolfoiKX65Xh5aSguBXQI8goehGFn
O5mDjyVUrxPpV0G8Y+60GZH9rqfJunCupAYLakkpJMtvgYMjTLQn0LZmZDyq3MT3
g4Ky0MSIlend2d5nqBeTK39w/E/i4dc39TXOTEFdRsfNNcHt44YOnP/5miBkjSxK
ADzSxIpPybRkQS8uRuLtc8REwgCkFez2wwKHaMH/S6msycJD6dlLfcc5oCzw13+q
oiYzFYL8UDjbvBAeALb2AiLLNPy+5gSGj021q4fn4n+BkYy0xvTKitnRHYw7DeVR
ic6JcRhxe+4HdqDWR0lu0NUFacl5jOEAdZA8kf14YGDzHImmF/uNwuXy19Fq7o6+
aL7ISakRFXMAt1/OWv5UcxPS8fkE+mXTQZ+jQs7ANzFz04zZ5/g4c76dluGl8UoS
gGqDeS+EnLF2sZm6SP9XdIRd0YVIQehuLCHVBYiEW0CGxZa+JVRUS71s+lV8I8lo
/A0vCrgPD27IS4a+Ix1G4VNndTFf+y1ETh7OTJb4GA7EKmT9j64XSjsXBWwfvLri
ocQwor6KlTSAWY1XrDPMY1hjVpm2wsgDhcIIWb5OotgaT1x2WNB0nucFldKw7RPo
MH6bvEPLjEXN6bf1g/hp5+53JE2nGr6Gt9OesVGAHRkVu8ThmlvrFB06GqYKoWX9
GH22j7Y7uYPwdSjhpyO2w1+RarmH4nNqYJtPRbcQdwr7vJGj+DgaSbnw0i2l+Scc
jbkvVfrJyi5KqBlD6OBOo5qpb2kTbrWsJ2cfVo7tzFsQ1X2++pBjd2zCNS7FhIiq
6+39xiaIxs4F0WIrWS6YUnooxXyX58/ndRwaKjz1fCgYogopyBqSt6BNVXp3n9pA
jjl/jLpRXv1KxG5InT5Zeagk5FpiNvYFRH48ZbCzEol6vRXaOvQY7ZrK41ujGlm1
37LNol7lRKuJCvd2rzznwlkaLgkviHZVvgSqxXdJdF5Lw1O4snpDJThyr54fR0qe
q9zluq+cNKLyxZRMTuZ09806xLxkzcO0PQEMWdcU2Fny/c0zBaDEAGtYl15mdNj6
wmzMQeGQRdnVBbg01bEIyNiiYTPtU3kU7Gu8/0yyevcbmBkalH7JBqY9HyjzHxTK
kLx2s/Xac1Z4uSrj1nFPIyBZmCGUBxqSe5JkSCW17xLjDt3tI8jygyEPukvrmruT
hzBq0fyhbfjx7yh7zPH4zvVqpgOIWNKXHCDymGh11gw2AJ9uBvsc34ZkdqD0JpIi
JkeNZEly5BTIMsR+FQJCX5FhGRms4jrZV3p2yCgRJ4fx0Lw7n1qmVxsxqhwF9P/x
vlRaaEdj/mvS/Xnx1FWU8i/J2cGPJ9AwQojgT/HcMGpK/W/O56gJTb3tpLOajFYH
lUwgt8GxhL3SP7bA9/rx+Lr17oVOfEoheuBgMZW8rjAD8R6BImBOb8NC9MnpjXIS
IaxsVUar93cv3K7Nm5PE88t89QA5HvyKFdbJz0P+XOfJLu+zp5/rBVc06m4YRHQu
iBALgp0n1sOp+II8HlLpk/+f9FbWokwPi7IVoBvgpmsn3yFz/kcngah3nyEuKI/d
Ci+1RQxdJjqP5stPzoilNP3sXmm4MYDONcqa7SIvewFIKqiZezBIF11ZB2kZaHZ7
f1XWMoJdQEJBUqAHvlYr5R2F5bt9UL1rClDKmBOVtBhO44sBrG92EMLGYraXwZNm
2pWJ5Rv9QfH4/WUEl1+wYY9osDBSJJMOM4a8BMnG1RlhmD6SMzfWuOXziVnYUl0H
yanmIip6H/e9qef39oct7QeTOSj8rnkkJ5lYpXqxBxkpjC2YsYtZrU2d1SUf3R65
dryFfcBX3efzhyx9Zvle8aBf3dYEXPVHah0hl9yHAaMNzR0eMjbd9zaIxzPfNP/9
6/r6rnXt9O5bgs4xzz9iZfJFcv9bZbTFjAxihoixnBs01L3N3JXQOv97NTuYzn9i
Tvi2sGMCXCkEM140E2UvHvtI6zrnrpsV34anQqqf4l2prWjd61uCgPQH0BwQ3R4e
GLKhyrR5IjRk07zGBOMOw7mjF4c8FG5q0xaQOv9w6PoPz9Ds+R2CEZtHiwbnz2IH
t6aDwLu1xF1jzyet/CjDf/cT9T0kdgncudI57iIATjD6P0fi3jT/lJ+y0oKJB7sn
CZBRS4cSShH9Ih5zY0x4Qhdzb++qAh6gZnoMWj844T/q0TfOdi2K5+9mDYMkC1zL
CulDYXL7O6OD+/m2pCUTL0dEZVBDOuVlYRtJH/ZG6IWWrK7ZOU2mJA3/OKWQ+V9D
tHIZAeXZDer6oBdowHTR1hMmCPOgMoVKhAxvp1ahjoxZ7PE7VGSmu9Vo4SVfbsM4
iEk12VqDoQqMV07BF3/twMdtmgevD4km6As823S10R9XgfsFMCL5RBguz0HShpsj
XqnzZiGzTmYS6FSBPCFAwhFR5AK/ZKADI4VK5MshelrgsYF20JSQ7bela7Rho9vz
Cx7pdKQfvgHcM02fBkKFRJNJqh0smSlLWgB7VJhVajrx8xa5uxEr1JY9xE6Trg7y
9RfdPcHOns/2qg4tpgG7WABCZvIT8vwaxOcoWqDtFFDlrWPKcTiyiPsO0D3J5bAv
/zIm1gF7+WG04JY4T97Y2mI0B0uT56wK5Ob+b4vm7MEii/SelDz9mfwVeYHhwNmT
yJaYpI/3DFDf3yAorDnsfee/uJAy7SymBPFHvtjcCxpEkh1oj4hTtEDmtUxIMawP
ZByQT7LtMNAA9xfOW0K2D+fS6S5KDDFuBYxSbPUGqVQfPyKT8VKXVipZ/EEFGK5K
Vcl4yHkUeZpOLzJQU2XRtSGi+pWnGYahhywLBTTz0mILipV9Mgxu1KPgiHdMYMmv
JUpEuraiPBjSuR8akvXfINbFhEz1T3uNAkfsR2L6ai4+JSIoh7a27ytQPsDlPsju
IgXGRTOkI5xj6opgKZw2lTNpvHyCZBlZSK6VhLMssZYEUZd4qu3yb52o0udC4ucY
wPa3C/PoLmNM+wVBUXYdxog/KZxpiXX0ySN8xTtinWHKfOoQXzXP+YBR7Yst6G9P
MhfecOw8NynvESx0tLWQBTNk6oR5KzE6qF5BRvJmIUPSANgn8MKfxKCzIWqh87dj
nEhKI7u2I22Kwdg46WBsnQxFBqZx8qh0fJ1qggVLIfyA0ONiaKfksOWUXGIewGrS
qjg5ASyaqNLkSKNRzY96Njw4Vkq2XuNwrIcpsOOoFYcTqrusSawgXchu1DajBZ7R
o9k+H1PR6oYWrifCiTgXWyNURXhPLZTWPsxRVK3C7NSg33I64yBZoIjEp/QYiFIQ
S6ErjeOX5jrY0ayCq8alrJLTFFYIaPk92T/LuwDaRJDKVbC9z0inm7bQMBRfDucm
cpMSPhNyRqY4dlAkGgGsAXKxgIlcwjjWGpSr1Ca/23/wtesAbaaFzYBx7Tlep+mB
DM1sl963pdzppwHrR6jN6ssAQX0eFK43RkyEbKMrqXDbNrYyDEWUef6rAg+uCJTa
G6pOU0PxmJmw3nRf2X38YYfE2BQvqDP4kq1F7SCkWH9ZAJ1ffebsONvRTfHjL3Q4
I+x3KUQ2T72WVVBCC8lN/dnzSEEaG0eJfclsz8Dg7GgSlQZCdAG4p0svPkk9m+S1
C+jp6GPKYT/Zqvi0ShvsR8faPUkx6wq/5b9F8/u4+UGdBUVHzVDLEPvrIBMioDuw
kqDnORQKGGvcNvUe/7W2FEvN73UdhtlcPDbPqTF2D9NCH/7OdgQWqqXdiMWwU8nT
UIGo3M/JjpWt/HcfHbrE+vXRYGNe6q/RdrB7EjgxF7Z2+OzR2XzTSEE2ySpX4eGu
tdjJgOJFfrNu6d957IhywSP0leXZoJAq8CYXr8pDR9+PknQ6CGXhSPtjyFax3TVq
3fiFRh1IztUzUGg/Ex1aW1qdn/w8BYhexjtxakxfaxnHfOMeFKSggJXpbH++uiv8
3zJJKG1YXDkK4ItOgNnwAnFQmeBHEz9BwAzFEwjmUY62ovAZ6yLb1ywm2IfUBdwb
Y560cVlZ+Bt7W+n8jxsr4y+pOCpaN2CTc5TyrqXKCmYB3ybR9p7HzKhG7u6ge13d
mv3mT/AXTfqt65xeJ7utFkst7Ek4PXnYWnW2vkYws9azka+648Hcm5En+/MlF4FO
P8mUdp81ZiGrCbF9iq8hixNMqIHTBucLI/ZvFzibOwbfEztuC0zVdeZFNRN2j+MY
7hUMG3gksUwerLKZiulCeCOC1ELO322XeRWAkaxT8u8WaxTt49q3lwrxZyd4RpyZ
BkRhHLZb/HUIX70KQRbBOUiOnC+E5jWxC/WtM1wMepsKZKREJB/iSqyA6LZvKGMp
qoIYQQr4WgcS7yZhhcMme0afqxV2qIfiuel2j5tn38f+w4m+lSLcTR72kYXg7m3z
nJKvPOE+srrBX97t08ACeS21DQmEc0EpExJBqpCkjNPr98RJhz9Epd64lj/awou/
2awxjSZk8KdpQY8Ji84ZOUaClrY8fm5Zm8ytmd13WwMrdk0HjcqYw16gyiXjrRgo
yOFd8slUZCo2pytL67KZoeqb0RDE29cZSVQd6UY+HZJWaVMmFmY6M8ZfdGV/csK9
bIPgeDuXRqe8wpy9/ogpRTAmkkcmljFsYvOatlaJIga2KUe6wZGlk72w0pqSSs+U
XnXR1xVbHtpWnjkuEAk68EdQSGR2aHqT2oTZXdqC3CgtP1Vu1gtFX8cf0ui6LnTc
RIxU/SxWN0vXxNbKoMZ8H9Kv8wY7WIHbfyGoTFBMKXq6lzrhQteZBPCQUU5MhMsv
S8FuIU88gPHdlTANx72UeGwoMBSsGpD9N8ELwpkhet5Tm4s/U4UJ0sbLckXrHbIA
L8sURFSLs0wFjjkr1r59/flQ/vURdU5Yc9AG3Qjj7TUVqLQOKB1D7KI1/AncSOhj
5Dv0XLw8mPUpn+zMr3alV8zFspJKQsMakZqj7IN16kUK2GVR3U8BoQbHeAjVV5uj
Zc6B99EmrjiTIVZaKYJBr14BLRmKdBGJC+wUWepoDK+QfADy9Ns73OOuxIbaJx3s
EXNCP4Um650wPcDhTcZcbVvNKm4dnQO0sQHac3mScQAeieXNMUufymUbJceJvjme
qSr3osHcX85mNlFsSTF28j7jWSr/ya29Bdi+UCfLYCD+Dawuu2EpQAI6brLyC2cn
rpB5nU0/mh2QgD6dToEtIEk5sYTHn8HXzFb2GZvy76pTPJFiWBwj4NjU5ljU2ibP
hpE2UMuU6MuxdwnJZZPZn0onQ7EpG4fcaqQIGJQg5KiJuTPWpcCZDroPhjSkb1fW
kSyI89cnjh7iWqsdLXy9pq0GRgCO/HSm9yRVUbZXhVN3Lk0pLTS2BnVFEY8lkUFx
nVHuSl7QIXk6naJi+/bCoj4pgVmqJg9a/ThATkf9dxRVpgEDTZRhrqHvjmItsztA
lbYpsropcpdeSVPOphj6xISpommlxvYoOe6uMLNsnenV1fRNhEDtdVxodX0wRXsV
8i2wp7H51rRvhUM/jSkG35Bnj4nj+Be3iPWRLZbEYqnUoLv7uGoZ17z6OWjfraVO
urtzEGaaqIMymIziDM08WxvnIn3DKtt7CR2EDwWPmCNTFUndJZ89StRRLGaU8pxa
IUKiBu5dOejdocvNjUXVDH/VPSy3MiEnmw0K4D8T9wP28+0INqENE7nqQ+reEVb9
znV1ow0Mnz51fcMlr/QjqJ3fR03lU8tPZsr/l51VYqls4NnrxY9JgNOZ4I1YGbWc
q0OlOVFvMjHNYGS+8/mtn02FuLaOSlPbyQKErOKyEoGUj6LX1DYWBstc3hcn/Eya
tsHyhXe0hQmeeCjA/iENOQUPRxqPDpu1wEiL9BWMDQSGgPaKDcI797QXRAS5CEwq
peHAbCzIjHrqs+vby8TtR6gpzMYtCZ7XDjQEkQz6A7aYi83Xnx45M/RHTThq2j9g
zXypxCNoiWNsKMHQ69Ti+MNh7Mv4hVW9mkLDVoGKTXouv2UG7vzBcHv5XvOQ7SLV
zd7l0TPvMLzU4Cjn8KiUj7OwKnbpoAKms+UmaZsdXSXNrGUadT8Y7H+W8oAxA6cK
SFZP9pQWRpPOHy3zqF9oIeVW0RAl5tExV5lTNXJGfuH0jAG8bS/f/RRVpNNrTQOk
m4oQKAi74Op4u3SoQOiCdQCVvVcBg2Wo4nbvLH6A34Qa2Yytw+xgAL4U/K4G4EFd
hxIYZ8ahml1xw+H7TAVPQFFNbkDQXkzJuGEDti8kywPjwnIkhrSkeMqaREydYS3k
G+Fglo7+LMXu8SqJZuIzJ2Di7EICslDO5Mml1hTM5BmGx7QiCEcIlj2+pkoCX+Hx
eMr6LuY6rIoWB6KpRbjEaLS3H2JxMqdTcz00y50wvl9aWPN13no/FXBHHM9Rw96Y
dg84b3Y1grNxW6GMYx+bBHw3RANzSY5GKdYSmZSdJAMFYN4/l2fb6QfE9YmkHukx
kxn1eag9jMonXEFHKdOQkPIGIwHKGA5CZJuiE4FI6h0mrCEwMiRgCmAerSiM3MAa
EW3829/4kOUNU5QUP5iOXQa8yQ8jVWZWGZWWa8Y26BjolWEDZPnULTAx7Cvt0aRW
suW+zVyI/x/P8o7+XS78LiXqo/2oF8o/8IJy87ELdkQz5/AmGyAbAJsWizUVEtuH
Av5OTus6CVokfT/LWmobJByG7icEFN25DlDbCqQwkarEYpsVXw3Yv58ak0FRTwaV
Z/fsGaEtte1uWkGypmlKtmAhwSba9mJMSkhnXs8uHUgwxkzcTCyeZZI+9X63GPAm
LTPDBoVXWx9i70J20W3CfkP+X8mWlvw1lNblz66WDe37EXm+kwNMly8+AFHfMWcB
oM8xjySYM0IrQoPCLTXaLGlTXhAvtpr3cCuuUetGw0TApDfnc4BJK8B4u5L+FN+5
Ja6KCySxFAiT3jZewsElBAw3+6tq68IYePToVpgwRj5ZBNxoERy7Wgd+9qCdnX6L
M2UgXZXGDSUHV8GVuoN+q/cXUQ8Mmzy72+WHoo/9GVgk2toQIGqQ5RiRUviZLShe
gDbJTy+52aZdLd6zM8bGhqzdj8YwSt02oSikPN3yRkq4kmjVKrv7HXW77YIrkvUV
PCBX+24fnVTQq5Xur8nD6DxhA4ZP6swcJjp95o7O974UqSAkmVLNMuoO/tAIBk6A
hoo13BFcAxPzxPkqCcc+3v68aY/FxQCNfrPGCF0S2OgjZYTBqC/OU1ibyohy7BxB
0r14q8iD+VzR5k7ihkXka63xenBQQWo1XMj1GEZ3KUJq1gAJM/KeqHNU4sL9JC5h
yJNy7sjv6wKXzTvtnEm8ABJHXXR1daxEG82Q8VneagyWpMEuLxLbFNlU7UtFMmCM
j1bIMz1aYUNWxigzW3ysSzHCPiBGqb7gX/vSgnBU7NnWGCH6DiCjQq0HsKuPKK0f
XWqe4x/ktmukSy1CXTecNizivIvdogpf31mZrIYdXu7v2m/c3khnbl1niwBCFnDm
nt6QMH3L0kdiU8bF62TXM2kozrvrY10eCF44norkCsIf1xvFeRDybywdrc+6l8W5
9HWdEouJXbo/jQfYLrIy7C7IUxTL04n6Qo/zyCeFcStfByk4pVIxJ4hune7FYHP9
aWfQ+1eYn6r486f56RDs/ejoQN2u8RIx6rhhucg9DBiKlH5SofRQByKInrvRTEqJ
ui/jFiIlBZ/PYXK8oJqHs85yRuDRBNo/WvU/H9AAbZVZ0WFi9IRbtep67j/J5XYn
CrlYJujf8dfRfTDDHDm+0kwO98yEuMGB7WyWsaZV+xLKuJfoX/QTsRZ7xzY/hcoM
0mtGGsZah45Oc4ZFi5h2rkFPJ7U0k44kAeoNfQ7aa6UZEmhkC0VodTVxwfzPF3ei
xWXtxyfhREpENw6A7upIpMkwuJ4cmX6gh1RYd+L6JwNWH2Zcmzr7glKToSxcUwir
bWduXNcgzcvucZym13NVTgWmbmvCRKdveg9tpFymJdIzwopNj7t6IumyUoYqDLfr
DTJBpBKOhjV8TjLsJyTJLHat9SR0p3LY38Ut0ZUnl7Ce/mw4i77PlGtn7oqa7bQT
KkV1W3NcQgES5YZO1fkq5WndmrAdcCdwWrFpNkA/gcb86bkT6FmrLSEwpV5FskRD
4wUZyc4mT8RiHyip51dwe+EnFRXiUYUT+mzeiipsjqo5nLdm61i8az6udANz7Fg5
eqd/uHj5M5n36ZrCz7ios6suBL0wkhEeh9eYAaLJib3czFYIkV4iX5GUAblv/6h7
HsRfs+BOyT8VOxTTp2onSrAWHBp8sfIbefmWbHqtHwIFK8jeSJrbugbJLvncjUFc
VGNshbFWf9CPqcZvI7acUE/H1CxR/EtE2KWtOouwd9/NWOuDelwvw+cv7dXspcEJ
+7bv8uPnFyPAUrGEXx9yb65tuidVQ2R8s8MkyvMid8/XL8ItacGl0soEfi4uVYiC
h6RG81L+oD9EqR8y5nCd6wc13mVevMf+hz4NN5EGb8wnm69fp2qHtZzu3f4JE5mQ
EYSue02Ec9/Vgn3bM4NcLDW9K0OCVdzhprV1a+++40WeQeayImrEHetEgi7TTv78
8v/Hj5Py8FgE2XjMSR1MYlZ251xOSRgTuw/dfXk7Ar3fSWqrAhX9+uRwdnPBqr/5
jErAYQzyW1A9ZBDTfaHxnIuL22uWNqOZms6WFKvmudvxf3YZrxOtWDsstwcZvHYX
ygFg16jaPK+aNZkOaTMUK46ruJ/qfhvfmGGyZQuWRHgcpgyuTYziXI95AbsOK6Q9
nn3v4wSD6vrMKnrEkMAj3gN3Mq09JlRbgMJF71ooIUcZHFuYqk4hwQTh27O7jyvL
CZvH3b/o++YRKMUDMBheYy4n0AvgvLF1jdpmuMlPxyEqJYgKiKmNKMY7vFFJg4VZ
zmmVLTRRyfmm/2lf9O/nNEDhjOiN/sKApFP9fpSYDUnciRkxvCroHjW8e7HE5PgQ
pw6+k0yEYW3cSSMrdbjAd1nL+uegYApAeIP9TW77/iacKEZbJf7D5bhB/IFHo5aK
hBeblxV3X36DIhC6uSi9YTQYnS7/8eOlOh050Rs13XaA7WlqLQDnI+/W97v6/dr+
T2XOFrIVKpf1nlBRVOX1qHPIi1ei7z9duoQiRoekdofvm5gxwnA0cjkNAM7lSUoM
3SJjQ3Tt1AXGWR5Fp36Ax20e7N79XLlxqtFQGyud+fduEjPd04KGPp7Tt5L8M/nF
V6Bd03j7TiH3pRSLRCi4GDjEEM6pi/6dREKZQ6qjtI7m9lyEbMPdXUW0eR5xZ+uu
gaUREdWLw/WjFsEbStVtw7srg7TEVtr9jDo3hWvZKf9p+1rq4gpPJtcADLIn6MPf
Ku+73wCeyzxxPzRkaNJg4KTLZU30SuPAvl/NY0ZVWrLuzv7BIXbqq/nklp/x058N
5W2ktqBebeKHtrDho7PLusDLoaGJkWkgbDuIfH5FYdH5OrzEv0tT+vCWu9VNOcsD
TANd8U2I/whPAPB04rryNHTy7jsYcJdIHnimzJmD642tNjql/mYa9ZjLuM0nh8bk
ED67Ly5+zUCV3G8AaK4sb/cptGU6YbtoTZ0XI2cT9kn9rMXQfPq2IukNGEuhBWUX
8CY5Pk4GyKKf4XlaGZkZub00hp+4rRSND+tpmxeBFfpnIZV3wkGumdsoACKX4Tly
hHVvKJ0d6RwZCldq+P7onCl/WWTwFaUbwLm7J61sz0cdBjQg/5Udkod1PZcYPVIW
yh1aAQLlmFk9sFkYOi10bRUShOJrBlq+BKQ/auP/vg/Z32pWAaRMAeD2VLN336XO
SgBQpI5eDTOp9yageXXRK8FJhNOOEVGqmcwxpBUotZSScpKfr+zjw1bB4kdM4tjf
SRFHjgAlsdzFUIlgP6kyB6yWCxFsspk3uyoH3sj0WuYlDbVXLTwJqHB57KlQr2xC
Elm4pZb9/uLqgXRk+6p+7AxoXrDKrtU6o+qnrNLFLiMhcJeLncmDZ5TPomdhxYli
v1QZ6bp+bUyC6vaUmT7o8So46sIi3JgpSngVsQ7E+5sUxcPWazO2zu5VJw9fxRG0
xSZWnWXaJjY3AsX2CHDuwaEeu8/Wb2rhi11lGKpmtaYRcvNAucgwFeuXJGYXZBeB
+q6O7dau9jI2FHt6LwyQ3bpFnKBg9kjWqG/jpLoDtwLw58hR3gOOE9S1wcwURl8F
74xa/UPhmLYttG17eYEppDx0TiDWTbsn2tewBg4Me+PZ26TTlFhjk1egRneL8CIO
frHlyHDP2nnFw+2BwF+MXxKjAzY0P72kI7y8pn6gv900OHL5Ql+Dk2QBDyvz0D40
JeAkdYEgzbA3qAj2OY03gdYyd37snXaWNcfSXFY1q0CCvUs/mI5ZC7RFAuRexVow
yI6eXc6EcY7fOQDZCdAqvSH1i6zDBUMAUB4vFz3CgQFvdh9hWKVLpCFH29xAo77v
riK1OxPReQ057FpjMujOPNwb3bvLFmNQDunKjUlYzi1GqmhnCVnfCGSLktgwVPcL
0Bn6TfTOWg1uW3T0/ySFsCA4qbexavXnwIIJsjQqpZYSBQToY5mEObFCd8iR4SWB
btamdrefrsyIaceMFG2RnMXh2KM8vTCsLefYEaM0pBcAUXeyTdVvGSN2dMrTo1vp
sWmPFXw9wM26hcXGQrQWM/SRGR5IusJ5skjVcdQvURGSciWaN6w7TU4RzLumxKb0
iDdFMZUrwYfw8i2cBoGmJos1u5d+0e7TxU3iAxlR8C4VO5lsQn5WURmmwQli72Ft
LJAEfAcrXEEWRxFPKWyWdE9XOeDA3DRvY5cGQo6L30d7qWCO6dqknhfs7DdaB4kR
glC3nXrch/15yPJOVUZ60owVLBPvrTW96X3oyIWG/Z3A/6irCnpcf0l5sCemouz5
AI2p0fcAwmGFV4x0HHSAiXcFQDRMZRLz6YVEORGtyIDtJ4Vj65cSYcMZE8t2U1XH
KL/R6iXOUXQ12peKumQ671rQ4sUniG9vTSrDlnF/GAcfPRIezIJ4fppzJBa4I5HA
Wr2DNU/hGMLA1eMsFKJ6W8I35ouDJOEo4drU1fZ7zngXL3S70Wm39QNjxdKcx58j
Sb3PQ82x5RFag/WHzudh118vx4toXR4zbHAEFATnwugiLtnOHwVn+v0IvOfCEq6g
TeEM0thPIBJBs2RxPsxu3MPwOrK0fm8qEgBqdLvIlZ8M3KZvqZ60MHRENMtIwuKL
nuIcT1OjdPune8lUAlN/sD4gQ5skejZVU2X7MqiSSgX1owVF1E0Ie7RFfqcboQiq
VEtW5TblltKwRqr975dyFRpdYR26ZFva7H9zLn6HPMuCyt4bl7q+bGx2MDlshp2G
hQB8nGsEH50744q7TyUGYLfDF1Igcic363Y8rBp9w4XPmRIte4ulp4wMcIILgCBD
qVYtSgvpGpef7ew54lb2tiw2ytlBZCu/9Jv1L/epSQdA9W7CSOy8zTU79oa+3kpg
H39+cT42Pfux35aeGpaWq2Aipbzc+MtdGDgqlPUoobpe7fhqVyEKvaomd5BCwfSK
kLvcEF89YZrKQNz5xGZ3opJjiSrDvOWXmPv3mqQlq5vHc+lnR4tZydTE7obWdwdM
E8AsEDZtJKLXSc0631EZqUEpoTjPa3kCm2in+T2eAAQbOJTZkpnpyoUjoq7fJ0VY
JjQw/QBHNwwnCjVL3ztCFqECHbADNJesSgMQYyJVZnmPJXq7y8CdSHAZhIQ/dLGg
C03rkpNqd265A8XM8D5U2Qpe/0/0SaQrbE4JTCGRqn/zYosebZsVkVzumiraIZF5
pqQZ8sneMigfNVuHHX6NUsclH+iHh1XfG8mmT8QFZ1PFQIeXvwSDcxIbHlW0E4MC
7YMXiPmEKu+0+K4UbJoI3yIIT3in+9orWaG+WCg/prUOer41m5surAWg34rDUP1M
XwU71bptd2HtY+O+kzQTvEZAF04MR8tEuCyQAKmNRAqQh7NW8N8wPLlyr05x4N08
bML8nwV6nHI+CAyI8Slqcs7lD3r+n/tpEqBVr7Gjh3UUwuLOlmSsgsmnYOrXWMju
iA1AmNeqjfAyyR11R2qYSwg2DHb4vPkQFiZxH5DyfSI0+B52QM76FEMW13uZcJpU
OHPFbs6h886hIU9UKRSMLUFIQmBa6vxv5umtmvubrqjKyR/GgOEAFZF5m8lpqavc
XtDB8cxwd/2n638nqTOfDm63jzPKNjWIuy3KXrZ4UdFoxR9+oDWZJy1FlD0vJjZb
lIOtZ0q+dqd8x+BbAeL3RHh2UgLpObWMVuWXE7+4S4ZfDxaUGBRhIsnvkJi/WetU
HLskVUGl9JaoKU5NFt0TFNBMpO0Np8smfol00M0dg3vk8bgNtsgffcABZCYckIPp
ScoKaAEsBGEToUyRzMFrPYMxkNpHWfMihdfV9+7ZN5HUxIXVz5v1RN1Fetl5YGYD
9PqVUvBbejDP9u9TsXF55wP0adkyDAFijfx/Wm1I/RfsR/VvKOAA1Fe2mTiz1CTZ
sTcRwjuKwDbPb4VJamlfL54iHi+Poq6F3eHM6FXGOyXclDnOqtsc61EFrLbL/b4b
FHNGROmvklOH/2K/zwnYQAa78Eon5epbABRqL/5XVHfRiFheCuKOJuKKmZqgJKnq
kajSet20D2LoSEeDSky4zL/GPXjTHQOrx4xfZJRLvNh352otfPvMmLC2T8Zcjizj
L7/vdHIFFMFmWwlIYkFt7KNOyS5ouD7zgGkfcoSB2BGrXucUufTf4GQrRy+9xCM2
dJvl9C21IsJLDSt5i1UqeGB7WbnxauJs8mNhnhw6SFSLgbUUUUbn2TRuZtqxL9BT
C9aZ4eIaEI9b0hpwch5a+Wzf3lXBNykdtjVlMgqvEBwxWiJpY8Q/3/4GfIqqRiaz
yJZwRyNZwRRYYTCzLW1yMZIMt0prU59ACj8RBKG9aij0mo0Nk0EIBXKnJoOiL8bz
yTHQ0cVp323mqVrbjtYxvOlKMJZ1SNyyOASBTnMpFkbktge/1Ana2YsqyxQBIMfc
AWYINdKh0UnuLlap3zr9Uqpx/EFimvsRtf0bgiqC0CzcIrqWDhGLiA+E9pq9cO7P
E2HuCeQPgWov8HOW3uwSs98sJcMmkyZONJPwPT+YqXH+OTWlxaGbK0FC99VE6HiX
IQ7JCZOh67ESs2jnav3LldbEmP4tbs0IyHj+jmz5R5OB5qvsZLjn/9KpCgMmiV4b
Iat67B3itBC5IMgFUPbF/ZYhG7MJnk6IabEtlGhjMMRwMk2skg7xhSlCkHz+eGU9
0VU2i6c0XQDRVuUBrC+XlS5sby7K067Q4oxGZzKwhfNsMbHhovmY3p2JHOaKznQf
KR1DmHuKPgc7N3lkdqcrb0u44Ma0HYff8fSy76csBPU09LQ6L8rfKmJs6ADAI7it
+U1FCqIEHRGFLM2Ze5XCKiu1gBstbtRgGpjAPIr+JiJe8R/5tXnH6S4BtNI+n1wt
vlDBiNyx3MYTjIbrn9BPIb9C1MyoDasn+Hz/s3Mar9Iehx0QmZzS74Z0HggjhuIz
qesJEVh+K5ZJTCIIDkNMqZ6EtvE9olxIDcQUvNph3G0OCLkAO1t7xDxQMH3HgDhS
NxPIA5sJ0EA0QlzdR/W5s8DO0a77UACkllpUvMf2JYy23J+kHg1+GINauOL93qzU
O89euEIF5zjheYDDUS+zrRwL89rg2LEsoYh+kqNUjSDjR8k5AuIng5M2Nl8waTO6
j0T3v7hXNb6JRlhwEXM7TzwusLvKBsCOuuWgO4wabb3WqKYE5MTs0iyYs/Oa9fqe
33q/nPx0kCjjMxzKwmO2YfhZMzTrkhr8q5X1qRUkBj96L1EYA3Khjv4kL1qKKy9F
opuoPhg6cT04lNrxgPgxMyADZq0aRU5IUzp1YL6oAIMZwIBvi9hoQmkT/M5xkJQt
l1VzzuIxP4dXRkIjQ0/SuE7XCnfwpZNq0dNvRg7NxPm20YiVcLA3UrqJN9wEgTyP
CafW+7eGzP+Bjqw43JVrAwFjr9qsmxVhFhM1e3v+cVJ9A29vPF69cYG8DINYGM6z
iLFCXoPMh+z2EVoCdRUsp1HO3g4jOZP6o8YSw4TwCXSuuGx/eshPxU5NsOLgHYLz
fQ3a76mHUGZx0nWnSSNS3hDAU6onHUzsTbHzeUAh5XQtaeuXELZvScLawOSnuKLn
XZKPrgb1paV+jSxIuutts1GZo/9SIhHhfNSuKp3yqpxxKiE75Rxp1azlk/DVVn8c
ucRDYi+ZNrTlCluNMP+ZEWYCSmU1IdduGIiPawh/6qBpi2y5hlrfZvrp7Kn8dl+8
jrLp7Qhf8uNeD0oXt2tgZyrZ8t43bzN6DRnfSW3ygBv48/kzYHNatsr7RLA+UUmq
tv5k1egWZqIMxUnKP5MPDvILEdHdBN/uQxBlTjpOxaKCSI/8ebztX90ZIA9fSr8s
lo582X0tQ25qXVmCnvwZhdy2QXsfJoLEHO1cbOl5X8DAWvbgVjPSaYcEU1gLUdHj
xR8eCc/x6XRluFNrTM5vG9eL/vxa33Za6njZG0NxEAs9fqBK+15TBuLrmqWg8E6v
sZd2DUByTB8QbQFUxZiaBzw4MFW9leowLWZLqp2Jh4BLRjJfIpopwwrM6WpTgqq5
r7wH7p8B6drFWgM21oRagE2rqSd5eNRohLFMYV8rfporFp+Q9YykL/CMzxqF7DQf
XDtV1YWjC71uQzYGIuBazYLMWFeWXO+8ysWVaiWxQqqMK+Nm6crY+8CSSrky7cP6
0r1xx2klXnf07dZ4mwDwSDEdvrx1ltXDn4Nw7pQKlxZhz3pCobvZ5l92ZOqxLtC9
eSLIdADuQFKpyHQfuUStkK+Mjo1UR9VrXZzPRIrg2Mm4cIBofKYn4qjCRkH34uvQ
M+N20bK2BVcDruIG7Keu841J+0domisXsoPooZSYg8/ZYU095DmzXOB6BVr9H1Xz
Te/BSDf5YrFBuIIXEqWNz3TsyKk7g5Az0GJtWF+LMsNQi8fewRxAKROaXXV6p4nP
B2xm0VXJVI11JiYtQdE762P2O1i4tcqj52DyX/83bS+LRxRQE7XaDU0eMkNq9W2p
5wptsE3FRF5Ln7OSAx+60upFH6y3YjJb2VPamcvAbyP2lfjs1MpbQwVRcqRDpfoO
WGdzG4SuCcxX8MUTQksVEKZw5wUgCT0euf377UwIBsnwsLzVw1TdbF0CZAeDQVP/
4skGQixlt3pq5DWyNKHDk9DB7D+OboMy06I60OENDZektYlTMCFU9orx7IJa82l6
ha9yp/CW2snP5fp9TXGcxG8w1xkVxe32RbMSAkn+Ud7Pejh6Sf05gnxS0SGRjmwI
zKjZFI0Rz8aYpRA+XgSDt+GmEFsDUjqxFlRosNYjG8LgaXyCtqaMP/m4SyxsPxUJ
7oYHpkZ/4rGlpm3Glv8Tt9w08seco83tOKDTPSdj/rYY4HFgj1x5avHL1fG6er9O
K4TdMuZ/lklo6m4hGEmmF38/RiJwbOF5PJfIH//Q6ZXD18xhPoOy3XLupQnxQgXy
tuaGvQB4M6W+eU1+HMTMKwl3/EMmuhWrSqXST97T9WtOzv0+I5uB2G0Hq8JGfUB1
yoJDEIpFVg2UXjN/TWM1sD722p2XWxVpfz7gFw7DxnZBT3r1VsXNrMSAAgmSMFT0
QNSMVzx20v6XVR7pY/JtjW8cajSsn4lqZJm7gOW0D5grFSa2c5hGIE/qpuZWmvMQ
bV2ydJN4gsc2UP1umF4lsPBaBLH7B6r9JB//1W2DyKt/5ecxmpOckrVTxSZVLUPc
89bQX6GSeVFouAoB14YPVTUp3Jm8af38X6GSLu26AYNRNi5xHTo7lels2uVk+Pji
dKm2lje0aczByS/meSLBqL4EGDo2H23JTycnzlqMzY+NrN3Qh5fXW6Ps5qcXwZK1
kWIO2r1UqZ4rWe9HRPdVY6eB3Fg1LfpYNcDTUeDmi6vbj0aH6LF4xiPm+o2pcdol
JbV+RZz1T9WSCjUhA6GiB52+A9n0fLLAYaOdpPqYBWgqmmke7mbXuO/nchzpoiwL
WkEje+8BtZPOeXvXuaezmPrjtVnjQZiQQfta5rH18VCVzV1M/n5KEp4UCrbH7Svd
wVDVFLv3JDYnzNMBg8Zzt/dO/VEwPdYxkpxjQdttiqHFkOm1RqAcpsBSmQz5uFrK
0z9QPYMF0H+xaB842ZKzhVXgbNKgi6cvkMfpP6TmpYIUBqo98zHac7qwv02zKtms
4h+oBNzi7J1YXdz9VD24+CARloY02y/vl4vQD7DY+TuBdkGs37c/tbl8I1IC4X8W
ZMkKmbO7ey0VmqL9yDPp1HU5ft0oMamSPOqU4z9Gtmfvbq9OK3deJ7sIrNMFvRHM
A9aFS/flHc8G0paf+axDo6Q/VPFS6pN9FcNwZIfS6qRKr7nHyhBUBmfIoVyz+7xn
GKNl2+ZkK2S0XlQQ9Lh9mnlrOUjpEoV2iKmBTFUnpJ0CGMO+8q/8cb20Iy1i/Iyp
PiwDawy/DimkyuIX6Ro5qSvtyUneUKUAucnOG/Y1KNRzzXH5eA/J+0/iQitUTgNO
i72sBDhCZDO0F6uhgrmpLDPh4OsQNq9UA3Nl1LMZZq+r6OYp0vtahQgBsDqFCgKk
kYJ1RpUJ+NJnxQbZnl5kSZSWGOWx+bDYHjuu0yZDSHguhVy8lcP2gGwcQg3NkOh1
ww1ACmyiYYFKG4C+gUhrMQNcbaDufmsXZ3Uh7pe6XpE4CKLls4ZDZvUKbojmvZ28
5m9vnP4RfYQIGDGmzmsn+csDyQEnRPjB65a/kjvbu7IJHcEEoS2CUawQfB5V6tqI
NTzqPMrunNCGz6RN0zSh8USOOD2LvWlkjiSaEeD7w5UefrntbUOzT/9nnYZXNW0L
5DV0i5JYId9AotAQ2aekdqwzStN0dLY90BMSzXdy9TH1ebVL+dZjMQIseGW4ZjTU
r57BJwJS+ZFcpUXxkfkceSLjZBB3Kk2h8h4RwFcwbibbF4MU5x+LGZFthih3HCCs
Zp+4DHRB2tQ8e2M8IoyDL758y0/uJd3Uof9LPu/vt/mh75i0PNK3fx/Edht8TTka
QFx2vM2gwF4+sLxvhpzduqfsUtmaqPIkPz+NRiVRXyo4Yn9AgKThdsjvOhqGkxq9
PP/s8ZkbwG6/y9Hf0PDoWnkWTwjmTpDvOFQ/zSLr/F2FnDhmUwIcyV3G4ujqadEL
OitV4gr0gs1mN+0ril+6+44Nr9L/DNu2NdNVEsfcEOIBVgY3HZT02m40GJlOGUX7
wUbqlubizCeama7R0GNr/I+UojlivAWtOVw3Rob9AH0M6h4IB//lCkWlHZ7C5ip5
o5OPXdVZ+vkmdj8s7IyqpOfsU9DZNtLxSjDID7ZG5loHnSNmnhpSpekV9zbDtMzk
pbygzkWyiWJULtAVi9vgW2DWspbwoP4FQy9ejD/AC/KYLEKNnJ+NcHtcf5qibh1d
/6cVYHuJkZVErhjMBCWpj9k7VlZt/xmrsem8HHwwVg/Pw2Y5oFBVgxMcNb9JooeL
hv35IQI9dJW/RdH89V9XCFyvSvSRI0P/+SsGvcXHlGLEe7o25BCuxbHEvEBxGOPf
7j8LPNdUHu7KqNQz3gCXzWC5GGayjaruPF21CUFndq6/w+kLe+CAZn8IFiLQ0UKi
BjCQz/rh6DGRZMNlJ33Ja9lR/XJB9VMPZEnURZHKib8iyBsBURhS9aHeuH77kooc
x6vJhL9TwuWq2t/+AWbGBobPbCu+9nZxuZj2b2Twtw5sRPMly3aAxi+DMUBQMc0S
NVoEXcHT5tiYSIattszc7Q6LZvJhWYNiF8IltaEjDmm/dg3cITsxUC2iVGUyo3Ut
SSlDPyzHkHaKWc0NDYvQyCsDzed1gkgAvX1VsgujwaHLCEBkQd3JQfAxHBaIfAwd
7RggQL8/zN0Bf0vedYUI9GrVEh53RmVXoUMyqwLOBbXI+5e0arTFXQH6k7ekaP2J
4gnXucPJqFAAYCwEuaCxSR1saT37gRpK8ZoC3iNbkuM9Ceswre297T5vunj9FcrN
JsWHFmlp2lsM/HA7D2gXGuW5hJi0Pa7+dMQVHMjjheYsLYfM9tGe1Be40/PDAKaQ
USNePH9hQR61u/whav/MsUtt8F71JClj4DCvwuGcHx4Dxgip0OL7/c8ZJhSBXDJp
EugdEILCzSAwLTqwXLRRMVVH3cF5rzeVtKNLHBtlSI7q73iVCI7TRA+HxMxQuvtW
E2oZxgQtTauSyDCXJGP+AOz+huWFXczp6eVYePA7lPeRV8fQ5jBph3OMihYMg6nH
6X5jLIMGZS69OYWZRKlcpN6boJgYXLR+K9fKm0qHiwgFiRyIOny2K+Jy7DAznKdK
grWgR33In2nA7ajhMjgR8p72e9qsWXcz2pepoWpJ8keKmS5nZo7f5qyULkFP6Dkp
o/C4jsEWa+7zNuPDiiJwlC/MS3p/wO1aby06zwMIMrvbruv42l9o7ThcL65W2ywd
qiwEa+FjdS+2pivk18N0k11Jp91ztmrg3Su8lWOyj4GV/VR3rrGram2YzpUJfXFF
QIeElRUY2OcSuvWsBHJmc/RyX1pgC1FWZtD+M9tSeIsxvMcy+jgNP2P4kbvCTHcm
UFN7rOZpxohg1vt5U9dZd3lV8UVUFe9bscZBhvHr9wj93pt0hiGLGscGPHBi7v94
37c8iFeQah7EaA6dgQ9Fgl9spEAF8mqq2zOlsWwUh4NjI9p66QNNIPgPnzIoeeYF
jN+VcmNNuubmFwvEgDvjt4WddQqDzqvFTrasJdvfaUuWDjzT5vj6wO3Q7f46wsXy
Yaw40gRk6jU5SIhPQRGbnIRgqX2/BriR6m/1GWHBhhMgmE7q5PC+A/BiI0rzYJHk
cBfISBYOnWveiBzQfHnmLPCYH5svkToxRVLYvN8d3yh4+8He01YHR23kSI670TOl
GPX+R1G6Zy2IXBUllLaoOD/wMOyIsRexzPw6qFrqVic6A94ze9z40tKn98RRAh32
4HQISfwNq3MIwxAsBx7FVahKHMc5T3F734IXOK8oob+om2g1DTE/LMoI3COvx/Uh
IuM6RVGgz+OSbZK718GWFpnwkBTGZohmBFXKSaiLuaWuVLaHGTfuj92KJExtR3e3
DWsy9xV8SMzFd2JAflE8fvVCc9AWJzdMZvpRsi8kM0CoAiGZ5k9J4/HUuI0HFqae
7WA2QASrXdWTso7l/g2e5rth7yJbt0HddKkyVhRog9pNaw0oC6nEJJGxze/hrDHM
tRYWqWShFiBG5qpAivtuRlwApSz2yH0gyUwp93TjNcfGhZ4q8kDdfKlVGMH84yVq
a6JPVt3MDQfUTOzxBhmTe7mnecmuq7FAhE7+yPiy8M1Li/NIkegmp4ZeNPkHWcBY
X2oyaODqD2Seq9vn4NSfm7y+JvWBdet6QWCZ7YZ0pOMr6wfZ3r7KAEeT4kR9tCq9
NieKSy8rJgoMot0C0FvkGj6WvLLGBPz+1kEYKvr4ktBMQ7cf33sQalfK8ObzcJQO
zM6WPqrXA5Hbx+QFmGCPcyE3RZDXuo1KrQWkiRrXNlMCcQDgxV1xLs+tvI8A+Wxi
FrMRcmT9Scvu8oJs3lHOLbnxJMI/4rw8vfRsiKzlIHqlX/jxFZvvJEAEqQsJY9A1
dqls12G6NXMNE15ytBuEZn2SgTSDmF89iDrpPbL2odzaVFxQ5UVk6+5HMl0t7R5+
HT04oB6g8WQ35xkhBXhjv2qT/836UpXBwqJXvtaXAjDEWw/a76EpKWJtKuroIaBG
b40a9hheryqBUdF0lOL5rXgE5q6+bvmCASz90rqhytwf8p57jaWNrJmugNA6kJgn
hzvfK3VWUql4zAl9xNvV3AL8l7FUs1zFZP/3fJDUPeN1rZE+5RqUwJsoh32wbqzo
1dpFlZCOoxBfTlFQaCAMHe5WCkF3QR/oEq0jJrA9Am2VjlAWGL/Q16Uq+vPnHsPp
qWvUsCiBXV/1fI+/iK7SbAYsuziJEun7oJQAnJpBktxYH2CUjR1Vr0GoQUP2cxv1
h9P0ZFgytL8uMfpM1jYahByGn7tkLtpa2AwC3L/E7LY6limMN2VR9e+wPDoxN5W1
8kKD53+lg+rdta7PyH5wFJF7f/y5WDmlqiT//0E2eOPt72u0SiXdER/agSfe9d87
oMP+uA0noRrt9BbslzcP65xmpG/0fd4bKs0ZVn22rtiqH2D7yBWAF+bD1M2mGkQp
jek2xDJhBmlQ9GMcryGZYEYfG0oOEhCOxQO4bvYHWq2MSvNZVPbNNUARBfiJywiR
NYvlc4rgYQ73wdtiwRtlCU5qbCsgWpOFuuuPtnJs7yvD6s9TmLoCiTYRpFXFGFZ7
HTuuBmD3flgE+11Tqzhjrf1tqO2CaJVdlHwvX8Z022UWKyzwaIUbjy65160xuPlb
VEcCeOrhOs4kWkvCWRnDgWYkRdk7dodyiNXNvZRGMNeGOc4bc4SH36I8kOwA9aUX
aKJc6ZKBxNJ/F5DZS7d6uiE7FvWFO3h6dZ8GqM9f2fR54tF4t3LaxkAgYh8EpKZp
+yjHbMeJk55niaD5MP6LWkAs4ebgvSfJkamASTwPqks0ywuhdIvkYrf7UqLduNDX
ucbmqi8fvmdO1TybaZRIL4TQRQNBWUdZJcP0dvpJr8E6Lt91VmFVLB9ifhBh5gLG
FF/aKKhg9ZrJi0vPcMTa6JO32DFczTTJ3wcL6uzO/jVlCZFMTyCCYS85gw1ECI9W
01P5zTOIio1xjvdM5MRkuLffPopswUIG7JnX2XJOiy4cYLrpCwvpHLCn4QGyU2He
Wi14yf7+xOuMkYmaoqvk9ZyGzBO18q1Ie6tTEqCaBRG4NIq8yUT17bbYglLHqGuh
ryG40Nid/TEnaViodyMawjGtwN1IcoB5Xr7DKBjHCxcOFgj53V0b5XdqGMwSzAcs
683N99pOXlCFBkOmYo51b0O2WgR/macQaoq4BosIF8Z8UfoKRtMK1e19dS/yl2Zy
8JlIr/UEPoEG1oG8gxTUxkTT1Ocyk/8PcPtuZVJc77cB1quOmnrJE70arWB2Y+Zs
PUPrdOS7i46q9gs1pqYieIqgBuHXiEkwcyvzExOzH47+8dFikyaUL1xZ7+B4yzfX
CGLABaBg0WVyW3KeaQHfDNZMiYLa6A/85gwOYOsYfenNxYpwyY9WUHZLjCZAFWSu
SPdUNVVBGir6+hsv9rH7BK5TrRkCPe3n84+MJ5Jprxz5/mz5LfOkZOw9a6/uBjg4
G4dwLHUJ/qFK6edIMcNhICeFHfwhdCkNG7H6075BBzfXYVDcMs+1yVE8F0A0wQ1Q
oMc1YhjbjfxECc8X1P94HhDs9l8/nI2YnYHuy95f/Xx6P7GOtNYYOrIPmfwugM8w
ieU0F3OuynRNSjGBFy691Wesc1+mdAD2DB4Y9PKDCoP9H5MKUdKwqG78WqT0g1eP
SmUT0jklZpbJgMzRJGDZnx6Knxspii90QYtiX/gpiz+ZCKSc67hEiDtcNXlapm72
KTnRp7LTuwv4nGSWZDgHXGOh9qiM4dKp+RPSERo8yW053VVmpeff23bBBIUHz8yn
1XDd+gGlve3P0mwPWMrIRW0XzXEu7MEKKK2WS9DrWW9MzloAdSlH1zBqSGrJ5IJ9
Mdxa2+AtE0V6aDqY6gxdPJYUhPXHhd7KH/Q6ZvoisNsqHkwZvi/fFjvQ4cU3fwYC
zBVXw718ZnZrOPtwHT1ySXuT5KrbXzNexHAcZQyudikuMOQSEqkNN9CvlVv3Tnrl
cNnivwQQBWDqLnB32CSMSqOwfBWvKwtsTPTmSdAdxV3AlmaZGPFY2BVCWjDwwTle
KXt5l0X0SulqyyOilQJ8sFy1CP1mfufRsBH0ju4p4AfOkJI69wYOEpLHqEDlMtLF
v5wMg4aP5erbpxvIVS9VGvMGJ44nD2u25SQ6walvWlWBifAT3TAy1naKjsHTYxHY
a7VAOUBrUGipx8L3QmJx0Zp3Kc4r1oLI+NEFHBmc45TEInDC6lEvyX8lhIG9i8WA
9ruty7mRZfS4CUHrjubiF3kCDf3DjE9GOqttIvN/injeX08DqeJJNGNOss/D9D/5
hUZo2RA4jacElqJLkJEgJkI9Mb2/PAmnRt4fo+bR7IP6e64gtC4azM4qJPHmY22J
Ox9uFUR44N6st97G7vpBgA/HQ7ava8+c6jK6VvoHwVPh5JU0l7VKMP02ql2Nsp/K
nh8J8rMcXMK3J2H7aseyPJmOp9gZ8Y7ZrXVYk+3Zs9Yu+DNrp3zssGxHoJWjMf5w
EVzBICw+r1r2BqjuTZ+IPghSBTuEPKh/bbE1jqoAfRttHekfDRU5vxuRr0XRDTmU
pdVUW5LMkHEi1hy0KfBj2gLtdCu8hCZTUpIEw6U/ESfqK292sz3i8QSxQXXkOCd6
xOZ8l3LDGwlfigz9wmMuF1t0l6ViO6lP1+dXp5lsRqNyVBQ4k73QPQiOOf7b8fe0
oVEx4KGBCD+QZqXBVww160gvzQzwW/+T1SoZB+JXcUYjEJBlQ5fGPZEaHrLm1O9n
LNdFlIxQE+SiSOs6zR5XJMrODTKiRudLMLiHLNRVEH8FtrOEPCY4jwxkUiQITAsF
/eWfsYMH8dzF759Gos4sDcu3rHWJKnCOFFuh8Zi7fTg7C6vxZlimFp+rZcWXO4kd
FDFh8S1lXfqnIBu8CD4j5EltCtrR7bmoY7eLYocru9u2h40lbHsNQj2XzvBhUC9A
o+mZbA56PQhddlITEyDlgOqP3HAskYCPviLQ9XzDANjXmN1qwshh8qHnPKzCk6Vo
8vhzlYywHBmNcHDRrtkOb/XuTYvh7+Oe2P0MEhd7Gc8duH3GK3mhLytdOMKXXTga
yspPMEV2EBuGDwNkleuvXIDjvL6QFOvesrsIKyCC+Z1ZXXTfo/c5MNqkZRbqpalu
ZUmRPMnWgwGXoQZZWlsm3a1uKaPlBQhcXb1qd9a/DrSjAnMKXN81pmGwy68fnCHE
viebG+dd0LKPrOAIctt2kt3YY7td6Vd35Ow121pXpu8+ZVvLJ0rMVwqIqx34Lah3
5iIJmXatemgqinLorpeW6DIhZgOU4y1yzn1eyGMWEJAvAFTgDFjpW1zMJ/zYla5d
obOKtbnfe4euGRda+qep7N2OKacxSkE3y5T3nYrkRf5VmvMhxooG46NQBBP2VUTQ
SzBp9crH6bGoweux+xepNkmrUxAzZ0NERWw18iiaV/x8euTpCZ1ZQmamQ8bhMP1+
upn5gXUETLYHJx+PGAO5Oj7A27j58ZIZd7sEXkDO8KwodQzkoA5m8QxsVVDH8+26
IaMGBw5nGlrKZXXVTZczqLnqgbu4lzKqUZyNndRGlhh8KDDuWp0FO5jhbBb7hhRC
uwfZ1DRTjwjILpCsyl1js7G0wtyK+4N5T8RtOMP0IbTXxB/2nJ7WniTdz7AIKa8D
B7y5KAGW52Y3oLC0TDx8RGkkvIpe7nTJb5q/vl4fwUwp+dFBU5PbZfMHv0xXYrem
OYg2CrNJnYlod1SbInhcP4TlDoCHsd1w1yIEdkMYJ5/NWX6rljlOFfp7buGaJ8Nl
2D7i6CgbwyMYZyL3oDv+7wOCh81qQXguopqHYwHZdtWRdRJH9FpgNSyqYxI4kF2j
TwAyF3Bqze8djm1SX67snU7qJMcEteNDkLYCccS7LXJSP5lHHBjdiFhohNVGlQaH
SGqSPFeIZX0AXxz3Q/mc2c9iRmWtJYUuD65CfKp7u8b8iT0OoT7e7o5MlCGB/Tq1
G/ZgbShrtFPi3WVjMqMBBuEMNYARmaYBvvlHrFCKPYWQUexQLFv61Ls4NrlAnG0E
oF4ZIbZIxdZEQ9/3mOH/vJyRuohXpUxv+tX1wlnV1m1qy7dBnmf0zKRECglfZkkh
KXXROi8cG6Sld6wre7VnF/3NUBEWmPQCe3Ck5qYls8rApFN0XOr8wER3lr86mzMy
ChKEYWmijTST6rOHIs0BjlqUW8Lh2sIQtpNZpicYxvT9En9zlnCSeJpgtSpz1Sd+
ovvQVnMnw4McaK9pBURXUsAig94iOMqfIL59CdECfSUF+xmtPhU2CNqxogmhYtxs
dNdX96LL7RnlNpEOfH6fMiYelJP0sJc6ag7vNscdycB7Fv2ucfUDX1o2rssWiMvQ
71wn6JpIL/yOByofP+fstAQBlX21+BdTECMT5f2YjssqyUdkly9h64c2J7JAtXqa
vEuuLkGu8M41ec7PDzrnf1WoFrKbvEYLQYQ+ycJ1TuEqmsMKjsoun5BSQN5wryCs
N1V1N4F4PEZTNd5sGuvg7yqgVNdvAkDWvCXT/7IiEEe4rH+26Pi4zLTdfyL3iYTt
3UeAUNpUrIK21WYP7S35t8smJDefSRSniBeiFqOKFSRqDQIERhesXQHnJD0Ftkvc
RiTbOrARjRy0fYS8fe1wvmfS94YuCF6Ikk80A+j+ie2uL3tYNmTU3CrI/hRCYnfK
wE8JF/PnHRt1dBHmIZHstNUphcBHAHaVrOYr6QyARQD4yGU+xapElOxAFmHlvqTt
D/jWKj6FzcF8S4DCjJB4RJMSCLW+BjM7MlNv/9IkXmRNcu+hUVBxeQk5bAt61XMp
XPtXCgefS4MvS9Cl7VFSL4wlcwBDTJANHsll3u7qjcVgH9ZP4dfFL/cazBchKhFy
NNgFpIIMHAYFQ5QH1U2JciPb6UP1ppMVypn6c5Dz1+w3aFJ4CG6Nqpwc2rY4T8Ls
Pq0Ai5r0xxeGJMDsHskBSWcEZMt6lis9XSXeIiIH5SLJ0F/ls6EbfDAusE/Y07aV
WQJvU33ofhUCNVd2AuGZifqWgpVNopwP8XtGNSBoaGp2t+clkepT0s/wyMiFzAdT
I5vsHGlDM1ouzavRhW6dAR+WAFEIS9wAfZ4qIPGoYHw5PixgoFiXTXiZVEwcENzz
2Mivl1erhZYbsHQ5AmhVWj6VKRdDz7+CSrXcIt/DVqBlge8ECq2jZcPLo1jY05g4
x7V6p71LwtmkoC8jxVJZqD+G5EB02pfkjDEcKGfmqaBbfAMTS8Waz0bqS5mRvPDe
Thlvb0hMFKyPRE/2SrqMEFnJCjpuZxKJNxxDlJfqgMPQffYnhsiCu1y7mjCQ5gdg
WcZ5Fug5fI6x8uoiTCtrc0aNcZpDLSbrg79/rQI2skOead5QccZ1RdU/5LLTsDLy
fy3cWe4r7axN4appn6DPyAESCKdoz6+YnOGEoTR1C05WNV8snMdTvJm9dDOHlLB5
b968voU/j23lWr4qeDF74L5VSD14KETPV3tsaHxX1wLxIeSaQn8W2A1SoR0QxJE2
Mt6YbTKAgeWhiiYbtMwwP/nl+biBXzdoCM9e8Oqo7NZfLealG0YPJSBMLuBqlbYF
wGFBVlizga2A8k4MFn2xHdkTlHduJ3l4PxlNugmucOQNK0UPYhPVq+GLQuPJt+gO
vcDfVbeUYitnWYs5sWmmFwF1HzR4L87R+ObPk8Wi6Lf3MCp+SyheeYCzS++Xhs1n
tXqXsoVK0r92NnZxdPH9bN4aKXKkSw6N/lmdKCGk5WIlymQSB0ODFK+AJQjmLgiJ
F5HyEEu9UcYXWtlPOmavliZDuXFnwI2q0EPR7mi3o1Hw8JVgNp83vU4Vr0cVeYqp
jF6CNc8mZOnewcq8NXMgrzzNmz2sKtMfqDGL65WOxDoVIDQqLkzi9PAvE1CUPwtU
O53AYXapAL4r0xM2r3jheAL7YRj43yhefv7z3j8kDvxjOSCb4JQOkepNMNfzmxW0
SUVsLoz+N3eeh17E0e+A6WJkw8pD3/KCrpDmR50MyZFRoHwL3fx602ZLE8fHAmSL
DPya+Psj3dnrlB6w4u9mUuIr9YZjH7nZnTF6XzVEJ5RzRug/19oqd76DYVHAPBOE
cAZnPVDbHa3ubk9mnkvPX4G5G+JN37A/rtzs61jv8bn1xoqrTyYYG9c+YhwavC+I
Vq+Db+sTaH1QS8XN/fJl3TY1Pw1Qm+pWwVK34Dk+MQHwj1XzbYNl5uQHjWY5t3fL
yXr2NHtXI0mbwZy5Qf/B3CLcxU4KfNJm5txkN1z1J+Xw8DFerOgJpiF6xvAcUdEA
UphfhfsgIf+G+KS3nuCb6GrzFEsafOR7c2tUqz772S13nq4PUw4xuO4w4F3YVjQ9
pq78Pd09cUkOkV/6CgdnQhNJaA8Al17x0xTHXvBMF9q8yHvmZhSNVGlU272o14zQ
SRCYN2DrmCMc0mlSq/HsbzuBsw9mxxXuXEuaNJxjNOhkxVnlP8/EtoOIW0H57AZP
AOii+AbCWnDMPZ1px0CGKuLGVLleCETxHnzmZs1Pl/VJxKSpktaLfziJvMzqQkKH
Kqnd2LedLQ+DxicKJWSQARou56MwDQhm3fcyxKK7hxFQUQLVqLpKNJjB+a1QpqXo
Gsc9uVp2/fy313ZwTY3zhPaUgRy9ZDnmPlUq5dZ70MsRxoHCbMR4u+WYstc2u3Re
9OhAl1si0SetO6GMnNhHaeQU8WZeVQyZoiGOMNCvOUNs1a/GnH+WBSI/rXJga3H0
EnSYwnafvX1DT92NVlq15PX4YkrQP0XwKIB8qd9565j4ycLxWYwk1aV1/sjartzY
QUZQPURQgqbgKqcj2Nyy+0nax2LFRc+OCiJ/WDwKHsJygUQMt8r3sl6WvrCsVDBN
h9e7wpzk0PxVdnPH98mxT87wceJBZaSzUkkSJ9KrRZQj6eZiIfDpwK+5BT450KRQ
JIClVKhpxjwCf57+mwzgm7J0xYD4RtQhhx2Yg2ZBRNyjm9lbEXc3RAPFN66yoQze
GemaSriajjzPKMdXuaZrWB219Ni9csuX3kL+gpjFk58CQIIjgm0HpL+PSXhMRRxF
bXxBcbS2ZiiXomrIcdLPgPMdOMfhRkJ/BVyB9CN/94H5by0JOp3k3H2dxeee14uA
JRpXfAGifAg02n/1tX0m7XkBrXK/HHUOCV9PcScX5hUY+dZg0Qpgj0MHoUflSHO9
sVR2xKUfR8HWlEr3y1E3iD0jFD9cWwbLjJROYBmtT36xMYHOKwRPSbrOwpM5exaG
WzB0eCNCuaLTVN/pS4qJP597iozAzTrsac0UNMJDxTXLcOurxrjGiAq16wy9j/c3
MWGcA3Ox7zmZ88kPMGvRMm8Vhzd1Kbzlx53k5bbwxoO2NgUA4qmfkBgU25269BDS
kY5M1Hnjbm3oTgan2gGpvejxTJY+OCRGhx9rOD3E7MWTCnfcsyarfvyPd4k+BJbs
YhUUgYwGwlbTTOccnp33v9ycDdSMDWfM5dMlWAQ+W9xcB6d9CK7SyaNLH9BXLj4g
CJtaWvs1FGbOV/XdlPpByruJqVvM1+lP1KhvkXY0VAzInH8rpGG1zqvdKqB8i0++
g2Pyr0L2E64ipX181iXi6DrJBU+7er2A3dsOdFbqKq0ujbyLGhAU/6oU49yNrZmd
0JmJzTFLvIOh2VcJa1xX5vFVvT4+YjVBXB721zVumbuD2U/V9wv7LFaK5X75bSnn
Q4eKhzaA5Y7nRUcXKcjmf4gLK7egxScqBUS8dhb/wSSnzq+2r6Jza9Hzi1i7VrMn
nQCkfDhTgzXVv5Mpp6ix9Ir/9TmXkKl5Oh2ON+BwtkXMCf4IOh2hOVP1wCkjKC+n
oMvIe+d6GfJ2N/hK4WMk/TzJTdlXNzHF/DecIpigc30JPHwTms+iI3BYSVncns50
iqGqeR/NX0KLol0sHmc8F9rdSnPfIe+EjvcwYYGn7GmKiZDA42td7U27zT7NuMhZ
0GpocKCZrcOzg6lRNy4TlLL9QRUC2wOess4UM3jHN/KP5qDEXyUw8sEC+E6EehGt
dDB8FMd5ximS5UtC4E81oo8pOfvP77z3iZeqMtyS3ikm9KDayjxXyznRTcLyhCW/
XtL3aosdNxJTdE1Ke/HmAFDQygkPksj2AB9emG29dFxrvW/NcRbeYiVJ6zY0A0z2
egBQUdpxBWtGt8LN5t3WYEP5/dIc+5YhDmR7mT8dSnAcdGZ26qTgyd6K5em4J76+
H6hc0JCE2wcDG8ZROABvIN+h93Hh9+X+STJyQZqdZa/YK3jWPI6L4A0hA8ZmG9/J
vbL5B2KnqRqwWBy9qIfXxmNjn4ZPcnJ+DqV+K2jxfIr80rABKWvPmjpJMeZBDjKv
bZABI6yKOvDeHAVKwKIPlKD5aUDJM8lDHahHb9sJ55b7gPYwEEzvUWmFPWrLBqim
0kjae0UqWKB/NCbKmbOIOYzGCorY0MTsRgh2EZEhe20I/CGX5DndomufvAmTLnhv
sWV3yyNREXEUC5JAZnssVh1iDOzOU5G6ischsW9Hi5A19Aj3MuKajDaZzfErmGk+
tEfjgVLbUsoHlt3IfHLVyP3QeNZJZK7gshw210xy1jxvMn8dtN4M2ix9bgoBMdFN
TnAjj+qbkmxWO/WHFrAe1t/kv5AWfMzjqWBJcKlZiB6/TzpS24r31SlyZRi96jdM
vMPACuXxcmts30WKIUqdjrLuuAmf7YeN3QP1e6ykiDGWWHdRtUhtOT3/m9poiDrD
JCTWJ556PPSioA97YhdxrkfDEGb7is91QSOLuNmm9wRvBlZbi3k/IrCikMpHshk5
J985osHaSmcj4jC9/X2JbNQBvqWF+crWudM7s6FxNq/PgmDca/oQD+9Cpmaj3gYE
L8obpWgUlfLobJLPnSLASdW89jPhF4Z5r6WyU/VwhLwd3dBy860vcCCaTplRhPaU
/UPqnDGbXgyfI2IQxqcgK4FmWCnhfRLQJuyzyFY9intn5lG1klAFq3T3ZhlJk731
gxFw971+DGIlGtBLZoDc6M1HQmNoPc8f70P7Rat5MUvEMZb1lOJXC51dZIcdqJ4m
V2jwpSRgxqti4BEsZc9q1b7p6JDetRBDgMP2VS8tsIRAy0/U+zsHUnLwSpzNDbNs
aNyWhfSUFErpDBaPMxGmNP+f9YHlUDXKKKqhMgUaD9CVI1sxRLiTKMcEzBSw399n
TMoiGnfsmPoeTBUf9a7iohJAUfdRxF7FdPPlXOEyKOJ762ywcwzcc/0NLJLPNndb
s46ibrcPUA0Iu6IHdSYLbUQzGtb6V5cs5GnsvI8Lz7RXOEBgQJ1Jl1DzTyRHmQnK
IlBLTgE8LeNtWTVwMCEXRNcUNF08WkQRKUIFPmSD+9ROXj5nnNK09E9hxAIMTGLF
NNFPRNV2wcHNNC1Hkb2po7s78U/ehWCNSt1g7AEFAkk8Gttldvo7GB+irvdulvMn
yEmSwpbhSLj3pH+NOBWR/tQVdKhZM9h+1lf/AQ9uZo/4ZKMIwSNaUkMPyU0GAI1R
EILcwX4gT/soGaYWrbcqVRcgyvycZRyudBqtyKWb7VcjexmPOcJFg8oirug+LjW7
fBWFkCeaN7/ylG0jkWd6fPaw0ldLHE6FFNfcJQp1gT/eZe7x7diq3jcO1Q8msxlO
b6FHLgjS+S05v0nYEjZ1r3oXg4lRosWTmzpzF8euhM5Yn0A61UZP7UyogmufrqnA
utho/UQxb3vbtDSaOGtIcxjz7NGQC9mtonCuw7pKNAeC53X0E3xbRQBxc5Xea/vS
UVUi/wP9alqU1Qat2BYRn/H8qHtgqdIRsste3oYajsIUHX+G84/ra8wBzTWpLcJG
4xXuBsuFvLEbT1m66zxvti6XqQ1DyJfWpCwrhDndoCwrcxaUbSg0KOLNGD7KmcT/
XjB5Ei4u6UgwqWRCquWji31aZH+DcSbR9RJI3y8rME4DhvU0yjhtAFZg79varjRa
lWdZ03c63zigU1dgbzIgzUpj6c8dYVmO1OJjkOCw1o4Mvx7qpEIt9J8enWmo+bjg
inbO0v4WEKxgpcaZPazTCjGJ/koOcNq54awaQHBY6p5DQn6ehA/IV3p1i2sePfk0
jHlNXv71JZHTOYPCdT9EF2vohvxjuZtN+8LEjbfLzqhVsZHXYF6+ATdvLMwPcTEW
5MU/O8/94oMcy9ekVVc/LuM+TDMMFcJyin/ZQHJJdhD1K9GtczFrOqF+zfoDJKuu
R1ORNytjhXRVevVZaqOpa2mf+FEDEKF7QpojhleFJtuiG56/rGvlDjZ7bbG0jnoK
000HVHZvD8Hj8+1kDWwFM/PzDeEtsDBURQD4RK9CHDunWZlQ+REShJ4xn9CaZJfK
tqNRv9qgQM+A7EajAa6ZVE2CeKqj+R5r2p67boI2i/w9ZLPrtQkdr2gCMgusOqxd
RTViVYjqOwHDbpQZaf4eHVkDpbNGgojEXncoRBM+yoaEI9Cdimk/6g+c9Ga08U/Y
Mr0aXQOgpG4PQ/ydsspy25MzSIaJ/fJDhdTxsVCEDzK4S5o9zQRMDFED6OJh1a0+
7eMu/PR2wmBWNL+Oti2gMD2p7RyMMn/UDYNsbjIfWzpxsCwvJvKbKv/iE3gX+0YL
WZsK3lSWeFBqWb0Q8FmXxKiMl/poYTRVb+bO1iyGqKwmmwqvTUnv5b1XdIA6TTyd
RfzWsARwTVvchIIZ24IAKrqOB0LHLZjcn+ZHtErlElw3NtZTbAr8pI5ERUlrGpz1
1pHX6gcuA7m+gE785eXFoSSa4PheTcs9QEv5Grbvyab39ijGF6wGqlCC4NY/u8+d
XAUuPR6bGkwGAxeiINWs6QgLRLCsuXSiU4gWxKpzc+b2FIot66qgRGqNW636vVtU
7o1t6MiPTzfEmuAGmxySRffPyeU14SrbxpKtoAro2ikm5ivR7mKb5ijyzjvMJ5D3
yS4Z5FYbsJ4V+ITj/VaMTUOA3y8TLhYn/ziCa8iTpunis3ut8EKWC5iy/KCFr4k2
H/nkgK3wmFDVcnGgrL752+o87K2dJ84wOxwEcwDKYp62l3wZyps6vuWkKcdEEkzi
vtOrLxx9g0XgkEVo2BDyUJHlburN/m4B22BfUNa2kEXLMXBtsxorDebOAdQtf5el
dP4oCbkH67h1ncWdVFmbq8ZJaAwCkUAFBxUga2QEw+jetFTqNbX679gD7F/jv0P0
YFttRviQbVQVhX5ydxeirN7B5pq+q16mDKFNRxfVmfVS238zrvkrNda1VlI8tWjJ
VfNWHJD0OinpThf/lnN4a/wZUjz8Zhhw3SXp31OYOjd+AclDXr8XZpWqb28EES1U
wJeP5h2/DD766toAyTilbfrgYeatXI12ngJ9cFYqwP7w4dQcdYabbZ5NU9ge2DL2
2KnggrdpYe5rCci7hWxS5k8bVp3SR2CXDgEwRtwEiVQkpYRMQ/rQM/GBg1s9lyQM
VzjEFoEm60X6OVrUjIDLSWC3bLsldyKKtKKyVy0gfJ/6MfxWnD62V4/WcPN5DdOK
cVUyoVdgXvQvX+D4NjiB2Ght2/aXtqruZoZtGiYJvKI=
`pragma protect end_protected            
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
SuC47TMNpIehplDIbpcbJW4ch6W3uOzsELsd25vJXWF8GSUMnf84I/bagKrjjlst
LLnZ9ba1JF9Pa5o+MWqjbQPcZwoPItq8ehMAO+r+bWoAB0/5r6V0Lg+7XgYldVFD
W6VrkqozrU9GR/z46md95gVcebwn+yY+xRhMimgvUTw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 366476    )
Wmj0fJDv+yyTWOmv9H/me3beeqdLOSrUubFakLFr/3mdVm2/wNy38l6iWzlq5ezH
nKCeCwHqJrBc3N2tH0JwwV2MM7K7MkfB9uxiW5PPY7keC3QL7Wl4K1qBKyXW/m2n
SbiGQgdQeNiau0l+XR7BzZbKnG28MMwa8V7tZCng3C5ZA2CIqDo9eEsIzRlY8jCZ
+F2NXuMuNzHZ2gNxEOUMoX3yRTTIxgble6JibsyjEwTcO6K6Ayc5IJzdIw/QeSgl
o9Cyq2+h8Fw2LWEri+A9am1JGFCofWKMNa5eYPzhVsgH5vKOAqoJC0kQuqFc1+bY
rcr4IgIBlQ3kFwLWLTp25AGxa6kWwSFrcdWYZ40mCI8SA3nvDBoZ7CFs88WzrNhU
QZFpLk/nuYrlvsQwREWy+r5k/IxoJ9yHNYadNofPS6k0uoyz2KNE10vIheXNHDRf
5UFlRnJWVIMYi1J/PvcbQuJtpHectpWajp7m7cKg96lq+VZS8InC1YBsO3aeirS3
9UoIzpGx28cwqJ+x1FVNdDt3Q6kklZdn+9yrS4xjmaZX+cPPEIDDYl9P3fx7OJ7h
aOa+6b0VT54rLhAoJu/30m3HBwk04IjR9gbSB/mw0y4qwzDa8tjLZd3QmXxwToT8
Uphu/HO8FFvIfFuojnTd00L8EY+xzTKQhRkqePvfW1fN4Gbtt+XdMxsBnXKzc5mf
3KN6xMZa2ynFip9B37iYK9rPnAOlqsQpjrYw70JwmFGAq0+wv5vEhvF7Pv2cW24H
knSVz+cU8Hzn5AeSnn0wouQ4ydi4VsAfPbAYqIwcy2+Mh+qdO3PAydqN6HMRm3ov
lEh5kVX+WYRJcLUxaQFGjyrKtyPUi8UskTTokiFaAFS9Ala6sd25SpCOH715QpsG
NMkILfMRpQQuxDvTk/U2AtGHp5+StoyOUO2g9ptrEyNBoYCkZrCM9B8mTdXBjlhv
uBneix9+7FrB5Ep6IsxNrH4lOCA431AjJX5atxx1XsgzSvsYXBpRVNgL7c2574YD
1CV1Rg1SsDhk8K4r+F4eL/FkKZgV1XHB1BiPzxO536ut1nLgza59lgpesAFmpW47
buDrzfWWxUqvwp2C8hHi7kUSK8pQn7lxMEG77XyFqt5qpeAQrkNVqNjIyeU7j4JS
UtYgeAgiRmrGIrJFmjdE8zdLeGVVoEEnzzonFXy4OwsK6SRl/vw2khLlegX6nfkb
C6dHH0yPJpHxJqGQvMF0NPbn7qvSo85N+BHg5uNaCzPLLZPgljK9zd3mRulrR40i
q5j5W2Q1ate35QZ6FBzNUiZDQ+FNzByioiiBTag3Hjd5rzO5gUt8I4x5okYAVrRg
XOSwhTDf7iT71KPwodVdH6jQDOEoxRiCmFKNlzOyP4daf4X7PLRRdBvt1NFnR9ca
5hFiTFMrq2WFvJcqvjsV9ozyu04hyd7DsnjibJ2v5T0Y0Hb3WwhmB23Vm6pewnmB
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
NKwrH8CtfkIAjuA6MZ3Ol8vSd8k+3OFF513OrItR2P7mjxrzzAUi/eq5IaxkXRc4
NkYypm91GxqAb0a4P05lF7mIAOAIGTglmflo/2Oaujj5xdWE2qVMqrws0YrlHIxk
bsk8H2rgmHIz1U10JeHu4W9AsW1vf59E7ixH1bdPOvM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 378932    )
1eBNv1KjJVt2rz43jHi99g6L0bWp4jGdOQtUYU4HinSjl9B3jDgu9J265VRBcI4J
d/I/KVYqVfrudRb+NRkaOKFkm7RvMs8dED5r36DnrAmcJsO1ZpxfVwf+wuQasXNT
zkw8lss29zbFANqFiTfCKZa2JoghpyZOnV6qYrkAd4UlaLaXIuSE4D50HC8bM4TT
QelQ8gZJ56ibBpVF3YuahhrvYDGRfysUCAI/UAyBB2iBVVRzUDVEDWghFk4iBF3R
Dlj59lI+Jv6KmZVu8d8jz0zVqKlSz95YVRVECDusZTyXPzJiOSYUGjnxbw9JxFLy
/VgHfP4F1fjQ/jGJYIuKF6EEBzrGXUWZA1fL3jmTwtnLHJmgUULvuCSOxlZI9sW7
rF8rs/BVvJyAhrpdjQa6qxDvVeqpshTjj+WedDjdFQSqv658Zvr+ekYLarB7LRDM
XtSu1dH8QokE/w/XfTRBwUbMlrczvYCsKWqYB1AP2H4+jqqhyXhXam4To2XEVirH
kNYfU/hYoCZtemJ8uql+VkFpnMhfwfcuU3kZb0M8e1R1Jb2i5waazPytVzuqNYkr
P3UzfCBQbyZ5hyGQwmXMSze9YheFH1BPYsysRm9NIZmmIW/E6yQ/S9z6v8Rg7PTo
CyJP2sHhSbtJXxyaNbSdghHjoKp51Jgp3DXuWsOOeR+9I7uVk2P3UFPt5B12vfgj
wkA7NR4JWR0JaMeGgxDMb6vz3BH+Iiu5b1Se4P5DHTdJtuYfntjYOf61eA7mP6RR
CKgIBqwgSEriA925bu9+tkE1hrcIkaum4NaJoeu8MVxV4XZuDZByOtYAfr/rSKKE
oqhOK92qRSsa5+Y9UhYDk9JvxY80XVJR8c7wdCHrTSPdKnExjh48ZKD2LAfJ/88J
CQ19b/qLvtFtXygRiYzJtHxrm7vVYBEWIWidN5cs6xm8ZgHGNkUguGgWOQr8VGye
g8/mHul/M8VmtOgUTUggkb4bHD3sxk2sVNGbRjXJCsOZGK2pxeMhKYWgHN5+VpMk
4Ozw/WcUUmsBVnKLAdQBbQuxE2Ef08s5hEU80aP+IF3wt7pejzfK4Qdy/pjXiRjr
Uom04vucJMjtDwKUhBAO/+UveI9OwRXxpCK66Nui2W1BD7tH4RCOLjouShS6dDvQ
xcQhrj1dCdQy53QGBXI6x7IuW2KXnq5kntEzBn5kF/RfEW6bc/WrbQlyyV9ACKNA
UTucuxObinqF4jgtDvaPsR3krNpEG0UPKp57LGJ++Qlf4MhL77h3oats9rpl/AGg
aoeZG6wd//P9g3EScsCZNJi2LDVu0LVtqnbJ3ehs5J5XRM1p1sUkNXUwlRNvz0ml
aIR3ByF7MgWb57DQeO0DJX1jnT8WvRqNvuQOuZgAz2JErJGXMeLW2+Bh3l4X1AYp
Mdul0RUbpQRVl5htoBOqpidfP/DfbOPsKtck1KGWKaQMyKQYyGC38NXIAEcclvAL
7JVQrjswZ1jCTQiYRSGBtzJJJ34XnxNecA4h3fHeCruWTHZLyR5ewnu95/cr0pZa
L3bi2eOnQUyMp/tfKN8mzgTra7uBEMxJYksFJ93Ev2lsXYxwJre4YVgB7XWlM7Hp
Oi6C3Tr0r5aDcztuBJwPrpPPv+AnYBDXBU8kN02jJ7tX7jvnqWsPbKMx+PAr50vQ
hSXO492mEfJ8377kk1jwl6bIAXlXx3kn365pwj9l3PKYa2WHj9QHyg/5O6Rjc6my
JEBLethzea1vFl7+1gu1rlK5iSXe43g8J87uvchM4MtzHem9y8QykKLO8Sz8QoXu
ZFATSofXFhwKTGTSw4KSFZA0jvmtTb8/h6RQvWKUT0tqdWXapX01NrhLEHwS1TeY
bkZuKRc3rec3GjlG1IxJ/UjUls4A069kmOcnxfhnNqfBZooqskhZ9mAU8UcG2fS9
YuTmu9A/xvRNpowfLNBiaGl47FEVbyFIXa75XD+vvoPzirgJ11GEvUbGui5w4iyW
OtUVuHZ/5d0z0Y11pdVH8p9PcGr+gGBYQtW1az6uTfUOhjakCm/O+WvIlMT4iQyQ
cEhgUZJ0NZWwhvwkRgfgUiv7sWG7wN2lbCSBwy5ugPjQTaH/8veE0uw/Q/xSf/B2
kgFkr+/1KFm532rTxPK+EH7GxfiaQFo+zHWZuwKN0WzleNbPQ8Kc+c2/iUfz6yBC
WLfrKP0tqJ1/ZwmwOxmhIDbVvaTP/HiaLaBeTRgPUcJas+snV9aZcgnKye8rCEJ5
uyKVglR2dyzZVVgLv4qJg2Kbcu0QLSIYp0SrpZvuGE4u6pBdQUg5RoF49znaf/tF
vlyYH90ptmp1bZCUTZEtqZbLHGL/rnuzUwz1lkvXI7hC/wtLbGzoVRlXy2ZNGMW1
I+FPS2bFORar0mU8oYx5FFVwUE/tAB1X+L99gPKLB96vLBsHmMT6GKNk8hKlgZ2j
aPO1ATRBqga6Ur38L8sqEz51qMKvh6McA/2I9KDi6Xz0XknjRm0nY75nY8BeBJa2
5Og/NIYy6dmGEl8b3GhewVV+PcVbDTBmYPSd1MVXSVmmzF/sSDpUpa5ibmiUfQ1/
oRVPPBXbW4mDGXr+BOYw1UlBDsCjen2wNmJXAK/QwzmsbGzvqxJ7IkerMebbxN9w
jDA9bUhQv1J0al4MvhQVdeMm2DohbH2nvuX5ED2+yURU+kyPpmSzI0o5LTlv1DMA
eQJOTzFmfUZTFkeV/SgZRdVZvbfCMVgtpC3uJ7rM+3drxHBhUeU9zY2Mupbu1czV
IgWH789qTKcauyflbtCAeJ/nGjTTtZgayg7Q6jXVNDHKgYRSGpG1rTCXH5V5upA/
/CvZeA88pHM3r2EUPhde0JEohRJ4E4giuSecU/h/SMhlC3JGTJiZe2qBmYCzmGPu
6V1mvXRyBQMgaHsThhzR36fwniZprHI+qQljWrCcpkmK1rD60vfUgBlk2x6332/Y
VASVj1DdJvIqCNM3tGe3cL52ixOaSdCWU31sPz7REpPYRUP1O712DyWsav9/NBxn
vGcEOIwMv+6ZXbREeVF6vK/j1TDCv73KwTY6cuv3BnmjZDBsC/xOGBLGJF2N3Tke
E6rTTcR1u2l5vtfMfmDTcHpqt7cim/qyc+owcdTIa3hpuyQuXRF6W8IHQaap1I4W
TXZc+v3qY4PWdQPFpundpQHIfupFXJC2/YBcZ7REzcXZQYLldeMApQ4aPOFSqpTD
iP5Anqw3W3XFboQc/aGBwhyQ7xI5CVbpRfr5xTIGEywypXcHcqN5dT9yO14hiRfM
hx+dPQR0Op58OqeQeoDrN8Ez8JM7DSPKPBg+QHUX27KE9t3oAki3UyWNdGN4Yg4H
+h/mUeRuiK5Yr9w0mlga5BOori+qaq2bbFx9QUw4rCXj0ykUuWYipkROY8M83588
j+a3hbeBj3JXWBjtTr7HuMRV95mcWSHr1Z2SWXEAV+GzIQka6D79R1lALdStH+3r
02sHCL4vePtxZchVEkzUvsRv4KC5JGTA1w99o4wlZaWm+dH/8iTn65AGtMLkrK8Y
yvy+XX938R6bbDAjTpmoah3j4sXDKRTl2PXAulPmYOn7cPBuMt+jFlQycUxp0pvg
Y/W/ud3PeebFDJTdIsV4uvKOurOMs/tTqumJkEz5/cFFdKaeM6RpaZUVy7yPyzul
AIS7jCM029QVrd3LN+uS0Xca4RvZ9jBHw5GH8VXTO3LRwIlz20HEgJn/9ucbE7ay
zEwwJPIWtCRpaDE8ZtkhZj04hHkGMfUnXgjNd7RGX0zZCDqSvUsJ44/4Hrs7YvLX
CmE9/wl5iBsj/h2exK1YnJH6W5gJuwZ/6aXVBzkT6qRsHfbqQcnvxMYv1JRdLhBp
0ad0YPX0RVZISZc5+qzDEGIqJYvAXiQQd7L3XKASIT6i5ASplZTa3bYvWyb7XleE
3LTipFPv6roVGg0KmeNPaG1v+ON4SQAWDUa44/mtmzjTc/LpHAfDzFT/+XTjckWA
Ei2D3v7m9fOiUxoRRn2FExb0tHgrv0ZujwrIcgDSKuBBYDtO5SzYvZ/9k5oqsZ0J
KCm6MRk0Mpi/CIzpT8YMWbBOO/dmDwatvyKqMJf7tkat0zoKLvWDyzsrbujYvbxZ
oK8FKMzxdCh8r0k5aJFCEisMNADlqiagDwRjxjd6Ae5bKpNmvxIGbqaKLsr6BUcK
am33NRVm0N5ebe3Y1rRgEaPhmnvbDs/kBwuurx0CrRO1PnidYsXA69WV/f4tIH+O
vmj7S0adrlxcOKZ5CVlf3HL8Rt5V3EnL9gGIs+cuI/p5/mFlqkmGioFOqpJdsuZY
cXUP5RoQNihI88Eel21jVD3TJBOO7ktpHRGHWoKwfqGvsBJsiEzyqQrN+mCxZ8Z0
zwHwuR9KaSMp2nXJirjnNjTbXUrU5HlEprPz4wHCQiUHPj57OsIGaBJiBY1xS8pZ
6Q86J3kreRPk3+ofYcxPg7nWzTxBk42DjYWarCpQ5dBzp5163Id88IE1oxki7vog
rtWzl6SEPBweM75kZjFFckbkkrzhm4KR/15+Q4v019iH68ssIYqKUFgZy8pY3kqQ
jOwwmpUIwXIF38infurQQ+nbAU6kxEXYiZ1mHaVDt2MCAcYDgRWVV+VTp1x8hMyb
LDhpnYrvnkgNKJto33kLKis506bdGm+85d3QktEfiI1XCbten+er3Xgnmsn+8ynV
DkNQv5KyfzdKw2nPHGakQIS+bKVaE0gyKmaokRPcw9w7+5iB5NUMdbCMCSfvNOcJ
hvQ29L6A5P9+8eKAqsRb8uLtgXh1RnRuCOKhOKM/2A0+Cky90pPRn2d3Gu+dVsfq
v0eLE3au3aWJP3ePpyZnMimyfkMT5G+XfW8Rxf44Velje3CVxWIDexCF/Y1Nu62U
Vl4J+rLXU8ZSQGUMSI376CqfQfJvX/kRyc2nPBRICotK6vi7oHAZzmG0jR4oxEZM
ioDpqSJbt4+iO56i8akfWaW3XKL/PV4kf2tR8yKAQ324U1b6IdkLb2dD3YOYaVyY
ecjkixs/5OvU/WxfCPZ2oGmLFpNvIbt4zBpIh8Ab03qihF/pOHZLDBNSqTfycjHe
nc2wwnSyNtA6yq3p3xgFxUPQio2XVCUGUTLM3mI88KhfjUaMyTiA+66H6WI1y5VI
e5I0GaC6d0ULizRfc4JPA7OjpmarxXU9qsTWM8sQy+zZoRf5VtMVCJIaFDTWO21o
6mimBg4dbjbeUbIw0WT57uJy0aP4bSqVA4x42NmzJOsLWaOojhCJjccnOPo/lyOg
PjCeQBAWEiMahVPvmMP/OrERT5g4GbkbyN/qDOH6mvyXlqjpkS1IXuX1rj1iENf5
YkrqC2zrxERzcIVOJz7c7eIPs08NsI3NA8sTdzMNXkvsU1tOHwN6Jhm7jO0EnLnX
fHS/sN+JUvqVarEilstXdsfsr/V9PSXNtuaqaf49U5XWjxLlHlrK9IcgxdLUhike
pOs1tsgsruLUhx+PNp8h6AUvRuvlYTjpUwO0kgBteOmVf4/LYvU5bL2+f8e4TYJY
5JFAxujFeqAcrFgL63x4AiqvL1ViDMSkJmbS3IZJyUNVB5BYFs4Yp/eURaClnCed
ioDV+2fe454cBUkEWUs8nmhgUgjadtNtfDP7i9WmHSNuRWjbq09BlzF0fSljJAO9
MbS6dcuSN48IZbi85iUFc49w8Asb1YYDFjA+rTAdqpHUoWT3wGVWnNE1bO5BhHyx
CiACEXymbh6lWTDSNoIcKp/BPhdBw8uZUzMlO1EnHQcb6DWMEuIdQNfOpKiHCUkm
jYrr///7fhPPFUv/ttl1ohyPlgCNItnKjWFUeof+nx+8eWNz44sN30DHVZJ+fR8X
nAUTz7amV4fe6PPX1YmOtIQY0XdwCes/U7dQV//BxHLLu/vPrD2pk2Zv5xXVeMn3
YMRjIQUW/EvnNoLxdfNdSLax0N4n63+lLh4AVvEQlwy5aRhnbxS9Y56p6XzliQOJ
xL/MmerpCVKmpXdSwFAjV6SbVAohbcmn0UvsmAhc6mnFRmlfD3YmFnMuAsclHY9y
bTlxT6ABLtcomO9EUNwUhA2L3a+FBn7AieZn0wIOITQ75Zi5M5iuBZmrZuWvsRaK
HaXrZ27dNQNJhyeZJX4pq3ste8KJlONhSQLfdmE5/FwOEn439IBRfFq0o21v+can
qHP3lchENE5b8xhLPv6r5UZM0CJ/WlpzezKXkXJgxQNf3NzrBnP3VYrjj1AojcUJ
xK2ttx2ud9jYEXONxqpQJ0KJ/ygCbmN38b2OW4B173HPlxoNHczEiOZMyS8HrdeX
WWfXmrG/xOvp7b4WVKXkAITDy3PnKpoo+z9WUmrd2WtJgVcnBAy/zpogedJjTY+4
YfNkZovdSDiWgHjrCwVmxs5tzeBk06pVnbdJjVq43CDKGvnigZTxjfXZGwgAqEI7
95KM5t53HNIgzarwiXf31XmGLOv9tKESViNynWaGyhdRCMgs7wvbvHoVnqOHHU5m
BDXzvlFxlr9u9z7NVulHih/zRWDcBsGEGKEOuvA1tKaFkHKDMyNJKJJgSk57uGEk
z8m0wfOyVUrYGGYpE+UNVDIzD4CUJCunLpmbQidCZ4DT7w6drkhU1gFH64Rhak0B
o2UPcxKpQ5gZghjs6oIigsiOZ3V1zp1wwFVjvOOZStWvqQboU7I1fMmHwVeoiWhc
NjnFe7WSDLMsquoV0KNAAZSA0aGrpArivzavshbE/VyJ+xaLQWGStFShU2/iu0Lk
eLbsxknubVmP68+i0hcofKH/9KvsO8Iehf3MZBlGrYmyIG1KRg/oPpoZ62kEXmV5
g+5+PgtviwMZ6j+WEzEmS1dh1h+9DCPKPC0pgv9sU1MibOR8T1eWFyNze55Cn0dK
MgJv198dB8Dxc/DDTfgV1nPsWYqwQoTpwjttQJMDzuGlVbJqoaQySUBjHMeTw2zz
U9VRS2bCY4kImbprfx4hDc6TOD5SoR3CKihFqUjkvgltQ6GW0/+2Xgjh1fga3zVn
tzwv0e3mzMbrOzlQwtF8HnEK/vmodUd+5DWArDZB0s3TH0ONt9a7l93985YmQ+Ez
1fel2R9TDNzUtcQEOJqWiahAGibSG28azpqTcd1aFZXzjg6RKLBr2z0TztsjJgjR
vM/R37RtJ/cjmoKDAKNC4KejwB9QJ5NIJwmK/r5fWXdCAQ+m09T9Iw+UUUDhu4ZB
NTsguJQnpfKccwVTCN9COhPp6+dOP7z+f/yjTG+l0Kr/jqNVmqE1pc5mSa1RQsdU
vqDwYoX9DwpbFPEpTcl2uFb186GasrfLWtVf8zjC9QdGofCDfxYodP65Og42vyCx
bZbkINrh4ZL0CPElw1tTfwxJOeALqgahx2miezeEOOalCB2Evq1DfhNG+BQGIGsT
72S/xYgM4umx1qvrliy4vdp91VqQkYYUJEFLwTu3kYg3pr1fdHVdHLFV22v1Z6yA
FcCcyJGSKzXlZcCFvYX92XOasxXa38zc0X3exbXPX8HM14GXG6krYns/utjilo0h
VQMsIPESpxwEnDhjnv4twAvSwExICXCkGy4cwd678agS+6Eiw+JcbM04Ple0xs7I
HUDrsdPJbpaZPqw5S1ZK0GRA9VKw4T0SNY2mHf59XigvlrbY5uiNbl60xEiund1X
7fPBmwZiLaPjY94654vohdiz6JxQqXU9fTl+pZQ/0lcVjAnaLES+6soyHzIXwto/
1PfzQmmrdl4vXqJxuYsUVZ/dOyCrq7g+78X36Jf0xGC5UKdri63dBEJujtU50Mix
FvHwOBi5JHsPZDPJZK9UsVqWNKNYsWrig01pprKeCUOuCJJQ6ugfUYkzHRYxqWoi
+0Y3H4drWAU4QketHPk4V3S34hGYBD3JxJx13NkOExIwjByv62RySoh33U0iFwaM
qL08inpEi38CHhmvsp3iDDBQmyJ4WsfFmQof4pKs/SX6AcHQkfCwwlnz9toZ2oHK
P++HsXE/apFw5llQcBY1aU8UkecHBF8g8FGsvfs8GgbOq/9InOT9ChreZpxCOOZK
grPwZ642x6WTQY8fiootwo/6usdOkJjWKuedJJekg5fjOOfMH5g7+fKrITRJUaAI
E9FY0lf6Z3iS8hUa0gTz5TWclfoMnUAvcQTXCl1iS4i57GHwrTM9n9cqaUU0ut52
cdNlx1/X7rSDvIfslTTfedGlLPhbbpDjUvPLv8tCCiSYxnLECU/vj3OlWPAHc3/y
ZLa8hT5iJZ/KHSmcPB6t1kyzGF6xrRfoxhAn3kYoEaW3gZWKuzAJ3tWD57IWeLOs
sEpl/GfNhnCYvwu57nTdpudGvnU7oxqQHSYmU8XqcuMk3N6s6BrW8VutNpP9n3e9
qvjxVW0/sETXRsQn1eo8yTMhX2OFDCTNT3/2Tg8fGaTv66R/nQX3jEkP0SUkpBnW
KX97tjJUqokbP9Fw+ytRXPc9OlT39k9KuhDYaYAQG1BMxgXK1nobhA6jCzJbE+pq
qcrr550YbIpUueoc6zHptXxj4mmicZ056W1vuFTXOxZnN6xGIqW5CyOIX20fPj/h
y9Q1GSUH7CroJu1Khy9sU9luSf85wEz6DoDzlnjfbz86ZR5xEuRirDdoecTSqQck
gqu1rgPHrcsEMt+BORdMrTEXvQ/6F4o/ygXB3CdMmgFp2GRCA047Xb/KXZAvszzw
EPTPZrPAicpEW6zqZHmwWO1SHgGru+ocA5zvsYHLQMmHHap0mwVn4Aba7qp41QLJ
uPhbW/H0ucucQk9jSvMcTMexHZe2vzF85uBeYAWLhoABBfSnlf733BF7nkjn01+6
sMQJH1jA/R+SSEMPoCM749CwilMtEk3f7mrPCIIA8/NH0qdOCdQKGuTJY/BUu2wX
C3prOA/5Sp+ourINnQt+VYoCxCxr8trQaalm2N+nAgQi/12LPXxniRYYd/0ytwHl
DwSy+fIMLgRtVilkGQ5qk5LjL5hvn2Kz6onq7JFoqDxrzlRqu5tLQwCeemdPz7Hy
CXTgBSPNL+d/Zsw4RnvF5IZZCjdmpF/Y/oZbI7soW+4QSIQTdqQUQxUiSg9q3E9N
SOl3lqB1akU9Oyf/RT1RNPLBlgVQFWC3OwMPrcbfereaEV6mtcmpMfCPTExLltds
VNs1ZrFpz8eMQXhQnuzyjKZnxL0MwqELHXwacduJBlmi14dXGbj7EzmGOHXPHhfh
zPJeGbpvrPA1ethjc9xnqexmYvvt/yCVEIv8MkrzGCDKe1HDIyM3AuYMFecqpnjr
hgf290Ezgjlh8Z6Du3lfYDpkGPm1HR4879PkWdWeqNJaVq+9rAgMqsiU9MBifRH8
IowQhVu4vZpwCd9hrRET3AqWuzdVVyfCVNKZ1HT91JX7r2VvypGkCCCdOqDv4OGl
T9sSndDkNu2EGGGlIgoo4+VB/EfyNYOT0BJXekE1IYZRJLR8GGP9d9KjdTtZ4zBD
STGU87QopgWuKZ2rQAhNz41Ef+yoJDDgOEzqebe0G/3/9xelZvV3uAHP8mpf2B6e
XbfLTIqBqgvB2U0dX41nFy/yB9WZhoJC/V7Bh88XVIseqZL3+BEzNZGKEVmqAePC
BDS8tcYLMBNHTf++v1TaHpe8UA9ker1vpypj55dhBmX4MGZVj4HzkZbKCTNIjR/0
tUeKo3ia2/HCwW/J7Eus9ei87/LGnimRJIr+2NA/8Lg3+uT/xEpykng6PHxwSBV0
Ilv9Ggjr7hzre+AYFKJ93XYCdaAMz3ozUYZzTPSFVj2fWpiFA86jPurmTPiy1ALb
KvYxiLt0ayaRXkQtSoKLR3HQv/XOKOXwv/2h8HOWHXhv59gwuO2VKqGacS603U0b
Pli8i2uyX0ZIAy5lhppT//qNPFADuUvjyQpsxPC/2avnfp9oDPpdL1olKd4Ou9Yv
hgir1ITMaSajRhbHGaKgEfvBw2T9ZdLfRyUW0lU45wJL5E4q8Yz0ycZ68Yf4psGm
IRG8aHxyZxFCuSL17PNE7fRlTrpmT1b6hmPOtGPgoGEuYwqqTKD/FI3qOR/jxTuN
9C4mRHHKclsN65Cguv/1lpG57dO5XnsE35KwH0jk917ukvthrc8k4UsAldvO+CHa
qF/z41v1R/5b7WFYLa7QJfdQeTxUFGUpjJozKz7LeFMBjKgyQoXj/M7QhAzOjfuI
oqL/i8zdwNUWo/wLgrIbGBEXghDCC+mTWCu2wu07G1bqApWyxPWzKm/1jYK9hznE
vEtgABHiG2IRNRphrJemzqppJi5YcRb8LrBF2AvK3oe2q9bSZNWdlqUehgHXW8Iw
iQFqnABe2hImXRZAwuFHeBe7pIW7tBW/WTMxjHOIG5MIRtiOx2B3Fl2tI6Lig7x/
pYv0vQq4+PA684/axl+jMHMA9dpBLPYer0qivsFBlkpa0jJnuu0VQb5zFMPn/SUm
L8awhxH4OZhixyMzIEoe7dC1+T2zLjej4c1H2wzdLYMLhXnWd4o/t0F0LCJz2jXw
Lhi/fA3ct1svTg2cOCdGNgRJjV71bLH67mrVU/I0DwgvkUJagi1ODljhGExwCul+
7FlKPzKuigP/uMGvyzsDY1Au6q9avUoRNXfbMuMiWl4gWO33y3NVnWg4pyCVbbWS
xIE5kwIep0WtmYrSDfOylI6q1affiTWIpej/aRtUYn8PIqrSZCetKgBndNPOJcV/
bbSlduaCz7ZgkBOTZO9q1Nz5W/3KOcGJ1Z2AnCOkIxYEWwjJEaGpuvhgA7s7gMB9
csr86zuetPzHBTDxPnxSKXtg8FTf5T2bWza/puSAydsHnpr40ecw5mwwnTP6XAaE
4Wu/fo6cGThHieFKCrMLQYxcpmGct8GQ0UWKmU1gSXC7XDuo1x3UmBU75/PuLxSo
XWWRK3wGNA2u6bI3mwfutcULGnAuA7/6mK/N6gobKTdCA4XbSUMIeMt1rqQG2Hmk
Un6CC5s7BXorJaZIWf4wLIs1ADDBnNKhz2BtzvFF/TB7eZLfV7y6JFHcK+XtX+yY
HbJTuEk/31k2dQf8yufbAIgFv8DuvEKZ5dnMfqANfCq8rIMc1ibOkDxQsVLAeGQM
Ou9Di1PQMg7g4xpZ6UJ8l44G0s0simKNhVPPe9QXEdzUl5eI4WW3P0/JPFPqND7w
7xUzDm85AleVbndGvruVc1rCchfwmKiUN0XFql0mA2aIJHxBJDLRGc1NYOgcueRZ
Xag1/29wMreY60A2KmTdfk+U6nnt9D3M1zfPFMbefFKR+7dqLxu4+sKf+Xw9/+15
zBQEK1knfPxbFc3NDaa7dq/WFg7cdmGeIMfj6Sr3lqzK1IS2rz2+vvEIl5My4EvJ
MOaCKwM4XY43XxPHtf+wKclNSPQz4F3duOuJnhEJyfgRaUKzUJcrZTFhPAZ58AFa
3gxBtqHw16g15Z5fEorkerQflAGxEVgI0bNJWCbDrsoI+G3/zayZGbGZTLQ4kqVX
JlrX/c9K5UamgWbUc5Pp6wKVKoQllNpsO2UFCw1xQzULKg69vt8o6zaucL63vIsL
V41OAYkmjahvIjsBwlxUKcfCSF+PwqfL3mom9NP4IcTwk5ICOrXpZd0wm5duNNm0
MYNlJ4wBdFCLrt0ZBpjXLbqm2xzEWod88hvD4lCE15yTNVEcm938AyRIKfbmHjC/
zZ/RXzZrR7B/EoLN+JJPp7/ryZI6HiAf7nzsIL1thddI+m4P4Fly9huClpzIhQNM
2Z3Ig6ZVbEMu/yyIXh4T+eWtF1wjzNKoySewcNK+4gXgOa7IcHL/1fMv/6mjA5bA
/uvL7Hwc7D/G1gPqKB8blaavrUSMlCHIpupStuVo9nsEdpAhgeXTt6EivpvXV4OJ
OkkAsN2QtMxLTAVdL58G4yTjHshqDAN/GgPX+NbVX9T7MZD+VNXRHIzI7oAXxCLS
4eFepBJSpkIJplf0sgndTIkTQNhjI0alLdeeWJQTOHqaeiU98hZLRgJERNozpA2T
TWHBqaIS+9eGX4sCiPSYjwU3U6JWg/X9MMwtyCpaa5MbyLz9qsB52z8z4JqwsWZX
7yY/neqb08n5WvDRBihDkzq4mIGyptY9nJpcHkwaKFcZnzmNx1uLdAucnqn+a5TE
HMlFmKGwMB1XsTQIsk0BUirfdTrdpnIuk7h386qlS+KrI2W9qVFovizVIwe17QFk
C2BKLVSfo7GcU4R3DhTc/SWwSLNqvZWHEsA79H1pT+E7UB0qx7E7fbmzyQop9GrO
kPMJNs7Pyyjl0v5U30y8r6Dnot7Q+mteuyFoVzJtX6UowZ1jXVF84I3vyrX2Z0Gf
21QaqF9dG9U24U5ptm4vQXTXyIUZwyMcTEx7jee0LqEZc9GR2AOTQcOQKNSwC3X0
gG/KR0nt5GvxGE5Ickgw0Ny88ugP9bAJjM/nlUNJqaWODvse2kAJ7Q5ZkPRRe0xm
tBfEapmXRQOeD+fTtPWE+QuUB4Gc4TKO7tMXlTkptWJi1HPlbX6lbpOSDMraShH0
V48z/C5NeEsGDpJ4a8JkmY3JcXNFQ2NNWDVu1hGeg1HwW73GPcvPGEAxiz9gNXdK
F/YXKCpMXgaVWjOLyH8GZ2RYH0AQxWvjSkRjZn5ZwLFix8yB8dWmoJIMAnFVpHrK
vt7B92Zz23mUtgVhrPlSxCNRNul7CAumRAT55PLQl//Dr6bJFDwVx+p+Dpc3nW8a
MF4eBzRVBK3/7L+9nmLRoQ5oO3he5NxHlPIC/NVGCxqiX208eYMCHDCDBgBn3wtd
VSEhx/FMvlEvywK6tQgA93qbENXZhagSBg+MxkVPjtu5STFF6O/UU5CptGSsfbsi
RmaUpU+di0sNI5gUNkStcW/Mnce6FuSuIDs9fL39bLjWjcv/+2Idtux9gpCcVOVo
nzvs+1uZJ/22Z4uscgYkf+mMvddmyCYwLLVvpk4CkCdBHfQ2G5rai0qdCir11HN1
PWmooZRdWoIhEOhluufArNaP17LZ7potYd5qTZE22InN30DKloSc2gms3pRibl6j
nUHmYCLBtlDtL++qJObCLnTozRjN3nU4dlfPkHLzYBzdLfvceRYAFbm6oozHLjdL
5dyW0OmdA47zKgNdek1uc7/CSFn64lDuRibtvCk71ISzdqv2IBUe86dXOI6rASpK
YBPcwsrlfIJkbcM9XbdkxhRzinNmni2HNP4OhPrE8qGzKWJSTgzhaqxBR+qotyQD
/d4yMOz+TDLMPfD7FhxIpbp36qJRkcgvyztIRkGjt7SSRPyJck9ppOqueyg5iuE3
cIBmsnQ19lSafMCphDzkDxBdrKf3rqh4AFZ4B8N6xyzPIUzBuQb8ubly0cfi1lko
BwcqkZK5MgAi5EQ8XP/PPp/9m06fuOtmfOyRrBrhykFMwduEEIlNZsPU8Wd/1RAv
dywe76+dNaUHfZd4wlp2sVYV3jQnuCLLQ43G4RV08J5v6yP0NBhTdQp7OWL0UOcn
BPasL204T2tzbH8rY4ydQyP6V4mHKNVsOI1tjCJBBqM96ZURMx8POBy893xSYZ5C
aqCpMT+8hwdiqQ/vlx/XtLLBqnXUgP7BMAPw8BA6O34kqS1WdOBPrx9Xdp0fuhxa
ksF0Cm7f+l3f/XIFJSh3mVtaFcb9Pkb9sn5asPnCglnfEiPsR7c7wP63xe5p/ACq
wkkv9Qkmi3nrllkanGkbN2GjkQQ1oIdbDpfHOjGNkn2hiHCr//uXNQkpS2DjFcbM
9pDuPrjBEQlrvWxk+8BZUgntbaNtC1itOA+AxK++zCzJaaBaQhHhEhRMfH0PBZvt
GZA5QXcaKEgAZJjnVbqLXUIRfnrry3KntCbijF862AN5/49RBbXNnSRBZ4isQQyR
+E62fARTjLBPISN3elBkmWXNoCmINx/+HmCmzUJToZXYgeySmP/WVgbKx8sEQWF9
zDwYjFK4DSIe8QrUya4UcKAlaw5XcBO/mJCvDuOniYMdiNbr3FvV++3Vz9jy3ZZV
4TxGihqs0fn2AIHXP45rmm5Sq82ywAfdM3jQyEa8N0AWpRaLoMlnR4ap95q5fO7R
YK2zn/btDhflazQ6QhPly8Y+TZHeUm/KkHDBFk2qRS56nCRUCXiiAKp6BUQQ4RJn
+f5aJVFJyPINUt8pevH0/AHOkBPfncRsvTXCrjLDWu7TGaCMVH4mjXfKQrS5MO6W
i11VaZMgMrrYFuxeMV/LHFUbAGrKuavLM3M1AJEOMYwZWkkAb9n2f/dZ+kzmH12d
egeY3+ET4XflJHRPG5bwX4obTN9ddf7C+koDedAVSlUpNEmuMqYjEFRjiA/v4Koh
+HSBocGGcI2q7YARCQZ6POyBLjc+Pc6HnuDEf/v9Uc+F/RelR8sBXpZUS682t8Hp
ZbFQf2JKHNPi5P9CEZRjnvT39EM/gveqswRKBcD6vUj2qprvYQA9EokwdFYLb3re
yIWuQQ2wmQqt7Uq7AVJf73gdRkNWIc8U/ebw6EDKMQeZ6u9rDAKoDb9YR7OZjiAf
HstgE4WXLwcrm5teCmxvGx3N8Tcl7MZmp94JjNgdHsAIACi1iJiTKsnevpSt9I3M
NnR2QLs2AGJsMYg+8YXe/6rIBXIRK+oWkNXx2x81blOGhkk0XfCVivEXE+YAQkTd
3iNqcq5Ud9uDsudGwe1z7O0EoXiwD7ThanRlgnZLeodNF4O/E+dluZU+8+wj0b2u
ci0ILHT8YKzNW3PrQuZbFDJ6nE6qn4UMO+Icqr5pxhiBad4zW22e4TTWBcW8xljx
GQeTiXMSXAVIXyZxQOG6IuF4ATj3AemkLr0YoOqo8KR9gYbuhn7ENEKDD5QtxchV
ETwIgA3yXD3lEXKAx5HsXdWTVZqVSnazQyzUWBFxb/4wE9dBqwUBd/hAm5XAXmKM
C7ME+ZHcMg5/Mlw+s8KBW4or8N0RdEn8s50mTdv5/kEt+v3cypykwJP094mdOxKP
8nYaY3i/6B7lO3p3usxGzXEiV57LfHwIMBBTUpO4bvTcsrZ0aG+fzUVuzdvvQFX7
A/xW3izXCqXOfKAVz9G9M5nb6wHTQlhk6tGNNd4tQu24hGXLC85D/rpk18R2bCll
aHJRbWul96mDYvfCgYMVwV0deM8hAo7QRtmePynvAd1Wj1CZhs/EbRBwqNrU79DP
SHDFwhPl6ouOVV8zjCyfBK2OMddyjgEeGcMYDMbWptqQzK+kIFBwcLTQmwnzfpgK
ysk6t+F9GnejeE7Qtr8pUy8bV41DjMDwYlhgedAOoVrLwBQ5UCZ1SZ6HUr/3hVIa
H6XRsHhkwlryAJ7nd/Sa7pyyvUHJbz5MAUQMF7Uuz0yDCy2rCtRaEpp/P+ePbYwR
b19UsAhz/1JGp/Qgzl1YMbWdXdqAmtVUWpa/dA4DEuyVdT79byse1V0qLiKaBH02
vX7kQcEROoSULhRFF15WJ+/UWzNoXm4uxwkP/EOxMOQV6xLTY2aBOgX02/9SPVnL
H1/LsLi2K3RQmxLdFzOexZ5d+WBZBE1ghLrKMJ2BfgB6EuFJ1rzInn4T/IbJGCBy
BsPXYBBG9os7gBQK4+MukkEN+6hmebnJjckJGBlbxQfAoBaF/H8KhJO9Jb+wB9MP
vhzllXwhl/nNtStiupXwYVN36aVitsrFwj2/eLw+PiPZ/BD4V9EbTDq5lJzL8r8a
YPSsXxJirkK9PyLOZwOdbrmallvTKUqAZ+fCxlPO7xDIUcfzFpnU05nzq7/UARCt
APLrHymmLQj5fGO7F5Zthj+phKtxLVlu0obqA4hV7wJRrwMeYruEspgacKg9LnC8
/gDFxwK2CCrDLXlo+FHZGE9a4OktMVBpy+FOw6wLuYqa1R7edWrpdIp4WdyMIVxl
d/Hp/yaRix9cjTlahqgCSb1KIoC8rFOloufp8+KZVxx08/ko4nwPU6aVn5L/UpCr
XojQftmGB05Y5FXuI3bQ/+wVSv9aDZs2F1v4+oxChLdkZFxqwSfhmPBHm4gegSBi
l941fifz6qBwgCdW5Z/pijeAxrmP+ZhB1k7yMCxCBUPwI+Vgo2BBzUZK25YzeRGP
WPDxpYB3PSPwzLPquJD2xM4I57FBJaB+KmzMa1ZSeoRAnEzjieoaKw9HmZvHQPc7
bpPuFRI7BgT9FwheymWgfcmkC85ewQuZelANk3thCoMREhtu+iRltOQLxfpIJh9c
7NJ6tlMJOI3Q5t7UpWIi3oTEPN4BU3PyC36TPn7uuABs6nUJ849gj6ruzIFjltCI
m+TD9EAGda1HL+c8Mu8UuXkiFfUpEqLQNOenOKGfy/43gbQkL0EK0+1Lcpkf2gfu
vc4Wf/GXiSPA2Qbl0hMtAMYwF45T6Uhf6xR2/QIvJb6sbZLV7o8M1pIj1dfQzip6
/ge5GGll8WIDhcByXyYZUzTf4bMK/0zECmHgkl53/50aVs2k3r8jmWpp2kAXo4Eb
gyYKX/6lfpFzycsXyx8u0wFEGjtdw/mAPpKt5VlqStZ3z5oPVkSzkDpYr01F6B2O
OAzJNAmlCLyFIGFEQQWQeXg6yCBigZOMyFtpeZ+V0jGjLq6MyuEN44UOXoG2YOla
Gmsm1y8QuNSD7yrf9p36NPFnh/5aum6zpTTn20k1gXiSxTB5n9Il8mcadB0VVzLt
PxPBFkMPErxqgkVMhDxFEUE3s+ROSPBBi9TmfFGPNaV74fXRZJMxsqXuT8AiHm7o
ggnMlS7DS/ZBesCUwX5A9aTcMn8zDJj5GK0DssSVQnc=
`pragma protect end_protected


`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
aNsZzBu/0MF11ejgqpKfs/+Dp9A1tpsKW+irHvp2xkGaHkJKTAyGN/DyDKWk0TxJ
w4vIIBXw2lgGBWt+/l6P4gg7n1xwVWQ58ZFGUbbu4kT6zNMywsxIa2G/aTsAgxfJ
0g6N/KrCg1gzrG3gShNWPAfGiuQyRAaYeAs/cvTLtnU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 379040    )
4Rqv383pbcq6jG7nVdDAVcUscsUF20I8/TJhYzyCVBNImfJP56iWuAdPBtSUin5x
+HuOK1EVw7Qbo/3V39RNZIB9uuvNS3foVVOAc2EbL7WNvvhoIL/blV64dQ27s5Ud
L+7Ijm59+CUsEsvEydSkgA==
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ESyHAazIJrtnRbyGkD6YtdnaMsXl/jUgG7KVjbvXIJUdquWpKfHPIqFtNnP/j54x
eyiLQrFIcn9isRoT4dUdMBuakTK5ZVr7NWsRbGAURNGP6O85tnN0v/YrWhZY/Wu3
HIBPvBhJ3+ZvUQJ7qZlC5TAwvFGUfZ0VS5ADcLdgiRQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 556360    )
KoTJmk7GkpCsHA+BpAGQcgm2jK3PCRgqJvxrTtzQJNpX6GP0yvIUDa0A07NZeZME
UtMZfXYAFy0QK7Dbr6nonfBcXPgMEO0wBXvuLVcxj9dCyTCg/EyJRQMiy/vwRCnZ
Od/GBIECr17qgFv8tiqHV1kgIXwoVsDgWJnLIpexJ8WtNixg2oM6bHsbJ9CUPj+L
SVv2Olb8Vc3f5RPgERNrtqpoTXFCqoH1xHTJfwhc0ZFj8MVW7F6wWpuuXOkaWdHm
TgLWTfhJVmKHjFEuutauvZCemps/sEorTY8vD35MToU0Do08eG2IuLLcMYeB+RRj
CRgRNJJQF72wB9S/tZlZGuf8baqZy4ozQZKCcKR7tLvIW36fpEcwHa9hdx4E+Bqu
Yjyq745LZTJWMNsL7TJGkO/AQf92BfTfEQhSD/l0HAlbfI9wZh4sc9dZjcXZWPv6
2sQKWjWhegK5IRipDZPaqSRMqqsatlpeuOOa3s9lkyTTJCTl6ou3YrVBK3mWI5Lq
sqj3FMHog4vO57Bsrjt8PARtgqVhJTdWQ0vtz81SW2+6kHxwK1d4U3P8p5cOjSXJ
GWz4tzwyOkGNvo+eVzEVgeQnGELiExBHx+vkjQLYTAuI9hE5BM7RgaxO1LGlgBZQ
GtQVUmwTKdY+nrUVIKPXItPtNHLPqf9kidiNV9vi2GNOWOLD6HxvdpM8amnWA7ND
mto4s2Ju95Ao3v9h+SjQ2WfB7jNy/j5J5k5hIv6/EaaPgj2ms7YiN2s9ioc7/935
RZaHooTsNgfbs69V22V31/SkcSOyu1kyc2dyvAIonudZD2LZzQMbJEXviNGR9rfv
y/n8t60QlQejtD0xz6fya24eFS6MTWEcOSmtig57vdtLD4rmGwDT1i+JPdLHysT+
s9OWNnW0D0csuUALpgEbKbwOHbXFxTauILHeXkMCyTzSTgZLcvGgbO4/TSyXlNo4
CB/gsT4+glTPvcG7VXZkXUvgYtK+354+JVWQSw+2X/lHm0h8bEo0nOg3wyaWLvGe
bkBU4GlZ9A4J6Whfk/XAEyEg3SKecV2124hPIbQfHee/TmhzEz6L9CWgEtVSerkd
ItLesCQq8OnzIVL9Whxzzr0oynw3V8wmbUrEZTuxYnmj0hPyfODBucPkvU+OcF+q
ADRe4p1zM2Y2sSSwUBlcQv9ngBmMpkTLNWuFMZw7gM3qhsbkyC7kwjB4nMZJWQuQ
7y0C/2lrPjNi3dINsoDyOzEz/IHnkT4Plfg7V1xx80X0zxEOwNxIN/Z9YsLT9sco
1nqLhFeE5a8ZZkhmwUAoUC28n+rOt+CQeK/cMUGnellDWqtznqlhn1A3bbxRX/MZ
LQJfBO4J1b8u1pE2sjQpZgiorrU5spTrbtn9NYZaHiZ0+CxUZn6BBRCMQpw3o4D1
QDm75jLUL44T+ITZEK5gBKNL86iABWNv/0QpBypUa3kIWnFVeWachORSSApHUJua
F9ivn3uHDnFMq7gQQXQNtw4NkF4LSqsU14WcLdiSxHiNd3OmOkgprzAvi/0fypdE
CizN03UouXARI8aZkksP/mP0+lKCZCUbUnOHOh35flsAhC2y88iyhOTwKaXExgTW
FBmaS/ALKI1K5OrLckvvSnFHu6I63pMEe1gTOM5v5EX8jC8BqmfNJpyojg51le+p
EeGUa0JAf5Mx/D2JgH17kc7awguyh3d7IZjJp3doySk5bNZ/huvFlm18dR5Ct8Ly
us0Wr6egwKHhnEAn6MO1oxzm/pR/N1YNNLj4Cph4DRMcBHLBeN2S8xQuFy4cB+2G
q3xRA9aKZbr0gLfpMiLnZt6+jrKj2jh8r/o/sI02v5lfbyHPK/QgiLPPPg+T/3cj
AYm/4tB/U3VTGmHXOqF+OhoqyO8VUuRl2dYYQXE9cu9ZN2bUY1tqje52n9f6Gkqt
hd9MkDwAHr8XWiEkXnS83WYzB6xQxQeo6+vnKR5kNZexdto9PQnS3FFIUAIXhOvn
UeQy/iARku0q32moC0kMUJ2+n1gD/GUOIfWutioF63OJ4/gUeqRGnOSPCqSlt6fY
Tp/ShNpyKXBhEZOZwGV/1Bo6Bd5RCtSJ+wuGbAW9N3QcYiT4PXY6M/nFdI10kMo7
uIcJsv8XwcQH8z6ID2xThNPas+ZGhWzuJQIKZXcPTNEVWgBkxD2tuv5bL192M7b9
wNWQMGJnFRYIOOlokkITV4vMd7T+aOspF78ZT0+wmH18mgDK6DStB4lviWOaJpwz
EuC4ULq2+6oKQCtrKCbQDK6Tq5//prOfP0YdbKGC/U0kpNivaF8dgvGWnIdKBc8X
BI2wvXiNMoicN86o/sPHo27MZSL96LisFKEAZHdmB0xQCkvMcetavDsY4yKqZ4Qo
dSm3QShPOB2p/W2Snjabq6bfnbD4G6EgCci3qz1WFmo0G9FK06r8yFYxeaHoqm8C
RRCrVuX3wfuftMfsiN2JW91DkAdHJij30DACaxlbl4sK3PGSw92KTYuFNBgHjTfv
XvutkzBJzYFZVomdMAiODTmlgWQTAXlSwoX+Yh4PKzEfu4ngVGqHBiRZ1Bk3H/B7
rsvcuMiCkY64NoZRr/u90FbOdoqczElixNyhT8tzXTioKbcGisgHGn9OyIcgy2bD
iK4X/ViZj19swGbyLqcmrhLKjQs49zr6DCOWlWwYvCdaMT+1E9z2J77n4euWpNos
zMTsYmJXOnhGMdK9mUlpavUtV3cJ8Yn/9y4pVHL2UniM4aHdSqe30lhJQg0vQdbB
Ngjp4nuiSt/IqfHe0JHRtho7lakF76G7+P50FE3jm5qZH/TmijkaU5cN+ciNoTDN
MFCFasZMTZfQhlamRdIaPsOVSgIFGorzOPEFR01Y40q9QowkWRSIeRAeeR5zLJQF
K7uovCormDzCnx5RsDJBeFrMGcFOObW/82FDPc9/dSVie3sOtMYfEoKV0NMiFq7v
yY9YlM4UY0pslvy0frmNHPiORPLFsxw41ZzkgEh3BtJXYLsHNHEGTOFVKBNqE09J
T9IcJ9n1WD5jvwZpqjiq4vrGh6VRJvwTilUEf6eJ57XvXwW19YKdJsqXINYFOy9y
kUgySJgg5UP0hQjM3VIfWr1aglWUwI9WiN7nJQLU93LENtVD6O6ki8fp6m+BlOgl
J+k4rmnLGMT5WE8KiXS9pA9pS0p2Zal/Xr/JuYvM4x1VpT3UJdk+wn342ealHRhX
oRX6OoIPhpZKxB+lrDBsYUbUEHkfpkVN1PJURByOJjaMUtUKjl37zpt1ZiOfj+Ap
6BgEnkQXanYeSgh+vSUkNpzbnWKVVEJSrR+VJVrzemBWb9jMIsOaExw91m0yEQXX
PDQbR1VxeCenUCLSJkzsBNXsTpBEEAo+OT74khSHnyJ1njr4mNuioBDpJZXKJCm7
aLvZzYNYHs5D9+Db+W1XecwbyjLae0no4qWUVJeYks+1XxlM3ND5Klo9BntpljD8
lFdxgDCKhkQD8TY0k/ZCY6d8ymWjiYmc4HiwLyLvcvEse8VO1OV33l8NrUtyvuFS
HMIgZ8sE0kfso8D2HdqY1E5Xj+cKm7seklrMOkcoeeCDBqeP4b15RoAQOAdvcOsM
DPWvTxKtYtabhngFCtNArhFWuwftPF9y6dDCrk2KLiXP6GgXlf6bvZpftbdMVzDO
M+qQqYYTH/KCTU3A0tqJUWkizBVhPcyAdwJ8t1pk/eK7CfNlp+DvfmdM91xeXjGz
Gh3G3y0QN5u5pM1uy3qMndXfaVZR+PZkMmNAoy5qq5VnTmpv8M9995SahGtbWrZ7
bnDTxnndbnrY8hUCS71aBqD666IrYJQJ0G5tKOiksIPb3nQUpDaCVsid/1KOucGx
77aNf2I9zPl5hFmCgj2EQHbaM1RypKQhtncoglRj3Am++juUZvlIxojGRCVbV0bD
8LEfKDuXLln929cb37NXl4thMK41q1PsVy0lRylYiU21OMIMyBic8aa/QxX7Op+h
s5coc0ljgg1Zoa7JqzI1YjcDNsQKh4SSE//2TScS4brOUfCowX3pK3Uml0DldNNt
6kLaXGnE0OHYgutjEEt2+qjh7wKFTtYkJ9Cj7DVJiSR9xeSR1icTi1Elk2qe0q4H
BM7hRSAdKa0gJtNRwQC4IqXNjJz8ZokGe9uL7AL0mKh2DM8pWxwwKRi5GgMNCiib
nB6gUhgSA1w51RjRfe8TcdI+LvPaXcQnr2+styVPPpc4SFDp+Z+tviJTHlKNnKNc
UtMd8ornasAD5rQMgtT6PD45yImvq5YXHVRdwO3E/ESF7vtzaK/izKZPI2bLlvy4
+oGOyFi2O1Gjl2i54cqb5+Tnjn4EjRFaiBfPuFfCwblP8IqU34mXd2xBODVObpvO
5yjnNr5emRUtfYrZxirSSjy5MW4hITWpqwiWvTkueJ+/2N/jhYU9ZFhsYoqYuykf
X3HA3tEdb/UGArGzitgP64fkISaitAnyWeM+vrPWOh0a7UYazr/FI5RUQws6eXN6
QuLCNLYhzwOjF4W6M0JwyKQWQ7ODH3VSUVFbm+VV1yhug3bB840ioQtIcIuOjRKs
DZ1kpyAZo6S+1OeZYU9NlWer7yi0xX9eZMJvGc8XxNVruT+MCOnWyYl1KGycYbmg
F8cQpWJZ9iaGXVWfnVFaEP6vy3YbSR9H8ihTWfu1zUG5gAbuXEQ0cQgOGw39T5bU
4xqbppcqbtBFYBa/tbAUD7ABH0sNrRfFcaxFum9HcjeJXe7/HOnlQOyYHY2Is2gF
RwOxkqqyYoruq7lI9uTaOgdP6AzUs84b9mXY+6Ui/9NeyaPa5YoUZ0Yh0x/TXQV6
kGXiLC/UASEptJjeMT3eEU/cDC5LSMkeS1nNgyHURjoTsfTRsr/mJ1VQzyXTsi52
M7i+k53Bk0XgwViOuMVi+/oMxh16g1n5pODsOtlmGEhdYeupBDZna6dG2UU8A8US
S6ceZte3/lpAyrUIG5fRLRdiUCvLKHKyf/bK7DneZpPHu+SACgZudfXz5eKxht5N
P1smFIV6Xkm3nqC37zP3QzbvDUhsr0/gMpNTHqlxqAI6crgpcJNuLmpXF0XT1sA+
5nHErb13JF43XY471S8Id+/EGMymjPA6CveO2efTZ+uoi7nZ2BZ24mXf4op1CddM
EnARS04mi+kKtV7q6QnUW5uCdEci5CPEfWuCG9dFnh31er6wonOepiUDOfaoMtCW
LfnRnKdCO86mNGKWu3x8WsfX2gjJRkme7KJjmnyvg9D8aktqv+rvCQwatHdzaoI1
7B+F5EbA1hHrCJOi8qjgq6Alc2ffz16XNeHus08X0WG+NI6lO3SPDupAEPQaITPl
s2uQ7CbMdGqjgQ2KqGyfnbvWnXDhe4TVigRFnOfTuOWuYp+0lCRb9CZtNXDx6AN0
Jy6myreMH5v5uAV8o9lSwIaLp42/AMrNyXBdIiM4UMAcR0vuwTIgu9std+b3FDv3
11bk0JlH6zwaZqr3jELSYb1m0zjyp/8SYfFokvsT1c+Ml9Vkx6xawQMZdT0pcTgr
Nu/bPkHSRjOMGtKrOd4kbI+qinVMgFL8HtR3FFyqj4t25zl21xZW7l+tZv3oMSvv
w+udKRfyFT6l01a8gpOFXZdR0sJIepFRziGToblJgb6Zt0Dwuz5oA9gvH10gWgvH
FHHM71EWYlrc+jDD0Epq6nN/Ao1MzgFwh0wZO4xFjIr+ArU5rNkQBeFwyT/IC4gG
NwZubZwF+jbfN7dccVnqYT5jGT9seMCIOPmf8iodm5oIBr8sh8pOOPWtsloF+3RJ
4zczpe12kFc2X7LfQIB3jkOAEgcdApb81HdLCIFt+QxAXPdgCZ1WzXxbqIXstBfE
Lw0NRZSgqZkSzUxkKStbopI0Wgiw38bfbcRJJ8GnVyYOAZsHtvcCO1K92QucpfEL
tJC/ulWOQ+ZxhPiG4n4dkMMrXJ1W7lic+5lYCY/mBBAMTC5ZgjP77N1Gj6rXFjls
DOTb0rU/DD3EMngTzwchcakki/Cdb/FiE9RW+x5ktlfrXyzntn7Yryad3QorHC/P
E1vXHjvfEl8Cv8RjKyV2K6Xa8YjDfAzpqUiKEyqgad5DWR7CsQgyT+ymWZXQBR1a
4GlbRNEAfkJJE7lkyWSCxO1+J9r/YQZtJFvVy+syjy91k/eoNJLjhlTQBbdNrNG+
ev5yu9vdaR4zhx/wCXpj3Dtu0U2s7b9q6As2k0VZZ0+IK0Rgahc057VkmqPXbdj0
PVlgiK/N7iQq1tjLvkpraT9aZ2eqX594P5VyipDeYBHgkTClFGdeqCcGxaf9PT4N
g7nDW1clE7IGM3b+IGm/ZbNsSEC6vPlBY9t0tlDAgHTGKYU4rEdR3t+wHEku+40X
cl9vHuqTJYC11/iQlHUqiW7a/+4utIiM7crKkNHGL/7qs2qgD0DfHGJ+OFk1Kj09
LJ241VmkQ3kqp3mZI2Wi2Vg/7+PeglJ1ee4QQ/ThqMvT8wooLdllYjDuXCoGxnBO
BeHEUC/s/lgMwUkEZJqf4qGCl23iXT8dY6lQjWXRRtXYUk3rHxObPDY7QZKiIB8Z
2juzK/kBKzp1RAI+yStdA4p/Zmy/wYVpN0YT1poeBJBq+6aQA9Vhbm8/9wSPvpb4
fH7SyEG9flz3UenJFOmpBb38ZeUn+ML1WXfabk6nTEs+qCIDFj3wBbsV3If9K5+p
0yR1bi1hMwVQRBkyrDvvxDusbL3IrC+K/QzmsbzU1+ntStPX3bQRtMC7q3p25xBk
ScV6UGoYJk8qStK5lapDE3a/69my9iPOseVUmDKEFSBc6GTxsImWLw9Kg5cFf7nJ
aJG4BmYmoRl4Q/bsSACdbq3lfNOQT00dEqh13upeGy1HcI+AVmZ1MW2mfcDHeHI+
InrJA4EDuKQhicfmr3wVRLiYNsB+lAS/DtXmm8WfHLFwkWeyguTd5vCm7x8Or58A
mtK+I/aqVN10NOV6oeU07essW026+kWXuyzfN0KSFVECPmLX66tUAkB8nM+8NOI2
IokW7oqt41PuqnxIyg8J7iO5u92ZioABi2hqoos+ugUw/TiRQbBjtPrkKZFrB0ls
7pEMTYtNBQSyuEIa7mVFxi/Dhc4Fi9dZAl6Iim0qy25i6H+C2Lp51xH16KOycHL4
AuqIP/NneZXRDaK/qSIJ9hd9Ep+Gb7aIPEdA42Fc2WozQCecNyzkDaFUfB6OlyFz
nagQIdSy+rJcxcVMXfk+lP6CceZSEu/AszdMreVMX4AbxPG5k9WMVObwwGliy4yI
vbviDfu2SX3toO7tA5ZbL/rnPlrFRDZeBOripElp+WuyUJoJzmZYPvYDN4uKOZEE
4SjWhUCUq70NFXQK9Fnk+ZGMkyWMLwXIsHbCBOgSPUouso4tm1x/ziYnlBJyhpEV
6kxqx3Ea1OWgKv6qM1Mr8UPGMdhIvDcuSL3MLxG9gairCyfEVCPmgE1dxFvHfB7w
kCnpB1v/W79MZYfjkXfCHnXeP8ahJNVFKv5Qn/E6U+j/QTa2ccQ/FMr1580tFbDV
9vXxZ9jyq3tGngvO3xlbwg5eV4tGF9NY7DLMO/ZrPQg54VYDp2+spIk+F5w1j0eu
vGbrOVVBHBvp6xlamaiWs7dyaLFRE3thYi7ESql1Prtpz1AOH5O2+H0MdlyPYseu
4NR23GJmu5W/R7UkzRhR9zzpKscRfi8JvecAkpeahag0tP/oQJU8t6y1R9tiqwnG
yvPvPewiPYUB+j8YZwkIKxtI039I2oiUCV4yJkCJCFumNld3evcasov6e0eb3Zwl
1cS5fFLxwefC3A4IP84FrK5f77cY/QvKUCNvkHJJrfYRrJltT7YkI6DJvh9es7dr
XoHYebxVFUcgQhQ4O3BZxAIK9acwhtlJwqOBNaAPD/g+ZHs6T1P0BAilTRA+F2kD
OLqaDMnXGk/ctiP0VY49nPaXOcPYq2Yi2ZnQZfhw62glU8NUBYLwsvGXVjXy4ta8
YIENhjLGTO2q8TYAPDPI8D01kYeF2a1d8J+MqifcHrNNN1lnjw/s41aRPuXT3OFS
Dkopk2ulE1M6bkXh0zuABTjyYRIrvHqBoIEGEAHkaEazNo+nv0n2vPpZvH+l3ZFF
tVDPDRv/hOPxfUwZCMmjtegCE47vmFdbtN7wtKGPwy1+pf9w5uKEnj3aKj0EQCjU
AAgKpvlBDGd5obtrbosvcaxR9+t+yXEMHx4nRNTI3grR+O7ElYG7UVz0RVj3k/Lb
1wkNyRNqhHIuVjpuFMTvkXpa7rTEbsfU36jnYdiOMrY7fcQDfCPha+NUgxhYltc6
goEYEdu69v8/o/4mn/80NWlOdD8xmdHuJrW81wF+tVkCwkPYAAenhG+iGg7r/Kzj
dp4aihIIFUxeRWPJFrirUFuSb0yXfFyI4Bmuhyx+rVwsYb1iDB+paHYBKhyWEAd8
eM2S7wCJySjjxHZNCdIcDPmzX7cbDNa3v94RE0zyecvqOK00yOBHf0fqImaW5JjA
WtRWzu+hN00Y79BYuIXsOE7qMsbi+Vgu9Y/+ex4rsN3wABJmpUt+abuARjtJgd6z
DTncO+5noeaNtdiPms+70NJ/XqBmlib4DtPhn0p8Td6UKbVeCYP9tlVspgiICvPl
use1UBrOgwkYfTy6N3s065wxL69USRuTW7VL3j+KxkP8xu9mv2UTvqrsTJLvUr+n
cRhvda/WmZgCDTANdbIbrGibS48fitGBRumC7mqsj8x9CHi4P6HDXwIsH8pJuR7t
bdG3SW20HqZ0wLV56a+vFH6AyA3Qdo3f0xfdPtVgEv2zHKh2suZUaK5YQXzmZEgk
hUmRqQnvwYQjENGOS6UJlh+mDoTkKYic5WTu2S9Giz0KLU6v6trjc5wxo+wf/JQE
pv7AqeoqrDkO/3dbEf+JVcflX5Gz3icaPPAzVsZEl9qzhyR7F2YkdnDkxYNkfUYR
rS2o+EnaNdu+FHOCEXZ27Jw3bSPmbXckCjqBuzJnFnV8zjYxrasYL6jflKa/WCCc
u+NJG7ZLvsun58kUc7gGcBygvUfecQX5mQ8ZpT2iqgRAGpN5rNs2fFV50ji2IfWX
zT0I6H34pk+TuK5qUP7QZctZrAolilbNaoeuHrmUH/e2qefQDbxV5DNLcL7VNqj7
h/sUnw+qlr0HOmNrG72lvymvM3JHGoJWTd42y0hv6KIoMcAWZiMjRwLKUYFVakAO
GrzbALxwmXQpHczwYSn1Nif2ENVmXNydyQlbeEvK4LF4G1sl9q1cZsjVqJTzLBct
oN9RRtxkXT5DZjNuImsEpHAFdof2JPOnvcT7kdCL8IMmgjKIi1jjtjw7NJvRpocc
NjuNSoKIObC9jrS5GqMDbjsMhkRNb7gJzQonoswcltd4QibsnQHpD2VBUDgOT0Lk
N81H89Go76RCAexvRJLWESimd3RjrTdZ90guOKHU9HVRjUlygweBUQwa4LH/N5EC
IjWIsrr3FtDSCOvV2P+ti7HOTq9faI82EvKW5c+tZ6NwoELzO4GVcwU/iy42nwtC
n7GNFt+KcjMXUCLbJBJCQfO+uuiaemIZfavrHepHdmutAeMTIsbJwAhZoL+m/Me3
DRMDexDfGtO7RRuanIhR0BgN6I+doiTGVnMy/gtfTHt0vfNvqqreb496xf77pqm0
jmty9uwyiDh4aAiF3GBQIL3bgOzG4rKCgUOkn0aPI4zqU6wl1qJFB3+1rMqx6N6+
SLJpjYTi0DQckGTFu9g0CZkw126z/43Zsc0sF5uzrxJpkIVNIRf3ydPFhBRn68Fz
B+U7sf5avxpEssVlvNlYTTQ1KyLh9jNRLcXu429syQHW2hikNW0lgGr6KuRC1ZAY
a2zqPEBNhJckGp+59huNmdd4S8mGr2hmiWtvjNtDi10eQpGbn8o9g7lnmoFEjToH
0VVMgoHQBJ2E+rdrZd+gq50l37SHlobJSc058dMqnfSUHiVVh43blEmDYT45AMsN
v1yFd2LooWjT8KeW0WOcQizRyWR5mHCM+zcW/zGpH+3pN21wsLmTIGA48fA+QkEd
tTzKdU4tNaMQCWXPPgXWVhaMlRvqBoiGlWAeJU43RnHjZ8USzV0NF9SeEYYRtRIA
j93/5Y7W3fVmyiulyN4AD+JALSc4Ca0Y7PJbnNLuzvn2rIIzMQYA3r4M7AqdETT0
M8HyX8RJmzlfIVOKAfC2mVfVAnbFVbJK3L4ihntRjzt1URWVx1cg/89wf9ILYB1S
BmXxs5jaPFx94PyeflT+BjxMfe0884McZmyrRZjXkxTNSNSLFVzzN5zW77eCg9ZB
D2AawgLifLZhaAr0bgnP9ZfvRrtFzLXJArZxdmzGiBLcpag36fu3zIu/7KiMGomY
w1BfJ41YyFS01pPpDH4swdFo4O9h6LMZD1In2Rj2WtxGQmjr7rxEba8/2AmDt9zS
6BKKYkvjplstua6fTgE+ZHibNgFc0YsipvJlzhqQIzAqWgdqv/4j+tgtfTUtQvx7
e6fa03Ok5231rk5Ft4Xq167shSJ/iPyVAsZOUF7r3s80ZAWtbM243fjPDOivVDkZ
OkQBuYekxxjO307O2RLPwaG9IPLFNR/R5St/t2xYU7LUZiWxIW0qEzd3Nbwsgt1V
v+FCJTngkYXzxhIyAtjAUc6pfdyeJdwDyngI09prjKcjpU3E9nvqmeZEGBnqNdkZ
AtswsA0n21FJADW4hKkqtUmKCFSSa+MdFHjLbcM6ktrtTJJnFGqD0Gu7X1Kc99nH
J8A+YvHbQ7HzG3oGxW3vRC2YxDjBTCZ53jZhOWaX9lvepT9s/yRWA+sS3r1brmgU
QsQ4mWl4wrMynCtJmJ8ArRCxXrLTSsHbYiTxKuAqH08vA9apOAytJ3ZjU02HApsi
3ZZu2h3J6tzmYkpwvFEpgdyy8SRic4OovNBiByIEo4NdW4N3GqGu3m9+8ln8BGak
gbTlTpMhrQe/iBgHSgthXSeTz+krtpckRQUx1XfpKnuZH9+7ds/5kFHeruQocW//
DwacpnXYoVaNtRPrmZe79+kYHc2O1sniY8awWXODSQSFFKMKcneVwmP4psuG6YY9
wxF9zn8ezptW29+0LJcBp/2zCEtwLeklwpoLK9V6o9LXvuOx4PbPIw7LA2QSW+qF
j5VcSVYCucoeJk2fZUQi4FefMzimzYO88epLHobj0KaGQxadZk5tUuvs77YUehVY
1mCzcsTJaSbOXUh9a9ihXZvkaOto41r+DJGDxVvFp1GjoK5G4ejbXSHxqd4+68kw
W8VwIaZ3TNdeoKLxwX1uCFmrsXFBpU7UqQtrBSOH3QgklpCiyIzT71rvFfqk5FEW
UXZyJYfESbgoKzvEDB92V27YhpT4zMu5O1TY1b5iuABsYUdk7LqA8v2kRQfAZ2fD
1aaW5VuTwGXNnzDOwXSsJ0PCDqVGLV49UzyQ2JkVh0zyDo9fYLBWcgazjsVKSz5b
RjavEo3bsNlGSu9h2rYbGr3S0ThfRnznCx5hUP4mtvOM+iYO6rVSkDsV48Z2cMDM
wvSq1wwtrOxHiRJwBh6y8z/Yi41/AlPsQAyrYeHBkTck7mHh4vOLLbjwIseDQVCg
cjjO0KrTcdXZHmdnOPc6fu/zC4GnfmEddFSXp809ZlsTM0VcMTN+d2xVuPlCajKA
TlTE/ldteyuMgC/KZ0MeI8SRLSXhnVlp9Stf/C5ainZi+/+jDOaCcD5Pk7MGiRq5
3iXU+T7ZtgSaZIaRbkY6zAUV88X38rrXtRzZKG8rBiFSzLGv1AiwG+5itH1BJzIY
q4Pb8UAXrZxfOmZFUcbwA/TrjD7PbXG9rN2gqKiAktNyhTDGvchtObQ3RaXzBQBo
hJa5UnulNU0wc8rhbH2JrNdvUacEh6T70DundyyN7pArCWkYr6Zp52Z0PaJ/7o6U
bf5v/yLYP5G5hHgE2ue/LTp1H0m7gNxVaE4MNtXZtILYxm0L8eY2ivUoXS77hLMl
uWDEpfIOnEVVhPKJSuePnaCAUHhoRcaJhUeEGyEfFTWHAiFQWpT6zyWnJStZY7Nm
Mn8ai+qmhn2FkpbHQcd0Wm6OojRghle+cCpu/UVneDGMsCPBiW6wjyvS/JXBOk2p
vXzXiOoGZxsYG/D7Z2IZpkOrqRb7W/mhd1v7L0YEer3+struKbxpRyHV1nm1Ao3i
aQtPbY9jxGd4/FQu7EydKCMitTbpQUfftud98FbxKQ1pKfRKuX8vARGG8mKVHHFU
XWsmnkeRp/XWL2eDFKgjUYbL0OoXBhUz0H3UTmbqhhmQMUgERJSIZV4YUwPTWimw
ep+JJwfmwyUjIZaHQ+EHr00d/uhOOw1jWMxOb/oIVT+5q6RywFWRCwfA1PGrLM67
jCSwurvpFg7uLJd84hSCCyYtj/mVwIhGEygGnLiHI+fGIaTU/FJO3h07bSzan1zG
lFFFMPgFPO33cHHPdNxumwpqm7YqOCpJCHsSNOyJwJkDZ/C+OuMCPx/BYAGcxEs7
do9MwwO4hifK3fXq1Kk480Iwhc026BgE764zWuBjbSas7+3NlREsiPa9yktXR9lb
pbUOtw8cdkuDJLqTiXdlUph2W94bub21QGwgL6KO9wr1uUwdebbOv6n38Hz4Fm0W
+wUOkJBFsP2RyGNJN4NGD/l0/m8KU35Hq6XF0tv/MV+AiCt+4ipbyaEueoM6vHTw
U9q/OzM5/y467TKV17OuAiuVJ8izAXeMQ8xA0rK5/zYCffIjBVUaAC34IKMrrLBx
/bs9X/rag70PZEbwGn+x4lT5UVKRRz+TKg2MOjk+aNyHEaTLZFnNJMqIiuC3Ijtc
rEaKMT0Co0j5zhew2qIR8Xv7VYMe56hIczsw3QI3NpRXNf3i/d1zHDTrLCWjTF+J
exbmsZq1Rcgp3q95zK9HRBEcoXAdehxQGWYwWqCAHfvQmcZV1wQmPYZan8GdJIpe
BJ5vhtzrs0qoYtiU3To3Gs+/m1mh9aPvqH8NjhwQ1e2rIBPUZ7F9v+eprHoNubva
GQwszRhudP9p3HTA67iVnghQxk0fuX4R6+BsXC7P288U6YR8LgUaOrAWMKiXngyZ
0PBJv4NwujCdU3Q6dL8YVoWaozHU89kA9KM89MMsQwARfRhCjrfopJbWV5/QG/ny
jdzEAxEsw6s7jLg04RphCPYcxrYOqVG5Bf2m0QPOSsFy2Wl8eFSBYG7SWMW5M0vc
Ut5GnHEqRLb4acQj0hYd8Q/O3+yS/hrPRc7NKbv4x777WMLC3U5TIl8VYha3Pl7h
3lRkTtLFzD5SaHUEXzt2TFNNN0RZzDXzw9mVeDZzzcRT8HNiIzb7WNSHN+CDKpbW
DWOYA65jYLILuKguVj0qB/Y1eUp02lA4vdKLQI9n5ouP6y6+WJV6yizp/9vF3h/Q
sB8LXtI+gdZuWFNS82aUDFmcKIHoEiqwKFHh6oEG4iv4vBc/V+RYKb/gXoef5c9B
lB/mwOij0nEBaOM0rMkTFyDMFsLT3CKJAUcwtKIzsoeEahrUKyaEkU7Jn2PDK9Vd
LGYnz0cFliUEKprG2Dvcd9q5FtRQVPMWKhODqKjTPOFr7teFvlEJfME23+wZQ46J
IgYZZrXnqx2dVcTtZBzqeZM1KdmMN0SgvTrG97zpt/s5dincTilhYHCXaAQ5vaAD
a1xhcuFeezvb2ibQh3yYd/vvJ0XhbNXzfD801GisbIqTb0+E61+aC+02s6WDUvlu
uE0GkHCUlU5sNFQtYs1MCxKg9MFKkHdETJq9DGOVkLwopbHkHFFJTQXDJexMxp8f
s+zAsZ8osBPGws5En/jpOnrtw6q9A6bjm75wtfGYZGXBNKf3ZyTTnTuQXBOfMMog
da4Uz95wglRnvoBpvEPQo8IqARnexBam6MWtE6CAnEFORBDsphAvl+Y5TYWG89V/
F2+6Vt+twUZ2Lg9zTuL8QLvb1lmklG2Y5uFOI0KQDddieIAkN5od6ujt7G/ngLlX
5gsspBgGS3NSCnBaMEUBXtCSdciR15XDnaiBPOK06ngBHJSZ0xARnbeMWTT7Ceqx
ED8fIEPLodAGKnSBQ7iJzu1SSJHQ0J6KUsrRJw2wpBd6oW4SAEM5St29PdYLSaJe
U4n81LNLzu+sGNSDVXePmPE5GyEYra8OOshmhsPlRa5JM6mo9p3zpmZM4pQ9SC2z
G1zfus6WTpBlmzaOXBgiye2n5CYiJqSFMnXL0SWcRSPfRDfamz9RU/CWfOh3vAeR
4kb1ukBilEETrShvBeqbxe2pl0v9xnUlq6lgy6C3T2apfkks60xzeTtUgUQLoFOu
7WEipLq56/86aA/fkIdJ5WbcYo9bpmJHbaBM88U9qyox/yvTvQw/widghdARCp2G
VFEEqenrGZcY9uWEiaQb8x5rlw2urePLom0OgofxzOYx9C6VJR6Ribt7qzCcH3UQ
8Q4NULJbvxVyCo9eG1jEIGWF7gdlA8vtc1WEtbk/bmdeNva44ZBIchmKTD4G7qhQ
AsXo7GxSj8CArG8TR7kH8DXWEOCgUsRirFzxcSUSTtBo4Ji1W2M/pUKTX6Rp83+x
lgOTOtyAiKHihwZLJ0ijuBnJoage32yFyNAwtPejTDz+p84nPnPcQzQv5peM1DfX
F3HdNgZm/BGjpxl3kLlnnj9BufBNxfqMZi6Wl6/rNMx4s8inTkGfpnAPQ9aqVK0Z
57rjwMV+VxAJs/5bDpLA7ona90FtkKtHXmdXIDmwDAmBoUT0p2yZIV253N6Rl9hx
AX3K/uc2fMS9S7igflStxygOdvNVhROq3/yEkr7TpGK438NWrNwXpjIVZwrNVfrV
yc8eLDO56qZpB8R12jkeQU7EQB7UVhcl+2DiJ88VQNAsnT2/TuK4LBJdu5eD0IGS
Np8ZaQBT+GRsDV8MfqepOcI5oGlBIOHbQewXCeyxQIlX2h4/+7HWO9u2lGjbCSDH
E8C7eHtQvuG6TaD4dFo0bgdG+2/b1pYnI8heIBTu3xpicE9UzDPqz8azjOj5Iqlx
AXJXk+L+ICYWORYkGknlNhmQmdVtgypvjqn+no9gse/iY46pSFj8fOwWHngZMi7e
FvP9Yg/KdupLPwxCzvlU5aJ/CnQ0Tg0w11trDpAWIKpcjD634xb8oFlQtyLL8A84
A9B4QvK45D+pdz0nQfcX77LyfVHhBGwlG2kPLGBIxdTGBqZFc7uS7tmnFPlLQ+CP
jUvcOHJVG9EsP7sAeyUYaoIzPwCAoZ+yqvIJmTu2l0pNv6L4GYko6SZA3YR+3g5R
BhhpvFSBPEC/0O/kBGzIxYYXBAYgKZWjVBwT0ckQjqQStaIeMFw5e0wmv036PXjH
Q5etP9JRLwlyCNc7ZKLwB4xR15gHMJZr2vUqWvMsN+NbYMmJvfCfTeiiKj1mctgf
w0+CcirrA0SRpt6MWL02SEXwKj33GbK5j1LsofYoMlD//7FcTizy7E2Tnhh952yw
mGLIDMlC3QpjjaGXqt22MVdUWk0pGs2UNvNKSJ/IH57EBEs3+zxaNe9d72ojyVgl
uLRrgIjBKZBOjFiPjJB627hHfo7ICDzygDNGeDOM9ChxI+BF6I46B3Hr/qEqPgHj
zAMPpOWyjGVBTaZE3MnxVeNMBiudCsB6EpUrhk+9Uubm94QsL4iPQJ2EFQ3KD1Kn
tM408LqymK+g9bymlm60/bfjziFGJY4uJHkSe7Ych2/98LEo4UIjntTDNzgZbkSb
uVFy3o3ljjYNJKTviCfRrouR8evGkAoaNR1dhwZxp8wFJgGHTCiTiA1jCm6xeVwn
wfgRSOMzsKEuP+1h7+nT4oy7LRyzLE0ZALD2hi9WeOtBzqmH6Ynw2XnzEj4RQksU
FatKjkpCOgpciyxlCVlCBJufjfHakuGOC4X9CnNNmHPSEGs9Yvku1+/7aqxD7B5D
3ceJ7CDaW3ns7TrdajJF9heEVzHuFI4iXrmeJ34VneDxhQae80o19sR60WTfNlN8
jSe5W048ugqexPLEOEWayMfhVreJASYyO0+C7buYB3qorTwuPKiEgI30w9ULTfeo
Z6RLCpfmTHjybWS/Axje1dQOm1pQAKt2BKkkgbexZYfWTttVlrWRG4YfLC/V/WAx
IvUmYxd4WaB4NQnUaMabvLCyh+YB3Z/sg8I6BXZvKGHhFQqeGcW+OSM0WI0f6dIg
W82VYiwNjen1/STLSV9qzICswHi0msyGAK4+cmGmdO81lQq8f59b+NPoBCK1iE6q
KvjBeRQaqXsfvl6URoiZuPtIBSbru6zhBU7Fwma9WgrGtT3NYyup1Q/4MTx5ZSp1
5lc1gNU/aykF9i0/NFhFXz8Q3Qt5KVXxPExaAOnCZWZ1o/V/6+9xRFzgBjwDz4X+
TgbMP7fmG0vMRmlAeBaRhR/G3fxLnbnrwaCw2DqPCqB9sbIoNVRm/spVhEoSRbSH
E97PC/bCTelNt3N+kx7f8Ec0+guSG76acfdYIP+kyr1r6PaUNJaIEYSSP8lLlpBD
e+WQ0NZW6cr5O8WlxVtCLB2u5/EVjbdVmS3r+51F7GrWHvAbB09ef5r+zSmbMqIJ
0FGX6Jka+Gwo/HxdSntjWgVd+BfBWdtAHwsx0uwqB+TptF1oeBRml7KMYHEyEgmo
BukrvYKEAWKb1Q3Wx3S0WRcNQbqNpGpauO34xLR7dChumrXRRE7Z28p2/9WuodGz
MoblUzD63No+0aGr56+IVz0qNe4YdT9D5+zHKtCr64B6shLdWZ34YkZK0FGZRu2G
63/GYzGaD1PBW4hwI3J/4HKPVdzVi+rlZ1sScObGqEvlnrmzN6vff8NOdl30N4Nx
BqSnTppGiAQ6gAfgKwgTD2+zY2xg0Yay92bMid6O4DE4qLJnvqPFauoGKfITkAqR
wUWcuHRXCnBRbexJ6Z3RHbvNtZCopbt6yf6vagMBTpk0oOd9Ml72dMqvU0czWJI0
YWbtytvGsc9b3ip9vWlTuM89wFGVnw4L5RPuxt34+MfIizzO5oZIQzSo3OShvjWD
4vToPnW2C88x1ydGs/McWDVYuIo9h5BGsCvbDW+3aKMrha1xDun6yUqfikzuGo4X
bIDkv8UczKo04ev+tdCykdIBDtEuBJPPn7GnZeVGTSzVbx09YEzGByxaGdSDYHNS
Sy0Qc96jkgDLjKJhO8A+Fg5nOWvlz9o+TLH5rthaA81SFYFBWi5l/6Ln0mG0Eb2E
ujPWh33/tVsJE4YuV99c2HfBmTkAsCnOI7fnLSvBaoGyEydawiQVRWGK+kVjILSk
F10yz2Xuaj0SPDZDIKv5wCuQXZyJd9/O0zaiHskWZwTAYAB0A+ck1ZCzYVVuzvir
8FDRUqZS7MiKjlcXSXQWSbro5ybY3n1jSrzJAj7Oc6knUSWHGTixAm2xOpjqwivb
J2aJWx+CARcHjxlfnoLFqZS1S96stunPWm4b/SuhnBcWA/lcijPY5Us6EIpxZPPu
W6CcUvW9HJ2I0lSuCAjMgz11i9KSks7Gu6U4R1/NZV/MbpJLiHWVtAsP8b4/ES6O
DJ1ZcRmgAPQqigroVbb2WdNqNXlZEQWkQDf783gqxnDVmJRo7M2S6t4u/t8pseAo
WI2dqRk/05A6k2Og1axEDI/S0S05869W+imOBVoA+b6LUtUTgfiWJVaFRfroz+Wg
8mfVmr+KHMNDrwjkFhBukz2T444Wp5S/VjwUu2+iBTCiRPDhM4tlXzvPzL/lPCG+
IabYtXx3C6hw+ewuJlKzOaTpDSN+tiNhcj9NXRbeFSvIv++dvLrjReIEE7ahlzvY
NpQ7y7jSRjXJHVpiIGnOD8xYyuHf6P0jLAnYukx1VwHCqZPcDp5eVPh356Wc6wUY
NnV/f8c9cV3gd8jCYGXoxfdP8sZ2ss8/RfEM5DBoNqEsLG3FtmeoS34R01lwV35p
KnghEcrGT7xF6S2OLuUcF68752bfIYlyxcMtHbcPghwkPwzwoZehFNaD/H49db2u
DyU2taY0vDzqIG5iwP8Hr2yYws2CnhcvuqE1fsMCS7VITaQwMczZggEWSHlRq1ZA
FsfIealJs8AtSCyMgysWDbe43jWImLaT0q0ml77y6tc+pEC2/ZAFMRS/QjcxjuyH
kTNv4v0JcVplk43BArsS0FHFOiyqr/xc/PpU4loBuPxvCr7KFH+Kk+PQzPjfxXfQ
wmRAbHiKpoxAT6tJF5BIUNYavYC0qOuy3Qzk7i4AxaSRGE+kLOeYug5pBJiEil4I
D31HbA87rKvJ/nHk0o/vt8INFYK+yMEV6mT75LArQJrSYGvvbcAL7ZgJDbiS7C9a
MSnIXuuNOfz4YhU2DCHKk0zn+tU8jsiwubrLiA4tNVt1Nm8OHvTMLQGW9VIs1FGn
TRJGqqTzIIgEIPzPjkCeA59FcfKZMjGHXTOCOZoY9kQ+7L2OKz1is8/S/9g0G254
x5tB2nMbDbHA0TQKjoFrqysMqsWsqHCosYg5Ddb8tjErP2uvDFDqnNEgNJ87NPct
zTf/QktxcQUfYIviUL1kz0+1kDje5CsMgcIajX0Sd1YY4kijEXdE1Qi/EYZUikXM
rvkRjPeoRp/Xj+SHl6M9cgi/mgcvUIgQhP6gFnEvMbVjW1HWrNaBgy8ROWSaXcYB
xfxG53jtAMPqr8zrBd8fmeDcAHTib8s68BK/tXY8+CniXXllihhQPDoUXaETV1qq
+CUxmMJ8zv1L3t+rqaJBT4CNJCT7PYkv7iTLNhzcJQDjt+aENTuDgJTA5LCo12eo
qLn0R+8HZHBFpg51xcqzLqgC8ufFUhZA1//AQKWcDIaEWC8+DNcR1eyny1zFh1/W
nqlJwltNqDKslQ2eMOBfoZlrLyrnQUqPk5Gu0fQFnF+Pql3QEhmI+LCPSBtr8F9W
8bqA11J9lcfhHPo0/rnlPYW+YWTeoPpUg465Qig8Jxqf5Ogt8OtcyeWhi8sqX8HE
3rkRuFDLBrdJWKji84LiqHiVicDhaaIA3zVEmXAby660yjpyT9pJaeDSbQDxzbjM
+yOvsSLdY+eJ0t6xu+9JZjAPPSgMr6D++ZcdtG7TWVkXqyV55orat2Q7CG5u0caw
ig5hDZe8Vl8DPlUVTY25CTb0DnfjDfEtei7al8UK0E4lfCy47kO4uVUvhXVfMt4p
Uqv27IfBakqTDFFBhWpAwqzlRKeIBqJSnQvz9J95TXgUZK/h4ZKt/Mjtt+Fp1U4w
auheqX4TsHxVDFJNJHLSFmFZwOniCrQyBABoOo3FW7D7RYTqdiGV/eDDXqxZE8rB
dOnsy6WddaEGKmrbmgH1tYiPJtSR+ZlEMZcswU5H2t/T16GKnEbXFmKq8VrgAsz2
fF5n8giYTRphf3MVB4CJd91gHjuShYppfedbwckIu264Hh8u6KJwAAU37hsa60P6
O4gpb9DvuABpIbv6FnqVcVOg6YSuKaIIbz5EGius0BgGrI3hfWQigJylWWYB4mr5
Vj+g0rW50Vtu056bvcZW09loi9RsQyruUSoHga1yFYdcF3dLEav/FWCB6J4sjtwA
8LbpiXPkpfM1/TN4ukSGjq4aK0gCzttfzafrJ7xolJpSkxj7LtatEnRTwiLBQkze
sXKcvpXsYO6hSc2Gz7wXpKORJVzm5ss/aQQWehWvGEI+r9qwmJId1HIUPVq0JygC
QzEjBVBo1+tyXeyUS3MBpY0gN7AbbfbN0xbpkxB1hEo+8/aB7rU5KXVth7VcKoWo
mYMpOVNthjzcheHJH8QIDCnPFUxJUsRFXOxSxa1+z9f1zc05zePrqTKKikxB4+4S
ZUyAnXxvrzBzHXqdhv7ok7VIuYX//m03tzDrooHjTgiHQaAoYeWPy7s5BY3Kxha3
we7AdVTxB2z6gS22+g8BQnUQo4h1iR6Jc9JfjUx+sEwqPHQ8RpREh5is8s5liNVE
GydgvBv8ZrdXw00CoOB8eyjKR9vM9Qkfjn01L3KGytn2zv2mEzQi2o1o1p7FA9EK
W0wGouEhObpMZ+2McZGyuB8nEX8FUg2RJdQunMJINHSL3ILq51WzIQ8MF3Yw+tnp
ut4GHBMlIzXhyuaJ/RKkWGCbxph/5ydlcKx1Uu1BvCKp9DdyBVxkbSEYv/qj+A06
H5H5Hl0ienNmfsEj8wF5LcJrvNrwRl5pVUHGfaDf77obTvkbENB9nm9scDJhifim
dufBnjetQ5Jg7twBvFn5Apw6Zke4pVH+cgxWgQZsS8gXJQZeWZqrPYmXV8pcG5kV
5xncwWegOXqXOimgri6Rr0+jFXwlsazGzx9Qqkj86fWvHhnZ9+1mq/s9YYmP2KkW
mygWbRZaHeyB441H/HZrRBWcA25CKXDniEwNLg5CWA/KQEM2QgyB/P7lAdP+Tz6v
ZXcTZXhgJpS68iwrpHMte499x8AUqRvd1+WOCIcMV81SxDak9gPutxWXLVFD5xMg
UMweB26eM7HMqMUt/A6fxodmOoG+K+aX+rAWyZbiTGxpqcvh/Wcfxw1mC6X5IFYJ
yVqsFUQs+AB47+RY34zCemHOygZ7Sf6ZKaL+LIJaGLdFjh5bGNq6hJzvgn7LDAhG
dTQjMfMJktOYZVAOhZyf+Gar4DSowiuOe/bVyV3d8AopPLavLliOUH0DzalKt2OB
e9prwhhrX5neoT4wAHMuYQ1Efym8jTlXpQpJBIUX8UWPPViYoFi3VZ8PfZGKKR3P
8xtB6BJlA4Y93jAFMz2SMzaZDkVUns4704y+t0ltX3B6tUYkQYZp5RsXH+9Bq6QY
Jcshupa3bXhB7HHR5FjUqjD7ET6GMgGAzMBHQ1lsnTXu/po7HbSLpmXiSVeuE3/F
Kuvys69UfCc58Ev5NMLCLhbTQwpvrrPF9ip/TtF338aDO+D/W0DrTL7rUBaxi8I/
MFvXr1lXrV1g8Eoq5DlqbuHhNwRxEqFcc9onIpvfmyRd2mw8WMFi7uDL8RZznK2c
xtXFleS/OuEs7HEIDpJhKEatUl3k9khlomwnBJiTkTxvWDh0yHlCALvhtMXqAXGe
5d4ih19v8ehA4pVt/UYv29RXWAvQf8j9rcMPDivF6SviTUbNems3EU9srPaXO1QX
fhYVoB/WKT1NO1Hyzfwu45erzLQGmCylwI6NrWuyw5YpCQJcrPmlwoc2JMgv20LS
+rey52Sb7jcC3y2vwXLs3EbPv3d+ym9/7AqZTYW4fhgz6I30zvKQ8cAEh0E7coVK
ecK5grBSUJpzlCRkB8j20qhg0oB1nB2tDle07PudUg1Z1AVbvZC+aqP1BYJv1S8C
RVXNxAylxVilerzw8CMRtVoy7WJzAV4ipM3b/GxJi6qh61hpQUQcOAoQ7DNfSTrR
sZ0HhuWKD+n0SDdM/4VUIyXENkJHWjidp7vyC+jAYHELxEeKVPth+FZt8eEuCJwL
Ug6bJ1YdlaEtYV8TSTeroBiK0NuAiJFAhfaFzSl2dBtycrXMK9IcoO30LcLmiX3C
XaI2gk/5w5BNUr6ZG+Ok9zSlxzmQXxbhRez/Y+YsYhPTkb0064jDpu3GNDY1o6xS
QJIr5Gog4vDC7RLRn0zwgYoL+RkRb2BfXxzuvlJrjFDReQKR3Y2S5HqVFAsTG6pQ
X9OZYaGOtqEQ21Fwe939pIAJid40wtyJk0KHu5BwuqmFKXhUI5g26SvTHEUb+MtV
a0QECviCrrVjjhHhrVlokNShGnrHLOUvuGl6ormKQeYwPPckH6qzL84GTCFsJ7mg
5gj81lO3VCQsSxui8jZLNd4CpjwRsgEREl6p9Jheb41X04eBjbhuHMbyQMG+GfmP
9ZN7CQ4kLSfOqtsL9V323AdMmZ3n9e41RRcklke6q9akw4h2wJBkc/FaVFq3OXWq
760wsaICENSZbU15xQMisW6vxnHIOqzNeszgIf8UtA1jWIRwhJgBKZuci9BcT/FM
0KBbvpd/KZp/A3vKR6Nq5kGGZLfuRAHtn/ImVX7GxWlZhlk9caNbbENcraLgCd0F
e3jJHniLiSbUdy6OQ9f8oSMsLOk5fjCfc0V+LV6Iu58HKZOE3gLK6jwvvhFpAicG
Z8lf+lDW3RQG0eCfeoeCRV4hm4zzWIy2VyRUlPCDn/UHQ8nBQLzBSWYUH+F3xb/J
LFWHFqKr6SspHAVZRz2yli+zmsZPBDJm4aDe0jJmEukx6WWvfWoMDQInee01V0lr
+vKw6k3WRoJe6wWrYaSW9WDkXcY53wYOYJ/ipnvNzjIid6qL6WHFPzp3d/obwxAv
QdPYhjV58qqL1k3GZ20ie4pdNuhhbTpVmRo+0wfans6OtKnpFT2mNThuA8GRqH2T
xUoy362KA6us+nA2lO4a92gqUhrdINBq2RPN50os3gCZfrgvogRniaNv+SUhgcL4
5meTU6f5AcrD2wF15Vs27hek+JjP84J8MQkh+h/k4Fk3tNbVEVhpw/w5K8I0aQVr
6fh07E28U9vzgtSsbpAtBLP2+QpcgHT+nGDXMjSMyWnMNVZfmhqfJ92VCZxMUQTO
Lm6jev9QpZ67Io093NgX/AsgygDxHJVPrGdcv9iTGvOLjusYYLQ4CHr5AGCph6Qg
a2WBdg3Qi+xB4rqX5bZNOqJy3qREIKQNjk+7mpXJuSNHLYLzkaI0e2OHfHjEq5Uk
M5G5piWUFQ+xjB22EnxLEQvm10Pp5TEx942VzfGdajVAYr64Xkx61EdffZPGU4oM
+t6mideCuVUrAZlyJSKxcHfNGBDRaXPNyOjOw2edwD1o9GXVLRMJ9mzI08HbdJzN
a2/W0MpkX/MrdVpb2Kr6nIxQp15QNleymeYWC8TC0t8UC2CPYAZUqEp9JNOzp6aQ
v5xCrTKOyvvhvBG96VofrUXC8narxHWUrVS24JqxaHhZt6Afl9JaX1RCrcISjjO4
dNLTm2HC0XrfZxEzNnkodEoxTLZ+BLCJAaKt1CjJtY6r1hOyRp6Ml+P9Hi2L83m7
IKXRiGxcEzOQDZwDMNNUxU+ZrvbuBMDbFzXUB1MQh2UM25jk9r028lBSo0ITANlN
LoqOjD14kAR3zl/fDKsphCNg0mTSmpZqiJZUIUONPp3pkbjOvrAIHQdfY3EbxoV1
F+YRDZ3B8AJLIlDDyF/spEgWRIwcet+NH2mfVxY1yKJmjrCodw/SjzTtTAKOL6vw
7Z6pm5T0jAJMBI16A4gabo39ETp2xt+zuusoiW+lnkNG7UGJtND7JgVJDE2HG35B
+3s9IUhXzR+0iSHYCiOFN3GfnHPtlnwCtwlfRYudNJTxXTgKavN9i48w+BWoRELl
5Kc498gDhpqEE9DW9SVhCfTXlaFDX7janSEw1EbGaF1DkijjxF7fwi45IoNAqCnJ
vwrsaYCIyiMy9FOXIRMq5rDvrLeI4HEKC61YwOPytnS4HTeiIR4yDGaBbJJUn6/d
FQGn3UHjpQ4OfHsPSjJmlwWCYr/0+wHkAzU0KC9gAR7wBqKWZxm6DV9XnRdzpv/W
tUIlaFXzwytBRg/0l1GY7BIscDs5LxyoQrA/04JKL+lGAbwcaIcNMULYiO0Dp9lb
a/8dr5m3OvhiK0jrZIvDFCQ3lZ9ZEzvrjAT0BL2BmpZqlsj4xbCO6OEsa9BUeLE8
37JoL4EXmEDTlKWgckctR0qwpPHLmawZYphKa8SrQnE3xFI6gF9JznSeev0g+wlj
vW75YhbyYiY00JKIUedStHCUPISXDW62hUw+dj/XCZSxLFfqLIxlfDaFuOyaOvrd
5TjMeeytaxfIZsIAAGflX9XI5mKV4KQcqDL5cxUYfHyDJ2ZGXXL184/5C5BOOW7l
8olFfOpMV8xrurW/Mnf9tQn0Ur7otCqPUvdWUbwR1GGWj3+GbusO2j2McQvKWwX3
WRg0EIu9VE+/ikGzrwB91JxkCJow9kEAYv+oFZjfTofijvgFyrF1k6xtxDm+ZHO0
AtaQo1XSEpGUrqN5eqPxV+S4UFOofswid529vcSfBir0mdCbXkjOEcfl5otQMy/Y
6LxoVSAjWUvA2XlgmuEUxy/34pw+x3oAH3rvFBv1yD//+cGj1O39lVmx+tgrBuQU
thukaUbuVxYlNGoDBmUTH3xzEVrQpkCORl2j6LNkuASdE8aS6GT0hwGgc++RysoE
jeXJ9pySEhN/JKBRsZMFl9xfYj1cW/cL2/HXSk05sBLX4BsstWIU/crgnwJpOPVb
9Fu/BZqjsM08TJ8nEZTCX81R/eiI8X9wyjY8SLULlhLYmcXFyjVt9F5WuZZ8rZDm
74HDErbRyCPG8t02R4MZLiIf/mUF5dvTzp+HWNlValCAf/rdiEhxx4ZT/2adm4iV
DWms1f3G8lQ3/YxDxibHLSIiMCgtjodkd8ouQokqL8D0jAig0FMLOJxBlyAYu36t
vB+DEOnQHjgTF8dKBRj4DVR2N40WznAh7HWkQBOziH9iY2YXJM4Xt5prcokhQv11
NZx+wZHv8Y/tbEIXOAbw5YhTF7ysUgqxtQj2ntj95bGxphxbx+bEhjZHuzHZqctJ
XRs2bLIaFBoyhB8p0F2UPv1uETQR9an8P9PErQtWUqUpehYTB9ogf/gmZhiiXYNe
dUk34JN+aRdaDp2YJ4CLRErpusT2b2aNT8xPcHRiY79T3hmgRsdaxt+IeDHS2bxe
y/kqdRBTEECpAWXVOds4lt8Qy7XuvAjU/lPfhiZwePYFM9UEKa1r8q8p0eBhUvSI
Cr7ugmvzvfn5OoHGy8nEgpHTBEHB9aSXeAiUDjv1YMwPFezHRLD58OE/NhXxaBR3
ZPHsF0MRhyYkw7iOHIFZ+G0Wlnw88F3VZWvPHYcJo89yiCpWFLWzZRpdYS9b/9m1
1tvJfKNN4Wt6lAwT+mFigdrzLc7I8ISCfVpjIBgN3I7aVRsXsdt9HVLL3DGKEoxI
aT4y9CiAebvWns72F7rImwQdnTB/3qizq0VUmbiCt49Lisf8EDv+L9hRrpxPBPjT
GMrq6CtNB9mH8dAvKEBCbyAa8iNA0tq5acvaA4cq5HjmDqXSYLAXhglPOcZpwlCq
E4PjsPdmNwRgb0qpPesGmoQ54S+z8gkWwQCsVHK1F6dud9KLUqSt6YgS7ReqoSzs
uikmxjhSYysZ/QhcMdKmZC2ztx6+rljps5RBxtKb+g5AO7mkiYoWfQvFH9ZkZz2g
t/bC5A/df1xkXPycYxtUyxV+3n1FzsXtAGlepAsw1zL0vqtz1drOuJC2zNBkd4vn
Z68CbReG7vkgRj2eDztK/1W01GpMmt14XgyAQUrMVuXxGsFgT4lw1vbI9Nr8jm1I
LOBpSn6AcjikaQ/oDm6fkxuNfs5OerPsNq8f7TW0U9CxkWsohVVnXtPoGWGFu7ZU
lrgt4+oZxpCZbNsQtDaLjgM8YclN7pkHm4DbB0FSeuApoLXpD4V8BVSGG/UEilw5
VeFpfVXYg8rT0sx4y6JwPEu3MwfzRYlY4huEaIPNy2bdpcV6O0h+axdKWXQr8LLS
BP8/mO+HwSDEG352wIQZ/1Smd9P6g1qbu9/dkUIAk5CJB9qpiNmevE0ZlZv6j/o+
dy0y0y/EJWzEM72Lorls/sR8RVywKKKbUWdYeOR+2iPAQi5JJy02SSk5FZ6Qdvsz
un9FU5C9D22P2aB9iCbAtueWUUBHaczk0RamG60zpnMfcorf3Vj6wE/55O+N27Eh
ZFF51ZKdX9RhUKnsJ1yk5yo/9DeJkHaiJJ+S2OZA9LDwHkWRxY0WStrDqPHXsExv
/qcMw5tyhS0iFcAvn20YionXE3/FRN/WTO335f7ZIH52TGJX813lBu483TRy6+hW
G7k3rJ89PUQ6JH4cYoZb6RYX4igDXuJ9uS546tujsZsp7kjy8PCIDfCG6B+ncISZ
qI2uNyDx967yiLBwRzoMapzpWQpBU1j3JJ5Iek8sAfTUQJDL3i4P9zgriN6Ote87
UyTzK7T2H/c7xFKNhTPYu2IqheAowOTQSPQSnLcStF0pH+p1D1Dg1BxAJNeXR/Hh
x9SVnfWh7L6Vcu3P9OLwAMsOzjMOvu0iILlpBkGUECG69si/cqmj15Ekl0JYiiVu
uHxUBXa1dVOLSHlaO+twQEO2LKgVi2/x7d74NkMuwDNpP3pm60mb0vZQiSTSkeGX
DRnBcMW3E8molovk8fCEYmQzbbGj4Zqea60Augm5QOZgkZXf0JR6/3pUwvzi975f
ldizPXjUMzoD8uwhB/NsNNFFSZjjFu4/9rjeL1uk3kAByLpFUaJinuAFD3MAx2Ii
Zn2GykgQnix60+spSlGwIbbRoD8pry1t+nWx3PlYV1d2MQn0YmqmOWEcgZqZg7X3
HM4O8yAdAK963bGc3+ZYiuHHDwjim6aW1wS0AiMPId8D8Nxk+iptp28IkorcGvzn
3Vh6bwpmL9NGWaMQ+4aAjJqU8i6gFheTzFdgxiO3d8OusmUWEmlFPFjVjAthN/V6
BuVjEaGpQef86SbbKHdl93bePvpz+4UGFps03dWJ+l94gnv+d5qGdkdXKSombrnF
DKZ3VOPAr/uXvpgoo3N6incaO6Bhq588MnGKHAN98sxTyLO1cnqmEJG6zWbspB52
sGJgjKD1/NL8RUQ93o4/wzzFaaNVlsTfYmJRy0PW8X65vrFJRpdOGUJCAhHZCrHB
Vz6IinuE2Jtma9+BEb1icnVXCrALYZiDmtdDTxh6vMAAjFhCG5O+6cuF8Y5V/0RT
mB4NuJPmp6NerN88480uQcq5OXaeuwR4Gkip8acB3v25cDwqYzU9lCkDTbk1yyRS
84Xlm8KcU+zq7I1oWL4Elxmn1BSDd+E7+uqJxBOXUOFUQPBQ0BqomERthpNmEE8j
1CySEAUCwYayERqAI4KwAfWuLWv1vY4yot4OH3tko+bwXT/7mdVY3VvIke0f5o41
6VxTXU6aRCysUcg6lAu2iRjUrOHGyOQiSVqUkZSK+pTI5UyGedD1Pg2WHaj2vN/Z
I6eVk+B2TqpFuHTP0SM4+gh2l+M6JNZyq6qFziipd7rTm7/nPw9knF24X3SY4Zbt
HCoQuXJ+qjwx8lyne4CsGQUZbdxY5zQYhtObPISX2phPfM4o4o2P0LaKtOf0igRk
0up892LgFOQb0wxoXLExVYlFYgW8gdWVWE2oB51ky6AowwMRmGpIQ4XcyF0SKiPu
qJCW0Bny/3X8SzLB/+wLaO6bQ46X7CzCn0Oy2362FxzdS5Hp1LmzKalkP/n/4Cih
o3J2c4KPTobCtjrTCl7Bm9wHS6DNjaH6k0x+BAXaNAdA4XqvhgQA0o3B+0u88NFL
Dk/ZqDozd7tayW9u7mqJC/ygmnrxPPbe12lyILuc8BCmFTdY9Adq/12ZknDaEl0N
kz2kyn3mdJYB+ca9hFzkDoOFAHVEbo0VqgvwrKXv359x3jm556xJk0HR49e8i/GD
M/41veOa+AERITyUs/o4ScbH0WlGiOq26PjsQs8FuVyF4r5uVYbTEjrAY9zxznVx
hp+2VH7wcdjZTwF8aalBuXEQGKAEFjTr6ZtqioPXENUOSn5EVx02YX83RPuiCwGi
CXJf162C4EOa9FgEbXuCVm1zRwzNVe6bVNpWaTv2VZmZfEKyFCfz8CtE6pw1EPyr
HyyJBnDxyNKkH1O4GF2rnklkC+fHVZI/PjgkDAAm84na4x2tE45sgdUHRInyNz/k
v48ve3Z/PPE2BXj5yhSLufjBanNgeiL/oRcmou6mREO9GDoO+jH6c2scQfOj5WD5
/2tz3b6HSbmaqpeun/TrNOlL2Xv7FK2kynO8ByW/e5xFd4vxmz1uSoObPXn2gqtc
G6bT6QH5RAXusNozSJQ8XpvyPCraIbP8KhO3sARpx3VYgU66MPSmdnnMJ4Ssj/jb
oQjYa2kagqlm8HpaBAc1upKDw+zkNg6w7Mfl7APfQ7Sd1CCuJ2CUMj2fLxb08A8A
b+diqMFTtj3UA5uDc3Ga4OChGeJ9DP3rUjSD6ck5pc1UhWS41bJLsl9vVAG59Md/
s2V4UqJjsKEWWfcJzC55Ydz2+/0jWJmIsNzVRdMI3aa6kH03DRduBGfAXfZ/CJ5j
lDXyXJJVXi3fR98z1FRYh+BezSFdKCSsWKvrO72z3Up1wfvAQrcJ7hTzM9mLYp4S
1/wvdkX5xlNTYC2wSBv/agn8voF5xS3X5iHzljTn2t98N5iTgn0A0qJUZvAnq9EK
ADzYPKDOQi+FskCZCN9yAyNQDrE8aqWpVPqa+ysVPpBTfTLMsXyM9KjE8IHHKHsd
0DkZFAN90IpFKVWzuO/EXT0wPVAgHPvPIlk5mvZ4HtuN7cnvO0M/+7BGmZ5eEuZY
syphTvxS0puEbJBt4xHaBaCQBdoV4hrPA37at38vdd111YWZcUvYeUydhpQUGoDb
6xJ1pRdcgz3t+wuu0o4kX4bCUTjP8w13hTK9QrjyXWo/xTv/XVL/l9g/N9nh5CrJ
SvnBW3L08mZJCzLFF0rmaAnAWetvskOpaaTTTxVDoJyC/g+EiBSGQlvf7jRxoVDX
FnI2t+nJYFXbeDCIfEwveu550eneIBCsslcHip37vf4oa65XFgZ+Wv3nujNVxq0f
+ZIMertg6oGRB4BTUaO0lQawV9QDj9Jg7Rn72MjT4ggWFN/lG8jkSTDgfvODEGMN
o2HJbcftbayhB0b578XeX6V6Z5oa/qRsJF3aOgKJBH2c9Ui0l8Y+rpOAORdNQGF+
fwpJG2YvXcLUCR4BuW8XgOs8tBGBlaQF6YiOVWhu+PGI2FBWUy1BDCGX+6uYL/lk
riAr7a/FJ4O2rROyP+NYB7x84rrJc1DBlXS0/+V/Xd5XXzkkH0N7X3hXOYTLXGKE
kPvbyRWninOP1gSPVln9WcGntDbEZnv219BnMGF+UHU57RD9VkWrbXNizMZDmlu6
euWaQ7GB8J0Atmp5lgY4wiWqKCc8pzZU8xm+FzdPLLE47bj3dJvqaJ86LT8EGBwu
m7CG6rqxc2+CGKXJnA+h8DSaY+7mJKOrSkEZRq+sjlwx0f5E2OfXMK67rNdwwoU3
iXb6bEBqi+S7NFGFi9JwCcP83yfvhMjjdhTX3NwqdwQTBqdXmGIx9vJnTeuC7ZFs
oZGcWuZkBrGOyeellVyNFeO4VUNdnr+FzV7RQ+hLRvI/rsK+KfxclOJcjNWJxLYr
dbEXN7CBHcQ6HqeGh6HV7b17MOuA9TWzz9E5Miqh2bANWvY/Eq3t7DnEfKBMQwzC
pvvqUKjCa8g++DeiUwaWBmY/V5uMuFxgi3WFGwOAvC+phEXWiX+enzE6DN/7kZNu
1g4RwJiou+0F/r5Qx0uTnnjlR+q0yySxFyTDmIVcJTvv0enoEMDEYBZmR0iR/k2e
1zzBkOYyxCldLjkNa87YIaFMomg9zZFLFna/Nkfx6+bMi5d71Gnpka5PyvhrTUw+
nMCaRV01mNoF3RxsbbB0pSlfOYNc2pBYS/JRs1D94aNdKr92MzVGCEJvfNF0ccKM
0GiEEx4pqpPhGPCWjb1FVRjywxxk6L+N9N3EEZwDgRq6c7lPfpK5udQaNlahSmBm
CqgXZjgWGXvHxJsuYKI9Xt0gJJA3P/rfaNiiA+WNkCBWv/P9RfaUWx1WcSwMCVuF
J2pNPEThTKhZmYuEtyrURdW5XFvXJ0tXAHHT0JB4GMAjwkgnwijFoFfdvhd3B7xN
twf3potYkSTk31foH4KxsO066WLwVYiH9bNPliYGAQ+xP+Rv68xcU88akgbRMSh0
GrAyPsFStelx44Ksm07f0damk3tieVVALww0oDactjZnpAcjnIo8nM8khDV9+skC
qox44QS2kM8XW+6J4cHut/v3m3HFGJqsqhy0ggadqMxFkd7A12b3BUFODbCZSMAq
G8FXtNKq+HLkPmh0vLeTRrtRwDuuEFPl29rT7P/9fhy/yWEwZHR7fayU58oYZB/L
GjXgVT3smYssqTq7S5Rc3jdI6kkHc9Kjg/vqY4ZdyGXc2A+DgxcavsEuXcEv/1NS
Pm6BPfxNZ6qQrfzraTRowDB2QH7uVsx5FNFUjX6sBa5AJZb+tHsLGmldpRzd842f
4QVNUtpuR7OkP/+BEoCOwt5S1lha6ZGAgmWmGddobMJoijBVYu2dZF7hqXvzsnW0
aNhR7+2hgNVZq5GjPV+vexGOL5qYaUvtjPO6xwvg2TjrCyyvqPm8kN1Q2yZYgGuN
pxXFCvGWKvLtVhP4lKmJTkrvU1u7NFERfFAmIL7Wb6joXsPaZE6X4X1uwgJ3pnXo
6clHoEVBrAx9/Syf3lqQRHxO5L7jfFHSYpH8vfm2SPkUHYbzh2zITh60rB0Asmog
opttwQx6ggGa2QoXbfsFNWJ4GkFwfuQT86j2ifU7aWHpCiPfPfe4M/HlvUDAaQ+0
f5NzPaMLp52WMfk3Gc/Tup4pdqwl13l8ymjQJvpZN+JZqsiy6bkOnZW09dgW4i/I
5v1yrrXp6W6sdtwEkSMz3CJKVTZ/xmsRxW8gjSJCkL/dZPJOrnWVlriSdiMwUq87
Uu0HYkUr/VDS5ZhGeg1eMvawuQ0RPtJb3AqOEAqxygCEGQook2K0SEfdB+y/W9DE
3GWq0EINMz2If4jSUnEbcccb25gEf2eJq9PqFmCG+fY3hwEh3ZO81MEhKCoIfwTD
kTy969FYKVRV4nSwpn+HB6aIFXr34neubf4TQ6WaPosa2z2ZMgRO0YBmTE3YI1UH
GcRzvzUDaj7ACSEbzH3E16kX6+kZlHJ6p6IVg0elKyamlgDqEk1NQMT15l0lvxpA
cwurq07pwJLQgmHhx4avkqMu7CUNu7RpNnW4ODyjs9fDg+RkalR2/J7eRnfOplZK
GpXGEqNkjqMmTA8fx0Y7mQo4PtsCVixPe15uWPC0wCl2vVzzQ2i5px54ZXhTcV6H
wkjHUxHCsqETOK0p4SC4WR5R1ArPCKWFVBbe+EsXfgON07NLNGN6M0lLABzpFHvA
2PiEeS4OQJS1Rfm00e0oh8Qb32m8j0LsKwM+Ot9UW0BAGFkwDLQC+XF8gGNWzL+N
KpBW5j16xReCMZJ2IFe/lJ9rZr+sjWxluTpEDPpGL/BV9uJxMnQR4WMkGyESNSXQ
BCdNB7VglhcG8Omzoqw78zvOnCtdEH7Wvj8w84P4JxZnrEGv4omvkE2wNL5FmF5c
LXHPYZGd/ozmUaUOQfIf2egjDba8XRmPYp5VnjtsiJuOM3fW7rPRlsUZq6GUPbNt
weGThtNKcTTGXBb4V1y+0G/mPCnEH9iXV/7JxqpAvNTRaktl09WxWAW0Beg5g6MU
hHk0vkGHNx8uy/s2iECb27FlL4hkD1ICghFqZVQ1vSeRLNcxqP3KhrV6b2L1wsTS
7Gsnwe2gjSTPFe+S4jFVJ6NRKOafowY++ujq7oTdAcmR71HBKp3GE6nbOtzeZ1c3
s7M1sAzz0E3RoXhGpnMHP8Js84CzlMxlUl7fihS8FCzo7NlOP+q7WwcHcLAfkwx/
Wz+6Ch9EJt4hk+wOy+7sFDMb1t7ic1u99qx336yUeaUESsOQ+ADoBebPNvZJw8Dp
R0HGmYTeEIfIZNX6KTjcFjt1WutA3xugFJIwCBhH1vnrcVtG3tYrrAGFIwxiIIYD
QURYC/rLrF6GbFONtSqiM7NQMYFjP14Jlo8euYSRVXsuPqhfDXY8mGyBa2ZDprl6
Zj5HZ52lf6nhahtI9cuz5fOKY1xbSGujjCu4koqpP8knDXik/Lnq2zXfkS/Ebn71
wed1pldqiInYUCWfZo3rYbEKs3VPSZL9jPstSj2xLoV+dAoSAkCjt3rsrXIFH1F/
vFdoaQ5I3ZOef6unr9BfvNWHdmk3x/SYpiIvGFkSMjiszwQVv6galYDnNBm2gxEz
pUKrKlhKVNFFec75QM6QB+wiRxvz44qKEfSm59dnMuQlMKQZAUzEX+t3BgHIpe3Y
7SpIBj2714RIZskWf2zVL4UuMh7312HtEshWBcw5bps+cx+xF6FrdcfSvUI9z9ZK
HRtOOV9F82u1QhcGLUIVcLyCGz2WuLlQq5cvCKNtqLHeQKnFC0jmt5vDNQvzpOgm
qbFnJVbS1F1oIfLhSnDdcjr7TkxVJDAEVRpPzv3LmQVG6ID7dQVRiZcktbb1GFS0
5VZh3piAWw2UFxMO8+m4llt36vkXwINZcI44HSFUMNuEiCI2vFsn+XI+ktSS3MTL
woTBet55Yvo6Lrm4ugfsLiTDyoSYjENkg4Vj10g8u7T0EfEy8pnHTDAH8kaNwLkY
w6z9A0ephorAEuLc7smWKEWmsA7oej75DuDebEyTpiyQQHnrUFDryhbcMNzDN/1Z
0qKIEX1RNiDWoFLG8VcA7bcsjXGqKw0S7kZ6cQFqu4QwlDlL9ZGIb585DsP3MLXQ
VOXIqGrx5NIx58E1AVVfim1W6nja7v4KvThFbVLgQF8VzbMBl/BIwXoIXO1GnMcA
/1R91tsNEn3lme2AXMQ9kYUOte5saReIHu4A25qS+wZAgq27+/ZVvWFivcZ/s7mv
gGwNz6WUKdDp100PF98DSU5k9HDtNgk2lf8ZJWAVUCLCkBQqOYpA6cFDJY93cZbk
MAF7J1eyi9qcH9JxFGcmiB2o2+mINS9b+q6edydEKkiQ1SMbVsP7CDOx1R6XHDog
viuWFnfsTicKDAOoyunR8XZ5U5lTXb+IsI7u6YruH6I6bA/z7jtZE8HpwA+TZSpx
TgCthaIAvvczr8n2wylG+KephLFUx5N7H8aHuiRD//AHPzlmz5XIkWcQ/iAsLXr8
TE9uyZEHYfzKA6sAPlvrCxCRSXmcufr3I7yp7LBbZvA3lHT/Cskzpp5Jv5lhACSy
kzTeh/04uLjXZcDSnJvzsNc9lY0cumn6tAjRxlJjmrnTVZ2Ahe6Skfd1HoGX+h6b
aZNJZYNasMKM2jN/XpYlMBu2kgJQQEv/ymfPrx392Ub4JpFczurgGvnd7KyEnhsW
ml9wpAVmLxPu99NkPzzmqsQATMCS4/Ip5wQNiTM9p5NBe5OBsy0IweSJQunTWI+y
QX5RNITXxHJxvae7ZKsknlF1QZ0dsFp6IyrbobPb0kC0UbZEtE9+Yj/fP5D+Kr6z
k0G8rANdjb+rPtn5urJRl97I1n9sf1fdSVWdTTTut+69Iv0Cm7utVcVLGe3qSI1A
ep9C+9cxjPqGmv5VCTOyD+LTyR0/qfqBoYrSUQhB9WzR3bkZ41gd8vsINUClDJeX
lCzCnYtBXuwgOPkvD6A8IzQR3GpwdcPW1F8n4Vays6XVv0c0ZGLr/Kg80Q/Jd2Mp
p78Yl6EvTRLrIKJfMYDTk6kqg/TwlE2sMdPx5nyVEG18ozfSxMhcZvXzyVynIAYV
GSaz3rsZKIqQrmnMd5rm+T1NEvl8u04XEmKSOyGY3eUJICTwE2Q5ez2rL+6a7Nys
OwZdTihZpT32V3ToU6iLJbvJm6kbmaFA37pJQ5RyhtYHk2XJDvTdo060Pi8NBP8l
W2fRPOIebMB7/VLjwn+8p1VfHgRUJ8xPpEWSE9m4OBbjw2NqmTArR4nmMDr/32wG
FD+NJdGepa7JgvyF0cshBfwxGnioMvUbNS94Yc7Xw6Dhb3sqwG+GLCIo3Tbcl0U3
qRzUnRsPvSuTdsdgBsnIdbji9QVOL47u/R6pjTCypGY57MQ9/2uDCOyCxQGEnDsN
fp0M7bezvSB7442nGo7DxZ5WTU4altNKeoW8WIQgo02iEJXAQBJsO+c81LcEaIOM
Y5VocbKjA20gO+wZTFj/pquzHqPGp82kfgWtGC3byTJioNeoDmL1//oua8ZXS7mF
tWUmf2GbTHA1KBqSmkYXE1weiSGxrJN3z/c5VcBx1afAKAsFXX2OCMtHfzocePjI
R7+FVA/Rl4MR2Kv5h3129NRZLG4kWFxNjk0uD1gprvdkUNRRGkpQk1aWjyhfBYJ7
ZCBOKwHPi9ybSmS3kH6Xmry0EeNW7JNERyP5n1OPRwhtuND0LZjVIw7X6v0FGm7j
CzoF+jgiXaH6qAvFLRCt0bIxJ5roiocUNEy53xrGK4nUXMEC72CAAogq26Rl5kEW
u9icJn1tbL10hvsa8XCZtkDUg7zt1ffYrC9+O4OIC/ysL8DSPa2D/O5taY9RMzK/
Bvye3S8YKVCe+t6pa5KoxWHiW1YrsNZhO69YFiNoqgesqzyCVzarsWSAkXCU2oPt
OOBabPacj7KwtewoNhoo8uZPQHlEl8aZaq7PmHDRS7rYCUVemdc2Nxfu2vZSBEQY
hAPEUK1leB2erIMSj8IJrUiN4lS1n9DMNvj2ek6fb7NsQanjEzEO+2PR4xME7bRx
AWu+0Jj4cKV5o8LaJOz0SQwuYjdzVYa0E10ocAOD/XPFf5rIPWUbde0RX8U4XvXt
YnzzXUHAR8pp9ibNXlpbmCGnXQnBvBHyRJxLo65ZyE3PqquVkhUga14xP9VIGJU6
sjnOQ0R1ETTr/M/EyupwDUAfmdI0JyU2/Mm1ugtslZT2NMBRSA0tklgalK/w5TeX
PweHv1o+xfgZo3OQkxyUzPcXt3z0vpqe+Q63cefCGCVD3HXuwezir9hX7ZpGTVQY
1m6QvTsEgv+xEwaaOes9jMG/B/7951AyESQfr99LXt4iM2kwYqy3UGdrTu6Iu+WX
8OLpiniVP8T5mn9iQroxOOYAkuyWJqMCm0dOPy4lHPBwXiDf1vM8q0myxA6UjLHB
YrHCasFNUbWml4e5GTxbiqc2Wae8f6402pzk4PJHb/wH9iUJLgp9Zp7GEHCbZFML
KSoWZ1bGa9O2vmbjqrz+RAHz4EyT3VXbyPdPC6j/oLqO5Dtjtf68Civkw12n6CKt
WGhlB4cbZe5mFyezYyJ/mTGRJ1DMTTCmD1IIF/2aK9cLafkJGgxxcP81S5jIo+LZ
l4+Iq2fX3UOlAz+9sw69eRwaqHehV+tX5Znh1zh7R8xOiu6fewzAtcl29sA998TI
6iKGezZaXZXWx/cT3zf26zlivgP3i8BFMDPgUZE/nF0nSdWHURFUmj4b1aJSoKrV
o18TkqO1gGbS337W0qbYkE2/h0SnBtAUY9JGDCyRlMNb3Eg0Xtg/mL9YllWmBrGs
kySsv1Q5sna+gpPRjXh8NcZ5jp2pROaNROzsYTVqn4n9MBhqstSBhEOjapsQDPcP
alBEt6DG9Ydkc+IguBIc85CZDvdJe9QtjKY6yKPCUaTTaezOEJudqg1h/7xGenGT
rMK0sdbWNkv5kJMDcKceIgMDrw5WTwHAZRPEOw2k3G2uCygJg2WykZEjjwzCWMq9
YC2gJ0hsfpzf6e8GMYB3z9Gwi4mbDqMS7Dz6EIbkoJSpGM6+CJaBXc+98Tw5CL3X
iVGXO2Pn+eBktgT+DAV+Hm6EvOvhGce8yRenJ9KPMkYLFTv4DPq00U0E0w0Ds5Rg
zztQOep7+30ueI0oSbLEKak05U1Vt3+tsRwGlztmLO/RazQkXTRbLYVmDiuzuS32
YBflml6Yl+nAwb5viirxbNqFJql3yQo5ixugxQIk4RCO1G8FuQhfZx2Wz3ZJdDks
NTsO2BQZI9EktB4zCEJnIHNRzrp+SwepZ2kpGZ54bUFrEPXYh4n0DecdhJaIiqoA
emsETv/RKWTItCKSRw8kMvXJCAJi7YuMMpSzWQYQnxMOwcHcKXm2GfAqu8txHr1e
CRngbZogwHLa2LwH/YXSTsUTsGEu7Z9ZIFE08R8dCRKg7Y7Yd82rQKeVFEt14Tp8
ic18FrBPzo7N1iFGOLPq65z79sYKYtrYTYxYlY5eV61RI0QNEdXXZWR5qATjyDcU
rW/TJOjqUe+rjjm6SxpzDg/LCgxW0QUsPkKG2+ruT0GKnOJUoic1dFUHdyM9c8Cn
y4L55srYHLoWcnUutXqVaaAQr77wsqnyJZJ2eCw21VkSWV2tHbhtGvSEMvkHWD0h
9pxxes54VneW4aQZE9plBGMAgNc1Cok8D7PiXi8IP05ypWzM0z//i5duaYMBtJuk
ice7Be4c5jST4eM0PfsRBfZds5QR1jhj17RsEnsr+TepKjKIjf7uZ6PkEADNdBEn
EO3rDqhF0nc0CPR75FmtlqWm+mq3fMsb3X0ulMVLhKJIIXrbf5N766z3QYToEX8b
5ySpaT/6xVlCr9vBC3bkN5Sc+OAy9uIMwxbU2eIW0+8obNaAfC0yVZWv4p9Pv+nB
vIf977QeOCvr4V8UfkLHXD4w1ua7kB1mrBjtvCXMyEus9szpVpK7e4O8zysTzFO5
qTu8EK5U8wvu0tJ8m5ye9lZ4nm9y13PfrrtUuQ+Zy5CHKmjyHdGW7BKIDYjaaqL4
jR5F8Q18AixtfllmAF4eA7tYeIigJIDXtCnCnhFajPvXXmiG6/8yUfB9PWGhBSuI
QuO2VkmpHtk/v7vi21KyC7FpiIvGVV4qrQKxtHQ92xkEUbNFmr8lDu2to28ei54V
phv1I5jj/qvDnskg+vCaf6yJBc3/AC1Nif6uBRCm8Nb7izcMxtrHH1leKY73Ie4Y
SENN2VIb6rCjEtyd0uy2JvVEgn/DCgD1LQkklrm3luZ+C6R0AGBqAh5taqojGtQr
VbF0zjxJabeS2YngCrjWQ1109+K0tIvwBmBuW7GNHhXyEO+qF5Wm+nq5MFFqy//m
tOc1a5KBMsF4fv/YitnI5aBk2Ahn+FTH/Z7yJhKjSojkbH7HM4rmTQ8qgHv3Dzk+
pbie4z6TCuOl51qdOwnSSlRjbBtwkExwwZgkR4SCC43RWzVI6IosIpkuGxnAJcZC
qAlq/KKccJ0qTdLDJ/HPWrMCn6iJKfKVZ7oCov7v7E13MuYfTfnYQSjYHr4sBxXP
orJXuxGGc0Fw8mJazSBd8CohOsn6nD9lai8R7Tm2D8I1SnepMDqzXxz6CCyN3Q5Q
CCt/Fu37nxBWuet1Y0l/dU9NtnHByVIvv+nCqBU/+VXKvgY1cQ4e6QBbeA+YhlyL
s1G5esMMf5DD9thuBTuVfRJ9KpN5zJL4Ktc5DTiCuLQby58SSbMIYoRrvDTuGeul
7ErBkASwd+oY9jt9sE+vzemh5bmZBMeQwY8AoLnDrgODxsxpvTPXaATTNonra4W0
89x/E80nO3bC6Z6bcQ1poQ4H8RFc7FY5ZTcRSpKtW2xwQqZAXIarN4WsHTxS0wqI
dcLezSHqVptyNcU8fwCenkQb4kb4zHF0xF4bFEzVRNAWtL6vPQv9DbntsFlU3nzl
ocSvjThZj3LpptTqyrMNQoJ2vU0VX8AhCWoAiN5yPJMkCc9bYoWF23mx1QZ0/Xxd
GGrm6UWjm10vxPGPgiCwKzRZZlJw/SuEA5J4iCeOPCvYbamrHwrL59uL5slo85Eh
Xk4g2gAGgwuPBj+NrR9PvK5CdDJbfH26KjXgjlsnR+iaj8ygQAQVSXrHMKrMklNI
pCAgmcwAiyC1fmPaWMPsJPJ1vq12nCBmWhOyeB6rCL4aU4Hj2QbbGNRA9rga2QHE
IdEtMX3s7YplYi4Sj2Z9pqz5y2JDjbPHOOXQRoUTKkDn1wwh9nQLlDCuTY9fc8/i
nFdfuL+RXwS+KQDxcQkl1uYuld0a5NimIuxXrNM8RMQT+zcbj5+dChqIGlxYgVBJ
oyROr3MhtF/6nLs2Hq0husbj9S2FxG3vS6WC6DWQ7jgSr+McZCUB9ensgrhwoNab
BWP4KEjgruOiQAQkGdzTz3eMICY4+2q8N0okOEVoMzWckBhK24YhADIEW+965tkK
cp2Sb6uQXWL4P+fyEOLx3Pi9G6wPeUbLVBW1VYbGB/mOwBA4jzepMK04cplHJDgs
aITDI/Ee37DK+FcHCU2LKRCNmFN48Va5aTEkD1oKv1PXHPvGe7VZaZcV3atFP93a
HYbwe7BcSPhVGN2JkosgfnNkpTNGSLXT9tK75sFvtk9He43VY900NdSLrAKGpD1F
1kVPjsIHU+nYWyTNpUpcWD0ngnZBT+9dkTtLy+y6N6h75wVqsrlnUrvF2WZMY1Aw
oMS4EymdHmVOLyI9s8p/SkEm3mofc3NxkjQ9ZaVBE4si2CsrWTV8l2a5koOdk4fk
Z+0KGKz5LtCifgCXE55RyPau61wziBdaLufuhMcZXvuYZooYbbgcDZi2jIu/c85f
Wvgl7sXaiEmu1UD7wFsrPB/+6xYv+cLOxr5jERvrywihe16TXQBwglZK8yvfvK4O
Z9QsDXz0X8NmsLh4p7gnGdLuuHxrZIxyBfPyd/PCxXcid6YV7qoLh+oHpY4Fdrio
yiyKWorXNHqpMA0eP5fjPcNAFyqJfgfMFCgfxy/YjSOECvAk0/ZyPmRFfhTYaUbs
H6LpQ44HRA9sbmb+dWLz+7OiOBvcOdMLgADeC/Q1bAmlo+HmMrhpGurCtUMgilV6
Ta6ti6Xz3VKXGT2wJILthijHUADhqKuQgDOHq4ZdHNMzI0UYBtaSGpRKlQce0w/F
PFty+4kp/Uno8AmL2TuutiFsu4An/dHwFMs+zyp311Yl7mrKbAQP5go85kEYPJ3+
ju1/4BckTvQjwnLVlNUOImLySviaVyyoFi2PIGXuOuONA/rq9R/grYD50rWnShy/
qQwFGxlk9tpH2Ge0Or0fWa9LZu9WVYi1zRdkcWLGuN+faIc3CtIKEb09QZJmcqwF
T/vxbIysw111Hx0BxBbVs4F8GR2Vbffaeu4a2M2QyK9FVZBbRx8C8DjbUwXQa2aY
p7346uRf+sYOtXP7giwXassh92ElHAbOLnFfaDDTfJmva1OxZSlY0eoC8j8EWobb
6Qvv1lvxlDoWu5V0o/3k5jsnfAXgwl8OzgPEBV2GlRHp+xXhqXRu1CcZfo4ymH6U
1fsrEz4r1/fIrWNsZB87gHqIJ9THnLdwKO0n/KNhxhOzf93ZLggzQPMuJsU6w6jQ
Uk7+XSeFqZ2M2tfdwic2X6QPC2/b3jMy9ZF95Rg4qPHUvogKqZjoVe5ymT9BduFt
u8/6/0eRxNQrxsPvLSKmzXugltJiFJc/iFkAwzHUVrOrH/m8+GZs7Da+2ClJYpN5
VFyxPRqtPv46CWXNlf8PcL5C9iZVhkUUvJe6YdmjfEt11Npb+ntXc3wKwaD+L0Wj
ulMx3xZZGV3JJRyW7ykb7Bdae8CzzzB6zwahRpcUT3F5MdWR+WSn9jF/vCntZDkg
AsnVVqFIX1bAi2GvAH7qLBgJ21MbKisKRfzFrYMubIFtVEFU1h6tJ4o5G5Td47zc
wjpnLdIGCT2Zg+Z062dECHOaamFOSTgji0phliuP8bM5eLQX6zE9lClL4N/qAYhC
NVFUScVfK7xiIZU4zIH20ppjsgE4+AGAb8/06xaYMuz38E1Jw/RZn0G4Be/lt+uq
t8PnQwEMwRBcNjx8Tow9prG8dsKvyvB9sqvFUe1CarzTgsPA1A7b9abmqKfLzoYT
BDZQQaSc8gbgG9moo50thk7oCEmlm/tkhl2jAUxAXy8wxrs16ul3gQeW9QItuaGY
AeBmnTvhM0Gqs2BJ4KSg+pva430p7D7cRPU6QFHHNAm0IoRw3uFvF/YU38UrsjDE
qZKkY4W3FQ21/F9ldjeCUGd3XJnvEPd3eIIAZOnLMpLmDr3MhpKZkSyDFpxfCeJJ
nXT/v9VfjJo7F+D9nGP/VZCQX4/Fab9daAFSojC2vsaptvJpkg1PUDqXSW+zQXlU
IGc3BlM6AHo4J0NUUWEmmsZFHn8Zw3ucuRRhwXRYXuCw4R9TIvLNVyqvSgbhfNeD
HN+ySvRszTPnNvP6G8zjn/SsYBDLyGFS968tz9XhsJBrFldxSgHCZSKDYCSXGor4
mlkPqcxQd7MYnGUxT7fym8qlP/Ay4Gx7ctnhodPJzmsz8fdWjaI5owXCIhK33j1Y
zVLBsbHDXgAVTCrjUJ0w4riwHtgNVxMj7rBhbkFdOxrLYhBg6mHO0TR8KDSgIPZG
9uM/JgVbO0TlPCL8Oql4NT95d8Izpv2N0Eqm2YQ5ral0a1VBpq6OmIxtLRi7xCbu
biV4yFPRNVlnkGRDjYrpgfAEAsFRr45XGr8YPaZAEjvg/ILZf61pQ+lSr2wHRA72
fcR86C8PFDhm3wLG6KF+Kx8blsPPo1Q7XBPyQcV6x5B7A3ZlZmqE3d45JJGmCCK2
jxh2fwBZ/EpCbbkMfv2truFbXDX8Go1rJ1U3tW3t5QQXadENh/FnTJ5hclfpgTqU
meMYeh5gA0AgI1ymF2Re7GycnuRHiKA528W6EjTAvUwcaGFPkF4j7bO8jvGIafN7
7TbukZSgrZC2rwV9N1skwFzwYfNfmfiZq5a0aI2oUjt8Dha7JfsiY2uatrPUaadk
cXtxqEdgcuqtCGU9Nab5sZ9HS1+cb37T6xKyJTxJkUKdgsC4JGZV2xpvqDOrJRqD
akLQlxJ0hTdO0AI4mHIkVtiseNasG5h+dq7NOMhj/XuCssA7wd7SK1Kq03Uieb5u
YnXVopUPC4IXB3OHxSwBnoAUhSBz3duZb9ctb0cn1q3RXrYMt3fid5pp6yrSqmzF
n8d+O/ujZo5Fx5hVG2Dv3w73m+2ioKmaQA4Iq/YnfxuQ696N0x3gWxU3mCd8ird9
uDbGWm9e2YOavbN42rE6CquEiO8GFnwSKfYZ3iq/x4/WxC6oQqwMMzsI4R6SMVle
g4bZooHOI4RUDPZDX0B6nvahKrFDtC827CUdDOiSAf8HefyEIEe09he3lBN+TFwO
iILfjrQRxxz6E8TjysSGRTmWSCOH6fgiUGpIAlAKnT0LaAx3+oo3Mimp0P8UE6kD
FPSo7XZ53yjngr29D6w0wAJWjKECpvZoVPDWODXxpObYdjKWVdsuU/DLzWMZVF1t
9vQ3sD8IZxJznnZHnbzlgCJ5+qu3ZBptmPNnV0Fjhm4eZssGhrXHnHVTCicvAvKV
QBCR+sGzJxo9ttRXtAo/bOJeWj/4RsnJe8QetEOOrow8y7t/qHMK3E1lhLsgsImJ
iuWnYZ3gR2rsSs+e4m7Sq81D1adPXuycPmYGYN3PR0W3fKjNveEaX3a9W1hH5B6W
QblWKQKRkOCo3KjWWaVYrG9oC+BHPn+jv8u6emRCULTtp5PtQZW+bE6Q18F261y0
8vkhPn3SGdgOz0fZ50xAl79Op3+lmpNj1r93a1fBLFQUwc5aKTr9MB/g58qLTzAN
4XymRxZLfLKXpiAB4LsU7YoanMAgBJy0LlfeRyADlqSlk+vACHrzkd/SRmaikg4e
r4FfvsemPOXElNyR7GtSlEvHpXyaKG/nXKcYFWxQhZPYI4d99A50JsSeCW2U660Y
Paid6h/psJ/1P4D8CCxP3z83Q0IOmawCDKE7JhRxPIMK8BrEc2naEj++LS0AlrXz
YHdoEcdffs36zUlpzSFI9kPazoo4ZLh3MoOrZsyxrqERJ08F9TOZHfKQHi5NB9UE
6Ex4ld0iZb0eejAyfSbPaYSo2N8Op/0WNbKPoN7Ofqvw4Sx09x58yBLlQRxkfckz
PWtY8z1RtJn2Q24pZfnYpRDGvnOQJQQU8B+6rsLLlxWizG0L6WZbxKVBFTxUiXPu
wpUAg6MNxncYI95zj+H+itsI5vFwVXsGcwnN81/kjYiNQtVgSWo4kgm6xQebABUk
rBcejCN69gIkm/111AdTnDry0ZjqSWSggN5ehVveqL6yB4/WZupgJrk10PH8Zhx5
Em67kzzoPmNyk3BT/MvhF+KFhAC28/B57fur5YX33fzSVkshHGGZMZZ1x984wMtZ
E2GLVJDAgVvMat2NoTv7XDK4f38Lu6qdJs7Xf0/U4ONvgFMj0wDQu2S5qfm0SqAo
5JIUCiFP7AEyAHWn417I2T3nsk6KnpdkqUGZ8IA+D/Wx7Lqqql7cF/U+Ovnl7Ur9
+UfOT7JCUjRX4Jr+OLpcNIrik/8RIEy5GLSI5+lZKim/wiVT5CIcdEXKOYHxwNSy
Bj6T2zAB0UDYP5pSyrtKEitGtG9ZHQbOWd+ZUk7zfTUz1qEIExs1DBpizLVm+7bN
KLdtTjl5s3E+oKK22MqUmohldBQho5BM935Z09umXPNEShoJvNcXDUD++CSnUe49
ZZzuPHd111e2y/3s76515ZDdFGbxFb9xt5EtMO8zWYh6M/trjoR6tiOOi6USMHg1
eNPY0SJj9gPfEIF4ZziV9qUk5AP77FGTHO9slTHhZ5ZDTS6IYE5jQc38WyP3vPUE
uBvAQVAuqLnXin+SMIm0/T4PZmdBWnJiaDe7bUfckSsCRe3Dn+vmCu4LhOb2QO6n
BszN7KgJEyOHt0hDdDHfhU3eBdX+dACb6Ea6yRsmGv8zd5zMxVNwIiZRz6dB7vl7
8U48l2qb9IpiRcmbbF6ENQslMfKF4qyRb1ro5xPYdEcLp219E1hPrQm8RPy0o9LT
rRnuk5KF9BHSAuSLCjYvGxhk5FgzAv7+lRKxgJq4Gb4VSc5UZOShV+WLLUDQ6r2N
QJlujTH5PSjk9pH2Eso0cB82jasWjHFj2Hue8mfTE9piw7tUCyacPHlIH8lKjX/C
s68cnygeAruOCDcD5QZuOfe4vANseb2W4uWPe0/eVxWVkVz2EzRapbFt8AsgPDGb
tBC5zUIZ37VuariSnBTNd3wx5ZtdwefqAYWKMTdwCIKck2XwhmnpOSAFoLF9DQPD
vRt0XV1hmlR6WYq2GtyXfnQupQdaRDGM1jZk29QIPPJIgCGYKwtKav5DB9lyhdFS
bEJ1ShmvZSa0SJzqX09ehdLfKdrCHgaZFdYRk4KfLrCYhlhmYiRLXpaM7695SPYQ
Q514BJUqE5XEIJIghSQgBVUFnZy+CzkWkjas+esqAbheeZwYPSdOQlFjC+iQ0yqP
+COvR2zR5/d+QVrX7ZZdtlJ+gDr8lreQaj2dj9jHDBHrcLLE04AMQdgFz29jpk2u
0MCBWWK+SQs9o8DSDEN3Sz2BS6H9xC2qD9ZvWqk2+lLcO49LhD93dILlAWRRsnW8
NoNkE3hxI6I8oQ2oQmVvYNHR3h6T4RnUtwnqm+LLNB3qR+mXYdHHpQdoKd05QSc5
V/9fF1rIMoyTEIFNu2DsQdMuMzAWS1fGYjwPetxU/zyDJdlZTfP5GGe5gm9WKtnP
4280P93JKeZs/D/4+Tj3XH72u/WQhyepQ0UUHq/CeeZPbTW4G6vjdZuQwcxI6CuR
E0uwmybjrRKdd4oOzuFb7pGtpOFrFSonDvUMm8e6WzjLi41TAL60qbalGzE4m/gl
6Oy/0BM+GjkTUJidjdlR/k1LXMouZUWZ/XknuEff1FzwuApCyckP6JIMrZLd6UyF
GU2j/adC37j0NYav6CJmsuTISRTa5wfbTeDYHa36icHi84wI3L9A+tJOaPMu+YXA
ivsGy+XOkNdYzgczOCTYEWg87EgsCW7B3P5GywSKF4uSwc7tHUaKZP5dUR896GgH
h00r7SGNr7Om9bPKF8aHIH54Q7ER4QyMP2e9ARGIeqRogfwgYqEY6lW/Mx86Pa63
uu8gTkmOToaft8sSi7uxFk987pOrkXXzaZUxjQzzzJyXnkh5V9fwdoopb9jndyIs
LewFhQ6FypDcYidvTYy2C2+/mZ+KsVWMbOAQyeg0k+DY2k7JUckmTFzZP/2XBtby
QIGjQNORMn7HRL0I9cAHQeSlA4i9ln/wvJdKNvqyOrV0LUAzGNn6nOE9vBV72WUt
fCJJUdt5O4oSDRutTw9bMLgRvdUfujk2F99Fh1Och/vv5vk3oWnV2xXDRAPI+CvM
Vqu0pORqjckBcWhl/su1tnktYuZ0BKinrtzLWhknMgZweO/FOiRPbH5FeHYf1+l6
VR227qHvLexsE5BjHwlA1jWWDZXKuL/xNX4mHhf+ynXQ2mkgA2AbEs1u8LaaRMCi
Jm+evGmh2pGtycjxWnhj6xrrkzP//mkbL8CakNgJqGeeKi0tv5wLlDQtogQQKBc5
FVAl3FAe1I+/CjCnMbkggploA1sTccfiBOsDErn3B2ydbztZ6W4Gf/E+c1yMF9aT
DLUE2Pv7SVIKltfeSg7sKGFnwdGzKqQWpRIPdrJTTeX1+/ju3SOya253FWidTg1t
AVqnc5BCeV0xC+XoLhjvoKT6qMKguL/LlDDDboK8SDgA516fV/JC8Wjz3hsWcplo
zoIZUiivppjODfAgnzYOFD5SsyWPdqLtDsEfdJHCSzsw3q7pQfjTOPl8CZQ/+7kc
zCX0mc/12pQXiLt2ChfJXDUH0KNIcaUP1AZBCwjcBjSmLNYs68eUInxvD9cTpwFx
lNWb56hEmjtx2ogpTLfjJWrjMXVpJZU5BB19Rlg5kvkoGQhJd3M4ze+jfYMXkNa8
E/+8Up9apY9lTt2q+MnMoNKCe+VNhY33GVWMdR1uOSnYgYdoJMmnkgcJNv7g8EkI
JoVxSwbfJ/PmeTAJN7m2ailtppTu3cK7TPio3i9mK8hiyzTeHLjHR6dEU+0i8zKm
eoPoocQE9HWuFoJ6Hl0qRwVmynaaaqLhNq8bMG2+RKypsLbn87jOHfbaZRCmaoyY
FwFrpB0O9Gu00QHR94xoaublqDQynUC+Ts2LU1RqVFZqg9R8gh0O1Y0+KlUTLSVV
aBFn3DZMqq6V9fkdshR7san5nRisxL6JlvgyZIPskmg99/kD6KQ2m8+xitPVVEHv
AJQ13iNICt0ZbNZhFvLF0Thpu4yX+6cZKvjgOGMZMvN1fYrECVkXO2naxhehO+ZV
IXkmfjX4M8drmdiqtg6fPQv/1/o3vqRc6RKRN3nHvXa5QT0SJ8NfUxelhdFWtzFi
HV6oYCrayDkmlux5GYAqv7sMUzCH+zKYR1Yfj5NfMrJjgvdjD9IzwOLyIgfllS46
QD7BQ7fEzxdn2DYuMLz7Ifq8uXxS5V6Z1rtkdC2nV3AqymWz09cEfqymYZq43NFP
RH76QnvQ7sP/z2UulXB2xyOx2Q+UmkRMyiaUsN1wKBUQrSM9JxOuXKBWgtB8wGnm
8/pXWJWdDjVF5Z+PvXkFNvvPzjip+A3j7xD2MrlzgFeu3u7YLQuHDfrH7/XVUvIk
MCappUE2kW7jwX3utVyq+C/jyiIcxyo325iWys/eCLgjoF/JAsCv3WZwNIozKeDJ
Zl7v5KhreRCcIP9H2aMiBgntZ9El+ZqL5NXklqcKtvHQpAqfLyAdCEKBAciOQciv
HhRZ9Wlg0DZSDU3dDFw81XUUo2oowfL1VLBA+Q+FsavvuVvD8Z60/KN92oRuGoRG
MM31aRBDgvqmma5y3CoLaSQCxH3MyY8TwrePVr5yzAs9jKBXiZLvk0rUXH+kzc0r
ibQWVIZtQWRIpmENrG/8cuyXGSESYGEvMpTNXk42jcb8A4OLArDobcwryHGB1bfY
Rp3McMDlRv8iti1dUuBtDQ6aNhTifpPnYUNBxFYxdVS5hwlWyOy5B2vAJqHi6sEL
6hADGO2N6OfEpgeknDHihXKsJXTDczTqxAryQmJeFDIHMEYdFquHVmouVLl+B1YA
nVJbJWxO3B8irAGgEZwS0F92rwBBzfqOKGaigiZoAreHsMAocL6OZwMWjpjQ4y83
jXbOoLkWM0/VfPdQj8ujckMgyBHBM94qgCFbP1k+tFKs24GHGGw/fTUfd1w+nkB5
M5ENlrZ9X9ixpuxt/OoIFVaQJeZ4gwBm9vTOk4IUWsDXIO4/fxnYkZUA0luQ1U1t
vc7SO8mBijh824Wt9fBdhVoDyUrSO2FyB7BzobZHqSEtKLcE4S3qZ5ZHsag02Ujz
FrVNOXnJUkfpriAkb4HVs2F7aNSN9cA/PjFiKh8radCSkNuUQF4ananknN0Zb21y
qyKJ0Wl39Xpyv7ftUThP8qyuvab0q196W/TRdugCm3QcsThMw5vWaatnSIUOFElG
zEzA7bmsEpwmcl7sLefHDECqtWY5KjU4Pb6nQ9S8SXeeLv8GoB1FDQITGkHI66DB
0cYGmjSKnTxlj3uVf+ZI7E4Q+6x2aIhH5Z0//glZc0I4+dd8sPae7D3RNNyOkSz5
qAdHOjndQrmmPwraFMYDAmymGHdSYRyXg1tPJoXwVNK9esnGB53ppgRS0FNtQu5D
dGP0Ed2zj/rmYKXQ4wlxEOhbUKNozQNSBUQgqv1QUwSwAAwDIS57rqpzxGO7DjNN
Gu0rKj50IJZjtQ3bPW9JjckSVs4h/QLJjpbhxubcal1Dsmd3VJVJcYIb5cPeiE7X
5laEGhyEwhBT+7gLNOypuq4VtftAXH1IfLO+1BEYo7Txb8Rrp2+9yo8OULDiVojt
DXKsWHzX1UTypJwTVIbvTbCn1Osk5s3Ee0LyIoyN+mKlujXEJ6Rxn0/cq5Op/pMm
97suPoyTj/DO7yRT5tEEKuPDXm048bkWhAtg3Dg07dM3JplE95GKek953XWapbHu
eRHRJPdhx+/jAVgKIPfWoiicSO9yGEyKMo+VQDXjnR/4HFgtilLxPJDZq7uHPMJN
flniPzG0SuEy8uWry8Rk9alNYlotowXP7OwM2mjb9Ngxj17RDRksvE3bX/Ioa9OG
TVYACvMw2x/ZAi0s7wn4XjzheBwDKyaHrC1s+Cs8GyqoS1vZCqka09HcA7yJ8vXp
OXgTjKIluWwFLozguJbs5XmnC/it2LUcxumvNKplLMlQClGTFgyODVoAc3JqxuOw
2LlixKsUZiRlZL8lThqthEtUxxbrruaLJRaUsW4d1nOGRsGm/FTq62CJRexo9CXT
5rjGb1jXxFgJLM6M9D+8BBLyZWwdmt84rcpNwsS/3UEDgjOX35Fyaf8Q9yjqR4/K
RZEzBv8DhBEFDZUH8TFgREW5v38SyeJU9n/jGpwELJXUTjdmP5lltWh5cScNionV
bI20hO0VV79TG1Z1WzF+QKqzqzbXVbJYRLV+T6wqMk0WlhGDUFKLS3ffr/KnIV5s
8+eWWVEdJrr7XsOY3pxtMxbQXbL7VlrfcTmSwqJop7Y7PI7cXP0v812NG+zI44Du
abvePUeSjfbpnE2QL8GjwM4Nzwb0HTCyNKZtplWiXYPvJi/LYqTuAsCxM+KCClMr
+8qyijXLBMzgFC8Zz8fPxaznODVbInz2ug+bJtugM7ibobtMvZrJDvKROqMOQu12
rQiI+R8a4pRk1LD/w4bsv2b9H6RvumTokovi7mPYjVc4iSyq66MkOpEUB7RrcMEp
6NPdKEr4YOMNoroWHJ6egtqOgAQ39HKLz8s+ovZWHYrSPilTHBktKM7AMsWfxBGJ
7NGXm4qxJ7BE0Gvg2ilLQQDDWW8qwsVu+mvoLpDFQUtY2d3o43GJqdyc7fEA2VBG
nIfgdfXuMV5Uhav4d5S0wnQvIYfm1BTPGPfw+t8V6zGBHmUlzwMXCkCQv1YVbP5w
ooy1TMT0cMgRQQlNqww/N8QQDJTQvvf7jy4srVnJaEaBuPP0SYoMmia8oIE4uiho
sVHkrfr/rlCzd9+YiJrF/VoMfpikggeXzjijLTPq7nljlzqwwlj1ni9g8IM8x3eu
0IwPDKH3rurWHBpGZm2IroguAcuNgnAZ4diE90KMa4Uf5gSzPsuu1SkC0g8Tsn4t
F51gw9MTfW+VVe4ch8fOJdYzVCaFA8g8prbR0c4HUG83SZ21Useoz4c6o0S1AX5u
/bRO1UVEZkGfm405Y3eeAmRtiHjNg37DSdvWB98zhL0gDEkz+XB/afMujhNkoVA7
F6Vt0FMdgDgIIqSSEpTZUejnVUVQnzykdut26l+L7pNh9LppbRYL2hFZ++ZMRlLu
BnAcikiqij6npOVEr0crEnEsp7TGNNcRsNu/J6WKJJaC3UrUenx8uHxEp9OWQetC
29yD9l/u/SSqSYIeVBzbgvH5NeHEaZbwRoec7oD8FSUKEv7Ic3itOHMEd6+s8dk4
lem8wqA/g8TGGTf1pyTIy6M/4yqHcCo3V9bbMwSUOJSDLKbY11rYmux2A68zdEl0
SAuw9n46lf2Y0zLLFNlUaRfU+r94+7qrE/sGZklpm6Dbm2tk56PZFYwtYrjU0128
e1Jn2p+1u4SdB9UIgCepZLZe+CS9ANnWXk78CJmCc0BqRc5DO0hpxwFw40dqV0h7
0qWMyY4KG3XG1e6EjKHCDLEdElK5v2ZnUJUwALUWr1CZF36YA11G/2fYurjOPKis
lZGyboFS+Z2Pp9xCl6DFbvQKkeoson+CsCRH7X5GhMI4cKa4sT/wQCb3YhMxxgor
EaNfclLPlOP40l0KdAECQdRixVdiNuFDgo+9IcjMkKUfvV7Ct6noyf5u2rXOEjqp
EBE1u0H/KUxhhLY5ZWD61sVB7JE1r8fmjgHhFMIWPj78VmL7GE6tVPzH2sSN6gSI
uh3aMR5XWz7dYqe2wYFSKOaC05bll/M+h63Jwut7jSMDbwFiMlbX3Kr/FZla/qA+
wylREBtyIjihwB7E2lMUVpbT33OwUadgAySaGhZkItuV2SETl8JrswuhdxyrugLp
zGiZFUt+a2kMNFPi+OFOZ2TAJtJLq8ptejRh01e+q6tcCGY2CdGv2hPX2n2hFXNV
HG0DfE1gfMSecC+PY2N7xXcp986RLTVejUcSDdaYc/Ob+be7284Qg+7J/TKq8OLF
qFYWCeexPdV9RSBYeGdcLWPTFJlYOwu/1B2Rid1dKZ4oIPKEFVwhhdj5R+ZQNNKr
FE8l5W+FhCMUdSw28pxcwF3gIfIlMeRx8hDSHzrsy8Kd6tb5AUq8QiNk38/49mYB
bsqc/ImmAqNe8Z9yvvd3YDJuE19XRKb9eieC3yG+CMGvD52ZrB2D4nJEy6pPhK5z
CZsbQRSsAOHFrG3H+Sctg+CqsurG1nj7pI7cG69C9tyTTRdzK4nEPmSE782Kaxa7
29T8HRgsJaSC5WOMBJXdhKKrhb28aLo02TkI8rGdfS/LIaCZFEQ4mqXfWscJHRYC
Ixkz4ibozoWLEiMUEdx4yxCSX68L0rePMRhfn6M46PzmI71JEcqMvr6dJBNgq7AO
RPAiFZuo9LLvq1WkTv8jzGduQqmjo55e46gtd8LO8XXpoOrWBEOzb3LmZCxDFhnd
R5wHAIvrDU4yKErv3e1hGs1OT7/x0t8qjJ7smB0JLluOhKyca70DYfmuxRz0SYfJ
+jTeC1y2Jd4NfxnMuGFQCEvIcVFjSZjRPbE5TV+cDUyVgh6M5qjMOD7XX35ohdPJ
dlrZ0SpR5bO4+CmtbHsNw1Yzh0oZGVPlo30oaxf1/vbyV1mPSvyNX6hANrFVYfuE
D6uQ6nFDZcjF40lmGmI92mOpo31U/LoPdgxH+n/LmOpkRgiHCxUoZdnT0LP5uk8N
cXMDe4nelwTFRWxBIIYozgob/poDsi+aY2rrKZdba2Ib2Hg9tORbaNOjMIqNHtn1
xojgixSVrUsBCeA9XbyuqPswv0TnVYILtmSgcAYb5xQXA76PqAVfyhZmugEUUPp4
kXFblYNC8AEq5fsC6KLSdyN9oMi+YGxtZBizye8R//Xle6Paq0Q7/JFbjO/0XGdU
74URnpar7LjP2CgMeTUdF6Ap5H2N5pqOZKE0+JTa4hS2hgVjmFAL5F+vdHqf7ieg
zcggl69SlPbqnrLutLtsEwY7OeBM+CjEQyGOLCjexyh8y5ImuHX85i5xn6074otb
HCOcX0LN+UuxqV7iANB4lPbPwRWZlfiH6R2UxffPTRz+G8x+zbHkJJFO3CaYvhn4
eMW37jFuFPRuTTgqjmZl5J3er9srQDHiaBTA1uejvcSmfeStCKnrgLxoQw7D/C2w
gUcs4BLWs5/rcAoBJsfvojE+ftL4Y99oQwmmwMyL+8PqowxcfnpYOOWIhvhUwt2T
thzVy8O1uguSmqhJbKiY6oVEzxOiZfHwcsV8ZuszstNw8ExVfuKqdRbIf3zwAWpP
3kJ+aOwEMTiyV0m5YhSCP6Vf/cJIMRV36ZPPgWQhU6ta5PDmc77MFtE3Z5P+TZyJ
9JL7Tn3mf+1WDrxv7IPDyOdAuFYz72zyoOh25iGj8MMhOFAIFHu6t6ymr24VVJA6
Js8MMdmkjjRZyEAMu74Fae2swrtZtPVDHxHJ8YBSetyIeJtDMpHulHujmoB43gyF
BwcJYnK9JsVvtadHaH1BQJTa6CSwH6dVll64ujohFq548svzq4IywNcA6RCQN7oj
oWXku1+Tvp8scFizX+dMC8vdvmXW3mgG9CHTI0tAGis08spV9qupqJFfH73Xi3lj
ITjRVncYyWcOCxKc+VnrT9QNc8crCNq5Es0PupILjRPQtozysT4CmLDl/eaGKPuo
UIHVEZ4upyMVtxWlsKtS0NTkrRTIFdAfhdTy3/4T57uCv6A60UU3jtL5vYJvnzxR
XrNRE7ydjgVD0h2h8UGSO0WHmod/x95o7rcntHP2JgnLlSXX6/oh1FOPsy8oQwgG
sUwKjM7JrP5ez8I7tIBw49BzKKT50ZdBGTbItHypni9ovtofkJJPnDUD7D/oC744
uWr35Stm1GC1/WEEP9H8EB8J5AvVM4RR9IX6ComVMzD5RKxHhVo2YC10xTMNjx2T
rzX33eSJYY7H/IBcGe12vi4T3C/gS70X3pJ2eeH5Fo1N4SLgYhX0WOywOvsQcFDI
33uytghGgssS71XJGKJiRiL7POAZdakR+ICovPljElNJPcmmfG6vJ9Z8O8Vih4GB
xbBnqoFSRr/XPQ8ZfcnE9NbsB4oqHwU20MckMI3GwDU3aXNyxZHYV/a5p633hU8J
B14lhmfLnDf7rXWWwoZdZR3pNyol55VrfGMNYodNy7MKe5IWjq8j1Xqdx+Dtp+0C
2XCx8hufYloqeNMFw2czKx2Cw8/O+CL4bp/zy6ST4sXGM0Z31OJ2w8/xBuziAwu3
MWr6T1zJltcyMLZfnRUXqwhT2mzphPblPde62BhMfypfOcOQmMlsfIj0EQy3S863
82N2p3SLU6YGL5GL1sqeX35JrmLoEUx30RrtQAX2TEz4lmZk3mvCNFJn325dVUTX
RcDEuVxxlnHiI9i4x7/Qz5LC60XxVtaYiOayQKQkxqgDNcEOhWWUU7xWuFb7Fq7B
ESqnLWqd6ospN5Zo2Uj98chrxQvzj0P9K68i4tgO2ypBVzIDVC6ZjyQq6IwiDR9d
AtqUY7mAtO/8hisDcOZj4tBE96zX49N1Ss4/71r6LUtPfdkFY2xUiZpdkiRqAahw
hT4SgVBy42kv9Tu9Gb8WqNJxmTN1mDETst/rp5S0T7LI6E0UlWx/yrKsj8Nh2zT2
P/swrcX8osLnFot5gHQnCJHi3NaCxZRdMWI0ew933fBQrHl2vXg0S/E5XWy7H6yZ
lgakz+bGJoWm5oxl7TqT3e+Db0Ez1Da4cT/NAKR/v2hJl2J/mzdvnrttBwQA2lr+
yS/KuFN1f/BWgtoVGcAtA4Vbt5jt1fGsKPv4ybBXzcm6iAecx5URSWCtXtT4wIcP
HshHzfSaTYHIMS1nL9oAfTZMcoHqo9vggW1lQW+8kXEVuuLO2LuQDLuGNMkLRtfT
SrSrULfd8quH7swVM8Q2eIzOeB1+x93Sbd0JIttGooYwr5lwA5LckipFNMssmzqZ
v+gt7cQnmry5RnXhRdqMmgF1CLWV3Zk0szcmXbKWeempI0M9Ql18hFvAPQ/sRmKb
u9uyF9w8Cf20FKVKu9OpoGI3JPvO+OGMVmzIPJIGU8AO6qYktn0wZSZhSKflTeU7
XJsiQu5NbvpVTU50E7oc+9MAPRRE+6ARSgcZyDzubd7UkmZ60AJQF/z3In31c1j4
Ax4bFKvrRwKIRxoSPDa7HAM4MaEeUP8gWkDk3ltn46wvTZ95+XQnHSQc8HPRQ2yB
8PjYd1MrAV3gCBJK4CXMuWr6R+VuZhfs8g3ZSB4xyX4jB5uhH+qfVTHSzqQ6I/vB
RbMVZWfkRMqnR6LrOOaOxlfo0R8ZZE+BdI8D7I+neQHzJDd4Wfq4FMRIhwkmtYmZ
or4jdxXI0C6BAnRcUc63Xxt9G5XmKItF9xHioBZGZVMppanUwtYAP4RKdl67Ykz1
WQJENhS+wGZd6ZImbtCRq5VvN7KG3L6z+5FR9BXpLx/EnHB2lBL6ReUUPR+0jGyt
EXPlWCk2KSKNM7bRldHQggwI4tZoe3ZKclMDJQGo4APGq2n7yT/vRVhQFBZP1589
EyvyP2VSopFPEG2J3QiziABhMwi10NN5A98HB9UyIGK9JrTcOG7KTfRCrjAOnLo6
WPv0Oa/GUfJQnKpnv69o1EL6uULrA0aRJy8qdRIFidjjkIot3bOPDp6QvBzefB5d
+mQGp9SpfrVd9D2OnNpcb+rMFkQYjxk5FBp1/XECKhCSzZZJkeBLsmXoAR50O/zD
pSTNCC3bLFUPBSOgUtEeZQTnP4P2QOBKpX2WAwlm3PVJ5/WM/4QUM0vh2HQwtBW0
FSBt/6NppRp27P8e1V2oOoKwXv6NNA+LKnmS7KhOdmGc5S4ihjqNjLyHb2GCWX9D
Mb8vLxfqD0O+8fKWyp+pOusmr0+9I6EeRuviHHOPS91vpd2FT5DCNUQ4JQ52Hys2
jGkw6i+lS+QX/c5rCH9mMD2mFnyC07+e6itMzQ8FaY2/3fBkJQ2UM7sBFGrbSWnt
g3GLnoJVJwAq/GJqYHlZUnughGpYmgk9tjBBzN2UybMOJ4lHSKERhmXaQZDhpB/j
O6oRJUDj4xprj7sdUhhLKWiFl62aSBCFOpke2roCIaeCuXhIsUbRdvFfxOrXqf2f
JrZ1MR843FYowCJ/+/RaHrlFoEhz8UoWiktE/IDpL2kPGUFVDO8A+ummLYW1ZxLl
l1JnEhSX3iCsUAwmerxhnVYW+dhWYshRe2sjTIN1+eR/j9M+UbQECJx5IlzAfZtA
11aTuwyGCLo+A5e10sSyoRr4oKFBYmrGdWTqKRshkEzIbpUUC6U53VfCbVfaDPku
Ze5LsrD9SkmgZ0zxe9d9GDl0LY5QFtMfn0eyD3rKLaF63MHaZyQEpuaU2gDrcj2H
FQdrrHzDRGv7NMbrTFO2vrlTDiIkwXWUs9djSHCFSAYQox6alCIGgC5o5uYSyIZA
VKdXWy9YHg1R9HzBUGmmtVekkVzSckZ5V7rlWk2xRYtSga+ne47ffw90fWxOCScM
DQcO9MldA1CQtyKkVqTBC+ARjpsmvlzzzPSp5HLvauRnkoygQHoagWQq/x4rxXsQ
siRFL/vTmA/UkWO87Pz8oQBUGOmsCb0pjZnFhBERhanL25n+UhmhL1niQ3GvIj7+
DkAG1lx9RUbAVdck8ndzT6GTFAApvDJld1Hfx3XP3jFLgE0gXXH2Wpdg/whBFv4J
4wQloinwLgI+M8AcGwk0kxSSGazHdWvsqINbyBGzo2TwYrdCIHSvC9/kYYDtw0qK
YDhm1mTFmGWfEZo/qos1NrUBUS/v7LGa4DUz21tKgvfppQgUe/HNYdWN6M6RZjnU
fT/IPAtSUy/DTOsy4H9Zv/D3Y2bajJgH9Iq8ucN/9+b2F6fknMk+EZvChYBgYt5+
TqsN8hBXe6WYf3ZBPGXdqiDFaHl3cMjN08eHN00wgGnIYpuOxvf/JhDHBIdFWPy6
5AhM7fsV1oX4JAFzvICQIbyfmCJND6y+VVpGhN6EModI1cvjbc/2plZ2sJjpuuTl
wkQA4Krxw9yKEBXfnM4AeCF4ks5lq2Rli+GhB3FV828/nL6SkmGxf+LnoQElhE9B
t+XkRCe8a5/ZSuO/0wnUp6YKp2GjXM55P5wBTLSFrVXKs3G2SpYLhAp8WQ4ayNMN
WpFD2CynYufsTu9fdmW6AVAI9Mx/uxpAeDx0hP9voME07f3OQUBU7Fl6ikkFBQ8C
a/4DKNtuaK9CYa0ynizmBVvb/rbk/XKTX729S7vQ1cdGwxOEFdvuSPd5StVdPCEM
kF5mGW7rHHHv0DzYKY+LWqJ9YVdDSBVuB4NQo0WzI2vZ8atavgCZKYWOU3to4rvr
QM8rTv1Tbxxu2fyy5pWcF8gKDxXE2WRdcqGMV0T1rBjcb5H+SPHuXA21CcfcBoAL
n8UEW3ab38XxStVhzz6T9E2wRdLroDMs7M7/qxquceihXUukjWJZxs0wERmNopGa
5LyPKH9P0eHE4FOMetQg45n4Ca/ClaJR5lrQHd7H0mF4yhV8EaLxVCguIo1cMXTC
WCIILY3WMdtUPZy6OzPDFAa3EjBqoDRIowtdjNzDZNSIf9TZJTAvr2QSMyQOkIzc
XW6ke4OYa+oPjjxWhValOOqLfQlnWfT1s0LhphHJTR7v7FsQuqnRsgRktFGi+J71
Pv/1Qle9k6ts/EfKSGV9tw2b8830hvJ4AccgTYgiL6SgrhkBaCINekqoMP683ttb
adR1BAGiPCz1uUUmdZ3lhnMp/5Q6Uk9FYi9VeziNRVBZVfBV7oWKxxRP34YZoRku
ZLfMRSapdgn4l+LaXm6liX4erXBjJvH5v/sag5jFvFnBrqvzYXUaQUok4C7j2Xzr
Y0aa2K8VJ/NyuJabDnuPsDJDZ6rcGszW+Yyf1s5E1wE5L2DELAFA4G8ur+gAz2NJ
ytnsaq6yNGGkmcbxKyhmariqpnTSegNQrWjhibXYDrbXhhE5Li25WdBrODeLlmXP
SaL0I5T8oIQ1sWkA0f95jaweAa6VORRHV9377IpQJqbT3shlFCjUYE6aQPftYz8p
SCUA5JzMggjnbmT1sEa51EI7jFWH+3l/aeluOs/VILK8KoOnFtJRJGjJFgPqVDqW
9FS9zs4emRzvSb2PqsiAsqwEA3WpYy6gaeK/jaqyTRQZy/uDPjGnXkiXDQZ1x418
w9KZ5fatQ4FK0m/IF65TDXIGWhxuJQFuD5ftiL+p9xgCKyWsfSt2G0hyIpPXPtQJ
Bekbwp1Al+pN/unxg6Cg5vfRcyuekow9VZxuAf5EprZ0Vitq+g2EvJ7zawJFfYLJ
ybHLrOpJ6jcSez6nkZETEPgaEIWBGufe0A7z+qGJFZbAirgi0+VROGgwkltbNSsK
Gf4QAdFsyAc/pl+6e+nFAyD1Em1J3WcNwA5dnDNng1OTzJnXcYHsOP/StfN/X3Z3
SyIuQiQvuvpxTQ2gILT3fW1bcnJtbyiuNTs4qeVUjkfjysdxq6AvBFWww1OxL7io
jnZbXrCYczgfU5bvJxk1uQY7PuhVLWvgHIvxuXAG/ShsDFVmiBuc6PcSx9tsv1zm
/LUJQKjW+rJ5BMhmbFjclCpjVZQ3ZAhZCy310oHnK/2Crn+aXs1TV/+NyronobsH
nDoiescamljnNnl/fL2lk4JwjIFDhK754kPgh3H61R6XzZ6m9hQ9cSNIRT5G5Qjb
Z3Hea7muXPDGwi+wzDf3u/8uLPhCTzISb0c2h2uSBNYh9xT5J5i+xmmWCJVYQxnm
24k7GEOwZoAXm6x0pCJRlpreG5YkRxj2vVAN+mx1/xpAREKAB7y7MRswGlYt239h
Y2g3KBzxwmDXScFZh0GfvAkQXDrm0zNM6+xh7r2ulmCOTC8Y5Y6BnwZme6qtVgGM
dok5txC7D6+Vej61xXWRix9TYqxN5+FuEA99pWdg1JSukX3ptvmi2KoDsQpuvLP0
LoxybXty2RN1VJ8bCo0Oy/6pM1U1b+atjmUe5BYjFQT4NMHw4cJ47kc56GzCLqlV
YGVRRveAxMhJ5gi6BEC9qPKo/5qjoL1QLlk4w8fXnFERzheS6Bo1o8Q817OfHkkn
eB89hO+M1JWYZJZvN/W9WmmWYl+SPGGdHaXGiGYOMLOWxfjNT6f1rXN1F1nQMpe2
acCs3z3dqdo6f0AI9n98uR+gaeC3+2iQIFedo4MHnqLwCMhmWYpAlmqd1nYbpF2D
B3+1ol9qOKkW8cvucYuHCzzGU+xzcjoCxE3TXJS5y5mbb2xa0wDRBy6a7f1zMfIU
9FY+TuN5MwBhYh2SwrUjEfBJF3UtTc4MdF7rogDceK/HLP6e0WuGzYyRjrz/9248
ZqMJKNn1IzFjX0NSOf5COAdDhkp58VkbQZWhsehLwyWQrcerTBhk8WTZTyz2nLje
jYfwOyZjLx1FluSA86qxOzRXb3SwP2zVRednzD9cNVPiMyXjFm5yBhu5raNgWLT/
CwTeYnmDLPgj0tU9b/MduME8vI69S0qo8C8SdlbdO8Ivk58NxXkIGAJLwHX4I/nZ
1U2gnyuHA/S0v1bE5etrO8XzXN6gRlufom7hqrr862B9izbOTZOjx+I8/m1mu8ef
6omzqgkGQbmQPdfeAZ1U0ri3VyiyJ7jexw8DaROvMzojQi3+7vlroYcK3zE/5Tii
pbYn7FZuPQ2GwLJ+GSSpi9OfpxL+SkvBUMLWiBoL4qpfA2aMpvnDa+btq1G8z9Au
nxvgyUDxrcSc2TWCn+1zzAgBV1I1sd5mMS1nvBycB4GHXs635wBd/XtDgNyqmnyr
Dl+/xO112LbQj0jRxMkY0ZIt3jnEUBU9sMutWYbC7PK6iy0rRmhLlGnRU1ttwo/w
uTAg+4zkiEODeQZ5pXYtyHCpsTzodupnX8f6hOlcQau4T3ad2AEq1Bo2xeDJKD4/
Dm/C+D513DGtAm2gZqdK9K2VelZqZh0I5ShNfJOaICtuPX4qV4T68XSMo8Rf+fQP
h6Il5dog3ZRbNTj051cWfA0+mFBH9lVkrz/g+bZnC1OR6z0NW1lOKHQAUSPZMCKW
AY4CZyDHsBtp6mpezweUwWepd2/xS0PHf2w28VXsb8vAAO81fehclDwRzbj8m7kn
4CsUnAVtd/VuvPCq/ZT7428VlcUqAnfAjlgsVVc95rS61r/p5Pey8OKxtEDvfM2u
GDMh9NVWUuGo5wlOzz5BSz7DZE5MVYgFGvl2r4/Koctv1m5DE69MJx6wH483uV0u
NhdqBRk/eoQAjFBFGmJ6Ky7cApP+Ij/yeYGmhChv+q0vtThxSQLPq87bVguMlyal
ODpbJZaz51L+pk8us66U+KYKLg22ums8ZJ5+Ma2sTJ/KNeSszlNkyHRnmPQpVMV0
jAk353LzDeJco/hDsQ83q3fesUHTwUZYWtEV02pUkTIqXedoP+MZ35G3Xpd1Vjic
DcXZyCTSQjPFZcSmB9h7hIl+e/Vlg1eBnuAI4v3Z/r0X2GVizKyqz2O+OssXXAXa
6DTvdOw1H+vCkcD2LP+IJKhK0FCJqa1fxyEjW06a836PyoUFkgYcc2hmoYwMcf9w
eFIARgvGQ9TpkIcEtnhnDBlQZ/2Frl+HaDMWFlaMqTGX6QRSyH9PpgXTC3p4I8ii
1ukl73UXUp9hVA0QVtG/4wu7hCg8MWxNzZvmVbXs37eeD6iAc8/RhnQn4yj2vzT7
Dm3NZtYr2wEWjIbAyTlNyg/FUMUGTG4bUIMkT0Zoi0d/Eb2N8V2RaAGjxS4u5SqQ
1QFlPXOgbnqf8R8MJDVRDsgGrR6wHa1ET9WWb+x0L88YvoD5dLecmkVqNFZVCg0o
bmIkmmfn8HXHxWn5Awo9TaI8QcPNsLfWsEP4gKERs9J01j2ooPiU4LA5SotK9575
UosI9CCQaWiLxFxjlmZMeagyJdPyzgpSYqvPYG/q37ksXzcM9DsNrqy2Lk53x4NK
oyoQRF5RaRmT3vCaP5GP87VmjuZwVb9EIJCH+4Xd0U19PvIEmKAhjdnm7pRxxlm4
3R/M9eZDMymJwiKKNNWnliNxaM4TdR0kEYxjDhfuRYa2ATBKpr6aIjWCPRgf7u81
Z5Je8Z8ExFaa1cFh5z1OztWxRqJO7Ge6kszCjMH1YMRXE3P6GH2qZfzBPgxRYe6/
Kq0dnwQXC5lmWHJ+JqxjLvAXEL+aEQwMv+9F+OQzya44avlilCWgJMn8w9GIw+/9
9+ExaVNypkQ7YjZbxgVZ4WqsxxT6rqxFZaCNEmtWbLemDLgLjucfEfqVo9237AvM
hCFgNOaCvXLJowpsDQNaK/qdM3MtBIDXef63HybgrkUU7F9n1sq/O5RdmV+IwfMp
jCc/1ZwW6eT//uRVqGG9QxciElymLDnOdYVAuq6oIYYEgaMpb+/7fjO0U7aUMSI2
j7/JV0hV4TES0F9Ql/mZ2T8+nsSDhaKlyC11Wj0HM7oO2eIWdbOCQUMuDK+gsoWM
q/q+aZr3Dbk3RjeHGCk/heeyFEfNHcP47NJHLx78XhqUBZutspLuxe5PNif/I/Vd
XGuzvO8u8H58n82G2MJ32zQo9YnQWW7E0AXOpLzImuQMXJ7VduH2ERDzWPFQlNWo
ecQ4wBFI8sa4708OjtPOBTFSdNNvJ2zzJ1SZkJ0Z4XukSDq7JocA521Px0DXsESF
qSwQR9MHoWU7Fn7hKEAA7gIchUOVJ+hTH8i4kcLLUpXVQktgP1/KsyMlXlVTpNTC
XtlsGPfYXSW7WrPtZIF91gUQlx7S5qWfPNylJwRA03HtZbTraQLl81PQvT1G/M8j
JE2fkkwJqzRvMEEmStOm1AJykjFn5AeF9rCKsa16APharUiEdrQsxNR3RDvSeRI+
hBoL2dff7ZzSOIfjJll0r7h36Ab6s+nzohOarsoZzxfxFgk9fwTF90lVGYnFJUb1
BnTvKZ+OqKUlaJL1r/vjnsbd8LtSmZr9fvKhuQDL1Bw0SRlPrpCcul4PBPI1TGl7
uyUs+amQ03F9RnuWdDyHan7kBYJ7ouhOV7Pxd8bGccB4FK8jxvJfopnfxghMSvwW
HEuI1XYyL0Imi72HWJpjpXgrQn0enW3xkCRp4xqNW7xxUT7U6zNcQ6Ugpt9iZXtI
fjaGd6YRG8uT/ngtY+K6jXVMwijFN+PQyTFbi81CGdHrzUP/Ij/d0KeDGrAE+8aD
FpkNzslhTKenrWlByee42aCGoRQPjx0RMphAXaArBljNYS7kEfGBUQ/erVhzvLNr
Zb0YUyBk1DRHAOJ6Gsq9mx2eFCwPLHsGgd3rEEwq2xc4a02OFFJ/Vor8Dq9QrGk6
Y87R7iZB25WIx6QysbF/jm99/gxKtCQTZ1hw+kWR5Eqddd4OhYACfhU+LKoBi3W8
31jJODzQtsU+UfoYXrWR2dzg8FbFtn04QrlhQb7LBdwbW9mCBj7cfcBIu98hf/X7
LVqk3HNwfIXyZb0I90yORV2f4PLxu1HM+2jAe9VGWjC2BwA2rFVHOMvDyMdZgDBZ
hpCcZi7Si65UulZp7ee/b0nTWgw1Zzidh0eEVKa/0j213aY224kI5IpCHXlTnGYd
CYzL2YfO92F+uk6JhYjeczxhOf1vMJUCe0PDLWr+ps6/bb2rHh/KG7m9GRU9TFKs
x7yivhT/PTmnsc8E2JBWqYzXfVLGDeqtgVnZy0eFRxIHlZF/EP5mVj6cyhsuuZpI
oCjrDBohmYoqCPq9O8ZCZIlVxBEv8YLv+qFIjE+ryPIkbNv0n1JYFaMFgXl2ZySL
zBgfmi3Or2BBUSc60Ht/JB3ItY7DA116RLU9m8RjZ13PP1pvtT4bow0zbXS1fAxY
sEIp2oRs+UC36NL1gAhGQBhHkhq3EZ3lO3ZQXV4dXjgesJ0t1PkkTWm6vo3K8IQ1
XTcsJ0OnYMOC6JF/RQGYDJ92QLBftDTBIZkRyRtGvWwyVf8I+vyrhCmGFc1vIbcj
UNN8OcnffJ3MLydR3zXEA7zYzpTPAaTd8oibvKlPOfRunCP/8EAT/y6DhnBcakKB
NLbXusl8KBxZqsw0nJCmJvTk6hW/k5Izo8XNBob6ZL5Rd72/QA/g41hzDDjlYCLg
3ZXuCnjmuThcJ1ErVuarXSJObamErpirSpl08JnZSgkPgT/ppEiJEjfJwFizhDR8
g1LZsm71e71bgz6E/CzvgjbZupW6UzXQgOWhFIv9oHvP+dqserpRx2/EQpoybfnU
Y2qB9bvYAzsAgeWIn4PC4kPjK5VgNs98+bx0U4tk+gG4XpYqpkkmCYYq7O+ngpOE
yecmgX9nSOTuwksZ5P4s4joCdf1edUUCTH4DEw/ll7wM0m/ktJIpm1zRgmwINlZX
mOSWgbDWdTloIlnDjdfHFFjPxO+oi1ycszzdLVNFKlNnPi1V1I6x8Cyp2gEsy3DJ
RUKFYjif8GSWd3AoX/rA/iJV2UB55Y+I24jeUKTOmji0XSQx8LittMNXEuI1mixb
I0mvpVs4bXsQGZAlI0Gcb2+736HesvVNoRSv+CfIP5Rr5QbRWrzuKVjeWQOvuM6M
oyTkC3zUX1rmE/kjNpebLYjYOqZlXvG1+/9NGLco+rxUtCGZRuY6f3WtHtbyXO2r
/GYoP6/nSSSRn4ksx9/VsJHigNFScDmD35Poq+VkpBYqwUJ8iS66rRXTpqdu3Byw
dTn/u6VACwuwgtjcafI+9AtToNF722zUbbyWLDOX9R21fOyssSQY01SGzDmp2GKI
MhCQyqM6STXmpnNVZT+eV1VY4NBHQ7d4ZPecKF6HSs1XJFAsD6kcNGCn/WK4H/gT
CEzLBcG0kdq6hJCqpIBAAPs8hfryb8hQgXn55SnkJOjWKGJtMRdnGYpRi1yXHvwk
27T/1ppSy82rljfNRmFpF8YzKc/XemCnpEfcvd3i7SJlDDCwQuEH7KmxTkjtYiGy
1rMAhMLzbiQGBw54W1Dw/zIwifZHzS2kzUoC9AEQSv68iHEM02TbL39r912e4N0j
rI/bfyrrPQpG9RzfvCSa+B10K6pNFDYdn2rVC/dz+NXEFAbLEvcXlW8/xNurcTVv
H1MGUhYYAbZED1sOQujL1aYhukJdQHCu6CMEn7punedweWNi+OPgeEyuD6iy1621
QWXHvz7RBdN+YdCXGMTG3elLL6BETBqoEMPTj6kYsAnJ6p351SWdgn/ai7rd5cE7
1iwhDpL5oRQfQ/v3Gh9YYevBOTtNGTc374VZba6WPax9VDx72o29lvD5edHmuuFG
fm2tdHFrt/2sOVakTb4Fk07TxHFiKTCrN6QcSn6gO0itAWPcVW22q9Ds5feT/Cil
Ca457QjF8VzKN21jniz+Vv4vuEVrm+PTO70qdOdPL3xQ+OZQSsuzrlI/9Rb45q3m
AdMgnvmZ+9IMnkl8jVsiFpTVR4lmphWZLmptHgwxbKd5uPpgtk7k0h2mxa544AKm
WJHEsrDNbpkCx9aFjLYB3Z/5tUJOPzindw5wjg+LjIhTx4wtdkh0wrgdp6yLObpz
vsRczZPK3K1U53B7AbtYTt6bIvIUj0NP/6TD91GzRtOd/AGxoLibJQIhWjzUCRai
65aYNZBakfKYf/6chEJ4D9J+p1dyCMsVddpLP6zspGCzcfgVbHzCopJ+SApVEv8g
V4m2FXDdhSInE0ASw7U7ulSXwXSOW7oRS/vRLcJc8cDGXaHC5QidBWsowztEDfw0
XnB713t7N/EUesTmOa3eRaPn+W11n3OFkzENC3h5FifnJoU6dDJ1LQlxzut9Y0g1
kEkM431I1PPthNl1mypqqBrM8YR2/4ODq2nBAsUQ8ghF1+f0VGNHjdhGNa/Jnvhz
lDXpgNNKYtGNOHAkXMMMcJljTJfflCV+ImiMW0m9gX9hNH4RvNNriWoR8cmvWSyP
4RqgiCwoAiW1d/L665U8mg2vH4qJQCVlJwGON8VY7CGEURM39rhFsax5h4b4Llym
QYbK1CcPSbNXcP89ZcVY2jo5HKPim/ypV73okTpESrHiBGMdkX6JxhyDmW5roXgH
wfVfEDrZhKPqKarbwufTde3RaS5k8siWR8xhwuST1ezuhT6fIHs/YTeZfMBfz3V4
10qMmC47ET8isWxbMz33yeUDKCS2IHyAorQOVTPn4qQev417lWkQPIfHvlelnRc+
qd4Azu5zdZKCogJDvMgZiIV4N8C5BdfbTlFREwCzRqRyCUT7rsm1kj5mKijCiukO
4NCybHEIOcr5U5SRqbq0XtK69v8Y1OnXHEzjStZSqwZnVyf4S8XaUa3q8gzoyrtm
B/V8E6AetfASLCmfSktBHsR19iDBW9za3RZcLVPBL6zkdlgqTV4EGTIy2Z/ogD7p
nlzgby+D7OJ0DTHMu6+Pttv5FczzVJG69m/X7oQyQjY2yHSUoAP7i9Mdq2monJzx
I5PhevludCV3bW3KM/3ptmaUOadNQ1nvEA7CUwiQ4CfPskDcS2w53SoIoBWXHzyu
gznqfPEI9jp8N9tigCEZs+R8f3k0oY2jJROWhzN3V9lCrGQvueUc6FvzSm3cY5P7
S+9Gg6IbCxJHB28JvHXMXjauqIKjEFvO3raAJ3DtLbci2f0U8so74jnzxNO9fPtD
fiHsvMm6HNqsI8/9sqbRmbKfjdBOFHczlGfDW3yRwpurv3p3qxlX6gEOzODVHkN6
q8h/EdEU3744qc8Sp94gvK925bF4Lm4DXH7A/a6n5/c5v+aAud0Pe9QCykqTWlCM
Nudh8jfPDhSC0eMbdCLQxxo6qMKO3TChGDsZse+wP1rytsuk/T1Ue9O1RCiXz9aw
K2s6lU0fc6fMEaKtdciCyW+YyzRlF+KH/Q/QKkXauSWDM6vrRd38Qe63avGMG3Ic
O5y05Ll2HG4xkb6GdyDwwkDoY0xmN4oJZ3X1c8uDEoz9DlgbcWl41JoDB1kr0LGW
YvqrvJKXRHtfSDFFK30dMJZDdZSdv6EKPSApEgZLfGGj59DBvzosTGgjXtoez66b
X+X2UZvWgtkgdaqeDSb2KwivadZEVLvNt8/ZY8qNSbOPP/7hnSWwGZayMAszC6m/
a2dE39kgBwlRu/0Nve2J95X4fQ/lB/+rY9M3gwkjbSZgwjadZwSq7elQnyhsZP56
NbjbQGELaaWSsRzgKyntcLLTwmNO+vSvZWD3xlgWIgt/5cVrDcQzkbabprd2MOJ9
WKCaz17bgseUZk/+6B9EdGcNbRdHK5Y9FkRG/RJO1lcRzXaq2beyDQwEwYFprOfc
ZXH20QOZ0ZK925IjPuaZbkcJ7r6rY59DLKAtq9DJvDlAy5wmyVoU2Hka8jzgsRai
fXCpdNeyKIM9fpriAJHDtXPreQePAf6padhYmjS+nh+7/nW8RTGwbIuuyh8LTAzs
UXgadhDePwwnmXyNo/9gkWavHsUqxn5hIQ4chuzNG8+h61LUqrH8whysxwJgiqlG
Yao5RmZHbUQprHlaVQMl00nBetoVf+k/eeazTEAsGBgCxCcG57YjZIl1wxw9Zxye
7yBTAV+LR6Z33UAx/Y6b1V5FZA4FskEbmZR4hbXIwU5mpS1s1mCXRGZpxJXsMi6r
ZpGw0/Lo+JRK/UWXf6f78/nFtwGJPTvkusJcw82ouZnEzBURZAF6jqOxv8R/QIju
7mCgkZLw91lMnhc9aGHKD1Dt8xUg5dxpBYk6/hPGpsIXhdqy98XpiztxlGSvvACN
2bQ5xu/znjyK+KHTYsUXDgYnBfz7Wc0j/aB+kC1fl2gXLwPr91BG7oN/HTjkQlmZ
0i2QHFsXtqoX9FDO48KKenPUpFEQWgjn0L+24xWbYTFJEwJT/GXIRNzeVkTZ8oi/
TBpy/jGPiZa/YsueRJSrTGHJC9WcI+oCRhNbk64pZ9+GOG4HJj7KubfgrpeDLFZ6
YV/9eId1c1RUc9JUO4mUe6G5LYHNM2d8rf16IbO/Io2/ArLVN85eVi2w74xbEvHi
TceYwrvCxjR1QO5lq1ZBc4VNqUAT27grjSu0kNqSTQ0doHr45CGv+dIORgwVLJvG
AvaRDgIm8B7XD4J2ThPAvVEAHKUdh+5zFnd376pOBXOl3/vYZ8IuP0KjlJdKKvaP
lKSqnCw0M+49t5wE7xOWDCKnC757dNZ0sMVvdx2mnDBj1GNEgWY/ycMCiRGqyoqS
pEwH5m/LtOuFtn6XA4cNeCDCXbmbyvG2soY3LYE7NmPwWZET8n3kbOMPxPjsePoM
LYoeLrb4KI/K0iY7rOVKWJnIH56BXxbWb32NsluBquULxL/7ztRcAqY7SsgcSJBq
c9rg2C7+u2y4WP+OBmucQGJ3N8QizmUzvRLiBthe5xMGvV8Qv5yHrg8fLr543KOv
QKzbdLFgfrxxvS+lDOCqeiSahnPFR6MV2oXPgAm/d3n4Ww7Kn751fnS24ih8lUci
xX9zMQpSF0lVlIcDLJbrhDtqMq+RDaVcDhX9MmRnncSero1229QAl/LCAVUjizCV
bYQLcn0raR9XyvfQtj4BFZECC8wUiRNqt7oCF8EX1QXpA9XT/VD4Dtz6zM2ekj5H
u4M77X+O/OujH92n1nh8fUKA5dXf/jTk0sc+HHRsbBHr3uBANRSrFx87e6S0v0R8
gaYL4IBdqq4J+9K+XGLMT+WNPKdm5BjawOZHSMcw/tfX+c+6+YUWO3Y3RS6cNolf
3vDZXlphvNPDqAgP9bTnVe7R2u+jWzLvuEZ4r+JH6LWAxC5skIbfwRK2SMpsLNKP
3L6C1qwTRgPD/vXLG8o6iHgI2b59m5ddwOyLPH+GtImR+7cYyZFMWWzXKFDy3MLC
uj3iIKv+pZlqX4zA5O8xo50HCfpPcoNPWFsDU9uYqJIBMP9uHmvu2PSLvtq4wQ3X
+cGtGo8ZqFIp4G5ZQalc5S42jYbFgqdf/FVCnp0Jx1zQjyuo8522dwVerYXgcNdY
qNd4lYvE1CtTtnz3wUiqXAMw/2Ny85nAedeaamqy4R3WfHf7jqrrf0Yg4kMO9c7V
3jv7NpP1yVxZI125C1Zteb5dfjv3lh0Uxshd6X/N5S+IXiSk1t55vRWphM5K12qB
OsCRo28QSWxETSQTXTgyLvk15VP91paU6bGjmXODjqDf53g06tajWl68/NOAnjSe
UZYaBaOml5axnbE0Sg7qgOifLfyO5XCQ8uv9nAM/AghxiYWeCMmFOqWzSaST0Wbz
vBi85SgjRkpj/W0fMzPI9j/jYMOGakBLyfrcDr2dLjQWnZ8KMogFriIFJAF4w0aX
Od5vRcn5kjo4mScLWJQLLm+k+Ry9GEiBC271jUzzzAt6kG+4nOPbbDx+G/9LJ6Dc
IYqxvPmveJp99umF57smqq2PjgDibCJ3LPXF8j+as3shHMnc/2w7fxwkkahwTCvy
8hINeHrDSNX2X7J2CxS2ETLhl2YaUxzauzqiCsk6caPRcqhPu6gM+PMsU7juVsoj
yIG1qvY68RIYLZLFczvPDfxlvtBzwVzyoOg5CEwQXHEp6jXp0prHmkr2vqiMzRlL
SVV5iZalPWdWsjCMGSti0a5VUSZMxYaOXBwVCXf4eD/Dr6uVtYCrEFte743hlo2J
3qSC9AYyTPaueI8LbuMqDfUUx24EHwYrtsM1crF94n8jP9k27g7oATkmbw4YOlMc
F892/ZZvMfhtvo2RYbJVzitUUyf9NKVCrqpCyAGBTgwA69RU2yAtXUE9c2hf8YYh
zQSjszB/ZF+MFlVvDGihFB1poIgf8VUVSVQg1Ywf6Uzd8uDrNEDF9oTZCilLs2qM
niUHfAwN+XtOUia3SgE3PkcbZ/U4W7qkTuUkWRqnw+gXQCzjPsE/hYXOs0FwEVYS
xCvqkt3AqvmaYe4nGY4aVcNJVF6C/mhhsJxc2r1Ufwk3muds6HykYSGX3c28vNL9
ZxhdgVEXbUNKxV38UmIHA2DLwWyrnZ35ZxXgrd1aneR1rDxDsg8RYNeOAZQRv3fn
cn2r9Lgm17MgbdYtCY06yJ9HvqUN+WRm2moOTBjMQuTfzZOFf5L1mdrC9yjtP7w+
to+Y+5y9K3cNodm5T/X9okgY8T/4qvcEEEgXvOYUnriKu1JV3z7nQxnf+UmE/WEC
kDn4GSVd+dxsMBxGxfoJgNsdVWOYDiWwFno4wSljbo6blJ937OcOnOlnr70bdb1j
rgMHtT6UnjX56UKdALhD/nPA76ZXL9X32pjKXZF2ojUmRcVQL/EI67OGsaPFglun
VoO8Keo0dViqQd13DDBPEKskND99Isi6Qf/5aQvJTuMLdSU9GLX4KO4mPfQURMeu
96qGshFcnTksLiKtEmxwMJ90XHxx5491wLEKX6LUlaKfNXRK/NXy1KWij7Wt7zjN
+EzI2+M0jFARmOBinZyFCiz+PEGW4MjTSlro5zihaqygxfnZeLv9Cek3HAJC5oxR
QzTM38MTuwGStO7/pbvQBHcVyDaYBlWIZvaxcTi+26nL4TLHs7zd201/FysnCPWc
wSrMMstaZVWiHaI9b7pA5Lf8ubvL9ubwiUGr6gaYd0gZCbw8YrfhSg0AE3mc50IT
zjJhUcULUVbtbYQPHbGTyhSGtdkk7F16ljfQzXKQV6J7nwZIKklb1B6qnaW7aOlv
11Kz/wTHjHej5nZz4bT85pzXlzOn8iCJPqRQ2nxwzEuTep1esepnyxB5h15gamMF
F8zl1xJ8em589JgzcBXW3TTLUpY5thHWh0wgvteXSs/ChZ85yGJFDcMMf3z7U7tX
CWkiCd4cq8B+w8zfbxpt4GOac6NUkZL5sYM8ucNdbR0fSQT0B0zHBcvbMf9FpKTf
HE+8hFuuDWreO9sTpxIndvWEFA7sJq0Og3apFuFx9Gg8QZ7gA2b8JWuInqcDiGA4
jgLig8Sw16Z3YRtQJp2RVdVLr4KdrVjR0buK57qoTz370XL3Xo08J54USKi3wT9G
yx8Wg18jbyZcDqP4HtTxdDCXp9zPXE0ppfwQC1DHGdzqVYiGW3hrlCQINOyL2Kjz
P4qBHHtks1lXK5eXS2+q2YGdUMV1VwkZNdHonXNNWn5A86omVyx7BZxSUD0QAew4
LcHem3b45zbqv/Eb7PVe+STj4FQ0TiyXdDrdo1I9s4GNBTP45mUm1jvU4aaqy8Ju
jPGRLS1aTJ/Tp9cqVkaV8EjfkeS5Y40kP7XQSM/e6klAqAqWT0V1D89nWKZeWc6O
lWHk9LlvPNy8p2M/UCZm7xwHp2kNfUGNOJnbYgtNolmjZ4K4EMr7Y25v/z+0qF1N
Ymvs/XaFJqfYq58G6mafvyi5JpBD2Jg4gvLEVV6J8zbMiZ+79MrSeNd+f/RLkfdD
KfLlqiBAWFSmXNhVUN6tCUxjjSXWJM5O/cAd0qaAg/nltlvsyMtXgdM4k0tDokTB
u22pO/g/Kl3knN3LpFNIojP0QJXbUFQKXZrx7Pp30jh3BEcPjiqyv73HrsAEtC5P
XhkcxFDsgPKiXkfI68kNbxVlcO9BMY5bgXzT7KXpvA8sFuRsq5BBz3gCZc1D35Y+
uz2cmLtPagP51OkQddORifwCmtLJiR2r9Ng8OgbvrM1b1B4Tchu2uMBPD1fF+pVy
BKi/a/hvGnV5CcLwaInLb6o8KJiSJJwamuqAgtPdVZX23b/70n7UxabelrG1G64I
KzvUEmirjZ+j5KJ7EbXn635tYDvL0zWaYlsigtXXOm/pPMzcn6SlSB/g445XpJYK
w6wGOi+mcM8UMOnw1npikHkLAsc+gNxDhwI8WT9544TggFk1H6NZd1pgLI0+DJci
3f78KscN9MEZ9OgmDcIiCudGYF8r/4DYSysaU/O89r9dfvPvcLuBU9Pt5ZNec7jg
3X4kv0sUmX9k6zUfPaOP0Lxw0W6miZ5p9HebrkT7o3X/OS/3geqGMuAzgwJuTohE
aJRxeZT22ZfSbl28GzQBlK4QjbXCWCkp+6fgdSlvYO+nd1KpW9kzzmkUkhrbkvfk
Itd9PO9CBXSRQ8dKpUq0NPlhyTRHDqy5qL12zjJXfCQlsk/8dRbS9eqXPvB9us0O
eyBuyLfP8f2mq25sEqGduNFh/qCIDChRt9PQXu3njLztbkbfRXESLF3zWY8To6Kv
KhrmflW3GLa7yz8qW2OdV5REIB2qFNj8nwJbx/2HZeyCGNZkg5ZAivC57ibEPI0H
Sdv6HL20/T7/AogarksZkHnTAQV8ro7CFWUHBnLV76R3u2aIC9e+mMNZFg7L1XGY
EoIsvBb4EvIGiH5EYsWkW8ivFRH7vhPXFzBxtnpCgClZdhnRlfGrcwY5ebAeNmw6
fEZpCTF0Q3QvyVOVWGfmWlIDB4jtdrBb4QqOY1WrOWLV0ZWtxfcDcJCjMu6Dt7xG
Non5ZPoAh/GKyyuWCFT9oCVjxhPzNmCNLPBKTuKeGg2y+IGwIDFc3h5CrEZqEExK
XGFBB32xlb9eliXpgA0Y7LK4QwVUraR/T/vKZsS/OMjKhs+zCbSSDL1/7LsLss6d
lXGUJXykvK51ikgDeCEQnoSmlWhCzbclAWQTDjC/Zc3TpuOc3laIpm+94Q6d/C8J
TRO13D/71/ur/okNF4PxzSFzTKeolwYNHAt33H39eL2A7kUGSGMy8QBAOLERUx2K
zCbYmTdHF2hOnpG1ZO6eoS1IJcWDJVZfsuqLB7nC+j8+9CPIfYHFqSllAnka4VpY
SqzFAyvNiXnEoF5nSHIsBAcaUGBhtZx8BzVhrmQ4Mw9xC0fo2/reo653cUx0VX4g
NSwpDUedEKQzk1492khmxsJfLRsPqLU6ywutdH3ySeN26mgJaD+Q4djJRUVN/iQB
tb9PdVU4ircD6JwKmqokyclzTHPXd1JlLKWnnarZ/Cchc7nIUHo3LJQZdX9XKI1u
v94uz/L78wdrSb8u/WXGteSu9NEqF0PdpN5MLnHnk6j+EJiUNnLuupSnF96i0P3o
JQKz6RLuafSo2yGRHuRY/2iv8z6Vj2tLM/Ztwu+z1TUuziHebTLTKfDnfR9ChCBd
vZH6hUzWycQXg8dqt6Dl/Qb+FIK5pzO8WdHvhVa21Rj70fdPlz3neu0iKpe/ynmW
rch5nqK55DDIkUVY+be0z88tr26VT/qU5KK+k2IgDht+APd1q6/sk2PcBghf3JZr
a6pVQLc7vmY23k5uOVcvdgveLBSNGcGdHoXGqWwMeUKg2MgvL2dKF0w/V2hmzgt8
smf9lvY14UKVZC7sKPkBAHMu7T+FZxmT4a6wY6lZvYhL8HpE005EjIkcYSQZOoKD
yn7AFkgD+/Az0BYKkTNv9k38LEjpmMTECQlsx9OUQ62flcv6FKHi1/k3WToy/FIw
QrFkPglu7FwXhijyBKe6z9PC47hkDoX4SUlzZT3fvyu1JXj3jRzp6GDe71hubcZF
xal/VQ24ohzf/puJn9XbUlMevLoicU3b5s9yW1cY/DNKdyt9Z5fhbmeoLU/cSWiK
qtRvSQoPrh2K1WmmuWc47Ae55F3YCEsmxI7WR7glmJD6jqBPk0V+F83N0jKB+F3s
d1UHXsqDQJ+Y5sFiEVrlk3zo1kXOzzcVQuLmQ9EOiH2CiC3GdBdGZJkux/xh7R1m
lF+Jbb5KWRLKUkjG5gr5UzM/p8ziaeL2pIRY0AW9E242Akw9JEYeHxbjC7fS4Tzo
HjIzQVQdh5TdsKbJrDmtOU/beiZCPGvhO6AKPHu1h7/O3jBDIvsTcMCgfDtYsa/i
umBKwzlN+RInqUNCxUFoAYfs5WzZJwJR40WhCYvdiE9CEh0Id62uneSXkanTYWpS
3kQf3inAX0vGnmmN5tL6AV6qnebg5PPYQUoL8glxH9GxpDnwKnUPqorunYC4Q+to
4fSOn5UHO3X8jJAcecdfLspPG2vVG1f0NSbHkf0ZeW8LgWDGvRZDz3vNDBG3803S
i8qe1WsRQ/+i9reGImG1N8WDgQUOZ8NBwr/qAHllAkm0Tq6ucikDap5PKttjfPSu
laIAhW2usrCLnlehm4fGh8qzosYA2toB8dENUAYWCxVeMQ1EioZrqxCKYyC+fsPd
I656BtSMYS06WFU338y9q7JTCCd8bzBKf0qX7j/NDAOnqGH+TYMls3CLIwDnMgIv
syq4IOFgCpfK5J9raJTf/DueRuZ3UeOY5lAjG3FNRT1TuAxQ7/p/hHwJ6NoqVsU9
9ddX9ebwJgAxa0q06oTpyXWcCodD9x5dIAKk8Ptyz9Du71BMcK0n2FTunc28Fd7v
UWFrHPF9Mh1PrJjU2pFI/vWQRCg863BoypLymj1OFIIhYQIXIdKvPRbVpTDtX/40
EIuHlMNo4UZBqnlrR9MsYyPrNfkCuoWFjuznyX8m5MeoM946GonNo/CDGxi6H6R+
PeDsqjTZ+bUC93fWUjcixkNKszVv0HMmgZy5QEXj/gqbVFTzZPOX3EaILAh0lymD
yXE4LnTS6cows1WdrBUVChD9yGDNai/D8PDMRi/qbUWcnf19mzfQD1zjROx7Fe94
p+c64eXTk3Q+Xupp+q+fiNY/6WYmhxFWCk/M8WoAZTvOWV9XojzgFQAIfFPruRAW
cIUFPhs0CWyhEExQy8EWmAlBN7n8M3/cZqxiFvvw6cdKpd744KJADKgMj/URYV1c
TsPFnhWZZhk8PxCNpqqNzGitpRkZhciECoTj/eeuGWKECBQKbfR+svOMegDEtqRJ
anlECgqzRePt/3HohVdYFhrnQb8nUQFY+xYd2yFyImD+BMQhi+/Ylb1XkbDlDajf
ZyVGc8T6DItz7QzHMCgwhZOk1Nw6u8ixaOlxKrkuG0gH14FuSLoVhpKSoYqCR9tW
rVw7zbtgpOvcAo+tgmbimvZ01IXakltPEZefXeq1sqqBiw4rors5uJ1qiTApVHK5
6w7HGZ354FPeBS5DLBUqYywYxaJXr+Kktu2csY89BFg3dC41swaYBXFK+RlIFCav
5j0pwDHNMAIyiwySRz0Hx6xblK08fkYALdfs66p70wp+1YBlM20woMhhoLgoD9su
GKanoAvlkU4HFgjZMjrLlCVB/ik49j15bpgwrgjjhNSiycqS5ZHnsk5fkOhCEZ5b
OQZQqnTEW4xHGvO9iphYrOf+ieGUWBaXfezTluw4aslp2MhTPnPoc/jPvlXrAcgr
J0DzQ8PLoIIalg5kCP5ReKXjOjNApknxhbDzBfyEfDvCNjG81id/zFvWDNfbbC7n
fWyW2bV9PDJREh3fKOla/Z+BOix3tcTD8Y/F6A1rSTHUObBnHQRQmvpebSMO3ob/
p+NImM/Su8Mt5nfFMozWLS+PH3LHv4jbExLazQJmCt/3L/6T7Gb44alT7exGFCpq
kHkBQ/AZTK/mUaEytezMhfa86mFRTa6iwEjkpzqMURXTejOeQXpjCLs0sp1aEvsh
fTgmG9XdP/bvYhxkNiB8BoAKbmy6dX5nMlK20wXwARvZ9XCL7ol5SrylMLif0r5S
LvN5SrbKqWpxHca2JFbSiANEcN9x2EvG81LKfO1i30mkTxjhld5AILbpeBPxt/Ua
wOzqO4vm7ySRNP3qNPya4xcU4r/H68zseE/9icMh/GZasCAHqvty+ObFScM3EI1+
Dykez3y8apoLzW8wKF9FyvfXPZTKrC18D6cX7N0HCNOv5FP6Do5eFq1dxYfIbDec
xxFx5QTuX//f+vH/ImEH9Gth/QqujDmCHsrM8zZwcmhxR1XEMsFKo2F188HYvIzx
9UQFL/XNA6vjQUXfHpu96s21en1aGB8fJ6b9KsNNP2tXtb3GU5TFlAIy7JZVQ0Jw
1/okByCWsBVWf0v9wJtDX/rA4NhtR2JIXYT/O4QTgg4gbOQVPg0LBeAqH6wLTrql
01PpHyKjRTwpV+qQLrp88uLOybTRwLN0HqS4PY5JmXLOu4xXaHdqt7NoYhSCASjR
NemElqeEiqOZ/igU1OMBJFee9Vpj6e43D0+9Ve/dtcFy3jGf1fqFkKxk8qYCVwdS
PC0VbR1X3WyIsxJia6NKiIjRGgKGEfJQKkIa2KyW0R3sotlwEluo8ryXdvQ6hUSX
t/puGWJanDqKsPgxDr+OEmqBMH4ZvpYXyZk/Yx0g1Ie8ydcJ3nSczA/z29N0rljl
cV+l9wCGqupWyBYN06IRcDc6aFKKRajeQGTnsvOUQb8u5J3LYxT1/ylZV/cxrtLx
W++lgHYgdUu4khYlCpOvd9VCbki5i3abZhF8+eG0G7nxYctpJ4XHskJnQHGLJQBp
rMGhH0hrwBBh6IR7vPrIi3QljLLqqFgN0jMfy63fajTXSI1/ucW7mkxg2pjY6wMk
TYgx/XXLIU84tbn7RDD+GCxASr5f8JoqT6xLYkMdpaL0Bl3TwsX7SuckkSTCiZiZ
OeaBNCWQxp1KkTs7yQHQQq2GFUu6NLmrXl5p6LxBbYTbfSQ5Jac1O+fShzSm2bsj
MXyZgoi3YaG8JeGIlja5CFzr8i0zrEaJJrYKij8ko+Zx8E+uCFBaOOlRD9qwepIe
uSzgy2Ex33cjrUKFANjcnNfgCgNxWguXkKKrdzePPgQn1MAZ3/KblBtzRmZFqapy
bKR+fmg8S+ryjOOzL9GdpufTD0DISYfc4lk608I0uTdlZodOBdwHIygvTMQKR8T2
lggd4wqbMix0h3SdF5fclCNSbaiH+Ixev0XwbzZPaxDx4ZEb7x3kORA4DfLf3IeL
BOaqnR6xIyiqOrAwG2qvD8//2Y3Gw5qpkVZC1kpJ6DmIbwYA0/3b+tEoeAlkTl6Z
aBDKtxufrzykDHoxgsLWoToMhl/I0MSohVknnZzcj1gBTjhtkJ5dhEcxv1C5HDUf
z4wMEAPXjHoHqvZyknp0QqKelXCw7SjHyNslCVQmUYoKmbmmaCBBPEBsz+NjGd2q
NnoYwwkZqXynRSrqWj1cTIYLAKFiLdtXJuIlGKsdgqw0f9vjUGrAtdrwXUJEGDWs
HH0RvLKJipnYYh898dAp03d4JsPHnT4iZDY6p5RDYLq5U4SbE7bviBLGtlzSiKSR
l9S+NzTKn0CHh2b/u49rYNAXjwYaVR0xouA7HPMSSD79w8Wt4tQbiPR1On1YeLDH
bJE5QhLyKDkTaZLRTCrdD96g9tS1nD3sEdNBsDQR630QOhD1L23xvPsBuKSJwCOn
rHO4Ehq6lfM/f++bdtO8YAVvl3FTJHDcQ3NU+dZU11E1LrRbRXxqumgHsFp4GWXn
pB1ZcF5i65xoym2KT//DxnNW+/bD7H/yMCMepIoNFzTXz6rv6RW3ChcwC/54fjbF
oTwB+lyxrvfaA5fs5lUcz4jViUOJpCDtGnC7IpFCJZ9twRUcR5UjVoTWz7Mt2cWc
kgSaeyJQmhtqAbSG6H5xckX52w3RpO5RWwtbYdvoWFvz4BxUzOibMGKNNxzWu0MW
D10UsgGmP1NqkmiULp4XwE0JdlgbBdMwM2By57qH3eAJju6vzffNYiprVdrS2Rsm
qDgWLbKNTRadoWDNQl4Z1qVBxELL0ocWylyOFp5DG1/Sa6jGXBOMV3nlhn1FxROF
yWo/fe7W3Ylcj1n2bReAJfOqFZ6rGWuGNVd3fW+Njku5R7DXoTRu2CWwoHAEOPRW
zyMI8OA6mDA75J/Fb3yXiIAOhlSd1KdkwK4pXtPjzkGz23op9jfK8SK8Yv9xyJ24
K7dFoH95sEtDCWdKjOOm0dz9XCMePtr8MzUunNqF/hiOHGAP9yeoDaeNuBtHXBQr
vTKk/jVLAT4TH4weEX/bMvOaMZT4h5EsLgVSeRXkckf9TXcxqOyqQIrxnVRD3koq
j3+EJFdYDP6zB4IIeiP3vwCMns/iQ117+I/GgqeXuDRuXRExxPiWx8YEWGWUwSuA
nVDdGufK5DIY4b8TuYcoNvdhYwqBOOxJRL7jXfBoG4rN83U0O4UyCP3bew0y0e60
R7jLRaGG7KDOQSxoNL/Mgra/+InE0li9uDDopPXEc+N8rzJjyHrv6UKbWZaNrC4r
XD7dj26IGFuWma1KPBQSWz72NdksBCXQ8kFoE2nYUuqvL6nKwWfdb0lTxGM3FHYP
k7w/Q/bgmyjkCCgxPUjxScqkn0afRdsVYEMzDGI2yJUOL1ckSvI51hROuxJ9AvV9
BWguf2XdZ589VW3bHTdmALK+NtjifvPeiXJ61sARXUbwbAw0Nwy/lFCYFe8UAd6I
NCPdfbSgKL+wTpoRV0KxCg+lu3T+L4EenalY6vQLimUhL9eEaboqEYKIZGj/TK+S
pxPE6Fq79ybgBiy0IZ8grFGyZFGwhuo0ybPiNTkFUMspgmDPV1BYL5u/i85gvaX1
M3NTPjCnyxifDeZA4SecZylIxTHUzUL5flKoptDe+Yi5xZ5NEdxuZSYH4xFEkSlz
1xTvVMWJYAD3ivAL67iwfC4oBVPpKmKXqYQs6IIuMTPwCU40hIEE0FP2junaqjnG
IwMK98iIaOQDJtJhuPQpdJJvyk2nCJ7z45cqYRF6H1XEDJEoThfmOT+4B4ysxMHy
N+f1fzDa2IoIg9MhT5BdwYJ5lOl19AHmAU8BV1OC90xoKTJ4AEUa5Y5qsQRJ3Kld
e30+kP3UuwQepYlwEA0Ixg72phgyB1aqNeTTx4q1EKfwcwbn4JWPaaQu72Yrq9sb
YVh0J4v8qnLiB0RM36tSWqanu8R4yarIe0OtYrCRjO8yafKRodmq9syd+tjMrBd0
fSzTvgQI2vaCGjNiWtcH+cSThUrqnsx1TSMphqsr5gDqzJ5xIWubhRqslgIvFJ+m
Ov3gw/+MusHss2EzgqXaRI3avwpcAh3RZDZoJabB9fmNef+GvxPKO1A6wKSY2Exr
VWKW/IQdci3I8j3uLr2iSUVfSpMfXa77hGJ5OoZa65BG8I2EnYYauGF7sOqbC4ny
yCTkjjS0gE89+XkcgjsFnMML5kuQMMRyknjkbcqiwvLbIzP6NbcfJad8KHalTkNl
eotkLUrfOeifpI7HocTtOa8gPonMfjeifa24DwVleDSIawAJxlh+vJgJ0rFirZqX
N2FR005EhGtKz/EPddPAEEYEdbgVEs8HNrUzrPMewW8BLufq8/wx4AyeYekKBn/M
4QOe2PBKuvHN2YFen9R7BlUhbmhsBI4DRT8UhqVRrrNI1lI/qI76e46DydxCYJwq
SIYFVSYLVuplqhGZpHxk7XI+DELvZeh7dq3zUH/ptyhPxf1S9QF4cdPexepKWrww
qJHpXlobpSCjAnlS7njWrX2kCc/L8i3brD7APXjzlDaCVroynk7th5ojdBpl1mqJ
FV1kJr6FubqbhhpnHLJix5NCwnb+ehkGDte0c58RgiMuD8MADvn07U2wrKQTs+J3
BsI0ygxId4fDU0JxEra8SL018WYfN65tCbEB+SfPmypm9PuXv+3g8pXEt5H8aAR+
krdHMxlnSBp0shKC5O+MCUbi35GyOpS0oWOMBoPam8TfmGwi2DaaEVShijDebvJo
G9skEdrheuKUbXf1Rhqrip0dgXwluHHmX4voH6TvAFpD7/QM5rqG2YS/R5Vogfbo
aVOj7OegqBkvUIcgb7UiKU5CK3zNaFWkqshBXTucit8zpNn6/vctxwyJ/QIkuZEs
DNnCDAmSwGbrIYmIJODDwBVDUsTUBgW534V49bYZWaLtbZFJcpKSEWpHP4ZpDLP9
RNfK1zE3CpaX81F7mSrTMLcja9hQdy1zYYSG3hHwde8tSzuqHrbr3X8iuRJMWIIl
p3fa3j0Mbf3i/trWAIn3Zw1Ns0kPymPA6l8C8Z93/4VQKHgaMZwgM5PV16OueH53
BYmpJm1sTt5s0kTEiwKKVop94eLfjR09wijQkfAVWIVEoCjteMOqiVR4gKF1vmQr
3B6Ca+DFr13cEwrPMmlEpMca/lnf2IsUW2FioMKbrk3gwx/gt74+/TYCSUT1T/wL
dT/GgqhbuoZnzAb1e3NrVXwnUaxCAnDEKiEBxraEdNmbBUDT1m1j5nOxWi6LMnbZ
/4OghQ65RnUj4cDdY8ViBHoijyvs3ViUW6jug5TolPKLWdjgeTux0cuqGncq59YO
XUHcNl1TVXUfE8oJwEpJSUwvp7XEDylnh58TcgMa+8dq0RVKEC2xgxBr0hjT3wL/
JjRMfyA+mTR8hptEzxxoPq3N2b9BRs6/Kw5nuUx7jXp/D+hEELymsBeC3CgiGaCT
xqYC5igyr0yVGjkKKmUnBDL4E4eVJENyhflOEFhgj2d7YWxjPJGkJxwhgGypR/Lh
+hsM+z9Gi/TsImy0TDUi7izYDlYa9Mqn+o0wqZyzR3wEiqf28G3enw3e3V4DB3hc
jr0uv4QW0FInw3srVkX9/2A3qtauqlX6g2RgCda953Hao8wTY7bHDsGR9F8MENH9
iAZFggN09tRdoQwugsH7Dmx5vFAHvFgkAnRDDhQr7Pi1FzNXjAxo2nbzJ4KKNVWQ
y+98yDJHGXx9da8/7SAL5Gq1+AcKXWxu8o1xtU/Rl80QOjveLxd1aOtvQq2RDgrV
fj1l/IXnQhJXsu3jjzVnq7+isEuA9sqljgD4j6fMcNVYhXYOorO6cWKI731pbZsm
iKCDvUrnpC3IlpeOe83MsVCgvvQtWchwy5eK4VF7sU8tmlexB7ZkCaQw9sjyIYXL
R7nwg3A9kBpeH0syFO1eACFbUgs0inLbT0RrFrTLJt6P0uyxS0Bt00RKLylGGZRM
pRLRyMl7BwjjbNP1YWA78/nSXmzvdShsIgLkRhsTwsNlH03rr4eBN2BwCKLKW2gC
0CMe7jZuKV7a6OEH6NSTgUfyCmhpmrRqsTaxFcVgu74AKAyExN9Qpc4DVpAu7KdE
KbkTVW57hiTZ/nDlyQ6librncEU/6rNy/An+f8ljQ2larxwMGTrNO1uCMDeXfEev
nV10Fy4uZ7L1yl1tfW2mAn1bvAjFhwd3XY+tNrJ8HaOoxN34/WkTrRQX5XwQ3uT/
d1f6gBdQc5zOWHN4E+Xvja8Dta6k/Eyd50UT6VzH1GDQLgT/6Fp/SFP0eNrWuhSl
V5pfOF/VXqW4QnMdJFDZve+7CY0TwsLtz9GC8doxEk2X45EUQ3hRZhIOOdN38Ggf
J6C1FoI/pCNEfbMflcSBiR/XVVCOg/IggREaGmo/P1VCuZQpsBHwxHXa+rjvwcDz
JFdqq2TRHsM/M9milDXsqbB6tbel+72wuwQwHQtxxw070JAahHqHs5kBqtJhnsWc
pyoPVrB8Z5tC1glO+fs52IL6TxFrEGRdnRny3HUytOaHy/DYAa1hj3U9XRcnuAVW
9fEpYAOY/u8m1V36zVHdcOGJ7OJjOg/UMI8nCQ6fLQ/Ew3ZICNnwLTVTDktFY7iv
I0f1CV+wvIZtYZcB3qBWDbIIQfApbsCYl/WR8i+oPMDORGcKM+7XfPyl/P/93LHX
iN8xqXF+RFKOgiRNTjhJMo/C6lUJcAXqZeQQPRkPUYI1MYlDE8eh5L/41IwGWkTw
doy31+1ZixywmD8TVqBZjXZcARWa4lmT6THRaQ0g6e+uPj1zxzvtI5s83y+mi3G/
J9c1Ypxdm0upq1HqWpAn2gX2qTbY90Z6yFcqq1c6SiCosv5HWHc5jwQBCD/Wjnn0
uwPEn3eBbHBJ92biIPhe2kmdSIR+VIhr/kNi9cnOuLX5s996ikNQongDiJj9DFtU
yo1l5/DF0+j9QGJstMu3PAEjwo+bpCheAyW92umfhHYuCok8AFV+aedKl/vqWLnk
hjkT+ZxICCRGR6U75Ir87yz6wfQlV9ie9rrIsfSXEoAIOWDzOBEO3Qtrv7gNKzd6
J4r6/o7e00ORklg7Tti7MUkhg6QMHjDrTyPHqhOp0DzMOEyfth9/hE46jfmVXTc9
68E80oqXL55rsT/f5skKWtd+nCPcB1vMSxBFUEWhjv+S5dTitWMBx43arvNSYlcA
Imi4kg6/HlYz/8Y4cEs9YSG3QJHtCfFi0pRPiuNK5ZqozdFP2HTyKw729DaByahU
e6HUQZqiOMx6crhEVtKZQLNYFJONA1ZUHyFx5Lzi3KpRsEf2A5KZQ+gXGWIWtjPP
xYob1Y8RB1Exsd+cClHEGCsRI8q7kjZPw//27UmdxWUBG3qCZq7z6h2SjYlrI4u5
BbK4OtstYCnI3YW13WrvE2yvgZi4ho1T0pDdFqjdabBTEob2TJBTm8LC3rRWOwbg
Vffv85pbeLhileINosUuk14Nd66fuSdFWc+QGgjmXX+CsAGuCSrGIrWIdH86uTXM
Y6leNmE617W7hzZ4OT9e9ANBdi37nAdFdVeoZqQbY5cGqQ5P4CzkvUZTLgmUxRrp
g55ciUM0KbDZKoS/cqvIpox7qm8poTSmi33V+bduOOR88+fuVyDUMIbdZQSBc1A1
zEQOw/KvPhWArjm9C1n0MwhZ2SD65WZ8mzYINZGUzxQOLgm49bbtatdejSaPrLY+
mBy/8j4e6941GK7hIMObv/usynN3rxvecfNHAoFHopbrJ4mwFqD1R/ABJsp5jIRL
P1VbbPVobQHqyEW8fpKklKS60DUXov0IjjKoL44g6+mdPI/cgIOlm8kgEDezGp1G
7XXyx3niug05Agc3yoaR+8eBQFHO7nO8IWIuctm3olXVnrRlNFLVXRiUmbT+n5C2
qNzbywJJ/PJr6yDHl+tKoaIFzC/DQbTneL7H3iab/WbleZVAW4QqwwjyAEvOik2f
Vy1Etgz2SjUuyqXUF/wXrs33MgJZ54fmJJ1pZt2+6tBIE6ouZy+Dykv+hRfcYmKY
GQGXdyydS7JlzF1E1lQeepJI/nZsrLufa0GSwUN8CZdFy8oKH70x7zCNOMpQ2I+y
aWjmLwKTbmfW1OeMVYv3ogoy98jPiF41zFa3ybgE4RpB85FyewIIrXMWXuyNC0y+
WogGbWaA1fpkUsnni5egt2kMM3jV6uWIpVeRW5aJHhHj8jSiHwjl+4GEM54tU8Lr
J5oK4WvJwjgAVX03xSh1EXF/Xk4CZlp8ijaxHXjt3RSbH38X+yEl16uNusoMWZ16
eGHwSVeTfndPANn/MdCNL3dd9l+U/dIKfz+JvRUAVSBIU4d9om95iButpl0Sd9nD
8T0H/W93u+dXt2RubCyIbgsU/J3yvSoofltNPoVKFGLU08iUvv0NrHHbWyEPYuEK
MEv0eJg4RpYbbznpD+WnKczeyjZ97qwJ9xX3+AQhi1UGWXvXSrsbJL4l5S14z9Gt
3jGtiojWEcFeIg50ad2FT8dMCMfs+f6i71Ps1tKGcuWkBVtu6ayh7RVfzcxH5bWl
dqsFDxNHdwRo9jdt7CFgDc6jF30ggIjuQ8uxyCJ1TVw9XO7ZwqPqAJ/A/3on59nS
MCL6UlLpk6tRu4FsyC4Oz/c+nwNEv5D5oVbMT5xbcuVEOybISFih8P7ujt32xrS2
Uka/Rk9zaI/8J5QV0YCDizXRD4fKHZIFZ4XzgGnJr6KAvDHALwXM9A/FxgENEwHU
1OmQP1KLp7Qh74qfcrKOL+Liiz/w2VII5TsaTwUm1uNk37YmJblEAZnd38Y560cw
YeSk3eThYsmUiABX+kvYyEx/EWXnDWezD8ZRl+NIoLDOsHV2EeS8eU3HzmlGV67U
lNmgnHsz0Pr6WpwHWBjMi/LtStoKdoT7Rhs03TPJADd1jWCkc7YD0rES94e8Rxp/
LcqWp+zFWsBLnY5GSrvUj3xtNlM28PDWIF7q+gSUTc80rodQw6MhM6zdqa+DinB5
Qh1H55WhqL2Z5WYqZU9WVi80ByfIU6tzk8d2pd4whluaVh2H8GXSk+SULRSGToCi
CqRXlElRVg+sUSlOx/5pSdv25c0gfyzQ5Ayg7hvHwAYgDYQexgejkpr8Dubnt+iM
ufYAXIcnxm3OPOyZsAFT3WrVlNFeycdJpun8OgR6BXGAMjRZy/JRktkTPy0ljZ4x
MboLXF8KKoGOD1oM+K0oAxAH9kB5HCe2dODfuDrFjcfZWU+di4qyhzNM9DlOlHJ5
kVWrddQAQXyhSc7ChgUUPf8OyrBo4IuVQorpMlz/i4CEX1m2CdKtZe6lxUd3y3uZ
0zLkGMuwfNu/GOvFBXegCJv6ovWOlHoxKFsfufQeCFsKonvycr9GBPoGP8W7sfj7
AI5m5xu0Y1uOP7lz4hV8ash3y10WGlAXM0EvmJBx0lEofiJNJfQ74hvE1qQGOlgM
XJiYpRR9IWEY83EFwmE1eC32kBMbBy8JUK8aaO5CBwH5GlsTSc0UMXDNFtAVdbad
4tcb9BNGS6lYHPsVf3KjwdcEMM3CUv4uz2xHmOwfy7kse49JULXgPVDUq5C40/1Y
rmMtitIkvEIEESX4BXDfOAhk598p6jJO4PgSriBLw/nnxGuoX0TtP/CfKmMHkeFA
oMJrFUKs2jK5n3Cae8PZ5CNvcIvn2C+Ttwg0AXjHyA+V+rHspTd9QYN8QghOaU3+
Fcd6cw/Jfyvgc/z4OGujTQzKAidZqDgSYjBXueoJjFjqxaZ3DqtC09WDDCRbmiVb
GKAM2yp5sAEFSgnE+1h62h3ZSvv73zY7seQg12uhH3NAnsmxn+UaUpTXe7dqTqzt
q1HY+g9vVYvseehmU7tn/CkflB+NP3AxZjBPDROTHzQsKxAlBaQi50s1mnCMVtb+
Dgx2k0GzFzpmWfu6lvRBF0KCfX8ScLqNYFW5cAL3P+b3zXxmRcKXwG0OYkHmmckr
ixZrY2HtdZqtTn/6/AW4R8PsKKIo7FVVMybEwL3hqunjOQPo1lKXxIQcd1pDSpSN
3hPakASC54YQkK5ERhmZsn3EnAvd6ovClP3ptLZ+aaKCZQqCFMpciKlPKUTF3R+n
v0VcG/1Fvv5fINdYtj/VNnXmUvlRgXqDvp09OPbp383FKUAOdh4KVf5+LIIfTIcP
tgNaHULlJ/8bF4ea1avHynP2wbW6YmD3g6r0Spy+TJ89wcVCD1WgKEjIS7tShibY
CJAWKZxEl9IsE0IVszvsIDD7pKJ/+eXlUykZsGM1RctvOGQVpmncOb/yLAdiIfIR
ibY3RXmU0459C3J8kwTY2xXj17vkMxteh8B4/1hwFT2fwGCDmPqGAEk4i0iOw8zF
8VQFYvvKVHvNaV0CUaf695+EeXbVq9wPGcqgA/q3Xzgj4wFA5nfC7W2QMg1sWsNa
x/dkFtICNsPsT/GYrhSEPth8+IYnVBTg/wiz4yu1KCL5rl1kmX+FYJ6VCJOvxgx3
QNIWQ2UmX3csaectbgGnqwsEe6W7sHXE0TBr2ZPSrYiBIfXWF9BPu/ywqX6V4VbG
P1A88eNiH4tGr5xybtfgyVMOu8r8zGQI0NQLQ4RMydWH3o+5TGfXR2+zQrnjeRnL
f05aL0q6ZyRkGOwpON08GUJWDk7AED1dcWNsIQo2pG/f+sT6o117szSsHsfeYByj
Q+CoV84C/eD5FiFUVVUD+Iut3XX34nEoJPWYAOzUgC6rZaiJGFK6hUtdTrl2QCLN
xmlcC0xcrlQyu4xnFbnRFioqupnAxELawM3JiSyA6OJ1EjIOTK6MWp5hwNABwAqs
ylN5X5c0mH050QgGthSakZXJvEftugO2SXvfLn5A8kJgy9sDWDeXdTqfUIv0AYBQ
zxGN3Q3vSvG48fakBmoWpBIJ4isqLyOCQvjH37Q69m+QPcFadTMjsn7yOyrVzuMc
lVFNGA0FQ1eGOTJ7RPxYE8LGi7AhKe6yn4F6Xa0Q2ZA1egfctMUU78Dib4+tNqYT
DbycvIJIIYQfEWNggXI7LhhkOVV7lUTpms9PlvF+AjHqn37mtPKKhrOKDtBUXGSH
919rk1EWiMZKy30ZJIlWG45yK5qR0wnkCO09KSycSrzzmmVHmIYk9qxEdKGRVD/i
1LQtpKyQ6w5as+GtHCO52QmRft64ezXsZVuLPg6VU6CNJV5LYoVSMY/9G2oKuNWn
qbedeRCMm0QiT2mLIbYAudIj4uSKT4iNt/8lcm3wwIdYsG4lQxszE+kVaVeT/+oj
IYechrmkl7l7zU2SXqzXcCyj+LE5L1UB0NObN6Yp8TjubEWh4D81/qXpFsSndIrA
9uJyL0f/yKhxfziZ536pEat5qmdaGjU7V87esDQkBtlOsdU7uWkKqNRf+MNlkoCM
DBmFYH9+FOOM9yM50akBDP/fVjGGRsfkch7bHyetryva3ulEgK665XQu9Pg4eUql
QCVoq9C92xPidgDE/L8wGF2AAS2RvyTHx5uxHL5GA6RT0qZzWhioQ5rONuGAo4OG
xaGaVoUH0FiEmDVH0tcckN5LUCJOvpoz+/kQ7+OmuSLB2QGeYZFZNoGkpGzFf8IT
5UE6w73Ex+eA942NMArl21/nugMKlG/UKvJHmaXQzd01pI7HFgS1K5S+LBTHBeP/
1zco26m3sgELl8N3B2t7zEjGIXoFAqPzCWsRb3IIx93DRvI+7aeEioNgZQ5jYE/k
9CxZLEyAFUw/wuy04aTvw+TQLEik6O9BfEUAXexzpacFiIW2Pw8bRXypbhZ/yjdF
xX/Fo659KPS0AmUPhVt3Fe/USpd9nNaKEQvMWkcE5ZrCi11kn7FhsIVqVPMXoKO9
cI/yi/TltPBWHZ+To+3eF7errkOduH3jT0ziBt2fG31goEWpsMGIhwYBFTPkKcAy
dpqK7PFOf9akleMbM7ifq+AL8Lqd6Ji+X8uI1rlyPrtz4ptV9SHfPeIN6k/CVG/b
lVjR3+r2nwODPac+thAnSq8GiOduDjpxIU6RWGS5U/NCKniyNsq4dWbgFLK1cLkp
HyiVxKPkK/DTZEELkcUbhI5OulRvu8upgxgVHa0XXBDVuvqM/IsdYP0k3Aodzsb+
cPlViN+/KG9fyfnDsy/SRV/ZJIVv1V7t8ACirZoF1FXRwoaMM/FUlYsVsIXBSQBL
dhX89dh+mj9kWbyf3m6u//VRW8kUz3nGKtyX/OCWIBvFoDucCj/e3ggPwsvWfJP0
gu864axJOpKn9iXyAssb4lGH9BJYiamVimecgTTkoYJCdpHtPjEDhxxydHNedPnr
nTo/3NJlvLrfmAvPSoc/LZy2YPk8LPcMgn3BHVFH8NJvwaXSzNMH6LDEzWjWg9aA
GvS3G1sb7Y4dCTfz7gHOwDntuJbB/VYX6n0a7SobOomtW/zf+2QwxIIeU+RNmuE6
6uWEdUN5OcUcaR1jYp04QyITYytgSq2HvwsJ/uncVnHQ1NEkyDjGfzSuM7HS3IWa
/hxQAP2k1/V+lolof7vo8o9x0mai5S7dOo4enLJHCIsIjq1TwM2AvzKhEEZmEK9u
7Vxk9W5CO+CTDlS7RL9x6cd5TAStIqbAW3L44OtiUjARw1pqLxbckB/IWduldfny
DuYuMqZceJWtS3NeSDCiFFGmEGhKC63QsLZm3kG2PNzHOs9qzMdZ+UU5PiH0a5xY
BOuKGzbFYBFdvGzkl6+FmvXesbnXrYGwti6fs2A2MATpsrdRP3HrzTdcmLuFtRRn
ADTKAZh41oKgroXUpLPepxvWOLtfMMgKVM/wAScN8XozJWG6L9R7bU7Qm6K16zy0
PAMaxX6CFsRzwzEKeitvbTHb/NnPr8LcXkJzrraZ5yVp6MMl1C9XAkv6EPo1ydfj
/VdfQffOJpNfYgpGoPTmezcG3sTMt2hLJyuM6WtGe4TkRJhXuPOL7wE9vRI0AYPl
cZO79Al79Uty8ia/g0FSIzhaCjuvfG8vjH818ma8CT5kTkOeDDN1PbqrhMCRvP23
cTbPzoEu9LsHUKpFPFNoYolTJ4OD5CrSpV1YQpRWtXIQdZQtto6hEeN2ark8HT7z
SZk4ECQWpXk0UPcsDpgnNMNmJTx8Q7zXpT5u1YmR4EC1OURdI6DytbHWagZ4Bgke
xDAv4jYpgfBp6toDRUtMrHkTBsoVbzS9On0UtN2iJZFjPS57P/UiQCwVEi+f3Aeo
Ei1/qPA4RJybNIa06idWJtKkJANPwkkdZpdgvhPiMGF2XwbMFU1X8N7OvpYylfs3
/6IhyaeE5vZbT5f3wG9UFIlCS0mphs6X/tA9ROHwHfTUEzxJ14Gxpu0Allg4pTDI
ED+1XfVRCe2YQrrhcIO45wChM2Yrb/pbnKCXTukjSFKJ7bBRqzXZyudJA2CMS07Y
7TI6D6J4ebvC885ao2N9hpJIwnOztmUBrfrNAEZBSwiPYWMX6VapYXkL1MmrCq44
PYZ1yIl08gHNDmVVQTgBy1c6FDkD5OI5XRR7eGlU75FJltXgQHu/UhKxgC5QMbmV
x/7NlB+xTfN2X9y4ccCavjGikr5fLqNpyYIjYtPdzBAp69Wic4qkh11EltrWn3Sl
HRjd28XYlE+2uXhucvx1b8kgyPJJ7Lfdd2MSNU+JkCYat13xzidDgW6hsufXg2pt
zUDudSBD/CRWoW4LuNYaEwuLk1hikXGQeJk6vA0xfFMseeJakA9U88guLk6nsOQJ
IZw2yaC1tZZm/iVUClUV01kONKOgE0k6iR4IyiLo6+9Ak0F39/B3KSZssbxhGgje
kpbjgx2EIuXXLnovF7drM8pJMoXumug8X0RE0Tbr7Ijw8BWbsOE14zsxwhmT3C6a
5xVnWO52wHtvD9ZsJqrsPPYLDU+/L/RDdwIU3XidUZ+zpdZlNsGdQP5MsDsP73Sh
/nCculBtybIw7c4CN20K8PaiTiVrsvjaW5mWIstf3EmEoy6KQ4wJeqPIQNAmIdub
57rz1XFsjC/RuHkxvffvnf6bTS2Q4LmxKFbHA5cGIqMyYkLwPtDGtHuic8KKZkpZ
kP/LSvyeB1PeT4FfcpQa0sRMhH4TJ+ZCdtumyHgbTC912PnPuatYnxDud2bAxOHm
Vvgk4kxNPgQRQ4w2Md+oDxYBRcqJ1y9qdhlQ6/QkZhbfpBPLq0yIytJ/WYGHT+uC
0sw1ecsl5NpbPRjgWq4XDCga4pTwqnaRrng9aMVluXfNgt4cHQ6tnetprqErsnYN
oNVOZ+tAa2XXXykzT+3GnzQu7Unom4JWKSJHnksTK6l3Mv3PnpOC6w1Gwo3FEkyU
/7mrvYTes3jRrYMLJhD4vSt7or8i4JCHrMExQyAuwCN7c/0JnefE9V/qyr7Ec8PN
1TAV2tnHJmFHCbEPwX4mYB9WNH3neFeF9m7LjSLvbgxq4CadcTJZQ0nMC5JW5S2l
3XkHC3imSL7WeYXbEvsJKeXZ7p7qa3fgTu56YtShPsahHGs6Un9wxzFBo5IINAb5
XIUbTK+KjIYXnNYBsesb/rTaSWKEeuSI8NVmMHV/k285y5ccClaYKuI0aAhQl2X1
ypzRZRZfcSN4XvEl713dkxnYCZhLnwbxw80bsZjMC1BJX+Jq0hSGemlqvAiMTvN0
c9VZHLgghW6hgrT496iTb9qQtnlQwexSJqaWw4BkOYRmDsppa9EvBmke/JIfBXmx
UFaxX1XtstSE1tDHhSg41zJ3wfMGAIGbWk6s+Wjb10uH1H6e3XdJOpE8E0/jSewV
zWTKgdgw+tzAFDRJxg4CaB4DJXiDiEEJEp4PQWG3C39PAqqgYW6bnNnngPEwxTFU
+KN9UHXjrL3mrWxbvVqrIhGV2lPoVzS9Jka7bCrraOeGWHRefLHoWVtMRpG6+HcB
lAY7rO2YmEtAMMWx7HfsfkxWhy+bG8e33SSP35j8iNvsjwyh/5pHKaF1vY2rKlzk
RxPRaQrqVjyysOzuKribrY7Rc/MfMJzS/T0gaZO6PZ3szxoigQhRqhSKMDr6x9x3
Fc9qFYeDRFUq513QOBG0nb47kdguHXUfRjEXxbuUgLvvsUZRMFAsMqXwtIiJ6Sqm
gB/6QEOskQ7n3a8Itw7swh0MhlUj4pyA9C6a2oz04E3+l94+ZYkDACIPDeOfbUfj
0w+NKXbz1M/noeVlwByv1RW3U/RZdxPaE75ysHKub4SYmS9rXPpRmsfNYMiLp7ff
L6ejmXjPHSs8EvxiTcXoRbNEJAUlvRuwo8vJGgKsWdj67x4Ky3fzy3n/ObRFvom9
V4X7dXfU7Pn/amoSL8kvW4HxDhOykMMDtiCiSphjBJpEnmwpXw3RjpCH9zpcR2AZ
dUZ88tfpmCga+85Egd5d9RkL1dnTv2LeKIbLPL1QoravIRHzM7SpT2CyAU78kOUU
Rj/JN8LnaYdSz4VsEigtCiufWGt6dGoOOUxR6qswe9xXvZ+X+7izlueTpXqDFU6X
uwQE3fugs3O04IUKjxxO6o880e+BDOWHmiaeAUsF100tOvTs9U4niSlSs9mCAK4n
s3fr/G46EetK3oEubg9xYX0GoI9DhEHEIHpuN6bKTJnfJoTbPucI15rAsA5fF0+w
rdoUTJQ/kheE3zMsvRMSR4D+tD3yx9sXUMdQSfeGsuENywfosIHblC/uZQklkEnk
rPXdF4Pu75SIMLx+Z2UD50lb04/FX99/SrjqlyOyhJ0AX7ukz+JvqTb5P0rzPvrg
PqsktLJrC3yII6D9YT4Q5MzIrLXEOtAie5CF0/HR29BGsZtXsFOVnSqBHRZAE1hi
pnoWS1AKYcTOfTw++DcnVAh+2wF6HjuL7cOcgQWDR+lQag5JOiibw/cWLMrCiDHC
epI6vE4DBGNQ/ZfIYRDs4wib9NrYlsziclTZm2a8WAzzP24mUOSEAn049/SVh6l0
yTv/Jr5AWArxLYSYCokGe2XYgpN5IeOvjqpaoa4gUcPeTcEFDi1RHsYvR/1KnzNN
RL9kYEx2kTVWCYysF8IsjANLvMyhr1BiatgFBWzKU7qfCNEe8Uto380QeF8XcLN3
pMGSzEg3U+bAHyj1n6cYO/5a6nXusysc6UDTNk2xKf0rd6aCxggzrZ4/8qlYb+pM
9nBCUdJs5CXqXW2Z45Ste8HDx80iLdevuSKXatOru52Gm84oGEh2cAPZiljpv6MC
jE11bIBJZJwBEPRpWDWeS8jhdag2EXlehHGkjqodNpj2jTcDsHnxc86pZcpmq6r8
Xe0l9oOUlrintL6jlfm2WgYX1PT4jKOkaKPpcEFPz2TzViX4jxN+8RNxnJZc2m9p
/dAqrPFzU6TG4DBUtTZy0UJvF6t+fnRVMDYpV9DuFCThsGqWXNzc4wBJyd8epsW2
hfkIWx5tpJvh/Nns3rYcSIcPhn48V9tmmNeDT+5msw3T+vQ+2Y5khTEwanKuN2+C
ue0gsDbWsNNTXq2QV435F/VOFvd3ylM7bBwYfV7LitgVkPt+3WeyuhvLC6g9gyDQ
/65FS2JK1BP42zzQwa+oZ4LRe/GG0DojwkDLc2AVcKdMZdkuG0GCQvjRopH3pQfO
nDraHmFOff/KMKqmfxGR84nFh3Hh2j7RyJKYajy4w6RRAMzwRwmgvo9R4zFXvqtv
AMzvem8N99uEXXz11TPGQAA1Vw7AgMFyqa1aAdngJ+rAsqGCwgKUvhNmpFJe24V/
1WMiDIlUlmxjKOAlzHQ56zdln7H6T1NNDgNeP8MrFQzyb8bsYwfP46iHOVA+Ltq5
x8htUYFmsre9LeVcBCRazyTTyrJgQ0M1525B2jOVlHwh19D3oGyKDJj7TD33FcFq
A4ckPln5ljYKrYX+ux6pXnVHd1rgAfYMxFepMpqm2BYRFf8WY3QYsBlL9fZ+MHLR
NPTg1jiBQnYG5xWk9wluQqHy+XmEOnOAl1uAGeV96n5SwAEznx7wTdEDwBB9n8fm
mlnuNKETFrXj2PXf8MpfVORb5BZE7iXn3iGv7emb3ySEHoIStEySqj4R2LV5vAwT
bmdwDLOrbiN3NL8/ZVHs4pBOk5AhHdacvj9GKnOZR1wKjk/OYwRJaJk/vRGX82rP
yeRWV0FNBNdiXcqu/u/hUPbQqvJP86ve5ItCIodUF3f9vCoJxOMWWLvxuVjcUEny
YZZx5g+EQGStOhOaNcln/kzgtPIqNQZfF+7uThKEKsIWDn9dtUzsluCvmXS3hJH3
eajBacJ7HSelkDg5yI+1eog9IaLwjOm+k+3l9/lJmNFTYTsmHXtosazGFdEc5h2X
OtrmCtivSavBds5Yjpb1Z9zBYdA+uPDPSicc5c4Hod4QGdWjLIatT7rVdye6foZf
c/vYvJz/f95FXAxjqIG8/lV19EH6nLDE8MgyKHgtSUEUxoY+bHvmRNEGxITIhp8M
BhwtyKjLt5D+LKG5GIehu36LZOnX1yu4DC0MVcv9yq2MRiYRYAYSg9o8FwHJNBDQ
+ep6OTNC8h3hQffmq8ypProeoCReS0lOiJYQ/SmWzaSL/87Tabys/amdkpoCB/iv
qFVbz3vpMdaGpPPD0nkgFceRov0hD8C6tM1eNSiwsYqas08QCZnBgU/zdVz7zgQT
F1Qpw8b5/Jg07D+UA3E7RIWGXLoYDtLq8sjVzmlZeHK869vZaTKqL7CHzzEW/Jhw
ua9Uj1C+M+HvKd8J1cBM45M2tvEs9TEumEvVAj2YRF8yDNSAwd9XHdFu1pmm9nNj
cKko7FDfucDc3oz8bUDrvC21sMs8bkednWw7N4awxn8WwJCMVBxIOAWKXm30BTKk
DXQMbmNSnsPLeBYiducuuE7BuR+Fftv3z2fd6Jpvldv3so9JUQQLan6DzgNIBicv
AhLnD2Dv75UuGWgqd4ggj5CwvT8gpNRT8ZqqVb09hJ9zm6iSO5Tu6/aKMfDI5ecJ
s4hzClzJGtpc6QP/HM7hs5hoW6pSMTibH7P1mB5augFdq/THZO9pcxxxMgA2tms7
9aV5z6oSOuzOrlE8yWHC/jhm3m7+MkKnhcmWZZ71qmflQBuAyUd064JMHDf0kXST
NwcNedXIBPXlBQGaD9uEZlavOGtIeagwp4Gdk2vcMgOgBk/wsSo8tSOcMaGycC0b
Dlh5vvQqTEskaF3tJnxSjKvcBu66iVmqu6HF01HnZC24dNEKuKWEeeXiRCx0H3AD
m8yawu4Ju4Nzs3yjhtA6VBhAPxsBEgz8AzfKyHVTZRej5DVdY17FI5VWLZYD4XEq
CBWm7pjTRmz4o+HCybwoiDY1kxEuRdkl+PWuuinS6k261Zh3bv1/GDbU+ReDpGYV
kEkWhIOY0rVOgZJpDmPhwCBhUDtBjzixPOwRrHqWA28cVomwWAth8i0FDxsie3AC
1hRv+moIQxweoDGP7GkAD9t1J9IB55UonKl9IuaMSZjtPZ+9q3ofTCijZwxMYbC4
67nnIOJxMBmoV3srVpzbFwVKMP94zfyKxfIrVOrRsVUcQSySAnl1c8aIacXYY9Ug
wq1iLDVOn8t1Fyb2wtF9pP6H/gwc96a6cUy71CM2abPu6Jr+N7Aq6I2cL8rU/SsJ
9t0GeNnG/V4JJhAnNgbeE73pA26s30MgHOTbDKRIyk6d26kFXjXWZuwJHkGwVAKx
vM0G6LaTM3cqkEz0/0tp5A5WwbdqM/DsXiowPkZMBBbqJY9ORjtnPMmFtSzDkAAg
ADVR5M++seUnsUXAwdI+YSce+ySocjDcAq+bUlkfh9PK247NtwT0U2f9NLOTwOfr
vARNO9fzKK83Sydf9ShCqEd0DamhCKGVn90vgXR5ruHYQIfcy0CBImJbXCBlv26c
h05fsxRQBX2pGOcrg6U0GamPw9Rd13NSuvfKcIG9gK8V1+sasRv/P4doVN2MUvf/
3TtgrswJAJreYTD7i+xNtL6TkQAo2L7UZ9ayeG+yiheV9pH0G3WrsRSt2VzpJnZP
A5wymSZx6+bQ/jDeSDqXKRm3oitXsmonhbO8nEpwXogvMZC8AWA4SUaJsBrzguIw
Vko92XS8CeUSbCrcDodVlnSwUg6BEh3wwPGF03WyUD/kgXtueYTcIHyFEWBVdP+x
fKmI+lHPShjhBkfsobuHNgJtqDuoHnJdZM03g5Ojb2fpuUjevrNFfpitXkHZHwVm
P8sr+t9xM/KMR2RN0jORZYds/4kBkyCQivhjxgN5Oau+wxDvjI9E23s4BJCC+bf2
ZTy4pgYLYwKlTEUIChUyiKrnDBbYsBB6dqk68uPNG03Xsi7SIHmoZ8Aju6NEC58S
lTuFt9b1LJuuMW+c0S4tY0eUk8ojsczfP91LPiR9lixv9SWJRvE4cEMLmbgC5292
6lOjmHpaohoCP+5Ang3QjEd5Jh4Of9wJr8ja+QPF2u7UgMUDevFTSPaMnDuVRdY4
VtMRgvPosdrkJC/AKBxxFEn/2E1TrM5tXLmq2XVlWs/Jx3Z5P/wNuzfiMfjTqjs+
K8N20rIMdu4AuhbOh3BRR/io3FdHP7TxxiZ1cq9LtDHWFyKQG1AXNhdJlj9SJ4jX
7caTldIuRnbkg0vguKqXKj7A06pWRfYwcwP1mkKv667yWc2p/gfL4cYIZNU5vqhq
MW5GpTdhUKOtsgMV39SnK0h2cPlD4NsQtclLM1Qk0P8DMurVhtBtlikRYqR8pwNh
V7sUATMO5NBiTZslivFjPSaMFsD2ZSLc6va52xvWXXP5AMyYSqN/MB2vZ/f8AgxR
wvmRfzFZGlW50GdWRBPWH2rnpRNmm2Os9JHsPyURgeE7t9EO2NEmv3tI+wfi6b7e
Ur89yc4yn54AKDU+pT8yg685MJWaw5BV9gMCGD34NpL5uyS6QXEBZbLKUquyFCC/
rOUVSxipPmkkOcs9/P2sPHgVv0dmuHmmc+E1oWxzRgQ+RW1x9l8MmOivPvimXBIY
FgdVNF6X8wvinbnWk8FfCAKbiYRzjHsfGd7FVbP+q1HSqG0tsP3tUZ19ajHf+tvh
PaGKF5cbqlJ0gqGeFTdqOuGv49L3Ygs9x2PRR2OdsS6rviYi/jQY3+YkBg6lnfE5
qwa5jf3OMnJhGpwk95OKPZgMvvoRPaKJ0+uNvMNYvS4I4MG0PpGbivI7ilHIgoHz
9fFl9pAeE0iDMGa3tsbw8fAyyLHUcS+2kXR9FdN1aPGsnXyQDAA0KkhE7tLP1yeJ
PD+7SZkHyQN7pYKC4EMKQPA32r0caLd2dPXPnr0Yw7pwwc7L3cYWYKpr8phvaGEs
SbJ1vDYRDcLOrxQitIk6Y8LKxItqeD3amZgZ57PHIkMLAJlq/SjNOe2w0xl2AXT1
bxnv+ae41qijqI4PBxyEXn35Fs8MbNLmBAf4PPYU9gkLkevbBlPLt2O++6ZIN1Bk
5VyLuc6zgwCW/WStr75j/yXQteDxq/h87pLz4K9WIG5xPwBnmPiYSrus21sEeoc1
XXf16DMYwQ2C4ML8EAcDU5Q3S5Zs+qM6a7X1dNVcfGf47T17Nk7kXVnbflxBMIpz
7Q+XD3hBJoZ7p4YuJjogEvh0YPn899nZMe5MxUFghJdPcXPzuN/By+Fp9JQtubNT
uTZXJS3Z1NT7ep3y7ogWkv3N21/gjPKdH40V+EPC8upTI2h+BQ2VHhndrqTVZoZ1
G8yx0imoZLkTqlwa4txXjydL8Q0fKdAa0xMcdPdmEiNF4Qx/mVzrIntUIrNRUOIU
cCvbMPB0MB0iHl+m2mNNJi9sXMiow6JLthqFX7z1sIko/WnXOliw5PMtlMQGul5z
x9bMVrXumTUBvUZmr69EmT32SdPS1IWOoizDRTTtIuvhimVIrOPVfGKkqRYXuuN9
G8cW0uamValqxPYLwFGebzcQ/Bk5fuxZgF7Kors0iHq5tp84lsqdh3FDYwLaTHri
prWKTJ8dIPsh0D6nK3gaMjG6HtszrXjgOmOQ6n71jcowQ74ZJJ8RG42nhUlAxwZZ
zOKa1DKwUYMzbweoLHIvV2kpBMPwNd10asieT8CB4GGoq8u2uuh6C2aLlf58ztHK
vp+ewASD7TgAJlVDxY+DiXQoIGCZYrH5Xmaa3znEpw9GAvXedahq7RE6sNZ8FP69
zGAbJa44xAbrQhxNynrJUm5tzw1QeRizlntuZh8k4eBoakCirV2V7cbA+b4FQc1i
aer8RLplboL3Ut7z3gHeNei76PJJgt+CGXt77bkzoA+GBPc7xb3M4ZNn2TYUHm7K
q9EqT/2WFrh/bMwYpurfuMNiPpspZhIs7zqKFIsmyE4v79X4VGWhzjZ2d4nbReQn
UxYdystz39z4W5ne0cLdPdfoh6yMbvptokiDSfi/PT1dQ5BqbeakrONwo/3dY7iy
Jg36MKKPbfwbo62Kz2aqyr9bqm+ueWeUXKuS4TjMBC9HwPddoBuzKr7HdrJa7QHN
na98QCgJQ5EM9Tl4CGuUVgg47QqTMgmP9i8dbKPDpVj6m3Cdr12vjrRbNd81RV7J
JHnMnr5/VhkIozfEqY25a7hCWNzMMpX9hme3W205EMWQ3gweB9aXbgGTprqg1eaX
wXDEo3xid+CE0A379INr4Mi9/Kl3oi+ZZyARR7tELMkVvDmZpMUzFVRzTPYbWZr2
nvDuRZ+FVxuRdQy++XJnW63o2E94Cg+V9xLinyv8WG4MdESvqxpyC+UlHDEpnPi4
scDL4n/pA+q8ruGxygjndzsMoJ9aZwF7v3qDrlnMb+kIIfWHGFIMBWDrL2KbdITl
fuh+xkMmXVpukh+XKCJ6L6Uq/zHGMPpgd10wdQY2OOeHLILVyjxSiIZkbK+X9V/O
wPjMtJR0BnnNrpSVraKXitNOirbjp1NokTjmoC3kFc+rFWJSsk3pRGwBZo2LsnaK
Nezh2U64D5hBT9YOVcxILHklLwJQLSzZZKC4v5hINGzJdDgrV21oUNVQmxQYqtJ/
89NY99Ah0sHq8cb6STptdKr8cX7qK8dxfctGKAiwIy6+Pi573V2VAWQMP5H8phrm
ZyAbWUjoRFxF2r09YN14a20YooMXlQcSBcRNkfKaXRG1UORCRgPKe6cnmh/LgbHI
ehs/WhP3vutIjkSvSQPwxI+uL7+fno4QGs9n9lQhrFhqSJzrbgjtCYQlBxHWzZRg
IWM9v2mn/iT3fNdmkOLzZnm+txL5XiFtOKAwcKCknSAsM8ssjpqpfHfQZethAE96
Km5w3c4n0jtvz2UfoegEryfd7sGsN+asOhkW+KDir3RcvIPr80IggOHsyus5yZLs
VUgE4dI+lWqLAnT2D3BZP5BhOJY9yUK5Br/2dippfvmKGSvuLhTX1Cm2TTZeWYKd
IvUTOAyYJbuG9RHNJ0fCSS86m5x+qCwZWDcY4Upwo/fqhZriXm9gSV2UYjDEb0NV
UDQJjnPoYK1gROaAPO9l5ycHs8+Yw2tSh9vhTm9eXk/3xtschsaVAOZmhDG6m+ud
ifgJ76UqDWojl9/GRi6M8FyrXSaGEAUAgG1lhbNM47xNKUECuJHtIBPtYA3mTNP2
IHHtExbUG7ehafafYdRoCIHMQ07snyeMJrVoKA3vj15M4Kr2d0Uz17KPPvnQ5tCh
kfMaL6oO2H1j23YiVgK9FyqAv8nhrHCi3J2Fhj/Y5AnlJZihdRXS7fMRtxbvDqzO
KKtWhmxBEHjUlztxb4BACAWcvIvcsomXjptAVea2Pi4BSGWFK4N3Q8FP0TnATRkT
DcHcgGP0WeUXUlw2uG7Hut2q8TjwTJaXe8DJ52eCZaEXUCu2mEAvK+/rvVQ4feT/
HxXlXsoOnVNwmT0f00D5lDY/S4+bgTr+dps3Nl5liTRe8+8f01KibiLGPz0TyAtZ
2pzP9b2I2CtGeJV/o8tq3M04JwcLJmwWzoqdNl7YROjpYlZy3x9ruLyGc7A5v8On
XGdfmJIgSz/8zoLuh4Wtv3P1uh0xkLvD2kihFxHA2pf2UvIoJ6U8Ax9+a/Gcd8Kb
s0uMMeTlMTE4mWpT00RY+1W9zxDWGMXzEr1tFlAFr97R273xe1hRGuXZBnLaYhQc
6UXbfPsetVKmJYAq/q/rBWob9UifOgUKVmqxe1pbgvHgrMY5zkOXLdyzCAFMsvfK
b1zCNt8IFR75/8kd5+FTRtQ3S3mVNKsdOCERo1YCX30HOD/8EoY3B8la+5hjFLuu
hX1Qcw4U0EngAixEO02+pgo5BuaRGsA6OAMVwmRWyOxnRwyr+x0WtlsuHbXIngrd
FhyPmOfAwJYrdrbY4XsKz2LDbUl/0XiRnc0eT8DluKSYlX2VE9rpQBxwem+KECYD
lU3vGGGq4XVbb/qT19PxT9fFAuYvc6r7gSUbMbfYVCwTotru35C0RpKaRvELZpMh
wqDX7K3kQaisUeJaG/gmTDto9RFiZO8rffcka7as4Ni+Az+BQ80MFgK++cds51JL
B9I2lCULGkfbU5HtQGtDgmn8/4jNmqnIqwEyFTRMm5H88aLPkt8xEK+9TB7qKlfd
9q3qDDWLdLwiBpysf3bmff/YRLNJQnU/WH0ROqdOuTEy4oMHRp4cpljNw9Pl81qH
bi0c8F9XMJl0FGv3dOImK17bbwiTvX2PiMJ3cGBk8bgohoyGXSgmL3x4Lba9xWDn
mIaNu08qw/s94fUzY8yxQPpsLwXeuzXJ1q9P+iztDJueQ5OuVWsFx89i+MTOnWkT
ZrMKh25KW2l6iYozPNsrj8sNFfeL4sKiExxPop08HuP1g7isNyL8/EDmP1/ObGqT
zNDUe6lureq3Sxth52G8XqB2zzy6rfjGnCN08QIYyInPkl80mtBCJh17mA9Kka68
NCUUWEHES0TtOj/KGi3J8m1HIPE06TXZtL7WCq3RQJbOWxC1rUlPS/fHUYLMaUEq
NADguv3lflledg7bhn/r2fO64Ip9YkO5JH8y2w2cne2m+Uym6FANc42UQEJNGByJ
nk6rQSaIsoZP+1Z6ILHU9SV2HERYY+AXBNsn9GgjjGXOb8wbeXMNUXQkmi0dms0A
oP5LD9Km4lKpHOoBj4Qn7MrkdYkENeKlQIPp/Z2Q/XWTms3t9mz7mjkqQEPLVmBK
omjsOWgdMAKUC+k2wjtFnyrRYLnr9cdtH4/aVWAIZKdtrYBXdesOVRCm+vOqCHox
37+cH5eWCi4ihWf5PGtJ7aiX7xfyhvMUVD6RoHIrNAT9cTd5SrsacZRQ0bUFPjoI
N8Lj3/CaCgx+U/4euqPB8RCBzW1kfuX82bRGeH8o6D5xE74FnKjLFbtDf+6jpmC0
b5ikjcqUYkG+TKbZv/VAb6dDJJ/izEqBRX3y2yIjKHfIPT6JWsh9XV5yX2eAopN+
wcliHZ0IBHcWVOKGgXVGZerEKPXO+AeZk3JLDabLzqmqaK5Le/CapeDP1UMGaqNd
TLnikOV88FdeLqhnHGdhfnCxeXxdA5+9b+NCvs0V9oZajt4N0JT1M1mXEGWkPly6
DyYLYNV9ta/v7v7v3nuqdrp10ur6e494/TYVh0ueqvvyWBMZ+gZBPmtZ45MMr2vf
7JzwPrRu48cmv6X9Gsu8XjB+J3QF913VYAL2Qus7DyNp373bVEXo25DUe81fRXTF
Tc4jXq7Da9w9NCt6/X2K3jDn56iu2sOrxtvlV8FCnbI5PMmw79DnjByOM96igAYc
tDr8cZs3nGNTGri8W/gzKjbxTEjTF+d2IOAv1P5iRCU+n47hGgso+H41ABupZ2lS
6Xw+fMAErigxRFx79FTJ1tgyg4vkrAeSq2pOGNefnybN5PD4cyjFWRWhMRrk45C8
m5257Z53yj0t7UYnq6VCibnaUJVc96tH/wbhQXWTfW8olgFU7yByHGtVf9WXgJb1
BUe+/8OpcumdOoLqs0hluEXYv0pXfvPaN1fU6tvtODIwBooJnwZxtE9liN8Paf2h
bnwZogp+zlrpL3+DakOJvu0woCcgYgMI2iTsHmYE2wE8Gfy0/zWDNNnbvCb4sq8x
ox3W1/3SSbMyXpiNzt/vZoZ8+C+rWvfaeVMRd++hiShBskodttuVJxUNKf87uC1R
RjCof86wHU+Wq5L6nZyg2yDKonCiRCUWTaOiTnhQY0aQ4Xa9rm3OFUMUyK6En9tk
ZiQcDnHzJZKrOeUF+Yk/G6sgzpKCC6KVOML0AMlg7D9nmUjdj5jx3bPIdhmByk9C
V8Dr5rVct6hSoF3kpjMRqDzbuJVZb5fIP6+ry3cY9BArHdCYw3Ci2WDCEfxMWg8E
LDBxkMq1Qnj8QdoUVkREQQEoJMNGulEnCOf3iW5dYxArHKHUh9PQq6Psvi76yFnV
g3P/6ggdzZlqu74od53SNcqO5EH2ZriwYI2KjB5YuWCeqmjQux7LNctZmxm7NE20
0MMtsNqPmY7U5euEXkgd2tsn3t1OxFAbzUneHnVS6iOhYq6fCJXH9sXkHdhJGVFb
Bs/PXC7wXwn6I1QgEpjWnLxZCvcll41e1ZNzvyAAk78q5gx56JK8Nu7sNat476k5
5WacJkJaqNDmg/R5cnFJqIVtZW5Xqx9ZU09SRhb/iMWrjqriUWnsp7oKWiQ5k8SA
gRlFvvmgbWc/u3QWy1nSVpAV42ZYxpiotpTPkuImjoEsE6qjZXTChoNolo0AAvqs
lV9h70VWYoRyjB6LKiGWOnTEOrG6HbP6Ek93nj9rf0gGXKZbbPQo2bRRk7B4p2a6
MX/Jk2LfekAUwkTmvaZvzLaAcVJPmJx8+pablSgh9+Mf6lRIqT02aYdH1T1gtbXT
5LFuterpdgAHBwwkijb2D5q3uKXcU/QTRG1pwvOQ1rM0Mm4IA7tML2exQNZecV0m
s90vDxFCaZ47LcEGbhcEdIownWEigJdhpHzdijfd83Yb2zcGDM8X5ueBGze3NAkK
URVJGd5FqfFFmXxYX4vlR0nZ47iKEpb3fHv5pE2otb5R91gMdqutesNGPEsQeeDg
TQOXuFSBr/SyUwHsNx0O0JjlLj0DNrKw1QTCJHyTTpOmozRuqaM+udFknJuiZWoV
yQ8dn9s5gh2AUDbMmBgOYcnCtK3Ra4kA75q1FfO66b7xreDZckhfNACYcKkfC2wp
MvW5SsCEyAW1wqQttyr69SJYnMm1iwg6doXGaF9cOzFLetWs9wi9HP11MPL+4UpJ
EG6ExPy8R3C500pC4D5RkuCxXUS25euvlcPr2Guq1N1mkYftqIDimBhFYvsht25H
9sCiGRiEDVQ0tBcZa9U63Oyw/cyVpPbhZ5xBh1gp9iXjOi8F50DHMD0qrIMQlsA2
ZrAglC2bL3E0bczjjj1Hx+wLclwD8y+tCy2vo3k5Qf9D1wdvxl5OU8onKY/ev5UL
KvAp+wFB4sLAKqvvUmQAYzEONK4qOoVyTWHPDg2WRvorFy7nxulaTdT6z9wToEE/
vW8/kjV0nfDPxzo3j4EUqM3uoiW0alHS/ydtzyYgW/v0PBL5fT6nusRDDReVpACn
WeWv1rq72bhBQEv3Gk2TZ2QJiRFqGW0LYY8d5HuT2l15qvHqVC5Q+OxCzlYYtDSp
lT7Y0eC2Yn/LtZPmYbNmB9jvUldxiElvgowHqNazf7/ydNQwbak5ORdRpyOX/WsP
1XYG00F4IBhNulbW0lf8bribVzz+nkTVSQJvpzUPR/hpEiimlHBdQl/yZITP9XBW
e13a2xxEogst1F+48ZaU3A23EaPu/wQh75HnaHUySivpbIjOS8U3HmxXzyAKoMwf
vN5pnidukWmPesiYrQpmFWI+aQv4qSnAtdCI5+sFrBkLuP4JItmJLZkiw9e7O1bz
zZ9e7dx4KM4Z6hi/TXprxXWN/m6bcPJhabqB3vGLZZT+cJjemb7UeZrUjJJL9o0I
BnrJmMU4dDfpB7Qm9FWNELl+Pn10YFQ6/lb7aQ0N/yVRYg/nhhTspwYJX4Zy99lv
gFa0OUBdzSm0sJ9sKaR7Sb9rM6xRIVAa/Inov29F+XgJRL+g2dCtEbAFtmsbkzuV
S+3aVYj34IS4SyTp/ywrnCsmdhqMgO2UNAETnCe1S0+oAW7iPl6BmT6trUUCNvwB
MoF0oW/9LmpBFqwI5LXe2rq5UBu04iLNpeXcF0ICD2xnuzcq1UJP2lx8228e+l02
iFgoCJ6FTAXx8v+MlL2GC7qf5GPjgl8CS+D3LAFCYciIwR0/zt15tUGGxdZbnS0W
xzA1wytcpqkpZbH06ZoRsnz5t93J7yCbn5mPr8LQn+K+KG+z5Uhq7oYJRKXGlcFp
Mb8/OjLS5kt2qSImFgkQB5OguQ+UibninoQPkABeMSRPyYPoKeJOk/e01iA/GZ1r
gjg2TTA4xG0aGbCr36XgxzbiCfLWkWS+PafS9tzjzd9oaA7dDfd/ChlrUeyO6T+c
Jg5bYNG+wlJsHslodKSapxkiT5yzvZgxy6jR6uDFVCrbuj6QvFf99hdP6Rx4RsWx
QrJuirNZcoEFd28f4QGt7tQqNfts6RkwOlMQguK66vhNZoksafsHIVlMHtippsUw
ALgz2qAVPSdg7b3oH8vNje57BsXCoIVHYfiAuueeqcOzfCnETNk+OVVwHBFLnzE2
I0OEKVp8j01Fk73fSBz89qlQSoS55IU0iY0I6KJvn88Qihs9nPgnCpvBsQGp9Vt/
Jk8KkLoTXIdQ5twVu0hczmXD4ZTpxao1LUsbcknNA/hJhBooNFrlGzAptDWbulS+
IyP9GsKKQQo5II3nz8UxLjl6x2ZtoyCBpWj3Z5YpSUX5mpVlgdjJJkKjKfpzKke5
W2JvsPYWc5ZOWp7et4LGhUEshjQrJUCJx1SQTrzEB95JRd5/rPRtag/2SsZvFXrV
z9zhIn9bAL9o5pLwajlbQOIiv+rH3xwh9WvdTxZaXsq3o6W8VQS2M+yQoOd+H3De
YcKOPjA4ThM/U+6NIADqXuv2xd+W0/QuC4VrxlOQcRMYNqIcThBfBAkKMe7QQV7s
Mu7r4OrGfx4sTW3l9zHx1lch+wJ9lefG9YUqe69+THozCkkqEnikjUULjmX+YahE
VKFBT/uMRHHntkrJzSMExE4baqjt9nTpadyyNqnav7z7DB8CqEikfoI+i6qzxzAs
AB0YHGHeG6WhgaOoimRvhLlgGb6TV0ocxxj+Ox/ZlzFtPLSiigC3M8hJD+mEp+uv
5wjcpwwI617aqsAKUOxW/oOnPUm/mXmPRY1sSP/vRCEuUp90hfGNZdLyZLnJG/9b
TEv/Czy9bwuveYIlOnXVq19zfiEPTQk8VnzuepHprgj76SeJdYY5qJ9SVpzwZSh+
JH1u8EfVaRrYf7XJZvWdxUysqxMzexKRcTlldYilP9XJnv6bVrN0zJfhgYai0RI0
LWRvxGhsPo86cbE8ExTRFJqv+DnYSS7k9zPp4+dM26UeKIF5kAOge87KgAv5AqDp
vTrAYIZydzXyCJFAioy2baI39BjuP5hibUqn3db80ivWDys8+/Qz8SM0no8o82NM
RyjMvV8bRmW+An/uYoSodofxVfY0b+9RueKMDD23SlqBKQON8t8mj22mExMSzpT5
zG9agEdqUcD3h5B5H3fB7s57/r17u599GsHyyU444P6VcqS1PFYRjEeUfVhlzfgd
SpjjA/VdQ8OXRsgEASgalrnJ92IZVOuucGeb6Q80swgh0D8Nyl88vlhoKAHdgE7p
1N4G8drLJP5KyITE3KqjGiK6VAup93RCbK8VPvpkVk+p2Uih648xWBJs2MxI9/kM
zHA+YRlXHxVWGfldSSKKpUJ0P1E97/JZMuisnqyt/0QqUZpQPeOATaqPpo83bFe6
ob0UmEQx2JYV/REmgiDn8n6XUCos+cMzdyEcVUXSYCvhLBFsCWr5CGxYF0gSwlXi
CDBuLgcLQ+xKu68IUAMiy13naChgZ0+XzLsmqZekwP4DfvMoB4tloL1cwbtimEoc
B4SjlkIeAPWSI1riDuAqKVt6vWozvEZE2TfOCFYwBrHyfW6FY5jsZpWXlTznQEOF
lpbw1pT0gL5vc9WcgCADjJovwb0K11n7XJiykjvYTh/pmUwtRdD5dA7H7PvrrsCP
bDvUGwEPaivnrQF1nPxH7AknF7LcEEf3uRpHaC5lec5WKersmnanYmYrzCxb/ej9
6gEwGwvtyTzlq6Cymt7GjTrah0PhQNtZVCvt8rdBfZfPnoT/ntzutC+fCz5due9A
FWITEMkOaXl5++jRX3snLUfy4QJoGwZ1qLLOj9WjLa3lGwSj3nd0do13K3eCaEE4
pZbK0zxNOX+2AmMxSYSXOswmgnrLQ0fn+cRr6wsI6i2vQqSpcOR++QgwqnFboYtG
JEARtWwsu36NS6rx9VUngH7v5cge63A5JFKAbSUUh5G5FVoHtgzK5JFh73S1I45q
N5z/sBjbhzNbjBw7SKUvvTVAcWW7QPwQVsw/U4WBe2/Wak36h+e6ebb6J3ES2RE6
eIErA+YPkg+ySbr6jraXi9+NerA78z5sWzXWRyiUccQ5nne6rJq/cguS7XrZ51zt
Q9YAQNd2kSjY+6pkIHMPBwiP4WYzAplo/AZgQGXwm598HGjUNuOeH3GMwlkiHUvG
MGaWy82TdlHCLD06y7x/hAdqp65nnTEv7BsHruNZblJPeu0suxq13yAFAKaCghX7
7UAZLGB44Fv5a+oz/0Lq8NU3qZb2glnIzFthK83baSEtpA8tIkv1jHlfv9DsQ2UW
4J690cu3NKMxlSLfMZqakD1Qdvl8jftigxdXFVXWQC+IdRXX9hKbye9yq6/m14cc
IkjKN1l6Ly74HIqkKdP4k/rezb6nOWpo1/MlYKWNmXld5/rmFJE8J+l0gd29kj2N
eX3iWQUH97LdE1VCGZtWHDmf26A3KNjdtkDqfVtI0CHdSP13Hc9IQIKKEG75Enkp
dgaf0iV1is+cO3WVqBqE4s6kwZFJn9TbY5QbS0U7r+e4N2p++WfJ1tCbIEB8z8Vm
pxqImNBlCcAH7TjtjJ2GsMMWPN91F1te1ONKxnIhsJjc527iRSOkaQD2cTdNmERe
5VBOeS2s42kww6KkhdKHyshewi0fwzHMI7cbSQLgjDbP0zx+YmZEHAVQoBrnRDLC
SwyAo8gSyuFw+Fi55VzxmeD2wc16JNV6nhee5U+ldyd2S0r0JExeCABSV1wP/JyW
iAID3sIN8cQyOIXZvULfQ9LqDIz8iLUXHzg1+HI7E3x61vFYXlrIIyBi/FBYzVBx
kCUkMXJJudlRGbyksQCDbmEKLJ+wugwz8x5cniv7qCwROo3sEbEHmbp473TA8tb3
ZfpBxwdGIKxwlFQxq0nZDz7x3dkNaqPOFvsL4+EA39Q7KeIUdAsqCjycARQJXeH4
d29qX2N88rvYNKCm1KFtMtyjF1nA6Gzsuh4gccxm649g3rW3bS+rXX691c2/x4m/
ezZLPGpLF9CWKlJuKL+77ZMjNWVzBWGn9V7HgK6n9FgNTfYgPK2JtU5Me6IbcIm4
Whr0/ENKeWQKKpHQkHnQ5eHUwm2IxMA1SKiy66DJOjbJSTJDuFAaHNEn/lpY1mK2
ul0r5NViDttdMCCaSDvtpqgmpctkEXJ5D/k7TNGUFCpQag3NxwM8F0p60aDRVmhv
XAsTliVYrd367n7W4L+CFQ9ltqz6LQAfqbQLpwJoAng1gWRwe5GiHKEfVV3CXt7s
GTKwYM3hbsrsAV+kyzlbXQ8vXs+EBQ3N2BCctL8eai0HV/vzw+m9HJ3E5BLJJU5J
43j0nR6elO6YurDgAkQGYRJwZf/NoEw5D2/KcUL/5TIs6DmXDjMjweYZAVeaIIiY
coH/t8NU36GzdWXioXB0dZRi59HPm8ueoZmnMHQWEF+cRYB45DASUTPQzjhkNQrB
wcxRnYFtdZ6ezIm29Ap08YSSfc4zWEmn+isk+50273vQZuMDXuS/N3m8f4eyZQQe
r7uwoQlxxsIAH1x6LX3NflkvuwyNTNkKWsPHsin+pnW62Uk3Mz2SausNWZ0ECkeo
9zOPAJMlrC4lEsg/ZHtydEZ0jfVuwREr+CyfeGzi+xNKnTXUw/gFwc7sRrzq5yJz
ZAJqBqAVIHmAJkVgB2xgGoN7lJ4rNgDYyGAOptaWg3j5V8PLtPm2zXlANyAG/aWI
At+RzNerypzWAR6KwT1KAkVPERZ3a5sWzU87D4KHl/YlVl2SqLADngKben73DK8F
jDwi2SPRzOL6SkPWHbYUeKfv/IAk1lixenQwXsknc/JUnIMyzflSVzPdZyuVGZuV
fe48EUP1nz341/MtOt+MsHpqt5Tz1HVn84dt/7RFItqgWezOM8huzX+jVDGpJxzJ
MOekpj+KosbE3Xrmo9FglnQf8U+oPLuH54QgxvQkFz+AFbFO7Q2rIa2RZdAr8d2Q
n61JY/0B8KcQ8b2/8rTreiMbmrrUCpM9QGHTALZ6/iw3GrA2bkVcOzz0kUepPIb9
ZjRBlr7hz8p0P/s6jACQhavD1Ga8sqhulCzrXmBX6GXsi1L3osExzUK7xcbm9KXO
GF+PrtOqOC1iLFP4BPnOZXdqeYZli4+ezOa/LvxebNoUaebxVi19hnEYdnUMs6sB
v4EjUjlMLOvSJrPAwA0nrU61+UU5TFvVf3sneWLOcWODQJ9h5GT2VNGQ/Z2tMjtl
v+9kOKCX53pZUc9PjNU6xUSxHzNKYkqgKKxY0rj9Y1mZKQpSZFi9QGO25h53Fk7M
hCp4WCf+hpgKfaaYYaad+ORzXpyvmvRuC6CdSX0qf2VkxLPb6UQPRyFBGAfwLogl
F2s57hxEFOkAx+zYFV3/Aq8W5IDASA3QEWyhMF4+LM/O2GW9l0fq9lpovlbSdGEj
3DAavI+2JBfVZLgSsK0JWp/I/AQzLVW2Di/6gz7+5jl5evYbmW7HZ/qYYueZ7rou
Xfybg2/34eXrV+1J5nEsj9KRNIJqRkZ0UKRYXq8m28PfGmyTkPmYdFiQum+1boO7
3R9o8Q+sH9GCA1NHeNkHbCF6fNvbetBxU3VZvTGANISYl+etT/EZI9O2D9eKAhcj
oBHkcjIaI5Y7lyZO4xaShhaFTFLwHhq9wHreQTn9bdhZHUG36QAYGeGAKXbDR2dO
JWmly1C7lmwwDQTwttfZQ3dvzMqUGlI64CyxCCyceE7SmK/yzFXCiZay9aIsr68h
bMqnOsGNC7aJ/5HjCqpjSaofnmATxuUtP9SvaUa+AeKLjCY3xjQYkBqRd2qb5cQz
Z4d1ouqgXuzQgwlPeFzYkNi9SIozfU/oe06Z9E+uLGwOEQUsn5ighfUaPAabIfcx
LPMnTpd0j/2QB+C25shUpz32tdRyL/TMLB5owwBXaJ/2gwsTw06cgN0o0viiZSXA
YqAEOrS9nFdlm6gk+tMJDUMFEaS6jLAiEKVIFja+05dAt21vrexD1ojZmfknuMBA
+a6zCLbNh98i3LC4OA3UUeRLQPi1aFaLNIr+95jf90/YanjCfCHQLJ8755Jnkweh
U0TZdfL4OicIPMZYnlUJilxRqJoV5/ApU82U+HG899G2T7FApYbC1PmAiSt2bUYT
oIrs1i91frIZqUilhHygnEt8pCE/xA8XQx4jmF9L37ypfUPxfHJazKhbplR98qAe
8QoMkG1noaBOI+6dnTh228Z0RJSiq7gp03GBm1s3rqYL3l2ywNNeHBFzECndu9NF
eiQew1b3Dk5mDG5C9PYdDP9crTvt2bUXUF028QfaDsNydcpJsBNGyu2uh38dTIHx
kn5n1v86+WPDH6vNiNglTlIgOiQD8s6yIyW3iDXxF573+xVy+/h+FWkxMc77tciQ
wLpvrRjHn/CwLdGtpTksEY94b2HZMyiVScf+CjDZ/6lbOGcGEZCMrVzPf0rTfOfm
m24tGDqJs0kzh7r6yYbAYl7/EXefYvyRovQlbvJo/BcWmwoG7ujhb8BSqZqAeRZe
Pr0der9VhCYYpSCBh6/naLnASowGhOotJaK5kJunmBtXGt29uTT3G3G9Tc6JUKSh
K7dHp5Px7KvacDBfd6i1egUw8HsnGOrQAPlmHg52tT86dWkOTxhnZXVnGCsTCIFy
xMpWlVoWBXPDzDAmNiT7NsdO/OntuUKtgqtX/xTOftGnvl5p9lSb6WMUNlQ0w3TG
t5CSdMbYUKPtiPeEOQ+rVB0fnuXGRpvP4kziQyIm5X50wQP1RrBZLFYPUXjg++Dj
iEYg8tvNhQaiekjiaHl1sHmlqOr/4Yon9lHbJgQhGTurwikxl1O3t6GUifa/A6lj
owX/kVHgAWSUwKYkuBdq2OUMvJuSv/sW+y7c3h9x8bLjk9KI8zBIQ/wZZzgDNPuM
xMn4sACNjKR70fMnyHxW4EwaigVHVGOHquEO6hMX/GxbMLHRatDbpidJVo8VDGIQ
CkGo61u4+UKzfSots9nIhLe7KmzqhwVNzvQmhWZkU+xv4tzQUIh6TdrTXjBl0eCF
5Os1uwHanmEGlhM4+KJU4nD44uD5UOhTmLIkO34sBgcfq7EOnAZZT5+9IMkumUUF
1CfglxQXKNOXWO6MuweEQC43yM+9MQg7TVa224zum1C1VvsPl14AXYeYyn3I1iGO
LxbnCEVviq46lm8uY+5me8pTIpZMl2xBlYIv/nrvRVY3LiCuex8hLANCo47apVyH
AhuyRhAEbEs0sQiwCo1u/vhaffytnrp24+i6cr8MRKnED0bBZC3iCSXUcCbsJMjy
phSwkjljVoVrOilfUdcjObbK2WfRv1mxc5dPDvbl8ZGd4pXXeyvZ9tUBfJpmifJg
XQMSh+FkhSd3ZzsyxqEfTqbkSDzfRHMfdQAm50S53QSkH1itvuiz9u2ls0sen1/H
CzFmIGHjr3tEHEG1NTOyUAOOiDO2C7f9Phz4AX9p9M4NDWi4Fp1LD3/pCGrj+GWG
XOFxUOwIFigjqGhzYC8yQSzhnokAnG5J3xfA5lNPGHOp04lBqzAeThtBqjsFT4tx
XRLD5eE19F/1Pa5pP3mpTEtZotacS73LFonZ8HppSU0A+rjySGOdNZ20vRFRFoW8
4UFTejBacecaMhSBZO83vS/FHSFLZWsXVwGRvl18P0+oJUa1+UEBtsvXqVLzyMIn
2QiY1dhD/no8O3kYDNmSTX45VOVpTBaqvOnR1rjiBnsIWOwVOLAxNP85ksNvnka8
nzWVCjnjPyW7bj7av0W8SD2wXzmIvNn6stfsfinmFCyFzZ69grFtDsAuKyg3PI1P
F9p1YKDTh6zt5zb2B7cAfpcoFU2mR4asJ5xQNQZYbQzwPY6VxfoZYYOs6tYYYFVa
3cMqaWTwD+hDoyMj9Zb3nSAtmzjTkTHey7bGfFeCMMfz3PHVu/0IZgpolwSJI+la
q8m0KqVsk+SSSUg6sn/M24y/I7LybFFabp3e2txMyXaoT3gevmuQKjIS1FmBMIyv
56KjEOiKtkJOS2Lq5GDHZWLGAJw5PIx/dczUFksrXXW2LXsyF9+Fodx4v1fto9Kv
tSopvU79YlwKXjPXHxKCJIulSmI7mSVdnf6/HGPjfklLOqrdRKrY6SxScBmZ1Ixk
XnIW7TXj6Pa+/PaRyWy7K9freL01aXzOp9yo06f0+HRG2C26nsu/MzTIwULUuKEU
KVX8mNzN0T3suAW+a259qHjZQ9zILK/+RWE5gvpdO5pQGenZFrJ5ECjWmwBb/U67
hvMUKePbLMioCDaWJJKjfZeZzd9GOX1jpKjvUlUEiSv9or1DHug+ExuetM0EnavR
MfhaBWL6Sl5LvFVU8EBISRJmdZokzyjSImUB8es13rfsoZxBHlxlaXQGRMdWMhEg
RQtxacpXiwphj1xrMjUdKtMg5n3QQ4zMuwqCVQLMBmyss0i1kNer0J6ax2kLCVag
0T84LJ789Arc5tBE9NnL4Y1bvhEDmlasa0E2LF0eyMwWQk4ESiboyTdBd1MDLY4B
glc6shtx8s9jDz3WFehzx+uhOXAfiO5HH8OrsLGJzr3w4uiNlKySG8tZBHR6xvCq
9sSq/DH2vQ0RyDt5T6zDuwQGxAW1MZ8TDVeh/9EARtTTV/+P0VT7LD89Zhu5fEEx
bX3KaSS+QysDYBkwxOLS3yEsZfbzOLdFh8kHRq4s9kjEdonmES/ynj20gl3V1X29
OWbgMLmos6MRLencCIQY8MKD4TNWSm71ViKkHWlUqppysUBzi4V9u9z2S0SkIaXG
OZbiug2Pm7lSPgdnqngpFP8cWJEiGm5Qjd56mfpa01Q6Xu4d3fimHETglcXmVIuq
y/muaDoyusvzOHnMhvMgpDIeL8QhCFBiu7Wg2FD2QnRzNfuel/HKmvvsQbneHsXT
jn3myNV3mleEpXYgOxSV39Nsh5RuNCKz9hgmp4ihl3vAYwALjVHH3fhqdzSX1xp9
A0HDvn1AjOeMN/6tSGQpIDJAOoksb7Q6PhH8C3/Y3bdu3ETYLiOoDSOIc+nd7+zO
yqBognqk7hWwvHDkxHD4oLwzcTWqEycEvInDFARQiEmoQLM3zcsmt8nA8EgIcMyh
TuGVY2ozfQJ0FOMFLsLBYnUYl0gpsq9LCuvKCQAsAvYxvtxQtj45WqeAg34sMvyV
qoUZFJ7d96R4DEDjlR+A7N/XlXPbQCBHmdbmrkdjikbJnMFd4iycT0sKnxrQ+KXQ
XDLWxiXFPd1YDdjgwa3DFfjzVg7UB9yfXu372jWcfsgvcjaJg9v/9hc2GyWICrqI
DKWfm19SAF4TIXFueRGE7DJgzXudDIKBnBDaOqvkfAYrRhG884mjl7Gzr1eCrM/0
51TCbvKA7WKRR8+0qV0NXQcbGuqDI/DVaMeW38j8Dp9g3l0a7fHtwpUAAM/cWDwr
OC0t2znfg8qqNG7bZA3b7NGb9/X/5DSbgwVGJ1pYzJIOyaX384BTGFjYlghOhA8G
yiiFrBE+HrC7Kk+0swwtABf0uNFsLKiYbcYElNwTHM9A+KjQyoadRv16Xsc/pp/F
MV5X5WMQMl34/imV84v/eil2RVrkZE+Iv3u6mLw9VioF+NGZsh9j7iH11zr/TIkF
v5Yd9p3rcpukCTJIn7wCGT8kcfwp1teRrmzHh5SdqLl7sjrmrX1qs23XdiFoDW+R
cLo4iDMSKawCMN+B0Fki4CU+LWhfU7F5YeqJ67EbyAgE9IpLcfwz4qL4duNuaPW9
vznEt3ufmhUNb/a/DLqQ6pHQYTuA2UDSkivkOnY3DWuCJqyFYAGzJU7uv6zUsvYy
cdlWAVfNn1wRO6dHc4KtEakT9fnpt2naijJUfZoLJZO9+KMmwvt1LNUI9V2as3PF
tzEE2X/VVgDQ55tOMS3eKnurX5Be9EF5VvVsbYsbSfGPLWzp0WyjCM8Nv9rFjD/E
UcOewwQM646FeXqAm+1TVWjYGB+IAK29aRGYQA3oD7NtvTMJIcOyG/hbhmtDka43
qEkMIuiWl0w958YsBywCVsE7yFc5iz618fV9D0XZo9eoXxizTIa3afVz1ytOKHsW
KlswA32bJbafxHownQoLnwdbuboVc4QqQ/GsRJLV/rfZssE/J8g1Yg0dqXG7WmqK
XZuPwC3oEbA3+FyDETWIPMc17Sk9rD0rQqoejwzsscI/3UAAwO1J7PmLOFlNt7x3
cGd1fO0y8TqYmjrZGEoqcGK/IoUPN5ab9AjW4B0r4XTCsTavFXdy8Wb5fOzZdauy
6CdBtFgi5GBjGfYMaJW86OToaHzhuBBYAAHM6xWe3Dv5tBrPmE0uw7rgzdBQMky4
Okh0DSTA1wU/O4zK4BRchfhpeGNmu5+bE1lSYs16aKfTSsKdszBa/hRtcRzbdOiP
6JsLYHQqv3sks+4EnwL1gfSimYrZK5stWgOqEhTgZz9NMx5aZPHfNt2dmxVOY/Wn
wOO5FJcKlGB9KOaPeCmR0kxEj2Fy2PCTWWOsINc2ZKIXGrJnJSBfD7nKaqbpfKcQ
oCUDvxJ0MAjwisIdlQRwh5i+vGkhtVQeeeNaIXJia+U6rSJAvemw8/ylNRP6dWBk
YBMYQyN+xQqxypn9XjBJiY/1TqSPhRRA61kIihz6tLc8U/sz8Q6Jsg3bCB51TBIZ
+NBhOPpoR9oKnMBlSF4SZQhhXiNppEuJGpC0i2V2G4rPehyXHNUhFgJZJqd/oN3e
U2O1k+D/EfODEwgxSN5IWcF8QihqKSWhmRytV4Kx3CWSzpu/5PVNrY28lKtinDci
vftb3MDa4SPjQR6ub1zJKqdWJKluZk4/gav0YT+meoiBonuEhHNXeTuN71+upAs5
jC8anSkHLBUvnxrd9gE4lVroUbw5OWLguBKSQIR5OuNIgkJoSfZh+G3bw6GmokcH
8M0KBPD4R0OgfzygjArpNOAu2IfEZvT+dejjWDvw1iBXEarVGJKq5gRSBca9OjRO
5nzSMZQ1fnT3FXb0nhkEgNWB2mrrp4wJ+hICuS8ukxQlVKKrrw5IycLcFfuF2jzC
KM6N2wEywMnSebM/N0xy7WQocfeBcsQ27x+loA0q0KPhdpYrqX5P5Z+Ksn+qSE4V
BYjxskRUlXt2IJa0gSh8oW/VxeUqkqpVvWhU7qi7RoU4t+yYNBZnvcCMJZWV7yj5
LEK+ELhbOgogFwO0bqwkpKqM7aVkA9uFGvbjalPTLEscm0m3kCj21/6czpVjWTju
qXOsvbpHVt93LH5UYSWgZUdJ2ztKO2OjnyOq4KXRIJ65qKSfr0XTjDNsi9GqaNyx
Mp866/v8D+wyveoyUhMwf2SPTP45y+5shUrFYe5hYE9T/u5OIAhkfBJ4GFKxyJ2/
fIl5eAtXzYBSEMuYrpsV9z98OcZ2bIsEa/M8at0iXbzLuVImPW0Z8Hnxaux7/k5Q
s/ib8Tas/jAihkvCcoyZWtNcRMI74KQaTR9WJxBJtAOSacJQeb8O6DxbRsDyvo18
Eedd2skd2dkFk9nult1cU54DKdbf7k3w5pKX1ET9HdBAjN5PFEO+yWhEpPIA8sV2
Bt5v72AgMChgunYl6SAl0GSkr7v7DLGCkFMVqTR06s3Q1OzmiIW431inuc6d9dcq
0PNG/3jtIsM/E43p1IXd66haGURWOvDpsHQE/2IwV1ywt7jBpToJ0+JHjmIUtFB9
ZaSjfcf7U/HfOzfJCyuwZszz55SaUHf4HbAIczkVCMHoDAZ92HdDfQoVYPmY0l62
00VnGsIwE70Uvc+xryl2mdui1v1OrwsNsGC9pUJtX/X+JGIl+6tQCYeiIutF6iJ7
+YCmDNvWuCac05W6KSEqlIygfsE/nuCsk0y+kX5cnHuvl2IcKT7kvacCR+aXPpht
Z4aegJQF6AGHQynycnWkNvhKQ36LoJMa3LiZ/okpxTy42rmxtpfeoG+zfocaVGiV
6RMgfrFvTG+TUSBLNs0SDXdxEQRnEF8yd6lfFDFwT5ULNpYC40BJRwCy/FH1gxAL
eObch57fvnf/yEfO34z30qWeTcZ+RBzufacxWaJUl5ypaah3LUC5Zz8C4s30NUSU
3grjjKMYjZn10xPWhGKPnUhUCRO0zIXPBnDC0/f0NPZup9n187Hjaw0neYy6HHzw
RWXE7eET0CyCtMxmzV7qsuIe86vjcqcy6DrShdwazPN/Mfz6yNCMm/eLmwaJsW+n
5jehf5d+/fd2oPnHuZ3s4cpwiEbrcVFfnEhOQDTiM8bzu54iYQ6iXn/UBqtTO0Qf
+Gc+ArDnS5w3KiqWO2GjwaUh8Rti4q+8+dCdw0mrIu3OzvR5fOgnAZYRGg4EhXwe
PeZAha9KWgf0Xoi3kGusnfa893hwSxUqfNQ6w/Nm92EDpqEJo4U79O+c0eGZUJjM
CrPBap2KvANsTC2qQ71LoarXOrA71+ceLcpIQ5S+G3kud7v10Bw1l+/vqC6hWxym
21SnXBnJ7G17cjtuy6uHPih4scf31GkHnTv2K+lAvmDf/enTRVbm0PBJam5qcquD
BgrG/3onz6e+p2kLugg02Z4SYMt4/bdh6Ab7m3CdXkRL1QZdPWvkaE7QfZuWtnLj
6n+NrIsIIabURCr+WBclgl5TbkEsHnP5JqbhlTY6ebrZ/GJKansvTM4Kws3XCcGt
iYqBkT8j4BUzeAjgbNqRFdNh1Ebj14H/PjY/U8FSkulpUTFqcOCryjuDWdhP8xiL
FuCS2iyhaMRXu/NrOZgqTGSW8PGm29a+Wll1NY1W514th4sRFk2QKE+F3zETOEUa
coV+l/fCH1RlUVUveU6cf2pXT9KrHi4dHCo+SIy1u21d3EVEZhXpr7DcGQk/4MhG
QZN08mMwK9qguSrtgPV0TWId/ekdagG/8SOWMdJTnt1E4YKD74c2JEQsxNb0zRBi
H5I9iRvmMittMmNJ3dEZyHrkZR4mx5+KnMK8EPc1abfurM0hP9H7vmYakmSdAj9Z
5lq4F34MlrJTwEoc0MKxsMr8bWpS8k0G7PQuG+lPPM4c8/qlq8CrgcgTOVtt5cLu
4BmD9PT023pG7f0s6hOQ8k820Qy0bS8ZDGKFS3YQwqT/kXDK3/Z8ttz6XWbmPXOI
ozKQfRjF7tALEH+/DVvc34ZVWNuiFBDfMMV5Inl+nrQGJcKT2CQ4A5j5UbvIR9jc
kQSEL6J2FuhoPMMT3fUEe9vUqjcmSCfiY3ul+Rt9zYz7rDTArMSTA97h4iGPZLeK
0Ij0R/2EBIj9YnMosx9tTchR5waZm1Ff3g3IEFlqS2xgWbISfjRQALdtw9jrOXUM
Mq/p3F0ixKy4fSPi+Yrzx6d36iNDUuzbGthcqNhNHbR01i/MwPyqqblc4ABTaJWT
VOFrObYIrF3CViVlzypWFHp6+Mu+7mqrz4NjpNVxuOszR9qSN2sKxpNuK6+D3+FO
jPVS7uCTrG8T/UrLzVL+kaMaC9SMw1wBeUova1e83Q2o/gL17wTHRnSzU8gY4pvD
Navim4G9JEiUHMX+35sujT3KRqXjoeiC2Quop38LOt5gWK0849YOUyz4/sOawZOB
EXF6VY24/kkF3PHyzNs+zFWGCuq+4QFWSwKlP4rlduLONN8SmfuuyNGjDS3Xk71x
9JVnY5jzmNyF/npvwMf3BKQSHzZu7fnjXWlcb92MNC95q3stzgo+ZkfH1sy4gJH6
uhQQgAARmzfIRBw0GLsPIXFozXx2PKiotiT0u/F9uUAIcji43jqdFiW/8nQlAnzz
E0WN32pm8PErLF6PEqohbgMytebo4SMMgqpLGTjQEWBRYCfX0GlA2e+vSCwVGKiw
KBJqs8lUhhawY80GxFQYL9o5JonPBOINftow5ti7ncEC4BUTn+74Vr0pXlw1qD21
9ZHCMV1mIwIu7C8MGKPi39pKFkfC2ZXYLVWWZaTP1t40nuIOZySbKoI+1RH9WRfV
8AYLQd5yiEioD1sCgxHfE08JcR9bUkV8nbcCthymDk5vPBwxtVHLUCnAG7AAeNYu
Sc1PXi7e4L89DgpweUFroJR4Pnc+0/Dpf0F8xnDC5FQk1DJ2zuKJFVLcwYZzgOts
gIg7k/00NGAiQIHJ4O0miaIWU+Tjn46JJU8G4gb8lBmXp3OwB9CAuDafYhJBsg9j
Z/floH1qz1sIixXTgcMzlHjF2DA+O+Ch1VC354RHY6hoCoefoLtRIbfmjs/ZmkN7
922gSaJzWyb6n92jt1EnvQ8bHRM4uHJs1ytJbAaCRlkWDVfJfiui01t5rgyL5AcS
vAzDFsqJr/Cfb5o05kwplDoO6DTd8emhT88QS18zdqri0t7rWLNAdbhngNveb8qY
XZC+VxpUtyl0AdS+W2geKXJ2VCb/ThJLQFSDxouaHQ5o+fG3IdgMcCMUGO/lZkkH
lhoygxGB8kEl3L8ZVhwQrGJLibKMDVvb7crXbvF3dSVLyrtQ5RJMqbwFn8V6i+YQ
eLc0gxQteHQypj4sKoQOE4nvLZ8QpT2etfhhjTcAtjFRARqusBQF8jOjY00ImOq4
ZN2y1a2EpHJgM7P5GW0+hvhhr7x8L9YiIhBauqx88y6YvKDm3MmqhD0gC+MoT3N0
RKTH1uDeuliOkdoFxbQC4WCMqEGktynNupbKNlapMCqT+E73eLOL08hpZe4H3tZE
GH2SZt4mvcNvZLUDFz6lHpxc8fd5qWIWN1/CG7bXTJtLPD57xSaJa3XYUGX50FGi
PCJbyatjwZC6SmeRW9u7ej10odP6L7Qegqbm1WWuWgbhA3kOhJD5MKHafdXhYT8y
FH6q3N5GPjbLA41SI5h6oU3uvsNY59NX7VHAe4C9rz4DhGHemGsKIimPvQQ81B/C
oUPfG+4tt3GKq7Z2/RczLQebKpes5F4K5tKIetGMTeRn34tqTbazQNwEsxuAEvuN
PmOht+2xpfHptdpdUKM9hT15rGjGVkuxBN+vkhdMVSLAoxbSXaqZUaKAj3uEJKvS
S+Muswa/tl5K/+bcgei0oXk4YVBr3s55MXWTsH1Y1HFwJ8RarWlpGgpKryk5jgjw
zj0GlZfFJDz3EdInYxkDri66WIxeDhPh/iCYTL8MqqFUgg90BhMZI5ifeYRY+xsz
26M0KxExJcBBCdoMUnhPvxQmDmRhSrhjv/obxQVSNYh92L81jKfTonLp+OBdXYLs
9SdSRBK9EKNrmf/uaTe/BuVzOCYNT3tDPchaUdNCbKojsTVs56fdrIRNI6lAJfge
HM2MddPlBAyMPkR4+Wydw0tG04+kP64lOAg0+VbqQ5DaeYZmgtGXekypDkCBLCzN
XRoJ5WqRu26ZQmO9wrLuWXge/BB2uJAqOlhnPiH54CFSDb+6dgdSENwZkkGlP/up
hCZeuaI4xCiI3u0t6TkmruVDKPnFWb3oAPswF5HA3boUqV2Ddp5WnfwRmMbW/vjl
nETfKv4rlRL0hitiutg7Yv7XufTu9A8EM6Udzg7kvX42tpp6+g8a9H/L1b8woeRD
J21LTj/1Jspm88BlrYJB67DLTxkSkG5dAOR1y+XB+L0r0ILArJsKz8vmZKVmlx8m
AGqFp5LDKunm1u4biA3DjnX8qGaDXK3QBxxDXqAeJv2/QvpBJPemb5k/ldCAImkF
XpGJ+P+b9cQi6b3U7ylxRxWUDD5QkyElmtSr9x2ota24nZklYdu05ghdJR1YG/pv
ReqBITY6WswkmzfpBEa7hqN4RdtT3v1Jgxl0DpgB3ii8AItM3avh77J88X2GI6Fs
A85CEUjevhk9+KHidFn/I6tb2HvD02uFa5Ej1+cXi6OWtoaNqGBf4zLjKzCCF9qk
zNOn0k/WgLlqNANhM/VglcYqyQHWGh56ixqF6VqSyl1xiVwiSliz8CFvBtoURnZc
jIaZ7DLByN69mdYLJmta0f5v2UmCVr7V+Z2pCRyuTW70vin28PyOpGBGC6rdo9iQ
BAcxz/gYLKn9KlGw6cctgC+J/HGUfojZpx0YiaHhbgAaGrzo7hYAUbPSh1/KWPEL
IyIHE0B+GKmhrsYj+9ADEdsgKQ+dK71TA7bWcsJKEAkk6VAe6SOp196tdfjB47li
PPmmzNPg4hGx7wFm6gNKyO+nhfk3Sw4onJgZV0DFbHOz9hd1AGYtCPGCnXNYX2ik
feQANwPVzrzlGWlSsSz2YAFi94IPg9D8ziqCg325E2XbbhXFVCU93Ld9sMu95hkc
CCGHB9s2ITI+s7XY57prLIpshRv6sgne9SkuMnauDl+xFz/+7RpQMnxDXjh0ECyn
Rx+cq7n4qfFQnAoK7t7Jcro0EWFeaTUrI0Bkun1WMtSX8YR5WH6dPnvFHsvfib63
PGTINnO//L5j5l5DIR8a2FEg2cJbCx635pbZM311YSYGUP9h3VKVu0GoYy+6MRAp
n+dLCJdiAljKeUIl9a2h1OlQtLVZc1FMSLUZU5HvwWXCBvy9SByyOnGP56qpaOBF
/6WyS2nHEvuYbi2SW8db2Md+24u4DTJKCGQWk5lMIZVBWZ13d/DMir+ntB9iQIVh
Y+dG24s4tSACJQp72JH4eLo5eQM8WR+8kdxobzXHRAf3TBZk0pDuQ2oBGooPRWYG
P/RSsdD+ALx2bvgvwkaJnXQ6Jtar26r9Vq43a3o4zkEQ5K8uSbAMMhNNREHa5QtL
9Tc1x6RRgW+XQSVJYzFLLXHMkJ4m/BnLx+2SS7amkuSHmdewrTbObG08qcMbNSoX
YYt9eqFkbfcvRvAZdMM/uTT9dt6jF1Q4OGZO0Op6FrHqfcA18bjakvpz9hSF5caK
97ntbEqjK7cuWGz1/Xv7UCKuVddKVw+i+4EsLR+qjv95WDagE4pdq8i7FrNCZvkp
nV3uLYsnia77aDSQgZaIsOQS7MyBwkNODC5SJxm01l2d4Cs+Hp5vuekGgYJ7hrkW
07lBnfr4gSKyP8/daCUyLbuCqt3H0g3fcwkgbXSJm1shIq94bBU0MmAlwZwzJK7O
qSCdRylLiKtTaRAk8hWstflTkqpVaC4T6umbw7mO5jsnpDkR6iXVSavmXyfxOKZB
l0zD0SU02in7tTmfOci0VA/QrCsb7J1WprtiJZ0sIrP0u7izOZzodTraASYFcEw4
9qJmEklRiyiHLlIJUX6H48uriJnaa0TdU9xDfTM6aVOkd45WXmbolKRUqkiZi+L4
hCq21T81xncwMQLeFcWATlMg23e1AzCetffVZjx+NU7Rr2cIUS0iNBIGJkAoLJ3N
XTIh36pTk4kMheMAQ7HxTc3KwKKVGsnyDY0S+BcVjP8r2CywnlIsTBCtvQ8yXWWP
EXpO5PVkj7HNRVomhOddUiHyW1RasOQwV0VEbP3nMJzlzRej11VBKKYNxy2maiZh
PDYjT7eunMi7vbejswl7dMAOkbZ40rFspiJ4h6VeTW2+HTm4PdioIjNz0FhYhKWC
uEOhXAWPo5F+F5Ak3RTwG1p6Uc/5oGNCvivdl3LOVdprPNs9QPNihfKihgvo+Q63
Fn/8LiWpqjo3gKfASr6cOqLsArfDMnmIp54+GO1O/6VuXbHkaRwv8/wUbPeoA3/b
tz4L35+pDgL3WlAZUF4QnyZpl/nGJHBN9Cddv5RZ9jyjK6+9Zj/HVWhDiVwo9+Tg
74qoAKcv7BKBRgrpY+eQYjjGRX+IS8boPWUnp59F4FxTrT7KB9LNmIesfCj0NMDt
ld0zR8XHsb3JIkIQjal0FelSsZY8Dmsh5FT05FjGkVUmsaVEgFwb115sxSsuvTsO
k1UCo/wngS4gEJkUjiq8Y4JPPN1obEQLThk7/Jxnkbycx/em6KmlldQm+Tfp/tSq
qb3Zzi4+Jy3PdFhyjmeTbDuOVDo3we3zKrAqsPq17h/sUBxnrBRxZhsnBzYMW0pk
0fJsfX+Ut81TLhKBcvwqNvedEPMTKva4Z1OHfceSNKJ5NpbnpeWN2WlsNgzttkKv
8Hm/sUJkKGbKa2a+vUO4deP6lb8ovHGl0LDgtVHgjDUJ6eQxPCMliDlrcq997HTB
iWYOIeXhRUUaYzr5E5kgkLM/yuqOQ7QzJgCUc/APvGpQ1f7Dc2MTMxtR4z1JqseJ
b7Z5ajhfcLZn6h5SVC9VDd5pDppnJ6j1sMpZh3Pg/jHaMsilmQDgrl4x0p/XCcQP
2Ow0MVn//M14EHqM+LiqrHUP/Nmj9HIVWBeUAFiAJsVewmGUlEUUpR8AWMBlluOt
1mPMFVSD0wMBGxlXwT9lX1dep0V+O527KgBJblXJ7xWVsGI+b2LNlrmNzj90GaOX
KzKVBUvhKiDm1hmndcH4qej2dpaAAhAZcrHYEb1RnZoYX2E7bVqS4PeTH1PBwGcM
Ki9LHTDYprVoNOcqn62gvDy1YUVJOf+E0ljnZxQ7+K5LXD961RwZQ/DEteohH5R7
+bdIlCulfB/9GlALmcWs8dyKQWe/hY0gkp2Uuhl8/aq+HyiEWDtkU2ptEAHsTgbr
/AVKvlZiXlouEAZSFreAkCRxO/plHxu6GL+gFtBZqEq4/FNoJ7Zro9TOHmeQGYrI
1QU1lnR6abBrNtYQpMBl7Ezphxt1LqVDQIuxqKkH1EaYqoEd1ejJGnEvMJv+zeKM
HSoSu/iLY3nu7LfM+03ZHAAzTnPSN+TE12yFVCFVTd7wkgVOc2UQAgr5tdIgneFp
iyB3O6ch0A/jBmq8kcR/6RJgxzeu3QCtabbEcnRrDyIMW0AeVhkLML+Eh6PGEy2r
fPjW6IeiGnh3YFtpRakuncAm+IoJrWh4a3ML1xOrHNVmkuFH9n/g97PN+rhSGhP4
VJZyUWDURQPk/DSKms/o91hW/IrmT5So5oThq7/sgS/E0wIIUPEIRQTXu234JqjV
e96lFKAjor2i/apYp8DJ//7Hxbbac60NmWANHbKzHfvdnUW6rcbpLg/DzpoKpB8u
xNhZWmULgQRV52pqb8NX7PbH+rhCo/i/XjHPqW0DPq/Wf9BID+2m1cx4HY3ST0Ie
MJXPqpdzhPwFt5ilGlVNY1FetGkUFgS04g6xdyuwwQEX4aUM/XDd76d71SjLfMU0
SuWh0UPItGaim3nuU3m3cFCo4tY9SlPjHTdoZnj1k4uCca7f+ns2wQ9NEI71idjL
SotpXa31eoKF4dKIq5Y4imLzBXlhi+wFgZvi5Lb9KwoUrIGrRG7HovPQzNOFj8at
getQZl0PAzv74oC2RkhmD32kCMfTUw0olfAyKq2rHRbihoL693Oe6zV3iy546SqJ
lY2FUduAYhvN8qGQVUFyreIE7qTf6Ml6kSjhynwVsnm+FN2TeDmTC4t9lEmrI+cV
tAD91+MJgRaFLsACCnLrRl9zyNwX4QBwVBRk+pYyYZwLXKWvh4Gf+kugT1F3jsV9
VA7oGrJsE5gH0Sw5Nmd8Fo3rDzCD63Y/zw2kjOF2vxLc0Zcd3agJhFVUd3fBGtBU
jxAdHMTRrNKqDn49iRiZd7KEAj0A0wv2hijXW3I2BqMkaXXpdZdiBbv7h89bPuKd
6PqWyHKjvR5UTiTEOlpDHXU7fewSMlzJnnt9p0gS7jH1d3F5OvZbykF15a65CfH1
X2MQCa3iuxuFkF8db50fe+OBfR95z6rtMqF0Yi9gr1euSxSfBUF1Xf7Mn7QlYyp8
ej05tVsOur2z9isqYz7IqXtMxhKJMKgWM7tla58ncRZ/bE/EsjeezPZgrUJV51US
GX4VyACYcnJTAH7tSKz2hfJLNN9e2LDVIXLo8R/O7lrEjEyTvGj/fDNZ5ISnkrLA
ggZmDJaSqWtrg1MXe1dicp7oSubnNsYcAOfDu+pxGf2DI8thm9/rur8EcNE7QpIh
2F0AEFSexB3stpmc03S6xnGEQpHrqmCYZP22dahaO3vb5zqlmQzzQ32SS+S8ENdm
iVZsAkKzISajZVHQUHK1lmwwFeT2JMvJ4iXapHNcdTvDtNbtXeD5AFgqvql1/k4B
NS2hAOeQVuo0gPNfKErMp68ODzGEUQOOTLHQv9lZ66CVVMFILiJVxxuX6R/2nywB
5DhFEvtFaJEgvpH4OcsJ+E+2gjsH0lPcLpy+PXQ2ta54Fg5PYZWyouIGYpyJCtH5
LsQq9pkkmb0Wm4zV3/3D/gZhTViSJpTyi0/v2mUnI8iIPK/ev70KEemkJ3KisNE8
ympDRkrcmVe3rHnoQZ2K177p8r6+lr1HlR0I2pmLMpE7Wh81h9lGZ6YAlrKK7U6m
9LVUSXfrPdIN10Xqt1yhlGckDPM+XnpbaoX6+lvE7aH/HdZAMcFHbbEebq92ZMBD
tfMMNvq/VLkGoZ6eQquff27WL5GjEsUHyUqOPp18q/vcsEmowNRApgvaw2yev03+
yn/Gysh2dJd7gCE5lfQILhKVmeV9jMDypXfMlXDAe2PlJ7hIqm0yiyq3x9uOgNJG
gxq/Q6MEId5DfQq/cGTNxW6vQV6laS5Uqf4RtffeRz79gqomGbL4v1eJtrkKwWoq
BOq3vyfuNwjofm9G6UM1j5lnwo2ctFlcSAiN+1mAfZ8/jYkQn0KyAwushYipmGZ0
tUuFZpRXpUaZTOZSc1gWUj2x6GSxNVBKPtT8m6QKDmtgi27A4oQORAltMz+WQYK1
UN3WDc6LllHE884DWySYlsQTqoHanXUa4ttGRA7RLkgChMz3XpO67643fCSqEFCG
Ee+KCCb/zkR5RoMUzRxvYyqhyKbyKccPO7gm2PHhWvZ/ey1GI+BoiuQKcqvJSoc9
4TEw57isC8Ms7kmDpcNBK/tVuEmVEU4QEZB49wbL03kYJWEVmiMRtH7HO4VYVllB
632Vsrc932c/pZXvSuNm088T4Ulfrf5w78KhcZcKEFp1MgtAEoOPQTK4L5c7GKJY
pGe9uKnAN33NBBYoGYfpVxpay1ceGZRkc9yiqXU/YexoboW7DEG5DyqXOwvybZJT
5FCBLmLpOxR6a2d0+dP3BxCugij8Jq1b06zI+POZkV0wN1lvWeU7+ikSa3CMxM8t
VYoc+lyRjumQx1TAsUTmm680+VOq93UgbtpXlNshdb/KS8tQJvKZK2nNHDVhtwK+
9YUi+NsB/mehf4OPYfE+xyVMLBTem9MeVaCj7h06QGkU/WE3uNb+OVlI+qUhf8A7
UN/V5jIRrMjD0607IyNmjJEytmsMLnJuUmJcHXQCcTZHwAO37ZwfPThSiMJmROOp
AKA0s7sBOzbKVTqGvIHYflrOH5MBhipwK4x+tMlushzazRMC6rxVkQ/hvXcpOtBs
9TLrREwDx/t79gEZzDbYlBpAmLbwpjELgp8vKufCFR6J58mzsfz79liOhoTGs3hi
02q+7+pNiA/4EVkRNL4bxC8mhMiclQMD0paeEQlsPHCXo4wwhf2Uhw+irnxOM3l6
JgXgPNtPJk424R75mWVJwREWfGhve1RDXOc2q1U77LHAYfLCtsR5QalfbGPPT4Wn
xMQfAMMDDywBRzAAol9ubZrOXz5YK43516nx40ex+ogT17FZN9kkrm6gw9dNwFVj
SKoYXEWpNcj3Qy6b3m1bdq0k46j+4moWZnayYRZSa56eCzFKQTs489YQ8tgB+sa2
bkR7D7cja/r5do3QXk1Ubp5qQ103iH2NXKV7kyIlNTpcZQcRF+V0iqUIU8dABtuS
oVYFwyp57MA0+dUMb8T1SOOxm+7Na1sZjC114n3yhkdThrCM9zxIyjpwWqKxb6Nt
VXTVXYADdegLMJkrQ9py++h1ma3M6Qa4dBUDRFny9e/xE6TW31HceUsqMoG3S+dC
uEarwVirykiDWmxvHm/UGb93yTJoNQyKxcpJPXG7AQ6HzB6mDHI6c4ciIAefUe/r
x0ygNnzGnBMwQBaU51mbyZkl1HQPPN77dt0ATeGHXopXKrrKiuOdFTQ0Y+5n/RMo
5aHdANkSAiNrJfwvuFAQgaaWR5ypJSwZ48hIw3FdgY8hiZ0+99vteqfnfyXFUeiC
fG3Oe7mHe4Ckw/lzwqr0DPTnza68F3fOrKgcZKS4PtmeRLMmeqNydk2LoSuR6DNg
cDKcJGSghjzlC9oyUla1neMxlJMK87odKYpIvX3pXAf6aT0JmZmKHDrVbqk07Qre
NAp8ajsN1hLgrOuD7CJ50V7obVccyxP7pEk8W1Ld5zPrCrR9tlti6L8O1UJsy3gr
/vLCMr6sbQRoy3g4GJkPmP6ee122MaNh4glHcI6QsjlCqrVqYA/49L1jFkZ0uDx/
jsoehaacdvLmjRhVr2hlBwVMLBXMHJIiJrkiybNYI3RI9lDXMhK3mf9QxIUhUpmP
O6oFHDxeLUiWhg+S9oyQIJr0DOMsn3g2FPKa52CteuUhj+yLKZbWYYsKA48QXHzN
4DpuI9E4t7Sb8K2eu+JsajQ9GIXeFAkqrN0cJHMS6iHGEn4SiMIzQ4J52tAnK/P6
JO8zzOZ1ypnCZbMPH8/CBIshDG/HxNgUoXIaRcZAYhsWHIIu/uLta0xDjDC54CnK
fDpW7jD6L2NHNIBYCY+6Sm5tWINsgI5cEkH2Q0EYSSiB7pzMf2yFnJAjI25W1Y3t
O9a73d6KF5c2BtB42JSVy0hOWDsMYKVlHmhi/ZU4naPZca5J/G+i0WbhWBojkIht
qbZf53p681hpn77Luty+KYym01s+pVyw4jWandlMvGvkvSyhJPKVqnDIOWa+w6cG
DInStHRQueCIUDO/QgTvKuu2II9O8yiNJmo0wjqNYC1SNqCGKpKfYcGIQwZ4j4Dy
BWOBoK/04pkWCj0Ch8Pp2vVV/O3ewSHzQytCDTArYO9wz2og4FyWxHoJrPP1mlBs
6EQrPB+WALizccl5bRZS5gqQ51hqutTkmTKmndw/lAqOo52dPGwnTSslCm6Erw4X
hAhsS479KHEaURpInVvCdoofwdjQTV8Aac/2Sr+Iatdmbk5b2n4utuOuH6YEylhF
PR5pGm3NA+YjwJKIk7xLGbL9TsQtiXestmARJGxoLM+M6u83xiUPEH8CrYY8JHWN
hap4FhsRrdkQxP0MzAHjCaQRpD4bVYXyxKewiINw7qzCMGpbImZCpuaGggPMavhY
YLc0LwrtAY4TASN3kCo6Vm7q5myqHjoy+s7+Z5k7OnOggqhfY8rzbzNtYbhkF+/Y
VdccI9PRdERsQ0rFSRmtin2GMfoxg0khWknZW7ILP1J0dUkVmtXZNvLBiJEK76N6
2CAfSCtckq3JhnXAYcSJZrclQM6uxx7F8kbQZKVpRBNXIUsUSfrjlzg2W2fAuJV1
O7ZPZQ9myZ4EdFYab2L7ZsSpe7tVOhlZTWVY0hzK/fRx9qqmXmo02EsHtLY2Fn6Q
Bq34d/D6alWNBD43MH/EKu2FoM9QTmJMP+NMWR0SQKs1kOs1jEBWA+dy48O+9izl
EdwybrZx/QFicDJR4w1J1LCUHUadiGdrprDKQNAlbj1IKekTCHc8uXKhk3jLoArV
+jR6qlRjybKNLifI+n9TSZERyfONsL6JeGJjCAStQ36c3U9pKh92Mq9M76SgRtOF
HSe39k1mNO4J/XGPVmhdOF1+pVSBJTX3LoTkL2NS4DsEb4IHSperCXTS0n8gYesq
Xlq03lpCcxFnDeCShsZlCAtw7uQ4phL+9CJOWfQ9E4BVSSFesud8EphgP68nkQbj
SxAPYDL4+OW6tJ1iGM2XOxCajk/PG2TqJgIAcpQxh79wIciJn0eOUuK556m+onnk
151YiNV+0mRZ4TcoffYbr2FaUwVk9EVQIuYh0hPXU03Gom2VRk4+HxCV6Bw2O+lp
WYMIEHP2jylyWipyQ33iHn3p1/DzL6yt3CjyFAD/lf8li0KIFQknLywFk5Clsj7N
7yGsTBJ30eJxA3xbq0LD0BQ0P720StEZ7lHlSkjvniAFArHERptv6Zov2ir//rPh
mrE1DAnzxI8FsHJPgN9kQ2cFh7P50wg0kmWceOyNszmDdpisJXGPq4Y2UIu8GHp+
sPn0v3RueLRGV2w6mJhIMxMcZDYSb8fxdMK4DM25I7kEYAEMkoaxVTLTanl7jrNr
xshJSRB6q9MHxwPoSQPr3tmww8atFXh41I9WHdwobxCCkstfXaLzFnwaeg2ZbkWO
1/+hlp4Ev8HpF1tAKx8Yt3ghnd+gF42t/ATLj0FXCynkxiqVvJNBC/1BwL66y1V3
tImtETM8ZNVpv7+hA/bcBuEgqKIstavGcjGnYTdD0gDORBJB1zk7nLglB6bShq6V
JxjLVebQuIgPw/HUg5S0EXZ18pHSYT2fTV0WyfEIOqkM2roe0BQRZ+Evh+FNRDcN
HuN+3pYCV1MwVfbAAw+nqEHmvsHXv8J6JO+IZEHrBUmpSeWRc471wZlA+mlIkijl
CMPw3npFtSbTawatk81ycYjLD/OjDbKaVf5ttZc+W6gjk5Bmpx2iPsHSYgPHxzwC
X9nw+F4/g12ZPvlpZKaN8SRb76SGfmhSNhSWUDpQpQ4Dz9hKSTNi1KvqqoGMAP38
yLDkrk4azQ6lQbMsHxzQp/W+uymvMwQgO94oArgnhoNaOpk85KGpqAssJ3eNnAat
LMdICGLVsP+8p++X4uffYacUCaTUvRjyIozVQkswUiDp49XdbYvHG/iEHrpbgo8t
4xNh5O+Wnt1lDF7Cfm++CmtU6XWICzkOvtwxShcYCBz+5+ESSrf0pMBcjVtbrYOR
IHtG5m3Y8QTNCB8YjC07QzdxiEYU14DjVX/Cx6q7YU7kYIhbNvh5eUYJDk/Aqy6F
ITMClKhf2sliEDy4bA9nA85GmoiFzwWuH5ekGLnwGgGxBGok30xj/unjtz2J80bz
ZsYUFCYrHcOppCxRO9kU8pljRJCHNOwDw1l6HyUAuHv+EdhY4duWM36Q6fS4KLyj
0KGjQqAHdLFcdHV7ePjTmSLQTtMlDLxAbJWJrftVIC0cjKE4Oe0V2S9v3ZtIx8YM
rZ0juU1D1LrBTAzOVv28tyXdF9Dz9fCzpIR5BSd1YI5yJvK3Yvxpa/NsaHWqMKT0
2F4RVPokXXShr8Mtr0VNOW60R4sxTZUBWT98VSpYtXoGPK11wI8cep+o0i7x92I3
WScV1Qq64zmBvUe0U94f+91hwLFajBM8e+2gPptiweLPJVPTNQeAMWOnRNNnKKjS
D7m+xZaMkhuzR6tRsaqloyqvZfxuydLcM8oMN2VktMq9dKI1c20ClFhgRti/lQKw
D/xXabBcRa4uCE0WYlW5zc+6stCblOQLwcNWEV5oAoReFE0g0hdLiLOwkwW4YAMN
t0EYeUn4pvK6K3jZv9gDsy9yti07/6xRsc5oMmpGzg1zHgmUUmiPjtaKmIyXl+ee
QIjMXkua0viYFyyaCeMXwIRh9+OjEecX45riH5MPkCpRm8KHyHzvcpnu+pAeir7v
K+maGT84YLOZYFdTWWjb5ADeXw8QhAK8JyikDytYjsD8f8rbSPGiL/hAHLQdJJ9u
MpypVvFz1P4+o4f47SRK0qwOId6XdK77aFNM9eWw/hmEsCvfW8lA4M5nYSETEOjR
bgUVEr951gMXhx3cELFFDJCYO5P22WQ2L7IwRVBgEW8Bb7OaSnx4lllSenE7HdQJ
oO35m5O29hHXh3XWm5pt0BYbOtNuvF+C/7rWhTn/t12zh3+C/ELlOwu14wFqVgWe
Ovah+x3a14ISsVVozGJa6569GWC9OpgZWnZh6+tVBWIKY2OPiRbOlLrqMAS1E3PQ
x5p7dKSVxy+K6+vs3E4mrYLxZmPljDfDl64FWXQbr7141eX9y6mKwolkItgQEuw/
QPtjyNeNB3z+GLtMFOe/J54Iu91DLn0vahKdMGjP5XZIjxOxfJe2Llvo3OTcN85w
Xy0IY4ZWXmyticWcIUPeboFyU4Ke9GuDU8rXrGUPY1SQAjaay53bLcW8k+teppjL
iHO6m9NxBd0uHiXv5Z9QPe7IxzN5PQP+qqufxBVUyd8gTwhkt/JbKc5SerLU+QTW
x2LsIeftsPmECX5nq6vVkr2SdTEmwHb9x6yd5OimQnKFAoJgo+/TwV7ux9y7y9sX
oXhEKS8jzPrzJdx6qVB3N0vN5o2pH5mzHBOIzDQpxB0/Fh0tZuJKQ0ngQIGOzLCr
bYG6oKVKMnKEHycHWd7TR1EcjTZS8PLFmasK/Qu/s8M3IHpWTNWdAOknLs2oI+Jh
lfLypGtbzgAFDoclCMtiZznb9usxQX08EESTRf+/Zijov+v+r5LpNYfbBLGyZdpt
FHGKJSIPeKVfgF8HnEmWC+QeuPFEU5HcvLIWCV8Bsmf09ZJI3Gd8lhDG6Wh0wAAY
XQFOeGa7lrKx/Rtm5lUPTwNexZUWq+CsrHSqSZHFmNjrDwBK44R4hOGzi9Hv7bly
i3ge4U8grK7rFSXnDxmgd+OhAT1cYHKBJ1qCWgXiGrXurNug3YUEjh//RvPbKZnx
PZI0ulHu4vkgB5aOZ7lhr57LIltRBtlAb1xH/fBNZ+NNj614yjDRTLRUpavrysLC
Flobrafzj/mKN+9Oxp4JmOGvRYkKyGmcJp+ZJ81kisPA3Lxm1u8dIPxGMt/XAfuv
WSmo/rrlssFkZh4oECzxv+TkWWeUVxYOUBiCS0c1EEy3h6uB6yMTJMFDzLeumdCF
EEfp29Nk35rF7w5AcgAW3dwDejOPOE5gYWHjNCTuFa1qRR33US82QTCxeRh5SqIk
7skzTdJBgmirnPJ4pbJab3zitW80SDmAzwYxQVejQoeI7duwtDUuqueZ8bhzHZdK
GOCjvSRqZKRRKwBZBt4jYddHJOHyFaFTV4QwW7RbrLIqIxvXhD31l75ipBsmPCT3
lrqQ4wXE80j53ZutFfsDISMyTiTLLBBwSySRR2kloBzXNcr9UfQCiNpCP5JXHPJT
kPcmBEcVS1GkZRnrdLAo4BKX+Jtzh7QeYgPxQK9aL/bURuyF1+aUCz26nshcgjxs
F2vaCGrBg61p5F879+Xi9OMt/YoOi7pizoahSCZlyr8ZMszxO7B2gSFidbqhwzQ1
pBWyj/L6dpQeZ4uwBq7uL3QYbHB/SaQr1ve1ea6jroNBD44XNQ9AqDrY9siqTvJo
o9QZNEt76inNCtn4JCtSNQO4Wx10f4wxPzxz+4Biy93zNfx4sGOJusfYz0H/F5vR
7WfonzwieNjitlErB9P3FW+MG2FVCtCe41M39qOLsimgt8t6oaFv6KqXhh49Blpa
9cINOe7WFxnt7p1GrEcEDqB0ZpKfTHYeOa8fBFSlv9DI6dzm3NyYebEYHC1kLzIh
adHN0xnzPOLfJONHsLJ6RaeJGdwKuRYdY7wyj3Vi7b8w4tYtQfRERkDw5vK5KUka
wMuoNYPELOpzbVb3qkiFp3RoTgCHehxep4Umph0Ba67yW41UaSLZepjm72l/CVt7
acyd5wYIwxOlHQRx2UtrtnC3fY3M+FFjyPpgp1T0Xi87UO93AGwDAGZvFcfnxDQQ
Yut1AlOI84ptEvQR7DfPpPM66A4lan6HKfk8ZXqAZf1vuz3osPixtccb/Oglkxvh
AeDRUoW/mYGU/jRZNem7dRxQ8ZZ/O4ai2nXwYNSc8yxuWkCMV2gaZPl5fmaZrDq6
yGsP1jJLlYv/sRIiciIkN4qL61ftYSDsaeq7g2i5YgaolMGvIGGRyHSux9/QLWEC
IvK5KYuhXZPsrTrwew5IM+JtvyZRgrDAzMKfOSbHso9vLOCTdylv6nNHzoYnDTM7
iKzL+1/lzpOTTgfGyCkclX54F7fzQwPw1ffUsN20GzlgHPZHASazA26LrHlvOL4f
MpvLJ3HP45t9bLzxrbZNGoE1mS64cfjOjnbxov5kNOsPgB1w5FMKkyxkTSmVJ68Y
IunqavQDzMPheyRpHbo7Wt2vL8aJ1qJiTKvwUzFc5T8M6cBVawbnVqVsiYFPTU6W
vRhSLXFPuD/DdZb9MwB08CYcHvpaqKblHOnuv9DCnYCbrjVA7scQNjRFJjRL0WtM
7oRQ9hktPWHSxwZJ9vUobzK7dcEf7hpg2HlhBU2mX9dHBCG8M0KUsxKHine8lWGW
lCg+fc61XLcrDs7Hd0mXTa2ibz3VT+/GwgLHrWEbf7H1wUrnGGn94U5q1+bsh+eE
rrhKKKVkFuCipDrFgJgsjc4VnaG7gEnCoFoTn5YfokOpXqrvG906Y4JPQYv3Wf3z
mvH43nqKzu8e5AlA9db1NJ4Fi/k/zh/MPsx5o2Dy4e/4VdjksLpPgx0kGOah0PMC
cv3WtnZQapelVplgdbp/7wTd5XBSmfBCXrkkEr67THJj46OOsp6vS7AT47hDrrra
jg74wl0ANdHCi7xLJCzVR/vKqnxiH+u5e0eVkv58+/Er+g1Priqp1WJG/5L4+nO2
LIuuerQOqgC6H3KAR/Mday5IoZ5liUDEFEncpwUM2Lq0oPlMoCkSxUAgK2SF01J0
Rk1y8pA5aPuJXgGjbdbGpnNGXQvGxsNLpU6iaZ62gVsU8RHLKiLyFpr2JWsi7GJO
cFSk5mD6xHcZgKKUISRXZlyfGig5rq57eSkN+Wv3b/lJlr7i59VW51NVid3Bm8Yh
iRYk6ja/UMW9J08ifyzpGb2bbobvghVu4wV3Id+Y5Ktm8Hg9H8lmRGxT3xQ1ljLb
9LWYXTwMmu3g5CNFrrOE0G11c79WxL8sufGPt6wGg8hUSFpCvYF9C8Vi4nqiE45E
HgJCSynPBZPe4v1pR8ar05M+GFTdSZg1MtVSD4LdSxGiKnNSYRqLAyvcpolvz2iv
7MmsJVjZhdGfeJK4yJ3R2lhAn0sAXIFwF6i2ktOGf5K3roKu4oTIafmODx3YTtuB
HmjELa5S1JlUPtQeEMtgwVFfiiZjziszeS0sdnY/c1P+bUrJ0NAPnaDnrt6sYbli
wmnq9bwWUy1mstfhA18J1ezk7ipSZupvlL8HlsT7X6liWQhk3rxMEHzKuEV8yfB4
Fp9vT0XTXxPUxt7hcDIhaiwBjtg/Hhu3EaanrTUJMQYp7DQl32JjSJGUws7k7tR4
+etat1Cz5bh8dAYHnk5jP5zHElKdC0dc2Yj30ndiHUmi5gQ8CQOC9+XNYkOU/u3Q
L30B9CdjEBC3347y/6djCTKEK/RCHEzoOTaHbSCIR6tYqJ+wviK5N7loIULJ3vS+
fwGm+OKz0q/w4P4UgwU4d2ij+OfSJFQhtXjvYI6YOSe/8ZiSrpXU1cvGALbhnWtQ
dkK4GLVFNk+iyjlGezfJN3ceMt+xxIfUdkWxyQmPw+P8v+HfLUkdPgL7uQqhJ1f1
WwYKOtbvyZU6Um6I0I3F74KWRa93W7yMC1h+gS+MctyZ6HkLCOUKWi5ZzQQrQVXr
yg+oubKChxqBNH9VvKLID84gpoFKrvfizTlvHd9MAcBnDZoCCnn3Rzf4bV08lZnw
lV5f0sM76sDtuje5dwTYMX/tpuyhPjSVDUZ715Lfh6JWcwaRDe7i2vxtLY5njlsD
fJU9HMUKG+pNOiaoNgcUdKqVLZdHOC9J1hhFxhBIT6odzNN9J90+cAL2SSTYmrqk
GH9B6VqFw8q5Yt5NbIhCJ9NU251I5HJCPyvrK3pULWh/ko8UJMeYX/gZnwyLiDZg
yFxpSUlXUbaMhFtXpWBzcVWVEvr/nFVFZNPrCSZ3agxJh/n7UV19jDSPsoc4O5Ln
/ED8OPzJ//nwpY2EqlIOVeGGRbwAASTB1mTEqAfZpywT+KOKD9NrLQTR9yxvE7HC
CCHQ1Leky7kXFpolXOwcCdkjGkTFLKCxb88VaLJlq1YCb2UiuX05Qhw2hp+6g3Yx
W0YU34DbqdVl0YtA2yJmNcCBumFCexDpkEl5Z/zBxybTelcCKB2ZS5Uzp33Zr6AT
UdkCWZ8n2OBYEFLuhPKHF19y0hltCT60gbSTevo77QlvoMRgakFRBJ1bsKcdbWRo
WwVr3M0QfoZnb/ZKclOpUh3VSmH6BaYARTJ2DmczxHd2b5HJiE8WitJjXdbN+QnJ
q87kR6rJJKNrDiMT93YIfUH5PHFPyoc4OOx2ouuHSZubzH1/e5XiqGXZQcz9RVI6
5QWgo8O0TDWjSzf8cuUpTkwW4ieEpE3u2n/Yf2NOR5HSPvQaneCTMIq8SGhOFHz0
v0CVRroSl8uty82HsRWrdj9IZX+3Y5XnV+m/VJAKSUrnwj5sQWicXb7x84C0QQvd
84RmNKg8lZoSZ98jh3jd0RwmZ7jzEI1xhH9TubWGOkpyoUMjd3Qo7lnTf4TBT36C
BZapYoVvq9Q17zdYbPdpAk+XMg/oTJwoBQ4JCAGXtunBdqFyoF6BjVhLE/wJKUcB
3BOpV99yHqaqRmJKMcGVYSndERjiU0nRFEN9fCqTxQUk1E1MFCEtLGMROuQJ+d9D
an66uQxMOU6YPXtijhyjodSL/gSo1HqtxwGJrWdYA7Ws9tZGAx0Ae4shbsflEaBD
HI3OhMS7W5Ehw07e8ZH5heTsNURfpXtDFgKr1z+96jWMTLrilUJmnhs1qqQTIERg
FxSuLaS5S8kveATjOY/TwCxaz1rCpeYg9CDOvtmFUcecIgoSGFnVnVfIUWTmPC5P
BmGnbf10dgPDraWRXhep2mF5LnObVlTt4zXJa/J8Nor9gzacgLN1e9uk2KEX/TmA
gQT7GpK9wsFKvCJ9R76hNTzlw2a5qf0z+hfD6VXi9HLLdk1sGyG7vpbwksmqB4tW
J2quCkJWEY4G76XEHscnPw4bjdW50r4+g8Z3cQWtDi25V0s8DFUm+cad/uUTUBhw
5uSTwARoEOvY/yA/Zp8ZEUAqUq9OsH/G6Pho/GIPIOhbIQ2UEhdmkj2eyERVfxtw
N65Yd0jlgiBx+rC843NTDcNASqBLzB4ppJK1WHoauoYnp9HbadV5cA+hID20d5YF
0cFTCHTbTL8XC5BSuA2DwPyXIvURUArcjPc5npbBFTY848LMMg8FlE43gVeq6DsF
ZWsA6IMcnwSi9nv3EEhwxK8Ook+jDhYpeLZq2UzgtUBJV7kwfQNy0Oc4MIJ1ktq/
fnZXT2AwZfUuI2EhnnwP2Lh0swnjvZq2a1d0zlUvmtYWD5awcRVZGJ6MYdoKxOCt
f+ZCbR7eDJe3IATD7vNPJEhJTXbkkjw8E6qzNbS7giMa/BCzl2ElNZK0QqdO8irD
snNZpfVhkkcXzxagm5FAryUro598E888qCWTyg8Ei6EvaeiBIPnbocD7IViZPgxs
uSW8WnvALsPXHLVdMkJcUlGkid+JNSj3LPOYLIZdc5nb5pPW+VOQYR5nDz+t0fG7
OzbP3M+q+9/6MbkAXnQurdI5wOiwGfYEYCBg/NHcQWd5YNDzOrMfkz0oHdXI+r32
Y2czubIREaYTbA4+Kr9y+50rUBEB7r+k2B18kaDtHG1p1GF5O2OzGJ9XEGrC//FJ
BOCUqDTbo/3labni5SWaULoeIF6kynOAMHPUk2120HBBRpqLGX9XfZ6y4kkx+BsS
pOngyyGJEJT+n8Ajbk+lfNACkV/nnREQA8H7S4+BBoAM/v6wplzxoqoVq361tmnC
AHwtXVC+PqWfUbN4AO0xrxg+ib85fZ0cKUdmgB2NpxUeQeAXoohxqFgjaCE7D/L/
F66C5w0auc0PifLRe44WL1CwOPOntddOO5NM7fHXX3NfXVnWMTzqR3rlic5BY12H
j2I4G4VN1gx2gDOLINBxja7IWo7t9s18kwPYj20XjSP6s/QY3+XbyHK0vbSDE/Ki
qJd1Wonyieg11mGNUozuDFpYmpaZuVXZSRVGOy5nD179upnrydwRlHl0RRBVhI53
cV7ofFyk2CymoebENFp0wEN8vZnndZvB+tBNdMRK3H4KoSvWHLXJAT9+gvJTFIH6
IYe0gmyr4Z+2mhmkWGS30vdLm41g+GlGCpFl4nN4C7x31JY8X7wCFRz8Hvt6y3iR
va3cgudI6/yZv+4JNLVlIQNAUii6XvBG4cxfBU+zwNafO9QIDq2wHhXhMhj5UCif
Sp+xswuSi5JqFPsf2Rs6eOSbDSS2JgLXvy0C9JVOLIdAEGJ9ihLiKUUOyR4on7WV
7RopvpQjVxLBS6u4qKlGnwR/h8/Z2+nuwyYfhvzQzptqAiBtex83xdV0BYnQRmD0
WOfnxg5HOZcJXeahRdAmyW5WHt8n0Q0v/OQCupr2rwhQNRHMItGRjQX+99XrAnFJ
70pmqJzthGxtl7jN8GkEGeUBJX6qIpeBUaltlL7I6L8baB9u6iKRKP372fNePxwU
27vZ59V98FzaM4cFqA3z7opebJxyHYYxfjLXxXGwxgUGC4nL1p3W3zgYfPrAETKd
VUUnxoRj2pngT+oup8s/DW8jmISklFBGd9FYQYe9FrhBQkXzV95VS12/Y6t/YRcS
E1i8oZfqS210/y2Y8Sot1nNZRuWqON/5Xfr+odMTyziBEE+oMz6COsuQTkTEflqO
j/mOM4/6ASbwsTa5el5W9d34T2pZ5kf4Q6DdogqjsSAtU8CPd5LCwbbwpdhDcFbE
f3o58Cl0W8sXJeqWTWEDSSdKi77kyHt3PZY+ix5whqT0cnrVun5By/lYoO/3RwFN
F0FEjVMvWrSmlul8d9/GyOE71ET0p9LwyaHNbsMj7oUaAWJslUwv2itfRaKN3Uzs
BneCW0t32s9DOXkKkQVHn5mAHi0UUA2qaDUGMrIqwDtjWWVjNxFMJYhdWrodT1Mv
TTp789WDtwxw9MGbHa0vIrvhcLYKUHUkFbifSPnBXDatgCvXuTWqB91DXbNN7jqR
+egNzFODv9DFlgRq9h3Hd5ig1BvOTHWzuo59RQawHmX4L1kRIRAh26D1jS5s6eG2
gbYbIM8mp/6n+E5VaFPs1bbxKfSSBTucwIwrbYlktoyja1Q01iHXijYYjg6rm7uw
5sKq//psmarUQsz0PRYl43uCt45WYnpCySYYg+cU/CkY53Il9GnrtdWOjsen8RcI
Gg3NbCJiDqYAFnnfM0AkO7nO7I7bawtgwAe4zhX8gtaQIyz23MvL52LYZX7rQ17o
amYSdeAgTqrl6g6+6ua34ApoovyYNLjvT5SQgwUEKWoqiwWj/Xn2T6TxOh7clIt/
6aUXsEefFj8rZoyYoL0ogJCRUTrrssDBJ7OuICj0dyYMv02guzciNrEYmmOvnf5E
dds0Iamb8uy8BBhfp9WJwRWRSGsJNyNOyriVWQLiTzW4O1PiZ48GRCujsMQnHEB3
1b/1O7LTcUHOyZk3TRbNYqWg+6iZTFlVMO3pVa1F7b10e9wZMd+F/2mQ1zwvPPMu
253uQMPxk+gy3GIsUfOGnhOdPf1VuZqNEQeDtHLnhOY+bHn4fayD47wEDyfc3igS
Xb0VxVUh7m2UkrlNXCQQbl5FJA4At36wUWcLmx/nwrh02gM3JhALHeWzzbvi8oyI
3Z24h+pFSdHMtg4PEnBMtkvar4/yWh/9IPiQga4Bl5rWE1hgsoMOFPVBKBzM06Kt
r2nRe06xJ8XYRYSv+3Kpw9J3TE05gC7oDyZQFjKbKhopOzQvB3MtUou44X4L5bkA
E+Vdv41CuaPjNniyRdqfPwNsRKxBI5Yxngh9zcIZufpnBSP4L4ngMs6zwtxjXgbE
EFgQIQo00X/c7rORpdKZY6/JXrFIhdWl0uPF8ze1XHAZT9hC41NWwe+t3rz3l7HD
t4PaAHPMawHQOPzCCGz7L1N2S9UEhBEonaZD4epjGdXZMSbym523r0gWHht/4ptS
IA3jjSdULSIUF/gcPZV8sAoaMgeOtIl7gzvOw0q1f0FGPVkrEFejqTP5fkrxFoE1
I1dkeqJDafYsXXVyBPos4urFsIlqtyRTaFl3SX1OD1Jv0c/cCTREWek8n1Jxr5hV
kxGxSbEbAbkuLw+GJXbiQ851el/hehndcSJ+Z534DJMUe3sL/AEusnAzEkx1Ojag
g80M9UDfaumZFl4hy0oYytzeFbtyM26hE9LAyNfy6+NfoWdqsar7VIdJEEN52LyZ
9PwBennRd0Tk8sMj1ZmKfomHDwwUfEk2NoEq91vP1Ow14cMW1Zgy0oOTqr3ANaqo
GeyrC/ZrTQcA8cYllgnXB6IntXWcZrWs3IMMMKoLK0YdHLBV2XeW+7gWXGTFpyci
AIZF/hKKgTdr7T8gws8nlm/xtWNaXb2+dJoaP9o5jPSkwJ55Yf58rSv9rpD6AfR+
rEDXKPvaDXKfLvamz20zMjx0s2Xq0sNx99nY5SCNtcjaZb9qZCkeaFloJsW2g8Dr
onDt/NYfELFzh5N5ZYbGA8MGhMWg4S6qgHNoLP11pukgKRo/0fUMpV0d/MHI0tu6
3OSQyiTJ8NjC2afNrM/XDuA5P2d6cWDC6+H02SxN+QjaPpk1mLnB9Oie4c4A2UrE
EofQS+fhwOGqiOJ+TqxMq7gNhyaMcWkLm8C/1f3uTWW/ZswOnzrMfH7frpLZBPSf
euC2nnH3x8XlyU4/zxLgkHJ/QnjGQ6KYyf+7/+5HvAJ7J75TP8/OhUxkJSLgf1s6
LB3VE/nEyogva7AiiNa66QJOrhZIfSA4NT3Ar58+SSyaqP5/35aSftPNAHgR+dww
GUCG3F1XfjsYOJU7Jnsp8ErtW2Eds+1gv3pSDkE30pDZFt1uql3XT69zYD5SkEad
4MwRJB9mlV2OgZv9RoOtYZPU+4maMBe6tA+VM41+Cemj3TxOxwdf39M4pC1wjZVd
CKMNkntseOD1FxBC/V5dnSSmBXPhmZdU/olnaTiK0nuDzTP3QobpbLssCGHXGl8q
FPbk3CGsQ5VkhNoBXFQJ8aB8NZDw4mB74WA8hUT1z0tY2y2c7vdVh7IttskiXd3S
4JCu7JfywfQPldoeRqGGNzv/jGuGj7OtfHmWvOtYYPM64jRkHZXZirZOLfp+KdIL
o4O5VW7PMoFxq593yqT60g0IQpN3cqap90SCJC8gAExiK9q7F3vLIRC5L/dEAXYs
2iW/EjZVjYdYP9U5lWSkNyOqccyyRqs0OgQV0jL3qtT0EWNiUJoE6FXYb0sWCuNq
WQcrDBlECcTU7mi2DwkhRsjmzs8II5vs2jAWrHEHv2+UjtCGaH4uD4kQ1hrckFsg
wXdjdXubCn1fucVudc/dtkGfjGkMbdRxhelQa4zoUs3SM/vnGfaHVZsXh+68PKl9
MnNtq5BsD4NWnY4mhsPFD3iV2g7F2zuhOayuM+G/Cz+w8OETHn2+bDjfizkXGbBY
t+zAgvSpmYfMbtP9jxnt/Dgya0ZdVpRYa2MhHGKdPn/mnA0P4UYfEHxGSfOboHC9
Bs2Pt9WKHltHprZWORfw4rllc/xDVw/WSaGle0055yHKc6A9S7cVsytBI8Dybfzt
Bw7rqJyf49sMh+yNiv0NapqBJ79x2QecO+5tUHhKtmMA8fPZTE0pPCYIaAVoWR7t
0nHpnYujHuZ5njy5Qkq1/tRq9yoceNtbpdsZYIofqKRGhMJcrBMQKLc5Myb+y2Wk
PHIfmNWhp0iJ/ORfgVspRldUeo8XNtuIUFZttvT7OG11vS/+k4MCUYtP875MbX2/
3kQyx4YhD1Vh6mTO86wIrtQh6QkqLEB+p3/t1W5QDK1GHraPPrhBgmRAmOQgROxm
GOUTyovAs/qHGtzpBVToiCRegDbAUaTXi7U4pIVy900BZkOdzAXRC4FkQjXypEXr
VK7cwQwjqfltqUrUresCr0tKXppRMFR39e6QvlzzjnMR564PsX4Ee0j/Da1xB7zs
3xxns1UTLLHw55HNmoAAlauNz7Ao2WHjdGZ2fQBjFTMWHJ35dm1SJriUdPRXzwHT
2xrTPJLxcLsEi84J+wZBHa4dOArW3nlW5OwSWIjD1Ia2X4oH+PWv8625+MXAqCzm
xcRFwQPhWavX/Le3MxMFjSIe1jX8rnpkEoIYyHJXgt1ddiUHykIFTe3ZgW8MQBSL
PZGJG07gWr2U+BCV/VIsfOBWhhIFPfC7s7AUHbdHYquID4qkJr16TZx/n70j9hPD
pJ6BVwlXqkQahOYMDYZ8I7Q0J+oB/ViMTA4PuXIRY8dnaWu6Q/tYLnpLsFmf6860
WxdhN3+OaPu8/d6RwxIiyb8eqBzKbHY1papw6NEw6xoDGLlkQ9SYQEEj1VRaZNoc
oo0ukdS/P5uFoCH3vLbn54X+g/ae/UEq2cgZrz6Oc63BE27oZHoZ3SnFed2HlUXV
QYmj6Gg1ReUqDWlvjSgKhPEh+rjlCJPlvkBHiK4wDg6wNTY4CFygzjRoOrvzGDR/
72k/e/u6QasU4OICX26NMMQuX6ustRYUzgRwZiQC3gmAVuz7UZD9FjiRvSKJNgpk
aR4F2DEnD0G6rLl67kQARW2B4iHyDLnod5G7QeoDr3UbakiEJTuVH7JOK7W5y/VQ
C0SIej9PKjMmoQWtpy2PjGeWO+bZtQfhWLPjXqaUS4qcSYii1P1P0geB+CQg/DUq
ee1af0mnqb0UyKWO6j4qqw6EdO9Ex1mrrFvR/2ZgWIFHAwDm/trjQs+uMdvQpnYM
ZXR1LhnomyKNSdIrrlyzrFAbWqi3MCIgI2gtPq0pqnTqlwrmJ67KKP6pbwbb3Tpo
eJN1cOg4NTHrPkStmYn8ZgfOyCnD4O0DOciyXiQ9HJGrzzG1CdcrpYuqP7v73zxs
q5YCNH2sEfemLb1cxdvIjxPqqszHYAVdBQYY8sX+CFt/y9V0J/VLDRsvSqD1Jval
vUUsNWmlOdJpJM39Y7Dh2IO/ujqXAh5UAC6RUhhvcCmBY6FfXlk8R6A1vIav/Q7/
vxK1HaRzL5tta4w0XlurWnLXa/x85GiQ7C3t/hkgqdH/PL2gSL3zCSvKZ7L2iqeB
+iVUk1egO4XqRY/bfvvBRx0hYGkxN3Pis4igE16HmJR7WI+5HvWe2lM4N921dGSY
XA0VRiSS1M4uv4LaBHAIZ+hj2FDcxKmHWhdJFVznjJIVRRROdI0sH04AOztffUez
KO5xkJ3hRh9vl15o8Y28wvor3XQ4NENUe9ezsFmeC6k5MEhe+QvJqRpxoPF2fEr/
ZmLo4xoNfwhJ+XegEm7spkc0gTJ2QpDEkYPaXVLLTGREJsCtLKQdonGIY5qinIrk
EQEKY+peb2Hwj//SzDO6mIz7ZsqO3EpEK3o69hkAycEULepntcJPKZU0vdevjVFI
+1ab4+IZQpFM8rR2ld2XGTUZNu3rme87kF3U8QAO4MOLAP1mvhG07m2P/nV69+sY
57WNPiPZVVcPq2m6nSUiW2Y52EEj6N9mPbtUsDHIib/xpdGVRM67QOHCrpgv5jYw
zsxnY1DACFTiDvPgg0+C4nP53j2njfNlW7FU7D19NYZoPAM8wkOh+BwOVFbhqy5d
emdxtR2ZPVORQIK0t8Np1RsnB7k9102gB0LXrtNTBEoHYMFSNDLQkLUHchs1EZhs
ZqFDPY65f/D1TC8AUBN8LDzdoKBILBydDRfMwZ05uc35KL34aD3Oad5bm25x//4W
6RsQo9X4pLL1s/EicDuolmkT5bhOvPS7WbwCcAKW3FUfyV+N9F3WT7woEM0n9DWv
gzgU1Rj2d3tDxSSydIRYjoZBsHMfUND+3nXRld0/0oJx+a6EiAchEp1D9mdgbVWm
A8JndhIy/urqmfRCj1gptJxOhN0QAMEe0BLfGtIrSGmDxz79zUHMUhTV/jEAzed9
qw02QSTbKHAcCbRg7FWeqX/pcGRQrAi8/0ocRVQNHU/gtHwlALvu62vGXf0LKEmE
8+lfKw7dbVM+7/mygamph3hxcTR3MjxgOH+y7pzRsQ5RxpBkZ2oxKZDwuf2KrxpD
Pq/LCkQX1O83NF7RBMZ0WMz1E+qhA+1fbnVHakVGxN8m+KOLvStewF0+uFqItaWk
SYu6H2B+69TEEOaofAQhB4pBwOqJHSNzUDadfNuZ19PALb7bHkCozvmkE27XRvYk
6HD8K/x9IKj+fC5gAyHtD6GrC9Bxvymk51ZOkc2d4cpvrws6DiUMH/UA0voE7UMn
6yDpqa9oSp7Egv8c501sXmNDokXweyUzoIe6LIkmaVkbVxLKNArYiTZ4NNxF0W0h
ZdnKjwFvHkob35g4uH7hK8DYQD9i+XpLDIzMy5OwOBPL3/2je5RgiXWdgvocUfSG
BR7OVt1xLx2v0cX/lJA0kuK+oI8XZrATNWOTjySUT5x+/BDjkNxw4JVxD+cYBPY6
BgNzTWyi0QTuayGTuR8XrePefxV56tbM9rycUxAZ/NcCJNjj5Kf3HhdN8wiXHF3e
l2O6TnFegn3OIfGkY0mIB3XK0yDlQCfCRHq4qP9/lP4vY6vV4lD9KIywYNIKy3YP
howyVu4kxQjVtnz8/An0Zp48Nm4Oozi0AyPY/QwRMJ1Eci7RObu+mJIdKAbt/qgI
rhluNyo9jOMjFpsqzqF1pEUxc5IE53FOTPAUQYnspDhPG8nxQoPGKxzA5nmXFKMk
WKC0AO6/bfyEP6rZBHiw2NGtpcwrdXieLfRZKSlxPWbBL8g+ogYqLVGdBv2+CJcd
ckthchyN+zQFKOKFXHAw8CYOczY9eVo9EecQPYBdl0msAcJnCx3sY85tqGF+srg8
nIDH4prZG6gjzpud1Ohw4H9UfA2a2aLPgOBNCN8RIZGRN7aZo/yTYNnFX6XzvOOO
14FvMdynVbaOUfFFSObBreiTHg/jyniDEyWuYbGupJDchnRndHMkZSXBNN/NqhUL
kqtn8HouEIMd34XaDYEuPTec882IrIQIOjQlPkxhuU/PeRHVwctlzUaNkz/XrrQw
iSI6zSKDx3PzLxdWW4hRLaly8poc6ZwUnbxZp+ert/APOtPEYksmPNf/W/yfuTOI
4poZnt++pasldkoN2zhcHTPV+TS5pmaVj/LO2Fh8ohJG+RBGRX3n8p7y2HFmWRKI
TBVCzEim1cVHFmLWcBk0rIcv3jAXsB0uP9yqFED5QdN1Cn6XnskttGeWKsaEH+id
WDM/ah7PG1WFZYmeOwN2kmOkYICD8Qzq1Zvb7VlJYOL6WvrvhB0HWKyp1+EL76jR
LQK3Q5pOhXtRUjscEQpXwW9lBZiEmsSswh45BCAnZKQ9SBa43Nkv9W3gPJYQw0yI
WRW/9zg2ZI0pmHyvIpw4u3uLR59YJdieq+unkI4gp7vxD8y9Vjg8O+qT5wCkbcXX
qHf4AUoc0b6V4kCDBHRJCmhIqKV8BOEEcE8Y1QpV2sMPUF4cDUoI29aByokXOAcc
8VDzL8U3vhOKamyT27vu+McW9RIuk9iIhMWy2U/hkwCHrCgwpEG/SDt1LPbIABir
LKvQNdCCCXbsZcsYzp6JhDTiral3nlMZTIYia/W8jdoC0rFh8RBi46V0OcdmqfFH
NtzwYySQjv21EZP0Qc8z7oEh0tuOEohfu5R6NU+PoDAnMmq59Xs1O5vxZrAWTUGW
OlLMqgi1MAf1s1j3O02Jlo8IIJ0kNmwPomqhsqF8grmmZOzYprven7SlWD8hGFAB
vVyOAdTV8aTR2MWtkgwkGbqYyZpKQ+t0rYFdlFHcltZafKha6bAVCi7GIWPslJo5
6S/+X+P02O/GzehCJM9wxPwHAds/89PtrFT4aeTa/OqS4zWp0D1VAkS4G9BlPINl
q9fgRM/zpkv3cLmwbnIqikIP0GTS5bHuZWsmEeOf6HEsXG/95rYBVo9eV11uE8Y1
g+/5lYoWbFF8ztfwxzV3MPsEzfpKwCMSue/5OQ3GIX5BLQNevCETxc0VDpDeZrtH
XsyrsCxODgC3QLCIkXMw9GgI0ZoPBk+m3hnPOZqzlODwyr6aygJnJO0DgR48f3pp
pGHQAPhzVbOoP/mco5AZq6GoGhkoKJpkDLbj56Rcsk7DnWRlnsP5TdaZwv/Bi3uz
l1njgWCe17e8f/Cdx00bSqj8KqsJeYBh4Eqd9gG1QNSkLC9dRppDji/qOzHc00Tt
Reclokvo4RVTQWzUK6ZKKasvuK8sn5dRsouk91zoRKFXlnAUHmiBr5Uf6BOvqsAf
cCeuIHSbqXfbTypqQgO/vi4ldw4quRXzxkcbarc6JAc8Jj11m91V0ygabQX1JEkc
bTqjqCii9nD/PGrWm/IuNKQly7kidFPK84peTcqGy+uQVZwTMgTBFiWstD+08j7k
Plzi7E3mB3biwDpnyxywAQ/WPcR7GuIntUCT2ZSexJeOQ1NJGGXuCaLTa6GPTBIo
M92E4nd0lEfhprN9j81R69K1AUS7fyky0pyjc/LpuXa0BnyP5YXzW4XVjgFeMa8u
Ga3pDFcl6BhT1NWneANC3MZsSUpB6YL1SnruUAejimK21wT61eE1to/7hbE4LcDV
FLhtbn1DocsoO4qhSfHJTDk1G/0oWJiNqBHfdFzpOKeUtvRGYN893DYU5Y+R5LSb
rvhmn9Cy9adZz91yxxaEctOOpLt4BNUbBz52c9IAwE8+veF+PZAf46tuXUH9wCU4
Bd/Cku5JyfTUKS7eD87hlLMhAY1kLZAsrXws2RrmNQ5cEt2jctHYDqDfX1MQTEIG
8wfVwWmKmqBaYxVHGb9SeXtf6//T65VTzARZuzZ9KUOEX6xnSoUujlSlQXugbnoK
EQRoGeQQKBxcbEC7ggBqVmkGFfto1oxvA90rJolBWbwpvG+ekTazLQosTOk72Ctc
5DJnFfwiVRvM91cQnu0ZpcLsFHbgrxZ/by5BZL5gMZDSj45cd+SIWDhIEc5A/vG+
TnccXluN0wmCEt/itGk9IVTY/cR64jKwjl1KM7PXWgBMzF/fXT9qOhSv2Uxqmzby
DG9k6rEPuWZKgMLh0BkmfipcAat7JVBeFT4b7tWj/2AAE4rVrgMb5HNWaakofneM
RR9zx2t2zVdaIgklR1ce2K2BmTFS3mesIdwx0s9tw1RvehgWz2vu/WqaSKCdnn3R
koTbMn81yq/pnhTyBHStue1yp1TL8Tp44lOj/KJrzhG8FlXWI3mF21B2d+e3IVBz
yN9Brpx4RGVljXVaFjyqdzG4NZYGI/Bh6dxGi8vFLFxYKCcFlnDj81fIZNsEzLdP
LeImJw8O/ff77essD9do+XEhvuxVrwu0us5ygb4siXJrhIJyVXiMof5J87HQsKb5
Vq6tpO9olIw2xOrfQV2IwJL9C5aD7YhiF8frZkK9NmIkoecLnqkfIUVI9kfONkC+
5WnqwLWn/c6F61SMnXn3dHZUqjFABmGY/y60habuza5mEvghYkR1MgkOqhXduNFR
62kk0VaVX3LgL8Xok+YbXAhWogGC9QC3Or0NVfP8I3BRhgQdKiacJZoibas36Pow
R7Jn9PVs4uN8BZabZXeOS6Y2yao5vy4FXaVSKxuTk4UZYXGb3vT+D7TP85USDSSf
TxCJt6TihGvKLv+TFYow436ivEZ7yezrE6VFJTvWkTzbYvnp6QALryPIr3DHtklg
3WyzviZ8bnVMPXClfpJXCjrlvvSfn1N0vj/Z2MfY3ONOSdsYfRtg5djjuKXnv85l
5L5ZG3mDhHQGanj9XCK6okj7xhrWsvRm8CLifTmGR38hEuwY9+3fA+F5jTx5MGZQ
HNnRQ8tCvCbUUZV4Fds+Q8neDxEHmKSSgIBiYO4W5mk2GsVTvtNx3c5V+2lw428s
59IJvFXGb+qJiPt+tZ+qpzcgbJmN6GrFMuBEYoW+artY009Jtzxwhi8GtrOeqa4W
QECZ5NRNIPIzGTNSkxz9DMQt+f63KmeRcTxMQBumTd6monO25Uwi2XfnTGK5sGWw
C8t+ggDSSg0yhn7pTHsJPo0GLg5c4rerwv4p/WkL3PLqDD9cftPsOXFaFbKc7s+o
AEYM6u9GPrkSS5vpwaOR697QQGydLil2SfNmotfrbX4BQ8j4ExrONkUUl6bqBEyT
X4nq6RmGZRrBKP/MXoyZmqozYm293WdMuO87bD+STUNKVpqo/K6kq2ks8HzxEkm+
FMq4Gm5NmHLV8M5mpd6NzsDm6DbXOZSxl2qaQKIjSjDRf4O4raHivGmmiqVGu+bd
XXXW9bJCKe+WOsj1GpB56f1Y0476XllPvboGkXZMG9RtNdP80BDKegFDs80uGi24
3r+vYZhngszgx3gYaeO+pNfAJJlT2KuHUVXciyWl0uqZfyXZ8CMKZ0WnxPqcl2d2
1NfWWPL0Uw/Kj2Sg6cHurD72nhBwbtECLOu08JTlRpzKB1DU9gjECq1qL9HMJ484
yPiUIav3rnpTtnUJEAiMfjADGSdowN7UijdzAQGtnFz4le1HKmASGCyBC4YQR24X
ulksmgFAQm2QLdckc/Hfo2cjYy+bkeJ30w1Br3cZs4woWr9JPAv7wLLyRLVbGRaH
/d8rKhkdy3WaPQEs9+eS44VTOJ+4Dt7blsFHFulTTC1nSfi4mCS9iVcyjjvtXTPz
ReycELONmj9YKyn9rqnv0iCr5l/pQvvvlrK0332BqNDSmpmFerFAbCHaz/0K6+e7
0sOcg+Q0FEwvMgfcocnxJwdWST8B+2O7k8MzzjIfuNhW3NpUthrDT/q5e5ibey7/
+NT5aKd8ou5XA19qV3H+4SItjLfOsdxjFb1y+EZR+p/TPNlX3CbxWfBrvfdzdUlS
jrwLgf+0Th53CbrH4UxoLklHgujA74MSdum4UUWQdTM5sFobyXfcIAI77I2f1LVF
y0qzV8xzQyPH74mLF01OK0JGzum6wbmQfmlQHo6Gu+/0AwnXZ8EyO3/WTtEzwjYv
jtu1uSALbL4UYSifpoKrXrDZHqiv9uJU6YJY4T+4q5p9IYUmhXgyXq2LQsFNUms8
hSVaHGXLnvSTN9wgH/1WcsojmU7eEUaZ4MDSMgX67qpVcx9zpDz+B8TKLIFNYTez
5DBHsJL44ZETn3N6hwa/7+c46LZAJbTwcvYz9McNAxpOPR/Ytph4316y828oYkq+
8T5qNG0RTdvvipdrYuA2RvXM2udeAVJ2+JbcA5tWDyyBDONrMaglgM/Xc51z4CPm
7sqxLRhhRlWLGP66u8VE9vDPvpXSAeeH3hAv7DBtiHS6y2nmmjVQ2Oex5MPvNFrc
fbyuVftoX736ApbthcB16KotrwnJd57yhtCC2a1m/cJ9h6ymqQGtUF++Enr2Lrgz
+QWEoYz4kxK63PASpNiWkXdeOlsPrvL0EbLXODMYSbl98Kc4RWD6lQo4uuZ4P0ig
nBG9VnpzTiOaYl5cy0XFE/9MaLoqS97I9Jucd3zmUPCg4Pl6JfX910sVxKc4vBVb
zRJ3qarRYTw5u8NHqJYaWhQ6C0rUtWBRajMAk2iCJ3uSTHJ7WwwSkuw+IOgB/zPu
NtXozW8USNrKPJqxDP9y2GZf+3idU2dixM2ciTo7fwHafQ99c3UC/kItU/k6Fbht
38fdPo4dUQqU2bQL3BGJJvfoKRMQmTusrl1cPYs2/M0LV5XYMuhCVwL2Nd0J0DV/
hhA+0nbuJhR2YXOIFAiZ/jZBTQQ+guTD7CGGJ3J3MqLA3KGGGlQRWZtFk/Y8cB2S
lT8lJJkw95RyG/ie9dkhe/fXnqWIzCJar3oy6RdSi7dO6yjI0vd/3kNmddqPHUy0
6fGS+PDEtE0Qh0OWcUOhdOTGjVNpKdrxrUeCPgdimosXSpg+9Lwwl8EgphcgL7wM
jO69pAve2XeH0S6LNOXMUM0hmHUL+Ta3TeOXcAsGkuNu+yx6M8b/rZGQ60vYs25n
cHziKog0FgBuFdMXL7uBj55nns9WP+JQAClDWBXA3OqaqZxWoMuhgCvucW8kUkfU
Tzz2vmWQizFlVu+8zEJN18qjdZyYYUNZXuwe1voW3ZerKap3rTmF0klwCrNHq3ds
uYvURuKm0gzQpGGaaOt6bV+dvq90uEcwPJWnNtgXB1pGCxmnJtunStpo0Rk8wM5o
FeGwdc+fjFR8Gho/gNTF9xQc0BQBAKBlhpefIFrO3j1I/fDiIi+9Nt8N6f88J9iI
/ph5Ylz4tHGcvh1XSBrWpR8bDE/8AiYu9m8Zjvf2y2wdw/wKuK34F9kmIVFrgGmZ
QCAPjyg4O91Fz3F8CppPgZ5y7QOcMYffcQXorPPdDbikJaGB5R12qFEAGdDATwFj
WSKJgZYpg/PCV2S6njLxiapnYFFMdGy5viDJVIyA/tCNwMOmhYnr6Cr/uP9ftL7o
FQwsQxOjkQN0cS3/TtrtL/PsO4PDnNWwMw0ih5LQKGbCl4D87Im2FBr/1wT/4JNj
dLXmuytlNXQLyqECcO94t+Af51JBy08V58+8YFTbV7wJKKhsjIz5+EBPsECAqKTn
pzz3Qjhj7jy2I2vt+O00o8smidA4hRy4YUDWUFWPvX+QBNkOQ7LUsvIKSSg7QVlu
2Fgm5FPGqQixThPClimCdiGySlbE/oZYJPd90KgvbZYBy6RvK2i0XAMuCn9USCcK
4/hFuZZ7TnaUBpH3EmmITxnYW6hwjtjWXEw9DzYGq4OQni4bZnXRSupLOpz5Js5g
PcnQnCAEmTjv3DRo351aLnyf5M+IMoXyQguhmRZnnG1OLXF+NZf1pqVHoQCf5HGo
KNXTYzY56VgrcR/BiqEYxlD84uaSp1uGacPH/8b6164gd104tNKsFUJhEL7Gd7MA
K0mvz9A9MXrop5N0y5aVOhESaJiVqk//JEBrhNzOGtcRKWY5bp6rMlLGLJmlzGMr
Da2lnuv6ejNWvasDNQoi/AbRGd3tv8GPegiXNDgzikcVXt9MVum5zKVj5sLwshuH
jGUMk+xqXDoUnjKGdLbR1AJXNEAHUp6ngMOvbpeaM45EATlEh0DPiT+XDy9YORc1
abi2bDIffN7vCoel4f773++YVvUXdpB/WInacLFDtykAStUZ45pbkco9IZHYPXxy
yZN9KOgEOzniEJMHPZ2sYZUCv7Q4oz3SeZrNVnH9xO2D3Sr8idBLTCuZbEo8cLlR
wuPQiZv+arGcjcJk3H3hB/L9J0mNeqsF/SsFFAqMtf8valoCoDD+2y8UKo2Agl4c
hA/8ZmckZcYMpf2e/ZdVhTTaUI4Xrltgli3oXxOHQwe6WBkg9rnKS86U6WyoPbNQ
mN5KnKuyxsrbWCnZI68DZDOP8lUQc8gpl3Qlb1BlQAA6X8OM/VEWjPBfdp4zz7/L
6G28l4/hBXeaRAgL9I9gGu+Q4Jy5ClXy2bDdZNOU4U7OGz/1VAMdd3QQgTnvRJqq
/h/+ksUGZqOedV/zLm/4EZBLGPVmCaYTdLcsRcjVJNCkzJ26w5SCc3Hn105meBSg
HJTO2QtUuKUR1Ee4aurJgaR3wb5UFnmP+iZ6pcY2WZ4G0HLrBfwHXbNV2HTshhjE
jjprnklLGldK6SIksbfsizegdFEHdM4xxUJ/poQyNXsQ0cxEMd/U6XeIxkkEDf1Z
bsKLAMZJZGtIM0nrd1sBA7QY7Mgy+eu/tkaCIbUf1/SMAhyuz0SWrMeq7rH3baQe
1+i3w5xDZGHHZunb1pAGXMeXsyfr74YXHFHSQeLn7KhuCycgacZ4t4y8/7h6xOtz
4uE/9f597akRS425cKiKW0TGlBvn5ZzdJiwe45nYZad2IDxnFjuG06GHiV37Xl+w
sEHYlOjK0F2wjVzbERZWiPtvP1nfTl3xHnjGw1niVuKqC9l9A9w+NPfvFFB+oUtR
+4bMJbHXmhZknMAvgDNvAWuG4ecToe4gy7YS7Pe/7ZylxUZMfRSgplZb2X30hur4
oieUhf2CBX6jZztIgjkRxMaErZQniG1hUr97kikggzNUom8oKxQ/Ous6U+k9PAt7
1c6IjF+AJeKQDZ4bm1ZOoqBqXOhBu2fHjjWj1tfB1KPvLZTncIWeqDLR+p0ovm67
dmt3a54xEwDYNxehDrmnjdyYtMDA5QddUyYMjqTgZtIUOn1DHi+TEs7uTxizQ43T
gZsXVzaX171Bi6SvF1Ue8OR4EiiwEGLhIJxTIi7HLVbEGHXCUWsTHi2U4B6Rx9TM
Ab6Q46k95pTNSFcWgZYYj4Cvbc7tPp6ZeVMxZ3fuq0KlWfGNQ3zOWazJcbpCzvVs
eR4Xc0JZH+tvLi3CACJXTg/twOTVIPkhTIroJNL0KzYh2n6fZpU1ja8z9afq2Vcr
8oNIMZuuXNJ2+kK+hMnN/0CdAdFSvehTfzc+EzEOK2SjF+Z6SevCnJ1XjmJvj0um
m8mJemY8CswSFyzpwGFedzh+I7PihJcuDJMe5m7Brbi+wI9nWFWX3p5zEYd36880
9QZoZiBfL5PbxNKtHkbbzclJxH0sizE9MqCa+bs2ct+JUejZLRGg+trKuFwDxWYD
q0YwcULKENmYMqOCAS/6LSVb8itgYlE7vXBVSevcBGj+sdCvPwBjBDOISvHJLetx
cad8fcW2ob0DMY4eEinEJNmhP5w6dUmBYTIJMko2APHn6Fgb2aHhVSTRi1qK0Uz3
RsKMvBMZ2QeRhxL0OBCfJsIoUa/n8x/VdGagFaOJq8VM2/dMcXekCUXG1LZW46LX
WKgpzUsEjPKWSZmpTMUwaRh5mAkN7w1A4OhthkRzw7K8hiY2eIJ5R3GPuQhKMpX/
yU7SFio+ZspGaK9I7dlMm9ApW0S5TQsjmFHG/VWOygheA6UOS+mEOh6jxY87vC5R
kAR0AceTnovoyJi30voG9seRgeiG8iIuu/1z2yCQbkxOyqFl9A/tfqlqGCo43IPl
83XQzfSAA6fh7iUjUxylnmgifKT+bkIIjVrtaq69Ob4WWdfiSeHdUasrVkQy6Soo
OfeM54I7ElHGMTOKcaiqDSev4hBmCaQzqkuoUN48koF80RIYk6nU0HRH0Z1qr9R4
BUqY8wn9QkXHYz3kNJNwAsQf1b/RMoqwYQPaU9vt8RMuY219q7NXkp9NTjnen7Be
BseWmZ20TFvZwvbXWfiORUJy7mblevpzjPzv/AWY0qp5MyN5h40ibc7Bkc3JvDLo
iZVBhOwlmi1J1M+jxUKI+CZRUU0QYX1s+38XGhs56YohXJ6NkmjtgZFB6SvQDDX+
tG/HONCrdj7RI7eY74hSHlo7bOkNbLTi2VKtVmnWGAYDfXR1dWSUzVzr4M3ttGQX
U9qbX1zR4vvl2wImCr8HQFSnfbpSgzpSGZTuXfz7bJzN1QzaJ0r7HSlPk4GNDBmC
JbT2sz8BTOeM2pmzuP1CJ20KNHZS52NJIDFC3uD+c4SRA7xTf60gkQJkgQcE0jeC
wUAtPQVUS2uec4ttXUHuoO/N2payCxQp/UYxq7YsqVgo6DQjLH/p4Oz4RM+EvGvR
U2tHaFwegNzkRRCQrao7n3tfG0PayMwzcR/zu/H+z7thoLBYOBPvnGgsukZKZ4Hc
Zc5ChpLf+mzQxkfLqLJuS2FiwhuttPLdYW5OOAnwuIP0jUiGzESv6R2VvC9h1S1H
XxDxtN4nmJkmLWak+FlSIepjjQ0UGcaY8gntFXi9Pp0HkDNluZX8Xucq82EiVLaC
LqjkkF4Pa7xgx8ueyKVgMHA+INlFH/AfKkwispgKLz4hqqUyLXDB7p1t47KPQcbd
8wLDqmGLZwqw1VwReWvGZVt+AhjLZjiliJVVnYm7zwhXY93gWUNqiGZOzlPu+Oth
4ycd+Zz+17NgjnvNjtpcVXHNdLQWAwBQocnE2OI6sBcd8OyoTNJUGZ8I0bdVESWC
s5adRYEgQ55UTbuU1SwloHFTfFPpb4fAT4ClgqsbwdY4aiTc7R9gUxPKgxnxU1Lu
xASQpRTS9YCbElwEfErw6R2fwkdrRp56EtI3Rc6UfVrTLPz1K4apkQjWL/Dr1OaQ
q9YZVkfAB8Ky7dIX/9Rv2PZXUsb+bv81+FrGLDtVFIEUKE9OjfX0DLBC6Mj8LNF9
9gsk346nBtXumFhcVVT+pgLk3k6Xz1VQ6qTQbVs/+GKaI3Et1ZeRrVWpVs9930jO
PH+7FnhKWUFFYHLcV0YrJvQ5oQSdcDbCWhcmWGkcxSS5BuPumQnmhOtDi+f9EbA6
wxeTBUKJh3sKsrj1AxXzoTgkSKpBMijDrDraHLI/8kO5nAiz2dJ92kPl9/PM8T+b
9NFehpqyNttHmhZkddxFXdm2DOZ+QJ5o6Aw7PcJgZ9lLaiocpnN4NJ3AyvGMQbPt
bZk1NV3nyLNStBIrBPttUsnNKMra9iWNZZG4mvdfesIufY+cT7VuHS9gmsZWenEf
xOL5lzNVvzSCo1rvURlJr2GnZgXd7iFXxvqzCUSaTiqG4DEn62Y3L5IRW03Qo2j1
9LevNZm99rkofpfgefyxQ0eKet74DENsPz5PGnaUR2NEkRBVvrUHpxQpL3sFUXSc
lK8Blozfj7OFXb0V23yzojFvAf4pPPKQFyRJe9B20Hu5F60AYO2hWqDS+0QaqoxR
hg1WMnsjgJnNltaeppDivY/1KCLdCuw+9fFD+Ie9oTjQNSyb2f5A/MpnR1vCiDZ8
P8eXe25sbiLYvP/36MdgK+JDVhwQGge1H+/Y+EcRN8RgB52cr4556F5bkzkT1fAD
APE0GdpMUlW6KcVZXCGeQBZ/v9xbulG9Z21XHtr4KAs2yypkWoNkqto0CXODmxXJ
KtySCTJ2GYGIag9p/Vv+dozDy2pKQxTtdQmmiHDufK9S5SinZI6L1jYcEJwqw1wx
o8DPwBwB9+nIKD6N5stldLa6TW8XMp4Cz2/48wTdScxG8lTMlEYUbFwg9kf7qXYA
8QYMvZWjO7qo5jiT56TCm/p29qgO/AQlY401VjV14nkuUskE+TwfTJP/QzMOedeM
cUk/wtsThqYvhUMisw/K7ue1wcHtiGQbCvXHjKA/BzDDUcBYlrJXh+VHtD2DbN4X
BoLI8buorJeJTuPSO+jFcOqBDlvtcSTF7gKe09nuUq+Ch+LEsLVHo3ewDRy6LVv3
SKa2a9Ioeoh7Q3uV94CT8Y0CMWBhn4gyGrEUOV2g8+QEIbCOdjKsIml0IJypTvum
ZGiZHTwZFA89BqGVxBQjcw5Dk2gUY0iQN1bQrIx0kNvR3McM/B0kMlJfgiJL0BPx
kuLovAHePkt+9lfdzmIuy/vqcrtXu9/sKWlqupuar2/YQXc0I/3A2zY4Cmo1RfOY
W5qLXuOt7cM0NwR/qVYliToqvuB42GkVIat4PwUFqNyqn5CnXom3J3WaAdhkXvDn
1TjQKNpjgYH4/11BPCMUV1bdv7yZCxmadJ/tArRweUXKil3KqVp1ITZY587zlNqM
Wb9xLxvLAWsCTJwd/Ih893e3Pu+16HRMCewrsPYdCbJarKDfjhlc48cqVEr6zX2a
d/cPHlC3no2hkvaepNOpOKri+Je6L+QeHEdc/ZxDGkvYDznyJME5nr+1lJGdi1rT
6Hgea6XDqlIesGlsvr3CzDH2bPtaFEbf9GZSrO/wNG7B/pf3bd6MKo4IurXI6uTb
MAg+8XJ1epCh5MAs3BtKEEllckSAfBIl2DXSJGaQOObpRW2tDRel4ovQdp0RWeFP
Nb1vjjFMwCOB4irSRFIeFI3OFkBUEGqoVJhNs9ysD+fQ1ABOoPn9I68Rqvtlh+7p
CWJYFJjR7H2aNK0v2oncWWEMBiizY5FJ34ZiHuAtcLM53JIkDmmvbp5hPpc2Qb2G
Hipb97ay8xCbENz4Tr60jLoi29oaNcvIzP1mE6oJC9vkzGvJM8bHJWGlwzt5sY27
o6qrv82+ZS5vGLI7UrKxSwzL6Nh37A1kfvHtOhUmxB2Hic09SO4YzYvXBNfMqx46
qtS43fWul7n6CL0y/OIxD9ECwi1BccKyCbGRkmgABqofisht6pz9lRtQuvdXyrwp
PBiXs3Hx8D/LW6elONBdK2LZV0RFdwX2sqXsEHaPQP5hiptbOUopFacN6ujqrO+7
JB5Z5mXSdbePrBfvuSxaGJEUAcn71faRQOt/sh/fydMI/5rdbFctZSaUruZh4EFC
FYDUKxDbnRW3C2McaeGKRB9RazOI2gOlTfe2oNeqE2lvW/r6iaxqNr54Rqdscq22
Wm3f5zOtVWXdkGjNlgV398M8bzGy6RyOgTO8HCvI7mX8rT9C/8yS/yQUZpwd4sed
cSp+zUtCfP7dGD1qcav2zmwGU8x/VBskzgVrmxytuYQnNgR7KwnCJncVB2YHIHxK
VcU40Z6hIwDdgPdYGzedTzrAODJ1genjNdAC+fbjsaGtm6xQ+q4PKz7py4ZMNtnV
Bs07S6WwWbh6a6iLDwbbzOBRVgXnnUHqk/wUIOQD2XAPSeklCd5i70jrbKfZJvof
fh46TIuY14nTfQqIKEgq0bcbnIqZhrcfo7fXNcUXPedeCMIRauoMxRMiw9GauvJv
l+Y6y5u7rYQPBcHHbzXQhojRtwnrM5bzpP9XiClXsJ1AR8PElNQURyx6rCFeLUbi
5L68/gSRhpi+50NpLMFu9vQeSaNG0H1+dtawFhfpLD0NKBctn7BO4BoXHiQTcY4v
8BymQtHsO1xo6Lamr87bm5stlLNs83/rJFdr2ji4UhONsfm7aYmCtCLw6cRYftGc
3hcQ1TaDJp4oPkB8wItG/tdGw1alYHEHQNvtx1m66H1LSTcIuVa1p8ONfQRWjoaZ
lreq9Wj8UK5WQPf5pQdM8NlslkljybigdCskwUXBUXBjVlHxdBdyPgqEJe9Wx9rB
wgjw2RQbKLunqw3wa1yHC+f7H69PvKN2vCnpsfFQGh+f2Q7WbySUHAvISYWTHSIk
HQ6R8MrK2OMRsvjf5uZIrG33x9SOgUYrlsDcJu+mEQwgTcGPzKoCxmI6UOMoMgoh
ksXbKPjZKxwd+l3zT2+NkXLR3APhB/dipNFzpEFHrXdJsTjgVG8VAYgJ1syoEtO7
loI/PYkBQbJHa3YGVAtFdFNF68mNtJYcVUeOVXdGzZ8OdKkehOkB4dN2veR1qHmg
dTJlph8suev2dhej/pI8BKX57kULK8FdjJ07xqpk2+eS9Zb5KtVeNXfVpA+036YK
s7H/Gobp6flWYXiUi/VtTPXlUeEKvoFrPRtSOB3g1sdnWttU5KJEBnw/7nkYt1+c
GXapx7CuCd11fmvKUhtEba3mWqgApend30MncR/78YosUX4ZAcMkwxqlxOMPeE3M
xX9CzsgKVXWLEe3gUxELz5wxnXSrDF0YnyIExgLd8rmYge/5xnlf40A1B4P4cx7i
gggbtPTqYR79ZseP1E+oWcAiRcy2lC/go1XvWfv8Mw2UjmeZ/r3ItSpmHuCKLsJg
pzlTJtyPtCrlcg18sCd0zsX/0CGEHUzkZT8JadJ91isU7wn3oWcTL+7J/ba2+o+n
7UDAvF/z9U+JEbGQ4QF4OmZ5KhZNnyXStw3PkKR8mfBnaL6gQBbK0SdumUbR6MsP
Unop598uwcDXCxsPJNqS4gG5kSDyvYhIaVpjmLbvmHwojGUUOCfUs9uZDguIHObr
a88M+QlkC7aJuXkkSYQotznyFucsqWI6evSP0d1mWdjFuYWj+SkxPcVd/NpiUuB9
JZD4PQux0YvvT7lJAZt7Pu9NQKDzYDwZgvzyMUpwXUZLMnNS+GCYxqOJmbtsmvbX
PapGBrTRqiDdLSEPbfEVCbTO/3xh9XbeIh15o5tQbpwhd0z8lf6YIOeiPXzrnt2j
GYVNIkM1JLzQogxSDh6qNa9Cl0biHM6X4dvTgrxKqENuD+ah9Wve+V1KwuX/Frdi
DMMgLUl4x2ZKnOlWjTWihoySmd6tn1nQ7tMCkNY3OrOZQuirq8fnU794sBUlYC6R
mlDihnJM+/gu6aGDxve4KomK8/4aSE4wjM/caCXMyQls8Yel4OXX9b44J1hNCEP8
btp3j8QZpXmId8bhPgFCiTOU+nVFMrW2VbNNeoXOrlk1SxzWZTPEId6KBXKZeX8h
teTfejbBFE0ZQnfybJvkWwUpW1Q2OEbWP9ASVYAOvQFQsjp0wBGzjR6LGjZ7ygXe
zpbCbA7ye93LAYzJELk82tBc7kVqCELsCyX3sIu11T3DFnR8S9ZSxOvGediSHOOA
mOSFSwacx/HsX1KN29mB4exWJrDk91UihvnAUOMB2WPE+vSi02YqpkloOXPqaoCQ
xtiFSiImtDuWc6cSUAdY4GQyOYRAO7h3vm2LCJbxl6fHyvYh6h0EiDYM/nHUC1GH
MKdKcSVNcuFcFaRnYCcG6okV9zjXxe3mIuy1/UlLQR8zb5iIefCzSKJxM1Z4W+C1
+NyZheT6ndIzxX9ydUmBpijhzbTYx5TOJbrNuFGiVASvQ4Boh7jw+1FnlAnbmRdM
whyzWcqhyIxVqIcNW3Lzx9TFWChsvlNM6VM85QW7R0BpjZkhaSlSJoat/EZfN+21
qyqKeTSljXbxaUdN2N6RnPb6t8zePl/7lBDHI32KUT44DuN4bnfAveKu6opRIeU5
wiNuIkOxJHe+mR4MtoYmB8OQq/bHCr820hqgDnomLU/NVAe6jo1RkTnroSwOZRko
ZB1jLLxZyizSwfqLB+ttOI5l3SLrX9CGXatN5em7Ad68kEewp8lVc++9OSpzSnNP
IfgYuAfwvxJVk7HBOBTJA6aCOfVljdDYseCXBIiLTQyi2amxAN4u7ABNkfQ/H+K3
ZdnFMEky0oHOObJUuT9sVl1qhEUCnjESFnbY9F4nSzsoqjlYL2GjKRVQp7au/OiU
VZALjiLViIVXG3/TIEJW1Ukc5ceOdv5HaYcZGF+NLe8q/7EKR4cK1mDAeWMov3Lv
0kdI8xY1eVmO8e77GTWvUoGva7h1c1wBbPFf8/z9HFOlXAuCE5VAfYf/1LI56hUk
70M762aQY4Yx1fZvJPDTIno6Mm41V1VSSN0ZZ8avht+BMSMHfHle4d05fOIslfl3
iEsCxB2sYELc5PXYWXAj92N/Z7KNyfIf58VUCJCyPP+daxQM6vkazjcTNTmpMdaE
BZWi1z0T0l+8W1K9Qz2CvZ43jrnJe3bqjwPslFrjT45mDH3T+tdWiCwm+MP6j5Su
Wz/wn8qAWAgpMyWc7AYmxxnjfjcWbn32BafbRBMJbsHRlRkYSdxu/Jr1R6G+lODh
WCi0hAMCNQDBFqfDgTJPQTIdSxMRmLKu/NlQrS+mAqHSrRQtidqZc8GLVdJPWIWX
fziEL3fN+zEohKx3ZIHxL3czdImis/eAnn4Sv5i9yWehthixaTeIF0/Gum3yAy43
GGp4ffT9P6MZyOmOXLyepOZO7x3YWNO25gGmLcC+PhNPx0LWVKH3cWklVNNm1LVL
r79s4K3XQHL2aLLDdKlKEg9rjc/lyMSEFxl1c+o1T6iYaXp591x+yEBVWsXC0x+g
VT5cMwKsycpxDkurh5ZHhvHsS3YqiTP72xBHtdN57DsM+sYBAwQsE0yXobpf1ZC+
IqxgxYtzQwgVQ2DEMLHcqBpEPIVgNjILSx22VeCpv7m+fY1TeTOrh+vNG6L96prZ
Tz0yOaiP/XJxaqgOzDrRdkRUjQnBvvVYFMVjnglzT5nANqLYG5DOL3d2oDKBpuKf
zswc1hFTF2oE3bjfci3LQ4duUjJJIf9FzZBqGQPjJvIwGUs0KZA1031HZlcwveYT
HuXShqDtMfPeurTPyev27X8h0oAbOfnjILRyZrzE8uybvA0/zY+DTk/fg+tSqSPH
PZON6LEodAytFjP2YZPCMdXGylaWRYLWn94zEs8vPoynI81sAkQBZP9tWP5ufAwu
G5n6ulfSr7Ix6OqsS6KG2+IfQ5bXScLFbTn/uRg4hLCpkkbNm8Qmw5SnEi7s20ql
vuSGQK97mKUMMdL1cycrEy2N2ZXBdv36OXE4d5lEJgrEcmc9y/WUz30AlXYP6wAc
1ggn/XiN01AGpA7cXo6YZJJSDaQF++Nea8I7ALhjl4sXz5E9n9VlZeNz8+ngHyMT
57//xe7aQhPi6+XSzoNFY2s4C2/oAAb60ar/KQevrobMD/h9R09gy5rd1Gklv2xg
p9Kf2Y3cFB1G4X8R9u00xtFJuBVbu/j5aeq75sAQ+2E6jvhWIno16M9JKb7NCbjg
F5j/4LHDSGFSDFLCqjo6crOOJ8YVPyfpfWAMxRhYTcXiQmEOeHsMB9RQzITbsSWW
VcNdOoZ5dmek57n6loMqbPcaWVtYTsm4vCaZINw1MZvpL4AJvpsJRj2vXKnJb9oG
E7bhBGiF7dkniGnu7c/oScuAgrd4zjNLBtHLI7hhyjmbyUojfrm32OnmzBzQ212l
R/fWDzG6sxW53+HPfVBVvVDFXVw7MtOnQhs4kNGR9iTLtI5oxwStepu/W1frcdxw
Mo6ZYeetDXS2RnBzJGKDBpkgDxwrcg9ZaYTXDUFTDRmh5uhFBnrrRo/rBz4MS/vc
+gr0DlB0xYZR8sUKszW/0/l/3NZMPqWemM4GdwxVQoEgWpLV2TOUESWYZ67ShKBn
n1yTUuXzfT0fr+x127gI161Zwdo/AdLGvJpP9KsI7yDqW521fK7SUt9/F0GK95YN
6sj2189UGHeTzGgxMkgiver0khgmaCevkL1Pv0PB9dcRkQtTWbe7xyFpgB43qGPm
dlqrvPOS3DrQDiPaH/PjYhZiIVHpFVYOCakYb0/zLYL1hbmxg9/5nG1KHxAHK/Oq
621IqR4BhStxumjpYLPXTg53eJPERTSw6y4Y+x//1L36arRh+S5ciedUSlgQ8uRE
v8btIXxGgzlR3+QxG8vH3DUgAQmhTN8wjerb9o/gEEsgeYxoGss3GU9582E9dlAh
0tALg5n3wA6KOfO83PLC+0PQ7Ni3xxsf1Kd69e99qWK++8od5SSU/ZoxU+4RYFy+
2c+DLLvg/3ENG2i9umv8AAxdlebuAwhbhX372DHhXkg/eSNd2bc829WI2UYgnQk+
sMdskxsYlvKmJXlgr8b+h5oTpXU/HwRg/r+Gbul8exGdolGNTign9C5BYno2rhNn
YiZOk14974ac0SpcIPlcUGA/IDfQro5Rcnagc0lS3fuq+eCWmD8tvh0ZtkwHr/Pc
mdy8dtrJuS96yNiJaE88OlJJVQl2QX+7zBddxZWdjQdK3MdVKN5Sc6wjYfsRNZYT
86HIU+4WD1xnL0dsw1VUNznHlabJYhsN09y8jz/VNGcS84ZWiB4XYM0210Iteu0a
8CaAgn0hmW3BcljL8FhqLUguF0U3R8qblDJxWOC66XWAOQm/i8EOvWOxP0QRCSKm
tTzD1NqVMnkcRruFeVem+dP9JEnB0YZY7ZXYKtITJOIS51eOUR6/KePHZTfcycQW
i//OVdDNbq5A7V+EJDVQy004mDqdHMCHe0vL4TLAyrbHo+Ex3phq0v0e12WCIgql
grrvkowB5ZUfNkwN0GlSqNaBJQWtQ4wnWAN7hOFKRSIutWllIdwgZzKtJANOLCuQ
AO6ZLydK4MMTsVMG8CvdY0RhvbhKQwR/SVvhKj+2PGyx+P9qEBhL60D+azME30Dx
I9pY/zeQxGDo/yY7iBGiDNaqcW6gAnWMjplsUWbDs9ZKlNZkwB+eGiUghTmkNiVI
kwkXWWnNToHjaVwCO47N10rm1gzrMCR9r9j+QT5noruwTcho0ldn+xC6Nq60TBRp
0cy24vi/je7AXXs+eGDV/o7bDDIVUFUHVeJiU+mmazjp1TKqhs7muCwaCyN5vu2n
f6gLDaFIRcNPd+Nl5DiTPuTSasYyjN47/48pk+GBdoqZjEmS3UuUL7XDik9Kk4pQ
NVNsk+hW9upMwgo85VrMy9NQgPh6ubqdf7PPVdPIKWPCIbcwpkuwDI9pV95+for4
rLqdF99Wc+T+0Fpz6Z7qKdBbjRKPg+RZ/CHxleadCdDVUQ4vJ2d3JnJrxOuWRBn0
FX8yd2UwFMUvRsPg63qvJnQOWrOAQpJBUIZz3NLC8LI+oR8jcr5iAtoZNSe7D/F7
kc2ADsn2egbN7oVjNBSXcaDv/juC6huiIqrMweIX7Qo7lejxROgd4uboDEWFoVGa
g2HV5f3RI36rcHyLb/Tp2OCCY/qZrdHRS6SH0quJyjGiPRrF2o+hbGLaAgbpq9t0
xo8umI9CAOmf4YBSY1zUGyhVpePqmPE4xZO0wUR1rfMF2Y7KkWL3baOhzbRMP+hr
hf+rNM2trJvR9v01zIlxEqkc6+0cGh9iNeXXfHUXyrZx5n1Bw2bYlypnzHpa6AE4
lDNLN0czo2RfEn6XGxG4S6KMZ8lG9svcCYRlRxNguHXuMa/f+g1G+ausmnSnT+oa
u++ZLvat5aHOKGc8d+X8pCM5jPtibZHAixIocaAz932z5jXn/T52+S/j8cGLGJSZ
NDP09Q3+oh4X+DlXgTUkMHiobjUgIFtsttFpiOrRxD60JVmUOlXdfev+taBJag9U
uh45i6d9c0LzSzJOrbceSGbeUiJTrdIOVn9s20e3gt/+qyGYfvfOOdKFnwwtbBPk
teKG6BsZ37N9oLuXqrpWxxUumih/7cVop80jSC5BMl+lMLGkejiDCvv02UMXAr6b
faxgQVYcNen7eAMCgpU0VDMNLLOGMltu/nMmh7Ctq08htGhZIeCEsHXK4CrnBR5p
8HlMz84fL+jB1graF37Q72so5UTPV3FDD1n6/5Aevuy8ENlbWudEZC9vQ1+dcVk3
ZoCQm5+/Lt6UeDPoL6x2oR8OyYM+9BoH9LQxY9Jn0wEdJQom6eiywmBZRb83fJfd
3cRp7A06bwJxVP33e+frmD84ha9XKoV9BV3NGm1ofamLwu1gB6S8b3gzwl3jxG/v
JZ8A4P/L3Px4JHs+jM78cid0PLnM98ppGErMpqjXUjeaP9CD/gRDgLBrBYiFl0qb
+ar/TENfFc5R0PLLLmFr8GuX8u/W/HOjgrKg+qravAkycBU0MHqm1JNHHv7GvBV9
j6pZCBRC/lxj3w0RzSDStzBh5MTZNJMLLGqsdNQbTqg20HVI20TQTl92ev6MFYZq
H6l3qlgo3Le+7gz71i8QSSe1XKkQHiX1AYZDi+x1KQElyYVTacbd8MA7NnVsMden
ObpU1BqBrsksL7fxNNu3V8CR3o2sGVG8KhTHQ/wR8rQlXMaCNfq+Nmf65rjFCFiN
Bu001Ntzo/4OcZnXA5KovcPJxg3HLlF/2RdzTtujFwj1IriIAfuIVJRjamfUefAZ
od2c203fYmRmNNp20H23I5kE49r7DY6cuikoBdmvhQATeMiGp4DNSmZjQTrQ7SRj
MLZpK89qEkX9tKcMURSFY5MIb0FW66ToCVPSNwwTZfOMRg1ql1k+Dig2yRFmIwkS
C6YIzn41ZQjbSrfEeN8xNeKsB4/0SnGtS/ZXc4cmBqPXLRB+edMuJYqX9eJ2epjA
0rfeo7WAAA8BDbAAknkMO56pYqFm4qruytJ645QsRr3+h8dI8W1P7Gat5LqS5i/+
6rfvcmCTbKxyYl+Tof5DGAp2nGTRgo0/8gfKIF0HhKhGGtszV0TfJURV3ZmSs0VC
rFsdc+hpF6Hcyilr2d6eJcKX0SW6dSeqIfWh7xiDKYjetYH7jWOXcRgO6eRyNuAJ
IDCzEf/T1WBJ+oNeVeXDCUDQfU14MEqLsjs0bCE8Y52e8KVLWCQKWBDYiD/JiY18
THbqxhfBb8ecrwfgt4EaZ0jflpls5uug0TdCQyK4arTROA4YicRNvOPg4J0CD4YR
MnFOp3QxFgmMGxv5rVJrJlhQZMGubyGEZ88DxiOXgrzsjh/FZ4wN+SlIYwR6AtQj
y0gTmrifFceBwE9v3hb1JepagUYUtj68E+0HWYqOttrTpHZxWEPb34Yawz7q0udY
0NL8Y5f672LcTA17PBDpfUhQW4pKbQIkxXvcOCVQuFSe1/dfb0AVzP668GVe6Q08
5rP6SbrRKalUDqJkJwkivwp4y7Zx6r0/STNQVCct08oNr9D5TJYrnwS9yGCZdQgV
doQ2pvpBr8be9b6PRVJLdiIFxkXFDc1TjR8yBZBSRmGFn4afK/jgIJxLYSOZRP2g
SjyWElhK0Mq8Pa8ZuG5AnsFJ4ivsa4jf2TOV5iXi/BX/fSWDx31NFVHHoWBAS08v
hL7rqcR7E+WcMZ0VLrWN49ES1AT44aWHbjzbgsVz21wIcYU5W3sI5DfpcfSJo75P
eUihkaSop/2TLBVhpss0MkWgVq+juQq4/cXKgXNRW7cURWAoilew42fGZYvCqtqg
0OXZaacrqkIcJTMfhlA6JwLtoldS5zTqoidbhRfDnhouDqVOU3ZbOi9cXWACpFV8
0p6fHM3ivh4ycrvHoUMzCzsK0en119mE2VJR0qOWhFiqI5TAfwx8A0P1JHljJpF8
yZmHADdkvHR8FUdOng+V2FpnTHQ7crM8pgGAG4yI2HfITo6ZafUebbxm15DQAzM6
/6OmjAd/JFSW0DPcCFhPSdViw+tabVWpkFcLDnVxzcgedw/RGB369SkCBAG+WvB+
8GNWXmKuTXB/D0M1CIIsywc4e2sVsli+mNVwwkIs/OSFByhCUJoWg5IZfPQ2/TlS
6m2fx/TFFJ+ZkO7qiT1XJzXO5D1PJ0pTqvjlt6e43GX9HqrMiaBNxdbZRhs/9S2M
xWSHZuL4ft4w7gSL8py+s0+fQSKk/lqlIYSe+K3vnkYY3OyvN5UU/p295I6H07BE
z+vy+7ozKPtWhR8UnU5ibI28xQ51ML/u3X/M7DcDNjDRuixPKaajLoPF2apwLDuX
9x255cJXTsU2X3c+3gc2pHPqViPYLza+vPVrq7MEq5MkwzEgFJrMLn7qz+dAClcf
/0gNL7eWC30V3Wjw1LVsDnhjyvXmOL2y3fEWvUDEVBBXPSXUU0RARq/cadU7RVOT
csJ+UbuNWqFMmXAi91A4fzCy3yj1A9+dxfm1gmXPtMubife9ElUfRsnKPUwFwiNl
hFhUcQwdsxN8wEQdqvvEtDYZJCyntTMgNYBL3PIvMiNYm8eKooYNmNRl2WnBqNCr
AGYZdOdnalnUWQeHtT48lA1o0+2BP0Lao0nVHILlAenUvmas/9lW5lRJBUi0I9Tl
/3r8XJCHXa5LjNjEDNOPET4SzuX7ydmAh5bSz/SXuqLwEMjfQfWLNpXMOYeDFJ57
+DmuB/7VAyinyDBdHoaI0v2YfF1/ybk6i8ntXV4WeO43ysAAU4W1MH8ZQGwUT8Xv
X1BJFeABimfWxqup3F4oSxipPHQIF1XoOYkq/me0R0n0ngINVtwMYsIP6Gu2rrKQ
maXCzoOXqd0VVTcsLCH/oywkMCNGG7HOnugHSRZ6EYqIk9sMZf5dwsasHehR/w+j
tijo/LcjKguA1o0aAtmMG847x/YE+LaH6pF3LbF+ppdSouGsM6EgoXSNJyWlQTEE
0Jf16433tYV09P1tgTVFtoK7yBMpnaiC0Bpvj1QUDl/qVdwYVmWu+p/AYGEZDCFh
F56G50HCr4rCnaZV8PhIwC1XGIS8u2UGgg7PIdD1nNVSCulUejBa5VmL/p0TRdlA
NObKGMbV6/bZB30OslSXrC5RWjSJqk/r6B2UOcCF1x0/vhgAgopYsW++1p2tUe28
GMACYvrxyZmIwffTEO513mgjxVEnBZ2HusYAoDQ2LLI6toUxIDElEUGbljhNfi6C
eyVu2SLb7byvyP9IoUSFOOV/egzevoZJ7HkllXiwDqihZ1scITJCe5fwMPy8KZ2f
Vx7ajZrGJ5CvxZN3TiGX4UrU85Seo7ll3ICldYy7UykpQeaNN6n5xdZ9RPeCKycU
r5ZCspiYPiYTOMTg2iWIZICB+wMyJuOpqQVYNcYAdsxGy4hq4wrVh7YIuLmuly3n
Vy7fc0LB35MFMFU+b3WFNF8c4M+KoLB4ehp/Qp9nQKBjDwZ7lhA88Z82i2NuOHbu
uJIUGFdOtyWhX8QonJdLBgUaKZ4b5wwL13pwbzNadShOkOLfFl1AY3/lNYcTd0nV
D9Vx54EiEa4I6zmPxLdQouLdN1TXiK2wrLve2nfAqIKuDBvl6IF8c+m13+Cfj8rj
p+rRNXdqwW7E2kcuRkd0oK5j4wNZgKYlyPGsLfT+QwNdW1iup8PtIL8mZ0BMNfgS
rfibfkSZLS1mnDYpYAznWj3ijrfMKVDNo0Rn/EgBnh2PPO7GKE9dVhPWaN+wXFCp
qU/gnMRQH4ONAwqCwNrNsQJhTz+MPHlXqndANoJvSpKh7bNQvlVhYAyiNFS6Pa45
c8OfnoKfqE0PxkqBp0ya0QhGV+DWbntEpY3GOUdGErXMu3+4yv5V0Sqv7THA5mN6
fUL3D+iQOQou0XPO/a+fVUvyvCHFKEpkVJf8os2Y3aAy+AuNiPIa9rX1L9Hv7GA7
R7jUVyuBS9VtcRoYKMMsA48hF9cWydj5UGgd1VS4MTx+BZMMnn5jUp9oumzB6ial
NHUJ72B2Y41TztQxc1BjbnX9Nm9K12veLJb9GKgSnQH48Kkb2booAyJDYQTkzpas
zYYeAa27fZuqeh8+vmcx8/GiGkqsBQOQM/iMARmjCyXUCSU3m4eB/EbvlNJGKrv3
4IohpMTR+9T8KY6pGXEINDPSgxdsPtgJkPtUBl+Xs+Tq+QVBvkOI906a7csA2r+u
JxcfiYkBz/CzWAEUyefoeFVtUfAqmeWFF0Z16UMPMDte4NlzHmOczXnH85k4BaSL
Z0tVl0nUNOy2Auk9714Swj6V7x4h5bF8gJbpBHvUXCX0EGbVTJKgWkHaktHeFxnr
MwlmXT/nbT42KSchsYVB48gGEj7A4oydq3UavbX7qJgnls0NaM9IB5O2HZsKMTpB
+fc6/9RdrRzakPTAA8QKLVPJtOGneTk+U3jBu07t5T7u1vdXuPmVk2F8K9LmmfTr
n0JAZjOCIhwKkd8SDzkVpLCH5ojIdwIJQkEN/YUCtx5kqj/JapaA9sbcZJRbAQKI
Pj/enpgTlG/LcuVNpEFUrXYQAJCcMU1n6CuLArjALdkvmcBuvl43bS1hnrp1wc1p
jziOLlebJvdJd9cHNW2epAo+X653xu52xeQY2oxUDTXUtOCnQzZqz+ACZgPWSFP4
ec5QV8tgFaj41XopqUDmYHmAab1/pHaTqGm9CqB28V9BXDbJOZx+Q/1VUlS9SBKm
CgM6K7xJ4x2sLIpspc2ziCYs2LWWxFc7eiWEiazyr/kZSIQNa/lgOGeI3O9zmdx0
X98HJGKs6u9VLdpaqUBODixj6P70U2zP6j6jEKXWi3iQAb5EI3GELJQNjeuK17Xo
ppOIfIgPXgIdG54V416l7NvEX4dUr50S89t2zE9RvDs4+GTtkTSiqbE5fmN+20tT
1sFDX2OYSRiBFihI7oRhpycRFYsp7/8wshZBvyFDOv3njWqf8reaclf3hDfLfwj7
bAiSR80pyhUV+Uyc5RFawJdAwAVt+daCJt3dUvG6NoRvZ6ULCR5+X7fdkXLJfGWk
s5R/yqQa3aTMToYMAKAjFoFXvgdIqHkB2eKfW791l2bSiHCfjEir9EW5hFDrPj+C
hLgJDQggsg/ltwTfjZCwptSOQhyVQpLIaGU2og20T7b1g26g2Ps7pN++oadcNXRY
M5rh7v/7lspDUnAu8KvfpN3fOf75rUWCi6x7l6siEEzEmeODJ/Dynpl5J85JF65r
sSKHFVfxFC7S00xlcckiIuDBjKK5S2bAoRXsTD6XXUsl/iCqM6TEkiwJlP2H/v9e
vd4OIpHX7/zz9aqj+RYm2/3iCwE+TvjH0HqdSrvlSZx7ijpHJEBYCT/qqyDWrqcC
ZTSKO+1gYAPlN3WZvUK2g1Ykr6RblyVl9biLHcfXtkKA3MNAsopWIXxzP+StH8u1
AdoUHZjcKjp5hhOtXR3dw0wqcyVc+LF2cn97fR0BdX9pZJNsy+627dcUzGbGjGjc
QazzYxmH59XTRy0A8ilfzqPwSPY75Cs4joxl9ieNlyn6acbvybpP8nLZ1g2s8MS6
i9tmtSI6gikTeFTMbBI/6t+YoXTBayY6/4ucfaYTcjicvclndcnekgnY75PLMFGq
YrfOKbozB+4SEXleqLC2ArCQCQtn42WKiF/aqJIxCNYi1SU5BFL7tZFzUgpFD3jK
yhGBsAL2PdE8FSzdRPAKh9cHTvmUNAohQzr2ZKCrn8HlCdt64iki+zPZULE2K6Bi
cvWHXlUCHpwC1NiekcXtez1LocSEAGzKGk41j7dhslreTjcP/AFResajSiYpMiiK
zwh1N05S1Sfs1RBf55kPnJb5CFrHigf7Tt10K+UsT8xCydcorjEyg10akqhtGNm2
yO44/lu9yIbQZvXHd9Z942Fn1Oril3q2QPSiYHQERwGw++zOWTjk1u0bMYSoX1jf
w5QRTldZQ1yfHKhIxj9DeA85WqunxChYFrH5pLJfVMbb/vx/SR/quZbLVXxu/t7s
xRKerDY2lUwb/fT/N+Cjrpflr/bncHy35cEUW+/7B5o7meI+ej5HxiCFBhK/82R6
0U7Mg/V+XTYo+GVLK+DpTdnLTlxgk9EeDo2fxl6sPzCYwDOHdLPS4cS8paHRr+qZ
BkJoQjm84JVD0Bf37u3mI0OdGL1CW6swnQ9WQfRsqC+0Uu8YjIN2m+vDQT+KXc+y
huhbnDD4UEyZEyr4yZLTLeVieoCmPoj/qzERFsqLD3KR0hyLOWnv2vEqAtr+Nt5H
y3+pdfVaYiZw49xIBvsBtWjQsDWnk81bBSI1ULZ61qovbIply3FcDBaoYK2xR5ti
nqgPJ6BNW4o0nhric37UKHowZb6l+Z6IlTFfJ/vNvqfhx9rb4MfKH7lrfbvYp7Xy
2FfQ65lIeClQNTvg1TicABkHrfbGG1hGdYQfD28z+9kmVAwTlIUx8sMmPKAVkSYZ
NzlXQ5gD9OoWPpXCyYqRShpvJ+8x5xe3L8VV29mt03N5KJCWfiq8RQYa5OLh3/yY
kB7hq1J5aPk1g3G+cMpHoXfxyB1Ds4f+k8rLKlGzqLP4D1VqJzpHhUqmbJqprM4w
iI9P1/dxh5DsDbgVKInUUT+O/649vV1zbHd8yR0mF6jm8ljNMWiZZH6jb98N1dlU
fdhiNBG5aw9JPYJTq4TEVk3R9EStWnMp88wDjQEmbj3wo9kmWaC4g31pwW0I5n/J
94ozyy2/YmVTigpQScWye4SdhlYgRoO+qNB3sLM5VNUVZ8ns6Z2yyqRyqNG5Hx1d
+yppZ3Wq4jiLYjwQw35pejGGvU6n8ZzyMDVhVh6uikE2kfoh23FfNldo+81jb0UB
rUiNwI+GhEPaFMtAseGfUbrtoefuyq44+dhpArrIPOrhOKxuzcAJfPBe93hMWbB0
nqhisrRXbFbTBCG7XQ4/KUjsb5M567l4YRSsmWtaNQJJy4g0m2S1N58F2sjJfGNp
+FR6mKHkhN4atlH/k6twXon069tMxHYAbEUrLK/Tf72ZoAb/6ntx2sS/team1VE8
8eNZvOZkJIpPP2v+gcyKT53x3U/kst799ME6zxXgRWxYgFwScW7+YOOIiZnocXYG
wkddNFIbTUf+WWcCfBLRP2pee5PeJ/P7nk9ik9+u0FItfKBaMGD1lGTY5bc8CLM1
pr/SV+dI7P/xlYIrfhiW3AyJ7ia10+29QoJmCiDs5I4B+aDk/ODwPtVUUHN9pH0b
LRF6i2hcFz8b0dG7DTFaOyvF5waqope7k5apH+AxtQ/ftXNscW1+1w/tkJW8hBkm
TOqIJ65ZC0oZf0a8/UWDtldhODEaHUrkXNYDk3C/JEPOPNQsX1k0nR45ppKRLxc+
mQvq44UBl3oJ6zcuyoLHckSD53QLhJGLg0pmAiDkNFxjpK5PGRdKIV7++YWiztQ0
mth17HZ6XNiuKvSVI2jStl3TValQ6hqHSZBvh2Tnkeb7M+xx1YtDQJNgjDzYiX5j
NqAQsyoCnO62amVBTsHnv2E35nO6VVCi/Y6P9S3XWyfe+PJfYnk0hYogrWgolG5R
vYNgFW4+CEBPCZsUq0N+fqGZkAgPXe7dFYHcVoSFRleM19kHsvmie8aMsWdOA9ux
7UJ3mdGkIDuR37gK4vU67njxoaAfzp43l1sj9sKlGSJoWwytOtZEtwslt+Z4L5tJ
bgHZG7v/D5fJV5TKrRUQtowOJ3xTj/rK9pyOR67433aFpc02hd3ayV/9YNExkQx7
gpcamKHbWMzaW3irv97kYs04ZuNE87/YTRHSYEsNNR/QDV8gzRjCFompxZYzlMkA
1Fsd9KXJlzl80FyKGSbIWsdYzMNr+9QlKDDDyHQ2lqsvAWuGymHQWk4tQCfnBneQ
EOsgzQx0q1pyjs44eM3G2E5eaKHWeV6UB2GdQGTOvIAsd9P7DroDuXjtUU1iVDdp
CQeVacY+FNViP2KvERf/JSMymjAyUr8i6o60pyzYO6Z8gK5+AZK/jewM/DoXr2Ea
s4U4pagpYQfYhjjLaH5JP5GeutsfTCAeC4QdqWNyt7hQihKnyDa/V3J3kGQiPUtL
PA1mux3sPcW6SBUaknhE3mkEc6JvAv4UekfGqNz4mM/L8uAyKCa7IaGRdKcpze4/
B0/yHKVtH4yX3mcntzfA1MU38ez4oWcsIV+3RUkgwrOxaSti/9fRoENO+9ahn0pT
hQRk8NcOKt2ILSTIIzy1f8LZgn+dE0XqMikc5tqMcgT+OS+eovHeuWgiIkw3nGJZ
0A3Yl9GrXcK9EC8Yu615Lk8W+xE6GDx+RftINzR9zwEUmtGvn+Q3c/husBWROdR+
BhaiHzhWLnUmVpupATur4FJ3JcsxFFcqupYtbs96FcKvCw2bK7ZvRZuTqLQR2IZq
/9hQVnWKP61K2mhpIvUlkncrJUoYSdgip3nyg/qT5ySsIB6UxBE6CR/mVYxv7E2U
TZzuNrPjHriSU1gbLtldaBND0OdfugwDtKraQp4b0a5x9obZoWAGrkib+vD5hfka
7oFiLR5Ni38mTtvBTNj7LIbNrS8MgTJRpV0OeqcFHIhkbYRdPQfTh8vUcRYSIaoQ
o8lmF3WzwDnYPrclK32Au7AQJW3v1lZqZS2hiQZy+sfnbyRXcgK/V5poCPfu8B8N
sZSlOlcgZymx4d37rh1gtqgiSfDQVtTIfFN9/1Gv/1XkYvAkS+aKfNdix0SUvcp9
VzbYmgdHTbk5eE2rzf7uQxRhu8SP4lVycQbR5Ao6cS4j3YgyM/one4GEzlrD0Tq0
m9xjTRys1j6N3BKqjW5K1uwCqoh1PkjohQN9yxmvD5So8Cfb07v+Fu/mMazpzOMU
9cWVKtdBOClqbF0lMuWj1AnsEr3FJxRSksJHnLDAJINtZlSbHnnNlBg5ARBzGvbF
TGiZfAJ94koV/9cxyO25R5yEemiMzbtePiaedGGbkwkkxIUHG0ikQMrvOA9Zn4be
P+RS0gAfIJ8i/JEFz35/anIxbvG13CFxgDHiKhnNme2+BLIMK2CHthCfUwteTYXR
j0uUQkYMkzuBtQ7HMrOCY4xYeguIEJ5o2i/q/nuMfgytlnlVTi8/ya51OfFArg+Z
57PSJHBbQwc7fkfk2GS37M4S7xjTY3KCnndZw//YiOhEm/BpZ1N4TjlhoqV5+avc
yFONMmMlh3ZwFPS8ltA6Wz4nKV/C1kCY6DZQnxuArpAptKPVeL+WvPOIUyrAduSR
XW5J3GV+wK7q+X0650GdO1PvfNO0t23OcbuKSGB1MlynpPVNysMEramuz73F6SvB
79FH1KNqggPzuspAUJ/V1y/WJj843a3bFtm/U7LI3+LzOHGcT0X6c66Zfd5IX8YS
pbdhhAvgeoGPs8J41L3Bmjux+HIus99DP+zT7XFrBuOxbQWF1fdIgieo1QEIAqzv
53XBV7ckNYIDKVSolza2Eq4pKGw63qOtc1s/x5wRjdKToWlYS5StdT9mfUt1+ejQ
aqcQkeH7a2PCRqrsBMdJTOmZeGtqIScdj/3wEag2+LcKontpeWbo2QKd3Fftj9Nt
96yNh2nzl4NcLl0jgbQvgHFM/NvfTw9xUQ9V5Ny7ZFNpLCkfSIqH/E3U6PEiJv0m
r4q2lElh+dAOq42KcsRiMrLEUmpDNBk2vlYc37hWL+8eYevNH20KO6VXShYbA0vm
kAqrYJYqotGvOvT0t+4pQ82tDwQROnQq6VJVZFzb2hN2lHxbr86JerAfqXxqURT2
DgwW1uHCTFGW60CdMSQGhTl+btKqdnh/QkgtQa3pNg12BvS6oqfAvcbtlhiwrYa+
A3BdZCUovKGGDtLJeOnTtz2Ihm9wvlXmKuLBrwuyVw3Ssa+iwOzHT/R6E3nx5nLA
0be1adt3h11/O6iuuFgkei9BA7B+JvViylBdG3MoZZA3sS/z2RhBbLWlz/AIkNFb
XOrwuKfNNgIu6iVDVHi+uK/C1mx7vHE8CEqsIJB/ovyTgaydQK3p2f2fIvykatNd
BRwvWMlVwWG/HiAFyiiMPOV3gqQT91raNPXt9yI4S4q5tpT64aLh4vknl3/Tchq7
VeFlJzCbYs2luG1fGDAnKYW2ZHxfF2qyJxrmxFRt97CVtoMAJ4xth9HoTBAfBDdZ
aDnjVBv4rQzJD3jBaC/KxKVu5yVQiGayMNWbA/wHXQIL7C5LiacqMtBIWN1cihuI
VA3NjXWmYLuusc8vLeWr+QZmmHmL3nO5sbH0Ap2EW5JCg7abtnATW+KjEtPmBEji
/6rwVitbFIM+io431HD8+sM4APhBtSQzn92/ej7ABE1xXqdNDIeDug16gxhUyoW6
pfmeZ5uuPiZh1rnlVg5Cibrx8xRKMDHA4xShx83qbTMszpr6TcmT52v+TEkOwXfO
cC1MWGAR0mhyowbVTPTHQu5tJh3NeXwnvRI7kmmtwsFHrdfI95P54UryoMPCXM+h
jH/pIEbDIh+mtnb0SQRsBZPp2RbvA4bQ+YcWfI8/ScDwfmhGbd5aLadoYCaew+6x
GRNMOSupInl3Slv/l1vjFxHOkvmwSd3PSFNYQxL0mpJRtS9luDL1pWszMsMRv3Po
tTOZskXbvbyLNvUiIOK1KBmk/aNWEYOtWw0D3uHXZueUBOlOp0vgTbhMs64T73hM
4qLivhpZHkOrz68lXyGKL/wDahrxF96PCxMduS6hpOMuRheUEjOF9RCe1FUEsOGp
BFREO6i6CpaswUpSgKeX9I22guwX5BLuWV+vAMyWSU5fJPkGBTE/6teU7yuaZ8i5
mSHE6PDMSMpcbjxOh/m0WXGP840mdJkGAuJQqywvRwr1OEplsRmgxvyr2yMjIDhs
Cgecf1A2IIkTLBGw+HdFDpHqzqlnFBF+VvwKKV36Kqa5a98FeB/MxHDzN0MX0Tgh
/mx9dIHrmnpkVsr6LU3qHh6Xq/r291PtirbZyATvl/lQqMTrhXYDP2GHYU7RqJxx
OkEDjvXojge5W/2xkgycsp84vS77FreWgXaXc8Id7KNge/9xXNRDkCsTI77zaxAD
4hfnsIYJWPIFYCTEtuxSYQUGWZIKNwHtuFvCqY7BjPSmRSb2iJvjp/Bzv6sZBbRF
+0axAkxO/U1haUuzOgtPIbuuQOWeE/mb7ijXKx18T4cVn1yqCxl+HMFPfVsgEhXj
ZW18TUPdfYh+H/ZM/Cjdb73kX7wCnrFKLgT7LXMPNHo6Jj2N6fbUZx90ehgXPrSC
xzUrgLkKXkoTofqKCSkEUgGH+CJGtxVT9Gi/CAd6OmmeZhYZ9pDVhTFlyLgJyyym
7I7Xx0nSHXoEPCC6LZRfO4CJK8L54Qw+uX0//k9yUJIuRrlH5W+QWhbSyuao9s8B
AfRtoEq7N7gCQgkzrhc7O9zA48oP9aYrARbT0kbLSmnFwN2+GOMQAeRgfxZBcE5H
qBOY0CzL+ttaW8fQcnx74lczDhP40ZFtto8RmyXgvheejccbX/Ed0U8zq6zjYkLn
/ZFlTshHQFJVGNq6THeF1s6yreEuhNs8AJn+hTXR55A5Q3PFZtOHGEdTFhSH8Eh9
65ZWeVFOUJDA4LfFlnTFiRDfbMxbOWCeQYqpPO2dpkLOO7kFk4a4DTtpAPbq28Pr
r+gSY9LKzvV4z5VjDgQ/1a2WSG089A/lvV4LVSlVDFXOE1CypQdUvocL7gXinJBl
RR9bvMda2eEukpmTsvV5y5/kB/vRPoaOY1DFcpjSD2YEJ+gZOo2yC9kB9Po+TM4z
n1f1HEoNWNiEXZS8u2PNPzp+ALACB6kLtYZ2+seg8hoI/PtqcfH5hG8jI36NQRsT
46DZm2NK6p3bDy03ogn/0+VSMCayxMlSmskb8YWhlv4DIMigS1sNZHT6T7pPDadx
ki6Vk4HBpVi4d2FBt0gWhliGZMgkyl50ibdkGMA9Pp/LPGKyuafcHqFp/0xZEuEO
UKTpPqymYDPI5/2BbLGHOi3wFacHKNTD1QvpVbWLfCUMJ1p9zka4hERClWZcKcLz
h8bpB7gpsbLgOf1rM8GhamlOC5/nEgQq6ooszC5YUKagQ1lptBMeVooF37vQL4CE
tnp/PLh2U1VMOsvzr71cs+H1U5LDkNKpV57V9HhlGAiiVm49gudzbciIlYnlOa20
Wr6iip0UP6MG46g9AKSegPdPxe4TXwpR1YJHEBPjKlO5WFAPzABuOJ9jGUobx2/f
PNJA1uq3CsEtaooToXNOqjNZbATB3ii/M/04u+RYiPOng7iuin0tZDSK8RhQCnoZ
pI8OjpuwYynouzkJxOwcHtE2fH+VbwEeXqdEcNKmntBTc+k9ECamYN4Cq5e56E3a
UCFc2ecCCzv9V1n6qUMIRCEats5swpireVkRkn4Huj50t6omO7y3htC4JC0JqlCf
Cl3aoXSIMdTXRgCDchJeu2PCjuw1K4Y6tUAlqlX//qRQa96DBFjgTRs3r5PsW8F2
Wru0SzWl06i70gxyM5cLorlJM93mHpglZ3cnE4ez44nWG6R+n4F/BnuRhp6F5IFS
/LM3SE10Iagkj7tr2rMK66Qs7wyQ5AZbK1L3VskcqBNBOYofI3OqVn51HBle6Dn4
SBpHaVe/XxSo2DtfJttUmUmM9P4ZgXywkVvY0AG2c4cu3sA9yZPAehKoDQorXSN1
njLLWbCLihK2Qnk/4WOIn8bWScNyJ1gbVOuTAVCZvP4crLwP2EUgGXizUYCQsTPv
L7UkCM1hIyZOMdyvE0/xkTcbGJzpInfAeUB1AKp1rxoJUkkTAfTLZG2kPEPszZ9b
o6sxyzf2TP83lv05IsiGmanPEkvtgsTvsmhcYB4b0sZx6kXHz39Mk+HzjAQM+J0h
VuzEKQbVfRx4QrwN4/8dNhWkDHV6sxFsB2j/L6yhh8OhKpkLrp2hMuLzHrmfnhJD
EmY/ea6qQ3E96Q/7uQvSrf+V21+GHHWL6Cg2QCpi+QKy6pa6T6xaIwSQiPwAlFm3
bNYDfM+XWS6jy94WV0FgsXDgPIVCnAfzA0lvojqoNaRasZgZmOu/GOqOpRmzsHXR
BOThrynRRL9XupuXKRpqip+RgTtxvch6Usqw+TFtKRn4s7s6kM46dvsqnfcI8L5v
NwSQxZDRqXBlvxblH8DxFt8Ar7utqMHa7o9J80oR4KCf29q2eCKCtWnGTrqvyEDL
teGD9ZCWme+xt4LcuJruEUdx31YnE+tvIbzYPiDBTbacxGVUVX9wTFaIB3xRzlwj
pZn41Lbt7rrxTOcbKyPREpyReN7hFyOE/1lE724YrJ3wpS1b3l7c59GJ5bxI7iFC
3RKt06PE9Zc7CLVb5j84P/8BDGqWo/yRuVcE5Y3zTHIG68I78UHvFjz1iB9zVeA8
UVTbLL2noyntC6N4krcaaAmIn8knXk0raGP6EyMhakZ5+VwNfgy2xnl0w7AFgUn1
2SQm0L/j5YSNUOWoVR2OgJcutBa3ePkkD9fDdB7A9klV5ckSyEKHZWdxOM+S0wSk
B9q9VFc374pioc7LEctKUlCMcRS/zd3COsMW0WatxlJGcQL2PfPS+MtOpjjqGnol
pGVel++qSrC9JIRhVHV1muLjYIwfBk/dHGZcOYc98PLR9W+fDXsOVOic25OdW7IO
haDB0at/e5pgLat6d0Rlc5v8c7dz1LISrhykeX7u9hql+IWSM1rrvVedzi0DL00L
xYiuIir3SA/+6LuboamiXVQ2T8tgJ1B+ovV+GgbsgrBh0KTPlK084NWfhhe15/G1
rCvivF2pXJq1qe4CRgVcT6J1IGTiwuxAJMdx3EpYuej7pnNQvdNh+X5kiME4i5/Q
P/Jn0oniFjZnGsae+Kh8PAM5PU7JeYk4/x00n6606r7Seqi5cuUpaBjwqskhgvLD
uujyvR9jPujQyzF4H2DPu+txRPtgVBbTXnpw7hNw3/x1rwA5sOgK5Q7LbeGDmAjK
mIKdBBIOEkQBL1HjbonUZ2YNIVd2FWzIGgwuyYLVTWY56h/D3E8UXpB2BqKDuvYZ
TACYJGdaxe7ZAx28WtYolfyN4jwOXBqIlkuWYWv+uyXr9IFwU+fwrEdSWaYL1gGH
pcVYQ+hlxCqiS+iYl2matBm3S93WVx0PmDyo+OlPqi1/QQIAZv39b+WRn3S/DRl7
xlhgpqMN1Ryw0iHQ5gJDVIQcO+KwL8K5i8cz0MPYpdDsAFV6qRPqgSWOHauABztB
TVXgGAeMDcU/xgEdUNs8Rdznk8CFyJM5+WV7xY7ytX24vXrQCik+DiXCGAGdgY1y
93JOrB+xLiqmrFL/CWnROGjfJfPShvMiwMy0NUTdTbW/UGliHvXCJYRA5WX8zloY
0hU/v2LD3Qa4nRDB/df5aoEZdX/HxxDmlwLebImpDGesAVDNB4hngl0IHW34QGKr
Pwa4lFKJOdk3RKeocohBOc0KVwCtyI/ppzcMO73OItaIt9yeMr0iZqfX36qMK6Km
Tmu4CbliV4A0RFrBBFF7PAq/UP7DxtUR8izrW9ef8g14+XGJtwCnTQ9jwvmQD2b5
+XxalrOKrVugLVtsgYb+zITf0UQqm1CSRGbT9eF9z7pa3037hBzHxFW9IlV2a67D
FFOJZivJTvM+1AvSWg1vNvy62p7u4hVD4Aeh+0KgoCmB6PB/BBmiHpGil79MuiK9
ZmmqiZeOeuow5R3awOSGbB3mGOMICw9C7PEPYGZOuC50gskIT5yR5N6zem55Euau
X4FVdTXlVQ/Zrws+Sql/YumyXKDNzW80yInz3wAevEvq78T8JpncMrvy5DRFfV1I
l7EPc0J4dW0ZKjrtMEN1Uj8gfiCED9JOniGY1oWLGDDNMdcZsGeUtqP7EnBHKm20
QiQ7rvM+8CqJhI4W0vthKOr7E7ypnPIsW/hpqYnZiWWOdUG7Dg2F6wqGbX0ki2jG
S2A2Nj1Db8E/EXY7G2HvEUIYyeLGRk2D+bk1U3lhgeAT1kfFe7CKviE0aasvemu0
zUmLAYSkZZ8uUt/3JvDCt0tkKQecEms0BjkVcDHmvtl6fMQ6oH4002sW1RTsN1vi
3HlYttaWSMFqozCrPVM25/gioyp3YHMHV6tEWhwJ60/Pr/OsNB7M3ax5pXeKshai
6dalohZRfO36C8381mGMiF7Tw7naHQ7Z04S7rpFjXeXLOISacdgS4bv8rLYwRnU9
AqRpX1uVTej1idqkB141EUcPlEGga8FVx2E5uQE1XkDeymDb33nXg2QHF8qKcxnv
/3IxW2I6/9sPZkUjcqIq+zOP/wRwejtuJRCzS2E3W/u6GWcjWXrpSbuS/svfH44K
gDT5G0wT8ZjdQkgSJbBXdjBwHAiKDtPgjYqxEYP5sN/E1uTal/MOeHRnaOl667g2
Hh4zLucF2dAJN5ddC2iYpGUFMV0GwCWFtj6z2MV5DLInH4uUiPsCq7DJpYM7bL5d
KbjSqi01UGRLb+AjDdende+ipT+AKL5khhiv7cvmGkwUgyQQM9hyCT6+bKEcIKqP
LiGJhI0wRbsY2OgvcqubCIXdypaGi1oUXN+MHqnFvnEnziP5xG+uemLlmgNQOYO2
FQALzi6NnDeaamklIfh+gcXX2KnNOqtb7k+xfGhL/eT5hqFrnJa3rf6bEwMS2++e
N59j0jMUApGtTb6my+bioEuEnx1bfa8GbUqXulyi/H0FxKLbzt6U2GPOsLop8SOp
sTrVO4jEBOA8dOm/Kvj6VkbloELnkSJ0WDnwO2RVwRepuTciJMoC/zNmEfREQsei
yzFyE4cYQYW2ovMZZZOMYG0VwLI91vyuhUVbWZGK1B9cPGmdtxZl5UCIEZe4LDNm
jCk2OuvJLIw0RWPIYgF/sb5uziWVS9s9N0pEsDf0LXWqd8tj0V8gb+XO0Myrs5Vj
JD/FUBtpwcT7DeUvvbQfugneJ+NubjxEFrPp6p4Zd+cKVq8BNAGpbcoswl4/xlER
VyYJS+7ZtvO/1u0Wcza8X355HyCbD2ERqOokxnoY1dMaK+TbhujYYwwzLzS3FKEg
vHPnj7lGj/epxHTnjodogpu7qWqBY1xzr7bw+rFpGjqXo8ITwjlsrnBmDyU9YfSN
SJ3XWSWvqfbty+Ns6XFJuSVHn8JuQZbT0jYVoyic0ggZiwSXMA4hXodaX4PtpbHa
2msqZMP8kqJikyavngqhmEXJFgbmCUvXlyd+reP1bzZLnM0Ejs7WJIYZO2uZLDwu
VLatm8asEE5RLvEVww1a6E9D4K0BRKPdL+Yv1p0QYieCpyfcQu2hq1Fusu+rJOQC
u6e52JaV/tL5t8jRHmqmmxmwPiPUKQEvbs7rLH5OlMU5Fx8AOqCt4WAm0q7rCSD1
QThUkBbZNa+DiQjEYwVbxu6SAc+UGRpl3KwDYqd8TI0pnWWFtS4qJu0DU8WEREqH
EXWpyQ323urvzTT5x8+p63EIZu90DCckjPz2I8rC5z2hnP4kVe/znH4fpZ01yBT8
B2DwHV5xysMgk9YnBdrrcCnJt7QJC9GFTRGO/ieTiy3I3a2VwrLQwR0KFioQWK81
DUzZeQ7x8IgHAjsDUXjvH6CcNHCzq0mgf8Dp+E1QShvk5f9645JCHTdPT/JVDtpt
H1ND4KBuqfja1OBrwu0EQ8GsOF/NSUMAnZZcjBVToQOmSwYQ95MjiC9NxGA/AwVs
PGH12M08gvFWZcEM5EQNEVB01SL0ZEM3pGlb+39nttpyiqt0RIhl3V91mcBUuMNl
gK6Pge1wk6bxRKVFJDgTIvKZn44ERziaBHr6uuJ9gS6FDYowQBfXvJgfUq+nyqIT
fiuowzh3Hi9Qd+rty5tu7MB2k+H9iZ1ZWOo4JYLJs6+it1RGc4QE/DW8AoOzlVbW
sW+g6H2TdvmQHgFRa5GO+A9lihm8lDe1kR+TxmWFHlaQBIZRsL/EZGvLk9Nv9VxZ
HeXFRK5Pg7pyeqLsgGkuSjmrOfZQonGDMqBjaiBNWud+4jzLlezSe2SDo4pYQOg7
wpjctnQzFTUVTgIeggNTJl2fdWBN+jyzG6Yp38/N800UaeuG/1+j78l1hiJ9+R53
ndAOT1XpLLBx0tNpJwqnM6/VFnSwhp6ftRPm9RM3579/AqLl2HDdof2JsVzL5Qld
xBpvIvqndGe1SK+Paq8zNYXqhqwF8x/sdc4ZWxsTnVrbMuIXUkqIs8BdIN635HhF
t7mVnbNZhZ7IgUB4TbQsiCyeouidqErZL8s0IJTwhjl6Mexh1Qz1gdmCUD4Mz9HR
PlGMce18b2uKt1lRWfP/1uUCmKKF0X0l2VLCNnbsWewDeD3n9tN0e4uTtf2vyBTz
lxLhtYhjgtl4DkKcu9IrZ3b0rxAQKbHi5HEH+0qO3heEwKwyuVJsVo/9C5sZM6iB
kbkp6FvZQrkDc9t1O+pfLJY4CgQUr7J4gwhAQUBDV+VjtxL+ssmQfpNyxHCBxdDs
JHid0wHMH74IgjyHtQNp4bkto5/f9P+DLUU0jS6Fdjwo5Lwzy3sNYW2Ma5MtVYqD
OUCMLvAOsYllWOiOefIvX0qsWJJKUNurV23yD0dLkWFikBqfMDiDMGHzDU/XLMJ3
7hLdxpfDEel4Lt9bCQktbUvbsfzdLIqHngp64AZ9ZpkNj54vyz8Fdsybglprd2Pt
Y0H37rWwrxanWUe0cpZhO0b+qy2EbBenYp1RIYXeyszf61lV7X+DOiFJ0VZ/HTec
tIXhvk3D16FjUiAiFeephrLYfb/fsJuXH7TCRXUW3JSOxcmzwNUJJcQ1/sSGp/A2
dt9TpkGiBtCG+OKDP41k2N4axGkRfoTjhMizrt52gbiqsfsUi/CppCTN9aXdsSHa
/67m7TzCNAy0QE4D2lxaNS5+9iRcqxooPWAomtfjcI5jkUBXsf066jJBsrO/ym1w
uY7S6HAlvtrlt0W+a6tmFJoLixB6betEGLWCbA3TUx5SGwB4i90AfgeJaY53N5Qn
457O08I/qg2BYHaGrfFH1KTj8WfmcPTtYyskyFruEjYNwc/fu1Sbe8ifsgVuN/Jj
C3fLKkdrq7JN1+hmBGAPwjuk5ncUtr1z2julWHlQq0xGiPBsWhaeS0SIzKaHONCw
EYH1U7VmdsDOtgl7da+nZkjV1vKbF68k4xzfY4tFNKkeNRBPZNHfd4qsgwkhI0jb
oflK0hM38YT6I1Anr2cwIZx3om9atzwgcY13sdBTI3Shh9pedbFu7BQ/4Xsd2YKj
hUA+oiaUmviD8CHXsl+CDAK2YIzYa61TEFOMMxOKejNq9NugENGAlrzWVmG40O4/
0oYQH/r8UhOxs3FXUfSa8aaY0TJ714sGA4ICPtkRQPdN+T/D0wN/zCGsMCN+nyNR
n5YRaY4qOwRu0F24BW9qj3CT+0qpcgIwV83htYPwBvVbObivKWhcE30+VX6NsXdK
nREpyywCvc0ijhjsgRf81H971sYvoWHpynDJ0JTmeek/hhc1zZQ2xC2C2TpwzOAc
3PzA+F2e5v5gmieSgyk2zQ2omPvrc57ET/bXxEesg9iU2t4xidmcaHCobH/EDXaW
qvjwRehla8Dhg34hCuIfVnSMpZ9XVSjVFz8Q8oRcvhnHQhZlaWsflxUE2zwg+bj2
4SuBClJ4J+qhY+5MH8VMPV6AV1Ls4oE6LcFxuEQVYSywj6zOVPfXxcnCbv1+0/H3
ZGy/Mipk8VeVqIg19Fu6iIQ6gY33b2kbZOPzEgKSNSpNVfATKzu8RxepnnG7j3ff
8v2AObbawXAmM45rKwR4oBAGMZZ7J2IXlW+cGvRDWIabkcpovvCcYECAD1mf2P4B
uhkZ0GSZvlY+agF96YA2XFqjCkh3psdqzXmqYOIHJTTINommXzslFpHixu0r9O1G
RF7fC1twCDjI/DmVlQJnzBbRce3hyhVl0I6Wz/8DeqoWhqDmQmKmVPt/msGwhIOA
rCICwxoQ5LtbA/fBjnjfAgqeXwDcrYg+DYZkgFQGCOH3CQuOti60DoAmeleX0tuN
0/2pkT8eOFs5LQM3ufSzcZ6YwUCF32pgMzOjzffCTnw7vDw7L+U+2NKHWgPuREc1
T5i6iUY6Tx8pu2X0kjDuJlb2m/RSfNbrDb5A0uLYwrH2oQSH6Ze+22OL/AYm9inV
VM9nFpRt8iSptD9wPIAIHLvhndzZknUTYlb+bQQSftIWL6zrzdX1kOaucsUopWos
IPH5s36Se+EPj3mQ44OaxSHBHnDU0au7O4cSMHhmhYCT0JpEbjzTSVskE2wRqrdb
zC1FnbEZuOyHO0k+ZPi+0sZrQ9SAodGLtFj9dqN1kzi5ElX9ek/O95yo7oGMN9QP
tP0eh7J7HP/JepfMJN3CJG1pNtrYzGcXj3b4tc5iD3nTq9jt20O//0wyzRoKk/HT
jHAeTPNqwR/WpLHBsXvwsfAluN4aYa6bQRlCO67tU7a0Tln+7yGIkZrpCGBC8u9w
vVyM2WIg3NN4swsMh7ZDaC22d5i42LjCSJJZ6YpKF+44KBLd5avBePOfT9R2oHCv
Eb2Q/Iu7svmafLSVse8CMJlTqEqx5ott0Tvii7AeYsUUhb2H0QMvfq+Sm6mvCv1S
Kno6xlCAJPnV95FykO+HAOiH48n64/SbcxXLZsA5OSflSe0uJXEQR+sToB1x3dcq
kbCBM8Fdeuzi279NFUP1g0cF58rLxRXWQczq6mhlQVq7PyG41ZUMeAmFkpeE/6BZ
838aKEZF5YOW9jUUlMGz0dHOOtrP+QNXsQOfs7KJD4pQqKhl6DWiXMzw17semr2b
ZSfgXjc4YDCqJUehmafa9uqAzjY0atlXd/xaL25Lyb2BV64VSbOfgjfaKLYuBlG7
IHiRPkymNZVJDmrluhU9TBYsgIhMq35YIzN0MIwFWWNvLhbXwdbIYzQSX5Oy3anq
jeNqYHqX85VSgzJLRF5iukRKIU0hNFbVxlL9p2uNtQdaTux8QYRZRho4HcYj1vWZ
JBOTrDCRMuOgNjTZlmdqD4u0qTLIaQktGv1aw3Zv8/6BPbxBo5swnpZFIM6Ty9BN
04833UoLYIqAaGGKBW2fnsJF28IIDAGwNBDPkfuk3MglSpkc0pnVmV9SYpagXjG0
dDrOhzZUQN5cZk5AW+RCutrthgrO/k9c47PvPh5/ggCyEhTPabjcG5R2Vkb6DjgS
dZDs6vPuFM4MZGDIkSV2Df2pt+gZpqXn1e7Htd8ZA05xCsVwe2V1DcI6BZFYbXp3
mkXMounu9afZkuaWTB6SLOBpdwvlT9L9ml3pyDSyjT6ayN4HJf7cYeLEJs5tvDX8
LgKJqpHMjDwNSmISEFvFs8+0MhxS8a7C06SQnwZQ+cJ8VJGTMMvdfa+aGyp3P7uD
zNOee4bQQ04X1ZGEoki//7ALhy/FhDWtPZEru84jpmlgV4JeHL+UdF8z/ANtDhsz
fBjSuCkJJ1fxnesTcIyEzvKwgIDFw5VTSYDzp88SOlcx6cgBhecchrWJ7lvltZC/
hOs3qA3mDgDv6lUpsDVx+/kPM06gf23etoTbPee7obzx39UqUZMBPDM6OCc1+9X6
4Lshti9XbXRr7+HBhrG7wMjZrmKU2ROO3PFTew0sCOvRguNK/M7jtjXZ8c3PCT3j
oMTE0sTJXkl+hrtPrF84ZhxEroyJwSLU16VJLEqEPSigWICM+YI1eg86W3HZKua5
o1Zs5cgNH9qxya5o5etPVdQQ778olDQef3/52hRDZAO63/kucwBBi8QIX9dSyhqZ
ypUtW7EJTY5hGXcmaHOjnhI536QuCCikEwBCwFx4O0Ubkey//3SbV7fDFF7hB3kT
8BIRcJsgxQd2PtcaqFIShefJN6vpfm+8fcMhPPuMBEZ2mCaHvaf4uRKUFOaTngjl
ah3ujtDvlpCQKONzJYwMFPWOh3MlbRU8ESmDDCGiF0hueyq9HrxRlOAOkXjR0zxo
eOn0Jn4p8EsfL6TybtvvVptXmuHFv9zR4zqW6DIJA2laeemh6yltVPVy0BQXLluB
46q4cW5u5PvgK6uILXKkln62Rm2m2DYpj6U9FOj5r240pRrqiRQg/47ks/MA9n9z
pW++XGAEtjfnyVXI0SHWnoK9rCvMq1ZSszYeNfrao6Mb7jLsqlLiMcLT9qDgWE6W
KCuTG+zGPm87tFKEI7N8+YvirhsLDQ4fjMEWI8pCnq/9yXjo+kTeLJHjzuJxBLwm
wmJcIRNlrQMVHvzMvBT2OQqwhGsoAVzuMFwb+9pmoCnnkYMVz3VvNvObC4DbD5FY
hHkz79TNxMtkdoMnKdNmfIwGgQA0C+WOPYPXILui+HwYqtqRPELvlUMLtLdEpJbv
ESOGfpK2c7zcs1i3a75xuR0pkW+FPKEHxMWzxZlF2eFX1eR1LkrsyW7wYBD5PY6A
u7frXEedU7C9L/GzzAoznA+CEa3pFhvMKRmQAxtoEZ9kO8O6L2aVJW18V9gJ0QQ9
pGrUhNZLqPkMxagprw0VK1/9+ESPrXrBwmKbYQZDGnMvHMakFVUP2GY6VH7RjK8D
OINbxG//214fAHOx5b3O1CucVC5imrpgskDaZpmn6gvrFsPiqiE0W+p0ov/s3a6x
BKSt4dNQlo5ME/vlxkQs1YWUher9SennCvoGc1VQcxKiX7hMqHmDPKpkrsadhiVf
cx+HLPQDvcl6jBJhb47+no4anqKSoZaKuQEa4k6FZyFrDhGxXcOYf6WTJAMcmFij
PL9WtPxhNvAczp2uTsuo54wbRVzVYfCcWuR6vyTEQ2a5jGFjEYKHKDm+cgOIBbPv
6Fh323iBRH0ml1hRiSpJD1tqMB25HEMajxnuuR8dUB3vzalMh70wy9mhB5+ItwBl
eVyu9nySZT0FOeW0RsGRv7BxoY8FuU/zMsZ8D52efTmz7dW7mS7uAQkoKkEK/H0y
XEKCllaneLcgCR7P90PMRTe8K6/kHVZafK4MXmlXEzhNZPoG7y6RpyupPpDoXiu+
ZsLF2J+bmNJXaTjr8zFP9yCy6wL/3JUvc4N3K71apkFFcj104sR65wGaJL1WXjgu
J6SdMZ9qvriyARqgizMUHWI7FdZDrUvbeQJwQl/NnBCfquDr/ioKZHF/fEegRUDx
0dnEgvjSchBtkrU7/t7q7bffzh2LLdQlLF8LrIOcrh+3Iyn1IdoQh2ovIr5q8HWu
r9kHQ4iM4vWVI8wMwNe4TzG2uexRnz+xpOPpUFw0wyj9mAQFtj8LUpSrkVutVpAr
98hGf5fFTrFFSSvl9DO/PoxvngmptFd3m2EOxAc2wkaeEP5tp71PIJbXC1+TFnZX
f7BjCZ5pqgHFNgF1qMLH9I9S/bDkMB9NfodrBq3MCtm39MI6Xlo/Tje+uZyhe9rY
uXpa0d/tq9i3ShBvxKk716qJ8W83wdOFczbuu/HlOyO5/kJiLSnE2GB7AGJe3JMH
53ssyRCP7yQ8QYiXAMme35YHJr16Hw2GZtuXz7Ea3Ai0X8VHJe1oPcdShvyj+vuX
ibzAlKStme2HvE1bdEo9ywZc9wnDL3OG0GwTt7hNNgarYWhQr8h8zp9f8yIvUkga
FE471rn0wSXnL12y/58fn4eOMVtlOyRNRXa1vzfbcUlbSHSbosfZBtT1UlYMFgcL
8491DE+95CnNlDb2uW3Q2xvNaq23fLWluCCtrz1KnaUGMm7/T3BKOfpv4d5QAj9g
TI41/IuS+3vI2ys1sZuzJCOwStPiAGhq2c9Ub+iyxsmKQx/XujvVr2/BiWS1Oace
A13dpgvWzTytWgFZOgvnqVQ+kHDdbY9+rOQTFviT2h3hXXmC0TQkvOIAz6S41UQd
t/NZozdEhV8d5sjldoa3DFDR8WiNWDCodAQXLS3KCiV9R021SpuLujTi/q56D2Dw
f1xiD8Rn9NvXHPDVZxi0TO5IiiOKGz8fzLzKDYLuH65E2wN0r9J/g6bU+bRlM2S5
TEpdWedTWgHGbAsuXiSBX4XDozduhhbwa6c+1JyPNcrRESAH8quV00Maxehbz4p7
1akHWk3HC+jG392KHcTjGbFL9t5wkfaELimbLih6kBHTNODpHChRRvFPQ2KF+QSM
p+m/OV+wpwRYPKkVKoBwVWyd9IGEdBuJ5d/8BFkxTTsJP5aH27Hws4ee/PHl9dOH
P1HS1mQzGlOYDYRvlsQHJ19Jbrxw9ax0wskqH7s3O6M6ORALs66Y7katISBqW55M
Nihn/bPUktvEA+dNl+k6X8q3U1l5qGFMDAHHQ4Y1Uj/S0nzLBXjuWmb8JtQUzrXY
+kZJn8LfhoMOS8sCHn+q3Vivy9VNq3qjaI3hZL9raDOxP5XPaZcDJLGS/GeTM2Ly
3+SgLIwoNJcrJCPOCTK4Xr2b9fuISG1kclxDmb6QrMnTgIMiPvHGVmBwGoUwbzH3
/cH2fjcDdlIFHRt58CDRBkajrnjLBgJpLhCYaNaN3hWruWwNfNzoYJMbfx7Uln29
4npOyGQVNJZD5ul12PaC3Xu+cYnAffpMg+cntQRmd67VDIo0Xp+aC5aIwbUVgALT
bQysmLjghwnqEpMdTNkR892ylnTZJwOxmaG4u5QXv69GpAF95QDL3dKBg1kXr/km
HFN004c39dUQpfwTRxdmdp+cCCW77VZn3H5Owp4nBt2o3Qd07p4Ch1pReThjQ1t4
/uuEdDrgkb9biLbnO3jXhEUIchY04fSYRmHpMy4fNqLaIxhfAt56yxBGXVzv6rHf
jRR9AP4aDopLK3fmJ4xmP0fF5Gumqzs5AkSia75aDqqEMv1hQShQyyqu7hxiQ8JE
eRuCKSQD5yYjJf7ogbZ7qqCcVc+/8ueFiJrfINcCG6suUNiU4PxFi1skScUmiqcS
EPaz0qvN0zr8d0pswoJdcRJVggN2V/6TgNYmMyfRHl0rm+35BE6prPQGyX3pDekU
0mgTqlzq0QvmByVMjobdpnR92C/9cTOIVpFnAEpjeJTYrWvUL2dBGY6jCdRDPDV0
lSwfF539A1/WI+8tupYNGiXGvH4fu7N0Z0vYGjqk/3GYsd5h2vzF7RaypZqIpd0v
5ESSBoQ/eZ09Sw1LswxLO3WeIm+QAy3Bnzbu1uV1BFgSx1S4r1k+hZz2ZNnJh2FE
WD0ECzdHsZ0lpHbwDW48nbaFu78oQJVSMXT+3JsQ88njqExzJ7sSGl5RlvZXViYJ
v7eyWvSV5hJ0Mkt9WenRuWsjhvR6DmfegYDVSf0xqsm9Ws0bwXATwzKwY3zT8cK3
52HYw7GxID2xIO6oeZIe1l5v61phe+BCgCd+uVwZ7SwkGGugwLT7a7nbXTolOZcj
ElOYHot+23kKsYhK/2f9CYZDdqkE5r+hFwMnYiqWtEmYl3HpufR6edM9aF56/KHO
fzsMvSbCk/Eb6VV8eBmtLcIlNdG0bpSXexycHeECVbzg1PBBV+jqJ6M6ZTPfKdsz
OfLHluQel62t/o7+7CXU5VPzFeaUEPFLD0U6D6VRJRxqWTJL5o9HpGYKnCA59b1V
0qJ9RGN7Rb19+T0KhZie8NhCsEwrYTi6XDcrph0cIpu8gmMKuxzFS4I+e2x+FuvP
X+kUednbN+/zwgStunVf474+q2r+Rvvzq/tsw4nTSI1Kd9AGufx+y5WyOJJXHf0m
KXiQmd/7RrZgLmmv3Gff6B3k/nN53nb8x/LUq1zjaGUoBdp4SpjjEMfNB5TBYplF
HrkAKtvZrDee+VuPBtGDCk3rW/6tbVcm+s6su8b3eVRLOBQrUHHfgsvz3wD1J5mk
q2wGlwE1TNgpaZ7qcDe8c0pRWRlIA1nLI2gXOEG5Hd12Oc6+ACdccfuCoL+at2iE
cY7me9ToaAcvocgFkXoHfqeISG+Xrb7jCDLN6Jg0yIhWGDCqEDUp0a8kQqFzJYRY
ZM9jcgfb3F6In7mxx66FRDgu5FhMYGafJtSLxjek1MfUzbEWme6FvB+s7IkybeXM
YtVOJUSDe6F+fbo+baIIcsjovBhIo4TnIXPmD7zsa8BfVu5LGLWDwm3Jx9Mx1VcV
a+9PSsxSc6OXkcCEjVCQ8LxVcHC1D01WCWK2/U+dQMIDvzC+opix84xBVw4OoyEs
XgJPnl2BI2LEvQpLjRQBE7nCYhqUurhNktrSd6Rjnn+T7xmYNXpkM/3DRHKWtbaU
rrbVquVjnV8IWGuuI4iKg2sgSMO+e4VWd8E1gML0/IPlARcA15uJkmgSE54kZeX3
n4VdtaCUqUU74h8PxurUkuc1YvL/9nhTyMWVfh5ZTafHF/KCAsKpRWWcjESwfjqH
KLPQC0PMC8mke5/RzZAndjeI0Gjmk1+3O7ImmD72gyRv0JvumLw8bgFEVi0J7OS3
xmdMut88mxQeGJzI+fPcgZ5S3dSRGA+HVKdyZS8TExrGjXY/nFtYzNYgU+7s2Pab
HL3eQxeY1bLis4wfu3c5m0VxswhY36BXEfwfuBqWb8DryookcHyhOpOveyxURw/7
MV193gYjuXTzN2R5rd+6CmSkVfGT3p9QC5QmlU1noRGlWKmbkogFX4kgM91nm8o/
3iEbFUhYMyhFFXWT+zibLPaX4B2qUOs1ntmozTk5P0VHUiAxiduGtNWTsw5ML818
Udz22bwgHRKkY87/bzAq5XCP6wTSrmwxwSttkJaX5MgVMJmseZkSnbT7SPQxsI8L
acTFMr9y+gfNqZd4kWpFmzs7bKlJAST+eZSqK24tZ1pLC+5c1JDpbDF3/8suDBBi
YPErmrFjXTDmW9Oamd5rQ9Hs0VHW86P9MXaMp/dFktHm6T8T8yM5MSd6TO7pwFkM
1EAhMezxgRIGMzFV20rqViwliP5SueOVcqmmBpwCmGImwRNWoNxYXEjlWj4Fpnrb
Yr1TCxo4BLo3z5aKPDERNY7U0Wbf422UeXtVtANPIY99X6Ae/byCm12rA5hgbcl1
qL86tSBkVvvgpJY2HxOhXG61FA3wNlSAF+yH4iHUbCWxFWtg1k4WsdRvaE4GKWgc
1p1yD4KeiGHOwGZwXRxYxoXZYERqdqwtImSyHWCZrhtXyotv022Cy46SyupIYxwd
HiRi5t4TrE97NoVWNzJjtZmCovCdCcY/FphgiobqHJGV1+JMKaCMoM/T8WoEaRfJ
w8C4DmVLglenIGElYd47E50CtkqbGb4Iazt7V+mMcSj+Kn6aMrvP8DTz6QyErfjd
dOfA/jm9H1Y6tpSlpk5juoWCfoyBS/hJt2ucXIv/cOFjCK1D5WQvosZfZ1mmPMZa
SoD7zJVwUJ3m3tpQQMjqOftvEoQuZE4CtW0At/PZaaI1UoAOk2Rso7hllSaPwbfq
zzJeQhl/Bnl99rSAU1eLEmsspB6WS9tM1/Mz8Ylno02qedWcg7Bc7txhZU//TVNU
w43QVhdGF/2GwtCGuy8N1vWWbtPDgrS6G17fCEV22rDaA2aDJji3QdlZeGtVT5fp
8KYELmbukaoVpSqt46OFy7worbKoNHYGRDe+2lRVeY5eyFirpDtzmFVJKjbdGALe
Y7jiCQX5e/VCBmAEFXMvlYcc9cuuSYhl6DXQvDNmsLGLWRJVOS7XR1ZGryK1umSA
PwXD5+iIfzuw95sw32EfqMubeO/eiXIYH5RLj9k7ZbVmDyouEYfcX4fvnH5dGLqd
bEszzbmwRAoO2TzkDSV3AsdcuC8Z4fAbwpX9JsDdcbK7kTBW0sThWrNE8OtQPeOG
5qNpXy6Yejoq9q0haYVcMY+6DMEL/OAR7CFhOX5WVlh3W8vFR8NK8IdjQh4dhMIl
+ddUb+qebS+c6cnSa+YdKjGTVn/kWt618uXfkjY1CyZJjKF6Pz+PT7uSJKFXB+6m
RP41tsJb6YClg7/tqmuEsK9xJJn0x5z7J1bG9KaXPPFxA8VwbkOJuRtA3Szo8HPC
YXvn9glgfBG3R1f+ZcHGKSBhfxMB315YH67a1FnQJpFnpozINKKZ41eH5nd38HCz
wbi123BI4ch+XrFWvXJikR110nudy/PilXNOLATeIVnB3PRPQtJgl6hQnaFRwRVz
d5EdCtD6U3Yjy/l/sCHX/+gx96pgENIVRvDojz/66dPcivn19BTPRrqnZfJGnVRi
bsQF1j+d9TXoSmP4j4z42e2gUgRAQo/vt7nT8F7s4hEuoGUXS19S6v2gtNqiDEeE
mNAOF+BYbVED75w3p3sNvR5l/rEaAb9uI4dpIUcCJzh/WucavcI0faZxxnGRFlfg
vSM7RJcdC6ifvR+D4zYYbbi4YOPke02kT0H6l6tkJvK/YMwcxiFSEaar9lBw+9Ev
kKFK2scGyq05agzVP0S3YVUOHHkHwnm5jFxa/MAa7qBZ8LVXaoD/VSEeClBVkN/o
4qnO2cVjmlOJgsnbFYkLbcWFX3fvGOgZBeiWxOCzDJYSLCCo7OJahrDx8NRybsAG
BS9UTlTQ75Y5lHZVj3JgcKrmHP//sU7gNsrhOLXlapBaa6FMZaJV9cPJCnLehbsq
YxLSOJFqJlrCKWvqyWd3e/xo2AdAPQLmWKAlWf/hSB5coCLODM2pgQxX5x7Pj1qi
ANcf3JD5v/RLqOF0i4ia7q7L7E0sc6L7s9ZwkYTO2K3XGzBEJ36zuavZg7chjMVP
m0GS/xcY9iMoTT4CjUyL4W32KA28p2fQQKM391z4Cj0KgIBSORlRYIuUpyIjCetx
JZrIdN9NWQ/1Ma3ftSIXVqjNQOSmuTmbglsfuvBu2SQuiTk58ngiUwkayKj6TBLX
Lxte6trnA2EVBX4r4MIssPAZIzjBZA0AXOJPqxgcDR6UG7v4vzTDP9/QbMEd03gF
nL7RgRdg2sSoxSHVbcfSejcNNa46s4RebIOdlanBGFPiXt9rksGV/MWCcddKhLVM
V0+BapX/jJAGrJkk320LvMBMXEUv8vnTQHlxPy8yzNT/pK+0G5cekghcB1FPLJnI
LgtkBYD1MkEtmWSEamCIu7d6TL6AbNq0Vt/+O2McmBKaQhNA3VzqnVx5wEgBLqKV
5KJzod2CPdg1TwjvuwCKV1EVhxtMgowG8qA7089hMLlyQPaqhmEPud3HJFu1VVaH
FXJxpsWClYkal9TX9ZnEQX34oKmiZCspKq7sTtsnJyrVvTQ4AEj42/iRn9ArRhyi
3Vnu+4NRmS9Xp2I8WdlPlZO17+UGPKuirXMaE2uG8FGKKGvfVuIitIA9IE0LTLty
BeCTfrf+VKeTmX0vNW0AOiGcGp0vJy+2me6ltTxU4pz2yYL4csg19J/lXlGkl+qd
4NSplmQtp1Hp5+DcgIgF6qeKOUOj2iLz+Vi7lf7Ny+g0ASTYi7SpPJ/2bWC8uoNz
b62IP93KufKe8XrULH29BMpuj0Yl4lW47Ew5Io18SvySyXxxpHcMUxk6YeFpBus3
GiaEAsJHqtoW2YyhP59/9dKd0t4FF9l0vmtK9MZ95X1gIaCwGV4ZXWiN2tG6zbeq
CVpCuO4PeD9XrJX4Lio0HR4Eap/gvwUNaxtT/cBvX6A7orhTVK64g09Fq4UfvxrI
uSN2idTJTON7IoF8CN485Ur3fByKt2kMxS0mfwYoaBbh/Vjc94lNqNmIPXQ3toUk
hUb7O9QnTKHYSMD0oct6j3wx7qcvyb3gCOQMosojQq9kcT3afYcvrC2jHx1824qf
AXQ0sW2PcrA0KnZ9fwURbq/qW6qQDAn76e/nk7fFmwrUFAXwTR6zKh8przrNu6Uw
JdBZ9h29++VvCUnI0+31XS5q8d9ztdX5sudbrI4tdFciE1FYHANgO98SzqXdO9a9
5DUGruhGPWopHE1kxhLbUka6EP208+fU7ZjP+GfbXlJjZGC+KPsOOs47D2JBbcLx
0GBY8T9hoK70ON+05BNCPCMLRcnVeopVZs+rYaXuW18aIlS3zjZNG3U46NJRLJdy
QmIn1uBVlZQpgVBqoz1fzPUIRM31kVdhoT1AKyTeckBoS6Iz9J8WR5Qxjb+Wogob
BJfztIKGE3igsgXZd9gO5A7PDfwRpKc0GCApGDZYM2C92h3D1usM4BaPLn+2oLwh
GlZCjxl3AIcHDOAxih+aLLgoF2D9Xb24ErjS7W/DdjI8K2vWZbgr1KyyleKvooEx
BlTqltsD3OsRPQdzX7uXE66doY+BsjuvZRqaCypwHQDi4vLueoeMHdNrAWVLMat6
FLcz0paWzWNOclAzZfiDUO5Y9LqXcecK4agvujIsfRwwjd4mB0e8zCMh0+wp/qYP
dAO0KlkyQCtsOBQdGE4kRfgsJdE6NSGt1etOpb2e0QlcZETAfk2EnT8+wvWtHg9I
5mV7yTBv4AcoirgUJB6PR5FouRAc9aHV19P6jIT84OntZJhuXcFPRevhkF9SbGD0
yp4a8xER/K4ajnoCaYGSYOvI66EiBDH/YoB/2rht9jNfT16FdWDM7VchZVkhTEYG
mK40TU7gZhmgXohI7nkPvWVB6Yg8Rc0ulY2dTghvO0iyhULMgi28n4QPrj/d+S7X
DMZLQIuXUQ2q7lCgupEtD+dWUHJuofACBjrvJjMxp2L59DHamHjYsFxtnWCa3A6d
JRyLzjcHnkssGFCJXVl5o3kUwqxHj3ryhr8PCnu+YoQ7DVAA3LEyYWmYl19Bf9rs
CEVN6GY+afEJ1bcp8P+4DgTF6umm4mgI4DcyYL77kJV8wYwxoh+vkZzpWApJH0ys
Agd5EHVfJ1LUoswCKMZTAqMcOPubAsGMOLK+MSBzj0xy/B7UDdViMCOejPrrbyLQ
Mg+xUX98oFjTvsDJ4GzOxFoMJ9qZF4uLCUBTbyVGmPfNOJvR6KkZ5fIDSvPVSKs9
ytffP6Oq5nJmQaY4mAkEMzfFTAA9kq4JF9ojRFf6oP/lhP3BxiPSIebYeD1gS8ZC
fFG7MU2ab88ZQgsomjADqxNd1tCHRCxSckf4f8DZd97z3msXUwyPKs4NzNmvs7hu
4J9cW2cUpKwO7X6zckDAG3Vk3kNTlEhmBCvDhhKjpBQ442XGvVf+/qr5BI+S/vr6
Vi543AiWhTPoLN3Ks3E7Uyd21yhxc0DluWUqzRJUf7wL61KIJ97N5ttuCTvBYv35
R2XX+YLCzLj8kpUsWpfpZfxowRPD0ccy/51ZbGEdYNve7oCUFMxY5Y5Rc44Lq65k
0V3iQiKkO9DduExumNLMs+VTxc8ntJ3J0qj8j07b3zxAmuYTZTxQG3rN3egUczj9
/Tj7MtQCzGuv5tOI+zmR6Pp5Yc+GyvhT3cxtIXYPw0mLj9HRmhJ/iU6dVhtN1rey
NByJEwiYpNKxnBD15sXE2JB9mJikLdgZKuTM/KIwo/A3iv63srYoWJaudZF1+UOX
LqLDFATOsPpfgXZ/XyivqR8NCMpchBGwS7Myccina7uMlRJXYMe/OiCxnz3Yaf6V
bgfE4sO1subvgqCEBcmp5w9WM7TIoSL7F9Rk97n2RF/yqLehPFBt8+nRhmxOriiW
hqmXUxMjZ4Agqq06rAnxUYyx7/CrMyC+xOVDiS+Ty2BLDgW3lgSPMeKH7Jf6iubE
7BFJAtqQIYlwpEDvWJCcKQluGYDxraKVw1dFSDNFY+xtaVQUFbMLZG8zAx8WUHo2
LYmFSQ+LCEZ5B9OzNEXWliRqzhZCdg5inyJQLKwys8d+zemK6G3EeoOWOw2Fw1KU
tkwcWyesLPE44gmNEppYkZ7KN/kjxp+22cprOjFbQiSztVJmREdfAjPRrR5U7pIL
EzeDrd8VHF/bIqakMagtGwYmnhUvUOtg9HJeyODlL0Kwe+V3YVbjOcNOOZJGliTX
isKBHW2br8iJHJJepYgd/N39zotYMVeuFvCw3nJJVSg6/D8UysJZZ3L5/FcjABiS
MNQxJF1W0bIXc8ycWp7aDc1lr49p4jE5ealeZYQ0MM5SSq9sEzWEdzWcrHkZTlYm
ec8xfKwGuAWiyaID6AhxZOonJRTNilo6K/F69JTrcEMcp1NXfWSh8/2jlu9vd+D1
Mf8xMWXtIkxLP4DXo04HrGL0pUDr4e9OR5DWuEdew+dP72rtb+7vAPUVu4OMcS9H
gW9mZ8ZogB0Cf7FzHTjzqNUye3wZ0uijnwjvNOtKCvtOTmDdL1EWcgJ6FuztJsVe
x4SortWe/ztsoTX48i05dpGJCAjmYt5Uatv5HQ/kgO56e7F408dp2QSu3+dENzkt
mWgR6DJle17xeKYiVFU38bM2Uzeaizs1H733iXaG8Zv3Y13xXphapzu7aW+mOugu
9JVVbOcjRW3c+Sdjoh7ASJ4FiCgG7eOdX2RXSXjUQo5bHJRgYsD/HYhVDtGnxeTt
VkXEhkW6heeaFK6FsPsOq9W1VE/Sga+NoygFobCs1qRcNHRW1p9+NuxgYkXV9PF2
22nu3Q5k3OYOxq0rTGwUjOl3MlN3iCP52Cide06r9rhiP6yp8upLZtU2NIKPKz29
C08iboEKJuMlMTrwQCsRM+O3tf2VKOAJCMhT2BJcyI4+GXRK/zacfQJgLxtLgZkI
nyK/1W7I8g7iulGxSBvOy3qqGIn3X97Fu+MDEMFCGGwE6urfMIRha74AvxPQn++G
ytOmnCM4ZuhhC+ApQVscBDbYh0TC5iyDrqNOPwaPSBhVia+bBvR9LKtrj86qJ9OM
7BMZ90TluoQap8oM8HSjYlWXMwQHe9cxz0c0ym4ZJobIICYsfDWM8ZoQufpHFxDg
2rxPiN0ABcnRuksP5wu0N+FpjOAR7MdpGWJmVJ4o0FSjYe3JD/xHSXBFkfY5Q/B5
ElKeZsn8f1fgO9NRcZ4ZzidO7Jfaa1pAgMm49dFoiMum1221yBJIcpX7iBMShNXA
NOGAgFJZY4SIU+lRmryoU05RfJ4BeUORmHVvMyvqICFITH9OlJ/ny7R+kB8Tdwag
+O8vP4mgv70p6L88I6+ITeEwD5MdEP9nTbpsxcSY+VqjS2fHAVMmddMwBESwC2zx
PgmCK+lrN8jRVLfS+8Flx8/uFjCCZMBA0qFrfVmD6PRRFOe6MHFAZ5Ay0TxVUb17
rmH0lsmdkvSISP7v91HiVripawvies6wUngkP70AiF7CWuFKSEzuJwlQINNApFpk
dhTn6tBBRW5LGdPj3NyVZrmW3+xWFTZdj3VJ6dqE7JNHHkyhKEgN3ZkuZ15ND67P
Q/1HX1Pkueu/WCTVz57UttDVP1ccnHZ1oTucVZ4YFI/nOk7HO4uRj890XffJ1fKs
U0Ph6cgYDlWDfmS/0Y+sSyrEm9HXIvjLptlWwPUESe8w8J1M/JMoWrU6HiESHdgU
jgAnDI8NSy5VLa/SvYaow8Xb1SMgQL5MU2fj9Ssbo6bwWx9B03Frlt3d0a7TzbCI
SPhHY7gOanXb+sqRNvM0Q0PCPBlmzrnSWAxVE0h6heL1muOi3HfSnQ1n1qYqa5wg
/oCbbOs8orZbWUSPPYNV8/BOV1UDqCclOd049l9XNpayDraLbYaodHPh/6NKY5q1
DZvEINghVfaE6rIhbVZ5QCmOj7yTIr6YA6WOfPHGjpAxng0fefIaXR0MjrqbwIP+
j3FswwESMdj8vH7+aoiZWyAqh+FcQUSE2zqL1W+gYI1uoWPB2cq+V2OM4kuAzyJU
ylVewJsy1mmh6Hug92C/JPd4Dbd6GTQBxp2E9lMLk+YP+LlKig33FGxQBDrRDynz
dwjrqqn69uM+JtN67UY9ZPXEOUFRaXzh6zr7693JiGyL/A1w//qqCBx8nt0cHSQU
G/+81feKqPuxpgBmm0Tf1sa6fkpADhdRTvaoTOob7A/X0wuA5HS7wyZSYJ2O4Bo3
JKInUauATa34ynlK2/gXvPXw0RjBLLNkxFEWpOF88JYBtLeZTrcGI1iG7G+JRaiU
oazplfuZJZbNilg3yv5zf/Xzo5L20i/OCgZgF6CJsGm1sOzIbsX4/1RfvRBdtBdD
Cy38iI+WAYxY1LuNH+tyxW+wNmVczbY8Np940Q6kqt0SQo5YtgpUmgv3s58Y72/c
Q799jdA2eatbJpVN4foulp77lcCdgOfU0WhVyBlMZNEXjZ9ptaEyKqXhanunZLps
EL9JpeXvPG3TQe+FRq/5pA1/3dwjXfap9uaOxv5PRhYNcsLt29ipWkHeU5g1IczY
45AAdsCHbjoRoRhQBMqJ1Y3/rOEJyM3SeISVZS4vOjIJX29Tr/xthpNmahG/yEVR
MRQrK2csFfpow1SChjdo8LrR2EoFZ7BbsSA+LX8nLaLlXDNd187wkDjDPSGQqW07
ntFnCc1ekP/A/aACFUIjlwPL2XV/0mKXbBM2TtVn9hbfaV3UW+YHif1tFDEw0hbR
y8it2cNrHPcnsm8rhEHTzMrPcEPul0jfAjadUo7eyEsS3kX3bpgnms3qMlP/5sJk
9Xtgx0PNeehnDAwmMWIfa95TP4TghBamHSmWDMtJOiwQ6Iuo+T5fEwr65ScPinO7
J+HXlnsalu+Uo3JE2U2zEwB53184qhiNvWGN4tbykyOJ3dII+O6zWV4EEOOVTKk1
vMzngJdeJfuisWUf+3/PLj14zZTmVXnw8cMWt18b/Yd8gc0VYElCw/S9REbTipAa
8TfJ8kKFKYG99G3CfKN7XgCTClchh9EWgKKNUbMEGoeDi6Y4QezRzsiIQdLGWJxb
ftTP0bYMEF1DkBjKIjkMeUHUoqMDH3S3RWJEnuZiTOnlZ1gCu86nsUaBACQIinhn
vF4pxEauh84wJmksDAT7xWHh5+oZS1GqLR58uV7pGal9XAGGd/i8wRSeHahvh5kd
X3iYrCC4iBPbupOk1mI1fitOR1yTl9RP2f5shoRUehzzsTrRCnKfEREQwHNTuqGD
wrIMX/qqCP9+WMAmgzcrO5++9qQV7guO8m2bJ8Z9tcNCrZsf18hgqd9CJjTAeS4t
K/KR3W09kkyxWGJNgZD6tjPBM7WIzt1gTsZ6j7CJR0AxCxWp/ZyslfVfEGny7KGt
FVMkQ1p5Eij2H+RE48rhxwOfkhTyhts0SlUuISIZHFWgW2QqO+pngpgSMZ4e7u6A
SoZijHzs2epyrv/rE9zfNn3zaVyr7NG9GBtBYOFZvca/LVlY1eLCL9zIafwOUP9L
lt5nsOmuoPCzegBG9ulbXD1PPsZPpxYTivO/u/8ZT3slAeHrRxVhrafPZilslngF
0h6xHPm80fI6P+tq/qu698MDdo371c4mIfWTv0HJ0zcpkyOiOxx1x2ophPU4WCu+
ZXN5XpyM5yk8i23/u5yzTT2Lh2dmS1d9zE5Rf3dj2hHyzDlwYXTuPQnAls3MurGf
mztpE0izKVdIngZW0E3PeEXA+Pd2USBA9cSpDgIa9U9MTAS4gPcLpWiBJ/c2FmgC
8V4wKjY56noI7qXvHoR4uGhMBnWB+5VathP80L46XUR4CFBqEdb6SGTRNNi/oIYc
smmmXKrhBwUwN882PMjoUcfH0SxavZaHJTvAgGA49aSOKtwwBriX2oxgMmpcjzfE
kaZ+vJxnlCV3jeHF8mQJMfnLttYe/2i/obrfAae/cO037C4BlqznxjuHx6GOKM3R
z3LBYSrWlN8a8dPeZHuuswO9NLLy7rxJzce2zZE9mQjhP+9Zl3pUKZC94a4wVNd7
lL8hZSmhV3OpfK3i/Ppo8qj59O2RlY6L4STd8bPhBmY4ck1HQ+pKSY/kEqR3rfTS
yijFlhIBEgEdNonfXvFnO0jAewhCu0ShhVgPymcvY2nfMoEdVR14QhMO6gUKenuk
6ztXL/SR89lLPE3Px82RKoMujF/+wBai5y4AI123Kqn82yx2TbEL9ItGmSGmysbl
n2KffFS+JQ9qrgnLifllke70yPs9wNqfxqhuFCpNk5xvxj/49l9JH9Nja+Nn07ts
gY9RfBPxPjyAFP7t0CGL+o3sKl/jGh+A77ay7O0EVIBYhYqkE24YHPCy3oOT3ji8
i4esytGPDj1X5bR5gbtXegviXN9NjsrlKnw7RR+tLhCa3Y+CU0CiNBtXEje1PtFx
R/01eUQaYYwoTiahXIzVr+cNPGNp0dr2JOV1WYTNHRth4N5iMZGTUcU3eHSkcKMi
DneDlX1BYYwlp4PM+kalb6DznMhuC2efbSvLfcal4Cv4nBmrkrOfvghEfYPRMfVs
2+l4P57adMm/0e+nDqtz2aU52qzD8BcEmR3Z9DgY97s7ZWztd2FpbMfPlKrEzPa7
W+d6nZugLPc5MCr33DocEXtifKc2u8oGzE+KaweUdAkRtWPnpymPVNg+ulTwzd/f
d4hjWALxmyDQWdCzp2ThZpU9VHr1A519wlhKKh7+tDZOvq/VFTVlKnq9bzu/SWca
JVYwKmOGu8MS4EnH9lo9v8WgfVLCiwl3fCqrpKRVmPUZklZp9tQ0auF5heKxa7Dy
5G+ZC6KO4ugdZ0kNhH35gMz6J++xuS5Tu1QVw9RVlWpm2u4G6ApFlFjezQi3ZBLW
+OAXMb/LIAWcO+LTJWWkUO7hhU5ypdmnoGKrhR93yPuSLPhrg7JbQWN6LJ2lbf5O
71Ny2BBu/TLZyvALW2LKStf0P+dqH+aWEJdt2BkA64jfwpUyalgaxvjOPbuWil85
t7B7L/ZjHkN8Pd1RTPbmZ/nYSMH23Inca2Hf93pXb2fOvCqwcU+vTwj/qpP1Gqn5
W/Oyot70YcINON6lZLi6TX8lK8OEVW/SF7VABh+NoGmBWIVxsuk+g3ORbETux+tr
u8moK+iyXWVRUICZLjSoeASIGzgD+seuxtHik9NDL+muDGhU4Paw5/PM2OQr2bDU
A+tXK9fLzRuIK3JpVbIqY2sxEHzBVrwwmkCL4YzCIQl/pwGnP/DyEBagP4Jp9ttN
8ni87mpu6OP9FlS+DAdlVOAGlhlAFbKrHYmL0I8hNRJFAJRFuy6iDNe47hVIDEts
td2j8uaEchWZAlA/S8jGU8r4Q9SHZ6CcCSEAge+0yd6kcLHEcSGVTwGjXBnwOBSi
fMd15jTCQpilQMcdvWPvxTfQOiXB0iBDt86H+UHzSKnu7L8thti1DfMjfTP+5pOK
0zvk7rxzt06PfuMuuAlz4wm/gdmHONeXVo2jluSoQskWd1+DO8kIxyv0QBAyIos0
FHEsowFSu3sDfivdxghkhH37JuajdbUhCzd3m5uOxki9/n+lTCKqmv8Mj/Y9AjH9
Iu5gWFpi90EUL5AfVRLq7uqA90Zw/MmR53QyC7vz5ITD7hsxBQUm6a7mXd3MwP2x
RwN7qsJijwW3zS3pHALZ9IfYcizSldWVNsQ1gPSQUlxO+RWqv0JEeSmUwa8YMO15
fMwQIs7gz2nfpxkskN/Z1AouqexASPNdkWeEgof/Q/AMfHqnyJwben8CPFX7T23y
WQpi898o5ODjqEj+8ogWWOt6T4PnUOyXxXD/g54tIQNLaUDeiNxaDVHV4Gxd6tII
OthLK0rl61m4mevuaD1Ed7hNyEaK3tRj13O+UGKjhi5mY55+PkTy7oNNHXTV+kMP
uHvt/nmb2guOp8481alSEB8QoiJzu91pPK/m4WyKL5N5dJpSPjxVKBHGzYSC0beI
GTQGpKspV6wht3oIMyEx+oBTQUok1bk6NN0GJIIRmk/zsSyo+u1Ug6eXSmvDcXij
1s6az2muysBY5KE9uGfm5XptoS5oPi8InHrl3WMIjsWScpY80k3nxqGDjjawxVdz
oh3fgGgtz+1XN5+bzy1fj60e2uFLG10tE0CmXMxaDiO1voY1XxkrVNDBoC9XNDbe
EKxw7sGCBIaXjyaLhgGErmLzervIR3AEN6q0FkN7JeJWMzAWqLODj/9xx9ovKDUN
dhjLeMVswY8KU9XTFOYhuImCIpZknBn94UVlOWEYnyBJ6XWghJdvTMwtNUMGuYBM
T8ZeOKX+/SBEsP+w0TZ4hPrRRIYkL7/BCdhcbHtJqnc5vdvTfqAu+BdtvSrUqFYB
LtkBS2/5Y8yBFxAcvptoo/0qLyd38FG54c/rFaOLmTXUAa0ZsuAI1Y61iTCI+OUs
+6Ug9st3OUhap0K/e5A4sFb6N4GWn9zQkLdZnpEUqbR2Jpy3SvMDrNsWWypghIcF
O1X4GmK172D7RozMQkGFVYQox0+snV+INzEUENjr7Qec2FQ+kp/ldcGgPDiwaosk
beT6Ta3gecYnT58aTyg+rpbsS7KFnnSa+GWUOl7M0w7MeRrEAoj025L7U1zeipbW
bjMdawOZQW+xUAqT/cdoS6dG49a2uXYeE73GHHM6ub0mDpXDjJvkxAV+o+xsKn/F
VBKKyIUe/4vf+Du6yEWdldZ61JtwMM7zOogcI57bBgWFZ5RBgGtSGdTTzn9Akgqb
GW16wikuNwgM4EP9PzMaa4H9I5PWNSysc/Dct2KM9oNZ7xBf4oB8oieNhrdNVXsj
7jqf1vVgtcbIDJt73U91XFCzzPB+7aLt5Rjdj+/qD/mrH/IbKN6HvetKyI/CRUdm
Ke+GaqNrhOSvWYzdtqmJBDXUwluyALXvvi1qS9BVXBCCitSTbdX9IL2VULpWGJ9g
i/P28FOf48n0zLbEDIhwyENdQ6KGESpwMBmTCQfng2kCHLz68N1OFPnDgOFDyPgS
uUWzxrgBdXqvu7+aQ0DwUprhgR6tASCfQjfrA8f8LVUcqNfWBvPqrtv/LdiJ2FIf
O8SV5kaFUa/8jbOWEgTT+feVec+Z72tX0CX5615krT+RqjOXbiDaaxTGO/JTrQKc
qeLLH0OpHEoVAGZe4RBjFpMqOuyZ/aQybTRB/9N+PLeJgRLZL3fiEYPB2BBcsfoJ
ezaTCtuNSv6c9TptpLd2wxSPG/7nI0jGheKNOF1udYXcgQiIh46y3ZNkL6LW0oUs
qnBReP3Vy8P6hIR728MFCVPOQfortwg9+vqVttdinfFxPqXc3OhMaZnNW3Ugdbd2
LTpa2P8zDelI0kOAWTGg3gBC1XJC9WfTGQPa/Ho0QxP6V3eejJ3UI3U7f55p3KSA
q2CVYHpgIejrIT9uv+MX4/aDlR0+UlywNetVkRCNTh9ViO6bfdad7SLnTkNNt8+v
ORlOikmr4iT05te+AaD43lt6iymy5VfsPIRex+nnk72ZQ9ZsL6skcgDKTtTqaov5
vzZV0o+8/+52hqp8mp9CfcQNKFFg+cpi4WxY2wuIP89BkKjXDv+uNLmuU8241vr8
Xu9v1zlk8TVvE+XwPKXIQwsKCdXt0bGZYQR+fO25fubvQJccqpm9cGzbz8lW6fM2
s1rECzFj6OBARl231S+th4rnm0r/qqh0LyCuNSR7pSd3R5bkEFDJhLsHv05SXu6d
2817qKvKt3m40QrEzKxGRzuOt/x0H4PBvfrEJX05LnEbwP5PiXUUMFJYwQNceMYW
TA9J7QCa6LlTBZje63LHKxHSJ+NAOX8gA8m0EryXGo5vslGvTmOmDRhA25vJKYMe
68XBngpiSRRDeEw1FsFS0MK4HUZekz2WOaTJRj0JVOR9qnTU+JBD7WLjalHGfKv4
X+rihS0zKhYGEqTlRVRaS3YXehLo31bUSNA8q7q2LvXyu9O+XFZPE1RHmAfUmsS2
ppTh8Et/RYY3w//ZcoRVFDXr8BrtCiGeBETmYOc+vXJi7TDDsFhFZl1d24xVaZlW
8bA6kRrzv3mDZaYNFdz/MavSIiXpQAnLwqecyi4BXAS4YCQyUG/I9S3eHMJJldl2
Fe6B3tVyQP6Dm6pO5DjhN7fTp2pyaDS3xM/8/TIuOpjnsKWswRDijxnzNvOHvwby
MJTRkhKW7JBs9Fj/jR0dqZtmWtmmWwbCd90p5xsjXmvZFwacKAz+7TT2qfsvPp1x
+Kf4fTB1XjzqAMWU7nPsuOGi2fEdrOM8c7/Bm/u8RwIR/oHTffAwhNZ9nnAt31+W
QXP24HdLaHbJJywd0aL1T81ttjB9xlpJZ5Mwik3u3oauwzYn3qaH+gXNcmK522+J
ZAmX00lN5IfCwo5I4kyNKXxMPS5EVowUx4GmKiR8WB73eYmlok0CXxwx+n9KNuXF
U+okOn/TnvJ3iDUzD3fEu8ZD4YsOc/O5aF54VkB9ls9ecIoR2BQWSAMJjKo44Wyo
lDr++ITTYAdu2NFKMdxtPZQxPkzuCQNGa38Gj7avxcii9JBwIwRiusP9ot9/++Ie
gBKIE4CD7+++kSER+1YWSowzSbMC1lRoDcgLnp9NZabim+Nu/Pg7ywsZPTIAHpl1
oL7oTX3kgqXNYHuwxFnfDJJOu4PR3THIXWXDAHbl0HZbgewe4FQISjxouPPcdPtw
EQWXITP5Sy3tGKokbjv5WmCK7Q9SJkrOxfinmV8B22KP9fsTOOc7EK7roXZCVr/O
xktjV6CGBIWLab2ueFNyJRPdzkPY7IruCUX70UrlLoMBSkoPwOBd+pLH/8yXeZLt
b1yYJP1Sy8B2WEf7mJLyA9EAJECR9kVOEVrngjDj9mKOOnzvqS/0AkDEK4RXOo60
Ty9BQIyn+cyDhSeaJPqAD6oVuw7VOao9hPSQwdZ/CpMO71lvqhHvlyNmAv123RqS
VL+QLrWc4CRe+eZ3DRtETx+5kdpeqGhLaJ50CkwGfpoD1OUja4bGvPHanvp/g4Do
dC0IRi8l/b2WUX/R4PmDpYbxMCHDhZ4gda6goKOgnystkMfnKhhouWvjpFT/oU/r
29FkKtCQaagkT+8IsODqAfOwVXM9gvPk6OuvM5ZfTHAEDqY5gTl478T4dLIXHe99
Ot+xjdxnOGVnLaxwEmW2S5mgqoUhv5MPQeIQ4okYrnDG251/qtPP76kBCs3/+gbO
2RGwgl3Gfql/e4fuyht0vvxeb6f+mC33fjGVP3Fi0x4RcnPEYgaQ42z+pcDzFwWc
7n8MPEAfCwVLMz6p6655DFdpGhO7QHI1vKRhU1jvkA8i39qfYwSeFtKB9Nsrgqdm
ONuGS+pSweBLZYFgl3VQHucKRxpC33yT5IMmsIfltfCLLHcQw42Z6NHR8d/7zPgZ
UazFJKFZhwayC0YUihY9MFtWpe8uekaFpeJgYDJR1ps6IhTJymU6KeDTR7eSTArT
j6By648GNplmcGerw3mZQ/vvbuAAAntVriqrA+6UOslGv4ekMgO6KPHdLdaODGQi
ZyeDSdplQgdVirntC02OGT6jqJK1SMvnI/ZFR2UjfJLaxmpAVrCxCebkSEGb9SsM
GBburIp+LI8NsZlKbaqfEEVE9vZ3vWjl4ZVU3O91P9nItTrYxeKCp7Qs/VW38Q8p
0PkRb/06uB1RA9R5HJYOWP+aA1hWzvOj9XC3i6am0j5cJdWcFM1XDpqeWojR6Wnl
W+LPLlh16ffrsbgUJ8DRQ+8Cf8JfT23Z0ApE4yaYnVk28wx3cmsvTSyjBiMY3uge
DUJKvlW2umGbLs0sZFmFPulJIJlT9q/ET0v/3UVZHv5/2Oj6vkBNw5Iv0ai13ng4
w+of8H9zbm4ykrTyYHLT7S4N+0D4e1w8/YIfF/8aPCi0wtQOh0htoPNPxpohxqWZ
t91cwKE6OwiSxykK8h5dJlBlSKkAOaGgZCns3ryXasFV/clX0HyZvNXRoR/62SPt
3lEyZ/eDklevq1yNuZl+zGQ0XOuOhDf+NhecEUbGLtKxdhpP3V3JNK4XH8TA0GJ7
XIxJlOVXsDA16SmWMC2MmJVWEeOtqmQkWXRT03IioxwbOb3XitrXMD7Qi3NjRb3z
dyoZqHmzdQ7STTBC3mMKUC6D5hEF3bGI/M0rHyILIJ9c9FLDgrkrVgtVIMus7E2r
y5drRN6k08u+ZniwXhxatMQz/q2/XvQfDpjGM05pKyWuLY2gYEVaJzY2W4t+JnYI
ILK8NY77/8GzsoY2rRmC8VUAxUzmlCkpDw2N1XH3LUamN1LYT2zR20NENkvhH6vV
gTDCe01haqrjKDcWC1xW+ZQLFwFcZ+FFzvwk0STgmFVakZ9O0/UixMjOE980JQxX
JAkp3CumVTIGmS0L0gnq8mroUh6GNIwfifMzqoswAWnGLAEDt18UsisXvJyBl4u4
vBJ4/IDod7SB6pGPO5SeP4/nWkviNEJbQmOUHkeBkdZc2VRDvAJCCtaFqKhP2K7q
zD9haKnEGOTjCXsXTnlaXpVdN/AfXUyNsUfM4qpBLv7JGu8ba+UJYqV3c3xTivjt
bzjU361tc4LXkXaQNiOJibE7JqMqszPGWQkSQxCOAkyKVwh/6G500F4U6S915qmZ
cAlbrlR6M/+hR2EkP1vvSJ/2kHb8ZEWVfdvXzgCIC15YlzL+drTS9Qb3yXaTgGpJ
KWXn4M3FvCqF8DSTlZASIEQLfzCBiNKHZKwqSMfVAnVvNZQvdycKQGJei1CDyLBJ
HTwGFmc/iCaRuyfsEFD0E5WP4RHppwuiWZ+Ik82zvJbqlwRP+RcVBkvrVXLLTxGe
lLLR4SaHogFTJle2fxXEROQq7RMXQHTKboaYnCN5neC2kbbaCqP7EMGTdPNahqWi
tQ4Mq1fUl7RfKKba/DAvOq0pfWkPXsR5O6QTlEfGFSJbTj2YmRw6pEtb1pGb1C3T
2jh1D2KWg7iDCJlb26ces6ub5wEE6N+c6XtMVlLSdnwQmTraG+5fIP7bb6ku5fbz
haku+NQDpL4q1pDGb7YZXGO/0Z0Qw3VEkW7t9olTnyeSyQx8lWQUpnVYt5miw5yA
laC3XT04NmSqvcOlzaGHgwm6rx2pA2DCA80ttegHJkwqxKhRg5zzfqa/fdvsZzy3
RQYO9pBzZC4785JjRQz2blj6AD/E5z6WzRJ7MD6pOhqGpSqTHcoc4l+KnsaDCqlL
Arg/5FG2v5shcVuZYOIPm1GEh/Ul3Oy6qSPJjZh7PDfqXZF9aon5Jrb3747w8/fB
atu4uPj2s+PW8Y2YO26R+TLrLcOx2K6Xb31uN5wjWCWk5WFSEZJbCiqaY4EWGx7d
20vsQX0gg5qHEviPGCFL0XfHGz+iFM9qZUOt4Ff4cOu9g42uBYsAT7IkUDmJgu3O
wkd95XupTcEOPRVqUT6t0VDkLNSbL5brGGw7BpR33Gk1jbtx0v+Q9mbOmwXg6B+c
xV0duElYiNtlDFxGqfUyXctVLSrZUMakugYL7lkar/gv7AeT/LxqOk5mXYZ/1QJn
tAXLvcNW4/xhIpA6Z9FD3xgTAI0HttX9OnhSp6N9MKaMDtZKiZjOGK3aGglHIIKw
G6Bwmi+iAxZEGv/m2V8hH9yGf0roAxtPfJInyIXrNKE2OS56eGiN77gf6iE5v0eJ
6c9XKQ82lABWl8T4FyEs81Hz9HOrontdipfg69vS0zqieBSpXYtkm7Ma0AoymvCt
GtSMpoVHrXkYa2jVSQEJv/GNfeieDb9qu9VIh+b3dJE0RQuE5JivKNLDBBVdkkgX
IAi00IUW6Eyxe5Opnq9vpGNtV7b52WfW450L8+6vwurfUBfRh642pkmUaVqUDg7J
rxkt+VrhIY4izPCZ+N5+KOtNiucyxYhBw8Yl/FcEY3hyv0GG8bQCl3iwvi1Bz+Xt
aCe0kSGAsz1EShGa/iJpj3xjPVpP3uUId5JJ0gqbiTXR9tpjwoVyIvAu9VSw3NHc
g+MuBpkdHJI9MpkZAJIyvX1AtFvcGhPwR0Bijqs2sQTXDdy9ELFAUZZ/K6kVsgml
zDviw+Vw+hB99AwfPeXVnMMdBDdUeefctLEFmF9Ofofg4JhzGkXKupSD7Bj3FsCC
XVcYBTD59rWUBpDIiSzDo/nVPxEOc6fKi1Ix+RRWqBOFZamfycDjhSFHXBje9jt/
DrIVVpyvqFIgEha0I+0UOI+ZX7OHd0ge/7sKU4Zcwp/yXpdkJhX73+8mOpDmVJjl
OgOEqi0gemWT7PeCxKZDKUnj5ItDQd+FEzfcJuvaHtRTyZvzS6tXi/sV8CgRlffe
75iH5CKa/rgjSLPOwvSDHihEmZgg9Oxwew/miTK4WR0ob7BHHzzmKiPeBTDcmUIk
VXMmG39g/wL2WNZ7zLDD0ftjcE4I7faj6TLDx0dEgt+Zo1aSfob1K1erQKBdOdWd
rINsVmpQWe0SucYUU7ZqoGBMh4dN6/mSGavRTjRaMOrbCLiIZwt1+XldLaK7iQmS
me2a5oVGPC8DmQvgpC5gIbyeSQgjXcKjvX0ltE7G90fjfIbodNNm2YPzzPKRB0LK
v8w1PAa2I2d0Pr3YSGT9aWSRe876wf/T/0LXbTsD4RmpkFqAOvgFTtb74paZNiYN
TjJ3iNsUIHNsB7yFvkTqKlNBTeYkwi2ltgV+zlm7hAR7swuBs+Wmhgn5jiK56D4b
BEjXw21qFDVRfwBtkjRcjKg5Mx9NZAQYEXeecPDn2YBD6wgYzO2Sfzl5Ee4fc0jk
JmxycE/NoqYWo3iqQDrc1rdv4rKwDs0qGxmvte4CrFuCQjGNmdbu1rNHv63uZoeu
qapfP+4muIoe46tyAtMM10sm3hEKo5AB5Ih4XcWYbm2BwsTdP0GF74+XCXm0dNCV
bTZ5z9ZuVtgbY6aP/TfJ/yR/lQeuqh1idT1wNGuxlpMC6jCKplTZfqFlb/upfSFp
ZI1gmn37Sl5hQc8dSCcshk+YEwGA6h77RQSfzcKrOD4Vb+9tIXwBzhpIgta+yF/W
uZqHpd6mKH32QeO6+7s8sA6XbVsAQMT6sUKQ3LAREEQEWnWAYb/pq8bm76Z7c9xY
xvGG6a7tjRmXbHJIPYFrNTzlaRKkP/UQH45CYFLy56Rm93G2sR9pSpcHmsRTaMSf
5BrHX+e+TfiRylHKAdYxnX6pBseVFe3Mu6mjylghhcaPT7nHq+BWzf5cRgzMsENT
qb3g3CrzclgI8i4Q2aqsc5LlagqYD989E1A5CQI+2JCuRzEQoOvct2EFeXPQtenj
4peTCXKHxBtgpFWJdDXPMnku2T0TGiunAnkKzZMXGDqmKIPyHO8AYgMrpAvuBThs
CUkS9ERXwk31OgOdvkhqb4FRMy9jWLrhY64inhessPRXvkxHENYmJlje3VS012JP
y20CZPPqdLCeI86k1YJkD2RKKiY7hRHg/Dk0M5HkooDyxIgMr9Tmrx7rg9lvIORC
rsB89CNvM2XfXiH8xoftXU5a4k9GIWCgVFhfe1eCoEJ1khrKjNH8OHCaVgi92lW0
pdynoNtvOP25m0d0vswxUY2CjoIb+scTN/L27UYqBGL2o9F6plBZ/g89+Zif58FG
g8dlHDYv9dIiedKiUM1wMX+oSvgjZ3vdyrdUSZJTjKikXRCei+uAJmtBeq1Tt/eW
Xbfp+Brruz1I/e8Eye0kynYgfGwS5k7Dk8OPSY1JxWHqd8W+aD207DXQrXf4/U3g
cs7CC/XRoNNVhn/zpda0hVRKDEXuV2wXdV7rHrm6u0HqkQ5GBcIyMz1Agosfx07k
73491wYEW0nkDrKvhGWyZ6bE+ezeGdzNQUgb85S+oAGIl1kw+VfnXZX/CiRvvEQr
iajEBKEGdSrL50hR/dL9aULSoULcOlpKBqqdr4TJSLgm0wLgXHDz5YyhCAbG8ifN
CgxaNnuPePE+B613+0kdJICCBe3QT+b+lXHrPQ4hKMmG2zCNdChW2jNjXsQxQq9U
0k2WTO9hzHJDS+T5fR3QDIcXRQNVsR8hhxI9kTP7xgjLoKIOilZcaQeFoFN5NIWe
x39s/H4p1LPm2V0EcaAD1WLSNwAZ8xVuu9qx5/W0tjtnQh1Bgt0KbRbD/HLm3kJ0
LkO1B+VjkZu6CWtECnxXvcwEgfvO+FpfDUjuCi3c+kDK7IBxk9mf6mDq7uDLUUNM
X9kE3/M9FOHkQlhj7o18TfxsNt8QFRc5wwV3uuJs6VbhssWRKB6wOROfWRNsvxU4
3Xp4b28qNlygXB7OVXoUdtwdW7mq69PDxTAvprStS91h2pXaN9i0CaOYTyltES82
ERTVoNdpE+azII5/VOZ9mob8Uw85fJcP1X4rP7f+DF8WgzIgev/zHINh07ZDIM2J
YPiUJULZ5L2Xdu33SGhkhuJS7R2fnjRC8Vv6SUbhAY6rN2f2EiZfWpeB696w1Ta7
GvPhOp51tUGgyAzrirRjLp+LtCXDFINXnysxYvtsvwzmJzC5LJq/8/+3KX9GiZPe
CHqdpPEzw7xmJZWmycbZpG/t2F79Mp4DUP26X/0CvJWTRSsCOe/vHO4ZqqDjAVtO
iX4h0pPmsWXljisIHeP2oHvKuJWb6z7ersuJz2qfjiF+3NKkU/veYjl6zf9MwNFg
jhmvI2utwIHC0nLrn64FH3tnjtWZlcCxIpT1cD+4criANZNxRB2cNrU5NT57cJnc
iFjC9nD05EP68rndYuZJfkdLDNiE4AqaInfKtk4eHUyqiDgsjN7V9k4nUcm/mSkB
We+Q3lW4rCKvOL3EYQxTBubU7IPcyVMgCehXYoJeJ/gMu6CsQqNj2lqp/+1ZzdJq
GzV0Hd0z33AXEo5CwDtj+MQJMIdn3HPH+BLQL7tDQESFV31VVRhrVRUDoGRnqjCs
Hz2hOuVN6FYRjz4WwaEp+t2rb0gVUveA60CvFH4/yt91KLWwiSkLvXFQP38urYX5
gPPRIwIpCnouSVT3JDjbhS/FLvXEHTqgeI/kuU23/L8HYGEFdkBKFlw94P4HPm/j
Mz0ALG80bcXc9mgJZfhtAp2Z/PdF8NuJdrTt9tvSVbv5YhP2RHskUI2/KWjXrjdm
Sfqw1n1MnvT317vqbULwtsP3UddRYKr1Be+JZMmWWF3DioOeXu1Zx875GtlOeBe4
xyb0GWWZZBhKOF6u4IdlPVakeX5RTEmba+xaxrx1ApxS4hZGBPqCkxk5TA0h0sNY
HvFkHuK3fA9J220QY0reRYmMcENo1vQqYI+yZd27jZNNPNFitQYrsXMwknznUqfG
GSuEX3oz7Rk9P/Xz/P6MVdRsLB++YEOXh1+K6/9D0MYLWPP2sFOCRz4zRF9hI6Fn
Eh/kNjR/d72OOqVsxvwl6s0KS5t3cJsPbX5m3CSPnFDAXgEbn2GuMO+tGLsbGmcR
9EtjLuy1Gq4a+M9t2OABd9+0+ggeKWkbBmedQv8m2XnsblYDWRRtqDR/86oVxqEu
FoHLPXHMP+EIqLzQbkGJt+P6O2Q6mIUzHDEfPmA93WVlIt6zlJ2XX3JLPvZiWwVU
H4QjkKP5pPUYQ8y0WViLZJd9CWg1FdqGxlM4VY9Ti+Yiat3BBw0mF4+Xx8bfBxRN
ULjGs+7ZRahtpEfGaMW5YIchgEMuBQhlQrpxQZJVDN8E+3AGYnb2NNApH+DT/nex
UYE62h1h0pEldpu24wZ92CfEecFCPVV5hs30pnPygPs8o2ak+PB4JgZTxcDnTNCL
xIIpkP9E7mqLDr0KniLl9S7iyLlHolzueF2royL72tozvwN9DR3O1POlUCj+zuhf
MHVDz44zq14NTJI/Nc8ApoLWHST2ZNfGeLpjwZwddcgpU2ElT2T+B+tHXhFNhkbX
C3ZcdeEGPdPOsvadITO02BDd7rIsjo1DP19JByYlQKOSYz30I6Ur9TeJ73SWU/9A
8mRWvENwkQm23oPgyAhqhFMLNUtHISavY2nRUZiZH1MAO69bUYX0AJyHGrQIZ0c8
FYY1kBfGJHNby1ofm4IIOgPJucvblcW/v6d24VajM8JNnno0c4GBLdrRvXzzk8Dv
zmq4GufzyunD1/AgTG6P3tmgFnEBI/pW3KbsDIKHKXUIRmuHuvxzmWszoHd6Qc8H
AZaC7ncxrZEFcbEzsZ8+qogmUK3eBaxx8/IqSbaYrP3/7jLk9J14MUtJvkm/Omo/
IF2Nedt/pMplcg0Z2lCYtXC9I6nJT0rpEYQfnt0tVa0moM06CuKGO/YG3FMAm6+g
yKvuZM1bNLTrZccgV3SLS+yajU9QuZjGV+9Li+us51l3MKZchgUEeZBu4ks+tTfL
VbMs3H8j/yBLzPtdL5m5cKLJ9cRUZUEffrx7aYE4Jd5BlbzdFjfxqGr94vtj6kb7
nG77DKV76E7qU7+OpL28uB4wFA+EqGbtkhHwMWl5EOfAMgv5Pl0jJPACIpWP7Dz2
JVc7jqmsd3GSfHjbCBkef3+4jU/pYuXfeQNbKFFJIeFba39sA+DG4SBpxCGWcFxM
6rwfSUFR19qqJk0QYeVRn/4VMjGLWeezQFRZtfRgiyx4/AwSiyYl9w8dVj3MOAEv
xXHkqPPu5tRMHG9FM0uXMHn0SJ/RLnwbbG5LtB6NeJSxfK3VIxALzdRnbLX0lLB+
TH3/CxvKNIcGjV3ly777NAkff0AU7mlXHBly+ctXbX/LgeQqb6Inqciy1wZFccG5
jyHSx+nZrDYqiSHh/Ei8VACxTVtx+Mirc7ubHyDMal4FCUEQ71a4xp9ozkmFtkBt
5UGdI2Yd3qpgvzTiYs4UChXJfamWMrnORZF8iRr19RUo9F8/+UX6sr1URP5PGTSN
xUN1S9OHubbz2rc8nPBRUDff8xdIZQJVzdpRnNknX1S5Wd5dBoF+QXK0KCTtMejB
Aa7FzkowlyB41pSTEof8OViDRUH8rT+VKfzM2dCS9S1WPpM0WoHZEpgzFejN8WRT
dPbL+gD0j5kIWCErf6HosAjhxLoIotzPly8sN45aQIGJvahgZYBp+U1C8Iwz2BmR
EzC5DGNFQsFk3rivWZkveRpQtzyAOt3t9gGlWTTnEmJBBYmWimtcDCVXMQlH/PjF
y4si19GYwkI11yXKNHyLLd8XkLOTpzlIvrSJKnJIbcGGw6VsDuV4xzmUkeLxNr0v
w9bzxYR4f5V09cDbMHfP6a2KVe0nWPutt8l+1p6QcsUq0zMynMkkAZfezqtr28bA
VrTqlrTCxLdJHvkE1g9j26K1mHNaIR/gDfURLD9qHgkKbFmCmucQp9L/BD3a0i4t
RG7LM1mHygbrEN/OXrVUFMQK0csPrQr/O5Lgld+Vr80Bw4k6tdmnA1eedFAL8+ui
qjdDN7JVBrDo6iBLPPPTNhwcV5KTXqDk40D4JXSPja4qOwquCu1ns3zH3F5g5v0k
Vq10QutNGCL5EsGyVyPq6io9XrjvmRgCABbVemosgotRGLVQu5hFTa7lTQAvz37Z
jgBT0JmUPHcAnzT2Fp37v8K4yI4tQJmBo5tONpLuxcvxPCPPHjSqo3Yfyu2g2Ybl
S3osjFGvs8WU8OCbEsEVNLgL9sCDJsNeXq3aHkHHos7j5GWUXxwuA5R7f8uotrsR
081ZNiEaam/1vEu2vjAgGj6uKrKDTJ+ifS10CUc3sXxR6vL00VkS7Cr9ck48Hx8i
SOLjqAGvxaBY4LDBOyCyBsJ039JQo5r3ZHCVMGxgFwEN6lLcVRWIxG0VgGjJ2Jlb
IIDD2JWzeCiR3DhCvuxk4+nEGeIe8jc1ZgtySTSG8Cf6rd5b8mAk3Ye54nN8lk+M
hwDatVraSOVfAy2o15hsVZtxK3g/9Zn4FsZBvdg2sH0e2usgr68pokm4YyRaSh9P
UQwxAmElAi1DaDxJN5qVsYkM+2RCCjEasYp2arvxQ/giR7tj2xybPr41Za6T6pMM
qoqXR+YHhKus5XmCP9stoAHRX/2aL/sw7P5pN/xJDzKRaaX+X1eCyqJUVbDZOR1R
bm1ynDK6hu2zgTOOPaB085JEnLXpvoYrBN+ENZy2amnXApQX6lQo8hpV/haQ6WHm
/dy9EsGtSaw89JGaiP9v+tO9BiMPRpj1krqBAOfRk7xjdWkdCNsBfDiMU8ZYbwuh
2AnXCIwo+f8UdDbie1UYMxf5voa1ZY8qPSbGnJs41qmAbO8bSvnG2Ql6exGMzrY1
iAlI9Jv2e0GVtg+xrzepMx6CbuR0A7CgZAecH1j9jh3CnJjjRFU+D/BPG5MvjOek
o6BTyP3D8Tuk9aEC0lvaHe801GYlj+VGmCg3hrKmnKHlQvlsNqPvTTTmIqQx3hEW
4BbGTRwH9uMuhIYOIoBgCo1S9D0P1mPHafRsyHRIgZCKaPtE0C1bu211WYDIjww6
MweW44Oo/8It9tbuC0BlmDZGFb2sDfeR+wm44WqqkF3Vov4KkJ+F6JZdxyW0njJG
Kgjlq+CfKNYnCztB3GKtQpZm5FzSyyWKLeFw+h+yTqcYBmIwvi9OodFl/2NacGtT
G1c4IMtGBlUa0S+uTCXj7mvv2sQ/V+awai+vUOGOx2oopfCh/kQP9IbMN9J1RqpU
PIceMfGJ2kv8SVMQfEHPVYn00Lu4LQG0OeVIY1wsbogCD21tETC+bFgvHcYqOS6W
yay1bkOguwgoa6rH163xJTBBxzEyZOO9p43+kurchG+/HaAmZTwBUWlFWd3GcIJS
0BdYN1OzPzuSBaMw0uxfjrEH7Fx/p2dwN5cyxwlrNk4k0+JaxU8q1wsOqr+sjHPT
VJ3hspM9/ZKp61x4ZPviFOth+LxlEsUO6Bkg2PLU+n9r1STCK5Z2RDi3cFBE7cy0
HOHynT4RhC8n7ca5pb+abuIqZ041M4TVWULKpx9j5pxlPZfcXnq31ze/Avsa3U+b
4pMHw3teKj/4Ss+Z4gu5mcyS6OiQSaxm4z/6xF5A0B+PvN6D7jRUc+r6TEjevWC9
sv+7JIUIXKhlBPcZFotFHcSX6makGu+CFjcQBbKDyePB3M3isbFxCcdU4AgDdOTp
SbIYq9JC7PRy433hxlAWcD+SOqjA+kGz8Z8meMCie71daMpltKjLsLdULD9gJ7YV
5QyZBUxeE8XsEknYO+OPmpsyOy08lz1q1crvBKpmer91oN2Lkktg+FDREvsk06pW
aTm2jd+yetNB8qW9TRL+hHJu6f4HVMAbLai0VuRx0dIk4vkpc/Ri42/PA71mRhR2
5JxiekhHxNaKa6YzyfiyXOJLwqG1fxDOnUmnsH37wWSBVRO0/pSOLPl7Y8/6S7fp
/N6oY3ro/F7llNuTkaRZAU1ad6Jk60g0XeRuQXAmAsJBr7UJsDzEcoqAoDiJ69EO
EUzZh6C4Nz0b3+VBK5LnAuK+6B7M9aRMntUWFpL56/shxryQr3G5DSQCH/hkimbd
fnXH7i86UYivXZtXazfTKhCUK+P9kg3DwCUwPh47MqCKvIlUD08JI4zSqvajW7WE
8EX7rxstB9cRr0h7oSHpDcXnZFjiekY28I0MIFA6vI+R8BhKWpxPaLgl74v9ojQO
FRm+okd9IVuSA9jZTBTHd3RQUm3+aZCbDPai1pKQZurJa3EtLzJjiq1uI2dXTRuJ
am5JTAzCcRPDIrs1Lri9sp643b69B9FJVyHmbqkUsrg13YGN/TWduj/piZKESElr
/bQhlDijCtXuE/WgBwrwJV4hGK36kqMfO/BsH8S08XuVPaVpVLcVCVaDWwci/P3q
vxx65pNsOJ+D0PLeae1AxR6kYge5pyEg4pTpMk5TYpWGMTzZB+Wt8cvaNWm1BLEG
zVaZPS46smbgAa1M1Svti8575quGfifMz/D7jI27LP0KG8e4x7V8FsR1IZNMqBXa
HOa4hBb8qwGNohgF4WnoounEAAoB2JHxau02XbuSRxA6gjxIioFVAnn/Fs8aFFUq
6e1QtGPkLYv2Jq3SfhxinRc7nSjZ8JI9ZJ6ODLo7bnMFJPUGqJWGOAFVKYaYLqrN
E5VAUs1xoMyCudWvEu/sDEhMM1D69TQLl7bwGvYdMF6tlGt4XWJj5QZvkhRuQ4A5
ITYQ5jHAhR4tyqXpAJGOHWTakKu66O/Zpv/pQsBVrR0pOmmeNJs0E6x8wI7wXwMT
8YqGIZbX+98vuIYcbqulHel+YG4OuUUPb2C/GQeBSQip3rypXgAsR6Vnmk7ja3dp
fJs3DLQxfG5VG0pQGzV9zQKrEhn02RAm1SkGYSC6DKz9xBUG2Vy6rwBdSF/dfink
bMRpLpeoi/1GwecZdFNMoOPdxOrIEhuO+vnTb2Km1gkSrYae/67FhaLtM3yFPaLY
M1uUH6RwRn4qzoo4tspdk8fi9+ryJfhu66T8rlAfgU0St01Yp5K05GooCRebWXVk
jdzq/9yjTds2XxSD2itKENrJe2epYECUPVcyuyucaqdreqwdKxD522DYQ1mBx99Y
VC3icB6svtW+kpMSnj1U/YeZeE3lKXQje6ZNtHd5whjrmA+08dOAxI9fOXJau2m7
u5AP+2gnzqJ7xnC9LMFrBxb2uqMnQ4qO/t3EiZSr6lcQ+OOcJcxTfiy7DiXY4oRG
nkehJv9VdgDuunRnz6b/ZXF9ndm4I0N5gfMnAiP6xuiX1a4ahih+rcOcrgnsl80z
7v4SPj/groPwNVGnzj4bx4IKdrUrYUu0yQBSbJwUkxOVLDelgT9ylfM2FmtTPfsx
tdghNLwZB6b00PI/AicA4Vv6ajxwRxUce4wUgeQjkYOTNFLNfPO6gLA2RKIqAHaS
FH4+1bIhHClIk0TIYvZ8uKYF828HNqlqy4FGYljc2ZHrjQ9rjErFFwWB0JDMccYh
nKVaIG/MvSDB/WdUwQkuTzdeoCTVdHSLJTxrAZ+8uQ9t7aflC9BKUBvmZA2cEJ36
7WT/T8jZMbdlheUZsUgUXERaAimkFEKcXBSRjSoHIb8Js1a9MY11yDjAVp+i1AxP
cZzY0HwS7O+0aVwqXBPKhDfhvJ6Z6GNdna+qe8JAdNXkRLAMeb9peS4KicZZUHsn
qJhGORlp/w6u5ivN4afpiyNO14YAXMvcBF4RFtFFM+vHU1H9ZIhj68tYJsSq46e7
yK33Vkfdwgw6DIltQcRLyKM5XZalQqCWVvt+i3z7f4XDQYkqNdQ/nRioBF0rYl+8
YdReXVVZMrXI13szM87uTXFTLb74Yk4zPUW53vPDO8tx0tvlmAQVOFKire1+qpzE
Yw/jLfYrDy/qzNFCgGNQ+rVtzuySXaiNUM8mjgZrg+QboOnmplueWDw5EoRoMmx/
4otAo9RBDI8kYS3WRONSc27KOFX8Zr5+0n+l0WAwIY64K4tz0DmAQ7YONJJ9r2XQ
yAzxQxI+083E7eaIBL8RAdRYguibkKVW9zR9tFZIJVRKTxKFm8x5r2Z1gG8a3Z7v
lAhwoeV4qu3fU0ckRNB/Y8MA68SfKUhxb7MfBcxi+ceW5aE3NXGvP1g79xxqHZQK
mMTjy+a6M4B2Ku07zvxurYdOF7hUTfkyTL5I7dpGhUGBKR8/dsCvVPli6EsShsJu
yq7601EqOm9L/Mc1vJc/x8uaTHtF0cQ7h0EvSxsjnd9nk+s6LUX2Z5hqOME3GAje
kJlg8ImykLMDegj33fReTr/J0lFeX2G4GGNUVequH0ejzkYeX3ZpCHqWr5wV6wCu
Gkxpmqe3PAQmKoS5uYiC5MSEV7suDgZW7dktz4alsZkZHCvJyMEAnA0gVIZm0F4d
C5dTKnVPLd9Nf6/iDqAZpAacDnVROPmNsk+3O7zULHYmC4Oxz3bkLqbmb1wRLJ2O
2khzvnXjyQVT60cSF6MuuX4u4ys8UiFmOn/m8ZG48pbm59f+a+kO54wrOp6oCuYt
fA+Jb/kOaaCMwvN5UlFTiLIAwWj9XDrSVD1Tq4OZt87g6gMddu44Vlds9mipEDvm
sRoE42WiJ1+syILaQS64Shb/GjorxVbrLOK7+FoH3+bgPf4o41/LAIGOi1no19Nn
Gy4/2Rs81BzHmrKobB6GRDYjYjleyBwRLAHcmRQMcMcDkMEFaBD9i9UK70O21bHf
xfcmuGLXjcicoX8Hcm3kGpFzEUWXM931i4x4uhD+Ub07qP1QaXnuqE0zju+I9Fg7
Ss+Cx/KJ411w0mLgxxusJNqpmeP0vpgX1dSEA/+TD0G70Rx0qZDGPER6mE3oS/51
9AFgdvEduAxZ5gHk9iuScevXFrldPLh4zD/zCQjOgvcAmfopgNBfwd0tCv2FU/29
PUy+ZVkQgus9o4vxFsgz6gewryLvRZ/Jo2sG6jIc7PpMEMkwfqGqXcbKTIRV1sIw
kyqsgXepUsY8yPmpnSUernL6U0HJW5Szx3dvvxClegUaDSI+m/4+z7slTjINZNCu
v3WITGgnua1SIiiFdk67W5Hrinem7lE2ubETkOwobXs5f0AmUkArhxqDftEDT62g
Aa4hTC25SMYR3JkcwD/kXSe1pb8B3W2r9dnli97i7GuGI642UGGZNJhQLelktOP6
FVgb/Tb3Hld+6IjQTAlDLJVoP0ar5E/gqF8LhFtUgCbCXr1GTPQ7VnGlDNkh+838
H17Hqn94XMFyb+NRMHmfZK8iGUN+vlt2wtYIBHleRdzOEkYW1kYER79lTusFoQpH
w31rNS5WPH1uEdJ/659nSLWedEwx04mmyJbvXzJyYB5MNVW8UMxn+DnySwsZWa4i
UT/8rLbzQi4VMsk0oYwtG+CXr3vKjeAdS2kWSVJS7t3rx/RjdG0FdwZi4Vwqz3eU
sR+fdYUktHUjwYCT3W9tsxak9eCop7hh+FMJjTsBIN13b7OESNbXq9/+uEJnpnyo
/831i4bxNNKBL12cpV9BJJcWCMwFoPKCwUqvCPIPtmS4LdZFBYHwfi28DZ4SKW5E
se7+ADH9wQxgNKWmIDxWXCnl92wDOHf7GVobKKbiD5Y4L5DDpt7eG5kAZs0wwhqf
0yyrXUT3T+eniZ2IBNncu6DxQ+amlknDG6or8NqfO6FJTBMi1NO8K6R0al2FF3U2
ZrTGqPMHctT6HhvLlaFBSwvzvzBFQ8t6G079Vi3afTiedEAB3BDP/aABr2UL7rtw
l0m0zNLWzY/b7ezzoQgJow5/UkZtC9C54fjJ+ztG8BlOSnps8spqab7hqpc9RlWz
otc+SVCCQPYx0nPc1q5P4i9ytWzq1dXHt+2Ur/M96Zq54eqGjP7qGchC2XWgmD8G
wczwY38+UHX2CciI2CyfG3r3YJKKE+fWuCVSIClltHoOGYU9a6262TOs/qJfLA5X
8TcpNyWjbFJzobWzD7aoLdbDGzQ6VLjl9qMJmxwtCJQRx2mYNIl9ekxW8/sRvbtu
Hx4uHyG5N2/xlIDSTPkZXLl1dEoAk8GNDvD7pG/UteP92K8Nf5Z0jwO5Mt04Qwhx
wVYjMCa0JS2Ah1B6aofcsYeWlAOFPxJcbFKi1/NwvpivupwbB07GX7Zi2oEeBILy
2FVtNp2muW7ZF9+vOLoPCSyNiaPSkRUbqo3VU9+0w3MySUi8xTnU9W+yKu52yoEm
L1UIdmopemWxHTjdWkh6KL/4ScX79CfJ+hDbd6DQuPLkpRxm8n6yZQw7BTRhU0xQ
uBRZwfVyV6RiiO58K0D+9bJywv0XDhdidwcRmNqs8kB88zgEFf8EF6bimWR5l2uX
rj7FbAGfeE8rTOQBMCtbYbN2BuqZGEOE4f+6GU4kFD+tDpkJp/fIVD1pj3XXiiPP
t0lqcQmPdivySJSwMPx1Y1LHb8nMWyg06W2lRPV7XmuvfrMPLSUMjL5G2ory/yGg
WCH6Kl6IcZiajhVrns39TfHx4iYltp/pt9IBMORzoN7puTRPoXWDtJN7ZPKJZb+R
qMxt3d7Bfvnv8r+/VXf2IVbAOw5afhMBXTzUTOek0Mvzchtkyfj3CkU6a9XjYg7M
sbTNhbx1HmkaacERZGVKUNiSr2xijPOMyy4RAadB7gA2BK/0A+oHt2ecc5WIuqBu
keOlyTDyFyVy9Sqa0sCv+mQwaGdQ2bUXUPRbpu0mHaNUpXMh7DilE4O1utm830DJ
bx5/4yx4lwuY5U21+GXVRJRYvnsTR2VUqJ8Css90BeEpPyiif3TO/9tVuyL7HyJa
dNCQnQEbcqlzosJZJWzxc8wumDtv4Y7aydJNIazMjaNF5T7KHcIhG/0A2Jequx4v
q99hYfGvqwvScYGZrRdo/VlEsgTC1Az+Xrl1oZ7zD64Cttedt0GSgV57bE7ZRjcn
WUIopTyk1kUYYNrtnmh/7Hqj/Fp9o0a7XmhmVeERowYYQx5CYnqfBDcrYntDm+UL
tipk8zXTUd918vnUq+hR5NHGzeI2jxbjoitoj5SD4CGkxv4jfSp14hZMpjc4ITF9
B0Ecc12SKZ2Hbv56/HOHckQB06naKV6RiP9SjxCtospipXdjgB2UERJMQGfBJ/sE
zSzSGyodVxgl/JdIedmu6FuvIlY0HMH4n7uLJSMmuj1HM5TQBJxXa8s20icFrCQo
2+pGpsJ9+MAhWiB11m1NxW9Xnnx/xGfhHkvPvnEJdhXnwVst3i8rLPTgFoj4TC2O
v5+40KBIf/d26ot6zuDdhp1uG5UQ/VR33kP5rk58rGKM7Eh4jdlVtBjtNkiivhti
ZbNA1ix2GhCt6pL0YSE6i7yFO9VimdqmUAokwc5bG/3ZtXiRgvr0J3GL0Lmh55Xe
4brGOI7R3QLbTdvkjRcN+qda+LOIHkXhq/vs2dpOpGo3SrvCvhvvBv641M9VPQr9
J75s5eLpTi43pwNJkOdbfk85XZ+s++DxowAiQuf0hdCOrO0fMh2/7eSDYG0aJH5I
LIJVWOGG3GZEKxv/fg9r0volN1RVvxLV/bKnWRfaiVm2pcZ4xtTOWXGu+pvCrKSe
06DeqRj2TZGlWgvLqHi6KhfZsHQHrctAbLa0gjeG6U7Fh1gibhRl3ntEUjuPYgwa
h/9Bfe2QO78V53Ul4R3U1b1YSFHBFiLQuD5Ozn9yOj2GHho4MroMzVTWsK8Yc32L
F51kboiNbgCIMaHShSb8pJJlhOB1KRy35M0lOs4rg70bXjH8jmi2T9fU3zrE8YL1
ajyjemkv/3dHOUFbQGmWoe86QKOTXUQvAxfxbgCXAonYqBbiHXDvGoK6RIoeopB0
GEGjy3qz9K2gQrbw13HZZy4/5ALDdxEZdoh0E5nrOH55LYV5CJxcsVzaIXyCaxEv
5jC1SPJ2QW2gM00V+MXPJjIfeX+hO8hSbAFUYEh/SkP8xMtzO+nT+1aVYKTII02q
Ks+S8T01sZL3mMJFtcD83iTwSWJm3yO0CII4J3L9x0YfhRxynIJykiuJt4vsD1rP
tywMHnvsdYvUak8NeDR36DX3rYJkF3IOxIxtoJey04/JQy6bVlSsreDNsxxfx/nh
rOYKd8647lPTlk7HJtgnKJimmMXE7DNJCA++xwrDsQxd2olvWEIM1TyPC4dFon0N
jcjVwFuoiGjBifRicISlEgWdbKibPYyBVU8zsMV8Rr5OEbE8uDRd/gG4nmtHwseW
H1F7XVlgM54iQl/twWt71PaHBWCaA/Y5/FUfHkBG+N/jT5rjC60EBgDECyhKdcri
/09qN7jBJvHvknBlyEzFTElg1+VI4C6D01NTu4hXTbtKgMOJm3N5yiG1Ej81YbC6
UdlyvfnCNzoEWmmgoVjuihbAbu7Q+GXM7tbFUH23RpKpoA1ulNegz+nZ1Yr8CN5Z
j9rNkiJxwFdlzToAETPWwtaw+/16VC4GDPyPDiKLS/d+rrkWawPPQTPoVu2Zdl6H
1xk1aUXFJa4OnP6+pB1s1OwLK7bn4uRolzocwx2iBrEV6jMrEqPvEdOR2OmpXYiX
Iifd7igGxcA4VP8/fnhmB9m6fMVLkxmJu/AUeNnPlGx/KNDiixo6PFLnKsTDQQYe
hbGABRYrB3kVggeU07/yBspqlEw6tgxT7qw84rsWW+G/mW2Ypi0UbxnVgSU960k4
grveqNYfYlocAUFiDKiMpBPY6OS5TnYFnQ0SiAGSpZ1trhciFnSMibFj9ghmAdcm
v5d3cXqvtay6bPJr43s3RAU17NAskhA7Z8xgp5UdOc1V0sGHGi9ERCDlJEtAz6ok
+sbZ6CF+1Kfl2fzkYHnJz1ZAeqjtR7pBFW8ahIwSltemXUOi+S+vPhJnjFlbw2Fx
nIsZSFWbDzBlcolk5yQ9kjwQFvi5fSmbmg4Xdyic0FeBvdZeWFf4xokRG5+KKLhg
b396bYTO7ll0CwnsODJ+hVUQ4w0W3jnMZzWr1jBWxWFdotMTrUUqn6/MjcVaJWKT
9RjW8RYmZ7j5qFc1AapXTfS3m0XD5F1YXdu/nit9VnU1FMdf0iCqPG8kuAnFpYfy
6LxqlmlV2DGHyeweRzcQEiscA6PS7TfRKzqzBRHAbICLlgiCQ7PXz2Yg+CIGW3Ip
0IAYy1nUTayT2GYnCLekeM0nfjMKGkk7LdKWWrcTULPj/p+iV1gvOkIPayhMe2GX
52rgOqfLlqMOZYyYtNyJzeXde7UJNvq1csTuKwBW4ALrybKcjcdt++nm4LZCOoDI
bRNfXsPu64hy3wceK9jNzWv3TtXFuxYyhJm85Gr14378iVWiFlJHn31lyHl0fBpl
PDov3qUEBT4QpeprcrMHa6qCQqo/dgaavuzcXnf0HnPgmJhVokzjM973q/gVeWcR
nGNet+zP8Nihgfexo1c5h+c0W5Col9Wdd1axfZemqM3dMXcfvOPG3QP8v8OX5gko
goeqIpJZEbOc4nd3mhxT0rjXf6Nikdhmw+M24HDBmjkjL0mI9B2Of63p4sN+Utpu
j0aVSLuEWTYJw13yyWSJOhFoaTMxhXXZIK5yDHWU0K6v+KE+dOeOzRaAPozKSk3W
U0El8NMImWB9nrpwK89VP+vQKDfsL1FOfZw4zSO69SYCo6uInFX1HxzzEKCVsDc/
rSlwu9Ly3Cy/jdNwoz39EL2APupOnsyCEU6Q+f3nLfloGqrO0sCU78oI8iV6KhyY
C/AtJZzFHj4QKoEOtL3j5PBOYtkiLLJLoZwvGIucHoSsoIsU96EVv0NuzY3W2F+1
5el2gf+RwhgNQsEyNz/hsjnbsEvY8WKinBJ+wKpkIUr8RVF5xhSi/vNQLYFTBo7X
HIzyhxj0tw1EX9eKDMc03MO4TvD17wUAJellEQa53IFj2iKf01tTY1X95k9N2ajh
xyY4z16jOJR/UOMHANQOk91vVOzevmOJ8BWem5Sm4G1Q9p4R5HXy7uiYfJKhiGda
5NexE/aTnkTihmE8aXIeBfZGR0ShQ2tfyRSOYUJr9SPgMr53cb2TzQZ8nfXUzYMD
szQPDBPKccP37Alyv2/shKt5jRv1iW9kfn4UBXpUQMb8U8kVtYcFGrr1dDnAgL42
Qk4BdBMfy3CwNHfLf8CON7YYM4gAsUtPRax9YwgMc0pEeYz7gTvzewMs/1x8jQnl
wqXD/DzjEdEY4+yhJVHcjIASMRiAmoBjBsOSh2LtraMLHzmrDYE8Ay9HBpXHT2p/
M2d5ELnX5UFduRqdiSGv9t06iKFcCk8OzBI8aOzS2o9aRRgSPOxgtd0CeOR3YIQ4
f70FgR/SVSk/tGzmi1dmhqURyCYxrJXkZGsGELLWIKTRu1K63wlBjJmalfPoG+2A
PUHmg+7vGx6nZEZZR5vor4phXJ8wfx3rqdVENrW2P/A65BxruDMMP1wPmyMABUZu
PkmRif7PFFsahi7OL3+Z+IuocP7pnkGJ+XwNId4xQ5Q+u38rkqiJGqU+DkMLX2pS
ouaB3umEbQV/c77aGDwtSBsQiTaIgaixU9TFCn0BPSWGWPBk8sxjXk+G04g8j9EG
GSgxNsA6xhefHl3thP7oduN2fXeWadr7j7XJhJePu1KC2xTW9iPaZ+8qSb6O/Q/M
6aXPiwkg9iEYkyH78yarWhYPqUX4j+dhQlQPUJk/m42OLQEQhISA4WtJVAF0KaPL
hgNN6jFCpNuhI4b6Sb+8j4t7mFJzbZ9A0gV/cgAU144Z0Gmx8hbnA8GoSyBiP2Za
o1aF5kmqk2d05MvRv4gDJ712itxkNWk2HwDExv9QrHyyYLAGE797K6zUYJZugoH2
8naz6nWuVxf97C6glCmN8Lxu0ka7V8PfLUNcFt546W8JwODtgN6dXnToiT037lxc
5aRTfHkK3yqgoDZgkfTTSu6cxABBdlMAy33otBqELWOXm+8o99A6ip624Bmpdcuj
VOVC33p2NUgN8J1yauvNRB1Jbtcm80fqEbOubVVU9IJso8PXyLOuVwCUZgmr+tgS
U46zYnNpf8oRXOtYLmG7O7FNdFQmoLa4ochTO2MASciLxWKFG5UNo8mAwhuJyXzE
cQ43jx5hnFaDAvt9+jUWrMY3wCi6IScYyPcc/Uu3krsKj09NaLLKR0D2TX0w7aRF
imG+Aw2wofXx+Y+vmtV50RzFJyOzMPcznrJYR8iP1W5vzlvfDFjCfTAcR42JDV6A
N/l6eMtP5/HqhBQduUCcwgCv3oyIudISO7pqoqx00DQE/BTxKDkr6IDUeRUGrK5n
Nroi8R2q8OB89xtxnK1IDtMUELpTkAWf8XISrRbd6p+Me/oXNN456ZzOVlZF7A00
JmQXzMEVkHZ02OPq41TWbnsjqX2y5Nqbj4cWNtPpIBg4GtsIcecChmWnhRapK894
zsARzAZruuic0KfMRtr7xeyABxnj6BLSy/g4lHeXysWaLzGQ97vUs8w2yItviBhV
vOlUkRBEein67hhUuYmhubhnuYHNcVe+dJK1xJdvSrK1tF5LxsFOHzHjlO2GMhrB
6UtasdPnMLlBWhk7AWiE+seGkz2RfCkMdpaiL9nYkJPXW4HRFPYxg001lejIeD+L
DC/pEdigl3ih05CpEGCE8KhdALixHDfHtGW3KNuvC3+HmcDOSs1zK6kA96olaL/c
cf5o6JOkf5QXLqXVZYrIIhrfhdFc1DL2svYNDRJdCrnoa35mHeXxnHc+Utf4Z1d0
8CrF2iJpsyUAWsxzY1aTgCOULHQnLEH1WA1+tR6r435l3773r7+g0184ZrCdWrQ+
ceugdiJg7XgYzV5h+32DkY4ugFeh46bKCXlPjWs57uMz9O1zioK/VJZIdhh26acR
ArsxrEI0Vfn6vn0ZP7rvP47IC6qCF55BltcXSxAckkPOkOsNmsiERQ3e6/r7qyR4
Y/UwryLinLPMG2pxM65cfBMKDpAXNEcU5pRSXp3vd9ARYAQA4SjY2fn+7o0ZfNNf
OM/Z6DMkZe+IDan2K/iqXy+JsssLVKqsI3Sw3JDv+u2nG8sm4vf8S7xBZ8UTHCu1
ERuTLTKxet9OjdAPzZv6dri1BHdoXTYa7olf1GWQrxfQefkQfxpK/14aO3Hwftmf
3VOQkpKhXkodHgPC39l0A/1ol75jXXf6FldK7DDIwt7iPUpv97stzvUu6Ybi88db
0ZDQ267VMTWqcv5kdv0XwlEPadKXJv56ME2J8JPwk1HMCpSO8rEDg7J7b60HbVoF
XytuECxOdOLBP8K6k5WV0jG45TuUJKLepmCSgeEKB1cPjMb3Z3ZiNPzz99sKLyAX
EasSx7U6idweXD0Gumk0FriqRPup+FqZqsgqdzclyJMuEU2//ry/13NCK/2LBaXG
IhnZx9+ezbEGx21PSOqIFX7X1ybqWMOiyeFdUiHh1TnsMCbsaAyDmFth4xgyhlZe
bxlW2Or5TjJ+7cusQYSGi2d3Wdf/HuKFKrja3t7DPlf9J2TRnueLT58rjilQNAQE
4Q0GWDA4Uhff0n6buCuDFghRvEnHOOjjioXXwwNLPmqSZAJBoB44RmwXLmU8BTDM
bkdh2bEnBclXLikEbD/5EbZOoM93mOQdDGPRLoiJWJJT9w/RxYxLfmq7hK4+ZvqZ
zWVplkMc4eatx1ghVTZWmZad2K1ONGxgZ5FeRm9INL9/vpzeBAMyQflvTitfaETC
6BQzsq8R/e5iS20i9bBny2vGZ+gEVE2iDwSCdvOOK8I+zc5pFiTCkW9n+ABjgE+4
7FmQUdcU8Uy0q1n8DdjwPBbdx3cQepsMuiAb2elfHI66y+skvcp5EXSiibPgZP4S
iZlBvPcrouTTwexrF/Wli1HZvv3m9CZfFQMDAP5nbJIySVcAOrvQDktvclfJtndr
llPYIrM1m0yBTs5NP4RwaP05fNeympf8Y6x27ptwDT1AL2MCm+pNgK96IgUyEjyg
OreNyq94GXsAR3yr8s9fZDgcRek1rfKvhJscrEZlHDJlgJqG2Qmez4MEgJ7G2euO
wnSTXlV6ynbOsudzvMLzKvvUXVx+R2MX/kaAr/PcPpseesFPfg+jQpHTwYQG9KOf
OLszRktWLHqtXlF15sKr6iVAbmJv7pxpEW/fDSeULgOjefgqFrQYmoPOn7ZPxgZv
YauDpoZjAz1EuyYeYcNJxqVAkEi3Ej/HWasiqlt8vzpScKCxCnMLlTZE07sXAa2i
z/Uzs5ELrTPxNDwMeqXX1V+7dsWU5r359ttEtu9WxQ/FDJZy95CLRZg9x0sSOgWh
oqWyCs+O0zMR3RNrIYnAP67p5fDz27GSm2nXtJZaaGenulkiuhYH0PsK7/2W3Y9S
7FQnVFFjGXbejmlTfy9PrNBzvqbwWGSo8LXA6OijBKT33vqU3yniCiYYIuGweV+U
UBb5X40nMnEsl69jJ4NitUkXMwnH1N6nADLaXmnA/JcBr7Mrgm0vdmyEeR4CaBps
rqlOJK4aURorsG6gHk2hS4YDDtlZR1o2LW5A4LtYKxjhNrJ+sy1T0RMRnw1A0c2+
O75L0y43wFRgewz458l+pvsYSxycvrnOZxeDom0zbN420TnD4n/Dmv4UGdQ20N3U
ZgN3bo+zsaFF1TinthZcO7b9fXReXlCeBcC7sKSDgBaPxFovT8OCU7MyPwoQP0An
H0+lbibi/JeQvveMe7Kjtb9Q07V6iPwK8WagTwaDQDha8YBo4aINU1C5ZwNRF+Y8
YLR/hR3AtANlv2lqb+2i+1iTb4nT4gJldbEgIQ5ZiB9We7+4XBvokWQly006089g
j86RyTUkFxEaE9nAVpwX8yPXCNcZFJFgFot9Ei3/+6bB7pEJGWNLg65ODSraZGbq
FgGTR2r0dw2ql4+8CfNEXF70OQGvpKPJ8MUBJLXOue5eu/jd4RcTrvasjtJALJ4R
I5Rp1h8nVNP1CEsM9/vy3O/V8Fr3AT6Qk6uXNlE3YOUiCDv2BLX2Y/SyIkxKFh9v
FkHeYa01bl1JTAhgmjL5/JNDmXN0oPtdRC2CQuW1vpiMoQ5qAK6ZVvFzEgtawWeP
0guYaGgRYkf75hrUYf27O5K7ag+4Pxy4CmkVBaI7ewkozSwDjwwme0pCuMo40hvR
a42NlR81Go71uQzcoBuYp3BSBRZElxe2h0YexJak5x02iUYIEpV12hS7UrzzXkGj
9HJb4YB4gLW/AgFs0IXpayGpvRpBLlAvuLRlEDAcCt94knA6HK0e3x9xbjKLEVS/
iJ5rgh0Etoyq06tFMhi5WK4Qoqlz1RkbdLzbX0t2NCSnxaQ6Hh3n781hzS80+yXo
5A3yH5z5D+iGZ30GCFZT1P0DlDJV3QCRKc1Rh9+IhhGKGizl6Q0rHI5DRzzmELiT
r/2R+CCi+JWv4gAvzp4l5mAt8eR9LmqAUzJ7anAG1lkYlOrdxq466IxkCsedrPaz
ol+3GuAi5tv2303thD1rNE+8zpe1yn5qbgaWqixKv9G2eSual6nO8WpK2JpRK54K
eo7wj8oa8p3nBEkWGzjJA1Y57Y1XutvhpG+FabfiZwQpo8akwY8s5wzyuqsQjrzG
TDBU74FPSrFvfRuFkjdo9czVfUII6ieR7VMjEhcupxzLS8hy7kpUoOr+333Yx0wp
2F+hwrARMugtsJ4TnX68I+o7miDuBihMXnGFAR+R+Nj65eReqwN73piwLDc9kRc0
9oe6L+amGOzI53BHLwSlAWJiTgsfjDHlzNoEBR+QMdsF8JZLRk0azcuY5xA9P/MZ
iOPBsVnwtZyOKocJRpqqmzkNej5yfaHYqY2Ukju6rUEHFDlrwlRRtaoq4OU4iVX6
6VtDKfR/pxuERimg8cyBaH9NMFI5Uhij1hHQeHpeEwB7c515u+w9DKa8DEqbY4TW
lBzp/tVE8JCV5EZr6xuHoVIaDSZgtO6eh4uAnHgNK4rsOELPt2rg0JPPNqgyxsUM
t8ZXZDneCbVJPYgrLBN89uwlP3/3Fm6+MFpKWNbLWKgYFT8tkDlda6FcatxZ2H3R
XolHdg6bBdTZQeNivPB/sdoc/BEHK/QdOsO8R4Gau0taFW5MHm0qFJ7gGaDYDUAB
N1h1XgJrV/3b699Mm8gDiEzyurQQvTL1dyVBjXfuoo/ek3/l19XAMxjvb5SpbcQJ
nsQMA5N4SKlskXUYxw5CcUWxb4H8CiI4tjrYzt6t4IyUr0xiXVN0kmdot+yY+ocu
M6aOeLcJqARl8ajZ2/CablnSiy30Dj8BKlZ6dMJvKHQT3wfsweDONWYC8SMZZCeU
UadgOGrbEny14LNrZOrevNmYz7bCN5CjlNgHy8rfdviAqwaKImjua3pgC7chD/24
bzds/plNNjWa7fmG3nQdwqSR0qPCT+s50hMRxBwgS9JHPT8yIL89NRsrp8f5AHwf
rHZL+z9arPSi4Nq+MEXYKyV/7jsMjNqpsFuu5aD9RYIVYCQcU+u/+hs5/fd/Crr5
aiA7wcqpMoTQrw36vmH5i8TU2AkScxPK59wpLm60hq+pckHZvbOTA2GaB2AJmUAR
94+XSUonH1AlWMj4D1CUNNobatdERLA8Bh1RgahMd3nyBpPeqR2vnwjMuSqxl8XS
Zq+rkXQL9lmL5wNtp3ZFUw0d5NFYaVKkFEzV0VWd8H2dYwinzsKrwDWNXfPCb5Eh
7mo5M2fMUEkOAF0TAyImh3Nkya8vCooCL/GFCwQAF8EIYFghKd8xWJwbf3DTwrkK
DCGLNy+HsoRToN85sIEhfwsgnuvQw1uXDlHRC3MgqgDg5NgJz9GaXr1QfJ0oly39
ciBk71I4NAdj7qILoNb7lASp3oDdlJHzgd7M6EG5kFosHMsxHYkJcp07YPhVIPvA
EToPXFBk+zIVJ46oYafyu0nDagGwyA8zu4K9Lw7AAMRtXTnieWpUYNYnHm8kNrNB
AZ/21K2tJcO3Y4ez3wZgz7EOeInNUSw657ZWBDDAO4mJo54Kzw2Md14k4/pQGzPb
cybKtJyQnKn+Uy8XU1EtKFR0aFBO+VXz+3eeIGhEt1n4JlmemOMEqRNvExoztVRB
XxoRW6dT9Gzw0uV/PQnYk4DOACSRdccjzK2hOsUSEBINAg4sm0tDnS62tdFjkdlF
lzLvWm/vp56Bp+gt/LMxToYgvySdTpd0+1LfTlz8OEEJ3lYl1BIVQxL/YXVZOA2b
kWcTYNeBHrVL5mFwpa7yhShQnPDWOz09w0SiR5Y5Hq5Yh3hIBJXuUfRz4PTGV7OD
ZySu4y9pR1imcy82idLUawVPVd+UjiP62kHf3oauY0cqECNzMJHttcMcr8sginFr
KFAYfTFBR6bGshQsYgUrnxVe2iNVBwvmPmvgyiYRDnGOf119dxxEu2WevTUfxrUF
PF6PTQRqzqcviVfgE+vT7lrzUTVdw+GYnXZsacos3VystlztK3LhpYuT9sttY0zu
VK1ANyKao6prD8rmCW1ZEfM+9vpiEaExAzFk6FjlOQIBvmdV3iEVdoIAVhyXotvj
N7AKsModmZgXVJePdvX8BASO5md47/gMsdOBKUjcwn/OjCOr4JLqQ6k2EcRBe5GD
/gBzRVlmsWen92qlOu2OkgXdj8BoHjasaG17SneC3DJlJI868oMxvGVA1k7LQtbZ
UWU9B3RXinPrhwyHE0LiYT8HhxhnVKTflQHxO3Ndkx8/n8dF+ILpGb0WnCXR7CRW
y0jMUXPKtg8hIG30ZhmF5UQGyeIwbiAGG9yWZqVVtCJNnuDH7Wrabrv++Iiuq7wJ
lrghft/4CC2l4TRmm3ras+6zoDOBMtWUS7FNGlLSBtXEUQHgFwCjAutcxlY6iu1N
n7RE3foE2x3z81ZpBWhhkbbVLAMJfWSzEZLP+cSNrvSajr3HpdEDI6KTGz58Mwnf
jU24Ti9hPiZi1cCFOJS/UwrzY0EE1iaPUO4YQDsXAeM8jD6qMwylWa6HkXH9Kh0q
62E5bBVPQaO2YKmep5mk4bYbk1dMiat/F77g/+D0ZXIB5yZKHnkomP0D+UZbWsM7
T+ptxT96QDiGsA4EABCrVk97nAUBzcLo9JXHcgJk8GprBEy91adNKiDa0vjnKxRh
+r/OT5Hh2xyC4ZX6cVejiRqK/JVFRNJ2Eh0vqHSYN4/n68Z7L6+XaccI6xbjA011
XtO62cJoQda1h7k8E7Hhoe7CLyvtoTzbu+jgZn1G8JDo5wV8ajTY7mdy2/2jCrGo
i21H3AdaBC2pqXBBkbQJszi0FTBB1ocpQT9sDK22m5i61fSMUx+5KItUMWfF5DTl
8H/7RKTlmUKmv1FVmHyxe/sGcf9EPbqrQkTILufbgH3AHEPBQZFULg8AOJNMf0KM
rkk5qWysj56fq9Kl/ra4bdZxAM4qV48wPmSP3vkETn1dnlERaKunHIiXlihiJhSr
PKGhQaRrrYbCjinVb0aGg7cT77+ieKAVEDppx62eFHZbwxS8OIeybN5DS8aFe3N2
BiiKtCmb2EG8BNbVEC7DCaEwihcidg3VfN9sHQKl4dQ6HmVhX3/uhRo039B6mJqY
kcvjFau3OqY6ivt2EbxMHnAU3PPMA5t5FtjWDQyylshxmRXcqAUjKanq3Jyo0EYd
UMj3MgOARZuLek9EyvkMW4HPqu1ihwjtiUuygYfApOI3ukyKtk9+ulpxqZjupUxK
MHs1Mtifn5JOgvIyHTnuisfNb8Ld6zgd/WddMmgpd8Tc3cB8jVX8Z4P/BYSmi5gY
zDk4a0uI88vTYi+CzFvh8OstyhLiP+RUrTRvkcJdmPLUz96WxfS3TmaUF/NBmjFD
oCrGzurk2+yhdNtUavkjeYdjyJl+ulNbehuSW10DVXiyQbSgCU3l+p7KE0hI44Qc
4uPSNp8H9cd6QcMpE6dCTv/mYfABl1eJcspt196iOxUJ6b/U8w+vhYIJGotTLLqO
8Rs7YU+FkoDU0fVRxZ8HI6lvrNkY7kilEIPyj7ToEFysQYN580ic7vzONlCu03Uy
n+kbzSp8QGKdqpClslPjYF1GdAHRNr7xMI4pgTJqePpcDGCWKbiZjZ+rrHlhZ8w4
LkDnoqV/N4Id8rS4CmgWJiBMahrPhoju+QquMqdnRi816rZ6X7lB9U5opck5gKXF
I5ifnx9CVkXw8XvBWx2lQjTk9fSxDHqLTTvJLKYKyzHI6VJg1mCzsaLfhNkZNVBJ
8lpyUufrgMZqe8IMSEN6luJS7iZVNWdD5JnsZSScJOkAd2MAIiS6ElvJQkjqxNo9
uKWPaklY2PiORdX+cfd8qmmdbtYwaPUtEqRa0GtUrXlBFiQaZchZScHZB5vSMl/H
fJfj/iRO7dTgXb2kRJqiAqJvIpNT0KBGNh699GxlgKTSL1uMnCrIUjn2znnVXhoZ
Puc5RHnby+1kcQQ5G4OtcD6vaSJcYWINmWg8HdMDz77zEh1R9G46rt7telUPiewy
DKZYdWcGGwqDrWZ+prNWHhtrCtbZ9r7vs4FkXvHsB8VzASm9u0+ZO4tpPzdWePfs
zPIc9zU3mMd+hiFnL+QznfMqbAKStV0lJgpYdaMKcjdsnFT9xHAHNY6mNw4nXb5R
CtwQHgOfw4ia9UvqltOSjQ/H9fzXhwWSmWH1A9qqMDRUtZr8gvcWmbXiBZhjwTow
2tl5DRui1NBFU6RxVK1oFT0uSa1gW6B6goL5GsEWy15pI8S7GLgZLV4oNfaG/Yip
fiFuVis1k6+qmKcitU208g3u5dYQj+2OZ2vxOXYeS+nOadZPUWzY403q5/NzFSwK
72wgo/BNRr/p+hv3N9BzTmqCfq30AoHdk9wuIdeWE/jMyHWDh2sNNKZxNGW8fnjU
cJiKrc7RjSP+nxiwcHQVvAvGOlBm+W/+nRhRnFYt43OE1a5Y3hXGQbvbavhePNh1
4f6JzSubVnLaa5tJwa7Kwk6T3ERNmM/c5X4aRjI8jBmcWcVa/qseqfn8HiQvu7Pl
Xqt/qa+d52QwoonAvusowD3NWn47dC90sJJ5xgxnRy7BLyaP/dGfpu5uSCHmLQWu
49axCQt827/UL5Dx2RVEFFJ7x3jkdZoDiSq6bqgi7bAFL1QtBloZCGKChTb+BwP7
guV1fbpJ54P/y8sPVmn3yNFxYH7CP+b5n7bE8BuSvHkxQugMQtSjEx2LJtiOVk7R
irf/aXaDPr20TAi8gVzdIKggrnvn2HQ3FA/zeqdYnx/hpHK4tVHlotg0wEdqXlpH
ojn02EklL0XJVkBV8BDP5Ap/9y6gc4npDXqPx1AaguPWq5Zbtzzxcc+AQv4N2GXz
qSIGK0JZWolaFujzYhCJK+inbQYCK7MuO04+K/g8atFY0ELy39Dq29ie4+4UG9pW
HRTndejoQDhEAxDIhFfSvR5aQXmRj5wyOrg4GQ1LtQZT+EdR52CfmuaDOK8PV2Ds
PuYJA9n4JSmUp9RLK77MElOLqkhyRn9imf7SGtnmDXPcSxdZSx/oWzPRuNwXPoqJ
VYDhnM6pyO7xaxQboaHrZUKS21Jdc3BtT2DW44hXKbI0+cS+cAKYXfbf+pUCVCaw
Bx5lo3W2af0peBqQl7t9L1DTIVcJC9s6dDzWTucUdXaEcduNycZSCUMWmpbi4RRg
NboqsaCREHExdw2bAgRtTfF2DP8+JqTXMiodkNnuZ9/D1ag5Q/bJ0azLo29Rcqp8
X1XcGnRvVS0Zwgqx9UWC7kUO00chQScipbwMoijV5ZlzMuxNROrGtho6M0w8LPt0
kMQ8v96vyIFUIdbaDA9RDxD+zutBDed/b90LiDgTu17OCyacNjRo4kywnjy5AoUc
sjOsBaNhqRvshT1ClAIoGbHlJKGgQNUWHCjj2UAlzj9+V+DsfdVQCRwEecEYR9Cd
zECiZ8NBDvrUURkGjsmWPkXfyJXxrSZlg6iTLFMUDqjlieMqb7sARJ68wgmEviaj
lAB6Iwgd/qWggJQX1UIWyvDCwD8acuf25yH5Hh4YuDTv0qnU+YOYJ/Upu/jnGJSA
1cc93O1DceRP/wiBOUz5F6c+XOkQYq+wbhWdT+P+nQWl5b1pm5VY7Nh+8/8KRnff
NHi4Zc+vMuO7ZIJWhSjwqZCoy0Z6T0sZ1aFhxqhtPdbLKCJx5yOcPdAqvOO7HKGT
2aZJfxCkALxoH2oHHy4V7JDuFh+VMSOUVAILAVn0IAn2GgJ0t00VwGhFyDPfRUKl
JnzUp4WxY5+qecZD2rnpQMBuK/SoD5VKoAJkYcda5ZtpyEIFI8YOG7f3g6yW5TBU
FEvVwhpbTkvSUx0nNRhjZXSrzj3Tc9QeYW9HZkxyEifBEF6jD0mIPetAU/XoBET/
tJNXgAXcEY8Ex4a17KiDKDBJLm51/3UY5U+WArndUzuL0+xctAp5qxBGX7VTniVE
LY+IznBLVAY17wnDSNQ0aIYHxh2OfOwP3iMhdhLypnWQfBNTWYCRe//rfXG7uem5
sGhqNPWC0+Oiroj9kEoKnIgyTZU7drCLb0RLj+f6y7xfbD2bjNwH7vU4n+OssL6O
twmmLOuYhh13X4mmfu+kOgce1Jy3aB5uci49Pn//vlZpKHjMcUyxTCP1r5wG8VzV
oYYE4+XpvAk2tOReEdKMSlmokXN0N3gGbeydliOVKPq5Su9RVN8FvH8JL0pFVOnV
H80gud1BhWDQRAzsEHiDeBXQ6AEEge9zZwVMX6HEogO+skVsCFOJRf5GcW8VuwSw
XoO6oF3+0cjhB0Yh/pHMjmrKcSeMsiL8hfWjvHNrqvpwGUl7HQJkjNhsEIzArXuh
afTGFFvpbTHj1hgJXrlg1hxlR8fVkvQjwRcEm+1/+YUdoCuoO1SLN84Qpnjk+UWo
rCYMxALccp9i6jWqHIQ6eI292gw0SjtYTpvzyhm5Iq+gbnko1XjJQlWT1j9xxxje
zf7I8mSMVFQ19mpL26CgZoHlO5VFF2ptN9EcA6PdJGVO0RConO51xIo+/1lWrYiM
jqm2DHk3pSRBl1+dS+Q9KWkB0nUMkjNzPQnA1/LkSBWjRZ8eGYIoVaW+rZ56IzzL
+dFKyHKfoRQZ/FgDQHQsmVOam19+ert0gSyCz/jJYgr1TdOd05JCgIBkVfmQ2l+K
I5fhqMKr7Q3TBGiwrdQxHv3qrhvy2Lew87Zf7JmS1aRwjEN+ED5nbGTM0HKdKxFH
L0OF3Iwj8qxkXrNYhRbxX0mzypjC63xmG6GCbR+JId/qnZCCDBtoJUOmGqcJ1AnX
RMGFfWtI30ZZuLEO6CGWZmq1TPk7DijNFb/j9Qly9RSnTcxPwAEGgdKJhfisJMKz
OLTqM8gwUoK6q+ny+52zpp3ESJGJqKUPkhcAGR5o/C3Tfo7Gt20LJ+swW5Lu9T+e
7Uh+dSE8NBlGEsafdp6sI5KM8kP/jG7sXzKdTJiydC0DOHp3T6La+P6mDwl91c2d
DHbdWQ9CgAggxw3vJp0sHnJjcAJOF8SqW2stj/w+fC1cyt7I6Si60vYE0M9MCxJF
i7XDANspHQPDcJXKKJGyksiSWrYsshCEq5sRiX1qRQ87XhmDPcP5tRZ2WQ+RxagF
K0wxaEXLHZrdCfrP2MRRwhuQB2hlzrlI9Gn7foNBNf1BDQcRatSQyEqCEraqkYrt
BZ5kvkb+38nNjMwRnj1GJfKMiZeF2GeRA8xZwGiFyKMp3luwjwY/0Ke+drlbGwba
TREMUV2JfyvfP1HYqImkD3KsRDaX25eZzpMFvUEDt6WexH9YHEDNvd9dnKsaADP6
yAcP9KPSxqjty2rFOqHERy3mMtXLc93Bvw/StcJ8c3eOsg8xuRFeVqhL1Iv6Cxj6
ud3Mg/Axm8MOAXdDMSFWl08VuH36SWCNOTmylR64wRE3d4qAMOlff/bkeOb7HR9Q
MBTFEJI75HKtwPpxeWmqjGiDauqAhH7RSyWbcrve15aDssIMQy9SYTAQ3gObAGQV
ZnTmhfEn5ygEojGltr7DmER2Wu8xS+rLT2mTWbRX0O2fpDcxLOS4sH6YIgwJ6QEy
wXuQQggrf7BT7QjAyokqGFujRUdsdjwGD1caZjfBSXH5wTyp8eMmJmaKIsh4IeKZ
rQTJhUxYmerjXCv98U1gvKXwNnDhj8hRsRdPWEvbRF7mP62QDMAu9jOPGPDus3ac
rqKAqlOux2DYGBCWdZlB3WUW9o33WDmm73GUeR3WAZ6CxlLkbcMat1h5LuW3oyeJ
Gvks51BaM77aKGsWsfDYZcuhlf+DzJkcHV8GJ7oE6+mflGSZcytKQsQquNovbHd/
XDiEBTC10eyor9F8FE5nBlJhE6MKZINbv4fZGwDLqBwRzHFpHOJQsewxr2Etyeu4
U/c0CkVeKW4aPST0GNXkGeE9wEBleoFJTDwOKVqkXX7s93EBHBHtoTe/F9iouFYb
3f5bZgfOzGgQqaNCaMyAajVmSE69rc53iFQ3dj2rUkz/DYAKxBEek5MYcvb7accl
FeALMMa729J2svG8bGLsMzngSbMItKA/qG9CJDHaZuCJOZ5gpBWJ/+S5jnUikvZL
CdUYZ5VbuvzqJcfJ168KK/jRfawLBriuhlR+Isj0N83O2WJg9Y2AksPrTMEkVwy/
bENN3HPIldcdq224ZN4knQsE1zr2X1YT9DiDQ+TWPa4n1/vCbp4C2/dtWEEsrIl5
K9fw2sj7QrzBrLhmh57KhqXzqaCjbZjKxQj1sliBXC64LSsghxwdHumv/gbT9XO1
yGpFHtKw4nAlezsS7ZrnuOzz+Fq2nbbYLZIhWt39Lsg4a1OY9lwLuSyC3stYn5Ia
JHZhlKcmvvdwNlD8YRhc6ICuDtbAiR1T+1V3MHkXarJYd7ekZ8JlOSfeLXJJrXhm
c/irt6f+UYNK+vjGdiJFNshCdMsyucRC5slndDSdzFkWQORJFa/RNugE0kQ70WSx
7Evfa67TwbIdYtm6mhIbjUQCIMTG6cKLZ5jDF49/D9hKXtMCaLUNL0lzbatbdxd/
9SM4bPFan+I9gJf0teKY/4tt2YdzeMZVsimeGNCzVkYzsS2gCmMODSptZa2oUFPU
KErw98+Crlqg0uvDhrDnr9ATwJQu5x+fK4b9ra+kQI8wyiQvU9l1bdco74C92tIb
AjjXz6QyGyGxxltop7sKPEn8plBnVJ1J95KAcWwXDl6mikoWyIzf1v88rqjQAIKR
azJmDpwjc4yw0SPHU6Z1iheRJEn9aDmGzI5bIRYdt980To1velP9n+Q9kZxHkzPk
9FzKuKSYkRjvY8Q1SL20yHGyoY1U34jDW7N77fb75JSIyv8TAqKpIkhRCt39YDR2
4ME51cycWEfotzLSoFrqko9zOqkD0zgCH74Qoy41ksNrD20MaieJigwr6KjOLAAh
Dz9y1bDVstYquMoIaCbkBGeYqbVW55cbXRYaUCqysGrY99owBPNlhtUdI1f+s5md
g+9ACNi7QEUp+Sk9EJxEkOktAY7RIdVXIqRR/kXx9SBrzWNXwi1ZtRbFjmnO58BP
2XIbs7obKOrqGG27OCyZrEHF6dIVFf45/F+Q885mq/+Zaevjaa2kZiqgXIZl8yGt
2wsk39COpjLz+MVOPvbtSNZCljA5oUHN9e1I+jkYdey10WmFAtSQZHJ2205TuWc+
rU141Uu/DjHx8Qtvts5/fZ21iX7D3V1ky/SAfh49EpbPgkhEll1IsYMgTcjGf1jc
gyyEnAYk/3X/08cA9mkltDbtlinV+NejDaCYaSKk1l+4uvtXbcSPTvEWbosOUMzV
QVeZGZmA2wAEdZvr4TTHV5zCe6mMmKAIm+7KNxCWQZGEDFSFJDM5bYorM+Q05OwZ
cfQYREMvq+Nn4JnkwjfjMc8Y6hZFaqqH7NMsnGF/81FCqmf9OYEaKcA81old7sJO
S+dYh2vcErzfSyZy/GLg34RxrfyuKtD4+QsmCMILZzR7JMnEH603vpOaRnc7mWtC
BvKMfAeAyMlF18r8zZawn/IlSaD3sFPuSX7oRVv45XueMYt3DkJL6gi4RUzK4twb
aCPhby76lCTNBv+nmw+Y0jZvsKLe/el6qT/0g9bU4hBwT9e1QQFPPCHAGN17qayI
beoHhtYphrgnq+d3NPRGclBAqxvrkVWiEyOkdVfdhot67xPUQ95Qa0WTIfI8vPrP
yvsS81hE++Z9JcWVhMhiyVmZyIq2KVIxPNMuyc2rCAbrqDZ/g4LkkZ1BkgMnd5wC
Ql0i0bYk07Sp80RK6qavSdhNO6c49H4ZTE7PKfMkAXwtQ75GeKFNfui8gqCkHyjD
gqMLSmhFFxlUg2EKtOzYEWSi80a0918AENQJ1Y7MqDCDVBpiaYxLKbzeplnVGYuN
sMoaz9TR753MaVp1278opG3QWmLwSyBB61l0aECmNWG+1QFODYmdQUQvTU2SWCg9
W0Yl0Y3Yf6aPSZrC8xMd4BUuiB+P0DOJREtNxdYVzBhA3kCA/XT3ZqUjT1+UIh49
Si/r9CBf7/sDEXjnU1s8UhMfaW5rdW1bZoWoF7XGIuUGr6++qCXMqU6uFXOeoqIJ
bSeFEOaiXE+GWTk/mhG/45WDjJOM6AGKy/G9/IdjkHV7Jqgt58IVAgH67Y6++Jj1
Uhjr60N19Dc9s6MY4m9wG6Iy3kjb0XGwHklXXI9kX5/tYgwcQ1TjnCyZpiy1ukEh
cdPhtY4McG2WmcgNnHSIvQCjsYBM4pCC+rG4emoVsAlhuyIKlyDhleOattfzlQU7
wYOsMSowwvVV84IZ3+EiU+fApd5PqFrM04TXqNCKkWWGu2oRrFeqRKb0et5ugmna
GDCfZsU0NCNeoQ7VHvX7+L5dhsRZ+aeTQ/HRY0uA1Z3SpZat6E/KRoJTQehGD7Vf
SPXY+cBOL27OYmrRNDv2lted8TZZMzPE8H0JjgBHD0XoJ0g4l6NQog1qF8iPxPkG
6+inahp+i/eQHpdalmreJRoPedixBo/ZJnjLTPjPFcu0WTw0q3nTMsGwEj7F/iep
IjGHelNd0qml0k+JdzFkx8E90fDeczicI3aeKmaG9RuydNruUc4OWQ7dyTOcRU6Z
yq5S6fX+nX+Le/24/6uP6rK2Hr+jXcRybrsGN6Exu2a8F7weus2utQo9eIcs492B
y+2zQLT796DbQ7P9HeUTkfUUrXNldhdPyuanFpGgXG4lyIvYrsfEr2XnfOkek6uA
WU52vU6IBEbrxAVtgWwVXejYMH+ZvQBHVEh9uS4D5G4X9t2TI1FnzuET7KUYNJT2
6qHGe61kKQlt+INKKISJYJpKCCX5duV83rnV69hS7Urcodmi5pZIeE5NWZujitU6
F6IZ9mNCL9MPozGOU+BxmlLIWDfDPFHehfOqwITkA/MTciR0fZu+pLqf06UjLadQ
Wcuim5hPmvv9dkvlwBm9P7TpSjuv1dATj/g95WXnSGvkoyrMNefGfBipkFhc+Tsi
mgIi01per8rPibCBAllxvduszrf0Sk9w+IuD1T7NOzSZjSF1RhnEjwDyYN7DpiBU
7BPYtG0UwUvhchKc7oiC2lO37s2nKab/FhjfO00WkCHFISa2qoJwFghHchAnF8rw
4xHsky3E+cbyLrXY6DE/tzBR8qo4VLXxiBCyXKvwQZa8vPvIJQejAKNQn0cPIrPv
cTcgxp6fVZBYBDchVwA/76CU/G7YMUwzNBIUyEEePzst86J9jHOVkAqcr7yiOSPf
bsCSp9hzA9t2Z92XzKcD01BeEGD8uq/4Rpv9QAUAgDMGkbamhPRTypVsAwTeq5yx
1OW3NYD/8iGZWfm0mPpmftWTQsGB+knt4Bhk1Mu5Kf/8KHHQP7x95cC5LfvXyxm/
tCkP8GC3Xaxa/M+OeVFPKbM8nZHEbE/aG6FRsbBsfBMdSllApeFLbp+w7xFrxsaV
2SOYDjx5R4myo+RtCVlKkFpgwlhfUMwAcE/MikMQFuY6ApSOud/VdsYrxT0aOCDx
2vhpquaQ378NtxWQ+iSof+hWAnIvdNu0JX7CAKuJISg+Ae1888+KfNa52G+PZOvK
6u2Bmu945td/lyolDUb8TQIAEC3n724Y0uYi0x/eFi0ELqaY+DGZ5L4mpouC++k9
nBzTX5dLJd7kcPlElZM0BDYX4i1d00cSeb/G5EhnYFsKkeWIe4+7IO4pV6/ZOr6M
C7dhpHt+RR6vAiVlLHQIPxcKxWFA5vx984g9sUpQgqLnGcf2ZVYnXYUivj8h2hCr
23vqTAsd9F989n96Wecs0fBDTFTKDjye8eZ9pSwdwTsAOt5/XdDphB/W57Y9Qo29
GVBUlHvRNf8GCWzwovx3zEy3My1wD8GBrdGprcr5/i7siCB5URqN1+5FUNRL63ZE
Ytxh76MaX6m4ppiMe/Wq5yYtsYRreCquo5zvnnQGeqHYhDeL0rHDvvsRH9IY0Ojj
wTidzM3ya9Y56iWIcQ5MDoeY7E9XZEyJqJWkcOUdy1/0mfrjb56wJLzBvf1bAsS8
FLmxHKLkOvEcUor3K8k+vjAoweL+kuaiG2ILmSpM+u//IbHBJVX5nP1lJZEQWxrt
0HzTfMwKIkr8E8eHqEL+falpTc3n+YHnMvhTLrbeODaAbMjaXYbJVNxTOPsCOSyB
NC/JJiw3W2tB88l1VQMFDyrEQMG2cpDI36YyyYWXTgTheY4VYlc4B9nO2jh9TY9e
HKwu7Malchf93qboRTOOX4u7A+6BpXDM3X6wPcFsHrJK7Qgk0BIjv8g2jqWe9fvs
It7Yo108ZGSYIi7cAxtRztOAucnm6JD5mH9vtR+fBs2jbOK/t1bVjMmK3+FKdm+b
gNswQr6vl+lnTrswbW2lZbj2Fa3bJUuVSOk3NfMYc2BxDj1AbIMi4vb31+OnYd/n
Oy84ZURZZoYGqHhkSzcP0AT8lt/35pFJ0WvkQpvw+wHLtj7W8Exigb9tu+x4k2wD
yV+C5DxEBDj4057XrWnDEnDZ0liTSn9gnveiEt+tlpRWiet+6brrMFDDDQzxFoy+
iJUdakdUHTN4t9ITwmz8tkjON9jdsu6JpkrmrLbPGp63vpku+aANo99BUHW4io7U
6kc7aMzoaBfsEfQdFn/010/k5s+aCTjptEj9UFhr5/e2wF6wh7lnhUMQF+nsjb+A
k8nPh3FWAJ5TBgOK4ezaEFyS+6QRd7TLOEZrvUbpRfXfL6KJarbEnws+WbG/85ca
jcFp3WSoFhPpueSFt+9Zz/GzQ1wlIyGYOPT4rgiaXEla4V2lUZSNY9Nnz4WhkMNZ
O2tbMgOZGCK+SJBD1oYt8XnQbAqRtYj0duDx//ccdidBq/m420XUMAXBNwbYky1W
vYT0RleDPXOLi/GV3+7Hff9oKjo07cIprBEzvn7sKz4AeUlzK4yzIi9MRwzlAWy3
0ip+AU91faKLy8pf9NYgeIRvuqIHzfJ24eHdtEppIXjHLuqF2bhSg7buPvTKxZ4i
sqQOTZ5ZAOyMYLmfH9v7jzXgz+v8GgfrSKaX2UO6aFcBCMInXvp9JVgu4aSdfG5J
bmnVOISpNU+XmJOo0NEJK6sqtJknHY29BswF8Itx3Ia0A3ZFfeAPbxebsyzpJsCn
jzYdhHRlbVtgP4gGIWhqQ7VBcNcp5oBdjFLKGgTGJHJvzvlz+XnE1sQ+PcqtjSck
WzHiFSqjzGpBuYqbL9vOjZpuiC3kpHd8yz5k9Nu/kY4Lid/p0TSRM63guZwMsKmq
PoqcCp44c1V/MuTzt8seIduwHaO2c8rxRzSYgXenKICP+i7sKqsqI2jeJ7yWQ1gk
axd1z6PgYtfTzpuFHMXjs+fsh4DNE3DtV/yoprApfkSpxwsr8xwtOBd/jVnTI64R
VZ2DiRTRyAA5Kpu8AcZJFB36RGdxicq2UAubgKGae5ekf1RX14Ck0zlY/s4U7FbI
CuxMlTGo3iSo5Cl92I7ZZJzDWbYQhiP2UVtLKaO5tUzCaa06YO9KqNSeqzS3n6MF
qhVIUd2N6yKs7lsA1uoQeNmxpoN/Hntg7EwIzn+ohV5WkGXaPvB8B7nHaTBXrcCr
zSSvmRvlGtIiyQEFqFf5i3Hzt9WGWLaLLLo3V4qqWAWFKSQ49wZvmVxTxenqV4kv
fA5cenUfBbooV753zBdVXMD9c/SuMkDtFGwgdnolVlSrs++h4jLt5DZgXfEG7deN
7vwkdj3ZgGdsoo3MxUMvYkQQI7cqKIaT+MsXur7XJE1SYyv2aMiX78SZiP029Q40
anK3Ah/lHda6rDGmWHieaiS29Z1QlZI5EyrFKC44jLeS6rRT6MtoixJedymZc2yy
70goQnQGan0/kcKDObGf5fEDqrfycEzAhGUZeSeMqH5n2MKS73OH/0Zt4rstBpo9
K0ifykhWa7RIqquIuv1iKmAjTbjhr3aLh2pM03Z3lZpO/QuA5/GBcgRUvMcVZf28
ktlgjC+S2K7Qa/YZbDw2PCIVvmQMmTPaBxxs1dzkwsLe6MQe6VupSx11qR5ImXVh
ryjUnuIfJaJLAKZrUL3VAyQT76n8yjuflrOyT2JykPyXizBaXfpYb4vtufDv6PEp
iKUaaZH1I6OBGFc31joMRC9BwncJJDvLIED8jR1wq20qCfF6DjLUfeg0C5etheX3
6LfEcwGu8BQi5Kju+UfN3BbZXIAL2kaNIZwZEm0B/2cURAdJrT8XWwEY0+uaSLv5
HfODPdpo2mHGBeY0owoYOqWhmaYno6rKPem3XFZYFiGy8s76oCCkvKOwGftVT8BB
TVHBYG8GddDEYHPmHdblluuGBQ+JLbvZcEYnQRFa5bXdjdE7yGWw7WyfeO/OF2El
M6Mq/pXJ7qEan7IeKUTr9df4BGj4BDjSuDtOx1Vtg+KXuCqzxmmHhgIy6chUD/1T
NlaIE2HqBjj55KNf3O0LYtplt6xKHzTAeHT2DM+TgotIZylBawRUpWsWl/xuCUaS
RX680+4l2qcnedl3q6IT8eUZiQjpSduE2X4KHZOo92u1ghPTFev/zXU1YhW2IXCa
6HA8dcfCRrdwBqaPREC+dmxRUM+JOyV9gPwTgU0w2zbHKSlJT0vdYLUPMpVohT2G
gRrtTQ/Mn4VZDTuaL2CMikjU3xYGy6plNhCQ4X+nBITWGDDf8JdIL5jmvcAUm+UV
FHZG/WdzXHnQOWEFZ47EYd0rwVenFGIgvaPziW7DRa3zZ6AgcZ7Y1sUIJvUhN1ZQ
425dhqRxOYrhumAJyQPIKoxOYJwezpMDhe3o8+causlVNIlx7tqGriwcfknn8lq3
aSQwGjjJgWxA1Vg8OXQukpiEh6ew//qce/3Q+0YVHzzFI4z5gEiem1dji0OZLEMz
Ox1WPMeRnlixViXOssQRHJkRytgJecbOnCQTkAYtR26rdGfKjHq61LXVrEgV9G1N
PXqI6DKT6Gs+UHVALKxWSx9lk8xoxuCAc9Dpx31J+cDBOwLvVO3OaG05/l9cQlwO
9beP8Pya1iTVmYDv6x3xdKB/yTnyZ+a0EowiVom+78OLMhYjuYoMxuxMC8OAPL2d
B/A8qtea6hZJlPJyxknQQ+rqoX3K24fdzv+DLjWUq6Y1plvPiqFLV0Bp7yC1QHKb
9AXma7fYxzFps72HhorhhUSAEdEP7+6BAocYTx76aPQWwdLVdtBpUKoVNSaZcHUc
ZPAuJOTc0WUQ/PtMXOCewHRU4+lKpRluGMtfZzcUoTBrhP6CC+NG+f6WdV4kV1bn
GPrlITCxcJiPTm05+c9V4arK3kyR69n2OkSDEEzB+aoxk2H/E14BKcozrTxwHWsb
bioTkVlBxHTL1ldZbjYt4IGIRynuW8QYphMvaOmKVz+EYmXCEM5t0BTeC2Dp+b4W
5ompih/Baq8B+NDWMrFLFjcbo3s8ZkMPM0bXL0836LKdrqGSW4OMd32PWENJuZRy
h7gIRbmpsg3P/FTETvqxqWVMG8RmxR4paUJRZbjB9N22b9cjGIjdv3LM0pw+Q7oP
20SPbJqaD56/nm7fj2EhbiiVDa6TA0VSrak/HO7EoNo+KmhDDM8LZvISVBGhOiJu
fRIf30bGc/BopLiLln8m7miPTjlwqf+ea8zyfH9IWiwjUEzYccR2dhbOUJSHME60
xEmILSclCl/YW+OMPDyl2fAlhrKinDFo7+Y6zaFFywSWgoMdO49/ZmhGnpUM7GsK
vXT49ouVn9mX/k4V4+wdJFKspcCcUG63cbCcFoDspXpsLhDe1X94p0c/G5iMeBBj
ii9uTZOmGpYA5PECxeCPzpga8lkiXDAIxWIP7FaT26VrsCs4Uf/XKNgFLk04DD47
jnx+kBZd9eiFXpd/1yoZ+VdGD8r/8CIkaVgfcS2cN3PfDqJzDpmpI7fLnlItZ8Zk
IPkNWHu+EyKsEFLMfxDXvFoXfag66o2BzjF791N+8Txbo79joedBK19tmJSugvGW
yBrROIsYJCAKzpVzz36V8wzaj0I0moq1RTKDYo6BvhS+68b0gIHzBYcGzUhup179
iZpSBwQuypiD6Sm5aeEuA0mN7GYTX/TbVOn6EBJvtsnCCgka2z8tb0NVTThy9Bh0
11QpIoydTOGOhMi2eFKuyk18yhpRJlp3ExuzIAECsfM/hJXW75X37I+qFq7FqG2y
8Ulzpbj5KzgzTRFgFzFcL+Et0hMqGVPBo/4rTHpWQfpCRlT5MWtEnAJ2znCdY//n
xTpzXsbTk6dlJLudA1OnKNX9p1jZZaPafSCY3mu9x5qa4isq5KJzM0r9X9zn6qwt
S0mY2O7y4e7pvX5PFnswn2UTOa200Ab1P9DTfrx/ieRBXZMJiOemyPhtr+Jjv9Mi
M9HVM5FbANFCSAPgMNM+SRp/TpEu8k+QpfXTCG4FJc8vVEaTGdB1ou7YGAcNqjD/
DzRWp1uFI3UGBm42N423y0td2tx14MOqLFIP4UeHeY8CiWE0aRBg6VzzvbXNqn9k
tJph9tU2n+b3HKPjI/squxFYxP3yos4PetKlelkRGkRxomKXkDUsLn6QpxD6uNPU
TTy0pusKNsW2TQbZ4lg/CqPi+iAe/blwHVe23ybPBMFEox/7pKguZEjIkii433dJ
HMp22fdtjGf5Av+b7gbXMMBp1mUoXuBLe01w2bfr2Qjw+CbfASHe56LFndm+1jol
PJ8Nd2zzZuVFpcv7wYbqbqbbEuaCMDBoX6+jQtuL+rvLYJbM8eUk0FynCCbl91kX
cJORzIcT9X6DHNrGXggFFJe+E+DsVMziMQjv6uMdwIqSvthCOh8tz9D6nc7PeB7Q
YhRnNsEpmk/1T465WvFnvSP9AICpYPT+Lqm575iL3T8mlGWYq/6mJ7YP04Ute70D
S6a2O8P3CnnsJwEeogVZCr7CftIHVBF07nhG0/g+30MP5wKm2fmiUB7LjqnIhjrg
4j4SleDUvaiIDD6qwYcyo9lNt2oR8bVMF38mqZCPuBFxmUcP1ajHZki7v7vAlpf/
H58LpqZiNKrye5D6hoAkzxDIfz/xa3iY6oxBBjQMWJQiCKgBKjHaehxYbRne6Rxa
6nn/l1BAvy2cBNc1YmKjf/3hbftw574L94oO6LOSA6MqPz///s3dDfMEkh0g0P7f
8kcNVIqMezkrWNlUP1KrCX3wBd7BI1Vg3TSLalGXb8Y8ssUJaWi/dD/7Vqihf2uw
C81/CrmNZdsbC5HV0uY3wrwq6qO0V685Dvuy0xt0eBdzfS+HDzMOuIAKCwefVOpl
p2qBe+Y2MCmgkOq/sllxuRhfL1swDa5FV0ynEczwmIUIdV+iVeuktF0cP3vgfWiz
UNX9K1PxE15TVwTyUvS1C/sxgcz739EyRWtklGg4eFrkiwPv3GffP4UAxaXy0cjR
CYDY0x+OYGQkMQzxERCyW4zGiMz5J42ZBYnlQW2moenJCPgdttdw1mznbPRkhUvF
ujKMv96hK1cJ0MHospwOXLEF0ZEj/Tw9o91mPTWvuMYrksZNYPoEe4PW6Cy04f/R
fSJzIEYvvaz4t5OO9GoQfXYfXMIKv6g+eY+iyffGvmrv7temEgn1s7e483tjRe+o
f+LIZ6PDwPOx+BONUBI45Rk154NzInd8gzTpXBMWuhKRMLdykA58ElJ0xzJq8/GH
YoswjcC+MzspmumkNQuT8M+cshtp0Yu0NJ1PLURBJPYJw1J9fnJWtwjK5k+so4EK
Z4VaVZuE0ysfAXRABA+3JyTHm6wMzZhJ1kJ0BXjTGAn7u+uh3NxXCZ8kcMBBXV7A
7JtCjMikrghrPsdciNBcCszKLv34fjhG0E8FDQlRrEp2PK5CW0hHLSTR84lK1q+k
lZEsP7Xx2UCJPXL7h/gEUOyNQtvJHLPyBwUb0uQ8uB7Rt1oUaH7JkREuxh3v5qtR
No1sSvvEBAZVSwXmsNoNZkFVIYGhzWsaNBOhTkjL5V2x5lBptPu7YyxEIclamSBR
9f9seZ227Wu3jqtgJjmo5MFkg1QIkviYCQWGxNDUNG6Tsptyf4EriUqU2v0VXmvc
+IV9SvgqdGkXRDhPyAwsfr1xIa+WiradA1FJ1mjaoyAASQ1vmzx61sPY5U564UMv
QKiDHakpRug3Xt1yJOu3GZNMSzHNpp42ZacokVRFJ7R1wFAFS6WdRuFegreAQZv3
SfNKa2lN8URXqz06sOB2sLyxsW++OXO5GMuB7sBCRPTHtBDt6gaDScc7Ra1GiSOb
hfhUneZxAXQNwFDDWX41fau8A4suQkyoftpGfoL4zNjkX3mINaORVqTT3KXhnEpq
KRyoWXnnqrApE5DbzIqK/B7kWRFKPkFTVkrBplzx24c+wf5EGwm2XR2AKa+9EVE9
87iuRQQRLaWLhHHiB+RYT5sN7y1a8aPlVEUicuG7+LQnMm7zfvc3S0EmWGItwj20
m/h15BPjCMZR9FZiS46fCSaZy0rO9fGkDZ3cvh0ar8C7B2aKGnt6tLa13QALw3PQ
6w1LyUkfupxwL0OpVAIE5YwRdg3jTnNoF4UbUUWTqA6LDa3VS80y6jokm/APXWfa
YCgsTDUJnGbwUG4RAEZiqqMaO/Lq+JDLELGs3v4l9ee5s6Hw5uDvNwINJ1qk9fEc
Y6bQCrP7SjD5n6nsWDQDu5ouV7GG0Bg81l3sdNvNO27H7vPrNwGdLNJzMcO5pQ1R
E8H8npYkBUIc9MZlQ6ZEidYwTQPIxsxrdmygbS71jdGEZJV+uB0t05PVpvZ46Gbp
YcbO4jXv6O6xhlM22qsQrTB1UJnYv2gQoD5yNJkclGl/7SmU2nei55+gPcJy54BF
P1MzsqJzuDnAjQHw23CcWkX9Bh48U4p+EEfmWcFqnpLohA8WYHMvXsDjR7qx3c9N
pcd89T1nkoVz85rg8hsXPsGCwsh7k/ld/kRh7Nfl4PBiEvxrJRLupSDux9U8Rapf
b23+Ha2nJ+NOXPaLIbfM0VhhKtaOTqvgK+c1zTxsKwN5JUqcr41CYsLnm2baBiHH
73srQZdsLvpXgodyN1i88xcxWwVfq1c/OZihErRbW2QB4agkY8kEkP6TqhUNHYOa
pII3Vatt5qv9Uz6TQGrAXyVLPZILaNxugf7U8w/7Gp7bxGwdIaFaMN4Bl7s5O5xR
oG0K/81E8rpFTKL/Z7rx0qtKSXwAoHEbHLOexGjpzu4XeVzVzT2hFnjBA0NmVZhZ
RzyLP+1Y677W2rydyPkAsmoaaMMu09PoEVVJHWdwzNmiz5iSnwn83WswUUsK7toW
IgvX+UwhBx2axDgjVJrRrEcPfSgnCpMbuS/qOX4FB3IvN0V7VOrUK7p0P6jpWi4U
clwP+/vMbH5WZ6AeOg4UrHv7uvoWl1Tl7yotGZM6YZ53xcefaiTWp62/TDOCgo33
0oBb4OCOVXY1Jj6h6lh7WUkcBUejvdg1uG2b5d+rSScm0krMq2ZxMJBBgtddcGtj
5ko4WgWbzSsX6WBE6gUgCYGTmvrNqur+6oinRh3Xlrlur59Ixsku/XcVmNCwq2gF
aBL+z67ht33HAsobzFcTSTYV7ert+AVvhLtJZydYh566oawBDHPBL1bnezHEtydI
r+m+UJ82OnyoUdip+Rcr1WmiaKA8SO7y+Kj7bw7bIR+nELDxgjwjaTmmv19q4/jn
1mFa8hXkfOS9Zb6oxy+MH0Cq4NVoJdBobbtyaPk2zW+ocpO31mAzOjU2u+5PKfdP
pAgpazhL1da307iT8/iXxMD0nXqq2ZeTnLDTh82AWD/9ltCZldf4xppfWzMpJhMQ
E5rapppxbYFwq/Ff0WAZCwjgvfVrZ5iNBIwuoG0T8hoJgqoIS2h4PXDcFSPXGLBt
F2B0ArgXoVeDStnCc7JzgRrelWIuejoWuNmWerKhyfhCyKbGI30EI4zNz36zXcCx
1cRB3DhUZivHgmH3aWtCidyfNM1LjvYSE7OFxa87ibeyywX1F/0xsVBq916BVmO9
uvACqrSsbvszTS62QbzuuNdniYWMiIm+d7xQgrRRQcPri8tkbGDo3v8rijg0VdC/
gWJvxDXXyohads4EMA1JOjeT1Aekbz/oi6EUiFwt3mZZZjp2giGE63u3RiBpBehd
f4GJz6Kidtz58oxOuwrz7oXJCXoAQ/quEWa19MkwfefORKlV13rzuDppC/pq1rBv
pF9flfV5AUBxfZ46FI9NfTOMlbe6PjKP13FA2e7DK1eUzJHjY/haRm8VUF3SgSTw
O5j7nxhyxHI87FrA9nAs9DSerMCanubp96lfWV7j6Z+vH1x2aSQQKcrzaEkhrW/P
DocxMnjekc8YoQ5y5bjB2acJWle+384EJ95r+/WpcHHGsT0zm00lf2YrBTtZgZ/b
UoairMA2gpRpTSFL5usyrjVSELWiLvF6U8nLlDqoMjwe4HqUZoKuJidW42J9ghbI
lmNl7zVlEpJAKSRXZG3ltG6vIsON4Ke8ZxuW59j3sLP/v3D9Iij4Pm8DBkTzU7nV
mIaZWXww7vvcra+kVyOfPo7O6dB5Y3vOPzcYbQ7TcW9tPeRlWQ1eDPR2XRXXg4x2
gZXTnyN82jcD9vn5y6tse7p+LH4ql/Ouyqd+tpNpAJCD7bn1nOurEyzTlJ/n+4U4
rB/MDu+KXOBrna//9FlV3sGK5uC1zircQDoxlrfewo2J4AyzEWwMHLaX1NFQ2deo
qbUY4UqxaG/Ab2wYtW9lsuDyb3z1O7Xcf9QORkbTCYL7Td545Zft+58D53h35QiN
7B7i/g2+8ZA68CgVAJswBxoo9CZTDiqCXQrdBx089MIPaH37G44cZ+eAJMNwax4c
0Qt/2G3uK6FLqikZLoH5BEZb77xxmliaQ1tcb6vj+fED5lQ2/XqSc1i577TIKSuW
IgFJ9EGtYl4RlE8fuCJyKNhdplAI8YArE3IYWNxl9A1abu1AZYf0ZjN+A5V3Ks4O
3+RK2NtqSIUIJzUMIw7nggiVKQeEeqE0HKcEvIEqZ50W92Fq2kA8TtHwm4r7xXQW
h7oB7lCtEsNPMe0fPNINNY1mnMRqkfMtCxd503HMsn31uzutKhq/hkKQc7v+5nkZ
GkglJbcSHomwvonZeJTig07anLbjZGwhosy47TgpOT7ZdxVd2FBsCkIuDWehHju7
GMcXoo/HebzUXwOYqBB/l7qrcQnkBmBnk10TAOpYgVZKXegjGTdywfX20UVKB3Um
vGchfxr2ZSL8MmaM8oXldZ07qIp8alZbp4GQKSxRNAKqWtASfypFo41yqxB2Mjrd
DS8yLLshIPTKK+flD1rMSPsN8BNuZMeUvaTl/qqVH5R/Ru3W/eDvYKt34xOZ6pUz
9sR6WLo791wd3hTM8VVm/x3KvfeoufUwai3OP4vV86oP7cCa6FQWTTYg04/CD1Ah
UUQrvHcI1uc7WJeEz82i1WozuUrotsUCBAtRZG0rML55qpgaegAt3YXxJg/uP0wD
6yTGzqcD0h56rHVxuuU0m4MF6yZHBY99EyGkQSDAIVQvx+bxn8F9Y0WvR2m6jo65
5S4vuam35S4pX0WcZVh6DrCB+Pka1IzHg0egTIcYcQS3d1BwM3pmjVEctZjcVU6R
WRZlw/060YSSOTZPDNiFZOuDHXED4C5Z+U/qekCTywlqsgATg+Sa8bJ1UgatJcA2
ZDHglAAR3DBGslE/+QXpWztdHMIcwaF1/NGD8lVnytYmznMlWgtngIkq1kWYmS4B
pKLs8ipJz8LW27qrfPXcyASoCmtRBhAXMuP+bS6+HLf8a6/wdVebJ2c5mx4gSaZr
aW/02DsO5bA21iSlvjjK/1/gi7wTmpGaJMcSJXWzkpxho27+aaSg/NO/DgTDctS3
/MFJDX/lq6e+K33tMEe7FqdixlvigxgtZxdiSff+xy9dkvDY0EjATcz65pGDsfyp
JN8jFXRBJEYPwi5Lcwf+5+3up4WAeQ/ESwxUHQnryIAXBUz5r2+vPBxGrC1vANgT
xH8hs0J/SbGCcq+Q9bgNc5T6xHbUTu4wzbOIiot+E5kzBGh5JIvRjQ7ungk2SjSK
w7sHJ99EWfJOFwnGOXJXe40jESVbqlsdLRpJuQc/Ljp5wqihiLbEo4fZyhColGAn
9MmOhgD46KhXI7n+9mSHv2oYGyDkRMCTcCUGnKPItptfYR7QO9iBuRPoZfccP4A9
FeNOyZeEHS/FC7JIhBZjH7TnHONEHYaKTnd1Ug8YIJxcScRCwukXv08b/qqc9nOQ
t9mYC2yWuUsCrmV9Fxz2FKsTkMKlB4i17qTWtpJJJ8OpY9nXjq1orXpHXy6IAHft
hkmbPRqiv0FKzO0R8pl7n4smNjjInhVY6YEm+ZZ6tbjrAS90tT7cb5h26FuQQE7W
byno/VPHkQsjpgmRky5onfK0KFLUCl4z8O4B3/qMT09mH5drK9HiQnPFYPGt70PW
oyesdFHZrscqxk7FtlxeCneHtAiISCbLlKHtJvnuPtIq1sy0lATaqwrdv4GjP10P
ltdYq9336KZgRAMKG0HJiwDJeE/KyYWCWtxvYKDZ5sjPTmoXNIHYeAzAtKQGLvQP
kIg++7fSC0REOTVHmBmPgKNoWFpm+4Zw/8IisHZvkWWm+TVLauq2NIQ9tkJRh8iq
F68DLKHm5n+Z8rSDzC7iA25G/b50kx2PxZ8uflUS8O5X8DYeidWZCV/CkEmoZchq
YZe2tNaRCamAmtiPkCf8hI54mvPHLLdg4/C7ulThlcslKHHV59oHe1OaSoBx7RrA
N24WyQB2VdoAzh2SwhUpufFBKDqdpIeV5TfY9Za0dHTpytEA2zMWsb90gBrFFoer
tif0grD5Rxn3VElS/Oe5HOwXwOnz8Bhshftr6dpNr1rBafA1NfxRCi8o1Se42mJw
b7FCZFwYomIQUL5quryP+95ZvNCbw18GNm/+8kLY8sBRtUc6d0mOUo7W0P775iJC
wWccjVaOH08aZ1EuPuHLH904J1pvm3D0OO9+gviLatcGSQQb6XITjKITaC838udC
cIEre5sgINTo27ZMUYs3io6n0fLjDrcD/xuccTr3ta84jZbjmggzy+NNNIALU57d
S23BcjTrDJ3J0Nmu7NIinP46r9rGGCl2pdqngmREDgilvXAqpvWlaVHQcLxrqfPm
1euH11mKUWYPYAPfV75OpjFhJD4FAsnK6x85xPkqJnmDxStyJWXH1Vr767cFQzxz
mIY4LFZH+gna6yQoSirj14GyL8A+piwKACFAV2FohXwuCNI9l5MOSN2dZPk33dkY
tYw2ykfdjofcBXorlAPFzXULTqFFcd9bdvQhztUWo/IEq89icBqwkq2fwh8uXTfu
GgcwxslxLSyg974r0nFreA==
`pragma protect end_protected

`endif
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
dlqT+cJW5DT5Gl+pbk0rOIXhgqSCJjCjiI94WWkPtMoJmIOjSfp4KqPmiI66FHYe
02QbGpBVmt7sW1NqMQM1nD3hykkDUjSKOMdW9IuxbDcstzxlGiRC4w/lpbmSRmyp
x814ss6JYCIFnAMR/n67REx0tod+6sg87VLYOpqi6y4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 556443    )
jfic22TQhd8srjpsZLnrY0MvSZp0tfxJx8PfB/pCe6oiKfwA02NCfz+lZHqA6s80
vGgmApCsmyI+Nrg3/thEZXW9Kms5axs7i85NUhDr2EKHINoyDedazt9wHTyYvOPH
`pragma protect end_protected
