
`ifndef GUARD_SVT_AXI_CACHE_SV
`define GUARD_SVT_AXI_CACHE_SV

`include "svt_axi_common_defines.svi"

`ifndef DESIGNWARE_INCDIR
  `include "svt_data.sv"
`endif

/** Add some customized logic to copy the actual memory elements */
`define SVT_AXI_CACHE_SHORTHAND_CUST_COPY \
`ifdef SVT_UVM_TECHNOLOGY \
`elsif SVT_OVM_TECHNOLOGY \
`else \
  if (do_what == DO_COPY) begin \
    svt_axi_cache_copy_hook(this.__vmm_rhs); \
  end \
`endif

/** Add some customized logic to compare the actual memory elements */
`define SVT_AXI_CACHE_SHORTHAND_CUST_COMPARE \
`ifdef SVT_UVM_TECHNOLOGY \
`elsif SVT_OVM_TECHNOLOGY \
`else \
  if (do_what == DO_COMPARE) begin \
    if (!svt_axi_cache_compare_hook(this.__vmm_rhs, this.__vmm_image)) begin \
      this.__vmm_status = 0; \
    end \
  end \
`endif

//`define _SVT_AXI_CACHE_DEBUG \
    //`ifdef SVT_AXI_TEMP_CACHE_DEBUG \
        //`svt_amba_debug(cache_name,$sformatf \
    //`endif
// ======================================================================
/**
 * This class is used to model a single cache. 
 *
 * Internally, the cache is modeled with a sparse array of svt_axi_cache_line objects,
 * each of which represents a full cache line.
 */
class svt_axi_cache extends `SVT_DATA_TYPE;

  /**
   * Convenience typedef for address properties
   */
  typedef bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr_t;
  
  /**
   * Convenience typedef for data properties
   */

  typedef bit [7:0] data_t;

  /**
    * Enum to represent the different cache structures
    * DIRECT_MAPPED: An entry corresponding to a main memory address
    * is stored in a cache line with a unique index. For example,
    * consider an 8 KB cache where the cache line size is 16 bytes
    * and there are 512 such lines. Then addresses 0, 8K, 16K, 24K etc
    * are always mapped to index 0 of the cache and so on.
    * FULLY_ASSOCIATIVE: In such a cache structure, a given main
    * memory address can be stored in a cache line with any index. 
    * TWO_WAY_ASSOCIATIVE: An entry corresponding to a main memory
    * address can be stored in any one of two cache line indices.
    * For example, consider an 8 KB cache where the cache line size
    * is 16 bytes and there are 512 such lines. These 512 lines are
    * divided into 256 sets with "2 ways" for each set. So any given
    * main memory address can be stored in only a unique set, but within
    * this set, it can be stored in one of the two ways. 
    * NOTE: Currently only FULLY_ASSOCIATIVE is supported 
    */
  typedef enum {
    FULLY_ASSOCIATIVE   = `SVT_CACHE_FULLY_ASSOCIATIVE,
    DIRECT_MAPPED       = `SVT_CACHE_DIRECT_MAPPED,
    TWO_WAY_ASSOCIATIVE = `SVT_CACHE_TWO_WAY_ASSOCIATIVE
  } cache_structure_enum;

  /** @cond PRIVATE */
  /** 
    * The minimum address in the shared region of memory
    * that the component where this cache resides in will access
    */ 
  addr_t shared_start_addr;

  /** 
    * The maximum address in the shared region of memory
    * that the component where this cache resides in will access
    */ 
  addr_t shared_end_addr;

  /** 
    * The width of each cache line in bits
    */
  int cache_line_size = 32;

  /**
    * The number of cache lines in this cache
    * The cache_line_width*num_cache_lines defaults to a 1 KB cache memory
    */
  int num_cache_lines = 256;


  /**
    * Flag to indicate CHI ICN Full-Slave mode. Set when CHI Interconnect is
    * used in Full-Slave mode.
    * Default value is 0.
    */
  bit is_chi_icn_full_slave = 0;

  /**
   * Indicates whether the cache supports storing poison fields
   */
  local bit poison_enable;

  /**
   * Indicates whether the cache supports storing data_check(parity) fields
   */
  local bit data_check_enable;

  /**
   * Poison granularity: number of data bytes corresponding to a poison bit
   */
  local int num_bytes_per_poison_bit = 8;
  
  /**
    * The structure of the cache
    */
  cache_structure_enum cache_structure = FULLY_ASSOCIATIVE;

  /**
   * Indicates whether the cache supports storing Tag value
   */
  local bit tag_enable;

  /**
   * Indicates whether the cache supports partial cache states: UCE, UDP
   */
  local bit partial_cache_states_enable =0;
  /** @endcond */

/** @cond PRIVATE */


  /**
   * Sparse array of svt_axi_cache_line objects, used to model the physical
   * storage of this cache.
   *
   * The array is to be indexed only by an expression that evaluates to an 
   * address within the bounds of the maximum number of cache lines in the cache.
   */
  local svt_axi_cache_line cache_lines [addr_t];

  /**
    * Array of addresses mapped to each index of the cache.
    * Whenever a cache line is updated, this is also updated to
    * reflect the updated contents and may be used by the various
    * cache access methods depending on the structure of the cache 
    */
  local addr_t addr_mapped_to_indices [int];

  /**
   * Sparse array used to store the number of reservations for 
   * addresses for which cache lines are reserved.
   *
   * The array is to be indexed only by an expression that evaluates to an 
   * address within the bounds of the maximum number of cache lines in the cache.
   */
  //local bit reserved_cache_lines [addr_t];
  local int reserved_cache_lines [addr_t];

  /**
    * Array of addresses mapped to a reserved index of the cache.
    */
  local addr_t addr_mapped_to_reserved_indices [int];

  /** 
    * log_base_2 of cache_line_size used for aligning
    * addresses
    */
  local int log_base_2_cache_line_size = 2;

  /**
    * Semaphore to regulate cache access. Components using this
    * cache model can use this to first get the semaphore before
    * accessing the cache. This is useful when multiple processes
    * are accessing the same cache. 
    */
  semaphore cache_access_sema;
  
  /**
    * PA writer handle which is used to write the cache data inside
    * FSDB. The data will written out only into FSDB and not for XML.
    * This means the handle is instanciated only when FSDB is enabled.
    */
  svt_xml_writer pa_writer;

  /**
    * Transaction UID
    * To support cache operation to transaction relationship 
    */
  string transaction_uid;

  /**
    * Transaction type
    * To support cache operation to transaction relationship 
    */
  string transaction_type = "";

`ifdef SVT_VMM_TECHNOLOGY
  /** Shared log object if user does not pass log object */
  local static vmm_log shared_log = new ( "svt_axi_cache", "class" );
`endif
  
  local int dbg_indx;
  local string cache_name = "";
/** @endcond */

`ifdef SVT_UVM_TECHNOLOGY
  // --------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new instance of this class.
   *
   * When this object is created, the cache is assigned an instance name, 
   * cache line size, number of cache lines, the cache structure and 
   * the minimum and maximum shared address.  
   *
   * @param name Intance name for this memory object
   * 
   * @param suite_name Name of the suite in which the memory is used.
   * 
   * @param cache_line_size The width of each cache line in bits.
   * 
   * @param num_cache_lines The number of cache lines in this cache.
   * 
   * @param cache_structure The structure of this cache.
   * 
   * @param shared_start_addr The minimum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   * 
   * @param shared_end_addr The maximum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   *        
   * @param is_chi_icn_full_slave (Optional) Applicable only in case of CHI
   * ICN Full Slave mode where it is passed as 1. Default value is 0.
   */
  extern function new(string name = "svt_transaction_inst",
                      string suite_name = "",
                      int cache_line_size = 32,
                      int num_cache_lines = 256,
                      cache_structure_enum cache_structure = FULLY_ASSOCIATIVE,
                      addr_t shared_start_addr = 0, 
                      addr_t shared_end_addr = ((1<<`SVT_AXI_MAX_ADDR_WIDTH)-1),
                      bit is_chi_icn_full_slave = 0);
`elsif SVT_OVM_TECHNOLOGY
  // --------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new instance of this class.
   *
   * When this object is created, the cache is assigned an instance name, 
   * cache line size, number of cache lines, the cache structure and 
   * the minimum and maximum shared address.  
   *
   * @param name Intance name for this memory object
   * 
   * @param suite_name Name of the suite in which the memory is used.
   * 
   * @param cache_line_size The width of each cache line in bits.
   * 
   * @param num_cache_lines The number of cache lines in this cache.
   * 
   * @param cache_structure The structure of this cache.
   * 
   * @param shared_start_addr The minimum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   * 
   * @param shared_end_addr The maximum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   *        
   * @param is_chi_icn_full_slave (Optional) Applicable only in case of CHI
   * ICN Full Slave mode where it is passed as 1. Default value is 0.
   */
  extern function new(string name = "svt_transaction_inst",
                      string suite_name = "",
                      int cache_line_size = 32,
                      int num_cache_lines = 256,
                      cache_structure_enum cache_structure = FULLY_ASSOCIATIVE,
                      addr_t shared_start_addr = 0, 
                      addr_t shared_end_addr = ((1<<`SVT_AXI_MAX_ADDR_WIDTH)-1),
                      bit is_chi_icn_full_slave = 0);
`else
  // --------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new instance of this class.
   *
   * When this object is created, the cache is assigned an instance name, 
   * cache line size, number of cache lines, the cache structure and 
   * the minimum and maximum shared address.  
   *
   * @param log The log object.
   *
   * @param suite_name Name of the suite in which the memory is used.
   * 
   * @param cache_line_size The width of each cache line in bits.
   * 
   * @param num_cache_lines The number of cache lines in this cache.
   * 
   * @param cache_structure The structure of this cache.
   * 
   * @param shared_start_addr The minimum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   * 
   * @param shared_end_addr The maximum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   *        
   * @param is_chi_icn_full_slave (Optional) Applicable only in case of CHI
   * ICN Full Slave mode where it is passed as 1. Default value is 0.
   */
`ifndef __SVDOC__
`svt_vmm_data_new(svt_axi_cache)
`endif
   extern function new(vmm_log log = null,
                      string suite_name = "",
                      int cache_line_size = 32,
                      int num_cache_lines = 256,
                      cache_structure_enum cache_structure = FULLY_ASSOCIATIVE,
                      addr_t shared_start_addr = 0, 
                      addr_t shared_end_addr = ((1<<`SVT_AXI_MAX_ADDR_WIDTH)-1),
                      bit is_chi_icn_full_slave = 0);
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
`ifndef __SVDOC__
  `svt_data_member_begin(svt_axi_cache)
    `SVT_AXI_CACHE_SHORTHAND_CUST_COPY
    `SVT_AXI_CACHE_SHORTHAND_CUST_COMPARE
  `svt_data_member_end(svt_axi_cache)
`endif

  // ---------------------------------------------------------------------------
  
  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given index.
   * If the index does not exist this function returns 0, else it returns 1.
   *
   * @param index The index of the cache line to be read.
   *
   * @param addr Assigned with the address stored in the given index. Please
   * note that if the address specified is unaligned to cache line size, an
   * aligned address is computed internally, before doing the operation.
   *
   * @param data Assigned with the data stored in the given index.
   * 
   * @param is_unique Returns 1 if the cache line at the given index is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line at the given index is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line at given index.
   * 
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   *
   * @return If the read is successful, that is, if the given index
   * has an entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_by_index(input int index,
                                            output addr_t addr, 
                                            output bit [7:0] data[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0);

  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given index.
   * If the index does not exist this function returns 0, else it returns 1.
   *
   * @param index The index of the cache line to be read.
   *
   * @param addr Assigned with the address stored in the given index. Please
   * note that if the address specified is unaligned to cache line size, an
   * aligned address is computed internally, before doing the operation.
   *
   * @param data Assigned with the data stored in the given index.
   * 
   * @param dirty_byte_flag Returns dirty flag associated with each byte in the
   * cache line associated with the given address. '1' indicates data byte is dirty
   * '0' indicates data byte id clean
   * 
   * @param is_unique Returns 1 if the cache line at the given index is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line at the given index is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line at given index.
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   * 
   * @return If the read is successful, that is, if the given index
   * has an entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_line_by_index(input int index,
                                            output addr_t addr, 
                                            output bit [7:0] data[],
                                            output bit       dirty_byte_flag[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0);

  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given address.
   * If there is no entry corresponding to this address
   * returns 0, else it returns 1.
   *
   * @param addr The address associated with the cache line that needs
   * needs to be read. Please note that if the address specified is unaligned to
   * cache line size, an aligned address is computed internally, before doing
   * the operation.
   *
   * @param index Assigned with the index of the cache line associated
   * with the given address.
   *
   * @param data Assigned with the data stored in the cache line associated
   * with the given address.
   * 
   * @param is_unique Returns 1 if the cache line for given address is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line for the given address is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line associated with
   * the given address 
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   *
   * @return If the read is successful, that is, if the given address 
   * has an associated entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_by_addr(
                                            input addr_t addr, 
                                            output int index,
                                            output bit [7:0] data[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0 );

  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given address.
   * If there is no entry corresponding to this address
   * returns 0, else it returns 1.
   *
   * @param addr The address associated with the cache line that needs
   * needs to be read. Please note that if the address specified is unaligned to
   * cache line size, an aligned address is computed internally, before doing
   * the operation.
   *
   * @param index Assigned with the index of the cache line associated
   * with the given address.
   *
   * @param data Assigned with the data stored in the cache line associated
   * with the given address.
   * 
   * @param dirty_byte_flag Returns dirty flag associated with each byte in the
   * cache line associated with the given address. '1' indicates data byte is dirty
   * '0' indicates data byte id clean
   * 
   * @param is_unique Returns 1 if the cache line for given address is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line for the given address is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line associated with
   * the given address 
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   * 
   * @return If the read is successful, that is, if the given address 
   * has an associated entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_line_by_addr(
                                            input addr_t addr, 
                                            output int index,
                                            output bit [7:0] data[],
                                            output bit       dirty_byte_flag[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0);
  // ---------------------------------------------------------------------------
  /**
   * Writes cache line information into a cache line.  If the index is a
   * positive value, the addr, data, status and age information is written in
   * the particular index. Any existing information will be overwritten. If the
   * value of index is passed as -1, the data will be written into any available
   * index based on the cache structure. If there is no available index, data is
   * not written and a failed status (0) is returned.
   *
   * @param index The index to which the cache line information needs to be
   * written. The range of index is between 0 to
   * (svt_axi_port_configuration::num_cache_lines - 1).
   * 
   * @param addr The main memory address to which the cache line is to be
   * associated. Please note that if the address specified is unaligned to cache
   * line size, an aligned address is computed internally, before doing the
   * operation. 
   * 
   * @param data The data to be written into this cache line. 
   *
   * @param byteen (Optional) The byte-enables to be applied to this write. A 1 in a
   * given bit position enables the byte in the data corresponding to that bit
   * position.
   * 
   * @param is_unique (Optional) The shared status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param is_clean (Optional) The clean status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param age (Optional) The age to be stored in the cache line. If not passed, the
   * age information is not changed/updated. Typically, current simulation clock
   * cycle can be specified as the age.
   *
   * @param retain_reservation (Optional) ensure that no existing reservation
   * which was made for some other transaction is deleted. The cache keeps
   * track of the number of reservations on each address. If this bit is 0,
   * with each write, the number of reservations on the given address is
   * decremented by 1. If there is only one reservation on this address, this
   * write will result in all reservations being deleted. If this bit is 1, no
   * reservations are decremented or deleted.
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   *
   * @return 1 if the write was successful, or 0 if it was not successful.
   */
   extern virtual function bit write(
                                     int index, 
                                     addr_t addr = 0,
                                     bit [7:0] data[],
                                     bit byteen[],
                                     int is_unique = -1,
                                     int is_clean = -1,
                                     longint age = -1,
                                     bit retain_reservation = 0,
                                     bit record_to_fsdb = 1
                               );
  // ---------------------------------------------------------------------------
  /**
   * This function writes into the cache via backdoor. Backdoor accesses are
   * direct accesses to the cache in the VIP by the user in the testbench. For
   * example, if users want to preload the cache from the testbench, this
   * function must be used. This function does not delete any existing
   * reservation made to this address by some other transaction. Reservations
   * may have been made by the master VIP for transactions to the same address
   * as what  is requested in the backdoor write. Using this function for
   * backdoor writes (as opposed to using the write() function) makes sure that
   * those reservations are not deleted.
   * 
   * If the index is a positive value, the addr, data, status and age information is written in
   * the particular index. Any existing information will be overwritten. If the
   * value of index is passed as -1, the data will be written into any available
   * index based on the cache structure. If there is no available index, data is
   * not written and a failed status (0) is returned.
   *
   * @param index The index to which the cache line information needs to be
   * written. The range of index is between 0 to
   * (svt_axi_port_configuration::num_cache_lines - 1).
   * 
   * @param addr The main memory address to which the cache line is to be
   * associated. Please note that if the address specified is unaligned to cache
   * line size, an aligned address is computed internally, before doing the
   * operation. 
   * 
   * @param data The data to be written into this cache line. 
   *
   * @param byteen (Optional) The byte-enables to be applied to this write. A 1 in a
   * given bit position enables the byte in the data corresponding to that bit
   * position.
   * 
   * @param is_unique (Optional) The shared status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param is_clean (Optional) The clean status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param age (Optional) The age to be stored in the cache line. If not passed, the
   * age information is not changed/updated. Typically, current simulation clock
   * cycle can be specified as the age.
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   *
   * @return 1 if the backdoor write was successful, or 0 if it was not successful.
   */
   extern virtual function bit backdoor_write(
                                     int index, 
                                     addr_t addr = 0,
                                     bit [7:0] data[],
                                     bit byteen[],
                                     int is_unique = -1,
                                     int is_clean = -1,
                                     longint age = -1,
                                     bit record_to_fsdb = 1
                               );
   
  // ---------------------------------------------------------------------------
  /**
   * Gets the index of a cache line corresponding to the given address
   * If there is no corresponding entry returns -1.
   *
   * @param addr The address whose index is required. 
   *
   * @return Returns the index corresponding to the given address. If
   * there is no such entry, returns -1.
   */
  extern virtual function int get_index_for_addr(
                                            input addr_t addr 
                              );
  // ---------------------------------------------------------------------------
  /**
   * Gets the address stored in the cache line at given index. 
   * If there is no corresponding entry returns -1.
   *
   * @param index The index of the cache line
   *
   * @param addr Assigned with the address stored at given index. 
   *
   * @return Returns 1 if there is a cache line at given index, else
   * returns 0. 
   */
  extern virtual function bit get_addr_at_index( input int index, 
                                            output addr_t addr 
                              );
  // ---------------------------------------------------------------------------
  /**
   * Returns the index corresponding to the least recently used cache line 
   * between the given set of indices. The least recently used cache line
   * is the cache line with the least age. 
   * @param low_index The first index at which the operation is to be done
   * @param high_index The last index at which the operation is to be done.
   * @param is_not_reserved Indicates that the entry returned should not be
   * a reserved index.
   * @return Returns the index corresponding to the least recently 
   * used cache line
   */
  extern virtual function int get_least_recently_used(
                                int low_index,
                                int high_index,
                                bit is_not_reserved = 1
                              );
  // ---------------------------------------------------------------------------
  /**
    * Invalidates the cache line entry for a given addr. This method removes the
    * cache line from the cache for the given address.
    *
    * @param addr The address that needs to be invalidated.
    *
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, if
    * there is a corresponding entry. Else, returns 0.
    */
  extern virtual function bit invalidate_addr(
                                addr_t addr,
                                bit record_to_fsdb = 1 
                              );
  // ---------------------------------------------------------------------------
  /**
    * Invalidates the cache line entry at the given index. This method removes the
    * cache line from the cache for the given index.
    *
    * @param index The index that needs to be invalidated.
    *
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, if
    * there is a corresponding entry. Else, returns 0.
    */
  extern virtual function bit invalidate_index(
                                int index,
                                bit record_to_fsdb = 1 
                              );
  // ---------------------------------------------------------------------------
  /**
   * Updates the status of the cache line for the given address.
    * Reserves the given index of the cache for future use. The get_any_index
    * function takes into account the reserved indices as well so that a user
    * is always given an index that is neither currently in use nor reserved
    * for future use. When a cache line is written into an index, the corresponding 
    * index is deleted from the set of reserved indices (if present).
    *
    * @param index The index that needs to be reserved.
    *
    * @return Returns 1 if the operation is successful, else returns 0.
    */
  extern virtual function bit reserve_index(
                                int index,
                                addr_t addr
                              );
  // ---------------------------------------------------------------------------
  /**
    * Gets the reserved index for the given addr.
    * @param addr Address for which the index needs to be found
    * @return Returns the index.
    */
  extern virtual function int get_reserved_index(addr_t addr);
  // ---------------------------------------------------------------------------
  /**
    * Deletes all reservations made in this cache for future updates in cache.
    */
  extern function void delete_reservations();
  // ---------------------------------------------------------------------------
  /**
    * Delete or decrement reserved_cache_lines corresponding to address
    */
  extern function int delete_reservation_for_addr(addr_t addr);
   
  // ---------------------------------------------------------------------------
  /**
   * Updates the status of the cache line for the given address
   *
   * @param addr The address that needs to be updated.
   *
   * @param is_unique The shared status to which the cache line associated
   * with the addres needs to be updated. 
   * A value of 1 indicates that  the corresponding cache line is not shared 
   * with other caches 
   * A value of 0 indicates that  the corresponding cache line is shared 
   * with other caches 
   * A value of -1 indicates that the current status need not be changed.
   * @param is_clean The clean status to which the cache line associated
   * with the addres needs to be updated. 
   * A value of 1 indicates that  the corresponding cache line is updated
   * relative to main memory. 
   * A value of 0 indicates that  the corresponding cache line is not 
   * updated with respect to main memory. 
   * A value of -1 indicates that the current status need not be changed.
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
   extern virtual function bit update_status(
                                addr_t addr, 
                                int is_unique,
                                int is_clean,
                                bit record_to_fsdb = 1
                           );
  // ---------------------------------------------------------------------------
  /**
   * Updates the status of the Tag held in the cache line for the given address
   *
   * @param addr The address that needs to be updated.
   *
   * @param is_invalid This specifies if the Tag is held in the cache line. 
   * A value of 1 indicates that the corresponding cache line should not contain Tags and the Tag state
   * must be considered Invalid
   * A value of 0 indicates that the corresponding cache line contains Tags
   * @param is_clean Specifies the state of the Tag held in the cache line. 
   * A value of 1 indicates that  the Tag is held in clean state. 
   * A value of 0 indicates that  the Tag is held in dirty state. 
   * . 
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
   extern virtual function bit update_tag_status(
                                addr_t addr, 
                                bit is_invalid,
                                bit is_clean,
                                bit record_to_fsdb = 1
                           );
  // ---------------------------------------------------------------------------
  /**
   * Gets the status of the cache line for the given address
   *
   * @param addr The address whose status is required.
   *
   * @param is_unique The shared status of the cache line associated
   * with the address. 
   * A value of 1 indicates that  the corresponding cache line is not shared 
   * with other caches 
   * A value of 0 indicates that  the corresponding cache line is shared 
   * with other caches 
   * @param is_clean The clean status of the cache line associated
   * with the address. 
   * A value of 1 indicates that  the corresponding cache line is updated
   * relative to main memory. 
   * A value of 0 indicates that  the corresponding cache line is not 
   * updated with respect to main memory. 
   *
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
   extern virtual function bit get_status(
                                addr_t addr, 
                                output bit is_unique,
                                output bit is_clean
                           );
  // ---------------------------------------------------------------------------
  /**
   * Updates the age of the cache line associated with the given address
   *
   * @param addr The address that needs to be updated.
   *
   * @param age  The age to which the associated cache line is to be updated.
   *
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
  extern virtual function bit update_age(
                                addr_t addr,
                                longint age
                              );
  // ---------------------------------------------------------------------------
  /**
   * Gets the age of the cache line associated with the given address
   *
   * @param addr The address whose age is required.
   *
   * @param age  Assigned with the age associated with the cache line of the address.
   *
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
  extern virtual function bit get_age(
                                addr_t addr, 
                                output longint age
                              );
  // ---------------------------------------------------------------------------
  /**
    * Sets the protection type of this address.
    * For is_privileged, is_secure and is_instruction arguments, a value of -1 indicates that the existing value
    * should not be modified. Definitions of priveleged, secure and instruction access
    * are as per AXI definitions for access permissions of AxPROT signal.
    * @param addr The address that needs to be updated.
    * @param is_privileged Indicates if the address corresponding to this line is privileged
    * @param is_secure Indicates if the address corresponding to this line is secure
    * @param is_instruction Indicates if the address corresponding to this line is an instruction
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_prot_type( addr_t addr,
                                     int is_privileged = -1,
                                     int is_secure = -1,
                                     int is_instruction = -1,
                                     bit record_to_fsdb = 1 );

  
  // ---------------------------------------------------------------------------
  /**
    * Gets the protection type of this cache line.
    * Definitions of priveleged, secure and instruction access
    * are as per AXI definitions for access permissions of AxPROT signal.
    * @param addr The address whose information needs to be retreived.
    * @param is_privileged Indicates if the address corresponding to this line is privileged
    * @param is_secure Indicates if the address corresponding to this line is secure
    * @param is_instruction Indicates if the address corresponding to this line is an instruction
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_prot_type(addr_t addr,
                                     output bit is_privileged,
                                     output bit is_secure,
                                     output bit is_instruction);

  // ---------------------------------------------------------------------------
  /**
    * Sets the memory attribute of this address 
    * Definition of memory attribute is as per AXI definition of memory attribute for AxCACHE signalling.
    * @param addr The address that needs to be updated.
    * @param cache_type Memory attribute of this cache line
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_cache_type(addr_t addr, 
                                     bit[3:0] cache_type, 
                                     bit record_to_fsdb = 1);
  // --------------------------------------------------------------------
  /**
    * Gets the memory attribute of this cache line.
    * Definition of memory attribute is as per AXI definition of memory attribute for AxCACHE signalling.
    * @param addr The address whose information needs to be retreived.
    * @param cache_type Returns the memory attribute of this cache line
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_cache_type(addr_t addr, output bit[3:0] cache_type);

  `protected
dVP.+^@f>TG);?7FcQGf+&Z;b&BM[dG4_<=DTTa7M9>?;6RTPOYC()=?>He^EFfO
ME?/+JLTBUTHW(U4Q.2-C6dKSYYZT/aF=Lg)V>)[D(66N7I&RG^)ga?@)+R0=RJ>
<4;L1DK7dZV=_WcZRaeRBHB.SJF7Zb8d/IAed.,<G[?E0&(,(7&]OgQ^3;g[]bgT
G3Z)CKc^&28T0B\[(,;\a]_117UB:P10OAKU=)Z5f-Mb3YTf7g9>97<A[/-fP7e@
Z+3XZF?)aHbYVMD#Nb(a#UQCfI5.:_=e40N5Fc80cGXgK+eGeGIDa[[[#Z_DB3FQ
27SX3EGG3D#MMML&R9V5eB=#1\PeXJ/(>HT^D=/HX^&INT,]D\@2XPY5Agg4ZTOTU$
`endprotected


  // ---------------------------------------------------------------------------
  /**
    * Sets the Tag field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store Tag settings.
    * This method must be called only when the cacheline corresponding to this address exists in the cache.
    * @param addr The address that needs to be updated.
    * @param tag Tag settings corresponding to the address.
    * @param tag_update TagUpdate settings to indicate which entries in the 'tag' array are valid.
    * @param is_invalid Tag State setting, which when set indicates that Tags must be invalidated from the cacheline correpsonding to this address.
    * If is_invalid is set to 1, tag, tag_update and is_clean values passed to the API will be ignored.
    * @param is_clean Tag State setting, which when set to 1 indicates that Tag state must be set to clean, and 
    * when set to 0, indicates that Tag state must be set to dirty. 
    * This setting is applicable only when is_invalid is set to zero.
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing Tags
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_tag( addr_t addr,
                               bit[(`SVT_AXI_NUM_BITS_IN_TAG-1):0] tag[],
                               bit tag_update[],
                               bit is_invalid,
                               bit is_clean,
                               bit record_to_fsdb = 1);
  
  
  // ---------------------------------------------------------------------------
  /**
    * Gets the Tag filed corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store Tag settings.
    * This method must be called only when the cacheline corresponding to this address exists in the cache.
    * @param addr The address whose information needs to be retreived.
    * @param tag Tag setting corresponding to this cacheline.
    * @param tag_update TagUpdate settings to indicate which entries in the 'tag' array are valid.
    * @param is_invalid Tag State setting, which when set indicates that Tags are not present in the cacheline, and the Tag state is Invalid.
    * If is_invalid is set to 1, tag, tag_update and is_clean values returned by the API must be ignored.
    * @param is_clean Tag State setting, which when set to 1 indicates that Tag state is clean, 
    * and when set to 0, indicates that Tag state is dirty. 
    * This setting is applicable only when is_invalid is set to zero.
    * @param tag_str Tag setting corresponding to this cacheline as string.
    * 
    * @return Returns 1 if the operation is successful, that is, storing Tags 
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_tag( addr_t addr,
                               output bit[(`SVT_AXI_NUM_BITS_IN_TAG-1):0] tag[],
                               output bit tag_update[],
                               output bit is_invalid,
                               output bit is_clean,
                               output string tag_str); 


  
  // ---------------------------------------------------------------------------
  /**
    * API to get poison_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_poison_enabled();
  
  // ---------------------------------------------------------------------------
  /**
    * API to get tag_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_tag_enabled();

  // ---------------------------------------------------------------------------
  /**
    * API to get partial_cache_states_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_partial_cache_states_enabled();
  
  // ---------------------------------------------------------------------------
  /**
    * Sets the poison field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store poison settings.
    * @param addr The address that needs to be updated.
    * @param poison poison settings corresponding to the address.
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing poison
   *  is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_poison( addr_t addr,
                                  bit poison[],
                                  bit record_to_fsdb = 1);
  
  // ---------------------------------------------------------------------------
  /**
    * Gets the poison filed corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store poison settings.
    * @param addr The address whose information needs to be retreived.
    * @param poison Poison setting corresponding to this address.
    * @param poison_str Poison setting corresponding to this address as string.
    * 
    *
    * @return Returns 1 if the operation is successful, that is, storing poison 
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_poison( addr_t addr,
                                  output bit poison[],
                                  output string poison_str);

   `protected
&(Acc;I83W3[;geT,56)&O[EY#\Cag^W+?>SG4[QM[,e;dT1PKIB0)C[2ZO)TZ6[
.;L/gQKYe\V_JK])T,(8&78bEOZ(>g7_-3:JCR4L.g@U8CQ15/(bM;gDfO+GFULO
e\U-2>>:+:gRTc1PK]P+cg(;IZM8eFZ,dNb8S5FXdIBE[/7a?9.42f_3@KT79M\,Q$
`endprotected

  
  // ---------------------------------------------------------------------------
  /**
    * API to get data_check_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_data_check_enabled();
  
  // ---------------------------------------------------------------------------
  /**
    * Sets the data_check field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings.
    * @param addr The address that needs to be updated.
    * @param data_check data_check settings corresponding to the address.
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing data_check
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_data_check( addr_t addr,
                                      bit data_check[],
                                      bit record_to_fsdb = 1);

  // ---------------------------------------------------------------------------
  /**
    * Sets the data_check_passed field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings. 
    * @param addr The address that needs to be updated.
    * @param data_check_passed data_check_passed settings corresponding to the address.
    *        For each of the data bytes and corresponding data_check value, 
    *        this field indicates whether the parity check has passed or not.
    * 
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing data_check
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    * 
    */
  extern function bit set_data_check_passed( addr_t addr,
                                             bit data_check_passed[],
                                             bit record_to_fsdb = 1);
  
  // ---------------------------------------------------------------------------
  /**
    * Gets the data_check filed corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings.
    * @param addr The address whose information needs to be retreived.
    * @param data_check Data_check setting corresponding to this address.
    * @param data_check Data_check setting corresponding to this address as string.
    *
    * @return Returns 1 if the operation is successful, that is, storing data_check 
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_data_check( addr_t addr,
                                      output bit data_check[],
                                      output string data_check_str);

  
  // ---------------------------------------------------------------------------
  /**
    * Gets the data_check_passed field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings. 
    * @param addr The address that needs to be updated.
    * @param data_check_passed data_check_passed settings corresponding to the address.
    *        For each of the data bytes and corresponding data_check value, 
    *        this field indicates whether the parity check has passed or not.
    * @param data_check_passed_str data_check_passed settings corresponding to the address as string.   
    * @return Returns 1 if the operation is successful, that is, storing data_check
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    * 
    */
  extern function bit get_data_check_passed( addr_t addr,
                                             output bit data_check_passed[],
                                             output string data_check_passed_str);

  // ---------------------------------------------------------------------------
  /**
   * This method allows the user to get an index in the cache which may either
   * be allocated for a cache line, or not allocated. If user specifies the
   * values of arguments is_unique and is_clean as -1, then an index is returned
   * where no cache line has been allocated. If user specifies the values of
   * arguments is_unique and is_clean as 0 or 1, index is returned where a cache
   * line is allocated, and the cache line state is as specified. The returned
   * index is between values specified by low_index and high_index.
   *
   * @param is_unique The shared status of the cache line which needs to be 
   * retreived.
   * A value of 1 indicates that  the cache line must not be shared 
   * with other caches. 
   * A value of 0 indicates that the cache line could be shared. 
   * A value of -1 indicates that the shared status of the cache line could 
   * be in any state.
   *
   * @param is_clean The clean status of the cache line that needs to be
   * retreived. 
   * A value of 1 indicates that the cache line must be updated
   * relative to main memory. 
   * A value of 0 indicates that the cache line must not be
   * updated with respect to main memory. 
   * A value of -1 indicates that the clean status of the cache line could 
   * be in any state.
   * 
   * @param low_index The first index at which the operation is to be done. 
   *
   * @param high_index The last index at which the operation is to be done. 
   *
   * @return Returns a positive integer if the operation is successful, 
   * that is, a cache line satisfying the requirements is found, 
   * otherwise returns -1.
   */
  extern virtual function int get_any_index(
                                int is_unique,
                                int is_clean,
                                int low_index,
                                int high_index        
                              );
  // ---------------------------------------------------------------------------
  /** @cond PRIVATE */
  /**
    * Loads the cache based on the contents of the file.
    * Each line of the file represents a cache line.
    * Each line should have the following format:
    * <index> <addr> <data> <shared status> <clean status> <age> 
    *
    * @param filename The full path to the file.
    *
    * @return Returns 1 if the cache was successfully loaded, else returns 0.
    */
  extern virtual function bit load_cache(string filename);
  // ---------------------------------------------------------------------------
  /**
    * Dumps the contents of the into a file.
    * Each line of the file represents a cache line.
    * Each line has the following format:
    * <index> <addr> <data> <shared status> <clean status> <age> 
    *
    * @param filename The full path to the file into which the contents of the
    * cache are to be dumped.
    *
    * @return Returns 1 if the cache was successfully saved, else returns 0.
    */
  extern virtual function bit save_cache(string filename);

  /** @endcond */
  // ---------------------------------------------------------------------------
  /** 
   * Get matched tagged address of cache lines with is_unique, is_clean settings
   * @param is_unique is_unique setting that is required to match for the cache lines.
   * - When set to a value >= 1: considered as 1
   * - When set to a value <= -1: considered as don't care
   * .
   * @param is_clean is_clean setting that is required to match for the cache lines
   * - When set to a value >= 1: considered as 1
   * - When set to a value <= -1: considered as don't care
   * .
   * @param matched_tagged_addr queue of tagged addresses with matched is_uquie, is_clean settings
   * @return Returns 1 if there are any cache lines found with matching input arguments
   */
  extern virtual function bit get_tagged_addresses_for_matched_cache_state(input int is_unique,
                                                                           input int is_clean,
                                                                           output    addr_t matched_tagged_addr[$]);
  
  // ---------------------------------------------------------------------------
  /**
   * Clears the contents of the cache.
   */
  extern virtual function void invalidate_all();

  // ---------------------------------------------------------------------------
  /**
   * Returns the class name for the object.
   */
  extern virtual function string get_mcd_class_name();

  // ---------------------------------------------------------------------------
  /**
   * Returns the cacheline stored in the specified address. 
   * If there is no such cacheline a null is returned
   */
  extern virtual function svt_axi_cache_line get_cache_line(addr_t addr);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM display routine to display the memory contents */
  extern virtual function void do_print(uvm_printer printer);

  /** Extend the UVM copy routine to compare the memory contents */
  extern virtual function void do_copy(uvm_object  rhs);

  /** Extend the UVM compare routine to compare the memory contents */
  extern virtual function bit do_compare(uvm_object rhs, uvm_comparer comparer);

`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the OVM display routine to display the memory contents */
  extern virtual function void do_print(ovm_printer printer);

  /** Extend the OVM copy routine to compare the memory contents */
  extern virtual function void do_copy(ovm_object  rhs);

  /** Extend the OVM compare routine to compare the memory contents */
  extern virtual function bit do_compare(ovm_object rhs, ovm_comparer comparer);

`else
  // ---------------------------------------------------------------------------
  /** Override the default VMM allocate implementation */
  extern virtual function vmm_data do_allocate();

  // ---------------------------------------------------------------------------
  /** Enable the VMM compare hook method */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  // ---------------------------------------------------------------------------
  /**
   * Hook called by the VMM shorthand macro after performing the automated 'copy'
   * routine.
   * 
   * @param to Destination class for teh copy operation
   */
  extern function void svt_axi_cache_copy_hook(vmm_data to = null);

  // ---------------------------------------------------------------------------
  /**
   * Hook called by the VMM shorthand macro after performing the automated
   * 'compare' routine.
   *
   * @param to vmm_data object to be compared against.
   * 
   * @param diff String indicating the differences between this and to.
   */
  extern virtual function bit svt_axi_cache_compare_hook(vmm_data to, output string diff);

  // ---------------------------------------------------------------------------
  /**
   * Hook called after the automated display routine finishes.  This is extended by
   * this class to format a display of the memory contents.
   *
   * @param prefix Prefix appended to the display
   */
  extern virtual function string svt_shorthand_psdisplay_hook(string prefix);
`endif

  /** Added to support the svt_shorthand_psdisplay method */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);

  /** Added t support the svt_shorthand_psdisplay_method*/
  extern virtual function svt_pattern allocate_pattern();
 
  /** @cond PRIVATE */
  /** Gets the address aligned to cache line size */
  extern function addr_t get_aligned_addr(addr_t addr);
  /** @endcond */
  
  //----------------------------------------------------------------------------
  /**
   * Sets the 'pa_writer' required for writing the cache data into FSDB.
   * Also this function records the meta data required for cache visualization
   * in Protocol Analyzer. 
   *
   * @param pa_writer handle to 'SVT_XML_WRITER'
   */
   extern function void set_pa_writer(svt_xml_writer pa_writer);

  //----------------------------------------------------------------------------
  /**
   * Sets the transaction uid for cache operation
   * To support cache operation to transaction relationship 
   */
   extern function void set_transaction_uid(string uid);
  
  //----------------------------------------------------------------------------
  /**
   * Sets the transaction type for cache operation
   * To support cache operation to transaction relationship 
   */
   extern function void set_transaction_type(string xact_type);

  //----------------------------------------------------------------------------
   /** Indicates if the cache line is in partial dirty state 
   *  @param addr Input address
   *  @param is_aligned_addr Indicates if the input address passed is already aligned to cache line size 
   */
  extern virtual function bit is_partial_dirty_line(input addr_t addr, input bit is_aligned_addr = 1);

  //--------------------------------------------------------------------------------
   /** Indicates if the cache line is in empty state
    * This API will return a value 1, when the cache line is in UCE state  i.e. both when is_unique and is_clean are set to 1
    * but none of the data bytes are valid.
    * @param addr Input address
    */
  extern function bit is_line_empty(input addr_t addr);
// ======================================================================
endclass

`protected
2d+&U2GPbGVZR+ONEUA3K>5-edFI[ZLd,N>LQN/YbA=82?(XM-\03)Dc3]0=AgFI
>CUa[Xa/6@F@Xf36[\NdB)D51A\a>&75-a__GB5e)gU09LI9@&QV&6-E4_f.G-Fa
BXCF;(J/3I)#T]FI]EYMf1[1CDY308V+ONGafg_JOOOfJ5REX;:Xa:Q:Y/7P)GX+
/>+)J[PI[=45JDRa;+=-I><E8(:/dL4UO5=f(T&K&WWD^>F)3(a^)KacAIWFAJ^^
f1@.edF=bPH)4K81[1K9b\P42cH.N/]1YeI/<FWE?X;2TAN#HV2IY5=D4AJE2bAM
+G=CZdXKC.bO^8K8-JU-OJ]>9Z^U9;#9f2]LI].VdYHEQGWg<Nf35?I:5?:b7,5]
bBE[_2Cc5CP>46F,WfRHM7ZSe9RNFL@M0:8gKfBAcGXQM)5dQb9+F9B/a.(9fgG7
=\,\79(EaZ8\.<FECeR)b5_TYd8/E<9)/Hf)_5C7#BAKGR)_,a7I60P+QSS:I#6b
TNeM5MH2[9;JKP[YeOHU>38.23Fb@=S40-<U=<OcF66\[7gK4T&5VD(=2<Q3I:YX
4I@^4#_^2a3C5J_[7dP+L^YFZ6QTfUbB]aH?e#-P>)WC/.>HTUN[AE,(6S:S8;LR
A;C4D7D8e7]2g<-VfYG9(4\,Zab:&OX/Oe1[-R7e??,9]b[Q3XZ,.HY06;6TB7N_
JJ4?dgF#N)07OC.MAeTcWQDBeMK[Xg]L,Z7aO2IY0]J<>D;R@41b=bNX\/&H?72S
+Sb6<f?c>8SbSCb73/9-(L^9SMeHB>DLM/]7^DSWGQe@H(FGe[L[EP&Qd-&=ZWP)
]Z51QC&GB=gV]Q6Ea>,L@/1d]K.W>]D^dL&gBGdZ:[^[5T]2Q=#G</K8D3.GI.GY
25eGc>Igb8L<QA8?_YUbXd]e\Z/gd<ZN,UgSLHBFg2(5UUGNY?d0PG,,&:9L4cTE
a22Sb^C=V0YO(<28e=Kd8Ya5I8._4Uf8JCDJI)):<\+PC;D(=UgJb((a&O;(,Gb&
(]Ee;<K4d)fKJHS8=5fD;(/g=OYJ;&XY.6>f84I.;1,7H[+-2-XL<#6N,I(]f6JO
J4aC5e,_U\e0Y3-ecTBBLH6D>eVYb_,&/EEO?#Y>C^BP,)Q):X@[Z=3P;@./<S[)
M6<EJA&c]1:6,81TNF#MC)E)PY]0DCfZF&)E0TTT=0W0UedDS:PQcPB0Nb4cTWN;
#(5EIFA3^LA3H5>b(EL</KN+:0M6IMVL(gab1@[7b6,077f-1MKQ<-Y3(/7=\_#e
DdA4?)fM>;YS^Z2?9Je0908[N_K2H@E+?OREHUb;GBM05D)HFU:g/S\R1.^X-A-M
F^C^bCCW@<,3(L9TO#/ZV/[?UU3DBEJ4#FUW;9ER?Lg]-J0S^B9DD9B/9eAV[BbK
.Xgd@9+?==534VA(f5Y=bBe6W;;^-93PTAF[:@a;4[II8Q_.U17M\Y=Pe1;/d8ag
,d8dRM&_;?dg_A\N7FA9[_S+Y;,aeON#d4_]S48cg0\;8QC1BX>Tc)7M]H3;;B?2
P5T024bA&@U3ET4IM:fZa_H67QEZ\)aV6>B7CBA9Ta[JT+(=JV^56&OV(GW=;RB4
7EWZQcZgM3XPT^aRIA-6J3_B_dUQOc36d4O-&2:g.QS&2E;eD<:d8.:Oc?I]cCWP
\2+(IL:U>S0KfbgUKQBEZ;(?UdXXV/<#e]0J_B8]B+O^d2b0OQMH^SS,Fe?NTK0+
N;@V781e76-f8)V9((FDW.Ye._=C4AMA329PGAV(XN9]@(LCV@R(,eXETLN;>O[Q
_KQ+;Vge9DAU&O>-QdNXeP#0USH2/45(DI>?>M_)>8aDgPD/F^UU1^?9OFdP/:JC
PGF>FNgAP/,73F?_(=H#bQN4TQIAAWXU,-,Q>A81,-_<2dYI2^JM_OMcJe@07T7b
4RG2Z5D6GF6UZ69A:bDWL(D<CcG1;BF@;g8:4G8I6,8,7F4:W\Q_O<]B#.SV:AT:
@J2gUDeF2)7IE/0IaYK=9=.QF&e0(^K4cXd]W5Wa;2XVeI6[c&L6=fC98;XWdO1b
OG(LJgY4_DO71)-&7bRURRC=H^#gOW;^c9D[a;3=Z)@28G/27ESW69DdSOOX6L\:
(H29)J9LYa5g/^?B\S@09#&F,<Z32]f]L:680gb8ZSJ5K_08&dDQfeNDT1ceD)J1
#,F/KZb=d?1\02@;[601QdJd9>H,^:#g?fOd3M?LD_d12AcI0V7EVBAU@8Ja_E[>
7Be9:_K8^GX@9U0;8.7_YEPecU\@KJOKTP==CS-S?]&b?_.=e&^7F;8;c[FdLV@[
_fe#=L4I,1T^LQ:F5\,JZf8_W0<dM?M3b9ZH1<IFR37?U71ZFAR^8@Y6W47#I&JK
:N7XN[#J3GY6fPITHO)MEW-d\.LU()Ed&\c7:?PRVV95ZaBC@K4aJ=\37gB]].6f
1L45I>C8//2W(-e0:;Qf=cfJFgPe-/gH6-dIVC8T4b-QH,<^3dD/X7S9,(e..NTd
0-X(FZ@Y^gc,Pc[LHS<#CE<b@A/4/W5b(E2JPGKOZF<Z7?E2L<2\?P3UWX-GX,WQ
W,J\TKRcSM&Q]OGK27V3K[JdXV]f4M9Bb&NAN8\bQZb#4&NE3f=dRb6;I8S]d3GL
4=0>a=UNZD.d]COF_H<+gB_=OA(b;Vg:FZC1I6f)1/.f2E16PW5,FMA/.6]JL:B2
WUE<)7P:+H#P[6]fH6^7?R?U9DX+/\KH1KZL4WR4HXdF=5\,FA\KEK6;,?C<-RDU
(:@6JRgQcH>.N5aY+34_CA^66d@df#OQ-#fGIbFO\gaLK-#DF6#.b<Y>Sg>#^;+=
(G@bQ2J/G,-c\9J.O@PNT@V08gNA4f9N;8)_B/Z=WF>Q\NOba_d19^UdcG#](-#e
(4dfO\SJ?_/DgaeTEB1AC<7^YOJZ.#(D/<+H?OI[-YQL<f43]a36?R[F_RH5/83-
dEE]<YW\@I<BX)0g]YQVGXdRAR:9d@Z@9eagI7H,Q+;d9LRe.:@Q6g><6?LXQCLV
g6U0?@:+NgBHPVc5RSeT&GPPYJOPNE:aVWGcMH^ITIP_CH33M4ASOVD0M)+5LgZL
;JD6Q:\@aQQXBNBUQV)JKK3DfQ,RQ8+Og;fX2HMagZVX09--R]\eB;?-;VHTQ[[B
U6I-=)Q/_&<WA)(YN-(_-YYH_b0[80WW7cANaG]g1c-2Z09egW0d;Z@g)1))f:&E
MB4@>>X6V(1#[3#4YE@TcabX_e/_K:]]2YbGGM8Z#\GOLeaPGM\cTU0GE7N.W7I>
DJ>2-c?Z1AUc9gIN<^-PW^(T?0?I[-(>7JNR1.8a<Y91V^K-K^YH08]:K;c-Ra+>
5?L067P>Q#(Y^;RX]V2_^2.M[STYZ/+?a.Dg&?U.DA5Z]Y7=Df,FIXG)=;G4.X=B
R=NC[X3(PQ?QXT4#87D5#LK1OM\]<SP0-]2]K6)<(U@7?fOg/fMD\)]d@Jc,?cU8
bB-ZbDD&)/?TT(K/(;01^ZH\G2DB1DTcU5bC^Yc(LU\=+:6QdMT\R6.4fLcX^7([
B+eaP,7^RUfggL5Z\+:gT_:-/ML:ZZ8ZggN4#3(5.bH<J2=I78A-E>_HC.SG(^ZP
Wa@Wd8aKcc)NeHQUe_IINC/a15UI)U]4]R/efa8\;?),WN/^Cb?X:NCK9fL.PfUV
HU@c+Q3L#e@@O4+E&.?=^LIE9,?g.)9R1+6TX><bL]aG&]OTFEXL]\f#F.?QL/JE
F=9J-:TAU-8^?PG.=6U]>XIE7$
`endprotected


// ----------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
CQ+4fSaQ,G\ag+>((]W?fQV?\K3XW#A3K\6:115XYQc9bfaW0(C@,(?DK-426D\a
V71(a)(ARXfcA_&LgG(YV_F29<GBfDf)&IVc=eT1;:,TOZ#,;Y;1:G;G^a:6T1EF
-(IR<86Tb)-5<F0N0W22Nb6JR\]?T_@d(I)0(KYJ;NeSS.0_YVGG189F<]75K=c)
3d(8K(5g:MD?/aUI]5YcDWB2E;EDR0MJag33dC_SHHKM?<AW(MM77eDE#41bKP/^
EM88<&.FBG8?-$
`endprotected


`ifdef SVT_UVM_TECHNOLOGY
//vcs_lic_vip_protect
  `protected
7A5ScWRVA7bSEg4_aW]/d#GbM6S6X;XM8W]X.b8L>Z3Ef0Z+LUKD((7DO\e8<b]W
cYM96EQ&]#>:\.O+VXY(7aKW7JeN/Mf\PS57fN+a(G:/#_W2E)TDMCZ]0I<5Zc:X
,3Af>Vaf\gZ;Ob+^d=4dVW6dff00TC2gRAVG/#43I21b?6NW7Tf96Y_:CLYZ-I7J
JQ+:7b0d^72?:G2c(B[PAd4UA=5-S2P0f6=@@.N3,_e2YdP4<f+?WAN=H?f.dB59
FXM#c9g(^e--ZaLSQ@CBI,>T08Z7_ZWgYN_GGT,#0BZME0PNZ:WS@O]A>C)L)2b7
,)SS?U9GfA094\,D55N+Q)5JKG86SDS5&B8A>]F6/)RAN7^;1a0R1Df<D]9?a3L2
=9]X.&L/:YcIT5_d+e<GUFO5Z8\:LP,QA+3dOFEec0O19L64\Wb6=,D04a2Ac&;^
FTH-D9LKZ7<WIH]R<1D\R7TG(8+<H/E:72TOcd+SJ71,(HIP)1RV=,5@9\T-)[g5
JD5IN024Y@+Ea]6VXJdc&XH5/O4a?4&MLX7D6,NCH7T\EPW?#<-1J5S3M<?&0/AM
X.?#^LV0G70Ma8ME8\7M\5>UZg3a2d>,A-AeXUa.DPEAT8+R?LGdB+\+S9_;LeB=
.VRZ+47g?WO#:D@Ab[2<\2[7DeZT(2U550f6Z:OTU-[FA4]@T3?(gX,^Z4T0Ud;M
)&VbCOgAP7\8E)ORRC-[[?:8AgH5+1=^f-+@XP\[8GbHXV8&HJfSFHgf-gU(6)#U
_[8L:Q1)]N5B2??KI,@ZI,-Y=WV)&IIM=D?KH0M??9R8B6I;JGP)B=A@].\dX24?
d])\0,FSe-MB3Y^:,\a]3bd]KSHUG)fc_<B+aN+WX8=P?]//WM[^:O).90ETBT5e
a=9gUaW^K95#CgTGfY)>DYRN/K&;>#.RO88aM\J#=)^^X;-H4@\QLB8[Z-6dPUP&
O/A,La1-9/MZ#-T4gI0;DI07^:GH>\g/Z[2G;L79_G5K6U0K<\MJNBYab_,]O/f8
84R_J2#>[f#X/g/FEAK6]g:#N)#-\>e>5(>bJ:0VdcS#J3/#1,bU@Je^1SNU/450
6:6dVZ.J@XCHa:9[)>gFD:5,3+(/cY)[K_4EHVX3P/2IYTGRQ_MCE@_;F_:VOfeW
[55DK.).[XMFSC6(FCV=b5HdA-#J48aWgS,c2,dW[-e>0aSBfM2:(#0#/A[V+W(B
;aF[,G2,T=A:D/S@af(,f<_d^a(M0cYgC:HJNR118a/.[>#dfNdQ5+JR^Z/8>&D4
g29(eYMO^F[-28I2EHTM(RDP7/B+NIE_QR<TFQT00C5FKbfQJ?>;RJRH-QFL^EV<
V1,,H,T=c2.(H&[F61f7HWM6#a2L+F1d.1)A_5#&bSc7Wdb8?AedeQIN]7N;b+(Y
I_Uc-/WREOT_^AVMb+DJ26S,#GI,MKg9fZdBB^ZV^)&X_]N+f]14cC/+QN]2LDab
3^)ALEa0[E[UEOV=LHDaW^Ie1WMRIYNI/,1ODKUG:XYEB.W2Q89UbT(0G=JY[W]\
5MHKePZG<KGEe.b@\Q3]N3g.0(c=gAB.7QDf&VHBZ)C2.</#d5_/@#=CVYa[a.46
0F8_T3&1d#24HE+Y01--&@NPAg<OIU1.GT.YZ.K[YEfAW_3=LS,:aKT27^B_?V8A
^/d;BN1QCE-2eFZEO(N&@32f75QVc0[(C]IZRIQ3V#.P?=+NBUeGG\fc.f&PD1b\
Z92R]HM8.@-dBT91^@f^d,L85Z]1N]C,@20IU7\U=+;(1>LHbc&,-L#/,BN+>^&]
f?7@a<L]5-(N0Q:BQN0J.@XX6L?&A,:G:\f5c2HC5_c=CORNA-a65M_6JH_.a2d[
MT\KJP2D\9L@V6^ID]3JHT_aMK4LcMb[6HH5/YAOgON^gS?WIKbY&T53)ZeYg;.E
D5?PXP;2X)WUJWe^1D7MH[N;Q_2)=&O10_&LAF1X+OP_aa/b&5#d8FB,RJ]b<WEO
)O#7g:WcLY:KFA-Z-^)AT?=TRR\:MO<-ab#fH^4P?(HK>;DPgV:.VS=Kd)\<ZH\(
D0&gMJ.\2#DKa+M/J2,L?V:<cY7-R-<WF:CZYZ?I)M-J;I^e/<ES7Z3B\SZX+.--
6@./(#]O&TZSYPGDEANW3)/R.=]Ge@fI2:ae)fK4678FgL6^d\2GUMAH8V0_SSN-
a#bVN:[;HK#FS];dOWV3be-=+>U4B5[7_CV3AH8I&FNL9;90HMQ(OcTDG4<6T)FM
@BKBC.gW5SRBU:,;6DYC;JNE=:V4W<(ba#?VB/?N4OUbM_RX2](B5SHFX)ZDM=cX
ab2b=aQ/EV1?R4MPEGB2<<\1EPM]ZTN2/I+C<+E_-FeFeE,CD:PJ.\CI<^9/HCK-
N78K2L+-WRJENW>B9Ge0-C],=;P:d:1R1PM]^6[bYDTOZeIS;4H.505Ja@224.bR
4E@NdHOgd:Q01_M]Ue)^FW0BL]V(0U.[XA[P:]JX3d4^-.C4Q;1J4\?J9KJXNeJC
gZ52],Z=>9ZYESMg]ed\>1,ZN?KFEcfI<&_/__g9P2:aHN\L^e>Ffa<\\/#)P2K8
7V9=\_(3#SHM:2FO)bY&QAE6-N.:,f^aU-LBO&-Y,_J#JMNa)ZSCR]GNIHQ2K]]+
+J#QK03ML#&af>\_Ib/H&f]=HEJ=V-,5.fde.G=FEL&3P0HDDOgU\f.5??NJ[;U\
8\9g&K\&:6.?<+KVfDeYL,;,R5&?(a)&6B6U/[(GSQ1KV0F>T-U\[OBSLEO5A(F&
Yb]OMA:V/?C.H(FK+gNe[,Q8[X+14^[EbB-_W^J45:L\)e9_@E@c7B4?c\NK7CM2
8,,G>>_SZ5e2U&,dJD0P4#,8b_0,;-WV.#>Qd2)NET4(J]Z,>)=6(3E795Q=5d:B
#W+])-1eI5<_63K;OcX+T;,87$
`endprotected
    
    `protected
c4/O]_H:A#LfE<d6g_V8>[L\;g_+?6\9CQO6IaJ,@P,&&(:g.OR>5)6C-?.1#N#U
Fda(D0<DP(VW-1()SL.:^DL\7$
`endprotected

//vcs_lic_vip_protect
  `protected
<aT(-..HQ#Hf#dMGA(5\K-60/I@+XfI99A_>0JD6X6KUWX7E&,8]+(dB7MbNSA(\
Cd2)PK>:O,7D]AKc^2?QTB5Gc\]X_45780<[6=#Y12M]MYBXI50]a77D8cJ938;5
4C#]^Wa_@(1Q_cJda4.f8A>HXIV2+#X63Pe]/5)SHd,.YPDM04?CS86c9?4e?26T
V_b)6.;QRFbC/L@ZeEXJB9;:IJ-9gJTQC5BVK_DWQI0W<^MVa\@bK2RWT3e<.6T#
T=FL;T8M_5c@OHGNL;ZS&U_9?#EIHUP(WP[+&X5Y[?CIL19Heg(5/MDI=L>B[Ta[
X^@@EI5E+1J/^._;e95Yg;R+EUf?&HXEgE8E5gR@Lg((&.fOXA0I2bE5TH\7X@92
1ZN?>OI=Q6S:+<Q2AQ7Lf:5T.5<2]bUC13C)C5MRJR;XR.XB.G:P/0BaeL&d5TH<
?/cAe]?;CBEe25?/[Nd>O1.FUVbbN)9_CgT+f3CC<F<J/PAZ,GX4GF9)1EeZ0;)U
Y;>P6dWT/+DDDS[VMORL<RQ,=1#B8DYF:_5O15]4#BOSOV]E-^RaBE2>DM2<GKII
_(TML&]+C]99a-Mc)cXXG_F6(W)#6VC9dF,^3,TY4W1SF$
`endprotected
    

`elsif SVT_OVM_TECHNOLOGY
//vcs_lic_vip_protect
  `protected
(eA1=2BfRF,JP1@gM?O\bB@.KKH-Z?N(5Z2b-@KbR4CeX.,JFLaD+(K.(MaU)@<-
-/57e.E_NS<HH[RHAHBNAfL2&5GXG/&I&0ZXK(,=IXF4=^&ZN+TS.O+7^)0-CWD>
]>g?A?YCH;OH>PF[QRXb[O#R=PaeA4Wa\ZZ5F,BR2eY)d7&+1?gcJ<JDB4#UVdCI
N:d.2EO>ND7c]e,I:L,9Z-dA_fO^#FDcPS#5@-3\PHO:47>M@TC\c>9]O#dGA)cY
FcPbZ9BV^SHT[Z7aHE;H>f-XNP-=:LY5E(.JL_-R2V_CON3]9HUP5]g8INF6.]OC
;QHYSUV,OL05GWcFV=&BF-T]Q\?XV)FW3D-#^,dbSRU.^/?D^.KQO;1DP-^&0M5E
_HfaQ)?_QZB;GJ/9OQg&ZM1KbXM7@bC-<O)3g#5?185f;V(/0HG#^7dR^S&UG<Gb
-GZ>W:L9d@<>4R_M0Wb,O:F:Y]]Q\VXO<9-fC,.IH=@(-_[KV943aP)NLb66Z1Z0
#56+/91Rb3HNJG<:Xb0W2S=_R.Eg9\\dOBUEdLR.C?&J_4<&5QD<V9G054JS3,:_
Y0HK(2fR1ZJX/YO1cQ_OO[),_Fb\)ZV_PQdS<HZ8.H3d+5+64V(<Y_IA7>QL+ZS4
ZH1_A;3bG]Ve/S(V3D840V@#dP_98P2WK_TU1AZ0a00=0J^BI,;89CQ9gLRb4JDB
E5:0/2#d4U[(N/g1M@9://_@ae2(^\_ICf3Q?^/Ha26,]5Ob/D_2C1G3)D]6BR=<
G8Ke9.C]JCY1=]NCJU&6.&0:0DTK1eQD2Q3<ZR_0J3:4B\/^41L87ISY6/D;V1Z9
TI[@NSe&\>PX?Xd^_C;^<f6OVH[P26AKB-\3+8[>f8bL\XdZ+c.Ld4IgDE@]HT^e
F#_S<0g9F20_g[+]DBIPV-g;014?O06V-6C0OB8LX?BMc2)F4:I>X=dOL^JdG@&7
[FKRMBDRaDR.Ae?@;6+Ag>B>1[V/]S/9B7,A9WCW\U=KK]P11Y\S9U-B:SD[e=O5
\J_28[He@^+EM&TF/SQ5]\N@]Qc<c4&E3:,WJ3_;f8fd=:YLAQ1YT,^5UeIc0NM7
5XSTCI],dQ<[,&O;@8I5SDTC92^1&\U2QJLV30J-8597J2JJ,.UME2QbV(^H9/11
f)Y9^ZN6Fd=Md,^-&6L2e9(PP4[65HD4R@K(@a\:c@#/<c=Q7O/8T[VR>67a/E02
V(9:WM21Q=QNg1,K?Q@J.c&b>7V<A3/(:/..QRO,XF@]MMeH2a^V0^\_W,ZBbKC3
0(5(VWZP(Q/S2]KTZ684P[]2(>P<<.;L[BHNN#D9MC8W>_49J?##A(a4DV@Wd;G@
]U2W3.27E1^\6)4GLW-6EHQ,MKf-Z3g]#?A;P40@K348KA/H?#S0]4VUS9WQ<cO>
@14,2:/T>ZW\#1L5^aT1+6.)4_-+fBM&</;#1E[N?L#Y@H]c33PR8?.&-K9Qg\TD
,-&WfDH4[1.^gK=L[K-6[fR(/1EVWE&69\6[TS4B5ZP]YB]e+YE[WK+MJE;]<GI/
V15>eK@,A\gV3F6LT>+PO)L4GNL@#T\WYYIO><)9[BC9;JLd,3>HWDDc)XHFH\P6
5Dd[)RT1G3b[TQDag,4?)/^_:KcPf3?dM1R9PZd<4?eP[d/F9.:QD_LT>PPDRAO[
HFc<]\0cc4R2R75KcIEB&]C\^39X1<LM/\VfQWB<S2SEY\W15,Bb?H4UdA]:FGBV
^YSGE@<AR>?<efbGgRLS-<P4?Y@\8]1G]2MIO.+Bae0P.Q:9\FM(ba5VM;X[+f.Y
3OLIX>KP\+[Z=g-LZeb#VI9>FWZOG[G2]\#G\LW;1A#88BKMA<91@//_9B.[MABG
U)8RNLP<VPf.71-=998NfYD:S(gV<06W<79IB[,SGXaC+d(Bc^<f<ZQ#gJU,e#7N
>TUa>IH1P;dA/b9bE/F:gQ>L)>TCFHHaZ-QB#8edPZY_^LM,;/=fQO##T#3LeEWS
9f)(]:]fV^D0fZa]?25:]BR-JCTL0CS(#A)\@LQe8P#U@eQO?YCZLJAFV.ReNW7[
Gb]H5NS;\Pe4@d5=T3]D-5P^;cC-@\]@XV;(.,VS_+6_9-A,<Q1]0;<]UFUa(SF8
UU>W\BXWEf^_W@S7@bMbX?(6,UWEJcT^.-]cT>]9+dYYR.Xaf:g-McVID1@&IUVV
+T]KD>FTgS_5()2c6?^Hd<PSS?;KE<GCU/=bQ)Y0[R5c,JfBe\)JgcUM:D7JCKZ\
B/_WARaNN^Q5^3TP2&J4PKgc4=7]29ZSH-Gfd7:>5@g@O108+XWO92-?2?3&P?NK
aZAPB&0^F4f_].5=JM7:N/59@;2#I0-CgW@/_>,D:GOG9VI1,DF#<XUU>6_Ngf>e
?FHO4+3S>(+b>,FbadW#XG-#QA7@(REdXHR2K6b0\ZXZQNgTD6^+[\Xb2Gf#Uda]
;52]\JWNRc:,\=R]+aR5=:@9>U]&6):I>:[fO8W2\7ZC_U[+Y&:3cU(SA2eMIPeG
O2R&<I9FUST7aS^(P@@aa^38G[2U4agOX;4(.GEJ60fT1S5@(cc0+SHGOV26;V]Y
XECANed8]=_AN:7#d9;DF\)Z3N-[d3>^R3dId/C#a^F[4A(\6CMH8[]1X607G-#E
VO.1<(+78Nc9)/^-Ib-#Z4HB\&QKAM1gHU=1\)\-bNA#8-Ldb]JA6\#4ZP(R>S+;
0ge.O<2QU@.SC:d.+RU483Y7IZ+-XOF;bg0Ag.0g49bH0^0;a]4;C5[^GQ&_M(fZ
d3)\5T?_N_].f5e6A=8R@_g(67]+_W9S:8DWL@D.E,U<Q4WSWIYacC.YFG-N[[\2
ga\:X^[Z5L/P61E6;Z20B4=??TDMY/^REO/D,G#FAW(>?\CJ,[<G@KB=+bPQgWSR
eH+^&cSO4(Y.G93Ug2O7cAKbIT(dYdcV3YR=#^Y3f+5@CK]Cd?F9VJZg44:=;_(C
?W3Ib5eRLQe7GdFP9Ce@.[\?Z_SQQeXJP0D72A_/Y:8_K>R\G?dF1B0K7FM^6\_:
6V/AN9J95N?[IQb@@7-GUK(.e0#92DL-,f?Q/K<=9_]@T3])Hg3S,0QIUMWWea(Q
T(@.U7RPScebFQ:JaPXc0M?./e=6CN7fBe2JXSK4T:YQM..ZC<c;D6;8Z_7KR96)
>\H60EP&JdcG>]H9.XH=Tg3+0X)GX<VDFT1c1;Ka=1#ScEGIS.+S5KeJ]e-]1L3]
H)IFU,^T[:]M5ES@1O/EI)+:B.7,D&6S;.]4e?@-Ig@CAb_/F]geWM?ZJfg+e=<+
4DI9^(BO)e@8PWAZ-]0>8)JW_Ta<4.A([7&gfK/N<Mf,S)3K-N>5gBKV_JaO(S.2
.ZKE>@++cAO?<[-K:OD;dSJe3G^[PU6:=QRBG4/\&ZPVNe[I_BRLZM?570MT4VE9
A#5UX-03LYZW=N_G<UY-M;:-RCRVdW6X/(A)L+>41@1aH#(-If]=VX1F8FRJN5c1
9X?U_Z7A@\]W0$
`endprotected


`else
//vcs_lic_vip_protect
  `protected
3bN_.5dSIX(<<D>^]=Ib9W#H-Ocb^<IEQC->C/EP54=<L^feYdDT6(@gR)VHCcE@
ZSWD@,])@ST8eg\:E)([SE5G^Je7gMNd)&AVVJ7,B>);VJ1gGO\.IAe@(]ONJJ>0
=Z5K</H,<[:YIPHdVXb_M_HJeZ&>SO;^9=&EHceNLc6,#Id[P36HC//gWT2CL;5g
B42CBNB_ZgdL>>?W93Q7;KI(>)NQE.6f]Q<28RV5_;A0:,+6OIXPbT-8A).EI;72
\/=,-P_Q35da6b?1_EJ8J<(B3H,F(A6YW0,+UFP6,>=F:Z,Ba,+CZK+7)5(^@^?c
68QH_&71#Y\/G[OAF1RX>RXSg]U(Y]-F8b9.bB+BCU<A[.T3,?O)e3g3,<a;4SWP
;2R<5YTM1@(8:DWI>>-B+1.D46e<2X<+72Cb,f&O(B@=M)+63.=gP#7T3GGN.fM,
^F=8ReRJR/QK,(2fU-07dD,67J9KfFP022#?:KYSC2^#ZVNcf3aR<A9JHaPcWP@&
NE5\Y)>[_XJ.\abT7W.b?.7NBJXZW@cD@Z)_SZ^IO4^503?RXc)R)VT_a;OF/&;8
SU_05K1]75&cW?IX3gJd9;=+=D#N_^9AN;<4@;?6#ZDd3V9Y6P[?F-8[@WX#?,NI
Le;C5=&8[30FaB/#-7KX?-5>gAF#Z_Wa42_b?;.Z<TbMD]4?VBd(NAXAe=M&U<(]
TY<b-YC61XBH1bef51A;UP5(Pa>eF>=QHR@#ff13B9_^HJ;VFQba?S8._D\:d++Z
.DJ0fRRV(?<7NT-,S>(][?K147gAZZ(:LCUeeXT<5JF/UPQL6N?NM<W=E-=J>+QX
J5K&L_Q;E\.?0UHY38RS,#,DP,JW+;@]=&I>NI:6Z#c.N@M740?4Z(BaS/+\b+fV
>cEIea,?\@g:J8#YM]Z^3cDRQ1K9410TG^WfCNc/VEOG0+#4+#?LVD(abLQF-R4b
4BH7XgP580+Q@J,Q60,e5GT3?EOe5.PfbTcE\eBaf@#E&CKaWU)O9R9QFL&BC\(M
J1<V#93#LZJ0/\L4_F?\28HXb[7Q3XbZ17P\De#A5Q6IG6O5IN+GI@T,=#afDJD/
]M?1dQgHc7E+cJE8UA;48Kb+XY:86DWX7/G\/1MD^DJJ0J[AT4#><7],)2@K[dVN
g2#H9aS&70EVc]:ZTW23(?E;M5R6fN]U8>e.Kd#.(/+DPd5_C_=d5+AbR+:IW.BU
/c1Q]fQTE,.8O^HF?W@ORK9&>T3=#cbb^9ZR./f3+dPRQ2a8aU70VK0FE#EP7+^Y
/1g)cFTa^ZR@-)HEUML_1@5HaD9A@;PZTV]cPLY+J=;aWR6@f>H18[INb/53]gRR
d6DX/RG(7g4]J\6H0RUZ6TJ4V9Vb,2:<Q884,02gVC)/19:X;ELB;202#O=TSW2d
Wf,aX#+e2\3EZV<04JGS:H5gHa+5\U<&C9\0@c/L7T2DUFCL^G(SE1MHdGN^#)@b
3&N7C7JO,D;dPWY[?):X+<E:aNa;X;.a/IZEg[d\.<c@U7KEA&BASf)15D4O\^9=
6CIAgbI_IeTICMdg:UZb=CMLd#bYS,@\.0T^47SJIXE7_H+PRJO+5@^4OV+&UY:A
I\GHG56SS_XC<]^Y#(K>PW0R>-:1NGM98?PB=8#.Wa5d2d1P+:B.:4@d&J12W?bC
Z^4bZA/\M#&+FODF<\T<PQW->3E5((LNU&@?5_VP<AW..Z[K/Qg\e.NADFg\6eEC
fDZV?.(9)c:4#@@;9T^DeSZ80J@1LE(<,E:?d)F=^[PVDP)6ec<<AT9WYM.E^,;^
E_[-_+/RUGUFX,fPBL+J1b8WRQG17/K8:[R<^V^cG7PTg_KRFG_:S?5+[?8@)>X3
Y0D;O=;Y1@5SPS8F#A;T-;:OE(C15.E+:5;&S#B8gBcJ)ZRgPH65BR.,Rd]\bSXP
6YIG3U)V^)667#Aa]8@B91V\17)C<DcB.Z\B\ZF,&M42.LT]@fK#OPE3fAC:R2B+
3_BW95H5SJ5LZZFLAf]JUNUVGQE.I^B2U1#c(8I,^_VIfb5YD/F34G_Ge;IZR^&?
)#[TK;g-D#&R>U3,<\9YNNEe3V>9SSNIF;Z[-Kd[(M@e6&/MWbcWafM.VWf)AbPf
X+[3NI.5#F[?M[(23.JU)Q^D;K8+?:bJ90YGV_H2PD<:1O.dJ2HDI?g.8DN&--TS
7Fd\#U1FPWJW8O#+#&UGNeS/ST_dDZZGCcY9;]c0]L7CGRg:+NUTY@SMVE5,9)]f
.KSUBTOa:=]\&f1V/;He8CSZd1XR&HAb+YGL^&PH03/.+Gae4M/2@TT]2+XNWPH[
<e,(&(9@NE.XUOC[WG>\OO]b[/]<PJ9KAZ(IJ-X@=LBZ>=2XM[R3T:RODOK66-B>
<U-2)W(.0g5aE3((.UT2K(:-8F]g6cXZIAT7dPR0.U/Y[RIbO03B9S.MDT\\c9?e
_+EAL:,MX01)IK,OV4>]4HQ0NCLRB>+L,&Ga^1Ub_2FF_<<E>GQ:3QI^GdTGg\#^
Q->[dJU8BANHf5GWM7@[aeDATVgK+O=8V4EN]g7<fLJ+2AWSHc@4KXON\Pd>2aYX
c.;4C<]3]Za#OHQ5S8[_A1fP:_#QZ;N&67W5F.3eW?;IW7D3TD791E:K;QUDe4fY
-fVgX0aO_GOWQXFaf.[fQeQd+a#6-<;[@ILL3=D;dCQBW:#WJ?8F=EVS(^dP=T?+
YQWCH-I8,6a>N)]GC>g;fA:aPRG<MA-FE6ggAS/1U?,L:CP&ZPGAL(9[fb.@Ed>)
X2S#.\M1bX^4MRUfeg\S.,g58B1fN-Ea?X5ebP.B8B^5]9:A8L[RG@9c^/6b/_aL
LK#T8:(D54VYNd&W.f\LG-d:1^26<gMAFD?gLGJ2V]PeK/VC5IC/L(ULaB]]gGL:
(5=,2/9AIcT43D=/27:MZGa&:7,^DI(RU+VL\FKR)g(@AIb8F1R6f2N3W)5GR-/5
)Y]E/W-D6g366Be?dX/dI,@C3G^@aC_S<AG74g,;,2FV9Md4TO4<D\V-eAZTE_@9
[/?DN&-^J)4b2FKb?Ye.5D>(3QcM^RZ_._?J,O\FZ,;X7+V0fJ3N4\DA,<R#/AK&
2JgMION1]9N?)9P6H?Hae+M&L<Ra2;:6YEIHDG/-M?d5^/Pa@[I@:)>,bbfG4ad_
c7?ARGe&SFNFDFCI=9E?0X0LSH6b&2fGWa7;##[3G)<(/J>91T.?AXB0[T\G/#P\
^^NG5;ZVGB(bEBQfZJ&GG(8+-->;@4fR;T;YQ3Ua3g;[8NBOBgg=#Kc?bgL;BITM
>:2?M7WXR13\Q\<6dT>0/172,4L6b.b<0+DVFIdMNf@\[+B+aD=7OeT_bF/Q;Zg9
\US<-@/+JU\\>;EZ#eE&A&+>@[2UGA.CbD=LB((2#G5/A[P>R=#5217UT40,D<NS
8/+]V)De;[X24.JGOEC.cM^^)/3Pf]<P,TB_[MT([-Fb+U][GO=-DB/6=33,[;(4
J>>DaG([OM^1?E5:6UE9?J31XA1D8-?I&].c[\Oa5c?>-<ZOT-1WU<;1.2>UY/W^
;Y9Q0[#@Ja5>G8<8c@HD]9)BVNBGFf=QUI>>):>K.CR8B:3fOA_&XR:]B=0J]Va6
5ENFBG=]/\+#bV<XRKe0H(A@3;b[MR8^LS_N5_/dMUFaAg)0]IU75?c:e.:Tf@K?
@CM&WL5]D#A4E7>A:IMbTL8eA]aA&O^?=85Z@[::@A7e2B5R(68#6S^)0L],1?J;
,OU90?S7@V]15B8JcQN.d1R8<0.ZXLR.88R+[PDGaYHfY;E__7cKe7:QRJaLXM>)
(IfTZA0;H6>d?0]Uf#)OEN8V&B)(XVNb@W6GI7=<NNfUUM[61MCDWSUD/M+,f1S=
b?.NVCc=Ve?G#GBPT=?df,/,:L<_NACJ5=H[,8]S6(Ke=_KE3B9f-M<f>][F\Z+N
_&(R8DecSMGR8@.K&3eF_0Fe:\,[Vf::C<<\Y4K7E(YULXK[)1BG<MH;E]JTS>5^
S89?9[a=P,UF+(^95_J18fXBR8#S&5=K(KgXJbF@_?Nd<\&15>-UaYB>b])>4J2I
IU95LR)E0bf1\XO\RQ6Fc5e03a[=X-HUT@OWaEc7R\WeKUSQga#/\=.6DKY[6/^G
D7g-6b0-R3P,PA<b_(9ZSd+E#fc_+4:>/FIeJN=0N1ELgX4=d-K]b9-^4H0U84&V
DG&b[HacJN?AB__9gN_cfW0(N52K@&<XP6#I@IX3SZe<Fc@:K/>38K=@\bQJ\KZQ
VWAe[effB7B&4E=c\baG:c0DYIZ:V?]1=Z1cF&;WKAg&dOOc[O>_4Q4EbUD@+A@@
#J94RY7/:Pd^g/>@AY>DPbM8HT8[7H7b/SKNeO1+\L+<b1JD#0d7X>GE3f5>KEIN
RGJ),YV41FQN_bEF3LV2YU,3(+].G:eR>,DV1DN^EV[:Wd=:FHC2d:/>8D0EDWG7
6((B(NZe2e_11M?gK0gDULIDTd@E8W<6J#YL=),e:&?Cg4P,ZTX5,RUBS;T2(?Ta
N[H^Q8-WX(/GM:f3PAUGc[58<eM4f[=I+A]+DgJYfCQN14Ef29[Nb7bJ]>dF=FS#
0eH)[I^+.J[;Z,,BPH_AO7]-MVX),L<[f^a&+<a<51R01_T[^W0JVFVJ,C;YBQRJ
7^2-,[)X7dTE;^fB@e:56J@Ug?<:=3NF&)2-2XP.G&>1@Z)=NC\1Ea14-g.79\#F
^YYKCf.=OF8QTBP7FJ]0:<e(\A,g?5AJ7.EXOC\f_G/e;]K?L_9OXTXcO#4R:2Lb
/+EW1S-E.GgO:-fTd;]RaQ2MV>:@4SNHQ35g1H5G35L.M<77I<7.D,B7(=]F&c4\
70/+cUFbLN^:>+D(6ZG:U<Q]8;K?O2T(28f(7@-0b(=FPKSd7U1].Ofg_YRf&>BM
DDD\<5;ICcY_.&1XZS\:UED(6II.X90E3bS8]#PI>,CCK39YF5JaFZ7[Z#BPOeSJ
-L?OU]MQM-;UFHE>4-f6K.[bEVP[23[=+\QG#<88.(R7g2F6S)H(6CG_8R,^?.,?
G9^4<25V;>H+9?bPNQ0WJT;6ZGQWJ9U5+Uf3]W)_.@L6Me.XF6:PUXDGUPR#1LIK
X-8&86d/@Cb<>eIRFO/UZR_F;TZ\RR18KPU,7C@TTA59f)B<^cE]7PeM7KE40C\O
/@]Z,#M[[g;].\N5d+PX(N??L,S_Vg:LcES5BFUIcZJES(YQ&SRB(ObJVV?\/-<3
ZVU7Ye35SMF7AUV\5SSXY,e4R&W7(Y^RZefZ&ICVSfT]X4[CgZ21&(cA,KO#b>;f
>G),4ZL5FW,VYQ@.MaK8AH63BF?-cgd3-&0:O(XR9>?Y-a6I2G0.9(&^3gb(YBY,
SI@5A)Ba3JWJ,]\1_2AS=I+)Gf#IN=C;7S:#RG@=5L:6ZMF,A,.=X)V<K@)6,B9S
TJKMH_gK/OFZJH.ZbJ;1,1SVfF/e56F:>IX7fJ0e1++<26A&;;43QcP]RC19@GZU
E=fCK.2(PE2?,M?RWRQA1]0a3N:R\FA&Uc.R_N-U=C-ZX>A^<1F5UV.33G2&eEGE
+:f)H1]#>U,(d.,6fSLS:eJ8eB2gA83fV8C=>K.#ZK<8&O(&gCP3PbBgV/,,Nfe@
[.[^;<U4[Q.LDe-#<&,QX2?#/gQC^:+T/T74XIcdF3QG&_a#DSBYG&?8?\9^1\dL
E5cO:(TK)5MDXER3^4FEV(8J61gf2\MI[P=(&/\M^I(@N&c_1_fe#MaBA/<B5VYC
0X@YZ4U]20/AN[[S,;DY+Cg@XeG:2-a]4V?aR#54F#WdVXS@ZF/ad/eN>:L.)Jb7
N&.eB?)a]<M01<2.PF<&c<HK1HF.CD@>4/)=;MM33MO)GGdc:B@6QP&KIg0HT+0:
)3[,RI[f79:2KR[8Q+OLC>)[E==@@,[^\eUCE^.OU\&I\DLDM=IKSSNb9a>8WO7,
SOYZbM_cRT90eKFe<J4&OG_,,#Pc:gR?=#]6G^=]DXKd/MNaZ=KFRV+9TEPW7P2M
GXG2g6Q^4J#OP6Hd(aA3-TRBU+CMb8cS,>JQ/R2ae8Af/^@Kb3[;[54dKb+NCAWc
bV=deN8TGTJZc1-PKaYeO_52G+CQ-bf1#,OO4D+^AU0:BR(16LZ]c&Xe]_:f)^2-
A5=HY_@1LK0F1?[W^L;]a0#@3:L0=DW0E6K.eWDV5M<5F7P^5:aUQe4@+H2O+M:_
YYY@G>Qgf-<H-I1fO[d5aMaa\G=,/2.g=MBdGfC23cATZ&7/63ZCF@L@;HAg2:T;
Z1O_M,T#P?IAgB92[SY6=bOf33RBRAC23H6:-OB-#(#5UI^Y\9P#/]TKJ=/gWESG
4H6S#@^8<aHg34_IUVV=8>Vdb:L#(?fOB-)IMOTg.&M_b^+KB^GDO4VOEVLB5eU=
37^UP:THGC3O_)TQF[57C/6SVUQ+0FCU/EKVcP_L\L(dFX_;f-XbcM/:.8V\.LY>
P?#fCVf8\D^0S.VS?_ADEF[DQQ.1.&1E07F\Z;?f7(0Z[:POdX#ZC_I^(<H:JN>B
^1BQ#<XK;()CaGc(NRXN6FNRUAU[@aL)J10_VFER5X+FMHA,(A[2Gb^3a?#d/79X
8(L23?&gM0KA:OYFVW+_7X/,R=HE>2a/V9g/f6W:A@B_4<O\9_D.[BUb1>0c32S_
?]P9.4G+3R>A>7=B3Fg,GJ478/)/3?^f>/PUV,(7SB+50K?<5K]eRfGHFFeYB1?;
]+@]44M9+E?.@Q?d_)5H3:B?B0??:_f=;1/-JFKU^^6PaeZ--XZG1QeN]2@Ta7;2
;3\S7J.;PVK8H[L(a(NcdW+MB\;P?ETZ]6+:A-=-[G71e\&d[].1G@,]\Q.&d[a0
Ya]#?PdTV-M62DGL//].CCQNY2gC;?;f>?7:(&+-\2437XfdBH\,bg]F&Zf>&SXX
;P.<g,>NF166+$
`endprotected

`endif

//vcs_lic_vip_protect
  `protected
G?-+EA)4>UJa?.a=(W,7\4ZR^_RNCJ]fHI_T;)Y0,BaX.8ESJ.6=)(>55U+91d8&
@H+=GEX=]AGQ^[@g(.1,MSL2<W^7Q)f1->W6>K;D65\DKG0LWP=fCARA3G?39S8a
0].40L_b0L7FffCE/X5RV]#NGGfFKT1e;?ZA.P@\B5S@?2FTCCg(G_e/:DOBDZ-g
Lc5\X6[-R\6X6Z.U3_UR^(MQ-:LUL5D#Z0E[^ZM]+ZI3L&7a570NM_[)1+)R^&Q;
;2SB-EDL-)84SGHBB#N#E;b&N[[1(KTS;1^VUfW>]M)YV)B:=?GEdKUVC76BT@(G
4W)483]>():(&JUfAU:<O\T58\Df&ecCQ3@5J(@3<4YGFdX#gdKUM+#E0+7XP1O6
g?+8FFC^W.CZa?0N3)]BZQ;?\:DOV5>BSeYfXO6bF:dNTTXC>,(9\<4b=f>a@2aJ
3Z;PFP30PUa;JP6VW<&F1N=DAe]Xg81V<N+GGFWXVS<I&NZCH.>VD(W0CYa/FX.K
.SLE<>NAA]:+I_YY>@D,@MJ[?<9d+N3I4cY:O(YAB^Y(A;a,f:0,W6E/Q-,0]VdG
ZTSO/ATC^5?H)S1YS#^]g6TJ4,P[54BTK_1^++T/4ZV]+HO?eXY:B\dQ&TadQ#9&
MB\8OQ\/WB=+73(M\Fb_L7;I;e@LE9HJ1<<P,6&db,b4.Cd1]gCP7@(>Q))/NRG:
PWD1WQ6?K0(95QY(U5ONBEa,^.DZP[?&MgfYL1H+K)OD7JEI0CZ:Ybg&9Q+aNQf3
R3Z,.f#O3-=(W6MPLX=9E1]gZg>YJ.8VaSKJE4\ga-68daR:UEQDX.P>2eP5=LQ#
1YM>e0D1RZ>?0a(McUFC36d59>4BE<31@ZYX_gK?>\2WBSZ+OEHZgdJ(RJ[:,a73
(SMg?+M0-SI9@f?,45,<+a.^;7f#,6a6O-ZOKHNeb?[=&4.]G,agd]#?\Ob.::&8
M4[ef^AGg6dGcC,V9K-dO0>f0O-T5AX\ZDOW5USZ3gI)SV_JPbN)M+ELE)8-#=HX
FNL:3>9)53BbQN8#Y.&c3aJb=eVI>4gNX23F3Pd0EL0fDAT9MWUA3O#e<BV&RAaM
TQ^97IZ-H;>b.I>0>=Va]C3?cO1JJF>I=N:Y/,:b@5DHg+#^XC[ZOHP:BBNNG9H0
^SMgPW0Z)<O2@_UcRR01\Wf?g9#3:]R2)g)FURC(=_7XcA;3GBcPKa.)6^-+973>
TVA;2cgC?f+]UHS,HUQK2/R6-8<eTT_D=V..bJ_+(1++0,(W#LW9J9H3\J,TXC[/
F)fQ[0;W625<XJg68)]2NKY_<<X-D<TJHIf<UXTEUKW)ZF6bX#(5WbN2J^WE=S)9
ae6;U5;MI#7FX)>O3BD[6ZfX;)@@DJVAG6BLC.XO?;J6g4&@b&U0A7Sd(Z&Q.Y\^
2V[#Q]U@e(e?Zd:[&VEABY/P4@,cSHe]F\,0H6V[DFg(:8D:.UTF_>=-:E;;ML,g
FGFQdQ95eL-FQ)/SKT::4=GDVFU<B\R\gQg\M6J1PJ&],HQ7SgESN-Q1()O_fO2X
^2MffDUI2W/245g65LA5Mf;BV3-4/XfS.@=)4D<EVb8W+-,LCADXCFBfOS+dEIBN
(,1X?:Q=B1C3,3G9J=TeT0G5B9W=KU#T_5c9;N,)(&b3ZKLe50L:Q-Ba2+X327SG
WD]N#Y9fE[gdMT/+NPZOI<<K/Eb:>c<f<7fd1T0K=??<(KN&R^^=4TJZ-aX8U0GI
+g;<TZRH>Ne+ZNX2MKE.F7YZ-@]LY_8a&W/<&T37L4Q]-YH9WT6YUL[/2J3\5=cO
3)3He(-/TD?eUeb6IMP&a=-(0MfC1Rbfb=VNJEd-R1(CXYW_8UYCecP:fU:QST;=
,N/YS,CS?cPDZ>B3=eD4H6aZTS-EBgEAE\B^OP@372H0-@<F4PM]SfE1Y@SRS<J@
Z(4&+CLNb<R_,7XOB))GRNG#Q^73][W+c]R6[AbI-(fe;:^NG58Y-f3FUO)bK^g#
?Y_TO5UDbY7HKfYJFEYg#2@+/eL7e&PKgTFK8^E-;d&/O?fGJ&_X/J&_F1N#O;cI
78b=)J&0Y[-GW<;5E>T4J^R1FKG^>8Q-&8Y3YWA?()7fIPUI>-(QZT^W;LP2c:HU
WZOSP+TGD;ED]NW<M67cQD[5:fW.:cgcK\TKKKB>Z2+#:7(I\>C^/f>a9^_Uc?^?
bS=\R?>R#DMV]A]<6:AZL>=cNBT)GMF6ITd:[g/0]ERN5_;YR@TQd1R^/7A0+J6]
JO@.760_We^dOg_E?F)@>^(?1]R6a;:K9AH&QQ+&]RSb)4B43a+_5>O7gGX(;H]9
J#J:-TUF]cR(EEDdBf@2/MGP>S)NR>+Cdc(&I^ICL6E&9W=@7;4B8gf^FSH(?/Q0
BT++XS+GASD,>bTa]]1LO=E25>dKU]PI_6J?^1B4^MdfX\+.+bC^3\9-dN>FgT@;
QU1\3Z0d9IL((Yg,SC3,9N,bK-dV;bE&dOfEQHP+PMFKM)[=Db=\cf>@:FG<2eg4
LOB?(:0,J&4);G:9C#O1Ad)M\@\g<09N_X^A#Wf[,+J;JC.F=B;3VJ>>ZU[7U7BG
>Cb52E7]@KMa7:H=R<Q4T0H@Y><cHaGg3(Xg#a2a:[B\(/9CY>.]OU<Za(D?_YH7
FD5H-TgLZB+9\4F5]RdV(AV(+8d@a;H,c4;8aO]K6I0S.?SIbDEQcPUfSMKX?].Z
b&,JP=Y8-OX:)L3ZO(5#5C&DZ,W_Yg=f)B^>^(]N<D#0^;X\FU/gB>@\=KE&3G[/
=bJF?/aYB5U\/J)\)gH8,g=H:Fe]7Ac,-E>b\Xe\S)5;<)6b)MgVD<3&+IM:d@VV
YecRa3)B<g+&[00^(WC=K9P7WT=1MRWS/?YNZ5A1aNMRM]]Cg(\,I[8^]31dEEOP
b3N(0eDNQ<7BO:gEW;@8<TA]Z:.>M=3N]HHgUP3#KgZId<H^ZW=GD,F?)_+RL@##
-WVK2Y6)d\Q\:@X\@#,4Ya_QGf[82NGIGK21S/^10OPGb+<6:0A&bK2W;&-a7Q?-
:a[#0S_cdA203&H[YT2[-=AWZ/Q?_=VeOJ+5Yf3^gLI)1]P&LRN))&=Y,CSTHURF
#;>S(-(KGGf,IHE)8B:dCC6Vc<Cg:B;OMRWg#cD>WT.+Vg_ZREaC4L@[YH.b1WYA
2^@[eM_g9P5(L1YEM_503OEWff?X:QV:X9CDEZ.27Q^YY;X.S<[,GT4Ub0D+XZbd
N4RLSYgX1#KOL2)ST92Nbd=-B_SR6YcWTLRUENT_U+P[33W-_d=+N:A;^[GC8<,6
-LW,a_a12Jg\\ADCL>GUfF8NWcgF15)LX9]@+UXSGJ\H?3TR/e@:P47D=OAG;X;I
TF(BbaQ),:Ga6_-\dRLT=EWH=\2ZY;&QRKO]:D4a9KZ39GcN</Y-dT@)+8Z)Za_?
J?GI6AI?#Ad7S#P[Ydf2\NfPNfATD:,4:cf5,(CUUMD)C7G34g;c&aTYJI+1J^EM
)O35KF#OBg_V_T:.L:Y^gdNeR:_4#Y5,6_93N/E)X#4OX;fBKe@<H#0I(D[0gPa+
]VgP2dg_=dI4(]404LP8IA7ScFO?[(aKI\_C\0bBNLXKG(B0(7Fg[-,S1Q#dE2f.
(]S02eF<4-L2V?0<bUV#L^V/C+MB?W;@XW#EgLJ#X7FKaI>9aR_JAP[5\C#<>(AV
&e\e?H=E&DFO11?3c-SH9.\#Z9CDZ6M,=6<#BCI,NN_T0FXFA8UVUGaQFe5]X/KR
eN;\>I5[W<-CA#10dJ:4F2bP@.RS,gUWM3]DcEUT8?3/</SGKNP=2Ha20M6<&+J8
Q<c;QY,.aYWD^B&0)P:2]Pd,3f8YMQH,=XWA^_EQ^+P(gB>+4<WXaYI?,\<eWGb/
\L[^2#G@IMeY>PT4Y2_VI_TWU7T>7)D.4,1A,7S:,#;cU-TgOJ4.dg1T<(]@9f5?
CE,-Qe]bZ??ebWX=5;Tc;e:98]0505EDGLW[d#c0>JB78Z\YRfa-.97,/.AA:&Ve
4Q^C1]c/JAX-g2a9HD^MI+cf:;DEU,KOLRCLP?T:==C+G=a=[[W?fA6:\?M&Q(]Z
MD2#8K(H;V\_P1C&_==HPf[d6E43e9(ObG_1aV<]gK1EL+/cMU9#K^ROK(77A<SW
[(bOYQGI39.b0:8;:#+GE:dDR<]@P_Waf6)R>0ccNRE\I__eX?^>2E.H<Z5f=A4.
Wb#0Z6.\CG@JPC)<Y5[93O8P,\0.1LdM#<;fJ<T6Pe@Nd20JO#+:JAVJ8SR/gg@4
a#AN,YF=0<DP?GHD-Q<>(E:_&E4=8[gUA7S#Ub0KI440C,PS0[B8MEO8^4>PIDW;
)g/U_g53BS2?YNLQY1G@c\+>=0[U)CEEd1b[QWVYQY3WMg@MdSD+8AF4=3bUFNFA
<QIWU;A,fPR?X_F4QND3=[:GHR>;c63&8,CWcPG9GG2FgIG5[.,9_WJ/QZ>BO9:/
&OK;?+dC)GG2VJGX6:E:LN-]/L(cVNVf:;O(@2LXOE7EIYMA1APD3JQE?W?ID8<b
/))K;7/e;RQJFY^<M?[C0I(L_XR8PN.-0U^H0,W>e]1LK@+BSV>.>Ha0^F_0V:.?
]L6V;+;(aeEV0BG^91e-841U@;>_>JM3W@E_T:C0feZgTLB?=D[DLFV0G,_FA#CN
)P4c0OL_;C4>7X^^K0AF8<9LJgL#7&#,bNH<KfU;BeRX<-MQL\/-<e5f-6E7FZ&<
G>Bd3]HCI/Z0R-)N>)1e:gA+(LK.,g?d75/,K/HA)P@#K<cVRZ<(B,+W,QgYJeBG
:f-Z;.+&AULI6Q-E#_bWFHBYc&fL8GSWPYB<W4HI-C-3c2Z_SbP0E3IUXT\F\M]>
P2#1I0g:K:+9U#Q6FELWQf91b?K85:KDX?H5??&DTJ_J?8J0?//#[F#_>:L@J)V[
-SgQBV)cJ<_=S0^I&95.PJaB6E4dQeeaa?[)JAd&DaLgga6d5(2D#B6edF]D_-?M
\9dd.LQYf,>ed+C?CF@TSP3PO]&GVSO94B9^N7Q.ObT]_a5N==L)Za[aTYa<(cQ0
M+>#GU)fDa>VWW5/]NDb2.1;L/+\P/FDG..K?>.&cH9Y1F[VY4D2D3H8XLJ0?Y)-
\<SW(KJ]EJ5C:e@Q04;VTcW,,4\F>:VUR2;[GV4JNT#[gC_=H09b2N)64bS?#^@A
Y[7&gad.)G(D8gA0F;O/A-g>KPU,]R1S1QL78/=17IHcXXgVA^.fgG&KLaM<e4LR
/G?1JH\8=QT[60/VSc=3OXD+50bZY5gT;SC_NYXN9d#J^0^L\-d\Yg&J,VTbC[(L
ccWf+1+7R)35cFH=589T\eWaNHH#IT(VbA[6MW^M]\EVMIX?X-PK[]KC]#&Oa;>M
TBbM&(6V4HR.Z58DOJAD:V6(E@S2BCN7>4=+30eP[.M6:.Q@CgMG0JE9T7<:<VU@
DKYBW,fabBK_OQ@KQS@#O:UO_BaZJO3\U>,;TV4;1<C>9Q^5ZT:.a;e0CgJ/?8MJ
H8++:2e.L?SHXML7+YWSf+f+a.2WVMKXa+RLDRCAKbCe&g7f_#EPACKXa8TXWNR<
^)1-;Jc#eR1<-(]6aG+0O7fQD4J0b<VJ[.a^[_MQD?>bZU6@.P5A&S]#K>Q#X2Qg
.ERPSZ@#&cgUEFEfc?7g^J[]+^DVb>B^HT-;AR+)MGFFDc-9K,>]L#OSeR#QT8=]
KKbG>,[D#[:B0=E,Y2A43DfXcc.YCSBL-H>Q<8);VXJW@\L(d=]bLAV#b4OQaOGe
If<X]H0/^d)G78MX6@aYM7>8@(3g?+gbB_#:d&V<>LGT1DQ]aI[23FdP>N7_W7^0
eZ8MP24Z\3,REVd>ee4F53H.NRR<#2d[&;Vc1F]J.<YU\PGb6>\+</\8D8GMN&Le
K1C05&(4&ASNa(/#+6^Z5Y(.+,Tf4ZYA\Z?2\>J(_=4TaIMOVXTNCLK7A/+e^c7S
7:??V,;[G8U1aY<RVb1bcQ]d,3cJfa&-Cg&=g@fEDQGf76?S?B+c-V;\]MA/K4e^
4RQ]/S5IAHg:&@==b?1bNQR<BLAe,/d[+^2P)ESTOgL?d@+C(#OC?GT/W^V_c3,a
.f0eBOS)B60\:]U(1>/WU0K]WMM.V+_?b?(:_\.<F-K1<X^I])HZgHIef.[b627#
WK##&1e)@NLBV3TY=F1]0@ZE_I^7/<0@Y+?IJd.f4V::+JO-)E/?I.35U2&66Z6C
G;G0]a7OB-?]DC,/IBe8PF+(DNXBE(+GASGT5=^:B4gI]4YXI(ZPJU^#(/>=]1^U
e53U(^&YH:6TJ.N5[]XAXY8+IGK2N+)-TGD+GQ:=-U9PB=Z6#.)3V15D)7I;2:IG
CL<MeUTIcI7/4O;HfP4?4S5_;O?If+S3,T01_Td8Ye)E?I=O]UFZbfIb2#2E[8QN
<\bY>X5_Z)TYH[If0Ag^-Z7d);1<];E7_SV?Uee:)NYOd_HPO@&)X\f^(,6(<bR_
#ON<G#60Y:FE4QfN13NOeM<3\M_adB1T^)<+S/V_Y_S.fBDY\3+\YBUZ-aV>HeE@
@a&2>3,FTECP&VKee;?U+4;ebf]PHBe=Fc;.McB+.V0ZLee/dODfMNHSCE=KL]\Z
?2YZT-UEbU+_aS\V-;<eH+g5>[5D.7@0<WKf6L496FU\11YSS>=_\3=SHF#>248+
QONZ8N:[3a+b_Q6C3?+]VS5M1I><7c,ONIT58-P/RK/8>EeM\8A49,a9#fNZKd;.
;GY>_DdN<0Q\?>^L\b4E)Z7;aP/4F.)MR9/RT<\H7;UITB_8,+e0d:8f?P;Wc:N(
Lb3;VN2JTF+GXf59XPGUce)g[M2:,A(C(E)+EPLUHBV4\;.ZGKV:SA6bVc_;8/@0
FY[f<<^b09-&HWK6+21WBCQR?HJN1/ABe4K-@)5e(H?:/OR./TW2)8:<XHG1:Q(W
D@P<Jg>0\3^@6RZD=U\POcI-:=VPAB0>,JdT8/S7W20N0C2+:dU5NH/W_PaZSPQA
&+66P.Aa,<J_XaI=J7VVV07V-.EQc=?#Pa60??\2Y<2;b>1(A2EOc6;T]?7\06:d
=K258M(9I4>>I[Gg/<)LB[baWa[KW7?RYFXA73PH.])&R-KKL;cH^cP<B15_V26g
K:R>#)FII7O@IU35C5df\VKcA_;B>ES^Zg-4WRB7]&/.DI-fI]Ja#-gJbbWSOVS,
YL=eQL1<be2M)U2\(XB0OeGM5X32Q1)?W@E/aC59QT[[A6AJ1G/5TV]b[.GAgJ=g
MDK<27)g)8P]-gI\PKfI>G<T4<R2]-1/J:OJ45M22caQN1JMSGNY1F(KJ39aS8Y,
P^?NKgC27M29)eP^F)7(A0>f8/,IZ&XdcPFZ@HSebHOXHE>@PQ3FSVXS?94?W0#a
M5:.R6\48,S(TC6=A5RT;V2V1BQ^DLMYVdG?/C6a-5R:aT=^c\S3_-F@D-]N1QC)
GY?eNZO+B>VDF0]8geN(JceC868/T2[N2,+_2c&US(#\TgP,;).NGGZ\6:g4NFR1
9aT&E^<),\VPEG,I/ReG(OWXEO,DG.ZB,H-7JO_agXfJFGE#<C<a2_eX>>3JAE+^
;K2FE_3_\LU_7UIEc77+W[^P?(\;R+]R#1(([Sg5I&&/VZYJQff,P/89\KY\B.AT
#HALRdg.A5Yf8?C8W,MY>H1<XEYSD<a[NC&U-+-8]6WeXQUUPKMg15-#+=YGgEc)
MQOf6/EG_:be(&(-b89;ZHe@LND&.f:9YDLF9^S97AANReNIePY]YGYHJ1GM86I(
Y=abYS0@c_GM.K:8EbUV.@+bVa8/#YH[[_#1W7e;Rd>(Qd-E5.@@32J7Te^)4KE)
+DR)@YcO[R0a9Fe9D:TR^@G;K,@GB1.I[WKJL&;/G@UWI(?0]=RFY^Y\fY]E16d4
5+>e^(_b<U;.FgTecUf3\X\282b&_<;7??b&bP(\;PEJfLbF[4dL77H<A7HLZ&eI
b,]4_33>)3[_K<61O<VX[4R1G&+deYH:@FUSS5R1^\AIBMNRFM6IN8PK8AFMB)P.
9RbOIS-JT(JbOf9QUMT+KL1B1XYMYfC,>g-NMFIT-[F+7=G<M:F5BWLgbY?H+.U5
(M?Qd\:/6RVf-\\5,VX^ceNbBJKaZAV^DQ0b&(1UE;?E-/H@H]4P6Q@<]NWO?[Ie
T9C4GO+]3/W>X[5.^YfTbBEeK_+gM[;e8_4<Z7Qb@,^SEU--)45X\6.2;Y,L)X]4
&S17AEBQ:#<PT76e9[BN.,^1G)9-e2V22)7e4FJ\S@\ZD7I9cce0(L2DE9&Me-21
PbC5D)0c@W&1<^bCFS[(/-Ie<SV.A4/00dKRL^dD@@O4P\KZR8P[S;ZJRMF@T+gM
IJ;/.S:aBZ3,KY&T;VWeJR3aA:LN,<ZE/T7;7YA_O-^3SA?.GVPJba(&9bE=I.g]
FCEY3SB\C]\/UD+Z/W4U>(eW.FeH25aW=NFMMC[F01\2MfZZ<&gc3HN@5c/.gVE)
V[4,8DE\>RK7<:ILK.C@P,L:2IT?0.AZ^JM[0W(A(Z5IJg0_S5HI;VS^9-B>?(AO
d]#VBIOa2)7OJ14eg)DQ,;932OD<O^R\Y8Ia,H#4>;T&+Y4.Pe@T3Cd<MT6,bCL]
IR+4)IT81K(9T1_6AJgcR=>A<\CJa?#Tde_I&\I-7#H#Mg07I2:#-(XSfJM.X(FM
\G-UDI;N4>ZMB>1PJ.2&4D>SZ9&EC9+.Y4cgEfS]92+Te+?4HHF&_R+L+@/F7WGb
JE1N:S7&RQ9@J75OCbYFJ[3b(B<Ng#(?<87bGMD(F#VQV.6VeR8)8I48N--O-ZGV
+YQP-W9-=YSgcZ7:U4S=1fA8=X^a7HIR;S&50[5Y>,>9,RI^X;RQCXUZ;Ub(B;9[
aeK3#L.HC58&\D=^LWb.5^Y6a/V]fSBQ#8F7DU]ENEBd+-0=5f&6E&UKeQeTK;&]
fB-Y+=HDEeK1-3NNRg&=G)9]gX/RX0B3E6?9Xg#G_&&X:++f.bP19P\cU/YSJ:-T
=A8E=)31H93G&)MEM.DONB(d2MRCP43&C-[U23T+9.faQb&P._)-RU^P+95^/?-9
5=;S6D2P[2W^+-XNI8)[gL7)g@]M,NPW8gDN]87T2]0Z4FKe7D\Nc0[60>S0QZWG
aL3URB.R_LD/-\<CYZZUeISD=Z+SL^)Q5Y.Wa_JQa/+WCLPLN>[+U,P#K,#bT5=1
K4N#)SbgT^T=PJ(2K+CQS6YeI@ALWH)IQ0XRNC2KNGQV4&^B:>#XZ6g/6\c:25:K
RMd.CW+8OW4=M[RL1CEZd89\J&EFe^G68/.B&=FF7XLe[KHGbRab23QVcFDGW4K(
Q\6_O]13H-3QJNfY.VI+R+1&]B+F?E^D7KE^K8c#]7,O3Xc[B:&A/SfG6I(<dCC)
HR&K\Jd-<4<+_)9L)WLa?V#cOe.JQGFXBEYFR>fNF6.Ab_bPWTK:SHfGK7S5cQ=c
59IY5?J(FfRg3+AN,ZbJ])U5\cK.[;V(M1RL)\@g1@S.S5Gc-3CN6\Ua\_d,1+A-
GgH6=D_80^KO(^?,gY@fTECaB.1?;:H?Af76G+T+^Z@<f)2.gNR,cWg]EfaI^C5A
0NSPW_K<IIT)F,8?-&Z@PD8SU+-U8KS,gX\N)Y_197N0D0\.V5dR/0a@>#=?V,KX
e+GHT9DPf32)R?\TKLJW^HBe5?gF23L,X3R2V6/cC\fabcT&dR&65B_.-;P+fGN<
d<MRffb:gcK0b2.?/1.bQJ,g77\-J:fHIgG\,FTL/2,ZY6+GSH0EY#L3UCfVf3P3
QAF;Y:2H3aRH\YY#VQO<\0&6<#SBOcXKc1=6NF8/X.QgJ+S/KT:0A9_@8A(:+)e^
C>,[YgAC]#7GSBA8=QHEK2EKfG.R=a?-.+F_PN4B^T:Y,Ef]R(A^WYGLTZFcTFM<
6,L<WTTc,CP(;XH>;.5f9P2QMYf/dV;P8]+5)=KL^6HCHC?d2F#7;.CMZ@3;g]PR
E2YUSGfKEZ=;JKbTSRPbeQC&PY+(Dg^Ud+3;cAaVRQ(G-49<-7)W42?U.6B_K?],
(IeeA@H18d=FM__O+&OOKDfW\LU_\E7A2Sb+?CJ@TUK&L85[YJ/]gb9VJ-Z.;.VF
<BM[4]JQ)#,A9TBWbaCH?Wc2L75&WAUHebS[G7_EJD=R@-]1ZN365+BO-C&N\K^A
<EV+IObZd)D39\#cA:c@fZF-c@ECGY@N+=9#aL9M<E#LKK0-LB(8BED0>=QWcdLS
=b__d\N@\+Pg=NMZYd&f\<Yb[+/Y^SKG^,90D3FKTc[2+VP(C,EQAPeaL77N9X6E
g99G/OEBeVBZRXgFTIH3P4Sg#TP59<\:#c[1e4#HH.VPBHE@0TX;70KS8.b.^.TW
++K><fW@FA8A,7(;OC0?\KCZ6HdYW=(f@LT0eB;7<ILO)B;(Z4X5JaS_T]^0.[_0
+e+4(,.C,A0TAW1_<S&&07N?6-)a(aKNUA;4\R+V.&4LX)Db,Q+69LL3+8905)/-
c)P;2)BfJb3#_,W.9&<3(/X/A)DOYA)H7^U(P^I>DY^571bg5G(dEZ@<dZE#a;+3
e/Wa+eM,.cZB@WV;#gM]-^5<B<4LGNZ>640aO]Da#Hb\LR4131;H0D78:>-LR54U
_E[#K@b8-9R?IN\Rc8CIg<;GM#151Ja[]Q3[WH_\DVK&ABeO=&OZK]I.U4-)9eFJ
3OC_d]<@IO&16gMKZR9AICX4Q/C+WV.V6R7Q&O?[_IT9bS\fPFXALG.BQ0R#C,&=
d)(+;:V-PT:GbP?HCM)Eg#961d(:=3T]TT;\:EEb4MgfaL<>/:Q/UD(EY+[LRY=\
BT5HYEBY;+__e/[f:,4a6#XT@TG],<-;[;KT1:)[^;E81@g#II4PQUC6_4PG&P##
O:EPAC3bXL&;=+ZOc=QH(4F1LbJ=9TZ@aP5aNd.DR^=9Lf<?_X7.WTSHPb><XV0\
=dP?(+)G:NL)L-JTH#070dHNbV]>R=/AI/Ue=SM>T6FUH\,[YA]PW>_)ff;S+G\5
ZYdKJ:1X]U@8BIFP)6[X^6Se>Nc4D89/O?7G2V3:4V1@HQY2DRK;<>LS\IBGPMe;
KXd^B\d[C02A_M^&Q(-4K^bP0MM@X0T]J,6DM4[AcIWSNfcPOI@C_(eD@KVb@7B7
9<_0MT[4J2-P?J=0[,B]RGK3(dKL0BV2_Jb4b@7Oa\ad/>FT#H6eLNW6G&6U9_eC
ae&XT16b9S5]<AOI0R\Lc8QL<+8Q?0YY4,20ea2TY+WgI38f.#IUL1d5&fH2[QM=
4Xg^5D1=(A7XP3AO<Z3WaH3N>Q&,I-(9+(YTG6RU,,[1dcG/:P(5(B<aB7:Leb0Z
Z)F;OYD&@:H7ZKd3dSRQccXQeHX2<d@[)GX\F0ge#A#=+.dR#IBN-aeDQ<df.41<
.H3b=@aJ2H-F4Ib0\E0NfXXWGE/UK\a:=D+U/W&66^8=ICTGTFBC_P9<BR:Pf3)^
;+\K?c6^50)@+a<C\KJ1/H3>QIK.EZE4=g3OJ^UPA(4ES1M4Te\3?dZNc\XJOW:X
Be@E^8+O/5\J^M3&GKL:E?.JC#=#:T@]a&([-DH7JC)C7e1L6@T]9MO0Z\<^M?C/
]NLNS8O4>1I=5B-XRR>=&B?1+>_(b5B6-6gD0eH,4F([U#(F>I+a]DBJZ3b&+7Og
D-b?F,V.6J5CBA&EDgW(6B)07/6M2&]fL5_7C(#Ie7X>,IW;[JZ-fT3>\EHa)Ybd
Kg<LUS#YF74E3,;.(QH?:[?&=>60FfHSN6[UXT+H^b;&S.BR=I?<V;a@T@EEFcN_
:CF=>-R5,BUZ9\W]b1LZK,S(#:B0^T_]=Da=.E-5gJ\3T3f]5>a,aW4^cX>gDFG>
RFR\TBK)>/VK0R2VR.T3d>ecJVH^XP/(Ke2\dU)>PL#W4A>-Y9?(K-P&(9)g&\S7
NLWdIZ:\618Q;SQ:_,J#E_.a8-S6X>AX_(\\AaL/c,82QW/fK22[eZ:OT/P&CK]B
=AUcgBJe9fd&+:e#YT4(b#7f8#M.5-B_)F4+F.,dW)JP)<38Q\dee1:HD,IOaG.R
.7N<8FKW?RZ\Ag_#_(&1fKF2gL-#^VUEX\/5Le>(f.V(@G\KY2:SFB5L3YJ?.QR6
ZBH;C[S#T8C[M,-MZa<caagEZXSQ6\M=?5g1,S5J]ZMdF<:XY.dFD5OWCUFDH.&A
]8Yd=Bf?Ma8V7QLGSKPUEIKc)^fY?##e[9b#\cgGZ1R5D_gU?U\-M+31:;3eTW43
TB:<eg=;XUTRWL&1401Gg4Y#Z?,?08NN(.GJY4-C1UZBIgaaa_UVZKQ?I(7SLfb_
-35?8S2[@NOJB9bJb7:A6R\:?0-/(?;(aSW+GA-OIQBWL622>DZXUM/&HNEg>01U
H[)d;JBA[OX:eVNZ>HfI^?OJ/Z)E]G#026W#GMO[@YCL?@QeSZ(1L0?X,BO0e<4Q
3DCfJGX/]0DgQY24^90YU5.baG#R<2Z#GbM-DeH?(Y^(U(C<_P.:3S4>AdaA1g^0
FI))ZC+207N>R2b&\4OAEDCISZTN#HE5bT43;==,NC4g1JQNF7_CFAfI^]aQC,Ya
,3L87cEb4<@&;F<2.JK99VfP]E,+gSC0OMfYXd4:S_??-74&^9e2c<0a;TUFGQJT
LUIP6TG:2P=XZ4&YEXLZMOPA,Y27R+9UgX?KDR,HL3fFaYgD]PJE9MB]?fdN,RaZ
E+&(S@=#JU;dDT\\X\_;K@B@\:@_T_2CQb7gR>ZU->c-@&UFHHG;VeaM2K+\-99U
a8SSM/8FS1^A3La?Z8)E]?T@W6;S.6BMPF@KNgFTU0?>-U[Y,>=O,5L0>>1>0.:(
2b6SZ,5V3T4SCbQaD=d,+:2/XJVaFA/G+XA>IZ<OfRR&.<N4U1V_Y8LO\c<]e5XJ
AIdZdNFY>C^M,QOO#f_WTJ-52M(&N&bZW15W#XYa4MY?c<(-)dCD9_f9aS830IL4
f)P[E1&JP=2[XBCY&E1Kd.^CT6M8>[[9GW&1HcC[5Ca=O1T3B2B73HPDGB,;&T;\
])F]:([L>,H-N=.(5/JIR8Efcc@g@)W[/E7g4#f#Q)-EefAC8AUMC[b3/;^Id.?C
c6P_aRc0/M.bNV8?5OUF^YKR5-)]E&44CB]PB^IJ@MNQ-VQ8(?,cf6e2>Yf6&2DO
K)6GS(,GgaHc88MF;:93F^F^,#)\[&(+I_O<G>F]Z</@3X9O;:>D\ZUe540M#F.]
)D0Lf9Nd+P/GeK)8e]DabM8,cfI;G.2YNI8C/.bEB8D+6RP6M.;bB;M_@,_)IWfW
3G\@cVe,cb3E=RBBT<9].#M4AN/XW#1TFdaf&WCHJYK-SPKO(1f\\g;HI/Uf,7B.
9K1/K4d)/#TO-1AR@OCZD?63a6M(IX&:L6KI@gLK5?b,)AI+Pe#K7NTTY9@=1R[a
YddbP+d.:L?A8#/V37gcSTA;W<U>[A\@[(#1da;XfHGW//>2&P0WU<A=/)D]gPHE
:86cLU338Z0TA^[\8;HFVcZ78P&C>/MT-Y^-ASK@,dI7g.]-OGY9\?<C-N_^F:Ze
68e3&K/D;d.eQ<<9\27BGY=DfJDON<-#5-?Fb:WFe;/7b;a_T=9(TUV7aKbU)PNa
G4^6EAMb7@b:[N/6PTbK_DIc\cOZHTIaHCf>ZN,_8>H:[dfe.JI(c]D-<)]&+aA1
3_aC<XOG6Y8d:JfC1NDW0UO.,8E^;S8X[>dL7K^:dM6D9FI<f+^0^F[F--cb5c1b
aN?fV:EP1(LfY4JWgS5_970<JC\M\W\9]UIHI6+9O>^05EQb?.)(cAOZeA>W1HW3
<:(T(ZPeRF^=/.4]@J1.+Z5QF)T_3>78eC>(/S9=L7a[,)NH;2H-79N+d,BZZAf?
JH4]#FIa4Y8HT/=[-;M(Y\(&.SG[/8>O3CF41+ZQ[:)._aCNYAAI::^><<:RdHZ)
P5^PfKg42B7A0[FeW,KRaTV8V+GEe^<Xa3YIdXY^L5KgV3?QOMbgeADd?OaQL@YV
17AO.ZHQIRaLRI@J6FHB;^.,XR)+T1[-7-VCHVV@&E<aG[)g>SVQQS0@R]T&:,1)
<dQ8(_#<NDD_.b&eZNG-^L7QA-FNSbEE0OJJ&-c3ML\4M1_KegRX9^H0V+N95,b1
eHG2A1EX&^(2ac6AWe942Nb#Eb<6MaNLbK;[&JJB[e0eHOOVM(gO8b#P=cCK9+1;
IObNC2d\C>e5N?SBE0^6=#.JZ6ZJ[U_Pc=OENU1+#UVS):UJ_bM[3TQb)d#ff_#5
5A=cA]e^Q9W1KE,&>-U-N&D\^T[E,QAT8V-UX6fc/MQ&)0,@J^?e<(@G3)2-B0&Y
[cO+8.I,1],-Z@J0<dF(B_XGFg1[O]X0OT:Q=17dY3IPSG,A.^NaKfc5CH(DS5PY
3N67:=5V;AQ6K>L-&gJ7F<dMcKL<fVOf1NbKK2=#UVB-PQYQ+VWE?JAAQ,7C.A^]
(:FNXR7/-A(aLF#e2,P6/UaRCUS^5K\/]>+5EB<6-&^OS(TfYVaWUA\ZLECSO9F,
XOFHc^NA)\.C;ebS+G-GN.S)@PCa6[H;,eXWeb0@IUIg;])ZgO2OPGgR[0C5b-,c
IOa/\]2XTYW\AcFQ,D-cbJ-+9WZR\S@5<V7/A11#,c(<1S\FVV/8UOc564X\Hd3J
c#1=ReWFC:2;A[:94U=9J)P,S=Z-16Eb)J@3YW<S+&_W&+28#edAA\C8E+:[207@
]=F4U>?4?4gGTaY@:NJH(S3FCF2Ga?V0+D9>)\\#b2:+C_1K^[_4B2K?3;>W1K8>
R&3L&1IJ<A2P.KL/&<8FOS;?T]eL4-?9JO]EFd[J7VfF]S,CLWQ/PEPUfaXdKX5f
<51_<aYdAdd,-X^cAETU7U?RW).[I\G/T,fUe:^ID^RP@XTbQZKA:/Y++T4BbI[;
U7/TT8LSK0GPg<FHQW3F7E0JVe0fSO-T=2AeTN:Fc.+b11OZQfPYaC,I2B0c/<Y)
Z9e(F8?-9eX9)[)A&^18aT?AKCU)f\P=dT=@YMH(]#3?SQg1DM_#>XBd7a/aTb67
FbF7N#+#Jb;>YEMUZ@V)F#2c0MIYfFR\5af;PDH;&,Z>NPTJF?[79270cF:QDA5)
[9:d+-1GU^F0e(.g4IO+?eIB=1VYFc2(E@;AR>F.H5Y+F49LYF_Xe:QZ)\CAO3&;
E61G@GQ+T&a;UK<)<.=Eg(6^VX3B@H2S@,&U<C:cW#+KY5G\K(TP(R<W+a[OO,+4
S6ec2PFbWF<LDZg>eQDPb8=HE4ZdAGU@Q<4Q7\3U7,(EJdVbF]R=dQ?)5e6UO16^
1fRc]B9;>c+2TWFR4JAeSN4^Z,)PKMYUBWO+V#W/F;gD3MCP5P#]80&.dE+J6Q0N
=WC7WbMW@0eVGEW[D2H^Le8Y/EDaZI]0T,FT;_=U@=>Y0[E?RGEXNfOOCbbIU)C(
;e0H0XF@C-g80]&Jd.S0^c?S_[4[WPYc\2dBD7\ea05/53:_M8QA@ee+01\8S+@,
ca<HcX\b>OUdT8,;MXO9A[0B5?_Q;ECgH#=)\D/3_;^PZb-N/;FFQ1FOdE584AK2
/[<MV7R)3S[DQ^8N>Da^/74a-O1[8Q1(4\G\YQa&H^N[AX&(UTJ6=GZCGE=N@F1?
B_8caTVJ[7.>MT5BNdAfg3;8:-K/:ZaSJQQI5E;KbEO,.gF)bc]e:W^]C>YSA9Hd
I-g]76LUF_Ae8H;=G?=._+84RFF>ZO4bc([(2:/@I,JdcX7YUV&&/[W]PUH]P.A/
&B@9[H@#+J92OX60W[B<d4O>@2VFA6+T0=2.T>/?KNR#2([A^d2+MFd\#B6UUUNa
<KZ#Y2Y,.R55c05GURQ7(OFHPTQHDS[];HS.EZd>2&d-\>:B^78Qe.F3C;;N_.EQ
e=[QYW017M44f=b5,S<-d6Z5.]>I3QLKW(39-Z.\//U80MFEHOeC[de-;d(7I=?@
PY;gP2gYX730;8QP84TbZ][VDF(0=>T6gf]E359((R_HZ+Nc=Y&dDV&J,@H+&P7N
22#SN)OMOU&7ZU&#7Z,1A\\8E(\-,3(6fVG^QSE;QO0GRabIY;5@?ECFNU^Z87[6
O]bc#VdD\_,Ge13Y9GB4+EKPfB]ZTe=9&,4A5QcWR?(EQaI4dVBVF8<31[)I=OXO
3E_F6.N?9/W)8gV;.+HQ._cX3=DJ^8_PY(D\:[2;/]H]?,/BU/N;>XIT:f=DD0DU
D4D/.RR20bY^PC@+IRJU1[&,2&E3/\[+GB92,?^aaf53g8a30Q44MTb#0I3;?A#E
CH.)3ZVUPT5Y[(2^(&HWWR>aZAA>>.N_EX4GFNJ8;2GR5bYU^KUE[g5d6<BP?c8W
S+,+-_/&LeB\b9b3BeP@PGT0b0BBWFD;.X6MQ4LYA,(0N@T0fP8fK24cI5VWO4LC
EV87WgbD85\aa8Y9bZgOXKKJ+03UA@C#SQ\YM6FS>_EBR=FRMcb(]\4OUY_Sb,IY
E+PJdPaLI/KOgM(a&0M5P/TX:Hd[:R90_UGd,[(0#c28X9Ce5Y/XP/GDe[NO0CM6
\NT_F3@6RdWcT8\Dfb&Fc:M4S,MMXKOc3).;0_@3H2K4DOWA5?&;-a>ZeDOgQ>CH
UIZg#aF1f7SD6Y1)OCYW^d8AQbIJIEH4&0]6[4O;9II-1cT#f(4J(#a.fX_YAR)M
bT<SeSY^]=]DLaK595WCCPW5B?(R;Y4)4JD@@Y+FI^PD4#gJ[L76;9O77),(P1PY
:eFMPCPJ&0\FY[^QF?X0T);&AV6Sgb,>QHGK3Q2geWC/2:+^aY>Xb?=3I8A6b@d_
(_8IP[=&+GFLR><Z14=Pc#ELT>&7Hd?U-:FfAU[Ybe/<F#GB+UO,Kc_8MNTDZ2[&
\8Y27YC23N,OL@0LaP2Q4W.#TVRW/cdfe1A6]&Ofa7T>1JPK-AO\7L8a0.Qe&ZA4
3FOa9?3C/Tb.3--6:,OY>R14b;OV@^fZ2,)dYFQN[&ULa6:5H8OdYf[5dPd?-WRC
^33\0]:Ug[=.9Ld:KdYR;_]W\=Dc(I)5BL,RT1SN>/f#JMb?D<UXEH4DN2>cT;\[
:Y;6>E4@?O;e,&MMKYYBXDO77.[1f.YcKM[@3;]=fMJ<GXTd/USb?9:1JJb)]#Y/
]_=2[GN;NP5G0d(YPN;d@ZP]<d4MgW@2VB_/WG@[RbYEJ5][5H#M)Da3LeI?gA=,
A9B=]/>@7Wb.],NMEeS]VObE^@TF/g?.,e(@P=?@Q<)XM].HEI&_#6BX\QGZ8#If
<bA](b<[(.@;;A.9GK?H^8W4cMPDe5U[eWBfS=aPM/&PYP@NL.<B:B[-P9ML^>NH
B^NMH(0Y?Y-b+(M.UL.KEFIR;Qb7ad-[6(NB\f5KXQ4V_)6NJ?S2&_X4]R@dNXd,
PGCF;M_9Y_YWK&-N+;e]U:(^WY:#)AQOF0?BCBCeKacSX-[6/)LF)OPPD,FI7P7,
0+7SNL]d-\>+cDYSYJXgBCGL<_OPMQfA,IE>dE&Y<7Sf3R;3(&#.HSNLU2@=6Z=Y
Q5AZ@#IW2fAB0gQ0M.PH/.]Mg[Q2:3_=1a3TeK+><.DOFW@>V.gQ\6)2:Y6[V[9[
Q-@MY8NBWfC=7W.d[TcH;.FY3O9CB(WaUbaB8\Cc]+U3/G2&#BgI#7_1Fg)e5F]e
\adV:&(&N;<@Nf0E8?B[Z33W?#+(,.Pf0V8T3-3E+Z6YYN,VRP#H3V\N^bG1B[=8
+X^WHONX:PX&<:)&..MeBg#JAODFCff2b^d)SaK25(A;J[7eW^fD)Ua/N1ab0^TY
.]]bb8#e\NDAH/:_L]?d33cD7[DP-S]_0/@63^;T^+\HO)8L4JIO]L_S/DJ2&V-W
1U<15Kd8).0410+;d5?T8?JP0B[:Xf#K9CPCTMO[f(;K@XG>?,fO15Zcd>Y.-6Xg
eD,\)IdIBNR61G4HS/8>Z_R60((a@=>1eP=FFX\VY38U\8WX2)3TWa1c]8@\ZVP@
_H8RJB..9aBEJL,@<NSK&&/PO\Q:0JC1UOR;Q^8)3?)S/Z^>M>Tf91#<U(_5J9eJ
-,=\aW8(=FYL=R]95g0(Lgd>-<(eGD)2;cT^47R<3XD:\fcS)L=g&O@Z\DJO,3WJ
cIYQL4)2J4(-J?&CX+Y(3UQ11AE3SR)PI;8W5H)/^;J8-\>54g6HI/IA;>^1eN0_
cM4UF0(4]&P=FDI];Q^Bd#N6PaKJ#?_:GET2K,.<SSGB,G\K\I.-42R>O@.(I@W:
2?,.@C+_U05[>^#CID9d?Bf\>Q,[@7;D:&#T?257<GC_U/;aH&W7WTf-PG+&]^Ye
13S7P^[A=R7KDAW^2J?7IU6/&=aH9W&_[N.\LSgbOM]X-)X(_OXG733KP;RZ9^4V
J1=G.,,e#R&_FZO-[Z0L:]f:bd(=UbZY?<&6C/E]eb<J@W_W:XSLTaEK0?S/D<a-
@J^)G^fb&\OeWa[JP3@aA<?cS]?VJX-LTb@QTURC8+MM_AI+N@1c^B>;02dW(]](
cW_;)W\^\4[DH>H<e1adcAB53ZOD+<I<^@1:(#ReU7Bd64/MJD_:ICL&8>/XI.4J
AL[E;a^FbXFIc6PfXC30C]M3^Lb<6,[9WAYYg@-P],4H8>EA:PRBQ)6F06C:/6G7
7gZ0[\&6f&JZP.\<GB:-D?EcS_>,cFSXf_#V<_DZXL<<06T>bEPSe3Cfg9Z3Y.F.
gbCO?CIC,O7L?TF9eW]>G:A@;#)DO(&4fA=/]IA,CW@9I\4g,_T2AQP=a\_^R(AI
.e;G2;8@FAQ);.bAK3gPCVU?TeA)+DK+0XQN@#P:.CQTCZ)C_P#J>c4EX#..=+OZ
3b[O7K6/MfI^e]+aa3:-SBZQCZa^aC6#Z[,<d0^f#4X0NPAd;cC\<;&?^>FUQbO+
fC050M?-B(@TA#9Jba/]VB0g,U2U)6<&W2IO+7VMTf4L2AAC[c?=-G)c_QDX)I&6
M91TTHRST+<11]B)T&#b\M8HJ[77A_A@:Md2BWB7CZ-QX2E0Qaa_&U.174X[QLac
dYYYHg<GU6_[-][Rd1gaXDRU]J9Ub1Ya:3<>g57<4Q,/-@7R8L=)SC+@W)@ASY)]
B,G7/74PG8S(c1T7JB\:fR?F;1cM/6,R=f:ZB+L8^I.I(5gYcbT2^N((6C)OA[7\
PE>AI0K:D<99JQPB4[WKT44FSR/(3-G7\^;bZ<[_V=GA+MBDbg[eJL?82Y^61e8H
(V[:]>ePOY#NMT2e:#eZ\8Z-DE(&9Ra]OZeXYNJcRT^ERVd7;IP2HV]8@QI/1?QH
c56A#MI?V:-cgc/&cPS,-T?-<@2),4bM=a,e8W?dWAdD)KDR9652,GAT59@?A\4-
Y1@\KURM-#fR-VT<K=#d_@)VRP-_T_e1845FF#2-F\@B[?&:61#[f=TV,V=c-[]a
Fab=cXZ-1KA#5=7Ce,#EeO)#C7PG?gC.IHH4[ZXTLC:2fW[]O(^(4ZJ)b3F[Q.c;
7.V(VRURNOG5a<OCR;>Z_^KLc;V@XDIWB,P=G>:H)&cYTI:E@TVMaSKd6b52)ZM4
(>M]H.X?62P\NaeFA<aDRTVPG5C:URd&J?5/#cc_555^@)Z_A0L>>E67;I]^LP>:
bW.UM5:K08Cg>FC9aO<Z:2\I6BRQ6[dE&9/8a>fe>&f)N1[,H9HIF3fUBNZB2]7S
ZG4b4T6M0]4Z[&TU>-&5]LU:5LGb8d)8;HC&/PU@]A#\dY1)DH)6N2L]X-]]\g\V
FJR+B1.VJ>&^:J\0G+6b-K,9e:a.PCdE,642G+LYZ3C6ce(@CAI.KX=EL?]ZQL^9
8N>fN0113C\6]Q\03\3f4+FDW0J+0-PN[(#:WK@ae[fC#A0]W1XS\_7>V_[G;DSd
NRC\:#F/J]=KG3L8/T@#M\(:ERJ?)M0gZST^T5UE@#YbLS>K:P-XM[G2]bfXY^&b
K/<CJF7_6;F#A8[(_T,>e.f-DC7(2Kb<YNH9LG#K^6AXV<.0CJ:9^[g?W;QK67Q_
;2QPBcMRJS+Bb&8DJGX#bJ-RF_+gd9ecUbS/2#(\AXCPec8_GfSYeA1[9ba)/KBI
X77WPY5?<SgVgKc(f)/_?J\^SK_UKbNYO9bg<g#<;dg#1[Y/M[)]).3\W(KNS^g4
)PQL.;RV2\FCd<-9E](T;=3(3c(c4BH>N6Y^XYK@4OVI?CaQ;L7+5:5PE@8[Kdag
):RQaRWOD-0KGHED6X5S_&NMINbd;_1fF4Ic]3P=;ac@#[K]:JUA4ANb?b1F;fA>
(_J@H59@VV2O^a0ZcEL&S/X[^(_B)Z=IGEL<N4cX7:IeS^Egd/+eP1GP++[=C:fV
@f;V+eZI,;1/6/+P\1ZE45UVAY0R)2@QD>G,DT#1&+_\^-aaUAFA7F+1^FXGb5(V
:7I&NTLF134+@bQIO]O#H=fYSG7S<_cGJa,6BKf_J3LWg;,0fU<P>^;^=/23A)bD
aFf-H1=0,aSUcQ((a7JGP4@^:)Fe??1M&R@(Yf].802M:<.c,aOP@fOc,(BCSbTF
YZ)D[<-J587#;40Y3g40a3JH&SPY,DL)X-S_/ObU=<RW5VWDSDWfOCFIZIAI4EU4
[71gY]\9@G<B&)e:(Led@_9eI1&\@e=A.+_8OX9S<BO(Sb;.Z\[E#_)0V\e8X?5e
f.dS]3VTS8UIZ^&>CYagCeMcKGC#Ua]_,XJaTGXfbM4^],<OcGfPBP-=:O3YHTYA
6GcO0P/[?2EMGMdB2[PP2//2FPfLO0OcZb8\8=\=:).\Y\;aa+A3R6YWN,Fdad;W
6<f7MaF[Fg_\bT,Y3b^24JG(a9N+XF+,7bX/FB[F[(d&Q6V<7fAgM)_a1bBbaU):
4XET^<+F4-L7E\OKdN4/G]I\Pd2AS5?EfKXU>FXB_\[;GT0f@Ubg>#I;&N.5_1c.
afd)U_4bf7I].TYK;\5aAMGQ06#Rc?:TC<KYLL@Neb/-##LI4?@=N(=];OH)MW5#
E/P:TfC#]C\+FWe)5c\73V[HJHTR:(^G/^^8=A@FQ.JD7H8H9[dAUO]M9]L>R7a=
CLM+XI-;YC[(2V1D1bH@DJAIO3(S1Y<f68_98+_?Sa;L@JWIcKJ^g&D<G@ZFe\g#
KNYVQIF\DVe,>F4YXA0##LJ.:U0[?RcKW3e36(bDda]TX;Jd9:>=V6>6+.ZYO;3Q
D,T^#.:OYad&S1Q<cX;a@O\7e[6X5ZDHBGRfN-4SO\OKW(1C))E;8,WJ,-e\(Uf8
HVIEe4P&<SIGB(@2TfX.b.2DR]_MON;)FO#^4[5^A?eS.Y+-7@<aD<_O5YGWV7fQ
F-8#V)<SJTJcC^?,+dH(TX\]eO16):;<MaOV4BgaWNQ9cD7V#P7QSf7&cV(?7?.M
TVZg3f+=B@;d\OZ-<f],5=7FOP7Re9D\.=;Sa_28Qd2EO5a..M8<T81KbOLY6//5
^L?LZCA@DMQ,/M9Q\UF@C_YK]DbeKPL3?>bFAgBQ36XF2AcJX-@3_R4e4Q(/&95L
SdC(&U3H4ZbV1SN:X/)@0K\4P4a9ga<+;@gAY78E)W]CQ/V?9AHAW]C/,(NVcc#B
@L)[IW?H30g,ORG]GaCC,\7P9WPB4eXI8#\/(YT6MJY9d?Z)@L+/@+SD?F=2.J+-
_0->@&aBVQ1D>\T:)_;-9g_=BEDA&,<7MT2M3@e^M-EdUQP9#aI^>:)\V7NO/?5b
.S&04;S_Z]OfF,/,3feeA#faX;67dcb\<G)5[IILcHS-g,Qe#DD2XOgZO=UFZ.=f
fe(:#[0CK28/dL3J<EQ\Qb^)/JEff6R4b:Qe]BA064\3G1I:FI+J:G_CIbYMIN6S
;MZ,#0d5?W1d99d>:8U8H+FTc8HN^\I#4+8T-]OCDN<.Z<-5YYWO9LJ+-^I3g/@=
65:3BKFZe:f\?M<(&[&]CK<SJgI[X)5OOa\+2D>;II+(V40cWaAB7DK<W8.B]bVX
@J/&.REFZ\68VXc>bXD\GX+AFU]=YaW02PH/7@]332CBdHX@A<^#d[XOC/fZC6_;
3g4g>U@U,A6XK_8\J^5=-/\IA&XB/>(00,3,9TY-+Ne=MCf2BNXS[e.5,c?eTW,F
&DUSaGe;g+OIR@HE;afMHAcQKJ#^E+WOR-V5AD/_9Ic^:)#9E=G-KAF\Z5]X0](+
Y(T1b1@<eJ:P>?C./ROaI.SLZVL1FYf[\=K[eOT[DXQE]gYf@bG9JWc<Qe^JHAXJ
T@<4L\FJc335\R^@]B1ZI-1#<S@S_T=c^D09O#<g.3)W/L>FcU=bf;?<7I/AG-:)
TEY=K:F9g38:EbCQNNM-<>;[:)RV.4Z<,C<DT\G^AUYQ6#E(=&_5W?UI#.<dU)<;
,9FFO(cY/4.-1gIJJ@F\[B(:gOHBU;CG&UW0Pa+I3VF@Q;W2(UH5.+IBCDB?Qb+L
DF[\9X9XJ>.Xd9J\QX653D99D1E@/:37[&ggOffXLUS./;2>WORC,^B?/-2cfFXT
YPRNd)<J7;_e:\NTKL=L?8D?<8f1BRW+P>H8N)f,3S:)?1b\Z&2Xf-<OX@e\aI<X
g[4N#f>L,NMc].ZO^7?AL4L^0#8.)S6]JW?FI=E(J5.0A?./38?=J>8V96^TZHbb
C;QfO&G<9EgV67LS]Gafg;H7=D[82;IRDF_5++<9=;0cLG6Z6]K05H=B@B?TQ/X1
E(,Y(TV(<(PE8Sa.[G95UDNDFd2;EPWRO#TBFXF<K?;>_[9>>IF3[30g&@9c<LPQ
_\C(98BFBXW6;[Z]VN+f#T_@60Q/CbgY_c=CDe&=JLX4XYQBX#)30B,WU[+TRGBN
g?3F]04D3JBAPVa?@;YHUdbN&UU#1Y;/LSH37_b^4KQ>NQH_-92D,9d/^^]_&&a5
M;=F]P#8600d/11cIP+KV>4HGOFC6.F<M-PG:8d?[<T_@]_G9I&O@D;+,#&BC+eD
PYLCKS5LPaT1BH1aA>g^7NaSE\/YHY\XCNJXU62^eBFG+G8)I.8gN#[G3P_V-BdY
g05&b+Rgf=CF(FC+gNQ=:?7C?PcE.GP4E\2)c1&?P&CHeZ&2eYQX/FO3POYWP3DT
EP?CV)L(&S6YJ-3PfSZ>KCBJ+d.e:cAUY[)<aEAS0aMMP?#3@E#.W/c-[W=1dE1G
d>9V_=(YKN<T-52cO[\8_.HT(5F</9,H9dceJ)d3IJ)g+Z7RKTa3\O^DW^:.dZK8
<8B</HZ5/_6B)gZ56_5(Fe7NMFf_QQ^0R:a:\Id2gOX)=\4<TX59POMCV7#&XH^)
/RJgEPg?Y7f_\EJdeg1[46Y^BXBLLH&J]b)1NFRW@:T^b##Z/N^^AN1=IW@[,Kg8
;LMP.e\Ja/BJIFB\Zgd+1TeE+AQ44+ZC1aA#=>/LdFc.Wd8EA)I-P_R_24NN)/X]
..M</Vc_I[Q[D4F2b@K&3^:-=++OP1dFB?V><;8\2-3-[C;W?[dE1C,K@eZ-a[J5
J_,W@D&US0N?X3SaY,)_@+,<68H(,8@=<X#TUO)b2&O(K#M4ZW]cf(H9KTb9/VCP
b2XR;]6(W:A6@82S=b:GI5C_TAQSJXJBH&;g/eET)9FX[).Rg,Rb&5TIHZV>RV0C
UGZfLJd-M(eHA4,=Q&?@)feS;=9-cVQ[)<7<\a/FI1_C100P&-;FgM0N#2:ZKV9P
F_2H1H\JOXUGE:ReO0G:DWU(O(BH)RJaYJ&6S>9^cKIgGTTUN@ZF;^eJTf2;gUBD
c(^Fg5B8WWG+,/YDVUNgYWQ7SMH^aDABg\2U[>.f;S6KXJY7G^c^^dGU4_9Ud/,Y
Vb2SCdFYAY=(#+_R;QdZ]<-Xc5D0_,X/QP^TYM#.\fAGbc-^a-7F;.V&8Yd\ID?b
&d)U\KD7JKLgC.7+=B\JV<ZS+=:K;T-^B&)=<57GP8:7OD3T.6;^ANM;EWE([ASY
MZ\:D@<;/KV@^3+&=<QFK4caa;(f<VKL=5B@f^a=U_?]2S)NG#,=9)8ML@\gM,B#
RLA0bP^,.N(2#>MXC+Zb1JZP@_[XZ5c-J,PA-&bQ#KQfWef6XE.:I:88dPM^<3)d
DedA3EMT7E\;M&<dF\;EG2KTg=>(N7N1L<;IW?6[@J9/-5P(GH7:[&Z@H0\OgWcH
-a=A,2b3C(IO4NB>b;F\+c/Y2Wg(f0R3((RSN\0[R,:K(2b9DOP+MS8aI2D.&NX+
eMRNaT1S>HSZM)NOJLPCVP^d?a#4a&,)XK@_(:P&\HA.@d8MT2)XKD;++QPACWbN
3;^c2U0P(72PIZaN,W#9gT-M/E71,G,1?KJ<6+Q(BG1NOLH^Kdg?=^8L57^KZL;D
=DIgHe]dE0I9:;c0-BGI2W-8,R]eS6C=6)=YK9CL2aN3G31a7\][LHS]^JMO9<4Z
#/U8#<A&6Ad:E-DC0,LTWUF8BfIJ[7KWM4SEDKJ./FT;:>QJgXG];<)JRGBUdKG+
7Q5C,bG+K&/?IgX&T,cC)&bPYF]QY)OLF;^;@6QWFC17e&8?JB<?1_2A&2DER<\?
AUMOd)R/4@D:a\TYQ5Y1Q[?M50(+T-:3(Za^G3f:-&_;?6A1)MH\:\UK#aS8#(.L
c5[3ERPabS,&Qa1<?<C9bdD7R=N-LU29(:ADG9NMB,1<BF6[#L)\,IcW3FS#EULN
K??/<_[P[Cc7R&CP4DF[ZNNGO&J^RK\g#B8H+_/.WH)-aIS#6]f;TH2V43^aH1X;
5TSa6F::/P-49X##<B_/H+^H\S/;(R+6)9;>?^5?N^UUUDf276FL5A.ZYFXK>UG9
P-=1Z_Z_S)R4+JVD7XONH;9)>]P7/H6JYS#ZK<NVc^1a?,cMc5J_B\#667.(5_CN
5cKfFcJ<V8M0I//[SAROJDBU_DIcY/d[7Bbg]eH9eCB\1e;,BDZE\P]e[8].ZO/#
61E6\.a0#LHe#/b=BG\&I9>:4J4O8N4CKWXX4b94e4JI#/@^V;P-.UHMQ:d-bg.Q
M3:-7<I+@?O1eCB+XD702+^/Zca38NcB)_4#U]ACgHg5,:UB8O+OG4/-,I?YRG1)
;cC1[MJ(Lb#AFa6Ggaf?F5Z(bA[KB0_>S+NLCNE0T?a.a\=d3dK=\HYR9AdW^C_e
Md^<>8:,VKI_?=FK-SV>SbE8.,N]Y7,I;0CH[5?Y_G_Md05Z9dM,0M;d;bW;1[0D
NH5M@52f67RHZfID=;Z4@Me/e(TB]e0GD]E&3cbMW581<;R1acLbYG(Yd=RgZ&YO
9>C+P]-e964Q)Bb@/LaVJ2F+8^+JE8Y2IP4L2VAT])>FgJU?HSW@E<0N5A7#S5V&
);1b.0HMAAQ)0H?FFALP@R2gMF1,V0IE8@6F0HWRffZTQOFda:8b03XOe0^]UP#<
7/HC8X,HO40U0Od.SIK@I/2M#WH;W#(-2@H=cccXcZ&b,K-5S;Y9N-Jae5XP38;0
+IgZVd5M-g(fOGf;U9@T2BHQ:2<;=(9-O\>):#,eZUHFAW94f2Z;:#J&af6U)-\V
^ZbO40?]_#^Xb7CBU,ZTTVTX<\3D\=N,64QOfOT:IKD\ZC(^V9&07U?Qg^Y=8T-X
aHZ/K@#g_5N#YV8\=ZL:D;<6#9YLX[UIQcZIF[S)<84EA,NMSHP<:C<NV\++)^0f
AOc>UD3[P?c9Tf:LMe&FBUeG=IRZ,CE_F[4]fY+4P&(A^H/GBTa6UMXd)dE);6<Y
&2AFG+A)bMbC\9EK-;6>6cZCB^+\XJ4Q?.\Rc0/O;H9Jd8R9+4LS.(\6Z<PF&&5#
,&V-:fX)Y5Md/g__FTYb:_ce(C6[gP2=09daAVf[HDEF/6I/G+3.\UN\ZTA73#XW
CaLBV4.I)gRA]1b#GL0AHK336UY1[,>#QF3E93Cg,G6ZZ:MK[G<L8SQAQf:C[QYV
5CA,[N7P[f/UffB(d)+:]U\5BMW1B>LbW#Vb\VT<JbJW>WPec\E)cdCRWa5+a3RA
SbE+P]RB5Qa(dO2=\94PUdNID<?A+QA&^#KeQP+QM@O0JFE=]C,32_N&ON4&B)eF
@=C45P,<D>XQ+Yfc4gHT0118<_B(^V)+JbMSN&eM0GfV4VgdQ)[38c;=c>BR9(AC
8CMaQ;R;L;-20YL3RAV6Z4GU+<d)g>DgB7cNgH_ZNH3H+U?V9F2TaPPENLG-.:QF
NKKDI>0N&9Q>N7Jf-E3^d/=S2/;\C34G;IGda&)IDL3>MM:-Nb(RZQJZ7c4G+-Ma
ZKb>#fQF=4>N>>L72)W:?_22]N&:6AMLUM(W6QSR\[G^6YMUgd5>FSGSaTKM:ALe
#H2EHdRGcVI020&GJ=;Z_U[DE=c2Z3)JLa(Af&KK82Z(U<)b;LYRL9#I]6/eEY+H
W7_f5b3f,HMFR_GCeAOg=H8Ca0eDV2=.DJ5>]6YYDN1J)5@Q?NFJ+AL&:f9,5C5.
dC^XbK;7WYV[1gBbUM9E,0OddEb4[H?G:+TC^g][Z>]NdfEE,c^CgKP]egZZV=^@
5W^a\7ARg4&f@I1X3LLO4ZaWDW5,[UT\,[;[aZ=Je=&Pd-E@NUYR&K19SH]:92:#
geO1YW.H(GFGBNO&83L9U[X6]O.YW@QO(.C,.)9Sd3?^VW?J/gD8+8#dCKe)9[4>
P04=2eRg(&:c6T;=2=SN^-Ob,HGCWC1^GUT1S._)(O)c_,^bLgAM&&W:edGXQHI8
PHZ>]VXXH5=H?[8X.B@CU604^05acV#TaHXe_c/=&ZRKWZYA4@X,RD(PNXJJ/^#-
&E(B;##JF>9AU?+1G8KZA_T(YGQ.A2RgG&,P<MZ^A&eeBE[(b/@8A4MEeX/YG^/.
F--AP.6J0_RfbV[5<ROR53<8?BF6..M=P1IPQ,YVETG2A1d.\:PP:dV<S_K(fNYS
8=W<((db+)g]YQ,J@_7RL^9;^WH9)6L#4?,X#[5QEcIV14?XW[/-BOPcaE>&g]_W
/,Z#(;>./c(20_cN&<=UE54T6NXVVF=AUT;1W@7Q4U4D/Z)7f0VZ0]HVbW45BUE7
MIdW,0R.L)I<K7;,#GMDTCae,F_G40Q6Y-(@]3_M)SNgbR&>=bG5UDQ==f<>LVBf
-Ue;SO2,L46S[]X/;[aH51cH7g9b-b+c;6^8;#SR79[&PS4e2#2GR)D@T>0<\b0Y
f5T2.3-PMA(T,/^I#S7(-VAG3<P_?Jd7TMNac2#;5S@-EeO3ge6@3JXM=>dWMZM>
R.XK1\TCZP3ESPa0U9T(=G[b(.)<QGad1KfYZC/5:Y-f^2.]3)D+I21KS7ID12#7
g2+6Y^M(4DD-AZ8E1,PS&WU(M)-X+ASg]4+N=9^O;]@SAf-;C_B??W)1;AN<A)71
:K4)P]YU+@Q,?7_]:Z3)K_.d5F\2a5&e?fIcJ//&2LF/>6@BbM0acPCUUIJgGPGG
cSNeIT>9,I:VRI)ZPOKB0&6(Q9(?/(UDc4&VN[TXCU:c[b?J8eB@)6NQc^a6dT^,
e&Oced/8:5/H=.B1GbWJPd)PdV)\6G+Z<K&N?Y&-X[Y0B,CQ;7WV,],X#Ob8V>L7
7Zc-Y\\;+JQUNfWD2f8;S@D2-K>:=R&M&T28A1I[+01eQ(^CS1Dc9=bJ3bC^PgAW
&Z?ge49@&3F<JZ\63+dQ2cKf)V_0.0QFH^P:@R_FQ-)3U&K5R1N\[P12d:A)P_YJ
&,Z8&44CZ>GCTNX<1CSBW7Ua_BH3T/,D_?\&-23F6B6>:HR:WT1.>OHaAM8a;AbX
Pf_.8XRWMLL@->a#9XNIT6Cc:?7@3dHb1d:g9aJ<JI[Z+U(g&g1>PV]X)Z:Y.&L_
7F,#^?bK>ca4RW83E7gP4ZI9L09\/@W76I5S]V:fC)KgP)6c7&Z/#1H_UO01UN;=
J98O4eNdG/FK7OgILXZR2?/XVM3g^.A.eb>DO:UD2.\DQ22LSdfJ9CYaWT:_Ta[K
/S8(F1S0.68>P^)&B;gLIB&LIKQ9.4[T??COBe-L;O@X:SW9;@^R:TREO-6TS[^\
:WEe\?AUOdd3I@@,+]]R4Z5,(fX)R/\<D05Dc(U&(;HG(BR(F:)\d,;+1UFIK&:0
aN35\c#3W.J]M6,#Q9JGeO#</)J]-C?Cg&<Z8,=[,I&fa0-g)3SG/f0R&AFZA[AD
6c=8==gc0=eLE7E36NV]b-#1b,3TY0IZ-G[[<WNCg_[)3AO-=cLb+DSMEW_-L;=6
,(ZEgOY3)8Z\[._B3,.5KfDR5F60+?g0I=1;4H](Y@,0WZe,OJ^G3fERVUWbOXJ6
T)bY(W&7KT)EgDI=5/&Of-X2@<QJG5.>bR@.4LfN4]\-c.^-RMBg)3S7;/Y-,K98
JgZHVJ7c7I3d?+Z1P-aDZ1YMb&OGO98U1gVWc6DNQ_0X[W3;O\ROKfK^INKSX(RS
U@G2Mg0<T:W@SL63+Q3<@aLO.ENE8>_U.14b>#IMgc(8R+Dd3e=L97?0c;P44BTb
3&Jf/2WLQH8e<G34;9bX2IM3S2[2A-DXU3L&;;)99ZK[T.W<7-9Y4V/T]VW=Hf?]
cQJ[C^OU6HI(7MVX0CT-1c8T-^GQM9187>GPBT<J,^2A&\>bX,V?GI[)O@YBJ)92
1@(EdH3Id<8A6TM\\2@CM;d0cK=KI2J[L.VfC/C>1g6/gKg2XLL\NNYebBWH<TXW
>/.b#_K0XbG-f)<>@3Uf5Y]\8b/JF&c3SXD2_@I<9FdM-25/KC7DYH&AH]e2RGF:
O(4=<f:K[AY:&MWBE+c,WNTfTaMaK]W<R,0e]4IfLH3=>O^d+W4[J6:DEf.36HY?
Q\61ELCf[I]UH#P+J086/\T\VD&+P.7Kc<\B-d.BQ_637O0,:]E0@.#.E_0eP01P
aP=L:c:+AN5\,[LQRYXS;eYMaBC^X,)+HXK0G,6HBL=gScIaO/\-QJ?+7gS+:U)+
>_a/b9c)8+D&&?XRL(@TD\I/):8I9=S\:3_=?0TD2Ob&1-?OI-,KCQT8L>F8YG6/
#K5J,D3A,B8>^0BX<<,8))=BCDSeZ;0RX<ND(g]?TG4:BCPd4CbNH66S\<c5=L-,
Se@0JA8f+90:R@eG3>(#UEZ1KJBWNb15F>HcIdLSfdQXCdISa\=5Y(5=DA@URX7c
TJ(6^8U;S_c;RX#<NB=L?^@V/de[E.IOQ(JS]UB0bU)-ZeSJ7S7Cf57d83a@L8[7
E:ED#ZDe,2KA.>6[D5H>><5_<EYb[6Y)1FH0c0H8gRPXTYI_[+7U#e]\+3KU(5G^
)#&]K<aAVRGNTX[.S0]#]C(PTc7X2_28gA[=2:.^H:g6?#>]Wa=?]+L?Z\\b=+C5
4f7d1V<.>-c:E+Z01=01Va<O7#TO\T[JBE^c#8AQb19_22b2.NBLH-SG_=J1>LNT
#)fHbO./KdMGGW3C[d&H7V2/)1>Pc3CAVD[_Z,#Uc+gdI7fUN/Q4E4VCJ2HD/E2+
:CEWJEfT88IHSF?@E.3HVK;W^K[9cGfPOBR]5g&1S8;ID.g6+dNC:)3ZLS6-45?e
\U;NNFOVFWa:0cU^L\L9^Pd+TPZfC]VHJ/6aEKcF)K;_dI6A#U+T(F[cfH:-?Y^E
[V:3ML1AIb9Tcd)+<FP1:SYcT8/K]4ceS^K[/#2L&I^>/U-R0bF:)C0<D<bXYCVK
,3LHVED<BV+5<5a4#D1,=>TD-0(^#N(T)W1G3_,>CHWLDA1]0+[@H+7CAZ4#<@dS
.BL(gZETO[MB81cLa:TSfd8WDRMWR35D\eGMcLB9Le=CXW3.YG\\89]&Q56A@7OM
JUOM^aYV((\XN#&D88f@RDE)3d48:0TKO#L6WOb?P:.(RB8^.=NEZ]>U,6bP\O0b
J+&f1^[c?>A-ge[6VEIBUc_XV83CQSKVgLJbQ;5Zd0G#<acM5bM=F&dfJQ^,P;K=
RPMA.&]HWB/d5T/DW4#F<a,DP=3(ZRK=TYd^\.6U=cTJ[6:SEO^]7<OL]VXN(;=R
c4cU-M>=c\,>DRg.?fIX=@PN@(49^-@H-&#I6N7,eLQYETN/4a+Z=#_V=bH(0FJS
F1SaZKAG.gW4:\.<;T;U3]TUM:H^;N6P.PE#;HJ=+M>2^d]5@P6a?N0^JHNdIW2X
ec^\3ME+4\-^EaUJ^Fe<WJ+W9\5?A9\M.P9J9a=(K8OFT<S<IMDCRa)4J1a51[RI
Re;V,^Ja4VNUITM9bEO3XSVEKS-X+?ZS90-g^)\U-)[H7I#S0-.].A#D)7FW\aA5
BPAI3CgTB=7R0?27IBE,(,JOEQ-_Xa[:0E)IVB5fDM?c-^\Y]BNK(,2W\gTId^KT
KM@Nd35P]J[8Z7cG7ATAZg9:YU\PLTP[=Q0B)B:(/2_@-Hf1cW6UC#9P7b=9O&Bg
FA..GD_HBRb/9G?0@>d3KRWH\U<<Kb4D-(.Ue:VVAO5)Nf]X>V/U+Y.O<?WTOWfY
Nc,CPcf4aA.;eTSd@aZ#)OT1)Ce5gb[e0<=.UV\+JcX185;eSfR.1P?/)&1W:G#A
H#A@d@NWJ?)MHa_;)f#>G+.+:cCWcH;.AT5XL#1(R+HgbL=b@+0S@MKN=8Q4eR(D
(-S9=I)E^L+7+7HRe-2:Y39F/]60#5?9ICK?a9?+IeOJGGV,79@SL6]LMO6b4[fF
bd]F>:1X5ZMH[L)U^Z;6T[7d\OPH&BVf](=7=@eQA[/I6e=d&4]WP68<IJ<(Y<=3
(N,R>.d2IK58KA,eBOfITIV8-Y_SZF[FKUWb^KWB6=M.P8J89>+,I9U9]+[/C]]\
I>+Y2e?G<5Rfe.#dSXQM+U6/^Y<5#L1VDG0AH&HIQ?/.:Id\^L+]?0Xf3:EcgX_[
cLB+56)K?_,MS4AZ4gQZM1D@B6.b6c):2;>\WUUMa46<1[c:@@dB2F/17/XKeHN&
M5L?JEgA7POKM?WP)b]^)_S\[B>KRSeM1#C&I:7ZLW<0cCEb82T\fSX90Z2URLF+
bL..I^Q:^NB@S)d^dLWMY=f8.?/7S=UQX[Z(Z.G1#<UfOMMe;FD#.f-f9Xb.A]+B
WA1O5S+<-,YQ^2NOR1Z<6X0CP@4&AF^ee-@USX8<)3<NJaOM&,_P#_VN+_YE[M.U
(D.XI[a>,C>IR:P[P>46B-X#N5O\+BABeTeEN8B^GAW:^^Z(V44HQfHd=N,FDLg6
LL^0;<-4-9ID)_2&XE/ZCB:UY#U)U5GPF+T>],\B=(J9R;<F/4Xd?cMW+HU8W2/g
L\L/I/,V/,a;KAf),Ta0:9\+3E,aXD9G#?814.UJ)AeYW0@F^6IXQ71P?##5ISG7
E>d^/fB<>I/FWQ1Y](YbL#Ie8XQRG]VU0QFZaAaZ>-3J>+c5d\VAI>;Y)Z6+g<LG
@F6JY;[0()Q]#(?8]Q1LWQS:aU925=5))(dd5b_M1)Z@]])13>dR5c131BELcIS]
<KeT+Bb2c]^@\LW8,RVBH3:eeRUXJA4TC&][R+5[KN68H]9EP9)SX9.)RK+a06O>
4B\;+a],5&J8H2/R(_MZ&[=_;P(PIG.Jg5G,WFW3FU+&a9BdQ?\IZSN+&b7aNV#&
92J(<8.FIVPQXJ+3ERJZCde<PK39EOOT(dV&.EBL2T#6bX0Z5DM+G=&1P,^b=:4J
W8d<HH;]O0F2B<13X2D9J(Qf2eY_b?:2SN3=H];g484JE]f7#98=.<JdW(4g?fRg
:G@JG1O6AeP1Rg,;._?5<b2,-Z7S<HHEdTO^)1N>[FU@?3ae[7@=>5EBW?W_,S_@
Jc/-(&d(A/\_.&T.#;E+PIYS3BR8?F4dF2\ZafJOPXN;Jb9.NTH:fUE<=PU4;VG.
BL=NM\gKY[;XD[bUeHTdH5c-A4AXbH,U<ZI(@H9E_a[LG-[9&[R@F8ac(a8XD#L&
[gNNL<fa5CXQ=JQ]/X;TTT;\c^]ZOS<K6S@/DE,B.f^^1De:]2T9XC)Y[CU^69]&
MI1R<eeST/=D_b#LW:UPO5>@17YD=GC[8109&b5.<UH;<gMK=H7dAdSBBV[:D^U7
X=Q7LK/0NI50)M@;>]CQ\KKIg/fAAV(8#,bXM\aLR.EEcFZd5EHK^8?<6cX8YBSe
/Q-,FF]_PH.B-b>ef2Z@.AUFg/]))VdCe^>BH7TBNTKCDF.M^gRJ^c<SCdE5b0&5
[(U@(FZ^L/aT/&Cb:VC)ZGO^b.]\0+#=UEe^FEM1aEe54G_WEdDZ)S/[&DVZ,Ugb
<Sf=T=.8;GIT^35eG7a;N/cBgY@bI0^>=3Zb(2_c#7bB.[&A;Y81/\)L563,#OAW
8/<^BJ_[&Dg_]0@2AS.dI.@L;LQML](JNY/APN0JF[T5T[,4XAeIFU,?P>MT<;&P
G16-OERP+W-X+X_VVGbDZf6]+VC@UBdTQcbb(93[K=-eY7G>g@@;,-:-C=?U^N\R
F_AB(O-b:AI)1N@UX+3+E4fDN5I,1B^b=\e\S8[F_Gg58P4E3K53gF<g^a28+ba2
f./a@8@K>=_G@:Y25=6V/93R#B]3SYeYO<^:SI3YF;G5H8\C.8)Y0Z8;;0V3Q,g6
B#gX_DUME#UbfBJ)7Ed2I5<A\Z:eTLZII#g<^]IH&\bPR,7O@Z[^c-GBQa)4-,1J
d_R7&3e?Qb1#P;7.DXJ&YcI6#AS9N^a6Cd+YQ;(Ea/7/aQ3E=Q+P5UHZ6+O\@X3-
:aYXE-JUH)20YA.U/WM[,[U]9#g1OIb9FL^T.Z&XX9.b7#Yb[=C)#A_MO\??^)QJ
G6&S398JR5::&HZIS\#./0@8)WZX[&9^CWJ\P/Lcdg_#^G.BL)^[E-2DGNME@&(=
G@]:C/OP,]LAS\[_3)^V.>/6.U)gXJ/99__aRN=TTg7V0GF>^Pg(C.<]g8d@@TDI
UW^/ePQ<#2=Of_C7eb:aMQ2R;)/cf>XY2N>O9&UeOAbE&)F8ee7>a>5IN.=(51bA
.;b543@^5([:B7P+eODG1eL6HRS?cERVZ5#MJV[fXBOK<ac[U5)=-O=7Yc:+MAVS
,eJ7WU7EMSL9[]3bH:^BF+)/K<7MGMOK:&FY1SQTba30LK<b8d)#9G<f:g<5D=8f
>-HDb#\]9HTTU=a-M9Z.5bM4_e]BVMbEA)H:eMB\]3?9A,gV7G.(5[f;=R6KBK@F
1.+4ZWe//)b00fb8X,P:N;f95,.B:T#c>J@.M(&fIJ0O_bGDgRQDD6JPGEe3eEG2
).dUcafS3b;3\&1V.\8=\HMZA;-dcY.+Ja^C<Gb.FL8M-<#_^dKc:4\f\G[BU22Q
e[2J3A-+BM_5X>HN#1e[)45X-S3#eK4R+XE,O+c>2#f4[8f5&-:C^2+DZ.J#HdO6
JDeD)K>JAc^>CA16.:],5CW([;3GYPBG/XU1T>XY(#NY]&gWXV>,DeJ.=03?Eeg(
_ACP#3YXG6@6MS1D?HZ3N8J]ZLPbfgX+^?eA_Kf]DCD;EZEa(^YFcCV#VJ<[TcP\
G3ge#f04R^[f<8NBYVDY^DGaea8fP[7C]@U<[1cC8P#V4HO-2Rd&WPWM;\T2gf\1
O=F=)+@Q/2;IXJK\\e>4WEd2(PXbBc[JO^Cf\ZE:TNL@(LGTUP4@)SZ[/W7aM(I?
>T_NM8<(6_)[R7?HP,DK:#5W[#^K89&a@VT_2I42D[,P_0,A#+#=UUAYV@5?T<\W
;C+ESdY2HH<_7e_fHeF7EUM,e.OMJ,N7,@19O0V7N9gdA3NO(b0a^S-+#&908+HY
]Ce2D[96CQ6;aA#UbHcB5;4<1-N72R\44_UD:4Ed;fCK[Q;fU/)3d_F<F9VL,<V6
aT/SDI)6I8:5P7VK#AR9]Q,gB@:Q[81;-WTXVN\H(e)C9,gYEPSK++Q9Q&]+RX\B
03Z^?11S]d(D;fWTON/FQ53.Y@FSXdV8Ng-a:T:=:M@)<]&N0OO,_R:e@^S,RK[3
Z,7<6OcT+3)_f=(28>]5(OE=B=>?O#g]Efe.6WENE;-YQ,?B+RBY>g;eaX^07TKU
6C/X#8.8&OV)QHJ)JQ0E&Fgg;Q7@Y33&9>H,P(bdHf]@XM[U4/6RXATNF.PSI[N_
R)3982YYCIE=7Ya6X?@Hf+JT1YL<-=JQ_b>6XJJ#,f10TDbEOO[81N@S^=+YCLFR
SUBR^_bgW3M^^gD(D9^@UbeD?)_4HWML6-VS5WW:>6)99Q)(Ma&-;>[g=9KfCJf3
F9I>W;CLD>8@0JZ3BdEdW)D?4I,@_9NCC(8D2I52XOFec3Idd2LLRF;0cRg#b53I
P3&Fa0[aR?^,,-eO<ZGYS8UM>dP\T4,aJ?.HM#+W6HETW#J[0?--:4K3>QX#Wa1Y
4M:E41N@H4/Q<L.7e9TRFHZP6W9M.?,X1fHRZ(eMMF\S6<&cXQbE6)IEQ:(2fJe8
E4->5>We&<9)/:CI8?5)B83L5J4[U.:DCcF_0<\f2Ta4Y_UP^#cb6gFEW.-WF[.1
[S@<PKZ-4=MBYRWN>0F3b&4)_(J8M=XOMINgDKBKE9d=L&OMEdUG+7KFKbK75fCS
gS;?N#a8O\W#EQT+cRe<CSX6,@-;?@IC1bd+3R9&A;:I/<(9,g?67YgG?LTUWEb\
4(8E:f9_MI9J-7XLb,N@5\07B<G[EU-_/NQ:[-J[d,-CJE#0@8SU6[,Se=N--(cZ
&e<785YN5e,ScZF@59RX6Y5+2[GF<L8KL<c&-O:HQ0BDF69Rf=([)9.Z)64Ae#-:
?>f-+0_R[E3QQO0LNX=0gWI?Y9;;c=FLMaG:2>ceA7@/Z<NU1.RSBG]).V-]6>+3
a+bW.8V^)W=ggSQVSSD,:.0:>CF)1BH7).Y41,g:W]0&<BT0+RRNVf2N8PQ_BF:6
3.H)D,=5B+3GL^(\U-TYfLS;L_HCa+2Q?+Y^9CXUX5Xd6@e.7L.KZ&a9daY6NCT4
b1a\UD5&-g0MPW<]Fa5CX?]D4PJR[.^a:g5d@B/\:CJA[C2)Y)OK_^Ve>II)-98&
D?Q(cRZ=XT@fSc=Kg+XB&D@;bO?,N\PP8HQ>_4S\^.LCO9/6#.-B02e^4bJ4LUDR
7&;N/Af?f7#(;32<Z=JV/Z)B\&aWdKW88K=,Z>3:V@>.4XC=+ddXRA/0Z^M/>1(f
?e.ML?fDc5SL4CH-:GaE0@ZaTIaP<G]EM>)1LV>Cf=W5&Wg,PWDFO_2TMR=X@_@N
VXaUXH^-O9?K=5E^Nf1>.R[e?J9D];9N?T+#;+_8NbDYcH>/1dVXbdYMFc,/LW0G
a0HQQ8=]cb<A9@MTE7(=\GM#[>1&7#F<OAfK<G#QI>0WX@Ra4#MPNR&H?BSO\a@e
G?^D6VSN.Xea#e+<D3WW6)>2)a]Qd&c+c/d/&U8#DgY\PG<//IWL)4T-b1#]N3J&
@c9Y\S32T&2#@e>&RUW3QJWNACCFK]D/[/)-7<OJN_X1]3cLFLX;M+1,6/56LPdW
.f3DfZT8)KVc>fd\BCQLBd3GEUS0WeR7YF>>)XHQ=8gcDaga3E&ZL:.(L^M[.#U=
P1FYCA\g?B6Fe5313Jdb>dIbA:(_VC]SaXB2H<F_fM;C(5gFY;UgE>T(U(d=B0b:
C.:K?,?TR5;P&@0Ob&]c(XTH^G[;__KC#IB<e@b4[3S4[d^fVLCUdbL=25ZQfRC0
Bb5^60)eELWMC;H:_fXX(@;U&YC6Y)/>O>2R;]bW)Y.E[//]g;=G:.DF[]\8QdS?
V)5eW>_(64->6UDcB;OL-(=WP(YR)PF?aRNB[[O\KI5L]c@+8)1?.?-]/]F0Id:R
)9_.Y]d2?93M4\7IWUBP+&0AL2>,X?V#)R&X:?K\NLY6f/,K70fIXKeZ94#[7]Eb
#:f,K3#^^(.ALW-JZK]/4;[<>;B1G?S#NQB_8M5gH_MR87[)AH?Z=QSbHUG>g&Qg
,6Z[8((beFb2Ag^:C9JM21UTSd8><6MFHLgHR?O=F)F.]Xe;_a/EZf]8_CM::K,4
(&^e\XP.ENF@,-__3+<g]ZIfG>5H..SgEVFDB];GI9_1&>I-:gN97F_f#];SMZ+,
g7#+Q0=DSMFF1[5a0XR+GL1ZI[V,_HCN\9ABZMATNJP2/WOZ:g62f7aN0,W2Y#,:
76#;f[-5(&GNf_Yg;K.-==&1W^I3d=HZ2McRBHH6D:Z(@][WH.EK>WW[=?,gI:3I
bG_3^a3:[NW;cc4\]^4eF#<^Q\c896#))/3<d(WbbX^C(gB1<.RKAP.6f&9RdV&-
^+>KEf>F:&&Ve.W\OMY0g9=Q_Qa(2Z[U\C4+QI1a\_-=gc)_^K42:;N8US-Q4eT2
-daf)B8#fF?2(;Y_;fJ9Z;<[]MBOTb3Wg,YW#H1NP>B(M>K9?2JGCEb<C]+Tc[25
<6a1R9AHI-:3aPE\::?]_NCXEb=5TV,,H]SV(R)2NNUZWL(_L+4;?:<,,;B6131[
Z^^eA5Q6[@G.6\U,RXJ3:4H-3b(__U/7Y_M-c:3RH/8U,d[dABQ)509#=8(<G.^K
5#).7@?4WDY36V4?-&R93-/NV4[D?eZ@)?L=H9dGaa:[fPFW&;>.5F;[WYJE-A>#
NC4Gec4A4NNc]_C[8]<>I9gUP,Ia4NeUD]eP3WO6@ENH#TS5[Nd^E#fY2EZe]>1d
H)g@^.]C;cIXb/JeVV]PT[#fKZ&QM&X)QLR-g(/Q#3#f6L3BQKYF&eBN?&@.Z#<E
J8SePabC=FFKM^0(7&\ZSER3eW&2[(8cV@3fUV<JP#P<\Q&TBecW[F]4C#4<5I?N
C9HGJ3-:?UZUG45gb&^-1,LWN=(Y5\ADQHXM,DZ/-J.ODd7e4Y/Z_WZ9+:MEFQ9@
K8)/0][gH_IZUOYX)AI-RZHVGE<a3K@STS64=(NJF-MK?HECaE8;FXKC7>_N:W:;
N?0Z_c-<SM^QYXX1]cEZL[H8;bB4562+8-7AHPH0&\UJeN)C^_fU+8da[Z^@INbH
GY:SHQ?J->ECKLbY/>?=4)Mg@U6W)D/,7bP8T8MKLTc>5J0c<--[B^>9eY<X)X@I
J2H3>0EW),)W&,AM@c#LOc_KE\,EVQ(eJVZ-O6Q].P:a4.Z.=)(G0=++@,+_#1VD
2@d16T7^^=[b#;.+df[;@9b;D#-&.?aE789GeF;ScYD[b>9+e36I@QQR<M)OOd]2
/GMGFQcF&Vd16ETb9&DVYgcZLZ5f<M(dX#>;:9.]_cO3-O-(I5LC-:\g;NXJO(&)
0&#RT<HJN]?C>I04;_JeEVfc-H#U:_#0OH7f(S^Ug2e?g_b#,;PD3/A)eJXg02SE
52Z\Y1beELIHJ/[9gV/HV?IBL;P=Z\XS>CbW^e/.BNV-6^>T+dED_(2X)0#aQZV,
A51-]a2g5GECA:B\V0O8833W+bQ<B1X_]CAYc(1G[+9a>OaC.PWN&HWZ2BJ]F#g8
MHO&)H]CcU6RYB\4Md5HH6Ee8155HH46SVQ>\NENaM<VW.4N=&\24A2B,KFX\<TI
#BI/A0&/#E<0\ZLf1CIga_X+(VMcWaBZ.FZ<;Se]8D8HYYBe6#WbVS^_-dc@#O31
ZSGgH;O18OLHa=)=)=P3dIBXC3FdK4)@4@dKd.3fIDS;,RFP:R:=&QY]S34,+4b&
69U5e;cLT7G(3Rcg.YFJea[&F/6^V_^>6[[P\1W0+S3H>c.?IT^S38=18f?7aJ;U
KfE4B_ATD_/SKAa@Dc#c#LbYRXIfBSEgBP9(_&6,VU>,CeQ7HV&I8c(e^+KAF-]M
3]B0S?8/S?RVAPRX+4OK(GIY[geYfP7X4L)69ecAQ@3&82Zg^?+)+;gXab1SJ>M<
L<5D1S8_+V1c:16Y4VDSMHeaBa<7a5]AAVGPdG_\IIW:3g@>GPTU]:E2#L?4422L
a]1;_7980&:\W;AVKNXTTZJ[EU#0BXc=e2O@dICXH?SOY+I&,aJ77MEZD^E2E8\&
UPb7OPgP:D/?A7RBb[YVID+c0@c-9Ie<YQ-67gR3W6?NIb0FA@URO[Z@Z)?;Cg33
\d_]\YW25A/.K[cK/9cWPIaWXPW)cO&\,,OB)KYYU0=7>O#W;HS2W)/>_W&8eFE[
]8[OS&;NKE@.X._.CE(c@X+&?c0dFRKbXR+0Aeg^/MLa)]>6H/FAUD)1([5U^P;#
Z6Hf@N\9eB&_.\3BMT?#1LG0,WA>;QA4NSEg2<G-W2ILTcK9#\QGDNb0STFKgF)X
Q:d8XL.]::];I>cc8?fMJd=5\??C/TOC4/UI9QJ58(fB]+OP3AA9ZY-BEg1#S=L<
8[P(1#S^H&N)/,WFHZM[U1P\<E&:T00#Y50\5e\>3XWJ&5:EL<LF4PE0M&eAD.L=
]YfI,NRQ9?gQR@CQ<D;[2C(/6^..0P:U@Q3X.;RBD<^3@Z+27+)I,@Z65fKfd3G@
IQBeESXb>OORQdG=Ya@RKD?C&A(72C&CHB6Y.BBTAGYHNIRG?Q:(aT7fO??T&J8J
&5D<:U=,Z[;&L6_D(4SO)?M(7P+H,gV_JfOT4WKfQ,:>E/L;fe(XLRVAZAc+7K:d
K=TWU-E1GD#YVLg\c.>RTE6Vfg]U2:@<?UG<QVAT&Uf?/;J[CTIEIEdH]WN;68WH
d1K6XZMA9&2eHFg_ZQ>V8b_?J.Z.\K7R87WZ9[_\OC?;TZ?Ae6,ba[@.3aR]K8ZO
)+@RdTeK@QXGC4HB6.ZGQ.^Z7UX0cA?A7Pc8QPPb95I_-@G\J:ALb@-24gH0C:CA
1@c3dG./O0[TY63>?2N/EJYeSagC=fcRS1#/T420DK/OF:gaRfg1FRVCM(1bS4.+
L)DG53W;b_Z&O_Q+FaEbE]405Da=0YHFeXc,W<V;Se4JWIH3N..G:&DCB7?N2?P@
B+:)-dcMN[7UYKF)3AOFQ1;V?d@QZOCJHG8fNQI8f>JB?[)GT=9:?@e6M\68aO5P
@J6eJJG[c4:.48Jd)8#Q:7FD\852U>,#6K9G5@T=@ZL62#eUV5;NZc:U_4.,Z5R<
B#ZC4U0Xe3/>7<A#)^F:QR8VUgRcVE&,;M^8LbQ#dLA#HM]F+XP2+KYI6e)>,739
NSZ^MLFRX]))a^I]A)R[>^+O^fbQT8BO9ZfNf2HP]KSK\9ZR-=-Wg>SEHX5-OZ;L
G(eHBa4AaE/LA,12I=@BM5L:)#C_DPHgdK@,+eWOJaW63+XN3U4[V?,1c]V]7,:P
6/[ZOQV2^02A&HV<(&[L)6dDVX0^CDLFJ[a^&3[f;_Q:0d>^eTAW/;JH:B=T,PO;
RI_L<DR:a#V<,^JG8^N2TI2MG?7\EfQ.)b=0/D>^S<>dE>-9U49dX+X/0;9^7W0D
D;CP1ddSQcS&2/8e(PIN=KdFNZ80Z.b5E2[/_.R3\3gKO;3WNX^JW/\fSWKZbSS\
XCf?._fB8EC7VQRN[>K,[CJ@V?;Z\cE>GF03EEdT;H531Nc#eWg+GbREA@YTPO,6
-30=3V1B&E/P?;AH4J<+.KZ5FV]?YeeCX7;W<.SR1]cc@T4?MRfcDL+P90.4+P?_
afdEGM,@<cLF0,:;b-dMfTG_b41ZbEa)@AdcZ)1UXCdgB-Dg]X[TCbE,[Q6b49>N
:#2GV,P0-Z?GRJ2L8?_c6MY]Y-8H>TQI@TOXCH4UF.ab+XJ+DWKcM9Ae/?+XA\_C
K>,7b=-W>ObI?OeFCd/UW#I2cI1(ZCd+DAX)dGWY+5A[-<>8T(X;_#,GaO9.(SE8
2^eNYGI[7AQ,R050#BcX,8a-,9TNB9c6dA]1??@5K8I^3&<[FD]_JE8W.9RceTMV
&E:7XU53[3P+BKQTV9fd\T5TMb+3U7<0GM4T47IYd>7R=eT6Ge>g+-(:aA0](/O4
aRW30&#dL^\;E,#C8;PA;Ma944)F/Z(fV_d91.4I62P?a3dB.9AcGJ=Ua)AI)G2X
OIME:0E_G+)?C?>5c:E;[N>P?^#P2X;C8:=^EUZ1COCXf(Z@>PFb&E&WF_5Q)^J2
304]R\PXG=_^.\H&&fP\-QX(&^b9Z0=WGV9(#cg&LB-\B\3D)<[+?a+g)937<DYA
1bZUS3&4AS7YZ<\[35-JBR\b4+GF7N]U/eQR&]>UZG#L\KV#>,4,+1L,Z3TGYdHF
5A..+&P1XGK+W5\5R2B]ESW2BBA.CFL_+E/<D=3Add[G9ZSIG.6SM.\A>.]dRT/;
D__(O3>\6CJDQd4-bWUfdT<#dSNGP.]4W7ZBDO:;ECDI-WJ2123SMGe.]J.9-V@&
NP/MAA(RR]ZfYL+c-JRA2XaHU8[/bGKT7]/eN@+./R__^L6M-FHR55UZQ[TdZF8Z
>KgS1;0_H4aW7Y;c,<AJPKO4ag8/XKHN]2^PH45<<.TZR.,;\e_CWV9DAg+FLX>f
QY(7[(NS;N#W5JI.2)JfQ(@1dQB/+^N6SJ4N^:\:6VAa@=4/Q38TIN71NcW\645>
dS;_U8Z,K^d@L,e3VG]NG7aIO(<g:\Q.=1GZQX,YU&DD8-SD6)PB5fWD5f(^F9G/
9RRc\COE&6BS7\O]25641(@3G=C[MfdVgF=9SIZbZa/KSH?9ZB+8TJV9;[+DB[Eb
GLF9Y8DHM=/?6^Pg\#?:HBgTN4SV#XaHNe5.PV]7)4O+4VB.)X==4\d#cORY)+&X
ME1NDCJ>6VeAg)]:^d@I^_XDW8AB(2c=(,DLGR4RPQ7U#)KU2CC6cKf.V4b]L/^>
c+O6^F#+6SNY5g3a;gH=UO]G-\C6I@?Da=F2/=E8d=4DgKH-1.Z;Caa2=bH=AYc3
I_>(=>#J)cW]^Z(Kc?^T7-,NM@FR&A>H(.(#HR^T:;NT&@DaVT-=>YWW2E.-)<4Y
XBE)F.,/Q6\Z:4&XOTVVf/^eC/f)QVL_:8O\(-U1@affTFT/R#UeD;aOW2<,2E@P
U@@7PQN&([:4;IA-C49E:U0a2GA/Z\^dg=SWa3WL27XM[RdN)S1:+>IJG_O(7A(f
6VR=F(>DR,e=C<;&e#GUGaCOKN=P</g?&Gd/5H]Ze/XTPd9.@9(bfIWd7:@cgLUA
TcbMdT[4:;9C5OXH0644fEO/4<MS#G6W97GMc@dHAJ+45a6cK&PWBCSPO)<C#>Z/
QU9X(J&1#A2P@T@;-82c[X&2,&->J,aagSN-YGKDVTgO.3N?gE=HIN440b#6^IO-
cXPW&b?>X?I#+-J))=1SICP/]Y3V>#VG6)SHF4?[@JY6\S@DU[@1=3,-f_^NeX:#
=db.<R101FJA\:?fKC9RACSWCf3]\H#0A#Le8J@0E<[d2:0S#H/[S[H3Fc?UEAT&
.cPUZ9+M).5FRT4H1<AaIe&P)X#J)?[_)BUKQcf4OOW/T6C_GLWCUgN/&M-aSWM7
:QcXb)0<XW]bWEd1&aY&?>cTHQ=)IN5KCK]QOSB1<UK6@>e6?0F3>?0-:7E=>LM1
O2&-KH336+TNFGZJf#V-Ra&(2[?8QB.I-7Nf=:>dMF#&6cfO&=E8DdQ;06WOE=I@
M7e1KO;V1E6gR0Fd#&,T?J_0QVKK=eO.ZDCSTC263(fOGPNQ2G&=(_=fUMaMD;D-
[:a_BeTL_F5R\#&I3b#e(UHDd^a3ZW2FP944<Y2M:1SR/eY\]BZRHB=:M)23[<^W
??Y&GaA4O#&?P=#:W5,LfJNFT35?4.FXSGSDaXJ-8&,CPe+g;_G?JI\SXY=8SB35
ENaNdG,EU1U,E^cQ=c=,V59S88FQ8+4Z]LJ/VXRD1#B.V+0^2(;?8aDD:OWO-/09
JFYeJS0Z-4Y1+;cQG.#FUF6ZYg>4-ag[Udbg&+4G?=DLE4HEF^Y6898KaUR_6^B7
?N6f_T;Eg6T^A^bO7E9Q3K]d;V-E#3.VEA+<bA+@>RJN/2Wc_HMT.;\2J\(45KA.
YV3U@@5YJD>OA-[67T6T+-4LT98:Tf1>NL04G@:X3(6[FK[0QIK[Mda;5-0OeW9N
d\[M0Q)9=59FS:L;?E-BKT5dC<Le6&YFae>[,3@]+FQ#d>\f@YIB;/K4\8a+Be08
bAW[XA\L:;NPAFbJR)H7]B3PAF/1PbQ&)IV=<@;]Cgg&C].cY.9.)]+AfW,PUf:2
^E9#[7cP_:+F#0&(WSCB&5WPWKg9eAU9e2,)FJD(2G=M-<UXH)=26gA<EPG2;Q@Q
bdUU-<5N6@.<F003.EcFc<W=9[1_QfCQ/(7T(ac_@aK\TV?[dba5FX=g.Z9S:-^O
d0#FLH)eeAM;NPb]T-#JYBdMY3O@^#A64OBRe,g0Eg&=,-&J(IQO275>gP&+GIC@
V3?L[,ENS_X-2b(&d>X<c-,/7DR>I/FBbJ1(WKUKE;2aJ.-DK?EgPPO&9>_HMbbH
TVLI.Z+_K;2Q+1cdYB.17&KVKM16--c9=VC;_?LBeFSc+/=#1SPfRW7+\KT<Qd?/
^[bDD;M-<4/X=D2/\E<a^?H[U8EeRWUMKVTJe?4(OJU>FSOIP(3):^0=fgc@E?9P
B)#D,6UJfd)S?R]L/93_MBEFDR9&W)CI6XI00,E7O[&>S3,-<e88b#(](@Kg@8a<
^.K#SVPcX#Yf?#^&SCS?<JN(/=eF@ZH(>[Y:Rg<;Rd@f]#;49QWaI46CX?HS434+
TTG:U2BeP#F\H\0_HeF6Jc8;LD))gKT&eY6K]]^BN9KRc02U6@[XC.FN?NJTT+g#
+^BeJ:,&_aVS2If1#eb.]T__L,>#EJX/fXH?1OCIMfe;7#:gKEGUWfY;cBI(VM>e
a;7O[Q-=N=V>Jf1J6AI99LKbI5F1LQ+b(P>#Q)5G8O^Bd--4,]LAP83gF7W^>bdT
g]dd)Y2b\[QT<gP<T<FaGPd.+<,9SMf3P,T[@Y94[CAY?=.16>#d^JS/85;LVWC\
S8.\;3&^T.bS2]YM\^D+,B;g?YFQN79,?A8^OQZ+O<H;S>U_.O7,PEgRB_&Y--DT
B;eaWDf&_C7>+LM6).d+MTY\Wb]3?DH_?H2a2R@6N&?(]O,K@MM&8=C33MB\JIG1
J7^XX8JDLS]5+DX-RI93dLZBD34.QR:[\.F<_F@Eb.M)b^^=d>O5f7G.:DQfT[9?
_HK@gID<C^MQ@f:O/JH_L6&N2ZVa7DU?XK;)^2+e1+#Y3[/[H<>;ME(ZAJ^B:YK6
\.aWb]@gO:)dbc][KBdW9:GU?#?YC=#MYU41X[BQ+,ZSYE)U9VU-6KFT-N0C_DL@
YOFT:>67S,#I0c@=cGCLfSF41XWJ:WY[gZ^NRc(&1b#W1S(bTX)QT;[WIBMFYW>-
FH4(WaRUPI_bCIN&\]4]]\7>=PLXN:8]b,JYW;U3K\/]/LU2=4S^./)VT+#91B?S
25&6OP)#4JKJ[1K07DGAd^aSOP_=gReAM#EH?Ka?]?NdH?(@_6@3N1cX,4f(H(eK
dR49aMSAT?PB/MMVP]5\O^O]IY6@8.86\SU+)X7E-dK5<L+)-IOU=d^V#O\TbPE?
,<3+f/6-(O@+&QTQg09;1<[-bb[G0^X?3P;4^]7c)9]6-J7)>4]^HO+_Tbcd:RH4
FZR&LeK?YI^J>TBLD^Ef.FaRMJ?=0G7EBBA<\C5b?]TD36/HESA4J]A+:GG/[[./
Z@S\a<V^FEbX:gP0Ca^SMQ-ATF-DIeP5XTTdJ](@K9Z4\YfUJ@AP9_:65>S46]_X
A<4<H5HM8b^>&=\XOSGC^R];2BX:ZPc-HAEZP?bA=)A91b9TK-5[F^;U&V)DAM)5
&GAFcb2adLFDRa]e=;UNCVK\N(,054X06&71-\CfKN)0=_-fAM5?^\I-1,d@F7SC
Db]f]_dT)NBD5N03)4C\Fd.-+89:(?9,PK-+3HXC@/B.U-f;K_UTG.FW-<3/6D#6
JOG#5HUXdY-YT[1=+YH@ce+AHR#D2QB:6@VU003Bf<L3B)I&b/05L5<J2<C7d=+-
/36P=]7^RDHWd6cSX#I0E25f\L5;fM\N7/7g>ca]H_Xb^W-S/c,@Kg[RS8QMIIZD
#B).4M;YM+49T^bUBf->=QJaZYD<RP9T,cBZe./6RC8AH-)\)LV_.I)X@?KPK;6G
ZJHM8(G5Q1;4@7:7,E-S6R9&(8d^8((:&8aOMAZ+2U_Bg9DC0+VYG=.WPO;@^c4a
Y):,1K4P8@9OQa9(0HOaIWg.P6R52,7,[>&:B4P)C;&#(FZg,2H356><<G0aN0MM
C(J23F9X<L5O@B2e?ZF]5C&4Af)V2?[_W,J3QcCU8BBYI1BFC-f\IV5-<4K/4g&K
VI=F=#B@94\#A5C=5@]LY2cd:FOa=,0)T1M41S5)YZACZA-16YC6]T+\aHYGWL:6
531f[E3I02JaF-Ob::ED_\dLd3/SN[<2aJ51-E0-<H>3/EA_C7MBFZ1FIM#dYXEB
_7(R/5/>#_ZD3]<gIM[=3T+<f?T0<TO(.e/S#7H?]:R8Ze:6.^Y;,&:AFONQB0Y^
#\>Q<FD+NRT(EEZ&<?+T+QY9Pe+]We5Y4[(_gObB.?J#(]8H#5))ZJLX9cK-M;IJ
IEDg3<g^D9=cO.47G-P-]^.4[BV9<9MW4-.Z)/RP3<K@f0Sce?^6CL4I];AFd/>C
c6\3#D68-43f=W9PJQ:ZS3O,a,U8Y)PS_4a_;?I)/SeJO8AKf76J8PEXJN46XVg?
I,3A3T^Hd)BW-Kb-dAV;d.,2&>HDBD2V@,OVdLUM)0VdP7[DLDf:N3@OLfEY?MDO
3OQUJO+C[cRdH+6P4Eg0PUNPIfAM1QH1DW>[E\C2.H230<&B4Te3(RfeIJb9A,S]
YX^UT^Uc:JJ6A1=&2G)D0KA21_7f&I5H?,#J2A^W5:A+7g2TV(8deL/?5^]dDQ6b
7)PRPAXB66?X/W382@IX@IK_C4be,)/<R#LZ1edO\#S3-?AMGS>Bb37-ZEJ1@a^B
KP=/,7FD+,eP1Dfc;R/=O8LR.SKfe(g3EE:9bGaVPGMO7:8-F@+L=c)UX/F1UO72
OM(3<bJ6E6O##]0LPePKJg6LMd90f]]>H(ZY]>ZRL4299]Gc]=,ECO_eF)1G0a0M
S(eH@cB]@R&-7(eT22[W(.Pe1M[&P?3>A44XA?c@/=^0K(]-81BKR55?&Xa,,H6(
\ZHCQ1O1gQ]X,V8N.]UPc@1+97NOCd&]QF2XZbB=g94@LH])c[\d_L+;]Ma:&ES-
<3JSO8MM^:8g>5Fe?;-WIBc)=[URASUIJ\D_L881.IdV8:1^AK#F.E,62aP1+H(>
&1;8]/C>)5/H-;T\JTS+gG74?;_YaZ-RaYb;+],I^<;]Ef23;JaZC,R;,DXD8=c=
XN<KET-B5D(gD?,IKDSHTaaS?L0a-afI?ff_L\[4&V2Ge2)2DW0WffXL#A>_@EDV
&2#94A1K969EZP:O:&Sb@aFMV,9S1-,]5gY8ML(7SRD^G;(OaH<;.W&7#O]EPGAD
a72GV_VMW.g/e,gN0NEGOTcMHWM_R+1.egV=^1bCOHPg))ICM@IJ0e0;)B(?3L/0
=5G_-+G15L68LBaE#bO#6QK-643dSE:CEUg6IIeV5ES(>1HIZOS[L#,8\EPQ#J,4
YYd^.;6BMTdb.HRJ#75)VT5NBSfR416R=7B)I9.PbPdL16(>IUCAX+CfM>(/;5.N
A(\1TNWXY9H2JO)_cP;\RaD3J1Sf#H]/C=f.27.=L8V,bJ:#c/,e:+CE,7G1;\LZ
-E5d5:&6X>O6=fd7M-eK2FV)T:GW0\aWQ)M[8WOD-G5c?O<[Q#Sbaf,0Y-aA#A)=
b@VV;VJ]DIKRd4/YBTE,1F02S=5e;;egLe].DHENJ9eD?0PeGI@-Y1]=#;Nc\2U?
8MC7QSTTXH+.L>PabH[8bg_W]Y_@/:Z0.dU3Z];++1MY=EHN2C<F:6,OgKXS;^^H
AcBEgUP(bY3bKD6K-.(>=_7c>7XV_Od=B?I^]4HC@5,MXNf#(-;/:.0FU/U)QX<J
6H@&fK)Y/E_:M52=KN46d00#.M>\_cRV=E8WEFK2WY/+)3;XOU08-\ce/CGOb7T/
M/XCG6:C^a-ceN9(PKM:.eH[gHePG<fPOT^e0LE[7KOZdf4M6^d_+-K=fGSFBP+#
@67<Ya.\C^^0BBX7?AL7a6G<=M2f)26I<.@[6<MSDB#=S?F<&A3fWe>>dMACc4\1
<3C6(46TeW:R,?]1RZX&&FK-I8;;CB,Og.d)5W@J=GCVW:G[Z9+(KS--MVVOCT9N
#A;F>2NF>SdH]I<=V.XNTd5cA2^4Qe05V]B50KfSX4T>[QCDGe^3;+).GLO^94@R
Qb[<IbP8A_[ddF9+4.,(=^;V\0PZUN>,/5a<MPINTKP,&_SfcNSV6:EZg3U#F0V#
bN-<[TFBe6f>ZD)1@?/eWXQ)Yd\]->Rc5KWY&\3Hc1-#f69aR#]N31>@D2VT5LgH
HAc?+AA<K^8?XeMWb2bK5T4N<\A>9+;Y+PITIX8gQ^9gHf86AA.2-=(8T\gFL=>M
2#A1R+:SO@ZLSPK[dD7,f-fJWE<3>(-(&EfV,fbD(26gD-IcS:,bB3,T,8Z6M)KQ
43OJ=1:HLfXgf[U,Jf?<bc3G@9=H0Z,<BLgSAA&2-&_A]Qa[NTSH1LQJ80K1K/c8
U44EBcfN\ZS.=a7/#_GBbI4cB9gWTKPT@.D0OfH2KcYfJCLF8ZI,(/A6:+]DYHNB
UPGNg)aFE52aQ,[?3X#LP+c?D,.,1[M.L8ICO\_W\5@/a5=3HUd9g=4Dd4O(PTS:
.M[EQH@eY4b;E3]DGc<Z8.ILd3DfA/gd:H]DH+#[8g>@]>D1]0<D,AM&S_R_&a=-
GJ&e2R,48=6\U;6)B3[1IWg-5.Cg=F+AM.I)80BWJW)V;GV4XU6CS7dXOgDD==dY
NZ21CB):(Q.(Y;GHO@+.1XKIfbFU:?IDA)\(I=G.9N,9@@&-0801F/J(R[d+2T^&
Ea[ZTa9O1aVJLQ41gN76&9-\^,Ydg\REO5Y?ZaQ^3S2\f\#A=M>YTa\5IOS8@P-I
ggK-7\PH>//,+IMG5^S+bb=@C;2>d,IAWF:HJ7JK-IWBVZ@b-Z:f=3d&;dZ;)HQ,
Y&>U,=6AN-Y:S)WC\aF&5>fIWb^KX&QH)QaLL))OYN3.VgP8&=8H,,XEAL](Za[9
AZb)5UU/K#[8QcGcGNO.)/a<(@WYN<eDDJ37?47F@R0T?aEb2[DJ6S&N4XE[9IV?
c:&).X)/T^_3M3.U5[,R87JF);-@bK-=3FX@51Db,f(_ZKEaB4K.]-(4+b8>=OM1
YY#;RIYD@IGYVAJ/GX\M.<eM6;9;_5;)YL64)[L2deRc7_bMf&WOIHX&/3AcJ0AY
LM?GI3_5?>3],RFRZ1NK?13+MX/]C[H/O;?PZX^+F5.S@ZVUBIN?Z5WN:Z4?92M,
F[#9;6_^a,PWMNS07J5F1MCK.cN#5Ib>K]4LfX+f_X@I&Sc>240N_>OT-=10aHc:
cEQA<X(gSR3.V]-,+Ie^^]?]gD92UMA8eDI^J1>[@R8LEPY5PL,U\;4B-)1@Z5<=
\\g,BI6-9^dbK=)^1N#AB9/Yg7a0]58cJS5a:PKc+&#VCWPVUeL#YHP=54gG-6SE
1D^D[c)XJUPc4Z_NA_CbFN3E5L[0+([:b<:&,..IC][FE##R8>B/EGbGQ9?S9YY+
;\&=,P=Z,.1ZMG_^e0-M5;V._-a^3O1\G>9J2]T0:T/CYfNTCeR?AQACa[W>cUDN
F@:HL@-3JVd?4I2CM17LN6\EXQ/7]>?+VYS_a,9M1bIKV5_c2)AF-Tec:g2eCZc[
UZK,La0;@A>UU<-/>XK&SD;\4+P2C/S.3;688QO<+Cf(b(W.D&d10[[f9C?K)6-6
K9NCXIQF>M-6f412<W^g8K^:?Sd/2O8dA#DF(+K;77WSEf5eF.33/2aeQ]F&CW9@
d9>>PE9OceZ&d,H6QJc]A9;<F#\SURK=OSZA3_[BHeeQ-V,G@2D\E5?=CZg,OLCV
\G)OcH;NR\U#J0M<:;(f(MA3>=F+/&DG>U3/)=g?TVKLW]LKRYV3P5T0aBF@_eKF
<M2:^Q4JOaKQcO4=YNgS/E.[)S?>XCAa3.Fg)Zd;H\N[M@[^J(.RMZfX<&#G9;g\
a#?eBPJ)2Xc[\a5J@C=?DcU5.N<I;N#RVM)deC7P9?JM8I@V(5IB0&-d.??DR(QC
9:=X9S:7=e^.Ud3Rd>_CN\2<G,3GJSY].R0.f?^^.:JPML@5G,.A8TE)_JNJ_SH5
G7(;K]>CeXZ1VZ@gH0aAAV#>.#NZf#;8,V?;OG&[+Xf4^]\]B?T[e571cEcX1W&A
NPX5eR.5DNG5QKU2a4<9X9a?GAeLW7C0SXWL9Me<#Ke^1X998:e5bKRBAB72fd/,
U4KNF5699L=>TMG]76K<eZ8QGU9X+J6=(d3X<Jc.3Z_)82bUJb,J(&c&<GM>94X;
4KEGAJ0XONZ^EeBc<XU&b.LOe2e/WW=B=H^c(]db98=W5KY[K.[J.U0+1-\O6df)
N3964I&6&1fWCCESRUD4bGS?OGAMS57^cU;[ML^aFN5HOD2+7GIF2+U?fQ)QcK1J
AU6Rcf-APTTOERQHR-dRKCE^Z,EN->&e)7aEd)1_DY+E=;eSbK7(/38?5N=9X=0]
6RZ.51O9:+O6T=Q8NJd@IGPAP++BI)@57bM+aOaXELNfc<6B#2LCYRa#<:UPEN\P
S\U+bB()O]0JOOBZWFcA#RQW<X\EQBe;WF;bd1,bZ,a<EXe\[9_9cYaF,7b4WP:6
gYK1a87I0.D@QF2</W?Z6519T3?;\TU8\ZKB0.eI95IAaFP4O,<P=bd2eG_Qcd(f
fB1Vb&TBB016WU8((H,cP2:4R<^_OIS=X17LcTTg@R\Z6D^c-27=[KQb_Xc;HBa;
V0P(3)JD>F#<aSW:+M5<[#7VI:OD7N3PU^E4Y.D,,4[;6+<(X11T6dFI:1J,[S)H
DV(@QR][=\2REO87Y;&KFIPESF=7X,I1]_G>_37:fZ90K[gQPCO4H88CffR\J,6;
70N@.QK]K+X&KJ/6O)fB:@Z2NUG@#/[-0g-EI:@=d;b&@8e4<]ENe#=_a>.dB5O.
I28SND,<Cd057c/_DGMREQO\?ZUB.IaJ3F62@a&E(G0AB?Q(_,6c2Y8Z>4a&DOEe
ERb/U_H<(9fLD[[?BafK1MKd?Ff0@=+X+Rg)6_U<,agPOW6fDC&Jb8T&V)3+XD1]
G9Q0VTE64QfXXJMNL&V&AN^P?T0N]1.^GNDCVD#;]WX?GB;QfTPVR-?/EMSYBR;+
KI66fDbTQ)_KB4Z^FK]fCS6,G]8\K[ea2>::J)#:7PD_6Y)+G9E\WHIZ,61[+X#F
#5GWa;WfGc,Y[Y<&e\Ge=M<^OVbWf?43S4[&R-&GET6XW^d.bf/;;(OR@fc;#Zg5
Z(Y0(NQ=D+#10K.gbL(@]9cdATY]TMAK7;_I)_cQ,2VBgf&bN)aY=+/H@,I_ODB+
LJe@693ZX3Fg.ZL;8YKXT]IA^OC+)\M@N+C3>?[,KS\8<>JUX4?AW[WZ<X]8[EOV
BTPXdNZT,6VeO/5I7Xb&+.:^=VA=.G=[3SNQa]NbMdEE/3b]YOR3?<Yd7<[CIZ]1
_Nf&X3Y4Y9]5SQZ#V80TDgI0?V(URXZ5.<2b<G8bQ5.>b>S2Ic&-1?/0M5fcOd[[
_Ic-WXVOUJfaOSdd5RdO:;A\d&>-FD/,9:POg,KV/Mf7b5:E>?PY(8g>7<KV72GL
_.C.V_2@_LAIHRYT;bN@5@L03;<0T0K#](aNH2ZUENN<+PHZYQ&XKBVR_^GXa&]9
CcO55?Z65=#g?R2EFY,]M;EP/79D)E9c2#3X8e#3^dVBPg[6dCXE:S@(J4JKd&+B
(gS#4P-f;+9eNUG>_GEHf>J0gg@AaMIG)TL0S;:SIId;QbAd9Q+cf]PD.ND^U@UB
[?1=Q<A7WV&5<\/LGfN(9)ZY/3\Wc[X1D=dG1_F-0>\S&aO#I&1YLQ1EWB#NJNe+
L-e^(21+^/2./4@:._3JBV86/L>CQRN899@+MU,ReQ+-cRRYCR4E#f+:3[<][?6_
^gAJX.cH18?@?:D:_Y+W8<GG?<f[LcXY\_H(>e/@9fO9PX@d<05+KS__bb#Y3.B3
QQPJ5+DAT(?JfQG+SM?)##QN]@K^KfKS7/610HJU1=eH4WJX]6LQ#X#e7WO2(Y?\
V37U=L;)0&E^E,8b.BE&IH/ICL&Z,W@\PA4;4FQY(5cQ7D>B\:@(Z-)/6:OS02H,
CK.K_R/S0/2BPe:,g/&f)PZUW+F+5NR+)5g<+H=d)8QW.E][+WBHgBe5@I2>geg^
A&1[2_[+XK&^>@E/B()5HX,Q45376>AF4DGR4B)cPPfM.KC55/FY;7f=-,3+@S\Z
4fU\=Q04,[gF:0=I:PQBATRSCZB:Y(2L6SB&5gQMee5.2?X05F<+>D69:a;a_.-#
^H=C:5e9QSOf(<UZc0a1\PL-=c;B^TL^7GY2W+9S&C&)L-B\fc>JJQ2gFZPZOZVB
;G>1JZ>]T/>XeBO6KR]bM<dW7bP]fJaMDWga0KBEV[>IeI8OgVE[UWY.4K-=be=C
E=H:MT(EYS?PJR2=_086361XXN5aU:Sg(cO[FO/W[F0>e[Ad:gfKb-(ZAHb0eWTb
ZS5gaUE2>?85>2NTJ=<Q_aLIgT4\4EB.;S796MP/J[&Y,KC;;Z^V65Nb?\^:VPb-
+CY57[1/1aEb+aL;@:A[]OB>g]#b861-QW&SB^5=.,8&HNBdBeba1V6Ob92X?e0)
\^,H>0P\@9e^^:#B@4T@?QG;0YVB>A5KVGC)HZM@9Z<G=fQOT7PVGB[1Q_IWLCRS
MfIT1d8#F<D0@f,GC3NBC/1=PECU?,8E5>N97Oe8EA;B2@(SdQa5J6>/@Q8.[SJ<
^<]_SVL1W_9EfTPEL;<,XRIeg=D^C88cZ#D3<,SD(>14XY&0C9><E=2>800bX(E9
,5c:3)M<MEN06Mf>_]HKd,XdSK7N9W^R-<G#;@:?OF1g\15T160V9A.-#L?0^T]K
@fGZZTN6eFJe[^_B/H@\6bKDUJDXUaBISN5T+(FKKed1Y&YND7A8W#Ma9AdZ5TZ-
#86#1);)/,Z2b0EJgDAI^9D<2gB0IQ.;d20JYXLFQH_.#XZHH/U)]#J37&ce(+Kd
I+@5B.8Q:CM\gTP-d1+Fc]c=BVPWXDBB+Zag^R_8)9Y)A\V&g(JFC(FcR6K1U8HI
46?W8+4I<=70MW]TMe_0BI2][MC.SAHS^34<<ZM1YRK\d6;S)DS^DK<>M/MDZfC1
E^L:<372aQRWgS#+(Z@gA_C]3/HU@_U<WIaZY4DaC?.,ZG@&_O(&&:X.7RFIS3=^
a#32cHS/+IL6WEWe(<ZAb>1WAZ83Ha&I/Wg8.N/0^/HQ[<bD-A2YJETT,)I9:2YO
g^?N2c+Y1SM3CP?[1)ag=<K.E>=(,[Q)-HV?>V;R],]O7=.8[5EcTV9GJQ.]_L])
IEea,L:DH_B@cO1+2g;8S)I</+S7L73dWL:=]B5LM\S7<96<3Kd0HM(]1ZMVX-g2
7#>]J(]f((LBI6J_9]5XJWA2<9F/\A>Y]4)U3[\KW[4&E_]0AY7RKX@]@?Ee)(]?
ASFd^6R+N6g0;@AeW>&MUOT:(H?&YE.,BbQ2);0Q8H3\d4E]L43&9[_E_Of?4QWa
4;W3(=L?Fd#]eO&8(^-a^eRP2<=57OJAMAZ5#>IWHLIBK=bSGKNgB&6+KKb5_>Y\
V)bZ=ba>QJgc_Yd/2MJ[]c7,6Q,dG1>@+M?X+d3L8Z:AaXJ+PAKYSBS[<Mg0:Af0
[.GEPI_81f>b4OcS;/PNEHM.E@O(N7_.XAXD.?FJ\6[H_XC^:D^3JGB>AM[?CcO7
69JSDY_>\9B^=.@-@=Lee6J(\STUS-1FM)63]R)972846b^0:b724ARE2_.@>/MV
E@]H9[&XC6T:U.[C+IL8=(7/^85F?3ZMPabC7Z[#.NFTRO7NNeE7>:\Pg]cC0gMI
+)c-PV2_W#c9fRb\+V,K/P_:U=bZDER#DVQGUKf(5[DYXM6e/)7b7TSMF,#=cDLC
#De9>4cS=+EBGDDH?>c(<GOWfHe@VM:I/X_TW4=IF)_;(S.MHBHZf?eV-=cTH7\@
EOV/7fEE/OFQdT_Pa=X\TP8Zc7XJ6d9C\OHdKN+V6c@0)E]dQ#ED3/)&-3<JH;=F
1/WI6g.VKE9_Q<LOI3_,>F.8<<AV^NRa2F-fO5IEI(]4:f)fU[IR2ee5S\6.1Yg/
0DeMHJ49NaEbKQ2)XIdI^[VA8LV3>5;L#RXL=3SF5?CK-9;(?^dcLT+/SO=[Ub4H
2TBT43,bB5O>?#M\(T+8U2V59=TQ2X?SZ\fW6#<_6?D;8M(^E;WQ[5Pg#<KC:CNQ
2/D1S0MT>9X[X@I0Bb0UPJQfUI&J19UC6O#D3F+;W[2ZNV_ESSLd2D(].-OQMIT3
e0JH^H7HdFOBFYKF.=6]9#Q&0F;EO8b@KG(Q\Q^/8gK_U3?4&[SFd72:Sg/a]B/P
H>1fN),-R_EQ3Cc_3<AYTB\g;R]gB@>cCMBG[M-0P5XF/,=()1OG-M8]NL1#1B.3
)NW+gA2<JSG/#]FD@TKf80Ld4=R+I)Z66Y=(>NcY^dLWQC5^>8Z02<&K?7BYfb\)
9,]8]C(fGP&&4/8XD]XfF&/N]Q)/BF=@<fE/MO4/SE7F[B=-Y/dAfE2N&FdYTIP-
R1#(>^#<>]4U_8geY:[Z[H@2--D10b2FA(2Q-=F=MG0LP[=7Z1A7f(;T2A^K\bMQ
a1]C5-RO<@[K)O(1.@4e]g30-_@?c>Y22,aMF&e5;E=WLZb9M)_W^4L#6ddC@FE\
G3-/+?9/a@G6ADbC.f9[G2f^U^WY3\=Z]1Vg^9-,M56Z#&=IdXg[MTFcaVYKdJ]K
KaAE09RcJ[5bF6UZS#9Z#cWGEZ86gYc0PK.\^K]4I],O6O+=(W2NSVV)2NP2GSd(
T#J5JH;@W:G9IIT:I?@Y-^:_7\=Jg\gEEY]-_[1_>Z[B]QE641TV;16@L3XOGDTd
NWb4@R?XLF#A28F;3,)P,_UAF;]N:<RMCF5ABU/Ae]eNREG)A9ZWXa2=V[ScQ<bZ
Da.5PHa[(1c&,_N[[J;>,:_)9==J+01V:P\91bGXKbX;VIb]?EJc(&U6TX,_5)&+
,7)09\BR5C#]0,TZJH@:g[.J#3M#>_GNBFBS?4T2;&8+KG1.E?fa7(aPOcE:\<JD
F978g(/#@]C7f7MMfZ5[e&RR@L?K,SMJ)2AMR8/C]O(YPHN21;I0Q0Y?]D9IMBGH
VfB_fI:,K6La@9,#Ld4J;]DCUI1Y9D30O=[2HOG@=TL#>&&W,@7\P.3/Qf+a@3X-
^BfcZ]_XCHB;7PW,17:K1&0b:]XG_,e3E-4M@0\[dF3OVR.ZDE)<d<+/A9]KM=2E
)H#K,6^fFg.RX.HQ?(5(_W7I(W[5RPaL.CPb5e)6W,7LWJ+M\I?=efI82D-5SYN3
MRaKHG64,Fc(MTSb[_db]+J5CF)da48;VU7L+[\&fO0D0fX^U#Ec]7+@B#PFD0K^
S/\^>Q8J5,eI;&3Lb64(J.Aef-3;<8bQ5dBQR:X3?V<g94RP77TBc45Z6?JYQ(J7
.>_6;.Z01G#T.5R7CK&,^R>VK9,L4-8c0a;MdINMUZF/]/d0KRUO.4U<Zf&SM(_Q
e:G^XM,@PD#0A@9WC:];[H:fd6Z[TBY:P6_HRG>6OHJ\M0)LQM2)WLR/>AgUPH3Z
2AM-1^3N>B6WLcbSC6=HSQWV(Jb]9M.-ZTQPQ0F)N/)DfDVUXYeD9Rb/4KDCU371
4WcXf6()Q)IXNR?VB4+CH^65)6Sg/5VOZ@?@()#X??gQC&T.NId+-P78YbJRP_PE
JEXXf(JN8L#0M(&5(6/4b&_4LVRO8_gSf;d8C[.(D&LBS@UR@[LXD7U[OTPcL+B4
AQ.bCdb;W#V@45C@&,Vf7U)_L0d+80MJ;aD=#=/W9TX,Q/c5,E9(&PH+&)..P[_)
0NE<&0&::XP0,a5)f7,B;J+M9,KU3ZY-3,1d_?@PF4C;0<223Z,Mf_Xc+L9VeFSG
]KY7+aKCL7QBD;.0JgHMAD6E&^#g_B/bF[R]G=#Y0P<Y(MH_N14;RIH8b&==LFQU
ZgN6NZEO:72.7E6Xea-PPfJe_3<UES9.Y9&936P/(>GCQR@b6Q3<4NfP^T.e+MA;
0dG60aB?8E-5[cG\c<ZJ.;)6.HW?C(Bg>W+6LJRNSfUFbZ<@XB?QSQZGIG>.Ib&I
aZ,?YaH_G>fE9Y=.8O6T7g[@@b&MGQ&M@O[Z-bJCG-KHFa-Q5a7M81X_?.8^44aO
4.CV22fWd]69Sc2&OOf0)Ga>^d1YE^/#T>V>#<]+X#6[-,ZEVeXH7TEJ1Zc36NI;
cLIUI#T1FHbeYRU+K;D@,-V:fIBeITK,e9=MTZ&1C9VTbGFOH:\6c,QYZ73.@43/
J.H&F7]V;OY_44UT>CFDG\5Nc_.:Q1CCFca#2?P);L56@G=9Q^A3DR>D(_bBV,c0
G6L5BgGgHc\3a=[I_Fc\,5\b?4KC7;9gJ#4NJA@&7C609,P,QQTEN[\T-S4,2(4?
dOJ+c8=LbT5d-YRV&>]a+QD@1Bb97<_?5a>)M4G3/21[8;VA#6P8YUVSZVJd]U3Q
BM.,L=#U.OJUFAW6^9[LeeMD^2?>K8564g2JBbJD6ObC6bMHc)][L\eTUL@NLf07
eHJ2W5XD>@g31_3:JQeeB?J4gWC7)gPPYKXT8?Gf]^C[<JXD^D9IK4ea:A=)b:CG
HP.ZGeKab)=Qe]T,,(eT5YOG[923XQ]CEdJ-O6cJ_XCM,Ca7T:VJO0F35Q@<B=B>
b4,[[N<P5RaO/]I4828+4WX5XU8EMXQD1T;Y[^OP6:3##S,#UZY1:#=+E3:ETdW(
D+AF?4\B1/1,C\/b)DLANROPWG[XD8GIMOKB@@R:G@g<IRP8.@3/Lgf,?,-WLcH:
W9PY=E?43aPJ2QX;&CK\bIPN=:T8O9=L<XS+,P75M+P>86)1EgRc<44G\U8.(Z+Q
(R07&#4W7:>,F]AdU(50[[-JE_3Me2#;F>GAHI@EK&f[H\cQIVe)f+c+&ZS0e>Ve
P/7SC#K2KZgN?9/\6\ff8D(PA^04e44Z3Se@/[Y,AU&Y+;Pc3[RdS+##@2Mc^F)Q
82R4c7-1\a(>>gPYVb7NAZ>N9^NSB:C<KPL.E_M<TCaHT9d4Z>9PC8#9eDgK]G]O
(Fd]60;ZCg(;dNMV(R,^WXQ22dT4&GO32[Z9\J@KS9W),c<O\QHg2/5S9LSA99_=
P&.K6-.^]:9Y&bJZ\Q)b&:]SN(F,S=@DL5C>2&8N<XXGYWH6@G2YA]3.=A(=9RKM
<;(\HYERP=86?I\G>-O?#9WUbMgE<<O+Y8,04[W;3DWUd6FPQBDUO.V,M1HLVJ+7
c6MV2XR5c+Y4;8]TGBLFGVgH9GT=OWQg6]S8#7,F5agJN/gG_+gP9PD\cBZ[Y6GG
R8fC]6-Q\g8#+5YLN^2-f8#>TQ1)c)bE]+aE3I8^@1eZg=9<=3WR7D1H(B7:/Tb)
:5SgD:P)T9-&F[ERSV]f)D+?c=-NFEMM);O?&?M,cC;8LM,20U.?;5;U9XCI@>?B
;KGP17RLU7g2>L0f<)UNWf4b@(=FbU6)KF^e3[F0[PcM281I9]8fR?e+LRYDgK<G
,O7GP\?JO=_>?D8_HBa&(fR\fMBg@N[\aAMU+aCE3K2&C+RI^=Z1?+46#4@?C8.]
#[/M6A8g]:OX=?HE9dO+PU8>Z0Q(NA\g\.UK+.W3X+;[T/fcZS5Z>;c)>1MIeH/4
C@8d\QC-IO+#1,[)/0J(3-?K46W]&;#cHC7Ub(S]K+@O029;C=&/e@-?PgEEA9fP
DB0dO;#SN47^?LZ/e>MH1OKK_ZgS-M>15+4?O8[.=P^KP\J?<?SA[TBRb,@T,V=N
W<EbZV?@TY\G4_T(E\:&@&7=79)NVd;R.;BN@^/6MfC0JA,.#\N0dMg&fZ5F>gN+
-e@GS<a,\R91d?PK&6\>]BO8dR=N68CUGAI=7U5XA3P(WRRVR]))Vf269gcH@P#H
+f-\Y7R.C:F:HO95OV[TQ0I)2(dNY7#Ceddg7N\TdQR4dD:YB.M2W\@EO[YA5W)<
LSg=gMLKLH;62eFD)50YF_C,dIPE9X[DA8f3I2DKcP4S?Y2QO-RUX[<.W?(+VJ6)
D\@_-=X?MFdcA_LY;0^6VLYEGLaF_H^\5S>=58CY53c3(BOaU77?5-0bF&M4[]dU
a)[cNR.W,LV=_@4;RGW;c;&b2:D3W=ONNOPb>Lf0RRA4JH6T)=Y^eG08V#Oe-(SJ
1,1]_0]4HGC1(cK,P)bD+9<5:T3)F,eBAL/U\<=:NFR48:-f&G]NPM:-NL?5.M=\
-:66;28TVdAL4D<#KO0DK60:2#VS2+^)S^9I:_D[=C,\X(/IE[<6Hb1ad(5JeNdZ
UZI#:P2>4K71TE6[W>(\N)f(U<g+A>#.+XQe4ETKaIGL?FNPN(0EeE+EdHPVBgJT
MCXa9;7TbdR7H,5LMPGC75J3XW1HZcC&,@HWe)c6QJ\<>-GR/&]7[?R1U6YA7P>e
d^49(RS-^aUP9aOaSEN]9<\)E4Sgb9;N9@&dO+a,.-)NP62#.:\YVc[XaL_a9;Q]
+&Zd1TeCTUeE[<BJ.\-bM/3((W84E=YNKRDZB:&\Z)98W-Z:,-69M9cPPGE9Ub@d
1a6JPA?33dCJ,X(=0LVY6+\d(@9gd+Y)Y?M,W<7SL-4QZW03V<IZX]a49a[.g4_5
gR@JAGJ9\/1X7PXZ[H<4EQ,RR4073-e_dH0VZXdD-eC/6?+NDO-,=A#I=4/R;J@@
gOf,R#-UU>S1+50F-=240.+WD1baVV6JE-#BP)dBJ+cJ3SG5LE#.T[:KMN?6gXL.
e9gNP)7?1-6Q@B?\+Dd47^E[Hd?6=VD?Ee&3XA#PgS//>#VVPF02Bc>F\7fKGG;N
<I)9RP\-SS7de[CS_>Sg]#1<VaX5efVQfPaZP.&/^2Vba_b/Z:-/Afc-GOOOO)[[
B9d>,U,#.b6M2._FaO7f<+M()&ITR1,,8PfOD7RL\cE-K00D<O@NJ:ad:DA/eSB5
7GTEf[&<=:12Q/DT,cAFL.U2)H_MSE=&g@9?Z@6O)+\2.+-N@QVJSBN/^SODCYHd
Qd9-/?S0Nb)KeKEA]NeM4>/[&QV(gU]6TYPg+NX=#BTJ8&SQc/8[fGd4&&\F=M/K
7Z<c]RSO<<7#d#3EA3NX/W=9BVeC,X,:bX3OeZ:X_BDBa:a]aV,>bYcMP1gYWG>C
&V)FeZ81\-Z9[1#fQ]]Fa.QEX9Oe=O\dK(J=\5FBKAW\F)^J8g(D^8g+dC0LR]49
UG7c483e\-9TFS@EFa71KK+1^7#E&Y[P^J?S]g(9@I]B?P-J^1OOgE98d0.:gY1,
-?.a)7(D0).,<0&5)(^OZVO7#\?C;T.H=WV4K7K?e7_P\1M=Z7dQ^2;I_Ha[>gJ)
WKfa:\Pe(>P(BFCYeB3P],XBTPHP+6N5f0)B]&F;\9O:cJ?5^(fU2>R]4(U6I?+)
5+KX1PCB77#K2Z+D.>T<Vc0fHY]FJV#(#/.=1NfOXg.2R>W>V#?AJ20gg]eC#gO8
03FcG;2;ROZaN_#EXN1g/&dELc_:29Va=UG9U>K>)[/Oe3g5R^P&6VT)4,.\.Qa#
EB25.55[T5NMJ,eP-(SBbB5>5;:OXeU9@g;3_8K=R?b07Q1XYc>OK;^(E-W61+@X
41^T]1TWa=-GRQ]=]5f>8d3565=4&2JN2X(:=-52NP:I5SI,fH.c6@3/+6[5.cZ\
fgZ68Z0a6&2Y+&AO?G@)-KV\.(R(4FdW?HLGQNW@[aZOSKV,3:N<EFC?@f^]\9)F
QUY=@CfCF4MA=UW^LLEQ[.&DfFNWa&,YbaJ9>YZUYcVF^bCZ^)G(TK^,/,J/c+<;
7aK>Y.)2&ScX9#<GgdK+.C>/=_X,dP-&HRgJQg16)fV44Sf-b/WMK2Z9O:+8IRBV
C=KNfVW+1/W.Q:F5T?fO]Vf_G^LO1[PB=9\=N7]D):Q@(ZbN2gQgYQ[[]RK@:W5;
b@\HD.EJ_+M/FQ(QHKM2,U2>M24=Lb66VVAAT([Z0LC<ILUTW.GL,\1/6/>G(NG=
5\<@XIYa3.OM>;XOeR;4UaAFIMK1MeO27G2a:D\0HOSd_DL&5749<F#(c&AXNY]R
7VPd9J6#R\^2_Y5_TB2<E;SR5+Q#Wa3dKS_#]ZYaK_Z3Zg<Yc^b\g+^Y\E9b5PK6
I6Wf9>B[-\VRM8BY-&4DZFS;f5S)ATg>R7]=PQU0VF;VM)M^2V;E-1@d&O6)<;=Y
JP=SIQ>;MIQNcU3B>7=^2R,AA[.,Dg3_/NgfGZ@@^e2HC&#D3;,X6aYZB(/AX-0R
bGXLc2Q8NEE[f2<54ed:XP8ZQ6K\>MF0>P3,>Y,\I98(A+I#BAR@=>KK>F?WYV8]
CXbNDb4IDe@#Yc72#8LPVa>B5cP6P5d^9KZGCJPdc,[&\;cOK()b^,-U6YWA?7,&
^Z#7S]BK;g<JFeQX:PN.,5;TW+O3SVOGdXU3^UQU[]IfQ8^;R:gU[8FNJ3(R;f9Z
X7JR8f:QIG1^]a055:Ze5#AAF>IedcAeM2=LE,3+H+Ib>68\-bOW2.=ZD.+1Q@4b
f;fSJ?JNCI:H-#\GABT+.Cg;4e]KOIKOZ?bF4L6#D7^X#?46OG?b+U>A:3\S+a0&
Re599=YP\<Q#LLDO/E5@I:B5d6P->Z1a7@A]FUbL>61.LMVaOE[HG4^U-VFVS@bQ
3c-^>BRE:ID\/aTILcMfbH;ab/(3,gHeV^FGATQH\SQc[T3KW.X/)#54_C8?_26c
DdC:9gE.;&=250:S881&PB3OPD_f2](f:86[):a(acP(#f7)^^(,Rda4<PA,a<=J
90CT-?f\VS.6Y-JA05[54^fEP(-5R3LOC_T^KL5TQ)UQ[&X]fEQ(K5Y5K9PTLFQ-
A7cI87DP)WH1>6D0GTJTe=ef)_b983cPJ(#E15VgTMK7fI;,bF/Q3P@=UFfWTQW]
Z#bgANBSb?F-b4eD.6Yd.I&[BUN]]:SXN#MQ78Y1@:93KNF3WQ<Y\_ZYg<?2@VH0
f>X#RN6f4Z#S(T?.DKdT:97^^EAV?5MLF[[d(LG+?V-SPB,-gTaE#L65..fU]_B?
Kb3?U#L>O<.RC.)F-+8LY@O/eJ/=)ZLbIdUaW(C>R)4M^],G25>R7;D4&;(Q;dZ,
D_>FT<L@&-A<7BO8)DGDXZ5BB-&8#J9<FA@S;OP6DF.U84T?@(Vg>gX0DDP(HVTK
RfQ_QM85XH:1T,c#6663TB(W-gU\CMgT[^:E1cX\USM]/3@XQ(RM;[/eQSA@UK,T
TO^U83&\\cG]@dJ,XPHS6(6A823;GG0:\UE2ZIK^\UPb<+1OUNWSARBMfMBO+9@L
^dCL(#DK#P5M5aMVPAIR5_>/Y.g(a]AZf+#^7EbHcgW=3Q[JC2XA<c.HgT]9,TCA
@Lbgf3d[^d:XSd/,E.A).Wc9?P7KF.>@J-.NG9G^7S<)\,U3GYc^XPQ))cHPOb&7
@2,_/D.:>X?gcg;X&9gcT<gH-dX64QW9/YFAZ32H\GQbZ?0Ha9@Sg]_QdWOM3&-)
fbRGg#@>1QWSMU,#28&,AL;?dDF7aZ+(bYEa]#0g8N=2M^afS8([3OaV48COGV/V
\/<1=8M9S?7/b[Jd^B;g_^B6f-Eg4TdV[c5EFXYR?1XeIfZL?e_gT(/JLFUH0;78
4:6MY8H+@7ME=ScaL9(:Z9AL:)RBT/@\KRe@Eg(=-EH/2Wa^?ffX:ca7,4GNTMGL
5CF:+GSVG2FM331^FUY7#_WU,BeMI=4]CP;I4YH:_JNRFR>\-A/FED7]1?,+I)ZA
_)1^@_3]905S8;J\ZQOF;g21]&8,Qe5G(?+WNFB38edV)Rb320#=IP@4IY[)EZZa
M5/74BZR<fgI\HTN6)#DL/U.49:WN+>7XL(CX7^>;PIAa5#M5;LIIN[/HRULPgQ.
W4&P1#FG/JOcJ^P0?1bLO[4=D-RTA:8[&T8gdO:]G-3T7E91R+8BXWK@BE5TJH-/
LV;T/aEcb]fZ+QT+HWK=U]UZ+fB>L\H[+1L^]LWW:YJ<Pgf/CF,R;L@V-fHLORUO
)-g^\c(2\U\g0AV>LP7/Y.=F[@O,,B&ZO[VIWIb><bBc?,UUPe0=?S#4:SfB#e;c
BW0E:0B;a8-<,AX7T+X2UHSW7>_H@CVI.3bfX&](Z1=Z[=G+@OX?a;SAS?3TJ,Vb
9@)SS+PEE0dVI8<fg\O3+<Z#e/1\AOG>W>2BRg=FCRb2HYP9L>D0AL&:D5:8\D^S
;MS[#G3?KF4_DAU8ZI37ES?#8N+D@eC:;:4DM.-?TZ(N.EXOFb5e0QM_J0.063]]
]#<./e:,YHcH)1[F-G28U4cT\?a2;KQGR<K=8T.[ULCSG@R[7@)30X:?3G,&N#/(
e)c.P&IZ:X]Q34C@/;(+6.N>gM2DI[6BSF</@dVDL[(E[(ZDY\@4,#=7gXe6KR>6
DVEbc,5E0de_=[e^&BB.J[R^7UTL)FdX][a88EcF]S>fG]g.aGI4.7DW4CB2KGKE
4THIcCZ3J[,JaYGJ(IM0E1=[Se[EGV;1WB<<2OX\L+#)X&fH7.)P:5W.R5:Y@PEG
&G868,^bMXd=)GQ_HggL/M3PO13g4T@5^UIE[3_&&W2M&#MG6YU@_[;)Y^A<G^eY
/AAXIN;A_\=+.+_<&153?+#]:@O@d??-):>ZWJ]/bYgK&D)(&<JR9&_S&+-FF<Ud
d+,KNK+dFZL][I^g-ES<CcT-+d=G@N\1GKgF_aQ;1f\^&8@^Wf((5OD?>W_#b)Q_
fQG2X7:3T/K6VO4d3[Y_e=0KJ/GCe.fAF6+M5ZA.22N1c.O4>C:T_K)C@\J5G15@
V6WK#<LDa)FNEEUS>b:]1WFbJ3V9V,E5]GU8IV;.?,PRUA@DA9^VFabR)H]BKP+5
:Cb6.R:AT+0:fB[I#3c&<:-B^MbQ?4L0+c98[FT@N_0-H\O7[4fCH[OM:D9U/WY^
>2E1BJ,1&[ebH>B,7b:IJ]-+N<[f16G7dVY6bY7g^RgZM.27_TY:SgWQ:Sce()_X
XR2MS:4GT>^KI>gYU6MdK5P8+QBZad>T;\V:;2e+>,;)Eb1#b(VF^LA18\H&5a1Y
Q:[2dD8YS:c\-&(]DUOPX].]ZPC/fM)bH7.?^.Y7L:LT6W\1,&0G&b&HKEgD]6f(
9K&NV3@TdE^1EJ04B7M.;X&HAGc#L,KY#H]J=JDW&S##H?0ALY2K<T?[=N6a7SBL
>G_\GdWC8.a:D0(>>X_3\8ATKM+@=AME_]eQ-D9UcSUJ[-7Y6.HMTT=O:E6_#Xbf
WFQ];&?ARZa;V6Q5e3PBHOAbHY6TNA8c,Y2c\dR(E81-aE\OTYEc/KM1Y&Xg;M-B
7cgc]+Hcd<O;K;[K?#FJC4WM;-Fa]24M,N?c1<^]&0NbdP<PbU7:D7FR7F.N2+N_
L3BJS:PLL><:<QXKFTb4?_:bE^f3bM.bZ@?HC6M^G4,=\2fC+QDDfJ3MeQ:7@)EM
>#Z(]RXc7+82,-[C?6<_C.BeO#@K,ZBP0E7?#AQ[SRIe\W\K&AJ+AAI&dG23EH>9
^SSQBX<>6PS^c2fM5H-A<N@H7JY.9.Q9g+cK_E^7Be94JNO>=GSRc(PWQQ&Kg<fJ
\5Q1NBYgZfG^Ia.2ad1]eU<N(.bR?(?S[@T@aMEP51&.QCZe<Y]BMH.NB2H\b]9N
:XM3fZK>ZS;Bgf#;+WGELZ)UCd7/+[290N7Q.T/<-bKPJ]L0D&:0F217^TS_8EIC
TB[<eMbPJF2(7fHBEb=S5<f7G^b2#U2MQZP&FPXP:Ca2K[H.Ig=R0X00X/F;FI4=
Ce@Q&C63g]c-ae=1LPWJAgTeE\XU],[e2&W_^XeP]@_#.9ZVGMWC]C,8&&Ped,F2
(XVDRYC^HBMY&W690_@4W6VWdL8XeRTK1IBfW@O;ceCb6(?X?;5XNSfYSa(>I\gN
5_;(<889BMX;T+-Ae]9G_-Z5P4>6GfAS.QDa-:@/5WC:a2ST9Be)Y?PbWSO+FFA(
:[-+TSAF89\f.:F#aJ;O??S)/VTNWV\S0E&g[D0Gdc435a3,&TCfQb=?@)0W5@<g
0\+@S20_;GG#W>K4+RQ1IE.+,9I])?GgDT;W-J9PSFDZ60eI<E^5<C1-]9SP#/&M
BJ2..D-M::e91<L)TPgAIfRW+WMX>Ze#_14AOY,/T?X]=&<VH8O.R&MX+1Oab1e[
,]6NNI;2PW^OCM+)+5dO@MA,bT\(#8Hc;B59OT^VI#/\b65cY:>4IXTW<ME;AfHS
;.G<HJ.O[W=YfT>PE5@MT@N+Z-Q)&6I2&&J0),:1>W_DW,=M:QCeEfT;LE9)J_QK
MFN&3HS8daFcF0@B8/gS([G:C]9E@(3<2\fT5X_B=g#E?F=K/QNB(+_(LO?C[=:g
9-[RL:b6:)HXbJ-PRJV?1MJMfE)E(U;e09\)>Q<I:##8BVaf&:E)[L5O1H3+MTQR
Q7Z7=B.P,F4C[[g@,eQVPH4IS0KXO7eBaYZQ.eJB87ILGb]Y>bJ\P2_1;-_)034)
14=[LegJc?[?9=a4DKVK1.S&][<B6eE)/>1B\1FR0=M)OY3;d?UD^)_g=-TgUCYg
&7Mb@QWPKf>4K,1BbAUL;\0B(fM:D]3^<75<WXWBaX[T9.Q.XX0E^8W0H\1UZ1Db
\OcIR+RMf<E&<YB8?^;R2TYG@a\UG(Y/G4+d@X.2^--/3R-6D81.57Q5\LDT:)Vg
9C(J^&6CQ8U&Y7HI[&RDH7LaV(QQ+NY_+7H^LfE2847Q;KIHQ>DNDI9FX8Nf_B/?
R8<F@f8eG+bABZ&(1/]d-CU32Lg>]]/g:<_Z<Vb\3b8-WYUVU2U=UP8S,TN(,Z:\
:-a@eA:ee[TGXf7<SP7K)1gG/(I(8RO,4OGW>g;&fUDV>V4Q=ARc6S)KN8)A^Ab/
2EVN]+]a)JG81;8>FR/,U]8YV(YEUH^FcVQ^9F)FfMA:WOgJ#C2G9\AJO?TFYJEQ
41.-_]&KYfN_d+O7)6]Q-8<Pb[If^3__Sa?B^\;^JC2Zg_E)XGe.fZ@+N2UNDCE)
=.ILA\5&bN2.PRBH3cYO3H-ZgX9[MDPT<9FLYNFRSDE=WNeSgR2AfZQc^\3MH]7M
6]-W])KXY82C.X8cFF<1PbbBS<V3>JAC<H0N#d5cS;WKOeRKO<L4D5SVE8aX1[c7
@9Z_4TIOLA1&bDV()/^0;(f2V4T46fAQ?b]G7_+H;AcR21QB2cI-/9Z>R+1D#W<F
<=#C.6NP2)fD8K8Z:bB\X))<26^;85R/[Q(#<UfTA?@I7[=;H63@[dMOVX[;DDP3
6Kg]Ua/QY(EVTXR?U(^_9?97.<LWcH9?OJ]IOeAB]I=3_J/=+0[bV(NefGb<<@.Z
E2\7Q3Cc8&-/NH,6?KP-77K7]T<HM[8/O4@-78>2,JIGQM<:]LRCTR:&:b_3adWc
<\KPg=8H<UCZ2][@63-IDV&I;MP<ECe8O[^A9EQ3:Z@K>ABOOYdY]Z6)ZVA@]&>Q
W3UM\I#>b^C]f\SRA.84F@M^@](_S<5H\@89H<=F\]bgKe^+&D@<J[:G,2^:fR@&
8JXW,VF>=NRf)Q63(2Mf-==@6-;(F-cC=GW.X;\J_@c2JQ<4U&0]Y]8ZfdHLgZ0X
WBA?[8:b9=B#e5dg4\+8X[@U/^E5]U#dd?(gF0[CN6EeU::R,EXXgEPeY8R1/Q0N
]C0.Iec#IV2G]UT^WfV2MfY2=2.+//<DQ9134M@Ba0POK&;8e0dTffC:I,XBWCN?
E&6;>?1f&5a6T3[]YVVWK2Y)+^THaVGf=.<4-O)YaZ.Vg2\);,#WcWXcfN:#))QI
J0NN,]H1/VSegPJWfIW+&^,?VTUMF[@,RJ0.-LY;K<H6D,DXMaW<\ZcRQJ?P@O4;
aC[[dA2HDR_:?Igb4Bc2SQVPL=6S9.+.)4X?7f3S&;-^X3cM,Yad7[19>H>6YM9)
:dc/S9OQ3XE2a>FEY8);K#SfMMW=VT_Y)-6KW5E[./.cJ:\P4U#2Y+&f?6W,UYfS
3Id64D5+DKYC]#CfAKe(=D1B@J3R/UBV\0K,CX;395/CT?):#J)P>F;W&>X-0a?H
)DHADKS?[D3WcO\/8V_N(D4.@T[I4[DCXYNbGb9@3UJPX)],6e6R(8?;S3fFggGD
\KRXIU8EK8C(I[(>a^,=6N;g>&[8JZ2Q=L&\JQ9f?F9(0MM,CV+aJ;40DTDZfW)D
[Z7T>\\1PaR.<W4Fd_4<\9Ac)bPM>JVU;P:@ZZM1]VV[g0G0>F^5Ab?^:,?ZgKOV
D1HJ#WUWIM(:<3QH<O)d^AfECUCP&)2DJV<&8@VReM:BX;fP/O[LbB71D06KFO.O
W:5+3:88I?<[IKc<\HaRF&g\g=B<NbMQ[,A+).?Bb7X4@[#gT8_4-4bMNUOG\)Ya
).]gXFHR[J[GLc>;AEJ.JJ=)#).;=_F0c5#ggZB.<48TgT4@D;TR4]2NH)QX4]bG
NAFeO56.J]@_/Y.KGb2B50:Qc/?\/)DbA7<.Y:?18]>[/KHbMGbRcZG[:+bGK(N3
K\AIFL,eYBAI,(Y/3EV#SYcaD(CZCW3&FW^L+;f#2U<cG_&:O2bP(E6<4=[.GD\E
VGfPA_9I,g22[-5]Y@^#<L:P7B1\dP,GKHL3bV.O\WBXD=<Q_1_bd]Ve>UE2MX65
^Y;(e520Ag#5M)IBZV?dc9A<D61@)4Yb7bFa8C.#BI\LV[e5_2cZ<^@53c:^fYO:
?ZMI#=e@8RD(DT2/G:a4:&LPKgH^]6I\SD;3#KW>&?VXMZ71A/FX&^=S?ET(0(/<
a0O;:5W4DM<Tcb[KFM722;8&bKY,?:KY0ZQJ?(f8Kb_7Obg=_aRN-@B80;P+d:T[
ReWLB,CeeZ3-M;XcR81@#)-/8?,:/^^>TM4ZZC,cc@TBfOK+8_<.10b/@4cRcS?4
7ANR&U?X)5DcQ:eAN&Ldg.SJ0U)FZCcY@@6K579X2bc@SQ:OY+&V;^>OA::16BCa
[(F5Gc?GQHFQ<9eA6(9g840LMH17.RVXQYd\76K-OU2XF,:U@@&Y,AICCRP4J]0#
0JU&R(GDB)XPa3^PB6,L_EY:C^K9d?71-LP.YD)TJGf8=H6<ZIL:3ES(DHF]+B0O
T+:[5/IFLRCbX2e,5KRJ#:Y07;e,a#5+6dCc.MR1M?_(?LYDLEE(=52W#(a^_ea\
cFT&RR+\O=7=H:UBE@Bd#P;_I/?47?g3I4HLQ:]N]e[;c=U9IR8F?4^=_VU+O&MS
Rd2/W_JJcT1&6)#?7LE7;L,<S8cRbV3Sb/&T,5M,;Y1N?ZC5(Y0ZYV6WU^Bcab]+
KKG3^C:NFDE&.66\AHMICM9@Xb-UMgNTbBGG8TUJKddKNXUZW3)\82^5B@E1f;VY
CMXMM+2+ZJY1_^M8GWTR]=A&WBS\.dZO=],==;Jce,/]K7E:XVXa0b?;ba=)>L?@
\,VKaHD<F>)^DQ=;.(@0[==OZV0?XM?I?0O^<ST]W#gbX]2H0I61CZ?eZcJ>O]C.
#cEb4/&U)gU_cN2)JdP>U@d<BYVVDe9.@cFN2S:,F)e3]IA0d0E=\TSIA=)K7PNP
6]9f+5E4#L6,O[,8/eAXY3agMN3=f4M=[(TL5<bSZU167Q++Z?@0FBgK^7P0?T4K
=:GIQI_4/G\YY)2Q#44MY@XEO7FgXa/<31cSgg&36a7Hga;b4B#1:e#=-)7J537.
L^-GM>>3/7d_Eb.Z@+#3XeJW=[,[W;.<,GR&gdZVde]ZINHL#)BZX9ZND-/8_\=Z
E[d&.(LXB2IM8L1@SJ,15@2AP,=/9NL@24EKD,\G[\WKZa]WC2f4@P?=Cb(@B70E
?#SI&eG9(gJNN[NVgL8Cc)D5EJVM>5+F?N,Z.NPL656O6HC7T.-CBG]_/:8c@XP5
]TPZ6PJ2G\1&cdaTM1R+Qd>a3YIW:M(,;;XN&c-BI=?&U5I]GO9e2?+\JgOI)/JR
/:;Ndg&e)YV.U(c5@fVF<_eU>J(aMI]aSM2F#-#)#08Z\g\d.=fYf^WGNbSWIcDM
A9@?8R@OOSZ/G4MJ3_b=aD2aYS2e=G(L?HFd10M;\=:2=VIJ-d@UcG\eKWI;HX+A
QI<PR)dLYQB5/Qe9AOCbeMR<@cH],IP\1]L[H?gS1e^gA&+\QHL707g.VH^&L05.
Y;?;F[-29]RE;_#0a35M-L_BA3[-ZCL@[I8VM>?W?[c1Ud=],WAPBa7_A,4DYY@\
@+HM=?f#DV;7=S-Gf&F[OWPB-;,>)Q#D?[(0H#<fEE2M9V:.eE?SWQAW>;GCPH\J
VC_<E2GR^OWe=:(6WdQLP?aC9D_V6Dg\]]+:\(8CDK&Y3?ON>D,.JS3(URWHTXf>
6DMbRA5_0P>C?:C9e[E.>LO\,6d7_V6E);)fT#TI[;_KH_Z@6]JcHN4VHXK42.Kd
KD>J.J<-Ze^:)5NZ<bF[->T#c.W5VS\FFI4.\3.M3^^O2096#U_<beC\gC,>G&U^
9=,d,NSEdN3@:c(YO&+c::W=P>EW1L557VT39FK\+.Ze-Q+G;gJH]U&T1:+W;NO>
J=WB1#Z1YdULTJP,GB3]D(/E9J5@++8b,2Z(/]RHYIe_7C)DaBRAcYCdFX&5:IXZ
REQ^6J.JZMQ9F1&RNQaFFdY:YA1HO1Ab:H#(;W3NY-Ae4E^WOF_T9N>I>cZGT&H4
<RVCX][0LX)YUML(U0?>72/H9fGIdT=1Va0SOKBE3Nff2VCYDUL/04[M9N55&EB0
&ZMAfM<L/7gS@^P3Hd?1X]2=8+OS+,6<]X<ZIc.Z8gRe6CKTT+_2GNA>]II4ICXa
XCR#8A9JI;]6Fe/_eU(\JP>?59YYefQbTdS:(EGeAdfU8^HFF&ET4_V((WHSE]<6
SQ[bR&8AKD74Yc=bP178DNJ\TA8YM;CQCTGQDRI4TT^fAX\V9fD,V21daa)AXdHe
:]AI)L?Z=f(@GOF,bbMHD=YTV,0JaYEYG<10?E4^D?>VNALX7X7.YB;d^+?F,<>c
FS3dWg-Bf,4IC,E@VS@)NYZF0Z]PV@>3Ne7DFLf/9b&f94ecLbfT#?D)=d_=3>.H
a^g8-G+(Re\;0[:<(-c7=5@;3>P=NAd,)C^++XQ&D#K<(\FCO?MD_=F(C&3TL+9.
>8ZAR5DK9E:A/gDUL6\g>T^Tc1U6VU9/+0/Z&438Td@H6V::FR?4f:YXg)P#aXO5
:dE/dWd0,W91>Q36R5+CK5ZNQ8/3^==)0\HNa5S:#4(LN0O@NOK\A98ME?C4PS+O
Yc<H^a8b[W8g3#:T&-EgWgKZ1((M.VJP]\b0WT_^XgK#<101Gf6QKaeN0aDI1=V^
;eFVJNIZ3TUdb\,@1CX=d@U/L7N<<>NYN6-YR;?[B8<Q7+eMe<DRI+&=30[ILO:W
,D(d9Q2P@[a(D=R=RDIZ_R8_76YFW6[,M\a&B5[E9ONWU(D1UXYK7Z^5C0f]#,1[
M-\8?(#-J?:U-Eb(:YaTD^6-B[4cLJMZ)Tf6XMADB+_82K^5G5b#aX+INZ0Ub.0<
-6J)>aKMcgAFEVb(4JeJJaQH60AM]\&?YPc63;U\68>EUKa^[McRb&G4C<C0fOWW
B[KbTaYO[F+3TBV88UE11C=G3@^WYJJ_W9:=21^Z]Z)U.C\6CFf9cWGHS&W470X1
0=(X/&=/PF\_70a@H<3N\RZMTV:H]gA?GNWSg:71296V#eGddS#^Y8,423QKc&]N
T1G1G4OG402ee:YEJ?EW-W=+W)/#+&J923^8ZS01\3UI?H^W_dZ.Wd3SL#0JM8>S
]V.MQG4X@6_?/DX+W^bC(]fITb+PAR7+N:0-/aPS&d<e^.G.;<R,#/S0=6_4Ne__
BeRW??^<)b4@=3a.FC9)M_dWABEU.R&CE1.-AXf7\A?g@#c\+6T^[P?8F@U./02L
N5BV^TRc-TC[]:/1@fZF-6PC@?R,,KM@@J8K1_J]38A36/M;gVN#.JgFK@@2O49-
N,T+e6J6,Y^003,/IfcD>5=4J&[RDA^VB+2US^:R([TDf@B=f_&N-c1CLNQF/8\g
9IeGDJ5&RYO#@L[=>>[G[NQ3H6CS=KCL;83<9XIEC#1H.HaUK5^NZg.^<3#e4PN9
FS9Da.F-ZMfeM6=-\S^A19\&#YAa@MgeFc/2R-;<R_<_#6G95_a1P/RVEOR4D]DR
-YQ46A9?Af@O]KP2[?+##dRTTg9IDH3@>BWU]I8U,_:6E,Q3\U@JCM6&P.#Q@KWP
3f#eM?JBdD0c5;78X4c<VV/4O2=5KHeA2)WZFJ4&<\_ERNPC/?3YfHOaXPO-bD7X
baH9G\R@V;&1<-U3g^U]_cd6BRNg_/GTf;Bg87K<bM)LMH1Y@J>Q(MW4M5S?WR(a
FG[?0/=Z>)>_60A4:MCfC)7\C#aC>DF2,g=?QYCB_2^XaW6aV@D)XL&A?(_5G.^.
+4Nb,,Wd2@J92?5VG2\0[GF.HH5IZ2)4,R#F+9AE.2NP6(gdLU1NT#YYUZD#IT1d
.S?eLX_A&Gc++M8-<U15RFW0H4=]bXQMW)_>ZGT2F3NWHW3K1gcb)D1V2@@&[/2X
\+KHDR@IdQQ@^UfaBcC:6T1aQ?FSfS,C^UB0T<W./a&NU8b\WE[f&+-937,J[--^
P)I(eNHW#X&aB<IPf9H?Y@>99Z=gS)0bcZ_AEKOL4T&.U@\K02XJ@M?>F:g;BA<e
_0-X+]Bf0d71e-[)Y.RgD?4J^AJBETUWH=_=F?[LHZ^Y>c-RXHTA/O;2=FY84@@L
[C#Ed;_[5LNY;)RegX+M(LfU0/M<_LA908S)b@.B.K&[.U7eWZ&.dVOT=1@)d227
+9V.eX,_5\;Q+O=K,KQ1A)9>C0/=OXE93S[9SIMFVE+K;6V((30;;\J8N53d4\#N
VLbFQ)UDV:f\O66)(4>T#[T-;IXX)gR9fa59K7@H109gR&@O[-Bc_T1V<(QTJN#+
N6(gO[^7R=-bHHU_#ME&/Og.V)7?@FCVgG)/0_5a;0VH[2gaf085;\4CB@Fd_f7/
MIS1?#bg5REQ^N)C]YOa_6C7<BFEIH3)P9fL<HG.0)&L[BU63(:]=RHW;(L<N&8F
M&.1C#&0K/+KYPJ(#.A_,-)>_UW?__bRYOPON4M0bW12BXLC0C^Pd[8U&.L^MC=R
3KX&OJ6ZUCQP4?EcL=VGN-MRd_->EZ19YAc[X,7;e#1C+K.[1fMf/P/N[60K+M@B
S&V.0Z\4a?T]LRcC65&<Dd0e=1_>b(f^0P[Q\@DU#^da&_g-QU0+TBf)37?06-GA
9U:F(a2_U//DA?2Ec5M^#RG7NGDMFG7976d(9X1Z=6]0&cAZ2CY1QKQDL:.=\aTb
D3?>#b4Z^D^7C9:/8BI[X:JG]f8_g(ecV,UXb,ZPZE-<@W^Z-6Q8O3SGaHBe9]8e
\MLM&dVOM6M<O<HH2;]2:GACFG;>KCS]>]C)^YGM,GS3LJHfGI,CV<>:[]cWa>3W
488[/.Q>1VT/4Ef-5>1QKfG8TX/\aU1ZV_P/\2gM?SI<?6F-P.1a.fVYAB.FOX\_
B0.0L84df>C:HQe^FB6PO6J6SBSY+1+Y_T34Z.4<#7E2B3)N\gFNb2IJJ7d(&>_8
/I<]3-[25=@O4X@BZ5.3DOd9YW,_#5f#OZ?KDb>PfI#R/,+_808dZ0QDV,E8c1=6
fU\/TK@A9A#:6RYe8:/C\([QO=^/P\<7WS;U,S+/D0(7#)PM6,Zg/?_baE5S-Xe#
/2\G\OJJT@UTQ)=,M(dD=N+V46BVV9-P23]&_>&aSI,::22;],,]N-e5M:^eD#7>
CA6>.FFAF\YKLG/aeK0(GO./=4b@Yd<PVDJ1]TY=KaL]TSV5(<JC86.a47I74::#
^c?KGTL-V211ScL3^\GSa\@03/8fH)cNGI8WX_;eRKXa6^LJ;^G9I,V7H9[8EI,g
#b[7X/Q<KN_a9A[G)gS4+ESU7B]=@DV<W9Q<47gW6QTK_bZYF#54M0X1,4O4IF&)
\,N<bM.,QfB-E><XfLB\.6:bI\;#9I93<-4H[BUU\e^)4WRUMdDRJ0KeE9DA=TQP
g8NH>H:YRLPH#LJZ8\H]1V>2DINZ\@c(P7.L)GNWVDAJ&26S0BFd/]dQAZ6FD+aD
8@Xa9+5?9D11DQ/a_63JcBYGA>Rg)5.D;cB9?G)=OO,0[_MC,#GM<-cLc&CSZa2P
a\J;D@?F.^QH.CbYaZ9bGVJW8ZD0#(6c1@>DI5)GIN4NdJG>U>:d.0.3SEeZDP4Q
<^EPOJe[,bP6Z6/IMfQdcTJdRZ@Kf0?+@N38E_cF_eCLVb.e01CK4Sd0e9]V[.RG
17Z101HI;IE\FA41H@C.,)eV2Z2ONU4B&JdOJV^aB6UV9VGFS3^GWTHC1-SaP/\B
cd)K-=-23)+W]CKfb_SHGfa3Z>fcP\M#_[8-dgE5=:KG5^MDb\/4MHOZ(,40:I^T
75A=.b4g,:g,QVR9T83FGR<K^/L/2)BTC#2O@Q)Rf.g1ZQ(];aPIbfbN-f&=-\9I
J6QU?A7GN/@FV7SIO2KGAH>d+WG^g2L1S<^E#NCb_3;]O\JAN)c62-CL1B&#2,?;
DY5?9E@QOD1La?I862:BIa/dP<8de83KJYM3)K7SUV4@-UDbe#Q)RfV0VdKU^0a&
+b>BH:ee.e:;U.=V1:U#=)ODMf6-OAILUU6<0;b[<?9;H1/f82U]DFV?M;9ffGe+
<O?4VVQPN8>cBM2J^8G9#19>K0+>_BZ<dM^;CC=)8\L\aY;X&G/\EL,^c;f0+POM
:M4_;UQDPQF#((N(AZ==E<LC9aRF=EA2;+GRB@FREbeM3QKYgX\[8=T5\Ud7LD:c
P[C1Y\;DMNg9/.)I5gM?3P0DSNGL;QgQ#_6b4G>f&W3-<>6)F;KQ]BI<T&NY.4K1
<XN7OSN6Q734;]/1SL;P#;(/<BPLa)BDa?UZU#:-[_QIa7^Ue;S?Y>O0)J3Ee8aP
H3&7LSbYX4>.HN1X+be)#VY#;UQ,;P/M.AA:3bW>@3PH+)I[]XX30e-F5.I9>XW.
E#2AI4cDgebEMa,f.^8PD5\AA74DZa-f@)dY;B+09AaH3g@W7-[9JPN-MXfaK<64
FC?YG?SN2NR+OH=FTEdU,TEKS&^IU-gYK&2f2QB7fgdKR#)H-V7Z63.G2eAG@6@:
MeOQ:N=<-ZTacRR>Q,^1OaURX0QO8B^]aJ8IQ:&LJPRId8_&ZY?/f1fG2\E[#C\;
O8DT49H=^SS12[UPC?(.7,?A_LUg;0/4cFJCcD^H4HL=8g/@S::BaJg73:QBE&V;
Kb1_SFIHFgb(^KBS\+^Ne.]A/NJT9+cW\6bM(WTRV4QX@74X[675.M:8T=MgH349
JA610CT]],6R\QN-=,T<3(J<&/f<@V#Y8AJTKGK@4H28J8-CGa=_4ae)UWg.Z0Oc
.]62UgS96U?]:8Z][XbGH_97NE)+X_^#0ZV_Rb1ALNO<0I0-R9;\_DWg8,VUeGd6
4);CQ;V_Z^ba+dRBa8adWcG:F.TUK9W@@@6^JV,RC1BLTb\=TQ<J>G,S^1:F_YJX
7XUHNg8a<L>77Tg3<UCFc-[(^&>)UR;:>7F1J^e#]X[X#N>f@/TRf489HTE])(:a
./=R(BNL;QI/TA8cP()?bNNM9gAd,9aMEJ-a[<]Ae,4P6dQ1CFLDeRITbI[L5[^U
aMO)7ZS-5SQC:3#Je@JRZ@fINEYL#N0e.[-6+gM,NVRT#3LfU+ZB8cX4&O#BT?2d
J/\a[8E;0P>7SXC#?-JWXLBa_c\U_3JWJKJG18MdDML[BN+.#(/D\2W4fR(^S3<W
X(HCEL/<Q(V3JO\61)J8=QG^^30K_01DW;#0<<5^H#Tc:2,&Q[:)TJc@L<U0<94H
@D&/SZ,7NV>4HS3HQ]b5Wg)CQ_B?d,EC_5CPfb8?_+c44UIb+V+E#SW\EKAbDJK#
?aZe5?&U306FM),\aNcZ,MWTJT).:+bb+)#+1KcF]8Ce)b&1;F@718d:Tg1BC7Eb
^&c6N4ED/VgJ^dR94:>4?8a.dd?b>PL.[?B.c\1^>TDKJgRM<R;0<;eV&42[R1?6
<PEF1[V;@PVT?D:4J/V;\73@dIJ^TK3fV31Q_;M\b?1I/9U,_D+9]bI8G#cb6]Z,
#Qf,ePOIP5OZf]U?.eB=bG5FP:2?9P0,3aLHS;OJ/dLa?d1e^^ea(H-??84g8L84
FDH@NHYYH@B/9@I@b@RdLg3)SC\_+2:M<FWO)C)@E^O;-H^_:(V@BWc83>e5DMPc
Ag@bK.NY5(X@Y7&C[RAGDa/KT1b=Xe\^>-F+>@+K9,]+6)Q2K[cN:_O/eC/e415J
@1=W0Jg/SOd;(b/+KBU<GYK-[[&\7aA4cdL3]5FTQdfM._SVOI],QD+7eaN9>gW9
70\]U+PB<[_2-LETOc-2A[F<g,62QQ=Tb@-\7A0).EUf6O0b/(Ag:Hd8CDNTf#+Y
f\[fQaaX&dXG&C0R^:Q1-;NWX)VC&QDU;Q_;YS#JGNWO&3?8W5]W]73L7A\-BNH>
&D/XK>D]g3B#Z32=1^I5B(_TKg7,\2A.@K-N2CRb;T@eBN9?Q++,<R1<+I/#9b8A
g\?W)NeaH>bR.We)3^-9Q#HHegP-Xc5=2A#&J+0daY@e2O<-\PP(KHf/Y(SeLUR?
Cd/63BEN4&cL\cHR_cM5G5O/W]#bKf9DFccM#5QfF+U@=D9,NU1K1=AWU[2:,@2F
4.]ZB=f5B1MaBaUHWY6^AZ:Bf5gL-Q4^P_]JVT,)H?DB]EXI+A^b#6_LU<f<Y1UP
aB0>S2_9Bc\g[)@V.QTf.RAKdd7AC4P]J]9a:6U-1Kf5Ad/NHBaL&e@O=@U[Y2-a
/>D=7KGQETdFgPY>/c[F9Y2gJ?c>[V.5<X5VN<^f(P7I7VQES<Y;eR@GA4:&^N<8
:NTT9<1f57Lb5@g&0AU8X4KOU+b/E\X.FK6IOAW-RDDT:W?f#a<@H]:R@2BBP8=U
+&fE?@]<J65&/c5:7.6ZI@+N^D5Q9N/\^A6>Ig4:H:c(WD>L[4L@5d/@MT#WC6?T
<]K3;:P7_<cP\ZZ8G=U00P581OT=KYT96NWH(g)T.AQ>O\RHN5W?H+@SG]?<#a6X
eZQ5#KWMO6[[6;7/LbYg.K5CJW,0B_-WR4(8fRgAI<Qec(AL@@EXd<8?+RVO_MDV
(L)dN8g-VH?[S.d3]W--)6S\9T/]0K+d.Y81B@<N.]\3gc#f#cA0-ed968A:Ve)6
S=afMVS88W#]>&K;P,-(<d7Hf/@DDH.TO04.Va0:Qb3J]aEV=XEUb-](>(N.0H)8
M2TAO(1.e]S@A--3)9<6SO2_T?[I#B\X?9,Z^<3]E+&;K;5YO(CaLR=a2c4[>PNY
.XLfMMcO#]/@?SDY]F;2>X>B..&QJN(5^A4H[MD;8CgDV_;ZW+J&W>-R(AX)UJPZ
Cc^?+?aF@9[>^0CAdC\0,==6IG(RJJ>HWK^+a@bU=)WLg2:9\dW+c,cP.Rg:0>PR
3WK2RD7gO71XM5NJ).B2CacXc?4Y/>Q#0=^E)Q_=_/a+E0D_01<_XeV=T;OLZKMY
PGGH(<C#UK@PEPR,KZ5@B-Z_J)9^@5HHHANe-<&+9J7=>ATRa65N0#_/KW+-fTJR
7Bgc-=S:QbK6<=L<0>4>9ZP;NHKfc0[cQ1)cWAIH3F6Y:916d2Z7OVE^^GY=Da.@
#RR322X+gB@O\S58g;M&:gL?><6_RL5/UK=3MYWKf-XC+D#5aaT2/M#]eMV5\@O]
H0I(&;5K.SAEDb/Z?D+0B-Z,BH;+eJ^;+U2?[a#59d\AI(@bALZ>e)\E\0BQ:Hg>
_P&K:_ef8=1M0LWBNd@L9<CcW#09.b<&60SL/?D\aW6=baI15E+()>/N7#6G=CTe
d.EgLdV.J[JN]aXWCAWT[9AEZ+NEN7XC@d3)+Q;#PbdA;#B&dODC@b<1.C>UO\b:
Y^JW])L+K2H0ZRPG>f44DKD__?cA@6A/4J_O6M:GN5<4J]KPbg16Nc;1->1C7,B_
5;JBgEYT_L;:SLU+[)e,CcI0ZS_@Eea6Ng]W,a#ETB,-DTdUQJH4aND\Rba\(WFa
:b-_XF=N>WOAEgF(BO]b.CZ3:WS0[[,9ECcA,B-8,=P[0R;-VePb>,6@)UE[=0b>
Had1(,Wf_:M8g8?]H=0#W?0:X(BXUZ4f5(-]O[7.M?8P(Sb:ZK?MKDWLPKXS1GV7
CbOV(SM<&4Z4T#),;CG.]&@]^BPM@X]G/MdEf1fBKF90O)>(3Y-P3#9N[Z([@#I4
PA\)7ME;16>W&:+aQU_QTB9gCLKUH>BJ,c?E:bBd?Qd]48U-[>(.Yede^35VYU#U
cOc?(3ITa/WLEE.LLd9<9-Z>CY/MDcO4]gP/(8BH.?VA)&8KB,GA\E/-7L&bL6?;
-DX^B\Fc3Z>WMa>5A9ZAV=(MZeY8U=(\IFfQE03ZRL.2>5E:T]E048H4@5+G7:;L
a-=\P]TVK_W4C2_VR.:\V?TU(MQEW_gPd&1TCQKBS2):gLYbb1MbD&@2WOKB6F)+
HGU68>fVGb0214R4IL7IDeUY>3YP&<fKgSg5K1g.DU[DF\[;:\(.0_;a2XL]3CFb
e_^_A^#_)&WZOK=&Y=@248<LAPRf0VZN<XWE\FO:;]ZISVDA01c:)NXD>3FS7I(K
c>a]2NAXLI1b-](85U0,XM6[gggB[:\>V3#]b_F_I6_THTM[ffSAf@gEW@0L)&&Q
7A&INGGKeXZaAN>g_7Z4[4FRF8^(W8)RA;bgfRd+fC-.54+g9M;8D9X]@@VGKX2Y
WBK+f^Y+.Z^&edZ0?^>><Mc=@>IXP>DTQF(4fSATI[ZX^,=\5[ZDKb?+<7P,:GI_
9Y7S.\bNEFD4]B[^c[1FDbTT;>R/-LG=f65_gP]#dBOY5+FL>XY:eZFgX4AbV-0[
D;0Y5D8g4[feWV]/=^AB=^;;K6N2d;<T1FD23LBa2=7/3=0F[F[\Z_7-0V0>/9[X
<H@)CCeL9A=0;YZ<XgEg1V><+E\V1bVCDKR^5e0MbW+8UL13d8Y27e57Z:247N/U
b[RM.;[7KAU<<ZMNb_&2\PW5?a6Q38FJ5GQ<E5Z7^=5FcM2SH14NY)K+;Z3.))QI
GRVHY#7O:Q)+LOFE@^\64I#=M<Z@[J7;_)257M/KZW-@X#>[d,=6_VT5S.c:U_eH
Z]G]D(e(A=O7P_#57RfDLR&K#/S@=R;V-LN:eKfQFWKf6:2.A9XLH)\f<DP7<I_:
_3XO?MDZQ@_7<g,^<W:)F(2.Y,QW-T+fE+=8,H=MLFMV7cXf);2E9BUUF#10HdVE
3RUcS#]5FcQE,\eHES72_d,.EM]Q?>g6KWfD[C7N20;EG;@gK6EN1)6L](NO7+gB
?O_R-_g]HM,:f0Of#fXP?D4B#HD5ee/^-@8I?X4+[A@V5V0+gUGVFGMA=2HEf6V+
LVaLD_6EV7T1L;I7JBHF(OK_6MY3<WHZ0Pa0Ge=g=FfBWV3c;fHV,&=+,4Z@4D;B
c497[F:IQ[_404H\[E5SH1T\NR4JLCYfF@>)1(@B,a</AO)O?B3eBN+_78>G9JW&
fV=<a\_E-Leg+-dc2@#eR64LCefY.FG,gQeY:f@1C\d3E>GSJ6J5D/@4A4[H[g\L
:AE@L,CeL]<@Xfa(@bM?/[5Y-K8BC<ZQM#VDYBE.\5AbAL_D#H4Nd7VV+0JJ6a=c
EZAMXc)f6d.Fd49=Id9Z3I5@dTfb2G_12N08F;@8Q#PQ^5(I>f/^5>NTaQ5TD8><
F:P/-d1D/_IJ4a/cD>>;+(9I+64Q52e@RXdd<2Q_;;^aGDA5SR3C@6;9=U:3&6#(
=(#H],^K0,a3B44_GE6ZT/=Y7P1#5K,)Ba.ZIT?0Z[PRPP1;cZ_QUg?TaTS7O)UE
3\>>9TY/(+@424Q;Y<0&8_&#B\(QVE/ZBML\EJ@;?f2GZDT<,UCPYdA4?bW-[Z=[
d5g-G<F_,=[[3:Gf5.:fG4:b=QNK\&W2ZPQEVA)&G#dGQfI3/)N-?G2)CG0\/NX<
XBg-f5^Z<SKJLe30;NM;TG1\((dUfMEH=-9b21CeN7c@EbR<B314geZB7KW9_U/P
):JE<gJB7D^bXJ8d>c6.-cfU@S[>W#OTc_UZ;,6B\IF0]9X1:]=N^ZD9>VCL^G1I
0FF@e@95Z<&<a-X:\L0Z^32f90c[)@[?4&@@PLDD1,J\O7?^5<T9?.,71AKaPN<I
Y9?,T+/9/??:AC<cYFaQPRaagfF]715b\A=RF0Bfd)XHEIFQQ,_\8LbPc1db&=BP
e&?>HEZ+Y1/YG4XEGdG2KJNVdLPcSbV-;e<-FKE&?#]7][YbEb)3\I_B@f=QW2Df
QA\<6NFUM-(>\]4V<,0M@8OfGeRDO.VgM2g2bM.<9VCH56HI?0GeU]bDFO&TWDGS
AT:LOaGF]AFWG[:5K6E[A;N_8EU3>8:)eK&VVAU3;AN\SS/.eDX;<d94>aaW0R\H
KF)JO3N?A4\<(PTBM(\f^#1-_=,cA;Z2_bfBT):7YY:6@_W@MZDAK(AdHTMfRNU<
a3J_+V(dEa-629MQC1OI\>O,C=.9>K9)F50&b<;BcK<8)IJ&4--:INB7B8Rg)U9f
3\VZ11D+(7/B:/[QPE8e>.-[=cQQY;/V#AO6+)MJ=Y?=Y4V@N,^J0[=de=eHd]7E
UQOb.W]\PX7IB&@Ib0LVQf9YI[+BI16\:[8LBCE3@Y>B)4;/HKFd8b(f_1.5H.6g
L[SS7ZUD.=FcIU2+fMAM;Qd:-7G4-a[^(Z\Q:WF=8Y^7FOWKF_J>O+EaZ&&aZHbe
/1_=?C?O\+caH;W:B-\[I6=4G?;W&4.ZK+H[C5fgZ]X)69A>_5a^^I.Pg-f[XRb=
YPLDA22>V_90JRKQ7;U5/G?e7YH_NL8B[)=dJ9df7IB5JA)WMB+=A\/Z;EXdLN;S
,G:7U5JU46fZ(E\XX>IST@#dfRVAN-)]=4452=NV?]?_8MKf80\\\05JSD-C[ZT)
;:#bROT?@\YBO6GA,CC?(C8JdIg9RER=Q7&VOWZQd]HL9NR.>H7#=KFYDK#6-8Jd
-J9]PM&B&AaA]-8BYgE3ACX?5K)YJ18?5R.)a_E@H,D9H57e.V=7QN_/5R=P&fXg
LNdD2FaPf@dbG54fUSN/XF-EV>1J.?&df_dePEHXbA#Q01V1dCd3L]Q7Na1D>O(L
3/@Z9IEf;f7G;>X;^RDJUEJZ77FO>SDQe_2EeX7D3O3[#2ST[5XcZ\DYcYSWCVHN
/&9#VgUK0/9^d[D)XLY.#2VJUOA)1\a(CCBFaWH-g>C;OHD.8Pa3KO,<a/,.=VfF
=O<Yg2BKX(X_eKVT5d\6O<S<?0:e=BW04U<VT[Lb8^IOHM4/]bb,\SOA?-[LfXP8
)+V444c&)V^H+.0NF/EI&H=#XeeU31/d@0QJIAM6bbf0B>]DZ(;NT)b0?-WHPBJE
FY-34d.fP@>?O6F0:8LSB/#8MG0P82C+:F\0=#[:3W^YWCSKf\0DBX]JgfG8DCL8
Jb+W8SMFIW(A\8b7ULR(8N_<TM;Y/DDC^QKB<VdMb5-PYH0cYR:Q)&3]>O4aG#T=
K8\_]V=BDf0\D4QKD<+HW[@[Zb-OXSQ+S+=:=a8V21<b/)D>R@;YW>bT&0U,A7H0
Z?OMJF/DS3)<eQ=?VS#3f<Ac1=)P]=\FV>JI&SGaQ:B(^IJ+2,W/+.:VM25ABKgD
)B9KP/.3A5MP42@F[0[\P.C_U=S\KeJA>c#YF^W(1X.J_GKX^^gdTBEg[=A?T?H4
McB&:+S1NU2VH=8aecHBN<PPGYXJH>-KKU\G>=4ERd3#3E3&\B\Md1OB.L@C+_Be
C7=#<3aVGG-]YHN):b@L2XWI_R#6V#LIg)1L7<FA&W:J:6,G3[<GWE_eeX&,5dXC
3]Ne7??G09)RW;23C#<#,fgeOagO.RY0)B?6g08]O=?HRL#:5JUB=Og(Z@K53._#
FIOBSCX.L0UY(fK73O4>12CJ1FZ7:@EB,AKN6NNYJKR?^;WgPT.UgZJ-YeOH3GS]
M#,>XERSB&Rd2d38<\ZgKUTV=B:EDAVIbLZ+O/7=DTcBM@^;6/8YE^;.);J_4(F-
A1EVL>+If5B8^5?(GK<E6Kd+gdH(O:43g__TB-XKO]E&;@=FQJcEL:8Ad]^X><AK
MX1H83[:[XRAa;/UYA,=YfBc9g3V9BM<A\WSEA#LaUK\IdWU/GN?AFY&Y?c7abd=
dbVPB6f(V;6Q)>N@,R=U3R#=[J]WPe/Nb4fN4.JT(^])6-D@>9bf3#W&_>(O55?-
KV&b_Hf9Pe(Ge\aHJFb)W^UL46T9.f;a:W>6Z;+C&bOe3[c-4^O-YT2KEY?N;WM?
J/Yf:ICR)<[89GJ#SdN?/+TAMQ6H=6-;37W?PBPN)UgRSZQB[M\)47g)>b@UfXZ[
eA#G[/e._:.W#=LbI-D:2P/4c73L4YG_N:1e4VLd-Bd6Q&PWUERCafVI0^Z+05,@
2;<1W:9U<\,6Y;b_W@PR7AE17\?X\=8GS:O@c6A0Ec4(Nf.>FdH==BH-DG/3ba]Q
0SL?OgHE&Lf@Y3aM,ZB.6)Q(],E3RLf@6;C/,JXc6ZfU\^8RH32VQ71g>I/KZ,Q9
L0#[0gZZQ<,<PQKVf<0RZ)25)QY_LM76A+>8+5^LE8?d_>1NgU&WD3M?S1;AUfg?
9<EA/dG=D.]A6ADQ0ST&@d547O3^8;EILH1b-BdU^@6;6YdY>FF8L,[.;1Og8(4(
L.UD.52_#;RT\A-BE:gB9NOTGYQ>&?c3ZJ)Y5.;RO]=E)KFRUTRRYC+,2O5OaM1G
PT2\b+^NHIHWR^56ACUGBKaN&9_#Q7dFNE-,_-W:<J1?gMXS6^g?J>MA#NZ\E47d
_Sdf1aC<a>(FY.U0_/D;R(ea6>=;/(?X6]V<=UT_U6A?4eD^88=\/D<f]@Q+]W&1
5[;b0SOQW,H9Q)U#f@XR6/>#\gc0[)5K+B5<^\f-(E=cJ;W6d4Ec+0eeSe0YE3NE
EIDP2CC5UNBOb/<?0NLL>79PBb-eT#UE)TR)[c0=GC/AMTX-5.7HZR;#SQ_R/U2_
W:;c\R5K2,HdB<K[d3WIM:.>,JcV(S58?,VX.),B>,:-fX&BR16UeALK<?EGI]T)
U)-dD#:N5R.F/XV-Z)]K5?FNdb73Rc2@58F<;BM6dG@.,Y]71->&EQbJ5V7M/T-3
6MRLP5gfP]/75W.Cd5F7@RV;80D_SVSSc(QF95PUgDY9Wf:+1O@C.K[3bbV[<Nd>
51_LJ-c5;_,cO7CF[Y:6A,OOa\VSMQWHS=OO1S&K?b-OH4eC9<QTR\/1?f2]6SaL
P1F::RcW8]Mg-SZ#/>LQ^@WC;Ba4:F8DFFN1WZ6e?Z&#KRR5^?>:5<],.MR?9)]N
9T1UXQe3G6I#Ne3?FJ;X..<LYSS>.U0J,V^=P:B(@(L,L[IA>Ag_5VUOW]&]IAcI
XEA3_S9[4JFXZ[58^b:TVK=P=S8VQJdICg1?KUdMe4YAHG3LK<dFZ;@5SKDfJ&.T
O.BDU/R\>H)bePU?/PHQA0;Tfcc4[BRZMH?(MOc2f-RS..0;\4]U;=]b7,IL--Y[
L:,cdOPNeXRW+B6E??KUB@KVT;5DeF0^BJ(_H#ZaX0PI)Q0V]NJg,V69)7K\f90K
b@U629=bW+7RENbB#V8_KW(72UZZSP^fcRaHO>8I^?:]XUJ6gYYVR>eGW]dP-X[;
D2DNRafHLC9E4MS^a:YF0/?EbI-7D,\AYOVc4E@8+Xc.<G?&95V42ITQb4R>0M;#
#DdPf(;Xe[75g8;C7M0Y0O.Cc0(fIE+b46]L^JBdW;g3D\4:E@Bb9a(_=)&;ET:I
7RG@@4(9eQWQY)B_:/dCHc[&_PSUTAU:,KF:V)[-1RX2^+49WIQ7TME->e<T&<NV
f&K?_bdTT.X:0bQRE>Q]QS+1NB)AfM_6IB4CUMSRW?6HYe;gX^::0;+H6-WH-\,c
B0@DF/#E^7R3?K+eVDcaEJKJ8O>IN<M.STL[))I<ACD9LK(Y7Ug\O0JcAS=fD7d;
@LMIMZ(,-H+H@IAc0aOP6#1GU=91eR:3++A.Xb337e4A>01;5;Y3OKT#,N.@+NW<
1JB,N<2Z+S.+G/2ARadY;H&<dO2@<J#LT&=3?J>T?DZ^FM&3e6KR,5A_=TXA_<eJ
5ATM-aEXgV1O[,+V4@:49QZbV0Yb>c>FTdK@c-c2:+E#AEM:3Q?6A8,3K99>gJZf
/(eFOA4E+e2N20f95+R&I.44gd4HcTa#\/0S(I4<\[U&<H+TM/QeB>TeSG;,9U.,
b)MWBHbbHI7CTSW7&R5:00bC>J_KBDPN]gVNTQEb[d2-cZB_.;X+KCM@AMQ0D=[V
O5,QAKXVOJ-D[T#Y;\>ef0T2##WP>5@I0DDS83NVW@UA7gCEK0.PMM8c<9ZM.3Ka
0):<Q7>;#OMI;<[X+&VENS,U/-dH3VJF:S)_HFL^ba\X=Y]3Q6ORT0/03B(Y>.]H
X11fIeUaC=R(9XF<3)+[WY3d:):]bbFQ]\_C-@=;&eW9K[0Y-XVS<g8>MWT(R4bb
>b9/fgPS7gK=WIQJ6#^ECV415d@X(eYd@AZ_8S9;AL17IC\Qe;7-NM>0)10Da4e]
aZIZ9_MFXJRRV<N9H)b.Wb#Q[Q17_X6A7?D\QUF4WP7S]JT[+OFF1IKT_QR8NW(J
B@G:T<2/L=Sf5G8_<2NbeT99;b&?)c,eMGad4::?CTL[ILS0BN.3LB,B1(O?XgRg
b5F&NI+eU0R(;B.(20#ZZ_e3OGN=e>#R78.8T,_3<Sb+f\1XN],LK._JS4@#^Z#4
PRPg>A^U-8AGQ2-ba22JU8?L9>KS;DKg]HAGZdPS9g9AV8Y\H3ZYfGWWD:32;g>^
()K5@X=L4bFJgO1Lf06RY_dVO4AW06H8O9Bg(MF0/-?+3N#=5N;.37<SXQ41ZKB,
O<0HT/.FGg,^aSc]P(9HQWf@g,[G&FS:XIgUT\5/f&Pf03,KC:OV#:J3a\4XVd/N
=f:C)#<>9GY?(:e->LX>c<0A&?;FRbQU#+?KJZVH_I<PPe599A3VW:NV3)GQOKT<
B?]VS\\D?4;6TBHgc64IWaf87Y.Q4FC+Q)8;BJeLAObREM]/JY4G[URPfAAD1M9N
U)Y:2CNS2.,.7(f2@:]13a&=LQN?W&T(\d\b)dZ4C#INU\HJ2#IKPZ_=;fDR9WaY
U;^JD)28:XNSd]KTR/K&R39b6D?D1WD]:@;8RLJI,c)X01fc_+KcGV,UgEBAD:R8
^=^7_Td(U1XUHA\OdSVBE4\c/>#HI5=f3X]BR8:FO#MOST7,82baXG90ef6Kc<7C
C0PD-c]c).B\2AGb_=(e:8&M(26WcY1+Jce:3cG>G:_6-TR\>C@bda<H:gd@;0?K
Dc6DcTB9)Z8R<#6Ic&TCB-7a9F:5I)R]E4T#J6ZNX^)V@HA028L-0KaR)<P@;Fb/
CTO,7=LOWHK63]a[Xc-)b;CXP+-UD3QGQd#>:+8E;O+::Y(^(g=:\b)&,6@#F,1a
]+dXD)?^fO,9.I[X_dB@fN:=ST=S.,8Of+V=Q(VA9&S&\KeOLbENO_c\8<LMg9@P
9_T7/M8PJ[?-(=:@9P9WN8fJ.<Q/:6dFeD4F37I_:-@-S0;B@,;[,cBBMUJR^9#d
YHIHCgMA\M=/NTG\e8VZ+JK9Fg8]ON=R<=2]>B5E2:)F?dMNSK#GC+D6@f9:;N_5
Ab)QO+75R60E54Q596VA.#M9CB9EdXZVI8141c,M.-FabX@U]H>VCF<4:8AbQRR+
Q6)SZ/afG@dKd=F).-#6X?4M1Y3R.)TN,HO8279aa+J-/ZE.&\eFAb/Q)DBS,PWH
.[gG\5^PNEARZZRS3LI?2WK+/CIWA,(U<EY4fK;N/ZGJTTI]PGgMfOD2bWfa8U\7
;1,6BLV?LDHaa@(O?S2cV#f)HR893\a,)SUCF/CbYR<ZN34.M#,0/\FAT.b[,9VZ
#4:.Z0gGW^1VC;eZAL,4f;\,KE3XVT-QE(71):HWNMaa?<?@RPET_9Z2f&b-1)M0
Ng-Y/Z4;c2MD--<34>-B7BbPO6KV#.20BRBeZN;d<]05)YeBF.VdF)TD;]Naf)X6
=Td+3M34RUIR5(TT+B3^LJF[X90>]WVYIO:H/J(P69J_Od]OI?HLb.?=AT7.#/9H
D#4HcCe#=RGZU&X0Z.dK>TOR;QfK(O+3+V5K31c5#PQf>BG.V&8RGEA9[N6Rd@fN
\DQ?=CCbZSLe+)1CEdF76gDD6T\F&f:BEQcAgG1K7H4cQgRA;K3>HN:T<TT.80@b
UeEf=b<gDW52@F;1?He=X1PaEXaRV8CV&f7@Mc?d=^B<)S8DD@>ce9<,3)\JfR1P
L[A4(2;aCR1Y0UH\F[a4+>@6E4-JZK=9e^VAG3K\165MOXEH3^G[B(R]Fa_@JU3f
#(UDc9=OB>39SE:;9L]PI1SCC:)=.I.71M-7+eP1:NYX(:g.Pd=Uf+X3GI8\JX39
.(0+cO\U2<\-206@S\(NMW3GLX6@0aRK)/g#SebG79:a,TNMOQ+7F:ge1BA^(G;X
=dK#[]A<b5UMIOLZ>I1cd7LAB[W_9HRNSSP2a_P(e6>Z9#[/:)dV+AG/>4\H.-9?
,cgL^<B/f(fZBTCG_-?W59N=O_@8SU=G+5S_S(A8_Kf2./]:[E:I+^H]X.?Z]C2b
\G(HYJ0TDg?4(H<IcPUO^UM\(/5geJcfd\C/^&dVZ,VR,6fYEB/SLP@0IWSAYL=B
6bP_1V0QH#,e&V&gdWYa7[1KefP.M^BIEF4IN^W#AOIcS^gP>-ZD,3BXQ_8b_/0d
HDg7^MMVRRc14c2+K2=<faaPS\c6;-,)7a-6f6aGf#TXQ^2-gf>fEaCQfXe4GM,g
Se-3>ME(HUN7b?KNeMHD?c8/E1RCc]+Z#=2Q#^Q=GV#Tb@K(]-Z;d[O1Ra4a;5+4
fCWf19:M<.f.>B@20f5_>cJ??;06ON&@7dZ.]Z4HNVMdA<]YF1NC&-;GGW8-:[V_
?-R]5-+K?D>9.R;Xfa[U_<dV2Ud=H_JD3Q:/K,J>T=YG.;1;:4@/5C<?Qcc=244,
-41X.<SC@)?:\/,ee.Vd.YMaE._9^Afe1M>]Z5F0I,=SgKcZPM>@Afb-cWK/d#L6
9a-a\1;-XCTP\M&DM:5#.<D@TJTdUFKd[eV?]O(86eZSGSLXVDERN1TKbgB.DDSU
ECP0.K(9cYP+OBf,Gb+dIO1UW=(EDJ[)45GNQX1b16=)/aeb9F18/+46(]=;_.\:
EMFcHF]1O1baP[dJC64L8UQEN6B0@e-2_GLL1HWGIRXf2CS(B74YXOCLC>a_Y_/6
UH(A@AMAQea:<A1c.X?KPd.)#)&9/0OSM:3<G5=P#f8cHHP&_U0FTN8fZ51eJE/F
5U;;C=>T@g1LDAIAU8LZaZMWaYHR@(VIIP0JSgM.+HffdPD[(R8M(=RIE&M?&M:Y
U.W&UFDUCJ?8>3J=GS9[8,-K(@cC)[16LJ;8GQY+)A;4GN_6D63C^4>D2@O2^?;P
RBO)<Vg@9Gd>^<8EK1B^Bd.W+/5IB#M&4f;[1OKc)9\94R+ceFM,K]]C2<0-Xdg<
W/=;+[=A22H3R#(EC3c)f7.;IY]Y;E)(>KV,+W<?WONCRQd?>K>-5Q[2gd9#>ZIH
/++,Jf6,A<I\OXdD<bS4.gG>V,0A_5W>\S<3Q0O,>8gdMBL6SIg,eIQCJ0+6SG[R
#^+#30P&]5Y2Qb-=0aUTD[]dDSeM-ZI:Z,7Y;_931EE]08L4927fdc3)QZG-W1@;
H9BSaU-Gb64fRR[Ze+M6F)OY7-<M\8<-A+Jg9MK-F=#^[.SEHB4I>9)XN(VXXf_Z
<#1V(2E@:[VD=-fIT_dEC^J.YH)NWZaQ;].VAQ+AO,/YJ:O,1<?Ue5Sf&#<9BM=U
cQeF1G_ADA^()LIUBc#cN[>;PL8d/X8(bX/KFDWJYZY^Zg0+A20/X)Je6Z;]N;(F
fT<BTPAIVeX_1/VCVUAC6a0[Z<-.dcPZJ]5<H?O(C9.6_<Y,#+UOF8(]#=0_SCE5
VN3)KW,.S[T:?&7J@Z5d7(>Q-]8;S?]L^DgX#a?dVXTeBbDIO4H)?2].&R6GG5[[
R^I<>1LAF_cMB?0;R@1R;7.E?I7I:gR4#A5)^43[d(+/5#<QON?@B<?[[>P[X-O)
YN8R2-E)4/V]NDUD^&5RH15@IfL=OebHI>DXZPR>R]U\_&F?@VJ+C-aCARXHU61@
@0d>#?1O+^TUARXQ:AT:W/>#4OX=/IFQ.ff&K06g&@H8LG8A.B0-IP)Y<AE2XGPc
9-9(;70MPTW?E)F1KJGD+AI[1g3L6=;MeBI<+32aLL=VYC=e=R.>B<>@6#YR-8Bf
WJUY:R??KUSMG?ZV?P4OfNPMCJYa5)T@&C^L0QK?X_Vd+JDfW0Ff?H>:OW-EdD.1
..D1_7OdB,PL7#FaK,@)9gSJFSK9/]97J<)aeC:GS41O+-9ZCY(fM/<dVQ)@/)>[
Ob_;)_Y)#MdC<6W2dD>aZ)#8\-2IQ[IOQ]UM]e+PS:f.1I,TgbE8]#ZTGU&C<06?
)U=HGfe1LY-f9FCTK82Nc-b,VS@R@BMR.6IM2GbfcJL\GZe;&Jg=N;e@J=OJ2#Y?
<eaUCHAF>09A/58=OZK997_T.U^6M\AX82DF>U72.07WR^;g\VWPXTD9&bPJeg#f
bOD>R<b?g]04<eW]gUUMb,<?9C=4^Q9EX3F1.EE=PWJGKPMOK7ZeYGeR[ZLdY[_I
,MP;Sg;&21L9cMC7@]fLJ60L]3CJd3@.bX?b;I1ScWF;>OF1()I(9]>1GETAU25H
0acXfcKYB;6A5:,65@GWWJ<XZd)gS#+_IA[;#K5)<aMAV8R2^@DG,,KA1,EH-XbK
FOCXJgLXc@EJ9+g?Q&]2gUe#f>eTcHMddS5Q4+PO?Af0V92<YHX@S+f#IE8J6Fab
caaXKTENYW)?EQd4/8O;;^LHe7942UIY6ML,0+B3]YR#[.8_eZ6Xc),1W-KE>N,J
K6LQ@D+>[7&F(SCE_YU9Sf9++8^Pd+LGb^0=cGKNI0YKOG.JAV<&1?XG+YN\aVSP
AeNO0D?T[eOBSCBebEEMIG@Y50OF#;O,9)A>WW&\6LIAc4@LK;:6,-V[DN6;F(YN
DfB^95:E/I9&2BQ02dZ\2LACDR8DfP2,,eJ_PW_P+1H9Q7(a)f1A&G7E\4FXLF:,
e>[)GCF@SaTa(Qc/8;KKN)/M.6:1U7VgY4-eTLFJMDBgfI[XKg;]8Ee[8+c,(^N\
<[8\4VO6HZCMZcO3Y7a7FbR-0b@SK@D:?Q8>Q2<R1D9-U+HL9;(c8,U_D4X]W9;>
e_69W4;6KaKA8L[S.R:ea3LCEW]<DZEfbGeIIB4B;b>\44a\J<96D6cbF422=1I]
&184[2TZ_^T]49A:/Y.OJ#.RF8V@aHg@(STL-[Ma#aYI<eS<_(_B3.JYFb>,3d(8
g_4(NAA9f28V[0K])CD8)(1a(0IR1U#E]C4U7V6(X:-gSN6VS^WOSHfBg:+]@R_@
0P(-C;46eB/b5P+_0Ke71&eJ0=:RTM.V/+,_?,5(eZb?2/YS3cX63(JB,5dRYT;9
c)?a)/Ub@@ZZZ^>^D#b[]fJHF)J;]R)J/]Xb0(X?DADV&#g)-0JGO?ZC5^Q+(S@Y
9EI[dGCV68PU_Uc.9RE<SW;45]]3IKaf;/#DK/,@^ea64[WQS_)QTAg9A^=.@L^3
+7\gLGdR5&3@(e;O:2a,20>7[C,&J#<OJ.Pf<=Y9-MB]DV4c[TS/K=.3F;N910][
SD))ES;9(4+2M)MJI#WaJ-HWA;D)KgFLBW?S)=>VCN[+cV2M)3UdAK^P62JJ#Xa&
_TSBGYA=F?INB>06FZa.Mg]QNW.Z[()BK@gA65(4NG3BPSNX0IWaBagH-6W.3;U1
d9_6.2]T]BgH-@^dCGOGOEV38OVdb;?G]3PaXJY8VZAYFgAZ7DO(bGGVX&?V37L@
;.QgaVR\I7X<D;F2Cb258T2E25>4__+H<T^(:=dP;I;]A67eN?-+>Z,d[FcGX^AC
5/YW-0Te(db@+P/R?U,2K7_\=-_,S4RP//.b585Mc>aI+FN>_S-DaO7#,EZY[IDZ
?JKNUN3SQHX\:BTV6#FRCKS=K7U251Za,de74C<f+GV(aN1(ZS8..TC/WDJa9=HF
+/8<8Q^cYd1T>9#\e)LgBVMH-Cg\0J4_,_+VeF[ca_#HgfS3J24TbC)BG3W:#\_O
Q-#]RJ@_?R/L)ZSR<aA.1b@@^W>NUOG[N)-f[b))S>ZM?A1N5BaW:4ZG[6K^6]0W
E75<BZD;gZ(D_8bC8J#5?&T\:FNMfORVUG+Vc)&3PRSSN54-@QZ865fHPJ=YRVO,
RaJ@Cac#aL+#AH(7.a72HL;C^I1[:gLUP0>-?Ig<1(QRTF?6]=JBNc?_@e3[#E7&
AN&OGB[cB8M3HTS[SRK6.W(G([]Z&?T05dFY_BP+C8#BeAJA>F+CW.-E0DX;Kd19
.==?SG]NWa8OZ?(-a2\7WG#NaECD@D5R&2TI:WCQWLZK@T]:f-\V+1:W\Y;5=Z(B
RL;31NTJW;B/[G7,3H]Q[OJg[<c+gVJEIX.7(5B-.,QV>@F9aV-IC_2#d1;4==HB
Z//]88D(/RCNWJ)80&3E7=gH7T]@D\V6YCVVHc9#gM<ecEA]aLLSOXGMd<B[@=WK
RN.G+VM(Ia]MLC+@bX;GR,-]bV;I1)OXT(c5F8TX@4-JWPN6GH7V/[2aIfW_5Rc&
U+>8W8LgH^PUc[V7-M:G5]:&P/E(&/^1g&bK9M:I:IA8/RKB_G-R&+1Ud\cAGcb7
-K7RFBN30\/MgCHGK#3<PF4O5S_,#,?NN-#BNAPZD;.eF-KN=KTc3U-3HIcg)Z/>
A_#@V7JZg:[^T#ZD+J,BL9Jd/,+=1YM\3S,V64]E&X4S:4R+FJ2P9d&J;^e]@5=Z
K64dY3c)3YcP1WV.L9dbH#6I7^c_+d5,F<5F/]19>@1NE=#.XY[B1O)H^K9(\Ke[
G&72.4Hb&R(Ze+EVVeB3[+Gb6.K@7<#^AR8^Z<7R#+fQ-\8,A:T66?b.E\4[K#(V
dE7d]72fY.a#K2#7>8_Ng_X7?fZE862ZCSU-#1\;N(;1OS80>(73d+MH>#;4W6_^
3Vf;B6).5HB+@-Zb^01LZ>(GC6#W>Yg[Z9(]]4ZW?2>69O)=&0?[;+10&#)6@_1M
-[7WF(A1@DBc;Z\6R+,:N.K/JRR1B2V=JXa<g7S[]E6W^6MNQ].A5XN;bIOX;<52
))<)P+\f]e(/VcfR0&UO,aT>?1c6gEI+S2_ETA:H[\AEVGU(g6Rec1I4Td=[eB8,
O&#+_N224K3_1S/fcc;ST#.LY4KbJUMS7?._2Z&6Ta3O]DTIJTf-S2>-FH_&<a.F
2?9^5N\HfBRgS(U>UR9acMM7&C,#4C_W<;>(bP3.,+80DY11:P5\CHg-eO:>F+fd
c4\dDMb)<(BE0YT)b#0FS-,fa9fXNRA,U(,8ZO7_0#LFU4,f^>S@deAS)VG5R5[1
f&:;.6HSe5V/5#JE,0TADNZ#F=3d+.W[,^+\b;OBF=ReX+5;3AW04(^fUga@)TEc
CQ5S;^&+ec:/J^0I_X#Q<gQ31Y>:]cSYY,H.RdJV&FYe7\@@+#SGEKV,W8))@SBR
eOQUdfQOZ,6IW]fP1<2QWa&BJ^L-L(C(,>b9:4SIQFf^WeK6]4aWCU0IM]FN\-J^
M;.f/>FZbT7b,Q8[+\)cDbH=BY3M-FHSf2).d=8-RQ<<N^:26<R0Ra86.&Qca[b[
[WULX(3K@]Z,<24,SZVI5&Ta7A02AZ,65?6F&_R^I6X?YdU:J(ES+JZ;@5W[P8>-
f@4ReNgV9XZJ1_2g?=V6#f[(J1PANUYHH]-SZ#feUU_KX+I+S)FJ</f<,4#<W>&8
_D]R1SfV/#FT]5?b\4^.KW-5EAZI7H.@?U==eg[OfC<9Ye]682MP5MP4&S)UD(Z_
KC.2g.SK/YD8JD[XTN0_EOd9VcM(309,28f2=+WZGfgBAc5:O@.<..^HI++@L^?(
RKG2KWEeL#G1B:bT\f3TFI.RK[--C.AH)<gU]S??21\WW_d[TAX@d-;U7^@F.M+.
L]N=/)MD:Ae,DV]c>>\LAZV3>VNgDW-F64WC[H25:0,C)5WC8#Bd&?T#A@<3#b7\
_Oc;8fDKW:6@4>-#;(-g81]c79AAESD4]NXg#=LP>XIVP7=DPS;,X&P+NL?W+6[<
e:63VO[S(5&Cf//C:C]/Z<cP-R#TRLFUgJ2a22W@gPN1dEK3Z64W@1_LT=f]VacT
YB@+1bUZ3?(M.Q<N,GKZg[e_0Me26O=ZfIX>?OYa1D=TAN_VWc0e.bJa:3OG_cR_
\-cM_V-D>M92,&(?dfBF/27dceR+fL)@CU_9:I=UKUeE;XU6eZc9M:)8ZBUdW_5#
<)bT)?aMQ0B0(W-,G9@C-g>[BdYd=^abBA8R2H\\=CFX^D9)0]5_>KBa1RX&cMK#
(_:/0G[eI.M(-\UHY0+UWL196K;dI-)85cd./>?5.W7/L@W(c6GHD,;O;W+7c_OM
AdP,f[28b7>1&S@/N(.3X\;HC7(BaCT7[CIb0BVfPM,6\G>/&:dC+RdE@M[9#E)e
a(53N&?#6><EI2WN1;+X#:VD)U];J8[NX[CfKL):1g=X6bb5)HfUf0OEZ#CMg3Y,
K?MWTL.?.e7-eF-WcL_2;FM/,PaV=]EXZS0,C_,\22C9#baA_&&AK)aK]_Ta3IUJ
3LKEaO0(=JG#3,4[7fIb33I=gNF\M>0bSMc[1W^caTPS9GCbgG56+6[<7V,\OUKQ
MUE5YFIcLMGadZP7c(e-)dD=Ic]f,\b(A&WS8A][NNHeQ?8N&f_=RecaNC)D<SW;
bZND5=6?NZ59(f-.fNfe(VcKY[]./,[f57?PT^;6VB)L2&JQK@UH[gVLHNK;2T?F
6=_9Y8J&Oc[.He^g(1EBBcIQU+=0e>]g,_:CS+W\W?N&><eA=0bWZPf^R4MXI2XJ
Y_\,HAF:MaM1M>1&38gTX88:WDdT=XJGdTa1+RW>]8DPLAb-,2M^S@-QaK4ca0de
5[>e1SB&FCNH>T78-RReQYQC3X,^8a2gbaEZ>T@ZK\@T)51[SG)<):Y-<g+AE,d>
?W/W:UGa@cO3-&\9\>g[8)3g]I/?SDG?dUGB/)FHU[,,Y0]QF3Dd4(86H:L(M&08
&Wg:4FH5B^HQ.S+>#ZU[aR3e9M&G@Q4UI-H(JFNege9-2([K9[A:N_>E[N3&MdLG
OTH2R)eF28GKBDc[aI9PCK647<ZFdICF0KUWfDN0f3c<5/-<FId68f-3/JANb\+Q
XMbG^MeC^aXGfK\1\d_QC)^Ga..G#L]_f&QB:;ID8=HBWO?)^6BggE@Q)P+\dCN+
P3d<#Ma]>)A9[R33B3,2_R][1<A^C;Vc41[._U.TZ5Ie4IOZP6\22RXOHH#Y#S0Q
fAF&\4R9QR+a.gQEeUTHO\25RAAR9^.gZaP5UZLA9.^g1YU?SL-_3_#WY@CU[_C2
J?.(/26WJM7996O)8V#QNa21LdQ:.ea18Bf/77?Gc<,MHISca==?bZK#-&&?FTOF
;UE>A^(57CDS@D(Uc#6Wa/UU@>R,Ab4ACA=Z)\.?_>AQ&P3K0fT+F1X..Y+8-Za,
-P1V]H>^=@fO)7&<JCX1714C85)bOLB-GG&NS47;+I=L6.--.gSZ.6ecT3.4J1d(
+KK33V^]LGCO([Fb=?+F^=\+;([Nb\aX6H=c^e9gG&SOJ[=Bc3+aRf(]7PPHS9Z;
;<^=P/NOHYVWBSX.-X]dAWTU8<?L6eXJWZXAg_EIc8cW>f9[]V.bd>6C5LI2;5)J
9M[bGf5PFfaFG\eGM:a_0@HH(-(&,T[VK(Be)8)^@NORA8U)</:_I+a&[aXM&0TL
ZA3/?IgE]U-,SFLSXM=@@\HRHHJV4]D?(ZXC&4]EY_#@^bT1-Q@fU>4@V,8ET9N(
WPe6_B^)-T2@>cFRcS0B7@Nd>398,cW2Zab&QNL-YWage3aKR@N3K<4?QG/T</#2
@SfbW)_\F-&:XdbK7<=]KA^X[1O:OH,b4C)a?9)9=@f-XW[7WT21#M6PMe(Oc>G>
e?6bLgF1I#^X1/EXYZV\;4_58/R\K4#bE(C?>II+eV)d,[CB7._&W_L>dW0c--W3
aW5=,/8IcJ,C21<KFde7b-)d@bNKR7]+QH/&^X8OV#[c6?#HV<#Lg3bbQdZ.Qf-?
>EEN&MTEFH8BF>T0/DBU84@X2c,d>33ZR3]/X;/b>2aY-HU7T)S#1V8V<7.N0Fb1
O7)a[d1#E<V@^-49/>;<:_;b<JW?P]:KL+E^]HbK.N??7VMfd8Ab(W>F&F]+?U]?
ZO\&a22L^2=N72c9#&AQc\b.X+#B1XHA.V5(70^MZU&eW-PIYIY__X<d7=6]E[Q1
cI^,@72OGPC#IR6@T^#Q?J(5X28,G&@LH3fX2P.da8]fWC^8]2Sgf3X#+OIQ^Vg-
^53Z_c#J2+[X,HJA.[H,.)6f?+JeX:QF<\39cR&/M&-^=SJZRE9<AE6G9d:9^DB-
gWN6)KE?B)JW6U1BPRT=\NAF#SJ@C#TPZS:b7A8/,/]:9\CPVaGHFB#_TC86^@6b
UER>T0-a\fN&:a8;f0GE1J+<5;YT?gG#?22^<5(B]0FD_/D,aMG0g1.d&-fY2Cb7
N]?S<]LFKL^QQd@U(L.^c]U;#a#08)P.DU@G<c<UG77I[YA#8?[DdLC(S@A1081e
4Z1(>?b;TYUNNNE?._9&cV2FNNEPYaIb^MTJDF._/&a@Y023\f\5(JbFWK-V?V2^
@M?G);fNZBL<M9^^gI0JcfB&1<[UU.Ld)KE5;FZ+YgO_eWP+G#7HO6D9.(B,]6Oe
]LP5,Z:@I5=SU+MT[eVc:f?^)?5IVD/R]Z[E=TXX=#9#L^0J;8e.KH_&&6TDSX7K
Q8]Q/d563]7D7XG#aUC7+T2QBOWMRI]=H_ce3=bZ?^cWZf?U#FHH@OQ9D9Gd@SC#
><Y2)@252g3I&B^c<fBDK,aMTJ,J0IGda;YJY#I@>(;/>=/gV).#CEFBZg2NSY>+
LXN8NBWB:_8VYQc-HGQA#(PC><7A]L4\DeH)-D4@dSB#Zb&#aQ)]</TB-9E+bT=5
O4>a&dS#MdaMd)-)M0>QR.GPLJ#Kd9c&X_&gPO>Q?ZF^5Z6/b26UOeM\D>XI@E/X
YUP7YWUf;VeCJ.b@[J?bA2BO>F5>g=CI44G1SEW]UP\S=]VJ097CU[(@N(28-Y4]
\UXa35W[PQWR^72TA>LPZ/ENFOdI:A4B\WM>U7c?Lg]L+38S<A:d[eN+J7dM<ZIg
3VZC>)SO,134Bb_d:XY0G<dEMK?1&AKG^\A[=]V/-_/IRUUa6[)\@e1,]TJf]1>)
F#NaPFSd[c+=BV?.2Q.bFe&=B>UAJ&aeegH+=IGVW+QG7fg,a)G/A5-QW[:+)RfA
9LbNUR[:B(OI[^DQA/,-U\^c<PCRHcLe&VJ4[F4?&02H4VTbE<f9,>E?GB;^SWS[
b;2V,9C9V>J=P>aSTZ7<0Z9M17Y?V_f(VKP)H;[R:8D,71FCUHed@]+1M\9&QDWL
#(gW]-6OL,++<c_EE,c]WV6<-YP=^QIHB+WN_&28[?2[?]6;H4ZBggcM0d-DYNG-
fA_6KcF\</]NXHQ#=V@RR3I]@b?EOOHU:SW3^bSTOVfT.77S<W,>X]BZ-\\O(PV]
P15Ia.F.g6,9:2IbFNM.WS)5;1MYUf]dXb]NUEMG>J]T&13LfDDY)ZTDO#?ZMK++
M0SD1U1B8/Zg6_1(72T70<Hf-X4N5/TeGKH2P_^^A-4eXKeUL7,8?F:#IIL+^R7-
UgFQfO9R?d/QP\#F;T?0dP;B8@c72[d)<&5=XN(PBQ\61,^R.^,]Va(N2<gH)_=0
d8e39_Mf+YIa@IgQ<XRT>A5=QG+PD&P_BB_.[1A2EJV&dLdX;Z=3M[<+>:^6-:.[
I@29<X\]J1_I&DHP;PX04/D,_S3Q9N_PUI0a0#6BB-d>-,TM2R,c[W=>5^[aXVb1
,X?TLOWV:8-8<,P597ge&MLg^;Ub_N5gQg4>K>WL:#U/ZS2[N,5@K,@-KM#Ifb#e
>J:7NN9RPL3^>H)d(ZfbF@c<FPRYRaBD:2(^S/&M=,0f199YM(0Rad35VIWG6DRE
0.N#\MA4W+]??FGJ)5-#H3RBN?B9>1OfQ6fKa[)<Ad;D14H9]S)<gD.FYSbUBAI+
/[,;ge&0H#T>SZDBfdY&Hg3dCH:6^E:<SO1XRK[EM],99FfGICS7/K<5EEg64/3^
^#2V>N^J0IE3BO^a+fL@C(D+HN:RNdIQ;Egf_EgP71&f+4R,LJFVK#V)TBG@67Ua
22JRQDO@(3bB:M.?b+b@0dFN;Q3a0R(F]_I_6P9HEBJP\8-_ZM/,/3VSbMU&\9\(
^KYB1E&REc33W)97=M5eY\QVaf4YLL,9D3>HT&IZ_FCKUR@N,b;+GUX;8.78LJAg
9GP0b?YaSe]910X03\K5]S6IJG6DUSLRP&KI4G]E[RACW<@6\cO9Gc8P#<7GfI/M
??2UQRVK,Y:I6<8NP4PP09\KQ8K,M:Sf4F=X+ce52(?CAP=VCBeJb]&dO&N0/U1X
=9#CJQ@QHB)06HT^F700HYS&]=M[W^J)O^a?7?3gBD0@MQ4ZgEJ01B+XN@BebJef
I>&,d(V7eW#ecfAUPKJ1OXDbDe6CBE5OVE8/.0P7]2P3g.BWO?V6A47KS6KSE>I\
OgR>AC-c##M(A&#JW&U7U)V(,_+KRIKP_#/W48:aR:K1B?cH]>D+)WS6(?J#fIB#
gX+OB\AX)V<MFVBO3,BIM(,(-ea/HS&PL7J\XOaW<-GcKaSF::A(=+8[6AXQQX0g
&A<<B+2dfDE7C/J8^_@?]^bH+I+c:Veg-7R;d0]&9XYGJ9KS,4@G26GQMJ2fE^C=
a?PCG0aGLI?8_QC+P.Z/5Ca)[>8g<(J:NP;W:Z8HTBc015.XAL+Lfg(7W@<I09cb
OEC\\/]:;d_>@<+KFIWNMY(#[5:7-TKI[)/YSfcJ/\7=IbD^Q?WecC9JW^Jag_:f
^dT@3HQdP>9/A^)4>Y]UV>G&9U8#^0eKRYWBU(e9@cfZHT\d-#RE6CXXa4N[=f\F
bT#&6^(T;0OOK<)0B^d_T\ECT>>D4:Tc7;XL[3BBL,JPbRUWb((c2:6^SX4I=HbV
ga#-;3R6MZS1R2DNQNFd/X_LYE)_ZU=)J^8GH[JCDZTTA([XF._1(.PL/d2_^LLT
):Yg4fE3:X^(c1MTJgdI^=E[RbeS_A0[PPQ83LYTeZM[A2,F?DVaUQHJ?dP@-0#:
^]aXZWBW7fb]J0^SU_^><4LPV96GMdKFU^MRY/)WW4?ZUg,O&3eSd<E9L_4GMa.-
X@,32LN#@I[,7F^FPPK+\_TcbKgF^I9]4ZC::8__;:]dELV=1T_Q[_\GFAC;1Qe4
IHfDdf0:XPa(<Vd:I]3<=OQ=b_4F(/YA5cSASOO+P))/<--f,--;AUaR>@DFR.G9
YJ5UCH50WUPW&e&J=cIa#L(WSMcV>[1HML^1PX8K9#DfS&81&&K+ILO&25=Ga?^)
CX3Je]3_]YG5AMcU_0Q+\7f[deBY7]cOSR3YP\X@0?4]B/#(<Z7WX>L59)X:LDFe
..C2@R)/6d-52DdSC#:R_=&&7NNcB[=c7HA>Z7;>VA^E1&08a8P65RVPeCN5#8<e
O8gHF6SWKAP0<:.0Kd[/Yc_8eOS<d=>2\._]MaE(G;^I@S(Y1geCCGC9IHZ.dMS1
\CD)4H@?V53+)\)ad]<(#31##Uf(EB.4U;N\-V]R;f>2=1T:adA\&4)[(B7FH^>g
KBYH++B-4X)g\1GMTLZVS?bBZ/S7d[FJE.R6bd=Y6+@R5]-gAEA@[W[T6<NU[-+K
(g@59Z_GH&#;GHOe@;B4<]:,Eb.4,,G#)eMcD^@:=Og<Y19cW#Mf:7e3:MVd[UG9
VU<Ng;H3]4_Y<3],1I/U@1<,J7&5IVQ)39:>&d^<+&U6\VcEegO<BBPC]GB)7;D=
,9IfC?6/^4;&[HWKY[UdA;>SZ^K6UWaOd0T:)FWXGL4VZ<D_K5:?,EgJPZE2?0VW
D83g+\53EQW^?L:UOJbF&_>0(3S2af/UeIa/b;N(CdM?^dR3+KUbUCe0,\2=9b]?
LEV1g3DBfF>eAJ_L8@Aa#:NCUD+1R>#g_M=d3Y6)B.Q1GEPA,UJ9bg0;;&Xe#I@W
<=(eG8d;@_PN\VbC.\a)EJPQ;=gQ,.P3U.Q.<UDM(#WXG1/ZM1A2dL?QP+7Y)c[7
40Z^Q[C2a501-4KT/D_JEWaV)UWI5[EO^cb&.Ge;O(A53Ic3>2==fE1_[)@g:_QP
A.;P^#e\7-9+>ZUe2J=O&[QVf^KO<2B&QaBA<_W.gAaZ-#D8RHL_L4FJ6;_B;Ga0
<QaE-F.P4\(+]Bc0S=]/\0?[F020D/BgH].2Z+Q.SW-X+3,DZ;>8X.K/..cG\:_+
:B>U_,>N#;P(MX.TU#d8?T(ZELaXR.SF[L1F[eCK1CGd?9_I91g#NH7E(P8XTJPg
A4TV/MXT2aIMF[KeA@EBM^<[+E1V>,OO<D=I/bHB&RaO6:T?BeP1M[Og/9U@dQO&
@)a0(YF8S_NU;,JZ6OC/R@ZJZH9f]Rb[8/WgVIFJO&31G3MJDa>baRXMRY>6#+:X
;4A,9>1X+K5T&P@-=G3QC,MIBPX^KGV<Lg49WB>b2e#=&YgaNcOB;@)V3d2?KX6.
fdIA&)G8b3FBfZ-.b3<C5<N3&agTM_^,Wb@PbHLB+H-KSJB[FebDag0ZIX,T+RN.
Q>^VL.PI0WCI1a:9D0#N#G)9F;TABd>R[.KYbKWaGPb9-B\=2:KL37Q\QBe;0?&0
WLd=LFGQ@7,[981\E<RZFg5<\.Z23]8b.5(-[]e>@Pf;JOf#/V^MR]TG^4a0K@0\
[^:F?4c7F-e9&6CT^,-Q^aP8RCW(#DeG;XXV5:&J9]gc>HR>YCK^\-J(9FL1KP7,
.Y70YPP:H?TG6GN>>@65Q1>f-1XHA02B[VV31#9AY(Z(&&4F+VCb5;UIXD;gY]QL
BI6,8;5S[CM;-/-HaO_d8XcdVF3I_e[X,H3W)6R;[,:IJ=^&e\d1Y7K1V[9;W1:K
5_Y<Z\FU)I@;>Q67c;-S@S=8HVV?]SN<P+XafAU+IMK8WLfPZc/R+G&DRRb:KVU;
>-J3/\ZS.]1>#dMD?/,1B6YF;CCLcXagG^fG^UP:#)K>NH)(dd]XPZET5=,AVL1@
57a4]F_6G6.5/0S=?Zeb0[gaZA3,PU923.4DaQ8+0+[>BPPRC71A&5N.K)B]5@Q.
LFeE=e\BO7&R]?)Jf^U4^[_NRXG5P+K_M<1S26(AKb^QGQ^:TJY73QQ4Xa^TRF,6
]U<3Ea^LJa<934K_1dHaIH?(U-e&^<VFJXD.3#4_8NYdW2@>>cdg&=:?#7LTDf-?
<-_GE5V#L4??,F+L&3>^&a<-S\,RH<):_>QOY7V4O<..MZ#+TA(5.Eb+VZ&.D=PA
G+&bdbF^)JP]_E;EN=#6I_g7;O,T3Q/a#B##U6KO__SKQ5,e4d:cQNOd<PPLH,1X
+\bWSL]Abb7;S;g8]eU^>gXABKJKXRf2FS)[O-^Q8.>]O4W&fM3T?e5)JN##.B[P
1[+Q+a)Z&)HIS[9_RZ/_?&5JKHLa<AWYJ1A;&N<\\1D;SPa;5NL6Je\[6-#;W&Z#
b1[-e+IE]-c&QJ02MaD0K#;:e\bD:9H1#T+4.R@E[2EQ2+D4+U0&DFc0=Da4(?DZ
^U3>dgUY;,CAA6=+S@DK_T6<09?LC9XR&\P;SFD.39534N:^F05XF(O/EJ^M]Q-(
1;MP;F);;0^V4RX7XP+-Q<?N9JJ,>:D5I]3fX18-_^,<=cN):4ZLN,Q]@HP-&@63
IK-Bc4POJe9_NUd7NVG.GGT>Nd47J.B/g44LTIaETF?GJLc\S#)Uf02d5QS>+-3d
Re=1B4KN[VE5cNV0:Na3_fUG.LPQ6D9PJT^:<1<-/>bQL5,#M])>AH/^=@^A2f4O
<FUG5HbKV:.W6<3U3M4]Cf;a)]?G7T=U2TO:bO4fK1b>bTaX99fC>;+Vd0:.U&6A
d8>FCOF?H24;ZD+/4JLgLZUN,9c#U[\73@<E&/eRdZ?)47\EOKQf\;5NC&A&;:<;
C73V]XA-.NZI.T0=4A&4Gf@+/<0a/0RRLabDSYT/#?fSJ9#a47JPIX2+A,;FK5/I
W3I>AG-49&Z.XXTUL/39J)ZT2/4^.H=BMR6MH.7H\[^/^W>KS#L08-P:.0O==9b<
)g=+fA,V8UZ&2bYX8=27O_.O>gFR^:5b\AV#[VJd<VfI#]6V];55V^Xa=d_WH45.
M\)P[)<BEI+VP\P2<.#eO+CF+1;+MMF-8SD;_#=B_0+E:ZaQMcIVe\Wd&Cg3eL[7
)<879HV?O?/1g)8McK9J=[XVa\=/.dYSUY#XCM@Q8,RA.]\=.OUZ1b-&fP03Y7O>
9E=fNbT&d<Gc,T0b(]/PL=)A1O5\KLfC>3BcS2+H3;IGbTd4cCZf3?3L7SKVU._#
Y#0+Y3>V.Vc.gE,5=2DYO7^SQ\+A@<7ca09;FU(0Df]bcS\e&ANM_P8Y>[GALH0g
U#VI92dDP<)0Zf[]MV6<;F.ZR7bK:,9+AaQ5Jf5<=;R+-a&/UgX)I)(P5/CZg_U>
2_+<d29Ad/Y/aggE2=2GPS,<-9agJCP:eV]Y_F7GVbUN29[,(]Q?#^O/S<VRV:OH
U:aT::HU@Y\Sb=+3aVB[]Qe;8GC\4N,063:>/:Ca2D(e)<3PDO^J&QZL=?c0Zd.Z
DXSRY-Y_)J\Z-X&A2NDMUd6@g@SaM1R\-<b5GJJeefBe9c2M:e0IEIYHFHLWTOP;
8P#b=ANJNPe+Ob]f[PdE]4WQSe11NZB79Z-,WVVTH2O7XH3AID_6?(YJ5I1#=IYN
baU8G8TP^N0/)AOK6=JY><2?IT2HeSbf:VP[@eX13)^bb6PgZ)g.:J&#I^@6Y+dA
,3+Y,N0C6bOfXdKYPMGIc)SH)-4[.X.JQ0d-9DWKZVV]LS:0Yg=D\/=b/9MN96.4
I0R\XG:16-:,>[3^0^#90_O7O@<e,;e206_9F;?<CMT^=YZM)=:OF8CW9F8=QE;\
ea3Zd128?/,TDa+]S\-:C3b>f>+6]5C2#U-a_9dd^E)U:b(#U)KD)U><+A_(N&:a
&>,OX77OX[08,c&[]&15Ca#PE1<;PAR/9>V34#2@/JK,eAdXE9>CCWGJ#;fP0\,&
T[_e6R/e.aU:GD7>aJIa+KFTaRT]2GbfJQAeQ:]b2L:^\CPdEaM1\c@69@@IW).c
4TGO8K6IGfe?5G9e+?1,_f7d23SFO]<JaX6C&0^.UU,=;Y&4fM?3A6d=0G21DXZe
S3?2JQPISb:ZI8^>YTWe&gK&KQ>AE;E9fH;1<(17VRM#-I6:(P&[+5654gT0^_fC
ZJG)PY>;+FOSZ<&e,+?U:@?bEB\6g=/:&]8U@<&JUeeTVK==IG(UBH(P\YF@;_34
dLL=eA1H;7aP=0VVcMWIIDMKe6@#,Of(fO4_&;,5JB&ET.7.0KMb_9Wc;RY-G^#H
1M/R?Zd/[_/Zg3(RM2P65NffWLF^LL91094(2f/Y7_:[a9BX>\]H.fP1.I,:?-OD
>..cH8.T.Q.YV#P&VW8^FTZ=O/@K.3<5+?YJIQ+8>S.V.d-S,)5?AT[O+V,Y-,F@
).P@=@C:]E3G7]fPSVYcICZI2Qg,78^H1H:R:-0<XKT+?ZC@\+#7f4=cT2S018M;
XeJ4)>:9gV>EX7?WgUeOE&W@/ZJ#(>[SLHCeP6V54\N+2KV/1^b+[=<A5=86&cWF
=9_Z/2/g11Q>7eH=54+M/RC_E@+1K(H^D6\Kc#?).#(-2YZef+F)O@XUL\41&/Mc
V+_?54CN+gIL(B(C^bfYFT0JOCa<;<K>X8>+c25]N+T2MZ_UA5T2@HQ-V^6EA1BN
OEP,d_F8DVT@@YTL[G@G+UB)PS_HE<[7?H&H\d3d[#VSSg^V+Aa_R,3#8ZSTBBLB
MIKY5LM\I\QM?bEAI]MM,P^^EcM+.)@Mf@[gTK^<VSGR2[8g)XNI38DPH1C2(HZ1
bS,GD2())\^V4R7(;/6H+.:<4VJ#bd^=6H9&P6>=D-I]O89>/YFHc\CGDW+PEePS
Ic9=g-WQ4X6(];[9CK+0Mg:J11JG;HeZ_2/JN@e7-+E=Y#cM6WL)S\C:J@O+2HSJ
D8_a<?.TH5E(+13W6d[<20bNTC_DaO)dg@dROY\850C]_:/N_@19IcNNfOa6?@Y6
9PT5ICa;R9+.=,f]]BHNV3G=Bg.G+A/5YB@\2V;=-3aEf_Zc--0U\IOH)KQ1HTDA
]+X^PATX)J2c7OJA6-FT+^7)T#EIAAK>)C0?QeG+f9HJK9ZX)7V_&YDV;T:QFW+b
]Qa[6O_0XA>0eAW]1]ZD,)KP4]Y(U629@bAK:C8>\Q)c3+6.R#JFP=A05C6<ICcY
&f/eL)MeOS#X.?.QKNOf]D80\U0/LeR5)0S5fH+FRaCPA,EUbET9A(gaBU(d(FfD
DTGeR\Y#U9[Q:;C,OS7;T=fbLB.PKeS96RCGa6f@0?f>92A<JZ\\A-P<IXX?IH4)
4gS;Dc0G_a0:3[VRK:Y_-9\_X9\5eJ7a@6cK<8IL^F_IZg396@GZ7/#f(Z3YF_8N
:a?30MV14NL6TcSE>Ge5?>8cU7d65A=4L;Q>@1C+G+;N;O=#.d9OZ_=,/BF_2<)J
T7C^-7G<(&>.X483CeSH@Y&M_L,I-.#703dF:>#L.<]#,fW9_^@^db/\7NdN1=.#
6</5>(HH\NNS5a^\SBZ2Q;6.aXf(I@DH4:2J2#(\RNNE&d#\A/#]g]Y>9RCLU1J1
MSKM_?.YOd(J#@#N08XU?KbA/4:_HRSL<K,[V7#38bPEEHb_.B76Y@EF5)<Sf\WP
+Y_BV:bEL^4;RU@..J.SFCc:RHU09QBU>\W9EQ3(JZ6RBJ;@@OV]FE=7deMT#7dG
#7ZTUX3.NgVeVMa#R\YGTd4E^&fIAIWA8N(AT(S:0c&-]dN,Q\HBM.9F=LcUf^F=
dNWdY&.c1?,A;IaVd7@3OQZI;#Ge_31>DD6)-E:=:02)b,B1a>JEDR)B+\eP&-Mb
D4T)OI:X(T+c=[(^\,D,CT70T6a;5N,.(P]06#07#\#650Td=L#Qa#RIC3S[AC-(
eee-B?9YZ1Yf?^\8c6]_cKC]67;HPOQMV6PRHaS^d=^TS:D4^9YRc7K]2c9K@Q3(
SU>TK#Y(=+De=)40cV/QaPF<)_#>:J[5W^,WJRVdHK.XVHF6eHAAL\0\)TIF<D8Y
QY,:YU?K\ZW,KLDYG?.I#9[,\OL[0&&VIK;E>Db=^A4;B/>=ee;^=dU+9f&==1H+
XQfS#U&F:4+PKS]A<QZJf#ZXR()=JP=HG2B^]:fBE+HU),f/14Be(W4YefP\&P?V
Xd92)Y0F[fDaY8D@J\g0H&E\GGfVYHXNV5b\AN=,NE=UbM8T;7#+R,8RcR37YRJ-
3W,4U>]]e(eX0E&@3XL]1H1@4^8SJW]?:D(4.=XSE@3/IR;XK1M#T_gXO#?-TN3W
I>U/DeV.8U6RT]SK>LY6(Dd/O[;[P^9-)^JWB.(H@)Q^YD0O6C^?]DWYFJcP)7U9
(>Y?WD(aM:?8<U6E#K,UT,JRb,EL^A2Ka^T,R5Y+3?8\O[d?Q]0J_G]8/3SgCJ_<
\V3#ES2]Pb&6NY1U2\I\8FN@aaBYKe=9VZ6HXW@(2U&XN6-<G?B6+)?^77S^\=9e
?\e@GC/H/Xd([S+dW0R83R/RR5]5JX=LSU)R6)=-E?<\21_)WGZ+E9KU[>MM(ee5
R(W55:>:@,+ONQ^S\1HYNS@VHWM#_)3-;)Icb&Zc_0@^=8bPg.H,X(c2,XbU1S(I
eUgLKK-:>:Pe9_RBH[[H^KFa1GA_BKD.C#TVW7b.QD@^K,@;-0FA^3?Bf=UGfSFX
2/,\IVQB9U;LC(2W[OK)UD=H6JE:R.J5A=&b6NNOH4N=>@Lc]0UWB9Y\=HAQDF3,
b9;X;.6gYg5VXMfJ2F?STPQ+-TZ:A1_A\E<-PeLa+R43,NARN.Y_X6GTDAS>/PJA
9/XO@S1H,1LOSIP<(E]&R(\\e<K1][RJYN_B#P)[f,+NXCB.S#I]XZ[7YYb)VOR[
fBGU=@aO2f^\S_Q6f>0\Bc>=Yf#:^0Z;4aG\M7-S^8?W#ARR&,L:JHTHX2,N6Z]f
HT^_@IT5LDA8_MCY9.1D(RBSEA421(;XO\^;ZP>YaVXVC[>f&,MQ]JY/F<XDRMKO
>G1S,)1,?L?I-QbUP2C_c?J[M;_#G;;#Kf)4@6\1@gc((39;G0(-cCC_:GY,(9L)
5B=)97CTS4IR>;VPZ;UXQ5S(@U-KLLeBT;X+.X/G&1R)d(/gWeG6ZTQA9_7AG2DY
78T#J#TV@D@_bR7ZI.07<W,[UW+UOO^OE-R(H7GV?<TBCR0A&M]Wf_1R&;0JVc9Q
PTDe:^E\OVE6&RZI18XO&MO<gGQMJ^IUGKV[\=O9:L@/JD(c/IPVX^OX+H/f]/De
?GBS)X\3BWJ(OdU_<[]dDTQ6#g3=Z;JQ5g>YfU<UNfg+/0/=4b58]LB0KeR[3PL(
>=OV_AY<gZBeXSZPcVfGaLV)]HQUfC0e^I39L8Nc+(5Vd(aD4GY]?].&B)Z(J>g;
TQW0\1@]0>N?5TKG;;6DSd/^0<e44d<g0(E@#W@Pd+FLRKEGE+EM/G;U;(J2@WK)
14;IH@c_[aGNT>HfB_^=5e6GDD(]dMBYC09L4.SO0;=^23LD<->4g0bQe-QI2MEB
05WR21;2Wb)c7H2(7#HFObG0FDJ&]Q^R/?2W/GT3.S?X(S.a9U=UbV\GL\=-[dK^
P<.cJ]O,O6#N)AZD164[ZQ=H<3eGIU/9&]GPFZ@JPFH;V#TKA41\YUPQ8d1bc>UL
KT2(WOa,QE&ZMeJ4()8:C,1#HK6X+M:8aMI0+&\IZ^4VHS+P)+:<?:dBPb8BGPL1
B.FN>fA/1\RMY_5#.SZ2JA/8(.^&9;,WEKQ9\2Bea#?GXXFLfT:dVL@VR:LO=7I+
4\[:JS>]/?7U&4L6R994ZWceI+Q@=MA7\4addHa(^?N17Y2TaR6H@9-U.M4EE@86
9Hb^_6aQJVg&HbDdR1=Z4;3E,:_Y6/R=^IfWg5H0/T/O&g@AXDf\/X[K45^L(RN(
VUUR]+<B.?:\;>_^/\;-6ad;&,(+DPDM9-&SXce>I1]3a/cY_&TB?BZ8Cc4\Z3b>
)C\N(V1P+bcI4gVWB>HWX]47S,G?Q<R&YWC<YcJOCVF7<YR9JA/>28I4>F8.U=18
H4X(\bYI^[A?<cTgW:CEJ36a^d.L74SJaa?ZOB:_eTROW7Q3g]#HeTA=U<VfFY@7
gCF\dZHGR,H.A>)a>\B[A9/E5.3V+4GDE(5<R#;daaDe9,(U;^O,5XDTTQ,6M-<_
EIZF;VK;NY>?5QH7AU58Aa4b=K4>?&ZK63T^3TQ>5(9;NaVg;dEeD,b,R\@:dg;0
.Q6e]>BFbK=(?Q^2R]KeP._QQ?P=,I./ETaD3@28HNHJc,8cQUM>^=C01W/77b(C
^Fc);^a&]:QUd==I8E=QG/V_34aUD#<Ve(Hg2+Ye204Y13^&<[LcK8Obd9I5;:.@
V26SP[;BDYRW14/B/CLZH0TA/QK=HHU#98Ic[Uf2U&C#0]]LHNQG:EJJ_QBUWKb6
bXSMD:WB/?Ne[,GYf1G&+TJDfRd=_+I2-+4FbHD:K(+@f:Gd\S8@5,7S0PQBad/<
&QR&VLd8W:N\:4.-(TVNYe8?0;3AD0ZgZ:/A2cURCAT#F^fRL)LY_Y2[?e]P#TM-
<Z58eI=3+\@;40/^/Fd,06HK_FEPX#7^;X<:b=EbP5R_1e1/-G^e3X4d^NX853\c
#aU_67G)U??LA=?&(PC\YB-Le;7Vb92&C.FP67C?.,9EX,-,@7?7-D-:NJeD)K_A
Q>5(83>f0W7S(W:L@OfgIb+4e3C(e<a./6=D^?2bf+]7b=gRE]=aGd\gB@ba^28H
F&b]cMIKc&dQb8N?T?)d&LK-F2A:c+;\^SNgY@dL_6fQ7HG6AWZ</RSXG\_L9,4G
dEGYB41VWAc;aA-Z@DP&)C</:^.K8f;+4eB()H,aNB:2?+H+0L-P)PBEb9=CSBB)
ZSL1KTFaDfHC=;]W)(/GZ+L.Z.)X5_/4H6D?3.P-L3559?->b#ZB1I3<TYg:>P^f
ZEg@[1f>?JG&aOG&:TY_V8FDHBZ>/Z-=cQ#d_#<4^9PWPE],Z=EXBU5DbZEH^fB8
31\+PJ(2-\>BI4@<fcGRR-<UUbaa1WA_8S20a1IJRIV7Ic6fFOUebHGZ8R]PbM+Y
XJaOAK]aA\e:94-QM1\-;[\V95]JabZ)e@/_RADW4?BI0ZBNO@/G.D2HT#Eb_-OK
XZBE/+25?98;O2Z_a(B&M/?5b,83fG74,(gL=].GO]c;g:9M16GH7c8eY.V8g9U(
;cad=aEXI[=\M,;][=336S6Jb;/>bDL\?cJa]Tg)d#)@E5\;FIgLJ3g,2W_XH>g]
SFJKa;>6U=>-b4ZOD;Qd)Z=@Kc(S6bYW(5_=/NW@<E9R:\)gSIE(\g+U=?PG&-T]
).U-2<D28+D:>g&TQJB;PJ43(];<Q<Q(0BZPO4M;A4ZAfM#+LO[-PD#R]e=-?NY_
_?T_cO&CADZV2c&e9fdDUC83R+eEW9<+?2JbCO0La1B#M=A:GWfWZ^\#T^\T:.O1
A]/]8H\[J34P1DdE[F6UHA\+\)N?<\ba1=T;>6.6?7V&1?+-M9729S6#JHLT6b63
@Z,CJ:[LG3&]DI6g=W[cfI\XF=@MI=Q)&8:.b^<Ng6WOGL:O_eZK>f@_ff,aBM&;
YIX0I<CT#2-=Ra+e;Z_^<PJ6a/[;56AK7RQNMbH\4[f=;6:c:V>C;dMR;LC#L+IH
b6;X_?RI4VV1ZR_F<7P@CH]O^M7J/6R?J86R>_JOfd:N8+.DQBe1PGMF&dOELK.(
<)0De&TOU/,1F@?5/:dE0WZD]CR6\Y(X:AX(BU[(eI/>/Oea24?RbQ9X<L8cDbY:
BPE6aYQJeC?eVL?bc1O/:5M885R;=^ORK#T_^V(0QGPFNMV[621&G8BS?2Nc143@
K@b4Od:4=:L3<&[YD=.1VH2(T_OXLVSGV7EAETS9LU^MP&C2]cGX<CFPUcUB4d<=
VKXQHVQNG\c/]L9cV<,Yf7STc-U>2:+0a(;<NW/-.[Ed6X]eGBBA0#/1H)#2#L=O
Z?DcWMIX-R=f:NLeX^U2LaJS)b(aQaCVY^d@^UM2B,L:Q>KY-HgAZ,EX^.c/T#QL
&a(_XdMbQ3/0Y^-W#F.V-Z-+b^VA?Q,.89YIBFGWYE)e4GO>U1G/0-B\DHGEUDa:
#);QRa&<1\&9)7JR3a1ca[Dd:C[3@EJc9],XEf.^]A,e6S(de#G<e[K+RB+1SRcE
1Q7RN@3+<J5RZ+Ja+S<TRV>,;O);@ZS&&+a9]3Z[T=S[eYCT__0I.:>B5,-,^RB\
dAaNT/65CNE/]LBJ8ZN]R;g)gg3-R=\e-48>RQFJB^LZMWM2A6(d<85=0-g;5-.K
=M(@]2(3]\F&(8gc4S5cO+/>NaI3+:<bT00_B1b3VL24/ZVf,8#O,;:DOW]c-S>7
I+8=YO]D8.PUTT.@cR6O_;\:\E?#=W:<eI7;I=/8&P5.a]b)+?YMYQ5WcR05^YDI
Ec5=8:Z?AIB)P9INU?JJ@)..eg0?U48:=;6J1CC_X=/_E(T2X98Vg]QFF]MS;0S]
IaAegV=P?[0LHPfCN-;ab/f)_WQXR]G37d.L8Y(VScgddL<0:)/9[[WD2?CXKg^R
Xbf86a,IaE+;XL+<>=9TKcWYTP,G6+\[Fb1f82M_B@MTY:9TH[A^8C@B/_93U?_]
WG27(D?F1@OcdOZ,J@EL@PM(0^6b,(F+fgVe4_4<HcY/E-1&?KA7LRAQOfF10A@V
MEK[?aX#&4cX-D,\A6IV0NES1U#[aZ0e-e;^&SM9KdB7+39DHU(HTK(,a5(IQCX-
H/218f6,>#J8[a&YS_I4;3.[Vf?IQ\O7[Mc]J@E<3C,H776a;]I+6YcQ^KT:WLS.
Z-[b+A:SC&&(09g&X;QQEOG+G/H6Z]I4IR=dc<3,<;XD/A.SB,8W#c_RA:7QfT5B
.gabVV+R61XXMQW1a<8G,[CUVXF+T-719E3:_C;M/?VMEBSP^3Q##S-Z<R<ZaE/N
-&BP-bYRWZ98dC/FS4P5a&(<2M^36KRRRL<O42X(Ya^&Me<4EP\2G+aX?PZ(Oe??
FbO4A2)S)bN]VaVVAAWF=&)dZ7Wag@YV<+7;?O(5R/KCTUW5:0XBKa9eefR9:4f-
dAAO_27-.F7M;=6W<29V1CH0/J4<^7,OHYK4XE_DN\<C;Z_NRbCBd>.GH?SAf-c_
-,X)O,DDBHH14Z#1<+ZX@;FSG5UZ01NT)\ag12/PB5ZXVU.DI.b/Y:?:,Ne>/]94
E07SbN@^.fU,^-_LJ^/.Ia5GZHG]49Z@/>:#(K#B@CIWWLcZ+5BL8B=68=[^<gB9
YPFZC@KOg_Y[dRA<]\\HZOVA>Z<Pb,]IG&aF:9<C[&1<SNB(C><PP(G/;+S>+<aS
SO>ZXC)b&)A(:.BS(a)X?0g2JHS=E<OT39H:48f^gI^TI[L-MFMg)8UJ&LIIB[&&
>4U2ec[Y#bF1,eO5eJPOEHCMB62;QLVCcL5a&gZQD?F8+B7Jga2MW,YBQ)+F0AbN
+,.T200.#f[TWXJM3ZSLH^e:GA<ID:-O,U13d<?>-3^;_[.:E&G]MH?=PW\@GV4<
fC@,MaGCX4IDC3(JSF+;V(;9gAGg<?PX).S2BN_=FXP,]_CDV3@9P.AXZ(KaI4A9
WM.2=BNQ^GW-Z3#CR\+^BcY#UK^)Q>DLV6gEIV>[eD\E=-#@.XWcA31MPV72-A8O
G@D5&K&+DW))/\,N5A=/e4\V@HOIg<UZX8]7Y1(S]G(@\be1YO(-KQ7<NH;(Z2Xc
7Qc#NZXGf++8LHKNS@CEWfO7^.3@K33X,^87/A;[PML6dG<-OT&AWHbF5H13+3XD
=9:bDa?;1?Y@BP:QJ8Q1H6/XZ37(.@:.LD^8[?31>4L96(b-L-G7:DT[f?L1;E4K
5::1VQU^EAC=8M27_A?L#Ug@34(5>L90?E.5A/9V3d?c]QIe^?>:bW@4SXD?X:;X
9;.JA<PcTDPc^7cQG-/^OLVU8?+W>)cSOd>;#WCAL7;YQ..FeeQf_F/P:-),V6&L
C^&@E]5(8gR9SS&+bTb6XcE);eL(Sa4deQ,&gIO[6<330^SLH;HaC_>5e61_7:/^
O&FZ4a(XaY@Q]D@Ld+gU4=O=#=LPPG/T;UK<-3+SB+:W/ddWX+=9,^GV=TB75SN.
I]:\]?7I)5L4\e?De+OD[VCAL4=IO^[X_^=\JSN[_a#UM6G]Ta\:/D2FCDdCB+L2
<VY?Y\--WI_O/aM+FA78?6E_K]Z<(Meaf(187[O&20W43LfDS_57KKQaP7><V7IX
AK5F[\TC8-dfL2DXKD+KB=+MdaXfRP.eQ##aIH0G(4EUV,L1X6>AcEXP&AeE(W(g
R[ee95=9375Kb14&+:A]SK^GC,<#B>GRBSX/(#;KD/CUFQ&S0a>b0>e0[e0fT@88
f1TK;TbAI_YK]3YC6Ue@e5@F@U)b5^@:,LC4cT2fGEg_80=5,?ZY&MDENdFbDB15
/7&Y^-8#f+&7AV\YYc:<_/B-Z;YTeBEFZaRK#6<E/E&AJ)&1=:>&Y2P<c2^^5K&B
4-YB<eME4=XU1eff]PaO1[I((Q7Q@7115#V=+Lgg@\?cX33#<gb?5-\dZUEO8:QO
<cLG+V2<eB)Ug(Mf48Jf#GY<gfL7+L=&De-]N76d>TeU:@WIg)<N>EK-Zf>5LV8J
P539;#5b8Y?UIfZH+)\U?WPKPS-+\-U.YKK&@.f61-,ZU,:2O;e2</1DP,fd6Hfb
&N)+U27;U8R[^6aTc?M4NB):>\_)/Wf12ZM&?[1Ua/RVL1@WGO1V/Gf:fI#0XH02
(5/(ZK/]3K;ML&)#A.<bPVa8LV]2T@+PAOO7N2dSf-Z^(aICKe8WQA;?]PKS5f4b
-;>DJ4_V@Q]XXZM2^TFP]d7M8ACV:a8:&/.P[M-F5;DBNRQD=I9HLV1DJJNK5].e
++V<?,7(OP);eGWUW@:E/KWCdb1XeQW>+;R712^A3eQcS3B.O#^\Z[\XSO_EH#5\
_fV:S=ZKI9T;6c:5;@OU3^[c=-8N3GIN#,ZQ^7GTLPH?R:/g+AE^QM77N;Ye0\SD
RS>8=4>.P9F,FG)LTQ\]4+1=Q#C:Z:5I.7.R-Z.D^5B>(X-V;E3+FWXQ^c^@5N20
[)A#&cXg#T.7\=?M7[59+X.W?=?3SG>&P/WD2KM,Q?(ORD]:HA>R-4GH:#DFM).d
HN_,#.N&BH6W1<RGAW[a-?X<]\DE-8Aa>C8[T;,GZPEaO&.&3\NQ7JceX8W;1N\1
TfgT44cN\g/.f=Y4/U@L?XPWT_SP?Ia@F#W[?IQP.S3R_MCD6c5))S.1&E)N?[eX
,0(:)-A8\XfdF1c&L@_R/YQ@Le-DI_ef??O4+2X^IGPO?HeB>e?0?,7>fNJbeS,G
F3C2B:dMT+;eY?,-#(,JGddf[b2R@TR=)\EB[1PV>f^\RCGIeWH<(W9,&;RSF>]]
C:f^8Ce^Z26gUGV;2NBL_a_+RM1g/;R\bH?U7T+g](F[R@5cY^01UP8H6[1ZUD_M
KKUM?@bG.IL>c+8633UR+CHCf&<LJI_eD8,)AMZ2e&]/FD#3,Q>2Vb5@I6;ZYJWJ
aLNe4KV<a>+&0OIMW<_#W3ZKIYQKTTM5.^.E[[d((/5_=,Ia:a69S(?)35\:3?BH
9.XfN@a85W?L31D4AOD(aKBSNC/)[;?HMf9#f7[1/TZ;7R)Zd9_T.g3TAORAU,T.
Q\QS2fFg^KS/[2DA<#->@84I;gKRXDLTc6F/a0[X+dROaW^=]Tgg@HA1XHD&NTa\
]CaRU[C)V#FJ3cJO@&T52A4^dbd=W2?@2)::Le<]YM;/AcG1<S5LL(NebeB?cVee
a=?L7ce^]1++OX,#9OC\Q]57@4^VB<&N67B9@@\DG_KV5<G-dUNL\22Na6J71;,K
N_DEMP#H66?IL&Ie?-X#.=4c)0WN4a6HE;FD6A,2Z^AKg4H4D=4UN))?HM@QZV&Z
Uag[\T,^3:_H(bD)JHBY)JVcceO_[2g9,^DWa_,7-f#AP9a\2&H@WIX(Ne7PSGB2
_e,D2Z_1U6>:BRWU4;8)P3\RaTKIF&GXMUd6NIX-ae.&\MNdS10aN^BF=5,?>cZI
eU+f8F\U+_GHAJDU_ebO.29Y]g;[/#6:)4gMCR/&.YdbdF:QKDZK:/Z0V=@\cA_H
WO0QJCN+:W/=e=:U^CFXHC+G=fe-F<1J&B^DK]65W^B;.&I35@BE);>fUR+-SIRb
3)Ia9QGZ744e#A@#F:._60(?>?Z()W)ON&HRLEL:)38g58Z<2V59BgH;0gYbX_F[
+,b@.[C([Y&GUD+J;<GSVXPW&>Y/RRJJ>4V/WeV#VUS3Z&Q^8Jac7KV-G7DLXU>D
_X)&7RID18Qg#-QPA.1Z]7IT/?B)<XLedEc&\0:,FT3H)<N<OG.#+7,,f_;=(FKR
S6N7bLO+7/WBSIB4eCE+GN;ZMaG-B;YF(@3dM)Q:4W)aA=N-\eAaVBD0bWbS=K<9
K-;d52e\@E0BK37e9.&.W[IU)6dAAET3RKT,\)Le(g=[bR<3bSRB2QWDa&G=&/+E
Z^3RIMOM-VU>Tb)#S.7]3E&f2;=9O\:VODJbYCTAB+BN;,@OD95#^:EgJWSJS94J
VUWFRQ1bc\>UO3H)aVM\GJ??XNOK1gGFW\XIcf<Q]^bI/K-M9RcQCV@5@.WX7-@:
M4)g9f5,Q7Y->fV205F=\5?8Ba?MU;6)]fN_c.Z92;L(c6aLe8^7S?7>J/F1RFMS
_&XXgQC&N4IE^K<<HXK/L>)SR\67#H:K5=_@f/5));ULZ[+BPG?HS).W(^;D4CcD
G0A<e:cAG)NdV8da+.TCa>3B1QHfQN?d([]#R>U5:_CXX7;-:F5)cMZ2.989BTJT
(PK@/F]EJ>1VGJfe\5O\[SH]A(688bKeM;SY3eIA:/dVAKc,1]7;WS&T3_NH==FF
10cBFK<9+=_e)V:8@N&Tb)3EYB.fCD/\M@F7X/G(9>52IgReBW^8Y&aK,G,/8#.#
/DV.STC.I4SB[MNU>L/_WKYe=HN&SZ\5I_d)M+8RLW/UZQ@N\\K8Y]f.\YJS9ZF#
@a=3=RZG&_d6:b.18I+Pf5VB2DdEX85NOI0KL6U^VLI]LJgKe>;PbXNHL1L/MZ(D
Q1IT(G2CA?3A@](5&S6.-R_+ZUYT/#:4.QQX9fJ?F2-J8LG.H:G8_-7:LP0e9aQ.
^WS3WSY5J_Q(-3E@I>PC)H-D\CFG+@>90LG8>5KB-dDP,-cfHVJ\8@C</d2XA<f-
I;(NbLc@A4dLFQ>5b&UcN?+C9L/E1MXa-]c5]TW4eYDS8U>)F+:B;Aa#ZgKIBI\0
5HK)g]XVA[Nda>JY..4+e@KXd7.2XHFDE[,PL^SJN1bRZ4-PYQ,Y+;AbVU74>VfT
W3ALY&CL9T@D:-AM]G3^X,X^C<FFO-D\Z4/4:g:.XQ/e<g0]D<CAN-R2?582L1G=
\6>gNIK]NL(g9Zg/Yc>@agHJ,U<,ZLK:K0b#H6EgW,5J7BU?8;c7NA8.f?G>AGJM
794B@PY-(T<bMK:gbU1XP8[U9-U[R/,9b7?(-_MfMR[6dGM0+Q>M[B#[Y)-2=V:;
OUcC?d1EGWV>gL8KU3FS93QbSQ3WH@TV?a8A/1cHODNgN?5&JWQc#LC#=L,SadEW
c8-#QgJIOZa+=AY26F.L=6@?#7=N\N7c?845?3&JM7=K.#OX\b&NWK(AB_<J7KEF
847QUb(QKXEA).)7\)g9;@).F:X>[fB.<QK7;@cD<EJ(L\0PQB15M3PRNMT_+9Xd
fY9U>;cK(^?[SN3cJNFE\7MQ&@JYg9b];7;Zc@@L@1)7(6f.\T&0\@bK<P<)H92>
W]XPf_TO8EeL]+X+7c1-TS9W=>WZFP=;]:Q@#\)LNC&@_5I_(9gb5W[\B_5ee6<e
e\8c[H+GYLLJQ7dL,K78IO+2Y+bEH7H)b(PM[6K\\T#Ud8K\c_=)8[Y3SJ;65,cP
90.94&a\:V?#,22WHC<450_96?cf[2I)/2<0_W^<6bF-[#^R3.R:B1)5LX5E\&\2
7S1CJ-NB>C[L[L9,8#NT1<UOK<Q(@V-H,aG8DBZJ9cG=P,CRS6BJ\Q3@4WE-+)@K
A\?g2CV0F7XY-_MW#9f9J5&BP3Id5VQM,(O^]Z1(.P+cg0d[2;AZ4IFX;90g81/@
g+H5QMX\@5Y]Z6OJIVSe@dY].B&e&R/4&2fQAd.+,+9H3d0H3\1.dD9<Z+6CLG_L
TX7\D&^9S^4DLSWQK2(-#=:;#/_D2/Z<G#MHEZXXZGD;A4H&JfE^N[_<]N4f=\H/
5PBb5F3<ZB2D_R0EAL#4361?Q+L]\fDUg(,\F12R3Y>8IQ>T[1-[CK8BQCA>d6>0
aMO[)N?>73NG,L,fDHSb7C]P2(VB0\[d]ORd?7=;F+MP>/Za:APcO:1N6/5&ZTG@
85;C5VUbB8.eLBdLNJ9Z6Re;9+K&V0AARG7d;eT.b6dJ_fQ46aXK;Na+2F2GU3HI
L:1c\G.QNK7/LcU159MF8<<7f5#OJV=gb_3T_SZOBb>NN^A?YY6N/TUY+KK2<Ma&
A74fI+:FP;Q_GEM+,a7aa_PQW6D]A^9#^]DL)(AG&0R&RX1(X[8dU5edUZ#@WgVZ
?8P/ce[a.S<#\/JDS,c-agRX,Ia\SZ,0HFXI&R253_&P=d&9@2IHO6@5:5aLD-<W
])<^JB.)+@;<2V)f^FgbagBMQLAeSLS9MgaW<\\?UgMXR7Bb1:?c>(;P&=F2):V0
#34O@Q1:/8@6]92(E-78Q2&.,fAI^M9=Ca^/XU6WU#Y]OagHP5GbR]BXB1@(cV,5
?N+aI4Z-_8MSV==VR3[Z7V[9:4>a.?HIg3D<0R./1@c>,Gf4;;?GPL[P\J>7GIKM
abX-M#dP)4Tc)12+W0(A_GT>-_ZbS9/?@7NJ8SQ4R><9/EMZ)T3QVA3DNB^CUTL^
O::[5f@9gLFGWPa;R70T5JT^6?d;PgU_SgUg?f3X8S;42J.-d,;QDK6=Y++)M;ON
60;)@^EDY8;>YHVHB&FJG@d:EgAY7&RbEOaWAgQd(T-6IICQf=N4\FB-eb+3dOcd
AKY,3b7-0.PE&/W_/c2GF#&gYbd>Nd7=HL:CB/3J?ac&U=\M6YTHdGTFF04\JUfb
=E6F>;Ab.c1FPX+da2cS&Xg<JLJ.]5GIOJ9U)UZMTJVHC080CEPF]dE;4#1T0Y#\
IG_BLd;M2U-HQg]U/R\8(;?_)+/PFa4bF?@DQA;4@AS]@5T0HH2e([fdE\bS4-b@
8a.A,f[[PKU=6Q.@dI?a&eX&a4[265\8NWFOUe7BE0FQPP]&JTW=2WdSQ<U9E<R4
5:ac^Be-.1X7;M_E[0&TTJB?)gQPX=WaDQKL:?=,45H9?.=,Z3VcV\I\G&J5--OG
,,0(,R0YB_2S=dY:YZDOK\(/gL5Cb6Cf-8d3M2IW;SF+[\_Y@#;_9D-8;7d@B-SS
.GgJ=DA?ff(E>2QTZNDbd5477THCGVdN]5f>=B\XJUVgHL[?F6BVL9=CKU>F0DD=
:1eB#R-KL13&;>P<b43BX6;ggAc8gL?T:HWB\S<0R=dBG>[H3aUP-dc+Lb@:WVO9
_NT+<Ya[^3=PUFAYZQac(B4(Z>P_1,>MN/7@RQ/?-dMUN2<[3-UJ9,VA\L,44BLZ
C2<a;Y--KC<TD-Ee]:SZbX3;]=G0VNe9gJN?8g@SOH3D_AQHL15S(HF\R9&LZ1A5
1c/Ka6558E-\Ef/&8\O&M4_0.c>&<CX_[TD)ecWY:,VH5^Pd_FU?^3,7=94Ag)>U
]T?[fRbU9D@YYS7^A_bV)XQ:>3/?TWI\\YSV(:0TNCET1;?;RdCUCb=a\>8,:1f+
4\f0Kcgd0fV^<)]AK;<N)UYT;H=,35-6@.f-b#&LQVcS._Qb\^C;^<XQ7N\+,((^
R95J(P<#A\JEL,7G/PdJaIeg8(SZ6gbQX3b:@[\c1+ILSKGSR+R>QL1RX/,X>LgZ
DdVEd&<=N1]/R/T<(YV]Cd36B0(-_VH-SfaZ35C0EJeX03T0aTU467gdUeXd8NH<
\236=5O<,IVFMKUX19d+R0,cNSS.N:V-/bNWbSN5D_F+(AA.@YH3g99Dg7^)HbG;
IRa,Z8XJFb24K4A/8PVVWA3Y.<5dICUCG]689DEQ.5?0cN3UY[MNQ<(]@<V1ZTfe
FbOWeb7W[^0A[aYL@aX&^/W7NB5QCIG/NB,@ZP=g4BI1CNJ)_B(/Z.c\^(N+3-G6
I5.XC0)]+Kd/cV=ABP(C?AF9V1)7bQFU)IZ@:?YAFFJ5ODf<JXION;@GH-&g\dZ:
&-,>D8)S-\FYPe]Gf(H8gAB9T8V_[9_&:GZ<(Ab:/5(,aI-#G>>)<M\c=eeK:HVH
GV8786LO#FPO?V=0TET][gf0ZeLX61.\2_FS=^C):EH.#dFUUa.cRB)301gDSKdS
Fd#5W+C4g>(XG-88f^]e3U/?6H9.c-<\NN<YX?K3(#NIU=d[;<ZD)([4<:fSf7#C
Gc?7aR[?a)^61=\\GS1Lg-E/eZec4Z9f@:1KV[e9cT27b;bIMbF6TW\GYW\^JSF/
+\JIfF22c)<Wa;1acGfBMcEW6P.I/=1=&I>BD1KHg?#]>H^X-6LV]-a,#LJf8EE@
M2.]3BJ#^=MdQ=A10[6aN[23WFe9Tc2(QA2)=C@GX3]1eIWKYP93C>gHR[(29f]9
U@UX])J5;4G3ad]L]baNIZ/[aGc_.LeBFNUA-S[Ff@DHb(,:1-c>XO@1Xd1QFAYY
D7-JJTE56NbCV.<>UW&fOR]JAFN/UB9ZNO\GX5HQHYJ6caL21^1Rf_A.9\9/>RM_
Q8N</H.VM,J/eY29GXF,:,8;g_@2&N9Yb)9^gG_3_8GWK+Z[UI=MLDH+-SK>9]a?
&HCW8[BE7;dS),:[=;>b?gd/B)J0H9?UX,V6Q<YfBDa[-CO2^60=4,D8T[BY]@SH
_-/]C&>673_;IcJDA?4&eEW-b^E/WIA>2_^(\fd/fDEV5?K46:A01OYH>;1U>IU9
cXcCOROJ)>]LC_WI#XE<JgGAFg/)U8>V)&Y3#bGL/EVHD^=Y@<:5JIL3(gV2-@;E
)E3W-2)C9DPO(CU_V.N82B?];J,OPA+dX_A^GLc0b8(=g2M8-1,bF/HM/S4N[-a7
LC<?U9a[&(PB[BFR1PE&E,C:9.#U9a./?KD&XIZ/6&X3W>LB]-?,aH4R_Q)8D&B[
BKQPS2]98Xe5U@/aU77)A06JGd)fB\B>8<YRJ(3c?C1B4.@P6\g<4\UWf@:@&2:<
\A,_-]14H03aEDCO0#0?RBP_O3A0aQL_(M1SAJDMNKQ[YC:\YSFM0f[SfO]H))OJ
^0+(K4X6+LX+HgP[P.=CS[L.4V^VIbX6/PSQC_TIDOf9MF:5G,8@Z1I9eB)NN2aO
^9=<(\2WE:[-0<E)E,:f1#G\+fceHf2F.F-98<[I-ZK8D8Q0a9AZ_XZB\+@<Ed@\
LALPM>Z0EH#AT@FgAHDfWV=DPe(\W8J=6H)OTW_FVBPbY&64:W&S6LR-SAfT2f]\
;+T^D8d32;M4gR.OW5X,BBZ]2YYgOg[;C,FY(X6VS=SRMC1PJL(>]).AOG/8(4IO
\QZ9_:\=331W/P65ME7g>8d=]X/e&NMg@RHaF]YCdQ<&1>9_HS:5,7bNbN]@0#ZF
86QM&VQa?&NZ9a#+3)9)3X<P8f5F&Sdc(2Qbf_^OY5\02@X^@<^Y;5B6WZ=Y?b:d
(;cDF-9/[7)\dFU5cOdgY[,e9@KOg,]P4_8FY-<T;-#KD,C<SE;0S:;[Na:)6J3,
0VY2Hea_(PM6SVd5a3Q=)8SCV5]K:(=?fRTYS):GQ./8;<;Tc3M3MD8c2[TH&aC\
NQD51FC)NP#,bZ_0,\E4?DI,IB<Oe;K<PULOB9W=gD&UXdYEM(HKY<E2M^+>@)4)
-[R+8V@\L@8gS8fXAfU(\aB9E0\a=.\W-FG@W3\^5g2\P.Rc<?15DMUJ1QKf9N.D
g(=ZbbXHM3J5-:4.Jb\Q&7L7IK>ZL#==4G(MZXb7&^+J1>@)=U.PS9OA_6Q6.0?C
f[->,AY3b/+RHEO&Wg(.ZgI:<X[f=(KVA)KE1bV_G1(@\I;&?&27d:gH[3I:RaH>
JP>0eF=79KM]=dY9VDW<U7\D.I]6\+/([Xf.PF3f;C7\Q4f5P0&^:2GO,@(dZ0^O
35WbGL.e&8@)J>AD]gIO\-\_5ea^02\#;[@W9c^XXf3d-&9[a9ASfZ5B7Nd<00G)
GC\M<#_Lf9fg4)]=e792dcL9,YY;]_,[Cc>g&^=/-&P[+C1[;3B\).>VM.[BZ7aQ
<]-J+.,C@PE&@K9@=6_EGM3?@7KbeF61Hb3OAd46WX7daDb-4NFK@FTeR_15&cB.
]@3#W5Z.JQ&664CN1VHa(RK5N4W;GHAD4+Qa;ZB#fKLJ)9Q][CEXg_GHS6M+#U>5
4K?(&<6XgB<2]-K32J=4._c9@#>79S8#AL-Ndf1M3b(.a[LF+3HH])<=2QBF0QT,
[&VOd^K@[:.4(JWV^caCW9=YdLO?OGPNM^J,(IFZFUCT]H1G&2[0YI.,\+[/,e0N
MP>K1SR41,<U4?K<]>F>BL7d71aRR3+SR;UJIb,(U7]?D64B>c.U>4QJ(J,&0(QK
WP@Y0d#E^e\0#J0CA)4#e5>&QGW?+9fWTaPNb^;?90C(:,I<>A#-Z]]N/Qfc.@Gc
\C]M5gH&_^GQS2N[NZ-@UC.F]R]b=c2RCQOMR9[]Y_4c8f3RTbS0)_cXBCg))@=1
E]ISAD3/7R\\]?A+;H2B^5Y8IFY6HH^]7cCP#]X-FaLP\57_B@aJ^A#e?&@:Qee&
82aONLA#f<0AEK9M/(W@dJ;-\JNg-1OPa#-Q2SUE3PT7QN&/0g-><&2TBI8AE71^
A,N_34&AE:e&SVC,/I)/;AfIU5>fSG7A/^D\^YcY&_AUgT2RD>^Ha(.;(X]B#If.
JZcK^BR_[X,:QVWdLPKO;1ESA,C1JbS\;.7=CgdbN-0ZF7S6A>dFJO.RH[MV[3#>
S=B:^U,NL\T,I]]N+Y^A1_#(U53CdXCK9HR:+O0#,/VZ>UVF?Z&1Y+IAH8f>4NA1
<^g.Y96V>U=C8KB<HY2?6UP)77de35JXa4)=PI/GBVa)Q9f6HafE.)5N]5L>,+OI
3W&W;/Q.[\#6FLC2R^_W0_E?65])(ZbKV01RWHLAP+Y=FE,L3+GcED712<?gC.Y2
8LI2[M5]4Z=Z3<aN@LM(^1<8ZY0OaD=&6<HbN?d[Z8_.LO.BV<E47_(U6RDd#Weg
N.L\3dB=c7<>TMSPQZ;/,LD;WKR0V^;94&e1#+8^GT<ST,4?aUQ_X\@CXPYY:\\Q
LKf7TN_)<Ac=AH&3R^4W&;CZS:V2MTWH4\F4^c\RfYS/K]1)T1/Ke-eZ7g=G\Q4c
VDfc\-/@eQ-;()_);5MWUNG(bVA8eOO/5V^.V>?eg<0[,T,(8O.U()N:ZU]gI<(Z
WO88WdB9CR@BH38Kc4E<(+Qa)0LfMf/:WL1@J4]WS#bg_T6Z(e/HgHg_5=KH.3Ie
G&B-3GbZ0/Y4=XbYbN;_MQ8bf^e/&0:I+f6CA+(9-MPYI=10?a[G=f4#Kdc>@0c6
E?AG;Y6BIaZ8I0FRYN_A_fP\H?dM<Pd/[;P]DMQRSXES_FO(cQ_0&LD#37O=;QLC
4?bfEP2R37Q8-_Oa;DBSGeSK]8G>:SI3UX;)g;#3I2I#XK.;e/6&d0\D1P[JfERL
A29A@0Y@2HaYR+1>.)R9O+#b4E9G;c@8A3Q&@RL_WJ5_2E6I)B4HTJd9=6dbLb@X
12WUdKYYN\3#J@>@KS(VH3fdC#=P0]?9#:eOQ1[.XAEJK?L\.V<X(BG#6Za7QWa3
f4;c&-faHW7f;Dg/7Q_GB.c-]F/4_.PS-CAG?OG[ce^RIdDATg=RM?0C)U^d]18(
ES1FO>-N4fO??.<._^SE66P2GU8=U-AD)O??Q4)HeUd&-2Q-S1,3<()D3N-Z(+<=
5;8M\FH;.6^P1&<&Vb.d[c-44;=M0N31fEPK):-6WP5d:#>F:=bR(_3EEf7(ITO2
+MCfg17<P,dW#[S@J)-70ABUO+S1@Jd?<6A;+F&-S)/BHAU1ZM;8aQ)V\-LSPT\L
LLT_-X5R?fMYcJ#E]CAH,d)c[,B6]UKRU926f&Q==Y,9_&>R(gBc[;:b^<::JJbK
Qg&CBM14XUSE7=R5;H?W_XK1Ag/QA<7^>=8.e&6c?8PDaMG3OVSFDF<SF6[S^T[D
J9/J.U5e[^=DV[GAM6.G<eY]:6Pd=TPUB#^d6/fAP#8b(JOVVV&JAV80ZQ?DdSFC
:#IdZB_PT_;3(Q19A1)]#X4]_Y)8SR^?=KM?+]17b[)7eQcO]c4c-7XQLG;O;2.O
>[gQ^53S(K+7&LYZb:Q?b1W2]Z5I7_A3.OeXV0/4;P[KIMcIM&+@aH<1_b-\@;CP
DHGKVYYSaU8+K:gUS7L2=OI3S7R+22_;@=b3(FOKXd191IBg,++:0,9/;dJI<f^<
GFAd8AJdf0.P\(8gVXEK=DIV/N6_LE-TF;TCAC]@V3#U1Q96RHF4Cde>KFD/S;&V
QBN6Z@2K]dQHC2_T3PD3;FUf-[E2(ePJCf.b=\2eX30ZbeGcD-^AT(\cG_G?V;&_
Rf2WMJ^CTgV)9P>MIL>Yf7<#K6_>(0B73J(2JU?TdK.gYU..N7V>,XL6a2)9+W>[
LA4]91\T7/H-a:;G>b5CHGEcM\7Q)/0?\5R@@EUfP3U?RfP\cA_Ga]W9L6UfC435
cM2&ZcX:>9?QL=E?=d3dGbf8X@+dA3X,c86YMCfP,,39\VK>8/T_bW,N-PBSND?/
?MfH6&(@e+M\C#c>+e=L4<#[0WFCQBKbH9Y7IGGUc8JC8_3ZMb(?3O/(.-3Y2NNV
@OASDOWP#eAbfUb(^-5Jbd=>9.,9(N&fUb=/1RDOCA4)VE,#H5b._1YF7K?gZ/+_
NU)8[6KZ6Ue:O5V^E79,gO];)^e=.UR14NV8Y7WbWG&]+WL@6\\7^8/14RNLLbL]
f5UV2/#?R.9C\fYVP_-dWJ;d7GeOgXf2W]=N-N-S0bbd>MY1R:&>#;5B,,-4CTDQ
3C)K/gDa=eA;8FRcd-84/W2dbO9=GXIJ0.MdLDfB_#KC]6.PIQ+FRN:3,EEXGg#U
1.K8^+6,,OcU=/WO+B>YJJ-E;VZAY.;Bc8DE>aNQ-A-8.bBN<XGCL0DMHW54FFf?
KUL9O&eE_<]A.SfG=:f1#_4HW;<aZ;e]?QT9N78]B..QQ9a8\bK(PP:=a<WLVg<.
S;4cO][(JOHH97#J3dBH\5(BJX-?>&)_B6N=O>(S)+c+.96O=HE__2C0N=MRX01O
#0N9,@eA=@#E9=bJ((^ZR>bS4bY)KGObaCA.^aEPF)?U4SA34HA[S7FcKgE8Nd]Z
@W^[)a;bRM9>eLOG.W\2MH5,=0;?g:53]fK1W^/5NMV>+^2<a>aUb;:]?RZKdN_(
.QCYCV8\?-9\A,HR,M@(d]B)5PfTRND<_F/Qb>.SO[3K+N(08@.ZT&e?G,;,[H_<
>[RX@TEC/eE@ZbQQb)LI.V0HWS-4:/[&](d:#6FeV-Ac-??U[6cbEf]9^U/]@[4e
Y+@7_1PFdMU52Qc+\&_D/QKF.YZU:A<#6(;dI(JO?G8->?,ARH5[6>P7KEU^=/96
(9C0^YVeGW,E:47dOK6Pdf@5\=H&2.@LCLbJ.[ZfF&<A87Na(7.(C9:9OJKE</?;
Jd^8#^dXD3.LZFA9.CMUR\:T@H8d7V/;GW<QB@)(=,b)CBPHW4GaDeg(Y2dK(BJg
,CWJd#G:7]UN9&H]5cHbZ8TS.0C[MSO4,Mb;L:Ud[+d,H#,XaKEZB09V2Ob7MgP/
=9A+dW_aBEP&98.G5eZdQ0)VX#fSfaaL:URNCdHWA))JP<a0?L6eACMNeE.HI#4O
-K.,[79^HA4K\W\_T.P[7&7U;^+CX;]N-eQRO6JI<V:bZ(+&8cb=OP^PaM@D-:c.
+EN^:6cX^IEd6dD\[aY7Y\&-,-L9^D#<]aRcAOP3EQ28+&QgLT_>cg/.K>MfH]IL
b7]0\>cU1N.Y^b#8f/ZQD<<\@1LFcM3.^??PS[?:]CgLV\=V<cT>\=gT+15IK=JT
IM9.Z5,),TE3:MGJ?c\??DGXE5NQIMT?X0?DW1fM(gK5OV3Dd9Fa?aN1,,E.IF;Y
0[AfC&fA#0=RJ;0)S&UT68JA<(S5A&UXTKUJ=,8LJEAMgd:?2+a.DcF=>3#ON#:I
DL8<?/,SQ;+Q^5.ZcOL<))]=1;-7;H^2TZM=[8;;F.?KX]RP)/:OQI_W.7]MEAP-
^ZcMJZg6Ce/&+d5,NYf=:77dBfB-8bG;#;a5\Z-MTU;9.3gbTF9PW\Uf]KK;FFGO
A)WKR2+O:SY;&)G.N)@gOHSf3(V#=1g.cDW9>/CM[cf]f.^VQ2CQP[]C^:SaT8M&
ZKB9L;;QG091;\_\)9>WT_]<)=<V)1];)&/B=_,+9)&+\#9d6)WcS.3H6@L3(R@5
CO;2R367Z_g(9EU8.(=[8S?W=QZW5=]HC6F/LB;=(&6WU8RB2R+X5GOD1>MM5SN_
Z\7EKee&Z&fYNdgRVacR0a)S@JTZZb5[UN-W\]/g4a,g)g]GCB/f<[)T;ICL](a=
eW&)EYD+dDQDOFL@JeLL7gC9g9FSg6)0[O:O)\e@/MU?BN.Y7S1U)-8AS/L3MN=/
_0\.8E4J\U2D2cNX94GZ@;&96LI[7(>5C8dKfZ_b2X9-d01B97CTWg=.Ofb5_@)#
QgH3DX^CZ]9VP^1[RZNGZ(YQHQ0[,FD.9QPC16/d+,dc--N.K-Ic.,2S2[QC^MF5
#+UXNLcM0M4&eC(J?KbL3c0K<M_+L=(>YJ&;Rb2f.:S.DHgU,HMESadJS,Ub#TPS
H^Y.R<YRKR:12KZAGE6<Z\]T&Ge2\14(CSNUOXR(G-#7Re2>2<cc<@a=f^]7dM/d
)-cU;@I-3BM.P2VFa5ZK@3;/-#V64/F1-#Z/RWC[-YGaAeIf=?#=Y6D(G&D/,NSV
.ZIO7D<^1>PQ2BQaXQ#_8Q20&P5+(6gBS+]1LVObC-)gKf=A+g4fW&#:6)gDQV,W
RE;a?46.2W#+aX,@4AZ?X+@gBA1OH_0g[7ZLNcS+eH=f?JBac2_.OT]-&KeE=]R4
K?42e2#Q#GWF_V2PPLAb6FE6BHG(7JBW3J]^V<EY<QeV7cSD]_J[c3)0bJ/HD.f]
B@#@5LDE55(;]V+GWFL.3\\g5;ISIf-3;G(.eK1BUYc,8:.NgK?[LeW4PZ?f]2:X
HN>?[-?U7f9@7#8AS)MX^(60FN/QMT@eGM:bS)3+_@PTf:aDFd2Rg6dCKKe>Me\9
IW\&?U[a2RS[><g:b-cbAR67Igg3+5\gFQ?c#cG?NLE;S4ZJIU;CIeZ.^Q4]3^_F
&B^/+d3DI7LEgWIBOPeg5SEXB;N95WVCb)D^<V\:7D+HaK<S)D[J#ATA\O\QAT@L
092+HI4DA\CO5gV-+7A^bZ0B(,CI=(A12gA(E488V0CZ:16]DefC@X9fN3-4,.bG
28IdQb)1[5EMFK+10]V(@7#dbLA>8A0aIR+cbB45]fIH+J#,?FH;]4-SfS[86)DI
\JN_4Ubd,&#&;e7eMBA#gg+9<af0d1+(@-Y],K[8)TRQ&?E(V#YFA=?CV0:U@:(g
]P1.3TXaee\8d6Tc-V)5#C^a^ZRKA^\QOZB]c,[-]GZ_-3T,]a<,/?#.F2@[9<_7
F;ERG&90QX3UIHd/C82UcPg7LDNCe<?HJD?BWb\DJ@aYaHRg7@V#L27a8gO+IM=>
0.Wb2gCcOOQNgS)?6?M14#9\):SO@X0I=>.fHT(R?X9?OMbX\Vbc7)S&+D&4Df7]
\.<?__P-FDJ,EUc6BT1.@3>3I05IB4T\U[:]6YAT.6NN;Y.LRKCKH&gKg&IcB97T
WK^&4]8Zf9eCATOZ@J77U07QR8f==cb8eM:DgDBHW(\WL+PJ6T90GM<;5R&]OBFM
e;#;5\?f@0Hf_#9\8R3bg7EL#8LbW[-4+0BH/;:0aHQEDBUY)Q4g8;(:N&;.3TV&
<+.FN-H.]J<LSDf1\EYS3^eFLc[S;dc^3Y.HcINC:[<g-FNeHD[3R/^/6UHB]]:6
fcE(B,a@?d8D(&C_)#G]0\0]&3g77420-CYSVW-DIY2+/QO)Cd+D+P6ZU+KJ@3>4
K1b5cF+VRQ^OP&1U_.^aO(g-9KJHc\4A3^PP13A[2dGLf>2=4^?aZU(JXe3TDDLd
UMF-Q(Z/:&V#bZ@P(NW04<M.+A-RVB<C/bbSVg#Ue3D\?U7Wf:OPUN9AYD8>/^OF
\05T=?gUX4O3=d42/0W@_T_IFcd1KG+Y65I+\XAHK;6>\V[X6+(:X<W#(@<PN1_:
U4V2GWSdCbWg2gNJZB^3+QCNLbG6A_QaU_#7#V1d,[#Q<>ffR63@690XV+FUFZ)=
1]Ka>&]SATJ)bQ/KHRM&?1V@7EbW98J+8AT91FZVO@4e9P@Hg_gf&IC5#R9LgE02
9\:=6dDcFB#dH\8WRG2)@-A=-+S#G_#/\#2f0/C8YQ6P^,;<bC9^C=MO+f<^E]Z(
DK>T5<,/+?8.OLL;=SHUbS2YJ)FXF8+>:<#=)6^DS7;N)7OL)@/B@H?K^Z3.4:/:
0)=LDD]5HR8=)gZ6OfPYfI/Kb5<=>Cg#eCM^+F;\-H/?M)BI^Q\,/JYB]M9_DJX4
3#SE6VZ79J8Ma1)UeIOYad@&FL5[)T@a1\UMIN5\ZMHe0WF=92(CCZa89M+bc=++
\8X:P@)N<J).K&O8gM<BDf^F>M)YD4NB@Td\\@=W2\NNTBU&:J&R?KA^2RL;]cgQ
\<BI(.5[M_N8W)2/X<fR&MUc4R#2Ha6NFJ@91-EPJ5b=<:?ID/MADO]Y.T.dQe2[
dedZ>bAIf_Y1Lb8]-?#<ZdZ)?V4JG/N2,2RO9Z4VC9</KT<2KZRIe&-_g6Ng9M),
AVg[P1#^Y,g.]])I:Y]L^\FQCOR-Ic&]]@ZS&degI\bASE/3?b#AE(J05M&&[)(/
^44-YgC(=ZAFU9,>K+.CRU?+N3ET3_)F)fN]S\HU2_^+FR@EG^FL6G?&SD(72Y;]
WcSdUCQff;35HY]&<geGeece5;9=G\>gEfM8O)IB9F^#c1Y</;=U49^/KPYKgb(^
]e;K5VIUa7KcS6HOgDE3G;K&ZGT-KSR-<7S\QM_^S72Ba@CAcF;c6,:N8P&[187B
@bST2K;?=H)&:fLg@LMe&>WGH@&Y]?S7ZYFSR-+QUGPJ#3N:;ISX4(&fNb2a7[;V
=XF207?g9G0EHIKX@K:A2;e]c?#[T9BQPDc+8._g(?+/<(b1F+FQa5dO-1<Jc7+T
MdKY6OfK)T-@HSHZR\/J98Y1)L17>2\4Fa6?Z6d58F8[(PSR0QK#EPfOe6+>_/DU
BHHY>fKC/Z(H?VH547PLDG+DOO4]7-#R&8(8IH1R;GH^&e9O+B6YP4C)Dd>Y;]C=
,AaH#9,@#Zb?KeS[_FfY8I&Q;,ZDJ24&<(@_9Tb6E)B#L>92<9cd?VR@YXTB.>SE
T5H4Rd>5T2d&Z(ZDU^LK6aaBa[[FDdJ_B^)48TM[O(\Z5fa5gUOY\#;g?e6W;BW[
K>=Xce(/,2LMaD:OIT>B(gM9SdP)G@[Z,W?S>;)gQU7XW^G_NFdWLf;gM$
`endprotected


`endif // GUARD_SVT_AXI_CACHE_SV
