
`ifndef GUARD_SVT_AHB_SYSTEM_MONITOR_COMMON_SV
`define GUARD_SVT_AHB_SYSTEM_MONITOR_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_ahb_defines.svi"

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Py4SCGY3mrzSXjGWNbwOvChvb9cZOg1HBQz85Q0UevEGLi4fGWf0TH1q9I8pS0iE
mlOGcE2Ol3oGuBZZUpNy+3wMOaQ9lomjf25OWylf9mp7skexG44l6PsSFgCV7gE/
3YHPPcFyArRx0V9DE3hweCW+usMGQ8BVI8VgBqrbjEE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 3532      )
cIuSS+SXiTr55+D/VcGx+00w27vy3sr9vl7+WgqL1pNRr5wKWDqThKqfzV8BN9Zx
uBvqAs3ZHzj31fFyXGRltJonHmalDMftztuN5DZ0+te1SKb5WOhglMcZwFJXdwoM
fIYSSeBfnv7HtHzeM5AcPH6izWFD6proScHoNrCZ+WPIYkhQspk4jZegUhUEErD3
C2z0e72GihvsMzaA2u8h2sbGR0qyQpi832xDsNZLLT9zzI1BCQ2Ddq/sQdfeMqmD
7JNBSUTR9gsyIffgFOVvyVNGUZGjBofTe2kGlVuSrtU9iH95j0A6zt9G6YT03/lT
+aILSyzeiLl0EmjaSDnxhGTzZZ69MxKVY6hJIUgwzjRm/E9ZXLggHm3n+doUmo7k
PVe1yN+RatRJZR2BDRIF2cc8VI9NlkdpxedFOwXMx9snKbPeChAL/rAS3VeFP8s4
jMJH8pz+Jd9qygs6VuiIWNW9FMPX5jK/GGe9QArLlalJI2eNcAvIaLtXHVSoNtg8
EWQWEMFdKYA024OSndiMrmFtRsJBhHPTB8luwa7z19fHfrHJ0nAnNQBw6KfKVWfI
q0Suyj+wF8iYefsjWzYx1QbIKudazYUajHceUZONyEDLu3MIyWy4bdYbfsNvcNaw
XDLlBtEjWlaqIAy8ils1GaHfx3o4JvA8OgWsHVffdFEPzwfhFgBZfnRci+VE7qMG
kBkqEfVa+L6bL4B/Ay7N0nt54p/ycEQyGT5yRQyK5IXO82rcr1I8eqM0QAgtMhd7
a0BFRAtGICkq2rHpHSb2HGfgq4MYeYn5Vevfk2MTSGwynsuMRc2EqLydL2EOCB6o
kEzi8J21KSoK59ZW10f2acdkJEfJFoK05vAG/xG8UFgvEi9UICeX/O5tLdnSnLd2
HuPgU7D5c9xgvMeqD5fBQMqBPKRB1L84fQK6PlJYpYboO9YB0BRzhD7ptmU2069H
rIGZ6y+DQJLR2B827bq/k8om/nuj37SOHL9Jr59IjutKoxSDjHCnhy0aZedaHLt9
nNXEQYtgDgLIANZvDoxrnm6RFZraKTlVHv1F9h/Nfn3kCDjkCyWsCVJI3FyeDWJi
Um6hGFKX9jx8+M2dnccUwZVJ0maEfzLHtAebYYv3fL1xIkFsOIhvmhOmhR7oHhOP
RRsUjXb3Tslbgc2VAEytxwC2dtPnHk9LknNzPllT9OpKOrhU/17q3xpnjexRGKMB
CmaeKxZtQuUdThskduSM3ssouC3q1TRzA+ewODwfRuHAqbY9hnt69KIZFhlShb6e
Im2nFq7q/UvjUgK6izbXYTQytvaMD7/mPjF7Aqd5d7+rP8OI3ER6XS2VpFw9Cl7h
SJ+YfpxpiMlWUpvnOc4WNjSYlMH9ZtoSpm+VMWKkJ9WmtN7OHFOK3eSl92gW6tZW
piHVKJ1ZPK1BxSV8IZSHfgwsp5ZRa8NrkdfhbJhaqN0XYrdWy5r/TUtlGNhlQGaH
ROJaB4xWes4iwq3LxjE4TnECkj6z2zpLSOr23z0M0Jl7YB0rR+BVEwowgqgtpL9M
zFY3FldJ04xOyDZlNz4/3NGP8ezh1XXb/Pu/C+G8JsdRs2QUkePQd8p0eS/RvIGB
Z41bCFLPed/v3Gm4gHT1LNU/VdBNoO2LQpUx1kmJwkTU3a4dg4wxQk2+FiG5+eyX
mwYqbiaMptDxgpi0nKe1g2ztHhZIav3UKzPsJIixmQkXhOqsEks27/FBhs24wYBU
a/4WeRlDRT6aw7yH1RbbmDXlz/j2ugspP8JpcxLub8kGK2ERAyPM5BF4gG2s4a8t
lgtqFOjuMVKXOoPMf1cuF1Ppw1hAygGADxJKGl/1f3MismofSJdPBUfgPWvUHFbZ
+YY76i5/rp1rtSqJQ8MdZ3Zfh7a6m2+B8aL6YY0+qP9VptAKJl5g0FIim5iLKdiR
3jRlmnSrUzMJZr8FHbzQEVy9cihr7i08yWUbkJYJQSDdIxkg2bCqriTscgOQwjMI
EGM4bEXYvru8q6MP+hbwycbZmtcocJ0a0ob/Jf0TEB+nJ/98im5WoY3pVtbwngzl
cfO5g/bu7cAPqG7lsb899gAYIjDVx0FCYX/cCLDHe51c9iJLw05EScwoJNQiNtX1
Cwt+k9fnBIflkrGgi22naOb6B1SozxdSOVpAENS0VlZwNNGtKuNnqmo5VSfUNPVt
e7lSe/XyOLM/GZAbnHKsgdeubxR3sUwSDGaJmAwl/AOs7VZ9C60MzpUqGjx6umyK
jniYpUkU4naDFpFnyvJqJQZ45rtb5EU3yTvJZnjWlUXNogNOml398oDAN1//oaiS
EInWDkqW8JKIlJETFthOS/LqA7R06BnRAa6pJ4CchKbtlFemhTKQZeGDMACp1/2U
34ozqgyKdv5PDcats2T0pHnmQuwN5nkWlg89wTM+C5HFzy9A5b+NoGZLeOjxY33z
KZGVZssNP5DtmQFncn72o0/2gA4J6omvNGGwqzJP2ArBwQ8SX6Y7rwyKb7LdAE/0
pSHSVPXeec0y9I7NdizQzN1rWRZwziCcG1/BOttN1CX9pUiQWdOeFJrxpCNvPcNf
m2yFmUkUKl3g2L/x9cxY30hOhGXkMENh1wCErypHD6HKAcntgOz+6mr6iIE9aLnX
P6QagsvX8tUe36R3LFdgmXpqodSk6cf2aDSkObdCxeJmgmZEXyPBWXHmREzDQOsw
fH+4IulVVcmclxEdnXsTi5acTCbTQuiWo4Ii2W1tnqrG/fUbiifwvsh5jS8jvaIg
+8v+yG2taAju3Y+A4YrgokF5trVeVD63Mw5AxV5EDPt9MPp32VQSNCOIltMEmwey
7Y5IGjIn/rMxh6ra6Ktdyhh+gceTKrHi/zddEhKN2QCCXm5Zjpj/ePHgeGC9lMnO
8OguDzTBj4OalsSYOHS1thXCaI7SLtk7AW/qVg179lfeiLHf4IprHTX60qHiNGtb
IG4aky/O+yV34BAypSN/7hdkFuh1vzY3eo8+KhS1CPoCWrkeX7DTiF0B5PMtykax
2E2RbBfiPIfDado9gqEgijRHxV/Feh6wBmPz1dHor/WPGFq+4q99PCmIVWywiIJn
Nr6cqKAdOtcZhIM9rdWX+ZZx0+irX9+onNZ2zHnrvA1wE4vbMbw8htGYrZvF7kiD
zzZ7Y8OjoSSZ7e3prBS+pBGiuZeT+nw6r9/1Jg9pMzfFqEhVlFx0MEDEBRZiqBbC
9BxZarTnPT5iONpsJ/lRNrCrHgrcygUX5DkamN1Lremy84dNErQbM8QoP40VzOaR
MnsgYd4EBbJz173pt6ys1ZJLmtM3M3m5eTbe2KHPFieudQv6xnOTughE5aRyJyqP
JREKj2MaxMhHmehweoxZPbe/oqPqE8oqinyGggFM2HeWBGF7NKIT4FxMDh52pB0d
1ylgRJXgMOAYE9FABdcb5j3fZcingIf75J9LAGaUtEe6J/2DUmHj/sQTXz07zdtF
nhTRiUou5YkmjMEaqudXtiWL2eVJqOJOWVsuE+gse2OhbSgP2tWLpXJDF+qqvhJE
YM6vtYuOP+I5H1TzqFPvjWunAU1ypGCbMjH8Co+eC0PmoKBrrfuUEGAx6WMpvU5n
O2yklh6rFsFbqz6f9y4yM0VLlm19gjSr5HHd8uArcmYVSRa25+oV+esJV2DH55jo
A6J2Ovw1HLxc5azBKkA3OSB5f4guehIS4ULDeA2w1YV1/euK3ydv4R/ooHf0XDCF
4bYLAdSRXWoZtjdCAs7HO7AD2ck1kcqb2o6gzaaMe+dxZCEtQVDJGRPS6fmzsBWV
wdEJaHHX3O/ssDWpTWhiM11JSldsA/aUa2UBcOgI5LbXDSdmo2bFFaD4SGzU/hmD
ZHuVGEbTz4zJ5tjsawOVDQTYKvCXO85FD6WcyiRH41vqgRKg4wn7CdxL7H51XgSq
6i1PXNgmxoV2fpWf8eCeAyiaPPa9KbUvRdGz04J9MURcqGYRX7QNBiJ57YDPng1g
LA1SpAPfT3GTBFrx6IhO3oBCdMkw1q6SpGoPMf/kzRxrvz4xIH8towyp7D26ay4C
wJOX/fejBVrQVyn9mFfMHV4zkw0oDIGinsfxESXbt0uRb28jDPzca0te41LKLVCa
pXt4flEbQpM2fFo6RwWxZ+DRzBWgTWr+WcNMLOj2zh+ui2UgyVR7ePR4JiKDpzwl
yLwre3PVU7PRo39nlfQ0RdipZRB+GHbp0IWGCeK7C7VaNNnP3wZFbeR1HL44xeby
BhicQvbKBmyXt4jGlE0GfYHmONEIOGQbcu64KeEJAllsPqUg+f3HWHxWhMQb2gEK
m4C6FPYqz9BAwzVvnlHqPA52kN94TZ9mLd6+V7l2aYtqo7n3iAFieMfODxrZ0PQC
aHHDTZT5YyXmwGthMin8uDqYFMJt8UVBPFsEwgbOVhRcyTDKL8RYERy/tpbYKq63
eVbdvzqJN+4z4RknKw8d/gPr6MFyh/2InBkWMMOHqz0LvZSwDJf9Aup7lHpSglTv
dQZLaUaqfDcSlCxX58602kneEOT0vkC+78TaGnd1D219a/hYVFN0PqdpkJe3sHKl
WBi5hjCXNWUAUzXGxsoOOFJM9sV7KJiJodatNb/b1Xl0B74gvUeWLOO4IL1qGcvp
jkOR8S8tSZSiVULKotiesHuZgOO92jXklcvaNNT9TZ57T2OqecxH9ui7Opm6HZzy
zXh/WX+qwwdQK395qGMSP1W/3QWVsDPjCamqOU+3jdU=
`pragma protect end_protected
typedef class svt_ahb_system_checker;
typedef class svt_ahb_system_monitor;
`ifndef SVT_VMM_TECHNOLOGY
typedef class svt_ahb_system_env;
`else
typedef class svt_ahb_system_group;
`endif

 
 /** @cond PRIVATE */
class svt_ahb_system_monitor_common;

`ifndef __SVDOC__
  typedef virtual svt_ahb_if.svt_ahb_monitor_modport AHB_IF_SYSTEM_MON_MP;
  typedef virtual svt_ahb_master_if.svt_ahb_monitor_modport AHB_MASTER_IF_MONITOR_MP;
  typedef virtual svt_ahb_master_if.svt_ahb_master_async_modport AHB_MASTER_IF_ASYNC_MP;
  typedef virtual svt_ahb_slave_if.svt_ahb_slave_async_modport AHB_SLAVE_IF_ASYNC_MP;
  typedef virtual svt_ahb_slave_if.svt_ahb_monitor_modport AHB_SLAVE_IF_MONITOR_MP;
  protected AHB_IF_SYSTEM_MON_MP ahb_if_bus_mon_mp;
  protected AHB_MASTER_IF_MONITOR_MP master_if_monitor_mp[*];
  protected AHB_MASTER_IF_ASYNC_MP master_if_async_mp[*];
  protected AHB_SLAVE_IF_MONITOR_MP slave_if_monitor_mp[*];
  protected AHB_SLAVE_IF_ASYNC_MP slave_if_async_mp[*];
`endif

 typedef bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] ahb_sys_addr_t;

  svt_ahb_system_checker system_checker;

  svt_ahb_system_monitor system_monitor;

`ifndef SVT_VMM_TECHNOLOGY
  svt_ahb_system_env   my_system;
`else
  svt_ahb_system_group my_system;
`endif

  /** String for storing information related to transactions to slaves */
  string master_xacts_str;
  string slave_xacts_str;

  /** System configuration */
  local svt_ahb_system_configuration sys_cfg;

  local int log_base_2_slave_data_widths[];

  /** Report/log object */
`ifndef SVT_VMM_TECHNOLOGY
  protected `SVT_XVM(report_object) reporter; 
`else
  protected vmm_log log;
`endif

  /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /** Flag that indicates that a reset condition is currently asserted. */
  protected bit reset_active = 1;

  /** Flag that indicates that at least one reset event has been observed. */
  protected bit first_reset_observed = 0;

  /** Event that is triggered when the reset event is detected */
  protected event reset_asserted;

  /** Event that is triggered whenever the hsel is sampled for active transaction */
  protected event sampled_hsel;

  /** Variable that indicates the current active slave id, using which the 
   * sampling and checking of hsel asserted for valid address range is
   * done. Also used to bypass the data integrity check if no hsel is asserted */
  protected int current_slave_port_id = -1;

  /** Holds the sampled values of hsel from all slaves */
`ifdef SVT_AHB_MAX_NUM_SLAVES_0  
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value[1];
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value_copy[1];
`else  
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value[`SVT_AHB_MAX_NUM_SLAVES];
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value_copy[`SVT_AHB_MAX_NUM_SLAVES];
`endif
  
  /** Semaphore to control access to active_xact_queue */
  local semaphore active_xact_queue_sema;

  /** Internal queue where transactions from AHB master are stored */
  svt_ahb_master_transaction master_active_xact_queue[$];
  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifndef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter UVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_ahb_system_configuration cfg, `SVT_XVM(report_object) reporter, svt_ahb_system_monitor system_monitor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param system_monitor A handle to the monitor class of type svt_ahb_system_monitor 
   */
  extern function new (svt_ahb_system_configuration cfg,svt_ahb_system_monitor system_monitor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Sets the configuration */
  extern function void set_cfg(svt_ahb_system_configuration cfg);

  /** Sets internal variables */
  extern function void set_internal_variables();

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Monitor the data phase signals */
  extern virtual task sample_common();

  /** Adds transaction 'from AHB master to IC' to internal queue */
  extern task add_to_master_xact_active(svt_ahb_master_transaction xact); 

  /** Adds transaction from 'IC to AHB slave' to internal queue */
  extern task add_to_slave_xact_active(svt_ahb_transaction xact); 

  /** Gets the system env/system group */
  extern function void get_system_env();

  /** Process this transaction and execute relevant checks */
  extern task process_master_xact(svt_ahb_master_transaction xact);
  
  /** Waits for transaction to be accepted */
  extern task wait_for_transaction_accept(svt_ahb_transaction xact);

  /** Removes transaction from the active queue */
  extern task remove_from_master_active(svt_ahb_transaction xact);

  /** Checks consistency of ahb transaction data with memory data */
  extern function void check_xact_data_consistency_with_mem_data(svt_ahb_master_transaction xact);  

  /** Gets the memory contents as a byte stream */
  extern function bit get_slave_mem_contents_as_byte_stream(svt_ahb_master_transaction xact, output bit[7:0] mem_data[], output string target_slave_info);

  /** Gets the address banner string */
  extern function string get_addr_banner_str();
  
endclass
/** @endcond */

// -----------------------------------------------------------------------------

// System monitor cannot be supported in the INTERNAL ACE TESTING at port level
// This is done in the tb_ace_vmm_implicit_1m_1s testbench directory and
// the tb_ace_lite_vmm_implicit_1m_1s testbench directory where we mimick the
// behaviour of an interconnect port. However, these task need to be defined
// so that things will compile.
// -----------------------------------------------------------------------------
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
C1vMu1LUsfi/Ck8twJ5FtdmhLM6TUeGKxM0D+Iip9rxxItwtgFphoGUMlQ+e5xAW
ZqzdQ5JK6Edx3CF49kocxjZEHeBq/UTXuLkVCk5yZBlxIdeWPmALxvVbbAzAN5kc
/5EEvEfh1l940NhST+rVypqIQGMwzTj5duZDCLscR2k=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4126      )
XSi1oQVw+I0jilaQ3umAnJoIBPqqwMVK6sxYHWYwz3KC2AwaLzcO8CimmZevjC4f
4vvokaLH0zDPNoGzahgUi/fJ88H3/m3IBgWDtSW/tsafQ+VdKvAT1bFYk38FBg/1
y4tbhDMpvijSRKMF4U0W0mbNOagRkAaHMDn0sEY3jSyqhPULvdN+QuU/j3ZD4eZB
FJLUQOvxQL2Q4KdOwMpvDg3Q9j8rBTVfMEMwACJfibjH6F5Ai8B7NZfkDwYiXQ/+
qFegMQaCed8Mil8nSet33EJZ4xuk07GJl+i9z0FG/b+fdgnNNHssdWBCFV7i36vL
PBlkfGy4bNgyW0WU0WRygXUvC5qNr9LfNZEXp5uKzqufnGbECuiRgP81xW11JEVs
EPM3wSq+wQ2Zh3n2UfJtdsImh7EsW3+rQ9yNlBeSfY7gWRkcHlOgTpgkGEfBAZEa
8t6C5FLnsVZD5oYzKleCrOpTQk0YkA+NbqQRebn6CKjjiG+92bluiUVd2SqFXFsn
u4qD2o1djdoGK7TTvaYIuCbG7MMYaX5r/a4CNysLf3A5x8NmlqA/7RumOm5U4KGZ
VsqWMB5b/evEtQTiJU0Q2WXKvc1YcqjHjDW+IkIQPWmHxlNQVLZy0CG0T5Ds69HE
iixfOnSf3ZLgdgkd5B2Y/kwn0WNKFFOKu7oie2Z2ZXhWJatdhWm6qH5qsHMBDSRd
unNRQGeTYqQDCXAfkHx9tkxcXHEOUl3bBneNEuomSiAhpL6TJQPdFYvVoEkkK0LL
sm5rb6ub7jPU3udGHYtEJscbW76slkGgt5PZQ5m5n6Q=
`pragma protect end_protected
// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Vc1wKOPXRV94+DiIxonchzObKEo4RIyKNdLrHLuMxyMeGb9NjMBDn9iyZmO3KhOI
MrtTHhSYRgmOktgkv1R0Lh/kV3C/qEJxam0JuIfdXZ1mKj1KGiT7JbiwwO6oAuQw
zW//S7bMseG6yFNuvbpLRxGIJSY1zMhZPxt/VgJY+1Y=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 27393     )
KbKFHGD0VAS8tdYIFftH7NVhCfm2+GqM+Qkp0Vtj83sclzRuZDJ1Rt5FkGuREU/C
uKU3ytmxqKlhPMTrbesGoaG6CPS6NrxHX79fKg5FmeZwxvPv5D7ycOQJrw2jO6Cl
HOuIzXFcWPK73WvlJcpNwBTBq53SeSbpRVQ/65oyPKZt5YBawJGI2XraukmOH1aP
beHckalp8k7GO5wtnmnGllguQ28MCl3UptxAhsjPjU2+/KJpaniGhLc8+zM4JTJS
YkXWzbUoq1Grb0hM4Vy48ame4WrJXHJBpVvREf2/72EnDxV1tqFauyObEj6vHrTD
0LSVC8v6GpGOs+KuwAg73j260N8MciFsPpspo07br+3X5Sa/Bddc+xoNSQbTzcyr
mDQIjt50gxq7tktJI5M86Ct9NSBUBiR/VjoJydkQTq3b3rVc9xgjMbdCcMz5LH3C
ZH8h5PM3uq7+pgM67F5bRujO/rKzQJXLHCXj32nHF1MmHq4fMwR1EALoiBmSJ7ez
SFnAt0420QQHAwBFJbkKI6YJgQvrLbCjXV0cB5ErN367TEeIgW4jUW/g89MiLva/
2rW++JLQyuEyasYp3gGnhBp2mHw0dt9naDjvHCym/OiSjnISIlSv8Y/SMHmFkn3+
ZQCCBssCUvfIZff4E6Kn4/SSFyo/RdIV8GLgGtNfHlOULYa6dj8dNzIOQqF6Og0N
fKZrbe0y/uOA87Gs0TxucRaCaP4KV9pUfRHcgBBear0HiYqWYAB7edFS2VLaIDJY
1K0VjpINi4mxXBUVqdozZ7q9o9GI4Px1EZozUZHaTdOoej0mfb45QHhS+17U6A0B
CAuRdwLoiJqHUbdqmZlVeRaNxMK5wOG6ugtFEzRX2USJsFXU+us2fNvOfpT1qV0e
y+cEQJzR5szL9vBoL5eiPPiboozLkbqSbBxTXrcAkJv36U+Z+/GQAsRmXnSs4EVg
tiDLyJMvwHDp5EK2RdW1L1trUDJ3Jri+UGK7jfhY7ZjxfOmeU/MZO9rC/zEGaqXh
J5w/zJXAdhkdjhuyk8QwhLB6X4H/tK+Kt0VtMrBt6vG5Ym6mcsvjmXNA/TPYA+2M
vpSw9FOLH0tmNR3iFdy23Ye+VgTyf+r+GsIddbMe7eMTKW0LXfhVzaU1vhF2VooC
uk3GdjDvbYCXT3Tq2+PdkiW4F2nTRxh4QoydXOOhNFym8N2l4kSggfcUcSoyfgnV
ozBATYl1wnXS5pb+87RcV7JXAKlG4nRf60OTZ2cqXfd4vhUucconTLv0aC0CblSG
Hkl+W3PAF5CiNkBzKPIinDNCeI9BZT/fk/6tI7UCqix+4M4oRRnZokMyLqXh7mTD
be6q8o7MTu7yhsFMKyg1c31TQmnO+KCy8sL/8l9K2ud5QuItJqwGZPVxgUt91rG/
3wsCmYsO00uNr6gH6iwajOt+LQA7o4Duhfa9bt2EA0hhtaO+OW4cg+fZ1iYfJDYc
k1whcyWJlLomYbCVsimT57fp2a/6x7JUoVP5YyUl9FYlsigcwL23EDIvxYzuBaun
XNeIIK3gmqbZ28aUUBT5lO9ADkcvlKtW5DeoxMIbSUb1fThZFk+uL6lXbDRHYcri
E0ypt04vppjJvZPBnCzo6MUTM6gYqHwt5IpYeSVQiLc5iiAR237JwGZGy+86PtMr
mE/As0Q4JR5WfqaVkynQqL6JYmqJvb9F6aUiCd/xc+2Z1ZT3VyJsyIGG6SU1qDUd
tazb1rrOAI4QGj++iEqVA279Ap18x/XGnRalxVorYua1+YCUl5mWIbxcpJTAu2Qh
92xaDG4G4thptMe4QkkCKmI+Qx51G4ZovsMvRKsgOmb8+Z42KsWdxS9YqaiRou2r
8pTJIA3dnQAdG3MAIN4IEXQSw/3a/uZkshK//pcfzTRIzrFmokjyryH4dfIhBHGp
jqC9PSq1YyzFCVdwkK11TqkWOMLLGP3ZBfPa/ETp307Z4rbgP2a/THpUhdRvSCLc
q5Ib/JtY0OSn84vgnSvm3/eP2pxf9YTQiysFFE3P4Gfd2F/cKrgPCOMvmsz8Ndp1
t/J30F1UusCiQCrrTScBCQb2qS4/RjnWPao3lENuxKKe80nIQinA1sktXKLMWTMc
TwhNiKQQFL36C+hJsHZ0qQKNazSSiX3b7gtuJdwhsCB+N8rlxhPh+LZYMZkT9jDR
RI27mkvbCHdFoJoDgMz0MNRsKVB9XJHDR60CbEW1oNZvDIzN+Zh4PhEwzIwUhDM6
9HLUJ9nEB1l3JBVPxINIlayNV5zi6/5yNsm6jeyOVkGxFs3eXs6s+CbbQ9DSgIrE
LAehjJIgggSVcaqy/1TgsghOsHnLYksm5huwRs2LKFUoSyh0j1XoRkaJWZ8pgnmN
iqNwbt79h1+pxEERVwQpGcxZCfept0bL3V92xyOoElcsVpVJfpv6CEkDa/jeDWF3
CON6HyNw+jdPQSll8wbA56fNzXITBNX4awCjCjflxItjNHTy3NDQtrFPB3KMjPwx
Ndamflk0Ee5MB2xARnaQENmctaoyzUXqaoUFOKwyhlWUAfUrrKws62qlvDs5y/Rg
nfZe2has7HuIGfkVo24LmdE/dslJBdl0qSsZOnTD/HaawgyUA9lCkPmu9n5bGTUE
KaXfZx/2DKFRoXXYGhwBT91Er8+v6jDBOq9YDioCXwWgWrfYTmVFCvzgq0gJ1u9W
R/028pCtVATInSWROgJbm8xq0Eq9KqAcfcbcv/Azd0aMYLETrdjTeck1saRA1igD
rwZEXvyHaSMkKVeO1FrcmwMwyYsDpnarDaMY/kWT4qRml6YXAbAQWBaEi90SOZXW
OFihm7bUCICzncdcqAAYw1npq7RPvE02izI9I4+Iov35kLf3NWLsRonFlY33eJGi
5vi0HhjUf+yP/xLY5Fv0BLZeTG+ZlfEQvcnfnKTOmfkmnqWYgs3y0BnvD0Y3Wfua
YZP4QNfzOWPSuwf19kKYemePp10P+1R22W8NcpGRrpTbgc6nNGvX16KXGXX4n1AV
P3WECedrcOTCMAIagreHFjTQFGZAXeigVbkKUcqzh4hQAdBsl/gdRyz4Dj8aJ+iQ
LwEYrd1YrtoR9JQ9nstItBz4T3h+QSN3PbFCD24R7qsPBEISzXd+sjpQ07PVKzzF
Fyd3r5vLW+k97QvthvnvUVoPM6sj7cdYiNrT18Q1MHWCoa9r9FviVXeTHSso1cDy
XXJEh8OIPHrR3Z6tKozrYGp22ZyUjaDSTBy6wPBCigJfuXpTtTAHlVpCEfiq1qq7
P/FjGQ56u4knbQ5tRtw3ho5T5ch4/7SRntfO1EklEVE/k7v7hXo0M4U81FCcATto
QApB0Vj0pFA7AlfzZccAcOQG/GQsOhy0ZBY71cIOD3xF+pj8fkffCvVi1gqFs4p4
3GLTtmSAAFQfN/nTO6ohll+q+/ttWBX1hv8QJx5EcFq/nq7ziL4hH6/EqcMqEeQv
gk3aVnbzLALX8BkbjVLXAKHwAuOqRR1WiqorMQ+AxjxJisVGsDuN2343KuZ0Yfer
XNyZaxtZOnduqEgk3cTeprww6HbK/EGaHFCgr+QOuURYFDnelyuPFz+1Y93TCUW3
FnoSRxlkj6HTwZLo9caiQZ2LANNt7U+87rqjPPhWqpTArJUroPyQ7Aq6VZe4Vuov
txwFLbUNLlXG6QeHkvDuIDCL05sC1PLJPJX3vw6uVUPLoJERcymBZAOxNut8nBXo
UphQZ9cJuKKKqV6Jv0S6EhhAtsaEMmxWhE8EimLIwFoeNAJIxZ6QktSpajQItEa/
ZFG0f0eVUiL1MoG9Sg9Lsc6rR/6wfwda2TQOnO5zc5ugfbAVRQSTbUDk2zFXa2jG
5TPCaY8eStAnOlEj3D/RUeSk45iILXI9z2rzl49DV8tGTNjOHpe5+4NDKyerqr6d
eh/ABheWwZrutWBxW9H89oxQHlyo20iAD0cqOJVLjs1JY3/paiz7/mdemxZU9vYQ
bcQt+SN2EaNCKqSq+HIJE0dK6oMciItGPUyrbCp8DDmCuMvGtdpyjcOoy781PSPb
h9Mo6naNtBacY95RpV/zNScUD9ZxjUwpcw1q7zYxcVrxQ0K5Kq8dM5FivTG53wUG
zfKoLwnunDDiqYfV9VirA+B7t+qFvfJXcDDn52Eg+kvIJvGfvSWaXW6zMVvdTwbU
CgHGphx2Pv8F3WZ8BsjTf1ovIjpYWiAez5D5VgvX0TJ+LWPI0Q8N/nblUgAcWabW
pDtnYttQmcUfIpqgBpbVA6txVAVETuk6s4etFzJ+3QFFW4ByYIp9tI3p+vijC/gC
mnYpDwy+K98Rzb/SGDlAeZdRWBO1f2oZCMmPrrNhUb2oaBmDGG7KffrKIQP11ivb
OXsvuxEpZTE++eC6gHqlQukgPDQubCAlHrVdeu3kvfLzum5HADpgibxBCk5PWJ1L
ra0mRe/PlJR6a8CCU3iwrXg8K9TF2B6QfjhjJbExvFzd4L1cgioyshoY7MZvZAef
4AOOXnMZF3GGd6s8EzdsGahQBA+EcXxs6hdnOsyk8ddGaWQgt7Rlpbn733z7eGM1
5MMvbDHIHiSy5bYCUJyXBii6jxyPXx7ojkOfU1I9aHyQtKUJMATMlUcpiyeKMbc8
8kYSms9yo3A2RxlvxVFeIFO7/QNB+XDumMlCpQkkfP3Ah5xJv88H5Biz3gRRhjU/
D1Dbt2WaKKdUNfbc5i0G+GROrKKeAxUaI1wX6h+zEHuFUZWffSvmXy46LVeCWyEq
ZGAZkRnYtU6j8bosGh0HV3dQzfMM+yiXshOqA5+pnaAT/prLH+LO4ghzgaX/fL3r
IDzPBJ2gHmFMTzfvX6WIGv0ffXn90W8flUpRVvS9ILrye7THF6E1gD8vleAUSKFo
iCBidE4KYt8alDeZrXlGn8/CyH0ZSofvLer0ONAK042MPIHjisHkTq8iB+AH65rJ
fcnSA2ylQ3WbCiX12XQS2MC/1F+AZX1V0fGz72PR+BHXezaO7INZVuyHiF3Wxikj
HnZJV+Bb242WrBQYEFsoh3qX3gmbe2xBDCGMtfLHejF4F/6rTDS+bQnT2RMM2PgB
5gLVuPB99N8xo+tMtcSPxrAI1zZA0w0ZJJ5ir5m4UAvAuMUcGw+M6NLrJ8x1vz7g
LT7lQHnR6JqyAnVK7wCOVNbAaBpdz6db318kiLCYKP7I1Eus5U0Wq5R30OkZYplp
xHBeOewB9u6mtbcOnYssw0V7aP3+iEQHJ7iWG1X25jTYHRE0Nvc/Rm2+nEXMvS/9
soDAFYJDYGHb0R7Oz4yiljkwU8qtLxjHFN8UrtKDrY22mgG1h4b5hPGjOvnlhRzU
XledWzfa8BhRnN+gHMZy31byH2+P+nYH3i0K9IiPh1xJyLieEDjWIWj6LIpLOEaz
tGQJYMz3BJQkOQmDIs9/xVR64FQl8SSA8CAYXaFNj0ZTU53GeNs1PJ53ml24TEGx
pHoVIXGuOvUwPp4L23aawO1hQ6mUIuO1eh3qy0oOTV9hnirAIqFirx13rXACDYK6
pC4rh6kFAQMXCRviFbEsdd3ZCZiESEV9+fsKdmfHmqZ7lPAEmuw7/PBz9zlfrjHi
dqyoYima7qD+/HV5e+8BwwKeCJuP5jaYnms1mKWix9O9DaHqJda1YgGJMlTDuQKY
8ApBHbN2jT/IKCiOul5MA5x4z0DU1h8YZHT37PAgw29r1dNpG8CjgQB55OM9/K1u
w3QhjAgSoW3Yc0c1B9bDDz2ZKbDmR1STD/KimwdToJro5y634lCZLZ5N7SCOEqDW
hAZNEmcOqHlLPpncQKhOaAyhEyR+KrrweeaYIQqoin8x5g5pjBWeRBrb8dlORe5y
Z0Wv0Mcjw6MDcwTAxloxAnr0POLK/lbaZTShDDX5NGKfcz6MVpsuY/87luQWXKWp
MNFXXh6SNnvpdzbKchgrJ8CWB8v1fWoZc9HvwzA09pnOsd18P+L9ODQ28gHLc10I
keW9TXxo6IVAe17BXM8/LL7xPuZLRwudujGtEU7S11+2lU0d+wJyrWztpDah3naV
kxnfhXFTJKeCxmz7a7HMMBV2QVc5uetJeifdud0N7I+f5CUsysRwH3Jgl15Z1e2k
+oHC/XNBGIAPDR2j+sVNDyRuvDaCubtUBb2Nznl1HHJada66MjiuVmssqDP9x0AV
ag5enr4VRhUD43JOnERURxCRNUrPVlePmHDpqjV6Kc/LeDQX6U308Rc2rucXOqKh
++MOR9ZPSx+Zgds9DL71IbT8fupypo3bANq2EykLYkY0IKfnjbV0oFV0lkke6+hX
4BLph0DrkF2d1HZdD7Gpv1/sKj/OVSbSqausc6EzxdFoE4Zc5VL0rB9JJOBjzSMc
6FBKxAuDFOIQXV5JAkRJdmj9rLl7Vg7YAsMhjtNvcg37VyRwAqqIUSx3ymFNK6bf
nPLQWO9sIei77Z+XZyEtkVVJtsFBrdvQUpOw9Nus+gOmj+na9j1/eaonjB69l9T6
lRyEaJNFVbXAuMP6s+yLOUVLP5mw2hH2V6Mdd+Du9MfcCcUEGpOOvYglIQ37LWyG
1oDDUntV32Z1jBmW8vwaw0Pi5M4t+S/uv8T6Xku8A6IPnbXaY7+TLx8Xpyztv/RR
22UwHRBcl1ujpsBXYU7c5WWIM/4Ce3Ye3SjOwsSnu2Jmhe3xqeX/2JC/S6+pK7gU
Mwj7ijNdyHn+fnsf+GBgzF6Hc65Dm0Q0F5K4L2OFmwV55FWero7oNRKG3dJF1Y7y
7TrNVjplsg1qTdUlC8nk6k7YZTUutmYZchNJnxkr7ort3CI/LR//NagnnqIB5Szo
rRoXPMHv0fYuQT9wmeThwFPkJlXiNILtQf4/A2OhcDYE8cLBYg236xayZIlyAhHQ
s3/jUxUgXd/V6jCR3007lk3FMVQSuLGmJSXmZUi19duq77ptGUg7lXJIZzPTTS0B
hHEWWJ3baWbvR2fxS956DWBm1rrBTUWNnkyI2FJgkZBg1mNsuz+WTv9328LsvelF
HOie9h7Kr+kyt7U8ymVqGgNub2l8Y8OksfvJuy7eFjA35dVLI6JPu8ze+zB8WTks
UL80NFQ/1COSEwCnhcE345WbpyNnsncDmg7CCWnw8t52kFqwI3ljmfEmnTHUjNJe
z8gtbgz/xWPAHnNlTYiSkzjgLHgRxQaaymqHQfa+3NmRnQ0qiGGctrE22T49ZJtw
0iFc7HfJCJIaqMMCnhnjVByYhe+hbzCWnwAgjWzuhE3DssioneoqiguCNdCiSKnH
LDw+R+E2PhdoYLhSQPxNOBTvEDx7e5VFcIQmF0S7y/BDBvLe64P/tuZ2AmePCIyE
ueVxxOVRZ8Q9w1A4GZn/jDxbozKAow0yIDE5kKTtiFkL3nSsl2IKKXs5yv8iPHOa
dZqmjRh/5dUgFoFiOlGdGfSsvWDuVhOPsAiEqJAx3+uWcIXM3k28i2Elcdu1vJ5p
CuO2Be3qPqhl2e/vo7wmetSA+C1INAYopZEIDlOoeOz7fBzi4zUjYbSv21jlGQrV
w8PtMQaKTl8p8S2Ge+1j7D4NaHMnhjkzuQG1SFYjfJPreQecS5BLazAWa8dyz9mU
35zK4diyxKZnhBb1CT/No6Oea4tiDs/8SkaKStvWRxAthEgrJPxtdc0VIswGdr5M
1C9C3jZWTfK9uwLoDNpu00w32PydP40GAY6duAu3hvU6F4gTD6MgT2w4jhPMiTI9
cWDnGPckNJ9MuuCtwMB82LGFEoHhqpreW3t7BwuQUAG6hYcNNUiqZ8TRYE1KMtPv
zpO3ffgugFtFmPwUv40VOt4zIQK9jEWJDSXqCPqeHh6ePfzilQypzTdq5ZceWmPD
xn3+dHaYyYSUuw4uj8KNyZBvmhiFaVNRmsY4GJZCueQ+WaH9LxYv/hUYzMXbVOz+
tTmrM9PE7B3F2lhvKpScgGZrpyoHC6fpdp9t9M8fWiTUuWV+lzy+QwHY0P3IWFoY
Y1F3Mf8iYvOavx1Hw4nv9c0N3iG7UO7ZxYvD2yj+jh8nveaBowEbnj1rTR4p/slp
CNdRKnLOkQmeQ3eNCjQutZ8aumsEKPvReQ8dwKzMh75zse945bdlsVVC4S4mU9Wd
ir8u0DKtIF9diNElAHtHFb9roDrKJwMM8gwukx+L/AXlDO+oDiyZ1c24aj/euiJh
EHUp0FqI8y7yTmMTfzesYFuKkp7OBkwQX51fYUxb/ZYN+FcX7yS+EqqC74Ofwelr
RSk81j52zKdeYioXBSnQLWf4v9OlKduq7pnXyPyYZhgIWdHeAiRMn5rLqoB8bops
AIPCOaww3rIf0gdMpfzqKVcWcUmw+hjSlGvyBsMBms6fCEET6GdbvEEKq72voHEA
u/Uk/7AEKdRpqPBlw2qboT4i6scXBDdebK9+vVU7MKW3UguhelRql4T9QBWwqgRH
FKgjYHqpix9AMbU7Rtcd95CO1YViDtj/adIi+WGqwbCHlAewyiwt2YAW5c8l3hj9
LcKD+QuVXGqdkgWS7XxUWD/q9OY8v/CqS6C84z8tmQl2DRB4VJEbnooqUwIisjJ2
am5DDAfliOHptAjQbVQOouk/WIh7u3HZrf4rCPLAj7vEWpo28gV5IbJHpmztI0DY
Z4DNgK2jo+vP2PimqIbFMvSfA9lhl0S7osf2PAkwAdnccHeQdvADuiAbIRRDJBbH
Ixf8OIWzNfOD/I2GaLDp4OcM6fofBzHJ0jK+SMsAKZNvdyo+kMCbA2YQyYWTYsTy
+nUjUJN7jW/DsiKGfWB3zZM4K3UxF4EuyCg8JvKCxWmzl2su8BbUkhgaB4kJtvHL
soOfMEWp8mkrS5yo3BRxDGv1BMYdga/pwJhK3W06YKiYOB7BCYSdUyhfLpGSOnZW
7sqB97Ce/jwLZAgwhRL6O32d/BG11dPfM/Q9hPoTU3I0MWrfI2l0mwHsWbQivteC
zEP0igFDpn4tYRiKQjUcuZDnUAx9YHMmjEh1cIQdDlGMcfgWpE6Bpz0CE3qN4a96
ohaA5ei+q5JFtr9pbkczEvnNgSj5DhWYlz0NdGGZlDsNMTfu8+M0xWy2/RIazzAq
iAyVcMruDEPRlIS869ClTQn47Yc4fbPMFauaCWgqrVcPgE1WPF9HO+Uxg4tUof9N
S0eWv24XLpReumViOIxcPxq6xv/Ru9ktAJK5Bsp4lqMV7na/vhtFggW0ivaMD7FW
uqmoAJt7ZolEaf1aok4JDrqD6Ctz3Lhs3CE76/UvQMBhVpz0gCaRlDLfueGpelHA
TUyi6yR2HueWpntGDaFeqZ9WlYYkNBCk93C/tLa10cKs3Nn5qzieSQbF8cnrpUbo
8vUoWjP1Lurcj2qoPfXHGmRPvCkdfjd1eooMEidiiz5Yfbzz7um1Umn3+522hODq
s/vv0YMAH6Mk0on9kBU9zweJ3fmuTt/oIMhx9feAzQtxMFzHGsN+/TPUma5DozFH
JuU2J4R2v09RuZE3bPMkGSNARd2TM6hlV/qt8t6HbdjkAcQkc57FX2wTRrUTdvj/
4d2V99k6VC0F5FsnTAB0XLEdcZh0q0/hiwMTTL9J4Qe5Q1ctZrqaO9JZP89CTJ+Q
adPnTojowjsyefU5MYAPbEr/dX7QkHDxDph03yplJwxYqIu0e6cjLiwH7AvrNhYW
XiLenE7Q/RjjjVCiHs4sZNtytU/TYlH9HpXQ3HDpy+DqJKBISRfrKYw34bNg0uQv
XQ4P+LpW2PH2YqIfvJoSNSB1j4zv/hKy7GOOPwjCiu8QLW3wFEnfqR0iAEo9HPLA
/CDTIHAKB/WS/BeJTGoCboTE95Tww3OIP9oOJAdbZQBp6Q7weKRcVgm65M8QoFF8
yq7u+VvzND0P0iogGP/agSkIi2u8GU9CjFJTs4A2jPpx6ewXFhLmt7LaeRDHNhpW
7MI5XwtRsl/Dd+srA9CEOtid7A10cuYJlZQD3M7iD9CMQU6AvZW1wZlnGoMYoXYJ
OU//zz/yhTPDEnhBY6gqrKICp6du4d2jGQqFGdHKyWYdbVhLfBvU/kM8pOL+aK11
UggpQQv4uA5t9dEbTgJx4qb7bGf1yJDGzlzhHWrUzd9Ke+Ds0XxI5Bv6fR5ABRjK
eSfXwFFcMxkNk8ULuZklmAIywLCMQMlymx9c6CHJsIvQV0id9mFeHsl5LpRl0CXQ
ynefaRD61pj5A2FaHtfS/gKX9SoYY7KiFdQwXIp8FAiX/mnLKXE14Vyb3S1FIJJz
GaytBErjsfgR3RbZdi/HqD82n+0byfF65AFsv6U/4cHbtgh0AWOsAgA/TS8VQ6NX
EtO6i+GhLGhDbGV+Az/ASp7ocuDgEXzvi0H9JkUMmshQvOOPAShQv73Qq7W8Df4Y
iXRO3r7uNp32OjkTNMR49G4oGIVCLwDvhsV8eGw0IT21BM/uxOIeZd0Ac6xzrIX2
W4REvRUzjQsXVV7zTdrL1XnWvKNZ+QrXH4VuevdJungtwqE2L7Ptc7G14l4h40Wk
WI315IUH0SU0t0l/veIU24xwO2PIaM6LhKYikTEY/2VbI5hwQgZXL+U1fOs68xT9
+LXNxfpud9n4CDjuUS7UOQutc8ID/Qb3/PYmgpCTTT0tdFNFZRinMy7P6XijA9zh
zi6QhdofesBmIQgVw1/L2RiHG0XpuQNnFsiZetyjwu4qMM6lRMxrr2A07khj7LWf
oHewUMYdJAqaTs7Hwz/FLedO1cgGW39X2977n+mG+H16uMJ3DAOAtZq4RX9MH7Pf
hWUC9rKLgGlSbuVKMoNI4MAl2w9lHgEIX7oCl9d7FQYjfrZ4JLAsSnPl4P6a5de7
PgBZeNjh47u+y15kRjL9UMgckiDXVHv5BEir9m4ji64z6oJkUYXzzymxLQbdNwhQ
0QdE+oUEraB9VuqCS+zKXPcxfbjCJ7wvQKRlJj4ajA94Lw+yf/gis5FMFIyaOHCx
K8aN7RHDWDTI79AGsbctHrdlvMJ984tPcl8WT4T5XF03WO74/I/LyrxrQwhPqSMt
aEB0Eyb5BMK/Yn4elLpzoTdHuTsPifascTOfpw1L8KRetksEzOHarxNkbEOE1A3T
yjVNWid96HpCTUgKXk0Wk8OWMp314cb/PboJ/r22HPsy1UKpR6Qad8eCgmC+ZJ6e
qYIXNi1/xK9IBy0GR+wqbnFpex8Gi/YGgdii+2ZeTUyT/Y2QG3mOfljYiM5jFg45
f7RW5Uzq+okTcTTV3Z6awnjGVhFG+U2o3eMxTr0apaRlk2XEwqozkRTloaOJvhMp
laTtRhnJ8x6Qs8vCXmbFO5RYy6eh3XRAkmoi23D30Mp990XvcEoWl/gFj0UjSFjX
6AC1Lh6unf9znHn0TLyMXbf6nGxd2q6ATlK/mk7gspecNtr6aOI7LcHWOBih8Ijl
zoEO6ktmumkT9briA0L2XENJAJXN1fkg34Jo4gauCAMlQT9JsV8X0DIcP67/tK5U
PhrXrnTR4QfnNqYfmGgFpr6Vxq2xbFJV9P0p7JU+CF4hgGY+mneXTH2iIzjUyu9p
r81BkyzTbyDXCk/bIgQzgkEM4IPK5TeuRaS1sKYf+E3QBY3eGigE5q1xJrYwAz3o
FYiiGCJX396lMY81Cj9HmqW4s+oMeZD/9Yh342xmLPW34fdxe+ZlFRcj7/QpxBTW
IO3+6x5+azi+Wm4Q8tQjht8QD+dtihBJQTIXY0pIMlXh1gQf8pYZuHBXCaQ2LnIx
phkP+FfxOkF6WOEJWZ9uG7Nqebs741ZENKFyMvs7CthSR++701TDchNaDjI4yxe2
F35wZDGVcwzHChfzFaCGUt7EaPjpsTxQTqebiUCEHWks0A1dyNw6wPh5L9JQQWF2
ZCZqo8vHsSAz4YSn/6VqfTBGYHVzbWaEVGfYY9OeLRuTAJU3hdWXF0DBqoxJMVIe
Bb4uA674zf+xLyFO+EVaQ8TvWT1t4sif3kV02qTkiu9KFUVCFODcq/oq6PLioRDu
b5BojXbgDbZ+QOsd0ccYJt2yH7YaFnRz96m60IwbK8ZniSMvriE3HI5kYxhxUdzd
N9+AJzI+np6Of5uLkxkZE5tLzPlLxTh13/onBvyOciF7MAVJJaKFJtqONsr1Omal
yd2+6oAxgItiMluUj3iOftgKEsC3V7OEoQ0lFrTJqz+cRxlthdYoLn3BRHHzZdSA
hPUeTZFX7CX9/68v21MMkmA9RUIZEBXE945dyl/2dXZ+VSqny/wQf+roxEeU4bQ2
wYpG60L6RgG3c0PR+3vUtM9xLXkww+HkVVcxnLCJTz5Umg+ZrXtfPsm/VqqxdNKt
nEqGV+B5ZcIDo4WQ4qoyHQd9blWSdvQrLv4XQTKAXtcr0DZjHcJwRqBT/1wF8Zg2
07zy+TSEDjn1RsrSKUTBkMVstVJTMx7xjCSUvi/IGfDIO5LFHos9z49fftXiNIs5
hTcqME5EZ4/FxDJnjW1GJ83UsoICiHng3+MF/srL7SRARaZ5p+v96o+H1U7ciVWU
A7WvLDYR/3/mqNmlpon4oxLgIRgiMRj7PBykDKNPGELMWNsbotqvr9USkCgL56RF
rr8BEOBskaCZ4V0IlqanugMUamHqXo9gm6lKQePaCEYdlJ8PBNfsUWAGe+XNzjSV
cCFx/FoO/CdjvMmlSztfBc+A6CUbtca0rzd0/JTncNHp8tsze8CFSH9q3fh3zr8d
jKswi1NT6U8w4IkiICXQj/THc3UMvGY0YYNT8wSahSVRIunbT1v0ju+ge5SPODiN
vUdHgbnLE0VpHXiA0+fBinw5q3Inc52p1qMZtQmoRBDuaJ3Le0AGiHvlhF3Qw26v
RD88Bj4ogY4Egvy0PqfaHuB2/XuzOxBuzC8lobzAFLIiM8PGkp6RaODiWtWl50rx
vmlqzG/ZK1U/Kd/bii6zBSXaB/ZZ0Xzeanys70ZVoXY1GFvfpZroH30QR0IZW8hq
2KN+z3CnBwlb3LZT2Yhs527h3KLlpwE7NJVQWvq0fX7/rn7/C+ltXeXDbgQZ/Kwp
8GYGuKrIxeHrRv2uK62+Y2vb7Kgw3oB48xq+3kqgSVfYAUlVSG0Ie/fSUV3XI5/C
vSaDtKF+LWzeO/KpKBNIRDhtYt2RLHN3ZwKxgRalw1+ak8KRHgLtHlP/xUBzj8GK
fMcqyzW68jkuPFr1gId8YaQ39eF2cJp+p6YXaTpLpPMRxdaPtFUlf2kBNYZxe2wD
IZ192UTjVUWPmwDXyll3fyX3Ot35gLhlbavqQ2/Z3AqQByc1gm+fU5lofYWFvovl
9gNVfg/JjFlPH1JDSEQMk50fo3+fSH1mJafcMOYv90UPqawYghDD2jCYdzJbkgey
mp1/PCzCaxZdZ0axrmvsZjO70q4SiIs6Hdy79dn37SW9p/OKVAFDH/j39TDjQSyy
pkmR1z42TyznmLhWfYqnrOWKPvR1cxNRtvpgdqUPZVyJb9BSUqTZGdv2uZ8Hyrua
PaPt68c3d0HwzZLl819aFP0qWgWwd1LU1/9Zny6cfO/8ie6nM/6EyV4hlfXZCAhD
JR3BAGmErZN+ZVsM4qSYQhYYKbyXjz8ZzjobPE6e/OtWup3i+jQFcBTTG2R5kZI0
wWKR+r9iHnIrHmxMI4LkYL1sEaNJOH/pRb74OVt/kFgvut6uzMp1UINIkp9P/9At
Tdykr60h9MXbsgn62nRlPLYVVOAR+IL7fesytsdGvP0Dt6LPnfxmrhffoK1PPPF7
AgLDE8Yy81emy42tI/la6EN6GlB4vMbgvgW4mk9tXe8/pCkZRBy6+b7VNuPT9tqL
mm0kdJLPtBFdEdfhgQ7bZOVo6tHZam3gB9FkavIh8eSQ7qi4IbvQ1TEM2krz/a5l
fhV6cEci3KLEqmjt+AH5tDx0xPk/ZZj2DQNHZEYMz2IMr+sglRDnAu5vJTbQoNph
/aV2P8Ma8EwcqZZqN0O2GxS2NFa2snrj9rPIyiTHqUyGqwbE/KCJ8FLiNGFUcisJ
LoZbl7Oyl5T9k2GzWLoOjs6i2ASdy29/Y4FEfJ2cIy48/rjI4nvuVNei34939Atl
VwBdnkjp1pOUYYkpD01j8lo+iYtAbLMdxXbaUiQZyhWDJS6pjHWoGKLI/IjVCB7W
O1/K79ZnBr0bMj7zOgqAZj3LS1bKjsgKcTz3L5lRRyxyY7ti8J4uR/Fw5dzmYybf
WztLtKWq5+FQUTBSs5oFEloZ340LdQbu3W5+JKdkCR37FfrLJHvpWeWvbD5nJe/k
N84Jw9NLn3Lp4J4Ef8HVwc53BNCiR9anSnzooJt8IA+c3iusplZwy3E5JnmeMDA7
fM1TFRYwmYfNqv0519nbiJWoU4wUk7teZQnfrEsBeJLCmsOtknRG4no9NHodRg9V
MV0JayT1ekqNNVKKY0ByDwLuc76oe6FiAAGsYLUl1pV/g0arGq0k7GUGTPU8hurE
gXJp8wKuh061uMHu3xGyfDgv01UxRqAdL94CsjFNNW8Po4kA2rCgftrZiZt30qQU
wwUMzOxGvjQb0Zd7hEOn+uoAfrmoqGBNqpy86VsY8JSQAw00B5IlWpOZgjFGtai9
aXnvAAe7+sKJa3tdfFl8oTlLvmJLTcpHnyocEsegwieWHlOhga2LNYGiATl0Erfs
FHB83sbwA3vBTKtnvv6AABiyiTmR6b4W18RBw7X1naXBR8apb9eYKgjH3HNFuvoE
Bx8uupjybjeiSqUKHckKvORN9Sn3UwLKIyCzMYi/cFtL/7zwQbluZLPSQAL38GBA
ivHEW7iVTARMBg/qNefe/g1RJwMORlDMLu3vUPeN+ivHiDDihGfe1oNuIaxoNwh8
0z/IPah++yy19T6jOp2R0xvfp678FA1l/e+mXFtsYYH8j8wQb6MGoJXfvoPijLag
bW3TImkm8CUNoIGXbhIXigUoTckbV7rmtLuHzB1SPdq6GuVw4u+Om86gQy1OSMow
SzlfXLje1alqr+pXUbwYXQGRUyxqYQLaOOI+seINOVuSUpVZVUm00D4wji/M3024
t3FM9sS/7w2HDzMX2fi27ZsGKrzbhT3AGeTgY/emCblSoQSLyFAFA5qQogtg2pyy
OTYOR6kvO8SM/nRcF0eSc01L5N1i6T5lebXd6gVl2g7+u1dLM4rvVUZqgTFGWc6y
DL5fBdB3pj20rl782dV06KRsS9joEXw8vY7Rz1yTrpjrdU5TyZgfvFZZNH6jbW/G
x0X/mUMRGQdbgPOLTwTJ9gAyXXFDrwPI9nAdBN5D2hBUxX9uYTzPSAM2xKba9C1k
2QXHBeC2WiZn4FdxEUqSqso2kGe9NX+HFxd32c9q78VYBmUefhVQWrTRZzDhRr5Q
xsmPvMw0OwARThVg3RSIqtmjYQZhm2XRP0k9WHDkldXZ86h0/+loa/SF/sxJ496Z
bSdxcepSuGdfkwW5xCopmOZlF+dzeugIVdVwWtl1s9MxA4YZ/YLQ0HwgmaWs3MnK
uZ4jHQ0hBZntq9EAwFX0dkYOzyn0GmXEv6ZqYYO9nzSU245kdu337TCrZOrVlt6e
/q7nAz6aKB5oNPanpVRE3bm2xtiKq7utjtpT/IiBV2cSIaacuz/VbD1zt9BfY1Yd
EAMHUzl4EHJtivpXXjhTFbBtEL9pXqPBbjCSLsJRMuESrcOu9bgnqjhYtDYfRP1T
8rWoUFCzTLtyvz3JwaaEYZ5ExPx3Ywbv9NiYcBsBnUTWmDrZhM6KlODh6L8ivqm2
XGT6IHAQqVnotxkrmEKrb3axz8YImn8JoPhtx48XVKsEiDo0iBfEkdxstyjfHk7y
nFa/UjKOK0eBh6N23O3xu7ZnIhzgMgXs1+qHONzE8FNOspOF5tpg+F5X+VOm6/bL
uXHSQfEeVl7UZ8LZjHDk5uyKm93hqUO7M4E/LHUofjYbnZ+MRZ43YOZsXJFFrYLj
AaLAvEk1DT62iz5OJTg5KVB+RzdPlAnsIyK9sdxhJALhEgN9hzT70d+UZ0y72t8t
vUq8IyNrfsvT6vFfOaMkQyt6r+VVye7V7oQNq9T3XQKtlZwKuGdy4LJ6zRvw5zxb
Ty/dFo8YDjDEgKvWEQm1aJ9Hy3dvrlsmNOR3n38XRFt0l0iJ26RzXzLQSMYFr7zd
wZCu3melQgS1lEhiBj5ABYinM7mbp/EGQykS0S0To5zjFhALpO29/Zh+Nyy4W3oh
cPtsM1ajyfBs/gqnJQihuL4NNFQR0rLpFS0jaat0FDSU8KvWlnEAe93xn/7oP2kG
5rs+4GtlKCD6MExlY4dTwcY79Y5JIFoQq9ENr4K+gSkZGQ3l7yUoS/AMwgiIg0Sk
hC3kulwEcrt0TKnqLseLwvYNstJ700jsZqnLGc1/xC8yB/w0erh5cgXopv/7CgXq
YUTWeWxrSI4XgvR6tmuHXBc/kJEcq9o9M1TNQwdHo0MnYU3CK9Lk1htDiNb4t0FY
mnPBdY+1Pez5mp1G9gwOLfsOIfHA2jJIdpuAvKJDkbfq+AMZL07tkHJtgRsNqEGO
G0ykvTjZjynnyp92Uu7egZBLNA7aLVnkfBKk0fyv7MUjszXauyxaPCQ7+7gvjvKO
Mj2EZAYOSM+IUgdhCxniiTz52Uv6f1I3eaNHcUXufxerldA8J650mPqgoD2Z3dta
7iC5w6EQVndFQblN0hzmOVDblPuiwNYdzPmazzZ9MxT8x8y3RkUcSfaS+xFTL+vZ
RtGkSVjDQ+DbtgfKlPsvW2MXZLYOGwad+RGXBkhk9Z4aPzloi8LWyC/O2ytAyK6d
R8bPMfOxwgf5YxnRrdBMHOvX3ijcGcvWr8ZmDmKxso5ClfCRrbvUiuA1h2Jl6uVg
Y0JeQvTV4b6A9Aea0+9daWlTkyFHlklwLbLziezqXfysxHsUeCTAsupldvfITUOu
jHBQr4IYeBUC+VNa3e0Lb7uflNycbEdOELhpjuDVvgQgZpovLUaDN3weEk/7VB35
HeKFe8/Xr+tLHVXwJKZbZqqLI4jo+G7WiKR+eKL/6NzS15uF5n7X2OgpQqtzM9VF
cFvFC0qJ2lK61MkxLco6QB8OavnWYDsnpfOYcmmy53D76sqfRKgptWrKkvg2Yr8N
RF1V6j55CqMBD04peDD7mCTifUTATe2UZAiZvkwUF9pk12yvJcv58QO8gLFFIYEF
aGggL5u/H/lumO57BNfbAY3rvizOUATwETdxtcJkrYBOfLohk25bwKsr0qyYHc3q
zGlTmAq/VbNtBl2tdTvVrrVyiXy1Q09GxUY99F13WDVcRjL4sBSUTEpSZrtmnShL
yb2Ts69g/tjN1thr8mQxssa6VMwhtfZtGfC+BnfPWCmNst8X+LM6ZGX5iz0CCGLA
R6Dz+pYmvnBpDfTemAjMImR9U3pTFesBtDphsOSyyC0ZMVjGJhpSdxcW02RUQOKp
bparak4suQPMj1bDJgCIrXmlNGG4f0nSqMMkeKeimpK6Uww800exEvgEzOrYx74f
MsnTOdLTLc6lsUNi4gghcMbhlTXVYxXWO77yvAxuSYAbeNy8SCnM6CUVaErx7h8E
7I7wuktAcRKsEg9qG4bhwGnhR53+DzzQMPCmwzh2d3X9KKiIO/Khw/W/Z+l+gNOt
g+UU9/4Z4XFaV8WBtcqKLRh/W5IBVww5RKYgDoWM6xOjs8SgKFz0NSVaNTqwvv7f
weLR4srtFVWmKJ7g/9vZGaTP/wNL8uaVGyqafvoXeFfyoTrvsqRmF02mTIJSTbho
rFdD2SFNmeOwETwcW8Yc74bKRH+ivAex5KCEOEH+6DjiNRfPRBVB1wvLAFgJNpqH
2s5ySdD44uyhoMKigi2lUmyXgEgUDLgcVaiYowkP4UUAcKtbPxzWKa+T6HJvCdyh
JGxLYA1w6SdTV9bLLdXzF2RfFxXsm/tzp3tFGT/+UijCqwaIHQMvyFh2N3G/Tb5T
rxqZvQ6wL5aa+Dd+PX1n3O7txRM+A2wF1mTVI/wXjyyOMo1sf1fmCZ3VZkJdtjmG
znIydfBKgpcNeMg90vslvuw68AGvsM16uZG8ODeq6lzlSqvCdiYRqfcZt7LGhMSu
/fA45KWjwgeTBXZKNLMB041kC/I50xffYsNge7MJ5nA5lJqHYq5j1WCE2KWJZklu
9kDQLuukdV+ElVvOktHITn2PwoLVXuA8rmWUTyPAbx0bP3hR0JFByzfhLT11QL+C
/2Ph9jxsbqw0Ewt30pid5ILyzMy7KBxxVfmVu7rmBqROWES8sXDSCbj2SIwnW+UK
8iDKuda08NKKsyNpY8+T82LOb3b2pwbfdzjTlro99peq5pK3cTgqdFGAeMGJ61Wu
p8ojNIRJLAgZWWLMxqXKP6d5CGUS4J268LGt/I+7kL3aI22FS6tFZNzcMSlSePpy
lruInD7tWNrsyeLnyv9bjpLWkuyEnnrJs54JQ4dUUyRTeWIHq/8gkXJY83rSmo4q
csaj7mKqr93bsphO/CW65EpG+YBRUbQ4PcZ0uns03hJ7AghlK99DBpQ4B4CdIggd
6z1XNSiIt5f/wtBgyxubVgwadHHdPo1ONpEacK8nmJtAPZqcesiYMVx4fC4i+T3A
fMSNg5TPT8B1ydOU7m/oVTVoA4oPcHY4TStdF1mXLEBtO4eYHR4GCEmAo3/Qk8zM
SpXzgDEiN0mCO3Zh4VnL48nb6GLNYVWzPRPNGYbo8CDGgcnN39Bd+P8NtTH9WHl/
lPV9GEMPUMunRdQ78WTBwqNgxrMrlW5eXHiSbjwLQNv5XVLtYQDp4b5TeEpR8+Zd
ld3wxuATdYLDEIC0dXG7u2mIPRd+8/XZBvfqqByKK6ngZowkHYthADa07gVAAAD6
sDS/5U/6mI33QKnlV8GflJAWcUy8vm6ep6mcWAlzH43VRMZvCqhemU11hay3/NQW
oSUPanpQfx5AM3fED7raDKXYuxVejjVmQZ0SCf6KRGb8+t1LNJ78DZ6VFbozyB6z
TWfViW6Dy53/C75EsVndTO97Egx/T3AYExDs0sISXJ3fhaSscKYs3waTxTKeMXcu
02Jz2FgPPErCRHCAeoKy6vcJY8EUo/v01GaZeZE8zA+a6d2iI2vmvKjSQvAMJ9zX
zV/O3Bc3jnWK/INvvNvJeF5oS4ZuX7/NLu/EuMjTcMCej0fJPbcKoglFEj417T37
CU81UwxcqG4Y+zdwxrFcacMGrteeDWboafHiafjwqxt8XeoNPWHSNZ6GlhEKVsrG
MXBoJZlVORtfVkkVvywBnHr9YAKVUjsID8i5/sEwY2RmHvUcz9l4Oj/SRQm0Yihn
uiv7l2dGUBIlTO5sDWy2MLUQFDhh9cbgsAYHna5hRoBFqmvPefCTf0I+UIr2xRAN
BUrfAQyxiLjw8gtj3hRA76i09L61sO63YjG1S6frdoJryone3x9VaQFIPCgVgvo1
azDABxLq4ryMbdjHar98oXThQTAb13MjP2fPzqvgg5Af5jCpC/Pesr3P76J5aHyx
sl70QSQc7DAbwfjMkBJAeB6JdCAZf3AWR9iSiThIQWStBlZFQGxK1BQ5jM2sDBqM
pE+jr69A4R4XhfkOFpO7JMumbbSDfOLwlqYA2QhEyyMZ3gCwU5JxTnyATMf5emgI
efsD6crQtsyToAaLrkNDBan7niVtalhZESdgWFQS8ggPzrSy7llykQNMN8F4E9xO
j/9NGTstYyveVnO9h+/6jZ0/l94i1xJTQim0Gt6w5oJU09RzWr9PMupDohBgGnQ7
3iZQqfis4xZ+874oi7ia0OP0Y0QBh/aRNX/Q96UcodKgdG/6yo46TOYBYzwUzN9n
cLQptwqcjsJDb5/n1QndQPwwyu+Jp1Fo6a9aIEtVYXEcN3LAg6RwqzW3R+QfxLWq
LlavyXfvTnm6X2Cvag06cBsKMhmZ1SRz4gjhcN5mZUw4BHUCyTy+BZ5yIi/IYmgt
4Mvy9tTZyO8GCYtaXv5OTynLXg4ZG1FwcBsxizLVgCQmt32Ix8HMAS8gwZzrXuEz
UqVHgu8t/rpoa4ucAXJUEdWoS1liNDKQdBdzVCgZBDXASnu5sDP3jHSgeGdfKh2H
oraH27xdFlYvlZNnQ5+QGD78awNuCyKqNcFKSC9zeM6njkQsSIIq9rO3odsZl+5K
yK+6KJQFyDV5T0S6ph91PnklSwVIpRaZ73d2bSS5J7h5Meo/XEr3Q0FUioYhc+q6
bZ+1yPBOXlLeq1VpVDriJ9v5pCdCjpT9sT6cZ+R7iG3avg33g3I363PF5s395AJF
4H3sKBQhNXejN53P0GGZhlgrdowSXxheNLz8jZUw3tgoAD/IrQ6K81XaP63gMajY
cropKbEhybasmJmqQM1+LZcGUhQL8quSJmvQhQsJGiY41Nfn+hh1HQU9bhbvZPg9
2kwUtLuC4XeKxOluOMFhhxhBpGMbz+FV9Y5qLPD6BFIIuZu/PryK0E2KoGhLj6wt
5OEVCvAZXCnQQMcGUV0YI026lihd3fHDyvDwoGrwiBzwWZXfO+XGBYqpWjfblor2
GRvWoDeBTbKWo2YgqjQJcF3/fj5SBATR67lqmofWCY7HBmLme1sdWCCLGBnFIm2O
51TjnhFISn9T8enfkhATBK7oSoGKWuF8kP/CuPTF5gmKL+NRzb5LpT/FnxJM6Y/g
ZJBQo56XRfbfVoqPu4gTtr7vI+4Ro/8QfYxd7ytBR2LLcjkM7f29XzyMto6P2yWv
iyWR2wXRwRw8LIgfxCTSpAxjSJxa4lXSPoMBOBoZAUgqzshKqwsSEw0tqZDZyMA3
X5KK1QUlUMQHuDQpY85rt2EazBcyNY4N4bkby+47mFABp004bInP1TxO/ggXeThi
sHoqvpXghZWY33a4lcXR8ZyMrRmKmUbtqtBk3Dcb5f0IwOy1sUJGwA6w7vnfTOus
QSza8PYWI5skXstjshTYKrcI/HXyjr7ROrhjKLbGUAtuJ/xxbr49xeX+nwc+JKlM
jgZ6BytJuBWr1d6Fc/tQKm/RUYejp4sy2rm3qkd7ZZrPJD3gnXtSGAg27GtMzW4j
X6X9vdKDmb9R6B4Q494vAhROee8M02G2+VUVmauUJa1Re0KL2P/SS7vpWjIGcz8h
/r7oSRW2pDLwx4n5uwyOVOTmKg19xus/MoNEafqwG/IMtl9MN91s2eq87B0uTB/5
Df+uwq9nedRR0vLGV0xK8ug1XHWEqvi7hQ6NmqMS5DR+ngcNk2Ch0DTgpeVgC7CW
272k4AWwNRa+ahnTDQ8u/7SSaYAQ+KcXzASJqnybE3/qFvJ667tE4OedIOiSGL8a
nodRnYMTQvl6jIT48NzP3vusJccC2b/AeswYwRRZkFo/DvmZ+7kRM5pTWQgsM3gv
M/MOgmAlkrdTQhBXvlqQEFk6jw2ncHDfQImOj98qxLFNxkru9qyCYPBCV9KQifQI
uhrY8tvyE9mSA9/eRZkTtgUnXXW3tT7/4mkUrivxTAcr9yFsCd4VWkiDuj3JHu+i
jlu6ZcpvcR7SeFfR5ddDJYU2POTvDMRXTIzbmUVMiH625ATdaTCFGXLWjtWViunz
aUIQtnT3bI1EBpFYTU7ZbSx1uV+2PWOT4CKqk1+0D6P2FHC9F+s96NSUF/oznlFx
VsF7syxUaazYdSpAXAazO3b9otS0fKYcOXf5O52NWuMl16RNLyUP04AIBlCrEphU
HTOxmtI+/RYcrftf+CvaMnSVl+BlXyJDhFQbidx64+/bnKyKzYIJJKnxPdLtgAxS
Id6O+6spylXPgmirexgodMDgmnDs4oCZkkodBImxgW5vetYQjxzJWLP41N2L1Usd
qY3oWCfzleL3nNdxl2vpjvcisi/afBKqk3WfLxKbWZUZBFUCjR+LPspaebSjZ4FC
8RubehmoHnHI0flB8BGhqQME93d1URtKmhX4qjZnldFOC94iVIOw9VXhOPDqYI4Z
uUGtxTnHazcrxg/PNOaplufKjtlF1Ri1PkJEWY7Sy8dh87OpS6/AWgZ6SSlnJz1s
pPD0hk8Qx8PcPmosd0gtcMFUnATB41ndrauK53XChf9c0c8hDr4MLbOQdngkwSe9
kdpvDJbKA6/+sDWduo00+tItxmJWclvtb8+XtvdwIgPdWOkVxUJleamg9aZIPdjX
uuYwENGSm4jiEz4B2pNMx0Cl9+/ikxZFGPLz+j1jJhrRK47SGlY4Em/qsHYkq5gc
30fCYvkWpHz5s6yV3AvDmh3NDLkvu0KGZJ0mg5zPdSIJAjj2BK505Y8Se0avFLr+
ph32r0ywFht8YlA5iy9B0rTDDAm8Q41txryLThvbxRrKyh22PrDSo6njJdXmOH6t
xHRqxSN/xBabFCRV1tpwvH+hbY3dUGZHFnGFirIAoP+wb9lU0kp36xBFoYyibciZ
46GWyjt1Flf3OdRVdPYrAhsW315kuFngOo7BJFfuDmk7eRNfjwbrAAdNKWrBiaxD
lZD/B1F0pJKc8dmT/71QggCgw2Rqr90FzTN7kgueLGxpfzzCoRKzwKBC6U0VcRaQ
j0nzh0p09Abpi3I1fK/R817Vo/E4pBtl5HFyT7zfob3ZEBjV9Y7j2G0/E+j/yaC4
GOTQIG3FyxhujpK+ZmzZ/fVQHjV43PRBh+e8whJt+tkVmfbOBHWXnjR/oh1SmWme
5j4tng3kfADj83RL2GgM9Fl83DgCw6bApuEpcugXPYM+FJQMCJRPSWfeEJZd3v8o
m97T5UKtxFQoIS58J+1PYg+b6NFgHNPq0izCbzqcC9Eei8Jq3HBOCaQMmMxRK5li
KvleqoVsTIqtywq08kiq2ZZFlimWw1miv7qGkVh4/Gp+RkCpCNfATJeaqYcJvfm8
h6f07OtZeSV5PPXMO9TqbOTKI8Hyw1YwZAGZZ9UnAC4a3UMhYFgYjaBbUBnkle3L
HQAgaKkDqYxADJRvZjvVy5wbR8oMQkNs+e1DVr1SMXwDSf02KyslSXHXc1U9iQV8
lvtI9+L0gGTS4P1BrdC4qrx7mkR1wgA1g6TabKrJxZJnS2Har47oCoruTVoiHBq4
Cr3XXVT+5A2c693vfOi6rS2//6q3VWAEDqw2FyOryDzsm4FGpsVgUgfhjzwCkPrN
bqsjJdwV9mxzGX/MQjXzFzAF0G6qqPGk8kGJozkgzqrYtSBf2nlJOnLxGGNNUXZc
xGYqPbPuukIJHjSPUV6Ljk0NF3j+70wiLFdQzt0xe0rmXU2ffGWlC/j5L5r0rdDi
njt5d3Sms6AuFBuBoEgsMaQoFTBD0mDFf01bvufpjymrrW3borqRUeG82hFck+q6
ScqSW0B594luFHWz1jyXLR4SwdahJKlv0R/7SCS4qXbvu3fLBf6alQoRHbKtJSZK
WpXOq6WR8wv1LuqVJC+8oL17qJCnaXT0Ac+UDZ6R9d5L1JCw2ulBsFAWfw8RU9YS
u1ILjGaOvYlUob0zQ2yFgfLk9QhQIg7evCZRsOpR4POJveNpBtYNpoHPkSncmlcn
lrvga4YRBMi66Xa0ufhqkNZBjTTRPkoFGvizJHr82uB9itRaumB5ERXcT7ltMeRc
4DD6PW1EOVoImr+XwQc8s5ro1lHOkGB8TXsoDfoomgY4Vj3M+RLUrCsQj87N39mJ
7FITLyS2PhwY9Yg0Unef0cjofsrR4u8B3K79CV7VaK0LgkvbVaOh7Cha9dyG2gGd
858LLQKwKzbDfqV26ilEbkldMoWPLmjrUX+5H18ZelSOv2LvbRdXtw1zEPF/kMpt
0y77x9uaN+jiimxUYikNwA7g4n9PVAUk778fjqJXXNxcDGuDmtJm7Ea1FG86uJQS
53wE4zD/ktnn1B1lPb0GBFPxeNWbUBGOTjoi8VSph+euYozGmSf0kmZp/5AVZ4g3
vsmO1kMYUK5lrpToURIG2JJaXoxmiN/Z16XIWm9d0u4ZEV5VIJOESNTNn33YLu6H
+ThOqhp23xJNbA7ZACv1KnT36Pjy+5xVlxG6Xk7bOArnGQJrpv2icaaQxnaELKLd
8nbUKLeJoX03Z1TAaU/+hoEwVkdHKuH+pK9aYrgG7MeSHjW9bzfWx5NrWViyXVID
0ZwOsyWeWATyUBLhZQqYiCucvbd1yMxivR+iLVzsaiTECXkUQS6/Plo2XNtzbWn5
2qEmsnQI1Mp1UwdOmLQb5vyX9cLreRBixUmsfbM74BB9+IY1ZNlDv/uCocdDlAFp
G3XlTyPu/4vFZ+56PK2ejqY/ucAGqcPsfBJyfYwmqKD0N6XXNvuiww3402FqJZUi
4u5oBw19KV6lku/vVQpttzGa5NPBDvNXSsAcY6fMu2mbgRqE4KX+EJzHTcuBnF1n
5FPQZJoHlE8eFRA2op6oEUfBQFA8egtBFRqjb6x43MiSaMhPhK2gqAn1mZwuxDib
sTJQsEVV0wFjMFjCU3qqGBjZQCgOIzgZQnGlo8CTd2nALgs0Ttg+ccUPSlEkuMuQ
L9Qfy8aTZ3/utNpdYdwjplR7o2+aXVxWBLNtj8u/tdTItGiefT8wyVLTga7qytdz
Rkv7ODWmGL4BW8BvnZLgLETPBnG7DU7vrefaFzmFSq8mnqiBes0vjdVQHTwclw95
5aTF/wh+eCcBMctFNisE/J887hOQQdg8KFY3QfXEvQX57lu2c/MoPOWelxXsOHP1
bisE8SbMintOF4qcxmfX3d0Z7SdU5pTZcZ7sOFL5QJsk9fjb8yXjxAkectN8nXYM
sIQcz72Dhl9NkhPI0KTceuGXdhRCw3pgoDMuA3byPaQSP2L+1bXYDbnGF9cBdsWQ
mtWkg0GZu4u0cMt4KfCRAE2lQ/iJ9FDSgy1spA7oqA8zQkH11bXXsmuPyYT7Fcxp
fjfesefgnl+xfLz78aYwwHEGYsZXloBfPNrd+IJONL3sw4YOoZ0UyyJQzo3A17X3
zG6b18r0E5+VMfTYOv4083jYxMB3LtxwMvtGk8j+dd7U16Lc52YFRT03xd6ImwNo
xuo9ieJSnEMMO5JJUgohuA94Rwctb7GBX3S5vEMHlNt21VELWegFA1RDql1CM2kk
LV2e/dmHh6Zue9bJIRmHkb0+6y1Ru8uPOs3wrKzIOJ/rmqYpWuAmiZ0WDFkTGKH7
0gRUwGkJpxAIFvU7Zx3WhmzyuLFzEc68NeWqw/YAxYq7Ly1DZ+jZms0GfJkGAM+4
qtq/eCeVA3n18zHLah1SCA9LI41Ehi7bK/EvRp6K+PgYA8joSn5qs0OxAh3w1Der
gjwt/sSjZoz/j2ymNj1SB66WqmbOPc03cEzhTuKxltp0onIci3/fXA6MK9jtaVu0
iMCzqslq6g6eyc6uHfKA51GnlmW5CuMcotBGDLyDbur+B3fBeWMVEraWusyk667u
YVx/2PTFOQAJLxJyAa+N0c8jPQ/I7pykMiA8ZQU6DBLAOYaCJJ12p4UDyVMU7jv7
GR14kGgP8KoIDHppEjdXoZQ8MV+0jnU3cZOWTbFbO+fbY9a05zMrmbOBHyaMVdga
Dz9MABH2W6P5LT/TA7M64AuK3fh03zpv+rBzzK8PVkWM+0dwXq7w0eDb5TS0lSnV
uEqcQXm0locpebUprnEqFMhEKSuQmiRhjOBSQk8U7UyMH66U7M0f3haA2N0f0eF6
GDMg54QXI6CR7KKg7Zq07A7B6qepf17OoUsE9HYTDC3lGOsukY5C6Kp776/gYGTA
93Rfl5g4u9WSWvuMTjc5Px//v0VZD8P6jsSCddlLR5A36qKZk0ZNAsdqAh0eTqUB
KHGMVb0mzWbNU07pR0BCpOJzW+9UBdmdn8eGZjoQYLhdW2MYVjOFncS1Cddd5Srl
AvIcNd1oXtl6csUyT2z+YmTTFkWRC5erzA9kc+VMlP9k4iYPsQwbrMn1nIb6zHLA
FQbl6ZN+PKAYNNlvZkvjFDYMYO89YDwY2wVrUN7sFujKGclB7aUITDsBOmmYNAtR
6iY0gW4e4fiInsN2SerQE0pugOydfkOHGE3NHCFMxonQCSUdBIxC6e0X2a8dNMYm
ctG7nC7Z0p6iz7N///CXbcfab7P2jFUD/MokP6ZpRfnmZZFLrjYl4AQYQbNONiC7
1QEvLdNYqa0kr8/zNiPqVMZX4DmAugs13/y+lNIs09KIt+UIeHZjz1sB5sx753Ha
D0dB+rE3kcxV3UHGTJ/e/kRlx4PWSLHdSfALRZhHWb24Jq2WQmaWtlY3ssQqwWUc
OScJDH46P7ZUxa/0bcAy9P7y5wCjgeG84sEob0Y0qv4IQQxL6iow3YZP9ba4Ou94
JCNo4+5UlIqa9oebvdYK4P/cjMdaI93KqECvOiadWDnvkIW22dBY7nsE6EfEFwu4
j7v8uDhHgnli+H98jJyrV7k1rL1AbKlkKNJiSPHwK4O6aw3cMDoF/Gkt2paM48ro
7H1htMAi7s8F0+udM/1yRA72Hp6+5/xNFg6RxV48dGPkh86p0WQ0BISc23Q1PXF4
KM4V1oZK8URqbQuJpxoG/Z46fVeWqeUIgwWKUWistYStrbfjNAwl/Q9ZeRwGbAQ3
rvjbG9nAw/ZNVOgOvHxz6dGx3z5/U/6fPSJ1yZK3Pk+qtaku8a+n3zmJxgh9aLYM
H+hz4VUlgs6maHdk38wpzzsNKLamAdxz2f+HYIGnPxJTjkculcD+epoSnAsDGiOC
WhXv/ao4q0ymd4UUD8Rfgb28Vcs5cCaByUs2dlCqCWiq6hdXnxixVe53G9kGTPBm
7NuU7BP1NOzvdWXFW+H2dQboCmpeAO+JEsJ+1+6TEqU56HCSLFJDd06BLdc6l2IV
v1jYfSj7mr5ZZ0+rHwLHJuRBW28biCICneEhwGju5uUHYW5JsfhSMk/Yn9NjxzYk
R60cJ25/tO3pMbTorL/kKCWrq7JS3f3bCcS1icL0hjmH4iJSp8vF6yr2R7k+VVPg
Dl0roS1DKF0//q0DqRkYMJmxOi4raJcKbsTY9ICkWV2T6pQn+xGvK8DO9QPLOkdk
iytz+mKh6dDcnaFeJWcTPn3+PK0F2lX8yGI9N42V0Hq/arT47WtCO9ZxCU/N7L7w
jyC0p7HPzkDjXKnddNSnUhSYuVs7PZtr8BCz32UaDwy0LpqeCoXfLZoMgRAGmBjR
ko1Et8zBs9MRrPq18xyVCMPScLxHJgicEGB+nTHQug16dGJRFU/UDpU0WZz6qBoN
t8P1VeTYrfFMcH8VhMwNz/pPM/f+9V5q/CTt081cV4lbZYyqk11thS/jYCtQnzD9
ARPZppd5eTjVrvrZzgH/vilEJMbtTKfnqqdxfmZ1VV11+eGbAZvNM7DsQBKN80Zi
PKW8k1cUJLgVHRKYxDjWj2sDYGZe+CwcIuCtGyrNa2Qj0ai6+lgfQ3g/n0OjYjZS
l1Wnmw7A6T8BiZ4SXJLbwSYTAg7Lyv63SmAYMS3bYTuWkGlgYK1mKY1nnNI57vJ4
kngYivy6kz+RqHj0aE+8XVfh+Qsgm+lFhRppCI6TM+d6S1rX4/4KZg5oL7LiuDvs
77oNJrdCODHsLqqUqrCnwHp2X+tvjU7f1SZ8XLkmt294MBxykocyZ90Oj14gMo/8
l1IuMNlvqq0G3DsKQq59djA3GFupYriMK1lUr3fsKRdhPqL2i6DmG1LzOVsMf9sH
QNzGmqX70oad7TntXKL5tG5DHBfsAENKGt+SwP7j6TBkCzSysbYdcF2/jSphqhmU
FfaWTjo7aWosTbSsIah7gnrRqZ5MzhuGLapXsld5CzcJ7GoMyzAIa5ciy7UQnEEq
G11bqqUy32Jw5Q7+L/4LL/LmN6Ysk/TWf7D1vMLV89+8127N3KAFNa+nskNBcM6p
Kfrqyy9a1VbyqnypLnlgdu++d/xE8jRZ1oiCNUMmRDttE20ZrhoSTG0Xszs+VIf1
d28NezBD/2cGR301FBvD/i2DAljG1p5XZNEN3JJL9v3S83sYA7RA4U7qD1d7jnmU
R4/bgcYzAuKMlnaMltpN5LBScJY0OxglsPIIz4wPQsmM5R29q2OOvvnHkFrl07fO
PoLVWs4l588nZG8XollJihQ8ksx/GvlTv5qzV4P4lW9znmdcjPhrpHGMZGrjJLL7
HjRTOd4pULErfcbp2OVS/Du3f70uMWzIVfvZNMt7ahqIzFNpkAZnqlpYoOxzwMJL
FcGe7Z6S0dbKtx4MCGnu3r+TIr1g8vgsD6ytLwzPAEOQ/gORBF2t9pm7NpxGDU9D
N6JPAnCHoZ1Ra6FxefQkq/VHCulQRKaAYz0OXqoPvAnoxT4P5D3a74QTjsG973oT
MvGbTvZbHP9tl3P3H9e3OSmH1kqXLWXoroP5b2vpw3hnOa4voHdU8yaB97PR9s+7
TUnjiyQZOb9rrFsVvudpzNmbNC+cIB1lJyRYBUknJtOFvdtKA6UNToDgk+h8FBB+
nEoKUsJ+YIB5WTSj6QaKZ/7JBs8zrx7dmy+ZkYcr87e1Eaqdfyq2+ZOtHql+Nvpn
xlKLX6Oefgh1G/EPqrYHugS2gYMuvNWgUZoFzweRmkpOoxfuNN7aT7lOd7Aks4/m
QOVh+toBvjAoJOc4B6zHeV1t/U4KkvzoGETN7Ugkj5z/dpcFqpgu2+6RgT1Xd6QP
u/3J+iMNjFrSZT2dCua3QIicghyBZKfvuVCVTqb7wGZvy76NCxlp5UsIyeBPViTN
ux2pKmIl56hKa94OAhjwARSfaOYtP096OxetWC/naL1d8GJ3U1SeXeo860qLXIZe
SslcIwDW3rzWJJaJ42CSgTqZqehfEJ9baSXdgj6KvBCTk1AlL+EWthOJmidVvI9c
y8/hNntyafZISILIzdBuYhE/urqcfebEtgjNumgLSWyfOLLUAXhQt0UZQBFBnKT1
NnacRAAXwvfRC4AmjdFV0aD01MrMDUUfg6+6CHdcA9TGb/OYxCnlgQZeHvZYoQrC
HBIuGL10SUPlmIiN32bgfP4CJXK5dfaGF+YP9WwyiFSoQB1jrLM7DNmqqNvVfh9D
z3wYSld+gyLKuhM7aVQ1pgPU3lKjrHXzhPIaNe1T08Xnyg0wRfnDvA5aNEkKvBgn
40dXxmMHGFcMv+sUixCtSzCSdQJJGlGaIiphT9goZ9wFQWxgcCsvkuKkbuy6d5TT
u5pPMjkEetUeuizDFGTHm4KS4Sh2tqf4j9knvvKBJVLfmhibmgVgaOlLKXZn7l/3
T8RMNKnDvTDxcT3e45JfU9u33IoXD4c0xix9Vh6H3HrzIwhuNHJPvW9WgibC8u0+
P98c2oYIr9Oi6LKxNPeTq1Xf1M5bQLaTIN7WoNZweR1Vd8m3NzRknPi+BI++jIjg
BQ78E2p8kTsD/U7NPaKBqiGNctqQNLtpedA+K26jrFpaKZGBVfFBibWiK2r3nOM0
GVeLu678WXB9usGzhh7FD5l4pR8vewYeDnWSl46aeAmNCTtxiHOCneeoLjvthXzY
DeZGjbTJY5NLIoFlHIsepubt8sD6Mu+SOEsmi/1xHhxzYPmvL5QEo0lI+v14ucui
/Uemr5ZDoWNfEyzIclRA2T+iqInN0ZZRffOn8TZV8RlSGo+rAjjt3Cs/bDFpqGsR
PbcWdenWwIjqEdb1n0cBAUB1ugoxU2gYWOd1Gy0j3H3K/Kxt0lzFGyIVfzAvafSy
mTQp3D3lQwcQdgWYDpoZQ42lktXuiztXBbAle4lOM1+hdf0TuHZRSzx0rSs9zngC
U6aNE2+//e0BuPeJ0MrFwYZapiKxw39DoZwVGYzT4mUzc5YObWPi8Lg5yh3zuX1b
Av3BYYTy9eAo5AkjYPNhATO7756T4q+rovTD5XYgbVIt9PjA9LERF+jwjH+wUet0
9CVTENiENYpwcOlrbu0uDv5xNlM5XgilCG75+7azdhkgUWMQRsDOFSM5OnPOlUyE
fr8ICZLrlKYe9UWJ74/Br4VNTf+Qk28s7ZU8dViaSu3pG8KcVY3R7JgdIbiwZW1m
3jfQ8+C2TMpEeYNVlEb/6Ozcl7cOceOmnkS1jH6RzEUo8V5Ax5sKqmwyb4GFHm0Z
NuTHS69ZMzMFW66oyjbs6QgIYDa0+DIkNAP7x1zPG6ZkZfC84FtbsIQcx7x8cf8h
5D5+LC7TrZhcmHkDkxLkyMS2ruZT8XBoNUGQNttz+DAuyKfarPBiM4E2yu7dUUWu
uLXqkMDr+PcA4r76SF+NlORea2bBrNWpacloO49AWi36jj7tS/Fe3JVXU5Qd7xXN
fvSuTlaAickBQfyb3js+cqm/RN7cfi3G0C6ZprLOjU1gP7Yef02/hS8TEvKye2aP
eOOCu9aS4Da8XLA+akkyaFpEpu/TwokM4wTAq+2DNgkD/oNk0apw85gk4WhJ33VB
wCqQxk+cQoBJuLlMQChYtteu53VoCwW9dNGQMkLgE3rmZuTYLnra7gDAE1KjWr84
uiv7h7qEViAsxPoNo7ev2XLzDrWAXiUMpeT/QXu0QhJwhb5ML9Yk3hk4i0AXKx5A
u4kQoj0vYPoV+GgUmgA+bsiQDJ8uV7B9FeamrEZE+G+yW28GiSboivRwOxWTieaY
q26qYmOaoiG+sIfgaaVLnTJtbRFuwc65tE4sW9OYpaiDwZjQqh+wHfOjN0K4qSrn
gjCsEYEHEZvqyo64eFAH1TcO8iZrNaNwAADCIiHmW3QKyB7Bu3zZe5YoZyK3jnC+
tjfHvrK7sTp/paEqPv/kdpsBMKWoEMMbXdgF2imHaxUFHk18qfOYZUrvSUmXGRGR
dVYOn14kwwBJwBNToZ1JNSKQz2o2q621jdfS7WR5CbZycL/gC0wu3PNAS/AwcjYo
FL34ijDopbJbl/S34Orhb91nBpPrkLeASCpejPxrlukW29U8b5ZN3Amju3MCa+Je
7FWTcKxwb9S+q0u+9caJ1sPiXd9K/40eAhTP7i0abLdqfSBAMka9Mql++E21FtDs
lIer03bwQekB85IgHiVgUj0vjX1ys632DhV4/lbFk9+cSv4LN1PeAuC3A/3TnoK1
Zjh10ESRAbViKjcckFcuPcOZXgfgm06aRaiXJCasRLEb4w/RJj2FnjkmQfEJ/7fn
npAguTFrzngn2Oao2X2Cwl9cl5ISdFbH4vRkXKCA8vhkJF6R2kgjwpZSGKIAScBx
1i8zloj9qyWHhmssYm8Y1KD1HeSzbC8lbzoGMLIvKoG4aqcUtcwWAK4P2OrRlYWo
0QUC9iLdxDX/zohstAq3qUidwiaDr3hEdhOiFnmZXCkLVIMHlULMZPy3xEVoByUS
lM7VHTtMZb1kHlMMj2UtS+AsL/Cp/epmP1a5x6rfuhHfutC1+7cm18BysB12/IS6
`pragma protect end_protected      
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
gHKNwRQRJjDH9it3MvWORxzSQ7aTW1siBoVF14HyMN61bNZ1v5CjqRhyZ1CcS7l5
A12F9uvgVulUmLv8AE2+L+tgTZN0igr7L4IYMG/rR0r7EI5kup4auObTg9KAHMth
a25NfmYRknDlQYnNhQ48gSd/qfJecVGBIkyj+oTNQoM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 27572     )
BL2wFfMIWC5Tny4LEv8CUpzdnJR7TqMaw38FrLk+CF9Lwh5j6QD8Bfth5JxW95fI
JplEl5ppMTXJZOiuUZkXV9abiW6iA8RIL+fpnGNVnO7x/dgm3MHQmSvZFyUsZsTb
NpVKjU1ySM5HHH+B2H5xsqSJKIe1/SRki87/4F62lbjABhOiKC36xlY07hI2/YCQ
a4NcT9jCSBXs+V89ANb1gK9Q3J1p4+Wj6Mq5SXinlBwUYlc7qpWTOnneNpD67kil
`pragma protect end_protected      
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
blCoAD/YKf2q422H4QxsNAzL8MzWeBPyOjfrKTsRdt1H7ZIu2EQc3f5qH6EGkg4y
9oks6ymtS21k0go3Daai4fl2met4TalMf406zLyIwv6PTtjreE+vElQRTBAhoLO2
pVdcw9mwjrsi+m+hdEQlpxFkjNojWj4RjDNhtFkMrpw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 32331     )
mImOveyh0OsqzSk2ZS7UPbZw7Ioa1nPFFHnBgIi0fxAo7Yq/c6OtcRJoix5eUEUe
gH9ENZ5jmaAlBJ1mz4yT2CduhYnzcB8pU1+g+FtdNZAgy2pFXci/2/y+wrmRnWja
ygq83kTmOIT49YdqugVS5ZrggP2gouJvyTIDZcWs3y4ZXUTZKu6YLkwIkrW95459
SFkvQ8MPfGaxiGhOYZ7j24sukT79of2o9VKElmDUyI36k67TU/+QwQIPsn+N4wV3
IuhGlYjwW++w3OA87+2uI1QkDr+46MFAfgDP/geJqMaPfXMFSmoDDRVEVX6lXCqi
BVT86usbbQX64o2Vtwl1cwuJGyxh0AFnSybF32lhaAbWyxdWwgoHxlJILHJeMbZO
Rx7N/snB0KfB4JT5bI+uKvGyB4d/7QH1YoDrA1g5emljk7IzsZ88hA/iSaiPfjfM
ZtqjqQ2hkjq5Lmiyr8VufC7jvvIiApIMU12x4yaLMtgDpkiyGUsUZtZx8ZPnI6kR
64d39Bl6EBxbOWiXTsY1AitgxGytAcutaV4Bc5nfZD4aOvy7u1viewv1acNLHbGg
HApqGGugRXI9snGnyBit3kIfq4+yB8k5xZpmpi/nREpCtCK6mWZxMbSOliRhw2qg
YsJsyfifxpM7QOPKLEI8jF16fU6UQIvu0p4SzM163qCFxXIfZtMwKgLInS6a4wyD
rU8+PmLjTjovge5n1CKs47lIxjxrXYHTYWHYRip32WewotMHbeOKYIjoxQm/wter
rwI4tkjnJQo5Wy/K0Wi1A4La88FizE06Rz+U2SKhUqmUrV3FmAb7hW7+sWyuB++Y
cT+cmttiGSk737/KBL4fbpRZxPGKmtIxhQOjPKkSUev8EMJKWRIl+TzY4xpyi0Bt
DtMssRhZkdihr8Bl8kcm+2vv69z5ktff+X/e1GB3ZnvrNv7GAz/poU+/DjYGAmMG
ctCOI95eGyZSit5eRUjw/Jrg0rSqUe1wUmX/Uh8kcRZ4W3mzfRCl7yf32+t+Sew9
TrFJaKLo3BWxkze6hWZtyJoZwHdNFZwtqrfaUddtkMRVwjH6SAxXZA3t9xfkakAp
MCMV81e+1QxHFNtVC86aPRjQ/qv+NCKKCUjUH+g1/x55zcx59u4wOUHfWjA3YRs2
UlqgAiHMn7dZlseKIFVTeGLkFiP32Azm5hbnVnOXvD/If4CbGkQWulyKf3xx0AJp
5jJFMUobaGDK4dSqR8382MD9HU6LyOQN0V2+2lwP/tvKpmfurn9TIwGdgBly9MLq
wzgEdEzUgolc5AmI+mgMjTM3watQhERs1h/IrG6WSyMpG0hn+IO66dzNPJmLqop0
7Bc8ljEmZmgd+objgU0sQJbUR2h8qIZD7DwMU96R9Y8gS5iltPhwvcNDEZFPNZdp
WzN6VrfFmADpIKqMAdRFJAmVwqJcrJEiijJhcHyN6N3fqQn9yRqKd+6yK2KL86mE
xDv9rQ3DAipH6VGxkvoOvE1bsx8kzIE5RttcqQqXevIE4JVFgFwtP6wx2hf4GSsg
okKRNC0yVp6BR6KYU4xI3LkWwSEZ9XYCDm4n37EddAc76krGmWejtAnxBXsloc3V
HB0zi65O4jtjYaq84GN12ADnPZTwHZhWiPKy7wsK4ChBGJ+Ol1btqe08RYp13thH
kuW+jQ5dorZxnHvAKUrXWBXuBm+TpSraN+8mRhlVxQ0KXrLjstl8aFjZdTYzts8F
tmZM61kaTJZXfmRUcbcQLtPGWEvJ9lis2l90ZkVGvD3V5cXHGpW58gqigAEokUzX
IPIT+QE49OIF2ZGZUQ8FLkaTrsW0tvbkFmoNv9HjBrGldpbKtx8CH2loMQGl4zeG
MGbCFE730S26vlkc1RopDjObcFj3+hzORvrr9euXUkK3nAMhJb6rcFvSU1Y8bwfW
vTFdRJw3oU+hIWrTFSdYaCqkQXEGlKu9qQzKZFyNEWJ3yumsYSLFVV+NLcIIivbQ
rJZkBt97Dc3VIDd3MydmOCNpnaMX28TP7q4MIQkDm3vonBZUtrKNA2ESst9kwYQH
JbLKmJPVyey+5Z5wCDiVMd4QXRyuF2Mzvt95g815DBxLMGu2ks64+9AHEmPo4IaZ
kB9x5k/uz0q698IV61hfKNFv6HSRCNnz/QL8GtAOPZ6gf2q+dwl6S5kfqaBXPMRn
/MllS6d8OlIJkBo/biVFo79FXq7JO4BZnToLQQm8p69yW6jZZ5ZRieK9Wiid7ir3
Bmh5s+wecmUXDxwfxlbv8ifZr617B6+L77Z4MlFRkdZ2Iz8LZx3d6dxZuRplkVe+
ppMfJWNCfzT5FIzTJg0xFgJZc7DupbVs4TkQkf5+xZATeArO8uZzv90iitRXT0X3
VjykSVYsIeOMfptABJ+9agXY3NEDvSUh1DrNwx40OmIY4MnlKqQOGUP3weVLei8N
35uJn3bx0zdvP5dS7uWmki86GyxSTcYdAj3Vkp6htDCkNTf+a75eihiv8AzoYZt6
bD571OXOjTXW+hWrth/4Yix/cvTPiz6SMalt4W/Yz3gtloOgYnClN+h0U/WcSyNr
rm9h0WNAMx5ZZcFOjS+pTyDzgg0VrKkn0mhMCja3FktGNXGJ0tdiM+rqgxW6BFGF
WpPmMrI3adO8kGhgn/AJI4fXSXXG+YNhrocXtxE0b48kQWk8SpBwvP7/hXy0yYR3
hmbiEB/tSPR64ls0bEdrW8tBArv/6o8GjK/+6KlIr2nG1F2aCDl7k+CijRwUjqaM
rz9ZvpNJcK8+BNVpVRKa3JQUBdnT9Xz1Ez+PAU0tXG/hUeYJyDknsTS5Ey+BkUl5
6deRTa6lSZYSkpPrjQ9s516cCMHL8C8t3QX5LP/gPQdlqV07yVMLe5GsWl/p3u5D
S52B6i7NHtT9bBWaQYua1FHOA1eKuA8kvJZ653bpyohMBw8Q9KjrwemRzKWQ5dGx
XDnAHI1WglQx/ckwFn6OtHyiUWuR6QaxbpHqUwGZuNYpmA3n34hmiVWheOvAdcNs
mR83/FEM8wTAsl3KYEyEJ5E+7oL8iM94n1zziIdTfHp+iGVW23LdthNicwBKBqho
CPv9ceYqPgQeUCWb1mzvQicgzhLv++bV+gU548RwKOwE+fkVaXMZFEBa4mj67po+
3lAOAszh0GXYckFhMf40QIYLgiwhRZYq79kbY7aDAMUqmUPglnIWNAfTnvhXYSLI
VdAb0Cjp60ZTVviV2jn3TME3kGJ4eqxUMiSB1Pcrl5SWPAhH31uuGAxQ4bUw4fRh
Y5vJwfux3wiXRedzlar4XQdIumWySg6+xtyshs1CkjJ3uVC7JsoOJf3DnRRpDIIL
77/Ka9BtJAbS5jq875jUaaFEPmeMMGN4crZMF9W+8YKLSBd1Jt5yDuf2Yw3tnDQg
XjDcHDx+VJ0b/qhsIBOokGW3TYHnDxyHtTVFjjzUaXRJuvOsiPMxmV+WluZK+Z8Z
OjEXm09Mn5iVX6cHtuQmCP0y6ZwlfYSfdKtC/yUYZTp0Y2QLpMpENHqhMwDDwEv8
gf+SzPrflStAAoIrFe+63al7m8pN5EKofZ5n30AzNDo5d1mtpXSa20CtJjsIKOgn
RedZsub2KgdWYyo2UuXgxICKSQHBL4SoZgXN5sX1EVCgDPwOtzRMqtHd848BLYXI
UNGlPvso6PMM3Gs00ctwmDycD7kYzr+K5D1VzmInz4mJr7EcEWIZU9EWPA2torZQ
B7mY5caUOVa+rayqzxULI8g2RVQf6mMIe0/BrniHxQ/qYQKb1k9gVpWTB6eFh0zl
8iHcRe10qSYM9F9ZiLKV36ad4FT//Xmj1NDpaAvEle3oNXiOELO8w5mR14Zkm6pq
eR9iMS8/L+/9vplb+pUvKWDRlB0Fkrkv9CF9BlxOlbbn6Eb9UARjK/lqH/kQw457
5NYth7/kwu6WQRws1z9TFbuVhhzrAHOIhDUz9bhYtnpzL0uugLCFRIJI0+Z4buI5
J38rpTeJuv6K1e/cxgcstwIWbvGJQm1eKnQkK2bOVOb4eWcm3j+PpTbbJ1DlHiJ7
lW6i3u+o88fOgvW3DBDoo+e1WoxlkFqkkFja2x3/R3n1Z5LACpT31SvyC/Tc6goQ
qBunX9XRPP35d1IgaW40M+RZ3wU+9s4yAZvT+eU4HA3w14U4tTFrXIBY2vzTV3mq
YAzxtL8rrToaf6YCluz9wCvrxd8qtCg1t7wQcDZzy5bYtz5DP36DB9lGmuu9AMUY
LRQX2PgbQ7znEQyNGAVn0OeRqLMwSd7JzyRdvQv6hSsL3WYldJxtYJ0c+tL1Nc3O
z4WZcGMdJxsTuAPEcANxtV5I3Mbvm5DSq3HMHlqNbtNGnzGmTaI32YBGtRu++oWX
eGfgkQdMDPU4r6AFnJrO3Adpxh3wnq1YYlS2LTE1Wsn3sViPX3wg6h5epLDio5rQ
tOevrAHE0QszzBnd7GwXpF+hkz7eHM8knCDcsqhAB2rVLFGJJHOXyIf5twggKqxa
lKgdLWKiJD08dtlGRM6dg+jsiEVruy7WcZ/1DWZUzoySd+e5zv/xeIxVaDaVT5WO
iybmRf2E6DgmrUP/TkISueKgZUKgOeAiBwlK3QJo/CvmolsIQJoeW6SX4p6bJQUV
yBk6slax0KPHJRuLpZH+fC09BkBqsLT1khBBccAh9TEURZHEySKcEUkzzHJzsLR+
94qIK877mqX6+DuS6McuhjkhfLD33YSx1HhIeVAHOESlKzgRthsbEiW3moJt9sY9
MR4cmFPTci7IbQ9Tun/0h15FLnMk+sDGYrqSw/Kwm8f4HRgOiDmLQmc+8fntAkYY
BKwwVN/IkMK96S1xc6aSA0oMIkrEZfvE/iJR3rOf3vHEw7Z8Nol2VI3MeLW9lZms
bJRWmr8uJw/Ev9nQwvt9mgWbPYssl9SwOZO2rRoxEoSZeCVNOAci1re4ihpnC6T2
GG5y1I/CtuWh3qYsE15muNQSNSaZKwMIOMonCUuDfdScfi65ojUGbjvsAmMHjzpW
Iqn5QwL/Y3f+xd1H5qnY0/OogQ/Z8Ozrc6HQks55K7/MAYTT+nW+jn66+qart1Xv
4QJ8wPP5DZxT0I5vXs0TmXRhi+xFUZlKdKYQ21rQFLyI2xzttU4dtaZcF3ZilG63
zsaCR4HH4AckJBMlJ/ozTLlkvD9rYr9gGpxMdswK4BEJv6nNY9UwzefHWqK008Ib
UnLVztgAMysS5CCEOg0G51AnM8oJXvOWbpkSaI5c0J9/e64nnShWGtjwIKJEy5RT
K6TTv8/l6+yZrgcFEaVMz46LbTIFbggEO9caqHV9zk73k+PZt+i8S/KMYiA4Bvlm
MOAq4s3DR3iXi41/iMTT3aKkYJ81jPrQWz5Co7/1dKUbEsSeueDTp9AuTLUjTyEz
wiTSQRX5n27rAkVIl7Txde4HfjD3HA7UEYte6p5olWZpnJZ2kozMbQjHBYp1rqYy
KAVDSw2UUYTKanUJzU1CCn5lRDPLwADYvI+NsVBgYIZ3L3/dFalcTheWr0IptcOX
8k3TTM8ZJ3GNy8NQh9gkod7spO7nHFsQHBKOxkDToOHHsjM54hnEksIR3ToFnQG+
aJiRHTWrOnRTbafeR5jeo1Cx6KkbEYC7mNNGg4mxw3x/CKgR6M7vIw9PBU42noRz
ny8GilRJO2BBz8yCkj3zMigkkI5yK1J0ZgkQ8A+6jpbx6vYb0XPl0opwQebaMi+x
4LucX5JsnM55hz/Jh8yNz2e5J8JhNCPFvR4VtynkvQElOxE/Bi2d/pzOzAPAbNfz
/1cQ2mSOGPUFPhDTUDeXGLkmGOz0l/yqCtxILieO42aOECp7XD6rCDhl2PB96oxG
gBI9dacKf/9kXH3X1IMMvGlKO8RxGtR0osM350aHEH6F+QJ5Q8b3JRQLzZboOMQt
FH57YDc5gb4FmhBhhKCb3JHvS/43U5XAw5jlNMchFeC5KsO8IfplONewVW5HDtoI
rZ8kHtMCxC/TGM771A3lrhxRzKYHE6dMWPjMBdXw2h8D+1ziXLEpCVK/MxNRh3LO
U2gT+I2IIBzigy2t67N9ZOPafwyFG83VajxS+U1P7LVLPNGeLYh8V4quJgLNwf5Z
qEm5s0Hu0IBEjwAD2myPZUMtp8/Fbb6ohlKeftA3u3hCUa8L7aL0GYZ59udlhPnY
bz+AAJRMYFZDgdtKAbLb4fnztGW9fk0NiFgkMGTy5p4uD83FY0gOHIHbN5cPG1Mx
QDhcRG8VyA88DFBZOS8B+5koncd8q4upfj5Kb0P99cRT+BWXqRFbscW8/12IsGGu
om8+NtjooBBgeGqm664cgHwM9lQgEHdDSl8HDKTp/FGfIq2z4lFQb0hqdbEl1DdY
6oKtmtlsqnxq02qkLO6CXA==
`pragma protect end_protected

`pragma protect begin_protected              
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
lb/5oGGdSwF7ca27jTJC9hHn8td3ENzKmUk25MXVRY+TqlIkzVQH5JgpK+FOrIAF
SquQvpt/BhNFwZ2bXnbjRYYa6gLMeMYyhvLB7w1Fmhrd1PdTcJyr2//aALqeXQnK
pbLRL25D2aOZHu4OmfMuBanxHcS4AqOmrHsxmvutR5c=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 32514     )
1xCQwTkMeDfV289G09Xn+YblNEoNePJhv2B5z01Uei44T7TVFKFWrfH/W5omlpEj
oLpbirFDjIB3D4IGYC82a/uIC1Mr2J9ZEmJxLYf4C7kyzAtHSbCpiMSJyRrd4587
XVDKb6sBFQ+HwDutzcmGs0WKoKuTrzELBQP0eyGqhRJLz2ElBAHygI7S7JakNb7b
V2xTcFLfqpHKCCHxOtofkwiRf5sW1kIjQ6VU4BEpOB2WRUY2mJB4Zl1f9AnJ57zO
`pragma protect end_protected          
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Y17sWLpfjBwlPo2GIXjsLOsMlAoci/F9SCIVvCkCqpS9tZfO/27Svi3Do7jK+4jI
MznrHONCVKCykvpYjJm/78a7tvp4qZMVH9qsYuqmk/ldFGr7wjvXI9tMd6SNzMjt
Gpf9VSJSpKXHnkZZPyZ+3i9KXbDqELO5oTE2ZcUawHc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 40372     )
xTI+KKVOu5Lap5T4rAMGAcmebluI6PgX9zT8PhUhfm9K5ZtwQZk56qcFq9KB8/Uq
5Q0ZSnFWxW9e7ANlYc3L6Wby3VnB2zRsscUNdBeJZkO3fbytJMrVkyaKx+c9jLx8
sOgU/7pVu/SBvZgtQ/yFPwyhfyexICqSuZGRboUQq8e3LBiVIFRY0YPkR0I3nqn7
aY4Oj2BexrO4eK7FKU9F9/L2q3jtyV8TMvLlqQow4I3B27hHvh4gqFv2C/ZIFDtg
0dIJpiGFD7Xg5s8qwg1CsHhfCIAKDeTDw1fhGFwqDd0Kujr4AjYFlJ83p+/EMtMU
tD7pDmxCROSGKoUcSeCAcFXD0pBTx7AZ/VrSECt/mhn+rTCBLn5se43BKlhncdMU
Yz31PEzHVw1IKTW40GSwlLrp3+hJ7ZFmIIUhUKswSImvZdTmKFI/i51vUx8eIi4T
9v5XLW0tEf+t6MvDbDTfmU/SdM2g7ograo7Sblx3ODCl3d/aOB9sPygSBYJz4hHi
Hp9habZnv8cpa+F5sjdbwmgyRGbHx0nmlHYsZIfyS4sjL94AVKQeCka49DGwGR30
8MIEVkie2dxCazU0EBvIw2S1R7Dbpg93+5YuEZWLXAeJq3kelHCcwM2Mu6Gur6Fl
imFH//Tvv8FzL7rKbj21DBBqJ96ETw2WphcZbXlJHY9X4Y8kfV8ch26FGubNRj7b
mYOgxrF5THBxEnQbcIPtbdrDlRzduW2TKH7vY3LLh5Fy4WDcQZOhqrsm/4qm+unx
M1Eao32OttMvgdMpYkcszwdu1qDgCQj/Xkofwuj+BFzIcaR7K2I4e1qLPDVT/9pJ
Etbf7p+yuHdL0G0UsMrAC6LCc6Au3gUNhe+NkU0DZloBQT75nns8cYkm3ZTB9RMP
LRQ1EESWT9m9/+0bqEQ2oq1llvSuMq10OysRQGZnCSJ0q5Rwe4O9XBrs3OYQyfmY
hgS0ULseeVQXnFF0Y37J8OoYoB7y987FsZgyXj05OVl7iWeCJUvQorFCszdC31J5
lv30BYakIAx12Aw96LFJQfBhl17tEjh8ouop/cD2oqML76FO7N3zLNbXF7d4JuFB
XsfwvA9S15e5Qe6boRYBy4qZzXQQrpM5OApY6CLeqdpHOW2/wFDnnWAL97FxNibj
h2MuVd3HLO//f+xt1N2QoWppnty3RV7AVeKHFcjEFoij02bMeles9XLEBWKqfhi+
SwqEwc5gZXqy58l3TRkuEl0dVGHuG52ngjeZ3ZDGGgZaUrxexHARR1gpz7FvHjvr
ZxoIRJ9ZS0z0Hu0dGiF/9WCRaD2/o4Kj5pCE/LkdfSWyOxPqlsOsyV1bCkKvM3ld
UloBucellQbEbotg0lL6nCpdW6apG9xkehRDFc+ehljlQSx+gEiTkFNiq/vM/OA+
kshXRTwGYnX81KcP+wdsXZyPbz0ghKXWvjdmAFl0JCPgSf3eoATF3np4f4XNUJ1l
NhzGtlM92RUdl4yo77nnExEW1XoEg8gfw1ndCwf8GXWm+Hjd/h2dEDa/EA16TQNv
wcWXRFM2NErl6/JlquH9aSqN011ecXt2rh+Qvm/m5Zy4hNCap42fRZnMloXazZcm
uZUNr5ayO1AtUY9zK7M/rTyyZRMlatGF351rHcLmBHjID+fo2W+OCWy01KVHOEbQ
so0c9L/ki4g8qfvyh/5VMZKkurjngy29D2lh71pDbMz9nOAZCHFXJrenkckxzZui
LA977Jh7W0WOFmG3FRvuWjqHHjSU/yB1XD2luYJQiPYJxgnQ38sI36lMcisBXTj9
YoKGMqfz1G9hhSUKqbpgc1dDpQrHScz6o7k37LSHAwNO6yUgEcv0O03w373/myou
NnpqTwTc93+Qei1wTzgK+TgmNZaXevWb2SHq4W1IvKFnKR08Cs4scPU2XNnPjAN8
xjci5vl76BkexpKwL7WmIixOa834j2K2oSc6XvRIoWIgJISI4ZBuxU4Sdvw4KRfq
WYx0bk8iJe/hmc4JcQ69ytjKmDtcaeSD+EDZKj+LSVuwmPTTBJKEch2CoR7sxSr8
gsm6m0S9aLb+c+AWjb5dZpWlhoDvU7t50jDZl4XI8hfrl5fBxIcSvBIXaPvu0xXn
m4BAFlhJlxJ2MghAl27zB4Y2iQGfw76PQphc3+5thiCVd2RPVT2WTrQ+67Uztxme
juC2Sa/5IxHcrgo7Kr10HGPn2PeHMWxuuWDE+6+K/OHds8okWF7QGwc5ZUuWHERV
1kkdFhrGChERYKVBY7w5/DxUgn6O1RWjuFPIJq00KZ+enPR9/swV/UkMc0BMipCT
+fuiriSUjsRRYVmeICHYDFu9DKdG46U4kZjJi7kvKhOVChZoSO9TvT0iToi0Zx2b
AbiTYVPqOhtcKtUFSBkPtsUwBRb5EBENpC6oH3m7SD9JrkiQQtfhohRk98RZFp/r
1neI6Q44XRla8gcBRfsc0NVuiSv5Tkdz19sVkGPSsLRux/W7zYo5q58cGTEyg02Y
Okhbo3FXuNI9sqB8o16rvv1BLd8Bpi99tf8toUm4eA9iOnMEczGCErWGJOu6Isun
m6v3GLH2pHjC6Z55I0HL9KZYSp/DHlK0UBE6BtZawDTv9TzC2TRtRGt768FoYrY6
TMos2OZROx6du6h+ZKNydr48Y0s1NS3ztrhtRx8O+0+5SKMBxHy6vAvEZAlDcepO
RuC4T292qm3kganXLlVaATkP/oyNjHstB5tuM2RyxekZbUi9XK9uADD670qZdJ8c
Z8q9OB+R8SveaXXlbCXjIG9+esjdqo4kfeIhXpTcYGBJEg2CZXD6b42SXqYh807i
KUMtjpVoAN5x4LxQOixWxziiZhNT9E9N26EKFvKXj0D24rojX7uXjtIsdiHuotMx
0989l/QY6qCYVu38VVf8crrVuLhJrEXhwuHYBfmaRx0wP5UDWTSLu6YcO26WNdvI
yJRCL3avl6fePJJWLhCSPJESG65eMSfvDMeXjkBAZ0mtOuaKet9571pAvTFKyNF7
iQvgRsac2x8G3+S15x8joDAwRS1ZZFLliFj1TcIPg4PUcWubeoU5+slnJUwAkdOl
hcs94Yriah+tm2PIYtB2sh/30o3uPNemVaBHNlL9YHeej5mqG0p7wbRbJo08v8hO
zIOfgjNmyN1ddu4LF71tUwCYEBDmFGH907ur/7fRW9f413zYbSBAXr6xBac8q5fJ
hlkzUQZVup7DznUg5gTeX44m34xBZHpw/VTwXZU7VPN3IoIPPzpMyB2pLdlCWGjU
pAU6LXjwbKnm1uurAMF3K19e/S3CCeVgWzBhH85Hja5vnA0zOuc4rjBEnK3OXXVK
A7vDQIGJckfhInWSu3EZ9YHwAE6NTaDxfqhva+f3TmNXIIqbiy8m1qEtzhkpCnN2
xabaKdrsNPQvlTnuQjWOqowuu5ODVg0nGKWJx5mkSBVgRZD/q08i/HI61K4ZlJ6t
oZcFM7hJ+ng8pocIiiLb8ScclX58Zt1bjyukOI9F+VPV1hTjkKCpmcFLZ1BqBW3t
q0dI1ZIQ6W23tUGyawMkGpwYEeoKWGAYgGyPXsOzv9BztcE6VKWY24YxMquvSI2w
atmbi6Wl9L0TeG76M9VkWcoTRvzxVm1hBTxVu0x4C8Vjq2U0sZ4b6+IWBl1cP0yo
6mdyavEF0vQDCljmZBLphCWmgn9L9EfPxrX+snzX/yTgIN3+v7sgXHQOm22C7qqB
ke9y+/d8AgqNMWDHmiLQgfc+MNeg64aHH6QOzeWU9mD7EoIk5p+IyPr5LLXr0CAU
K5aDt2DEA6yFwbZqaHGlAyDU0+58ICJIu6ohULvg6OAh1liz12bBu71c6/QB0JTm
iDy2Zzt0G36KvSUe1XtXAmJVrWxyiQxIMVdsR+l1BOHcCwOIuTYXs7gjcaMdO2FI
F5V1+eX2uNibge2OuOBk/v8OCow0t4BwPZmWM6naR479eIXe9WlgN2RwMgh22FFf
d5DzjzMDN8fT30BlHmslRUVf6xcNFXORthGWZjiJP4pEehQeCfT7lEh9biiQ0Qup
5M3Xn/fm6gaBk8YI88X4pbk3znJi0ggceGUYg+XebR/Nv1JudlYdtlffKYulhzYO
u/WeZupHebuENYbeAxKlALqGzg8BPTbpWRvvyI6/7mMEVV8/Nyl7X59ZFrc8HwtF
782pz7IUljDVcKuPjdB9FxiFA2apRaqbeJYPSfr9Xsi/0wVke1EOPxIct4s1IjZZ
lUAT+GLH0IksPs5RY+OzaKWsZglfSaCQKtiMSQJz2UtFWlYZfSocfE+s6L8Qx3wz
Hb9FE8ZZmhAmm9Uw+tv31dZK2UVE7sbnqpP6P6VRA/zVG/VV2oIwRvXtibRAV2H7
4iqzAWoqgf3A78rFwdozXw9Sr1Vhr+Zwm2R/5gxBYoWkyjS3aiCFFdq8R5Bw+/8/
UGi4ihUUYkYFPE6QFHSgyOk89DVpH+cMGHmFNiuiBXSvovticYEYB9uiAPzngPR1
GMUhpqtx6+gS1UiOjQRcLi/TfN+24QzdhSPFMkCEDAp/+ckFAutJTUmHqpSNRYQ5
enEusfh1QF28DE6cYJ7QzjIJOr9kYlMIEHBE8WIhcr7phIjCnH0tegezU2fKgbR5
Ku+CdX5XbCa1CtGuzGWBpcg+mOwn2xdttXJLwe3jMpoAay+97ZBRVviE9iXE00UB
KUpivqppT8yeUmO5c4UVgW/ckKDxcQ8KQkb2V0ItctNspINNumhwPjEqv6MvZQn9
lyKmWXx8sWu8JeeVndyK2iW2dP41pYnti8v3OVvYZ0xHFtzQw2RCls5ByAmXju84
DeGfnJlBODVP/VxbfNpa40snsecDwHfSrTIz7sYM7sq22oixGI0KXAe9TjJIfPCg
r9YKSlfXbFkF8IGdZVbWiBNpJ/zU8IfDZRFf3J6cK/rYxODtkQEqVEy21fcztqHK
cepk2EpzmX67sylsLMxcVXF219NzaGJDymTUbc4rdKoEj/u5S7g2IV2qEbUSWi5V
weGsf351n9CKZ+iHWQQ9rhz//8ocyj1y3PSJkp482NfUHHGsJkrEcn2j687CJOA9
tsiII28/ZwP2luB9ifzdgw32/tyuxJ8ROEA2H26z3Rr16ZhK0tV0WeRKdNLUkDKE
Xop9tp2LBalS9Uj67NuwsQhS9IkuDT+M6JzI5f2KgFgQxs5OYiDAXNMRwsmm5rHd
hQqBejLK2ihrqkec7X6ASpJBPTp5aYc1KLxfClM1VY/o67ftHa8HW5pjrxWQDinU
Aa75TYZkM7GkylmBFFzXEQRs3KV8qE0faDJeij7MTvhEwUw/SVYZLZWbqsk9qYej
43mDp9NKVgoUpAk2+vBhrNP3KjFhvxMR4XpdIpV0W3yylsUh2fs0EoI+OjCzOtFQ
z98p5rQpyRTmpef8pyMlph4CmdKNy+T3cZgxV7mIi8/hYdjny808DosYls7DDOG1
OfAO7t0LlUOIJGTVdtSszp5vy2S3mP0Yq12SmXY4EjKOK/QROtCRgUVlxT7BoAwt
GIlnpxyitKUcaNztPg59QbF+b9GQv9+JovCQffw/1bYWMqao9zYaglQHClhsT3yI
yFfmZZjehu+paVmxMo9WenqEukRI5xhdulYf/MuR/As+a2iezGblGy6+Hcla0EFV
aKBV8cNBd1o1A6rOsDa75Gtr4TTQnexDXXz1+ryLsQ96Bogyt2JlBLQLtCdGTJrA
O9axJP/2lMDuP/Cx1bNNRZkd5NQAe4dy3nX5hH/fFNIBfBlLi4ffr5nNvcxAVyl8
jmbynP8tqfJNlxbiOOQoDMvQhSZ7iXWMroFj+MFtkQaymf6EXOocJ0mAgkLolknN
mIev+b1ZS7TKPwDbwxVgJENzRVJAzEweJEDFM2mQBxZkDCGTlqxz7SuKT7AAQtFP
S58IhSz20hdW5aAfNfz4L0Euy4m1pWJBFoXGtmHyw2lVjnfD1/aKh4Xnsq1kLq0u
aCO3tPSG52P3fdszya9ZMhMxKF9g7IIzi6pwJCtKQYFgUmPXyEvEmQEAQH+LV520
9KvlQrRaul8/kM3Mq0ZIe5a8WtvapUIVfY1TZe+E/MkgSpLCXpx7qg9kxaKgaQfa
suYViljAeaclXO/vr3A2jgnRTva9kNzvDG7l5WnroGnxVbeKE1dI9TwMuxZ1wHBE
Sn89o8jg/aY0mw6QYre52jvZ/K9LwKAranHaBV+Z4qrW8WeXlg4msXavd00nfj9i
93we+KVhuLB9JicJQJ/Cg5kVATr4RXS6ACUYGBAyLRTADRoCtAkcVU0oFHVewbsi
Y8h5skWmqqGKg5QnQiAbt2IkFeR5F6iDkCkB8TzBYNoShqeXLlSeETnrLc3nghdf
bkIteGmCHGrYV3hkFhaYqVHzVwxTfbkl4lWAFGqCY1iA3c1cTczVNElFEdljh3Ad
+Hx6edD1XTkk3dYjdyu5DtdZ0fpuV1P8W0PWQce/7+rvz7MiDp5R3kQRyoSnljzL
BxmEIJTozYKWIMvUXeN3ek/To+XW9S6YKGtG1ZXbjByRE3K08u6r7DQAs46DLolq
EzDEKv3tTLIT+pKvQTTRYHD2c5QM7OIHOiS+mro5o3QC/y8H8my9/sCYCoshgvFF
eKmK60m1nnXz87i0U0D7cboLttmK4atxd3/ak6JoIamNHXRiq/f0u7LbT/D/m0tx
olmRfbbgbJUA7nSsr9WlITdkQo3PWvD5qEz83Io7yTepExhz3er6EHQZSYD6WS5E
Px0+QwfnqAvME5quEEj7d/4SnxMM8+FWCjVTLjcakYEwIb4Xt7K2XKUbC4Sbk+IG
ZGFfMOho7M4aXaa8T6g5hURpo66DhQQlvQlaFEoiE8na4JIbpB5vhYtuc/INpDxP
QbyRsrOz3bo5ECVoPSG9ioNsyUkZ6E55jGF0TgAFxB+bHV1iETnsG03xgREvQef4
VFF4FIgc/s1XM8jEovxt90UNOEieJ3YS60G1h+W2u7pehbTzIWargooGzavKvacC
4ydhqdZflvZ18pAGdNJ2kbZAYCm5am2SO7obW/fNGTOMpahLXiV18pOLQ0WPt2q9
/hX2tS+zTe3HJBB57BJUw8elimsOEY5mXI7KSVjHdfUcevMvSq77UTxlmK5m4f+K
13YTJ+f3wUUNAJdXmbhSu/wRxtIVI5pfhcvux+nOmV1HwBqBGtVaBA766AzvywUi
gVgFUGL8af0mibjEp3NFqM1AD5yl5S7clTEafJA9i/ticlyeU48GKcqSEgh2i6lv
u+H7Rav+/8u/fA2pz5HfCe+OdxRROVVPEiSrLX5vmUWUWduk2oRp4TgsEhMC9/xR
Z6LQBl90FUiKXr+1Ix6WIOzmyuFe3NPcO481e2Ka6ZtWww95zOCZHxoyRWzCj5AM
Ec0yOfXqMzgKn77VhhGVopPyx0ArGeGwgVf0mW59FUBu7MuemQlavo+yi/L8tCw+
10Fy8OXK5xalj5brWFOVGo1Gl6P4xGHSYIfuw0MecAvz3wc1/UbWDZkLxBp8UaA5
NLVSir22m4tZe0lXOi2ZydPm3sJZFXzJJ2ba/lfGrqHrXfNkTtUnCFKsjjrICsUv
jnrS1r6DqKHO1m4LKYdnP4O855gbItki9SHQ19e4xFhj25omu6d5cUlW8951FWVN
uELJMVDOUauAPyqz3g+lliVoJp0IlZQJj/fU00t2UIkQ2Tt6qF5hMfRH8VOImt3e
nkFRJlpaxorC+6d9b92XJ6ixn6VWuFnQ7mdx8y5u+A0VaLtYxQO29Tk3Up+7NBDm
rb9M7EpZ9tX54wgNCdtcIipygVSn9kg+zZmwZ/4T7rrvnS7ZozPK0vzTho/Zucu0
1ik/f4DVm5tEFBZKzntCUDtsavBb/nf4YnkoO9PJZY34xGcT/HgmNzvBQgP4GUsr
UXdO8A+GeqXdqJcjYKifax5HXeAI6QSjn2c/UCmkLECAxbBSYyXDbdlq/whCu9uL
iHdse4ilOXepaHPR+Ux3EVz/CDFKo9AZWvnaLxjlC3y/vASniD6euyjUE6PEYTdh
g1hHgsxid1W2BkUMw6382F0zxyTe/emTV9JdZtLVm7Y3Rtyp9L7Tm4iG9ajcxP1L
vfACmqJeBWQW2C5Fa5YX8NP/xLkU7ZY9hQcyd/FPSlinKjTuDaM5moBMQjhTgo+r
WBt0ZywrHF2UmLVrDoBa32cDFWdCP5KTwaQs3BLgRww/DCb0jzHMWdxFiazFbm+K
DACULxtCw6eb3z2plM6WNWCB1mEwrDNwzgzc/ftyI7uSbyZ25NHtmHc9OTNVljJQ
sVOVdr23D1N222hJCtaWRnkXCGT5RQCUcmY/B3TQj/lKWsKz/AQbHA5a6qLS0w3a
qvyavmkxQHWNjU3Fe7ddD3EXXV6vSReYUTmELvcW8LlbFu40Iu6THxZvZRyZb/3e
IkuiPsfbwI3Rjf+XiJHCCsATDGXSHIdSG8HAuBG5inDz2Vd31EVF56C6ShkF4+wM
7OYzI3QwiJ0gdlmwEPBRmnJUWWoMnp1QZFDB/Xq0QD5NyCqhsnIQJyBB44+U2nLJ
sIx5toTnlZcOaZI11v3lcP6zSgunev0z7sebr0EoEyD+tV69AH+ySNX+/wmcCFm+
HrgXDalLLMHt5jkS7GaNTqggtAw4ycrKX3s55JYtN7Ss65UxA+BP25YJQK/OBr3Q
gz+lQsSm41TYSqzzMmi4mNKVrFZAI9Di40NL0/bUFFkjV4hmM2kTEbMvLNx6wPCy
zFm1Yb0UuyaYzFo6K97WdEcBSCNi8R1gwa1Icm4RDYzKY8K5w0yENSXR3eW3oWGh
3VAi3yUpD1iEq3+lif6MYXfyWpUH7VMLag2mvcdn7lDUm6yzFaK43f2AEdp+CyHF
jL33XNa/tJfYdxNCrJ5DDFgzFvXG6uYW+eZr4DXsilFrcSQiRrJ5ot8Gx6o07k1B
9GFbEPlUEC58pLITCifLvZs2v0+6F5KoM5osXWykiDgvtUsFO369eyN0k6jwOqfL
JdiYBuavd/ef4p9tW8NL6mBzFtXv1G4Um2ECj8siiekSJLFEdnbkQ3iVpcasq2fK
+i7x+MeSxnxfKg/WcN7MkX5y6at2KOVyQvvz73cJzA9Brjl9axserauRHNa4Hg3o
RY+AEVerMtj1MwKp+WgPP87X2TwpxIKgEGbjLNNeVg8YFOJ5XMcOtgWJVQNLkOT6
R9z9zZN9Kyk6ohztd+7svSgecmF2JHe72JlPTrwhY9GUw3gamNeUe5Fn1LeVPPV/
OZRD7PvkCOyQI6OAPPOwsSK3PWbFwKWfywUdvmBSUrwlM2zb/obyEAo6y1Evhv0Q
oQ3cgq+A2unu7k1+kcuBefduyzYZuqKHWiYYdxcWuarFsmQvaws1NNhOcWp+b+5a
eAr7BPPmf4utor+fvG1giP6AqS89EuoltP+C9OHBpqcV3VZYKzAL1tQcqiOOETp0
/yGdAaWXFp3nAgY4oAXLmUM9dDbAQHPbHFWzCRvm87gxHF2YLIFeVUkXBfBkuHTF
Wp8Om2Pyhf82kHpkIuIa/DZRMcTE54Z/0P86rdDEoDOY46oxt6v71HWM4xiSnU7f
u9/I3gI9bYE7HmBcjl4BWaxti9aT5Is4HqksorZlYQFt+q4MwIBjjxjZQDFq6ioh
EmStpC271I0xtuSnQTdbJa9NUXEgISuxJzcQr4V/Qwa0PlOCP5OFw57I5PtbO82z
kqMj6ut/DQ+GXK+Fg84HAKw1+Py4TiAe0PSH9cvmuhcjFSbtZh2lL1sJ9BLIGvfZ
a/MOEXxe0VwbHS3uKaDV5BQgXLhFCLOXKT6BsN6i6/Ty/xg+V5YyIv/X8WfNUfYA
PODwHUFETFMIBufEiBkMLtKWL+VXsqZA0Y2a5M19rGAqV82ULWL6cnEnft8izIBi
0r1Qn/zB2gwsg6m1ao0PDAjDegxEZ6A5Arzs2VDSDA28pSf+7o3Rxw0l7Cev4N5Y
liji91WOoAFo6F99OS2JfuPoW0abrqkJd8kFNMBt3E4YdRmMLn4oHO2TdvGI9EhR
9Q/1YE9HB3tuB7TJPAYGdCs4I5p3qH4NTUpAEKzSKYC16kQN8k31ZKtoDsJko4XM
uRBiAaZ4SFh9xxYxw3gJADi85TxqFGHL2HC2xL8wEVO0ejSuxdHzO9oHOVWIZ0h0
nEcOIYBOiPKaqE2Y34NWzbIT6gACt1DNENjwvMzLwKvay4lLkaHPX7p/XtPz49xc
G6hsT5JlUGg7PgoKVHR+osEpvjyBuXqBRDPptP3Pe3AdzCLjHGV7/PGBuwHrXkW/
yj3YFL72bp7uaT0qe6ROCrM/Mk2tZ6cVCslvaYRlRuexJl5pRFQh3wsOTG68x8Yq
JdODEtmGz66IODQCBy6Le7Lb4FWvN6ZvGajYDpdiiZtVe0m8jr8D3+cUFFQuscNk
bRkJi+OWcAq/eNbr3FppgNRKoPa1qwzpGDDOSLzKCQiXpVp3OHoFQe718s4/kogk
JrUucqcSamlVzqSYbSQaxZ8dJXXB7T14wODKGyPkmN7nMN5R0mMdWoV7/+C9Jm9t
`pragma protect end_protected        

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RigC50oXa3De7OXe5LYZa6MGFXgVfghBSRORlzwv8IDBG2VdiXlKzISkwj0fBBLJ
J6uEZ7C+sP15/Pnfx2ImX+WOzsMmPmwltJqxiVDgzokA+k8wGVr2i9QAqM0j78Cr
y/v0paAeGQTnihsVeI3DzTxvd8wCorMWUfdmeJFzl+w=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 40712     )
gStibPmMumVFkoT8vJMocYpJFlCms+IlSDiaWBdoZb938pr8hbv6jTRKj/QRSKyv
2YXD0i3qxOm/d0zpdBDZvxpe7JHic1xJtLV/2pkW14YX0MTJZmkbGsZ7v9WBZmVw
gAALNKqH8U21UixD9RzOs2vfNr+UxGwWjw6vLxozXKbMVjCN5Ekec//7CFnwcNeX
BuXRoz0auJdM804LZcRkd07mPKP8UEPB0uiO1MF69pkxb7bVxaPxNPCaiHEKd9hu
xUkVEJXi3DkicG4iSwlX9m6GlprL+7LSKIrp7V9/Hrt0qdtRmSluuG1lY1o1FBZA
A+FEv3BCvJck728EaMv6tgS6SL386Stung15QdBwwSum2fi0hgvQdcEVC5f9u3++
C2dojlfZ/zGISdKtzZE8fz5ZTqkwWPrAwdCTVMqZhMmylDEzD5wBgQK0sQsTokpB
W2+TVcS3toeVHt9vfYYcPg==
`pragma protect end_protected        
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
hPIPRk2ehIiG/kFahOHE4xsIL29wVorH2vv60cHe4ZRgS1t+RQAgqLwb5tkkKZIh
PmO1XupQ/pLh/rU9Q03Z6brqFE8F43PEqJ6CPtK/yGgNRB/OyPRUY8bCSBvl+WRc
/Tur1PYefO7iVvNBzXR0S/QTDYXsZYJ8r2ERFVX/73Y=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 55524     )
0/OCgEeYzf02Ty9CteoOJ3g6lAy2z3wvvLsV15nyPhsi6dfyDCvVZePvCHsX8YGB
F7KkenumnGL5i+7yJJCJzs8xD25PGJvqfIAdRlzGuyVN8l6Dudd+a7E7sncObWaJ
X8EqGLmfgTOFtP4H8yU1VdS7MUkUFgCmgiVxzewmxNQXDmpcYwgK8XySi4D5h+zc
RFBnesdVvoVjB36MCn/W87waD0RKQtMF9v8oJSNrEgG9tQ5l/R8Giaar0xuuZLCI
Bp28RkEPux3o0KynzS7q+FuW/P5Y+E1eyhd6QEOm1CbUWqptWNp76848zAQSZ0vg
Nyvq5d7N/pOucCgg3hSVUtucyr35m5W7XUdQshniTHkRrmWEmJnmsmsLNRilZQYm
GEAsIk5Suk9ZWOvI78H4DJWqAZ0TjupLYJvD6TuuUSF7n0z5taHPNoJq+wdh04Ej
BdA/EJOtLc7c67pCx8FqTJYFxrBpnbTx9e/RVs6z1MC1YF2LPa7m0EJroNQRwJ3i
HF0VpFocSdEEdK838nuljZxaEVbWsFdpjmVj1G4G8QDnbUEa0N8Z/KyVsZwnQODv
taretHWWQ9J8VUwSXNqnOGxaxGNHu8IE2PyTarUXWumEp/S5nuOWpjKAMeBN+JCw
SlpH3XtpcfowYw2hjzDrDT28XFmcX0hPYge4cnP5SGIBPl6uMzsyB4hbOcwDOGui
6xXF54ktUVlf7QcucjmJPauamx6XoxeuVV6M8q2y3dcdKdaaicEIS+4aKCN5M5Hp
aJQg/fMhyc7ymBuyfzfc84t6Agy5X11DYEy1Ak9nM+XmeUY0c9kwEYvrACBBmcTv
ix+oSkfnTZbpG9u7fB8cTFjbsl521ORhYbQt7UnaGW7UcBsmc1EfuJtrnYdXSUZu
qe24aNI2bMpcshIFiGTh6OnI1QUXHyuQPSDC9/lw0ppy0UffPD0RdApeoZCgqZIR
osYiMoPcpRP2CGvccbwg3LlbbzT5rw2Qd9yQevD7D1UCdpoE+K/7iywKmc4bwBDg
4Gt7f9dE9cva1Y4n8yJ9C1Lfkk2d6pcuKSM7wWfSqODckiMHcDZJxbdk1D3ipcgt
W4y1P35sp6mmydlIPOVfkNK97kKeBuaRkbegWYr1w57WUknYtRbhII6etu747L5N
uHsoyr+Q1cIQ7wMINSieBDiqDnPSV5wJ2NkqOyxUdzUkkWs2syHichOqjFrfS+X8
66njyRk+rc55N+fw+v0W+sMKLMc3J4buaiMZU+PtIuWu8IUWYDb+ah19NwNW3w5R
f6pq7JIO0zDsoaDVlTnBPh+dO9iSkk1z64Ie/a6GnJcbJLaqlzMdEiqOUbNitK0H
ducaqMcqVNTVpO3cMC4LdJt6njt2949HJIZAs+cP7bVuYzcd47CKkov6HbuSF0el
dgIS6YO4KHL69MxvPD/GFh85VrEJDaBV4xf9GcQtfZ4cOWq2n/7YyzWjkytSDzSD
rJ6sH03EYKm+DwA+3jRA+1TZiS2VAw/Drc/RXsTP30QPUTMHDEaR2aX3zLiuDksg
Se061538FDl5CyoGz5LmORaq6Nzje8+PF6Wqb8Y+fJL6whLYLFdaniYj/2S+EG+w
oeDQKccaeKG/C9Yjtaoro4X57PMyZw8t7vqGV87pWl8Y0lh6PqSJ3x6PI42slYJv
uWuAQKztW+sxqxlp6Xt2+dJklChuWS2czPUbinYbWfQ5DH05Y9PubYFv4LtjS4Wm
ONzOr97BjAQwrkogPFe6tDj0buBWtFUURjItPY0xQi9mJtwcwYj+h7wRRhvI68vG
imRZOg0vCAxx+jJuMMvgZGtvcdSvQGHuiUBggS11M4xoOWkbcQyFFeZnhuq6hJ3F
G5/hsH+tAFInY4XEci8UeAlnpFi75uluV143EiTsz3X9c14F3tB6T2pkfTByBzO/
3uMzX5pLoXqcYY84DwcAMBeBA810/cS9Nfw0ynBVeAGivSjziXx7LKQJS/ICPRVs
RmbrI51vaulcKZOWJe+G1sB+jLrVGEd1pznQnF1Sn7wZwrVnwe2mxVMQvMFgIaoV
FN/FO/c4OLZgz0mw9UrC60ymqeZvI///sjwDXyyWQIKIB8crKfXJWNfqs53bMPJV
//z8IJC6xGsGUIwCtrioLhuTQtNk5zdaQ1oVw/IdPFP5kCDzyPqjEnWHW63PgnlL
xwqkf3ZOt8uSyJV2g6eFiZYju5yXU5CpfA1jNGCBpY8zdoeOny96NK95ZRoX7tsE
plGwD7Z0FTJt1BjtL2X6sgWHZuu0xfeTVf6Hpi8PZHX6cHs2qJnsF0U2w8Io91hK
t5pcPMsGjoMjXEYd3cW66ylULT7zRX4RdA9edGCha+l6cQUVPELtMnieLCzwHIg2
mA3/e/SahKLhCJ4OP7hllcNR+/Sl6RgQ/ctbA4HD9ChGFvQY3XniIR2CHqj62jkQ
6eQvFV56VWesCR5daAdIT/J+qDVvFI0VkcCXp3Z2dXzAMANXiGIWpjLKTkRkJh+M
9BxAMb1A547EGShBR91Us/DAYkChIN77V5NAwUgRpXjb/tSL5hxsDsJvJ553q7g9
op3IjOXrKLLl4ugTCQj0Dnqd2Et1SHclKoJCYRo2myUk7Y9LXrJdD19ENQyq6eWu
zN4jmogMeTH0GBHZAzCVFPGQ47wV3cx+hyvUeHUy07uoqvYDLagc/dXBewUv7P57
4LoDBJpd1XlAcQvXyBwhIbK1TNti29L15NDP9sDGJ4thTKyj/MIM+jDEc5xc0eUR
hW0k9HCuwF+QwZ1BT33vu4tSjsfqTKalk5EB2KREOSkA++EcUdK1hJ3+YPIGhX4C
Xj4Hs1gn1b2/hPvIsealOz1tuNtqD50GYQWd9omoMwE/W306VvFKqD2PSBpqqlkE
cLQdsQ2F4K6YLONVQiq6jsLW2x7Qgjhfo/Dv7nd2UWiRtJfOZFndfBe+YC187VYU
myXkt5H7801v/xBoa7aa0tjhy0UB4lDND90vZCRA/BJy/MGHg2ZtcabmgOcwsk/d
8uOBx1B7BKpMXAMpZ1dg9uRSpXBbduVzJzPQDTihpJKDDgusmh2bRDWsQkNKOlzn
EYegqgefdLFpm3F7mIn9elyvkHaFxM2ZjB0Tm5EM/3tbGyDG7p39i8cL45aQQQX2
KKfMBg7WCq8gMTwz/QyorrqprLIKELOU8NKAjXBxUIFE153Z7uOhav13n4AQJ/z4
W+b/+4yMItXnfYBzBG7hVsjnHthGLae2p8uGUfNE/v4ggEAEEciKWjkNYsS2mU58
Mutjs0yljEy7XjJ0J5lHijAn9pzl5D5IVdZ9ImMr7QJdwnUwUbAqKPKsuKGKiZuj
/outZeKaVNKmuSPlfw7LCEpLVx+3TB8yDuEsMqUCihmcAUukDj24Fol1zOkmaoeX
HfhFmXuQrc9P6y7Hhqw5IS2g1fE7NE+UQDnX/qBktiOB0tqTDWUrzUOophO3Vlrd
rEh9WC5VvZiQ9qOEbdeK5xxE1v12hLaKQx0BrT+Lj4X/VbnwT8rUaZn+mWJhHTnl
kqWVuXz/nvg74klA1035UH3hg0Oj38lDjNSrBvKOoxSXawph7RGrFH6Z5JOOeiwU
CTI+z0tE4uotcx7QoPBIugmmEEHoKrl6Szv0Tae1LPZc9xPWcwtySPUyvnEK6u+i
Tein4Abv7dvCEjw9T2pm1fG7jJuLMgfx6SgLTRNydzpulp/cFXEzr5BSIefavqlS
neIBaO7odbtdriSa7xPfzG1s7wa/g1lrb0waIFzuSrJDKhcxlwkZToS0Eu5tq1M3
w+Vv4fgEvDd8VZ1L04J/PLwW+ac9pB6MoukSg2OulJYkcS5mPJhZToVHdjZGysCk
kngdYMPtRfb7db8kLMGbQ4nf12PScKt2rKd1yVjejEmek9vieUKweLh7VDvA8FTK
p0DmDNDECec30OvbyoSWhl13KBS/7uGPj5OONKoxmy4K4SYoMmvVt86fJKw4klPE
ylhNUWFz+2kvd8os30e5m1sgGriTsERlNRH5QkVVST55O0z7ML+pxatFpKjK27cB
9JDsWewon8ZU3T4LLfQdaEi4pw312sxzHEOvKf5HxUIpMGSqO7RnHSGionCgaldR
rcpQ+v6/XMywXcHcVOmvya9n4TkGim59n3S6/dmiYu6wg4C0XEy6PZapVB/7sMNN
fzmNwpyVYJiuO0ydV1SWondUwglyp0yDsZztQp2acwQBsx+gJfaXFfq/M5nplw3w
XseBJTQWvaKk20xZ3g2jCJum6m3YAr2NbDnhrsFVR0xp1itt5SBp6RBhbmEdGoaP
l27nEYf4PCudIM47BwGsrMmjjO+xKqLWNp26lXossjp3T2lQOdX4bg8/nJzo3y24
/1xNa030oWnVqgP6KkhK+1Bb3s28GaKoUSSYJBsiQvolo1N6WmWgjXUs0apf6kqL
D39788yxWZHWJSM+5VTKHx8oy/ZB2dV4SgBEHnbd+v47gFkKPOMG3kGknyD2c/Gm
K1LXLvgv7ErYOaN3GCLQ6CgAni7mSxJhDTTKS3jgnVBnybsOR9ZEmvYKWu3uyVcc
YP6NSLzwDb/kERj49GSOVrUy9Ex/pmL1/hMynNpsvuA3Kwp7B5SGp5RAqymL98SP
uL4zjMh6Pe7wXxePVkszp9iJCSSG23i333d95VEZ4fvPqJpmSQXaQ2iIqDWpUZry
MznyqNJZwoHnyeMw9MG4dG0CC7eZ6CwOLYSKtk/d9UtZxQrauTDf96XCIogTmoe2
TW3a1LYX4mn6Kff06NEprCrnJeJMg++EDhNLy6Q0ZQ6KDwgrUDE7T7Kujxkmj8bo
FzNgmf6TbC0QsajFxm2v7ZGyCEZZ1UvB9uinHWw7Cnl4pd0QAvO5IkvJkKrcsHJ1
m+m1o3fn+40HZG7NQaetI5xoSgIHSu0bpacahOdANHD2i5IPD0CdIo5m/rIRvAKa
ih5bH+GHJs7pECfhXyUoLMdZ+pUa+eHps+QVru1DKArIdyH7x277Z/GzWR87vyvz
rws6zVRZ6VhKFvWabhiajl60IWOEub4OQb96qOiunI/LhcDAoiCZcMobqhZNIne3
gef3cJP5YLhrnJH0g6ZWcrQivSU8/+iqho3IO6d6gW7f9rppCqpg5k9HSSOnMbj7
T5zq+Ag9Rsn4KYT2ves8c6edMqYTGbvZD6xidAv0Yy9vDGjAFkN5HW1pwSbvz4pW
vG+v9NwF+7nW+jGsVtIj7HaKVIaK2G3Iz/dkkL+2RYNnWVs3EiR9iqvF+G5lK0o3
LdbGCfZAHaVwXf6jHvzoejqOgwWPEUtbkD8GPNszGWBWZr8z+tKWiithVhcD5B0a
ExbtLLn/x+WOFHdqro29jdmEHw71RoX4aRhBN4LLGH6ZlwrGIKUECAj3/mywS0eq
ASFNCpZ608l9ENLUUVi994kFAeO4bo6OTqaZfogek6fGdl55114wtRJmnMnLZFnN
QlarfMmaBqrBDDSvCiHd5cduPJJfEIjdYnWzI2q1BqEGb0UUe7ltU/6zMKPtqcVR
qjjGazhtsKj0wRa19OkwAY0NBAAm8bgscmWYkuAgH+63uZjMHSpHrHHR3w8dDV5S
EqYqGXSivSGuoO8PNu3teXXVHxOySFTp/Z6N5N0I5bD9FaHUo1+FjNgjpzcCf7Ha
l7eH9P404gYSvNAvi2BLG9SjqDT0MZEqANFHrMJyEykqmPm0lkFMFJD8qcxUbbIO
GNFsAWAzv9puIHSh9FqH1iGQjSk6n5DPj/7mhJe7f+si5dG6I25SqQ4s6TuhDtoR
APjzKN1EONTVWuEjlOI4cgFwUoxxnRNhhrhjA4HnTa3pDAevGN6Mnuf4HCHb+cEV
vlPngTXAgNz16FWS0qMvezlGF/c05CUFazjZImnLc/j4SoHzGngP/F+u3fgHnQNz
eUUQEmSse0XcWvd1spgKLD7lmvxkspmSElueHVkvlf04oShT8hG8Q+Bm4mqHsZi7
doeM/Du/XrQF2QJJ1Es4GjnsPk0/jYgpOQXn4CSYyC2lLep7bCWouhY+M2oHXHsW
umJh7wPH472Wf6GCV/MrKCvYpLecYSt3HXl7gmffnjpT+f2yu7uNFlMS98d/9sic
pJ8aRZBB2Jr1rhD7aRvhAq4UfJFQ3hBXVHvtaSc5P7nsTgmlyVqXoJdpm7TS1RGs
IEITaFLaGlfvIjkhOVFj5KKrNktX12FHeL6oVOjRXFLZGjBev+VfSNOwAHKkyetu
MMKZQMR1n78FKGoaesAPTQwM9wOleF45w3A3mbCgn5zScWEbcHU4LRPMYSKLS8i1
IZSKaHol6ijXurLgcE3XArKrxkFtI0KCgiHbevthSCZslYWF1Wbr88DA/S66SGe9
Ucbl6iIcwaGEDLzoLHJWw6m1IJYslvPt+V1vv+gGnkMyWPYjoUWEst31fyrJjYna
a6n5P5mRwPGYFczgiSgQ1pzAVwlf1bpOhKm1RH88hle/EOO6dKEDUDUqXrsvT+ac
TONMjzZUv64mD/92BUKtwiac6AIadbj3w7pjJdu05LmWnGelXR7QxdQ3AurMN1sB
Clnh/swRg3gLxJKOXcyrng1TRSLNDWGnmNcDgCgIAHxdYh23ZW32zSK27OV2U9gh
EjhdZxBn3Rym7ej3+sP2MtQPv3SclyRJfnUk3BTshdrOB+jY0pY2itPMydC90iC+
w4iNuwevYikgAyu3WfSurgi/9IbDYvwxTCkAwx3+zrQerig5gMtkqqzbK96aF9I2
7nmEzGQv61nrhvnQaFoeOOMBPnhgmRyMx7Nc5HupfI9I97sKEifmnrrNaQVvidkD
JFqGpNIDP2ibQzF3GbFP3NMlrpBEFHj5ttiGb/1o0zKFRUJ8CHFCxtAEhI2yofT0
A7JDdS8TxSIwfVFdMaP/o0vUYPJH+Pcf0TV0yOoKU6Cw24djEOW0p+xr1dSCUp3q
LPce6UOMHII6Xy/qPWoDHucuTZBPft83A3A72mWHfkGvdoi+KdTPcQ9Dbun7RQIn
IxDsM5YwnY8x3HRgcJ6gEoLGH6wdEyH+0YS3XT3z5b418dhwy0kHaGrCn4vi9qzb
b6ntwjl/NIMdUAqh+sa4iEP/Lv9gQG5r3FSsOPOYu29XT052LHUjtBwstiWy3rXC
pFloy3HxidzHGcGGcSj6d7DmszJhM6qFEeub4Rbu49NmN2ibgu6A23eNYZ6bTUbF
MX5CV7swsACLUm6Fcdgz+Oo8feytwrsH5z2nFQn5/vArLCQiqXRSwbwwcwnxOVnU
Tk6VQRjUJXDSpMmcO1xhsB+2aPWGn3cCbBK82Mq0uoFqklAdI+ttbi86JALQOu5Q
t3NjiyB5A8fQnc75TQm9/69S4H43W0qiffYqA6GULLv7P7UAcEZVHzqvYOWBlS8/
2xfWhx0gMlz/hKEp85ev9vKqy+xoNb+JVT7i2p2UL6yJmQnPLQmFtk6EBeYWDmm0
pqIvJKmgCSoEdXtSP3Mw55dbVZA54CES/SnSVW6IpsgvsqTaaq7A8zqi39/4iWFf
Lz7iuiIrPCFb0qBijbRFnbVLyjwt3vu927c6mK7fPGbbmlP70keNZichveNWAj+m
S7ch64Uo0MqnFS0hpEyoVSCYEHwP4yCAYIZ08HwCyoixxnmoymFCm1LnYGI7r05G
95loycs/wn+ptleGeoEh/fxbJAsBR2TUm0VMLdWuxQufPbko317M6KyW9KtJCI5f
xagEfLpFxpaAFnewGCz4pv5kpZ0Xqa7S4JC5nLO29JhG6BH654ZJK3zEYGhmTG2v
tehPCa5MLyFMPeIrUI5E4YM+FDHWkOFaAv+ZJGY+T17WDrIhr7Ne/mlQhTFDn4z3
iy9lZh09Whc60afpbZZFipK3GItN5Ma6ZbYyx47fEiJtdNA85Xuh241XcPGJPdSI
6Wss1SFWPPvbmgc77bu5YArGOvQw8eYQbQwccI2nkP8JnIspsqTVX9PKuvYbO4tb
RpyAknnzW06fxRlIDFA8gfR+p3kCcPnGcmWunxipZSJq/q4tby3+TNEsO+S++Cc1
xxZoY5jNde9NYQKIPZdCkW5PZjVXJES97e7vhTVIAt8whJOZiC6aquzizXjt7pLd
gvIrRhMYQ5NZkda0/CULEaANI73jqajDWaHKruCL25oIUoK3z8Q0OYCGh/s2/NBd
JI/VaIQoJnP+ab1WXfT8cFVtwjGzOdw9Kn3FYFmYv+GjKW4JkprqjSUTkOUXtP44
Dak5TpbCGGFC11/xg3969RJr7pAFu5m1Tfr+pJwr3XXW+zZOJXJCONJDZpHMNn96
23Ak6tsz01RDa1HMXCfjJxvlKBAVNz1hulCUbtdyp4rnrBrXUFmzMYEhoHYcn6OS
08JdgTnns1nDJmSXDAQeATEwoVgX4ohqvZ34bZQsrQ0qAMqByBRMTblWDJRuur5b
lY1JsnJQ0F0OX7xwZUIFrZsI8/kBFWGvuAT0SHnnj/LTruPKBBu73Hl+OH9WtCe1
GXGS0Zn3yd6hutDICCcIuFaWKSsuh+NA9JlfU6l0ArxsaJJbDd9cF1zUM/I5W0km
6PpDbkyypZlYf6BPTilO+m6SdRKiJq2QF4CL3m6X8eeLnUwxXwBmYecpp1RTgZWI
DbtnoO1XKLG9j+z6m6IhrHgAtyPziGZSXZjj0rheFZlywz7B1LVJvtfwTBcdP5Ds
3L1o1NO9Bo+nbiKI9DU3Tx43o1U5kRsum19KzQXJ0qkOs/FUTKbIPlC4Mq/jMJxR
TSy87w1c94Wmm+OfuguvT5HGvpPD4D+VY1PEwsLV0BTe3IrjU29EMIFzCb3NW8V2
GCrKY9uoruHRApeQ4O9csEfrLawMEbQMK082vInQTu4LlJkMGBv91qzwja6hNzR+
GZjDE32xKUnx9Loo9Ed/VcbsU18P+dcYjh3RGIZJIhE4/x/nsgzV2MI0boE5qnZP
ZNpJWFi46gUtseaLf2bRfuPzD3HWEzECv8bfzcdlhXCvTpswEyazWxfRltFsN0FP
jv98/1hLc8dEVwEHfCARKu9kCRHs7bRuVKCcNtAaJTxs2/ObTVXPEVtW+eC9ULSc
QQac0EE+6sxHi2wJAh+o7cjeBTp6KF5kG+aJqN7a0Mkvhx7HH7bDyMas+L6nlKzr
7SGiwvJ9JoTJEIe/eGgfxMeAQx5+XoutX45YLlP3jmFsG8o35XtzXUQpy+9Tl6/Y
0EunxOxF3Y2eerIamwd1BjESaig16nnR1TKZe+q69Fd4T0aS4ap7wKV8CQ9cMRjg
6pN/TKXruxZRwxdUjOt8VlF94WzB1PViLoEpf42M7YaAQhjSf5nqSvlNvV7gupE9
rgT7PLrknBU5PdXZFuJoAiupqs4T5X8sAlriaqU0lkST0g0Tf/Gqa1mF667StiPc
f4zjcnm5B3CpmVOoy/TMZ1N3yz6eRNbl88NSOAv77nmT5W6qbD+KbtIbXjIX+eCh
r/XQdLfmyn+BjxmTQbKVzcT/VO7SIu5gAuh77t8JQJpvwb4ngsNtqkxsPCqdgiBy
XlwhUKCbtiMbvjsDAwa+I87/g/DOwvSlY4gAs61HRHKH6mttH6BFt/b6IHqXNR5b
2NCs6/BR1ARhrsrL6YDrw+1W30eej2mO8BBj7arasBQudJx8eqMmvozfDal2etxm
5yuC1aRJJ36SPriZ8Ikjbm7YglWVyfFax3Pt9kI/F0U5KQqRC80fai/63XGN9ZWW
ze87EfveLDtdsJau7In72IiFVwweWsg3R7FIOTep7DXIU0WueWBDofzNxm+IndH2
gdV96ta5Y7j6ZTEkVdzrl3aMjAamC8Vqg/qPZksVsGe2KKz6ZGqEUgH9TOgc0gJT
xUFTnG8nsI3bXZeogGg5Ys2DDWpJ+n/2lj8P3QYJR6UzxGUbd1D70A/G0MnBm07q
H934kL2qk+WhjeqEIzhSMc8fdrj8eQj1MRcFJfSf9fRmF8jjQQSSm7jpeAr5EEbr
+ZCBJM89UG1XZd6fsa2dWBYnS1vjeLPdpeGO9L/rjzL5DPHY6Pt+aIaJKIzfqCQd
YiBC4Rl0otkEXpSVi3/oCA9zvedTVP05wCwbXD0U+AAq4rU9sGY/v0R+r6QR9cjf
BHGULfa4wEXyrU5VCPACtVdgErKYFMhCM3Z159ZTNYGG1ajm0W9fKiabc/ddrEdO
UhTSkJkcRkvNOW8gZ1Y1n/iRNk+q3Sz1bMYKev7gxJSCuwiaI3hd7XSuhHN1KWLL
Kncn6bbvCSr1eXor/LOyQJo2llwp1/VUyJJTLwOlsgsJuMaprXFwm2Ox5PX4LLve
PBYFpS+l5E7515uxt0NKmmPlqtL7YysEII5MiaKfQoOGASq6ZCT6yxnfvnOK4wn9
org4b/4aMDoY+i/QnL5mKxcJBMzMy6XGLavUHxDYnH6DwTpwEYF6YvE5+T1uONkj
/JOffE8jsH/+ys2XZ/0JkHEVpdBg0X2+lsfAyOrqVu4fpCYmQvzNPt30Z9oIXqTV
hlA0CHkEJ1uSrl6qn3HmU5drMTd2wKR4jDuJC01KDIQenKqYDUDSUu9CTWQF8IOe
w9jVagJHVRyqGFJaR/rNdiG5jAngGCC6T68+2bbQ0Y7N+IUyK1rmm7Kng2gUaIWM
lbWdQfgRsJvA4qYpz1C5zS5t7vJ1Ww/R5WqD6ikc2Q8zilr7buCyot90cWKYKFKB
u0RNZU8ZPGB5N0ScvnW7m7LK7d76AGX9BGKw98j+eJ2yhgtnWaaaGEcDxS9ZSr8i
eZqpFNqGGPNp2SfheUFMcUeC9DDjOJrxPBJUwQlQFRIvaND23iThb/Dx5TICBRpH
C7tcwcrjgs9s8D0Dr2Ly8+Gd0UpITklkN/Zabe25WtB4h515kIzDPhYpdNEicyZS
ltP9gLJacwzNZV2kUyf0177J1Aj7Oarg0To/mkK8x6ERkgvJax9KngWPnDDhiuei
Cx61zn3Y7M+3m/p2f8mCtZz1I/RxUOvkgltAny4sbm+SUrOWNP8OhBKrYvccM+L/
Cqe5ToMYcvn87VbLa6I1uxpFXKTFtXv3UuW28OGWF3gEputs0ea7gfmLm0AmMHW1
2nGbmc8BpgxRD4iNoin8V+jwlHCADnnAZ6sx5Rs+OA/7MgWTmjMSmrU3SpRwTCEr
UPy2kFPrLYtUZei5sc3AQv5VmEj07XCWHIYcOmbUjp+3VUyJkK0ssmZhLd1T5E68
nKmgMIzJQfqJQiIXZW9+nLgYO5yvPxZsvcXiRp9mOyf4Hk12u+cZxTL2hi41jLvg
ujX8Q/uI8mqYAlPeCnYOmVqwfE5hXJQdFmxJ+K+2hL/gGrJ1qTDTzZ5SJ6ZxkMGX
uA/ozKEpUnLhZTNAHnVL9JzK0Px0laUumvrGddtgLXp6/tuEvQxYA89i5Y0w+nOc
emZCUW/5LRpF2pU8wXvHbj++wdAjbFurz1zcZE+2+s5LUIM2GyPojxqrJ1k1KsPY
c0tzxl+YaBsEjf9VzjKp1eIVFi+LvY0d4Xl0mSUzE1/76gsVn4ot62cJE63o6BoK
feiJEoUT98I0yJUQ+sP1lYvXFKhe4ioBBP2mibpkZFs09RQyVDlHLBmOpZu9Bm0e
RGcIYPYyErYw2dt5JwoDshAuFhlo1O133T5C4GqBz7GMadBZSspvX20ECnWG8b5a
a3HapzhCyLukif9/c8hxV8ft02EibsEbaLaIvlZ2ikj9nDjDByiuzunOz1qpTv/4
+6ueOB8BlNxczwexIzT6fU5pe2V3a69rewGiXGhFompw8MVKkIwv+BFNh9Fp86WX
Y7vctPHXvlfirtIa1FdbUxnMI0CudEB9dKKpTA7MTE93p1ouM/vSc28RVmUjkqss
s5/n+HxLBwc0FslaME8D+ySuda0cnHG61ViEa7gyHpOJptalN2IM245oG+YrdSNJ
vN6sOVo+5gxSu7tnzHekBan/gZ/xGbIA5LxZqMNko4NRC6XTpTvercxdslokH5dL
P2i1BFjTBplMjWXWe0ABBLVwl5ldnBQ79qALK98/ks02ai3yVZ2xxyaw8rJJan7L
8vWkoI/O6rx9lEz+wcOoCsOTQpuT1/qdlstirkai+Z3amfnLiaBUXWmKTay7tYmz
6l2fr3GIlexpmGQYDRxZhc9+m/7klqvpbef4wG6LeQ26cH2Zsf0wK5YXtbNKyVdc
peZqLpM+JFff70DOq9eIVzphDwFwh2PAAZdnwlseK/FkZNb9QJtYnYPvPy3MeLLh
Js4wHWcXhiKDbytpdvsrc52tNDnEE14pHOgskfV0NfnqFpWQAPK3hNW3aPP6CkHY
MoqXoLReP7aBc0ABTnrHvIZguI7NFZm81IJD9ryZg3Wtui0x/D5fZznpKNHI/xtx
tY2hP7XQ6q+CYC04DmruYPFCbUtKU7Pyp+SPVXw2XRS0OhMLvj/zK9l9zsX4yds5
ZZ3mc2Xh8k0ZqMLmfEI4JgWHDIrE8uB2MTA0A2kFqzzl1j8BRCzURFXJl6+j/b7i
8vWu1KdJ3SPyDzgWfpOaW47pX2flQHdLK/HkfmfNL2TYUsyBdsRwpUN1kZxRTjTr
5rrlnX+UFG75yYJcj/2UF0+NWsrpqdK73o+bsUPWVLTmYL6Nbj0VVzslyz7Na8WX
TCmK2QJSJMj7CDxwq8yM9vaAXSy1FInw5+UCuGCxZ+6mXA+p8FGlky0lio1YphMe
kYTdSGit1aGPYvDn6NREaNliZT1Pked4hQZXTGvM/fK+EFimG56yPFEYh/t1ItGz
jiRnHnOxeZ2DkKslp7//z5Ii2iwzTbfKRV8F9lf64xXWbCBrzvcbNpL7XVSSMXUZ
dR1Rc+itoT0+QdEZaFcTsedhRI00znLZJrELKG8LEAlcjTrYBvf7aKtwvYGkLWcQ
/YfPn/IKYcaZHwrpZ7jpLvlLSMuHR3vNGuafP9KHx+G/YzZTDOBST+/TEyCAYHJP
9pa5c3fnXM+KYFiqqekjeZVfPUrVF2cjWUi/P8Rsy9vWqGTSVRG7TIbs4bjlsqxj
E/2l1V3ct69B+BkMduITLi4qHmSpyKSga/XnFBeHmwOHR9Piz4MjL522kfh4JP0q
NGD7ltlmNQ/2x98hho8tylXN/iJsDIDj1OAftO99m6b37rqCqkQLXxrYy24XRM9W
B/dJTTf8zyR0LOQuxSiJZ5CUKEGIX6uCwhPvNFntAhVwlHRKKkJRIQ5s6lqGms2G
IcfvTbldrBs1UK8hCnp0Uk/42HDlX2uU2JzcPhRMzNL1QhQrk/nuj89K/RL9O3uT
K0a86PZvx+20SNOHCGmcXihsQvvO5LwBpHenN9g/D8FRUcqDDA/FnCkfK4hAQwz0
XdduI/L4TXFRGuVle3cp6ofiz+Y8DlJHu6DF/pGNPYZKhtCn2fV8ErPEEJSc1iKR
mVck22bjDGCwsZe9nc+SBPBUzhmi3j67fCZmLlXuXDNxq6KhecXYh3wJ4Otha0jB
3s1QVgDBtjpeysltHB34CfXLVC7jV8s7BuL5J0uG4OO90nLAWCNreOScVvKpamp4
aGTL7D3vYqO/L5Vqa272OTmSHDOVte7N4LgCuxDfzDtjQ9DOLRNPahl1mtsOqM5q
oW4SxFObl5McrvdLjAsqVc8txPVoxKHXJeoy/+vV0KAxgTuihSm55rXNGabGPOCq
RAh7HEvo577rPedAxGrXdkQNylRKh205jr4FiCyIG9gpVmD1Cg2hyzUFCR9opqXY
6yIyrmymdksW7vuSrfTYHM2+BaNalFr1DHWVt2Ctzdavadunk164y8DduWVn8RHa
4iJfaYEdCwDTl4QDwoJIMxEodAlvp3LqzCqQWWPdN+yQGQpZ74zADTvfWiacPZu0
ITYowFrlyclDkukQd3EBQnZFkUU8Xe4ferVJ73HDJSHefZ9APnjjjJJd/ikUwuiu
sBM+8gtkb0XuB++7fG/T8OcPDzn0fYUOqAi3KggGTiyi8ZxS6wJhDCtJYaTQuDHZ
/91CtHc7UA16aMnlFl3CvxA8wtu6+X+NQbSpzoIXg+7/YZ+ZSgA98+TBaWZGSqjo
injRAouRhvk4sS0YQISFltzLHuEncTC6FZVduK7djK71JCQRrCwxC/X4B8yBOOmv
R5PRFXvBzBBVBFM2h+O0Ra+qIOAlkywUgNk410aQ8Qzm2yllcC8cf/9HSogcDuxQ
xEAW6QBkC8OD8Gks9AhAZOeiNrfOc30s50p83hW5hiVwkXrhrjEl823dzFX5uoAn
2t5V9yx59wFRBtvqCu0EiNqt+38X+w8PgQ1c9xeYoSZp7SRKpPKIqwHOxf4QaIl/
Gl1laNR6fBpYgFHSv0Yaukbf0lWinK0gwzsF+SZIXmUZWNeaFIad3wTpUcIrcWQL
uzpm0WwKA8RwfCQa2gc0xTNELS04bHvoyuu0HpswgjFb+zaHaS0GM+3BzUhYj7Dr
T88JfoAHQk9yAPOavdc8FX327XPCzLtg/UmQuuY7LnWmjqsqXLzKF206VaFidRhp
8NjwTUrkZv0VX6VTUmdb6abeVdoC+6LZRrPujbjNoWYPC/Xh/xwsKItgIJZcHFxt
Y8taeCv32+qMf40+CXoUPRYiqzIIElPxydMgfgDm/NOgkvPC8g2p0DhOUCaonLnp
/0wKqeO7UkaL7XW+5tn4iZZkLPGCEhkUy/td4uFUC6B8G2hRfuC1wItlGjJKbShf
aMBOUrVPKvpsxDgRHh2aQgvD7k/iBVJGZs/6ZHYH7ZzwySlHuOfiWXPczNxBlyl/
56aldKJI7aGG7UI1xDJD2g7Og929e2oecU0I4QBN4w2ZHq6AY6UBi7RiawMzScwk
9OHxb6nj8CeS7lMUtskrPJZWGPLe8giSO7sBexlDmJOc8D+Vp03lz9n9kTL3ZhRJ
KgHGholBo8GTpEaNspdshMfl6bh/W6aiZzwaAB7FgvrY9nC1u1Mq2XyvscSR720y
27WULf4Uj3f+eE9ASPWfX2nUKjb4Oje/4cHZLHZFd8wLlWc3v6VBV1gf7NLt3fJL
sRGuEfVuDT9WZYeQNAzKNOluC47HjARvL0lGLRKnbVSNKX1STu1k0ueuY/ctmO+0
ZmIdajwu2p+0wU6aTCDEQ/m7r0IVDEoeTDP3V1Am08zNWTGCVyj2J5jnBbL7gUKl
L7k68LPaNE0vWg+3brTSMavXl46Hs/jNOXbvpfH3c55J0BUA4LoL6ABQ/dXH5+4q
QLwxvU+JAMSgVu6w+L3kqmx46bCAALrtGgfp/sMuwL1QL+2H+xFIQ2arCSOBCgoQ
2aG7vmxGtUm8Rd8d9cC7/rLRJpv4tGhnoxKxeifdU10uZPPKVk7mSAKlknsQZlZ/
9/zNSi5HEr0Qve0WVagUdiGA7aqhDBi24kC4jdoto7YMdctkABKzH3YBpRz+xoDR
L8fkiVHMU9TTKu/L5Xt/K8h2D5JemNFtbN945TyoXkeVFEDpOUOQCgPf6Z904Efs
r0haIEdiM9j5Mm99LPi79gB3mIsBznxEEOX6Si2ohv18O8IW9FpVVPcEFl88vxfv
unnvSfozQZ7ILcJxAiR/o3MD3zZQwQt1nCg2y5CO+Cj+xeKadrO3bhbm6xD/Rsh+
LdZQ1HJxBeEF5hB8GUP+AhdvkL83XSg0aG6Raxg7BEAdeZymN1WmEQgsf0WIvoLi
Xfdj3C9XKXp35oDPpyyrz4GiTxCPvifO4FMoKD8Qf1sOO1H98Qr5mVN72EfWjCLX
aEU1goYWqgl9RiJudj1XA8PrITFrilC4pGBiHlgoSjjdbamSKLaMglan3RsqBu19
kiSH/+qqxE8CpkdNBFbhsWm0zOqbUMYCKzDIVal27rMnbj907GI/K4XZttkxaKfz
/B2TGce2DDC9vfLenN3KnUwbyatQ0qc6bMnKybsUX0NjW/P7N9vaUXvPw6nAcxn+
Tsos1tS921CqmAFj4aGQVwzvtjI+rpP8n7Hrdjs4Nas42zD7stCgkdAWJnS0CN79
hBt3O2bgelG4TyLZp7o1C14HbegxIKeO5DD7ed/qcXmzT3FmVIatYMTYd2l4JkUw
PtxB+psDJA42/xh2EYgONKHgN9ATh7EwG+dEy8VKnN87gYarOus5kkap8jEAyN2p
FaeDd2fqsGTVNCg3P4iCpZfyRjT9vD7z/K+FJbOah0oMhMyBvIgnfb/EoxOJLp7K
xmt7zZFyuz+YZydzOgmGVVgwKbeRQ6BBYWobsrqSo1rh5XImS9sQ+9HMVZQO2Ck5
Bv0WThbeMIRmuIPXeo5da71nvnMDLGTbtPBUwSIO2sQ1Q0/0oSiGlK/F8k7ubW5Y
NF0WrvqJDKK0Z422+5pv+492251ePudA2CXd0Q34rAzWE7wNEda8l7RsBv8PEsRf
PLS447XSv4lo7Evl2jGulxGdpPCgcRS1NlncXeEiDrABcN2a6QB9yANn21vNjsiB
FQxK3d+sGtDmQJ2rbZcR9qIQJd2XYiZIQJA/HQnJ0LkNoD02jkDou1aPCz/Z0GMn
ANNr5qtk/6hY4Y93D1LQMmTmHVAy9HagaNpKqxdyL4UKOa+pgXUQaNW/BEx3BCW4
XxtkHkyk/vdKu1PafVbQ+W+h0R27H2gf96KFGmNSR68SXAqgjqjs+Z35wbXG0mj4
1LZLLzqe3QQLGK7pgyYdX63aLF3yuhouLXfp31bsdEWYR1SUrYd3RyAryyXQwjcv
SoKbz6DKpe8qdn2IS3W8txYP3ddWNp675RD9O0TTi7zBduwC/5kq3Bx1V1HaA2a7
yuA/Eh1eUiUL8y99kDV+EijEpTGWqFPFGd7Qq8neWfHjCctJ+vKhHlftDu86QHjA
Ob5IG6H9CDf+0E2PcXTIqxzGryMqb4uNYnJiwW7+uNvOfCs6e2BzR/27c3pTY6EN
U/7oUOV8rcZtqVfI5JmjQI3CydLTjJFXQQshiZmVWHL2LOWTRaXE05xXAeyf0vAW
PSUV3WHiFJx8RR2Qo+DaiHOxgSyXV8sXRcYCtMQ9MA265ekNnaKDesUNuEcX5sN5
ZELC7v9kCEEtxpU3Sl29e7dO05E1lSkUAVxkmOvr2MtwBdnWhodYaOOW9Ev1IDrK
yFWbBi+zM2OWTj2WB7nBUTFViLHUpL4d+RNgxS3Q1PJVsvgEi9B+gLz4w3nAySGD
NGDSQ1Qh8DD8djYVsPNxtNtPI/S8WjZW9oZ4IcGPi0G0BscWCQBUP6G1MK75Nkku
uXmO+vw6ZYi7/4QISWxHPDAOlVZi8b/ipt6tVeetY5FztyKmaaNkblBT0t46rGMq
6Wz04R8mreDZm0bojr2ZnWs+DCFJWxGT0fnkIoI5MLuQeqb8R8x3fFLD6fDXdZjZ
2OSgvkLksNlNEJPrUErhAJA3IAKbAhI1HajQKJrHXr3y9ae1TEQV2Pnbra6gxpWb
mG02vglVHoFtssjOt8raRNaQRK1NwYhi1AfJty1GZD4ma6Cy3gNjXY78iteF9Jsz
wVN+a/S1f74c+P/RtmGOCAQO2ksehU0SNQvdB4NtjhpPTEV/UNMgRw3HjaB9TuzS
gmIatI5IWLu+oLC91oVozJ1aqHVzEz1orvgD73kRnNcxnr+07Lf1ufrEdZ8B1KXg
ozk8i+ta0zI0Y2Dd/kk1BjWXJ63LOikLGBNgStieNAX4EDWyse4WZNv45JBycTde
qPV6DB5H5NUuO1r88qP2zQFMP3mmyNtT7IENYMbR/Oe7HNuai24YCJlwMXl/UotD
5qpnGbGGytnHueYU/oqSCrXY/wQSR0G3humkB+nz4eFAJC4pSOdoqh4DDvsilHJQ
VbUwhQu4kSACsEBjsESSKiHPsQZK0qnjgaqS/JKbBBOSId7iTgwsYdnHKQDgpkSU
exPu37iogwRRNRu9Ng1hf75XB6QRTGLxZqjmR2jNYfMgThXchyyDaee4JJaKp9/H
N4zH74exhnqjbf/W2cdmglduPdklEYKzMQZlKPjEFhMyMCvqDrgi/pLHiqOgY8pw
EPUcqSR9Z56OEKlCm/HYiwc8F/oDyX98YRx8haWjyZwhF7TzESRFgjBeQgzUXt4W
ooDSwUCdw/cKpsoqr6c07/uzbgKj2953GTf9sYzIsqjMGJQj51TT6xhLeM0p0EiA
Q1tJiAZOsPsA/KiRtPsYewb40NJEpaRd62MZytXHi+jxbHWNnof2FFO5PXRuU0EW
+asiseq+BtfpQVp2JwgCk6lRlkVleQsvZpQ4LLaAz6RWsoltOh3Kas5u7Lo83SB0
61qtv8mX2gXNqhOlomAtBAlh3UnbQs6doFhonD3h9q0OL6VhbODfXDurX65Esb+h
dsGeTTSjkhVRgPUd3qokUDVpxt5yBxbY96Fs4XbR2YhOoLYKiP98xdULB1S3h6vz
hkwEV8OZEJsxMBvItU/EcSj8wDhC0Xi2coYM1xhhs4CedBYZkjEDsgkKKgK7ohTz
xYMEYZfBb9ZrlCLVg/caxuSN8KUECkwzdNit8dctXuZHLA0UIwvo8KhMSSos9mz8
U7oAAIBKQCuo1JXDo9YV6qP/atVt1ELufOivygfCUlpBBfpgIgnt7JCGi9yvNpPH
HHbxUV6cjsnqcPdl6t+62l5b+yNeMD/fowTBXbKxSvMiincWMYeNcGu3s4aCBbH1
D8L+FmltyCZamrNRF/pebepSAJZdgD2DWN4fajhBFNRRGfRs70I59nw5LbpIE9i7
JIIA5GZlFd0rriRJdo8q0wkCQn7c1ImrbbFrDQ8a4DPSKqFkGL43o4un9RwncmnB
otu6BA+zRSlm87KSlo1Eb0EmR535cIaXW5OZDbwwc4PkyYiyvuMKSDB++y9T8w6M
pt8k7vXxNQQVVrua0ZHonpqA3uLDdFfsHOpr7RNuA3nxpvxC9zdlRAvT6UTeUOVL
8koM18lXlmTs2GzcSRWOTnyc+CFJlvAMdk0B6BhJhR5oZZIoQSs2TA8vX1DRrydL
UJQGqZhVNXTjMXULI1WIsQnHxmwGHh9zkARHVFdhOx5k2A49KJIRAXuQFB7RWltF
u2BVCdwgA+FzDJ/xgg5yJz01cG5JYa/LLgol7oCh3+KpdelXbTT/Vf1+qAfOCOBJ
kKkJ3weXp3rRW5+ehQraVWhc7ygEkkO3aqxc1E+qV0EiQ5HfxEN48z47Bg4sw6To
baZSlLvyai6YeuN0ZOVsrTP/rkcxNx/GvZM9RnY2qHMPl+9pnDRIv/lWVk7lazAu
1ajfrZ4spGAYrwem9rYBGkTkOoEPbqj360dkmoFxTzc+fxM20hvzMKYua46uXKFb
IN36sLNrJPY6acLk4rrc13VDz1AE9PPS4yJW2Ywb59oeDR9R9KDkcoE+UeiGG2Hf
63RmyqCRvfQqv3DVh5eEoJ82AoyhIFTrpQ0cxBQTZ6sOZBvnrSLLvl46f5JsONU/
Ss1+bySmOnZgyNt1noWdsmBX6xSfFf5srwUtIC2rT+FLuQ9GxQafNLj+NutEQUaz
3PNIBbQSEGoPlhbLwO2mjJD+a1VqneEgoGZHfkZMAqhg1RlA/Xe3jBa8TDCU/XCg
LDmJ4hnWzS7MMMOoBbs7PKERwxs30pJ+pz476v3hv0On8RkfOo1mFZflInPZzytt
BWrXvDVxp6/FB7jGD6fCXCUl8T4J06a0dWsIlz18IhO0DN5JGsRmUlURiYbHl9WP
m6zLUQaQ+vPDRKWxtl6+Gz5Z1VgJt2i1LSiHFYABMLd3mcvTvohBthj5v5+08uDa
Vd/pkbHkGyx77MLaK5bdgAdXTIj+bCG3zTg1DKoKrlmCifM8tWznCoMR48OYF80M
2VfIsueLOR4dyl07znxoUbyZW3SF2OUQ1CMa9cN49f2LR65hERGwL03q4E1lmxxh
nkS+3m+simuYFfxYNqytZRy7hVaMEPG5DEtzwkM1rCc=
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
fYPe2mcuS/pQtv+1F1eT3AohnNRrfymKavxZntC0FvlnjEHqyStnx2k9lUXO6u9k
OThxobnOF7MnjOPl/OmojCSMJZL0TgWIDo9yLyg1xnA4V9vGrseDQbD3zWvS5QuR
/iO9ECgw6o0HW4xzKcidE0QB9Eb8wo/bKv4BvigG+MI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 55910     )
hAnmvvsjBhqxgNLjVBf+I8EAE9FvgDNFAbwNQR1irl0PsbqBUAXdcf39IPjttCgm
oRSaWfoJ0pdezb9nTunez08l8YiubFm96rl9Q4Fs3iJibOnOc2lpzas4NE3KfJyb
xvXaOFg5il4BXxm0bv+nFosMCJN1zOaXTFfOEU80KSD2685TAqC2gixoiLnAVUBP
NVT9zQwf/0Y+hhZwc3TWzzcyB9PqNQh988SL0O/tGdfKADwlBGOppNRwsv75B49b
4SMr22Q1Ftn1fbcgOEOJjvXz9MWEeHlAAHmbJcNgginQ7e9gE7YM3fJPiO3wjVqs
GrnFg5ZV9TxdPMgLpgKeEP5X+B+Z1TAGJkA3u8SZjRBWchZKBPYs5KXXIAb2k+5w
kwFYLTOyZ9uCXjsIxQCqmHxTqF7rRlgsI2xU1Me3Rt/p9MV64TFu/BmgPUZ4lFXh
KVsndYbcvc+sttmwTCRqjlWIiVgOuEe29J2pHcBYQAEdBgqu5kRruml6IQDlkv1r
Cg/kHxiUIE2WPeS78IWC6Q==
`pragma protect end_protected          
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ip08lhIHz3zbXxxTUNa0FoV2Db+CfCVYYpbWPGhdOiWM6oisMrop6sqWxS1XunII
sUg1bAWQnHh4N/xEk+9SJ4WUFvSv9ywMK44PrvgP1HQ7aKZ9WZnckrq0Fw8jVRuL
Viykkblmj2OEMhLC+vspjmHtHbUL9jcEpKhQAIpZTMY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 56207     )
7lpmUOP70H5J3FdUxAE0KLHw7Oei2qFoqlBDG6sAU9Zl1/G69jbQ+TqsL22gE1vt
HMrc/iy4Yc9Ri4gDuUgmdbhxNwHcI8tpe5Oz1UccPexbIQlQXskl1d50na7JjQ/l
3A4ULQVtJ5P3HooEvNIwmN4E43XWlowKS7DG165BpQf65XteYzb4SHTd7CZ6vIpt
+bW4qQptM16Zzz7n5ZnyrlwMsvUhkXmxiUj1BcX19+xuEwsZNJxjdUfizhxCsdC6
EEp+MHV8LVI6m4HmiV3UgDSXzoqWAnNllapXhFBdwUwP/7uD6h7fo160qYyk7BWn
j/jjunJNQzA8NH/TEwIdA676hsL1fOrG2QSFTZUOKGiGA5z0bovh+glg//WPpBgE
IjLUKFwDpfHpvAuVzZwFOA==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
dIP1Dt3Ad12Tns65mKArJEyDyxAzfk290jLityW920bAyl/Aq5WNe0li1ZW4/pHf
Gq3bQlDmZD0eXFLutnSqpcEb70d1/7Qz7JOiqOjEXvj0xH9qr08rBTdYCFqczvT/
SDY/uFcQhCA3rQ+88rHIyK8BWE25bwAieMvOEHf5d1g=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 56558     )
RuDjPt6tlL08JIyMqd2Hrz0zHP6p0ciMWJgIyAXQxnXDdlmVmCKulmffIQ+hSGvq
pc4b6M46G8d0ew5+fKO/8eY/w0gSR93EDAJspdCsY6rfbh/OZsysTxJ+k7tK1/44
+DeG6a/F3epe10fz4Ky6vi4XdX1x09NRVasYTDky0cwmQ18cmkQpH9MFUqboYJer
PqJ+DzDkT/zHekGSXjIMZxNVROgSMSZLxceRjb7G4/GqgqfRoTQwrI54ejmAaAdy
qpAWYKAm1YpjS9ukG49S8Az6tYZ/TItyuBg/JAeg05k8ZoKqR9LPhpMiLM/unXmF
qJYo73BKtGPnzdOvl/wKT7+/H1XFJ5piN04S25AFjN+fIbplRkhm8VgiPrpYRtpy
Q2kldVjiri1sXVMZHOrRrWbgqI3EU91keJG0QYPnqzZ0+Zpcs6zgGG44ucBnFAxy
lBBRdTAmhUt/hHwDVy9N8g==
`pragma protect end_protected        
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
L0szKNMI7x/shd5+2P1cpCBZwsB+Ea7a1lBVtLAkG+4C6EbKPOH+C88cwsAiTeRw
x2zb6+OqnPqTLeqeithaLUpEL+SYA3oHWxYHS0SXiJaxqBokiKpAco+bz1ssy1pT
jd8E6pF7867gdyj82HqJdv8i4Cry4Klgx8snSPXBSjU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 57653     )
qbxX+YUDywWuew64nDBC2WXkjE5ABzx7Y6Lpno/3ztaTiSiTf6d3KKG5lZTOp3XN
7ko4ZQINX6LQZk+HQ3E+RXoQh/dN5Vz8rfrXX4yA//xQsxREs+Q9JrJ94xYceeqC
9UsJcziiwWasXXvTM/tvUAWKeE65b8wKETFvzi6E9Rk2EGiSvlX0K3vsqNWCNrHn
5QV7ODPdOX8bLrEIdVfOL4BsFjZiyhiYH2xo5CVkZqhx3MIFxgyN7pWqmmkPEytL
+4DEQHDLKsyBQwSxVNdH8TRibqBJf1GgH+/YON4Kc1W/F0QNcCnY0VuUKdLD+MZk
bSQIult2AvM28I1abuPUkbHLzzQh7F9GF6Ji1vox6qucqcxc+rb7oFMbKJI8+/Oo
vGyOPtMnOviKfEvz3QulJY4KX265Egh3Yy2aroardpXoE5T68xxQ1kjHCsWbeUjy
HpHjbLh86P01Ami7D3maoDiQ45W1jG2Kt1/gIKs2xf/OLiCYrZE6jYPibBoRYhSr
jRIIphflkgXdfFOqmWX2cmb9/3DoQedlurkR/MiAuMf6AwckOKXTHo2DX2LpdTIj
jSzGNI76K7UPRrvwOdnns9n+W5FRn+h8T3/C+xqOc5d/WRHjS+4RZrk7ClKeKtXH
nMBnabtobDXKV0eSjQutfindYMelQjfJNnOC3PoU4vsF5kZlBfNglBTroZ3k6XIL
44ll1ZpUGPgB+Zw5blU1OLHO85e5LkV3/m21hvpolK/rw8OjP6MUQoEceue1/NYF
wjewFR20gU06wreeKwJalDV4tkxK2Zlk4p5mQJ04mpcK7iFB7ykIRyf/37tvAKdx
mSS10ErFd0vqODeAsbEgVAXCQEUnlHgW2hdrRLzVF8kOLU02L3qxIcno9Xs5CrT0
gHx7XSX8OkJXhT7at+JWJGHxiP1evgEmnXWG9vFpZN7EfHRyko6JV744J5nNfjTl
dVSZAb7eyxpZlW8yE00u/qfEbMbalJTi4zRO60XP93sd3N1YW878tssQZAgnGynp
DCF8CatUfBEmZcfyR3Msr4vAsnwB8CrtVgRLCwGaQwVyyVAFa74w/FtB5MBxLDpP
wsF+yjyhzpEXX+2YcWQBos1GYSrj+WMS/OASp73KAvZHj+dQScuizfZwBrZbiMiG
kXvYZzWogD6RDrqhrCxBZzkXlgXa7GanexcFh+oDP2Mnk4Z9Nsmz1te8J3N2ldbh
dVsx2jiRCVcQkwPxaEwYcVuYbiPC+xk/JK4PsbZJiLLuzkKKLzDQGP//Yhlf60II
zVlcwMrdc+0IZgqd1kqVX9gQXzJPSuOQIgn2m8ttwVDbc6ZBmQOe92jno21eQ1fX
5KPrXxTp54gXc6EA9zptRWKsaFbQV5c8rB14A5agjzC5SuNdXiskiytzbDriqd0d
c0WrKlw20iJbjYGIXBB+I4cxzuW2zfnr152s3XK3BfyxDwS/vIwUPwmnbSxc09uC
`pragma protect end_protected
  

`endif // GUARD_SVT_AHB_SYSTEM_MONITOR_COMMON_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
MoPYi2uWaGkMG8sHGNkPU8oo0qSDPbzdaeIHfrURinTdoJfge7BBjE3BOhCfgDI8
2g5dPPWJCEo+9BXW5ErwuSCcL8LJbu2AjTNBIhPzAUZLYWxQR++opx9x2Yg9AU3G
nlooQC7CM8bsJXFjo0JmBPOdAKHGY9cG294PMjfCXeU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 57736     )
LxlaRbUuN9BbgjksS/8os8W5MGrrN8/+QoVDM+HvBJzdb0udhEPbZFaJUPdRRrqQ
RDwBYNVFkTwUTQOEgwnKp5IAJjgH3UyG0Cg4CeFnkHPnAlc1lQWK24m7Pen9tXzS
`pragma protect end_protected
