
`ifndef GUARD_SVT_AXI_COMMON_SV
`define GUARD_SVT_AXI_COMMON_SV

`include "svt_axi_defines.svi"
typedef class svt_axi_checker;
typedef class svt_axi_port_monitor;
`ifndef SVT_EXCLUDE_VCAP
typedef class svt_axi_fifo_rate_control;
`endif

 /** @cond PRIVATE */

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif

class svt_axi_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** Analysis port makes observed tranactions available to the user */
`ifdef SVT_UVM_TECHNOLOGY
  uvm_analysis_port#(svt_axi_transaction) item_started_port;
  uvm_analysis_port#(svt_axi_transaction) item_observed_port;
  uvm_analysis_port#(uvm_tlm_generic_payload) tlm_generic_payload_observed_port;
  uvm_analysis_port#(svt_axi_snoop_transaction) snoop_item_started_port;
  uvm_analysis_port#(svt_axi_snoop_transaction) snoop_item_observed_port;
  svt_event_pool event_pool;
`elsif SVT_OVM_TECHNOLOGY
  ovm_analysis_port#(svt_axi_transaction) item_started_port;
  ovm_analysis_port#(svt_axi_transaction) item_observed_port;
  ovm_analysis_port#(svt_axi_snoop_transaction) snoop_item_started_port;
  ovm_analysis_port#(svt_axi_snoop_transaction) snoop_item_observed_port;
  svt_event_pool event_pool;
`else
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_transaction) item_started_port;
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_transaction) item_observed_port;
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_snoop_transaction) snoop_item_started_port;
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_snoop_transaction) snoop_item_observed_port;
`endif

  /** Report/log object */
`ifdef SVT_UVM_TECHNOLOGY
  protected uvm_report_object reporter; 
`elsif SVT_OVM_TECHNOLOGY
  protected ovm_report_object reporter; 
`else
  protected vmm_log log;
`endif

 /** Handle to the checker class */
 svt_axi_checker axi_checker;

 /** Handle to the port monitor */
 svt_axi_port_monitor port_monitor;

`ifndef SVT_EXCLUDE_VCAP
 /** Handle to the FIFO rate control class for WRITE xacts */
 svt_axi_fifo_rate_control write_xact_fifo_rate_control;

 /** Handle to the FIFO rate control class for READ xacts*/
 svt_axi_fifo_rate_control read_xact_fifo_rate_control; 

 /** FIFO rate control configuration for READ xacts*/
 svt_fifo_rate_control_configuration read_xact_fifo_rate_control_config; 

 /** FIFO rate control configuration for WRITE xacts*/
 svt_fifo_rate_control_configuration write_xact_fifo_rate_control_config; 
 `endif

 /** Sticky flag that indicates whether the monitor has entred run phase */
 bit is_running = 0;

 /** Sticky flag that gets set when a reset is asserted */
 bit reset_flag = 0;

 /** Flags that is set when a 0->1 transition of reset is observed */
 bit reset_transition_observed = 0;

 /** Indicates if reset is in progress */
 bit is_reset = 1;

 /** Indicates if synchronized reset is in progress */
 bit is_reset_sync = 1;

 /** Sampled value of reset */
 logic observed_reset = 0;
 
 /** Variable that stores the exclusive write transaction count */
 int excl_access_cnt = 0;

 /** expected exclusive read response */
 svt_axi_transaction::resp_type_enum expected_excl_rresp[*];

 /** expected exclusive write response */
 svt_axi_transaction::resp_type_enum expected_excl_bresp[*];

 /** flag for received exclusive read transaction error */
 protected bit excl_read_error;

 /** flag for received exclusive read transaction error */
 protected bit excl_write_error;

`ifndef SVT_EXCLUDE_VCAP
  /** The current fill level of the READ FIFO */
  protected int global_read_fifo_curr_fill_level = 0;

  /** The current fill level of the WRITE FIFO */
  protected int global_write_fifo_curr_fill_level = 0;

  /** The total number of bytes of all active write transactions in the queue */
  protected int global_total_expected_write_fill_level = 0;

  /** The total number of bytes of all active read transactions in the queue */
  protected int global_total_expected_read_fill_level = 0;
`endif


 /** Internal queue to buffer the incomming exclusive read transactions */
 svt_axi_transaction exclusive_read_queue[$];

 /** Internal queue to buffer the current exclusive read due to reset of 
   * address by incoming exclusive read transactions */
 svt_axi_transaction exclusive_read_reset_queue[$];

 /** It sets ID to 1 if exclusive access at any monitored read location
   * is failed due to current normal write transaction to same address */
 protected bit excl_fail[bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0]];

 /** * It sets ID to 1 when matching exclusive write transaction has been received */ 
 protected bit matching_excl_wr_id[*];

 /** Semaphore that controls access of exclusive_read_queue during read
  * operation. */
 protected semaphore exclusive_read_sema;

 /** Semaphore that controls access of exclusive_read_queue during write
  * operation. */
 protected semaphore exclusive_write_sema;
  
  
 /** Timer used to track exclusive write transaction followed by exclusive read */
 svt_timer excl_read_write_timer[*];

 /** Semaphore that controls access of perf_rec_queue during read and write
  * operation. */
 protected semaphore perf_rec_queue_sema;


 // ****************************************************************************
 // Protected Data Properties
 // ****************************************************************************
 /** 
   * Triggered when a reset is received 
   * If a reset in received, this event is triggered prior
   * to the is_sampled event to ensure that all threads are terminated 
   */
  protected event reset_received;
  
  /** Triggered when a new transaction is started */
  protected event new_transaction_started;
  
  /** Triggered when a new READ transaction is started */
  protected event new_read_transaction_started;
 
  /** Triggered when a new transaction is started */
  protected event new_write_transaction_started;
  
  /** Triggered when a READ element is deleted from active xact queue */
  protected event active_read_xact_queue_empty;
  /** Triggered when a WRITE element is deleted from active xact queue */
  protected event active_write_xact_queue_empty;

  /** port configuration */
  protected svt_axi_port_configuration cfg;

  /** clock period */ 
  protected real clock_period = -1;

  /** current cycle */
  protected longint curr_cycle = 0;

  /** current time */
  protected real curr_time;

  /** Async reset assertion time*/
   protected real reset_async_time;

  /** Stores the last sample time. Used for calculating clock period */
  protected real last_sample_time = -1;

  /** The cycle in which last arvalid was driven high*/
  protected int last_arvalid_cycle = 0;

  /** The cycle in which last arready was sampled high*/
  protected int last_arready_cycle = 0;

  /** The cycle in which last awvalid was driven high*/
  protected int last_awvalid_cycle = 0;

  /** The cycle in which last awready was sampled high*/
  protected int last_awready_cycle = 0;

  /** The cycle in which last wvalid was driven high*/
  protected int last_wvalid_cycle = 0;

  /** The cycle in which last wready was sampled high*/
  protected int last_wready_cycle = 0;

  /** The cycle in which last wlast, wvalid, wready was sampled high*/
  protected int last_wlast_wvalid_wready_cycle = 0;

  /** The cycle in which last rlast, rvalid, rready was sampled high*/
  protected int last_rlast_rvalid_rready_cycle = 0;

  /** The cycle in which last rvalid was sampled high*/
  protected int last_rvalid_cycle = 0;

  /** The cycle in which last rready was sampled high*/
  protected int last_rready_cycle = 0;

  /** The cycle in which last bvalid was sampled high*/
  protected int last_bvalid_cycle = 0;

  /** The cycle in which last bready was driven high*/
  protected int last_bready_cycle = 0;

  /** The cycle in which last acvalid was sampled high*/
  protected int last_acvalid_cycle = 0;

  /** The cycle in which last acready was driven high*/
  protected int last_acready_cycle = 0;

  /** The cycle in which last crvalid was sampled high*/
  protected int last_crvalid_cycle = 0;

  /** The cycle in which last crready was driven high*/
  protected int last_crready_cycle = 0;

  /** The cycle in which last cdvalid was sampled high*/
  protected int last_cdvalid_cycle = 0;

  /** The cycle in which last cdready was driven high*/
  protected int last_cdready_cycle = 0;

  /** The cycle in which last tvalid was sampled high*/
  protected int last_tvalid_cycle = 0;

  /** The cycle in which last tready was driven high*/
  protected int last_tready_cycle = 0;

  /** The cycle in which last arvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_arvalid_cycle = 0;

  /** The cycle in which last arready was sampled high - update is deferred by a clock*/
  protected int deferred_last_arready_cycle = 0;

  /** The cycle in which last awvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_awvalid_cycle = 0;

  /** The cycle in which last awready was sampled high - update is deferred by a clock*/
  protected int deferred_last_awready_cycle = 0;

  /** The cycle in which last wvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_wvalid_cycle = 0;

  /** The cycle in which last wready was sampled high - update is deferred by a clock*/
  protected int deferred_last_wready_cycle = 0;

  /** The cycle in which last wlast, wvalid, and wready was sampled high - update is deferred by a clock*/
  protected int deferred_last_wlast_wvalid_wready_cycle = 0;

  /** The cycle in which last rlast, rvalid, and rready was sampled high - update is deferred by a clock*/
  protected int deferred_last_rlast_rvalid_rready_cycle = 0;

  /** The cycle in which last rvalid was sampled high - update is deferred by a clock*/ 
  protected int deferred_last_rvalid_cycle = 0;

  /** The cycle in which last rready was sampled high - update is deferred by a clock*/
  protected int deferred_last_rready_cycle = 0;

  /** The cycle in which last bvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_bvalid_cycle = 0;

  /** The cycle in which last bready was driven high - update is deferred by a clock*/
  protected int deferred_last_bready_cycle = 0;

  /** The cycle in which last acvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_acvalid_cycle = 0;

  /** The cycle in which last acready was driven high - update is deferred by a clock*/
  protected int deferred_last_acready_cycle = 0;

  /** The cycle in which last crvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_crvalid_cycle = 0;

  /** The cycle in which last crready was driven high - update is deferred by a clock*/
  protected int deferred_last_crready_cycle = 0;

  /** The cycle in which last cdvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_cdvalid_cycle = 0;

  /** The cycle in which last cdready was driven high - update is deferred by a clock*/
  protected int deferred_last_cdready_cycle = 0;

  /** The cycle in which last tvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_tvalid_cycle = 0;

  /** The cycle in which last tready was sampled high - update is deferred by a clock*/
  protected int deferred_last_tready_cycle = 0;

  /**
    * The configuration that will be used for the current time interval
    */
  svt_axi_port_configuration curr_perf_config;

  /**
    * New configuration submitted by user which may have updated performance
    * constraints and which need to be used at the next time interval
    */
  svt_axi_port_configuration new_perf_config;
  
  /** Timer used for performance intervals */
  svt_timer perf_interval_timer;

  /** Timer to track periods of inactivity for READ on the interface */
  svt_timer perf_read_inactivity_timer;

  /** Timer to track periods of inactivity for WRITE on the interface */
  svt_timer perf_write_inactivity_timer;

  svt_amba_perf_rec_base  perf_rec_queue[$];

  bit stop_perf_timers = 0;

  svt_amba_perf_calc_base perf_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_write_throughput_calc;

  svt_amba_perf_calc_base perf_min_write_throughput_calc;

  svt_amba_perf_calc_base perf_max_read_throughput_calc;

  svt_amba_perf_calc_base perf_min_read_throughput_calc;

  svt_amba_perf_calc_base perf_max_write_bandwidth_calc;

  svt_amba_perf_calc_base perf_min_write_bandwidth_calc;

  svt_amba_perf_calc_base perf_max_read_bandwidth_calc;

  svt_amba_perf_calc_base perf_min_read_bandwidth_calc;

  //vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
IoTEGdolf5XQZmvTJTjm9SGr/23gNoB955cMuqnJdeU8Pv+9CtKkCO+wRbN/Ac77
KvxVCSP9t9qfCPBNFKpIPpeYAkDtc88p/BsFai8NhQqmNCkgX/+kNB08Dn5zf7zE
NtlGRjlm/5C5itXIzPlqELEUUjj7WMzDJGxPgGgh24Y=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 335       )
dze2qE0R7M4yw9RaK+fGwpP3T6gSlvNno86cXvgQPyvySy07ZlXaa9QrdoikjEMf
feYcyfiVnaSjCpv9yV+b7cMvObTvw/s3r9serVSytCUXhBh8vosHE39O1t9KKvIr
4L5Kql+Q4/9Clz8dLVOEPB0NZzryGiQ3MOVwfekS0mIboLzhtv7wYujyfMOJBAa4
xtRVOChbCWOGRKHLRtoboFuXf2nW97m3IybyY7giKZ3AybhKRYsjeIrcSXR2EyO/
v1bKAW8qiKTfSjcY4y0v60MJ0Q2cbU1C/tb0yXY/UTcxiaTXtLUW4NdxeQvcTyt6
0zz/wwzxZltopmaPjrnyYWbE2d6BawegcnL9RSKgwtlLoLFOS+AaCZxxPdIDnMRZ
d4+LAyUMYFKSnNPaV4dIXDrL+PzbEvF3LKC5IbT6l99M7vhTbymyFjNAvAAGdhFO
`pragma protect end_protected

 /** @cond PRIVATE */
 // ****************************************************************************
 // Local Data Properties
 // ****************************************************************************
 int report_new_clock_period = -1;
 /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /** Variable that keeps count of number of DVM Syncs which are accepted and DVMCOMPLETEs
    * are yet to be added to the queue */
  int num_active_dvm_sync_xacts = 0;

    /**
    * Method that auto generates DVM complete transactions
    *
    * @ param snoop_xact Handle to the DVM SYNC transaction for which DVM complete must be generated
    * @ param phase UVM phase from which this task is called
    */
`ifdef SVT_VMM_TECHNOLOGY
  extern virtual task send_auto_gen_dvm_complete(svt_axi_master_snoop_transaction snoop_xact);
`else
  extern virtual task send_auto_gen_dvm_complete(svt_axi_master_snoop_transaction snoop_xact, svt_phase phase);
`endif

  /** Returns if all Snoop DVM COMPLETEs are received for coherent DVM Sync sent */
  extern virtual function bit is_dvm_snoop_sync_complete_done();

  /** Wait for conditions for DVM */
  extern virtual task check_and_wait_for_dvm_complete_conditions(svt_axi_transaction xact);



  /** @endcond */

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter UVM report object used for messaging
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter OVM report object used for messaging
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_xactor xactor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Detects reset async */
   extern virtual task sample_reset_async();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Initializes master I/F output signals to 0 at 0 simulation time */
  extern virtual task async_init_signals();
  
  extern virtual task suspend_signal(string signal_name = "");
  
  extern virtual task resume_signal(string signal_name = "");

  /** Initializes master I/F output signals to 0 at 0 simulation time */
  extern virtual task default_signal_values_async_reset();
  
  /** Initializes master I/F output signals to 0 after waiting for a clock cycle delay */
  extern virtual task initialize_during_dynamic_reset();

  /** Initializes signals */
  extern virtual task initialize_signals();

  /**Aborts the transactions and writes to analysis port if reset is in progress. */
  extern virtual task process_reset_for_new_transaction(svt_axi_transaction xact);

  /** Sets the configuration */
  extern virtual function void set_cfg(svt_axi_port_configuration cfg);

  /** Waits for a any transaction to end. */
  extern virtual task wait_for_any_transaction_ended();

   /** Sets the clock period */
  extern function void set_clock_period();

   /** Returns clock period value*/
  extern virtual function real get_clock_period();

   /** Returns current clock cycle value*/
  extern virtual function longint get_current_clock_cycle();

   /** Returns current time measured as (current clock cycle * clock period) */
  extern virtual function real get_current_time();

  /** Creates timers used in the model */
  extern virtual function void create_timers();

  /**
   * Sets the delays in the transaction based on observed values.
   * Calls to this function must be made before "set_deferred_event_cycles" 
   * (which updates the "deferred_last_*" variables) is called to reflect the
   * corresponding values in "last_*" in variables of this cycle. 
   * In the case of bvalid_delay, bvalid can be sent before the address
   * is received or after the address is received. In either case, the 
   * burst_length information is required to calculate the bvalid_delay.
   * If bvalid is sent before the address, the call to this function to
   * update bvalid_delay must happen only when the address is received 
   * If bvalid is sent after the address, the call can be
   * made when bvalid is sampled (as in the case of other signals)
   */
  extern function void set_observed_transaction_delay(svt_axi_transaction xact, string delay_type);

  /**
    * Sets the "deferred_" variables to the values passed through this function.
    * The set_observed_transaction_delay function works based on the "deferred_"
    * values of event cycles. This function needs to be called after the 
    * set_observed_transaction_delay function is called, so that the current
    * cycle information is propogated to the corresponding "deferred_*" variables.
    */ 
  extern function void set_deferred_event_cycles();

  /** Checks if the handle given matches any of those of the active transactions. */
  extern virtual function void check_xact_handle(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

   /** Checks coherent transaction. If data is available in cache it is retreived */ 
  extern virtual task process_coherent_transaction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Reserves an index in cache for allocation of this transaction */ 
  extern virtual task reserve_cache_allocation(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output `SVT_AXI_MASTER_TRANSACTION_TYPE lru_xact);

  /** Does the necessary processing to end a transaction */
  extern virtual task end_transaction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit is_removed=0);

  /** 
    * Updates the cache based on snoop response assigned by user after 
    * receiving a snoop transaction from the input channel 
    */
  extern virtual task post_snoop_cache_update(svt_axi_master_snoop_transaction snoop_xact);

  /** Waits for post_snoop_cache_update() method to complete if any activity
    * is observed on the SNOOP channel */
  extern virtual task is_post_snoop_cache_update_done(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit check_outstanding_queue= 0);

  /** Adds a new snoop transaction to the queue */
  extern virtual task add_to_master_snoop_active(svt_axi_master_snoop_transaction xact);

  /** Adds a new snoop transaction to the queue */
  extern virtual task add_to_ic_snoop_active(svt_axi_ic_snoop_transaction xact);

  /** Drives the awakeup signal during idle time period of addr channel */
  extern virtual task toggle_awakeup_signals_during_idle_channel( );
  
  /** Drives the acwakeup signal during idle time period of addr channel */
  extern virtual task toggle_acwakeup_signals_during_idle_snoop_channel( );
  /** 
    * Adds the transaction to the internal queue. 
    * Blocks when the  number of outstanding transactions is
    * the configured max. value.
    */
  extern virtual task add_to_master_active(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Notifies the slave that a new transaction is received from input port.
    */
  extern virtual task notify_slave_new_xact_received_from_input_port(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** 
    * Waits for a new snoop transaction. The monitor uses this task to get a 
    * handle to the new snoop transaction.
    */ 
  extern virtual task wait_for_acvalid(output svt_axi_master_snoop_transaction xact);

  /*
   * Returns the number of outstanding transactions
   */
  extern virtual function int get_number_of_outstanding_master_transactions(bit silent = 1, output `SVT_AXI_MASTER_TRANSACTION_TYPE actvQ[$]);

  /** Returns the number of outstanding transactions. */
  extern virtual function int get_number_of_outstanding_slave_transactions(bit silent = 1, output `SVT_AXI_SLAVE_TRANSACTION_TYPE actvQ[$]);

  /** Returns the number of auto-generated transactions. */
  extern virtual function int get_number_auto_generated_xacts();

  /** Returns the number of dropped coherent transactions. */
  extern virtual function int get_number_dropped_coherent_xacts();

  /** Advances clock by #num_clocks */
  extern virtual task advance_clock(int num_clocks);

  /** Steps one clock*/
  extern virtual task step_monitor_clock();

  /** Waits until a valid or handshake takes place on any channel*/
  extern virtual task wait_for_bus_activity();

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_arvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_awvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_first_data_before_addr_wvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_tvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Drive the idle values after initial reset */
  extern virtual task drive_idle_val_initial_reset();

  /** 
    * Adds the transaction to the active queue. 
    * Blocks when the  number of outstanding transactions is
    * the configured max. value.
    */
  extern virtual task load_active_from_master_buffer ();

  /** 
    * Adds the transaction to read_xact_buffer or write_xact_buffer 
    * depending on whether its a read or write transaction. 
    */
  extern virtual task add_to_master_buffer(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);
  /** Detects initial reset */
  extern virtual function void detect_initial_reset();

  // -----------------------------------------------------------------------------
  //                                EXCLUSIVE PROCESSING BEGIN
  // -----------------------------------------------------------------------------
  /** It returns 1 if there are pending exclusive read transactions in
   * exclusive_read_queue for which matching exclusive write has not come
   * */
  extern virtual function bit pending_exclusive_access_transactions();

  /** It checks the transaction with the same ID stored in the queue */
  extern virtual function void check_exclusive_sameid(svt_axi_transaction xact);

    /** Pushes the transaction into exclusive read queue after all the data beats
    * of exclusive read transaction is received
    */
  extern virtual function void push_exclusive_read_transactions(svt_axi_transaction xact, string kind="");
 
 /**  Removes  the transaction from exclusive read queue if any of the data beats recieves a erroneous response
    * of exclusive read transaction is received
    */
  extern virtual function void remove_exclusive_read_transactions(svt_axi_transaction xact);

  /** function that compares the expected and configured RRESP for exclusive
   * read transactions */
  extern virtual function void perform_exclusive_read_resp_checks(svt_axi_transaction excl_resp_xact);

  /** It returns 1 if transaction with AWID = ARID exist in the exclusive_read_queue queue */
  extern virtual function bit get_exclusive_read_index(input logic [`SVT_AXI_MAX_ID_WIDTH - 1 : 0] awid, 
                                                       logic [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,
                                                       output int ex_rd_idx);
  

  /** It monitors memory location for exclusive access */
  extern virtual function void check_exclusive_memory(svt_axi_transaction current_xact);
  
  /** It monitors the response for exclusive write transaction */
  //extern virtual function void process_exclusive_write_response(svt_axi_transaction excl_resp_xact, input bit excl_write_error);
  extern virtual function void process_exclusive_write_response(svt_axi_transaction excl_resp_xact, input bit excl_write_error, string kind="");
  // -----------------------------------------------------------------------------


  extern virtual task wait_for_cache_update_post_curr_snoop(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit is_snoop_to_same_cache_line);

  extern virtual task add_to_master_current_queue(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual function bit add_xact_with_same_id_to_queue(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,output bit[`SVT_AXI_MAX_ID_WIDTH-1:0]  unused_ids_by_active_master_transaction);

  extern virtual task update_current_snoop_xact_handle(svt_axi_master_snoop_transaction snoop_xact);

  /**
    * Creates the transaction inactivity timer
    */
  extern virtual function svt_timer create_xact_inactivity_timer();


  /** Tracks transaction inactivity */
  extern virtual task track_transaction_inactivity_timeout(svt_axi_transaction xact);

  /** Waits until the transaction ends */
  extern virtual task wait_for_transaction_ended(svt_axi_transaction xact);

  /**
    * Tracks suspended snoop xacts and triggers events when they are ready
    * to be added to the queue
    */
  extern virtual task track_suspended_snoop_xacts();

  /** Updates response parameters when supplied through delayed response port */
  extern virtual task update_delayed_response_parameters(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** returns a single unique number from xact ID and ADDRESS */
  extern function bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0] get_uniq_num_from_id_addr(svt_axi_transaction xact);

  /* returns address part of the unique address-id combinatorial number */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH -1 : 0] get_addr_from_num(bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0] num);

  /* returns id part of the unique address-id combinatorial number */
  extern function bit[`SVT_AXI_MAX_ID_WIDTH-1 : 0] get_id_from_num(bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0] num);

  //-------------------------------------------------------------------
  //                       PERFORMANCE ANALYSIS
  //------------------------------------------------------------------
  /** Main task that tracks performance parameters */
  extern task track_performance_parameters();

  /** updates the READ inactivity time performance parameters */
  extern task track_inactivity_time_for_reads(int perf_rec_index);

  /** updates the WRITE inactivity time performance parameters */
  extern task  track_inactivity_time_for_writes(int perf_rec_index);
  
  /** Updates performance parameters when a transaction ends */
  extern function void update_xact_performance_parameters(svt_axi_transaction xact);

  /** Updates performance configuration parameters based on a new configuration*/
  extern function void update_performance_config_parameters();

  /** Collects performance statistics when an interval ends */
  extern function void collect_perf_stats();

  /** Creates all the performance classes used for calculation of each metric */
  extern function void create_perf_calc_base(svt_axi_port_configuration cfg);

  /** Gets the performance report as a string */
  extern function string get_performance_report();

  /**
   * When invoked, indicates if the performance monitoring is in progress or not.
   * - This is applicable only when the svt_axi_port_configuration::perf_recording_interval is set to -1.
   * - Returns 1 if performance monitoring is in progress when this method is invoked
   * - Returns 0 if performance monitoring is not in progress when this method is invoked
   * .
   */
  extern function bit is_performance_monitoring_in_progress();

  /** Reports end-of-simulation summary report, checks etc */
  extern virtual function void report();

  /** format report string */
  extern function string format_report_str(string exp_str, real exp_val, string act_str, real act_val, string unit_str);

  /** Gets summary report based on values in perf_rec */
  extern function string get_summary_report(svt_amba_perf_rec_base perf_rec);

  /** Stops all performance monitoring and kills the thread that is tracking performance */
  extern function void stop_performance_monitoring();

  /**
   * When invoked, performance monitoring will be stopped if already the monitoring is in progress.
   * - This is applicable only when the svt_axi_port_configuration::perf_recording_interval is set to -1.
   * - Returns 1 if performance monitoring is stopped as a result of this method invocation
   * - Returns 0 if performance monitoring is not stopped as a result of this method invocation
   * - If the performance monitoring is in progress, that is is_performance_monitoring_in_progress() returns 1,
   *   but the axi_port_perf_stop_performance_monitoring() is not invoked, the port monitor invokes stop_performance_monitoring
   *   method during extract phase.
   * .
   */
  extern function bit axi_port_perf_stop_performance_monitoring();

`ifdef SVT_AMBA_ENABLE_C_BASED_MEM
  /** Converts an AXI transaction to memory transaction */
  extern function bit convert_axi_to_mem_transaction(svt_axi_transaction xact, int mem_data_width, bit convert_read_data, output svt_mem_transaction mem_xact[$]);

  /** Populates data in memory transaction into the given AXI transaction */
  extern function bit populate_mem_data_to_axi_xact(svt_mem_transaction mem_xact[$], int mem_data_width, svt_axi_transaction xact);
`endif  

  /** Enables/disables performance monitoring of each metric based on configuration*/
  extern function void check_performance_monitors(svt_axi_port_configuration cfg);

  /** Enables/disables of all performance monitors based on the argument */
  extern function void set_performance_monitoring(bit enable_monitoring = 1);

`ifdef SVT_UVM_TECHNOLOGY
  extern task write_to_tlm_generic_payload_analysis_port(svt_axi_transaction xact);
`endif

  `ifdef SVT_AXI_QVN_ENABLE
  extern virtual task qvn_process_token_request();
  `endif

  /** Tracks the timeout for the signal argument provided with its timeout value given
    * w.r.t to the event or status provided in the argument list. 
    * Mode will be changed to enum type as seperate activity. 
    */
  extern task track_timeout(svt_axi_transaction xact, 
                            longint timeout_val,
                            string timer_name, 
                            int mode, 
                            bit status_equal,
                            svt_axi_transaction::status_enum sts_val,
                            event timeout_event,
                            string port_mon_name=""
                           );

  /** Tracks the snoop channel timeout for the signal argument provided with its timeout value given
    * w.r.t to the event or status provided in the argument list 
    * Mode will be changed to enum type as seperate activity. 
    */
  extern task track_snoop_timeout(svt_axi_snoop_transaction xact, 
                            longint timeout_val,
                            string timer_name, 
                            int mode, 
                            bit status_equal,
                            svt_axi_transaction::status_enum sts_val,
                            event timeout_event,
                            string port_mon_name=""
                           );			   

  /** pushes an exernal coherent transaction into port monitor */
  extern virtual task push_external_coherent_xact(svt_axi_transaction xact);
  /** pushes an exernal snoop transaction into port monitor */
  extern virtual task push_external_snoop_xact(svt_axi_snoop_transaction xact);

  /** 
  * Returns the number of READ transcations that have started  and in 
  * active queue
  */
  extern virtual function int get_num_started_read_xacts();
  /** 
  * Returns the number of WRITE transcations that have started  and in 
  * active queue
  */
  extern virtual function int get_num_started_write_xacts();

  /**
    * This method is used to get list of all IDs which are currently under use by outstanding transactions. However, user
    * can choose the type of outstanding transactions this method should consider while extracting ID of active transactions.
    * "mode" and "rw_type" arguments should be used for this purpose.
    *
    * It returns '1' if total number of unique IDs currently used by active transactions, is less than all possible ID that can
    * be used by an AXI transaction. This helps in determining whether randomizing ID field of a new transaction which should
    * not be part of the all the IDs currently in use, is possible or not.
    * 
    * @param mode Type of outstanding transactions this method should consider while extracting ID of active transactions.
    *             Currently it supports following modes (defined as string) ::
    *               - "non_dvm_non_barrier" => all transactions which are neither DVM nor Barrier  (default)
    *               - "non_dvm"             => all transactions which are not DVM 
    *               - "non_barrier"         => all transactions which are not Barrier 
    *               - "dvm"                 => all transactions which are of DVM type 
    *               - "barrier"             => all transactions which are of Barrier type
    *               - "dvm_barrier"         => all transactions which are either DVM or Barrier type
    *               - Note: if "rw_type" is set to '0' then only read channel transactions will be considered for non-dvm
    *                       and non-barrier type
    *               .
    * 
    * @param rw_type Indicates which channel id width should be considered.
    *               - ' 0 ' => only read channel id width and transactions should be used
    *               - ' 1 ' => only write channel id width and transactions should be used
    *               - '-1 ' => common or either of read or write channel id width and transactions are used
    *               .
    * 
    * @param use_min_width If set to '1', minimum of read and write channel id width should be used otherwise maximum.
    *               This is applicable only if "rw_type == -1" i.e. no particular channel id width is specified.
    * 
    * @param silent Suppresses debug messages from this method if set to '1'
    */
  extern virtual function bit get_ids_used_by_active_master_transactions(output bit[`SVT_AXI_MAX_ID_WIDTH-1:0] id_list[$], input string mode="non_dvm_non_barrier", input int rw_type=-1, input bit use_min_width=1, input bit silent=1);

 /**
   * Method that randomizes DVM complete transaction
   *
   * @return A handle to the randomized DVM complete transaction 
   */
  extern virtual function `SVT_AXI_MASTER_TRANSACTION_TYPE randomize_dvm_complete_xact();
  extern virtual function bit is_in_reset();
  extern virtual task         wait_for_sampled();

  /** Checks if a WU/WLU transaction is received from the sequencer while
    * there is activity on the snoop channel. This is checked only when
    * snoop_response_data_transfer_mode is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC
    * Needs to be done so that the WL/WLU does not get ahead of an
    * auto-generated WRITEBACK/WRITECLEAN
    */
  extern virtual function bit is_wu_wlu_during_snoop_addr_activity(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /**
    * Waits for WRITEBACK/WRITECLEAN generated for snoops to be added
    * to queue. Applicable only when snoop_response_data_transfer_mode
    * is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC
    */
  extern virtual task wait_for_pending_wb_wc_for_snoop();

  /** Gets the time at which an address was invalidated due to a MAKEINVALID coherent transaction */
  extern virtual function real get_makeinvalid_invalidate_time(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
  /** waits for transaction which has been blocked by other transactions more than `SVT_AXI_NUM_BLOCKED_XACTS_ALLOWED number of times.
    * It wait for those blocked transaction to finish. This will avoid starvation of some type of transactions and will provide
    * more fair chance to all the transactions to proceed
    */
  extern virtual task wait_for_severly_blocked_transactions_to_make_progress(`SVT_AXI_MASTER_TRANSACTION_TYPE xact=null);

  /** waits until VIP is out of reset */
  extern virtual task wait_for_out_of_reset(int mode = 0);

  /** waits until VIP is in reset */
  extern virtual task wait_for_reset(int mode = 0);

  /** Wait for start event for performance monitoring */
  extern task wait_for_performance_monitoring_start_event();

  /** Wait for stop event for performance monitoring */
  extern task wait_for_performance_monitoring_stop_event();

 /** Perform master signal valid checks during reset*/
  extern virtual function void perform_master_signal_valid_checks_during_reset (
                                                                          logic  observed_awvalid,
                                                                          logic  observed_arvalid,
                                                                          logic  observed_wvalid);

/** Perform slave signal valid checks during reset*/
  extern virtual function void perform_slave_signal_valid_checks_during_reset (
                                                                          logic  observed_rvalid,
                                                                          logic  observed_bvalid);

endclass
  /** @endcond */

//----------------------------------------------------------------------------

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Q+PJda096deXstvFu8b6cqctzpmXIVvB+a4oS1nLMkpZIO46pTRj6/Ik7f4WGOGZ
vx9itDnteIAjcc2As6ZFZBw4vD2Vwy578msU+P3np5OrWYD9c0IPLCdlNAajHXnl
6Tvq2Kv6RGuY+kkU1cBdky0G1UlpyLfOTyVLPqW/ou4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4101      )
QR1yCL1OreZcnfPUkxWzW0iaHKYacMnaTuzJ9uDDBN63r/82U+k5nR4ZR0YqT6Tq
M0ElFB+Chj/y1DdMGfDF/iZxVTcAKnb27yQkO6TKztqVO8Fyh/C7PLevhUTd/6mR
T/fJBVkjAU3agsLKrw60edbJQ7kQPJu8R4Pd+9DvQrw7RJIU80nPUfJsUH5jB/Rk
aC9WETwFcgKwsClm6GE8d5X8nR43iUZjREFIuM/Fp4To4i2e7g3UGODwslGWRi2E
uWgYBxB2pVu8KU7UUZiGnwypI1mDNpMe0HmUbbU5ob+ynAivh523hZcU7pvscEbq
XJNb7inTlhkmudlIbvDEpAiT40EzLZMmj+b5eDpPh1ucCyr2k8QRVr363ocmG4/b
uKEfnMko7bmEXVw/eWeorQFmb8MKYXIGe1lB1+9h1ON5GIsjUCkaqgFrjSFAlk39
yCM6gT4TiBD/BQBQwb7IMIJf/eaWNJLjFbrx+Rp5jBya7gq5WIYWnNBpY6K4cpvc
PxFH/wPm15y6zaUA1L3uhvjfwtgtpy4sCLzTMo1N/SOrIfV4Eo7l/8ABhfkwc/p+
BUTZSrS96nQDPxmGpu2MbfYilZuX3Nf+L9MeqjoqdG68sMTmKokKPVr5umjdCl4r
Q+5ANSHq1cd4bhJ2mGP4r1F70yx0pmLguFavMlv6X+ixTBOfkFwBUU1myEvVT7hM
LhKh7PmhmOYOYk8wJyMPK5xMwPdSxoKn25fXiaGqpbElGHChxnzhlNPKR32C+CXS
Mc86TqIBs/RHc1cRyXUyySjGKKliXgGlvge98AHflo1L41Py0uQli7VzkwDa4xUc
kpOwxrgu8WgbnL5Oqv3sAlB6rVuK87ELM18TtEiVPI58TI+f2ObJ1roL/h5pMdHN
wrccW07UK3IHE2f3ZV+w4DiA+Xx0mUs3xoxFJY1jnUr21vhmauI9Y+c5M/+1i2c+
63fz1KWsDpu2XpMkOprJW00YS4G7gPAICImNNAa+HSIYkxkbe3xgHXYt1F75UMpQ
7aVMJoUst32/Hz75pQfNHHXHkbe6OeY7xoNHiT2y3t5xs5PfVhpcKH5ry+0rosd+
COaAjXjlh6lYQLWA8fS7y9sK9rtbgFJPE3tIhKFX8TJQwY9MbcPAYt8S9CqyrRtU
xJqjb20d8VD7YKXf/DyBTahbe2ZWPBL66AK9tODCCioS3Xyt0XNco5575YEKvrhj
LYj2C17oofxdf2oRGatPrFRct1jJSlJjsDqOYbtFtQdeyXWVAs+fKH4eVlbPSIMD
IvX84muNMn9onZnVMmyPaXK0E+T6OIbBAtbnYR7uaAmaup7JYE6QMVgjoOaptJFf
HR3JpDd0YFAGN6IHv0GsFx8Oz1FtOjsxTcrHjMLTamSQePe0qhd4eLdxHm5or9WL
OqbAurrbx4Nxr/e7CacUL3yBlsToXiT0hOIuWbm/Yr19rUja/Z0UMk29GKyXLaj4
yu7UPbU/fZOqcIj1pH4xNQwt2/8kT0K0YQvhBtaIuXNqD6BBFPNN9T4j4G99yVUp
0Gcj6nF1m0b5bEjq6vEmv/droeMx4WI2fjuPa9vIfk57jqyM1JLuNtApOm407qcS
G80deaG/ozX5fMDE/y1hddLNfhigO+GoocAE7fNqizIuIVV8tf9N29Bflcsdzjdq
s9BcfsdIQDhO2V76Nm0mj2NbZ/yN3uO5+U1xJc4bW3BKNe7xYbJoX5oL4DdbVNM+
C/nsHWbCksLSbdin7DfYTxoJDaOvjMxsYRtgP7q9eYYhaGTPcoH9X69ez/Ur9QL0
62JcD4S5+Xk3qZhv07g4w1hGkwiHDWNaSWFp1D2t6244Qu68mCv9cN7SzrT0bmU5
ezubBUIP1emyElhq+ktcKI7ZKoz/hEWJyqGtFmHRjTSlwFA9ZUS2B3CyFvJTUT10
hnoA7RZgJKc3My5ymgWe5CcbbKhz6iu8XG+2NYwJ13hAz1itf6n8boV+JR6GzXHl
rjy2aLK0DeNCvR/hUC7BCeIp58xEgt/tav+kU5lF+4rFOzOiUJ5ewIkW9V8GhpDK
Uz4HLacpz4DAIV9rETyIxrLlehWj997kv24h8Zc4iSItVLLu9slUI2elynrIH8U8
jKbMWpOnCZ9KtgpTlNhwQalsurL2mZyBKgi/S6zKvtGKQtvbj2q1Jdf5jZ4zIKod
m8G3QXuCFcivC3Hz1p7DvOrhFXWysImjBn74qvW+rb0D9pFkgrKZ1IHKJiKj3rW4
M9Eoi5qMyBvMOwL7yENEcRXYoEsWgtHVv/a7uXMWuAPWGfOnoxCBTJSEUAxqnzhA
ZAcXqi/aBpPQl5/obgmluyQWIghZDkkb/ZhypJHZjVD0opGmQyYtpKY5ktMlmN4m
I4M+FIt4HHGL23nlBOtzqHmct0QTgsfpyzNnkAIcHx9owu9J4aM1zMYhcSSF2hki
Ib/k0JNNdKhXa0H96SAKKiBNOnJwWmCMOxcnHDgDNSYQI7/e3akMKMGlTVKEjBRZ
ZHu/oH+cUqTp1UB2+1wihbWP0qfQR50EekdBUsPyZGdqXP11OAnrFFgnlB1nuiCb
CABrUZwdBjUgiK6bhPiqkWz7ir7X0zQo8Qq3vhL6TVIvDe0VvOFoJ8BWclOYE4Lh
tHtNZ4Mnj5pci/TwUcSbtZHeDAXRm+rv97IKWlVO/5nYFnr7XYXxNyiMfOePmxIT
y84/ushqCHUbJ8HcBuhPlbwhcdyHa0wdD0CwnvK6DCVtbRaFbXMWBuWqX9DE3CIh
lnVCCpETDbmjVu4QRJ8cpJiSucO/Ik1rXMKuhRz/p+T2E8xgk80kHgWbG216hDEQ
zudMW94zGgfOQ/YFzW424Wtl/EUuCo0fX72DYiAeATIvt1fkUoYVDQiYyuGBjO0Z
rZUNV56xWRQ85W4S8B8803rbneurIlKd1YL4a+T0CkbBJ9vjt3rs/BmY/33fcD1e
pCvOyRXtje1IqmVgYulSVUJfoVAb/TMamUjdetS7q89iGRRCF5kRbpRuPTs2Ugo1
mp0UcpNgXxkf4VnAvZEQu1nJBgkq1FDWtohg4SWbxZ6PRSSFQNMus+/54BEGh9uX
yD2786gt64OPzrXWrIa7E0Dh12AeP7DOxz9c3bXQTj1aDZY6OWU27DUEBBGx0Gun
brf9YcpMjRacfFDS34GjQOo/fe1Ud0q/q4DxiQtKwoAFKcy1dJHxF9BlgF+2gCJ1
HzJfAapabNC1539hGrkCKjHtZ6m/ZqzkKcjCy64gtQfZAmnBE9oV6L6FXzYFoWaw
wG0/iysraDxPg7JokTjvweB3CpxG/CV2gjr26oe1PyhYUtcybMsNa1GHaKX+hjSG
NnNEgysCs7zQrUTOK+HzTIIXannWDNxDXguLF11rjQ6FhHwpl0GbdkDyB88ojGTh
vSkkMk7C0w4tecgbaMBsB/y8QxF5Nj7xSu7BqxQr+XFlRrfxTDJqoZoCaSefewpP
BeukYjLtKhqbcjnHPEhBrlDJvkP+fBdQunvmLDfbH+0kNZNb/RTLt66wyH4CwnJO
XRLlMzHX5+mxiIRoRM3SZlpXPadkVCNk+HNy3qWBRqV+WDBX51uh2AmilqOvXcDH
Akg3wverlFCrA7fJ7RGi61Z+QioRreWMYx1pyw6BooRy19oFvetHbZHe2yW9Lew2
0Sa2f2X+ix+QjWJzO/Sx/4NZ3xrLOTInGRpROKMKzoNyRaVRfpfeSDjWq7K75TwT
WJfw7PvOQdDSX2KBa/EIz+LIpMJkSx+EZue5Op0AWhd0ZEX2bHvz7DgY80O/0KN/
QhR7DyhDG377JhiTM2b8s+0QoSupVBO+kQ9lzXy3XEgakCLSrlHRA8CzfrcG2S3Y
MqFl4MQ+nGPaiOOSSd7dVDAkTJnibhE78pqK3gyYIQ3hIS9+7xxfGh6UoCapsGik
B2fFy3NMy8GpinMrkx5k9PAX1q6nd1aFoSJRsGbFrL0govUVO4cv0FAw29TfyQbE
ziZbh3B6oP0wyI+1S0CivVQ60Kx0epVZvXN54YHKFsR11wjBcI+Pl2Mb1sChCNh1
JXKpPPieeqW5aO3B9PLgh9Dh5/Ii76KhcuUf+hyTAkuGEnuAy5kJnqUTLQYL7OnH
7XM5F0IzuLWA1/KAh0Mwp+v8Vm6j045c6BFEa/+Gc4DbOpBRzSA6gIG14P48/LE2
MrLFnWPOYiAakZZT4vVaC4GdTcRGKep9ZQqvLc2NhW2XpU5RWYZ0W3uYjAPk9KGO
f+0TROKIvTFlrHBa9XM+aLky2DVDr66JsUkaBSmzZHOkgKjoz9w0oUZneAS0MUQp
MSZcIjL2+43ZCnpgol9nyiFKQZ5T54PjmEovL7hprgLDeN0VBZz+wmyJesKXlDWD
Tvf8XSWdaZwY814CA7lm/AWqf10hHp8R59oFcTGkviB3N/N+v43jWxZ28UG1DTHM
S+QvFuoQ1FMJBZzEbXRgQChAn9MhzmJhBfGrvnprTpMO1xstxqpoSfuvY0YSuo8U
VlN0VEh1q6mL5iTL95ZjsbbfANV3AYjQLMAmdUXVzN8TTOgvSqMA+N8lXdYo3FIv
vDrMxsNPhjkQstnarZ+7YF56V/3y98l1Bu+gZhrde0xbspUv7hCWUxgn3p+VUCkJ
zIS39Ciq94L+vIDVrKxs1hafABcJ0VcK7UhFMPdoYD3PpENIa45k7QNm12jzA/vM
kP3r5t5meZ0Gxl9xL1dmKICjGvikEswpFobx7Yqb8VLkbX4G4JW5FcyzRMo2YmH1
EdfDWs2KKRdvmXJukNXgINDr1OSnbNfvUErTGWpK0QkzbXRc3vIW5fduiqNwo6sr
FPfzHCCAn0wnOYGXFZwAE0HZhi0ToTtOPKxjhb0P5OPXpjj8KPEG3shCuaLgqYOu
5hXh3TDhCs472HC+lxyQVWeDZlXbdE09XXIlN/689bGKbCwo7hsL+snZKXoS0P0w
uUiqZ0Avzu5J+f7i78vzozAx/4y+TfUXu0Fl3zbwh7Hz/nc/FpdHx8WdlF38QQQE
/F59v19pgP/IB50AT476YR9wvdwh/GLPOfCCtRuJUEk=
`pragma protect end_protected

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
bTRx1n5KPeXMXnL8bsO6X7Jq6eljGk5nWHYYLD6x+XE6vUVDxSMNOVFMyEJXmfQV
xwKWCBm5gMq9BxNGzT/rtv3FW6459Tmy2EQe1JbFHqKWX1rdY+QVTMaP7NqScn8I
3CknfC9Fr5Rnn4ngtcwD/h6bOiDzfXZkLe4YFPaCczY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 12356     )
tX06OaZscsNNmdconCqw1PPdISppuDC6kfuCnfhUxWYgklCoyaNrQsi6Ekv7KU28
sJ2dAsZVbPxXB+X/Cf0CucHj5D+yvBVIp5k4R//OM82qNPZFm3HUpgWzkUDZJxGZ
xqDgWYyuf5DNEfWwUg70L9odHcIeT0mR5mH6UMkkGNgkI5/v8mTt4N8iEtvQQrSq
xahNbfQTFh5Ba6rCCfjOJ9pEnGHS8OS2toYJdZra9HQLDHqIUsxIjLg76CJBxLfM
gfhOek2eDFRPIcJ0Wp60ZxvDi8CF8MopA1F/Ba2bt3iATOyqjpzDAfkIAFjGDlq0
68qC8hK9cmYRkruAXHupt5ptxfHHgfk9uKAiWsYwSBV9K91URqpVyuhsXKiHN0um
yCnDsXoCmmWE1SHmfC0ENMpGV9yJ6bk/ogj+F2vNpYYMJjLmpNUXbHBS7wqyrIWe
fiIIoKjh1I9KFgGUMrcZFmc6ssKCM1GYSl249omdXzq046gY3eNGu+koSpRfriua
16N2WUl/JMtzot+OzQLMCxtL2dZF9WVD58elfZ2pyvz41507lcO50r21wa/sdwKO
OGKuNnveJ+Ao07VWI5ZOgLJRfspvlWa5eEJhj72DOsMTnf31tRdP9G3Dv7DVz47W
mJJx45v/k+Yzh3T5A3t7RmG74PivAbc2atcLeAtxokHx+GxuorLiP+MhAZ0qYHOE
SoWp1Xv77ZpMXaG7bF/whCGi6nmqcEpUxXAC0B8sIKZEwi1V8nnvXZVXVIlSwaup
e/EoaPs6HAx7p5WESEjk1n8iuR5P92w4+j0/8Bn1BzafqfuEGJYI3L0E0aXPOQKc
bK3y0Gp9Oo98+BbxPUyZa7sRag76EvoJEzrvncdtj8SAqpIt4HhCfqP3eWIzXsV0
+cCxZRaeOjWoi63ako5g1DEAfHkk316BtSf7oxhETH16vA70VCOZ7vd1ulfG92aV
S9r6e7XqF/3M3pDLZ0MoittLKNnqA6GxGR+dUUaF2EC0kJs2p0ZDe62yoFhZeiYV
KHooZfX1ZR3h3fxQsWfAs4r1FM2FxKvMVWAi+s8LMMk5u79/JXSolRla6C1eTxBo
HtFEKTU4cjcpcg9K1KOTO0mhEI2s5DfF5HP8NgN9ZXal86FoB6nJ0F8eSn8RNit2
LQjuHxPb+sEV4BauF+7Te/qv2vH3VCRVgGVNgGtnRGeSRtKYeyBaKnMWvkOUA+oO
3119jcnXM9sP3vdsaSJ5uDHHfkRZegqgtsA0cwTj7zE7JmXvUuBcMNNUyaAkz245
5arschcmUCiSY1HBAFmkSzgPRQ+Vg91icJ5FY4/v7W0CcpKYC79lxKJMALwPGlpz
T9wR1FYOe1J/8mA/IgmR3QfTa3D9HvgmvlhQWywD/X/gRkYEl/HnHSRQpApEjf11
jXOtzDCVvfKp20Q3zJD4BA+UQO+B/wCNAVphiq0hUlP7KnT/KcgcAIYIKO5OlzzP
UK0uIlftF7ThWcov93uDDxzuQGdZHzSZPMnUrkvYhpcc2MVrt80VlTZZxKBv4qaK
5bdAhHV4dy5a1yaed3KmOmA0xqr4GmQ65bMrMUQrX5LLE6gmvE9jw4OGZjX/ULrt
rDSw4DDtaFFdmO20fj8m0AXDQVnZiJIuM9Yg6Bj/1b6CNFRSSq4Gqv9YlK5lsnJn
XLk43QW8AjNqlQVZBbth1Db2YFQJYgFMV+uMyTcIGk6lXYPRgZV3Fu8e8dv+Ium+
gWnztQMTBwV+Wz+Vy10z1fSaba3a3XfPU/RCHT6L2dry+D5DT+afWRS/fzZB7jw3
EXz2TXrmzrK+3QrNl/jzF+zc3dlomWeN3DnVEg2ThzwHhgOsyLieeqWlaFi2a1J1
VeWXLs7ezA4Zs4iGp+UwlL9bM1KnMCQvlgTZ9Mf4P1WH0o7xQwF6IDapeRAx7nQr
1mZZKvcJPy62PTMTc7+FHQvp67oINNZRw5Ug3XfXGXb/pFbxC0sIH/m9KXTmIcPF
6jEx/0C8zm6xxyW1NBYX0hIewTpAk9HPdvfm5CntmKyJ8lyxNX9f9QAKdSoGN/W2
oZrphobF9n7fAvKXZ91lE3wZ+8BqsUl5JNDAxF4ABEzP4MLHcaifEVGxgeyAcBAR
rteatOkZ0Z5eyr0GlZK5SjmngZ+zAKYkIRphVZZ6MiscoStak+wtCHkyYs33fMud
TdC07n2fwacTWh/XdoIQOkrMCnY8p4YHihbB7B9DyIKKO1wQKPTeZhRu2XdaLNaV
L4uYlIxS4L2dxoAuRqJEBk9TVwq4ICj6t9MStztPeEpR4u9axtMBYY3WexeD6w2a
1FV843XsN9B0HrzH73RGRhRHDWWM1wv9gPF7kzZ/06RC75OWSkS6nmSfx2EWy7J2
CZwJYHmG604JGD+gfesVsOB8ErkyIOK1iG8alo/bAvGrUrWhABHcDt/2zhx39Nhd
WSK1eWIG7dxwwDE6WeO6sQ4/1d2bXrAG5vInQ2dr50RQ2ue+VBUoEnP6Bu119GvE
GHonifNUIDqj5vhNgKYiM8W55vdle673OtpG/5TNpBC7XqiIDWZanzTJqpeWmguu
obXGjt1VAk0DSd8SMVt8id6LyxNvow4G2EIgnUjgd52SuieYaE+nbtfSSjdWYqHh
OeFkPTxcUyn+A8S7fRYtfwEM1ESvrywOjjGYFl0NCJAWE5r1oL8Tb8wHssxcb7mg
AxXtdkKVFh67K6WGPiaGmTjg5OOM/ySgwayln/tP3pzF70qVMgAq/Y/75XKhop0h
HGCGcxk3dH1NpWGv350IwKXYze0/zBVxPc6/9w0uEvFYrPoxBePX+4fTiOQq44R9
EWZ7gFwf775CNMcTbF9BoozI7lpAzmWaU8X57plF5P8ZLKrmHjOHR4vAu2hmBzE6
ftA11HeCW95gKbA4rkB1YH5QDCxsFOqlLxjk6p3jibU0w80p9Exnxm6d9eQ/6ZNm
sWLPk0CrPHu60tt+zwvNoryIFby61ji4Pb5s/bAaKceZtTSpW7wQ2SRMz2CJwIMU
nZO0Is64OkXV/07buH3HmyyfcrvtwJMjaGa12tUSOH7M/KSFb/FQEECtrwqN0eEq
Nd7rEuJRLHXzpvgKmchUK7aoY7QLVHSxmIR4FpK+xentofnb2QtvWDtYvpPkVRi+
RaV/pl6qN6JUPRGLYPRTgl8nsaRdQZAVVfkT15hG9dN9Vc453abk/v1Odsihd7hx
7flehzQXhR1V/6NsetUl2yUPGeuPuSjerStj0uaADlbYCaI8XtcOERPr7ZFUFj00
DuagdhgHX/FyJKOR0lf7wye6OsIIfp6aKpghWzWMegw79VVAkVMWA+f5o9Go+K2l
znMR3Iy0ts4VATJ7zNA4y9id8XmBb2JFznkRt8yd+IS6Bq3QotLgTT8LYbpoDE5i
9jYM13t95YxXj3B809CS1gn05IOqIXHQlINo1rv06cIs+rYpCGlZiUSHWt8py5Fz
H4D8TlzOdtpH2fmLy55kqGmhljy+c6If3vAZMIJvEb4sOvBBlstKMWAULKUO3NRr
Fhe9jZhNAHimhIsSedhbC9ali4NqRzEHeu5yC+P8O83ht4q8e3WUah+6NRIiCYUB
i7PJ6xA1MfHx0w1OlSWQwoG+WZ8yZ2ZYLC9DZZC5z7/JjwehChvtLw3d2cEf3Jn1
hKjZyt4aCxLB5SAJ3UTqxoF9UBz44QLqbZlc+5MGpbnmyGXAzB//CVoDY/IsV2jF
SOfbc/4Gt+0ZGx5+iH4e5HBehOg1tCKs4DQ9+7XtaO88E0XaZLMSx/TAL3oHq2fT
bQCB7/Ud5NJqP61g5obh/q5v5LOTebYxj8Jr6JWe9OGjWb6k42r73pspyJN4zfGv
RQczEwi16qZAf7tW3xacZ55u59wzoPCfb8orrr5lcXwgVuSthb6LekjFubZcNBiD
s0klmoTsArayfdXrM0Vn++/pjfpgaJkbRg9i+ZoOc3viBO4VXEwZDRgCnYk0Z7TF
kYZP09IenvfdLLPmbiAvBFM5/N0li8WFlGyzJv7KESTtymVVRXU8iti7O8HmfdYi
OR+SnWVxzll2XQ9Yhx28mIZuBk/SR8GirsBPXkRRVmgYt/CGo1kWjIcy7pKFIA9V
6rA6krtxYfCKaVebW7oU/F838YamnzWFnrvIOTJoIFD4Jiy3kKadbN/7ZBotV5yv
D361+dxYpFxBobDoZtkLvFYzaQlssgoiDHU1hYIaEAFSvBL9E36h5ynkR/oFGpA2
tWaPJ+1xWojlCYy2YESPoHx96ycOGy8RO9ArCxffp3psLPJsY3vQC1dMx9f3rT7a
A/D/YG1p5p6HrMEI2k4Rh1XsIvl/fKGwKGMMX0td1esVbRXiR3oQUfwFSJK5rqxp
ot3QSM9gUEq6G1Q3PwSe4nhxazRd/AMLT0U/vc73orn6FeSNcEHhcP7BisMLfXKL
x+/TztVHZoxQjZD5EPcRuB7NmYz7M6ShkhF5jJwg3YG4h7R+ZVWlEaKKyFKtGjpI
G/9BTGpwOwo1cfOMdCXOy9/U/3kB1YIoURY/nYvqgQfxDeo55ifHKd/Tvgsdaq6z
wdVFHwJQiuvCKxCuqVmTlv3upd7/7JHVuIdR3+T8trqUWYDljvi3xFHkgC1OO0Cg
kx50IIVC0ML9GEWVCN8edRzo4gAnrjq3/2zD3DS1Cnbgun2SkxOLextvTtdWfGDm
WBTuVFYIPHBuMg1hI/4DHbx8yYBWJnMxETsupuWENWVCgeF56uTsRWhAY+s/BR26
HG4l6hYg/b14xyr9D+oVCGRb3UDDshCPAbzJONu/mXM4807H0CVSIIsSXMaJGp2q
o/vC4H3KdRLj2cyU/AR0lkwFT+Q4XNjimqGxksSm4POQnHykES7DuedBXxFeIXQr
j6BHYYFpJKU2xnSMXY38ovlPKZqOXOTM+UiySrrz9pyq+MnN4JkFhUXxW1H/3Ijp
UqCZYenOwyIM9Y0hudC5bOYImHuCS+ltWpYie8H7CzKyPj8vbMVYv++s0YEp9lNT
aq/AbpUdgL01jSUIbmPnCvH110Umy+BKEiVxNOa+QdX4mX+HieHuRNbmawb2ZOoB
0tk/HUrSur3c4ReHDqGgXHy2E4mcVTmX8Yth5bQDqwwfkOvYMsmrcICSdK9u9Bxw
zhjA0ubT6VvD2U/+IB7NZW6YQIBptWbrusChJLgWTnaWtABozGhlmOZjDmD/qv/s
RjsrKtEodfAsY6DFFqQ8u8ucSVkkQaoVOK6DL4a7+MoTE9HuwVhlNY9JExaNyynQ
tzQ7TsPqF8VXN9AKild+b9nH6cLcBDQyw8I98RMFLvyAkaTfa/XYKe/Bt2SaD6GG
yOTyv7tzejW1fdfwdktwkrv6WGe1GufmQCyds147sovxkje0tY7LUw8PAyZWmf4b
tvIDlZQ9jXy+qrS0YsTa174WzNwfy5Q/BtUVLMzwbsJEH56nNi5Set8hU2MJ20so
IlTCVFtemMzymFzZy0T/kR6zUDfeMml5vZKOpSWQj/oeplVWUxH+IvcxFiWwUzUs
C06AiXbnl6jn3SXzR2xsLJgSt7K7gxUfQVk0PVaoZd73KUPhN9/49v+8TrYnQ1PM
1/nYK80B1ITub+wmuehUpG53bvgT33OK1XfjBGanxFc5MHQP68QFe7Y0v/qulLlJ
i51KkKhU2dDSzSJ96f843coxxVE4tgXRTYikLDBJhYQmpH7ulGgtrXhV+KrSf3LY
q/I0Cd6Q5pC3jHJefusIKwlueKmfaIgZ8mBX+b2UAY92j9APSR9wpG0gCUPiI4pR
QaRNA4F9FFV6lXRLmAqutfWmtxc2KdlFbD5E1hNdEtXFKmNqhaVFSR3gNoMEAlqN
lA8zhC3B5IM9WBAW98DXLVRyv64pxdr7vkWeUdGaG7Wedgdfoby9jADhHbZxD+VC
WhJ1hYxMSPXqP9tT7SJ16nrCpwoYLRBiGLBN1ltfm6NjQ9biO+DbIDGcro7YBKII
dJI7j0U6z61xFQNiyrsu/sKJn/wDWmsJY8o4iDgAcAYIPDlidjx8yps5E2/XUFOH
piwZrSYi7mRMPCydZyAB+yLxF4lys7sJXlbj4ZyAvZdgNTGiXbrjTduRFQuvi50j
IJ+wZ404eiTXjOGSiNSvHw5qa2Zd7intiyoLi+FV/Wjgw1Gjb0zVz5MeLCkpKEKr
p8+hgqTpTnyDgkvQGFDeUYScQPOgTc8DEOHZfXfBOxv69CyqPcHs+Yt//lnWssB7
YqLQj1NlKLQLeTGD7ObTqKCQwK6aXghsJKIiTnF0r/qkSI2kVxIpsxHqH3ZnrfKA
IM73Ntxz9tsl6qIi0yDtFWndYAegkWtI0g+A0yyKY5akHV2yXGtPHTFr0WYbkcXR
yM3866rOxfa/s8tmSBwrdptgXswmG12nTDobldUWkAlDoFamGrcY0nMK4Ij6Ofa9
KtqLPePSdkq7N1G66e/TUWv2ty7LgXU9AjizTL1GNreDasUM6YyTsC8gMXsdTtfe
y+Q+NP8xRni8vsNB2PoFmPjJ94c5JDz9zGbB6bCrgO8EL/xaymOMehkQF14izg/r
GVI7ECf1BqrT+6PT7UGq3fXDY/ElQe2mCKFng7jp1ZZqA2NYOD4upDfHttAYP5Jt
u3LFwxzVOrWLg+PEt5mLDXDRRQj9rs4U9704IMBpSIAEDrBp+tUredZ4pr5ABDQ9
Ly59o8OR9kX5wcY/OMHG9J/9X7CClqDpxe/+yJ6gf2DCCELcu1cno3GhBOvCrGVM
yArZa38MgQihpEeG1+p0BHBxLM3REuj188wWIydPiw6vvDcxANk3+5IixBdq/Z1P
lnrCc5Cfrup3vawerqGBbZ1Y7j0HtV2Ma/fhxja60tTHBwMOTF6td9OzNkRChSK8
rcDM97KlntczlpbI9H+hdui7Ca3bPo/5QkoFXzdFernBbk7trTr54+rskGpVPzsQ
dxbZw10w5LgQa7n3RYtHwbJ41FB7orvbYMvs1qSRktGmvzge8asLitw6qG8mlwsx
RikUQWaF4eIR7BUn4k1jzc2NazMn2sYFVwIVKXrRAnvVdJzLmLt36W1dCcNj9Xp4
eSvgfzUXGUDsEti/ru1uDeoYm2ow68WTDKV+91A94ox6JSvRlIwPtlU54hH1xKY8
vf5SKdvWn9KF0fR6RoHOuLknk2lvgp1Abd15/IpbsxV+PMk+4HrGnHZDEh0XIEiK
MTEfrUrnBeTKBjd9uRPq39Hn1KoatbebhjmHg8XFSfNcQrgXRP1c+yIbeqrY1hJx
YpucK5APisAVvJo9V0gv3AWl6Fms4ij65IoLfTa2itTtJ9Afur1YyuKthp3oRnte
TOtxiSDqixVDZZDkncDHy6NFrPcl9DPjbtrnym7Ym8geIz3lBjD9mbOgfj7zFaO0
Md9yFsK98AoQ173OdBF0b7CTc4OPCiw+yrCKmzxl/Su+2UFbGdMaP+tuZFJPQ9Gh
VbO0YSrHGqpRonz2MFlsnoYbJ61iNVZ8xohrqzhRKd/4+imNG2GXpLGAw+mlf7XL
uUy6E7TSo/YfeY0rhIGowjZxnAjWsbaH9IqnyJJ54nm8+PKTMGEyBOhAsXwrenwA
NLoqiIAPuqofJTENEXmuVGWZNrLb3XWUm76jxUCf7bvabbLwxpQiWTV1QmH3pMUk
8ZAUyCrjsCq81AWUi6blIGMsrfUv9Jgyy8UwV7q4KGc43X7m1Yi2WV03XLdqsq7J
szGIQ2MzoZAMPdxWyV1DTVeC7FNV86IxkzdBsT9vB68Rg2VOf5UzjcbM49qHGLuC
9lSZyr7NfsOEt+zo8Hrpp1HeQvvc7jCvYjKi79xx6/tEc5tbFVvs6/sOUR+txvLr
nhqTKBN1LfmNPcyktOr6fbxNxyIJ8XQ2FhhSsO4agb030iTO0hFH5tvfTCXyRkE1
c8lKtDUAl/qzUlGNXkwbkfgULMEMVnXME6jYpFdW8ndmzI7gx9KgftHLydnSstWY
zx7x1bM5OfaWmfanLkiJXa/hjf0XICWk9Jf9+NdMHReTFMETs8Vc/RPScmeAqli0
5hWQPGqEsnt/Ye/jdiBaHcc+NT9VdosFoTT5MmpZNux1R4gbVb6HolXeWUsfVfhd
tyCl9N3B/8s2CflRS/0kvgSwMZHwGevE47vfa1GMGJrgrY8g/eNeA3ND4u0AFRJZ
hi9GJONdU2ZZy01CJn6Al7YtqatjEdG5GzntY0qsvI0sZLnwmxjsj8otFzWixeFs
QVXIRLpOsBsTM7LSla++x3eDKY7qvE7OV2ACRmIC7G8PCgv0EtQRDUQPGZTSBL7s
KdgCpxXUXwA0Ap64h8DJAB0wdWLkJ8Ra69dStMyUNgVBy7l50YGWt+xU85IA4JfP
myQ/PAQcTBjZhARVP0r9MxKOzdgkpuZhyJfgQNsmMJu57JzZvPiapxYZ2KHNlkXc
VUCtKze3/pgxfAbKDRqen//TgwqQJNKIEHdeOF2RVqu0LuABrfKfXsYdSsFfe33q
qLYeEiUV3eUE6Urdx7j5qyt0SviNrBofthcLtF5xwWoT2ICcnsCRpkCUnSwF6Qa2
AOMMta8pb5SMbr4MA0KQ4IX+0AmFF68+lSeiLA5KYbTMBdR1Io5Wbt5UJmRrJENL
87eA5BI6MxL09sw6pzcQVQXlkbGmxQw91Qay1WrLo4ra4vtG1w1VijQWPxjPxXhZ
hlpPIhN2qNYSQAQDdfCfn6coW3JcWR35vCXK6xkJ9yZE38PnZk+L5aQYUwOZZ1KO
2ykoSQAXOFYULj7CA9B93urjevfiveRrgeSXsiLnz9Eu1yvGoN6q4pGpehfQLXaU
dtJOPtvpHEeFp8SOfW7Wg6gJcpnuouvbc38g1LzDbdhGu6S5W8QsH1doOT7M0Qtq
Hju8mLysn7nm68zBPFBJ/F0HHHm8wwJwOLdiVP8D8s6QWuGxUZo1kXxJBpolra0z
9QZ4oFK38RirbjLIp6OAduYbSDNWEugFmAXWpVwlX62ooyEC5T7zCWyTi9wnMawp
2x1CdWuaCu78hjMY96hNU6/ERJMqjbqYX2zV1NoleaH/jlOoXxDp/5of+2IntNRp
n9sL0wsRV3+KI9AJ2QxrUkKMZrjxOUbZ2gyhkA5T0bLlaeEGT4BlKTR2uMRUdqNB
r2sRA5x1mD10qFcx4k16N+FL9sIcl1FBsBoe7FXBAX2nDzg7MXyx/5O33TXCuSfe
8gUMV0hwnYZDb7HpwUga5WKCgQ42b8RJjPg880XRBEOAEkuK7c3irGhSV7ex9wrJ
9b6zsLnFaRQAZo3oaK4lcikKJqGq0+AoGvWTnI1bgaeqmIhmph9eHgxFuoPkTjy2
oHPkY8MIAOXPUME2PG/CoG1AyvcHLydga+QQBwveWIK/O4aKNFK7xpOhhrZ0bDT+
ymt3/V2+mVI0h0noMOQZTYt5RbvsX+mDCDgXNo3wVjv9o96pxad2q6J+YlE+yDzB
poSfBqYZNF4m6r3mIlgn0LrBbk2OfD8HP4cETUqGVmsS9pJzyZBArn0ePgF8vXzH
O5AYGFtM0vB/6AlPYDecHdSRmpWztqbXBLP6R15NlefFjEQJlJTSx6vWY4/aoxT9
OBn4ReIcwwMl76ZLZQySVdHz4M0unhirIwH1E6kA3vjreRw8Hj+pV/2kdKZHwwpp
TpV33wZqIC9LUCSgRkmFoJdmuAFj54vn10vuH1w01L6KSEHY36J65goJtHeSVj41
Obnt9hDzmWyCAtLN1uHqHPWXhQ3M2z6IFj3kNjOYni3LPzJaTDbaeLB9ee/OnJIV
JxZJUpoHNQEgV/zGXtPzE27oidFQS6QmcmPq4wOVAw2qxlKLaP+XyLBlWjOnl5iq
PjCzb8tJgX9z32MDfpxhoSvZcRwvshLUog9dJ0kodAOIelGfmM2Ed9aDCBmZx+vt
uJbaEKORatbzsyZOw+jH0QCmWQOHLKxkZ6v75igq0mQ2CCNAB19qWYtjMgoDmcha
vReKFXtJ4XLzBiSwDRyFilq77izKNzy1S5LUTRfJYncxFrPrOVf60FhzP9Mqxj0A
0QUbikjPEiTKg5ugwiwWcyK/zc2IzXrpNlSOat7Xq49IlDDJdt4aAjvXOfp7AF2g
xbJMRGNyZWFZuZtzvnPc8NI45V5/0UgDYf9chdCxrOB9KN50q74P4dozfpYu/gUb
fvSSaSGigzdpebvc3Hzp99Pwe9WJJFfr+robzYQ2lAGx5fO8BiIhE6TEXXQ01P7l
QPOaIc/5b93m/b3DOxWZxK7MFqrpcfsUjdd4ucmY4By9VwKUEEAl/pRSqk+D/vbK
DDC3XNs53llyTzARX2kcZ6XDLnNFHGyIunt+5evuD0HudvorIFjozGR7Uv0GKWHY
ZaxzcdqMRmmwps1Y49xWJHjrultNe4Ctth6dhCE8HyOmePl9PcAfVpblduO5AXsY
IRK72JUNXGTeHigDc0co+csx2d6oUq72xLdHZb2PjVB6IYfJsZYK/RTl2KLp5BUu
KoqbozsqviKH/a37OW9WR2I+oKVVIyYDGZE2QEtHYYQhAwIb1ENkP1NxrY3BM2+B
EJWqy2j3xisKdVqNwJuiUvbGGAZxiNfHWwQVJV8jVCKKC4FtH2GMIesEwSDBf/Cp
YWwUtKTV/qRe+7mgETaZ/I19qZrz+8BUnncCGJAe6JfV8d0PUIftlhaiDgzLnviO
0++y2Fbz1V8VTOWjfoqUh9qTl9dq12A41qeSL/cZR6E+n/eKSE+zxXTISSXN3bLo
q12uw6s6NtbNfnHkvVzVEYRyrhHo4vPNeO93QGlCQs7ktoaMOLUK6bOGW0yO4baS
e6m1BfRqH0qbtoIj1DulvH8IT7G1w6CXtgsQ60Rf6dWfOkArqDp4zHgzf2DyQU3H
ALL54XZboWOG+SSpGoc5UEyd6wL7uUK9n0Y/73DHirsatuRK5U8YW/SOdnPEFa85
RnSFJZUx3uZ5oXH6A7zHofeWtNB8V+ffOt7DUYI+EThFttoMoXnJhsS8lHCi1bf+
8ZybYJxyzY0mADkj3sbXgawjvnpLwMKTWSaxD3iDSR+uF92XuUqIZqFXvOzrnPSK
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
LK1+pPRfHHgj6dZpD0lL2iG871knVdEgRMTLRGl2jDLirCFYxXCd2fAbLnu6FoA+
wj01TliYg5wqd7eMXuT6IJoCgCoFlQ0twV3FrGwvz5zVJgxLBNDG28g9c/TQcQHu
88YhsUeAWGlZTRguvP83nyNaJx+yKX8qfusHxGVvhDA=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 12497     )
NXEBWHi+Ekbp+w9nza5jIn8P1l1LV7nx9yE0ncBA74uEkHN5pPt1sVfPyjkRBonL
Pk7t9TJgn+RxTd4+MPo1dcv5idsgfmWIGDVNH8yr+GWoNOTWINvpcvnTAHOM05Xt
w+jYXGrHTJy3nF5D1MBWBjgVyUy3g4Ei6y+1HaUAz0HR0m8XflSnwA8SYpJ0sNta
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
jc2abQN2VQSDHIYE/zVJaEqqW44YDynspGOeZe9gQcEpZjJ6ZpN6V8Fh2UBuAJIh
APYzqZiLGlhEQG2EvbtAQd2+Kq+my1HrzJQN3/0a9DSSwvl2T3dR1ydmkpNbMrvx
zQ6fCu/HnuPBV8Qoox0jgbtwE0Y6X0IkMj9k5rzXsns=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 79714     )
vi0XB39j4E+/oNGKefxpNsySfsr+IIL6LOx1ajltnzkiD5Xjvc37C0TJw9eUesgf
19eaDBDhoh5Vzyf+23eV4jCX5HVxQh4VnitWusGyhb6IWQj7vxx4yiASjuBH1cYk
kIPwXLUEFtlSmltd/TICuj8Wo0DbDk6V0Ch8vlscvsmFMmx3fKdl4FMcHinOxsVM
j1Bsi+euq/Ky4DlFs8xLepBR8I9vljya54dfDOq6765wftLfZKMp8AlwgZ0jn2jk
Gi7SE09kCAMXGS1Rn7yhC4y2Qascvktv0ftqjyJ/NAjIqjfcChy2dRzhX8bpd9cj
3Hr1NDkumZjeWSKcKnGjfqwkbTzPHjA3GlsGMHHv/kIjPOcityL61psPKzu4FzLi
+c/8cyF1OV/9tyHycbN6VelSwKhL99K46YWr39ZieEL5PB+BKp3bzXlofhxu1CGA
xdcRv1dB5cd9nUK6rtmbB7y7J3ZASD5AkYytjGgCcq/pNFGDwHNUEv67CPrCJ3wl
Iye578Q6iVz25i96u0cWkrOB9kvrLgkVPRsaXIVfPQmarjSf9OrdPDNGhRHywMd+
55evjvR4UFRWYYLrlqOBUCpvRgSW2SbhKGbkhsZ6822+xlt/kIfOSVODbErO+5WU
wYw5+TLZ9epf+0n9l1++FaqMsBVm6E5fKtmW8A7uPN8crqkibkdHTN+9N/kuynDD
3gzFzzmq5m59ZjP0pgrpmqrln690oiw+/w5eVJuunnLKOewyDmGEWtAoTdc1mNXP
zKOHFW/the3Z6kkQDElVfv0svL32MXGphi2/GPzTZMlWKUuToauOaSoX4XHNBHL7
BmGdcRuoJloc9/XPBuuHLgR15vdFp8+L9tni0nFFiAZOjymtX/dCPymkJsv8B+XB
0OlyIjWox5Zfyz1/9KlgZIzFe6vFFKPuAdn7oqYDYS1pU3Ke6M+t4C1rEC7U8+bj
jFIjo4hZB3I2LMT9P1ZEblh6J3kHL3qKYerl0tXVEEWdBh/ceYRHTaM+rdIO9UM5
lSMUldwBe8H1FKJVQqmyJU0wyuxSxVQJCuRHz1ybenVUvm6ZrvJDTmtPupXwGV8i
tyq8YfPJQA//kv1B0/g+Z9u6RNNWIazpF4IGBtBut7dmczh28/c47LU9m9NBOLV7
z1cbbCmydOkc0+uxqaRiHhW21UtUuK4Semh7/zajErjJ7RrXAtJW/VegFRV3/OeS
gvJa4smqf2mkl3MCBSCkSGbqIKTUcg01JeW+Tit4eNt28AJP1zlOSD0aclzTCXSj
9UL25sgC8E5oTm/Wue0a1jBLRomE7bYHb7s69EKLOR7gm1wweNl3GAF0y8PyFOhy
of/T9Wpwwu12jtqC6JtQBFlhjLZC2JwFfGCMPVcewGnmMYo7h+jC8fhD+3+MT3ei
5TIpz8PUIDlZ60jJn4In1DY1ZrU0wdMmXoA364VUiP0hgo4lciH57v2NOJP+gHGu
UurlEUwGw532rjjyLxqw688JnzCLFWPPGwBsHqBpRyZvnHKgYioxpe1Hz4CO3H/A
ubS9NKmJYsioUN3UxaXXsqjkaaZRdzwvnNj7a0dZ+raJWqZ1315+F5MzpeiFvGH7
sOnuuK5PFDrKM+BaNpiiZqvKn3z+GFQmelHHLLsigeqfeSjZQHjKmTL0JNVh4oCd
uvwx6pHmAPDj8SsQymn5wdRzX4tAPfJqef1El6zfFdvg3MmgQMx+QBJ2b+27z8rM
6KM9c6qjDosK/QA6KzmOQqxEK3xFYJsKeUt/UR74el0gFIREGjXe5oPuWnz5Gw4T
bxsiwuRe2HPA3dxXsqQ5pZYeE0J/O7zdL10fhn4Y/CYZ2eHpQmZSLPZV1PNeAEwL
ygkK+Y+KQOHy6sYwBIberdIzjHT5vFXRqfXThwqH+f8rEh/VPrVyg6UKmz8QnH7j
qzYHC1wu/6UhPqsTz01j+qz2AeuhLCC1y/9pO5nHzbkKHNTrEY4tRrpYB39IT75c
s2VEwUZSbiItDdNG6wBrbQszl/SZlslOg+ow8MigMCjv3z/Z0mwdl+jrCeKI7cXs
vKY0roGd3T/XQgUtdq/xGGM9VaegY6NnUCN5JBZCeDsBRUNhnXSfaOMUd1FpykmR
M/Xa0MNpxZM5dJ6aNxSTezGTOx5kmEMXsPd1PMShPuMiVSK82l0/kxHEOaW0Vo/n
Ua/gPzMov6zeYDzQs8cOgjWZSL4bNz4FX/Q4erYNfE1tfUcJ184FjGHxlEsiVhvX
18jYzoOGaA4OJX32V33+AUtsKuG8zbFz0LMSFeo5p/QkFv1iRQz+Nrp/QQL27Z7G
EK8C4RDNCrR2h5e1/MChOOrZOshvGOMy7Qw939tM3f4XDDKy7ToJ6p9dm4bPVw8Z
WCMzWnHrHHP2wKm3IXGVj18362iRrCnpwuc9fZFGktaE0vGPgNT7SgNtyberCOX0
2ykhbdDz1BR4hKOJXIf+E37Uic/gqFAJJ/0Mx1EOAAvAGwVP7ttCDNtrbxnvMrId
m93sYnWejQ4K7PfvYUBTBTGi0pqGUsarWZJ60XqfhU2yXGkdzVwaPeP6R+8FGNlX
IWeGIwsakx7CotItxS+NbA/5bBEzBRJ/rnPooWcdjyRKM1hJ6tvRCkvBXXnI9vHm
rKdLA3mrLnQE7vZA8gogSh17d68xFxozI4OOOKilJexyoxvF7SWUxS3snen28zE6
W29FAO2akU3w5IeCKCgbg494HjRagbhwMsh9f8PKU9vvJMZiT++aIdDODneWzRsN
VecCCrIY0z4C55sa+l2kDL1CX3bUaLZvhkex0E4MuZkICo8Ac9yWTDPThhdBlYab
caniMmMMRPZ1wM/KdYDRJsS9Qn77xIDro+bEkZYANJizGz/RKHklVIzAkZWWytP2
NVV3s+K2hdQkK/phnNrsnDJmyZurQr+YdThGvQsDDNN94o5GuK8weLLrAoUBGWe4
pxvMPEXQY1TXFyGe9YRJOQSLDnnl+m9AgLGKTusRgIXkGd15A2Z/xxXG/Mg//LWm
FZmD34s4yhSHjQd26aJy1L7CP4obVhHA6j9wK2Lq34e60WQW7Ny4owvuW9Js0ybR
6HSboAj1ZG6oXwv28ug/yBCypBZ7McnJJzQY2FSj6AnX145IO6rD9JWgOwuoRBIV
OvVm/Ht/xg1F/JOUpspfD6Zxl1QX6TjNPrXAWeDO6Ko+GtSYaqemBo8TvIYTNQa/
AxbnG+2/S6uOLpyu5A1lVSOxJFTl8Ob/2GukyxBy7mCbkOnJ0PTG+l1xnamOlJC8
xFLuafq0WTNa7BTlW+SCBK06/vHrDW+g1qtxJEnxqtataWgKhtkYFHFYZwEvxRX+
RwBzKMEJqMNOWdUUc1MDVbRaZZ9dSg6X1WCvVw9urSesXG3AfHqIHI2E2FGHZpwC
qlfxMYMjWeu/4gWn52K+o3YI/VnyPJaJVm3vW4ZSWT8IRjv10zXznM6higS+lXrZ
4Ls1tdv80ooFC8aSMBM2CvfnehfbCnaCuU6vKla0T11ASmLimfvT+WQhS8vzfu8i
n3XiNoo1DwruSwzIgS8659whvaAsobZHW4FL7tgAb0Yv6SUxcqVQQxz2LAC5DYDI
0jBHC3DHJVYGB6Epx9RZ64nY5p1mErSdJg1uHsvLsezci2H8vscbfDcspr1Ajqgc
5dqMtUpUfOeIgEbfQvjBGUjDCpH7kbHYU//uCigb0+RleUgi7wzIz8EPV6uI+Mkg
YPJk7YPnf87WKFYP4LWmATCbg/gwrzTNgK1+BxjHk23q+kyXgZeoSfdp2gC4umlN
LBTSP97Y9v48LOPr7YsPoueWnhj4KFd3+HMvkGXEI2hGz4+/iOB7Y/Isw8yGBSxV
/tDLi1IKCZw8lHOADAc4Gti7BXtUWerge8Qb7KAIZ/wVX+Xdf6kljjUEDrJG/Ci5
HGINYeNC4qmCUJ43DTkpDuwsJXHzwMhVgeb5w78t8NNx9FbNUKYX57xlfgLq2kyo
lrHaGKjLPtDgEqA4GOVYkr9ZA7Cl5UoDBK3aW6IDOcYECBmVWR5W+LsHAcDBHZjG
CzLOeOb/BqnB8EEv4rv6/xD9KpPNBqWMTvwoVopg9iN7JAwPbZytZO99YDR+qHFU
STdFei/i4V8omrhaU7qzO52ULzbEPvFCpNWB7y7lERJCazAud7DCZc0diMp2n7gC
0st/HcblUWnFPoghYSi758Nz10lbUf5bK4mhoecT/Yc7c6j1e8Smw6CWX1T+kO7U
dLGvBDJm35AivnKqMrhHOqye+RFx3jSz8Rs0r47XeEJhnvXvvXrP9a2ChQJTVKdF
PVHoUPlwMfaBzSunWnP0yIgO+t69nWK72jtWSx0S28daEUnMVFMJNfixvNrP8pre
rhUGjosmuwDlxXQsfmHDFy0HTrqh/sxjUbeMKHgXwnPrx0Q8Fz0SWKjP979id4Ek
S9TjjXLUICf29VrSBQ67tcZItPkVu/8YbybL/5+RiAO4C01p5KhqAoGXZEiJk/VO
McMfZNPfPQAs/7WDHqa0g/5lupC7xtLXnOP375HQCfyRlLCP1vGuMrlZEz3nqIgk
VgqiqK5FsuiBwf4X/VXsbsiqs87UlPuGpSSWjGNUGGN/YzyJ9gWoJTegku6g2A6X
t4cfnXvcZC6sgKYxsG7qki1dklhv8pa1HyLnKmaiI+QKARRf/PmwVxQipuo0IMFH
6+nECq8nyt1Vsyn/wJCJllsJep7dXuWmt/q5vaPk1jJvnb4SrceyGZxa96dE4y8b
4kWP2QBhHUwzU9kRJlgFnTit4S3llSZyG/Y1o6+GqnSQiHXc9RBCKowEaS/8lYZb
MIC3TFmnkYbbX+s6jmH8SFGyYwMQ5OtoPjC79zzMui0GPr6avU5DL6J6Fi58H77o
X4TOlA96x6fF/dJDlqIBMs1aQ/1J0oGwbl/ZdDZeE1FYFth6TDFgH67Prluad11F
K4RG5A5H273YHjD5x/K39WqTnt6INsvdxlSM7Dti04ss+pO9apVFJk8OBiX+Lgpx
pfahYRuBgSY0CdahflBN869omSxxmsawVmWp5lgmNUg10fdPmkxdihwkY2IXyOeA
Vxb0TNgW0lFQJ0c/jNl77QI5cREfNUaqlDs6Q/ncdjOq7v66/KAt2PyaH6Hcgz+7
pHIgc3/W7Vmmfs2GzEqLVbwkhyjoxbISfjye9nRIFneLgXd7pcTx+R7vr2SH0/43
TH3vlO86pSXpMW51EmezTmE4pPRu1LdHZfLXEvsL2WNLHv5vUUuuOI2YbR3ctt8V
smABYBfF0TiUzp/ZWoNgtPg+lsjZgmrHCrYeFU5bhkmeyT9r/36VLGfuCD1zyp1a
9Ok2dMjQgq/G9MmawCO2bgnQ56ToEreY74jD71rG2i2N0/3fB+Ns5uWyrzb+UnDL
xW1WPBFytim9XBRzpTwHvc8cpgl2QdfeilzHTYUull2yF13GgO9u+mgh0u9n10gd
WMyKpkOVp6MiK+QmlpNxgw+g0VS9Z3UL8Y28+ABa0zqk+lx/0A9I9iMDPlClWIOe
YnZMgrx503zoT4RXWmvlYjbEHpelXmV9oC+uR+K98Z7XUBWwEKC05N6Z+X5H8Loy
kd+7HetvcWyrX+CdoqQhaETjaNhLFysh7E9oj8KVRS9kYoP9qMjoDT5pWGAdgba6
wpVyHMwdsDyuEXKy/pkJAkmoQJEeGjUudGkJjcsU5bicChOS8uu/PDxOSbgtfjxO
lY9p64x1EgumaFLnGGS33UNC8tRZqFSsz8bE87UA5GTh+c7CzKPi7lazMOYztTf9
fD+tlAuLvCLHjMLtz+M9+7fyrQViozK17BBz/sCXas9EIahmprweCLy7vY/iqswE
BNT8amYTYyL3ctFveaPjtKJXqTYGZInkHJ2btqmDROiIV00G/VxoZGcjWrt8loYf
xmGYBtGZh/cLtaieOO4sfqajfkcQoidH0ZV97zkyHb0bgOjELmHxMtApIEaKY0ss
5dPzbGIAa3H3J5+NHEr5OvzJL8RUM3B0m6vfRgW7AsHAHBHYmBQjCzSFbSNyv0em
QoSa3o2rwG5XOnp/mzWf1X9dFIrvKK0NkeAbCiLRoa63r86GHpHqbR+ApB4BB8s3
B5evX2YgaqmhqvsW+Ol3cnbi/p+QWtaK04NANwPNH3DZSZWh9rCF23pNAqXm4SJP
NXpY/cveOPpvfs1kM6SM4RliR5HbOdBQhXNi72AuMDVuYTQYbvQ871ANAWqktF4G
YnCOJberFpDcwnYoY0OhcGtgQtc5luyjCqTob3DbQAMhd63ZYgd1HCZ32K+nI+oq
Woa9PxZ8fYx6q7bsHcRQMUIcaWmgwr84nc8AFD/2ZGOV9CQPBPOeBJuDMIYSNhSK
wR/5Lz3LIM8mrkDL5xH6z8orS0+2R8Bf8eMJcnLD1IG/y/bePvJvV6okispwPq9d
dmmbEWdZVkaJvdSI/ZC5qIsZZfN4z64WbzsFcz4/GQKb2Melc6SFJNtuKy3K7WjZ
DN3Uhjv8TzMZHjrzBmsgUTSPlaxBW+b+Rx+4uAZzqjqoHTZcipNvQqpedw1ESRHC
B/OPbpXCL7RY2NNye/WJKo03e+2Mb8Woa+5zIFDIyqBZOzw3IYJ/Nu1Bc/tfXDZ0
8StAAHXo9wy+NiG5vLVbRSuGR2RRa8pxJi3Tj6CixVwj92p+7cZR282XyZTzAwdk
aaF+pVjH9MNdEDzeZXUF46EXen/yfb+33DMPIvUPqTtV5t90n+YCjyeMckVWGua6
QbmG7TWTFuxvG01d2EQyhDPIYaLNyVCckrxoRriFKNkHxYFl8GQlZ+gTU0I58Gic
sMn/BUxE7VlzyYbDoidGe9cCo586MXNzHt0k704FIk6b7yDvHvRT0oUuFs+bv2Or
roh3YoGyTAgveQY+Q7bclKvWVMK/M+JPeBgsNgve6zatTi4QhAn5LUECOS4zrN5D
RMmoXmg6y+jQnVj69nVKykJ8fjOlf4yv2ofr75Fp3uUJ3eE0Kt9RqxCVryZ3LA0A
2EJ8RBSR8M1qnvprx3KQGEJwxxNKXpBB3TvGhDAA60RB9JC3SrHd6l4H/1xavZXr
jH5jWRAILZc2NUszQ9kkGgDsuaKWOeW7/Cj9PxalOzjnvFFuk8b1YmEFcVRnwfpI
RJ2oL6t6ShwE9nukYSW5gAjjbL1Ck5W6fRDJbcdqdYsXjdg7X6ZkF7/fFKhBW29I
Tr1Epy2eUXreNCxoSLNGGB9oEbhptKSqAAHhiT2cHs3gg/VpDLsKUjQzz/jLShZY
b+pOMBP6MDxOiWB0aYOKIXonmxyDqh+cAs5OEil0AulxM9LzQ2QJBe6EYCgWu1Kv
jW4VLJzRplOk5F42SGyYR+B9JfGyFzSvm8Drj3YPWK35H2biDjEj5cGfMsMTyCAZ
ptqfKDwq9aXIMhCvA42OLyMuhm+WQnw/gtoBavD2pz0dfL6/g7o0o575vZ/oPyG3
07GZ1gjoAGciYe+6eMJlYnYDTr4KNaNe0MBihanAGqA+TyYSL/4yNmLoOGCC0OuT
uscYsdFHBjvyzQbVh2Y5qYp/rTq0n+TBw5jZBnJIbWeXNGX+AyCnJ3jOnm73mxnf
cRrWBLKfylNRSF8jECXu9riLkfXKjEgdj03YWDknW6J4A3iwuNY6t1oXJzcu3mdv
9iVbP79ZXRxxGJF5ZosxiEfsaG6kGNWxhkfTdzyxSS0iuWp2oqBBOAy3UT2ssHv+
WG9H4Hq+enlqzOTqUG71HrQmcid7ma2IgNIZ3DRawDq39X/CmYECrSPL0G2jbQ/0
I+D2dgT3Wj9osn2mo94QWtcyvSiCeKpnmXNaSvCd/ZxaFK3qDmOnhlsByG+MU8wN
xmQeLaH8McLAesLIAYQIqUDXtIWcQM28+qACPYlkZjRKK2vpR06Wb4n7akK/SdNo
K3xXzyBLxb8kxxSAr9rAqZMvHQ6R+KGzMiajSmwrOPCyoAiwreyyllzCIaX2p07v
QCXRZRKjoa7tmDQ6QwogtZDVjQYEkA4HQWypa6fnGnswRKiEwx2xU5IOcvKbx0Yw
0R/AS2rzAoxHM8ctSQZdfud8D6rwwETsKjBtVEjCfr04qhPJW+vCxA5VvdGj1pIx
KKsQkFiFqA8+HPN5U4f96MIsdn3DZi6HxpLws8s5tU+9xtxt82kYoJR5H4mOCh8t
q/rCw5Zk29wkDkd7v+cUa4AvM4Yr8Y+hgavZvAq34nS1zK2EC/a5rB+QsHpzIuLv
JIXGLjlVWijonnSFC/7+M0nvWY5NgGratRxF5yiBMHB52+Uk2vfnoS4lc60VCV0N
n8B1vX5kswK5IKkNf49SWvq4Rb7pPxweUyqxdMSmQYf6kgJzpiOpknWCakVJZoj4
e4GSISeMbXZ34FjjxHI9h3egaIyV5tm1t8+UeVC9yaqUnQsm5xWIJ15G/IgBuGI/
ZsJIRxqpWdy1V9c5kqQ1qg9rQS6qKG/dJp3HDoWlBLRKMuPtU/uv5b475zniSta2
cwABNbWlnkM1tPtpkLigruztFLlbMFot6rom6Fd2krKDhFwwHDMKkUsncl52RI1G
iPOP2wypSq8wU4FJ9AHy/JbQ6z/g6fBkjASJg14I48xrIznGSiUN3P+rTQsoh7tZ
sd3UlPloUvmLGGEHIPOwF8yWpxt5U6eL6ZfYxL1T9By6jBo5QiDl1ppjLVUbBWr5
fUnJL/FLUdST9k+sC5oKfjoUQHd4R7kwVLH5P3AvdJBMNOsCYyxCKzjtMzkmkRSX
KotPmV22Ip2SdcLy3da7FKVmODg04gI0NhBOUKitBV0uILbWXR0DvcvEw8L0cnAk
takLvn6uPq4M6XXkV9dj6LZJW81wtS0gP8K0pOq5e0dFlbe1NkXE4GEXpclxC/qK
jPZn2T813eGdBN2hAozjlvlJ2060S4dAXBIF9aks0j4HYBVr7fXHXEWc3goGjgP9
AuI+LV1npSMMbA9gHOceSurXToqPdRuRbDniNuAxj+op6WR7nUoZpcWKE4ZSlxox
j9i/mB4javxMICVj4W9lcpBouYKIJg8xuId8kGlyLTS1DqJ58cv2LEjeteM53UjK
ir2+TqEKKBhCKh1yMiE53EFY7zD6UvTIs3d+ONs51rG+MBcpKtejG7AtiV7JZPYk
LCoj1Ks1WNVn43xNSBU+XZbkbmNOBc2AHvyu8EKgPiz/OAmnoY0V8uxwhARwfEXB
uRC6tl+2/+w4w92xIWaLo9SgAuTyQkilcRvUmpmLjRH0OupMRveVb5+rGOWym/wH
0T0kOQHlZb4zINgJovnZn3JwbrE20oe9ZOYOvlyq/ZGTeqILodHoZKAkEXcLdWFo
Fvi+d3KGNJ9RAR3yNW6MFKAGDmYAEy32ES/af4PGY8DSJxfYMgT9bvOvNBpN3xOZ
wRW0HC+5eqsfNzHj4nFQcWtn5V4LEVt6M0mMdHRPwMNcyBO+9FUUV4Ej8sSHKmvT
44YcJvgxlDj0bb8AyPk3FqTun5BsnrUVmo07x9n2j3A7vdt8f7W/mlqk9ImNGJ/h
2CE+shteTTuC0gpf4pNWE6P19/hDf2AF5MB00vVZjc79UqPkUpcJKWRupA0QWIO0
G4DG4P3DYb3wND5X7ehAqP7Edz8bwDeo7TVPoIW10XciPq5ZkZu0kvJ0oRomvY8m
bUvH3JPRyR+pZVlE3FqSKnps8uZhAYWXV5xqqpH1VKaiBa9V8SwBnXEMps36nzJa
HyjpyOzTiN4gsUgLO1v/qB3/J2vQBnR2XRhsiIhGy3R886NjB9CDcI90ftsM0ztB
mUIAGvsJWM3ABwIH1Q/XlCQhZ23j+dkEn+JTSgMrK6vyEc4FjpbBMeZzKZIHcq70
s0+ZeSEoHgi1j66M++SpE5jgXvNzgqqRZp524qZHHbXCvFFdVS6U7Twt/IfUZ0mS
zrjEsSyFKeDUj7osr9WuT71Oaw8NQdPc027iFrUZ3zc9Q/ngdhFpGLVbvs9II1gG
fNNIa2UosLJdHDa/4jRLR36wAEldKds9qlc0YJJiDYpUcZzNXfzMNpt+2TByz01O
U8MphYDro6VgtTu5ncKRm2r+bnyaAPHZAku7dyR0/oNr9vO/Ee0BIB31cICvumeN
pv7iAmHIjrTaBTYbrjLs0uSwS0QBSS8fdmFC6hGqWuH+zyjOgF0ujpyLy0Cf5Zr4
+dYfxPR3AmGYDb+loxNo+ahudL7W3c+y4SuR1Bkjy7oVj3KO1Hqzzb4wiVzy5Nq6
bwIXikP/pBJhCg1FA6zP3EMK8eBx+qu1KspalZbtg1wZW8viFmcbpWzFa6QMM2EY
5RZzBXWs7a7TtNyf1OB34quK6HMmwgw0PCjThA4IqutO9gtFD/NB8Y32cf2wub7I
VhIAN3pRGr7FUty35+hg6Yfp0YVWHk3Spc9nBHTfref54kwGPQKb1p1LUzgIAhS/
nJVDiegbyFe9uPIHWpi3GSuXiVmct9W8K9uZset2Ose0YEtd8qyjNaGZWgXYNW4i
bzeJ+hYUNuMWfy8Rbnx0YUo5Tjm8VaX0LBk+7MyA9jX9Vx2VXBw1Jo2Eacl/6jRg
XwCNsF6LYvWTn7SoYd6Jop2csU5Ux5TGrRgN68oK+kk8ZTcG3okNYfQt6wff/IRe
5stSfXJxPfIC1Ie35f8gOUtDn/kCrsB839EQCTWOrRdVCYb3j1RvuR5eAA8DprNl
vBdxLxF+FBbM61/xNr4XIQ3jSPn4kFQ8zkJAl5Fq/7uqvgTsn0DyeZETP4imlx9t
M6JO95he+88LIANzH1hJ8pUD6D/vZvmL8/OH25+MaGqwMVRwy+DXArelHshv0oxa
Bbz/m3Kx3s/87vJr5kXeHo6zg+k9KQ8C73/s6f3sRNn8uNFCWVr3xoDgRPkJQMu3
ENWyCgcZWa5MphenS2gnuIh4Cra78w9V6qGRK1u8re1tQ/EUqgw8OeVeYa2cjFPR
ja8gN2z2sVrFeVTPxkZVIFF5xonaNEj82XjoRAlfEj3OmxERU3Oz02l+ePEC6wR7
6A3Td+PTZF+OgJvUK7EgVQUBYKq1Au4hILo+BAPWDfqVnYKpMJcPEZORUgUcFkjk
nF/R4u/jx6jkfd0VesNscyBE4YxLRtJLy5UE2VRlQfh0dJrVHBmLPoOKqvsZdUl9
56nXaWygP0AGY3rmMaIOU4INWLXU3qJKXxAtuuVh59wLThH7q6eRkyh9zbl6a71q
gGXQ2Uuxjm/TPM4GODPH6ic589WLCv8Bx063FcKWgfMB2j1ERI7jrKJ4XLUSSzYK
XS6ghgUHgMtokUdCX+ssyx1J/dHgtPsUCYZxhnNETl/mlzD/R7kZRNDT/xcQ19ww
udEqwjPS9VaALd8ey9Z5TbwV37z6SS86SrkarGxuncyP96UkyI15PYv1xsLJlgZQ
zipJYNK8LJe0DOsKNZ5IoyR4XaU8sosl+sJqAhr9b9cy/eXkXQlozyvAGZQuKNQm
eBI4rYOoed/QvckQSwHIPWMexAEJLa002c/E+UOtYu0PIWRchfp2tITGC3IsmTTt
A+Mk8GVnzdkvAj35NvetAjgI8vaL5rUNl4oy4Kj9viooVn5Lpa3wgyUqRvti6x+s
ooDW+n7zZGoc+jAsDFMjOajR+5Rt4uqmd9SnL3fDaYI55WgRr+dwftyB6mwWdqiY
TbfuvYUFdludm6JyWbEBe9qCNF/cMht4HHwvOyOwf6RPenBpt33vs2dOeaqIsyTS
cHlsaX09NisjmluiSoctH5NFVT1vfYdjGKaiQC8JUQHfSNy6csbEWGlVNMC3Bqc2
uriVVc8mSAMHLoDPSy0AVqDWL3AUfH59VCs4AsAkD5R1x8W6mkLaaOvEzc1BZbyO
VXImXe2qpAvWoVZWnnKsWnKE2j/EibrkppOtJZ3KEwgO+jHiMB3zhkz8NjdoXW81
cA2CXZkdbqRAaxcGzt3wGFaRPBPngSN1GV6RqRlrTLDq7Y7WOyVtz8y6/TtyZ3EH
jiVaiAZrccfg/fuZIUjZkY5RHRBESiPxuh0eS/MK44IzNaLHqlR42L7jk8cgtTMF
L4j4XoMBcMKN+8Hh1VgC7vXQxRHWjoQFzIbzyj8q4haVy+PdOaVMRCEQ/woJ24Ur
lxUxQfnmk9HzX3U9kPut/tCHUfCtmvoRT23M9Yz+DfPfv/ulD+Yj6XqN95i1ldHS
9lMeD1Sbk291tLPEtqovTvLI7i/UeB+7I/BLPPuzlRb+/M1IyXb0oYQAaGsfqnd+
CMt2cf3/sMwthXPustdD5Nd1JY1aSQUf0B+cLRgAtmEnEwpyKsA2JuHvu/qNLdj1
feKxY/rfbNzFZd26rvlZOZoe0LV7XzFTJWP6uTz9WVB/6u48bDZXNGutBHv6y6hG
itfnRFPa7dJJvTnYKLbvvDmcrRceiecE0JS+e5/5NjJWwe6qkNX5aThGS67g6UBa
u9CAY09JO48YTw/jgtPmqFhqjk+XPsLU2WeJeg+oiUPhVafdqtvHBeJPy3asDdBK
BSZiQgLzoEAX3Jx6ZpUlxS3RNnrg1blsE58iJ5OmdD0t+5AKp7aYGSFBOfCDWSq0
TUStDgs7zSIcTZsSl6T6FFTkblVfaX1qr/55sv3/RvrcUmpclNZM6HqQ+azE9IqD
vbm7YwvjMDYsC1w5agLCDd0OLxHfyly8bFIGHcZVDrkkAdnmhb3npd2m/3gWYfPl
+rAwfFagaR0PyPFQpXWpv/UtgJZXIPS36oRUOLEDEfD6Svjj+4ZAdJAJ3vsUkTkU
VtKsaoq7K4ySLOm4MXQyHddmTFnjzlEaTRLm/YGcMW8l9760eyTyDCXLVqVeQtcY
UeoY2R2GDcj3Vp5DAwPugYEhpTYBOdYjvyf0H5Nto9lAo1TQZPVArBf5zAZ07lV4
tc/h4mYEcu9M9/SQ8S4pW45jRAYg6TDupskmjadObjM4FKkzI9Q27SGKZNvKNGQ6
EgygqPpxCew2LyTHD01VN67BYmdot5wHGDTlNGH1MTHdXb5xlLIc8w49OX64mri1
pz1r0JROATNbJ1jG2nCGv6HFQXZJDhhrNiVFHEOr5WBUCXMfFEyovx0X4PuZ1utg
e/L517wLWVkrp9jJDyp0Sh9XUB0vf5teM98O3lXc4y8V27Zv2RUFh+uZw13LzaEk
aWL84a/vlQghd2S997Nw03ALbLfGDWOqsY+elV1tY0Np3tUKiIJCqNjEb3ODCIII
3hjhU6ZXm0Hd48PsuI3GqS8hZlvl2vj3xoaQUIbnp+43zuQtl7jK1ZZ4P4+pPvmd
QmMTwIcj2fQKl31+V+PJ1XIzF7EWQ3MLaRV64y8dAavDdBYDzmClxyGz7Vua8BH0
+ALUSzJoQzg3SbVBtFnjpU6W6NoMvAMA4emsmPnFQGGW2S8OWlRICiondi5emCpw
0Pj0KCx/pp4c/BJ1M1NnnP+LNeG1xsK8Rj1BzY5Euy4H37w5TYRKgUqpvuX3CZi4
BfQiuhxIlxYcrNLYIxLWqncBfbIPp0WlLWkV9CTN2Od7mW9UOGYn2rwoHgeT5Z2k
6IRFrduqGw3N5c3wd6141P2H2JMdNgP4zxnL8Sj2fYkEdJz75hvP1+p9ziGN9VjO
SpjZJIrIZlGpGpy9zjhzsZpyAUHVuHuNA00R6RorCAvJ/pHNHNJLNzCMF1dFwvME
ARfvl4FKtPon1ubaFz28dN2frzoVFMhCLunzig2HYUZVl8i3Cp88IQ/TMc4j+9Cz
rttmLLJeXwzgWJTrBDnbVYWqDwn/Aazm5/GAXgaQ55IolWGYXkmdZHfmy3I+nPY4
D6pRhuGM1j4Tl9GkwkFYrxDV0JzznW8uLCyZHm2uShsYJzd/tY8GS8Q2qaXBzIAA
onrGBz8lDWMVSmahvDGbKKrajwJtc5p/6nGCsa7vgBbSi1kOvc9iHna0nfaMYXun
cKnH9WkSVroXC74NbQgQvqjK21PKQGPp1Iy2q7etYKPWrpbbXfeXYZKdzFcvBLzh
rcuIan4phUSpig27ye5HUVn/GVqkEqKn9pMeoGgsR3d7dbh0cLrMheXInlj5Lopi
4Me9i6QKlkb7B1xWTMRhRDRWoEAVAsFQUyuddDdQWELPJvicKcXKtCYVouSuVkN5
vrE3iwp1bjJlqWDGZM9QNdwKoK1dVfPjOJZgE3Ba956okn4VFrWRoI+Sah99EJUc
J7ZIkEbTgc53i03afeq3zTosrlRCBj6FxDDCQ2Ikt7pVibIMs2rtCFrTV2nPfqbZ
+BPYOhugfJkHSoJQK5Nr2Ec42SqLxFPYtYCJolFAiXN9ksNuV/JK5QHbXPdM2iRv
zAq+kVguspi5wFt1eW0diTt7yXy2MNb+owcke811hR47m/sO6g/nR+FpMILvFb2B
LphjRIFUecvteW5FDeJujfq0Zftb3UfLqbY7GbID8iEDBVxSZyOy0X0tJQrkANZt
wfeTqwxrwrty7VxLE/0BTSKxC6KSIVdD2aZOM66CJ67Cw+5ETeW683WtXbZHbOqd
hV3BYFBJtnXczptvUfunV/YjqcdFPROPl3nsEYvS9ICUJVFg/r2jxNjd6KE5jSe4
giqUq0srRA3FjFntMhUtjFCyQBrBffTS+bEETGq6mlEycfN2ZkXLEyn0IoR+ltgX
snZdKMDUarBH4Y22XhvQiFAgp/4haiK9wcfv4e/V+yaCqH1/OEr7bjxZFEggF0xY
zlQ/VTkfa/DgWp5nohbqfSlvi2Puz+OXCOO9/lZzk2mngt/WKL2+DdLzQ8N1fY2I
Efi2IkuHbc1LeLsH6tVhDY1+KbhhYTvc0LUq4cOp9o+zpXKb1fGTT/jr8oypextc
Kft5QaH8LgtnTkhlQvYK32RoES8xXjfRfUv9ZFte4pTQ2JiJiUAxmooKpJokZre6
VTnPMn6cB40T9VUUQyvGnmRtWVLtk2CmxsONa7xM9W/2nMKENixhZgZN+hGgLEz4
qeaTX7u/BGvIFqcRCni82q0uQGjK+bNJOciyv3YupDWmVwjcwKykoK8RXFthUalf
HKBOqmAf0Uf7Qy2T5VR2YaMz1vOQxUO0Yx/cI4LAAPsG+zFn66+njssgaIYQ/TaZ
vanstEfXoHrrm9roBUh6+8owpw0kpEoHg5Kyz6h7veZd8T23Hp3iMPOMNwDlOBhr
xi1G0xVP6yuEXP+X5iUmFF/3dIu06zlz8bvz8z/SsqB4TKgFO9MRFWE4SDxeNxku
0fyEBSzVqkOMtOnDf/VQKIY6mFg0XqFr9wcHE2GRgIf3+ZIDkQSIEm1krfl1uWz4
KUAlg0l9v1sOX3FHvcIDpoYL7mnZm7fHwHjAq0+ExWqrJHYak+PQMVG44IHaqROO
ue2xvgG0zel59jzHToT3VYpaHn0U3+mziduHpPhJPu8kBalDX3fJeexttQ3TJhcY
3q8PNRn3cAfbDoeWDfjRxTyk0NZRaVfwwMPy7CKRbMT1dp34C9z6IWr8YNIsxAns
Th3+a3VtkMY+la5mO9SChIQNuu8AoJKQNhZdSZfzBDvv5nF5Jdv7/dWvdad9jkKV
a4I9xGzoVU4A9BiXvKLYNBeNvl1WwKcudST5MmLQWJMPvmiEPOImoW89teXRtzH6
aq17XjplqMm4am82HGzVsdiRiZWfEOVrkatX5geg6ts4PFS+z6Fwd56w9NlykiI1
buUmeHB8tyw+TIycr2vNtFvIlELvcxOVd5yC2YQCfEUcDj1TWAlDmNgMmhNER8bI
u91JUBebL+CZzMTDRvkbzSvwX97P9c5Nj+PRGn4xq2hZT4GWZV7uV5HIFYLnukq+
XTV/WQSOCesF7aY72J7Pg5Xx4YaOoncxFAYfYUkAwV765kKmmWcYKxIs+Qe4uwLO
QMpFUH3M5J5+zzBoWf1AXWRauHVjQ5wyqBeixDUxPht5q/k+NRUzcTxj3CyG48Z4
USTKGv1LW6iuJesdRJ01NwjtVcRZvbGtvVd5gQGcEA1NWaJ0IAl+4JM4DG3DhiDh
fwVUrNelbVnQCC+mWEFiFT4Fd7P3N9y5Y3F+jU3wFIaXMa15BWbHGVB0oxgkBaM2
K9fwqSCThBQrKu8baJO+/lh6AnlFu8v75Y77/59pYLlqvCBPiAUhk+e1621TJUBl
Yo/EV0BNNVv/30HDn/ZOjiz4nnSlUA9B7Hij2Y0+OJSxaPKf6ifiatd9xr6UjXoU
abvx4GavXthtSGCToinqxGdRA1cT/1aFfba8ZUT9CaQ3M+yjiA6KbyhosCxT5knV
lPeZY3lh1su5tT2O4pXtxq91XPlPLi0HFdQuH6z2/unysjnjPS5yC6T4XSgDXWQR
VzZICA+0liJvRIJdAHeIiphlDprMdApX/nVK5z7ODMFf+ZrS2tTavPcl+5q3mi1r
741WGABZZrX8OAn2ySme1w2YDKbzPrDB4Zsp7lmDkWlRAU5pWoUF6sFnOuXzu0Oz
1mOhs9izLBn9DIXwLyQM1B5eofRbryyAcAnUpgz5+t45Wy2OarCSQ2PoGTQblYoV
nH2hJFRF/PN923ldjxnSp8+KetaVOgLcjmDH/lhp92e5KrbsErPvhRbyf3WOyq66
H658EsSXNOuZ/vekx7x5+RvOTz4m873O9GHYtfjMGmYMkeGfe0tE4aCSkaMdPo7N
DlCV7cphECp0qT6mXcrVdYRwmaKdva4sIZ8Lh4m3O0z4zfzTYpLtt3FH08aHzzY4
6a/Aajfap1np2xp1TpHe7h776ELfBCr9i9diKwasHEHiGbwBHgVqG9ydrAA2RBfw
Xp50UtOdjB0RlJthUaNaGJazdJ7k+0o7rCD7eedMtwSxH/AfmqfHhgH0/Udda6tF
e5lAPlIRLZVKZvSl2D/R0RBNdZ8WCfm8Yk5D73HIc5m6TJX8InKLKfBD7l4zqWLi
tpXa/3KV8yotoJYJh+aUwOJlRY8hi03fxU3fLqhedE6DrDhUPqtbznETVjq7X5y+
Em8YlqN/9k4yHH/8CARbu6XANN3uezHOFqQ8SwQfEBKWxDws0dViqXYcvZRB78vF
5JHAPwaGK1RgxWDKxdOWPoWrDQf4p7zFaWl4+FkEtdt1zoXPbt73hSJE92mCOeD2
ACnPNnHLJwMApJmP2Zn28ljP9PtS3QjkNs3yT1oM33sWBcq7ag3EPfG8/sze7cUJ
b9n1rej2yMc5Tjyt8qRdmEJLvNDEqNr7zhv6Tq6smOeMGJtowhxhWbya2XjR+Z2H
5aeQgfqlTmsOPXrchoA7fnccj/05XZiyhibKcFQF8Oaq6jeKiQWBqYVGUBEpSn67
maeW6ed3FXFtNvLxp7rEZe5f65plPKOj3F4qnYVDj8jC63w/xBzb9np5AaVxTW7h
1WfkUF9vKXnBcG0lVorwlEEgMRwPVwJoCq5E6mVRRjDALh6emY5gwoKAtiWm8Kpb
R/k9lRObjCRv2LefX8JW+AobmeUHDfNOtc38QE8Vg6TFiDg5M2J1zMeyW3FAZdvJ
6QaYlkEeusjyf5oP5qUCKJVMfadfqGLyZplsvUb2HGDRxiqpD9ZDZEZN41EEzKLE
BmJIOfXm5Wa3vftvtzIEQ4d+xi00CdZp4mAygvGrSj5Lk3FP4fuIT/bn9INTyjSr
1toEp2ROsyYHBlUAoN/cLSOJggxo5l6/+YkRntJ/+7V90CtAe014sV3sOTv3mqWj
DBpK1WMA9I+xLViHr1Sl7q5f+AdW3wTcnoO/yHUlc7uWFCOHUYeE8afPpO6p6/vp
8wlPxmKim6u3S9M5O/tINFXzNEqblEOV/4Lkbl4k6ADO+BPXrPwHVwvIKaC5PQ3B
ZDeCtHfLqm4iV8C3cibuK6KvRmMinfooRLsj4kE4Fs/33dV/gAyp6TXj8uEIi8e/
Fn/jcw+mjG6NJCqX8Zb/zWKyOJ3EjN0QxBlwCRcfgt+namCA8R3Y/pnh9J+flc1D
eh5Nm1i3j+5K6gKN06vlN9YRhEb/dgm3vkIJezVEibLWy9RDKDPPiZy4LIo7UboW
lG+Pqb1lttLkLNxlpu7Je8REm9WO0N1TK/NB7708jgMQBW3y0X40ldUm5yZ4ycHQ
hkcSmOKwZXurjDXoTFr5ZmsqWOQCrTKeS5sABUP5TNyPuDptL3Guzp+6N2tMx5AR
SUwKomaI93NRj0WpFhE+T1ujdBO0BDQNq4iQOdJ4HswfkSOd1w5m8jUgXqVAaQaK
hQ1pVWuJkGuB9Uui0UPrHVzwoDtIdFR+ZJIJ5MUk5uFpIy6pWKQ02+Q0jD+Qz6FE
KYWNTV4KTaD34SGzTK3+sLvF0bpt6eDImiJKpip+S7WMtKi7ZYHkfxND8br4/xvx
pxZ/wRo256HBJbtIkmge00hv15LcxLbqfv5CMc2PBwqDG9MFnd5bELP4KvlvZ5MD
ZL+rrZL4MBTgjbdL8hdnk9uMJItp8TOUvocOXhnRZgBrvl7WtgVk4IAtrROP+RyR
8SpV/j786zK+BogB1Yd8IPTOcU+U2emxQU3WsYCTXZq/YUIEe1t/xGTKJWc9Mnsb
PnChBoXbCfReEH2HPFxVef1mSXUjzi//sy1hstvVx5XwK1VsmPOupdtJYIW20qDs
wX5k+OV0zyyk9V8Eny9xJxM7uufBGooyHW4GtCP2YVh136JNDE9zN+Wb2Z4qF2uQ
CrP5aQE0NfIPj5BxiZ0vgrRiCHpLig4lbK/oVIpQIMFAZxt+LGqqORYriIKaIFFE
jsJkGQOnCQ33bAXwrkF39OKgPzWGQnxSwN5MEeKKCrx8XE1VdHwgOFy/OsKqdWgl
aQyF8mkjhyXV7TMJnu4btnSmDFlBkmWGk+SN0Wpn3PsGGBKhtZ7tmyjH6b/IS2WQ
n24lj50JrCPmBlMjUa4EAx/++S3lh2Do+ZVBFmGGgMbOj+mV+ztCuhRqExrRVHwZ
fTzVuY/DlLV/OXGYqA74u/NKGC/OMdNpHPQedq6JZgZAlrUfqyphBzJEJ/nMaDug
+EdXbuH4JkPuqY9dUzO8PX6v8FsQJi4gKzHJA0kf12LZkVa1dkOWM8MkJ1+aAA8O
o3CwYbzJu00bax2vzBh2Sq49Z6xudO2qh71joTxzTq+elPCEP3S+L6xpJyTBbtnk
hHmOo0MDuUG4qN4D06GwkNuBRRdQH92/EpLaNRpWIw0CctM2ivbR2ApEhWEj07Eu
931Wk5L1Z+EA/RcfsneBSEUIbxYmOhLM20NcnfREzfupYZEy8311AsAi4Aq1xPx4
zoCa/v7+ToNmTsRpZGb+gmpCtvoP8h69KQVLaMqXPjz0BfosZYYpIg5BtPj1+x3B
hxpqcaqMHcGnGDXXtjCQ63mMfKLepYGaxw7HDAxFl8DBz6eaeFAqfgqapPIXTjY4
QkPN22rXAnRzEPKbYKJKpOL1aYbLS69waKRwvHCD2KvLaF6D5kn4CiY6+Itn/HWP
3k9NgTDWFmbtRIyaAuBtkvdc+ALQIdJCkV3qq8A8HijlJMV3s143kIRG2XwLpqc5
ehZ6FyuU/gX3nxHZ9+kXSbyracc4TPi1iGlqpVlArt3FZWKOgFkhaLqpXpbpSyRq
WMpNSqseP5zDd1B+trl3F2Tg/Qb3W2SKYTkWxDehdqSirhqWNQRxQZ3FuxuX6c78
AIwFow/uUe/xxW05hniKb98zFSIo/RQMI0uVftBRKDwo4ATKkG7wheAD03Kwdfi9
vo0mgqcEcuwYPiemTtv3VU1acXK0T2NnezXT+xGJiZXwOZpP4J1A3i3DzKc4unNe
+Y7m4omuanMoSakmAoql/+qHzTWniwwMa9RJGmAahRfQE38lPqI7PTm7IVSE0E2K
lrtRPC4SY0RDBhcOpc+PNgWNLHwemYgAyW2fw1tZAUwxtx7dfJTkd+s/7bVlupRE
52n0igYRWx9jrur7fcS5RGtfDuWXrohj/Inj2kH7+rkDbPvBmcrXw+NfrbCnkpiM
Dz0kvYYx3TA+Ad/JixYVuazN9+6+DEG7Fo8ll4Jfa9Wr/+G3ykjF1JgTYapgRWbv
80aBoPHrbDs2HyRFdCLyZjjJCpnsU/WDGlK+fJ3I87J9paOedqtqzmkZHK7WB3ii
mk26O5dzT1vXv6cMZ3TZwi2tghHJm8rEpJ8sr25HhQWZp6JPFe4ahMPrTj2oe9l7
flbf8J4NbMgmJruguQ08ibVjdgCd+NFyY643Yzi12hPObA4rp/RmLB3bWwtxT8au
OwoZJ1zc6afooDPPtJPC/gpXGmJJqlemyI8YBKxTc6zm7F8TGMGBSFNWTZtz8fwj
Gn+3gugk882SVxrm6hcdKxULRjCi8zJI3oQ/Ag4NRHSfM1TtiTecPdfGwfpNT4Em
ywdSk3z+FUZq5O1md9Yo/zmHANFlGjNX1FwrJvey4KlpZ5oSRdYSOrJ51k2b0CXb
7pJnBYwI+mVfy1GneSvvqBKc8KmKWanClt6TOH1m/aTouQFtjFRftnsYgCjyqia6
K2cG6Pdlkmc9jTgwUSBI1dj2UPI38FMcN5UIiRg2NWcBLWTTfwNemYUvPozEdLKs
5lzg007KRc3qxFRVpnBYiewAjZL4Lz3i0D81lJC6TPuwER2MaFuez2FOloa+t5hB
zqajmZzEnV3WMPvShghTvBT0yMnI8BT7ty5APGrOYCrT+qi1dWT11SU5lTAL4ETC
tawnzjEitoE6lXCcnkhkDFxya8un5nbqxPsJTzMcHDXZZ/FqXA5ZmJDje5sU7G9u
2sdAoTXGuL5AMIXFGQ/RnP9xpYQmDQ3XCkwotM0GNKbY9Dq3wgIXqxozrNmWgedW
7A+QqYfZdmoQduqNSwq3XTwfxBFMBtuuoGzHrVoBh1M5vDAM9miYYew5yVlsCFyG
Mo0Da8p9Zec9p7U84aVJgCdYBb0IhQIuwXwCWVqur6eDRUfUbkvGEIX3dCs2vu9F
GZaGaIHjdQ1BAtzZqBwrofPS7USjXxzMYc3qiHlURY8rMu4zmapKJyiImzG7UWUW
YjhS5NmgwF+RQBRsi17yYkbsHoIa77U9r5ShtZiZI8odptZKY3CcNN1+ZWsZ/Qdb
WwPbehifwlVz10UviZjrwSiq6A0HgLt43HpERiISAGcEblqT6gB6KEKi3LyA5v14
qnEZViBgS2Va8BCy1uUbVDvofE0S3G+mNrJo5F142Kim4gmMeUKeZIW80O7yi5bn
vUycAzVP3+31dwuuWfHGP1DByRFxHedsAfIyKsS8dQipcUYih8Qs5bGL9uo6M1i/
ZGlG3nCkAoZ8ZXr7PrXUfC6YxIs2LIcLlMVguY7e28JtNqvWlsbv4imNOlK0uv9a
3/XUTLOpUu2rCEVsEFh30fVN5Pm0sQ2MpCoMk4QVL74WXRr6wVeIJtVe+4G1JQhK
CjDlFV1LNTEpM2oTJ2FXV7n8rKbtN9POsmYvXpZd6+ZQ/+JgPoBDJ6tnUpKMpWSK
09VdpRkCu0EyyfBMh4gxq+wAoBlU4XC4vDZrvaV3XUww5R393FTB8N/9lZve4ib8
axp1HHCQu8/27KYcED+ygNlbfOlus5b3pXseRjEKgec2+NxS7ld8APnY3x3mitXJ
XMeKFOF4+ZLyB32w5GIyzrivAAdz3tFfL4zAT2KupWkq0e+uVY2TOgYP7COofCzY
/gCdBrBFIlQZKyGSeLP8KFNjGqYoiUMtxTEY+svA2noJBaPLkc1siqOJiet7izGA
IFTHFuiL5yQu6IvGW6YvYiTYXlpJqnuwnK2+JLdVaKAvKUlaN9lKdO/Vh6V2UcZl
6lM9wuwU29LQTGFznr5erfWU0HmtqAZ3Rm3FvvLAghSRlibstpoJydT5s+wpnNx2
rI68PfWO8BAnRQGK+ky2f7TsxhwnoBDwxg89PNg4N9cjcaqmtFluwJepoLkg3TFc
rHfzzv+N9bNpNaYoeDooauBtIYMnFVfmBP2w2xUl4mlhtDUXz9TCmkIdIFCfyqYe
kodnWLd0p8sLIJIOs0lkDVIRneCPAfhYvzE/+N0qUn4CiiLYoPzq7E0o3dq5Mjc8
300x2WprHR4X3/WqyHu4pcyRSRB/eDRrUI+RbQUIcYdN0i/kTkwrwn1hI2XBCdMJ
rT7lJN/frdd8j93aP67o9WN2lIkQ9lQVdWwolevAzxdb2T1pDOcn4Uo89PD7yLbK
e81SbHARARlrn2+VE8RIdvqI1TG7jQnRYdKEc+AQ7WwHVyZIDaLS0WBicQkR6mYR
wlREP04HS2zyKFCX7d4nx5WPJudfXcsYolqgEoA77aREhYNaophp5TCU6St66pXW
iSJKhd/0P19gCTwgNJ97IT7t28BdDsgaqtW882OA284ftW6GGtl1GiwyO2Md7WQg
mu4PHc7Zh7uOYJzzrVSa3Xg5pBy9jt/xp8W56BmlRlBf+zbqU10IyLsDhvUIOedZ
ld13enoNVu0LfFiHIBK62fRFCNMCzQf6eJmdNuMDeYfJ6MatHewT0nMRSYoKblR1
CB8kTVQ/52MLyLQHfKUx8jCIfPggWpfp2lSTwFYEecVARpgAJPGfnu1ZEpxLHlK4
+sISnviPsb1A31Z8VTDV2xSHfPMoYE0QLqZCKEk8wMCcqNohIgr7ayxFRVBUPeOi
sgdt/ItlJiTA7aAf0SogHDV2hkcQAlOqVGEZR1JAAgX2Lsw5rfUT0+zu27/N23MW
Gqn9n/AM2OCNX/RxwGrHH0IwcachCOq3aXHHAsfbyJEU0ZA3ta7uDBl7b/J2wB6+
me9T11NKB9srXvkDOhJx9FGmVZ/0MyRXLHPQbi1s6m6gtkoWEI6qWtMUPESbDmqD
tpArx1TWzmQv4vZqisGYC+v7KHjT0w5fan+F3vvf7BswsnbF6egnLc5Jl49R/cik
n/OF9Zr7J7yd/CgzgDGl2mDJVAfhoTnPh6RkXIw85zVFLjx6REmtQ3GugYV1EzmO
nXUWusSaG8cU/0+RbFIuK4hDxuJak18jnN7GL9WbYiSE/xMOByBGSfntx5ST/oIA
oXe9J2azSZIQXFB9oPbZ8xxKQ9Fdy4XHvabzH+I6yk8RE8MRV6tApoqzu86V/Bed
+8FVojq+ke37zU6TS9plr4Z/0uVcPFMjT3r9bN0xxDXgLWE52DYYk7uT9SmoNJN8
aF8Kx4RjN2R6BaZG4QNxmxWLHRZBcp4tJFZB3OYCs+2xj2edEisdS8oSs4QjN+5p
wYD8zsxrU6BF4GJNwgg/AKWXzn+mC3zNPa7AxP8y1idHqHmFUCobW/li+XMhIno1
I8lMevEGfFxx45FzdLWnJ6CbutF4XAjeY7CbtvJY9DysozWGBRpw6wkPZ+XPb2tw
oloZvRb3ofhn9Rj8lGnuX7OWe18Y115nTnmSzhyBsSWqQwVl5dVs88XGjk40XbC+
+M/0IR3YNU18nfaMA0n+RgCWSDXfcIBKwAMNOk6HsMMOIjOhGa+bLD2YQIgWCIh6
aphQBxWksmFMGmG9TQG4qwyXl9/OraRnNWDxXhFCmR/JjiH1qDirsCh72tphkOOR
SK3ezOR4xDYMI8GXdStvPRGAWIuOseKo27pJu2xf+SreJX28j8xAPGxc9xQpk85i
Tny0edh7SfBxpVZNctrcrHQIqlXQj54ciQiXcIUPlFyaO40Gc+o+Pu/y9VidvSyt
xrS5RzFQIjm/d8sX2xGKehPB6ZQsnVrkYSht0GPXZaWj67ggTtvmY/MV8cr39cDb
B4IAsx0gDFt0kUak48EcGIRqHbf3NCGeElFYbCUTy/h6noPbzU5iE5wm+NXLFXa7
rWWmERElE+ItqTVzFUAeavuYI9uMa+S/nf/HVLAsksNZElZ2Wqnyoka1FAQodq9a
mTPRa5Xvc1cDxvLdB9289ZGyBhu65uskt2P80Llf7l+I6dNtTFeFBJgRPDW3EHji
BMALWbTReyhB4L4YIiie2hAOHboqdnOl/NdOmKhnALwCoGB8YJZ5GaEiATIA8xVO
dc5ZHQ1LB3VK3B2qSkuIeuiA9pJ0b1RGH8b4tr5omoBHjufV2JMsvtYsv+TLXAQi
hk+XHPQ+w4gfiN1Ux7rmQb/4wrp/o4WjPfxYJXQryemkwh/Oi2TcLksKKR0+DOS9
+HNSn7/qAyP0G/sGSrJ45bwY9ze4Imbl6licwFVt52TUzEMEIT8GegF1WvAW0ae/
fcZOnnadEi1nJ/vj2lDRq2VU8K4pTpPYUufar+xw7V6Xzs1UuojRuvDBUftnJqcs
8SxBq2T8+2yCBdbdUpKCDzUZzGx0WwUo1YBVmbPlgzX8JxTR9OkrzVMuFXUZAN0T
XOSYloOAY+4LxX7BA9rg2B8FPp6LI3+0bB3mnHU4Vj+jqbWeeWn2Z6YQ/R6trrnI
QgvWiZE7rwcx/26eA4CmjxR+yBVjEQZ1PZ66VwVVUSpS119MVKV3otZfJMHjpJA4
NPnKJHGaKb8r7FZGXTaWvOto6WkhC5G39YNeaym0z3673VJibYdDo789VbSfjHN5
9eEpwQ15dvGg0UNPKVvnvV3tuqIri4VnqcfPU45d71of+MxNJiyyBENFLD27jsOh
DAAGPqTGA9nl0KYj4A9hjeJqKxkD3TYNxp/nn87gwm8LgaaoDPIOq6MGCP9dhts4
6+GUtj4xYjKq88z+eWecj5HtP8l0pcgNNTHhh1Yy3yELH0Q7cR/F2FOkrPP7RvH5
k9TRLlYtV9geEWmecn8VgctGoJequi2Pl2TH2rpjuHSJ5mGV2fHRV2hrbWaO4bkK
ShA5qSAsx9cvkJwO6JdvlI1S8K3hpWl6Hs+WGaaazLN7T04c6fbHpgDcilhtIpFP
o4UmxrF3ls7S3A99Pb/7Sc/4CX1+0fUXvZwSiSvhMSREVKgyvH4INnoZtXnD5x2Y
jgoC40BKr2zXzlxk+wp2z3+QhPyA+ERgylfzhK8KuFn1gywJ3AVWf+Bgb9ZOXVwU
9YyAAzjhaQtMPhfLODxC/xRpewM9khiCQXq4/qPk+yQ1JovgdlfEbvN1GVHWFkXn
UsR67PmJiJ6UU7y7EZXLPPvg+Ly7lPPCcKE/NgUgAc4yAG0/qifC4lkKIHIwiqqv
zu4ozB7DJGUr5StjnkmGFLaXEFn/aIgrNgLoOB2OskT2LnBwVwN5ziIXnfkgdJA2
53SVtFayS32GwKWxDGbZP8lEdMQd7Dky4JTeRD5vcm2QQ/bNuqeXX5MqptdZNkz2
2Usx/6DNqeM+UUFZpnBPfPIm9PzzMZ9RbJ6nxd7iRy6QkP3bWodqLWg8We6NCyVg
X7BG/tftuRO1F8Jo6fVLTyqsHSZzsQa3G9ZHonFfjnQpfEwr97/Gk+KyaCeQppoS
eWPY2xWEJby/NtR+eSu9OJHYimmugKw3EIBqurE20Zcbc3JZ9WY20zZFJDcXn4K2
IYkHQlZThSIPD5LCWOvtrYszJxoBtQsKAy07HAXBbgGPtWWwy3Jf2iMcLpw6c/Nw
g/8w8p0FG1OdGMKuc9FLEuqd7UHxCf6eplHQGJC4TJPlDgESseyFDMqh50mBPy4u
Nfzu94IspZtJFzG3se/l3dF048vrXGI0y3rVNPqEF0QcpnUxP0EWePEQmhNhy3rp
SJLb7deig0KnRn3y1YwK7CIfX6ptvgNtzR0VyefTKxTmZS4bJ5scxQdyrpbg9clc
vYZGXS7cU9n6Tnoi8i91O6MpIyM7ABHi0aEGTHOJDjJIZKlABZM2Q2B46fgimg2w
v6RFBnU75VTNSyxWPD0ebu430Spr2+X/xgTJbR1ZntE193knipOhWEFrNuqsO4+R
t45lrcNqqbldeRlbf910PfpWWQL2KR01GsYDR5lt2SGevPxH+8P8FWYNBhs+KYyy
juTnkoNMQLe+yYU9J5P05GiFx5eoOCLqV+BvSeNFSDm2smsfYo2jFtj5EiTdKQY8
ybjcTG6Oxt5qzMSXxUwQqz3amenhSg22KeJLAR9dxk5se36Tuo9j0/sOk1flAvhC
SkP5acj6NIEnno1jcVj7r9KrV8MvBhPqijP+oiTYwMQSuUMDMC/8v4G1BDzlywbh
t6NBqN5F9X6Y1zZK2tHnaq4qH3KXrXv4cdpGK8S3vOd51gKJfFWsQsdoumO7ksBv
rkwlwtfxui5UkqTEC5/ZkMRgM4UoNhCFNzdvC+WHtLyGLzHInyC3cXTNM7SP3nEw
Js1DmT30QJ5+QZ7DFYGorY8i3OgvZxly1p9tysY3rBrztU8JPT/Ge8BQ/e0fDYS9
6zPhw7ddJqMLFLLkX4rgCxkEBlqwrQz4VPP7m4SwBPQi0NO3zIBDXmGrZUbe9pAx
GYIEcnVY37JwlKlbdAjuTnbqM6EDtlUsTKum/XAAuimThg2XQdB4vQazXuNaYWRw
QofSxSmelNxvD4Gjvc+fmnITZO9CffAx9+VHy5En8FVBCRkPmYntXOoJqsEuHAmN
/DdGFIGk/NMadySAHT5gtInt+T4ybXtqwPuCsePV938ehO5kcnFZkiJLQiEz0RrP
18ZlB00JZkOIdZHnrZ67S9DHoI1pPC0VLrtjCkRQa31Wv0c1lAcZUYJbsp4917h/
RjTpCvuNUyhtqyA39DlMFQOMHKSSRBUL40OItCI6wu0tLtdm2j6Rkq2nMA+U5PQT
VjzBrpiOHFzFDZikvugSEpBOloI/JadTLF+2c+ZFiplvumicFm3AxRKhU7nPuAYI
PTsTA2UFhJLpu+v4XN/m+W8R12Ffphl9kX5pvryX/GfpBzTue2YQu/N3Bt+kS5eo
SCQLvf4XK0mrYJvJv5gVYEF9vUnearRSnkruHLTB2LJH98RHYd4HGhRnIJU/9MUr
fGK7QwjID9W5eKVIKLGEqt8x32SRP/nvUXkPn+jmXiJPJ2/yhcemC4fYaAECLvzS
UIzKEYgJW4x5lG+YbNNuMYPJazh9vqjULUXYXonl20czFaYL8klzcMEasqAzEYWl
Z9b1TybhKl8I5NcqBTzWv2UCc+iaKu0d6F+0ZDItmbWV6v5Re6zYfU+v+rDFRdIT
OV6BbSe7jypqi5dTGMCZbePAhWjPHRVl+ZiiiAImdRhH57cCozaPf+Y++arIwXiA
jKznC9q93jMEegz/sRI4Qbfuy1/pEzE5lnJsw+RTc1wQXIszqurvIiLTYqAvVn+F
3je+IpT4YaAg2z9wpze0qW0Vz7fbJ8LfS0fO/SKAzmP1JpxekL+Dp3YXzEK4kMxQ
htmfA8/cNkNxm5swbjAQWdEsdbc73lbv33NS4hdP+vThhS9xv9oGpgdteL3fZ270
wYf+f7bUpRPBBW+eK3USzTpUoACkvZG5Ets70p5cvYbNkG5lO0JYRgQxvByMpWNv
23NoLg3zDJJTAqtkt25vQ5cm2yJuGhkBcIylJQRahmbrgpC8KZU5emr9P5XrD15R
2Kwk2lPNQkCAejcE6ik1BNwfwDOMtkkH2e8vN59W48j/w4TSJxgknF5mzDIblQ3i
3K1kiU1/v7wXMH1yFp3uKY3gSQ0MJMjr/w0Nh4nWd5ctyqki9Zq45aQgfcV8AIWh
1eOGF4HSn2n73EXOEk1kuFP4QLZadpH6RKNn3cuneNxrVLRGMUoLzF1C74GmhygV
sAeqeQdECUWwh4Lx9Ku//w6FIa8XW9tPGZc0irvFNNGb/AuJpRJZN97QEA1ntdfM
+v7hrz7epaW+u3nhCevq13j+feywn8cDQhQEhIJVgcTI/LXGSElY4+L5YO4MN1Zk
ctyLbiXjKVAQNlTSSaabxSY4j2s0yHBFHno3zshXJpp+ByjeRD/aiQVeQfBin4Xp
TNJ7mtJauMPZj/WK8FnWg9v4njsajItsTdfru24/KQXoRoI5wEaCrcnHPm6SpDh4
u+ZAEHr7zoo3+/LvKrIja3p7e5+Uob28rb3Fg35J6aSNX5UVU9Tob6U3wySaWaRa
TFJF41Lbr5J3MnkZ0lni5JEXr5cF48g13W0Bxin+xXKJvg3NmCd76pyWNgbGKW3e
YjdA2OpMUEW1uBUD7RDXBMchjMXA2joUxbCV0XH5GNHuk54b+yqUh6GHEtZPJMh4
3EWxePE/z7fINF1n4TSzbXAabDAAFpZ0BXq4WKR0X714Ahx64aMxh1/rOAzByder
lUxTVqogedqbb2F5Cq2Jf72ul/7Xhzk1rw/2nJstNKA7TvqV/uP4MeqPOqvnN4hv
/rR43U+eaonpEjfW1sVc8+VIvjimgPYxtaUJg3wuC5bjvArqxYljukzcXJ+ZTCgQ
mNW8iLJEspWSLNpSXMnhqHZQ/yQbvrttkmC3H1dTUcl8qZ/AGBFfjHuW+82hvb94
ekQTO59asuT859TK+/0y4iQkUJGugI9/Xy/v6hLzgHo+K+rcL+wWG//aKBimugwR
cyJV47qqoj+NnbBbUkcfyjarr4QHapAUPygKrbKGtwTIp6zoiKUudOxIAE/PI3Gj
1qKqph/sTJYANg1ULDnBK9Vg9QewJuuiwIqQI5CVkHKfSc5IqD/WwAm4XTMU4ngX
U3UBu2yGOzAHwFU/cgjww7xrh/8+qqDicHfTF3KmTsvtcXvXSW/XIB2yQ9QkvD2O
yowx1k7Ix1/PUEx23mk7N7gUnt4J+wTfNYOjBkSuuvY1xBjq+0x9K47U7ZRAlYka
IAG2sOFxdIdC016DwBuuC2o4y23eR5KPJAoQX6WYNMwv0bgZzqw1dUQn9jYpBG5N
SqsQCplB/4iK97hEDwLy+ydcvC8oLnExAL7ju5to8+f/CeqnVcaILVkvE2duyANi
v+mhrA++lj2WOR8Dp3mzZRMPki613i7FwRUtPzfYf7GInv7CwMziQ28zS6alHFZm
TZvw5/i5j2YRZRqevt7K/YXnCNKzVoEdvnr2H1MsDywVeFS0VC1Rhtyze77M0+vM
GkxB5Bk4nr3DACmwh1hKTd3BeTUUnT4koGfJKnp8Wuzw1DGrRCdaUyqtQdA9i3tt
tsBVUOcZuUmFJ+CeWrzsz33jzTcSysBCJ2YRhb7YSav0H/grmVpKkygCx7/f6MVH
8cAeqKkPup9xiAdFejjc3KiFr3k16FRFQcWXA3ReiUTmOdjBoyhnIohJdo6cqojD
FFnqAvSvqqCKQmbfjP8W9rX2/ygqXus+TI7z8Mea0AdTwQP9D7IieUjrhelLEaFD
/oDjVyid9nGqyeb1CdoUsrzfquEgxk6lCkQRsPYk1sq2By/ARgzA2SCexJxXv8vc
flixZHGJrWZxVcKcDG/SFSOj9bIW0FxlqNgur3JFXm1rWHYvdopI4MtamlxyzKYG
dZPuXNHEVK8e4FBMl4Qqj80iclLUSkLO8j2iaLa5UhycVLauh1jgxJw1dHBNWSX+
/lljV6diRsfSNadm0pTyp0/bb62XpuziJhZ06FmNOBgtCdRSUA5ft5dpU7GTmAf1
VdtUCIoSNMK0HxvmPaZ0FMSTvdT2jrRt2tjsaOJO+DndeszFZt0VrczyuKOPJStp
yKL66uxIqMrwj5Jj8BrbqFankm4bSu2ysG4CE7UhIwbGJKDUZMQPTfX1HRwd5NuJ
sf3vgph0W9//Kv61yBXxTgGHzuB39hxiPw6OoBxF1blvYG1mG0yv4cWrKq7sBceo
khplDGXJT2KElI3vjsXYlHp8hmzsWhbRrXycN0g40l9QBX7O4OBWdQXKup2wlYbg
G1EIjNF805AkM2KyR3lb5pcHwFtvQXVFWxcKrekKdFyEdyR8/xbLjNSWMP8TJDfE
DbnSwELuwQC3L5bhkOVC6ABc5EQLXxiWmp0HrCSCqCskrvUy9VAdo9wj3T8TtRDH
HLMvGKxFhfJEp04/O8prMM9ecJJ7QJ5/y3wK+n4KcT/I42k/9J3bQpckMjFQcwEu
wXXvy7omEV8wTpctR7KHYvtvQNMkQKn/9bFZ8JazEjcKHJRqO9UtqdUusURpm8f/
QiDnxSK4UFceOvpMEdbnTkzcCHVS2tglJZbgFFD6P8bpz14XkDfqGjIwClaS4nGW
eS9bFj7GwWmfhto55AeExk01RFx7+TVgI1s6a7hVoi+aUvzL7MqcN/tTkLvga3vn
LHbg6MRxK51JC1UnfQmorCQEb4S5lfcDGI6QW3oiPC4jCtcy1Fos08Wa9Q8JEVjo
XceQ/1XrPmDAFDJboXZQLowziwS6aAjQIzHR8gZ+R+3IwSsSbNVt+M4IzOAMuMbd
MNDRif8FNBS05pPEckjL6bI/RCpcC57xhWJAYAUN/u8UZUyN2KxsVpEccxqLBfW6
wP695e5iuaNOknsb1wmt1foMTHoPWoZYNDM17v+I3y9YXbilGZg9CRy5J7FDkxDw
83s0W+ZiEi+Ti6ZYpR328Nz+Qh5s+9sEaCynPp/Xcev4or4s3xSjpm2P4gpcMi21
AfHUbpBXxBokjak/u/YiAgyEStxAZXBZL9IVSqm2Apdb2xNtRX6oQ0zj25icRo85
WgKBTtznInayEQh/OBOZrsJ/1MYAnRw9lo5NvQMceY1lO4NEQJlzLJfHQ3hYzHzi
SxsLlZbpvCk9463IBrRYuyo9Mvd86JwZeActsNHq/Jc0opIshwzUIjrlOqPqTMzL
gM5DjZc1s0cCOIjZXrkrLt/j1OAoQFurVSHpe6zU9B98tRE+H/EhWC0ZP5mKCz+l
BuHIiLABCxPrh52t/8p+tyNK659JvEEvZRyA7x0CHG3uHJHNd/iYQMtS7MHKz7jg
jvRYcZOOC6CDjtaa6ausJfS/nbbza1H+ODN01oSXcngk03JO5MLa+ye7m3vy1jPo
OlcqlzmpTwLL1OZ0h/4TY28t7Fr9/CqXZxrbXd2mTvDuCjaERWmMssgyVf69sZO0
81joGutAhKtNVVYZGKxuYzrGGuseCPz6E9sR0lYm2KCbnR18KdxoBGvQbgz1E05W
ltPNA37ymZ9tq/JwcFNdX1yXCvarv616iq0NbStjissDvbvSPTtJSS31JHNgaxmd
K/Zw1SWbxVfAiyFeJSvT0YuV5D7X8xvzNer4z7j4jwQuNJFeYO5gH9KC8oWIaVv1
v9O/rCs/eEFTsxci14WSixaljgmoOwKDaoKFIjE7FalwaoLmoI8ALCZZY3pK09jQ
EtF7LISjxvNRWtz+M4sfm+1vYrRecexyBKSZaV/6OyGyuhzT02egkj6C2z9cZFjQ
ZZU0e+ktqarDlTuikj3cj2G7b3vijtO1w6rxs/dDuhj9NwmR/TqQLZvKQjoN/JMh
ep4785+sL4SZYYkrglZmYjymG8W2Obfo99Jz9pW19oWV7hDww0h7dwYALkm+hAzZ
gu4oYDFdKKoptleTpbCvY/XvgQzYbegDTAAPJlC7Wsnv4zppwIRFZQtEv5vnno+m
lZ8ZBSfQyPLT+w0Wp2sAOwJzXl5+3lHyYfm+Ew+9PeCsOwb0vzmfiA31VSzFgdy6
+d8Qd7XaSGmbc1cYNNGAVjApEia8JXyomnFcq1vuB6Ej6DFkNq+Jl3u7rlEZSg6B
5suDMbB3PG+CHHMPVke4NnDX4D4Chdf73yI2ILd74eygwxVb3tUcFB8Is6CuwyHD
5LLYwlTS2UjyHPTtqBMNKCbIax1JzNqQudnzM1AVILc7iS7QUazKXbvGFieDMy2p
zy3dogmQTBgHeGJMLrrg9mO/cGoADyrglSRw7ZLjX9iGcDQLZ1AmNJdY58tJ1bQQ
bJfrrfdImb7IdfTQ3a/JmNDaO2tDy370uX28RVu0i2o4QM9CTbgsteT2QDp/iPPV
ubSj7XfukBoBQRTaVUiJnavqcl49ehKyY6oYmHluVFGbB+n926P9Las9h4xuNSjA
z27bRuBKE4hzmfYf7Np9ZNms4fGBWaLLIcOcUIOa1Ny5Q/t2iP9HGMJBMIdLulWl
Y0KJgu+CTAPjFM3lBKSPM2UBKPAumuc8K7fmPdAEx1ALk+0hHYAWtfe1Ymi0oxUt
l79lZPdqaNyn0AgUzNHYvTqFFRt6Z6XVttSVKHM8RzoSWx1A2vDMbUV6XItQXcuh
37lLo0vyNrPYq36u3BnEuZIRSWouM3CU7tzeFN+WeWQp2LrFnlCgVTVMhpKgBtVc
pIDZ1vv1Tx8JqbIsm+jrY8iBMEKojkx9ChC7QTEK9/IkiqBAJrODv9zdRqkc+gWH
aDnHPKmcSHs1NsxIAmYlAQKHHxDgpvELOc3VDP88FcMXh9PzhS5XH6rM67xW9ZIS
9uuw61uWx6I2JxRog+Loym9cuab+fRJg5dFsHRfzdhe1MkEx/GCs6lny1XnjHKEN
kTiS37M/GzaNFvAXR9Q8R67kI3Q87MH7PYDtu8k65fCe0gYgFEd4RiPvzl01wJNG
pKTUQ3zBUoxlggIRF+0pqdUQ31lpaTz6HVTnyT1qG269QdCVGpPimgKoQGIbGzeT
P83QQV8bO3IK+PWrV5wS1rVHdunF5zM7uNcBbU+6+0p1Co+6Z4noNEzaUBqDHB5W
1A/JeWuJOmGs50rnrqlBKPELxHAxkR/v0almWNKQ006KRE2zgjxJxMGkOwzzKllZ
aB0r8kjwPTfAdYAu9glghk3ebv4dRkzw8JNA307VjTtjtpfRpUY/iOscIi8as131
ZfebksvMOqvGA1hlTGNXVYJ7VRW57yjb/RPkJg3h5V4pMdflRM2x0ocQn/5ODNUd
wDkvg/bBiestQYaJv266tb1bK90qZIIOMnj4bQaAyrIhIUXC4qY0Q4tpRqf65bZ6
YulI+cUN4eAvibEow+4rQ9hY0jXRmince2Fil03cDtKPYfqzeCxKzqXHRn4ht486
O5yqhDpVJ+PA70kgpkIv9f38rNjFI6/VBkpCoNQ8cD40HdX6sakun+jpzslQmb+U
5Sx6NuXm195Lc/rZvpKJAg3hWYzvhPLnf+p8NsM9GD7s0OwDCtGXX/S5zSDDMYgK
99noNCPIkd5+AjlGZbN9EZTZbi7E1JX0siAJZBVPwGvC3k2BNNlV5ENW1+6OOv3H
RkIVfe9dIjc5a9N7s9TyXLKSTT/EsRpXy1c9P0LDep3DgHeQDH1uALXLIAs/tHog
uPKc98JgqdkDug1h0EfRH97bqZV/KGCTRpHdZJW280B6JAp6PQ90dGyFyFEHpOY3
TFUUdloEAMYpZCVQiAfBI/UuqYapivsi3PjOXvMCJV/LNqORiyPkH+vh5zyEtu2n
KXMdhWrJfg0+J0qjx3IxwqBPBKdil7r7Ug+CLgX+rfae9AedaA5kPJPqlDgpjnaN
2ltA77bgrOZK4eq8rrtKXNfUszkv/LfK8Mve6XYm3UNdeOdCf30RHO85dbaPHe1O
7GY8utLcoRVTM45K452OSmSHmHLn+8xMafBhfiTs+T5k0MzyIpGkmFibW9VSGwYn
4qsWEc6A3HE0xOjzB8s44jYpUIaMc87idn8vUYuwzSlt5q4079JhdUztf7PrLxxY
2JnjQND25WABcxB23iVppe2C7L4zr7/kzomkQaJ2s+0CbUTddpDx/DzOKl8d/EH/
jt9JeJZUiFWB3gGEOXqaFqyXRZx/vLxvy9CHaZcZuSOqBE4lT8UHNznUh/iwjWK2
2Fj8ftSil9CP/YcAHoPhm7xZa6Qhqpu/wHQlxzJOnNfSLB7RfVfzZNzsOHWOLbOA
d86NILCE8icvap1bGErWoYqFskatK2B0bguPmtDXeNrbaPmy+nFT+KfhGqzszdeQ
uw90h0E+t9q7IfEVanvCZELKEjm5SLutkoA9MnT5dHD/ddQHVIlhpARhqao895Xd
JWbE3QtedPNymaiMvRZX6XnGuh4CaOY7UWWSBh86CZjsIJXn9QwiH2rbCnaGtLD4
rOZz7NkGkZYbwoIxb3zj5Ar+JdYeStu/T9oBbuQKqhO+2spd59ii16tzoz315Vn3
Z/72/mc0cBDQBOZSQtgppBhFdue2R0c9xulBFxcJOSCwR6kJzl2Xc7lAosKJ9OMp
tIZDG0eMDGxY1fcmQKhHKDeeWSQuwa3LnNxsPHG1e/myk9gu8QrHKIwXx92NirKf
JvvkpF3EjWocVqJsoSulSk7hsESyVLtw8uT1cQm7iuTBCzuMsvA8sMsOeBHDrCs+
Kw2SzhqwODdF5jniGr9cSIBVHLBCt1RdM/5pIaaDW0Frqux9njVqkXQjBgHyq+zW
hIQi1YtoSN2F9gWeTKqUc5xp6SanMpw0/fdySkT+pc1fmVZt+nDQ2jMYCh3MNek9
0sG/3zFMcnrkTBlyYL3fXjxW9hGWYxQ60Rhpy/ms/2wPsVSzmtigdto6rBGFwFkm
5q+tV8j5krXTjuFBmVxXOK8RYhIpn24LrOs/b/V2VR9WlOw0NoUHOqQEMCeWKiiV
LVbW9IwC+/23pFpRPdu8O6fpqByxC9r5xii14dTARr1HbwnyjyWplKfYfPSC/VvN
5PvaROc/KceTu/JHK6rl0NvHyNfWuDlgjg98Qf9M2ZOdYFavyp493UvF1hscqv9E
hl7mq0HJWlktUrYq2X/abFUwJS/D37yWYFL8Y9SdRDX03IcefyIPSPjBUclU2PmX
wTjFqONy89xwd/EoAHJO4V1YPNfZ3+EryyHyYbzCB/gas+vWvhGoOAaTcyrS1R5j
sSfJKxKilcRuKaYLFZLz4aXjK00qJfV9dNG0DJVmtVmHtfXUecnZJvfAZ/OzYOX+
KJYSeaBuE4foQZFvJ3h7Vp6EhqIqqCEqJr/jzHMzTXKpqGgigDCD48WSqmE3hw8B
gC+5L1JawYpRISA9bnAm36Eq033wCriUUbtB1a/DajjqiaEUNuEvrcp0C263i1+x
MYobkMJMirJ6/N5AJwcb2okWoE1n+OJBLroSj8NC4wy+fofAreh+EuHxkpn3USPF
xICigQbtB6eNIuFWW4guW7AwN8UYvXJB7HKZf6giou37+zKXfsNYJ1w4fcMsz1jy
aRFm9zaKsOYnCZibxZHsEbVFgwFnx6YhDT+RiUfxFk/WHoVNlEsMCtll1Z2el6Hz
giP3TqpXsaQ8vB2no80EjSsMW/qNVB9dhZ8qb4MT5p7PnckVe6maQAKDEOklWheN
lbbubEEQ0/dIx2uSyLLRYDsHVlUeptbG6EpULlkB+t3a7ojntoC1EFnMoc71Ei/o
WmzH+zGrCequbko8wvIJy+iWJJl09GHAIuTdR0bSBl1tkcau9rT10jmBrEUAJ4EJ
OYS7e8m0oNVMPZFiVaxIVTC+uZJH59zMGltnxuoYw9UtqbOYHnlUFMOJ+5kfov7+
2vM5GluE7emjMfs8N1UAG8YoUb44PZ8lCEeAawBZnlS5sxHqQu7OsMkp0CaAUPq4
tYBaF7MwEJwm/YSys7O11dqXTH9qQk+DfHy8AjA6uIimufcUPqGm13wUAIGa/poh
SC+5y9H51r6bnpS75eTMGH13zXdz7V5S0NxXiFiyBg/xGR/iZ2qNTy3pdfwwO0zJ
hhp4Nt1GOvVTAoOIlHd39fL9rkzBE7sb/sBrcItLwEGgEdArAPKnGUdkdZ/Oynkh
Zsis4gX+AqQ+wc5iOQvyP3ryLvgWMoKhupS3lNYPDdOqmhnUxorGzjzEuxdj4EQk
fB+HrlLu2J5vtfm6Q5urcmBtbcNrU1rA+tLd67EKEc/at9T3TTJfMh4632B3OpKZ
P6bcmR74JNwYj0evNdewdOm2+kI0FD6EpkXhTGMLcHCQd/IgSVenWIKSGBcwFYo9
sj5b+MRyq2joiHddlAhIoTkmsK8cS768NyhuoxNT6oNGT/t7MSry7NFXc8Msvlq3
ygG+uDGuYzM37+KFahJfRNQvaN4aDI99c/VhxK97wKlkDqcFOGxW6R1hjjaxn3Xg
hwWtMsbP8VwSSTCvaVzO52/NVCKS844P8BNJw6tJ7e/U+5cV80LKVxGJ7lt0PtGo
y+KbFnADl2nV4GDcJ9gKz+Cp5ZsWQ35YjHKZ2n9hlnLCgWK6JXNEmU2jt+Sdqpor
xCEs8SLkXeLsEhPVJHMeANBW50ZK6iTrMk6wnITc1/bSM/BhK5m9bv7wHq5fkT9A
sRBhhlsZu+veaR6rxhBUb6KdPELQgPidxucc80/i53vnZyDhPR0TKnV2I5u7MadW
FC6vpMb5AJwGNxjFuEppK3dQdtPNBvehDPtXnRlcmBc8yTDPt0WPC17azkXkDF6p
VYmBNFy9i+374XJ9U2+SenFf+Y8ntUFZ54Q5zX13rJwgwA6jHgR3CpxsrFzPLNGO
1aiBFlYJRHLxF3aNiH8pqJphxhzJJwohwZKFeWVwkWEUx1/aw+laVJalzlzz47+k
+MU8EQcqxBorHfBr/A6r4gU0b7Lt6r3fvbGTD22NxcnRUbZc1lTaYH098bCGJ63k
qUX2jPKDxl18wkC13ykG2EKNDVaPouTmxLgoLnjgS5kaWfPPJ4IBOi8YpXKF88bi
yYePTSTqRDjQVADgy6wX5ns8qZ6blwLhy3hF4vPICtHMIjMfUwAzpSOdDUizL9+5
ZqcvGw1It45S8nGqtEN8PY9jiOa76fmCYL4v3CzLg5tZGSFkUnL2bPahrfFfBQQ8
7qm7o+/rwEHja3Lyn5Ru1PovKALW+2CXC8+u8BsDWmxAInI+lUiULenrbGByVBNI
a9W4tr+tMC4mzZLarAnXc6lGTtDTVjb97mWbPQtPPkxn6nlVTRWQEDuGDM6eZxzc
GbBv0Rbv920N8puBVKXkC8a/cm6otq1X/HoL8BjUnixu4To3jguCVKyBOH/cLC8Q
3Ly2IOq6G5EF1npmNLFBIKp6YCsnAmhbCVK2PAYWVa8JvLP0XcBzQVuVfcYQs5k6
rRLUMnLtMgNX9jdbOqHVDX4Cznh/aHRKMt7a3l+5RA6p6aGLlaBKCR+aLFyTzYs8
+9hm11cGRGZcOuHmhVKbwduqQqtxmEW8aK+tdJF2E0u0zYBQ8gVyIwN/tjz9BkYU
q92s1+UQcNmnx56mAsFJEavduW8VUW00x8HvMQ2JH+C8pQKP8IvsJL/IOD1xsBxB
rUW2qCMZzVfYzFy38rDxKkZGVDthHrNLh2MBA2km9mSkLXYg3EHjAh3nJGxAAOpT
gzSD2cehniTQVgt/VXkKlaLJPqGTpMg6wrCMxuIM52hywfVirsbQF1Wyw6dawAHH
WnZm1J7HdBkJlvVb1PN90hCal7G4LKQbMjy/ru4AHmTLg+/Ay7CG+w7C+iIV6zm5
0xn4r45qrHZaPMhi1y8dqGOVMhUFWSLtS6erCq9khNgdYIELnfKj5OfY0miLAAyh
z2YTcpg4xQqtDcrzW77OCfPp22xGYXug+esVAjRXLwh80KZlW/8GDn9zw0SpQOZQ
HCh9OosDuq1+kapVa7RxydKzZfJ7v7OCLHa9bIkJRKReOlMvbTiBXOKoqsoFwBRP
LSsBdG8FF4uEKJjTW1AeNiFDOzvFWJZ+wG/P3E0vuxvJwbjE8SzdW1LprSUbWgSJ
O46bYCVbsh71GhZmGjiBYSsm7yW2Gb0Iyc1T+hLhHhfVOEjhj+FF5zclUV5IGNaV
2R9yXNTYNwwZEWKLH90Act7IRae7ZdNacUFgzz2pBx8nLXbGd/PRPkhhCFx02KSU
dFVzTHPk3zS8e9HQffPEQ1tUtcPe1Uyrth/MbA+juBc2TPiWK2ID7vqXmbfN2lk3
+OfmJe1T6iboWcAtoeq3iWmLxbrh76lmv/mx8t30YHE6yet6M7zHpGQ+7odpBvwb
l24ThMKp2pDLukj+VSydnvEce1IQ2m0zBCFvO+eGc7UHRXTYCSsdCxkSKsA1JDh1
w3nQFdTRgcKfjeiy09F+0z0KV8npkCh/Z46un5kGhmWSaJQFTWL0SSjXWiIa9aGz
5ecnteTe1I9Bt1NLqYAl5dOGVGyEKC9bQCQjVnZxz5cbaqk1umByGwjLpEbETBCd
QQ4XgnjwecHl+CWznoUagLDN39V7sc8HpjE9bpOqBsDSBuOcDAxvSgzfT0NzFNFq
n8DV2udxiPakYm7jccS0VrVYkAj423W3MM/iFTWFyETTW7qgcocCfWSJqsqhf6wD
mOESem8bKoCi+iqGLM9m0YZrUhV6POIdGb8BwT25MCthkiFLziZf+89q52bAeY0Q
7I8cp6KeWbuSaL5inJJVEcjLOcNyQctVtR6uqX2w7sOHHnYqxlDcNFFlfxfTpJ5A
pTLHxxUmX3lH7tX25issP4Ah05nbO9GeS0G3ZpqGeTsPY4rSORcK50MUpRbJ7Rp/
8TfgNZHhVThqFGXoZPphkzW5xZofgmEgbWqG9S6Sq+OBrc2ko1yiYZgV9KCERYWT
XiJxTkkCbZpgMR5GR2YtKpa3dRU/rOqi6CFfWw5AB15ogHD6siiymuliXh2GPTW6
DOzlwWxYbPSH0odJQLsrmV64SoxsiymCANaMQBTfbTz8ZRMCn5+4g4LPskGnBP66
0bUHf76Age5c2gvWMyGZY/9Mw5lfns13jq2cxsMWJaBaj6qPwyEf2zOeFJk7+Nm9
UC2kK2g2WuKG9tL/SAFLggWpruCytQEcfW4j7Y9faHqflsCD5gBV1vwxo3o9L123
YMRtxyrHQEtUTvgbtg2P1OuvprmN3/h7juK6ESP12j67mKCOrx++KxkkKOP5J18Y
PNXbuHFOePUxpy9MDD2dhNU4DzNzS39b7DhOUe7ag/ldetTIt7pfe5cyIk9liW6t
t9sKblIKWQSjsBolrhiPxzWyC5z9rff2wIRBNE/zLIM1sXK4flLx4ndRTeNb2cNF
65bAgQEaTxyAqYdIBFTAEu1AfANAsjUXF2IGubb0Fe5sLCkzqnzo/OMxDqp34HZe
020bH8axaFek0g0HkcCnTHjMYvOQ2jrWdxnly2z0zFNixGxh66lG8ViIUgiSaejT
Njxd78QEEKIAT3f5UxCt90iDOWyUN+U1T9o/5VX4Ugvpup2gtU8gt+6rXey6z9Lb
+VCLuZhvgVieor/hq+GwOK6KRzQlPlwcSuMXxOme0x9uw7QphpmvvyWxuSq3nHHJ
JzdjMqqRD8InteELfXVHk/raWEcxbCK165+5QxaREFh9E5bcVbGzybUZhwxHrSUh
0y2h0ARAPibDfeSAEsZskdW6L2Ix0Jatgpi6BTuKhgrsub2AfkhpuLS+/yvatL2v
Q5yaat3wtvN9Rm/qJswqsZW3ucihzaK834+SctKqKNbZ4UQVqlLWbMd5TvCAFuFw
Q821TBs7u3OersZcKGDovujidVaaU6wCWYwmFSUVzbDk3WCvd4QL51w6oQyr78Q4
1f5827bP9LLWczmshjF09wn1TeJSyJv26aAPbBhUhWVFRHuL4KktMztfEdVtMg4U
JTGj6B6TeBRGlQeryMZZD7pWoyW6mxCMwkJpQgpyrwn+xbiXB11a9QPDfOqOYTJR
Qhd2gN2gcM6+N+eGJf9ftC0D9go0a40FdNHTAuOC/Qeq/rVIFTz60zCSlJ/uaCCV
jGEONWcSEpRn36RZVH160dp9IePJxjahbB8Nl1tHLDF2BfLGvo2GVkQuf5899O7z
hBscozAiC92TSQVQz32LLdo+ItHkEgdW8pRQrfwUvRDFmZY22b4cz45Ul9fw2dOD
X2O7+V5UIvWkAaxsoYDU5YbH3AlumMmu4HnD4ozPQWmrv0kQPqtBBPVdLiq1ymc1
cmOnMnR+3+X7pZMlQATnEKLYzO0lLCEhWs6MzLmqKUU9r/am6f+59X7zZtkJzd5z
XXdN2UTdFjS9UlspUXN8aUVPDq3cn5b4qdyzQz/3KNG/rCeZxjcL1pVU3srMI0Aa
T8PCXqeJP5ApPooyJ0N3kD7q3VTKeYTD74dTjZlhDZDPYmi1kDr6vCYEkIeTh5EF
zzJNJFNuklSKBryLOmeqECk4oJqmALqX14zjwZB05ToFQTLm8IhrHfvTkIw+TgJX
fSabr1bz4e6UXWcVOhAVkhZ7zKWLGB1mWUnGB/3kYsFdiZ9mMA5pypVlUoqr19by
/fRJ1v2H8SBCYQwcgIIcwS5qfm2HaaP9Anb5SF44bOF2uzXQ9Mzipo+AhbCVOPfE
59xU6gdbRRS2r5zcX2aMCj1tgmFzknebxZIkrZUliNiwUSX30RnGUzcS3+JOLiSr
LTCwbU7atom32+Se2trX4EDCcUH/HcG8mfUJaGYIiaB/8R6gwbyzzy1MyJDgk5UB
AOo+4QJVqI3vG5jmLChCYzFEKHPy6ptpq5wWHGOLNdtymfS1DHyZoaRgaQanvkVb
3r/eK1To/7b+ruWztCS8gxGdsesfNuAvfSKgjcRoB212tRC8GcTnUav7ZIpHENRu
jT9pXfsrfQ43huhp9ZFWrKpGAMr1mW9SNCDx8ya35kvIwSZDJJyq7RyIxG2C47HZ
N8eugpV9GaNMCkK1ygflr8R+BejGHM4UkyqLh/jeTm/y61jQgkDhzOfma90rOBXr
+XMVU3/cvXH5W/700V0vl8L9h6XeEiyJjil8c6+tX68qGpM/OFmHAdT/a1tftffz
mmRGoiw4LUGEbS1CSFsY1sTZu5fbt3oC6J7bt2XbEkXpsOlMYDf2Q0wmeM0yrY3K
v+6i/FkBJiVuFAF0974kMg5/aj25yTwiqRcxGdQl0uV4qGQrwpNl+w5s7HlDiYyE
K0jA9I95wPFIFE0fgKcjSf2C2PJeFlG90u9sUoPC1TbbxHxVlWYAoN02zFka7PAU
qvvlR60Ac2qs7F/Y53nBIbe62Uj3R4xveE0nU9NLtU1+cv+K/GLyvIeQhwEopX/B
7SAE5FZPPlB1QXZSu3fyhPVXakxjA1GELmCP3+okIzg2BH9pMuujed3LBARlqnog
AQcLlUJXNPwx2KFes9cNxuN9Nesomca53yeHFXA9TiBjAlS2IOtorlQ7FlK2Za3s
h+FLigOOodm+HWtv0dQmzZjEki/zoS8I/iV0hTR8zFIl1+KVqdHXDbt7E7KyzxO9
ZXRfvzknKZVUgYGxTdXwZzTsgoUIzYLt66UXcTjR4s8kwX+9R9iEk8as3k+4eNrC
XneP3x1MJl+r6DWATy6crWLVWYukhg2HL8Hb8n2TglXDCCzlxOy6NTf08TvntsH7
T6ZCXzYt7JvcfpQ7BbDORALdaMfsSFGcQJKCp7I8QXVK9Wc+C6bgGgajWP6yOTEO
CXJB5UBgROmXP2rtbV6K2KBsdDMAZfGY4uiFIvNn54T73FlCivmGiSsBAQsYz4sq
mTGQDwXYzKP3qpsha5cyTAYAwWmgYzzHemzNne8g6ULv+2AWbJbdDck2kIX2hly0
SbFAB0eGin7b/hZWAld3Ia1L6nJXI/9nFgCb+65FyeNvqAjUUnfu9/04Mamb/NCW
8+khEK566AJ/cTPrThA6RQO70q/iuX6D0EBYy8nme8AR4HPcQTldPbRK1L/zKI2D
pUq8CL6B3VYvIHae9d8hfGZW4aBxjH9dnKqzitUOMzIPyu8qh8BPEv6uV3VJAwRM
LgD+XTXInrYWN2d4WSa9sMHLTARFyDG6NZ5ecLl9VC7qiUJ9mJi0j0FgD1/f8lUo
qWVoWYRyDERVr7RwP/wzuzIHicsZSUp61DIglR1jZpnhx7SGKAiZe/cSEWcGaPtT
Fhsr3tM+BPgZUTYIubj9wl6+/dxaHAyH+h5uGLqV3bNh4FJ00dJyWxb1SR7+Xdox
BrKjJ4CgLTSgAN4yucQ+YqP5Fl3mz+Ktc6q5Fm4CzQhDxr8h12pZuC7hrjKIt0jo
v7ErYJnlhDQ/Fus0r9I3oPOFMHNCeyfQtMeWWzGxUcQnI81WhWm1QODi6zu7WUTb
w7i54PqdCbLxKwLKBcBQsdmg2k6AQfYKHHk7Lkk1zerE+ZAy3g2lmVaxnx2F3dLY
9dRVF/Tvviq0BWVsv7FBswI6SMjh46OG7CeHgdf3pWTNv6abhN3UvUQY99F5iLkE
zypFmRivq1/2WimsfjX4izb3QABG7p0Duj+XXlMqRRl+Z4/Jjbh1I3tArG7nd6/j
R40tkFnUtfyBtFeo+/XIeCfH4twdwg7uQR8mVSupbUDLymCpwk0XaFE8wA9e/ljn
1d+VOG4M1ohtH9XseZNcWx1FBF4/pd4muu42gERQnMs45BL3ksQHhC8hZncTQIVq
D0i7cYsZR3jkG6NVlmhbfngrRliD5dauwiXVAfGtDbDxxt6yhBah2wW+kO6Cbtnl
M+K+HD7s3ERTDJ2W+0j+s/GQw9397EsiARzfkvDoh5tYyNFFJ8yS6/G97N1WXAZb
sw94RH/Mc4Iu0cSzRKFlTqVz/3TJIt6SPzxObh4/C6Rfd1/yxv3nRgfpVi2FIGV3
FH9Q5kxYxLuctkt6qy64Fv6sQEuh1/bzkGQlScKZN6iYP1h/Gk2ELUh9LpwF6XyU
YFg1PXZBYwQRXaRJuMsNM/bQ+24QNfeTVLQHuG/4Nl6SUboQ2jhtI1gWyjSsXQ8/
NqJclQFuZvVoQA0jl9ndZ0R43K2ZAAk/5RnV2SjDSbKzwwI8jL+3zkAgPkEMqX3M
JWbUc4ItYxV94T+Jq31uLfAC8NS5fnd0H1EIRymqhAJVEtDlxL/XE0Wl7UgVkz1j
J3FuqC1l3JIvNsHZHC1FNYPhe4+IzrMxYpoxSI34bf3sftR7X2PrkpBg8MZFwGRr
F/vJb+fs3LIpenePoQJAuqJ3RRRziuDC1Rem00Y5u+UC82DNRwAI2jMnj2kw2Qwa
BteV3zDUSDyPus1otRoqhjLT2FbUB7bYuxyMyXCVHfY0+cY+2GtpjVrzmkchM0IT
W/dEKojwBzadtajdmjj8f2NM9r2c3oW7Q+uFNWce0jitFGlfVSIwX9YZXwA9K3Fb
OnDsrxWZgukZ3G1K2hpixj0aoQR10iyIa4Kk6KheLTIbJKz+vDtpCE5CZOZSJMvs
Vae02/SBP3FdFQcU2OQX+R4wutMFAGJwgTEoSWmka0c4WzfPnHOtE0lA/K6Wjx7W
lxCc46Wr62fB3UREMyT3/XKOmO2+4zP0Ef7Vu4SvT+Hv9PTYXaeeqPjDRHNp48oi
KRrXfEORsKzN0j+2KHFDsJkEyMzgi3HQ55NPzue1JBPOPTVs9OMe4PJOe6xUiF2a
gq+FTqTcrxgZEaBUNwCt+ImiAGOLX7m/cV6cL8ev4SXXLEmVC2V1Bm5j2a7kcsz9
bw3oeqj/ow9LkzvIpalDaVqjJzETAKoJ7Oz3URJKi3WtlfZ64W5WDd9OYRk97YJC
2dZeH1A0NopDvMm8T5Q0IYfkE3BNA69IIoTZoh8FKHLlAV2eRwkF2VLaCMfJs+Ry
UG2cAPoVDUmANJcB+VbtaBU3G7GLXBTgxeLprYlerI8EEsdfSv+29TN/Od3dp7lW
imxr6pUt100Kh0x3Q63PHEYHMCJHNEmqTyb2Ftz1qzS/qtDv/5tt6ZbZUG83RY6b
8ijcdqD/mh/wiFgz0SKH/jq4QRDZ2KWakSNKxQVVXle1S7OEpYlYCw4hbixXWmz3
6BGWF896PfylogAwni2TVBCirvV3EMZB0BA15KzVlzxzZ/FW2VcAtTBta9L/zHWa
d1CpWY1jO+PtfU06b/K9scnRlAzUrAKLUB8CQBWoEUvK8pTrpJC/tz85D+UM6wME
QCSNUCWytOVwBoAGN5vy9H9S+9RPNwDy0VuxJKlBLnlAnGDzXACgo89W5Edn++cn
lCsH2OsPtBlMfSnxXDu14ySjstfXlF69tLqhyxXUZGPI/sEzX9GlFc8mzCF4E6vo
wFSbvXw2gINBhiFKHcpOi3A4jPEbHwOfp2PgA2yzbta1V3yZHcXTyqYgq+nRgegv
o2EPIWxjTaiP+1JW2gfyri3nb505uqCDffjGodsnm0N97wRB1BPpav/MvXwHoC9H
dycVtpgcyRTeCWbUMhwf0iQLxdTp0ReUk3A53TyQfqQLPLYfYsbOr5+qXtaovE/I
31hj9yQovQbuMghXk8TQadlcO+k91g4jHCf6SLFsGqxLY8MjUn0ZtXFy2PnuIx88
3aHV2Fp6QtRL/1IjCG8uFM+urn0f9QianV6eTL6UiMJ0DEOVjAGxMRaUH4fESmZe
+ntlGBEOxdof1v9ZGKXL/yQ+S6rk8wHoTKDnGzCqb6vYDiJAT+cyvm+TMDqalor+
TjXeOiL76prQYU5fg3ttdrgU6rq8/GujUh8krsvpxPTRIWUbM2dPXfBKm3q0in7D
bk7y61FrD4UPhi8WzU+Nwq6vvd4DeRubLGR4z4JH9g/C0TCElXErgmPHpNTJrCA8
HcILA/oBvvq9N5zLNqqN51YT3Bl7KljCYF+OveNW3Sno6k4QlYPVbYfM/K0iU42k
3JE4Tw4DHBfe1QyCfTcoD831UE7uZ622UU3TEEWGZ40yy2094XLk3TSeIwuGVEOn
YKNZDG5t9OxoG6Cacx6uEPkVC/DfRJf6ekRk/EaywOAucrhSDEtz0t5BAdQ7I4nF
PyqjnzhMiBIDbQlgYlhXZlXWGWqedFcQ6UH8TqOyjyBFEKyoX5lIBeM4cmSbfA8x
vJkggMvI0E5K3Yg5KVEsINBIVy2EVkqbkHZqPD1/8MVXfN2pCfbDvjYSFKEuDfmT
IzfkZWgfvmON6tEd5jO8+pz5w3zr+/LM3XP4nfbDprDksdE2yXoO1rSfkoWcP6yv
FnfPFWhyGTTrZQSTvwewLEtkm8jkG1U4lXjqBQEUANvG2VjCYlvuP43UUiFm39v4
Vmykr3zI4qvl1BcVBlZaqVk46RO87XCh4QQ8uz3cpe5mhJ2ISrf0n3sE8Xnpw+ep
rV8wwKmCFz0DyIE+uS7e0YIHhDMT8IdAaxuzWD8LAwLpI8DaV+nI5abcsz5D2jRL
4vf40keVg5eZgEP0scm5tD6k5sfcqIKY/lIOgxtfevjaV14xYIk5esbI23+F9pNU
7fju/cAt5KHevvcvOZGvRKxkcT8u8JFFn1Mz3NSTuen1anDXCPXJMjlSNdx5o4ng
vNZJqELc5LGvTeyYjBv5BEXptYCo/zlz3DzdAVdlf1Bn8AC2QGxcp/a2Wyzgb/Jj
5LvPSA13lDK4b+V5VTZuCS2MdJePAsiRk+rYWC6CI4Zx/jyTqGNKjdkfgbO0+78H
jdbHiKIr2wK6hzsF3a/Pq5aEx8NjKifUA2NnKoMscUQBPkZLm4O7dav/WzccOw4a
pSe3gONJvILVmyh49glmSiwAODhKaTvOc3gAy5NAOjuWBfS11cYwdU+GrsmqONCi
9Uqm4Yefc0/+6zQWw/k3rRWkq+K8Elepx4bkJ+47/hEuDrkacvrIgGJAQLov9V19
304OceKLHULMUP1+9shzlHbPF8of8UitrPEqK7PbxSkPKkZR+Ib8nZjQxS6GA32G
dydLcelXmiuo/2pmzdNyWMnwnZ6y3HGVfnrq1HQVTGbO76VUKHmHreMIyBNs24Kh
u0r2gs9P3VE8zdnOK5/GOqSwHbxSC3DRt7EvAgCIPnQHP2CDygGS8F4Gfke8Xj0m
q//j9/KbBtXJRctjFZepdLEYV54QytHWC7fz/v0InYXwwLZF1AJZzjdcn2AgH25M
fwUSpQ4C6mG/E8MoJuEhv8W8ydIci2Z0fc811rxyaUe3bLCg8l0eQDaR0N15VOcM
Dw3Tb3AewvyeAMh6L6Po0PidgWqblNqWxqkA7dT9Vcnbw66iHU4EirRc1mzHSSE7
BJpACw8t+Dxu7nwqiJ5Om87qDn1+QJasJSwIlDEk+ubhQxzEcTrCRdWn9+It2zhm
s2nv2o0PX8l2ZBpAwpHKNvUa/9lEWuZNFGaZS21pt7ZbGwj4PoYkb1Jg6KivHqFX
SR15/gPmPmQpl5REBVlpYfVBCjkWGNH6riRW9coRvWNe9ClDhoYJ5K2PONX8SQoX
BSF0SWZk3pdXdFdTzR/ViiGQkuq+FamHSO7Tfiy0vBgU+j1wMV/6ZcqbP1PPQxUP
+2X0gf6hlv1xda0VH8qIKKr2GAIBbqKRQ+AYuUKxEsR/c/jRF4ahGe3yIY1pt0cz
PmmIybOIb/D79JvrWxGUVqiMCg4z8T3n2EjvoAZS+gS3PQmly6uOFcqOeXadDFlP
j6qii21eAEKvvaXbHN+1WVTyNsQrITZnwOpEARkS8o4A3JlnPqtjcjpM5pXqZpru
apHK4rOdPkq7YuDX+DtZxMKUCAoNITFV8AQDVh2Ey/Ejb/45WXsTqb2w/jnkQ92d
fmOKYnkgAG4TzFbbNwmmPKwurdcu33WKsWUCJZvRHkImiMGX50Bp6xFmMJywSMmN
Hf9dclIWPrXOU8qTzet3xOcAv//UHcRu4AEdnAiHbL/JBd7QVhfJjQ6z2bDLzBHu
ux6kvhTAtw4GI2XlvhzAcEkF7MrYbqezVQNeuQiLZ/4VudCj8Z06kB2wWTp7OFIb
ap/gk4KB+lddarkmi9Sx7J1bGyuW3ftXPIil5XM7oXEqiXtPYzwrr++SC23ArRM7
76l4O3zSfD25o0xzk/NZDJuEsoSmQENclX8+O7jnWj/EST32UsBge7KwjBkz3Swz
aK5FPaCDU2FfZmpXumxGTQi4sU0/SKIjslcQKOv4IVuZwQHWUuMPN+1DjYN+JqMd
mZy1Gh8AmxcwJbkbGsqjIf5i3x0u8MMli65qagIKUgdfbYEct+u3Vh0P8GjhNwxO
xF8r8++pTyCGwRfvz25uXYmItE8Hqaj1/OMjr1bh/CWYDVAYjRfg1Dhd00AitXrf
glNC792P4eZN5xgkvicYgKIDTg+hO9ANG31nqb89ag7iFQqeQ9QgniLdLzNllOzE
DfhkD8zGGfrc75DpFEUHn2pGEdn6JcrtObX8TLQAXqCtJze0Vr5CKDim+oWScrVj
zcBoO20NtA5VOgHXwfVUKKq0kXJPuS01VJ3Eky19RUMJgdZOgT3wvui2A1lWAaJk
rKzBafIvspMo7Cix5GNSPc/2IC9P2RcEvqk8B1+vL9ciuCiijKccf5qhk6q8MTld
lpmxxQp8iFsVTWaYB84HZqcKCIvys0YrLN3gYdH6LWJYaZrjAJIId3xHt9wnLSDK
+F1+ZCKnLbU1LUqPGCzB5ZSVz1xFV5GaRauztFSS2/T/T8p8uqF9oViT4HjUJbCv
3BY9kzETUFrYGo2d+Ly/uOVzG3SCZNaCbC+TkzrHkS9B1zCsjEbU00t1IfY5MTkY
1ITW3ZTu4TonSCtvjaHgIkipPh1MBSkfES/nmbYzSjPD9TBZYg86c92YMjIvVL73
Vewtr647IQTxdcs9a6iw0DGmmyBYkbrgUoHuRAnfz/s7WI9bfEA6nu89Phz99SeR
mf2n34uOPJX53e3Ir2EaUR9uabM+TY3tGF6Ar6xq9EUCdkpzqG/Zvsam4TlUx6aU
I7wFDvYEO1Zpmfo0C1xsW2tbPWMJafcitF5wvXKxURkkNX7w1Mwi83Z+MOqiqXiY
xNmAieY1Ip/VTtZ6iY5/x5ylkKnRXAr53+nw9FmxpmU9qYLtPCKA5DW6lCBbRHTz
mUXaaFtjH91rMG5zmnr6ABmVM4A/mQFtodkUysB/beZIZKiV2rsSwK1DRhJ5PfSI
NdSsz2Vx8gPQUcvY+q5Slfe7QZHtsEmn6osD25JnkTLO2db0VyX2arZPjwSFcUwb
OTBBEL+MhUpmDrQLG6erh5f1UJ7B1da2RBHfiUR21YH52Yr3xQfW9nEYUrTFhBeY
1E4NrKyEB4fbxCi+JVMmK4EtpdqqK+N3RqMyjLdMCqlKQKhPRkJ84LpXHUN6MUO8
/44BsBXr4AomzoZhrdhPZVLHppKrAt32hVlsIF7jMnmpv2IU7SYfwetGrMkezhiK
Uv88VN3ZLFkHP9yu5DeKrGB08J1IxHc7djnFzwPWzsbG5owNxyCAgmMgk0RYo359
qSceIGiz0ZtYh00OA9Gtmp/R11lRU++369bJ8/NceJmGJuf7LEU2Df4yOvUTWAsb
XoT3QuJZ2wgk1wv7B1gvADn7RNF6WHb3h74hgXjbIv2NUuw/TVIMCCVnsxwACV39
Fp12lAs7NvPren/rsXFMN1ROkONvjGWHVOa0pTXCbBO0BXpd7ss1ZDgB9oGxYvGz
b0rjolKmiIA5btYJNQI1fo+4CkJ9BbUCibVnMtfWPu/VVpoZvB82/8V/xwMuzSBk
22fkbKHJbD6KbJSQBPr9arc7lKdM+ylLJh/kAnEiinDZ6gTo/5K9gIJ62Xj/Kzrs
9TTtHarlEqoqT83xvtmEteG1dWmuilAHmE+Lrj7tlyDLklDG2mlmSXKtJgjLJYQh
jAHQXG5wkvhJ81bOC2JatQOo19teL/8MhSQYexrSvUalHeVcJgNzAyDv+8eMsr/Y
K/AJIq7I9/Gg534GEJMQyhLtQep7v1lacdWfyphKTeLo173c812sIMbF7kZtwf0M
T6N5kl9+FvgjSa6BbgdwM+5lBG6prH5BstP+LXHHJjgB0pEGmzPcvN6Qe2fp2+Vi
dW78DdNL7i65OYM8LTCPsuW6QMnrD+BK4rKJtjQ3oY6jE4rDCwUkXTfPSirpMDJz
9ckhoI7jMCwuXPu7LIkCn6MZ2Tx6KdWciHMYkFB+mTpBXblfQGaBe+T2rfqYfij1
FeIgKT+COOmIOisueUwVFuE/cpUKJrXwGyj4umRu82XK5YBnHgzP0/6f6w0IxBUi
tX3fclbGHC9yXNEqJNIk9tjdqzGyJtYgAJo/qx521YchXvkM3zi8SrS/8LCuT0Wx
5dZ4w1hWKaYDmJizxgm5O9LC4dNkq42LA/ukVkIS3S/Rd4Tche27NDZWbbGKNqOD
MWkh0YiOkyXS7i06cR8O+I+yK2jowEfxE139VtaLgLRaYrnJd8XL44rLEp7yCo3t
ifOotAm7nWsHrQQPogXpg5dOto9sQPmn4i3BjbgrIlrky0Y4q5xRmqufvNrQey5C
nWSrWb1C0KUC54ZDljGe2dqTYbjSc5qvj1RW1pbbBK7RcKDTEi9+Kgx3OXzROF4f
xmxTDXgcq9CY2An8+g6DHajJou6ULsfquoB4/55FftZhajHa7Mr1rWaRtAwhJa/8
w5/8gju9llO3WmuQ0zHdStn7kPQjXVNxyT/+13K2Uy6+PGnpGmc8lVmojvEZvyiw
PVFEOew3nPR8wgtc+TOLI+YqEU9GtpGDguWgFIGQq9fwrLSudk2z3uebmdYU7UjV
mRDFvTuS18W692Ojj34qU4Wvo3wgrCld4Ke/4GvOmhrewoIo6PpaF7PkfJts42+q
IQFJKwZbUQXdqHlx1q/s3G6ZyPwEgSelWZB/c/eLqeA2mCta/yQy2D/OnCVlplgo
6rFOxKoJqH97CyOXQIaL23sU76LK8eqlwd1CDU3rSd+nao5nz+e+/OkWZ914QNSK
iscie/tvQhfm0ggd5j08INzRc3kMka9fD6dmDDg6xq7heijVQu0s3b0vXydhVnQv
GXOjZrth3lG/r95c93D3okqdi05VseYJ1lE3cdR/GFkIri0RqVdYM7XOwZ5L0pIE
gRcTPZaXBq1zN99HEgf+OMk/R0HzIlOJl4KlXzQ7lzpTu06LHASAG+pbFnMXdwzc
8k7FHm613jxYHhapzugk4ho0X0gdEuDKhS6+GFI+3S1CAt/63v0q/1vp8E4a/rTP
oYSkxJqsYxMLAevL7e4rdLMUFGdYL3HxjrAAje4tZcTXoqnMRu7/ltnlQsGer9gK
x3w4RcfpYrpf2CCNUkrJjclt+FVNhPueGsLrN5iTeeJm0q3hZiaJEfFCnK1EZBRN
0U9+xcUYSZKD2MvpWqkZoDxipkU8uju5CAAzyeeMgrLNH5bzznrP3oW2nMQkNUvg
0nKkgGsdsoL6CqSNvxy1otAP6Py3zpiiwR3vQk4LXk6F1/S1joPmkLosvA8iM+LP
yKxilCQCcreXc6nThMCMwf01OllT7uFVXVlkslFv63qi3AiH911FBviZIJfrShGF
RXoe/PoiVBHloEj1UDTDQjYHcPsHPZOIzutSpQx3FLZpGuhZuWp13w/y7aRKPJv+
uUy9NlcazeOG5peKaWPVzB8Cdo0Q6rKL6ARm76FJTqT8ecjCIxKXzuLuI++x/7+7
4dwU+psF2dVmVL7Z+3PJyeFtvO1uLkbQWkz4XNYUEuOIK8mo357m9Hfo/mnvkkgn
PDDyGlVE3SdC+Eln/QSCnLJYORtahMVmOPpNRsL4omvN9FF+4z+rmclw2fuVmpQo
Ool77kaFn8yAA9CxOdsQI1MEs+qxBqyAl5eOui9M8wtPAYnwYvscaSi+mRv2uwbz
CQRrNsydMbxWzo4e2LaNn08l5VPcbBdOQZ+XqSwKZCVPMtyBrIMlcptk9VP7bDLz
d0hj/HPv/wSq/0nOKJcMskSsF1rlbL9+wjOyt/4Quz5Cjb5d/8WrBV9IuCPxKff0
sPc105iZbl+JN1XpbasRfMadizBZe3YIMDFWG5soTHybEqYQw+P0+RJIawz+n99T
/r2bTDmMg2hapfKzs06bS6EoQA5Q2D27keP5H/P5e2nmHnO/cvHQ9lrOtQZ9mgw0
LfeTNfwvy3mGQTKFa85Ndz2wGXYN0VCVIdn9/Jxh5Jfs1EIQ4umjYIYERSNPAV+k
Iti6I05WPAcQXcNVwYADBTmM2Y1rbBoYnh1vrLGuNWJx2PwEsRTUevYDUOKbftdm
7ShKNcc79RlW30EQTqBIVdaC7auIHGaMDeNPjApQXZ7yoBJHCAIBG3O/maS8Q9iL
sKgXH8wTZ5lFHcY9iotWbMb5yEndsPC7iPwMRnqZHqQKIAI+GmeMN9kUiAKXoc1x
XHsiiOsPsRTfsQ/p++NCuT1c59B9n9rAlUBJ3cYUTqIf3G35HNV8mlqK/U40u1VL
5L9WMeApobnkIq3MjWMkqiSY9sMMUFFh9EJvMZlA9w+tO+Zhi16aamc6hE2/0Bhq
RHzIlpzj+dXkqJChNEIZv0X+vPwlLFpAP5+BtmjEPwvwv+LH2y0Njw6BMZpoZmRr
uxN8GMIw+N+Ux1jO+4sHerBWfD8yjlmauUbfWNWWxpTmMM/SQ3LhyKPaxON6KKXJ
biR4+M9IXY29WZ2NPVLUxWx4/VeXaloguRAnCju3JMwUodijis+IkxNxF0xAUq/n
NEWc83I9ouTJME3dal461JzTpfJxfFTrKJ+vKSlVP302d+G/QCpqsisLnpkOBJ7v
vZKiehmvdI1trAk8MzGUGzlphnh175D3axGSu5QbZNdVxwqqM/mcV4lpxJQkUmYZ
+7MBRPJtioLGtfB445YDwhojbd7/e3QCkHR1OM0D5mu2GPzXKy6V0EIjRbZPurER
sV24ebMyNn5fL+MLHBBlGtipBdCK+W8jCApuysSqKpiLlEpttnMkzViVDcTc4A+a
PVAKq/KQCmj/Q7+7cyPmhHbnMuHQlSUKamOtfe6N3Qn5P/f7ylbaBV7puHYwoXis
KKbYd7WDncRLZpRqlUL3S7md8pAUTV2OV+XaULOXzNmJQ7FACoFEdZy4+irXBu/l
PYDIr/QwtV8DtAoufF/qMoiI/0t3INSaQuhADT0ofy/uxVgnIgh+XVHvTwmPdb2E
yVZ5pYpvp9MRk4hMlIwr6V5EUB150oshV3tvgdJkRBazhk497jfGR/At6QzScMpW
uk9cAfvbqCQ08kor52/Cg4x1Ev837yV+l2i2G+Fd0sB/rTQ/BqsD1n2dYDNmbvcB
WGB1P1YGLGMC6/Zp017ByhAWC2fT79UQFHpFTA/HWetC6whDNm/y2qQNet4/zu/n
mJkI5nR+bPLUdIcUvywXMPPmX8+WayXG3Ph3dTHyvWnHQK8kC+pYMU3BNzA2nect
nTiDEoOaYMG0oFXvWV7gxBrVIkT7+rJdWdA6GWmhh70gAYUkH4NDymcj/b+ZE7iJ
7TcBaDwaxKBKzNcAZ7UR2IFfPqHzPMTbDKOPj8MOyzYP4QoUcsMfR768NzSrTtwn
yVfyLNX00BUOCcnyeRYlLSKOU4l7jliux2KF5ciVl9wK4DI10pQ35wMUbrX5ve9c
T04dt5JR9ome9YBWv+CH87iq5YzL/yGUur88vsOd7bpwCjB/cewkJq/TKRVxhBth
NcEruyVwHJ8Ovjsgi+f+M9l954TeZjP6SVwtsfzH23DwZiOVxls0FXWLl7495+ac
Lj6E9DcnJkbAyZQEXooqNGETw2viUl/xEx1/5FQ5z9xgu+42L+yc9twyjavS0dJj
pcVX99fgSHcYdg039rhiMHUM2JNJ4T7uqFyxJXzXxa3y1adWv7/IS+bJU8J/Wp4H
ye7REOi/qjNgUp5DxPAIOx25UcJqN/S5yDLXNVprBCg2YHIkPd2EyiDPtWuT1OoS
K5coC6SaxgV3uXit+bfoC61S9BMDXR4MoZShiH/eVdFlR1Lx1C3TyMFvJOjIB4EP
326AAH6ZfTFo8S+k4K9PIJbM6O15ufagammDsyaFbj0v+5ZxDwf64/MYdCuz1y/E
QMwvlN1nNAHBZ6mFpfcWnLtsTNoXz7bxp3C08wf8kCmJZK49kLZC7dhpfXCUYIV3
cKaqmx7udt4UgrqQfk0vGh/aHeg4p71kfUZMOlNoSbxQDBIdkZ0/Bnb0yPvSwFUj
kIl+ZS/cRrcP/ehyB1zXLvriFuj/bBBfw71WxiwBc3H4+mgP7HTAoNP4zfXniEj6
1e0Lns+pw01jtllp/HSig0l7gnY7sEp5mPkZBgVa6ew3EgflxxMx/6rssTSNcPVT
F23YVf8i1wHvp8n3iqmFOEEd8sD+nWmzNnlrqeR6mdBp4yG3TGp9CH21ZsYcWcsB
4vO+kCODcVd/pOpHSHPW4cxskIFqdvcOLes88VWZgnV8dUsDixQ6SCR7NRB5kpxF
CDTCZD0EPcj3CpmJnqJXpsukBCgjZv1V7xfxmoagmqqZzVuiYVEzPFv4O0cQaBBl
3vGe6oPy3sw36JHeW00y4NoDRp4Xyhl1wEPAdVNDlbHQHn8DsWCIlW9Ru3eL63W1
blreYxSDgk5frJt/r5OkqOaC31eMfVUAlLI1JSbcaeA/C3DlGbXey4VDskrQxjo9
mf2O5gVq82G8VWXSUy/Kah/shAnfiH9nMN2cd55ZVoM7u2iTknFiKyx9z+qenvZQ
n4GytlIwcuFN9PTeIXLqKybBc0DBzqxwZDVIxD26+3F3RN69C1GcnmyCSS47BLoN
+84bQgUzjI4pEBZS4CQmiL4e83mo9VFIq/RjxXUkNR7Vq3jROZWBvSOqk95Vl1Ub
51Ej0NfMN7ahzIUbGvaZR1cSNweWO0JBVDDaYG1eGnX4I5bFSx/4EHSyMYE9M/lH
OB5zD8z6q1j98bZCcSztU1DICrpT4cOoaJTFpagYa+3Ho1Tx2n7exSoEt26cPKZJ
weMeiIGM/ZZvYhV513BPkoldfcdj1oVPvb65Gw8aw2Vsh2ZXMdVvSas0tScEXRkZ
ZKcpxrWtkBteNspdr+z5lbd9gLiG4kEUIc4xvAFy5GghYhBQmFhtMU3T/zmV02MQ
CnAzzL7YOATvoZlrJL9szJhkIn4wxY14Hk9VWq45OErwJCG5S0ia+5Fn+ze/rdaE
T8bopyLX28PBBNa/5/BG/XCCY43mRzaGWUREZ4hHJYhI86L3JvOwHz1Dx3J4GGwT
dyBqFIWs/Cwy7Bz0UIcmvkFufb0/atlVkay+cQWtZFcWDsCv3DOyaiHoLWdAkUxs
WprMRBxluHWCheP251CVns8iOJrVv9eHsy0poejdPw2dHuOaa8r5KdrDQpc+Ud48
MuW9X1zjTFuGT/hKwUjtfMpVIm1lZPGQmQlv8hOgLdWPQbR9CG6qsUW/5kbVdGnW
z/U24IRee4k+6e15sefFR3tGDjibQv91f/zFDa9Cd/r2ajRvwtAo8FQAAjOr9jUh
huuX3Gc9wOCryfxREcZwvkLYyV4KmFSw1Z2URhlFYFNNgaUDspYNo29kjKlr5Y+h
NilRahjJ1juESNNut6kjftv2GxVcXDsCK95N/otWPdlXuWq9tdfBw2/MyLDkDxxS
gLOMQvkZLs6Y8+B74ReJNS60K3sZsb+rIziA0mjOKmE8Jqlh9xxyGD4g7bcbdoZa
wr5UdZLGDovSsXbXUH55cWYxugOASInu/SEsT2/5U6zG25T+W5B7SLB3DXAZHL6J
vaeg9iiPvpid8BZoWelBK6Ph6G6TUHiCn6FFddzDujAGmbi7PKk3d1NYfUg9G8Pp
YTYkFy0BmF154Nu/GdViLQsuhtYYzQ+OfD9upbz4pTkMNF762G396XhbLWHeAB37
LWNpgpYMeH5SLrxItUu6HXp34ZcAsGKD6SdrbMJcam/swar4r4sQikedyZXkTa24
XUOwKvARyQr8V4fcU2BN/Q7RQKQKAYHgPOQG8pSd5ntQQcCJWS+nEcQMPN29lbe/
VpSJlLxVPZPe3t2UeV6eeaQ5tnqTt29l/0sf3IxV1uQwwfupSCKBtp1sHB1cezeK
TqQ3AOBJHcOMIRqV9QDKJg3xagEmf2CcVkfhvA1bvI6HtRjZH15EQyh++jsizyyg
6mMnZ0K6gDmCbRiHgIxvF+xGy1y/zY228YUAxQnEznpzbF3wVKTYCnKr04gD51uZ
VyUG/bZ/B8svQTzewCwqj6sKBT4a0cmfWLuCBkYMKQDysQ3JCw8JG6QLwh6kc5ED
xwXWrtFwjDlSLlsuMxLMJNzxopx/EaeEeLySpVQmrBAVfB89q0u+LnDCfjQhggmV
+VHH/Jo56Ra/1+WNHhpWOU5KGoCsbAfSebCIbb2J/68729nhAl16lWc1djOPmNlm
8NVywPD5sNybuW6bZ7rDnBmo3b/aEQQLtvYD3S3MLsOg5EOlv+byRZQ8eBwcUl2K
oecW7Br8s6sGizqedDrTH3vXRVywBSfZEgDdE3tctBEN61Nuwg/RKZkC7CuUgSau
HnK8BqFKbagQ3UueDCIaihOVybzaqyS45W53UfgP+u3RHCIM2eiQjPa4ecY8WL29
9+dPShfieJiMLqS2jlCJoxICtSjsOg+jxUCKIKCPCMrtVq2pL8LepBsS9Br0Ry7L
QbaSTt52GapUG89BHk2jfbIuyAm1++RfVV/84cfbSwB3rLrT+CQjI5eiOGC6aTN8
pQr4dHRocKZGi6Xhv7fYwW/XeEv1jtqR9GU24AtKAkOk5VEEeAxVNDL5OuipbsLU
PA6NguJqC4SIg6DHeMhV/JfliOLkpnmH8+/Yp78C9qTKaud7AaYN0++GRukwfG4h
ky/ywHwrkUkscc8ZV1Sk1td3BTbPhOJDhTm0XGrOHvLIfufcsPDbeI+qK2AhGXNt
2HNaDJFNx8YGM1oZUmkcojnVM282yh0+y3fXq5PSiJipgxRLNFcGlNw4BV+B2HMo
eHQu569k4Bn4/mCZUur6V2ye0U9z/VXCqqwb/l2pEIJeosiW5y7Y7j+Akin8zicU
YAfwryxI27sZd2UGRNvNoVJ/7tYuKHsBnBNimHfTDXX0oXLyRoNsxoKs2X6lSkdb
fckFp6Pq99V1RZzN+8wOsmK7iRgMLfTgA4p+ZNwzBKFfnziWhxBYqZGgiEKQdVLw
jHLuhW+NNIxMepcKc4QPSQ6ZHq4gmPypv1r3PXwne3hUaccpItgA1IuPY+9dolUv
F3NrChvuv1ry5mNqKHCDWghtEBe4CkYeQSJy7eq8TnZsmQi/O7In72uZkJFXg6WG
YsIYUf0ZoDUoHqkgcrGh3u0Ls2nWqcxXY7z89hSmU40QPyCGRcTXZy4Vz2EnQNlw
dPBr9wBku8UZx8Zb2dujEQtZdigmNesGlESCvnej0++sS7qFOAuiqNkliJ7h+ZY0
eTLkhZZLBn2LLGyK1Ynw5AtG9on4RScKVIr4U99+UTeRBN+ZZDP+QTVpW7l9t47L
FRygaZ0yZPiVtE3LIZS+o4gXv/pFzb7fSPrDoNZi7GYEuSR+fEvtH9D5r22O2/0b
Z3bIh2Me1adagg1RTsA/TvMViWU8z6+4AixT6mP0Op7gBLfLU/tB3hHr2l9voz7W
z/AnQBaHDjFw+n9Dqbi38jll2+T0bgq2JVJ5dDSeTJy+ST3BD5xtCjXgrue8woH7
Xhx4dcr2ZK0pRrGuZAOfl+auB0DF8LBWkWo9Mq5zqFloUX/Mt84TtteJHplwiheS
TW0LZMtqlm0Ls1W4Fa0O2PRfKwf2Z3Q9p/A7FC6dGAEcGwoGX4tFhLMpo9vbTu56
IrsQhQuaMGPQa4LBM+I1seMQlMgojk33D7ICyZFzMjm/YRbZMD+4FuuEE7GSS0Ya
5tPKKHacVETah6QsF4xNc9pNKfZwS+yxWhsOppmgnhWm7z17KFzzdFSaVvjqmWHn
e25Q6jKpcOUM/4UOnpiy63/4omE3S7eH2yubprNf42EIwzu+GB6KqjmrDgnmRx2m
yw4pbC2y2tD5+s4f4xepZ8jwtWirQmk6T7XgSG+R8HFF7a1PxXtP1/Y0bPJHK7pS
zBiPOYp3V7hx4DTA6CWlWutNhGYAKL1VpO9f+9hRcdyVJOt1CPA8htssOSvLRgD/
IyUeTtWxHs+Sus2zs4wdRkBgJJPkxcnb907DNVOCfcq1Jl5TjKhUT/OgF7TqK+Rq
OmnIpNn1nsq7MqDQAwps777X2upbyA7gm5+Jwq10U9Llw3yELbtRzKXCuudJCqCF
CwU0/+aj11kwXbZJilSvRvrOJ+f9MoWQxMxPSJKV1knNRjCc6uQpcjNu6fx3vI0e
msbr+vUG01wKv2/7WpJrM8KAOZfH2g/nFfwYBAIXCfAJCFeIKCa6B+ziWDOsb91Z
BbwBxs0gP8IH6Ix8xzABr9mbfAxfg3KNmhoISD1kxyqB3j6pTrc1pd2k3o6n1DfC
hEumC0yLMrr2Oti5PUSgt+D9DNQjZ1fDytn8ICmYmmwce0o0PvyPJX106Pt2XLJc
5HwquJk6guJh1F2U8vwdQr0bI1lx36lHGu2POHMEFoV5ilBP55Daq2csQGqFaxFy
x83hSb3EDY5qzrmWHK2CBl5pBj5zi/+CX2IEATbm211/nOj8qc7voqEO6q8O2AYn
ikGG/qPof8lyJLWpNMA03LCpvZb1FHwXmEArJ3COHANiWFPNViO4QJtdQoqz8f3T
H5QvWJw5i0TebPQNc5yXboHVbGWJvqBFHHuBq0obBZCvrLQUl/ph3NmO9WUclNGF
GBdby4D6Uo3mWTWD5nlrpfWMcGm8ipzqTU903XLJyZf/FXsa44m/yTG/43b/mvgX
3V7TKd+8zlvAB0tSh5O3K0mVcjBzfvgaco7uCr0kr7YKkMcdP9AIMUzYBOOcuRTF
NSmsNnFZwdBFSwLDAFE6dNNwvgTXbNjDKM23/kRVdpfuxJS8WGjUXp9vwzkMexuZ
lbNjz1Fig3OZlN3MpZuxFyFwyQw8sGYXGBetaPUVNimYAu+jw3mxPhds+IU2Beqz
v9Kjyl/niZD/0ebJUzrR7ZTGmd/sRYjidiuGsaogJzZlUG90tDq5eg9MIARqXwEn
MjjCwcHPRHB5mIlFizi5GEW8xerXhgWvnLdJZoCD4/JpfjkkNrKlZvdx8e8Z4HmU
JcpDxixUI7mu6vlFVsm+eG+bPaGtZQSi96YJYmRUxsJjI8XSUgbLSidqHSQ5lPkc
4GStGSs8860RJHl4jVJVuaqoHcC0blz7nVSYnie7UIF9oOdPlUdum595ntzrVCOA
lsPWhoW15BTlyePv5ZQkOMr283dcKcSED17Synq0pkxlExqqvP3NHNRAfQknt2GY
tfpIQqv6slfDBVcZSeR6W6PCxp3x4uQL+Huytwd0s2xo4OIIXo2OK/8kqEDeMXqe
wHRPC4Ji+u6vHRQdM0QQJ9WsBfkjqT/efftXr3g04ahdrC6VT+AomoXFFmSvqqOl
pcjcHC44pYlPlOaMTT4KDo9iigd/byYpzsNnl5IfG5VqY0mrYA1FenyudqavZ+tz
NItYW+tGvXOgvtTVihIXrbw9ffgDr1G9RLxkNPJzW7QSCFmf7AMQZIP4NNJTT2sM
1B+PpHgbPk6f1gCWZ9zIs/qcQi+so0P/eDK9vynR0oyf0NhXFJaeQdFUCO8Mn0yg
mH2hgLDSE8K4CwQhUhdoQPoHJgcRVMq64WCnb0Rm9Wr9NFYaJfpt+FjGNvj2X3lG
Ck7RIHWyFLre5xi2V7AOqFU4DcMHpxYxRPcNWScUGxoJZxa/0KZSRCkjtQ6F5Vge
9NdSoxxSNtbEAiTOvLwMjxPzQpB2uhCmg0IB4Yv6Hc2dsc7IB1vQ19JVPOJtQ31F
xVFcklbueXsETkA32icTB6FvS1S8aA9bqDOv9/9gS7nzXaDL5zorMg7+wCOJU8+k
z2jwekkdXS8NRYkeZHIrX9YhASawv/Lb7DUE7GFVZU9dPCeyb2MRFskh7AIn53zz
S0vFPB4JnDkNy96wV1RadearLdGfZIK1Oiz0KR02Uift1pieWd5+LPLR2GqSmgBY
GMXnXvkM2y7nRaSwNtPyQCPMPFUHZWQv6jxVlCGHzhiU6YczVnZaTHciq8Sj+KW+
ZUdmHkbpgiYjQfST+ejta6nBpPXuzKGSHMDgnuWneg433Jqbxii7rt90vXqQvWj4
fX7UT7g+FR69rU9/wf7IL5j/dPKEEFmg3/DCyfrq8Ubjgifh+A4eEdulgAWI3Osg
Mqwtpp+gaT3UUEaFbiZMFU5Sh3bJD/2ZYyXF72WNNfEqPeCyMzvAFCWiw/Qf+bKn
vFuprt+EbdA1Wg7vPAvGux3tz5QEUxgpFn4HJdxaymKe+rBpQDWbqrwg5Zg3BxHy
ZFh9k9EQ41c0u6GwTeBm2PDZW0o4x7+rCKtGG5K0hIQ63bhIEy+N0EpImVar1l4I
NRGCCsujoCmgQ14Wpxavuyltp7r5xj2h3VTCCBXdbUA4Rp+03ZgZNShOYZ0lArI1
8bu4sAZrdGWThHcgpX4A/RlQOCvddpAOrV7p9CgHfi9maxKm0hma0XxSoSgET0dV
G+D256kXePO9f7cQEhtSx+LP0cglwGkQxjvPdh4ErbsFhAx7jaZ8848SRa4eKNF9
0xR654nHZi+zSCohA0EMFtACPOG+E9dliym2NLfw7coSkkYL7sG7VHBrawnIT+Hp
iL1yF3AJ++ZHGTyz2g5B2tM7YBtieK0TWvfBQIgw/E93mNM8upkKyCxWcQ4ZDoN5
rtBXpz/nGv/6BjjivEoXn8clmi/j+nN+V77gboHEFQ8L8DaOiwEfQ8Oh/0nHVKPz
9gOdHKK29ii+i9ZMmMOQxCDKuDIWGz5l3JkeefSpYl3YYQpt2Nc5vQgBHAQCDPgx
8P7mixLwNGkdNq/DsrOfis2XxzfKVSfV672kRt8Vtp8m1tYon6u4ua3DGnGF9g1x
h2oDVEGTUDqyxZD2ry657KlJcccR+8eG6T1d/ZKAHDRoTeBlnE05C1oJL3d7kOFj
a39yLbt2CEfbvgLfay7UAjs67sanNxDE5rHFFQYMIGakXSikwo6ZM5iFRJA6T5EX
yoQASJtrwTiD74V9gHogJW27xwhqeobS24tM4OGMJDEGXnSuhFcnpUm7+HDlxohA
skedsLDplEJ/2lFAg99iJWYhNf6v3RZS13GrisPcL60bcn7jifZw+zPEl/3YFhjN
VfWgdXasIkTRT5ljEKAqoCp76qOAKPrABYgnHYgS1yFzklUEEtBG3akPNlGqU1yD
A3QRtov8VgnQi+179IbIGKpgBxFwHRD76UAzc30vul781fjwHDWqQYlsqcOXjr0Y
6FwMbLONO+AfCbZuYtON5VtCUn9jhJo3Xxg/MRL2rYPmMQyBN4nUDZ+msfQxq5+2
nnvV98vXnfGdgxAuBibrLnIBMDOzWdA90ibXLTLe0om66H1fwH4+K7BOfd0GpJzd
/OdXKddv61wHvGfXdms4nWjTMh0fQk62Us8N7fvHW94CnCh4VspskWii/+GEdU9C
ZDa4ccf8z4vktv5RSi65X6iMdCtVdybHXlAzL/FqQkXBrvSucPVOT7eqr1nHqtMx
thp6K5rNi3oQOCePsYdpeVpJUD/g0WCPsFXZl5QIpVaL2Kd5sbUeh6ARltLBD0QR
IY4p7TYxzmoZXGpexysSXeBWHQTy3kP5WGpbUEwmkMcUtwWLV3PKHO+Y4B9/WvbP
qEK3K9Lt7dHla5o2lBL24KsL9wyU3yncO0atFQPGW801FMOTSaLOYwEYqzJI1gcp
0ZfBsjlTHDyp0kziS9d4tDZThley4USPeI8NeJsegLkSluK43/infaq93Cii9vJ5
LuN3oZYLLsUqqkdHgjx3Xldn4ErAAGJ8MkUxLwk6NdZUqxf51VEyHPsbtxAa1IJO
kVN8vDVI5aLXEsSkqOzEeTLruSlkqI0yw/j7uyv0rM5130h98CFPvv2Q+QA/v6Aw
ufo2GedgKR7A+sd6T4EkQyUGRoBdsrg6buaMxb+joDgvB/rm2o1yqBiOQkoTgtm3
aB57B/fNIEr1iZQhFE0gxN9GB92nIBri91wZ5qZC8jjW5cUDb7ImWiILemA+Za2p
bjpkTDDxyMD4s34xjn7LbHiTmIiD1NMofUhewIFTi1+rjjD2GhWusZ12d/6sSbQ3
YKsZCfvh/q9+8dOpAHXCpGSgMfxFxDgbeW9CdnQXJNjEt8wgZUW4eU5aWVaJZ9hh
Pao/P5TIK+URq5HbeDHjsn9K9qRP33TNx0r+a67Uf5JhneQEFr1Q4x8RnBaxFIZ2
4DCwr9B5GKL4gH+/NGMfsU2gDXMqSrONH8gTGojeHKvyFMkjwSs9gYIr/nBsOq9D
bx756RhtgVf+ml/e7pQk/EubgwGfpxjlHrYArfvjrSZX9k+CKMuDKfcxnKLSUv0p
MpUCXQx8jZzdv6pJ1ohj12hR6D+FlGO9lzCNttoQFbzpbK31S4+0ZFgg3iPtUlTC
EuwNUdadIF8mg1bikB4ewrzU0RecFIA1u6gyWA6r4sgjpiclTi0c7zC9LtWRpr/Y
ngkp4bSyoGRHEkjIcfXc9d7IoWkci719pvg5KOTClYD9PNSE7PBtYPXOIFRIN60N
jgu5W+h/bsLBvs2SRrZqDd3PTerpRnep2nDVhN4VFwpfonyglbPFEJQ11o78MbhI
5hocDP1drbMSm+acoHQut/VcP3gqqKX31/ZyAzY1zMb67XflQb3Fw1S68sBNvVln
qpyzO87s6sMHxgyQ8/kkIJG4F411Zmkl6azZxz705SzKjjhWGPm1PS4x9eDGI0pE
Lixj4tYMXhQE2xAcgR3k1oAJLBM+KMia7xX2grGbdk1AXRhlUvE4O0MY3ZZsPqdG
4CnLMNTWrspPuvH1z19aDEgU7NR61ojswiBkiwJisc1TEZRDfYalvM9pHEEP/p8V
61kyhhP+QrUNgsjQtPlT2PmP+j924gyVQexCCEWlQzRdwtaAj2d3J3ulP2kQQo4+
aFtebPYWkx5FiiblypAQ1xIBJudV5Hor7rV+LtOp0PRDbEj6Ezp6d38nwxZJKEAY
S6u5D/16eCqzsp52VDIyCj+XaioN+xeEomIYd0+m3baAE7V5uJJOcdUdUQT/iTKY
u/ibIJgW0bq47vwg56RwxZyvKXQx5uV0Y9VA4natU2KDtrian8Ca8eB2znp7uSBV
JlrsPlKNHMXDbQPdo1Jfuhhq1dx94K8gtmykYhPFZmR/4FIzeesXX8a+ACPutcqD
2go5FHt9PhdWgSrsQ1ml2ho1P+OEzgFsBZ0mfpZRY0thzj3wkNKTdidMGYGj4Uxq
yUpKQZQJLFkF8R5hBwdmHj6qy+HciT0n9vDgHyUhmWyClPn08YRVAvDo8ODhJ5g4
TXVd//r+EWAHz/1ZhtcMWUraU9yegh7lhjF6nx5z+e5BSt7lu8WTlnEcKFwfzysK
TRJb0VQ6CYvmhLiGLw/e2wyMW9ZN5ITGw73nDHhKiprnNzbKpCAYkL8l8RiIqW0N
UtMpGi9rPqFcJoN4pAoCgaZYmyemOwOKNfxPtSIpjRTaI613KGR7x+qtcwFgswBo
VH1qXTcvu1SxjBviwgUWMEwlwiUSk9fv68fmbv/m+nissmKWPT76n/Z3ZHyz9ZQk
/tvrNjzK71N8qO0i3lHf7XeMR3NpMD0u1tfMOpi5dd1/pcJ7OGGrKkG/Te4hCiuw
Phr23urQV5NQPSUWDx0sPcyKKNkTfATVQ7lV4wG4VAroQ+r0j7/AgLbTWJo6U0qL
DVOxRG0hJ2nFFDvPCAR2O1nXeK2YH/3sdDqB9rpS+cqEtno1xloFP0lLkgDrF79K
6mJlCEfzl8zCukrILXBhi88sy4NN7dgYl3d/n0T3rJc2JRfOBsonHa1iZKHeHD26
g0JvCBAyyS2aCPuBZs4pVRCegiTtfqNgttiPrtH6zNRb+mOXf6ST1nqMJinwsavu
keNHXbVszFh48apI9CWQLg4x/kLPa0iYFl6H9q7Yt7TFkzsa93+VbQJbPIqGouCB
A11uLxImU/XysczcQjoWsPnQhSrDupjv59qbr0GsBUqnkFnsp2jdCH7NOxod6A8V
7FdPVUF8t+VYX6zGzoWyeIGwA9T8vE8KATR9aAcKVSbpAQPvxP7MCj1FbQ51Jfgb
kJ+5QkUjy+8IfPHUpbvnDnuJc5h3IzZL5jZaDj/pCxrhy9HWMrn6zuX1pkVpdTsS
UcQJ4xL0tp87CmkXKOEhIjc2YspRqTA4Cqx3bP0VvF3ipLw3KUkVwC0ydNfUWNv3
G0dQBJTnkCBf/sfGzbqk+ufZFqcjWshUkm3WLhMzy6nh5cSLwb03sOV+7jAbVWCY
9nIolVw5kylzS8go30HoGk8aAVBYUD1Y0+J3NTjRktEWwuRTY8wd/6GnWNfPnN9h
nu0f73gWO3/HOvpFIiv7u6dmeUtjrAYhBKj26jGp4gNBphfVtxwOGkN0N/xou34b
NLe9aAWCpPgXkkfctcoBdguVKXhnP9MpIuO+M08t1gR59wL3SmDkV6OMTf1rPphX
rQTKbhzWVmjshUFG7RfBiY/lN4vHzip5ozTs8NV1wkseP7eNwOdeczkd7ofNLLTx
4re2wwBQJWURFMdKizprjkg+9veBt9A9qgmUu8BIW49hzvYg610D5+MbGmJUU5po
b314xbpxNGqhL2PCsYHqCTJamGM9+k6a1dSmPG7JbuS5V2J2Aj1kaIKYNqkpEKxW
4rLKn3W5bY3jVx++P7cwzoRqes/YvWxs4pxqDp/C0qL2WsleRXNcGNR+o7Xd7ak6
EA0bvP/8J2xYx2EODmLDuFMla5ZFBGKk6rqIC3E/Y8WCLYR/QF2nUpu4mCG65Z6f
17MsgQ7angK+xM+6qyLI60Q0kxl2DDjer/BV7LeXIHSXvFLRtwUeXCNLH/TJGQnh
nJohi1VkQzzjxD7PXh/Jikv0Ay7wleDEqCVA5xGCd6oSS5FOyuu7CTygTrEvjpGK
c4VLES6nJqfQIO10/BUR3uEgJ3Vj7QwP3RBYiTM11BAMJ6gih3t23wvj5Jek1J7m
JMsHdfelF/znwkYyxoZxaUQQJROP3EVEVeATZLIEz9gd2CVAgw+6PcrckoikbgSi
gL2K/gpJAGBcLR1rscThJ9lENdq0VSpB6IVlQzU7Bqjuf2Bdwvx8D8eA5nE0IUOA
cSLID9UizNyqOWekVA4Df5zIujwyEk7M7lEcoh8/gVtShxh2EXEL2evL88pyiQFk
u2rP4zDUlIcVkjTHunKav5V2PAOCrI6OoZrcgffglwDouVpmNSem5PIIAueLmimY
h22eDr1JflxkRggzhLODNzBfwuWhzzNQEojLlJVG6v70BwBp6DBdGVnILTQDfcON
q45l+KoWQeL5qjnNO/AY1sSJ1BqcMKi2w41KiEgc2PIvg+gAuuspURjpmx8Iu2Sn
dj3/hdtUaF5yBNkVRKLRMOmI0nGDNnkTXwHy2zo83B/oZeVTBbRevS1BF/wC/dlo
Gww4W3LXkFSiSgc8F6793NN/MMZXaAqDV1HtXeAt6s7gVy6HASWH4Xpgv4tjJkzl
QkrVbBrtM9O4JChpyeXFwJFGnepTK0AycUrM5WsQxo+UNygyjn8udfNLJhyMZvWW
n9F1A6Z3iS2JVa1uXTmVCYZmCjvD62Y+IBP9cuJtzFyy2OHA1QWE8LQzfVqD4GN0
MiHotXkJUAnrdL4Jnblde8vP+wKUpKuLmPWj+pWURMAZfrOyvgMiYrBgk8mdSVmF
9aVg0pQTcmMKJ+TZf62N9ox364Q9SlUzBuDtWvaYMrvndOuXtVd+HR4Pm56yqd7+
1mvyss8bnZj+rmnAZ83tkBQyUKZgoSfepMEj24glqpLv/vZHRG/FkeDV3xjY9j5c
gp2+R+sjNnpcRPSYbyhV88EUk8PghTiVUtaFjrTffOdxQFyZhfIt+WgF6yBELT81
iOndw/JhAoPPBhFkMkg/yB/wKh9B/sgVyce64uceFXEry/kBWOZzb+9wb8UoG8AI
Hn63goj1E4Vk5hgTlq+fzXLvhjOA2iPHg3WaO3zjuNy6a7xpX03jEy12cceBICDr
2C1to+Sbqy6H2PRF6k6hGtFKtaZSQr9twhs5E8Bq+yLGXZQqG+uU0Ob2AMnjruwn
lQRLpTFV8UaSiT7CHrF95A83pkCMaqi/JfOcQEE5hzyoX389b77tpwmM96IzCeTH
qALcxNG5xEiyRB/VfQGosVh66M4LtTa0QahdUjp78XJKhJfFLMSffL/rKtgMO7B/
SUhdwcRmEwvu3x6Emze1Du/NB2sefSeOR/PSwX4H6VGuCbNEG+gQgkaymXip61xD
AjEjz7jWiB6AJOkM5cWcvm91/xzXM+lULyU63Ln9e3TeC61sdW7zUkmhBivtIpFf
3DtMiYi+Iygs8y1xQMF6N4vh2p6dXttquQ/EmQ/wN/hPsRvsdLnYEzyji+I3Q3Y+
D1n7STqX8QtQ6MuOs5MXln52oThiwKozKluiUxCUGX4YuFkL+3QU9klrwSOb9z7V
dH55/IuKRA3GxoXzAmse1i11mAo92euMn4i5leB8xUDzyZVVqW4BXpsnAnDRse8H
RECz3gpYxMff4fEHS3BfoBFLNdwzFG6HRmQ1kKBu5WP8hAUT/Z6EkGF03mSgUa2f
/MfYaSqLq90+Vt8kid1OokJBr+IoV5E0LRUENx1yKrMF7YjinadBJW+6xws76+ki
HgDtlMgm2DIgFQCj3vo5m30kpVygnV/lvE+C9xZbSzHmbiYUgJvmlv86lh+24kgV
KxW084x6fJmmgDS0zJkwPlNU+KxqbA0OG9LijMtMDMyqii6As1TdnYJ2NcMKNt09
agu0V5hGHL3ADaTTl7t3LI4GDkGYaWULY8W5cfy1x4jqGSk91CBYQoY8x4/kgGdF
vRc54AgkS4JAovwr0hs87NoGd4BGtROeQZf9UNTVkO+QMZO9dtkl0r4IXsCA/+oH
+XSSu85BPAyEXcedFu3WagHfH6XiRb5kuGD4klfbEXIMVGWF/nKbzLtbEMSSQZY8
wMge4GgZ6feYIuVgYZNrTvhjzjxCyqNqZgG1AVD0cOUpmCjBCaDPRn1EsfJPf46s
8ymc1czSYQVrSnCWcBimp6ZiR9H4Ec4faV0GES/cCPBSsUUffKZLWK2X0mFq8ula
vjKvaT/VxpYUCscOl5HlV+prFc67P2ymuEzsCd3BJUU0Hxdsp8rL8QqmcYiTs7Nw
srD7G1mK9WPFAk6zLDZGOmmDJaW5Lo5/vGSfE/CwwZOAtztAf7fw3+286UbjVa6P
aeK0ZFWC/YC/VLDfBLjyjpwYSQASFurrmnKQ5yJHqfVpDh7fLztzufZJnUx+Onfv
C3S7t6J9OUIftZIeLwrERb1rXUTMqnJuFOHj0w6d/qlS3sDGWYX3BQ23LBha/4s8
WYh0Ct4wFSZTv97C4zSGTaKbCr9MwtX3XyK6mcKMnXR8nRATG5bX6Dj+emrq38YD
TDVel4YQrxGJslqYPLZroqn56fTpbFf78n6o66JtG8pOVKg7zBFVOXqEPZqM8X0s
2DFEmDiSFqL8VCfpMc5b1jvZISSmiIz0EgNAPWot1TLbLbz2oH2FaRDrXDHuxdD9
fu3pUQH8Yo9TTnpBvU2UdXhZVYdnf4iyX+tYq6l01AUdwdHRiJ1Q8DZHNMmmK2mt
KXdgwRceXhSEVYmuXhqd6SGUPIoxRG2oqDFRGxShW52g8KkyW2pB0ak9kigbSKLH
WMniBnb6/8luIu0G4CPimNszQsmKAeh4FuEGhIoG4/58P71ieB6+2Xl5n20+64XP
rlziOttR1Uk4wgoBCQuykFN9a3fCuVlepfuvVCkMAymFg6Aqu1UwAyk9HI5FXyS2
CrtI1LdxnIz44wKurPWv+p76h5KEysQK9AjXpXgLh3/qSWEQrNLshxMxCGMmp7PO
67eyDrshVarED+Fh4TddYVq3tKhyLYJVpxYe8zPDL/X6UHCdcpuPlgy6Ypn8yc5q
gHqaQkIB1YnnvnGgknE5ggNWOcFpxLK1r13LqoumYJ/5T6OQ+qFatb5wNxE1Ygtj
IvFxFQKFbNQYK1Qbp+kFGXpQDkKvVxsXBocBBadsQy7I8LmaJTBLEg26jB7gEla+
k4veIVcHsKiDsqz2FJfmjy2ayFxWiF5uyjiGOQep1nx400haadXftwib/BY2GzkY
9F/Q6E1O1LfQJFr6t8IABo58Mj5qVH5lIXHVhsU4xU0PGuAzGhjD+g8IaRQAoBM5
VrfmVaD4lASqqckJat/3CT3w3qfZKern3ikYx2R7MuurtdojD6WoQyZN8pdlK/92
REgJmyaeKu+jDBoupJSsIxojxE/ZtLWFpeKMsaQK1/QxDAHNDbNCx10cExWyLxBs
v+AYJaQPj+7zDwqhSqDYvYEAhM+DpJbEac3MiQ1tJScg6Mq6W26qradPJYaSy4Fz
xSeBEcqTov8ne7YBHZViH7hF00rP96WlB0/hPU3EBB1tHZsU8Bgd7mWRD3nbB5MA
IpdUnqs5+ThR0ylz4YehyhVRZem4kiDJ3OTmufFOOIkpO3tE2OQeYbUe4Vd+jYkZ
E9t85yqfZg/raDReqqKJczgKyDcMw4XV7OZRyDnkrWkSYnoWp+06GMMNT9k/UoSA
FeyXRoIIGi3FlY91MlJr9XJ6JuYap55mFJi6Unttf+JQPl1dBjJfgHZOuNdlziak
s75PvtmhdeJfnyk6a6HdQU1ntH8cHT6XXqjbfWN76L9MhlPGAwwaC91jeYgUVKqj
xVwN2B+1paIUgC/51vUNdk8Qq3KqZMnVpAv9jkuA7IKuQTG5l/0G8R0+NN2K6GMb
K6hjpbcmctM5juhRgG+VKZyKdrnF/g/tphHjchp+YLPWg6ZjVx/ur7m4mZzkWb80
sg25++rIUiLEQE9GeScG6dMDH571UFfO8xuMBQ5pF2Id4to7pBM9sO571hurLFf2
hwF0epvGJ1IV6nM6E2NUPzR+eD3VqoEoqvBEuysmkNr/1jE6feL3ldENCCkAka3W
XzUILqQLdv0PBSmIrOLbreRHlJKfNecRiejhk+/sx5sITXACMzm7c1FRIrxpc2nB
jeQp239E51dUOsDEiNa8WmPgzbfPRydKh0qlobkyyjKmZcxC6QsH/w0i29JyCqDg
KLAg1cl7NQLpJP+mWEPGdXUrY4H8QipOx+b2WzxXPCn8kN2leFjVwJb66gXwpLs9
cez9oQPJIPLfcj8dT37tJbkVW8S1SUym0dU6mU6Y6In5Jpnpu34m5EgmRZpGWMsQ
oM/o6T8ytvRfmtzJIML0KMHs3BWH/ctP6UsRyFM05/fLjVOOE517yIX6bHideLU9
PkA1K45o5rDuJ2cMGdxPsm7ooTbs8RvTvF1FjnofOW2EbNP/h2oVqqgHhXVU9IG2
d99l8RdPawoDRzypFIvyLo6hBr1S/y23UiqaIYQkMg3vKWGJD1GoPQX6YZa+XaLp
2EMBn5WIF++Sm6qokSCRuttr/kz2Pm12Dzez2Z0Ok9yoHakk5++1L8l4vfXzpUHX
p6kytuRYRwKtE2oGKGWCxQTwphbdHxnnEDnVD7KfO+vXAc51M7Mayf4PIaBD+zHN
1SHHmNsPmH0UY/+QY3J4nDmxGllb1D3yHmvz/5078wnoxAa0su6e8cIbfGYy6BTc
4ksZMR71ISWQqjVw261pTAygrwBBcOzObKlSIj8Q6/o13B78TUr9xYHtHg3IWbfM
0GA5DSlPLXzqxb7xdBhh4RAgOkqGEs9jy4cK2+AKgp1PUZpE7YH7NhVTNFcYqDyz
Ygv7WI1yByxBJujbtGXp3LWNqPerdp2kQuu0Pq6FlXd2QJmFbO2n5Ed1q/agqyUE
drj8+U+axUKwYSESogxxa9t8zZZZ+5EwLhAKTTfvYG6HDcRm1/8mA9cRbDZe+EX5
kPCvdt8ySsOjDAh2W61A6lZuDhGlGeITEZobl65K1/yzgaEy9LzuUfnT4XKze9XV
KWoShK0sA1SCqA9/jCf2zE0nzELGKVDX2Op0B4vn3ls6uVZ98pSslO6NQYVVw+eB
oLLpjd0NlyozYSsapkV0b/fZCHMifOn/HEUMWVW8I+ocL8sBZTQtyNoqHD8t2q1n
Ja7FZfxxBmozDNzO0BRqJUt3z4+XuFYU8nclRfUEu06j7T6dctkTo78jYCOW35Mc
d5DHqZHQwAy+yUsbaadiiWBSkCbS6+n5aiTVEFMlop3c2ohLc+x3VYo5ZSpMSOd6
D0ZeujF2wrRJwpml6mfxhbxU39g1HYpVvzczIzOux06ra3YHjxUEioJW4ZUviErH
QH3AZN1jK0iSM4076I0syLtbkUfdFIssgRczN0OU1z5wXT8yDoAwo4ySLsDjc7VY
slbFSlLL9EaI2GvqqIO8zxuwNXZwMDuVkbsleEytKHQKQYSci3WH8EzV+WIlPTYC
v4kK7wEibR36+nQQtlp9/kLC7LCnht7zUg/Ldz+2dRCp0gBqwl79O2qYMl1DX09W
zKV4/+7lk13x4PmbfeeUqTahOsqofpVXwMRuLILq0PGcPSJWv1guH6yWH+GwZCVK
ymQPClsrKmAG4YoGvgvumnKyt5nHPRDIGtl9amevI4kaDGAM/YT4DYGN4VlTACHC
jn1PBpuRk8TFIlUMqTKaJsCfwf8UuAuLSLlOrJ0rW4M7YC+UaSWzn3Gb2ykWv/5B
qu5Bn2PEExhooFnUkTt07Q/n7Ntf2T9VN52KD5L3v1BOAR6e4sxQs2g6oKfeqqor
+tNd3uPI8YsiV/95zD+Q7cbqwHkBiVe6HHgtATcrP+dnebG7MIOQ6knrNl0K5Non
41sN6/qj3lV3/uNa09d5KT8NQVzikEn9ewgtRQ5L9vAjrCfD+5Vg8NeyPj8jgK2v
YLriR08+LTvrh6eC2lwYft3xr3LYjsW1+KRFMKy6yq2Ff+lLQ+ZT1BzoHDJMyXOI
UdUvP00DNvMN1J8E0BuEqbGA5hiaWNqcyEOMpgF3Tfm9SxPVeRpknTwI72VXmQXd
pSKpkkDICsRUy9qs2vzAZU9w/axfS7Z6+GDLg58Fi1FromCjsbnFsnTixGy7xO3j
y53bg5S22D6IkkMFuoN+khktmYCZIs+sTCOxF/REnrT+XVDLwbBLd7UzYjCcIt9t
Ph2hchzw8j6ESqcPyAt18Qr8x6RPbarVTe6Nye7G9G5eHK4IMgcSKDjXuSjBXgnJ
a4xnCfnz1jVIkRTyeRfVDrWb8m+Gb8U92W5fSO4RdqbkSdSbrQJAyz8R5lvX8T4T
Cer0jhBTUIHt7CFV/EHwdLqXz5gQQzoAZOP4+X9TYQi9iqzVxb4FwDsOXdY0/Kbv
szaCva0sJV6DNka7uXuzV6KPpFnXJG3lVbHBrop6M9i0iSTNvfOvFcdrXgr2cQ82
CESxZKa1Vjw1/lYGDOjO3LL1m8dzujPVJreLJa+TLxGbTw7j8irG+ulf0A1YBeqT
SjYT4WAH+EqqMa1NEVq0NQBYBwxGP2GQEMWRnlp4GsfOvslzpe0ZsYFyiWD8tXij
Fr4i9mOBXuLc3w7KiTHvxbMBfcg2dcBGLQnNAwtxx23YSXHPQ26h6SC+TizEfiHd
3UZYnOl0BEeLy9ms0du4TolPOwytrkRPdjkQ57SGR5iXMKeTXOv699LYJBETS8M2
BdrJYuUa8D5UDDuv+hVuOtBw6gOGnUFCIGEqWK3s4w6GATO9txJHx5zD/JDe8IlR
FjIjeKS27oH9ikRP0SfRXfrAvjxhJjHDpthU6AHatyt2KcskFPhmlrUwKxg/2a66
yvLBB8T3wYNV9VNwcTmawsHV+bIvAyQ5Dasj8TTheBKe0IX7s7l7n1yn8YC/rka7
d48PhncSRq1nfRtWBvAcBEwdjOwULWYYGxMR7chQOlJvc1P/OizZhlQN0AAUAdYI
5L+BwAVaBH5qoq57fMdjVw8Rd52aVywvBB+J0BNSdY9euJhUdfM9yuNQaiuBC/T5
n5gqZg/WM8yumRdt4L+JiKnF2kGFdSxWtgDMGXSWNWutUYdqLgG3yj8EY7GTmgdZ
KYEwQDHOD+onNPIPB03S+YD9UuqPe3U+Men2OgwZiVT9vgRgTOsN4Rv52gMXVMcl
U2Jtn4AbhZb6IWcNziqMAVUYS8fQXm3Xg/1z6yVFThq0hURdMob/6wlHxuRFayoT
VIIqY8J6lRdclua8JG94JvfWch2h0IrkjsbHOrNtl9AomlPNLGImrpmgb8jrEvYu
D+x2DH9DnF9yk1R7gKcXAw6Tl/7zZX+KvmY2B1LhYamVpoguyNjZzxL3Kq62wIkG
LR6MZVWpy6Satsg/cAVlPIXZ3aYexP/vrj6h4nrfgysZywwMqJgjFlv+nNAGamwI
k+uYPKSmujAWuUsDr3aopEtf0c3ghxcrAlJN+XMfJij69aiDdLOrK+2s9X0k9yPJ
qJcq77p682MLerjNE8rNkK6JKY4hj6dxlHfTudXMvE39KhJU7cgAmHyydQm281sW
TCAkouY59IrF5PDc+Q9SEnYjQJBHT9TJlyB1sCRZUVUfHhSF846SOx/SL4i5JTy4
C891dm+bnkr81VVBm+5MWN6xGyD9P3S63XQeirCAIjn8M7X62vyQxXncXODc3ZqE
NFe2r8JPO9cm5FbkvCA9nYIS7X7pOV5K/nD9Ly7T0llB69a/ynKV4/dkUkbcwcXo
6gzY1m5R2JZ2bhL4VhTDcI9MnmsQp4t3FsJGt7UTS4tXfIt1ztragRA0eP1H+XzU
ppNrsEGxiaZAo74NuSvJ4vJV5iF8zzS1vIERCYN2kw9z6UJgHHMhipo3+oUAfZle
f+TTUixRzx8LlUfWFXXKYvBLiuGbiwehXXmmWJwYIr6x/NaS3a8PeJREgXin8R+J
ezUczzZxY+hlNoByQmbaJZEhF2NAiZttEk2TaQhyHBkL5vYtJHqxL4/dQN4VCr0p
CriRH/C6X2kb3mkuP5jJl4yCUPN687UqRo93fxqpKG25Q88AxBaGsEwZWMOgwAi7
u2TTD1H1OkQ+y+oYtfGtlv0SDXXOdb0Fa3tcrEeBqWuRybCB9Oow/fxO7Ql5N2iE
oOOdGzPQgikUbHrmjpNVFGYDpqTXhbPkgX/40z2DmA/6aZ8qT+yTsBbzE6pPfuJu
L1VQt2AkeqcVHS02oaePIiUUNe4A3mXXzwd7wH0lJCixfYmIyFeysFCQ70In0CJp
Zv2stS1dU7p7VVcCufJoIap35DHMN4bEcWfgjv3Ntp+Y7/Hr6Ae/K6Axz00Oam+6
Gx3FENz+qEJQw4mqoBlhDTrpbdQceaNCOha79P8BiETOi1o9Eup7l87ysO+MmqyK
JNOWW+52xJpqzGOYcFAfNfM3ekLG6cmXXRx6SQcAPPhAtfSeW3yuKxrLXvZMNPov
XG0vRHFyuybTp6EuyNSe/X4tB8266xG4aqpHn9RqETaKgskhJ3Zx+P7i7QmjpD/v
at315qEccd0GVIOE5EEHDWdrQuqp058ZcSK3JMsu3MAURzX3ZklYCa4PVkopIbEX
rYPS109w95w/Pun6aozCdrSFgQn3abL8QT3SaGe7x85qck8/fv0l6LroKGleZu0o
OtcfexH/a/nqhUCRN+ACxhm7SoZ90FL8b+eCF/mR8iz0lZXoJC15QfJN4EmGEVrU
OoqYGtnn7XURmAYF6dWCk4cFtOy0avogrGbgt2zlHClhkqE/2PgRcuMpLacKOhR+
U8gAeGLtZxqu21z6XwSLFhLlKLp9KchfgH6imj9KbznHRxIYW0FWm9BLBFOxxFt5
nxZBO4geU1jzPT02xRh1xzZLY+3tlU8g/VlH8x5AGbY3Rsq9H+hTlt9AS9q8K0fq
S+hw3cuRCI/BI+iUaES5OrVH7wa8VE4glusQoHJzFxLhRjX6hl1uFwfLaSBbp5Bn
4zGIbk+k83HwQnhvAZMwSgeGJnrD0JwfokXKc8Kms1FkGyRlNGpwJNmuiI3dLDKd
JItDsxYOsze3WjsGX9TZ7YITHRUq0sLIAW0vr7a283tfGipSNL8Gtf5LfXJ4GyUq
QrxMZRKj/g7DujIPNWk5zx4GhH842qEbizAfX5JwP7GDpF9neUz3tuAxrpbeCkA9
vb7qTwQkk6ZpRoP67aE1Aj8I3m/CgrPfo7APKwywVA3/Jn5xWGIJvMdqk/b2sCDM
NXvclAaiG2So2PytFxQ8+iBLtT/Lw3QYy8PKxxP7iB16oQLbRM1hzpd5qiLC0iFC
HFeHKvk+laEZ8bsnGtsrlGB3+qrY4VXlx0vO5eFyu0Ne2KvqSwd9aVPSm2u+/AKO
pCGcu9LywgIL3r1g+Gr+xh3QlOlyWl3E3zUuphsmGylK+/Mq8jJB5N2tUoZ7Qf4g
AgZiDFdCJt0hf1tlwUSFNjQOMkghlUCP6qc9iT1/4VBZv2FTTclXprsWiAl8tBz9
EWFrz/FYQ0sFYN2t8E/F/73W3hnOWrMPFHvZNDOKIRbvTzweCmPo6UDqA/txgmn9
DNfBRCvpzGW01RBiYZeBswtZqNF/VLiMpWfur5Z6x19+bUL9JMQjwzDeDF7ziBIe
QADtbHf9CXKayc7QSC6+1jNrWx2x3qjXgKgWlW3BYpRDjZsf45iAJTICIzY4RfJ6
4dKCCkOFOojitr3uiPTRkrBz3BvBQ6muVqxDJdxsHd8b07wwtYFzwZ1l403y2vfc
IQXEbjA1xcqORinNoEsq7eQ7hWrR7EG8SEy/7mT7C8JF3jNin2krp03h38FTW2md
jyi3Lopp8AS+XvLuE2Ct0x4R7CavAZbLyra4k59/M6rgogJMVQJOcbz5/OWbriB/
VIDhB4GPjrxXL6v+kjH0phkUFkAz4VxQ5iSJThfHqRJc7L0z1dTIxIGwYjXcTMqJ
Jg6qAIa3UNASGyuoNYcU7lTBRkcRYxboiFP1Q6uY1vwCRydW9IghC9YYppqLHlbo
rz4zVYNQ0biNa9+aqRPTPaIpLg3rYRiJESU3/9E5/zCq233LXrIAS0cWaY+vuzBs
jQ7s6OMQ631SfoKjGRshmVd6PPSB7+pjNuTrvDVHN6PB0kHLJt/o3P19Isdglw05
bauOa5ug5lShTeoQFD0VLmDR9Ly95iNZ8qTg/F+ExOz3GPwHudz4JsGjEMatjess
A9OZh/jGjh0LgWVPrHspB8GRMwOP48dKprcyju7mdR8cHadrUWdxiYUV/RurK6wm
b5NMKX+4QSz8u9XMXKpRXeYGkxPLfLIyeNlIIPmUvPWZl/T593u1BJBMboTfT/N8
M1igI8d0LbP9wQzE1q6ag1TZRZ5qu/FWZOA0gpv4w3TDI1DiSC+ZG2HK+YlXXHR/
ea1X7VNZygAnQtNDfhIDuZOgKYju3Aq3bVOXmL39LnthXtqTymnfnPbn6MFsA9Gx
eOqAKEFZ3rwzbgih9nDxD7YXNAmqObwe8ZsEHUZY3E+Io4D6Hr8amsPoaf/sze+P
NeNm0t5uy1puAUKovCkEVmb6wJJYQG1xY6aQW5Ko2AKtdZpjM6j+Dp8zdaTNWH7Y
nhrubyU27pnHWSbA10QOFfbe7Hyc7zNfzE4u8FYQtgn5XhdshyMER4slcFakuDMy
rGpmsxgav8RlBQvwrWMvTQXKaT422C7zNpDaZKp0/YqIyLpWwX3JqczUQS8bqCsE
2apWr8+goTVYhXry42oZvoDuKxHsqwR0Jbm9NHnAMO/QA+j7h0CHE/niFNYlVNe9
mmgXCZxx2CKvNHqoNs1TfMc/qrt0a2/2OtGds6mDXjdNfG3I2Z0sE94pOwZpg83A
rijjzgS9RhFNjto/U6wQH2CXsAM8fwkGmFiaq8+hoCE0humfJRQo2uYxuwgCkQBm
BbK3YTTsTcHDyE/2hd10JBEw3wNCNqhlZnYi8BoN/Jkm74/AD2sQo4+kj9vWzfL+
DJ44caVCLe6exv2XkZ9rQaKLRJCuHv/uL+AUSFi6K6uiCCfza19End9XT28SPuFk
ObmRYDZMtJJRpbJjESuHmB0qy0zZ/WZb7Hqioo7CTveleXOkTpkZvjoZTg/Oxf9y
Fg3l8ypxYiQ+W2SF8exKdBOWOVdgzIlTjQCELzHvRmb1Q5EO65nHsBYeh7r2nPS6
tVmIR/gad6ZWgqsEFLh666zPfnzy13mlRj1Awjh8m7Kg7nqgDtS5uTDpXCa6FtT7
2gRqBug3gFoU51bj/mF9nh0BtNAVv9FlQdUtmOHGmH+nTiUtt2STtZohqWf/GPcu
9jlESdJMM0o8h+bOvI3YdTTRCdquc2OjLRjjAg6s9x0mleyTw+gxgnbOq+BH4TbV
CvPptua2YMz7QhNMhN1jMiisZ2Wv/t0YAp5SMGyw75kiizNLYf8tbkg1QzAggfU6
oE9XRiCdabjfeFFnbzMHrPGRipQVKNrItmKd/bw7Vo2xK58VFeBI+eiVm0fzQLoZ
96Ry3zLN5Uy17uxAo4BBs8ujMut0OfNbdJIiVFUUA5xUO7mBmPpBcSjiy8xOpldk
NDk+iYT1tmTl41IUi9YIfWLJwlgw65IvMlcbLiEf8yyZi/kWvN5ryfvcWCU7wu3V
U2BFIe45oiS7QgYAQ+daCMzVEnDlZj+agxSZnpk4Xg/fM4usQCc4JNsT6marp81/
OQVveY2gxqtgkoDYix6/Yyt/caN9VnaA4yrA4RQ6vbuNGNMtOb/Z/B1nKBUL5aOb
IhO+4QMAzEoJITYXb/42cVOWjm1Wm2QXSDy8ok/YwK00e97zZUJQWbJLrG0sP8za
/riUHQuSGXt1ZdRy51vmXu0fEooXAklE4KGgEXkn2s4gokbiB1LT9pjQ5oS4oRGY
PQ16VhhWJ4Ap/+wIP/Axbro9m7ckO63fw73mLnsf6s4M6pk0RElweBaDcI5mCkBc
CRzjtj+eGa/kLB2djf/QJHIBR5e43CqbQzn+8z2+t6KNfEkrx/j4Bh2gEC0hOR1W
SF4T+xAIJgV2+ED/4nPUR3+J2YLQbv3zFX1ROqh4Pbw4i8uwoYwHZw9IwEtpe5ZP
SMhuqpnm3t47POubqGMncTVgF4rLeLWjFFjOQ5dL2E2rAizXippBQcKlviVpEDAa
NFM7Q3fCAK0hJImbZ6RYirD61MzDwk4nZJB3hlIrG+WNdIFVXT2W1HhV7UplTZRh
o+tkqHp3paolYfffONP0NDwj/u3uINiH2QWpNcN+b/ZTYozNXav3TH5KL7VrpZay
QkTQ1VRQebGhMztNDKnbUECXjylNleatWkD3SP1DUgf7oVhNGckEfVbQM1ediFJ2
MbG6vKXoLXxg2v+M0PtddUgSmCfEhpxfu6cc6ofK6zGMGO8abcIPscNRAMlnUSoD
bQ39iVAkSEM2x/kFf0pewnDN2IP0r3woJ4vyIe4hsvjE9RUVupicqMzlXmAL6P8A
XHV9nFMEjrzhispci3Zqv0tgTCNxSmtX6sECcVQg0rQclFbqRCsTRPB4FFvEAeMl
xNP8+iC2/RrgBrkn0jwHecfqjHLAvWZmNTfeVx4xwLexEup40i1qCey/05Fe9Ju5
QaZ9wssu3tjmVdrvoeyg8TFyoCTZ57L7OKQvfdMUuPUixZL53k9ciVyJDW2D9Zvy
PoC4324hQ47u1IzZDfl4rGTWBMlCdIWvvQ0PKcNX8GCh0vZyOsZ9+STXQI8te/H5
G1ZpMaDGmgYRLpl0x8QmntaOfRzvq/tNNUiqYTg0BCehmwJ9zVMpr1yKoE7ubgF1
1DsSsIIJN+pSSQhtgDCdN/NSY+EpAmEZ6f4LPDTgQtC89sm4n+cMbKymSuHY9QcK
KonpF/cF06JVRtqJWG0/Nl32iA0qSHly6w0+6RASGOXsjws7/a71nBkr2mgtZXAm
m9OL+FQRPOt/H8+FBqYoAB7yRccNxljioNVe/XUoZRNWGf38gk5YvmTmfG+9qfqi
88GBjKFrE9b0sx/po6tmnM98Wpyzp8swe6BZK5g5qqLyeKvsRx5x1Po/jaNEGMtv
QdBNyhZhLncvjK8PERInFsT9AT9isNZ7KnY3WxWa8nBQ1e9+YjKGr61+O+2ayNwS
nh1VHgZSNFhMhl4YtBwzyvmZ8wv6o/s5d67+932tDkC8yztpEwSqCGdxiC3NZ8N+
7xCH+JExnt1L74/x2ol3M9252MZOZT2E1jHuUAYOPxos2cfpI5Akra5aGCO5Mtp8
/R9vi5KvjpWdmawD5PuCLUT15XJRPXhtDkIhN/EfUwEE1bS2NA5N9ojO5eGBSJNP
6bevNVhBiqgFf0AbwO6GZvLD0g0UvFshz7wTpG/hO8rk+gUBBSXJF+1UHPAl3CdO
o1+KePlwz9oI+7me4SXo4nOpoaO8vS95lNDLyJ6zTTE8IpP+DxmcVTAYbC09r2eS
XQEZ1f7NUG2g/Ly6qPvF7SRCEDQVF3LM5sR7Mj8q2hLaKt+C9WitIXefK2bgOp8O
9TZZsnF+YLl777wE1ydA6fGgHat9dygFuVUtiuuEqGpzmxVKrf+sVqMcOwOBHnZ4
sYzpfrSXQgbtonvsJXW7uk4li7TTpyc2sS6Gx8H2pPjLYPPadL0thdjd7aRpTovt
COlmj+zGu36ShjaX5CVZO5+kGoqhdzQYdnUYokq620mFbxeY7dUuKAsnV8CzTWW1
d01tzIH71j1vtAKirV+mO5ZGtHWKbo5cmiSTv6PLFpLCcTjFWjdZaKOViRR8P82b
FlSsqFOK6eUIRJe+DNvnsTxS71E8TA3iBT7VAi6cyOZL+Hcip5lmzAfHcAUPjW8O
dxPzbkuG12Kqe5l2hITDA4afJeIrxJ4jaj+B347OTRpHFaUhhcscWDOjjwU2/uvo
EqGR9HLtQ8Hde2+AnQWwtCSJKUdOFsS8AvaXFO9VjyJ2A1QMNLVWgiaUk47vZRHk
HtUubMmrb9nyO9wSiaiF2WPk8RSUNra5AKo1V+EchPbz5tn99WretdtUXaynQfgH
JKiA/60DGZWAGDR5nsg3Qzau8PV68Ka8UhRh5u0rpHaauEq66MRoLmyB6waMRD4u
pR1gMKZQ3ZPP/G3fbImuduIRWL+nC82vJs/GakByMMz1jpgu3Zi3n4OIKgnN17Mr
2YWfvUp1gzoBXZZahvR78knxo9nLyG6HSgtKY4YQY6TEYfk9uvMFlWeY8tujv5zv
2SBuYLGbZnk7LbWlLCTmmgp2dP5fO5ogv+GnsXv0YN8RV8dqljkzEhaQ+xrW98SW
LPgxZwku5K25oZL31CE61fhYXv7PecRxTCRJCf+D0pYOV+H6UdLYaulQNklShOaA
DT8eTijwjI2oIPjqdYzGqLIr3YlJKbo28xUN1/JWWE4k/nMbPhTC/IPJqFTqCQrx
aqQsdhUmtZ2Vj1KzykIX0eiONB2bJzd0kf/c6UQM1E9D06jeZ35RCat7jhkHa4VC
pWPom2dX3UVJ6foHuZIRsR7jO8dq3YG1QTqqKm5H2iPr30WqcuS3hlj0FB7E8igi
4CxNmQJZxLfmwBfqvzSQY4oRMqAJuvtga8CCqNavOBCPqbrfaXtecQBrJ7YBATgx
yIfE94HhWFqOkX8fJlmiRbi+RYQ0/R0jkm37fab084lCLWP+QUdSOI0wY15dTIZC
b2u5IX67Z3MIGeJSFp9yCD7mEx3/fIIRL9iWftInxA3FtMu9l3y6iYmLtIkm7x7a
SU5xXRmHssw7jnKoQxEMmSI16cWjHGb06qUQ7Ykju3J+gSUw0WuaEbX0Hm5PtZgi
NzMlqdiYd4tlsZJocOLx6U5KsZacMhfFnr/7AVPEuVD3v9dyWwq/1nl7fpyhRW4V
15WzoQPG7Pw9mQMuifzy4OTvXN6586UGBfOe78pesKpioQi7bXBxTIVqgVEzGjQl
I6yRViwobr6ehqO6Jj0YQB27OVp/Rf14Ie99BRnx2Y3TFXfK8ZHi/sy77RvSZ0Jl
HK96wUOFieJi+Re+IunSO5UnCuqddQmTzCSDL5AoqBwgiEWx/d33TxXLP3gJfmUQ
kWhInVnrjV93FVayohpGgteWd6DCSiqBv2u3FpjgA13u+Nrt0mhSEzkeB5hNYZC7
B8CBabW+9yLNBpqqn2gqaqThbKCsjfVxDTtUnsDPQDvurHxh4n/nBvNZKbApprjU
eGdSxAiBDPxcJ2cqEYHJjMefnIKoPs7nqXO2ndQ3oA6NMxMa1cufySkP8HyiGiKg
/rPvDTQoF3sQgcYhZMb00BCkvRybp4Sk4X20i86J3mJnUNLvXNxjrUobLF8NN0E8
k+QxFPiS+PnP38pli2UhQVSDiwjLOJnmfx9KyKaP7PmSHIdcPnuIygx+aBHwH46F
ok9A+6TZ9X+gMNGxCKnAx3p175uwg5mmN8asv44MhZ8DStndQL8bDxa+xduwTFz1
47jG4VDB2tNYyG6/3s0ty46ChTxbDS5OKEKwH/vgFl9+fgJp8ehTRIrBAOnVpWnZ
kn+v7309E9yLldiCH5ETqeC6YhtfMrmpmE+I4KDDaaAH24TBsFxXFOH/TUy4CRBT
+fKrUp4OnJO3odWdSvXzfvaPGB/9HmWCCzz+UxlG10cxPALjTo2vb7UcwFgXNGes
mxLyiWIoYdqBLAplNqGzLuCaX681+WtVrVElE8D42BZ/60RodzQNwJhQQmw70goJ
Bg5XMS8yC1JAN23D2inBmvFtaPBbSZw83MzmSe7F8Mk13wXVgxs2Vru5emP5Sma7
zkrIr46IW5kgx3pUnTGmoIrwYw58hrYjqg88+bfvwIJgrKeGPuxlPiQSEoDR1cAz
uZ8NIukaNEs5XhYMJrTt71mWRXOX/FK6TU/4S7IoUbzbT/APBMUJ5iVH9sOXtBAB
CEmNpmAqm8UuCAOZrQVFLFCg6ptyPIYEFo/4INC2mdhFuI90zzz03WegJ9pG6vk2
9aruG5Vt7GHROLK6n5QlEhA4iuWTPf/rIbDjUZRCPvphTXpMCAfSfLGnm9YVTrvK
X3z1VFzxhKuTeRJtU0KEN2xrpv5kjNt4McyqbyWTR8FrUKv0uIWXNez7bVTK/X3R
W9htWJo5KoREqagFwCCpVjkThLdM+2vjNU7lA3eviGPc/aOHtxOvlBTyREuItVhD
CYwoQi9ewKVHAnZ/pEVfXOX5AG+nXk3a8Ik0gYlcy0SRL1DXPJdAVBdJ051zoDf6
RBcMnEwJnNx6mOJQvU8uw627hMdZJS7hpwKg49bJ+WRlc7H+RSzPWAkYlo+Om/Yj
4o76urFGE5V3+Py8qVqszzU+QnSjxSPUJ46+4p2GhmpX3GJRq/62Nic8Cnb1aYWB
7BSVeawaxYOUr6D6NI5CBRDSal5SKYt6SNarKZcyFmtLxafRwPzvTrrvsAd1sUyA
CsNPpwgRoFHsYstWWpkf6w8mT2/EcW4o2yV5tqmyiOA7gTWGoyuQy8PmHFyR2C7U
ncIFR5KPAKPukrzpJhZ/p0q3EmB99i8zTkMwAbII9iBtgJXiQo8GwXQav62AtFpu
dC5GJdsRy/16+E/FvNctE5/mlpoJUaakLaT9sGt2iIiK7Wt4FUTvkhrOKj7IA4Jk
caiEoAsTnE7GQLfgF7s6n6s6qhN9+qR4KYTo3Rxnba1o/VueYpsEoWp7esArZFbQ
ERRyuoO1Obgz7hmoZ9tX4flQ1u+t3a7NTRi73YTY9vC05zWumJxlX5s3SM9d9NV7
Kbw/8talrWI2osdOTh3m+d1+8qSyu0Cc3MNw81UinGUHALP77ImHOIooVkTYrS5M
wyf1thX1n9BFaTMSrOV7BUZhUxqsoXqjHao2wDC+o+VPJBwFrAW6+EZ5JLH5ZHwk
aSmEVhZ6Vc3yixEbpr0ZN8CTMvcJBOmN0RhjSpVlpAJXVXB9f1Ye7gcMUy3+zoSs
VhkvvTzD0UYvWsde4P7IBBdwwP6xqQ9FeezwKPWKVjCzV6N5TuU3A3o8kyIfdcAA
DB+rxN0bl63tbw84dXDAPHYKEMbD/oNVnDg7n+QiLoX1s2EonDF5uoEin6+kBtw2
LtEV9FN4nlXO+zF+6lJyqLX6aQ3bhqPGFxGuGZ/tS7eCbcwSV1Oid9KqFihJXqLb
KpzSyf/xCyhYLlKst2Vhps0GDcbBs/tMWaWPcYjXE7WLIjLzv9av2R39DCxPN2q/
8QuAkfMcmOGy3YQxK9an90fSTT/1k/NAhoupiyzVVcHvL1iUN/Z9Mgllf0/F7oAJ
gRQxDivYHwEmmMDPeogzokPgJC+1Vu4zuSkOMbDG2cZaP8D5JfUU5nGgi/EFoVWZ
2ovZc8Vg3uMkKkpKFej9n8kUjMEeqLCrq4R6V6Oii6qrFeufypZ/Qtp1j5lSi5fY
b7psfHdbRlJVIKUnPMFKc3I1Gj/cURmSUpjC3iQi4QmYaZcKR8xVAetzx3AZD8Qw
35ehYirmkfqQ3QamHZrWc8QMl6iknkgA5l/9Q3b52PuJffJ75tG2QDtuygR8nspt
oKQPb3lK8hvnYvf74FbCirxcS7hEKx4JbdONwbQH4UMC6kWf94ldU6oBW1Nu6tJQ
GswCIdwyv7MA87MsQAtfzwhiC3XSOt3VXOiXSx7qEouseAKB8oWDdQQAvy7gUFTd
LuZX7m1NWdq8iBUeSegs3+Wdc0oallgtBhl553Er8l/5ivnYDJ9LqxhQ/137KWz5
EmGhtPhAP6BfzU2gyUSZXum1woelrj2YgqkeUTJP7s7epaEfaYi35pt7kI3fs6If
NfgpZdY9/3bi586zjTpDAwOfgcBA40zq7TliB6dEigmDDDB9fZ75rGaeh1AV/xVl
vcVRgO1W6v1trHTTn2kHete8xe2BP7VBdajDLRQmI5WC0cv3KKwh4wy9zGh+q2bf
4h+8YN0H1ZbftHW5S04Jkcbe16St4SzUY3wPLSsnaGof5K+2ulP9+W6HjT8LLJrH
VExMGWR7eW0RneyeWOwSq5+ZMvbW5Dknp+XtjLl+8aDJUO7fOfgtDMK/UMgIJMYh
AJ2kiaZ1x1xkuA+7fSSeITKHI3f1RB9Mx3QNJ/qLODU6QsztS4Lq52/HmMpMVS6j
8W01B8h0IJuL3o+QBjCStab9jCfcPDNa1NVfF+U8kWMZ/syJ4Q9f319v8/zc/KTg
ND16GOUyJCT5fNgMwHF7p9tXYTtfRXgv1oZxzXgBPrW4Isp6vV3p54nIx4tzWCQL
jHTS5NuECs1VNULFZ4aNL+v32O+4oguLureDGkTuT09TxxWJXyblfdcaZPHP83xf
9JJZz7yuDXA5CMNiHn+OGoqR9htEIDkxpKfC1jtmekxfpK8bdN/JNyREj8jj1H45
0p/XDjvu1Dza2cHVrctOQXrOgXJdpSYu2BKNwUXZog7bvaDMYRP7xqLz+uTfZpHi
iNDG9GIRAK4D9Z9ZdsRYv7rHj9/1x0SrvT5NCIOIOPLsEatTqSFIO6/mkZKbCY5A
OVBVIysKRXY4OOHKTYvTrbofZYTbRAjGl6QG04jaTcvrv0f9fKdWFXH5dKlI/30N
45SQwXr8gsVhZ/5ncehSGDiLyHAMFKw88aIOhIVTpYSzahV59ecSJUwVeDT8gUNo
/CYNAl7zz206pa8n35EMSEuuRfG4UnU88gDq9qbA3JNAFs8wYKylW4MV3P6cqznS
cRObaj0K00HSzjO+Qht12rlqCY+5agd4Uaz/lSznU2WEU4+wDZQmy/CRFuxLf8PW
NGZhWNGAEDCNwedo0kXNhmZYdbb1yBF8QzklDUVam38HMtLovImiqmjhp+IGZsZJ
kuwCTPCfTYFeRaK1cDxVnTn6GlVzbFFkIwPg5OkeP4G/1RTkP8AVxxXKxFeH/x10
F+R60PC5btODlEjO9i8OY/7XIhbPjoFya5MBedVZI3BwIvS86D9f0rCT5lRJ3fAj
1X2EaZAPJkV9Av3Ap0MoXniAj0YzLr23tT3Q4guX0+8fUg0O+xvEdi6OIQC42bQW
PvhdtlaLfvhVFs6HTex1Lbu6NGlz4Wp7Qqw7gGMx74irrKlyY+Qh8tKMp99c3pZK
h+yf8DKvP4DK4oIEMrbQOnJt/a7FFp6xs40h0UgT+KCOWZxpSzm+VdLHa5o+7nNE
56WJRSJ9IYtIlYXFdof3J9Vz34aVg0E7UO1iDsK4NDexG3nnU5vTBsoGddxd5uy3
wEJsiWPylgFSaV7mebPc0PvCOEi1vAbhXFjFFzW0FKdkNPTibEDMzgOscBugwO2S
5JyVae97C0Pnyc8BbbpiH3XRoczDEGmZEGBKG2Ge6+fXDFE5uM4AlnwbpwR/I6nU
IEuNOK2MDVO3VfXJqLsiiufs8Z0VJMf/ETkJ3OWNCS8SpnKiYxNuYDjWLkH/HKQO
Q0dPO63wXq66lGbR7N7WkgqL8DKZPa/GTG7/K3OLej/dV6taTmhJrhYATF4sQ1Gm
/uwtqhmaIXlMhV0+2ttfREzlY6pEYMRfG4dCuix2rPEUdBi3c5fKn4OnZPWSuady
lRqfcwQPXtK3wESWCiuPwquNjzimUXmhwxGUxvANF7DUc1myeopqL7v4LOmycJUP
tnr/6l1zOeWalAea/QZbY5s/pzZ3NCqkTYAPBOYHz9kzCH5FBOYRrXcLSTAbEPz/
v8GTKAM/JczSHn71VvlYU4W+h1vac8WVafGirAn2/N7U7eBaosaQsG+qn1zpdT+m
R3NNTvC9T7mQBQF92hPsYtNOSQfaZH2/YJCZbp7MYLEDpkJUwqKW/Cwrn7Yepoil
q7stxIiMmi+l5UsqjO3Ld7FQ7WvPmhUzYv7fprZZgj0OuaxGYEP6UMVgftXflpNo
bI2I7bM/G/Ed45K1A0YNwD4068meRe9taaI7YcKRcuvSZt/4rdunTnJjjAxwyZYD
alkDZWXBraAfhPmqUJlx6gdZxQFzw/waWFfnI2PcQVJfAVLzVJHMpY3XiGbmCLJ4
vGUVh8ew6kq6E0qYvklcHNidoIly8JavE8+ZWX7EGDDDLvfcLD+6R5+ZHuEAFzgj
rvVihIeG4XoYMajzJpOPVHthpk/03kJ0iSVwcrfa0tLXZLKomICrOPPvFFfTVwfJ
V3Kq4sbRfcc25nnyNTEsz5y/AEH7wHTimtdAE2A1rOviZhCBtbVE2hQRltjtPeRG
6TQEyqC+oaDYHcCEuNx3gYY3uY/85VRgwccuZv3eH8ItFtir6+ZcS6GCSv/0McyR
LYzOJ6qg4jg9if0YWcmugXX1IVDMOj26/hYGHa0C/sYDTIDBMuoCNmlpI7ObbIbt
RbIW4rYo3ItJkh+TkkKTVfh2goWvOFSsoCYVUJe0WD+w+lVhqCWpJULkpkm9R0gE
LPkC9LKbLufXyyad3GpWufWV8Tirzp2PNaV3JuoysRfeXMqbzh1nCp9nBWdlRrmE
P7AK6/zufveprMR8hLspFdBBRsaKuAleJ61TcN/TTP42ayacAlIh7+Brx6cKa5XJ
FtfAouWSz4bJEqe/qbTZPBDclzOmqCtcjqvDHdTn2wN/LbjJNhS+URARf2RT9U9a
Mdjv9nQ9EncTlQ28Hn3QKTtJuTQqkEkKzpk5NjRokWhnxDSSYf9DhausRdBO51zc
G3VNyjx0ODk0HfCx5KYZP+I3DZLCcjKzXg3UPcZNan6b20thdNLIIeQe3Q0tPIrN
IiQQWd8uMRsKx7r4ZM3n4R47SPzK+1ESHI4DQuwOkvqKlwconN5z8rP+Lm21/o8l
kjoo9E1aljaP+CNUs2Z8eGuntlbWi+8Cpk/Kawav33QQMnnVljV7Mx4lHEcYmnbk
mCTX7sbACh4mIoFEypB1O+DgvX7bsLglpgRBYvQpoF3HvF3So3Uetz9WUESPuEsO
55hmAfhsPiegPFMWQrNoW3OSRs88wZgHXU+jVKb2PtuiA5RCqs+WFpbw6T7P2jJo
2/otvFem9H7hA1R9QXx6w6eTzLb+DeMG4VLPy29C5QhwEKNOZoOzeu1qRs9l53P7
TD2QGnXpRHAAUA8ryer5lFhpWW2zlutEzG+4IirG+bfL9VXGAWdPqj6g/jptCQqh
CkfNNY0iHvfxlnpDgpmcGbE5cFdtQtNXCfGkSZvxjBNU1VOVR40LbIVvrT34MAHl
ur9t7+JeGSb1IlWj2nvuRyTt57QX52bQU5YB5MW9JWhTS8HySiqU10Yfam8Vl86N
4zTVymby4j9hcwx0hzKla/PRStIm4vF0Ynp4F0W10p7/4kh7IrS9qBK1+cBS7kO3
XEtKSHHxecRDDRe+nWAzYl7Vql0qqCHG2jwgRfl7uCDBhVpkXCG8seWs8y7oARBJ
Y9yF4HLsYV2tnbxwqiq6hl9tziSqbTGk/U0QcjFTFkoNBIHVTwBlwHm8HfFy0zxV
W/Kp06tpGVdc6jBKUBVBrPSxsNsRT75XOsJPJSnBzt4QBLkg6OJ88rcCkqSVjv42
TDSek2dvGxNo2nPeFjZZjnSgETdkqm7aWwK64o6odtdbwAmqGMA3pEngAyg5HwAE
sPHT9I5Tw91ZrhmHEGPDOn+PpO0vknB/3UKSA9rFm3S9WqpaiPYBTvzAtWqzj7lT
AviWZDB0d+3pJnb0SkM0xUcp+jHzQHv3Crxb7BsmucEdQfrDi0rO2kZJDgAOrL/J
YwQMYIcD5nm2Hg929NU6d8QOlWIlMJAFGTX8O+yzRefz8AVTP5ez/s4EnToiY3E7
GdZQ9hDEnoc7CjN3diPIzwmyWcoZ+Upq3wDEXQYidcLDhVtZbwHUX8HG7/s7CLUn
S+R+mzLyiiSL64T1duL/L43bTOVjGqMBAkjLbrGxz2iOQ2CeNWSZ7+UMhqNJgRWr
nt7eCux1wcdsqYFP5Jl7GpTKKzObsUnbyTv6AKf1wEtGr+aDzFkR9E0fTHCpxN3n
C8EhTwKYyUUvc8sEcGC3KZa/huKZ5qLqfThaODF8YXukqOZdE3Xza0tkimxMVgfM
mi4b2LMJWV28evMWSSKiXvWPSTUJ7ZGMaByDSVMQnhlbfxCpMftVFbW0qs8LwC8a
4fVGQVLDqOjeAzWa1V6N+KcWjg9hs2TFNoEQ9yFuM05jq9Jx+WRCmOv6Z3EM1ZIX
o3uyKIL4Q18wipPvtwdHpMKBWrJdj9rhVKFklWhHwwHHLXvQfwCZPDk+Wbiepr1v
cV/5fum+VWIPrCE7j767CGMfhDUPdejQIHijbhRF5Gmj8YK28Jw5zi3pTa0xzFYB
BFFmQLb8Jxi4fbdXGW4Nroc/m2ey6IoGfhi0iQJjgkyJ0/43lxUyTp28X82JV4U+
tMiBnTJbqIn2n0v/qvZ1woQFoS4UsfGLHbB3/hUm20SRk8U+PZk4QWGSCCJpYIGJ
jowCRSlEJXEm4rVOjg3GkFjjZ10gVZKteqW1tK2enr7kY7GTYsHxddNIUr61yMuu
71dsjl7VY2mpCbUXw4LJBMEUCR80kxVGYQrhGkS3sGzVMqUar3lx6FiPbEdKWfqx
RxhSYHDqMZPvdrmXELc6oapJtqXNzezEs0F9f21EAw0c5riml6sAlDaZOKzyPbHH
w5mAQlaSW24h6rWrGOOsq00yMXykgujLDt4gsQ/i14u1Mz202JYtuinNqfayD0g3
E2hbWIwWZ7eRR4IYnrjbdbWLhhbmA7TwQywY6LN9Eb6W5RTK6CVmm7uNIddCkrPo
MWf1jM9hZLYb6OJ99r0HjF5vuQbQ3lUTjX93E1Yhih7nxdQs9TjNeZ3qWDCeXXoB
GlDVVLLNAJQiSXuzdQc/tkxDkWZEOs8w6ssTYHr7h9MLtE5wURZfF8dxlS2iO4hW
M4uYmurw+3cO/vxCCmEJS5Q3CH3KehtBps9vM0vmUHpL9PpxYRiMRYDPU5yyrOxn
7pICCfERsc+vyIuHKx7hguNPrkt9WkX86KkTy7rbGuiLRBUDF43mv5NQ93pruazA
1CFvYOA+TGnJmFDsNxSvt0qXk8xWvKlayJqIHbFPDuawuMa5oxyyEB0rPa1vc7JZ
0QtKXJoVlqXcZ6h0m/NZ5Cx3SZOUey+CIvAJ/gSJ6BXRedQzrlJ84RFpHi7iE6rV
689oNj6ESDEniHcaU3AkBbSLPGVjJum58pQ7kN5GrTGK0FPXs7cvjE+kiRlNxS9T
QNsxfN+3BNF8pNsXgsmIjpEhLPhMbqLbUKxQwMd+DPwBSHVibi8PalYI7Q59L3sR
snFudp/aqb/+NfkuX74zvi4U3Rc+Bok4+7Zi8ug+dHek35/2tOeCjoDbC/bgLQ/L
XTIhKPZsT5aFG9CJOoLKkg8qdWfYaFj/+Ai/7zCqlcBwZWiBd5I9gOr1U5bqaqVW
+UmToHScOgi0wxli5UsGv0ifarPKwA6q/fIgQ2a/2YT12Je+wav8bk1IHbCtGz/t
/qmA+GCY/yvYRSCrT5PUQmPWdt6/dJjdfvJAbvS0dNa/TP+udqVN3fHxNvFmzWHn
XTdEKx5Elr+ssS6FxKf+cbeboX7ZeQLxhm5VMpTusSfAjovxg3Y6+qanycORIxlc
EthSqFARlsTLJFMW3NjBHUEc9rdCFskOhJQ2a0OnumMD/+du/C6kBAg1pZD1GstW
QAjz9AS6bce+OS8iaLp+aQvUAvocPKlGBnpDm1UCxyMBjvORotaK7TsmoEBKKJ2a
L8pPUXreYAlgRErWWGT5Yk3lcqKINXiH4lGgeJ61GCkgbea3/BNwKochphMEMwsZ
r60cyHzBijlGdjsSr3B+UWUvxR2nin1xN7uTNSMMIKJ3QOa6mMlrNSg3T05D14be
6Mh3TBq5J6Y8s08KBdp0d7SYeUJMd4g7y+HbHSbrI2l4ioLQ2qW+6Yzv3e9v178Q
Plw+jbJkCKSRuMwdL927PwvAOb7fVH5CqG91OiuGanLaFOv0/Jws1QKoibQ4SKZ1
Y68aj45gf+XHu5UEgnTn040UM9iaS80N4ZB9m4gNbs6o8UJtFB3Pt8dl4tYLcLce
DZ07Ad/IgXUia4+PiqN/urD9EsXTCRmQtPNsL9jx2uFUL6c3kMui/BVP8ZKB8WG3
IoRHK/Jqc7toSFSWisfDyrzkg7HO3F9OFh+kjKcfcJHU9u9OCvs6Fj6E7+LSyg6U
2hoCObPX2fl9+R3nNzq09DG869P1XBPi12mv1RWe3et1+Xe7irkyrAwPvj+iOjzf
GlyKXrnLbwltlphFk0vjmcEJFr1iaEXtGG433ivVDtde6Pel+uQBAnG9+D9gp86q
znfMBQ0BQYVoKMCXxRYq6kvjcZwGxc4KC4XAXqgXbfYoGVwVscNOKGhpKNSzVHgU
9w/4wOnkvn0wvoBFpTMdEMQrMInryX1r9RmQ0IPUx0V6NiiYYT5QW0hmTO2Gk7L1
1k6WNmHbGj1QcF3HYWImXFg0c1PazdruBL8rKLZ0+6xp77QDT+OI4kjLXQlxLaem
wKya1tqymDc/4VCNZebLEKxh8seBKfz7/evEfJaf+R5CAqiB4xbUrjWg3wOicC0C
Cg6LZWEBsJn/uCqaxc6qB9UVVYsqKru/uBH5cbtjgc14/v8ShIakn5M/UwlaY4O5
pqKrDrY++oztUG+pQbqY5FPUFvFOjr980yvmcsAhlU1ROd35Mg5thcj/1BG8JI7Y
+9YS9aNrtDGhuzu/6rlgx/GrjMFEoPuOEcTpl+qad4JGDRVL1uQKrR1en0gS8kFD
kxdYubQTp3RMwKTQhTaXne/Kmq1YcvS66Ht8yoUfy/sJqfuLXB1BGmlp0c9wa/20
Qebh0yxZfnc0QagLWPDTSxE8J88HMgsQpijMf82YV2N9hCUisLmLtCjbMPn3tDOl
A5etPAEol4FkQ0oAdjoC3WDWGrw5K8OmPUJnCtQu2w+EG6eOist0cWkei/fGAIoG
XcptaHhsNH0bh6l0gzKi0kzLjuBYc8KZIsG1sBCYpGFvFN1UUjcrBvwTNRjSMu6l
G+n2D6WC88lWXeSeNT3Hk292fxtnZF+QTbu/wf9bfOZbd4hR+MzMovkcN+j1hYB+
PxBVcI+6RS1Fx5St5pS/Jub72+eGo78iCcBmoOE32CuSXBHOIIfu7f+YM8J+HD6L
itR7xWOo0IHCEUDZWZN08l0xqaQonFgwaIopfwR/sLnJfCry2OxyoU1Yt7s49hBW
zzpyEh8IbrxpJyrl9J8/3i3KX9CBtXKoN3H0fO4OlDMoIVag3o9mjK1M+Gk8JTbI
ccUtLdVOyOd2rDsGCtwHTkiq9fXDbfEXwCVeYr1Y5Jp+PL0iLMF7RpAYnt/twzFs
NZfA3kxBExB1JmsyT/VxxDPhl9hzbUxiHwG2G2f3ir5kNQvH2TIvBAcEp02bUAm8
H+EqgjYszHZcfC9qhdFoqEKTdAGhafefXOj3XER6j7J+1dPBJGW59Bq+qrEcfOvW
u1kead9arKiPh5rOl/jN2ujUytz1WvR1rNXyP5soaiDeO/JaMzKYKmPZeo+m+rdB
WZiQ4JtT21kzGb4vHbFm483B1gVmsfSaW/o9/lbhpnNuMMZmEPvqZnvnKAshlu5h
L/KhH9dWTofkmrEOCQRmYd7XqEn8dohjdFwmNpLRzpv1itZgZFG0m5eFRCBV0fy1
77/cnSG7zdhzkX6/ptNoEUQSLeB6vqFz9IqUwHykWKF23v0/hjFXhGrEbfEvbv/f
8YGX+WCtDIYmz+qNnwIs4TPaRQTLt0dXEyiF2Brk+FL1WcejPmPt3YFBjFRyRm68
wnxh9Q7Byw3bfG3U8cXHQpMyooFU1R41l2AjIP9Wb/K4qx+u9VoScZ+0mb/VvPiW
pyYMIveG8ADswv70DJgj9471aek5pQYv4uiq+2+4H7XHJDJFM2ls143ioSi6hf3p
3mRPa+HAKRyoiej293gK5g/pFwSuWXIRbndJMYyuTaYKxCgCWsEkbuD68KfaRUK6
v8/Av1XLUzlO+rAZN0Sl9fwps6T00u1ntjc5jpKNvW4P0F5nrDpz/9vlgcJN7Wkv
4vb7Fb44kRfwLtLSie3LHBpzLjX6Dzfzwl3kbb2kkdnt9lO7lvudWDtOKVPmrNpT
/yW9cdkCfChIyS9vKovRx6pxdI/8WJIS5SK8SFWEP4CHWZTrUuZP9KOWslzoub3x
q1gL4LMsjTzPjJX0hExN1j/q4SbGrUpaoUK3xBWB+Q2GnYic/exgA1g1L0tlpGzS
4omf9zSmRLhofne3oi9PevgLlUxviTeiG/4SeuJadzVrRTOgdaYW6iINDq1JRQMZ
an3szPoPxmqCcv6y24aaxM6AnoqSFgEKd3EmAv4D+kT86n5OE7UjZQi4fMqjAdqj
JZ3MLonzyfotuNxNf4ns2J+ZGJpbIo77hSJVVWxAgw6nOYxhSyfvTy86iLPVjLqr
1/oeg1JKStIRIA5LKMFPeiws+0DFxF/nF5VmQhNTxXmHa+NQwOXi3Oi01v8s9pKR
+yWeGvetPCsZMObGmRccPwJ44AUeY0VZX+EINYRAMjKPctJzlitIZnnITjrgKrFD
eBBfln6Uv21Y/+s/XAr10WWdlpg7DRm4+ei5+iBkzq7fZIuGjyMbDMipJfdF2FsQ
0NYMSCmod2/nsPPw5TqnImjeOTYR+j1+wPpfFajnRx32w51W8Sc8c3FDbtrykFaN
p6NTC5sUvdkkPHBMO3orc0TWpkqdCEd7W7itqpKHjfRkLfyLPURI7Af0Mn7VrwrW
jQe9DWxSmqZ8PDaqAgQHJb2FdqFQd4MHFpLRrHQkzPAO0RIperCz7PxYdYsg4nWR
eM0fCHpwYxM3g+jYW05zTAEcxQXyByh8MdUY0cwVTPE3GrsSmrIZFGfal6IMUgaG
hfpujGkQcdUDg4UmSuYN2Kvw2vxWPtADNBsHivKcrsGJXuKYd/fShRDCwFJ2Jf5P
h87GQrgTQaCfPLg4YLDqS7C5MzrlmC5gbLPCz3M6NBgAFTnbVkiapnMf2zttchbp
OCfo3Z4sFPOdd5dxiJgvPYrANpqq71httvOTx0LWvd4SLzOHiZQEZDA9FrKVZMFD
ABxYDi24yPGdyfbSBpwrj+biRyk1smY0E8Vq4dIrz4I+vEtowBjhSCnhl2UDMmYI
xodQ8cgSR525O3Okr40Xl9Tm0xjg9T8wyTXGkrbM3S0=
`pragma protect end_protected        

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
VnX5yMzl5xtINQYXkCMJKJT6+lBQGRROC/QuhFeGrpuVbWrJTzv55OzK8CL1aYR6
f9MAnYGVrxWa4e2TwlpaUwvUIiReLGROEr1qQc3LCWUkAY0wrnhNJs/2tGWHa0lk
r7jo5drKlErfkc45/RxzFbxRonfNA05JSPtwNvi17ro=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 79873     )
77vMr05o2l2fnbAJK4wh4rWNPWWSCAseFObUdJIF1zpIktgW6TDeyzKOxjAuVRyS
VYLJWVEFa0QC9kPrc6NLwt5C4EAreFT9cbkAu98LfO4Cb6IShx6F14XF8Ms/Ry6M
Z8h1I6BErLUOKHA+QB+HuIpCsz08iYf1tNnCweMmmpmTIMSKdwpV/7EwffZvnB8J
UhxHWKvwGJmU9nLyYV032g==
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
GrdLhJYfHP9mErPT1BmA9GKxJBJo/43/vgfTu4jEiu7gw4SXERbZyYc/xOUonqzd
jWFFfnP9TL/qRC1pgFmy3/wFmnmfk4RM5gSB9r5RVslDO0+gO4sFvF1TSFMtgUJU
sRSFOuqEeTfOp3+rMw3KBWHmxPigPmySOILo1VWs97w=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 83289     )
4nXBHnd1hELXb0qMba83f0cKz5R9GmiUEK+3jcFk64b3HnAbLm0d3pAPrr2xecmv
/RYmC/F3qjE1b7bbvzvRmV6PsZcBAkmnEVgl/yYB18h9n8zQWmFqlU/nMcAPhhwY
9UmUVH8yDd1WZpiZVq1HgQfrDaN1XQnAPTDjtjPzcKJp65Xmlj3uSn9VrY7hNwTn
Xuo571jXe1FpgIOGkGSumQXK6UxFRonm8zNuPZPr8LEwJ3hx9foExCoznf1WREP6
O5lttqJXNmiRQx475GA3//IvLClLoC+ORnrL/qrW//tD0kyXmzdjbn9NsG2rJgbg
13dFEY7BoWnfcwY3ZyTXd2QToJgVUDdI2DmsgcDERFw6yDnnCeWSL2igMee4FYz4
J2EgDse0P0L+VfNh40OFHyhUWnlkTwXKwt7ysvVgeixUf+mQ21KCOizEFW2ohrKu
G8xqhhieD7ZZRtPzCEv/e6MzwTeufe3mz1Iq+a5u32Mk7bYuSEcUbqw+fHelGTfM
enTxaL2XDmU9Q2NCkT60eaFneX8UtdAzD1LUclMpCY1pnwCwJbdGbYLIDVkFW7b3
Clby42jXDPjGdlWTpJoYK9ApPbMRhrH3CXJH3TQJqQVJqXLSDrNsMW5pkpTO83QP
WznfNeMI0N+XOi15bVT1Xb8/hYSYWCqFIc8UJ+UiUml28Uo6xgCVQO8ZDDQE9nMk
Ryj6P2r9VFMJi7TMaX1zNREhWLbf2jMnr6dPTQumO3zi7C6+2zR03E4fyJe5SJVS
x5jVpTnjYpuRKTJij2GrO0MfUGnzp5WCukSzkRO3R9QuEjKpiEEcNbjWGP2zArNN
XX8WZcELx2HnQdDSapPutVtPsfcsO84Yn25aSR4Nq1Ij3JgLTUx4zFRKcVjRKBnJ
hU9bNVtivSAzUAyBRO/23DtP95sWJ8rSMUYKTj7L1MNOERD6ylQwkPn4Fg0wEN6A
2dpWoIWx/musdwSv+4VJspX6rJ4iV6sHcRWrhNpcmohU5KT8xvjD49FMNiXdcS2v
0PP6p64v1xF772MtMJ8wX/Wlr6xpon3UG/8k3QFWFYo/x9XUmkBT+WS3JPij1i6U
SRd9SMkRFZJLBHgjR9cCWMRbNxw6A0780NlkZSjZuN2t046gawoT1BVZJ8+1m2AE
g828tgjh+TKpoHBUANtF33Zliz39AI1ChynZsRv6c50XfjD9K7YZp1m1lzSlYJa6
Rw+/XgEysd4QqX9BtJ4f2ucwCzWYaq5E6g7XkobHAYEiRb5LsGZ9DQXPv0wp6FA9
Ff2daC6ZDne+l5gvwY+bSJtvO6G+rKppFtV4F0g1GyIolOSiHlp6G5iIr5wODSX9
QAmLcVERPjz/KtKG6r7cGXM++d5pLNGc/TxeskTa453HjPYa5x3+hDaO7o15tbhY
aw51cKRWnbkWQl8ntQW8i87mJE9XoRsOgUXl9T81uoYH0ltj7XzgUDPL4gq+K2wi
vVl0XxN4e14rQVZfughqER+TtHL2w+lu5DeF19Vh1Cmlr/kl1BoynpeVDZI29Rmf
HtR3nHmN9cLiUDv1asAV2tqx7UZZJCOt9KUYAJ3oMgV5M9YhGYcaDydPLUMlIScX
FykS2R0JSBX+CMAT07lDpK3VvOkxz2N1q2CkX90gOd1ngpdDzJS4jK6aQOhLsRAA
+N2Dytkbr/ypvzCqIlE3goBRusfRLjmHSIXeEv7MgRCl07a9rXLe8uYuvH+XWsCc
CXjYAI4ZZWqG/F9EZeMjSm9YKqE936ga7Vcgc6dVaG1m9I5fLWwLUc6Mf837XfLL
NsgWY2DZ09hocHcYvLqJsaRaVrl/tjcTswnkI2VCnq7JX1MszvQ3wcPjhefF+doc
vONDIQhDoDfVWLp1BBLUIt5bTcf/1NnJXiM2S+WBP2Rt0fwe7/vYc1+6cDN35B/z
raohJVH4WfeWkqjmJ7kSvt5ETcnyHjnal9SUyQT7mU1gPqOxydWFYzYXqw63X32T
Hxy1cOxCvYyImJcWoi8E9TND+9PyF7Qpwvn0x1k4XQcNJWLzwOys8T14nMr27YNU
z/87jgtD24yexEgfqJYXUsrAipT/kSvdarEtxEu75453HGvGAXXNb+jY5d9aYgDT
WIWXd4yymRqWCmYPYI0UC+pvwFrcmnxaA7kZq35W9VvtaBgn81WEcvIInlPerJnQ
LJbDGU21qH5iN1TDjWlRZFTLZDwlu4FtN6pc3TggtnDldkQL8Tj5FTDZ4mUoAEMl
4O2WYWbDegkMXCBUkMAcdONP/egyhH0xyuEC6s0Mb/p0IrfkiXlNAeDZrCodoTtr
bNDWmumU3FOCB0fI0aNwlXn2h4eR6NeDpsJ+PxaKZ3zMwS6zH0Na6Gbv/wF37tde
0yRcF5PcQ9PMSZgRdEXHk2MOTMYT9lI/bvxlER9r287GsDazm6viJ6NMvZNNljdA
BppYiXygpYBfb9Sa2kKe95iJkKU4ZeroxCy1nTwredxUK1NphLqGUrHTbvDkf2HV
8j/HYXhy3++EBNhH4KR8flwia3aPqWsbK66S4WXSy4uO2EK1gMJD79aqd9MaaSDS
+F/CT8g56jmwg6EW2HWFzVhqciYyGCz9EUsIOzcbcP0qcGllkSMRx+/ERKCVMGjC
KapgwhXVDD+cWJ3kEbLfUeFDavj+9BPAyAbBW/SH3qwkLLAyd2EZ6/ouJkraVfFi
HsNZdV/YR4auk+s/9yNztDf+UQv2fbKMxDSc0MW6ziSy1iYMGTAXPuwhhabJS2A8
u+p4+I34IfUdwBSG4tLrs1u6VZiV+QrVDJ8xsiwkMXD/My3mVMV5JB2ydo6dzNpt
9L9MiWcWmtuP6bn5CLEaulu687pbSjaxvoOeu7jEWqbHyhd+LmkJ4pPeV+qhEWld
JYNcENYZ1gKALisIpOEsSWTKBezluxUtpT6D9wj7VNwXJb8fwv71b1K3QbdzKCej
VyonWivpt5l4PhVltsbLI7s6pqCS+7Uh0DHMDOwZmqhjTtvhG5VmTjuum7YdlEhb
gQkJTjkWrG8yhtS6LPnPkCGckqi4TOa2UhzY+0Bw06Mxvr62G7mWgtql7FP2EYe2
7CXq0z+ep44dgU979mtQWv+9heGN0qqk79zgIZt4twaLuqGzzpdWaAem9Lqe/3sa
vqWunQkt5brZSzAmZJfkWbCkY+0/Z1O79Y8VBtGdSSD+zFOR5T2b0KnXiAKtPZkm
fQXYsuwnVVvdMf4nMlaghLs1GM7NBoii2OGHslvtQ6NpKZNSpwksnwfgUKaaWbtM
5YeLk/IGY0DzLz68fZ1c4VM4MgtPHMCYAhLLCPf/ysVfOCAazvHc4zNjkKOeg2P/
hNdAFKFTzina3eZxIkjd5tX/xCjyTqjSfj/Y+Zx79ooo0YLkThODfoRtY6q541Uv
FEr5PRMu1R5gsuOeg7v3A1d6Y1dasNpEvrDMNE7qu9jpV10zpsGydhhjo99XfXmL
tY4enz7tC0wKXhZBpM0dhD7H2WGA5bbQOUf9LGzGpy0lLEzIMeNlbf3Hc0Vd1zRR
H0VmEjigHAU3wnr80wLWwEfJwYmna+2EbKFXegCwg3E70O06fI28U65RjrcPmf29
bKRuFAZfP5iW6dC/GEV4cqPghV1KidChvtZIvc5G846VkM2lY4F6iiSbZzsb7sYd
KML2AgAWaO6CD1UP3yKfVwyD/2OvRNuVPtbpoXNjHgftHfLAoGBP6nZHNePCmBMm
K1AloJsV8hRHLMnQKt6FubW4X8p9RiSNAtrmH0uKCZ9Ps+5eESp9fi1q7THHmwXe
MO5ypjY8R0ZZtTkN+EriBwYLmHkuPQksndlmKWy/gMDgej78xs+2k2nWLQBeeCV6
wh3c6Nm/DqzBMOC3jN1tJGhV6idfP5VlJnMo13MIA6P70x0dLonrMqGl18WH2NxA
3kbOs7KiV1fzZMjb7RuYtjBW9kA5c2vH7htYzcIw+dCqtiizHyel7olnkeC+iGn/
XeusElc9YpbQqU/seUuU7VF8fz3FbWX7n1sfmPP6w7KF2mkY2F2hcJnov90KmD07
5/yOiuxrhMZ7ZrTDEF0wsSqK6JJa4OnrlFGBVG81nT6v0GgH5jnG8ogJRZg4lCiU
KmGOphoyy5oeMNY1b0ZMvmPo3mkpx+bJ5G0RzocA8Ksj+5UOIfhV70VfozO5FVFz
lQxYiTfFPfxNw5pUpXR5OgPYhwXRrPceeNCuYhM1p45sWlenUUmgHsTnSDBIOnEX
vi3riHS3GPmbAWpJ3B5yAOAdKNzlbu3932ImywB96tzjZU40GwkERGuKy/K9ZqC/
mMhCz5VabQeDe0aiWeMf84tEmiXmLKKmQe/+HbT97NQAnJA+MnkZ4KiNmieWfbPX
YTFXMqvr+F59q5vTt+vQkdzDW6hl+xTXaE3L78MzI0BJByFNyg2eG5Nlmo2/5VzH
0LBZNrv5eFACOzPj4hBkcoXHSaMEi2eMytz4WeWb3LyqbShWHUVl2/ygF9WjL6mo
ljHnpoy9HUAqrCPtPtzJW2+l7Vk1cPAs1yr4Ksh8TaMzV6oGSWLkyY7qPKPf4Mpo
m+72+5RKpqwkElxe0g45Qw==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
FoIqEOqqjgs6C0AMa91VZUjoXeNxKHFqQnWo7seWlmXgeg1kdsgcKNa0JzGeJpoG
VQQLveAwkRy00jxJ25Zwxzx91s1QbXSuQv+DE0JqXEHFj1gGgu5zBZasZe0X5Eou
YNSvHg24uNu3YkO8jgnT3XZhfOZWNU0rTzMQ4p0UYVk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 83487     )
MMgHYe2l5TGIKf5/SbfC8pAncA3NmhTI6lxY+qu5ku3Of2B8Z/8dXug0Y31H5sTX
6+mlkvX9m+MAegnxthtB0ftp3Fr5TuRE2eCCbloLpTKf7UAQkXBDy0Er0URuMNbq
oLk8FyTHp4L0PnNyCQ9TgDzkE92ee2rV+GMvgYa4lvavx5znGZQts8Bd4UERkdVF
k0eQ9uPbKQYGvlfayN0nhqXCy1IKTTYqja6SGQWMN2DG+bPgLYUiJpekp+D8AMZU
BCJ/wasAHk4Th2aLYMxHfg==
`pragma protect end_protected        
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
DXnIbWXpE/cAKhhpR6IlAqa/cXFrDvbnGQVf+lEJmsa286Juylb147DnwHfMgdKl
F4Cf/HxSXLTcFAHgUVEZLLCQsO0upfXKavTB3hQ8qmxeRIdrIZJEsf8SMJvU7bni
NHNcMLJFrB5GgotLJacZ6Ktwtbw+fN02stKXFPF+p5I=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 172262    )
WhQN2VlgCdZQBUpOBNUxYAF1RdVCGW+g5zhHM0D843rCeOvSM/vS/9Y8n7HWEeE3
DeEa4yEYoVwz7dKTYt9JrUDg3Im2OwdRousFsHjl4vkQN4g8xVgAozYBDcykcS0s
i+wUr35vX4gP6Hjf5pZKmquZkmuwlmYqYyeii93zdwIC42ditg0wBkByaianbJun
RakA7rFMengyym24QRsqvIveYt7F6tvNvramNF+k7mx1Qxlqc3r/q8DVEPMPy17Y
YgqRwc7sC85kCZyH/tSpVCVXA5c4S1gw3btzD8+eg63cF5lcXhyAQ7Vb5igxe9Gy
Yv1bGXFpJ4MuZamsk8WLk5R9HcStZCDIhfCpQg581NyGSVrclFek1DPg/I/Bcy+R
2tAv7CqUwc5vTN8yYzZ23eyCw3niMRC0S7jwepCh76g0pIadf9DaTWlhEGbN/W3T
MijDG6ufFX+ZH1mkKvmapHodArlHHPol19U1R80B9V+yCM5RnbX7l5/sYToSELfV
QjLZKfAu3PsC7pNFzxKzUeChmGlG1uUJm6/Raq9SQPtLAY3ePTJBAlHs1kYnx7Ih
9iPvi8F+jt9MjhOwh6FFuz1aGZxx44HMHQpS1AfTipxwewCDACiyKHjrmOC2uppw
0EdEuNtIPD4HMjUW7mosK7SYSEW1elQ2nHUPuvIcZXxTmU0EKhaP8guPKoc2qQPt
gTxF47ptz96bVR4Z1vJa8VIcySVVFuVXAeENFbvBBgmIMxdlO5VDHHK+Md+ixEgs
Pll0XHVxlVDvVwn5hktCx7gHTK3M8dH2kILXddhCmiopcJNDGHyD7B/eSWi+EWfp
lRN4Ga+tps7MR/2y1CpOAMUCNkKNhyK0OPlE103jPle9jJl37dGiRUkopQyU3047
WnkN7Zkqa/JPtnrDLh7kOUziY/U36LB2ce9t4wDIEzR2qv6pSLmP8jStezvNX8np
TC7KBQauvVvw/QQARSm0vPbi8cqhrAI4OXHqdLJ1UUZ1v/zu0CeFReUfass1tumd
4P6ys0z2FeJxhvsl7JFOW3dWNP5GGoHr9sPWgpgUjRCL3j8B8bBYSxprgmCsG6wy
6cpfF+vIeRqbFG3Z/BD0LyOjRMBopIusg86xhywapHwCVmDN/2JCF3zdJXt0t829
VIKwJct9/lBI5PU+/4j8s6T+sncu6ihrgKoeJUm0E1gkMVtB42eCDDOUO1fWEzgQ
Ml4QQZv+tj1TDszMyNF28LnbrS3ueHHXjQSyigLT3EP7TxE8bYgPnzXuEl6w/gGN
16h43uiX6Ma1h4nGsLUX1nmNVBBiFkea5INmomw6bzdtjVvUaSYhpRZE17bAnsOE
1vjFf743Ifnl9ZyocJGne8MvT3o5kmUz4f+ok1KszPQx7OmuzYNHWgS2qSwbKFam
b4fpha0CRjmtGPbMaUrvOTchEsZKAgJCtEYyQXtcGLHjYJGSpfPOdN0ewKflqKMN
q/7mL+zSO6IyevlBZSsmow1BBeTvrhvwhI8x8QW7gUMpszT8c3hMBfberj0J+KhV
A0GGK5V1ZBfj75lu+IJuZ3YNTcTu4urEEIDTv1gfC4kkEhiiEKl5ooljTfr4PELJ
ziuR3ErlFrtzQRodKqsxrZ4+dZIGEM81e88qI5bBsOS4VxdEivknOusYkd98IFs5
Vh/4KY/S85I+UMLZZPXx3kYCdCaOumAKKz/H/cC9wEBDkYj3yRLqKA7iho9YBSfL
UlaumK167OjkRlZd/jKbyZZxKj7HjlATnkl3DVnito0HUSfrLnXfx294f0Ax6wUk
2mQh9GjC4gUMx6zczmIws2lfnrogbkK9q9sppIw1MNbEg3GgpZe1gZ91LMW64oyS
fb7FQAk84dzWd6mv7lwUzaBHSKCy0QaSV2dT0JlT8Vdn/AYFr29SHeP62pvx1cNT
bGAq8mJBu6+sYcgVjyFGN/KN/Px7rn3UQPMXGU/I3AfIga45DRMQffyiZR5nhlQw
7QUlHRgRmDQAmXOojOJlhkd7jayUhPn561KA/ssJ59tJayYPs5CGye7BiHY3Gqjt
XPxBIxlHgF+yEjBpzlMULQH+tpeyc8J+FSLugyl/qjKJ30zWTz2ax9rcRhUaIAMJ
6Q7HQxx2u+eiUj2Jnei30Ni4AdVxyYPAdyyegNjkHopyEnJ2WbXGY043n/nao0Z9
QhahnEOzU0dRdC1Ny9gGmyrxaGJ1H3C3NFWL3Ih0D+mDIc60frXs5/ja9EdnAApi
CB0a/FNQD7qbh5W/ozVQwufaLTVSGCygD4OaoQali2iZqp7fPSI+A+J/zsLLpVKI
3rC34sEbMhQbfHAtZo7iMYl2QRACyjWKYkpI6HxXhOK4sQ6xIPjLkeU/XOMbHvAM
ZuhKerMxqZcN0Efs5XleQ5d7yg6Kuy6bgpmn8kfYnfEkvQVG5nzUPDloNDRfyd6Z
icyOLvLQMqBUZFhZljLbYvKUapvAV3qCXrGpJeHVBclpNVFgnWLPEtxBwjCfdhqI
KChm4dSWuwjyqqjMLUdWdyxH6pO9o/8l480fq7WeyOsz0JWA6+nS9ll0r8yP0GWu
105q0obFeiLQrQ++UN/7gk5+t+y6k6JHJKtKQj0ds3VM877HyJPvJAC24OmvZv7K
MLRDoN5KtM0oRVSrNoBZxlax4dPMB4YywESu2cfXoWK1u+zUF/ZH8rlvpjYd74ud
q5jpjj6a0eBZaTNJl/oedd4kXCUpqy83J7wMWnw9OZEgtG9CQhzRACEfyg8tSz09
zGCxEq0VcsGyOFUWPyVwRyfnIGMOfx/Zn7E7284jnhJf2i7D8mGkG+lNi3WqGyVG
vnlB60DPt8AP6G2JWfRSZK60F2DIWIE/3wZRKIlUXy8a3EKGvJBBRAyIeM2YwJYO
vdGkMmkKTxIq9K9P1nB5tWV2+mLuwrqr5JBImGhHELhFJxI/9ts6uXjHDDw/lHd+
fhnZUZdSeZRWKto6+FnxQc1xzasSVu4UXtHaS2Z7h96Xe+0CIEPaE9WMzQStm19g
saxSbxyaKIMZ3biY6pGARhgebMXPwsKJTVAaATIsrZXGDUE06K5jzuRbDkBsd3Hr
dWMvLBfzszq39af69x23Y+0HBwF4qjGbmI53EO7Vk/wASF0Qf2CzBRUyagf45k1y
MESG0hB7oL8PJi8aMKivVSSlOzcO9cfc+lqqg3LCLYFQND7pevQMXWPCNltKMVMZ
B9bSkUjQITeg1Iqt7Ixl3qog8Ho0ca+ePlV9yidA/bYg5X07580dZp0Wd/AjcY84
ukLdFTztY3vYC5DTeyrKtaIfFsjgUdijQ8cZXLRTBX1RRxpjNCGwSWLyQ2szvk15
bSnwDFez7de8EVYOnsPuqPGZ+C7lxHCiAGEVo+eTPSh/HmaTVbmw1Hr93kciPtYb
4qi+qE2vDaJXZmhczS4EfyLeo2MZB9n+WuM3HtgRZAT+Ds+wYSiw17dE4kTXwGNw
7o8Yz3R6BsLASXsQQyckyZIVUaxif/kJeIK+gxJrlH4DxtDFAWTQxVhRuO8xB1aa
jLWL4PYR8xiBS4j7mQWKP7tRdV3kULVHJnxdTh5NVIPkkx2jIhQXa53SnyzYOYEa
tedXw8qY+IGxsevlcv/zcu2zSbjnG4HAwZVfXpYK99yESkPz2LshBOsoVOSXCMIZ
Z6CTKKy+p46Qs2g+YSsQQpO6nIILeqv4+fbTwy+WxjYeUzsQjzcCUIhHH8F1jvHP
NG0/sBbjouT7ST3im6L3vzMD5ThULvJu1RH/lWjvgfadvNG8cIisKhJq6tnU03Wn
4rV8X35lU3qxLfLVo12BMpxSDkcw6p7dyt9ITMsio5fd52od9ijtE44UJ2wQFuDv
X3/Kpf1UNTe2hH53Fuwepj56ummdbevLToLE9LvrtOq4ZlCY4shlPKaglgMQQKcy
diNKmKGTZM2YLlMOsjyu/xEbAWpjRdyWWTaEGxr3sEfxx/JI908YLe75q/x/hSUI
VYlcs17HXDe+ugB32Bm6FKVh+pFXpu4XLynp9Vn0O0+hzAzMN2P3Mn9tT2hoFstn
hLjaU3S6JgRL6S7aaUFFbdfeNjQIdOOgBZ/Co1FhH6DDujdFtpUYte9qtraVtMe8
ylrxTuio+MaqyPvR5wP1AzbhKIqTqtYbBJWSmPVAIsi2MV5XfV2QdkCPRFfoqmbj
f0wy62F2drURtatg4D/xsjVOIxLLTWIYglkekBsHgMkihGqNs+rGPk6YA/cT3O5d
IRYm/c8wxHAFzpceXSTb6BhLpCp7/l8rJk7H8GvQ48/YAJkS3nzTnZdSwtV5PhWO
Tg0Obqru5+GXPS/vdsw67agJm0D+KHgFMYcnGpehmnM5rHcsypWh4QRP2HMNsLy0
WXDqoMBZXjCkQUIwdt/ki3dfKm3Nc+ygDH0nX6gRyhO4ZwVJIGI6R8gPA15eBYr/
ZSUVQRaTMXajzDAiiWIED7y53PtFNZtOXbMbn54dvedEO6g86jJWO6rgPoHxIFJS
uH26bTteHuM9XS1skKDYdhdaKIICTcfKwlivXJ3yAvq4OLivpBpsQBiYQWbZ70FL
/8mXWx8nZWRRUbYP6I4RyrqjZMrFVOmjkecwvC6QbEsg+Z8Dmxrt9l/P2ESLVjBO
W9/Ve59XxzF1leJpPGRL2gZlR5muZYQPcur+9/2Xu5ffrcsgXTjglyIiJQTwL2e9
iyy5JL6ANsv4d73L1Rd+HOqe2y1LHiU6VlAikaidigp6ThUhJUEJKy3++hwb1A0w
ZY7bVNjM+vhhDmPlGcArxG2rEVNoJh9KVVLOk288Lhn9lzUBFz2AZeODE/eAWaR9
FcryYZ2OO1TeG2k/8ko1+bRB/DfV1HPPHSEgjCEKpXfczhI/ZOjL+umnS5SQkSFm
ak1R0i92xpmocrCtnO2SthFPx75QL5e1UCVrouKLYW3lenssQVHTTPYl0dX5WACu
HCPFTnlGiVqDNfXtQxiWKncDHH6B+niRDPcBu93+VeGvg8D6Q6C3nZd22u7pGurk
zKqaMhXViNuEa1szZNi/1C82SmMyW1gB10xZQWaA6KyQjrjylZkfN15WoSIO1ayZ
JPBulJhIDjCBs9/DL/t8yt89WwK4DpLuUlsaxv9Zw/nGIQkSOdGhfEBqK3vhb/mw
ezmlxGPQiUyQ8smjsqXkIDC1dDIl4YvVDjrR7oRHJeU+Bn6ohCwvRR9O30EIEYnw
pDm23vcXDE1DbkSmNacbTx1RrfWT8ffqd7oHsSAxJKwlWI2pZGX8gnl4QGMIX0GW
thocWYoaI4LBZeD/Psa5ZD28xZiDHE/7PcOvhsxlZE/06v89Cuwr4vugYDU8OCFY
4a0/wM2cwPlWtCbqf4ZRv7RBszORECyiiUNE3IBPNK7KLp/K3346G4aojterXECo
pXQ0P449+u9oNsWEBoOMas2zinRHV1AUfeGZLmR75h2Q+PsAxT07OyRNyTzyGpY1
O0sYIZRIXpQ8MacsgkAW0yxZc881mSCiEVSvWIqli3Ow0bMQu/RIHc+/nRvZTEhq
bz61gB75hvDIr8d11/LO8m05crFR0eE1X3UQpjVGeT4lpdXaU42VhwS87LjTljXt
WUUPZSHPqCqCCRclFPub4GGeumD14QZP6NJAht6yPwB4wjBh1PE4DykFej7gCLoz
YgIAIsNkAUIx2sKHKWVcBHWQ5WGujQDzQU6ONy+t16hkuc4XVQ2MjAsqeTwjOlQx
ZUQzSeSiF9Y4YJ/NZXyiZ5EL1tGcYuc9gEpQK91djhg3iohnEYH2JdT/QDnepBLv
SPr400mi2rkE6ma15Locy/JJT7nPcyaXqTVmq2r+Ps+zX7VU8MUiFeRAdeqWlPKk
UL2Fondvru2M4cum/0/qmFR8l45pr6CBgLzDL56BK+V1mJVgYMKVnW4X8C+VdC7k
Xz2x5OCU1HDKnfe7tkXahTN/NSOGebtYpGrkhtI5TeG2o1IEuNQj483sbRf2TLQP
L/cj6+ArVC14UGqNYbFIGvtnEEY54WszppTA8H+sK2Bs0TbYSFKK3Mid+GWT1zqS
D+VE7pzSGo8Hc3b7ahZj4PlPda276p+QNpY8g7OgJ8HxxuCaxAjMbihIL31vHJ83
PgrqTCGwsqwW6roZb+MziIxoBsakjbxyYQ5HKM6xkj4oH8vhQA1TMbtvwVGYCynk
MOjMl2UNOw6+NfHxtc1oYYUo4gFrzcHJY++XiqCra/N8lXscNLnNSHLFDCMhjWZw
7nLc1GoAHZMRH9S/qV1TTywffOVkpFj9dcU0W17Yh9vKrY7dNZcljxJAH4vqOu0X
MN8FGF3+aa9qrk3CHf3+uc6wxYnJYQhVeipzPhlVe7C9TrrcOJtbqMJPJI/0TiK9
KIDnXRvu7YeOzB45CtVBrNtd1zYUDLOIQnIaPdBsev+Hhfepc70K68JkXJmkR0U/
fDrSPLjWABzcI2o/M254OQHGHwgBm+ftNzOQ2MznayiCxjzxitAhJsiiCK25eRo7
8hV9toWT3fnDvNX3JAXpHLMeykEPzO0tBNUoelA9u3hWgu02QyQ7YwdKgVh8MFf8
6dk+aj5hyyRdYtx6pmoMHLzKeZNN+wkqJp1Ik4eDt53tAi2ovDWPVIySd80CgRWK
JC51JDnyaYzzGLkfQfRxr94/SNoNk6h9emcb9s1qXc1cd+abLM+nYcyjTHZ8PppL
XkXsDv1o0LNR8rNsYaNUNaXyWP8WIwkBqjVN0UjwXd/K+0VVoBW78h0PRvbGL19y
4/lirCTS6BOOwgB3LoqEhLoksHGUJl83szLdTtH8hFM7x2NJdTY4tu3GW+qWoGzc
graG156VkxiE2Jhg5mjq9mqeZR0/U17BPwtmkKi0cG/nrcdvglTgLWmJVHTe4DZe
YzWi7hSVnRh51bRlpJFe9zdxGwGNLVsaBUwKEGQi6WBAx7tWZ7GKSJkS1npQQwH4
R6fCoOnfWuPOplJarLXSiYoqPddR1tXIa1KmClLGreZTcV+buqUfq3n6BXitZn72
UPo4vnD9NsZoXKQdGxrKqCU09tTcjUotNWyma/I33Q4Dcw6PnsJHh4UE6B3er6d7
ehDXtGkJwIfWpV42JAaVoQTQFkh5/xKcxxZWfqELIFADy1fWWufE5YCcHAFueovw
krAnLS2US08GDOyYHD2VHmZKFv0uWybhbs8QiEw0bXjOc5hNr0USWfqqdJ5/VYMC
/lL4QIOwz0E4E1ifOB9Pe2gyh3D1hFEYnyMhm3ZQBBJPxp/Le2gMy4FSCR7ocdFA
q9JJV/ImwK902LQJa2ZhI4g5L2zWPuyNnRCpBpc4OP7Cbf3IFsxesRIYDPPOULBj
XZJ0KTD4w01nqzv0BuMX/TvZ+/g5QGLOlyY1rs4cjsn8HPY7vJXjiphCoqEuj535
aE1Z2BE1OjYjRN9IN19xmGjR2/EDoyHZHeCmm2yTEXwecID68IGtL6O1QVfMclr9
F4SlOIjPJWLEJ9KutvkyN2oLIk3nSDSPMk/wC8CLSwcDcaLHu7BM5zAB5naJ/ThO
t/yN4nfd/ydbMKelsERcCNoTDkKf18DNcEzclGFwf24yDEdIqBPJutNKaBYicYyA
LL+WhTlx3cDD4rg64wocrUugqQCHp47iG0hS5CRu0pRP5Hw9dGedaNw5ztlNXpFT
rmP45z2nezwRdlfQ7K3woMlrb8pYKYpwgCIswfsLPrkF/mTiI6K1OkC0emWyoRoc
fEkx9Li5Q5e4EXKIp1FLOOgDT35c4lhyK6s73y0ZHSPVcvrj2/yQfVGKCP3D54Mv
xdEASsO+SJg+ERbqHWUgmvbo3uqG1KCkgUxbgdPDBx3hbEFC5+tib5+YFarWLaHF
lMWbftxV0yLNygipkXJHinRxwTkaTJi92nRiTF/0IN74HLo2Bqx6paHnF1P0frKF
47g2DbmAi8vKcBU70XoeT0sK7dqhjIpD5Ro3EupH6M2EkXJRs1NdkPSN28Z1hA/9
II6u3OiP9/yPX7PKWpVnFrDaQLFcoJaTCwwipyxge6COx5JSHJ6BQP/hxdUh93QG
54LFxhYX0bsw8CwYz9gz4WsZKcA4OuWqLusjF+GqW0K5w4C+o4wGufP+5QUfqVgp
SGt8XZpqBIJ8/q0WD4y0NkOxOPDrlKBUx3SrBFWkGQ3LTqhGZvGdrUZvExuKe2hU
5R4IlI0XkZ1/LazuYUby0wchGzLMznRNDAZTrcYHm00oGE+XsZS1Es+n+pt+Vv6K
BRvkGYXU0Fr0SmkVGEL08ve4WGuqbFL+YO4CWgoQGOpCWSVTKrYGehgQH1qt/THj
auBiZQ2hEkC7id1XPC8e3a9jw3zNCULh1lrWdnPb2m3Xgs3JQAASzE9UlDTWXVV0
PzhJkO7WbpwzrMCDsXr5hMEJw0TmhmE5swTScQdxie9DAc7xnQDcwgs98YrxUkVC
w6vlifrqOZjVAMP09tz3P8zcX7S63S0wzqjhEwFvJwIIQVwMwiVZ3rWSgeLxZH00
v1Pp2RMX1u1YXp4wZNdPcm1BkcuQBqELrRNuyUlyuCA8VkRif8KlZZ6470l7PxHa
z0Lq+EmsG74C4+mNdOsK0c+GrsOTLeTjTgWLxX3C0140Ww/XJNF1wHmrFGqY/NDe
CGGBWmpAFvH+y3tVMntagnMJJntQJYOk7ZshBAixg4mLn1aXT0HaRC67kvcz4z5x
ll6QdJIu3YN7Lvx58aEbE1UDbgmOqdHsips+u0RSzGkBVwWgqGELSvpBAknFT6is
FnGfbxJ925H/M7iBkpbBsNhXTmjRfABXayq/3yHRW9+VIzUUR6eMfctvYculz6Oy
rhHzHJBqvLYSmBAuT8LU3nQ8/720vapEsgHFGlMzzljQlvkYAHIkimxE09QQXV02
hz9LSn9KzjllnrNKIA1qb/gPJw8f2ebLBw4J1ecJVIoUMsb0qHxte11UJrdaEAVA
OUyZ/AOgbfJEq+HfYBT3iM/pcTTpTjR6ugfPJTarCY5zG6bD0K0PCq/rHZ6sd1t7
VpzoEhg0Vv2jMG83+9xZF7eMP+witfttwcc3KW3vDVV6zztLExIcKp4GU10V78FM
CJ8BJjlw1JQZsrccpnI3s+hSFYHRstP4Rtf4sT+n60Ckc+2MJ93UPiooSVN9OO8j
IVJjVCTLnJmESF3IYMrpAVkECyt2Ncnn80p/E0SdJK7OpVprF9oeLlem/J3sQizV
SLYZZE5+9QhWomJ2FhPGTUkR62ChnE72g9D2zpgEd4LrVwlZoL192DBaJktE5M/w
lkxVo1KXfkU2I34E9MALC0U7rLeAH3yRT8G6kv4bLj/VPDAZ/t2eNZ7K+61s+x00
viOcpvKyC2xODtO0GA1IhZggW1PdxMPruaEbXnB1i+7PHc4TroSKm/zyBbuInM95
3xFigdlXaWW11uYWXHixgblEgUAe2TkrTqVXDsMt285DqcA4yANWey3VnxzrR7iS
GsOls3LCzleXwTdpzWmAgVLVu8q9eZT9HVZh4N/jhz3lO8XFgpHOPu2cmixotNhx
27uDrGy56YSPzl1zgE53hn6SE3lIl7I5IX48xOp5+Xbd5u2+v63TNnfomq8S4+Sr
uauowADjM0/G+uxjXVa+uuTcNP2aUwHBUylKqaIxzpMuG6wrB3TzRdBhnIq8n4hs
WSVlJSnLdu+LAvY7z6sKpJbiDFLTU8ERyfVxFSkEhtqKkS4ZTGfTHc8qcb5UZmDB
Th2lg9r4sBNwabwSqZa9xKFJCUUNyXjjzgMPwwqPeEVOl5B0jnuuF5uMnYvWJupn
dpd/Ai9AA7vjpRgeKHxeAR42RE0UcJXVYzzwYEzi/hf4SNEVGdIYCN8U2w7wwoFX
NvrnPO/j8ChvPTihcxf0fAFoQ2jzXHD9bWAdIHkwYWTaWczuQBXrLaVZ+pWLZtwz
UVNPghHUFkxP841DMiwFo1L7VFc6WP/eQ0YBrSLQkMKH2hlQs55N3/5g2fca+Rs6
uQ4xMdIeK/xwVORID8xSRfxzEJBKu4l+ZlJ3aTcyP4o6h0zEBZKYNkgdgAF6M6PX
YME28Hh248cVynQxXKcjvgyMkDmMl7lSx2O+aDWk4ehhlozg5fYJR79N9oj2rMzo
/m90iKoFI8fUVnThqTTbrIjfcmpoOfReDj/Uy2QLi/f3EmJlO/d6CijKzPIJLnOl
Et6pFoEkSwWfApepWx2xX08ll8laF80+80IbAsJkT5kgRC+YY2OuVlK3e19lA/jC
7DCdEi7yA6lJoDtXi8lW/9M/K7vOEQNK+Q44BMUY5raJqnwHdidWtclKhfuSslei
TstLGDiGBMa2l3Fz62MB6pqwBgxW5KQDfchqMQOC+ihQWA/q35jyYsXrbo5UMzXz
Of51+opj6bRWvedtVw5y/Mv2R4KGOZTa2kDXQTGZtYVSTMcLZ06BHiUBMcouTRVr
ppZevl9O3QVognrUV6aqGDvX4XWn8IwJEkG/dhXV+BugnEzUx/jCgqAxYWmpKY2y
07eXeyZZS+AO2BLjd9O0TnZGdoSFR0Lg78OQHzVe9rGNpYD87kdUowyA16i3c4s5
biFAfB5u+vWzPZMKg6r4hO/gHZ35ve8sM5hTguYsqIvlAGMX6Z17aLjSnmmDgjSN
OUjxHouvQ712DEncVTACOBwwGrX/2jxgYpUZugGxgWY9DnTdLJFK9bdtlHhEHAvp
lQfHI5cR9cvgHqSms5azyw2STbHNxS8+5nHzBfMfbWAbISmip0ooHwF3GyCdC7+C
lT0dTAayLMb5zwrQH/JrrjkvvZWRTiQ5PHpO1mnKx7cQ7Xy14TwrF9Cc+YRXOj+0
YTqTbzFxAX7kxF6Zqu+OxaNmwbjp4L+Wd88KEKN1vjO24raCy1K376FcluEyP6TP
DRpsOlRyK4K+gZS/n78wBBhoWtn9+FdmOHObff5AsdPsCBwv0E4kIEb87FsyKNZ/
I9ozXkrkekL8T6zI9u21aGY+OpDo/owkmYLolDYGomFUnSgSLwHWZMezhfCUHKrJ
V6zjRzcqw4dSoOGZFH9AvvOXKpSCOKswekYy5Kr0grWwLtsSMon1eCYs9gm56Ef/
MMmw1u5G0XCvX85qjyj18skP05JEdhgKs23OnkmpGI5RNqFFWk1P+u732ehkrbfP
vIBQdhbkugjFxgyhy2MGCtDAivPHdBzkf6WfexFQ/Q+AdVM/sXNAbQRuLKMHrUx6
FzpreAg+pfipoAMFUXgG1w2jMw/xz1+Zsh3r6MYxbWDZ0uJG4T8+PljzYXxOcBPu
L3YfQ7t95r9YBd110ydKDpBtvrGQhiowYyseqfO/Xzy1ukP4fJ57YgePt35eEXZM
VsLFisiUXQ6gjlKbBlgFU8XaaihJUTBIdSZt7rJLDnvJSBOeN6cn/SdU2BtIU8Ts
eZMOiledaMMGdBW9C3CUTybh17WBL8pzmRimj/4L8tj+VJ5aIDMp0sTYSWsE0HDJ
38o7p6f1YHaNqdKXMizboO6AMHpedehh7bOlaD6zcgQy57s2bp80jUVqghFV9IV1
+LH4XwHTBQiX2O6GygyZ4CKAG9t4Q5nQ+CB2VS5IkoVEkveRwdoIOl5K/Uc2W8Sv
UdH9oUfpise9e36/t2O3xDGwzoGb5lG73n8ApBg3iY/XNXTv3x6QFHkKW1uJtdvX
LwD7p+w4dGtUU6mjIeDRVFoZZeIa3Unth2cEwthtAZ8Ty9bNkxqH6W09X04unfmB
Qg6nsbxpNuAyEV61vjyC04DbZn/9kikX9akiZEdBt18aJ1+htbEjRfk3nO2OddcV
FrdozTTNfD3hsL+IP3I4GTQFD1SGwqTC8Cip6ANwtNzkrrhv6RtZh4SyUmVSyZmI
Qr6zKQnHcgOTn5/6d0qHj6Dhvc7/qDoYxGMh2qSeJ+WGmkwGDOS1MXQr+dWhgN5y
TXrrAWDtjvzOftiNBRFoqBb7GWfoEgBPVh4K4ZxG3PmvGRE2Sh3bV+8ooXuOTvHI
gFOJzBZolowprbWNXrGwyf38tKQ7dxopsuTGH+gMWbOdP0EGjCvJ0bvjc3JupXEI
C+yyqxsE7vwRKj+4aaVTf4/am8IxGi8h04oZh360UlMWo4hC4uWzfg66fiXhAccH
Su8AfehpHB6wg6v+/UuBQgMXThqJH9WvCWXdo7K00jwYrhbsw9Ef94XXdXX5c1WA
BFs68yQv36z+oSVww74Cp8QeB2YNRnp1quNjt6hiQ+RvMwYbL3nXuMPgYIckZQbL
eLw4/LadDJE3tzYtD3dXpYvan2qPUMEk1CyOCPQ4MqythLPIBp3xPGFWkITe946V
ZO8ODLJvliadJWnJpGhTgrLluxUWPovX6VsaqoZ8S76bBnKDVTXIVjjk2WVHK2W6
BNrdSd/f0r7y7T1xsTdBnb2PCfMCqcK7/j/37oPxnaKRiO+G/jT47nCkOZ0JV5Ux
ExYYUBuQ6GLkxqV7HrEJWqQ9cU5T6MEfALwZJRc2gi5izk0zEFXRL5VKhFgPEvpr
XVdBV2YWvN0DVHCNiwxH7SHsnIx4dcFpHeGXHwyY+TM6aZp8PRor38SUSD81LtRR
VI2FCXBcXNzgX4VJmFCyHuNXbK2nPMdxCNlka/vLaLJymkzxay0QXieFYCl0Ffc8
jl2ZMlQ8KFNtYwIRcLIH+VvyE34g+N/Mp9wqkaDMXJWGG5xgNQvb7URmT3J4CoHI
OPqrAyzlYMS3qaFKQAt1LWi2xmiNhIGdFiEdOqH95CzKweTjIWy6jz/1pJ2JsPUR
JsZXbPfgS/7UBVWL7KRpWoeeh3AfmtXU0bP7+/GoHRcismH0fJoWFnTC2w4+ISfP
fr9Sp+kK5FKdbychGSbRSLt+IsJ2dveD6d1LuB2cwVVbBfc6Ujxm/WIUcQIEhPlo
DtpBnGund/nVrZllFoCoMW1ibBC/ulrnLofqTtgpjVZsUFB8CUXFpPrUh1/MuuND
Cd0VVqiIBw9QTCaYgDPmVyr8Baxo02bwVDdtaAjfwBCFA1/3zj0509HCaeUoTzfd
tdHXndwMDzW56WhapzPeyNDHh5erj7d5mwL5nUxmw2bkL+E5X98VthM0721GNv1Q
xXiTgKh3fB4Rki1D+iAdeH9i3qzWgJgMAPJidzoJgS80jsa2fgzHuT/tYyrpeeld
k8a8Q5bC5qlsL83j0o5LTiOuZ1+FVjOIvZg8PX/IOSCCLKzo2p6Sprfqf9aU6FNa
ix7l4sMobvrlzLVoMS9hX5epurSfHUkVXwL0QDTpD16jvoA7ikq0A+XhoQreOwE/
yoQmk8HBTEkJjOBhu4CyqjSW6vFAckEqlUxNLh+OgOdrzas2eV5/EM1nBcYcc6zS
E3XQ/l92qgsPYI8545AawNy8OqEbrlDmiGrMu+1KK95Ess8/XL2jPqUCcI1RBdqX
zL8Zvzzt0L9Sil7RCsdl2lgJmtsFTpuQCzktb4ZC8nJzTbsuDtNDfi+YArLlHKgQ
h/zwf4cB4hU3F3xf0qMqamxyTLUlL2oDzmWn/QcEoObO+zAHIdn+eK9LWUsq19vi
ZeRe98GkNdM4OWZp+kM4zWTI3XbCq9fz2XNFQ8or6XXid4YlTut0esGmQdKbUj97
pe6plMiliz3xVsIwytTdmHcvUnrtcTWEcUdieNbDUurMZn4O6ENTd899czt47D5D
rodi1nEyXI9vTQB/l9ptpk6Vgu0uU9nsNHwTt5O/hxge7UdwTHJPCDBThEO2Qt83
2wxKsEwp0UoPoWTdsNBGuum1aqJt1/mok2XuTvBx8ldgiGh869IcZa6HhkCrim6G
UnlmSoKvgJqJPRIjxqqFOTx5CL9bIBZ8WJHzmC5rhUqofKX6cg6Vnk5IH6aksqPm
CCfIWtk3Aw3GfJD5nTX2X7XtBatW0Lksk9hLNIFnc9c4Wjk4ErMSwlG4qIyxfkMH
wYe7NExXaMxV18+4NbshmdLN0XwF3b+QzZAwqSZpUPdO9bQP5kEb3QnqfcL7BvzU
8RoBqJGKdr3QLI1zUMiGJ2MdqibGFtuYsFC2Cf/F0lPZAX0/GvUNG471wVRprpH8
z6UkPbeSQkJtmY2vOq7d7YC4i6QOiRCbDq/+ShBqw0qKaZwviwFt+g5AlZe3oE9U
rlQntf14xNgJOu2VEbTwC5D/TBn4g1HSTsAzsi5fYpX9Fz+yxYC//5CncqUdqE6T
cwF/7Q3d8Vl7Io+0In6TZ3SOX7S5Ed040eTZnmYlLU9H9TvqytNp+DhwnTIm4/VV
8hDC+p+lYSBBsQ7DdmqLz/nzgqKo8ANzn3VqA+wXbG7dMQ2CslC4MlU15Uj+DXQW
9LABbchPOKUSqEf56QdBonuv+6MgcS7dE5k3yoW3MnM4LLHmhSvQ7Zlw0OKIIkcm
jtNIo/qDBHX9YbSu1glXRjr5vExIUdiDlfzK5kZPvORYvTio2dhhjCSaPhGUIXqp
bijkKZvB/n4001cwrhzxwDHDhMj4dUDWELk+gJrm4rX2qop7TrDbP6PUQfGdTKB/
exPbODMObclnDRp6kgPdLvqxcktyUauamvzUY6dRgX+XlopIQ39DPvuzY5FHNaoC
uuq4LdfchYg5F2Q4ctjy7H37P0q9mUVB2hp43gUD1mqKg15ULJqj4JTsMvTYRxjF
ff/vH5EJoPPo/7FWEE5OsBX8unc/wOiYQBbT/cHOZ++U0T+cGYKk6RfffvbBK8Sc
5zUaq0imzsMxxoQC8wPVIMAG6j9SmprpmciHyixBsUau9mpUa4w54lmS8MxHnAgY
owDAWVZcgIm1DRckuBVi+wgc9zis9lH34qYuBaDOiAE5ifYQ19kXBuFprtA9PROo
NdRdO3uhUI7J0Pn3BocVswRYj3SmkawBsX96FLPAkLli5/TNitgtha9isJH88uQJ
jQx4cpA4DTAzXAMnsEle8CHTStNdz3JkwtniCl6Ugx+fwd9rSz1Aa5doX1gHUzZ8
CZPvt8ojYqpl+ufEZ4JnmcvDsIhH+nIBfD50Ldu2jG9gFtejp6VpTjeRcDJyWLU8
+jjlrFfZLxXZ2B7k+HHa7rgeYm5PL+HQt+NT63rNMwqHQCRrmONjznNixyZJ+fdY
/OOKgCYiRMrVXOVsTfgqQnxQpji90w0QPHLudbOu+cYwWKWf2CF4kv/tgmkz/e9s
n7hZ3dMfKi/q0bVdAtCA4V7xzNgV6RtbNcPtM/3h7XnUx/iCfW8bty+W3mG6LqHK
qQDLcu3Qoi99uwkxvmftxWnIYvWUlratyt9GmeFrD9iN/4d2XPlOP0cxMscpiQS6
TBgWANM96wVE732BdAP+lAt5H3BYhc+ns3iS2XjykthmTPudh3XSTQbhR66RSoX9
XRT9qDcAlo+NW0QYVcAVJLgaaR8g2cYdOj8LQyYyt7/R6Wu1VUg2Z3zdUIYb38nD
TJDn4XSUk14IBM0Cy2aCxU3wMjiVasjQSmrEGFLPOCH51+9Gwu+Qj68AKcBQ1jph
cyE4Nx9CKAZgkuEVFXVT/CcLzDuy2iobvyYiunGUOMvuRZeCc8QwI4j+nWjl8xP0
691FUMOoacmn8Krc4BJO/PMIhpG3MytShHI0bb9gZQZFLfKB6vemS6e8STJZRqEj
k0FwGZvY6e31x2yyJ4JlTtazZp7u2ovT1EDpZkArs+OQJdPSN87CHKJpsfHoGID9
dim3AJEv+dDVHGrHLMSPFi3RXRlquMLw4DVMQ6goQueDVAWd+o+t/QFrIsUWE53T
dV29OWTfiqRAcwyZHNCahTShkZFVHLD7fSoQSXDYZiWYFXhwhUNrH7GuZqJLk4bS
vKY45adh2DA66ags3GfPrFehIxMeAwiibK8Z0jnqidAGRkC8roUae4GDY6T6GEfO
uxZ937BaHhI4cxnV1SFtUsg4fdM2bLL51YZH7aTReI6u8HCrfDIvFYwoauaYU4fA
C45HcWBKTZaezqNMC/qG76aP7CX1YjriQyrD/7dUjRku+Px+se/PCl9V0quFotei
Mabo2FxYAngju8N0CogACffHBhQ8awDpZCCPu6fjTAELnmC09jwE76/S4G54gy6h
4E2kVhDaQBdRsc/86J7N+WrmYXjNFlt1enmFt2uaIHc5U+WhDx50QkIA+HviUb5X
oWGC/5ky8IdnmxvCxvjlqvZz/obrR+UBkeI8wqoxIJdG8eYgLuXkACMGAo8CHpD5
CaX5r8KF0l9Ga77bFwiG8+q+QnRn3PVG3vqNQ1I55/HscdkK0/GDrhQvQgxgy/F+
9ZHFrgdafXuBZD8dMM2wP11qZFhgqIUoIZDd13L0CXMuoq63w6gQ38X45I+Ej7c+
BMB6O71hJWJKf8rMy0hy715aNQDxMb2kGXiGIi/wMxnX5IezxGkYU5/H2i0YhzoV
1GaGsGPRO614TZOm076Id7OQ4oq6MGPqjcPA74LZ9M425kGKfckTqPx0E1licBbN
LhM/+IdY8QYo9cdsHahQGsWhyuXH01bW52QYZ6pcCrZ+H8qdV7S27UCv2SODZDW6
kgan1Oe/yHb+Dwnlk4qUwZQ7hzZw1HIywv+LdwONvadcoZW9sx8ewD58ItDn/DZH
dahZ7JBmqRskMA908rczn7v3sAmTd77nCOfA2X73P470QQ1BmGZ208b6ApmWh1CJ
oXxOXzgQuZSp5Qbvy5aXblgqmskaFZr5bDi49yLgyckQIdrWV4gcyUJ0gFHW892N
feOvcQAfG5pnVjb6HO0qffABlV1eldYCH+U5EOq3M1n0eAOG5YEQhrbZBMDEgwE/
g323ufnZ9WzvrVNVd+W1gWXTedCQig16hso1qMYxBKeGZ58hnYk2oi49jOUIlom0
C+i6TA6Yz93M2oqOalpSNR1ABHis0e9PahCXhtkygk2D5lVLflM4b4h55PxoiXBg
93RIZKwCbmIQiLKwCA+P3IWdIUO1HNZCKT1oNNwFgSIhKx94ZfV9Q9YeAiAYaora
96tE3nUWd3FM6J66GEXYR+aHXegaeSLrq+R6qFgJX6myk0/GyJ7Opr/jdReXzap/
HXpkfilnUw98gGAE+5rkz09capuNRycKWXQZ8rIR+33+P3WsV7s3i3ZaD9xc46NG
9zKh4qIGCHJAK0mDl5UImXekg3KcUJdaxk6a5f4OhhTaULIgfhoxcl98vC8d4dd6
/dfTesEM4PVKOz4sPCqUyj/Z901e1nhapyv/nhI14khXQ1uj4aXSkAdDcwIkFP6G
0BHI9kK/aTqSAsbs4JBg5Vn0336Fr1zyzV86mxr81RAxXRsGEZjSTJLOnhqoE4Tu
aeBulIaSe7u0z7cjMPQoHe6EBgmnh4iSQ40of6MaRuboNiiUSftR4NxlGIIUL5s1
J/9C8MKQkoBpRXEr/yQ+c+TBS8JTvv3MDmmMD2Pe1FpZwJOarZJpZsGmQMEcpPtt
F2uAzCDVy0s1mBu6E4tnEsWlbiJgcV8ZOvLLV27VknnpMBNnMo1iQWLfaaa26R5F
bY+VfWnRYMoUgTA2y1KamD019fbBFWPZnBfU5DqZ4p19+sVVFHL3B1DL5ItosjXw
7NUEHSSdquc0ai41I0Ee6Ezl8dCytD53i8g+xwwolCm/OOmviJC1V2pTeZVLCAY6
mCOyuBErvXZYTMA6vbt6SCctRDO1Frokscl6jUyQn6rWHpEEI07qDK9163uQQbvw
1ksOikn8tIas7lf6txWnkLiYmtKzQGLx8mXnCYJq4CMd1OhOkkLwtCf1Wq7N1/Aw
16jlsZR9yIkqc2U1bn6bbbzaN2JloMf4AcTRVfOD1H7IckRWPyQcVUxOyHcrLFya
CUoHrAbChTdbn68DUFi4UlY7au0XefNk6XZwVNgMjPGvDTjTDQQQWF+RpWOwDicK
Gsxkyp2C5EZPqfVmkxLNEIIcLyODP6De91dZEs9xIjqDncALu3qeJjUujIDXRhTc
cFzJXLp5B6lPq46kHTA7Hnq/jNDJxo8nUW/vJRU9ASEoN3cVmMsfV4ckYzq/pOZX
mOg+I3K6XrnaSfLH94bOnu1W/Y6MBfqK5nj21qLL7ujvdwcZa8z4HDX0lEKNI1TO
ZrESxIPpjW1WIs01tL+b1PCDeD8Mxjhdv/PCs0f78QiPuG3JSwn93P/YD0xknkxX
MqMMc2ldl+DW490gpyGVZzl0hDMWHGZGJuz2SYqZyHj5MIhn8CJ6WfbejMXZsP5g
fnN3z0Sj8QxVqjrILSwM/jPRLA3H4+FTd3H+/JgJDDiy26/vyMBrqNJyemvB0QJx
eYRdFaWBDAmfIq9hUrvE2xCCYUgl6NOnqIi4Y0GcSnrdKtz2blm8h4hy7myEFOGh
/Zy1qbl3si6XhA8qekc02zLrLGGZO3UgV/JLLJFbuEj9jDiECiYeG54Gk7wb2s/d
PAsiwGgbPHdSjFMRS13Bh6lVdBosvxUGW0znjRz7alb5gZzTDYIY4b4rw2cxwT2I
buz+Angd/WG2XU8pEjBLEHq0tTVuzLNikUFvyhqUYW8NAB3XFnVMBwkKEvA8BBhu
QlPT/8zCDyP5/z9f0CwStoIXJ0n4lwXuMKcOv7WE69UnVsEBvrubBwzswEPKvPQ/
PTaIckbPWzsYHZ/y3nmW41826leecCv3YgdkTfGc1oHHCCEtF9FTPbM+Hx+Pz4Nl
R8jvB/nU1C7QaF9pRViriXW1V68xUA6BOXO8I1/ACoegLL+Pnf2ozQc8qhwF8Aaj
zf59XZSzILfTSLdEbBh1rrXf3+omLBIbgFpAOrw5ax2Bt8OpdhXEagQp4T/6MLqb
zCJBj03bPjovEs54j7W/rM0mFz9jCNUVts9zwUlfIVyaLVOCjL7qcSBtNMN3yb26
ET+GDdxQ+jKKe/EZzgLfRiOab1svrr1rxvwoJHFguU/HzkNQSp/4alhxt5aWmKqp
AmPZsYbkMDAyDhfPYIfbz3zuZOZbdEJsBNrtVGv1tGxFzZk0PPO0u3Vw4TtMuzad
aoUpyVky/I/S7t+g85hcIXN/j+7zE8gdyZ84xnDYZHoKQvYHmyDpq6Av0tB5xEAQ
m3YxxSbr2B3W2BLypkvX7z2TsEt/3YIJxsP48N+X2jX5v6dD+yj5KZYT7gzzdDxc
+5+Z5MGSfreww6WBnpV5qOnfc5DaIKNvaeEAuBWeCk5vp5BC34G0tCJtZ7E0Bsov
8nEYLjqml0qTqrjj/XjW/43IxoClSQLgq//zIgdC8+dtbdGOYyHZWxQ0EJ08AtB8
wiI/Yewll0z0lhENTDr/YIdRIe9IuSrSmKGfrqjVg+GHxUOzOliDF6OjW0qCP3YI
zLMOTpcuO2cxcFUC4cJl5c5caUNq1Jtpzto31moyivU9tBjKSmXGxfubnI0MO4qq
vrZtGlMotJLknQYff4ls0terUaxn4yzLzIc3DkKo4zVKJfXyw83EwrVAvD/dOiZX
I1kYRk4/MqZGieASO81ZSG+PzHbbNxGCB+7PC1BdWZ2Gbb/8wVaePj0sMUUzvrGX
jmPHqncWQROj/6uegZD9Bc1OG6hOglo6nqXh8ICF853SaYysJf2layzqwloEPzeo
nw4qY3JGQ5OAhgS460BR4yd2f4xr1J/4+bGwnqYR+9euyq9F6LQiTiI8UvJq/L3P
CMqINBnpsrL784v1rm3kM9CnE2aBkX/7zDbSPbGEAvnRJ/XrWtEdfXBv2GkBvj/w
FUo4aqhsWKyuq0eiyZVDy3JCFVHYfWgbsuZZn7ZnrdPZphx79LDj0CiEQkk5tBGx
WcDYBCWPbVSNvSm3llUHZcRQ3eHd/FHSvP5NgHIdFCb8q1MfVA/BNygUmvLw8Pn3
yI0PzEoqwFqWffBcavZUTViLa1g6k6VzHFG4pWDOZD+LuGyq73iUChWo8BOGy6+3
kornRmYq+bZh/s8nSSlwm9AUOr7cXrfNOep2yufmakp3B4R9Q1S4RNOzjsvk5CHV
nJnSPMO/tu8cN1mZiXK2ESF+K4ztHOLcXZYK7D439DJL51jigg+3Aqc2/O91KT1g
sNrIpsj+RBdp1B63YlVAOP7CYnctCoN1vSCUNRxdiWTGMA4AL3KdRLZUYdlKJ9Lc
AtpE0HLSqZMNhdeZmBW/w0+qqGHA7tp03920GPP2VOPVdmyVStFhO6YM0u6MTOKg
s8jXRG05VIXfGTipu2KTBlCtzsGV77ZbSCbgN/CnFdG1qUQWE5VMIvaGLRQuC8lc
09tnAjG3wP9FFS9x5dZBOCBX5Ec8JHU9BOUVCW4vvobKMpQGWYWLldoocwcMCRZo
EbcGpoLaLd7b4LrL++UCQcWX0Vk0O/MOisxJgoKAvzBDJTZdnIT1nHSInW99MH4E
e7m6FDyGCfAw7tRm/cOMNj/+Kb+Eu8bjhOKjuy+o+loFIbtNHIiLKs0vofIdJNp/
aYk20nQjCyvRcV6NTJeqa1CZgJ7fw5w1+8X5o5ll0zWe/t6d57XkL0w27vGNO8Fj
Kn6SuT5MlrsLVsyZFGo388dijYZKNVo2RWA8XY5ByWf2vPMUaXeT7CxChnT6ic2/
1J3jHyWxwVvOq52vdiL2pz9LmF8OMejI8P4lKPVRsKbR1zi7nu1QYR1Uiv9BBkeA
Ui2sc9X+egCyWAgd76eEOEy6eO6BgS1NbJzlUXEpsTE3LnvUPPvXScEKYzGhLQas
Pc/2vfPoItZy9+6ZXWcz9EKuGDCpxR7pmmarLGVBhzlQNPH0XXd0UCosijMUqJaR
1OWQGXlETegnBDuq33npdTFIuMbsGaCs1CxmSpzXfLwA1GLYJhbV2HVQEDF7L/8i
bF7Cc384EYP+zOtBF9aGvb7KIgI1UHj3yV6XYBn8l6MURAbFLT489L0aKfLXfJ20
mFsUzBL2iNboBSf+snqCMNQAeQ+9qcorqew479hmWt8VB0oDAEUp7zoPgOejTjLE
0Yk7p4aXJRsdsQ3pTTTehl32A+anGbbiE9Lh7sZ4YYRjw4gAN5s/9iBfKvRyJXm/
MPAYAg+7Ceb4IKIGhPy/Pit6h137fogG23pnS22R6bg2qcKc+dLQxaYTlJtSbyFu
PeBvIoZLPr3k6jXkVIABGbHxOGYnGNYNsh60Xm9ItYM/4BlsSB8zbLoFQKyiuu+b
wsgacVHHt58EY3euPyyJoskKEZfRsUMdr4TrPFtz+SvAN/TyCm0RreIx2YvBkn/6
0nvogT4Ulpvz/gUuiiDhSScL97Gt/1/xf3Q5UpII5SIgzH/xL34zeEEAiNVGCcBp
1/CwHNYoMXlurSQ6/ktt8+MpnAn8/A4mSfK5GEWxi25JFV8iHcSoFw6vjS2riVn5
QEiPUdPXlDqVkQYwKvFZ+7BAfgRrxZDWePc9964jImIwHjowrkXwFvKTENFWwgmx
LjwM0FAjDqScVckofZ1qcNOlTMFAk8WQQWidzVhT1iKUnJJ4wSJtoVye7ET7GNi1
XpgTZKn6f1s+No0vPo0HimLCSfg23tmayOvBQjzpFU1wuID9aBgq2Ok2S2tRaaQe
EptzUNcEjBdKyTuS3qpwsZxmD77QyIDgsSNhqdzqwnIftSu+sTMLXIzh2nbKyIER
VajJtHACPQ2WJo9miYn+iOU186a4h+FHwCrRW13XK8kTWKeZxm3La7DWDYg9ANTV
+pyeGhD3hL1d57rjqOjj4EZNmAfa2Lda5fugf2kZcuMvrKINJMH0o5JKNEucLHmt
2e3h7NSefE9X8aMdcEq2w+twNTl7uULYV3b3AhqvzAx0A2P3QO0VyF/nPeKTGPpr
eABIZ1Lojlqn0sZ2fZwB23hZHfvAqy2QSJidl9sCzGrlSYjsKCwKnfJIETcMhRMW
ePYs/9thQoNeWiWpcXPsrj0eEilz8pXKTI9hnqX77FCg5Nrrl40RJoyjs055m4Xa
ZUbOlcc3w+iQ3VpHVWenIDhyW8RlQhWGbPabz4LKC8dHqk2/dF4Xrz03by+GelKC
KlyHB4tzUp1kwuPzPUaJosyWICB5vfBR7kff5MEUZW4F1ck+FoAFKocI3LMcJyPf
FHdeH93s7wg2Ups6/j8jiFWwIZbxLYxrcr4lCxvZ3XXTP2HLC4aojNf/W7qV++qk
HZ0Neq38kOVYfBIIWiCCxK2cJr0VSdgnBFWUepSmdy88OEhFfoFId9hM/X6/3qKX
h6Dgl6d5Kv9LNwrpaEXqZHDJbHoiVHVNecmx6oQpRJ2/aymxyopE0x0nb7Xs0X+J
qNcpfT5XN4WQNeq2AUt14D2/6b1nqU4VnrF/go2FBC4e5wNU+8rSRRldNshdS7rV
RIm6JgoDLPCf2i62vP9b0ac3NX+S4bk+hExtuEELBRAzmK4F7x/sByZHiQueA9uI
tAyavso1KOBKQ/SE9JVm6AWkuRtfAcfRahvh/N1CIrdxeSqoiN8zBu3dey9aBkZV
fAN4pgEnlZeu4BaLLjFSekWbnrACvUuoqHIxNDjO5Brl7uyA6I9mFBU52OwlWAUL
g+BWRaBqFXsfKoXKZHd00PvKrHJWIUfZyypa6oMEsJBFQEQ4bDRHuyG4rCHGRDun
E0yDokBNWlirn0G0+4ERDqigvmUR4LQ7FlfzZrf/z4oOM3EPpXjwgWtsZ/Zrx1s8
v5XFAw5d/Xu6BZhOKR2ytNVfJ8MvjUAfu6B/5bK0N7x1JYXnwE08hvkTnN7TIj7j
3zu8RR3/rXTSEGnV2SNGWRQ45cu31Cel7MhAMIXvP7be+kkf+W2i4OuV+fQ8Z6L5
j3Ef8AJMh5NxiatDAd0dYSVrd//qdzqCDuTa4GSTSiHlL3YVHLFVd1awG68GsXsJ
bVROZwjYTwlaCIJJcxdLJdl4ewhpd9seyh1DTL9h06LuSbtzcKp5oSINVGy9bZfo
TeIL3MjABEOaptPLOpjzcs67GVIpw3mRr41hOJPQc8v938UqL/aD7zAhcDpA9DAt
ta/m1fmPnWk3RVb8f2ahbvV55sLwDMstHyy2EBEBIWgEMZ8fS6CBaRNMtZ8Mg2NB
sBKgJBRm77NXlgIzmde5HhjSG+ZOsj7Qhaea1gh40xJl4APdGmvMN8y4DZk5v3gq
ICTTM/D62xrErabpOj222lCt5Y1yF8hTlMd06w5NgrTbgh8NG/aNSGwOw2NEHvAg
Cc07gEzyPgGzbo8OzUtmMjIkrlp4GuLPJUm/aHZEwEaNVjYrsaks1JgaSjCgf7gC
3+no1Zg/FCjv/rkGMiUXQM41KaSkUmMrxMmw2yqjYqCYfS2nBYyTdnlS9IEz1FTr
zz/4XDqVfLUtRqXVbZ0edoVsJqCp1APDjpbOYOYGeWXpSpdD69qF1Ly0K35Tcfm7
no0Sml6rZc4gbfIBE+dxqbdk6X/LqbHTkPVSY9v13nuArkM0nuaLwBuBbU94ru4z
2jB2ynnk5zUEIgRsi4XaCUfUOblNfKyTCXofev2S1FHajNJvXlJWot5qmBsyGhwN
nuUXPZnAr7JTmdWY4V9WFsp0EBSJK7k3/nJBPrgzksKkYcfNNtTODFzy30eSUiqp
oZjsAKy/jz1j4cCrBeq5JKMqVi/iH16p5tJhtySCjOLAe7B6TYOAF9E2JkyVjGdj
WgvLWRR6t2PX/Ne+VQHHJcFNbWRZJrIYVVeGNC82n1w8V4sX20TaKKZpKAol27cR
UAbqnOZHSEtcOHNZZ/y33bsou2n/sCYRvFnqrRrLWsUvW9ZisPt4zebRYppkCwkN
uiy34rOSnxVlfOa9mNSgZL8RW8fWpzUre/0vnig4f8PKiE2yrWebqEFmE7L5PZP/
/glSr/GEEH7Pv4WU4Rie3AGGUznSsmqMJOsXcNqver1elWAYkwt8QQ+2yfyeQU8T
6PSHEzH6BWLuGGcrE186qYXX2oz0GVi/Ocm6DKIUk3WaCRqIdVKpZgXf8ix2rzN2
qrMyk/DM68oC6oMiLW2YDMU52onWi6IMQy8lC6kESBHJlWrdsdOZrq1CI+mmg/Sz
vFzR2iR1M0sKaTGPssVNR500h0OCenff+PIfksfGelytTDgrMIBZ+bC69bLJt/1D
KMRbNs66yzg/eT3AqLzxbzawioFiG0m+s6DM7FJlr4tGw3aLVjj2eNK81ZCvnRjq
X3hbIbW+UKTD4kdQ6I1ZJX9s4ljzphhwDYQKUyXOhOKSnQNhCqWi6PAookkmhuoz
rmWkGqKq4F9ToVPJ7znjeCaTXHOwgBrabpuvacIZ9aYVgZJDYAq8c1ifZ/3E31Se
GMSQVRrYIcnsH2Rp9p86VlytTOtDpGSXfvtaTxFTcvERuhtw9vy/HCCsQvO8qOGP
+AJwNVY1qCa8LKvK53J78MkaMbQ8QbFd/opQn135tKJa4o8ViQcGNjp1CCU/TM/O
RXnKmKuET8pDDMKFGRN/j4Wb3IXm7L+xwFfXAd6ZmyCIx7yPXymId0ljojzqCVtd
+kEDuItrk5EaNGzsHiagDEz6RO164BvnHT8WGCxyvALdT7nA/ImWKBkCy0Ac+NJk
9DTrswPxvqrdzUdsZNMlUrGCDjV8/D8NsC2BPrY2YCoOeUWkJWPfN5q6m203+DcA
GKWaEocQjSfi2//r0fW+seOF7SQ+9mS6jKW5+NPKwT8ldTM1igekLJyUWyV+8zrj
K43sfDqyBooRkaPc7w+uvJ7jFT7bLKMGt8Am4D1cNJyERf9DSKIkqtKeuSYckRKQ
6958rTxCtssuTAmC4uMdkb+/iClwAEPVRFmaJYSCzKdkVlJZbnT8dJk/v4GMGu8x
DuInxuj2aKHbM8s32aNToQIaxOrECg9yCJen+PZi14frhlN4GkzigtW01AQ8xTjv
H8nx0CsL6KU2jeZOcYQ3AMLU3xN+X8hejVkM5W/0X0ccRCnvks05arrXQp0EMtIm
OR1cqnyf8lFV0XsYWtvaCnKPJCElO1qqG7+RAZhj7xrUFqKB/208IRMiAdNb7Xv8
ITl9U8WnHYIMGRtQSARCA9l+Uo8Dep+7TEWsIvNrI9yZTE4Sjj1r1YFGht7kmANp
eqqviioocJ3pYI4sAyDzfOgVPlNm7x3rC1CM7dvUL+UFoYzfMg23OTwSlnDZkXLu
D0Ro+nQNkfDZlo4sbJlqx+FVe6C5psJaVDSbmoS9NxqKusJY7s9/2tuQVgS5p7uU
Ex+yB6ZIKiwmVj711Ev56Z2bik9DCW4JFdWk4irOHvn+XCt1YkCIVu45T2mbwpy0
2/pXQiammWMpIwyZ8uHUrlNd4LMIONbJQ0kunT+eLeNSoeooopxAU1wBiNDyPGxl
Q9dMXi2T2LXo9DZVf/LhzVwVTC1tMbd2ABvX6z0Mh90EWdmI6A4sT0OjM1d1TBbl
uZ47vHVUS1h8ulKOr7TwLzR7MG5lP3lO1uwMN6TJomcH1hDoTsaUrYxw5yjhBP4w
OTeSeVr8EzDjU4gksN9d+uqKqzMw+9l78+CCnKZ724aE8IScNYHXFNkNDcZmpab7
PzdXYx2jnhTGoj7U1QpMU/2rSKHMN5fKbVvmGHFQBgcm++lLoEolk/3HcAsDmsaG
vbdOhOtrpnVn3E1tPuhoO2aQ18kyqUzGqbjN1asLk19l6ZqduI14/e6wQGFJ+yQJ
rA7Z+us5cAvwA86u9IEOKl+IxZLSnD5emlOii2zoFZ3ti1L4Y9wL/NCqTnrp0dks
7R+GMAIH5x5WTlScKZMrMsXpEAJavhLl7HPhXO+crHocrxpru5tx6OXE9N2peMwm
x7zBxwMXdx9kxefUs6mqugDXvMwfkxG1GuiE72Ag4ccg4AwzhH8IbSPN4Qsqka5+
boNcA0fhlMcoq69VInO0uqBC15pPVa6lwUgQPrdBM8rBFXy1bQ5eDy/yKv0mQdGV
EmaWp6BO6ZKnZv5gPXN3J6weW59SLIPDb9L/JT653zGLnaggbUsvFvJipsvXtIW5
USp6nkC7rYBQACRdjBKszCoCXzVusmvKoWaSguKOQhygJkwZmlU8spkYA4UmaxJK
3WQmCZR51aVzli4wOpbFXB9ALBIKLjVZGvgsL1YA3LUxa3lqDnLjB60ouzhoDF0P
IoCJst7zxasLwQDZML3+UivwPuiXrnHmZLExnNPiZRrNYIvnJCZy+eZu1XdF/izW
Sy9HATf5SdfhKVxfS5Qzed/WMza8uX00sw9Rq3FhuFNy9Xmq9NaeCGFYXxOS0Flz
ryL1z0+/9Ani0evJ+fYlOzhJFZ6Gh7RhUqcNet1jMkaqYz/vqHmlBOHXyrjbkeVr
24iZYxumMBikk1K/yOy3jotWXHQJWa7Wyu9typ+cCy5Rntom3eWLoo9m0vkMfE4D
ndqpPoXeXPUXXrPtRdJCeIt6tXK2jrK9CNPR4gZLAKhxT6DKeaSOhqmj6DxP3ksH
QMubnZ0vGId9IXvn2zcSueNSX0/1XUYjyJs6mYV2WxNn7oCHSurx/PqssUuMDJbp
3hpr4Yo0QFel5gVP9ioFHIFyMt0q5MbIp2Ahpc5fULhhMswayL/EtOZ9t3tIbDiY
EHwnNXa+w2ubJztwaYDe3jTa/MYClM/uftrK0aoVuIlr52gl+3mIrT2LSiLOdSfJ
8vmsdPCDn4uCwLEdXNpQ6vysi2GiXxDCtFvQnwvUVDEeywvPSMghORI51gXh4vhC
+hPgZ7r4ugvjnU9h/d6zjd2ELnJRWEtoIk8esW2VXiT5eh9R31IZm/GjbFS2gZwF
7s1iJBcsGGZhwIu80ji+A6VKycYZA9JyXruucM4q8ugJwhfVX6hXaHHTbziZSMs0
1rOtDoxvc7azKfFToQwhz17vNM9u4ib5InqXVdHqgE/K/lbImWLEnJL9cF47wPlA
CoIAjyDj0DUKAneWEOcDeH2gDt66jPef8T3gSFl4Z/M1rbAtJE3BVzhc4xnNHSIy
pvHfG4BZNQUWWwfnPphTjzkPALP+RMIgqJmCQiNahZQXnAbT18mG7TvjdZudNt+6
gGzD2Hrsj5+SRIS84q3epk9SZCwJIdg3KpLdt9tLI11ApYFfYWu7vWRmc+YGqlmp
iTExOlyY/iiR5jqKnBFGf85smkO0XHYUrpw3ZQAyMw0yH+bXq81HILCpEkuHSfp+
WPWyE00MVRlMgoOR2bFLOgY4s9Wn2S3Seiu5ihOlxyuTQGshVuARp34BUsarZDae
aHfWRVg5j1U3s1yS2z9KW351miFv1yrRigqW95nkFeY4hr1d3tVzwOVKSv/ZFArV
mphfh8QfFefZU8/18rurah6IXvP3rGPemQM8L6OE8DjpGsmSmWZtMTegTHSuIXLC
XlppQlUb4DcR46TUrlFN7zEm3wR1jLBbNvDP2IvmDTUumLIlUMbHFMF8JkdnGmm7
8DO03zEkb7WiE/7h6XbClSa8vKbB3R3bYn+WtCyBGKmSMe1jEPrfydcsTwC5/kOc
sNg3XmUQpA+SYYhpNIvW8I8s99d7+ZERCy/RRZQI5vAIZIjG+DHLcQs8OF1y7VF0
ioKqYiYmKsqYdw6orFING0Du2BZfchz4OtK28fuJlku7HlIKYS5wPD9n5zKFPuXj
XbNpcmZAaMJ/zcMTabJZyXHTe4mywX9zB9sdookKsTskJxwNsbyc8FAwLNDNCRJ5
1M1c5VRcBEhWmqRTh77eV5gRXu2d6Cc6+HHlObaA2a+xpv5lRBiVtYuPfUTWfyJO
Tza9dsidAOxdGFKSY3X60aCYmvtr2gx21cfI4wMXFPUGy53NN0O6aEwjM2shzbdA
hCUlXfiLnV2vW1mDF3hgn2U+1V0bjNdrAwnb/9cSZm3GecPWRhDNG1hXVvVcxJA7
9IpdozkpiqaPfWgsPaiwqVCpX2nyPgLdTZ8/6XwIZPzX+24/b5aBWB0AQmDpF2Uq
TRKIzdwfpIWebq45WygWMQlm+l3twh+NJzsU3v3fDU1L8rNZ+zJNM9GiSbKEqA8v
/zuxp36xzGvF4aSf8jCZPK1ZDGox/2cMDKWqIAYo5S8gkK+PsHcfzCHo6hFEANQO
vLw1HdP1yJ47wuTvFkd9em8MdErXDOvuDg3s/5xca5diINRcc+EAp6vgUpZIDXHP
8xpX6Qyvamb44/Y59p5j52gwizu/QttVZb/0aXCKtxdPlI4umZom2NsX2Zp9ik/X
EkSGhUOM6aaC2kecryjF+0UEh1P6Qj8tEevzo1vjHpDpGEc3dFFnlOj/dwuVOZeD
xKmcuLg4xBNB+ZZTvUBZqF/r8J3UGVS9nfbtUKQnkhQmfhgePNDtQga3QBx+qqzN
Cy0guPBgpjQwiFHSuf4PJ9rsQJsfZVgHHuVqjHLSW4lgkcMzPGqxOg18NKo+/kW6
eXY8lDnwEs0urs3xORne2A7ZZ8+GZ4YVqLvHU9Pfc1cu5zPeuA+AGYm9brSh0qB/
lJq9VfLzOuPHRuDoCVgrhTY2bFHr4OH5QOYMiwy32aMwLos3EEPgtvOFbAUKy3dX
q7Wmq51KjdzQtvuASsOngnuHiLxri3/DoYAHPVo7WxbqFvhkRh73R4hWkv3MPFoc
HiWIG3Ep2KNw4rokwJy9ANXPMJCtHq7hR2xEF2YkVNv4QiTwz6wzbcgU3gixBVzS
6E6JGxJyZuDczu2dZ+FMvSCe8mxNflLPgrkFM2qyPY5+0ihwUHEvYn+Byg4Q7Ywp
N1H7nAzkcUMhl+vvJCollv7Dvrr+A1LzOsMpAy1P8Jzg2mxSPG19Rwm3DbVg1mX6
1xk3cxLdvNnWGp2MDsjLvAEViSVa84YqxbJLp8nYb5EzzHyhFLC1wzmu/GNG5Vfw
iPIqaDkm51GY9o8trlE1QsczpIQoKFnsk1HPDkpVzmVuUUSTVrfKw6tzRupY3nq3
uFrLfNNTSO1E+JayF0YroB08HxRm+ETnPCxL12WQyXFq/MiS9tD8hNUpp9DGQeXA
G8szAKEH3bF/+na6SQFmOA71NCvXWNBCiaKJ5QXWf0TZ243UqPpuObl9g7q1XvB3
pOFGn07IIXc9yRyGLEG/dtc3tvGHbugp2SS5SVvYYPvV+pxb12Qxk2sVRyNJUoNF
PcDX1YGTsZdzdv69f2WDgQ1era5byBnphPKvEM3gyWD4J7JC1W7IMXbxvIJjcLpD
hF0ntU2sVCB7gItO8h3o3R5KRHgy4qvIhBDyDA6xbIz1UuhIiSQd2DX4iqDVVsL3
xAJkXXFPsCeiveFBhf5xZpe/hNKZklc4DzfIbT0qqgjD91DNeHO9YJaAl/XkYhhj
9KVQyXGAZxJRAODKLdg+7i9VkGb9PzRuCwu+GB4chiPq6rIjCthGyTa+5IZ8fil6
TlEn2hlQWbyqBLOuAGiaAqc7HWaynut7dmK6gMZHZ3PdF6b806aJB4xCsYZvXLKb
9fasoLFSchpTbsfTR2LUvPkbXbPFx/FIcsAKsyvqAhz6icoZPkGVU4gasWt2U+XQ
Edp7C8M4GGAUKjMIg/b7woA2iy3nCXrslbZFTriAoCFL4fy7wvwPFuET2mxksR4J
pxc/Y8llsmAJcPcT2KX5ldJF8AdzlTLR7EB0jdFhc3ufswgMETcdBzJ9m3674eOF
TcQGKOT0TQsVvc+MfuYadGHfvAXEscoSPOOgsoRF2j4yQ0klgHzmxtes2xmu1lXw
TbURsUyV3d6m8/NdhtuPm246cuuFyN3EqXWjr3NGRtwK+79azhmovQ5gpDKyTqjd
zHSS7ePSWG1ckMrtOafNU1Vj+LIxFvWbVwPiO6o4vAI60n+DUQdjLzjkKzoqqXqQ
tVlKWN9+DW5hqegazIaUqxVQtJ0hKZdyEJf78NGOd0gh3JYR54LTWw9tEDzIKUPw
BVDm8Mtfgm7lVBoQvLZEuicxKBbzslFU3YM50Hz/4gfhL54Jo9QcHzy+KDKLfh9o
qFzMGePfEqMFIPaUos6uTqnfktVx0zF/0gzC3rgdwbCDHlFKWsjKbnyq7yi/Bii4
gHM4McDTkhJY/9yxaS6K2C2kW4v+fJM+0FnFxS+VoI7q4d7wy1FWzO8fF/jLEiLQ
ZnHtfbJFk6vEiReRbhhEyF5/dV63o2JtaVoNWgHkLileJHNk+502YC9Kf7UbD5aL
5Hn/zj1F/s0GktwYHHfzN2zlPlAZ5OiIhha719tAFXFzxaY3TUENtuT7ISubrpMg
THrq57XVHChFj6jMY8M+9VM0vT9tZqe01SiF1zY0NzNQaGlabBsv+rdB/rurxKM4
8TZNnidzWq9oHusysEBR0bpIQKbQcJx7HUl4uzeBC+VTvS82J9MlmMVx1/ubtke/
I3vkhXIwTr1MMy/9Oh+/mzajUn/j5IxlTqzKswJHaTtigxjW3Z8rahr6XRM7yoNb
Di8XMjdZpqA42pxUVOalwvhZx6i2tpNsl+rL5aWKnUoZQXd6BwzD3ldtlABeW0qd
/w4ZSkjCKa7TuypynnZ/E+td+jwaDHPYQz+ulY7jlUPwpd6AjhzhevuJW+SZgXwD
SwHifnzt/XdbqEk2eaSf7x08RgQ1PldwUg4guLdvfl2lCEcjeJgJ/mjsgwzZxBGk
fQ4gDC92AmfHtiDcQE/z+tqv/MZvu2fE5b5kKJ1AtKnyQrNo4gROcwxLENMstzLR
PebTFTMgFuYE/duc1F+OXKfexSeEhYVt+q9fSQak6wQF4cEbkosxWJ/V+OTR/rRa
FgeVYNj4ayPuIJN1ngqP7438Lsrp6baRTAao8g95Xy4Z7Sy8nbezCr8Ak1Rab6Fw
G4/ZWbQP9ykXElh1GQ4l/upHjswTDIRxFLNMQEaL/eRZelNLzY2WuUgYPLE6+7qK
IrjMFZ8mBylVR8ACNgQHvOuxdP75wLSqkU07U9OtI8G/09xo/sgONR8aU1JeALEx
qY3BNnGugKOwu92+OlFTlJBNscvotkaD2EjuvX51pKBuy1EU04LjiynD9Af7dI8T
Q3y6NN2se/QY9chnxUl93a2KHv3YYWu2Rv91mocfMhOUVRBoSdskzuUhgjvgGxXr
Kq8KG+AimK50yz4PF4EZ8RhwE9GdpLAg782z4bB599kyKZsaN9y7FMKV1znLzGhD
LoScbo89G1z/h2TNftlQvBurtlrwR9Z7DQ6WD+cuUKjNsNxUVLGW9C060K23sggE
noQnJEpN3CBpljjtknkz53AcRzatLvcbNlYywaTRMfU3HcQXf45QH01wN5jIUQEG
qkpjTu1LMlIl7HVq6tkHPsdolBbw+44btbM7qSnsSyn9g9B+Jq9Q9ht/l75KMt3o
sffKjg72Peymm6bPX+oyp9abXqF6uM3zIqqc6nfOkxDxjAfDMnGWHa6iRY0Ghjx4
5sf8jfAs+YG2iqp5UOt4LKQyHyOf6zTslcdTKx1yZj4xjb4OW1Su5uVmHCrkkOx9
M9X3BWlygm0ejtJfWbwTSY/d/9g+Sze0mOCs58ZJK3t7wCPeeXSiI9DxICJn/cNU
ntZ1A6rdQgT+LTB4RPpR9gJFnT8r7vNLsk2dM4XRhX/OUHjz8uwMxBtEWvesjasH
yAKuzNdP0WzhAl6g+JSJ5prYlkmmFsR/Q2M1xQILPkpBL94DHe1bwPKtc+0/E338
wY5a4g/Z6Fn0n8FtWoU3wXZj5hTF61Rl+Tzi6Y5npKFIzj5ikFcwVxu0GtRwIuO6
AR5TiDGYAM9tfVI4e66sx39aEQZgbk/wZt22xMtmPgtgvaW4Yasnljp2M6fs1Ff2
Mr4YQYBoXNYpp3XRYGUrFwrS53U+KZHTWmA/oY2J9I5oHs3WbfCKTjYrR05yT9tl
h0KSsJ8LEhGBjTtWFy6TCacoQPE5pmduG+DTrl3F6feTSVccttamlMu0Hme+SJ9u
MDUmo5CRZT6dc6Fpf4HqxRxctFlrYwxSU2kSwKmIU4o8377xsZparLOBtejkGAgC
fJZAQ9Q0BghUsBvzqxb40D3iGq0KK5KxJ0HkiFPetORbOyHai8vkLYXrMj4Qa80x
4tRI0eaYtDzA38dFeO6qENS/lcStAnLrqS8irXV1DcrP5yNXJmXyGX3plnSt1p7x
ChYgDg6mOCtWmDQ+o5STCqBNPfkQ5qPUKUDpvtHr0PmB0mBqnqXvSldCtq0SDIXi
CNkmfZ2sCFb/L5eFQtygEErBTXTI+DItDo0RJKl8feQB2tQC+aUl2dZG5vx71NqI
4p4w14rKXWRoY6pzA316am7C9bVy9n05oGtmzkSh6qN8YipITSm//dVy/K4F+uue
diWRPxPCJ/ZKsmFaVj43bUcykx64cZQKC+VHQsnwTwtiRUOJwilspr3RgkoeqMQ3
jAk37nkTbRm2ZsWLOSZM1huObGEwkxbHl+SQ9+VnAkzA4brPQcrLCkXC1PQokHHP
5ksCcfUwP/vWmuZ1YFfKfaYgM8duXoVKNItExkRgFnKD8MErqQqRgBnFwCFclqtD
tyklknFzbbCyHPAP2p18WMH6dun14LDe5avjBmumia3y9Pwp48Of9PL2rvJZXFXH
wG/w4g0v9sxuysHc28Ojjy+3RnZrmMs/Msr7kh+Edmjhc6D3Vvvqil/BrS68SOTg
0AasmZx+qNyKEccGyCTITlG4cvAIMOXWGyROX3dL+HFiP99qjwWGlzp9oidIhgsp
0RfiRxBcO8ziz6s9RZXTAeI+tHj7pI9k6lRSZmjNmodsl6fuIAFmkk5O2u5oxR/3
2Xhqq2zD/z9DUo03LyziZKonJbGjiJaVzxcFgd9ZYvE60JJRYgYgTFeGlpRt2rNj
O1loA9ealwvpaphSlWe/p4TlnaqdDzxPUMXuaytOKuw72ZFf+8JZC2Kp7C89rPL5
c/QjVcEDGqkBa4z2aP2GPp+DefqqJ/l5MAYDKv+dUd4YjYOaYwbZlPDqRRdPo4U7
KHu/tpyCvWibDl/J0abCk0NRaImqGCjW1U2jjJ6Pxep3MjNy0PjUUwahLjc4hIDi
Zifn43gREBCZ3kCFq7X+38skw3jIK/XMqWg9slF76JilcpwmTUatwTKUH2hDSNs8
QJGjwo6T+1AK+T41E8ltNevkUeVaQGEvVATlZuk6lvGJbXASdMIDd0b0MlszrsyY
eSvtRVSoW9Bm4RRS0t+UAuODa8+AxR3eVAK/SqWo65iW6NBclNEaR4zjvhLBKiiB
pYyucwbCOLnZG7amsDdBnmC3fBoH40b1pbhJIXJPjqVT9YwD4lVHoAnzyn2/gTQH
RNVzYiREm1SjwP8tfKlB02CLWjtLyA7cLJcsg2Udvnf6WUcyINxROoNt6BBkIWAt
kVPXHjPmejaOTo+cMfhwOxlQ28+mUp1qv7CtXAv9cv8CLSx2uyFPSWKNOUm3GsG7
wRkgHcVJP74srL0Vs1PUBWpnEeMv4zP+ey5xzy7wfc/Fd9hOUwONbsZEc6YnW89X
uVpiX4xDlPEYmrQeAE7Wikhw4Aqc9vm0ESmpAQNojKjUWBeCnqr28X5m1y2JYY/M
+BV4rCNKC29OzWz9RAe8m1rNwM+16Hv8KcBt6nS2wVemFlQIgdB7m7+Ol47cDuV3
IXvZu6helvk0tS3MowSppNQsC5hr/v+AR2LcPIlPuFTOTPaWgZHzbWxCLMe6X587
7OpQ8ea1A45laDvinjWO85D9mqdTNUiwo8agXbXrZp4YHz4VKfeQM2swAS7jObRI
ZJC/itTqDwm2NIbOfnotBcWvdWjTgRzdpn/JX8c8Q2ft8ktYPIk9jkC02gUQ7Ae/
TMr7PcZx/iBoG/1bCxApKumMjiJ9pIftmTlBmS1eL42c9lEscsNw4zOaA5OIDjHL
r2tKkuuv+SkSgR7cBk0jWNYlIsTY7AoaPgYtWDl21K5cROSLq3JSMPcSCHueE2HW
lX8j6XbVNRwKH2rb5etruexO0bVkkMFewE7ZWAwpFcP4U7Pgv1A2aBGTZcuMw1XU
VHAFKtEa0Fe8EELKrTcrcxPMF0ImXPqWua76QQXevqVwZAEumpsnq/RRBCILbo4s
fYX+2tJ3ysD9eV7T/wG3WLHTxr/TpSfoXwMX1lzSf5XaqQqo0ojw8rGDxq6LXBhP
iFBMN//0vutiTxPh8tadJYXtl2eC/Oph/Clet9Bqguc01ZkjHo+DZ0sf03MKsgTJ
+8P5zb9FVKzqKd7E7ZWFesacx7/yDHSXSRW5mkMLb5I0K4u1IVk4eglehdLojuLx
fc0NJQBqUhvsk9p0LKdXsO2YGZvD2W8HC4vmH4u8OCfi7hUri+qZ3lJ62MLFV+mY
mBP+0KGNTzmcU/meHQ4+nnL8rlMU9X/prXQR/MPQBDKtCkP+msMQDeyxlL/OjAKD
eWePtUfjouRSfE+W1gm/zOPEQIb5LDSWXp2A2y567FoyK5KOWC0yCw4ytVfF7v9w
sp3lY7FawAuIPIurJ6YVExn/lyejwO2Ebos3ERl+ZuOoxN1Ysy7EQK5WXqF0uep4
0VJHNYeQoAvDUDyCtjfU6fwqw/FIiwZGaXkQmB5NXAqVrovWjKeTllRmsCdmqJ+c
1v+CpXRnBhmFJQhbrQcfMqv9axxlEzc/bwkoPQlLWBUXCW918xGEAfblucRx6s04
ygRhVcVyM61YEa1gpTpNaK+/XcehFM3YZ1wfNYl52olbaEtWS7FYL8dct7vwGcM5
zo+9Qvox8KMoL5XyMOouHoq9dDfTs74E3+cbaeTDzZnkAkGNI7haIoSD/yQGxtfz
+kXS5ZLcJscUjmSz7TkidRGO4NpOiy539cuhJBPTGl1iwUwIhiLnnTA49jQdUHBF
5D3T4ndc7kXotY5aJiJIaiDduSSqv/BHJjTpOggAPu4nhYsB49obNhuQXcpUsqt3
giHtSjkpeMiqmCoAkj3odWNprgls4ty1hIIf/3UxPeN/hxsgSUZcl78qBbx6Z207
BWXzodZSf0pz0APe2oFxC/ckW5NtRLZJSeFSyWeYd8R8YZfAqKVl0civ6hfEM846
07/ejTGoznrqQ3T82hW6LJQw1wopBe7MIWIC9/fQql29dBtZv7bcJZENOw35Tj/S
rIbGkupPiXNBpnbnzCocPZxGvZgrBhzp5+Ly9J+00C9VRr5PUoqzr5qLqpicyRz+
jWaPOGXdnmOOpoa8a/JRLGMSO5vHnavKOp8JchESpVoAbuDXPtANWGJqu1cD76ca
2GRnlS1/K6liY7VWsCQHtxW0tkjT0ZnvrpV83huJYP6glm+AYNqEFgnykrtgKNBG
rU1CLQSJK6mblawAVv+NoWfeKKIeeFssWaKvVmIpyVN+LtLg5/3bZQQmo0b9rjU0
DAwqig8KGI0s5B3BP4KJelhJ2bEa8G9thELhISD2Smz9/bIzw8pABkYjedyqUVgK
xMw7cpiBz0VMdIpVLgrmFyVaDINLNep4/YStjR6e9gNhGpyNWdQT79SW0Od/klxI
rGqUmgx4vjK6eq8B0jPrG8L8kiNm/MCIad65bxHW/Lz003lTDk8+kztB0TfyZ45u
+ajLOmm9YJFvot3s0EaAo6kAzKy+MOm7ShojoXqQBunn+wTGTWZZg/GhgCOEMY78
osBHloVoUTvcNFdXP62Uz3uFMleNQPWdsGAfN3mlch4VxaDPFDfOUFQczFm/SKPI
Lo9FO06x/hi6XuvWBXEgZy5aGFCyo6DGgPG4RSq0GOrFZ8KQh3QWhhGr4DAcwnoh
sii5GFg1D1bNQ/ye8o+Gak5Hn6pqm0wKQPAg+4Tooq84R2piKZOmyZ/+3hX0XN4o
UbXmueHy7zCzMQhGEkjpT1XW5MBdpFVnjdWztmLz3KAZy4lAu391UJISOVbLXfeq
xw/B3WLB2y2sUUJGcjV3PnZEarjfO7e91yYThmlba6tCslh03A6dxvo3ZpjAtciR
NX6Oa13WWgJOcAeCb6F6dDy58DAPheUYmoChhxM9mTpRvVMVVzydwNMsZEVV34Wv
jEXUe9sz7ZuhlqLovRjRi25T0u7DrjT5/Y1HSVQfBDioVSHP/WUNCpQl2Hiy4Ve3
XWnryjhIbEIAqb8ybQfRVO3jgNaVnL3N5RbYOwEIW+OX3MU9dBItmP+oeelMi6yx
ZpQ3B+I7BKeJ0zja4BalJNhuug5CIbhyob/vakwEOgnCOZQGoTpC4N+kp+rGL5uJ
XaK7jYMZDG5KmA8XSvlZNdJUcRJP3sqWcepPXjdbMwRpsMX9wMjv/bm+4PQ36NTj
wy8G4NskiDJ99kH3R4lI/Q23fJhmhUBAD30br31bYjknWoUM7PdefizsYMaLNuw7
gjZ60LzbGjcRNavEA1U3TplS2F6VfjHLztyeNtTI4EPoc/8NoL9wN/JrH6+85r2r
XxoxYMrS3Do0DnSrYyPgnBZVpXtV+1nQU6/VKBoCrcOCzx++4GdAo16ledsGIXAz
amf1613UQfC5OzpF7QthhZgVOjKEyGyepEGN2TdmGjxMoZUQ65ItesbmOX702WCR
ZHH4X5vrNM3PlJsD0OTSPBPm4uTKkZuegq+WV1FxKWCjzjwJImi2uobaraxHgegA
R7WB8cGRo8PAZQzYvb6HfjkadLk3+Oj9lshP5E5y/1nLU6lQeafik5JTIe7oKtzh
pWhmeFNlMgsHkEB7m5F2L+54F9sPXcIQgHK4+jX1qAWbOmvtGvz8W/1E9IFzbwM3
LSOj+0ObtuCmRQ6Qfly5AFlwcpLlmtbaGVYee/AcRpgyUF8InaTSE6l5kroOpJ1K
c/n9GCi7X1FIRfIs9TRi12Qo6HkxQ+jU7zPc96ljY0CoMuTcdeaA1I6zmvf9u1Rg
17IjJfz/HY0wuO6dybV5NT5ObCNY9b0Ite3S7wRx83miggd/k5/yNtcKjOyVxYsm
FUnJfSPh5hdkRKxAPjr3TodY8hss4KnpZP8feJQqrG7AJZa3Y9k5XlGv5lF2mS1n
nAg1Ub0NqmkviST4nhdR92eW+L42P9bUxSlBQ3Tom3fiTEJ2i/w1TIGxRxtZ17Jq
ELELCNhheQD5P7Swqf1mE5QYqFVsjMcwbMdmcYY0OYdVvlBI52Q1c8rVuwHgtGxh
RK8V6gQOZsxVZggRfb17ArCcjEmezOY+T08UigiNMRiy6kMwEizJUmo3fXIya6Co
W2cFB1NS0MZc4TkNEWdjzDAaTo8t3ejsXuj2TGpxfWV3xx0V/t27/osihG77OQER
dQFSPeksecXL5XEgbg6nvB6ZpxqwVDYrXUnR/q/iHVUPAdvUbW5jZgo40wGyTEtM
m+eEYP4VA+ujplfZpQ0zdpxpiiOgp11rFG2AdbWeZMcWgKLunQ0XU61unlHgQHxe
QstfYxxGzoc0ObKFnIfzkpkyALztQnArzywyRGXf/cFE75pVwAu2UhWTUX5gSa6p
CLXI0Z+c8IphL/WBCkmCVVahOQN6k1s6iP5qfTMEcHHyoZVaDlhwbfs9QmHLmyOd
L92zzsT7JGx3oHshtZzAli1MU8E1/3s/NxTbxucJhGiLN0+NrUFye7GaUjfFYVev
BUjHh3Pzq3LwktA/tHwPxOq34n1inYfoSO4zeESvJwHwQ0ZEND2Qubk4SU9W2nsl
I4STxVN3rOrwX7w2SFZLQmvDCd4JTSq79Kx86LanAatPIHGd0ALT6gCRgiP4fOnu
GuJF49gIZuaJv48L4eEa7QEpXhytDjbVS4+V2QcmQwxto7uOvym85eDHV5Kjxgtq
e4yDUpd9xh8eE/QgNiHWIPjV/8nnIoKizl3dTynDX9das5RIWRQ9kdbrbH0f4JIR
/RV5Ov6xgq5IsV7MxyIeNkjVLWg8/Y/HdbND+2k85rRcxGuo7qxbcbMDQJTeOglH
2E8qV8Qw4AndxpAt4gmhSs2SimMfpPD5ir22y2aDQHOcfyd1b+qlpaMSOCuAFYzR
CUNz6TXCncL217ZHN83M/zwE1CXjbEo7mwoSt9fdyYTGwx2bwCIlpdEjPvQZwFo0
Fw6kSMI/bg4yIvX8OHfEufhrgTYgb7LgEzSPQoKuSRLCmOjwXEd/2/4gzPdMGNPm
oAu/afPv95zBHaF0mkPYeNEpQJ2YjjL/qkfpIgC5Z0In3tNRTqHZ6kmjQfksIang
yhR60b278JibmVQY/5ZLqu9fYBe/+u0hzyH8EFAhLa8bAx91nvy9Utgk2FAYb8/k
W93+UyypHbvoz2SGreIZmfiNP1Gizpf7tBzTTBDsCrqubteZ3DoUz4uvuD4w6j4q
I2ajYb4/380b80Tu3rB1GxKrHGKiYsJQYh50Nf0vZkb+QmDx5KZncS8hZsfq+RN8
uW43kHyxDQFAw/011fKgaaHUCzHj43mDA3fOVKhk49xJ9HtfinPsk0SQX9oJVrp2
cVyGfOvLCVU7hXi2ySflRIsilt7dw6fbLhXyExu8QijniBNeJlClKG/GwKzbT8e7
dxilreZbrBjQr2ic3bylQ2rCAzpIektm+l18qqa52ZIMok7l7SS87vGSB31qz20v
w2J0Gvaax/y8ZdoXCqgGeQUak+Dik01S5eRukNPTJ0gcoXmvqB0z3Tg5h+D8Ep8r
z7GaJKccAqMvf4K7UYQYF9XmH4iu3UFHpJ0aXKtnR6PLDeaAeev627rtTV+TaQBc
Bo1kX5JL1uSxpN573wZQvdBxG9oqq5JRaB0sGLTZ5zdnPWBsj8lC47aT4sjjn7rc
PUcoeamTgbjn9m4ir9kM6PpY9u7489zdSdU5S9VKXXYVszvrdwuPSCFgsAymrY1j
bOGKkXicBHf1yJxsdq7b0edrKe2hbR/sUnaeeVKgpSxZj7Ze/AYStOxYFTRi1YE0
vNofhCwj86ATN5uHH4nnauLDhJjhLbtJgE3S2tZ57b4TZpbxr2wnwFVIHuNLZTsJ
ZZO3nE3j2shAnirnOunAs3/0tP0g1ylCLQ3hlAQZLJf/TwTASZIoOa+kSH8WuGVi
mXWtoxl2cuM4ZO/n/UtQM16Ek+7T9B6N3rgQ1OWCMWB2wQl4+cwUIhwJfJmz51JH
VNrN3QMtIvzuxpM3ZDSDoQhZ1bm252o4Hs8I85lfbBx3i/j3aTZZd29ILJxOh3fN
uh7p+sQYh3ywvJa44ek7tAtvt2UJjNsgvKlzrySwHuiM9uqehqtJzG2WD1ZmwmmI
tQXMNg9W/7BosJOMv8E8DgsHPd7tY+qznp2BdLMR6Vtw2LsPs2czRxrt2JmbqKbh
7CjXZrXJ0fLY3VBkpO4uyPSA6riidIXSYGT3bwvs+/E9j+6M5rICxKYGnvTIpVf0
dhTiaD7nB7PXea7Oa9+5AWM0gCZkstjMQN7afGBK11ck98XzLpdi0S7cM12TyUpl
vaw+ghyudLegD/+dDIIdZ/hNmO/6DJHaoNLl9IvbkCrUfx6WYgsjrPm8/rIVHCkc
BCFEc5oYHyZH9uG1kj7lqlp3JsamvCc3pFqr7Dxta/gAzbiSb8np7IXRq8N4B8sv
DRTa02ifAMIWQAAtM+Wat4L36Zm/ABHHaYkCPsi04OPYyeEAcMTgqa4UYyjNI4Ku
k4tSbie2CV4yZ/FuG0oW+yB0bAuMapOH+fsY0Y6p1kA2V+aUywKlHaHiUheuNiCL
k4gqm6WqF264reBiFItrfMJY73nrkt6zsLJsgfH3tXTumOMXP+x/TyI4/x5kNQCp
BIpfn8u9CHdtpF1A9/JcqB+6rZqkmv6Lw/8nKJ9xOFGsLaEf3YtiIDX0dCW2FWAz
Vl9i5UXv0o+x8lmYsos7y23VU6ModNrbgNx7DaVxVXHYX2mMXDpeEdh7Ep30qnjR
eVSUCehI1F3ajDWlHfv7espRlSFcOkiV1l3DzkV35bYzzVfB2FMxXYweeCZOEA+l
8JKcMfeq+iaPgLHnkmiR2RvSDCH2ERu8IsZMW6iIgIB4OSKj8wWbj/7+JMqTpg8Y
BnyeRDCIkBCZWSEEr9M77fyI6XB7ba7qgduaNfiZe9jtZgTV8AWeCGWhhXja5pvQ
o8sMD12zHIUFO8hyJZ/HA054rgNsEWCi7b5TjvWX9aoi8wrn0D6rMMbQyFnKRtU1
b75MevlTu9jNcviDda8OEZsUw7GyRiAs3614EnH8mEuokMcbieeK9+k3Sxg6fAoC
Oi1gDqd3d3jQQ2vvUwjeZjg+pX/Pl6jk7LBv6JTn+uRdLT3NU+HYmiIbXnYLHMIc
/HZNcV2f1fOEItYoCA9Sd6VAZEoIewjbOAv5tCu/hXA7qQ0XL1NDidpgCuf4XiB1
pEdN4Y8fTDUl0QW/QIazt560uqcfwdsvmAWehOS4yt2Bcn00kHhQOKPcsOYrvo+E
Zj3dAjlMPaXgyY5qv5O3cR5k6oPqjCPIrO5NRN8B+02H29eez6A6ZRQgTxY4fYkO
7ZQVRlz7D4BxTSqPvIfNy9eqOacdY58dc1GLa9DVgl1YDO0BwNsN5dSrE9LEDMzl
sOm+cN8A0DX3cd/j1cBZ+Eq2PvA1oH0MmEe2Czfso63mbmVFK4hfidLcWOIEGQMg
9HfKAmsg93owcDOGmnjo93cWglQbz10R0oj9+4N8WBzJbS1+UsolWsz8quYxIRv2
lnjHTo06Xnjh68Y7qxtzMCrHKPpa5IIUUxr6kCkQh4yrBKXVZZOfQlPgRNuI6vvR
4GCWQYCFUpe8hyq11gDw+0nq2wjLjx4ug3owGKXZqCMpdL6WiGbL+pHn7KGR6eAi
C4wMYiy29Av9lf36CWOGZraNbq7dnFO9JC9bR0BR4FpvEvSUfDfMNmQhgPu5oFUU
O8he3EpblGxTKauGeCm2GnwcC2mnSYC6mDCNTEtny1DhyIsnVC8r9WzDvDZczS3t
pS61pEF5ucbRtoiyA1bdFAoZnzkvwww4GHFHdEdtaTYVD1TBLHRzolmneTjCSltA
c2NSoPb3BCq8nLlnTt4LhQWTfkRxSN1y96FIW5s55lx636GkjKsINBlcsZhNppiQ
ErWk6L+qQu0BaZjPW6F8zsC6IUO6fqStzZRgJYCkXqgfWEQW2n5oV/5PNnoYNbld
Jj6HAGPHvCJjl6gwMsAzcXiSg+BkH3ZsNscCdxZbMMg4yjqYcVUDqX247d+flJOn
xmuSWAm3V3BEqddpmmvtXF+htpoOWheaCN3WF8MLZVyjS0yPyeueaYpUESZJvWGe
9iWXMmOJ5TA1XIL/TzwFIQj9udnBoyVMDAXg9UqZhipFgt3divyGIjT3DVsfhCXc
oOo6CDoMh23r2anIFE3R4K2I13TvgXuIojBOzNrnx0SO1XtuQQJoQ6fgQoJJHkOC
fQGsjT/sbThcDx9fgTny4vzLXt24UDwPRw21R3oimGk3nMbUHsBw3gOYgez47OEt
oy+fNH1F+BfxZwzbbKy606yI/tn6BZgjX16doU3SxEzgpqzCxebMMIiFbKyS0+lu
cx2BXQfu0w5bskZ3GhabJamYoRdxqiONig9U29UUlNLLaJikUZDQKipDqY7vRnuy
Ih6fAjzCsWXIVUCumTWOJ33GyAub4ai/znXaVRx1PXFPA0rh98NmlaYV7HTwiH49
r73hdddiuZmK4+F2Y5M69vXlX7HUD+Nn8XH04Q8h9OWxercUjj6SRtX+5LewB50+
buvenm1OuikLciIBjtkAHBmDhmWHS+WNRD2uORkMl0wTNkNC8QWoOvsXGetUeLN8
/bvZz0Fyq03EImkxSeuyeR1NB6n8+DwK3DKoIh91YTDQZ8ZDd6jYbZbnz9AQLk2x
ZgqhonwSCm5IMeHVz0swswEhjR0ei341SDHA+5t8Qbx7ESts0FYRxDLemRZ5UGgR
qrstJVAqubjZYnLysAuEy97aw9o0Q16FOLsvvd0ZwxJ4ywbbRBAtCYgHld9bOPm4
a3n11/ipr3tdarVpluzAamqzwVNl+evQ+PRR9rgsAjRdJBxeMJdvhkTJ/389rL60
BAlnB7boD5rozKODi4MiNlRiEwxo8hrhGLH4zOBUwChSFXASdTkJ8ZXOXe3Cmwzz
jO0yljuGAWrFSrbhu1UjMb0h2I3JUHPToHigzNDWnhqCzxi1xRCTvQTYOMoX3/bY
FVYjqQ1/zejSF7dOJxVhjHJHgLm1Y3kxft2Ch7+Xq57HKob2KwwA+mHsY7K5Tbtr
xqIQbABT34k0mKbw75gI/7YxRE5mxMiL+ntr+Z1ICjvrUhitck1lgWoZF+qYxAJa
T7F7b303sTT/NVpsMwc6GY1IV+O6mJDFtoVhc+sPTbk3mAX0Id1mHgL7nVLgzJVn
6bsWnTFPLnrVPqwaqIt+d/rX9lQCYD3zlOCiQ4PCyaOA5DYhWqLe9cH65kI73XvR
tiqwjC7Vb2RNHkagJq63G3pZZ/fmFm4cqw/0Wf/LqkLZWbMeDBXa9tKQw/C7SFHm
H2NdLfKsNMOCu7TwhnDiQ7vv8qkSwbeHus0snC0pXhL+AMJ9XTex5/ydIEGKGxQ0
2tKNAOJibzoc/2BLgCGBEg/TGVnrOc2+OIKPkV3TVVJs9SwKEAMXkNDHiID8qFrH
1eXBP+/bnFCYLEjQjNdHcwHRQ5ON1fHor7kzG8YbGHYcaS9ELr5yMgIfUNTEfQJH
YYfGXTDo3ZXke470DmtZwnT67bECxZfZlEt+nbfJI/TUCn9W5JE5DT0R5eHLjeY+
3R39qsYh4WA5J6WUlHCW8qTvt5KsD8/UrApTz3hotQzhNtDHmFUNXVf/ncnocEpF
qifOnYPkhV4yn3vJx3bXQAjE2SScfz0jaiRuphbkCl/2Lgkgdr/pqB72b05dzFK+
DFzlBfhlEQB0X4xq4xb31CFpj3yXBCwFrkwUsOdnESHaWCnhFdz5UoSQBpZhVO6b
YssX6MsJ5zvjEShqGMyyZVVCL1ugmMATNOJ+RZ2D99kn1W0wULFCSQX/lTjMzYnV
YnyLH6pgH32uRWTiyMl7ZHSkpJLhyvkVD9fvOEb3anwXarZgqBsVgN7y5zouWCFU
5La/B4NwfcvOIW0VYKHEX3wAf7H0Dy+2SucvrbpPeUrD3WENN4YJ7JVVPmMZYf4z
5KM8U4JyxRmzYc38YXft9JlXelFa0gGr5VaeF4YXKlB0Sm8AB4l8SWVvmBEDfVMH
AC7szn+4aO2KpJ8nC2tg1vUG155LWiB4YlLyBuubeJo7av3/x2bj/+TKGvSfbUFS
41/Tvu6jcoyB4Z+KQgfBM4yaImTDqiBku8Q+AMug5I3pMjcCnReuDlG3TAPVOIls
yUBA2fS0EmDoUPHW3LFFL5/r6CmVnJqytjkzB8kxEub8ns8mErZH1gidO8Oe8aHz
KLnLpjAIxatAYJBWw8eamASIDbS9muDmpymfBcZyakw2WdJycoHuuc+l4hBg1ZKI
Ehk8qaFiTVA/C8vptnmy+oXqYfClDvhP1GJaXHu0zsaolJ54iYUhD24gVWdsmiJT
49bt78PjvK9ARRrmkkB+ofhqWCXtXFQZYVHcO8BOSj5WNF3e1SpyD7MmcsIBXaVU
9bQbwOK2Mbc1IGfQPZwSSZ4SyBIVN+erIgFu/XxkvJFxTd20xmWOqLsn4eru0STg
vfWhYYjMGm9ml03KcyD7f0mEBWztPXomktNhGqwDkjpPNR7F/gzE3NfuYi2qAqy5
M5m46LnFrn2i9j1K1s2DmMceNEk5zif+env9OKDxsp24+Vb9x2VgO1EqZ+0yhmTY
uupeOs1BLjV4SqS4TGFsSmRYbS0ON9eDTjrLtCWD1bqca7arZabyXR+sKQiOmjy/
Q5O6p4rXEBJQFMP3qSeqoLLNr/bMiJeG6eHHmr5UR1T6KtWQ5FEfCxbUe5OTg9b/
VaIukecdMjj/pzt5w5AtRgwLr/oh5nbMrNaqTRb+0CasfIzPWkQA68vfnF5yWHBe
IRB0wd4TYPdj62JxjII4lwHn0YWXYFKmQrWsphiUkRiVf3QV4FTrtudwYqpRKb2K
y0hQpE3sTkSh53OzpFqtmKUxglJnaGlUKmjvEYSlKr4Bzu/cbucG3Dh1vE1CUpnw
5ocAs8dwcX0G3fHWVRtfpCZbiJMNFHdW0U7Gb3KDb0z7reH6FiIO8yedy5maY69N
1gHyVXwKtI6aMA1DKbakdco/VCAQ9xdPoCNJ4OgjymkGZRR9V6bPBX9+FL4kVOGz
RZFSnfV1HR9egq2bvDH0FlLrQLk672LS78/p5jlPcRqWkBpl2yl6u1Il5Ts8X6nf
WJQguHSKuC6bB8uWsnf5uXwkRiA/RXqbt015CLrZobSuV3HVVZ7cYL/TxR05DZPg
Co6GCB8jHm6aR30ILM+urUAGQPPt9i1/Z+x1hJl6ZAchixxplBEyZEJ5P/Y3WrnL
vVTg56ghxiFHDXSpO7hHdcZzRAVKIX7EV2tlFCL7Ks/eS7XucYwst8D8u4dxrGyi
YIfR70Sxunn93Yomz57sNc53ZnXC18lnMFW4mj/xMb05mTvYBtqS4Fls1lVy6a3q
HpAAaCmiPf/xm7zYYNjTclxjSeqMR6PzZIY9s330BH/xQT6OvIz7SfzFZn+arYV4
9RU05e38X9lkNxJalB/BZQPetScjdF1s7o9QM2D1mo9C8D4KlM05fgkOqsJeKHPW
5Rfo8HW/h3z0jKAGjconOBX5Nf+icCELCPbJKdLQPmiXLHxb1xpaLCx9j/JffnAU
SIMqVaD9ZsBm/5x8UqkzEPMnWXyNkOHV9DmHbM5SazPdjCWAbje5jCOd7S2/1et4
bFu+G0kdHAp4UMkdKLcAVt/dlEnMDppPr9jI63fZLNvj4knoRBojNePz/KEhN3m2
tXwsDYKZhIxGJ1OYAB2U15hUgvVK3I0Bp6c8YCkHz8dqLgjVcBtiWwQe2P09Cgod
6tPpqM4ohE0w24sQgQ+dflKGi13CZTAjfCiFBpV5UGURxXzvTWSkMWP6hgCIbXlG
WvITDjTZiZAvYrUk4tXaf0omNeKO3rnyT0p/slVdQR74qCpE5ffc9VvkVUDxGm92
Or1qP4H+1QiM8r0Iw6fPS9eSjis7Dn806xNtKMdeDWnsxAltlVLKrOQrK1qp3fm6
ZEG3HN1+w827YEgxHlQLcuGNTvLv6JDM4UXmWVzInBZL05oSuspGT+bVGfqRi7vX
X4Ip8qcg/o6w1H7bXV7260uiRDy0zlUQcRbdEFMz57yvOc5l7gYamvU0ngEazbOe
s80qa7WWHof5KDqwv7eEgkG1G2kNU3qbMXC8KN6SoSyqHSqXUznQ0k6GQyh46l8W
nBBi6ZG93uEufIgLkOGth+rb9HYYuVI0F9jHp+0fE9g33dRVqyD1D6OSrstxlrH4
72E3TbySAGod/kvIphjbNq2gcqf8W8Jk1vuOHL+OO/H8+ow2osoRRKdZEKDShLFz
S/BgV/TXhILu/wP+XZU7a+h4eLOn5HLuLlOkqBxRTigBlli7O7ntp30PRUYhXLuM
o9KSE+0omlA/B9F3jJM7f4PFs8Gr3qOtwwgK9EcL/IVc9Omt+CjocXRo8NHZVDr2
ZTja7/CKPXw64qrNcL3GHCVHa2RlmvqUj5NKOmwjVqfJdKtvkjx1PxFU4zjopjvD
qqCdqk23f6tbPKgZjmo7mE7dUdv6kGeQsp2FaO32T50m7Nr26eRlbEgjrlRJtVLX
l4tq/jQ4neY8rV/S5FJcrIchos9To1dQSOMv8VCpd8TcFtKacx0Lh+OozDlwgV/v
mGt9sZFFgHDDiBYxOrk39j6/jFSNiXH9A1ohC7MFUWpCq/2+2NhrURrFEFAM7sJS
0U4u+kHYF01rbdfIFRtRROVlV0/Ow6vThM7gGRvEV38SZBr3TaIUdT9LcuqOwjSK
JC66C/IobWm5KQE+B+4OFnVZz5ohXx0r1wRNf8AvHLtFwQzghJYNycNgRxmG4BqQ
NZJyeH1T/6q/UsQmsmp+JTBC8uBKiroYjyrKKwMybAXGbdDYESc7Hxu9Ca9ZWsgo
Qat0OBz2bP9Q9++yafQ5SEK9jIBAVy+73h/kMb9jRM757u/GsFNa/xLWLQmvgPhK
4ueRyteJp8NDKZgn+G4OCfBIzS7ogAnkeIR04fiahDBn2pzxod4IQqLMK/T4GqPK
WS3cvBI7Lb/mdVL5zqBfs4ll3SeenNKnQcwoD7PqgwqlQ/8ObJWa25UIne8pPUe1
F1n2Y3XG1XBKPctswWcNoi093Zn8/JVb/Ekqiipjy2VuPNVUPqV0sq9qt7xHuOEM
JlZAZyJuB9K1UY2Pi68HE5aiAhoEvJigznI0mA3UmsdeUwDfTDAWOyRWoIcaXhhc
dwQzYU51JYYYRqoZgy/pQtMwVXOOc7ls1tAFKxELXYSb7PUnZOTq41CFrcb7JG6Q
ZgLXF4R+qn/PyFV5lWuPI/gUz2FyJD+bO3Lrkrz4aaH0cBbUiF8wu1TozAlBk9IW
aC1ZtoLSQJEWPmrTi3j9Pj0WCtzxP2ARPoBg5ZKkH4WKJc3ctcyG/9ReJsQgSHTu
kHGti0EEP0DaSNHxqPFcVZMQJhqCfzYPqMFDZtEkNV5PDZVgKUC7Jj2AHaABteT+
SDMtRQkDu+iDjPB+ptDh2YRHq1YopTB3j/Tr3FdmSPuEJzxen3fNtuyWpLrOVKob
I53dkJyuwsxzZnYrG1cfmoiwab2OB+lSn9PNrpM8jrMzVmSJmKexgDTAlGSfoP3j
A5uhDvllVMo/HU0rMTWQTqwLTLZ3fv5olVI4VwoFHEBP+heNi1OtSy32kvjR9MPs
OS6bDg30x4MvPz4eJJ/nqSmg1ntLRFTcxDUqwGGxRKnCZVVmHBo+QhXcXtijpwW7
USt/7inwiaE1l7kIpxHRXBzI77HITNR3BtUYfuQibcCepEYgCWbDLIW2mQrNcWjr
/UuKiLJczM1F/mJKp5pdNs+KOa0OuDqPHczzF9Gd16FFj+vbUHVnpSJ9yL0qn9gK
nC/dnH+biao9oBVl307+NZFLQz1AWlPClExkmtK8bt+M2E8htRDV7LjqtB3oSusi
XnKd2JBtUildyTpvnUJb+vOgK8WpTDTE8Nteq6UpfhAZhetx02tzyrYuR6qnpp+z
hf5/ZFqT+/s13bI8nwcJP7CxLxBDuM/6GuPL65fTYJ4JF/fQwbIwIk1Qrw1fEtdU
ukOppi2nbk4GQLuwAl6E7fc55J6LceIR+Zm2kqTgRJoXnGWXmqaEwOaVVawxjTBY
MRXP5wOAKCHfkXcKpaQ2N3YMB3Imb6RddXL+bcOXfQhQxqVo13a0D8lxzjGiul4p
S4+lcTdaDm3S2fJck3uNlOgbHZ8nY1GMMf1yP3rJI9jf33TZAfhBqu0bZlqJbmAs
rxbgaaLLML9JS/z5c74dKn0PmNrn7GA8LFpnc1fXi83DPZhFyLijLtqoPAaFrRIk
YwWW5FgrpOKFOfJxd3G7/fjXkhe9CiHH8ExP7SW12dX3v9VAWq4Tq+P+m/K0SfhL
FJGuhCDHsyaxR2AWIzCfhnIw3l405XdDta1pQBSbhP+Z9h7XLzCgEDIlkbpB5Q9O
gaj7iowelFp3ZNV+iaDbpn5M5UI+YQ6o2TF+0eqb9xmYazgiVybFtS07upZu0gfY
esMz+Xt1R2mP7KUNdLPyGinexPzaq9tBKPOOBej5HMR8I3T3jce6sNK7l4W5XlgE
dkcUXZpPVFkScVSFDs+nJbYAV7hntlQKanor77JQrnFiBW+k1uD2N2WAFaXm9v+o
XSdW42//JJRixtYAZU8d1Zo4stGLBVEcnpngq+Y+nXT46DSFuY5oXb90BIfhXvRA
ylaswMNb0uFtmkztNrIjweEkGTHEamoJCKkVlcUWIxySbFLksr+FiHz1D0GIFykx
UKp0P7dvWucRfQ+t4PAJlhJMWotiajbC3ROoTfcIAs2BmSn56uUMPNqQdTsnjnSz
16iuRb0Yvfwm1FMpw0IKVw6RbU89Y6CbUsPqAwA3FJXMrLdJR0TuCFF1wlVBKZoA
DA9Xpnn1UWjNYYo8A9vpb3+WpIJZbvqzsLY23ucOrbjck8w+9rJVkSQ3xLbD0kB4
Fr/JNifoh9ZzEy1c019fhJV0YyFQ+VS2uYTrO5Ojo/L57izsRJ4PHzdmt5N/rLzY
VmuzQ1/btWRSiNXPzE2NyiPHDRb4pkbmBMpCOMJ6iYmsJx8rLhgwcrlVsY3+gtHR
p+AhoEsZ9qR37VSrpvP1O0UKXzP84XK1I7JXYXnRg3MVWDxTNzj+KtcLAubk/+bx
8Qf1qtAjz+4BNTsVnchkyIR/AGiUAXYYPDbZe4JYKuFUDQX1zffmuF6Rm3PckNf1
qJvfnfiif2ZKtc+zIgHbCdNsBpiSTHGxzufcExd9KO29Grsf83wDNM9saaK1kOfK
DZlk/0JJaRJYhdmbmcMPRUbVpP/0ivLZns8R+Y3k+t8bPpfQAccGMATFaQGmWdgU
rQgSJMRIJHgPof6nfe2ZRwWYi5kC5eIuglk8NbJDRR2Jz4QX5EuO5pmGqykqJPMJ
+EefWGb0tLnoCfPwtrt3KPcUEPdHrUW0nLc3zHjbW75zGFE5sDF8670RiEDksxOI
+vL1+f4pUXWxoMX4kSLpjX7LuSqTA++v5gcbOBdIQpod9rxUNIMxvq6l6lo/AnZb
5QYwX0chCvgQVtm2rLTLSGKnTgfql1BKy/YLFag/KXm0Q+YVahrl/sOQDTkSPIUM
P97M5dsvfJeH5m72vYQCxt3NAHQduXWATuQHyxwvJAFfO9ocg5rkGCzBHM4lKeXD
VrNolVYdqkIWVyF+Nr4taD+eNSsAjXSnNZ7/t8ssa1immIhsH6FGq4bKdmhO8DLr
fCNPd2EJUAevjc3bVZlKN9iYZVvilcNBgfpanfzktkFENOEGu8W3gBtwymVKk10u
s6i0mvAm4joihOPtkAYIhwTYwueobodGl+aCBFdSfZEI+INBJfXu7rpAQOdKY0cf
INK7JClwjrQIvTbOC0DnXmtbLghawpDlIDQuzE5nW6ySBcULirWWxYWSDhMXCSUL
X+g8WHd3HP88ibJAyrO406Lsy1WoVTvWl+o985W0X6qOVHoRpkbAaQ+Oyp4hRSa4
90r7T/aTBsiApeAjzN9NzKVOq+ODnpvjmDam2GMVuJ/iz/iod39/+p1XULRxOQ/R
cH9FteR40HdTAbmZmdffT7q0CS9T8+SpySwM/ucubM1uoaB7NmIV5eTHqxdWxjJ/
glhwrNmJh2bha3ZR2hNIvguGMT8ybViW6S9danL+pUc/wwNHAnILZtf9RcUFmbv1
xQpWvXFdt8SQdIgRqCKVjLC44EvH0uHwMWyTfUzt8/+rvLd/ff/Mm2xS7OVn/3gr
HRHgZcKhG0qmHDtKcQmbxqxgzrvGlP3OqfI9r+maXRT1o216lp/Gp3CIRiqnjaiC
96E0Vd6U8A0Ucuq0iCDkDy3LzG5F3m76jEU3JGBp8g5qPvyebmlJBVeAb60ubF7I
2CgDHlvdsWwOBwoHZ4pC8bAFFvOxLMABtJzVEdFSjLcN93s8bp29o9EOnwQMvtGm
u8O4+lgYFmPleAdoDBXvSqR0cE7WriFp9YAHjp8BAG4vfa4uCLBMSIyZbk1ZeIO6
zZgoa/8yAsim0fldGs+4PbY8K0KBfqABX2R/xJ2h1ObS7ZMwCjzvTScAqcvOiBgv
X6pxeEuicuFAs8/zTfCjwyRd/B4cpl6Ov3DCKRat5NSdPkqa1AeXG+qBHlVs8Cyj
KE7KoppAd1OArFLnTtRlI861xOOp0ahnZSY/QaBcHM6vYKs0nd4Dd6gm6D1rtqcE
bx6qK8mwOdrke/Is7jbuX5zCKjDiM7n9V8UB7Kef/dLxee6l937euuvSVQACrLTM
ns4GLqfhBMx9a1/yXt6z1BpwXm4v7gn5bmZrj+ruSjRXQdpsEi7G3dBJNiLtMJa3
2kmohSSeCfn7YHlAzAIOTXpRoVshyMocymCRft6xz37Cvwq/v//FuQNhc4fhgbY6
CyO4EzTquYKialoiD8CV12KFd+Hx2FYVwnAsj6+JJ6qd7ftEntD2Xfo6ELClETVv
JHuxaV+G/RsTBtREv9V/Le/SQqXkniTLXA2ROrMiDHtGxaSUrnGKuI1/ZsWT9IxR
6kxDLLVuqOdvigfOU0edpaIrTM51K4TvHr21R2pgPFvEWGnx5wbr88OqY5SJPYZs
cphHr+5CHK1j/NGqWXlkmbsi9d8LgjB15kH85ZjJsvrkiVKOPj8pD3eYtAOGYxM8
h6H6lQZVzav/XLRlj4kLsVvyWPFHLi+Nzpf+Y0yt7D1hS7fpkKb7hh/HlYG9E411
6jDgTyRSYXi2B6eQyJ4qIDZmwSDa07cZV7W/lQ/EQ2TiJS98yWK4jLK6soZLZatt
b1vcvuLoOkT+5AfAbqFfY40KoHN/bTaEvjF1DbSoJPirdcmK8nkt12ZMrpzrKP3I
e2VDYc0OfEtlosHUoVBgGu0ueGFmZXJCRYaeWUsmHX2IZgyTHnIUKR2EVm9AXd7f
Q+06FDkIedKiZpTVFTQd3JVHyj/ThrQesbDUQmbahWzKuhWemS4KEIaWBzghY5Nk
pdOScPyPU2mfBtNmLmk2BVAzSPIeO+MZC8WC4/E7X3NonsbCTCSVU0T3RRPeIxdu
dD+noxgtK7Vf1zXdWPEFP4zMkS0/WTbSPHaDR+WcYfNC9R8XYpKdysHHZc5wjeCm
yazxd3Ap/h59H4tAPxRog+etD8V94stx+YimoYzfxd0x2ghual45tkd5B9fttiyH
r8s5b8pxO40S9zkR/ihbVuBgbWiz75m3exmwmDaNJktChZe8T9WYj73m4bXGaiZN
OreGlYz1sV4B1dglpTh5AvhfYOE4ygoGuyQnRXwyEubdwewDJviqEmmrBU6ckwJy
IrFb1T1AfzUYGI5Nf9RCRcyXvE77Yj/kcOZAORJhVID5fJ9uDdBkGdQKV4CFfjY9
9daWDO44CcVTwV82T7tpD052q9fzNYbwHH17dEVpv3ecVucxE6Q7PcZUJl4peQM+
7EmoK+hJryt0kFXrr1NgWKYRSajfvjo3L0e92F8YNCtluqeQSh4YWH7efGzsD0Lf
K1jdvQ4pMYbU1tm98IzcLlafyLIviub+GJhiSdQLzYm62Ny0gUcx++GrtT1KVVFN
+Fzd8nb9qW7R7bxVeVt+dL1lWWrUtvI4PTjRuCTsbzftND3vITrFc8B1PvjIUlio
uSvm6cCs71b30kdCb5vZyjboDfagj/lmEl6TXYXtknpyT9AOcm0DRmeFcVEGAID1
rHrUDAhTGfMQMqzSTdt5Aa6ROJKqn5I882y80lPWImogtzYHiSPphYzzob+W2B+v
hOZ3lNCA/pLfifQtV3xzea1dUqlGqwp5fp/qISjDcWR0sqVK6p/lhCrTHOTC4H5U
NN0abYtxqBYh74I3HgMI4uPsiBa80OSUxpwXKcYcys2xp1NPEkA1dTnSGA9paHD/
+YVeG05D8pSYwJUzmzB2KAthkJ0xTJMzow6Tet+Q+PlPO020EXvB1O7uplCF12f7
7Ir32VFZroRHEX4ygnIzYKedbr45U8JUH8s7kxPCUSqaZGPFhUxWC7ISc+hC+mvJ
BXhfn1dU/PNXhEIX/YqW7eONiSjfXwsVKx38HAxlhSDQfh9ZiJXv58+tu23yE62X
sMBGSsd2ehmO5dMHprx/6wLp9n9/YwI2kn4ROH5p6b+Dpl12I2i3P6TZ34DKO+re
NV4ITMxhNqIs5wpEGDZcPw4VLE7JC0u42whnoVsmlgakuQDS/bIonY4kmCM2H1c/
7rZf+b7sc5Bx6cawMA5ucX1hV1OPjeNaFlBfhEMr2QIXQI4UK4t8j/0fN4m9ID6Q
MWbPlMLKCXBgsBvB3BrKHXEzZeAdgMzpEdcmwf1Dc+D4RM1tt41YL0wVs3Hyx9cG
H4u4Us/Dd7OSn5t0h1o1bKPWlimylzIWz0lhzpaGh1N75M6JFZrRrzDiczuLZ248
hhsoIjxqw8UIeum0eKd9/OTIbo5ZLhs0W54w453JDvdnwfBPB0ifwywDn02DoVCq
mCc1Y3eIHiSd2g3eSElOLKmz/6yZcujOPW5OiHk5ELRyJ72I9IIosEDEqIqW8zjW
5ghFTEB0ASK2j0xvoIOHlZQyWN8AXQ6agnXB4ZYKcrtK5cGLJXL9h+Kuz4jjWbez
VIHaH0QknKrbhMYWWrFf23hYFEKtyrJtt14oyenkRlRrp1z+osx+TFTQ3hAn4zfZ
AGBC5ZwGaQf7qs+lH8YXf/ebGDl6DFGDtXInbzSedy+PJcOxsGZl8SlxyroumeRn
ES/kMelDO5JhgtyJg9CAXdpA/yOH26Hh+5nbDJL9c92g+bL/E504To1BXDVPsk8S
vmkcB56g4c11194qJ+VyaGOKqkbuwPvzdEUJPjEbGRBD1BiypEXKptpV0BpJHdAR
2pblNC+9PK3M78vKAQ9+BA6LcBBe2UCTQz52SyJD69kbwQR4/4EuJd7GlFU+GDAY
ib1TsyWdhtO5PjMe0z5tZ4J3B9PEYaYHpa2GMNY938S0IxW/waFrcMl0fOh9duBp
xmT9Nxu3fxy57npD9kB2Y8d2m9bu4Go2q8WahG9Fvla8pDqUH9LCNbKO/4gabvN1
k49J5lLPkF5Lbd5/Nk+TJgM8rHK4eupNsob3/qvqiSBgFYCwRaoqMW1JYpFU1OhY
qn56AXwByhJcnxZ88G5qBqrJb0NC3A/74AxMYSwDWynoRHQUbvwBYcu8qzWhr9ZD
BWtmcHKNL7Xoqz4rZqVTDS400kDzBo5CwUPfYMQwmeN9PyHZvIO3Dz7AHCQCmwqZ
CAOysxiNgmxMbospkUPAI8kTMILgZnkDUVoipkXBzOjgSNCgORAUgOd7fllR5iko
6Q2w8dPLIAmrKpdRUAXjKwfHLAEI1DLxpP/yaVghTjP3W67HobawZjipQ6oh/fSa
ZksFX3thtpnjV2+sk8WqQAOOfTPjGhOCAy6Jkx81QFrEzE908iZUeMeKZpxcdSPH
HlPQKDRGpIHU8bhAeV5xDMK0Ku1Xjit9/awLowlntxkIPrJgA6xGne4JvCA07gEG
yN5bm2aky6FeOCCSZbY44US4jFvw+QAWEfg6hsGZSI1AdUQZKvTmjErhcaWMUEfK
jvU9txo2xTqUYQ9nbt7gpx0e2ksFoo0+EuHbbR6qo6oer7tJ3PLpOyJuABwqZ/vN
6/dkj/vBLWItA221FuZNqaeGSNsHcPb4cUrCkxpbuVmqAD/Sde8yzK4cTK1TEXJJ
Qu/1/2HiIa+n1wpxjbhbnZqK3opAGvAYVyDlwejLrCuD/8xFEWXAtSR17GCOhrrn
vChtGQ3di5Babija1E3OTZ/KK/3C7pUVUIsfzGyPnu3CbmMYRDEc+Q+Qo42vcJku
B0/8O2YLMAmVwqn4FTq6uV2PXV1ksPL/T87QEh0E56yuTBwGq7teAe6jBLDA9qo5
HZlciHz0xmbsG6Jj2mbjD84RwmQMoibJJAtONEMdfVl6F6hxc6TJIwyY31UBh+9k
ktgWwCGFTaVBGM+XVq+Aa9tZFy1HJJjanmTZR0OLlunQ6DG14Gr3D/84FdGYYa7k
e8FjarIwQrg78tP9zkRAIGDVFCGe4zAAvxkn63aWOYQdnpLUR9GtD8mHEQzgYBdy
3J/2JznxEDH88B1ZWCPpE9oD6Bd/JseP3oLr7nIF7uhp2l3qezJtQe8eEfKU1uCY
EKhZG0i4SRUt/IvU8wH/g9OElguyRRi4qbRU5rI7I2NvGSk2N+5KuU4nIZgqOZjo
Z0MkpjDiZVoeepzpLBJxoq4LRRRzO4G1EpNPHvBa1dKx/7qvmY1eJJfk7wMg9SBg
DV8mbPhqcwPKuipW67PMpUuI9F8F3f22CF0aFp3tbH6hDO8DVftMbakZhXQiQcIX
I2wXExVHN7425bpnRUEqC1OkCIbJHxN9IEZbDNJOfHv6lYB7zF7VNUfOrO5XzgJG
eDVsvvZFxvMzvDpEDUqZCEpZ0tIp3lw8nMbz9pW9pqtGlCQ0Wts43Z6d/VosyYY0
oT7ZGoOTOlMOqImrD6jfS8ZjyUy+JpTKTq1EGz3tZdv3MToiCLpPKhq0qu9U+boU
ZUuwYV6IJBZNkscplB3HQr8tPrfs8c1pm884BZIY1LnS5xBLcnNlzLmeMC/W0HFJ
kkHoed9AGh3M8tdfCHtQhcUyS67d8ArbrBxrFpK0486wDft9imaKsAdS90iKzUyX
vNgzpZcR1t2poVno2Aw6nayMItcW9vkwuSwCVKHeDxavBo5A5nQzuYgsowv3spOB
Nak2svvQcWd7obbbroJyaRXUsbloOxoDtlAWvxaCaivcy4kUzHrAwDhOaH53ViYP
oxO3NXK724Eg+p2ekngaJSqETtTQKTR3Fg9gvg1gzam2Iq3GLDYRaNsicOQ/jW7p
FR5QJaF9wV5CWxexyR9FDW/HP1zXaE8nNct1tJqtk90zn+dmg83Wu6INUEefDVqO
mO1WBBfsF106mid7VzzpFNsYTpQiFY3mum3OSFGYE/fUchW5vd1OZWPslBnINFXE
CY8tYL9MrutsiC3zLDEPn+iilbT3gNaOnHmozYeUUk3cZXci31AOqaAdKfT9lOma
v5kIQ8iRM152JEmtmQb498sxj9S1R288YL8rtnONErK1YIujgtg83rVNHxhi9lWt
JKiKdhIZ1UOT15ZZKJIFJ4FzQX80IQKqoYdNyoVuz2mgBMtWvCS4b1/LSqAvW7e4
AAg3PLrNQ4N2l+37dFgoKsXEKyJggk/Tyeuva9pDy3GFrG5QFILJXP4GfMkoUgDt
sJEaUfpNWfNR5X2fb00UDyOXy34y66/rEoV2Q1YaumMGIWf7Yd+gaBkwN0GXROJU
sNDgnThPhGSEZqdX/kdlB1SljjaQGp506B52KvO8o4wbhOrUMHwb+AKniOWal6ue
Jvztf7+jNpPOppe4N2PJ5oqM+2wU03CH39FcSd8RRyVg+m+JpNVHYUtke9+p/h07
zQJXAlbQyka/Rzm3br9mbTvUwuxl1iSjskH2kDcA+segK//ogvvyXFfrPnSXn5Hh
c+McAWKyEonje/G/1A/neZZhGCl6i7XqF6lpzKaka/3uam5rbShCuYtYIRRW3v/6
cllczhL6/5r/LbDztc++RExFUgrGpZDNi6ZBm7zR+7IMKUD3KrbkgvUshbzI2wZp
h1RC55xchI8ga9OUfthqU/8ucvFft2xgmaHRKIuFL2+pom68z3m4/LcFGvtA2dUZ
9ifU4n1TIjCtlCz8fuqmhIdZ+kndSqAPBZ5M7nSn9ynnrvBcE2TVYzuXWpUtuKqN
aHwAB4jukVZghD2MiRIroCUXMV2vNxQcQ6+EMiL+5a4BFvoMezqDsupJTlwouYzG
z9lO3D7kxi0dgWqELSbqxsiHqURaWbRCGFnGI24mcuXr119Wb/tlFRZ4bYH3Ztwl
YLkxgdfht1Md8F9d4wI5CElYDCF1tgKKQUrKkctCHpQlfJOiRiAd6NmW73kLxLQj
E7Sqv9sWLLLxuL70w81PuGNYi1EN4SW7jqseVEnhsNXsze9WZCHDR3Gwl61d3rND
h13BIZXKM0gTRH7xMD3w9KU/ns1waz3KU1Z2l+Oz6UfpQW3c3m49ePmtu0yns85/
oFOBY0OGwY1gdHcYlwcHqWrSwS2UL34stw1UnVBAzQhMr9w6+r7O9X8Ou+ndpMpQ
s/B/ZETvBwMqqB6mmqOba3zAhsGhONE6Jpxn1AzFdmE9fw1IoeX9jCDsXsou+k9B
Kf0Xh3lU6gaIvRKxMhsoRj+n5y39hf7Ty3+TqFlXtNZBMTv5EBM33cM5E9fUJXW7
pSZh7cYeQ2/Tjvq1YyJmzqtoCTXEXTxv3N8baSeqAc3WjJacCbB6/htTQU36xrhk
UXC0LcyeOOBjwQ/LgeikKWWLClrfP8AIZJGQOx15z5bgdkqlWOrlN/6dHNiRh8jR
hRqY/ji22B4i1phyb2IyP83mIiS2Mjzd34OnHTWS9Uuh2UFdHsT3eYj8WFtwAmE6
uyw9is23HHNodANWTCMQx5SbaziGjB6g1NntUXPSN4xrTcAF7CFMZX2ecqPRb4/V
ivFB94NOirpFnc2YrzSzphaR76HJ1NKrU+p+8Tp279XAJCqIcWjMlpFyNzhs4Sl6
PR4/LKfyhXCcgKdEgUR4swPVlom81kG1MqUY3/sf0GtPHbtmqSQH/fptPTsjxvhx
g59Iq6yJD+K43noaJJx5Y+H5Dx28E42m5P3xHbbNdA5kBC2DeExWiQ4ydsYIbg2S
SEyu9TsctwXU0+1Medao6fIxjjBPGu+RNetx3BGIvIoPRyKghjMBDx0/ZOeyI9JD
8U9x2fTYVqDiZPeRf+xUdlxKzXIKaG4T+x7Rq/Myh5KLJmHyo9qoZmEmSrgwItNu
8z3VSeKsnjHB8rdOVubhOHx8Bul0UvF+lD0+Pat2khvOadZbBuHqyGXlemMnXgNa
f44JSJq/k19WmRmyLBAlXYaVPWl9cGU/qYtHwDJ62ba326Tpd/2qnC0PICnEDt+K
r3CzH6LtmazV/y7G8p+F2zG6fvoF7ccll2bYBULVL5awiKo70LjXYjV/Fycm2t5a
Ib8wc/txo6ThJ1BGS2mQJptoihr2VuzF/sjPOtU4hiqxj81TXvZecoeUIpfqBUMc
239PpPU4SEdqit2jL003+ZC5/vQj/xlQgEP5BuvKsHMqtIuP+d+za760KIldKgQM
H9n45olX3rKhyld5u7FMGp+rWTEYt9aJ+B8eDn1sYkLcTGVEy2XhsD8X9HUOgoO4
Mq2xK8SzGReTgdfpTB2OYdkpo29uYfdNYG0uPOV5zFPkpY2PN65OrcLhgNsA1/a6
XUjbz2FfGZPTuzS2abRI9uX3vG+zL/PKFbltSfXIZ7n4g3rHmuYmLmy+BFepXxPx
zGKmsb9hbmF0TASTgPN7s+xjb3RRMUFZ8f/F7L0CyC7P6d0YFR9na1WYnf5oQ0Y+
4NjODa027S23XuGE4mzVKrZHzttj70gl3INOWZApNzEwCnSAJPVNXWx+sr7SOhL7
H1nGOelO2YawTfchSXi0EaSi2CvWD0kgFBMmJAmkqfXqAxSbYNqkyE0c620jfSYZ
RaDOtYbvkSbI+DayrO5+KhKhsGj2X8t1OtbEKBad2yziKeckd1od8PWI7srft6LF
y5P+wn+SKan1XFJAYYhwAVQtKO7kzacFYlzO3xS8Bqx26iDhNe0rWIchquyx5gGU
tu6bOUiDG5pDZq/KznwGlaZei64J26AjrG8f2f25bOBZNiAEDIdXoNA4WHQeh0hi
kTLCKZET93gdH4TbBM/grqL00jp69yc1GkNo8TLst8Vcj2iSI9bdGXH+PY0E1bg4
6d4wmVL9Y+hNFaMAx1IQ+fr/C5BxKqtFZpcwmvGFxsFYUyfibCI9GBu+6frs+H7j
fm+W13+X0djc/bJdwomrdsenBjERLxB8Ey7+vpCo4prsCVM0YgF6c/mI3WqEtb/a
EWfL7qq9U8NeQtNrz/xxl9tkGaGVKLMv432o9kL4bF7YT9yCiBUd7jlfBcVb8uxz
9ZNpVc5JIUGDkuCT0TkSr4TcQPrE92XCG5/pbqZ4NVP3h9rqV+C7YetlaSYSMsmD
IvKf5qoutrYgJKYueMjnwgKJmwSzcZM0g0xX0Fih8bFQdSt7xI+wg9aR979bWK9L
Fc6dcI4wm705oSkdRB6GLHSUWkCbwhGG4C8qDM3JB5+ws2Lu/xUUrU+Oz2c6Zqg2
6oe/1oSXErhQDr2yJccl6W0/8fMYy/qC7MOM3ECNxjmhQY5gdi5+b6i9Baza7O8L
9Pljxy3PNvlNr+LuK8J7xUjsZLlF5AAV4fDw1oyUYAHHs3cV77eF/HNLtdCWQjDh
BnRY5mDL+ly8HgjGEzbi7czPoHcOd5m0+pH99hO1H5g0SS69g6rziaPISsyhkMuo
SyEpLNhzaa31ges2J+7BeEkUwN0bzE9n32INoa0M7rtM+iiA0bPClY9rTofL2iR4
EPT+vvb4H2tgnj7NltuuqyN0xBd842Q9bTKIXe2wPNMdf66FBrdj1RKViy3j7q9s
WcmO7s2TOUV81QBLf90Rua9z3Z2Gu3/n9T0eJ91u+xOedt0By3eLuLCf99d9bjqE
KejaKivSjum/ziimPrsuTwrX8rNJw62SeigRt7RmDCQ63dfbCVgLZ0AqN7yHBjg9
+PwAt4LJx6Q3qIGLad1FUGlTe6Wr8m+N37qVSm1N+Bg4LmldE48TxuxOsNrxfIy5
v7Hk5OiNM0Lc1THSx/ZUJakRlET/PJs/QO2ym/gqolRqvlHl4wD6t7pC9iRw5ndT
NmZl1fWl7iEqMGRXTDOqPAMgwRWDPmRBdBS1DrSkuiI2/VZjzv+edINTBnz9hQeB
+tjW6OnItfVUg9sNQAgtAIg3KV+7X0GL9lO3eg399zVwzkX0UMYgy5FyumfiubYP
6xpamfQHgxKrskMI6LcTcl9kibTNrtAjRYb+H496fYxysiztDazvhj6KmQ+wPqZL
kHSxpdrT0SEJU3PHSXjOPgM9+LSkXMmTls9aOqvWe6uT9bw2Se/onwTsmRWNd3kd
dYvfnvP/+M2kccK7+fFCM5/9WRa1UF9fJphCbYIOP4SMg7qv9zvWr9QFVvHbqSRp
OyjUuOekPrfMnnR1kO5rC09Gi8hGL9U/X54cD7g/P4adBTtZOh3+b/IU8dUx+82n
F58k0LF+Uvz6LxZVC4/K9oKPtdCWFeVKTorfNXnHO7CnISqUFQuV0JqmkrBOuoK7
2Pbem8KMm9luOVCj7tVq9YlkkQ6B3GAI4bO0Bb3EbOwvaGEDyKtKH7io+RgNFTU9
T92fG/O20WZEtuah7aWLKEJTfVLwf2arep97PMwOsBfBXkSrdO4Lo5Viqf4J4H0f
SBcllXZvx31+faeX3GURKR52K+5KFEDCLgE2ak0RGF6+niIqUSuFi2n0dWIR5ASo
B72F9E/R76WmEmyjSXkt7LFijVRcjf/++OZ6rfZP2U6b19ByOAT2xmla08i8LdvB
4KKesRdLugInPu35SIdpNkb6co5Gs2IXPHXHBXNq1c0s73/ECOd4E1MFGdNiiSV+
cN+JgagjVtrZKy54tg8jyTzL085mWPJUTHwc8/HdRRqPe0BphyKHYw/2dnnz4KrQ
ZllZndJnkOj7hPY9uijA/7ZDHyBRkl6D37H54hZI5PJRBqz2gZFW+3XpMSoy5IAd
O4Xl6BDQehHAVoV+wLzPUFv69Y5ek9DhJogl1wa8DqirE4XjAxz4wTDR60F8kRe2
4Fqcr1RL5o0tlWdyLXgX3smIqPApO0bA41nuBtf64m67CrwbsuSlXf96rSj5aoik
Oaa9ZX801S55c/hxeYMq+825KFx4UZ8Fi8HEa5SwhV53mVVPna1YiUqtpl5g+eOV
x8Plv6hfDDk1X50nQFyuCanXzpKlNBsItQnxkmO/l3IvqlCpY8GZWozS9cRy+Tia
pNcRLJI6zyA/y4TNdehwL5+6PgcjNLDumher9N9d5GlWFvbWtBWa7SjbpG9UwVDH
z2uFIomgwLoPD+lqYGbxwrSG5GWoDzN4d9KJ6TV1lrtq7BXYZ7ylM6V7G3LwwpC4
gEaOvHjSV8qLN4P9oapYJWTgHgz7snIpIwQkekeYqgEEv2cVsOsXg/tSz5hxNKGb
lpnz7I1nuIJWTI0dEIr1rGhMINwsTomdm6WcXMSRVsPsP+FRAPgU0LG3QpnZwJv1
OVUS9DddVdpqvOUK+eGpeesM6VTiELRDt9mIZKNIiUE1+Dm+ug1B42bdpvy6wuzA
sEsFcm8ZCvxxgdSt8k0PaXeGClyOB2joPljIOrAyqocZbOggMoNdNdxR+dgeurMY
fZ84JqI0g7g72rvMXacHS7q99Nq9Gmn19d+IZ1aa2DiA3h23Ma/300x3/lqByrJa
HfUqmMjJ8yLshvO9tIn8R3zpiytA9Axm6kwMc5H84UAUMIjdkPkshFjqWFEms9U5
/f1CXPyBbiDCwziPNfw1ZDCxF1cXikfanP10DOSvuKi7TK4hcik6aDtIXLbtwVNP
pqTDn9n4jJeyRBMKm19bORDhbvz8wwYZ9UHhJ//COGAc1nIr2VaDjdVCLry9QFoJ
eLvi3EhpIV9K0vcoAXc3RQPSZJwe4rnOt5dKjlmGFRkUwwsKQciY+tQI+Y63wgEb
Te0l31sPhrD2DzdUEqWnUZTEVwtGMCgah7LzmCI3a/nxNsWuw5FJszcYjVcEY2Ud
Hnuydf0N29nui5UU+K535SgvE7e6LNODdqUkmx2cdfYdODhrLDPGpXkAWfJeEpNU
jK6UY/Q+H/O+dlxSYBi4tZzWxRptGDMJKSVfQ1Sx4F3HegD777SGCnV2i7KMPmCr
Br5EohWy+C1xTwsC6it0NrWn8xEOiF6zPebIu5BiwlzcXt2G9O+cBPWzYjb8Ls3I
6B2z8nBD95/97byw71Fdnq1YkoGjfjjW639SaNdya3nMKIMHhK0XGRA4QgV/O8bt
CAEVg0sxXjgk7jGiFFg30eWhlj8GcdCPAVnWUe+dsLKc7bt2sKOr60G1rU/B02wo
l92i71vEZZUJmPrUvatEdy/hJ7TpeQEUfw5Z2Gidnyyefw6/vgjsKv1fuV31qhbD
Jqry6QvcYli8/HRZT5i9yO22uxpAonS0g3tck5DjCCEzomfnSXBq8wndJ5+2SQrc
lCXwcIK8CIYA/sj4j0lzmzgKuZSMsRO/Pd0gsrU4S8xiaITc1JtRd5fLfjJuDdJh
9H4Iq726zopunN88HlF6WhlcbWJ0KcltVQxjfISq/16GN42Cws+zyTQVNZhKk6i+
HkYQUHVO04MDSJ8jdBfs3c5TMlfleZ5W7XpJA7NAxjPYu70BMFO+IMKxAX9wHbJu
1WcOH3ChwEQhP2zQvnI2oTvOv043cqMxeoT0tvUxjw+KUoDuyuOUAX0qge+y+z2X
LtZrWMI7AgUr0iXpLApYOAQZA63AKnQWkft5zv6/Vgc7Op6suGV6HsSSGV/pXvm+
juAdBXTmMHj606LE4wmiDhv+BRj9mf8XQmMZZPSahlqcrfT0Lq02PJejr+ngSdnH
E3qFI1nSDewASLqFWSIBY4Q+xZ6y7bv9ieDHIFIM4N/TjzHNb8EUgjs4xxerw81r
Vb5hqiNhTiD/me2CxQyU3MgnOZWZxt9TYBS8AeT7QYb09Wu1YXAT2b9Ye5l+Mu+H
YZKlxZSq0TjUZ2YDT4tHxiAFwpRTV8tB78p4ZI9rkBuWl1wGWkCfXG4TOU5K1u3R
HQ7ecqQWaKObTntiJWoGquHPjgcymzW/Yc/3EFncNgudSVvXkUFaadmckOr6/JxZ
T4c16xMAhF/QuEt3XYS7VMMNJJSZpVZYI79uyCgS3nqje2QoeMahqCNhkbE3kNlD
vUq3IuqLfAuK8+irYb5gOpw20nXb73bOouBCEeB5tiiJwjXhklU2wLNlm+yrBJQ+
Fv8VIYziM7dQdGrynTea/4GDj3CU2mEtaxmJNk7FT3k2SmtKwEft4lJquiikYI59
m/KgFr2tIrxAx/VkPKZFOu+4b0pbzZA6Kf9MjprtOOBfqFPVxXWhrmnzAPry5XJe
Tsq/gnyAQxghaB7/Iev/g4SYwLdA5QFkaQRkmQUUtbmPuc52PPCSnUV0LTMYgTA8
aLYtBaR+dF66llmXaakQcO0jHUqH7lW+2hZ29LrSiMEUS0/Be/r0ubiTC6YCC5Nx
UwhlUJL2IS4EpdIYMZb66fRFvLnGWg2xIeGJ+abJlQ9oXIhsI87K1+vykS+pwJ04
2McFQ8vM3kC+GCXt8L6iH8PvMveFJWagsZaDb8V9GczIn/Rwnm+cCtIDcyx+4pxV
SjLTqJZjdI1kta3WjpqNJBVjHtiH0w0ypqe9UL2aiqFSqIsaqMvUFQnkQemrJXzk
JIPlfJyM5PJK5h9CQ1u7MD68UN2scOdWuGguiYmcpLOV3h3e66jUiiWnjBwzRNIs
zw1fS9mw9pIICIQiv7ocvQslOcta1kRkipa98UPhACpqrRt8AuinwxIUDQshhFht
zPFyF+lqf8S8MlcD1iUUfcGeMk6icj+Uc3yuY/ECptgqbbXUw4/2ZSFb/F53iVQM
0OumC4UoEWFrs/Sr0g/kjWwW0qQ7Xf1fvC3N7QOfY7Wpn2xWDXCqQc7Jd5FHVLxe
b8i+9PwA+lYU4rgDZzQy+pU+TGcEmPKaOf/ndEd7imnreOMJP+t+pYR8uJgRnHe4
82s01WoqwErz7DARbQkJsBFC5O4O9pSzqvVcvxr8tbyVjIG27p7bpBgBXI6FeB4C
BzJLB5WWIB9BVBtkoKyc2FkmO1k9rqmpACP+c0IMip3HLv98Q0YdEyGBUkaL1ied
vm6yqpUFIY8L/yp37gbphGif/XBRzRtJOpEAdOwDQqR/wBYrVyQTGauWIBqtFHk7
zOjGYeDCp7fVtA+1k3CM12kkuD5418P3mMvN44d+78V9NZ8NvyhZyzhajxAPKvvu
vKRQHNo9G4KT9Ql+UGZ13Gf+OwrBASEZDm9CCpdQHOSO1Xck4i1A7AXCZS7bzjRn
YVNUp4H9e0oz8Ih0lHhaz4czeBwIcJyhNcZ3vCm9sSe4BMHsezbQJ1vCIA3b//CC
DJ7ltmvnrnYSSlSzFAwvQHlnHJzQnXssIidmHOHDRWd4+2EzGTDHVgSfKZ3F+asf
u2nAreNi9WxUZbGy1mppJxSXhX33MRb2mStuN7Hc1/WDqsEwg4ZlYGqPW+wmZF+s
bPwpRVqW2Ub9lXqpa/2ELVb/9IunksE79LbvZvQa3o0jgvnPWSDxkEYzW0dKUMAI
L7AdteX+p3NT8MGxwSorRlxxlix0r3BLZK++JqwkJamrGXqR/GCkmEAUR1VoZk6h
PMzrZI8sJwl+4TNow26KAI0x0WkLhNkKETrEkbrp7s4VgTPmeLp7U8LdDuhX3qPO
eaiAaaNIFISP2UDdlkLzUxXJd9T43rloMFkMcX5huaEn+hbg9/7gOPs8jbAcZsGU
Mbcr7UoZiJ6/D/KSlwab5JEa5QNYBd5D6Q21xMpJ07iW4cJba16VQETa+NSHklrt
oGfpUO19S/n7yfO/IOyo1UrNMg6Kp6/7CtPt8DqxQQ9nZy6R0VOatzNmVc/6fcMa
9PSs9qTHGgjnoxI1exRT2JuThu+v7oetvIG3OB+e+/hcYybgtYFLmJ2OMRS/C7+/
s2raMKc1cu3pid4kf4mBT8WrYab/XLmlTlhD1AzRrUlRe7AcYbWkuA5cM2EvRnCM
fn65fwmKS5tP17jn+GuRsT9IE4X6peIGbgVd1uWrmZ18CLRQnNSyhrGEOpOVwBY0
zgtTscksbT/tljvdtm7nm5Tqqm4m846WkoLLqSgKlY0gVNqFrhYQ7+a6Njb15Oi9
bhKrE2sRQOSayhAOSFvx3YERq9n4wM9ZYs8GklcnVF9snp57GWIgiKYF5e6gi7oR
RmSOy8Rzl3NzFI6FpxJgRb7kXApoT/boERGrHBKYLI/9Fwc0m5eTgnz5U78DWB+B
9OYsXqSrek0XGAjY9XtZx7cRginSya1qlxOwzsMD0tFIiEGTX6JY1KN15OLFfR3U
guRy7P5nxEKt3+eFSZbA4dFtYNnWIB8Rac1mZV1mpSqafcOa6VnyTHYlHYwyOnaA
pP83Fh4p4dXNVOJ8ekhC23D2x5bBtt71kHPMcwoSAHhIQdjsEOrXWwfKdgSAnZ73
VQSaCPnVAlN0UTk/d6oV/xUgnR45We9J0RXkyDT4imMK0vCmvtIxu9vXQJhflI8U
ygH8DvE/lsgK4WXE93L3xNzE2WJXCjmlcR+qghgKIgB7jX2RHgmPIbcURK+VgjIv
Vu/Vd9Hky9M+p3fGmvWN9fgWwFc9iEE068GBN9sVKdRF1Igjjf9cjAAENBAkILLX
o7EIKuVMrlRew6Socw2BDMYAPFyvkfOceSUNSNeHV+/mHafXHiaDrvC6KBbZLWEL
KCYOjuvuNMjMuUlOh5UhrXgozncQSS79B7wgPzuwfgJ7XxXPCSyVw4EasHYJse9A
hVc6rVfxY3St9F/IH5fyQJRXcMBUyFiXR5NMsa+6m0d75D4kT06yFW7R25TSHXZE
V+vOMZVw4JYzPsiOldUkJVVr1ktCc1dDZztwK+MEh0KUH6OdXHCjKTvRFO5p2nu2
d2IyDuXhR1NUThgJJ/ljatiVEljSqcis57PV4GJvCSr/VTNs99DwHhUNldigjm5C
kikq8rWdSlvik4Zg9SmdUnJ0JIt8j/rjUqagB8DmwK/uCRQgOrDDV+Muz7kfyk2v
djnbQWgjNZafF2phbYBvHzQB9s7voUJydkqSOEjG/g+dJVZ/pssI05GLAUHaqIf8
/YKC52g+BtbjHXSpAVRL8vVffLtGHwxHNkWfrfnendXwUQFDAg7htH6k4c4vOHK5
e4cznpachzgf0N2pUsO3LYqCABJIRLcrnlXuiDL0aUmmhv5/ZvsM0IR6MbaFW5of
kUuuAQkPJhPXREZ+qSkVyYaBxrXDGA5LyYje4IqPi6hiJwwBaL5c7LlfCDMc1yMW
m7EitcLZOX2nSBdXarBWKzkP+FyWMYmBH9LLhaGHZXFspTap80an7YZwP1FFzeV4
Wqde+DBJLgaLblLLEy0FoRuU8Hu3EEAy+xbn/eS+RwSatQ20s7jiHfImMuybkvOK
2BxXbXxPU0X/a1DCBhUwLe8H+wJF2ZPUT7WcOhfv1iTwXxrihzzUIgrk/HCXqxs3
eyZGBzqzcCphOrK1bR71EOU4YauFH+lEIrDYSixh3J0GCtIhoUjTVFkcBERwFZ7J
kBOGq6pFzULGdZMuxXndWEd6kjH//mARl5qZSDKQin5/BUxdQrhKyLhMktldQ7G+
mxhgqFahsL/rSlknxER3Fm2EifbzF5H6xBTgJPejxKFgg3XO+VH7eqmv7wiqqjnh
wIZEsLJUoMWunkW2dSz0lbZcLzu+WMSCH/6x2HJVBHFKIbtrP6W6dB2fEsVtyyVQ
fTUfldoQiWhhMOeQQG6epZQygx4US9W8etOzK4X+d7rULP24ocxI7RUrVHvn5B0t
Q+WczY2qRG6OwzNZ3Rq4aMDk46cowKsa7jSGet2+/23pgXFvsdM/46Sw+W/nCkyc
tLlyvzY1iva+EdgCzlnUwtIdKhbuGc51uQ2Me5keORxm30aYtNmz2dtPCY4sU+4+
lWVG9wEuL2aYZdJO5qeoFYUhrIujUBOUnLthk/ssBkwiAq6UzpB99FaoEAwiaSAV
fnc3sL3ml3JjROd4DilINCiqyeItHSrcwEdmbfqVR+C8T8UwlVu2ja469VBimgW8
T5dA9FeMs2ppMhL0+KJDu3Pd4Ctx02xFYFixn2hUZz0yFuQVjun2R/p/AVZs4UUF
/OEB5C+CYsDjHKPoqM0ohKXPJCcq0NvGQAWlK2/PwdgUySr4Jvmzzq0c/ikWRFD7
TKD13DfSzGRAxT+qfoqhkwBs0ftpGXYaRMIcPlfNi87P2Z4bUtE5azHBoxlJi56m
Ama+6TAsxh4IVlD23pjiY77usuW1NdFugfjf6hQVPfHyHfo8P/Pd9rin53aBxKLD
80HtlJjXePXkRKHoWXrU2HNnrp+L1HSxTJP1ei2s2bbteNYtZUbd8Xc2x8WDVTLx
QjP22j2qVZoCkf6dSregbzQ/YQIf1ecFr9MgcYH+Nl5CdhSAo8BPshWFV2XjZ/O1
vcPld3QS8kUynDc7HK9riVT08Y5aMyhb6G9byKqPi0/USlJF70UCb97Vv+BOEjqP
PCeSyI5iEPpgLaHilx5U3mIg8XOkOAhpBpqBAj7biQ9q7tTMSrm7jDV9LSxTKyzF
50fpg7b58gtqYWOUXpkH3HeIOwHoQx6AG40tHCruWsfcxKne/Rztf8nnZPZt53o9
C5SNj0nzIh1p/Ob0jDLo0IbeeiaSkht1soFItEIo6F51giioAN/W4clXr73yhVkK
B4dhFXJ4uJSFpmjmnSx/9mUrxqtjQnNsg834Y2ceQSS5/jV4cdiMYWYlbKbM7UAh
aHjqMV1+1QMo6k36fEWS+HzNGTsfDNON0ZWtHkli5NRCS/gesVNvDWGBwVU2RHhP
4oQUWtkKV+2digcPGKiTYiUVZlrQ0pDefV+YEAN5+xYmr7MsIGkCdzAkWFAkV9h0
e/e2Vdb8/DlR1VBqSa17PjpYGJuyPoJVAt5KKzYGLukvuYes4/NALLe79DRjMZon
T8k6FmHKWsIP/TqM4Ac8ag9PzK36Rif6vuB7ww/MOEygkK8e9S+Nw9nz7c1VV8Db
nW3eBDRUBmUKEhUCz82uUdCEMUucMLr3bS030kGkfxAHBGg6WTf7U1tTTCGPdf9+
OnFdMVEYmyH8k7wLTheFUb37tUO72ASCkQMbr7SbYeOK4ZawIh8X6RySQE3dAPvT
Rp95raw99DMDNCoRT2OwCkQFIVgHMCRWrG+T1wNtlicMRm9NTG95njvAFMIALLMb
9Bd+Xlo12SisWOe9QpmLMfMxQurQnyALP3f96tj9Gg4Gc+irRH8M4WDtzNypJrq2
ZDbSptHKhZAl+cdsVQ5woh8BIu9ScFUAD5azVpV/7swZjOboigDz0jcG1RuMjy9X
PuzELDMyXGMnSv7opZlPvWWbXg2cMnzR6QHGWhPMdtXQjTcv6xyvgI+MI6v8Ix+O
VxuSi7Ug9isCsVG4F2neTEpQkkfmquWrTwtvlE+g4THYIpYkjegL8lMO5yMZERZy
X+TPrKm+LhrVb5yJJPoenv/HpTzA9Tv+XK2fhWjeKEpckQbr9lGaSRlWxVKBzvRz
5l91p20UVHzeSWMoITudmCEuyAHYZvfyeWTtsO5JtZOCg0GFO+RlNz/iiFB3KaXh
H4E3RQlMQJ1CLuXXe31XoD+yeMmL6GFpS9L5Fg2Wu1Zt4qfPwzmZTlS40iyIqVRG
ES1KBvQ7JQD1JKE9knB/sGZ9xhBuLgw1BDsV/moB2cneJiwZzmI1DK1EFeAp/Lns
UZ5o+Ja9YngzDjX1Pgwt6nMgAAxdIBSIUCxgjKK1nXbFcUPbVkIOmfEfKVlF/5+E
Bl3M8sGnvDaEOtvdWun92Cuz4QbjiePq+PJtdvOKlN79sohBnw4c+kG7gSyJXVbC
stVx0mR8Zs+xGfzvTosY4BB5UkRnEBRL8jp5o3ztbOMRUMOkgS4KB2C9kEV6KUKm
lrkZGW9LOEIfS1gseslVC/ADSHiWW7dm7z7XcLidvDm3OfLVV670QFvPid4CsYkf
1MeCqRKnIYUo6LY0d2flcam1bimKfZoF0T7j6g0u84an0phG0sIkoAJoSaVFl2Tx
guj5pykZbn2HLDAGrBm6TSpi6vVhlp5wyFDtAvtzo0DNy0Yz3LtjDL1XYNYzQ7uD
vPpmAhSgpfBKTY1SMIuc817uVVSTT2/opxilKDF+m77WZXLl/I5z3TCvJ21GMeZx
UT/0REuNRL7hyILI0WlmA5BG6JgKsj8hX6/dYYkfJH9MAhdBGFSeHWAIa2Cz+CyK
yqHL4ieA1Bj0sZjc4GTJsws3QRpLCsjndgmUjNNsrtfMiJSBH18G0HA+3xbI8pbN
x1xjS6cgTm8crEZPDwgSI6FDpF20BUKQcjTmJhLH23m1QJq4HigHxuEXMhyBI1FM
NbNTEp3Z1v7Gvhf8S16FoWNQ3GZO+lBImnEg/uz5voWxQ8Z6bi36DJE6BW9qCevw
Eo7jlu2GPpCo03weDSLMIQLH7DVy9zn77zLK919tGh7G6T9iW3LtGarjG9NiJvfN
jlzmow3MnWtfG1UoTAFuk7X4UFM7p/PTpkJGfKk6vl5WO8F7sBjaRJcbKzPu4jlD
/iiyy4Bl5kDgkQWBSND+7KiNV6HsB3t3o3e7hkBzx3/Oy9zlOD/jZw7oU1jTvo/v
OJRsa+zt2SNIEiOORoYDzXZJM+L4esMveYETKFE0K1Ptc8606MUGLUIP0v4uj32n
16iKBiopDA9xSJNPXgf9z824wf/sLT2p/0+N3zqRI1dlYcvXH4Toriqy2CahZ34C
8tgP+tj1D66UwqtgAtjrDUGisefAgtkWZCvlTlWRV5eFVF20JYuNDvh9DY+Z0QFx
hZrCe3KqaRYBSYrlUocWaxKuNgTiQyDN7SOU7c2c4sSsKGGQGFMFSrflzwPgE9hM
ufnFTESU/FUhzt+vl41i7xpNZitS/abBFOoJA+g3utzuigxKhoIEyFxgkgirFSsN
Kitzc8fkyHmUZn/uSjeSyY2WmRNKZPoEGZzVjjz9C9YIcchhtOsQbYcEXYMKpowg
uxzpenO9B7rqZY9mQlxic06G/bx7N13hZxzjBXNAqZdhzYOa9VvyFLT1bnFsrR95
v/zgpXULrTXU6R96srbNDw6NJS3hso3I/5IJf5rqZyz3G/rop/BG/cE1CUdLAUjY
2tlEVbY3B1hiMLQxsAkg5TFOmLPsMvUIP2FFypOFzSfDYrMgbEoX1S+tlr4hFYpv
R03OH8UHcXzgOA2wmkyA0uINW5ofNNTwL1UzmWc4zW7gacS4zJ5k12liF6jUuAg1
TcgDA/K4NO1zlQoSJeyaDGBouXhZUgaKniifwIPcEGFgh25mOBN4JOX8xDDNdcJ5
pR6I8a2YvjIR7pRx/hqXKm4MxTq3EBN0fxa/i6ZHacEZUo3scKkwkUr4bV+Bgcow
d6NdGGYyMdNQ4ZIZhN+lV8BXuG8hl0MGW3T9Z81QwQKjsDSojvpHfcf3noelNht3
siga2uCkz6TuyMnQqwEJlneDw3/P5oFiWtS2kqfc+HnXOrj/vhKVh1WnvhzJmv6A
KXrEl2nnFWqS695KllDtJ5eRTQN+HmS5WkJE9dYKdt0otfOcPxE4CbW9cq90QlRB
PUVetKTDr05ozu3pREvmaVc+YkTAW/6QyszMFWntBQIWPRnrW//uO0dwAIgAbIMr
zXHkNRmxahHxdzvJ6b/tDNPNm4Y+Zfx03maBTLC7VwsY0NxKRGk5V2Phx4gywqQ3
488cuy8W6UR4iA7wpk3yYL8O34YL4jmoKob1sb1Br4YMABh6YsZvKGQ7paa++H0P
INWjpNU1j4DJpiicMiCvgitiCuj0Z9LHkXnBHvZODaw/AlvuJ2AhuUeGPjD3ACfR
3HIi7XhNrdjikcgjIe3OoTmpTgpFKFEXLMTisTUO9Z4+3EHrMri/FOypBRwhDQJ2
rz9nO7H2m3re89LN3tON9VulMJp27GvLKn0ovtp7psbc4tNpOqN7drdomcC0xZvR
MqqPFYGCgQrDZPOsYTXAYixwQWf96ZsYCCCeSJ8NXIfCWXEcphfNiW3alZbXaRnM
yXhF6dm7OpxnIoLWuvmum/Mk6iauxm6kymrVwTfGOAW/cBlzpDm26StyNN2RXaDw
9bNXlFNWmRUUJbzc0R07u7XuX2mNVYEZXPdGkvVbNb4AEzeC0frbs6iBGu+MeN5H
YP94k4qblV6qkI596fLZMv0MPcHAraUpvU7bUJAWzeIV6SH3/QeSJ79nYHXxlThw
2tYjR/ETHjtefnlGl6h3za3wRcusxahosbFljV11q2CH1mi1RcHuy2YDYMEHwH4i
OvUHyAr5F25qDp2jFRARCuAxZoYuOmZu7sdR/1mwFyE4B2yIQ0k9l0jv/f16dYtO
hVmo/DWXw0HaKwgbS0zhrt6Xq3+SMKVtQeGERNZ2sCVtPX6SiU/mMjzCAzgoFPmr
M3j7kg/J2mJlAJ95c+I1y8P70S87NJo6BlNdO3wIQYlmISzkCinv+J0X87p5ghyC
jPTI1BfqlneBaQn3BdRgXiEDKfYP85noqimuewE86WLH7E0lFis1t7aIVndvFhkl
3ku+4WhrJ2oOYARBcBSzv09dXj0Pmbw/eBrPZRQ0VMRM8K5lMjjmKAbQ8ftcqaCD
D0FekYNw5xJj2XLFiYVq1Bk4Jum8SIvRr/XMI06kVRRDM/Z6VqdHJFg2p8Rrx/6K
WSiYs8VjBY23a24RlEumMzubBPQz3LWlkPzHuuzrZ5j13r17J8dLWRfpHOXB5i/E
5jlxJUtsP0WiFvK8v7dFrs6IhQUyvINJv5uhLJ4IBBNaM0RoWD1708hFhClycG7/
5mzWngveA/6qF1HC7zF5ZZmnAobeA2j043t+XIB6fRMdtZ8otVCA7Z8+LNOh4sm2
fHx9U6CPYcuXusRW5OnMGoQdC+03gQRvV7wJqDk6NRuPXuAF9E3CM7WuqpkeQEME
pZWCBKQlMAtu+vbW20crBKmyHuS6hrBQOjnageOK1OaEsWjbDnUDHX7jqi8QFV/Q
SZRCnfKx4PMIrmmp3DyBVqBV/RRiLFxTkC27NMebLdvOXVwzNFeCB6P3Y/39ENlZ
WgkFGIJzvK+gU6nqv/kaO80NNrv1cxgdpnW31CBtYNpkZ7ZelbwrK5BF50q1qLjP
8UxhUS6DFuJu73U0XpcwSsI3p8QFHBsBZ+kOHmIRT1Ra4auWz7NlXUyB927FctMh
A7uZinjXPD5+TlWVzR6duOfvQuZHRn7R2NnQ8yC6OV2l+AfZ1AYIZOifjRDXOUlJ
7/LFl7LBi2ggTGBTwkcaZkrhcsYdzKvxie3MfrkUAbv73SipR+4VVtxWL2AaZ08q
vE5rfimKe8bM5PA9mrSdU4hJ8obO9AF71anqQYGFmUNU5Gmpvv5L5zgzeR2wNuet
GFLwPL7F/Hu3UxauW/8qG8P+XIpMOOJQmRr2wCQ1xDeE5SeXG5Dqn3SbFmWuifGA
+Wb7tsuSvIVmk1vg0szWuxCxuXKkmMPj1cE4GjfbcUdcIYNx9Li3zeJ3553r61rI
somNYR9Ku53JGnKKo2cMHw9P/uvUHErBQdutsFnLdRQP9NyPBLK3U3vbaRMKDTMt
yJacr//g9LReUvO75FT5jRaaCXuKssUf5EBXYoa0XiXrJMhwzg6Mz+0mWMDIyS7H
NCAHyTKCn1eSoYpliJR1xZD0M7T6gBz6wlttk+JszJzsAixGrGMrUnv6yIbs3I6v
pbRLUeEgJMtuOSUeoXDYaH7fYC3jx36k6cnyGgorxTtsLRjOXBxTvQamTFycE4kQ
9XiK+72HjQg4JQkIqG3P1tP+hxGZlsHFkk80Y8DitFUIfEKQMpxqN9IA+VQVc21t
xZr4qSWaGjtrOB0AqJO2Gcr3i+XgnTDIlS2xxIeo/5pqdSuBS7IQO+h3ZMyngKc3
DnoT48uGHcmCFeOLlYWzacvPBn98din9ujT/R034pEvVHiUN0RsAGEmLSPuSqKa9
d8Qm9tQVbC+wgLsXWH45pMIM/EI1NOK2lINHyEop5qxqg58AnvS4BKb2huZwwrfq
ErrtQGvPfzMeP9te4Az58ARzLmrmu9eS7YfHONu9c39rBmLC8oj9b7Ofv5TYWVvK
uHJqQAXKtLQGRgfZWPFwJaYx/Fi817a+Zp9G4FaewqIklUhGsxmUNIvZr672ZZCg
m3kuUxJnuefgUXcSFjgr0T8SnWZP+5qmBnAMlh3pn2CDxnblCnvQS2/uxD/0sDTS
Ch7pApJ4/AV2SZaHeFAl/3GMbIWGK3jJ9wr7Xwh8ajnHBG0w4EQ4/MCJXoooBFyt
u5IYQC1gIpDKcNrVjmvJJUMAF9iGATCr4i4FtPqa8vDaez8lch0npWHwizz1/Xon
pm1AdY0ylfu8RYXtLYT3hQ+m7brFL+qvWfe8jFZyDZqGXWdcf/ZRdp5UNvwc0AaZ
sDQ53AOz1N657kA1X1NRpzSfr5A9WlCrBdCuiotYg85f8O1NIrG/jcyGbvNSF5JU
G8KQeFUsCXzeIQjm1XtXLVL0qtKNWOmQVryv3X7wC04QIdOlsVlfk+Um7woP0OGh
Ieq4d7XYXSmeXFZu1zFtBbLbxJuyLP16IZolwo2PSAm/DsWw+10f8C+A1WNA/7ex
az6VigQVuykGQ2/R1MR9dEkJEi1iVVaKt1/q/JdyvDu3jvL1RtbrEqJG1orMmrIC
j2fObPIkWZHwFvCkH8nnDy5AcWG3uxBemrvKkSxWCo+HmJcWxBzNzZdXmhAEkZNx
OKoxlCIxiizaRTtBjzE6jwOraoYiAVKknLNtFORJce44HR/gSK4NKroipNW3bB7I
T+xcEdEuPNwjzssDeeM2sFnWQ5bmKDGSoue0RNjgSzYUQ/lPKtcvgqElIAnNGBhe
hQGmMhzbegCybSPzRNZ9aD3g7vHRoA0UIOo7yMP35rSlrWah6i4/mSP42vW2HtLR
5Rsb+eFH8ndk0XWNgwougL/KT4V0LqBOxMMMtRS5q/qgW97rvURGBjNpuXz2HW+T
Q0MnL0wbPOOM5SfJ1HxBJLgTtjvrClv9i0X5cZMhGGebg4XaLITps14HZ3GTBU5C
jsOJMEICyM41TFJk8OVI50a4nc4nAp+145IuwmT5cgGIKGcXZEARlEMrQ3bIIDnV
Wv7NQgBjxASsCvCNijZUz/k76UKCdv02EgcYG+fHrzrPGPqpmBK1z2g9wwTFLjvk
3dOst0VBoZfb2FGlw9b+9qtpEFwmhOLhB7TyGGcQ3brebLvjbRpMe+csGKaWdkMy
PoHkkZ5kTGI6GVKhv2vyPwwvexB06to1PWN1MOjpEPuE/2NMU3wWgonDiKepO+L7
Ey8DTRNZfNxIB/ggjJJ54kgSP4XYUl+6nI1QShCvnHnOS0vLgGCwhfLRgcTEf5Ow
g663th5Sw+VsoMBSvHj/WxPkB4nBYdPHjyrBkegrfSFfmlE1hlIOsfFaPdXrykYd
9O2opY6xBJ2HnTWf8JUPfClr4SjYDONVWaaRU87xh/C4OxGGA4CATmusmA5B0zTC
XDcbuRS9WOoQbjRH3KacmY4ArVR0rlsRo0AELC1mbbfKDrb6x/S5EhcZywTDE6Dt
LQfhhqwsVEhJmdbN2HuKYLU4KH2reEVkLzmuIUh798GvjVkErQSvqC0cyU0q6F+4
0tEJP4p/LJkrMYHyGJSuDJif0+kaCokO8XpdEAhcNM9dnCd+VHCotQD4LDLu2Hfx
oCZVdpF0D1ojv4dmlssqGROES3bNGXwO2YKD7Ry8Mq8gP/iTZM0sT1a6i5z02Mbm
nwfZtFf7YfSWYoFFmep3fM26k5yGzjamriL9YpBBciB0Re1lOr5Xc1Wx9s9M7nEu
imvd969MhayelSG4PaBL9Z2hwvQptI6V8+KP5GZgcew2WQVAvfCmg0B2sfZ2E2vv
blxPqDFHnBniVGXai4fXy7k1NCFlZslaRA7468Bjmgz9SlS38/EOr6wJQ2lQX9Oz
GHlbCZuVf3PqQE1T3dUM1M7wrW9KsJ+ouQIa8rx/PqA/UGgFTZyILNhd7i3xBebY
bm1yy2VxHvmTvRupm/HqClIwx1Q2r0HWpfcny03FxC6Tl9D1vhm1LilymDPrw21o
nlNAa5KAtq5fFeG8nZD+fuGNYgWzAxFuK/GQbcgxLvUYkVGY5GrLGRQ57PTcWpsG
Sq9BlBGYi6ufJ20ctyddSau+B+2o2I1rodC6+5rJMUeyFWx3YFf/ENJPlU6TVFny
lrprLKsUoY8+rWMIJF1Kr4rktVMKuweitZrDSa+SXmQnHXjpHTYIXdWTkMbG4swa
cZjENSkLhs7zyE97OMsQhHH+zQo4oYkVOiioAKwN+4EqeAxaqbC8vZscmBGEA7iv
29kFVowyrx9qXc8vNBv+QDMkVEWmx0Vz0Tq1bIVHMzY42MMawdM3NFpdJdr2LuDM
KQ6TGvfL80X/uTBpZAwxFyR3Pm2MHdBynWAoQaHRpm1M34dLu5QS4/UHUTlb58eW
hBxhMrs5KvnZVvSSAvdq7IKdN4XRs193faXOZ4XV/EDn3VUaFeORtdyJfQboL4X+
Ixy6jame/pB0B9AhQmvH4VVyuuZbJrsDgYRr1DU2XhXSYkKeZtKewHYDhurH10zs
3bLwFsfDLeLBKLh6BrIwPllsHl3MVOCTajKtT8+HXb3SE2DtJF4zA6Fu4o19H7iy
2BepK1V7/I/gye7n3KdQ7N+OjyYcL5/HmqZt6ovDpgG9XRLDPqPRXCiUX0opyT8U
RsIighNcymDOOlyKfZtsjphdLUFR22ivcllEIHq+0+yZkN8FODI7BaAfkDI2z1YS
cGVgDXpdSrsfhM4ZFvu4QtkMxnYcCmIO/1p0zmjqKmwibBDDr1XiXusD6X8cwz/d
xFyK3DnsgsLrrNH6fnklPdwEiEWS+MGtWP4H4ErSzwgDzC8mYKlvJYjhRQVujRN7
GtWlqz693/LAsGC3sNX9Ma7zX2XVtDjPsQKIhpLYhvwFHEseZQO6ZDYl/yQd9hmq
hXI3pBGiDK3VdOglrXHVZa/jnxIfv/EbzKARs/7V3tTgBn/fi36GXPiiqpYCSryU
G5SDP79a31RLQNpV9GYvB5gSq8EKQpPNhRVNJR4JlT+Edqm0zPJzyN+RVRmmOHDo
fwNtNLtBFVH2MSVGNQcsB/IO08Sbd6ypXr/4N7Ar01eiAFPsrxP1/cJWsy4hGCpN
OMQvqMfvXdOqUBGckZRfCebynSVvxHxwKiVQRT5SNVOM3UlZPtIiknJV2ZAEPTpM
Fnfjd44sRRkHlvKYiwTYxYQG8eiLZEZQOOaHMHGMN1f1qDl2oU8SJrO5fElOAUCG
BjJz9wH5rnhLfcCMnQQ0RODoK4llWpNY26Ddvb7d4/yVNmI1GqnqQfTiorjB9cu2
ouhy/KTTc8b+wGsR8yv8egCAvDqNImdZYikSRVVne9hnC6E3cxb6vAgt9wNmilQs
J6RhcPGEvCNvD0kQHHozjmVtGM0w6+4OTmV33OguDc51Y0RSiX0N0dTpWX/Zy3jk
YgUkRHURgM5rrr9alYRTxnEi+E4YzYO2GosxBvkAqocX1Rexqrq3fy3AZcgVEkCN
JB7SvFcgLqrYRw65fY2pFUDFe8xMUszeccl0iLDOdW93u/1tqsiUY8kQXI91UCoM
mdtbpmDbuvaJLYW7iFc0KwVIhqSy5Vkcqo+WtOgqk3wKC5JJ9bJvic7YCN8oJAJH
O5lmmQEGygAXfgsB5KOwTDK5rikAQgjeQzHs1Jj5qXpwtB3TaylqHpMtir6CTPst
Bdigv6CryxTBKfBJck4iQsrriackRgAgTXdE6mc2XlMaLX7dnKCYfrR7EPhio81d
goM1k332VLAJ7CieWE6/sIoHvG0xpWKbXF33Cf6gWu+Nz6bOUoLAzjPauxnFUwKS
JdyvnItqoXULph4JYVSaZ6R5D90EIqjWBc8k/L6DPsgumqDX7cPfhsbEy5cJf3MO
bAv8IMjipaLSI1/3dyaeNwBaZEDfnk//czWNrBnySZwtfkLkjl4uyvOJpcgDCCJZ
0u+J6fdQi5J4Wu1fuBjeksZHFKBsWey7vKgO/zMz+Q2tSG8gq+cmDi/vHKXxS/dx
fDPEkUL7HiUC2e15TSoZ1EyGc3yFYWZrLBtsNkIWOQqRBhGG2l8EBiVqmAvTWqyN
SwjjP5HZK+PfJ57q2hMXi7FLS3qrT3y6cyVikORxadmhOOc1JATqJDLxC61XIO+i
S0FU0svL/Yk1Tj7HF/VgZEUSXch8pGALh6WD5JkRzeutr3TaRssKFzKYOfUjitMp
kdqbZJ/NKI7wslv6rs6GVzD9rtxQYqrFcqPbbCLdSUAttkUV2PxaOykpEXGRtUBK
DJlojH9/Oevx1dr/0/zwKBsUpra4qegp49wckXCnjGPcn7Dyu5rm3nAx8aLufekx
sSHI1pwXoPNgxFQjcHylfCpwuO1MAXbH05+bSZgMlD/UQsgdqUpGTPAnC0ZHgKoY
VFs82O7VbCeNKgP6xC9qHvUy6A40NPBHxr/CfAB9rOwnrq6q2LBqsUdZxrhYCP7d
qfqtP+l1vSWVjbbv3Ox1jRuJAkIxLebkW/qOexcsHfIMuwuYuk29HEF0go36vUHh
pVwbnuERbad6+vXYZyDP7XQqJ4vkjPSq6yWw1/VF1v5BZZXE9BYrTHD2q9YHhp+X
LfttZt0C/w2E++k10nXwZONsxkjzr8Sz5IZ3DWiFvtRd1FwAE4inDBDuhPJnxIfm
BlmWE78jjefodT+4dYgeV/G4wa2ekWm/hFN3omUm/gxx/Z3ubx0snFNup2Hjr+TX
Fyevy0TyZVRCRqttz0DR6J6rAiUAIJkoFEVMkev75CEtaFq4KAP2pa6puFgtW9Q4
x7tIP1rUUMHWD0rWxP2p6I9RnX+Gtt+qWTf4WkN2K7NPC9DjTmll4Ek1ZTPpFhGS
6ryfouNqi8p4HwyCcM7x9RgY15qD0Owu+c0PgmVs/q0w9XrcO9evRShhjUpGZ24q
xm1pdonw1Sp60eHTlvy0Ku3GxnJm3AElISil11iAUATQ+T+IrBA18iqc/nnAbcfA
9J/mxFm+UIvrWV3BNn/311S6hvVb6EYJSgiA96Z0QQl/Ap6AJgu0KPGwPS88WNS6
bZPiz6217FXzZGli6o5rWhX/1b3RWyGptsxJXU59qUIBlqrRtxLGcgXjOQ064cZt
l8Mt+QJ2NY1p3T090zn1OBZZ8OfGqmgiAXU0WRzO4JtKMmDkjreDLCR5B3CTGTRj
iC5YhcvwF6+JoEGHGgu8dIPIwr3EdeGWPrp4pS7YzToLVeqtOvUBqGhYXg7DemJQ
Y7KYaE+MjF4upzRoJn6N7Dm6Ed9IJXgg5++IunOMyMIPHTBt9DZ5iB0YfWyrPypx
UCKYfrOk0ZeDPojmawSEvgbir0T4hsDO174U9nXzDEnnCyjZn7MSh03ZdBf/eO5p
WE+JWKMdJTD0MDvx9KX+PH6OKHheWiN3FNvmjogjHx/rkYa+pNBy8gDIC8dA6eIN
QNKW/RytYyyKJOHEX9Yp3ax53iqaWuAWsxk7iNjSxjikQuu6gkLvZGy+B3vRlwk2
B6/Dy2BDIWHdGrrjcZlzY8mgPqLvDRx4Du6oKRZP7ccU5ATN4m+PwEfhYSOHD74q
VygzSAZsMRNNTUSb4XhbkberPI9PX4PMkTih0zN6qsbrcNCzqNBKxvxyPMaIyEZk
Z+Hchs0CBl46DKKgoACamFOSy8ve1a/T2kqtDZTPP3Elv54f3KVr8UHRxh3Wa+J1
bI9nH/uni4po5t9aiSJf3bzTPMTU4/YFZrdAgjhgsbpZgkrABIUEQVyZPhgPv0u3
YERh/r+nky1FmSskkvSMq4zQzx9u41VyTeNa0nu35p+lTh1006umRg5e1OOnUf1y
5l26QcatM4mF1b+a9lQdfhUukS212FL2PBgttOMa2csBzy6dQCbemnTY6gHWR9cS
D+ngk8teBHI34m0tYuV35WZBk7Kymeb6tOArjELtt/BBvWPjQuui5KHLui02wX5e
3w3dNlfCvoPffjEqNEaXfrbES1jTMvjdKXQJT3YQavk2eKAfJ5iGGQQDw+cuHePv
hVHLD2ZO2tg7/RSt0I9SmkDF76kprJX6HUqgB26Tc/VnyQonBV/ims2bNmevyaL3
MdVSw4ltYR0N2L6nLPGBzKU52t9hpP4EBmaaiINkP/e6/uIgd61nj3GcFOAH9pYH
6j8FYBcuIJBOMCcZX5Gpfdz5SMTo3aWZUiRekYg5iWrnmFgGAKtn1yn2VjRkGJQr
t2haSjHhYPp48Q72qk3MoziMXFStmLB6ZdlcHqfBAnTlcB4siQ0/0COvUOU8v6n3
HTsw/8UhdJaQgtUgi8chZJLT1PmBr/9CvZZnAF8A5DSnS1M1znM30jWys3A8D2/s
ycK1Ow9Bh2Hodz++/IaYeVz0yPdcyM5uKTJ2CvWVKGxtD8Zduo9DM0EGG5ACzh15
kSiIgTpl1UzEEPnMFhdMzZZ3Qa5XUgZcDbja8ggx0+Q8tECRUoOPUw+QnqZ2WGkD
bmhUXsVEKEd8t3DKlWXb5Xvo9iMZF2rHEswpk1DL/Lby7l65oOP70HjxRUwTNXn0
eBgIR8QHs4WajKG3B+1k8WjSmqDPNttsFeUatgHMb8crK0pg2pwljEZ0/lP8nt4w
GHMPfQoDc44ETI5wRG5sqdkzUkqIHuIJpiVcRO58BuDflzHgoflHNjjPnm6V/juW
7WGw4ZZTPRwhedfB1V0j/shfMlIPORE4LWbV3hjuKd/LPE0JKohe2Z9GTGalu1hV
LNGG50QQBfeGBJbVcAFd1zhBvDrmXp+V7M3TMnJrT/OBhk5m+b0QLqH23tHiGHL0
/bSQ16PkWy+UkXnT+EAcOd+MtRbqmQzzAiVq8PZQCNUK4nTAkI0GyssvZAzmXVHg
Zm/0gM+V+nRjzOQDNmBmZCvJPUPhu+9XB6hVVytgTj/2HIcqQ+m1MJCErKkIy5qL
sJf72SWcSLKArPWb7/3QzTYhE6jDJ/Yj1hZshb1+DSrTi0fVR5nl8pTuZTXa8W34
SfLGNRSmB1CYcY6kD8KVUtTlf9NZ7yTcIHAdnkE5GLp8OKlI0Wtic9aq93bdWi/h
D8agDEzjPqa1L90mIZKvIfglmoPMh37uWYpqotWnfyTU2KZr9C8mZDlM3ITtVHzt
hddY/N9Jx/p7/VBTEcCCTRdCYDe0ssIDz7IJMLzsFQd8dlcofO+CYgwl5UbgwvN0
vbdHqZnH5V9lWxhX8zP2uPIPBrQsI/z/c8NROa3NbWzGwr5o2grOfhr3p6joIK9H
4hldzAkp5AOT0dtQ+wlWztPAS1i5bVHoWdEqrJVb4W7gDfANmnERONhVtBQVVDkH
gwfpgGYvMr4nkQ+aNjGlonIPAi6PE0ofZ/JTxUQ58RSlM5qjqQCsqUnXcCMOJcix
mLeQyVIt85xEjdoII7kxSjCpFvcMctgc7mlRAQ+WxmRYBsqUM6CysAoJy/RVN08b
pQU8Nk7yM1X36zFV6MKmXCLVA7fVaGnOivNfrUWDaQDv+4XnWTEWXkhDdx/YSyDa
yUcaoG0pp+Hx/BOk9sZITNWSbGos0WDwxgyB+oN4a8wWMX5YrrNn3EAcvYzTRFYz
iTmPe0xo95UlqaE8lfT0QX/MWoGFMB999WbjlPu7oZmApoq7ehTWSj2eJwB5xOkG
HV11NY/UNo53vP4SUaRo7ZDVaoic/LZQwfqotJne3ehTrOuOGRcVOhRlGICIsVx4
Wqfp5N0viWvu5prEg2hygEi7aP5oiwrFjwnbyYO3sJP07f9Ef5QaCTp1+Fn+g1xV
niSMCS6mXgjE1hnDbE6LRBxsjwmFBzcH32gwpUP6pm/ffDUzLuqUKX9+GebqMYZU
YfYIOPQ8MKjEjV9JtSj9ftJEuAGy0KvJJJyQGLywsDDjrVNFJc0533NKNyNRvA8+
Bym1455ZaYXq+o4No/mtHf+36Gm8TkF2gsPxEHSQmX7DaHOmStesnjzi9+pP1Zc5
8WpEiO5vG0oCkQqVqll1LYE4cnA+T1BB3X60RnIl2YxSiNfk14OmKjOxrcYUncjU
AT6W6OQ9CeFUR7CH2Fu0BC+ySKzeFJAm9kZY1wLmZtIBNxTKzNFBWpdjOo1p1dmI
rknC76rvx9JFUtAzJYctT9THKOiyBluM/as4P2NjEw4ezxsIWuCJ1hgK7gf8np/N
xf5asrgK1N21xcuDzU3fQPHGCK24jJsy9HlxxKAHWMpUP8jW4WvF05w5XSsJxOl/
Gu3xct5HqtPyXQKJGpGsEFpSafxyJ/T29ZOqN65ego9XUuykrYaSFw3fiCINMYrb
58cYE5BLbDxO1J8dozc8ay7ad7epN4Sc8tApzFkMlJlRgtJkouKFAfBd9aHQro+9
fQq57r5TxMja2a1fxLL/Tq9SVke6ZcgY8R4QbZ5jS47YpOCOtKBHoJmRe2dDalA3
yQ9FXHLUMNYJwnGLPdUR8d6lGv0gqL7L84nyrBNSfy38wgWgjLIbIMsyLaYosiL7
0yMPIJdfgJnDIvZMBXPWPxvRHq4981f1G1alBKoE6xaECoNYewRTDe0qmBm+f3pu
zT3ESGcSFV2+Iz3DSc4+D0GVrOe5FPsSaIuuJC98++mnzGiyCaTsN0jrF3EXwlqI
0pfCFbC1/7ys7YMr2Jr/XFHDj+Z2mcKg/QR/XKte1PfCvlXmMTgzvYTWSsJq7obN
tg6r2g6K5Td43sqqc5zZ01PJRoo1YcNXIO0TYhxd5UR3pLce1eN+egPKMEHK3/DI
+4UW/yqSYmMpflFIj45SqZSHclmRevqYkYC+/JqJv/ViKNk26hUL7Ej/LNbpI1U8
SCG/qqdxRHkVe1nUyaOvX3bLv92yvePtEzypQIHeLCDEJALTpAFzExtuzYSQeEEU
AmY9hmAt1uq06Ac2UZUogcoIjr1jZEwNSoxrokYQhLVGNFNWP1J2lTlwvBoDGwhJ
fN4D4XAu2p2THiUwMWA9SNiBpOn0Pm2XlONoN3ZQPC6TUnpRQA+PnWa6dqt9t0kK
qPixm7F8ayJwbuaVBh3eAR4RK7Wm3n918jtfZvHNNfSSu2S9/JaawbUEYYglegbd
ml+1d/jDuj6O84D/C/oHz8E3+upivf+eQxMvKTWA9b3q5SlUZq04szTsTkYuqe95
EiBlr7vZ3FsEADccamFeJ1bPhsmXN33jZvU0yAq90i4B5wliBzziOWm64+5bhzfc
NrxhkS9IxPl/kxvZ5RPDCZMd4/tugzezoFgqM16E5Mp0RMsULllz63GgHRWMUT36
IohtWO1spaVbl7vGdFxCeKUVpe00ufePEP4QLW4QW7r34wvEyhSXj9+oE38d+Ip5
CMu2olWvjdAh6JX+7Ld0D7y9RavcFHh4h6IS/hj+aSaIVyKvkJP+RqjjaC5KdJEz
mlkCGPXGVfkwPNb//7/wPIodUWf4uvQvMWJ1T8EqSMm1izCNnz3rH5gNNk8a3gAa
2/x0DUVdGmQiyeQQw0bF1SOqn3Y1517YPE4Nm5VtiRCzIGZKPmPnJL7G/Be0dsZP
MXWhRzJDcRHlrxT0LQBvlNm+cqrCk/Pf6CyIXfLnfGSh/mInQeCxGtd9YfMwgLAS
6kWQUg48v07YPhW/P77883VLKxgkFTwF7M5PHi0kOVjnxr4kPI9knZdrxjvqQ4sB
Hw+QVjmJKMjkAKzv+UVuOC7iuZVwAM+H5AEDY4F34Rw50yyjIi9DJ/4mShc0Ne10
S06bGpFS8j5bQwdNxEdQ9fghFSfAJLsG+qlEWUpOaMEgPpJev2xq7/fGadMwf/lW
MOm4CT2lKZQK/1bylKFDEMgb87yrxRIj0NEkHOyK8hnvf0g8sJ3hNLRJDrl0WqQr
HaFk4KDCormLIKra1RbWa/RbA7WS6Bsf6+Y2k6SVGZg/+DwgbpSK5uiviW1Esuwj
U+y/3x3D6phpXGLydhrV07f7J5kL1USaVzNS3sozJatnQuqneV0Degm3h27gRh8n
QgGKSZGxnrIApvmSwuhvd+fbnroh/CF2Qw06ZGqvKlI4z5aoBoFyv50mXACI2ona
LsJdUNtwXCdEDyBmRA+iwZoTXC8p5F2LbYvfGo6wXgoSplk3Axx+PDJqJRtUFEn9
adtbdX6rqljYIxtMQd1zUBSqclg2TWMF/zzb8u4If6nUa4dCTt78UOiFVFhNLOKw
WZ/O0+sjhRQFrCK5ZWMuEFEbOds+Krj7kgJ1ywXwilNVN52rfzd+NlbOULkaE0z4
OsKWHCMCpCXBj2G/TxcqPFqYdUrlobu8YXoWghLwqMXJ3w+VG7B63wllSf9m20zU
lyljXKh4y+bt3aS6UxltxugskNGyF43EuTtx3A/nAEHkLP+wER0k+q8OT8VBnz2V
hoC8WIUTwfro2pWIOASztBeVI/mzHzAAJjmEWD7zjND7Vqq5uraIWrZ8AnIsg0Gw
lUsstwBxTiZpTLyycrFV8wfA4aXM79Ykd9AHM3fJfeFAjxcULLx3/xxRWh+uAuet
5iTtvLLczoqyN79b6V/v6pt8Trv45f217A7ODLdILSk7vn/WvIbvhHLmF6cGrqz+
Btn2S0hZouuLKyGJVv8xgwbHmz7JX0+msYL2CgbM/iKPJ7g1LDcYuP5yv3YYwiqY
OPWB05cKvm6+uS55PKhueEUjsJ/meSApkHl01qFEN7D2FVV3gOELg/rCEHqotFBq
5EZzcd8d/H/AO1NylQFgv6BeAjUIwIW4H/Z8Hpb31ooy6VWSrfFvP8hzBukRYVRp
V7bYIrA+9VfuEhPtISR2s3jCynCNFGkDaVzjHv31J7jXPuJXLPv/O5LtSRtjXZJ3
7Kw2EX3qdqjEE8YqThtDSHJXaFxILJYeBosXNyI+3ypi5/7RmrOunwiALAKql4AF
GA8JTDmSPdjAwMW0xC/WtHOiGV0IrLQaT5TXWaJudWIhl0ZWP0Z/CHTJF+zKHYnU
KOYZNV4LAA/FPpy16GFBPzVsR0GScvgMs1tj6a993VAogD9EacdZpOv4hefDTswP
aSS/EivdfOjYQIsAQxpOnECxJCQynrwe93JyeAi65ZFjoRPBXQJphD39/w9pRuvy
1IgdHOW6/leR+cE9g7+3KhSR1p+s1eJMmMUyRm99rsbJH5aJPmKOZ8woixVcSXAC
1Dhb3BMRmplwkV8SkP0FvTGOwnUljvpnmL8novUYEWlSCtTr1rJdc5lJpaYt/jTM
GmrCcLFvP/CR1CipjuSYDpthTzVjW+xvBCmEqxAyiXTcNO3a33F4OWBwkuEZ7k6Z
2twSE10KOOXyWhbwdVUuA2DQpiyeywI3/TtVZ9G58Ae+UgdC9GViZXWy6reorJky
zejfH8tieg+lqvdBQX0fyCa+u/fNdDXZdM1TEKMz91gtt7kyGNCcMHb6ymREd+jG
IPpemeFT07mjKBwU+niOr92dOU59hXDbVaSOArEZZeNlKc2/TbEeJqJ+KXiudB/i
kQTwJ4ooZX1XyTFIW++/VC+dmPo53UGJX+OXdjNqljnGZAAd4m5c+PVq3kRqPh1k
kB0e2vOFQZNOa+L2fvHRHjBvg0tWGZpgevGwby16ztSRbY+RrQ1pS4S2yhgEz6jv
RSS56wLCzm4PAelhlScGJZ8mMwCodFezObg9FPySqBWEH0Jm5BwYdm42Stq8axZF
INc0KVh0OicwnwjNd4nlpJE3/WEoODm+k0Mhg+XgBMCjyoufbFkS+rh6ZoaEGYv4
B4+uwQw+A76G4JRVwzZscmlbv8V4uFrHpoeIbobFbPM1Ziu3dQe/PcZFLmfhpBsA
M+X+baK5RY74F2OCIybKYCyJ5ZN8MLR5SnbbT/3vjgcjYESrOtTFz9fFYsJs2GhH
8zDQYB8T/z99z0AY1fH7089MtlKUS3EE3tzfntUUSBMY3FiSNwaME3ihKvYDcOmH
Ft4YBWHVtWG/yG2ykKfiv13pZOY4I3nk9xe8F182FSSczY2AamXGciPzDa5QAZvk
fpsxG5SrsFxtb4VvZ1rwmlp0d2HxHjktjxQbd6Sp80qoT0B7qoQQPZZKiVnLZCHJ
j7u2Xdo3QbcnsBp88CMi8Kc4v2lFqStJb82mdNDFh3uawe/DyuMp2xLC4YAIWSmh
Wmm037uvdj3gTnin0FsooM1SXpmPGBh2w1FxlUcqSUs+1b4807hHcmuLrElwzxdC
COV+FXXD5b9oSGwUtmGy+yV8UxPurNm1VGkWC1CS0Wrf5NbnSJcz1PUShtkRlk0O
9b6FmoiBxq9CsN4dafmSt7Q3pS45MFcreCid/Newumt2dmDu/4SGgGHlHaM0VtVS
bjwvNVOB3YeTAp/pQIpNwfE/2oEMW4CLCDfUfYwpWm3tE6rhFXh+RV8c6biqdDj5
HzaQWSZQi0CGnqN9G0pz45m2TTqoYYr3bz/Pl5zqFJxtoYO5xCrPYNfK8m7mzGh+
cuP5BMbP61pY9Qhd+Q3gTIKfnjNvGo8FDJu9K1p0iZ9ACv/y0FGkQ0C+E02DPfqL
Y0NdxSFe5il4HVM/N9/K2MV98Lev1elhsEe6g2bK4tvq0+IaK1oneRHtVMRb79br
YY0E5fXP0XlROaTLiZ2gX8wfbuJjdK28rxwl3pS30mA6pY5r1INmnqglqFoZfzvE
sZsIh5Ocf2I6HisWmKWCfw9v6j99sSHrUCODk8pVspPMwkq5Fxs3w2Mut0+Gz0ot
TNm8tTWF4l6R/cMAYTQo24F+4kUbsWtNSLVgMNG1SniHHHViR1r4/5AEp2sC3K10
9+f4gE26g2a2OT56WJw4EhS9MwMmdzHQTks7Thaos8IADuDAHp+o7KPiAD+vLC3H
W6KW4vbA+ZXnCsABzO54tptsUPnXIOvoME54PoDplAoBjkcy8CZ0hfibnUB2QeAt
LDjNfrrZ8LxMjK0rJut8aeNT1/j85Y7USwhyrLgIiKTwvxGpr4NmSSy0dPXz5xVe
t0jxv5nnD4c9/PIxEOjP1t/U877WcCc8FJ/jk65gzR+KclTsdstQOixgoEQcz+NU
5wjKoPV//VQVWTgfX7u1Ds6Hw6fRY33uzkgGaUi+DO1xk6IWIaahzbEpyw1VRhKG
yr66VFlTdio4KYzjY/EXiIKJcZ9P3TtKbZTqS4Qss/UdRvVJDhCxgj7k83WyCw2f
0oq37l1bJwG3Z6PLgRTexfJkS//g2bhXJtmss+CNR7GBSxfOUGS8Dxp5K1PRJjJO
zCI4uNT184hjXzbBbgqlCMV0byH4iUJoX2W1ko7EYRIUOeIi4oJqaU74jPuJ4hjc
3M+szHlhrVJpv4cbJIySi1hVv6xVhlmtpHBSDrcLAwone55PKQlCGoGYmDyE8kZm
pYpwfrHI1vFIayStIL4eA2Jz1h5xxQjcdZXZ43mpyacpak7Et4SUDE7K0SAIgBYh
dOZiRFSxMloszMmkCM5yEGBrbs2Rz11FB4tXNql6eagpcIAGwd7H2/aLMoTRJtT3
PkNFMiYC1VEwE+VqXa/Z11pyrKaIDGJhtdd3s+I5jXwVaVk1WEfR2TgIaLwup6VQ
2qMdJ9ImlrgkvcotOtHvAv6JPVkjugyntXZl3w9VEob9Hdv316WquERALUfXlYem
PmQgaoXc93fZlOTpw7A/7Z9OV7EmK8rN40+rcfthrDEXeDVViveo7l37rU6ktZZ3
cfpxGMvgOE6cSyCiuBb8PxT8FjxqNaljxv+tWmcWdOhUp0RvTyMWUe/wb04Ht76L
C9+4cR3gtChqqQkW2PVWi/f22yozF3rooZUnoKGqWvdl3DRTVcmDltPwKs0qTaHy
Te+3RwYdGIk/WOFxtHpLtrpG8vo6QVI4AcfkpTmFzpKW1N22HensGEoi/0Nihm9q
8Z2Hulo3lruyUVVjYoPJWYJ/MplaUIQeCgxa09wvqJGGmqsiEiZduWeqN+YvU1dI
13bz28NriYZjUt0cx+wcoPage3ss5cTpW3TC9/KiOgMd23/xR6KAajE+O5ZzxeWG
bKkoyPkEoIzqwWVCCoQjzRL8OhLHiaw5Xza9dPUoXysI8kehGjoyXErSjf7dFB3A
EPdNSfhyFbMllJtBxXbTgZyeXkUa9M2UGyYsleFnrHzXygx1T+jwhKZUrWwPXvau
//N4LNi0gTWeOw4d98k3BoasyZHGAgCYYs8HOmquqIqt1qrGsDLIDTD9P9I+ZkvB
c5l3jVzkldQ/8AT0hPsawwi3rKUvhlNaaW85mYRItOxY+SItpTC5kpV1qlbEPnQc
TIStOBRhOZ6rc2R2ux1EHS2U2Qh8V00MUH2LghSwHSf6lWW0x0EM8we6Ho4t+Rjp
Q86Su2DwiISphSRq5u8f4pIKuzhRJ8qdN/TKwQlwic7KRVexGHA009OlJIekB/yR
VPnd3mOgBWD6Qn+dOGkjKWEC+qZSvB8V24TTo5DGNBXFhMXp6vhZV7Y0hJdMQbI7
mqOnTPxyRRAWqZSBe1ARmhQdJ9wmIZ4/B7Kb59QPM5fhGJNNkDiqioG9fCduDLGz
GVrfBH6+FLacMp4ZTtzTR4keB+RWN8/9iwh/y66y5uh7KuVKLt5IbB0NlOL084UC
liVll6Mgp7kC8BPAZsFnmoHcpB9wwFb2avbhMzUXaV2HuIh39RdHtv0S94iFFn4B
1OGEp5CykkKZYeWbmQXCsrwb8A3qBSE31l8QdEA4dgxo7efsgQvqDp2r10rmLFQs
P9V3g2DW92UzQ1rnXZGjBp+LczC16VvhgDlWE7EDqIeM52Ig1MWx9uZzGQEMETKe
F1goXKNjzQpY2qKWMXyssnVSL3BLfIRqnv9+/tj5cwDSWQVajftpVdET3D8Mr/es
DHTIBKhC54kRIOe9VPyLJ2azviiwN5Dww/RxPH5SDhCSth2oAj9ZeMDr8h88Zz3J
mhCLfdKPfl0YvqM4iqJO31GIc2ahBA9W7+NYQG0NsbQDqGUkThraGcAnq2hkfA75
7AlrqIN7NwtApqz+2vNrWxow67ct3+6IGxcN3CS1bQl8SIVNEzSfuTewPUe1kPqP
vyu8RRVgArx9m+k7K+KroHGYk3JkjVDmkcutBuuqcJEmeETR5vFg7Sk/Sd1J4dWV
gZAPi3GArY62EsTOKmOE203vQWVR6caodec88RDqBSq6u0G8wnluge77RUySyQpJ
VOshz0dtgfbXXc2AvsOEjiCBba0NL7c1t/7anmSmOK7FItvcD+41iRuG8UT4H2A4
AkIDL85tMC6q6kvjlGuu/dFAnLNd7KAExmtY7HCnfBVJ/j4lnNcKakLv56v4gTUa
E1iFh2i3jBKYZA3zmjXkVDyQRvtVCvjqMsmWQl+7y7KlAFa3GJJd+4OW9idaaIxw
OmcUZ+NHQRZk3q/rN3kFHTC2C7skF/kKW7Fl5Y1NPl2czOyORR9wLv77KlG1XRCY
PEt96qfqnRNLxpedhcNnn32Su66/K0WSR2yoaGcwJ0l+60hC7QM30FItvsXgmnLf
nQgjL1B/nZvHYkzZTsI78Av6BP3CxHG0ut6VToWgZTbw5/mAIXtCgHl5WG9toHmS
2OIdQRhaQJhsICzP6VRx990hNivLbrRDlX+7V5tIYoEJgdlWvQko293dxGe+xi40
qd2HO9DLgFJfxCaziHQKB+nsJsMbxHrD8uoYdt5Q52wJPE/MyCtAI9W7BRp5ohz6
Y8XNmzmb/hZHmOY6zAb5F8ymLUEE63xpfiDN+62Iavya7S9PBbI0o6SNjBAe2cdT
WoblvOq6iee1c5ph+5c8kot89UXxziyVxw+baSzxfnp+tS7mRBHBrxDAOq0YYjw7
B8I5nU0qCpXOe2WZxA4j3pIJpiN9Cd9P8Uvi+3Vu1lRE9eoEY9HJfOuhi9Wegz5O
i83v4HRP5Yk8qsSgWpy9dDsXrD6frGRByjwOgsI6nkvJhVSOEZ1P1nGEd8JMjtpH
SlkQAnJJ9JY7AqjFWWUjW0fEcM/0mCHa9930aSFLcebZ5MGUtVW5HgePHKOl3cAE
S/oWr1sEvRzo5UNdyB01VF5UqDAviRxKdAllNgO1GhOM9NFLoiztB4emW3XeTgDL
2MggIAY7Duhg1Iid4Bkgtf5pDYEpZqIYA7VLvIZaMBNkD3Sp6pKbqB4ziE7YKwQc
tTOLkFyLFh1TJoZ3ChlvpXCbpDYh0id02O7PwbOpele+BVSpI/qDmRnrimm+h/s/
eStGGvcahwY//Je25+CI6DJdPwJtc8i8+lW2175xLK9e6w42A0ZZaPWpylV/q9Ly
Ashug6nVsEnWorM03avNRH0x4NspV1iqilsFSp0P4cIlqEiNfrO2oV2zZiNEyuS0
JCjkv+hZSiiOxXdbcCiBC30ePJlVzCKtxaw4XP73QNsqqpvD770SzuJyL+yuNtJq
DotuHuVBcLNWiu/G41f/yK9RrVhJhFQ4j4AtcWHBRruE9L+Sb7+KsUGSyCZai4kX
WxdNGfHTbHmpHHc43B0p7d9uyIFPvDJb1SC2evWU0syyKim9p0/Dm5BbmcPsdUug
RRt6rD7J1BnfXYrq4gOZGcQrc5Dylfuas/mrrxNpHVOBZmQRwpNPoyWk759b25wQ
Zt2Ay6YekyoUGvmcveHha3xJvLhidTmnLYc+RkNuWS5NM5K0C8SVFcdAh0ep/wwU
JLseWzXPQfENkaRa36V2vpK/WxNs3lB20gDc8x7mLgeUhTwjerx9pTmbRMJeB/70
jJDiIUQwB3fsOETdKNlT0lI2YRdsu4DFW0Wa+xQLlp77Dvi82yHcp1wRVuxs0q1v
Ns4cXxXiyetcNIOFbhXRnMnR9Wdt1MM5+tjqFKYfXoE5wHweeGAqyCd+WigNDXq9
OYt9yfPJtHbz4Fa9g5GfMZAsXuubpWpBvgXoKijLlDgEbyg2RM/VLW3OG/hrguFH
x+zHkFwMAy4T5eky3M8WKBPlOcKLZ6zeMm2fDaMIy7NSVzlHVnbGNSEy6pP9z5nP
S4+ZeIlXrFi7HYXNC51LFPpHdilNd0nw0LHfJGQMBaJFfk6KoNwLcCe7JiOz9EfI
0VJaGwpy0uSymWhRg4Eqy/t2gDOp3wNqYNpFa9QBRUOwf3j4vOLSVHTSDrXpz6l3
09D2hd7f2rSWeWBa/a75SHCeyfyF7pzqM629u6QHoMK1QNvb5yTJfuCjDh/414Rz
BCHqHlFXbHhjfd2GYkhN2Tljl9erY7YcMjDE44/G3m+6lRoPlThPDc34k5rBW3Tv
QtN8rWileH03yhFx49fAGQyEv28nel6SBL8taCX5LmZwsZxcaSBHkjXHxxViJYmg
te0NSKKFwwtgGF822bhvyOVaECd9HRSGNz4gn5SDZzjvgTTnW5ZknEs/mXbmhJpM
Oe4cmb8oXtBl9QLuyHFzdPXyyXeV1+VNTQxCbq3le3AkT9P48U2SiUuterIWhtG1
vrzOW0oJfYpCXdGS5Ec8F8VdGSKegZq/LIZUYFfLCEkwCWjxDJj63VdCt/Z9E8uI
w3T+eMP6s6OTsCCFqoZOZxOPURq6jJ9In6NyCy8wIRJcctBWJ5sy07nmcd3PI3xo
znLYtUtnsHa9FaEFLdBAuIJYECQwUD9eD+/mrV3FqguKkCzmpvndcu2O7jmZBJqP
Da3r8kAyj65YHKmdKjHEZ8RZtKhyhhWKPcCn5gb05y69RCp1ciasqXTBYqTnSq4W
Xz/jFahktEcIKO7dqBI3vYA0KpZiiygw9EwlhxdeDGGg4ITC6I9Xa355ML6nFKGY
v9XHRM2+C+/3lJi5WU2pOue9j7/H/k37lbhfxvNvpMLeIllAdTzevOJJTe7Vz2iB
aY7M5gM0h1wyHevZ0iaecbhTaRWbZZw8FwWZ3uRHvi/JKZtzWnlfLN9cOPGWI0O1
Dde5MMKTJq2lRqBeBfmYX/6vjTp53u/E5rW7dqnljxBEYdD5g4QY8/d6HaLxxVsq
lFccBYHsssUMaMJyplO7sUZiSAXBDz0zQL4PQMzi3/4L/AcM1UMlK3MsvejOBapd
0qHxpuMwo6r/rRw/QajZfzGqri1eNqPof8VFmVmw4x13amybE6BwAr3O4p0JQ/Pc
X4wIJGc+jonEVUuuY5EVvVSTkBAa0k4z+2BE5BnazrgQPxo4WY8RUoieqdx01Inh
zcmQJ4LEqJCTo2pJwS/QJDQ2NF5nWQqZlqhkNdAWWvuc8dJICt4+odMyQcICBN1A
/alON/718LPw/pHq0Fhscduf9kS9y4ZeaQ9QsRdkT1d/5JdsEz2lmA/lkLeXjCTe
W5AI9yjADpOq8L2/BbZNfoxXO0YhraGIfLms9t+fRXLovErgFspJAsCU6D+L7s/R
NaMamxm9eIQKwn6os5AKKXY9jKeWUcM/Hszs01d+G8P8wPTppa/2b44szylEmAGq
k82289xAJry3HV7yL09eyM5iLa8LcUZ3mtVX7f55RYin1aVgXVd6cqfRHCuljo+W
pGYNBQURIYozt/Rh/5zW42+Z+ucgiJObO1lVIlSaz1gF+G2Hv2o1VpksxPgcqDrH
U8U4YEWbJYXJD0VwqUz6Sz+6dwiGLCr+BB4X7r+1vb99Jc85Wm+cBieR/Em8ohCz
8N1PatIKXTIRHL36YAQvPV42EeLpUPIIvZk4iKcb9ccUVfHXkZXJqChMeWz91ysp
elsee56GPdpHPKaXIdjnefKDjt+BFAPOVUgIvN//rOU5HzvJ/wvoSI6z4vnhe2nh
OXY2CLqR5Hv8Hs2hHf2biu2EQpE1Cxl4gU0Ec1HNjrqHaYAyTTfHActR0bKxrVsk
Bc3TACN6RmZ6bIC6yST412cfbYwV+CYGyKkUmaOVMbUnlYrqn5fy3FtfgmLkZ3Er
rSPJaNWSvCtZ7F07zXchz8BWPW7XEBaGvFNQtNnyhAO+Ul9QXd5hbCIv3DDpZrnf
I1/L2VBtFsynbZSaHipb6vO/8iVcCXFhgblJTrbbGOEyKl9bRQ5h+CndpXoupfsn
eHDNVG4PIHuP8D55KhC8wlLPXT6S7aX2pexj7dXAcBu8jIlP6WW0DIv7SxFO4JYx
ME4qhP94061nBqLsNljsUhukJRaf+1iUBT8H/SJU5+nGFDNaZI8yNOg9HBVX9ktU
kgbv+Dz8RWm5avQyQj7J2fMy0eSgroNET//ZNajCNjeCfUzgRpd4l6vOyaZPo3JX
gXo0jyqpwy3UdHusFOjZtQi6Vg5aA93WQGFkMy3z6zJ3COwbVG4eMj7mJHLn1bR2
C3IGRqB0GENNsFAyWFUkRLJThya7mDRWmJFhZmKVzSn2NLMh+TZ4CFTvKC2ckMmc
4t0lmag/qSzIbdx3qM8K3V5/vu9I18S0AEL6uDzXuAE9pj2hOUMc0wXrqFcwPj8W
Nwag7Egko5fr3ppE2eKp4ZqUuUJRtO2cHaHi+5IXWOhrVzZFjEn2EZYG12zeEIjn
0yJS4C4xvwxb/jsuKZI65IBTkuSOoR1qw44dr6gUM45S1kjHolN64zde+9fuaTcI
34zUB0p10OVV/WwfsJQYc9hVqaoyXrl/AaKIu8u4RtNzVQjYUPe5uDnNB1xC0+NO
Ha7uxwdZCoi2yqW1rROixIOArolBCI3W5J6N669LBU6PVUhuVlJOtV9Zfsdb/TFJ
CuVhHKREcRIbUvjiR2HPa0mgvwdzN3iAoMGCWwdznZHaL9wVa9Q8Bzpvq/drNF4t
/Hiva3Gf8IbDaoaLNBDfIhGn8mqxKkwI2LSvKs8tbc/5li5wdmAgyeUxa9V/Vglx
Y0wUXavJDlgLKmCNUYNLnojFu7gbXgepOxNjGvgJDMHJXStzSi2snWFHOpujiFxz
CLBs7rxEFdb5LpjIOM1+Z1A/TGyY8gEvAf8kctI62M3nQBN/l7oi+HMQK+jFdJd5
97EbxZqsw+v8fUWi1jXbXvUnCLnWk2qHgqLbLLnco8rZq9kjMAXstayxX10COPTj
DU2ydAq2HDczLGL3WCFPH+whnE5K2y2tPZ8uIeLoRR2b9zz0+d0u1CqOL55Y0fOt
i2sCboesQ1RV9WCMXk0VVeJZ03Xh9KWMdzCAXr+zIVdMRsmy8pQfWV91xRKUHve8
r5G2hDVHN99wFb74Oj8AP40A8aQjlqOq+JBBNb/kSeA7CXYcGibVt6t3WVFJcLuC
Fc44VB4eGE3L2ZlmfCSWFmHfmChH+F8EsFu1dfl3GZd/bx31PkSyu8NqnZQ31w9d
vR/iSpFpyAP+OfEc618tYvpw1dyyNKZxqPQPu9oLGaNL4aQY8djrnchvg4BG/wX3
L0/T8NfZT7dPzxsRtlyanSS5huNwU5v1JLMgusW0VuoLi8rF2bSTR4mX7nanWYSw
Ihm8hyhxksZv6n+pTMyPumInK8ve3bc+grxlxVAnCzWkJU9QD/aVExjiTqw3pQPK
06unXTEoHUcMKP7qXP5ERriyVLPCzAowKtmauv4NIV/1KeWGbHJLjuFCjh7GPVol
Roz9W26mlEtr0XDm+Zlu7J9Ittrr5HIBe2La9sNiIwXrxG1dsgktOO+wp8sCp1JM
oKcbSjKRvGbtAR7ByiAyx4Eu/qzp03fN+10L77O5uCfRJnk6qcVkz911Xk2ngd01
J6tienxTWXYKgJM1twaVdrNyOZ22H5DSjOdtKMfzCNJoKLNaKBTSCOKysf4IS0p+
c7K+7O9CWWYnbhTbQi4FSbA45pJMR9xJah6jFeCPCKgJ+QflBjXwUcdPtUSYTP+Y
C+3g2G8dtIhi/GFs7q54XCLMsuFLES6y4yAG2ypbCGErxTLQnWSuW/YAQ1m0pSIs
SDXioKTB1i9+8brWalLUAdI2ITZoaU5EpjWN1oRZQZG6WYphMzv/E2zV7qdjlAX2
MxkIKXOk/qZkNwu0ntzqyto6XMBXhWT/UJedZPOHIvpruAiUZT5ASIGg2WCpboYY
gEUqv+hoOAL/ON91/sRR/r+mWjh9FY0+OAR9/lxs+9ldM0MwBa0W+0QRAYLlvj9K
7JYtCOQM1ybSzHt80QvnH0n2uiIqu38SX9V2Crs1VsQ5wqpfV/NiALpVS2voKS2J
l3AcwxuPG579/ZlomZfuvG+uK+FF7YIKUrUARO1qwL0cT/gEq47pbiOb+mtNLZJ/
7RMDx9jsCebYgP/XgZDr07FG1XnkM7YWR32yNrlI3xnOxxr3YywI24is4Sin05HY
mEkWyj882YTaT1FwFhX3vgXotOlqu6dHEQwdqVMTWcLIvFrQuhLR7qgMAMjMXJEC
28DjrxhmvJcFOzfdWiP+bzKI5of1qM30VIMSCgZ5JanBr7MTKaXZpHDKEQaAG5CW
Bolb7TFpDaeukJ+8NTrSRUiqiVlUj94iWC9pfwrToBtx/ILku4otFDuuq92SUOuy
U0LYlvrB93p4RLGXqVCJm+zLGuvAwFzCnoq6xnVsrUsjU73xBskioPiAAVcQsS4P
GFxde7XP3UEdeYgQoyjJHvu0AtmfdY2C2GQ4YcIqmJj6GaXjhQg7xi66x/WC3Wm/
++TCrxjiCN8DyLK+zJtgRT1o1EiY+61GBJ6zC7lUpL2KirKxijiyC4E0C9FesS7L
/HhMr7VghD+uSWr8noh6TvKfKB/gpR7mwm2h0GeU9HUfFyrHWXhDhD+ArPk+cs5t
caYDkSSVKhOXzH5SDCDf3ayLopHCDh0SHyTaa9L3jQ86e5eRK2avk+TOKTFpxDUV
sEJ7mHAEbHZ3lusIHVWBfzaBQEUMlm1qO5NF4h8HdxuOqKhxLFvLsinxvwVfG6vl
3AvBPuF614FBv8V+WaVMtFFmBJ/rasKs70BDl/tl4qOoWrJ683XU1gawAga9kVNu
ebaee9RQ6kSWN+OzNxP1FFLpe1153yhr1j9SpKooKHc0CQCa5qfGNyIdwTkdO/nZ
MMRKnSRKT9wpP+s03nBa2SaqUBwjw5zJaJd2txP3vDk227ei2irOD3FcC7TV/e4X
t/zsddYWdtBrEiV1EAdOYll2Iahemg5LoFpbbCkkYmUPFqazFaQX6i7BgXcuv1re
mtg0SVQR1Vmq+CP7Xkfne+Hcqmc8ETZhhuzFVo3TgSokncVId0AmhKnGLF2mKgxZ
xLHNz19hfvdfEbVC9VPG0+Q16MHCh+hLXp9TwKX4cHle2ZsKc0tB+fzQ45oZPVgs
psB5T7MXPM4zQ65Vjqs/1+RUvBkU93ElXBNmOVpfcgc4gsiVfcnojWs+Tq6v7kMI
cOjR6rCMSFpJLQWxCLzT8mu/Lw0Nzke8ktVr0wxMJlQWgdsm/TNy5tDEJUzCXMSm
uH4pMwvlXoXzSlUPGzKA+LSkix9aTr6VPSHeMRfg73x2cYvuyW5WjHuadK8yLIw6
3T/ahqXAXLLepJgrm2VBfuBJjjldCgLQ8jCKbsYaIzasPBQwboMyDtu6mbU4f5MK
1tb0sNociD6X/P66UGpyUkiBtarXfw5GWPrSu0xA1Pg2y+1tYE3ZX8Y/kRNQnv6D
mb2sAP37OQRjTvpcqocUQeggoP6VAsBxznA9UDg1uewkUtXwxUh4FhfZkmZ3YuDL
shh6Qto4lzhsxy5vIYqEVKCjW/sA+pjKAn0u5ZFmxfm5LaunKsph0Vx3TcU+S4Se
03eOLT5bn5+3EwtWdfchIByOq1T8AoJwEdCZu5TOG0mFWm6vGWJx2IV7cO32Eq0d
KNBnqqqQU+m47MXN8GFHQP7hm5GqcaBRd4DTlQDN2c1UT4326YBiKFnb1lIroc/W
Cd0pfE7EMy/lcZyN9e+eJF45qOKa/tEN9HqemORJqZTm8CqAGUPs5ndhl6J/xwjL
2AFz+rhXq8lvwAnWK0G6wzV1GpcbOugIeHYeoG2fH/VqzBqpv98/eDYbF1iTT86f
m1vQ6Nt8HyWBYSP7p9OygiWNXjMbIDkvT5MYeWoGFWvShM/pqQJXxaeoXI3ZS2oS
WE/tMNXK13p23sy+wqn6fLhQdHhw6REDQawsqGExMEPBRXXX9rKtt2Ntdatu6zFz
j6HaFmI4ZIf5ifWeWWb1NPdZtBajvPUJK8ZnayQm49HzSlT1Fplj1qo8p5TIhiuz
893R0LaRGK5uXY0VQQxTHq2bg63PkMHnQdH2xF9xXxMjA2Hzkpnoe9cFGIVjouVV
GNoiCBTWqq4JsXUj6ZI9uYU9DsohXA393rurqYpHnD006lF2v/ZAbzn/8Nbm2p1B
YvPBQV5HxIQpmhDW1KwuvM87R+uXmZTnMzEPFlwAEBDiR8sqnyeeXdPdyB9ZLlpO
x2dkNxM8lCLHAnbx74BbYH2ek2sHjDv04XEbkYvq79KRsLta2MsviooNFC+LKv3K
8RYGquIeT6EXpf+boS2lx5sgvJsNCTS/axbK7Gmi/lbl/UdtaVKBJ2SRxfWACGAO
1+oRPu1/OnnC2bTkH9K2r7FZ1KLIr1GwSgCe40xByY780YhHL1dquqjDvFNZ16UG
hYNZCfNkOQxWW2RqZ36GF+oJuZySDwvkpwOBDL4Uz5iFZRvVuNCeyvktkMeiteXG
gWPJO+95efROiwWlLMu/ko6it+P9L6yieFa1SiY+l0A4wCdsp9dn6NDkQjXLkhKV
Tu3GW+AuMVWyE3agedDr5+wnxwstgUc5i7uzRoDwA3wgNw8LX70/I729W++U6mAa
yI1JWdAwcHn55ctIq1Cj0bwQvAZhqnLbd0Xq7d+0FsB3SmYppoUDJ/SixAnlA4xK
jsEZCSknF5Vicerych93lz5We+MTLTxKtxf10reclFsZXszhLOAtPytndHRiAa0J
I/loCvL0BgETHgKWDVumbxuGhO1ZDWTvHq+92yf/NCpHs8YGlG10Wmrx96wF47XE
lJGbpeFx8kOTj0a+WlUoZhnrhmakzJSXzRoIADa7MG+hAv9fnFFxpGH9nn5kI1jm
7NamkbgGb9Vbjr7QFmMN3Oy67larTLpEWZ26W3Gsvcw8B5r+cy+BmOedbw5xz4oZ
1T/Jsd+5VQaVlJwT+dC2a6fdouuhkSTBJrcjT8QPA9Fmo94GBPgKUTKb3E/28w7K
X0tWWBDGOiTAGocPI7Q860dXhs7fXsdL+jcvpNkHIVk3X+RFYLs7SxK6XwH23Pcm
Y5nt/9bDSbRUxMur+P/+rSV1pzzWbVtgEJv0MUEYKJa/1gP4RUF94Gi8jUkH/cbq
6GCun6dCwF3juIhNnpqnXeEuotByE9RbbquAgyOn4WZppundyk/Xq9en+vMk0QLU
Qg5oHJWgUKSpYgsd8p17nnhLKQS9doKWqTFrqhZ7eMCJkz188tgDnp0c4rgJ/K/a
ycDLfR2vhIjtSffcGfuSUYwjJNYhpZqYsGbsBELRl/GOIDXtu46wcM/7nf0Ck4rt
x11jyMyaMci2LV4XHVnDugW0nhetEhxxD1LKdLSnFAC3lCtDv149B+f/9J7gnTMW
u8VIUFfoJhjRYlCms8EgzkDV9EuGbZrrGhZ+6UXhnCMg8pgMdH8j17N2RsrlDQYL
qMVuDQmqBMBIJ/V+HShpbk6SnzfNhSXhtNF0qIGZ91loGXvl5S/W8t9C8WM/OqzT
ofFzs4GusuiEaaTYyENeeABjEkbPoW6Fqlm8DXHEgdoRIJa8m3BBKvSCDGKKAKSY
iWVkqQdSpTpi9FrHB6PD3RcXin4xgqbTMEd93OOL9nAUoTjCCEljcyhfPEo1RigZ
cjpU9YAAKxltaAP9LF8dBXfP3zlixgGF8uYb1HbqsztMFwRbkW4JS7UguOF8Cs0k
bjoBJ2jaemH3vrx0JJ0bV5IwHZNv691jmWTKLMkLto4/9MuOx8iYzMRRYNgHnBEg
ujZzn6P6CvFGG1ndmUwxQaaaeeb6icy711FoKWWInF6MMuyNPXaA3XsOV01Wuhuk
UOlZUTtfBsZ8YcyrhDhM5Xwjtuj+O09GS0Mai9cY71BXQ+BwITgaDoRy8l6buuO6
Vc1LY4MM2htZdeDMO3vs2pP6WT2Hs08/1YZ9nQCsfsu3XrRwmVhnCxO5EOTJvzm8
uY4gtJ9mlIcb3ZOZEScpi7V7J8yKHX1UeTIK8vwW/TCplVBE3VdNM05lLA/bUAR2
o9+iRjd6pBS2PwBWl3EfdNrP5Arak1ZfAssdHPWAJ/QIv3r8yZVOq319elxCirza
BqF/czvWMQxHcSQddb0xu63OJLB9zUsdRJd+2p0X8wEPXpylhnbruqWONdRtzIu6
S//eWI16goCzI+iRqgNs+5RMncTed3mn2Y8omrnvGBVjlimhlY3sL3XFtIyAevdT
Anp9WTqVYquA2NWYKcnUhRu5LYhsLaSIJAJZwBtV2lk1HXydRCoFGX1JZ3zAruZF
aAa6RxeE4FPW8Ro/fR6XX3F7oCus9zpiWPw/hSa9/LS18A4sMSNmeoJcHVbPQfhp
JbBCFWIhyNeOvUBuqHLaq3o59ccpUhR/NuVmVp7tOrX/ybHpWtLUll7QWfBRDhLm
fLZGne4YnhMNJVji7P9ZICkWzIbUy/FpU5VmE2Wbq3k71UU3xiOHJqSkI3r4fuKn
XVEv0iXy8tU4SJTlMa7LyYnWNy4sCTHz4SMFHHs1Gjpzvs/w5HM3fCgA2WC3c9Mc
g3kA00FQNwxte9HbQoXnR/Ay8OT81GZqAZBzJK+L3XEucX4BjxzO3ZV4cj0gU8gk
p/2JUMZuozVxY24gyZNKg/NuCXDwFGXXvqVIFj3B3ceJTtkM7QR8o0onHqJWKC1O
ZdyEqwutaX20V3wiSgVOsFH0NKsgmJovOnU0HPeFSkAibXMZo2LR+QvXxuTwx2y9
wvVdgcI4iZweQgb0CSOY54S3qGDD2BWX1+c0jPC+9/py+RoI2htbo1uGfxp28Zhz
jvoq+e86EVbfLKD2J85EDODwrBuAmqaXk9WdCY9K0MveJQaww62S2umlF55wWbb5
x3zGcxJ449t4zI+LWD9VUUzcdCBSwlQsT4K19HHL7SAv4Qy8Z6s5RKLUPdvUn/v+
pRm8udlsiF1Ra7I3u3BppU7Qk1C5TrTHR3uv6dQggIwSLecgElWLLugQhc1CzuXQ
EdargzfdTfT6xemddlYI2SWXh6MCN+czliG4H3kILisKvpeF62oSXSnFa8Sa5uKs
sT+VKGMLXAmJUG+PFlG+LOXEksQ6G74+AdDpB7PMULyMagYk3241PYoGNBt1riCq
r/ZZnwR2c6zsjj7dCEbYK+YWxbqr6n6E5GJ8c6wkZkv7TASAemgoApxOyTt/BHfy
u3nu+54pwEyWu7UMD9t8Trh7ppqFta5en6Cqhj7R1rREA9Ep3zCghpTtfkzwOvSM
RMpfoMHwovZ99b0+5FOP/wvR1WkQUV9WLb5+ZXLt8FTukrEHgOvYj3smPSwZrPL9
AUJOO/tWLsETcYuJtAdU7k7pdPd0+B6HsUb5bMTBABIaN8m027/RxLsJ0CRowwAt
DbH+YNIiwcDV77sDr+ypV1/sPipECbItHgISnZSp/+yqpOl5MpMnbcCactQQTdr5
ARhjcDloWxnu8KAoU4fbOjjV4vFXVdwzmIHuTxNGEwZ6ZkYIvMU8DfnERn4Fmh1x
7l/fF6t/VLv+Zn8R12YJTmxt+4MrG9zBif2rLZ1tqr9xsALTfIdubE6iO6j+Jq/a
KNlr5MvHVlhXGQeB32DjBGsPS1jvlIgOdOYSljKP64MdrnUqZbly8g29PKGtwddj
SjNhYgLqAQaNgEuKkqsyntiZD8LcGW6avSUFfgjwz4tEsc+2Wzeet0FMhap+N6oX
krIYe+4A/OuefCLyznXUpM4VB91iCRmF8b4od70O3+rOvRjVRiBE3ZRSgH5SyUKT
uykmI+N8w2LXvPaYjuPSt80M7YcYFe+2FOHjjbI7qaYHU+FUhcbQo2z0xTLulkiY
2cTdL3X9XLlyxQ/rmWZ6GWjnxiBcOjLNoXnPzAbMlJ/AtwLMZRZxUZRW0OzCWsCW
GbeQ1Yw31UB5MEpfvBdnI7KxgNzC0U/iHKx9Y+TP2TuYk9W53SDFbYT70NSCR72K
t2e1g9Ey9mJe5ionj+pQZjh4mXWhXMC0aQR2HZAxyFShMFuyBMGX07RhcUpCFQdT
BVi5ezBzeUn5XQ2UsIUPzO7Ev7QPWlMJmm7EPb2LKKIbvMRg2oL6ZK+0oJYhznhW
niZ2oDoORBjB3aXRP2lTUYBfxd3Qa6rHi7+2TkdKD+0VRFoQ1vo19rtsg2muFY++
wUhTV/SQjJcyjiFwtziKiZARslCro9ubLpEI8uahTC5OpYJTwGXXhmsqMo56sFe0
Xbz769nQxwiO3gMbuUHoSIAQzfxnpqFtuIYO2J8/quKNcNufz/k38wN/VqTUBJNh
jd5o1cQzY5UsvCGlJFngj+vGIqt/igaYVYUFov0o0FFdjwXR6r8AIdjRyA6W2sOV
uGMDks4dr31oFG0RC7VQBPc7j+ZKnuJ/iWrPMDK+mOFz3nmfNwmSR/iYpD8VZ6cm
L2PuFvsjRvgyG3xdYF7Et1SaAtGl5RG3/MDByHCCsa7DTR2M6eOz9F+3IWyi2Ww+
YCBEH6Df0PD0+G1ti+LIlgPDyYEPgxaJyELH2HADwDCC5iXrUY+eiMnDMpZqWWvy
UzJ2f3OpWJ1LlqDc0+yxl8FFzF4ObTswesge5csJNBIVJq/CrmMkTu2os9TAfjHY
WYF8+Rzx8qVfi1DhfyZdL4IgnH8qWBerkQhdfusL0SYL3vkHi0hfLHR02qg/rkvi
H+VitIqoKXvB5hMDXuBym99sK4rm/1iuCD85V//7rjOnlZAODjeml04pLcCoKdrg
dXmVeQp+G1K4so4uVDV0jxomzQJS6wtK1QyLl0v4hyzBGUlaEmdowxYallRWeVfs
tP9k57t627vTmHhoQN5OfeWPvd1mV2LApTjv+AvHVg9myyq7ALo40sL4wdcxk/73
jieg5eobb0ImlAyjQ2qeQcQaJyGP9pdYbiQL3nWNJr/ELfOtZtnG7sQ6Qz+W5Zo+
ZVOZMkO3yQaVf89IdBkc6WDZxanvAbtMmkgvnl81r5Fna8sP8iXQYxGknW4HcoQ+
mJtYsXWsthymhODkaN1WbN3bgkPYhWRjpbmm9TxxOe/LwYLf0EcSP0dlZw7IwUgY
RtSR5/U/O/oJZQ+/TCNFUgU3UMWtWXR+OFbKemjlSZN9w/wt8wRa2FYzOaN74Yva
cA9oxp8dTKwZiwGVJBc4rWmJxRA0VjGHwTG+dMDKLyaRdGv0osc4D5RephCamvVr
2TGuGXIy8k6h9O4BfTZm9MWfHzwALCZ7mXvqTqtiZpfK6eP2uBcqXHUcfYg0DMLH
bO4sQ2OiVDAAfX3A4OCW37l7PpCSzRtVNIBVSz5/4RcchhOWmJoRjvDCQz22he+O
DRFfxTZ7rrNMMMcTUk3GqZbdIj+zKyLmR1v0jdJu8q/nfpcSIPyh6w3XhwwpLX9z
UBxwQz9dksEjvvz2pRg4T2SQ70l9pOGga8tKd8Xw2geRRgPTvtWDRvsMfIm8emO8
K/dC3u8n+uUWcsMKbszLFZhYuyOgW6pCy1h/qYFNjFSvpUBsWeicLb6WmBX9YiDk
PwRL8uSPRFUdfmYxAzViJMgXE9NPpGtI9Kg1eT0Z5isaeCE6xtMwDs29x3jFnMeo
YFh+PFp9VH6TDh7xlUbxHF9jfKqmIw1WTKbUChKTOgoAV8qEkZcmMvuAnSiMAE+z
RdNheMzqJQgIjE0rvdEIig5DS1am0HzunJANqRSUJCNEA4GKVHPRD5XdAXnMbKtC
hWmPQhuRrs16rSmHLHN6B0Fe9IS+6kKmn9NxB64KKqyc/rUuYRWirBWWrTGqdKjA
attaRT5WaGSVHyrB7l3DysiKtNupp1N6ahTkHAiYgyMD192TlRfcNja0t8Mei/08
cuZPyj41JElVG31fX3ZEzwa1c60NYDVeioA/sFyuQGYsRW/ZcFeiN5JVlmER+BHA
aFzRHa0iQSXRIdT+HXx4UAKUvBIzEb06R+USqypFAEBjfuhuQfeZ4AtSKIRFxc8p
lg7WEvVimmnw/5dZbjl2n7uSqANUqDD2mzmm0cWKNZMpG4S8jR21RDKDtcpeKVCK
QgDWoYrnq84BpLlq30kKOV5pJgmHibq4Mwx5mYDsIkXgLhvk8Gogc+D5He7xGrnt
+jpMAtCJe5L7NhNWp+SUTj78xeean078r24useHRN9lUkFgRHZJQIx5EDAT6YCNv
j1vV5BNEvCVxtN/wf5GNmIXH95W8JgnHj9WzsOjDvF3D4a9Hg3aXUsjVrVxfvG46
2A6jYsTTThBbJDFfq0UHeTtjLlmxpVyJ688ZrmnG4yoho2c/I9nAfJ5elktUds1L
VOKTfxQATkf7sD+AELGR2zAcH53LugG64UwDzG3WHSnepnkqAGPHuM/55ggku882
t94Wcg/cFhYwbKZeqvo7ctZhfUmcJ0e61oWmlKOH46DYAXYoWjt9WkQ9D94WyyZI
dCviIdBLwWisKRahAL3xw463rC/7lhNLF9KlWZl85sI9UDUyfL9Ou6Xmq30vwanI
2xsR6+1kKSC9poQs54h0z/nicLjv28P3IwiEJUcAKV1CrOuSD8QkduusWk494HSE
dNsnQFHrFUei+rTILCfBtKzvQxHQ0y327xK+spbSyd5Cuvgoaw/sUfWolw+fQjGS
O+m3asELBR3n0qMqNERRhGGsd7ZIzgMcZHVRqM+AODmXbCx4CeHMi1zXEUPg7zH/
cXy86POK1FY8dko8sxb7piAJYqJGqQ7wJXafYqczkypV5k2gP0AuDL4WqtLfFVcp
WK4q5VjhVwi87kjheYEGd+00GOLY+Cs9+XxkWOr/F824NKQVEg99tsdWlc6cGQFX
7qOAGGONH1/YrymRBvpHtzVFh58716hQ+N1j/ci5m8u5YyjnJxY3n2Ge+bCRHfxc
URbAU5RYFodgIU72RB5ildnuk1oWwt70o8+6bYLubKoAi/auRoR5p2KisjumPG0z
QpjXFa6ebcnraJsb3cjvrgySl1AjP7FtOa4aDlJTmBzr8mhaquGc0w7U+UWGUTmP
LJ+vlJxGWhUeX8a4sEIsElHqjzx1H6DkX+n2mGuTHMV07vX2ZnMkXBEZuvhkecIy
5/YQWyYcH/0dJUjGKzamZf8/Yvnwo1EVw2juauOw76CWj31DybcYTdFc0V6SAPj4
ZCbwZdI31M52rxPeyxoBwRpR+GTwWaGqezx7CXlnDc051Jnyb3o7AQLjDyw6kmjF
GLK9MsikAdw1lPc9iwGUjHcnlmVUQiF/xkYo0+gfWK2zANt6DJSQPEUudDdt0CDE
CvWwYAZtOzwX25qi6wS0zPW5gd2P28Ai3N2HKyMrZBy1ecFsbG5iquC5zdesvl86
YZ9m01TgdvtpOWxOGoWM/UzInjzr33etJJWP+NKFKP6CtWlgieNF017ZTeDuryrR
ql9Ik82pGgDNlrMFM4ORZi8Fo+KZprqMRZra7W+qMEBg30mNRQjyAheNKBUgWZO/
aFMHI2sohtwvM8NSPEUcT3VDceN83W0SNdk/dXsJoo9Cv8rBUTIyXfgaMzPFiwYL
6x1V0rvL7ORxznlpU4+kWRn9VRaVFu1cwQQhUxQ61Hm/6vmj74mxulWFlf1bIHxF
yish1WqAGOU/vvqeb09C0dODZWt9d4q02CTCLHG0xPIynpLh7DuWaWpURXpMUGfP
kYK/FHxfWTFRtRmSYWNhY69tA0j5JLy5btKwfTT/HJRa7c/erxjMc4zam23YyRbj
nQ1mzHuHL+lITSZl27kqzsNSKP5waPFz2SYfomVUjeGE9Uox7gSqdo1khZWgHGqz
IWkd0gaUJik8ETXN5+xvaW+8oUV3B4eh5kFScNYSWYUczzggohnNk9oZ6b6i/T3s
WF2371Qk8KigrmK0LdYrgYVu4ZFr5EEvKKQDVwYRmgHiibrIBbpUL/CJCdFg/TxC
FYXlK5fInx1sGMY/hEm4VSysIcrXuZBz/u/3K/GfCvyYJQrECvbmelqXbZnvnS5d
XnWSvuapnikVQWR1p12AEWlTowkk3ZPeiZCx1ezZbwhh/UU+YK+WaTxm9negfjlD
Vts+ypu1UQFBoiPQkQARoixMOsxNUA1Bpxeg6kgSPdfJrJzJTUeR8udl+HBpWnh3
pLrQF6GNz+3tK0WjOd2VCLwxBabzSHGPcQJsACSJafXGFcrXY7h3QZqQJW5f9DIQ
UnOELGmyGnlqjHl2FCSZI6t2Js7BWzMwvJu1495NdTqRa72FIAE+0edSfJnjFWKP
MznhUdDeZQMy8NMowBqk+t8jIN3TawfHRDwBGWtyyO16fGbfm/mEE/MFCMC/jRki
okaBxGVGgRtJW3S8vWaTS21bky63XlM0pTI+KWNy0ZJz8sRU/1SGnzXy/c/RBHkl
g9n/yCi4Mve94sGpyJfjzkiSqNNrYDtLMvRkAeOJX0lXHOH6m7Y5RAUbus7Dnj4n
aavtGnH2UNCuFkw8gfuTM1qruux31WqG4v/nrQrqgnZg/KJptxF8jVnqG16lQ/pO
JKpsar9GWwKKd+beQz/qb+jq2uUyupF/lbf4rU+yQh+gN8r0VrgRM/mYuGHg+bOl
WUw8bgxLjVfjytMPCtvcQlNgARpQx64bPQEx93bUt0Xh3A+xnGmw4xUJrZXcY9oN
Pm0czVxe+XOE8GznmAWShp2KLru7irog+4jXGqYdKRJ6ash+dDtsM/ch3j+qvJGW
e4GTn4WC0cHAreEcVhvC5y6Tl/BQ/y8slEVr06cG/OQDEmCAndpMTF3mmwerLQsZ
mvcgIJ3YZ92X8nLRKfeXDXnJ2e69NEKzmiz78fpxAhGDSznp32S+WdO1MDxxKj1t
xFTGfxljVjnOby2IdOrHVJaD8OcargWhfaUCUMS1HWABS3/2iV4//r496EWvwEVy
GiVnxEa6EiGckXldYP0c8InZyLTtldrfThzMHwwwnSwFdnxZ/JFqgyZkcVYmJrkJ
uZZ5kn9fN8xV/cv0vuaxevkSCbF6TeL+y6wy4suluxT35bT3lZ6RFcJIV96Up8WA
N2LVg58kHLhMb0aO5uSQ19TUbDnRJIMuGp6gfQ0/JxQd8oJ7dq1MEyDIu1v2blta
sPkDNy1Hp7GDZtdvFEoZWPFntHimOrvyBbtH7tA6bEful7R1NZQVPkn2jHqK2eAl
L2drXBlqpyU10lh7kLS06Mrx/ap9P4onsp4pZTb26eV+h+/jot6nH25QhlNX1cuw
o4w2dj+J+Vo9iLItraOWXwccuGt6MyXCYds6GKIiLbhEOX/Ip0s8E5SG4KBbDItp
qvtdu2tfigj+Eybn9pSVjFARrT7xZSZv9QzM7679H3lDfDSZulE4Cf0Ufg8eJJof
p93xCAgJXeTYLwwWTSu9pNnO5t7P72tkv3sqTjHkPl4CPGMN7baF8waC4X4EayJZ
iAVdvep6q0Cb9HReB8yluVCmZLHvihh7IrlclyRp8N2O/CKGPu/HedtXZ2DmhWTm
3TQbjECaE1KL9u6wRIz5sEf4NXFgCXXNydcWgxdMLS8/32q2KNWkZmLFscr2yENB
PRZ7UrLGh6bFLkgWAN+i8U+9iFDfVgy1vH9i173/33BhFsECL6PYo04RjXx4jSt0
9thG+Q8i39GJnJO99AQ0B+xj53KrVGS/EVycWBEaBqgJ/f7NMe76/WxlACSnAEQ1
1J+8rfMe3BKwd2arIEgsdIuVaKxlRBwaOQreua0HepP5PIFTpCKg9Nmwl7yv1ZSn
/b6u6b6mKU0HWHsvqDyFHlGaiacnz2qdLz8GQLQ3omEWUaioHnMw9dhvdYRs8kGP
zJIpj5BnWaa4K2gGZKm9BIpLe8nJf9s/s3AR9qK7ry9pG5xS4zPFBj+DFXeZL7dE
1lnpagxaCdUTFqUWSWeE8wTqFH8AodI+pmtxX/vQ963qHyCzdBwXNc2X8+7VxA3q
uyzCvOOlUOWxY9k7DgXaN3wny9cx43zP8wj90gGXryBl//tUSmKsCa7yJnt3NONJ
a7eN2ZmIlHrSdi+AIlSBjQeD3/CkVninkMnA10nVdBF8dF3+Qfryyb6izpGa7TTV
EGYlhFSVEar2zKAsl9cgYHJ9MDLfsaVjuARM155ToebXDRhcNLsExHVjZ28N/nIS
wKp7jLNWC43Q7zRPedggD6uhU5SxmW0tie2SUDQ/BgN98gt3Ybc6DN4cpK7zb1CZ
mjXYvAdPTQGr2N7dEg5xz7TjzWbN0bKQY5HXVRlxFw/ysWEl52GtwpL976vWyMC/
aJobMy45rIFWYIm6tnbGw6+Qcs6ZUFL3mi4Q9JoLK2ejqXoTcp9BsCrTc7BjIg0R
vAIIaYvU99hLg9jzxK7LHKzedaAJjuLhBrmT1YQAwo8/jv/iLlcaRcF7qWXgJcfL
SN6LG9IDW5ZMYCrStMovgqlNGojcm/wvkmWO+fz7h5iDfuZAiMTjiexAuaAIVPHj
IufIp3Zq7fuwU7CZu89Tx5xrnTaZv8SGKTm1Sz6zgM1Pm0om8ddMAsSYALAVgqjN
+Hh1FMs/Lfl9LA+WIevH9jiXv/h9iqpnVWUGp2ZNtRDnFbc56dNKhgnKEmhrRmI7
S4r/soGFEUQTMhjT3AOJKeC1rkyTggiaEnlUkGE15aMJsbWEtBvUaMEypC/AH7cY
SRCDSpMYu/cCyZdJKGjRcXTL+vFrfDtgYOlORlsrRqkozE4i/6mCycPAktW8GpfH
rf2ReHqmhT8ewK92X9KE3aFGiqRWPC5K0ZizEbL5ygDtCK/axnQpNjmT3cRkPhH8
PMaKgwN3TvjP9xv6Yam+mRhq6GEcuuAS6vHg6RizXb2H3VG8NjBGC5lCGsrTygqU
lTz8tRLCFMmyFLzf5+5luXW9ILKkxmCtmq/guz2oEeEr9pZl9y5eoYtcHaClEenI
Z3O8lyI7AQPWFfX7uN92y7hezFcS5TnJzQTXVosYpy24TFsu0cr4GcNlBdRiZoeq
+Iy8YAdPlL4Mu4wDRGrbgKux3b5WpYUWMybNTHMbm/s8aKbwbxDqj6XWdXW4A+Km
kV1XM2H7YzV7Y1IQNB2E/UflYPP72QkWeGpUPtd8a8kGEwOtyw43nK/2B02Ip+DR
Y3RaUyvrNOl5ooFKlrH11KSC55ru9/uQfR0wju9ZqCIXHHCN1dFBksfK9HF1i7h9
dCFxxum4LvQpiilzhwdawT3CwJVowqSU1n13cJZNIBn0+2UaKkWCb3dnHEl7hz0i
2JtF5NRJv7bnjOUnfrGLiFPQk2pjKXNeeSirhapQTfHXpssnJ2IjZ7D3hTscq4/O
mx/1gLcikf5oODTBwWgGV5Yeb8Z2m8Nk7cRFYxcNzd65ptci+noSvkZb4PS8DE3S
WNwZUjTumQEPc7Kbr7SmQu72/9ADWRY/3CSh/BLamsgamBP7bzkPzmitFkhHbXFN
aJrzK2lVD41WVsj7DtLt/pTqzjC1DwggdaY8wjS3fxoGN2AiS32EzEG0TQDAnkzR
aQfAKQUEpJ6dmALgWMg//xK0zNnfqYPCMMiT+lYQ3WHgF/vyuvClAr58AtgihqtG
pVciYJskkFBB72sogUP/BSV6iKeFXGy6y3oJ9jYZxFSnXHG5MQnw2FHP0pAZ7j2d
R/iACOPfCrZinkiovqfFpVziY9VIOZrsSHFrErBwtuWNYnCm1KEB85V3ocUFd8Ns
hLlcPF9SEHxD/XXBsn/dIEf95VDnLjn3KsW+mW/aHVdt6+eAdokPV+yg/m+vRiFm
cTnAXpb7VVpIlEG+ndvKgwKEr9wLdIKuR+6Pvagfzd352iBgsJaCBzRijEDH9iC3
0SPazDsuNOeZLHIGwFj+dWD20rozosbHrKDi3W2g/DWXtZYXpNQE2GgYXzDDjIUf
aC3EMSg70k9FSt3iU8nAehl8Q1FsPAjJXQlqhdhgJEEIYHlRG+PXC2zh5Uyr2acs
gJHg9QBL+9KxMjzKx4xC1bk7msNKglUXARgN3eNkauZ97g/920w3B3ndQpOiFpvm
v0YfbyIux8ZW5wbXlcJhyiwXLMY1kGilwzhvH126qI/WTUUVl9VP3li6H6WcWnMm
k1a2HK1iIyCyOtTvRK8I/Wb//1VyGRDtn65XTPZZV65Dh8J4fhdRj1JThWYpOOzD
irs2r4N8Eq0wyv1bJboDJG/ebClfANnxn2blWW/v8ptzTN+XCjLBYyr1l4YZe+Sw
GIss2o5LuUJ5VkmwOQhdoOP3XYEJItpLNgx6BC7bo4Js777xkHGqMFaypyl+otAK
iH76lqRG9sJM0/HX9RDsyOJ3ol1x66Ib4QQbMndiYh/U5OKUQlr+cTTUUHhMKlV6
naWhpjf4UjQGI185m/AARoBAYavBngFrg2JG//BzKSbboEjBs3F/+5d4MPCWJJuL
V+j0FFx43b7B+A3OzBqyGHa8EGJscjpsd1dWSWRVwqn6O4wsX2SfEjgqNC42XeQV
O09p0pDslidfwQoaIdv55jDRnqIco3bt1U2euar4Ma+Q/Aa9ne2at0iabpDcZ2/l
+DEBzpnz4cKckKPcVV0LtUcPpuu90n2/2d18jNKVFHiaWZ8TApBjVfwYfsaSKu/S
JWMl4q7/rsmWsoGxwMqaHtHBvZswYxe/l5FHK/M5itCEitoEIHjTkYTKOWljUBDK
MTzsFtGWFcCfDx5eyID40zPGuYY8dFcJ90Cl7/A4mecQWgjbeRbV2UY/yxDqn8sP
hQe9w8gm31yE/k0Y+AjY4eZjTjWJVKFc+hN2h3vBmosXLciULQ7FRY6X5uyCw7Py
bLjxZCsOQQiOtiNGpzrhKwsPePBruBi2GmvMNPs58XL1kAtLJPyRF5Uzkzli8NSH
m7Vq/i+7oIqhelj+8nu39XcxnT9PlXGh8JMF0bSNgSrIq7qZnrgKBLefC8wLx1Kx
pkKvPLsGfkTyCNaKqTpzSVun2m2ccGtXFFEQbMy173NaCYGzw4P8Svn6YgIu9SmN
7ql/EKloNMNQuapwLuc+2A69JWdRuH+JTpRU4soD75Y6/cr3SgCmD4jJGf4w07ff
V8jraGCniXohCpX3LW4r8dZbdtvjjdUAadeJcqtaYrkGmwl/J7nGg8qkIv4CersE
JRB2QLEysgysr6hVDwHYeT3R4khQHNLWs7EDcJPXEXEPPz+e3CN/DHXPSfWwvzSx
SefTWSAufUVRpkwcnPdusGPI4rHrOYr5QKNR6nbhVN4OZi0pkMBL4aMUzNmatmFd
+vztv+Zv9v4ROenxRI3gtF7FiDL0xJJORzx1f9baOmXlfujx8rRBhfZ9E79MGA9R
V5b5yDwnwrpXxN2vFeKbPjYb4oWbQes1x6UZmY/FdsGzxASDmvnu5IiTi1wT4dul
0LYgGAgVrmuT8mwJYZL/zkZ+83P9LcY/BfZ3KER/wHzlt0pvbJIlBF3Ycyb7J5Bq
l5n46npe6rMZ9uWAACC/LnwZjIEwpLhKMUJoyACYkaOb1SEhLmr6qTR3hN6Dj0ar
ID6DUMMKAnAyneSUvEySGeNDds2J+yT8npCwVQd2Xv2oDs9xCj1DubK/pXr07H9p
Ja4ptLM2ZI0FmgFz5ZgP05IUzBYVJmexuzKIJNFjlZOvWYplXDpUZrLS7AY7HpI+
6pJN4g3OHaK4FeZiXka+F88UleGKe+txgBftk0YlIshL1mU12vnovyX/2ZX7TjGD
H6AQyOP8Oh4d9l8LbV46582ivm6CNMH8mZvbrEXwXy34rRsnugGlVY4OzZyp4lQ2
iMQu9PSqnuOINsltzn7qiWPIhRZW7MtTQ/t94Hw3Fjxk0lSkqgAQIjrj053AGHtC
cMpRYmLtVDP/geitQPqKsq+dGwG5B2YbvTY+eVBuL0jqcugN7CRWeX7QRA1v5DQg
5Mqq68gJ6nB6Rvs/UV4XkSdD/XuGFfspjJjDvjGjfNNNXc98e8oUuy+bieEGkuFQ
47/UOEPX6rFZ4+hPxup+06zVgRAPjwHBbLMEIIb7WQkp9gPEegzRrNgxHKchOnYW
ww52ZiF3Uk/u6upITiye2Vj6R/g8ZmLXDAB6pJmbS2qX/EEKqzLgQbBOu/2NQOrV
qmn1MKQwH/Qo6PPWi9UWv108J+L5oJCiIJXAkdiTi9RIib9i2rFNfUUMVcvJE9EJ
ag6H8TIYcquwRwIs8tBN1s6pni27m/RyOdqmwqPtOq52XIlWyACZ/qfNh3XZohL3
KmMSRXE1gXhtNvH+rr665/GA8yB8XXs307f7c1KrGuEmZqrxotrDg4RNiZiuBmHA
Uv33MXo0zbos7cLkL7cbgkpGyUZa1B1jvoxu6Lmj6d+o5B+SmrLtV2XL5JWGP1rF
iGLHJGIJLsg+DSq6bRFLxHNscpIANJlHaZFtjTaSxY0FTBkW+/g7h67nQqkV27fC
7rQ7NfMVaOsZl3RjfyxkTOQBYLBL44PI7KxwvDtGwMFCPApEDrkmVoecrZdzB2pm
4ASybSw3W7+F2EilT3a6M7Zm7J87/uaLOJVn76ikTAwJF68e5Y75RiIpCvotT2iE
iMoYC3sTAeBN3WQjf/8T/P58jrGX/6TGABtDMB6cyNHPt2uYwMa3d++O2hz3T5re
CB9qcxgz+rSJWKefz9bjfU4G/FT4oGe6tun/2WgxIkXVFVrw1Y5+nju0z7jYdBNm
qUNzk5htgBgC7dQiFJbiJF2tP8r9IhQkbsMrk0GKii+8dmg1wFqff/32YTh6mIAs
+UgoPSJ14ZVqRXE214FOR9bVIC8XAKv+gbQvoSe/Pz2ubXmV9+3twR5QD/6cgV6/
RWRjUfBY3teGSX5u1CFb35UQq5Rr9EIq//FNVvsPBnDB0AcJx8er/f+IXcDExv5+
orieXb+Hd8nGpLME/vHTmu+QxMvAB/i1fBmmlsWW4hC5vN0VchHkuSz6oAeZXtyg
ttDYu+epggarrk77PTAqsVzNHVjGBy9kNEo3FOTTXyo8bqVyHDifN+XP4lpXzfo7
cm5DeCPp1WsK3JRMcsqMZkrvqvisEh4K5mg09Y291WD68vy7IlwdvLfRV2bgt/jV
aewmUul2mBRvr4b4AhzO7u9OOuPXcwAPNF4YToPeDzrS+OgAslm/GzY30+KqYL5N
5ewJFcFH+K7AgLQyxJOLhWGZwqeCbI7mZLtzg3b4Q9GKaWbgljW5iGsSg4h73CyR
D5iF5Gk1892K0qToQ19zkWgRDXRQAmlxV5kDJ28l6Cjlest6qtXk40NvAnTReDnt
oaUdgOkiArco7/vqp7r1KiP1XAudsbvDePqHU/24Kk2+yJWluIPGVz9OyPixxpzL
W+kRn5gIjSmhwPrwHRVodrJWZzcT64cxamfJvzyl/WDiYKa5I10ZTo0Xp5ONo3kP
46HaQvmarlnZax3H8hLnQl0g9MXyT7JXhUHbLrVZXN1m8m+PXOanq/3aIHxxAjxW
qdrrcC40sH7/Bx8Ff0FOaCodTjlUaTreUNLvyKpPmwdR3x5BAIzWAG14mGGxXXhL
/1PYF4T0rud2eKN+jQkBJjGJjCZFFq0/kiw+o4Lbh21xaoQLfk8l0idYhY9De/RQ
Vp45mRArRFvG82SVahAKqqZxHTynvdGhViptNE+AV6Se0wb7xhxeXmyzEr5uaQpi
d/bGMcSx5mxrSZ6SpsWU57xj56EIMXu9d/wJa7lZR+zcsmz4qNfYTCUbeylMhZNt
8jLtgH3qTgiFpLctQYCfIQB4TfYEFm4KFyYeBqXbavhLRh60stXm5YH1ckovOrwi
Kh7+8VlItOEes1CXC5czpFXlqB5E9SWA0lTPZ4Q/mpcsu54bT7NxVWl0ld1zHCm2
tFmYUca6Ui+XWkpCwLoJxoB9OPWlMP62hSvrbnAdUPk2beJkkVUqmD/oNAkAxaev
WEomHg5/MLl3Oa2zrLhTrHszMBbpdMXj8ZW+kbj/Oilomegd5iDcrLG8lzp2Clsd
Xlr3aT3ESBaqCjAmDjd/bzEHt0hVoPFX17O1+HTxr6+pNvBxwyAmsAHjLP9ggZbl
XlAj7kmvlx5QfzuWqhvJCHEM215A2k7LMdeDtDlup13QzDd+SHzYdHldJazzV/xr
n32QC0VFlAQyJkC0s/ZIidI5jfBCskPIAVcmvRKpYA666KqlMJIIyvPkIc6YubMS
i8RRgBiyRZrb6Ye1Hx2X4CMggZCMNPDf4sJokDY1qmKjDVDV2/KSGpvVCH9VaXb9
g1lr6V6ct6Ivf8hHIt0e5xlCaydrvly/YxkdIBq1aXO/TNXbxoohU6cQbSH4noqs
B5wbBtnolt1MIR/NWEHRqLbV4eLPneiAHDvF1E5/WDsF5QJU1p8p3Nl675mlhwvz
ciLRvh0nvS8IqcTw1WNYumxZtRbjrwhUfmbn6TjDdFJ8LQ/IKj9kNGaydeMG7Yey
IQSZjcRJOTfo2XRi9OamP/CGSPQCpFSULklmQLfEg4DAsu01dZ35bQmfVUxvpsaV
5h4d8YsSMlFu6ou0U+SHcKWNeRKVP5zv3CbfZzVARIWswDyczn3vcM/LTFnqLeJe
Vg0TSmhL/37M8TXAStBHwssyswwJcg+av8/yY2/ujL1rUcEpVF6XX9Sk05pnrECb
XA4vuffrluPL4Hq0uUdqGI1nZhTjLD+VflNH5oNbViKoeVFW0O9z4IXkTM7H3BeE
1Ak/PN/348sUmIwb3F0eJNTC2bDSrk48q8HK3kRQXNisswkLbqlAOKVWL+keJvF7
/tpEv+gEqLk/fLrgTgPborvwlPWewprGBfKFwSIv62tJCQBsyMgpPA5rd+jySPf5
33fctS0aLnRFPURcUwB4gHibq7tR3GrnNidq78RbilzEE2L5BIv68FapvkcUp9hj
6i85rtlHShAaYinNyjBDPgVNwiBsZ2i2gy1uhRxiiKARVJy1qVvQpwpbY88FF2ME
0s+3Hpmnw9NHENLkf5iXe9WrIEYFbNtjxdRZ1sLzgYA12KbDcwmvuhjJ7xyGvD9L
dUQeTRiMjgIWTeayOAFEeV9cKf6BXFz8cT7vujj4mZ29wZ/24hAiFy2w3KrTTZx7
6AHpsiUGjpLQF3xYhEUJiEt1YtkLr/PiUER76cSW71QAN9rIKZU/zTXtY8vldgic
aKpNN43HqnmPZgg+lMt5JySmtTvBeM5MUx0j2+sovnreu8f6Zsb+mbLHxtf1oFaU
mNGwTBlkc8UXrgrAmXnBVuNtlad44Hvnrl2ZvuMyFA6FjmOgbLDLB2tYln9XogUJ
qatkiJ+Lbq5md5E3HZ+HKb1yI98Kbpwz5XyWI+yIKsa3UL1PnHUoEdFIITYvDaAa
C+ZMjwQYvQgKgEQC4aVhELfIUyD7SBZjrPwDSdX4o561qVZSYJjAKVtr/aLB+5cQ
Eo0OEQHXmVLl7HkgADKZNgJOa1rJMKk5f5XuP9Wi3RxhE6MO8/h6T+B5GT+Y/vlo
1SwNZc6y4glEQdVSEt+bcyqcd2NyCyaSS9JXDhYz44pSn3G2pUfzRDThYbVtff+I
GquER0+BttAX7L5/PjYLzwNdeMGulGbkBbNizjdXJ49JplvOI5dFoFDr71WPcWxN
eiPdNk8q1u2b+G4uECxhxQOcvlDIht2ZGHOBLEMGZ3RWg77FCU/x0ALnWzV8uh8W
nOBIkLzr0+twJ9RojRd7/4wNS0UmcDo3e6SrTcwYyMtfPnRiocrHIA5BeZgP38u1
dJ8iLpelbHk6bJvQSKyWDboUgE6IXixnbJNkd5o1WCFWHnPapdxWiOGLkUooMRIi
YgHzdYtLdjD8eL/cdULjWRnZL5uUAXXI920ZnYGCdd+dO7xei/wgEHKwhpaGgBSW
JCav1mptQ/jD46lLtAa591kfIRHuQpZw/NujGarrbk6JWV9Pg6Fx1/L4ddaDAqtR
lrDnC6kDuVqDYDhHwO3vYQfjIK1WgXqlgj+qWrrFDmMUtEIzLcWLFHB8T7VaEMVj
C3WyU8ThGST8CtnIGeoYaxTt7Uts+bFkB86KWjj2a5paAmjQnGAApfLaowiElkVK
zQHaR0YaKVr3fxTF+hsQThbf2vjL0Y4jWF/orHlYkbpFvnw3Pl85bnIYOBQTerT8
C0HZmJSyz9qEgYK/AXQVFbYsdzmnvJ7VIOpwv/wzl6hE004f48l7QvDiBg+TczVt
xO3hiCKMjOh4swMpXnxcXaM0y8r8xbX1W4QnHvWGxiL54h2k9h0JMt86XkIRm0uQ
xuL5bDdmL4A3wrcbnzH11SZjb4l0LfM8xp1cgxzRtoDkC4WVJZtuecC5FK+8HYQA
wmKkFre1ASy2xR71ysSQbRWosLyvs95sFW6JGY2xexzRl8qvit8T3DCl3ZHopU4U
NJH31eJyFGFik6xix4ysKPtJ7qcPHryk89HikC1cZSlV/i++BlHJ6xmoOcFtCnla
b528eX9f6jk6v5kVhLK1CKn47XfNoUTilRG45oGlFpROfdjNm8+MCC4iwLuz3kQU
Y5XgZf5xBmSnGL685Ojbwc2RdigLO8Vd3NEmY9NXyufm1NrRW1+s1RH/FbVEvfXr
cCrTDM9Lh7ZIulCwBjyU58WDSYbGmPuz7SX9pZxMQ/lY8Ky5+ygpwXAppLC55afK
Zn6UsIfi5vHwGKkJi+SnF0jokNzQFhmRnjq7h/dNE4Jy8KIKCxjxCoqGQ2sq6WFX
m6i+nWyxsM7aUUekOdiVxNeVdyrPOK17SnqNSnGJZx1tV01zyZy216GfcgoA/zWM
Y8T/NvzdTaoZhOU8rSkAiwB/SmdGGeYjkyGuYZghLCacWiI03Jw5QGtgMH2BfJR9
2qWzlidHrDR7ovuB5LVyYGJXx7vJnkIWeWnzy6AYHTbvld6bQek/GTj7gMM60zQf
IoeU0HO8Ho2I1lCk+qZTJcndpufvqTxBYqSEkrjkczJoFwGL149tYFzfdnMntJvZ
WbCBUlXoACNqv8IFrh1R2QoIYMLK0Gf/BdkIyzvXXrT+AK/u7RPc8aSxp/i37koG
XJOQzYn8G455ec/lfRTRV6RrPzhzAFhCOfLwk1tkbEnuPtcMzKhL5c0n15WmA8gV
Ga5uik6lm3gM/9zF9cD2UOCq6FLP5VC1HadowRGf0YH7uwZjc00WHixo6xudWHYD
yDJgNNSIwVEhdvXl8/NPTkNZs/HSIFSdUMsnRzKniD+UU87keRWzn1vNqpTs9J6I
mALGB8ZKBNRuYP71wDyPQTIKajEG9wHlQsyMAF1SDTBogU9iCs4eHVSmRuXcn2ED
7TgagPWWJazEYEyQi2k8VGS7B43xgLbdAfY8k+W/X57boHxWOASkmoBFyZb4Y5Ml
JTybU3U1O/PFGRZXWrmXm09D92CRyNkLtNLMEPdP16L6UhFCgO14m15URb/7oiAL
ojHDjUr1E6k8plz/bycAg4GKcOBLm2Z6DtmcmIptRzqDA/05EqwyOcR/Vo6k1NMz
/nbvd7c/aNLMkLjUMNHv/dWdVqLk3eLxwcOquwXBXJNfjt6JjaEIS/a0HPYuivqm
Ghy78LjWHpqJyxz4Y6HwxwpTvmiHUlQtakUPQevysdFSA2ZUyutdyRo6pJqZKMV+
++sS0/c6wOQPXHUj1CYleF9aDNadojeN7idBVDmLXqOmNgK/bBrFlpAG7PKE5RCI
sCAU4jfdQ+rktdMm9t7CStJlWJsWMI010G3x7LdpJjS8/3vTdnjef9Xk30JA06R4
8/DNZ0rRwYFxLHij6H0fEcbKnRC7uvJoOWfqmbU1EdB4MrWS5cu0hHO2NxoQKjBO
TMX0nyAQT/c4sMldbzvCLM5vCHbNIeks2uIbT6L9Cg0tssIig+8R3yTYdiFZn8nd
O/hPYar3I/J6M+LqHyGl41Rz/20n+15ESmS+nkKRPj1muZB/bpI9LZEslTed7+lz
KbtBayMrxcHSOvaJp7b7qFQPdLlMrKdWHhr1RMF1am9Wlh2TwBVIbZcz31WmfqjM
8qCaqhBsSSAWUnwklAdynPiquTTnzV1JlwlIBe0IPpstzNi0kY7UM58rY84jtrwj
jxTkltnE7h4I9j2wMv4Z7OOvvS6qrjcWLQAeZgCyvexo+BFIlCE7JgozlsfRBBX9
I0XtYJtlU1PXVXpSBGjtYbYYjidf2kquzlW6mZUL96RmJ+CXGamgasW0B8K6Shia
YKysppioQvw07p1GXtxCBiAdV00NBsQ5Fu0ZsZ270TEuwOWj7giyIoO721AlWBAW
R7sEQ0F7USvFz/PMCHxGXEECs9Xsw3oEmakCm710iSblaUF2WJeyFWXHYCZYyJK/
b0m5SjqIYiS4kfOTqBt9mckiw07JxImdNFVjcMG4KZhKc0TAngVR7nqwFpA064y0
Qog012VqXTKZAkZP5QaVKEfpK6f9qB+4oYZchJBRdwkSpVhb6R3BW/o7T+dOPCRQ
bfnVibFq8B7ACfg82oPGCmLL+kqzl7mh8M0Yzds8ON7/wJH/UWeqZgKTTt3wxAzf
illIfn3paEOgAOThxl9+zCFCG6ta6neYZWR3t3X3xXyxEN1mshCiTr9FDZOHFSkd
sVLo8+inVt0iyfd0f7PD2WVXuav9QEg6CfXn4svBBp3QB3KTv1Wafi6vEYX/XSfk
hmoRtgYuH2QW0BySTxatupRuuKWxpTrayIE/pYHC538OTZpftZ35usk8Au3tQuZj
jPOO49jnwdCNhLQyDnKJnVHaTL7x4S1XJ/R4Fg49joMLth8Qt3FAJtl4weSlsqkY
bDB/j1M7t0jvQD5PuJSqDjKkyU22/3hT04P8aI/naPimwNoGUk/QWaT9GcPIm5y5
ZX7Syis25aXnC2cyoxpxCwY40WzC/kfYaCfkdAmWxkD3Z8hqgouxEkP4yKdfqwP6
NxPmxERj0ajlMe/HGGtUYU0FyP1ptyAU0jJaGs7DN/Ag8F+H3cjh33yn0z0K+S7z
Jv7hn5AqBQ4d6R0Z8+5jfzeVjMDVkCL6ZKY0rAnQHwtGesXfjgaNphX2sNlB1WS+
5NDDWz7/8NdZiV/G4Dv5LqYhVf3/j9xvATOISm1MSp5YjjUHV0a8bgwtDQJHldVG
IOvb4KcEOrlX60rvQ4lJRgN+Bjqb7N9arNyPdBTRte9Bg90mr5PqGEZpsPUfBxiL
tK6eimcEigNCm9DIt7LFBoMB2tbETI8g/xly0a5EWp4Hbrkp1EB7hR7oANgCCI/6
dgcxaTPcFnayiXxoo9L4nsfNeKO8Li84S2vxMzPzbXOWp2jTo7a/QZI4m+bFHkj5
g/AxmlWtFfepXvcWxnfyHNGQQQJR4T+P9qdgB34wiMCjIt/IJT4kIGAlMHO2r8dD
rF3s0N1wW9JelLfrYloYUd7v+Kj4dmnoUHWkab/T5lyH4gaeNKsMAMYrSmfSoHDU
qXSV/wN2pbsKr0lkgg65eJ6WjD6ea++PeiTX/y2O9TPnUXK0HZbAw0IGNAzq36IX
xN0/7Kzc7DjiDcNgvdB9o7kDVT6NX7pEUmvUPd497y/8xy1qRhxl25MEGQmlfjj5
NMV5ps4FONbr/t6Us6HY8wUSZkOyCOEgwljMu78z44Sz8sZNiXrhvnRelrLOLO/G
/dSMOdY4chUMf/IHuW2iWG4eOjiUmgxBZRCtfjE44d2kVlVfCTuYQUfif+I1PM6n
GFPiEuj9QUm/c4BEGZC79fz73bRxBriFLw17milpKPpZRnBs5tAqB0nufa2R9byk
BXwq4+Yq5oBGQiwrHoGr3oEi9LtBIIFoQ06Mwqe9ARKNMhytoZkEykE+uqj1lnJe
IqwDcWgyiJNHuOFZng1qrWPiNmOhv2lgraieL2Oxg80x6majWDBagxUtAtSnzMr2
w09OdCFA9ZOZrH9rGfsT7EUqRId7XdcCWYUYrlyIcvFDhREAIsW53vK3xnfZ6LOa
ISQPU/kSgxOJ9z2+8sRs0AYS9gcbYZiDjKqQlMZRaE3B95qAy9OLduUBBDnL2ws8
EFHs3bNe/bit7Ix3+X7GHOxsprhekFq0A1msllKvpAEbjY9M/+AsQXqV24CoLZw/
jX5W7ejpWkSHR3BfF5M5rS5CW46kN7V9sCSb26VbCYEXzkwXsOZxCOIn8Vz0SkLT
+3QhuiReuYr+Q27cTEubIetapsadxWJXQB9w/oKVrysIWIyFbv9COZ5gInAdYQN0
NTIAfBTPZstEVmBlF2VSg73+mdRJKp4xwgE2UOn9Dha8Yl0qNHvdJzrt0j7pYrCp
Q6G3r2M43uflKq0j29GzcK56mUscuFr2wXpo61rfD1LGelav3HqA29d7RWw8RwEA
dx7abHQEanykG97baqtnPgg2xsQ6VXnnQXsbrWIXzDc8ovCDb76aio/O3V5pDA+t
TCB9pvHuFvtJrxlpq0/HfNcjn85LU4+DFincydfeq7dyLRa4W72CMfURkDHNLvDI
qbWqJnjLmBKiAMmEW04yHj7WrwkYhcMIUJH0YN1ZGeuLM/FO7T/diZBkpv2B4jpR
VoPy4SvCZ9P0BTF6jiJiB2/1pSpJC2oKmAMnYOBmq5s/8SfutLcSpYWTIo5KJ3li
oWnidJD8cDM2oXieayWLqh44gbuS1w1DFQaZojS3sAsbKL4LkFyjqo5KbqjU8HAm
cio6T6KJt+gOx4lxw1zfKkWjWH3dBuTQxNBJYITXYixDY0n8nUAmxapmhkAh49XC
JNNkVcdtRBgdTTD+cV0u1rxXMR1CyR5hZxgkbBw67+pCc6ucQtkr4gAHTYBuomwc
EM/n9zPnafsZv4pXq29LiZrNPxFCdRUMvd/5TItQoPOoZtB3d0qdjIwBhY6LKepR
Z+qeNR2CWKWUXjtzIxOphaSEO5rOKZJvXHNiMlOkKI/S26IqYpZmtzC7Amd5eCtC
IEr5xwSpa8iYF0XPEYlN04fUYG1rMv4IF73W03OsvpK6yLWjV3a95Xr8lAJzszi9
LSpSVLdLaLhPVfC+Ua8EMgB/K8+M6zV9Ycc6cBowEsmVBAaDS4QhlYRvInbSdDyv
1zwQLnIBUNd0ZZ3xumG1WHplQ6g5vgEScwbdJpcirIpegsmynD/AjBcS/ZeJsl+q
hGtO+EVYmd2GGPEuBoB43pItmNUBX8vCJJKzF9lu8jHYg6XB8RqtIU1RYZv//S3V
OQp4/GscXNEuHYiToVsPhTzdetOvdwYfC2AIvSnFIcG74N3H/MwFPb4TMPTSFOD0
w0dp2UzDcO6ptMKhk9WHJhV6mtWZoMX/7f9J23dmvp4bQ7V537PZPyCX2j4gcuyV
Ne+avJGuMQI3bJUE60vEiVZwB/XzaOtGVOkEtDNR6IVNqdQt7pWEshb6UUlT7K2c
DSy6I/VpLqAge77zzqdMdzYzqxr8yjSAfl+QGuHXbE4+dh3+LS1AKHukSodrVwJ2
3NSi0YrqvgohJfnnxexJfPbxfMJ0jl19oArjYeFZcllx1haQoLqqs2/8kqaHRUlM
tqJC8qfMLCiCFmea46XgkoCWr9p7YxURj2AV4mbpcpNVn/7PIVJSiE6+/0kixs5u
rBQUsLcAC3+SbSTMdszcQo5k3DkL7MqgoN+UR6Xe82az3rwTvS91FY/gSAzmBU7q
WCTeiwWaTzD2wMtn4BpQRSslOJONk1SsC849eCi5KaCWCcw3dz7uBQGiZn974+Nr
w9GeAlGBKb8SoqqKZBs0B19bNWn58FLYqx0kgEb/qzfkLt5LMxG1VIbAOZXdKFU9
Jw3lvAzDQ90T/lyEib3C5xOT5rw/9eEaiG2rxd5hNi8f6gbPzy3XAePM9M4nzPpU
TaUU2Yp9DYuW7xwwmj2J8aquwD9R6ZGVQudYYYHTcgaNFURlyM9J3jawWblLCL4U
yvMZ03P5hFbP2x/atlxcVfbSdHCrSWONixcF175NsqU0NzlcpAXPKWQDFvtdMTwo
LSle/pw9fjn8Yj2mJIE/CWfoewMjFCn35uETdVoWmtjJZda26p0VXD2icnp1zF4n
2wF9g2z8EuEaD9HYN6E3Sh7j0yJkQhFUzfZkZ802PrJDZvSH0U5flApzM04BoDVC
qAwvyg9Ge7JJxDmDn5p653vUg0opM0rvL6rvatqoxhyUeZc6Z6ODESgV2WmrBZOF
SB9tXkOxfXcehgWKKK8XohmDsZMZp0qQ8QyFOCDxDQ2tN6Hko928dVUGB581v5bG
4KBhZVibtFbIgaQMGmOtoGyM47I14Wt/VkESAe8rhesRrHEWWvt/WUwk5AnN9XHG
0/DEZZC4NqWeVXliiGKV2DQyYYib/upcDNBadExIV+/KBBCHiHbOflgOCKXXmdBk
sIN0cGzDNQSdw1WSWpsbg5ZEJ4jZ3bWml/PXIg7P/AIG75c4HPK2VhiVi0bX7KJA
X3nEBPIx2i72KjeIvd5DHDRC34rGnUcDMobn0fZ8Ggzng5Uu67o4Ojzm5usi2ZWt
xsyONhNbdzqItyCHUfO7bCj+QTkuzbJOkIc41qYi8gEKl9dnoAf3iTO5pRNmwRiZ
Cbsszx4Hm3Cvs9G89h8UcWqtipebjAVhnG6zNNHtoz9aEArYqMVxxgJcv0dCOvog
e+3sMv5WWz8I0YEjLcoZcjPS201v3rc+bXzGYUPtgNNQI95mXZltusk5Z2oxgmRx
EmiEYy4/kq4dH8+yldtCsa07Jze+0m+oxNI+oQk7pgP3HWuZWS0W1Xc5MhhjbxX/
1pE8q0ea+hfXN5PpONZCxjNENWmklbdwU8TUpHup5DgrIw4z1KQKMbNnhorMBzRp
bLcuHaVeZmDT5t5IU3TkWBJK++Kb7zRmbmHI1Lgqga3dut87VfvyBS0Myg9SnaP0
onpCRkkY2FiO/HD0l5E4kv1m1/G3QaYLW724Ve9aPsoghCxNLxqJplC7abX5ZnNP
oGHq6f3pK8puYVzTc6gVFsF6rcMNjtkFYwZM3C22Exj4r+c5qnRnhfMmWIE3ukDe
B21x8Fq49ObWfGyxegoMnV6m1wITlBYOB2TzyNRZHlk8xN1bxZL8OYLHknvvBl9U
Lxxr2WBJMWPC8hEvAAmLl82/a+dWfeWCdIjqbTB4L26NL7BWXB7e8RxjOn37aVVv
WDl0KF1sogSU1aQiBlLlPYrIxFMngYF+/vRA4QTCZH9gtyk6nteSyLOP6+p4UMs+
/ONqKVHCdJrQPfaCdY6Ec7uhShEX8leplTgswafEecrVa/7T8z66f+Cr8sqm6DYd
LM2KmrO4Eoyc8NOFn1/rxgLtRVB4W5GBOQDaweBuhU0=
`pragma protect end_protected

`endif
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
L4EBOr42s7NbOQP1A8IGEeInYl1cEmGybQGFCXnMCbfTj6K1IMLYfMZLdTxdC0mk
Ca4Aq3FXGfnDN+FHdi6fOH935W+ma9ioIRbrPDPwSKMEwHOuoiSgUSSCHM3FMtC8
B4zFydik3R4LfxPQUkW3Zkq/dH4DQUhaL82DAJ/erTQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 172345    )
85EqvXPxvCn5hIQK+WcUHGt2VL9/0Hs+BZitS2AB+FY1t6LXIHG990beIXXeDzzL
Sti95tW4aLELKm+2bIGJ748/6LRuu76m83AEMPbLHste+F0EjuULZAUG4MkSR7Dd
`pragma protect end_protected
