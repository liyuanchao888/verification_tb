
`ifndef GUARD_SVT_AHB_SYSTEM_CONFIGURATION_SV
`define GUARD_SVT_AHB_SYSTEM_CONFIGURATION_SV

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
c5w4xwH+ZdRRGucUkDkIt/wma5YJCHfMjcEc1d4tf0cCu4lqm0r1LA6eZpxxrxMo
uG40CEyrCtwRvoAESkm4ux3IVu+BGGCri5OIVGZzSZIKzjD0Fqnach6GjhtO3VVK
WP3SZyEL9CMkKTAgETdX2ZVsQpPFuqtOQKAvk0hdQSapp1HuGskYzw==
//pragma protect end_key_block
//pragma protect digest_block
LfKWcGOHecVlk2ySWSCAWAWJ1OY=
//pragma protect end_digest_block
//pragma protect data_block
3PMHzft9JbGVmhBg8NGZHB0bXgNddJQpCUdnju2Qr5Z6szcvrEqfehzzsSOmqXrF
n/AJzZgCx/DKkcvAf4ksueWyrWiV5nx+PAuz3gQeTmbvxDdX2HEyssRnW/ae/Rr5
NyIy9v6mU3iGZO3PpJ1r46jw+oacqdMw5PrJgNyrAas5wBYdvaexRkQ8LAo3/PPz
tqdiHaUvcPg4Ec8gn+mZFf/HTh+108QBv0DRVunSwn7dLRJzWX+OIK486QrlbzmU
6zyrTVnC12KQ0uTcHvWJe7dhxW+eatYn/vY22LkJ79N4FK0VZqp+d9dl0rRWlBta
Hcst9TNrvNq/hVxKuHyyS7FmvwFfgsH6JHij6xfU4pBoiPWIMKrs5l0kDGuTd0rq
03q826uk0cVPqQYksJByqAD5IJIA4I2e6wDf/nB17dGNgcU7tDo/jYAa4lT7AQ/2
PcqIo1z+gdzsPOCmMbg29wSSyHHtCdLCl22jeVNXCXPBePqknbYDWYOyW5QEhviX
aSurq3IWtRfc+Qr4KzgJvOylR1NEEffRUMQ8q2AN5PSkjXlVhvQs9OT25ACAvBbZ
AbUqFafTHnRnzAdUFtRE9WBiKLz/ooUDG/j0fZ1khineTYFpclrz80tWJdMAS/2S
9/bIZ3pBd6cZ8L3YFb4trKUAk9rb0OZ9K9gYQXeV0Dk04senr7+xyZJxDuARYe/H
2JsDBlORobHVVwjK6qoDmm1yYp83/Ie8YtImdeC/hbJWa7jPZ3oc8X3SQVL6oDY4
WjZa8d6fBgjHSlGgl377K6qBOZIM9M1LpDAP+G5K5DMOEPzpHuXi40WRkOF936EU
qF1k5lUpMY80Btlsrj1N8is4/0uXTdnOTpki9fcw4nbjb4uIEAxSPFtvMQFIegxy
QiYTYiYf+n3ZIJPajB0jn7JF/igOb/3TfPnofZ1QScnnp9RtlpDsdcplgLS+5lzm
scWj+qV8bvqnxHA16p+rSosLtGWeHfBFhdBM+gxMc1ETBHvHxxffw/iBX27RQCuy
2j5B9ThplPprzmS8ryfnv2VVS2rjMN2Waa1qMgH79LzyphHGABHL0npE3/Jvig52
/lfLE2d7AKih8dfuBKCp6eyUAbo4ggDzILlne8HCbLqOe1xo4huKyO6lKEWxZW5n
lLNbK9fkyak4D4cj1jmw0GY4G4xC1PZfctZbws4OUn2ndeSinCQwgXkl0hNTbsoa
V4IKlQtNKG5+AYsi6kiurrgHGMA9JQXTY+BoSpedgn2cvL1LIm9Jv+hb0A/Cjx/a
a5CrBin+gyh0jm8+zN9Bg38CvJgTJOFledNmAvbeOrVASNbVOjnIMQ6KSq8pAAnq
LrGIBUedak+pK+31ncytYfTzCABptckRyfarhO1bAAVg0PHw4R91NzQvStNIqFbT
zRHc/gy+u5FRJvUSvVklv8cF/RzofiWExgtrrekjj6eqRbAR6Si7v2+5+RsSRAJ2
q/uk7TBOJI6g8wCFGUz0lUBiOcfVHWuhFhm4OZlGH15uAmZ/Ed611HWherfxnXlW
ltrMKsEe6zbVfOjbdjOkwkMKwE+QfuKrjirnyaNXJ5So8s55u8JSUr4ri9rs1Qh0
pF856cjVmHLUAqcxT7IhatTxFDWQCTFk8MT8lhJyp9o=
//pragma protect end_data_block
//pragma protect digest_block
xjdeylTfREGQv2ym5WcaChaOF1g=
//pragma protect end_digest_block
//pragma protect end_protected

/**
 * System configuration class contains configuration information about the entire AHB
 * system
*/
class svt_ahb_system_configuration extends svt_configuration;

  // ****************************************************************************
  // Type Definitions
  // ****************************************************************************

  /** Custom type definition for virtual AHB interface */
`ifndef __SVDOC__
  typedef virtual svt_ahb_if AHB_IF;
`endif // __SVDOC__

  // ****************************************************************************
`ifndef __SVDOC__
  typedef virtual svt_ahb_master_if AHB_MASTER_IF;
`endif // __SVDOC__

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

`ifndef __SVDOC__
  /** Port interface */
  AHB_MASTER_IF master_if;
`endif

  /**
    @grouphdr ahb_generic_sys_config Generic configuration parameters
    This group contains generic attributes
    */

  /**
    @grouphdr ahb_master_slave_config Master and slave configuration
    This group contains attributes which are used to configure masters and slaves within the system
    */

  /**
    @grouphdr ahb_addr_map Address map
    This group contains attributes and methods which are used to configure address map
    */
   
   /**
   * Enumerated types that tells ERROR response handling policy for AHB Master.
   */
  typedef enum {
     CONTINUE_ON_ERROR = `SVT_AHB_CONFIGURATION_CONTINUE_ON_ERROR, /**< Master continues with the remaining transfers in a burst after receiving an ERROR response. This mode will not insert an IDLE during the second cycle of an ERROR response */
     CONTINUE_ON_ERROR_WITH_IDLE= `SVT_AHB_CONFIGURATION_CONTINUE_ON_ERROR_WITH_IDLE, /**< Master continues with the remaining transfers in a burst after receiving an ERROR response. This mode will insert an IDLE during the second cycle of an ERROR response.This mode is not yet supported */
     ABORT_ON_ERROR = `SVT_AHB_CONFIGURATION_ABORT_ON_ERROR, /**< Master will abort the burst after receiving an ERROR response. Master will not rebuild the transaction*/ 
     ABORT_ON_ERROR_WITH_REBUILD= `SVT_AHB_CONFIGURATION_ABORT_ON_ERROR_WITH_REBUILD /**< Master will abort the burst after receiving an ERROR response. Master will rebuild the transaction again from the beat which got an ERROR response.This mode is not yet supported*/
  } error_response_policy_enum;

  /** @cond PRIVATE */ 
  // This is made private due to known limitations. It should be made public once the STAR 9000993130 is fixed
  /** 
  *  Enumerated types that defines maximum address boundary limit for a given burst transfer.
  */
  typedef enum {
    ONE_KB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_1KB,
    TWO_KB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_2KB,
    FOUR_KB =            `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_4KB,
    EIGHT_KB =           `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_8KB,
    SIXTEEN_KB=          `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_16KB,
    THIRTY_TWO_KB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_32KB,
    SIXTY_FOUR_KB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_64KB,
    ONE_TWENTY_EIGHT_KB= `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_128KB,
    TWO_FIFTY_SIX_KB =   `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_256KB,
    FIVE_TWELVE_KB =     `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_512KB,
    
    ONE_MB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_1MB,
    TWO_MB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_2MB,
    FOUR_MB =            `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_4MB,
    EIGHT_MB =           `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_8MB,
    SIXTEEN_MB=          `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_16MB,
    THIRTY_TWO_MB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_32MB,
    SIXTY_FOUR_MB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_64MB,
    ONE_TWENTY_EIGHT_MB= `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_128MB,
    TWO_FIFTY_SIX_MB =   `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_256MB,
    FIVE_TWELVE_MB =     `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_512MB, 

    ONE_GB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_1GB,
    TWO_GB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_2GB,
    FOUR_GB =            `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_4GB
  } max_addr_boundary_limit_enum;

  /** @endcond */

`ifdef SVT_VMM_TECHNOLOGY  
   /**
    @grouphdr ahb_bus_sys_config Bus configuration
    This is not yet supported. <br>
    This group contains attributes which are used to configure bus within the system
    */
`else  
   /**
    @grouphdr ahb_bus_sys_config Bus configuration
    This group contains attributes which are used to configure bus within the system
    */
`endif  
  // ****************************************************************************
  // Public Data
  // ****************************************************************************

`ifndef __SVDOC__
  /** Modport providing the system view of the bus */
  AHB_IF ahb_if;
`endif

  /**
    * @groupname ahb_generic_sys_config
    * An id that is automatically assigned to this configuration based on the
    * instance number in the svt_ahb_system_configuration array in
    * svt_amba_system_configuration class.  Applicable when a system is created
    * using svt_amba_system_configuration and there are multiple ahb systems
    * This property is automaically set by VIP and must not be assigned by the
    * user.
    */ 
  int system_id = 0;

  /** 
    * @groupname ahb_clock
    * This parameter indicates whether a common clock should be used
    * for all the components in the system or not.
    * When set, a common clock supplied to the top level interface 
    * is used for all the masters, slaves and interconnect in 
    * the system. This mode is to be used if all components are
    * expected to run at the same frequency.
    * When not set, the user needs to supply a clock for each of the
    * port level interfaces. This mode is useful when some components
    * need to run at a different clock frequency from other
    * components in the system.
    */
  bit common_clock_mode = 1;

  /** 
    * @groupname reset
    * This parameter indicates whether a common reset should be used
    * for all the components in the system or not.
    * When set, a common reset supplied to the top level interface 
    * is used for all the masters, slaves and interconnect in 
    * the system. This mode is to be used if all components are
    * expected to use the same reset signal.
    * When not set, the user needs to supply a reset for each of the
    * port level interfaces. This mode is useful when some components
    * need to be reset at a different time from other
    * components in the system.
    */
  bit common_reset_mode = 1;
  
`ifdef SVT_VMM_TECHNOLOGY
  /**
   * Enables the Multi-Stream Scenario Generator
   * Configuration type: Static
   */
  bit ms_scenario_gen_enable = 0;

  /** 
   * The number of scenarios that the multi-stream generator should create.
   * Configuration type: Static
   */
  int stop_after_n_scenarios = -1;

  /** 
   * The number of instances that the multi-stream generators should create
   * Configuration type: Static
   */
  int stop_after_n_insts = -1;

  /** 
   * @groupname ahb_bus_sys_config
   * This is not yet supported. <br>
   * Determines if a VIP bus should be instantiated
   */
`else
  /** 
   * @groupname ahb_bus_sys_config
   * Determines if a VIP bus should be instantiated
   */
`endif
  bit use_bus = 0;


  /** @cond PRIVATE */ 
  // This is made private due to known limitations. It should be made public once the STAR 9000993130 is fixed
  /**
    * @groupname ahb_generic_sys_config 
    * Defines maximum address boundary limit for a given burst transfer in terms of 2's power.
    * Default value is ONE_KB=10 (here 10 indicates the 2's power ie 2^10=1024=1KB).User can define maximum value upto 4GB.
    * This feature is applicable to Active/Passive AHB Master and Slave Components 
    */
  max_addr_boundary_limit_enum max_addr_boundary_limit = ONE_KB;
  /** @endcond */

  /**
   * @groupname ahb_generic_sys_config
   * Enables system monitor
   */
  bit system_monitor_enable = 0;

  /**
    * @groupname ahb_generic_sys_config 
    * When set to '1', enables system level coverage.All covergroups enabled
    * by system_ahb_*_enable are created only if this bit is set.
    * Applicable if #system_monitor_enable=1
    * <b>type:</b> Static 
    */
  bit system_coverage_enable = 1;  

  /**
    * @groupname ahb_coverage_protocol_checks_system
    * Enables system level protocol checks coverage. 
    * <b>type:</b> Dynamic 
    */
  bit protocol_checks_coverage_enable= 0;

  /**
    * @groupname ahb_coverage_protocol_checks
    * When set to '1', enables coverage for system level positive protocol checks
    * When set to '1', enables positive protocol checks coverage.
    * When set to '0', enables negative protocol checks coverage.
    * <b>type:</b> Static 
    */
  bit pass_check_cov = 1;

  `ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to UVM_HIGH or below.
    */
  bit display_summary_report = 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to OVM_HIGH or below.
    */
  bit display_summary_report = 0;
`else
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to NOTE or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to DEBUG or below. 
    */
  bit display_summary_report = 0;
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of performance summary report of transactions by the system env
    *
    * When set, performance summary report of transactions are printed by the system env
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to UVM_HIGH or above.
    */
  bit display_perf_summary_report= 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of performance summary report of transactions by the system env
    *
    * When set, performance summary report of transactions are printed by the system env
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to OVM_HIGH or above.
    */
  bit display_perf_summary_report= 0;
`else
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of performance summary report of transactions by the system env 
    *
    * When set, performance summary report of transactions are printed by the system env 
    * when verbosity is set to NOTE or below.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to DEBUG or above. 
    */
  bit display_perf_summary_report= 0;
`endif
    
  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. When true, turns on the 
   * AHB Lite mode 
   * for AMBA AHB models. Lite mode has only one AHB Master and one or more AHB Slaves. 
   * It does not support SPLIT and RETRY.
  */
  bit ahb_lite = 0 ;

  /**
   * @groupname ahb_master_slave_config
   * When set to 1, enables AHB-3.0 features as per ARM IHI 0033A.
   * Applicable to Active and Passive Master and Slave
   * Configuration type: Static
  */
  bit ahb3 = 0 ;

  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. 
   * AHB Lite MultiLayer Mode for AMBA AHB models. 
   * AHB Lite Multilayer mode has multiple AHB Lite Master and one or more AHB Slaves.
   * When set to '1', will enable connection of more than one AHB Lite Master in a Single System Env.
  */
  bit ahb_lite_multilayer = 0 ;
  
  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. 
   * When set to '1', will enable AMBA 5 AHB protocol features as per ARM IHI ID102715
   * Applicable to Active and Passive Master and Slave
   * Configuration type: Static
  */
  bit ahb5 = 0 ;

  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. 
   * When set to '1', will consider / drive the BUSY cycle only with HREADY
   * being HIGH for AHB3 / AHB5 mode
   * Applicable to Active and Passive Master and Slave
   * Configuration type: Static
  */
  bit count_busy_only_during_hready_high = 0 ;

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** 
    * @groupname ahb_master_slave_config
    * Number of masters in the system 
    * - Min value: 1
    * - Max value: \`SVT_AHB_MAX_NUM_MASTERS
    * - Configuration type: Static 
    * .
    */
  rand int num_masters;

  /** 
    * @groupname ahb_master_slave_config
    * Number of slaves in the system 
    * - Min value: 1
    * - Max value: \`SVT_AHB_MAX_NUM_SLAVES
    * - Configuration type: Static
    * .
    */
  rand int num_slaves;

  /** 
    * @groupname ahb_master_slave_config
    * Array holding the configuration of all the masters in the system.
    * Size of the array is equal to svt_ahb_system_configuration::num_masters.
   */
  rand svt_ahb_master_configuration master_cfg[];

  /** 
    * @groupname ahb_master_slave_config
    * Array holding the configuration of all the slaves in the system.
    * Size of the array is equal to svt_ahb_system_configuration::num_slaves.
    */
  rand svt_ahb_slave_configuration slave_cfg[];

`ifdef SVT_VMM_TECHNOLOGY
   /** 
    * @groupname ahb_bus_sys_config
    * This is not yet supported. <br>
    * Holds configuration of the bus group in the system.
    */
`else
   /** 
    * @groupname ahb_bus_sys_config
    * Holds configuration of the bus ENV in the system.
    */
`endif  
  rand svt_ahb_bus_configuration bus_cfg;
 
  /**
    * @groupname ahb_addr_map
    * Address map for the slave components. This is used by system monitor for
    * performing system checks. This member is initialized through method
    * #set_addr_range.
    */
  svt_ahb_slave_addr_range slave_addr_ranges[];

   /**
    * @groupname ahb_addr_map
    * Enables mapping of two or more slaves to the same address range.  If two or more
    * slaves are mapped to the same address range through the set_addr_range
    * method and this bit is set, no warning is issued. Also, routing checks in
    * system monitor take into account the fact that a transaction initiated at
    * a master could be routed to any of these slaves.  A given address range
    * can be shared between multiple slaves, but the entire address range must
    * be shared. Note that this doesn't necessarily mean that the entire
    * address map of a slave needs to be shared with another slave. It only
    * means that an address range which lies within the address map of a slave
    * and which is shared with another slave, must be shared in its entirety
    * and not partially. This is possible because the set_addr_range method
    * allows the user to set multiple address ranges for the same slave. 
    * For example, consider two slaves S0 and S1, where S0's address map is
    * from 0-8K and S1's address map is from 4K-12K. The 4K-8K address range
    * overlaps between the two slaves.  The address map can be configured as
    * follows: <br>
    * set_addr_range(0,'h0,'h1000); //0-4K configured for slave 0 <br>
    * set_addr_range(0, 'h1001, 'h2000); //4K-8K configured for slave 0 <br>
    * set_addr_range(1, 'h1001, 'h2000); //4K-8K configured for slave 1 overlaps with slave 0 <br>
    * set_addr_range(1,'h20001, 'h3000); //8K-12K configured for slave 1. <br>
    *
    * Note that the VIP does not manage shared memory of slaves that have
    * overlapping addresses.  This needs to be managed by the testbench to
    * ensure that data integrity checks in the system monitor work correctly.
    * This can be done by passing the same instance of svt_mem from the
    * testbench to the slave agents that share memory. Refer to
    * tb_amba_svt_uvm_basic_sys example for usage. <br>
    *
    * If this bit is unset, a warning is issued when setting slaves with
    * overlapping addresses. In such a case, routing checks do not take into
    * account the fact that a transaction could be routed to any of these slaves
    * which may result in routing check failure. <br>
    *
    * Configuration type: Static 
    */
  rand bit allow_slaves_with_overlapping_addr = 0;

  /**
   * @groupname ahb_master_slave_config
   * Default value is 0.
   * Used by the AHB master, slave, and monitor interfaces. Used to disable HLOCK and HMASTLOCK
   * related checks when AHB locked transaction feature is not used in the design. When true,
   * HLOCK and HMASTLOCK related checks are disabled; when false, the checks are enabled.
   */
  bit disable_locked_transaction_support = 0;

  /**
   * @groupname ahb_master_slave_config
   * Default value is 1.
   * Used by the AHB master, slave, and monitor interfaces.  Sets bus endianness. When
   * false, the bus is treated as big endian; when true, the bus is treated as little
   * endian
   */
  rand bit little_endian = 1;

  /** 
    * @groupname ahb_generic_sys_config
    * Array of the masters that are participating in sequences to drive
    * transactions.   This property is used by virtual sequences to decide
    * which masters to drive traffic on.  An index in this array corresponds to
    * the index of the master in slave_cfg. A value of 1 indicates that the
    * master in that index is participating. A value of 0 indicates that the
    * master in that index is not participating. An empty array implies that
    * all masters are participating.
    */
   bit participating_masters[];

  /** 
   * @groupname ahb_generic_sys_config
   * Array of the slaves that are participating in sequences to drive
   * transactions.   This property is used by virtual sequences to decide
   * which slaves to drive traffic on.  An index in this array corresponds to
   * the index of the slave in slave_cfg. A value of 1 indicates that the
   * slave in that index is participating. A value of 0 indicates that the
   * slave in that index is not participating. An empty array implies that
   * all slaves are participating.
   */
   bit participating_slaves[];

  /**
   * @groupname ahb_generic_sys_config
   * Default value is 0.
   * Used by the AHB bus. Defines master number assigned as default master. <br>
   * The default master is granted the bus when none of the masters in the system
   * are requesting the access to the bus. Usually the bus master which is most 
   * likely to request the bus is made the default master.
   */
  rand int default_master = 0;

  
  /**
   * @groupname ahb_generic_sys_config
   * Default value is 0.
   * Used by the AHB bus. Master number assigned to be the dummy master. <br>
   * The Dummy Master is a built-in bus Master model that only performs IDLE
   * transfers. In the AHB Bus VIP, the Dummy Master is required. The Dummy 
   * Master is granted whenever there are no other Masters that can be granted 
   * to the System Bus. Following are the cases where the Arbiter must grant the 
   * System Bus to the Dummy Master: 
   * - When a Split response is given to a locked transfer 
   * - When a Split response is given and all other Masters have already been split
   * .
   * A Dummy master can also be the default master.
   */
  rand int dummy_master = 0;

  /**
   * @groupname ahb_generic_sys_config 
   * Defines the ERROR response handling policy for all the AHB Masters present
   * in the system, when svt_ahb_system_configuration::master_error_response_policy[]
   * is not programmed; that is when size of this array is zero. 
   * In such case, the setting of this attribute is applicable for all the masters. <br>
   * This configuration parameter supports the following values:
   * - ABORT_ON_ERROR (default) Abort transaction on receiving ERROR response.
   *   Master will not rebuild the transaction.
   * - CONTINUE_ON_ERROR Continues with the remaining transfers in a burst after 
   *   receiving an ERROR response. This mode will not insert an IDLE during the
   *   second cycle of an ERROR response.
   * .
   * This configuration parameter does not yet support the following values:
   * - CONTINUE_ON_ERROR_WITH_IDLE Continues with the remaining transfers in a 
   *   burst after receiving an ERROR response. This mode will insert an IDLE 
   *   during the second cycle of an ERROR response. 
   * - ABORT_ON_ERROR_WITH_REBUILD Abort the burst after receiving an ERROR 
   *   response. Master will rebuild the transaction again from the beat 
   *   which got an ERROR response.
   * .
   * Configuration Type: Static
   */
  rand error_response_policy_enum error_response_policy = ABORT_ON_ERROR;

  /**
   * @groupname ahb_generic_sys_config 
   * Defines the ERROR response handling policy for each of the AHB Masters present
   * in the system. <br>
   * Programming this array allows different masters in the system to have different
   * settings for error response policy. <br>
   * Note that when this array size is zero, the setting of
   * svt_ahb_system_configuration::error_response_policy will be used. <br>
   * Each element of this array supports the following settings:
   * - ABORT_ON_ERROR (default) Abort transaction on receiving ERROR response.
   *   Master will not rebuild the transaction.
   * - CONTINUE_ON_ERROR Continues with the remaining transfers in a burst after 
   *   receiving an ERROR response. This mode will not insert an IDLE during the
   *   second cycle of an ERROR response.
   * .
   * The following settings are not yet supported:
   * - CONTINUE_ON_ERROR_WITH_IDLE Continues with the remaining transfers in a 
   *   burst after receivin an ERROR response. This mode will insert an IDLE 
   *   during the second cycle of an ERROR response. 
   * - ABORT_ON_ERROR_WITH_REBUILD Abort the burst after receiving an ERROR 
   *   response. Master will rebuild the transaction again from the beat 
   *   which got an ERROR response.
   * .
   * Configuration Type: Static <br>
   * Usage: 
   * - Size the attribute to match to number of masters in the system:
   *   sys_cfg.master_error_response_policy = new[sys_cfg.num_masters];
   * - Program the error response policy settings for each of the masters:
   *   sys_cfg.master_error_response_policy[0] = svt_ahb_system_configuration::ABORT_ON_ERROR; <br>
   *   sys_cfg.master_error_response_policy[1] = svt_ahb_system_configuration::CONTINUE_ON_ERROR;
   * .
   * Note that this is used by master, slave and bus VIP components. So it is required
   * to program this attribute appropriately when different masters in the system needs
   * to have different error response policies. 
   * From slave VIP perspective, the indices of this array corresponds to hmaster signal 
   * value. For example, if the hmaster value is 8, slave VIP uses 
   * sys_cfg.master_error_response_policy[8] as the error response policy for transfers
   * with thi hmasner value. <br>
   * In cases where hmaster value does not correspond to  master index, this feature is 
   * not supported. In such case, user is expected to keep this array size as zero, and
   * program svt_ahb_system_configuration::error_response_policy.
   * 
   */
  error_response_policy_enum master_error_response_policy[];
   
  /**
   * @groupname ahb_generic_sys_config
   * Default value is -1.<br>
   * The Default Slave is selected when the address is not within any 
   * allocated region. For non-sequential and sequential transfers, 
   * the default slave provides a two-cycle ERROR response. For busy 
   * and idle transfers, the Default Slave provides a zero-wait state 
   * OKAY response.<br>
   * Used by the AHB System monitor:
   * - Set the default slave for the AHB system monitor (-1, 0 to 15). 
   * - The AHB system monitor will not perform the data integrity check
   *   for the transactions routed to default slave port.
   * - If set as -1:
   *   - The AHB System monitor assumes that the default slave 
   *     functionality is embedded within the bus DUT. 
   *   - The AHB system monitor will not perform slave address routing check
   *   on the default slave port.
   *   .
   * - If set to a value in the range 0 to 15:
   *   - The AHB system monitor will perform slave address routing check on
   *     the default slave port.
   *   .
   * .
   * Used by the AHB bus VIP:
   * - Sets the default Slave of the AHB system (0 to 15).
   * - Always the default slave functionality is embedded within the bus VIP.
   * - The AHB bus VIP does not sample any of the slave connected to the default
   *   slave port ID.
   * .
   */
  rand int default_slave = -1;
  
  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB System level check on Default Slave in the AHB System
    * - When set 1: Default Slave checks are turned on for default Slave.
    *   The default Slave may only respond to NSEQ or SEQ with an ERROR response.
    * - When not set (0), Default Slave checks are turned off.
    *   This is the default setting for this parameter.
    * .
    * <b>type:</b> Static
    */
  bit default_slave_resp_check = 0;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB System level check on Decoder in the AHB System
    * - When set 1: Decoder check for hsel to be asserted will be turned on.
    * - When not set (0), Decoder check for hsel to be asserted will be turned off.
    *   This is the default setting for this parameter.
    * .
    * <b>type:</b> Static
    */
  bit decoder_hsel_assert_check = 0;
  
  /**
   * Defines multiple slave select signal feature for each of AHB Slaves present in the system<b>
   * Programming this array for each of AHB Slaves present in the system to 1, will enable multiple HSEL signal<b>
   * By default, the multiple hsel signals are disabled for AHB BUS, Slave and Monitor Models.<b>
   * <b>type:</b> Static
   */
  bit multi_hsel_enable[];
  
  /**
   * Defines the width of AHB Slave Multiple HSEL signal for specific slave.
   * By default, HSEL signal width will be 1. User can control the width of HSEL signal for specific slave 
   * by setting this configuration parameter. 
   * This will enable the user to configure different widths for multiple HSEL signals of a particular Slave.
   * <b>type:</b> Static
   */
  int multi_hsel_width[];

   /** 
    * @groupname ahb_generic_sys_config
    * - When set to -1: There is no limit on the number of rebuild 
    *   attempts on RETRY response for a given transaction. 
    * - Default value: -1
    * - When set to a value greater than -1: Defines the maximum 
    *   number of rebuild attempts on RETRY response for a given 
    *   transaction. Once the number of RETRY responses on a given 
    *   transaction reaches this value, the transaction will be aborted.
    *   - svt_ahb_transaction::status is set to svt_ahb_transaction::ABORTED
    *   - svt_ahb_transaction::response_type is set to svt_ahb_transaction::RETRY
    *   - The info of RETRY responses received on the transaction can be 
    *     retrived by calling the method on the transaction object-- 
    *     svt_ahb_transaction::get_retry_response_info()
    *   .
    * - Max value: \`SVT_AHB_MAX_REBUILD_ATTEMPTS_ON_RETRY_RESP. This is user re-definable.
    * - Valid range: -1 to \`SVT_AHB_MAX_NUM_REBUILD_ATTEMPTS_ON_RETRY_RESP
    * - Configuration type: Static 
    * - Applicable to master and slave agents in both active & passive mode
    * .
    */
  rand int max_num_rebuild_attempts_on_retry_resp = -1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to check that the bus grant is 
    * given to all the master connected on the bus.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_all_masters_grant_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to check that all Masters have 
    * requested for the bus at least once.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_all_masters_busreq_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to verify which master is requesting
    * the bus and which master is getting the access of bus.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_cross_all_masters_busreq_grant_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to verify all the slaves have been 
    * selected at least once.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_all_slaves_selected_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to verify all the slaves have been 
    * selected at least once.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_slaves_selection_sequence_enable = 1;  
 
  /**
   * @groupname ahb_addr_map
   * Enables complex address mapping capabilities.
   * 
   * When this feature is enabled then the get_dest_slave_addr_from_global_addr(),
   * get_dest_global_addr_from_master_addr(), and get_slave_addr_range() methods
   * must be used to define the memory map for this AHB system.
   * 
   * When this feature is disabled then the set_addr_range and translate_address()
   * methods must be used to define the memory map for this AHB system.
   */
  bit enable_complex_memory_map = 0;

  /** @cond PRIVATE */  

`ifdef QUESTA
  /**
   * This workaround was put in place because Questa could not solve the nested
   * foreach loop constraint that is in reasonable_data_width (out of memory errors).
   */
  rand int questa_data_width;

  /**
   * This workaround was put in place because Questa could not solve the nested
   * foreach loop constraint that is in reasonable_data_width (out of memory errors).
   */
  rand int questa_log_base_2_data_width;
`endif

  /**
   * This workaround was put in place because INCISIV is unable to resolve the 
   * hierarchical access to field “num_bus_masters” through bus_cfg in the right
   * side of constraint.
   */
  rand int num_bus_masters;
  /**
   * This workaround was put in place because INCISIV is unable to resolve the 
   * hierarchical access to field “num_bus_slaves" through bus_cfg in the right
   * side of constraint.
   */
  rand int num_bus_slaves;

    /**
    * @groupname ahb_generic_sys_config
    * This variable specifies maximum address boundary limit for a burst transfer
    */
  int burst_boundary_limit = 'b1 << ONE_KB;

  /**
    * @groupname ahb_generic_sys_config
    * This variable is used for checking address boundary based on configured max_addr_boundary_limit.
    * Default value is 'b0011_1111_1111, which selects LSB 10 bits of addr ie addr[9:0] when ANDED with addr
    */
  bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] addr_sel_bits = 'b0011_1111_1111;
  

  /** @endcond */

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2f9CaoTY4+S5eBDUbBEODq9sLyDn4cuutyMcgHlevE5n98GudIm91PPf1I+ltvvW
YnGAD8eGAU3JM3UQdRUbdtFDlK4dNzhXHatI7KVfO6T+LZm7A3OsTgIrv60h5v76
Vab6TTEFDks2DYfr/gPptFwch3cRcxcCDhccWxvNTfYXBCtIyUZ31g==
//pragma protect end_key_block
//pragma protect digest_block
i5YLX2+SQE9cqdmivEvYaN1fTFk=
//pragma protect end_digest_block
//pragma protect data_block
HekrAEBCG+K8zbfE9pujJ5j1OHsB1x546iVnL2NkCmGdrolP0JQhdfQ6uAJBpaM+
96dwQ31SAz4JPrq/kcxElMNlHP5VRV/kWKyCxWeHhSot9Wq4r2CaetI9WykKkWgH
Q0jTTXibiJJsfPqRvRbTItsF5/rno7IF00Tvl2yR1DyhuHVIf0fvAWJyFozArmwv
n8rirrcPxcw/Yr3xGqG3VEKcmdChiyIPIhvGCPIprliBUggOuKYE0qE1AG13dyHD
838yU6Fy2BL2M4/Xnuaoh/D3SdkteYMBk6asWoNDe7sJ7CX+AvjRQthmivpXGxe3
JBnaDK/O2dnDg90Xdh6phEcTfQGu0fjqoI0lTEniCMkYPxbdO68utuE8Aw8lQU2H
xu+OX97qAUDrB1HRbdX0Zgt+svKlODJTYtewUdtZv8lspP2PdI5FEF/9a24qBaqx
UbbWR3j6KjshSxz0RKEBvG7igdDeJ4hoEqTaNVYJkut9xD8KgwUfHhYVTXVT/t6y
l64k3+4dKN38lIh5GdMKx6bHAgqvFro4GlHH3+d2QqovLR9w6b4hizloZ+JKNdvE
yeUQcEWwSePqUw2h5lBNimXCtNoKSvJWxISJ8LEwVJWiT5jZSYTo+iqMAn0Vdk8r
lX1RQERl8TH8eonRc8SBQE2ZY09lpZPl4r+CinIsS/SBlhZYOU6/Q+NrRoTBgWAm
gxYSK5qlJ9gawKFeox5nG4EBBX/QEAzkFQJzovDTMPXUN5JE6amRMhtym41RKhMP
So2i7vyqDUDqP7fCgttiinFE862VNbJId9p3UnB7Y9eOjA9v9PTohYAlw5ibAyk8
Ng1ZxMscslJG6lI1mw5q98OZKq8lQ3Rw1c+TNoMwXHdKumZ2AdCmSWd7a9Fh8YRh
rfNY0ZhZy7Kmnwk6TfTEP9ZJFfcuUaCpqgzk3I6i05P5cy2q9BeogU+7egGgAqOw
UVA+5U8sm5NAfNzP/6GnuWwFlFEP4nehJbc4JrSS1JAT6siXguJa8FLElSSr7SWr
18dpg1d86F+ia8Nju0Iv1hg5M5HWQyjHq/4MdYTifa/VH1BCO3Scjz+LkF0lY8qy
231VYPH8Nl4tBhGgFJfaEI+L55Aj2LqG+RaZjr4T1PJtRMdw4uWffzdg2QfUFube
snSs7YyVcWddG2taY+B76GxMkh3GYTuoRWavHDVYlrph8lQT2pZGK8R9tLUoZmr2
awaUE4gmEYhie5eEJJWFQVFckC9Y1pX8scasCmbSW2qXr1IWSWhtzrJmW0W30a9M
xbyYoKLnzJ3/aCBUDjuSAFV1iBHxyMeHpy9ulRHCS5Nex8xrxr5oAsx8Bl46Aeq/
TyYTz36KFG8gnLWiun6m70LwWxCjlJJf/vyn1nqObMzM+jSv+h993XqbLPLFDqxz
r379Gc3xCJuLKCujk8hUTQLDzaqSGrw6igPozs60PCQBzSPBjYAEJGJek5aF8aqT
GgfICqYkNGptf0z4Ix82ty8U5ttV/hb4E0FFhhHY8HhmU0eBcgdmYG3qhiuLEDSl
86XWtMKo4dHsh8HIQaWxMJGDSMe+a7g0/qAIozZ/oZ4aUh7zaTYInrWU5ZAYV6xa
MEp1tNfDBt03TRzLevBuxCj7RkQ1vrt/6gaPrI655vxHWs07QiAOXPd2josDHsUo
iMWbfiad23nLkFn5nLAB8LA7uw5E8fOmeweI0+y8uJ+gi2+WMfqmv/xVnWu6gkyu
pa9JfHg3ekNgceKoesXfjXwWze0lbUaFYB3MWvLqK0qkEEZrYjlnh36c+ERwm8ex
YKxw/EYsT2ngGil1gU1etsHOlYp0OY8D//oKoRW7erUDF4JUwBdBEkb74uaAMXzf
LcQNFdLtiTiYzYh/asYXoCkl6jd40qVFzubPjy5mQgUFNSvGToUXUHxnFYXUNcyC
yRrpXurgfdZ7Z5WdhWvih2WZTAwuTcxXfd5h4kgKUWTuzI158jsRk1RQY4wpFqGT
hMFmFYmf56dK6QRxmxn/F7LHtcdDs5iBa2VtAm40lTvpHQXSRHXGzbzCV8JOD/EX
IT9cF1Pf77TXwseYdvAJGtD+x1By+UG1xRCfRdT4I/w6ajJ0l/ZKKJl20bwdQl2Z
bH+Pz3EANYAPmPjT/kLS9OGfSdhB1PV5+HLLXDZKOptkUGtbrPy9IV7GmOpkzfnz
uH2kSKrJzkmMCju3g+CvGddCmgem8FGtf6tmqNZgHCbXsKkSaNWmrHuIZDHHTudj
PX7CHW5pfe6d0YkF7DFyRsBrVGmhAGnad+EDgupxxuQcEAdJxi4zpyPxEmUV0vXK
dStmYLMD5n7tPZ8vaWV46NB430SCnsiYN0iGA2VZjNtVeon/jezOk63B+VRSi4fk
w8XV4L8ShFlrpfDuHZDV2f4R82OLjw9PH5detE5lPxlZ24c/+q1gisF7AMwyCvE/
CT7ftnP8+s2UtaRZh1U/sSJqyB3FWKmDGz6T4Fl4HxQLgIrABz5//h5ZD9OsV2Kc
xH4qxLYFCXoW1bosjRgSOC21o7Bbf8isptnEC3s8Ma6WI6F1OcXMNYT3yOB4EHp8
YSRYiMgxFgB8s1NBqQBG6ADgu79NgtSkZKch2rkCNW7BsZvX8y7126c2g4DgSeq/
/wd//0a0Pz3BgQRZ1FWAWz0GQfVoLDJjxT1+LDc/do5rVqJr99/BBcJhvrVyBa/g
oFTqMsJJtMXJkDNKWMGpkQfdpQxMVLX/Lb/knWo1zSNprl3azpv2t5F7luvzGVzt
0HOPU6IMA2QvHhmp+jwwaCkcxaHe6ik7vFlj96ucMihrBbMiCme1lC8s6gvi6Xfx
HfqpO36c0WcjLiFTvmUfg/orzvJGyzrCL5oPSWxcb5PXafFMrlNiY0y6247L5Kz+
8zt3zyhhAnygnnzxXA9naa816wRza/wk5YFsCz+wvfLMnYAsRLbBKSUIpjNm4P04
YNBw62uL2CdEqreFTkr1Id5BLWufL686XZWf1lCSrt0fTGMynYpTszG4uTKp5gM+
C/UYVOsLZKskMs5cV9N+pjwLu6WiP0FumdxmI4RToYpe/8/r5ePA18GqToX6ehKQ
KzBkvg1ZK0hI1R/Rqs2DyIeqGsGksheckGuXBsjK/GL5JxBFWZ2XuwFaSTZEx0+V
J7yLGgPvjCp00mzzpUjjHXTKzq0RDmkHhsGbtwC5f68Jz472b3wzZiVR56jrnteR
eJ4HxVV9zBAs+cpDJup7yUsobGVwfCuHa9Obs3b0s/vvdOuF7mT/gtS+goT8Qntj
4gKob+wV0Xfs2ys1m6JZC4fyKmfVhT8Vh8Zz96WNXI3cRJIG+z8ga+WXJwNdQKyk
dJEIUtiU97eGOk3tsIA/BQcn5vX3vZfAvik1hsvP3B+R/EMbzBg73XU3EibsyDNK
iDdKTc0yajSCx0mKiqP9WNJnV29N+zlgLLV2bFZ6570gs05Y3ctQcWkIH5x9qgIk
YwhQrEnoKrFi26TtrLz0MI9+UtbbZ0Avv0KrGZ2FG1pHs9P4pTS6TKYOY+t4nJ2n
DFrxgpkCQ0k0WURf63RgfLWVfzOqC0MoeMnfxJ2TQYKrS46Nz8K6vHE66jHhKkOl
YGhy5QOpLmAqKlv1d5u3QbtqKW74UvtiTsqQVoDrNiwfAMdTcRn7Zg3de/hw9/qu
W25Q2lGt5f1zk6+S42wm30FFgOIHhbX0VimHIzsl4nijx8K3yu1Q3ObcoLSzppsW
uw/Kbwju4M/ZWPVJvF4AuVWcQmhWH8/HAldcMWWa8VBtGf3/VmMa2DmRly0HRLHO
x4zmMZ4GZX109DMr6a1AO6moHg7BwItASz3PTKMGVJwSbFe49H7lVRmsTXdTtrIe
HA0uZOC5tPLvwTx4QEy4BcWCb9w2N43mBQJGsKz4CYgaeFIaU7lIF+F5EOoblQ2G
dsMshrJwlRfQkBucHnNqgNNaID1Xs0TSF0iPIFZJ5Z6OQtq6eBTexp0p+6Nz1JCc
gOraN4qri07dAWoX+qyI30EH0q2EDJCyahKrFf5xu28tdQkevrk+Mqsjkps5jUJX
IBnpSuvLGpUePBVqeMNExvtfAy1QxAxE/7+npkeFE0FhPuFAg52O6zdX4TcCD2uO
AB9Qjg1j1HEdKZONN+SKk6KYkTI7uc21aHRl+oP1xXyeq9jIj9dlhISUZfQ1H4V5
tjXjs7QiRgfdHt1IUeJspI9a3zgkXbO4TNmFuGil8UYKM+KY1zUjuRsFvBHqz/0H
h960FOYyRGFdLQMy11TxYgRFFwg3ouFNfEct2MM8zZWmft+hUoS+OuTBYB9/VjVw
+X0YM6pUgbg+ZUsz8AymleGm3W3rDlwsQz2bSs8SBgk+99FLGZIzxILobjO0MOz9
IzSxo6YlTbS+OWQa74tUl3grucOT2TOVvzv9MD2aMtbw24TpTT+oH91Zdqks/VPz
XDJ+WCEisjNFChl17y2UIz06Xk0KSOZv7XZNSAFXgVYn9UC8/+DF/VkhAdQdSeCK
1ERRWUiCmiA7HYuutDgwVi7yVHJu694QHj2w+PF4kZm4kDQSrfIkM6lEmkXiM8uc
ZTs09jJDc+ixIB4EGQKqc5VOIkZEygZdTO1N3H0prO54fYSQ6nkJt40Ji57m4hND
M9jo7lVISD63LsrT+Di7VzBEaImUQl0eyiC3AXfLongPweRRASaf62BLonr1Pg5a
DQogufGVBqFjg3ZlsQvurvPvfsR2tOVgDxeJ/WKxBC6yzaxUsm2ja3wKn1fQUWwJ
O9VUZEyvDPWxJkQKnwWZMlLBiXuuxmUO6/pch8IyiAi6F3RhiztjEegjYPiQE+Uk
rBuLgp1AQeFpTX+MHx1PtkIKSAh27ri4CheQDctn48iyTrtFC0wB3TH1RRIcJhwT
VwVJ3PNwNFuG4TH7AIWisJMKFOr8WnQu+vb26E9UE/jy9XeI07Ev/gBkPySYBItq
PPhP28DPq5UHfGyHVeHBMQYDi3D01eB5obBB5AR1lMMUXGDaHQGs7FPW6dlaNJKP
+rPOSjhHxzF0UnDzfv18Qrufi1yWJNd2VHrOuBW1xCO4KwwK8LlZ2Kw+4lTpFiHN
T14pg4WZsfAJBeP/e54WN9krA+8ADlwQj07FWNZM3dv4iQeE6g9+Rk0qNetkavhi
xjoJb9aX62ys0ojK9EgT4verkkgvCGVb0LZfrbmkC3jchPgPt5f3sbCgHT5mrKK/
RU8+5mvrCaZe6LvPqUllRkC30X7VcOfmjH9a62NH4DouPlke2mtZn0/dFm6n6PBy
tGzwINjZ6UMnQ/PtB80EhoiQ1bD9XXFjGNeakYMOUcKE1EaDGklfXiH5QyDnaqwt
me6x2EwVsXI0JH5UaYB1z8TtA3Z9Uhh6sQ6iQHaLhf0/JYVFlY12Y1YrYJRYnYxZ
ENQsDliI9M1tg4arremc4mPpl3Hnq0WkRP0l8OnuasOkW2ACiHZ0F6YRTDQ6Gabv
GXM8YMIXyu6ed8gQePxlsa+rLCRZKcNSeYlZE/6KvdqbhFO+fAnkZfB5N1AHXe1J
tnI63DxmV4nwAzJCNVNsLLc5YtJm6ZonARv2H9hdGItljKkOWzpXQxiP+VFSnMGu
UmPqf3oG8GHb7R/UtqqFVMvFbf09nHFs1aIfMEDzp5UeB7+R9rNHSsWisLMf2oH8
z5wsK5VAqGA/PPdeSuaG9EiQf3IzWVrJ/gv5LpTOlxsozfbUuKsD6c3sD99z4Swz
0wjvoIJJglKpK+T8p8X1HDCFJ+RGiovRYGdiukd/G5od/hWssTs6lOVwQUC/OsSN
oND+iSU47UmAWCunLopXyFVTddpAuYMsPNqX1c7cEoLlBRldG8djIWiy/tcc+z7y
62KofvC28IfVfaIHiqGW31vCIzN+LRGvXOzIDim7thXdU3cyTwijI28Ys+prgQzP
knCIYrdmRBtH3TBiy3qWrJGu6jPzRS4dMfdUtJiLByTl1qZ7uAdsmU4VHUTZHTbq
V727qas6vsE9/N7RO2bF4UIphRXF80JofBpqvroNDLPOfALk6ummfl0lZ5rb/vem
ZMiCl1g+OrHl7Ik+Xy4wK9YD8X89HMDOZCyu9hgS2ajGzyjhnMyxzVnzjPyC8NjA
1lHgPPpv7MFYTEVYfyTI+gOXBMJSeCRC888A4WbvI6ZxlcuENX0jfTL/kylx9He/
KlOwfRlDvTajI2g+LZvJkULjdAnNMKMb4lqpBcrTyHP+uHh7fHzGntNXnfTZn1Lu
GEqFXvv3AShPcGl0Y7Omju/w0Z6qg9CDIaECafGRhEftFw0D1uV/ue161/ZE3l+3
j4Iv0Z5Jq5DUQt5Q0iMwUo68R96C7uFfK42a19Z0sKokVHvW2C76b4ZaEGML+nmq
HtyDTPM80dP7/zTFMTV8LLgrW1I++ax8830nNjdh1ow6Q57HipTBLdCQ5BME4KIs
Mf6JQFbodM+o30CG8yVm3kmjgFYR6kY+fCDYw+P4niMjyLfYrxzQX2wwv9GxH3V9
gafG31DmEbDz4JVMhzbMRHmgAcFe1Cq8BBqRObFgYsJiwZBrym8QtxywTBOdwEGa
/tG1CFC//DBelNUdzwL5vtgBuZsMFdMf021pdtqqmMiGYsVmy1/GNaAR1tbNhnr7
/nOwTFFzoQB16M9S+GnNWBZEt0t20446s1JaxoahbUgUKgc9gssIeokwpe96RT41
YP12e9cHh3UzcjSgMVM6XSI6A63Vx1U8Xl8O7ZK1AIpTIzAzrO3xhoRQE3f6jQBQ
YPGdwzhEb5/cykKwPYsWeST0pkg5ncXrve8pweG4Bsz0u6SwoYx5v1rgCIqGYwCO
11qMri/aW2E8fdDJnK7Xwil8IcSwv/uFM449L0JnWetCUflzTwRBQyxnsVvB3/ID
T+G8tWAZTavBJpZh8U9h6zmnc9Sr9PIKsUDYg9yZNCTxE4wpIRfSaMKuLsrAxPL2
KIOolcZhSIoim15tCypGDLyZ+xydVrcGXG9S1Iu5X0GkW7J0b3DjLJ4iPBtelmP5
v2v0zotWl+jrrb0e+wNJhAD/KJ4x+RJLeeORAq2zEyTR7NY/9PigV35tWtDN0MQh
AfcOYYKxx0T6oWokxgB/cvirTf+QJix8GzbC+OgCqByYAuSqvVMgLpz8H/8nvzHy
KdxqgePIOj88SBPONRzVtkPaX2rlJI5Q3aNhm9J7n+I2Wj6p92BuwuAVFlnvQbNF
4ZOXeopzZuhwdQc9716ikd/3e4d4IoC3SM0wIL17ZlMNRKZnNbNYte8vFtkQkM89
MBGInikGo5s6XCC1zHMEF1lN9FF7FVmQDopulaHMx3KixihBAin84fE+VjS/cDUo
JsYlmdHfMNVl4gkVFGudlJbWi7eQiw7DJXxQOGGvhpPKB0EGLATIzDXaRerbeKpR
cmpg5s0JURkV9bgcuYuQHlmIrt0hMK64kgCaKFLHuFDEqRpqXmsX8s5Ro14w0beT
lxItYTNDnV9hjGnzrs/cYBh9dtpL9hcH5vO1rWdfRVttz1U2y1X4ibwR1JMSXvcF
ur6yXkxOMC6f89jjwiG0bvUZPKL5Cbl8NPN+SQPlsNx0EKFX8BmPMwvPRlYrJ9IG
7QKARfwMJ2fRebqV2RmcG+Vl4BYXR5TzcJ6cVI1o5LnTaIQxv94lxWajxZ+mtFfZ
+UEBi5nPSuFYlkxdXUzj+cVzg1UGJXt1tFReY3XVhkkxSwNEypcko3jS8gqq1v8a
stvBlxnUVXxDM6chk0ImXjjSISqp9avunipQd7KmyhU9DH8lbLMBg7oAZ0qZo08h
jEk9X+o6pcHzy9mK95g3NlbKPRBVSc0R/UEUbLSmLJ+2P+cZPtmDo/HPKTfKRp6M
CjLAiBg3TDY0rklIfHMpnLsUbmyCMs/yzNwy26rRT3mmrZK6E8YRE3GkThWFDDmG
BoOSks2V2QzWnaObm8CUYozKeRsj2/StmBTEYoYcnc81iOjgbRUH6xzYuFP0+cfr
UHDQMtc7k10ejdQH2G2jPrZPoKPt9WJwAtfABZE0iaZzNbIrPFc1rbYuGe19LKzS
BTPiKIZXVxEIBsD3AiGRrmVTeCUstSMNtoYk3Kh9XACjygLkJiLv58IWAf6pGsES
5NL2euK8NyAk7SO0ga3aMGoSIpZE/fkszdZ7Xrmt0nCdHO5QiSLTCWBo3jqOcbes
9uKA4ozMPWOuTjyRsXRcEo7ctvcy4tFGRsvd9hn4i4ABWhX8sNA+PdBE+hqqlthF
/JyrPo8SDUm7Qmj8bI8kXzreeJOIHZ6GbiBizrpXvbJA0Yx/ypdpUDplBNE7upen
mhHd2lUAKXMITm5dBEu4HfU/Uc4Rm5Co5GUY0sPDADDKD+tVZCTOT8URSJdWLHpN
jCBvEroMonYOFAthMC0Rreca9fjElkB4ccjcVR5MMiPY3jrizc8uqpwJpoZfxY+z
FKIpOKlWuuz3kdLNmKXoh+5hruunseYO1amq8hJnz5AkWVEKi8gbS5Jjy6xIr7FK
mCZt9EK9lF/ROLGqoyQPams45FQvzY0u3+3cDWGs870L/abb1SLgFNsjkp24M7+K
gp4mkyZJDJd7ff5lRdjiVAuMY3oV01rjCBgnCTtycnU6OXhljcZWjqEmRetueRXl
vwrLbDCY7RfaimL48Juq3zoNMnRiPZL5EW8LY6HWof2T3yzDWH5ZLZ+yo9O1K9ck
oN7kS/A4ADMuVCH2vkcbrV8Sh6Qto6VuT4pn49PfEExQ8dP6+mQqCBBT1K4HgJF/
Ak2Z+m9mMozzmG9C+8zCCphsOYoZ+VFSFxZSGVJtkQDyJltQXli2fYg9YXfN8fw8
8XZ3ImwJM4rnegdM/39qVdVrCqoALsGXMHyUQf7rG1S32o0y9OepkNExjULsL5bR
Pc3Gp2nvvd8fEjBT3QRctWhegYfFM9ctM8nE6QSwwjFGy1QTBeNYxKhuot1oc2xE
M1cX5Ag2fwXJ80oJCkLqnYW9vepPOyNq3YCPkLop3QtrEvYO2DGaHJSsf9l3jmib
uDzM8p2uNUTdVXKWQ+Mdy0E82tLnS833AZ7nmB40gUshEGUw3jpv1I9oaEkFhv8a
OcbjyvsnWeDRYraXaDzsDB6kuJdSilC9/OnayKdkZrz9QT8z4COUujUixQfLm3WN
7P29ndN7VAEiVug27OyhNcncJDpO8KGsP5d4dmlccvHZsJGGJb1DjfFXPdOKaHBi
waSfxH9Z7uvFGp2U4Or2ZfN9OBhWUrd0QbkCoPo8s2N521B0Zdl+uC2ftQcLP0Xx
52fkG1/f0ufrBlEiM4GQ1I+I/5LyX3tqdvJ5xkSQ46xgTS03wnUukA83vp/bQ5SU
0NPeAgy4nqUrt73riW7nItRZpnT0dyfPpogqTVTsWwxjJ3KIkk8DQcwRak2dlP+h
EK5Yd/TbOJUMc3TO7oe+ivfvcTTIGxKYvDgJEBAAKDL8rLjfXf8EDEkhkZKudBzZ
ncROkhCcI9CFCM16XHV3res5FMD0/nZFhf1wRZwCsT+IBSDmBwSZnRlEpgQ0NZPq
yyQr0dINDE/4EowBmvcEm65I5nImEbXzPr9q9iJM+DGacLLHp8LZV/bg/F6H/ENt
JNwd4AmgGOKssY80MCjKRHgjk+73Lt1/Bqs4LJzwTa6V8/GX+hHWp7yFpFqrCeTP
BOoekzGLB+opCUf7pDGh+S8fu3Y+AUujBddi6COlWtAe8W4luXPptrx7lJJjOM5h
N3yp4XoYgG5CBA84vezH4JIHVDPcgOozHok5ioXYBEp/BZhfP+fhM3PzzfKN1ek7
QqqdQjakkTjlUTF83EcW082HWGbhjrXSQXorxa6AlUfnGOMoVdmJYfwv+v6vnWT+
99LbI6oD+o77hx44rIWIvRXbK55reoG8WsY2GJTkxSebRoAExIC2r8w2zCMwVx+2
Pmucbaawc1DPZ4Ql3wWsUmzl7/A9g9hj+o58b3tTm85L56N363c1cmnCeFk8jdpQ
36L93YyyEVsh4cU6jqTgDhudoiKAG7ABkpB16Pk4hEXG4D94RdZH72M6DcgwDSre
Z4nmIjNuKGE0K1h3I9AGZ8yJr7U+hlVAyAR4iY0IwxwR3Grun1PZSHj5A5qL9WyM
dQ9ZNkyC0+v75lxP2OjOCc6ZTWzhc8RJcK3wjp17aLQjs17pEcwqe7GqroZoMCuo
w0fpsJxHV1EuWy8ZR+XZc2+trkPdt8dRpyNFSfETrn1altUD/S6hd4wtJ111cvsH
ts688XiztBvh7QVDftxuy/6C2/n9eOSZzghqUWgIE18yhTlj/yIqMvlk3j1o2kE/
F8nCPyOwquykIkSG5cDIyTPL/hZzOxKTJ4QDBBT0ZJ4BrqaU2+9dAPzRlg6IEPAy
d6csL6MZL0ToxwnXTetzSadbh3G9tBZVNwjJ9Oxi8D6QxbAtlIdXSqgWEISqSBpr
sUdDpcQiumY+s5pRSUrrezFa7YzOgQ3o9yPKxgAnJjKr1tGtVRgvQORha229x5xB
dGfjcS120GctaxUuQziJJbdFbf+5TIj5SeaFSjRtCdHNxq8+6rWXaO7k49IeELQm
Ifm4wVPKIoxzYL9KeWAh9crDKKqAe8QfciX/i3VkImx0Iu4XNJm9p62D0b6625q1
jKM3vl4zYeCVETy/VR+vv2xcXofrTRNzYz70PXlzEiKLNq24iHeFwK0tAeE2AXSO
x0yS6nAIY86t8/j9356bG7vnpNMEnt+7ov5163GX901dRiCl5VF9uxQ+AtXsh3lo
xDPr/FU/T9XWFnLY09oaaV2ZO9sYunQc1NFJYv7N+oCm96/MKwnQUx/K4DrOV4Yi
XCsIbRx2a7+t3U2s9RpeNMgN76rvYJPmJfgDGXwPnrd2mrscJmWIkuDL2h6yhxzs
zH3xVXuD37piN4GyM5+45GwByxv8eloj8yHcSZd6b4Qoy1VzvOEwsdJWySwhO0j0
s40CBsTkx+/t6em0qJ+qeHiWDpMpV9LHxjXD3lDHkNbIeeQ/sP0n0+nluUG50Vpw
MYSaSOZZpLn/BEbm7U1Kvk7tQ0b/BmrPwDQ0Vgsk+nVEmV8gW9QCF1bRk7bN8wB+
gi8ntWUNgjvn5IT+Mfss5If53EtGiL5n/yh+i/tW086cuitBclWEDlmYMj7abfOi
0oMqmzSITUh4FF9wtEmZ0U+/tHvA3IXHArvBPdZUS+wOHdwBYa4JkcV4BAysMEbc
9JNjCVTNbPDyDLytEG2EWRV/MF3TCNBCF1ErOd6vn+XINxsMKKp2Y3JH7eB2jFcE
V1NizurrA+FHOq5V01s6SUEEI11gPvmdb1lRDbq6b9uqltngqH+0RKl9OMikyOai
z772OnFThACmS65M/6JbGAM9sRPO/3gJj1T/VYGdPniP9hpgpmR6jIeI+CdczIz4
MaJzzPFeD6jCr/8jkwj3ThAmTU66iOIaN03dWSHuoEsbJ/CxSYrFx0QYFWZCENH+
tVvZTvsBuSkHRU+loizeoqPRHOhCvNRiBQf9M2b58H0UPsIm8cLaVWUEpUZsnLHC
OZ0bmHGaUxUY3Bld0oZXsV/BGyLQegPp2cZ6YcJtsUh9QCUQhrCE7FyHVnxOdi9R
UEGgC3rvZgcFRS5oXYNQtw3z1FFQKtw6NdzzrI6YpbylJCQpkyv46OHCWYsSoyq9
Ue5YA5XKYXyHPIPXVfaHkyOsXMPJ35FGPzwv6JOM5rrdBNO6t5OznNgcwQt6YoxM
sFJ8Ogn+NfGXb/V8a+rKXEd4nD2bXq6CV8Kyeam/7f1kP90CK2NSvQTmwNephvDY
DbI96sjFCC7MvodkXSI/Jw0HLjdKcfpC45/QMHZJsUGddOiH2aMCIChnGQKbR5BH
RSNECFO9fU73Z6Z6V23ClYMt3TlW9bkkroF9bWt188kBY+PesIe+9o+elp0/TFRA
BKcn3ZXxTMOARBScs/3QTU7+nHPXAIV170hulTJ32gU504kqKmojCml9Pex8CU2c
irCMMKqlvqPBCSr+rO4LGwnSW+dWW0NbCn13LWal9aI+7Bu/S46wgJZd/zLsVRR+
EqNiBE1LbJzpyX/npH2Yi4x28WqivDzcOm4HZ66HzY1UWCkgv4w9HybZ6lCOy/fd
hx04dqIPXUQFw4ApFFPt6g9qLEE0R9SsjOPCkeRevyhK/iCWYZjxfDIRDnCEgxWo
zS/HLP9tdN03v4NkIBRQQGLX6m0NPcTnMIVNu++6K468SeG0W7tV6Wcdfo57rhX5
UFsGc0Vq7W3mD8NMM4yF/9VNMlgJRJvxu41vIEaEhEI=
//pragma protect end_data_block
//pragma protect digest_block
LUNQCDY7f+sMc0DfnpduNnrd4x8=
//pragma protect end_digest_block
//pragma protect end_protected

  //----------------------------------------------------------------------------
`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_ahb_system_configuration);
  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   */
   extern function new (vmm_log log = null, AHB_IF ahb_if=null);
`else
  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the configuration
   */
   extern function new (string name = "svt_ahb_system_configuration",AHB_IF ahb_if=null);
`endif

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following:
   * 1) Allocate master and slave configuration object arrays
   */
  extern function void pre_randomize ();

  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_ahb_system_configuration)
    `svt_field_object(bus_cfg,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int(system_id, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(common_clock_mode, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(common_reset_mode, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
  `ifdef SVT_VMM_TECHNOLOGY
    `svt_field_int(ms_scenario_gen_enable, `SVT_ALL_ON|`SVT_NOCOPY|`SVT_BIN)
    `svt_field_int(stop_after_n_scenarios, `SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
    `svt_field_int(stop_after_n_insts, `SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
  `endif
    `svt_field_int(num_masters, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_slaves, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_int (participating_masters, `SVT_NOCOPY|`SVT_HEX|`SVT_ALL_ON)
    `svt_field_array_int (participating_slaves, `SVT_NOCOPY|`SVT_HEX|`SVT_ALL_ON)

    `svt_field_int(use_bus, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb3, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb5, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(count_busy_only_during_hready_high, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb_lite, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb_lite_multilayer, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(allow_slaves_with_overlapping_addr, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(disable_locked_transaction_support, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(little_endian, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(default_master, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(dummy_master, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(default_slave, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_enum(error_response_policy_enum, error_response_policy, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_array_enum(error_response_policy_enum, master_error_response_policy, `SVT_ALL_ON|`SVT_NOCOPY)
    `svt_field_int(default_slave_resp_check, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(decoder_hsel_assert_check, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(max_num_rebuild_attempts_on_retry_resp, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(system_monitor_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_coverage_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_all_masters_grant_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_all_masters_busreq_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_cross_all_masters_busreq_grant_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_all_slaves_selected_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_slaves_selection_sequence_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(protocol_checks_coverage_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(pass_check_cov, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(display_summary_report, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(display_perf_summary_report, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_array_object(master_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(slave_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(slave_addr_ranges, `SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int(enable_complex_memory_map, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_array_int(multi_hsel_enable, `SVT_ALL_ON| `SVT_BIN|`SVT_NOCOPY)
    `svt_field_array_int(multi_hsel_width, `SVT_ALL_ON| `SVT_DEC|`SVT_NOCOPY)
  `svt_data_member_end(svt_ahb_system_configuration)

  /** @cond PRIVATE */
  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();
  /** @endcond */

  /**
   * Assigns a system interface to this configuration.
   *
   * @param ahb_if Interface for the AHB system
   */
  extern function void set_if(AHB_IF ahb_if);
  //----------------------------------------------------------------------------
  /**
    * Allocates the master and slave configurations before a user sets the
    * parameters.  This function is to be called if (and before) the user sets
    * the configuration parameters by setting each parameter individually and
    * not by randomizing the system configuration. 
    */
  extern function void create_sub_cfgs(int num_masters = 1, int num_slaves = 1, int num_bus_masters = 0, int num_bus_slaves = 0);
  //----------------------------------------------------------------------------
  extern function int get_num_masters();
  //----------------------------------------------------------------------------
  extern function int get_num_slaves();

 /**
   * The method indicates if a given master's index is participating
   * based on the contents of pariticipating_masters array. 
   * @param master_index Master index. Corresponds to the index in master_cfg[] array 
   * @return Indicates if given master index is participating
   */
 extern function bit is_participating(int master_index);

 /**
   * The method indicates if a given slave's index is participating
   * based on the contents of pariticipating_slaves array. 
   * @param slave_index Slave index. Corresponds to the index in slave_cfg[] array. 
   * @return Indicates if given slave index is participating
   */
 extern function bit is_participating_slave(int slave_index);
 

  /** @cond PRIVATE */
  //----------------------------------------------------------------------------

 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);


  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  /** @endcond */

  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 

  /** @cond PRIVATE */
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  /** @endcond */
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** @cond PRIVATE */
  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

  //----------------------------------------------------------------------------
  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);
  
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();

  /** Gets the slave port corresponding to the address provided */
  extern function void get_slave_route_port(bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0]
          addr, output int slave_port_id, output int range_matched, output bit is_register_addr_space, output bit is_default_slave, input bit quiet_mode = 1);
  
  /** Gets the HSEL index of slave port corresponding to the address provided */
  extern function void get_slave_hsel_idx(bit[`SVT_AHB_MAX_ADDR_WIDTH -1:0] addr, output int hsel_id, input int slv_idx);

  /** 
    * @groupname addr_map
    * Virtual function that is used by the interconnect VIP and system monitor
    * to get a translated address. The default implementation of this function
    * is empty; no translation is performed unless the user implements this
    * function in a derived class. 
    *
    * Interconnect VIP: If the interconnect VIP needs to map an address received
    * from a master to a different address to the slave, the address translation
    * function should be provided by the user in this function. By default, the
    * interconnect VIP does not perform address translation.  
    *
    * System Monitor: The system monitor uses this function to get the
    * translated address while performing system level checks to a given
    * address. 
    *
    * Note that the system address map as defined in the #slave_addr_ranges is
    * based on the actual physical address, that is, the address after
    * translation, if any.  
    * @param addr The address to be translated.  
    * @return The translated address.
    */
  extern virtual function bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] translate_address(bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] addr);
  /** @endcond */

  /** 
    * @groupname ahb_addr_map
    * Set the address range for a specified slave.
    *
    * @param slv_idx Slave index for which address range is to be specified.
    * Index for Nth slave is specified by (N-1), starting at 0. If a value of -1
    * is passed, it indicates that the given address range refers to the address
    * space of the registers in the interconnect. The data integrity system
    * check does not perform checks on configuration transactions which are
    * targeted to registers within the interconnect, as these transactions are
    * not targeted to external memory.
    *
    * @param start_addr Start address of the address range<b>
    *
    * @param end_addr End address of the address range<b>
    * User can configure multiple address ranges for a single Slave as below <b>
    * Example: consider following address ranges defined for 2 slaves in a system<b>
    * set_addr_range(1,32'h0200_0000,32'h0200_FFFF) - Defines the Address range (200_000-200_FFFF) for Slave 1, defined as Range 0 aligning to Slave_addr_ranges[0] <b>
    * set_addr_range(1,32'h0300_0000,32'h0300_FFFF) - Defines the Address range (300_000-300_FFFF) for Slave 1, defined as Range 1 aligning to Slave_addr_ranges[1] <b>
    * set_addr_range(2,32'h0a00_0000,32'h0a00_FFFF) - Defines the Address range (a00_000-a00_FFFF) for Slave 2, defined as Range 2 aligning to Slave_addr_ranges[2] <b>
    * set_addr_range(2,32'h0b00_0000,32'h0b00_FFFF) - Defines the Address range (b00_000-b00_FFFF) for Slave 2, defined as Range 3 aligning to Slave_addr_ranges[3] <b>
    *
    */
  extern function void set_addr_range(int slv_idx, bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] end_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Gets the local slave address from a provided global address
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a global address into a slave
   * address.
   * 
   * If complex memory maps are not enabled, then this method utlizes the
   * get_slave_route_port() method to obtain the slave port ids associated with
   * address the supplied global address, and the supplied global address is returned
   * as the slave address.
   * 
   * @param global_addr The value of the global address
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *     mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *       indicates a non-secure access
   *     mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates
   *       a write access.
   * @param requester_name If called to determine the destination of a transaction from
   *   a master, this field indicates the name of the master component issuing the
   *   transaction. This can potentially be used if the routing has a dependency on the
   *   master that initiates a transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @param slave_addr Output address at the slave
   * @output Returns 1 if there is a slave to which the given global address could be
   *   mapped to, else returns 0.
   */
  extern virtual function bit get_dest_slave_addr_from_global_addr(
    input  svt_mem_addr_t global_addr, 
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output int slave_port_ids[$],
    output svt_mem_addr_t slave_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Gets the global address associated with the supplied master address
   *
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a master address into a global
   * address.
   * 
   * This method is not utilized if complex memory maps are not enabled.
   *
   * @param master_idx The index of the master that is requesting this function.
   * @param master_addr The value of the local address at a master whose global address
   *   needs to be retrieved.
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param requester_name If called to determine the destination of a transaction from a
   *   master, this field indicates the name of the master component issuing the
   *   transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param global_addr The global address corresponding to the local address at the
   *   given master
   * @output Returns 1 if there is a global address mapping for the given master's local
   *   address, else returns 0
   */
  extern virtual function bit get_dest_global_addr_from_master_addr(
    input  int master_idx,
    input  svt_mem_addr_t master_addr,
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output svt_mem_addr_t global_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Returns whether the supplied slave address is legal for the slave component
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to indicate whether the address received by
   * the slave is legal.
   * 
   * The default behavior of this method is to return 1.
   * 
   * @param slave_idx The index of the slave that is requesting this function
   * @param slave_addr The value of the local address at the slave
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param target_name Name of the slave component that received this address
   * @output Returns 1 if the address is legal for the indicated slave, else returns 0
   */
  extern virtual function bit is_valid_addr_at_slave(
    input int slave_idx,
    input svt_mem_addr_t slave_addr,
    input bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input string target_name = "");

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Returns a valid address range for the given slave index.
   * 
   * If complex memory maps have been enabled through the use of the
   * #enable_complex_memory_map property, then this method must be overridden
   * by an extended class.
   * 
   * If complex memory maps have not been enabled, then this method randomly selects
   * an index from the #slave_addr_ranges array that is associated with the supplied
   * slave index and returns the address range associated with that element.
   * 
   * @param master_port_id The index of the master for which an address range is required
   * @param slave_port_id The index of the slave for which an address range is required
   * @param lo_addr The lower boundary of the returned address range
   * @param hi_addr The higher boundary of the returned address range
   * @output Returns 1, if a valid range could be found for the given slave index,
   *   else returns 0
   */
  extern virtual function bit get_slave_addr_range(
    input  int master_port_id,
    input  int slave_port_id,
    output bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] lo_addr,
    output bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] hi_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Method to determine if a supplied address is served by the default slave, or
   * if a valid slave is mapped to the address.
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to return 1 if the global address supplied
   * is handled by the default slave.
   * 
   * This method is not utilized if complex memory maps are not enabled.
   * 
   * @param global_addr The value of the global address
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave addres.
   *     mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *       indicates a non-secure access
   *     mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates
   *       a write access.
   * @param requester_name If called to determine the destination of a transaction from
   *   a master, this field indicates the name of the master component issuing the
   *   transaction. This can potentially be used if the routing has a dependency on the
   *   master that initiates a transaction.
   * @output Returns 1 if the address is served by the default slave, else returns 0
   */
  extern virtual function int is_default_slave(
    input svt_mem_addr_t global_addr, 
    input bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input string requester_name = "");

  /** 
    * @groupname ahb_addr_map
    * Set the region range for a specified slave within the specified address range. 
    * @param slv_idx             slave Index supporting multiple HSEL signal
    * @param hsel_idx            HSEL index for the specified address range.
    * @param start_addr_hsel     Start address for the specified HSEL index
    * @param end_addr_hsel       End address for the specified HSEL index
    */
  extern function void set_hsel_addr_range(int slv_idx, bit[`SVT_AHB_MAX_HSEL_WIDTH -1:0] hsel_idx, bit [`SVT_AHB_MAX_ADDR_WIDTH -1:0] start_addr_hsel, bit [`SVT_AHB_MAX_ADDR_WIDTH -1:0] end_addr_hsel);
 
`ifdef SVT_AMBA_INTERFACE_METHOD_DISABLE
  /**
    * Function set_master_common_clock_mode allows user to specify whether a master port
    * interface should use a common clock, or a port specific clock.
    *
    * @param mode If set to 1, common clock mode is selected. In this case, the
    * common clock signal passed as argument to the interface, is used as clock.
    * This mode is useful when all AHB VIP components need to work on a single
    * clock. This is the default mode of operation. If set to 0, signal hclk is
    * used as clock. This mode is useful when individual AHB VIP components work
    * on a different clock.
    *
    * @param idx This argument specifies the master & slave port index to which
    * this mode needs to be applied. The master & slave port index starts from
    * 0.
    */
  extern function void set_master_common_clock_mode(bit mode,int idx);
  
  /**
   * Function set_master_common_reset_mode allows user to specify whether a master port
   * interface should use a common reset, or a port specific reset.
   *
   * @param mode If set to 1, common reset mode is selected. In this case, the
   * common reset signal passed as argument to the interface, is used as reset.
   * This mode is useful when all AHB VIP components need to use a single
   * reset. This is the default mode of operation. If set to 0, signal hresetn is
   * used as reset. This mode is useful when individual AHB VIP components use
   * a different reset.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_master_common_reset_mode(bit mode,int idx);
  
  /**
   * Function set_slave_common_clock_mode allows user to specify whether a slave port
   * interface should use a common clock, or a port specific clock.
   *
   * @param mode If set to 1, common clock mode is selected. In this case, the
   * common clock signal passed as argument to the interface, is used as clock.
   * This mode is useful when all AHB VIP components need to work on a single
   * clock. This is the default mode of operation. If set to 0, signal hclk is
   * used as clock. This mode is useful when individual AHB VIP components work
   * on a different clock.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_slave_common_clock_mode(bit mode,int idx);
  
  /**
   * Function set_slave_common_reset_mode allows user to specify whether a slave port
   * interface should use a common reset, or a port specific reset.
   *
   * @param mode If set to 1, common reset mode is selected. In this case, the
   * common reset signal passed as argument to the interface, is used as reset.
   * This mode is useful when all AHB VIP components use a single
   * reset. This is the default mode of operation. If set to 0, signal hresetn is
   * used as reset. This mode is useful when individual AHB VIP components use
   * a different reset.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_slave_common_reset_mode(bit mode,int idx);
`endif

  // ========================================================================================
  // The following method must not be called by users even if they are public
  // ========================================================================================
  extern virtual function void set_num_masters (int num_masters, int kind = -1);

  extern virtual function void set_num_slaves (int nNumSlaves, int kind = -1);


  /** @cond PRIVATE */
  /**
   * Returns the configured error response policy type for the provided master index.
   * If the index is not programmed, svt_ahb_system_configuration::error_response_policy
   * will be returned.
   * 
   * @param master_idx Home Master index to be used in the lookup
   */
  extern function error_response_policy_enum get_master_error_response_policy(int master_idx);  

`ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the APB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the APB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif

  /**
   * This method is used to calculate addr_sel_bits and to convert max_addr_boundary_limit enum value 
   * to interger value which will be used to check whether transfer has crossed boundary limit or not.
   */
  extern function void is_addr_1k_boundary_cross (max_addr_boundary_limit_enum max_addr_boundary_limit = ONE_KB);
  /** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_ahb_system_configuration)
  `vmm_class_factory(svt_ahb_system_configuration)
`endif  

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
z84mUQhy4ymSTZDeXlIhpRms+i/gN5mRdTSe9t51YCQmOXsftZ+g7lH0nBzd56OB
KcIOSv3S/WAKXK8NniafKw2Vca3ORBOQQmbkGQ9aByks59g7vfmir8FggNhiPHh6
LSpq0O1dB+UMZgCw4g1x2QBMDefU0c5VmAMK4c9dKoCOn7pE5tj6Tw==
//pragma protect end_key_block
//pragma protect digest_block
QdeMxcyjBUVWnw0EJM1SXoJKC9k=
//pragma protect end_digest_block
//pragma protect data_block
6VG4z4z7snQC5ndkx79oN0PfG8pTyF8Uz7RwiRu7WGJahOcydftW6L26aE9cpMAp
2O6RZ9m+f3Cc+XwtzALaECquCuN412+o6wbpuNYuPa23O+/WCekM3S+Vh5a/ssQW
wc2qLt0ciXqr9ojL9x8A9IMmNb8pZhen/d9A7FDiEWT6qQ9WUOX+yv/STGwL2zIA
Sicg4xQI6IeIsKANKOlm3n9moNNacwwqKQ185VcYqHtk/PNL4MZrMe7/rP2gsce3
m4HI3DS0/7m6rHfG6WVrXWPLq+OC5RVn5Z7CSiWTn1HflyxeB5AdB5F6rjhdHMzv
dHsiB+BKGS/pLw6C6yEH3lbieym1Oiq116A85WEfCPG3BuGzhMznxGDn1L8C4Nm7
DYHdCCB5znsXkrf6vDJIbYTk0f1y+eTlDSyurbXtdBRp9IiDcgV+1U2m7BZbE4wy
JxLN94YF1yzeMGcSIeAnpb8EGQnK0av8TOtnPGV7s2JahrTJSSrDNwxYayC9tl2S
Q8Ytn5a9VzeMEUT5FLHm/0NABatYS8DJCeKiN0kT4nXXbfYOp+EgdzvVIqB+skwn
QnQrvDvGucxbEs8mX5Oebs6RCFnx/A13/CofKHdrHpYBNAiq3eIvKvSAlKRjhWAx
0Y54OtdFGucUBJH31PGnfi+3M6xtG0weJD/CcZMp+mqn4kAFBpekG2FPnsCjs4bH

//pragma protect end_data_block
//pragma protect digest_block
+ZH2RvFVyAh3Bev1YfXwy7ljfW8=
//pragma protect end_digest_block
//pragma protect end_protected

endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
OSLVxsXlZS9m+Xm76mnlanSP0DO3sIGciTI8FNNzM6+uKhndkBo46Dyrmmh4J2UH
ZMfESS3NxUiDXqW49evpNzNzRtZAyZI8+fect+PuHtafMaapAl0eBfIZWXBXyi/3
ekM1779aiZ8q/wxm8zEBBWCYCFvW8Ug0tp4LH4iTWGkptEruuHv8Tw==
//pragma protect end_key_block
//pragma protect digest_block
nNCJwJbAjzR/u09iO4OHgwf0lf0=
//pragma protect end_digest_block
//pragma protect data_block
MLKO4etAjMwKWBtatwV9bq/62wK7rfhS66ey5whKliuJBFoD3N2tHZQ+VTTqug++
O3ShKwB8kXAvfliG0PyV/ygPARCkH7pihWHpJdhwDA2MIbEZTzW9XxMOZ2Kt5QW/
ctCceh1SYgy2qj+H8rpx/rRhtkKduahhTErc3tWJM2lgckIg2XOXrIYLDiylLt45
Rzw899RzVRmTtKsNzozuBIkpAgHc/Odri3J18mfBcRtV3uH/p31Kjg8y5h/6vbAv
SkbjGaUNl794hBc7EUFJyShDz9YZDiyhZGdNZ0vR95ArASB4hT8O9/7lrfMNrv9n
hr5GdOrADdcvQp2RsYCBcc3qP16XOH6NNiVkiVvD6b3DorcL3I97uMOQNFRHGEPj
oYwXQUhNYZIj8YhRf9CXBJ3jFVjGvufUt603atJySCGl+QE+/lez/cuA6Jac6Afb
+ubq990Etcnzq2bm1ZtXQ6jPnLv0NQYqoVMz/tDLRV5KO7NRMZnwvN1T5fKbBfvj
5sVNix2jLi5InlL9b9JrIGDw+wViQrybss5d9F2oyAV7D9gZ3FOmi7yc5OfVyU7n
nDbzRQs+uDnIpTHsX5oll10U7f+dgj1DCeGDMjQ4KVCgP2kKVNi+Qni5shefLD+f
vYtTwueQ39iCzs0cl5Mgcw2fffUTY2MEgOf81C394nDDZxQkDYXqPRBmb0iH/4kY
dzBgowZB6NALu2jcWAHlV0RK6lTXFrQQLr1GWB+c8pp3We6or99Q4ehBA6pO/C2N
iA4Eg3CgxYfK8FJUlsfbAApgW6HTWkSICdLMUHF8/RQOAMaiBvpibRkmn6C7/nGR
4CMv+9mprL+a2lvLVmCdOaDCZbmWxUwgLwr3W0AtMgHSzucYbbi++CGao6qX56FY
sDM6lV8alS/q/8ZV54rmymU3tfL8YECA8OpUTu1ivisybM9AInyeG/JHzlW8sDCE
HWhwTdM58h5L5LfNsNaBEVNLgdIEU2h1Vl6f3wa+CkQydaVUIP+l0ncBd3TWaaho
8t26zyvB8YB7exMbZrnb4bEg+cli4ndyAPxAB1G0X063jVW9OaKmvwQRM4AtkMdy
1Dj4pqf5vOzt1eVaN0qtFvNlA0zNR0FecbZa7LhdFcPcBmifYRw56aVse/1P+89V
rO3Wm8blnPJn9DK8ojSWMG59UBy5mMbervsSUnCFO8FKhPb3LVfJteRS7aRqFN/E
Tt18VaJ0GoqFwoyMA1m/aJjgpfe0yrc0TIzPpl01SYqPslVw2/QmuxyunRKuxhOH

//pragma protect end_data_block
//pragma protect digest_block
W8NAsjajcfJaJQuyV+UKNtZ6aeo=
//pragma protect end_digest_block
//pragma protect end_protected

//------------------------------------------------------------------------------------------------
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ryyeN2C76UuuPegA3hho1SBGmWz3KXjpay2ayU2ihPFTxzVjrgg9g7mb3CPbQmLW
JokxOA2NxqbTGssDbF7X5Ceg+owecLS/6J0hx0FhWOjTtkvZC7Cp/wgj2n+LPL70
66Bj7Fv0vhV+ZUE+W7AbFeBDBsp7JBmnjtSY9QRV8UGZrcvuMyniMA==
//pragma protect end_key_block
//pragma protect digest_block
wM65TdC3G0X36fwqp2SU9XNn1ls=
//pragma protect end_digest_block
//pragma protect data_block
ooBL+b+IhimkdWKnKEfJbpA60g0+o2O75WeC+8Mx8DirWgCOLOBYnszgBp80ypZu
nKLC5WqyN7e5H47hQiZ8FCYPlTJbVtYzuxC+fP8ocKvHu6hXczCoVjc+0og5fKio
uoYe1l6FyjteaxCA9mW8Nm78Tz5I6j95qAtBi6DEMVvIbgXdZLcudXL7BiZLDsJx
pYoGfCj/ypCcDhGt55iXWtFTBhHT7XP6F/du35pu3vkDSxix1qolk75IQP+zf0B+
yH4PxQcY3YsrHyMPgwBbg26m4o1+o7FfPa7FnbMPu84KijiVF9+a6IKu/tI+99rI
u9omHORvyYjRhzXg23/QDWYJ7afOHt5FqZzyYppt64+EvH9MMyYJUtKyu3kBhfsC
4GlvOZVC3BWP7330BVAyPF5ejKyZ2tBKg8wevjZmd/GwuIwf+B4oTDfRe8wWZQZr
LqIyK89iHBO8HLJBbte/xgo8vMDGLd8W0XwUS3DfRoXo4v0XC9NbZS59ub0XGhUl
tfjzRlIvqQcYQShCXB2LR1YlTTm06tHAvf5zHzq3oeJsqyRfs4Yn5j3kmDML8JMe
Vvl0KbOxpbc6rZkgrIMH7qkDADyQ1Fe1nS/TLhm/I0ylDHR0F08XUol83XotIjt2
XdOXh90z8gXyGg6GuT5QNg8M2k3ztJV/VFRc5v6wKblQXSwgFpccSNr1OLX2uySQ
CVFOyY7FXEFKrujaXvCGQxsnJHB64cfl0ew+DHE/MafpRG6SBUcP/jioeKIxoPFE
b5Keb3bKDapJLYOKHPDhFRWE1MYFEqoi+uYrJhVT9LCyr2GfJ7nr123XGJgsAXcv
RS7xEROQ2qGsdS0yMhb35PbUAJGQrjwEZ4vL61UAM1z+xgi0IW5s99sWo0M3olAB

//pragma protect end_data_block
//pragma protect digest_block
ft5wQyTukpujVqmitkA/T93DHkg=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
6KyHaY7KNs+5q66ckwwjQ+5bDN2yGusBlAgNSyt4IzbvrzVE/G6y8pj9IJRckl7d
/JPk1oU42PtEE/2VEC9QiLIZ+Rtt/Wn6X7T8bR0ix6spwqU86o/mmen8h07439z8
YCst/moa9gJNrZIrXhG/eeGG1PUhjt/cdRsLeJkY0F1AWes8jHuDOg==
//pragma protect end_key_block
//pragma protect digest_block
pOhL8bGmjif/xRKvstmw6b40wrQ=
//pragma protect end_digest_block
//pragma protect data_block
6OLk/jqA14eCQE1QKv7HXJ/m4H5TF6RIgnYl61iUDfL1RofcaLKxIKKzQ+WUKHU9
nUzMKL36YyrsP8JilHvqsnSHcIdWCyU66z3xIpjAVosRDpVSkW1zWXBzIbSo15qq
hAKrqqg6WfjxVAEAP6Zhwu0nsYdvjxnSjwrhJPKiBKHAG/vRcvqjvJyOC+ThEuj4
KspRuS3tqtKjXW77M6+FbTyvuDq/yNPWyco0nc8ieT2R/WVlI8HxFWuEzhuRXbV8
F/prPoY3m64lAkKtbJz+Fr2m3b9QYb+x/jOjoWzdaSCdXwCHG918tBmewUABnWbN
M2YHSYVapvfBZCD7CFWBWZTV6Y+cGwvDqrycfrtd57AmCe1sl41SY91on5zAAPYR
0g75NfV0nowttKyfORscvvTH5VxADGJALNr8Caf8fd9gnlKHI2242/jCM/hw5zg0
JSSq+ZEO1/qVYBV27gcdQbdeTw1FmpEJeb85YOVToSHQrMcEW2s3WYptBpvdp2yO
25LmYpNWa0g76Ka5alrU6UKL9VXVkltmDdR2zjiGrkQzi/WZXgGEWFP+/zltU0jq
I8VUvB1u3GNfkHl9XRANpDGAlvCIKFDiqatUz0RZaS11ZfsVSnkyeMtar+m3AZYb
rrgT4Icp02v8JyRwMj8m+6h4u5rSAYZgsnjbNd79qzKY5gqts+6rhIhFo3TFOUt5
VyP8KqujjwZKyuxU6SOph6bQdkgTErm+mW9n4sg5uYA/O/TmmihsLvB4emEaZEBx
ARuIRFOsW7PMJdCSOaffpvnQ49v/T5MsBR7OncAnkAUwq2bwAMxp3M5Z3uVFfHig
gaQHtQGB59ig/OxH3Td1A8m/Pr60EEpKVOaoNUJ5i9hMEYOrMGY5/KVCbiG1IphH
WgM3gyEw75bGwxEUlbiacxkeMErDj0IhMeX3OiWK6r/tihDYSP1nG9N+MRq/zTKj
bvNwEAip3SG15S9Jl9gKqCleDFPgxIsdSWuQaRbHCeJII149GSaaUCMUEITe4Njs
citbQeI0zw57wy1OR1/0Dwxa11YJ+g+PRpJ//slnrigFUfQbpFolKEoJgIMWDxj0
THRJaLNG+HbMniR2vCNstClPyX3LYjnSTQRwaA/n59BFH+KWqTJOhsJw7Q4Btty7
BBvmlrhGXBHl7Z3GmWlG26YEuhHOAAo6p/BpvjTs3Y45JshxXXbeZxA2YJKJUMeJ
Z+dIleYUuS3dVNWHxFiyPOo8unbj7pc0HlUaYH7uxHtePx3JNl+KRqtxlvnQZu0g
mEquRYTv+YPLue1+XCjO9Amw2+a+vaKPcNVR/yu6ZcdI+yVI0K/xO/fx2ACJ12WV
irN/ZMb26RJ0bmahtZgXWlrflw9aZe7TgWHGXZLRP5LgUlmrdgr5z9JRgbOL6EG1
RRmYNid7/dFPkfE/IbSSCpSP5fTC7Ig+eLnYdCiHAcUYcgugkIsftkIAHmkIQf8/
GgGXGyhh1ErEqpQecfHJlWbcOVm7voun4WSk4C9G32ZbusHjWeesxBoi2zBCHtSY
gFV0Jb3pgkyrruc45qlKFlBq8d7FsRmxa7TJ9eHsTOgKvYEbts+kFxa55td9l9x1
kxC+4S9hTAVR0+UJSHJh27Vc4dSMDefsTM9c0rHhvgZlAAVYTK1RpQQ9IhTarO0h
ANf5MGN/f8QmfdWuEeP1gErDYZehLrSHlNUJ8nDdtBO3B3n1mWOYNVzdYzG2r0N9
3AXs5b4hT7fr5cKi1iFYmhZta7Mf+Ei0Gc7NsL7vbIXi0vrLKWBVaSgEBd16JWKc
6QuBII5Qwnj/irZr7VdnZ0hlT0vEdJg0h514FiFPrYq5J5jFXzusfhT/TguhQtP5
GpWCtXVtbb/2J82ILBoH1jrPIhPW+PLJD3lnHFaRGQuHYAzDjeQ65VIlahD57xQE
lv3Dlv5e3N74yb3voPFltS6T7XsmsD1PPdQg6VbL+clTvLEUBR1m49UPQUCcpKxQ
S3nTzAjEQT7QdesJXXKY9Q/Vq2ytkZWWL5JMoT53oAPxGpxRu6F1I3zgZMN8v1YE
1509d93iyhbQ/cY9mIhPqQimWLEXJ/Zoy8/P6lHvCYxoAxXq6Cf9oUjQ7cTQLg+y
jMSAOmoSaEMCv3cl7aDjh+KFcH3q1SA050Vh3POadfF94iAffiBj2G6YVwgD+Aiq
+Z8yXqKI5eFeT/abJ3Jii2gW4bzcejXHNbw462cqvnuC1p78HyKsi3ADkqs7zdcE
X6sbBAoPKQJ3izvTzlHQ6KXa/vRgD8JfNtoXG/3NUHrHOee3M5CQ7huQYP2IA+EJ
U/TfmAET60mhhDotym4AbhH88H06JumArG8a4AHtxIdsudnMvnJOSTy7FvND//tA
4z1Y4aCH7DfLKeUkZLU/sa12ER1Jh6M/uf/ISFYjzK2MSGxMDYNDIE3I5Rz0eBWN
K9237VsJucCrmCUeH0gUV3OD7vklLbCn/Wy6vnqKukKbyqxOSLsYLliTO8bsscQc
wDv9Tzh7t4SZSNKO4rAszqHh5kQeIXHwZDJSVf3h0vXJ0SSLXxlnqwkNVYkdSzDg
RDoCbRESAuryXk6yP+4VUN23wQu9/MTG4piyn3518AIq1i1lLk5Us16HZH+N8OpE
K9l71WSbWNYqFmP1ISOYrbfAY3kEaCKcUOGnzBDmgbmu1pG7RyMCUGVIHNR6KzsF
g1j5eqsdo2TdlxOmgoqhrmRtEdBVN/XaNzOyMVdkq3QixCkf7068nFy2Sc68oYbG
X/pDi6TKMaM7mdpKN789U7vGW3/hxY993aVIzYoBxzGJHNAYNhOhwgBARaT+q6VK
/42bnx7VvRZMYg16eoa7LBhGkcGrScRgaUgO02R4h0KNaIjbWqzU0VkMfupH6NY3
3cfRPA5hmL4wJ+hYEH9Ta0m15qxzbCW9RgDR4uVMpYUKOyT5mkdsj9HDu2mZQbGE
NfnV9iOFuYn/rSlTMtrLsrhxqgmhRjUJRmAPaxHo0b75onQfRR7HjXoGYrg9FY4w
fDFU1QWokF6bxY1p37gy95L5kck9HuqqJExgQJgZU+NJgwYypUMwVDhVw8EZvgLH
a0xM92XGW7CkI1dpEhAgLdRvX7/h2BlfzOMXqQ04eRgICwHs3FH+TsEMMEV0bU+1
eqzbdA5kiOMeNkol8GFiDJyOL3vXyHv0sdhyz/IEiIXYkSOc+G4Jbl/QZsF1kTjV
Gqf7GwTvF3HIrPekOLGUd2FJDL/R6omlrWJNrDPDyU7DRW/90XZUeUCWci9K0avX
QJ214aRoJx8MdApWgzsz4dJvqwkUTMC+Uo3LgFqqJhEkUPI4VXMAaN2XBGFCH37g
E0LELNd50tcJUXYf8Sm/p/BrHjxOEdL9ixkMzNuVoKqIXG8YtxjgEECji9WN5IPT
kPMpxLxKlomH4dpmRjYEZbLSnlev4qUfnmU8EYXHY4z2ya0N8b7ILsabtt44Njfa
0pH9fc1oZ/cpXLBFNUICdDn8LzmOk1+rGpkmckfyodu3YLs+1vhpXScMYupYYnuj
/EdtdjmVnYfih3xGg3ddrmxcm/PkMddMq5vs61asNOzZqKGpTnc/lZCwmf/9f8w6
9CZ7VtQyb+ryVrvrVXkRP6O1tvaCmZXJi4dDFrlZSPfU+iRji8FPd4+6S7Jcxc7O
a3P9Ats08IfV0nEoohYrly3kPSpEv9vFHkWBC9W9466RmJzSHxIHrfhFgoAyHmP9
/FA9FtBW505vas3QKtMt7anzo857GzDdPuodVQsbMqLifwlJaaKYO+VUPR6GMQTY
FPO1iVZi5FM2VI6XYYOQwjC8D0sLe+QiL3YDwwZ+10H64+v2GEmeEe0/Sq6mgRoM
HnlAEqvcNHKUrJk9Yt0f30AM6sqdcuAgHk8KmOSByZ/NIxLXDd2OlmaOfzs5dih0
MGwvZZJRPuokVg9H7KGeaQvf8nuWxzWuLRHTxzm5E6L0kpYaQTtCWk4tTHBpyqMy
PWrtX80G21uv9nNK96fWXjPAcaS8DZcURaVS43N+hwr+tIWBeRUWe/IKgEBi6QpM
7PszjGgELeos9KM0Hx9KVAkoATD2OQscEbBDzWYPhTIA43XdlFzf1sZS1ZUtX9jl
k+kqJvZVtwAHhbj5r3PS2lmBlZOXBX7WOyaiGGsl7tjoI+FIMRw7Plm79jH9bb1n
mW+h1iYh9dEhGOOkbZG7vqlDrkLfcSNa4j3zVtvchjCYiPI5RG/WPetj5v28EtdJ
77IwG+G8U0X69dU2qHMf9jQ64+ZdlVsnt/a2AsHGJhlyqZ1hPMtUDuX7f/tag9+k
V9nJxb4Woef2aVyZrESK1ImMkabR2NdeavWRvPWi2er8MZx/yZDNbVpVMZl3kain
NQ8BgFnIHpEV+8pKUiTSiewqvn1eB1aNI9xYE/61j9YX4lmlSLRqwTIsREJ5ZRV/
ZDi7U3ctE/JorSPl4CCn0dHwanrE5BMwGprwE0+94UhLOh+tVhkyEw0grFQ9YteT
2AaHOPLuE9YQqOyz79mtPFIpctPTSZDrdzRtCNOngd2O9/39XgjJJdyG3E3v4537
rNncsc4pPTng2PH7eMY52ROrtH/TpvRAWWr50N3lmCzYWg2UxeQpvmFoVWtdi0Op
8p+//vTggwF2CsRVjBZwdNziOjlZAN5EDxF8sT/YT7flP6u4YEM0o64hI6W3Pj+r
VvRNlnN46vYBGUi5F+eBSnDmTbO2CJJWspKewY6CtbIg7xtqmU/ugPdYWgvcHFJp
n1DEqrRUueOm+Dq7yPKxavU0GF4Zf7UfmEACZ6qMmjTW253CBJd8l+b+0Be1/n+5
w/6WJYvZKmbL84Nsyt+pUjZNyLvgKlAIunyhiR75RjqRZQBYtOYyN1GEokNbEj2W
/pIRrMemlTahXejogNwDy/oyEG0QBa2maKAKeAYUE40wWe8N0OaPR5f47Klhg1CP
2tcVb0sS8RldYWMNjm/WbEU7O5oi2Y1aeRjbBhINwunpHN9pr7fmEONdxY0BOVA+
kfifuhpJRtOLDEHP2dKpskbD3u8Okno5HbfLVHPoJ+cgkCd/io1kvgYUQNexX0iD
0OTV9WA3/ePm9rI1DJvy/Xr+fBK8VfGoHHei1dLigptILdcWG36xQOZL/CfTIq4P
F3yVY7FhDypsOLwQArwwp5eHjsZ7R4thMZF8qREbB1DAEt1P/W9B6Uo6hxMwKr7y
T4sVMpFr4eS1ipsWVS4zwgUU1jh0IHbPABUYLNSJjGnqCBcHSukzFcpQqshxUslR
FfFMHBsjUm75rTo8DY/ezGn22ZGUWSgEcZJgEZdAFCFYOvSxcj3l6JEWOmejXeqk
YFsqwMprDHNgXZenbyRWL4+7/3Qb9uBQ9zTbj8JUPxE/9jez7YQodGwGgFN9GIL+
SvWf/WjUh1nDEjy21GbFOSoUlMMMtIrBECV53UXDVT3zujkq3bEnIK5gfORiJtHz
dV55tXaTN9nZGz2zIRigFn6QDv65qnTHH75nCf8uHiVvKCdX3thoyp/NH1jGYzwA
ab7m5D1qopVY2L7ymWa1vgylSxnwG37bhjf+qMnSpzq8uPJ7g0PO9nUsTdQpeRLS
Lg2NGaAGhsp4oA6yKDCa1TdTtrVn2UMaRNH1hKyr3tvk2UBR8TSQGqbeRvxVRDId
zwSJ6an5/6qY5eO0k2AZO6FHgQKx9qHrcd5k1fLpN+1BV5THbcfeNDcEYdTq19GW
FjuTuCd1rmkpLNbXFdf0/pfjQVbNYked7p18alQc4lUw7f6U/+UU7U0AgFkD8nzb
9W6BD5JkxeX+1gpmxsn33rJfZOxeg02PMCGcf3x7ve6wLnwVC59Z4hCGYTso7Y1/
rNsLL6874hp4oep1bfHGvJcWDMfp2JMfgIbAqTzZlKBj6oAZ8J9RELYCVMlGoG2L
AM5qsA34U1CyWdZ6ss5joiT2zH9zXY/x0kjzbUSnMxHX64V/jRmy4mIMbVdTcKgw
iHxn9PokpTK+UbIllr5OpzgxZyDW1kyK7oND5veujrMfyDQ+HZZT+WTNrXuAc9vd
s3TRKT856tDN6yTwLj+kRi+r7K3X668enfVmtUA0kI7nOsZcaqUHc9/RexFMfjl9
/HZvAIbp+3v3nPlC3k9H7odbek7SNkFSE9mJQTXUiKrAfc1sfxQsEN3zdbjLzhmG
Bt1QJJ05WS/4RhGSkh8dgHJ0bLjIc0nMz6H70znSyhccPJBPzehVin8acJZl+Zaa
abuA2Ng/lwqBhEpNge1RVNWGUZhtFhMAdwgbxRZdsXimgtxsdWZRnMMwLwqqTb6l
FckJ+aJ9eN/7PmSIQILihaW8Kp8NgxI9zyD+pNrtz3qRcLYe2Ap+sfqr+vS1JSb9
x4lUtmlu3DMH1M5uHNtfFgWZ7cbj/IvvGoRo3u4+5qbjy8k3NSL2g5FY6OFbjNEA
HSLOB/tV0T1Z4TDVH0AH4bhDP24eFjFdBsdS8HnART2n3OBFmWrv0Exm85fHwUqx
K/n7oE16Ca08ceOuOxqmRqKZC9ym95y4EcNF72tQqC6WHf0vnzQmQCD5EfoW0AOl
YGx+M5domWYQYYHqs00M7MOf1+M0r2MRjC/yFHZwEOzLuifQNHk43QGlrowfWteh
p6OyfebLlzDHbmHntsyF0gUXtvKXv5jtxIKrIuhAjd50BU0jVNnWtS0TjQFyi8/6
hf18V+WESAeGLWIrrtC/sRrDUMrExQMmvdRUmQzrtJ2BC+h0CI1BsunxTCZ4E1XQ
JM0mY3Bp9jMzAHFBN3Jxh+CcqBPSnsztgK0BPjis5he3d/MdvQSGfmBAUR0uGu1v
wO/uw0zZ1EeGrAVP3WIptPt0VL/m7MxiL3/piSzBPr2v4Tymukhp7an4ynv5TZHh
SNw6fPjTck9p4lbZ9Y2tlElDo8jjUvbQXJAyBwaN+H+KtWj9GZyk3cy7NmwhjH/F
5TmUae6vn0WG8ijoIHbD+UoHzFkf8S7HFzEBmviYH4hSeg1+/HyuAHzQpgAt0byP
IEusa9b/zwBMuSPMI7SlPP1CULxT194vJta0Zzh/xCBMTLODTDrlzkGIW+2+U86H
bWw2vvVvutETs+g3Ed7zjKyNNeAZJHJnGTUhIdpJT6zS20hqjwi+PVriowYGcFh8
LXirxsfPkm5Llxa7q8tXyqTf0HSiSIL9PrsI5M2LjbIbcyWDyXPX2gFVmPaQasCn
q6LIbClqWFMO2CW5IE2M/NhI06VSlpKF91jtORO113U7rmSsC2hJpXb0USOWpAz+
OaViAyL4S39rdFAHxG+gSFmRASkMCnrN+BBJ7Zb7wMFc5JbIDVNoQjgY0gKqNDQQ
1WPwCujI/4/p/6QsKJDTOr6sbTgXRgA/3s8EtkelnI+BrXWBr35I85SGk0FUalTD
f4IxMEaAcxtWcVyZIHEbvByLNe5TU33uZRck1Ljii9K+aB2BKajnApQsLLm3jKFW
n/Hvj8EvzXAROJJCmpTexzeesJ4skDolHehBJ6/EVrYc4vhToybU7P4OljIAh1ax
zgWNFZXlx9kLl7QM2Gsmy2TChRtwH/GLL7TLJW5DNfOK+bO0lyOEZEJl7YnGJfxv
w4tNC3WusnFzhaFktlF5tSxvluffnSjXe1/OF3z4I0k5p4/TT3MKbu/UM80RHu7y
c0AMTTXfNBx1W2h9Peq40oh9VA7IqpQrCt8NwU8Osd1uDp7Djjt9mfWyREG4xHgy
vvEo0MjMU+K+a5qGPz/D6H71ZSuIxi5nAWRxyEmESwwcHZaBRv6rtGkCdi7z0YhA
jPKhCwho40GLz5bdGGb2aWiAoS5mJ/kMN70ip75TIHZ7yA9vMjtyPL+U4CErgoE3
3kShKHBaIGlmbRn4TGWwYA3xwcuzlyI5jJr74bpf23+Zj+CbWwde8g3TC5O5d3zw
PVUW9xJngd9Bk1zunC1HnrEf3izl8rSiaMuGpO+xC4VxDOvO7dAW3jkL6wGS1P4N
wX8hYnop5c2pRs2g2as7mMpSXW5gwVCF5hsacd2J+tSp18Nl2/X+Seh/sE9FvOn+
2D/VJWnrUxlQVFfUckEqA27vRPPFkyiqeWDSUOFc4YQ+x0eMx3Z5KZvubiPZec/4
5QK4p6WcNxhb0rn8Svw6uWXm5OEK5KvOsZHJqim9u7a2flpY+5y844ugeyzVI5y6
fONU2vem/9b2eqiSf8MUUyaac3GgFoh4QY7uu5AYTdSxyy15Hq53Wdh+66d2huMN
QyTI6wMGhB6JidSTBnpFNrODugR8Y+5UqgGeZLZvHUSQJBs4Cy0hMJ8jhSxCt/Eu
VIa6ud4P3PKu78awEgKe0chFIcxHUa9ejbwpUudHFa4gBDhKvukYTF9yMVyqIafm
rnis7N2rIG8Yy3r6bPr6y5NYKzAaCCqlnZVcStG8zMaFCnMoWN4pvYDf6ek6m5Ja
d9qNs17xAGLAaOfgNZbdKSncE5mHAfDiZWX2fHF4isJm2qAjDjFQJadCbOnJIm7p
qoa4IbfxM9s4dKGrrS7mw7ALaQnItpJ86fdlqMf/1HeqxtqqhK5U6wD9IYVGS/D5
t03plP7nYVOS6zZRffX/r6xyGKz+Td+mZI/jFH3pBeRZHKB8BFkheP4BWmE2TiGa
IgyzMawd6ZHnZw7cYpAO9HHMfLI7FoeIVhVhgOqaS5lRwC8mCZtBVTQnYe9E7ocB
vFLWdrfyWFxGY/D6ie4QnKSwN4thhbikIJGqtZIQN4e4lvSFHEOoarna1CcODPK0
Iz42I2N8RroIQfb7qm+0Y/UiDkNOg6on5iSWgJK5OUu2Q7e70G22f/o1/0P4WTlo
fKhH+bIoDmDggpv/b0IASsothiykUuYE9Od5bjIG9nLMUebSdf12ydUoEbYP9jh9
1tLbGVtGwGzrdH5j96fPUt2AawqSJg54HR+X41Sqi54PVLn94tn6EtSclSWFwFft
QHh76sQvZbJD8m4qu/0LKE5Br8WaJTJcb8hTQsv20f3uz7xfmObzi4yi7YF7F5l1
XNGgEQxV7jpPn8wsUCOcAv0FIOI3GA/gx87SU0G9nZlmB2BKD6zxX2VWQtZd9d/2
KiurFNr9bs/nZ6MEeK6Q+o19VL1BLaOT5FO1LbnXVo691gKHWToNO7v/OaIubX8h
UDrD9XbiAWWxdaElOR8tMqyzj+PG7JrmGxpXNGiZI79AUEfL+q+rZ8m6yC4RA2by
gHaqGUj1wriS+G6TIelQfO3xLWQg8Ez6G0rqRSNtC1OIdxR3L6dgmrY0DJ3n0D5S
COesTANXgA/871iMt5wr8z8XzTnWFWee/wCHZWT4i0Bl58QlSjzJs7zc65A3oIWN
yjSx3sh+NafzQRZ5yFNNFqnDeO+JQ0M+x0S8Gzyq1Ih0elwcrT7JwTBmy0qQ+V0n
P/MT9Dn2oVU6aNSjnY03F4yok1Mxbu/0PdANP2eKBCeAhO2VvFUt97bvgjG90kiH
bsdW1PJ8alMUpgSyim2k8JL6/jPLSHqRYzoKtnZzGma8WI3Sb7eyx5g1aqVdzPOs
hcIXpkUUlOQnoMauaARdmmChYij34cXe/ecMrQ5wHgaxnGJTynYg6hee0RPExx3D
Yx+idgNako4dDs9MzbeCMywzJKsE78WaQTOoBxEg1ee6xaS32gYTDxNmcBRnHAnG
/P398Uh9MFq+6zNFXuFumwMDAm3+2SWgXht0dtO89PJmOmEYV6RRc6v4KQl/nf2M
dOWVqtKikQshTvqIhv3btrVno9PdHdzovlu+O2cTTgvajwsiGFGNPqVL2UXn9GZM
pLUmDGzp9noKu6fvnwI7b+8P3EFRLOmmFxe1mOlOfpIHCcGnxOu2ZqWJCiOYFRiK
pI9UXF5n5YO2L+wezsAgneAomIfvzAyyyzJcOPzBwnhjcLy9zNgwa0/EOv6azS8i
mwjkHU51BNVXPIAFZ142zxYNUoh+GkoqVmWNRN8vmIgeMxo57aROarwxVQSXd+hN
l3yTYE+rKx6QSmPu/ofy84u4yJaVJJvUVC06q3yhn1/gfKQZix7kXrWFVB576VDm
P05eTvo1nzf6nyeCq+oW5JT+HPIbvwpk3WITow4DnwC+6w61VrPW6aQgBFvwTlqp
9Q4Dk7mXKc/t3jqgH/omXJalJE4k/qJ1pMGiX0BubH7w1naQx4aZWeLK48bpHUm2
MA6ntFN0UcWYq3bktnepuqAe/7r2x+8VEVmqUjh+j/y4QHr1K2HasJ9KUalitVNz
iUJSQ1kMId7BT9soa2JQ31YWFHwAV2tPEwurA7nMwN3KYC2QMAIt2xnQiOZGmypy
Cs4ba00Ehud8LMzSEqwzQQpw6JQaKSL9iD/SvZBwtlYjf1MxH6mrEjimNh5MabmT
53AtdCY2KGzWn5UvW9f0NW7t6AqcymMNSbLClfizAERLuAJA7/XxO+1nBLKPVbQm
jirkaI4NiQO7AuCMPL74NQ9g4SnNJbnGyML3Vs0j4N8ckgkP2mRf6FWeIVJuaF0g
KAyWiphjv3Zal04azgAjvIJ9NEBdWRp96vPgU0DGWusurfsKhhM1mbbQZ4T2zl8F
pUwPrVkeMEH8UyQ4EYJP5EfJNTcaZZjOFgx+D0DBwM3Nf+FkIi9tk/q84C+JMAFb
7F9aCNfIjR4j70sm6wCUCkXMLI7oVxQJW3wcNQ6Tp6f8gdPYFAB9KQ86z84tu+Wv
mw6CP6FFpKVTVjYOCYwJALJqDbt9HzOznxxwCsLWLwY5qzj0ugw/eHa2yaiIPjg3
hfBzKnBtGSauw4JQVQ+ohz4qg00pOCmU7m0li56AEX0K1Okh+Rx3BnZiigIAMYr5
l1xbTRRtv/ocOLdrkvLgnxKir1QJ/ITerS44oNk/PnCBqxirUMRPlinT823V7iId
MLCmkvT3QA22meXVe4CwHiPGA5AGp+kqcc7/bkGgSoaz8W2w9ohL8ppCZnmoAtI4
9C/y1T+DUdtMgP4anOk0YN2DbqKGdK21xgwjfUDvutkJPOXtqYMU9iGWQuAj2mxX
DdaHC7qdiuVsSLNZISQj+osttYvIGLaN+1XoBLYDk6/ew4AAL3IVD+xHI97BlDK1
m2iPumrL7JHHDrlbW/5R1lXtauN49+abjkTolHls+yeaZDIkMlGsP0EvlFg5kNjM
pIvBu49fVN2fFN+PhYbVAQW9L/SXhPHYUvl2m5WPD5JcIiWxz9l1BsopD2tUWiJe
6VoUGorISR11hKIVlgohT5U9TNh/kzelcATbCTCq8FFwY4JQfQ+HRU18Y9T4eFgm
T2pZR8XnzXFiGKjllrVnUB5th7sruPHGKRd07DTDHAiSWONfvFt6k58cCsw7GoP4
37hf6uWwdLWJPWhJvX6MYsEAazK0vS0Ysiu1uvbqJdexpgqTVEFCHpcrdu6FUUFk
Abo606E3p3E4y+xWMhcggFr+GOqVfxRSsmRjBoMOJ+Kr6D2cz5QKzeuNYIRGIbhk
18+GoJOvMbKPLo69P25O1kc49P/MTqbhd8JlD/SI/Tch/bRz2FqV11Jb1R+E0e9W
mzYf34W5zVNuLh9P+Q+qZhhcczvM+Gnh/f6gQLHO0VP6dKrvw4GHqVFNlb0T7BKU
bvutI5AuuJo8N5TZZc1IT3xrGFF+afpXN+vEXKQAeBbC2cMSaVjnghMYcJBwVqNl
HYvfjeLmyzAdQpkc9pKQ8qMMHy1g+2cnAsBEVDtp8RoLF8OOdNmN/0uIqLh5bvdz
XBw1Jt4k94ZgA5AS6OHT84ULKUJNfgErODen/570tzLOEVFE9nTecTTi017EZmAW
9NecqO9/UcOFNfwXE23FR0osDo0AttMw9Ez+TS9zCHhGoT8z9XMtQ/LrEd0s2f79
vsRzLJoK8+A3GssJetaaOV7Gp6jSOh/4QUt68MtlEwou4bIc95V7udTzW0AhVblg
doRhvPaxuxlFHZR8SFDdNkRBuadczm7+s9gJaMrdDAXsnPcObkmrCKr6lYMXgwx6
4yOF0i0h77jZ3YcYmq6upixQGl7ds6ipLbPpqtewZbkLAaplIYiE5LtyykFV4Ses
qCRGOxunyHbKrwv91nCZymbw7RjFADDUlBVr/mBIvA2yXGJ7maAZc1I1QsXt85PM
rD8fdFdn/Evu2vcmaIOQeluWJx8g+K0EijqbBkwSVfK+VI8pAzrr26R80wx8Ze4F
q3CnG+2HzDUSj4MMnc6fLHwUlTAEvT/K8aHCgnJ7OjLrfvGDSK0WWjwsSvbtv7yl
V2h2Eyrb6kAtC73AffmdcH+xKiY4R9XmcJezWhmaDJuJQccCSPu1A2h3kBKXjGAc
qWNE9JMqNIimvxtHYu+l7qrbuXDzrN1AuUmqDrs50TxqXeiMJqjKBIbbp45zOYm2
14sM297KJs1xhyfB3EbVoJTAupRIifzYDq85LrYkOTSJ3ba7Lnvep878tdPgSK60
bREWG+tPqJGHVles2S9iPnH0IE91Omvj0x8kk2aGCa7DSvW0LjWIp+gzrGwHwUnY
Rd3WCmMPprJfgFbfDXCwV7F1qFenT8DRItjuSmKxfPTglsmf6qnArMRJAPQvhRnU
QJ9ylvFeGSnWiCLy3uSZdtiIypMDjXirESEN1ufgKx+j5Blj5d+zlUzXclSmelb+
Nbzjwa8r1i9rXL5+v0WyfJuR46E+uRmh+PdRXGS18ee4E9yBxsuiZVwAhpyclVZF
uCcadAy8ZcXgxo0u/k97riFbR70uLQB399S525B5bV5kL6QSgEEXI4hGmEGyUdkp
dTqjMbWJaECIJgRbBoP/4kzL+TKUIWv2UmKc5CCRypMGt4o8CdQxUWLvGhZuDrBC
zWghgmiCtrsDifhJ44FZl0JRAGRzkJAtu19sNeDU25ml+iBV2bfJeNxHBTP2hsNU
UZ4IhuFOQgpJTLA19CzkokAM2XObiDpQLAt7Atiu1iBufcMSGqXOTYu8HOt8Wn3O
8st4sQXEcVjgjPyiPhvCbRtaHkCodsouJVTDt+PZeDbfaFSat/Fq2O1QLYjvCItq
+wjpSaImUpjzlbWTbpVDKX8TidMr+nVtc7Nt61vNObHnADLuWuuNbcYFhuQaetWn
vM/Ef+zOpZVo8fGVAfq6kd/004chKZ5FlaGGclquv3vmjSKiS9RWbUdzq5caBvVr
SfCDQJwjOUfc3EEFXplHROA9H0Q/3/UuadPyiqq8NBq0RSxuEO4uvKSFrLYzfEv3
aXSYiX9inlPEiUDKXXVS+eQD4pBLACBURbvfjZtc98QxeY+L+1UI0kHHHHRonAxD
JeTRDEGQl7sFWen3cYmbN0ux5zmoeVpUcYIMMxego61wXmeD03nn9eoBDFZ/aTc0
J8aTszPc3edulXy6xoUuq/Yg0ia/Ddp2z5OyDtrWJolHpx4X8EWxSsSnAnSFcX4D
J33pEKRcenLdmdmmINYawlNeWB+s6sp2wFsXpEs9fCjnLWf4dX0jLtF2khufEO52
2NbVXuNBXMmwGpGnXuff29Em4KA89iMHiRfz/GcEuTjm4V0+qAtm0aL1N2QrlJ7+
UiaKQnVbycBhVXao8LeDT41Uu1b/nRCJ3OaehGM+udkOeq9R76gEFvyfyBiLm5iv
lsEcbjK/EzUSjArEbZ/qwvNiyxefUy/hE10MgRBmQji+4/F7UoaWcvroWnRo8qlk
+l1I09X5FSx24JfVvg0PRzV+KX+8tundXnwsoAS7LQh4F7C2yHzyaFl+HA2T9hex
sNaCt7rE43hROZppn6WMiwCUUCsMPfUqs0cfSp63APAKajCLUnL/EkpNlN09/0Dl
no+G7n++h5d/rPp3AJ+p1aOHiy7ULss0Dk1Ff60vI22G5+GTMk5n9q68IxirP2Gj
gVhYAzEKIq5N+RncEKsh/TuTSpjRyBFjNC+/9CGMZv5T+AzTEVo6Im5ZtC7FBxgi
CVMphGbHJV9m2YO9N4XNVLXRuVf38XeK6814p4Tn5oLDdVdEift7C7vSeX67pWQ1
JTPHlbDHb54KJLjsCDJtYUnMirdfP+HptwZwV2ilLehHqrWm2W9rr4kBTeTmXPQY
zCllW/os74Cn0JbQ+TRCMK/GT++ZwplFqcbZgAmq3yVYPt28Fa/fvampzcyXVBF1
FkI2462U+rO1/DiOPEbUC+4DOVtbaWVjSWEu9/GsfArhO2mVG2Zy1tx9DIX8Bl8t
3AgwxcKegfD1ln60a9jCycxV/20G/r8pd9o2qQVdul89PukQEi6cy5qPPii1p84b
j5qHgP1lZLxyM5reidZlJ30VfzlIqcOhkWirj09QPlggWRdQsqvtH5QkH35UvL9Y
Pk212VvZumUte+pzbPGmNq2BxxZ56bkdhhrD6MTBEKlU+My4RjI4uqeuGenApH08
TEC8+qfYiHg/oGwGiyYcYge+Wm/kZGmaz/O71+WFFaqLWvCEW8HToganznKfqUWC
AMR3skdBCgfdJOJk1ISIDpehA+kkGtAhsr6RT9d1mV/xqB6uSXmzBkLHCxNCJOre
VxGou+wm/GkzPtwguHkeOk926XgNzYlMD7An0HNbMEROQzUXEyPZXiBP8XD4tVpO
zwHiw13hVT5c4eg/trWZ902M3Gido9lkunjqE8OR3ccXHintj4k4HPVGdFQckXbl
AJxQdY+/rj+IL+OtZIVw8Vt32uKHXb/AS4qs7cn4jJuMRAefUjKc+3DXDZF9T2r0
WK3d31+HRwHH6slC6JBYB8PISj5VpMmVk6hU5WUrQc3RrJ8mJdcFZs4DRuu0tLDr
CvzfaJq6R8I+COce2OjB3r/wDk1ryAI3TC1za2br0WYfCB/uwXTGzMsv5Hnftk8C
C0igjx+UOqObKBNNYUIgIAMb39pfZF8gxCryx8rSfpH9cg5ShVnFeX3k2Mzo8wd8
tdf8bnoXPhFRP6UDkGaEEwkrEdiGqxKGMdGolVuZjTqPjvyc11l9lnb/rK4M1Y/x
M/haQXxWnYLMRG/j/fzDUJtZhIj1YDeh8lf6qhG2vYZM5PznlQlZrZ27lCG9tCCV
bZV9l4fyN3rwkgkrCMykO75at64pcR1XYLjD9O0hBYUvcFGf0dGqhvH1w8FH36Ay
xPp2aiOKrwUUlmAnHdZ8POngb3VItWhNu4yn2fsRNrlQoZT1k9+k+LvqsPt/Ztyz
qnuPAPwYW2nyt/KKi1U0sD0RCV06a5l9JSYqutZkOotBy6kXQG57S+NiFwkFpPGZ
ral+lTu/fXkU/yzKvu0o2+bBSS4UNOLQblUekJhXQR0BOMlPDXvaY0xrh0UxX9Ln
HmAizRx0Z8Vui6J2gSsyyFQKDoPtN9aVb+tqXmiWUYrl6LP5Kgg6zlCSbvimKtqL
KdZNITf1FBHsxhxdkuSP1asWP54YcRze6XGvZAHAW0fpFQ8vuAEdYmhp4JG4i6vJ
WNUlo43JHUg7B22e+BLfJb7NnYU/KijnOtvFzd8pdVmAzHM1nGiqgi0bEpu8x9W4
qcP722WwsS6qCapYd7WLOQro0T8WJ+w++GGQXHM4J+oc3WvZT9v3LYCPehumUCtI
rCkr9Oz5j2xznNWea7j5kANwsvxFj6H8Fc2F2TKyme2bpD/3ghsZ09auiHtrwiqc
Y2S4F/M03Pf9IDa/ZmYpgVWFDnZuUfhdCMc4ovhAqX87DELTCEsy1TPLJtg48NfV
+ztZ4cyVdSAvjh7Qzmo/BQnx+hFtgMk4m2hTDyaaU2zx4IDvJ5d0cmv3ifx1349F
cHnfcXpqX9TklN/RPALnAIjZS8lSrOSq+FOZWhSKKQreIiEXwx82BJvQHhbv8Npo
hbmJkPYEERfLS6vNfynP8SFJb+ki0NarF9b0MpQIPogQ844xuxbzz93Bu8M3nn22
DsNGHGCOadqFc3BiCGWPMANcBCAy/Ot0dLpQUc63PUBoo7doxMSGwvDNF7XUTw0k
X5RsWtexq/y4+1oijukx7HmxgC2kwfRfPBQR940wkPv2eh0csx6oGwvqh8lgWdTk
EnvE+mehhOHoy8HK3+xG9SrDTXcnyLyvMXjrtvoT/2ZicosWPegVOoVWhSpUMlBE
bZBm0TIVAGdUVNLbJEaKcSOAGOUC3AX6oDUa67DKxdM4iseVRrhtpRhOfc1lNnur
cpdrpUCQeXus+1GCN5hbkIuEDr/W7dLC9Fe8vFojKUEm49yjaQfF+x5eubf+9E9V
dKU5Qrj1+zaWMNspq/BmIzKCx7vrHKljhdFoggXzqlYuMhOaZW+THSWckfH+T4i6
nZSFLXm4OSkqZ/1m4S+E3UzUzKkEjpfu4WbWj4lAgs3TlHOGFR2X9U5+TwAFQUw/
w9fvcIx6foDN2U5P8J7j4ketefXueWaqNF0JbWwJPr0QRSn0MSHfQ6SpwRVEl1YO
FbuLt34NeMdxY9l6BUilfh9wAgavlqvzZ3rBt3WpPL7THxyvdzm2cL504vu2/GZY
W+VckAoe0x6tUW9RbUf4t4fgEZ43f17sfI5zIe85Ew0eK4rx86xVjHyTaQk7LOQh
2TO4jVyL5bHdTrqBKum2Cdeu0Fr9Ozrd7WOBJjbyCv5n6UexRMgtM303wh3hs/rj
ADrZyi0svTmsi5ARHnTkYYHoN8oXAhSN/A1md44pH3waCJdCxuAPid4jQ+cHHCcb
QJO4a8Gs13Ol9irUDcVh2G2+arW3aWN6wAPA+NiSy3GzN9cCVg3roX7uFpeVvYKk
ZTeDW4YnNjl675BiEs9IjjLXY2ZyiQ2+wesy+S1cOlCg/dOoPOlqsDz0ncmtNLi1
ny43TeyGsQBZNB5uWboJtOmO3TGGvZwso8AYX235ZlejgAojfO2RwaO3tjd95uDX
8fGdd7oGQFcVY1thkmBFjkhoC7idgRql1UDIhhPyccTGpvdbHonljm0dZy9icUkO
C59qGEP490jbY7iBRKLKHrSqID4+786+VFq7h/UARnG/zReXGJ+ZlA6MV5smHDHq
tj92cQI+1dnjftxa0jGKYPfKFA1SS4VOjSuhDVFwrscdFooO6BwcolSrMOSnjTIq
KQLhgTTSOxbxFmnhZZnUV0//72uRJRGWtoKMRx1Vi+5U/n816t3tG0Ru7onYilVP
dbIL2Pz9uUyG0zAiFWzfXgzVwRcqvJT97cDBQ9D3naOU0lx04vXYiJsaXhWjmkWm
6kbl2rtUJYGUGRTD7irbTTEthXLD+Sz8bzO/w+dJd3vu5NXKC4u98HlE18/LDFUD
GH4pPMTlaHHcjGOWLwEcT6Mcs++Sf92UwDpa7sTIEHb+Twt5SA7HTY14Y25WfTui
c5tx6kaUniAcq0fMNyKZm7gkeATazEPL8GWQ8OT1yWX8C9YjG6zDdekT+pKeotN2
h79VSuRWXtu69Mcw+5p25n8J7YF6qZyjaEdTq/g7tp4DqWZYhZNoVnyADYhiFaou
Xw8OjhHEWUdomUjL3agspioT+KlQkIfURvUu68q6rPWZQKPMnf3ohv2ExMyNrWp0
+SKVZ/pkAnE9c0clbVMT6FHh9PfPDBqOmR6JJH8Ekt0q2E3qhyz+dn/9FFZetDOD
cK69xxTWfXM5sbrSg8Yj8AlmIh9fJ4Ljy5EvYsVbN8mEK9dAOM6SJbnnyzri9H7/
9c/oaGdBzoA5fvT//dkfoL5DHWj02ssaqQQDhYz7y5mhph/MZYmcnGIVxzJgyTtk
39xOOrs386g4gwn51frJJTj1qgmBMJU38LQg7prNxuA0KwEJsWW8gxexeOJLUDcB
c0n3YozmXfLZa5v5Duc4oq9RTreihPd2cjqaf6LSK7g59wRySCv+Rsay3yoDJMg+
XbUxCxubi5GDbv7i15DM5E42kSroEJC2D5h8+2vBXTNDOje8ONYGH9YoHwb827Tr
x00nCdvf8xClOzfKar5axOQOI1q1NQVxS44MGvBnWLZsiJpoTxqJj0aEhdtAMnyc
qKqYb2Z1ui1i2Gtqwi5dbaQFw1Gl+sz2Vk+cT+1nz//ZfN6CPi9m/CI4PLOmAcC4
bt9KZwMLRxgZWjdbitcwVY9ry6VKr8jYtMpFhcNdlhJHj59yEs2gjzzNnKfeVVzJ
4Cd3QlxFlWBkDCqyQQ9qYbKHppsP5BWJMSByGzvQbMOu7kohzMW3xcxo+h8LVmZ4
lm36Kxe3G2UkWuwVeY7Vhuuxy1qqrb0ISvn3Ba7sWiDRUqzn6jkI7RHfePM8KXAn
bIOf5NQLeveqfmBkK8rKTZF+amSYqrimK3gvLX+Q3GLGCFCMJe0SOFAbbUpxmmpW
D3FxYGYCK1P7y6Oey1TQ9NVZ7iK0e66Ne+WANKXeuzeNcXcWz6AUEdeZ3tSxTsrC
Zdef6i7wBkU4zuFoySUn+DsuAVbfO8Lg2iWQ8oRCksrvpVEuKV0iGGfjlE/93R9d
RWVohusBemeC6KBIHZClWQNrNQfXLw1IG2bgUyTK67l4FY9nI1qN7+yqVdLbmyzu
6k/uRySSA/0V3jIpqdGgc8KsTiH7W+u1FtxXRah9fx9cHzKmh8MYwFKQFlRQW3tJ
+x9qdJ/lxc44+eG5YL8CkBT/JIzwlCw1BgQ2hadxldWcwLEXFttK3kvpUzTpaIC5
fueO/b/J4jFcvv9SsTo6Ywr2x1m1iOYCGRIhzNvsfgkxq0vn+x5J9InpXrhyN9ST
d0w+5KBZLtZm1jeBLiMSsD0ERMVGxKaO2bIQE+6L0YChrsukUbvkEMyU6WpMPnmC
gfRLsTFhQu6jpPgtqvgci52B2HWjh8hKioqov46hnqbFqbpH/jLN68KYFYnkiFbj
n+dkiQZvbdsvOkjXI9k1CEYt6q2iNDOkxBwt2eZQGm22T/RFS6rk3cDE8dL8K8pw
QNnlCm6jTxG1nWg/YBSGWbSZms1jk4yt9lyVrbxIIiiNvMQu4Qz5p8wlHLN59R0g
KDQNuf6ICy1tsZNwAKE+Ff6H+T+ZDscNsJfqMtz4AhjKhcRfuX2SaWQVxPFtjjSc
034PhtMd6hm9oBQrHGSboW+PsOWs2f3yqGTrnopVmgIGMr36LecdZt3cPkf3UN7m
sdGHNf5Ps+k7C42gvE3KiSqAVWxsZ2FpAwdB+fhvMwOYqnou8f2G8f1gt173VrDS
fJXXXyjlBJRoEXScLIGIb0IK4anyoYurg2/TL9RTnfoHoeviNC2Le2cwFbBgE/gk
ZY+6bCAr7Qv3F4WMwKlm0ZQBr7pWGcTdewhaPkyqcsQIV6haLDvODSc4A9nwY1DA
35qrdbTfmU+ZE5AkLqBaZ0hqQk7TXOxvlne7Y4GCHGEt16qLaaIiaYyLA3sdWW/3
oThdZJdeQMhMC6QmLrybhtaFz8I46s7XO16d6YnCsyMkLDEJ7Db8YIS7ha1RQehj
PCHkyhMz0g67+fndHMMNRqEABu3VPZUXweuqtyIGYChslIeEey1HgdB8njyT05G+
36HB0x+DY/LpJAOI6UbbSRhdI2W8XF8BcaRfi2mxVkvot1RDCU1UFTPnJySldSjA
cHoRdFOlpOt2CJb+N4g//qk2LQ84Ua8sT8tbdlbUIZyp67h2VjHxw2ryz//0oSDT
bicSiaOUV+YSYbXOpiBWWO4f6IRDR1O8MpRJ8sBiRL4i17dT5yq6WKwQm4giPmkS
w+SmgP/d/8wJv1zMhauLuKALQQb0yCo3jveclyDwI/rjVXnxcfWNiwlANFDrrrAR
9RLJkS0U+0GHMHvyiOzZ92pZ5COqk3Adh+V1iIqtJVZjyhpq5Ah362vPOztzuHbh
2B+t6n/ii3pOQdHT/6DVF/3x2/MbcqNhFaJywApqkVzZ/0Ebo9dsFryqYJITvdjv
m9dVsLUSVGvKodHaf+kAggGi1gyFd2ZOmqwi/oZy2s+PsDGululCDTCo3ycj97Ec
kV8ptIxGqVAlvGYtJt39HsbFVyVF3Y2NBq8C9BBausc4WLe1vsrycimzrQMKALz4
iJZ9xc36WyvbjCTTKahs/XxVxI282gSfqWTL1hqrCYZcr0HMUL6JHcjMJ6bvC0pL
/EjOboQdYNM4JfPMi8urVx+uoxXwc+q3qSm09QQo92ObRgU35UqtGDSCrLqDnLgt
ua1XRRrAWsr3KYzw9a6MhvVWTmlLVeDG/EGd9qFy85ugqZDhg7kY6whSzC/qUHv2
0A6JOdpDQQjUATpbH2XUhYf8/79NG+GWcBfM51yxJkIxg5mZeFKJsupB2nK+4m3E
yCFFT3hf9A8dT8qu3FaOk7LetFW+vuk3HGn9G1nlQ3qF3F9fS0n82JdWHVUgivpI
2gaODCbMD+wKS/tHXRT/RFO3FQOBYWVoJAm6IzdwwIKM60EEu+qBIbrllacZbmgX
qC7xlnlyd1kpz4KuwfdB1y9PWnzkwYGYXrh4S90VLQlAEdct3dP7TcYSdI4brH72
U8TRGeFMADpzKO1ONZB8FFcTgwTFDxBIBXNG9H3KRvwlFlDCx2cSX+gY/cQE2Mgh
0CmGIgt3QJLa6un5fdrb46xoCk6K3+jGMAJ5DJGYLs1fWLkZ1R2eY2KidABOdEFe
+UdXB3QRwSHI0dp7nMrlujaRMm6IPzu3SG92QJQKI/FtGzA9DAXY0/D3eT/+wgEa
Inj2bOjf2hdlEVVPir8u94iAgr+ZRD7Mos+xa0wl6WmH/ql+qzd93qVJAflmq39d
Xrll+zWQfwF6pmgwWlobmn81UyYX1iBBZ6mVpKaf4awX+06e+VsDRgPP7eWPX1WO
0TwtPBJ470PiZbio08BlvtqK4qIdctGaNch8SGvSXu6P03wJ0tS7Oo1ZGuU1J7rv
pJmx+cC4qBzK43vsAA79qnUiBnwwu9qZA+ydNJKcdrQaLBW/GbrIarSGDoOSENdZ
egyv+k67hBhMWsRFtQjWL3gpJbcltJmvyAmAXlNi8n9Ims2Q+XrzgPjI2DWIzxuX
iuR4Xhz8tZtZb+BeUDejxfryoX2r1ThG6w8JSg+N7aB5ybau/XhRjzpdH6EAmuUp
jmeywbj65sFhpA4pVIyLFpBeTtiX8AHReg7gpXFc3CjDg8hOT4Zhr5+hVhwi3Q/1
5eZ3QEFvDgqA0NIHtxSBOuF8EgGMxFMUQKAx8ecWWRwl6ewZq04uWuYwvkDNjK3e
Yh/wCNjw8XirkrY5ahKl/gJPSZUTmB7a/lOVbI2wlGm41lV9xOl3d1giabVV8KT4
Mgqmisly7AwCBKqHYayyqLCNlLsSssQXbZyED9jFcd/T6jvAPGlz9cB14YpJox1G
+8hfrPaX54k3jNWasfnH4yGo8OG7y9XPc9SZhBYq9M9tu9rMB0Pgqmc5ttKj/hiA
UM8qrGQp3xpkSCjcWDcKM9tBNQ0HWCPIEMOhlRvfYlZtump+CUXyfrgikpskHrXM
5T8/Z+a2qwfKIpzJJc9OoU9IyAdiwqgh/fMhhGMCymGHZAtWYxwj3KMqeO5KE1HX
5PBNEv0rYr7mSqqFZ2SVVv8v1n9gkwv2BsECXdyS8MMxywanb6ufUjJ2+3CsmmWZ
t3G7+cZdfTn1AdxG8tbfA9+fPxWcsELoF3whdwjfoYTIdg4piPtTnGXh23LlMF/n
4vEtnMGZgwKmiBfcoILNrVxikWMjNP5ebiWJDqt1CxaGnIhQrEDPybHthnhj6VgA
Dfk4gX544cDIhijcqoO2tdCsWpDZDXNtg37XRQF9ERlTMkA38ajCUuPbRYtHPjJF
/+PJxJMVgyRkialc64Lw0wpGxmbnjb6Pd+Mls+EQRJrvfWvyEKvsAUkasU3JmUTl
miAUiunPySZm8xIB5x/WnMRvCzAJsEtUurmUKjtw4Lwls2gIMMZaq3Dx2rb8jtrC
9slzRkOCYbuJTAD3vRwJkYsc+sgWDABCi3P30Q1Q7qUKBdt4cShJNrOtnbYoaVVC
DhRBllSOKTBzGTlb30ZYfPv72wqbk6MKBnLVLtvV+SCyGNG1hPAi0s9kbhkh78VD
kVLdjrNF7OR8PLA0WCG5ea133cSiqVTi4h3HhPtCMgPwzw2zDwpO6Wa4NFZv2PVW
5mAPsJtMycHvqhwfEOs7uJJk+qgE35l5JkAmvpuzhIkXZNDb6PcxMWrC9HFd7fhk
4S19tKokwNzNclkMuQefiie56Fds7pWeE1fzquBm3vD60nxEJeteyN20O9zaYXYq
MnmxuS75CMeV6De9zBv+OM3Nxk9wQY623uh5JY2ZDYYzR7OFjmNmP0Dup+iabfEg
1fE0dtmOml4coLNn58NzqALaBEHQi25BowwFKOiHP0A7APELUlPGuZDKvvhvRVRM
uUOFGo96j7dn4k7/vynpdEzhHO25rhDiFN9+Qegp0W3qmfkJEuXNoMPqDNf5tUnM
tNzBa5xUg5TAK3FyBeUqtQKdQ66pZX0zalc6K/KdZEf5h/bDqHtbsitq9vPqDRDA
y6U/cnBmucnSXaFgtxMLGJ6v3wgckXim4XASEbki6RRVmfpMZ9vsaSTInMONsSA5
rYn+pmwOq52NFfoOLDfABT1FMgtKHv+b7YBkVklee7j4K1gXslQ3rv2vbqW/YV/j
TdqntGAqepl25+kcVcMumNs/eiY2xt3NkmlBZ2rIsILlsG/4lKTuVhO6YUVyXEnc
0O3dgo712m2SQbAJj2NOsGfRsRkW572Wugt9osb7Tl9PQvNupdakWLAKaphg5sTP
vpD+9F9CthZOLG59NgBLS5jSLijGPEibWwu9bFByUKC3NCo7L0jXdSiYfjsFuePV
MOMUxvzI71d6s/jZyyZ9tDlP5ERoFxXVJkG8esr7A5kV7S8TL5+IgmpF6EAGd8i6
uJy5QA4okiZDbp7400U/u7qadVqXjm4HA3/c6dSibjpair0qc0wrI5Pv5QkPsF2+
ZbKXWAX4YZ5PvskM33MUnlrMn8E3thuCIaA7yhAcOrOEpBqDYB7xC18I/dG9sG5l
TZZtIbjdNCSoV9GBzm2s7XecjjzT8C6nf71ZMPEZ/TD98Qcm942XaMrSMbJso/Qh
FgzI0aZz4obUZQmR1wmZ4UwJzxj41BgADXv0Z/hP9i8UQ/XBsHjemEUIYj1slEtd
p2P03cVXYkEN1BMIdOqjAaPTljRo6hlDV6R4MhDgFXSYwCx/88DqwRcvAlOr1Ciy
HIr0oicr+DCdpyGFjdSuMla5xp3e2iRq2isKNyE0fkWX+c12L3G2SgEJDfYeiefc
ZWhh4OIW1Do2pnVn3NWM5NcA/FiDdSTxtFgw1QJsn0nbplpYtU0SEyN866/331tF
vrZjHWJClG8dJHv9Mu8ST46AgG122Vk4n8wUIqQP1XDxk0VQjZfQvc4TGFdKoatR
CqB0FTT9zEgdfJod72OrRjvEPQW1bdm4IhZC0TWziDrMvMKxrGgar+O1qbPxGHZt
q2SMPDuRoa+/GtgQVAZmbR3YECdnSRK+MPqRSwLGliwv9Vgvc+TnQjqW5FeO0FmY
nId17hxdA1HNG+20Ck2zwxsVzg+vT/ACiAjutlQ9vlGoiYsrUx4gtCn8W20MdEeQ
/o96HV49NMULGt22N/0FTJml6FQkOwgrYrdZyB4iU2+fm/mhMQdloFklfsF+kUxi
TzKn8J0HFMg19oVsX+Yne188gPCGpHKPqdImr920qPJWRSfVWZDmeOodsfPKSO8e
q4vuyCs3h7pAs9ATJqOUQA4M6QnI31LJOv1cLXuVIQ+FdWSGMnth4cgD4lNccPD6
79yCWhEygqUj+2ynDdhLdDFHvTD4tocwTldN3dZADFgfnLZl2Six8+1cSREZV6Zj
P4V578byCHP33qp1ibGynTpuyBbCP/EgpdN1Xs9afqR6MujfqmfXbtxulbcCuJTk
g4SgPfBVxID1mhiUEdM/BKbbp22Cr86Q7OqvJ01ZTbouKaqvsLgyCqTBE6JfhXe6
I4yenRJlOYncZY4sIUE9nZb71XR3hoPhhGsfJpsmr/ofrxIbpG+/2cVq1Dbdi2LC
UFb+8oXwVSlZR5z09eRRBi3LDEpKg0pKA4+BHvRd1JJy5O5Y4yvNSGGBje+VWK5f
k8IOuDakAYjfby6RDqdmSPzAQPBeh//UbbAj/7U2POdihckApaQ/Xna8KWC+wne5
LRtCF5+Dp9kvDjtcDhUgJPuYU9XALRZ5F0/1f0xxHPESBLUCF9xnoAZu3+ifwkvB
16tw4axQ5TBz19DrEGV6ky1mkAUv74ZPmPyuyK/cxCZPh2kgTQLRBhMLV6SmWk7F
ZwwmMBMdL8oDB9vwFF8A3OSmjEuGVM/amgJgHQShmK3M3PJP+PVkQIQrApBdnaM8
/kdghLacj5wgHdfOKafw6AtAOC2yin7NURCyxcRAIIdoUaojPNvtNaw2RGVPEMXW
WcTzwa/FYIlFcrY9srSlVaeSbPjYgT1TamszItiJmOv97CcbiOpbv6HUHZfrCP/o
APkRD4LfuepMJ2y72Q4iawS8osoRUX3ojOnilmOXxadd6wv4Th5h9A9NUVlqkvJx
n/Gi3cwLqtSY3ZOaR+zm+GIHKnJDPvUYPLYyWprVf/VplawHyu5Fi+B0gFcPQPN7
xNB3AyfUFKkcBH2T64hJMF1gscBwSKOqaqqts4DF6Rwxps4tuiGBFuU9F1zSdFI9
GJsPF996qwTpLc/R4aEFaBbkAHqe//zSRsTGBPs2k/3AcWkudWlf+VOuBQ4Mh02f
05taC6V8sbpaYqQdgeo0e9UqhEzOO7w5TAu3GaFVNeFRduNmlCmvEMzP375ZHv1M
RkAUYOuzTfTjTne56adeUwCguP3+LnsY7Jubo/6pw8WD2kCyPPKgoq4cDICozyeC
/vCHublfoTvRUXShr0fLV60NEXieqRSIIkpr18ZF47ONJzySZkVgElC3myR3cphV
XpkjI8tceeLBjrVzCMzK2o9WrDvqmetA4ENrjj5W81bfhmLgxQyQXhJ0TGzbA7/3
I022Z6HDERldeayFvWoKPQzqGEZ5d15/Ho82PKyJT7/eO21pSvgNB8ZI7nnnG2Sj
LImm0trcaHAqp9DbnYnCFX1tMRDaWwzySTDDpcEbRfs7URPnfJ4U16qqvv9TjkF0
gRHVWny9wzVaTVrwdNbmMZFno8Y7Egmjt/BZgJVnT1Q+W9hdX9nIyYwTHlWksw/+
aDZOS1vw07OP1NDmfTXEbot2n3c9VaJs4viZkLsEqE7nJk1Aqm+QOSbyNjGt8PYg
DdPp54sIb70w37CahDPMdOyvkF/65rd+R36qd297F+NjNWW2unXAQoIsjMZlTeV5
K3Zj6d5FYSDT5Fb4bls1Z3CoPRTffh3xlcvq981x0PWpvTVrhSlZfxHPhwfQtMzi
N6JmxRF1nTpMzoblE1EFVKRpOwLRgM8mthDg8v/geKaUjhWmDD8hkuqpqwdY0rva
Lt6grN+sJvG7j6KjD4SX6mdOuwwuPESOM48SBFiJ/amzrpdo4kE9Ed7zWKM7ejfe
stPwGVgH2zIKxSe+j3cOiopQ/K31Bazdcib3VcBUfGMG5o+jQELIbzrHvhJnYpCK
attpZmK8l8GI3pHyBWLc4eD3ZjrtxRIyDFn8wRkY8gY0Psdt83szyEDYxOm3AgnC
JtBYyi8KdmYdmFuGiYhFTFufPw7f4BQqPkElqZJ4D09cgBxgbmIToVioODP0NM+w
/nD3F4Pcn+JtqWYXsRhankVMGFkpXeD2k7kXEZe50wIq/JQCRjwESU0u/2p5TSYZ
eXIn7J4sWmWcRq1H5GdDEMPXm3twbDShpBjaNR3U+UlcI8eQ5rXde69kO0BQdhFE
8B7IalKP4chwdwwk2kXZ+BDcd6lU1Nh0h4M/EZ2iFxdXZy+2rKrSVHpF9uL+WJ9w
uZh0RZni7eAi/JChgKhP2g4FIf4YBU3EXpzbzMpcH68SqAF8FB7EDaBSBHG4928m
8sLaOSL7TIR6FUXjtQAVSWTPpBPzoI+AtAHOUKfDYlwmIs1alIVgGnlIGjkWBcS7
9enbR/AXlM6oeYZp9+tVI9YnTGhOfLspW/ynOW5A885d0LZBYxNUEjMhL1xWt4cK
XM0Js0ye0s6J/HxUU6OQPHTo+MU/Tzebf+PANwLq0VSimHiRfsMq2CEldWmqxJIT
vCEkkQHtnYWoS/bx/gy2ljcxyQwJ9Y0FcR2b3ExRRkCBEb9Aky2O2Pi+NojiIvGx
TbOamL+PCZ44cmSBWEO94Q3f207Bc9maLD2Lc6BvrAcJWEB2Gr5Upr7YPNZ81Edx
ufN2yXTh+aRFsaab5n3l535nqQWpV6y3G954BW1RlEhG8BMgVWYMb2ot4J03lAte
Wkdp1MiD1PI6PwRqEV0xpo5n8zAKN4PIUpiCl8++RK24IUFr9KCLxkmZVITp94T+
/AHHHxHxQUBHp5XNkPMCVmV4oWAMdjTN9y7hKHZMtVHGAhRPGHeQnQmvRx1G/xG0
k59snFb7Das1cmA2F7Y+f2uiBCZ7UdlPmPVzKNZlpnUvaAsMSWT3e6wPqiKonSn+
COuP1hUYMmkrhumLVJSqZHUjbsQCZ0DgBQPGFvvA6DcPDx+8zYjHeWbbs/lHDvvS
PBPsnwAUTde7Hp4mL+FTDkxdkcgRS3aHm2QuQcIpqTLJ365dfTQ+6p9EXZOJYhPl
G8nxw0KIfkseiRxO8wyaL6eVRW6UquYqA1VdmYgkoyodnXkXSi7NmqvwRdKN7pZy
XfInJvB4tzdjWBuawoCXk1eiL3Ju2soDbTYlQllsxMAac9njbxUbUsuJmAjtVwuX
22WtF07Je23zryP6MVsCMjwvk7jD4M0mplKR+5V1nU1Ws9AAi7Bk6F938ZAm8sEz
2sBboGLoPE5V5s8ebETG1SymiNGrCMrCGCkaiHPkUX8rKkux/8HXSDX9ARPxlSyS
n5fwf7FIkWxatoL2ND/b925irDuztZ+IGld76ix/qQEeOJtR9zgR/n5jhaSuSaGd
6WN1+Uu3neg1v/gIUF0hD1qf/PtBqAzveximG2DU1S2AjwiA2Z8jyVxey4cEa00B
175LsGOzYw+LjLIvk+tQ3miOfm54xWP8lStpn4eVaC5lMZ5qCWhi1WUrsKwtReLm
qrpk6xKOrN5tV60gkB0zogR3Cy4sfqGEuBXjvm4flUcCA8EEhKG9L/DBaj97EHeg
hFwcCZmdwDJXxa3colfQT+5IsiXSecMP8JW6SnJn/OPpjuwutpBEn/Tmj5lF1kHo
wUAsvFaP0vz0xrAz2Vx6fk3iHChCjhLk7GFvW5sc1cISwEaziVGhl8139sFRGfbC
KgCfoZLZ/9s05SfdG8TEGp3qjR+Tz9up+0/BMCYas2TRW5Po4SsnHpgvXlGcZ5Ml
Tm5b2NRWcmrUHlXax4QDsZO9dqi/Tg3uZhWhP9Kth8JQ6ZLXncR2SmfDbdlq+oPR
GFSTTpfjhMbVnC+lBdyx15xMqBIFHqUUD9IZijmZ4NFG0zx0HouzUVtVOIg7uksL
JApla/fcTbcWQ+6WrFRe7zm1uVvU86f2YgNWnTTzUhqkoU/lhQ8mkRMrPES8HHz3
7LALhRYBGwfwxkcfOuV8Lr3NBETsmkQM3wwNVg5XUHeE3vAOnMWNuxHgDa9+joDg
l4ahc77P3t0NT8kFnF0a+ioTI2/iIbKgBzR8g8d0amuFD1qtZFG7Gc96soPl3ODz
wCEkVI7+sAvC/3dCsn6FxolxlVqPlftzmLfKOnAg6In5lTS/Hy753XbA3AWCvSfG
22QBlr5drGHL5lzmFZ2BFrj+X/gR/+IRJQT5S/cf8DtW0s30BwheY/mDjzQa+HG1
iRBbb2QlDgeHCagGejjaxILUZaWDQyZmjclmmXbTe9hiTR8DUCTc/1gzD9882x5j
O8JdRwE7giBZawhtmdQjezgLwBFhqJ9b15hZ4zb/rD0UqVGgzKR5TORM7S45ecJ3
Ewo06tz0V9ZIMfnLAI1Owzv+X8bwf8y2wZhBYU8chaUPIFi91jaNKFUO4os8Krfd
pdvpivCRnVQlhaVmlCAj4RIzD55W1oBLuqDOh0Ws8q7LaK/68tgy4mLzJ7rz/nKi
8/WVgM9rbOrXo9zgwVFlX5LujCSp93iNFtN9xuvXAEyGdbBwR2z95iivjqHUNqr5
LsIcfnM24ZmhlLumjJoXh1vBL9lnI2PWPSu03dpxCiESSJqIjjPmB1Fzw1gnz/h/
Ph+n7FdfTMaGFUjSPTQmkeEq0VTtjTmkG4TE3odCu+RU5j63v6iNfbPozhbGW4Wc
zPRHb2DZkitmEJJ2kotwFe9vaYlQ6s4t7OqaopHm099R3RA1RzeXJrgouD02oe2Q
4nMhTlT3bgkrqpGIRJ+DW02XWlbo8NgfFlfJOXkFCQ6bkJFLG2xNiTUgN7mqwRp4
4VIw/NwNMW01u+Jg23ezddC7KL+4MsIJ/ye4ok3wXcYfMok7znMMvgsvz0lFjRoh
vHY1J2rf3m+QN+wRHeUb/OkKAcRnkPawkaZ7VqGxxTJC2AgAQpYICPtv6RYr22Qg
dlinJ8Pkpj/28GD4Xq9mE0psTfCowdiMX9MbIiSzlEZkJoBmuq6bOhIjQTgUNUrf
98+PWu7W41Lger+jSB9m0HRpHID3znK/+o3coTrPGM4r1C8dt/szsZDQoc6Pcs8T
ysVsA+/jCMXekwbKIZbMRNt8eJup017Vnk1eEkUGNRW+dOjIcbxRXjZtbb1GKQIe
UIAwcUDhb8CBMZcHyKhWx59mc9TmZ7wJJ2pSc4Bj9eRUQdTU1sU62jnLSBcF5h6V
Qw8Fo0GBsAx/HAqgjfUqbwzMvc8spUpOvkCLl/nEapshM1nkBbwh+1J9JOmNviMr
UkzAEpOlZV8FtvTuxbpMqcBmQ34c3VIuJGHYHmRDDHqivQ39jVo1cSZhtpBum4wU
4Ir/DAslKkxmzenXEvlkHaDlSezQ8H7XZA81/DFEID5rniwMK1zRmAeKgZdcVO+6
nqUSZBjyJxWs0420996tAW2qffQIImKfKQXHJ+gYvD/HYdhjo5GF6N6cgGB8Ag4B
8P3OTsbrH8Xdx13FHjyyT3KcUJie7AE0K4AM499TB6HXPHqEGi0E1VV9xMj2viqu
V1FkxgyMpbtMAVhaQEKjNEYU8Kw3FHC3bEbRFD49Pi7cMT2VaushB7WGetWj1sYp
vqFnSQNbZCvIpPb0H3apqenEVOUdH1LYlUQQsVW45rTe33ylGemj/bRJ6JCnAfXh
4Z3J5iaUXJhLnKnSi4qPDlpMEZKkCl1ofHJkDtsm8jI82u3ZENKAN9vjOwCwTvzP
Js9Vpc/VLGmJZuTwI9xeT1Kv3d1vztCddPBsBGi35MfBAY0jwV0hFeEEtbwX3yo+
9h0lvb/AXNheE2BgQngdC1KbFKERX9fNI2KQB2d2WunmrTdkBpQ1qqV1oH1KDahr
PeYhZRCfhQzljQZ01K+wJmY53Jzub9Yxmi/CSBw3xtOfLQumcaFSEkjHPt/hA8nS
w29L4YQIMn0I1cx+BXhtzAjLN8lhvURN3NQ/xZUAEQ+HQ6ZI8TVwsKS4TsQbefAG
9cV6YLGgD4gLb4M/5irgYcTFjJ7GtmbEPdwLbbiLQGao0YPGRZZIes6bBLOb/U1J
U2GnLLQ8gAM+1TmEDbcEmsQYen/qkvsVB4Dzy19d19tA1X0mvwUfVCqffYgSXAv4
913V9wLzNtjaEKAqka30nsSODt8J8HoodXhjjiKdwAVdohjLNRH0ZysQvIiXLpGd
uPpQDh5qJjDlhW/5pWbg/iuD0DU6lDRHV0Qbwf3BkLG5MbW2iCLsOMGtdb9AVr8O
T4Vq00+htGlWtExUbK4cbRYx+U5uOlK2Pg5sFWeQ/olpAMu2cLveYds8ExliCB1j
3vngePuR1NT5cYAkLxPtVBSCMrkFC36BvQesow1nUQ0kXSEotvxQjHibM3rulP1I
O51XkfyHAlPArOUlATkxGVnKsD1LasnrEiKvc4eJyRiJ6jXqjKn/cqMzADailxbL
iCTINgoaCJtlNmiaXfWe0NWKYqXBym+js+vzy+RWnL+qCJEsvqsYnB/TRc/3VMP5
qpuJyOiNoikYl1fgJe6tWbiSnKWY4Qa+VMdTsnuRlA+4AldtENPdph5v+ESBE4DH
EF4Zsmh7CiZmBq8JFI/W0xeMrXED6DWftFYdc4ZboDeptyVrTQt13rRaP/aLRJPS
qKJGHp4nV9c7Fduk+P4xWkAHyMK/WuoyYiEfIRYcCxwdZ8bg0vlnqGAlG7DTim37
QfI6ysGFXAdNTl8+a7T/eg6VsQper7W1X/+Lol1M7f398zL1tjbomRsF0QoBUDO+
iutyabe1C2b9OIQf/+YhoScP1mh6ah0z3OcKFfjHVuVtTWMo8JgBGplfsL5lNcsV
3Jns2xdZ5ahxgmsrWallPMWuYsSXKaNhrWP//X3pRahnv0kwYhITP6nulJmDM7L0
oWkd5rO34sXJolJE1a2gLHW7Og2ugWQZxOCctrJWS16EtNc6/cX6TBkjdgOqnXMV
/hpKMXCeX/af9IOqUpXr/OIafACHhqh3//06eebUBLR9BpX9p9P+aY9TxcPWjrdP
hDXoBCyiDEqkbPjQwa25pfw0QODr5ZVMALIWFCVrJ9ro1bywljc9f2hGPB1QhvpP
KozDxVn2zDWyBazAiid3gt5SUoQ1fhRn9XEpwZLYB2tYB8RI45fRtfFOe1lhu62G
bx1LZzCsTb80TU9NHHwPv1ommX03hqlOz6oH8NKV5AEDVRqcxDapjf6ZbM1q1t6d
UHI8lUnbuJNj+9nDKIaJzGu2SJuTpRe6wDj/wGTe9F1g3wckZgBdlDf0LSvmAzDc
+0zcCWIL9Br1RVzoffngHo7xsVtbEpHoixEtHLtrlPMcql+lBl5+JsDdZS7ueHKR
Y6t++TJ9Qn+qwORlnZ3L1q3j55hjul4zQp2EoR0tEmHP4TGJaZgDcCdoMmWMEbla
qXSR5vWPq6VRrRQC8ZcrsxnnI+EM3AE6kIM1IjmW6AwGSd7EwX0w7XZv3u/wgRfW
s0Pm12cLUcG/zOWW29sWsN5KQVj8cIhUJNz7Rc0oVzTGcWiQ8I82tn+Ia2g38Dh6
uk6cT+y9QVUIQaA8fEe0wrc9CgU/MJ3NnWff0Fb5Zi5Givl6OY0NEe96Bj0qtUNv
sf3wgZBQHrHFffLZVijrtnZmWGC4/KxcMmwlG+v5KalzFAWRhSoTn1x5vbjr55oH
RuA7d/aWfmYs7SPnBQvA5HDRcLmVbr9vExRktDTqk0grOo0P6k/6O1XbYznt9ZDn
mB4P7x4nJOWFHAT/1g/GRqvUDf/Yv/yTNLQsX4rIulu4hshjEH9KZsGMbyoUt5Zm
xBteagcsE8ZVfNmxQHpU8ZEPBFgrxzGktWrntP90iew0mZljlPQQYI9fcXpV1Tc6
SpLOZWcGV6GfD6hrs2vwcRsOBJ/fJUr2aXyo9tSthtK0HPnLWd16u/B0o8ez1Qgu
oimEOx5Zmh3f8Ua7UqWBDxJGNqIbYts10o6/P7CwCKCs4pq/BOOEYbPypxik6b4X
aGkUomgTVcuzfPgR9a2Cp2rQ5YBJag4YqxkHMKsfFOBkYwLVpb0Eu4+SkbGtRFPB
xEwcy1HzafsrIyrotQq/F9JULJihI1a7/FdMK2LVxeyATku5TqwEpaghsDtv3LYp
+Nh3lSZfPwDwm8Hrhw6jzLO6y7EGYPvjIxE/l2uxLryACORLUtekFYbntRlud9DM
1aNch1wQPlWa45rYRwjgVao3UFucroN+LxjZLoit4jlh8o5etBqrpNngE3ccZLDG
BKfd0NCKJQwic84e8+gLByPUVpynNQ96LXOPp+ROrqCoxLb1OcmlBesJBiKfReye
IdG/sc4VahPCVuOEsqy0h6LxjVFhf+MbvtZpprPBnCUZXsHPVWH7pr40xRvk3+jJ
eXcy2D8Mjz8TcMdeRcuMXuxiadMPCfOfdfK/V0KYSP3uYU1klkkJfUqNZyjOSiTX
adcTDKifRLQqxEozvix2ECHD8o0gRnbUijoeaWt3leL+lzLwmZNuY5eMFOcBA9BQ
ab39fCEewmlfHKkLo5JjWtHdGlU/K8v7v9KkPyJxL+P3+QJUBCZEHn9X8x1gSAfi
/9eoRuDATKGBSMoaJYq7AtxTPsBTRLnSTNlnoukQ53jRTwxjTz+ovkSzj2Kq9OFG
1Xzk0yG6ertuhTkNAwLf91cKaAUMcreHhD1GZJF53B697qpYZtKYVa15pDQNBEEP
iU9hay5pOflijuuNZDhuvfyEFLGdxodEE47dD48bZYihro4e8Lg6bZfUf/2bBUnW
5UckLhpFZ7U0ix35Us1dQBxzA2PnknAsbscUAQaeAeVJ/QuJ2A/DAOMlshxqXMlt
NxeDxTs/AyqYktAWJKQ4yndKDKI2xe+DbLQsM8PTvjFnxRmrZKeXGAbYt54IwzQW
qHbojQCMeUohSisyoLUkRDGPFk66gCmPsjoAqaqjaIJO8KytQI5yqqNzhPrYn9YM
14R3SSYCHXZbk+lBwmAG9k3a15EeJMBJZgENZfVv7nrX5YBWxmx+t5Pk/Rk96FYX
eMWAt6izSBy2r7W1kQnidvdE2rcBgfbYdQVC6O3cwUsCSxpeUu4t1j2aRz47idEh
GhDjEF+uLidwUm7B5aRAiCdtIgpcL+iyIUyS1F0GqNsH7SLSAUqAMqF8UJXEgIFV
gCR5yPyTbHZLA30JCRMMicIZE+atYriYUtCxPhGmc3kzwcdXjAJDpyQyavr8ui88
69khQY//Ltd0NXYYXAmshQyqlVDUaYaGV13ADgPUzH0CF8zpiuw9AtUfmNw008u1
Ojv6SGYK5q0oLHwLkawEM0vBv3GLSk6CxBTN7y/s/0xVrrQieyZia2CkiRLc0e9Z
eNO4NJy1yptvzkUdoBMQdF/G6bl5b9Mg0NgMdSQNZdcigsFP2VBtgToZIDmG7CAg
xFnfOsoO6+h6vK3dyM6g8+T/dg2YjS715EqCjMnnTkfI1d9bokUu3MXjRqMhCjTr
RLZbYq9v6xfvjDLdmuhW7vXOHVWHIJctdxTXIpTVozRuY6Fbdo2J0L+O1RkhLHSm
VeZriUFUSZ3UoleoPfJY+ypE8Q2J7GnqWR19DTxBh6iJ19hoQnX5wi7CzrZGXYwT
+IpWNX5g0gYwUchH2aGWC25yonb0Svawmd9ENv7XkgXA+D696FIyjaZYpjKt3Ova
r+zW2E5WX+PFo2ULXhSdw3N1a45bXXlab6LHf/gW1HeLnOSecWE4tpH181nIxcQK
BJT2x7RqPbxC1QcX6uQDRwGQmZukykBJaR/sKBgCIUQCAQOiKCFvzfg15oipI3p+
5cF/a79jg4lEaZ6tPFVm0GE0xvLYPSVS/6YXU2YwVtZvd/3Qa4EZdp8T8fQXiADk
G828wQhnKi9UItGWVufH+PPICMSARB8VtZ1kYESTKUIFSBByDGjHXTJ1eTn6w/z8
fVWry8u3E3UP7Jkk8lRAtSjJdeTeKdrlp8XqoIzV8F26oMOabqs5mdFe/ovtRIju
g2MN+DtF9e11mvChaf809ZmjnZDedlyBG+SubBF77Pu5nESpFPHl6LSNY0o3JGQ3
2CnmMYhxEC+ABSWhQ5JzUCiSy0J+Iuq2Y8MG/6nMGFk2yQ7UERCsax75eQs8ZDXU
ectN4oszcfAQTOQhknwv5ExcVjzKaLXi6IksBpOlNRhfSKBayvUfq3wfMwNnedys
fxPP67iKxMeMKL5N6cJnkMOtuXUdOB1q50/q1ovnB1xPLMV9/lhU3CU6MsEwV44r
S+Ch+NaeK+RJxcAM90u3nD1mA0oWz0PG02G65yoZ12No5GfWiv2L7jCFLqemyj7R
v4AQLzaFzJ3sSLZmJdh0amMaetaMnWZb3I3Ie+BVqYSpn8WBLkWYZWrfOEvyAkoy
1ZC7mqInNNDv33k+R08yNmOFqQ9zlBLBBXnbs3JUwSKntNm3Jxjb/THNozK1JwKE
6cGaU2AlOOOtJ3pKd2+mJ0H474ZePG/HgcZuwOisllKGQMTJwnNK5f63zPYGnRGY
gwBlc1vOj4kaC76xuDK6TzKHMNW24rdeCOtUkd/nh1q5vhpvNSTcJ/mwxRGOjaA4
0/j+KRcAGLym3DHdVrZxYgDF7Mpj97dwB79E+fsNLlLVwldxCJcvR9jdFpsp4AAz
aasRoguKqzY2icEourqImKFEK3zk4G20ZvLl9rM0HJz2HlTJLIKar8tkeI3MuyBQ
Okd3GGS6LXrVwsG3ATQFvGeoZ4m3yuR69j099rcRb0+06LA5AxYcmrmCuXVQDucn
ftYn8QA74Izi0k+QmROIYlkqMdVmVfY/VVKXY76DTt9pz4RwZ3g6HI8iIjFkeeq6
JZZw7ntptAYqz1++FMe1YIeEmq6KLyWh5PoX+F3sdHKqu2CbQpEAG7zBNRI0Vl/W
+++gHP6/VA4wBAIl0882ZbwX8Sq8BWob6q9RpMqJQXzfEqCKTTFAWSsi+oVNhC/S
y53o1tBihn3vbwAnSILlwivutqmbYSlNkdJXl8X+MM8/XGFkFLyl8hTXAFe1tLif
1Z0/CPu3LoDEb2/J18HkN4btuXBjcw6i/30zkv405i8d2L1AjslSQkU0hOGXavld
inMSOtLGweKgs5U1P/C7xO9NGc5Vn2cmXqGAOOl0MYldffzXEm9M4p15wF8rFQPg
ehuD2mhQF2IELDhS3ISn9UJhjFgipXi/u4uoAGgpLnTWV7k6dU5KhzOYwhbBVFNa
lRwRz3f+pGWZ6s1m3bf3OWxzT6mAK7/tzkBmRXhb10R+Bswd1WKFsY1RdsLPAye0
NN3c4ShBE3EAU+N2KN8YNsRCfasWf/GjVIiI4986p9v8kMkY52rmuxxw/7pJP4ZN
5YchupZl1Da6AeH6Ncxwh28jGJI7IrfmA2DZYqVQLnhne1SSluRZAog2CBTNoq5Q
FThlg/safkV2hRU4zZ9xRLzbvqH/LSKj+bfEv3t1HxJLQlP6w8jPOTGm5Sswm5/V
CF4ItLFhrxNbWlwrI0c7WjYKSXNzi7SiOfEhLtMI8bu9m9Je040ugZkSa74g8e7c
zK2sBIInYqbdcKea8jgc7K0LUgkNrpObUH5wzOnQVgC8UlkIPa+MXK4MCa2Q3URV
0NMyAX9fj9cACNzYXMkfwwZQjwOU8wuh1AfRVCc5Unqk2DSKeyMdO9cQpky7ldkk
hWNAQorLRzTYAcZQjKWFwwNDdB+kwBbWHz7+yTdh7gyCMTl+jVyi2t/HEuY2OnhN
/X+BFiYxgXBXLTPmx48GHiuOu+yoF0wVvZwRPa5BLKbVIgJqeyRM32cOdw57jpNI
KL7BQ83WD+KKnw7qx1xFdkFVYNnQ1IwvfdP9jaoC0pj5NK3IYjAorHHNtGdHOIxk
7Er5gXdvGWC57pdlUasJJXm7Ar9KJ93W+JsRTXDhfGFjiwrQYCTckOWiB1jcvUpL
rWEDVNv91IzVm0uED/DWKbYhT2R+qLQSFpWuzPVuVcOEetVdo/KCdyyr4J+9DwL6
x91NSebF2q+8Ssv1/HJtqKedoNs7Axni2R6Ynxl0yYxxKTaMsHvqHflmmVHEyuwh
t47mTnBLAtIBt+tsyAvDPk7KRt/85qg/5DVWEKoRGVzD5ZHFK/sfhY2B9I/f4Wh5
kKsah7L0BetafCY1qwdtEkU04u9UJrwLPYiytyw3p0Lcrkw69P12JO9M/oRc2bjT
gMn1RkLCC7Kfi9bLERKL2yF7p/TM2knHm6ZgseLBrWp8FyQOzNUfBkrmCNFzndhk
Tg+xIr/RokLEtGm40FYmdd2VL8WIaklbSL4w+kfUDeu2U+k9a0jZ+CKTL+dPoLBe
zKDT3nh/DijhmZeg6mQP9KI5UgKWcUFgTiE7KZQGEAdd+Bw3JEuQcZ109HcMg3k4
fXzfTi/MblDIUaNi0Mae2Y/7MiUb01IAKsJzu8L3Mqe88yhJwsC7xv49et8g5vh1
clI7YBoS4V9AQY2sq4+EZG4+EqmOUyaL5wnjFP9ORgCVrN8yfDF7zCRUtBp3nkBt
W3pXdi+WB7GvkcbgJsvhOAgY6qXgxO4t7R8bEh2GkdjFJj3lDnWvmVUQTpzsdMmn
r+iUAZqF+MDDlJ1Nb+Gh9vaqG1dzAlwRDqDJswmjr4/OnRSV9POL9HKlyBvMq+2j
rdgnsgx0JeW5sL2nGMa6iuzDLzKSg+XKpXi3VwH1u2IAtSpO8iH+uQHvCZnRiYpj
bwLEBerEp6a25OZ+w6PM+80VVffol2BQvyDqmH7Ccn+6U09Hk/m+3BsYga8iR5KN
AcWc2IWcTP9Az4/btu7c8VgF/2GtnWmmcerUiknQ+xPD40kzZULCf996ensVixqQ
oY/7AWZ1f09NXMVZk/Qe0zZF8mNaxTgwyAxcr+L4iZrkF+lWI3hnsoMNl8DsMYOf
MvBOfLSAv+hW5OLrSZVTD9pHp/KNPxkfIHi0XtJQvs3JKTv+bizerBrAmKsq4974
mQFXrIQdWVQ6c9Y0qlkfsJmu+DM+2VNwzhvxl/Y9KnqUbYq7xOTdRUn5MEYCv1Do
8RCR6FVb+RGBBgR6d0IAqMR0BSr+ntg2JEdQaCkbRVjGWAi9D/83opJFigIj5D1U
TVrzogIuvFFl+YO3LBKtM/QNgrRUcibDZxndKhNnZ9T0QRVJa+/pPU3i8Y5egBje
GP4Sp3DnT6620MDj/tH2BMDueMowqWxWxS/EkdWe8HlwiV3UjRs9tVeUDxP2+WkS
UtN8tgwUTBR1bV4JMsyz9xY4/+zHazyp2naEBol4H71nacCoLT5/qIv9iID/8OOK
BSCRoRmU4zYrLDa9GAj8J8PKu2vJ/uUZe5BQX4WPwt6cbOWnCfwUqnaLo8GZrpL0
mglyV4B/Y4rNLRl0FVH6bZb1SFIkLka0zBHFjXpmzSwsbH51yqCdkhVTF4iNoTfi
d/SiAQSAS8BZeDocwkD69IOHmmu0W4l9Q9gRFsV13kq+uyW0KzHK3AZxdWSMEANw
AUJqWzxQvlRzq2A24SNAkhhaIE9JoV8DYZ5/8DKWdSicM5bori26VxYSJ5TKLn4J
lmF79vopbBWphsqOAJYQdN1pCeiKvU9JLVljQ6CMzQ1U4Thho+UGcooRj2dgC7zX
a6+1hdCob9LOCJokaZrpr48AwluEmoL5oYTEgOLP9iUyVK5rvkxyYnpB5ugwz8gM
J9kO3Q+pi47d11i0voV2SllhvsK/oEBPJ8lzdg03pQsOFySUDeiPVzOECIlophGs
r0w3HE22ESUuAbB/J2KePxP7wbczDcspENb7aNWHrPVnyQTzutkXsITU7gSF8Izq
eY9jwWTPs9/PtPkHClsWT1N8pnLaXFydxyTnHaJjVtxqHzWuUUByac99kWRHmijF
i6hylxmdTdTxOyZNHC1tpn3e48UxBXpKsArec26UwGqlteJTvS2O3+mcQT+FjGSP
89cXSxLvFPLEF3SjAYVHOmhhPPg7zPTnXolB3bI1jNXkJ1iF3HL2edjKF9za3fnm
TN2KXf6Fr8Wv7yfmslKKz47VclTZnA+lU5DZ2eqwJgrtam+11h07HIpGgOqdhiat
TDosCzx62RslOSJbEAqyGWi4zpB35WBMAxsj8Tk07/g6xNmu4ML2PFAGvQD1N6Wa
sc1HqGjS1IBC/8Q+Um6uIewo2+Y/riQNi6iU2pBG72PC3Y1CIaWgwPB7l4jX59xp
56MU48v4VJ9lOKrMp/7DDwgJYrVBFAZKyyYsyolFLFP60bwxSm8RD22sEt7MDZYb
cq6vNg3z0yLXcYlR4uUTDZsAxKPBj6DftcoqTCG0LS2HVW9GIZhx/9UKAw3e8hf6
a4fqhQczOi1tZUaLjh+pfkDqL2u98s9GRIzK2O9LTRw0rtDhV2Yncres8ofKDtmm
mO6tFP64RGP9bKsZ+kaI0p7gdmklU9tbCvcL4T1Vi8DS2uynjlP44dc2L5RRckG/
VDe42WRenzPbnekfv1B67j1Uv8C8ymcMPfRtAcI4PjpGOiYzHZs9hHvafcjsBrev
15NFSq+Nlbzup0Uid+Haw8OxMAOCVHvoxiPvDhEunI6e8iqsHWlL9AMcwm83JS6q
AYhywei+phKnZgJeVc1g4icuPVo7GVvky4+e1j3ilPZt4zjDFWk7Pbx7XkdtCoY8
Qdi8qIv+BM3y7VgUVFjlwK/hRgMjjsP6mbeZSPvZc2uMw4wuaLu3WVKbUH/++QNR
/h3QJQm8qZjvp35+LMSc8cZkkaUuJvuXtxKn3QM5SawHaUMTyx/2W6PYPbWk/or2
W3Z0ierCLAXIHxHYDthTvbq9XaSGnVojVCjY5KJsDWq50sCE4ofGblK3n4USE8hm
w2VZwmjwe2WFBb/so0JXK0LWRzW4Hhw+TzF1EEvGpybfz9MdCQkw/Lu5IkwznvdL
wNWbBbBbLl4MbCNkWwFulLKWEcixQqVPgn7kRcehnp3KAlTDaUK/mk08C27S6B4y
prCHqRT4S21ABb9fCsymvBeCgvxaDtX8bRCSJ5lSUDVS0BVANufu87KukPtndpbD
8+zKeJQEjNJUguIIN0TLHz8QUWXiY2JzD16c8keA+d2U80UFJu2qPAM41ZM9HG0J
jxVX2/oh1lumpJ20S/Nb3b5Vy3IucED7L5jcXVhusU9aEajzNNIRJoRlQXu3MwKc
cqLEzngaCu/C/vXz4F+OBxLolaxLjtYd2t+RirVyvd0gJNbb/oYZqNO3fEORO6KA
AO0Kw2QwMUwo5pcZYT0Nd54oKJHzraJ5lYTycs5MNP3fw6GMajYFGANYuh+5FpZJ
HiLNN0RAZDsWyd4ftxGv00B1zO7e11Oi7zGTxVwwO4AkeoEVLfpEsatsDxUBCOqb
NyZrfv8k+fo1Co4u50Azd0yueMn+biapYfy5EdG5LYa4gCI9EgM1Y9/sVBl28hIF
kqT80PwtbkO1XuESMG2hZXaSmiQfEtcK6RZ2Ke2QtiG2W3qTby3/2VS69jtZW/Mt
F3oeM/JINpJq+5EBfZ3c57v4KBhJuL71/LCwvMc5tpaGioJB02xjuT0OGO0duJcj
YRwosH1qM0cN6b9WK2Tgk5VrzR3IfFlJK2zSxviZTGT4/k/JLqO4eN5phtDe9Ft+
aayd40cgeNk1gswb9ivPrtYWQdt89T5xRJdjeCordzqh1TYgWrF+uFnl5107VgZI
fU6xrzAcxSohs8DtXvo3HZo7zumS6Pk/BhIgugavW2vUldfaI732wUIun8wcC6aS
A3HDFFEn1+FW7vN1BlY0sOBbeVb/sCJQqcWAqdUymTSwZTWkLZnOEuH08UVDPd5/
kxfMjwneVnmQxsv27b2FNi/sBIGDTA+QFijEdXk6lyJqkL4jXY/JIKBtg7u7kFhz
u0T7MlPFJAm60JjA3wTcHdtNn9U6DfooM1+ZwUfvvFWVoF6Ia6JQKnXs/zLf1sTz
VsFOq6RescZ3WxDLwktLKmwwbwxcM+ir1F2IcHXRi6wkwhyyhcMS97/96/uXooDg
kFHwdILNPusJB+ufNJKcDfslLWzeGS1guF0oUOm2B0DmWzbRJU9tJTQkSp0p9zCG
w9wzYem49qqoQruaGxpv4baFdK8QSyF0F2dM64OLpzRf/VIHoMJZeDd1lnOVy6+D
aGH2G4EC8hKtDAzl6mn95ZeL7F2tW7HeVi4cxgRXqcyu21q1neQZy7ABbKHgJNHB
ZtGNqHDY4t3guKkdRC0m52wT3YfGnwOGBFOvsHNgIT7kJskkDwqq/eepFOLzhurc
K/5tVejA5bvsmqnrP4n0YV63LeieKnKdfSzm2eqbXP/ZWmH3nC4TPcsEo71GIlyb
evXx/Cf3IJWiH43AL9ou21rroRJL2/Eq+uLpCaVn9FhX4hzEbRvgMAiFWV5ktd0A
nAsZraqAS+sGcDz41NMp2mOE1/H3NhMnE4Dh8Z1/08BsY7wCMrNI+bmcIb2yNGJy
4x405BJMjWw+xhzwOJVFFj5ekuhA86GTtRpk9AvG/7HZ5iEUT+9ATtnXMrxCzUtR
EPp4UMrxWHyOE6TnprzYW8cCr828pfmyHjE6D91qDL2STEusLDBsVly/lDeleDQJ
wZIdrC5fQhJolAkn0kV4n/4TVqAb7k9BJBMu2EAc2jDUTbK48RRizAeBWV43u36+
F1ZvX9DGuw2C6wJFU+pP8Y9ztKWezbsdN0rTByF6qFEbsyyj9ifEcP3sRt8H0lT/
/T5l0sW3C+q3mkglgxGm3seot4GrkoR1+yZbDw769lTzPstBa7zkLGF/oCh9GMhz
Vz0qzQDkGUePCuXjHOv0vdgMad3X2Iit01yGVYubb6J9MDDzQ3QmA8zjrC9t3K6q
r0FIgYI0H9110HeZTDuCQn0qUn6aSCLXcQjwbrKCvDnTvWMAFINctZ8VT9+HLFIW
4+gdxlCaqmV0xWLz7TaHr4itc+MZfZyGJGRuPznLmLPSd2rj86ywy8Cq3+zAN37L
W4OUpJUYnsW+BfZXq+OmY8swPB0AwrM5opNcKvPLaEtNGeHvSl6aGIJkqmQSCak2
FW6CBD9KuZm8RW9w4d/SUrlAt8ZFj3gxTduEishJed417kY2BhG7HlwmW0tJ0FvN
O7F+wuMwU0xL+zeZEi/2IisJ3js/dlpSJ+FOVJm1RLrmpFLtLnNWgoOw09+Hy2Qq
y5VEM2+C8BoqYk3Z0wVYShAujrqL9UMR/f5PJTS0GyJU6THh+Og8z3S5m4l1Wy6W
Cdfg14TkOScoy4EiZF8/yPncpELN7iRdBMkyHXzTExW51FlgRTrRxNEyZDG5ZMub
haN+rkMqxK5mjgGKaX8LipGxAJyo0dbxmm5vo/tgwtXETBPbQVZUfJM8Bab5EhHz
j9J/5Xox1l6edlIRIm5P+kvbO7XXRHYXy7J4LSx/4Y8P8Vt3mfRNRGyVkPB4ChUN
8TbjF2Y8dodQ+k/M4Q1bNRRGJ2TKg6NhOv9ugTa8jPMWksDVog61NCzfMSiv9Rau
VxudHwz3kdQf1GCuHfNoNcMCX269wx6xPp3NQItuO9rcrwDWCHvIyS80eHI54mk7
EcXGeGi6GaAhh5fYo9S39ko6agk2Daixb/iiirTZMOFFkfb77BybB7o8+bTxSgws
HVtEItSrg6ZhaT1zO+1Jviou2+SQl+8fmE0gqjVh2zy9p/iTyHrg/Y0AYLJvarv3
xNFsWhvYYEYm2fIUwKTJo0zTVdp64gh53M+Atma5ijTFMDjIjnpBiM0v8jus+Lga
/j+xrKWDEc+U7JEfqP9byQBIbgWEDIu3ofAdLNHu6MdnGb0c7h9WRScO12VERSbp
PyOGuBIp6m3b7YdglteAFXJhC5LLU8v41WiMMBfniTdoo3++/34h5kNpi5QbUO1T
0HwqMMWU7g3xXMPzlRAWU4IueI2cPH48QZzEuB6yH/X+FiJz0bjoWHSaLiDILQK5
J0exN/fkZVVjrOL/O4+gqVYnSKE3RlnS2i4YzDWynJGhH5uch7Nd5svE3DfXJ6gN
yhxGm5ngzSJGxu+VCKhjWS7FGfArZyCGr+n7TytpjG/W5zi4Ua98EIQRjYT2jbbc
hs2JX6yYT0Y3IKJWMoy5Z4CvSoVoouY/WJaSO9NNp+fzHYSlY8TUSOTpA2dV4Zhb
l8uBaWOsKYBVwJcD5sgizAEhNMFLU6zFcbdB9vAUvmnxDeScQHoSe2LpQD/YOg6a
doWfFdfQGb0KwyL5jpiDxk85qw1qYWzu40tGpevLugwTw84pfzgWb3xEThJ/QiC9
LoDEWLGCOYRzsLx9zecjfVMVV3gTgqj37MmusaX2dxUAR1yMde3N4BQq/Q4Zi0Ka
c3w71djf2ih71EsWcYf9ZfTri+wsE3j4jIu8PLkZXW3nRGomVRgjnb1AR5891UyH
mk2Gf3JjyFc/8f0nk7buhJ3ApEicwIyzARENZxnBKYGjrEmYSh89U706bBiAWeBn
e8139ANixQGya3GtMXnOjuXREwj45XeJPVJWOo9giqmaAGA0MX10RQ/i4qtE6Vf8
PMvQwmEuxyQwEgAqUcSdSLsgbIz1M8aoUp5KAnzZP5eFqNSEeyCSOWDL15Mjf0sL
GcENqeWEj2P4uKM66DAEoBBghg3oCWB2rAExsXYL4G0pJ8ZkhTw+86fuPrrBFIkV
40BY6lRKyrT0tK5QyQelDy6z9cX2c95YE7VY1N0wXjtSeReBprKJmj7IsA/mcHoA
Q6YS2yKM40F6VIxLwUZZHIvvtWSPmstjWIWEyDS3hB8/vcJ16rXu2S/ol5jv/Iv2
1j+ao2qAiY35mXi3xkbPjjRBB4yN4Oxjee56YNereVWOjytJY6BhyI3IIjJkUSHT
0c1zYHLyDMPLLRt9p5EF+oABvXe6Vz6LMftJymQXOCl2CVVakrY3NuIs/lARn0E2
BpmsiUcfTXsmOvze6Eu+Z9mg0FUX7VVwPpxbiyLWUBXyj4E6zxhuUmF2QfAd0o12
7rAdn+dBbCwobdWmQHi92vavBBMTAxP8lcYZujt9+Oevw7aCkfGQmXqe+1BWbpUZ
kmbk8pafMLgU8L5YNnZhzOJmwNbcxQRyVgFrCHW1uBGCpetvuf4lgIcBluGoIAcK
NlGAKb3nGrMI1qGeoCytPU44KkrI2WxQpZHKx5VqGSbQTeVTT76LSH7slWQ6IE68
PQH/tAQNhGNSMmuHRSibuujMWhVJ/N8AvCkcZwTe1XE3QcknJZ6mBCPOvjJkAyyg
OWJIbB10B2figMm7VLxGoc2foz4qK24Wc7Zq1YbccLF02OqhCNet5wufux/ncHcq
I4i3o/MTLfi9FP9+HHvV7U0jIHBTpF8X8SJI8XbgZIFtMqugxcFN84lG87dGYBWo
lNymXM52LOW5faWBmR/aQYnpke94qR4Hxyp6L2GjZ+FCQfucmP2bDfEmF7cC63+o
xatFCHHIRWJHniX7k+82v/XW01L0QQXuXm9DlXZV0vjbp6L+3L519fIgEk0r7WeG
tWRme6B69+6DlFLLiccHsTquPMX2QBNq+b2jwQYsHY62KDv6hh/FCNT5RZ+UQqeQ
x/PIjk7s/B8bVZGfIz1YOx/GbtDsTd7ssSbjDR4kiCb2gc3KheR7Gs/Dnp5y1N3h
EcPvCwW+tXAokF/Ffwo9u/DmGOr4bsw7b7I7Zg2pJ0KT0U171rY8yI0etfaOe1mW
ahRVKnZ8dyRwC8GfJfx2eoZ6r2T4rr6vSU5tHdPI+ZaNDpaLFQa5Gdh7AyGlxUVy
GVOwBjF09/Xi+tUG1qc1hyJaizeavJS6uDTdsy4jNVpRl+fkr4Jj17i+c5de0Qwq
CiDpt1N0kXzcfr48Bn0zAL6at7BosxEdESlQZivA6mH1zZJeQn6BCz9YtSMKHFxU
AjE+5DHslQnWC8eXIyF7DtX3ItdsSK5kw7q+sRuXzJN32pCUjdnw7RMQmjW/9y3a
M+A7GYHb4UbaxGp7BunY4oZ+OHr+52hOM4ay3dI/al9u2K2nmRs15ynRgVhhF5Ky
ZuRXfXwKtm2ULYCXbcECDO3hf29SZU3TLfE1zcs5SAsbwJa6+m5fXpi0Z7kl1lxM
/jWzzkHaNRe7M5PUbMPFkaSZb0GcphieNfXHu+xShpshquv8y/pFbXomjlthZrKN
60U2d5wUFCR3mygIGca7MPOTvWjNgYVoFwHjHdjGSULBmObdikOmtPNXRUtNCnPX
xo8nBs4A7iNnJfoVkU7a5OPDiTEkLSIYZy6hLVGydnPzJvbMd7mgzu8HX6dXaOwE
cocGH2Cqogrtr+BvypzOkwsdR98MWu4cGVU3D8wljf/qVc/uI3n6qP8ZBUMFMVHa
NT4EkZ47YJyArsRNWuqwjmkIdBrmXYPKEa015ceva2wVWufegdRtN9WitzKNa9/N
WWu3jMHj6mxBs5vcJ3SrC6FcydJhyKLok5rfmfZELeD4W4NAmZ67d03CnrWHL36r
hZSRRvlPO2o1zSiratC63I6dnBlqcCATWyEwrtM7dtBOKQImdG9jMoi5bpaXWTnH
YOWjBE8dtW2Kzl7lgwySoYCxqGB10ier7JgW4wDPbILWNlwx2C1ipmFHv+jy+heS
5WaTjzmMd11pU2H+J626ya5gy+aGFwfDsjz07nEf+Q7kvTzlZnLLTcvusbBBFxM3
oSal2wnwRTCYUiSbTdh+MKcQXfMFtdOYVSysmSu/CQL9KGWlZBOme1DjkvzY8587
Hy3nmGsQkL9GPwH8Z8MdV4iIVqVO8tvd+RW5Mfbz+L4lfcYr4bUZ4UFXencKodxy
CwK4RSMBt/ckw4YWZo9z0lEjyEVQ09kI+5mdfhSz4ewBK4nxMbXkpXjOAkHX02RP
1/xv8dObh8tmsxWTltGd4pDdkH6bixBjBF2/2C0A+IgWOsc5ninptfdGeorOL2C+
aSuN5KG4i27tI7V6Dktg/TOZWI24u4ZXYHG/PYHBNaqAbU/EzURVj/97LvcidB3W
Pr71/u5w8wPxoB8UICzwmyi5DYcebJBXF8lSWoW3ojlze0MQb3lqZcP637u/xc9r
6BHNW1cY7wzBhQWX/QJ/6jNmeGHBi9tiuCiO25Qb4HOYh/aCBib77TjyxXIj9Iu6
5QaUzzvWkE7QOXHsTVFMafaWxC9uYMyeg66TAn8jhU8fDHFN7H/krJ+euMpCrQiB
sqOiqx6qGBrNEQO8qBsc9gZTMMpF9m3j3p8EREZhAockQUExhXHp2x5UEEuddFzr
WhK4jMqyuqYoBVZAKAXhlkfFvNlFrmcVIL+j0rMrTDSJj2wS1RQ+0fQyAAdU08MZ
AeGzoHYJK1kIxmwV3Lazp1nGe1OzG9OSlXI6rbkRev3vyeafA7a/VmOuLQEsAGaI
OFkJGuJCQP3RQH5L/xvJdoHqJJcuHnq7l0aID1rMC+tw3kOKIvkU5uRHYKrUBwqy
z+Yd2bklzr2J+0iY6C37M1HTjlS1Qn4pERGbI+juZy2vS0Q3Ma2GB6gwhB5uS+2L
Vci45aKJbnXtpXxoynxY7FEdlfuJarrHsbZ/UHy1R5XWFf/9bRxrK63XAzEZ7a6v
dKU7/D7Gq63WpvWceWEjXMOEE6mCWJo75ftp0tyXjos6vsiUFpdYrgZWuGs+PIEp
IyqkAbFHvb+n2X5W4uIFc7MyzOps+M3MWrGAa53LO3m0kmkPjqZAFldnO4PQ59YC
plBHnmy+2laD20DUZZI1s0W224zQZDfdz3/NkRXISL//66e9uhmJx1u7iGrYC6m9
OOn7nGRYNotXKZ/jkoewn6XDW5XI5iHKS7iDmFEe35gHg+YrUm9AzGg303frbEgQ
CBTNohkEgPECVXONtN35CMhkrSFE5k41aVBmITHypDqi8wQ4Wh4NTThJKeMAdI8u
2BkFbdxhjr+C6kZI45LgsgNhhw9cJS8PlQQl6fl1Tia3uJkACftqVXB0pW0u62wz
ZN9wSDMfmJnIUUQSpqOd/i4Re+kdCKS8XjFVtHwDS7aXlg3tXSp/mSgLspLQmkt+
il6zgmaORG3Dh5E2nbe1ifUicJX+9h3dP1kR5UOeV+A/ldO+yeVtsx+HFTtUriar
NLk6WJ206SowUccSmB3BBN74aEfG0HMB/F4CkHumvVNTFqVSWiDVLX/bVEOPTEhv
Lr9YYZZc5UQ49gItpwQAf5C7eWaBFrJn0tymdnrAIw32Fug3GiLAveEgEvmhw/c0
R9VXcXwEyjR14bVs4vj4j9Z1n9MY4Hkt/87WJakAeuN5TLuW6kKtIT08tlK07tiI
8QSc32dSxdBZjLF2c1k3izDyKk5Ce/ZOEgExyMm1pOZFFHOP5251h9c+LoUiPAsT
LKz1hvjeHcU03PYAkS7KO/ZLUdcsc3zopGstZxFJj/pkaiENN/zq5Jlk6ac4JyTu
znmfwmqMGQBR+ilvHiGVM4AKJWrsFLUdwc9ewwXIrVt++2IfsmJTksgt+bPe1EhG
PCKNc23eXOFUUzMOybhQTJ13ouAvXTCqP9aScrMtDrZY80SxLv+Nc4QBMB0vHNiu
QcalqQO4KYI8+DXx9XUx0fgMPq0K4i6hQq3NyDtEc8AS8/BZFl+knsi8p6kgavi4
k1FYduCWX181wnFnlF89X9IC9nQiqP8s2g90fSsX6DXYe/yQioDRRCBfK1vTffkV
eDcEQ37AhW82s3Js1DOo+vceiMNDCpznBRH63SUf29dVEAjJpdFS6e/8ZiK6116d
UsyCQQevdmK14dfpp+2yhLSqdZ5EO+g9nUtouIY2gnVfAtLkWJWS4H0jgrhxFMfk
Hgj6IgR0UNBg4R9CxZ58BT4NymVo/Djj6F5eMsFOAsXgLjgxYcZtkBjl/HrNilzb
+3fXtf+nBCCUWs+x1Cwato1zQp4VHD1kJSAZy0DEcBdCiM2B6JtU4y7VskW1uu/A
hLmKKkuz3u5p5KbpqhgVeujnzr61fmN/7MCz+3oT9Yee3nRMKqv2riWbuHCAPXFo
BzcGtgabZcW+b0PRGOxbXVqyrVVorMQRafBAuKtRhSJ8mac7k74YoSqL2byB2+Wj
Lh/ezNG91yhWWtHl3HySQ+YPLHPBphGYWnht1RehyZ7ltGBvKgeeYnnKitkphUOj
cVYkTwTHL+v05Lo+/Q26luPzmGhNwDqC8gyfypCzpeY9e6Ynjz9ZdZmPvrb2dEBv
Y4BsL2G/j8+O85JGPXSCYI52ulqWYrQK7iETVIcmkUVuZNhY5QelNhV5fuWU8IyN
FMMOYDEgK2lR1uW6gkzWsVAh+JQgpF5QgLsiQzX05nOkL9XL/5dKondLseXy6aX0
Y3TLWbBsNSxwLfAKHmopRGOQyIrZnZz0wbL7ouKvA0cEvm6xvZ6Q7ikjAnzCMq7i
nsDPhVoII7FtvbmMcvTyBLkpxPIDWGDJ3MgkAYtqTIwoEm3GDcdcIeZbbNHQUm1m
KjIF+ioID63BMXPuUtlB24fEESfJwDhV+HI00JzgsWvSn4L75kuy9yWI701RPBfU
Owh3WdmTdeDP3WuVvySE5v/UOMbl3slBU37Xdkrx0JefHZP8vUzMObx+5DNPtZlm
14uBp5tfAe04Fk1w8apIqe3KUozYpwv1Uv3PyLWbqxUQ8nV3YDmqQTJHlVQtKb7E
s+8kPjPX9aB4J5d6Wl3KORb6mnAiJnK++goswgFbg3l49dsD+iKrSA7UR1s3gd0w
KSDoXSk9t9QyfA9fvzQs3n3cG0Y39+c8dYlZtxptHS0R9BET24yoibo5+Z6r8gGj
mzHicNwe//sxlAHI++m0KloYBGPwt1oKabLXzDqCAf7/A3yj2pGH3gM2PwQGZI1E
/Ux4ybvRaBK89UBPvs/yjKFUX8UmJwPfmOwxvpDsND3MF7naac0XdVX9PpInkiDd
skW8zjz59V/QMEOB/VyVMCAJBI1lSM9kNPa0WaV8nHK/6h673PhGcwXHpQPx+rhR
hmmTG9dx3upBmXV7453yBhcOAWb+P/uhOMBL9GoPqMqtaJDE1lDw7rT0+DUMNthq
2QleACMnzBJyxQfNg1qySlPYia6aho6ZodlSjbPO8atozyo9av9T4Q2u2fA7lWKe
7XQL7efkZ/ETsBPP5/j+VjTYiAgU15Aap6ZyMBe16vL+/WK53BUEeCLISbZzquRk
TlnDM42qVg353ll5SuESvy5xzqNKRZK3CVzKsCVYk3Be5GIJBqnKno2BToZsAf8k
ocB848S8VaACYF1FYWiTBu97ktxzIozEeU4sm5WCPWdvA7IGZqms+FkSED0g4flH
y4fjBWN1nahmgjVcFhI0/HtSBwmmAEwUIoh7IAp9y80TDp063BWsc7Sxq9wtKeDN
d0S2eN5adjw+uQ5RO4BGyCuyimp7dNRl8+LsXvRdvk5oby3O+q7fXZgkZ/tOGmBB
/Ld6+5CYj0NEy0TVhiD1fQc3uO361STUQXPbwBfrU+Z3pGowE3tflj4miWSW5IPG
LfYDyI2UNZ+J1JLHMgX84v2vBv5AIXQsjunFYwVnfsiEkL65wWGNXSboifa1uWAs
h9S+V3R70qx2LArglx8Bs0O7SQXBncaH/J+/Kg6NfseH2jy+Fvf40sw92nmGedOA
LV5Ce4N3FvMSG6F/kXRbKHFDJIwobT7a49HU2NN1sBRpy4guathfBTgdhzk2F+xM
vTlBujBvm59xhts4UZ2msMiBY51bOc3eYu1GjGhNgNcRrPEfl/VIEWW1N5Nsk+go
n+kcwc7CV0KAG8s3pxX8U0J2LmetoybzaKOkli7uPbOsekRvlqyYTyWAnWE7SUoE
x7KKVk07sIwa043mTekm7Dt0eux6tFriWomEcHY0ow9czm4XNdoFR6fM8WGEGyT0
t2JoQKRCS4KYjWO/3FD7aXgN37uJZ3DgZM5G3s1AiGaBCPlOocbGk3JtZeHM1JF9
xx5h26w6BxDYtuJBXn45WrE6zHsbSU5R/QCDXWHUVLF8Tul0MsJUjowMNCE5FdvJ
mY1Ju3JTJ05+YFPhNM11fyFonu9hreSpgteoio2ZwiAkTLiu4LpyvHk6mZTDUY0G
SphNYLHM4hGcvnhrLxKMB4mPXaEylkNqr4jqA1nGO4vXGgtpLNyTgx3kuR2uWw2Y
9Idc8jOL/RuTU8oZhi/WyXPI/mf7lxdstCMCYD92KwFnAAo+4o1zXZRdbMx2OvbR
yrV6SBfkm+0lTzpFJ6KHky78eF7XfJuFIGb3UbAPEVMSQI3nx7zGaxgZqzI/lX9G
qrRRkfDKYucAiOETU6QjBQznlOMyiQHiJQPkFkFqG8U/toogS7pAghaQJz/mdwNW
BpKWd4Mw/gWivZRlN2KaY027JX3elxBgnIIgm9E5aoKx91KTjh9K6kbfsIKqvpMN
YNYEwauNW0u95Yml4zU4wVs1dQGtEGi/n9sAKcfJFxOW9EN8RkA/S941rkqykwnr
nmdCMLPA55DWG1gfPM8oHiMJknhwYZiCB0XSQvjnU90NxeLi3vjyahZs/+2uiMrr
wpns6wYg2twOO3Lyxnnd2SYD4r8xAmgzpGUN28036uSkeSeANDhHfCIUs0EHo9rp
Pz0lug00zupmGJjPytausRxYqP9v4qVD/gNYonBLh/FpIVhS949pWSe6fOtoSVs+
uoW5DDLUONw5lpeHSpvnWDIDKIOM2pgzk+pg62raXU0W3i+Cz96NA3XK9RvkQw/4
z2BHWAsLyGQdU7edshk4cCZGn+JCD92mdDV70RLPsHJ+jWzUQrRsuUyWsFTv0fUt
FvG06k5yGD9R2/FFK/E+JVLexjoAps9Yc5PgRp9buhMDdwEPdEe9cxOU66PhDtoE
v5Xp/HgzEtCwq86UT8UVUgDpyvvusWfWWF3UlB5y7o2GV+Sx/sHBcJ8dCiJA/+Yd
hPPphDECs6Cx1t+Sp4G44Bhw9ziKzyjdPusD8aHgXb4MsmUoyOydqe1wntBQ6zDn
tXQJHy7TF4lr5TonuWEm+0xD8HIWc+j8ZTH2elxMX7g7vu83AM0IZj3M2jAEoYSC
pqs0lYHTuDG95f+9IS7DQ+NVmivCucx8FW4VDnoVN3aLw7g7owfiTejxCw9O5Cvj
M4yjtWL6FQbwKDeKOnv0sBnKlowS9/9n9sZeBqdqgxrS3fIdSm/gNyTWSj/HMAZH
HEcMw/b92+/T/HO2zCLtz3IwHPji6+AKGgIxhY4ZSfn6IAzc6K+W9I+XM676IEad
lkBKZl2emxn4pHtHBEG8tvhxmSKnj+K88m5s76eFHIUt6McBrHNj8JeiE+eGU4Ge
dxDV3LLk5V0x14OB5lIGn7gYh4ODhIcwSotnkY4M6CKydoRbJqBTbjRa/1Ruwq0I
ZtvfrY/7qkC6C56x2O4QEsCobG2v4pJx/BRNPjHmEE6APk7eLhmYSe6T0q6yXb3m
YAIJpNiIEvnzz9YAntDa8Ddfdde3gncbRtgqTKQ5JimQxbydhxfPy9UG4wNcSBZp
zqlUUHEiR0AugnpGEXH9WeUPQG6mrwgZFEHf2gvYtzS2I+ymvwcrR7C7qe/o5s3G
sk1AW7bCHs9cd/fvi7c8WORJKmV8BBrS0ZWuuqd7tVrgRIbfqlz9ihLEc1whntzm
yMPPbOzB963DSVjJjTGHWV+6aJgb93Jt3krbMrCZkLKXMwi6+q+P2CgtHKGuU2NY
ya0IopdRncvxvYOhso1+a6Xujar6yvNvmoyUgJky07UhIRI66C2rP/uC4xR51GrK
S0cPafNhOh+Tzt0uvfzKI2RUkWsntOkBc+eipV81yCVWRruf8iesh6u66pd4FAUs
eFaxqv+yYxmGk/sOgGVn88FmE6A5RoCVKxpNZYMb0aryVm6ruJbbwN9sh2jh+0KN
aQOCAEEmsV8vWaY3xOPi6+o3L/rJi0YPMUB/NNCGJTKUUr+WDb4W8omHFMadQxyC
mnoRB1lSRkhpdo4iCyJ7bTZxOmmFKsdhTE+QpyZAiv8SLCodyalT7MzcBogTWXff
1ob7WpXYg2ttyIDsbI7c25VAeFe9b3vdtZ+s9jSbvBw/0MfLrGT/fzGX4ySO0jTM
9zaowVu2ZgBQhCAuGd+W3yhuBU7aYODhnKsfXW9i5N2wdMi24GUSyOOM4CbaqZAN
R5T1LRvNT/awkXDtJYKL6bO5aQkPk0jryYXvuq8+9xcOmwux6LERmT7Pq9ZmhX+Z
zUT8+RdycpHy2zsuwr+bD/bq92urlSpJBUldD7VPmVqJ081EGG9BYg+gFZYuv2yZ
j9QeNJxlJtFReuOl/EAoTAozzTSNJqACLMUIqUj+Y3jz0d9CkWhZbSlmKgOssmBA
apIXWdK2AxwsMp5JkQA13tloYrg/1DOtcN7ekttxImv1Dg6jrgIfNSDi7sssf0/w
Rudf7gqCQtQJPxiddOANG4nZhSUQFfV030cjI4vTmp5Ag/NeSJ9uNQhnWRDz2W4K
M0y08dfs10GPAT//7eR43wdBREuyPXhfBhqDGYcybrdqsDLwvxk8RnTEpnr/EvUB
N5jC2h+VjXMBEcTCZuewco4T5xcSyOri6C39dVrb42SIlLDGOxUJEOujYToM418z
uow09CNKoeQQ8Uep9qqn4Rq5Vv10YMxWtCIfEBgeOIOBsCmJqbOApNYcnTzUP8Iu
bP3h7cbty1hoitLpiSxJzxZnE1EVK84apdb0RkTw77mFaKk4wWkTjzOB6C6cAlHX
EyOeaeNQGcigwIJSUIYmHaBQwyRsui6oH1DMji4oKg+Bf8+hhYQByvWE2J4CktOd
RoTfxlW/uDzw4Yg0d1D5rpCAZ9VJJujX8FcaT7Wd6jqsJualsGdU4eutxYqsyzJN
fl15smc8Mc/0MxJUMj0qY6jDYnHugULaX29aAKDEy3RFG3lVSBWkrtOrP//MUfD+
D+gP1Pq215Ljl6kk2S5mZzSZ6HYUI1by9YWuElr1rPMEozcK03TCWbW9GVr3RLcP
7GZXMV5VL/Y4jEgK36zcFUlQsXusSTd7f1vGSSfi+8h+1rtVa4FENm/iM6/ERwsn
URPvMOsruDtLgjwBtMTerpEfjkA2ZN0w45pC95UJWYT8gDc6ZjtS2TdjiV+iHATL
ESNMfcS9Om8/z4/duHut46/ZM5xf+2OQahXEtdpsUhH1PiSSaXiiZSmavCPbPhqK
1fUaPHQ/WT+isHB3uG2dNmd0pbBUMK3RGOfvXBgo44oWgF+kDXpCPIWWzGVqSuBB
83rewEiFGZZuLg7onuv8iFRg0zWHytfWVt9bLssnyna5pcC5b+GrE6vtgB2dyeax
CKGlrLLnW4e1MGG3louDP1rk50ZG8AP/wobbxa+JZ7ZENI+2kUDZ36HGNRoxgfRc
Zbw+pmy9H6emahdQcT7hGDrhYmNK8UBbST09pme3GISG5PGi5k9KykOIbYJuw+/g
VJ8N5gbeH67RvBQSl1s31r+XzpcYAb6Zpwyye115czEzmCYV5vpRbkUupDv2wg69
JelPekKg/u4SYNeHFnpaIaVYDFer5bXtPjHcG1Q51gyaEJtkV6Tj0U7n7Ewpwffl
nawvNV6xtmC0ftxpbXB1WtDPsdQOSxL1u609ai/71nCvGDwmRNtnMTQiHXBzrrcL
dGcVAkYV2sbMsQTGSS3LCo5Msb03EPnOIzGiBwr/sRbppnAzCAObadW50BjM9pgJ
yuBLiUBUiJPZ3MI1+eeOMxyZo+8ydXaD7U8mfl6G9vBlkZkxS0o0jD2A7ESl14nS
j/As7ZKIlgRQ40fA+1Cr2pDC4QgebKnSVlbdRephCMjKAnsURkm2z41X1eyvZ0uC
0BXju/HFLJF5vb52Dih1LAodQEXJ9U3Yw/LV47xgY75iLNM6GeAUkuSOpiPiy+GU
Xsr3hmjYuHn3j9TSlc53OL7AZ1d4G11inbOR4n/m/WSgbxKJzC5FHAupKNPF9t7e
mDC4DC6IYiuXr+Ch02OwSr3AiwsAs/3fT4uRDooSFQoT35kOmQutSxbUOIZTkZwR
uZDc20yJECgHo35MRhP+/2Qd5mF0WWQwtrjxzAF0ECJGwMJ5ImIYaj5qTR4fa9ih
SKf+2RPErHawdXTEJ/jsYaZXhFz67lFs3QL+/zrLCsOGWhqYBCTPmFEtNFN7jQFF
TtlPMA2ASxIBtn3ArZSZSOKKsQXtdt1ECIjKX5Q5h807yz8slOEH6ekX5LRT8c71
w3ERhrQbQAxCBgDWN9YMWTOG8kGvvRMQhn5jtkEtwLNJZlOUFy5ZlUgA59Gy67OF
GHd7TX0L5GgHWhPqzePXRxEOgIAm/BRBPz/AW8UnTt0/2GZCbD9YeZaRkD3rBW0D
7tdPIo0MBtCQgmreVhgTihpplHBBXSDw0vHYR/FLwPJ4S37QCmDUMR1QW5A6s5AX
OfVcm8heXjMwoCbTKcm22dtcKyKF6dPTNHlHGGO1UpjBoBluBjizEjOhkgHz5eXN
BfCSS4cckpNVSy6iyjrBM5zCqOwoBzPdTOYgbF4wDHQ+oC+g4M/TD+rPDPhMZFhJ
rxKmh0ufnXiA/6ASHz6hkvKqToU5QCFw8BENCrSbSUwDsJ8POh4ivXbufdMJmjRk
KbwpPLgq5YIjgn2X3fCdJIDxl8CrsocHvGdYDKmrUXa9tLYmH6rU0Gu520uxFKPe
qnobqSg/RRppGg36Swjp3119eqjEAVp7Nj4oagjQAOK/nBHqGkkhD0wEKobdHaBd
FyMWE0e232vEdrvVRWz+FLbWg/ldQJab8xqp4LQ3kiXCYdiLugGjU5Ov+gF9rvs2
NolBf2KJZFBCcNY7OPBvZeNqcIG4q8NiXr07Cq5cDvzUjr/uKYEw26+26sUNogeF
VLd9/TM/GQ2KypgZNvfwvRokEFwy9STzLXOE2GMcdqhTEuVos83prN31kgVzdG3Q
cv0NJ5xG6rQyzgAsX9ryNA1FKHCBhPQQXHjFuIBlw7s3ZR4EVcfV6r5vcI9l3aPC
guLUk0FEcOWunJHMBlPJdjijs5FTZj5FiuM0aHuUiAjUVBvivU5SBXyiY7agzLUi
BQ3wXktNTVmBfzKBja0+VzOb8xCkRDPEuPIJndZhzTf3kCahP+o1cjlEG5W0OQdR
pSLXL9oOvjcepOWBft4cHALz6hbMdAdpe8q0fSu8GVdlAuE4JoI96WJhDG20TPv8
tIra/BTkcz7pQvUnhjnjLdqBVx0ZFistpA6PmnDiCvQtHYP9urV5xQwlXb7oEkaT
KC6vf5aGDHeXi7j0qwgcVadS1rAJw7bb4gAXpVZX7OvULSOJ4oIAEhsyB/Vz2P7F
/rplC8wHIXOgfZA3B7iYyMVuHiogDl8Y3Rd2q6YCH+qiN5JbhAT76XFNEj2V3A8m
rGVHSvgKg/ctYR/syJnieMX6uYGUOOQDo9Oz0dS5MskCHJ/SukbUr1TJS4zerTbV
ck6tpr0TZgeyqD4bV2D5wW8OcgyuA5RwoHtj3MSjz3x8o6VOqTmcj9G8gZjfuYTE
+J0TxmDzQkbw072D05Gcr00hSbFPn8cZzyoDbDRBP0HEsgOFdaNrNNEh4eamXkbB
oY5/J+QK3lUdPtjByXVUQIlp8oqzp8wDCYcxo2x6mQImwf7U8r3qpnZ+9pl8gHPK
1Ua99lvAKYJdygniztLPP6jIxxJqyqC0X3pp2ESWOLoJgWtdjO+SU/JPiv5HE1QJ
nlNJeKfGdnEj8oIBbcNpqhrmFYOn7MVT57V5+d54QfICLhu5ObW3sN0v7D5nMl1s
tD6UJR2BK6x7UJfk3KYgYV96GRZNc030/Vd4wuHhAo72IR9kXTiUZRg1A7dUBeP5
EfFpS74nj2iAb5+VASSJzSfEfBqYqAFqK3S9XtydepxRABoWkfaZgY+u3a2dLWbX
W2Ia5qkSEqlrZ4nxSNj/X+mOcwOiypigf+tEmb3A+CV1HutmRsjgAgeX4DXNTvZR
7YRUaqqAUeLwTlZNmHCdZKz0C6XKe30RkDv9BJDbB28sfSMlcVYckwtzQbdveK3V
3Hp5TZP8nMLGmTn/cS+l/kkzRxPBIKtIQAZBHEzNtOhGZUoBITgdgAfDU4OB43rS
0O/zreE+4vqnu99hDLVMB2XwNNlCY4rjHXCWf2W4ljaPON6JEIl/JWm4mXUpkvAf
Bi2tTjnrEbeCBzMn+U0UIuvqMxZhLu7Km4/tMLgMhiOrBXjlXGPysKldNv8MrSI7
Kore4pN5eJDHBcNcdOEZP3feNIP11R+5IV5wr79LirY0g95Qd7ITAmdqGlawftki
VLnzC++TKx6yRnGGB3N2raa3Gm4olNjineET4EZ0QF/6892J1gOYkZNvc0rhJobZ
KAVarNorDXhYBwymx3WtoM5R5uh7JX7l/8vu1bSdYw34gW8R/apWJPNiAe325WL+
xFQsv3z2bX+to0Av1HE8Puy8uC0upzboqwkpNPGBsq0oAqCTCBeGONse0OIb1P2l
iRmwy5LxQA04iHNPTZEU3I2RrXbt2RQczuZZORrNqV4+kcEGcBPUs5rjeVZ+E18a
dpYg4x16BalLZKK6xVeyiUoWtEyaywhPgQOD7s5ei+BEbqeNPPb+j1w0Rdtwrbt7
NC37eY1BJ0R2hTZlVkXFl2Jw9OdLg0On327MxiFQF79TmHgqHFasph0OcMDSIkUN
Ltm6/noqr3Y/qLGGUB9WCX34/6F45YexpaCqY0nNqGwRdsZkbE38icQc0CGRQKq8
0t23T34ucTcKSk4vsG2/YtZWyjx4t/50TOlfLB1grEne0ZcxlS5ceK4F3VneJo1r
t+d6bSYuVuOTMf8BO9Z3nJ3V2fC6Tam/9NHZU6mgmH/vWHSFD0uVWgNmHaMOq/Nr
4GWMBDTMhg3Wh0CDoQ3YI0i6lr41f66XQ3rxaVUl3kCWPyliZErkZjj8AveDZ0ru
mD9eMLPwI+WAYqwSDoN1YRuthOislBhz76mNBtIwxLgRMmkwYGAQEhTVK2smlMLm
DyR29yWHI+kfrX+ydTy8SqcA1km7wqdgDfCx3ckqkl/hcvmeTaCRrzFaJ0TaTwPQ
dtcTKtdx7ZjUpY12w7vmEpuEFyWACF5IpWlN/YYsSuuoijf/jk1XdJex+/yPkPCf
bCMk+hhBAe0pxpIQbJ9SNlPRHLWLl3d68S7kc0Th5Tz6oNuMUKova1kp5NpdHGtU
ViHHvPL4mXEpnfjqY3/JYdZE3IIVeaHIwfFS2HefUITjQ7Ry06cfXSPD5iruBZXR
lidvmFPQ6NRZqXiTkyp/83Y4ZlYdB2hfPVHXBxE4FWzMt7+WQJKDL1vNA41B4kh7
ZGr6/ts8BQ1jN9dvLosW0Nx1bWQRq32swT58ZhkrR+TheGZpj7EQxu37kJ1AuNvs
KC8vMYNT7N7mSj+L4QUOcdBuDUz7xZdAiBRy53Swiacs+4MVl1yDwR5a7/cEigzn
UTbPhrxSRo7HvdF1/8xfNuJJL7V4mAcv/q34Q8XB3d3AIYMAnrCMW644rZQImO7c
tshz7WmJ6YUXvzZ/npdpPp84kUW0wSQ4NB56E1T54D0MnQ6O//q7/b7fmghh0CJh
u8AnQY3CLS5BztuqOMpRLd/Qz+rKLSbsFGL6mWxQPIYe+KTtzf5MhtEFoigPN0JJ
rY8otXbIUkH4j7u4DVYrdVm1vqSI3zwMpp0DXFpf4CMPE9FZZstjA5g6YpM7/cPm
tb9gRmCn43JwhZ8EW3veQwPDwh4Ur4WsiRtOhXGMMbWfclrIb7mvyvzsL0cP8QYe
7tGEc5hpfPyNjJt8AQUTHub96gQrCa4jB6hrP+SshV81067MsgUlQVeBlubAkZhL
vPIjipapPxI/9xrsxk6ss1s+2aJZn/PSM5hXlo8/krs5DgnZmAREx7o3Py1kVolj
0HwzmsRhnWYuPSsvclQ/j6toXozqmN23fw/XPCX6L+eZJMSTKWTv0D9zzGNSpfNr
qGS2NBR2uN8JCp6IHXK90yxyHLlRto08c6VPGrDnT2uQPYAY0kBmcVs6aXunInqF
C5i6JhkeT8OUaU8zPO6ZArkILLLqtk91bIg7E68eAd8vLFieCZaPS6YbFPoUTMjA
iclhdn9ktR4HIt5/i8sZWwy4IqQy+zGhYMt7Bf3L6p674CDYWg2ZGE8CQ8aSVUX7
cPFA0Ony/bsTnWxwDqJPya3WLvLsP1II7vJvr4d+aLkAD1vdg2Z5UiIDOMKZv1TL
8VSDPMkRY+TqnEf1FqiGUPQ7mDKhlfX/xPdo0EyhccJaSHDj64gS2UHa0CbuO5S2
A79YWsGg0E66+AJdcC1MG4mAr+5z/2Uuh2B1oqVSnvmrrMjtF1i/HfeXc3M4k7lv
I9bEXzUCxN3KDQFA4F7hc7tdJk+t75Iv8Z5i8ZPyoTfWOwdTzJeSH5SJnGplYsjk
+SD2+0kklVZAjG0kcUnam/ylPy6zkBs0FNEoea/StukhH97pXYQ7YG52aoecmUIo
UDsPKFEpJKsUWbpSkuUaN402r06Sm8PSyzBCrfQHs5Pn0iqQ7cgcC8CC0XA8P1pC
lzPnRjA2FrM6hsTcfZi/lKh1qhSUfes7iCYPyvhrijVqBfdB1Ma6AZVTivTOzsqA
SPQyGfloEmflfVSQa3FAU3nDXSSU7J2VtWumErRIoSjGLP+vKCWaRJXtO8bv/Aho
HAFFCSzZ+8SEMagyNBD/4Q+W/9QZOzSgAdlwFTioUr7KEzF7DbNJXTzOPahzpezq
nSeLB1eXgvCMv+4+ho9F+m7dKr6az7LPGg2nzgvKh3H5K+M/iklQ7+JFAQr2XKtv
ww3n/9g8Xx3/5Ib0vArQW6bw/JLxclanurNF+O43jL8pm3VsgwQu3vh4KqMmllEl
4rMfM0daDchM/F34d5iSDdyANkVn0lW1QLxiIuREFfuUoFznEx3fzmSmz/a+dt8s
bb/sL05pSHAwn9IGJM1PMSp8akK3kywJV3TWXixkBRh0HWHh+22NyKK3M4VVDHL9
9EC3I1QSogIK2Z5Nu/cHVlP7ERt8d4CfK43v3otKoBQQziVIIarkMdVgM8OaQ0Z2
vlb9c+HYAES6Nxd1ggU8T/Tv46ng66O4ZReFvxEYznZJ9zQBaIm1eEmVBfNGEilw
SRfS5UplOE9e/9pjOqAGxZ2dvIHIqBLkp0/oF9bCibcGcOqW+B0cxdq3yrD8ws9l
q+Ej47xGZSwLZBJcd3I+INA/P+AzTEe7EdmA9fLxUJqxLpBQA/nkYhoqlfRiRCgD
EquMYJ3wY9D3iOy4GO4SQCFifZGYys2C3JA7I2bVJCLg6nNnTzQok0Yt5SPKdSgp
pGZlEJF7fTyYH6ze1FnzmFf34P8X87gPQ4YB/tMp/VcgNKuTRdi8xcerSNqPO8+p
utd1i5rd+0Ercd8NmtNt6OORHyqhuGohheLJpcG9Tpeep38W/Q3RdULQMCY4duNO
SZHmjpIOKW6CjkfH1GKP2PrjnJtHZdryRBHBowx0HOqWvgvPCFoo7icFR4hjZo4x
HwXoXtif3jeLjwZCOHn8KxMGTBiVkbe3GP0W3VZyYp9UvyNb/HNwYfZJcuHYE1Cj
iWECkxfHmoFatsCANrvDIqUWV5rpWuTBO1P3qYLj5PTbZwwZFVXNVBXhOvWQs840
0dzg75GH2BgDhdLVigh/BwECGwXYXn3Q7c87oDX9ifm46GcJvxZixWfA+p4NgT9R
Y/MTsnTwrtwZcFWM9aZKzuxuB3h3DMz1K72gU8a+IDhOSXaQWGsPO8cCrhM8uyeg
j8jaB621U80lqfespdsgg12VlPZMS+YOGljk6ScUbI6xgpLnEoKNqGGB3S4ol0Te
uKpRSP4Pi3EXPnausSVl+SFOKzLWdN7XfTopNPy9xnzrpSDBjgqBKXiOM5YRqr6h
c6BW9kQcipl9rA4k5xAKqkTZR0Mr4dF7dFkIV7za5W/zKqYaedpB8F3N49IOya+d
t8CXGP2dX08flgAl8e9Xo3bXqQcpkcN7//UlxfbwbNo8BfoN44osJ5zGvw5bumKa
IL5XdwLWQkyx/2kYsvpgxm5F+2YJxLg82/5wAwhNU2KsTdEh7Gecbc4Wu2heeX5m
oE80fdRggYJ8uZxPniOBTjU4PTJPwiyRhzRHQru9yQzNjr1N2RoJpoCp4iuLXPzt
TeQOKhzUCOCJFfqW2R19b3g8+ITsr39OiY1hewPW2PM7PK3RpV+nWlLf3y5mHYhq
to11tCjWjMITuf6gLIzpFgBIq+MnL80YyvW+v2IdDul8mnEBxTcV6j3l7yGr9E25
1slF06Gza7G3I+T2bPnvEzLOJDc//aKT7KROKrnT8bo2whiNCUOVOHnix9vO2ZCF
YqHLemEe/6C5lmexa37oLvoWsA7Lyk+Jp+cv0AiI+DbHuXbhQJDkzh+PTPxOe/ed
ygQdXytmt2yylatHPlFWeyRwvpmwaq1jQlVLedYpxhMAyMwDZCHXf4sdqcg/50YN
7LM1eqvLkCCGoGmduzC5RWV9pzosLIIt2A7fmR2HoaUPpvmQg/fERt0T7wDBBmSm
4jkJcm2/VmQIJKh0vQGyFzXAZkT8Gl4MhHqjiTs3KOPQTClAXCBfQuNAYwmnb1ib
XtOIG188A0blRCVMepQE6l56b1uiaQx+8PGi+fHDoBxudx7k6a5/+nsWMfCLmBMp
q5e9iU2hUhzJjo0OV4QkkJgofobzz7DcUkLKRH81lNTG24o5117tVEHsKfOaWDbI
3n2eobgE1l7OLHU4ZVt7efIEnCtoPPN3gQXGA9Cz6tMMarHZAFH9ZCPYnmtz3A/a
tgimkuRMWTrvA88BK0+WPoSxL5O7sn0FfKv+pN/eL4TVOAtD9PGXXDowQ713rX7m
t5vlL2a1jCY4u3jVdmLaX1q2kDOD3cvgOgr4PPgvH2Ual+7Kszz5mXErcQzp2Jza
YdBtp39LE2msSR/Re9DrhgLOMkM0FfvxXtW4Ld/5WFFgxmrQjB3RVaLpr3NkNSDm
R7p3+kQMJVVHRM/Kxk5SfN6oI2Gw6jXY86gMojejj9kLbapnmkboDTF5+E5LV9vS
M/KuV4IjH5UApHwGXaeA3Ysa8HpPmmImXc1S0RUcvHCmT5WXut35tLLXApcmD5pI
z125EzbYLa6glAIBr0Qj2q4A3q1wIanFwPu4AhdRSFU2AcY1o/REcXEu7Rl2nE/u
gwsCJPtQsKCTPrQelGwxICWpAhsJ8s2faKDx/CE6CekZZoq5lpxs2k0w2DGvsZCt
n6lbPxmxKpL7a67g5RnOjU7RvgoC4sfq7V2/j5thDNSjMzo4DfOIoHoB6h0j8opV
JiIl9IMEcOiDSeXeArabfRrxfJ1YBUcU/zhCNE1zSbpE+0RNaesJw6V+0sdAQ+qH
oNHPTmjeh6rmyR9rCoXcZv2jHEF3kMdyGLMuR/kJ4gaP3M1EOnuaoSDfprGQ2SFw
VjGyWm3iS+PgpdZWCrf7LBm1tOjYmIVz7MdzS8A5ukBCXx8fXui3DU9KQ4rhAbo9
w7QEqr4EiNrA9ZCoHF61WjWo0GS8ZFbOaWzXjn2DUS+K0cbGGiNa+MtlGxliCZWe
773Chkzb1CsAD/OU5Sz33qhzszBvmqZUoSnwUpU5c9H8CF9WjXxisWTeUHy4UTXS
MXitGzau6dMq6rnhFAWlTia/lr4y93FaP3PQaTMQ73kBmN+WM0rMuZ6Oi7O9C0qP
ycEE22/CyoCDLro9e8IBW9xm1V/ElSIyv+QBZLjzSQFJe/4mQTVC7/f6ZOQqc9yZ
iimXU5agDUzsOyEL+AeNefbzLbsf/Gq8iErhstJGFJzZdeGRzl72Ps1pNRng6Nn+
rMSQVbvncVJ9dTPcVhyO0xjQIB3xOVvqojaDs6AwIssLO6XFrSbtNgQ9NZ177QQC
IQobe1FMDR1AgLG7IQPcGxvv0jYJuwmQBg37F48gQlg3NsZg5h2c3SGPVbqKg+Eu
UdXN6kofQb1o6h5rBOYKdoImfYiw8URSCq4Z72UfztN1lIAcUDfvZLpi57LIdcbI
NW+PjNMMwFDhJ7WGV5LVOX3UXY+otPSyOMPVdu2F5ticSPghu5mPa7N6yHNYy0aN
DKK4Z58MeJHPiDJjRE9xvtQPzRg7O0q7cbri0y0VJguVWI2Ea/LxjsmJbccpYuye
e5zDDhduo7LEdttyUTVOKSx8eLzX0ass1Gyqu13WoUf4NEGajqIEzdSNTL3+xsG6
T5p0zx+ZzEMyx+3KesrpLTLVCKWjKFfYcVMtPiY1vL/j1bqmKIDm7En05JOS3ocl
Uj6oDJ+cW0WzVUv4eTmkXKO+jwCueb9fIt9jmujxALm0S60C+Vskb/gz1zaIBBzM
pAd5itRhGHpsASoJGT3UsaFacNsnqZ2iuYiHp0Te6NlQGe+lsc3nvMtIYYVP2u0I
wcHURSYqfhg8zUZT90B1NnjuHW0OXscMWm5BXISIIdF1D9+YKlEbBCuVskVqZInv
Z/UyNMsQniM93ykvMd1Qa+9U4EqUuEf6DVhEFvP3We9TGMfiazPOHXt7XyW/Lxoy
x8A/7KX30RKngEXXncbU9EnKUHbDUQuBBtxCRYtpyKqn6PHyggeI4fN2He/Lz4mF
sRrCpE3UpTDziXIHNKnl1GF3O6UjNjOUVeAv5L/8d7ZKH/O/zqauKXZ4Ksdb4ifv
m1pBofPHTj1UFonGdjN0N1XReQv0joaAlkWF4YDwCvQkcYO7z2yoeRHouqaIw0DO
N7i6pX+8YHLg0gC/JGj4e7zp4utTXuS89XkZi9F4DUK+cSkrCoqxuR03KCftTs0j
n0wUgtKK1fEW4Wjh5nr16g0+/0d76nVXNYvd9CStSupgRL7l65EtPHltLH9jCIur
MM88z802RUlK8744+gnrv4KmHlDg43aBgmWQDBbIa7utKyN+Xkw28Hs7t4OA0bF2
OBQrZiytb8c3H9uujyEkYpQpHyOAgEQZTRJtocgeiU8OfuVE7p1CqKMYzjC1YSfz
l3HN6nzJ1nR2aGEQCXsK1dT0hEg0hZFXKkPoPs3UgZxtQMi0MVuoJCTUmg7uXOxo
vohjAxueKRQ3/cZJ4algLkOSYZjLieqZfaXb9v0GrP5NJBvXJieJot4ssyT6R+tF
hOLWK0fJCP7TYScAIKK9TQi439rge0YqiEm59FB8S34WuT5P+Hqoe5Frx9iATAxV
Esmev4sNkDNXVEjy8fVrQfTU9GxNjlQJf1d8W8/ptD9pfrYeIjR6iZbUK8aw6aOl
eAIiW1/DqXgesS3/iv+6qg3gm+JSELgNvNm4qyweKqsVPaft3oyvyvd04pBdK4IH
p818Bq2iZmYjQxK2p0viil+95f5ToJ4dN0TW3wT8d+uDagepffDh/rfvY1FMC0nU
UCcHJ7JcoPqqPkI55QyAhFllI6mnlUzXamt7VIZ1HOWizrYZbhyU7uI4qqSXJewo
6skNaPe3O8YsGP8odfDe1f+RG6CWavYkaGtPyKjDSjsr2b93mFPUOCRV7xuami+1
g4Wri1LjqYJJh6wuE6un+m2IWBuFUHGaqpkUo/lLtPpqbVGN2tTvGc9pCYGH5IEs
THdJj8kUArgdKaY5KTOfGZ/cuKc1hd4dYEx54YWrYyFmejGX27RF7eF+oVuu17dI
WCOQAD59QJvLq/bAiGjNLmviJ5RrUsJ0aCpB4Jhni3wlK24CsJe6lAA56n+NZSfV
ZE+Y1qlc5Q2A2EJ8LrAs6wzHGKxxYJ1GMgyPtLpNqtFR+NiVilxfCzt24u4F/LPe
Jme2CHKiETtfzbDl4hjbziEJ1prdG3NnP4jBdHr8YlcpE97gwGaaUx+1w96Hfgvl
AsTuA0ai+yekF4dVFEX24XMlc1d7SNSGQ3Kimk8e1T/iiF2FX8djmGCkCfsAkiEd
aFnkG1COf98hu+wOuKd9LIUCb7r0GgAaRmbECvXUZLDsB0GthQio1E1O1LW+mX8i
VuLKIwP/s61T+i7iAYBDhQ03P6vDWIYcoWT1cNfX3U5yu9HLnh4t4pz4p96AgfvH
kXtk/GgQfgeOjXfo1ywcF3yiV2P08eu/lkn9zzv3/PHUiJZp1QeQs/radoEC+uEj
fei1NbhNzSB13w4kCdl/wgQ3z8LCVrefVgGOyr5AdGI4ClbtkzPcbx8uAEN3/k6a
FPkVwM4/SEB5ZCsEGNlA7P8AEaoPqHzgCBmSNM73tJqWKPfKUqg7oh37k/u2NMTp
ENWf3h7bempCVA8FLg+jTG/8dQIEeT2NPvLxukeHNdUN5U8GaUYTxBM/6cbAG2Ta
S5jTruc+K3lfOTzzKLXEU1lxHImNwMx2GQC7rb8GbbZrYqsCBjsopNybTadu3+xU
0rA44UEklkcCvn1zEshDz2tKYu9vYcNr6wdPXok1FbIx/IwiALt2Hjzm/66iCENX
p5CSnOadkIRPAsVPSk5AdsdIXBdGKz6nSLdEW9gRE4uMAhSmptErhKvRh+Hu2EeL
VyyKacgbgDLPTzmuAMQ5CyBjoncr7VVwEVWrntlLfp1SA2+KUxYROnh7urEguYDC
B87z5AUewVABnC4U2fmY/CnMMHLxJlj/wkvzoz8Te3gOdH/GMLlVMYzMeEDe6E1R
xaNd3yPFEeitz3SU3WJBSEbho4Ryn/NPoPb2+UDMG5mKdyKYLX2+WZhTxAWzFOGC
SQw6OZYeq5aH5BKOX2bSw6qePbMWHJJbdFAltqfiGTZ8uP42iyyEK4OfsRuzmbjo
Ggxees+RGacU47i1cLb/9xBx1LaWFXreEdjIXNFv2Sdt+KRORZ+xQsJEzi6A5v6Y
b8+X+5qnEt0AqL4SSeDH9umXmhRedtPd64E1+cdfMBmEjOrrjxlND3eKwwVJ6dwg
//gT6u5z+64gtdtfU+kQs/87z2hgTzY2NydBBshtbHWuAR73rjDFWN0jmXU0UCP8
GkXTXjlWcNcj2RNTVZs/n/5mDkiRwwGYipLtldpZ07rGDY2TulCM4efHiIdSFwLN
qh1E2t+lyqPxctf/1DNBGXmrrRzIin/WjBEGQ9JhM36kqS78o2LLvJB5mQEaRXtq
w0LDMwq6jcqolMJuPMwwuu7EOte9LuAJMYy9uKo3cnW61YqHwbcBLW0aUvrOn1Cm
4vQS75AZ4z8yM+wnLHI4Yt1qEFTGFlMP9m9J2zFhu9Hp4RQKrK+lU4qsDNcekLb+
tkn+o7tLzKmzqowG2Bq1Qp4yJlWRJZl8l3k0VDu9DfWJl2ZpOYVr/Tw4xgXjlTGN
tuDn8PKNl1zRP0kzZX+gOp7/bGWhUhG7M9SNGPI1qI/AobZs/8gAoNQJGboaVqUg
55Q5DX1EkpmAuYvm6OEVWLkZmynanQKVzHqcsiWgIMj6E6aBMD/RFhVtMQok4Tn4
n7mZT0vmONaH+sFNi6XBCULEZv1iLb2MU5Y3HIsRGXAMcGTHMBY+yO6VdoCC7roQ
LM0YQ6E5mDPErOISBeG8p52KhmIfHOT9Dr5D2HW6uVcS9AFuOY8HAuQXsiu/ps1G
2PNOb3CjcmuowZlY73dcjKDEVTcFS4cFIeCbT74fHeEYC589s7dD0EyPLB7MIMR6
d1KqZvRjVT8Jj20TukrWU/KoV0Lio9EmwjF0YGU+5kfzfKxoea9Fq3iCVncaPstp
l0bbzhvkAOsQNDv/D1vRKVyZyjlOX/GojnCRGKbYySP959iIfuqtcG6Fba81+0Yh
XYa1eVwtJ3Adsnox0C9Leree5pwVOjlOCQ6FQJzsFLpb8nG/NWeJGM0XgOjw2epu
inp1xrghW4Tg72cPlOPzZK5vl/4lEZa/6QzW0x19Pm+I97uOiL+Csaxo5gRV9eGI
Nu2fTb2wJOJa/y/E/JYZFBJgUtJecxbpOmXv6jKqtw47tT3OLGDri/LpA9e4Dlmf
iruUBI12itp6mdCamdmKI/YZFGb35gRB0jzxfEPl5u+ElfU0CVa9mpzXrxxLxzah
yTsUxGqYDIgh6sipEPG8aaRaJxJIdz9Z7NzMaA8BNfx+RPPcd421BADo7ayZDd+P
aDZ8xCAx2PW8e5QY5uq0t883sFayDs7O20RiYbuLA7pPvjjjPPTCWEmh99j2yHNS
OfTT6NbV+Xa2zD5sPytxHOTktDFmpcacF79hmSi29SQXEisaTkFhPSDbSg4sWden
7EDX7qCdTJNMVTHymIZmxeyWvBRbKjDyHKT+N2rhN1T23xexPB/pvJES1INqRa2k
A4shMjJUzOP3WDn2g+WNEOpbEbuBO5AIw+zcwSMgyqyyXdYTsEmII3dgv4uj9q4J
/aekk23ZBuAxDYXCrFrjPKauanzCdqJTyU0tcNAzZY+WVo7ixeTM5YadjQOm+Vww
QZIkC8xKKB0vAgmc6FS4XaHPjSPEDoSSY3K0vRKq6bq5p/UQzNzOdBIUHurwp+yQ
gFGxjZ1BfX9Mw/rKSkkLrkHwZdr8tQUVYMRt/HST4qto/xNEEWa+8UtFFo9tW+9E
mNxuAUijKQ2kYXog/ylUOTq6nokPW4RH8pE8W3N1dkUaGqd5K0+wNmpb4JcMIkxQ
VCJ3vkW+A1+5lUZPzuHc+6jMEWbp5zYDUCOffZzOwod4e4lPXr5+NhxB7XIG/1A4
ZLTwdMtojJbbGeXNUqF28XV2LWOHuAtXMTfVxm+gxIgb9W92eg14AUetgBS/6yjt
quJsFyL0n9BJnKt691hkhIw3I4E7Og1b7Qlj8Vk4aDBdmZw4KVxJ7G1iKNWT8x6d
VgvHUTtyHaIpUoVpoF68IR0+/oEBvlnijB3DdvUegzaTSL8YRT8Yj8q9421i+0WF
hyca+OJ+nRJSRtHqiDWHHoWmdz5ImJX4T+vZHgTyglpe+mYLwWPDcsNogPlca6Z7
lnIG3k3Hlwy7O10QL5k6gs/AJnj9xHvh5HaSLRw144tUGyuJvwlef19EyrGu26b1
tyb1RccDGzd35ycp2mfvwHJ9XXjSNGkppfJwi3lwX+XfZqD6yyvqBQ56vRfIrxVF
unV9bU6qLgYReoUury4055Nhej8VBkUGd91t7C5qm+gYsV31TfvPZD/He24mEWQE
p9utByJir8IKKFd76sYwMDSJodSKt3OswpHDcqOJ6igU+OCDn+OUBWqPlbJ/KGUz
eQP6gEWOkg2MxB6YbuEnkQgSzW+6+c78/uSPkOYDHZGCkEUG85wPO0eUTXITyV/Z
L4cv+qxJbyq4gTJYTGxH6O3S8cS/jUxZkObaDmsI9VyxIPhDAG1WFtKmG/Qi/+kb
BbAnA5On+wz6zxtqHo6DK1Luki+ZjSG4c9SmG+0nCXy37c/xw/kMdJ2OWD7+tHKC
H1KBB+7+esEN0+Gs66mMcnQSiHN1XvMZi25AsdCaf1B/0hc+QiMFyWbn2uDoFqn3
ZZEIAhHduuyZVTuhaWoN5Igd1K2TErD/a3+6ubYYn23NG6UOOOY680cClCt2LutX
cBxgsoGGG8j/7SXG5we11SEeB95aa6EicuVL12Rx+E+v9q82x1t0eFwgiLq3CFhi
oB5b9dPkIcNA/YYn5o4pjhUt+a5tEYC2sD6XpFh2YSgOldSMOlLGnGL6pIUHRezw
X3pOy267slYlBcUBEPQgnB3npc260gRtLl8xcgGUrjSm/w0MDWsXHlglC+icmKbN
wsbzHeypc6j+OJZpPI9fMDjQBqKdOjngNuVbV/ZAM3894CQPJgmMb/yaCvguHuOC
xt1Asx1I6GpPCc/mj/DT4kWxku5B+uJg3CzXK5cK1TL82QXfylUdb/jxAtletJxA
Zv/Wr3joa1PysjIeql/zfPlw+yiHcA4ALp6rTrwYGyzi+tH+FMB1QnCOZfpGk4bj
ivDXK82KgcGPQIRdwy7OZ5oW/HSck+qPv4meqLDtkY5bAWf5LonyAgIWIAg1tr3k
RSadqUOT/BpuGo5T8VdW24ah6imtUZoWxuH1UrbFRKI64LhDSWZnUHtlmotFfufX
EYCH8rUCZgct7BynDLBFUrZ/KKdxSHLNn+AJRWPcu1/Nb6hL1+zCUeinmzkd0TtI
AnfrBXjvkKVb6m2MAVy2b4o3a4Wc2n0d0RWt0QEHP0T2ecCEscW+R3A7BJ4ory+H
CZeRq9oa4lTUwq/YBKMyWWVkmc8gY/Rb/wwnT/Q4WDlU+480P3SEpUeTaNy759Qy
zYWxp8pyj17OIIUAkcQre3kH+vzdRoiqMBbd2YrxKlEmdTDg5sFSWbe2mpzEUtr3
c2ppxcuLekkDQMDWpcXJ10E1uiorpKPuipGvwwtQJJF8sbcIllfp+E0eLiFZgqmn
eNNHjS3AfOnfKVo6ZvKbjHuw9n2wqL0qrvSz9OAJNN5/xkwPpW0N5mAcrQLPP0QU
se9Bcn3U0nVYF3UmsNQ7L7oIqmm0Oa1xthozuMIEfsxP1odcT+yA4eAk5sc/zdhV
cT6enac2exaZDLqXDbKZY6X+JHkNs5YCwnyjYv60rIGzNznAbkSwMWkKqFFAVyvY
1/tNcrNxif70UKAACyLqKHrw8Jozmy3YhWM6yYSSFirlW+ffrYciwq669l+PNGco
alNfK1CaF4hVdRCmo7AGeQMhM4XlZn7TFvKi5OK8xH+O2yYn6OzRwTRf9cUH4Nh/
S17y2Mzcv3RajQg7jaQyXciTGkK21R4zewrbZBuQzATEcfOiHXKtcrsMI26NDhLN
jZZFSmgtBbeMqaY4O5Fl/xezfN2D6GwmOHJ9ZztYhfp+QPhVqRfFatBm9haVDgBn
D4x/VCC4ULBKjqzHGKDrLM2gjc5vqq4jdMgUDiOKez+0RZR6wDvIJMQX6bz8GOuT
lJ3Ormx+2q7mI7wSu6Znnw+nyw1ceJprFgWpipIfU4lU3Z8rccDXosDRwEfS0Ufv
i+6p8kp9pk/JvN0sE5PXs6enjrDJcsRJHKFwNOYX583OGqsRwT/41e6tdLjQIyi+
WbkuBpGbbrQubErWiGTA/7hdbgnLJmMJOGdZqoIjhoL47bD5GOdcHVdQjsyfrl7g
mYyAuPFfqubu/KvawZR/mzL6QZSJ+PcXliaz7rMmr7mTXk/2V2cyoCtL7EoFnLQo
AT3UsEc7I1KOJxwDZotqP2MtojGVfrXWEnOeiUSv8+mr6UsdLrsjwK5LGI34hh5+
lLYr6W/25jtE3CL60tVcXVmeSmatZLDce70BZhXXrcm6KaTVLRAD0gwnlJ2ugRxI
pYsmSn/XkyJW0wrBbaZoB4ERrK5co0SsRyZMAws8j7KMH7O5USJ2GEtAdgeZVCpb
eTAkhC40ySpXlEQuqdfNREU4JzztZLTqLKGjTANnTbAI6q/yXOc1VTx6uLDk2/Qj
TOapkJCga0UCPV8otwUOugGQYoyBGPNL/eUxSabgYBHLF+wKTOkSTiCUE29Tb3Q2
Nk0B+4+Hp64XpSYbXBaXGzB3STld8HSnWk1ANiMPdeJMW2bq37mUwW4Qdt+KdCfm
3H/vSAY5m6SLjUJCTs9c/PcitO2yuKiKmjLgxoy5Eq8L1PwqOIwsZ25ib+PzJu7g
WEtbOjJ1PYPSvkTGgrm9BT2X7mMfu6GYGPMpBChwp4lIiPNZwMrEnU/HqEnUcBMA
FwDms/SR4dTEaI9kaq47TTn/aObneLFSFnRdGyezIzN495q2nz6JMQke/RtZ+SYZ
7M6uViNfH4qE7DDQ3125If6tbJzRwUosQYyxb6+1Ra/UemSCr+TnzlYjJFkI3Ub+
/JSUlBKjctKHi8rSnJwmNm91tJfAwqAKB7f4xDQ2KyjVvVOlOj1TPWyc/UYUmtgC
GvocgS4PROLUBDVPsjitExKiPYUkhVzeE9jY8u9FeUXA0y23jZiOp8Z48ZM6a7bN
gvVdCEzTedJH/pC8e+zsOffuhpf34oHvtEFvk47+S0/jSMLmzzfnk7yh3QkjzbYA
di7XrxpMl2vq05agLkkqyKXRyk//zkPd3a+z4pQZcmM/CDlTNz68o/pQgUE07afa
nNrt1UGVaN3CZ3diQEDNIMrWhsHIYmGW5zjfpybX46yqZcOJqCs8s3fxXZy+hSEL
+dYVt1alAS2ztQMqNGFdhuXkxpi3zEuTVSTdc4zbZyEyU4Kjkt0CBet19/UbkqLn
Qf9u8l2Q/pBlhTrE0NgWpl6ojuBNMjF0rWsObS94F/6r6yhamrTSgS1xh9tIBrF0
XSKoga26qmSwMTfAhrT+/Dz8wDOHii1Zcgvrcju5QcrsiPyTkG2wtHh47jIqJ4gA
20cX7jpKKJceCSxeh/3P9aEucjj5jfOT++BJsdB08t6AskzFKpIee3ND7GZLON9i
VooC1MkRb8YCuldF30g+WAsKqMgTy4z23L9c6pqjTUlT9UmS1w8LD8UPqd+sKR/C
yAkiCU0m+yhMZurg2H7ej76EIFiOKe2pNcKvZyi6wVi5dUrihXzccafBwd7rWnvZ
LXfzBzuR8cnkxVZ+o7m8PWMzJ6h76xWkPw/We7LuIDcSaX0dJMTNzLVgVtHld0bc
RGdffiInWNY+kVIsWXS2oXD0BC0nP9QVsULfU7BVMxwCxbt222SUgwFzrn5e4z9Q
+vaJmFA2HCe49qLcMU7XIiR3OJ5xDzmkgn4p8qGteNjm9/JdPbgZNp4jlCBVaorI
DmkLkynMpzXXcfU/xBd+SzVIzaXmjDoYtcg0X9NoGSVjPbN8PilJewIBS2VKRjk4
+1ZBpPq4oid4ZgMnpGDpq1ZJXDpbTyinGxUGxEIRqUNdJ9y8VM2ddZ9FEvGwnDqI
yNTqIoRHC+oYPbo0d9wsIJPYUKViBw5YrwQK+RrlexjkUYAjLr65hSHPDXP6h7TZ
bmX2YChZPcJBQnkn4FIRCKftbK7nym+LOixAUZemuVHohxobR0fTiRYPIl7YWtSz
equNiGyLNeNGmvdLSMMhqQnrmGtO41bK/dR0Fokp0MFRboSz2XIfEuXP9SlkeRLM
S82Cip0V1oQMrbDFh6i7QCWldJ4Flkh/SQloKJIYUCfQO5DPJ1Lqw83YbcSTETpL
s6AgeF09rYmNxynRQ92kRVq4XiGzSZYsRoScyp6y5eVI5Y9CdYl5Ab9fe+GIr3nf
MDntcRSqtLggnRSbMeZBcVwY5C7wfkvOP/F9wEFGapPAjOrLp1tRWIonxzLfz6Y8
hWbx5TTXFh65Ko/RgnR36pxlMLGhCufUtGWfXCz+N4h6Ith2LN+csHjfb8cNghI1
ynku8so9ZuSQjgMFB6WQlhrUoVVnzYTzIPLKqPAIGEiKg5A0oaPedvw9znF+y4Bh
UNh18LQ8pHOjjdzgaExY2B69L60U+uYt/dsiZU5OZ1mLKqNR5FKsoji+1kR0qpZf
xSRphz3XCXxUUXHnxwbNWqF0rqXLcuDqbXERzTRRVrFb4VGfKg2fZ3KPpoHNcKdp
oBMRr+edQIggli2KruvijZvLYXPQTUuMJ5hu+42HKuvwCeEBl7yOu/fqQ5RzskZ/
MHyR8R97NN5kaCu2/oAhivI0xZpGD+K2uIEdCXM5DnhDhfmZokXR8Qm4um/aG9KU
z2dzPJBYVHvuIEeUwMhrjmTVhYUMLVO8REa8Hy77IRk+qY/IBCRBQAJDPZwORvvi
Aivo07+d9zG/Z98jk663EGrAuXoDhrfaYPOkiuaaMcLgB9RdFqmEw1zW2CTQyxtm
n/2Xt2M+YN1zXYjbRWr0F/0eNFbhV1NFzTfnOBD7u5SRxgGonFb6tT6RME6nTYxW
0yKwrP/OI1HdYWnonE8Dm4WUaE9N10ixPzfNBQbyEgeYwzcPLTR2rdCcbWaKYR+g
jEN84sLaMzY2C4UmZN72py9e3g+Nb3eiR+d1k0hDRoDaSbxNddW0tYV0c66EByiO
eNB4aUOQGsni2Bx2tVH0TsGsIyvAufBelO5xctNgpgm468LG4fEjCT9dBubqFESC
d+NL5LBS9RZ1Bi5FxrKpq/VeNcuzyLh/olDwZkC0bVpQ+/xnvuczeoDi2ipBW65s
pk63yZLsILfWnhJCzllY0Dlhq8TAphQqnQ0hzhMDcLHkICKnQ8E1HgOKPGONTvdW
Ye0HkKS/KcN8fINMOLpET6uRA7Gzl1DwCsQCaLiJXjA1mgzfrUTZ/dzhBsNfnqH7
nl2qwjNGDyGsRPSS5DM1+K5C1sF1Ws62iTAVfhtJ+iLzIFIhN1k/ON9zB1Oel4VR
pSMoaKnDTWJbDmtrDIPkFW85nXf5wcdyIBuMlYL7k1HJg+gHJJuI6jzWz80vLf6Z
mgVL0CaRdv/AzDhi2l4X/iKXhF5ZLJkDd1tMKmy7gfjIKgnh6Z0n5ICeMIJQgsaL
JlEKbVZ3loaDOx+MvlL9t2hqIBsZsV0IJMpp6nJpOHr6hDroZz/MAaxpSsMBddHl
f7e1rN8eHRw0az8Lie3bc8ZAJBx2Cy8k5Co39q8ZeKaKBc1tArr3FtqFC1yqarKi
f6Dyh6ZVti0phNODmY6FwzPw2lzpJANuCR/JTStNsGh65Tslukyab8QU7rzVI4qR
ht0bYpqz/wkxAYEDrlhj+yG57U69shQxsj9E7GuBFi2pU0ZPbxw0tTLXLmu9SfGN
4sIKKQT73nb0c84MuwpHNuh/ZyOxz7QFO1UlW5Su5YIQJWTwq8gsunt0zfBJpewx
xq94NzFGTHK5AuF0+TVXMoWyDOSALOKsveBRdQA8Ct3wQyhSFBemCvAaBcxneAUN
CUCHcs6MnGrV5OKwB/greu7Os2OzGE1X/3vvEgOnkJI2xCrekloXNZ51PbCr/rAT
daxqDzqRsI7marepWVvoDto0VpBgZG73YAmtGFjWX0Odyc2RSz/z1Poj9PrYzfkt
MHyOodxzJa9rQYB3/8yJAFRO0btPNsyFd+hHmWnHaSKAf2phJ53YoUCrXs/wcJWp
Su+fw84kXIp/d8WkSbQGHSXkKucoCEsiSV7x8AakaCOpTgeA5xAlZ8FoiWfR9T3Y
TBoDvjne6iq/SvlcFvHv5PpoQDWrRghu/BQm5mjvbKCQlyjaQILcnyrQPjW4fUeh
B14mi7YYB3kQrsW/9vrSzK6B45tiYDIs9ArieS4r2hNXM7J92bB70A+ZmFdISCYP
M7oUgaL/YU31YZ4X6q6olAImDreVLr5wjMPkTQOqzar87EAaE/AlFlQcp1p7DZqP
31Utmgjsj2iwl7CcBQgXiRdN5eL0PODyxhCKRWAp0NFa1b+qGZhd0HzUaCHDurR8
y/jhoO9kI8VLZtrNA4Mrl1M5RCBplPDTpY0Do3xhMwUEHKSW4pqDekbEelLAWqrZ
vcPQJwhM0R+EeKN80kwCEeAg2AIgtw8pwWAYZZfDuKy4MNtC2cNNuHs2fA/gdWTg
re04bJUoVtTFyHs8iXGRqH3FZ5IoBWr47EG3E8mq3cG0vsp85AFUpFdTwd2leCf2
rKFkOJk2eE+XIy1gVrW07ypVUTtO+k1WT7FIRGQSw02Rx9XXdNnpLhxIlPcMx2sO
DSib9EtrCi4i3WK6z3KwH1U6CArBPV2TKir/HpWZ8Li0Df5jLGYAYNKfeu8EEEfl
1vEV0wIV0Mc0Q5HIB0k+hpN8HaoxFINedemAcWUIZkYPYzZtYQLE9ZV0FZ1RXnj9
1zCQIkmDGVZt6FQV7YCERmfT+Dq8hd57AJpiA9tB5MT9RIUhWii6M9L6PZ8zKbqg
s+yPKudU/yjXXWyVvhOtlmcVsMfNrQsIBcvo3YmU5C9XyPkvuFWcsfZ2QGj+5t2o
BXJ5y51xzwMyH+AS++et87Ib75LXkRE0Quke+dd4/epQeBGBJ1stNh+c7pHoMHUd
4njBNWef+2BJ2408PiqROeCN9UG2Eq/5kNCcZO7hjUr74WzoNNzjBgK/l0cuA9SE
bqXp/RrF1t2TFtHszRQ6D1fdiEsdJjLFAUflggUUcXFeZ9ec8z+QJyuya2FW6ztR
XauhlmVAAKc8uZrWetNtyahQG9qAy4Ikw/ZDIAChi61Xbc9T0qtxygvB5UNHhqZ5
5oyASJaimtyB7H873Pv/Ew8QlNChnYsLJK1fvFQbaaTWztI1dyjpZh1rf94A8UAS
K19eEqDLi6PSGpyXzBa+m1ttG8lXY/Il6xP7XW4HbkLGkr0zyfHqul5HArnUUaPU
vNcA+N0ZMfBc4ldi5bLXCpp4VWKA174NWXUPUYE60YJfNncXCJekNQjobEnBR0Gh
eeiozCu5VO/1vtCSUZf7ecGHjffaoR7uw2Cp8CqYgPJzzvLqGyuJ71+yGnQebMZO
8dELVriDbc16bdUXQCfqBjyxfGWUMseeHfl8hJpwTTsb4tde3dkg66j4J9Kwcn69
/wgs7OD0BVkuyKm02cmRPWyLuLIl1DKAGHbJq2+z1ukuPylVZVQZaGMK/b7TE567
2YITQair1GuBVLBgD8CYP3P7U3SgCWuwigue0sV2qovgkeQCDLh3w/FOsW7+370o
MBYvaArzZWYfzQA8xkNMInr/dRsVF5v6MAhrYgkoHqm/m82EHnirFrvF0BvdkbZU
uqoYzpO+rCW4BUlD/sVd5o488thMYD0sE/riFfQqeKjIQX+J3dhMNFryM2yjn/7s
7LtY9sfrTSWkeW1ZqyPNoo5rW/fIFXETWGaxLUacHffwsuyFGWJRYCtwXXTK26JF
j/T37FNRnHi85og6Tn1yCDINdW5OPOc6+Dpq+4NWJforU42i5KNja0/WQwaD7aPy
5TB3eiVqe5iWFDqIeQLaVsEh9dtTdmP0kjcmRKX3MEBT0oILsgLHRAcGnv0HlhJz
qLojAjzein8I9kXNppTCYEBkt8240tXjlql/1zQ+pWMxyYx2Wks0m9BKTeUnQ/Yr
zKMNKboXcbJzS4WbG994v5KD7V5EYw7ruRw3IkLXr8XoDXYWrlguPb05bxVwX+Hx
QvtyR5YOvP0JO12dpS4o8JC3Lr3dipLMCQK/n5sbeih7X7/AiKBTnRmhFzTS23df
rY4yaJlTC7srRVDnFwNdCHIspVDkivuJgWdeRJzzW24G98rKLXqOeenItSQdpUF/
J5EtPdVROrvqLdTNHgk1eGRRM0aJR0X4Dy5CMSmGUV4BZ+cBWB2JPyRWvc6k4sgy
58l8GBgcRwnP8/LnpLWcDM/FbNEwvA5o9ffylk1jcyJNkriGWNO8jURCfiR0Kn42
DYAnkB+cTjcC9xfopV6ODS2gF8g6NOcS1ymMbRj+UGE+gboPqI0SaAZMo8m3bBIV
CarE2Z7f8R/fdR4xvoGM2m45fm4+kFTYcX5Ox/Ig/XhfdXFGpPWJdIZBZNXRQTnt
a8opdD6uv/5gRRkm1RotDDlfZR3E9X12R64KfiOW4Q5eZPwoJfMOXfk4rbzQFBmI
eW3AKDnG5u6bjOktVjVMHjl3qYR/PTgkEkLnPVvaYIGlbVxAJnv8OTNoFEhituZS
cquIZMhqKe7fRlJFf8rchSGjFOajrdydwdxAMoOzMINHh0jwJaONvaorbGTUV/tE
QNL5Wdb+YqgW0DcK7RjAW3NQO8xCQUo6Lc/1nxgGLFzp85YSLzxJBjdoisvV0R6P
oMcqK/bgd50m81pRJTJV5Q0MGEjKu+bFiO6YCkrr3FQxY0v48Bu1wOflEnYQcPmD
IQbQ9NOXaYZAVJmQ/m+Ist4OQB2AulmEpuo6ZP6pM3+4LDhBmZFj6V5I+I7oVVHI
Vr9j/srFR5XQzaGAQ9rOtn13uuwEd+2ZJJOPpBMcmQcSnAQQ61b5w8ri9Gr4ci6s
bIG9EDDGjCDCgE3l0zZALFO+0vhYCD+aTuvR8qM2et92++dlCSKKPGxOLM96itxV
ChlBYy1RPbPOkpHevXyT72c+jV5vKc37QhZU8CBG7Bs/wLv1FK9AZ0YROscq7E6U
iai7qSO8K+p/3MwbyZ3B6u8Feg88JiBJu4hRvt1A0uZgmh1abDKYXGG9jvFgJuCW
Zl6fu2aRhww1IGMVPHb/7J6GZT1HQAG6xc+yO+OqSbXvsY27wnFFCdGV1U1luwWY
LXPMGyASl6Notyjjx1LZQgeHsAZshBHwOxf1ijwMIttz1YTwP35fdnHsjMvVMglr
LrNobGof0O3ZiY1MenQ4b5WyyIfKbpY7UsQPNjQiMrv6zv8YdPBZdEBiOiOXEqhh
SndRnJEzL5Q0/L9A0rA5z+a2JwgkmrV/nrOe8BKiD4wzJTwLuGK2npckmONapPHr
YjNDTp+3fq6lPla+pv8aljz/LSVxINSzJWQ/8CkzEjVpFwjHKBWukeyWyw8zZB2A
JXIv1GQfdhnllcpZ0HB1luXh/4nu8tHYKO+Ll0xy6t8bnrYx6BIKjSOePvi+ZvXS
7P+UG0iF4tKd37cYgdwe5MKYtCwYR/vyitwQK8P4ssS7m1pxbWyTg0JYa67UXdoT
4Jc4TZOBe7rLUwhrMzjr+qZOKcNwtmx/sK+s9apcY/8LzOFldeCeo+iGhKa/L2+2
ZV64tAR4iRThFyLgKrGvu6Mp2yJyHnjMVoatmk9w49F2ff2uq28kS6x+3mDplnTD
/s4BRS76MN+I6A3KoYMt9NlXOv4hP9niKRHAnBC06EJb9X7+rqvykcXi195aStUd
Mlk1Lx4AXrk+pXmZZIf8UL3zfGbc1ez3Jweg8CpvIf/JGpWC3ZY71lDgGr84x7qS
8hFnTv5YJRwbynJA1UotdfOgiVYNImJbKAm9BPfuew61SezxreVzvK7/Giwapw+L
5dsOVpGw8INZOwkwiEQTMa/tgFxecV7JKPkwmmZsOVagbyIr5Zqgx2jx3Gnw8D7z
q15ppxtBhvafhAIgE0jFvvrFG1ZXSsDAbv4qq1a8MShcmkXKDM2AySn+DYNasJkA
Uhxu0FtHzn25agUY35iOFxB+xEaYGITBuAcx/9ecInO2pl0C74GQWu81LC71rcfP
D/+kggsfLBzMX41UTtnM7Tlh5qVhsuPpSo9dUjjzfhNI1Wu4RorNqLqP9qK1fRGH
w4QOKbV4Kht9pOHlTja5Sg+845cJ98qLfjrqCCfggMAhPghsPHrKj8e2vpu1M+0j
Dy7oF7ICi7zAw5XooLPGAwYJ7O2ZjKI+rruYQ7JMV+OCQhDyfXCWlNU0MLgwFa3/
d3Y0DboNQ3dHpW4vlGowJeBq3XPNZVWOrUUfmH1YsMgNtz+c1j5ju5eUSqrUXMKi
AnS+5UfdPVLeD1+0heCvZFOOYbYe6W7v0ugQ64O7BuXXN1UGivyeOrzClsOI2BzH
2GiswnUcthkvUhCuLHXSLzzCQaZzG8FvIzGc/9ErByx1zGyHtbrnay/oH98Fhieo
VV17p89S3RX69V2Bp185DtTTEn9fj3m5ynj6QYdhBKnZ9E2vF9Df23j8tR+NcXkT
cu4cqtjuSBua4rmKLK8sx8XLD0nKcejduZTMlVORBSUpjFuqp+q6fJZT6mF7V3ya
cQiadZ8jzHMYJTZHvNaLylEQ8A6/jJGJg404ldDcdGUIfrh7xoBhNXo+hVWlVpdo
z3PZ857zFEsw0blzB+l5qRvMK2ssAtABTcW9ZE4xlet713MQ5BolTcsdHhBHZ0hP
l9OTwUFOTwEfJjXu49fUr1ITPy4uVBh8fZ99LSE3ztVU1ZzmrQ1JI9GnMvMVpv5r
Q0eWyFhOsTZQO7whnZcM0Ch8bFLDlY8QUmHRZL1wd+xeIiYtrMRDKiC5xT4OM+vj
cJ87R4OfoPOZmRc24r3vQFARNFiNIkTDk5y6rNRW5hsch+/9RAN1o41KmZrjO8Hx
Vl9TXgcUch7EcEqdg+FVa3JLX56UvF/6LfN+7T5/fWBi8YBmn88ePx0rbRaI9RnO
fU5h9j31GrL31Vls5rQzBRek4seAzli6H0cBJHS0L+NTmqvoyPgpMkdKyrU9uItx
xIx9JzSzGOS1VQwG2mgvWF6eLr7GxmZFcSvSiG/kdgONi3ITMuskqzaj/GUcjhjJ
gMLMjTR5ec7QoMbGbUbngTVzNJtRy+Nv4Bo3kbz31ooixDqz4OuKlZ2LP39HaYNQ
r2YpRQu4VjBV/AcdPalXyLmLlXFvYM4f/icdjex6etL7u4IdVwHnQyqoB1S7w9xN
Ssb8+QaLnvNf7NhxogaRb3WhiNY9Wo2bdJ0IjXK4/OzuUIxXABP7q3WMh90d6mA9
KjjZ0VwEKnKC7EojQSQhl3MYUZ/LEMwV3RoW+YKBnqwUDjg269giNsV9hU2Wft1V
vePKFJcUVSN8pSM1OFv/Zsq8foX9feVncbm4xfwIWs29Hhqm87Nmg/8aZ5OPJXnS
Esn5RewSJRDH7Aq9wJfShDxS27Sq3ol+S8xqvEfkmO6joO5V2FG1ilZJ7MQgnkfZ
TdVYF1nslzGtVw2DlXiSD/zU0W1Yiq9aMTCAP0vmJQ19huqRsXUL/zBJ0meyDchc
FrgLDxTCF0jGdrynaioC0G2j5ve2NBXkPPztpP51aMbY6T0pZ3Ehjf49y4kohr8+
VWKqANyufb35RD8OTxdDhIY03po+q5lvhAQfpNgYkHxAab+fXwMFnxBkEFSSSylN
KYAi1dHbhlkAD7XBNypcirQGz4BfUEQmKNjisK4Sx0E0NppkVfWAEdr/HMl1cBEA
tQFDqn5AIcIFyxDVQnUQje4WKnirAJ56bj2GMqzxLzscIuWR7IoyiUO596wg4wS5
S2fiO1jqMTVeivLI1ZmMZte7Hcsh2mF4drlpr3Jo+X3nQsKz1mDGlsyLUC0O0Hmp
ozudBumvXt6QFbvZ/ffNQ5xkT1G60pCBh3sjabqd1iWnTWUNNJgqYmjzWnqydOkA
jP3kSqb+WR1n1hTJ5VYpXNMKeN6TEgmy52kcgzK83PGS+VTOfCvUu4u59yldFsVn
RBwnzh8mMPF6Gy3xQ93QX6fTO/9Gt7ieoRmcE68CECcnIBvPwOYsQoqqNqKm93kk
3hLVzhvHPeDFpUHG1m2DVu4mPE4n3jjpRkL+kZQNRMYUUcJw4rcKkZ+iA55u8IrK
jOd1osAyvdtYOQvE59sNippY5VC6Vm2qWFRrJIguru3pIo5cyZBba5e29+K2Gwn/
cyGjObPW7+JS6ggtdrgw35Z+q63qagBbwlTZglovk8tQIcpF+55BakuQQntE8ANN
jTleH2sWQp885S5aLd7mrO3hgFfUG0XdUcoVuRhmwBQ7TXJkme3WqFvk4dcXOdfU
RB5ORzZw4UxF2Gxcv9UAkEe/7pAaBxLozWhAkZ/z69Cc5cZOQ5GxedwvNjXUknws
SEJknm+mqmh3ARClcu74FY72lDjSZGiy6glgk/AOFwJ4b9m4S4vhkYRFgU1/Z7Yd
ttCv4HMsa4oOgc77jk8PKpvOZBZdYh37X4RdSelmE5TvEyq87Jseo9tQqE55albo
aSMaFIKkk50doK4JlMHcy7S6RZZbIGOdfMByY0yhqUP4NLrCcLKHPGG/6AM3YtyH
Z7y3CDK14801gj6mP1mPgRm0C+2wTYXP0VLlnzGfrWnDmq4WYRPkxyGoOhCo5EtA
RVQYfxYlfnYUMhHNNrB2Ba3SfatwIO/wcIqUrnTj5nH2pMha79QjKp9gBiLvrSOB
HAkBzBVAH4SoQc0MEdDjw9o4SL24HAkG4hPW4eKGO/WAlmn5sz97OSjmX8H++lzY
oLm+VfexbdOhr2fv7dKSAA7Zbk7rAtWgfSILPTijAEjMgZeD8wHFfe7t9AVI5b/0
RQLDye6cghjF4BZGqlf/sYRUkvz6CpWgyHs2M3Hl4N5C7EtcKTW5ropR4HH7kpqD
IIRndVw2JvhzcRif6PnMiGhIn30Hs7ZXLZGnnNkGyeSnNdWkCqB1HEkWq8DiJktV
A8+lMs145eVyqucT4+9UFwbbx1AxgoelpVLwRmn65fD3h0hNwKLt2ZA7fKzHhkye
y59r24hA9k4S/R/s7+2A3UULsuBnoyRic0vF/XDIrx1i5xDSt3cwknJzb3gAe6OH
KPDZdgBtQXVmSsgZZ+ynnsm6bkfYwGKs8/rOz8t2HhcmGT2dRTTJeZaPa0X/FJAB
Uq4lj0eAH589oZD8DnxKpTA4UG2Ue/g5NlWw591jt8g2AaPeQIQBci/RGDgG+/vU
ys2HO9d05qCQx3Jyqnuu0VgRcmi/DclkSTSAs9Plbk5HTrGtbeoJ9RmX/XbY7VL1
hb0bJoJA4J28ai+1M+rNwXb5s7p5ETh2MyKn6ZINqJmVstbfJTeIJCQhZwTOQnla
ckBog7yeHAK7LsKkFiWg9nOc3k4M3wozuJqkGlvaUn8kKIK16QZCxPLbym8+AFcm
D0w//zz9l2Sq+Mt0Cbcj12KaDnKG+iATT+PjlpMbDIpPOwDmB6+TN1w+lPSXhoPd
s5LuuZtDIXNgLAAX9GrwQPFOjQLhSNv3/R12ZsfZe+CRcE/7bseKEWHSWjol+9iQ
vfeTLoowChPu8a9nylLjQ8puMR0u1d0uhZqxQrTMtE5CrX1oTi4hN4jho6tra3fw
7PMLLQDG4j5icSb3rkPFBkDf6ywx+LwG2VnyVHM+ywNC9ipRmi13KnVQkIgR2PLi
SobWjEbXkJyRNaSHB7QBk+k5zoIuOUA3VDeCo8OrrfI7JembBDMAQE0190i7G6kZ
IwPrHyOHsZP1DWuO9y776RJFYr1H6ruCUzqV1EIllmlNCNPm33eo6txhhnKkD4yk
wk//3PwH4hFh5MTXJO7uofegE5uYEu/+3ADWh13lhlhptSLtB2sIp6XbA9ShUk+v
6l6yAmp7vmtBLEJQnN4pr4QUxUQDzLOV7/vAF+mJwBMmMKY07d0JI/Whr892HnND
uuZ6nN0P1jdENmMwI7dC8t2YVbb8Pk/wpFaVOmNBpJs55FAp2K4sbW5lTPdlr85V
WWcxJfYArA8FsLswWLrJnthGWo1dqXuV1wgM77N3ZLtcHJXhU+ceFDcwz9oBfwOP
1usZB1KeUxtAC/3Wqt5ryIJRwHPA7y93qduugiosUKiQWjCaw+aooADl2UXMOyZQ
gk4YqPklmCD+gruzpxQ4/wXkufrJcfZ0P5lb4r83Ukx8slHEao3Opvp6kunhL6ZJ
RCKzozWz+YalxSbk9vQi7vvp3GcmX+egOwErZaH9mvN1e3Lo3ScLtHAN9Gt8upPt
EoTT2znBi/Y44Gk/57TXDGiLSP4YQqrWFM4OYePjc51xePxOs960fg7PlD/2s/mR
8NUTliUy426gHvxyogx/qJmAGY1VVMIe7+L5WFLKtrBiQtCcrSPJ444tdUXK4Gc/
5EbgS676ZPm8ZDP+1B+pzJmajod0OwrGSvWynM+AXl93Wsf4ha5Unbo5THgAsOQp
7Th+9Vir5zdr8X6RbM/Tw83fHohm1//SIZHKVDdViVFTGbrDWPKCicYs+kFgidnz
isyhWRbTlk/M5Xsl8Fffkaol97/pmAp6Bw6rAqf5d1WXgFSuQ9hc+sCzKTHmEz52
A6c8s1fflJYuF/57OYDc/sZBhn4H7wbOaDGW24aJWzjpK+Ty9ZyF9A7FHleSfEp/
0Bag1VKxlylcjPweR0t+ng7qxmnO6fRDY2514ElWm2rPr7dzz+icVX+obtSj4P5V
kEfjE98aRGDYT4t43D2wikKERVY07zduyjb0G1cV5yi4zj20ercVYEE4B37TTjef
rOxfFAvWDqWMLOncJtHCvjqxrMjl3Iy9c1MI6gs/RcmBX5P4SC1WKnYnujzb52pq
MDG5DaeHwFBLOnypIyBp0GhZKF5S84E3MoW+Ixw02BQZjJJizGQNqMOgXDI3msal
qGZES1tH7nvCWeLExlqPjo6xTA3maQce+7VqdcFNDzxrZK+eIjmSJxZSYUJtotwp
GYKUI4DUS3QWqvIrxRE5pGrbgFxOooyofmzXKeYEW/MPLsN4GvYFHGXtQmmgG7cP
s5ZlTUamK/7/w4ExhXNm2dVBhkORT6WX6pQKB1Z1q99UcW/EN++KRlk8ZDzpw8Lx
ryBWH0rkULOW6QVsW7NQwNVzmYibOVl8h2A4jHbIOHAmPwWWMDHbwjMSx+V9iY+4
GGoC6frHPGNfDr6uys8JS3b60yqkpH9kVaW90UPh+DZNOwR6I9CUbG1qy4Z95AAI
6M3/I1lhIZthshiGIqBYTN0ZucflzyYJs6azZwubGTlPBOoCE7NudC3xbzEefwvD
aK/ffFPZXzkys4qb9WkeHtXmx6jBPO2tMbUK3VoF9QfBS/9xP4iMKfaj35bcbgd0
XS0+brTSvXEQkGwNY4MdXT03gE3UAPxKSwkIvzoOWOSZIcX2tYD5pLZ7iXPd1E6y
85IchaMOnt/JPCaCnI+Y/siT23WjzB1WMuFFitmhOBFueXodPhI76klNlc9UvgGX
vQct+lv+UypzhOzEYPQKNq3FB+q4Ed4ly5rYZygxC/ZvPlZm9cL202vH2UXZaLxO
/NTpfFSDDqynN2khoUOABegoW8cqZoC8StCAZMJupwOKHAmqwiPswwK1Ig04X0q2
EEU+YCppeVNIfokP9UkZn/vkJXj9rtdybgFEQCWLVIs52W/DYZ5KwOi9i62T6567
h4RJg4NGe6crls4cAfCztHbxojvXAzOIkuRQ+8huce1Z/kwCo2pYv94MJ2ku42vL
6jMs4cpAZqvxas/vZTF1QVp6Rnsf7kyJdric8ccyIvn3TNG3g4CdUgTnvmEohTq/
ZnYjE6mJKwD2FEftw8OPNKZHY5im+qVnhInzhoOAO1EokHr/j0YLh/MTT/HKQxJ4
LBKmlZw3RakoU0snPuEuHg2Fd2rAo/zE7wXYMGfYNuMWkFBuf0p9+pnbMa6/8E9x
1byMmzFVhifiu2/hCjaiUrMf4g8yjqAfMw2AEf2Dp2rWfeaG+554uy0niirH74pj
R0WDwcSc5QiLuXQYRb11288tPmUQA6iInzlL0twRiGfuxMeSbd8zPMba/I8ksMxe
4uOGJRHcvy3duB3q8RhDk0goU/SJTjw8FOiJO+GcddImCsdyFkui/yYCeKFwMq95
9gPwnHJ7N16Fm9erud/7iyiojWF02DmhfBZQ9v8G2E6aNmEI8nukLYegvGReQmzI
JbkXXf5YQ1h3Wz1a9C9cbEuvS1NsdYnSUZW8iWoIrQ/nvTmlCNNhol7g35sqdrww
Bvlx5q21MX0zgNDrv6477mt1L63nOXWLZl2psY6Tih40th3FMq8R0apMbBwdlusR
c/EQVkElaqtWjxHrcxDJV1RaeqGQiO8iWix2OJq+4UqWSoVMuDRF96wE7fSMctoW
n0n074HiR/sosHbABGgoQ8HQorklECJOTyD4PfnapIDFJQZnpi87YqQZ5OqK0KBK
U9PR0zhWcB3cRfrp85WHFFov9FKf7KSnLZowDGwvW68O4fmXt5sUFLlVz8EENWf4
qovz/2p71On/aFtGdrVagUqCNuE9kTKI+KX0l8rE8z1EuimRulVM34T+IRRoBHV2
4dSGwmwKJT8QKw0EKGnA4v54grf5eKmvPWa2/abLKcD0OqQnrTrkNrhSGoVhmkGu
vHOpm9l/J4ZtC+rGRs94Cm738lFf/ur35C35WVB48ptwdyf4K+uA+G0LRvIPXF1/
6IDt1GnSrhCYt7n1y5MmhoqnfAOtXlPNKe0uugJCppJ1ZWJtTXDs/EjRa5lcMydY
Z8EnD3IWGinD6Tz9geBgbG0H8ck9I7aQt5fPm2rZqHxxzLPRIOlxwQl+NydaVE4p
3MfIojv5jzduteaWjeG8NQeiJDVpFZnYTCWt+wfgX7XqTAKucbxHxfpmQ2umNvob
XwKJVV6OlDQmGeYkFypbb86ca12YIHyhvZ/9vfjG+YsMi5dxWxqq7NIeBwe8k13I
Yq3aRf3tq/1DJxcXAVtGn1Og/m0nE2A1Px82rNZBukIXo7OVIfgEt+enLaIaWjxc
42ibFqCJ//yXLhUc1E08FGL+D6UcXlDz6uC0FyuknAnQJBZaZezZRf93Od5XK2nJ
or+hG+p5vakmtYHCoa1vZaNMk1T8ScAv6RUisVWgpiVDDawyN9sYgFcuvWidAil6
B1rFlm1a4HPiLOvB6VQ7TzQNyeV3RxS2YvG1K3x8wcapEIPia9N98YSDHFP8AKex
N6XT5Ost6wcO2PLqmtNo+8aKs+Sy5LAQPhlYpjM6fAlPbQso59bYhDN3tHjG0x/V
gdRMonBpiWaT46LbZISuKCgDAWcY4My4KNyHbisZpgkfwHc8isRYm3BTTeTEO82l
pOjtxbB0vIYTuxWaQ6uOwBF3NREDREqpcK63kvJ2wwg4ZCNOW+8fCOKddOrLxlfP
7lh4/iCydUZRjt6qhl+w8OFN4FzwPe7G04Js2hYwd0W+6x3UmWvzAzyH9CrIrHvB
7T3Vq4e5mxPSN4Cl5nR/7r4/ovzxbULb4D10JozgMrc6HMakftk7JTSsK8eoQ9Vc
llkUybPUrPrh2NaX0bAko5+dV3LMn4m455nuI3Nsvs75T3JepRRWzYnSe1eTLJHg
qgVmWVripwl0Jtcf6uecKa1rEHiROwkMIVrIm01OwNf9LhiOAKkuxyJESMDHlXJy
pXLANI9Y03QfIqZRVPthZ8Zc3FPTxvvao6QBE3Dg+K30dfZq4sfKimrqzO5f1tQG
EO10qTbRly8HzjDHDlXWxK1ctuFnGdG+nOSCSJI7Ixfr7bypP27nqaoRVYlrmkgf
VlnN0nkc9jZD8PmghW8wCrshYLutY9oNVU7NRv7mf+ROUOUx7UI1epwnj6JgVVlj
soTsuKZJYtzB5KVPS3PyuyUzVbuJvfW6lSdAID0N/gB8Kyl8VqTRJTRodl7Xq1ic
488FUi/2XoppOVW/u7yY+PQDbXFgOcQtY7OssTJt9IidxrtqMndo4Rd9ewrjDTcf
z0oQh4sZ4ZSYt+Eda7bLDoi3Nl571pW2sbo8zJ1gq8CK7kZ8f9gKowEuEDWg9sbP
jFf2k2QZbNFgrWJJiQyDIbOnfka/4wee6tgzYd2pHWXQqLSWjJSig9fF+5BKbSWK
mw4sQ9PobkqkZhreEKUMHwhrrtT99s9z8jCTEpxIOnZQzPoxZa8ErR3u1gsTwMkB
vdZbW4Dtm/c0TOpeGXP/Z5jglg/lYiFLSmlWvtku3bCSsr9TDC6+vGolDDPRaRrr
3xKcWsljsVgW89Z0nOBj0TGctPFP1OtmU5FWq9AgV7idAZBJg4d7LQivS5XpnfBg
SiYvLMFbwMtASLiTEmTu/8ou4w5FZ3lvOj+C08GzQNiKGHw84z6TJJpdn/Bk5+Tz
wZle+jQ0e+cYDJw9mAlgBKMsZNAsroQlZq4eHvJla0BFlKCZv++YESAHh0frjwRk
IOYlyg6y3ChjGtDqKQaAkaYbUJXQ7Mj/EfBJ7lABpdep/gcBQa6FUU++/vgdzQWt
UWNBzOg590dMGoaCKB+sgsRDVC11mftNp22eUoXNTwQ6VQRuyk9LW20k8Rw2ezEV
THphJatmd/WNsdnPpMJLAAYwQbI9qMgsuCA32R7nqrvaL9BPNeQjmatcvg5zns8W
goGlB50n16uhbW4uJVtmZItPrPOJfbiT5q5p1VGd6MLKl9n6Vxh41VLtD8FmRv/q
Nhw2d59uoL+h+84l82zkm6PcmoloGAVL0oxcYEzvUfv/UhMI1w3zyRUkdlGA1hhn
Q6rA+fymvWXy+pirK7JQTJt2qPlLSZBQ5J9Vy7QPLxkOrZQO5bSCY524zjb3SnTJ
r3O62k9yLq7uEoS5lGVfZ4Wk51xCBgjt6h5PavN/+NudMAiWv7J30CiWtb4UVmad
NkjSO+rTkdm8XxgNC1fHSY2w4LV+HpJJIFbVbjXuM3iDEPhnYz6IW6VGiYu3XqRl
StQi4jOcRGbyPQSnp9wBstTYwvdMrsLunKwrfpKTyS35t4ppKRzrT1QPmQH0SCTl
wUAEy/Id924Y5L2mG75i5s9FRiEbjJ9YNw1d87umW+TsgPpgJK2rOlgUzOMreUvM
itMNPfOPfC+CPdW0rnUyNU5LYqqhGJ3m2zmnVBuH/P+igHXH7i0JbXmuuSxwCuM/
1I8LBP2FbvWlWVdkqwpfWVwjidF7iFBDyqhkF7eYxKsYV6ULoY5OCMCqFLqkt9V5
fCmf4YuMW2UesIKSR7ATosuaN3+P80+zlxu4SDcIRv/kY8LbIP6vNqUrMBTn6N1k
i+hR+XcxgZvU7/x1Bf1eNiwdVHg+UBzBUcF1fTD/Xz3n2V/qr5sOqhrM5gYtqsqI
4EiQQ4jWH1AkWIMKKWC3U/yjAgl9gIyIe3T4xfoPm+KRtBs/8Qh/Dl1aXzTm41KN
F5n/Dc51BooJrRqYu3LJtGw0xtxAtIlE7US2wW/DWV7UeWSaqUTs9sLTKbRvO6oG
lxqHNwBVKedwdDMSXzTtqLu+WOlVos5Lmpm2WXoSItNdyqyENmnh8wu6c7q3gJh3
iSZ8w4ab2vbhbIpX++82Rj5C192QTM/wEXMoYSDvbF7LDoYZfq1Xn9VxYu7GMrtC
1pfVXOpeuuY/+NRqGxRQgsX5sW9HEp4eQdbBSwjX2ivXsX6MIBiSGGCL6pplk1NZ
IOrIpWXwqqzA24QYDvS7aPiA5xFwYqQB9nGz4tyI9jp/+AhXuqgEPDnJTQHMJInY
L92MoAcJIqYHs6ClQw3+qv7AZSRhgip4zgfZi6iGlZ5qWWjgcRbqTyPpX3h02ett
9xrrI+++rTAnURNHizXjKieHumUJnRjexyKLxzo1lExt7ErZuhMNY/eM0P+wKiTO
7IE74pH+2Xzt4AMbpcYHCoOBk+3CsGpvZAehdljv01TIGqrOGfMzaRr5ahqqcFyr
uXNTGt2NuFk4aWo9MawC/sKz7KFI8hfEf07qI7LgP3/lYFUWuByP02SdAzKHk4yg
YiXjNucdgdFdXGzGFH5kOsitMykhU4VPdPAmpRuBcuM/wdhgx9rs3V2rfPIUvIYO
hC6oIeh9jUPu8vZdtNVPVMgCw1YWezPbNs4wBfLv3IMVMey2S4CCwDsA/CNGG/0O
ebcReHhN61W5p9IaiELThCDXD+2JFL7hT3+iBj7dcVA/wb+DKVM2/eIFKz/aZStO
CHg69y0sq+Eh4/L/YEgDukRq/GXJs0WVuvxfwz2m1dXyIA/LD9GqE9r+jxOwlqtH
PgKA+0xFEM7pNHcRMfbuZe65t643vnegSjRerG9qmuock4ytbF8LpcvJg6fl+3jF
WRGtuvEVfAu/JoAR3uoFfGHOFhHm7h30cs0BWONEzFbJGL2EPALNefY5zbOnLBBN
OJ6HvFyr8EguBkx281zniWpsWNfFiOPw4MgKqewpPxJ5nLqg40Sqrz+9XR7/pfAY
OXIWI6RmCpPF6syJmu/3X+3UiwBbkwymJXbc9A0v2fEImN8Qp/QWxEMZ38dJhidn
NEDuzFMk+AG104zqetzo4biueiNTcflCXTXBhOsa5t7qk1MNJIMjrRks0DL3/Im/
tRwYmKRZ6fAgInDSO93G6+12ZRszD8pwCdm2eJHNhlLMpLt7gdnN1z19v1F1mQMd
us39ZEyWogoIc1+d6n43fRHQTvaipklsCD3e72kyUWMeJRNjuvCjSosF6kzLKFOk
O3rTQiaxUlepBG9WeFtPbnPXUmPhLG5ynFJz2JqG8UuaXV8+Q2PpzJbUB7OPghaI
He+MZ9QEQgNp6szS8uZwbRy8q79E4nVAoqqOximdCS0f3RmnK2x/CeAgDZbJ4HRR
1abp2tOGt6xGqwe23ZioeObuucZS1dgfm7+143cSYjbOGlq3yncPPvx8JKD8ATbw
NS8tV4qRsAr0Zf+MQNlgsqpdnC/+0eDMUXl3T3D8i171t2dnt5oYidFbOeYiYk4l
J0xqoMS04BSkHc3fCub+pW64Anons/rbTvBPstCBjhAF5/exFczs8u6PEqKB1Nyb
EN+AP5f5Ig512GIwzqVUvn3i/NphSNV9utgqogCMuV7A1AXF+qqhZu+Vzz8Y/rfC
2ssDVQWEYj+slFvxTqM6Z59JreGUUF8eQr5drlFrpKPA+feywYe7F/EmgWtwU7N3
JIO3x3n6JwchzOuJNG1NPKj/bmwbrNl+Z8wexQjFUHmE6ymdS/XMgY5ywJSWiIcf
JUvH7ip62mdLQQmh9fNa0vMjjFLAohXknclwqbqLCOyo44h6nBmgUMSUGEnt+vei
FxXpKfHdbvd4re1tJ9X4ElL7FZHIEDbVHATzjBw0TamwBjdYCaz2BINSIZzGm1Gy
LVBorO4ouyW/B4blOJrx05egfWrpf3RjCLY51P5vg9Sg2SF5FVxAmS73XRcxPyVQ
5XBkydNL7weX2GYDv5ebpd5vdWTaCpqah3zE9lQgZjhRdWC5CZaHUmk/U5PipX4k
0yC9P6xyeCOB0uvu5ue7J2U9StMeBCrvpKxkGBDiTpk4NvS2WNkhcygNFo8O8FrJ
rV3sZAUCNzQTu5oEvLThjDLSZEJToQW/611fOgPPhHwQkFEjF5hx71uD2Oq6pDUN
TLjEF9HaFbJrsQC9zouDaCGghNcsbEqp/U76mnMIIy5z310L6bHBiOMBDhXMgLCI
b826qHO+dOixKhb1lz6WYNj9YJnpdu1LXvnYcEf9LYpT0czybc3PA4QUv8LI7QM0
7uHVt+oK0csTPPHB2Ovjs/O2YRvZcOocgs90mjDX2McaqUwO6ZGprYrjwDRTSnJp
HkkoRhC2pzUm5j8v8oBQkkYPQXcbEK6MwF2xAqwJtJr+l9WASIS4+WHmcAuk8CE0
/5/3zNq8QyZWGkAGd5RsvhGMWsP2sBnP6ZuYfXzbrs9w5cFzJkEa8ApUST3jqOJO
Y6msYr/rRuhGAttb7L4o2jTUtemaDVfd0KdgO0sl+OX+XUI7Gx8x5frU9B1sEkJR
djkh3eSmglTFlrl4w8Q7vbEiDcIQiDDGVVT/9Si0y0MoX13+/CizAMFBh5aHDpFX
iQMXifp8d6wiakGkX+0ZuWHWgg1C7GhvGQeFO/F/9uXyto4uJyBm7B8dqtFRGaGa
oSc1TPnu5x4fdfOvApllGkKCmoq295GHOWuk/Hib+rPRq5CJhgSweKURc2/DDtrQ
JtSsxmNNHoM+Fr3vYT9uTOH+W+dT3mbECJwwYmfUJea6rvV6gq4bJm26bs3+35Zh
4iUZtYfPQXDM1AfOrAuYcR8dsw6Li9oXiz6kvCOv20F8bgu9mzMaqMrYtv9MdEW8
j0eZ6ksNUKFv644za09U4kYxi/BwgO69YcFWDGDVckTXszbKNInYJ7rkF6F0UXnO
ZIN7S87KS3UNzYozMswa4CAAtnqbNMQmRBv7R4tItcL8dHHvJPonKtnBZyUNQqkh
GMpyLAbEMo+LUb9nedOD4VOfG9zdR3TO8jFaeREpHxM2Z0nhK4VqE+Cqx1m8z/K4
Z2rtZ+KgWqWHi4G68Nn1iiKn4YEknJOA0Ir2TPIluHzvFXMnShWd2i9YnGCWGj/o
K26+cHB5PDM21szFdRxTtsLVXtWQ16WIR41qh8sg8rCt4+hbVNjUW351wI6EMTXU
neq8KMTq7Vp2jK/j74dU9gFJACzqaDyESiHFFB+bF4F5HJLJhLSxmVSWEZ8Gln6S
DGH3FSY1cBEdSKFQz2MlTCPQ+g0fatPLq70aD3nGv3UEBFxpoywuqGUu5D/F3GvS
EdRdQxzPEz3YSMJoqVu2gjyVY/W7wjP8bU1VN8FTW59AqSi8xAGCAthdBgEy8dha
pO247m47zIJdpjKqjH9ZeeSz/oF8eZb+jZPWDvKzWwKpUjzDkNthPl9vl8Oh/Kur
b0ZnJT1H9KAcqQntjUDKRB4DaHQ+mxM/iknuBt5XsPsesgPiesH3LdsfgnkUUCY2
rFp1pmzRnFa7dqFaK35PHFk27bGTsdTRUJFrN0c1G/L3OHk9w/sJVwg/jXMGTS9/
GU9qXxihbbTPsgqVtpuaH3PoIYyJ9zgXhcPRRQdQjg9fZhuuo2pmMlENzuk41Gn+
u9QDGKbTt91QMimzM1M1LZ7z2W4wz3wddkYh9ym1KyyCsY2nxnprt8ASA4PeCR7v
R0LWuwqiIir35e7l0DXzipIVuvt8gwkwWAbfiFahTjBWlNEP7oeJkX21HyrpUHg9
uqR5KMwjv/1WuL9WbaFEmBPFeygmRErXhAz2Nl5L7CEaNFZxNKn+dHS3aaOePK7x
g5OFXkseuV4nItpr0sg1EjIVBXM8HKNo3fquX5ANy6YszZxOMpuFa2XY5aQGC2NQ
TCbYvQCcJDtvOSvcRco4tQ/bZiheM/F+iAkU0TN3UFRa9hlYNTwZHnEOmZimYgPW
9wYdrCjcaR0AyLL9J+YX3isKf2+7+BANRwp7ZpJtpOVD/5WOWKqVfsEYifrEq3nd
nqtBNpTlGTYd1z91E60iK/rh38qwNxZ0YECwWrFhZ84sJEguw7xIEsWXrrmTPQuJ
o0WBLqxE4bmydK3lt0lZc7e6/+3qBSBtY5ZoSRAGD7a0+tbNTaXA3bN2mPfH+Y7g
QPLDZRdz6waobOmH6gKs44agqWCIJb7obAYhobpSBfFmzAztwQxa7f2vFeL0mO5l
AQA3ARSzqh40ocDXiM2ENYhSDPKL4nwayEbb2wHdSZ2VWeTyvmNE3hNruEaf6yWh
j+GksAKDC162fBwkRcX4Gr9BXQkAEOBcnBjvU3Q6ujdPfTJEVwc9ZbJXid11P2SC
40JZKrEbHvJFKoRlrdSuAkUcKNdeSoio5GItqYq23bAqiuLg008Y+q3HrNnBnbYC
z72SjxXx9vn4/+Z7z6JkMZSRWVmz6UoUMpLU62sRhfAzDjz031HjRUYwGQk1kvYM
aqhEBUokCuUaRNhNULIAiTEl6cf3Cy88+zXfG12+T7L9d7wIrsOHzaWw++FESKxG
PZg5CxwyrveSLDVACg5R5ZiuOIBWeOl6BUgPUgg1juuLVaft6csc4tKjEjcjKXFJ
9Lm/n37C0RH9/qgptx2n6DEW8C6xCvf00T7TGWP5ictr7CCw8qF+a1qBN32jvktR
wQSO73wuL9UYe1xZK5vcNv9NY5H3/j/WI8e/cUFcaQU3taCvOqCp62c7VYnrMb4P
fRE+dp3GdSZpYVdwE5KE0mCYCNMpxefHx0Q7yft31dRegvK4xxqZnZnW2I0k6Oz3
ikByg21ZOn9YLkQSVO8dqUnP+HCuR/sVmQv4F8tjHwYR/szyWYyxR/mnpp4ptM/Q
OyhsBtcayD/bo3abLpkSo5dPyyOawGjEeilb+Rg+RHKpsmaZ9aU7vcYegGtOnalS
nVJaQK2356fRgqrC//uCh8hO3YG/A58IgW2kSAYoQbxD1y/RvXUI8w+UCg9REkwl
9wL4RUwIii76Y/fF6oJn+SmkLQdlzu5YfHwnfutlPzE5PQUImxM14h7wteReV0U4
cMaXwO3DbxGvgy2L3uJYNL9pp2FduCGXwDAvOZPQ5CuLIGLFWSwerWOlcfzL3tA+
ynsLOybYrRBUBtFIjoIRCMVqEenHrZ8DZc1nMCKpgWrzi/L8ypD2lD/dwFCwq5a2
qTh5i8pTajt4GMJ0YwOamdRjogGsxzRy8VTiH8hlZur9tcM9LMypJ0Y1hqKmvZv0
PtSoppeXoAA3dnj5ZNXFPdgz355STamWiEBKn2lfaTPcE04wQwDy3JSRAbUsEEoz
G8Wi2hA+qYkRuiq7wiLtmRYdPkliSfj8aBoT7goAQc26O9/a22ucnteibk0n42nw
+JvW+GtgrFZ34gxxL874NRc/uIywTS6oWf25HiCQoUAQYc2A7FyDeDJqZ1KziqCq
A8dxkInXe30XstMIqygSL47+VnVcc2aIwSOjE5n0vMe+Sgss5XDqki9eGvrpmjwP
7B44DbAnbAfQfEVJZ8pe28VIfs8pNE1406OHaUmHPalAaeYKZV4Gp8ETCRJxquRT
X67G7qu8JkE2yo8Id6som0UHIS1nssRR4EKw4+OLfuTE2ZzH8Dx6yvhWSnHv0j0h
DNRIZ2Tz0WNSU5pLMKWY0JKDS/p76TtKMgKpkAq03lfS4qBPIJQIfoZeEIsmQn5T
PrBjH5o6cB583X5aTOpIl9/pQJCOo/Hzdu5tp8d0q8K5TadqjhGDoPCcSGPcrvRt
3VlbWaGRIgve5gsb98Fol3/icw2iHWZ/XwIKBdupnvtaR+61i+B4feEaHeOoo7TA
8DYThXsCBvpqhGirhy4zjzsSM9nH7INl+7vUP1skodKzfwP4XhEm9O4GEI3BokIT
9d9vRQTE/UWHddAgc494WAFdphCJORwhUFAWMwnqXGbIBjMDyt/vvhbaAaNUv1Gt
4OVB8/aCG3AbsgJRRN6LhwJOsKuhTOJJPiZDG7SULywNpQzmRPhVH7fHDHMZ+EvD
WMautgaSXpBjio8Ui+Lykhm3EGlmdX2HodeMS+ZpTFGqAyz1XS3EDuY61nZ+B7aa
U8jWBPuMZFgqzSSqK/zni2WDc+jZ6dvyDRGKxl8Ebwtsfj1+l1iXZx/6LKxt45Bc
roMVwUSv4uu+atYRPus/2LWg8OL3ZDX/6b+it1Yxg6NVph6vO1NJOQc/18WJODkP
cEUw3PK1e5VEq9fz4+pirPiba0imkJxwptB/aK5RKVsHq6TfRlbX21vK6f8WGbvY
pZJF8s90YE/WuEwKwiQVYGfscTsiR8aphiVQBnZAMbKRpu4Y/3fnIuh5f2slk6i9
GOkliyFAtrJ1ZM2AUF4GZgj/3fj6BadBeOSCideB2e/6zXjUdyvNMRCTPCqr8usT
7veVi5ZypI2oN7IHITDR20CXSkcpxs3dsy5jfYZAPZcye0EkuyR5NuoGvXpS29Jo
EZECWN/1OQg1Xv3+jZXnbxo80HBVP7JgOqulpFnr4zPH0jn90+JC7E4rZ3elTsQe
M4m+WHwhkZ/ye8CCNV1YUm08O7RSEeeCRR9m4CKSPUIhDo7a2kx8Umq0NY2vphFN
nSMGUXyINnjQtcql/kOBrB1LOQTbH38x7nUCPjPQa9gms/0BL7oWaZ2YxY6fDFT2
/jiZ3c3TWapU6FnjVl6lLyR8KU3gO4v5AiS04v84Gv/o6r70XCRTs4PnAh3iJTgT
Pm4KzKYcWe7cFLkM2tQsioRqd4N966iU+Ae2jtXGv5LLsxjV5ziv7urQLOntNRvR
zAyrxMq+mn0FmYwpoQwTy0BZxMPBUKqEG7YJCLvz5gH8kBBUjaunPQff36HWhZ4O
QDV0CJ7K8sr2zUnDb04d8SYeBUuYjPSXBr8/wOnBfMIwv+60duiI+aW1fgx89wxl
6Rz3lKoBZUfYXIbfOLTLyf4JZXnD8xwv7XeoXbvjLYc49S3K37R4/0VZrSwINnf4
ICL4StPLk0EtPYHclH0U9JJR5EuflbbK1BPDYW9+i+ySSKB9qg/yxwrFhI6dIKZF
8o2yPIdXqzgjO3jSZ10tZFktVl74kUwQhvwSZFTzmIIz0/yZF13hcU3lQ5MHv2tk
NOu9bNxhIjSaKm5f9MxpSmpUd6QBYe0Xk+Fb1ejfzHOMD4eajsnjptZy0y93fB6W
WVG+2ZGGX8AAajb0blb0wmbJV74dbFIRBW/O+Eg4zwgikSgdPoDxx8nLC5Xb0bMO
X5hm45EY1JAGAMAqAszT7yZ8r1BjiVxWHMrzEkjT4W8OP7Fi/OP0I7ckN9LOyIX0
DqrDKXslkfjy7z9awrg5JXSaEAh2E5zzP4kUBssQMyNSaaGe0R9m+CpO9O7AHaXz
wcNs18uiCGGWj+0YoO+xlyeWvFofjp2RfiRVrWmF7i867k0y1TuhffZd3alS2Xn2
uuz8q+e4G92yJFr7nMw9nLX8sxsFMN/Y7FzOPLT86Zswmf8G/eCUSTs0QHapPnfw
GiNp2nJuM9LrmvrtrkfSScA/QHN9SCPqp+kPzuIfXht6+Q+iOS3Cv0Fvx70izyDK
33VFsQQbihtuUcEX1eE17Gv+wYS8EoEClevbQGf3MKhaHkHyAlxjAOTf74c9P71M
09dUqzHhK3cxCiaEXQdyNXHNN2Qtjzagz4M1D/xew0UVzIF101yFiITlAPOaEpxP
5ube/avHacAfXuUVo/10wwdeo/+u1EZlEtlxbMc3tM5pV4am9mjWb3XC/YoG888G
44vCXuvR7Fa4QWNcmZlzFShxgDP8zBqqf7qk/aWSv2mz3KGI2e4VjuJkHD8TPgD2
5eSFmy4acz7MSD2HgDVZr/6L2pWuNZqFc7uj20lDsfwv7qvq9wRpnL0NkM/qHhGn
AO5VhWAuQ9lu4FMrdFCJYzn5uUBrUoJ5vMGsFMkkdPWe4zBbOPUeaOh1JlYaYQs7
EldH3OpUqTA35zdO8g5roGmgHJLv4wPwfgholfTJDgvNliO7WrDCaNOoLHv47PNW
wGjATkTAjGyQS8A/q3spWEZiwu12cK/g+TzxSAaak2GN6GSW31b6LsKBXArlSW/7
rsRxEl+KMiz8kBDiAavztAQpK5FDZBcqGI4+UuBVl4NmutbdJo53BXcHDRU4ppwh
tcPEvt2Aj1FG92Pl4aq60llPu9bGd3Zqo95Hwnm0R6MnWevQzY8wun5NXhk8Nv9b
tHqRTXqr21Qu4YZQ2/t/hWN1ApYmsa5kAhaJJVqKISqR/BIKE5tEkkzVoytTe7cS
JKB+ZcVQJ5cn1CdF/ffw7uLlymfZ+d5ezhPgnB+EeJNYpalkNxEwYoTdgJwMYao9
4BnptMdKhQCqkq04pLZoyYcRg5l+oQNSO+3WhrYYwmrUjgGzw1oy/4P1VKRMzKhV
RURR1u7ATKfsGRIVIIgIlY8bUEkdRf8GcPMVL9OmMS+ciMziPwot77BLE3tijtRJ
T2aoRIRq3/3yFMJA5w94lsoeINvGWzLBs/kW5Gi+AA4X3pmiH9ALxL0j0H5XZ1r+
de41I3dlGDvgRgbBKz+9pTJSPx6mTHaYRQr1ZaN9jTPMyuULQ7dyrYJ8BQC+UeqL
Ob1tCRxo3ZodIiQoREPF8XbKaSzjKcyCiHOmJBcKpiy8fyVyf/cVFKW8VW8jJWym
EOqFlmk5DT5Zl8poqVzahmobgg9oqDhtQ9l9IJe67pd67owMPESqSk0cPQkmcdrA
r1+iC/YsFESWj2BBlE5mKj6+P7lFH3M/lrv+rI6srcz6wHDRhLiLz1JNKuTNXULa
MffAuhLdyidx+f3lSQCyyKtoroAHeP7XcwWF17s24BQxvRZdKyZhAVX//zDOJtDk
pZY6Rcqp1K6rO6Ri++DQuvAecuG9LcVmEh5iU2YhWt1HwRuFKs/z6iPRTYAS6WWU
XJOzBVS2QSC5Fe9YzWTbDCxoOFEMoGWkkT3VQdrA2O8rcR8nByRSwcN4kytj/iny
TfOcY/+LkkVSAZ87XuRRQtVlWbqgOvzGJ9DOngpRp1A08C4GgsU/jKwYuRAqeDnJ
rblW8vNS1x1uSMfuKC1gm89OVpiMCabO1jl8PxmJigO50hvIUdmrUCpR4Rc97vhh
1RM1mPwdbxTHn8UTOL3O8hWxTKPZ37DLPJw+aIKFrzN5fqk/+LH4OOFGClOZ2XHA
pyAOUHFUOZjmfO6N5D/Z4WP7f0X2YoT3diDQEwdJHN8N88T/EcBfJsW6VW4s43YS
N0P+cqOBDYU/ZMyMapwNEMVBq9pgxrGO9qgAEbbmA5SLXpEHDgOp+MI/7uPaoZ/K
CZNEQIW0vzDFHNCfW0DX8La+n8JgKggzdhT6Vs+bZ5seNNGvETF0n4vIVPty4vD6
OGcOQDzKquM/dAmN9JTQjspxsjQgrfprNNZVsO/Rw+Q/RAQWmP0Ud+gDzfrkXukH
ppzeNZ14NpceXBBcONOztp3jNb0ArZsjPq2RnzaLq1snqRbyf8+0WQjgd+o1WVE7
j6ZXbda/eV2v0cVahHtreuUoFfJEAPvJwFWER4Ahd/qSpIj/KzlO4Uga6w7N84rl
znMP372V6Ft/PA+fb/AXFMUjAQbu6/yuGEaNdh0A/lweymwwkCSpMza4YiwUOian
ZPI+SCm5fuZ+SYquCLYWNcZrLGU9bGvTIwJrPZmU1BPXof7RH64Rz5Fe3bjAPAxy
7n6LYilvPIOxTHQZAPSaUHgnaF4BI1qymqMZMZHv2qOvS0WjVEhDOO92SWfYOEqi
Q0rzhctL1HkMNj6YoIHtaZ/oT1WiGWt7p+NhVlPF8Xh5KsJJ9uEFn4MV6oV2HG5G
D8t5mDCGNuCP3NY89qhZFuGwd/ioC6+aTmkJH1gNfXaY3FtxfAGOuwAhfK6HsFY4
o/2vLphQjyWCRueStQSBv8n2s5Mdu1EMNy/xzB/kBd43h0cQS34zlRFi1SmUFax+
/+G3sXPimdQ46gvV1p/QzAn3BplkwO1O3DU8m5wkPUNC0uFtvdLTF1TBWF8ZIola
t+QGE2xfAw8+g08tLfS0Sv+E5PjgmpepQIu9Pz29LVdRB7EFgVTJBrNiF0yF60KB
wg2k9Domt3Rxo+R5azjzPH0s3SMS6J7eCLFoNhfrZsT0ECKXQGAFMNcQhVpdT3Ap
aJx+mBGQieze7jW4tMLQo+h3W/X2YmT4NjXW646PhOHPKlHxDUxiZZtVMre76Fpa
EZagJVXcCpo2uC3qaIK5gUQ1BpTY6JV1srLzl3JIGgtVfO1XxkddAQlAztlAOz1K
SU4ormqFIVVxOYI+UF1OGnmfUu3Mz85OkoPA9NCkQs5gev0DrDcYiNKFE4DSPK8u
nj5UraYKo2p76UAmeUW6nX8KMWiEC4p4/lxJU8zc1O3TPw8KFVO6igUXmwGvz4bM
gEu+cDhBizYrXRkkXm2enpYNOK6TO1tvG7yFxSK4/OATb4m/59igMveAGFKC9835
OsgwB5SlOa70qtxcrGH9Fl00Bo665YpPNHD9KHT+fuXMkMUve9Xq14KmvooLY+Qu
XhRUynpTSKTYQQYcmpLO89iR0oVqS8/bNgbdg/g4W5Gps2q/BrgakfygAHWUmn5A
+uwro+dl0LU0fPkD+lc+N6uI7DRm2jYR5UyRMB5xijSVOUzvmud5lgkL5tfrnJrL
cRhbA90wJL083DH5fysfaJ2lepPSIxUrdrdangafNDdY25vZCxoPGmDleCo+UVWe
3l5D7hbEd9GCCyu/Bf7bs8iW+IlkAVVgk8WJ2HDbhmYILJ5u4IElnE6sqb510d6H
PxaCw2vyCXtd/JCEgIYeueuNKoGzBQt88gfRDIVIBcFe7CR5NxMFVLuQ/ceM8rk4
zqXr+cLb3prHZQ02oCod0LW8ZEkyF6iI/PMucMKHDpGsdxnxVRdHw4RlBKinmBPP
QpMrXKpznjhZLQYc8eXgW2m3MnV30YUEAQ3+xNYBqbwLQ+3pJNomDcfNj+Ndf7B/
DLOinhYo/+P+bvdknGHO+2ZX2kSf9JOL8FUXXgrQeNLy22iDdlei0mXUgb/sz52v
wBDjqzA8uVpQOmy6NZQgsbKoxs1LBw0XKtlXQxd3HaeCj52awI0ABp/saEqyvcuz
wLB0jokxL2k433QRWzoc43qIZr8UNvO80CAvqqSorD+rmoC1shudZrD2Ztu+V8Gb
T2u4VQGFrXuaOuVaSynTyM2B27izRFQCFYzH6dYH8YmXi5pL4tG2GHSINocJes+B
4P284fSyatrcfQ+iBW9fJxR2S9u7i1fsiJNcJRFIr+UEw6a2AfZYShW3EOZNhHnj
T6Ks7RvpuISCIq0t4t9mJdvelk1y/EDyM0DFtAflp5U7KYMOM35cLXdW89O0hB+Y
y4qQhVmQLYFydwXMYwgVWXVnmhwgisKJ3FNsFiIBfkTeewQr2swv9Qv9v9CKTE4L
6cs69TTPMkA/2zGSQ/+SPMpAKtuJrea5vDiGPk/4QvE2UXvGNoDt+ACXaWZqzTuq
sfnwMdA9OkXhlfobZ6HsBFM21P9xXjjoWV4v8TCz4PCtkCcNUvtPE8gTOwH9y72D
BbXKS91NFtrwhaxKjIaVL/7GI2kjsPNLPleSfSkzTvAIeEm8u3MtEC9Wr4zbnGF0
xXo4b7pWPlaoKiGLM6bsQBmrtW8BMyRo3zlDjsWnJC32zHrszCgluwk+ftX061ch
K2YY954rAnDJmRRMZD1Hs4kbi/b+nmpwvM8xH9IFNLJ1brErFDRR/Jt8ORRSItCb
Jyxxr4C0JIPsmtJse5915aoQ37vc9U9msE77vTk4g5xiTN5zSLK24PUvIjtbRjkG
BVxCQG0aCt/DhwBhS1mVUjJpSQhCqWbCAL0eeT4xlKq+99McYqp5Biz2oZGLZyuG
FWhoEJgb68kGGjajAQP65jNwtx8oOT71V8NM2u67cUrGP4sTRc1+BtqkOzTK5AxE
7qqq6ceNDzIUEtqav58qjOzbtDj88lnWm97KSxpZJepTMTB1HcTggLrRcGG/KEoR
Sk9dY1t4ClpPm0JFtXE9GgGFtOZktduObX+Z0SDFTHyymBkj6QuYWBLGg+wIYIuQ
ninsAxvyLsQb7MC+Qu3q41ShEh3QLn8Qe4lIWs4YpfstYzxysLq/XZQbfRQM2Slc
G9cn2fnOi0YoZxjtYWrJGj43/E7mP10OiiV1yLqIdKecdAJCJycLfa2StNn1K2hC
vbW6wPzyiiDuUrAjHIGhjYdOdp9x+HEBsir77gfD0to2YQc2cYhaJlJLwFyJbJK+
btgZgkXqVm6adBYZfZ3Mu8nRSP35/oZ4SpafnFD49fYfrJWUS8JXgUVlzkC04OGK
QiJNoVwUv+6jIZZEbykJbYbZ0OmJo/I4iYwHgWeCqFGXnCk4hjB1ILj6Ohm4aDqR
SuhEsprCGxVawtH6VcH+vym9nh4m9klPyEoZjtyWiKn4Ji7ZWev44MwbvdPG2nic
JB6uB2JeuDTs5AxtjaTGBd73Q/+LJDocgJPWNDFLQyAbG2ICfDVxgiYaHbP3sCOL
gBB7ecAAdRtfIXcsB1IXilPABe2Sjf9ymzmzcH/SlA3bA/vjK7L+NiACn3Vd6Kie
+a6evpLPmgHA6sskK1h2MpwFxT3rzptBpwHHJDeaECIvE+44I3x8tueEwa+9XGN7
s3HZCDK8uYxUrMSpqx6z7H8BxvBH09FkO4CFKlp3qb0+5WsFtxB7/T3F+areU5uc
b2X/mr6ZsBv4Kfpq50y8Fh1iJ7F6jWzF4yz8eRR8lfsAYKiE7jL2EUYnN+EWZDVL
M2xLddc2ptL3yBWrQTPv9ZK1jFaW6PONclwZzHxQw7kygbhReYH6hpwpm6+9Pe/Y
kaQFi6hOCmsdWi3NT/2fez8UU13TvDFky9YQk6kvhWsbh/0jrtWBki09Bcejnnwq
pqx1dW6QBtAIjICwKENOdpHYq6BWpr4TEZznbXJnvJ25JASgX4CAFZeNX41qV8Yu
5VkR8mqiHGHODAr0DqklDu24CdUC/rKvZ5BnRCw+NB4MP3Yjo4OpO8q9JOHIt/Lh
9dRnpQAs9kCgFoXcXq9hzJ8dC7yu/xvTAmLlN0wEQSzjqxyRZ8w22bEOidKGP0FC
Vrmha0T10auj7rs+w3RnHaiNqqzohIbGXpwUaJV3aCZu5LaIvOaxV70gEeYE1jvN
vAuyhssGA9rn41kdfFMyMDy30Wz61FxKAUc/oecUY8Cb1kD8+HlKyhHNG1AETus0
QjVzOoISCZPcVkA89sxODBUKEH03lnGhGxQIOPppV64F2gCzHuq3eEJGUUD/ZO10
1AxU90gFC/PDYoHzD6dIpv6UPK8+I7lVWUUkSObo1Ak2SgYRj1pbdA3kfGRza5pP
/WeRpBHKX1nLuLCbmq0VXzLU0BfCpnovGBv1AN1w5bpWK+toJ7bkXmK5Xy507y/1
2vLbT4oIcpLpzCcaC4viqcHffE5uR2Ygo8dNP5jgOD3DBwvy4yftlTQEJKZ/H3xI
urK2XyN9+r4zsa9vHn5lfy6cQv7P0biahHqdxqlqKoDK5fWUNN8y166kNrQ16KSV
t2R8HS039D5QtuYCdLZdBjF8RzQ7kRyZ6AU7EWJC7gXoVMu8ynDM6vRoCBYcIn4g
AwBH9zct8Tq31KOKXY8aoy5PKcFZBoZrvSBxHbucAFKLPxyRXKgB/8YwiZqL6Njs
1kRAhGbcS3ZnKyOvsbviaPAXU69/An/xkyAgR1aHzZCfkB+nPXPO84+jh+rd5kGh
H4sYM6PeTX2FL7xECy1/sl49gJhJXRoHPInxWP2Q+T94plhpWEQQ0l6reKUi4rX3
rDp41ch0BlFl+lnu1ootSlQ2CD4FjIlm+2GGfvH1gCS/dcPaMgRuby9sTNUNRGfh
4rxqawNQNjVeGpkFZmhss14/q2od3Z6rewgPFeGsX7VPaf14dEtjEcRo6XnsG2XZ
43tjGs8MqSqrxjNeFtmSZb/5cQ4llSBiC8YdYJBszZpg/9yB/BisL4dKqzDH0Cx8
sUzS/fbRVBXElsYtUajMC+1r3GiiVYqJwtVMZiJmsdWJygcu2otPwtbiFYf/kUAf
3VI+nfTLe5IGjreuRonNxyvZL8bzHgPVTItrmqm8JKQ83Mxqj0F5vuDR8EUMbE5a
SLpTrSU0aVyQAdoF2N0pqmVENY6kGuSxeiMstmBZrtctq3DwC8OVppZlxElVDcHS
ZYSvLNlfJygbU5LHMvJR6I01w0MkNERQ0Rd1DHYsj636ud3HNY85O/htYXgaE1nb
ffCk4KBTTjhbrF5nfeXlPL94KyTK7EnmLfhrZ762SCM1T4QRPDeOUdF4eaJQ95lC
KUnr+ga3SZtcnwBmCRYaeiYO2ohFmylL3IZIddFAIMBswFtUhVdHkKy71DwqNAkj
8fKklZQYTv0kZpn5/0kKCX8L3zHtk7NycxwngqbY4lZbg2Msj8kvOHqbfbiksNyC
BypRqQ9qxjz6lzMl+J5oSlQtk+Stwgv7TD3yFRsITTeGcpGHzI/wwBewvTXuJfsy
sItuliW3DFwi2ZRygsglCQr+XqwYUONd8qdI2f0cR7byFKw9QeHLnOIj42F9McwV
8xJbO66lMS2NX02OWopskza2R+z3oeAtsRKlx47mFCxYcmzWDbKhKAIky7QJGxOV
zv/7zBd4eHngmMxAG2WA8ST78NcsCAbYAJIN4ufW+U6/FhMc/4RUiwzakAZ0UwlH
NSyPJzGVHIaK6y1B+3d192RBWOTVLkfIwUj7IX4WpRQj/gpuZSxxXLLxdIpCxs+z
nZardTlnQI+POpAeqKODmgnDcYBQ1W2YkVBodD09daytqsomnVkG1RywHdbfcFV0
vd3chpeEBwOU66CCe0i/eIGj+G6aNv2P2iTEpxxfBU66oluW4ff7HsZOs/fKGXWt
9cq/ty3w38UZ2zGYx90bgCkMrEyRHNeM8B5YDRUa79UJ59/yFr3X79R0eweU4JOY
kR1sS/MzCat7ktgChdFVLj1KFlEZbBIVwYfezlRsR1gc5B4JybiNWJD8eGETyX+F
FumzIyDzjydPGhSyEmds943eykq+9KneWxJciQ7cIP7He6q4gNDO6PJWsQysHJKL
ixgCI1ojfmWzaTgc5ssmFbaqt2oZNdClls5EuZjPNI30IXeX4GKgAYJ3p1pTCzOj
2uX90cQF03AcRLOSirSWSyFMiqy8APpsOeEfkZ35aP+boTFAQXV9fHTLX+KVF2z1
X+nZFSORY48v9pi8CZ+LWDlBAkvdAGvYDhlTNHb74BrAd+fRTdiY88HUEK7U0GPL
etPxNAMPjvcgTMyIPSw7yQ7I/d6xdH+fAlyA4IJ0Q9QQ7Skf+X5vo2Ub24Tg5ujN
iukIGTjTPmxw+RrTOR7AnkIk/hJutpc1y1DMdepctXMuzssPeC7aPs0w7qv60uEQ
zpVKdaCMSSRL/0v90iuKt6rzrkv/GwDn/fM2MFK62GBLleGjuK+TQV1ePZ/f2iQV
iqdSf7ClgUqqPBnNetAz9yaukacGe1ckjK9lOlxDxsj4wzjfZ/qfcWNGTA7jw/nl
ehYSdufzRZY2yl4f517M/PDT8vFIUtJW7YXO3Pq/LaZKErzm8cswpMeOqCQsqcfR
yfsXEIHFxpXf9N8RjEU60PEOPfzn0wsijDjbVhZQcb6k25ESAmCp5/Wu3n6iId4n
PpZcU+hWlkTlV0HFP3rNrGMQag5XINSQDVYjhS4uNH/YJgoRS4pefaOqn8Zlj3tV
s8mnQAOmqgaZAZiAmCuZFlUywUHee16VWur528zYptiMmszKcAeJgKEC3v+/i1ym
Vz1KUFKxQRlL+NaxxCZRXkYgGniDzBeXteaYRkY8j6kR/wHGO8uQE7bRIOG+0D7f
Fx6wh89wQLZt5Bz8a+SllZQzVZ/VoInqGyvLfb8MfiNsx9qld3bJ4RRX6D18wkRH
IgUV0S5qRWr6SyDRevI5i5tNZOcRk09I56NtuL5rqnJ/lodSirFe00GGmBASCW6m
FewZJ0yKi2BCkhlN36lKoFLoxNkZqG3j1BAomUXTIvBtfTW/yUs+S/fbFFWvSWTj
lNuhmqPaDoDgyIix3IGqYTHXiVpGYoyjczQy3g4YZZzGZSjQWXeyBD7xnGWgzWpZ
EMyjFnNs2a8dlvgekzhHI2hQnBR6kuQ6d420qqmwZ8m83CYcsqGNSehq+n/3hgLn
7nrdGC0gLKz1rtjKPbpKwIxkQuR+kjbTsOHysCI2XWoeXMIHT7/Rl7XYXpdgOuTH
3EOo1t9JHle0HH3xgoN9/qzQq8mwmCWbQz1TODm3kxNS/BvZbMyLKh313wMc3pEO
wMG5ZpzArWnIf9wlF8TdtXFZlRnxeZ+7eS+vM4zfhRhxz8qR/lqLKRDkeLfWPrPT
kUCtjYwhoO9BpFUBVCHlfsi5iF/lej4FXvuj+ty1h07ZhspyazuW2726y2gb00wf
L5jLfkQNDyr+kWE7lJ0mI9gzIAzRfm8O0b9gzALWqFIfRv8fK6EnNvAaHHSun/ap
HFjMFIg+6Z+BhLMcZtodUURM/hm4Pq8YFkqmkiGcaAJnc7BppQ/oMh1G4ztdJWpu
OEiPH73u4gH1/fVPgSowmdm9Rb2xrvP2nAh0Ee6WPAm2Hs64N+XDAKkXog34nJDF
nVkB7Yyns1lbXXSdRAQSLLFemrtlYUrky6x7hGA5OghfZM868iMo5pMy/OQL0si8
FeQvwcj13VDJC3hjpeXRDGZQvWG0ijdbAvXadEbTGXnmbR8fSFNCjSTl2leGpVne
Y5dn9HYYv2ZqA1GS9ILUvvOy9Py+fWSe+8jmsJBJNbMvDQV3g10yPdu4xsGeg839
Fm6FFMkEzq+B9ISYP57upQyhA9nvbh9xWMq6Ro7wiScSn5YfE7yRqPtLckjXUz2n
e7zIJkdlrDKgfU38IuF29S4LTHu+HK1IoP8e+wOSkibyrCuSWTP9Iqt7sWCkzSnE
dzMOsFsFof3VAIgL7AQEdOHO9CmbFPi/ywYrRRxwHbKWVpaD0GkSq7uBXHWD1PQ7
s0MFUwytD9e+AYcGdq/ljhcMrdISqIHqV8e7KyUaRmCOnG6KcDOwffsxtuDNBM4g
S08hVkrX6mn7eC4u6W1/7uF1+Piq5zHE3bLLDUN685eGPYyLrlZG3xRGEdoMe/Xm
fGsTxsQmVZx4oOyFKqRNEsYRjWnFdZMWZFp4hy24OPV14SF03w4IR40pA+Q5SvWD
0vdEqcCBOOlVlIxKfYGCdwM+WI+Vjdh3iK+VuPhJwTCyY8miYpeaTWL3lnZfMt+c
Wb/loYWrHK0dzjk7e46htq44covSnLqWB2HVGf455eWzIpHHTyyJ981WtXfLwcnb
898JIz4XSrX4xy6AidyXi6u+Y/WVDr2DJHo4RcNIv/bLlvgQE7q4fJc/OlfqdDBh
yDLgTnQLboa1iwNaGakAIVav6hdZCtYQfnGYMn9/AdkH/JQwUD57R8LxUfFuNgCV
NfcR6OmeF0EubmcoFpqPBu0VGuUmwM+b6poq5u20mK6K4/qFf6142WjQbUb/ww+T
elOdQ8fz9tNVVwbn4FT+4B1ejFMsL94oAmvmyP3PrCDRoSYy1Mac1zJdC/RMBebV
udesn9aSgopxhT4Z+qRsagJ75mHbnwx5e7KNMv9RzH9uXd+O23UmwD14PMgHgxBx
UcwPsdskloP4wTAe0oZwylKrwLwUW6qh846LXS3BzPI3vO3ZWhSf/5ZOkowzWpdd
0Fiy5FCWtLnn1N/ZRQ+7OppsJ6vVggLpoG0u+HFAgYMCc4SMQ6aOyB/aQgUQ5VJP
8R3E1JIKpzuQC0IRpVwtvUxqFTdVEoutWUDx55b59IT9/h6/9HHpAqOEXUX8Pm5x
I6MXDyRpvrJJTn3zQ8JpzzCa7HLn6DCgvsXfJrJ+MVt9vqi5QHdNC6Y/QMpagg9Y
7RiPZeZTvrfeY9mnNiF1fvArMy3jcvHIsaJGlHFun9Tbyut4VqSDZN+MG5KJVvRi
8SnRadJ6ZIjC2UVg0fumdKvr+FHbqutVUy5C2rwnVlJzsMgbkhXSTHKlxInAZGDP
6ey/fqGBnXjRlkPpqnx+ZTuNzuluRFO7kgVz8Z5D/2QPtHDJFDcToeLma8O8BzGe
h5ZY+dy32xmzMCf2PnYS3kIkMWSXolDs4AVHAEF76zPnB8VRtsRpyJpq4z6PYCQf
eaHyOOzT5REKNvo1JjrU7kvqqKYpVRaIhwgbqtYRuvEPyKLZkjFP3PoW4dkoTkzH
G5bokPgO/hLkaDR7aUMDRTvjwiSFYstdkZ5orbHPNirrQAAgIO4Gwb9QinDPxY62
DovYqUsQ/ffP70lDxSzeNxZ3mDqbLzTVUai5h1DXuoupoOIavBdbDEQOM4eCPwSx
Lbu/ST4+JCk2GSVOt5INacTooDs/3c4CoMq2fr0rnW/RKGjhVWjQMa1bRbqgK7+h
jzunTXd05LGFVfp5VQdRDDidfPKVfdg9jUsZlYLIbvWa96SCHKZ6nKvI0gn3eufe
09IBSPFZLSE0Hbh1nMbNOPwqUhK1mOJJOd+0RV1Xyxnb7f9gJKA7Mkw8OAgRKF5M
4e8JhE1bXLMDztzS09h8yLUSKlo7Hwtm0c8vFv6SV7EV0YMNnk4dfJDZQXR1YuhI
SKyRdTA3KXt8fk7rYJdrC2UnbwPO7WOlrhbEHwi0o15bHLyZc89ewonMTY0bYKxH
jWDjxno7fGWEIaTo8R1CZjcexBPsQ3vOAlBi6nXka2XU+LH9iCw0Nz/rVkX4ZIVT
2cCQzJLcMz4WFd85lz843zrut6wFepg19pgif/u/uJ0LzX++TRcVqIG3hg15E/4Z
mek4v4OVjMNtyyxUpiUUI38n34ZPAbtt3SdPX3iARxm8+JQlLP7pF7w+3GoupD/u
8u0TUw4a92c2wOiQokvI49lem86pO0pp2HEVf1OOveUiS0Xhs/kFBiTh0q8OH8z1
WKsdmBsSSZZkU8Sz/CPdSTmxN+8A7uNsh1GctYMioqBVMbTXB3sB0m22jhuVQjd7
4krVZCWAkO0YOfnaM2VVLeD/J1ZC20FvNQdo5GUPfF4e4zm0hpMkiGHzqK1IrPFV
E10PCezbz5/mJpD8L7A2WDcA2UZx6la66imZDiqz6Wr9dxiP6lYOHiZstT6JkCgu
yXUf/N8og20oAnd54ukdDNKjvWUiFZHnJJrXbFvcGlP/Sfvr27CRExpiFZAPQzHj
1C7xE5kfIU84nvWaJmCeucSX94JhBj2fJETnrjNy6OyL0yc1h2VQxp/hF/5QRhOm
07TCXwenayh8T5hlegiYlfaikoV9yiqNUZ+2B/q5H5ZvsmMDIw21qvt4TKRtitow
BVwa094hEsgquGpNwkLd6mN+EXcLDtdRJGKso6SoKzT6yV2QOIJyc5zWTj9y2USb
ONM5ihjb1kl7x5kKsoCTe6m8mZHTGUux9T0CRCnAL81R7mKD+axuB+EHRe3rjHN3
5bwE/OQomP/ptPvNhVEKMUB9ghiyJEF+kVkN5TqPro4RVrMobvhf5ZETlsGc0/XT
cNpiniMh1+rJ+Rf8+2STb+gRhHmqTfStkVNzwm0ZWl7wBLRNN67IjCA6ZkBozk0R
2FZ2/uh2QFNFn+fUwsijGle9rHAkYJgdQdDRSyxEB9+Ub+6EPXdBUVq6SQyB7vLx
ufPQC5M0a4kwksBLzP9VLPMtxcTJBAQptXJqybXFYBbdMbT5smE8xBx4NmvJm5BS
THsciRp9kaqNIjmg23PORuFoMtLeQdIzjMZ+3Qr/WXPTVCVuk9VYrMnXnABZd4Ib
aCj6wwxsaO0eM8ngWAi5wY+7A3JnWZq2HFqqp031/O87zLjORGIYAWDgp+2g3g1d
DIivCdkl5AGIGGdf7fB/66cHyJUH8u75E7tBbHoP1csVBZrsdVrdE949Fu5LoD/Y
r1KC0CO/OLggK5emDQyMJHmVfp9Xq2Tu8ZeZV4qO4Gay6wF1shqLtGzdQfwQp92h
9Rc2M9xGbPFWzMV9SfguPeXVJL2h44V3KG1PfM47NOixrvUzA4GSlT2HejXOdbm+
I5jJWXdPGcuOSDNNEAeVezV3SP0yrEPlITOX8JGjX1fxRli9KrIwJ0qZx8CVsRrE
s4P4vSqjXUWSDhR61/mPoSihuWyx2t77CCyCJSqGwsvJeFLD9N16AT6VT/VonEEV
3LptRn2Q+vGrwL/J2iN222uiHyDAEQrhy0Hj8gkDsWOk17KZKN5/qojgIP55JETS
e1uKCqcq8CzmKD3yy7vcwHxqjArvpPW85W8oZcWygfVFygQvocH0EPNcs80m/uKP
ZMoYeGel+77dTRSoohjk+sSeW83lLL6eP/qdlYNAjAhKl+etos4Mnoxw720yZvYz
PgiRdvsRohRiQS4yzhZSNnPPuSnJJeyLq8pu3cEba/oSq5+bhduTX6JlhjZ8egjV
1y3V+a3cyhrDzqRT0h/8gL4Un5KaP9gP8mDKm7TDz/Sw4f2hAfJtWY1muq3cOjWi
eZTS7XqZqwIr++BsW8XObZL5OIFNg+1fh2MFxdvz6lHWu4JwL9Jifa055CGqrkEG
+SfrTA6673b1w2sZUaEEdrix3um5vPdqYMsY1aft8IDh73F6QJ4qShOhyeS+1dfk
pxR48j/NNrpTSY2iYw3+JiGunr9oqN1WsF8A37voQSMpA4Kh37QNFtkDgY4pH1uF
fyk8PyPsNHrAmS9437vc3n+b4KwUq/dVBU7Z7lEQO79XULEukHIVSDNbIzByNGWE
yvLUPWQcYSfLfHSXMW2VI/ghVfGBox012dMnmmmAmLpS9pMLJxzxBOA2+BGw4RZV
4vrbKXRVvKSRRs9a+9/VmcJ2HEu0sq0YbkUCdqN0jzP8LdHIc8yuEw5Ggd4LVqBP
bZ5m7I3ZWayU+KvGzsa/EjR85+pE30xA2BfofNnvvkoADEeZH/O+xmagkw91qOrG
v2MBlG14ymtIXHCm7pYeMObvMvqPRiT5l9zzStCd1Moylx+gVLOY8u5ub37/U3a/
wCLoHYuw4BZ/6yH/hZc9gSWJjdeRa+OEdPR2lQwaicwu0Dje00SRtX3OiP3WIPPO
M7rRZIHqif1Ic2LymWdPXX2pYao4CGh4WfQZx0zWPMScTf2TjLn5H0DOQXu5wbZ8
jm09Dk7K+rcJ59IvQnMKbUMu9w+wqrDu4vhFfYnDlaHRmkbdEOMoZzKuiphImhBe
Fv/rLIBgJJ7LkeGTcpUCltji2YEVZtXAaJXZWH88xl5h6gf2zjEEojasCDsK2bTy
wUv73i/qbA3pLvqKBJhWCD/OsG2KUk/BQ/rk+hQRBWZSmL48skj8n0mr6z5fyA7l
CKAAqA+JeKyNuTCuPypEpHZL5khmJGsAumcn8TdnqfeYzXAUhdv0KU/L9JmQUz6y
88JkPmujQiDaRb+peNDi31fZzD9G/MRRkg+mldjUz4fxE0rKZOYvIi0IsBXx9K8H
74WkxgFlgDjSRtWBMSC7pczRFz8E8klymgx6ZNdGUq1elMPq/dOcLdoUFTtzTpMU
ah1IiOkQbOnn5+3NMnqaqIq99RD7VtmAtkp6xXrboMt3VD+5YG8c1rpdK9cYwq6E
f7YiacvvmCodphBHmrhxQn8QmNMI2F4qO9otr9d8lStp3QvNZ1Q6I5yWlUeugA9J
x6cnIWkhE0/xqIf1IgIem1zoBmkd7Twj6OdrJ8+6Bs+QbelWHCk1BSpy1EQbnqcz
qCWV5OIs1/Eycz8hWpi7DJt+k+1P8T+6Alk7NwGoSUWJzUuXo5HGqteCO33nNIe2
iymWfLi2GDCrxuGkdoeiFTLj6fjL7fg+KvZifshYoLjigOePgDfVJVQGU8q2NqIK
txCsetCU+7L6ivrCUQFjiLPWaSxNHqn3MH/FqQ5caQ4/fi3YEJjgSoJQmJJjuttZ
lyFBFUc9p9vzh7HbluMlkLIsG9Jn4HPWUU14SAiFYpEzRUf+OLrsmsSXKu/KVWyx
7FTRK2bNTe81kv434wRIoyvRggtzHz8LCeMAKOWZNyzdNyT6QhbauUL1h2gMUhv2
Vp8M1Dtc11EaOqEieBDc8h8RRHPfn1LTvYsmgdKuqPbSYbfit0lkS9uFU4n32G9V
lFFzgeNiwrV1P0wKokxY711kyS+ojsrE7y7Z++s5MwwYPkik6aRHM4sxfqJhyn8d
zj/tFczULTxW5monIDrMbPGB47Q3OUF9YcWFY+sk9Js6KfViTH2N8IaxyRr1T3Jy
eONBoxmpvRPRRpwFSJiPaFD7Sv+1abDlY0vPBMzF28hLLuWrNwVLaGdMss4hEmZ8
BpiMAsuwTy/nbEAA72add1dXCktW6JPPOQ8fFBy2FD7Ip+3mjINu4FORON24mdw0
+1CR1s27C/Jb/Kcw6ZHMeLnTRwk2mtmxQ7XxfbQvtC+OOHtXzRK/HQ5kelKWsFeP
l6qWDGJb6Yr4BTjRaSoXizByMfCV3lShyYHeLyR2Et/cKXXvX8en5lvoM0PQakl1
Ikw8i/7Mgy/Clf7EefuOyyk92gbGutRq/+FCkyugbaF1MsrtDbr+Zrivr6RWrt4P
AZFMnbyFY/DsAwRvq/px9jnbOzXXJAhCUwo2kp8Mq5eUBisUwllflYHvFFoN9Zbk
+pBaXCM0LrfCy39lFnJ/wumgnBIWlfrX+yzwU1jUhuxnkjnouC3qf0W5i55pw/8E
KNQfmbTJvmh8N6Cj/5jEBIq29nLlCeVXaHHQrmaK0rra/4FDeegG5oLin+NxMEL7
5UazBBjkNllTGtKz9rvn1/H/qLE/9FFceXJLEjQC7liHvOJW8C61PiHv4GrBI2ai
JISVpbu/CkElrYdDCIkZbby1b7z7R7IN99CJwLpOoQZjccgeYuTFMGCGOeeqCfll
7Bt773n+/lJgwsGsG4LtDOVVHtE/dAPdG7+AL1hmeXQoynbW/vm87VjM+6vTGBM1
q4tuLdSEMW0bwSEFgV/LIZ525MZkNGmLc+5+NPWzPRRmOCyxjYRGgpcJyicjsQWi
fMfjBOKk7cijMOg5/uEgMYOXNssBL01tfkXs+9S60WyEy1/6MUZI1OVRec8I4F7o
J4iz6GxAWubu8E+gvzXKYBpmXmxzmgpDmZOKvsjxzRsjQ9Yt6FRCkLpHIrRnodrx
+meXI+UfpluA3HMj197rHKLfuiUrf0tWzecKWJMLcIGM85dz4bwt3BPR9X+FUR9T
2Ni0ObAiBk+lcFqk8AZaspU2SJ/XTfTMzcwsrF7L30nx6SE6bEdYfSTHfmcUDj5c
HcBBVAhuyHv5dQtVBf3Qlg2sIDLXO30rhsJRnGjNWs4bRRHQq+nV6OxB7mzRNllr
W6l/+CiR4rse9CQLt5QjcgY+fKWkvyRXdCN3h2vVpyQ3sKzLFaKzI3hbdqY7EunX
IgSHJWmJq+Q+ew8coWJaQOaVEW7+50DWdwOMk2LRasNiJplJyg4TDym1H5G66yJV
98I8poufbbUF8nqDdVe1KT2FnZmFW5Gq2Gx/UEsGFtW/Px2H3o7Je7V4mlXUYLTT
602R5eNAA2nBj0/s2SF6FQTHWGdWK9Bk/BieNd4uwxxMbI0nUcRJwdIWyjlvBLTl
2IphNeL1unuHev9gHihg6PP1rpetGJvSo63v7SCG6AV9zWOQ9CNIMbeLFMfSCRle
6xfF5nZuTZbSwKM6p84i+ww7Bzr9Qkw8JSc/otfUsd0xqTVMlBA2jgss6jOLxap/
j1of8jHA8WUuHcy5xkMfBZOGb2jr2zAlH5m7jdUoZRGAgr5O6yDUiqzI8KniU89j
Xex84l2T36fW13U9m8HtWC1vP7VdguAcJEXBWL1wtkXJnRJih6E1Qiep4Etie3rM
AJsT0ysbG41E/8yIETzgtbgHK+ApyP9jbXs7qehD8v5inAj6oBZ0XAxRD7P4ilMU
mmEA2jsKB0n4oJoZ+Tzm0YjwO53pFtYhJXmisKtpz8DA+mP5wFOCCzyDRJECK5e5
ERszaf+fi9USLOs4wNyfGmtrkELTYABUzaT9Hh1OdSdwUVt72yni2fUxTz2b1WbM
g1m2U9SdthAmu0WTMcE31YYOLcRfXxfpCeWW5iwBV5uWnEYUOAXExmWZ93HuAM8H
YHqyOO19TTb0U/Ad/YbczA2a4jigPM0vsDuTblHU93JTgtPg9DTjLa8LyjF46v5J
Xn6pJ15vO1PbetpLABiCNGftIR4uUaeQFWrclJVJKQ9qZx/j2nwcg2nxxBVd8/AH
xnAvXv+dTTo3UOvfeo1hJo437pWudbKNeUJ0CgnuCRdu9ytSSaYuh5Nz+LAfTohz
QAV7MmG4Y4+rm/Y8oofsuV0Y+IlkA11StHlPLSlNHMT7vfYyChDGxtHfjrp5l2eN
5Qora3yP+53eSNz6M0wvGbOszmmiWrcWaCYOPQ/Mwjrg0ZSYklryt3TYdu+K2ueF
MXSScPObWJH7ispWYxmcAuBMvIaSKpY77gFgQHKB/nNv/R+VKxSlGG6+kypkkHlQ
ld7GDGlvuz3rTO/Lg4UDuxs1LR2R+TBUGWpLag9rvP26qo8Or5qmPD/uX5BqgPgK
bMpiwGHImMnK66QOnAc0bu7LA/EM58OzM5fEjAd4ok392oGl+zs2yk/7URfk5SY7
0dB3ipbB7FdRtxIP1BuphR4bs2/4qLnitMhaazeDBSDqQ5MDwUXLUVE1R4WMr+DY
1vx/OKVF5ae9PyZrSyvXinD75/EqKQ/FvAl6DznFHRgVEeWGqQ9ZdglqdC/5FODT
ZkrsqNC5+TnxzzDL2sTUwrQDBposAMwZ+nnsl1t495VSdPfAgZ9GF9hR31UuA39W
X30XRgHSK7S82RlpqHARzhleyOVjydtxpeqBvwl3nLptitbvpOxkRUPgtOXlStDU
UOrKukhlMpNAR5jYCZCDL/h4I74Rhi7qOae2JRNCPetsQQJF84Irh5U0B2n2g/RG
BBfL/rGkcC3evCUjbcTdhEIoB3UiVHBSiY4cEX1FIjPpG58kBrLj9obiosKKovps
kcYy3QG07sK09e5RmDd1xXyFK982SipiqOZinIGiBo4KRJFcfmLgspgF97YInhss
Pzsxhltj/PeKmBOhQI37sWWcxxh/UXlBSRKHjmqWOYqxJmd50/CbkvR23QX2BVTo
A8z/ChO5/J8+yxeAkHtYG9iMAPrLwnANk71jKNzbLTGJoiTSRiIyInfvVuVpqdsA
R5En7Lt6TseFP54ioT/ErBfsErpQmJTi8rcyf9n2OuXS8licrgeSzbAy4qtwSG2m
CmiPaUF0OJNW+xxo1AwgtoEGzvd5w5hN5uG2dDg7n2Pwntwb0cPklWTS9HdbXF/J
jB+VlBzDdv3fJCMQz+y6HhVWlfbLsKrZkUZvilYQyrwGDAAMno+OWh/Ke85jySac
2Z88F9ua1qq2qATbrO+4GoeACuImMouzP8L/u8jAeBcu+C5NRPXAg3MZgy6r1OW/
8PP1AO+GMdzoOsemQw4YeWZiUvcsLRZQqI5DwRLDTaUEVq62dhv64SKeC7zWEai9
/3+gPpxI9avhNrqSQQN9xo0xJ4yJ+Ei2f0lEA9NOIVJv5/WjRyzf3KF3lKP9Ofp2
hJW8RDPZZK3u7fKa5aSxMMHdo0rrPxkhO++3TrLKa08bzizoIBdO2TIS9EIhC7OW
xVpX4APJAd0uc+9tKMl+W+2yTwZxIyQCqnAipASqTajI0nKYylXpLda4H/ezcyk3
p+an/4j6djyzKp+zY3NxMgNGV+ywiU2nZBoPVMQ2lmv8oEgoplR1rgX7BDxJjGCj
P8aL/KYKq/elZsSPMidz8rQMmvQJc6s+GPqqs+GTk/5tnZmqucNGkwO2JNMB3OrJ
W80rrt7bSwRASSbSaZ0ghasIZFvVl8U244nh/7zd4RijpQC67mzXWxh6ws2Ubbo0
hvCEc/dCR47tjbV/Y3aRO+xwib4kiFd2PXUjfOgqTfgDX7bSCCHfCaFx0oPoqMrE
ABeTYL6fu1ATrPGf9bk2r7yBpDhA0gcLyhYQKxtYkIy9iN4EW8kw4totPIPoDP1a
yf5tF6AgQpi+iR6Y7em5XZ1GzEoAckrR/LVfgH8teGnJdpfx0tuudQ/4YdRLSKzS
9ApE8x0eG19wbynJAf/cMOXECElbbjx7MQaaT6Wyyi11vx7hZNxFdbU4yNQyUlDR
B6nUIVXMPMhFfKzMUOOX68NSISJPwc2zUEeBatyJgqIae6rC+D3AiONfWJOuoV/F
DtLwAwSSJuYF5IDD9I6AgTlWd/I5amB31+wwsHEa/t0kJjAAEC7ExCXOfaGeX6gu
4S+sEe/0c+DWniGmZ1M81PpRxiX3fB0Ok9cffhgvS5bR+RL6uy9lBsuYx2WrYoLK
Yx62+TclxChEkjojndadhV0xVWHmhzL+W/HuJIX/KoxEnay7dmXMIR6Ju8tIThGa
rLeY8XTY+ACnwh9gRCKShlHHl7pdl/7EOg4UJQlnDyhgwDRuqEoE7zzVyFKUj4QR
93zDZmpIPXYB5RNiBExnavn0Rmab3RIY+5LXwifQxwOxMf8Jr7OW7moGJby2l/Sq
Q2mHyricEzu1nzBW3IUQHO6nKIQ4sJqsV5zTanEYGdglVfb++GrdvXFtvHra7q1e
1xFsRfcN9qc2+E1iAQPLEf5PDKGX7plss09IdbWynyPDfOtGPboXc1TKEaG26bBp
G456pB51fy6CRQbr/ECBXX4IXe0OVIKenRPiOi5fWX+2PNKVOnLPaLxq1TffvuS4
MBaaesOGCNJIK8g4bLiU5l7GIV0uJma8CkH4Rw4gW+YEJr8rQ1zzRKhyCPGC+DFc
91IsVhKZOgIsCFBQ9uln9z9IgIefmtoNmbQAvLXWfORyxyIyEZpA5LaJzoj2CQw7
5V4nwP/H8pg7m5X1xE0pZC1eCLk3TACaGkMs86ED1s2/oYiOXRlNq9L+zGUa2yWD
nMUiG+NfnnBuwqU1PodtTmagpQQXWSxcSCua4AQvst7aD2xr2LbeOkHCZqbOSqP/
dElNajaG1mXyTAWThq0PNq+Mhb8EQzgzFSHf0phbgHJ6x6Pd/mmy3QHUwxiUGgPb
xDfsUefAlN5qsaMRfuGfwJQuYg+uCvNWI9v3cn6XBIv9tLnHNMmCdp1FcE/BuEzA
RJEY0ioOfvY/xB5TjG1q24xSyNH9PU9Z/3qbj6Ay7/IT87CD0ZVp62nS/t4yXgeV
D7xws7Nd3nWKOeot9cxw4iBaQ45vAdGvJhYl7lI2z2vUJYbDrHber2jdTYxVACpo
IzQdLJmejcQqsJ2/bAJ3INR63SLJ2mSWPDI8CNeJW2tjBFtf8s/DSs7NfG5PlYeM
/73Us9fICkdQug5Y78ouCrEX+5IyFYR/ud2nKAy2Rdrfb7DNsaGAoLM8Y8wiyBT4
+pcbpI0nc8Ux9bOSI7TIiPqYWtgFLtAYrmywTEWulI8cHEM5IpiSf4HDjjUeJvx5
4ft7xEgCzjv5BcUNA7k3WnOUCQQOhqpcBn0UGxQosTNSGjESZqZt3D5mktHNdmOU
qznySjdAz7IuDkvaGnyn9HeoqMGI9d/P2pPntSZ4vke8DnkVLdqiyXDx8uLQyyLo
WbMt1oE0kssW+6+f8uDAz3RR2vMvbFgU9ibYA3Wn+L9bdtAkb09ZcAJ+gdNskGQU
tnBqalNhqhGGDifH1DgH79WgSp4GjvI896qe9ugo81SZhEn/GkQgTrrrRJ7XBt4j
z90vB7jJfZ9rTdNbL/CYZVtGx765WYd0CwrozspBh7uit6sg4WFN3wqRQnkbTuS1
kzbtV2CueuY9jHv3pSwk3FEei2eO9CISb2OZK0QUhRmLDq4/CPE+oUDt7rNCexYW
zYNN1HuOqCGdJ3p+84l5tlVCi7BPJDAF5fCXIwdzNo3KkUz8vzg9Ev0PKwWQMW54
WuYguEF1+zirjVqGgvB9DjhV5Ye8dn4234aVaM9bS+IulAYwdjv5vZaq2xIeu4io
VyLQBmXlHV9S/4dotfGKDudD7ZxzUTPf5E/XqfuZeamgo8m7+/CvtIpVkO53KfB6
zBiCHXyhT3O15hpimAR4ibFz++Q9RP+UMys/iu1GGCOdHKwgC9SUtUWcTveJyl2K
fktZgCc6bkaMHSqENNC7Xr6dI6r8SSpxMErspZMyZXF9apYDMWIXXAolyZ+01bDj
wRkhjn8QdtknWbJx2vA3F9khZBgKGd2BjbVq1HuRPSdqUZG90/7jNENMp8fsBXe/
o3rrKl/zxMqOCcKUhqejZKdloYQjguZSso32HuBEUbFkMlkHK0N9dinree33xIv+
3ODMSIF+yzQdBhduiL/jKtbQLme3QDoSdpW3bbtuRL+RA7emwFfehc5iXKnYsMO6
Dvu+2i/0w3tUp1sYPFzzP0usNFSOaipZvMeOgdZojYs4eXu1nY9pV7P8xcAzEi8g
ucZy8aHTSly3H+eRYRJgA76E1svjEgH2NR5atUdp21EeZzkAFGcZ0EiJ2KuFt2b+
zrScJF7GJsBQfm4ySgw06VDsg2JoZsIqa/uK+uTeQacCFw890y6DKiwfij8RuYMi
7y26Kt9TcU06RleXsvgApBDMgg0Vq6SQhXkhSOHZ8U+k/ocssz9V+0pNObzpS1io
HX6EeqssZwQ0cbsKYHmCY4C8MmtDCnmp4f/yBPRSsrc/oGn6TRw/TNbcasYm7kfs
AY5wuFOkBYybZmjmXJxObXvQ0ogstSXrNLtezkY6PWxynrN1uTyNYVxT2OqsFxoJ
cyXWjff496pbbGzVI+iV/yQKvdxtrGtlI2UAmMF5Qs5n19ctNRKJe9N2YS1bxbjb
4Kq81O2D4qeHes92qxIPq0qt9H7xDWNccxN+JGHSNLgneIvx7gUmeCX6EEjIAE9N
fWLMypTXBmNg4KlLvrqjA+78ULbtcbUwryVLIEfREvzsDwweA3mO6+ryr9TNRKPz
Rg7q7dP1GGd6OWUyY2ppCKUMMR35EJQBWhtMQHL9IV9N4Y5nRTehfitySUDzcz3E
Q7V/m2yVBELZnmID98frp3b8mtVpX/tINpjXxm9R/wyZme/r7IjwD8cfjFjU6toU
2w+5+8zfov7rEJMJ1eBm7aH6UZpTTKUa3G8DFL3L499Bgtco16mUA2ossL1Y0zEs
NqcqyIxQeYyf+gd1xW1YUYpocMFcnFXfP4/8/C8fJVqeSZwf4soX1ALC1x/IGCUJ
NG2RIDiotYj80QT9vx1S9b9ED8HEIdJY/3QJ+m8+vgVuQA31bfDVvrixDAXxoqHG
EdXHb2Mexvu77GEQv6nY8TTBsF0LkXxx6bQhygNBEXGKZX8XQEABkPqunlIbwccF
JPzdgz92wjQWjQPR3enMul/wHAxxjLNyX6Qk+2o5BXxhVR4GcEjv7c+kw33U3PTz
PF+ZwAQTzYc3G0ZG8JmLAqGJ2vy5iVe79JLtksVQUx1cj4nEe/AZsSnQrkXjEqXM
YGpSA6fjclMvPAVO38e25ZyzYif8UEKq9Ps/Y6LBFygh7B3tXHeOOvwp5P4XFPZN
Ch8RXAU4JLnCV/qoAHDmQOOS2TZ/j29Hqsni/K2y7gswcgCF3NNncID+s1mUGft5
2SV/fyDGD31cMZbMMpwj8ws/LHKI6NiTRWZowMbaxiOMXi5IhgOiqg4PdpPzIM7r
0vHl13f0rp1cvWVzBdY3uXk75c5wUz0j7CNN9oNKcM8JimyfRTffWcJdoFhn2Bwo
mWGuExFcxpPg9O0UqM2boXhbsaMimAEMABQhgNQ0pQq3eRAPmb8qLhqQN0m5eet9
xEQ0QJZeZUpFHkAAeiWVHFmKEptuy5Vg+RDsKFYRz/pgmi0Cv4KbqbDnLHRMse6A
YW5A2LOp+oAjMjocWO9el7afYmqz9sy3Rqo5JfIHcDV8XrzrUV9Ef2VJkXbKviPi
Wl3WoEQbPm1qCR0aD7vaDjytksiDh1VqFlEUPzEMnnJogQqPnCQWff6U/AXp9VmN
JolnKHu8J7tF9902ZplGQXyflh931F71gnEJ5A7jDWsBfeHBpav6lRKMPITVg/j9
tGCagwrzR7k/avvpES2eE2NufzCXauux+SUScNzlXKTa+Xi3EO7ZdCw0u7QQ9LyS
DkaJSskABfrh/o235xdQoLelDXYyWNQmbtPfOGOMB0K/FpiDvuwmsOB2gLwj3Bi8
XYMs8cHozBUwrR4LuKNqePtKEoyybiro/YROUNs3wW7s+bwwh/+dDsq/s5CMwO++
/rO7CZWh8/BXfYO6wwQpFEMjiz37ELTNnu6/IcS/aJQ5HJVoeCfbvHsBpFmjTh0v
f+haFvhI/WRTHw0VAUqrpsoxdKfoSPRs/T4oUa/XzG12rjqbDtMjCoV/gitd2EuF
ivOb+QkNboqiUOhSoURCLc+DxTcw+447mCASBFV541zyGheFSbuUmwdS6eYMCJ+F
a1psClWvkT9a9o8cdpcgZDCdTIwz7X5sOkNOWiUkiKDgXSmc/5+xHmqRRoyJH1VR
wy0AotqrYT8KW04ZqKcJcqGIEu+arkrnM4NCtGtuw62Pm+Y7woi+wblDR5L/SpD0
VOWFXpxQCWP11JcCOK7p7ezNyRVPqRQ79GcQ2KupDnY9i92f3vbye10OVtyhP6w1
3CpCaxgkxZjsaK++NPeV5Q0Njlzdl2j6Xw2VisS1nDpH2wxbzGH+3STc5Syk/wzf
M17Jb6thM4ucKnOlWHsDMEWw77ZSyKi3V49+J16vMWdZwtkLIOLai4+p7l9cHa3s
IqR4szLS56wqjiA0HOGdtPU1nzGLbcbuGqK5T7ejUb6vcrtgyuc3j2nAsl+heCkf
zpoq5mHVMpr3TvUDxCXSDVBAPsyQA4xXjus9JYAsiVYc8hCiaJlmlpeadiemoh0F
qXRKRDS1kQcCpQ1TUP5V04iRucTc7k8d+/0IIP/clLIkENNHtCqKjnWPhXwVTB5e
rMio0KMw7RoyeLKt1sz7d+bG3IJZbh3QeMggQFcMq2x4ZKY5dMOYgFfRPwNpNWji
rjgxWpufe+cswCn/2AwHvYYLK5GZHsI2oPvIb76fUuiisruYqFYvIpPtMz5o0el+
JMRjegfF7wPBtgGX6M4qpPuRCxUu5TlzbYMVTEHXAhPcBkAcKhqp0NHqx6lsBg6Q
14vrcia5w1AbYBxfm/bJUrBFNGMfDDDqB6C3RWsYNQZdGpP0P01hqhLrhL0hK5k+
Rt5L4iuRo/JUpdaI+zEV9GiIz0cCqrrGyfDqaMyh+xd95z90pHryDU7YgwiD8DNi
lpGo1uAPYIUlzsJOqXDwHv8tkuvyac3PqAG+hJ1zBvmQY4zSNETrQd5xIDszmQwa
LXZbiTd7zsGcoEVw0FDdjkET3O2D9sMZ/AIS/5XQ8SmAxG5PRQzpLG1H91XGA18u
gyMtNp14yleLWndcYdGZTwlgaplGEWeVdiljKYskCjUP592UU80NOr2vNdmrTV1o
lzGyYKS1In0R5hC5qt3/pnQa1/D2eUQGx1X3tt9ms4a5e9qR3WfnTu+gv9o31tgd
xvBbP/bpuwyz4xok/Lx2AuQOsfTa1kNYtPHROh7iDqmW7abq93Fh/Yl8dVLI+1wL
LYjBRKIFev6KCrIbDLNVsmvR6+NQ1+GrgQW6VhOVxfu1l4z8L+Eb4W5BANY7Caa0
7N/wgwA7gqhq+PXSYVZp8qbd4shuK/bZ/5HV3jr7stX/nhdom8s3kPEiF7npQ8un
AkenVRpA3a5yGLkcTDzu7m6QCA0LzhHWdBRkcLRSK9yh7J2jOAf6j6v1Gzoke5nt
1PwQ4AnoCWkAYR+dsCJeKYlrpdWkZ3pHh7dACfLdyMelrI8gTk2/n3sAqlR5UzI+
u0lsjMAT7Mw/iJkIX7OcONNMGwU6mbN8uJoVWtCtp/ytTBZaW7azJzVaPKUHEbHR
E11XXTlA1LpgeY7RO2t8jvL4uxqbejh02pBTcu7sV5HnRQrDRt2/Doc6cGf/FlKc
iDk7b6/4lS2XDycAexm+R1keARAu+4o2zLPgmORgKF+QCIDnSL25/NEf44PK6RRz
um4sqyMosySF8qFxVEZeKSrURhkeolne8aY/wAyQmd8Vq3CS8UEvHz5l6BGNgQpG
+7KV6r3APSTyFI+u8zkafhsaG9ArXPLzd3/8chXB1h6UMeJwMN9fYj73gqnNZ8VU
mW6IV9Pa2RUzunJQQ169n+KywQj+KWpep2np7ZJeIo/z+pS9hvIXqhp3loF/QoKb
XkIsPuofw+rrhj92RCY8rGIIYiWcbNS6d6lHFg2m0pCjlbV5DzLMHFEs9hKkbQcI
jvYU5du1X1aSzNx8fIXDYHdJGNjcz+BykjTrXswkzjfGTOD0XCQAOD00Md0IZj0w
nD0Oeha4uRMCW7W47YCMTXeqAqPkWmCOmlJ4psAC9DKtceIiLXK8xhfvhkG1Q3nb
dCqIbsYaPdvmayjP+HJUg9oYc2+Hphde/xALPGuQhkJuoorOcfXMTsN6B/t2BAsD
E+7GaQIdcpsQ2NZ67CcMXiomJYLQgFPbFHVW0GH2m2U1W2BaX89eO4DHakwUTvel
/8HkKZelxGMUfXfQ+HLVd1r2HUuI3CfdEYLLoxD49dBr6SsYC8kn4KI37uQAw5L6
13/TXlCz/i7C0EMvVaw7xijNQZLKDDVGetG9VWtRkFHtq6e4pS/9f4jNbllPHbXH
aJnVXByMQabsqgt4q+VwHK/CM+T5Sd1IawO/1AXO+ETt4LNxuwWAzR1V0CfAXAsL
YZK0ksjsnPuzCxCqa3PV854ynuNKpppf3XqmTncaGqXrzbUe/Q1KDhGOfXrzhKbP
YrsbcZu/ExwxTqXyDkfXFfP29zmDd4Hd4Co1I/LqDZMbZbJ3leBPqOgmZMsrc67b
kKp5klXNIntooqcxW397Ln+yQO561nEKAAFdnp2oYMX7phnqo0/8QlMbPbib/JT9
GfiHNC21KOO6+xeu4h0v2JhTJgnxe51N4rJkAlpCV+IA2jnFNjtpm3kiB6xXRtlx
fzyRgmzpbRmkkWJPEK7ez+X8056IgizbrGj1pyWrPku0mSjX9OCin+4LhuJFo3pl
5LLIyybwvlLPn4hjqQ7Ey64TjEoB8KRw0+OGTf8yZd28S/pCT3mmEjMtnpX4P0SB
ZE36yHJAHVWE3U9jdwTEd3htYrNmT3rcogaQn/YJTEAO/C1ijaRE/eFCYBMMhKRU
6udQSJjN/Vp6d01a/5Wh05UZUNIlWvvZfZmuVJzuge9Q0B351Nd0caeFjfU4QO3X
O3gzqm9H9hefe78PXsqDaQxI81Xwdf5TOzFE6ombPeazkrC6OllnNXf0MJIjkVKA
lVfClKImMggzXLmvydAcRunRhFRdQXHsWoX1zdutIxvQbGOfEdXj+qxWqemEhVkf
KtsHtnJBjHesmO2m0nIPGDAKG4sLpd3c/FBXSimqIVh9I8KQ+Y1342qNU5WXHu3i
9SDEI6X67nFFnE+YwsLwJHpbHX2cx9Uy/n3Xnp20fEp1iR9eYu/oBnG50rJFx9jD
jJrSy8x+f6r4p+0I1giweer5np/PhHsUl/cblR/4NXPc4/1FX1lNz6jOP5dXjWoD
GO6K6MFgjzS0AfANiIZz/YRRRirZhxNEAwhjPd5hZm8e3EfmkEn9hhLct5Qx8b58
dyKmcHFQulz08eVkXgbsksMed0mQFYv6AvTgaUx5+rh8rnlV20sXqRI/ZS0wYWt6
NsDisxW19BJhLy6oyC0RA3oaxeDbeyL75PnHhB7e/xBvpplnhBHyCqbRktTXb3eS
1qUq5UMahjPj9ukcHi/Ed1NdnegSHM+n0Lxp+j3TgVuisd9WZEMFYDsx85H2QkFu
5NBV4Gfr2j0VwnEqzdkHgexsYnYmIN8m+WiJjBjA9T5P1rPMiDfPShy3EzFzWRe5
RN5KcL9bYBcleTapkRsC3Qi3jWbk/ZuZKx6o6W91X3KiIzHhvjQW065uZCOzBCLe
qv74ZsKtSL0wr2L3J7CYJ7rWK6B3p9FN6k9RcysX/jqCSaHglot6rQZESHNlP2lu
AQKBh3sqtxlT/8NXFB+ChkpSPxUqFKn8NrT9KPj0uEVS5l0bqVW76GQM9iIicy18
ZfF23iA6ias1FiSBjcree2LAb47QSXb4kaffdyRbYaGJO+0YzKa4VN9m8GkBhGQF
Jl4/TnmSlIBUNZ+K5guIWNiQV5fLVTyoFUh5JS/1xREqwX8wL2h3GPAyZq5RR7OX
2xHwINR5v0kEwf6UjppJuL5NS18TMP1roi5QM3CZ81go7zi138JL8Hv0WxStamxE
bMf+Pt9R3I5PAxdUWtvS5CRuEa1lCahPAcXrLQ6zCYI+zf5pfGsDtfaV/oHnjHSI
Ku5fZP6g4gt7qEC9YVOp69y3t2TIn3YJlgDRj6+zxptQDz+IkyZWiPWyoAxQLIZD
/OUlurWVwdk9cz66xOyVJ593zQSwXOW9JB7Cy5GgD2o3floTGlbkP2i6ztP9rmbQ
Kro5Z78E86D5ucndRbqaIL/LohqHQ6ayO7CjBcuNqJqRAGMz29mYIeFR7z+G3TJ4
EhdHvW8ks4c8XXKuEAGcmH7pKzBNM/jXhMYSDPaK2bcdSvXWwmhUIzBDerJAbdA0
wnEuJRgvwBLsi37DP2gKsfGYRG8OoJ4aHm067k8O4j/f6RVYJW1QFZHCfslS+b9n
JOnpYQSqcf2WxOQfcGPj6U/sIg6wUoU8oKHvpqoBUPw2AphM4Tgd/UkfykPxm69Z
bH3vurhro8qiB/gmlnofKqxedxK6HeL3icFTNK1hgde0s7YSc0ADZyeSE272k3Ht
awE7Q0+XxrqswLFp6VjHfSlgGjYZtznejBqHLNLzyx9fJtj2O2fRD43vgD4JJRLa
dqCDJ1MlRlOQgzL0SdWIsjMdzhN2YN2flVC4NUbrcMTGalWQB6SfR3xbBoWgrn3F
MpTNcb+uRKyC3Do8TprvZMrsFVlU2o7LKfjhltX4w/C7UivZHvlkIwV+LMPbM3pU
Lu4jZ1CBJPadIveskmIw2dom23GyfeTiircDkg5U2DWwlKwqVEdzK/OULWpvV22e
njWUQxf2dSj0gh5WL00WaOiY2ge6KXkE/7bcuzeRCPJqbyvKuCN1yZJ0WhQz4tA6
V9VCHep9ZUOSS4XEiRjO/CJDsXHFGX8GqkZ8PXCXBFr3WlTWEXayxaKabmFrNxA+
31VmUtSq8WjzQXW9cChYPlGe1oqtrKE9ooMp7riMrjGheq7GvxxdFuF4KjH8ufiI
E39H7kCrw3M1RUXS8QK8OIj3sUgdp142+hzhVJ8C/NZB4eo3h+OSbFQ5ATKeIAWL
/v5yXDyvO1TvnB2KgQK3Pf4ElIWxk+xWko+/oeP2AqPMgn4pQOm7NYLwAc96TNSL
BkJ0hrfgSTrcGPWQs5sSJxrmfRTTLPk6Zuq3dsvkoEebRfWXjt1EddjzvB9CvQ40
A0TEkxBpvekUsd7uwr8SGccvSaTXLcQ2b+gGREJnUWnlFM7iMiOQjWFnikVmUnUH
2lWmHSNvF/RTZ0FgG5ppXOWjQO+ZUl/1FlJx3I3DeapyqrwvpZLjTcaP9xOGffoL
tP6VBfOBWbJsdnacj89mTR897lh/QxAAITHwjKBEnQ3R8VrYXJRSJQnagff3HffJ
c+WFvu3YnoWbMbUSaK8N2wB7w4DrD1rcNtkr8oCO/00O38QjxT/73+H0txta4ozo
wQJQVLQpUb9bRtXksjl7y29axBIwV/nvSsg0fru5+g7i51ks6r1MAKAZ2rClp+Mz
z1KLl7vuO99eNjOcNMYbG/HifAOkUPNXh2Zp6ca/r57R96p1+8hAgHNVtTQAg8Xl
xeJ7rsggPIeonS2fInt/ncUQn25atxyO00idzV5/Bztf0QzCpqT08cBimAO1G4XK
PaLgTJa4TS1fODZ6Dlwf0RIe01+0et4k328Uyvg8XfZtbLcCwLNlYLNLYPQEblZf
Jol66y5cVv648rTNL5GRmFI9vTHLgjKSJRqfwixnFdZ1dBulxYAiQgxJ8IqdOS2d
oOLPmEWJ5s9VfJMyemdR7WGnpEmG6gBj5PbCCIuxV9tOe5Ojp1qe4peD0KZtzS9o
gOkZj3RjAN41w9Tkf1a2cuDeDvr8+AgUxzqHAjPkI7uN8ONf421UL33g9sTbz4hd
bXj3YYWRXrHdobvaVhHv4XTp65hOeOpt4Ts64q/x01aErz7x/HXwJxSzMRm3Zkeu
AGF02wHkSgdHFJs9Ug4PzbwO2cSMajvBhp0TKIk+Jag3mH3M88kI0pb83otWQQuo
c0f7pWY87SOy8eOSLx0oLziagrldb1eIxwnjW5t1OebXj/W7g9waE5hjYYX8VCMZ
QJ5n/fOQN9o++117PP96ZaowTn62SxMmINAlPX76VthXyIJCGPwz6i31fFDc0FTL
Wwnq2Y6ZCYO43qntAs47OnC3j2uML880kLNLQw4ai5MDknjkRmeTkqpcF9QnUJ7o
iVxjArvU8eYGBCbZtxsTLg0Z/K1QuUMERiWHo0NmLw1fMYOMsOOP5jA7QCunVbl/
cAGeU/ox1pzlfdl39vR0XAFKvoylKmz9c7eit7HufZz/r9dPOPiDcRJ1EIyYzlJO
8Ilq8frrtHqXnVJn3ga+zBxiFNOTI268eqJ66977fj+F6plBVd0FtLV0dptEipd3
iKIjeWkuWICOoquadYvBIPFB0lCFg2fT7Nk6lM90umiYV7FRLxR0d+Cab9RgngkP
FZYykJoqNniVPUqzOsh/YioTJZmgFgYSms+jfkqpYsFLemPtQmZ2csiJNbMxqRee
8/VF1V2dtvL2A/Ilzl1ORNC8PniSQxH4qXUGa3WFvlZkl1JO6CjCUyntLy84ySMf
JEKxZbSV4FxnSYExpSawcQ5YYmAOp85M7Z1waoMy+FFDBLlkvh5C01YcR7OyS/oI
XqmkYIymIjLpoMNO6baDQtgFecHVJx9AZfhLaq4CtKjs6VoTrYoA0knBVT15cdPM
PsveLgX9Y3d2OZIB1Vui4BHRwNSMVtnwpx65xUVCD3oonDuTaveoI2n4zsuI5gf0
JB5sHjSXhNW+Q/IgLCq0koIUE7V9ws4ercCDWChWkMJJfzbY2OsD1gw4NF3Zmf+D
ppQnea0/4K65bdkCj10R9m9FLESQwpVYWoXXggRFIRRuvVOobbKjZYt3kYOec7Sw
AIg2sr0Ehitw5OwN2BKXqGnkkPTY3pwqQgx1x3X/NShe5oeNY0wkfwlHRb4pwsXZ
7mVgCc39Zm8ghNpJypJIrWamNKUZGVfXrfD3MnzNCJqZJArYKL3mcWKwYJIcq+DC
4LDNbkBhfJVrVEFC6m/5dUbJ69FJK8BqJFhlmG2Hoj6uSuYr1JdhOnWvuFV0Wt2u
8zJXXd0d49f0TzgJPOHCGqt/V3vQc5/u43DJ/IXFDIDTZs5oK2RMsTnL1n8sPSJi
iHwvy4hWq2H6hsHkXPs5Fj349u8jPpDkfzVwniwOpaIboSVTSolRK9cqUCjbj18r
8dPd6YFVskDwddwohV2lSDiVYAQLM9ANitXCuG4dDhlv3ABGZBVB8q7fxxMZYULw
QSJCHuMjdZuzLWpPdXKUG0RJXmaPrI3kcaaEScXnhSZf0UbVZ57pbYz9v7Da6goY
FlEjAy3MeUuHxspHiE8x9q1M2Wj4fr3WMeKYN0Js1E9XCXgqINMS/L+mVCAOSwIA
gpQxAnwdkntn6PgpaI/Cy6DopT8o75Q8RNn7bb9yI28zJcsmEopGicl6LxbFOYKz
PAo03wjDaeKCghh6F+i1GhaCnpvddMZMXCyFezpQgoXBgCdIv+D78M51ZWH3MlU2
BW4oLL8SXOXthL8k7GEG958kYRWousb3/uyct5HGR4xrJYW6dtYOUExnq5p7hhlu
G4aRfvudOX8fNvo+myPkl9eaOjFluPl0/S+f1M7u9OuaRbQv+gzbsb/fBhs6eTwf
ovCuCv0Xfi0u9GNzYna3Dasgu1TeX5Ed7ZfM4dzqKmc2t2YQvoUy/Yx6F60nHaVp
+XdcdY80HuIuL6vPi4STGu4Gg4JDCxQxD+kRREAOjzLWllYiDI1XpEhCr7UQBTi2
QFyEvzv2rUK8TPcAE4GUEpuf01ufh1avPKERWxDl9c6FrQ4CwxgiyKZqJRtNnWIZ
ZLM9HWWFVGF8s3LxFId1m2x6Agl2MQH3Ep/aMpj142GXeMJb2q0GspguIDSVU0Ak
+ocwXMFlvemW99F7/OBk53FXCyBze1VDJ4DM1YMxwmv8+izbLoTefUCV45qK+FkT
qx+j+DXHgxPFssUeLaMz6DkcEaea4Sl6FKQYYIJEHTH7LbDhn9YV8pkpM72FLF2s
vTU8k7UkZM/7WNG0BzpxicjmSRZD55hH+IpcUIUa01Jg0wB08yPganLydObyxaWW
6XAYWa6oza4cEMFA4cMrNTumuITlNdpiRKzuNePj7uIOEvXtbYTZPnvWIApVeuoO
e2xbM4c6D/2BSn6yqgYRRbIoooeQglckbZYGuMYsOuni1aP23MRkn+7uxlLKbdC4
um92DXFfOjHGFLrho6+gIQboeoi+IYjwLxxT0VW37nW7HMPL6hKoEmXEG6khzGL6
bOZx4rcqUl9Ic0UXhicmK3mRIfkDG1bPIm3pVkfWlic+9dnPWoCKn6WpONVHORrl
yas+g/4RtMtOQE9qE1oXV6vmuZCmOcuZMlam9dk6uRi9oX/JVBM1bPYcT5UmToQu
mAJZiwUzSRTwyPcmF2XfWXnERn02QU6pl10COGfFluBccUm3JPMevEhUPuV5YaB7
lrfeqSn/OEJ06gOdl9gow9NJ++BB8OcIjmvXlRlFn/OhVEXZ8nBMJoMASWuUCIS1
TC0BdVVRq4tQwHFYsUfwjOQ5dGWkGbLPIVncGuJlXhRJzPo03NIROrDEiJkWCZjP
SCA0YL1vHoe/QRbHwgpMFnF/0uTg7w8NUH5NzBCnT8kkNMkpBZb59vyf9bS1j87g
imQCocitJq4PZxkvPESQsQbhLBLNl5zZODYLWJrkU1bpVeXWk161gzuTx052Ps6P
RQtEhg5S3wPWvJVqLOlQlRnTlK5MPs+b2+Jqc7ZBkTGDJs7w8jSh7XT+WMa9hUuX
3AAhCtFvBfECVYUcrXxpyIhR16276z30ABRZ+Xtz+m8fyLIj5EosVvtjLTobw0nC
j7yfsOyzJ55aLRPKgSFRU2zmvejykw//nlCxRBQl92yR9R8mufktwyL/QE7SAOXv
0GyHxba9QqTiTpTN5lAQaYIOmMoN2wPqG/iRcxNAYZ2u8+lDfmgB5ZlGx8J+5adq
OswHRPOSm9gY6w2XNDiH9RiNb4iUDjytqIMRPgNoo09OYrtYQpuD/C049fZvflrz
Unvq1QH6ZDAGcvbX1z9JEyCOQKa/dVtGFrPET8bLrOJuLAr38oS+/RNjpw6CFR52
G+51lnG1fSHkx+S7tsJd7d2jLRez7i/zrDq9L4HJ6+aPriTnmUmnFQ7sjq4FOCn6
SPi/HFPHSUHCel+tIcW4LoaTItAvSO8etdSSklqmp/F5PoYEPIN2RiZjojlfvi3O
HBf3qa1TnpIZx4L1Zxu5ittufiRHJ1SETtJfPRmPxa9KNpis87E/YeAJOFlVAW7l
EQD29KD+zISnwoiwV2nHPubkD1AZmD2Vc6Tkg5w7owba+I6JPuQ1Fc//bWU8H4cT
n9E6AAfIBb/SRilEP5xTPLn34OMvJUcUbaoM4pvumYgy4KkdruHzVu0okc8irZOK
LSnCJAEWlZFtTTgZZQz25BATEYmGj71uWg93/QGbepOFG3y1HihQZhxw3A+IUJlO
k6+apbQhgYtfm3XomcAAwuWI2U5WHKjb6VrqK2vPVMNzRU0ocVk0OAxTEaDTRLL8
sqA47rzO//Y+8iYi9Kcu4EOkI9o+u9SIijExObFqKOL8b/0EtaEGloRPcY7Y16Ue
dHjwx6nP03AgbDS4rbPmcf59M/8IW8wS/Od3Qq9ku8Bkr1prVwBMMkFRre9dUyfL
tjMyzWKqhbC+q0CgxMh94m01SHp6u7hLeWS9K6OuYgu8uw9s5Q/tz5ekL2xdjKy9
lFpR+d+GubFkjDoTHyaRVGngA3YtAeNqaZj9Po/P3IHHCybemPrC40+PcObr/x6T
MZexgydD3J0NQ15lMoC0R28lgQFNJxgZmMDDiC3sFr/9w7V4vz9Iq04bBQcJJLa4
6tE7SjUSS3nP9l79Y4cW6g9ZMWK1E0aDCvBz3ixigsD6WEIPkF5EE8NaDQ7iWtxB
jHRHTe9y/BF0w5Bl6GGfzvygoBkHoHEe7nBISkfWxun+JbOV3frq0oXKnoq2Oz5f
ne5d6Tpxj+meZ0tWo3H6aSwkc1AjULmOQHMG+8Ivg3gXqG8PtujQQDhL+dt7zD4O
Ty/OtBLcFJwcdy+Zsdub07a9oMrwEA9xn//l7loJIsBDImIzNxXmxBfVR6aiFW+o
n+GUntmGXX//MrI+GJw37UBlMR52rq5qLMYr1fJvjEWEthop/OtnWGDVnL1POtZV
O46lJaK3B3TCovP4GmXsIEDWC+WKm+Eaf4hDlJVqJ9iYqqFjuJ+siZY1otv0x1N7
lPasy28pnAFr54aPupafxdvNiuFhpin4DGQNKdnrzfE5T33lDtmTqBHINmCruMHn
UWHmqxkP5Yv7JS4gM0Hbw05ItpnFb4wQj4MwJiVf1TQUrpqcCxNZk9WgGG7VNfVh
4dUJH0fEQ3SfJ1+E5drdAXnxgGghSCsvvRhyQ1SuC6FA7z68f7uVeZ92lh7Tbyuc
mWG4saXmGQ72abuDzvNkMNynZhoAl+YtlCgZT8V5JGGLdgjdagBY5uvfqgHKP9pl
t0J2vwNMfwtvYyuB8/AcEUpkDNfUyVLAlot9cfxrZFIGZrEThlMMMEf4iwFGJKcX
UjEsJ8ueyGX02ad461Gv1I5Q+EAlzabzFFz6SqcZ1mef0r1zEM5kyukr3/AKqw6i
hdaiR6KCv2mPNonN9YQg6J8E/AtYWqOB7HECzN7xXbsoDj9dCRU1qoQOQgobuGEb
1Jhvsz2/aAOvsNl7y69gwq90G1b7PR0hiQ+aHOKQ3SSRdaRohdpBHeykM8EYwfW9
EWSg1UcqoRpPGTzc+aeyo6h8xjAiEHkvi6Ob5cslNNXeDXwNdxkiXJZeZW7ZPmY0
GvYdLguxtcOvj47SaIcmC8dggX/wU10r0znkOlcstVqbBrHPDBiKL0cFnQI9NdiQ
qI6wOaEeL1jHG8xQhQfwGextwyfTmy9IhqVSnm+on3dH6xEUh3EBLQgfKNW0NHLf
e6jYMOBaTHQHJTCGnRGzJSQ03fi77fDij3YwdO48UTQLAUSS4o/hOofDRWEkMaC9
LOkpsu5Zn60+O/+aECUIKakg5iqvsRyz+q+dgBt9QfVIFdA3jIBAvaOg6/DPafv/
1EVsCcWSdObadrsfUM6Nq8CLsMBEpuYOnaRVcjazGJn1eRVZHSzzDyNMfCMey1pt
8+sY66srmj86GOntJSHXPvWBT6msDPkvAqqfE537heWCtVyOMt1ME8O+ftoCcToX
dBm2oKMITBZiLzvt9kssB2wBTaJEegsKI8o+bK+CDmIoYUS23BzQ5oQf+vYyfbWM
g+AEN1cY2EzGHTsk4XSJqo3qc3NwJyrQBu4PVhCpPUfzkWrFa5KXDAK7NrrL/243
mf0yeWk0h47sntHHxVmI6412WUS/FkkadLO6WXvGBGCS4nHSwIjBkt4BopyLXGY6
JJnTmfpZwUk2AG3uPfT86KlCxJcaNVGJK4SXIZ9M7EMtMZyctL86GwhH8XOcdPK7
tGOXo5IUPAAx4+G2lenjJByYDxfaoIrx5B3XT8zjSCgZ7SwSxEMefn8R4uap8UDd
XyCO2IfqWDaJv0A6GSfSviopR7biDMPlRP+4BEUlm4w8R19g6Cbt7vYQuQjkwHuX
JTANlmC2wGG7DV3uQ1cXSYLgTm/c72Hvi9OAD5pjwxb4VK2Zt7S5Pk5Tv/rgmueJ
skj6scQnJEIa/FR6CUqsJJ5JrxRTbFfXn9LXWoUugwxTlL+dBS7TULeIoc6yd73B
2HSvQHS/uuTnS4Naq5KxOfLee7t9m2oUaMxhWiJKruFyLo52Ach1AoVFeORDVEvd
k+56yp8fguadgDMRrD+Ta1PobJ72uC6NXi8UTZEbG8vH0RsuDDcoS91AANRi9rdv
/75B9EixA+XA7VAlG8j7DGRVaPbUjmxEmOXq9eCbXj5oUOfR0y3F8FvOgNgbCae/
JOnOahy0Fnkc1efh8NWCCDMZ99hZF4jadYcXSXaTEY1T1JqxIYe7Ir5clkSI4gCz
hiazMvSDIxbY0II0sb6P4gla7OtkQQY3PiydB/81ZpaOULEUKB9dBkW6KjVdMjmk
EAN0/F6QgxYFQaGeYDvXIXK9AZezOGcS46lCvMeYUprhSXF7h8m/mS7Pw1kw2aDA
Qf6qCcf4sKYmH75bWnKDJPLuyjPwKcYL8Qf+0ulrIatXbAujJVMJXI98n3gFNglq
f1frVp4vKQ2bzDQZRCNeOK7PrCwk845LClQwrs/6kCEH4cvqJrpKLqgzshAwEghN
eAd1TpTUQQzXojIvsj9jH6D0rhtv/Z9LKhnwAQE6/RC3qetyRYlv3S7q8dNNni1l
hTPSAvyQP2kkVWZQFvfERePLf+R1s46Wx8xj4cYgl+OUp8AY/Q0c/cmIFiSw6cLO
x7phjk8rh5RQ+ET526VfUEPZP8aUyNVMFElHQe9cYUfWg/1oUS+CYnYIOy8fSQRF
OIe5v1QP6+C8+54H2l2zEE9LvQMn4lnPDZuCDp0mlVskZ+MtqUoJhQXqY63NjsBv
7ghqjWLfzdt5BQxewXK9rwGaLMsJ4cfB+5rwCrdPqPMZ1a6Epm0WCUILOwcxZ6N2
umBq62nrSi2cxkIV3bJpHhi6vLadEPixunOU52pizpSJ55+c2LCVStvWxS3OzAAV
nIZjy9PMu0jjUcbCOogPrUjWbU54VTkdvzcnG18wOdiZvBQnwahTx/Pe4cq3/C66
6IhrKmtmrhdbHcMUUy/RneiIVEM7F65I7tLDuhAMUy36QgfNnrL1Dp1yaxBXlV3p
ghnCkMci2lwFhU/1g7mvQ3tJFzKD2PDDjVW2cRPC3jfSHMmFelkr0bpt2EqQGiWj
diZGxAPnm+rTTX6wPEtc4J55oEveEsFznsAPYatZGLwqIPv9HgrBeiEksEigH86J
7AgOTGzb+rZBdhwAdFjVdCN3XH9Fk/c2XVqffe5DUusGVvou+9s2gjZ0AWquNf0p
5CX97gC/nqV6UbihEyb5VziuaG4ebK9xOU+xl/TQnjk48DE8CBIwYPqKBNCQiecm
oEMNW/F4d7YJ/9jMiJDwNART0SXOega5HCZSdPpDIRAL3BlFR4/BxOLpoVXY4Qly
d+v+/zE0zO5AcEVo4XScBxChA442TDv2iIA5ya2gK/jBVnnsgU0nAMc82RQDMu3f
HKye6RmfAi/59/AiGIYe1k72s0erJbuvzS5OXQJ2owQf3L397sQ3TZvwWyBkeGFY
Sw6pfTu7fIKLKh9CRDXfbIwkFYoWpv1WJ98mbXenU0w8T+krwm/q/DgZ0qOEc4qE
V/S+GvPZLGn6aMLK8kyJAAjQM9jhxkeMfN5pxKr4mEumnEow3Gx8xFGMnbf/i1jg
HwFB1GTVrnsWgNjRspR5QmgVwcwrEdit/mt4ilfZkE2iGfCJVJSwYx5nJ40CoIUs
KOm+Vu1WSS0w6VXWfmoo8TeakxhENp8kZkbbAAZwd+hsVwTWEcuxc1sJiDYsyM6V
l0Gm86asc2I9/0zG2UQr1kqRw4Xql/vKzf+nRuqt0YrdZXIV/upzPmypVHoZmrcp
nXiEmam3yTgWEkrnATYG3oyZHrlLHbWO8tiFzW1WruLAjpQyEtXPwevRSQn6NNxJ
HWknRZv8rBampN26FYXO6fveF1tsNOgS4L99mGTrjbTD7nuO3yAg4FkpriEZw+2V
GnwWVeZdZWbcAIeauU2XpnoglggfzBm5Vktub3Y/2PlDTYoOYvJ9mAlhiv9iVPz1
byIsWzaeWm+JWq1QhU6Yzv8DlBfTTfWJD2i9aOqDEqxHGk0jDWMB9GbSvn7UlHUE
S/iNhDB6NtPZPqcuhfmC4uS411BUkEpHJcdrUj3584f18lwmefZ1Imn+fj1BFMpj
IwSbGRl1KctGlU+GgZwuYU/Jy7Sr7Y/+Ax9mksCjyNz9opakrQaM08Bw/pXPEZVk
cUwrd5jteUcZDx4+uEliz9yPuvkztmbzuY6T+WLO7zUPncCJDIHtgsJKcM5lvtgf
DU3HifV5qqtis0Lhh4y8OJgAAR8+cibGdSADcEMtiGnPDQcfg95oUnYvRGjzgMea
H4nxtuaqgJqu52PwlvVImG7VeFSiypTURjggRdThJp0h7RDRXwJyBPzrp5s8BGkj
MLUzqwbZeHe20jrG/whCrKImNVm5qV7oVZm6BeXP1olzY7k8FDcB6UNas5hNLa0Z
eD8pmoDwtIsqhbsh2xTHAwSJMSSTQfq6CaNBpY7GRdvQReCqEVCVWtDwUecQX3Ph
jTM0s5yp3POxpeH/Qv7Yu/g84ULOh8GsUWiAJ+QxjtFkJPJzIYdtTVzGBShH/gC/
01idyMq+F+xtZOjnc4x8q3Gcmyignvn6zWnncEn1FEfdsfQkBU1MBuv789O/6m4j
mDx2Q4wmUi2/aKx0Ce7/Ks9Djt8SBF5hS1BvbR2kCkOQs4xt/3DcxxWEMmi/46Hv
CrvXqKkxZbGZl6Myoa0/GPi59Dgmkvs2+IajWW4TgSh/Z8tRLxte4pW1UvnNKc+X
ktFFXGo3y+RyqiYUZrTfM2ktL3Q/pjAuomAF2hYCCNWSTNL1xsJXFqtIjkELGWSS
5G6uceNDWQDXm5lPeNrmQH7a2DHRQoIaVQM0/HCwlJT63bPU9j9wKL/KB5GlyZN7
QOcPWIWyW6kWCQVGM0vn1FpMzHbSbEwb0cSUeICcylKYhiRp5TzIezY5jUGmRa9a
ybRY2CrBQchCfJ6D80ZksIpUuwQxee2XvklF7SPlKMty30FKWvyA3QqyXYe5RH4M
V2em6D6AggcpwS0lktW6N4ZQ8J8VsppgUD9QCB7Ge98yna88gvsZwWM9Eki6s32m
uU1x72n9p+nlanEcV06x4HEolyuMRmeWFuGdmEXwyJpaPRUSll1LIWF52eZnTgAc
sN/W7Fp5HaiFv/1bqryPLAIIc9wbELfc0BtoukzfPFVUDuLVv5gVFf6I5WtcElQl
30aowmTDdq+WKQguxW45B+A5xXpo18aHDcW+A2bYbQlQCYNoH502+m8zGH2mK9ff
E8hj2pKUEC6CjowGBo4yvM5zu9kBTiiKnWrbp+j2fLdx8A9ejlt4/A18O1R1o4JP
W42RludXmq1VhSaEHr7rgrZ2lO9akUgnXwsCFRpss2OJg4CGlW4RIpvtJCpj/Yip
9n/UmsM8WXGwVc7rKR9HvAUb9/qIdhrR++0hEiSuAFRNH7eK4SwbysosR6qNUEZ/
GqCwoiySV9ZzXr4IYmlITPJ2Eft6tIza23hHrHFzub3BaYl88Xf8WJmgtG2oJnuN
cThHARWkAl+lh8jmjwiBQuLkJr71Q8MXTlUFyk66Rusic26g4DF63RhPh2Vzuk/Y
tQxGoLm4wfcg9UP2WpgYPj/xsAeiU0qK70pMCfgrY/KzL2V4MGc/qd+RshvTo2RE
8wxdJi8jTekAb5Xx7DGi/DZ8QdfF8qfrdeDiLk0OCKCA8oPtkE3X5Dpo6K6206St
iPW8l2VUEkPh9tjN0GpRn6uG9WmOBGWkKU+CjYkO4QBPvl66p6DfNfCWbsd/Ya2f
Xt7H1f/CbcYv6OwL4YEsO82IUa3l58puw6jRijan1+9/T+myohgQ1zB6+Est4Jm9
0Y3+uIN4X9iBg0QPtDcBkijaYOtd4bL9KHM0JPZBx3aqnSPMtY0PTDtDbx0UJmoM
WRjwn99D14qoqnMCrDX6mjxx3I1FxKnle94SYIx0DFM5nOGlBpIu/Rp5Pmmh+X09
I5xaQh2YoKa4JmVoKcN6LZDStIbQzNHN9qkMIfgtegLxbldTvX/GeG0NO3pt0uq3
HUtaSXV4WnarIG5upG+tOLVJGyc8zchKkx0Ldkb+YGfDiLKOH0lcXyurdfbvyEwZ
bgrYbiPAqrN2xrronSc5cp1GjSZlra1x1c8AQfRqq/nAf0z5RR/Dl02iaMIlasrH
ujVeWvu9MWe8CvU+15WNs26sFCp4FnWzp2eN4aEeNE+a0KzkSlqk/DS4Zn5hUel4
majzthC+x+NqxIqSdhU8KKgq+6/XKOCRQf71D/HSlWowuSUaYOxyX2yCSfCnUvM1
WNbn/QN7xqxOkr/5xMSmAam3HHjXWASKwFIRMD+CD8z1fkbqxlvFbgDv5pD6gK3z
Hy/lvUFLrflZkzlvFSxc1nYxTHaIAy8uYlpYf1eQ6fgdnXBtEhtQw778gmV70MDT
qVOyuNpvKVRKhmRECJtkHNaS0VdiNeTLkXzSUPUeasovrppUDcA6WTTbwsm5He+e
wZWKuTSauBl/LXWve6ucC2bStIVjVx0ll00WnF7qen7JJgQxyPcaACuqfSHOp+2m
Dy2dNGejqJcfmThzRd62MsWSimo2jNf6Cozlvlti772TL/6FPnHOjWkLkjOegLG1
Wg5dx5ZvzHLL+E/wWgwIL+Rwfgw1fSlay9m24ceI8yg3xlsA/HJwmSpqCsUUuf5U
VKl0cEZLHtSYHVh2V9BG0Nvi0YL5OO4Wn6zGWCDWo48RXn+U03r53WyE1lXgT9kg
eteHZDVzYOAVufXVvsyBTUm5MocqUkrmNBE2XqsP6ZZN+zZC8gTNko8MF7Ulkd40
hhqIgnjwIlIFJWHppFS74kEUQmlCmv7rrMmRn8C6bTs6Hn5W1EsLL6sBF7VcsgF4
oQ4ZxusrjDYvgVAG+qrxbI7N/VcV/KFX7ltbhk8fGyJQrfs2jOYaTZrbc5p/4lFn
Q+nIeGZkx/DP6ZP0gtXekS7+vpxSQuR60mZmGcc5pOD3Z+TJpMNUX4TR0GspAGHu
GF58+GZb3x9Oofh83uEh7drr3QQ6uCvNTVe3dUVBMXcclocVPETvGiMhFpC7zkIz
ETuDvGHm0CUmFHX2D9hjlw4PlKmrqyxGWfW3+xYUSgVZCapp/h80hvLbFgCxrzDl
NCqlhqze4NgV76CNO2HrbzLhsMb+yLvQJb6FENJLh1Ikc89RLBFAPxbju0EUUN9a
s//KErLyw8/iTaTUv76I6ZviwtesyDoJVJhC5KFWvNbEkWIaD2tjoykwEDKmcND0
tTiuDur+IBgeIu+MO1Ul1xjoHoqQfm/rfJSGBbf6OiTivXUm8x6WrdwyPbsCxlBU
4lSvzgVV6Wg5/dj1NEkJ6K2JHfRjdFbgvssMQA35pXCZCAlKlwJRbF338CLzD1m+
Me//NmescUkZStXGenMISeudPicyPgENbP2tP3W5JpggQ+AxQWaFqEoLPYibU28a
U9q6ZboFPSzQ6RO0PK9FdnIIYTgwnn+lOh59vSlpwKdn4hGNVSq5+Kl17afOMYNR
usB5qKz0k4gx0iEprWUd7zZXu4+nuslKc/DOhOYtuObyGeejUhi67cH7Fa2aGXLU
GsZxK9hdmRvWjjKB3mPVeP0KTwKI1VnjPpJEUh2XA83GC1H2YVUb8HVHQnfEilYz
0lnFIXie650Qyxu2sE8aM1F8kGhSzjSX9ia+Yw6LEn8qaX2TBmUZZjOmTHa9hNcE
/qk6hb+Xo6oKeXtagOQ6iv/jL2X+V8GArr9AAaAJAJUoQYEwj0L3nPa7lE5thg6X
Swin5k3ZtoA1HF8l2F9BIc1eZNjbrtvmIQFBu84GlypXTrw6cII/DCPB13o3Clxt
jFq08hSn7rQsI1sGUpV/gvBBJLYxMjvgZsHCbOoeJhlO8c+r//k+QSJyNmNhZ8h2
bTIL+zIFvftsNuV/j81u5XguZJ/0wQKY90VkzNF7zbVR+dcjNlbK5+NzRa0eWqA7
clwKwLKlYEXQ5oXZkZxq38nY83Ix0iLr0Zb9F4f9Hzyx5ce7AsfdS1EAHjy/TNZB
5FKn06kRW5Q4QAq69/lFTU2NTZIgclyjrkPbR904HR9nDeAfx4nG9vH3hv59t2W2
hVy7jtPRI/zRZbtJUcAMDLeLQjMxoGDaYmrab1LO9dWv5+Apb3QllfojP49vSDok
zBrmMHAxbHDy4vdfU9pOmRvLizanOJHOCgKkaEf4bEUz1MZ9mNL/qAa4xHvIsBJd
tIB/FJraTeyWlX+yT64WHt1E0F6h34swFSzJ6VXg+faEzNG+pgKXcy+WvJPVKNFW
8xSa5ts9l+tQDqQx2BRCvBF7HmmeDeUgpar5WytV8z9VKb9ZuD33iTYe2tjPZHxP
qXMwJrhnaynE7nsL5/Nz4uMQh0eBExtT8Y+HddJ6IZrRRMMmyRmLXtzBjqb5hTXG
wzOnIRNdfhCyv3A/YTShZwAmFN9qid91yeWYcdjJuJm2/S5BiNf705V5RJaoRci/
zu8pOS0r/NfILC+JqKigCee3xQ4RKADprc1GPat2MWcw4XTwS4/yT1s0mxyVk3cM
C8yijELsTs3eLPxqgmjmXicuGpmKsHBEshBeWLv+rD2AGFxV29OWHzAqE1bodbWm
zPOjNN5aDrTOSBS66eXHjRvENf02WufIq5TgtS/lnGZMwLULSVCitvyRNk5uykDb
YgLoG4n8vUeGofZhAR6/9KiFp4MosUDv19U7l4FQKGE5JXrOmFMkSNB8piN9lu2d
ptD3Dg9Gl2J1a37MN4gwT0LI3DqBiZrOeaflxr6iZ9ERo8uXIUWzqs60Wmk/AxA2
Y12qibid1ZBpTtsQQI1GiOjD5zo9bZ/ZpfyQaqzGM8CTSMfwGoYMT73qsE0ulgmA
2CBOS+vwmDkmdzGPik6kAWTvTBkMgIovsBUFE+G4HQprtJ4iMnCS1yfwWqq66qbI
x5S3BVuWjbKwTjP3eI8FxLzE3nq9Pyih+SoJ1a6KJzu8SOj9nMHKdMMmVOy+Icdr
iIU3J7/IzDgqjk1aXcAdNevlBUmGl/1YpqMlgIUJ0dcaKyQqgUMWpLyAHS19F/Iz
IeW5xD8aIP8dy4p6PtCNpTRHTRrlXAk+YKKjmEhTsE2pBesybdFOgXGJdSxluqNG
txwsuLoXuJMbwqsAUC5YiGqWYsAvLwwLlys++Q1rlmN8XnzjQ6dnlvdiJGJ4LevS
w/uNppC6ef9Rf1hSaW43T4pCPchZk2/T/TO6Dni3VJbHNEoTbg8CZBaoBp1CdaZ/
iSQi0xQ7bOxNcnCUdC+i1+BepgFtu5O/xzfI+AsM3WZDu9EgPce5HYh5hRiZ43/1
nm/aKrtVoSaYzQ2cy2aJG+BOA5dB7LNNPwzE3bLgbxMYZjNdP9SLXFx37Ui7tiED
QprZ/yBUjQGXv2fKIrqRLudfXI67EelhnupnIn/yL93xaH0WHbLxM6EQ7h/+FCKW
mJ/fIv/EZBCmwm2DFBKd/0yZklaWv9oyZdRAxRLnrT+4dfRcsUlLvNN9EfagYMnw
6we9xM5m7PgC1P5LN9oPqzyD0Ios+EIq6ncoM3AJDPbvNnf5GtdUFGuWtwlVgde1
A2AsNJ+w2I1Qa3FfnkVV2ytFDCZFI3OjsBADdK+SRx2co9XjudOsZV3bimlJspyJ
Gn5LfYkB2OF7tVTMaE5zrnYcLDGvO0kxEFXKdPabOZiNCgOmlg826Jq/lzwwFBxT
NgKvMXfKHtSVlLff76tKf5CRkUkEmI8vmmv+31NeewJ37vaWdbJnXI2XaK0+n3c6
0t+gYVQDozWVtIlnHoCC2WBHhoWBvPj1XkvRdcQKOsS3PVLV8n4xObhn1RnqEofy
WjqBW0I4QoONAAIHm7agujkWqEql8a+QR1hg3Tc/8e2zclj49Yq18CBdeuNXfhTt
AYpPNMgAzB38YWLFte3qDIa/T0EuBMa9BpHQGjJEAz5wJVSZGzaG8aXe15XKyCGl
Er1XFzv3vDZlYG3j4yujG/R0W396Tk4IabX6l5k7ghGYaf0slfUDb8EBv6CY0/d1
DoZgO+J6wuvV0Yp/0y87l3z44BwTAjLGUQ/brUoLgBewxfpuT6A8aJ4BhpBTFo1n
gxv/kN+rqOT0eUHd/3j8yjNwgDxHXpSzwZwu/tNPxj53TRwgT531yPVR+NE/uzXv
0pEEo5LZlNEw+AiYB64M5YyKdZQ/4KONSE80iv/w8LdGQ5YoiCEuH/D92B2eCw0O
WwiDtXrYxX7Z0bdKVyM0VueNjyCPY9/ZQdcVV/Q3R0NPTWfjhuBFC/3povrDvyzM
uPC5t+WSIEM+VO0KlSOzAswppu2XQUpWiBcjT9o4PrzOBGi6D6XbwU0yzGWe9rh+
lH3Pyy8p2Q03UQa7HegspeceskcW3609wGKbvEsWZtLxki6/AoVGwRqfOFWz1oI1
LOuqLwcjMqwh7yeRYlBlnkBT9YeidHORQ6KH5/4N8FoDK19DXSa2WNXrRSWGgQ9f
3QPJKcyr20jcWBDLpuKxsiRz8pNnuFeov2xKLx1hieBR8OtDunf6kLVmeXxZehnn
lC0LL1yr4ggbEEXaSDjpCau4WLzTO0PXPWqeZG/tnD4sgtyl//gWzsHt8qgyWpnL
Iriz8QlnXiFY0r0DryGHql6snUNj3K9mtT09C1jNxZnyWMgX8MkbYfATicOijfyl
dk46kJyNzx5wKKQJxf6mX7z/mv7l+MfXBnwQ/jCud9am4oNSF+TCQTTRgFWYYDhF
8yNco4h/2QpWyV1Wa+wCATs/oy+NUPFDx884z0jDE0nmm5mrb6iXb58AYE6721Xo
GJYutJgkwMXeSIZhfpqED1D3wnEZHDUNxuDUVxHJBeaOTY9ywNA3d4KFLiFapitS
5xp/P0LzWAOQrnQEoZ16OofRuBoH1sS2Qjt2BK16wOkpq9uOhoCvkn2PIjVF5NX/
w8iR+fwXHKrp98FcWe5l734lCTkNcJC2rGiDSYjl7Er8ExWREe/sKpaZMc2tkEnc
ZNrBeUY0cpk9sX4NiCwRFSX4/zO2WgrYwzF9sXS3HgKNQHKMYlQp0EDq8xaxmN4X
xUjjmrUCjdsoUV/cwmzFo8wILOgHD/bD0D/jfbOrO555PP9ykHMA29ZkIUfSIOHP
ZdYU1tV0N3f8J5hruEAhBbyxGWFiSvB5Ee4jAlMoUE0CbUaDtKG7hMPsXEGB0x+b
L8Q2en5KIZQioVmfmgLh+NU2j0BdTvSBsHbbbrbo/0DPLwzUuzr6FJAq7fm48LX8
3Qv9vaIP9nfmxaXkwnUWJwvjGLRMwUYmEXPu8dhNObeJr/0P8lx8O+fKTSMXgSn2
tyMRS97gaSZb4A4o8yD13eFcbbRhpRv/OgobdqkwVqBxCRTZdo8dzjR+nAPPQOVo
oQKhzUZ1MFfK4YHnQhu26ZpdhhMbeINcQ7OKoe7K4ePK1YcAetZEnCsJzwoaNvgM
XAzisvdBl3BpfYDjgJBaF2Ye4eARoVo/DSeeKRwd9I4G9+wXKWRC+y2BduqwQjC7
mn8rhIp+K4Qmdk0uMdHLRpW6AW7ivLY2fL9V9nQ5aYlLjEXDdna7PMbn/MrkHQgo
IZFC8rzsVNWWWpNDQFwftRie2y21ele+HteBaV5DBHyna2dhXcPV99yft6rbglhV
JZVsZzO7hUmpwkUz89vjjYxbXp+ra1sn9sUEyBcB3jtRYMlq0XSflHzvLFgi8ivy
gZSYCstAiMn2BCszm1G9sa/EWtu4ZApngZquk7lKv32XJqO/u5KjPetHdyPdvmHL
O/c+sKjaWPkNig/pe6S7NodQQaZE4ladEFDyFjDVbq4BnBqIDRoD8K6PLaSVm1C1
xZpNWkA9bOSVqixVttxb+XnFU0d9Az0rueM5L1g6TfdhetTRbTAhzxBl/6goCFes
L1t2ivyp9G/wC/ebzCerGz5bjzwGgSAFhfgWbv8mlsAs0dWRQeXbDNO1XaVLv5XL
WXmE94RIKxitmBGasNi0FRf0KOE+5GxELXzXGIYjhjs1SH9jf5oTAcFXhBffkErL
ntiZQc9bb0+y0iZu/YrU1eqH4WuZFQiZFM2Z8/Pgbz6QeZ7FoFUAvEXQtNGBbBvj
X3RjbbzosL96CDmabJdc3F4Art+/qp1Xsoijs0ib89g89HWkQwt9ZOA+LqWM2kBC
F1FE3wy6+oY6RCwoQ5hz4Nl57IhBPjQ56qtgo6tW45eO6du5dBJZUEOJ5RvNyiHl
oczJSynMvckYIs7P+H0ujpklqN9nAW4+oCqpIm26IgMO3WIrhgzIXd78zObG7GAU
o2f9qogdG81tMgYQSkSZEBsP4isJJhAWWuzLXchuAI6HPwrOPRPojW0boPAIu9AE
EgwuHvJ+EdAf8mc4fJ1GZ27QlCub09gMy2Rk+4qBPDSzoH99hz5B7hctsB77uJrF
nEahb/Vgj6Dm4a39jhTFiRD67l80cefGk6XvFdfBFioTt1hwJ/qty1hAJzgP0ili
Uqao9xxzHsRnml1nd838QXIduL2YMoilQ8MBCCZvnGMCKnjoU4AtfjU5RuVxWurj
iHY+/V9p3LF9zy8yl3VfYUXxX5AxvDmzcbt9bmu7QvCid6FfenHzsZpUbllu7d/V
WsgRaXlFF6LOIab2dBha4mz1Cd+19X3R1Eo5Wsbz76yFd36mCuJyZlgNhuIaoRmc
tqgeMq9obXKboqZPVfNXY+GNbB1XMUw3pyiS7iBVPeQGMmZi69vz1Pmm1Cq49sn5
5gFW9ZRHLz/93sfS+rG+VyKZigjKnVn+zEMqkoyn/HxOSyrQ5CzXh6l6MOfq3/4J
43JQ7pvt1MJK+DqHTsS09F19LYsQcGqRyRUILWfyCnHUNB8smrTXWMH/Ik7i23ta
Q18UX/wwrR2dJzLUCFUoSmDR4XrqTTQvbpa5j4+ITFt0OOp9IJtZ0pYhEdblD6FY
rufljlvN5CLiFtaDZ8GoDzzO612DbZoQjqgLy2MZn3pzCBQdGxVMIUw2u3jvqEP8
PRmlqGrOScNz+QR7a1ukRHgUHSvK6rgquvDzUKDHUwPH3ZS7ACgaKCiKTCpH7R1G
T4z4A4zRStHDfY2vDv8Qe70w7CQ3LT/A1tXOrmhgWOb1A8BNeNJDMjGXnzrXL3Ci
k3Y8C6EPe3udMSruPw4nMNNjzm5C67WnuGT08lRetDQiKUf+iFo7MyEPWmfG227S
8o+jibKG8JwMF3xN5UjelTFBm+Gbd2sE5hXEcy4Xgf6hUmErS6LUdfun1Be6zTO7
60hB3SMBH+FF1dpx1zj+drNWSDpoSQpim1lWgd/rZGcvzfJvhLQqn54CEfSiBtA5
9egk30X15kgmMLFIhNa4FSQKVIntHuIPOcgiIWtlymdtDdP67RtMZflIYI4OofLc
fF4P/rfYQ0yxOoSnL3rBDtFWgJxv8e255iADXGMe9HA/jkQBXvSm4C0M8QzxYlQR
vVo1dr5JeFlAWgXck04WVFm5RolQK9HsRPnJ4pLR9B6yHxzkULkgL4hBTGcWzEaV
dEt0O9wyX7aPmCCPRLaOYIlrlU9iea8WFcuBggjb8ZcgDJEMKWXdy3DBQmgvLUcK
1eTlhkzwSj8AtREaQWx/eAixMebMEAqrO6hqJg4THN2/rbN1BahFqLBy4uW0i9x5
d1uUcH8eEKuaPqQJtytVBPDb6jJvj0rrsy5FMRa0HAoHuw9TGrsto3wlkejjLNlb
lfxk4tcgQo7Xmmw9OUIalRnXhrQVbsRjG7wBMTA2WLMwIPd6xPLr3Y+VwBOnMWXI
EWHzFOmHss1CIdcBVdc3msNmeMmmlRgRg6R4bTdi7rTmT6a5OTg64EAx6uAVo7xZ
C/nKfxt9wIluY+ybFfAoqfPjHOuFODXpQu0Ksx80DyQDrxATroO6i01ThqP+3dzE
0MXkqq5LtKE3A/4oDzxC27JE26QUbx4yUYoureXB7yq3rV9CFfIIEukX5BOvKAGy
zZJoTvkCLDmjJWiKWBLLgGPb+LKJxL2xHI0PFTbZAzWsw5o4IzQ4dYkyQQE8p9UI
pNBMamJZ3E9rY61tYlA/q8JHd0vMEcO7pybv9ajlSSNaQxJqsGgZ62CBiD/ppJ2P
roM3rXJ+w8dudK+0nPv4llROwkmVK6Bf9TlBYtgSxC9sR7Y7FD5tfecnjF36tx8X
ZMkeybke7bi3rO5vroBqf8/HBiJGndhsAzn4uOb3gYIQOhFFWgVL9HdSwz0RkH0L
4UAFUtu7gpZZE4jMmsAT0+2ojPyC9p7ZOBi+d8K4OW175Svl8J7ohSmTRsh5d6Gg
omW3QqfBBZE9XM8LL+FWAIUUw6B17HoELrzf9FPf47qdwV7WY8QfK7YPvXgQukoY
uRJkUspgn0fm4JXCA4qlqXI7A1r8q90WUldMyjnUz0oaAf6dAaXyYxkOKmiu9rpF
vGgLTJC8FLdOCqe/FNPzv42X8esuTdSjk+7gSq/8RXXwZ+xx07VvLnpcgDMqt+bg
XCBAicOqn9XHUiNeZhVziu0jbFRq4+tGAgaGQo1cGjbVZ3jW2zd14V/Uk+XEW1mF
a7Y9KcK6KeMIi9i8smSECt0/7doxbMJpldOVRwouI3ANxhjhw54kMFTkQgdRoi2x
FT3wHTT244iQFaXUFTAWpdrtlRyxbdsRWfiRygGHP8F0uP9IrhgPqB6Rs9jJLtNG
cj3xNEoSqKM+kZPp3qaoihCWjjgBDcabr5A99y9TA2Dhx/Aonzx28U2iW5v8avLh
n2j49txJfM52IVyLbyRxSXMsRLXITlaK+80gyIkkHlIWw6ST4WPAtwinsXT2aegC
7qHazox6/Xgw/vFMXy0lHtnAOnC76Xya00Bae0br1Jpjm+WOHg36aJXeYzAjc9+3
5kDJwMWL28BbvkyKoqYGVUvSzesbudNFbyR6h8cIBsSl9pGoWScMm8n9wfUG43Ib
RCTdlBpoCBbH/+TcouEGUhmf6lqUihcjG+EcKM0ZX6zdafTEvB7xhXFlCcTRSfqm
6rq8O5DOccfiFjxte25vvrajNSXx6WyxJLU08JrTk1akpctQ3xDRt7n/rkSPMPkW
pPI1KiFcBYr0aHTzKQmUU2FDej7GiremrzpsDQjYW/gvKH4Yy1Cq64EvnnCyVR5g
3H4FyGGRSpPJdAC66T/C5HGkZPHwKoNa5EM39NbFcYpvojOmk1px60Mpo9MIV8Ig
DXxooGEJq7dmEocMm/vuivc6iIamjFtolKe0ugPWqjQxR5N7qZr9w+oW+cUiMf0K
5xhfZc/K4dRrYWk/7n0V2XVBUv892acM1m7ZfbByb9fp11/uCk9QTKqD9S4OnXE7
4ufW4z1YR7iNbupPy+f7F5vPYB2veSKw5Lgy0LfvvlweeVgpABVX/AuGPYvEu1Dg
MMcANTolfloFn8LcMFKNA5nmujOlOKI86RtJl6Sdbr2MQUbhEdpud2QEUwlo+rpT
9E1Blccsq06qsHcnLeJLQrFg4c+XP/x5Gbm0zDRUILN2BbNzHxegki++rbbSYdYq
KDHPQbvtZMqYnfnfvMNAGbzIp5iHnEjOD+rD1EpC8fSkWCBKU/tvTrXtnvVJPGb6
jSDD+uHgiXTNEC1PccNI92rBnWnuFnSo+p5qr28umpvRn0ZZEXjmRRrj/lk3cmgg
V8Ji/p3oIzpWid7JiRDb9iXxVXdczN9vVXU0gbpturO0r2lnCimMcCt68Ynuxvoy
aZOGWzSsYI2czOBwnBEuiM1gGHYYI3YDYAlofJvbRoJ9/agbJWhUq1siZckE4CQS
J1/AlBUpLiM9LjpD0cyNDeqL8vft3xAgQ1RRZilMx4qYRKFtO0N3uvW1XLSUT/4+
9f62jNbeoxwQexoGgcXESDq0JbVvAMxENG3JIk7uIcS5Y5pwVfzUBOOL+fD6ImQo
l+Vo753Hp4KxMRdTu+hdJrgN3IOhJYsCq3RXAqdmd51kJicwwsYS4S4A0kjeZN7p
8zxRfvC3l3TVFb2/3L7tsCn4qk3+pFhZH7tVHZ30F76EzC6GDNnJETnrlx/kwt59
kojX49QZgbq2WLkqF73pWAzZ3/FsCctlq16C2/urE7sjHP0X1TCHI3c5tXw6zPM5
sTA8Fpg4FqKSvHo0U/H5PK9hk3WwNdG1/AgwU7K239QCt2706V5riKo4D4XFXOPS
/pq0T6i+E6J5k7Buptrgf/2SG4AgnSO18PJN1N5TshtHgfDOObDPOoVNbEjBSolz
UV0JwC2dZMo/ImDa2FpZPRacurBdKAff2DkzuW8gAk3mL/6JA3J6IEDbYhsSL7lD
YrUL2Vs/5UEoeH2dLqDsIfCCfV5UloOXuSYc/10Tz2vRE4iWibhLjOAROkczLKX5
sASCzaxeeLyfR9p9ZGNVI2KVm3LrW/4cuB+NWGDf+3lXbWI01Y+SwP0NFRnsiNjx
N0bib3hhR/+sP8lNWIsl/lOM4NgG9bgfqwPiaudHKic66Rb5N4071Ro9mNQDq7FK
Q/0bVql8FI4YLolKsD7l07Ios7NMh0oIuKuPfSgfEuAuEUI+TmpO+/UCPxOwFrbY
2Won2a7cm1FvJcTzhO1vkmAjfu0dkDDUwNfeKkHWN8Z1ggUEwDRB2Gp1qlGSFI6z
j6PhGQgGbVR/Gfwt6nPjrEn9Q4R6g2bhezcJYk4qnTSfZRPfgiC6DnQgdPH8pUu7
oganTqeXh7dgI8vVver4IMJBsSDKe9xV5DBYEGRHAhsownTbhm5RmA6H8jGCYt7m
r4NkkuiBGt1IRLuscG4pAq2t6R+qRVubi4Kp7utC3WPJIlWnFzB5IV/xGWcwMCVm
EbhiB4cJn2xpXVvYAz7O93BNtofRXvYoTi4PGLmZKaxE5pG83WIknMN7cDBdWP4E
jJmpOTOVmNJc/Ov0fF3XeX1t7kYEuoWOZCJSgBQWbNlzu0N3pfXKdGIG3duwHgJ1
heFu5EuuDGSByaVhI/Dn88/GTMESau94MRsEc9Y+MxSlgiaR6ytDoZQvNfM1IG+p
rzvchjxv3LnxtCQOIvLiJ2QMBcrdpYba8KzdWn6vgzdEFKQMCsZ3ZgiES7Ui13sP
IZ13+LolZ0Oe+kNTqLEANV68wBYJvG9HJbFXbwYF8V2pteXQ7rw3b+QaOrUFDoR6
JDWiL4i0zi68b+1Th96RqfG9ycqIk6evQx62Ekrezt9u4rSvGOfrguXodUmhdVPU
/Di8QvyFIJ7FkAQfHB36fsSIj1fPkvYiG0x0DPTDbJACOr+C6r1WQ2PWKOYPl4Sh
PPMr1QaknyoAvqqLIN8+8F9CQ6oepMo2uDiD08eWwReKsmtSgd4/MUeCWOo9LMGy
62YwsZyyB2C4QP/eOd3Y4q9rv/8+YJ1F91/p1JNk9UHGUC622TBxc8S+S7gus2ox
cWG8CAhQUBTWBbq+I3K+AYcSgHQOKTZKGf86eclODnA5lrIqWzKHQItTzi3m/4ID
hLnxYBIj2guVEhsrgkO82LN85jEcVcdf/Aaq+DQ4F15++qRhlc4VcCXmNu0z3WMM
ARaYkMLl/LMjptaBNLidtjU7wfx4x/SGn6NnFv0q8gsbL+Zh9DOvWZuhRgWtHkR8
UNkGkkrECR8M9s+lxO7zANoPOAGmOJuWNNmdLtGD771eycQPs2sZYll1u08OT+Y8
fGrM4M2EwukrSL9/VkTyAXjW7bLoauN8nLBgukeyWiwsEFiSGbfbIivWjg52n9s5
QNDXnralJSHpQELucqaOMiZ9VAjg8M/GslYWut7F3+85P9KfA5ncPSW15IiPhnue
0lxNyxqMEmLC3x0OQrzB0+RDOk4oprcy17YvytN0MHfkWnJ8AIfyO7vleXMhrDXs
DcIZQQDdcX2FYF3fFomeqlSUNdEfuNizFdhYJgnbk2GyxwihIjJgjWxB1kjZ29QF
AwafdvML+u4CU1AaYxeTFSSuv6qn0zuR/PkHYP+gqsjp/HmIaxC+Ym9UcrssewO2
bnoIM2xsrNMFzMGhURMOjDHokpqoEvfoL3XxeX8n0OuEEU/SrZscDx3NrcaPP+Ww
uw9I/+orebXPnW0JL4X5bdfGPCDP+N/7B1bwnAxK9YlgKUn5yxYieZLX3ODH3P/g
avKhU1lFbAduCZN6LBNpmRVumpMFBph2tjw3cFKcoN/YedRxpvuDIgJkkUI1jO7V
mEdKGnY7Qenu36BDFbWXvNQPmLDxQ3qQAGad1lnO95w2UZps+4Jxuv/WAofpoken
ySQN+e9QRkDRpzeg1urNgEOZ1PL8CE0LgDYYnXabDLM/s2NNaaDqmAgPNmScaYgJ
SN7YLRPh9+JCuM2YpgTE0Nn0MUTd1K+ahsBWhKB1JIdcHnJm/sihdrfNE08ZoscT
uNrF8IAOwlCCKoZSaOp3SINT+sqLmes3HAE7s+1lMjtXgRGfPCh3Ie5HwdlKf9kO
cKSqBujo1JojPr2ASsUuol3ms+1Inv9CyrDou+RRF2NdGO/O9quVGJu8FxQSmjjq
ZIpGy/W/+rUY3BM5newt+26E9w6YPbM22ysErEyoLHtgf0lbOql0hQfeiFMSPLz5
PtLrTy1yiT2/Crc6zgmhG6rimJKr1lMhd2VB5rMyJlJm/jnVXgxg/PnwTLEVxeuC
Aux0tfjClBzU6j0obAAWlZNMgAMiWUGQ0ZrwFlQSdpKH0hri23pCRL+WxK4B1mkr
C5n7lPf4G8ROER6GvS+DvC13Esv61YMzS5rMIhG7AgeugqHdgLzDqkILXS8GwT+7
dAUgVEjQgxYxuL+zwcGkGekHAGG4wOo78MBeeIK33FfdOs8TrP4mN5K7B2tAsVLY
vE7Jx7HF9ZM0xLXHXHX30the4LEoDB2L+xdqeSRGpWP8kpXpvu6HCcJGHf4ueszE
FR9/TPqgb21VLg5sStTNfrb1rnTUPuCqOFrt/rtH/EBfIRZ7YMedKT3XwNROMNNm
ETN6pd/hMk6jU0zqL7mvTXX1/ktyq2CqDvCt392j/yElqKtXnp2NPPP387yMSM5/
xRIPWcLXxNZfsdD8On1+z5FEZE+RxtJ/1SWI7oayReZvKQ9ZCPJel3kKaOnXNJ64
fF6nxZgbrbE1XZ/zxzEvprzGb+2c0suFbBrHOAAr7z7/ek7IDEV2uk1hepTv3AIQ
hpwELh3xOjwVmUqgsW1YgZ8XMW8DHTe5hDw+uc0cE2rWiVGlZuc9u7ILc5QxmHYz
kxv8fuLSGbI9SoXX3aXR3mfYEfPz3fqLRnF+E0n8oEXq+Z+Se9iAhnQfWmILx0dA
Y/3p3Ywh2djSgD8PwloOz8AQlMBJwwa9pq2fNxNkPOhENiMTHHE8sKXZMTbKYILk
u1px9bGdbMbKa5APEWlhMRpDsM8QpSZuprCjOA7j5IGK5np0CYx/t3uSANdOdQlq
6u+5AViNvacniwTJtnytiZo8UNcKcczQNBXvQGVF8nrdZPXtkKjigOhok8L2YXLc
VVWYaXzQgY7/84H4q7qZY7bteSkwcZniUellS9B+pact0WiBjMJ9hk0HSFDyPAjU
v9szpoXhl0pbWnUE+1FbU1jhb1kO1y7ooy+gV231lpIQha0M6tucn5Xcd8qhQrek
Y1MCavyP0to2ftGF1nM3xAb7/CesCoO+UVQKOIW6BPamiEntVk+WSvTwjq4cfFfm
rID3PgPc2iOUrIZoYVvpzyOepeKSrqNdpxQ4KFQoI4ds6aDsjkEk7jdWc/qhlVkk
4KArohEDI1F03RfkjfTCKlgCxjk7j6USiaril/N5vDm0cp49j12acqXVjMNo7+oa
jUCipOK7tweJhP0P9byyoN5s2nV02CtjBGXurUT1pZezb5m9g7DOt+hm391sR3NE
onTiOfiMnMIgyl0LOYajYpeU0OXUGbqNOvzAHszyFmGFZCBWJcVGQHdyhTU/fxjg
L4QuhRjd74xsvKhrpQx09j7uUxbm0xbwjjEdUqA4cWWrKp4xay8Yg/h2pUTj69Vo
A0asX9+1e9JdNEj/TB+1F0Prhvf5APe+dVDo3FmL7hYeTeaZpWxzXZ15/uZax8sg
y/yL82sbShdJwxcja9RODHvONqgI06Ln38kM9ONtJtKTkS5BJA6NrWkUE5hlmlKg
bZ7+IfCkvVPyYhBw2nniU/kMRGXVGMJL6GNgi2EqsE6JaGQUlivdyycUZ010yWMJ
+W9KSdPm9me3hIvOYY6HEdStWItWbag0Ty26sCzqRHr0DQYH8TDu1ZXSJbOpYyZv
4JG8dRfw0m1nDW5iaEW2olDjYNRvnW2XL3OIOXp/XjPgfsmrqMRJL/hMaSirNPa3
pjJeHnL/HL9H66ntzdSlr54wpU3ZFLwpf3gUiN5xnQbKgyVnzQFVzpsYdCCSZuRc
YHGXkG1ouooXakdh7MGcwFcnq1laPuNQpBnzEG7kcBFXH0ZI/g3gedYgPe6Xx5Hk
toROQnR/NvTb2lz14wn6C1Naut5qIEAxnnmvo8lRzrg2l/4DXLJHFPxctpyWZPoe
MP3ZLOVG8yzJ5WbelunWUuOhrxC6bRH53QWlA6zuwV955sZFGCPHiXNJgbzmQ7HR
61NbOvwKPFZ0d2vpEExWZed6cuJZnYISHTLG0scKXJgcfgK9tbkKWouD6Co8MqMw
W+49cG9+iwgJjVzlTVKjv7PNfRj6u2rmnznIVcIeeXatzvSAidDtl1+vvnN3ohl1
fR3fPfFrcBuazzEMv9FWGODxmB2l2IU8cAjTq0nVJ7y+p6ieauyUSY4Vv+eCqKcz
FtG1q+NPhFO/jS6mfJ6OA9QYoZL0kOr8VWFaTdQPJpox4f6iFfVeBv676Uvfrk6V
WpdltUUSDDOgOFal3JtKafcet1OndrropOcfWl5RlpZ8JN/X0k/BiChRc+SC9/CL
AjTzq/cwtFXWDUoilo21OVduu7AA52hzhRDG52MxCdI7QZ99Dnff99X/OR6WwJJv
A/Lj+RMY4O0Kr47j4K+VI1ghBO6okOjPrvIoHA/pGqof6x+tr+hg4TXPWR0IOS57
xMgx9EEHQWuPeYbGPXkpf/Cen2b907Xidr2vPnofqAHAMi8qaSigLrfskwKUn4wM
cZK8CxCrb5gOGVni5ICJJJPDv6Y7SiWZXAZCh8/aV/Hjc3Aws1E/IpBYDMoxl6dQ
Gugm5JYHT7M5M0dp4tTCHvIS9/vr1dAHSSTZ25SexXfaVijqlS2GYRpvD7ytNVhJ
dWryF+4SgSfD+kAo7fHVWD0oq4vuzkvzWg0wzHN9mvmvQJIPWUYV5doGvP7yZQqC
x/+rNSQq+jYDtq9pLCu3hlqxUxn7w9DPvsafgmOqM90QynGtgTo8RhzqEG50qnH1
GI98huLU2ZgMs6eUyrI7jvJNQVQMbr0h9NiRMOgAy0zaeU8+5H5Zyc+9o2ycfkCp
2sW/V/Xx2sW2aJC6+0QDEGUlxhMDToLTZ4tAEFrVPLmNCwUSIuhSNcvXvgy1c+Hx
bllKosrBZAIZC2a/Z8fI2LhOafJAYDgJFK9eKwkwE3tWBugDbSUwTojaUpsgwRII
dy4LbwO+obSgMf/neDd3rIxQat1smzqeXMCswOSv/+noB1PAgusQ8fMf2s7lOq2z
KupwpDGJn8QNFzdYDABmHFT5oQXEwMIWdo31WAOB0Gz+9QCDwsJnYwH105B3jg7i
24/S0yOyqAhAyvSh8E+u1o2UzUIYG2NEt78v3pj3HDpP29E6aRQQL4qdtq9j7s4w
zP6jOZLbf19HTCdIrv+uFhOtGaLkU8aZVqAtVC3EaAd6zeK79kMm++91Uy4DZhev
cKsdC5lR/ePeQPFRB9ZkARmZBOlh1HTrzvgWqCiRATDIqCGyHyDs9WTIOrAR26qs
TNhjfoWbegoD7pSsd/EhvDunvFxpJZCdShEUv8nqwb/WeAMHvyX6dMB+to1bmeuj
/kGW88KwUomHf+cqPPxPeYrJAROzPugmNeOQX9GZK6JrPKTxTiiFlI1DIe7h2Fk5
1p8JtBvB2ovaxT70ImhXrw5L9mwdVkrQspBftrgN7M5XyDZxuaGjUQrV3ADBSCUH
LYdlbzM96tTt6cK0EgYHUl7xzolDGKhpf61FV94Tj7G0cGpLrGGUg5x8sdt09g52
ny9MaOTZ8OicOjapCwqNmiWQtmG5MDOaO2Gjhnal4gMmrq3LN7hYzvbTuwL6hfEO
P8P8b8IWy+/81WvpzJaW1wehCgo9FUlLMReUEGlOpAelx1aw/PFxxtgB5E+P8BGE
AW0LO2lTStOkKCUDh9AbWEX/dtQUoqQ+iB46i268vF5QK9SUUjFDpswSaNV9Efoz
MMGzGhArxHKu+I+IIyOKTLGG8J7FNXTSn7dK7jjsJ1rQf+eX0O5f1NB1fR/hqqgW
Fj387PCDer7wrUk6129r+5hOE30HPTZHWHQy9ECigBTOcxiBRAMYjMBNZXtGHm9S
VSGTXUOhCBGREt+dI3hT+GSdlelCr72k33hLt9Qk9qY/ApEa9c+7Ng9aIrFXNWg2
+Y8tspFfDPwhA4VRWsEUYlBCwBpvgzmibV7hw6F0KXuEWPZTADn3SmvP8x/nDnp8
W9T1CF+TXTxrK6gaoDZaf1YMCbvnXcBOjighldBNqVgG1G4PUHUQZ7OID3/0GH49
xXULrJ3JPeS1HziqckeYTQfKjLqmm2mXI5tS28GzzhhJLAYpPntmRt0xpxJX8H5Y
ySFLzTQqRACFINdxVPo5SVrgyP3Bm1SHOa7wqOv+xEmBu+sGGw1pU3fxvqmb5Srl
1BA+ukp03yosA9WkiMDIOFcbIhX60iYk49Bj1CpAoAsx7usIiAG9Z6H0XztEXsRd
+le19Pz6LmQ3tLuQ3a7umyVX/EFvd33MBaR/FssnJ7XAQl66ZYOuDsifXw3Acw3O
zzWzEkHcCa9NVy4Mf7Y7mPJtLdr7gToLJwzEQPyYbIDSWz6zMlnVSaZCSFB+AAem
UOai2I+vVElV/w68QFt0jdHuQSxPkSfbFKxAahWrZaCgwrmihMqgEuAg/KzebPrl
3Ob7azH82ApgfeuorbgJ9/zobOCS3VSq4W0IlYinIdE4neBuENNaPgzjifNyKy+n
H9tejsMbFcGBY2jvW3tZZv7KLJImmFR4CLUPef8x9NzdTgRO5L0BDg39a5CRnx7S
X0uZHjLVhlWNenwb6XIMJt2vwNb7WpFyyzxKLM8bsTfZzINqD7+KOR8GsTbAN/Kw
5yASdLzIcVgwn0kDQ/U2Zoe5+Am2smoG2LXQ1aJ919Z8BOmUgcspw/ZIxd+vJcEU
yHh2naIapmOjzGxcfVXiMJb+MMJXjK8I+N2RNZWCbGqgqJaljMhT40XJjfuW5uYg
bLZGQ5zB/HJu23TgMiZJMF+DuA1GzsXSA/UlnpGgeNnusELUEbmZR7psaDxSfUpE
oJaLVN10BA46VgoTQfssuRESsw94qZQraHbyOFiW1cuWg8et5KGIeGQvd8usYR1K
2lTdqoJQn5BJ9DnzvPtn8S5Tv6EHMAcVy4SaH2VTWgYN9vDmtBLvwDp++DXMTCsr
2ssm72TtkgYRFTK31FRS42aqx4g1jwk8r4ZAPArqWJ1+y1YgrVaY1D1Uc14gZ0go
qLocPlGbOCzfICNEgKeQQhjhAfCbGspAZr2K1DsRnCztUiUBrJ4tgh4zJiepnOHo
ndCbayBH+T+NK70gI/rzYlCm4nTbrhtgcm9aATDlFulIsU/6F3U3HOR7ptAy/w67
4jIVs6e3eJYnOP+tFN7D3zLnrBM9vSI8bAAVgfM4ggUAaFaUQpoOkaxiLHpvx8xE
eCcp5wvLVUZuvYSHfkHTYuEszBWn/OXQqkh44vhAPsomFHoKD1+Z60HniJb9cY08
eLFMu33+dRhngk+n3/FsO6rFGFliFwiDYYfaBKXWMjYysNlxlzJDLGBHYtJFE7/k
Hz8iAVSYalzsCy4qYEXFWFFS1NdVw+pQqx10LGUq1/iNUlZZ+tLsJmRl94B+xScT
Pbix/8ld1rsVYPkH3wQAni6G4lO8qcj0cdEvHKqdSuDseUN4ABg0J8hFyUTkLGIO
DFUr610ngTTINlrZMjPcRvqb2Q9/lS2sGnuPI6uOWt6M5pYIKuVMUgffkh8wA/li
MKpHPUYxrBRaoGMhAKGrE/UyZ942fzmwUC3KXlAZ8ndiUm9m3caam2dA4RQV27yY
rR5f9xivoJr9RqKDeNgJLhPh52SObjqtL6kel89n6EVZHNShKYzeUsoppDSGNx5r
SQyLYhgoO28hWBugavKTYlR4TSHAQj9aCmuLpwEzlZIqY2A8qlH+/+XnWd2DV5i1
NOLT+JSjut0bDeYfpQ/Tf5to5GM8sE3t96rbY+qyQp5/DOMcbULQ4uJrf5E+Q0mK
7KDdRHCgd5TfvhiUqtfKKbVpGVJut3O9ztDArTP/h1UsILJ7pNEEW+ZUKgEBbA9C
TCbXAecARabyo60AtRr/7rjge2ulKdK2etl3bIlMDsipmhbPLtmvr8O9nPeckMb0
wsQ6BXW+rODJR/qTjq3HFAP6MvrISKC+/jFIkxV4k+A42XO5JBnBXQLTR2wGmH6A
4LciTsSRQTK5YayFoetueTDs565U8DeHLJZJORu2+L+uUu6aO6SklLzUwDTqd+kZ
yxsCh1YfqnVIYaDyVvBEUPKs3VfJS9Icm8+XSBd5jwvexar5lQ158Xv75o6TObHK
vr0b4IaCvhdEYT72pdma38GCqfIDMu5gik9aOvC27ieZgLV3xrR4EsmTmZq+QUkx
F3wBLWiI2XcdyvgGw2yMSkWViMWjzyRXNYcWPF3J9jtJYgWnWJ+T1t5SmJ8z5HKv
1wYbsz+OP9hORZ8O9HjPgIOexwntmJqr0inCZmlpMxyBb99JZzEfuS6BKj+zwLpv
US48g+EyUKudRTndHpuPIKrpw88qQqE8ZYr/Ny7rBijT37MUeeMrog74P+NzipA3
BDvctcM5b2MfLqdi2ty3QwBnlvRKUI4XWA6hZcYc+3F3tQSm0+Pm/XFOJdy4qCW0
MOsqczIwRRkiruFonxDovwOcjyXdw8Zq8UGLRU3Z31o3kfnIyKfgmyW0LEoHMRkn
x8kjUhWLWg3pyz0bvQuSmvF7YZ6zc6hHXY8nT1at1waSWWQyWzmeq/uTFruOhzUM
AoCTCCgzUF77EvYge6IUiRiJL+DPU+PuIfXDwg45so6q1JZSFAcfufJmZ9rfDfIl
jXDIFZU/i3wLCsun8halIv/CFhmgPmp2O7i+/T5DkxV0Pa6rn2LGSo6lhLM5o/XA
IrPTxeqg29v+17JvBj+y9bqoa+U4yox4M6GxKn95zWSzhe+KLYGM34KIrHB3affJ
xe0vvRYaRviz4lgOsx8/K530sVonSKQyaUVL1wdR6hjOfPPzg9SK6YHimOmbJ6w6
rlUTA7fNKobnBG7sK8dkgFY9fL4C8aEDHYqE2ZBtaLqRgQwDfcKc0VBEt/G6BFj5
kGbhpnEAcNnulpioFmXHykIS7OtpReCGfkclO+XKm99/b8eDdBLfyx6SwqzLZ5uv
tlfiDPdJz6TDLDSO84ea1vGppjASUrB0Lfbkd6PGED8f2qnKvX76UkCxW/ZWct9b
6wum7hghT575A+NGgJDK+fLEPo/somQCdYLws5KsWaG61nGwA1Cuc2pikAFyAA0/
TNQax69e6KoKorR+Y7XK7HnCRc6hKC6yEzhWYjVkAglI+cAMBLNzXXRF9jEaJqpT
ipG84sEozbhGXnfZExmumKu58FvRh0HBUpGfspBoKLpOsSOMfFoPgu2Ri0zykkT3
Q247+f6/3E92hniMeG0d17PO5zKy0Xpdk1JkkwY+9g5Q/nuQZ5xMzh3iCmRHT/hx
5L+to51QlP5DsqECqtMebAS0VFW1oHopEGgiVlyMoh+0/FHn+1d+IQu6JAArqvsC
xmFD/xqfy75rUzto6xDeSan2YroG6FYg75dWxkmmBFQEIigCCDtgNdr+vSZSQ+u0
QlWc0P15V7/9JrRZjhWKSn4Uhpw9q1Tfay9RUdldH5VtM7E83XCzzdjSI+F/oogH
4e+krbkb3n0PUQfs0n9i7DeeEHtm14hHOgpJMEGACC6OgWkVDdXhnofT2nC7ZFFz
xqc5gR0xGYNmctHVmB8CBQpSKmbARbOv4tl2J9u3YGgfat11O/D/OWR2U+rjFOk3
ZHRo7IESffKg+6UfWiqURKvmo15Wti5cvIJvwN9R1n71Bvkow+DwKQSme7eFcMkG
oHIS9j24+vLa3az3H+FjGZKF9nhPsrw/4HIQkM1mt5p18Rz47WDbA+0izaAQMEf/
rMmCbH+pNgir93kv9+XaFJ5+Bb5Ck/lQCoFjT7+HDdXBpV0abL30SB7qK2rvf/0n
zHxkwH/+3hmPiee1T1xk7wZc3c8IYiyYOXP0p22DL5+4MbQh94weiejoJ12k9eAb
29vrFjrEoAt2z63eBRIQUesAp6/SmAF071iUL0T22aZ/xxBa8SoZ7un/qdpPGSvq
R/7NXJ402qfpoX1B6+Ggv84go5QhBr/eM9V5YkLXck3CoADFTyEWqUrbi8/PFw6k
cyFAu+//ZitZORgpkgN9VXsGS8Zi+JoW5l1fFNcuoD6snF3nUxaPkU1TyUEEZnuq
DTxYYvWcV9WQa4O9wvyH+OSS9yYVOLKmyk2ISs1PyW1j5UmnuWtyVgpiimXKswEl
s7pRAuSr37F/cZxrc+k79XyTZLhGf0686qlS4YejEv+UYkoX7+0QQKS/udxhZyPN
IRuepYxl7S9vgI32VtM0r2tASPGsRfRxjFOZBqK2dMowHhTikKrzTF1+7WKwuC/x
w2hK4B5tY/8r2E3I5j/MZAUneQm+Io58KeHGSk/qZDuXM7QmrESW+wY6VHOcyUeY
GtcJ4YAOEHF8WyPx9qDnZOk9SQ/xb6RRKrnkmw+vjyJLdaolj9ZNrh7YMuJ4PdyG
aHBE1B8iNXMGKbcYH4uYgk7XEiWocV3Cglgl2fU/nqywWrrIyG33qB05qs9XxqSq
4zkUYxNwiJ7F2lh2umVQ/spd/lUGij6eFDgRegTPsz1ukn22mF+8LxeFVkDkaCFX
sEECS83i10VF+WxF4DfhiIYWO/HSg6MCPOzIPju/6zrC/iAUA+y86FKaJlZSXcIX
PVLA9n/priQCS6JVMxuk6jIM94E03X1Skr5IWlxJWTMgCRNgw3UJk2h2AghbYQ6V
BidTUe2o7KGSeV7OAecxwunvFWkH7aAkd6/up49O2zDvQb/6WYqTrgPrfl4Us3fc
4xPbxjZ10SgUmp76tmJ7tnwRYmS85GnS6tnQI0QRu8clGqpQUQdWBAO7vWovU3vN
fV8HNk8Q//vAdmqSJMqVnSlGkpmUGmNY7P/UDwiwFvliRR/VJr7NbDzd9FPp4nT3
LQN9gDFNAXS2erTe6vNP4eC0pnSV56Wo+1wTKcxG/Z2ya0IGqHtpE8JjOiH2IkRW
UfBcSHLG8xZsXqSMQEcj/nLhPdJrPf0Q1qwVa5wmhT1+Xldv+5MXYtfkP7C4Pmre
ZOX5jvBNNfzCTaIV8uPIqBjALa6fr2OQQA9kfKeqnsHZcMvUsAIlchTrBFzuU0Nr
iDRcerSgD6fTKqxZHVYoajpKcbZHEKwIVTx34FJzE55AF4JYzYS15OOpOl8RcT1W
C+v7GPBCsB3Rt/S0Gci2mHeubkFvv6w8I83+DHlYHodFLE/NuLxvbH808/yfbchS
e2o6HV6baQzupG8gyY3GPpZSeqpfM0y2YKgQaXwKlZv2ayI01xFpkr3i4fFqAGv2
d39q1Pj32iBUhfr9b7zA4f/AxwWHMMCXsNw7BawW/xd9uqaOaWcaQ9MVHbqX17CE
+Yb+0+GMJ97WI317MIhYnTHnDZzfuXhLL0mf40x8+PwqXbgIEjx8jNV0p7rl+qX3
9oJIP2BMofnS7JCbUPcg4YqR6B478gZ/BB8qq3W6fjHlUcT/rz8jbmb93jCSJkBi
QH6P8FYMTkFu7njz9cvm+HATSqIyeah59RwZjSPpdTYwH0c9zGqV8C6lxN4/TkHJ
OPlISpQ9wCXWlC43B71ayUjYfXylWR+FysDsU75OpZpSAcvH4TLCYafotCUA2frm
AJCTVPtfbEk9SfWxrYKq32MRjgUodoKSXi+spNRrSg3jWFcbIJXh8oKCZS8EE8X+
p/F+MpH9Z5MSRI1jL1C2dkU6KCn9ZQ3Op/jN8nnhf8YbKFGcSzLbq1NADDeRVZb8
4UKCXFKjkwRemgQXFrGDL4wHS++mlfv8jOrEPq3n+pj3d08tAK2UKJvEc+oAerJb
V2nTCrSScZU89SzFAUX0ylQ3yYU+/nLmr8SdGyh4rfY6o7VOerieG0r2hLDcwjT3
2cqafZVUzr5Me7iTs8PqY0h3bzyKo6kXRUk/ALoczGXO07cMkGRpeOn/KglXpYz4
gKeMisORBfJVEPKMWAVWuo87tAD0nancDmiwtpa/LAgB+1Io/rLOYU0jpq0V8uh8
ioBrYzasSZWIfJJLcEYnQN7wieu9WSiMarSqyqX5Ef+RUoo0e+D8D9yAusZsXI+T
ihZk6ehPKIHu5Tpt8qhxwMdumUP7R6KEc8ba/u8eNUqFDBZrNLXqi9ZFq1h+rxFc
rEfQAAEN4dGw/jSLuetI70OghKkT66OfmmURikoj2M7r9a8Riw4Z4mvseksRRI4T
WX5MbB0NSYWBu7+OEZniByEMe8gzlh4a+PJ5CxeQp6d5fAsVBuFRu1JTCFHuyUcb
Rr6OA6Vka3iOmKrVR5A4TlUJoIapPgkgy5/mLRIzq7+zn657Ol/e+xb5hL3cPbp9
Vh5xSwc38XFS850zmGmdd9yIn8J6ziY3H8ZTKTyJECbJbAYboEZ/EUOZ1GXR58JR
tqvgIA+h6YIxaX2w3vCew4cCN2jpEuG6Jiir4MBfQLuCOIKt6cF5kEDg7bUjmeXV
CUa48bi0/dk0LJH9k/hFolECJA+q2Z69wTp/ueRr4Rfy4Oi00fayk69UC37kXPaw
oYWbK2z5S46UYBnRMO1sDXgK0f28ScSwkOoUau4PWZjEn7cMAwPa1BLwoOEXXa0K
QZWctLCnUZmnHb2B6hJQ1nVQdNoPCniT9cdC1Q+uaF9WOMvw7VmPaKvA8lyACEOA
aA3Ps96scxKyJC0nTxE6GVG0sxqHRMRV3T+BlnsXc8t3QfBb/SnqZgFplmk9MQ2P
mLS5x3SVRljJw7kIma19+nHmVXczXpjyU7RjGrVu76B/cREFFeXaN7ed2aj9bNHU
Oy6LXXvu3JyUdnEQWYzkFMqAdz5ldwi5f39s2Kk46HJbVDZc38Nn2hRaE1inuAsg
0oV4WU/J7SaPITYQRoA/4/U3aC+0XDVoQRNRf5jhHBiS9njyXXNDLOy2kYdjej45
YjUNMn/HoKXbM5v6VJidx47kp9novCwMvaFuSYcW+np5xLlJCfUI9gjxjbaVVuVu
9QBxxKUMzVVplM12qdHwHxV6TRhxYdV+u+9mhalmqaPfeADMXZ2+RE/ya7eJ8OX5
MwDgtPoM+9TPKRCzvi4bLGYPIFOe0fthzdkEnM8YGKhJrEMrx36lEyMDIibHrFjw
DjgiNukNCnRSUUwOe5N4avK+cuuRM9rND1E1jjIiKJGCuwiGuPq5/oBu39ytEZAO
UvxTrM0Dkbc/vlqNm7RIu3mex9OLPJNii2aAWzCbqmO0NSVI3d6/Ys0zeVf6w7bK
GtMCnI3mpQeTdha2MqFUjxbEXYOHFJPt6jOqjIa6sFSJqLcbNkX3+MJyXjxfl5ad
ifHTeDraE3LDkfDtYoWv91XlP/DAokkcwoXkatTcaou21/9sbuuz6BaYWwAJ8IXy
w8T16sqoebVnlxcYij0S31iNp3U5T2JWt9Wjgv209kezDWd3ffCdg4k0HUdS6STt
ldj4Cnbg7X2lNmMVXPWO1EWHPTd5rQN6gfkl8pVUbXZgz5LE0Y0crLSnaMbNUWOS
dkExXqHXJQ084Uv+hHVxsD3aStAHlxcrey50FP0ThivDNH/McDgLTCbhQ2MDsiwe
jPSODc/joMg1MRwR754TCept2HQnSduI1cL5xTZ6nrgdIWVKJtzwUbyQchz7011i
3CmBoExWVcptqd2d/Z6Mc8sahr4AafVYqdELSdV5F7v5jGNtkHHUxrv9m+cAq4ow
p2TDe6kPjJvsGeTDHWlrlHa/+gslPIKeOqZM5OHIYOjkYlaPdCtrzbiqUSGcH0xI
nu7DXZwAVwoPwoS+mHA/nud6INJnNb0ALLVk7NQSanuylEotJ3oQxCkrduO1MHjR
7ITWvXL1laB+O0LWcc0LtU/w3zj8qmFv8XBrQ0QJNHEjyCWrQKXEK2gRggbfKQUh
5W4KfwbD23avQHUTDy6wVpR9ajlDjqQBdO5ZJ6SIbxHwCDbBEz6RdCtGElsULeiO
6RtxVcAASncu2vTO230NRxH205TLoIJP4fP3h+R5OZ13zdby1jjFNAnsokJEuUuG
8H/58YnJ/xtjAZgV8OpauTWFX0MdC+emfVRwlaKUpmUqoh1hD27IHDh+ASp5fj5v
A1EbfoBY+kMvBQiLmJ0xmIkONQkRxLX7KurJgHUW7U2MxeRxHIlFqJeosqQRf4Cs
qhHqbNje53n6W/mi1lKUagj8DUYTTGWxvGVIWIkXtap6bbK2IumdnZmOAdqqOoDp
lLxJ1JTNLk0dSaqw0ZUTQrhAMNeUI1qzy3FMD3EOgjImloZqNUIcKzp7pHaWjhaj
p9vs4NhakUnkXeVoHNLi3UyT22ZAzL3znjxdyb/Xt1H6HiJVzUZKGLXI2oCxkzjA
aQlZ++/k5auYVqLpeIvXpKoowUXerhgd20ZhQm6w9j3Eqzi6IqFv0/v5w5/SmQq8
5ezYq6crru4UmqHJ9X1LBYtQOJL28CldkH0JMGikis6dmVTIAQBem7jU6yuSaDYy
5s+xdVM6To2C8cULJYCXvjUOm4WPB0yBiqZnoq7ZQonUHN7jejGoTYEV/BrnUVyP
/i6HJuK9bdq0y7lJu/U1OQFzNEXSe7H8oA7qEJ3/nsRbVpmRwWMilg1S8j/zVOhg
Aeaox8kNzYZst3Am5rilElBF+cSA9IHUcloUqyranLYrSkhbRxs09aVjLr3CKePG
cwt9RuSkD0CaGmU5/BSOq0+J2tEeNSnnhakneP1Rf+7RCTFLmUWXI+8U0Lp0SDhI
xwGxesSTM518461Q3k8g75evBVEDJ/RFlyAR0075DYDeeYJDXDTk2qtjLp+NUhuS
i9kENcMMccYoN3LLWwsWA7ZJQwL79Yq9cKxYvPc3whx+DCTTBbnaS8cHNqKGUD0S
hE9sSZEJjJiFQmyMDvNHM5Bchf1DWKVhdw5dD345BEe5THWkwzo85uYOsQGR/Ap5
2D+sAFGYYj9XKgAANKkXqHikIfAi8TRBQnCL8jDRxKz/u2dmB8FkVkqgoaxZebQj
1Hzi8Sk4tJhj2TdfYqD63WX3zyChptkXbrwqcz/rGt8w9UBTT8O831WYxQe+AIPd
anCDtaQg0pPt38LBIojBWLDWhfPe0PAiYyUj0VwmIuP7Q5vJ5D8REGPD/M9ONOM9
k0iZGvdOYMsLfjEu7PFkspPy/wl5lwYSCHRrD9AxUNlWNm0CzdAV09d2IdZXtcOZ
zpe4mOGOoQIfuB7OHxSB/WAOmPG5uGVtAKsXNfVIo9T2krNivqZI6z/O0sSpS34S
ykoK3Rno6vdY3YXCVue5Hr4Q0hpLgDiBk4Qpin+CxGuRr3gO7fXjua9/AGpwB00v
OU3loXM1lVBsiPpyggKWLP6Xzok9zlzn2dS4kRSnTWKl5mUR3KskD/fM1eXkF9Rc
P78FNLjBcocXqyCFGWjNEd9jSIJjUjtzKDYt85WkRcbtZLVnb1neNYSy1IGf0RJ+
PvrRMoDZWOa/uMq/cLp53rw4jSKrUjaUMiBmKEUjr2BPTMdwus17WG8WtUotrwbO
NvDrafFWLi0atQdmBhn+827r8Wl6FIZWZR/Bl7r/GtExZuYkYqVxWARWRex7/gdp
mWFECqX0aTiTsGbR/UeiQDchqObKeqygMCxhP6bT2+PR8qbSH+G+0GnwPYM3l6Wz
j7N3GnDzP0l86hHJF+1XfN9AtC8XlqM5+PdlYHsMj7QHRynbt/uzmTIh6itVq/+t
WfqJqKVPh4DqNcN9MDyTUPtmyU48+4rdrw3MM63xkw/g/X0CnO0mMruPCdQYIPBJ
SjNOlPDsTiVPZKZPfdm323b89mdY3tjvg/+/5hiYr1dX4VBotjEEvO0uJzBYQ+Px
6tw4DRwv5hCngXg21NthY4J4OxPGkkzkuBYu1Rvf1trT1OLlqNl07Xqx7v4SUg6V
5p/FSWalIBE6VGfysS/yEiSV4VO16PSk1/eihJTvzsqRvXf7YzIToLejpmciBmy9
kkkQ6Leye2t3jQ4G/s40FUJ1KU3gF0mOEKD63o44xPYmpbALJBLHvoNijI0ph1FQ
6SYG6/1OYhqhix8Z+cQk5GlHXspgTHp4/Tw/9csXI0yKgSHQWZD0EaitgfbjCT+j
ILdWxYx46ze9eRDdZHblwuI30VpthayQjs1fIU7NaWQDGn6FMK2q/r8/AT2tSpvP
OPNt5NgnHxIredjPW5cbSghiyEUWOlyddUY+fIWbw5gBN2SSqTtJi4VfvB4YxtsU
RXPgs8J/5bfaLbfPfWUL//6ctEEukRYDoFC4iVI8CyTDItV5j9BgZ8ELB+xBbj2K
tLk5V27MgjvmecwVr+DfhKo+QlCTSvR1E0ci0C5/QiLNXDVTUmyu+p0fGLmbapGN
bT+VQPEhUXtYsUjLhKyL216dQgX9LBSNyv3UJbQ3i0sGnMcAGq8j9DTuWJ+kb/C/
eLtp8OgCJhvUwdtqfZrY0Psm6GU4/un7S95LueJxLqLglnyvFzXhRhji9zSzUnw0
DUZ9ERfp5IzpyuppnwV0O8K/RTKNA7NNcOwQlX00jH7kQx/7AkSYSEVTdRClmRMq
UNcnll0KwmKDZ2mgmqxH/ITYlWVh55TI6LtY1gO095CADDHK1mtdMbqTh8xVdk2M
RWsIU/UUNvnyS9pQzxBZIWS+zgNPkHCQ11rHGiZ8slvQE2bDxzP5Mr2ywUDCGBIy
Wk3yjd/5LHDcYs0HF0H+b+ZFZ/NCRrNs3H9FzdUbJo3hPXtO2hB/FfuOWIlWJaAB
bnwDIqTY7SfO/TNl7SyjdGz2mr9193X2giSAhdEMmD7NgrQuvqy+37BluS7r/plb
UfxdrMMm6eBq4zPt6vxOIup5aS9GoCHvCAVEjH8sxFA1ra8EDy3wIPjbcXWox5nh
gaZfL3iSnmAyBQeilPX+SYWJk+Xe8pFt6tQVEa4wvFB8X3+2em2TP/vf6QFetl38
uZBrQEwyech5sJUR/kwjt9A6B+/azpunVuToLGgjQjW794kA/SZViFQe7qvAw4g2
18WQohgZbkz84H2xJUSGRPDdoF42OaJgOr67n57uH9Ud/0CCtdxMbT3ynZcpGz4P
rQmuqRwXjSZdxGt2g4SCpgqfyzqJ+vtxRUSMvPptUZ3TH8GMWaDFGyq1Ug5ARr4o
nOOoUR1fawKpWLYn664huiQYQ1StUjGxoCHYDmZQbcvD4kMF3Sj5fR8b5yGj5qPE
tPitGCYJ9bOj9hjETe70MlRiFInS7SE60/MRwoKr+6ugqOciN1G6dPLlnpud1lxt
PNn+rzGG0KsiOlgv+mThu33cPhECrQ5SdGitYQd17ErlR8lwjAhz5q2jv5HCKHEm
cFxN9ZfmDR6m1jkTKmqIptkZ24yzfHaDBvpAZOCO+bD/dt1oQyzeexOtyUfVlRHm
63JX/pLEaA4YohCi91m/RZhWiJvLqTYHcBtf//3xmS9DQKtc8TkcOig+FsoxBboP
+u10BzF3ZyNzoDoXazhx8a7nQEbR47lKIwgfgxX/nR9Xu/VrIP8UOXWMBIoN5Dzb
MwPKCA9Vj2Ha2mNd9XL5+UTWOXbzPwVyeu0Bq9WJHbIQ4jADOLuSuzhGGmHYefWZ
mv5WPj2dwdIfXG2HXqEdKfhNZ91GOQOARMFXbybmvarptfFCUuwV+nMQQYraNYhL
RSsjJMEczNmEq75AlXLZpz+9eVKFVFuZ1gHfoU99Qt4LuIAgmIxZgEvIFvhcrqkd
SYpvQdGFOEORdbYe3XUSEEyA+xaBzbWN4jIxDVVEuNIM67mKrzIKwLEy0Erut9wh
6Hbm0d3JTFANOHN69NhgIKGmVlQSp+wKmtlbifrhsy+U3HubiMZUhMfIEzaiVv1W
r4JuWzZvK5sTGTNfNm5nambFdKZ/2gYR5HntZXhRvdum46q5wq7+pl55Khf91mJt
NoeM1Jc81ruGo9TtPYjYAdfvr7KeOHU7ROU3q+o7VuU77Lc5ei2ggB24GJptSrtW
93PvUul3ekGomcP1HS+h0CeBougyIV3gTIrS4JdWRMX9wiEVpQsE9zvfYuRFUZf/
ihPxJb171sey+FxPe7kOOjH1vwBtTaYlKeJZYfRqdIa7qtGYO2jM6ZsSCQElEnxY
BMKZfykjjuZgFKDAQqjkBEO9GD2iHtG4x0xAHaitOfjhL+ugagEfztyszYR6Wa71
ByU2TGXvHMiUo4+veZinlLFoegwD0qPNGlxPhm7neKD8G1pJnFUjG79uv2LfeqEv
k79IRG3L0PQB0DENuUaxwjHYW3UPGcQ4qvwQncpbumjZG9FDiMzGgxmQGipEeclk
0L8ySHAhqHazh+q1FWQ/6L1V/hiv4iUO4DuM34q0KQjzQh9ysk+v23WFAkgD9wcZ
N3Ifa3aV72nss5dCgzGNSlLo5HjPAQ4a6iaLz3WQmh4mKXO68wz3LYeGEQGw4jE2
Wcj4mVLCl+eDd4aB9uOn3MW9x5x8Xu7iuY/gDyfbkBVZ1hvjGeLRumG7tsMuUiD5
pca/xMlNbdR2WcdP6S+IT8x7EfskjUN4vw6WP3uXShz2drbCVHxzmbsmlcE71hkP
dbjFAp1bYu0D3HzHpVeP9rD0hyWlIFZRXz3xdSUgcfWWBrin0EQun2A4xdXS9x7U
0o2DBtDvDHX7xPxWsekWKkhCrsUebWwfNmODwNE6StzfnHegxGoSZ2UmYMem1EwT
P/U1w59P4N+N3ZGnaRsxCntJb7grE7FLRKurgGlS5r/yejet91Na65UyL8RcdekC
qr9Emp07/yvydzVGEsA4J+T+KFfx6ecpnu+u0wV9lVAF2uJMkKQhVhD54UZIi2iE
BqbHmecEGYvMJehLm7o3DB1uK/In8hIym/EYvVnhQAFCAOHlP8PR3MMXBgTmkxhb
sed4bF+/ni6ixOv9ud6MU4xR74F2w5XozBpa8yUvpacclj6eREIVXu7jbqkC4rxV
De1sgvaw77Wl8wV8Pzatspdy25odLSa3Gwu/pC5mkfD3kt6wUFwE29I3PMZY4C+d
X6v0oNVOunNxVu6dPrl5Tw==
//pragma protect end_data_block
//pragma protect digest_block
AYZlBTcUsipcIlCSLkqYxBbgoBE=
//pragma protect end_digest_block
//pragma protect end_protected
function void svt_ahb_system_configuration::pre_randomize ();
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
B8/sepYcpaIhyi3AHB34M9rsKP7wgrumc3Aq3un/37txc7LNa43fUXCjlWueXPnj
JbOJpu6u1f2mUkthuWRL5mgCeUfgirYgKrR8zu7QDRSLzzqhYTFKVyfyPNT2r2lk
aAHMPi3WZCMiCF6FVev/jQ5CQx75gCkLSPAwC7sUFkbmCtG5pBkEgA==
//pragma protect end_key_block
//pragma protect digest_block
Irgx4IOFxb/bk5IKNLA37+g3bD0=
//pragma protect end_digest_block
//pragma protect data_block
tQfwyYw8rwOD/DlCoRH9CK32zNFJE5NISufDXmP+fMJbTSSmI0R8joxGZyr4WLQA
3Hxu2w8fKNacqeK4gHTM3gqi/D1q01F8gL1LbhKDrSWOyfIc0rBKToXSfw0hDPTX
fY+BO62DCYqvtQtAJqjCSpB5UC+H559QWB0863NPhb7FQv3gzBYPp7uakJ7TQlou
Xay4NoBmFY2aJc4iFjpRvtTC8Tezhei9GyVVVfkClZ0vJ7m+wP4gTAlkjUaXo3r4
BUEoKH/zRIA1wABWanMSmoUMsn+mnet8SEhp8GxcdfcaOqqV664tE68e0+jQEKly
4u/LOYsj+U97d7hKawkphLxpQfrHxnI+Tt3UjVqH+d+cn1FOPLU+JeDSX3M8EvEc
9FTCbGHrif5seP1Hc3m7RxOqEIIRHWZXuWytNHTJCf2aQi2veAF2kfw/5ReQEnVf
UmrFQO/4zuP+GrgUuncX5RU9+g8CrgJeb7jnG8ybn9dDXN0epuWr5y2rnioBGM9t
47mySiyJSmm2eZvCvIRMXicB4E3eY777y50FNvILLry3J8U6Jt053YHYFFvu3++t
dv28j/jkD5DuB+fpoloh/jtCZdqvPRNMkD4qIc8oobnPAm22EPBQw8tDdwZGwax7
S3rD4LEzN2mCFYaO/zWk3BOshvDPdXonDlWNDXA2MQQ=
//pragma protect end_data_block
//pragma protect digest_block
9cvfInUneD+H7upUsclE4QFC0eI=
//pragma protect end_digest_block
//pragma protect end_protected
endfunction: pre_randomize
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3qrW7PZIFkyIxamj/nSZriEgobmuXVIK1c9n7NzOU5oqW7d7B6iX9hUmT788X7yN
4NCmYR9LX4F62Y4PMD2H3vkANsSQtDrtcqjMdfnrpfe1k/7f0UJDoEO2Kok1w2Mk
THpzyd5//gwu6JdlcVOnfO1mWgb400WKaAJVqCMZl9mt+jAQcoP7OQ==
//pragma protect end_key_block
//pragma protect digest_block
Q316v14YGVZEWaZMCSWB+hR64SM=
//pragma protect end_digest_block
//pragma protect data_block
bilklzFxzDtPjhVNu8yXLQZpUUArG/7FyQKTakXzMQzExQztjOhViRAAZGo8RKov
6KmVOHVjpWkMdQL44Qdfl+PyoIE7Ln+ADs+XMiZuAST013JV3GtD72hkw1BuOt1/
DkGU251tjFLJN8uOiNBF/8OvTnTcvTZnlmeU01iyC7kgvqlZ+n6Pgb+gifH0ueWn
Bb0wxmbVj5WnvHQ4OVwgyMXoipsio1435Rupw7TnEfrL9qgj6iQQRTeCaURGy+ap
ijYqXYFH3seBG/VSwNeqOmKNuMx+GppLgcb91doEbo5Lilds7oAF9phHfymsgEKg
oL+Yw9vU+rN5G1YVcASJ+TtPdhZVEZIXK4Hku8DV8U3aoLQcHLIZcLkwZUNdCZ9q
l1JWaKSmmKZf6/5Y3S5+gNaseCNCJvWRBzhIrHtIOHkX9oHOhHnUQJbY9pAGhjKu
3HsYt0TNvQLHXR18P0irjZ3XRh1TCCqEicXRM8xRkKuAy26kx7wCicIaRRIYBKxU
Iumw5l582BCRP9BOiIeH9xOfGuVKl+Q0goVNEwBe4nU6jLvjzw9z/lycVFGJmfVV
EfVXXHgbsmeUPNBdTZqbJ57Jw+/SNi8aByZTq7gEO7Z6YQjCciqcT9AIPNjLGFd0
e0uLOXQensUxJQZAehAUSEYgzas8UoKfwqDRm3gCMpY15u+hLM7/2+0esixBd7JW
wTatMdqabmf/7Ty0X2ZsOs9lAfE09mscs/PeOxl5PWlOGvRanJ6gE2m/3qfvQdNz
A6asAzOkCTQU0onmeJcoC6Uyc1J5bQfecQftx+j4VrWPky4bmc3DTIJQXVMGhYuB
DH8kuzYvEjX9LokuVPAjk9/vOcaHUd9ZtWKEabjoctNwiRD7M0oAKPSSsc4KgxEC
D8a5811CvDMMsM0TsdSsjEoHJj/FbtE1aZEwtdixC+KlkFqwRS29FDWo9RtvQKBu
UYwDLMKYXeuIyJTeg/zQCJBFUDgLMennw3jYYoqc7xwWJnxfmO9/BheuzmCkMVgJ
12OugZafFMQ3xkjfrwkklfoeMyfLDmtGhS1XUdwII9fbidw4roOSRUJ9IhY4ZCmr
KsvxcTDiLQ102nZXmTF5oTqTCO1MiBhlvfGABEGpnvLcw8oIsHUJHyr2sh7apytT
IGtV+mzZSfkEfZRhxAJJgo/ZnQV0UCISLkfmScowJuYxlT0pBbDBJjutxytD/0Jb
yXtnm1lNqNefbu0VkIMQTjNT94gk/1zbYQSAkz6Mv4i6papigX6bnC3MLwyU7gsI
aIPwcNKGB/aKD8zOimeQXB5HDHrUnwR1PVEzi2aaHBYG96Dios2wwigIWud30NcD
j48y2G76ha2fXqnyYTECke47s2G6kiyJVuBMykAtFLs5ASy4YYepUkA4rdkkdEbL
mlq7KmfsR9qSUQapVlga1Ek0fvGrg4CNzXxEoo05Q3haeZYRGNs+3+KEDLmfExzl
r5WxvXGqAUYpzRslKLW0a1aNdKK7jVAAc/uFASsO7yFAiiB8za/kTeQwe2f6/7sp
sLzfZInaSxTyrEl+TtlVsJPWv37JoUW0dY9Oc14aevRYxWy1ehbwNt/lHwfb/I0C
z5np8Ho/vucih5N+fydK9bBEvPIfXbkIYb2j7uDZUutiiWW7ajYQzEb8lLdaUspa
OEe7Kg5MajR2xFRsMc3YIoeZh4Pz4xTYz/9Tp8VxNaY0x86XP93S4Q6dQjoQpUne
fjGq/1sWDZ86rY34YdQ5cdgcjpkW+freyDOqAg6aQn1oNHeI2S/tErjMppbacjhh
luAeK8+BqDxRZ5+Jt3xi4x+zidRl6vXm8yQGMDCJN1X5ua4YlbJqebSmUozQUVkT
6IOlAz6pffU4hBfg37LknEp3DTUzgsHwh/sLAylNl43U+PYZ9Ner5yodP7PLQ9ea
F2J77xrUYu1nHQ0WdvHr49/XKn9hPPI57Mepw7ObLyTTGVg9XcvgQBH6dLs+c0JJ
5CbkQ6I6FCiB+cwS3V6tLD9S4x+EvNoGA9dzF3x60e/mN4/BeyAACxKaSsfTOrmQ
pkb4BLJmr2lEm6pk5nKwjnm7kckzG94TebnYnr96UtJvLBoxhDS1X+laQZCDfy54
WWzH/yZFbzdaosX4Fm43lpq5/AXqo0d0PRC9RSggVbsL7g+ZmvB/H5a43AO2+qBR
Vrpw3h+xAM1uwCR5g2CqgBYa/+zDp4s78p8GbTNHPKi2RjHu0lLsh4XCse6M2jZx
Zqg1Ju3w/Th6YHDcjlSF0NJ3M0RqKRHAukk/2z1hbqP+YFrisKUF3CJX+rUW+Z7+
CjycYPtlt0P5VgI3wwijr4rDNo5K3hjF6XbSEgqFV2sVuWxe6QOvCa3Htt02C9iH
AVyy5c87czhlq5cofhA7O8YQCBUIDttP3xncH8JMGiWDBBVmhqP6K79/N+5hjSoq
7Op+suqFiNJEhdSfI8rrOvNm1L2blDFkTz2lI1t6CO010OMYffuUy3ngrmBIOjMw
Jxjh0l9ledIYI5f9yxEGDVg2Z9bfeAn53p+O6v4soItTnQeH0UNibQJXCpfKr8Al
jC0PFeKGh31BsCOSbP+UD8ECpjBWni82K1cMoYAJwOAGauJvzQSg5YBV//Tn28XH
wWLxDjb/nxpSLikwubC077W2zwx4qthepVF/TfVYB7CWpvHTojoCd9V74JFzpAcL
+oolBdeymnHpgxSFlZE1tsaLTeQhZM6oRad4kWEIaOepu6cERuGmfVKUkJzxO/Pz
h99qMyV/9LNpsDjSCN9gkaW6ns6iczUuWL8AY23YGTCSMcrFpOKtY5XvQ0oMzrvH
CK7zLbzog7kGZWzoex5a8CpVdzEw+E5ZMChWHrAm31ypznsq0qERGGjuXN1krgXJ
FuNADL7PQXqLfeHQAknyfJkI62gzlyYr/DCjSoQ0U5jiB9B6KPBt2K+LZLsS67co
MQi6U1gcgCSrMik5u1xe8Kt3+Ou3cbSARiIaPaYxnrD2phWC4WG7i38BQ+7BI8HF
KLV8BIbWbik5A+AWvLfZaTxU3vXPSElg3D3rJBGuTIDuLHFtEfSSQKZ4na+7t5NZ
Vdy8AbP3H5InPrBJuFduIn3Lb1ywAFtcIXc+VeiW5oYP6d9+fc/qZ5xoRxNjJisU
ZoZiXdkhxYO30V7MSRUOS8AGkK0TpZvRWoKyWdm47XBtNi4rL4i82v4Xoo7NyWMw
o8tID1YinU5zRbLkk2XDGbWLCqd0bNv9y7oX7RG1ADXFwCJoYcSe16Q6YQo15DQr
QwfkWyV60NQ9Z41AEepJVsnkbSV7bIYEZbgdgK2vOr0A1fUMRgnbFLmUrU6hR+84
ipwTKVG8OS1siWqB0v89rrGExgM8w7vN1hktLK9h4hsdJmtMXbl77Nh9aYwlrwj2
OR2x/fKfAe9zFBM44KucXENRXfCCYzzmw4musBl+pmsdPbstxEtGEP56DnidCD+K
3JvKKbvgspkMmkkAXlKIBzaleqcyX1F4dik/y3ALqDnlo3uh0G5LnflAuYxSvRWO
bD/tr9hCk2nivbneEGkNGbz0kNz+IOQnzfyicQNjxotGirmRqgl/yHcUMinLKTKf
ReMNFA7ESKC20RppnUCLntb2syIcKxGhuS3OtWBae1SVRa8xwa+xZhJP4SmBbPyi
JRxVssdHMdTLU8Mjcnhyl9JY2DJPcjWTVO+odfKMF/PoXiBwEEDuZNAX8VnEv3f6
Ug+U+WpKfn/JhdN153rfbQz48evIbuf8kdXo4ubkkxuqzeshf+7dARO0q9BRu3Xo
PHkB47uV+cFBBiGdhl2PhvxC7zq5DEjYb2+Wa9TqZfOMJ2yxLbdoKFHlhZQSgkem
DCt283DYd5RmfkvakeIr/JJjB/TDmB3lgzLa+bIgCIW+0meDCsFllm0yp25ECQLj
mvPD+QXgbeqcevzBDcFJfBNr5srSA3Nc6f0gKdlxw2cba2EJtdpf3llShEjByWhE
3NnMGEGcBlngulbDl/mdpp4PmXqPDSYQiDDnpfD2UCXKF1IXNV76A5gLL5jmQW/L
LN/sCJFMB5ft3O6UbCPMJcP9Xq9AhHVIc7DNZT+Bw7/SlTPri/9lZYwlKAv+/I7Z
8W3vutFa2ZEqWO5PESxE0A6bsSQcGxmRhRzn/UeNn/4q6pNpyxtTxoSU4aYOcJFC
IZR2VpoO3bzIuSefKV1f9d4TEeL2Xt6UNYyELswV0fOvgr8/mE9titrDhC2Rs2OE
zLkWeIcNMXvcbQ4BJb+YRjuhvd9zKxndjwAsr6/KyLC5IaErrNjphn+FtIMdcfY/
U9HxIDTrFzSE796jRQW1L22GbLNK6R6U28c9yfAt7c7HFDYFc3Uh7qm6GCtbf6Of
Z0EZF0KWusvM4w4A3DHiXY95rwOzg4lUtH7HvBPNv8/pzn6jXuE4TpfLDiPT4PhI
mt/u+tPEkis3PAWUsAMyrLdwTooHkEGHunjvhoJ6NX/x4ITFp16UpZj8T0x5hAkk
KgSAJyQyPC8GOx/m1AXUMu0brqJe8N5+zPOCkV81MxsTnFjXfX7DP3L/U+I/yVBr
PDcbXGRYed7yi43tamCgLen46mGJSJPWS/0KEVFB7Em2HJrZJPf79mSC6Y1kjj9F
nfGXIr7Pywsszm3pm/6YsjmlLrWz1L1HA0C3t2HOHpt6FARC15L0YNFPIPl0PNrc
zAUvcUz8t5hAS2W2NdIbYqWu4j753hQf2xtb1d8yr5aNcfmwOcIok0p/Yh2yDbQ1
UTrFHNtOuwvLObMM21ow98G6MZYDizP3tcoYiXeiYG3sCegEmBO9iQ4Omkzu/fuz
Pec8lyvU6yAyqRv0JeJ1KTXZk5boX9V4nnFG2Ijx2GWlwqjuw8EgCChC6yT2O3by
98AxmFC0K4wzElfEi/0MpRW7ZCF20qnZO+Q3WDmo8t+TJUbzo2Nnh7A2I9IFKh4F
OVDQ6kTXNRInQ+qjPA5u8kJOrYqG4NUxn/phy47WX3UFx3qEYKFqy/PZFM4TGtLj
FdGrpUw8Gcz/OtZzECRv+lHe2y0vfeEd45dZCwwya2L1v5TqUfW3zXAFUE0M2/Pn
N7SS4pd+7o7qTowqn5iHDmIZu7BMz/yMyp0fbxsKbAi9nbaLN+5p2A//Swtokx7K
NNRcnB+QiDfIJX2dG7lBoYHw/jgSuGRb3B45PaYmexG+Ia3z78gnhN3RETwai4tE
SogfixW8mYjN8PA7WfaPpVtzpxlkHCruY7c5ZikQQuBYuXMqWPo823JRhK8MxAUR
e/4rueiCtJnr1g6BUy6VkYFmPWgS+9Od9sQN+qviwcPCsQFx5m/yOrLFsd87cmIH
IbdDG7iTyOoAMDCMisr05mkMmR6wRSyXWvx8HsSOrxBiW8yaG5fWyPg0xhmqoSJZ
hSnHUFPN/Y84rmUfZv5qb9lnFjOsdqh9wFEYB8QrQWvyGgF5waI6X6K1cXy8of7P
EI9QU7o/5tsy2us6/pIaD1uApNMVJFM/8CAk9wteRflutCwFqZrMRsyOQsAdoAxK
a4mvQwz/vA5h/gi3LWaOyENeM2GMDKIat8h40MoyLG9ZtpF36/7bosBeTLaVCvX/
8YV0ITeZtYbiOwen6ZCbJznhfiZn/QldcFaGPj/JJJZF/oc6Pn9pkpjGDIyROwML
yhuBzfdOi9XHIpbAcsHXoVB8uShdiXQZBxci/f0Nm8HfPglYUVNODgvWfJMVB2SN
00mq0B1mLq0u2bNaA9H/h5suwVg66BtfmPMeKaWZiZAksL7XAY8rrIlOdHofOg+Y
+K8Uu8bkwvinTVh065FMvQxFz5htduol1zHn1nDwBBLMJ6mzA2UPUGwDpYTPAq46
DkH+H1XcyoRa9jL/cnUrQrW6JyI6gxwigqhBRgq62oiArErDpUnJXpLoGtsVrUK7
5r9GAL+vuG8+BTjkwDUnsK5WY3wRsxavrfwS+/8W9qbNu93xkL3r0lWhU/KbFRHF
WnqlXQ+3XqE9+oBqxnzu91l9Ol28wZtXsQqn2lySDJZvGJhkhzyv/kY3d/QzdH2G
Ycjko3ilmL+O0Dg6/mwWZBSzSwKBD8fKUdW7+uByU0+g5Zsy+cMNk6gOaYfruCsq
ycGU7SrKcpIszswhFltOprkHM2nUjepQX1IXfZk8A3oX4uWYQPqojXuWJR5YWtCO
MHXJeVWhxmVz8A9YE4SI3GocH7xIxy8YsWlzZK7pFY+aD89SuBRVwzEJ8u3mKvYY
JiHu8sAqEayiamBlOynUG332IB8n5U5MQoKvtX1v/P7ZR0DaBdRt2LqwNaNTWUni
Snf9sbx7HlkOGP1eSe33HrTDbYHF/BEoKNjxGRcZFdmYk0SmZSrnQanGvhSiktis
XUIZ4Sx+XGY9RHDF8ME68rzdEEm6DT2FTyRLGdmfJjwcyWC5O4ipGw5J0ltrVv2U
YDmB+kGlNrDa/WiByuKHFBDUyrq3P83JsEPcwo+K1fYviw0NJSN8P933jS/KuYJL
ZOEo0tq/dGW9yEdcrfYxHP+Lx3riaBd/ATP8EOD3vqkE4dysR962MHwODvi+n97G
geLP2f33u/SvsuD31gXPCPsg8Hf7yaHfy3pxlwcU9lXWRg1zYTJZxl2g9uPtzYyN
NS4jQiollXyEU5Y9xUy9XQSgpeKMWNjN+GV8C9DDuSXGsJsoV0vob1vsB5xw7cA/
L26FQPPua+e325BxcjNSFd9gwWLHAxEYQcdW2fx0GEDWqf47pFC7xv0sgahB2P6j
q0yFqNbSWMlAuFu6gcpd+XGmGgdLppT3oxCDHJt1vLFmwffmq5jhsAZJOSvEsQhk
Dk02E7ALEYc3YzmOjxhu+ahkh1rvhzKKF6Fe76LzFOyuy9yKUzmVWn0ACQIifiMR
Kt/t7J6M4cbXImsM34KqO1pfAcXx4YZAYNRdUUQMTqHiCmCQxXXvG8GiQWWZNsjZ
o8dIBuB2W3AHj/WBt5V99htmKoxPAQdS8mJbde4Gj1sHJUaomMcMAOdKeRL5i3+3
U9YDJI1lNgHFKgko6hQMM2H0Gf5VCo3WtZVhUZPFLZ9vHezCBIuGHciQTZAE3A+e
rq8/zqRdbw28YU3M86YQVSJyyRFDJDt1bnLzWFHDK/EbwLXMp//GHNOO9V63xTDi
T+5XDplsedqbhnMbmWsSPb6r0ZznaRECvZBayqhmLt6dDt+/IMo7yUzMgxc3XkuA
51Ydhv1DX40NksW4AIZgL8IXZfyPZHySLJS0EKMHlMhVLSxkyODqHFzK2zfHbMDJ
3Pko0sgGttZP78RlPUv7PBqXjbYlQSgg986nWYB3/EBbvTb4NNZvTUk4+ofcl/CW
lzPlLN/xguX5OT4LCKbKmEtMeJr/Q5P+zNA+v/90JdLWhP1Fe39394wsAOabuqjL
7Q2i+Er+RTVPrxFA5d5pvtyCh60NZQQCf5yOFJdUu1hntj8flRP03w8GlZbP5jC+
nMNi42ZuIwKaIKJP0IHa3PzA0CkhNBevWt3WxRqxGUfUw15SAJNEvCPccQTu5AeH
TZXfTNICtB2YN1DP258LzC1IrILzWVGOHdidXei8bNRjyh440iOZ+IP7QkZYaHF2
Pw8Q7OqRxNd92S7s+bhGh73vKFcwqpITFJCC9hyDC3Ia5CSWVAxhpqvV3OMzfo02
tnkr1ya4SR9wYdKJSp/kpz9bOjC8bdDyZLXb1NAtVr4HCkKK73q3anxpoG4KwhsR
wLBIUk1x5SR8aRzbOlpvlW/YAKUCX0dM4omF3/d+50lYXHttKNu1WtGpw4nJsqhd
dW0Wsl8EcNNpG5UpT55X+WaDKsiPnSwfzjUmPkAy4wUu5A3t/8Rimp/e+DwF1sQY
Sl0KkwHn+YDbJ6R62d/5WKw8zN3Xrhr+Nu+ckeAqvfyJWqr2eo19qlpDeY0dlPpm
WrhkZ5infi9vcChCZu+Kv3ETglL4RUzWgcWK71VKNNce1cAdDpwm6i8y26dQo3BM
fjD4ME6cgUD+nrMsNru1DefO6pYCbOHFDka+gr+S8OzHKy9lL2Wqm6l6RAubZN+H
mmqLkmq6sC6FJWfqMtr1PaZYMnfPHZLbGbERV5WMOf9Yz+joRiH2Xz9awioC/d3p
Qdxwfnh9aNK1Qv+G6VCMgXoIDkGO3cgz0LANhvxTxtaupIBFjy96lQFxtNHtINyH
5UHkR+etA+22lumPV/3ebHO6i8Q7ejVPMTyOsyIuJ2NjBobeLEOJIu/CUV6zTTBs
OKqKPK8voTbbvTH1sPFDpOBCCa2dmDelaQmqciRAfbbbSXfrcgxbkR1Jp56MhsAs
Z4WE3EVTXSVR/qClt5D+zg2I9rUPdjlcSxaWCKqxYk/OHxpnx/nY/W405jkRLDwH
Pp7Plgurt7nV4PM89lQaV+Y0bodMDA5xywRX7Ro/26uoueHRVEd/SSf7NTe5voxw
5hFir9inUrNntzlQ5vhF+ipf4YLFK+FstnTI4RctSr+k7SUMkuTzEW2MXLoec24z
RFW9XCe913MG0Q4dG59jaNiXIVfPVgMbfx6CBv4RcfGy0UBBl3VkFNXNhs+wgFyH
79lDP8lCHuDM1hiVa/vVDoWa64dpNp8g5AqaJqpFpH4K0Isnhnu5ORCCh2AyedNU
I1/A/FYeLTN36Y8LHy/IfOlmQ/6L1fVvbfc5E/bypDjNBZmRiXBSYWBXokM5lIvo
J0XgqM+PTrTtXIg8OxAsL7fLF7IsuJxuw1TWPTiDfnNua8i2tQs72domAdt6XJ3/
3KRePTDSYQ0Ikrd84HUJfvSfU44xpqYxO/SiQoMMVItC0HQ2AilaiWu1mSYaPZkK
C4xruNXE6xouA2pME6gbPceZPQ3MkOqCBTPpjHdSZAy7NSEU73yCcrHDWGkFAfcy
3A1S6PYeGpbOtyH4B9xxWOgOOU+wi30y56kVJMCydGecw39TkVnnKvqjGSzv9iKY
P2hpBUfIcr95jV2BumYl/t3ZvvHEf5MN12sc94Gh4rCy7KVR7AQ/dtuz+gIREIS9
4XmClowXWfuERJXwtd2oDQ0kpuGxTRWBwbiIFnZf+tnWGFqmBCY4TFsE43Pccv6N
CHE2xODKo/80g2e+sVQGPYPOS24q0z7lxkI6cCUBWszXwupMPMeqlZjacgug2HjR
h4pu0jWnMmTAP/GKmUQSpXPBZxcumuyqKzACTzPoUojKuiBuSRFUnji/qJriKqyO
yEW3uOkaecA+62MUdw5jCMuMSfAEd1VvH1eYWyP1cb7fNn2r8dTz3eqOuMO14yX+
yUPbME3uX8/uTL1mZgIyO+3OgXdANjN7AvWaTZxJVO3lIDujHIwR9u01NoxLPKy8
7WrfkfNkkKwQCSjvjC1s2zZrLATj3KKLyyza0fJvpKvJ6MY8699Ky0Ur/fD381U/
BAS7s0iYsQVbPEwgODXjiPtZas4lQOelrIW5arVz2mdL0Ne2XkVHywYkud7qhfh1
LuGgcL8mwLelzBnNTylb8PU1j848YQPB1X2B3EVdVScamznnR5HFKRDW2Wv6NyqY
A3UnEvf7v66d+G/aF++76EaFpINq1OuyT5bWBFivhEgPHZk2+C0nGUvESw8Ke5fk
yhEADKqxTOd36EqnXsBAm2mUiIO2qXL+hbtu6w+3qBxw0LUZsoyuR+RoiwDr7xBw
fKWf3NVleTyUO59Cqh6G3PQJw88VL5zZB7JwOQbUmEcj+oBEdi3LoUdIOFyUbHSG
ohgoJpCj/jUBRqxHbKaAYG31u3BzvwIbvy1bCNp1ej1OJNyfQlyk6O43Vp4Hfo84
1IqSI+lMqWJd+lNB/jZNUDu6jTb4Z4jyd0ocLjy6rDRoMwtwQSIZbGXL4I6KCeY5
xRGJ333RSJt700x0oTq7x1saDUjbShDz94nWOWXev9ixQ/PFGW96wllCSyY/mOax
eLso3Bs2s+LEJDtU6o/3R7S2DHOKF1ekE4kr4Z/QZ5q8oUZjDktlSFXI1iYce0gL
hgXDqCYpKseqc0jPRnrOCqbiAbM7NAlQoYp6QTVOJanAZPJJw/qpnCV4DHgkXa3/
5dgsuqAZ+dRwDsZrMGphXr2Fq6DXD+RnH87pdRLFNUE843pCeuhbPXKLgomPyHZk
c/cZ/tvCtL0Ulb0CZWk/LMsNanQZf1ZwqfA89398vFTqB5/YLetI7/cHPRBLksmX
48HjuC+jxIHMWci6r0BuQrTsHZIWZb9N3QJ2jOwKPkKWM3607FEg7JqtoR94NyZ4
qE6+SZyAV4YdLSxb1Iqr5DkslNNUz4OszlxkA7pR+LPeIyj9+OJb51bfTtypGKfy
ZHXqJl+D9DSCePyoE2LdIMLvAMG2gSorXtYCjWpW9U6dChvnyCaBVJqUMvRPSRtt
NIYsMzqiTX1cyOl9UExDpNAxAfVS+Wl1lJT87Q4xm7g5H9Iqa2rmhD4o35OJHwRW
q/hDCCDqemr3TBXgnzoU7HDAqluMzALsHnzyUQlIqGfbYiELC5D1DhppLOFb/5mC
N3WnMxtJAwg9Hmm4aTEUknyzWKQxuGz5/uFVC3OJwV9BdoW2rLRLxNN4Q9VVPDO9
BlEps7AwJYI8aHZMvTHOFyaSy6rYfuG3kgOsYhZdBmy3dl7zygTYTm6xq7AeB15m
uCeQGnjLveVoawIGXay/LiyZOPjCHdGNp6HfAkSaSXE4hGG5VtN38DQmDsk9GRG/
yCUoA5k9WnlLw4lNqY1W4Iel0srbjnDWuHNm170iFoaGduCKYdyVqDwTAg/25BvE
l76FaRNQnJwFnyc41YDVY3l9Y/k/XjOb/MI6UX8/ZUdpjYEGdT6hJHRBNsxl4/jk
Ocm6d1+kpXTawov/ig/Kwx1qzr+Wj4VrjpJurBxGWC2ij5jI7vsvTCNn24JaxBTT
i26yUBE1A7OQ7nnH0+BQzs8jlif104zpMk4NQURv2ns9aFCqR1xV62ay29zHVlYh
4ze0DVXrlsx8vr6twnbstDn84A3PUhrDenPuCoxu2zseiGAFBA44bVR+kj6n+9ev
FQzrc9dtohqef3pRybzV1XvjTHEzyeYVnuBU0hwZf8K2GCgj3as5jXhY7IWXTftl
WYgr/LIOvJILLz15mqz1BRXTwvSszCD5JO+fEJlcnoYMysFsHBoV6cM6qxpAvE85
MHuLH6/5UfvVqIgG0Zvre5+ZonI6L78h3cTYQh+/Whl5zKeekEwN7Qf6SdFem8C3
KyyioNYxchQSAlKmbAiSBtPgCMOtV4NziGwqM8rVxXTeFIA7RrjablEJNbuPpSPv
02QxRdcXSy56JLL4ZdBo1BPfgsLZepwEKHc6AwSRHOkBfmc9LnMT3e+M6KIqWlvc
7QdWfW4TKi1t1drN6HCNMo4CuEQG6/NDqr+xLOy6xPSfvGH/fizLCaQfMw/G7cRj
BVIjE+tfSrP4RyaBpzuWDmsggEyFQHM7cgFxqLCQZtNX0Ay3Hq5vfVZAJlUI+1lB
E3dFA6Vdl5fpCp3LJ7Mel5nHba0Qv9kqIVduKI+IOAslkLeCip3uXfaxo5wDGJwA
IE1WBzK+I1clTcdeTsWF+GOFt4REsUgN7O9cxPeHCthcbkhWJShrfeHtZAkkktPS
eNCzCvziNEzVjA/w9nG2vPcEb0+QJ0x0Mp+5+gqagv1R++zPO72xnc1u52fvrKrk
507jUDadsTG2ZEBaTWcW7kawL6XZeofzTFuHDiIX5mHAsJSKfhLn1hvCaZ8UjkMr
Bs1i/0ASTeAVXUHN1qQDyvz8kyqq1DZM6PJQKIX6hlrZC6yt/9u6uMgs3gacpEIo
HgIewzyEwM4EpU3IVAMN0XsLDbvufHlV7XGExPof9ytOB79nQ15LMYVb9rxaN5KN
Ml90Yd+f4FoLuZL/ZLfmPQ02/UPyce8ZcIa+H+ajS64ItuMKnn0a6vndf8/Iiq8Y
IEtlgwrIwSES0dFMUE/YKU7VN4igXxf5rQTGfI8YWShhou2Wf52tQqv9PzWt1t73
fDjjjUjvFzYSvf6hbubjsK6KCOHvZU/zIu8elDQ3mPLXrbTudHDc9f2SN4Z2A4Ia
ChwiYgzYUPnupdgsNy8c9DYxwm5U0rAWJ6LyuS9469XYZXo1Q9QVRptoiFRwdb3b
vF5L4edVoJqyxjt7+voVSJAzfBuhFQb3PsP3DkZ1R4Lpdp7PIMIhwszncniR94ul
j1hf8DJzAyRHFYVDX41cQbm6IuquugsTl/21WThqBOiFMjRgqDl6OIHyBxFgPGBD
khDjyHJIeJBYhA9Oq38Ba0lgzd77hqWjf1ngreYFz5KJFOfR0F2iTzm7rnBiad1G
WGh/a0RpGzN60tGYMpMx7MrGwtX3zZrIXZ5GCUjm5o5J5UQnYa8qXo+HgSZyRh4O
lU8eyHa8aqwgUW9KWa7Ei5LWkBU1BbI8DTKfVwcOPu8TbSAfx1od0Z7ddHAxn0we
idVM8Jh2iXBspCjt5f2PnUsXuf6sqyWmFICIFoG+mOBjLmHhdwoQljt/z8p/15Oa
cy7PIGHi9kEpvuhHPpPfum0WgWGBK+EpgKr4c+b53DqFPPRahU52z8vjS2uGAgD2
MYed84TQKxX0Ztu/d/hd4+AC/d879eiTewor5J/uqy58LKX5MroviNM1lgE2e+2g
ot1rbwRijs0RTkvIfB7SJUOtZyPfqtEDAPd4vBik+tDEEuYWkTnYu2Id1wObHSxN
E2aEg+dYWbbevyCueNHZ63mmOq12MV5ZWt/KWy2lKZMRWzzHyUEbKRDgV9vUjySO
Rii/fLbHtFLn5ofjZEAvKm3TTIY8mXHQcl1+dFDSiX+hFYRzKtmATnfhzlB7ppfo
owlJUxQlpt+n5twznj2YbPZmHVNRiiLGEWIakOsC/OfyqrFjhp8SWUzCbWwR9OOP
ixDoibi4kBaRaIpytnWMBg5L7Npj1lcbNDeeobtAAVahK5/XXc60SGQaUUPtL5ks
2K2h23ZmJJr3UtdR93iZTo7583pfje4tbzaoPAmrq0L6TJhG3/ZpUlqHTAcR3WDk
onLSJXuJ3+HlKEYDEuooJqafEVsWRZjPADZje8XlM2usSOhbh+xiMKytZjKu8LKp
AgeL+OC4nZ/BqSXxjGaJPbdxUhWgBmViREQgH7sV702O7ma0+xwxvSPbo00vPvWt
TkPOrQ9ZVYvoJwqMcmPV/o681TlmjvMG94MkiWD7BEldDBt7ElK/GJQ8kyarnmE1
phzv+l2UFZZEmgY5t1AgZmyJLNCTlYO5eSSrrTimdH0YGNbnz8zyasBSowzeenDl
4ljb+p91BeWV24zwONQc6P9vBsHKRPqyRutGCf3ofRHhaRoYdz9pNYW+pErsRsFn
AfOIqod0qFD5vuWZqFEyZp/yHfPttN+1fK35v/8AHOW9pMdBCTNW/iSjY2vklAqr
2RDVyePHF+A0XmchHp2kC/Y06zOGgbyRZNtqKQ5aiIQ1Gyo3zB6LxRxDAjcJQvPs
kDVXSu8etCLKwnYasRR2GnpE8w0qt1MBsH1GJ2YvRfRC2M/tQalsC4kkcpfRyKsz
XO2J4BlDUsIVcTeYQXfMLxiNpto9kR8hwq5GnNdOuzYpvZ0PoQbjOQTKiy3iv5dP
zDK2KFmjkTr45gNJFVPk7R3pwinAT1k+nmLWlXfAAmP5Df1D79J65PR/2cTkFe4+
1d0aVmpU4qtXN1yy02ygCgeAp4OO7jCaesU9Q/jtPgoGkeXALfhH5lpyIDso3x2l
kbpY6LGOmcyqlMc0K8BEzr6OduL6vdlRtMBf7uuC/mWzUA1R+AmAGCXrUwndEK6D
DIK3A2lRY61OI4Gkorn1uCwJqzcNeLHnpwhqD1XJJniYEH0eSUaiHt7QtRstYvj+
e0qUwxkokAjQUBRFU2UW4KQETaoQl3fm28ArGGgAYrpjBhnh3NKkYhn0tFLBQUPG
nHG/3tfOSvdDjHmppMkzTrYiVajNIla7DJ/WYXHbc3BDultIfgGXKiuzeQuRM1+k
NqOL1zTsWcIfQBKMiRv7DffXj3xxXVDiy4NKPVHxy54wv4iqk17je8OqIVGkfwRI
39HOBcmzrJWVBc54whnJqA7vx1LO25+csJ7En/CQbTsCBdx2+Fy4t4kYL/y0UQLx
YTr1d9Y53xOEltnP9qPHxhaera0oS1wxCcN1R6e4DGiRTf3BLLBelAJ8NrWyrosC
/gV4gMFDpviQvB8Nhv5po2eBq8e26+v8hB3fdE5hGtJ4nKXUuTYqlrvftkr5X7Ly
5KbjQ8KJn5mKI+McWNfQP9RgaI2PprTBVPV35yAR4r85DFM0qLZ7RltX3KN+TeMx
Rk5yngm7YijGWk5i6SDlWdqtuo2m7CGAhPkc7Moz+oB4Uyp8JB5lHgV2fwc3i/8w
GxbGuz2olM4qimd35C6WG5gXIh/FEgGF9TrwrSdhrRYCkhkkfkmvrePrfrptT6Ho
SomfQaBAi9uPPBsvkuXuqyu+McoABX+xidQMACgMMgiCe0B0pq3KwwE9nfBzfgjV
GIfPDYldJ3JHIaDS/ytINnHzhqLq6aSZ1RB+3paCmiGsLM4XT13H66QZAhPQubLB
2ZVeJNctlTv+Y1cpVpJv8Fblsy4x2gvzzDXMv+APGoZ/EspshuRNWHGKcAlEPlz5
NSLoFVmLmpeDzT9rIaDGsIvva1runLPKxzJPaW7C1oAT4Lbfn2C7IOksdjsGo2Z2
k1DlqtAwopRcnHe5R96/AOb1LZ62B1ete/8INMZzyibbN0TdewFR/epqx4ti+nXC
xmusziG4QmsM3db8ynMrlWc1mjXW6Trein+FTlq+kcn45XUqozT5OukuKzh/uRkT
R/dbcqyB+PTI/ep47+/rcjhZfkfepUEf+vTp04bhHMYix9FeGmvLfy8ZOul+eXq3
3K/nc7BvwK+Ci8JA17w4+9W32iG+V1nAw9NZCR4Ncw8waEmOUMlgPdUNgERxQ6lH
7CT0Yng0Y80mDlhEGbmovhtn8u/uM+bOY00s/mh/2W+u/0x/SgOqhYeGAw8Lr+o1
xdwUFrklKDzzv46VRTQdi27dPlyxfpoEtavhFxbcSQIPrAIzrUUNUahq4nYKuxJj
heU558RFhoO25411CHYPNLatGBe+jPdVsxWZ+WGja6PI3qqp1+fba5jxfhSVi2Me
nY9C0pylA9xzUCcMBMglGDkPYswWaNAOkPc87Hbgmfb35COAJqQ150YaBKqis+QG
bluFMs+o9tB9YF4Po5lDvl8TWLQsXp9ZuC7CR8HNaz8LI/kJ1J4CQupsh9Ba5uSv
jJ0q50J9f/X+DE6I+VrR4zO/3k3BPvYDpQ45RVvuEFN2rO2QNBfs/Tt0SOLRsFCo
d9VyVxvrgZ6y1u+/huovoykSHMgipFSbsQzYmoJ4GdljQpQ/AWOiWUE8h8mTgQaJ
nEukB1TsdDjzyS5u3hcg3LCPr3HL/4A2SLoh/y7b1/FQMi556InQhEjCMb1l+a0F
AHivca/aDjN/sau8LH14Oe8lPqbjJFEZSsikIo3shMIzAQOVQJYZRIYvY8H+25eZ
q47wKUKiVsrzQCdxJ2TexxOdLmpU6sGzW8cW27In61lDb6klMLE6T3JTuiHGem7W
9pBUmo6y+pL9UZ5xqFGLt9qYWfBVnhY3SdO4ds/OruA+eZ1eGCqJc6zcgR7vBMh6
SMkD74zVXKhbZphuqKqLe6CXd9FWYRT6XgO/dQR0YJTCRqtCTgPChatdk0o8F3K5
5ki9T4jt4rkU1d47DvebKuLF1yi1e8us3JGwD+NGRbSDJdjAVwjWOCUGvpLn9Mtn
yz3FJ6FlU291rSPlT7d4qIPJDcZhQ1dCk/n533XY0TXbePNP8Mmth82EY0krrAHS
BBpg/eBOJ8ZsFHJo5qmPOsk4splvP6ZZeH+Jps5HdB0EIHEkRQp5tfFchzzZHTcj
BEWbrbJrTqFH2ckif6mKWDXCrL3upV4Rf+X/3P4VSSqBLa84ZfXCRO5Md5p7W7lj
b7BKDSMZeHhQXI5epyf2KMMbOaXR5i76hRQx+rTzAZgOwBuKAFu2W1TadOhuRSQy
oD1/oRXkQQLFu8x5Sv/19gBIRmXxTxFAkZwOwBB6O0/fllLA2cbkd3QpS+Ud/r04
1U6m2HlmTs5sbHxtJH1nxK3UYHltV+Jn4RR0IfcpNxXkmyWHp9nWQp1KFpDWTy+I
3YfLcLJD6tdvijL4um0z1vjQPyuibiXrEN0gl4uRHoeq/FveHnRyQq/xlTe57DwG
Ee7JwtAPe41kqnTkTE6LR/iWdDBJxc9H2MMXMMyaAdwvKlECI112ZMZqAKYsrO5V
zOCLgUhsF074uzcXS7BDiUSbZkHMzP8D8aQT6uYi5ubUoYEWRS6x2YFZFNEm2f8y
xVGlr65scKhVkcsb/NXeFwTAuNQ6N7awGBBSvM4cQMp8Ds0DNwbDNizdCCj+G9hv
5V55oBORlfotFaUuCvWp9hUmf5sG6wTlmmqFZ4tRYXsML0zvPAaVAmTzXz2701h4
dmY7qbi9+sQJydNYdxatQuoVa2xpn2uVUMvUbDPjuTjbonkiLgsQ6v8lF2QNTwBc
DHo1ld9t6hessuxZ/Ux4+UYRG96pYtJCx1+Tqe6xepBsgoPAKCxC5RDJ5cNqkzNS
dYGhGcZma3+gLs5MHYA/kv79SDwjuigD9E7t49BeyUtlf8OwdcLlzmr76JZo3nDg
udCCN4UF3c7ucUcU9KVvexdVGVYNFpVhV3gafdEPkZhX7M9HFGwJiOJ9Lp+VzMhW
GHyJsYvW4Aa5kGW9JQsc5QvZEXEjq6AgmMCapTjnr4tvyiwjMr3efTuTTocQNKaJ
NeayjJ5tRBMNas2d3QgOSoEboPds7Ot8rDltW/m8nUmAq6RxdYPCKpAkBclmB3bp
k0xwHqXJfxa9ebtnzZhsqNsCFl447ywc8zVRoB2HbuLkcZnLjb51hnmnOjYQzYtf
EyPfuzqj/HEmpOJEPV89zBtPBJ1AoZriehp1BOh02Jzqc25zUHewQTzJaK52qW+o
9hueMawhTwTxMg2odg+fqIH4xjoq1PYpBWQ0WQJYgQyTVWAxUwCnl+CMHMrfUFox
pWTpg8/1Z/LxSA3AxhU28UDXIkzX38eUScf96sGaLQ+Mg3ofnBovaSF7Cx7x7u+y
WD1ZY0lsux/DPmPdNt6nuh6ew+DW2izRCd+rPoMLgXQQGHv8eiKh9EA6rN7PAhyn
Qqu1q8+l4rFDTLEf2lLlDN/QFSvPXpJJmSFuByd+tnM+gA3VVYVVTrlI0Lcg6pbJ
KHd4byIIYF1yX3Y3DVkT+tulcBBHLs6DlRociaZUmb2n3tTInhyEifRMy4o8ij4h
Kc+QtrIYfXfjU4puFgw0SKgEiabLMbzw855S+iOWaXW8j5bavP3yxOh9IVAp71u8
bjtJ2AI94WAE9Y17TAa8lrhpt7O8p/oGREY3J93V/TaJwGPiZNIuAHOvtTgXFjGC
Jnxbeomp5KkLNRbtSsCk9whshRgNdTmyNOqymhYt/VubW3atnm5eIerxnPQ5xWHv
QcgLEfe9SDUiP5KpC04EwqqxBozsYQQQFNDRxywLMnGffv1O9sV5+wN5bZkWwF2+
a99JJ0UcsprTu6qzuWWUXFcFVCoNnqT92buM0eQvDYfXIq7rOnuoGJnYweXMiVKk
kws68TIVBJFJLRzAcle1JbUnn++Z3bpvek1u3eayMqcvzNMnEGw5pg07rbj+NLL8
KvjNxU28+3siGTMRGGjyNrG7Ei4fLlHTpr0deILDjhe+dyFwSbQkKpa6XQBM5LZV
yclDuJZPaGJ1ReMK47pd1L7YwEtzLbTOm/Psx4Z2bId1N4PBgqyS0k93bMz7YuUb
HbSmsCEKeDk5YRQ60CI414V5u0Y8oeJr+ktJL2Iu1f7FBsQB+ud/vXnoFigUyVF6
EAdP3ZytJ9ZYZeXeXQ9CvTvRC0I/LFQqToGlm3lcsC0fiAYeQJE0FQtYMO0yX/dE
2MFXzLi6nEevKy3pjDFZkX2JaA7MCKkcIxadCPNyJdbZUReU/1TScbPniKmqOJUy
/xavc8Z8wVMcy7E18iGiWmUD6OkoKk2MGpalKKLKNWTxzbO9MWm71FzXewDVSNTk
4WW2Y4/jmE0rQ5U7R7l6C8b2pQ8HqrR1Idbbhz5vsoy1x37/rQySofUVPizkhjlR
aF0swZuvvjjmbg/utudFp7QfDCS8UVhAr28RvbYYzXsU4x6OR5iAFGyaaF9Rh6zD
RFvNmh0r/qYYLnoCnzNAPNZrX0GJ1497vH+LPS3gnOJ7qSR9eE1Tj//wIUwV+ork
X5lBVlYoffPG0zfeW8gxeZFlhM9p9mPVNjFX5dmPwLpuf139LGM2RHQvCxTf3+GM
FHAnjup6fWkKVmgvInT7xtXFMZQ+BLp24BnN/KxVbSNLVbJ6JQWSx9cV+w+v5UlP
WrUKl38WMdROgMe0mxrUTU5v6u7W496/tAPJTIB4/FyGPnnmrSXd8WVSPc+xZBGa
T4vzSeHLeFfTCHyqTGV3Wio5gAUM8duSqy97dWwZOVRSHC26Gvu2XmrDmqQY3qFQ
4pkfIQZbHvy2Gq0uBZiVazkQr43j7m6QeKMH4dKe7zDYZYksww3Jm8UBArDKi9p1
PM+mjWfIwV9NKm3Ct/f6ed0TupGd+5+4wNtPyjkr+11a6xFmrEYoDBdoMjCsw0fx
6zRnKekQZN3l69B3GyWI9c12vXc8jwYVL+lI4Ac4osAv2kwrkFynomMp7s+AdbN5
O5zaLMAH43s9+LoCi/edO9Iei+jhPiYBvdTIEopS3e7/kdE9zd9iDjP6rx2JpcHN
JnFnOcWn3i27Yp2yVwb+9Rmp28RxCPh/+xAXL5UjY9AsWlovOtYLlVQPdjHvkDP7
YTMJKYQp2UjGgNMLODnMMo6bbtZ6p1mWHsuwlrQw5jYMEl6OjL+cdLk1p4yJmI9e
AubrUQ/YI6rAhZMQTV4d7WLEO9UadvKVqP9csvwFyXw15awSj18LzNZ8Gxqdtpt9
du//HeGYgBgQs049+dsbbvNdw/uonmA+g3OPMeBrM6QfpKgGQm4wKOkEwlX8uwau
/uDg7vAWLUmmTzkebG0TIeuFry2tLM1oNGSw63jHYYrIs0WK+w8kz6InK4ASX79k
4kLNBaUOzx1Z4nCkf0P5t/jJQViyt5dUr9IBwJLgTv6UFYEgozY5ZDfETKU9uc+4
YXkzBpY0JkcPHjGEdNmYhBPNEov1suWeQD2D2XvqsjypQhdxBLdWaUIs4FVOgWL6
bg9oVyhQhVMgO4nkArcXChPJSK3oaAso9/6z1GQzQ0wDkav0qKfMaTx/udz0UWZy
hgn5MFEW0K6ofBG3VKz5uGkseOydKHqlbcsmLYNRe4NlD56J6zDDvn3uTFwOIbhO
1HBr6rVNoV89ZWC/rw6+a8J6g7drqff3ytbQgdM8UM47SgfPa8J5cVEXzeKsN/1R
SDOQXngQEDJ42CFpGZpAhVRvxw4RCwtBe/C47/qi/p1kMY5NtP42cF+FVYv5ZuEP
4PidQ4XZW91c5h7WZDbN27+5VI0XjIT9b7lxM/3uhVM3C2JH2Wswm2yttzzdeZ81
bK51dsOOImmU/ejvlPcsuH93ZR3wvfACEBNh7c4lMH5iK7P/R1RIqGZsHv0kVmEo
9dGQxle12yDszXCkCV6UGzww6iQqy3yN7RvAlC05e/gklgxVIIm6XgNQ8S1+5c+S
wul3lVDUxL+2RnRUcMSIgHRgiAZzX6MIGgIYgtJcMiYq5nlpO5b9Cpy2iGCZkEPt
Z4nJfCKNvIhRpq6Wbm2cSMdEjpYS71eciDNDtof9yCBsZTRR+IbS7eaCQsHIzbQQ
H0G9hxWbitOeiPjA6a2RG9zYNWzGUHCg5EwghgbeDgcaOGsOqxi9T6uiW/kqBeNZ
yL/s0aAhaIXSq48nrK4o3Ci6OGKKB1YUDHkr2JRv5udowaIt7cJvf5770i1l6pM7
7KT9s7e4uwMEYV7F7tzcQYMsXQKxP7TRJbUtt3eowHtU2obFgwTBT3NK3OoQIPRA
hin6z9wgqJct+TFLPnmU6fE5JQgkShAuxCfrr196cxLx0lbw4FQNO286rNGimj5b
rqSRNHIkpJtTcbj8Bd6pRz08RdL5NjkZ9iL9IuJmFdgkqNE3uKCDERwOINmFuGn/
hz3RzaudiUIV5EAOPR8pZg1c0i1G6bMNKTDN4YIeRCH+yGisP6OWdlBTKhHCNAF4
Q1fbycsWNhVMQ/azYhkZzFcSbcMn4gu2L30lznnzqT11fcTRmnV4I7/kyre7Fahp
ubVr/uYqitLKz7kKe1u9ZIvXcr9/8v46twMK3I8W1DTISpfuzQHysuNWwoHW7qTX
NYIu6sT1hYRF1NnMup7gq734jri8IewqAR0zvJrgm99/LSH2SfyGO9anwh0e1p+f
OlAKgC3YRjpJsZPmsCDBTEp4jsn+54mkAdPFS2Jp770h0/s0TowipWUl1L9KUmtV
X8z2j5gOR+zVyf802sIBJ4i2l+fRr2bQ6x6x/DcGTSQO5E9cdRxgOIgd0c/bkNTQ
THMRpeO3ubZEY3WxurNcntG20PJXdXycH7K2mCjXXfHZwHtpOKeu+fAPPZnl4r+d
NmVe6hk7IbsqZBNEZ9jJovazXiWnXIgBOAW0DHVT3okKk8k93O7bTczkCq+/Vg7P
EkiEp706CBPkwWNqZQlEl7/K5DAPMuFIPL6zeU1BF74H68UJu9IM+uGoVp9adp3M
RBGSf+5Js2VPHhTSw3IgvAzyCe0o5gLNXO99/WpDGxLMG5j9Upit9316TX6x6Eze
NtuTEhw15wLJlGZKIK/7fH2FXij9/sxrYVPLVKEywACJxdFaOJnOZh/x8hZjqgD0
cfxf9+xJJsZa8qxcUNLk4hf6yRHlt5Sf8xwWIzCE4NzUQYXwcOhBvyXlsVFY2dQL
pwEwWZJnTuScRmRL0k4VjgTOOpfmFnHdILbME3mY8FJssu5ybK+e5U9DZurrVTkm
MsiGz7pFJEiX2LW25wi1gcq609ovNFXxmRkGspI94k58Ru32SNer7q7R0N0stGHx
mxrprbardTwz6sZqs0cb7wEpTZVRNPqTkRR6uAxNcHLFbLZaQVMAyw0uzZ6F4zho
BmH1BZ/HnRrMxlZ9SwxcRzwPO5O3Y4M82H6l0ehIpXY51DHpwj4m7rYSqqh/6Zge
hp3pc65/YFc8GRhNUAJIe4246CaUdw9d65p1M6rZOTjcKQxCPdDKa37vFiElldk9
sGGKYONgBZHic5lucwntVlu7sMAFJ20OSHWB32gSeab3rUpxuKjXBuiUMtbe5q/R
GcYZPTr9adBHItCejNJIgmZlTezuOcBNc/cVC4ERqnBp4TijtleRAcjY9jP2W4s2
lGa/JlNGld6cvrTJDrpR3e64HC7wa/lRgqASvjAl+QI4POBWhCOMSyCA1r4ywf7s
NIUcZRenGOs2ryKAubNkJPgspQBzsbfIncTII4odXgdPiLx/drvkz6CXy9J3E8lV
a92h9c+gDuQGMsi3BZkdv4ZJNbmGREYqJwDIVuaYEsIq4BFlA2xV0xRG/NK8Qq4Q
EI7D2hCeQhb1a25qAZJA1QT73CEdMvvOX+tufqGiWbL3SZE5z1Paod2DWp9yQpqK
reoZWexVUH/yEW3qHqZYWp7EI2nvvg9NrvZFRCBu0uyz79c0fNfczoBmRRkw+96k
cp/1SBU5P/U8G/WDetjV3qXk+cyOlQbPnRVqHchkcvHWQeGT0DTmBxLBmmMYIOxy
NjnOjdOXfUFAkJ2dbkvmylXViwGVYC9hWRhz+A5Jnn2ekeF5zU4XAEC0AvhryVZa
LG4h9RiEpFY7B9Ggiy+ubS+dxS+d3Fr5yzZix06eHsV7TFvAMweGOsvHYDSHoosc
97rh4sOuZw1BKGw/yUdKv8GEsUAETor+cggZ2LHGVHiMN0TDnLJJ8l6Xq7usRuKS
JagaM3cBy4KOuU8T8+UU3dNbCU4g86wcC2mGsDPmBJW/v7hdxjRDpqkAKsbXHLzJ
LycpAGYqFIDjj9WPSljLjE01J+oeq0fYiDwTv4urkmHyhhcyNdomgyQgaq0NW+n5
oP+VHXrWVGk82cK6xa0ICZXK7x6HLzb0eL1dsh8decVMHoH0rgBJm8H+13DBXVm/
mzK0TLG62RDyW1qSzfY2JKSUsJTrg/d/uSBRNt2zvXxfvBmbNxRixMZf/ZJPqeqn
EvpQYM255uxE9id+SYZmA0kA8EVLwaQHF8Y0eauEiqKKQROdlgwwSms3/QxvCr53
zds0DI7yOJlCpSpAxk9bO56WHnvpWOkCMc4t9urhjb1IpGA4f4FNmnCBroAio5gI
Z/kbTKJZlNV+kD8yQtoUPxmWoSg7T/FzVuKZYpqo8vWpmxiSXQnw/LdKIKq7NY8S
F5xRVF0LPZZvfTPvMPGWA4q7ZW1XoPylp7QGq4I1x1bhswGBroU7S9A9cgnq3zIT
ftkl9MRgvGdYC6T+5ajP9Q375ckgDoH1mW3tqFIwKEKVHVJNp1JegSFGzoSbE1oS
g8XsQezFjFWcXrqJ/eD9L/BPh+xrTpOfsl5GIDHIwFqo9brb1XireLtsxip1WC8Q
vZiVJfTLblD2Xp11p/dorhBph83cjvDy24tBQSv/QHbv0bDBwuv+8nubEHSMcDTV
M4KfT9DTPl+zlCxL0/ec9WWES5eNh/b5XLXPYFmEwWYGaoLTb7QqonarjS7N4ACz
xYSv+EvxSJFQ48GlIOaWtrabRVRA1D7dfgp4zhjWUdoLJUL62gpbp0K6PCc1Lu7G
sy+MowVQtc63imRYymgrNM+rc5A+GsNCr85ZR2C+pJYflb06XiagkjFbLcPQkpNG
xeUAbhOa5A9bxNXZVDTs6fdYxp+aWN+l7fPXEoN85aykOOwjWxBeP0oXeftmQP65
s0lMG1PwGHhJq/uI7uJ0IkukhBmLmuRoODm5fa8+vCRcYMKVktLAlI4eot4ebeL5
49AfX6Oxg6SZ7XYchid7Ax/rHSby21hEiV2UkSEMqEdO5bnCh0KCQhotOh6yPRTT
69T7PxLaASGEh6ROWaFI1jel6A96RZmotiJ0L2oLzNb1HuVIJW7gc08q91Jxl533
F3VTe26pVcDYLOXfKpHHarepZqP4yi67ghP9tqFVE7o/FgIsI3hGTzUIYsOLR3kz
k6ZNpjNO4SrRHQus/4luSBE6zfPtg3m5SU7frf2pwonFPBt0ihYO+3/zi7ZfLU/L
WX8US5LxKZtqn1cmFAIWBDEu/gWuPNcSKsYlVb2QB84FJ64y+nSom78vyahICYA3
VERvEhO6WuEbBuP68j6TIj3SIpt7x3lUGBshUv/Vh5yM5PPDEiZS22Ad8l2co2Z2
qzVETwbqB4J5UWtdRypE4CkMi00x7AyKNXUNFEzgMJNrZs3mKWx8cC4bhF0WIZke
55ohuphDIXCjj9jszEGRNVYZi063qSS07hwTs+JbSHHpsXVHhelDs6t1kIAc1lJn
Mqg7u7XG8KCvtgcOc78HWQ2OYmPAseS+Zxqo1Og2oo5kzKLNCWpUHbBYTDBmRHXh
CDBe8V/ZXLhV0cTGljEk4F3IMbRpcpjLkkfqSyOX80uZQbx9SxDqySZ79mq7GIXP
ZygqbCD5vdlr/L4SizxneP+9dlYdHsTsGSz5kH004xcmiocqdZYvBnlsE9dzu6RP
fO7l11p1Z8778UfIzUSk+elm8c25kSqp/9dzfCzF0Ds05zMwcHCbob0HAsM3AXrD
KudLoRTOxAyW7iN4/yirOKnXWAJOs7m/+xDZcc3B8zX0n43Qi3GsxfWZ4lE4lg0d
Y1a+2+7fwjeB+uGF+t8LyZs46a8f0vD0YD9Qxfv4WcblZZ9ldKic04sknIdtPiLY
CflRfI2aXiIdaGOBQYbqWn1qlt5A2As6vWcf/BDHizEBY0/IYpWlIQHPA2j9Okuc
4kduGdcNHxrO98tkfGdrbCYNdKTLzwvpSbU44izPczgR8noPX3UIZ6RUbZJDJWn9
LYf70eeXtWrWIVjtH/NyIV96inqRwvz/Fpl5MFLQ9i9+p+aRtDrPSyNcKO5E8JLI
Ly4QGd7qBtFOcMViiFJp0h7kV0UB9tJj8wDzmke+UkjvPgziUwDkpT5cVP2g2Ngz
eeNGii9W39wF5heMrjs+kpToeCmoG7koTJpjGAZLzrUbWe8AA6b+xdqLaLT9g8//
p2DBdC+CXPXtLa1MHoA2/JCIHwjY27T3L+fcnVPtHaj+Yudmmc/HYKxMs33N4w4O
tGoy9dGcAIqkLooeYt19dESFb0B807HZTVrpdiBZwrh0Kkv+a+dbd8ODpUntIhSS
1v/I7ehI9m8RumXp6EYJl6bVcMkVX9r8FSarJ31GUmnGAl7MOi64rBYPMUkOj4wy
6Ilv9Qclrk0tf2n154ywjMkN5/QPhbQrIuZaVal8xaBuDVk9NBy55X5FwODbAroQ
MdngxUzIuL+xwsH+6mfrCtGfCxd7Lt9MgBRX3zyu9ulaJR9dTq6AxwAzkp5TA6sC
vdeLFKGo/KIDj7q/TTwQepUVr0jgJNlcmF4Ek4wlHGDofzhM1zGglK+ZJ+aKbn5+
S1uWWrViHxXGuQIAOIzyqjO/yHiMI4HbzklcSEmEE5LNFcek+f5hGe+4v48wWVYA
VvwfKLE+UhhYohb9zzDHcZ6Ep60B/j0GTdSpKx3ax28Vx5oDaDGZG9MldrrYMxeD
vGMc50llt+UqGmD+VUgHlvhR6gsetOgyVrCUwp5iRxlnhNQeAE8nZnEkcRuwiTc9
XUa+zA47TLZnQhTrc2RO8TFZyr4pT6cx7NkYOs2BGBwOd1LliPuSb6PIl5BDsmiR
mglYFe2UtzZcXbf4CPDlxxdUNW3U7jfy8wTO6kYeBmZ5YqplpOnV1mZSeipsUTmP
pkJz8e9AoEzBVqcPPG9IjT5cuh8cwUPB2Fjgi+/pnakYok8fOyt/as2iqcmtm9Fd
+2yRArrA8NTUS4pfyTgGQyMVIxdN+xEfn2RygUdBWOD7o7/8Wa89TiYjTffENNlW
IcWAQBnf0/dDtPWtF8EDkBgBeDR5PjVj5/yqsFQsYv9vr4ufklpPmz1S2jDQ8bAg
SVnYbqssfhlxJWF6rTT4amZGQb6I3kUIrOed+J7I39f3S6TU2RvcLfedS6Cf7BUd
OTujiqaKEoMa/OUmkE0cRCgS0Lc++bJy+7r9YTH+yTu1lftda+LSZYLjTEp2zX7h
tqoL4CtYOukG0uYwpdHV8yTtEheMcT3TOZ81nBfYMUz7YAK9lHE00Y6KpPHN0sx0
rHOXXSQha2/xq4GTX5DJf441azxjwUgRLF9gxkclKJA6VbtyEwgSEnRhxvlCkq8x
PqVzL5wKW6qSxCL9jY1QrWTtUEeTBLEP9vdCG5mdIN4pHKaiP1asUu+V4VqwVsPl
G5E0G0QiaOJTa5ciBHjgik+WgWoFHKAmLiaDIUxxCCKxKK9DldgGxbNMtW1TIb3N
pVhgakWIb9k9rwU7R3uDcV+KO46m82qa3PDO6fYu4kPusrm+qN9p+fipfwLjbrOd
xASwcxSpYPjH+EyM7mJDzRuo5gajGn5k0HMJD5BCyiiJ43rXkiqB7FRTnn7iiWbA
z63dws9F7uAunRy3CI9ED3V5Dp/m4T1DZoFM/GJUkijHPZtpSNZwH6e13Qdxjnwn
YORozhN6WOISkN48cveNgs9j40O6QuQuQkwK9ZQkt1tKNic2brtC9Uc99onvCl5r
Cld28+ZfSFoG8aJUEZc/dDfykK/LtvMiF77VO8ebZy3v/hkoz9MKfZRtC5UTOWlQ
fPGqyNMSrSF7NKxUTuaV/b75jjg7t6u9jBLh0O2YoC4pNMCPqfvgYVRqVDgITvg6
t19Kjf5GZrf+d7OdskvAEBlOutBfp5dTQuZZB9jpYMLQUaVRjo0kA4lhJ3HP6I0Q
DKk75OHdzkutgRLwwqPORxTqtEQ9Pd1VbMR9Gith+c75cXpwwfLWxxuCoCOVbrgp
VpEvQDJDZuHeE6gRqNwsFOTIwDfjG+JHgGicK+GyXEQVjxyrOBUbPG7H0/XzZAyS
3zWg48HDJC9mxp7LdV6dd+lCC1XEfYGznb2YqgEMqp5O1omq0yF+5AiKkabZm4VJ
kvrCRUKcONjv1a8+SecEkJEHXzbOIhqAkVhSNkbemlDS+URJGNv0S2eFmwBtkB40
2ED/d9f2a94uykfmfISnFQVvK+IySXjadi8LQtTPRASTl3lI3h4LeIvfrAze59F4
nal9m9DXfUlfPXl7MCltZGC9TU6R9G/ZGYtsTehbhdsQIwHFHRjPYRDIGRLJ39PQ
rY5S13ZzSuly8aysjkN+okAjGIhOvZEmHQTpkY3KGK4cTrEdNYD3YiXp4ixKPnpt
VY+v5TuhjN262UitSGKtcaMzSZ4NMC6NCEk9x9nzrpc34JxyZKP69dydp4yP8msM
9HEN5Xx+wfxoWlhtz6K5pHY9AcsTEL/cpA62YnxtpwWFTIWl/RXc37jG4oyVaDn5
0op1857RvGtFqs6imGaWDQ3ZXrSRWFVyh0za0z2dlIBupD8emZZ+PtJQ5XoAbhbR
EaYl2rxpOHLacEvjF3Ndc9XDIW9q74tmTTUV7YM2hhYsJpU5ptd6h4VfkMlPNB5e
w/FDr9Zl1F5GPVr4kkinazTXOeFDeINtyTLbAmi0wDKlpOqgzPAqOgpTz3j0VJsd
VFyXg6VjQOqNod4MIAWVxjPvnkNtpXZdB0yNBlPv0xb53F/RZNjp+zba/9yB0wUF
dnLB/DLY+8FShb1lCn08oxiaGzI3rLwuZ90bku76Q45o7EkNUlTIs//EbN4Aw0v0
uE7t4DEBv5fg2MVu5toeaPYOQbh3vxm2eLVSZmz5IjXDTV7rtNSP8fuEB88KoFIK
K7A6HU6ZkonSNa51Y4r3MlGDVX1w5n2zDfYUQ58M8NmYj7SbtyU6irX/YamNUSWw
pOTwVrxfDVC8Q5pPjzIygjsRcJVZpdgl9vI6qBdChp3Hjt5mgXV2pwNHYRqktVyD
ncKmeIWrZCzySmeAzv5+t7uC8Wca0JeYxuRlEYRk8ctkRBJL/APSe7FaI+8M3aRA
WqHmP3yyVQhXv6/1ftAhervdJ0JhteoTLRHVa/pcpNkVJfY90ZDbqfF9BBGyXAXi
0DwgUK3KRjN+NoQK3pya6/3lvH+j/cJ7HsofdrdSNp3PmS3u+aVIZER1d5/tGkGU
IfVsCDbWvylV5FRPWAbeEZYIc7HF/iN0WuAoE1zhsblpY/waQViAA//tZwj3Dvb6
bdRCn4a8AGnWVKtL8nqhQZWqCPXmfTxkR33BA8zIX2pmDsZh/m78UwYYM5MLhMKD
jS+KadC4r9uTvsWAMtNKanghNoF094uqJArOL6PXblRcuWF1nhAMUgERXMD/qVgJ
Qj1WTaNxJxjIi9ab4w0xPf6nIzIO4HbRGA2M3jQfFYNdjLoZ8D40MUUpnUZn5bWE
8CjA0BoFFoYIHHITcGEt/MLsj+kq9ISmRnUJl+9PFh1NJooZWwgzWksRrGH6q+Ws
hN0PoTUhOQdUYRoyKXmPF+ayBm+EBMXJVA+xqnnZKrj7ZwrcxRD7DxPmR2EGZsg9
qd5ttxWcicQXW9hzGRCKLjhqi0Vbwu6NVcFjfAmQRV1vaJYfURMzpMjkEgFterfm
OeDOkr3EJY5YHLgva5PQMtCFYuymdiBb4Z8hjxfcfXS0aOFtSBJXS2CTNSfdfOoO
cy3c70mOt8TWR7R3L7A5unXBx1RYGyPIUL284FDvZvFkO0JpGuiR4uDJr2X1Tl1t
Tk2NkJRIICNru80vO2EfJN4wEmACHnOTP/C3+jwNO5pNNyXkcZhgGgq8cFDmdPSp
OPQE81FVqy8rfD0vyqQ9xfZXRc7+ibrN27TkwqU53tl/8ptjbQ6s5CHanBZy5Hke
yPSSodcMPtlMo1R02R58c8jDddnY8EQSZ12ytVJ44ifrCH16qT54pWbtkvgWxev2
vhbzVGpziaMBpgkJzhvQTUWmfbaIMy2b45jXqhIiXKqZ3ctBLBTOSmZpps4hV9k6
FVwkUNunerrJF6lLsAv68tCUcL1YPS0CrF2M9kc7q9c27yVNRKO8eIVh/Z1fHStk
oixGeGMt8GsFxhObqHc8U0lScxHIhtsIBbqiiwnVHCDi2fjQnuUneeozuuR9XzAw
CQJ6Kf50x/TiVIgPisLyci6L+KldWScDJJ4YPccWavAtkRJ/vGgx1ldNSODCwHcd
UVjiiFpBRAHP8jN5e6WXUC3L/IhevjzyQIOtlReO/kKNqI3kc2KMYq5P0S+edP//
ZYY+HXlQ0IZEaph+VGDU/oSBnxpufO2FWEkvlMP0cII0f2OI73S2MCSiPA+jfpvT
d3EMBuwp7WAd71KTRTC9xbe0CpAbitt3FFNJ+34iEyrESaHbI+X+kC4H//gdwS7L
s6R83eAqconymCt/Pa7o+O40gYGYpomdcnQQswNLAnrQpiI81BhtrebqSTJXCvzh
hS8aFbF6mgrIl3wIHogE+mqImx4BmaDxBOlr9fPNFgkub3FxSDcjh4Z0TrIeEadt
4pPw+5dXQD3jVfj7NyBXpQCZRHXgqZsLNj3vumZNzWhucHFQFhiXOMY/cOJWTmlv
4nSzGpBiIRnLuXhpAN0AuVoGEL+1mOReESfg2/l8C31MJ/EgBoyIVWoc86k837ti
uKM6jvXj43dKhBBK4/FKo0WH5tag8hcP0FmZEYdKYr7TDgAZd1vqTpEo9Lq2wE4r
moDhMu/7VPGT9b5b2O2Vz33o154BZKOBnvmomm/zcMxqxhsHaLSJUQFQmsIZlAib
H7UmqlbwAA3BhCYIWKibImqeuxcrl6d7tCMbW2CQHAz0P038Q6u2uOFytPAlR6zL
2iAEkBxigAzyo+GMG+MTezlY5YfE3hIpWTOZvigEvC+Io4Aa/UT3YNWv/hbx6w+j
0XvL4uzskKE5Q9QetKFq+VwkoYW6jnQeIvprPQJcYcu3gmL6zc+WkBeUKMxFNn+z
o7XaA1JNDtf6dBJe0RAq1RXo/GNJhN9Hq3TG3xgIZKdhTi7IG1ZsmOdqcE00TyUa
TmoyWoUySIH0XHrZWelsJlmM//7fhVB6G0oHnmS5duzspnE8f/c7OZhrY39ihrSd
K5ySgR0gl5GCvenzsXGztSSXInFRq0dP4sMWgCLlxUUDgheNPFFI4pg0xKvThgYG
QyM40uukaBt+Bfyg9u2Zfgk0TGds9fQa6KNAKg/QLfM2v9yBsT5U/Xy74nndM68d
Sn18be5XGujlL4pgYiQUOFyaVfpybi8oMpvUHhpVYuOF9keGdyO5u/nvSy1J+CNK
NzUVzRcQUT9NKr4mCqiiPfOcxZsZMMAbWggdUjO0G8lG7Zxsc0GAG4bOqfeA3Wr+
toEU4bucxy1u4EgfttyoDbX7vAEOgRRLk0cPI39Ve0XD+XQC2DZqaH5JINZSL1vv
VZfWHJuKgI17cuJr7MlRJ+Artd87QYkxF/7Inxrd3Tt+MEL8fjaBtosRp05o/Xbm
EqsnIuYsplE4Iz6Ry0C0rP69tcJm5fGZuEzubvWARHbLBa3N74m99zrFRUMYs/WQ
+QROivpFwCYnbY22smcvTJSJVRThS4eCrxXb87M9m9LUOw6Ees42A4BJ3ZGfMJ12
kplR3JkIwepsqCo502vwLh1cAaKwDDq2gHaYf7ijwU27lvQimj8M6iQATONa0pda
c2x/Wxn3WpnyDSKokJEDNXVsKX7YKKHDhkbriYicF/uFcr8vQfMKEFLoXtoi2hZ9
5xSwP2oIKZ9CMleef305x8wUS73MgZ3OiuSwYQt/Jgq90/3CGNbTtUUcki0I1kXE
MwezYYm87/o76J9GZ7GQ4A18OJ5466cKNyL46Jl2iRd2aCDe/TInk1shr/KH/89d
UgQqCt4RIWT6P/U4q+pYmYrbSB7igRzqgCNrWwaZ6N+ql23gqqQZNpKP83v8JCiT
xL6FGsNyCC+8OhLbUYbP+a5SlztQcEQC5AYMiQSorbWh35rF6Y/2GYQriveWQfo+
U9BF3NmnGIqxp4lG57H83tF6DDVHAVoHF2gZzasujgT/nSoHTopMl7i8lADSy6k/
HDb4gfO/TvlVCECJ6Z1nFhIWsvXYeDc07kL8D2u1oBlyN1xT+g7vvaR5ei3MBdYa
xQeYAkERMQ6mTNwwhqgGfDkbkugdB8MehnWMJ/9gspcwZrSxmj5Iw0lgTqz4zPJG
6/Es+oLJv6+MkWH83NteSWklbt3RuMtJuvdbEo6/KQoTcc5OYHv+ghZOLCOtb9ki
96/4UjUh2VWa1CxyMB4wN5Qq/8B52XwBumWTj5oXLIw5nN2t1fss1B3Fp9M0n1OE
Pzv+Z80eaEN7oDf5I0Nz5PbVdwjd8R5lfzimKIXVLaHGagAh1pVKgJBZ2OEfo0tD
FzUZdD31TLrRIbhtWcVok1yvAO0Kjk6g3QUGYOb+h/+21K1WSZ5lw9ySwsmYys7Z
mDZia+wRgBh2S0GZWwyMZsBvLr2GjOdxHjYvn4Ygs3hTrgP7WT+SuPHA4woh6gbe
Yhc/eaWHQzWpjREDTy2fL2ifmGOplzc6AJhF6WYsNqqYpMV7O8olgyrcib+a6L3R
NsaBqb6Sncc19uL+9b3OIGyI8kXcsJd0L7ODJ2GgOcpCRfrs7MpLObap1jyhxEC+
21drMlKghrPt1xDAXbi1Ta9yz4b6FLLkbPhpUf1N1xAfc0OTixILp2iFavadoRi7
Y3uSTATGmUwA13gN6FJg0skNjSe/lyXQuuafBmJ66XQAWBG8jSWoZjRorX+SWzUq
tq4gVZSGG5lzICJ36oTq+XbpOLOERKBXhBzk+H2injuhifg7RRAmJE4IObuvVkCi
o5dz/3hSRnSeTcYOChzrQkipOGK4HAghaqO21x7FMZTv8Ds7TCvx6Q06XfRjultd
+O9cJAuM8r/ij4zMt8YKbnYjFWCm8nwUtPDyCz/HsKK0zNrXsgzcF87yV/F+fI70
JzhWXpGqHinEGxoGDmr68VQcxdMP00UiQXtyBN4BaYJGZcQOBgCf1d+laluYltm3
wSczlRIQVEi6e+bFj9Jhy7H9i4Gn3Zin1iSlpS13k+SgoQySP4Tw7oMaPYyBgzlJ
pgg3Ar3G4IPgqD1qd/QlJa2Ube37Bqud9+ub8TeGNaCum5bQSNBugZIY+ZjlAC6y
CXiZpF186ePtqLm5ZEAU1VGBFIFQaFEZs7jjnneP+eWeVq0Ejl/+8BwGI4fYOKat
5qXcEyuExf/cBHb7T3/H1W1kUDOkF2hGOsUvJW5GDALp3PmBNkdXA0UTRODS9OGg
aqF87v1a1sZQY+SLBtrGX2wbm+RnG2LFzA/63OfT/5lcIr07+UbPoYA/vHQZ2lRw
Q4HhQxS1nM32di1kijQi3Jrc7/FStfQJtCfhALRoStIVnO1aVmkO2bISYDxfOD1M
XwcdxVYpUSgD69d3HXez7P8kXNLo1SLJX0AjSkIjylniIH5KwxXgEJTYNMmadGA+
su8BKMBxwPcbJi8cKPcal2quKzYMZgjE5BwSTUOl5K879h9cHOvIuIe8jx2pfc5Y
1hdJ8ZTwHO3mqXCXiYI7wwZK+leQC4eQlL6rynEBLffWPAtinND0w5TwErkhQNg+
IcRR0wn1cftEpmYr1yLnETBEDR7inJ5/Ex2NLa4UTLmctLtmC6uqVPQDH2p7IN2u
elojZiD26QpnUA4Loug7v0lQegPFRAgowFIn5KBCMo6modPKRlr4Wo3jnXO0Huf+
7pLoXA/+QR653UKVbsG1MENzgRLFcPsN/PHLz8NyV5pV/DRJYI7y8vUkRYrvRdTM
Twh/IyTR+H/SFgtMyvmaYZlKqsp1k5QKRyu8TcDqqUnZrcknts9bYU6DX7OyO/bZ
gCu7SQcwfK2bmgA5Ng3r1fCPelmQs9okMLC0YcYVhiHqPf443OKmJAP54a68/RVG
4YXVoVQa9eH3mTAsbuWux2ncCiLX9i2MxWmkoYEznLghs2siLxIXh5BROGBR7fzP
Ys1iHckwCUuJvtzMAWr/TKG9tIDfY1Xw2L5mEk647p4Ts1ZWnBjzMSnC4qE8O6Cm
/pqY+mygvAwrU3kEa3NDJTvXV3Rsc8jWH/OVPjXl/43gbSAFnjvB6rYLUvU8qgWC
MvfbBqmQNMBExxXX/rK4C+RKcvbfGIv/Kq0XHOBCiUXBp0oEZfnezriMQny2ikox
hsXfzSnCj07Zajcj13uQhrst7HWdNO4PSAWlmwTq0FqRcilrFlRfFLKo2Q16MQxU
9GQlamDvVRwCMYWtW8zLG53S/ZWz4tC2C3xfw7N2ilIOc23X2/3fdR2KsJtY57RO
yY8wCUJX7bkHnd2zLHNXL3pEsme3KbWpKLnEZz/t2PxzdCBXoPaIXGkBhRrjGBtx
095YI9c65ykjNr1GCmsB0EEt7AenZuf9/V5KMjhM8jxE6Bfkos+QrjRt4WFNJzBa
MIFEuEj9u7Kiw1Zgac5hNz6yLpAbAeZD0PfFYIdd5rtC8UTtkINO2wupqiWPDLPs
ZUjNVr3SAwrArsy2w19orBG7xN/m9mS4spj4BSrZlWFEN3D/Fz43jJcZkSUY75N4
xdwpFdG1P6AMBcNJhl0PTDA+9qDEMm0QhpV9LJjueguRtT+Tw8uzDM8fGOKxELyb
yDB0vVCawuZ8hTjUKWiFLKSqPM+0hpKKwrG75uAnXvohuWXApOoBnSo6c68diISx
xLlMCIjet9xjAbWq8dbw9EyZ/SSLXs93LIQW1Bpb/ECzfKbgAfR/SiHeqeKKsCz5
EGSOVB8Zvh5+YG8P+PV8yFK7V87c8bGgIwA/QjrVv0MeDzSy+k18t1n1/hAcCuGr
2LYd/cRfmJN4+LG/QL42F/7Am8MXegdP6Wu+K3FDTSgoy4w+fxE7s1pyF7xIl1j/
4GUOO3kGMQtfLiIGEx/4V/W1Znu4Lf6F1eVpPqvpdoNJmg9lRCvCWus0IH3+XARj
qaLOyynBOMdDEYzvPiNLFDhQ23yYvWaCQ/Ywvl50LdTXV6SVeoxqsZsIQYBGRjKl
x5PzHgzpqFflkGyOu5OfnykaTMfN3LFUSKb2cPFAjiSuCLX2b+7Uf8PpTBdriRLa
YmHfXuQCQTcS8XlvbMsVpxzjZ8PVPLpmnZfrEtWW3G9ZdLiLyPLPqr0hXvPo0ryy
/ntolfpzK1rBnJU9KNhi09VtyajdnKPgfiuGUW5mxwbg8UaHZ+PieeRfnxRpmHvV
hZYO3/wscDtqTZXCLIJKjRFoAGQBFtiIsS5InLBtWUMQ6NLkLvUU6DK906WleMtZ
fRPTUfPMmd0mauVAh5v0Er8H9ZFKGMz56KV0Tnhakj5vclv6SKWoDJBf3mLpoGN0
Jrw438SEPD0JNeAg+7bKUyr7kaCdQQZJubHV4PpPqSHAwwhjrhcYT1+dD1pSMFIY
lao+2tpVYQoYioqC5uTDxy9jnai904miuc5fyLdFu+ymyeuno4NdNB9dWJx9H4Hg
dlTk+TltXvkKtSOUpXs5Kqkdp9/XdLuhqy2C4+92lNif3W+nr2SgoUmZUBzQJc0P
7HpkBeiUcoi/y+83uWTXl7cHrGwnhYs7DarqBt5WGxOWq4p/ZzbSwivNOrBoxK4t
AFvh0oFYmSqtXjIg1fiaatjMVFrGU9bzk7Q/SOKOKEtEfTffHiODKu2Ruq8MPavo
unyljPIEYtI6l6/AsIVPbFxz6hUuJ0nG7iTgtxgZEsg6uFH8yoAXF9b/dIh5hjOY
tAIhbz9c87JiFk6304I1yrqzMaD9Mmm08+oy30EzqxaeGk+vlhIWRipz5AIVkOY1
TRHeaYA/HHsFmdeJPPmVwBXMZ7R42NXLk7CIIMRZZzOdqF3fnp5tYqt1gHxmjoAm
T/L8m4B2hDrqhbxo7yoDcAXDlsKQdErit6QrWQToyvygnB54wqi2J0B1239ayknb
CeRMNfCcae0JVLxxt1klBUAGGhqvEvA6Ov7eg5tabXI8p+nCKW08DZvrXRLhfk2V
iTp1RCIi71lruOk03QqPs5jNHREUtCdMb9bwssp5ccYkY4B9O2zs1eUi4mz60a5J
qLOaHXpo865RObUX3YVNCR+y4mG69+xu7vSUeSvGXTbDVOxT/8adzQPap/T8kkx1
Xnme+Z20L8PDqD+i8N+65yCVUIWl54B/iorWmyPkEMdDUATuwlw2aRELCCtA4U+f
wbdsLsaqcuy4pLD6vDzaNS7OIFU6Fr4Vxdj0RFh5rwYwQ/fyR+lbmH7FKX9h2gnp
kkpNAbnmti7IYAg6gF+yjTDKhIe2VBPL7LF78BkovJGK3H5bYKMDy9JytDi+siY2
4kR+y+YMlfTKfAOwlZB+fSlKoo2Yo5r2TjmJn+a8wEmEMIjEaXFwlD+1GqiimXEt
cfgedNwFTIzbZ5uFTC7kcI/z52cbPXFxjp78yt25pN3wYQTL9XC4J32teyilfx96
TOF3ILNj0MkutwD1bMIsZsLFQERaDMd8x1hbR8YyzrATAZEAlUsq85XxOPQHvJ0r
nyv1kcUaVp3bAKtAcOq6oQ==
//pragma protect end_data_block
//pragma protect digest_block
ZcvEmNyOnuPR4AFgs4kWSn3/ZuU=
//pragma protect end_digest_block
//pragma protect end_protected

`endif //GUARD_SVT_AHB_SYSTEM_CONFIGURATION_SV
