
`ifndef GUARD_SVT_AXI_MASTER_TRANSACTION_SV
`define GUARD_SVT_AXI_MASTER_TRANSACTION_SV

`include "svt_axi_defines.svi"

typedef class svt_axi_port_configuration;

/**
    The master transaction class extends from the AXI transaction base class
    svt_axi_transaction. The master transaction class contains the constraints
    for master specific members in the base transaction class. At the end of
    each transaction, the master VIP component provides object of type
    svt_axi_master_transaction from its analysis ports, in active and passive
    mode.
 */
class svt_axi_master_transaction extends svt_axi_transaction; 

 /** @cond PRIVATE */

/** @endcond */

  `ifdef SVT_AXI_QVN_ENABLE

  /**
   * @groupname qvn_parameters
   * Specifies QOS values that master will use for each token request.
   * Each entry of this array will be used as QOS value for token requests made in chronological order
   * for first token request it will use qvn_qos_value_queue[0], for second request qvn_qos_value_queue[1]
   * and so on. Each QOS value is bounded within [0:\`SVT_AXI_MAX_QVN_QOS_VALUE]
   *
   * NOTE: size of "qvn_qos_value_queue[]" array size is set to "(qvn_num_addr_token_request+1)" so that,
   * at least one QOS value is available when transaction is not configured to request any token and master
   * driver has to make a token request.
   */
  rand int qvn_qos_value_queue[];

  /**
   * @groupname qvn_parameters
   * QVN allows a master to change QOS value it has driven on the bus, while it is waiting for grant
   * from slave after requesting a token to send a transaction to an AXI channel. However, this change
   * has to be in an increasing order i.e. changed value should be higher than previous value.
   *
   * "qvn_num_qos_upgrade" specifies maximum how many QOS value upgrade master will perform while waiting
   * for a token request grant for sufficiently long time. This means, if master requests a token and it 
   * is granted soon then there may not be any QOS upgrade. If it is granted with some delay, then master
   * may perform few QOS upgrade. If token request is not granted for a very long time then master may
   * perform maximum number of QOS upgrade specified by "qvn_num_qos_upgrade". Once these many QOS upgrade
   * is made then onwards it will not change QOS value at all, even if token request is still waiting for
   * grant from its associated slave.
   *
   * SVT_AXI_MAX_QVN_NUM_QOS_UPGRADE can be used to customize usable QOS values. Default: [4'h0 : 4'hF]
   *
   */
  rand int qvn_num_qos_upgrade = 1;

  /**
   * @groupname qvn_parameters
   * Specifies QOS values that master will use to upgrade any value it has driven on QOS signal for
   * first token request. To clarify, when master sends first token request for current transaction,
   * it will drive QOS signal with qvn_qos_value_queue[0] value. If number of QOS upgrade specified in 
   * "qvn_num_qos_upgrade" is greater than 0 then it checks how long it has waited for token request grant.
   * If it waited for at least corresponding qos_upgrade_delay then master will upgrade its QOS value, 
   * already driven on the bus, to the first entry of qvn_qos_upgrade_value_queue[0]. 
   * If it so happens that master is still waiting for token request grant and it reaches next QOS upgrade
   * delay specified, then at that time it will use next entry i.e. qvn_qos_upgrade_value_queue[1] to upgrade
   * QOS again and this process will repeat until token request is granted by slave or number of QOS upgrade
   * is reached to qvn_num_qos_upgrade value, whichever is earlier.
   *
   * NOTE: Master doesn't support upgrading QOS for tokens requested in advance i.e. it upgrades QOS only
   * for first token request made for each transaction it sends to read or write address channel.
   * Each QOS value is bounded within [0:SVT_AXI_MAX_QVN_QOS_VALUE]
   *
   */
  rand int qvn_qos_upgrade_value_queue[];

  /**
   * @groupname qvn_parameters
   * Specifies how long a master should wait after sending a token request, before it can upgrade QOS value.
   * Example: When master sends token request, it will drive QOS signals with qvn_qos_value_queue[0] value.
   * If number of QOS upgrade specified in "qvn_num_qos_upgrade" is greater than 0 and it already waited for
   * number of clock cycles (i/f clock) specified in "qvn_qos_upgrade_delay_queue[0]" then in next clock cycle
   * master will upgrade QOS value taken from "qvn_qos_upgrade_value_queue[0]".
   * Similarly, if master is still waiting for token request to be granted by slave then it will use next
   * entry in "qvn_qos_upgrade_delay_queue[]" to decide when to perform next QOS upgrade and it will repeat 
   * the process until it has upgraded QOS for maximum number of times as specified in "qvn_num_qos_upgrade"
   * or token request is granted by slave, whichever is earlier.
   *
   * NOTE: size of "qvn_qos_upgrade_delay_queue[]" array should be equal to "qvn_num_qos_upgrade". 
   *       each "qvn_qos_upgrade_delay_queue[]" array entry value should be a non-zero positive number
   * SVT_AXI_MAX_QVN_QOS_UPGRADE_DELAY_RANGE allows these delay values to be easily customized.
   * Default: maximum allowed delay range is set as [2:32] clock cycles
   */
  rand int qvn_qos_upgrade_delay_queue[];

  /**
   * @groupname qvn_parameters
   * Specifies how many address channel tokens driver will request while sending this current transaction
   * to appropriate read or write axi channel. Even though QVN protocol requires one token to be requested
   * to send one transaction on address channel, Master can however create a transaction (xact) with more
   * tokens to be requested, in order to pipeline token request and reduce overhead of token grant delay.
   * Master can also set this parameter to be Zero ("0") indicating that it already has enough token and
   * no need to request more.
   *
   * NOTE: Even though driver requests as many tokens as specified by this parameter, it will use only 1
   *       address token as transaction dependency i.e. if no token is available then it starts sending
   *       current transaction as soon as 1 token is granted while requesting rest of the specified tokens
   *       in parallel. 
   *
   * Maximum allowed value can be customized through SVT_AXI_MAX_QVN_NUM_ADDR_TOKEN_REQUEST define.
   * Default value is set to 16
   *
   */
  rand int qvn_num_addr_token_request = 1;

  /**
   * @groupname qvn_parameters
   * Specifies how many data channel tokens driver will request while sending write data of current transaction.
   * QVN protocol requires one token to be requested to send one beat of data on write data channel, so Master 
   * should set its value at least equal to burst_length. However more tokens can also be requested, in order to
   * pipeline token request and reduce overhead of token grant delay for furture transactions.
   * Master can also set this parameter to be Zero ("0") indicating that it already has enough token and
   * no need to request more.
   *
   * NOTE: Even though driver requests as many tokens as specified by this parameter, it will use only 1
   *       data token for payload dependency i.e. if no token is available then it starts transferring
   *       one data-beat as soon as 1 token is granted while requesting rest of the specified tokens in parallel. 
   *
   * Maximum allowed value can be customized through SVT_AXI_MAX_QVN_NUM_DATA_TOKEN_REQUEST define.
   * Default value is set to 544
   *
   */
  rand int qvn_num_data_token_request = 1;

  `endif


  `ifdef SVT_VMM_TECHNOLOGY
    `vmm_typename(svt_axi_master_transaction)
  `endif

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Random Index that chooses which particular start and end address entry from nonshareable address arrays
    * defined in port configuration must be used for randomizing "addr" - transaction address.
    */
  local rand int unsigned nonshareable_addr_range_index ;
  /** Random Index that chooses which particular start and end address entry from innershareable address arrays
    * defined in port configuration must be used for randomizing "addr" - transaction address.
    */
  local rand int unsigned innershareable_addr_range_index ;
  /** Random Index that chooses which particular start and end address entry from outershareable address arrays
    * defined in port configuration must be used for randomizing "addr" - transaction address.
    */
  local rand int unsigned outershareable_addr_range_index ;

  /** Indicates which domain-address-range has been used to randomize or assign address for this transaction.
    * [0] => '1' represents address belongs to INNERSHAREABLE domain
    * [1] => '1' represents address belongs to OUTERSHAREABLE domain
    * [2] => '1' represents address belongs to NONSHAREABLE domain
    */
  local bit [2:0] addr_based_domain_mode = 0;

  `ifdef SVT_VMM_TECHNOLOGY
    local static vmm_log shared_log = new("svt_axi_master_transaction", "class" );
  `endif

  // ****************************************************************************
  // Constraints
  // ****************************************************************************

  // **************************************************************************
  //       Valid Ranges Constraints
  // **************************************************************************

  /*
    Mainly covers the valid ranges with signals are not enabled for AXI4. Covers
    the state of options signals during AXI4 Lite
  */
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
La0ehAlXXPTICAU/lRTh8ah4NA2rsyppTSLJ9yrXo8eRTky8dAhcS/2n0zZ5dMiL
HmmkLHE3HdZLq6hw4ZDRcYx2X5GOVJfteNtGUQonqJ5n7fGfFMYeRaZNiPYazwcI
NFMXvFim/uz0Uxxg3n926cIfgPTrZ84UksN6m7nmdUR0mRmR+Y4Ghg==
//pragma protect end_key_block
//pragma protect digest_block
5uMRBvPHbz9jgjkZO5EZnfkkZN8=
//pragma protect end_digest_block
//pragma protect data_block
X8o/5weErdgGVUIaUcIexbhJsIoSSyFNPoHs6yFo7Z4TdN7gvUFic3tvQ/2mNFYP
kO/U3S37GzPSTG3QEmAR6IW/yG9vkUrG0KWAHZLEmvCsOgXSMcOCwDhg76oWK2CQ
xRPBm0psoSocl2a/pF0TlWS/WGl5VRhBn6di0n50syJOPHUmxgMvMPrp/En2+thg
h05JXTMZlt0ci4aPsngsTCh+LZjS1MMaKoJH4FPGTUOJpUAf0MkoSHspNxeUkIBR
J79WFncqvGM51Roj4iKv0hWsMQWES4YasVwpnBcKsf1E1LljomHRhRK/2Hnbow+Y
iJKQlzi8hg2uo/TZYDmQxXB9cgrM7jZG/Jo7v0NIjgAbTIHDYizDLUcVDQU1c/Ug
fHSRASWcKpnBM9127tXT8oRptM9d/Cxcd9Mg7dtGEo/BmCUg5DVpmqXFAp7Teuic
DBsWYGSmnkm720wkbDm2VdHD8fkSNlQkGS1QZ0jkWGfcs8wK1zzGP2gYVFUOQSzz
u1s8RzhG7dbBE7sVevmo47ilukT8pXFFWLbGIufJCkQCMT25tO5u3bd1IXdCMoj3
g8vHRE60GiK2UeqXCsQIZjbdbOd3z5qOBcRnjqyu5KgPf3erMaj6AGLACDUd/Ez6
l8w9d4ax5GLwUspUQ+8rvA==
//pragma protect end_data_block
//pragma protect digest_block
u8Y3orBJZT7s9nnyHFgnjpoF2vw=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
hxAdskQboCEWphyR2wQ7ryxz4v+GdDzHGsUpEclaVcOrX86tx9MAV0jrODbMBHUK
BhLUk5xRNebgpPgRVLPjnMCmWFeDCJu7WEK8jTHNzjY1FdqrZEzRRRpL409zHleH
tKjhcE+S3tXqUy6E5OcrSxAtAS8D6qVb+5uiBj09bvPfUDpZ83ckrA==
//pragma protect end_key_block
//pragma protect digest_block
1TSZpykrNSjK32GL8IYsKCbFZBQ=
//pragma protect end_digest_block
//pragma protect data_block
Ej0wtCGYI85KbMRtUs3OvFuCaEH8yK+w+Fl3O6hHVMwmBJCACZN89hxD71OOWss6
6aiQS6LfHC35iA5QDOWi0MbX5CaB28x0IQmWoTx3UNXiL/ZOwyc1yXQgR8jrgSbs
70gcoecYDoRltNLqFcw6HQDjnDbPyDSV+UI+cYVPr/nwx/tvzFYsqDis5A+qjvuR
R5XGN2L90K0NunHSoWXT1tMSn9kA7Tnf7CBwSo29l4DdpkEJ7tl4JZYJLJhJYWeb
aSy6LYmijmv/eXcymianOXFkTgWc90K4zcNgUS14p4NwE0KbMj4auGHhM5sH+ZLq
V+csbtjR6nvD40qrlINhe0yuhMHmTnaextsyIarIySKv1l2AbVglYgWGX7KfG++6
0zmU6g0zSTSXOTzEnt/nqFgj8tS7Y4ZJqHvKtTMnGiG0AdzYJSG1kQdGIztO+PXa
h2D2AsqF0tEnMXqavRIIVN0HcG6rDxQJPP79kkrZT6+8LL5231gmNyxg84z3i379
9TCygLfvMvaf9lDNbGQZ0kdLuwrN0KkYzHE5AZxKGFSfyiBOoNO7ImlwEXhUPZId
ta6wvdM3klJZ1t0r2pHWPN60nSYEkqLmnz9+50yoMi/xY2LXrgMZYeBC1+2Ha94F
9c2otmME09NUAt0kp8ec4AmlsxU51m78mCD9bRRYrfPdv5IdApv8D5WgLNl54J0p
vb1lfObF9j9pkT8i1yzFF3L9kq9dHbmVhAA84UCLeXG22kmkq17kpZvxF9xcTQvk
787+ZNjNA02E7UHrchRNQMT2gUXOxlPUmT4hhPnMCYF9XI8FfTIYz5csF0FPpqEM
rBuiCG2vGRxWc6HAqL6OHJ6L8KUwur4ggr2etvrzPdNjIOgW2TegGB3jGx58x/MO
RPNElvrP1TyXaxQsmeYgE5e+3iVR4VsDPBD3IXRiIDllAbn2s9SNvcnPqcrqMpGr
6fwoHpFc94GYJaGOiDhVlVzlH1qzxQaqkZ6P8IqbAPm6AmxmneU/hJHEgP9Q175E
2EfjYnAsixauHHlB8jd/VI4OR8C5p9sjDhuZRLQHF3zysR9wGCqhEYrZ8XYNb219
ASQONzng2hJTpF2tHzb7WpCjgNU4ze8E/jcLenjiOS9bY15CiO7HVIwN28WYGbQY
9GET8xEloNGMhETKVK+qM+b5Oo7k9LN3o1TzmUPPKhyQeIRv+Ohqe1zBJGLFucav
ODNJqgOyN0Zgiqhl7gGfI6N9aAWLZxeTW1JOfo4aMF0w2gLFI1oM6rIE3Q5iFUuB
a/Q5N9buYwwaFARJNuA4dksj5XoFlrnmcjD+6DfDhGIcK0OBCpfplulsyXiIOLBe
bLLiuJggYGskuLzaj10vVoPZ16l5BDK1hgTW2OckpIQ+1KKGrhMEUa/j9X83q3J2
WQMB6HEigSYzuX9+h/FC+uRjtlmY1hJMoU00kojU+kCuLC1TRA56pothYo5qXXRG
P34OY/sU9DY7Lxw+lck5pmfxEn+c6zCKMcNnOapyz7UmvMUFxeDgk2sLfwLvPLBZ
pq9OfHnJ0NQOHQrwWOHDNVnOD8SjsFW+F9crDt6MfoZ+mdp/Msze29Coj9DFhwYG
1eaP56E4vCcXmldNo0SLYFy/Y/QwNw46c5PG0Q7qrUnGk2A/lBuptl5XdIRxIyF2
y6CrOoZef/Y9hK8TGo7vSbqZEJfURkhqBhxZnNvBQ9VP0+bYj2UiU1ZDkaamDktc
waafmyFtZ31DgSe8eebQ5uEZvwDh1zdXqn/5u+ryVxEkBwl5s1eyLd62KzLpL5+v
/lyRHoO2mqiu/VEfZBFtr3CoLURegpWPlfmOhzyPpfWhtEStcHKRehKNqS+9RpvX
pxNOLSucgzUCB3sEWj9pjSAe4pml1ZQkHRtjUjgBKrtxaA63hJC6ZSHDX/aGsq+m
wu6RD7YOaLsd4H9DqrjYH+NoFHnw0zkYNwMDqUv3a+/5pFmWjdRUrDZ2NMhzcXUZ
CW9iNXVvSkEwdmMlAVFnPuWIw5iJbSdI3lTk6y0IeAwiKNvEJfgrI9H3RE0gZmUh
P3UmSgvp4Yx3ZyUPt03iBez+MDtEGo1npzvFv8fTI0O9I+i4BQM+t8WmsRtgqWMu
yjBSqY+nQvvgKmucLSs089Lj0D5P82FEksBwAztNvJ4+dEoBPXosz/H+3hXX0yQq
bsRp4vH/s3rwxCgnxlJSBDRkryDPvto03hdgfB5A51GheH7qNd/kBIhomd0bkP55
cIzwYfRYvZTgmRVpbMwRh7F1R40X1R0KDwP8+I8WoyEeIdsBGCxxISzJ9X0zBwWw
xaNK2RlNRyDr1IoiVnJbtq7dB82gyU3AGTqJOoMTEQPN8+1z/EXJJ4XkuwwViVdx
4rSU+iT5d8TGBxT5K+U6ndg4GAtAtgJEHV3BS6SZr8ZNEzMC9w5sxtG+Oe2CxWFm
eqUBEmJIyRvNW/Zn6yldeUcZ3QSfK5eXYFmZtj906iGrQEn4LyQmuHSnGJkIuPAZ
4BSlN+pAgZbDrIvAL79xrEEmnj2QjYxh6W8yQ32K/O5WWx8sm2EUWwbzHDHBzjuv
VXvrLBrF6NBZQuVG8HyFF5Z+ZhqQQoxitr0AjRTI+Q2JRQtRPjCDOps1YIe5z8Z9
AQcHbF+gYgfoiMMJcRQ1F9UG+40tcnP9gctf3qOcv+Fubaylq4k8/TdeJLmd9yRL
QlUoMukWqNhHBJSbqtMefxABB2/lYh2fBbZDXK4jGiTZh4c4WBLDQcFsKq2/+pwm
HjYU6s1e3za42xC6a8KtdWt73vQJN7q8Xv2LPo8iiD+HFOlrdz/lrX1NT9ei2A0B
zrJpqDIM4voOcxizOTTjktHwsG36F+Djgh0OOTcYaE1ZfETAaGn0u+OCNY65HLnb
lxa4shHGvvhF3AVIzGIP+gisgmV0SD7lHojhwgh5jdB5MUsBkKqqVKMbsqPyd828
QDL8BCNIu511iOB1JQB06vaPb61hNewcTZx9xwwXqM8YZCZVL3mSgJp4WCWSRbP/
X3ZbP4BGMirlYoo+Qt+UWMso+i0ev+QoA8AEH5QQpjXGtEYsaSSrHr1uyt1v1/nv
qH1oQ5034adAO4/BKfIK/NrW6wyAY/HKZ0FLi4gBct7813eUjFig1O+LrzRfS5sJ
ikLAZ84gTlyVw7MZNnCQZNOWZYQP4hmfgOm21ZXVsd7mTl9t+QKiwQyY5hEinhJ2
hHfBwOgnrF2SaQiWcC+JrVItgPy0R2Iorn8e+Do9sPUuQjmKabXy+lxgNv77aTUB
fENy0OQxOm22Bh1n0TYEUNuFXHOCHEVXbvqZaBJubmB/JC9jqJO4RrW1QT76wnWW
jJlByAt41ho48I8asPkVZs1fRoj9Aey/6rLO3tQwKk/2pse3Xmi+MWT6jdErpQGU
gKyfqEMJpkHtzn5CM8AR1fVMJN4fURZ/cJIGGtsk0Q2OowBgyrUg1pU3DZw30odT
MCwsH8cIR9vrxI5pbuc/8yfJ1HOeMr7KL0ReEBkcLDyicZLWDdIAjO3tUHjfiv69
5YRRPB/61CYQ9qxacUAM1Jh6H6aD88DHnYMUKxn12YsID8V8vuRqcDuuFAS6FY+B
GmtXjz4I+vadXsKppmCf9e27tpoL9u/WU2COfPywoISr+Dwx0KJrwglESrHP4Pyt
Zev8wZVBpd5tt1YgBIQ2CjVhoiBKHcfE/bFqbXeYqe5ses8d37iZthaoxPMmEm3K
wfgK7M4pqTiN1io2XH6hXDx7lC2YJc1UK+/4roQ69yDwTW/njPsr1DBzAFIzyfVA
8njn3+LZK3lNsbotjVCgDQ8gxEyvIWhGlduX2P2DcrRF8npGaa3QRiW/zAwsP/dI
IRgrMdvEmI/8euf9uyZUxtxwRLoR8Zh1Ma04Y190snXoXdUdIWhZ9D0jilrYF/Ej
jZFxDgX9PLq3BsTh+Q3QLtFkhBDcyL8A9sdkjLTFOrh69FXM6gSEVRgaCF/9+W+Z
vjlutUXemXm/l1oLeyc//FjACqHunuWagqvDUa188U4o+WIDbO5+X7OWNcXtfbpF
5BEusDaTAt4ReMiuS/FwVVFPvNofLj55VM+C8IrX3ckwQ4r6uy+zceyy5teoK2HX
yRNPW6LyVwsed1yM1CwOTFylHuDkbHByD4nWG+eRe6D40TS28rSUefSHo6KRuGh3
SuR3q70x+n1hIMpS7H61c16qJ2I/1JiQGtoExmmNsPeA6rmbp/qnOhxo4vQvB4mU
vc+q31ITJjqPCM6G4FyP75H0uG4/uMMdg67kBcfkzYDueaQUoAu/WcY4Cq1+r6A+
F7jvi1VAxi7HDxP2YSkD7WLyVQpTOWxtWegT69J7lrGp3NNuRwJRvSeUNS5zTwpF
AXQNHTcsM+E8DE/Ev9BQF0D01SVACUSWhRF6Y3gWFGQkI3zCoBFmvFENrDkUoL4z
o8orx2wR8bcnjq+RBI4kPoyEix99HwHYRqKIAK2ZT5ztUOZDpmxiKlDNa75KDD/i
Ve6TEPnLUMAKl5nt2af1o0UCPyJrD9QPei8gQycYL+xjlrr5/gywhsfRE2TiYVzg
GJlMumgJUgNIim3c9E08CBKtRcL0QYwa9HJAuBHLKzyoYCGr6lZ90DeHFv0FUa0s
EuVEVfBb2/4LawWLe2+AjEl8DHBUEvivm30DRwABdgTKXo50JuqBXN24nZSkgMOR
MmPVNJkGYa/OuMaXCHmltO/G5OL0VTPiQFY5//hOmCvAm7X3pTrMsNOftF97JW6A
FyFLiqGwGDutA/hKR/xxX8VyBShm3W4niWGwkCs1g0KSXTov0PmjwOkflo/3rCNV
D08nhyb6yUUceckux1bOEkCNl7881ymivV3Rd1TTsmVfSiiolTkPTOvacBCfRbYI
WNfytMp73oJgb83nkEt0HwOdJBCtQatK0x/YEduvaFkQYvShxcVfJYxGnQddV/D1
UxRLGZ7aS79E1TgXxJcUWokcIkAaCws6yLAgaxIWtBDHZ9r1yVsFzdz/XA91CPF7
YSz0B78LiAc6wPTvD4OSXxoIkXoib8y+9hBVUdOFzNv4DiBQdKeV1fI9A+bd119a
6bFPKzH+cyQw8IAApbry2sMnCxG93zP72tQzmQIBoeHEXAJNoifs2lNvlluXcmdK
5jOQ19czBUxO8PBIN13bhsxCyF8pGBw9tWjGwqzSyyBilW7g1Gt/jiOJLeAayU0M
LDbu8uQbCEEmnY2wGeJnUSG0iH3onkc2/NkSmdXGJH8ZDLyIKoCoJW8mh/ro0u4d
IgFRjglLvu225DwRapN2x/ek8fM+dslkp0B1M0sszuMDAo9iEUdY1yMVMjVHWP50
1q16n7FQiK061SiBcihnFLACaSuXNq8wbrP15pE2Nd8npwa50IrzdvpWXk0TiiWZ
L7Q3RZv3uTfoYS6wv18R+Q39uJVjDucW8GMpkQM6V4X/jYAS1iuA7IwU6hKfgX3i
ued3Rt1T0fOwgRcuJr6PGdjvtc7zruOitXh5yhmOh4OzJRO8YuFxHP9Ifb7mmi+k
nXHFSS42Cg3gJzE1iXdX5JAA4p16WpMgG7r6dwbp/5UgF2mqYnhbZI2eciq+7Mg+
vg3+9EUjZ1LYO58kHyxAevI551evGxPR9B47hWk6BRRl5QgTBpBtRo+NnTGrBfSq
VWiyM9yZx487uRY9ggaDCSopp/M06xrH2kF5x/9KQ/ne2MCi2FiTzGQ43a+Iorte
Dea980QenxMULZFVLA0FrTE1QbWU2QJPM0wqxfBxGQVfJwqq+5+2+UU4C2m7KyWw
f1gCKpCRemn4lgbTZLbFkEkaUXf+R6PsKgljc+oCGl6y3LabRxZ3WUKK0/OmxfoE
RK9Ungpd/HqJMg3/zl+PDfdHlw0W7+rMjWHbMIvDSZ+DsY04GHcR/wIfESxTcF5y
7BDw2oMlO5AnycqbuNLBQk43uSVUcStaMrWt9/VATuTZtx1gonhzGQkg1L/L1NLJ
RtpcNTawPfFJed6XNDVnO74+wUdB6GgW2JRoYtdy67A8Ghcf3Jrs8x7yyhh4M0bF
bfxV8PXf2QmBV5uZaMveRj7KPX/Vi+z23KfyBAxtYMA0nT5TOwJv/8eVB8Lh4Ugj
Xji0LILXc0yP0oM1/Lp1glk2EVuXbK0r3RldQJVoJqr2Bo5qpxvcoa0PW+3A4MSp
YLsBKchogRW8E4j5SsrtGayLL7YLDmlXfqPVn7fcCj4nigQEmThqIKzebJZ8tFcO
8ZAo1sMQGc3G6bGbu+te7z6/Yb5IhOQe2RYNZ9bFUzcmBS9HL1vIkpcH/RQzBw/V
qcCYbq633dd2onpFCLM2if0nWzgrn391B4WXgMVoJXCyhhgMFovQaBhYECjbbcrc
MQ5IYWDSXIVb6xx/9LKdr7dxQUWeSM8TwP+bGh9DCYR4Iy43WiPpUx7E66zGl6Bn
ahZdqQHKtLGrVi1lOfaG5wWDEndrmGavNtJgMOJrhNOL3Cfo62PBKR8AFELvbjIh
/jKL9eKEuNt0rHEhTUJT0KFWoC66iiM5kewisHJrvJH3Z7xNG4CtYt9MpQnll+UB
4rrRvPoBNGQLaZkymj1HOZ84EPxBkcKEnGCt2liUxNiIvA1HbVBqxrLezjaP9/BD
WzZ/Thr3+5YXKtm1BNw9ZOnFDPcr85pkdxF95ZFR8YEU5QfvS+QY3JR73XHRoh5U
uuMOgMl8AOuB7ix1v6WUO1GMMpw3Bmb7PafrWRxESr8++DArjp3OMyEQwwEx0tPM
Qd3yrBJQWiJnU2ZtMA6LeDj0yYocICo5u5GTyD6L2Fbzb9xi7MPrzGXuPW/PjQMI
WxxJHHLIYV8DSOI71LCk3nZ1JUWCqQZAP7c0BRRYkF3CRfX2+rmODyNAHQZNWNzx
ouc7FGa6ZNWwA1FphyvAP+wa0YWgvlCgQ9JlDv1P+YXH6ZhavTHN3pYeZwONuGm7
9Xpx1XLJN4llfA1YJNzuTA4bKDXbWtwuCduxbwJeRxPoM0E78pN/Bma4hK1q4gKW
4P644AD6ZVj1lN/42iMSsWWAwHyriLTg/Dg1a799yCFWcn5TKLTYfkWVIirbbeDS
K/hVgvqF8f6BIHfh8/iEwtaqrftG56RlgGuxwTjan2KA7b3+mSRL8qyNG7ixH4cc
iwJOJEr9DXsWOZE2aWG4/6xRH2/tnCI35C+1QXZEf4a86CODb6K3nymXVr1X0OBZ
jjNowKKNhE+7++/PGkc9gIRO63eug3qsehI/rptc+umyHRI74nAoRQGqinFS8TtV
mp2Kpr0FEUtfJzQUZ2FJgM/s5WssJG7sPfVBMhc5UnFaEr89kMbRrYaFjjjqfrEF
7eh1HAa0BeT3cXQt4W+nIjRWlYn6VAgXmTJiEHI1Mxsx5cah8rAM1miHqcKIzLOK
mbz5H4KaEc4ZVDY7HNu0kYilg65aUjHqLVkiawY+2snNfvEOzsLHa8GKo6xWzeVE
sKE9bAgSKtRYxqNw42eMHU93j/IO9aaUQrV/1GKv56qHJUEVIMZDg/IWChrkQRx3
NvqCVuFYfB+20hDlk9+Zk/p7doArrrB/ODflRKm016oRBQ4M95BL2L4zb6OSHpcU
OJ4f1q6n0dso7mq8UslmwSGbhU/IQqYumo5OHh86s6VHnAp7oXbSl2zsM6thobp6
UThE5wSgNrs/p/mRZbCSnUZUfhNDLUJ18xsVpV+N+eLDHa46ui7EjSIZ5c1ZGa6C
AB+0hoJZxU1Bqv9jKEhbi6vAp8qqQPjdmi1Zm65Q3mLzjtRFUhtplodaCosJdyX6
ZXvR07LrLDUpI0mcUPpOwfPBxWaUiS/kA/eW0hC/FoJ9+iJS4vDG5S+2sKKqhsbl
czv/ficywol5MjMEDdRyRIz79ZNhN3SB3lahWd9XMerYRuKWma0yMO63keXPyEkw
pEdmgRtSMxxcN87mlhcKpMg3jU3QQhuAsVR2oMyFvPFYn0EVdwOrhWWKj0W7oSEw
NtjoKwLvYhtvwLuM3MUBW8Tfct73ti1TSL9UqaeZhL6HcMhPit28ruHheUlNzygD
blQ00ZE4hdw1UYjRB00istiAFItLPQbX/enfXKQT1C0E0hMfYYSqJpVRs0PT5/6G
kaYqHOF/ns5YR7GCFBTUJ4I5EngdVbJj6Yf2P1g42uNcYoA3iZu4TZQptEqFqxF7
M2Xg1cPN/nGpwKfmHyWCyUwyQiGKSMA0aSf5Js1R4TQ0BowMtr53MiicWUCUcqI9
BVuo6bijDL71lQ9suCxh27dnxhAjWXJPp8xM5ThUxIUnAIcQSDuqkhzoCwwGynTy
TdzzIOsoe6FPY9mO85dF0YoGYTNr6TBwCnJO4PGSFrzpcGxd/SzYvKR7C263wTWi
6ys8WeJKBZcWBlG8+uuhRhZn35P9Nvd/20RTdoZjBrgK4RqmV23XMREigQwutKme
UsJkO+XxxgGBZDfLxL9PHn1fbZI3AgV04o6l1zoKmwVecYmx/LfkxAy548RkEp9+
rDrGgQCnxU1XU3tRsCd1l0Xo/di6b6ICWD3M+VcN7SFLltO74NkPPIuM93aQsix7
LLBUZ2jOfj2zql/kY1iophS0N3qqpZn87P9+8DEjrdLsLvB/bIqFi0JLi5h92e0j
g9bXUIh6rIwnRZiJks8wtxA2t7x2VIGSI820MKbVTFw+jxeu0xgoFaeAWaWJ+wgO
lLm2VciiFlDj0biU3oCa9iuy87EeX6MFJHu/2CwhPx17HmuIhrnYe/nQjGE0bLQS
dTDdQae4qwNk9wbU7FMxtqJ+p6bLCBlNUT5XljRH0O0by4LJ0TnSjrp06GfGyfiv
z0pOU/MNP1erDB+ScAU9+A7PGuIIcO4tW7KJNawuEGb/ySgBwmvTUSS/NByv4ZFO
mTBHfWYyNCITAKaAFGF/tZMdJYusI3H8MIPTwvd+HaesrshC5NMPgSeqnASCFOfJ
xeM1RC/C7ah544SCOSpy4wCGJ9dkO+GhB04gPpRVsebCtQoUrfEE9Vhffk7IJOwu
HCOPsnGXbQ50+Mj6/2T9ak/x/OQhjT2+6wteonJfEyQI2hF9RnrTKosaw1w9JVU+
f9B0BArIOv6VO330ohOn+Yq1QxDCAOhQwkueM5pgnsAIQ3ChA1NonbDfcKeuNYgK
mclvBeiOxvwk2IR6B8Y399MtR1bMSl6ICziUKYeNteaO76VdAZHhH1qHDMOXgyg/
ZwV3qO0FYUHdwYiIvftLaAmJ1dj++TWYwSiX/7MHYYw8tKLANczL8ySBmFmXdZdK
OjgI7h/D0iUPi9GPfiajHTscTyTG7H5VMn1JE6p9v+u79TRCquJtlnFDGBRctjKF
Tv3ZVLFifTw1SfUFOSNGGzoKeEkCY530RF58HOE+3sl+QjNvXG6dFKuQtlJe4VUT
uHMaOqlYxFcmG/2sK8cXlxcnE9c99EAsCthZ6I+Ac8DFyCEtBaSpEVINBeOnDL/X
uBe8o4y2ru+7ZzstVMaS3dYl/cfdDU/m8dmUJQIGuXb1NVT5CvxtxBOIx/ASGNoo
h3RK2RUz8ZncULWaBVOZer4SMHC7RRqM774Pd2tnWX8k5aAqlPzehcHlHeVoGpSJ
LmZymV9gancWrlaUxJVUjy/W80ArrHwuf7CTInaFolIGlIIt3dJdQ8q9/6gWY59F
hzsgbndjnBpmq+eXcB/NVXpAcFHzXwpdEM/MncZqYHC6liQYUUW9f/gU1fS0PYb1
kN9Mb7RkbdStY/7qVGYCztR4GjbF0rnq+iAjkBiyEspHy3tK70JL4kEm+Bmo2R/8
hcQPIMSIgkv37/uULMqUciX8MrT6pueDcFh6I6ZeCtkKKQCgOkNxGKXVhnKt7EMy
wQFkPMa/XgG1dvmiH7aPja1yLMRDf0nLpFS3yRU4M/pU3ckoXmfZ3ALKUM9Rp146
lvIxGhq7mhlbQC29KV1nf8ZbIzPi37TIkbq2pDUDfWoJG48Mk0cTATAteXOtpDlP
Q+1xH164OoXjQxwknMtFEGZqs43Hr1CE4LMK1ey04tgkLH4l49L2N2rSWkTiYRgr
sfQ+q+VyrT+KsWWjgrpOeWnBPp8fIIS3wkc+hXsge/++eeZpZT3RtbT2wIwMYDhl
8vzjVnCE9gK1klOA2xqJXw+/dceQvw+xvP+uts/od56XdnEVbegY7iMf0etoKX5P
FWhQ3u8MVF9ldsCygQMu6jEOEvw9FBCnPdM+YwUZTYb2ZjTsO4XRYt7O0MuOnlRm
qhjJkzqpSNmTGLc3QCTS658U0urSnnG+NG9sMSivJKTLXeBC11MHQ9ZxyST2iaeZ
kqjk9uKh3OGeh9mNKlNyIH7xXpsyWZ9kZ84emOtmx1pij+QjU7fuD3RuZRWm1eii
6lRYaIbgrmKYFuVbFt878+dyX/jXf2Ns2MdfVoC5jK/zOxnZQHrKp0pM0jXeG72r
CyJBT5sMNTnQYZPQhIDWRYknN2lWkA7MurainB3ijqNRoBWiCQn2nwrHugtyEAbC
Y2gk+p4yRSq+STJGMEbOqdUPnW1kVhsgctyCL0Li+aM2xplo04YQTGFgzfsvFKbw
Qs6Lue+e2aXCIAV2eWMFTcszDkFoBfE8eyVR/5Qag1n1oBKxg243ehm6T3oMfIVQ
R9P+37cmrG34FRMlT3scgEhcQ+WZFp6KccoKFhE3kPFGUQVUqkkAGd7re3lxDJTz
31zAyR6UobfD7mljl9K3pcKs20HsTxZ6JPUk3b4+DLTCDTEp94oRKhRm/1sZFwBP
pGsDZ9d91XYYgnzOBxYeEZntwNkgFGqyIreRpzh32kYmutt1jE2Ef0lu+gX7KujU
EDtEoL88zTBfrmQjklp0gBX7DjWB1ZwWqGnSopTbeVfuyjmnp6ZHzWneF53ifHRe
1xSDipi7vjKgOuHzbLSDpzSUVO0ewR3t+x+rNryNQr4FNKg48m5Pdl1TZkCzwulf
rX1lUYW64v3ubWMbWmlxvDOUh+LDlXqBvOId5g9xOud3fx6ccuD7bXv/CArkAujh
fWDN/1nhJhNAj2bUTweRCX2KNEo7LH7fNFNsUIkpNUD8OItjkMhZAsqBM161mVrq
ySql9ZGYIK5bSlE1IwFEIvx+EIcRLKhLA84pAi4JTwMu82wVCw1BGV936A6HCl3V
4em3khJelxCdlI1WuI2hySGP1a+pnAXmycDSCTKu/m+75HHtAcW3B/YaXdDeBRqE
sbLVbsFgfc9+fTNWnj3IBl8d5lhJl362ppWR4povLMOg2AAFV8mwaNboR7PA+1cF
XizIptjR9oXgbQfgrVXMjvtiY5f8qOizV2m7uuXKpe2S0vGeDJJFiYFwv65MCVDD
aqt8BGPKS9LQuua4wpaMNMygXJycEa5a2SJpMY8hbizjHMz10p+KhbcoKOwCsa01
RsnaB1PrqYHGYuKS6LG9/ceGwUK+wA+LMNeVElZaZeln9e286W+yaa27XLFmDWRK
u76tzmXOxRVTT3yZYdFvX6eOAUqq6AFdFlKTdqI165YXZdQd9xaSbo1W5EPO248C
jz7G+QVPOtDQWS5VXRh+ljTUjiMesI3KZZkZHjPSzmPD6dcDay73sDSHpwHlogRg
REt9BZvFxW+pXH7Vt3xc9zqv+wm1vM6kDAtQBI+0Ydvk7nF9F95dQch8qH++Tmmr
L22jhRvg2Qny2I+5TRddAmFfAOJt+uh5yTtDxiyWYwg4cflDyO0R0j3xJxrY2j3c
txGnPpoBRcsqxfZ4cjfCFOJwar+xxQRKGdIFdV4NJWrgXH/s2pBOwN5vSTuKH+Od
73EMEchTadwzjZkvnolIeRp/wRgD1R6AAZg8fVOvc5yPt2Tu2HCsphPgne9VguTz
r4pzav9CCqLhQH6Pf/Dgvl3Pp36P39KQkYkT39R88mf1mTS5FZs1WlT7MOCCv/b+
F9547g1D9ETUiQsqsagVgtYLd3ME2OHNxMQ0PFvPUYo4PlKjB6VphGWxwkNdpEd0
AlwxXRO2VjpEZYjpNQg2Jo9bb9SoLNp3EiTBU+CaOiEnZ4R+LyKpeGnlIzhNj0L3
D0E4u6hOEQZ4Ma6KkjU/R5AmsbWXpq3OvkKw1QcGF7BUezeGESbw44K+b4ykOuNw
FZi+vazWR2Sz71T8TCl0uFQrtcwGWxCAvtCYbUqHivuH7EMExclBcKKidijXo8jm
0fOQvy++V0AJ/mFhW2bEXhiyxVqO/Eik+H5XhoM6pLmDcBnt/2VmGe0eSeBNUEWq
LPjjrqKEu3IOnO62xawzxUkaYqY18L9YmnSkspN+EHEQLT0GNbus0LS3d+f60ExI
5n/zwCGeAsx0k9liUb+YgHFzX+B7H4qC+8uvGWLGkCXGnmqTTChz+WsbVRUSb7YT
qEaufKRcY30jRaS3tDIO4Ubg472owUyMVlG3iU4GuU9NTtBX+bMW49aiayIKo5IA
QrAbMM5DPC3tV4mYnz71f25gjv7weOMatcyvcB0P8XC6I8sQyKBLi6eJuphghGot
ECqp58h7wjjF8IZTXaIL9tLvqRqTrEsB08BA8Zj8LUNjsOpjoJkE6Fk6dPdSXodf
rNQJa/BKHT2EIxLMMbsmLBIKiJkK/TSmplmxipgv2oGSO9gA5vkMc/g6vVgze7wy
3SXOtdUK18/N2QQBb4QqvJ96gSIp+veiGNIVSM0n195K9heCrIjbjydGxMfaWmxx
2bLZNYx2z1utvJPtVU6GdzsQlrwVFPJxmnZzQ4G7kG4L5Fq+lHf1hYz/jpk2kdDl
Sk7XKgcNfCOCeWdsPU5hBaHu815Maee8TtPQ74WmkrYUtwz/XPMv67H2U2bppr7X
h3gD01OPolAJKix+2JOjH2oLH9mOXIPNLb+8Sb71ne809P86+KScJ36q7vqUN1wu
9JinVC0CccYZA56BEScWJL+DzZr+LMNMjk8phC16VM8rY8Ef3sJB0JIKilOYetOB
uMeAvMMm/j0qVbIn8Fe55ThqYDIZgTMZO28b3SDg8QBCqxr+/ItnIdaZl6SgGMEQ
BWLKfei2KHlyGkOHIYR/vFyf2xVjNN8ASsx6gZpIoThYElNx1h9UthhidmaBEYdz
h4FcukjJi1ZjJGSW2qkt2l0DbAhF0omnuUG14ny4MUcAFfkjsOx52Cvqm2/2piq5
4Qmg+AzB9hUPNYlknX2996ynS3J+hTZPfFGQF28fE4DVj/XCn3LYvIrZ5la9AEPx
6QXowuFrVxEHZT0bZcHZuzcynoF5R3qvZNS6mTH/T3GPGRzNrNR80b7y9V9RQy9p
35DxJuDzxajV81n7CLS7HKMWVJdPBTMyol1KsZJQHYKLecnCtiaVGWNtn1vqOroR
h9ZQNdMsaZOvPPGcNGrdchsfbfVhCx9MBmaaX02qic4WUxvG6pI6SlyLmZcSEw4q
KIEo+6DfiTcd/jKXz+MaWp7pbYQQo8IhCJjAgDiguNM0zbTj7o8Ftgk3sCrFfeCH
pZHu0eMEKqr3i39gXup7jyGg0TO2HiwbZu6ZkpTcEy05tsIg4LoemeqLWU+SvKmY
TOMWtmH65WVEtupKF8BzjxO178OfMKsnq7XDl2SEun52aGouNnLZ8+Ri3Jt2x7Za
i54LDrINMbRYL74Q+tEULIwy+Z/q7YxgIBL7TPMOYH3tMAnnQAjMbBAVZhJsLDvJ
p8PG4pfNdiXLZT7jCkG5UsyiRkx5Q5/t1eSq1h4zlm7nk/aClWlud/5BlS8Iak/2
W/2gqMukfKMMRtXzRjQ+5dQKKpMOOF4Hj8qJd15djdrfTrvrI+24acmBpS1IUB98
hKa+g2gY0/R/QzbGFxvLGBh+dSSRDv0XtVIbYfSFUH0Z9ZEY1gjDlC+i132v00L3
CPyMyDEpYoMzrH0YnVai2oQ8gbK+SdO15YmD45gj2d0lclZDsaqk1Owkn8Z+/D0n
1cHPp2KIqeFAFI3Qzs2+th2iogxNlOuI1JAhvCPck1/5g1z3v1hRDwmH/sJTK0jS
5Ka/XZ/d9fwE0iRGSmOj+KsyYqiW9r4UrurJ0vy0N8lhvX8b8e3t6WETmCikWMWI
5UVseU9wuX6Scz3k7nooLJLXujgwYyHjciolUe8BTk+sBBmrfKT28aJMfTBXXiQ6
q34JYDGvKClqf/dCs7RUdZiS6b6D2fc0SslGkGkcDK0ls+FnLPO83vSrSJPcr1cO
J+fG65tM+ARC/ztQxYRP61pSzSklhwSWhg9gr+KKvWj/1dXPk3ZgUD/BNdwYrx/z
0xVbyUeCaaUL2JiM2o28YlWCXWM8hRtLmFvXsmFN2VkksKpZvloTygDIixcKyY94
cD+jOzivOAlqYWiGAGou+hWxoV8dQw82EgyWY5Mfu1F6L1CMjkw+nkgNCzl7XvQ4
ae7bYJooynqfLw531O5soxK26zSYxylqRrThC1Soytq2jU2wt8NEvh0vwhPUKq0Q
23mOLSyH08ZnwF18D26jRmtavi0sZoMjEFdWY47nOsS07bZVp/3DaxwZJuc/BTWR
9AxZ4w1Ou4Yq+wYeg5A7s4/Qy6zN62hA/kspFwJ/JtNRVEjEpK2fXhktUF8Q0/a+
yIDXd9bM1Wu/dwM9Gzhp+IvtoxaIcAEpH2WNRyOswzzoQ8CaulYXAZZn9u9DSXsB
igUmQbvk55hqVuWdMHRvLOzHMjtBdr56GzUmtCtqYQtsv/+AZ7+36HCXPgN0pHdY
BBuC0jy9A3KmMliWYiZQrzbz4gLwCnMj/ShJaLkgWdm+jqdRpebsAD1ZwXUoWnTs
IPd3eUdx7fzsYFCNCz3AnjYqs8LcBIjaAkStVnYgsvX55gRSaVq9WkL0s3cvSa7A
gQGVk6v/xuGKJWJCsbKPwYbTlwkZaHZm6Wzc6uOcfZBm+kelxMYEcsVtSws+WzSV
FjO840+vyzJyyL64t/hn8PDnu04Ci11HaP7jinep/zkENLWgnSc1lf4mnLsb7uhv
5gX2dM7eRvSnbUY7Tggr1C9fdI11NqVaZ20ST2CFD145g85cZ4GpWP3VzHA1Bhho
p+U+kg93GGcDlm0L33RwzgrtNJpLcs+eVP7KbGMMiJEYGE2y0yf6jC29UA1DqNfr
BFzwWTmJ6HnKZNQ1SS0f1oBw95Wm7o507KNNPz7EQ5HHdC86v2LE6LdtioNi60F5
3FdqhQc9Xsu85eBcDTgSzBrMrfM+W/XuNvuIbQwnP8ZhB2xK9BryCT5fZhVPbp63
+N5qeys8IEQtTYO3GHtr0/+rXgq8rrcNn5XRPE9ykn8shLVxWbM74SllQcmz7HLd
cEBqmF1W4Lv/7nvVP39Ib9CXbzzjrZptDqnOEBl8lsnfOfFP6XegPJ5DOukF043N
cS2QCc+8W4ncCHEWSyOOynBkXRS4hK58ZNYDkq0K4KnnjOG85TJjLKRBo9sfFzEL
mgCrQQ0P82Ui+P0qVVGzKlB39NfWNmzCYbtkI4f7MP+mEhmLS5Ai4FvOhXHRown/
OUqFTeIrN7BngoZIKeAohZ/3L1qlElozRk8bpUxO8aaFzDwt2C2JHIGEA4LCVtJ9
PjysqVB/BtQ5Ihl/cGlyfubLthOwQSXKeqnAVhQOXcYXP6aHj/wVAdlKaJX+Ir8j
RVa4zhJIk7QksAv3YS0QHmUgDWKAibQriiAL7yS9UzHW44APz7tPDrYHhsq2T8qw
oyirKnGlgEYZvP7eu8SN4nQKQE3sCIkMSfjmP1v2a7ZVVVxj4dwRhg3JLPCv1SF1
qYxWFIo2RTGjMKaw+nMoggBIXy1/1xdgrxaqEw4nkek9oVRg2Jj/uOy+lEU5XgHW
9+9l9k4puvs5OcguKpn/drunf2mu1NX9XCGYt/2GoBWXGkH1+QPFJ7TfkiEdfrjo
S1H25GC8gBmqvIygRfZK3ZPAFT/69cjeF+sd8qlnCrQAcdPsljHrQawPNIeF2Uk6
ZEkVAbgs2C7nt17S62LFGc1oNnd+uE8vA1v1K9wwoniL/wyRl5WaaTNEQOl53CpJ
UNmHjnDMw/7ygYbEK1r+ow4saSJ3xaFK2K+KEVgkVaP23QjODsXYnHOs0dZwQQQO
F1MYBjDjrN+7WDnitMUlSKMDa0+c5D4IJZgo7TR9QwYp+KWs1UbKfHRgJdgezVZ8
QDs/qmIxrcl1pZbNRWdmfl39vu8Fm+ylsXFqOtdoSFqm4H2XgYVXW/+HSo10hK88
LI3KkdB5WXrwjKkXd9yZDQWSED/NiMLx4WVJm0clltAkixHtGDNDcaK7hL0SSDxj
nafJtZUX7jeNlHx0nByYP4IA2BfQ9ccDBHtvyZADWPEm8nJkJbFQp6TeEtd3uCTC
9p5n4C7rk+yFoBqpixQi/Q9UKWV/LW2sEs5FsMa8Uz/y+UJDZwx9zPX1ni6ybVMG
H3HkEhdIoMwQ3EATyroKDixq3CsRf3pmUEygAIMjA9mlNCfBq7DR+TKyPg4k4yoX
A38RH1ZpE2LiKafmnZWFndi5OSRyDgyjtLR5hlsJiHwP8888qFBN3cPgsCzIN5gx
xfj88vpM/lrGWxbLoTBCN/tMw3zAKx05bSJ/7t2eGm37jN2C6TfBhWg940lKZuqq
SqoiKKSokLrOEBL9jM15Mu9uv9RGB5pfzQkauvW03CH5Sq4eDFQhf926qOgHG+S8
nybeJS38loU6yXIG6YUk6g2yQ45uH3Y0/OgdnZ+wTWFQDOL7FKDGawB/zEkdG7hB
bUosBKpcktSbkaon8tPX3HbANC+HKyo3Ccqze2npedyBguTMHAHv5Xz24ewXAOLW
wfSAW1cyWPvKFp0ARZtvSYgpy/2idwZ7yw6WBnl/F+vhJu9Lg9TXlKrGrC8+ji4R
dVO07g26u8CR6qntG+/+Z3f6Hfp7Eyn2VD24ZYVj9VXd8cd6YZZbQcYP3p5dNynv
Vt57X33IZSLrGB70kn1Lz1UUM7ZIVmIgp638EDlarauYXSUUKF2r1w+I8VhXDgyb
Dy73/ISVtSPDUdYNMwtvcV7tjPU7i7eTJYTwpUUPI9DCVSpuXsiAIyVUbrUkt1gu
1I5F/JzdldNUHsbL7YnjE37cHlOP5MkSWTkuJmKVeVfPf6wpRcnTRgilO78hTiuP
izcqMgH0FeU83Cvt2gBaqtHmZXISb0zYUJcneeekAAPBktQzmJyGwbPeTmf8a2s3
spvaY6x5ExcRBbTgTy8PjPXkCcS+ZKMJkqeQ4kKu4CF/AN9S2Jfx6/24TiUuHGt7
spBlCvriE/GbwwZ75KaMNeWbFXc3q8QrGkr06v+GcqFhpNGKHsQC9uGPLdVhFnFE
jO7Xn6xABNXOlGQ45/dzxW5dLQ7BAv9hSlodvYkNmxHPbXMbss0XQhTZnQNHy2Ze
vpELfDWpvylnToZWMmwKG40ZFhZskWI4Fy40iCQ3VhWXkE12m2921XIpkFEA3KI4
Sc2D34kA8/qSbS8UUHxyo1QLpM5seZDXI8WsQfU7pPzwL7BvUNMph3yP1T9IO5Yy
gXaGG5DooOtCj62iqVHMG6L1pCfEEOxvbCfsJKJRgI2lScRFQXXMJg3K5P4czNhy
XKlqP4xM6Gth+FZd1OKhzscDzJxvevMSOeIBfMWhp3MlKvoqX0el0h5Nk5zIp3H8
eO8b5YzOiKz3HM9gfIRP2nyZbIOvQHMKm8OhgRWARK+zYEBiZyhOh7PFtE/TKsHB
9F+Im5BIfkiVe656vkJu/1ScMBXPsqY8X2taS1xjmK+348xP3u+3mNmL4f0+DPbD
ejny5fnGHRWKN7OtQgx3eo7oNIkspuMAUHNcaX1AXw7KiLvGRg7y5HGqC9BDe/+v
DnuNzdATACBwgCrl28bupju2RT+4paa9DDmJFyEXjwqqBZ3jqV3Fu+zQC/PpMZVR
ml4oaico8pUK+vPU0dEgPb/74Q0VsRXPDQsa9zJhAQGuBf8AqA3jaonXXs5/H56c
hn5LUZmjGhUakmz/bt4C2PE6LDCEONzg3J4DnDrEONQvk95LYQ6CEyijf/f504FF
5gX1SIaZ0DXZSbdBQ/VkwZTN65SQR0dEKqamZw4d2PNVROq3Ou5tyCbxlaNOMZNl
O+8EfYgpzUloYNk+uB7u4NyBzMypuggdhvX6AbCg/juhpRENVyJUf4euXosiMt6H
sePBu7qaXim0frucqr7vuZeF/Ed0kVon8A2XuqpHU/+LydJ6tFqEECeqYoPUUDbc
f/lNoDU03XqapFGHBkC4Kw1MbjnkICRemg3FERQ0KOaGTbP3bgTvIAdtaz9mAuSJ
n/4ddpJySvz+zo5Hj0Sq72ACV8DeL84UhdEAt1R5M61Zr8f6hKICWukq7mUoXOIr
/VNhtzboEm4As7ZXDvEupkDjkvNBuvTtTts8lZZDo5zPc2tIH4u7fBG5rXs5cpbL
JIyp6I7wpEFN7AgMOmUAjsazlMFV/KCXRkr+BpAPtiImWS/Pge7CpSy54GnyJwp9
LighQnyCFaSU8IwdKJbjKmlh223c+N6CBBIpgqVgWE6rrhKHUNvR6rsYfNeeJ6bI
3HDe9jz7aGP2F2R+nxAGZQlmeNaA23HkH5ym7UFCY5SJvMwXA/jyHG1XmCI0MGLC
n3OuY8891ppayTPcLB48fXLstbME9tg2rHMv/4ep7AegZlNp1t2dxR2+Rpj0n0VU
enB05q96214ZA7ZLQ+3GBafLWwpJLYBrD2tVJqb2YLSpa0FuYK+A6+wA23FaXNV0
zuCCboQcII1ZdBT194+J9+39fhSSASF7Que68RwOS//HAnpDWYSSxDRifndnCFtx
0BZk3SPcmBPTcGNlJNi1CI6ETFUjk6kQZuAG0bKEtbz1w6DAVRAO9Io4RiosFBaz
z2hG/LIeKfVwR4WJcv7dYekQxvgJMLdZf6Rdz965xwxLBulmFcd3Ywaz59ndzaVw
X5gmoB7T1mI6yMSNMYENMRD5W+OFfffiY0G3/kxMghwbQhclbm4N0lrPiCQ4r5yB
SDTUm3ER/i1MniKnYWnmgNfzYiM/5zlBCMHRc+xst+Au09uUlVEEY/WPj0+puksf
ANXWLrmh96zMwQETTKd7loniIPakEi86ZRlGj2bAli3Mn96VhoxlUVxMnHsc6nSZ
WpZZ+DpUxJ4NuC8cyVNffLgkE98eG57nWef7KC1N+8nNJsqvx2RUeULam7eNg5aw
uH1eE/y8uIlX6vsVDxnaQh2enfnhhLcRGM6sVewNPLiIxEvtDzIx60xJTC1EyAo5
eTLJHfOAFNOvt2pyaYs4ZCuCusuwqQ5VOGaI2vWVGTn/iL2v5rPAbLV9m73KM35g
IuE5OYWZjlvp+VQ/KiQBorl9SzkPfD29DI1R7sUOO5gbTzouLrHezGkkS3D6o49U
YCUfhXmjlRxAGYXjaW9lQB4y5TeYh3UBFidjLnwiSVGYLotaPoUlnrArwTrsnJD/
m0LDNESUEiNEWP6aEGmYrrhELEneD10c2gYhYtdAsDhh+xA3Vjdieq096WZ/MjTF
/PAX0dkFSFT+AKwsOhaUSRNf34LIf0G185xVxQfcBoM2N9yle/kHnyQombDOBiyI
sWSG98pLFnYxx57G07SIhP4oezPAH/vihTh3OpwBVpfkmd4UynpO4PyAD5D4Swlt
NK+bcrR69fbcq+XwfcQuQqZszxcZJhP/KJQbpW7eg2UK7W1lzk5UJsh5rFsLrUNN
699RBflZx8AOhJ9B+q4tYrw8BzC8dfmSDQ53Rx/S4XXmU2jgu57ApcYepOA+hGo3
DFz8rp06VlQxBSpinna42gNVTV/2nzbv1QXtoJ6HpIxD3A3eX8J3l6FTqdz4vUF/
9J/fb+OpSYVn9V6Dp72TR9hvm0IcYitlJbpNT5MG/+3rbmP4F0LAVEC9oiNTGpvw
yX9gbXck0qUtK3aAIMOrRXPRdaYGrouhG4fI+bXLWYkIyfjhN9VkkgTswmPCSmHm
d4X5FabVTO3dm9ccIFgwxv19rtmIZbaZhoCyNX2dO8VRZnVt9BvkAmYowfzlhFsq
aIcxr+xC7mmp761VjCSdxoaaQA5JTtuhBmgUzNYlwvh/+V2UKL9rSXOsBBg95na7
/F2TcNchHV8dtxDL/h0HBHdsDGLDhQd70tF7WsC7StLcpCD47xEW/ZkDAi53jKKi
QlrShfBlJH3utwy/7JfqBOL0pf9K2x61MCo96gLnLDRyNP6LKMIU0wtDjJTPULJG
P97VXGunkL3wbMSfyFiLLHzm24My40G4y4iypPZz1blGH4bZDDB8y2LhpJTMajxF
T3bmsWuTfUKeXfVnRD4DX0O0vyzhfW2hNTPVBcS/ghk/AxUH3Q/o3ltpGAt9p8aL
ZIGWoxkK88Yq6bXRTFauP9XzYApZNIe5NfFwr9WXi43Q6tGFZt0PzObDx1zsHyJd
X8v7F34fB4AOOEcrIprC/n1TZ79fYlT7jOTo325bGbm7LH+mOjWjdNdaeqemi+y4
nEc8y1YHv5y6SS+Z2FqCn28ZF47jBSV48X0xiL+6NSSXZs6gEsT6TirOFrWjsT4q
CZsBjzAOTFHa9D74VVkGhRsOobCGjD1dJRmBqArf7yoUezNoKVpDGiILn0BD/RtY
VZVp0DrOhM7slRnl0rCxb+poBgq5WP6wR4OpNczfiZXJV0H2cx1JB3YTT20IpCs8
hGx1eZf4sPeMf/HyqxBHq5DRlRzkOwpQO5wqpasvXoAKUwuk/jK4e6/Yu0g/E/mo
3IVaOmSOzmN/8Qeqezg7fBkGmhWFiTDXr00IzA/Oz3xaU90pR+j85Qh0NDVbgJFb
DKkTIkQ/UJWGXxMI79+ECX8KzfO2McwDb7R2O1Goj6qGZprTdWLni90FflXbltqv
pcjRr3VEQbSTV1gmtMA1pLVUoCQ8ePEoTHm/0I/pzAr0waSwJOzTBvRH4T4ND8NN
A8ZiAot6V9RpyWGYjx+Z/dvhS0mQYFayUpwgoLV0EEmdj7//xhvfG++d7swqSWzT
c5ss5oew7AK10RtUduMG4r8gVVxgwL4NsMILw+oKMIpx90JoyxyxLLrxW+ECndxu
LlAta2y29lak4xQA2PZblARtSBpwDzfsPaBRKTXJ+97NWw311ePoWLb5su2wPQ2i
xqqxCylJR14M+Diim6Xeg8HkRkhwTiXb2hsWm/vMcnBNLI+2h+qKLnBszTdSGGFc
MIvmnt1d8jn90JwkCZ2C7O6IKoo1mY7swrsX+NK69lR3cAzdPfMbhtphkYCIHYXE
q+gHYuzikWnMKoiZmyrrdSQu+Y76L7rc85kfnxuGealOPamn2tyJ6CIA1aoZJQ3b
GIt1jsa+AxjwRxN3OnQVh+O3eqEUj/zcbFLSf7ZqkBSSMoRs9QSwk0KiwWCjuKhe
1jdtI4Rbq89Z6f1rmN8TuP2B5M6MgZZ6Abq9n1+NUirnWCRqM43SSd7wWtNMIq+J
96ioXFJYxjhjwtmkHzrtQL9K9Fbak8hoFB9sk7ZtX8zgUmPxmKAQ0eYIOj7iVbQb
dSAflJLjhLorNk4rbF6k/ZRaiaJGNcep1CWjH5ZnTeSC0DdITmEWLCV3vdqAxADh
IDAH9BnKF8QqOU1Bdjo3wIqjz3BXc0MirASBkzOMIsOLBJQte/AGebKrpsyPHuMq
aSvpq5N07/G+Xa2zs5xuiRRxHPdiUsezjERY5BhH2xiNXNajGXwuIzRUdS9C/5k9
lZdaR+MY7QrlcEuihfXccX/z0Hxya3p2oNJ6sXnlbtUbqv2K2wfPKOr6F1/9B22F
jTW1UR5STj3GWB1/8NDJ9VB1AOZ7lNIVr1gd4LR2moOqJAmzesmT535zZMTLp8jU
pYE2Uu//RBgEztL/nAJ12HfEhAfi5I2ZX15N/nKgat3E/+O87TQ7F5zdJ9SSHrMN
k2ND+dIAiI88yyjy6S07+jHzpqsMzJZxPcBF+0S436zbPx089uLHe1vxbIWsUYzM
MGmigwgelExoirea8TdLcuJ0ZR9ZOdE5q8HiNQHQT8WtOQ8IRErjCJ9ZSKILEUvN
XvaXzxFOyyYVB7SUJwZpV7soM/oMwu65L97JsblOAUuAT4qMIKsinI3O0SYmbM+S
OeNbMyFdpu/NCLWacR8Yc7ZRdURjYY7Tl5E4qvbUavnHOItn8ZxrH7CBS1sj4qAm
pSEwmFI/wiKCVMWumPG6mkkfruQ9nm9kkgJ50jK48vMhHJsnXoJXyCahmydteHjG
6m/tv3SuVwM1cScpKiUOqImRdIny2gbCsf23KRE+fMEr1uEJn9b5wi/cUmXj41PZ
1DDRKnd7uVGWEQa4V8m5N6gmbWaJ+1b7pSEXxg6v250LGxX9JbUJxUArHrIev2zM
DSYw5QPEjblX35/ZN+wYngI52+PbUSO7VSkrlbNvpg6qxnva6qobrgacmCPBBrJ/
b1OQoJktUUKg095B68Ax+772JkKegZMmRknLiS5gmY2emPw21nF3qceOHqNwgYqc
tHJ1zF/S17wpO3bA77wPqMTW7Usk5/C/0p8UwQ+cg68pTsRFak3Xzessb6+KNQgN
RiIG6EtajvKGzgBV2607gP+kxhnvn/nM41oEqIWKtkRbxmKcyAeGKTEckcfqQRcJ
50WVfzqsPw9ep1ij10ihRwvkxPIT12pgghR13DXpS1+VrOHmr8Znxxy+GTv5v+kz
rzCvxwapQTbShucfbm91npCyYllkkjEq6ATvZTAW9N+lamQfHnsNgOAGqzc3lIGn
shNKNNe6g7ST5tZJ28xFrQw2QeO8S+Do25R25WByg6jqC3dLKCfabNBg9E2uSWiQ
O0EgaTeTBQW7e0rfdlbzJ576cVVIPX7TfWkawL3sZNNe+JUVYoGyYq6YGD4dk/Zp
D6KVQZPMueuyKi7cJFsjjKvywjOichneQNYF+mg6vukuk1d1rFsOEhm7Mcnbq3lZ
HZo2T3Dkd2QQIjNNbvNYfpalNjQ0FF1gM+Ey7E3crL/peMyAduO3dWmIj5YMdeKo
TVflzFIPdXYgJVdWR8Mcl+nueuLE1VN8lJfVJVEUzF44Mh/jNvEa1hWmDfWE3npD
0oUuaEVzg2QkeBpvLBAS889Qm55CEckeBmRTUr86PVuPaF0d4LotNQo3OIxzAg0l
bBFCDFuQRoA0j+EGjbBlfJXqZJTxwzVEvOVLIjjAxCvowSu47FmXT0r4OyFZmuc3
9uUBSyN2xA7yBQpKN5YsB0MUmOlvExIW+xP7BGZ3GMKyd0Ar1DJKojFsmZKANCxq
YD6ENvSMxLWlunk8Js5fGz/pitsGv8KHygGYGmNDx3FpF1eI1f8BXnkkaFZinDfB
Pi5Ow4wXVWemoHTC1YUZtJ4uCu9/mddyDFKrccgLiuzQEgONn+yqQYrBGltfGsfz
wF08qzkjtcAp5y3JdpMYiX4v4NyJ5+0cm6ih+dULAnhRkaKTy+V5VTXIlcX9Z8Fj
PNgAsN1VufSuhINjYKTG+u4YhVAInzS893MNEdrxi8ESN4XDuHgymuAVgfmlIXec
cQOPeuxgEkml0757xgoBVWY77OUBwxNG3Z53zvXrlOII4NtXyUVPZYwOJaaWTc2A
v/Lz/0CnBAtpULLJFGg4uTI9UmJNcEMI8IVvhjakMCraDu7YhzzG1wjhgbSSjUVt
QjDBJVlNIrjHGcWVr3FeaQ27v9FC+ybJgNqbFT/9RYNjiVZfQIDsAZLe2FLgoO00
q2rozf78qhuURc86wNfmvUwz415HODRRlAqUhQ5CL9tdSYycnSIYzCHocerWeQ7a
N0P8oapz4HGG/0v8HwsRivs693eXJEzb5JZLhiB3dePWBmPb94mbuUy/EoykQllp
gn4q0HCOc+kWUvwcTaXi/zDQ7XOMl2ebVdetW6EDUrzKcsahwoDYVGC5rNFLb3XV
0uyA6COaX7AOY3ZGN4JchNfI5YE1yasjMtA03yTvrVMcQmZSe5xIAe7+6xO1sjRO
gXdXB1CdHUJYvldTFVurWd6Qlc8xRKdcE6mqQBFtw1vIpEntakL+CAQyf+Yh8pP9
Wz5WF3ryCd3ioNMrgUy7JP45/nJ3mdXuFCpaoZKukck7d5+aaudTyK5TLxBH2HaU
+si/fzOmnqQTTH38SEeuEl5AK0dyv9IcE9sf6Ngl/2jeEeNtpgxF1zx5T4w638nn
BMBrgOAzJvYgFLq0nLomOBFhW0EhTiT9hcQx/sRxIcsfqFcM5Pc+7sGyW75ChzhE
4JT/2SwnEMT1t4KownYMYpc/OGKUjlUbfTrLlWqoQ4uOum1rB0DvuJXteW/VosQU
nZK1+Oq7DnkilMOuWfLp5K1/kBCWq5VkYxJzPdxH00gBDF7g51hKrJUVBHsKjrQF
q1nYgL96fAyzGgbaCct9nX/nz4utf6c7YGE/wnSbBy9ZNml9XrnZM5u5UMs9OtOA
KpcUzfAaNoyQuHNq26mA+FmIog9ZN/MRwrJP+Ah3GbH/waAFNlarsy85Vlh92XY+
EOye/46/Q1+dV6FZvLav2E09PbBuZdTa4vNQCBZiE8R1PTKcr+qHfEIE8cDu5Oag
8SPkwV9xzx1KECgM8J5xjmr5pP+hTY8K49uBTidze43/0RI7JAK+q1h8rN2r02gi
gpjOXcZie2vHW6LhIz63wDh2yK6OjteKhoVjzdVQEnnZpY74ejRpGjToX92hPJ/n
UfMPEBZSAOzRjiXdnRThLbjXdJZ6bA3uOBf6CGOJA/aciy6sL+fj3QGx86OG+gD+
hzmgVWWsUWFQnOyAkd74dcd8YlsslTxxLBTR0etDcywn/moMpUzoixkPAeqnMEft
q/kU2IGiqCfqF8edcax//WBqwrDApwcRGI4HkBiiKOwS5GIUSrxMyZQq3TxAzQSZ
2SZpYRmWEzu6hZy9i76Gp6L+NNN6+a8H0WWbPL1H2i1zyKlZJ5vaFkFeSC0XgJAL
MH7SEnhcfyfdh1975ffAmq9ylziLrQvj66sTosI60BNuOgaA/xjLiTjvWbwPqXSe
d2yX5bdVIQgsNExE0PAJIHK6zsIqEfu5hfC5UMK6t2S/JiR77ZQmr+cp+sz1eYay
2F8Kmz8iMJLzUS0dYVTT2PBOoktXygkLUDPmwsw22zEvBTwxsWckbNcu9eTu0tks
7MOoTFVI+Wd1sHxjJrTvQNlzvRhHcK2owkPVjpqb24xxRMsNzwcEa9aNG6cSgmR7
u5aiIYyVH1rVEGhpKnrw7PwUL0ZD61CbH/KXJXNXHMkAt09WJbWmDBUuSARyGvBK
1opQ3ey3cmOzJ5LWNzGdhQZbbguwuTkkKfRK2XC/KprTXnPoDs9ua6JI8VD/X3ct
dWF0lN7bemUvXI4xq8GpXDudfkcl04tZijlOEM1BIi3T4eaNrc2YQ1QAMJvwYi/D
ABQz1sMB0vRQtmW4KINPMDaktmM12Clfg3/0Mi/AhoDyJBcCurrzSv2gR7rV7XRo
1rSqaHfzQibM3TOjZz9CstkC0/Pn7o3JsEaUTJw5Ipmp5l8CULvHJg1rWJHyrd4V
+f8dJydEknV/8TmsqQPDrlXwp/PJHDiQ/T86DpqNr0xBIliDsHE51ZyAH20TgdGw
/deuPstTCayJgkGc2q6o0eReXqcToesQ8AEZPvC84I97uo0JUqcKmSCmmcgO17/Y
KJZsHZjyGeQldFgWU0Klu6C1+wFvoQhYLrnUIZpmE6VOwIlWqC2ER+PiaTeGfapE
74fFqAQlf6arhSefWT8/6w+irJ+xORyzYg/6baNZSCT/lkBmpGy7FC0jP0wUcVZL
yUalEtdv8QyETtBvLPgVqd8flADSvzPrn1Ak2ag4nhnFZdD0ZiUhFM72vGgQSuzc
mnBcAScC4K7VpwVjCpKvv7UE8Ya+rzfn2myguIRHEU7PDf0vwz4KlaHP1ZQygWw+
5aF01V6XA4Nx8vQ/slbnlDE6oHfRItvIsMoHLhdthVsfC5LJ3qTIk7Mlc7tVlELS
KQf9faYu0dnaY6fOfoeBfZIYCrax2VeMIHRqIysrGtiDRX9RfK1S91tAhbWcxEvY
Pwq20x24ZOvS17jOUr40q/5kcon8waS51FHBsJKW2TPZWg3yP3Iz0KGlq3IfV/Go
mb/YVtU3WROdt3uNL83C2wQ+DwX90y8QV2a4WP3FwNhE0l33kxKokMjmuMeHNdIB
rVW7rq+K5fB9XtjVu6OVF6fycasYoOqIz2zoE+0wrXwiGVnRFGkqSvuB6Nz1vU6u
QgcEolQAJhoM9DUE0U5Q30VHpvKF8Ss83WBLOr8qyzOxkSech+ecjsyiZIp5VkR6
hECLb8S63boB5uQSYy+5imfBmRJLkV6u49ygkeoyfBvr4xXk8+jiiDQ9OdgB5pzE
KhjGht9k4cxyOwwYpMy2zFGuKfXH9y92WMQAGNjPPGgTAok5tm23zwUnkW+6nQT8
U0igjhAZqYgsdCGp0QQMa2ubM8IKYxwcAcGsp4Z+XuvfuESGMHRZmPppWPUA+tyy
gxRDJe3+yWXJr8n9yNSwWvC5SgoWeFqY0ZgVrG2pbPPpV34ADrgDPE92aJ6qbKsJ
sS7gV/u5MeRAuGIvHX5A3nupSO4xdVElX/KyYpAp+yvTHxzhjbUgKqvpaZFPa2Xp
q9HDb15f5zh1DD8Um38stHXfg1RSkNZmjOZpA4gXAEC4NWxWhyDTxh2oA9rCXjm7
kEABf8bMBxzrqu/bwrzhna9mAKsk8QXo4/awqDBaPD4/kgwpuu7YDr/xN+/jU43P
FmFqd0XB1973Fr40xv2x35j0lDMime1OIZtsdm608iqsr9oG1/ChqZTYBsV+JOD9
tUoeY/ip7TBkeT3k2nRP7DB4bXPPfRTDXhy663kLuBqZtCp/iMFJrPY4TOzWL1ye
oYe14tkH98hW+z95BN2ZKuO6Y7K+slPQDm/bB6L5rRl1Z38jqdUH6V//m8qsxkGv
JvbU9LM1rJf97sEm/3rBhJ+odK+Ip3X72jdNNP3KazEAWX/WtSAp3WHTuO4VWurH
RyFMZqpI8RqxZ4vLkjJKlEDMDUNkw6UJRvvZhKwm9qaiOvEL+sp0Dz6fXjBetRU2
Y4Bl+7dufiBcsH0o16CDFKvtbbjcK+pdRMLwdoYsx0GzWHzxEuLZelq3tFdFppWZ
uGxXuqTK/EsfYLVrVyhlgtw4qzpPJEAllQOYViz020X1aH90Pm0VO0CEP0XcIaDZ
Z8Rg/OMJoCprZqNoEy/LGKexX+5KYxHqgb6KbikaxcWmq2iT5AD0sBEU1UDtr8WG
ltLJ+YyU2zB8WeOvAqqQDlbehVS7StxJHRttB2vc5asdsKhnDxSWyftWD+31hcMl
49I2r7GLAMJAp0X3JfIisi1uOYGr7G2ZT7WHAsAjlgqcVdaOp3h78rw9HhwXNPn6
lhb2NPYN2NVETLXX1ITXCv0uDi6SW5SVnEFe0b+Jvb2rp7fBQ2itrSrtwjfB0J0F
/OVYVUk0BaeL2FbnPhFVQSlw3WAocXb8v74CTzhbRNsyUCJQR1Qywg0RQT97zQzs
UHRCHfmgM7GEI7OQFDzxx+CkvXvt/zBfRfsfDUEthw+QaRuYTq8dgFCBCq8V5ifq
HXp2F3OrveW+0M7pBv1TUyK61VEiR/tJLqKVgkI8S/GO80xdI/xzBejAHZbsHfgr
VisDp4kn3bwRPuAk/7EbnQ1+bZylniMECXTp13tTvgavcNeoRD9l3eeJA7hW2BT6
8D/bJTTbQB4YJoH5WZRIvIbeFH8qkhFVxAk6bN2h18QlKJGrTpynnXRpOEM23esc
sNqE7lkZYodVY8b2esj6nHvD+1mEBAHIpli1tMZvzbeKAKsdjhooTmMMgsTKs80l
s1fhIHUj4bMDqN322r/Auou7CEiwLWLOn1N158AaDcSoTNyxlOhttxjA83MIC2Jq
gKE8QCsdGCAqeV3FWx7vpfbtc58eu7wxb8RujL3faiH2NtXoYn+sAIYEu2UHCzbe
tCwdhEGSuPHPlriOP5ucM3IywLG33sEEcH4ogvfgpIncQWxjyo1UW6a94Zi2Zkvg
31d1Jjo77B6s4rXdZxhGADS5laOjfE/NrTz6B+5XiBzhBvsXXXus/l/2SB6UCqas
3eC1MKOz/VZw07uS5eYTK2vJ+nQ0MZaEsOtmvx4habV0qBFLH50alJrTPOYOqAZ1
IfNFoACwOYWiKcaOCGKyU4U1PuSfuKNImTtHd9rQ2UkDnuFpMRV9RJHN+QLIUgdS
zpao5xCNdKfQrbH/2GI2O1UYM+X387BXRemFhju5jOkPUoGgVnU8dUUeHBvWcfSa
zzwrrqkPkkXL1EdieVd+xkxRPrruvWigu+vmDIoCGlwHwAynBk//2x7P+TVPs6YW
CdArp4ajrTUuJPwNsJXfLC8XwnpGtF09fEKo5+gPCj/34JYDk2Hw2lEEF8Yvsk0G
wzSNHcG91qSLf7WVL3FiPZkDJLMVPC64sABq6WTxz5hvvMvXJva3M+Q7rJzmq+7l
3Q3WiF35V3fmPsXAdtghyrO3FuvkWsM5fAspx9kU+E//0JNMVy1MFet9PdTypk7j
aQCRWu5InyPLIaMEGnCZthXAoZ0gIlxjrUBDWKD0atGpADq457ZEseUuwLEn4mfC
cYxEH+v6u7ueZl9uWzsnenaizq45KLMPfgD8fok4NHi7JCQkEwIj10iVv+HOgnAQ
p0VclaPpxFv9NQJATH2BZk1FrTgeIXwbeXDZnV6VWy4G0l6QElPk4srVkTngvZ3D
Rjid1pNT/OGrvdqObTpTS9HIQ/znnxomilaZHtEys1Hm84iI6vXcwXKpB7OpSv0T
ahhbmOssaV+2YPfDN8suVb/M/QTR39M87M9MnuKmJ1kDShCWYRPGSnvMW+tzJdMi
BdTZxnVwkazKZeLcpQpsYn3dsTUYveAlCs99CYHFNZk+zyQwKuFP7UIDAGBp9lmK
NhJ5sA2tECRgB5rNT+ruQtB6O7e0bJMVzrEH7Vn4bdRc3XnR7zsL7gF9UU4tuCcg
jNgvhrz2Wlb8ys1ixLuNsWyLkeXTbehxPsdP3t7fLAt6nOxO8byrL8Jcpg6r2LoI
I9Ll+97cK8azhZLDxkS9Yhbm+3fkfEwtBa2ffNodlHG0N4IW7fOQ6chiQ+8j3zEd
S01ozXQikgIYGV41p9GPMp6nxxUngyFKIF/Oi5TJuQ9B0jhpiY+Di93MTee6CwMP
fiiF2wgW9aD7FSG0Z8p8kTo+llltmCoqpTbPIcap2VhxlMSB3ceZgabDZbqHB4Mg
EEgRnPSmCHlF3R8wRlT06nQlsxrsWqe0ffi4fxfDpTSrg9j0rzZyzCX06Q2PC7p2
E49l8gZ7vziiwhMfTwd6Q9E6tdDq9gUHBGyJ7RXiMjFAVF18CewabQ489pC6KfdA
6U4bdk3uZaAvkqZMdwXqbaypafjCJkIh/BedMo6G5Vy2H8nLOusubYq9f08O39nr
qUmdi5Phz+577saEe9b3kLja9IqUCDc1dELhSoIv/nnn/8x1SjhvnRnHoya0V8b8
6u4iRncH7MduZXsNhCVgUH+ySjOSuKI2xyZ4I2KzTgUMEb0po5XlolW8etSarjE1
mfWw5LFmRzbZmOJdn2SQXzN8zQIS1zJ662k/d+uNN7oAi36F/DiWMKwS8rCt+X12
XfHObhS0gwKdYoJKiIktU1JH5wct4abp3QcRKTyTYZD1bIp1+jb3h67mU8hbdmlr
3Cj5UxGIPcJW9a4v6/S5dufjDFTz/Tc5zwp+7Zv7HQrUVuR0JP9blf0Le5VdJ5x+
emKY5wXzo28h6YL3euAg4IHQaPJpQV9BiFXHT5N27gKoA+plyYHb/i+97CGJfXMo
o7i6eTVAZSr8FZT0V42rz92QS1UjQ3TrY1rIB1kNh7iBcpE9TubDDWyYm33+kQPD
vAkFkLrMzXxi8wzmxd2THn5ZpHj9TDCrMpxYX83fHzQ3Z3s83ThYHt5y5ht1erhg
yJkryZ08XE9eqXR1HOa0/mBpQvLo/fMgyBYFnQcbTgDetl8NecBRss4p/0TFihAS
jd0RttD9W1Uvr/N4QcUSIYHGJiczwPtwNufNq1DQoqGgTssSe81bKi2GN8gCQl0f
v9GydE9JaOw85eDTNIINmkh1jvKuMXCxzBp69LkwrAn3cUVI+0YPSHRNb1xWQXHb
ruQ8DgZ+woFabiV1SOGUtthT9uu0HJ7nGUMnOOCIb1AVf7lVoeEWgrMIETobwr49
CvArY32iWcEryDfOU4Z0224HKUCeSjZqKVBnVmYoCCCTNWIXivw62Gn+pucNhrNp
yPKNXxTtl6xD8wJn1mOVjd+rinr3841kxN+xS+VF8v4EZl5v8BJ8VTJBk727QLzH
hd4f4OijJHNAWEILI34ZycjpRbjOl9M5Zx3Sa3tlYfwUyLNriigEfCz1aZA1Ri1q
PsIZ+4QwxcW5hGy4gtehgXgfEX8tHQIWeYE4//1F9dIocVMow87JEWVXQhQVGfOp
4JRmKv2+veHXrBAjXFWsApEfhPYnQ7wX0gZgFhNjsAe9p6cn4Dvj1tXSRBtKpf/c
+MI0bvqZqSNNdYW1A2dw5xvAxRbSVHEtZXeaeO1PKZAyGaiT1Ovr8/MCLkmmc7OO
Lgs6JaUWg2bZouHKrqNSuuH6Zq3tFIQ1P5Cyu6hFB7ufLJVAj+p5sa7Z4DtciN99
XL0kmGVQYj03ppIKsnNFfImybauYv8UKWsFrgWzSuxdeWCNkZO4YHD2pnb1DAMze
YjBiq/FjZl4pAyLGdGwTWLMuNiMDwlHE8j8Q/aZxpyZCPtzQw7uAd4Nh5j105Apw
+3lsE42iNqVh8OTkArAqaEf13tpPU+IsPMu5s609qhx2iMH8SIiNu3Pk2T6u4DHw
kHbVZn/HLgxgKMdrXfMWo1ANCylym723kH0rOzULwrcUaLvqvNABQLizphVtuuHg
FMxoud8EOAeYXN1DtECkgw8+idi+fz+Jz778z5HFFqQiWT3dSdOWw9ba8iwIyRW2
Z56qA1lX2cPiHr8TYwP7PVyfhnI4JBEg84ZM0dBpXUXX+zhU4Cqeq+GXfLOWmmc2
yZMxHz+0rnph2DkirzcadRO3HFjk5kFlTzHklzZZUKMyRVFlAYD9vAafP054C9wc
iivWGSkkOQAgdPeYJCYAQS9nKdqHtu77yaVkZrUalkBcCTSmeFcfs2vr5zYawhle
TB2bKD0a0NYobpR1v5w3z+f9xcmApJlzODgOMJ/U3p0IEgjvHf+UiqOQVdv09iJO
+8K+KJo1v4wbREXI0ASDDC0OuKSFxtk9mbhma51Fa4MSS7RcYJXOoPdglRIczKry
OcaG9SrZzdYrUNjC5GrB8ITQw2EKnx/jExvlX9TZWMndBYdhwpfH0eZzy1xspQ47
86zhrkcyZpnQZlIp8mCMC26eOA9cAauv/3NBpdxMC4b3vuBvvhNtbvMf0sGdnItU
Yd5UxttPTMc17JBR+PUognS4mSLuxNLsxJcDVu0kl0uvVH7HxtbUAmNuXcOaAvBg
6IlX5iDL3v8C5GmevgUwRU4i8aPJYc8KkIdkgz4mYLDBeA/iZVrv7E3sjScItM4m
a/evb48wDwCrhOPkBFvlqjf7+3F2J68oj7nPJ8U9mZXmomGc1uhKJUreRYOycjjJ
VLWwX8jfDeKm1DNFYiHwOALbDejXGlaekEfnWuDmPEn5YPWK+4OzL27TZouYiAmn
v8dGaVC8iYbaHztPx0QBljgXmXuZlc4TgXzpFL79CIsPspiEjN26zz+M3oBmS+hN
Ky+9f0zq4zp0PKaz6zWHm0kA/qyJuM4IZpJ4dxqj5GRDNBo/5lHldZoly4mBItaP
18K8cvktg5uzE2RcvttnfVTXM4ahgtgPkRkdnA2sNh7RGvJKDMuy0RN5fazBy2aK
f8dOn6kQ+T8gSvC1kDAJqYCh+3XagwxDDahmnAXc1x92iYdXzId966W807uA7/i9
5yCcQ+g3bv2UDUYjv3Rtgnqm2mIw5qdosOH6pS16aIcchOCscuBKOK7shNrVTphm
cv4CkNHacvMWbvmXaDG289mROL1QpsPTNzcdsOw7hHx5zAdA5hG4v9aaSl9cBM6N
ZoI+VS12jmhGbGQm4Yckh9bVCrCxOiHnrEhlYHwgPJHT2zRPQW5fWxoX8ULxcO54
0vqFXfHCkDfVwJzzx/49dEZro1lsR13YcYBOZaspC/lq+8EbVomgtYrE4svRqjiH
0jJbVUOHYxmSwENXXFYetK+ieBwWyoadkpwTgnVlPDDS8kPasSNoW2aei5SjqdBi
LF7rPXBm/ch4+/+PG76K7qzgL/xuqhHz3f8Ct+Ltiuu3tEwvYNl4mXt57+oxh6g5
0qVKGcSiA3jvIMks3RRRbg5ki8/sniehnVqd+lpevef0r0AkFEK5KinVn8id1obv
6jBrHXQ5VBVhKAogrIL9BJ8t+sXuH4pRmnkrUUv47xYcPs18yh6vPRV0DeFf3kBb
Cf8eOi0a/6JgqP0PfXFqiNtijfg0GpIZ7C9St865vt7jTqTOzXMDTF8ThbYhljnL
Jm44tlkRL3ngyqRjn8CJAgHh8t8VsD/aXoIbvbEA+AUXoZG/geUIpxvkLEBInFSS
Au9fVG5rrAvUi6VKAEcKeLmYebp5/hYNnqZ6V9a8euppE3ZJdlt0NBx0LedH3+kG
kFxe6tcay8L2e/Yic/6FPKUTS+QOaV9wsAtTUah97cweilBMV8C3YCh54wiDu/AT
tTwxc2Tv+pPFW2GpeLaWNRkVD4pXLAoePqH81Z35KaMOSHinOnanhUji6i5F85dw
/54YcfWruYeslk5lfQ5dYynb4zIuNBCtpIv41xIoAJXjcA1HZXTNPgEHAYFWvK+b
eG/ttnQnCIlDSgJ1649JO+wlidaH7GbNjJaJSKjLsSnGgZUQPfyQxX5bkhlXy1FT
jxU3sW2rwDBLkV0Vrca8u78Y7N7KzADzrjKY7ioLNQO1dP7wsfpTn7svnouqHBgW
HmY/joQgnHRQHnIe+elXPz39sIYV/EevYKhw1oRNmmmdxwrVtuP7KJwg4Pz+0MpK
BQJiFTi9Ca/D7VO9We2OJr2ky73a0H9A1o+7IpOQChN9nlmFYY7ZnRs817XeL6F9
7/AhK8+IQxNbjVr+WNlGNxZ6KUDuhas4neV9y7CHbu85/4eeOMUjNYYWqaWKtHYB
6ZdOEnuwn4PpkUr9bOai80oQUBAPXLlHnAfccvRcPA9fp3KI6KAxIW0ryP//hpeQ
/BG9xWRvqSoIyPtOI+owwEaGWhG9mu8bxA5ZRdN4KNJBqomiP/SmnzOqB4EJjftW
XQlNBYc2Ypho6PswQmSFGZXEtOaS89uno7XshcoXaX8zp4xeKaTwPagXrfDdFroW
Vz7AWiKf+09vePKCyhlIDXE/OlqlkJAh5vx8LWKrbA1kV6D21G04mMX8sS0FutsI
Z7jo4l3w0p3aVPHYikh4HmzkVmIAJdFCAx0xdumZZv/6+21lRAF/s5+nzynTub2D
WbVAwpiBDr+rUwAjFH5fdk5QPdSt0vwZ9Ktiu9WpUjta7MkRDEA+TrVR5rZlbDgB
69ldcNBDxtqYHCnP2tjsNofAS//5hw7oGm9yy51nWobwjOgFO6dP2ni1D22pQCjX
p9scqKVMI1iz8KE7wPlORpnicB72PzGktDZA+I39Y1soDTYgkZsBQwWP1DIoFP+j
ycd3djR3PzXOPlec1/mdX2tgUyqXe3UZnwmJL5OXk1R1cMoLa9cWBLpNh4WRFhw8
YY2n2uQskILKWhlR3/U12QmMP8zmRIGxnSaOMt9lSm4xWPTLSk6QlgWU3sGGnhZv
Zks+z+g+saoFS9vPO4nTiMu6Kq+0UtXx0HGI1q9U+5VkxOttaf1q0HIYOapvQHpR
VNoPO1zp/7c24Hn/yag/yqZl3Bou+2ErmehFqqyDX/GMK9KYtTHkKUHdDj51SEvz
85cYDzAYOIMoD9fx4lEwBKrcM8rC7a+DJ2DZnoJ0HkZ8NWL4TybUSYz0CKzg00qE
5wURnyDer5/O1qtKvqJJbeKpWkATNpbH4zfOwREq1FuKN60ZJqa6Y9PKoC+dNjjy
SOBdRki/AXbVeh6r+GKvmh8xgusGyIWAGUzHxUZoJLWyrwXzCFBqn5RNzZ9q2pzL
Vm7AzqgH+3QKRNqnjTA4USBwPepzz8am8G+7KtyA4QoziJTk18AlawPYb1WK6NjM
xiF3vBSjvmV3yJoZ8j4n1xu0ppKdCH4PAgtUvdcS1ANSVJTEKSB28Q+l/FmRh0Sk
rhXzwdNEnM/dPRjOMZHfNkTIB396TfnLGcNvOjz5X80eNyQZnv/tABRgvKHr0GV1
Pe15j3hQcJjBxqfvlBA69kXsjFxGM+7Uuy6h8960VVG8gdR1ZvQOD6I5TGY9q7T0
amLP0pgWnA4hARbe6nqipiZj/j9XTP43h9cc5FuNKT3RPS4fh+CH4i9q2fKF47+E
+1f/fAP4ywn/VGp2dSrKuEIuzpNMw5eSv0eecdKnDMHIWuBXXsEJfTKDnsAOEH+c
1oI2opN1JgY3DhEU8CtpjsJYucit+FBuEvaoFKoP2pam/Z2swxAChpZonZnJBMwP
iqvO/Cq3jyrKhrumyeggi3axmndu+twDEKLRiDuaQyYnJAxzSe40PA3HATI189yA
Htuwmven3DRtXD9cHyYwvSMFbjpQVPCF7p45XeknCd8HzQs2qSJjOwdSaeW9i07L
ZMkKGTH4VmvGIq/eN+mEHf8tUqxVNo73MvHWdNLxznsh2aG2QybexKkIjU1M1Qmb
CJPX+f9x2Ida/oZKPIfiY3MD70M7xCwx+1gqSUaHYctFvDLt8pQ+HFQY+EKbTPY4
BIIi+VfmDl5zqQryx5mM01CA26UBdCAm/foVyqylbMClRf6105r8uVaMZrRZhiLl
2yldytHYZZTGJg45mmWWPjCjWBU274j1mvoau7e14WRRt5poDc2fx89vkYPJN3o6
cnx/az7xajQUHiEQ+zopSyZ8b+2lArIA59pH1zc5u7845MSdp01TN76MUaHQc+qz
cNyQGNBhkvU+erO+N/oTgtDN+jIB/RvzCnH/VSBMgaYdSl6rWMUPKxX4itbvaUID
kzJ3aibU42b5cu0H2UYx4kBih5Y/cngdxwlL84TjQa8DP4jaR9jIKI4A2ZcjHVkc
2IiLrvQQ1tln4vmRN2+VryKHujjvSkLR/6bdPCG2mjIEAQFTiT1AzpaEcYU0JWV/
BUM7A5F/CwrHEHbgKt1VJFMgxW9hYrVo4n2Ue+B28W2YF+9o6n+iPaoGNNltJRMh
/7hVmhNDxg2mlNbOS6FSUVk3XsmdL3cYwSSChvcg3WZ3JVTcvmYXDsYctVdqaBXR
U7v0PNDQmccP7UpDizW3YDOiPHeLRyGCJDd8VGhvkY7v66UAOXuS1C3AElFKfHiy
u9Z6Z2Z4RIclsCR7VCfHVJwK7J8VS6VYmOX2HKGuczpDgWT9khQaArt+uZDCrtoU
/eLGqWtR90i/LtbN81BNupnvJJ/lGVzNT8Dh6ExE88LqwENpcN3m+vO/Qjaeo3rI
5PopyCWEJbEOD2xhTRXYMis0qKlT5dvS+SHtDez3xgsYt+EcwT/XjCYgspHp478r
EO2sQqjtk9qn0PzNsXAtBQQGw+zsP28qQwTBItsmWOCkzOpK+ltLXyEdihMeu1Gi
8VPzQx7Hz55eGl4iINoAsGgYguGbYZuYFxXseZ2x01JnnFpZP/+yfL7xEz2+EQOy
Me1ZFFC+HNBPiycltoCeN/wmsKdJv8BBLxyuBU49SPYjT2t67AJP663/srXywyMG
8ktyoIKl2Uze8gNAvk2LNx3WZmInRMeI1gQDHJki4qbGqMgIcL5wpZWs+F2xvSI6
EGLFCJBCnrgcoTBKkM/fbXbNS0KgJNj56i0yuKa2ohjGr03jZBp4oE+tqjsMprtz
rhzS8JY8Hu6CAlW8WdCMuTIAjWsbFl9LU8R0jROm6m89XrxMQtr72Ms/7ZyV1LuZ
pJwwlqahyX8lF/KSTLygfvdi5A17YuEtpJIVKKWOLVv1JfwY9attpCa7HzlJkIWy
nvYwraVpM2Hp1tEudkfvFsjBGD5lul93UexwyQdFeSsoUIqGwLXmQN3RcFwwN9p/
5PuyGcaD7jnhHk0hJEjF66YKAaQDsLI+Tojfu30I0NdPBcjogMFKcutx7FmAQU31
g8FFluUcwqNu0xCtQBIcqgTpdt4A0XemPKYJ4VJlswqurtsu/GCSaQ6yRbPrBDNq
kpeT1uzyYrSraFmac2UAETE/5gzag175pGfdnbbsIncoSPvHcGcdT5eLeRMXJD9C
IMDTrdoMv5Btk3PwwOKZ6TLVuq6fGK/HWPZEiJe0H5Nwpfo4VFF61wSwmqbYtweg
JAS4JuBlg1cs85z7MT0l3myV5pcfEpqjtNOfW7uiGp0+NNEy7AMyZVrGmgQTyGJU
P7rYfkND329RM+uhpX2zWcw4oM/C+imW/MR7ONfOOZuIDUKiQw504c6mXg+VswEV
5EaGIwDMc2hShnJ7z4dmqA7Vir31BXL3K0r1A/BKohjjBbRhE42lVbe8ZSbjb9ex
Ai0vj/YIqoawwT5+p5ikFexnb3nCQp6ZlkQZQbhCKQ+wxhBA5w+g82t2cwEduxm0
iZz6DE8FsxNtAGppIv5Y+jggHqKzujUolZ/vyd5yyGxyrl+ijdOQMoO7QmeH2cAJ
8jHamv6V41r5Ve+383m4La/i8li/0rv1QZ6j5QvZGH2FBGiEe7d0wu70IeJ8XXOx
nNFtv8cYAmsGIYV1ERQn53o0WMoRX6gE7YTluxIfca224lhaQWAkFOlfZ25PPSaq
JCwQgcoYtRlzIIuqJRbpEkHVQvITYaxDAgywf3sX1fZW9LfyIXf7fBkyotnV4Gd1
QBNiLTdZp/OJBAhMifP7Q5Jdr9kAx6XQlksLMElEzuroNG2prtrqhNVfGBU1YHxu
y00uwiq26jfOCMJu86nHV/E72tYkfl+9odn+tKdcdoc+SXi4WCY8IQt4HuelWOqh
GlGVqiazJBA1CY8wYcLaJYEyk9L/JpbLL9WpITlEAqV791428hcvqzWwhFiff6a+
hMRsdvBR1wxwJu1gpjwZgL+vZaAP8jMVJIqF9i3yx2MIPdxOVU+j+JlRpsx6PlXQ
YmsXw9LCKnlg9R4ojSIzqFqY2kxIQc9gxLSZeH77A89sSbtEhrl4HXFjboqc9gj8
iLxhlP7maG5kaevlnKbI7dQ0UBy51khdJGPDXlmsbj7dcAL24rrbSt+DPnsQUPFl
1Kl3EJoCt8HfShB63XruaSP0pc6CImvKBve37+jN9e/y6Vx1jDs2yKmun/pa69+a
jKmsmkl5nCUwFmyOXh1mDd/XSM5foaQ8kxlegNmhvEIVh98MWcsqtBoGLvh4oo+b
ceoMaV8YFIsvvedkKyHgBpQoe8tgi9cFi0ygoFJv9QJPiPVgAEogBakLyy3zsqCp
pEo23GleTBKyVc8WHCapQ+FH871EreS3DG4IO6Vgl6znRDvnJoXnsNyXvAkSP4KS
kW3r1/zLPFzEVVgyZDLIIRKa+ICAY6HiuBZZX+vbq6m9V3TSaCzEG6fd6vqLD48p
hpCVrkpphDZduAQito5h4W+CasYoj4qLwSb2TulSIebCZthb1Y4hKj0x80/jAx7G
BY8CanxSXnRoemwTJi0Wr0JQCB7f6RnLJPXmlcwXnlxfuR1jQNdClxRiELNHODD+
LD8GRpbPWrRBdV7Cw8X+uwdS64aSrBu7xc6PK8rR0Dhu7ixxV+wp99/mBwlfJu8F
0i7itdqLhau/4Dypx0O3JS/Amu7a3qJw4nstksBwhkRvMOGA3YXwP9lJ7845oEpR
v6QRoRgqZOdTQuWxhfOT8/xSo+pXsp4yHsNxqOcQ3WZQCyBBLNBLmSGJwBNcLmuR
2LMzL8yihCvhoTUm0j/CyFQTvytWYeW1aTatclyM/ivcV1G7OuCVWKgN2qhqvQrd
bKQJhzb4Eed0yt98SQ2YdVwHe8dbFOedyt257HaT95QxpsYT1sXZhQuflz9DtYTb
WVC/p+hDCXJLvMYGEf91aNR5oVtggEbXPeDYlEKc1bGoqLAp4lxNZjL3T5BOSY+H
0o65NbzOHp+tgBRHrivTXyuBNjM0thK5ZDXzbIqNZZ0UQD7OEYQGaOr1ltshjbr8
G4BpEo4e1L/3DNKjICJ+zL2q6BsNSIZPhvFb5HCJ7FUiy4FdSissSqGU/QaeOa7q
rQWUADrMopEmpfwEtTYItbKi2Az219tvh94YU7NZJrwq+U8g1zF4HsaAqCOTTwEt
beDBEka7nHg02p4XUWX4nTMk79DDaRNB89luXMMTSGpuL43ESK+0P2UVfahpVZtF
fm8ULJ45mWUeNxYjxqXpUpqbf05tDtRMvFsARZkh4yy1gsP96Iw67+zlZpl8S1dw
iVoll5RpNphjLlgq7qno2ovrmkEgGoJXcsYaIk+AiVzXRgqkQFxjklorbKVaM1F2
NhtxHgaex1/d0Vy8qdbKMsD8N3RvIuiT7NQTAdXJMaj5GvsdlgfsEUNyUf+LjPr1
vne2J2cCtDkWgVSx1vLfch6r24oOJhVrI/Uuivt4Ktm9OHmhUHDGxi1muY2oWjcq
Efr/FoSILPkoIlsc2jenscFMaph33OHcoFl4Q19MXpEnFVrwPhxVjYggC+K4FGWn
AwpkIFZFfRkFeaLM3DQrmprEqHsCa3X01mCEUk7lH33EEw2VjO61bt/GJ6wJ1nw8
FS5l55SCR7fV6IRqfeeVewNYKewNvG4HsE83tpAkv4rct3LOyfQtq7duMQ8aidRQ
xCrZHNRr6IHP6d+0bwp8ICQDdZwLKA+xTgtffj/dbCjVx8E3JKsNAeWzK2xor135
2Fy6EbuRY6dtQzwlTArNkXFDNrLgSjOL0a15KKWAV8WNZMTRDpWbQZcK63McOh7x
0JcBy0KxysSei9ZxgBdZBkfwQUQphj9rac86uqwbDm8gqYOuZxbHKiwKrMKl0eAC
cxCpLgMWCVraw2d9Nu1qhitFS8HFew6yLzq6YC+FSb3cBb3Wots5vgDjAdjFj2Av
J5FPR4Bj9dA61rKM+0dSNHrAa6M2OwrHRy+qQpxVsX1MJIxf2JRVBIli3bfzawWx
LkwniLbOaMdulIPxKia7LDjmz5PKIrmSd8s4RppGYvJr7HcFM6/LrF6eLz5LlFNt
pjnanKA1qSASuUA9mKmENjMdErdoXgKm1/SkB/TxmUbCHFX3EJZrwOT+3WURhUkI
z+kW+rF4b6DHNhhBXEtEUviGyPtSNmqHwj6WJvxd5lkmcz0Gk06dEA+L9QcGbq7o
nV61FFBRc3CvzoEhLC81NU7yL20G2d1HkRixX8eDlnVKWMRAdwKbVN8sd7TgFJGK
Ma81DMrj/3G4a0TG0pM0MWhTJO4JL55PDZYxhXbgHf6Xyy5/D7DV/m+1ZG7hkp1w
p7NUejZo8iYvBJKAZcoYtIa2sayVWpMHR7lN8tgNsG5JYsLM2nZCblMCcHz4LwGs
yGg4y/FEiqiHqEhYkxfE/JjWe36eFxacNf4o9j7/r29ZZ+NQJHSktqCFkudwofTc
kFDW4DT5tzi7PNsPQUa80t8V6fy0YibHR+qhX28qYk2JAIaTQT+1r41pNlADnx1w
ay7Z/gngZg2FRB4v4gdAmn8AG+2EYlBF1/rB1KhL4wAP1DMSMRE8eaqOQGQUUeQ9
k/YBeCxVTzri66Lvltft/v+i8hv49lXQEHQAG9P7k66FCpi8kTcdeYXtZeIJix3j
y7yonMcrjqzR2Hgy4K65BT4liSOYUgjT0ia5Cw8l9iLUaCNUbInThiQR7XH9eSu9
Zovwh8X7ro2ucLumIZRxjXLiYQ4scY5KFT/valZi6YfzW3GF2CKqZud3J2PoyGYT
LpjWbMRQtxnF7HF9SMxhqWyISsx6ETTPGlvr+03DP97Z/4aobuUsL1cwc7Cdy5Uf
ZAVosYUr08ZIOMpSUwKxOGSTv/wJtIsRXMTe7bkSBHHPk6WF1NhHke9ohpFc0CQf
HRMSdqTXbJ7XP/Uii7eiyHDnKfeGgq8hACJsS4cnYXqSEdp6CvY0vptL+EzbCQf4
ztFhBFbHPwkKIGJN1Wix6l6mYxpj4XsIGDAbki+k9yCrdWKS0dDcGud50byITAaa
ojpQf0GATLOo2mP/Z595bYw5tgu3lrZSjkHNYB6sOuRLi7D2NAUgjHF5YqDZtbl8
wth8U/2vwpMez1ycFuCPQZCtoKKbhh4KQlvBsermG6f4i42vzNRI8cz4YBwHtuTv
YxHK/ZljFFD37GtCo8UMJb2HeOaoEHx9SuN0PyfNxrPD3syspHktqEcaybyQkb8l
WMQd0m2n3KTYcf8AQQfzIXZx9J7/3ThEEabqUNrBuoIHa2vQ2fh8QXnk3E0u01uA
kLcLlTpulwmTBndQSmFSTo5d/p3JjxDvjT50CUX/5xULVzzX7vcmX0sF8f7x9TNX
6eGoapkqOTyAmFGRrvMXr0GPzf3c9DrOIbWS0YP1vF6NPdTUdexda/RkrbeWnhCf
SulqXPriwcUCcje8CLKxTaaeajRH4gcBYdQwxXhHvTl7Qr734Vq9mhmzGyyyNTys
ZlM5eflnzI2ly58I27Du5SAJ4u3nuyirIxLg8o9meiZ8u3e7HUtGp3uEix6bfkEV
khtaiCsi9XnSmrbR6c+rJSbJWRG2Njl+Z0gkDYIiQN7hcRMC4TzWFdUPhPRvuIic
ZdYSw1juhcI6x0gWO2VZ6IGfIkbvlXZsj0MLqeycvfuTX5z0oZltmpcrP74/9fGi
w6e2f1Pr7jM+S1fsALOQoTM47559pFNCzwA//Q9Qt0RnnVXjzprxFlwEo9EurCoP
PgeiSeq/Dtb6skt6F61jCJ/VC285G4Ca+gKnfTh0EoSzAfFw2B050sAPR0bfCFT2
obFvyWg7oLln71HSBRL4jU3p0XY2vTuFxVnH1cNGIY/wYhO15LxTWvBVoJqXDbz4
AR10CgasVHV0ZzTjg7rks7DBrsALSTVBvTw7UwqxZErBKhCfVPhcxOUXnmENiVoi
dTPHSUxecmkHKquVpqjbgvbnw1bptj24pMNEfmYSmmH/Jh+rGsLqs1eHALMYwxJ9
PaocCongOMudd1HebuF+uvMvfJZxOg/7Q1RfNRfX3ebRN0uo4l4u88iMpbhPOpDK
3ka0Td+WL633KwR76ozREH6X0VEgnDkBX56TwSDHx1bZE4SfVrgnHzlNRUkLqgEC
taU0ix2yMId48kNOosyAdChYMTVTQ3OoVV+6sdZA1fo8xDSmkj12SJG78Nex0LHT
xdRWmzO7obVCHi5AtneUjcaL0P2vf83NJkZogg/JY+p3uZmn1TJ+S2bl/J0sxzRM
7dbA6Qpp8VdAK5pMQ17/MfgFsj4rW9bc0DOuJcOBcep6RBMt2FQnn74s8AkN5Znz
OXTimlf7kwx36aQnUfIvzV8I67CbI0d7/34ITm09agx2BZ6rW3SHc8VmPOmWuHpV
uOTT8vrskOoYlOYTOR+giMoyEszcKPeVbHobs5o7bAoWXruG7XyuIHThecunwrej
MhO7y2WlkknFrzBNWybb7MkqVpOlonjRlUuwpdU4wxZP3kbw247p/y9JAKBMiuvC
A2/eLVbjbbUpW3sI9HzE1+xszakWSmfS9YXh9fbtiM1tiG4zo+9cQqBYRR/MSAbF
BGs+sHbmtFXxoI5/DZVg/oRWCZJ6kx0i094AS8rURASo3pNYcWuwW5o0eg5zYtDX
8BEDxlukl3qaSBUmHlVG/YGAwLlPpBRQn8a/JUNi8z37M8CHlgVM1JY5c7MPOnbr
//NgFrrkKeaXdYRt2HRJjckRRSilProywB0P6qbUdYzb17hPUiFvUG3ECIvunqBz
4pZiMDA8/Yo9izKyx9ZUSUc6ZbllTo75dQ0YFt+Ag1snKoZr1q/4De9yzM5aSbur
KBLfJ0RzpNsc0+TwmtaUsP/OXKaPH6OlOgdxdJpMUFRaEzOn0Qntv0E+SGkX4yE/
w23kCvbKFTCWL4kjwtgN1OgtxO8ID/8BF/pGRNAjGjz4vnsjFow2NRJZsVEmdEl4
HNCSTFmTDsbuEFC9GLEXCRv6WrH53+FWH0zS0B+JTmLyK9V1nK13XjyXFd+HTgSJ
Bfv8sCQONZarJjFZXlOo6oKlfpA+Azm373EIudlh4FrdoFAzkvwzy/dtPT4nEBlZ
4awa+gRBRcgvP2zJal7D3/vY/FQiskT0hbhhviOjz9PnuAQeJKXciiDiS9MbHJ2U
V6kdhLhfqQOopvRUZ6IXT6sziLBFlhEf1XsmR4+ueZr3R2ah+8Rp4cQPg7M+1U35
lzTJxup9i8v5DNxWnIyTOM7UN4nGevIbXfgBY4YMiwj5/TLKOy6kTkb1z3s0CcWA
Ac7GpiCEHLOPYhXvVhZyNiC74H12QCVrZcN5zmvvs+xO6EkinVfTCO2wB3e5/hhq
p7P4lxX/VaqICfmDCBeRZGTa3hSueQyopHx69d46IS9mQnN+OtwRUw6jjm84fm+6
nO8gDMGIU1k4u8UwIWM7nC5tD930IR4hJiQvgRmUH6mP4npjlriYZuJ0lG3/fJeM
ZMB2KrWo/yVS1PEmP4k6bkNQ+sSNgAkHERbFvzPmxVGznj5MaMAwiGRfJLYOykX8
G7Iv/xXd7iH4gFIx14xbzwtAEuIA2mJJ5HRt7AWroQTUlHom6+9EPo6Ewyzh9uFO
IsdXgH5Sbr0wOrA0Tot1ot3LSMf7ohn75IsCn1z1CS/1BbUkc0+dOP9808Yqz9YG
knL7M+dWnsPlU0mmTDEYXRXUulecwN7V47hB8WDYStuHBOPmQGCmATujar28LNfy
T7zTziTPfJc3YMzIGDyzraxntfKlvZqtbD/C8BLIqOSFZbeXgS+0IgpsR1xJ4xCg
jcF1E5qhrt3nOYvzxjR+5SvAGzc+ZHUNIpqU3AeNAN5GuS/fDliiQvUVwPim8YN7
4MA6XmBt1Aq2unau/GqAnSSJHBvvZlShljSxBiAF9GS/IUxX94ax+6MzKnUvxrpT
i1xq7bA5XoGUAF3mQ8jn/yxqU8rsNZ7jQZhY9yurs1MVdMk/hlmJRL0oQSYmc0yk
mzT1OtJCubuY8kay/DBd60F0I4YpklFob7TqQY5IdHeSXobx70kFtYKFrxp8Zn3X
CHkx2S7Zpxmj871sDv68nb5CaPi3kHkl2cpwosSoqHvbCoGVx4h2/404zvKiO6xG
mRTBrwvXC1vJkLStDKMxwUPxRncXqsIa8rI/+U4baBceJB6E52h0TfxIRNqzm/lF
HreGe/hE2H5qv6LHR2iirVD3yW3KycJblEgkhHd997wxXMgFuoYq/0Bm/mB79zR7
SH9pVCmseRh+AXBkDTsrcayR0TXJZuphADkOKuti4bS+gSWLcM1MQVHja/WXm5wD
GrOBUHglgX+5JqtQIf9XYdPV3mtz25SSFJErqpUeoI+RN8ufXo7QRY+qWh/9yUlI
Tr0CVhPzBpnzrqenCopDBjCZFfFykenaEKfq7YS243BXxyxHHC8vEn8X4KqcZDBF
oxotjd74zhwkbNoU0TbF81J7PjeBua+PC47iWFog83e/p4VFtFDwOn7rRF4seKfv
qE19/CBNP3URR0eRgKfyKSwXA2QvvwNsJpCgjj/oOjY2KKdzMWZNRAc1A5L/wC9p
lw2rVmIuvXfvtDJeGCDCQRIFUZAU2QJu1QBweMFtgrY5HACayJaOiCvF470KViHs
Wz8GwoTMZr9c7UOfRqIv0pXHBsPCmljU5T9tt3WEFeJYzUCZ/G+qCtkIkQ3lNfWV
1asDrQpp9nPxMS9DQ9YDt78P2ntk9LjTib8qgoH48ajzN33CuVClb7/vzGHXxLxx
2rSF3CU4PIy6IEMzicL/Y4LsqtRVKq/NxT89C4JrfKpmoXHx/hCXAvFRSFdv0Awm
8ELiQPcNaRUKCDa07lxPbFjTPcOzBeBnb+hofZ/DwAHu3SenV9AT+rPkAi9eygbG
c6vDngyAHE2Wq8S3u+w6viz8JBOHwF+QjytJapHPsxus2LfX6CViArzqAj+LVTnI
eFspKiWwRaEe1CGA/Pl8hubsl12rlzR4ojHiNPlj/y/BxCTav4S78QL7LvEaITCS
l2BBfuUFL4F31iWZHT+a0d3YsXxZUfP2ku2HDA9PtUuWZJmad5p3RKwj4XkdPEqX
oOjiD3FrdK5uRMyswHD78VILULLn0uH1urwExsPt5l5hRtFNroyTOGhGuqt38i+S
l5H30xBPnb3ws5+sIjBX9HJUJB1jDHYXIv6bol8FN07eTmluRhdtzXgOqOS9NKd8
jDxT45c11gKDTcF0djLk6bZQCaqZauWZ6VtcUMlwNmolFcwKeiBbwElVfJpa2WEY
RoGn7miBUMZFIhRmA2cH9LfyY2dN1e13QLB/+UKp4HvMTNPMGOAhV+dzo/O9kjt6
GRhP5DTBDODVuJ5Udh/a6umqZ7ER4GBcSn1TOEYDMRQ7sEyw+d5gLzlInBeEsw9F
efKE+5yqDCCA4DzBXO20iKIDrXTGZMMGjfnKrMpEk+7MOCX7lH2Ra+dJmoxww5Cr
5dufzcy1Kq5i5jPfanoYWu1/rURWc9RJdjaz/G4NEtxiYsadpGsPJtPr+hgG/ZZA
997QPEMqDumL+bhszzTeS6BbLPKeMQBOw14KXfme8lZpwSjUmmirGr1geQy0tEyP
qd1zZSJNwjtukEc/T7uqKwVvKp4fnQrVE0buZZ6H9wHml/15EnM4q07BGnKaL/2F
CqVzCjQX1BuqrdJ/LsqVAmBnRmq9pYXrQ5pD4NHCuKz4a/pVHIFDJF55U48bnOR1
krOI3ExBtr8OxuNV5axPvb3+M66O2nVY7qyyJiVfifQgaKvxdiuey+NTRHmqJtlt
oUwe+a7FZazFGdLREclNNFO/MBdOq2VHWV3RiC4N4ZUbxdEl2e8mqjnZhsgw5IvF
ObordKRIP63NtdpNJpOloFGhGpllcBPzUPfoQ61OktEoJvDmrxo2HlsA3IphTc5R
C3WIkhkdqY/a+0UPiGCPUNiZAF2XXHXJQVHWBhIYEaD7UMZ1gTnb2UQ7MOjw4e4q
ncIN/SNTTs8PQa/M+44e3xzFIoD6QtXMyf3QQaHi+ztjodLp31hqGLk6jY7hQTIX
3yapCTsMaaMJN4iuAB0Erd1ifkp2mSXfGP9iYOcTBImxbX+55Q4rpRJHXgutaVir
YZnkLpOmlr5BRIlhY1t0bOljtb7njJLaxqvIyE5V/UQiuTlK3AlOrNi1rUjNv+WE
Cet6LPl3wappc9Q+rhi8BijqqKUTj1OG7rFIBc+soyQjlTuXjn0q/bNwJi7qRLfs
OXCdY2gFnKCMFLuH/BanTOJ6yr/JWNtKKVEBg5MS2p0S7AP83E7CB24ahQpTmXXa
InnVWGM3W5jtqdVBG2Mg/gW8w+Za3DfVTHtCYoXd7gMRApXg4XiQRAcGPibBvXQK
14pL54vuZCQOj9JDtANUbo+29XYW5i+SDcHT09TS0it+oFvkbmCJp58/sv4Oiden
qhEDTGQ5nso7nktig1u3Vgm0w45B+Hk6d0ugS7xtLPNuFMy//UNU8tt2liZmw2Li
7Ba1NFg68ER2qI59ApgxTlIow2+JRN+TM2AopbjEOlEJHg5ylG71xxSfEG52aOS8
xsRBPo6FiKBb+vxjUPaFCCh2SbDlKRf+frqYZ5phBViKdfA0rgOD4buKKgDKp7tV
NKlhzCT4noGJ4LcGumrhX6+KZ3Oy4d5vMbWKuqVWisMRGfUGKx49lX1dNPrvn/Ob
pScV5OzDW2AfxLiK4wy4QGuhreK7T6fmefxByecES5jQnW6M+/O7/Ai3F2Ebj+ZD
GWsThe8U+yUyKeP9qmVsIuBCNc7pLIeFZFegqANoHyFmJ3qNgznF+2r24JAMBHko
dtIqd3CCJGfds9OwFOi3pNSpLfMBnsC8BHoMC0DPCkc2GV7wk/sDuRmkqGAV5gMP
/vnmup3Qzk+hiymOAUf5N6GWfpcltxze5bzCxwykPnyetX5rglgIT8Vse2oWrFoi
zMEA0uA8xnAu/8ivsd9k+lgqIXLUQ1/VEkDy9hg83+bO24MeKQcUSNRQJxoLBfAr
1wynlUXC6GBx+rsvqM3dQ8n3QoAPxuZyJiMGyUSt75aHUQ2mXNj6O7YHvNJKs8my
SWbTUcPT9up4iA9T5T0yQKmnaOODRS726eOSDkdNa2DwBrb/RCOMfJeTY9UoFYux
EXHuWmbChb+ILKNgs85HqKHUp94NvAUwHrSxEUS55twQ7W/k9T9WHF+BqON+i30T
81BUVjHYL0uinwd4l1Vh9g3I4TJnMMft0bG15zZVvqeBuzQCqfAp/RwU3oYVhFyA
id3x+JB3k43wUWcO29XSTHrwdd0SG6Vz1x79d8PhSj5GOxKeS7AdTPNyNTSudhwI
G4w53K2ro+ahPK7QYJvmtgz6pxD22ms8bven3kJsghxhorRHsjcRHoDCvu3uoJU3
2nJ1Px0m38UC/w4zQ6PKnk1n/dDJhWa2e+p/RkkIhf1nv02TYpVRGSvVwZS21wlH
cCaMtj4ExW8Ff8AWzWOXLoI/LiRqu83YkRCCpPsHVfksb02bcHmuEFtg637I34pj
I9C8UqH3XucrtXavy4ZVzn+XldeZkEBbEenuI0NKmAKOZ0CzPqkrj67OcXA4jkUg
jUMKJrZnGy/Or7LKgQCL1Fo9eBb/OAMLBO/sujSLMgLkDp6XSS/zCZ07/0SEELps
wp19QRm1APB0+AwCSN7ROOj3VyRbs9mlYtLfDD2ULM9ijGB4ZbB2YrMXiBVmwlYL
plFmO3+0rNfZiDyIsQJ7kkIeAeXHCEbc1GJ+nD9QuEg6eLN0Xubf/DUwCO4o9bFF
Wy4I1bOrZM7XORrpUs2UBg3mLnCnrOVAvanZmVVyL+o3hMhF68he4DITc/ZLW3I/
8QmZqVwCJYy7to81scDidbKly4T+umq466+Y9ytetnsnPUaFw1sGWu5+R6juaKtc
oqRTORIoujzZqOJ7ob8LipdenngJlz/en3Q0DVPjXbyCAMugiVJU/t1+gDjDBnjZ
gXKnFAhYxVxyAHxChpJ0fLHBnA/pUuRmTSaCdX0BxVnD8LoMFhZVhaKa0vJBBRqu
v77sSX4OZfisiX8rCvbJdOiatLN9LZq2MIOYe5srbSonFLm3IN+sXVNVlCpeBiRF
4oJJUDcxk3R8aOmk3e0Gs4OWBKiqTXtcEKgX01rB4xqoagt1i0J9cFCx5tSKi0KG
AtrwkN4cfyDdtwBPzUoNbdY6X6pchhv90Rab1Wzuc9MyaaKC7zGPpTzSl1vLb3Za
NZSO3MKvILdAjzBHqBfTwPd8XzBrqHKF/qrhOjHdglu9sGP4/tF8auj8G4AOaXC0
JnKmX+ihY4f2dJ1bOBKNT2VqZjmzkFDnTaLe1Ivrdp5GopJcpVI8LqUsJ9lWMk2K
RIkk3PeknSN6y3OmhwDkjvY9cfYBS58MPfjEUlp3s3b3Ahpg2LAaai2d8p9G6Sek
DIazRwCsH5yJYLWMu3HuLHpYk6RG1lmlDzexI/Vg2K9dTF/TlPrMM1GUsjg996yS
cUHFJcCWzDLKy2LGYpZp/wL9wA3P762gYw3705MdXOBVBbzEo3zaigJzCJQvoNG+
42hIhzqAMcocJgsaLBe38yFv2A3PqGIcIyGTNimMhvllTSNMQWyAB8nSw1Ram0ze
n335YFsmmIVLYCJAXGNmgRf5m39rLSS6UcC/BJuMYILiP9I6pKD/MFYcEQU0AY3R
hnzykq0OcwcxSwSeNhqfzY5dN6qUpFqsqcdsOgRP0EMHoviVIpPTy8qlZfJ2ywun
8eenrbCGjmDNwyF+u/c9GptGfYyD+E/ZtXIvnWEbYJVFC86g07eTIIfesFr7b7MD
qw5kfB7tHYiGW3ehtoWJX49mFX6EZhDN7VT6brLcFDrMeGF2LF7wOsyOds2BRFWY
Xb3YS0feTFRQJO55V2/4zW5CJ0f0P3s/Q0V5ymU0k2fRw2YieTCTfTwu4xqhxxAV
OSn6QGB6Tl5XshAzl/ADL+0SZnEncnts5iFq/VdB+S8sEUUU4QYHhizg4cQ40E1i
VsU7iFYwCIoX3cexwQHFf28EjDsDJCTxdfvCAvIc7nCRyRv6TDd/3Tqfm1VLYFus
SIWBv8wTfOopIV15PYVRaBWotj6CdR8dNbVYxUlZFXIuVGtEWu6Ka5r34KBegDy7
DzyiNr/plUwiuDlfcCFepIumQIkMj6Y9ry6m71sM0DwAHqeNEHRQKQh8JCAgJRci
NTfCqKnNzEJO+92+G2+x1oaNQJwTd1UfkvP+1erRqy/hjugJ1oUM2h3UJzO6/qmA
/7n4olEq1RuxSxmvK+uwtM/w/ersiChRhNj5JQrMo86lXKcqp4SBFMW4E1r/hIeR
6G7K2lITOETaqkSzbopBX+defYDwnGFZDLNqohfUW/tQBcA1kqH/YhuKGmF7LtC8
upBJrKj5fWe85lnLwGi/EhHtCzzYTpD2llC0IUe6zP9/uXo1nzmAvduR1lvAmoE7
HssML59OsnA66fQG0bALYTdHqlW16/CNlXJeFFF60gcQVgW7WBT4u/mOGmyWjc4f
3tDwp7Eg+6N27f8EuZvbiRbVcFxHe46n+k9VFJ5+wh0EVOeDAdfbYn+n03mXl3Y5
NtdkAxkeM5bKEoxCuhlrLEMciis6WBVvmDdr5BAYvEUH7Uylif/+4RudWZmFs8Da
CKFbZsNJxKYESEj4VVDUoym2ZeYyrftYRsXrItgejeCb3pAhCbIWMg1Wady79K7s
EvdFLjUzJiKuwxwJEmYFvi2Nl/xMKUuLwBIsoZBlC0JCRLgTn+a9oPz6MiI4co6v
pIm0GMicyDQdCb2OMB/Q9MgEXqxGFWkNb4QZ5VlmmpJqkDi92X5U1JxUJDiYeAho
PtVJ6clmJc0A0HGLYhXJDxxOZ4RqjPKJGd1wQs95V/Zp+3aa3uHTj4sMqQDm1d3R
pS6o3zKVWdEMDBVVGERzo+wSbU+3bzJjCgR8fYSFgOTB4Vu7VHLI4ajGj2pMnCWI
NZdw33Wdy4irm8JfqS/CNFncBpko00X5RyInx6h8tPtaJD3Bp8E/kzsbZKmV6D0E
c3Q8Ze72QV32z7v/r0LOVCHdGdUH/tYWPjyDO6SFNjEd8PP/pSKWjjmvUo9/lUad
dTubcgxBbxYXitxjq/Ye8zfO3mGSvuMHYCqKNAFYY1gMTY/k+ymAFJyALnbsAXj/
C0IjD90Ge9q+w0PtlUs0mDYnDR9PTqkM6wVUT3rngMrflOKXjrVoEO1OkYQfbNe8
oT7YyDunOOA6os3piQQZC8tE7CpImQV3t/Do7rJqWDN1dLLyuR40FHxGjIpuznmG
fyw/3aFuOV4vT87QU+JFv+aQt1tHMTWzeJTYtdWlfjt8SFzEPF0XAvXt/S0Im+LP
2BjCXlgwlbscDWp4VzUUsHK2w4VMX16kIOLqMHByAo4oPbTWCnJVyFLfAAMp8JkS
VW6YCH2hcwcRnBYp41BsnM9YL9pzcN6RW7B4v3oed4K/p8qTo2+YlLpc0GjTtznf
344oaxPDWeSkDaPtmlCO95fPoFM5snLYFtHnaP975dSWCUQq/V8JH4hPJGXn9x7i
v8svfUXOV71Ul2w2tW3hvM1P6LgA5fknvxKvwQWPcYbbdUwie7TYlAmc8Jw+nIwZ
9T802uIADmMCtvDZNqapGc4VQAe4iahmU9YoHU6Xg4cKm8lC2lKi21UmyeIdzI1V
xdyxSmrMSxhPHVYpaM68w8n0zn+Pm9OHjHWXG9KXDIFeXVe3pdvTtMj9mGm1OId9
DhD1Hsx1+hAlQl9j4lrV2WkAiJRiPWJjk5vxN9BZhDQtqQ0ewQH1T96mL1iYpkzz
NIu4jG8rLHadpxWxERLXez3TfmSRhAlY/ZYCHoEmp59dyptFN37wd4sny6vdWnGt
gcQ01uZvCXgC9YbQFiL67MyTdGFGjHBIH3PCsjQ3jLBtFQVRZeJwuAKhBmZSbrLP
5uC1GvZUEh1/VNWiTLGYYznAQqdbICoqwrcSCmiQwfsAeODEye8EpcItqrdaVuB9
cIWutYqzOE3fAQv+50HwQWz9GsQtaC9+SGubv8GTZRpaKsL2GEsyLc7H6rCT2Bve
HPkZap5ape13LeCkG/g5/7ZSxU9Pl5+nFO3t+akL7O6s1Bl7gQN0wpQCGL29RWS3
PLX+Zmq75mgX8NgEkrNscaR2izPEJ0Td1w4vAhu0eGgncPbAvVjco7OwC8XIqgZI
JXws0T+xDjz1HGPjoTqg/UGgBCcEZ5kfKzEGgxFKnO2ZvogD6RidLdlbFSW4cyUp
Pgps2BvQ17Es1jvZn0zFaCzXVdR/HXy2uNyTEy32U0tmaSE0P2oNg4CTW/nNcmip
1G7sSU1yQbS5AfKZkAMEXxxDhzSmErk9BRefnmL7D+hNKLWOoLqibo29tIAthKMA
k96MPZ+m51uxAGJzm4j0qhpixCuQG5uZ3tohwCYVLVJ5lq43NnpI+8MxhzMCbzzW
6C8xGpRhMlBgu8VeAILY6DUTMR14+aBWzzmkMSlhH14QJvwNjnaernaMReEWkn2X
zHVQazt0pTdQpHD/hOKvjkZ0Cmy6mcb53Ntf5mGVTlUBW7hnOsKT9AFV8hn6co0D
KRiKdGUcK0kPxbLt6S1FKdI0hlAAdTGobtgsdeFRmfY63cMtDS+pxNyyzIU1jPqK
ccz5BEcyCGsAKHvsUcREDXEsWbtgVqDtvJ+Qoht0ar6ASxkMt5OtrcfAhWO919NU
81u8IY1EaUh0Bp2aouToPwH+3qF0u+dqDcsbLegfQRKMoCM50wAEMKI3vzLyoHfC
RqL0WWWoz19Wbi4vbJvTj4LAZwqduo+G0WPzsYPMrXGRoVEz8nPG1esYLrzmVleQ
yus6jvt2FP+3TzY9w7e7pTCc2onWNAhGbqsj4aFIEm+fwo6j01OjCiJzEjBQANbT
JPo4F2bXibbmSHQZpRjsA/sc/s0gEXxlufy4jOVB3X1/yuuRHsqw+6rGYrz1y9+4
C8cIFeB5jKCkU4LrSvjH+Ao8lutqhWkR9f4gOdRccty3Z6qzaDoIt9QPNVLhFEh9
LWWDHv1kFcV7QZDokdvvDb02HKd5+iLL9AwBZd0dm3RYplvZJsrwEm2gJBLZStqa
DPZ+kp21u9mpj0FEDkKO8RaEIr6ZREcB9R8JcitvAbhMhSZVYnd9ONcNTN3uTd6d
2UlEikigUlOzUK5WBdlJbNpCf/+G3nJy+PijSvBEdvZCPQBviqI3Tm/Q06r8z7TC
KO2oeY7LxfbvC69XRlpzHdcTomLALMkgLTp+6M9/4fEUBrELKJluDEEf91ICrGA+
jPDs/2qfFhk0fvWIZEiO8hn/kECZcel1QNvgffhwelCeG44UPI+rCjT91KAayEtQ
mUj1tnRGdOA4gIh6AQi6x4iAAhwOs9zifQPKJyIR9lF18XfVvqsMQwKelUUWYqH2
6tVdlisXEkeXPEYRY66xScJQx25qW2gMuRJ11d5t1sbBJkmJr902PFmik1oTrP2y
y/JGMr/JyuP+Ui7KuEl/UHnxvhdRL01GXJyOpZD/++D4L2aio/SMngkRSw6hNrzd
ANI9CY/SoJEVz1bM9Cv98hdxYujchI75TzUgDp8N/OtWw2Xc0g91qKxz1eFP29Ja
aeV1ckwmKKr5I/sdqRCo3GbL/OaJnCgiu6J12w1QG1FIT2RKPia8ulwJ9zx6U79D
z85oxSg82oeeRHcjes5EDh5olkzLGRWvKmoaUsPosYmEeeoigP3RO4B5FkPUwdU9
9K5wRY3QWKlvdsTHumSgH4FzcVSTdmuQ6BuP2Ze8Zt0ojWmw8YBH5+Yrq3L+99Tt
gXqEkZONRA+niIQpXM0r61wdzXPlANM5pndNERW9tWVjVjjgPPiimwIMgq4SQqZy
yFKQyUQ15M2+7cTO0F4CTqiWDtmrBMRqVLBgSwsVNn631PE92bciLm2nxZP1GuUf
+HY8MOZ+iq4lfuzcR6yLAroJqSqDSmUGZX4EJ6vnYAAqDwe+Jpbo6xjtsrHeobJV
2EJMiAmJn1SCHW6I2MFtCwZezhKCXgDSL5pnF9HDMIAUup2PohVLoCw0Mp3Y+gc6
9L+P6gehIPw8V2AFO3d0VHb5c90EDlxbL8OMOZEhY9HcFqDO6BZQXIB+EEQ2b6t3
Kid2qZkhFFlDqeMXqrFDcn5QsxdIi6aSTmHYKz8ZZ+E2smQa/ioEOw8VP0ivF5Ji
ghlKTafnliz3zS+PA8bANMLQ2JFYJRttRmvuWCTfG4DdXoffMINKYwQbnuFR05/v
YdXQp5HDHAn74JxBOPH7HjqxoLDBOJnEgEeJzF3GdYedTVeYrGrNu43gKDk2070H
7cfaFAgXdicBz0TsfratbykFBEZA5DsZzrpfmLS0nyWKD/6c+VoiJI3MIsOKihhr
eLt7ob/rMIowxKRivJCgStxZ1q/gGDd4D9cVhNwBrAVVVQuUTYXSHTW4ELKAkMuS
bko5TtMyvM/NOzJ/sZ7vEvugCT2xK5u9g7wRL+BCiBI8Aysnfyqyk5qsIZhaCIS8
uAcckmegX9WVTdlGf6C1/US18OVDxKpjVqE+5gI4GJdHczoY9UtSZICeOqGZ7Vfi
cEpMWuU50WaepNquOzyyil+UUSQMd5Xke4jX5+WZMFFI5XuiwZi9931wqhGbIe0B
D1l9d0XSMwxUG86uRyHvur7WubLy6t2OfFVuh6NeaFVeWR/rCbvWnPl8tUDZRiTu
6/W2ANlNHtFp8WWT96DjSch+LuDevI+t0K3v5QBjR11lTRYhZxOhp7PktA7dhPM0
P1B55oYSK3usgoONDICBoYVsGjp5+INCzUNpT/x+e2CuSkLvBr9cxbE5LUuv+oMm
Rnh1a6pV3Brvg9b5lANdbue/U/9HoWcraphdUBduY3d7pYPzqDmYkQaWugPsv4hy
taOHcLSEXy0xaDf/AZwOsr+2W77DEf5rE1z8948v3A+cf+l1OrJ0vKhq6zEugyNg
fJc7qylY+rkP1HqODFrMxMMOdS5Rc4mItKYF6FD2Kz2x7X10IpHas6N1NjPt9zwe
MjMERNfmt4M54xZ0rZgEUhJ+wcm43apu+Hdpo71Yebq20Kmpg658KFNibYx4ZRDf
9g7slJwQrjVP6XeZhcOQhFbbIbhcVlg0sUqHyNU/vpL6jBbNiPNt0tSW568CsOKo
j+dYJazyEzzFsY+qatz0x9xgublyEjcAXeOfttOiYtaPeLn7wpZMZ9PQzSR7ZX1g
uAoSlI43oDDR8rOb52/GaBxKpSA2A1RgXl0V++/vq1xvFIzA8rUGvDdabjbNvaeA
/KhGP2cI7ScYmVz9MT9fle33kSe+oSHqPXcLIfuf9oiDzBa3snI6nAMXimg3umip
qVCTWUAAatsX87wWYCmolQ331qhbk+ksL1dZIusVrR0/+ZRlOZJbzMulJeSILQ98
ABVjXORggJ3DGoJ6NU+hS6xBLw3waH/8IYzc/1jZRwv180FF8pReOniSxgbbFmH8
+/9jU5opeMtIw9eDVra+7+GgDcBK7Od2A1lyuJJuPG40EwKvQM+86xBcMfiB3ZID
SN3P4093GXbHsn6QHhQwUP3yVEU2YgOMIC525sTk4/Y40m6FbFOueStgjKvFsDBY
AVcSWrHiTP3MtlXG1X6F8izKH4ToSyTx+sVH6BqYkG1+NMitm0P6rElCA0qXJV3u
OWAbWnK8RtTO1oyntbm47cVwKZ3bLDOTDT7+u4/cYpviF+nvuzczM4URlNf4ykOE
iTs9TNNNqwW/C+kZDDKykSZh6vN7i3Lpw50rGvuSOOiCYdm8asM7JGaAk7KDpwEC
2OHkC5rd+GDptdC+73rpyfHz+DDNKzkLw+r/E3mqchcqBnbYAahBGnyJ1IyIyPnN
q0hvt+ENZaGgzdjoBT6Jq5gLEtyiKCVv6K6pmidxK6oig+pdUQ2aBuDBQA61Wh3Z
5N6MOCkjwxsSCQudDuFT/+xevMosc0n/2moZNV56xsGPfsZmXribbC6LQgYyAGkm
dESRSybCuph8giwkw4sl29qc+51+uvJkMJYf/AAeVwYDL0WTwvaeLHNngDqnTMSn
sibh8HP0jPpDi77755ThTmtxRR1vGL+3xJEFQMgKof5k332c/oXaOGkayvvt7F75
/FFkm8+Sh96u7FGMeAHheZ3UuCyQiELRxzAspcxhVm+OgSMPzVtGT9ogcMwZvmlh
pU5k4EjoxS+7sL/QTve52KtnaWjX5ZGeDLC443ye8glfBMC0EtX9HI+UnG3D6j3u
V/fETJtD6/nCtX6n9TNd5B85C6iOnXz6IdZK9+RZRf2uZjmgGj++6KmS93qSctO8
HyxqXZ712/0Ekhv7bEz6Wyvxs/DI4BTs19WJ4Tyuf5VIQ1I04W/OujiZmy9oF64M
Z7IfjqEP/XAPhTgzSHAC525CAimq0aGrpf5ulWGscRZYskg9OaynTUKrIITSaWVK
4LFZ9pGM5qD3wT+XECJWPz55pxcOwLqmZ0YZuKYpN8iryUJGZR9H83PhmNso5g5q
awCreKbfIQPysYWx4iFQFFPBJTMvyjFLQFAB9tKR3kWlx3UIcb5onoLbmDJAc83y
VdnwKlkXfRYMz4+eg50s0yr65ISs8VcwcLYQ5cpp3WvmjEr+MZHaqCZLvT78nFXV
ZNOex4h8x4tIB2njcviq15pa+vZUaa9UrvmaRWEhycgjbQZkrY9oRNW77giW5H3F
MgcHKWekuMhlqxVetP6zWvqcuuf9kl7tS2QXN4jU8G2IXWNsyDid85xWpXegC/j4
1qQ3KynGWxrcUZI2T+mHvIHY22rZ2wW0TDY7tTl8yy4/fya6U8Iy3QvV3o7S1DsO
EXA5YFDNuD58cKdIRp9VXnGkwuN1Wuq8feZjgr8H0P9iuWdQQEMXYObHGnNHUk/C
mnXv3J1cY06pLdd/EVshoOOo+Gp829rW92EE2jZaaKdNPXIa5FwT57oa7HzMidz+
GuCwEtUEWTST0TBFTL0ONUuQOlwGtph2/8LAjk8llAH6X+VMWVRQAoaaYZF+/5fb
9eizXxpsA1bRS4Yx7PrC0Ogn5B+YMpvQgPyq+lnZEoTfUsi8INj8AxSb9Zp5BEWE
HPq/a8tuCVv6I4VOPQ/T12Ql2AHj/k7F4wm0rIZDqjUjPxYNmLHphlbljcPvD/Hs
xCODG4Q3I/NCVuzouquSjvr7Ox/VAUd4maeerbHIDVMHBa6DHSydmv1fvYf8Ru7g
atjRf3OcLEJHl8xFUXxyOgzfYrN6NQv4u/HkYChjakRD0x/MFZGbwKZ+NT+gUbeu
jePBxN6EQqflMcriR0NyW/UjdI1FekRel8lRzHI7+HMN+BY5wAfsmymofCczCZOX
mVT7zMSpa/aIRN30F0q6isXW9gDuJmUmuReoi4RrYFoOOH1Mv1fsg/1DAMzUBsHN
cV41Ydmtxmmakvg+n8ZJI+O+bjCxP/Z3Zi9VcC5yQ0sg9IL77Vmmz31bFwq7R/wV
scmrdnoOa32g4GDA/2sAPuo0fSOLfyURzgArQe+uUOHrpLagT/pwGTReiZbHQqh0
zpvNTUEaKPTg4AqcFDnPTjrFKjQqjVLKRbSS1TyZf/oegbPbnlYhexL4Cv8evgnE
hdRW1Iqy1YHNi7MXusP5M72ZuXVDiOxe0uF3EVZCOchudCtluI9YB810tIJ4sDk+
MqosPyn73c2KbWMxa6dC4vQzwlqHvou49Jx4Iu3UxM2v0hCGB6yJOThbU6f5FaZR
Co/n9hrRlbb662iUnSc4frGFNUjnVkUaNnCOCvJxk/wF5OPDTGNPqFBG2MIjVwm4
zSRYwQJOPcFIsRmerwwpyoX+3E0SaQ/xgU/vwe82ODcxfhGLv5F0eLpKKWgUYUkg
mXvCy+LOv2uQY9b0rbJVOoS33QwVpkXMuFsIcExEFKrQTiXUofe52yug9O+SyGgy
opKAr9xu3tXo9zXJYEAwL18w3nylIY3sNZODhCY2YAtPn+U278h/sleqsh+JuV4q
+AkrlZyfwQtopbr/huW0yD1AIXKB7izg0+TeCYCfY/vzNb735wCCjSzg1B64oaU+
h/eRCUWm9PbRYxaasSYqOY44vdcd+VB/id3D2ToN6mO+09m+TZU6i6j5ouxQUsFH
y/VZ21lU3fYegfmZUmazufQpYmgWr/Y38f3Gnpb5kN/Fd/LKxmoGme1nROIVTxdw
0nJ+eRfBBq0LKxl0Nx+NY80YZsTrtwtWIrirpBcmSgcJWflLcvzphiVwQ3QBeNl8
p+CBgIJoXzy74BOr/STfzctH4ylUbuw8gdB8qzJk8bvVIQpaVKuEk22PtMoMMYz1
XJPPb5GWvmzh2AmavI/tsn3dxHd7KQihCEyevjWoLJq6ExbKKqFqXWOvvF2N0mfO
AuqC/6L9+kx4+FDnFaeqkQ1BaYv12ktdxFkzODn32unfO2ibcSmheOglbhQULn8T
fxEIuFnquR/IrW/h3X1MGS8Ih5fhgJK8+eOi03+r6hLZwlhI07yg/ourIn+kMBSg
wo8iKCs73UjKPh14xBtljwoBbWqAZx1+lxk08xa3kDj5z4gFmzdL0GyV0HQZ2LXG
DLEpsgBxDAU/ka5D3/ehaPSLEU/P/WmD5wAn65JLWfTiD5M8SnypVAgfYftXpXh/
Xt/AW5mTmii1RgTA/XDhjQyIYjstwpzXEiLJbmiKJ4kefI1aZFV9UgcXPtdfBnN5
2Ksu8IePONXRsUIEITOutlOVj3KwCq4TdwRpSRwB1YHqmbsrtCQAJrTOEgAPrUlY
wefR7MgQopAiWfGy+bxonYIH9gM9sO9cabDjBjB7U74U4uexXetHTjYHu5mFswXh
GgQtLLLRELYH2YgQ6w4mHc0PzNLTzdpTvfr/I/fLUN0LA74ihe7SXW0O5GSbnXQU
rR0yx14gJSgQMkLY132Foh+7jXoa/fyzknGyZQn7rZPf8JUMj3ZSR587pCJNfnSY
3xA9ufsgkAEvK0GYMHB/SEBN7F8+nqxk67CBzBdpfS6hqj85DfOQe8XZftI4HOJB
IlRT0tbxehTUjN8TuulCP6q8t/0uliU+wxGGoHQektUSk9FIlqnpY+XtKfHXi5oG
KxaDJeu3TjsTYLTCsZZOG5GRLXJav6M9u/iZgW5+fvSdLhUwT78B1sL295m8F51n
vXO/6dYcTTnzKFXXBWzt08CYoER7ZrOykqBNtUrDeE3k1iniVH9P+tWRUW3ccVWp
A+KHrNAt+hgVYiAgOdY3i6Li5wF2et7VLo+/CiYHwj1lw5qgFBBsNVACPtZgvuFZ
Th1UgTGx4hlmNyHgy1wCQbfjfGG7mz2Azo8yoySdm4Gk6I+9KMpDHohfFTAKJyA4
OdH09XMXcYr9DYcWZoPFVV2WJsmEVIIAdYvvsmpMxR37glGuMjUoj7GOnkXFWPrY
QuVsn5L4FE1Y3v63bf3pZHeMmI2qTcVFs3eh/wPnOXAB/zE0Qs1pY8S2qVh4MjRY
5VOirk04bfI3uqgp5DHkILmfL6w51HDasF2ZMHvgF+uipL8PJ/AlEobTu5Z9FYL7
R8BBqyptRMHRfaE5uqoK2KaY4OqGTal402Y7T+4oYS8cMySxAPKKTw0Lk+xRAwtN
vJZWqqWreBwUXsV7QG3CjSQY+gLWiXemNAJP+QghzmvdAOVE/NFw/qvURzSYA38t
2b9Gc2TqUKdglpPN/mMalpgXB58RqiaaEQk9I6gX18q482iOFzBcs1aylashCYlk
NwWvIS6K89H2tn3PVLKKNb1b35x4fbyxsLUA1B+EyFnZY3l0a7HnsT8GY1wyKGNo
LSXHG9DXpnM7/Rnk7jA3bONa/6pIMUjQ/ZrhwngORmLfEXBLnQrPega7/kChJLrM
aFcIiX4yXflQDJzYadXv2OctnQaGe4t9Q067ZSB/Trpucx4iHf07x6DnyiwpcOrs
USIUZ9Ic2morhspPwp+Wa4QF1N8iq//+qAaVUKpmLIwDgyxz07cO+P3+BavQao75
/nIGKD/x0qUmBEU2oQuLqMtYggy3AyUQ+C/zPZdWse6Swh7gfVBnmjbU4tMdeGhU
BcFJkdcHiFg5JVZFcOWk1i4RAygzY0KXmXQn2xVPnojqiO/FJ2WdkDRY3GII3PFZ
sirFZOh1v7eB6zokSJ1M9Ti7dn9JURE+ENPNF4Uakkh7I0axENkZFSEqbrfALzNz
4gzgoIo4vqaa0LUF0/AMnOQS6nAZTPot9w5KSAtME5C5bO29QXiqd7rjsTdkYeKn
R0h8oqoqGzjdzhTu29R9dM9HB9AbHBJXMzdYwGSY6weR7a66tUFcT6JTzmwQOKdT
EJFEnLPU2mR91RNtbmYP1JiEygk4XcuyWCD2+xgxZJIlrCzVES7F7Sflmby7ZERH
yaU1xtV7W7kfVOlIm0vRDVGX3+V7glW3MWyzfZShfkLkFMoWf3tB4TwpLQF44QT9
6vn9/UnObb7MlUvQPg3WEQu/PzTChXv+D+oDAN5ECc0ceqxpSJl6WPaUkoQ32pY6
h1+9kSfXR0eKRphHGWy3c0PemBUUUn6K4iHaY8p3INnciuoOwBL4WpG9UmFqc7Yd
966EhtVMX0syKxT1O4SHKjeIuB6B41f6UhkO8lRcLQU6DOQnMACoT9UfzLWJPKXy
V4cQe5N9Ls7QAwJSrwUIcIqz4J/JkJt7rnkpVwKmKLg46ELVZwr85a1EyLnE8vqI
jdYK2gfIbmeqqibSAR5ibDzsFO8G0HauWnHLrIoD/Az5U29JWtEltTBFX/93ivZT
1qWB48W9LleBPoRrw3kj1tFF/cSYkazU/tnwSlbPHM09UXwUsEN63unlFD3+ObA6
X9N/9YEaLbEXg7b5t5+B0zvSGXE6U6Ep50QkF8X4UUUGi5rZ2eP2rFln4+pMhfo3
WFWzYS7cUZSMN9EvLXx6mCiXbpsbQkzD/kTbyNnwlsCPyia3lBjTVPjpTwzK9w/0
MJ8mN9OevtiaclJv1D5AlVhxhMMujBZeNA9TGGO9VW9C5p7eUo6vREvIUEjpvEr4
1tZr50xh7uXOZ3wYt1LUntjCGD6Wpm4NIVQHecfpC5Rtu+DVASCeiuJ7pMGaJE/f
wV3H0OnLw6gKTDajqXH8iNRzjURo04aeruuXhFF7uRSoLXUWA/l5IUKxyBTAMX3E
+6z8DEATn8cXXE2uJixtfXcAqwTRt1zhiKIK6AdCnz6UpBoZKEl3ttkJAOoQfIeS
184aVRfR53tNVVAJuF73rlB1rKQOOZYfvQKGBPHdRvY7z9SNNiUloTLyX1F9AGSK
CkGgPupLAoIKJowvGlVCszQ7It/HQlZ1t3J4KfoBf8x3RNQ/tfeL9rmge3bRYb5q
i6Kc9n3+4CZZcdeRemyuhxxadds3b5aMvbQQqPiD93VYVKZrRklkkNkPAQm9nClF
4byq8n7eY+wctfYUI/DbR00jgEXTjyeIO0xCEbnZMozrXTcb9uMmpgjJ8ZeHfjJT
EjYz+N8qGACdS1qR5jL1vuJSbhe/1NSlAhLbKimkDVvLSGM+/Qd6pqMnFlHNX5Jt
zYI/GfrM1BjSi+ecL6CRUeMQC3mTgGQ5xiRyO1Q0KAU8Jamf07m5ZCY+9JFORPcA
fbxODBpIDqCn73xfaeIrjPO6QOJK7iRnFtnfuWsnnNJWMiTMsx5xb99EodclO7vI
z4MMrDl9z2upF+vWBy+IY8FPwDrmLrZcVV9Yx1UTfHsfunKVUqjd2e0TvBLo67iv
H6IkkDyevIGArc/lcyb1sRnfqTW2pVtnfXXAgty/iRWJOcyLDIZBPd0nKDVcKVHs
nKaD8GwbcvTVzJWJQefCJQOHF/50WhH37P3rvBQVfDVZ9yKxKRRw6v1q/rm3kX1z
XdGCGPA5qWLVEWdrJI5kKbrDQf5zxG1csp+VnONL8HHqag8oGxZRm8vyfbNZaaVx
GvuaO+WAfdn2kkyFNLzTSNtegpCDby3ImiVWCjaVuXdjyx/zY110PMYRGm3kw1p4
pJUP33agAuTC6BHYDJCYkUNgSHX3A6tpseC5R7sGyHoxevdhK4OCKyYAUugHchpy
kqFS6t9lb43mA+ksafUUhzhIsJI/x875e9GbhDqGxNHupQ7fK/38nsHJzAQkxrP3
wZNc1Qpvmv3qTcYuKbx+ZGBst92hX7n6+/Hq6ZvodZpiA67FDOROtN2dzJv/FF7I
/pK0qrYnIyYLKELdsja8dX0O0+M5R1PMs7c5wYNXBMHAqOIUJ9Ze1R3Tr5oaHrzD
RJKvEMIofMuc1uvYrNlr52fv8RQbQqfUPlfs94lzy9hHPu672mvqtpAiE6spQvPv
GHdh2FzBVvUuU2S1Wzk7V8zGQDs8G7DAyfqKP6aWOfODDjEk8ln0VTdTT3W2EQgR
Y0hpdE8alMkN9eLnyPGgaNYw7sEl/SSYdYJb8XvPzUbXeHw0H2nVrOApf2TL/AjN
CbaLIM+AVlUEAl/bDuA4lI6foQK0QpNWgoP+1YG/5mRlfgGnLnjJNZZ9LfoIch9A
NMIitfMNSS3tYZYxOKF+5up3cLBEBXShJI7DwM1jHIIziYqH57wIU+gRlhUgo5U5
ilCZhadIvyVOh0BoEgOv+leZRovzvfSPf5lkQ0CuD2U6EnAwvj9xClc2yIoHPk2f
S6IOyQCt6ZuibJVZCsW1tzRrmknLFXsU6Wcwot9FkKbDxguliNMizWNTJeEpw9K5
JILMrofsZXtnzcX28rdVgozFgqOFIqtsijW0UWyCEMtkL75tI5v1giEIN4oHy6nY
oUIPkxs+u+fVqRSqFo19EdZvNpl++VhBwkB0xRmMbsl/ikZUaQihUfNGGmm7iik+
2X0ccx3Yj25FtCCzwIzIkg/BFBEOX5CcgC2ZWGgJHztUWYKrnQOrh4kPUsGE4axq
RY/gVHFs7B5aEIyJzlgNPh+3M4I7b/kDt3zQu6gbwglKbdVfHEWfeqKihBYcMURA
0WjeA+X+57ctcAWm5+VV6itXjZgEZ59igi4uZSQPcgPO7A+ekFh4EDIh4Cz7jeoy
nzIDLyqjTWicMrbAxMgUO3HiTeRkp5aLJrytqKO26u5PdkXc4PfSu8ZPUr6VMHWi
gSbZqUaBDPxkjWz14uq0bVJ2d3/lh8aQBm/jSk/vrDdwBXhrgZygw+tZJ2zxh9Gw
0qD0WRSw32zbrFKJ9xHlrsn1l7CTfDzdpM1gg9qT26r0mC875aqRVXlSARDkUhCn
8gKzaAQYstAwnSCyN7j1Df8rEthJFF5HyeVnc0aCOMT7MTOEIBN3I2E+JYN7y4NH
HbwhFRVacMY8zGAeZJhQOVYHJti8fKrDMXb4eCECQr9cLowQJiF509EChdrHwuBY
kqJh99FF/z+z7AKFJ5jOoRh0ak00puGUHGLnc6nt/uk1vXXAdY0gIbQuSzSRfCyE
BSu79LXIIHiWtY+j7GuCRAaQ83c0kP5o8cHrIo0APBWBCN8rfL76yfkYV4yS0JYR
xP1TH2IrnHJEF8XFyZf2MqDl3zoPfZQjL0hW29Lus4sp+TZ9uZFklDhE/xSY9ouD
6306WDQaIgMNQ1qTSJTsf72qC0xslZz5xprFXeqrXj+ImMXbx5x0ssBv25K+3ICs
G9Lbc4IphFVvQwsf748oDKQvmltmRtUspK7tLxSaXjQqWK6qo+vEelyByE6M60RQ
Mn3Y0TfCH5J9WiZLiTYhsPtgSLj8qwYqmAhowGFdZIfQxhiAcaDEyL5w8TLLME5+
cyEJzHsHQZXM0MmVDja07iK/ELl1MJdawMjVz4cxE8vNVgmjDv3iiAd/yRm0jUhg
+0awkLg02VmHW1pBaERqpuMgY5xxdQ7DUHrWTwzUFNWY67jNvVjlXbiB5ciMpI0+
aoUZ+F34qI1nkwoUbROi6NkPWrBPoOt/B5Gl2zPyVB7EUQQiz/jjK71JT4kNnrI7
GtwqsazoVDoIcLydyi7GRvIoEQAzpZjIsTQCZOwj3UXNcgDNvu1t5NQORdgurElA
mFoyn03RHi82A43JPY9DGSv0LplAW0M/piPTxJqi/Mz5/9id9dU3gIvW/3IWpfOF
HLy9iBNnM8VaYwmAPr8Cq9BSJR6a3G80P9u4Y9KXpj2xa9ZGsBsMg1xf3vzMfJeE
5aqgS+7ZG8bYJ8Eg2xF1MxjCTG/X6lIaIunl5/o+U08aeqz1o90JG/nr0oYiNJ9r
DmR4+F1VhSIVvFPM9zLC5MJ9Jx2N2/cZz1l3mgs/s/qxDY5RKgUNv5XW8tDsoNaB
rXCYxF4b2p4gpUjEDcP0ICNAVjpNiBCVnpjqadOyuRus+UEA4VKLR5PYH/Wq5QaG
lJZ/bmLmkNhpHqsWGEaV+v/wjgqxHgIoEmeo4QzUu8G5aIvfVZ3bOoPKxUbnBF14
gKR50pVU2j0mcYRS65QBZvqZ42E3vuYsQI/tHhVcvR2WGUfWDw0iw0m1zKsOEG+R
KRoSxCijCU0H94XwHeteERAadZy2rjDOJtf/y/gYsDUqARQO59Pitfkodj8B5POU
maOh5iCOngMClfgArZ5LE2ainM0V7CwjQuwNb1ygH16KUaRULmFXMFkau0LqoOvx
Ts+Vngm8/Gpo+4LCf/0nLJx5QkxhUiZy0For/oy5ay7lVQNua0ytB9A+L3+8v/Iv
uD7dd/pQXqvBcqt4O4fIEKCG/mLbnbq+URHZjBpL6K0huGQ6CWNbnBO0tbL0g1sh
qnq7OAdXftdAGLf1/9as0Gzq8kR5RC/dhs3fflUwKO99WMZAG98yOql5BeNcqdA0
fq9zmUkKNT6RnKoaWP/t1iCmsVvVMqFiDhqUYHkn+NcrufkVsKpECqfXIXDxO+2M
nYRbX/FmUAjgI9WqPOB51wlggsAKgviCg1YsEDOhe6DxliD8ktMjKdyGfiGOEhgJ
4YfqDSMFX1sa/v51w5a0fxt6RyquPxldnkDLuTGM0LGI2NsBd6vzbjmbhZELGF6i
6zVsUqQnVamV84tgvIyT62JyDSB4iFF9aFB9jxuEqzRwW1X0zzvKif0KyLhu2A8q
OfOmxf3oI1+r1U1rqQTUP1Hqz+AewBgrawuTl27qvBxJXvfSerOWM+Do43J0v4Kl
K+Dw4wgAhCBREOWJnzCPj30YtQyBQEr1hJswI3fgEA+uRvnhBfmyIuyhgOJ4UJjc
jNzIGeXIxCEIluN8ekCBQPT7gU6DqeQsxKG2f3JWK4I1hIns19FFA+FtDLArxuIG
rse6L70zh+dmIzCAbKc7rXgDrbNeaLz74MRMH1YTSy3QKM/lzP2ORJ7o+eqICcw5
8+9zCsd0VxQLG/mCVZOtZh6QFPYgq0PswTbxAJSFGkXohT4BtmyM9fPO28Rf3LR1
hz8GtldQW3Zy+fq/FDM6y7ZZ342d+FFxcjMFwacfHNSrHrh3q8Yd8ClRF4cEr99k
PCH6RykJWaqF7rLVQob6/9Iyq/2lHb/Hqqr6F81iSWGBo82SMM685LPdihVWMkj5
WoSm12YwZwyRyzHVh51lmdFpAAoWGDW8PMWWGn/z2eWF/ks2yXjLb3/A3031V3Ku
aoTkjy3DIAG08lMApLiZ1IuZCP87civmjIdWoUBg2tehwadhiesjOcZxcVOHsUpT
FwuhGOTp7SdEGbXFhzhB0dUOJNXQONMJwIwTNZhG64Rw9EL8bhS5XbPx99pm0mU7
Ni/2pmoRl16BOOs7sgM28jV6RZ8qp3FBGyBuNgw89YVhfUVqp8qi6l872pyJNNJh
n1X6b9h2vTmINUpjYzTn1FyAePbVKVA27vDdx3DRaAnTWClliD6V4e+2/wyOM728
lYxOaUevbdR3Euqm+HCyVTnj0qMuJWWDzJbYktbE/38y/UrHekd7mg803IZJ+vqU
rS++KaxdScgk+Xs7EDxcYnwtAtW6LfUJ+MoIr7+K5yG4u/kl6hxZI/fdBvePJcOv
wPmElCK/9jwQMbCAJEDsSp+Dqh/oU+xVPxqPgCpWWrn27gm8VTNpLEEto1UMrQgI
958IB0Sim/vR7ZGqbeUkwZsdSZqP/h4qecExxHTTS2yqzxOy1oLnUTVniaTugW9I
/skh2AQSLGl5nj0ODtdyTyHJwTL2bSX7BiVRmiwP3xYfIyvklpx2F3H2YiCslIhw
yYQMHdtctRPnaszTqaAOUQ5855bQ3IABlpJ2hHgDj94XJIv+f1Uu4f0tYtw4QVi0
OyXaKGkw7bxmRtZEepZIB7FOE7KbLLVzuD+gamXxjqg/f0tBBane9hSgh6dTY6o1
/E1ntjVRimfiCN5pI4BVByb4IxZyJbDC6dKk5tHf7aWiEbyXvmMHHJmSZhEjRKOK
LGvdsfHKbHTyWdn4ZzPVnL4DD1oWsrcUbRs6qTeqHVwQQ4+NLu9j6pnE1WbFBwxh
z/bTT5Et2Vh/CuRTW9+YVYqdybEROM3nO9bLgUEKpKoV7yUyyIsaX5S2S1E/YA9t
lbfKkWW8Sc/YeIfB8y9yiZDd6ExdKEUCMczBqoKBZZzs0XiKrrhzw5KZa9x5tqUl
o8G5YbARwJurnanipnz/W4vGGd7z2B5Uf/Oc7hNskNcrGksX3p5Kl738M56b1dIy
nCDgLLQj2SJ7dRrEAoWa2R7zpA7iagt2TLONBXJ4PDVJzDkHdLuK8zm5m25ZDnA+
dRbsaP5xoRVbljUWmoC8MMw5Ee/Hfx2eskrj1KJREMtvIYIOdgGAPKZCnTjh86Bg
ZBy+Rr6WfKqL8emUqz2Z7ICoDyA7KFlR49uZE5/MEfr0fa/6bbo0zeEgCaI+/lmt
cOkQa5uGanZJ4fTR01AncXJnmtvdjSZsUgKTSXP7PN5FYbLwPN74S0DACzXF4weN
MfZllWVP7w/0STEDrd48pKY+ZOJLka7vWrX35JywK735AgykecB0yfsZSyMADllJ
Qar7oA3mQl4tqSe2lk/y/cUthX82nr+UmrbzJySGsW4MVPFuXOrzumtCOljZ0zHE
Y5UGjLIwnQu0JB3GhFVgGO0PUnSQ/C13Wjj4PcwvfexL1Xvli7sX+/enB0nJQUY2
XYzOrywr89HWHsD4R/Y5RumiHcxMhmEoTXJFXo9hBRv/2O61zqdCnkuRcIUbpARA
f5GwH1ZntdBgtRARAmADJDYHCn7vKA36eWc9iB+TNQBxfbFsHOvAxt0gduO56N4x
YL/TBO3DdHo7pImPal0hr0CdG8g7Klsxn1NCfrneBkAghbDYQnNjUTQcCqzMc41t
Ldk5lm2d20sPaT0o1dZQuSsn7uJJLy6QigXqxijppRGvgvuvcMABiLrr8ft+i5d3
A1ZVIZTvd3LbzUHLHdQ0lxiwQJqB4jRJY+K86pxIzFq8ekAr26Uy7893uIMnasN/
v8vObx5L+mGHDxbtsEnLIwaOugu/aqyReOcePCGn36uZSpSxBhhFTzcmvoLUJsMQ
Vh/xs1NyIt43D3sYmwbgOOkO2JpBEQy0jMxZbaQhuIzwxpquAPdMVb+l5kmmGnpT
GDz0HoTt0bpL2rApSTgGpFxDtAbsIReiEn7xBDxhz5KWAod0jWZWxCToFYo5RKSF
/FYKU0GTK6DXpDZEXovIScL8FghOAHA3NVy/HBNy9yCoeEaC8sWQErETZQZHKpWN
MIMT2f4XCpS2I9a1Sh/wF3S1Dk0JCwsl7rqyp69xre/XlVHKwdOM1hoW2bR8bjJW
/xhHD+GoShGsFegYjBgj92ZcFHvkeZbJuiXXtV8wrnuwlOcpnzn2ZYY4e9wyUqRy
cOdRhlmInswIU8wOW6T9Xq5l7joOYL6pMNO+I9JkXqV5zgXM0eCwUbWPTv1BDgKl
7RbwCxairxbkC+xmDFhtduwf+gE10ob6Z5ULiOB3AO0pPr9QHew32jGAj5gzKPPk
186EiZU47/k8IXnxyM3vrh7NWq+Oo6OLw5+ImtI5+S1XmKXGTffOBCHxvu8GlOB3
P0apnCOFlmVHjRvXgNAIXSAfGWJ2GL23wf58313M8NpaqSKr/hqQcm+HQ/ZNlvkW
YO0T+m02O2WVOWAmuVZgmevySkYQGNuTivCTODa4bBpUgbAo6na68uqiSc6EASb6
xX4jhcnSJHW3ChKwp5lEslF5OycOQeNVAHpih+zcN2ZFLnBpVVLWnaxrjkW4L8jg
jNUvX/qPt9fzWsylWU3udMV0DKnSxZGcydaO2j7pbgCw8Na8CV3ZIrsNjYeyeThb
8bUPqxMuT2hB6KcKamTnRl3sqZ3xIyV3cPFSWh7eqonHUoCSC4AxEFPyrPg6zEcH
PVSkMCU+jaReaZ6e5+yeJBMXTXcmu8mfO8AfvZ0QIEyWv52NvhY69MSkZI/80ECh
ZsY5EtOBARx1p4luxR85+Y8mwztewnd3GzcCDffspGcyxz4fPSX85lfFxp+T3yxI
hg8liBcZulODTYHQGMyZqtZhCzgje+YQkhTU8wcNvt8VRi/DNOJDIQqwkrDkHSRf
MuzH3WJlhfjAZujkYmWzfjYB/+ALbgtKzT3xApmNVqSe2QnWI6l6bY7s5dTNFYqo
/xf2uYmxvdNx+IYpZGpO6bc/iNgwiI5SbQBvVJGzjzVNN6+DNWyO+4ojWD2xizCq
d50srqFErxXjCO9In/GHWfs1ucQQO/3U3Wt/OQSUbYCR9m+ntDyPT9NSfZcAwHaS
A06YMp1QCK67rzUHWWc19OK4ljMDTriw+D8KsxkRVzDPAHRZh3OeUxW6CEOklqZK
tv01FJyqd18O2jIZU5sCwC+DmuUl7UnNtxncJjioiNk8RsJ06HU+6F+2v2VMnybk
BcFoJmVmJWXipNrJkkImNrNKoW54FZG1nDAxJUhiYKnb1fOQuSEWXuinFgQacy1E
yAR0VZkprm+FH0nq+r1lQa82pVoM2wis/CLmJITxJ1GVLp4auZNeYDzaIB/Ms8dQ
3MbNFxdOrNzXCRDJcoES7rQcBshl5wjp5AgzvSj+XdSJTZrFVrnhKprRptGev4mJ
NIoYPlZ5zid+z0bVK7AzZSwBmNWWeB+ByAu+qAnVS0+hsPYbqIFlBKYnsIRTytoH
fbZOZ1qiZ4PkseksrRSgJv9NP8Xehqo0qG92LXdrGbCinLiVjbeD4wsFTyoZlgZl
ABheWNvY2aNcnMg4PIasjpzjfQDjkhUXAzdzUUZQjEyjixwuWr1/Xuzy/88uQccz
8vVapObxQr2MGimGqI0EOK23btwyTw/ib5IQSaPhpRorRBsR9D9giO8V7RFjZ3vi
GmeIsn4Mw0BUu6ATg6Isx/+xn2bdey8h5udduRip6OiSKxYQ6kiDsmB5fZJX4QHm
M7t6VyXNkXlHZaOqP3HPgDDrSkulay7vSieFfoth3Mv43LREEH2hmaG5mQaS8i2h
ln5uNt5vmWYHHlZvMdXqWSjJKYKKB8eoUCUeHED7yF+ubNTi44fJTse4yXYBD1Xp
8xmqpdAlMTEsiLkT8slUu2WCzHAjWjScUJINZ5Q6N9dpoGBWE2YV50Xmzby/outF
HOSd49Cbb6yahcsHyUyxmDqcJw8/V3TOTX2TMo7TCYDM6ePVRdfQ1vwY9ySHcaej
0Mt6wArtXhuKCPwJBIRQCXz7LGY531HFJht7AwkpYPeBqdQn4QKWdT+CC+dFmmQm
2yuhVdHDaHBSQk5zwo0Q0Jjd6ROiGNlRNOdCM6a9l65690rdKklVl8YUieqSzNZA
/d8fOBszmBpKjasPhWSIE6PVcv1tMdlIj2Rj1ZAuFkpk+lEzqOPTEhZOWeyQ72S1
fETzq0X9w0iDqwXeZfdEl0P2neIYl6eLpev9ebP9aKMWNht9M2bNgV/tNhpe6SUD
VjWQ8s7NLhv0o5Q2Yz4pLaKS1Mm9e8/oROE4cbuF7z4N31bYiRloWpbIkZln2JqU
UfsDjr1u6U77a/goAsbhlPN4+aamec7n/yt7s8ENF1MbLWr2C0tPeS0q23vMEfEu
UWrzx3Di5OZt4T5frLKo1FuEcDnAlOwPceljauTCilxb2zHuGQ0P5h5ap7mkgEQs
kQCJqvUpvqBkV5IUHgYZ4VAVAX7/uLr1fYd0gkF/rXvOfGFEsSQkibK5Q0ORKLIt
QP2fIzpBuRZys/8kbuze2ZdQ0gsdjh0TU/z5jkE8xIzY6qrbAbGVa3/q0q1d+sBK
kY3QB1ukBIuej+Qa71dn4kHX1NagI4W/x5fBYoKcz9RYieoUiiIrLbEPyYEsK5eW
UTHy2hoZMyvvegkfC+zwu8Rqy9X63tilDzYwPYfPBoBZnV7ulyewbgRlgNtJHs71
L99SDJZKecV8pkYU2QhLrbG/oKm/fxwbSPG96L2XdA6Ths0yfeE/hAKM6UZYFSnK
VUNqU5s2pEZuTNwi4YM4/YH3vCaSTS8iZ6trjTQpy69OY/FhjSgC3TmgqGGeeZgI
uYHzt5AAmrMKjuNK35hVaxDBnFpODRiV0q/m1QrQMcsPWJUgL4fnPvO3kMHIzUJe
MAVXw/HO5Uu8rLhRgjuqE6HRT3vMRdRUr5KmogdoPcn6Sxk0PujA//kFqj3XbAQ+
37AWGeyRbpEFZHgPhdDI42M1qqH+tU8g2SZwNAueL8WqObJ6zDjd90q0tNu19c+/
Lr29EMXLirJA1ufEcp+27CnsK7P61zn/UbCpyNLXW/y/i7VqnxX1ZgXYGHDsZu7Z
Khg95QwCIvTyotD/AU6CKR3B+Is/d8avgFTXal2GKh+ES8JlqJJYgh412sDclc8/
t80xSml7LoyWsjX6Ygmw9kta/NMN/jhnzOCuXT4VfM+JVwmQsqL3VEMT2eklpZOq
iYQpF0tK2tCK9J36XLY1B5NL6jMExJIMyXUpSC446AG3Uq5BoKWkMWbMqjNFZxtu
CRGq/oH9diymjjyVuaCSAfDQL+EtSYUNoMBe+C8zcBwVwtFNal0ULV69DtIX+Ap0
MrASiTxCWCckdQyJT2pGP0mX8JfS1apBXw1oo0ACsKxLPu2+MHQfnm1/FYtcKozs
bmBVU+GTlCqtvc1rPY4cuafk9PcebFVhZc7NiXG0cfDU+YpuQoX3mom9s8NKwVSs
mOgNKxD6521Cr348UnBBSmfwXLeiEqlW7pH4uJRG7fDQwfHWEz9Coa9vYJgRrAeJ
nmAs7syLwrQyyjWgpViGmm1pX8AJjrdlND9IEJKAbeOMDzG0+wKM0tdtLdCmM2Q1
ToHttrj+HBREIySiSv5m8B5PIeJe76ysq2OW8mRJrHXIhvVjDinxF2zOEEs7vOsu
DzT8Kz06g5WAtC2RKo3QDUmRUaoH0u6VqYuOjqgjhCPYLfxOnuePSyKoDRobUmWL
7zcL+goNWH7vQWThdTFgHZlSOWmL8MKfmMCYGQRmOWeI85jKPCNgMtPGfUAFaBLU
PNROD/8pZZcSvn4yYllCdMH3oCQ0UA+oarS9VP6gtE7IobGOPuU/adKEqeBat04o
XFrAHsM7Un2b0fbDrqTWKyPuP+92LyPFnFMtA3Qt73o/ZAQ61KcpT8GYz/PSbLFr
PtbLvyA6SAj+8M3xnaZXLPLKdqb7KqRFEZGI4PNH5y9yo2jIvTA6XzH18qqqw6TI
IddvN1VG+78twRk2wwNb5EuAyWI/y4d63MrgQ2a4x4ctLt4BFseE2NA74MXB4qlx
rJ+UYK6f7T5HrrkO1Y9P1nRSIh5oEwyu5wcJ59ViWBJpvmzOfQ5e/YhiAmyjbyjx
WF8bovIF/iBMKAbQa6unJPwa6X+NFWhhVefoHs5yZqe3VWMrGdsaNdrDERHZY/dC
+7P+A1bNwtNFYamqFKwuGM97qew4Hb23Wi8UlEdogh1GNA+ae9JIKKW0pwNGAd67
+Y40HpMFz4tWswOwHwUZCyjKF5jSo8xsNPHwjDw7Kg84XAg42+ayTzSZrhDzJmw6
qw9+EViL8/Y38i+3KkOIedbaCW0kMYRaW5noX7heMgUvCjjRn0qcdjWn/lZ9ohHQ
4NPaUxpCH3mWs/kXw6TenN1uW4G3oyq54G/ib24zXst9jKG72Dan44XNBoSUxRqO
Caiw3Cmk4l0N7bKbOBXHh+7rq7Xlf/MtL7oWhF6Pwk4aT5qP2VWKrDoalFBnRdVK
zxgXBmN6DCOaQlHsTq5rW02y6K71sfu5GmMl1yrOP45Xqy0v0Hv5TektOslng9Uf
YqHWvz1U1S8LKlOSsDpKlCd2fuUwJXovdUz2PQnRpLROMIPCj9ABe9QpJGCUcSf/
I2GkvQrOIP3FRt5XuupShUg5gTRcdDgLOfH2fgAvpYwG/Eze7cA5g166FJJxQ3Kn
/JKxyKqHX6uqplHPt9fmitLKZuRtqnWWheyRx+iOsokdZ5H/9aToASmCRmJgYhir
lU3J53qjuM72mZ2ip8ilPTpBYtruQ3dJfhTkJHqHQBxial4LDNCIEfaCWfClSlEW
wTRf/4td7KteMm+z8f8m3lC8u7fvJjwu6n3bkRQ1GdrJWgB4khpYKREUAtH+VzKZ
d/WfGw9h4zvAq89lmZGMMliIwPBoH5SJ+CUqqg8m1obh38FEcOh04dtcJevKiWfK
EvDya+fHZKjO4J30/4HXpd/16xyCJLk95csn3FkyCQ2IQ15o7HWZ7msPVQ1DG4aZ
EueCJfsIfkBOq39f6a7Y3QinCfPSuaYn9muMBb6zNmTkDV4FkVgErfhZIYYYfjjD
BjL+aJK6tcA08WkfXP8Ieh2AyV3f0i/jgtpEqAIOb7NpUL7opnomL3OjTEO3RpFF
5GcKCIrfCRt5hbMejFb6UnDe8E3Ksh4sn4l51GItF7Aq7WYG1tvPH9hXcrqFY4Iu
v71S0rmaia9gLzJHQ1Oa3ycu+G4/1x+G/ADryVZfqtySEuFZ1OfgEhZQI60uCog1
/xQFlIHQDrqKCUKp/+jxW7Etnd92cXGOsrhwgM4Fs22Ih9e09p2rGZ1CCdZ0k2k0
sA0CSLdrGWhsm4Unu3SN2/qgX0luHJdvqfncD6BSsvR1PuU5TAlsLoWPUXqB/+oq
ugocATavsyPHlr04Ve3ImPVwe1Zs3Hy6EakmFtXrvLnQkA/ps6TNfxDjxgUcYBBO
niqroqgkP8xL5e2JJM07Ny9wWf9pb11/502gpAJ1TxYeVoTELRXaV+pNGbtxf1lj
lXDPZMxr4T95aoIiLyD+4heNofK8USMZKVE5KFaogF9EGzXoNh+gAt3CRWeM4+YH
2MYhPCXmvNvJFkXGaqPmQg4lm7X4rWgu1TfKRaNRS6aV4seD8H8zvLY+HjyR0XGj
WUJl169l5PvOIGKikHYLvDiy/5EJzh1mwHvhbvrcBVSiOXuWEbWmRSS4gIla0/y3
XNd7HSP9JVSwKEZBoBNWSQxGnTM3KYZUazKZp4DcbcwJ/VlS249N+qUrp6ltb7J5
aimQCi/z+4gU+Md1bnZ7KchZc2Ut8OWilB7nDmCQ0Vsrk8mpDxx7TWEicMFyq8X2
hI8r/GLmU3HYAH26qsgUcjRH9xLRBtvmuUT3W+IZBVjssXrRpPiLfcrJsyjovPr2
KVNGAxO0RXbJ0Pft1MksHHCaErFqPmOe47ceSgjqKKYeZyo6mE28ja7GBk+YeOs6
a6NPgh4rik/1ASXvC4JWRClx6Ji0soAE0R48xb7wlIoVPtkv+XRx2H4lsoSAUM41
O0cUF9dYYOQojfpeQ26A3J28iZxS8NYp7HFPAcrq9BjdA+CSa+CxTA6qLZ8+SdU4
RNXWp885rY4WxoSenwXgwXEg79SMRwxieyv+e0+AFTTPW9s3m1YHI4M/InRwihee
2v2h0ipWYDXvevK2xDcZHxlUeGbMBCz2yVCV+pmwv1h7Osc9poPTd7jt6ztGvGDh
vWC4j7ZvZmPIO6pGmUpjLIl/sHE/21gjQw4xnjDCjJx+p9Gv+EmjXYByT2HHxdhQ
0cTqQNTUoObPacCwwgNTITyX5z29/njHN6o95RNO6KaYFbkN/MbGB9uaB2aoLNWj
7RJ9VK7XpGsZ9q2XtPiQIJ6oAKD/bszZeJ36QuUJ3KlIpa47rk9x3rFN+PF53PW5
sbJHawpobXG3trHiTRJ8hFRmXsyT17BFMJjYkLGi1i2/lxnPZDNHdWjAoPMMBwvV
d/t/7ZCmYkRmNtt7OPxHrKRWTQ1QcIcjxjHmVg0dfHW3n3CNfqWeDpglPi1KiX8L
4nkOgpwV9Dtz1vWe/qWU/+2JWhPGHt66WgP8Nf93BpKTd1LJRFB+5mryyUUL3C7Q
NIq2WaBbiCi4ipJqllw4Px3iNMYcPMBz42+8uqfA5b8uLdyn0tjnSHF9srhdQmil
CUZixUQkkrIkNj5QUZQg0Nxv1eIaYYPht8TFkINauk2eNLa3X+1DkhtuDAcQZUBl
xLoKQLD76f+K95/Ra5AO2fKdknf1FatddMEl3aTv596Sho6SeRLG4m2pdjy2LqPH
oaQzx9R5hhbpHFTq0zKZm+8kIshHvbjaUCxWQ7LSr+BF4i4dIWli2moZfJ5olmai
o0rhAvMgLglT26cESLRKnTu1E+otXD468Vm+/sHnp7K56kNLuD7MFNW+PPB/833n
T+rozFqGgnHm8TZkCLtE4wNHdhp/Ip6BEP4WeHL1GEyt4Otiaa81YsDuRsyNSQgE
v/35ujxM2+OrAKEtB1bD6YhPMWeuIwGXZSCFxqCBzql09vaLX6J+Ax05AVKlr4VL
4HVlhiIx/JaSp3Act9ZouVatzDb4ui7Csd26jXEOmcTdk4z+ZII3iLtwGfot47T2
YlMvc9G++PAi5R6gks11wgiF38wV9OtA1nPR+HVtmuXh/t+Z8cahp+LzkWHnnbJD
k/Rs2E9rr68s0LdDs/9aUrhkWYVCSbD/5PuLv08TQG5O8Oo7XimTuKPBi9zTcc5B
AXbhoa7kgo131a56QmMV+gYUhq0NRavD1opqZn2NHnf4LSmxDCuBz1H9V5INAYaG
xJ9JKTwuYkGz455lmFw9cnFBWtjgMwOmwzFSZ8qGESQtLKRcPVx+Q7muItXfMfSJ
OpbWQZFTepHriLjKDfncB4Vq4LEqJ+a3ZPn21lnKNkPAZEAdauQzBK9jiqn5t/+p
Uc2j/OJYLxkVwS+y9kI7r9J2nV2frgxayh7Vi1m0an/TvHcXP+v7TkKe64NVawnf
uxrhcIZNtDbZ+RxVuqz+WbJ0xYfVTZmpzQGvI58M+ePty/lQcx0Wk3sqlhBhrt/8
vBtQvJOrayfxoMJcnkhYIm9QeSu1509C3j45pJ9n0vxzZ7+s6CZSHvZXRBI9tTCH
dEwaOG6qQ+5nOhX1sTJg/bD7kumedxSREmT+4lb7TSFzuqNEWg26sAXh3pfOW5CI
4rrOtGU1zapzvRYZjRTadVrJ61cs35eBKtdyWL8yEBq7tnaRia1oQHt3vmdAzNM4
tDaYvFiN9vq2AKRX7d3OyeD4RCdLUYVtsQVTUlnzx5b8dXQu0FqSB9clfbwb5Y7z
HUdtSSUsqKIXsdd2MgK8ONsEOuhqq7fSmnV7sy86GNX63+qt1HxsXm0HfcfAGwx5
2lUZFiG7w7Gt0wT0AQ0HxrHyObKfeTO5qU7vZJkjFs7YqPTp+PuCiAnct/UUekH8
1QfoSydj86abZx362NL6WUHcGx3KlhIMahDSqUK4RiCSiOwDDXhTalLr8QRoPSqk
UU2ALcqotqdgMpIjKxMF+/eeAK1mnv2DRATddPuk5hFkHv7rLqD+3G9G0Cj/52iH
PcjSRuNeZQWmfkMgpdt4hmaxKJNhwKN1gR4L/k8Pg6sVvcPWLKq2bImpKdcutXYE
HZg5tEpae2rA3TKz6sNf13HIhqOLgNGHTPigxMgVrMeDdzpk4ki41f3HsF4MMWVV
jvRorA6bCHKMXSoFWEj5K4mEfdW8jMvJQ1V3AsO3l8sIU8RCgHuCjWwo7eGl0f0v
/TRYNcgXlu0EUEiUxyI91/swauAyOAscaNMCg1jU3J6c9/xZiLuEsybcF4TccYRb
sfopq+7FBKKrOeitfT4e/FWxUK5foW1KmwHNMaquqMNNSs75Kyvx3U35rr406FQo
liVsdc/hmxXXXoGs3F2JaFARLxVPz/ewyzo6kSWKMp74HcBHvpcPsPopXj4ZCze+
b1ssbHdXg3/jnqYhpJHkKONDdj/hII4tMqrtJHVd2guhnjgCqeIjISV5BrPeb93w
sbEH/XDdE61YS6owQ2b5Iy5NzANAM+T5daprTWDq3ukIVCdgjWMepzz/Gg07Hzy4
cFrfoORRwBbhrhhf0dueeEuqwyMDWuSZd+GdcURDGj4KR8B0xiDVP1MauIly1XmX
JAVATihhFrgk/a1F5yOukQR54kpIzsvf73xL5Db4UOwV7scBsRKaK6ChGKtngVwt
+25p2qxzRTApeWsYcyhBvJd4o7ohSKNalL6UPWmXsTloPXCQmEwvPhxqbGPSlAuK
kBEOqM/27/zImMPOAarMOUW3gQk2jOTxdeFhi4lkyjXwubP6bA6xFV5Hzhp3FEc1
ArFzwyeZM9nIQ1AEcg++PuDc3U8deCJ1r9Fxigq9gJSvigjIef63Lh2+jF/DaUjW
JkusDaKsrcLr6F223oEg867w2BcX05vD37oq8/VRiVz6XIDupPw4zfbdzqWkS+9i
gNLj1ecnoayaRStC66oPBMQYjhvd0FHTrkNstLPJ88T9Xl4dxtrAf1IZWGHZ6i/Z
nSlFejMGJq2+/8+pNcXBtFA9KqJaXT3qum+JFYBSdl202aYrTFOYySh7KuVjnRIl
VPhWimXHXF7XoGLrqBjbxTfyRGa1yUP9E8tOYS1Br32AYIubWa8AyC97mWbUrY9b
QGJIIruqZLbt0IDxT19XVw6GZ46PDRZ186gp8M+Cin8QXRjeZhmDIb42AqeU2dCC
1KhYGH6sXtkHv4XR0DnysVYWy3JTpbpTRVHoTLRNcyd2jRX3b0o5mPtxeWJ1IqOi
Lvi/fvokuaRsuFUMJjH4pxDWRJmJji3GwMIoxc6GYwzn0iXTUIVtcJ5izLGyGIpN
ZBuQ5eRCMygwv0okp+J9zziCrJJeMrFkAuVWGVw7aZ5jdV/quEFhDZEMaGBnDXZY
F9G5sv/nvyTOZs6jGELRQc1jrTcB8EJolb+/T+TeTb/UZI1B/aqCwQ50a2i1Guxs
u0g4LhUGCi2EsvaA8nVDRwRvD1hrz7mMkMNFC1zWhpQsRD3iwk0zTt4ka2voSzDL
nkPj3G6eEGL/wvFS5smUAj1XhhFUgw+vxk4Gc64Sa3dPIdAhmgn7YRsRn/TARpTw
DBqFwI5sAhJX1j9mWFPDVkqEq7JT1Jww4yTuu+rjNIaZDnUf+PJMNCGb6u//eGCj
l8YovXOHXb5GDhRMMYuf1BtxVBg5rzUJE1c2ZIKx2G+cw6m56qGJXcpTbIc7tcqg
VLwLrMUOMSUPa/TWH+AyFTEf0r/fr1x2RUOsulRwkYkxM9seD6I0weBB6F0qlgyB
MhO76CRP/AGGBArsEzSgxIVAeMC/ryTR+ssBCufuCarbGWV9dNUbQLN9FnInknlF
zyGJ6h080Dn4Ox8WwMLI1l7lN80h3TYTG8phFw/+LW6M0O4IAq9fubvKqXcFLCtk
Lmr2NjiOrinJxXf7x2MaxZT/BpuImu9Cn8ICI/Lw4r1zstmKIp9yuVt21HCTOlvA
v+9m/HasSNUaFeclHzfLYRafPuctlT0espfpFRpz6iM5fXM9TNZGpCUQNIXtSbs4
bl36d0cJOxxj3Id5TdTNLDoMaZfS20pA85cpXPtkzI1bLVr1Z6HPPGgjpHPbntuR
xBVpnP9/ukHypFf1ynZeYh8f9IkmsvSBmazj/Ruwl3iw7iKCh6kGPC8d2nJCQw13
pNfjLrMm96+zYt6FWE8mNsY/swZEW96hd6xSaM9cNZA/jm0KdEJ0Lu7BnZxb8Jdq
CH74InJeYoC2h6+l4J0i9gvBva7pl2vLPnb3naVTD9VS6WtLLWR8GEQ9PJpigOt3
45SRrpqXA6GxMjHIN5YpdUslmhStQ9VXy4+y6aO3HZwfQy2Z/HK917PMq8Wn8un2
JyJvJnlV/1VvO6JwcHrEn2EtpVg/QbdKYLtWLdYCGrpv2AMlvatsk0x123Fd4TrF
5a9miJnhPd1hFU6UNomJ8hRQPG7Fb8ohkno71+ncbmRa6xRKxb+SWhidNvLgPsPI
WPd1mBRTkrRuy/6TbuUkXmEVABU2pMbIIEVeM3s7C6ZXPhGnwlXz2LYzpnY5nCK+
s5j2RMWDEyvscbp45QZog9Hk9Mttrg1ult67mig+lNy2aUESgCHQaQ0sljVqAynq
aKEPK2DlIe3RZ4pWnOwQKxOZX5DFrw+s81dPEmMzki28ILaXCmN/Lpgu/2mJzIX7
43ZkpJ0/VAnJZ6eZuXceQFORoGDc0refQnClI6Z6JciFT6PAGVf2gPE7Ebv9oXgR
032iq7KheOUARhTDCxPu04dAyjXPMwXF0lbUWrGAN8lymwNIoR48V3Pi/kG2McwP
u5wdQJ3I40iyuRVSO4s1wnGOTmzkdHWXXy6wgTy4VGwA4Azblu/LdM4f+f8fDhx2
L9xmlCn5dtuHAg5Kdjrec2gu86mwa31D+CWRMsaGPiC4V34uIzC4NHcWLkbUiGhC
jx56OXBEfO7cSuMP9Urzzym3RThx4Eo+EjjrY1LlpObbZXpa2CFJhzTuVWNZa8iN
kb9UtSS/fStyGA+KE1aONg0QlSq7BVV0MaSUMwe6eSGslqj5H+EuCY7tlF80MANt
z2QM340yiXnGZPQL0SUoDcLgP8swjVDFRLuFX9CWVRgUHV1btBiNhB07J1RNYfwi
uY1eZVAw727cTQ7Wp0in/dDv/qH6Zoun3s46MvHEQrzxKgcG/LReZ8mjHg+F8xgf
A0ZlEDxJEZsOzC0RCs8EAbyIrCMB36f6SiM4LnZjVrqGzVHNEjQnsWa3rVqd5beH
fzlP4dFbZbMQszwLDr1JMAnlExiCr2QCe13fEiaL8N56rf/Q8pyGdH4SA5uvWKIU
Z244ISCRbERxHz3mHHjEE5El9OEcZtb3YKv/NqI5pwSvGtiLAugT3ztz/PVv08C6
kPCOVQfdNqLQNytiP3MZVp55dk9zl26o7BdjKyX+U8x+OCFqy+39tKe3gGS6Oqli
HktDr+zZs6msReGWeLA11Qpfgyw5Tm+IEGayjJt47c96htN48lP/4Or8ihnB+v2M
r43oBTqTpwnYja7SS19NKIkTTZGjRVd65fz2BQtqpRw/HbKXoU+eO5cMEweou0tv
J+OMMIsTDznOqxuoKMjNFHns2S2fndywge8QFDJ7vxs5aS+Cp64hnoCl8Rrqe2hF
LpGHg5laQW3V+ttJmCM+XhP/KSveiZiR7x32w4P7UhLCHwYnF+L683I2SX8xP1os
H6/N8ppbGCyySmBq3bU33LYsEt7+0+QfL8lTTPLbwAO4UtP0Aj+ATHoxsaG4luzg
+d+gzxQ8kKVjBqYMAAZ0OzHMkjK3uCLo7G2w3tM+FCKEHPYu+wQ/VgnXUvnh6XGt
h0a3uDo/uRZcPPqtytsYlN4HJ8TDi3MlTRy5+W9eNfwkgwoqz7393k2qV9vL2aYQ
f7S2f5mqThyOeTAC00k5m0R6alKgikZ0O2Ia8ZCXNtP3VkSJg/RV+bQ6micpFq6+
gPDufzMCicvjW8xK0CvN19koepmD0G4xGiQ60ohcASoDRN7LALvonwfRKCtBdPie
+cAqJqy2229wvUIVlmCvx9Kex/Pe3aH4HNz4740P0HWcrP/7QvZlePeLbQaMt5HT
1Gj0dMzjkVBe0xOa4vydawLbX3VC0l1anFuoFP6Wb9AgCGeAbiLXwZeYFEtPdC+L
JDGkxeUlvIIQlaHQB5a4uDd4DYyrA/BHCeflIUKBlAPaE7yv3UQ0s6jIGNRg4Nl2
B+rhlrgcZCHWpkX/d/ngS0RPDAzWd3v3T0t/0/fFc7XTnFHVBY542SgB/888ISTf
TwaZZ1dsE5nDhOpFz+YeWgQjgGMKPJ/zWoneORlYx1jBCBPSLk2X+XA21Byst2b4
Rk95MwGN/zlbCJnJdMszjxTC1zAEithKCweuh8bzwsRGar46sTby/t9strJRRdPs
jNX8z8Zt1C4JYPji4Fpkv0qTfQbh21kR9PWJWb7zq4NrRnkOECaP/93aqX4aubkL
oTFj99GY21dgvObbKjOYchzh+H1g9heRHNkfl4sGXkQ2cXCnWuTgPGzd/jJJloAg
rBRPIm+I/9AI1YDfrvaJAAPWEuS3YfpGakpn2jBIwYAqSedvSjcSPriF8b7OGkAN
R588AD/2AnDCyx9OQ0l36T5UZV7yvfsKAKjd5v/B4vIRKQWThin/qLEBDVpD4wdb
kgmxaK+03n0wBqMMFbXtXYDxZZDAyn+viL10w4hlKeVFGjigHG+hwKnjruw5BXKX
VeTSE9tlsnSeUk1JIyPwLCgiFuDsQLYG1HmVFWrrRRrYPMaYCLJUpprQ6dwehsSl
C4J2AH00Nd8DkiT5hqkdH7xbIwbSjGIaNIS/6zVtnRMfvepX7EozsDHUjiOVo53P
nkOF7EeIVb6z9W/lTjtIqkuWNC/U9jvg6CWgkpKLIFvq5NxnWtqozYLfzCGHtDCD
67rleeXfl1eiBy5Ih0K53/Yeo7uu/Tu8xn8lwASxotk62LHKVSy2E7Zy/P57gOSt
nKdBG9jTxahqImAr+l3/shYsu95TmjW2gNYLRoxO4V+CDzNSDFrgzTKdo5/rkavf
q2K5CBcCzxq5Pcrj/YDSqz8GcLjCHi+FGNnFWZFQsXXGiXX3xpOA+Liibu68eEu/
DiD3oB2x0psNIW5D66F3k2+YwjOMvJN+Ze0XxA+Ei5NzR9XS97EblmzXeqHngFJQ
qaPj1BEEjfPGy5Omk6ZSizMCxYcOGbu8b9ydfCAjvkoogv0TKoJVqnxM7PAF2+nf
rUYZr20BV/niH7JbtdOhfo9+oIoIXQ89b4NkiPJFtLwZ3lsKipj9I+/wbVHNgLpy
wUpJGYMmEbcQwVJxBRmwNl64kbW/i6rYErARShMV7GNCfwMRZeqlD2j13gNu+qEn
3b3sC6eHkZ+j+k6s3xMwbE7AR4Vwm/0MeBypr5oOFXCLs4u4gV0BXLjJ7pVqwGGH
rJH0ExYZpyHwMVY6hFdkqBY5PXhEUFyPRhYGT/BNaGinMJzyW/OTRla0kbju2Xrb
O84j0J7PNuL/Zd8iE1J4rK39+/gvSOMt5k0Avg6/N+m48f03T5THt0Xk0fxMMEqI
/Sa7O25ypmWogH3N0p5oD4FZwJh/ZcQELk1ME+/dU8y+wEFt+xFdvDxuZaa5TxP8
6anjLLCIxHBQznpLo8Eon6vDdmBXrHVTOKXCWzoc6HOoscm+uElyfXdiFzebUuEZ
Pjaab+0BrU4YYCEXT+cswj9e0/ya0/m/2qaxGBxyV+RXMTjlXo+Fy6v0ZcGeq8O6
mF/FhRlUir+9T/RGkxpNS9EAsq2/+jpvpgD54WwQ+5RQLQnW3lNnF3aqtH9xNb3L
habSoATlRRoEOKSGemLx1BLJwnsTu3TyhREL8z864GQW7JM51fuTqf2Ykn/kEm7G
WMAvgtzadGjBURK1kTCl/8FTZXcaZ4VvnZkKJyRk8r4ab5dB01TzVaOzJV6LCNG2
cZ60l9yWnyd2HkAbRzcNCM2v3TlgmMup255J90Xt61fq3EK+AvMQyYGTXfNRc+8B
29uMgw3T8qLVu2+jC5tx7WGZWD74ZLIB2PxTfq9qUjq5Gnv6R81p1B79VNPpgPgF
j5VURbQm9Tve1JHh77+cfCF54eAZz+Sc2GA3rYEFxBmxY6dF+HxJfeYkiQTg7FD0
c7xzOgkG+O/zXdYE5Kh7107aCJsYpNRecFsCoZqZf9u813Q1qvls6HZenJyJJAvm
xRX98nJChUdb5UQDE+h2tNIpbT3ccKXZDDJxFJyGp5RfOesTNU0EvHzpGzyjejIg
wQC42ZfZ8bE9gw577rblsCLjLPrmfvD1h1N/v0FrhNyqWX6Q8WC4TehBFx6/ZwxY
MblpZCLp/iA3J0RswGHFEnsHW3k6Hw/bpGg/Y22KpTCKFL/Kf4QBBgsT4uKQ+6CJ
tQttSy+YkJ1dwDjjT/lNY4Q0A6Y88ULkL2PXvTYVPd5kfboc14oslm8EWI9bOgt2
hP8xUhcV34myp8iQ3YXe72JMQtPmf3j/3UIOqVuOYebIE6pTrluOIGCB+NrVUz+X
WUTVqY7sG1GAJIoNB80nHXV2vvj8XQO1E+2vgBFIzYaQOpPFjvaqAnqMKP4z4zAy
j1yx0mhaC+Ra53KY3VZDfU5J9LmrdGbwGR600wnJoCh4ggse+iQLa4vh7OvhiWsS
vYiZHrYYruI5Zc+sctziEie2KESfoQCK78mXJwesgSGW+I657CbtbjHYy6tsJaCr
JlQEKBpBkUrwuYd7k8FLuJ/YWLzsUVryu9GcP27cFN94hDGg1lopgXvtfXd06p0Y
4EgjTvHl9msC7msxbBbw11Ont9e1iQUNMvkg+tQusjWmA9iiJsSE0OhfaAFQRRz/
QU+eKxj/Rz9T77UfStjymmK26sLYK+YRxh9WShsIDjhHuEmWhBZAg+GUEBlu/Gc+
xVNXJzz/2izB/b6OerMpIM7FFSNpXaTHX04+SWbaIFMkiaStWfAPtWAcPVa7oktb
lz4xP4PMbFJ12Yr+oQ06cyRn6MTbBgOi3awVGkCwE7MHya8P8KaDP87V/L8BKx/k
QaywYpiQJrsASRS3AmRiK2khDphLdeItvpxP1+tuN/G/ZrF+8YNqrOpyK/yXHVuY
jGGBxonRXWIHrOHeYSETe2Hk2t+aU7SA/sRzWJVE+QKrvVxIAvkGRbNUPd41hz2n
jD1164CXmcGNX0AylXDOVt0Snl3B3kDl/V7WDgWem9kBjnsluNdw+y9oAr2QV1+H
rE8gz8pzbE2pxcOtNNGGOCk5tx5Taje+Y5/EFYpKA/xnEj2rAovVF16ItBzEj3V5
BFiamzEEClC9H/LhLT1shZBXMZBqc3mb2gV60RT7tzvaQacydvg0+dkKuL5Wrb5i
d/92NNxShPc74qEHNsrR6fauuKOwZqNRQw0olPzGQ23w8/tfEJL0cmfQrjK61aV9
D8Bna/Dwku3PL3GWBgsGe6zUo3pnkaQfYETDOHlvMmyVkoqoAv8TxZEmuijT1f55
uq+8bLXQgRSUOeHOcIyzh1RQ/9QOINiUpmEIADZm9jajcqIcnR+ZYireC5fo5QlC
RHfmv2rcIEnuW9yl/hpFmgPOUtpU2wJTtd1ZwTZyHwtJv6hY2Hz6II3Bs7nlKhhX
I8WDCG+i/wE7HpOJSxmXwFEe53jgKqC3m4BrcnR8ywcsbs3x4eqQC1iTIYdo7j6N
lqJ2pzCvCkY7Jtjl+wbMgAC4s1oqDCYOcfrI03AOlpCxh8Bj8a+pgWNSCN8O9I3d
1WFnJmNh7wn6of10g8Vlsxp5zyv7BET5QiaLGMsjm5i3DIC10f0P5GH+I7j77sUz
5JNTMsp5P8fkpgkpBPO7kxSXcepQQ72516c0sJO3WF9NzYehf+xidmtbm/yrtxge
tGv0AW7IoGwHiuStb7Z4lJ8Ztb9o2PnOtKmJmA08JaMsFHGgDBq8kh2pLl38eZ8n
f1GJ0+Krr9Uxe97d9RYektDqEsVMuwIAYMjj8KkvwNCtzylNHsuiMU2wskGvDtLO
+1Hzcbs3UMeU9LpFquWYYd8vdTTrt9YdTyJkSNVOy4IPD0L3O+JzqsystbUIZolW
GPihvmdVAzd26wRNmnVk8sON7Tf55sa15Dci8IWzLAQtykTF7AEO83EFWI/Y3FrZ
WYquC4sOQNGlb7QEFe19XtzM0LVKntxU+afgN7+JiBQiuU3RZR1f7R2CLhDJhL+W
B/1uOfRtth8t5fr6cLSKgNifXbEO7+8nJlxWevDsl5+L3qIyx1j64MQo6NnvGZE1
2ZnSath9JfYFOj8vzSbIuU2wU3w9GRnpXw0UyzyoW/lpQVUEAY+4z1ZnYnwIfm5t
pqe35WjaLbtaXWwjWMCxnLZNhHlAp6wamuaZ937DSFOxQjyiEYc909WHd2UtCeSv
Fp64uZygIQmTCavk0E8nEfwccJiK48725uN/4KMQEwNch0Rq+0EEHwS9dhG9tRKt
F47cN3L6hbjEAaQWZIptaYPayfzSfceodIl3GcWb4tNShtrrWIJ8V1Q0YzAfewmG
/yF3bYk5tUPxWywYYfbFxaaQzleiLu2CYF1OhylatpthYmvlmksbr0si7bvmpBEm
4TKoBTgoRCCYaACUIxaL7NPOG+EMIwFGIO4eAbOzrAVXIKKswQTNxFmtJe76+FW4
c4lXZShBqLMdlOnjHNFVeY80ryYWs8jq7f+q+E9c5rZax2k0eA8ceN8tgQnDx9to
2fXaKxD7SIiKiIAs9Cpn7HC/Qa0Le905iJMc8K2msHg6qlkk9m0ZcziIS/WVsEEv
tprQk1CorIHf62p+oIhOIdEtYfu2T/7fr2avUkByxHKTgi1TgUGaErnxXubdRhj6
q25LbagcTLZv14s4SPr0aFbFCW08TCWruY8p+aT758LVJdPAM8LsxrTrhtXFk/Ri
GEB0uW945KvhQ7GxvsADSaXEpf2eKEYvGNWvIFCEUkgcdtrSAL/U2q8x55Tcq9Q/
wFXgGqTUbIeoZ8a9SGv9WOBXuav1AMMW+eTH5J/Z5aTYhVWtkXzOZMcotmT4aOii
YqyhBD1Z67wYspcQxpJUTcIv/ofjxkCi0rYZp3OqOUuVlH8vRMDhKhZn0rwWFnoL
NfGL9Wq+TBrXLxGgD++ba8k8433eimjT+VO8TwSqqaxZ46xkNz2o39yf5I076L00
Bae5jVuV3arO5ldiGkiav12sHYQdiTv5+DI6cp3vvlWzWzU0K95PHgjQPfvQOKAB
3G/AxFMHVQZq34Z00VJ9unx45kGpy2ytc3eWni0VDDMpbdU3i2dVVpFIdsALb+PM
Z+JoumcqKvkco04Ek3jUMosAoGyxoEenTkiwNB2qEAV+AQkrbEbP1CIgTjtbcq91
5Ys6M1WCj9qVchwdvS5BrerYMtiPoDhhJQMZ+ox1N4qP6TaikiQLuoUtgu7kXBc1
hlDOkooDyyYvvurihjFa5yFKShsWRC+X8KROrNYssxCDrDWSnx+IVghlVCIFrVW3
NVfXC2aFbbdigZsgWtWLpWbk/uh/Dyz24DW6MQb6IEfPZxeg7CEcLxNU89/peKqK
66lsjmuFzkRgSmFiEPBLS3uNMCQX3Qm5dMlvKwiXNrfuSkgtlt+isyxk/ZYsoWzy
G6H59NZVVpK954BpgMwBgpvr2hBvCVmzy13DOTJ4HpjjTD70oWozDHuTONFgRrIm
xZatbyienkbZ7SRiB5ZmR0Kiz5nn8ymMQ4EwLnWlXgq44tWMi6WXvmfXic8B2I6/
7PpG5u6sQClZP3tawG3UK50qDD7PiR1+6VdfpSntlwUzOzhAtDlcLKY6sq+P/WaY
f8SAkiUkx3CIb6Y5G3oMW1JUo3QSwupMUe8pd1zYvhC7mnAoYRcqCGr2Kp0oLvoF
HE32V/dgp4Ff3JpMpUyoRS/mEz3I/Sb19e+xtx1CrOWucZBbnK5Bkty+uo+mPN2f
eJ7792IQrYfsIbrdwie/H0jbJ43UOuaGwnp94Z+Kp/pFrv+aK+qSH9yj+KHIuL2Y
wL5D+p7jXTpLhDW+XEA2uUTdhcbonLRm93JS0xYb4MPREQtfEpueXSKCB8+pP8xT
6xFcZQEcLqMb2qbDvaBMpSxGGBbkq/h/0+F2HXbDs86PAJKLMNunHfl4VxjgYqH2
9m6Ld1miu3iMUvTGHoLncNVuIBhlfpgzP1Uc8dyACCrLL3ytUOpsvtc+yNZ3LxCz
45gguxq4380rnc8ZUYnnj02fUj8Yvf/xOfzLVvxI7DeAaEZLWD5LvBc5kmk2XrOj
29IXVNiwjribs4NeADhQsSyIh32cYO713/RWEjE3R92HGwwCQnCwMUK9K1SDeL90
45YLDexkSMDoDvuCNK68o4MejI0WvOEXrpDVroX945CjCOdoL2eBEEl0e0YEqmyU
xOx/5ox/jhEmc4NvZw6207asePXabxYtqqxGXWkpP5Zr4GrNNyOFYQE7UWBUH84v
FBxLmQhZWbTTINWDs1+cJedA2mywscOnzxgl0M0ikYyD4k2RJyxNpNMtlMWb+Pw4
VQ0wBOmHP+emRCFbjsrIOUVTHzclHQylg8qnKXaTCqh4UnjYQhsbLQ01xpU+CrH+
44BLLYpKS3yqXLHjQuGNoLSUyu43GRakWudSyQnGT4oukUKvTdmmQW2T6uxlN0/s
gVd5cKP3skXn4n7Blbv3Vv0+emSmAU8swV5QPYu2BXfHczEvuBkgln4eJDheEM/h
Q/HTpFVEdNX8ckV6PNLWHjUlyzomsbZraJ76AVnrrg9vVa5nfv3Ag8UqzZAdriRp
oZYHx32VN9CncWbvfwtr/e/E2nAhsDygntTPmwkgOJZsnFrX6zXamBf8Kc4v6f57
O1YfadlwBDrN6kiEqE7NGb8xiCkTcXzEzMZioZRxVnjy0CrjxJ2iHlWbuTWbncUp
m8eHQsUgIS2lbA1qGJTmKQ==
//pragma protect end_data_block
//pragma protect digest_block
bGtuPeU0+CCyrQsIayG2i5zu4ls=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2Wir3zjMF3160n2FT7gg/Pk4SI1E6RBLFOgaxWrGC5tulmQJYSZN6LOcSo3gOjtc
DLg5nAM/S2exP2ldpqEyuLGboiYoa9+DsRwRoKTo64ivVdgWuW7Kgil0GfIQOelK
tXWIcaza9XYcRASxyU5fsPItNm3+b6vKgYMQ3bX3iLnGsz6XnM0AUA==
//pragma protect end_key_block
//pragma protect digest_block
7+BHSXZvInGF93wonXUW8HZHXIA=
//pragma protect end_digest_block
//pragma protect data_block
BU0gvjbW9R7tn1Z5AFNBKSqFWfLWTzvX+5v0yUGJct6c0iUB4jz+3wfTIZUs5JcS
M0elH/Q6tlxhwUDR4NUc3ZxdGphIfmZK5hB4H3/WcBqqG2S/Ol2uMKNLp0bC2GWm
TK7PnjLeTEvLwVC/4ErGaJkoDXTzDbcZ/SD/ThCJHrWVwC2WkjV1gvc2t2V4SWSd
u+Eq6z45KLxJECHUpVp5botYvdnz5KVddw3Bs0rV8rS/FdpQE8U1MoTkJifTxKLl
a8Py3zieL5dF6Gg7txiEhCUKJrKdd2FpRIki0fvOb6Uz3Zve//MIImGBq0jevTZh
YK9NwW/Qfpb8nB85WfjyWaUy8LXAhX8iVPi8QH87GUrv5QQVsQ7gFE5Lf6tl6y6B
te6KU+wR3dRK1IQmdsKHf1uDrgeeNGAphOzycjz0cIFOWhrtunET7jb9aqxD34qN
qLJ/sgnrzu5aw39OB7Z4fD80F1kcgXYTQJaTgCUsBNamBxs4bT9WXeALM5fosX5m
IiCYwPRBxl4cj9A0RG8ax+8Mu6VHQAgTMPvjyAEHs/I+CM6cAHn9FIbG6oXqxMzH
7FA0XinwJDRRTxtF5IhOUg==
//pragma protect end_data_block
//pragma protect digest_block
/+LuzrfKS0PVu0GOeO1Ftehnzmo=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
LJ61AFmLakEq/w2TIP2hxy3jmHq+V5MvEn4hj1lz7bnUPHqRmgN3Rs+0bSuF+AZr
Ls/keOnEh0cxSLTbJX8L1I2G3pwi+IrvYpM6+FIznOxewvs0iNQwMC8WC0QZN79i
esCPdkbLB+nGik2nq3Wyvpwn51VoB3EjAnIMjNHoVWa/XwyOB6bieg==
//pragma protect end_key_block
//pragma protect digest_block
CtHG8zczTxtvoFaHU4Kh4t+eyu0=
//pragma protect end_digest_block
//pragma protect data_block
EGfCBq0YsRPa3fyibU7CsxKvQgazn5VxCw80IK/qG+Q1+pu2zzXXkEiPSXRYoLTN
R622yv/PW1JYkUmEkmg7mzgSxImfECWUWJR7kTuCd5J1BOvxHeMQVXao68g7oXF1
xG//BIN9G+ZVBvNXXLghqy50MxlvY/3O7qReHtZEHhZqEXLTPScYBGboXawwc22B
3qTkP36EEUOG/WvzHMD59VII6obmSeEwulaOU0Kw8iYkebcHxP7weqkJGYxhnu2e
cRcRtLH/C9D5YG78HnzZb/X8xWIOTWWgII6Jz0o3lxtVcrHugj9E3fDtwFBj07SD
VpEoQPygEGjzphkxkh9I+zK4Ex5pKNrWSPCB/1Mb5uwhoyU01SN6BvWdo4D8qDlm
+rkjUwf111NRS7Ph5PuIdhDTyVhshQ+IQ/GERG3IlyLqERHkpppMxcUYpLS+sLzt
x+NRZ+aImIjYuztR/AUMADhUbMfWw2RzNiFF5HPuz6/Gv6mpTadJt3raVwe1oi3i
zEjt/kfO72hT6FtEmN4j3gD+wi6IGy4pVaXJlow2Jj5HmUc8GIFDXK/AgaUZA4dX
i3hbGbU3hYFjEtJGa7QTGaD/YlI4oWqfztnmQ82Bi+0rSkA14Umcx6uwu26XGL9j
op580KT7dynZsTPrnNRc/Bt+m5KyZ2JMVVpeOSCkDnvOs64LSt0CsKhnpCcrzt3Y
QP1i5eXHBi/8tM7kAVXvT+fu4nH1snqHvGP+yHb4FGOqR7XVl/5DjfuCiLiSf86J
TZg5n6kHkxpc81tFgH3R8TgQ3kU16p1FkG+ZXnZwUL0oJiJBlWbsWMWvzN0vEm9V
Bl66u/qviBSOA/RJh0uaGGMJHgBus+jTYXQc/S+p0Uy2QqPaqbrC065Aj2KcPj+2
aOh0TguZEBSjBbrSE6rBNz3Sf9FPSN6Uvvebb9HKCvJdXvyqAfTRdNAidheAhtnE
ze7k+I0vDIHffF5SJqQDn5XeAyES7cI9jvwtrq4xMivHDLDhxVB3YCwy7hJLBm6Q
6L/1cfhOOnor3PC8Cm7JG0GK8Cye76JWjmrdqDH+PqoGyBdqmkvb/UPsbCwNnch/
IwbvQA4EO4vwihQdVJXRRvEXre+tA1bJFPaqQBdukfkaxC+2Elywbh2oE54A/ea9
PlZtWkQV4itKww+2AWw5hOO+amTXyf2quclFdOBokSVxrhxh9yI997mD8ccYO0Mn
R61EgQ0KO60aOw8335075F5dWGBp2/mN35kxIxDj/ZRBmR/evtyzfo26GrrdXjRD
VdldHyz5Km3+YnTm9sN1TeTx9G5qIv86ZDlY6RwuGLTPKWpnwprcucz4im5uUE8D
VxiOEKUz6GkV+ek6QU3LSl75mTqf3bwujet9sWmMT1qfXPWJcmBnrijZwsNCMGdv
/M9uoloOWoRAn33b1hPtkaRZ4y6I0HATawSn1NsvbqGcXMq7hTQbnbS4vZCJ5llg
vb3xvY7EO4RbEDmkEfEkAAkhIsITMyeeeGzvPnhOVop2O0/WgxU4qwoZS7K3OasT
dragWDW4UsDH5GSC0lr90HmpJEWnwKOxI2edGdxzNSobaUKRfstBoh1PqfKwdyOp
9Vgjget3wS3DT+hC7cHVgtkT6eQfIcHuSjHQe4nMjd8teYA/AHBnmsk8ElPRumSP
9uo1PP7BlQVcQoxYNgxjORFG++PumTw6w6iSti99zfdTHbR7nLLc7KizKcGzXZqr
Un4YjSCPQpb/EYkWBWLy/eSH+FEQoIDCTBYjnb5b/MdaeZepRVcEzdypSoruwWO9
PSS4OyYSEuDPR6rPWg6fpvCYW1dsRicAaFFC22nswJXdULkuDYd8KEY37ELqMa2t
3AGHk/FimCOSpeILKRRhCbW/iccqYmtEnXCRyAtPDAI80o42FpQKZB5+AL/WKjlj
5vh2EqdDMKR/G6pVEz6IuwylSRu/NBVRp15+6+X6gyB2g+ZZjj8ZKFWduJ1oBZE9
JzK8yy5u9PMeTrknH2CgilZ7oWZoB8zRsmsEdKpR9aymmZHEFZ7NACJkLk3eWgmC
CuUPyqkBYM7rHkoGHiVfgOL+C2DXrPrmnKvmIVFm3CvVV2prTM2AZsQA7xDydPzB
qxw5mX5YHLtokNiR89ztyZSCCFAH9ebAcNLgLXBIhnk2FkllQwyxT56BVHfePO79
GwmUpWwI6qiK7fylE+QX9DE3acApPBnUDBoCp9CeTV8VKKIKL74FX1Ls/Bq2GQbM
+0tGp0+jq+Op2COkpNt5Nnnq/igzUC8pvhapRtU4DAb30tU4UVfXtRcDJuOkLxSC
81QlStVixUQQnxHEXXK0KP2Kee/lxQVYX+rzNxg1fknbemLWTQdofeNdwkTnvAQ1
iV/smnyCsw2pb1TIUhLj1TQ0DbzdK6vgmrP6RLjrwOwQvpN7d1uZ/uVReIJi8bkk
1WJxnleQx1Nc3zVF+A8/VA0ZluAuDkkm7TtUAC885umVuZD7czStFYoRvRb1en4n
bO+8iPy7PbY8DJSZ1rGhm0P5Y/Xqz0NlbaHnGhJWLAgXOUDXU9PD6lSRiQvLDK0t
1WEKuBa4USeLIp6kYMEPl0J895mDkJdzuPOMh0Pbhh5ssjQJavwGHajajY47vma8
wE06Xuu2IYVn1GVY7qIgJ1STdsS2eipsl6gkmMsWL8nrhBvrCg5wHAI7zJQ5TJ3N
PFZKw4KLGAOcyxIOdZFVpNPH8hfRwHEw84k1QE3KAPjW4pGUamMqsVH4ovWRqmV+
KHhsaDS67Pg6H5ej3J1FWsRID102Mic1rInEcPTKZ3vPlszHZ8S8X4EPLaJzDMIZ
6lpNF6GEYXXnFQzK0csf+5pHJN+YSS5pZfZ5SR3zul+gljP1kuqHefLDKOTEqm6I
0SGJILEoh8BKmwd4k9PP0z3rtvfXzfzGwo+QoNBLuxmCsSv4l/K1wqJ5gfnT6i+1
ohFp0YOvz9bi0N3/75HF8bvEv7dDrzq84JussP/uGTpy8kG2HscxEiiJxxQ9Bsat
nMu1jrVsASPac6RgcWAI2E1/Z1F4MMWSNd4/8RTCNkuJm5Mc8odcGlx2jgPZUgL+
9ZbCM8lnZZTpbvks7dSOIlYpBXLSppHXuRNXy1t8QWYFSseRjaeDH8hZPoEZjx/p
a75Z9cLmJvD58ktBROwcBvJLplOrVERHNtn5momHkrGjITvdFOZI1DIW2gR3EOE4
9uxV0LETguc2dkOkT/iPTSF6/ND3cqYjIdZ384YteasJfJMgL63Jzrh/5sxM4SqD
PfaNueCa3k8ZnBcWAkbjdMEXhR/KSUmxbyVwq0YMUBDUBZNZF5U08Z2Zt5OkuYWv
EoVuHY0B80t2hYJd5HCrBOTk4rt+EH+pII4BepMdq75ai9nDgP7jZu5K+eM3y+EU
6tF5vYb127GI8p62ksSfO3FzLjqSHTeKyGqpulzv1wrCjv8qDZIvuF2zDdZUSP8f
cJsB3LH59L5hKtKLgx3GDKEz2386xsiBzp+f8pp+oZJ28jfV8kbU5Tj1Yej3AiY5
3Yce1tTiMs0bH6/UN68d7CfS7ipVgWyCjuOJtbNCRJmF9cNoDvPaFqQhIi3zEFKk
RfSPpTdvxA4fOYUCcHCJKS761Agge2swgxS1SOTrFU5rKtFmyYSBQsbddkkFjNSA
ggQX473nQnIvojrs2vVQYF82cFOEcLXFhZgSEf+Gahz67N7Bi2p50uyS/gOhcyAc
68WuMfG6p+atbGAqqFyQwLg49YpqdImppw7BCAn2LBd9wRHcrQlhh8FGZQtnF76A
2j507B2CJx/7+RziPqKfPj8ARyFLiF4d6qQM6HXV5rDThlh2l3vZVtbTol6x4fAB
Xql0q/3//zJQZ0MAhevZPKzQR3NM9klKXUymHo2lFGBUn6W7rPbBrsKy0pGgBz0L
pDxXwg5zNRDu8HsBAfeOyAnFMybMQT26YYyx7ui4Ozv138WYe1bfTKIsj0SuC9wU
bF/BgpsZDQ6Tdpy2wcIckafHb88iACABCp+/OF1nQlV4eDvcDa2MfnOPBmKrkI1j
g3Q63Uy/il0KETw9dF1k5YX3k2Pe5SBdTA7aOg2Dn7nAcGEAyh1/Agmcr9yxQft2
dOyTthwJoDUK5Z1NvwHu+oY1tcVHKMG/zZAaPtOMBMdFS2eIjYrZzAlO/t9lNnrH
2ZZUH5ukskgypQjCGDSAsrmuTD0MOjbXw9KIzIzg3XLRFIN5SkG21fQRjoOVAGPH
48OXMVrkHWudrdciLc3NCOZmaah7gG5/Oh4qFrwRp9CBMzHTEsX4kiJOPXNCk9J8
5bF0WnC3KlfBg1L5BpykHhHouqfYPMr89G+F67MeygmTVk5COBr20rfcHWkVqTBv
ETcgvw6rEQklShnPeSWG+gQgavtLPO2ORiJGqd1PPQFWyiUp2HwjXNu3Xx/bLY2O
CPJy621IAF8CyLhYIW1M6ggBQ/Ix9zd1PCAUK/C5aF/asXCWqw2YOvz1KdbdzZaD
7mzNsFRy5c6ZKOfkgZQYvOPFFcSO5GXAYjngc/x8vOjRZTlaUpqC8HlOZd+Opb85
ImkKDPmzywI93QAVgiUe3UKUlHi51AY8WuSi2v/eXG8zKD/r32M482Q8SN4PRY35
drK9/28ACAKv5SpaLnzPjGbRjtwcGrlek17yiM5lD84SZYdMJ8kr1DU68ifPJxwM
q/YzX52/flMTdq755MoQKckIYR8z70VRiHu9+qUgINAkNNFGfhhV17ujpfEdxfK8
hGRqK8sv+5QeLMdn2qbLWBIR8Vpwp1cWL38y33ldx0QAze4Wg2KhcL4o6MzrQcPx
hl6mYYVlEaxJYcB7kLJ52x4mZ6O4BfC/o+X6IIomLD93exQCgpkb30n7WCR+sqgw
aqDv7E08+9WKBwJZazgBE3JV7byNVjIzP11UBj+wnM1c9icd5yx5QzYN6oWpycb5
d2xRuUjEwyVA7CyeN/lvlcU8pjzGZZkVU0VCmLyQqZdhLEVRz6nncAS1QM1ok8Mm
omu33ofAF8dvXFmUvat/z8WJIYekNYcjhtv4AZ9+o7lekmjD42SQcsy47yomZAEF
Y78P3oJ3jUCB5agvfKU6/hFwsXHqq0g7X+gwHQnNdVicjqCKtNu3K/kO4naTJOEH
hjV4pecVC6kGRimMWc+nmThnELBBWxbEwcFRJ5OITiHCDyVDh+FC+Y4NrXpMwJZ5
LeUlEtf4UrrkZq8hxq6xVCsFnaMfCYphE3MsgRq9/Vb1frcGrhuPh61//XT03PO/
9Vd1T9HpSxRxQufFnLTozz+X/J6Pr7wZyOmtiLw7zJgbH7ot282yiZK3vHOCMUq/
WSccguu9Lq3oQ7kLcw+3yZjTL2MhjfJG8veURlKg8/+0LPrncym5v+midKHcw+gf
r+p2tzmAos3rZp82gKL/T97d3oi8HQAJ8cI9zAR9O5+hhvZ50V/luunMLGiedCYN
m/VIk/DAM2JnXVEjUwfWwJ5do+ZWBnr99PKd1P/RCeejyeoKbsB/kcZljp1c6my1
sV+ILyPpFkV4uiLXjyDgiiDfNK6uino3qepUZJqa/8X/kVd/rVeXZidy2QKQ/+zy
B4pKRoHyZgGUt0hNChrVI6Kdsli7P63Dpv4TX3X3etDFeABSs8pxyxJLo/QMPFGa
6n230zT23wAK8VrGJApk7FCYr2PV8UHcVJv+atFAEojmc70MpKpRo0l+dfjlWoE3
MPEhpkovBiMX9KeH4LN6LTZXG/tbLDeDT2ztufBQ78EJOplkwLlTGtBko1tNrxV5
wqSq7tQuOLZ9OkcXwUk+8j16XrM/srk3dAxYP0HFYk9USPALrcNqSSHso1OY7gnn
Fen9Ly7wg9DyYC6SV/7KmRzGsdBC2fA07DMVKDSSfjRFzWg6lmjWpq73DaTROS9b
ETwQ/Na1krC8M6IQvBqyUzMeqKjuOKtcyOVL14FGOuAx1S9kfnNgOzFQ9K0BCT7R
6K/Ry5MwyiKV2bFT5iPkLhPKdLZQTzxCZRWACq4goMc+gaKMd4ubcvndua7JgBh7
LGAO+dkaCTUPYpgkHd6Pn3X6Q5cT3YlkBbj3lLohWqVAqdjDqkewb8924RwWjmbA
SkF9AT4v9D5ZYaM/zhabGYRgjz9ricajMR9R4y2xtu3Gb8tzsQO8YMmMf7IPOmkl
Yjw9rUhH0Sb+WWdZlBhppKSzTgesOoCtdUYOa7KD1aawul2ife74mOdIQA1eSuRW
ina97ZNW78X/j1frRLE3TPsQ29EkWTmzvCHnUzruGKWWRSxp/q1VeCRkqDv3zfDD
YnWPDAFAvauiCMUDcWIy1q4I+YV752/QtNUd3xFHhOk1nmed4DN+nWmc/Ty7uVst
MNqRC8qMDli8IxoSBfA+6lKPhCY8EDNMNOWDYTjs+ZD2OHpxPB5ZKsq0213qLGtM
0UVQyajxmZUq9JZr5MEGDmkn89+TbTJ/jupSJld2qRcTn32MLO73DnYvVxFzQl7e
AWeX5oS03C/sUv5C+IZK0UsjJL6icokg/3RRu/gxeiiLVidEIywZl9b1mjto+RGT
2OmTMpMVRuZ5BZZR0PNLFaXYymg9+iNcecmXdXzYlPtkl4R7LdjM7cEEKB+b+7bh
OqppO8whgd0u/kir6OZz2tBIpTmfm2uek1h9f+ekhJ0ApuBDtos18XjRC4FhgDfr
lDdnfMx0zgK/Tct6NpeQ0wB8qIhD8jxUUtQbv1A5VgNpeY/Ubx/PBdg9MItfWvql
tQjbW+hU34prAg/knh8UhhT/pEnGiWKP4o3+DC6ckEIhGDMCk8MqgSLzFuCWX5/m
1q80iPydAO1aJyMrdepMpwDqXAHaIGOigCExN+PLJB8hReK9ZNRJZ8fhhID9XCQ1
T+Qe70xPmdZ2EOOwYRpSM4drdVxLpaCDLnzxlcPXbGvMPH37ZCbry7MUk4B1fnWm
wjOaJ4gmDdLU8FdPbWJH6wZXAC0vgQ+AlyJkn1iEsUA5TsDgEPE7+o6bsXt+6tOF
rsvkhbaa4AZl/DA0BvcXvm3XNuONDI7VkScoL9qMC8SIK7pBtXkj92tEEiWM4+mK
QA3QoHD9ikHcGuMRYz/C6PFqXQPO5830i8j0Z7tniyKdyNVXj0u/4qoO8CjBr1xI
l86s0g85Ir4Zh4z+0AiBbQovFEZN6SIF1yoTQnWqwtk8UWSbBugcDOsI/PKoPPVd
/UJdERMeV3e8+kRQM5lKHye+PTUFG70GuMwE0LhZT49ZS7n8cBOWxBw4W/dma70E
AjlU08OZhdIBm7VZ9tGhT3zOdiYD6KPML7tfUTaMHueeuQUbsM3cU+bG5HSSO7Co
GjhSX8JGZ9+kLd+j+WC2LSLDtAI042uNPmP9fDXjBKOb0Na91ip/EpJ9yVMWdgw3
GTT1tfmdByTpd9YJ3BKCpmxSribNbP57EsNKZlj6GEChQbZGfhavIrFpoVePQAT5
QYETwkWeYHaj3Ca2hKYKSEmzxNWLDibHTmImFv0Cuap5BWYQ3XgMknxnVlO6sxT5
OZsKPpoxTdyTbsk06cudhhaz2o2uLY5PuXUpsQWKOicaBvi9opwbVw3mL7zSJN26
2ns72GxkhBkoTkTyLNvSTWtYZhPznvew35Tl5rCNDqzQt5u6y8u4pFKG4tK9wFYd
77hGCVW4UgMzY1srGVUMhwE6NrTRFwIaebsWAzM2xnu4Yuec7nQ1BrJW6cIizX9U
EuOfVakIstIP1Ihh+L4KZvilRrIkFuXu0mVfB4CzQVNL+Q7AGZjzlO44nmbwrmZh
gae00A6Yr5R2l8AkjF1ng46vxYjVaW/OKJAniEX4OBehOVtlQlM/MwTZcVdDulYP
Y5Eg74J5lYD3KMDmSWyMWppoTzmPmqGlcInx0kQWzJoWTGSTlZc0vXRgyobX4hvH
FSU+ogwL2xli/m71TEQYlI3vclwDWxc6sgjArz4CggCTnB1EAvnDTx3GCDIOCWRV
PUAwBgSjCB8TItgD7LVMcrmfoIZaf3OAQGBhtIWsoSy3FPNtURgZc55/Ld+32y7g
aHeSAzTbSJPR7O/GDfrM0Mrep/Y/WX4Hk1jIzBViFLjb5Ge0IUhrvPjJU3CxXqvy
4i++cj3c2j/aIUvEQxMo4PbJvJTLt2Yuf01KMzqFJwVwYY9rSL/6b8RX5y0HDgiK
TtCprb6y/3XS+T2DZeXuSKTJILW0lb/0QyL+5OGQLODSPN2Eu6wJpivvJsIOiejt
6f1FHcmG+LbPrltvybbTIJvXV2G3WvbbfQ9Yq/eTkFVwu+/SwxkKPewGzImet9r1
sQy8dTTFkOdCzPQQcO1TqwvNULlDXnfBWc4vGT/DkYIuNaScs1clABx3ADGZpBOM
z0bQ1x8bBv14IV1Kplp2vemS3fdUEGPo3QB29qL6A6eHjfwB96kzWPOsakN3/0tE
lYjDpTuGV7ZsFdU4G89ybbzrZrAbGSCIo+W0iwgV+MvKVmRRwwY84/4qBrrAJVZk
WGcZ/2NCd4vTetcwsXzvuL95wjRCVnSf4ccaAyr3nfUwd3LjynETW4Fk1jUbwsvf
KSyV8FA4hDIBsrDVxggoAQtwr3jexBXhOjAmeZ7URaG6Ho3C6Dln+wp6ya8zSZIb
1TPFkydaCktAhdqyOKHL18sItSvKfAO6egoiewHNZ1Td5wUV/ooSbtEQ4IGLWutG
gYN/DW4GzI1uCEUrCox1veP2OifIPjj33ur61qY52ug5KiqeLAwaqp8YQkoeSDWp
5poWZiRAqJBnfj4bY0Weuf7Fdgc2GsKcsjrgPjLir+d5qEh3LN18XaFF+E3EFWGy
WvYiLcJCQMAEAtH8LOMMK/5KVDFEK3j/kQVs6OvBVt82wY38PgXUvSSx1BoLXlaq
jkOiQNaTucLgi1jXxGWpRZSOUGbHrkvFK7p+IYWhPSUMAdBN9K47BVE5SHNgsuDm
cDQPfUikq42qcvugUGAk/tgDK/ncWDRPymYE0cRzcbMgaPAPe3wX/s0vWR46l0bB
tG+bVNGJN1NHU6GsNXUpmqD3QKN9Fu4pWA8bE4Jng7F8f55Yzr5xXW2u7nznk6j1
iskuvlBalBtye7S8GBZGBc3Z+u9hVoK97IgU/P+auvgOYwZXKKpu1hjxXDjsVD5D
J09pFawlBqXabU1ENexLnTemXW3bAM5BF8GK+lgYE99TV4zz2MVbX6nI7t8eLQzz
cEYfr0XJwIKzx3C0gHKAVopZP1j+EJK/FzDa/xlWAEKpfkjoA5HicZSB6Zr7NEBs
+aUJQwqKg1ESIxqjwTSUeq2XKYGZQwP+6fQlmVuEUbNNyH2fuD7MjZnq2x9sJmTc
WIA//xp2wwPuNUzIlyPoLlONpbF6KrK+3zwldqgdZjyUuZ/b704LcSeoHE5G5UAy
tvC2qYjRZYaVock5ch4EPaSaRvUznBfL6p4L5tjAnkhXNJAi9hcDCSJe2XyEAl0j
ttcnum8Svo5H7JHv7kCI4OwHkXmOYg7Ygaz5/lBAS1kwaHhYsvpYPlDd8lhsu1KJ
wYWc2n90nuObsKYihRH9NSsVtbZ+MWZelUPcagHnC5IBHrak6tp+QMtOIoRI+1s9
WBgz+1ybR3jztCQYeXsoC74jzrAu7YRH62qx8nPMLZYPrQuZwDjlf70RhmStp5c5
RM/6+neODki97QgcqonywQlLZC2MSuJGzLjUnuIzef0YFcAuitqWD2j2Z2Petey3
LJsivL1tjNKoJcd4MBvytjjT666/JByGqu1C0ulzOR1424dYlS9JWcm7rHy3iMni
LEJkrGhKDYmVFDSzbP+5RFBxPJf1MXVIyb8WroL5ny4YtxbFxj1iDmoV9J0S3s4K
k28ZKWSNQC2I/svTa3ps3VIYJalYPht26OE4W88R3hLJ6NSyCW057035Qr+dhti2
3Q7/AmPTNCntR5ZHyvPLpctInUEQY6onw84y6s88/Icwjxt/9WJbxa9ZtdYprPVN
oFgBfKHt+wVBJgb/esLLXRXT/aYJdHirQ3Sld37hZA+BTa1lVUXJQSEEGpn3ZtT8
EOi7IRd7lejpS/40fvySJU4SaY5ichkGatYLdGn+sJ9UmxlIaaoe/8LIrMrETBBr
LzfSir3g7ms1YaaEeBBIYWKeO2MeBswJPoE83vsuohLrfXYsWMICJxSgl2+OQobW
f/Yn+vljO9u66kMMIWA9dnadIHYeZL1WQ607GeRIU2xWDcHP7uMw0y1LDZcbc/Yi
9L0CUv5jGQw+0iKRXCW9JsjtdE7GEDtLBWL2S4RD13vNFpFvYHekvSYhobfBU8GZ
iz83Y0LX9Of/kzeAPbnBN1fl8AT8rjI8l1Jj3rb+Oi93AzBU+Y6mr7kSD7xrzh1B
yBnnX11pNYaoqAHdwkLtoUDTr0RfmLDPtcwZ8vg8O33m/yUk0i8lS6t36SqYXRVF
gUfq8k78EPL4g0H0jEipVs6L+g1Ov1uaBqkL9N4+rMvfn7ZkHT5skHu96G93sE1G
TWhaQxrhyCszaqze0hw4kl1gZuxKvdwg3epp94DMM3vWU3Bj4iaYfFIGVQvPgKHJ
757gPw/jhrAh14rCaOVMTfqFcslu9vZhHgwzplUeZ8D6ye9KBBPYXHKqALepvPB1
X/BfiTkXTMeiGbGpesVdCkz6aOnfHk53BXMJP6rpXWo0OQxmw5KChy9bZaH0xmQA
xUvSJxXphjEnGXzIinZ61itJ3Ks3lZuY+lwMBxdV/tl6QoXrSNvXUapp1/opzwjq
eES2cpx0OzAJdjqDmnDF3l/zlJezzCm214wZhc8+fpK6BmXb27H2rreYsBOSC+Xe
ikhDg02Qg5AxwS/xY1Gnzve9UEXGy0RebJsQunUFkXEi7wFhMs4jY8yhS+v9M3uS
82TCanwKrPlKZnaiEmvlHmSPP1celfNEpGJ4NllSVBqJFP/dbmXQcWkb9tBGXhPx
510ZdAMPvV6Ue4SW+8/whLACuagJH2IedPioAOVZmi3331RtNy/m2Fi13lERE3+y
resfAYl4isH1v8k46uaWp5X8oDmDJQCOCrE9wUmZQbHy7RikwxG6wElB8giNfkGV
9jtuud9vQ0OEXa50/3/xbNoijY4UiPKOym+2PHYsmJCnuVWB5eFKVfs2njGYhUVA
SvVTcuwwY0P4ku1pk1o1M8Ht1FPO83iGYJKgWFkU9I7OfcuADZwegY1jirFKnzqX
3x9GqZ1DII+wlRAF5WuovYzzHejRZJVHiiBSvgbWTaA8Iz8YgEOq/nc7DJ2HT86q
BpXZkHIk1PtE9jaOA+glgBwePh6xIEn52EbR9X1/x0T7pZfbW78KSQK2+zWsRY6N
qsg5HU/pbKXVj3CbvXsGg4AFVg/LMv0qBKvfSryw5V0uXPnhrKNJjQ2e0OyMfrto
+2uluFZQbLDXToIi+O78FIaEV5lwM9poYCEdvmgNyDQMhzld5U/9NQwFpJpNGiTv
TMogTImSveY9iGtckcIak3MXhlGZPWgpLk6PJW1nNy/hsglaTNXrryIN9sKNgmko
G+5nxe+9oeeQi6sIaOXise6mISc1lZX/+B6KMrRbMn4NnrOXwGEorLGQhegsTPAY
BWJo+qRycfiJZCYCBt2O6INGprPcFZULvRyUP0mGFL3j24+B0wiaZVxzAvP3+UY4
9wm7naXd+YCKPqQ8GHfEzy79Xv5gyagdWcqLqfksazxC+/DboDGqTRPDAW/4lcNf
Edv9/bzyuQdXqf5oupPvuajc6+3phHV2Eh4NAATpcqv+AYDMpj3fZi4hSPjYZOUO
iruGxU8QxWoDiyuuavVkyxgR2d6+sKAWOe1jVvd+XruDqvWplCBZp/NmVVZgrP/h
AJkkKWGKo7LliRQ0I5F0ABMGyN4OvvilPqJn+pFqbIWkgLWbYIZorLaQD3lw9reY
Xxtsvwy4kBXQCXxX/AMvX85PnSBaWJ5lKz9VxZUU+xkgs/TKERH6pHFtZ8v3oDY0
JDRb0CALFY+IcmgI52mhZaSAUgga6QcuXMJyY9e0X5r2kn9lCB6wYdzugJ777xRY
fUloBQx1xnrYnLivW6lBJHKZOVOb+WHTrcysy3qQ4kWpOCpKoUwKDozpzrPKk+Or
dXwKGY+NG0Of4kHfQOjPFlrw6sy67MiGbiXOLbHc98BaGmJLTvb6LMWt8SG9JIEx
VCq8jp1uonw3fSZjcPk5jxF+TMSc/DvB/Qfx9ZutmoLks6H/wqEAQlBzd7eY3GyW
v8F4dYEW4hmKH2QNhEiBEamCLWUA8EVdDIlUIRyfdly4ZUIdkAkrlcGIaUmpSWdp
7xJ3EzxNwo+YjKVTeoqFFPbOmdIcX2DjflfslqcNfCyxK1QkwHL4ip7j1g8nomI8
FGebpsk1HRtiELVWK5KRDgzyiscBJDB/Vutzcm0UdazmvbRBlUVBju6zTdInwepv
DZ2/OOcikTBlZsOBNY8k6/nMoihHQmRGYz/XlMxK2HOEDaKheLQViarZW4LG1y/v
782Re5bh7cPIE/FZ6vA7NDL/rd8n9O5TlMj4wPtFBE7/gm9IHjeQ4OnApa0tDsbA
foEo0kuvrr7DYrKFABH1TeE5OSORWkfCzr3GszGR+SGn+hWOQiYdG0UPRqTUsvWG
LLzn2rbEcIx/be+mTjqYgGrcdH6hYsVywcRCTLy+r6ia+YH7+1dRZKoa/Sbhw4jT
ZeMj3z040TYaqYDMJDX+pb2K4b+ulJ6f0fkcuxe6Lov719vge8IAuAdPv8/lvnpO
HjHFna3MEIMKENxSxQFDKrucOwfeBc6O0dDinVI/dtBM39BLnDrQqIe7Qa4W1+Y8
f4gGquUc2xS9qtOlfAapAJMkQ1JuMOqaLJJptO+Rfej9tjM1J/x3k5ibhQEei5Td
UdWVlxZfKkbbG2M8z0I3SD/XdklEhVDeUR+D2FbYnT3ot12m7teVta9MwVawMMAv
4lKdwb9RDh7XtE88OXwlfq51e42Yc863zBcaRycWj8A0Lt/XO2jlPahCbcz7cFpt
/G938mz/qCNHM6C+iSVmiPKaqizBTb8xxkv2B+Q86t/0iEXQB90HUoXbrVk8m7We
Cd01r6H98DRXSWrVrPIIp3zEwwIdj1uL99euH1PgEvq/FJNMuseqZ5Ww/5wHYlJ8
MmZWtSgojDg9AdxTUhnJmHD6hIKdPHCLSUwasVNyN04+m6PQcuo6H2TvGpydhRBE
tnaq3/GdpZNtRf1I9z4x+bnb2Z3WkFRktzZHf6rOFsuBy4t6lIHRbuNvfRIuixrg
ed4I6csIgD8X4DXgljgSi5JMPyDngxsXN/VuCub7eFxH9boEICuFWAl7sVZyjPgd
0H8CtaSyRBTfMadQRNdP/6ylGckRJ8pOTB2EFVLBykkOpX3vAFrdDPBmI4kQQmXE
mnUYa1Q12o+Ze+Ed9xjAqRxWQcfeq2a3uI2ypOSO8CaS/aDMV4m18rVAGmqGyThb
tGUq9iNurGNxbdDcARCvJB0g+ceFTTBq9x8QUrHl0/uKDQcJzFbsZw1B9P+Fk5wk
kGqK7hecdfneigjCUmWfUwaH0JIffrleeKNYmN1BNO/zOmCuqHM1YqLz3uLTCr74
F1YVEc0C26QvQg+AjrTfLXJBh7yBKAQTBm6FxkPMZ5/lgFLy+HqcVtgzgX70BFCb
Aw+MR8ll685B460CiZDTpIR2nxt7D+41DDUh+Wjrn82OWVdZx1rRM8nqOAPIGaNp
afqTdEKlGbaQrZ/9QFvZvCFuyZqh0RSGISJbzUDyx0Wyj6DnobLT9+J4FBmeawb6
R9E0b16lBQ0j7PBBUwWHfqCaZ+Vj2nSdH70YaluBQWjkvXQ61QlvxJjKoQeD3dyH
6rGFuQ55VuWs3DuSVSS7N7LkUZvDfYnINhU7iUjgbrTPJSJFTzUfe498MXUTsrmn
9yTWYm8p0H3Q37ZOXkoXw7FTz/FVJGyP4uKO/nTBxH/slJdoqiJLXzt9XuuPE+PW
earOjLbhvbx6v8yFG5RBxPfD2fO9M6RNJvpOtADQnmwaLhi3vfCvJm2mXtgTAbV4
ClnsvglEU8G8PJdHIpM42FuHk6h5moXEUiQvLbAp5vE/6rvjh/TqsyIG55fG0Q1u
RmEUeeDyt2h1nSe/6XLTYDDjj1zKmNlET/XemIBYYYEx+M/zmZfVL+R6OuDS4SyD
/eEAtFJAcVwGiM5rUeC3reG792dLchJMirD+3Lsuhtz67Q2i4yIR9NmQL45BW8h6
4+JVuXK8a4XR9pv5X1ctK1VaZxCXMDBhyuXmWiS8lAOQ9U7Hzw8nnolUGl+NF6Gs
2jXnsj8Ho+acBK8KL5BE6Au/RJrhB8/7pE3I3XX2qfqULCcCdTVxFzr3pfLncIfS
pQTKmyDIz9CPnR75OUSQcBGLZAsZulgVPHmq9sEfH36pS/aQBm1psHJPGS9RMW2E
xGJJoN0SIZY1augsF7dR2nvhFAbiOOSI7hmNDZT8+x/defV5lfRfp/5rCotV8Wql
1n0wEa9cM2aJLBxxamgWSKmgvku/4r8kQThzckcp7iPV+loLKldx0ZpqZmHHPIea
/OAwp6BoeI+ftv04M623SgPEWfLeR2OMirDkKZ8l8B1iksvOzqngens+Pw0OaSWI
cu7GWQt9Gr173LqL/byDmFIvgepEmtVDxYur5pdKZZR4cgd3LJWMNqcimY5m8W3t
kEm7NEf0EapMGrYqO0jgeZUrk1BfYaYnWAdStN2MP7z1ACBfUQb+sAOhwB50yopv
L/O18dZ4nI2xTX8mdOcdajmxIz3mRDZlAX5fj+aeJy6vCgAGqG8PY0V2pFhk/+0x
Lo8uHBu5B7MQzh+Mv82MazZdpqfvP+cJNwCC98ZYOy91iERipS+mS/ufI/yJwqYq
WU4anpu/jhmjqTBEs3eXSc6PIJDHggwXkYQ0ccb8uG1t65Xl/NKBTL6V0vEgg+hv
Mgzf8WbIVwMDmKLwM+cRVcAVo9qYC46+lqundAwmKPCDPGUEWEVmv8lNREyb6+hZ
fzcXuZXkZwkVNZR/LMQ3AfK05IJgpgdZ4Av5eca3jRgrUr6wvTRKGy+8Oar2CHfU
SgRsRjFgpvZcgqMX7mTkC0jmgcPY2X+db4UPeGd+1/i5a7wUUC89x1e98INHjDRi
b/8M0IddVWdYYb8zoaBIura8SOPDkPNyuQB9wokzdNIxsoXCWaffRP260v480uhN
Ll2GPOQPQW7I8yOcIbfYgeCzdZY1y2BFAm+ohnO6bWfKbBw/AewphBvg+/iqe1At
Sg35GRAkGFJEb9ZCuDaCLHY2VmGIXHkSaz6eWZVST4WkJW7amonXyyW4uickXysA
oV+TgY05JuRGxYXLeLC897cpaWAGVd9LHZvsyGq3YAPAfUqRt/JeLKp6Z717wScO
HWpbigRTtcCnaR3Cx/YGhE5qUGByJaV6EB9/Dgpcx0WKpX8EzaAs4jT+uLgviO2j
BhlXbROO/rR7dGfsYLK/6ZhmBhRj0DuGNRNpFt0aLhkn0qTDPnEN8pmOpS40xriY
WvRzKEdazTULu19iGGE0WrJS9bTjDhRmyKJN+4U44gy7+C9hG0dBOk08DrXfxjBb
RqSavnKHXLrwUfg1pPXaaEzsP8O7xA7vQS6yDw+m9FjP+yARksRfH0TQvm8JUaTS
CIxpcO3dM4Y4PGkNHw8o+3GMwdPyx6LEydfov7GuLaKEeX+HYBFOiLPNYShlGYqc
1Pv/DU5CUSRQOrzlSQb8Xcw9uTLH+GeU4E7vm3X+pCb0LUm1oDvDUPjNWTC4gBbt
2YDicfNJ1+WPDFPT6DrJVu6DmN575LD97YJOpVtxuHX2SbsFJBvSs7BM2BetEiD5
4PSM9lNmzpwuyyoq/TsxEyZNdm2gqECOScBvnDUj0vgiWP4Tdjrjl7gUBBwFuYcP
g80M3+ZJohuAzisQtu9LxF2pVwS4ekElVEffxLEzXKYG2eUF9ZhnRvzU4c3yz2J5
gfPbnsDzwVXRh0D4O27akejU0PzMNC/dH+o0rh+Ua5y/ZTiWtb5cDyoeh6kbYt+F
n/LdoL2Axodvl8DdQP1xOciGTXUUi1dKdMqZY9wFqSlzMYEOx4XvHnsoW0Fh365n
rmDqR9XWzmsxFkE6gqSul6TaGDWjzK2mR04GEOUNcNA+w9K1HO4RCvzWdEQZ5Hpr
BhaVjndhPK4LG6cy9sVNYWBwPzB5N9kyfey/noe+JszGTml2YySuCI1L/y76zmKr
6TOAnsJgRL1b/NF2oAcX0YQc4q1LyRt2YIo7LLVa8uoeB4/rSCRhivbdV1gGyy63
zCQL4SYfdkn+VEPyrYfXIuKzBB31tA5UqqsZ0eFuX39GdbZ97aN6nQH0DgTogwZx
099qDDM2s49XH4t0mWF//LW0O4xnrtYR5qryUGtYhDj0ihyVX6R3BgaLQhmXesib
mChbYTPSsfJBeVgepg/ODQLpsFMo1UYMK/NUyXE8GCfiJGEhhtxGfqV4vB1lMeDg
TCyhfaxcZ5LA7ykgFNBTN6dwrDNQkjVIswnuLHy2RwcCu/mlL19hukYjBhiTvcgo
uAThrQyboypNksC0ucGx92TVud4da7ymruILCCmJGc1dsWyUTZw8n5bG7Jzop5XW
WeIxZNXloOBH9gecZrMJRA2TIeWeMJ3elULQpXKx3Z4GrWyT0p7C7juELLUqVA+v
nsIuLHxHagDmuRj7I47/fhcKJVqz6lrW+HCj25Y4tH6JRgVp5yryw063B+PbcSio
Xop516DjPtnEGebdRGKr7ihYv52zeR3w/DBUW8pPPRxS4Ac3K9dw9atS1gFPmen6
wdoQdnCwY5nHgNcDrgkphifTkgUOVen1hz98hf3YU5Uo3ANtqoIGPQJvkwAvbLLu
z0+xltYv+LD0oAM4R1X/f+H3CKlD7GrH75NmPfCynp5Ez48vNapFsCjvTprKyYrE
Qdl1xzDsNMSnbdjdz79voQ5fNYxKhjfeQJ8siEVCMukCTkAYPrRgsNWHuYsEyXi1
4q5MxGPqUGBvMvdNIP9cvmydoFb3jIvMNvfDQs2h+Qf38bpW8vbaRr9jm7YIZYTB
AVeJKfAd/xgZBK7cSmKJydAPk3wdimswfDO+GaM5qter25Ud3jfR1+aggaSZtfJt
6BLnz51p2PJPtyyPMUJbOsx/vhcq1D2D47aSRlzaEsFjz06pChxaVKcbaXqRKjKN
AF8R+K/48gZrTvCQ79kFgpvzxojClhxv4N5ovHhPvbispZShxwpCUU/I6TX2KhrL
1GFs9H0M8Dpc/OlqK9t+xpUGuuJ+sSW9A81y6u6ZGfQgV4EYClKKeHJGzsO/GtnC
d9e55hGQVQiV/6Xjb1wSv/lCrwvh7vFZ6ve/noNIYif2YTn0Jq6REIYiEtra0Ca3
4f5A8ur4sI+Ikl5zSfp0exNbj1ggjNnJHC3Fdaa0E3+cSoH36v9L4B7JXxv/SFt/
c9gGAu+T21zLN0Cc3DJ8OpBcdQFQsclhjcSJ88YpGAZQF1c166FzDIMyqb3zHJe4
Ec9G9vkyOqkToNI+YjPV7hSUgv3N0837XpCu3IY9TKG/BbsRvS00ymDw49n6MJFf
xwyUp/TOs6Q+owaARq3gTApy5b7CfJoezaa+o0ZXNv/NwL5mhnBR7jPOx5LnGZHy
zS8srwsREMUR9ySLYA+mv+qyVP357QW1k39luUCX2X1z7ThJQlsE9fPUoFaE4BvX
fF6cKr2gzNdYbKhVkMqwKK7Ob+Va59n2UQQYfVuzVqnY1z9zyL3eUeFEeSj69zJ7
fB8CSGGvT0W65mBZNAjf/Jmcf5OMmmBRN8S6QMNQGZZdbe+efjd8v1bVklMf2SPi
S5Se3GSKVQaFoPXXp3CFEwukzQ0WCEwG0Rpo4QS6L6ccXQ3QEOvQoHJSIn7GiviK
p9kgM/sQ9uH6W3g6zWmsIfj9zdRLR5/jYM86z7yPUYrNSHz4q9WrG3syaIT111Km
9vYucDDPyzgQYAOFxTDc4uw72cad23i3gaQrB93zlpaboPDI6gDde3HWu0HlfW5u
/3sDPqY7UgbpZYRCSybz7uBSp+eH+1nnB/0818uHRgbjVe6nXr0pZNTDAMVgIvz6
plhPe4ft0KkkDhA1pYJFM4EiA42xA/k8FxlVvKRnbSiOY/Es37xeUEJc56A8taOk
L56uaiCk+T3oPXfoAYQpZ9iLFhusVLBnGZ64cTmq0vmprvRxRbgHCf0h4+NXZCkD
dCsRW7eJEI0eZT4fhU/6H4VRCcqzgB4F0BXhB8Q2dBSqMroDokKovfhh95fNeAYy
EOS/420xq3a78Cmy/NK/xHFV7h2/6ydSrsq0fhxRGPE35pqjyGTLeZKypYhDVc8d
YAhrUfhHgdAFGvao1vLwqgt8GLBudUosrNoDuU+N6YjnBcGyt9dbwNkVrBt2GDay
JMjklg+X8EmTZxaV4okeVKeS1EozFfpNv61LrAaxff0yPqZV+LbFZ8aADem9qQ++
sOOVrsMCcnsviaPd7xwbi2ExGWveYeox/2TFS0oa+reg1SDyE1AO3TMU0P60uqvX
TKkZNnNQcDQab7IpBKEd1ThMDdOa43niLxM0/d1Jj2WodBCW9uCoDXl570EAtYG3
S6di8G4XF4jxlSfH9+eqp3a+kGHLkFK5t9h6JWAlffsCK+1FKgvSYKEHvakGSEOH
DsZDMeYEgURQ72qQ8Zz8q0fIgI2outOiULm1CvCyz/PuGq2YT2LShB19hgRfspzW
Cu0iPjlO3LR26EhUzm1c0Klo01mOp4R0sw2im+aVy088qW4LDhIPqjce2kWHxzB2
M8sN7uoxXDG+DU+N3BaQ2FaGfCgS0jtTpHwbq35l4k3n9Cs3UzM/eeaqFNNNXKUw
avshn6w0gtvJN3f+uIfOUKIJ+8IqKYfBfyUZ0DoyJKp45byHSN10ZDtGVmSAGrpr
GDnz9n06KDJUx2pRClG/vXffqHcADf1BHFVplWPLGxe6a1LkRRgprG5Zegzb2TyH
ZhkuTSrKT8tohYy6Chvl/wUgaGMQLaPjdd8mBLNCYRTMFscmDKg+7Ys7nvbtalkd
zENdddmGX8NqJwqhkyxqKt3teLkcn9SqermiBUEKS2QT2ZpTtih7gAY6OnQmZYd5
42zg46qIKUalabS58PL6DzK3sPdT7DgWWBb0fpSsTClw2FEKjM1nDj7AJo+/CTuz
p9cGI9PfJWrQMPsVALNZZUdsheTcT+tDCWO3qqPl+WGJTBOa0HLt3Brn2JlLrbhs
HUahXyYCpfR96FEzXgABf4FbtFdq0mGjY5TTuClcPt7MAGn0hGZ0hrJLRMohJXXP
yjcwn6cXKJx3Y/Vee/RBHL57Sx3F3cqzGZXPQFb41L/Xo1S8O6B/uf4Xlt+0bF64
LEMFc3F5mT7yFKo6ZP8f7B60VUOHyo1WPQ5gz9a37khwnUDqstQY3uve8WHXcg0d
IhUKFhixRkqWeMRzuH6rO2Ow6E2ITNiCYhVkTI45EJkJZtRvwB/p/AvFldAt+xrP
UwJBUhoqhO7yOLYfw3I9aB9p1hep9COWP3bB2g0saE1gOXRpaHgebMoQQ89qH5Yj
MW/7k5k0CjoFH9DhrFaFQnmLxyFqESbD8h2VJJWUxQcvM4KFSovk9U6pZimS9FXp
4KcqpLZtAqh/tRS630K65Vp9RjzqIWYZXMAdbVkHm9SoPWKLsJvE3r63VBO46Wth
qNvHiOiUf7ALVo4ANomLX93M9V0ORkKN+fkqrAdebbfRCJQvX9J3wnqbW2S7L7en
x7yQavQ3ylBoqgp9+G/Y7OR/X86RJIWFclrh/VOQovkaS+SxG4U6OGtnUYtekn7y
EzkJr40PAuu4FcqImraks0d8PqKwR3+ilooNbheMzQQU3CD+PxJ1qLAi9FUFpAML
cwbHjKmA9QfFKKZRa+Z8S1P95J5SlcSfz64LF3tlgVFUSt4fP60Dwh0kage0etk5
TAhC0lWqJ9A6/8jP4IHVmb9M7UlfyMRQmAfhvTb+kREdGb0+/IDmBv6PyctuTh4N
B6Ok3nSlztZ969PRjR0D8um6Yz/36dSgab4cGC3uxHW4qFqrX4F6ii6EzNUzzHJW
AEC5Yr/EyB3bWYHHeA4z08f982axXtsh6sxWr7ECYgFmYbJn9RmzSiIE71iLfSOx
drgH0ng/nWvMyTtRMUC2bSsGb88I/0wK31HYBWVKVAKetQfpngr0yJ4ko5S1laB8
pEQHihgTHbl130FoXWhkZAnaQNhIWd/vMEv4A+IkXYdk+U7gBwLdbjEogDXeFRo5
9I5hEsfc8EATULLItct4d5bTtlsKB6YqozDGFY9mRRyuv+Vmeef5hnxVbOuKA6s1
8Mx/E8SZLv9CmHcfH9Kez/aukiX6gQdE5xJFD6851a5Nyf8DslqookMdxXwuhXgK
WhMW4RSeBxdafmExFX8+cNX6fJB83F9i6tYgrJWyYpIGGcg4J9nR2rthGpvFin+3
zbOXE4+4Rp6TjJkruWJp2L4fDyBhSD4u4KaNG+OuxuQaUgwTFytc+ENwcQg0b8kM
YRydparM8tr9W0w0I2nsmV0rivSedUOiYz9IwAYGIYGCPyC+TikSchy/3H+JUP5A
tx+6XFYjOJY9z69Jek/N2NGAKVrrCjitAHanZNHtaQhvXwrcbcJncinOsdBC0Pzg
awq7KYT9ABDKcTpZZKAtGClE31aFKPMHMsS1ngoIEUm+WUZkZzSXqCNPRdstzI/9
48ecUjRLkc2Qz7n+palKTYWbDMIA7IVBSbdimDCuCsk66KVplduFZ6M4BHeMY2MT
Q1Wj834EqZP31hST5yql0Y8XjcebudJ8vRWhckgL2nSoZhas+SgA9D9etvaj6f1f
Dq3u/FB6rHSBAV+sIJHhwfE+/t9S3wWJ8At/g7TvXpE5Ud3DHdrLNk9G7zDOW8SJ
vkbyckbSsLwcYvr4uZi804IGuPVAIwi+pk8AKaIs8Dm4Zi5vVdYs6Uzioa8cedhz
flWuvERRNZSJdWqNng0dgFjsIG+SZm45PX+BFJLmdLcPVYm+xcgiQDrAPcWPv6pB
k3T9bkhkasIBJNGAdbDF0hU4BuOjKyC79uIUDMmYavcYITp/YZdiwWhxJu2puuzf
agZtzs/t/zvukxM1vymn+q8xOJdUuV7AhLIpucj3abfJh2C/cea/5SHifjWyRf9Q
8nZaMF5UbvyXkODb2b79fGG+Ytc1TNkl3MYcZGPQnfU6Du5rB/7EuqNILohFkZBr
ooTPK4nUBOprgXOrWdDrzpg0HvidILbhHMn6e/XrIoGiZ7g9M+lFDsuXZxFA/aNQ
H0AZDWmZx/4g9QgFxur5TaQUjYCcYcXfbfdUsgDHsXUKfaIijsDE+HIoemsDqps6
YW116zqwsOvIiskUAqDF63tvGtd2VWEQKKaVstV1t1nTkLO1xuag8IRx0g3lk3FZ
uqGu6EauDnSsPznOND/zbOeThYGQwF7Gq9dUg9f8YEm8ujhjii7pude94Hi1Srrm
GIAZ+pMV3VNoQbs4IMDZnYi3b/RySQckLOny2TZgiYWyXHVp1ayhK+UCyy7d4rKf
0orCapmkBhl9axf7LEOH4zATHidNVNc/l/PPj/pJmyIy0kSxbgmH+nhUUdVcDnJa
EAOskotpRepGRg+8JtP21qKYdOILQjgQ/gwUMw9iUiLYQLARGDeGqFWztCJjqqBN
WGGuC0grEXg8OknN59RbEoapdvsFbWdHnxaoZ1cT7vLi3uL9fZgKe6e3wv+MblZL
qyBoXeMokTkQoaQ1GfgWC3629MAq8nXYxXdi6z4wqFwCaCqOoyJACJKHoNYHl+5D
tFRKqfnkU7LHNxGXwoJjyl4opBSlk3aaVz6bOaTtQlfOKgddKrwu+/lYjG3R2RAw
8MiRqfMZGOckWWP0cDoaRZnt0/4LKvHhnlZnHjs6TyhLYOauejTF0Gha5wOXEcZd
/wShkiMUhbxiwLrjMd0wVoQZoBm8r3awCHCQBa/5WI8kFR6i1EEFMJqPTJUMhXhk
X4XBTx/ips/v7oqpWNgi8lM2Psmfk7I7QVfC+BywEi9zArVIdHsBOhcD1b+HYLri
UByvl7Hk4HDqorKpQVEUVFY+Hh/RnywZaZlId5R0D7qGnOCuGnw8bH/Sxp+SfBOX
ibPy0n1G/p0TEq4pkW7kINt1vCrSASaa5k9y8cAYZzI6fOZdg7SBYfIw2/LS75ZM
NgpmsTPQ+XE9fBldUsErCY6QjfoT5VwqnaLsW3gHp84l7ejEHJQSTaOrMpOpQeoU
A5EoknYGQWspWwJ7XpqAJ0W5c4peiacUr/mDh5OtgUyFqEhiOtEEkJvl8qnDH2R5
nCiXfXq8vYZq2EflUM6QZ8mGqMDMkiaSynZdAo3d1xeYyL09esM3LTwCckAAKZDp
IzdYX4uIncnhncqrbOF6nO3v6cXh+Qa2gLfph6tNCSczy2uhP+tHzioNUbOymBar
17ZJ4IHaRfoXQUyHTZBBmfGDJZBJJ/Ms7QsJaynkXL1S+CivXJYE20UnD4XpL2Lw
Tj58HR7dwbcV7i5hH+0+4dZakrDm6CbgGog3TAYbiVgogHevhFbTFTdVhQdsrDK9
MumUxJHTxcFKZFUEH/KDOJI9XXMooTIc7qk9k+YNjGn8vn9RTfx9NSclWRlpxNYD
u28L3Qe4dlMTmkisNffIUablk8WdMbPOhxCbq5LVsJNR/0hb+USJ2UZyzPIIvTmq
zcYMzT2nC3UVoFThssWLDXwHOmOLtq5y36y9DrEYCJAEFM1RJWEsPp4mtCEjmlfo
N4AKZs2xyJNsjgpCUW+BX5hGrMz2QbNx48te/OC7a8EtrcBYQA2mS1MjzqShEMQ8
FgzDNPWd8ItmjqJl26oZOVwJg46oJRqDll3XMaxewcmf7sqf215YBPAqVynU3fd8
fZKxGbRT6QNGERLSfHShaWDRGYh+zvhElYz/0jSV95YlfaegfHrjK3c+b5KQyEtt
YwrAcay6DiZHeuuYUeJC5Afwr4hWHSWLhxRiaJRtLovpkheoZAihGBW9Sn6AEu+k
rjmRLzcroBfEiHheZsb34ZwiFydyDN55Ri5ZxgTnJTpoCU3aZhsXlgD/l1f0UydB
dQvNlOiJSTXeYoT7Rtkgozg3no1xM7jmsR6P87WuI3JiAy9/lkL1BoPVLJ/saz1x
vi/LxnETIW+ngEaU9f7tLqArMn0qF6lfg8PzClxSFH+rykXfBHu4gkLhli8fb3O6
aVlNFgv8BQ4gObdNxJ7DylnoDGP3yTHYAGHV9HT2TSmKnUTOJUjtpplKNx7+C16w
YxDA1TBiP2fTvGoylLlwt6P2VnKP6eRQlnCYnSR4Ar3POgJzXZ/nqGQdBWmictz2
wBzWjxiVM1FNM5R7JwuqKTIdBEWWpw0TsnEzwdi/PHN++mjnjtMSZ3KzI0bV0W9R
w8ExVr6upiwZ2TlBY48UHu4HeBMS4nDMukw9KUeMQESV8KhWRlEINFCuEfiahK5q
3QgaqION0Imt9C4MvtEoR4c9Ht0PcFDvtEW7LQUbOE/ojgHhjKNxCrhG4P9cw0fC
khmUsVXKR+8lwCK9K4C/gzxvyiCxYbEninXl3Wee6Lp5VdlRfLAfsvglg7f20SEH
KB2h1PiSEBNkI5isGB5T8qqGMVVQ5koFthGB+2u54XLDSu7V5DQp2D5+CCbgf3C5
J1kLtiRFCdxWpQwxc84Cp8S0p+lK+Sm3L2/aLttJ9VZpBsjPGXWYPrP38BlM99Q8
1ew/w3hiGr4SFcOL6O3uQ6NkS/T98WEZnPOQNnahNFSVBiSwGyNvFhDqNYVCijie
c0iuDZK4djmbLQpeRNTFiwEuAFI7pNCLu3kOPXlKzTfN6dT0sbgabns26U5XASDn
949hJLXsrRBMrmyshUX/CculxbF5AAWb9vMb1Ygxsbd2tBKHFcd1hwbjJy2AQSZ1
HHHPJQbcewt3weuNiftJv8Db83Fbz4kbaylw6rHahTF/20x5t8zpZqWnM+NB8zRX
hwgbXiihkLqOU25gT8Uek9WfaY2+hLoffOBNJwttDZWfR4Ue/8JWxwaxiNvMElwR
c8mPHXfqYjyXzDjVibr18NXkTcU/Y4gSwuLx4VgmJkyCF4sj+U2tewJdI+cggsfD
XXg7XU5Wh3Qe9YnI+c+kXVJdgEjN8JBh3x1d309P4K726neMiQnK0n4kL/Iy/PLz
OpkSpKnrJ+Ev7dPEuuLbYwV2uah9a2ySpz9iQYNUWQFkDLosBqF9/pjZDDh3GaWc
Fh8ytdtg2/GsHS8wi7QRI11wXVYg+hxpa1um9MP99fnObXChFWrVMuUJ1t2NjJi3
vZ4mYhK+PPsZRTdKo6hmSUrrxk/KI6DfruYF4E2LRPUPu4lgyVukGpQa9PBF9xbI
Jl08uREDD5kZZ6fuex/x5D7jUcUFvf9Yd3ZjTJFiAHN1pXw5wL46GOzJyrjAYb7y
YL7JqA/vsEuF9X8Qf2DhSJ9FsUYhn76AwFK5meForEwhMb4V7rjHizQfFyWARwh4
Ov37adTBnFoG23erY23v40YzwQ6HjpGXriknFGlytaQOe1HBGvJA7ah0h8EQLqxC
+Hde0eC74fclAnTTxoz7/yBfvNYtAJuYTbeuJKx4ogWzaSN8RLOR6sswS+Q57ULu
xK+Tsf4mcrvG1Vm6jErYTvS/VNEj7Msb4rLsSM4zIuXfZPWktO3y9THSUP9nhzEH
vv8yBgFQkqyWHX1VEThoVbMq0Tdop4dAmrGS4MVuSs17EYCMEOYQgaG5qoCpV05Q
6o/1XRqnwBgnG7bygX4QdEoLlobuE7uTvkLLCVJ0k3R0Xf/5tDPPYwWAgY4kvHAM
jo316F4eb9essLHew2E5K7jP/vGs80tBuDnJyUhXpm5GUdecG5a98dCcQ1UjgIAv
h59NxQc2P7RykE43nyhamtthy3Fdg3AkDLn9x9TIbDYVs7O1UcgzWNZDPW0bDuum
7Ar1q2gRbW6vA/h09SZhaFdJ32eiIAvUTgPPNj4WltJj5dJQ7XvQT18oEb3hvGB5
1xLwNTbixx+kRrrmFqJLHBKssro15/jHyFcbP9s3b9N3GcP1/VeDOWGlNOGmHcHS
LpprXV9qn4pzQKrT6Q6YBSxKWBbwmj+90rCdi47t6waJw4iS2dSYiKGQ9vwTQ5rT
fMAzMssiutCu3cB4pJjmFJGYtpms3mEayzXitIwDZLiR+cHiz9BcL38dWmKsDVzC
gsz6rfH7hvFCHtjPRVnZLj8LC1P0ySOdKIb57y4yZYTQF/jyrMY06zQxYjZVWhio
gasoGh2nRUoasPRx+PEPGfs+WkU5U25HNgFSzmt3j5ePUTHEgP0ZAqstmPly25uP
ixqP+6V+k1KVRiXO8ZoCAi3tZb20tQzLiSPIPE+lskxD6ZzQ90mLSQZd2o4rZESK
f+UwmklbMdoF8NmQDXpOEwWtQTBOAD0MlTDB7maz0vw8FGvUArEMxAX7n4byt2Ad
Iixfj1ySVteUWK4/EolQZA5JgBFJshaOhI+33pnnmQIjzhic3UQb7rkKAmgQmVgc
XT5q5XK3rGl82fzYV5OoWxjJ3L5QwWlFDVB78O1z3NsN0jk/J8Gh9+gVXzP+F7qN
JKjdQwrzgEQ2jPPeRH0V3RMn5uVPUs0TpMy9w1fw03OYYwLPZPrEZUF9z8+4UdbS
WSnjPulvBPtsPuzv4mC0xMqWHbe2z7MClLrwGrEEFFxvM3M4vyS4Bz9UGadHlulu
/mEC5SW/8uSHLp2s4N3CRSlL1R8jvCX+Kxf5AlkVeVywIzphs8Q07FFoguVSApad
GZoJjGLBK551pgiHPUYMTIXUS1AzpO5BU/3kIs1KJgan9tEr5X56pq/fIhwDgir4
++ObyqZOQ1UV+TqYwTGj/9BFP4p/WW/1OCjaaGFCx2i/z0kLHOY0MonAbNmJKkBq
7faHpVP4nRZbZmkBEOJ4RzvaKpHr5mNbZv2NNaWhr3ZWo2UbyzI+xFGNYVHGLg0j
EEBwjz4HYoMep+HAMqb9ge19puW5XdAi8o7h2hseHExlPBB5g8u75zG1Xg6h+T8c
Pv6HF1gxSwSxZ5XQmUC/mG7uk5MEzq+pY6xejcPW2UU9l3dkG/VoPgyCcRp5L4rG
3xoct+lhEut18eq5ejwaPf8Sd6jLOZuoEgSSdz5Wz2Oa62F7j5uitUBrJQJQk2vt
7Cdrv8AiOW/9IZ6/j2Ufbnskh0TNN1Pnq9dNteqWhJni5zkdcKoq8wlgeca/JHNW
EuJrhrOsVk1Y5mhM9Bt8pFkIvnSs8iHZa0iWByce3M1f46GZnzMjYlbqoxd6JOLg
NVhK4nadhJlXfxkWmCyKHA2wYPhKl3X3SzqTFpWvrKfmh1swUZQZdzf+7Az+4P/F
oWwrBp75yDZTSIH/KXbnfDF1nFtQVmJPgiXGZPGp+ifHMGi4pNxpY2D8tRulYgb4
3bxbDrQLkvP8A2FJ6oBDwxaBQLUJ/0Y5xvmdMYAfj+9LKDyZjTe87IJeaKChBOFi
G3YgkpGREAAUxHczzK+v5WFLXs3lnaCNekc18Bq6D5mFsQVqU5yo8sv0ZWanBEGD
u3377DX+luw8ZQSIz7M2PwTyrFOVTQvu+GVkcPW89YXQda7tBkE2WXh3cvW0Ph4a
6T73Xy1lKb6AHy8GfHygW4rWT/j8IM31YcCu2Ut+RQwq3sUisKAnnKFdFOwljxwZ
PfVfyGIXZJX4Pmhb65WIq+uJsZGJ4Ul4UG0gZWCC1rf1y34tzapA9PaQE1Gr2qp6
0qMWTrl+/4YAW/cxVMpKoAVw6PMm84O9wM0CNIQa+d8hKhHn3pRwB2CiYXkH1Cjt
mHTPqTJU90/TqRo+MEa8Mu0MP5B/UBMUOy8g1EwQeMavtYZA31QFIAKnypXsI1wG
OziMr2BSNK3EzUhwvTcNB7NP3cviE6QQDlcAzEXOA+c8ftf24220STzolwJ72Sxq
T7Ex3oApTC/PA0BZaITiervcV/bETlEJ1Fy27oIWMYjtJLaU6lFWBST2vEvscRl7
Jjkz6gNFbWv+yzgApzYV+bDvI7HHCVSqXbDY7G0K3pRFJR8ije2ipDxtauxOK67C
5scg2HR/del9uxeR5UcGspH1//KN43iooON9F1vcxbt4QIK4x6G5mKE9NmIq5nIG
bT/eFLPCpcxSe9eHS2LMf7I12CFNAOuevJZHfcFOfnuI17wsUwSdjntkgbXqakA3
l9ghlIoVZ3+eyNhm0qYyMP0HiY3ZMVtea6x8G9GJSiAq0gREV9QM2W5Bhreo6BzL
3uDiec9P94//6E6dd8FOCLDnFtgFf80XEYdRF7RchipcFLszum3OWWgI0zWoZbGX
ZvoPaG52rYwZFeNuGCqqwvp1nQXXelo+5oPRBMiOp3tko95IGY9UFARsrVyhtJvl
UauTCYFkKaRlUwvrNIeLzabkgiy68Yc2/6hccbdNT7RHfbuhwu3PKW+Tevsnf7lC
hgbzh1YGoJEKz6O+nmQvlpvAS1QymJtd3XLalTyFACs1/s4dDhR3EXri9UZRZrwS
e9yfYufduMgHPQ0kHSbx6Cg/er8lO5y5gwpmxyxpKbn51e7vTEs86pzERQ+3bNbJ
p4jWEZRqnGwr+kwcqkma0CpalwE8/spKUvjOZuN4flYecnNYuLSngr66yxTKq/oZ
N7/B2VeveRTeETIVsRkhe6/AFYbogHFD19TaK58S+VEnluaB64gmNam+W8LaMawv
iSp9+LYbWqg+k9e+Rc8XyCeExt+kOCTQJJOIkUiTsNtYpDG+Eh1a08N4kHLGFaaa
jbi4GXRWHRYFnQl+LKoL06kFWe3ns5pTV31AFyD43QiKGoR+p17u7YWP45sCLfQO
dWGsWuTQ2wwFmhujqzzG7Ewcrce7HSJvt04JOdmsQXdOYIOqb2uwPgsCKLn1F+NA
3b3H/Xo3Lb5UBp7EF2kyvsqSb5+DJ4DXEEhzn3Ztyfoj1wNXx16U7Y1qnef2OjIg
akFjDYZ0fzRTeSgqzPqj7+ChPxI8dzOz6u3yakJx4muqn9tDQ9Eq+9kyNdwOSDcX
kRGWKnrCmpozI44mezF2JI2L716KJrxvMX467ybbf/1QF8f/raRD/aAT3dYPkR/H
xzJtuFPDJA84B4y6SKIDwOydrGJ0UP4YKEtU6FdEYh818RQMrUiwSeYqzPH+HFCl
JvDDxu4ytg93wcz1+YBNORrs6kE6j07X87kN3x6Y121vlHV9+SgVH+RlyJhi4s2F
qz9QHFIiKVuZgkGPColpxLZSsd3iVJsmsXq7mR0jV1ipAAnovURAeRFC0z15K05B
173Xnx5e9xm/uZlFINQxcRjUwudqT3Cn7BNkCrHpXVC2YJYLmr6wk//ZKgGu4nZ4
V8TRjfdLf1hyRO/8gU849tc7xNSAPk1LYYsiuvbFSKZaglgw8M0enySPT2oF4l79
f4HZ7kdP7eqDW3f9m6C5Lgxo5Jn3hGHq8MHfq4ScIEIIk4PuBmHGpERqhWkhw/uG
EMUpsrOgcp7/P12wem3rnU8KScFa1slk8PtsX2tao0Q5AbKNHgJo4EKfz8ODSWJ6
JvM4OT0gEjV+Qm8PCWWOGXgJoJAh6wiyjuNaLh1ImBgMGP03Yogt9Q2CfHk6epy8
bvczljVvqKOxQjuDWj2jPmpKL5oXXTEoqQq6PLAz3xCfySc8qtsp4NzmtU1aVZbE
Y8SmF1uklKELSdnrJ/zt1vSVXFGyXQO+FBwYzM6xME5Le74x8/hnGUeuJVz2O+xo
mttetFzkpWSCD5d08bvUv8y5ZqxxlR9CEFuf7hphLnsOIddAeh0hmMVOddqAiUMU
jX/gs9uCZI1LL8aSzI7Y5Sr4nlFFG2MsjrK74Ats3OziuTiSY3Ht4uVL794o0P1u
WkQOMqqSVHYi4aD/EfH7UYaPaPBwF1DPePkPEa3nTrdp2TsL9IvgJEThEVVPUsLG
LcPVXUT8b2hy3Qd9UCfFbk9VMSV3E1S4KEh6+TUFEokx6nv0tThSzToBhppLtG8a
qrP8UxMJjQ+aB/GCjh+z92HNMdeLL7ihOxRDebTBJQ0SFhl5ALXgjC/Alggv/zM3
B2e2+UKPU1vJOeb3B9GYFEssIYrD8ut0UE1Fuq3LfSuSHG7ZH088vpGqoSWjz8A/
YOPmC01JQUs3xz43E8JYr1UuBcPl9Kb6GzFEKaGw86PmOB+7GIC75exZuz0LUl6g
6oNIv2q03E736j3QTlZ3cQ6l1oiR1+n4XtAabPROwEOjl55jgzvVLx1Dk2un+37m
xbEP4jFTgmWg2hRBJNKtNVXLWaK21GUBfG9vczfhZmKxrZcokaQEUs5IsY6RBPmh
m3USOvtLptTxdX3JneEL2ReAmUclco6OH4dzltumY0MW9e1DWc8ydggS6cKTXkqh
zU14keHmiGC2uh5QvR8bF87FQwIUgBEf8xcOb127aWvpKeFSoTGghjsFoRSaobwb
8duqcBW3uZQ/8BkMYSGLK7fXZ3he9nxyf1yX7C6yyxocfgLuTZTvG0RNFXWxl/xF
g77Z+oJ9+vDZxT3tCmVCK1sCbHJFvh3c6TjGNxBRqJOp+6C1EDGdFa6aCba5zCns
B6wOlfD10DhXaALBTE8tDrTaTLAC6q6UCVhZQtJW+ObVLiB8IT4CTgDiMsnc5SnZ
C+2n8YnKSqD0B2c3ZvBjupPJjuwxY0Mvcej11/BRm8w0lUaY36q0SCtIBFqe0ATb
YuTUBCrRz35dG0FUm9G9QzJctVHps7pz005P4MCBSCFagGqn5a+XP4/4VXJ5B3DS
Pmf5zmf7Sx/lCLUXuBNN0PSbY/pYatA03vM2oBjIb2zpf8W6Krd0Kp7U25eBX9j+
2MCRnKp8kj3ReNQ3UvM7MtZtpmOw0fH2ayegakBntN+l9Hohbh4Es+EXIXX66OZW
QsBnbuYhBUY3tX3/XoG+zBhTm6YqM7+en1S9180TgaIxQ/3LZabLgYSSujW8PZLt
VbeRZIbE6pGU/nIy1QxGHqwp8LpXL+1eiKRweestGZYW7u4NmDX7vClJiI5+Fi6Z
hWuv2LQSRcui/umqHPfZeN3Wxz4VibkesTyHAAdgWBvxILuXtWP+sbU5eyqeOSbD
0IyTU+ECG3QjT2t3Y3nwCP2tqehb8C5K5TUYKSisNcuez9DuYg2VovUix4AQjMtW
dY16ny+9nanCaQ/kaJ8pH6r+4aV9yHQ7jBHD/QlSNsaKvz4Yqo0wAF4AXSHcAwtq
/rKQA0MsNmad+3zNUc21ds4Ixj0ESuGcP56ONxyWwqdgqEPYI+kvWEGHBpOIjRoZ
w+coYqxQG/xzd346UWyjU0sp7nYV2ol67x3PmrbSiZIODo0129/OrVyMOw+UVNoK
GNu2xkF515Y1ipVXRBmeadJtV/mPivqffFXmuUIFv1hY/sLfumDklHl6Jzwpn0FJ
qqVmlCeqqlGuMyJQd/UBbG1GJa1AbUKhTbnwLM0ec0lk/eNCQRTb3w/G5wgYJ5kS
KEw5g3Q/n9Ne1waC5sYC1eFcxnDy6TYEIvCSryFllO8v3di86WkpQafG6TP4fMJ/
6KyoIgjcn6jIsmW7L4jCzTcnLBG9WY6XAWz1QTeilHO4PNlPIcx4/Ir/xAdC+PAA
rpx9Vndj78cJMeNQOZh2mhkaPEAImG6tpHwIT9HBxMAbRYUMZxZwg7VyQACOoqL1
JgYt6ts/d3Q0/Dv+LeI8ZouLPwhHttaK4P3mbi3Y6mZ1fVT8QmPHFZoaEFfjuE5O
zVc68sDAGe/7QmvqSd73whx+MYyx5sFG7rlsVZJRTsNwp3sxn0OlIZOiT5wdN7t2
2TD4ubsIzAIOrOZfJ2W06ZGuWYK7LAtvwpxUNUDf9nqRSq5XmaHoIV4I1k4ZiJAO
YdakrZxfqqwZo9C7OO9tuGsEyH0bIId8jwi6SHAfZQi0wZnrsrmffDPTht8TFp6b
LHwlLiv+OxXnI9WTb2dr355v+81LBMBmr+0kVkR/JasH7tAcFEAGp48g/YXGq5Wk
OlwtcXthACbWPoeUtWHadwLnkvprC7LWdrC33zwTt7Op8C0ADDELmLxNtQHjR/r4
z9iWQBa8KfXjkPbiMzzPvpaGPy/b9EIvnNk+gjz0CLx7ko44l5K6W66TxwvT3MJ4
g1VsLptu0mqRNbA9RzyweKL8nBMI33ngRDr6UVzyDtsF0zs29l5ofDXn28xbx+bO
ri1lcWEo/JLydN+YZzS/nfLX4nTvfdmVXf1mQphXgdM44jKEN1T3qA88GcoGfOs2
0ynC+MYIByWmUl3VzYoe5tqDgX2dcr+EH1UDxvkVgt2bZo6KlMyQwcMNveCBGYqi
ID2mfpROWAXrJBRcASsvBOfaRnUn6SgPlo6TWg8+hqJHWwyzoyVLr0ksUgJmMKLD
LXjXIREoxOlRgfsJ7T3De26rkjZP/pH8kQDQfdrGJmhKFq/FO64nnieclbX+v4k9
8ilBxEpEWvOFpXpiN/Uq8jIWWKWg4CobCsKGR+XzhYWsgTNjJzNxHYe9JBrH1uYm
UTApYksCOwwBBo7lFPIKz60ETmYRPv2USzUZU+S+m3phR84P2EoNZ0ecuryyHJNh
eTr8oTBhrbO9BCXvdLt43f/MD6r+dgSAHjCCwTRB8haPCHhC69sERYAA35YV//LX
Naslpsc2Y7YeCstzG2t7U764Zfzn2yoo6oaXkaR3uW8vfUB4zPAwKJY4NzfmzUiK
U7szssS/hsBDO8VGW8QsrYeDtmyG6tn5cifmOXDOXDIxp8ajk+FHITK+twbvYZm8
94sEBKNQevOV2FQY6a7jKLYvo+iOlU83kaMKXHt5PFuCO40NMXqNOuiDMSIKkFXK
HrelvmlvVilrv5iaBCggxHFMOy/nokBLPyBs+V1gj4649OQwQ2xV+T87CljZwKKj
baPaXoo8yaBMniPzmkao+mesTJv+DRYmwn5CWnxkhQIjufQa14Z3tAYX5fYOtwJh
4ymxkgsLvf0biFlwEzBmD0HTIvlQojeLTqLdM+7SeRUWFJ4XGF7w7TTLdY5RnDNH
8b8oGp/K7o0b1VMdX5oWCMeVB9IKECbVvzgFFu3LFSIrMsOAvgbk2ZS9ARYbaYG0
1H+qzSim3NcLuoBS/cG/vkKCgDrfWYUJxOJYzhOCuM6BDBqzxB23LM9lyX7F4aHR
nxYrwj8fOQ6cVQGVkJxGeqoV4UzGprmp1U06v18hthICCj6uf/rqGG825pCLxKRR
QLITofqi5Ccni2OkVEWvXnu+FY2PXpYecKjy//VDo1uzf+aRbGOvFZI3++ItiYCB
D3YOwrir7JSib6avtyK36d7L19dguRhOjkbv7k0dJqgpsMPuyOB6D4Gg6oYF6FYr
XBj/wotDEme0zD5Rx93Ta1lGAGnPwIndy1ov+yxGqjZodABfqxVqEBuFew6tDabh
HhTbm6TdOig7PtFLHtaomgOne46cH4TVma3PtgtLVBplv6nTn+OkIOrvsSTY1lAE
GZK/4USiF+UXQjOTzgioG3A7kvIAShs89rE4TOZqM1io9lSiUj05BA4KjnQhDikX
l7TswgjF58JuBIaOx4STBrhQuOZv72OjS4WIPe7+NYX9UUpus8wniuH9Bs+2QRMJ
Rj0arlUglzgrB56opgoVx9aFhK6r5GAIhZ9wnjPl7UTJTTQPeFIPkmsIvs/JAG1d
0dm1cb/EYy+gG6TiWBJAEUWF6VEaZFDWOgpJQRwmWFPOlhU3iapr4GHUtqyJw3Nq
9fy04zNalC+KmIyBfskYP2QkRncDvv6XhgFFjuev1NNWoguzekXz9VAD5XsZuIMd
dkrMV5AeAIF92rnPOTHSVzsN6e6jND7b6TuBEzOHOuajAkAiSFGo5pjpkKEgq6Mq
Hh+WCcfIHXykC3n9SkYHkMiYFjWi/mKaT/lSgMWbjI04QwbjlZMqeLYqsfzR3gcs
S8rDzPvH5P416hdiNxKrj4+DiBs38BC3emJ0JBylaLdON8OCfXq6ilxJArNHQVCB
HmswGcjvprXV4XEnEV6lb1vCRlpKWQYEn63y7xgH/e/NT+60tdNXGjl5RrLV+h/e
rd735w4Lm5idqK+t57rHnnwJBf8wrrgiH2Ggb/r0WH06XT4JXAPXy0U2jMLq5fwT
zNYSmIWkz15nJ4mJnF29ofaumUXvwL1rLlwSKAiIUuSH6YqoI1FNCz1IC1rRwXL8
nGlM7AqpVwOoc9EM6hGjgN0B+6areaKtSJbeNIgR5iIGd7/LI2V33IuA6IBB0odA
rgCAjB9rwksNae1HXOGgxabUFv34afT3noSTz8kd9vnwxt5q7Umx/t8/Wb5dS6/p
c0AKPHocK7l/yKkhj4B6DEVgZYR0/DE6QUWyfYyOZ/paAnXkStpzcrMTu2fuHNBN
qvUlt7BUbuXQExkgPIpS7THctKeurIINHtWd88+a0zeytN9ziAYZHxxi6Ja/S70q
hFEwXvRxxB1E+jpgbRg0WbxqyP21r+hteqZifqbHK4AUkYI/w+LEe8Jpd6F5EYNy
qeE8v7vsRVy1mbBnmPardfpuh5UG/yVsx1qw/RmQoa3AKb22AwXa6J3iXmH3O7gy
TBBcvVvft43iTTFo9R3CYyDa7L8hM2AHL3IY1qs2tZTnPvvTwjd9fQVO8W1L48dc
DsHtV0e7OfGt1m8lCXCWU1/Ma44MMl0MPecEpMqDHFMCSfKmu9knxw8VuabppRfe
3pNiZ9M7N7sO7Xaj1q8vpOtQoecvUnwtRKHcPJxIhE6AxYzUaSppYgQCMB8u+BxF
awvqCMhrYJYFhOImdHMNviIffx4cDcC9FXh7Le7SM0/psCk36/ospFubGrUAwayv
CX2pIZhm7fHWRaS0G3vP45TlIhcyo+1+3A0UDpyLZVGAeqNKxwYFoTi0zQNxBm6G
1fVIO8WbFfGJF/Y6zFx3t0S/wSTXbrkP1Nw7NFPQdkPNgEMC42xHl3tswq5kAxz0
eDA/TdEPyO3p3jNLsPvw8SQzeDRy0Ut7mZlJuun07KcXBN5xIh3KesYqPZ8oTOeu
Y9RCrXT4h3W3KPDnjUNghavOOoCs/Wv0VyC3z0JUXT6vvvS3rVBqF9xTjilycVk8
XTfQMTPWJUDeht3dph+oy7/WipXFaZT5p/qToVIs7IouuKsvaVmFr3ShwiTna/0K
3GVqWZZhbZXIU6GMVrrbaAoEqX7iPQ9OKrcS4MHTdNPU/jQppRcTrLQ2RGq2E2n2
lth4oZqkG2CnnyKctlJpkFZwUYMTVd02CEgfyBXPFfPCo7spI0kXyjknlFjh3s0w
IGy+P6II5zGorgJghnsfjXJVJJAklVBNtiY6FchIRwn8IPQOTq552Bhr75EtrGaX
cNfCI8u5/WBQ4K61/iw1YF3a9hmK9uf3bcguyS5KUpuMdQKYwCbmIPgDf+sCd6QT
OG9GHjluZ/wmrm5RQ/OYdRt4n6uDWNvvfjgsAqlmHXkIsffhOXrBlRbvTK1hrk6T
6sW1gKsVaCVCUjQ40s4fg4Oe2PiV3oo7HFNrIbb+KdlcopVTgyTlN0sDTS14+1pv
24WtSqgKx8iMkMgUvvNSISHpFHLT4RTSSA/ZDT9npkvErqcTXEBDsw8XMXhdu4WY
B0WDqEpWQNnes9uogZzabvV9Z5wJslvimdrtzmRh2UP/AimB1BavGA3g3f0UQAL7
/DnLgb0btFCQRdzzgxFHaURVRtJ6WrdQ/C6sHN/022hikUA1U3m6zSUbRnVM6Uk7
3hXU8U0BmARsLYoMIfM/nQgZvv+0arwoKzee9Pn2Q9UQzMxW6iRzbpCiGBmwKrKJ
c9sNzAdg4LDs/+A988wI2/I7ljrUoiWtb00chA7nRnxcPKIQqEsx4RgOIfLUQ7oZ
eRSsjTm/gcyLxwIPKWymkNjfj2s1MBXr2yyMlIbp2JFEbO2wb2csr3FTWcHiOYE6
jJpyo5+uiZEiiEPWmLSmWf0nb1sFT5moIKvdwF3IHqOwDtXMBYk3JlWCh+c6uCHE
/8FR6BFzMDls3SY7K3arCSkrnRg4eP+eD7ufG1FCFMGn+KWr8f5cBM+S0sO8KHkG
km6WTMifHl8qox+43ts0U8RuOUl4XUY3MlmNj8Jy0ZGopD0Vj8gLsK2a+H0URnhv
0noRu32P6o+gGNhvwUNwEkjSUktadzvg1NhcS9uwDd+FvatUZipqoD6I/Ww0uwME
uiqFGzWFARf/WiSSwoCDaS/3skxHBd0JwKBDp9qLwnLHmmRP4p3aEmBs4IAzWPzd
y0oiRTX0kn1ui5FPLmM1GODZOw375h/ZmtpXpcS5AZUAkLtwHOrqD+31syKaVSI6
VIWTGIPf6fM6Wgvlhf5QJN2UH/JbRemB2QMeh2C5Cn7+84kt2VcSLalvagN+msH7
velf3U/9GKfEASL8ykPn6RZxmLRgy+9g3rZcAJV/2+vulsRVXX5ZLuegrCQ+DCCA
Kwny4GNMFSjP2wEDqkYpATP4t2DrrPpcAKA01goJ3VwG+/JKnu3X1LNhRN+tep6Q
bDcw4w+IdksADho5Ps8sFZcwaNot2oGPv/uqTlyC0/pZj0zcTGhsSDT3kELtGHlo
Re8Q4obx8yefJuf0lSNO/ScxabI0uVOyzay5+zGM1kGKURTj0rRTwSaLTXRdm4Xc
A4Gf34oAwIuW7zOUB1fmUGsijWGDCZpb/IXOVj8rym2HwbTmHInRMAfToMumlrWU
f66q0VilNau3NgddOnx7Je87ijaZbp7cfrIdMuP0ixx2oHpSnX5wfvxC0NxtYcG5
rRsPti65hLJXTvyXpTvL8w==
//pragma protect end_data_block
//pragma protect digest_block
P83QXyROc9GtSvgdl7KxOBgqndE=
//pragma protect end_digest_block
//pragma protect end_protected


`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_master_transaction", svt_axi_port_configuration port_cfg_handle = null);

`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_master_transaction", svt_axi_port_configuration port_cfg_handle = null);

`else
  `svt_vmm_data_new(svt_axi_master_transaction)
    extern function new (vmm_log log = null, svt_axi_port_configuration port_cfg_handle = null);
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
  `svt_data_member_begin(svt_axi_master_transaction)
      `svt_data_member_end(svt_axi_master_transaction)


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode (bit on_off);

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) Tests the validity of the configuration
   * 2) calculate the log_2 of master configs data_width   
   */
  extern function void pre_randomize ();

  //----------------------------------------------------------------------------
  /**
   *   post_randomize does the following
   *   1) Aligns the address to no of Bytes for Exclusive Accesses
   */
  extern function void post_randomize ();

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();
`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Extend the copy method to copy the transaction class fields.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

 `else
  //---------------------------------------------------------------------------
  /**
   * Extend the copy method to take care of the transaction fields and cleanup the exception xact pointers.
   *
   * @param rhs Source object to be copied.
   */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);
`endif
 //----------------------------------------------------------------------------
  /**
   * Extend the svt_post_do_all_do_copy method to cleanup the exception xact pointers.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function void svt_post_do_all_do_copy(`SVT_DATA_BASE_TYPE to);
`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(uvm_object rhs, uvm_comparer comparer);
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(ovm_object rhs, ovm_comparer comparer);
`else
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare ( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );
`endif

`ifdef SVT_VMM_TECHNOLOGY

  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_axi_master_transaction.
   */
  extern virtual function vmm_data do_allocate ();
   
  //----------------------------------------------------------------------------
  /**                         
   * Returns the size (in bytes) required by the byte_pack operation.
   *
   * @param kind This int indicates the type of byte_size being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in a size calculation based on the
   * non-static fields. All other kind values result in a return value of 0.
   */
  extern virtual function int unsigned byte_size (int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset, based on the
   * requested byte_pack kind.
   *
   * @param bytes Buffer that will contain the packed bytes at the end of the operation.
   * @param offset Offset into bytes where the packing is to begin.
   * @param kind This int indicates the type of byte_pack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being packed and the return of an integer indicating the number of
   * packed bytes. All other kind values result in no change to the buffer contents, and a
   * return value of 0.
   */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1);
  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset, based on
   * the requested byte_unpack kind.
   *
   * @param bytes Buffer containing the bytes to be unpacked.
   * @param offset Offset into bytes where the unpacking is to begin.
   * @param len Number of bytes to be unpacked.
   * @param kind This int indicates the type of byte_unpack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being unpacked and the return of an integer indicating the number of
   * unpacked bytes. All other kind values result in no change to the exception contents,
   * and a return value of 0.
   */
  extern virtual function int unsigned do_byte_unpack (const ref logic [7:0] bytes[], input int unsigned  offset = 0, input int len = -1, input int kind = -1);
`endif // SVT_UVM_TECHNOLOGY


  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>read</i> access to public data members of this class.
   */
  extern virtual function bit get_prop_val (string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val (string prop_name, bit [1023:0] prop_val, int array_ix);

// ---------------------------------------------------------------------------
  /**
   * This method returns PA object which contains the PA header information for XML or FSDB.
   *
   * @param uid Optional string indicating the unique identification value for object. If not 
   * provided uses the 'get_uid()' method  to retrieve the value. 
   * @param typ Optional string indicating the 'type' of the object. If not provided
   * uses the type name for the class.
   * @param parent_uid Optional string indicating the UID of the object's parent. If not provided
   * the method assumes there is no parent.
   * @param channel Optional string indicating an object channel. If not provided
   * the method assumes there is no channel.
   *
   * @return The requested object block description.
   */
  extern virtual function svt_pa_object_data get_pa_obj_data(string uid = "", string typ = "", string parent_uid = "", string channel = "" );

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB.  The pattern is customized to contain only the fields necessary for
   * the application and tranaction type.
   * 
   * Note:
   * As a performance enhancement, property values in the pattern are pre-populated when
   * the pattern is created.  This allows the FSDB writer infrastructure to skip the
   * get_prop_val_via_pattern step.
   *
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
  extern virtual function svt_pattern allocate_xml_pattern();

//---------------------------------------------------------------------------------

  /**
   * This method allocates a pattern containing svt_pattern_data instances for
   * all of the primitive data fields in the object. The svt_pattern_data::name
   * is set to the corresponding field name, the svt_pattern_data::value is set
   * to 0.
   *
   * @return An svt_pattern instance containing entries for all of the data fields.
   */
 extern virtual function svt_pattern do_allocate_pattern ();
  
  /** 
   * Does a basic validation of this transaction object 
   */
  extern virtual function bit do_is_valid (bit silent = 0, int kind = RELEVANT);
//-------------------------------------------------------------------------------

  `ifdef SVT_AXI_QVN_ENABLE
  /**
    * Returns index of qos_upgrade_delay queue which matches with
    * current cycle number provided. If it doesn't match then this
    * function returns -1, indicating current cycle is not suitable
    * to upgrade QOS value. 
    * If there is a match that means current cycle is suitable to
    * upgrade QOS value.
    */
  //extern virtual function int qvn_qos_upgrade_index(int cycle_num);

  `endif

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Mycc1KOal4XStkyz2V8TbJknUXyM96KJ1lpMQ/rtuVjLBWhfLhXSRVBFOWxSwa6r
eYpZdTu+vOLZ5LO7jw0GC4OX4UjdWG7JTqRwcjFfBmC8aHVyztaXLyUjJ/vbF4lA
g8jdD6pf7iT5a4+Y1mKv2X01H6gDOlTmkxGM0BQdpK+ucbYeTBbP7g==
//pragma protect end_key_block
//pragma protect digest_block
RMqDKKsIBW5+qEyQXaUAwonDIe4=
//pragma protect end_digest_block
//pragma protect data_block
is+mfep3W3q8imD8RLei0IrbXrY+E1LORulElJQGY17uUQ9geEJhDmJTRlnk3nbC
+83HdZeXPsM/Ly/0KUQopEuijFhIn17bx8KA9zIlZCgwqDgIiHLvTizLTZbgea2F
BaVii1XUgpaeP5IeXMG9gYFRzoDputSatZjy9USaW+/hd/3r+OqkBcS1VvDPmR1O
bJarM9dLLdcQyyWBEprme66cO+fbf6fGmey0pqhHiDXTt/aw/VhczCNPF9TnID4I
JDtN0J2TbaXbZKaxNFjRvdaXfLL+feOajGG0AAibCLNHX7ReXKXbS9KWaPp6OWgR
/wGXMlvpJ2aNNgmzz2Efk9gSxXXiGvI7Z0wl1Qu6eMLFPrk3LXdTYgRfC6rOTIrx

//pragma protect end_data_block
//pragma protect digest_block
pONe8ILqP5r2/IheGl5aACO66/I=
//pragma protect end_digest_block
//pragma protect end_protected
`ifdef SVT_VMM_TECHNOLOGY
     `vmm_class_factory(svt_axi_master_transaction)      
`endif   
endclass

/**
Utility methods definition of  svt_axi_master_transaction class
*/


//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
7UyJTC6gqw7RAZfDQXtJMRS98+NVeYIKkaeHVY1UpEOFa2p30hTdp+EL+8rRuWA5
Ne4+bDHus3Jt/Q64uK5dHAfjVb7mLOb760VI4pWn5JwY7RYcFgeIMlWvj3k0j7ht
H7GKAQ7mehsYUXjros1ALnCIDez6yEduPsozl4vBwJiGg8hE8fY8Wg==
//pragma protect end_key_block
//pragma protect digest_block
BWFKw2YUQLVlaueZxL3PiqOH2hY=
//pragma protect end_digest_block
//pragma protect data_block
9NyIY//Y+xTTTC5SVhTBp+l/IbYBu31KWUT2TML+4JgO/6xxCxMxe/yFfTb3a90f
wDqwbCyZrKZxEw61arlTOhP3luWwV8ufneS+IApOEXYWneUdVU6xYTQRKRrcpk4O
DQVumFmDiEleera/vvKQyo8HtN/ZXUyaNIX4hrTGt1VtU14loLNJpg2fiOEcJbTV
eDmA35H4OxewSIHovAKfiKjCWaxh06IAwO0gYMiw6JMgXYHsoW4O90PjHmQHnOVs
IUcGZY5eZGq32W/qfDHLqFBidstOa/NR/vVXBK9NhZL44nWd7ec0/56nxEDwU97o
VONCSX38qniAQKJCmsKaApF88yJeopOi/ndT89AMv1sI3q0iamUAdDEBatTtd171
/DfGeq3XrnelrQP+ZHzkaOjAX+gnke9t3k8lCuaWlhOXWzKJ7JX27fj5ttw9qImm
YKeLPZMVAlJDJ30adtlHug5E2hkmKFcjBcetuG81u9KJ+5qRLFO+BzD800v+98NW
0pxGBVC/MIyGqDxBcT+gvmpZ2rG7VdKofznhzmlVCCVCpqqQInxEJxKgH4UfaK+t
Ppj+Y7pxdPjppSqGI6IFhtq2xe5bsPSQOQ5aamsXvT3OrFjCristRwgOkFinvzvp
KoLtZhd+cqg4lmJr/09r4bl/+SiiyDvOKvDXSr1WI7T4snxKuhyjXLS0BQ0rjrmq
xv9jhCaL3c//t7wxYmMvHD8CFxyQF1YQFe4EdmVRy2xBv/l4NJHKBBRZ9jR2hnT6
HYp3dknVgkkL+IwCxhHb2AakcJI/UcUZc4DIlRfYdcnwYjfpFHU1x2kr07+rYFj1
XIBNJemYEIfNYEkyXZoTYjRzMVPI0MXG8Y8xJeGUwgX8P9p8SZnmTpbsnTm5lS70
acLDab7xYBeC4eJLXvFBzO/dzMaEfovPKFuBmwXrdj15TgpbGGauq7jSVnHfqupk
X24XAoPmO+zKctq9HDTai0i57B4MgIKy75gEYOwLwTXtBpOrT87VQ1h/sNWynDGU
PU9/yH5pfE2IfkrZuLDHXMiTc+Ybh4rIuZcV8h6lHwsUn73Dqjjlkmpuk1Kw5h07
mDMYYsXzpiUnMSId5PFIToB5QyMcvifO/4QtNEOyS67Prxcww9ddqEmda2oPF8t6
rKCAFwP4PhoPvU1AG8RMYu6WnsCl/VKjzbVB7z9gJ+47LdDq2eMYoc+W7SKblaR0
4PBFZhr9QV1t6+3J0FE1ImJWGeqimR9kwp6atJ8PvFBleL825V/pKiCNMvnWfM/s
ukuxkDbfhDEUiI4UYbbnbPQd57x1dH31iQT9MWHYUt2XyLL7N1ESJYKbTmTUxQVe
Mk4G3E9VLzx/TWtCDPad8/P0QuOIT1QBdhVLd/4BI/+Mm0Bkfn4wSUKYsai0hdi3
0nLj8SCoLt0izDu7w2dlaYlf+e4RN/DnSqC2jaHcanuUnZgLTRbo68xpA54xRJHw
DU5zWfRE0eoatk3VDCyxfDQqA7Sb70bGhTJ6xejlZMAswyaEUx/OEwJwgoZ4UdhZ
Zmqg0kRwuGdfjkI9avdSmJFW6IS2OwjZ1HaK91jlHF1lruWaKUr2pHxhypc9YKFT
axaddwGdt0MSpIvv57CdY5o5zzoRotExupBcpIvMzGPNDzu6ZKE7FvPmcJ3ZVTix
gKewzSp1N8w/x720wMV7QJR4F/eoXnwW1+a6MKLnZzIpT1IKiSjlcLKsSwXQR32m
yZmPxImOMhdjmreYkKpfKS1QXVO+xfa0gHcP0pVkuekyQyQppB0VRG4tzcYHI2EL
6RW9qG6HtuPlZ158XZjsUEoG9gEUgguUvECevVi1a9O0r6QZZYxBiH+t0KiAjXx+
n1UKuMnTLLh17ZllE/RZldB/bVSqk51souS8vlPwm/fxgpC9gtvTMUXoDuzh4tb7
1Y7svxlo3ZEW7zCQjdaqQSORUfB8MlboXGWR+b6qJHkfG39bYbrYYGsCV6ziIIGJ
S04xNYCvF/aL5+T8Jcr1FWgbLjT7KChICkNc4eugT/m85R9Lzr1SRNpfimCsFBEF
P1yocu2NQDzxgWdSQBLGsc7ZQv9BkxhXi5MtWKu7KuYuCbzdqlqiM4RGLCSY2ENj
mN2GA7PgxPeAogUaQeyHJ2dTMjndquON4WgaGxyeL8i7lQ3nHDLqeJA4IcUWFrV3
P41wbpLBnU92VsErP5CYQTpaf6RVL7/j/iZZDn2sBzoybmgoEeDp+j/1xw/E+Qfr
czUF4THtYsSFOux/kYuz5th4NUKsFJzbUZ2HhOo86X58Tk0U+QvioJRVj4bZbyud
6VY+DFbOpqAqJcoM2EWH4zV57+TrC1gL2B7Y2IkR6XMpqfS6Ap95p7H9mDROq6mB
Al8NZ8OOdyv2Iq0nJ88Ts0xyG6qZS8x2xGEV/sEzdzKhBfcOZKVA6QdT9YkWYBVA
V4vYKbZWbqggjMTRxUo9qGwYzm7pZl7RocpjoitNPmweWhiGnfKnYxXNRqDdbJXl
Xjcu8aHNnyyxuz6fYgDR3FzapW4tLI0z1wZKqs7fu+8DotX0ZWMN8s2WRzUNIjuc
d/T8xe4Hln+EU5PzXj67+hl6CTICoQNqR6ee0Qpy4TPrf5yBMl1C9F9mNVrrGXAU

//pragma protect end_data_block
//pragma protect digest_block
+u5HwcmYiIAMOFHOmUyIFoHB1Io=
//pragma protect end_digest_block
//pragma protect end_protected

function void svt_axi_master_transaction::pre_randomize ();
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
bjVxmb0huX4Rov3ChP/h3/O69j0DSuM3iM3OKSv5wFOXLK/QDYWTiC3R4hbtbptr
hvZEa8mf0HOvAGPnNrS0qW05RMpnA8YHyR5fDr8zY8QoppFPmKvmsVbhEVSrUatz
3drNJUxp5hZOqzgO5fZxitsuUkYecILUvv0Otkn8QxpvvryVUGF85w==
//pragma protect end_key_block
//pragma protect digest_block
XQfZe2F2KLt9uHICDppEIwlF9sE=
//pragma protect end_digest_block
//pragma protect data_block
1QQ8Zl9rC99XReoxZhYAEWmY29Tgubz5uXy/zlIFLZeNsr2+z/6cG1yhGRmtilGu
ZKyRmHN1OBYthdnZz+DQxmm0TC7Ip7aSKohVezCcEKOw5XI7uoqrT0iTO3rHdi6B
izqf8J3Ge1XBJ0QUMZhJWdtYjeR1zQx+G4yTaRGgRtdfU9mdm/wLSxJsLYEFSPWP
MhVb2V5bheaG71j0twXnOVXnJv41e65H3vKN1+gdsMLEyRMSPgL8Bvju7dKjT2v+
UUhVbOdU1zJYwvYHlWTigHBPMbziabe4uR6kLC4s11xGVOv+V+VoIY2HBbmEToT8
TJTDcrYFrwdx2SduMUSjwdKGY7+LPt/VpEtFuXFKH/Gy98YmDjJ4TslUXcCfF9dx
iQ+xgCyyBB8Q3Jmme3t0WnWFO1YDwarZU9VyPFzOujH3oEYI8bvEY5sW3tbhqTOo
h9MpwLrnWBQOv9Du63w/4+E6462XnocwnaYrlGGdBLzKtyMnSIkIoNhg38viff+7
Vt7/mueSyVbFYlGkbL/DxlIKKLif+Z6gpYm1zS+ZDIgflWwMWQE+JB6CQyaAzm/R
cd+4ib/MeIKP+A1B4qAtdofOr9KCHvC4QJ8Tt/TTYtFeR1qo12HcPfZK+4/Ud7hV
ouVP+vw1CeFgNqep1n1sph0BZKw4iZF0pRBLtXiKFrlfi8SCln3oEZwVV+2ztQXs
MZMrok6kQdMc7oGD2ADPVamiIdHDwfj3FltACRWNcqT4zxUxLdtT0R77oWfP+J6S
z7vxs1glGItj+8IEM+MwvSzB2znl9tcXgF+rnMh9zVoV52y1ZeQjEvL1ikeeKMVB
z2Y/7Wm58acWPNYM/JroeT+DAoIYXAQA3ekY2+qBTXbl+D1JzNT7lXVmvAWl4b+k
ZJaPQx6+2RKrD0CbB4VyINQgVUEPBRRLtsQ3pdkI0grQcZnvDbhebzeQ3y3T5gu4
TDsNZgnIhiAI3SDscPY6hNCEJW9+vLRulP5hBDe6tw88pJgaNylCmwdfZJMdYIPn
jVgt20quseMM94BgLyvVKwo9NkQjk8wnDnjUM6t7iQpM39ZDsUpz24axHpo3byp8
gBAVGMP54dvaUQTvM4I5S+fhWj3yxdXCG7pWFC8JnslOqpdFOwietwqmDmDEsM0M
LhU3P35998v543+x70RNqCTroKfzin8Iw8buOiwaVJlqi3VxDdbjJn1sp1bWZnvK
wBtT1HRp35ihFZIFYLvSnK4R4NRGPtxsUo4iWfwtDz0TCbN527CTDH5Eb2n6g3Gy
00yjcfTE1yTS1O1JgfzTFAo1/l9o1RTw3ihQEQtFm3v4xtBDtys2pUWe7ASQ1oQ9
vBwp34QaDzIZKHkW/pm01fvqyZfHb1RC5fzYcv2E1wd5RDqG7mXoUZFRWmcIAciP
RyKesKl8/7npn77YIHaf3gyYsY0t+zXfszfxejJzZMwZh25X2TPT8ejnI4Uk50Dq
6pAJeyCQASp03+USjMYc78oJSnO87bHkiUgm1FL+DfGAMQhs51dFZnW7VfkZnMp2
DLHHbMtyu+H65SDjs74uO7hKT1+uCkh02zDum5h4/Ig5jyjnFRlcxs32MAIODQNE
XdOU+qx4TO3KPyzWpdjiRxWPyThUgd4go1HmiY0QRpsETKFx0xyLRFq9SQ93SMae
rd4C1WyAUOxfuptg6ijdRLo/Z0dLIkts7Q4AsKsyabZS0F1RDEnT6vt2XuhGUwvi
DAGkZY1ij6BrcYrUKusYzfu0+tOAKzgVwRNDFt7c8XuTEPOGPijjxWMBEs1q05Ud
PCHfCxan2D2oOTzZNiC2P+kQN3ZxEtnldGwn6qSWdPz2hfoZ7mGSBIW149i7RXPN
GtRuP4zTcNOreyacdqFuTToeBhw8fRdbh64z4FUe0gPCqI2DD/O6Wbw9Xp0wxNhO
TvjuV6gHunQZ7cgpaLBrOESLitO8J9MZ3UVpXt629xZveWR9ogajaeTueqG8L5rj
1htgX89QiAjQrL6duosYx9rflhsKLKMAWQ4gU5j3DTGlLP4ovzzmdTlOck+zKDwq
FFOAyphRKA5Pf++WgHEpvcvpHOlbziiAbaF20lMy9iQQXA3LMU7nu5+0sX04EK1V
p35Xu5cIiL2CUc2ghL4m0hMK1aGCqWsoZ1DdAVElpUv0uQO7uN8eQUeyoDjoSWJz
RUi3qAMSbRFi7uJd+kB9Ue8mbH2xjThSnWsVRX0ojIyso+cXlnKHtMm49W3MMMCF
kE73P+lCgb+hRFHIQruiA2ZvcQdda2PulUVsekwO7qRgZtFFN5ss3TxeTE+3EuG3
EH6ixDWKJg6qZkEuGkNeF+IHWrrHHBSoOXILi3CxnJaZLfmd3aEMgRixhLKCPV9H
/4MG8yMjRW23PjN4LrsTKyy4IsKXAy4nUbl9L7/w/7R7WvF6mDgi2qeMqysC90pO
qgJToW7L7mdt2tuajI+/FxFfOkKoL9USQtkqrgVVsZhDfIhymxqvRYdDGTec1d5J
FziF2EpBdIhj2G3Xk/heNW0Kplv/OmuokHPQJh3iExnqnpYqjVt+B1+iICZZDwEv
yfUOIFG307+Uoj1EyuEPIGsikSCWDkZ2ZJKsSY9DDYReGAiCwh3b8uIdol8tiqob
er52w/s44dRaBOV5No4PIjni7KjqcHlq3HZRcRVXZr0r2EYqkYSxsAwdgDBzBNvI
mbfzwRXKQG+E09lDrpFfhEaCdnx6BRac1sBjdHnMjHnY2MKRQaFOsUu9TCOa/i5v
Gp0N+1o7Sr1xG5OpTcXdJEpbw7g5IbWzNdPxdUGjuye5Rnh7uw14G9Unu+9BKSPP
LTrTeqmpVm8XCmVVDNIHVdKvtAtujmrlLU9cie38UxpBXUz/puLJxNPliQGzVIzH
B3hHpIwSW+lIB64A3APZHT5srx7sBt//gTSCt+86xto5keH5D1ELeDqr0CanqHLD
d1aUbT8yAhnk0GjBG5YGaItpyTKt/1H7hgKJzSFzbAvNBtoRfRsVbEnTLAZhagut
YCCBVDtu9reYJI9SzrZp/M/bUr1Vht7JfTTHTsloUnRAbxOdFJh0mQDrvIPl3Eoi
bgha9rwoOd9MKS48sEObypIWUsOU/pkMrLA3r+2Q6mHM2y//x/2ahd8qhKQfw/vD
VWW8J8g5WjUv5pBBB85QKJQGGAv0u+OjmTViu+PCS5lqJwrOXGCGiTo+CU4p75jq
vMNnGQSCF1NWq936BGlGJ0K55DP7g3hoB0pKJfn/GVK+4AqkD/g416shK7xX729A
p5iQXJyS26aaqL/xkTLYdCxdwilWIkLAtt90LsgREhi1SQ5iw3i4Wfb9pPO+Jetd
aANq9aXeibX7B2EGz8O20zJAZZHowsDFsRmkEZY10uaSYkk3hrUj8nnF3q43MSMD
fKj0ZAU99nBkrVyyeeJjPZ2SzJd3m307dKO/RcmGTiQaIGPPMhTcIXenpmhEKAPP
5CkOHpB2N+PHFqRRbU931YD3yaMpKlz7b+/sH5gmpKcfFvUVw8zG1/V/rBBX6L2Z
HcGNyvFWBpWUWUQ1M2wiAw==
//pragma protect end_data_block
//pragma protect digest_block
8P0RdOfkebLfHYxuIatlLJCSKaI=
//pragma protect end_digest_block
//pragma protect end_protected
endfunction: pre_randomize
// -----------------------------------------------------------------------------
function void svt_axi_master_transaction::post_randomize ();
  int log_base_2_total_bytes;
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
WOmkUBOzMAAwbsMqxlHwSbVLEOp6zf4awflU7bi7Mt059+Vj60Y4s5hbSJmhYVDg
Mm4h5p9ojpWEqNniV7PgAPu59ZlGIACfsg8gXly9M+fnah2GrG+HXt4jBsPftxBt
LFauBHz9HzLGPZ0nhrTIm8UkMmC8pARF5ZW+kIGKgHdS/ti4S6625g==
//pragma protect end_key_block
//pragma protect digest_block
P8O1rpHixsMN+jvgiOlYcVqtSjc=
//pragma protect end_digest_block
//pragma protect data_block
jZWSxF9WzMeLMRAXC6jZ0VhPyUvQRz9OZByDEFyU7aOO5LdEA3GoIRTQOwzJK906
pfK+1FED5znUVKsqXbDdpezAcfQ5nNifsrg0uMWJ7cYMau5aAoWLdMgxRGVOctoj
9W6awA0gCCUI53hfWwyiesEWywA+L8x+azn66sF78j+87NI99T1n5CSXzTF1efHR
0xsdKxBzzcuPaBqfTrSTKYsYr2ZiGWawKV+CGuMSbv9THxtUU4iL6hrDP1t01tFi
Vcs4BbsWLRu0/QPtcLyIgb77rrlMfqLR+loVbt7BP9Q0mDSQkuig217Q9B6WWtSV
hBALAjLLDL6e3tcNmpxtQVaSDGehwyqccZqcNSXkymHlK1szJlqc3m8rvVW2aczi
0w7M7mFg0AUim1Fi0HslxBbW4ipms2xcwtpG7oYwU2vdXT6ku/6beae8Y5GnlZT/
HesMf7yv7EYQYJVccQGMJMQRC4FfPd2VUOV+fz+jXCIK1dPXXlhkgYHAZB2CQwfk
xdxnOhhlGYyRIQDKDLxzlxBK2PwUn+Y0zVHGhSPE0wwqOoym6SuKcxbr8qPy5C3V
LolqQb6sAPBtFw1H7Z5yAIPS6rWmIEfiTqfGcrHJ45wdub06VRWmoiKam6RPXuLO
xQb9n0zMFUPFqpS3j6Vx/pW1fuH3NTnCSTBbfQU5/mW9gwDXvUwVW/LSbysRs39k
IU3161q/CsGrk7gR7dyXPXIhG4/43lFb2XgzzAs1e2UfXVxCmfiv8t0CgLU/qfvt
KSHI4II1yXw+l3mF+sb+Y9QGgx1mK9SYD+a8ne85/90Cvehl38yM4p6C68yo7kE1
Us31bRTNvOdJ5Y1+xNzrJwMXLShWoRK5juyhJ2bFc22o2o1cLByt6psUCkg2jVy2
UvAv3Ib8vHIINp08F0u43e3OtTKdac1/m/K7YLVA+HEjVegx0juIBVG/0npTXZO8
A3ZfqVxvgz4Xzb2vctIJ2Gvt8CBN/mSEN1yPYbQ0DQFCz/evw9c4WPPH8AtLJBEc
qP1tmQnvBRg/+KVnzQITl8QW78v/EQVTKbB1A/6u+Ov/rzVitYJaJ8ejXyOptN8w
Hju9tWFFlR2KtZatQlyr2ZEI5H0TcxbXkgK+t9J9uIb766ceKhxNWdL2E1CDB4RZ
73t2miS3ECj9I7vmsdIkJyhRiI/c9WTlIlLyWHNewUnpeSuK61gJz0OUu1jsULP7
bl+3MPwgK8ngs1T8fKpNwA==
//pragma protect end_data_block
//pragma protect digest_block
NFvRRDhthQq0q873LnCr62Lot3Y=
//pragma protect end_digest_block
//pragma protect end_protected
endfunction: post_randomize

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
TkaG9M+uB4MQwYZEheYEabexVDxN5u/vIQLpAXPqjrJUDqxe5T9bTMNsfJbaJK+5
165RfXUXZiidEIRcAHVYrNKNdr/ZFpvso5xIQfd0/PGkd6s+iPpC2qhfzDi1C2AU
tz2h89G+UUfm8XLszCvLlL3Lcph4VRW6VzAxRzE5yiQu41Msfm8wEw==
//pragma protect end_key_block
//pragma protect digest_block
bnYYgDjEPEJujWFpSTIv6P2KwhU=
//pragma protect end_digest_block
//pragma protect data_block
Nwd3BAdqjYvWmidqYmO/daDdarxuTOZbcHXSTcq9H5k/L3p5h3w8oZaoWq2cNCkF
GlUAglQGvwKXjeJcoq20Lxd7DH0uEQshTqk+E2rcm5n7TZw58FVabO5tJ08B+LAc
ofG88Y0zv2cIwanWf4HoRl+p9kO0OuqGXPoPvHYmy7kL7i5G1KyAPLw8QCjCxYQj
XUt3WQOv9EjC+cI/mZ9DHI6nIwJa6npLkxo54EQyTx8F/udRnLEbEAMe7zTkYic8
K+l6Svb3o7ZCuufswgxY87Woebd4Q11koel+KW9r5z8bSyKWV78E2IxxmL7NI0fw
mUpW5WWsHfGpHbK9AyfTdCqL4njDFTz1kdHKg/GSGC7O8hWzvo4tVGbvcB34Sa63
lsWuxIKnVdb5duE6UNLDBJ1W7DpFIxq0ffa3079LBLRcn5vhJav+LQlKQq3bJc/q
v0qswi/eyG9dvxbVEuZSuqkkZ3J2VzT77Ai32FSnKKeu0PFw7QJwbROB6kFQmoAP
iIfzXMuDNUhnK4YEOm0zMwIVjaCQjZ95ZUgJhz1S5smyNC79B/f3N0JWmA7+3HmM
PBlUBIPW4isvDViJpn4htQVqgpPMmgLp26p7SH+mgp8lMipQR3lDDDE/nTOvvtcQ
23eO76yjBrDwa3XP9XuR3WW21pC7swOCPPSq3HjbLg2MFWcuG6s+WSv/uduew/mM
ViO/zXRnuQfCiiPElZgauMuvEHDYmuAf89ZFzxlcBDFuXNYrWcBjLvUQBGYyPj0g
nneOoKBPE65hoTD7s5i0mZipGQ4uX56s8l2qx/2e7o5eSOhTyk0zuEY7XnKWGCZH
TeA5nqpw90bCh89GVOm2WbF0WvjiWX5HH1PEIxFRA5qNCb0H3WDBGqrVQ/x6pLtR
d0I6PmvqLVxyaZDSfWBXnbO/WthRkdnDt4XsSBIIIw/47Vrs3jbmOcno4M82yc6M
7dJuiw+ATdgkziemgX3FU1vcdZdNXqYg6bK0hu9TJYDRi7g+XQuoOroJNUYBsPp5
asxYaiCKa+7ZhCZmV183I4JvCNxFvR+rg+tMe1Ozl1Q=
//pragma protect end_data_block
//pragma protect digest_block
IC3b2YjTaYlWl0gxJtv6pk02yQs=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
RX3PFVJZHt+dXxgJefuSOWu2yfJhXD8dAx4K45E2YpX9B24VXex+j+vFntb2Z0qh
li1EYo5vcyiSaIMNVi3MdBBt4Bd6AQCkTCoyxm/CIfZ4jTRImWWVRK9B3QubrCuY
fb9DA67n/BwbQM2f2MRcj4hjCgrAPG5fkfIWKa5sz5LyKZjjo5MylQ==
//pragma protect end_key_block
//pragma protect digest_block
8kso+uOraq6rowwcR77zPx19Mso=
//pragma protect end_digest_block
//pragma protect data_block
yFhy2BdHyoqkGJu5dM9L+ZuNtoh7MmRBxkGuo6XRZTZttr+zTOv3XqSkCsJTs1vR
FBFlh80DJk2bqwTLIOeg4rvDowiskgSUcvEr70yx9cnAFqFOrQmMv35DFg4bAaFu
O3D3fx0jxv1JZrpYo2y1CW4eKsPxXElpid8F4ZFlFChbEohrW+Aj1tPwAFkP2na5
8NqA56kYUQJGWTqB/HCdJA6lPR1SsbXMrJdbZ6YDVFhKn+8sdxv9Rd4gKB69QAp7
7eOe4bP3bpjuhsISKv6Yj079URZVsvjq33Y5KoTfGFwgpQCaQ/dGhMpJDAU+N2r7
txTJXxGAiHZs+VZ7oRn4UG7ppIBiAfy8fxNWn1Q15YA=
//pragma protect end_data_block
//pragma protect digest_block
TrKBt8fTyftBMoKItj52ue8udu4=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
uY88Nr+7hpvdHW6zwUg+7W2lxDwpDZUyJd4ckvo0Htr7a2pNDign4j3eQbNPZdQB
yoamQgy9zzwrVNz9AHVkmT59vpMNrimVZaqmshEB2xhSGxM6BgXOsXN3REVELaJQ
gjm4JPwpo6JGc91hjfZIOG6brLElhhvmDNyt27KTYT0BsVK/YYuIvg==
//pragma protect end_key_block
//pragma protect digest_block
U0VqyVv0sNjm05LBkjlWl4wU214=
//pragma protect end_digest_block
//pragma protect data_block
Cu2BeW0wa3q8PTBCY/zMtyxsiw7czdP9CGkbnPExWdpC1vdY4Y2gB3lrkV6iZZjo
LR39ODyAdq6+VzRCbapRMZO0eGFCqqNYoUCUdn3FL/7bcZzzVMdRwRzjJOgn4O3q
saA4vxs+aQJGTE3s4njEbxunojzENhYW4xRSFtyFcMZTcBHECS3j+xRQdt9tli4E
ixXiBdHuOZ0UdcrR4Vmt/aTYSRV5U+hYEO4H7iXOUSoa428iXqB4eZY4/oBJJ1mi
1CpBVgZIgNMVh8anyNdNSvDJtLdRZsU9/N6E75bkXydv+w81NKzJFj/NJJhGTMVx
HRUBe90cx3YS/NQGJ0WRPjuW+g47as/n5EH7QQW0nYj1dSYZeU4okBFWN8QH9fIL
Z/9IWRqCvaWyshgYJHuWNHUh0wEevy2z1YFre4VDyxqs2yWijFjoM5+II1ehq/Br
MFzZdpgX3L54vOk/iaOBVsZOglh8ua12Cxahy2jlC1Vj8FLLeLDxiOmV7nAGSa9m
TAjQBKREjvK5nGSnOVNKWCzytPevCZu8ooN2SL0gOfb3ZjMBVdzpOCNhHKZQiVSy
9LUWs1SxG81GzZlkoZ9g/cqkONqcY2mRxztjIqQ/8mshUFtbop8cg6IGwSiB1Q4M
61eGTB/tS/7fbwQ7Y2+Ue50GT6Cz3shCI5B2xSz2K8M8bd+jyHdqArLERXEa6/mf
eY4o71T4rRG708IUByEvzmuGhlQfpLFtszwI3tOUh6FWp7o2BQpx+2QyOz+JO+rY
sHIoo0Nt8Niy/Mft4Rb1DJOSdbvasvDHCg1wLKx71SOgxrWttQkyPaWbSxnUJrBW
Hm7useZlz+gtMctdElyhL7fSOpwMt0/Xb7m0Rf26ujC2DF2ZTey1rJwdF370WT73
eGfhlmM+HA+RSIv6t1kf22+oXUUimC4F9hzvvmZQ40KmTAF/nXGz0Kd3TN+NVNSD
4z7gfW+4/qmvscjrW4go8w4knUCESFXFbPxZy0urmlVFiaZx3S7+YQVqPqfjKIj+
C1dbpOp8inAKEj9YGX/uO5Vq7lTYYARnW2gSecuzjfuTG4rC8SgjGEmaDtmIH1gf
ToqKEiHV9Qc2bf8MIDTzcXlLzOU3ZKysQdDvB1JuAYWj9DFcMpFC301wofxsqxMg
hTnUVu7H9H5ZOhQyS8WiNC709yB3mJKzbOKpUUTunkYmCNK/4vcPwO3E1pLqUxsq
5vZlANWuXWuIDvYKndmr+4pz7n+QlSt5TtJqIoKkkiO5sXVm48CjwQzOZuuEc4y/
QsDD9GLwryDP+9uVmuNFUsT9jHMRQKCYKuvAS0g1nntJj2g/pys7OcWOIxsQTdDn
0+8TZyumfeSmRYBDj+a4GXtxaHeB8Qv1sI4KqcHrQzVuqPok1tC+LYAG4/bjXs0f
C4k7gWpq2jajyoejjyzzSjnsbKMa34mjrNasnAXKZcGnNpiMSuQfbh1lVUBNvQgl
uJQTbOZalHiPUjig4yZeZ2iL0ugh8GfvILZRby8LBdwLmL+1PZoJQXpTDHufVUUK
ntQClp3U8zlgFJzmdBoQCazhHQ1v4nKO6ujTQilvrmJqEeJbkte+LtMdJbreyraB
LA3ECRldOIOg+AEENLOmhvqI9F7SXEqgJ/+2WTponL3uTK5G+eS21YnXr+35gTZz
NS13ofQJOoiaHdfMy3KAigUtJv+0cwoz/PkeqwpPgzmex2kBKT9DydvOs1s/tq42
1IfVRzenrdgbdfzzY6aBuVCeSXqSVGmPE7jZ2lc/+Bna+gEFMOnFi0ipihaVACke
rYRtFZvqFKfSNpJuQ2eUsZwi2j7dH51Nbj4PGcRVUwAQZnp8dYWhyp1BY7kCTJop
KxczA/VJJ7HNi7eSXTMdsRG5I4QQ9t5JL6WutjG6HOXdSndB0R0LRBR+LztfjCuS
yyZ9gT6QkeXZBWBQomdomAHM8zyTba8R1/oiuIYvdOP/nwPr//ugk13px4PkHS/c
UAXCfqQDmi3U44tmD2rhhO8XGpng1PiePo1u4R7S3KhECg8VhPsgIjKOL6h9zYUD
agzE/Mt4dRrJQr4Oh+lfEXoWsBTIZAHXnVpNXdQdg4PAcOXEuaRiCLocK2xrMv61
76GaJkYW2tM31R70pt7ttqyBSz0W+FoGV00EQ8GE+I3WPp5MKy7wHJ6TDg95p2Kn
C8G11xDHOP1mjFSlltGr4TcVsvhaoVIZmPhAMX+xRzV/HWRt1UgRYBfiHY9vSeVF
uxmrglDM/P5iD0SD3QAkvx4mPg6rej75mx9aBaOIsjEkn+WT+zSzAXglFWH1Ky3Z
aJ6RHpPOOOuPFOgrV9QCWz4t3UUlikBMXggbSSIUmB4nkm8HlfZt8wYusrXtGEzk
mi80ebl9SF3DAE4lTvw1fD2V2UGscxt0Dg0E2o+2nFdBVPWN6SK1ILMZ9jRnjurZ
p3HjKmbnX/XOgCANhr3PEFr/iLLB42KDcF0DD+SMeO/xF75/5eOFg+uN4/I6i6fJ
RBwJ2FvkW1K7hRLwvbSgS3CQrW2BB7DlwIgdoTKFk7E2BwKBqowqmEUxZ9/j7u44
XZshQWmkWgaO1Cg5pATecmUZWkMgnlZ6+IlASJQlfclEpaAPNTNQcWc50Xn8bTZk
N9QA5Xau8ysAjCXsPKbCrtXCwswgMpRR/YJY2p3hv3Fe9PRBhLDJQ4GYWe1zdxlm
Tp2gAqk0Bs1KPz2vz4Hub3/bMpTYJ0aX7hRD0MJgdKEJWCfHPzlvenxdqdk9RTll
4jtCEV1/rDxdpl10KXvezaHZWSZhtXru/ZDnPfqTNqYZAEqrTXKdxQ+PKzgX3c7m
m7MUiH6puD9axTr8yc+0szY5EtJ4e095xL9R/U7xlM1ThR9z4B1VXandKrn5SeVk
KukakdvnsvFkSBvbGl2sb2BXk+EUfJVUEdBFQBDR7pSpjltaiTIQd6dqkEfmsjEN
+SwEXHtpqX7xJvZwuIVj6HqPj8IEBocWuT/FIJOrEtN/Rag8bmhddLhiDtTij+yd
jzfXBpRaKGPSXQe96zWzMBn0sj3if74eMMIjBJ+vbuY4k8ijv9ErOkGDMH1Tqw/f
diHu4J0jhGqvCr6IrSzQt/NGmxrDworvGec5lTPPM4EiotbI7Jw1TVGI8l9XJHUb
YcFvfh/Noc0lTREVBqb3IbAGck6ext265G8n9qr2oBqqNcFyclusRB8QmtzkP1nh
3CS+7B7PNG1oXMV4VKjiLvmFpPL/VAwWr0tdevz5n77arxFD7tp72EMZfLbN0JaN
kIiveaHd62MbUki/mMdfLzyBbCWOfpF4+3NdmMnZHmzhgDFG4O/rNbgAZ/FkhkxT
I5KKEBgzP+ur9faWaCGOSbQJ4/ephbdwbziSijNc9HuBR7VVFufI+7vPpZYURu0J
H6QY9XyjjCgX4xUQ9gL7Vghf40EMvwnTPmP2EIPbVf2OXQkEPhCwsf6eWevb+nHB
R7gmuGIM9eu91MRqZCRhSvDj3nf8Ha8l8LkfWQAmOVoJqI3570dRLiSXIFWRelk/
Dw3uB3uvPNbS3aVz7mebMLxBNXlQn0uEWGbcVKX+fQpt/36OZEID9YkDW+j+Nr6c
TuUjDx8grJlxu9E+krXdDiP2iEkCI+y1FWbc85nS6HXlhIm8E2mMVcHZJrX7CoE6
K6jinD0POXgWfOCUieK4XXtEDlf4scUzuqf9z2JH8ADrHxEgbwp2gZn8D0CC4YLw
M/LF8Icx2YHLo4q/eY7LNsypWibcCpsZ8mYPlfYu3K8tlKa0Oy+jbeolj1x7be1J
G7h6jp3HpG8quq31zxkBg1lqOur8NWzvhJ0dNqlsQ3E82p/L/Lg7wWhRA0EFTWPo
5OgQyDKRRAuABfwyBdXoY9nAKdq/3DT2gVx82r2THiR1TXPa0zYCNGdvFE+CAboR
SrXc8+I/wt6iw5SexXaJ22DsdIfG/PmCsNoq15OQ5jWgYZrhMucxI2FxIQ1G7UVB
zXgIGe7s2SK+4Eqk+AHSEsunw0GTeWKGhECWgH5vxsLH6aWuJ4h7SJsk96zL1uZB
E5lACdfBFhlGOZ04Vm6dVcmZgwFEFgxRVwCrKaRp8dGcWxHuY5C1MB2ddiXqtvyO
mxeRh3U3RCS37d2+eoFHhb3WjNudZ6BRdYmrGTBWPP8Mybvx4l6ba7KfE53b1qf6
n31hY+wfztnHu8BBdbMJhz58ScLlI9IFXnO8ZAdoC5Dehr3QjpyPOwBPb8TBzl1P
AzxFnEJbZnRS81MZnmJs3YWDuoMjERXk7jffQQ+Qhl5hdDtxQqR0wfS4ljCOk9ti
kJYT5WC1Y2gZiotx4NWDLi4cY3KCOM2AmCdcmm045qeKAUnAdfFd8Gi+r2ES90FK
Jqc3WFDBjcoefRYai3J9Z8EYGXwsR+BXIcTIL0w4MupbIctHohXjiFQLIuT5w/jK
zr6BbeVsiotfot/EaLiIAT34ehfk4HjKPPKIuRZbL/HN6ce8+SIn+QDgOkXR9L1b
afllrbbhWmPjfj2eala215HVWRswjfVMqKD6yN8E7mWykpgLUq+Cpg0RKhbumpYh
tRpaZwVY0RNVtt5vW2yH1Kc8LABLloBBaY/+Lcu+esUsTB9KGkZFkS1ATbFH1jJv
JKkLO8StohxUlhc5CGl3oWASp+6tP8rK75X3BFFyDMD62wFFdXShraB99eMk8L/D
Phj/InACgKzXDaS5n2nYvEPJRw+lJVmg+iDlFKWoyTsAis7U/7A3T/NQyoHX2whk
mp4UDEvw+92aOmv47Fe3Z/WR5rrzwOAOudNvqycHhpuBk3j0TTh1JmcwVWzRfKTe
v+UHNR68ta69clISEBfId1ZM4bq4Yexv5J6hQbg1mfCcc23NNm22KqRi03sGcc3h
b4dywwhOdfKSaczJKMoKfRN/+64FUx2aAr8Ze5f5EIVqC67vjFz7YBaIUZQ7QJ7Z
ZztK5ayX4DMc8iPVtTOgPV91GPDq0rKqfbf9wcadsGQgflxGaPaVGFytFzB/ebZ5
LhCUuBmsMiuxgGOZ6UV9VrM+17u5PSTNlh2o5DcXAjPT4WDIuL2hA/8decWTAZcu
1xpmKAT+yBftJe8pqHHyWGRUYgWdyzRd+Nj4DW/nOW3IWs+XdizUKKo8InvMPUlr
6ncoKMDKeWSW5DN72k4LE9wxbgUCG4DLdB0+mMkTdDUCF62Cairoqqt1iF+qd/v2
KKeD7GWJt5rs4WuV2ZaFvA5lNz5f+v0XC/N7RIMYd/AsqqUQVhlKejt/Ehij6YY5
sfSFUqe88r9g52ANLY8qrxolR6zdcBkoKOl8A4K6I8V95xkg3j4kMp/jmrwvwhUV
Xu9jq7Zdtm28LbcKhE77sCtgDpwDbB7vS51qJNN40XYrRu9Zs/Nc74vC1+CS3OBM
oreJOac/cICV6/odrifIbHqr3mHEoWB21J3arIcwDIex7ihoHRA9VM1CLGR8morp
ZXk4rlFG7E8vsnSrN2p6wsNuD5Xkz4BEeBSaToW77SqiLc47mMjNcsB/08dMGg5b
XR0oOm+8F3wJF6ob4dTxZPf8vdMWR+9Vjo4TeBDctkrNXuBi/7Vcx3ah+iVcgUES
rRO+ZTr45lj0r72+Ixuj03Pc0NuuUnl+yZNwzGfYPtnZMhNCce2XzwX09+ecDVTb
dvNY56hSSMHvZicY6OvdiIukYSAakl5JWSSU+ILI6JuD8F2V+Fm5YVmrQUYEjerx
GlJM+Aj/lEyGhMVuhMPhr/Qob3QG+FYBV35gKPL8txsp6m0HX0QzCX+iItg11Dv8
k3gYF2lkYoEA+UlhTDIk4Fkl8o9Chm0lel3mFcmh0err9bmVTU6foEqG2lCQ8X4O
fPTM6otzUpeHvnyJWRjhs0rm9cuToL2o3uQc+X1+RYog+QjDSRwUS+M2/g21a1RP
V3eDBlD1Q9+HLNRchEeVQtKcm0OwUmRa6BM5sc694XbF249Ucd2nT0+NJy3tSb2D
Q5e2oZdAE4GZjCnjetbvbje9CL+YUD67MajgQxojZp1bziqleTI4ySD3Us+Jj4uq
UrIc7RVFrvrshTTlqgb5Gg6VYXv9ttkTAHA2mhtlUjlDkRxZ7TqTxRhVfX1SnrXr
SYeRPVQ/KrWpDU94CN0k9MepuguIqkeyRkrIilCLzuGZfjtCNjeoP7gZPHV9HgKn
InumF1Q5KyQo40d74d6OKCNzL4Xjh1zWe/3xtQYmMFduMMmmwPJlDkhSS1WHUiEm
k3MnoOwsUbFl+sswoLpF0njVQsNG6k37ireBNrpZqtfeJP7O9xqkVdvOkBI4QpqF
hQTaGQbHtouxi+ev9nlta569hRHyY3f7EObxMWdc/WQOEaZTOZASFWrZvX+yJUG4
F968mmg/kAR2C9M1RnVux0lPuSANqe0HRHKAHGZcwv6zziTu+dYOj4zxM15EjBuJ
MYioz2EdV71Z/ar9HlyKrXbRZHmLsWc+QaSCMdDweAE/tQTBbxIV1dfktJyZLbms
SE5iEPlCEM5vUp+NdaN6wUKjKhOemNpVWwMrc05IiUVv0QjbBAlBmfSl/rvYaGpm
HaYmHjxxHw19KrEzuTdsbDyc5pOJtMx6FYaR7e/KiuLvEz/uI9VQUg2Zjxg9g3w4
K7hgOiFtBoQTgQ12IxTgBJMjVr4zLcNyi5y0GWUj5zLQsMWJumPp2jpbiZh7qN17
2+ZkwAgLxUwv7g1/f524osZW5AH+tGLYVQebZgoiA7rclDFYGvYP9SdZnDuQ18RB
c8GHengFcaWsg84MxDLBblNtF8GkMic2gOb08kHNP9/aZ96P+whEbXc/q3s3Xt+i
J0f9fgctWMA3aT+aO0wI9xP5NQdkLQgvnYhE6v5QN1NjE3pluoyZmK1PEUNxNwR5
MysYNxry+iKPYi0UN78PRvAjGsoqYR0+4DpJAsoCEAh5zYaga1Iygh/BEDW/slA4
2O7+MO3/yffZZW6GDmRH9UsUpQ+xUoP0fOaC/oH+02ErO63r70canIjAvbBnMAu8
JzrLdFXtb8fLKuNHx3GmKighUKNAcmq/4u0mLaY3ey4XpI/xVGYO12ayyyHCc56a
73odC5gCq3T7Qqam+BttOerT3b4COP8cHvO/n2VeN2vnQrCnzW7b/Hw0PxWHJI10
HI+ugLxRXG+24GpHtJ/dERHKHpNocSuGqC1WvkU+W0bPgfLFnObiJBAl9Ope+Stb
yK60hBH2DuRi75sia6GKSLVdg7xKaSm9W7Xnwp3DieBX7RBEmq2zRyWWrOCX7DGY
UhjLHac6wl5AbgNi/BAgFlUnA9E2JjGFYZ/ho+dtSzqBb49hEhw4cjt5WQU6WEtj
8b/OKXBAjqUHU5gmiMiEvGzpSdaCZpe9udwv3U3X8HPqtKnJyi/ctEGbW9n6pMGF
SMpZnGcb3s4qUHBQ1LeuyaGVGjT2oLRp3ntEDlti1u+2IeX70tsjimbDaEF4G9lu
BE65EbP7xkpiDkyej16uRKSZIqv0/WKQQi2YOenBfkMjPJ20PWJoxKqblpHpcBxs
Mym+wRxaVCcO0onQcLJfKCEEUnoAY+Zm66i/eYtokTuwPFmcHqwjvjWQWo/NCu7D
rtPfC0mHGAtbBpAeEq33hc+UsAxad8W7mGW7i3BgRe2Xx9gEg2ZQU+BBHjyRiqY8
YZto6p4fCkeFrHSvjPZAVUp1gnWiJN8nK8K4edaQQicxN0YzNAfL69/UvgIIBAUQ
5Bz59KBPw5AA8ShKLrMhecuBqD1Im1rgMMYIFBE9aVmWh4USDFAkiRJOT8D1Vdr3
Na53Jm635Lmhx4fe3ZNPRHnsACbcM5g1bd20weCQeWE2hUbKw3Q3RDD5odl7heE/
kGEoFitHgnkLJhwNUpH+3W6ChyYDdxKsP7br5geMmxyIZSUkEF1QbV+pwPD77t0G
fISz1de1UCg5NBOJz06VZgrfiyWoi2g0BXXQIYkFUuISK/m79oBHpzzr/QfJLy5T
DQt459gWJonHmHEnDFO/5Vx2y7U8AtKkeaJmPPF1QBoflDHb5WMrneLlLvJTJlE6
hjjfKf3cickjrZVTP6qEoF8660ITHds5Mcabs26FqKuvkVBiLys9u6cRBC3XADgX
UoQk7/63uCHw+AM7Zvl1mzX9//2JqwMFJ26QDQpejOGhCfwJpYtdMGuU+2swg09a
2a77Cwl1HLeaXyJG42nMxMw7LYrGE5BDbwq4c5yNivJ6OnVf02GCqyx0tdFFAyL2
PCiRYPlNY5QS5oEf6iFAwYxHuyrElBuGTTIF6eZk+VFgx6aTGqpoClaBMsP/VV2L
jHc31SZsp3fBy4P9CQISych97G0RPEN2a7oNVE4RdsoF0D/rQeORRbcjhEmd8Ik9
Pq59WUEO7V1thEU5zhKbb81ldo4TWFkY+u8dBABX0fJZ/s9BYq9FcYgfOASwajBb
fNTTpMgdUya2T0BJJZxJXWHFwZWulic1pg88nee0w3Au+WyKfKKK4aG6QrP8Rj3A
4KFNOC9roWQDhxZuFWhn1na13YgSiufYa9pLBC997NO2K57KkHohWEbTCVk5kLkW
reecuCQAcTje82yZ7MMDIxH8j+27t0OLfIXlk9Rq36MHva20lw5eEw6dLwbqAphL
bKmb31r8MjYG/tqRhZw7oJRHFS7VXIHa/HJY2tRSUabcEBS7yKM58dJU4N2LrAdP
tlwWa9dh+xd832eLUYiiLcFOe4xa/hRxYt3ycksb8IaR6Y7yVQvitPbuHIedXpUF
IriF+bHSVVr87uyBL3DugzJ0j3C1P+b5HAqUSuPrab/IsON6OAtmRgkyYbOUPq0/
y4YAUwYo58KBSFo6jK76QB14yTHJjDELPDYSXbxs1kjeWlRo4AebAXh7aU9mJ5d6
h62cBuS6Bp+gx67Bk/zwuf8KDEXNQ2cRSy+GDavusXxHka4qxMwT3El8fd3ETbIQ
gwv+EQYSZN688dq3xkxLRF+sDpNdC85WB+dVXL+BSBQC9472uPJUyxNFJLaNf0Zh
kSp47Orbi3cZoNen4u52mKJJscm0TP28CHfv5GYJwIYfFSFs9S1kgYF3c5MFqLcT
S60rc07jUGEbtAz7+jQn9E2AEnOi2xLuX11d6XPLi1wdIbHS6szwb0gsGs14jwNx
aOBVlmYkI3CO4rl1of5FxQI9Iok2dCvF+oyecCANlOGnM2yqPMXWmUOevhVivEUr
SMbx+IZVtFMRAxGajfEXAdVXmV7xnB4jmFSH6NIhW900/5SJpl2yAehK7cQ01GVk
kyyQ1H4Tc/U4Sj9dOV52EDqQuNnLVNl0Wowa6Cyr6SXjY6cCyC7OsePIA8GKEgqn
SbxXxaD0iagUhF7YAfDdhOlkCia6z9HMTosZ0ayRX7dT6PzK4XhdPRqkqxfqRvWa
K7BhvjUYMaLNZ/mwRNxpnSWSfsQs6SEryyG5Sc1iDitS5H8PdhhATopCTVcu76jd
Kg6o6Jl0VGW3PAQpojIhsXRvosnMVvRWqlsCkXp62hKeY93bH+YFg1uE89UWoQSJ
hjb3il8fxXRkr7rYoa7z5jXho1URNVcIVttUY/HLIYIbXGUVM/9rc8oiTAYxtOQ+
cNk9Mq10Ys7kJzOZBwQqmg5rSfyeZKB8e5tBXw/mlpbmVZaOQakf7Nbogwzh9LR2
X+43m19uD/4BmC1GgKveMWqg+KqJmcPpUn1b9uxLvxRg6MlkRD7XyBxmLDBUfyj9
kEkG9itz8OdaH9n1Ruy2WG6IaulM+lsLTm3bIsQ5QVSBUE+qD28IXZu50736glUe
wYpYmUFvajnHuwziV7BJVXMQelKHPqA8GJtldCTc/zvJpQD+FN5hMjh/f+EUCRtO
L1PekbrxVIsMOgzz1hnXy55tInNbIpjtD3vGjl8TkJIBQ0VOpmA+9eoKjQAwUyqQ
lhFjaTDuxgGKYoDCMLtsgmVAY0a7q/KRIsSRTJM8yIBw5+qE4d4uO1X247NBb2HP
25W5i7I7O4k35UUmeSTpUpkDNhmmNsAgDFBjQodHItLkUWP/aLDig0ChFXjwMb7y
mGD9peITAOrdE1QCOhLh3QX3basf+4hpoW759++RrM0JNBpdhvAD1tUwaIvX6CMl
zofBamv/wdMX7aONONyYMHGzOgjBkLmUrM/qH9AqQfGL6EJLNC6byZHJkRkP/Dz5
TsvgCcoPTmGivXoN8cTd45Wx89bwyWh5MkNGCTPHN4yLBrpZ7KUOKFrlERdfJ4dU
tlTu2PAK7u3uiRs6xvYQ0c58DdAoU1nyqGIvLDgFzEMmg8VpcwechYs197fGkEYA
uo76Mp2TLgHlNDnO2UPV1dHjkuxx3Hr0KZ90SRFoFvHSrLVqio5Md33Zo0Ew+oa6
p2YHQ0FBMdGayYAX6an8pp1NklhNoz9RBqGmEYVP3ylgMr1DKj1IOfcglzoVJbgg
PZ0VtQkUzkvIVsCXnR4ckpPZlSXQdGuWZmmlMbOwpjko0aMec0d1hPlVvipYopev
oxQllkKWtgZASdQbnjFUy52Boo7NPcrptRCNgL1GIVO8DQ+9HM/P34CmkRbz3F3b
VUZHtuLEcSXnr/dm/ln/5GiDmP2pdiHCmdgCxfXaYdsSoNXLf2jcPJtegokCuQJW
cjppWTGBhNFL4HYmtCe8J+rz5OSsE/VCvaFcUvfTKLGHDhZw8JZ683TODrn47MuX
McHDY2sTM2RUYN8zYJekxSMS2bSMb8n3yxq1qEjaHAlOKyyF3cX68wfwI3GGpUW2
v2A0kI8cg9J1bTzustoZGiKy+NxaaonIIlZWV/V63PEQyWOzg48sgrOdxwiUICYN
G4APnW/Gbsa80hdWqiVpvt2FxX9tqyuCHgjIHlGKlfGkSXdxpRauiFGUdmmJtQie
2DfCa5L7+t67M9vSQZN0ywAyIsxA2OqXY3o1b5TFqFEsib7pvX624S2lcv1aHMzC
ytl/4Fl+UWGANxdxa0af6yy8zWk+uH22gl4ZM6JabjX6CuFmv3GQbRiVxd8ccKis
yIx0oUmlM6v9xYqSJZsfaJvVlgiJlrEnvDv+cv5XTrBBfJaTFiLRasM5PvmURolg
1wZ3teO8YRlwOt0gz6c3L4CgDCwkv5IJxDWYJXenXLU45yiEr/jEwUpntxximICl
ii7T+t9Y0XwE6FjyRIntwEOe/6x7ebVWLlnHhIGSJmurekJP6F67L7Z39ptShHJs
4QTvLfPFlbBiPE3OuxSiGd9P65dhvNOqTSo8ohgn6elCO+ow13vKO27Z28m2E+bf
wgSbOx8nFssVfWhSEVXgOI2z+0FvoT2/n5ow1uNHK+ZezPHZd4grL9r4SATOaIeK
sy1GDKZeTto3wJpSJ7ZCloNCrga5QVlDGZnE3GJCK5TlL79w3MVnFJcHXGkFKrMm
iAJMsR0nPF4ct/3I7FszjE5VYDMXEZT+vpPbTlri4axJAAmooSzcBujdMSHOFaRk
cbzM+fUrNqiAQcb2vesk4vztPAPE8DIN+W8tiPo5dtJ8yhLEQngy7Z2AuC61GezE
XxUzaX2Rvgtzbnn4dBrk5NiYeKhTRpkDG9xtiXS2cCVhyL6eersIA9evNryIe8ZJ
yisfI72n/knLC7Z+vKEcELaGz8GbF70+m3DZvimdCznTD55bfoZEY8F+EyhARhnu
EquOYm4wmhH02k0ruzwFibi1cS0bVHtvmtjQTsvYW4S68jyFRIZHWm3IfW5UqMo7
ZmTMo74Mw8pe9SXg/XyTq1tbqJEdKOZDq0ES9JtZZ8/0dLVo6vJGq03kfyvVQcHZ
Q1ixon6LQH5wRLpYTdjLtyp1G/KIhLDtWvt/kVCArn5yULEX6yyMxM6RyNeUjbBB
swb40IDWP5GsiIz0XvTUugNJ88awIMe77S+5wE3CP1iVXF2QKAvZ3S9u78lqrd2H
ylhaKfQKO+48lBYF9b4gvHyg8BYiqpABuq07T+HPqE89c2HJu5/0B3LAqpeeEXkR
tg7zaTib2rlRlxVr2Ilxru8opmBAGRBmw+4zUjoRdFkkzOgC6vF5TQwLG+oudD1q
r/ki0H2SAN0dpaXh8/bALXHIFCeuBjZVy4Ef+YdHJxiy73UPNfWjKdaqlONFBuqk
gxBl/31M6ZgaoQmW4KrWR9xRJi79pGacmNcMx6HeHPIHkbYQoivnsSC3L6c9O+8v
R5y9sxzumk0EQXzUgFL9nhAfBQ0giHi5vtJllQ3AZS8HpKIemzkM3UOVnQrdB8Tk
IgbQWlkX/Y83Y0+p4+BG/3SjjfzZmCHB3vZTTYVWR7xsjrw7wmye6OuamDU9Ui/S
rAIqVoEPtQzD0MPp5UwkSAlmjpzaI6OeaL/8DldWQoUxeGuJBCV4ei1ORMlVxPu7
oEwmtvb/MSshpLG2wngOe7YuqYfTmNn/E6eQD3O/8hYojAB7fVgpqCGoI8VgW1iL
HqmHdTivP8dF+I1qZB1Hk7A2+g52ROTVjj5lROUOIbiNqesZ+LZiqKtNYrWe8r3g
oBwGaGC6sjQRo3BXI9JEgHaa/xBF9gBL5q0KL2pd5uSlQWaWTPzPn6FnWfKIZPka
kSbIu7a0VudIqma4aivL02u3GR8Z4wPO6RBN7M7Lp8aL47Tw3lTXWFdY8rkHeXU5
5DvXDqfK34bb6xNz4EdbJajBrUhVyYbTRTwkgItiv3UkYQX9PizCOfOlW8Z7wC+8
QwS2wbToLecEONVeUj6ktKWexJAFtKCOXM+tWPHb4RLuQrZXn/PaciKkN5fmZEZe
h0EEPX5HvPJXZB21ZnrgP++EPCasrapfL4fN+2Es71ki54qukvXmFJHY5KW62L7p
fvnE8AVDBNsJEi5W1zZpVxLNeOEBpS4nlf8SyL5+6dsNGlg5MXfsSvRaMHcGljdn
A/sE4H4fAtuH113Q8upua10r4odWd6pBoiwbRCD3YR1yXyz1kP+rF48PREzwE6JI
IhZEgESaAZzPBSzC5U+sHbSyUbGpIC3tH0JKs9V/s++VDFNjXTSp0y2jhkWq9fRd
qfvn11nAzFs7Y8mgTCpR3WBSiuftXSDELIubCDa3qFIwcuWkNWM03bdhSXwKPTBR
SVtghKppAi4WmtO3y4GJzt4QrZ3dTbhdLXvSSbpSrP9DBEGPPFzaOLHvtUVAfyp7
B9jt0ESw6pkNzwEasrkSaIcF9ytPC2hnBE0Q0f3KlXu3ZWsXafYIKD3TTm9xsiOV
FjT5Psghi3ChQov9G9Cxf2YRznhNqeuo0wLHPo8Db+dPUkq+gV5odZCXHNLz4qYZ
EaI0qwIzaYw0c0/j/WyFNoGMVHVz4ZNhWNyskwEG7Lya5XkhgMUUCBjwH4u9EeG8
qBoaXKGD43MMq+Mk9OMwyKpckndZHuhyPXgodywGLv+tXyiuMOSSdUpbGMtfih9R
/JUK2g8kUTrg7kOudqzywlPyyrIcmbN9TTTTl/dIFSp6LE+vQQDQIjZjkYBCxWlF
E/c6jHHt9COz0fAG+pruyDaTZxd4FS/HDzwAdjVKVMz917F8enOndqbUNZVuGaU3
tVNjaP1cq+X+eIZPig3mtYmBr1Qds9BIW06A6PfTrbpxBIt8qv3Wr6LFx8o3XbPs
gQvb/9jvCxG7uTxSq08vj+MS1qmxmKKIvI6GJTxKgQC3VAnu/A3ImWhk/R2QBJae
XC9PFpL1j7c+oNY2ULfegYborKYwIWpi+umGW0afRJVAjuniJrMBdOosJoGbtTHo
9Xj78CV+xoZObWhRggM4qZd9UXf6MTnYWaNK29x89R0bgJ2LjCZIA0LUb7XcbNT2
9FydHH1nHoS6lgzSLrZmQaVJnSvANYcUyKR6/CYtKqZ3SViaXws/XsJTlHrFh5dC
1HbxWF64CsXBx28us/NivH3Uiv9kUsbj1x2bQK43R+vmzk5P0Ddz2mczj3HkIJyw
Ddi+/G4ClzN5/S+PArtKXfZI9ERY9HxY7VfOJHCmBg+hm+NN176w6BRTZvm3p+PX
qb9iNlYkMo5yMSTocLr68vHL2leem12FVU634uMdJDJhXmCVmpdN6J0mxgJdwORZ
LK9Mdrc/KhZFeLaKZx8tRQWv+MelejUF9x2MOC8IMwppLv7b0wt9Q4niPaSoppWa
nu58FhrM6Jsn/3pX1eNTwPOeXrXMA82sRJie/Veqln9Gq7VDhBJMviQY+CLxoLIt
A6O/ti31UiNhlV1aEjyL5sZv6nmLiz1Rbj1T61entTKLQT8JoGyQyDhigkGKcO4O
7V9raCk4T7Is5+ewv/Y52n56ihjYkoKTtXuUZtIECW4nxWDTasU0aPo6+LNjgwBs
SdlsAFgo8vlOiKE0DqKSuD0HKHie8tsFQA/PZwt/Y55bU8YaJttOZ7l9j702k5Bt
B/XVliFA/HKAa+C4vTS+pOib+etN/YVVpk/cjhdkmOPprSzDq+op15zZ01CHeEfy
3KPds7JXBWC++yJ6CikHYOG2mXIfMbI5sbTOl2LvZX9Sv3olUBAOh51xQ0E5YUoT
ATMpUvbWyFOXLXVU4SNigfYCXfvfrnp9EYbGcafuQLMW8C3jtOC3t7edsGa9e0ws
r9leEVL9uyTtJ0ibA5y5u7BKclyx8PXvDo4+KSM12VDO7Uo9s5zl4hNuEdyR1l/e
ukggA9zbwAPZ/coNltB2UfYstb8/F5Ptf1aNnfk81KKJ7kPptB+lczPleClHG252
FnPNMan2efnwXMTHiUjtkkznKwxAg4uscUDg2wXFLy9vWvYVHBYve7ALxR2LcLVO
lSAVVCpAo+aZMK7ZUgBpJDx7d3psZw9CWqSCEWrcP9np9vBPYuS4/crG9l7urXAt
AB1XN7CNlgtubAZesPb1UAKbYOSwtpiYdc1lZRGj6KSqxGKEuaml3e11mT22Oex4
38hRlXTXCVTVTZgH9QyXyuAItCq4ozr5fZyV1cUulCWgoro/Xgl8wp0bPQtOZF/3
WcCB0vpwbBaWTZ8e0IRJ0cQvB3g5wDn3SEndS3jkZF00SboUn1ZBQjCPPNUVi6TV
9y4dc4p9VE0hKmpopnmfJxYwqK33Nj0y1vkKgkCMS3lCXK0NvKy+cQV4Zt+KFHds
x+MsxOs4aBv4IQUISSmCWSPnuk1dFfjeXW1IeBZlH6Tz9f2jbSaq+8PizKlUb/Ni
3nNiVgAUTqVaLN2R4vry5Y2yvUmUORBI/eltIgCPvZq43R/jG9slh2qDyUQ6j9Tw
00+gQGSG+3a6jDwzvW5RSzIrcNKVkEoDRpQWh8wVBNUX7lwh8nKfaXoXq3npoTAG
Jzcw8HsD1IQB2vwI0KywgRsVQdVsrqQqiBAETj/YR4Klmi1BWVlQC3Sk6RfP3BrJ
qlppchzmJV6HdE/wf+K+fV5IP7RqFrdvAeJUMjLZMqXJfhO4h+ow+jUSRBQ7MC2R
zfd3E+vVqVddYXKfHzC22GXRvMi+RAmt2tRvgdig4dapWV3TLCPeGcgq1ApfoSWw
SSJIM/0omRBpZBUcVfqS8CQfLeVKbN4mTkx5f6q+roPCv5pqWwY6Gp1auZ7yVau2
YbgVcOvlyKFzAGFQ9+2sSvOBxDFpxl5cx2lveiwng6NiUOdOkTvMfWbNnwv3f86F
NinSgESoQtWCgJfiWJhtcbgwnl4nUkQ85ExhxoebIpoDtBDNDOcszM0zAOc9tooX
OpgN4rjjBybEcnL8qTXTlpWl5An2xDjcGMtTETURDvcpZb77UfUDPCUcHSwoDwIU
GLkAnNRbQC3tWGTatz8J+VuV1+dUSthYFtRBZzXpYETvVIsnqf1LXy+UfuTPtb4P
nJrmVzVAiSHqIzmotwXmq14JMm4HNudLgnWIacZZc0nTKqstmrwoL2bcLSCShjic
ZJfPTGPduDl/wpSXme/BVuj7YpQ4IKKb73P4kruxwUYsrigTahobsuYLc8ZIzxBA
WZvbY8XUklXJ2bQBO8P6nxnpHAey8/T0xiB8dNpNgru284zWy+yspGbubewv7mR6
E7ixIrDx7KV2wVzz9UlTFphTQ7461FyaePq9MJ9hxuvb0eJ+Qa+aKZAoqlW4v1Qn
SnRF6/Y7Dhu/AOUC8z1R6jiCyHPMeNAyqIUbg77r5iJFiIUJA7x0jsE7Mjay53zh
KpJfxkW3nbUvZywCVYen6ippV1UhKg7n+Qwc6+NK+zTmv66wprAXsxiutod6LENI
3x7/8XGumOI6uGdOTa363ClVWp9T4EocZTdQQHoGkrq2vIg9rouli5N6Dv0ckfXV
Y1cPzir1cpF86PgoX5IPkc6rZ2zDFM62fIAQWWQjjdLqYJv7AioJl1sZctbfNwl3
ofNNKh5DLfwhpsLvsLYD0QwV96sysC4RqlQGeIjWDlGoETt9BQy70vffM8XkEgz+
ygCjCfImd0GuUKc8gSZvurmo6jUG0EdiA1gl8y+NWAkEjoRh5WswkB5nrZq7fylv
EmzWz7pwn7hyDx/dUW14WWC8WXTRzm/bvrK/DX1xvFI59YjswbveGGMLekH6/58Y
M99PRxBJPfEjGdOcgClZmtE6+IcfnK61Q6coDRx4STQEN+DX679l1AYavsjMCdJR
9sqKz3b9pAa4iB8qmBVFQaRKeRDjKdN2EmqqN4egH/o2DkuxElklGr16+GdRUYX5
NU9lCVFQU7+6Evn0L90olvnaBzIz75/y7NdIey7DKGVJ4o9cO86gE2PAYJ4RyYzq
lTA5dEZ8/rZHeqZBY2b3hV2peHO1s9ekgpxa2BKtUz4n8sLzYDpQgERwkmjY+g8L
lOcYgTZwegzWj3+xRG156V3K7CmoCO2CpMNqw0leaMHehw6ySZ6zy/288dyhdG9I
8WMzpUZxLUCi8GJkxxsGckO9Ixe6cHKhza2l2BL+yJHS8ql30tP5cOfuLTTydCRF
+4S2ACd2AXYcd0FqgWH6ypX93M8bGgaEV0Bk3YdMzlJbOXabHVQcMeAOpMZX/EZ8
rbUKeVHNn/P9tA+fC4Q/pYENJYBeefU+oXd+g8HNjCWDplAyYZsJ3wnVKBOAEPBS
AbMzeLi2+gTGb81WuBGNTC/wJ9808oXdc/CTTATTEjSnSKXcEBvjQZfm03v9Inep
4dOBz6pvEdml56Vxgb1pfMlM4QrwpFiGUm8TBolmB6g0mvfTwuLGBs2rq8oCKRjK
Mqzyj5M1wHlze0Qy663AbUZri/f5jD45rJwd8I6abFByo0mR45VnAwEcbz2kGumV
HazzBs3o8qrQbmK2h5YASR80Sur49XQImG3Vs44otA7BmMp9ZySko7yU0pgbl+XJ
wrWnyanmtMQzzjTubLHPCEYC2LVhMWdfm7TdKYFJw9XSsiAWBZOXA0suznt39NHl
xMEXKUQr+FRpL8Wr1gtzEzBNb1ITimlS8Z6kSDPVkQHFJ6IoXgj+/n00tXI2Ko8O
LW/VMZrj+GipmrbEXXTLnIkzZTwsxJy8any8jqf7ceUhp7F/IUP2AOz+0OdESYyq
l+nzB/xJf2Z8NB3FPKC1Y90yyz1ng3hd3wZrVhZHNESCepnYCwWE9Ofmg0LCeOFD
i5uF+Ox/XbLiM55p6exjQnGrIRsuIXZfrhovA7+YIo2QaTM4VPjAnFjxPcbcZl6V
X3gmduLFNGFeIE0lQpx1IoJNzTRMf6MtCixDRZhsIN6iG5/9ykSKs/UGlXA9mVqf
2s93jvgX/2SS/rwnND+IuE1YDZ6wwvL5G8f+e1QjuAAkolzz91mjmhdk8ObjldZy
3GYbavo/OkemeZhPMWy3PqkMVzIi0SdxkHPH5TgZkrybDaHks5ArynOJ2X0HUQGP
stBcS81/nBsowVZCpsnckzxzgHvab8SepQvxR3BWXQFqcJDNvU4mJkQ429LvDg1L
N112Yqoezu7IlOigB3Vtj3uZXSw2V+CsHypl2M6gV81HjGjznPA2hFyRg9O4j2Jp
cCtCGbFcORUnLiM4dsgYwEzbYa3yx8+kglLn6KFCx1aLfsC9GIRJFolbHJWKDz14
EOpA2EkC0xCOgr25EPL50kE8Sqys+3dozXLCrQEfGLTs5khWXfEizQDPIX9Tt5zK
ypgDAxjum7jSvHMAFO9Ii4g5OnDTXYyNUsPDZqi0vyNFplbj4bKBmAaRBGyQIXfK
24lHxFLaFnL5DfhvuvYMi/3o+DBT3JoqZyXa6lkfaSWN3d32Mjd4Och4F9Bi2eoM
DjCCh506mpL3fZu2cie1rDvjUQc+dGJpWMK6gT2ZUMqe3T3odCA8u02Ax4Sv4Rkk
+wp/nS1EOXOEanx2uKXigHnwD5D3VEOS/NIIoyZ8mvPL9/ShofrW5rQgqFi79lpc
UDgJm1CqOoDrgLNr5lVq8IcU8ShBEyeByQXyujary12VX/G8sk8C/L+eJvrEuP6j
f6MnAlkL03Fsykfd4uz/L38UGnvassoEJucCfgh2VTfnHQshjjHgfoa+fKHZB5Xc
UduLIJHK8LrAzDBhkEaol5yBKhH212xj2sYWSeYIs6gd3hnETFv8c09FNWu8YE/D
KecPgPNgIEcIIfNKAPWjP5RHPU192jpCoXZn2YH6qeY1DYMTLSjbo7/bYWmYebz+
d74eQuhLrVurvaUKwnt1rW/blJLV1JGptAdAAQlEqxJcp7rFDhC8aa0Df6+qSo0i
P+AqmkmCNoxQWh6cghcukW/cyr6XS46/A24Hddr3uY2+qlBqTWRLvzrL51A9F1BA
TiRimBGwKveB9KkFvcIu4c6E9wi6oyJVfYfPWh3HJnF5Yz/bSqom6wVwQow3xa59
YNTeEeomDsh6jscD7gr9atXnE7lFss9yU484yqxxANKHqK3o+crQUiyW5MGPdcFv
iSJlEO6TSO/nL0kI7LfwP547U1Lzyx0paOHI90gNR7jRJdHsi7NBeKziq9I8TVid
+V5X622FSs8gTCKqxgEjsbJHbuN5/XU7dD+qwxqgDI4LZ3BLk24oLGs7p08gkqxL
x29WbwFQzDMrrZ8cmXukbWffiyDzF88Z0KDgn4l3INW9Koe9UG4Dfm7L0yY52tWn
fa4H5RwBRMoGsCwQ5YfQqdtcqwTVUkQvKZWP3VsSngqcfj2CTBQk8o0BIL2OUj7B
NBWkbEwmJ6eSAJzPfsBGvgUN5+WxyxZ7tDbidTtA1vRiQyT6Dg/t38618taWnN90
j+1c306I0/N4P1gqWhdJv3EgxLnPIFfpDIAyD5hLtt6TybrjHwhIZgXILPSHrM2O
YXWgIhgYmnw53MCVnwPgYnnwPyeHW3AiraPyqKqp3hlPKgxQO4mw6krkD85zo5mp
C4Bn3J1oA7keijPNJos/9dFCywo7oC2vZIbNfI4J808wbyQ+4jhOoYqhU2dGMzch
7pCrhtKxZL1bKw+w8UQYqer0tl5UFTU6x9NnDMsJk9y116iQh4/BGIKDMx7LGcKL
DxkvYLd/8L/6sDhiaOl3BU79iqtfb+qJmkbbVndCWaV2leIYcwPIESDqHNaefX1r
3FkKDh3hl7vSlfP1lwe2DdhdULFrDOtuXcp21/wJ4mUQ7Y4AYYsNcSNyvpCUKlnA
U32mL+PscK0bMa0BP5V5nWOgfSm3yN1Vq+wF6HjJq7OBJrJkSo8Z92gw8VPAim+A
KArPADCt3vwydhkTNpUuFdxzW0jPIRfO4yP0Yq/UnsLelqwyf5T40t9yXGZbSFnn
o1ipqAaJESJW5SegbdnPRlK155ck0dV9irT1d0hA9adMyC42QBahmMQ6x3OcOFGz
M+NqFC7LeL/X2VdzL86wh58kuGbKIPpC5HrKYuamWNbkw9VdtMZSmv9IO7XEofMk
MkB53khLK/DC1ka+d4o4ht7CtIumqHC1seuBMyLGuOO1RURbYaIHDK1GvODDWa6Y
5mT4Fb2hImYy9/NG3lIE7KwaLV8XJNyJH5EjDYpevKvtxnuaCsc3tWNwYJ+zOyqN
o1UNSN7/4GYnW8TqZ/LTpPmH1wFfuc7QYcnUk+3PAkpPe9xNZG8agtmwNJ/7brRS
mipGOH80syqG23rAc+Qs5XnihHKr/nM3GMHStbyrNETeCbhXw8WYQ3hy6/kJ/qyi
BIKvObphrRW+G6qp1GJCwFJ4vq1fP3wCrlVfrJohx6Hgj5Xk1a42lTsyrrEk9wIT
90dGcxkqbR5vKqs95rgsfVFNekKZd2sVywz23ItWnDofWp8/4Ho91mu0/N7YpNFK
9D7thqeHASjKsuqqlNBRyCpFQgNrGd13uA9794iNHczm1h0S8/zlJzzmj2Efaqhw
WQvLw48q3Z5JVN9QquN2IAraXRgD7SiWlinyGQN5hHKNzgfAPEpHEFXHmlxbhcoU
K6CYayfDCexvvIqX6iB5488k2zys23MxMwrolr8W0yVAT9VnlhbN7d6EN/Zs6rRV
S0V9I93JTLz74IlsXGG0YjMYAi6qj7k/FCSfBhFcGNETQV8cPSZYssOeMelO5qTt
R8XC3GqAhX0j9DcXZ50txuxrsgaL6mEmgeHdh1GtGZVC9kkylgOCK5XvJgPESBWt
dSJmbps80W+EutcIQPnYQsLMHfg/in0ghdEddrOfCSffrDnZ3AppdtIPffdvWyEf
OjFKZo1VNKhOoGAbWIAN5QbCv9SF+9HWimGQYUehu25SHg0Wa7n13wi753hXd5Cb
B48ZzF1ERtAd4ckOG7myE6k+GRIrDUaTD3AGLjpmovCbfWzj3T+ZJD4gQosvaboz
pnh0NQqMvtvFEpGlcW+P0rojt0DdOMmTPztFBQAl72SQmGJcssFAiLgxSwMHWuKA
08cY+s4tsRhkUt6/GOCoKu+qc1MpTDe9OcAtnoUmA1FfN9KuWENG12RUqel4SqWr
mtaeEUiVbxNizn+pu2f5D0olGqoXOtIPJhPbxTXKTqfUI1XBsGqQz9zUYsRhJ4tm
HR6C4ngwX9p36DqZWk0ULycG1qUE8Ri38QAGXHSp/0oo8cM9tlj3JGRIZFIuyYQU
ckl7uOJeO6RKjfIxCgaReZmgsZYD2qXiF5VtQeyxRvzqkpDyUXlOdMQmJPdA4sbd
TadASIwJz29aXrtgxb1jP7DZhP7ef/1DMVZmEr8T/NuteK1LEriJZT2C+XdaJUuo
YvGcyme7kmONjTiPsZ0S7x+K+9DgOEqxuOt8VrhccRNqyThdN7rNt3zfxnl4Pkth
JJwegkLPPP7cmREx8JPqExqwwmUfh/ygLnAV+uAyMA+Oj+gSRU4GHxix00hR6z4F
dK7gq6Z1oSwgnvN1kSJQioIIw45YsBHsRcit2aS25D9n26fqX/KHmd8LIcV/2ZRN
AkIRT1pvAcBXSofV6y049hIspHiCGWtdcd4OfSucJ4OnseSlFQ4XyHMqRSdAALj/
7DgkMERbCa6O1S6X5+vbWLUYi3Jmd9Zwrx4KHkOxClEZrfJEY/Aug2/6puWPP3uQ
brkNL0iVhaZCWUgpepH2xa1tYYPAy9HgT6039E7cZXMEGdQslJewQFpiOmMtxXaM
mWBhxIyhdG2Py3oWSKPcQUv/6roJvtbZChAPmLYRg8nZCithlq3LTaPQ5tHr1YM1
tcKqcLxMOKWUL+tkp5W0nLmnDrToJWwiX+A0+iMefzKdOUfk1Jzec83h5nc4mBFG
v3tZel4a5o2jEmqzgLKoHg1joexZxOjw72+uJTdyyI+GcVuFUKmnhOFWoDQIQL/b
3xa5H5Mn+hGerS0zwXyJ4Ej7Y7zfcCduQO4vanQO9lg/9/IoPmq46xEi0E2rlqsQ
nzzvNZkX9GiWoTzoP1Ug8GEtXpN8wlxweymMF5jWW/FyuWvUxTUuW/BTUqUuayGp
sgmxn66vSjGcJfGSvQhxaIy8VlbPSsIAHbdACvVeubrfYnYWNN83zYNFpyX9GuHV
dst4KH7faXlmVly+UsiegsDYYPgbmL8FrJm1CiX3L/TrLp9qcJLvUTxKRh9ShJP6
xFLbDHdXa6CUJ7SsWlMU80rWg8k0oEYdPfGLFRm3kM9RDfHq/v8XTAcgC5C+G/8n
+HZloyVtzaipzeRYZe9dS7f8voeo52qZQEQcCZPqB1X2En6aOdczl1frtkAwn7pM
JcXTm4zYYXkxOhS2dOOLnl4+3nRZX9ukD3veusauuZsn4p763gIc5lz2u4ev1tuA
53tor0q5l68bnM95TZgvMP74kNrTbvPKf+bf9fnTCbhoBgrWHxwpFflYoI2WtE2q
fl0X9syVrJWnyclp85vjt4Y8eYSdjfhaNKLhh64k35wBPhzZgj2hZ2sRDjyhlMWd
WZXAOEwoXSGSDGtCPXiXSaFQ5WSpV7Bqw4qO4Qwxk5RlHap8/cSXaNnFnNWDIi7h
9u27mncF7Jtte7aMJD6Pf2Cl7obAC0LN84Ub3ayuU89lVNieRplbSalyXSHa0brQ
Beg2qeOzlhpTGFO/3S+qNMjGO4HEj2JiDSL1twBlB46tPIKMzIBCRANH4g1Se8+j
wPT6SyF8BBcX7eL3IdlbTVvM7aLt5MpcBjhKEnn2fzQBeq41/IH/lOtBP04A/pIq
G1qK8XZhdDGZUt+CWZ4xiOv3fg4+ThK04Q6pVNDcsvBpc59PtOSxOq81bZlJ2A6p
HXK5W/pyOopYdbDmaFz+UCNsNIZig5lhC4i+Q8YkD/aIRdBtLi8cBkZFE6/0tht7
9vCYsYpO8WuGCDgNoopX9PkZGkF0+7QC/w8r2LKdV0/TdOogHnyp0WP3nUoxnnQh
mbzV/jgoz5+0kAefne5MbGxJl9iUQ5LUELmBNuziyq/E+oiVZDIsZVH/4kt2Y3Cc
vWBQsOdzoCylZ1TjuQUOaHE5UEmeAQu1JmkWlTe0UMHB6O8WUeY5B6y6SCzjNeV7
Xl4Nhm9McE060PRwg5rxYvOr4/VadMvJ8dB8VYc9XONDd1zw1mdipFVLslYcQilZ
M/7P4nHGD9aSwESttmz2hkLXvwB1ja5I6jhCBeGKHCG3EhUp83/bR2acVueIS5Ez
ySIOr9GFILL96vrHfUEa8z6o0p/zKYIPNFQtUusjt9GsukW4Pg58IlBAgO2kVeYv
+fZKWOfwEAxRh3WbaPgFcqeRZn6w2ij5iRyWQIb7RnLQNaPQqKxTtvqWdhsAvKU2
pjODkHwZjC0tcoPS9RgqhOwG6ketdpaAOw6plWG0PJ8Sw/gTJOAhIesinVmm50ux
d8B+RtTD1B/3ElxXTs82dD6WoWVI3H94LrTqG+6PxgspV+Hw1T0zciRLdO2vkYNY
fTOVA6LMUyf6Cn8th1GbHV4s7C2HVk1YayfXjr6EuqWRKqbgaqTIWj4BPygLs5UY
uBqm0OWuTTR3VbY733Kx6PH21Lq0i5YeaVkFHmb0iWBy5eRswXSPS7bHvlpiwivm
1GBzL9xoYxR9FEgdaeaJzkaT0FXML/wFGP6QleTPG68hg1GyQJ0uh7aCVdz7Ry0X
QIGstjeVY1SoadPtwnJp9rTa3sTGZIe9/TadDNNwj1dqcbfZ3+m+xGDSpOXETwUI
7u6/gqDOxyMoAfWBrFNaVJLitz9+PVzAplM1UcQujiCl6gDbbZotxYCJgDddfytO
+W02zlVdeSacYuPP2PMIeSinqcx0jD3KUujGwN3TrD87cv+aUPSLIct5jh0jbN2+
x7luV339ZyxLd5YjB/7iVLTGErE2daP0ieN+fc63NAGaxuuSwX63s4AtFtT5aC2L
An3Ri/dSOXyky0wWVOrQfdVb5qYhyHblGjrUbleo7p1g8vR6JCV4UQO+1uRab0Qd
h2hXNq4I2uJsGZs5eq7bc0HSnSzuJk8vAKntLfK8Xr+a4HPJjYIKESWIhP4LJKvb
FNkA8nyUDwxtmOtNKprqCZXww8fqCXA+j9rm62pCCqwMFYy59px7RCoJTAUFs+8N
96Lb7+jD2UKl2otvwIZM3eQDsLX/B2JTIC+un3DkSBq6qyWH8D3j+PWAxIXJZl0M
yeoZhwSAbZYAQs+pqORumagSu3l71R+TAV9P1Vof/KiP/PI3ghv5stCrVkmlPgr6
YUPSrG4eaFaKKhCt0wIbESXB7t5ny4RCxlvHhuppfWcftyABVjIDazkP1+r1tDW3
YDsg6u3PipSc9NsHLftacIoojP4b9Ka6tINl3PCz4Hpz2VvAMczB/fX6daZEEU7P
Sxutll7YAkm3HeQEEigeHYLx+U1jeISXrLwbxxm91txtOAH5ngU2bRsy85AiPKEE
+qkPGtTXaRJPcBHE1195RPAnfE65zg3X8AwrxcJMpfDCajJbr0+FoKK8S5/dl8ih
ffAiWLlwoOBgq6Wqdf461wkUOZnF50Je7lDt17jTJ8VgVmfp48IFtuSbEF1HOdYB
VKyX1KqzFyjqFyfI58NaSAuJC06OZVLcNAK6pEp9kiw+B5KdgphNonvFSxkITZtw
TmIcC0KMbyi5e/K9fFI4BKntXRqNdB9tSqzrShA6YHjNlSQNbrtNEQvDoy3yhF6B
1UaIiAOWkdhNS0yMABAufPdFNMOe78RQpK3dzpw5zQ/vs3HNEMEPaftn/VoKlYBu
BDNtIzXv9mIzeaWV/g/0JoRjosNhiZg2fLNjdvMckTcdaQiEcN8MVD0tlX3gdVkh
t7m17YN/r7tDClF0hTWKOn953wA1oNbiLY5NVcf+Fmck16miwqti4kX7L6zzgm54
pAIT30jKrvYMDXYxwto/gHegZMeqLPb7MCgubfoG1ZNaDPCwremCq/nrJhNp/B2M
pECMN+xkD1ZGZFRu6ogcBsASVTdxydBzkzOmZ2OjB4H2eiAmuMixK4WsQSw01bD5
enoGkrgxHCJlYLew5VfM9V9M3WU5VONbsyQxv2DfEkEO9DDwoZWtYxXpNiC/KIHa
/pI+aQjlohtk4+mU1Wx4AUD4n44orYnLdQmBsOs9xEg6IFzUDZhHvEZXqwed0FPk
HZFaZGIIhhx1iwV0GqAcAFabQqg4UH4nCFXsFp0PernsRPyJgmXxWd7TLcGWKs+P
/s6Dxu9aKrKmVfGx82tw/KEZIdTi1mkEGqPAew/o/FECmvpo1jIRpKjrgWLGxcV0
R8Dtq1ayFUkShTTN+Pk2IkIvZCfet/tc5BPbaIzBbj+wY1JI8tHW3k+z+RIs5PBL
Nkq7Sf788Aeh2823P2Zfp2PL9iyPdqz5qwK7ZnCsyvX/ft9dddpvkRjx9Va7yary
Jk9vMiTwXna+Sdy2SfmT1hPdRCXEQXeLkLKKcdldEOUU4fdPgf4XXWi9xMJ1W428
l1dDPpZbDu92dwQJMLa6N1ntkMQBmyVGGNlFagbQL1O6iPkiA68q5EOGfzzOywPE
vVBXCnkkSc53c0I1SULNxgxpYxHPbzr4DWdgy0mJI3yaQFhWV5RYRL3gXw4RgIrA
MqaDwbwJQbpePYm+DxoiPgy2JyhPK6S0ezlBj0E2gRqanOqaOahDNeHJNhn0YxK7
QPJCU42F/LZmbgr9T14R29ANse+Vl3Rl5y6Pf3L4LNMkL5uGmwHQjRu4kdFJOJwv
f77boSDFw8mRyJ3q+Vnhtl8sKQnV9zDg5/vEFUU8swRxB6T4ZmS8YtYUJ/p4LF9j
aw7dxXxBHMQlzSfUZkT3TjWVk0go2dk0MP12yXuoio6XUQ3lHNn0ZUGJf8NOiXkO
9n8cRNId1YNS8IWLjCfKFHplLehWF4Y0gqJngMISr0uW/xNW3frG9DYd3bMrYJIC
/z6giPHPPyjUyHW/c6YjMWsFw/tC+Od4DDH+h+qHzgOwakYhLi4vh7qi0INLfuaW
XoSJKfZgJc/IuEE++ZogkFSL+jDxW8JpQNY1obvnGEQmWy96DngcKbPOIOqUGOQ+
oE1w7LP/i35wX192djfSY7EVcr2dVo1jw5mo+dUJPK2jtJj5a82lbgn+nH7x9Dh4
EZj46Z5/IAjWXe6rz+9+quMPQG8N+sTAcwWR35wDF8iWMn/CUZUKWhl7Fpjsc6KR
j4YZfZ6u2+GGFO2up2sPCNiygZlgqDeUY3tP194bO+q4OyvPGn3bNpL7iLwinVTh
VWTVsqPZGXBOiVNIkdkqKRtitJ2wntwYLnV0o6Q4ziC2ib5hYuk39SGSlnX5/tIg
nGN2nw76VO2GQpuH2Qxhf8qePbRaKW2tCFdJ80xpCpxx7svUZWXUabc/R1xHprDW
3IlVDVL5GH1o+7GIlxakp9YwDaGma4J3TAVOp3R3RQT35tfTYRlkD2xywNPybq/J
pUTm+ya8kckfzEQYRiuyKd3tVwafxpgcv51694UAk8F51dfspYaT8vH/73MPwFuG
fS2lEmhMHNmlYbx8AJ1sT3k6nctICkIYRYAoVnbeWYkoXiUKOcDFJ/K7YriL2FdI
hh3dMI52c+ouSambY42J4GmvykE2RsUs3DJKUa8FS+WMPMqoPxk713augSIO7ENK
zd6QXmrnqUkDIcen9EENrkwJvB2RCsKjmdhfrauXIr7X2f5/96wlrLqKc22bi5TH
FrYrLlkaGuuDD9hdcFinNxXyagp9jvzjh+sG/FEiYfbmchdtvKGyTXN8KPxwaqau
8INFRU5cowFBUrf9BU8eR5hedYu7Vj2j97dQEyHhmCQtpUYe3IXIbctKsPrzOHeG
ZTdTPmW9JrPyiCLVHXrq/QaWlpdMMZSAhqAVABMxs5LDl68crhA2KkTAzjU+JBJs
LhQjTqFMuCyQms9u3kfVgMUrbRCC8+eNqezXeERcPuyqunvkUuSPvTnVAHiKHtt/
Uhb1AaYCvgU7gl1nJ8Znns68CjP/iSzUFeM9l4n90cxi1S6RsdIwyMiud9c+Mlxr
dvn1Nhj9LG/tmHvwFByp5KBFDEKHT97/hev2Cp6GN1yDVHi8SBwJJI8HycLp5TLv
GhFEW2GQLfsh+i4bJgQmVbLHxWX7i5LqBYVWQsEk3Zp1N7sLdL+Pa264ql5nu0KO
v9rcU05KkgOPuWd3Pe/tJ9Wnw4B6vhMUM1SCUJhwYsGXsqPEb8sMvWOYF61LAgVu
13U1VlIbY2bXucjEJ4MYXc8Ag5iFGe/0oLAfvS86obdPH6nSclbGeIM4xFabz7QZ
Ke/PmPk8CCICEWrFEK8SRPUHo5l/qR2eFM2zIMKMX5IOvZ4a7YGSCXIiSD2AHXZ/
BjrQ8N+CJNB3uekp1JQk4A+oK/JIEAjVSVHjm++Fr1ZaRD5rp3ul+Ius52YQydey
cG8UPH55WpRv5TmQb157XvxwQ7mNuQppftSEUwTmqSEw9YtArj7tPLn2BdM0V6EE
yABcmrvPfOwrtE5ZYMrzZ+Z8Zzq3nAF7uV3IC37CkKkQAg4OnZhxibf3j+gp4A/d
OWSPYUvbPi1Li47gDBJswx+TWRKKm2Q9a1GNAqQdiqu6GvmA/pWgaAuo54634/2I
gzqaWruSSHOrECk65A3TpnKD3zmtTq8jLsvbcQyfMDSDs1SravagUFgEEWQFkQ5/
cy2dvcn0xYYWwtZNgl+I89Au/Czc7yUbZD1rg/gx4ec8tbPKtUs1ezF8roYeFImT
juQ9Z1M9XFcRlv8zyPfC49C5B8OQ3nag69debiF1C9BG2z6TG5DycDDRVKD9kYV7
kFiEnyEha1teqU7d9HQLYsqd9X3MVx8vx6PT6yf70XXU/hPNjf36iJJ0j/WLlHR2
MNoDuARHAosgn5gFcCuy1EkBgWQxFP/yFhONH0wj/QG6jIU1QJOBKNooMQB1sqpq
pPESWXlT3MQWCgX42zcVrau/sRUBmvUa912Dmo6yYtQSlSjXuwlqjEMN7NCpONnB
y25PNRQtmZt2mmbwNMvprbZlqAHhbpTXplV5cZydMk1Q0MfrNh4QQkrjnYIkL4Fc
pSFuTnomNkXZJA3cdxtYVwyHRi+p3OHjn2XV4bWhhVV2/glCYH/H7/LNtKqYU0jl
wiSsy2WVzTQb5CQ3Zj2zRudaWLl5sp2mybUx094h+OW1lYRLgkIcHlae1ODglP2/
GIYgmeTQgADK3hVAeXDRYNpos5ZOtSwU/g8HEb7GUZtt2R7BKqznL10Kts0Zm1X/
t4LD2iIPe8gVq8VW7xKIvZsUqxd/AGrkwv/8WxgovlHAhCg/+qVPzO/P1rW89FA1
BFn0I5TKraj7pLCC9ntslU/hmku3LMMLYtBOxvze/kq0EZm31dUMEDFhuk5bo9SA
0iVUJLA86bQn/hXCSekqfBdi2S4OtZlNimrZ8qaR0rNsjDKaH55lFS6L2O6bTUCd
7bnBBN0NhxZl3sbrNO8/Hhb6LLZya8hgU+mF0cjxGneXqN/yQgI5ApQhzv+WpuDO
B3uupCoD4kZcy0wDsejIg2Mjjo4dsKhj8GWk0UlPe/N4C6uaAHrioNRXAUDUFPld
d3UgPJYoqSYqHo1XMzry5x6FEkLAPw66oRQYIElT7xHYFISJt8Skrv5LP8UEAPYY
wkYUBmk66xJRnosmf9EOm4k1XcLsnHAxnApPwd0nyrM1wGajIFBoNRAM+XNC1ndX
I5aEty4wKBtA0vEyZkpvRhheKi2i/r0CdGoxJhOldedmcA1IIq4MZEPd0/Lc83xg
sVtlM2pX0OOkvpZVYdjyyWBqHti0BObuUx7/DDm153bdQeFsOynjiRjPAETTR45q
gh+mAANXAGmoSi43MoCBdCuRqyX/HePYdcj/akWmHvCoFasPEtU1K/m6/AYzuaj9
LKnSkMLgLRXr6bbcKHKFS4ztF5jkv8AylXOyI9ycjzUyXEsSyUOcAOM8ZWd4RNWz
RujirxLJuqKm9UQwQm8nWGyoCFPrI7/zS2XoE4wKvRzSfn7/BA7BtQk+3/FYxcbT
swTEdPc0oTbe3H7aeU1GhuatyfVrl/vLpZRd57O+8IZOYDxkxHxMkJS/msbd1azf
jckr0tgQ1wAujinS8f6jf9BKe2CCWtVLwJYSeUmqwRF9q9TC1Tyoe/E6CuOX61Ui
Rg+Fs5Ofufe0zF0JCb9SO5QniUFTj8uE1MVdq4HaqQ82z+2IJO4ggSPrXZ+3UJ3q
GAZy+WXRI3XGgqxc71poLETnc02bpHNJ6CBoffq2QfzLD1cs2RWC+OzwfKnnaGcR
tSnZKO3vL2NfoBKUYKQ71Oip+SzCOTp2jxzm//ccqpMieKcF3HUzPspvVhahn7gi
ooVmXoz/lKNyZE2PLuNmTau2RHGyEooZMa6q2xyJ/2xI2ImK6sZDxZHX0cRHtOWl
s7bWeX6sLPSRsSs0yVWiCQYuen2CZOPLMvfsphMh94Em25AnFAaA+yT82PPN6AmH
HQ4AxcNAaNgJh2cj3rh+31vBaskX8d2Yg6LNkBjcwrfVTeSLLVnrTjjgYeQGeuFR
Iu/IFX0qCaPRzQrBYL1OrqEoWDe+1WlCmxjEDXJzZVyKy1Ed/mFxqbM2dIOxMHLx
6Q7ekA6nur0mQv2KiVnUWErQfoNLc9R5VhcgOqgD7T+eSGsGTIOhgC/6Qg+GjMSH
3rVjHOsdctkaKe4v9K2Hnd7mpMcVcsJjqq4s9IBkdNuC0+ny5TvHhCSvAYQrz/u5
QVVu1gds5dubUHMO2i5eOmKq71FEJ0mML1647B9m5d09yIdjLdEJTXaIbQHJpvUL
9v8qNJvCSsONYY1dppMTqaTERW3uyK+B6JJhHGZ2z1+3Dbzm38vethKR/ZPCHOxb
zdMIu1OVXazzbnYAkQPvHdOev8NnMeJFsT+hYBK+AgGr3EBbXmfHv6Q/QyaHmxLq
Wy+GpxVzbZYeOqtuEm0xp8bXnJzXLwq9n3J7wv53DpZgLp4mRSErzqQ5vMjA422q
JarlfYpdgIGL0eAnkT9+pE07lcfeeh0cRSABicmxKVWoQjnINIPbAyKA13FMMtwR
vPLpuXUkaH9oOHbfzIY5/nx7udvk3igo0huzrfUuo7rAHjiVl+dY6UN+vAesaOdz
ywPKTQ1VRZGwzIFk45w66ejJ8tXPAn5Ydew8L5iltuIPB3t8jXhFJwQz6sU7RvtD
yQ9keJpKo89q7spjwmHSIJdUQfcDi/OZfHIrJRX9DrmY8McJIcwZ7jA0yF5P2eDo
aduyJRErvq6+aqYu6xVDdRPTRJNZda+Krwohfk79EcXiUdARDmD5wQxtDN1WvsLv
8ahdHqrpw2R8s0Y8i3LKtsS/URucxBF2ipgQygKtjUhDJM4S4Gf1f7KLiYMD3C7s
Zi5x4EVKL4YLBL16peR85dsrsZFNK0NItji9GmgRCZYg9um6jvLc32VETn+ViLST
RDxyOh3pUcKeCDmqJDhXER4RuO5n/x8q/jxMaeM43KFSLCWWE591DpH0QZrw+QlE
Y3XE1iPfKBqBQICbcMirOloKEAjEIM1zCY5PvwuALCo1nqsDBBdkoVK3GW/mHsji
f/CwuOOc0BloEJoINBU990gTGoHfRdb+JiXPBpPn3gfvQmbydrCGt9eg4XEyqXbF
y5lFv+JItkexQjJzX1h9nJa5hAIHeX8wBacTyOp1H/+CRt6N4dDjHec5FJxdvPRW
Cjh4BKHg+X5U4oPD1mDQtIRm8mnT2SkOvYLM2iWGERxp0VAw24D7iIu11nAvWmLO
Q/d/gfV6+zf6t68VegEuHS7c+omtxLs/oFk4BW8jyEbnriTNQWyBFSsvhugp1qGX
VBaKZXD01JtNhmxZjhdxCwQf/W+BDmUzIILPbzNApmanz3eDw+LWvpU8mcdz7yLl
bvge90Q2KFk2JlqgfapHvcIbeiO7851atZEHd1zqANebLToz+QCPeI6ouWnDO++k
VXZ85O9wcuhGGKRhzp2oXU9J/mRDrMgGTHPqEgOaPesvMnqGM+FeH0bhGTcZjzA2
LcgJPx9kwY8AeqfhpWTHJKUrsqWAuHck+veLfRd7mCZkcEbd28Sq0IWUk2wgTXrz
4gfHL2Y647HMmTNO3o0cS8uwmUEpzBdLAT3afoVFy+4H+d4shAd3tr/21OutbSHn
rMhSydyH1OiHdKbprhnzjksn55GDBl5DuU0RQY0a8z5GHF1/v3FAxdtKa8aisDrO
M1JLBct0r4ibMV6HerSqevRJPNcdgA0WfglrNZrrlsGtP07f9JRHjTK60A/4l3/D
MZhiwccLxtxm1EeedVIFQeEUy1FiuqqkjHkITpxq93VtPOGRqJiKxLC4OIM8oY7/
Q3vLYLzffBQ/L+e0qHy+Rjt2Xwko81vckrOdTOqxF/rx5KrGTUUI2VeDJQ2gbu3y
ZjWnDXDQSxyNkGn5p+Ql6VAlJRIyhsj4w86sFo/WSGsALDDugwVGjiZdikrbnPG5
wgoFa8iw5rL2vVbn2YRaW5jzv9qxSokfaohkwh9SdpFgpnC6w3+WCKYEKsZc7/qw
etn4giqOg8fE//bRzb2dLqe9tMYtS0I4Wh97rAAlb/DSckv2uwOAbH4EByJnOSDX
rERXNM24Y2Jt10zZlCFDz0KvWGR7W4uXmalo6JQhRZx7bX3sZOnv2H6+vbghyh8R
/etuactmjeiQZowixKseIzfQt94oN5iEeag1katI2ObX7v8U1ScVvs+TEEwiC0eg
vchRaD8lIsoIX3vR+Lbjq1UiOlgqs3QxJxQPXTcxAQeeo46j+nxgQF0dbDUEfD2C
msbcRyWjAQqUXVNuktPlnP9meJQ2s0YtpjQTAZXCcVyW3pBn0ykZukzGPxa8DYNG
OO4ePkp3bOFtn6qhYLRHwe9X50N7K7VVqxpIM/U9BQCkxU11BOkbfQWfFAmx+9Ob
8mMdd/qh05Jnho/U5U+zHT9MWUwcJfqcfmjIzLAX3vM1MmK4ObGg6H+TSu/QfHcH
425ocBUmZKeVDM/vWNultCylofYrXbTJYrSgR3cj74AqYCFgHjl49+ZBty++oTLn
wzYcJe9e7GFS0xRMNefNdVLCiNe/gTvHulNtcY1jr2og/bFgfAjNDyC2v3bgP8jw
5pwSNEc3gRysmrF05G70iXVO569alsP6nqGHa2WkRW71D6P+W3U4cfxBPSVPy3P6
PxJNrsk+zydnRqzRk9uSIukw2IHYOnUU6QwaKRw7DQ63aJZajTv5X9gp8o/LGqmC
yfXiZyEtQha6D7hSYU2ZVufKz1SxHt+uCxseP8RkiBEMbB6H9zS5ek7gE3Qz1+bU
DgNykRvaVd1ccuARD+8hCakXU6HV/1oeIKCRlQnTcwyBaVsCzlF5xU1EVPNN+Qp8
uaBlEjBg8/lHbLOm0DDvLe1TAOLOhRBT27SHqhI4RltKkdlkYOailyyhcwGGC/an
Yk258G4jWS7A9Z53x7LPIZw71KFL07sBJPUo3USYQpwd6+lVAphdiEkaxj7E3pX7
m9VHqgOinXDnUSAG933UL582XYDhXQnHETcwConhGOQCQT5QF6i9UUCOs4HH0NGM
AeRbX3q3izlGgqOgGETLpPItE1i87JRuik4AOpN2JtsI5Ah7ArRYA8R0vcsW0Acp
wuXfmw7gVemWrWfsWZ9sYmHxA4RQI3LAaJOrYPFcAD1uwGqvel20mlDkjabxExXp
nUVWi6a2mZ5gF38rBtzePVqv3sd4366pok6LtKlQrDMtr+9uwMHEhnG00maQg9TE
jZUB9Fc4+gkCft+2I7OM6WTI+Q/qBS9pN1PSLOkAfI7URaUfBvh09NoJuxpozQll
1f3tNKj5mjeNrwNQEMkRBy/E26MSo/Yzc0QxFIedI+EuXAIyvdDTI/CCnWho72VZ
pBSzK5G/dKMl2xEn3jdIaxSX9/R2PwqNFBdsRsEczC38KY0b8tkQ4NC5zU7x9cwO
SNLPqyRSyOupe5DKJ8V3jMihuWeehdfd2GNhwn/W3I0AW/t0OWhLBTOcnJ773eIL
Eow7uRhRlsZZrQFjtR06ChHGrUf2Zfhck3YzMP5nO9hvFXF0FRCNmaLp9yrvki58
eO/HnZKmz9p8Nxrrv2G8TlZHo+u4fqvNqMpFrdlQYjAe4fwzBbYF6LU9MABGQSS3
FbSCC6B6fz/tygp6BHH3NGJUNo6SaYd4KpjPxWynZZmgCFK3Y7C7Leq9QzPRXMpz
nQl0CCJ2vND79NSDW7W60qwtV0qvcpOO/zi0/g0fB8hFtNDzIOHdSSZdOtxYcTMr
7KonOv6hi7CWpXcn6FHWbN+y+Un2fx2pIMzoPph0Bb+JjKHF5KDAPjJqCDYriIRD
3UT9xqwnj3QxJcPjfT97yOTjPgAx0bpFdJJg+oM7H8vFrsEBjQl2dCEnZ3VVKSYd
T2cFUSWnirigZnh9iuaVypB+mSU8ElKBaTOMae8on0VpFxYPB/6aO3sdcl7Rm4Er
S2ZHOnF8QNLq96m5c7mqWYnhUKNs1bzre7dySC2gDnc7DYacczlf9KB/GZdnGzMk
3OMWDF+GqgW9cHHkJv3BxPVXG579BpmAoeTzxeGFd/WE3ZdaF/8EgXUMT5HMnQKT
ByMyp5EmA34Cf9HCJG2mmtQjWz3KD3+jcIrF4y+EHkHYAV1K8PYYqhIJlDCwovG7
ehDTVkVNbglkBiY7o/BDjcDmdBgUCX4yy/t0C28QTgjDB45p1wph+0wrVBygekyx
tpUlxU1ZOVGot7omWv1SqnRZWOgPY4u/c/kWBTHwQ2SgtXOWVUNfWHPRmXYNgFNO
yXlTD07wYhbogmHOj8mjYikTRz7OgEoN1LH54+PXzLSdWEqk+PR/QOMTPwXB9B8k
79bvtCfWXYZaCY67BVKKniTMA+FS7802Q4kiVWqYFnmNQRfeMsJ/f3k99kVvxkR+
8LmSt1tZC1PZw2O1xXpq22I1ksxZPkNar4dNWXKEs+icDeHrG9qVsKcTZ9P0Az6U
++ZO1lDQ3vToviOb3pClxnywOM+5qn1AUuj/jyTqEs0AGZPhx3lRz3WsRtJpPLZM
J069n/9eLnPFGw4trCyWgyBYjf1RDoZ5Dqq2M2HePjeD7bQfW+Am7ZQNwzwvLfko
OejK5vTtJA9pVcMr9HFK0nyqryPuy7mhNnHwzfg1gedtVcFnGBe+kAewNaqDSLdi
zKcFE0stghEvo7Gbecj6SXm1S/u0W310Ve9/PJjicSolmXGL+MyTB9FJ2iGkNOff
0Ho95NU78HiW2IH+9MSOXY+Dmbbnrz4/cQa9ajcu4dJeVBCdkD5IAnzcrWCxkGo9
o5uOiNdsN2TzHaF4+vqQOOl0EH5TUJPpRJpYvVzxgtlMNVSE0H7X3i2HintCwG+3
Nc6eVqFwh+QFwmBTqUtQh+z4RKkvcrMLyblyH8zOud13OhUUUm3cN4BhpZjT6FEE
ufIup/wfVJFBg8mNSjSDTyKCrc1tVMxMnaD5sxjgAcx8wNomxK3b4cCoitPqlPsg
hvLx450KUHPvzPPj50hvz2Y9Ao++HIAWT1OT0JrqWxjsddOrdqPBOmsDiEQtbC6o
Pd1l41VHmOy7bBwQ7CYhrypj2bobXGwwOm38bsPMKCwO6pTAPUonhmMyS0IOrTOm
DwFdQoM7sQwOW908+zz8U5opZmCEdLqEVEBPtP6xKXDQ3DKYRvkvNqU5m2Vw7d5T
sZWif4hU8qF7KXO235GezlyXbGPmN/d/vkRY4+D7OOK9OrAmgpuL9cjXX+T8/nfD
YY/HmP85gBWERpRN5ixamYZlak/9ge5Y21yIVvgb3XYBNne5usyh62QwK9vyN9IB
C3v1xNLC0FV7fKLSyZduQlYj/Occ/k5h8ZsulJAxcV6sEuoLUWT09PohBEfsQfN9
+AHGn7XTX34Pz2VUNgBHwUL30a47zLkeBowKzzmCqCYlMsY/jtOCbi+TfAZrKSaV
QogFeH7cAUQEN73HuWgqIqxgCl16hLLeLLm54226bq3Z5Z4iJQ6ieO3jACb7nPC/
ms6vRjukzqb7fZ0cOB0aDriobWhrAUpUUCbQdtruunxLXcu9OqUrwrjfRqTrE2EW
5WhdseFTdCPmaKqcg7kuN40L8BO2YoXHe291Z917nv76mgtDFFKCJPZYDb98Aw7k
AGHBfpO5HWNwBItuiEwwNDhkh0/44kkr8YAk+MMY9jDz1tsVjjm9fpWAtLPWDWWk
NFJ8kyKiDwP6gQYDPe/23CrKX3P2LAvyHEI0DQGghKcW7Qr/taRfllsNCxlSMpQC
KgDXDfoTv/qT1dALDIaHtDev9LEqa3IK+dpe9f8nLBV79T9SPOBVqEI1JbMj3Pkr
4usAhsbq0mBkDVwZe6CAMOU5OlRCdTERHOv9vEH6gfuMBGnH/T+LEcXKv+NTNtFg
SMp4Oz2+IBywGJWmlRGvlerwSOzfm1sxmgsjnVqG2uI7HJ2tXffPXnaqX8VyFug+
KytV2MCFBjYgeoQq2wFoxqNARnuYliBLOxfiv15M7ZjhcRwYc5MhQMdavOjyO+Pl
nzHVu/39YRBNDVNl/Idn4xcrBUvGmPuYKOxpEzqFHO1ua0tjWgJKltUsXGleuc/P
Ep5K2ODzIdf9ze4cQALdXqssmVlJy4+6wUQGkWN3SLWM+rVKmsRxcCQ/+IKBc4JH
PGCntvUupMsuPbv0L2vkZigUeC0xpKamwEMeNHHmW6DwTzENNLkrKIiFdV1iAb2W
/KkgkTKQxzhkbY8aZPbT3FLt/7W1B9M1flrqSvQK5qHP9EkqGXrTDkd2Aru0WRpb
1MkKGEy+3ud9tbdKYPQa/uU2qfdlZtzaH5C91r3ym+lbHDbLnzOTi8oFn/axmb/Z
SbiMcS16Drkkoooy6u5BtUgWITJ5lJbgPQbdcR+U4VCvBYwyRukZqXQUYNwoKo1H
d3h1JeqnG10lRQ9Kkc+F1GsEFu+NKNcwcYoeq2LwtcoKsXUD3lPO1X1Xof3CorCE
/RslyeWoJQCrMVStRTEHxWkzwvNSukUPgI1zsBvxYbNWEhmiYB90swbPRovwfnIC
40Lhjj0DuY22oTeM8ETCd2hkK0yV6310rq2J6t6/NXYZCTm9r1fNX2A0ZWEUHSLv
TTnJEn926P8oiSCWubOts+CN4SPQKi0d/P+F7qxAVuepwHr1vXiTBk9Xys4EECBm
TXEodcDnbeVU6KuMmAIEjK+BxTR+HOREfw0XhQdGYEaPIFi62FeTgAEvzly5nENB
766QS53wtUgWvO3H37tU/Zg680z9tAPJ3r9jVp9aI4+xMEmdZp6lamKUVPDyAZHs
fpJgqcv+cfZ7IsCALXbuGNI/0MJeHN3B0aE/7SaFUjmtj6Kgtxcv2J6YYAbaoy7f
tE24lKqyUVdeaPO74l4Y4PX8O0gJYNtmdN2hVc/gMwC6eYHW5oKQG/My2Jrz3Q4w
Qg/fjWChG87OMx1pxneLHl8/d/XmrMENQwb5Qo+EiHQyBMiel68AEc479wnvTYMx
JkntIixfoFDgsv3iL/DitsX5Q9ZBijT5sXx7XQPIDThuTclaYSMod+50XvSKRT8F
A+n/Kl198S5PL0XXnrXAmBvAt/K7ZdYn/zYCGf1IdzY=
//pragma protect end_data_block
//pragma protect digest_block
IEv3mHtWQySJlKAwQmXKvO03s/I=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
x/G9xJbhGmYuiBLI97JAmDnHAT9bH2NUlMLRqHXm4Sa6PZo8A8e0AJvizjLDp22C
8PjGdJGD4kPhZr2fypq2C0B1q26Hta3l/qPmcK9AvSuPozPdePyAXkVTqExUUtPF
EMMWi74uwIUveR2T0pqK/yu6YJtE/vBtiAlm9wrpAJKvEFfdJPauGw==
//pragma protect end_key_block
//pragma protect digest_block
2vUOyGa/C6HFEc8E94kKmD1PYyE=
//pragma protect end_digest_block
//pragma protect data_block
LLbKWS0/eQlumsM/dEM7o2ZcGlcz91zl6l96eqR266dTlsuXjIN5OcoiZAqi1k59
EZ5Z1XiH5+Z/0PryfFO9Opb5wWa0aJUWVqwPaEo/9Oh8jA3xjdhxyWvDWuhM5yYZ
X/B9EsTbohBU4FhCaML1cIZlc9LQ90EJtIwrX4WlA6Fa+hbnM0ClcslHwo21Vdav
DMVakDo6FB/TgQ5vGIXUIjky3p8PO6kqYZ/Z3oauMeVDikBaOZa8YBMuPbr46/QJ
iJhoPon7fSQSq5UgCM0J2od6Uq3QIFkN8c5i5hnC17kh3xG0d6gEEOXt8HEDcf4C
3uEXAXgbxYIwCLhR2C3oBRUekF35QMqXGH8Gm3X/uZbyv51zNRPC0ZPKm74E7GOf
z5qeoxQSVHkngzpE7FcYAg==
//pragma protect end_data_block
//pragma protect digest_block
dzfBR8bMWdBSHUuu+Q3dJaCRZXM=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
EDlEOA8EAlc2ucNVkOSGZD0Z0WKLaXOtHp+7nqnSalcZD+zK7hG78RL0oAxidFK/
TmJNfR7v0+Hkqh1PnYx8ggPo4+NHhRq9GtgdTUaxpOZ2rAP4DB9E9oyhKQvGQ3GC
8rodg/73ljP7hhiPwmtOIDazyCfp44CecFQVSn0cQDof7SdfrWCEKQ==
//pragma protect end_key_block
//pragma protect digest_block
4t6I5c+SGjtYtA4fgH7QmDTDGxA=
//pragma protect end_digest_block
//pragma protect data_block
ApeSUteqL3A6N9OToWFfQ9R6mgEYNANiGzOLgD75JVHBUMKFQaaOTKo2DTvHf8MW
a0IG7671YZqd8ibpnCXK0MUpxRyOdEFWxfW9hfCy+XIilNG2jS/VCiUn2wCa3lAE
6XpBaMRaQ4c+5TfU+SIl2xJtXdp7rm3KI0A77SJRM4+bkToFZUhHPrSgZsWy2tNZ
ap6M+kJEB4CPpBmGZEzyWyFm58aHqJ6F3uXl1Gh2rYS4g87a3Mavgzv468/ZB6Ea
wVujpVvUD4x2qXmNASSyKvWvgTfAsYx6QJcJudLFcX/0/Avhk8gBdK3zZA78NG8G
UiZr3eYGZfEYeSEpGDju2tr3bl0FEoFomGiHiC3rtJRuIP3g2ZoRlnjTNG6enTqE
MnSixInFQ5sI/rbRctD65wsWm9TKhdu/cIOf5MiCws4teCNGdfc8ZdpN49jImex1
/wXqYly701JaaVtNlkJ6+UdfWV8xYu81gjAaJESh0pE7FZ1y4HHVqKeL4yQcuVj0
zfPhdeI7DoOI47rTOj+EPnBZmU7b4HhPVZU+0mduaRGtKcPrD1axffB2bYNK7rec
2fIDl7sh7ttGhoAxvAgI8yi+SSlGESpWmDm2k9wK/227naXTa7ABbScyCe6IvDI9
GTSr3b9a50ntiTMyCfdcMAL5vWd9CA0HKyJCDigk10d+L8ha2GrdBNK1gJdFSUtG
1bfIp+LLzZGYKQnPrdu/Y9QyCC7eoTBdS9AIA5rjLcI3yPr5vvSe3uFo89qFlMvs
ZRDFHKuc2dlu7QlgMbgmNhVE/S4ne4v3ToPLSP2WhVngCz4C3Ki1PeBAIsRnbNcs
E3BxXNYO3aQr6+AaBsnvTDdol/k1d30768uyAp9B+5eg93VeFv7tgcgviFhDJ4Is
YPjRiZ1j5NTcwsQxGvnbeqJhRN1BAmP5FflPQuWjRHQ5xukHf5jNBOhqgKzInVLf
RAXXsu+YgEOpSctsPLd18Svj5Tc21T9V026ZQ/1Pt/KKDpnwaNEpJ/V6Y+k4RMcj
7sBrzC4e122mVnlHjlTZ6/n8NDncWxIVzFKNuquP7YFMgZx+2gELuTiQEY/dsDEV
70YGkU0GQ6+erRV7qm/ICx9OFxP0PICRtMsgNFtGuEbfP66FIEttLJl0Om68AsqN
h4hbzjqMNsea5Gc4qIcbqos5u2fCKfVPgVxDII1cYRKm8LO40Ukzr1655SzgbUDP
3CwB4MSZB/2RlwnJ/Fn7NxNMRMbdlWB7TYSczUTcDTRAzmVjmYkCBMyCEqaCe6F5
Qp8kJISJYrnjcvSCycdKG9h9LmervHKS3W7IvDO8ENX3pGQYgWx0U5lOS4rEpRtu
I9tNlH7zfPiv0nGyVOIEKaEHyt0VFoYIzP5cssEOuOf8TJw8BJVW5ek/ss+ybXET
umJIJgXzafHDeH1YUgTmWqofMoV+Jygj6pdCTiNCnYrGwVqBaejg1vAqKsCRmmq3
nDFSHkZZuTSf90XhwEAO4Znhqjm3YFPhofiZ9jy3UEtWUuLmv6pZ1Kb9BRrrO3tN
cRNh8K4aiueH2OfaeY3/f1Y8oP7E9Mu36GRM2Wr9VfEI//83bmJaeitfT4Dkkl+S
gR/ksmi6q1s1C41wPhTMcj/WURxuuBNxBO6UmFYy/oTuzu0kr3x891CkpGFuyXWT
lO/JJfMxldz1XMFs/Or0pO936iLyaUypYTGCHNB4uLBwD6MvVKx5BWzluEQph1T5
ciRV+5EnJIihadU3LWcfjvwxRBKQZpvBq/hoT0J9JxC9nTFEdGAkCCT5WycxcYY+
KmVbiSjrFzr2w4MavPOM3HDO3jRfw++aPIC1jvsLXXkGHKbOytm3IzMcQ77nFg7M
ttCckeNSBmuPhVHdlDSZvaY4ASvvFU/jFFaN763ENPFB8oVB8r9TmCCOMspt0Stf
nU8O/Owt1sIb1I+g0RLte/OofM5FIEA3QfZPKO3cz1QU482rqUO7auKluoCl2qIX
Z2tC4uezu+wNgDUpeY++jx20RE/1cWTApGr2bCiljutqqUEFCRQ9TSh9F6oPnrjz
Sj5HEIvF6jP+HnvZ09bGXOG9MYjaB9+9sWMUHitFkh9Le2OiXwIpMdgurH/OeWuc
9eHnHsEEuB0c/2cRURwhhHBnJAGAUNsVgTDO/j8IIZ+W7W+EHLY79uKcxOIdLaI0
YUo4Yy0m7kjPZMKOdkkbIJ9olddU9dfVeFUmrKykdGe9U3jZ5KKIcyidE6agOAqK
a5LfY8fssNKAk606X5iKUcpADhrx1j6TJyV6Usqt81za57ySYYhK1GeyStmd6nTo
uwjuvJO9zKIhRiYEw+FSWV4I7nTUHGw/kAfyZ3jIkybfMMiaRsrTTBbmDyDqJI/H
IHZA0mcyPUnDgiVRM4HGfAh8/tGN57qjgnXe2ZA3PAyS8/aZAvC4/GGlkcz1P/r9
zJ+PG22BtU7YmTIMGVTZ8twWzt3zWJuUBWX9xhOPNYV7bdhHDa6ngA/Mnk9YGrwT
Ngn7w/eUk4gVKwsxEqZPvewFbMrjAp4vaaEUM+cLvAr6lru+cLtekhWYQ3yo3/C/
Zynrh+Fvq2l61HRCLCKQKOgXAz0bm8odpDwxEM+2SG5xuSMbdc++2X/iSCASZjhd
Gt6S+5u7xbKhr73CAWn9nvQV7tlcsqwFPPypbzgGVuv4pu8/BpgTYKV21SP1VNW5
r1wjehhfhrIC1J28yU9mIlOGV31BE5+CSrxkvgGqkAAszJMLCEJfmVm3c1+9GSc0
/Hv4QRUSYn5E+qqGH4dBUzt4NTlEk2F2DgtTmRKzJRYszaQXWoj4bTcDbzrZtPbT
NyGXo660/FxDnBU07Vy4o59lM1Hef7KvFQLLL6e0ieLbX+tpYqsdkWEkoF3qaOeK
cbS19mNkuznSv4qbYgsPAHUPkXrWP9JZwdbB7onWe7F+WacZGeirUO8ml3JvIguo
2o6hxh9Nn6PTSsi65jF6fY2Pz1hQ37gaLe2LFBnxRShR13jlUny7Isd9PRbLJIaY
DT8PIH0Vov18NrjU7DJ6AXcr+45lMu6LnTE4DXXK9oHb8HFDBnrMPPP1ClhuWXqR
7EQJLFO9V49SH2zqw5/3JMRsTw7/n/7le1Ty7Qsox4BCBOfpNyeIIDJIdCr7zLDU
KxQXFoCss+srLj962+vW/I+K6/wJabzEwE2rXhmmyCmqDHt3fW8GS4+O3IG+5L+C
ZOyQZ7j+rUwW43uvgFen8a2UUy9OtrEeWbS6/JWn7rwIfMSgOY7p7MKbhU1dIHNM
C8tPcc7V+QS/InPo3gDOq97jROWHZr8Ul4JbyNwokX3h3cf8a5175VSxkoJOqqnc
BkhjtJHsia0RBWnsGCtMEzQSQsbAU4uPgL6ZuOsva+5q+rI6VAcdknnmvq/utCUp
qmPWM5U0ucZ3m5ppqqZ/L9+YpeGi527esz8Xae5pIMHROWIpEFV+OUL85ZA28g1g
5w+6KmJcqnIUBLLuKiXAsv/ZP/lnp1yFJbGWSmhSmtOmpmf3lTbJMxgPV5EPeeS2
0LZQAHfMeimR2aOKivHFwqFJpYDDsbHelGjFgWfb7xG1iRBnuKJL6XwU/4T1/tu3
TlrdTgIrKlIvTjrYMxCO6OT2WVf/EJdEyhoNRDeqKEDQ1dVI4z+SzBM99LMHo+ZV
faqJ0OxgvLNs0wKWpH5Rmf5Krh8fJCmt+6NErRRc/eQvWz51JHXNNxYGgtw41NUZ
/er4h8ZCJcHrZkgRQMWKU067E2k6J8uTpTZKpcZk2SJmHsFSwV9OQm2qUr7c3/ER
MvfFt1SwKwrPjyR0jcoYtuxazOrkC9StkGz59tm0UrvyDYBatA6tiAEEe/Em2ZF8
cRHOy5JSQKny7j7ZwFE9XdUMWUNFFsc+2VUH16UsOzMuTej7+nHqiwoUI/fHLtgA
XFq5uTtQZyGmL//muNU4wAZGUO20nPVQ2RG7/09m9kHq5WxkTuZrrxhXE9+5DXS2
om1P/r34i0HyL+rJG4JiaigaEfePMaARiXcfb2PxikeRfOeybu+HvKrzDq7fMDqA
2IMHKPtLddn8Tk5QOPe1k5X2eS1jKPZ/ijjzUPhQz8m9qmKVtjzTB8LBzXqD3cZQ
fzeU9zmrc6nWihIsKc9g6F4Q/RCj2G1VNds6zShYRsggwBofBYsS/fzpiwwRWJBV
cPcPkYD0Zxbpwdd6ZrWu7uAmmLiC2e/evk58WjHm89yaCGWovuqio+o30l2HJbpS
BosnMgcQF0fNn19x43OnlhEDXMtdkqc/7tJPLmCRBwOqsgrPaPwTIpUr4dk4SpAH
hjyEcbNAoKaFhVvj1PiVvSNKr+uzWgC+rEFQiEtO/8M4N+8yGKXvJfC/5VhCgyZM
4e1HAT5rmDCokP3VlIjhOycT+yzxjHzx9q03uW89z7T2uHQvZrbITQkZygZR8sWQ
jPgyrxipAH26WSvJYjvxEL7ccL99XHd/w8/XY4ph9jyIVMwCez9o4RfbspG4Zouk
77p3U/154ANs2kY5RqpmfrUcoHWNTXPFxxItLZ2YbEKhnBdDgsrFN7pi9S/xhXIr
xJ3nq+zc0s0WozVyzUdJaDhIRfJ0oJ6dQyF4pllV1aNkKnqZQxLLzs2q2+1cxysp
RtnZEtLZ/Go0JWwimV1epYI1ZhKf0TTeBTiVxydR/JBaJ8vKi/rm1yZI3qP9OkqG
uCcOcvy2IzIyeMMx9PgIxMlZLKkKS7KxwbJBlI8PmjR7LjtSL3dD8j48sC4nwp5J
Orn/kPQqfypbD0WaUUZnqmUUyAXecq2aSmGqgRDqxGBe3fuKSXr9ZNKO9Vmz8wyR
xR8xRixkzQpyJBX7fCrVMmhbo6J4nW3DvE8spePCYWrDBAAfE6BJtJj0S18ufqHm
lNUhKmrFBMfeMOAa6GtaN+XMF+FmzvVPCuSc340Q5iRHSc0oC3jbyLSTljyguc52
5flSIJAInv8zj2AiOo4Okx+Bg6IKp2fsG+hLX+UkQN0uT8+v7mNq2AfLEh9YK12T
PwdGgaj9C0jgLvRmOcUwjrUeHOzy1pXE2SgausfbCE2JcdE1gGz7sEwBET54pAWa
3vdK8y8pGflKybG39P3ujapTawoPXNAH3SHSmstommN4hVGPOt4ct1t1df01kIEH
hyIXunoDzXboH1SCk0DhZJ41E7/I06MQUBq64asujmTuqPIdGvSRbaTSq+MQNeh6
5e8XbeX6Qb19BqYTb8o2LJ4Gm+sHS7vjolCEv2H3NTUVQJY41S6LpclisIyPwSHq
8tLOPO2a2yj9UvT5NR2uehML6RDOn1Ot/fBd0c1R7FVyfVKk1plwYp+TJy6Bidtb
gMgtgCAPfDBpc0ir5HAZzH8AZes+1yjCynnBnAqh6Vc2OhHOuX9yoz/5zy4h4CdZ
1/4yJiIsTQ+XH/52AqSlxjWa7mem9G44vNjUGjZ3Izp5ZdO3ZkuHrryUSY4zJGwS
TSx75VuRs+Q05SWekJ2VDcazetOeIwbx2E+5CbLfGkaLF7DjPYXpuE1ea38ejFC9
7GIXn+f0VLBgPMENgHrPLuHoFvSdPcWRWOVLyUnha237+TIzW3ePYl8K5m30RR+R
cx04c84B4DhCoZPbS3+EF+4PvSOsduTJ1dkVKjTyn+FH0KdIkjGlgKBd1X3frinW
VwUqp4x4ultnxpfy8DX9O80Hrf2kD88B0sG6ZFj4lNyH4BoxWr00y+eteaKMkYL9
F86Ou6KHr22LmHzYKiTLGKnUtOqnVXttpASZOiRNk4T8fEFgrPDSOIWEO4egX4hp
cWbgkayajjUME3wBeWhnnG0Z0Dg6fRdHZflmVW5ybWUNhh7dl72JcpOfiFncx5qM
C1hF+WEWKDnboELeJQY8hKOYKuP/sLs2MsGNkWnciKVdt2FICaMqQTBTchEl/+ex
Ums1nicIip43VaHuKc76Ykh9NJ0LFulaYudH8zc6Xkwjp+8xTaQk+4PGEOntmb7Y
gQeyJoN8Z7sUB0NufShht0aiIyhxm3Eq253oEHy3AsruUlaf1iS4QV9NyCluAxXx
oxO5kWIEs6Lu9gdL6a+ry8SadGNDEm0ygrzsRnMZHbzzt8//MUMUO9C+28plV+4S
Tfvvg8+5FJdnZqKKDaUTdMLuODA2X5yzTRbOdkj+UteP41UBe4aFEDEU6jjqCxQ2
UJ6i/5pH4sOtu1BiXoVHHA/WhMZf1KpdSlLlKNaORFCZo+jmAAjg4YkTmo2+nnN1
aWWXjUGXNiKeMkTmHaVqYmHZt3SLJlaO2zCkWMRiiV6XwHk5TZSZdj2+YxcUdSv7
DGvhltmK4O6s9LhjfqWHyw8UfRB9pufXau8ElWNX7VzZWdH/Vg6hBwHoZRiSX+oL
xybI8h3SoJekFrr/dedxWj8ZuyeVNFSQBy88guTyJ52MisyOiyswgk3Ucxc2xTrA
nsuNRQgK5qEb5aiZOCKZHwl63X6Liq00hLi6lDRJFVOJU9SbRS1kPMl4cQ8O0OVN
NjpLPViRP6p45Wb/DVJm83rYEsbqkuVNiPJUYAck+JPmATxSjgd+idDsnTCwWpk3
QQ3eZVYFCp4tc3XJQPrKZiOifgPoGSXf1ptrkDuHRHZHnOYqjZt94VX94QoNUtFa
86zVEt8SWcDti0C0LYF1DwJz0hznBtEUxfTnyIjIXu4Xvlh3/JBnO4X5aeqq410A
UYXLjqMjCwJaCEIz7XhP2x+YjUXdCciiAcKG4HM0P9RjfVB5wXSGTjYD9+zSaYR/
NoKXUnO2K+3a2c8MdXohZ7of4LpF0vpGmP/IgGJJhmzOVY9yF08WtbJ0MTWCLUis
maUbNiUWjDjzXNM2FwJFMukDsD2zvUf1KBTUPK0JfUxNMy8rp2qxCQlPonKQDei3
OWwQAI6Bc7Gocvuy60SqygTNytkcHGFx83I5XEMZWOplEorar3TorB/akvNuZZu2
iu7mspfIzZCyrs1lWp+BL1Dy2eqy7Xk1BsQH7y40ihXIvt2ARmvuJpjbeicoymIG
JLVr+OvzSMjujkBDzh5Q9C1gBcb+BGKuTPhFeFYwPW6mA0LM0BA+L5gnDPjFSEOR
tQsFrF4sv0xdxe5i9j0YmAQe3SQFtKHWxF2nHV9lew73yzOvSUdM+DCOu7/zlfSq
CoSXT3L6Zv4Lp4U2+HYJNG+P16odQ6MR21So6wPbR1x55A6+8nQsLB0iRpiseml4
l0K0f3P0P9MxixzMt5jnWpqsY7WWqZTc5HmsdgaI0T+z5kstKRiZXnG/U0jnJ6Sh
rdInd/ArCTtD8uMYeiIr0qSeoqRtQHfhf/PVobOOaR+VZYuZZxwnxWFLnhvoAsYx
jNkMe6TX4/Wia5rxBuQlIn2AvTOJciPaQQUks/P0ZyNgVBREyw945qyq20MimMzz
mG6kcJvZBVaJc7HrvLGsL8Ha4lt/x2Ng6KuIZ8UF6FfyXf12oUvPV9T77WaZTLYU
nVCHE+DkRDk+UKeAsgX1wOh0i1JHFK74OqyEk5FGaJHXLFzGvoZYcXbkKT6hrghx
m38F0naC0vF5w1hLhOJF8xCS45TmlVzycyvKmo1kR9gbABjPQYGc2OXGLLUzP2Yx
D2S2DlWhLAf4imLNMITXz3ebuggAX0GQ2lNGqYKQ6n/xiWG5FV16eQbXZjTIkBrh
KdnF06jJSTiUqFYuM+A9MnD9gMWJYbGREt8nT+yVDRZTNFBC1L1t1Wl6ck6XgIBl
1EScaqADwuDYC1qpU4KLNoIAgP4y65MHAM1ElDr5rPDLQXAH33VaxgsaWRxgN7o9
B3Gls3Ab9T2j2QrIU3FWAlR1SF09V++X+R6F/fce1kphFhpYAm3Q1bh5+GPSnMfh
zRqo7HGWhxHp8hK5iJI7ujpuMSu4O2hkhAiK1/3kTPv4y20TzONvJ/N9v/JBfmAn
2hUr8IRmdMLW9O86sPHYkLTzy+aQd49bHgFHLUu4+3hB/KPwLIja3wcn8Fu0Epra
eKEaVG9e3Kbjxe/CNUSGGXvJN25lkkCp0cfC5wUL4StL/M1cWr6x8Ze8FAJlABXm
5AQGdPskyaSjIYqzdGGNA+p6URMOe8OIng9EfbrUb+lT6o1oTHkAIN5uwon1jhGc
h3+EOfQvw2XlvfdqbtLQ58Y3g2sw0buDFSPbumvz4CecUiDY+cBWRlRxTpEIGfhx
SXqmQS9QloeEQyjmn0H47Wd2qMNcteTx7z6h+WqZgXjAf67IjH6Pmgk86RgnmDTQ
lBBt1K83ymyrf56WtKpUDIAX/gE1aDzdEInPLtq8CIPcIwOwM5QYCd4eeG2C6m3d
D+y8GVTIIaP6xGGL8r+gLkVGuEkoGf7nlWtBGadMMi6zoVC/SMkgswbHYnLHgHQ1
YGhbjST6aVQXDZbHZlni4uruJv9Sv1PHgN4qQh0jQmTIjmYffiMRhMsQRxoKzifJ
CTxgJT+aDOG6GYD/7vuS4BdmLgW1KWfQ+xfUOvTzm4QyU0zE3pFmeAbFP2gLClNM
LeRLhUicysOR2WngTeXC/B9zU3s0Z8uPB9TAwuCAGYdwblo4kzm0sHP1bt87TkDc
rii+OkbY3fbqYoNRLeaSePHSC0eE6oJDoQcgDt0GKR/qFmQeh3PoCx/ugQzZfwUU
z0PPShUf/Xi3RZNm8B+GQUJXaB/FhTh6qyoXlLOJLOXRTF/t3tU7azLAFzTVkP/j
dEqLlQT/QTz7TYJchGtRxfLmFlWLnwS5krX1Naq5Qev7owCmcsC+wmsWfCcvvZga
VgTOqR7Sm73wGP8BKAe5CZI7SI82VniommUDjaRqQRUuO8nx6RJ5uUdrVFH2ahON
NbCHqZTIGRcV1zA2nIFwmu4SZlkA7zdzlxpDtMrMa1KwRCcoHMzQgMjK8XHsZouC
qr4iix7p+UP8dHU+09/TFyqdbyeEVYq5YlEWYqwMALR0KX5ll0Icsgof/m3k8f5Y
qKhCHet6+pA+zcmYrup115snwNuKRMHIhvjtVQ3FMCGc8yRb8BcHfKNL2G7fEQbr
wJ4xfVEinn5QjzEif5R416wohrJCzVft5NB+AJ4NozBIO5sSUj/PMTYBPWndLQRg
YD1yFbpkISK+jLRYmfd1SPja3WLiAdUDpsdsc1GmhPVYcRu4fRYIE7bVM3izzB5+
j7H1tJYZ55WuVmDkiOrGqKGLYmUhYAPMQuHoKKyYr6Wsc6cGMtDSjIrRgqSyq//Z
kf37xPFGF4B3IxkwRea81YI5Ey2yCxsEITzE3s5S6Z839wyVyhd1QVUXdc8T0t3S
aAAvCDqlFAiEO/OpsgRRHAua937XpT/2SdB5LLp+1ABPy0P2L74KF5U6gu4hE8O7
emC7kF/beRoOp5FgdvXIZ8v/FfwYb+Osr/oI7AbTDjfoAgGSpauVE96Gesajk04A
uCZZcRrDgE9n3MOCKFgTJuKvgFuJ01t+KS9GgZMd1oNYdfi2v05epL+s7xtUv8F8
uKIn6oJUviGOgFEt814YxtnO7ez+3xBaK6ya6lJT2L8TJcsOAsdHy9cpIdGvrx9u
l0CAQgJESA7aZIue2H5uSgcEMMO9I8O7PJzsCQpAApoacHLunIywqvcBG6MD6u89
Q52k9XQxoysZdV1fbZD3POayHmqGmk3gMQHK+rr+M73caHoQE8lhQUBUiBdCDsjJ
E6rIfN/dfE2vk83vIO7zH9+Mk1z22T31t2P2YYgFUSnt5+3V7/+wDIjmSU1BM5ax
IEDnS7uM6Jxisy+ONjR+Hhg4wv32GnCNt/Nm1HBJ1WNuDMfis+PP87FXamnpTOiU
dt3aDDWD5aYIVworcKX8AGFtAUo0oSnh+g0nK5boKOvLmAKLZZRW4kRWnR/+snN7
34OTemAexhle7djAmvVMf5htLPDunc2TKq2hb4a/pU4lXZcus3nIIDc1OaEo5FYz
VjmndgG6EIKuOa0o8x2A/wZ6BLmyYoC+u90shAi6eM+4m2thYYJC8Je/ao0Vn0pJ
gi8RPMMNtLvJ078zWm4Ufv8WOzq0E5je6mDepsOtHWh57ZzhrlhJ/ne7eLKx6PiD
Kd5IcIo2YvKn71p+LQUfFDi1AyDexmywuYZJgXCiOUFQH2otfzEs3nuuU3TCwSG2
bp0MnaWK9+E2DRDFi1LaDw9bPGNdkKXi6x0t8hW9TWsvjx9LzL2b7jew5d9KAoNB
iXjw2AKlLXJ+uxI+s1KT+af00yWwu5WT2D1mMCyzYbovnSRdoia7K7dhZjmQKZP2
4JHr4Cdt/g+Mho3ya05WjeZd0HexQDif4kcBNhFUu2zOcfRYP9R9z/MqFSc9ZVod
MXcjsD/ynRKQCrWmBgHf8CWUj0OaWYIE4tIod6wSd01ohhMltIHqonQckkrxw6xf
C7X2OXUXmcHkCZrfOXtK82enEbI686ibzKfdAJr2Io8sCAQqhlAsCGRcDdRohDJa
yucr7qKpVwf1PHUtVsBPadcAmv1oZBSM7bLkMMyen0hS8ZK21LoCVRVw1sCqsx/r
J3vH3ilAHuq7C+azQ/RsURu8Lbt/9fdU0xQP6DrwJjdT34QjPXRGZbisnsMIr5WK
z2YAnI3l0YvZAwOmjkZ926gE0tM7QofQmdda074l5g1NqfflB9GEs7QVRAnXl8ZX
SIwCbiAQz2xO/DNnujuNdXbi0DfcUzCkv60SO6Oqw/FGoajaYf7YuUhS8W4r9JMp
ldlEqH8xm4fVHHyuwucN061kmat9rT7/KlkPjxK5GzF71cyypv/C2PMqMVSff3d5
wOLom+YOTkxD9wjnVP8mE7ME6ZH8kB2kT3uXgWE9GjSn6AFjAzmPa9Ie0drDCC94
QNVbMctmShNG3YOe76Eg8Hf+7HcoqmARPVf8Qb03T3QS3swWcnIC/fE+iPyuT1l+
BjSAAc5z6BTEYdLf5+VW29n31DEznpXsnH9hMKJuqVf5tmrsQ4pEIPYcdxwDGuo4
FhQpl68uKO4MFL3rpNxkgEb1w2plWrsT1B3ZVKPZIpTuWblNaFvWfNbrVCXQ8Eeu
V+NzYKPgGpAySf7H1erob59fZCklbLqwhm7VAg5VPyteRg5aZLLFrShqBriwTvQt
6QZjMO2hOpdhrfZxrpquqrXV9tFRwLsx5u1m5VPPxwo6xOqRtZF86WxFdvvVNihk
MmVb9Fg2W21mE4ZzuH04HX9Mc8fP8Ny1nEP/H1/coAK8a8hh2UmmJaoUUk05OjXU
UAPRpOZdFzxoV0aBr8tJrYSKxmo8DpwbyaWmVDv9+R8iemwW+swBmjPqbNNBWVg6
xq2AZ/cgi+CRJp1+cPiKmNLehQpce2qpij3C/TmKgOs2+gHzD8AXiEFCQdfmBU1h
2EA42C6Er+gRZTcA+4aYQJt9zD91Wa+xHT26851hoUcVgGCWjgVe5MaBE4N63b6V
PEXqQnRRVaOuAMmsXYK+4S0khqSdMBBKUG8qNCT6miKI2KvKBi7Q9oPtP/tacO3o
yGfhZldMTWrF5x4I9bi48NYa4wKcvskX1EyT5WCc4GRvZGfcDiEylqTULyKb9Qtg
AGrn0OqGkDHk7b5wgk8TnO3NzyGaDfydtbzs+hwqcAqwnxsgjk//Y9xtcrE1SkUO
gtXXB8TeMjWJdMuUtTOg6B6HU0d4mBC82hWSdIY7oloLQXfx8Lk+XwmQlhdNJP4T
92mytxpGPVuFFyX44npo+WQHKYTT0xnEM2BqgWo3RRxxjLIB+CDzPhlrudNPctt6
6sPoqqLri+9QAPAer5DwL4M1RnVfgid5QjxW9z4733UmDf1GWDpFkvbQd+Tfx5Be
Gq+6OJtVLBu5gAyUDmbY7e5mgx30M/9HiW6BblETFlnxI2n9eauhRUi2wyRvKTQt
GlZKzz6g+C2Vqn+oSCzEcE5BrWnh9G3t9noEq0WYTJbgvns92GW5szgVZsvWBHJq
dhSVdd6CbQ8YLLgwDacWfWSOYc/QbMbwrijQHVNjQX7hS31/jsU7tJuBhtXk/cXd
VlDQn+eUBGypDrGWe/fYxfX9mu+ul4/9foJHh+XGVLIhu6oAtJJNF0QBmdchVVde
LD5WrliSK2igtX7aKG04iLtjRhinEr+4u4D61h9vRMTf+TYz4NnpJTSiiafpAeHf
owtaAdvCAlR2RzNWHUn4uVuZnDwKrWfPL+I8GdeMJeTwRU00qAQeLmxMpUxkVImt
4PqtFnS/GiW6i5PuxisTyYwH0LrL2yZa4HpUsvmGI2Ch5RpcEOICpZEVNeUlUdl9
RLL7C0IocedbtXEpbyXfbTK8w29H7j830oBoOoF8gtp6Ynbubrip72/DdC+EGM/t
j851ydnXRNfpm9cBwcM7ax5hxFTuqmaolcJV/jVlc64TJOk9eNw8NEKdcjb8I+B2
ojRpZ+NxRQFKvcvgaE7ruUVExbubePvWwQfwqCzDKLZPOWrUKdO5x/fqmtvQR8Jj
aERjHW/n+7tVuFx+XQl5lfGA30WL3TqDgWig26YmLaY//GPzNjDJjUGXGWAMxa12
IJ2hbEDNkZZRiH064wMNmSapW55iFOm0P9mmv/R2MXIaBuh/wUM/NH/DEUwj9SDm
A0lW2IkuUgTTp5vQ3M8AXV73eQUp7Q5Ko/Oq7zSKNjrYHkBJvjJsA11pcSovjR32
cVOMMl3sgFaM05xjYBtXfpL6MOY3sQiUYxpOgcVtQU6Fgzl01iuq+lC++CW3oAcv
qbratOcqINQL8LDbY6hzUcEzxbisEpSzISypvCMxA//Csvs6Oi/iuoioX7wSjlw5
V32vwgpb2QDogEYZ0sA+AzAL6pghtYtxpbTZ2DXQ7y/oviDh6aBIR4oWggbMsXxY
eGvfKlVata8Vw62EEZLh+HpYHngIu5HynYtPSjHHGOsDQxO0wqlzl5hQGrInT+6b
U9R6zQh52okdS60oDkVw6EeCBVPxmGx5udrB8cW/r+JA11XvsiFNTOOso2nM3lzG
SP7jPs2flXiRxcftn7y2XUdGjsqRFVjKe5/ooKQZoKznbYV/tRuOFBEa+112f+xe
WX61VtQZfIYTjHN2VFjuWteIxM8TX+H2SgoYR/p9d3y6kLHPwHW/u62PqRs8WbP4
V1dgoX3vCbygkEYLUVdB76gfVjIdwuxO1nlnA107yMKNgjWn5aeCHamQbyCpB1wi
Kgtylqh8eIa769bLQoijl5H5ZqVNc2ukORR+4pFtKyG0apoGagXt5zir3qfK17q2
M0xWAEjdH0/hj3OTJwpiNj2WFKiDoeEGSMg8HRBdE3OPGzUFLd2QXypatPLl0XjM
SN467DPdv+vj0eFLyQRaPSynE8ApmFB0tGRc0owuLdgt5WxQgMSZqkGh55BGH9MX
1JoX6OzI2B403A+oDcaKWl5FPixx43I/SPllLgYxNtjHb+WSOFjHK9t2kqkeBQo8
Tzbujkjk1AKUj0QZHj8+KqQLtYnbDm2shD2OrWqRVN3yzRjuVBr6oKdi1N+xbJ2b
xajDXhfA2K1bOGUu1x4I8TpvX7wx9Ka1VSUIqBA99Qhq7N19FdrDxTb/V4kbsoaq
V4MZOKWPpn18x3hLVlXo+F51k1I7sxcUhcedn2jWxal8wypV484Ooqkc38pBfF3h
pkSxaTLbuizhK+wGCplLOm//dJ2iJdum42nDJyBgZATa9Lt49JTPFt3BRe4tuLmk
fUCQJljHhNy4t57N/8Ae7tAQg6myco/R02lA+FguCkXhjDlcyQUVt/Ow2qUTHTaH
hrO9A/yyfriuUYKRs4EmjnLh4zKzaZw3LTII6C7APO/EzjdvhahRnvqBlRlZkc54
WX/5UjJgNIzra5ZbgzJwd+QrULPQw0tce2McHnZRTYwWAM3OAdRUQqF/hlrptfBZ
wmBgFB8QwZNOmQRfsUIOvAZb56Lu2HTi4KG+C1LWM+vsBvMfT492Cm80Z/65dSJS
i9G6NhOLdLQkijfy/c/r/bnvHRkiZRX9OjpK4SLTjjNtNUhhaxHH0rgciuCZoEKl
8EdiBiKaPxv/gF+gRWHHsJUDmhCy8UJ9TyQx2y1stWYOIjkrtp5gsTZr9kUtRd4z
TMV0wRrYI0UEJYzgH+Oxxf3+9etL2lY42tve+96Z+ETrMzq7BeqH70fotGgkwxTh
AQXnCq4ZCqU+3zm2AHiXMh+5xR8Ru001JVnemCqHADdOOI9kPYC7QeMcqjaSlx+a
0rN/psEmtH3Gu3prXfguVjYmFMXm8orGgh1OpNNLiMRaDj9gkwTN9sfTwcMof/7J
q0kGlUDx22L5Go9ReabJf63uk+vAgczH90V0O6hGO14myzY9J7lo0afGtOkb6L+W
WPYx8pZrET1JSHIoYQ+nc3xbu5nOdrF0ajoccywJBWw5Hi9i+pBK4cGQ7NZJ4Kut
ZzfewB/n/PSFc2mO80IeRkSqrFClOSnMZNtxY/1fUkrzknc7zFZ/SrHYj+l4ewD+
f907VbzYZ8HDcgY2mCucsqoR7C4mYI7NSYDlT1n8WshHGloEukoMik/F5LehqDnn
ZX8h2SSaZ36WQgaBU8chxz7S3wx4RkAe1Sv0gNrpx6kiG92IopxLM0mFh7gk0PSg
XzE8M4PBgrxgMe/4E8ydqN7TcZvDfuBJrT0zNMhmCIKNo2BwJ7xXD9Z6qrNyJuNF
AntcZlR+xivPGDK0cglibEqsxXPOMHjxOAo9bcR54WyHm7GN/45M1ccLReUHVtZl
dzaIWjdiFPq4v59w6X7f6J0gQ5ydFpx9iMZlRnO4hDwhcARKXa76z+lwBzbT6J4l
due30G/L/TOSfvxXv6L+o+p1MtZMhn0JyS6HgK2l5NcXz18FxrMoZfQd0/2mNy1H
8SR978Zivro1t5jeuVcXPw3xTYlFugpUeh7bOl1wclEBi+s0/lqTVqjLFKaC38PK
V0DL6dZSfoKlVzhw6nIQpETGjZa4um4aawf3khzJ32DAeH0snPqbHCrJvK/r4RIC
meJynRjoYRXnTX8kQ+whQu4ZJkvCCSE8hmWKzQUCEOd3ubdG5n47ECM95FyLWu50
ykqlAQ1SC/n1ysER9QaiBcVqU1fve/d3fNEmgzEs9P8P9u7YE1NuYes9Vxry7wgw
Rv13KBlelZuWh3lIxN/Tg5QE1AOnaEdpjaHIDvcv8xWlt2JFgcsvHV43pyyOVecg
7cZf0/wzE5MW524o/zGsRGN/zzhG71cXJ/UzB1ox93Dn4NE0ltAkLuK7rRVvJ69E
q2ghbY7KWoo2RSqSojzti3k0yc7F0aSt6mt00VbD+1Mv+jOGLuncmMbLWp421+kq
wkzVgTLNs24tl3UNMvbOFeEhDpftjxyXBkX4FvFTxPUl+RX0KTESLXBspqpnH/l0
4xAs3hS+ous+JzO91MypX3zHRt9ODvG1wy5g3QF/6veMXiVmouAEMWRmeDqvgXUs
E47sukhFX3EBSE+4PgYH78rMTo61tYKLkBPaUXdnlUeSo18ZhpX2qs0WXfzox4A2
Oc5sQeq3XUUkjxRaHYTEdo3oeX9Y1GhaMEvtJiz/RDb6Qexp6JHUn+n34k7geHlQ
4vGMpOvdMLayJsqNkDUAYloJBwIHrVbCa5t5R0gnjCJglMjmpgDM2y3j/r8Jy2F8
gDwOwBAF25FCbd/Aifd/M0alyPXjPLjkeYg7OUWtB6dc6fJlIGJO6VDyaCc/YprU
TE3YEg6h6Uf7wO3DFMUoshzzXKo85ilqAptOQxu1sy0x7b3JkDkKC9mjvgdq8+Fm
YTlIC717WOz+ErNXrtiu4nWXr7+oMRiBMNhh4C7Ln61MP6GjtFQ85IRm/ozt6SW1
4Y9ifozBVd69raD5QWPZfEu6tRRWsxDu5SYLVLwYApNj3cJFjyYT3otQuLIr17h7
weqOakwwWAem89RaMqKfmy8r0cNjKRaq47XDsR2tXdfmgTQIkYbxTG0mFeC1jZu8
9irrsIjjORbeGCv7sGC0tLWiGQzHZNWPvGBRX8QJVTIHCBi6+hw3HslgLJaMmlKd
ULGk74qyZe9/18jV3tw18AT6vP4ZuzVvY02iY0JSrLjVpBMvLV/wsozO0KnwhyDT
N941PB1SFudSKBHSopUzPQ5X1oAa4hW1VjuS3Mp8az1rlcnuUbSi2iXzJoMUQW/r
txfyf+xwxRoB4EcCuWfeU9RXMtihAuj197bRhDrOZ01Rfufof09eBQ6njqMMrleK
xnjXzrN3NPBSimpC6UKpLlErNN5XxCTb8OjgTJb/gjbyZSvrJoDbCX5ji2od5utm

//pragma protect end_data_block
//pragma protect digest_block
4eW7y8e4/FZiDJ+Q8+90dsIxmyM=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
uR/xMDKq0/B2EZupw0EGBJ+Wd5PzjHo8A+3m3qL97pzWesko6EHk9v2Rrj+3q9ZM
5+RjUyFTSUnLsh3ckJyb1jnb+zM2AyIrJJhQblLxljml/x2ns+9AYWO/NWhYIjOI
sN+ULinrbanV7+zDIK1EHZcw3ZJgMnwXrDm3GKbsppl0fx1zx8BlGQ==
//pragma protect end_key_block
//pragma protect digest_block
jkFFkLG2AujXdcc0himuDnGR17E=
//pragma protect end_digest_block
//pragma protect data_block
5AmODNa16JqCBhNnc2TuKSFE/PUx7Tg5zbmC//M7pm0Fwgq2lDLbJrfl0R7Z6RwY
zoNbd4Qi8y0IFiEc+5baxmvFN/JxTEbQmDMoDokRbrhXBCTXHbrLZKckNgEXIO2c
zj9LOVLvNHpWeHwigL64dr7Y3RgPbPkXPJ2ytGmuk35sn3anckXquH5bvNjOuHAp
Zd/94OJFsGhl7ennKtsektPQr0AKehid2TsbUkcGCbXoiF+IdyKZWLk69BRpjbbG
f9APKZGpbBYSF78G0EVDLO3AyCf3zmI/iQd8ubH3FFFVXxRBJMJdwxmh8X32uafI
R5SOKM1vZdjNK2JJ/eZPbXMwA9zrjAZyFPypJ+YlFHH15v50S9nMGLcw4MWeLOu5
8ijb9EV9hf5azz8tC4/D/JcUU28ugOXFMkPdYL/uiqpuPy+Rq6zqSbEU+gg50l/K
F3CpNgYZQYMNl7JCpmwhcQMaMogAvYtRuoqKavTCZRV7qXHUKmTCaMc5I4uthJ8D
ffH0j3W7eoKSpPIsaA+uqZiXfzNCyobL34sfdwYpr7uD5M2vkjd8NKMO5rx51IRv
vz70oEu2y5/U0i+Ff9c4N9B997KxOlDP41h3KSGDgVeJicwyVQXa9YHx8uK8qBF9
Movr8zfhYtdPbGpsWFgCY0GUlkbO4nJ2pwXDrRgJWsrp1dITbTV6QcVyIXIFkkYJ
RDu6crRRRG2z4Hn28ml1882gCw6s9HSKCh5mz7IOCtSggFBDg5tWhFMnGSeSDDI9
MYf1MxwEcgQYuX/+tcaNHAMx65a8QJxqKGIkUzZYYLPFkFkJFF8TS0mGdTcpzKSL
pvSZfqV/OpKaWbd7znl3v/kNFGAsJR5tQFy0dDkX2JpPVYX9cZKPPgvSsbgeqaHt
v9uR2IfNwlrHRYfhKu/csiYg4g70MQdFwO+4HL5Yhhmxl68Rt54P3axp3716X1KR
zhKGeRXy2bCe7ow0RUZu5KS8n7xmFwlnPQZQBcHfmC4=
//pragma protect end_data_block
//pragma protect digest_block
SZJEqjYxfTaI4itHDSfCyC73+z4=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_vip_protect      
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
xmrMgATrg33xm59rqqDwrMSwnJwbFACu3mpMYbN407+mAEivyaphzesdQx20I1Ws
tRnaJYuWjvcCiRkrbjYjI5tZhl49PIOAUYGlRbLf3e9Z8pk6NpNyT8d2f26J38s5
xNbrLplNhDTyYyj00R2LHz90bpgS0OukUp0rLv/hovnH7yu41XoLEQ==
//pragma protect end_key_block
//pragma protect digest_block
qOehCy2f63XpIW9Zhfnse0DPXpw=
//pragma protect end_digest_block
//pragma protect data_block
ziNpIG19ZTo/Qf1UHjVpRmOMFuCJXq/CyKWlL4taDt8RP8LmwFfeA3THYK8yql5F
MIBj2g6mE1uatSZr3DK6eaig3HlhhJGCrp1HjYRhZVXuKZOpEbnAiOqfLdX420R9
CB4ZIzinCUzTIVu7paAQkUgQbT5lGeS/A44T5Qi9qHjD+gwgIqTjFR6thz+TrAo7
0iVKyVNRClURWOG5HrCeEzsLp9Pe4+4X7vUX4LiG/SIHaE6XNquBOr6jwxXL7ptR
4GwmfXQ7x5IXe3Tw6RvNMJvg2mXqtE5fz0HNHMKZb1gz+j4pW74ZFk/tBlPoJcUh
3jT8/idq4fWWypc1va+45yJtLOrhgZqu+hbrSU26KtleHzTwWhaHkmNL6rHObe3i
IwAVi3NNtFyKRosXAM8tpEbKWnue9dkA50cDYPpIp2E7W6PPsNafGK7k3aEv936y
mFxA4WZUleFWM/XQ37UbFmG4YTmFgbCmDU0SnSEneOdDu3N8H1BTJ/yVBxSHY8Td
wMZInWyNYioznf9UWr+6H4KEhm8CQ/e8NZNrj0LPmcI4PplTxjZErw/862PrcSzt
g7eh8sLYjDOfM2khHO1JIqrXtvOH5zfdEWXGROiDe9zJEFHGgaTEZD8nL+ELY+VK
EuG8bUkjxog9X5HDUx3GdLjqE1V2YZawkAHWTt3kKGJyIicWNsu5jKuSN6EVVn9B
E0Ucz7Xynt3Bpi+DK0gvRSglwvnbavm2gFnVMsHnZ2FiGImQlApXR6QqT2t9R/4y
trln4+KD1c1QRkDFxd1G+4Qj+2b5mr0+Jg4CgNGRDKPJWcPobxpQd0kgDHW+q5Xr
IplXfhTyf37l1cgWSMEvD24z3ah20YMHy/l9NvwybOg0NifZ8NsJ2zjifF/0VJ2k
iiyBK0YXI8uyaKtJX3wGUR+pbX7j7UaybPrVQb1mC4e0Ie5zPKy4MWbiDfr7c94+
HRt0/a35zmoRQlA23vVhztY7ibyufj99x8GSGFEfxWv5/ClodAjHmN/NVqcZPZ+6
Q4yWLezqWyXTzYg6Z5Pz0SyfP7eFO0R6czrvWMPWE63QYNHPQnz9z46cKuBVw7B5
773lsuP+SOuNpUuUEjxwsm0uY7tPoWDsOt1sd0I8GIbpPtfLkwGn8afsXN6/rZfu
0MjyRIGn4URLzNZU8sHfj0b1SqZM3ggK+uLxqGm1b8+5W+FZ1xZDiCgy0CBezB7U
A7Kw+ugZzLOApkwMWOU6C2TikwSTQZLwl9Veilo2QYGTsOIgS7bnx9RkBWrCJti7
lmMaPDwK7TtC2snb74ZhxI440NkAbohmaby+Y5v9II8X8avQ046Epsgq4TU0VuFn
CnMuKR/0+59S1Dr4JqCSrTBO129+Nj5BHSEqN0XcG0MQhV8WfT0HWFh1FW+OEk7N
wGk7kL2zY5PZT1uUgmy/tqS5MwXFG8hatPctvztEi+IcTXxily0Tjik2J1RkXQ8A
Bz8ytP7vB+bddEi9wh4B79xxPCAdge/+kx/5w3/Z1Gicu+58nX7yFWbUQcUCMuHX
oQodkK30GUhmV53faK9ngKlO9Y5RAYGmZMHvF2lUn+EuNIoW+mrOR7jk/bBC3pRe
bqe3sso5mQEkPHadAh61s/iUfkhB3zeeXpBMGEVGPIBvKAyvcktizcxysb8hMd8Y
kIq/FbxToSV93QMKcF9MfJMJjNaUxjbOJ/EsbsgsAGEwUmsNDifd156VWpzhASfP
Z0D6ETzw3XfK+y+uzHmcoVrgChHEWd1yRxBJpdsf5mwS70lWFV/4FsqmsLPhZAGQ
RcAl75LgIIYMZ0v+ioITjka0Uyxy9JY5yQ9x76XYInpoKSKOWVQmTbRKvWy5WFfu
uIB4sEtCUVmC1Rfq5ARULrKV6dPRloj416VrC+AuoGBYNRgsjWttxWOxl6jFYFc0
e6br1QAvkuXsLLWmcRD2ZSg0lvf30VQfyVO43bIC41A56FbMkQI13cYvxEm0vLv3
+/67Gj5aPfxOYj6ByWk8mGHsssjXZPfUYaF8TBaBM1Vkr6rwSWb0QmcU8Ua4TSRb
35hUECYEOpFfqGgunWSob9E/C0+vyZOo97p+nu5hze9nuaqgfFfjMCGhRzhmtfMa
yBu1XGkIiTAmaOd/PRsYVqG7cgGBSUGG48TjoV4QSoQzG3QJLuSkXJKgO9ADssMo
duMVC2J7m4cTG+yTQYO1BVqyKdmHQ7FTltVUfDftzXzk+AG56FVtpXz7qlFGJpVm
/zDgBEMQ7j119DtQezFJEec+T5aNFBCt4qTTlTdSdbKnpVtG/pX/xrd2vfbGexiF
nasZlwrftrZDchaXoG7HAAzaBZvyRtfP/29qCIqjo2G1be9gU9QqNAAQTyu6F8JA
jYtMWC8Zri1gDvXR3GCv4l2fXp0gbobUGJ/CtFtn44Y23MwEtkz7g69YIAxc3mZC
O2aJbqPegBxwxmj0BXDrc7bgDQ1ndQwvxWMH1ed62K3dmYFLqaTjXEqTZ0L1AX+U
kXyx/YD8Ncq3sYdKt+CAo1Q1WbrTj0b40j7vziwwT3abfly9mor7PNHy2U8dY0ME
ubVHKvn7kZ+I/KTctneGXHQSgyYcAQQRfn/Z617kAddU2BWtqcCc5aO0Cw7y/riO
OCcq+V7Bwg/AcK6qp1MXPtpcwb4cluHdVdu1srYbTS2OTVd/pD0TqF7SvXJ1lt43
OOgDNkz81nZfKhn02JE4eVOsrWIjoUrHCDozYfaQy5ZOhTYpO0OUULAP2pJNxpCv
iiM+w1nTew3g3Spd5X2OBcrTXOXq8Qf5ogMfSplAmL707Wuv0cqhN+Hnxz6KY0t+
ld3PUcsYjrpVhganhCuksNbpjxBoE2wja3zS7hGDDDa/5pz8NsL2G0JAXlQARQob
Os6KDHab9Vi0KEM/wWaacSYOQyIEBbem0E23p+ulKobLz0fMsTIkTZHfMjLnwZxt
NVGknO6cQyAEm1wLjT12q2evocrDVzQVwvNN42SLgerhT+RELla9NHMpZZSU9Bqb
1jC3VEMMH5V+XzN0ZZPhb+FCvH7SlQfKDVssAp0p6ETzUNChREKBC6EFjlf0nAVk
sRl8kw9mEHmnwIK8mQ2KHPdDlzMo2qpWppLrVTXqcFvghE6cmNWfUv+kMLSSfHxC
c2EEWEgnqgnGe+7PYkmLFbR5fkrz8XnSPltg4kwMZm63Kn9f0s/MhpkhW1Jd1BeC
8gS3jyKXUpXxqkaki4XR8oY/uP3pu1ZTvprBv55yG81SqJ9pAqsCeSooQc8zS+IH
XYHwi1XtUCG/IP89CHTfZQ/6u7l+HnXS7X5ILUB1TfGsI9/9PDYxBIxs1XrYF7R0
Qp1IGH0us1zDR1sM25evEPvnwPEJD0BtJAIZCbWnEitm9Qtr0CTnP6odjHTratlZ
Eycqe6S8SmHNdsotGmjohdVOI8Q9IX1l47agQost2egtj9uR+sa8JywBMFZ+/btr
BqYIcVN2CkEx1et1yNw8VQ420PVelRbYI6E72OhjVWWk5UVoAc4sZBpjHucCGcRk
AhyTftXcPowm6GreFqMZ70EE36i0hX6OottYmepdPmpfb7+7NzjJeZGZ/P2iE77o
vqnWGgX4xlvVN9MJJLI81gKdkUuSNfIFU3ppbgqNr1SUjkIIyCqiIrqMoPuaKrN9
uraEuK+siNub7LOiYt1sS0nVgSl7/fQ8uAd1MnwNR0DIaWEoWWojqwzxE9lni7rS
qTuOJRCCCIMEubfLSpAHE2o4UR8xczIZx9YIu/e29OL5JIJ/8qpxta/+ssf2F27n
UYbnaDiBwcpoH4cnOTFEv2FSK1phjzJ7ZWn3ZDY7RIq6YYARMb4AmAfzlmm0e6UJ
zQ4p6kEyNr7n9toRYuJorwZb1k18IPaS6Vmi0fXNwbTe/rw2Ec02sZOh1j2wRigP
ovOEtPgtfmQlSxGAvm9R6RKlUrHWEu4+a1KD8WzAOfoHYw9ya2Ej5nTXYlA0XAun
9vfTazG+yCYagHAf+b69JenvwWmMgo4kfrumO3X8EKDwojnDrniWm+aWHEBGCMSi
gdHrr7W1QcPnJ/qcucEEgwsjfuUkbj859zaqMwAwFcRYdF9507AZ05onwAcR+5D9
AKHV3Dr/7BsUl0YeVDz42osFti1/CSCcClaFpgcT7C3nfdhicV5ynPRExco//W8q
fnx2FLv4Zo6JhrOXcyIdmTd2AUAQm1QN5WlOUNt8wIgbeeQumc3QrpJX5IWPifSA
uticopFgRPb61GHQotG2SNKlrOXrOZaFPNn/9kKtskQIOzdiBw+LrQQ/YBhcfqek
Kja34GXx4VZ4xj4pvWG4196QfkRJoI4Sz2DRFdQSviqVl8xRqkD4H/L3ufmVe+2N
Gb1i6HEoTfqg+zzhu+tOxbhN1kvKwV9y5zfK61p37RVcePDBFpOFMGcIkdsJniOB
GkkYrEgYpYGdGZC9dZQ9yfp2zqsnFxbNPVeZtS3rwKcgXz7vVhLY69NIO36n5Y1G
wTB65vb1FGGwGD9KuJ3I0MO6saIYuFFsqf2CiDsHTSBx1QWiDqxK4HVxrHEBHljQ
VFkYvNYTUdp5mOiQh7cdHk8TazmlVpBvNmKHHXjESLWyXmsVdQujXKAmMJdGzcsg
CGg0lyZHk1ppoK1n4Cfr5N1+8zIga9oaw4X7xfH9Eti+mH5rpy0+o30qWrc+BPOE
a0cAfOpf0ZY0V14vjPVFdkQ28cQ6FSftMfcvManCTuMQ1yvcDk6QI6sqQ89SRHHK
ZSY2KaR7G/2p51mvzu42zisydiIWkzgsqetTHUYCM7HgYjEWyxHN+FoMB224ookX
PDWM+yiDVIcX02N94kVG+v5lcwJvzRS6SREZWsfucrpVJuyaI6rPbniiA6KhmHvQ
hTwL1KwU3dlU9gE6NuvVrSTbjpZ4Mpr6UMZW0jRbBWhJdyqpSgp4vrJIZ53NDh/S
Eq5H+Lw54h42Lw1vUtl5jvmr88ambOAn+mH7/lyLSgTKwMLtOSMokF5UrVGLF1Pz
daVTDysM+NLTOb6QjL7jFfM4OT6tZHcZtvU9eiDl1SnVf5SFY0a92LTOxc0ZKiPo
L2hm7OezA5TYZq9NGowo1COmLgdtRZWvgPvNiAwb4UUdk0MWuKclXcNb1odLFtLz
dezxixUgzJMKHcOp1P33/4YX5OET3ix7/iyCj56d/WuPxbsxriai5Ah57rwUq0xU
r/psiyD3acJv9GVDsmZ0tefcKep9RD1b2fpu17+kO7WK9ApGrDrryXpBqJFRxdri
qg4AW8mf91q4p1F0NcfuQ6ljnCmxcu+W263P+YJXmWVGXYQ7RSk4II9BKX7cY8hV
LMV0yIMPF7/vl7cV+mzfQ2NtKUIO0p/04b8rnCI/HbMkSECCim8cqP/NtLEmej4H
u7KiFUdTpPxIEWr5v1oCYtrSefP/vj8H9O1vsrx+OROyxrBSJ4+Poj3lfg0uqBjy
/av/WiFOOPonpoEokysbGeXWwyxk5if3EiO9uCcvrflB7uQfkU74WRVZUgpC10CW
RwtK0+JLXX574s6kuocWhQ9bBTYEmDtgjqZW04Rpk93tPoP+XVVD+P6Z7Z8kL4+8
WXQRiSo44TastIHSJBK2i/5sDXJ1aeY9g/0yIKZO5ZFH4PnTbHRJssjTgo841kBu
2931Ci5i9IcbpYSST8Uq5oYcLOgImxsYH08TK4UlYizpAwUpJ2Oj7w7wtppyktZ3
JSL1Hf8DPqVciEeHJ9R1RCiZmf4Pe9UPwuAvjdr4jcWMeQxs8OxtnAOuuvqOK/e/
aGD7F9JYxJS8Ooe+0J8KRvNiDfxeROWXvj0eKYet1kNGri5hswzpMaYPxjg1GGxj
CogCNPPdrqlQVUVQRg18bc53uDA7sem4oCIw9oCCuXIvpJj2calml5u9dpr5bvdd
SGKp1HlhuTxQAzR3t5/Nd6u+qafdauaM4arS9r5ijRagqMLp3aGjxfhcsIuQFqtO
tApaiFmp4Ig+DQjaYnGBtPIMpOG0XQGUVcmGaGN6/Yu2xboNV2V+kz4WBtHIpevQ
gUaYtOgPb/RpwqRmuk6JKCnYImXIjI9hDWdJ8fXARAyXdVeUaE+y5RRhaE7MNWnN
h1fF9HZZ+CxQFlH0Urxdwzez22SiucaeF0FmfDvaoNnJ6DMKHG2O315c++hnRuCh
cC04ox/RgZRa/3rhsLU8+aAqQuh+z0hstXeDkh28SwXNbsk1oHZo13PKylvooOeW
DMWOkw2/LtTKA3GHtcIDe9yX3xIb1SJ1iAp0ogi0mAaM+YJDjLtgEAU3bmNlNaJc
JgQpr5b3QEqsUYZvDpRyI8gzrlIZdCzkpqDoREnpFMrPO4DspMTlV1mNcQFO5YVZ
FDRxDUgYwFrhc136izh1c72Md7s9cB9wvHhvMQt18DbUNHjITtvbxMhfk1lsp/m/
ahUqmcdIVVD0mL4Hvwbj32PnJdRXyYhndhZgN/ckoX9/X+fezLZk7d2g3ENhBZQ6
B+KgqldxMFyDI1ubz7XdMWRNsfjEfGVRZxjlr/7BhLUdgt/kXhMtXWfXEt9vJUKE
bBO+PAWL5vz8Mva5fYyTaupZobANHKO1xnhjwPeja6FNngD8eqFtBNc+PxdM6Ik5
h1POTWs85usBo5xzeunxe/FT0S2KzBBUJFTMS68mkt+shRe3D8CHNi0d2ssVsWmh
dlAjv5/MPd7YSuDe/5JJQE/hDuaVZjZio7DxoddHLIL81MvfPzq3dXhBhvQV7eqf
j/Fw7ZY89rgmJAQLhk8jgY+A2LqzmEukD3LyhIttxFNWoxJ+ZzYOMLq+4Q5LA0gf
z8YjF+/LZoTAxu0hlzJB0JgQk3iIkyK5A3xXrdmMjGE2UCOIuft6tAClNaoEMxVC
Bof03EUiVFxCFnAXPpM6OhVR9roMcoFr0o7C4ta++YpjwxwoA+cOMbW5Lzo5W5R8
yBRUNR/bwQ8sk806yE2cK74bBfX2x+JiPvf5fFVRflA4jNsA672eUqK33hFrGwug
y5Qn8qAxvEXm/fxbqrbw+QGbQvdYSi8f8wnh8HM7zGnqKLL389Y9oAoW+b4sI+SR
x/vbZjuBJMrhi3d7ZfiExL3ycYbENK0Hcl1TEYeVGvBDf5ZB/PUvROyPbsqX2FkK
aFRy5F2gujIKoZdD6w45OVcaa4z5TXmjtbHKw1hmarnXqwHR4rWKSI84ec7TQmsn
PZxtVdw00RyXi1kgsutqKcC0H6ipMxLLWuxKawmaX7mh7wvWgF5nW1Jl3Pq5UzFu
vRS8ofYAdY5Dkb8AxfCmAmR8hxURu6SVLAQHV7JTOfOcJndKVJ/t58mrF/BRIw5H
WTdFoSAigzzP2KMLSahudE1qxIezPdH504o+cpqNKm/f2l1cm2inv5QH6Jx8bo/j
0z0+1vtnQhB2C9xBq9MI/gyOpzBBy+lifuvfJ/HTd6u4l8zQbyFVO6ycDxG7fsyf
x9EFBvIRcA3/6MZB0Zj70XTAOhzn5ua7dm9ShKn8qQvM07nA89c4hJYKi4EsApAs
z+Ku69bNSA2My7NlxKZ49lymlQEkaFI/ys1yZZKTF4xVlFvp7B2tiU3EQpL3C4gy
ZOPG0qdSVX3o7kLPTvSTx6Tm7FN33aFp/9a7mpa44DyE/0SquuASoCKVGWCB3eXM
EiRZbOrV+KxvU9pTSFhJafCon6I4uGVAw9v4zL5/lVkU+KI6JcRBtTy8wi7i5P8K
2m2rryHXZacYqc9DG70BktNrEJixPot269+ar68ypmuTS68gQtFelqvkukQ1g6u5
dlbpFlYwwjGHovpAxBuHxmQ+MIiu787HomAPuXZ5S0g6LnwzlNHlDr0s9Qn/M6tt
7wUgfKHilUyL49ehtuGbTPqJq0Ri8mq5/7wZyDZ2uwTFE/h6OPGN3fbFO4r0jYgY
Qy4X+LBKygaU8tdaEq+JN00ohci5Gpuq/H7FJaQQ4e4HE8Zwy6BIGZ2EmrSKTFhF
WEutqkmJ31ZbOUUhvySWBcuvFI8IOOkT3tzt8e/q3OjbAgzfr7NkuuXWwg29O9ta
iJOSNGKYrqSGdjbk1gD/V69WLk19eBIBEAw88HVrnDeAUwKekEU0NJaZX/7wpSs1
TcVyLLvChxA2361fWGtlscXMb53f+Ii0gI3YEsycxFpaPwlm2auYHCb62zaJuncD
iGaMJz2iNcQMS/mSq1Uiz9unzv2QOi2fuJT7VQWGcc+T0l3IyKFucgSvEo53cit/
dGij9sNd+I54w817d/Ba6XuT4Wxl/AmvQ/NxOUwsX5RrKkkdlL9GeZcVpfC9gaNi
pXCx1vVQfnsEa81Tu6Yyzx5zk2LERmBBhAcboC8F4iNGqw2PIS07GmpcTYDj/mWb
4jq9uwLNkyOsMSRQqiALCJxtFgD59/n9YQ4ECCQ7Hooiqc0EmNr2BJC27kvst6Wn
KWwgynnugq7iKjvxr6kxtVhgSb6QIPRdSUVCvZ8hrBUNUFQqKJSX3JW7p/AmudEV
qDZrc2A/ufMQu8OTUJvngi/VF8KWOtenxpcs36hTUhkCY2/O8ajryKI0IJBNlvA8
9QgBJzVXY89RCSb+7YQW2ncdIPLK5nnVKe9/x5x00+yhLKqDQIcmBeKCzkdqW+sP
fmaB/leNmK9mFYJ6NeH2kO6JZFAGs0yagZXdtKlWiLXKyMR+zOfNkB0ULak5rKbD
IslV2CnFF4QTy65LAN8f0Cf63FCaUmYt0mMk1urEd8zO765f+2/C92hhr8Ju1U5i
iigvDk1FCjBWVV+0kkGOvD3kOy7ZqefR7JrKYfLvorfbQDDp6Tb8KvdcRsPQjx9A
okJWDxAzu2YQRPceAAnN1e22BfVeZ1pga/kTiEdDfr0aM4wMGKobm+EY+FPA+HdE
VLZ+0lXT8WQthK46AAt7Tx2Vbz9HpeoZHVqIg2YF1Tq5FZ/mIUxdo9MTE1JSj2Od
qp8hp7Y8YO5vXNHQ3AE5mSlbYxIiBiZiqQIauaXe0MxE71TYPNs3j7Ge3tA0VfCt
iZWz8RzZLhuv711Pyd51oQjegYHKuUHbEVzVl3xSvA2s75btaDGOHdgUAuOY+SnV
98wuJZPefYJ5xjT5wMzUEzO0FmWuvIoNJePlYmsbKq69dt8uKXX0e5GZtyYN+3IO
JF0LN8gjTtv8KW0zk54yEcNVigh/aEq9kiuoiQcue68QqU9ZX7EC0dS0/YI7CVwy
KG1D2H612ngW5m1mMYlffJadFPRewt/aylazcIT26suAh/vA0Sd/IDBOPX+oFvi9
iO4YWS1reH1lnHCxdS7SHqM4LuZDCvpkk6yke0H6qBiFw2Ti3mwsbV06n+lbK8qc
IzmwJbBb46p0ZQ4xUjQti30N8SWQifHdsjzmIQJYjfOPkn2OMwbgb6RmuAVvXXa7
NYDtCEKLCHjcbILMT7Z7Wx+q6sK79FSCoY+aDZul2lusslTN6eckhm960VZjvkXZ
0EY73FDU4U98IF+sesN2+LYtdRdxvstU3c4dW6KuA6bX9nz+tM/asVckyfuvBHUS
nt9anGQW9l/VgzQZdqRw2Wv6iXIWQQSrg7lUqpePaguXjMtDZ/3zU+rGHjTDY5SR
sz3ztwP5g0UDtNyBfAqcv07FkOFaTo2C0Tr9MlZv1VADm4rdPZIfAX1K5y60VIH/
dvZ0yq0bP+m2J+57BivXl14Ckuvt8hx4OgZr5jOn3t/8/GuyVj0X4X7gDJvnwyle
qrjR/pK4HtaSs6ZG/2aVt90M67gEIWtArUA4u0xo+zwk6HhqmEGSGXwEST/2+4MD
oqqGjqlPcskESJ75VdmkvxU3yF0kNLnZRKZw4b/7kh4wK74Nc+pSD4lmGNSQXnLy
LV0t85XbPsSLlYI0ImPcA9ZAlPmuUuGVRupn7FHuoXejMzDUsput9CcrG8S3KExB
VjI9NKPnECyRhUyQi6MSNtiRa0hJA/ByD+RbywJMaS4Us38/8Lm20yY02SUGlm6H
t/935QgPJ1p+pON3sNDtRHvVVjBT5eRhihJarPnsS8zr+fOb6PVCzvT8pgQmomAU
zFNK2FqiIgvI7VwIOrIV9NgUThhaPkp+PMBO9UDCV6UHoNx/rTOVOZasOr82O5XT
gbivKzIHNvXlkh+6Cxn0LJy3uhx7pzHBTpeLPObQQ85b4sW0nSi4ZrG4TbkzH56i
vHyKqQD2tSFdjw7cpKqB79ItiQ8FdCHTmCuiTCfbTYaMjcKUZglT6RLc3o9BmEiQ
QVo5pMV9jNZEcXATyj29amhlQZ73W9W98KmGSauOnXpNmUtjxNlzWZTzpDwkX5/1
VRBzgvBGT27k4nImaPosPruO7HCyVdrCosaceRFOcnqoAW3WlaQJbS1MG7JmDXPk
IaSMNaybfL/G6DIj1tH6IyACRL/Bmc4E9NkKl/BV69Uz5AKLXjE/s910CHL/MF5C
D39R3yWMCAuztbqgvN+0l8FSGt8CjF4eXLfLamJViwQA3mFS5DUaR3Xr4ZbaL++2
xEkAvSMbYfC5eO55muusFqIk5/NGuxAVJnWq8qU4fSuPIPMtpKfS/x+Vrrner1G8
izb2HALitS9JNGE+hh5efhjm3gbPkkp1HC1+fWEFbYmrbN+4WwGpqMtWJj9ftTjq
Lu1agrxRVDZohGx7lfgCBxIONAwz8VXjSj+xQJh7RBrPNsYK/J9DC8GLUh2cHBsS
6BwOg6kh7bC3A1zMDKIhqutrl3tG52dmSzrcXnC79D3YuHwgRujBcwgCBAPUHFlo
6IUsS07h8KtVDgpxWiZUhgYrFnydQ0jpEZRnlsnPnrVHJuMW0ZjYfvz01svqk0mz
+joKyrqqaYKVcq42aYVhcUQIMPyiOpSES+4wFKziFzmsrJngS9OHAsePtM+uK9QU
CKyH4bfbt5Wp6+y0PU9Ye8MeHwqfjhXsxoQNb95kB3NWLAZo3DTktQArc+qdppcT
gQBHGun+ni181SKJojvFF1U9guILTXoxqb0CN2qkmdJ6I1wu3CoodeJK0a/V3rx3
AV/T0r1FH44ozbN1A0AEOK3DDUCgvTL0AlyydKlK7WCIc/gJ1kaeSISnJIv/QOPv
GrCB9eXL223I67PlpvvrLvaUbVjUC5U22Iz8RVd9spv+yzaY2gJTBiwHTj86r+Pu
MlfXXnelc/c+GRxkd8+SIEpOAA8h4b8nJdM4O9wY3pV5oEduhJlnFng5LuM64B14
jHgFasTLbVZXN/yo2I86yetLE134bJ06O7PNKvslxwnz23Qvc1219JN4bXK+HqzP
FdB2efmLZy7UBq1xnmE7f9I8jpVJ/uZ8RWl3XvGPR4nEvTWSQAzMab6bzUSVdLhF
WvUItd7YwdQfdQM45XsLcRvvWX7WecOHYGLMUljUkcI9+s3nU/AJ6ZDgFx/43Bxg
ZYepNzpMOfCSihqYocWcdQom9d5IhhlA7JxAYjTNKQ0zPqZehCVT8knGdipAMgVc
udyBbjkFC/wiHN/qJp39cYPhzZFrX3aV1hiTxUz77HxYuYFkeg+FiQXP3wgbYACd
gTpX8bOLdR9xSGKunSd2Qe6AcqXC/b3efDdE3kPD9QyoTeDiwk2Wr9OcjM3MjI5j
Ui+j8QTv4oANbzBGqnYg4H5D7ZW2XrYOqdddItI0WLmccIlEBeWK7LgScy+MSZWI
6Pj0ozgsNbeWpA1gurfBwmw1MMdGbIpfhcXeW5Go3X72Zw5yfGbMB41PMwG+hT73
vqza3ExwoBB7SX8voK+MHxLE1dTfpO3Jp9nae63YLQGn3l2EVhcv8hF85PZBUcwk
EQXye0/ZhRKc4oJpkx+TSkb/x3L3x+Bec+aFwA8daOAi8cZq2iQZoyWyDSdMe2uw
oNwWo+6amqd+r56mhCyX6S3nz/hf3LCaxE/88yok4yGka3J+JznKmzp/LOmJNPvn
h5opy9CHNwe0iJ8vHBawcc7DCuQ/OjffWI9BxKG1FTY7k40fmyM+cZa5mDSr8zvz
pwr272nWrFPTmqyPoD2s6Msvo/0XsstDYuowX6wzy6dA3auxJc80SRl9mjb8J0Ay
2BtkpNt8CCTPjy3SDstVrt5v5UXfVRcT0rCJJBf1nbt57qNLh6ezJnZlF6DGELtA
1aKsmAH1CTFAl5d6HPuOjDPIag8LfgxkkkNBnhr24OQDayH63E6Ku971cAHvXugQ
Hn4a7Ra9HSgJr3p6uUnzwMCWTTOkqzUqhnZbJOudXX+VNnw6vf75KavJvt5a4V2I
ekRE7jwAWJ/lJo2XQjU6gkk5XtdhkqqRMGIYj1yHfYiRIew4g/lxe7M8/37bsuBp
UiGrB2z7iZEx5CeaMtSiy15d/vr0lKBDdkW0R/iAgRd/IhMQTtIcbCr3lXyZ7xHy
Rday3B3JJOpvB0BSrwn4d7RkBBlFWgi/jYEWp7KH6g0EL4vMM1Vwr/09lx6yW5j0
izT1rcMiVKAMD07vu0rPDq/BaGWZOSrrRpQMLCapo2bsdGGSjXLRE9ECenLywbq1
DkaBksgOy+/Jc7s6BN/yekcK5Qx8SC4C4BLUL69DFPGoA/6BfxtTjPm6ERkzPvUm
3pp+POj+aLee3W2vQxg4jfoJhLMlhTrUZ/RBr82/LSw6ErQzxDih222uyGqMq+UM
bD3mi7tCRCpZc4hRBN8fg2hyaXPG2xjc0eUDl5qQKx9cGf6bF92a7iKaiQsRrZcd
cs8oLMgqLCt3ZhCOrrDm9lK+JXHy4rzYdQQIgqApgfuVQIvPeDP/bVdFJS72zuPj
om+O4o0zoO2CpBQrAq6+i11gQY685jBZpbPJuoWJrDL/2UazABw/Igi/IXkDceZR
0J3MgS/MGW3LQd+TPi+2XLUpTfKB1rQiQiDeFRKF8anK8eDFjWM9BCPr2TiNuI6L
KODSjFXDvyNo38klzfZTOzz1F6HTxqeQRI3A4mRe8jasOXsjyE1veoNJRI4NqU4y
pO2GjR0NTIyILKllclDOy6KpGIx6JOeAQR3FYBBRD27R/kaa6QURKMRy7aL8ifOQ
JjsoDo44h+1N2OpguvUFh/Sa7ibP2pGxl2WOiIe2yxY+eNDOApGQbuAYc+ex7ed9
5ixndR5ZW/DGbhdLougnOekjiNJwGWN7Z1I2H/x5ebc7TrGBPLl+Wgeu1VmpPWd/
713XuRZSH6olM1PPT1h25Hfz5ivN3gVctjBlTLm8+NVNG05hEcHniV2TLzV/bkFd
VUQA6vuX1LjBskbI8GFvGsmlnlUsi6zaiUMr1hBN9C+wau4Rle1bgWfooy5MKtcs
B1JjUjThBV+l8TeeHcNv+tpmp/vcVFv3BChxr+gJXP48EA70k09nYv9BY9fYPXxF
4n0w5H75hVGIoefLWQNWLV0IUVbLCDH93PjHjI07ZNNy3BMgSRk48zh7lO0k5IdV
5oXg++3cTlhHhwvYL3qexEed76ZKqmyumesybjH5krvPcy073mmbG0EDwtgrnIAO
A0I988la29JcKyFCJ1mFEoZFG5DhSTQUkJSyvk7vKhTNtpy39tqyNhDeshL1zBfJ
WxK5CoyyWqiq1jy4khML8J2HwlZWBNSZ4dP0nHXRgXFKN0G+YBXrFQD/tY+b3m4I
HgwyTU+gBvZz6cQZ7MOpI/tFd1qR0ptYoFZ003Y40l1Bvy6sqhKpqvt9iTKheiam
6ReHA6T8n1VQwdu/qwIbj70tdJqs5zZpa8ddjwxrgnMh/NTCFHBDpQu8aMqWJwkk
qvEohngUbfSwFB3PyS7DUi0MqBsqVT+KNaHmUJHghp30wQaBQS2VilEtPmjNa1sR
o5nuNMy9bjW4oQxmrstY/J2CPomGjrXOjEcQPkg5h/SYsoePLEGBWmO8dFKOLCJ3
3k1wBli8jnW09BJphIp/HehovIu3Hv9m+TGUV44x2SVZY5qAiSuXeAE1twiAipUS
J5KE5bkCVJB/zS12OxsYXxJlN0xci1RhyoxEzq9wyWr5oEYfKdlWvSZowDhwLFCa
huxSGIhxgbZ2FNJQeYNXX5YhKVJE3TAtLaX2joOYZ1HhAMOkk/WYg+dXIHVHvRiy
pa5MTccQ1UFww83EKXF8SUF+eI7wR0GwEbMsM9RRN8FSOED5neqXD+aFZ+BwrTD5
4sFy4z9VM/3SAZBKau8rxUZxDJUrVlhHOvU7IEz4SMkMz0VdRjkl3rd4lI9hPTYT
BqzCN5uhQ90/WiOvVfXkzKu5K/ttDHcJynRY2zWd3f6SQEzqGhq1797o/aNxEhEp
3XX6QYc3zXqy7KPXVM26KhiuuS5rjpY6++7sU9j0usfMqrlwliaaRFBsFHUARMKf
Scb9bdRSp/eGLTEKeDBmtuAOT2AhGsPy5RvgX4Ic6JMMSQNnYG0NgOWIWBwXZzLs
g02xiBcGWwvqaVZmu0PlPz43fpBs1peGUl+ssbKNGpXaZqfgyl4ndWv29/kOKMQ5
NWOyIGkQHB4dtmyLSB0tEoN2S3JujRnF05G8aAvcMWXO4tWq+EWC7xtCI1iHXv0s
HyAikCcRw2XJ0dxjY/g2u6GMmz3pxFvk/8DhYr/aZ4ERyh9Vry2iDHIwWWT0sYXG
/pf6bPQP/P9AhzOUxnm9yvrvw/fZx03VguLfMkwIXLl0JGceKC6b/7ku9Cbe9rwY
TGntsykbLWBYCJESldooqKaCOcquKc8KDBBp0H/LrvFYF+TUTNO3yFwqff1qcDnO
12JAxTm/ryDYQITDHtBe4eH4pMdRL0AInCxfHOZoEiZJZGnDBzMqrjsUl2S+LVYH
HCDUsn3A6vYsENQ1QCpdNEmHGDsQEoL5YaJ2w93mhWYFUk39QHBBlaO0gADgNg6y
DTxaa3gXjSIuq/OvEWY2v0S5G7zrcuorh8tEfnuRdBt2n2b60SSgTJAbX9hfe/Pp
7zXRx/gM4Dp0kZT6KfAiBjzucfY7GvivfwM4H6Dagsg911hJCBBkMcYWQoXC3Mto
2wfR3mPpwm1NG+wUaObDW0DdS247C0E/Ey6KjOJNwhWcFEgM3w5wuGBeql946e6T
qH2ikcHr6fDd6ycZKBf90f4hT5kUUqDIxXHs8axlyIOYGhabsO0AhkWErcnu8EE8
Z90r+QQ2VwvZSwnNVWGmUaBNja3rYWcOGxxIVv8ED1WcL4nSO/y3EYODGsdJ7vD1
XCd4ym9cKzx2kIEEV7AH4VR3SSiD/3Bk9sJka9/SXmHggTLYu2U7s2GqVK3baLqk
t34Id9gh7sjk+L9fUsPFFvwpwnVIHAJ8Q1PC7TNbFAHaVmAJj3LM/olhpUaYixZV
vGING6wbuJ0865ev3xilwvmbQiJwOCScD4BMC+9E7gCjk7wc544rAG66WbKznfhA
dCcNKqP04WHyzJzGz770/+6s8gePXddriALglA8L2UQ3dvwQ5h0ABrWe0/8OFwtH
2iZWTzJGOXziE9gQWvDrK+bvFsSSsZHZE6j+mC2Js6azDjCVEeF1nKMm3/A2ha8p
4jkYF3i6qU54kZjhqjw4768SgwfeSk2zn0Btd0CXOUDOUr/PcMnJ00bXZGicqhSm
EXi7pCMn0fi/LSS9oswn4EAiNS6aV1tVgCIYllj0kuw6Ezpl7LfFhD9BQHyRIW+T
5IS4+WCEWUY03nKhYcwY9vI83xQs7u3fQKDM6+HXA/ZQcQ+o9YNXct7ZZJ4CIsgb
F1fOLmJjwO7DV5OejfeAWq7M54VYiHmIza3cPSzcbufmoUoWKP53iRFNffOjw8Fm
IcRH9CCCBsjJaaH4qluDTTMdODLRyfoteyNOZZBMbqsGD7+JYIy3MvuKEboWqowB
qIOjnqQJwPN6VoQl9oSlkZ9cgZBg3Esq9pBTfkfKI/nFyuO+HoAfVkZlt25W/kjy
H/xt6E6Q7Y7aeXB84RY/PSQ8JdCtBH6JdZUSviXhhSJ+ZevuMDDLLYCMWL3HzAU2
5pJHb3zxAs0NCB1DyrnS78l/8cojvYg8OHiSFuaFWh5NV3H3Unh6rIpeRLqRo+bb
8B4JMqcvDvQ3MT3+ib2JsiVMmrJ/ohM+vpZRfhfQHkUF3b1K05u+93bt7Zy2zzv/
uTsa9HKHUjWqphp6p/tFoP8/0GjcvtUZpePY9sgHDFAtQTyg62Qyzx8fsaHv8yy6
tDiysDMSP96vrHK3eQmzz1xK8zeGWSUOm6gRoFM1J22RPzq2dmeiceoXE7JPNvpF
J1BLpdpblWQDFrLxV3BcpAEe4HLe0FmRsPfVuwGvCvN3PU50BV16ShBLmTuisUes
VMrstu8nvemwseLYVXf741UIMm3fCekezLUTRqCZbi76UqqH4mWP+Z9ekVQvc/LM
w7B2p01e9E8tgGK35c6DBdoQHywClspUWlo5W8XCgooRBWSJtvCfd8U3s2hkaCxr
ZtAPY+8kc8IEU/IKHElk2UVwq18RhAf+RB8uspUNFaEL1RZLRgDUhoLSgcwcJobO
+iB+08X8QXVBhj7zBdfqGlFMliHGn+GD7q4GpG1CA6iyY9lqd5X+waQzuNptkeuc
Vg0peHAVCyJ43TFjdjVB6XfeMoY8qb28rf4UuLD2Iakdhezkg2AHSyBZIGXsu7Nr
GbPISf/Cq+STqx1kmY48jirzzGGO5JG5ZAgGhE70zMGXRMqxtcQz0fx/UTSokF/n
tNyMFSBCeq6bDmp/RAqtDEIW2X+F7DeQauuno6ZBSZCGeAtII5M87KdGqT2fz38Y
QB2BKebnsiPzUO+6e1mkomyKUh7Ui3yiW5KPcQ8DKxvr8C7g/v3kdO56a7EaxQwY
gmazaNQZLPF7fD0GvuPgvgwwkp4SxS2TO6jW3zoz017LdV8cclD0+IpWSveD+mwX
FBWT9wvxYou0oaiCNBua5Bf1HnWfCxUvUe51i81yd34xBUu46MKotygbnjXfv/SB
4HRrtTuT9BAwRSwB9hHDM1V6OBL5+mbUPQ2U63q5xH7jSnfbFR2XrcEsiWYotzaI
ZP7R/Ro2XYVxfnZ+U5Dj0hbDPIYApT62BFT312hSkqKjt9n9KLgCxwfo41qGB9jE
S0sq9rjpVXh1NBH6+niVDGihlGSM8Gp4yFkCRu51aBRLlnIBbfk7K+KJ2A8ETlzs
vtIl3BJmQ5ynCrUVRtw+PSSusUMM30uN364z6aeTgpb8ApQH8YD1qWiiiTFW0GT6
ejo+IX2ftvaiQNYwXqS4H0APXhHwWb505j3YBecghb6LmGk1eLHnvcdbOvMxckFT
ElwoCfKlHZxUqBGxRa0wcG3F5R/AGgRJm3CyikkcWb4/aQIN0qNcOVDDZSTkZFIt
c6GoB7r6oDXeiwzTioQsgiXQFyXx+J7IIC8uVimkrNMpxDENybJBRezEq4OyGUlb
nCXPV+JtaUpXhHu3dBmN1+7e1jljg3GVJioODWbpgkEOam5vlz6WaeaYUjteYhRK
QWuBcvtL8es8BprsF4oVPnTW46yJkilA8GgSEqj0vB469wW3aw+fFgoKhiSW0J6M
Jv7rml3HWfBoIsl20dQkfNUZdwwatva9bct6k7/R+C/zLoUcgfPhi98Ed4jHZgag
1jWX9kJcq5N7w1lJ4Uen/aQdBbVRZZ1/G2dauIod8TeHH+Bf+3+pDi0pf4+920Ok
Fa4yVr1PgY9yzaxXTCjdhXiW5VV4OtHa5XwShSdmRTqHFONOuO5ygjA9nt+ahL1/
2B5rSvHyUMZsnhI0IoOSxn+A0NxtdG7d7l2V4dzSPX5LJCk0MefT4/cZKcnmQqPK
/A8/iamixxDl4f/2G4aHljpYXxBcSqQRVDjY//8IjlO8GIOTM4vnSVw+JW60kRLF
UhmYKrRGY6HsUQZ1BxbWbsWfQXQE1dJKANXaG/52bVf+NDxYNBV5jZanAg74l0qL
ce8YfhMDU4k9GVNe7ZqSpNg4qu/+YP8YpOLB3tS2YabngW8ssXNJdPwJ5JF/q0Fn
WR7t3/lr4VTPylUrBHX3DqQgoPhe3zogTDY1Tjt+RkVa43Aa4ScjP4YvGziCGq3l
/flcu2ynHkezo1gIXyAZOj9PvE3LU/A8ArzyNSjKQx6LwlhjVEJYA2AMx4bVKQe/
zcS0thOaAFz7QIC4rJsW2MK9NFudYIj1gGeGoIOCjbvulLtun0hn0xggkDigcyld
+7e7S61rYJiP2WtZEnV/ET4exsx/R4JcqDcBGXvRqrzY9Zwph+LM8wjPKmLzSw+l
UHZs84YWaqvzbpFELnmjp8MNi8gZKcm8uqwPwa/Kv6RCZ8pcKiucMWky7jvGo63e
DkjpCBKvJ9zrcKBYZgirF4d2TTNCD1Dd+QejGia+Ucw+gxIVUJ4RIVJEO5hfTtj9
jgFivAABLP8EvhWIv6vbXmfjhFj9k8hMFLUCnw25mWuH9/sOc34HJyC2Axanwxxh
OxXIpTroC276lcL7K8wB/Pbl74zVjy0dOgtQE6a34FAs/mOK4zdCgQ50D4o62c2f
wlAYk8em3k48W3Ywhf/Pst0cb9JMSoAYeburwvXdT8Ei3KTK/yi+DOJzppZhynRF
qCq0uNO/27a2ojlUfHq16Gt1zMtLfuAEO4mcCPsuG8CrH3pMwe/2ldA/+X3sOnQd
AyPBxR2hzQDDuG1nCbBHjl0RCB7KBYB/NCXebuOPcaTU+5Y3qUJn3L3GQ4lD0+QR
h4y4BYKUome8WIoOUJy4xeAuErSV9UiiwNFJ3rqYKIdrX8RRWg6vLFbMFzM8GGfA
c8SN8zlXSB7YhwCZvDPpUknwYgO4Hd9akY5vnauXJfGCHmyK1Nouw6EVrVyH9+DS
WFXMI+ts5Iz291RHYlOxDruP+Yt+9QAi408sRgaDa0UsRN9BV2Eib+1dMNyCCCO6
+PATYOxFXbw6YZQdCt/Zwuf53YiH7p5Cho8WMqaRgEHC3KTEBZGvvzQe1wKanNvz
ltsJVNLd8lEW1zplATjt2mnYtuExex5bt+vYMa3N704HfW3hH0rkbwOh+cW9pEGD
0a0caL7KlU4eSexurbmHfOwRCkPUKLXCzdTfZN53xBvOydhOdyB7sGA3NifTvh/Q
CsTYc7qWanhVJqOAHCtSXCHL9Zr5Kq7aXKGgUcdecJpZ6H0WdpyK33CE7vvx/hLS
LR3DV2BvCJdwtCHKxA+C1Wi34pEOYe36cCLLSjp017mS2jcSEjWif7eQGlFB/snx
LE/bColSr62OrjJD7NlVp2dd+U3ghfuZOXaW8NwELDwlensrZmtk/6vDEMko4JoU
mOfFq0wBNohNj0PUO+qrPLm9AT3ZB3YinkiymAS7Y0X2X/trM1p/m/kVX9gElKQE
8BLuZqKsWxwfO1/8UghZyqJDi7KN6AfmrVA8SUpwb5EsBllCeQekfqAbLyU54Gwh
HDf2FSYHiPMIuxQlIu3a9WhnRb7X50nZ8hoyIJ2iRHad1rW0mvQfIO1/ezTnomuD
XL9PY4BqUcmXngMl1yR3rscm/xzV0bfa4OB/ZyKxD1BFxM/KKVMfdO4Qd2lD8YIb
0WunEP/MMg5hKTn1nI6KaF+r/xUcp1t9VzDjknn4k/Y5BtH4Y3SV5ysI/d0r/U7m
BFgSQ8YU2HD/z5LfoXzYnhfl40l+GPRRZABHQYgDhdg/Sa5ReiaLqg5Djtg5QDm5
cLaePMof7NQstIMZF/PpxkFUJ48Y1y6O13I4jn3kkgLOqOEjIdPcEEkpV3XTH6Eq
QWGElkQ0TTpHTZtmbSFoN1jfDKeW6BVI36w7+qWHNVxn8fgxDLfxRlr6lIrfTQbb
tiBqgZnzjt6ObZPw1O4jfOJEPpBMCF8aM1Jbn9xAd6ytnL1NgUD1GJJ08HITX/7i
frZyjep9eQWpO76S2FABLDm4mqULklwxgLbbRVQU0ffeakt2MYz8lifmyp9KIQfe
jvHwj4ljJ7qsdNffrGNb1d57pfAALdMy/FD3M4NIPXsThMii9nzVbUS8J9IH1LxC
y6t6E8Dy6nOc2XeS1rmm2zQl6wYIAiiTVj9x2EGN0c+DdYO38dvcGo3Nkcvr37Bq
rraJAN8hC1cOK5VYZqJCgB/hKHErnbO31jgUKihHMkiGZj3gu0qo8cHFsRVT4KDO
0xA5DdEmJRz3CfM9/7hYofsfaORqOIMZ4rwVxFvz5ctQCBFgfG/5MXqjalKRHBpB
I7WRWJ7iiXEdXVmSTRUklJGd7JiDIadDPn9I7vNiY33k342+b92I2GLZLBCyFL26
DVwgQtTFfLoLHBS9P80WThIESUTdXnQq9AK7VkXXJK30ooGcf8a6oyHdMkYo7w2h
ISzrtdMUAR12XyveHlY01sqDk6fBWcTz1kb084wYNaOlNWfiODJj1buxVOR45BBu
fb6jLWGBCv+D400/K0Ay9G6xJjTFlyzxBwoWlpr5Z6PM1jzFaTYMg5344LBD0+55
WK0WZRoWJb9A/nlVVyrNdV/FYVHF+fsaED3Tzom+evX1iTgsVUTlMhvnjEsM576+
nc0TjohIVgeLazYuNSOASPvf9G5Wqifk93BmFXFWiYAAOZ9/T3j0XdT47MhsC3jN
GQLSuRGQUwb3gn9CVZMYB2WOTzlnXq3Pfe1tA7BQeREQnfQsvMX7RW3dBb3okRpy
zpa3XfTn1pgaR3sZ3d0ZQqvcGSRNMOmYu7kZ7uoCbMpNTARQjW4k62VvOpYGRyku
8UXUPHXAm5eUVXf9k8FSl6zermf12nNGu8sKJ1FxLlsCxze6Cj1q3L/pfiHE62OB
c2xMg9xDhAYowXpq44PLAy9sFwrktFU556Cmd2uFDcnLeAlNsMbHe3T9DBhA24+J
hoiRTNItMz35f1wceFAy4AZpO+SWESM/TjW7g4AaK/jQToMW3WMdxaM8kcYW9doC
+Ai0yohmw8Ct/y5bckoKKS5phAvkbhYhMyhZ8v1fq9e0GfKPKefE49LT6hNkGg9E
5FnO0xHa6d/Z9cMTDCBB20cutkNQsawdZkjZEzDRVPbZRw09Ol4SpcVTjAz/cB1S
juUifKmWAeeCfQwRhvnEZFe/QFjtlEWDEFXbXKEY5XHsmJMNKVcf+gl9f7AXmNR7
y5/gAIplm6TAaiQ/fNrFDRlQZuorLHUcX1N8izlqgVKMO9YN5rON/FRzumxOBDZI
fo3SydtkwCaBLGD3eOm5qrXr1ZOioqhRjRfrr/Hnbb/gBmRf+dgkaWLrjWgEpZGZ
0JlwMBY68OMprL/IxD7J+Y3RyfNjeCRnIR558k+v3oqlRPuY50yTyt7C9QLSL80m
nF38t59XEZX1NMBkh+IZldWBCI4Lx+NmpUnvYuZE4AQ2tGaTDSQ9G0aIg8055Oy8
683wYIZHljEjS+hsb9z6z3F+chI/5F6IcivjgPKMQ4g0FPXFdo9a+9WiaucvzH5Y
XpoiQ5SPlw2prhRZxM2BoPqvEldSDSYmAwH8QPkqaKSOkmyyDjTqr6+2ymRi1/c8
sLP7vLBXYYRLdapEP2IfoAIidYwq4SCq/2mO/VAGop7tHvOsbzRnzsCB59nFH8Ly
aOyeALNpSWDjRpzQOuaiN2ZT0kkd/B7PypBIUcGlhPw/ZcVdamgZxN+IfNQpYEnn
DrsmD4hCG1wTBxIhTM564avc+ghGsWcQqQc9wmiD+i5JQLRN7Amkmb58YJniVlAd
gxrMn9j0mz3jJuuT9aSXbIcWm3BbI/Zam6HfdQgILLibget/a8VaH+BWsy3uEYOq
6h2koRidvxhMq7vQdq6tfU2Oi3oV1MOEV6AcyTy2ReYoPESHNP6vEvZACQf0geFS
KEujA9bJDnAP4y1rXBmdlflKI2SKldBUkf4iKstI7dcUAstfuR63nshIWCdbeq0/
O23ghWzFcM8+nbQH57ErRnzmGxY56taD6W5Wx2hcAtFqIZZtbE9lQXd2DMkCnOjm
pb2XwBahotHynSMhReGj3XuBOYbW7g1T8DjJ/xv+Z/GiF7epnUdCXjBuST7agKBp
wZ1f197EidAWbkiU+Hc9RtpG/abSt809SGxPws/QBd9HwPrK57bUHlaNjWSVD1pT
FAzJ9dlkLn/XE8wp9q33/s9EVAS3Y1p7ro3El7KcKWhJYrU+sXeLpkkq6E1JZl2D
P3NhAmwlf7zMmXJfkkGuFcHHwM/C8avHF2QwrbSGcE5PW2z8dErFRX5tmiK4kGyh
fMoB+o1/v2eV9RUGcwmP54hD4YL8PXi+C+fDe9VUjB+hVcQvH0QePOdzh0eXHkS4
Chl9n9pT0GV0B+kyVyzN9BM0HHkV2diaCSVrF5sYtI54N+q5CiFPBc4cbsh3A3/6
rd0M8Y/US4xgSHteu3WVsJlHt3BVCzxbTLbBZPXNQrcENFYy+9HlymY3o8XDsr2x
FiZD8Hc/lBfi0237Me8vyuzrQHpGUvtfKUoeVUF01dHyKBDS03W8czNLyPsCqb+w
r5Gzm+zlWdyq/cd3kogpW7HGrC1tdO7e0NBa0NSao8kUx8JdMWgDkw1EQRqQlyQ+
12ExtSUi08SoAtIahmsR7aHXcdveWct8UKlhfcAfH0rkfgxbz4vMi6lpUWLjHDy9
Ys0s28JHzMDrsSv346+Xwz+Eb7ajVfvc+d9sHD3NizdQ2YUtBq5TOB1atHaZmIWP
kovTWJgGs2h6Htm+pPPbsAmJN+BxduPHaA7T94wG7DQIGChJE+t1bD7Pcm5IS3IO
cM+H6a3ZPiiuy7hcUNklWcSPbWmdAcvtMDSCLLPFLtOWx5EoDu14heCt2V0QInDE
OWH8FX5cl4RpN8ypbVBXA/eFxu1Dg2Ks5opjPyumHR32eCyWtAaJmN6jUwZHr9jZ
nEyeuZQi09jyQ728Jukme88ZzjeBQMtxh1CNT30/c8KA0UvK+Pj2FPuLP/BbwOVD
kLs9lFymGYSr8V2pG19p6+IbX55ePcV5uZd1ecTdXpC3ONuv8NIkqCDHdIr4sJI9
HYYzZ9lMS4y+Fl3QFow+sdXUkXpPVvk7Tav47gZPYQ/CrOfEGGSi7/UP5DwP1MFQ
i3F5HZRxHJhmqEbmdRZK+UZT4md5TkXwitWdWDOx0uZNurH8VpuylcITXaejCAsS
aAiyMN3RCwa8a1FHmHdvJJbCaQIgyJ+hb0GXaIzcuJE+e1iiRKwZMOVIV8NbI/g2
BCxmZ2gZQpju0nU4vnmcokEsSRuJhlXwOqOoc74hD+UND4/rF2atzwqo+7OsdLL1
BuXIySvEEQEEs0F+euqCn2d0tEMONY1RGaWyMytywMjwOR+w7thnbsTo+uwSR+Ue
M2RXiYSeTgr+0LzKJDVIoiuH0OAgymAfil+lzJV/MvDDqaxJaqvkenUn3R6DZu1B
g0P1KwukZwcvEsokBEPLpUzpPR2lGOTSyXkyPtj6YXq/AnhuXrkHIhzNAMuHKxOA
bjj8glqOy+C9bDuREiZ5irMXjA+W+v6VMflFTSg5VaHzrnmuk40TrexaV1kCD6Iq
4Sa1e5R9TXoOAxJeUe810VJE73LgXvTHdEvspKWmF+tkwIbPFcpoEmF4IZlMcN5u
i1/LJzHTDtr8r4bYti4foh0gO7l2Jz8JbWn66Zz7nWx0H5QSCSnXrMotoKTX3IEL
TSftsEsGwxiMuP4nixIUbOmwvnp8MV0pJ/lubVLNEtZs0MK4wlvkTsK0eZ/gNUXJ
CuPQw7PVhW05f9DX1NYBYIYNWLCdQqG8thMsz0z5mIYDY5DFNwhna6tlH2wDOlio
lIGDbut0dKs3XnApqKSGs6aDTzLd0vhNGeCBP8O4+VJD100Xys45HsJYdUcJ5S80
vOJQU7S+DFrnF9LWxCSbTvAYamp4SvisdUm/9K0w/lzdD8XIHj5jFemz+ct6YUBN
w+F5BfBVaqf+UOF1wA0P6oq2WGe0L9paDPWyLNPub6g/6hD5wo7FL1Zw1JQeSccl
DgIMto4dn9Pjlgng+llwc6VruYQkuMDne4YOg/9OZuBzEAHnAEo1GrVwfJslSXgA
XkA4xd2nSZHb2ndGmdw6F5B6GqV8tazkkFRpk6PuRG5SMjCPyAEalMJGEIpZM02I
RzAm7HGqZqW6hVpQgWAj4xnYpQOHAq/d0ARsi2ycLmZ4ByPehG2ZmWDS53RuXzjl
OasnFsrQexqP6/nFV00WBg76hqRYDWzrsXDZG7FtKEWQEcJIBBx7udwHYSn/ivPr
o/1XiqOLZLZVn4HwRuLFsp22aYtWE8QTxC6Eu/z4pIPUMvM4jLcVEkz4iqgtmBDe
t9DN1ISCGmgfOVw8pk9rINIjHjG9EmyJL2875qa8dBiW4SJa2MxymXD8jTgB4UDg
cu3vNqO6PV6kBSMBgzrNI/PX7F2UCzzWkkG2GtbfwLwRNjPopK6BfcbVUzaf8cb+
OCrB/Il22fy8qMKmtxpxG2R0w67ql5poVHOJcPSQY8bFwGOOO4K5nki8X8Tw0WJg
752BIebELz3tNGQiBYf3gLErG8YzxR1A6FIUBfbSTdkSOPLysIsvj5gkxKi7yJCO
CIwvW416/8ajdISuh113lDWQIODupbTbXmUj8HTHVoRAoZuhgJq470qVkCqiRCrP
538LsxMQap/UzLict57LQKA/h5iR0kYlmHAVwpjAiPWqC1IlT+Xz8O3ewTOqH+I0
AxpgTJVmJkxrbqPU8lgUUsIFayVNwJZYtbc6K6hpcCSy6bQMFJrUTFabQbjLbCTU
C+b2LmtM5PNfmuTbcC7tOf1cBwepY3rLQqf8ERkWfKlYwOmXhXpFzu0bRoSmxa0G
QjUHWAc4PCqA0cPWgLPYU0jMtCTwV3faARjFQmz6Cd3Q6CybkqwxGqGn3VUJSGwN
r4emj+cwYZhLtgbRa1eKUPkiBoKJ0sEwcZDzo51xQLMOQ0Xtm2KSHr35RTd+luoG
KfLDqLcZop8VYAPLIqaATlRzIK9aZxaG4DXSZPLpI+CMgmDNF1RIuxlzVqIk3u/G
I9UJtWbQJ67R2Pq8Wgs1+PYo1W3lenFP904WJ5DDox9uiIrTUA048HI484Vx32Ut
KMI+GuYX/gemojEIOxMblEPI3pBHDNeZkYuya2FefHIPLN4ZRv47w/246btXQWRY
zxIv6fTNl/7v9GFtLAwvPso6jcRRqW6PCHZEvISh5t6Ax6ILHmL1vbkqwQ/32Xfr
3m2zq+WLWMKncFkvTP9axZUqx/ueZ2fNywqIE1l9aE3EdRkYyJj9/jfEXOQ+8pcD
TDgtAvPpBQSiMuVy6ihHEZ0biMGvqqtMU+C5etq/GbAG9G6pcMoe5S/CuwM7+NwI
Pn2uGdIIYFJIVDjyk5WDOKf0XWUtH0Pjk5dJqsDdYuFFibpBLvPIBHL/KFxnYsU6
Ba+dP6VaSTSCOwo944nHzbAKYAOOSDFCawS9rP7O1rVcGPubXycJ9t6OwkkuGF8/
8b5UaMd4YWuZ0rOm7bMLgXQh4J0cdIRuRLiSLRQdMwDle/c4EaDyFNzgrhjrvq+g
a5K6r2oqZNUg/Xjkc8lYItCx6s8rKzrmwmEYhUzmAYFK53N83xnf/TpRYNsgKZiT
Z9dMjTdvMRfdPzmfxSZi11Niw2dBA8D2K8FvCOWl62snxjwaqEnthO81w5AWeCgd
j5LXQtqybw3sQbghBsGz0w69KFZrjga8wRIdf8Xy4g/DkGmz6Au5y8UwEHrLgLc+
CHOWf8XyRe4Cy/rjENhw6B8mu78+RiLZByUukwpTQ28ezm/cLcfTbGnDGiRYQfEs
YxsVVVZO7Qw2KrGXL0JRzIbbfqsHN1rTk/H8K5kePM90sLc43PX8eJspsv6kJbkR
t+oM46WOayDdPMGn1TesBt4rEd2ODXVmCkRc8+8+k3frAJWUflq1ERTzp4AauKyP
+TcCattiWDw7unMkXm3b0IrLAUtiC89mVdX5EPMbpu46f9AK+ne/eku6r9INP/5G
NaAEOjzZA/W7qzR4HNcP9uECUqLGL6XxH/6a7Qm8ZrPWAYBdo2DJFheJeGnib+Qe
hCBhQo2MNW9bAk15Iairu9tyCW2GpfmUdzM4giCsDDR1cmvJjmM8gWg6T2y/JJnl
T7LN7WHweyer4OR4vaRLcfTSm6TN0BVOQnAbCzOWgzgI8RV3/jOROvfQa+YEgxn4
afTJiZ8cU+PGgR4w7ETlK79dNudCohRaEODY6Gdiqix6BW+Lyex4n3yDPuiIPKyv
ZK1Csv5oO2KFnlUJCd2lmeLfU8yjgFDk7t1qC5aKQE9tvaH3RUCALXdJm8WWql3b
YgT5XoOpFhUY27G7euMmYFv0XVJSlv2mL2pPbK6HwE2CyvLttmkB2cX/m8RcyxSq
UmkUHmgG8QDkrVnH1h2Td3us3M61Bi94ej+VYIFPf3odWnyMpU45HLknNDPhE32w
jXZQUm3DegqBA2AXUaPeHL1WHOHOfbHIL7RMGvy7m1evxp8s9k5hQsoSZBVOB04a
g7jRMavoGN7IZT0J4+2Dwhib3jn7kx0a4PQ9Yan4dExmW7CdbBppNcHeSOL1HXty
ORmZzJl9gn2+CCOx72dt44rolm13RFBOqTOlNFm3BIXRLJtnOxn/kP3R+IQVCpg2
28EUfKWq0SLpdS5ZM+LuT217jL1ljwI3V83IiAqi7c8sh05UNNMVv6EI+LHIfB2E
2wLTad3NLmFdF/dmy4C5Vs+DXps5+0e7pzVbopqRTSUCNCkRIdYAojJC+0bMGcHo
R+MbQUgxKnfKbWCyc6goIvdEV9ahgdC6Esh+tf57KUcpKySIhx5Ujao7pg1E9hQA
X8Sj0f1OPSq+FVE4wse7YHxxTXohzvaEa251XEfEVbWH3+H5lqVzVh37YypZ6+xR
qE8raa4g5i3mrmhfBDzEf1FAnHtQNgNC+95WjOt416fLFbcaA109ifyEmq2uZ9bF
NhV6VvHYLGWg7GF6Vd9w7LIPKxF+48mOyPNXAe6X0BKtYfGnskSgLCvCwZtIKwH/
n5oFSUTJEMsTcoZT1rdgrbPpterTkBLkL/qgXqBF8/KKa3KwAiWxZEVCw17zAGJ/
YMUKnE2cBP/j7MwAnYbIJW4akz1QIqqae7xob433cotg9nJEcpdrJtfZHCLNTWE8
g3CZ+C1ynOi8nLki8LcBFnwnFS/NF9d0BkYmbIOr7o2K1oeJPwgRztCQTYAMXLMt
Bzx7EA29edYVaLD7DifjFfLR3wzFirKPE6TTiG6fXBc3a1mnjXz5E+K9mB610K5q
phS/+x7aFvyw1VPoXbyw7jlQ7nynBGzl7XU2U6fekFaR/DjOVmF+lvukof8brj0D
C/UZIeBs2yH2UjqWH1gewfLCXt9Go4Mpqp9y5i/uy7SXuEvz5Dw5UpyaifivFe1c
EtPGhk18qcOCVu4Jtak5IXqaKN9M/K94csDX0N6F2f+bkJ3tULqqVbswpEiAVpSx
Ce/nWZUZBNQ+QyKbOS5A16AB5rL3+qKUDjHaYs18KoEO+RSoymO8Blcwc8mcQuPk
aH8thmRwgK73qxs3DtCEXv4Z7yWckuMe/214/9jlcJJXjoGrbIq7Gakh5+07iKVq
BJNsC8tWeBykiucM291kVi5fyDpVHw/1Y9+pOINZPAxvwN0i0MH0AjVPFtppKBmx
KyiGcNsNwxQrLUS3IvicdXdQti8mcm+25t7BMqpT2GYRPTnsDtY8K8htIh+/hk+V
Jr6X+RCUXN6BqYvMUIub/dAVt1hHeZLZTcGjEtzEpfywU2rzdHOaz5tGHs0axYGw
AnllDPz0hS7meuSo2tsaAEZToBW6KiPi8DoSszwkZLeF9CQQ0YuMpR+0aRkmqPk9
1u3m9Zbfr004MFUDXc6NGK050hGrkDBbCsJkurWvLVIWsA0zvRmLOGhsLaP4lZdo
46vSJ/NE/SR+oLGRTD3STMxIuoYdFo91AR2nLLWo44HmGhvme49f0FbQgW7rieZM
M8ychLPJdzby9G97OS+gzVENqmaF6rn4GxhZpxRLLW5iT7Qlp46J/hWgqUSQhu/r
zlTswpjCgDQ+O9qBzNEb+KP/JFozw43IMZ58LN34bejTskE7imCoivHiqltTYeGA
SMC2dNTOCYHym9tXKQM6zTSDcssckiCOsRtb5rMDXHqmwK/+sb/SaH2JJamhobBU
pHRfPcYotpQN9BMMWtmPAw8c1kblo0Ob4l2zJmnKUK/85Nw7+PQ6M06LWBxT2M4h
AE4DhJDNLqJ11yCo8nYjUMcX5ZinPnkW/UNkTCe2Lo9tbjIWnvg/Vg1UmGpKxRWh
qwwG33whKCO0jSEmOBXUBqaSOiwgWdYFvmbR7QosFcZ+T7+72Od2vah5aqzywFCo
s4xb4qvMn33+MKqf5q7BVkzUqoN4Xr4SQZVcdF8BngngWjtYtf1GV4tWcyZGHmW8
toHwdguYi1Wf0G1vmocmnpfvk7DwE3QLsCbkn0DaQOE05hLMNXFizalbPs8hQtj9
/PngxtwJOS2m4QpZOpXkv8rUFKR1UBWRlu4lpFTg/nkAwihm7EvcLimb6LBAas93
EuKgy7a+M4KIWM0JO9kpihT4goBmEA9M7Mb+FOWUw3wDId7mVqe6RoDrp+8h5GsE
GWH0YppAwfX5BO2Wc5qGwYOKVoWFrc0hUT8MqDbqtGiQBzkurQ0oIW/17tGPl9aC
R/v6FQGW0r9NrvXhG7zkkFpG8GOB1PnKGh8VuljKcPz3Q/+eJdMcZ/RUvH8xKHIo
6cFBmg5mdCS4NdvrjR+ed061X0PGWYGn72guuNIHE/up7fmnkHC1DdWLYmUr9v4h
PpdCSjdOyMqpiwTTlAqXE34V0sQv/31SqDOpxLya4IG+i4pi0r/JAszHmZVIwKl2
dYFRCkr5R36L0IWGB0zCMclYsmw+r1nC5ue9yuShGgDosVWdpSPxqtiSyXlu4zMT
9vlpb35RIcMguaKKaJ9T+/HzRnWCZbTISmrVJsp45kfNRakojMtIgp/zfDbf6T8f
fDy5muqM0G6qibbA9Iug+iijsL3QY4aU0DPdeSGloglFchQFLUy5qULNBJyHMLhr
HbPPE5SNB6q9r7WiFJIMElHE9SHq/3EK9VmczuQCOoDXDuFsSOpPJ8MSRIywGWym
4zt7NmmpUvNfBUD+h6typ5TanGI1RSzAF3l0GUn/Xjykc1PE3m2AUPnTzF60RtU+
8vRDGe+ko8btmWuYHb3mKqZS6NRA9tjlFJViWbnFLOnQYs0KegUYHSKjvop9ZccP
mKxZnPB1WA2TK4+d1q2stuOG89X4ybN5ViEcOzI4H/DxRi3u5DMy+x1RxK2mryg4
AKjH9gojdV0AILU2QHOpBFRQKejsnXRhSYCg9ODP5hAeAZQXsltGJ/G7OAXc8Vpw
QfdGkmj8DwwWXtY262eQKWdcCpOFv6+D9AH19aVLWIZtMMW+DCJElx7rEqbx4cWd
cN9B6d01O2dkmCJFoFdo+eRh4wtEzCbyC3aZeTFtdOW3j1W6DTi8nL1Pixd3pNXc
i0JxcVL4MAAUH8dOzcyOyh0dggM11m+BhC6LPwFWOUngFwvTVlbF5APSJkLPcpMk
1XNPJCDg/ZKzNyh3hPHMthjqbmNYi+mlEOqlvkstNkVVscviCgSwNjV3uK9iuzLG
4K+2RABMrX7TTmZE1O5ziU8Vh4Szn99IBpwbHUNqvw0ew0ZXVh9WxpJ4LbmF76ba
8Ds01i5pbDBnrIIblPsBHxOnucVLjZuEtT/hkxvM8lSmSTtxGgReeaGIdFTLWdPz
Bz9RAUfpsNeqklfQ1OKyxJ0N57eUj78BKzUsWz6SsafBOJTc+fQffjl4mtAjhDW2
EBV883avO71XytkKapUOujhWK+UzFZyx46BfISYvkvNuzVsKrgVt6O13YzuhEOyf
KdzGvE1MgW+H3Jv1LqvihpUD/qozz3QIPoKBzOF9ckKGXed0+KFQwXLPs731TBvy
lGYddL59IyIXBARWq3B+glk9HAD/bvvgF+lrar5NtdcxntHUzXx69+5o5aJM0LIw
jHe1emQI41gpdEDz81isiAG747IbQwK0AwEdh4/f47kDnfp8PRItORF5uhaZzFQc
GVwwMbe0GXYZnkzh0kJtdfETPHdClrl/EdYWgW0wztNHiAYy2ZN4f+El2woxN1UW
AOMVWd1qKKrK9wetgXoAWbqvA0iHOFQ5DasKIHj6Kj1mR7eSbMdtLF/CW9yPVG7i
rPgt3de5CBEOl9V3u6m0UKJe1DGdHxVBISvNDvOT+gV4G086zqOm2TY/O3INkwtM
LXVpA21i+pmHtJbzICC5rK6YIpwOhodCGqGZiZR1HJwyYFManEY3NSxPyOAJt4HV
7YcCyBlCP/6a5rsOJnyMenN55R9nsR5U5+e9O3QoqTxH0lDMsSgtJyoCIU/Lh9uJ
IJXZMakaRljaJqiAQRrqRVNgW4RHHqzaT4ex0xtUkmLU/CGQAMN3HSSVnJXQT8/Q
UMHgjgBwp8qPIyuO74w9lbf+FdCwt8mDp8ELhpEEjbmSAxEK43X/d7Hy9lXrDfRK
hBV+84cTw1YuZhft/mBqNsWB1Mcwxp+PFK6QzhH69k+rPeS9qm4WNaOp/C8E9Srp
yeUxrvHtz8DR3mUU3FVUE0PoqoaDUmzdzcd5u7qOI+eqPZT3eIbreSD5+3Io9n+J
eoZybHT3USj1I/zRpBCn3NZSo3E0CHlBaHg1n52XgtV84Cp21Om/JBr9ROnq5uNh
DbEFu9Pzo94iscSH/Px5Dv6cHGuDOgaca5lL5jM+kaE1YtorcipPoTl1YssW5ZJ/
3skWZuLs9shiMjQOSc1oC7jTjY0puF4y5MBqKjPKs/oMx777cQOoCZ9Bac/rFoxD
p+TZQuTIv1QGpNGpUIr5nuUwDn4A0BnHtzHOd8YuJsb8ivFF8kTz/gh4sG4dL+JN
qZcY0KqdnxB9RSEmpug8OXuK4XvQgt6FIK1HnOPV4NZTwXCnywXzjSpLl5S6cK6C
rDxqkz4lu4vkNNcGFzge/1fLJEfEC8Pqfhy/5rOM3MwE74EQMpW3EiAuGIOZto+Z
0gxWhClxYcVVzgw9aAzKV/b2qJbn4dKLNCiq0idmV4hDijtFhL99+z1Y+/9c920C
6eoPojSoiPo7nO8U0Jym3AbwzefPLHlKCJpnObH/hGmSSA98dh9aodLspHWP/W3/
aPogT0ryZNrmtRMLmOsLyD/86C6ruhepPet7eYBO5eMppNXRJOgvY0EkFhebjmDj
LCJsvG5VRJ0SIMC6EjmTa4bZUWkKAscl9iCtJO6iB3fCyh5Pao97qx1yx5FyscVs
BJyBUZ18pS41eSrZbx8dLsRGmy39aFsXmmbZse/6Elj6sMhwaBoaa++5kqas/ur2
KkQQlCAgIZw2hRriUwxFpljZWLRl3aLGpFIkefIsneBoIppeGgLqlrJdgmUxV3f1
H5zPnVQ7xQSNq1oU/3Oa8TzhXebB+Bh0AWNWOBXDAKkEy32ePhK1uBDB9friFf5Q
ivHnZMvEzAV9pWaGhsGOeixtuvmCJuLMIwFrRL/jWgAiUmD3Jzy2MXIMWMXezgau
0GvD0C88uKJWMgE5ccrJf9KeTiiQ1fe+xCzUeYg97znPHyX86ODPBQhPPrK/aqUr
6OW6duCjkcF7bWSwtxEprKyQzDN2dtII9ITXwSv7L+oSGAHj+QyXzgf2TIWHw294
yS+iBaqCv/vK6wnAjC9Akv7p7qVs1x0tJg2dLGbOIGGY6Exj2aTVZLXmMzfI3sHZ
1dPIbYj8A5XZZ+o8rXWg/Y7huv9Tsf52dISxF7gF2M6bCEiE6eRVt4urZActSj5Z
ObjYeGSKIahNPMLXKw/Oi3tTXMnMfavCIpmWAKC212DGSIm4l6r0boomZvzPe43B
gxq7qUJQOk7Di5BT9GhAdB+UN7xahpDkcWfWIkOpds191NXgVOf3mJgla4JhsZqc
2R9VUrkJTRA6W/h2yCRwVKuMns3C1OVoS/5/fng0y51Tsq06wYZTM1F/gJ+4YTMI
zKXzkV15ZG54N2bepSwpjw1lO4F6Da0sOW2FJ/zwznKCOk4Ms1AxAoUh1QkOP4R1
LpAfOPt7K1XyqtbICMrbVOl2fhUMAgOEeC+DBdUap2WMWjrHTYmytdtZlnEq9bym
DmUCg8OZPR17g+MU9YWLQ2hJFiP8zq2wvqCOyLfBihlMDV9iH/grJ24MW3z4R+io
yIto5TIaVe3olNgH0Vh5UgFjPHxUMLmfHYU7exEyjLbLtRXDPKQJrEj5+D1cKI/N
OYAprzTBXjcQ+oEmpgWAfYFtegCzzEbmQTRO//AIzROISUNpJJAnXBF8lufdroIO
0ZeDNryLmg9LPWXMdvLd1pT9+THJ0VT4tZY5xR1NALIBEnCwg8Mzp+EkPbp90VbW
gYkzf0yb/moLPbiunbyvR0ScAP0G9pzSLQ4xee7WL0DEMtCpyld9qgAkPHTTck2T
uWoC6ndJ6WgIrTHe6EqCGpqBh7FnM2KwpbAAoX8ATAlWwGpG/WjJ5scwOqOj+7/F
1d/vuF97aB2K5JfKzqJ4mx6qNqe2SvbNB+ULKh5odc8NAx9xsBjGkHssg85c/mWg
n6iUtKPaGy+bFZmG55BVaHzkPLxu/uvkpPOe7CnXPvZhFDXMS2Ba4UUkPjkx4A44
UOK/oXFLGLMvqXjzTbTSXZIv6rEQtnbkYPD6VwfGr0tTSsN27SYgcSkOrUdQl20M
SwS6VIKIsV/70AWJPd4cxEzcUDXEbSVd5oyI/8rA0WBLB8f3TLgXV8MwDBRgCZuW
30Ju3Pd7r6c0OaVTZL7+dHxyujoX11BKsBAYuGu1CctmzTgHI9M9+zluh9ypxYl5
TuUb4v+7Ts6fI6HKUX5+tR0xlCxsg48tOTSrcOMnJDIQGK5FEJLJfQP3QWJP/+tQ
/I7RfLONBa8G0eH/Lt+6PXMvC7+P1CfpEIKbyoKbP3obK4INgBzrHViazW+Kf0sn
iUAd1K/hRZUrKGCDRhPs0QIiys2rmikkFf8zJE/uhOSGwiyhqx2gcbec7Mp0W3hD
xsTmgoD5fuvd3bhwEc+QTwX6WaOvLM+S3lwRrjUW0XRiz9o9xphHfr26zLXJpQpc
tNRZNM5bXsdyVsiU8YI0hhNh1qWl3ihFc00B1Hb5AQziXYnJdlSk1uIyfua8BeE8
7oiN37e7ozD6BPB+vkZLxCSJjgDPGOCnH+pR2VA2PApw+WD5z6miNPXYmqvXfYPW
JnbhwrWlcok220vc8B6eqrS/3ZxCHEyCx1bEP7PX2v/53G6ptczZjyiExmO/cBVo
ek4+ugW/9n/fzj+bZThJBkKcviIWXMCmvankRaMI/syOXPyXkFAQAiYs5tLKhZLN
1uaLThIoiIuU86sSRLY6IfcmgSQCzvRV7CpLZrEzYNF8iP8ulAxs6evjK6sk5PbO
MJI+IVmafWHKlQ8sckiNs1Fjow6xZeKRbqy65A3xi65rmzFXKUpmFObiJvI1DWS7
PDm5A1LUPJ8+OvpmspM8hTph/+AI5htKWTa5W7c1vr30kZZhIM7Vvcg0plEhr3r3
7vKxW35cjH+BqkiVTkL3ul2LYHIK5MRrL7fpZQ7xGSE+RDZa9C+5dbKTJIWbKFqt
GJktd8e3nVJ2mf66uwUky0GR20h2YFSNMuqPnJy5396RFS/DjqBJZ2mxorVk8tEu
B/VQv+mPQb2LdxgfyessGrm/fOptC5FuiMKKepSrB9oqp4PV3eose81DwtUiYem4
F5dhvfgkvjjVgxFA1urAjuxAsDF8Jp4Yw27jwkOxq4kF+zYYK9y3UKj/pbvyR0Bq
f55F6QtcqNFCZ9qixd21kjp6XbNQvrNu9SaQikeESTOJ4/r6MXVrXdZcSGUD0vNw
Gyc8X9f5oH8wV+csxyJJcO5RLwQSy4M67nxWA796scBlFnkmXvLuyz7lwI2cymK7
jfpu5mxinE3zOLjYl1mMQcxOchKW9/u/kxffgpwQMUZ+MgGxvkHi9V3s6l9RcdRf
mFnYDEhzYGrSdGUhFvI5Ww1FSlBmOxz9CYeswK0ntCWHOy2l+m56cYD4xHJqraMl
z5x5KTaP2UopKLJ0HM5j5xF+zTx9qi/S90zps1k84tHsYIfMfziUeNdLbye5q87+
WVvZx+9emn75OR2FPT7zGikTxBpHyus6oqQ+8pPF9tSdA/XJKIdG/vBWsYGtFDHx
jhZPzxuy001E+7iSA8sEGSKGUmAfd5NbhVXVoAFe++wOoCboqM3D16lWCE2xFz5m
c/zUigR6Rbz3665V2CVywqoCk9xX6p4DdX4uULWKkpjRVonSuyszwjPdXc7jHIlB
8zGVm7sErcYHghUivsar+JHNUYqX6Gb/NCxfpRAizdmUA8wrMVk9a9rpf6tQSdkE
GHuyFiDv4FRIqZS3mXEORK/89TS9IWSf3c78wRjblDDGLH/Tr4rWo3VVbt84KidW
IyyA2sbVGVzJCp6vA9wVjDj/p0nk1TN03gujw0nCMMpyR16cxkh2j6tDmpsYgFCj
YFetCQTwgjdOSb70R+Yf0TF1hpTTAb2Rg3dizBelDi1GorSFMmYiA1iROqIk3p+Y
UK83hwYbNwOlTZ/Fi5eMMYDPm9uz1X9pvNSWqUohLl6CAjamz+2kDMt1iu3RXMm0
ruy8rbS0eArlAUBHu6GZhHEng+oKv7hajYTUmyMWbYhienoX/Vqw5GPUq0elTZyI
NjGV8aujM4m5CbqtfvG/oZwk+R95upSkL0F0+0SQ+LkHIyLxCutix22z+lbd32PQ
akA+rDiR+axckCRfNbWs73KawF1JxSJpvbkPVY13a8nD/54AOmlEX/50gXLvX1wc
M1REiWWsJee28KjykBWXqzq7+yKCtGeZSSkSQP5W6CmkwbpXo4Wlzu2BfGyE67RU
UO49a7UFCh1Uw64iZ6UT+LQYso6+UQYk++HoamM86I33AGYN1s/TfCSv/XhFSnHr
pgfuwZK7keGO/f8bWtTnGg1sONLx5dtQuQjJUxR1JIb4uxccRRnYKfjJmgEOERs2
8QCmi5CBmcnLebtjzTvhFOCvBnP75JuS3HGn2eea9mJyoo234redYj/6obPEVdsY
hPwgPSMHF+LwLP7NlvQwKF9lhReh2HRypCwpLK+KvK1cqEGCVdKCN9/uDobz9CTK
DhLcN08wKvvA/nY15Y5FnGDas81pQlVW6t2ZS/79/VGtSLASTYQDSAJrpgMApndu
ZW7xqMMN3NjwZiJPD8KgGD8hphS4DsGjcAYEQLgpH/he4NvRmbaAx2AKxBOAfxtj
JQcEK+gN8d5bOcQl3ZTuf05HHuHjKt9omGlh5VZLoyg8jvWiQOufUIAediF8J/vC
gy1wiGNOFu1HGmXzgoxlmrBJNfYQLuFJiMfT5Hh/QmNS8719uZY+kLq/jjJGlWeD
WQbQx8+T/odAW2tqLWkTMK+eku1iVInEQUHQomYGxqggtSoE+0G1a5URFe/EX8FZ
Mc8zDqX2Pkka0xwsycQWO5uaMR4kZEjbBpVmag3BhaXhSrGvuINhdsHuaGGcJ+Sf
6o+PeIFWu4IM0m8eS5p8jB4OOpEEy8oqKG/TfH7OvVXX6Hn1lUmW04yfTBWSCc5B
iVmSUSeT1ILG1/0tffVu+TxdbaNr1IpC+FBdR1Z5p4h3MsRK+xnUlEEBOSuim4tF
QRAuzxLKJ4ta5953YPc5+SXT2/oarSlrdSKJarS/pTcAq06SzjkhEi139dklfULr
9qFHNRUkK3KHsKwjUKQJCDzOTiscOnUiwT1U1f+shTQxRlJcQabxFCEqUJSXyH93
jcqDJe7b9HTJ7aek8sHSfmNW+ED6C9mVPolbd/6or+NY2qSCl0bw+Invg0VA1qVZ
tUXCzwYEv2gyMLOxgjOn8hYCA034XNB1iSz5tv9PR2hnnFsjXb3ifd3K1HGXkdIb
n15tK8sxQ1WZbMEWI2Gg+TQ82OAvbrR7NL5JgCBGUrrip8X97/RW5fZ/xX191grI
uUr8Qt8yhJLx9RlHdXjbtDmJDf0vCFnNQwOCDGupDDWyWfQ88iCeA2x2MZFNXWAO
4a5U+0fCPY/UoHOiGgI7MgmSp1KElxccS8+t/pFbLGlRD6MBiRtMSu/qpaZOKXOI
nbSglmsuBGBh0VW9TcrTUzcMyuZ2K9kvHhl9S0/nfqdQ6ZfNtmisutcxWZe98SLf
gbyjfsbMo3ISb6SYdApUeqeIMK7nAKs+N+ROOV7hSO2eW6wTiU4+3FiGmhYxaVta
kEYc1R2SQlrHaAEVWWK6ZpJDZj/Svh1Wr1VgwymsdE/eBl6WDbc7T6la2Sp/KwIt
hS68sBBXhsDHJau2rNYVHAegM7ErhgoP4UsgxukJxOmwLUvdSfCZWZTi50+S9zFU
16dgw4f8hJX9B0xtVZ6qQ80gUTL6+3cDrXN0f2qy7bEVQT/zYGlMvel9FSWYtfQR
A5BZrdKHR/X768B1IHnk8eFKLejsf4s+T1Fsvj7rL6XbinwkiyOh7jVP9qDqC4l7
CnAn1teSfcMTLqcO4Lz90nxtM1a70R+IUZJ19g6Q3wZP3xepaC8/n9uVNM9tl/M7
lAyVFZ/p+O+/2mCU9C3nDeB9iHYmlEnhYwuyQwQnCoPynRqcHF4x6UuUjx3btVf0
YZXkQUVBoOj1gDeMMCn9AvAoO4wEp+4utTCSUpoc9guGkCaXnhkyf1/k9R7JMoGc

//pragma protect end_data_block
//pragma protect digest_block
4vEUsWpbNIvF7JDT+J2IPxMJfLU=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
y/q93aTjYOOST8bAA97RFheqDvr26tXpACVlBPf3EdjUh/q+P0eM+tjIKJRMvM1F
SKr8DjdWnckZtfuR/56tngDPfFvUikuvZD/D7LHF1dMuu5EFK9ylrGG5HdwK5Hxz
y392kf7/h1/Wa7Wk3WRY7+Lqttnyy/OUsUZR03hwwyMRk2+0/Ur1Aw==
//pragma protect end_key_block
//pragma protect digest_block
nAe5QclWyj+gfHZT6xYgXzQ5LQs=
//pragma protect end_digest_block
//pragma protect data_block
CFlCsRC7t2N7dHu9uvBwyI5S8CGocjr1+/KGqEGZa5+LTylrUHP55HEXdXVK6Dno
UvSK82rd6VqWet6npSl0QEcsvNdCFObFm79FBDtmCkIlH/mmK4wxrnw7u99/csgK
LSED8cFvZ6RoyHjR93y6kSV240LH6q1CRQLzhk7at+KwayFOK4vU2MU9YrSOR/W2
hfYAJ1xuMNenw7tc2s+pRwRV4m5+IPnQDVXlgPvKqw41dP6bjNbWSF5gJCl10RP6
L9HxTdcH1IWZIdIw99lHBZy/itFWppsU6I1FB0u/vD1WDKJk6atpL/vT2vz5QRE7
dJrNuVrM0Nyx9ix/YFX7bZ93aBqe+yX+/6ke2KifmiJ5dP78sCKrphOK24q0d4F/
znlOy2qPlxTFr5q+ZlTrbuWSCa9nhAmnWX1pPyBAkywRLkoFgPdZrxy9D/6PNvun
DUVrSJaJKsOqJSXI6/sAB7yL+sNJwx0IJpXHnJaOT0OGgO8LTl8+FB9pzI6GZXvH
rddpOgaCtYRBlYOEWMUay9Ws2YLHYJ+aC28KEY29+bTFrToeK+NP9NKjwBsyRqy9
zNoQbgsE07qmXhzDMXI0rh3bqjz63LtXgmpXHaNfXti8Umc06/nOEj/OGQlV54Wl
nAdUqYQV+u9S8PWIUlTHRMSE0nAFVybIb2SxY31/3XPgcQLlYN6KRp3w5FIxEk0R
dBprFFrgasNFi5+ewsZYDXCZR8B667UvmvY52GxzI09X/ok0vLMoH3oXSw+SrqyA
EmUoaWELo2y8Bpp9z6emcPjA7xwzUE335d1PxmZxDy8=
//pragma protect end_data_block
//pragma protect digest_block
6g3/OzSALnVkiAJSsvR29jW+jnc=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_vip_protect      
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
xuJU6FrGu3pwjrRYLJDT6KZgD4nmtRIJdl//kHLbHqgPHG453JJliH/YIBqYGsvP
jTa+bXznO/pB3EFnmSposL9UZw4qMPRY+/4NdhXHb8wWXSxzCnOYPh8Oni4hNHch
TnTwNW/lKqHXG9RXjxvwxtUXRIcow7jvpm001n8i+/e0okKVzSqeTA==
//pragma protect end_key_block
//pragma protect digest_block
cH0kzLfGLflGXpjPakEKKGZyX6k=
//pragma protect end_digest_block
//pragma protect data_block
Leo0NnoAwAdNodLjRBJbe7W4zgd5Jwl12XYYIuEebcbJemHWiGZwwf6V1fSsUHOo
JYaSGcfd7y4BxRAWT+2LKPOEmxLWo5FJodElpFeh1j62JiZS0I3KM6+CIprf6YPO
waoNo6aNZgvY4Du+Vh25p683m73WZh9Lu3PVwOAQQ7DIoo9EyiQEXi8kaK3XYq8w
4ItKi7iUoTsJ+b7J2d881AcBVBWwDym8BaL8jalf0a8WRvv95ZvZFQ44cqP4W6V6
mAvomHsUNedcHdNbnCWlfitDjbTr7a0vzg2Xcn+Jv+QbW+UgkPn+NtCGmLV9YV3Z
P2oTUwdgdLNWAn4vDOfo2FliYuh6l7WxR9F8tLmUINLJLaTxEh6XMSvgZ+n2/R36
W8Uhb3gpieFI0q/snQZfqLtrgVn6ai076ZWemNOm76LYH/BfgwV49p2SYwvQUneG
o04bGZ20pdIYCcA6YWZ9qwTcMBCoGo9RWeyMhAh4Hky/3y96rvyL6+UAfxIC4qQY
3AQOA+AJhoi9NTdpmSv6bnhsKxqVx9CXM57zJ/AGwIOSoCC7QhRKj21dOKX1DdvQ
usGUKFjaragcc8EMZyjwccIJbFMzZlA6fjQLM0EGb8sJ8wS07ilAT/eYXPWW2LE4
1381pQkfDuma8HoqCE9xZzSy/k48kHk1aFiSqcK8kngkSpM8V2Ik/4NiTUy1wtNw
EG9dAcdLxcvGK3GdgcPiFnkQZGieRPSJCAQnkg/0Mcag/w6oEgPscbECwf7qVZhI
uU+eSxBgttPHrAzDBZ+aBRl10pG10NhZkZAhm2k091+NU4SrelK2M7eAVFjnXHTb
f/h2+wTr1NucQuXJcJpVdXDUcKA4rxzrEDI9D9EEEDOXMOnKuj9Nukz18VEqKLjR
I+bLZi5Mut5wXo/AMP4nT5XmZzxXw3lxXW1HoK82bkkYnivzpytk4cegthWtqMw8
gtzgVp945SRllBlQGPD8o7tb4UgHDjOfNpUfe4j0J65+p4YqUHuC//E2Cve16eNj
fp9URraco7joSOlnCYjwO/2mAkAxkjtx2LzuBHx6hxljpgjnCUfv7O/TA+thNzkS
U49y7PoIli8do1gzy0ANxWAlvNze7Wjp+1Zx4wykGBkT6Yy3a2+c1XePxnTkRQ/Q
EwThcGLL+7GPUl+KjkQFMscYc3E6U4Uv+H3cbTlcveoSHpwnK6DGTvEef+Z9aI9K
BawNw21NYB1n9OvPGKaAFHrbK6CMN31OiSZ5tZl6+DqzEwTnbW7Kc8IsMw2Sirfi
n/ec14LJNfdMQa46DdJkC0Llm6uZHBvlKcp7AX3AuYhYx3sL8kp7Uzx0csAkhgVa
SQUVVzH5xCyWThCTjYKFEOzYxKiw+swZ84W/7L/c5i+Ex8HxA5M+KHFsurLsacyX
DIu+fStj0iNj77aE7rNascaWCfP7Cuu2wHXSGxcZfDosg6cyzUhs3DfQE+awZSg0
subVjgbUO0DRGqp1gFkxG5Hd1gm7wj3Q9G4NZbi6a+R5lxmLztf/M4J9FtFcGquS
FW3STFJVC4QXnhkNVKdUX8bbjThlKqesgmLCswvD0qNL7Lg0a0NLNXpxAjoRLPS0
KCIzF+APRMqLgOAtWtnE2l03cET+w1TwoKvLYbMIR5mRSHLmItTiF2kvPAOfG7qD
3xCC7W3HepR2FCq5TTfoQr1ESbkizuT+SmbmO7o14KUvpprpY3c9Yjr+RQ3cbuKe
hWrmkZm426gbJnnGRo45yJ78wZxGUK/82SbJTV+sJlcI65sC9cuINgNi3kyWUAm1
jqysnn1yELWUVG+7Us5YyMflzXNj8IsR5qZ5d1GfTw7mA0rOhoj7j4nU/0Tq+pi+
t7Z8awSKmD1ltFRWk4kG9849v7epHyu+AAckWwFfovJenRuthe+pns1meRvvg+m2
HpUY7yxmRv319blVwY/4MAlgsz/AzDl5u109bvKTK2IVQGWjWJY4Y31Vh7SsaUxf
IeX1tYyS3npJOBpY1FEdkBvGElUxwspqnBNVFskkVFWtOqNr6S1T9G8fqn81OoSZ
oWWeuwH3WCWh+ab4BATogsXeoiC4A2GrvWZF0yW2gGZdyXYjoFpW2mfFu2rx7hUR
oYEU8IXtY7F8oo9uf8G9cxFtij26mjp2M8hhVDoANQUtPgvQrKg45GdRsqubqM23
d++HAR/Q3iO9JFWKt/CHYTI9MqY6xrgPabBMIIqeTUwI60+3QDbU2k7IaOM+v4Ua
8P6YWrzu175WlMGZerIPHhU3so3m+88ABhn3nz3DOlVJRJQmEG2ean46Dl5MaO/W
za1xhFUWTl7F8GNGg3NKr+mF+KcxQhW4mwFSlaefOQOHc4jU8yTWAWglS3LdYDZW
AOcuKoXmHqSMQsB45LrXMW8AsCfickQUZLDlFXI1+w/MjKShs/aIHma9HhkRSRPk
yt6qEozAo8pnmvCsuh5BJbklR0TofVa/FVo2eoCWA99PE1LBGg8Nkf6buGaEsuT/
jjPMmBTzw+I6Wp4xZv9Qi7Px0h+1HNT2m8kC7+1jstXk+KnVxk5ePzj8HME45oLa
ULLUwwDJMnmH5uQ7AAFns3Dup+f5YZjRyvMKaIbk/ZbLGV76Y38YRHro3pzlfvsE
wEQ5xn0caP6CW7btvv3LTSzOHjJwnT8Q9XOMUzNIx2YiwH1nIYwVSA/VUP6NIYoy
nu3CrP38B8OlUT7vCbSXgL7RloFcz+h1CWKtPh5hNG/XqGIiQ0JvrpN1NJGyTbeu
M9vJaMr/TkrkHYbjBZUazT3kKaKBKr9RRgJUXR5Qako2rQwf5a7SzjMtvF6gOaIk
XvCHbpyX/RqIYgRfQxUedGtOSdqiuc6x+Orf89pa8A9aDQYCoV8RCrJ6TZ1AdxcI
XseXGdcJRph2zEP48i2T0C5gN+mXsOIg2yz60+UtpZX1NfaXtAAUjoLjLsETszyu
A3UsjXcnMbWWvIq+V79ZgYY+bjEUty4w5KLI+O88QsLXXFaP7wP9zMZSjgVQk+Xx
1qwGtFUh9mKhxKXlBb8IobTc3GZEC8GI7hUUZ2Fg/aJD5sNmvM/azUtLhY5g3Rjl
E2+n0s8jxypSYJDDjp7fyH0mdXVa8cJnHF7fDAbU9swcnPKUIioNc+yY3M8k2Ak5
PimcyVVyE/7buT5CfGthOvpHaw0pPzkC6OW6ItDhuPCVDjZXxrOmXJGWCdiH5XAf
78E9iwpvCJERuoBBSwVRYoxzPQh6U1Ztw1iejtr2xhWlLNl81Y8oXlVVtfkgS4Rf
JCwS7/haSF74MzXwyQLLErrrjHIooiByAEOSmu6x/D9JJBntuDRk+510tb2OHhzB
4lDTjbN+nvPf6087IgE/xbwBYe//9bSXg156S7N05MDGpVY2g7v47FPXcvfPhtHQ
KI8IIELO0zfG/kRNSdIdqiW9Ex+6m4MhoDWysVwD8nhKnUsoTT6h+bqFHZsynjRD
DeFpLCridAeR9SX7SIQn4R30U2E3Xg600nS3BkCmyyUI7X4VIOHcGI1OxtNwmWET
zMKwlyw75TX1rGKtNpglHbBNHLxa0yjl8nXHhm7o76FnHBB5lMyTj1SwT+2Qi6s6
tYLOwKUacLmeTh9du5Z9hYkyBd2+a/woV3g+pLvzpXGctVAKK174a1aeL3b5Q2WP
4ikpx0VC0QOYdLOu57HH9T5EbNVtYAeIVfP5rphqVF2lX1vwZJS1b3va+IWmXNzE
KcUt5YxtmxCTIxer8xobhK0fMZrvdLc/kK6AXSsJ4TmJqhUjPxLYL0Txt/CEbePC
jg745mBiRLGMswk6mbYr0ZgUcW9KNBolnBdQVA7WSQYOpDr3/g/4uys1vxkkKjVX
0xOezMZaTRqcG0nxfdujx9QpwBWmbB4YHCtmwpFvy4ejFSfHr5T17oJN4Fp9PH4n
2w64RgLK3Yu45Iy4vatt6K7sr/Xh35oZ6hx+PPgGEL+6SvEJ4n1XYujmbmrYAUQM
/xMhdJdPmThse+udgmiOxekhqTtuwkIBjDzJB7yavNyr3lQqN2sUgvhiNYm7vqXM
R4KBFRvmGnZrYF0zN+qbuWTfd0/S2GmWqL4t4EbeOFpRRGMUGK1udqqu1eccaD9u
mppt8pgLvqMpManRfY5JXOQZgnAecF7EJBJ2jioHjUIwKA3KWcWbhvdfRlqbrMRP
wD94v5uftC1bTXfDZFGbdpkkH2YQ3zpI1/Ijs3iaJ+DdXGJFf82Y/uNL363wCpDY
/GkP77HbrjS1EBfhuzteG9N9v0JZS4FxGJ7D7JSDb7USuTuBKx2mL2EJeFnnFeVx
5UD+pRWMpVhgXMz/cKS6eRp8/C0IpVIwCeYgl4BVbjJkAfYlstObDuccYBl6lIt6
yY0vtM7j/Xv/WNr4X5e2klwNpeYBJEdMBl30zsDn8jkPkONkzcoPjNl1OIKXN6rE
nmLnfml9QRScaplPJOVKv6ZbeSFZJ1H7NpAvUi5Amudd8WrMF9U4HhbUHbCJHtbi
kdGoRg2+zVS/3mzy35Hpgh6nHs9MhSDt8g8ZsvOcsjb82l7icOmYx6c8660bdkoB
oppd3m1owX8JVNAi8sTqGM4LdaaKQqRfuNtdjQ+wOcYjlgFVSPemNSdiPi8Ny7XM
btUS9BzhsMh5WlN8rv+rWJ9LWhlM+shdnGD5U5p0pzSkPh48gIPVI61mBqDpPxZe
VRr24U8NkuWatHBCEtahfR5rJXkKg4iF9zyMI5wmRmV00v2Bp/mCkw0WSs5d9t4x
da87K5ODBnexTp/ZLDYW50HrldGqIy6yDxgfB6L+u/R4dr0dRBn0JzXqniBXc4rx
JxnXOFZmUJLKzO2gc2zol5SZDIiiuUPLU50ciRAleEvXf4/vjzp3qgS7j151n9DY
t+jESaV+ZuDqhUggbkGTgXjLUvD6o8dydEVUYICTCMFHK5FDRotO4XocS3D+PO7e
IONo8JX1bWGatSJBIe/uAb+ixXG4az4jLA+o2L1ClQfzYDHuoiA9Gk30hfHjPyH8
Wd2C0prvMafk6ifWJlpSQIdTg3oXBaYTbZxOhDl+zvZh6xmn7HIrBdBwbiEmu20z
QmCdev/LYPCJjGJQmfHyMBmKpY/xYX+w7LoLCM0VpC54/Pk0b9Hz4O5WzxQrjwJb
WAWx6nyiIbHLTcStu62lrFR7dblWRxhO0Wo779+3yetRlETPwhxcgJ3HBlUMB3AD
NBhdqKIF4DuQH4Y8/umdvZBzmzEo3ptdkvursH7y5+WMP0uwWPXKXYlpAJKu0kNx
rOwId+AwxZV5tvIoBDTadm21+VSG+9BQKGkcfhxf313a06ioXUECewDkdGJqH4nD
b5iykGvBM7IHkHckV/8ZxJX5NOhuJELXRqt/j1EpNXAVZ/uMvsW99U3tQuG8PorN
h3f4e44MVUgYta/wBA5L9ep/68G773gdmB/Pj1J/jsSoJ51ls/raxdk38VO5c1eG
50uRGE3i7wNo4j23fhMRxfKKRHnUiodiiRE2TNt4rjI5VVVzv/1tql3QtzBJgU0b
ekndESkYFTlRQOLJDlcw1jGJi91pu9H7/5V9lsNnHLYwEB5nIXz0Yfv90VC+kkZN
YmdLkOIx9GCcvSdZiLsANHGB/07eta82dgR7KJNAyTrONCry7pejDQCwzfk24sw8
Ipw/gtSJf3keUDGY0KKCNB3lBAVjbWSfd2zLyO+2Czl0oo3dOjBwg57WlbIiiOIu
sS+jtKRENXCmKJGwFqeOJDUusILLqetLYXDfj+NDmeH/ieJBbudq/jyBC3nQrZEu
3znPqux4Hna+BvdX/h3Mb09GGp4ZTWV6t00cGbBOdSepe7nfShbpgnWm0zBCr23R
WLE65+K/NJR5+4ti59aRZCsg3Gyrh4MF+qGa9MtVnhccRfbRqI7Vj2JHcikdwhay
H8ezzh2JMaEsgOLGIl1cvye5aEMy1jJWzMCVan7WhQfTSZFsLP61BJ80OU6SsujX
t817DsPK6AfuQY29Iu21CTkVBOmrrWQbaBft1SErq96rlG95lwgZpoZflo+shsVf
vVLlRyUxqQ9/kx0tP5RviI7SD6Hu8C0EeVqNLKabQzG0SrKQwnRzgAgt6AalVzQA
yHH/c7dgNSDKTlA0lFtApx1iYGhiMsN6AeRUMwupNBB46XVKYnQN8k/OVv5EvowS
0X7mmXPbKxgHDd7yrgGuUNQXIkfTu1QoLR+xmbXKC7F/PGPCeSMql1EeWWcjHjLj
9dPfmxoHe3ONEF6wKjVIMkDoDBwj+L6f5BqjFnN2DewubNWpW7hLOhvenPJ9gK+5
EUiuHlIHShU1K5nbuQHpt1UsWNhkmaNyy+X9HYqmpVkKAn+wQ9BqqwWR4qaEn+7i
Nt4En1B/FeARxFv2oTEaxWlfDw8DZ2FD0oxBPbm1CjFwmXSwdUdojOJo3BeDrAZf
n3Phod0KzkpTE1PLUXV9/hXjJM15RU9rN+b8XkIa+k50LgBCCp58eVveqvC+QgrA
TuTDg43BiYtJRLTTZd6WzCjMKFfPVtZmCQQq5DcEdX1ah0KY2Ba46u9jG9DTWtSY
mCPCdOcwyNxEIGS23AvDcVENJE4VPrgPn+FE+CMN/vn+d5NKAFpbF0wT255zxn9V
iTa3//ZfYXUOaioYbRL1LQfi+Om5diK+xb03HQyp4FF5wqabICKaczJklu36BYhS
CmXonE6rabGCxD9ErI1250+4iL5KwgOe/dwpxRAKYljON4s6lDPxhbJsBVkfiTfP
1YSyY1oj/ZtVNopijNXj5+BXkXAQYQ1nJn4UGnGMjVUNIDMdpdfl+FVO1/xKxCaJ
frxb/aHUP9LqCC8/M77winK9SMKYZTP2/ohKv/BxNoksCIpTOBUItazVSwX2va7Z
JHpNsdtZ0LPD8cSYUkky4creZTSTXQ2Zz9mbOPNU5oTKgXJRpS7KBoIgWkK84M32
lMV193ZsdXItNONEuRk9K1azA7bDKoqOSsRT9WnvmIhMjciernhXXG7GMuHUb/hL
fN4SgzlyBkq5V+sscKeeLXgagmg1lOqexdOHa4nGd8BWFll2U9agi+vzSN1I/LPI
+mX7L83Rrg3BbukIb1KcHVAHGt0yFPa1S8hxDYnk2iWJ3orrMhAYQd52ZWorNP9M
DiZ847QDImTc9vRSbwS9Et0e6F6EoWfdXAmorp63PROwdSymyl98buI62DImtFC6
EKQ9/viVWagGF0H+pQrCiBDaDJoT/FHW+sf1imN3wZfx/pIV5mAmBqHhYwAmKBOj
ZLOrWkgUck24o/zQ9Zr+QT20HVM5wySMG7bzdIRarA9FDyASihup4HZPbMnML0e2
V4snAi7sfqs3CQ8PJuAYn05Dax/ZDlwk+GE3d87RGgQsdmGbU8xZkmYjjsbyZc71
m7ROz9IgwjYZ69U5pcLvLdL4vStr64NlbVw/W8uR3RlZF4hrOsawBtQElYvyqVwv
xiN8m32qJTL5ear7D9RoYnT0hW1WkxMVS/3PsXJJW7s5yqJVnOrKOyHWh5eP0du7
Chpc+WsWAR3Qr+wBuVVU+5qpKLrRynwvuYvWneihTdLm/nLHWJa3eShmwPkrgsx4
n69n4j8KZGJt0nWDhfA/1+cvlkh6vq8Hr/QO2f3/snjV2TiHq6tIM6RdgmtmywrR
zhCMEAOq3bKI2t8xHYqAyIHNJC3cjNJlEuKAKWZ6R51qtkBSnvhA41bAAxi5sMB3
lhMSqXg3rX2p3SSv+Yu2ozm+jCIe4hBh9BXDSaARrnUI3Xl1Y9/6EhO+66Tnu6Dm
P9XwJ+3V9uPdgyr4DmxESREMoyixEO1G4F4z7LPZWFIzhw/vbLaCigQur1t2dIHm
SHZ6DaGnt39A0+J1u1E52cndJbSHGlLizyOX5AGmZ2udS3mA9LCX5kOXNFe+8/1c
i+Hhnr3BhFUBGKfJzh2PD8uyfBYXgdW3U7Ah6g1XvcLi+jjYiV7x/4k7KcyOy7R5
HH8cBbml/PF5NRedxUuM4ByxxbuJiwsKxawvFWZ0sbmk9zWEdikgVNsXqmYvtcjp
0nztGiKEWDOCFM6ByJmrJVpio0nHhl/fpX21REsRcrYsYC5qoK2+G3At+OtRtjbA
ZBCJNKguz1Imdm3PK5qPwCxlksM7m6JYobAvTlVn4BXXDnqmISPoc/jUmRRe1zqT
KJtpH/4IXqa4h2UYB9oa70IEUHIpN/JYRmPsVI/7InHa0z3eoPOO53T0aFumrXlz
X2K5jM6RhPdcgCOp3hv5c5BxB3/x1JaUO6OiZum8l3lYUfincwv0JL7tYhO3q0UF
Cydg/s9JKSGlH1Q/Lc8GqFsjt2uFaBYu6rvaAkUB6vINcxXqC1N0WYcZJjkN+WYC
xbbwVWju2N2kB8Iw7b208IBsznytKuSdAEUf6mI2Yf8uPQWxGl7XD3cBHBzvD494
/LPFHGBFKISQ8+VtL4rkTeLFoqbI6BKMLcEfeUx7s6tlwvaYCCV1YUMGrMgG1xV2
TNN1nFfz8bCgVijuaJOeTajFZU8wZReeGH3q2gSTxW516FuhMWO2psfIWr024D9m
SW9YrP1w8i9K3qc32OZi9m46gPi24cMopyt9XjBZkpO8JdPMNPEgm1mhT5ma46xb
CuUhyX/tYLlVwVBso7jLSOUAxFOOtQ81pwMH1D4A3Y0trUTXZu9KRG2X7oK1BRfo
0spO16cLEom68eVzwG846xMxNvRzFnMpOHiepO1r0VQRCJgiRMigrUmJCuJwqgb3
eh/IwlObOlZBdwtDwXn6/JfWSmiq9rh71UjkE0txxglAKJU6soSPVHOl05djC5Bi
VhNSPmMrTQpcd7QQNVsJCF/L2zdvwWQ39O/8mfuHy8DmDFbvVrZ5R/d7lHtVCtOn
gRE1Y3utaT+ecKdttbrEnI2TkmB00KnEFdqh3RA86gfGJ+yERpkQBFoTZoAXij1v
/dmcXQzUhooo/zvMEUalr+T3mm+XZHmmPPfLp9bHPjobJPpO+tqzszyy6DajowQu
DEBUEIKVLJLPaSRVSLkQwCjISTmcuke2ONNVEeyarZULJl+QUAWBv9c+e0wtn+3K
rOA3wOTT1NRFyOGJAMdwc871knnn6UHN1FXWSNoIWKOPR7ZyEBKKnqf1G3V2hxm2
XF9pyPBc/QnK5FPMfDazFRZA4SEBcFL5GebKyDYAuKu7+npo6LDO+Tw/74H+Amfn
1bNCaJmi45sXxbkzOQiL557zjH2cQq+L7zxhotjccRIEeOBYwpr7897seXycmCK1
qgTeAvYU9mYs5nJ5HVJFEZPXz8ZdSyF3JdN+yEM8VSc59a6MYOjZ9q4lFgLROd8g
gc+521a73f7ghzOXtQcTlUBa2RfSDBlWeg0VanW2jVGVKgQHHZci5NabL9CxG/Rl
u5Cd0hjnuxD+LMowUDUPCQVK0I3iqn7r3NxYXpLHLznESl0WauFy5kwcTQLuFBhM
/3ssDv+cIfV748FLkiE8cv5yM4WzyN55bnByietQiHG5dCazlgV6UuKBBt1GObWy
CI6MsxdE1uoELNz0L/V6TkoNBc7/++R2DQat+pUqu+mgXs190QbUq5cVa7PoiV+G
IR3wcWhS5Dep7Ep9ft6u8bYjy4lVxrB2IM7TpvREGCnBH05u8RvLUbbMEe4XV1qp
C0p/MLgsQ9UjRKsj0g+kt7e1ypgH1PKBRkfG2ZVlHaia0+aHrRTatv5VB7R7Wlxi
xC+yiysm8TA7IBndKjVBIZivYq3qcRLvbBan/TjyDeOjXQEhwm6U6tYvvF+T1CUV
gb6P1uSmKoV/buoTPR1J3iHt8HZGlghMCeMJWtAGlPUvWuKJ3zOHU1NnzmfC76Gl
eyy4VbNqWRkN7GymODNcoq6cAsm9gsrN/1usJ13Pa9nh83YwT3azCFL+0OiKNO52
PZSsznr8uQrIr4prv7MgOTX9MY8J1/KEFDZKyBHw3+ViqbdT1I8ZEAB4iBN9OM01
XlMZwcVK32ekjtXnxBRRSB4KOOccevD68ledivn+eLGF+U3M7UaiOjJj43cJiwA9
O69VhNoBXw7PT2Bv6efuJFZ02UTxKVQq/p0rwyr4PN5rMy8/G2Xz8W3tIS3HGcYj
ugIAYqzev9OkmJsiKeAgeLoc5AulLq2COJFyqdbDtO2H1TfZGH9/mO81r4Zt8Bwy
7j8qkxeeBpetsw/kvazxtTPK4NIt/19Z7hXETDJE/+kKz1qdx1RP+cz9AMA13xXd
FrrpwbTuWPgrvC7Bvn3YFMIGXQjVZCayEplSPS4szkPvob0KbQOrJzMg9I/w5yTb
8FUENgOgOEHaikof1ODKUNjXueDE1lJfBBNVFgnqTFjL2rv7aSqQRBCLBOQ1Dts5
f/0yHLV8FNwhtvD6zAlTeNLX03NPG3kSinwhxQ8v0AlqcUXUyNmoUL1pylxuP65e
tlYR62Qn5u9VBZmZyt9EaTE0ksHxm3WW/MG5WNaA2FyfUHf89eCP+FPogmAG9Rf4
gjmOJSEGGZSyr8Ju5BvESkP84zJ2YHlME/KuiVlEGYzu6qZNTRxet770Kg1XFYyj
0LwSjsTRWEkniZLuFOEbFBi583LOkyf/VAthEL/S1OGZfaIzq9TDrpxKQYRzeovV
Qn/Mheljq+vJ1xLW1XUiU1FtYHbbh/Rl5/4jPE06YU5ZwJ6xhFMP4eF3Gr2ftiBt
kHXiTc9YvhmdHBQFCmPqpyBXQc1tqSgQjXZs1h9zdBb5Y4+cenPX2pXtw6WZEQ6Z
jo313XnFZuNBhHuDslXyNlqvG8HdlKlgtV4nTcmgkRwo+8hGhWJAGZGnqIuiieQw
IzEujyg61J3CUHn9Dhpvx/0gTAZk1Afra+r+9plDGDU0eG6kEgotucBfhLw85tSj
z3wYAQoYcYqRyrflmwt4kr3spqpwOFZDCB9INGO76ySDWBJtGlJS+eKdwL0AV9SS
B1nZxo5NBQJiQsAtcGWV/Tybx9bj4WZAE/fo+CYunkTsV9Wn36g29te3/Td4aaun
XqTLAzorP/CearRQDGMTSfWzFDojgayXZxUUsVKE9vw89NFwPlRHeKiuYmoEKPQ0
F4aWQ4O1d06PN0i9QPrATiVLpcGDPw3a8ThcD4qOCw3kBIqAmk4JOa7J5JPK+Ore
zBmYDCqy6+z0XSDdroUB23YS8hJ409ZQXATfvbJIhZ2O2Q2/ynKI4BEPM4Nfrsm6
zwzXVDcnDKJ/OTHzyRTEvd1lkmPJ9qm3Ujo/8drBe7H2xwLAR7TCJyD1XIBe/8vA
Da20oMj2YSmmAfaEPhTLjLt9132AMH/gJoMBdVKQXwaGMGSLgQprpv1xmGy08+uu
7V3S5u1Y20d+LPHoHgVbNN3OdfIrJwSajqlUf/YaHBi8lx7eF1+u9GmmfQGOY6Ko
PxbCf7yMEagahlM1nxSEcHQZiyZEmmBKY7YxcTZZ9vMuMr/76amBwtTDULlKp/qB
UD7MfjxwY9RarKgTwCWz57TDfOBdfQe/M2jzL8B4+E5dzxqu+m69nxcZywyaeHo0
1Qj6HMIfT1xvwsxNODCODoqbdpbDxF24jPEX6PhVTTKdmjsGv949ewmMHvX7Fyxe
XJpiyCPCPiwZ608mTvwkEuCBG/5VF55c4xcgKU9D4528fo2DD12YcGlUSQiMi1Qw
8SC2VItLJ7ubBZha1KWJVcrljP7rLE+pOJ9+UbNGbh4QcEU8X3+pZQnZv+yrHDw7
l5E6rvUyscMhOgZUrhiBYBnG2MLHhJhZoBFxpH09UxH1DayVGWkteWaQM+0JM/3G
h3FspBT25lbM07I434vAd62GNQIFJ5PA7Ql7DnlyX/CuuABoptdX16j2e/Uny9WV
SUA0XPXERLrMjhvXw88lFWfPd2ZCsv0JDw8j81T4lZBqTPWCUVH9CXmGe/p/s1TD
vHYasgMwmMDfQB5Cclm68GfcFClQWsK9w5WaEMA15v0KAkYSbiSFfDJm2oOqNBE2
Oa7Cr4nFeowWgxK8NV/LEn2vRnLTDA1dxRYsIkvdsJG2I1NBoU2BU93V3yYiB560
dtmgC8vqyhJi9QCFO2OkEnvXmgTHRnHHrdiZqBb6tMFlW534449eaL9hXASEVLAh
X7q0YfKb6SKEUpmLTbGt/8RmVyEG2SWhgejsR5gNBsR/7H8I6mghZa4KcB8/50aU
W4cSnF2ke58Hzjk7uqhnP+1aT6Lxfxn0/5k9tebKrAi3Vue3eXffcfJtm/AwXRmJ
Mnz4mCm9FFTRlQAhX7uw//e9MJkAgKzeTWFy//f3tltEw3BmnK2jsrCBTdW1l1XU
w2cBSqI76LkK8dkVyuKnAS/pmzjwTzE4p/+oHmwGVx04sNZzeVvoJzD6mj8yVt7+
bhqP8y1MJsgEXNGCebctK7a/k2xR9DJYoLk8NHCFKjZlppQ/Jf1eAyDkMWVc0Hov
ULLH1/gsoEhXn5Yi8Zlu8mmu73eYd4D6pvPnzksDYr+k1vENAhBrJzg3sNsxj4PS
+ZGCvp+MQ7gGWA97LG5qiU6vKNM09fd9T7fdSv+/dEgjSgxjXzCqIyBqVfZAOXCg
rGxp73DRxZDmg7LrNcP1PFznWYadziKeRE0lYfrJ2lZU9NJciSydP57UgtVEYZyS
de9Znb+LBrGVB2zsGgZzisLA6UVdM2Z4dEf7O5X+32cKc6jzj9foDtNQGm68MaaL
CGGYqbdcY2XtrviCrWhuAXK4NsWrJwc1KJ0xjDEFpG6IJGtAMKjsiDJOyt0njub4
FUdRKAq53zA+bO+b4+eVQ+xrqfjidutWIsnry4Vr7v3ugYKFSLTatfHC6WmnxrRP
JDL4D7yis7F5xRpgjS9LKVBPOqbw9FrpsKVenZ40lCRsU+kJ4uKboPVJSwAdrEQk
6DTJ0oDo78EG/B5CVkmKzUOL+IQEF6g3hBrtnKyvkq4uRAOpEaUMdu1IntdLCupx
bXBEjF9x6xLyMXrARR+uwyzzHdSNjeZCFtGk+87DS7HdLTFhXzVLVemmUEBoEHaS
il9MVQwA3JX5/YyC7QUhht7nOJ/soBBmHdkOraV1fRUH6WrW83Up7rxAYnSq7ta1
7c6m9V7pnxo3RCKtkhM6E3osMQ5X/zRIiXW+ZaPHSn5z3CzwQOx7aKpbHsppG0Xo
LYr0WYnhzPPEd1NjQmx2c4A2crAKlwiqLsCA2X8F0dNcIYNXfv68bUX7OjnTiqcy
ACNbM4+yHAed43sAV3sTuzX3e+Hg98DYa1CrR09CKyc8kCDrhacEu5IWVllPXjN6
nLvYTr5exm4StsfMeEBF81RR5OjR+RnKPL4MIIqWOMsT4nJ9D2lDtcrwO0aPoa/s
xr9ExHgFH/XnX2AYMS86yUKRpgY7AR1at3neV+JyBK1ChYxe/MVu2u3HGWYbHqJB
0tb3bQFxewTMkOGVd1HNbpLm1xo3xwXiEjTPcjqWHzckSdhK+ctkm3y+KvqeodGM
y9Owl88L2Z0tkHsUvb5yxHfsJyWQX0SxSBwUP7LHOr+elKvy87TEordJzl4l6xou
r2EKUwobludK8fMRdxwYdDmzjA6RtN7cJSEdphNH2sbHw1f++DYubdHCoLsb7dLv
ghxxWGZYiPp6I9uppjfKuX8oNDpdruLUTvrtK8sl5CANiSHecS2M/9kfi0vUB9JP
LH/SB5Po/0Bd6RvSY883zdJFogZ+DPWfeaa80vQtYGyowNXlrd15ZTp91ajpb0mH
8CzN3SMe/3eZkWXHndoohPym7RlChcb0ysrzB4I/ndmDkLOu165oODuLeFfHRYtA
aWvnRBG/WrIonx5QJGvqgjMbOy5slOpNWpM4mpF23bcbPhhqfp4dC/TkJedPQNGd
YLaS9xMXl3Eh5w6ujUga+wro8qkW15xr2UDA5RSNw51qc2HnIixf8Y9d2Ptxjaqf
jmJAlf2pk5zbi88iqQWAXqOFmeyL5rtymu8aMKaI3Nx+oP2FM3vxy9mLx10lS3d/
daXVvNSNVu9D45nnwxkM+Hj78yOQ9Ue5HbKZbmgDtKf+G6JtSKtYAJAEuY7uGLF0
jasOwCF4EjNV/yv9el4zM7PullDdCqQGF2GvnWbU9a9PT7jUJZbLhes67qNgkdij
RwjhWOpaPOb+Qqtf0o0YzhiAtcAajKbfe3UiUwAm8p/3aycyhyRdfC5WSOcmfQUD
52MnfsgPo6tiKhjRf7uASPIQAPRqFglxkpAi1OJH00WMyaB3ga/Q4+JUe7Zg+erB
gzpj8dobGS3fQeCd86oxTWMjEpoSLsFV95BvSk5EJFDzCyYqar/+YD4zkdgr+6PC
TAqpyo7hEz573kSDgRaPRHjk4GzjJZXcJSjuSpXcURMBhC/STzvCKFwKYYIXf12O
uenLhNxCZvB8slyDHBrm3If7FD58ouOr7Ck2itY0FbqP0ofm/ZKcToeh89n5tuGV
Q0rNHFyIQxsIiG2sQpTMDpMrRgkZy20opQU1PzfGRfzdYU01Y9wKlMUxlMP0G0nI
YLWqdELbuDshx1TKeXLq44dqz3AZYLI3SjXkZVEIRvdramyaPmU0VcAy6IHJ0GyW
580NUIIdxEqUCso2BJ+jxlHIGm0zTOkCS3VKEzpdMhxUsO2r5YMXxZk+TQw4fR9Q
YdWRcGXJMs0zAv1DpTKqAL13GK/BKjCwT7k658Jrq18YEBt0JLvqPUQ3r74R8/xA
CqotI5t6ubALDW9DhWMJsa17YKdjaT1F62sKOrGrIaRqPf/fe3GrLWMMQELPYMp9
Ho3xECd0k6mK3yaZVLY9dXQDiIJQXo8JAnhZyitCe8BxMM21N6D0cOFH+q6YABtx
uZjNyEGeZz0sPy2YfKxcIPqfztJPxKbN9aW6ruF6b9tCvDLbqpuODByJwNxMZsNU
nNjxPUbM50RG34v43pjd7i/pRYZhLnXAHFHy6kmNAq1WfR5/W1HSMd/aTqElNm8S
mu4dXoYIffsAMiV5Hy7S26DUHLqR2yFqhTK56epd3N8gu1d4Dj7WLGXVTPZp0RlI
pXEXI5c69K3695KXnlchqHByhaoM++9mGlVqieOOOOAOQf7on3clfcIRgOpSwTeE
eS/it17SLiGI+5i1eVkq7rQVk7PRW0sryv9QAQuqac1QMG8AKoFi9GnV3niw9CRe
oV8VWD6OyQHE5VWFVIavk0lHbyHNMG+gyYCsesxE+I+haTTQorzs7Ia54GwLwczf
4fr4iMTC0qM31iGvfm9Z2MWUleAAp0AzgCNPWrBO0oQ+dzmXuXArBCBc2D0Y3rXi
SWNeLqkVpARGOPnjpidu8YUn/mml5JVDAB+vbfL8NDYHc6z0WLdM2W9y3EuAQE6F
jvAl7LGAKU/BormCTMbHGv8NbZ3nBV5hA9Boc6qwXRd41uTQsw0ojL+f8ai4k7EC
SWQCvFGsRvvCBOhFqpihZQxVNjOlB2sO+lEn6i3OPcKpNqe2N1HKlOTl4ih9fYcU
00PKn9WPOeEGNrcgj+ciDkJfDe/dj3gjbMUOTVcKmddDtYg5dRl0BCHDV7lZokNd
gKO+Mm8J4/rABpOYSb7xcJGa2Ys0BuP4pHZVuMAtDQq22VI5xue2UdHpDYx96ThJ
DNV8K1qEBx4u4KwCqAztS/NUrh8parWtLto7tQQySGbDj2XeD/+dWizay32oW9vK
WISSaMM7nra8Q8dyjMJ40dzTtHeUgk4VzLG83beFPiohWoHnKvTaD2WAqaOATBSX
2k3feWulQRXCqbPZGUzeGCTRIEcL4vqbGjbtNKv+O1CatU2XdV34wS0NiPZoL1pa
tq7NLjDP/stcw+8fh7KmyOA4crLpNtPnFVpdvgI23cND+KZq1L9wW0bWhuzymtbL
ffxgL2215l1Gw9ghjogIJePZov31ljmxEcdKOyL4lQfXzmlJsHDcTWo2yYApB4il
rUPymUe2xDo27Z1PE47nicKBmF6p25O8mjIMk8KfayXJJxKUtMKIT5j1xVqx+qSr
ZrUWDoYkoPGM7nDZ/mOsO9nMmzEJmZUN3g7SEM97U3mLjIoGJdY94idu+VAjyudL
l2K6A5AjDI2cAy1eLEGBrWpHC0QxzyQn5GvNvF9E7UZMOfZU/adecfv5/PmgkGvU
UwwtvJKu4TRODlXWi1m9cot6z9Hp0y1npLTc5lzRR/o51qRT5S6lzm/Eve2pR0GN
jgKMjYRTVbeBsTEgaU7htr7HwfB5HzJSUl4EIHbiDi1lI9fYxaTGx7RjxAjSJi0i
tYdstwPzh14/0dexvQIrjHo1eWwcbgzk9kYbHas0aHlxHFhlR0U3WYyoPNMOeCg/
152l1XM6aHE/kgCOM6/tnXbG/2puttrQ9AiEqttjtnV3HtO7mKd3ST28zq/0KtPp
gKnNTsDgyLLvCXJPuE+OLA+7a+bFIWFV9GD3gzdVeZ6hHdXvD/skWYdUS9Sq5UDP
TVoJC9JimYWoVyCTGNPZfUz19M5y6/GfRuXLSrl8RSg4Td5cdrfB4BeOl1/Do1Yf
2wQv/ZUs7emC7C348gnV1hlmH1e54pXxZs/VsVefSb3zmVxTfbqL12JKYNTR6RKk
aTr48y5BX/6lPrsFigbQWaQWvCL4Ju07pU8Zj6TKLSQ7UEip+BXgKt6MGb8BfnP9
XY4kXD2axnymTEdRuNqmE/BGMjZr+rFMSELdbCG61UmjaDGt2SkwyIS0uFBvso2g
SFuM/qHzZkC1lNnn8/5EsUX/z3KdvgqnnKirBrwrl1SUTODlQGRdpzZ1Q4PFcnNi
WnaXygQJnrnoJ+C5OJIwjQh2jGfRJOsVtuW5bJuMDigoMuNk+AOUrKAkrI3dX5g2
JjCsPcPEJc/Ra7gev85+dg8Zk32GvOHbshlOubvcTOB766+1aS/RMFSYk/7KHPuK
Bg5C9lASDOTLUSsw/F3tJe7fHGi3pIowM8Vp1z36JwyLOmwiB6RAlt6EoD1BoFAP
C9Cw4Ia7lO7ZLNVt28jl1u6ZwMSdJYYTW2TkBn9QLWeFEbrou4Vi1DIeWmEmPzSV
GTkUB9M1Gq6qLKDJVduUbkpyFQdzp/LpTUEewhiGWbU9835JB+8HZXZkM53ZqQIz
q7znI0RwWw8uWMroB0H+RTx25258MI/71EStH7op7MFdvZJPMJpjXip8PK56TgJ9
X52FzvwobjJTL7yrRVh83DWuKra3XI3Y47Cnh8FKn0KjT5z1gQ8SAblEeN0bWUFo
JkUOYI03+w8Zkix/QA7r2D+dp/TpIiL15kY0kvvp4UWVrm2bqEXCOW6JCd1yydEI
CU5Am3JIJ29XMnYuDQaxeZ6rlAJU7VklEF+tgt3mBB9lOlpcWdozwGS4Ywutt4em
lptb6bZTVWiQd7Icyoyq51pMrm3q2vYEAVq1dpr9r9IuEe28Jt0nSF3WpVRSfx8I
QJ5v1MfKWvWlJRGQmqN70AbvgrmYLHb0HtjJy2fAXGtNp/kjk4y53webS3j6SlzO
f2gbQK29GPNZiWALXjfg168bp9PdiIEouFn+4HUjIqftrAlAJSieu4az8GrhOBeD
KWzskFKCnKZ7YP9oE+c18vq5GWExRPAPUriaIlqzw1O+iN0iSRqvOVwL0N0hUchs
hYORtisgB3tJrUvTN87KHCrW2NrG3MoizT0yNNfCSTUoD1+FgBPr0hTQOkBNp6Tc
4Wg8NOk+ubk9MenkF7oXB7PupBuaKF42IkWjzL8QKY4KHnokIaPtZaxu0ON9WRkX
4ffHX+HC1rs3GemICcaFrlb6hQ0Vw6/PlbEBt9A/QAKxgyJ0Fv0eVlo3L4dzG3Zl
vRHvmUVTybhX7ehrXrBasXWVo9ou0YQmgl3hFV86whGB6Bk8XS36NZMNFE3FH5ZS
L8ryUiMqpwlE5M+4nwEFcT5NXhO/7IeJIDiVSHIk5B3d/ZE+ROEYFTsQsBPDRo8Z
iw5y97hx26Qx818IDMtN42pycdl0ZuNzJvUDgKkUzcujdipYT6pSWwGcBokSFA/e
3t+3HxEARoEtQep6gt1Ay6+4jhYQzYiJxx6mnVqqqqGQ38C2P2qzwAVxp6bFvHCl
VeiGX7+7kJE3DVo0++qZ6ctQ1wtEG9DpLgGeBRfQ4wdyF+aZ11ZF45ZPga5QFKB/
VyXRepOL2/EjzkPWV4qIKQtUBVKWsf3GW7xBW8HMHiphzXBHfs8P5P9M+a0LCOpw
iH2Fc7oUIjGgCkXM+OG+xLKWG5pootEQQEdiK5gsy4xZrqUYxWUozSr9NUwXzaLR
eFPUTO9MpQbVMjYmvrv8rv/CuUKDdCW4oG+G5Gdq9FCNkuFWd0JXVdAWQpGd+Uaw
PaaYYB3rG4ClAO/eXmNYy2TtDcZFfveHhb7gJ/KDYmUXhCeKvCPkCk2/KFHaP2TU
cezkf/ZuJ9mi1iTh1Co4nDJwkdEu3z1koV3MvzpTIwwPqJSEdguAym0xw1/yOJaQ
Q5vq9t/WAlGNFiTqsExmC3Mh02Qm0x2pqg/n3iptGNfXPWZkDASe/H9gwGXGEAgU
4SvlYN27ibEotPokVUHzHEYkWs4sYEUrj/XDGT+6/MtSdaIl5I1dqUnXD/A7Wo7Q
BmM/RUoNWxB9lCG8BLLbGbtEPTlrk6BzPFy6fy/GIYVZaQvmIRZHoapGoqv/icfZ
9NzlPhYa24UJ73auf8a465Kxp3P7eAy/gk6SZw513oJSNZpjGgK6VRGADAWRwiaT
PBmO+aVpqDlSiQ7izXSfvG6cACzbjUVfOSUVg6I/O1SirWcxh8skYt+OcBrtkS5d
/9n+mx0xApsiLHo49thAHKAgH+qphwYy9jjtEHTS4+7o9WTcGvuOPqnXHVoxV4aP
5OSaEZjjdNrbwgb/vNGEJyD4cih2E256Hcun85OuqZFnDe3zHnKBfCCQNl8aNtKq
eLRud0TzH5L9nIrCFufjWPFvzQH8U+Sa0Fi8+diZ8sRtHTPGJauh2ibda3Jkk4xd
JmGVWeP2gnECei99B+e9cOb7phInKFMPZ4gV6eC0m7a10tWPULBLx4elnZGgecKn
DpkHxc0Jf/jUouo+sVFqNeoExJXDWE00GmzfDKhxWlFhBPaZK4R9WaxOysU+tIAH
1wCTUhViS1El/3rSbHyMwUFAhCbmR1JKk9KOSG21Ij522WUiOViyjQcdP6cLC2TP
peTT7ahlzpQoRbaKdVSHn6CMuayoOEngWH0NW8lSJTXoAeI2ZcPLMtryOx0TYkFn
i5qA6R6TAg+PnRj9eVWN9CMyBoJaJKMOt70y7LXGy1PLjLZtyT4vXGlxsFa3/Bjd
/7OUjZFLDWE8fVjrf/zrVSg+WxNSpl1VMysuXjNT3oxTOCKIhk2Too3cbB8s9jIq
dz/Y3iES8bbJirS7JPhVB6/ale7N0yIGxfBFVq3u31HhS/MnblIoQHD43nnnXYPZ
KXRbzQyrW3mgoN1PxOOB0CAhWlzQwghxUkzTIKnx2/n+fzowy6nxq1nrNgF5rlV5
+cgzTHQgyn91Y9qXH6Ae91kWMyo6in9musFQ357uJKDPxNrH5tenq5cX4tIW1E5g
K1+I9X5FNDTecQhcEd+W7LtHCBtnBdRTImeoFINujtuFkYXYNbjhUv/drNJAlCUh
lSN3jPLzlOquidF51azLcECjMgTmPsPxQMf2PPPkNV6peLCGAjKS6iXtduedV/Aa
1OKWCjjI+QRHnEbQRc6gF/dfz+znyVpyojA5YzIpEZL0qJ7slS7MchPMYEeECxju
slspF3BjjfMKUVtIZMLjIRp0m2knvHWPeNvcb5o2UVovUuN9/JMhLyfuhgqmUHYe
fJCRI1OUpvomNJaEtpv8JhY8wrtS0kbxiskb1wkSlBfGbM54CnPRfAlb9ZVMXjTc
PUi46NyXB/l6utXaMUR0TWg2X+iS7LfzYUK3A6gIR0OGWeXR7Z8MO7T1K7bmWb9y
ZvoGrs89ZwdSBEz2EFYmBX6AG1szgnwM3SH6KfbHR2G+eohxNcXBCri5Tsh2Q+W3
LnL/wgZ4vz0MqkO3ueyur2KWa33POLKDoorkN9DEnnZ1hjU3JGNWkwriwtMXMaZO
gGdNZse4CfFdoKa7XM6vWDRsvUlCik7QJgEfmlkm2cfZ9JwWvGn4m9MzySFMVH0r
aTuU8vhgzlArcjHyHs+MXLGZqraR8fy/4iQN0HR2ClUxE2GvaSP7sPxt9SO5mKap
X/126c0l0xFb5V5HetP0OMsffZgV0ZpIUfFv7DfEteJTfo+I0EunJrSABMpi6TFi
/3/t7acAe+atS9SPgMiOjT5VZatsmbZyW9uzQtmrwKN4qMzcb/xM+kOOQGuWo1KN
NeilTDbd4+4J3r7Yjk395oB/LhYTNxs+6h4BG3d83kRaiqyUlyzOmPLo7PVAkCTF
5EOTVkqvy2DH9ZVNdP1t3e6PdRRTUi8iW2b+6dYXdGMB2gB5Ott+0Ezhvj657n06
VlhXXjhxPsYFjco+Q48oSXsV1OSE2wBQc9lsk+Ms/te5FvjubeC39T9Flej39y4P
LzhNj14KCs6M7ZCDHeyq65PZ7dzLCxSnvYLToQF4pwTUpsbuUdU40nLE644RyjGe
8PM0HMm3cf5LT1L6O5EghUq6hlf1qYhJjNB4nLZYZuoIy3FAvJHRvJRgkJgPQUhv
77mr46qk2EKIsAu+RyJz4mdYhlQdJGnQMFoEan3OiCX2EJzmSSfPGAttXLIFlc3k
WGa4pmBHBpkwKgixyJJ9aTIL8TGzC6LaXPRZ6ODyrITBhQFYhgFhsnrmov/8MRzh
zY/Na/dPSwErtGTG5LmNcNf27njigF14vkpk9Da0x7IOr7ybK1Z78EvWKnnKG5wO
ZYNKv3/jIg7O10NGu+N4GkvbKNDMJeA4gjKWXPw6dooVUmISSZrm25ACvuqVdFf2
g9GxOcsJrL/coPvdbmd7ErChQiZmYC2E2Vb6k6csG+g7hVrkLhubb+TbHYw0Y71T
3qBPBbTgFqhBqFj8dwz/QtcxKCYdsdgL+D+mHcWw/noNSCJHceRLLmI+7U0K73w2
NXOIu07cYaz4ccwQWElSZjCsLYo0QMzpUP3z3isuzEfU5eqqCPh4MAfOjlgsx+li
YkodTpM+mHUZ5tvD1ikn0y9OJZ7AVZwJpnhnycEuyLIQbXT3AVynNAMIKP/M6A5k
RnDqP1Yh6Vf8H6dwRn4ai1+DmeHsF1CSTHJJu/BaVCqCwwz1L9CI0HWkrkNAoxx1
+45bCIqRiX3bQSaC6Ox+WtebPT38SBL+22hzGm+KX3AGWZdZ3DRaiqLz7X2CEaRL
qCU48/jf5u6pJGv5vIGTkrTKk9dIvl3UuIdQejfBwS4cV1L7WMfG02E25obyRUvp
GnMG6QsfUJ2tll0GoloQQqZrx8RNHGQ0TPWX3Tw73hkxLsHbFu9xhh3XmUF5oI3C
X3usJQsju31fzKDTpp1cIOq5E++oQQCSL+yX1CpNn+fDdqKVAiiLk4+U43/6Pur1
v6KQQ3jY4LekbO/w3SvBmQPLkV2jewV1cEsT93kjjbEMjfGqZ9SocITTQSZjtnoH
kNpIbjYBAHuSfV+HPb3XBr4ToKIsF6QQ24yU8xONcY4OBs5H1U4mukuZUBRzPVxw
wOShWHoxutItHyzmdNUZLjNRDG4fIAQ6M4lIWtGrm7TdtGsGg4WLRUAxDRl8KajC
CA7PCpRsRa6EbyM4Vs3mSiYdmsXpFn6mexR+NjFoz7vZ7qeX8EULMGRNNzFljnPW
fbLSAX7TcJiEJQ2kDBEqoCVZZLPpBjKfCVRp9DQ7ZdP/0aAuFaFyCkVg4czR0gCR
S3nSNccrJY/C1xgM269XzlPlYqSu8VD/Wtd6zmYZ/ymXZ2vzG4nrC3IiS2fg4djO
zUQ7PC2OOVgbHbc5UTqPEIcm+eiC4mh1yR2yRZ2LufgBJWXAwIWE8td/Y8+kzyCN
miZj2/Zveizy+2G0X9mTtRz7LChOXXiEpdOZ41DMKljgRqDHjBX5E6ndgMzBWeTV
NABTpvR7UcC/wJJAuX55BIFDOfDdzd8yFGrs6Qk5TJ8eVoppA2LRtsMFEOZ4Lcjv
Z2Nxq/Q82rbY8QVDBcrORsSJMi74ToBNUnw0lQIoddD7J74SLmL9IM+JD4AynXZE
0IxDayjkQxPPpRysHKaO3RNbKN4rbQPO4CMLRw/H0FmCkye2XLwC/B38NSr3Iz8a
IDMEYNI4VhvQD37js9zRIiLaEeNrUCsFHdNIC41o54Z9XVLkmErmkp10aFeOCxqO
yMfF/ls7raZu/+At0hqJj31oToGXFzviJfly3SnoXk8mbqGw+2HpBepbtJ5h8oue
n5TEszs44q4ZOEMoI2togKk1k6bAIzwYyGP00KzQ9I0mYamhprXLq8qt39hrnmVj
1A4Q8gel0c6py2vWgygaJrJ5KYEocQ4XG9eaA/LC5Y/AjbevibQUwRhksSTIFasK
Erm0XBwJwZsxIH2mt7iLXofoMW0OuRrhtsNDnQPVw14/jjphLGprhIu4FanG6iD9
Gnuvlfqs6TqsJTelNA9qA1HaqbYoz/XGmhXNGAjkBbAoQIQW7NgUmdJAmQh/wlXJ
Uz8uk/iU5EYKHEY4u8lfJdJuE6WdbAkP6c8V/zyaUi6QyPSdZL07TbxlfrwkNAj6
s3RlElXneNCjGILJ3h7V6qWd2dt21CS05Yngh0UIGdX+EouhAhpWX/PzxOf1YGbY
xRvtnv3DLIeRj9yDDFtoULQGzm/wFFDv6U795dmKDPzHIKN2Mg9EWSv7mXiDRmqg
vvRap40gLal/Xx+6W+rQI0BcnQvl8IAORg9NbY6dBNKhmF+gabQ3coG5F329g3jD
uYyTjwwL9CmQ2d8tUSYLFABRLcmEeZkDPcjaEmptRIVQxEtWMH3vF2HwhA/JqNgf
4BXjof5kf/fE4f3BT7XeZsbqR/2qgWoJnwgY9CQ0LggN0blnB1zRawdlUMCdcLhI
2TMqsTKywPDCK0zld15CmLIUV6yEpJTkOOU3AApOXHCYiN6tXNmjSxP8dgnK3KAh
5lDxbJs2WgEfx3ZM6pJDTHcviFHsbkyS+YEMqkTTkP9XUvn872F3d1prvgJP8ZC4
ME/GRrBEs1pHted/6ZhF+OhgfUdrkxYjDoLjFITxAZZJ9pFYlOh77Up69QZ5eo/K
iWTCEmIn17lBs7cRUa0n3EXg7EXMxDSpvfHles6Vnye1Jx4I3AIDhS+cip7G+Efc
3UwVBZK4yw9kvox7boHQg0zmFMWeXVg0gk2PGA10zbn4uOpZ+/hB9siop1bHaTrp
13OHxgxYO94a0Vb7emeRur/n1JksKPNpaZMoYmeOxrbhHxp0qP0FQ238zKmIyRKm
FWE4x3G0K5Ru4O6ly9/+NQCcFD3n1/0RvemcioQ6Q7Xj0F2ju3/Yi72JPOL//7Bn
JmW9C5kgfvsRUx1V44HfNEd3DjSQV1B0SqgiurkEdpdv6w3em3zGrBoJaqAGEpM9
Mne0jv6UymSS1leG1dJGmC/IL0ksD3Qg0r4E0ny0W4YW9QYRJ3ym2fe35wQ8WEtO
Jlq+BHYRr6vrZsnGIgfF1CN44VmO5PwWYW+ayIyhzpaIt76puPnUQnLIkp/4B9sB
eq7oy0RuogXgvNbv0zl7w+3JpJWc554Vx+4EemLYXy7b8IgOIctho/BKoVmYOYV2
/FK0ebXc6+AKUvwgvhLiSNWZvuZACL24/Zwsz1ZZ5RuMmSm3yM2E055TM3BTl88+
EkDwKtn4VnsTphdrZqnSTbqLZBnRzjVoHOXxif1xu3KArA3zlx4z+QlQxYmnnqbG
Q55c9umfqyKGaiBGkuNWPYevVErLi8sn/bWLB3BaErhj6+w64icDNGW6cPtAQe/1
pODyXScXSBBFvbvA2RdRVQKGTolUFGNh3omnH10uD8zWIEMhvqmg/TGLraoDEf9C
pjFHprMXRJ6jCa5xkmw+j4dsfTsC2iVEcQD4lbWgtTcOyFtE8DxJlTiUNWPEobOi
d71WH3MHz3i2UbBN2l1z6G1a42y4S6oaFLqXGGrkGGKA1cLMjm0fTFS5tA2qvIol
9jFTW19epzOdbegiLaHn1WBjj2eA887gec36qt8XCv2ZjuEsbCJCUlh6oTiBjUyV
c9QLF0dSqBqZ+zTQQzUSHrOIuiDV4Inw20ZL+6b5XdSeFHUPGMh5w8qXScBZsh/+
JsP+tUd0+v6HQSWG/UQxins8ePtpmsQSlQJM+gZcETVvqQTCK9iRA7I+4rTPAAc6
/VZPtMnSBVA40LkYjHqxnlquBlSKUo/KheBY89NbexnQvQovpzL6z2N9Jj35wYjX
fkIqGFMIWstPYLi4laSGxrCUMm29KEHAmGvN/Oq6Ro0JgK2rwlphkG+PDpSyDOKc
Mj0Ff9Ex4kdxapr2LV+aKJGTcF1XAtLivQ/gTgRcdXdmDc78gwTe8ujbmtEjmBqt
rOV7s+uIdJJ+mb+WTK+KmRtAr1FSnnkR+LxzG2n67X096ncdmzonnfRqudFBRKxl
rg0KjBFLRAQcPw/ZRYE2Ioy1e/JEpvpxkFCnwppxcE1hBP5ym9M/n44yTHhb5I+M
5RSJB2SP08f7NNESjn0eJm4aH7XyQd+AmVEVHOdCq80pOnqTane7Z07+aEQ0X5GY
0H5DcSu7OYw57hsyVbNhwxwS6gn5Bhkdzi87h22fLYU65hT9NevCjrPGHhIeT0B7
de4lSBr23I25cWb5ccZn8T/Djc2oEEuwCNOkL7wpHWoCpHK/H56RASePz58ID+Ey
HppogM3anZTrzDfN0qIjkjvHLqQBddvUh64LKeP8a+oJD4qrmUkM6WJkePvCQdg+
tSPO3toFgbQUuBxiWIFiecbNJD+0gMicPJzX4xDhD0Mo7JYA4iTmzUJh6OtD0z7u
GIquD9RHW5hNmBuKEhpH+XUYKkbMFxo/NDgjUfuW6cxOB0H2WkAPFcE4tNR/9Gma
YhxywHDc+ol41TpWT8OWs/c9/wE7bKbiadqa7qE9pccn5eizJvOLGYx+N4NCm+NG
FcloQbmhTOtVv6PPsjNN6G/9vkBy8mlrSbooU6UlKKwUjZCboEErGuFNWiur0u8i
tJfLSr7CCYNP1jVLUvuRHHTnMTeUS8A3E+CUH31Zb3dcGzH3mjE6sj9fXkph4/G/
UbfeXl67vnrDITWUzVwvPWS6Jdk4qsGHI6Kd2ceU+ICuWTkrgReA0UTonjCvVoBR
xeq39Qz8wvgATiu0czJ1KT4cJD+uu6M/YaTk/bWSa2BdmHIN6NvN3jhrHMCXfGBx
eH0VZzk+v4fqQDCHsk7LFfGxtfW+iD3e/v4cZo/Ro3W9ezi6jmXzAmWfS+MPyfTA
NmtS3XAdDA5YL5pK+K9oznW5owKJEBA46QAAmXg/hjeUKw9XOQRnaVkRWY+lMqM9
x1YMJr4C7muinYzwWAkmrvSI+tS3wBszA0t9bdl9TM27LxkSn4JvCzDFI8hB2CSz
2UNRBtGpvJdGqFXLaFugydd1NmGaBIoK65TWgtqIZ99+6w/qigW/0KEacelFX4hA
xu3i9cUCubm2isnrXZfQB1nmwZPYBvf60bnrZG5xMSQw00F8YVrc8R8iv9vQlIm6
QKFCyF7TFyY+4sirX9WbfiJJHTt2EVRSm21PIII8SmUQFFky6DNniSGIbChcSdSa
g5nNjxtB9JI530jFyfjBA4D6js2wUucNg1AB6jsqBuPoD7JmrxE26TTZ8AtK6/4H
Q3FoBgDaSFASKV3dilYvWcUE0N9JvxMOxMUWXmcxuTau8tdDnYOgFcGgswOBaSIK
ukn43/27fDhGd41LDffpM0y+87Z6aJvr82vR2MBlJxvUI5VG4wRbNXbxYDM53GEO
ONegbaK3892/YzeUv1AYrzYvxu5KUSvAtAWBEwqT1DVnbI5O0O8EVuVdhqWzIqJQ
37agJrDw9T8yKQ1hU3+lgz0n5xDfqzifFaFRN3FomhJ/PKWwiBFOzLkyQlpTBNzc
66+5/jWRKMXpKGvNcrPvS108pv3HbFuC2zmO5BQvu5QSpMvoTr5Z8FN4eOB3zlr5
r3x+WsdHgGwn6pNxJNpnshurV8fY0qPQv91noODuYmjJExvu8G062YBnJnaC2zq+
y6qvvNcxdeTssM4aiZpEaXVoeYS6WrXXO93WknZTwf9/fwXJMPmWadN1XisYAtDE
/shZNGhNNrB6RcSOkyfj6TPy4ISHKLnN0Ucp6LpKWYA48GhbtP3tbmT0imWn1BvK
DA0iAGhPCueehdt5MYokry3+Ifs0PmF/3r/8cYH4jvWBehOKz5K7Hro8MFVxaE0x
xsrZ2JK9DyI9Ff72gxbatDBINo5/j5AuectkeEK4FOg=
//pragma protect end_data_block
//pragma protect digest_block
+a/N625IFVhtNboxbplNiLA6L1s=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
1lNYmmipQlGbs1qqEvFl+WGecqAnnCDlOKWWm/myUkZSz0vLPPRKanWNJxyNydLD
Me83UsFYhMJSqVz1HhO+UMapwhXybuqH+lTrMs3u+eYp/9LahX30a9zlZesU6noQ
THHmfVmNJfxGvTtLgNg/DsC91tETyk+HtOVSLQVxM6TgmIFKj0osNg==
//pragma protect end_key_block
//pragma protect digest_block
KxIMrvNyVqCimX5DlKP9v0rqKxI=
//pragma protect end_digest_block
//pragma protect data_block
0Xo+SWtXCdLKvpfvY9FQk444GIhLo9CyAxdEd8aABx0VMbJpXcOTK8l5152JYPy1
rqSl+JITwmKQ3FUtCX57C9uJa3vM11sGirY1zcOPXRjJ9dW+L6FNBwgx5U1xDO6X
aVTVQdu4Kw2fgFzevm25a/Lyx1MinIxdFv+g6RaSF98BtBqeW3fQEU0UElVGaFjT
DqhdzwofUmmoCVit6rtaqa+apsp2kB8ztFqdhjCRjOIra/ilf/RLhsQAzaS/QBDD
UnlUckwv0M+2xG02UvcWMcVxEG1s+BrLbXXalhuY/pW5Hj5m+TnRgX0FW3UMx9zx
UHogQaMdcv81eY2IcDcjCH/Wtmor42xHaFQ5KOx4UZHmySgaftVJTAVyg8NdqmpV
2Gr6polJ+ndpM24+ltEWsuwpOLQwrvnnX7ycQu/5AncFSYGOAJXVvIUaUT3W1/Ck
tYPwNHi3xQRijewdrQxZAKMZLTXaFAAmdbgd8jlk8s5UFtac9QlhYXd4B6+M9sJP
kvmx/KzChzSLLX5HFU2WL6tbTKefiS+VST4MnxzfFtuVnvVzWIOIqPyrN0GcOXep
pYSb3s9L+fWHpfY5gO8ef7FhWNzZHkPGIvMQhAtzTTTq+P938s3DZRrUwPQrhWP6
sGIFYRjwG5IWkRPYzwYEG+cPblUufGlxX6bQLiQ+H7EnW7EsUuZALj1o0hi0rNgP
Re2iNcWxAvBTb2SOWnzogJWdsDloOzuxRelC511IMKr5N0KKigmq+E+5e1T44YLA
8j0JQAZ0q3+Z8YMRsDTupzhYBFlz/vuAc2/e6jAB8mFK8ltWKd6AuLhguSZ6ktej
dL7gL4nmOgYtUeMalbOXqVbrDCkE9/rjruHtswdftfy/wlGosf7VF/Xurdr1S8kN
5q1GZe9wZG3feUBa9NfrbjpIAKW58vHqzM7VlxqpqgocxDE2n2Yw/U8k0euub9Nc
yV5G9LH71UZYgnq3+UuONdWlaDk03nvH1BFsTe3bh6Y=
//pragma protect end_data_block
//pragma protect digest_block
c/6AuGYjJNYouOShc9/zgjw9b00=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_vip_protect      
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
G+w4y+4NAw01W6K7BoBg1wlS48HTpSX36u8UVMVtR+JZKI50mnfwNI1hqVi8KhJb
PqKxE6QU4EhsBw2uEMhJXtecUe6MEJL7I80XneYK67OH24WOX6N+C4CCtFyp8V2W
uAQrKLcN9p1miLIbe3RaN4fXvbrQKX95JRotKhrRzttFEsB8CpmiWg==
//pragma protect end_key_block
//pragma protect digest_block
rsOHCX8/kMyw1Cdkxzq2P7aqKY4=
//pragma protect end_digest_block
//pragma protect data_block
53YzcMBhDXbmiLETAOGxQrnoYjLll6PUa+ceWTQ6ZLfhcgGhFb19kTVVCzbvyOM0
MUvT7ZW6bMnNgD7A5EF7r9kWNJ4fTjWQlJcIWwqsy/nTZ8+FFJRseeg5cjJow3G/
BehoFN4gaj5FdbXrlYMMQJJpRrmDq3Xep2BvmwKlGMGVJEDdE7DW5m5AmPlIZdYQ
mexP4XWDh0XsBMcEa83hWOBLI+y9/Zs5ua/3vO3tlKNUNsaAicmeB/YlYKWfmYX5
qrwdEo21IhDlTVJKQ3JrgR5OtY2870t6zvgeXkVWs2e59EDGzgaC9KCBTB/xzZol
ZrLeAE8UV4uxHfiEQGij3zahejuu2jQuU8ZLZ8fnkNtZK0gXxuVsBgUwz8v5PYR0
ADotaJvbkFcqzze9JHil7nTg47/rBUm0DJbKw/CGmNyXsXia6V8jKksOLcfsyK1w
JR18tEOreBe4gwtSztvEcGQRBGv4qAYTrsPPkA072Ip/mdjpV+KKlelcEsNcHbgL
51hDIOTJtrWHlzKjDx5+P3P+5mjXV2lfwOkMeIa26VFn0Wztm6PozCa3mjOB4oRg
8v5JvDGve2ebeUpyap84/eYV1S7QaQqd0vDATHU5qNO9zT7oAT4/sBPi4GFzKXTq
FllEZykB6+zJzRjyGfA226RwGF8VqxZ3G8sd8Y8O1bnI9W7YXoXFGScH8eGXbupw
wBwTuPuRdd4YzFLEaDXdE0Q8pIL2VmEejCYDgFkoFahGYzESdHR1G1/xf1n6GVZw
WrITnHy5v2ffCph09k1VvhqTnfnPbhYVdAL7rZsTotpYqo7dHOAbV7D6BqyOkYPu
kUxPegAwmRMXAvE6HZHyvwjkXXzIFk9qi3JBLV64zJ+ho3thK0rjj9nXa6GUmygO
RnJekvWxPtV3XXaEvqaTDrIGhABgRbqlX2wYFBq25r/sFhuT3EUHMrOXApWIXtAe
sPaKUwNQrss7hYa5RARebWKs0hMCPaSYNr6myrqybbSgh7OAsWnPtqT/Dm/4bwtM
jLFSLcf8fqs2QqjRViFp6RzUaPfezHb3tO5N1LAAcXZbkTbgyljwNFBP520TiAdH
yZER3vdlMW0j8R2zaNM688dI/hbgXD0cAGeLpNIkDyU=
//pragma protect end_data_block
//pragma protect digest_block
jHBLUx0ftSeL/B/eRXaTD8HBULg=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Jzny7P8MGUWo4Kzt8ukhAXeI1FXjDfGzHRYEVYvey77YsDhs/iuZKBoZpBr3/Gol
eLa8jlDWhEPklbqV5zyA1AY+NtkzWOyaeZorptKz0PiPekX7hpPFxSBZKhvUP5nA
N/UpbYw96oNNmr4qI9ShumJVXr88HI8NNnGJoaat9ZyKtPKhHHqAFg==
//pragma protect end_key_block
//pragma protect digest_block
ISgIuP1AANS4M5Vtsir010jSsKU=
//pragma protect end_digest_block
//pragma protect data_block
LWlDs5aELXBfk/4vb9xVWRZALJoAncF6QxWG7f/R4fpbnKJt/3YxHJ+majfQ3epj
KF2Sph3BApVpxZDEvA91N7EJTkKznPtISxnxM6yc3zqsbotGQeQtmLVv1rBz+e3P
3yBnBaE9KA2ZLdUQv0beO/V9OlnvENedoOPoAuVdu2a3M4CvsuP6V/Je82OC2Wgd
raf+w3oF1UVDjATmoUPEibQ05Qc0oDOb3RUU61cPRAMt8DOqbzkdrf5D8rqpXyfN
yT9yaBDLVasQQ01Ron4lKLrh1sAP0e5rmHEwI8gdD1EmHHhHWofxN0Bm2DedLyFY
aigwGCRInTyD5gYVwEUI0kEePAbSx2vQVGQSj5RqZaEhUzDJnRprvWqfYLYw1sHD
BqGxhBczMISic1QA+nYR6PA/IOhmbhrRvbPLbS5nd1Tnt4Lb4wkZ9UPT2X5gbEfj
8JeVFCVjJEGfE19e9PkCAHmNYFAmisbJHxDNc+S2BSx0b3J+Ebq7VU0fbchRm8LO
i3xDYfuZrjc/WhA6mgOHeg6aZdeXIsX8dW6h6l5lohxrEbNj1htvtG8cLmOuF67d
OfBfLbRQRJ2kaPvNZSCfCmtFQNUadHgqzF2Qj6vWmaId+vzezMQfCAbigQbG4Y+s
CBsClabEWd4grrUPkeaIFoFCG24bR1OCPaaX4whCfGfcnZwW9B0CxFjldTa05vmM
LnrromTMif0hDT37iKyREln7BGYtFzcSXRhdPoiEwrObHUuQbUOSkCb4yQ5MAY4q
c0fxcxhTRTNlyOyGiHV9btsi0muNe3rzsfkviu4vMpFrQBsFa5RNHg7efSitAms6
/MGcDsxNwZHQ5IPzEMe9oNYpj7uCJRD7IeqeUKClQF9xhdimvLAhxtChGdZhAAWX
IA2FBhQIEO4lNvz3GvgCtvO7vk+84nB6WO5Kx7yeHUbHdhldLnWLZH8dZOO3BM15
J5EjvVXjcb9wo+UlkjIUtH2zXajWCz/9NK/4RVtAK6BTDsm/1vDsphb82Nwc0v3T

//pragma protect end_data_block
//pragma protect digest_block
sSvNyPZxPxvLdDvIP947HhuziDY=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
h+zh7QyrJLoE/Y7YM4tjz6EIG8gnBAkpYW/fkB3K4oyJ24saeRYp9CkMOxdDqO/J
Xbo5oocifDRqdM2wl9Gj5MQwlrdYvs95zaghGgA97FioPydRx/V6DKHGgV8fmyeV
e3e5Fg4HqFMwkUjP2j06sqjA3MGto5mBkHrv6kHian6iHlZe0tv/IQ==
//pragma protect end_key_block
//pragma protect digest_block
0CY82M/TXUg9+WSpog4MdS9bKYc=
//pragma protect end_digest_block
//pragma protect data_block
vpfOQWa/5hI2BB0Z/VCu6tAaDBbhEbBP18thoEExyvpzZJmo5I3dngDDaQlbZe4p
EB9Simx0nrxTK7bI3usekmUSNOb+R6rHkl3k/fMAbJICqTkQWibqgbX4cWt5Niz/
Bkhb7uOkFZ5QKk9cZfmobmRQcYGBcnI4y7x7vgtIrA7zx38jIp+QpKsNhHUZrMvj
yGXG5sagkk//eINbRChnAiYxwlBhic+55mwWV15J7906jEIh0xCdhD7EwuXFMZs4
SG6MAaaIMJDvKiZQVgUjfw9zM4VG246Pn6svfHYDsEKcafL4AJhxP1q7kmoxzDQb
SS3aDlNqmuOyYjo4Vw3DPrfIpXST5Mdseh+00BVij33urtVIHhMFLeNYHgolUSQh
g5nmqjw2Juu0SdjSADUaK5eSRPMaxE+ee9pPVfJaqbPH/3T2smlhFMB/0TSin+Pm
xcto0Aiad4Jc3KScxUwVAwmu2Mv+IqDLjR2cgETuFDcTKTwh8GnuMehHX1yoc7N1
XokAU7eNWFsOrAt5GaUXhhTRvHn4TeRWPW+9T0Pp1xz4UvLAe724XUXDsNHzPdY5
JPF44ZIw6zAVVfz/YVB9x2dnlJrsAWBeKlvy8tZ/ake8zRenUvQC3cCsY0czg1wA
j212JBjkTNvivWaSuu7sMZJpHd2F9rakeJGaCCf0GMnz+yf5hoPb2r6E4A+MVdsH
YvP/fvcK7gRJrka58B/ShpFKGq3gkN3WBkhm4RH/0VRRfxtxJXvbECgaF0La7tU2
QEynD0W/t+aBp8gNOlr1SIA+rphK9rJKDEDxLoTiMuONvrElHrsUO8pPoayw2DQJ
57m24e1ju+SjZ2zmkWDQGycnie3xE0SUsf239B9yoSfHRMB3IlrFi7ax4edj2SW4
ol9/YR07dU6k/wGfjNRCyjmZ6tzajrH6qDdY+gdHnt5X0lb/mMmJcR6wTtDhCQIg
i9MJODWLdrNPYRz4M5astjsdryPI/cnpJnXaSPImDJrfB0m2Xq/x0oS/lbu4y87s
rQ3Hxg6lJQ4pEdPx1IUAlX8IF4HocrlZJHauAKPgD9oM106pwpmg62MUeL6WIB7S
HbFQSscBT2cxWi3SJAElY2Kry8qXXHwCQZYky4BsBvxtWSSVnbcZYN0X3lLwrC+m
VitJQhkRpyRpQphbYJcPE8A87OsUGtpc4XC0Ug1SKLgWVY11Px3KtxdjfKos+pgq
ArZ7rFZq2oVcO/BkQpzqYNSwfoMRlHZazq76R7EaKppZ0erAY88LldcpoUuMzx1L
gcyRy+SYdQTLmdyZpYytNhEFt7I2QVQwYE2VNspYsPsZ5QSm1/3ThGBPF5Cmq2x1
M03dh12yXNrGEtWCKvwmZTRc8wmQPGPsGc9XENbb/+mmWPdkRAZBrIG0voqZPXN3
58fiP971R4LRCK+wzzX3SaWPl3qQJUjtEo5HpttIZOv0nfBxGkrNzM3Fdk4agFV6
DUVzm8VpaoGvZro65eq1crLOhXUSIsFlzv0jwVUC/JxQ41rTukV01G9j/W5Ba0H9
Hl271dDCA+O4WyBV/FpUYZCJxISq2iMYb7PmahLb8huud6S9RquReWTBR+gEFL4v
qRuHtrvol60PQlRK0PrDqD2Oa1d2lZL6ZQs/Q2EgEHJziu6sMpk34mg8LEtkjkAC
wxgLpMfFQk+1cwSvQWkMEBPOaipWP/KTfncQ7vTacBxIa+eNH6St3ENDkDG+iZPI
1osVaahdYAcxYUzQw1DjtipMAP3Fz6n5hJnXf+gQGr4B1XT9Bft9KULwuGSqNJ09
o7sW1VfBcVTd9/fI2KXKAJYvkUnLo6GuNqfS5VeQwv+UiAfmouo80QldatuUGWSQ
7ndQj7f5GtXQT1PbOosKdRtImgDKjLD+Hox08AyySJnKwhKoe2Wl++jbZaBFL6K7
Dh/dwVTVzLfpN2FqoMRWuCotKOtCpMsActAbPpVgIeDd2xJLFsRoTasgRaGYeJXa
2f3zkqRhnuG1fXy6ZJ1qz37xOtZOlrydD/kGM3MAMXbzSnCvQtjw57WZmegFA7cC
Z3asAiX5XhIV1VNFuNvicDkPSsUpCpeX1xwPRYtA8f48FT7gxL5ULE3uqPFg58OZ
6eGmVmZPtou4SByoow8XosUUkFSG//s5h8HOx1Zsh8j/KED8h9ABPgx2TGObU+QV
8Yzm6BPu4t/7FmUadst8wVPsKo54Ck8w1vAJ0G4BE0wr0FOTi3QdrW1vK7NNdpU1
ZqsZeKh6IgcmgG35ploVN97tcaMlytii+mZq46VwlPyBJVz8L1PwYl/0paA+Zg9V
yA9hh6HrKjb2smQOaIBB7BgvYtDLSskdJKHTf4z6XdSn7BmbH3FLSpcFfch3Y1Nw
1bGOJlZKh6oLkU5/jQYBoiXwmeGAvJd6BchRhoAyu+BsQ9ZMGEDNHRpAPTOYxDj1
rx4QUZIKOSkUI2oFv/VPheAr7+xlSgKZAPprlDx5geLfSUt8PJ5LSKuvSeU8xDLM
BfYSCIFI+60NdecV6w9lOFsmcOy/TmyRq+yldJcIPsGbT9EHTbTj9urhz5vN7hZu
qF58gWafdpL+UG2cj0ueoZHSa3kAEUIYmYfWiwpv1RmU5hEOFC+hNBlOBPbvCRaD
DXVwsmwqzczk7VRo1GU1AvU2ugPR6LuXS0csVaVqkwTCVCF0DUaNK+tHIz4zhaFu
NN5P6ibHt+7jxvU1vp2x3Np9lSOeHP4PqIU4ZdTyc8McYy549Prt+taN0MZoGHMP
Sx2zzEPMNi2GeCicabbodUGHkCLRdw3u4TcX7u7MctWurPsAwaUHZm0N1AwFanTc
70ocisAYPJjRo3h5ekRB8CF62hXI2KORMpi4O30xfJZyNz84i1PxadogWriNeGIg
itSa5qcY0s7nkUYjLfX/SqEcEeFHH1Y8bOq/EkY6fEwjGIOt6Yz+10ElIXR8Ev5r
iQHbDI2P1lim+tRMpD5myPrun4T8rZ5ksE9qPEC2/0E5IueNIUfq45McHy8qOUxY
r1EhigXXpy2sGwu6b5+DoiDVFa0h3OboAhJB+otW/DdIk6fgYX874eTSo0+dwqF2
qIkC7MVy3rYsl+9I50MvH3XCwwJfqZa6lbJjHYKIYjQKQiEkgOUnL3gaAp8lZKI/
enGgE/C2y3ZI4TmAwW1hLJZKle19+15JigjAhcVC7LZJUdiHR9eWx/79n7ertFNv
Vc4TBIMfnmksPvte6ieUrtSi12ZhVhRl5j35IZIuYg5nc0x9sUxNNKCBABNTZylU
Nw0zDXgUGslxQzN0m7eBqh/UIEaPMMdWIUFiwlXZ6V98tqcAHIvvmrjZYW8rLyYs
Z6qpTgesRCaHVzteEf00pe5xdVj363bBHscRn/jZogL2dmF7LpJVnAM9bx8vXza7
xU8RdO3WMaN2kxl4a+KOrN8w3Ymfy4NLgv2dDgD39pswXX87fgbQp8dnUPh0sR6H
muocXxksrlkSJW9IC0Vx/RJaeVBGL3qeWEfT/pqM+7nixxfFlzsa3CdJPDvblfLh
du/xmFVSQYmILDu3ebEdSFaXCaeoVuiRW8xV3QHp1gRmcs8n2rtiT/46xBuRNBJk
3GlZEzkNUagsKA9Hc2XyrX9abUBTHAKF4VhH0Wbgmnges7cl1QWrLOjgJ21N9CXA
pDvEjGxIbKsyWi61P9HXwfPTAU8atZaauuhN7JnenEIq2ILvLWDmKsgvIWvNh1bU
DrmadYCpaC3FgtiR7yJWa9QxGR/nocObfMKoHSfUd5D78ka5StHTvqw/gC5kWUfp
KT9EQBwcf5gl2g9UIDVB9mwiAKSqgs/v+Sd0o68SJwayLjaMrr4j/CmOA0DLCOU2
rG91hgkMo8xQjtnQWeK8IgqQo5UTb3/B+llX+/QfJH/928vcWZyeL4C/oLR2Rxt5
84FzeN1J875zkIBEMIZWmFZOiJTH6ehOUP12SmSX8idSyz3c6t1gweYD64u+Ha3y
SB0fJ5lxRoHPLHLqBMvi/ChDc8Y2R5t4GqXUaciYgmjeuz6Yp1AKDM3u0PqleNIV
aDQXgfTPqvgp26OE7gvC+mMendk8VSHT93jf1TUhOxAzq0UHkO6eNHNf8uaHoj6z
3t6dMOa3SExMgEd+jsmL5bjZeUtz5utXBNKApujcVesBZL89a0FbnpwX6zz8xSXu
EZ1dRwpvo1ykEeutXvxGN0n4iWkyUHAYe+dpdiAfKgSzVojp9eNBGe3oOhp/EZ6D
kGdKGF7KRlAY9jaKMZ/wA2BMO4x7+CXkVPoci/kAO1CxiBdJei2Rzg5k8HUZAih4
u5pZYqXcwN+Vd1aOPszKAnloQ6H5BN6LEzIexSLX+HHSB2q2mfSVEml4/AFl+U3R
OaQI7L03X8+iktu4vLXoEK8f9WNZnRsfEjSVxENyLyPCEpuIHRKLs6xp4PELO4JM
usK9hoyutTcDEycVE+qVX5n049CK/fWYSTsTqiNerne4LuWnIA9zaFnVaoV+Vp6E
Sa0t+bvAgtzoDJLLS7v+ynZ3/5K7zbN7oPYdKiFUi0Azy4Aix3aram8rSMEdkzB4
wVaCHi3RAvna3xrCz8YHB/oMLZrXyv3nwPbSfjNBX5cErswahBe/SD0Ny4YUrbWM
Cjjgzh3BHwLCUh7VBMwcJ6ACYtQxajIeBxRu6HEjbOflpaOgIIuXU7juRsU5QF3q
OlhjD8cuxkDg9ewrv1UPAKoyfQivdwpPYjYG+Hmd1HLYxmWe3+0DI6+7yQHdyr4l
oF3XvjtEYY0jY+bVR3DGGc1B82yR3sfhSY+HeM4OHiFOTJqZlhIBXWA7aMLRn+j5
GDFqDD0V0pvaX5688tGDVRtc5sIwIOdTTTirIvJrZCAO0CLPHGbKvzljuxNJM8Am
D6Kswx5BqRKgM1jcchLX9qMDhzNBjtPSDhpAaHmx3cnVET3Zo4dN+kNUDp7H+SKc
CMDUk2HKqSpx6LAsx5eSM3rgS05ZJUlGtv952VKLYw1q1HQUhmU6uaI5QeuseVG4
/lVztW1/nz0gt2R1yiB9AWVJabnOxZ8seKkPf2kPmoDAsvF++Sf9HtPBirT97GTX
z0Zqrw0hOHMfnjxJC7Lj4Syh30HAszsubL951zT2tx2zse8U027ep06TxmaGsuvY
gK6oxRzZq3OwX25l9Gg9jL7SfNmQM2tsiecl/vpiCoHo9E+zFNsmkuvOZQ4xJSyx
UHBWcP99hnX5GFFOLWxXlcI79z9s4Le3yXTRr8aWyaWBRovVo9C066wKf6tAlIre
UxXd1Wcr04C4bugBZZ+lz4xNBdEfAJnti11+fDJmMTBld5zd4td/quT3JgZiMifk
VYnXudBx3uVa31drXvTsdKqXY2SeDcjPy8ypV3uCUqf4gzJxrW/6g8hf+rv9HxYQ
ZOlZSx9A+z65aeNV89sx7DF5C0m7NTl6EhNIVA3oOgEFGnW7LWvGXubG7k4kFZFO
DcOYLEIhA45EBdiC4wJeKPGgo0TwdeIvtiNb/azPuXP8LCEoUSsBxycll85HYM2v
RtwXKiTgY8KskJIefBJpM5PfqpPYXRrDTtvZSJt+R/9qMLkIwFaDj890a7JeojGA
/9iKTwJ4NnyaW0Rr+LFHoP04mGI7DQQpJKBXPXRqRzhybHPGQdbrbiPwQEBHGayZ
Pglg/cQd6TKJyT6WWJ0FrTWZeMrAaTns7hba4PoeG326j1wbqqGkvmcZL8AGs7qB
MfUMTGwd5u2DgKMSTTCUDEMbm4PAXJePMHcCIsEZGmn8hFwsrg0qE3MzFkQFy5rH
s9lERuNsdjp/Vr2kDMQePvegKKP8HcpRrEBCXepbvN1m8e0W6DT9tAvls0O4Ez/L
JQe0LzNC3BsuXTmTHU5svlf7fPxn0VpN49W38vMCoHdkqefv5J8hlWcfAjy8WXVE
mMBnYTwraOWTvr3Jb/2YT6c84fJtY59WZ5sCtMYoAEVkO4u3FnXeIEPcKLG/mCvg
txxUTSd4vrCQpOTwNyPhIBilRnN5/pQb1/zGbCQ0QLwj56TOeF8HVtFvVwWiObD2
EZNd9ba07ikmpGrf/S6Z2OQ0hS/RWg0Fv7w0M7m8BuHE3kZc7KEyyNXTO7SL0mBm
yoA1slL4hsMWypiqUd481t8TjQ5pAv3gxpNElvKvaS/S+/7W/kMZuaN8zPJIbjAU
u+8gSfjuMg6CWg6OBTQJHH11p+noTASAtXhKB9FOIXVNiyeBEO9K2P1mhPCJejPe
YXVotCxNpHSZA9DwPCGjSm2ayxeMJjZjTZIgTy8njW6rKn3TSjIqoqbQ/45Mn8q6
VbZCO7F+4AKga/AMFUPr3mXpceWMijGvODHAn3mLTsYDn56HIIQXpytJgL/MtI6y
9IVX82qOWt7lMwlOQhf/KTHkkbkxPU1vx4rFELfRveCvtPRW1mu88ds4bMFsP95w
bPw2FQL1C3L6sv4oSyN5llm0YVVAs1YoBE9oqPHaOXp9/xs8BSZhIgP4tbPaJRj6
6lkpHBHvn9/V3SvhJ3E8DuPX2moABTpB4w6kajBy6MRFeborWoTdON8p6c3XZlp4
pVZFS7MZN0NK37NSEmgYO3uQzF2VXVp+T6aOTLIKKH6ZPyd0735rN2S3y6P0LVtW
NvjV1ldzA19ufzu5WblFNXBU/Cv1014xj/hIiBKD/OiMvS0dLMgUTGoJSwWdOexF
QEmPlDkCmSWxgMgK6je9cwks8YczG4NG8eubY4qRkoLGiA+5SxGM05aKC3f8L2Na
i9/olrAImwKuxLn/XWEU/DtmOPV83N6FF5sK9YdUpu2DSDYK9pjzo0umARekWxd9
mqX0GTtIrKsMLrPPdD1TUdHJY0z4RXdVjQevlTOsRqep9osFGhW9B391AjaHElm9
sPPCm3NCWMDNgLF8Lg47BieAtioHgBOyBorftZfy3osfrwC6D6EAnKMJbBP/D8sR
/4LlhI3mDISLHNF+KdWa0So4JQhgcSsCd56gEAmH1ehqhT+yAOb3QaLOxhhtMflK
w+m2xC/99n/fD7S4pYCvSBxwEs3jEP0s2ma41SUnwMqIe1e1/7KxKLYYZxaFnMR8
n60D5ygYunyFQfuokxQBqQdzXjh/S/MfRWDqNiMCXAqxb4B+SJI04FDT3kEGRWj+
yuWZTp0ww3LEHSsFk1/PxwZ65orPie61VQQXA/qKIZwMbz5gs2pFwKIrAZXzstGB
rYIyeZ8mCDOuDT+HA8Q2rjCTNAFEFErc+eKd9CxxgIGs2uvZoNEpi9TQXWPWoyYf
c9QUXYaENsn6YU2fYexCLdvEdRnKsXdYWgbfdRmjIdyJngh2umMpvZqHQS1BiKtT
xANqeUfuUMBN9lPXZiYFf84byf1EmCZI/wvLmhVCTmL3BmsgLs78Jiq/I91LlxOT
vmsn+Tf5uFe+pRYN/lLK9R9JOlXhzcg8pjGr7QW1bZwuBDQSALWB1W71oPiKAs1Q
RcoIc7yEvVFs9DB/Me30N7CjyUlHhSklGgniPPX8AMzUaCcsg2ElejoLXkNkuAq/
/DdgVPQMn8N3m3Zz4B4qpVh+4HMIq3C8vP4zcBwnRI4wEFzD7bKxN+DinLMzjhTn
LT+X7W7g159+oC+e/8vjQmeWTU1tTQae4N1t8PM/zAxrnCPInOS4zpJqkCQRcAfV
qwQjyluGptsfMvLyl4NqCZT57Ho1HRQWmefC2ylgOIT/MsHH1yurQ66RAyb6p9Qv
Srv7H49uHEFcFbgqRkxNLhgysIGGzkaHFRW8fX/B5UVRDWoENtWKYYleDzwPs2XQ
GLaWAfj0f9PkEthGH4APhgCCyLRGUR5fg1MTmnvYwMsewGjFr7MO9HWnBM9w1Y+p
ff+54xSvMH9fd04+lYEQct5scOkRkO9Y07/G7oXWJcp42UGns3WNiGGC6Nuvtgp4
+8ninig3iRGbOwLv5psMyHMSyxr8kvsnSbp5yrVAyN2jvOBreNq/CdS3kZ0tb5S9
eIivCW3H5tluduXPgQuoKq/74mrGyXpgP4BdIAUSdMnvG4gbfl8xF9G9SsLGBDHy
JaMlxNOaR4ULBOPpL307j06A8mlbOdzGMB1w4YQ6khFD0uA4Q1gCzey+vKIc6CIO
oqViSUfVwu0l5xGxLOEALkSZs1+OANcXqq5ape3r4NCSmb/8EzCFALDlyH41N2Fx
junk+Cn9JINwnPD+J79mfV+JDKgwuS2h1ZNqNZ3JlpF+k670/SR2eiIi5caVO+mo
5NwCNDZNyLJejDCxmTD9BabgLVstlOV+hSkaF7ChXz8R4Il3HDhMSUCY5FIwAuNG
2x3WvROP84xfe0wf8di9huldgwey56Cy9n/EDWsCuRo6UcoQAyScb0Z6VP+hUIbF
ov4HZGGPWYyzAe3Xj7cbo5b2mU0qqwcJ5bqP8F0HFOJzOv5ou3y4lcMWrz38Ekun
lJPL5ckxznpZrkPWXUxXPIkejgfi5Hgxj5DD4jszXdMSnjeXWgX5aw73RvEDCusb
Q92MgBmrN8eZwfDNz9rv9qH1D4Vk/YFGb9AIydoBNwUEcNNrkD6s2ZDf5qyagZqD
modIi0we+agayDPPWAIEGE19D8BZKVJoATQ3uQkQO0I5av5fUn5c2bIRzo+U06G/
+NVrf0LSVAUCFUvwpyy3LKvdNedceMYPLQacQl6VDGvw5PiTe81C5psXtemF1HqU
VDUW7YtHIxmWh97+FLfQSDXcxPmZbp7gFcn/jSNQZ2rn5m+ypaSdL6TFQI2x9Br8
B8nCbA/X8/WhBiQ2k1DyuOcpXahQdriE6j2Bh/oDPGkiAw3Hn/AaNc6xNeh5aDVN
C1WqvpdlGnWmU8saO2Ww0l6u3h83bNFoJrW0PwcUT9OAEgPzRUkYGIThtwCbppIS
PY6ghP1UunSIv1TItjlB9jXK7YvQUzLlo8HdngJAHCOuWgwhYGw6ecmXoUg3z6id
jLsFAvDEn3dJK+s6EB0adzOy1knLg47fvtUjnVG75xvVubgOiRO+ZVD0S1J2wZBQ
h/fygqGQZMRwmaS85ng0Ao3MaN5tg8Z4ZkzoUuMpIYpXdU1EX07ZdWKlgU7+Tv8L
JqhCDpz6Czqvgkfuq4E2dreGR43OSRziwhPurrErDnNhy6F2t8PclioqOG/L1AOo
MRK1qX6Te0tEZzX88C8J9C8OC4mpUxZL+GqZiNwEWh+Ccckwe/KjRqnwxtULdv1L
m8wY+cAyNZHdCibA7XGeOac+4YI+Pykgv2MtjN1/vk9sbEJsg70ghoNZRTxvLSqK
MBmwX9kLAn1zV8VOVKP38bZ0fJBV/HITo0krFT2RjMaHl3e6ptpcH4KeC07wMGht
c9aGj5uesntunB/jloLGKS+eEYguHcACTfePmaLL6h/dP7YO9RI5Z20LZmjQRTqq
Jax/Li7IOAbWlfk2uTBZlkoi8+jKhY3gFvsE8+1ADKx5Twf+f1emwQkpE3jiIojK
MO4WM8sIEyMaRtUDHieMUwKUtvArVyF9eafkX/tINvgp8GRQl/Ckdqu2JyhPKgkj
zzeHqhN8oCfKp5JSacMw/hbeISssBCsTlh9vsOdvjLmykRec+opN0/Cmo6JWF+18
atgfoN+hVdCFbfsRr1lNeH8mMJ+1TKQq934jbR1BPtxoXdh4/Tb34kAWuvY2qZZj
FaEsZhARLh0t6FhFYEtawDlOWVdx1yq5Z5MX3tU/wJAWMoIT3mC28nbVmPBR6Kwp
NBf8bk8kS+xlDFQFCWmqW1+qPm3MXHCIQfadTfmBe78KBVf0ZySpv2b3EcMGkYhO
KwMYS3Zs+moaRJjtnjLgtDIVAWrc+6+uH3y4QUQQWORYO0TdCgIp7BUXmUZcy3L+
Ez3AavTcrAoondTogGpUd/eyn84j7PhLmHBZ7G6uMtzUUGd4cogO2U1ptx1IpTpj
1s/z5THBnd7k1w3iGHpwSR3swbiRcCpUTMekFN+xo5YN4uwk3Bial5dZc47Jm9M6
c0KR2+alTjjMoRwZJrUW2LKUryRm8gktxax54zCwKqM991ywUTBGaNSOqZ32dGaI
foLbt636SFtCQ4dLdFE11auYrfUV5uo4YnXmgtd5sPDZPnfGeUaR5x7IG6xx+/MX
k0kYQGx5ZEHxL9xrel03s5hPbWMYinQ1f760Xwzauk6WhQhjyjyWIXuwTWc1CC84
IGbNzsVu+3GTdY+ohN7eySNcB7SzMSgm5iP6/PQ/SBNyjYJIbpaz/FbJPKKbumlF
3ApNSYiIKcs19P8m4Lns16uA1wOreKBXAz41XEe39jA18SKRNRUsSvTjAUUUE3k/
0gKatxQ+V7ycVGY0RXePUubX7FQfK0j25Kxnewv+fjV5MS56uvo7SD50FQHDk9bL
sVWmDbVuU6bzk3xFNNJYddhEALsJIhVmIyVYcW5cY5GuvC+KUQ/TZ+xfRvVyewqj
43VPzr8EVVbM+9DqrVLQOPYxp8uxkHYj9MYi0lDdLzxkdKC8k5e4ATTdlx21hX8F
KJhwP45SIwpz/U9wsW20vHd7YT0eg1DhzQLqMtejVoLvC/7VfHkyLFDmtYwxMUiN
b+Vm12qmsnd8NI+hBHm1NMhyhW5WUo66lkGVGA+iPxT87IBMtvS7NaYcLYWLUREK
AfGHIM3fXJSvqpwyhjV/tAE3qZN7pwzgFSjcFVhFJa5THoXkoi9P6CeG/M5LfFXZ
30Nw1j9IhDhWiH4J9W3dATP4oVQ//x7Tc7PbA3WHG4zMIU46Fm3kyOPRlce/uIip
HcdpRLqJY8Ak7YtNh8zFVxTcAfmFpfwVwWWEJxD/0H84PAfOrvynY94oNbdCMYRF
WFYEo8WGQoWwYPXUHqUxSkuspgvg9Cuu6Z4sO/PuiIrzUswJZQfulJo/fxBbnPIP
mEEKqm4kWDLwmrrCqHKXH+ugiyKPn3fqbF5g3e5ObhMohrUXMLH9UWuteUMhs4Q9
h7zagAolxOJzsiBx2kcPoOWLMVCK4x+S09f1wvfkdohL71v8Q3WdN8NTD/03Y/s2
SYLLez9lhXTYaPuq8B7lLg4urXOgtcyZTK8+3AgK9xWXfNXVroltcQMjYY0HfoDD
Q69eFNkK0e2q4WB+MJKgl0vUB1IWR1Sw65z3nBum4IyzBGL7d5piR0a+P6qaoLjK
gE6eN+cK7xduy1wJfmLOSIoR7wffLICPCAmoZD1BbBOcAZCRvCdSqSksAIdakeF2
VfcP73IlyiNaizfjHGqvQN0QyzFZeoLg4n6VkRQ7N0/Yro0HcmwWG8XeA+22VOee
ciEIEbR6xsjYHKYUNB/h01pIoeYyZHGsTHK4AMh247lqtR4tsIdMEvu8Q+uolOrW
ZpJVp7VRvF6Jd2h3qNwVm6s8awuSORIYEURkn5UwfEToYd3ReX4br20hXslbzBPu
BOwBF8rvlsFUa4TZHwtTKv69WWnRn8J4hBJkFYrTaeDGqdChksUL3iVYJ6jFUdHf
nmeSrSGVCXidBNf+IaLEbHhRU+027OiplBRAj1Jioan/4iRlBz43UqO6QcwqqrQp
wBBiwQtNRNSTiullj6kNn1EKgT+6iSD2rO31nUGibRa3sVgyxBbEDB2WesTc7n3y
iCV4Hv07eBvwdyYJ8QOOiz1iEqTtkCSTiFN8mqv3iO9u+rLgbEkzbp6oGofjb2VE
8YgVEUH5puwkpu36+kte2dii2ZAN1nlGiNVrPiSiaVBVPLIC6QmgQUyjzdlO6o0t
sGs1rL+wDeUjYcSEbpOtpoincnW1kUJ3kAQw7XEFqTZBwUuIuu+zL9YdSH0pr2do
INiKyaGwEbu+9nq7a3ccn10oyB09cWlqOztCQt/DvzaA7quMK7AIXlzfW+1SqjPS
dm8m9IUi3fg9PbAIGuSCH02HP/78aO7EEAjpzE6pBKMPdsdJyQB0NTSteXOBcZRq
b9ABVWRCawpB3pPUq5W4TJeHSic4xO/CbZ8Jexvq6nQ04KTXm1WF9uLHc1cHIckh
Bb1cFDNLYzadp/duTfvP/oyd/Krnex3GFSf2d9RoBRGCy72BDTO0RjhatcYmduHk
NqaKqTN/r3xy7ey87mu/dntAW3caDbA1JlHuNV3jXvh3H6hGDAJPmJKczAoAp3F/
BxOW3Dsxfc3Svy6Gt/dawdu6z37zINPegfdNCOrEYTNFoz2RwsyXwbGwUf/9y2TB
+xdOyqSphuvhLLaYfy8idAWGOhAQfXdrjDMMSaFeZa+BmleEk47w9tOYDOvyp4sP
oA+9CzkUMhKej0OB03PM16UDGlYL9foZ5Fok03echIi4Zil4tJQGzixe+HjJhIz4
tCheFQnIMPjR3xaR6aYSTwPEXU9f833zjsOGqJl80yGdRSKxtZdhcxTDQtOB23tj
SPxHkq2sxJ7oBRvpmIiM7sJhftyEeKEicv7TRhVPJkaJUHwnw5ALSZs3BC397pSM
tfSq6XTrZJAK9nfAAySVHw+FBjzB4gEwh9bcAokWkLn8+pPd1iiEZomA6JINRt0q
Vez9N74MNAhK8Pn3zLgYPI1GSRn7684t3zmnS7hiy2GwvsELRSorBhiuEC3969XO
eLAcDW5U8VuCsmeT+HkfFsTJ9y5/7P9LYnPV9+YiBG/IfHxQAx+EIlRsAEsi3V1H
2q58/XcVXZ8010C6FlK3YDJhZUxF1bkh3E7/0iSYTSzY7SdfKyPqoAyRqFt/SFda
36KzPA7B7J/t1S4kfU0W0atuwux7f7R+qE9XVyGDEHNiE64ffhhfLHJ/lIkCMmKi
9X3w0H7SCbA7CMOGGt1l9OeG/Dk2o82y2aKZXUXgh3QtxERNyBRS93toHXgS+e4C
ISPWxCiInSsOAphNTzIhI2yumhpwz6spvFeb1jbuITFGiXBZ3YqjniDZ8Yog8n/n
qs0RBpAwUbaAKmAuCGUhfbvkFyCfDehAKkVDlvHhkTtFw/9Wuf78ln0Dx7IfY8VR
LU1LikFAUuINw8QOrUYuuZxX2VqdTJ0wUsEBgt+wpob9kdX37cGqo6iq9X2WS32s
dFpWlVqMJB617QoDAIIQeFxgaa418GrO0Xh1l57gBDDzelC9+pXdox/B2XBGttMK
bPEENUjAoRFpusopvUc1lbaNz1Nfso6JX8T+u3tJ923mRqZdHJ58jzRH6ImGtNCv
JkpLIpt79cL0FBqfvzLY4/Md07WHxvxgQT89dKWJ7rjEId8Gnun2KFyn7k3E+RLr
QRnu/47ieQ/WSJbN7GgVRVTeBrHv0zCoS/fbcvjwakJS5Msp5qK3sqUniczA8iLp
a6io0byc9TpuUP/bcj4FxIVE+6QeU9krzz32KJmCT4sQ4M/b/ogbkrrmbZDWXhLs
ieNFdOfTKOjXknbwG33Rsfrb2vhlI8ht0zLi4Ljta4IgnO1d+5vfVGKxEM26JGRR
hS7qmpW0X74mFFf/TyUe35tOCjfJxzoZsUxlv+IWzFiFREus2YogCY4qlsD29AYl
CXXeVal1A3QwyVD1JUDvHIl6R68p++Npj8gckIMMgVLxsYEw1yj6ttb+ZveoNj0A
vzDrE+OBtVEdDSwnjNpWdGVHZIrZEeCYfNvVQqe1mPvWrAKwyENyJfbYgWV58AN5
TElIRGdLN6+WsTH2TI5Jj03aVopEKJsYTtETxakA5Lxcd4Y+g19AGEDXpVRdTPux
igsVk1z93q9Bs3rQrY6S5zDe6kSoGzBd4n7orFE1Uec2jVdsPSaTpXnkPms7DsYn
p3MEu7ovvRNXZDV1n1nEM9wPAHTGFzgF8P1cap1bKOIdEaJSdMkJGinlmdAYZ+uU
P98tFOMxRngKubSKdYhF4BKCYox0HVjG3LYVthbsBzqUiLNOjUOIxkKPOQuu8CED
tnRYg9qR9sHwbOsYxDBjvqJ333tGNtDDQ4NGQ2M8zR2iWAxmTnQM6JkWBHIC2GDn
wWtezG1FN2wO+D3KG26YFqRplxfvJkSsvTNlQDmRluD6v6mq9T9WZQrYQ6lBWtBI
MbzYv61BNyE0DRwzDAi0Kq8ARw9kxjabXZUM7wzQjaBaJ3zLA8gI7dtbpDwwZhLu
ICofGSsGeScuhX4zVgq4hPeGza+aLjvvSIMj9k/hq0JXUNfAbsKtsxW+c2TWIuaJ
xeuRhG5Nj/+bpPSu/TXwDIRDxu4sLKZBzBxQJ16YBo1mS7t5JzXGcalPmVrBORtx
+zTNmhw8nbqDJOAag/uTbuven2/JZKuMeanHpTYleoY4iO5VPFjY7s4jgOw2EWah
A20h2UhPRSflCSicpMz+29+jmcOSwl4oTTcI/6+6AAK9Sc8P4jOCDKwEtduWEuLE
PpUtGp50AsBPGz5s8/RZ4r0BW4w2lu9AaaOPoqwss0F/tewx4nX3tN43PylIwfrA
eb/CR0k2DTSPIf8y+Qg2Zl+cfHfz6OhQZpxacyFeqLOR0adw0ug5jKYhHeRe8EeB
7bDTxxgtMrK4dyhdm8su26Lmu42nTytjRXA9nwn5UiSrbu6BNdfaTC+YVKtFOZyb
Rc8ecy0RClRcPfxryEl/PTOXXQ2y46DPZ0Ka+uA3Od/TYpl+bs7+m9M9SNCHJZSi
muM02dmjyE2I0JcogveOdKP+Ayy1vCeo1+Cs62f/HVrAu3kIDPdB4gbWN/rjokb1
1ESXqk4UH00+cZz45hitBYo35Y4yTXsT6FVuwxT/wNUyJXurIuVmEgdHk5JzN7t+
P9LDjQR7/VhADNrGsUFtbMXnbNV7siPncH3GUA4tnNPDfVKITlMKW+uYmn+Duz0m
N631sXLo0TdJAtXXHIkusAuxkm/UywXCmBkHnMc//HqxbUhQLhL0Iq+ppmAX2Bec
I/0M4whlVTzyDOrT6jefoAimBYkhvQyauS6UapcGST2DScHZ6vUmhTwrdQOnR7dU
sLniBLB+DdAqV3G7GAs4mS+EgC6SB7EYQc3djeM8tvhKCPCXPuKd+a/E8tLTpPvB
YxY30Ug6/NQMlcHi/p5b6+xtYjM2RngzGD6+oDS3YXG/PQxUunDHLtKlqkr5+pg8
NgyOfYznAQNbnOqnm5ZEh1QRjFVv7RoLLQTbOHYSjx8gcpvhMCTf0GBAx9I0zj1x
SMA8yV6VeBXUj6lMW/BJLRs3Riu6BfWGdc6Q7M0BJQFwjaDbiMVN0tUMzfews+HA
NsA3iOOOnryjw6VhyVBo+VR29wZ1Dta9Z0bFPwm98TRnA4HL7FFWjebI//xjKYx/
7tD+4Ht1NXUuoBFjCCLS9xFZv5IoEUsfiTUOAKOcNZGgr80zZXJh/8s8SHJ1gyJm
7G9IEvMRLhSnWTlDzb1q5riVdJPYZ+ltSt8gKsyT3ztArHGCga1epq50/L62LATF
9EAmpCl3cH7ukBS5DGWTKB6cyt+LOkwjiLxAqmYMUneTnOGl7sQO8mjmaihNuu1t
kCdYnJdZRPabRftjHrGUBS74f0AGqKqsK0yAOj9y6dsgpIpGV3Sq821AwkXKXsij
aR6fwmSYz+etUsbLPB9JwsA7AM4zTzAucO/6RMM+zME2V9aU/D/0gMZlBZsF9F+d
wF/aB8osww2AxG6ZPcSS2y4/+CYn5Gy5nY3X32vFxVfi0kDwlPYO0I4bvoVv9gGL
idOJrKSml6e0DqdzrFR8p3g5rrn88b7DZn9sMjFfHsFCYxtvXFfYXE5CrFZG2FYt
F4pq+hpQNVXYY/6UiRiHnvhGGijqdkFN9JilIklZfDw259CK9E/O/QsSaAHYBK8Z
SwehbmWf/txhuFeKi/0PDyJqnWUMQJYZ+QgmtP3ER4mev7epwDw8ywiH7GhvEftZ
kCtaEazs0f9UHJhm5Luk7PixKD/SPegMKeP1m3iK9cu0deUcqoMrVj5TK/kBU+XY
QBfuoVrC+dKpdZy1jMrUhi329DXgUd++2jIUPccsk1ZNsUMCszERCgSS7gD5ozN9
B1eKmxe3JT0qi9iiLH4K8r8iY0Ux8/Bd6iwDy4nl2q/7fBHqGOm7cxzNTo8OEozJ
Ybfzb92+Xpbeie8pLeYE4jH71eIBv8TLYs2kRlRl4chntpKUv/YajxfEFdUtSvoc
KiDVyPJJYfFhXwbg+cyRqSE3uP2UZVzlAepRkPac4lThIQvi3yBKwtpvUZYjDKIR
KCzBRCYhYr5UuuFFl64mQQRpzi1Tba3HoCSHQQxUhpqRxNxGIK+/xgTSL0+ronaG
1ZzJohT3mVFb9hv1FtUfHPFCeTMUoFRdL4WnIxXD0mPijJ+5i8s4aIiwzc3YEEBg
o6h4N92i930xA7ce8pJ+SNHO1xSsAh0yirpeqROQRLHhyVkmHPyPi19BIzCQouZm
84cXufZQ5dUPQbkuuXoUvE/4mfGFs+I83odZN1+1v/88UWINERIWMARbGsF06KHO
F3IceEYy7elY8gDhEMqe68tXpYGTzkoGeObBdQZNuhO/wEMQ3vQvCoLL8Af6qTFr
yAhbtcUvJgZZyLRCn/UgLIsaUBeh1YirKOzk4xaIvTWekb+h83HYlYwAC4xfmhvi
H14bTHH/AbtwnCcNjzixrOADwWUMlikYs9t/0vurK5lR4INGParusCcvgrY42fPD
RQkj4XznRkrkeE74H41ubRksgY0njusjleSGS/PnjbOneRpz8qdkTn/LUF3iYatr
04vCgB1cKbxCxsMdf0sQDShxVzxtyieSNOglYYn0g6o4npsaQxQ3vbvO2jR5u+RR
xioRsDcPpaj00U06OHw16DGN4z6xFb4RfKgPvEgot7P0c4ESvGjL4B0uAAsvq2w6
yEjDqIMCu5oiC4vCso6bosFadMbH9M+Ljity72dh/CUQHggwjWMXmoqY7D0B53uB
ooYkE16HuXRz9hi47RGi49ek9XKaaxouYsYR6TJFPOyY1EtgMIO9JN6tYfVF3fky
oIAqqdJjWNkUJsD0Aqf0ZPY3XsRvEiSEhvBqX5qDqDLFCZK0fLG9cKK8dbU/t50o
7XfvBdiLeZke1gzAtBmCqNQvjg5QnCYn0NSn8+Y1MtcGy6Hy5kEu9gW8PZpJ8EGP
hf/Guv+f7Va1+qS4jHdFPlrC1Y7afNC7M6oePWsxWs16MiX0zb4o67nV4XkLE7Hq
cKPCFuZNFEKfljnMABkp0SZ/9IYzd2KW0NobKLdmf2/gFcILc1IQA0tBefmejKch
KG2kAkvTNje27A/p1F190tzsDmWq+Leyligbv/NcM5utaU4yL1ppTxzn9mK5nlA6
FtIGbIRiUl3slItMA3Pzi0dD2XiS+wSptALI3VjeOuDerw/PPP8EAkpWKsHc3O00
s37fV9liTYy3prLmoEJS9gisbTHGsdNziGS6009SCtUmfD1YKD1Z9iwAHa4WNwF6
vHnTaFVby8a9PgIE7ivY1D3K4QzeP6rQFXA5jkuaz7HAJjkgfB957D6BcIKA1eUT
IKLm06IyrdrgD8X1J6AEy5X521H4d+iCTl+sxxQuW8Zral+rmsObRaRu4kFw6lGB
bgStrVwuHBgAphbBsWY7efxDDoaz17lcjVAVI5hwPiQvq7Etaq7zUIOj4eMBUjzX
EAekyZcGMWsQz77lAfXrOrEm2igDlcHJ5dVrZ3K/HQ0kd9ZBJSf1RpbjZloE3hYp
ttT9IdHLbmCGjfGRuY7ftorV98gHXBbzn5QQN7gtKhyqHbF1Yg72Stp832wIXRjl
tNKjk/cAIuTeXBauncgFtYTDWh06Q5djGVA9kP1bOvJ181Fn6vZniXEulG+jdi6e
PpoWKq7b5OemcTwApHJ4P79K60IDAeKLpCRvHzmRW9+/OBrd2EO+V550ItM5mo3i
FsWfJaEh9R+SRKI5ZFeF9U/bXGXmk387fsEkpe7BSUevC/slJXnyR5XnNl3AFaFF
fo/MkDIeTxWVswJ82Fo760P05rtn8UxTxAykPed6/atHThWfULQyu0WlbJmudTWz
NHnVmLuGtlM6wOG6IBwNpNHzEHx5rsVlwW7LfwiBKxApArA6lKYWhGYEbS6z1CM8
50HMvReThKlvkXpHLoQ9Ghl8hBpItTZ9fp9sbt6LgK/FGhh/ABNrLCGGCRaQXlqI
3DP+CMDQdMxfQ6UnVTySDh9t2We0iF0T0ciZgPTQV4vRaiMqeIhjZDvfKJnppXGE
QyP5Ibift8Dowg5oPL3sIkhgwT/JLC3pK+2XdIsZFdFy9Bt7jQIzXFmx3Gg0SYYe
5GMus6cvZc3398RVsQAMD84LhWcADqKWIDKibfcXvKBM/XQ4RhlmIAd4PKJ80hbQ
lz6n40mjHVoxouQMkvEaiq3ksqTLbiU7gejYT0gTqLVKXkciTdDtAghL8jfyfJ2Y
/TNJScD0QmuqGagSGww9msuKDJWthylf09EFrIDDZ87VYxFVGOEsbE80pYvVQNUU
F3clp2GV27bPFXmugfnp8JZbZ+ETnX5jeR4CsdNNoI1Z13jW+mydNuNtu6Go6l/v
Wj1AhG1gfIA0TlWR8zx7sHJ0jipkHBRdiTmwXLMr1+ZTlqhGJUP5HsvYVEMb6Kte
sRI8UP9hA2p2ykNVRj2JVWbsbkf+Ar3AA3vPslKYCxsEh0AojnJdO3kUL5Fp5CbC
TJydTKmJS3PMFHazq1vF/5ocptQI2PEYgOUQlw8A2B8a3fLgw21VB5dtieQERAb5
otBB297tFp4urBuK0fcrTHrHKSPrKzh0kkDakkVih05+Ntl7zN6q4xvoi0jCxoYZ
qGIv08IDWJvsORQCw9DsSxAU7NU+x/t5umbSFgThSorC5x6c+QztC9+AksWUkEpl
piJfPp+moA+G4Vm70YdwdAIQ7OfhGTzJDTz/9FhOvtFg5vfoqVPoTeVeyKHMAfTq
v99AQKuc1JpwVXC50ZRHlZdvR7edL2w9ni9H+c97HaQqCZhMewl2Z8vKT4cGt2SQ
ozRaetxuAeJnZgYtRUJDJn0o1Wo3Zo1vp7qY0/2YRvCd+7h7ny6K0ou1VK99AWjp
TybR8T4C8PnJSlGwRjJQM47mjn15F8aYktxhVzaxPsmJkcvcqCyPilbC19Z6BWAb
7n6udXTvCeL9lmFh8QFHtKn8tdwCu51MDXlKYVaFvIFPWEzIedPZe/aW63qXIAr9
SpT6HatZzAGh9PGbViWyhfC8Mx25wcbcloZbOObdR+8FKMiyxL3CLUvLMQPiy7ds
+7nwWyRZHE9/f5xdKGLuUieknl9/qHgeDYVP5JwatbqUgFe0s++h2Z64jgeAlw4/
258kCqz4sQD4FeBPc2CfrIKMUWOhF8UnvBVOtaQ9WS+BrN3OwJb+208l1RNwZjjS
Vrb2qME0y8BG+1NVNpDwfTDBjPNO4WUMBXIe5Pm7Nwx8SsPE2NUWp2frXHApzDiV
aHXCMyIFxgytcd6kauJQmKzJ7ezek6vzIiiS0+t6rfWkT7Nx1iogywngNRRq7DGv
M0pu/hCWZi4b5OWryMECdAXhuQGOpFoaroV6l28ehRmgVg/Ah0svURFCZO+KLgD4
zZJrutg/mLTs2XKEbkWu1iMvGWm0UCBofWXS4KFG/hQa0EnKYY8NltF6H3KOaS3a
bnHHHzgqgHcc5Himu75Y1OWw/pXf45+iS3LQ4GMOqytkjpVMi0n5bqgsu+H9dBsP
yeCh1ln/moAz4NzrXzNtp+Z/UW+Om1aQd9ZGDH6yCX3rml5k5TeEb+TxMa7hLtBr
voLDMV3wu9JYFii/FBQ+uI1L0COgkg7iuedLdHZ9iWSFcuX23mlTEmDMhqt3c+qY
+HrG5HD6+0EldAe6PmiPIQsMCCZs4omKCwWifde+vdJB7zsi0KJQnXs42ndgkNWW
N1ktRIrh4BzR65LSt59W9JT9idFOVkLK1odxfBcoctWBCUdmoPZxGNn+MTi6hUHN
5fvkW0qK7QcMnIWFXLM/6cQAfaCiJybt/9vf1jhWSlwJye/hCoaQVI+7Pxz1dDSZ
RVz6QOWip21LHOpGXqNk+VkTLuAZDfeXP+GIXq4+ReaktBW/x9P2sMVx7Y6uFHrl
gI7+ImHcpcS4DRv0dxcvddzy2NioRigEKzcGN05F3/FU+Gzi1W/ieynYR14jcjYg
He0MjPOz0TxOuZ5ATHnPLGJoiIR7UurMMJxS8aYKXLzVH4d5NAo5a8AHXJlPcxhg
d5fTmw/W3mDjeXqwtbajhwyHVCL0alWETIVk2Mge8/LLId5nCi3PSxlyplLddRIu
zJNN9pBhf0zMsXZGpmSgWsve4qWBnLVwXGONwWjIphLxE/GGPYjdPRbhGWBfrmX7
lvtVOsSAnOl+8rBeXfkHEmoKIY4FAYGxou0dZWGDWfiVHcAoJVBrmSPi5+D55plU
VVn8x3DXc4vBHK32069pZCWaZsCyq3ujeIQdLdCopevzDiIa5wYoqy1wR8MYXHh0
SqtrQ7ztMQQJ+TeG/ecJTvpsaNQrCo2O8yjUUSgUAntRre6x0t+mWVLdDNqmRxPe
0olwD1g3OGRrOyQkxa4cVc++hdJTpvonTVZLUs2/5dne+WAWHiH77qj1BBHiaLYA
rx4Y08fq6304ASxprzcSmGDo+BUnZE9AELPxzTIgpD2TYLFnAaj9KX3xJiA8H7PK
d2JgO3Cdy8dyBO6OGbbeXXDZ3sREvBxhoBq3CMqB1ioWvkS6L6sypZMFu6fGN0UT
fPcP9Eb+MDFwk0k6NeqwU4OkdUtavtEWyEFvWuChAMGd6mDWFKPES6GghStBkRx1
xYMOVc7+2axs2c2OSG41N8Ym3S5j/L+WYW2/oxuZNQiL00VZRcV5wJj/wj6gtBFi
wNaxPIHlOpoZUFNMBiX0t8KESGARzGmPqkpfK6v0fP44yOmzHECyx+h1fKEz9o30
uGIOwUfdWiINFt6qspHCTb/lLyivvA82kb4gmVt/sPhTUv9+BHtNixbhQGFzxMQj
PiCWrOlbjqZOEVqws9+JxQh9Vw2R59oA4Auwej9itY4dGF/MIZOVeUJJD3j2yfqu
4J3Gkbg75GoHiNyLs/vPh9gIDUVFHYUzKIFAUng9DG00VHjXkHg76+GV5I+RnWux
GBpjNDD6gcIR7rbIDBqNiRwfj7OAIB96BRCjP4gNa8o7eXB5mBfvVnm6yc8dqQPQ
/iWpth0kXeF9JqRA5yvwfvFYfiibGaNECN2GsrAiOiRI6JgfAouo3sNgFiduf5C/
dXKvh614ZE+yt7GQVmHll7wHCwzu5Y/RrXcSfXWLjdFI9SGmHfEIyYCRP2HVsemP
pffx/NVQumsTEVTv+5EqPJmrzr/iY8b1S45TM9A8rA1Jicq8fpWs5RqrU21Na6U2
MbAHXd26LBrsUDi180+coqZCi23I8uu+9jnGoxP4+xULJeY3dJg6IoiqV7B6JZZ3
IRVs+skRrmphLEPIyXatQwqaZhv8P6Ky/40358ZwfaVZxnCWJCxxFc9RJP+7hCHe
Z1B2BtN5Nb11IlAAvFQSmn5dUpsPee0EZdSk4R9ItUiL4hQoiVahMP3Hxoa2rdNv
G5RgCBKguo4s52eYhkir302me7m2spESd/KesnOPzBKIsmSpSsgnp1OP6pbrUpaX
2pGlEe0VkTie+g4m98AiWEuTlN2Sx8MhwtuE7CDfUnFgpJlpc3VfSMbV0aMFaJCW
eT+4dMlTdDsFcHMyoDxsVNkjt0Zip3cttavtJgkz6Eayi/asxY4FfpYAuCWJcsji
9M/MQlFxk164LQMpan/4wHhxnvD0+zgbQlsG9Z1+Y/MSQVPz46phOVJ/FzbwzHjt
diPC5kW4D06JC1dJ738Ioevg0Rj8yLhjR/y3wcknHLJmnhWvc0qJoulnTjuOROus
Jibsk7pfaGAVnLpsY7HGogqRCJaKfWQTeCA0Gcy1zxOTlQo6RVwlOH09AgDOCqf5
WiddOVRHoH3m9UkkzkCssitmJrRzxZbPWqhHjWlRH4fCJEfWF05EK5/GNXmiPEgP
VPDZ/RWuqosRvRurWInxHMe0PleMq+qMKWee8nJZFDPrRPXE+tOUIb+G0aCG7CId
eU0h5WKlJDZod4sYFksH4p7XYHjQLRe6midmPg23ErdVfFyuQHRBm4Jf3v8bm5e8
CQpewWHOysEqouWnt6cI1YJh4Dk/mhQ9cYZbh7FPQC8RWESysztde2OjgEthbKXz
E8pdfwXPqlqQTZROE+tleI42ZpODS+rJgZC6Xus8SiRn/9JccmJ53aGc68F3wiVt
KlTzWeaqpnXXp4zgvzQxYnlDJjq8ykgIJ9vkPpxlZzBzXJlS9PC1Uc5a1Y8PcqzJ
zC4jVROH4QmUnGErAZ3WuLmMRkrgK7IPJ3x4/Ztw3Fb+iRRygzViFnDNVa6e0+Lv
oTgSOoH5yrE+/yOgMLGsmoSAM+Iji1CumMyCcUPVdCSFebVte86unoLtngqI/bM3
ZfHzgC/toejauHmLxl/Q3r1dE9Z+AzWdVlUfEoKSeknBcTLuNlQ8H9uKVCP+KBDD
HpiIi7V/VjilDUwnGuTyZQ89lYMTkTbRHHW0LuEUZbIB7Ch94tJ81S6L9C2qEVsS
PwQRbSrpJ1kvc1a74VdmpDcs4zezRJImOHKV90pGVyeGQvC0FCQKwjjlbO60/fxV
AHiYvWuOjtFLzVXNh+uPQg7+XXgaz0kgkDvTinoox4CNru+J044LsXNUqGoAdIx0
oxet9H5yPnhehI6HV9hdFhjpQzpoZkxIqxoKe2O4Wm9BXMT37f86w5EP+EkVqAoD
ZIFVXo7V3ppYJS9tPTa6ESE9pzPRYbvtls5CBPuYnUIs/QlfdY/wx1JMh9WjfdDq
ew8vvM+m9MFHDo32l6LysJbKH7SiMcJHjSxdpck+dyzQ8uDhe2GOeW9ISN8Ajubd
lTy4wntRlIFh6ZHRr1zNNOYYI8nQUptbG7s5088F4JFeYMyn05ediJ5kXmMyd9n+
QN8J/eeVziW1G8KEhrZ0EWl0lBFhh6VP9UCkXGCmSPojSO/PNhkmKV/2MkXZQULR
kzcKRGAyeHk9A8yN/zq3qKCwX1OPo7M6gEccetMBZ7xlbgKEriyUFodrtMIZN3Fz
yt+QcDk3qcs5W307wpXZn6ldxeOzcHr7fe6eCdA/MSBZCcRvblmpwOoru3gCd4RE
ypwXWf7bI6X4A6jELp8VOjQSGRRTa516PiRQBG58+ZzDRhioe2R2nLRS8Lp7OzmI
ocPD4qxMoS8kVxLlvhlDu0PddbpYIox3Jg9ESwcegbeMUbW5tQIpCR9JJVB75HDB
dH4Y0c/KyNiz8jk2H6ccmpZU4DO3yguGBOQHT9HpxpPmfpBZXxw6izhtDjtC4oMh
T5hjUM1Qfh0Rs6PGKSTgUosMj1Ft+YBm3frihTr9SsZdUVCBB++1svJp8+9ZaMnV
UxC08dxKuMJbz5KVAd+DPZarinfxkyqky1AWBHb3OnP3PCmtROH6VQKCwE+b2DS7
8i+y6FEj6ylz2+TO4K/DxC3GIHML4nRMMVZf8YW3RoWy4ZsQSVnteWacSBpivRBv
tEm9MU0lcO5/efMAqOnNvvXJVnwXUhGPTsGGDRTXM+nrR4PnCySMwBnW16pLd1kP
aRNWi98VyAvOV/iHgZ2QIeslvL1BLN0t/4o80WL5S/eDVvVX2CojArL0GD055KGs
2xE01mgo5tZfffE4NewkVNbOtddLI+VQZ8lSJkJEElCvJOGHePALbSajj+MzVW9L
agTjZ2YbrXC4Hj7uoNMrncRsLvWo2w9b3Zizr/fQ6B+f8HUxg3yEuF35Py/nQni1
ccAINZLezpE61QQaltemnfXQgItFV2CFTt3QnL34fSZtDTI7aVqhwHaKnydQovpJ
tWdIx39gJJ8dQhAUMUPxhGPKugxOLngqGi/iHFBmj5jVr6AvLY9b5iOWcxPzS4bS
wF+fyS4KsJst8wCHPisEXGN885g52EgCnI9fPQ8ftQy8dAqF6ZlXOcBYb2PkUEeD
cEkBna6bXhwVa3KBJ5V2opbSlRSIjA6FW5RiJ+riS1sph/Y3uVSULCrX8VFxAKcn
1ECrFGjgSB46dpLluluE5LKNekucCmNB1qa9K7/kYqCe7xw5OqGgsJQTMvDJo1HS
Fgm6IPaYx828bgXvbS1mS+srv8Zv7Of5DCjt+R+/FbAoRrW1PHUrbl+swmNj8yJp
FzidX+Mz7cQ+REc7VryCfq9zE9TD7HEteOKYTeixwD3EHjTlJNhtRU4ZS/Yl1JtV
z0huFAWCTu/brukp/wBfO6QSAgoRWFRzIuNrfrId1TM77MQGReqoZbXekO3+zCIZ
80VUDAZ7bi63hK4lg8wzNQp9jrr5qaYnIDw7MM7ZFBpE1Jehb00yxEA3E7r1HR5w
DwPqJiP3LROciSr8O/sivvJpTpFskGEeBpcP+VXff951BfDCkg3yCh6UhyPXcEMG
YaAbcgZkwP2KVwIguVVBJcnw17s4sfR9Lyp3i2mLojb4CyHU0BKMbfihbSGMYEAa
tUGHfFVEIGwJvXXCVXoOx3axgEImN1vPQTRTRRO/chSjYDfYcYe1OZgjjcst9GK9
v6TFvcNr6LIIW3BSl0Tz6nEZ1xZY9GFwG6FsT7PVV8vdBDiQ8GUe019KkwBSN2G1
sWRxiUSgP8Y+YRRN5GW74rGzcA0igW3tQJOonTjBseU6cq/yKZxtP4sCCtE7nFZv
GhPNOdxNnrls1e3QKKa0DQvMh0hBXBxHXzS+DPSTATRa6GhbDripp2C/I6VSGgCq
vBH8LcFK+GzCY981JsFjsz6mbEdsROQ4z7vy9O1g5u7gNBgAQQRppWHPuhvlza6f
1M50jsjk/+WQMW4I/VFXoNkn9hT1P8CXkUHyg9t+ptlGcNOvWpgBFTyrc79SaMNR
fKq9s3KHNYi571PaiSHnxXCHp+jRyQTu6LOeN4/FAHQmP6mBgYS0c1IO3dBDQJ1G
JtySwSYIPcNPiK/hzfSZ1yAQx9g6Bz7fI5MH6MEIYzaxtR3+AAsZGN4E/ItQAvLD
OsIBWmsBXKqgn30b70UYtKyjI3dHLd/P283uGGm0ef7d42uUCJvT/v53AAGbGit3
RR1nUlQGDJnbojc9Nf8affwyO4AU3boXCBFIJhvL6EUHNMgWzshdPF+tumYbRGtF
7/zCgDsTXyQDBTHFNqYeXrWKvcIzM7+tKYPZ4aoNAcFTYt6VWWx/9TY7TajtVzc0
tRgjBa4NKwDTVFSLeF1iUlwV72ybIMmPJ7psByKKoYROG5zJmEM+nB7fx4q4Oora
Slbk+zDQr+QaV+FgVj1x745rudH5k9xf7G5H7cQE4/1ZbVFwcE1vxk5lZL4/tQVi
jKLPPiA5MjDcPhdMrfLAfT6cGBnKegwNlT7mZ15SWx1ea4MVV4BxItl0uNm35xrb
nzWAhAprpfxdvkcUoju7a5sdocZ+7qj5S02nJ9hhF8oBbUA/bYUoWlwC9B7p4ypu
nSqbw+DIm2DvvoQS7EhfKPCPowRJ6hYk3+DMFVNHWb175KwJkxOZEnDOBTGtqeq/
hrEY7mSdiIlTIGQ3LrajJlBGEIkRuw3sH2y0+L07V2grpE1NRKKDzkExpDBNf/Nd
D5jmKEpvSaLhqT6G/0UabyM4nnPYlCJknPqOTMlMEiqRuy50oO++wH0alHOu+Obh
gmQ1w1RUMeW1Lg7xDqQJibCCYGcklUQN8BvnVTYGTsE+/zz3EwiQkesh9V4bA2mp
U/mLGuojcPTBGmslVmIyjbPOxvBKVYhVGFBuW/NcwBxLvLeY/kaXxQT0D3nBrQYq
Tc2XrDToVSL6nZdaLZ8Lw/giOS8cb4X0CrgZq4zd38E4qg5rK05peDWFw1JM/Bww
KsDOtyLLq00ct9OdIrttp/4pFsMN1vhpbd2KIVJsJvQuQE2kLtn08T5at/Ye0nBa
y0qxNsDd5IqRkHB5RsrpCy2oQB13pHQZyu/1/AjEJ2XZaZa7wNfZ3HDswZjOq2N4
aL27jF//My8+FEyRkWOkJ32UQ4jsQL+eMvv/I9FgbC/cMckO4rdvLf/RbdAjtVEg
uxMNvcO1vSwyherdEr+MJigdRLj1OG3HFP1CzJoiuEl02n12CqPWtU432e68ilD1
MDzePfRysgyFGTtkR9eHy3wpkk/xEdmorEomZBQ7mHXXzWmYluF4UasyNDn7qI5u
Gi/a4TcPlvI8pCPEOf8GaJ3QQT9irWcpw3tdDMd3eChMaA1pjQJipgrDEuQYGVUP
yaJgKSLLL9h3gl4lmg2IRdYxLqxqweiKxNbH9ogLVkEbNU7Vgi/s9u/attuS8Qlh
xWvNaBqbnugZ/E5NXUbc3/zlMfJv/TcT1+N17bhRWvWGyEDTGKFIGRkd+UO7+Zj+
Jn2WpU0X1mHloLmUZRmXVlToj3YmoUnRn+9uKafeoxYWbmRC+lYMZyxdILLHgF7b
NYI98qmxA/QMzM4EFhhzd+gLmeRPTVsCuq/aV2RWYrJYukWsriUG5f47oqoDoUzU
i3EbeLtH7TxUZbVOzT+MHEArx7FRWBUjgIrmy8p50xiSAeBOB/oLJnLLnoHSaFMN
GQhtnbAxdRKrqquC/ewQ38Rz1ve5uLxRmxOX5qXAUB0mL7kuDFsqCYtq0jMmurST
ubzYNxz/2+ysklpvvn4xhyNx0M+mZcjqs3u1MhpT0KD5rASZIi3IBVhnkcmtv9GP
CnGDpkPvp56C1fNVSjif6nCmeHy6B4EVeqYOfwEbp0MOPrkNXOCRjFxVhF4CUQjJ
btotqNraOXNUkmqVeDji9y7nCM0lNHSpsgnDLICs/ttVElLJNy4EQDeyEtKDlVrx
mjmFLS/lImdPvge921dR5cgCQDEWVZ3Rlo9b03XTGQ/zyRAMKYvUoeeela8MCrFK
UenBTWy+flsx08/iItkTl9YVh479LBwVW7OA4y/EqxYbdjIZD4Y9b2mf11w62UDA
5uiFS9g625yi67ofpMWrszYqiv9M4F+Mro3JFKt8JrzjiOrmzqEh1JDhZNdLrh66
MDIusJk6ENu3JO+lLOFRVopZFV8CCJeboMmx+Nu6HlxoR9MPP+yfIbuAugOo4L3J
lfbPU4bRp77WVvhPFtf0tC0rIAt+pQjFEVfDSuGwF7dL4e12SMHGMJ1VNcNz76HZ
Ziqb39wWmHKj+InJKuwETU56wzMHivECFtlnAlc6XAr9dTqauiKtkA0dRIoTqv7y
Xa7ALf2ga9HnV65a+fL9nnOoj+AVl+GMx17TjgswBf86AVptjk191HE9sCR95y0r
pNpBfGkRQ4pVOvrn8GMt9La1UpGL8Yo9cyFv0z5fVjCnDTcuE4zlAQgKn7dcxOZq
3WKMiqgiSyZCXFcH6YkR2+g+RgqLpd8lwBeTKiieU4UoHCZ4RUb4DiHPjf4bZQrn
zg9A/x+pCSo2ZZTzyE4p46D79SRTcn2ZJKjrSqtHGPtwwyNSEOYEtmCEVK9mC1cl
IaDjBjvytgm8kBLzK7nuj7/ZxIm+Qp4LkRiDcKXg5sh1Gw1aMwyCIVmvp/1JtbVy
plfvHMj6ZccNmcHrIorGz22ehM/k02RE0cu7/rGcaFwn/eU+Bas5QSRj20e7Jrw6
cqNR7J9QyywFEye2jSPpvd8xEMgay/Me/ZW4bbHco8eJUWtmA+zEKy6ymQD5qyAn
uIMKdLLLI0b8FU/8G+w3/d++DvEcGwmpi8gGEYFwznktxTkutBW0SVf97DLYsfri
mvHXeIlEcaysDEYjqIOfpFcyUj467vq0VVpCZMcs+nNXYSry3QIVupwZK3zC2KUE
vvHp3FCw5kEowoJVPasDjNpsEiDREFu2H5cTPcTcyMXGgWrQOIQwGS+9CXg7Yapa
p6Y6AqdII3DvznQQRmbaQSvV71FGCUzWwEX96+DAuCxXPMaiqGIwORUd/X7kIwro
q920XMnPT8+jYOHtHRuX01PLXYmS/kMhdtc7xb/QVrta7cn7gx8s0O++fCxc3OMg
AaFLPC6+vp/NlKdxRHrPpkR73GLgrO/19hT7Lt8hyKdF0An2+mKnqcGq4JHrQ7cT
dwWWNpsYm/GLf+qfRSipx+68WlzjeRytQddTl9PVcoT4ZGKSw02aPv5zaDYo+C3v
KamDiBq3fdKd7+yoG2DUX16CiNs2Q6kM21aJHjWsr2BlJI+OgUfmQm1/DNRix2IM
bBH6Svz1Xn1hFOb84hyUl1ue1adU7VGbf99nGRFrVyjUXaums2PDSqxdrSL/YSSG
1+Bo354aVAZRoYcpq6PsJxSLCPCPhgM6MzYBrnIW7yQsdVJnIm/q86hBmLgDwH20
P2TlTMWomXKa4iivzOOcQ+412IIx2Q6bxRvcb0zAvb4RANWLYQFXgj79dfZHdQcc
V+hAbAJHg/yfZA3huoZN0d/xx3aIk030/Qs5eI5h6xGY9X0bNoEVOc4XdXbf7V1D
PvdVOQ1m/hBIfI+O8QriNaDbETiFymgIlIcni2Fsh1OPymPD9tLxbw5A2fyxm438
n8KeCCywi3wRE0H4fBzKnuzYKx0OcwQhnmYz9R/iJHqA8m7CRAx9+K8sfDlopu5a
wm5A4aBw1QavSg14kv6VhmK4TVNgoyNqt83H6mubgBDR1z1yj+RPwjrNS4+MN76c
fpCzUPymp80pygaCKkcRSZVi3x1cRjf8jAyKWQm6eH+PkvKnAOO9PU/a1L/fWPFo
rEzL8qhUqimfuEXTX4ldryLoHn8A3UKimHT4hGOhfjn2p5kZA4rhgEz4m/IsxNt8
Qg77tuMiHk4jJJ7XIoYOt+uiiFq37ErQGeiMG2hm9C+PLxMJYXT+/H7D1kXPrfEQ
Sdz4bMQvzU4cpu8ZS696qM76rx9cN9yYU0+Usd1HBeLGSnk/ydPx/hLuA7E7Bpxh
4364DRJgH7x//BDQVwCTMAXuPbmb6fAXTKJEOU6lRrLpamRfh2b1xBEpNJV5jSOW
sfgVgsheXvsD6zgNs5x36nHgPyRBag2F/m8c+1wBVFBe29KdPgFT/SaBl3e/z667
0zeLmBQB+i1AgkP4eYowfvJ5RAWxGjoEt5BJN7iYVeoBLF0pU/hOR8d2ijDJkyHj
lnDMuxyBSVghmr+BwotCsVBL9jySRnSc/1WthLtAZhzouiY0V9olxXCeDO3E9mEl
q6TwLgN9g1YbhKlNikxdGrIkJs4X44N6R4e+2U45c5IB6fSTTYvP4n6DpKkyeKpv
Nw/3kqOYaR3oVVpU83VBmjc53zBU1t7jd7Bay8abJ5i8a6bbjLBeqzU/9GetzHbq
0O+UgkVaJOCS19Uaf2SpOfA90N85MtU7OzluZKcSwAhvPSCYEfOWuixVhyqyqyo1
Bo79RpMmZNzdAyS/H+iFMquBCiofNbZRnWLoRNbmOE43JlAM/hxK/MG5sRL5vrm4
fNTpPBm7fM40Vox7K1kaf3E4bWDiawPwpYtsJJAdgUjP0rE8l3vD4E68dtk2PHSG
ipeAesJvvU69iMSsbAqC8Sa6jERgjlRbDMhLPTfhQIOucFDijWWP1B0eQo8WzXKH
m1wkoT7otIW7u6FWNs+dUzmrbOg+eXEA7ELlbU9nhgbitKrwJODqqWQEs6ha4G2g
LEo4brQjMYzq/QqfYLXju+mJfjEcrSkC+CK0qogVBki37FGuyb7ODeDl2s7keeMp
9SmHi2K6xi+qGAxKCTNvajX9x7Sp/3q1J+G94S6GlKifWqE4gZt5vM2VejtOqniC
yG4RDD+gMkdGbU1ocITHe/gJXZIJUxSzRwxWhNLZbZ4H2yUrsL7QVwLfsgrd/9Al
JXAfSHf+G57OpSvOJby/OcnbJSZnc4Ec4A4Mm/CcQrUoDLuRucaW07wkr3S5n91r
V3PB6Ukr5jiQldCqBKtnPy6bS1cfACS6qd1bFLqAV3Pq4Ftc7F7I5q8ioO9jihLU
1UonUtIBPpZZk6BFF+PjfRkO/2S77QowQ2RS5f8vdet+oov7NpJ+JhWRn+A/96dO
wyt4BzdvOlLB2/LMic3pS1PgDwhVEUPvPewmzbb7KQy8YuXofpubRvElzO7yO9wb
hgxYXzeSM8iHBiIO88G1qm3FjYnlSfFQVcI5CYjSQRjMcT5f4QgefOmR8iKtpW3y
SS6vpCmJP5tYBTjFSrU+fKq0dS9QW4IqmQhxu2uflcsnbhYM677U2iGLXxJAbJak
BznsZ6mjZgQAnw2wp/+0BMRK5D/CbjUrZBkk5QvJzvR1Jgdze8jbGnkMaxKp/wgq
NdyjqVG4I74ocbVJTP3/pjk+7GlXU6/m9unYYVtWB0/XQsDVRHy4zXdNnwZG+rYE
FEFNqB3aX2V/Hquzyf24YqQsdZzMhZA1OhY73ymyFbMTSfNM8Dq1Xmr8s/lIixLQ
xYvljHLBNnSrkE95WXDvZ8ok4023kw31rGN3gx/kRJ7sRuZx0uRWhp1JRN/Deqq7
1Y/HbnnqJJ/Wc++24IBR+leVU8zsLaifwDYoJLW4+Its7biWjUiXDDw4FMUo6D2x
PEObz+xslbny47ixDyR1+nA8e1WVUgqwDlSOVB/iSOPehPzmiLt9dM+3MsvH7gct
JNuE7TfmmmOnGHHYHM0rz13543T77M1zNqLzJr+ZrTdrVlIftcKXInX0XZHy1qzk
W67/VjzLU+bACTUHR793RI8XTYM2xZDUo9PYtP5kthvjwrmZFJ7WxbIAAjgttKRJ
5L1Tjjxcs6G2qyhJrWfOPG21JIXDJ82b0nFzITQLi20wNTv/o/Wf5e6QvvqMWKfe
WQ8SdWP6CNAhVUyVXSUtzMcEpEmhRRrX3ulc3X3lVj+yDaYoME/msc9vXg3I8pqm
uJ5qS2ePpcf/F7RSzlzF51wlVTrcmHKCqKo1Pb48RCldp58wbCq7FcnWjJWoI9oF
XQLP4WmbrNMVz80FlBrrek8YDRjOuH01sJ0PIBkeF6EEtRA8pSJ/h3nRkYhITPIa
PACjDocouf4B3x0pbIX7OXlR2SZA/H/1tt1KPc737iCbItGs4ZXaWJ/syiMsTXEq
6Sd0NvjubAE39KES6f5atbKrEBk03rq38S1ZVbzFNtfkJwDJjBVKvg4ff8BgU0xU
3A1MJSDUBLhIE3Tytshnhf4db41gzRwncvXNimLXuXrJrR3FrqdI1N81kHTIEugT
ZdN+2XxQKqpLk0PdCJWk51ohDEJNCuJ6M6xwWgOt81TyiBfTkx3WPAsMG6gmIoTj
89EUAOB0QlOBnf2pmWgqS0aTvJG1QHId0gMthIwWaq1DMzlP69qlw/Xrcsr9t/B/
hMqzOcMccHQTe1sLPhv5Si10f0+qy8eKKWwqUHoGAM+2lR1uYauU1w15ZfF1cZpk
tC6Xey1miMOMRsaAxB19WKvgvN6L7OX1PldvMbfIFEKMHrVAF1aqweJaT/3cjPc8
7Lqn86Ogu7EaGi5T/alAo7bV9kE5lHvTRshHJ90sZgrQzt30qhzFJh2i2s7/dVeu
UYFN4mS40a2eYzlglo3MbVCkM+gsAorwxzOjpu/8gb//yJb4CJAmh0ENq+2UQTTy
jycKUZA8Z/N3mwdIDGQHyU+AJ4i3PKIsSalmnN32DGY6910+F3efrHCpzQYGaW7t
bcJrm6zSObVpCAqe3omqox9pZsk3G5ch0B/GMp3qUGTbAMZS4e9dsFP+vZhGw92U
VmucdHaZ5xfLMoyBufRpWOyspJ0x+dFbaZRW+Vfg4pE6PyCBSy+OJBv7f1jQHAru
r29vY7XrtZmN01AJv5XXhLV4qRhTtIrin1bAMouyuFIOvoDh2zbNY6Fs4V4WWyUf
U/NEUjzUT1uk3Pcsvm1bZfJT81S/eSs0xdGXRoRdNCjA8FzNmx8EtEs7MvQe6jyE
iWgr53K/jw7jbrh5uQ0qdZ8J0f5bi1Nb8NAC7mjUR+mvaG0y3ngqjQ+PEJATxSTA
hiMXd5MCHTn14RJJBno0aDdsbyq8ZmkQtEOpzxJM+Mm4YvKX8A0RByYMnHQX5K+U
yKTiA2nVVEfnHDocY+jUw6UyTe9bYk+XcC15yxQy3gstHX2woNV/HIJ0LojhEt4a
z20Eaa+BMbRkKFUqfhVMJkhj5ZwdtqOmgtfwcuU4KWQkoa8ONFggAam9uJ7p6xT4
AJ+wxmovWge/5QjNcepSL89WMISeu/wYT5d1wwlbk3x0xLe+SmozCrwyYdo5tWD5
sLNlXl1tq9naFYNtZb61emYBe3JYKjP99g4PTgKbS8cNh4mhn4tICCYKGdvq5xff
1/JcKtJmpR5RBhjthVNfQjlgNn5DUQClo1/StenUe15EcYrDkIxZp2CheAv2y0J9
jHLLjpjH83+u5fba1ypi83hWWjesSkjlvPainqek72calacubm0/t27jvWJIT+dc
ltWIKvJNLA400zj+JQrdvOPkBhggi6ny3vIoyH6UafDMir7c8iDGNPPG5KPwieWL
yyjd1RIQ0luU2AmeoTjVpkrOhyKjvr7BmhsXXJSGKQFf4ox5MtWAlfXk9bC1Ti1r
tujn1Mga8CRgPX53/f8bjxgUiCqGUN9aywBN0Cl6uIGz8wg/xxaXO7TijVjIPKZ+
JH1QywjPcZ8gXlcFeCGc4rjMhlhQsly4oGZfZ7Gx4GD9Txs2US3R/mgevAUCw84x
h8wrP9uV2I+0LRD4pI718uPGuWF6CRT4+VlFD2/adkQ9rOsajhAq9Niq5mUwL1Ac
4IDZUVzM3sxh/EVEoyNjkkO2r7D9DaI1hwYeBDwbjAE+0fNjjq/aXwjkM5P64Dla
U8UnIL9+KgAuHMrrIo2MoT3kKqbSDEsEd/vTJIivRcHmLwhDMufbdhA1MoLIG0xm
KQ0i08aIZD7K+drsonUjMiG/jXTnrbKbs/2Lqm+u22JQD57Sz9nKuDZo+3j3m+Xm
JDzNVbVHxJKWQ+Le+3rPYkQ6g0gBy5z8zEgg0b4f1CGXIretNhomDs/LzYos075y
EtwZUkMavXLvBTFFpJtFJ7Q1WEcw/6tVgDeDGWA9eO6To3pypIJVHSUD7hW8Ac2X
0+U0EFj7XHqKYFftq8Ox6CHEKVh+ZsziV4KPecyvCWohbOZlKrr6Usa9ISyOm2+8
2zzxqbfCKX1HSY65ZvOn5C9RJyWhWvqvDziG4kZo3SSSS2SdDeuNsy3UsX8aR8av
f5y5Q22vxZ5kxFRM0BtdiKbr/GJAWjzSrIJEVPVhKSTo3b7Blg+QJYomZ/VjMYxA
N61Kzmb+MX8u8hxUMzpurXwft9BJnVOiWwK1t9eoukc/e47otHqnFrcG9W0KnPVh
CeDZQN89Yz1Vq9JVZXSTfFduAWuWFy4kufCou2iEOcrwcYYT43m8DwHFq06WfrWJ
DxXDZfhTTjv5ZAiUGTHqMGn8KJNeewE3LRW32tqk1V/CxW49TwgI18bwybvXQgR/
jJnDrtpkLjVnUHhRTYSxzU4mA1RJ26t8poO0ac5Q7WcYkTvQLpTZi7wQkMP9CaKo
XriT4+AdO3oC1+U0XAsnBI2PejBFf7yO/n3XBVZ+9WLA+F2Z/eTGtPuNDRSGpRwp
NYRPfogw1hkKYo7Fr8SSPZWlFj70b3A9xhc1IuQ3B3fIZuXXaWX88oqNJm+lmzEd
ZQH/QiGFKPBuvPo4Qjv8E90rj/xm0KGlBiPVyUEP7uSjXaSiTCIUp8lUoS5wVq1l
+9pPKicjeVuhc8OO1rYSwoybJxdt0NmN4DWoKEjc6a3BKWVmgGHYPKxH7KnTynML
VVmdJMgcBgUv01+TQ55jxf4LWFXkjBUYjoQh2mGsrm98CeTOqf2kevu7a+3naglj
t7xzWNmNg7VtACoB9chE2C+WwpIxXZ64o2aBt6ve+Igb0f3d4QhZzq+Ve0ao+i+n
gTi4xZdUSJAjZRiqp6SR3A8RmdOvF4sXVj9mttUPm2V3Qd02CAL5em4dzaRghUtS
0wFdU5bnLB+wGEEEItW0enIfPFZL9S2TunbOrZAKJ5fm5Z+FgtomksWod0eKF0vC
tgwp9V85th0RHKprHkmks8g7Rkp9eNENaofIqJGaOxm2oI6WzVsjHZJumsKvfWCu
Nc5nZOEIgvWxN1PguewUkPtM/35cngRxqzuA5yY9aFEIvdyqxhA/eosD8Eq7yEvK
ubGH6wUvVCdDJ1SGT33JMmjOP9di3bdEXZ8WJvyeZ36hmA7yydAiKqRd+tbhWZ4s
SdtIsNhAq6O+B3BoWN1fqLhr6ecmCfhJ+/MfExhv2jP2PNHf5xJxMiRpb/7Zg1kE
QbvAMBvPt9OWR5gxCu+5EtZBkv3jEAG7oBoEo9UUtoTvguEwG/H+dt2mvW+76QSA
r/f21cTB292hYinLJXJOCJMHkzCpKIgVJkzqtM5uGmxhYgnPLYV6IUggG7mEAom+
NHxFCrJAGs+QMyCFnrR/JfyE8IcqHvclHTKLGT5sjnqas22K4IRJy+rsUSBUUiT6
D//FCY32irdL22ICGUM3hK1DZK8yvY+8B34bZ40ntPQ7LA9BdhWAWiOGPDlC8IWy
B21iHAUfrc+zWDE1kb9SsxSeg1LbMfs90JwuXn6ydAfYO0RtEpOxsabxFPNGyGiN
iZfTHtGGkn5jKzB5sJ/DyR09b/Xb+hIAx419jAJGgVK+VpKXM1B3b/roOO2X/Ows
T3JpiVnWvKL42AoO4r4FlSvpTtYL9bbl7jzQ8sKXlf5OeP/N9YxyCR7/ovUq1Yzv
d5CmAE+D/reGGnQVF76IJA4GD6n/799FvbDKldaSewL3fi2Vce25WgTimhM1/Lp6
oPR/edvwg4ZmOqlPHHkG7tPJwhSdkrc91W8yuuVy5In9sPH0Ma6YsypcH/2JWeIZ
wDezjgu7HY9irkT07rxBDVMNrJ/SoAjU8ls48etAJqJk3HxtrhkFNNDEn2kUKrAc
/H3g9nNO1CFOorta6uHntb7GGShlf2DvFwq4mrfiR96F/EoEHNbpcs+t7quv6EeZ
wrX3shH8HRI1o/7BEsLgrMJwteO5sq7oVI9KCS56RGsl8kwau7IitQBwm5PDmtvi
KlasNdjgvIw+qkmB96U5YnMviTt79ecYg6j8WP+/6WJNo/NTNUmvIHKUUBbu92zD
LAMr2g5I8H2rUh3tdIPOdF5rMT0vM3Oxy7wyxvTCqCLUO/yMR3HX9Sim73QRxiWp
sjfawZ1yaLPIOu7mtHBedKlx3ZW82WLsuQt3gzhUuhmyhEYDq3EKYq/M4IkE6cIG
gtJzDwJW5LaEBGHq5LlKk9wEZ03eFiyfpxuNYgz2wKijKhhkk4AmnVDsBZc6Zx/A
rZpBtLzmv0Hghnw6xFgAXkuU4at8CKogNkQI7Xb953slwoyptbgsrGekPcE/wJSE
LxPX4GqBexqlZbiP++SmJCan3qx/kPMNJK2hac8kcScP/ybIaCJrvgKyXNhTuTXP
gTPKnooqDi1fGwE67hbuZBx1Qsz7gc0hGRCREpZeaNWsrYCaackpnu99wR82HYrn
DvweZoLhwGFa/K56XmNQJr1iEVykq/CRlJ1A+XTXAsTZH/Psj2skVxdVg8DXQ1PR
1M7R/yS9YCxJgs0Gfn2Ko7Re0+KQq48ywmpImL9HiDqyCDMwlh7VJ3HVqI3mA+4/
YM7Q9DXSoFBT6rx2gBJbEWvtHy/oSOCsINBpQTyyWRcR97bbNLHIkJ6YKSL6uA2t
HJD23YOELC6qjkIK/ax7eI1IdoOPvcNv/HCzt+BjIJfZiqmibbFhJDabw/4cFd29
hvElJpAfRiH58u4W/K49oG9MqE/+x7XqUBjThS2eumuKyLy81ANDmX4a/hmKWE5b
Wb2ZyHwz8Q0Y7v42rw9RfttbrYUyZih6Qw/3cbwagUIQhe+Ipr+P/QTID7SunhsY
re+dKkmhHv8OEgIgIFcRz7H1FyOwco8LNxFqW6L2Ct0mhnuEQxDAcTDnZQ745iJY
UqhDZM91pNyml4/UvZkZ0flqr6a185XQqed76h1XFHU7Ue8luOogxBQRx7ZFvpEG
2sYVI4pbV7QrDipUQlxcd0J5P7jbRMG2LBj+RXfmrniFF6rw5ljy9C+W0VpDz8e/
1ugqPux19/wBrbSBsMc1VnrvjydJo6mB0TMetGy4gTuy97Uz8DB1koxdqNBq7qQ7
QWvoog9C8UkCWvNKvugFIWZEsAta+zf305NgadRTfs0KG5lgTq+SF+n2UDCLhGYm
o10XpIpBmAgj9sW+OQP/IwpLq0RYbfg4xrnOrWR/Qbhh94xPhjlgu5wT2L0fe8JA
gVaS1N+RTEA+iPBLBE/atQ3UUMBEt8Ml7R5/v57bCm95/1/f+9tjdjddFfPCGFdQ
EJ9CEuZ3EyczW5YmuihimoOriJ6ogoex+QT+QDxqu0GQPzzcSOYTjc+gTvxSic9U
jM8KfkGp1tFMUEpUUDy+sNKUcQvybAPQ0+5rRyc8fl5v6y3cyl07dViFW2bdRjGr
OheYniTczcOJPah/slWjjtKttgl3ROlkfnhAurQ+2TWhCqYAjHTWOCB4phk+Zm/V
V9g5x95bdRG8SOAgES0LHKBREALm/ryZMc/eUjTXIu1Kbo2dacCKDpG4NYMQkcjB
Td4Wf02CurpD7ElA3IXsGu+s752TlUgJW7pjowDWyAnrUunKyxdou9lWuc9rmzTp
LtVQH3GY46mL7WyN3md+qvRdWDU2aDeniFZE1o9504kLVo9MPNh/d0Fa/rb2jrpJ
TQuLPSHjBVbaVt5X1q8pzK8LvM860dhhgqnQEdmRz7xAAq5xBd9J9EeCbWwakZfF
N16K6smrONCO39jnakn0aSaS17E/9y91ar48ZvaKvptNzJC+YOKghI+z7tb6Jja4
Qbxgf8GVIFxaiL0tL/GDFR2bBtvJhgrZydBuYdh1BmwqdGKr2EW3Jr9sixCFmNPS
r/eYU/4NYgvpZjfcf7iu2rlI9fADbAzmAz6jBJXGNOipYibKBAXBxnqJiBHG1zuD
4Rhy/O5g83IZNHM66WZf+JvBOsIOTc2+IYaXYD97vpC2NBtgiCJILmRRWEWPv1Lk
GfMjv1BOwpcOmOU9xifqfA6ztiAw2byBUWjt+aQd3gCeyYBfiOCGAlUDM+tsYuUi
dEu4t9gVc3Iya/X9PS8TH3m2IHbaAlI+vjs+Lqij+oswov5PmhnqvChSGsaR6nT8
idcgB2kkZ63PvHuBdt4fIiFnzLVVuSi7p4C9e9E+Mf6/+4qyv+Ras5ZPRbdWurml
CzonjmRaEUsYJkmqRQlIrGCiWoIP4Yca0QfsjYeuHcup4IcM4jYNYMLWbUl7ECPj
gTzh+hmOrXuhes29uGicXRe54S536bEEGQeYdgM+jEAES7LZH35yjlWHJVuee09z
UJVmo85xDAKzzNuVv4sRa/Cl8VWkH1EJHYWyTQ5CnRjgjheQe+4BrG1PEXMQ792/
4S7xc/cfhabKJN9DCfqj5NIFfVJZgUBRoKYzg3SZYQhTahmzm4PLBYnNz60omEFg
gwrNEmYhOGukNG1VN03k71P+SNedQWorUXaGov5gK5arswvmEaM6JXGci2VwgYCF
pv0oQKzwxw11r0KJIiHK/vuQWAL6iaPKXTfRVOYqbl3xH1cKLO6P3lYG/t4RUMqN
vmgkE6sMhpaTW+B779qYXVTAE2UnmY6IA2cAcky3vSlJfmSk17fHhvuCEYyZORaF
z+Wa3HeaCfYaes+WzJo0E19CYoCuAKt7uy67JejfxOUKUTZLdCDlkPFrMNLCUFvg
DYHkSjQj6EM/ZirNj0gFQknupZ7BofsdpDPzb1xSIAb89u3PuRN8M0s62oZ47D3a
w8kI5LBMdCJWBjvpmmhSsSs/IrExFQ3XiemdVU0ngfZ6LMJWAO5uphTVOIpyFJ/w
5Qp/srKU5dMUnmA1mKoyocfVmtTMKMjd9xfnLxYCgwZJ2RpbQw3oplASoXeGMwGq
tamI/6n/o4MSA/SpNaz0daCpH9ZKuELJniUy8AIY+VhLJokhbMOmFxOBd1H6mcpS
g1xhaWW9N002xg6oJDPYS+KOJrEozpUGOOw+Okq7t7LsklTRGhVwtV5F+kW0QC4d
fZj5PQxzCBft4reC26IidXHewrwy5uhkagXmKs/PNtPiRcbE0Oyk9yBlbFfByZDj
PYOfSdmV7B7UPQ8511b84M+jnfuTWvByG6hp4Y+I15Qq/GjRR28I9U4cW+6SPUU0
Ge5uzqz8WOB8axdkODY/McbkGtkV81ZgNwtY2yPsVZLdAoBC8lVZQDGKD1r1zLm7
h98Q7Eu/9BaGtL9S1+wVAgQC+HAiTv/gm41XontKBa3LVZVX+X5OakZ4qF40hPEJ
6Nj+BHv3AbuIiUJzMWFAkMCxR+qgI1qvkxQlK7d+bRhA2Usfh549Qwswqu2dX0b6
vw2EdAslXmUW1NPKc7vSMO2g0Pac0TE5xT4XRHZIthgkN0F36/i01RsM207nG/vP
REmS6NYixxt681uxCLo+bYiu3YJDdjmlvD64TDjtagpyzVZV0mc2bs13ql8hFdcz
k2K9jqJLrb/pdmI7KIDUAKYunfmpCezDfw4AtbMK3b1383Osb56mfY2aK9Ywgvhe
6ixtOoCmDmuhcOBKAtVGuGprVUNoReNTVsJbRO4GFx9Xtsdk/bhNcVMRVoqLvTbn
64zaOxk+LIdvhTa+GN4gwdNNIUeSRWJYNntHONG0raTkG0P3x/J4Qv4gPaNLGp0m
7JNpQfiwpsQxnEe2Nk9j3yZ6ChDpTuLgoXazYWt5I5CboNoeu40uwXPAkQLgpc8Q
48xuIw6zEz5Oge+JjRBq3xGmQ4sHD9W5pjItOtgOagziKvi6ZHjl2O4ncEgmvypv
0cvaV+zqlFgPt96/P6QDG3CbuuOgPg9FxnQjBPFHYmZZn+ooDJz70Tk2wwT/JI+p
qDHdcmQnBp0Ag1hK0fI/eJNE2ipAxSgRyVOPKE4iHOJkoatE/HJ7MZtQ82b9wPtQ
LUOuxhv1AlbxwjuW+iIO7/spL11V51NJRzFvbqW4dJufx81sXIwa07eXH2Suhwnp
zs0ADWuSLXo0yVtMC9Eq/Kk9qqGtLi/E3YBhOCLtsgfUV+JhAiLQ+M6GmnXBc5Tk
TJUJAf2OTi1TPQ6Mrl7uHxIVhL0atGWZjdYxKN6RTkchlutRdZ+keXpDNXWzULQM
2gUUNylmP02bExnNZjOW+CDqSXEOpWD81boc9ND/ZWGp2rT4X+CtSpaLeKn/7PeY
wXKo0EIy2cdGpE25yFfku3GTqqIkARrLNj+HEgNjxi/NpwarnOjiGO0i7q5EdkCY
YCx7p2QCES/IobSKq5UHKW1ztMpOMnI0sWA8VhPEeUDKOg6m0uTnQRyaU2GF5KhV
DG8doVD8rGpKzD46i1rAAK1EO4KtlK/IEmRdWCEL247Q5akElIT+sF0CKGybJLM7
B14m7YsLxP4HbaYroKr03HKamVT2W2yMX9BzSRBURcQ6PpLNsvqrI5WiQz94joyG
9r24BuOc0OQDI5JESPyTl/x2VIjnJqP0TMcfkWA1ayGJYQ+M4dnNpXz5yAIZ5M3e
J8xP+VtPcrOEDu401QamZgPfSzH+WG49AlpxXZ0DNmYXCKDLJ+Pe34Kp+5u7abR8
FH0HS6Oz3/DWZxGQITkfcW9JvFgmUzr0L4p82RzBPZDzLd38kFs6+ovU+6WFuePj
I59T4g4+Ugc6d6zfovqXNyDzqmQ2E67CbzuIzIBxgf96gW6m1cZUkybGZQheWyli
LIkzn/HvNAtxPS78oq3vGu7wOaOGtNylVk3O8ihz3DkNQl3R4tjgsHgD9zXnl3lJ
aZ3V8bBxy7wbFk/XXlRHFh9eU3Lj33uJ3ZgGWM4y7TeFIr+dVx07oh5xjulCBuE3
Bg4Vv5k4uqIr7zGcpZ2BxaagMpWYJif97DmBDp6F1+ZrOdV2A2jd4LI9LAavWBZZ
KfWghXMfmX9Z/Em0+2H7EUtTAnvYzWy9MTweatVG/JNRe/vdMgOT15KyezzFm67e
kv1V3eYqpQajh0aqnqy+S5DKTbjJWwdG7kdl+55sJIPq8p1bXRFuy9bYIIoprKEA
K7IHWvOc1ezGW9RtLIDgZslkVOjKr/ivSWNqozZhH6UfvvTXrlB8Ucdfi0/NNX5o
vlY2RtnvyZVOSLGAdGaf6RZUkpM8mRLDsIiSCaorOit741B1Mht4lMjjSQhJxGVJ
WgK19KLfSknZTHKQNqPt0pAhr9+gx+IAiq88KIp5YjejG40uOzK7sw8HmUyVmhIY
buKMpE/q+lf3soax2zlIXlNIQe70G/sGS/Rx9DiCWVgYlJ5jAx6yDElMfwETJKi7
E/+FeRXFc4NNRFL3k9juWRpgD8+HihFmzQLjDOxL07+9mSFQbMEXnaW8wBKJ6jqo
uiseaOP8aIQ55jrH7uNPtMjgiLx70n9HppmzHqAR1g7j9dMpMT67KAWFLBkazc9K
JsUp3pwGuMHOFy4VINv5mwcdmjMZ2kYYAKaP0hSQ595RhEZFhkRTe7ABhxnqZJjA
oq8pma1GESR74Wd5kiJj0nBw3JVdRftQPk1Q+Ad/+2X/O1G6Li9OnejENrtY+WvI
Occ1xRnzKsAuPWmknTGaxZtZeLw/CfPug61K1jJPlQJ8bQfF94NaVc3BmIb8W16I
rAsa8tf/GFLCAUqcL+KjKy7BeygeoAb2KB0DUBe4LC8vM8X/6hPSnp/7SQ7Mq8l0
UEUYfwaVUHMxMY8JEM12xoLln7pFpoRFoO/fQOHHh1s9ZSW+zIukWIKPyFeGRg/g
EdBHFuO/i1GKlSoluOUuW4T+9crNb6J29IM1gy/0dGRz1Pc0TOkB2DTtd2N6Cd3s
4/G0m6YPn9ZRKq++EF4SqzQn2XEgaOIUwk3EiEcWp+Ws+4XkYcroktM91+UHTYU/
4sYzLJbHW6l1sWaynimRTatnPWJNF8LDmKO41vXKCXgID4Jz1EJggPMPo/9pgRnU
slMR15euR/f/tR3YhIDicvo+mfHZ2PoAlvWu26NHRPQ1BbvHTKfJEPLvmOLSedx+
y7taPSkVhEwqTKoIw+3RzVrQ/nZ51goYz4rt0y4wSXZ6COvetifB10in6PzROQ5b
8B5H/GoX2mIOdNYdlPmFb8/wQ+BYQrRg5WlBWKJs78w218D99vEGFe7iIEFb/bvF
omkcxJ5rO9hi6X7eVYY9e04e6I0+gezmo3ZQOwtPIpynNgcsUPMnPrIQq6fQhLoJ
/q4as1JmAmrW95YJK9C8XOg2ldrbsAZVAFa8Nzhy9czasBQKESytAz2bx/8fS8oV
hsBpXF2wPzgmgcAzzi5i9pY9fWT4bs4D0OvLOjD94a+9PXHFa8w400dfZ5eSpZXE
7yh1RNXXOhPFQ9bqyWhVJAh97ruCJqHfxne5b8feJEHXr/b+TvMEoe9+rWT4pvSQ
yKos5tuE5wZgARbn6r5EbxHVYlBI+KHv3LloYfpyOreGkn0t5YX8msw3D568WyFy
kNOVDcRQCu3jvXEnJGeItIImSVfqwF2F6pwMMNLAlc8lDI6DNvvAqh/5O16VVYx9
f2vO5g5/tT2ExKi2Jn9RI63TVLjH8Owldt0pxElaqt467U0hAnqMBG5FVmFb7wCE
S6IXTT3uOA/6FU4Y6kx95VI6uFv/WNbP+sDboEUtmIb/f3WuBVcz4ovCOoIxIXNA
HT16EKLQt9v0CBr48eA11pLYm9LdlXkL7+QwC1Opx6k2n/y+yeGkajEzgiU+Kywl
vTJ1SrdTZqmJlCpjjJbCMIDMyf7Y1cMRyH3GUFRzbU4BCcbppfiWzEHOIIJjME/R
ZiMioGo/pdr4/NT+xduNfx77PFmvUyAfDGcbs3cL2A1EK6XKSXR/0zfmDcSZLTyI
Auo1D2HvLD3F8JCB4nlXc+W+vc9AhWSClpXYpa2Fa1oke7D7ycHpLJoMnxOq1nLo
d+Poy6awDxo3WLIpAGImwggUNSOAxl/m6FBH8vmzOauzIaLBSp0aQwATD1qYQ0WY
UvFcwGn+URogwVFpegT3lk7+B52LqcXSRVRlgbg9LOrnT5Cdl1k+qe2RC/qXhcIr
aMToWkOSzFjQPtdZR3TmnjSaXSW095ESUnsSnCn21FrUdsY+hqBu3iMqguJhvZ7t
fl/aWp3oi3tBKt/G4yPolET6K1hjqcAunUYIVfcDIjPsdYvRw1E/QYMgHZn89k99
6k/KQn4mcnHIJWFFZqR5cHCZqTqRbd85n6zX/ZMKp8zBavm0xGKdv4DaYSRAFOPo
MZS4KhNIagRAhoECRQAw+XSNMrDAB2azSM6uxDkMjpwnG5WYRqk2U6DcmT7ds8v4
5ExyaJLCvUDtNXjf02NT3VQbmh2OFE9+eHXcYZcKqF6l9DpcOio1cSuO62eInciB
icdt4uBnGSEO3yZjmsZKBOX251dg0M7Xuq9qFG65ki7hCjaz1zmjc2ieuOOo4FTC
IltliEe0pw38kG7D7fwSclwEhi8WvAPUKpd8XXhpI2ViQyiFTaqzpVAXQs9gWy9w
FoauysLmWPIuOsHntwQU6Pfl1oxz+qv5yspEmdvPHvSPTtowvGRMq1tXg7qdOd9y
iUXyyxcnVjhTiTZi0vV1TLe1USBqz5ih4Pk/RDzPlPQPUUA/cLzT/iv860/pzCt2
GU1Y/Fey7EChE2cCc8hkptCRFfbPMsPvInopMWfkv4R9tGSgMlAIHnn8CZlChwD3
HaqG2z1VikjrQFt6bg3zLrOnoPXWKVGljbwLer7xFrT+xfbtXxKyrEI9KwMUJxK0
15FDo6mRhjTKJr7bYKiMLXlzvzH7YXtN4IIv/osd0ZEx83jHKpfGxYohsSbux2xL
jy/nMRxHz/JOmDQ//LJrDATuHmITxk9zs06MWCgZsPIPCXan2C9MRqFBUERNIS4k
3sjvpq007l/Wtx2iMvKI5FbOqKzBQkVK2t31VnxIz+tiXWXfQCgbq6GeDq2ii1Ir
+Jl45gZULs7zXHxko2gYeH4H7SbfL/z+NfCNMEB+eQOd/cNuBdHHkgP43f5vPjES
hvaK1wt3bO59bpEs31+mXVSDe/u/062NwDdh8k4KDq1CFFezvEIZ6RZgjezHIn1a
N07GFw6PAu749dsMgNKjFYlOjaXdW2Leu8nCaM/yOLMJSmbTA2neDiU8VKPGQBE7
rTKKz2v2HCfQgppNgPdKMz26cG+igbD2h+ffwjccDl4Hj/7MWqRVVwhwjFxCX2BN
RZ53BJaiUUoWBwOPX+FWpkwEVS8DpMrvDWF3PKWDqcO1yQOgaiWsjDxFV/JHp/1e
fGJD5v9ZP7xqr4OGaDyQSfUJ3h9xcBX8Upoz3XblzIPeqXPYeJ/jjc+6RVlRJgkn
hH3T2NKfv7uep3gSB48WnI6xY9iTkIR43aRR6cPSWMS/LKB6Qaeg976LHQdXZOuD
3piJumr0FW4/HMCF0DxMiX8FfqwYO04TD6a0q6kNES/zUaQCVwFuhXJ7U0AXv0io
9YOA50sZIpC3YQah8SCOLwRhzZFxsgXOUQJzKh/DW0IJqLfc+kEmd1HlkMoKikMP
9C0X0HXDKav9H6QpDn49so8S0zd1cjfLH2XsCr/Nc3Ns+U+sXQY0GtINR54esoXS
o0JtcANltSM5mQTaxTBcWnEX40jzdYnnKuE8+UAk2ejsXQ/LH1JR9lGuc0NPJOr1
LDb5IKgPbTGgRcoBs/1trBSiN57CZ1ZXC/16/dMoriyhRL95lEQX8M6PdICJcigb
cxIKXWK2D3KgZ61wQyPT/DzWJFdVSSiRBjmW2n8JW5fBewpY6pMGb3wp7546wDzu
5xSDIoCdMnKyPu14aCVZ+7vgjFbxv2KechPrGTr7D8LLhGnz/ZlNcGdojNrpa+Bo
5hhtO5TpQExeudO8dboBBiaQSzDEf1CYVy7GNjdYBICEzybUTUt+xaUiplNfPRqK
dN9mqDiLZhQl8JfbYAJo5iQFAbzwxc5sLl+jjQuDrJOXn39MYkxvj04afkXV0AHi
6iKPxcs9FqHDrlLUTO+oCu6pbVZ1Q/vyupJHaORQDGk0sKADjO3DZNr2x0WXwsie
7glrmCC2Sl8HUmsmG7IhsBpvnMo+GXOEcScHdBq1+PkhIA0y9gmT/ucjVZsMT6sf
5Zj4oSLsmfBR1CMsfwVkidKQ/3v6pAVlU8z7O28Jcagks4sZW0iWKEB0ljwBiaxj
Sbjate+CuVeRXKjj7KcZp2W0raeet+dLEvPLUtXdS5BJ8/xpGLouQAlAuGZ85YbG
8xKTrtKD6AXtF8+rjJwWVFIYkgqs3SZGX8iOCkoN6W2A3Lcf0qHDB3aHBNG3yTWe
NYQ+gUSBLI1zJdyPnrqSRVOsrRgrXwb/TVg7/G8Sib1UwKLtaTE+XjmzsEmqYWwV
NkGs5bBHjXQTkp3MuzhBV+tR6bZCIhx88tyY1y4Urc3miS1bdVp6GqxZanFIiHYm
LwYdRI2qZ8AwKXP2C5q47IMMLBvNGYU1befQqqF4pJ9rEnRzXqCPRvdExBiKcuPH
GXgEuTdPBbcjkz44ne3kWC80E39EODscFHx5XcDrjDlklH6UacubmuEAoJwUtmfF
g9LoA6ZpS0DjTK1xRZ1JwLvawaLDu+8+t82mAGu0qGEuSU98/TQqAu4jivFmD1Zz
za4Y4Tgrvd11t7dqYkQe4IbTfS/hBbSrpKkp1l/wDlYd3wWsPsCKSDZcvrE8ksjO
gtcCLOx8ynHdxvFonPhIcL37Zt8TWGdXZ7uhj9r9xSI5tKoEAXyj2DmBpOjfwZBo
pu4xWp2QYvVuJDUokcy7fl0FECrknApmSqVysz8aMf0Ubawb6+7GSGT/xaQWrw/F
XcXZMtpZAustEoJWHQ1IA7PvOVoKqcN+GT3lBS/ZyWVvDngYqZ4KnsaGwjeYbSdb
nBufGH+hJyQP/P4OXs1WXrULcCxm8yyAfhWR/1RizFzl1LVGtFeTVd56kuG5/ApS
TEM58oc97GUk5+dVew0GOvi2pcjXoQNb9JhD6a3d0wnFtZZg53bluAVJDtUNt3PN
J7loU9QRGZx/YEjnP1AYh3nr0EQeGC17IJmAUjCLW8qAxOqPd7mAlsSnac7bu9bO
J5tHXWw6ETqWLPAajbTGIWTXI+lZy9R/mHPayTN2c0cdJwJYRJWi5lVNdmQaY1E9
1A60aWpk2MEjgFxrHTbPNXRMLioRlyL0RgIXKWVS/1fuX7y3lavMP2cw669hFV+C
GLqJnsT0rdX+Cg4q7rJmyrN3UsZCNPSQC5za0xdm395FspPQXKhBGqPaynA5LSzn
p/kTa2CWq2owzf2bvtU+Lhg5T5du6mLzft/yw74yhHEPG5XYkJoeR3eOgFqUCDzU
8aFoJmHLSMCv1Rh2uQUU90v644zsDStKZXv31uCht52PrpOsOY2POR6vrDfBojEK
cVNqs1+JKMxFasXqG9NJMh6W5H86scChOVImfgwg4SaIuWwHKk416KO3JFbLR6YX
V/dPL20ZltgYfjX/GRsKj3nQWZwMnhS2hbJje/im2aKlEPk59m3T6NJXAdd8aorT
BgrRBQV+5JK3z7QjlZUWE/JJxJWPlCJ3yj8/Ki6oWK7aVSwNk7bCZx5NmcckoQiT
SbO0Nk+bTDdif9oo9M/W4AgfavOW/FDqjZ5PXGu2gDVT6CqrOGSL2yrJtBfshAI9
tJzsbtexWqjMR0imTCFV09maf1Eab/toDl4l5ZqMTJUKYiFWgPNHeBJBVovD0+e5
8TURZsz0t55ypqDD9HRwp4YLItJ5ZRclarPs26stES7AXgBbOblpKpc4cH95Pypp
0rb1pzLBOgFIaCEnLI55JV8ClSmSLKtzkCFkj1rDcgNZJYCZgmcszvzKWRKZu0lq
QnZtweVncibUfmCkYwVy59p6A8urOWwoQ7o+3mXcQOOYxmx6f7AoUZcXS6zvJExD
lqCP0GRuRL0HiO3H6ToAi43n49Lb7PTke4d/21Ye3o7Jzm3Kf5fMjTwUseJGz7Kg
h+2iGO2L7bJq5gX+GU8NhRYSdMWoi7A1CsGpOSRaIvaM5JlPQ1T+/5EUj36XBTj0
MyEo1LSKrhn6qctwxGyy0MDryLAecIJPZPsFD7VkhvbZ1K6ir4oFqiqhIWWYZM6R
HXkdrh4c/C9Aj4b9mRAJ7DkxnAiFPJXkeekVqbxfpTzqV1Q+mwQ5h4j4XDS0x/re
mQR4etazrgoJfUVJJ3zJfOFKqbmL3NYosOID7ziUnFSr23LmGvU9BPpkvr7XqBGT
l3se6TI3NjUBTb5QJdWxupuG9FifVJ2TmWK6ZcdAdeg3z19Jd5SV4C+znN1S7oJg
QjujRP6ls3GBQ3KD/OOIvIQLbiUGWbAPkUd5wP8FyI7oAAyA1wzFxjXoxxYgUSo/
LcadTdyE5ooKQpec3WSGaoQNhUXTEfSVQ9YYLO+CRMtk48rSRysA0KSKiiWHWHnG
DyidmTQrRIV6SEIhtJ+Fz1RU0LVKtGOC+m2aeYTd8T/auFSR9JI8b6qDnTbl17YO
VGc2jMPD5vz/Y8BGPLrgZwC8xqejZxacrlz+z0TQSKtqLqu46Qq60L52MYqVztJt
2l/iTTWr1JoSYbwwKiGA4ZrMDMCXU59qKCrjSn2Ac1Ta4JP19ZTTZWRYdCMMEBYx
UPxrkfb4herM+tr6Kb+Hkzeugb0lYSoih23VyXkWj8MOQ18ldSnXb1vD8dq8juZs
4ivXz6u3UE8+5poFz5jkX2kCcnD8I7Kc4oOOctJVhjRrMQ/1eImJNLBht/z7R1TU
7c+j1c/WIgYJ2myKDmGfk0Umd7XjCFx9unnbJW2AXFICzzX2YusmHAf/FsF4+av1
2k4xXd/hR+O7Q6TyWCSvi6whQr4pcaMXYMoP6Q1SCzXz/AIwJL3WMjbzQFq0NmHA
hJs+Qm9Xl10zM3V9Xc0TkNVpQ5/mRp4MWxvNhLHLI7SfX4tCaDCXjZXr5rrF04Cp
bxl9kUALnq58JUDmvykMB18k3mxtZdTvKMJCLyjAw/j//lTmJ91B+qMoVbKTc9QU
rAR4SqTOGKYz8VXOpBHVH09S/VRzapVJTefoEv/wWNDh2kzyrbl3SWgaYUHWJPeD
xVv0sbjod7CPmkwaLwL9XewxyjCFVZXEHxiz1k5IC17F6gCG5GMQN3kBRGLJtTIJ
QVWIUU9Fn8aj0b3r88LuDwG4lsB6Q6upvT9R+aRTRr3TIOQ3jSkqhcQDgdOXYkDW
5J+9wd6vxoat/TPYlY7L2QkecC2l0WYHzZbg75e66f88BgJeTGyT1GFO5SporAMo
PZNmerUPH1lLNw8viOKFVR5guCNKjvEAREZ5CRgidOvhwEQTi1m64Hn6ffV3/OFG
nswVcZ2HSyIYQk+Z/GFRb/vxELtnjWKqZv6udt1w0MPnEWzpKhAeVxHnYK67gEn1
zoId/i0XkRnpWKv7E1qJr2cGn0vdGCvWUKh4T4RIySpraYeBVzSx4Je9oBOIxE9Z
MXDtMjI5gwW2Fq2+rizroP6Rzp1VBVofvOA8Y9lOE0aKnBO7TP63J0ri9wZdqGuK
8CBpzjE/cQqBInP+0XxsBbNZ1EDCt33lclXsBX+f5juagsI3yOZP70S84UaNx8w5
HKuaPbDttbK6nyNEZm7DtyFb46NBA7f9fZJ6arBJj4z4qhrktiIJkdYOCVLUPWye
zy0bgvA9rmkiaAsM1Yw2O3+8wpL8dVIzg656GAOMnpNDO/DHwbMabdGI5PQJtDe4
TuWk+rs48Rjv1Nkg695K6MXDgjC759A0k3a4oVxKNnYtPktVi0FUkx17Ym0gT2/Z
dW3tIbKh3oT6FhOHQZr8UO0mNATmlpb3TYrZeKaVkOEgpc9vZ6NzZCwQX+k+DMpQ
LqdX+deha6B7auXVJ2+TbbLqQfp2seP96k6P3mAmYUlRKMMT5Y7ISQejuUFO9eq9
4e1QUVwUW0IuJJAd0fA/iADbO9wTSGxYqVu3xq0l1k8Dx9AFO4wmS3O14ogmcmRo
yYGV2bM1l6Gke3bTEU+WU40Fm2RI5oCOYK48OdQg8WZAct14zvAVRJ+p3WyoomRN
OpqUxtUjbewOGFnb8Qt+1oGiq4hYU6O3YUSEkMEqArkJOb5lqFKA1AfkDpzNAtd7
RRVnqyKQ6ZQ3jo90R0RUrLeuCnZOKz6oFCGYUViLAcfkWhWNPug6NieDhaUS34JC
6pGsJmOvFSOp74+bV6p4qGlEv4wgh6bGxTBzrOTs1v31Ki//nv08ZZ62RpsmElWB
dmtV8FLMQa89nWNqZag4RzubYK3LMiLz61YBnIDjunRhY4Ihcq06gfZsWW/BM8Fc
5wk1zUyzVgJF5d1/glX0YriSQhI2iRXJmbRpydRx/TfIaQfrty41bA/wbVuniH6j
wvoSV8bc+wYMVMdGHQVeMghN8E/38e3aMsaT/OJ36ByZXqpp78AS3Qmy05Xk+uVX
u+Wz264wTXv01AC2uhfLA2lEhLtMQ3QMel8+bdR1Xs0QtiR94//+fzswLIWpk8OZ
xkKAkieFbdDogaLLGCP82XHYzJsI3/ih1/d5mz+UUcgqbCcLqYfcBOAXGNXtRjWh
LDT9T+6IYhhyYM7nGzRcqYaBir/x+mzNqt8W44/zteShmlmDWZIrTcgieUWD+gFU
5gt9MGPkuLFIBIudV0NJQLiJZqvydDjjFjy2E2NrQRBWij3vA5yTXITdO7js1Fdq
h/yb9VeKMOtIx6kT1kBuBZLD2S7Mym6kvWI3NMmXY/6BiSSl4tlCRPrm2Dzp/BSI
JOYShh0u+u4sQVES5akrhxhHfdz1vYv+wnOOzQ/C/FF2QD7Poy7a8LtLtwJwZX2g
9r0MkSSZppZWOVaLFFywd18E7RBwaM2izbHVVQI2UiBqeqfFA1DFk8NYg/96MIAf
phGhZdMlKyxSedIQ7CDAKSPwkoIimgvMpoYCpIvwjcjcL96WTIjN8SWtZy4Qw5nL
K02DBxKUah8Ka+JnneKQZgXW7TNKHmFj1sOm/eOFZdY7P4K+/x82wloMRyeLmG5l
D929i7LPA0ddia3WQcB3bjkVGs8+s33W12OdgQwi0AjHaAVmPHlhG26rN9oUXk+G
/AAp6Z0NMCh5AagNSToec48rbuYKG3lDQUGHlM0a17ez2ZVzQji+Wa63YodVAXXD
q1KXX5AQ8tN0y6FStWrxiLKuW+PHZR7pAWJO89yhQHjSneeo/SlMDGHyhStEHK6y
6rQotj/FdyalapucxPHGlMrq+ia4Y1Q6ggG84e3L9TdosYOr47PCgeph19+Tw8t/
yv1xXtuhLNmDbdfxd28OsU3R+jSlYCufXWNo0Nd8QGklhVCIiueZyCrXA3t5vqdr
oflZcE+GmJUjuPXTqfHtb/1Da1B2JE0B3VOY6RymO6xy/gGdrQeckB09xAhBtUIh
3gJKoeyFzWO0pxbqF7rtX+lDhiJ0cUj3RW4YKoWcvfHcCJAXoUGSKNhXW4vvCNxg
thLFMHXJmB833FAyAoteQfwqTd2eHUUiCnVwsGA1fI40UHoPYCQ3hptOhRUKsNB+
5srSqGiYPYVucrSyc/o0PajAesvhHjnUcs9rotObqxgDDZEF/MFov9AFrCG+4/Fk
RuDYsTx67ymdYPOmflsa75I9bCAY2ZIRu50XmGcqjbsX6GmiTE8Qm1MGZBdR2q+p
BMHU34E/NSbvcEuoljfyXIvs7qVbRGQbqTG5AC5uUnOZ1TonHU7uxbgV0Y367bGQ
poBnNboRygQm94ExbKLFqA4fP0pnQMMA4VNBjpiCWwDBTQZBKwlx5zKXr8UhXV2u
v5+/nOgyfUHFkCWsUB9OkpuYQIG7Jy3rCLEjiHzpH586mCEMOiUlUfY6HM10m2zq
vcmG2YebFZerA/vzdqZb/nKaWHyRppCzIsiTl57TQNIjnL4ZBgA5sblKbD5RQUdz
ymOzXLzQElJOl1jN9Ycza3ceod9NCY6omFhSxD2XHWILc/SEuhUH78njkGcZCSeJ
rzu11tW5/bhdPQTdPHGVsHPl6h/EuSRigonHpANBAFdf6YuL/NLm+2Fxltt1DcMN
WZG2xTt+YN8qTgVjE9HFY2N3713H8H55b70MN/CenzU4z+WZomUCa0C1sUOQCKDn
gZcGCNA3O2SvJxTGn+ylOWP8Vrjbq/IdnHNemqmY/nFLMlvtVni/lSkRgZYcW0jB
T1EqhodxeFHHjRhFtlsxTwvPj3TSOPcPWv13Vn7OIGKSdZR36Q+hoiSb0DTTD1p5
LqkrUcdjhLPzxoAAit3mpCCVdpEKWkvdl4n8vATu8msH5ssmV2Nae9SB4YsQK8/+
zdHx1xitloF9ILnAHscG0HzN2xFzIlimhMrzvADQywSjUFZgdCEqzw+aVlP0pqj4
KCrsc0kBCVPTlo+JrGebvmHKkYj1NVafzCD0qvtx0IeEvYrrNm0GXd+kNhxtFZ2+
FGU4og/IBicjff/gqpBYuNUGExWYxc/gcqYIUNymEA+e1DwuDHZCX1LaDSlBmJ65
R/3YNePp7Ta1JB7ziy0Ef/ZWGvRbfHY5fUnMh3VTBBcoE58MI3pI3c9NTSwnNyMR
zlSAkfUEgJHYxNi8G+LOzEkhFOo0BKilN+uTxyqcz+x1tjyqNCjmDD0uTnXQ405b
U23QtkH37rD6rMQ95Ivs6mi7momwASL0WElTA+fzqv7B34jW5Jxx1HxzZ1/UwcES
JYT1AhrRYuO0yt/dPn2xippAYdVv9ngS5sST37bSzuHtILO43fWIQIMLXibPZUE+
k6Y89ErGL/SCKRi9OGG6c5BNITCh14OnLRBHtO6IJYC/M1/ujj6Wmgd4r0eH758s
Csg+8/FwA7VS4jI686mKY9i8Ro4xdUoqn41JhHnF3DgS1Tmn1aw+C+FCwX89WxZD
dfGxbYx3HoDIsSA8Qr1znFVjJfiOPOBAzkdhnr2kjXveKeCE9ntvxjpjHQRLL8vA
ap9lmB53Fctu/N0sfB+eOo49ah4fyY+4YOP+MmoYgwLlgFACtLWGXBxnALTy3oWU
5gBBQqLtRYhBo9Trjyi43Z/690bqMAqKhS0850n+uwlNsI+d779jLndCv/3n3/Me
4NE7hUdjjBMtLhz6PZh/tRHx0+Jb0GsyYgjiaHe2fqPFLzr3ND6e7Snfwl5hCabV
GgDdB8RuRjFKX+ISuSU8NtXV216DmcgP7Ds02xfrrVX3sH8FXXceA0RYLcCokkDK
Hy0jFzcRHVrRqYURxCSmK0JrhOzUAz0dRKn8qgrnFjd6KzoWbcG8CQsi8koJ8be+
wVzdPmEqATNdl7m8F+Zhl9nhL0I7JHh1eAHOCg50BJ3x9/8UfLKp6NhETV3hQRqi
NA5PE1XhfktE9UuG9t7Bsb0uWOxcB/erX4tQ5G/abYygO4S6BLC1U13uBygue1TN
OYfFjD6zUdOHI4wFn8uHpAMJiZ3NG7Lmsv5XC4jJ5mXoddfdEnmOmuZMuCqVQ1aA
0o3Ik0JQVMwvUnKBuvmFdsuKNBwOrtaHzZcfW30EYEWB0pnZDiFByjZRkHw3nlDL
VmFvBHBWP5Xqek57zoRMw/EOORFbhM5xmgI/Ap0RkxDJcrWrlXTpSwhUxKIgTjJo
Q1wBfxhMbDAQBSED9cKVB41etnLmqV8sJq21nSuwknfwxu+HL8DGqFc4TOTEldut
6Pqb5Ame7nMOaF9jUaHVUo9tcm4b7LkKI4XxC2v1X7bRAVsxBy9PS8bG36zvpqE4
F63uXIvcZgtGvV+I694IA5whMqU+Dp38FQ7ho38F4yF9P7fwy1AzHvRQ/7sT94Tv
pNxFIHbPfjic0h4WVgz9+xvsxvyQ3CGPKvt0wlUoSCXW4b903y9OXpmDQ9s7K4A+
PeJTr/GdAamNc8aY2i/g0Tc2yXAagSMjPe7LRX19WbsYlToM33WS+jN8NTVDUEip
U++jj3+YMBgh7JU7bXOmTzhcXSExerqGSyw4cUwdolF/BKROoa4bMKPx3e9ko+yp
Px+alefEJFskvCTf0p99yV6xT6pCKIlIukNL3o+KIgKvK81aAoIXmj4GCcZBMVdo
XruuKTYVOYd5TMgraZjbOLIS5anWmsZQLVVSjMBmna2dRyzTBaUHVtJ0Kt31D4G+
Kml+Z8P47EanwRTJJ/SyVNFcDz/FX8wauSGCLXYs/9drnthvUpyACfgLvE0WN7Xr
a4FLlvdZiXOelB7ybTsS19wdSXep+Vlo8L7XdMUDPtM/gtCe8+kCIXLBHkkXGBos
+6ohdf6lwNnjF0CtZpdzUCvO+ljNePmNhAPgliCSekV+Yxq/Sjdeif6yGM/xAEg0
UZCMdqN9P+5zbjjSfIi6MrJSMEZ80ujuRQb17Cnt+4ApO3y/x5KAeDXO+RVD/M4Z
J/Aav84y2ICB0nLQA3gkMbSTRd/v4CttH9tgvUePWxpVWT400jfRpdXBKyMCyqPI
mtRGxLeL4PyP7MUW4BemlgcSpUqMSQfiZ6VWuVYxJHeVS3BlI1RB/TyIyfsTzKFS
eNRQpr9aTAPskEqwyFb2KPczQctuYaFaXAnCpVCi6jKm9usjcnIMdkkT+fgU73ZD
uX1i/QPTWs4qM94sOQI52mjEFMGmQZF1EWYE1i4FRNX/9WxL4egNU0U5eo58Xox7
dPjcK9r24NKo+w4+kRlXQMQ3X6nXPxkQYft0NKiF9gq2Mnum3WMdqKP1uVdFOhRr
ypxbR071M3wrSN2hF6nLvc7M0wpSl12dYv294Igso5IC0SVmPJiOTJldvMzzrcFU
mm+ZuLNWkJNoLKpZow+MzP4SjsJ+/b/EYPOQFPYivdMxeUzKzpsXzYLX9q6wJbNH
v5kXZEl0zddP4VcVlXsnLAYn8asDs2j9OsImaegvb6ujh+7pdeUzEi3HOYGQSFqc
pDxzNeDgzvsOByjeTwnkTyTxIqgNYo1sQEJ8on7Bezetti0QoOD3XhguMMaAXNZA
z6L77YRmDxL1pFyqurfQacqEOJKDVcUlsTpPhdnnpF0+1ZIfG2leLjqg2Bj2E1nq
Z3/yoVYDYPqMipbF/1ljKlnbG4PnDl6ujBQ/TaOqPi5rEon/llL4VrfU5avmX2Fu
noi4hz4QWa7StyneW1oRylV8yMKVcC+Qj/tvvumbvuPp2CvG/eithABReJmZKUVx
+UQ8ivl4kq3/4gipWJqaVFRVFo9qThLcRP4lbe96t1efjXI9u7lutcczKHPy7y/f
098GDZlGwiuFeTTg6ZACnOExq+5m7RtxKmkL+e1Q1gdmVQC8N6tqR08vmATHS56B
c7c1zWC4nXcvnVFSF/X8srXscNocpm8Ss4I/CBjRJEaKKsIgSkmmgLM0rqhJKYID
2Z7dMfEQU3fvzjshoATYpx+pbDZhe1ZBEsF3taq7Y2KRYOhicRKWqZx98t6xwWJm
L2GezIZshOb2xE19AqYPFRNvEVKOs+rluPlk3gEQHSias/8f18bQ63WqksN58l6t
uU9OSid6XB5EGvHEUuXQWol/sNtWZBOWqDwDeliWMholgBTH50Io8n6vpayhZWN+
mWxZYLOc+P7I4G1fuQMsX+quGhTbqav7+jNZH/xUnxWZEwJCjoAoB6rtl6b9s/E5
miyc3+dS0n858ZQs9eX5mpM3jDzuKE0oozqzcLn5DMl32hHwXy/Zt2D1WJZEOvfG
vWIxsMb4MRx747ytfChyaPXQNCSW4s8b+6uFwSHTQ89WRN3Q91jGqiX19bXF3QJC
3BPJ8oN3Zf10wAtXm/s6IOlOXtujnst00voDyTXg6lHl+pK68LNihcjUhj28R5A0
oelbHDZ2nNcvL1WeN31fvVJzGML86Mx/+5UXWUd9h/07PBFxubVszldzcHxZUr5o
yQeM53sFf1m3wWFcn7jxv8VZF/PoL3X/sfaD7+jW9Vr+bYHcKAvpf7nq47jjNIJ1
mB+8Xuvcy5y9MRsL5BE4DpUKx5HSm9Vy5YzQSWBArgANjh+buQA6YbasvN75dsGK
fIr6JbSXJeTBtt7jqi5wcY4vMOPQfC3Jkt9leegg5+iW/aLYggOo2CRFo9BfToi8
XaWoOHDPBQYp8BJRgzQnsQT4JKrY604QMR+Q8Ww/sDFQJPwMq/8GbXAC+aMiVMD7
I3k36nv8o7YleJdQLor7AmKqLwQY9EaT6OkDg/n1aJwnCB7yaz0niDZ0wrINdkcf
r58tl6CvnMHnyudpSZV93Nm5bTE6PjIFvcFF2HLIsJPmn2+pUzjnOP7pNxoHnV2f
nOpknOCWhf1beCQyozj9hA==
//pragma protect end_data_block
//pragma protect digest_block
xcO+BchTEug2jZ3RCPEvjS3TVn8=
//pragma protect end_digest_block
//pragma protect end_protected
     
`ifdef SVT_UVM_TECHNOLOGY
   typedef uvm_tlm_fifo#(`SVT_AXI_MASTER_TRANSACTION_TYPE) svt_axi_master_input_port_type;
`elsif SVT_OVM_TECHNOLOGY
   typedef tlm_fifo#(`SVT_AXI_MASTER_TRANSACTION_TYPE) svt_axi_master_input_port_type;
`elsif SVT_VMM_TECHNOLOGY
  typedef vmm_channel_typed#(svt_axi_master_transaction) svt_axi_master_transaction_channel;
  typedef vmm_channel_typed#(`SVT_AXI_MASTER_TRANSACTION_TYPE) svt_axi_master_input_port_type;
  `vmm_atomic_gen(svt_axi_master_transaction, "VMM (Atomic) Generator for svt_axi_master_transaction data objects")
  `vmm_scenario_gen(svt_axi_master_transaction, "VMM (Scenario) Generator for svt_axi_master_transaction data objects")
`endif 

`endif // GUARD_SVT_AXI_MASTER_TRANSACTION_SV
