
`ifndef GUARD_SVT_AXI_LP_CHECKER_SV
`define GUARD_SVT_AXI_LP_CHECKER_SV
/**
 * Class declaration of each of the error check stats instances using the 
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 * 
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */

`ifndef SVT_VMM_TECHNOLOGY
//vcs_lic_vip_protect
  `protected
H0?,J/0N70dc?_4\&2=cUY,-;:e<-?:^.aQ?B>==&/-8Z/G/5/&Z7(RA7@\U@:MY
>@)KJLE-YQ6;L[QdWEVTfD[8a.1LGd4N(dBIe1<;1C4\FSNQA==S;?D=E=L9_CRT
?&>+RfPI4CM2]0/\<aN@9B]eUG[C+LRERaH:[:R:0-/<PG:HICT4J4HS1:DBK2g/
T2WfW#N#D@/;CG2JS.6b#RBHT0U8(5LRRTT]\G>GPM@?Y\G>?0_M&R[;:,F;EMRe
g:R1;ZQNTf\F4b^MfF=V(26PYFe(]=;&ZMQQS?S]=A,6Y5&7&fX,?KBZ\\Ta1<T7
(dT#eTDL3FHM1ge4Ee8YROQ8)RScbJeaWR0^ZaD(;]\144P51PJ\4fBgW-@&a#&C
;IZ4N/B/acE1IQJSPW</+D[(d;fB>3A0)@.HQ^,N3#(Z\LJ<\2Vag0bdY)T?ZDM+
@dC/Ra@K;3L\<]LK\\:.8^7SbNI9TNOT>S[40F6^3\M20J38^FU)6,ZO<JMJ.BS[
:0>^,KbCg=;0f3N<VO8cVUPF(8_;(V#I2a)W2bJATX/5Ka:[ReF)SJ-8H93a@;M^
V]:61;VULbEA>R6#C>)6D=NO./K<](cUJZT^)?-^B\Y778=;Eb>,G[@#W)T[09YU
_Cg[OcX7+INc386EIUZ6&8K(d]/?NB7JJTcP/O4RA#6]R<B.[1&X8ZG@Z.8#KN]Y
@bHWW3&FNCJ12-+ZSK/=K?/?D_4#JaCL>gPO2F_PH;C5)E<dfNHd?:&cOMP8,;Uc
d#0N4D>QBe>W34d)PQ9E^S+D[FI+G0:<=W8eN0Q^e?E/IQ#AXc1=,Vd>8I4XF>/Z
bSB>AZ6@BB#TTFS--Nbf6Z]9?eBcKMP8CN(O_>XW^.CJ>JX\RXb0_NFe^aO_7L1a
S1Y^DCbDg@(>-1BH\<B=\8Uc:Y(eZfW&a08[Z.BNa-V/D_.;E/FR^/SUBg_GVd/4
[.E^&Y5d[.Wd92&WXCb<L3_/ENS?7-Lg6f-a#H+9SESXJWE=XD3RDc9WXQBJQK))
_.(\?BDE+UA&R()b//,,e[:R+fFZ=e.#Q@>/15fF(O;Y>5E\^HLYJI8<FUSRYR=^
,(\eE2<L]H[IG,e.3Ed-(2219_QR#+.\.HKTM,fWFK:INfcDV[(5ROBT_K^b,FPW
376-#5,98?a/GBZZUJS4HHcCEA=Ub()KO-^9_#?/E\>ebC[OV&N\D2^BE1:BBA2>
:Oab2?A;;,DTWb7EA[DTJ=2U0[VUYO-HZdQC>c/VDD2/=(MKMJ?(F]WgFUG1HA2H
(WB0FW-OF3Q>W.-ZBP_P0SZS>@Kea&IUaV1UD/Z<.e0G_HM0D>S,XMT#]WcK;U==
gS&/>0GI3P\;@Db4QF3aCYJWK)C>+YE_QJBBcT@<DXdE7>\9>A2Pd&.AP(P.[]N-
LE5J[36+W5?e/>\Fc1cLUT,SNIa>Y:W\KALQX_bL7.9AG<;W)M;63&aJ]dUO<]R@
NeV;@^,M4c4[<MZ-Y&Og8<,1UL>E9/0WT]XI_]J\c.47e?a):Tbfd_SUE^Cf,)6b
0a2<F[d^,-eBA;Tf/:@](.Q>276f5J;Z.W&&[H;OCYR<g.XWVIX<O/S18FMN/G9L
3LPb>I1;Nc_RH.a23=e<RAdc+Y@SWDN4POB2QB(Y^f[-[&3BE<e9<Tg0>Y1H9e+(
19fV>aYaP8UabZ?_aa,Q;A@(.V_>=F.;^F&f0Q5.FB.cSY[0FN]LU8B_W.D6+RD+
HN(XOCU@+b,DO@.M/]KRNFeC@(Wg4;)LGRL^FMW(AN<5KDCc53,U=-_36G+,OOQe
RM,b\G,2@(NR8Z_3BDO.89ZC@6J5X#T)CLC_6baXZeJ+U9\(ea[50M5K]17ZF)Wf
#e1?5GIXD,S92@VF;.Q0\,3J),2:<-#FX+W,=_56MW?)ZbLMeE/M7EPg-[QNKJee
QWCS\;VTKfJF00@KM#6JR=\+T+Ef\]/I7W-BFI0FK(U_XYb.F@GS<f\@LN?7/EA0
=;L(MeXfE:DU<2RX;#HE<95[d)>5/::\c@]be&ZYTROPR51c<KJ+7H.B)d-(XgGY
56bC2=T9WGJP\HET<f1Z<TUMV\\,Y9)DS73U6FR^,:^W5><(WQJX4,a>^H@Jd27Q
PQC6(+6a:4b(TFeNfb)JBRQ2RD0IN=dRb&dK9_+\J,@UB-H:5^V42=eDfdb>CYFI
X_QYKB)K^GQUZ@fQW8Xc-OA1]>J/PP.=A5.\7MOdFdC-PeZ-6AY<.Ag]5I@:=XUC
^Q>Z-LF4S54e(a)Oc5.K\E6OFKNNOTW912^5aLg1NdgHWdL:-7(7U+EYOA;=5J6>
Z-g^[S5/aI?B.BH]1I<@VAe2-</T8HJ@\@URB..c_9(d2)]bNJ&@/3.b:-3GbBOU
D#W;B?O_K>2C_cba6I@G&JKAA/Y3GV9BVbU,dI_d]X]c<>YY2YbC/[I-DW?84CfX
4^KDNX@BU^4,?9f5<WR52SL-U&PcGe6&4FN+44>g[3S]BKfXQfdQ;]&PZIC;fcHY
fW1)d2d_^_]2NP][5)6cDZVPMTQNT6?c3gc=#-Y6Z/RL(APcSERDB6AgIR:fQX/G
ZE9ZR.d6VS2UJ:)Va[PM,6:c_1dSOWaUVId0[,UXJD-K=JGOC9EI=J:U/R6;0#D3
OUEd6,EQ+YUXaR_6e-6B6f<N8VA;/K=57L_6_I_)<JO[:;V0eg=XfC4)-0_((^-6
L:=_cWT-F4P(/N+e)a\>;5Ya3U8Q+HRU@<P_:DeG&S9C;^<-P1#02##CU5.>(S.9
E2aB8>:S:P(O,c;Ie_2_5-+5<4G@N-Ff&D[LDFYJ5W_Y:(W8(d^Y&dbE_?eHLWJ@
12gWb6K#-ADV<FFf1\<I@;LRFdF9A@<91BH_?UF^N\T:6REP4Z?HM(a:6BcGgQ8I
>O;Qec4Q20DFD>=WZAXMA8X<.WV=W#JbHEM)8BL@^AU0Z5J(LNcS<:9OC8^@Yd.,
,XAO)_ZA:#[Q\63>I;+XD5XIfD53YUD3U1\Hb=E0McJ=YXEX\KFF03V>e5LKBS)4
:Z[<4Y?(V+L1K36VDa\Q[>JETQ7[AH_4P&VC:U>a.P@2L7\f>N9L<K>fdKV6Ab,A
?HJJDb-AS<-Q-ME>Rf\>:XFf?1\c-4=L?BTb\Ca_AER-VX\BD;10</>fO$
`endprotected

`endif

class svt_axi_lp_checker extends svt_err_check;
  local svt_axi_lp_port_configuration cfg;

`protected
8A0\EOJJ6T5PZaCdI6J6;MTP]a<DU/_/8I7c=6IGYe-GQO8Z[=3e))g)O54I@CY5
B86g#16#2KQP,$
`endprotected

  local string group_name = "";

  local string sub_group_name = "";

  /** String used in macros */
  local string macro_str = "";

  //--------------------------------------------------------------
  /** X/Z on the cactive signal */ 
  svt_err_check_stats signal_valid_cactive_check; 

  
  /** X/Z on the csysreq signal */ 
  svt_err_check_stats signal_valid_csysreq_check; 

  
  /** X/Z on the csysack signal */ 
  svt_err_check_stats signal_valid_csysack_check; 

  
  /** while entering into low power state, csysreq has gone low before cactive going low */ 
  svt_err_check_stats entry_to_lp_csysreq_before_cactive_check; 

  
  /** while entering into low power state, csysack has gone low before cactive going low */ 
  svt_err_check_stats entry_to_lp_csysack_before_cactive_check; 

  
  /** while entering into low power state, cactive has gone high without waiting for csysreq to go low */ 
  svt_err_check_stats entry_to_lp_cactive_stable_till_csysreq_check; 

  
  /** after cactive has gone low, timedout waiting for csysreq to go low */ 
  svt_err_check_stats entry_to_lp_csysreq_timeout_after_cactive_check; 

  
  /** after cactive has gone low, csysack has gone low before csysreq going low */ 
  svt_err_check_stats entry_to_lp_csysack_before_csysreq_check; 

  
  /** while entering into low power state, cactive has gone high without waiting for csysreq and csysack to go low */ 
  svt_err_check_stats entry_to_lp_cactive_stable_till_csysreq_csysack_check; 

  
  /** after csysreq has gone low, timedout waiting for csysack to go low */ 
  svt_err_check_stats entry_to_lp_csysack_timeout_after_csysreq_check; 

  
  /** csysreq has gone high without waiting for csysack to go low */ 
  svt_err_check_stats entry_to_lp_csysreq_stable_till_csysack_check; 

  
  /** while exiting from low power state, csysack has gone high before cactive/csysreq going high */ 
  svt_err_check_stats exit_from_lp_csysack_before_cactive_csysreq_check; 

  
  /** while exiting from low power state, cactive has gone low before the csysreq has gone high */ 
  svt_err_check_stats exit_from_lp_prp_cactive_stable_till_csysreq_check; 

  
  /** after cactive has gone high, timedout waiting for csysreq to go high */ 
  svt_err_check_stats exit_from_lp_prp_csysreq_timeout_after_cactive_check; 

  
  /** while exiting from low power state, csysack has gone high before the csysreq has gone high */ 
  svt_err_check_stats exit_from_lp_prp_csysack_before_csysreq_check; 

  
  /** while exiting from low power state, cactive has gone low before the csysreq, csysack have gone high */ 
  svt_err_check_stats exit_from_lp_prp_cactive_stable_till_csysreq_csysack_check; 

  
  /** after cactive, csysreq have gone high, timedout waiting for csysack to go high */ 
  svt_err_check_stats exit_from_lp_prp_csysack_timeout_after_csysreq_check; 

  
  /** while exiting from low power state, csysreq has gone low before the csysack has gone high */ 
  svt_err_check_stats exit_from_lp_prp_csysreq_stable_till_csysack_check; 

  
  /** while exiting from low power state, csysreq has gone low before the cactive has gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysreq_stable_till_cactive_check; 

  
  /** after csysreq has gone high, timedout waiting for cactive to go high */ 
  svt_err_check_stats exit_from_lp_ctrl_cactive_timeout_after_csysreq_check; 

  
  /** while exiting from low power state, csysack has gone high before the cactive has gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysack_before_cactive_check; 

  
  /** while exiting from low power state, cactive has gone low before the csysack has gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_cactive_stable_till_csysreq_csysack_check; 

  
  /** after cactive, csysreq have gone high, timedout waiting for csysack to go high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysack_timeout_after_cactive_check; 

  
  /** while exiting from low power state, csysreq has gone low before the cactive, csysack have gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysreq_stable_till_csysack_check; 

`ifdef SVT_UVM_TECHNOLOGY
  /** UVM report server passed in through the constructor */
  uvm_report_object reporter;
`elsif SVT_OVM_TECHNOLOGY
  /** OVM report server passed in through the constructor */
  ovm_report_object reporter;
`else
  /** VMM message service passed in through the constructor*/ 
  vmm_log  log;
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_lp_port_configuration cfg, uvm_report_object reporter, bit register_enable=1);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_lp_port_configuration cfg, ovm_report_object reporter, bit register_enable=1);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param log VMM log instance used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (string name, svt_axi_lp_port_configuration cfg, vmm_log log = null, bit register_enable=1);
`endif

  /** @cond PRIVATE */
  extern function void set_default_pass_effect(svt_err_check_stats::fail_effect_enum default_pass_effect);
  extern function void execute(svt_err_check_stats check_stats, bit test_pass, string fail_msg="",
                               svt_err_check_stats::fail_effect_enum fail_effect=svt_err_check_stats::ERROR);

  extern function void register_err_checks(bit en = 1'b1);

  /** @endcond */
endclass

//----------------------------------------------------------------
/**
AXI low power port monitor check description
*/

`protected
ZNK?VWL@1)XNMHG.^gEe>=/I/^XN^C)MOC6Y@dQJ-17T.1/X&BL,1)9UYS92NQN9
1b7Y3TXC1G[RW8^EL5MKdfP<P-]KNXKQ1EK-2=Ng;H9b;EY1[]c9B4YDN/fAVZb5
OeB.96]KD-W.+6eP7e?<P,eDg>TE1f/K^(T)b.Y,\+B_P==CIWQA=#0EXd69U1g^
^GB^6eP.Z09Fd.??Dc5-/7^)H,67<C=@RMN)U0F,#Y:Gd;61TM#8;&dd]1\#2JEN
a#Vb/<<gU;COa/&3?NLGZ=f>GJWda]Q8X<B9Q@,J8N6&Q6]6aP[6;-3eUe+;0<W5
AKI\c21#ZHIKKQVL4P;gW<SV2&IN1f.?dK,6BP>:_5@?VfM\OgKBIC#V0e2C/Z/N
XSRLMNZ8^K6T;.-W0NI2_@Q0A(_KHL-eCUAe0=1+/CU0A>SB2G/e)&fB#W12TQSI
J?S]TD@d(g.?DfgbE_BaMK+QESU(H-f/NK?#1\A,Y[:N+Qe2G#Qa4C(MBHcE6_1+
>>C#]Y@M,Ec1X?Q<RXFBHD</DHNQ3<\_E;[\=0PI+8T,deD-F=e#3&SS^DWR1BI;
C9(IS3Y[#U>\bJF>/#>56AF>:M4JeZd8R4??H^a;N(><8McC-JS[G;)3>E74AZ4^
9)92@RXO]aA/0\29A?g(aP_2g/5UaU)3#^TR]1eCN&C#_(HAeQ7a086M=O&6=+TD
N982H+^AZNH^<Lc1+d5IM=<?<EW#c)L655BO.<VCXLb+S6)+g3fc+_)TMK]:1<XA
E8Q1f#SQPcdZIJDP+5J=-S3X0;WZ93EVU1eZB74[IbR2OHX5=d#aZEOT)EFAT&,@
8_3+1MX0HAAX#1c0.L.OF3_+Q2e&eV-.CB.Xca(OcM@7c<^A7_]ac=R,MA8DdM8M
,UNcNHIKJ&?>_DF/_05NcfaA.6]J>KgZ20f3bO56A^#9N[34[K/)B;2/(JP.\)/G
NOO&]c+UG[>P8Xd]&Lb=gCeLbQ^X5]-F5LQK+W(O[&FH2.L91Z\Z7X_M45A8O1YF
8R<@CWZ_ZD/@34^/7F7e)U+1EZ(SZFE4\;9<V<K?[F.L\TA#:82NZ]28+KIL?[]=
^OE:D9a.XTX[B)dOFbfc6b?T2E2XV+W)d1LZ:Age5.fC.ZMLVHZbB-bSR+@eR9_I
P\@gDe[;Q0b(G3dGEFF=BK,Z6MW9,>;)DK6036D_^B)QaA^PF=DOS)DY&(IeT/fC
Oba6ZJZ[fPPUZfQad(EGCCd5e_\UOHWF?YKO3NO=KTMC@HC\aZ35Sb_P<8-ZN4]N
cg1#aN>Z.-F<,5a][OMZg51(;&&gSK2CCegWeXPM^,EXYQ>HE12)gR>UKS39J?+d
?NDfMc#cg?P2N3RY2@],TDPge(U1^.B&GL?59+S^=gDHFBJ7/Lf1GBTT_gQBL1;T
VM/^O0b7-P,\2YK[4gL5>OF,_(_TW6L\\H\>[:H#>1NGI\6U)0&P=Z:gF;=<AHZg
5IW8N1X-g=B_Fcd]57J632B<ED2N6+?OEd[7OP4Q0@^UQS,-TTY#KIU[\H/G/IS4
=<Ob3=,\_F_VY&.EOVH@]QOOF70?cVXFX6c#X0,U/VG[+A3.@:MD=5FB78:+1V?2
:aWB7]JZZeUgb3;M</RN9K)S.5(RN,W&QY<DU0fcAA-8;\JLdAef8B./,f1JDe=^
:T3_3+KcX3&X?dF&7)1dH9#U#3[D,(].O\)^\2XL^5J+0fK].\+\J\9J;3NWG-VP
Me.:LaH&9DEGJg<2]Y9Yf\4PF^3_\P3OJ(c86[EMV1(+G$
`endprotected


//vcs_lic_vip_protect
  `protected
.8\7>[-L:HE8B.5#:O=L,[eXPWdINfIZ-S4&>]\O,.5&8g2ddf7L+(0=-8WR+[JN
,_A95I)e6+Jd&f(U7,@N<F:D;<8/Ed^#2WF4M:3.M0aE:^6<Bd<VEaKGD[[QfQ>\
f<B1g1ab&)BWTN70V,L=8bP?ENX8Z5KW>O\6J=8>+d#)5G5;gSe0Z,;EEUcCMGeB
>[D^V4cJbSLJa?-+:c[Vf@V@KbT5Og/a1>J411Z/_97C/5TS+X2PNdR5.XaEF[Y3
de?#.D8\,8Y>=f],#23YV(b2S6#ZBPM,aHGc7&#gJ@O0F90I3,Ed,5X+34+e[FC6
P.XD(I-B5?5Xb/Eg:AfD,G\,4<F]Z-@Y7_PB>66&&PQ#>#VH1>C;MQgX2J>5ZfJ&
JE_2)=#H1T9CYL4_63Mc3S).F/\Y1eJgE^8=Y\cBKNcS,+5dE]U7H_fBGb6KJE_(
V-3K\F_O,LY09^5L8-2H/WI(NKf/2Y1&#&4SKS;IK>R:a)We#&0^Z<Vc4[PTPYMH
@I3\BSKJH,L_,Z_DW8DE;E,EI2[J[AbfIOC2_DJbScbOP7[[U,5g/.XNSa<444Ya
HX@0ZMG2TY=F2LIC6e_>?5891aDR;QZ5ZC#I32+gZ3=TWAbHO?NWJ,MJQ[IFX2U<
A;9C(Af(KZ4S6C@DODeV,aF:WGZUBP2,JQ8eM0X>6GS>-0,CPU^c?^-VVQaFHSS,
496NfNN>T&\_X<;)V7V>&J56UY=4)ba630A8U0[J(]L>B5R7_=AW60H>f7M04Bf<
g:L0e,Q(WB+:Xe1IP/;X3/ZQP&[=?2Z-5Z5A[.2SU<3Yd=8P[TX7X<R9b2]c#0FZ
_#_dHDaXJeMbK?)>\6DfYZ;#I#7Q:H;5;HI)bAXAO3.)eY7@;VQ0e;45#N(_fAH.
b_/Lc#-EcSL?EVGJ]f;JQeLTG;DC?725F);C/(W]F^WM(_IS1HX_.dAP/:-Za?7Y
2>U/Y3B_dQF+QXF(YFX.\2a]>?[5g5:3e0/PGg3WQ(.d[>VNX2G&Y,Y-Q^&KHY^/
J;G5Rdd=RMMS#4H4>)a&U,D=C:b;A]b_?N3VN^V?ZET@4.NUIB1Z@[_2N/(gdP1X
C^PF=2#S_S?,_GJAY9[.;VKDc7?GadEHdP?/425+:O:3Pf3D=0\UccbFHIE=R5B<
LSG6Ef:d@^:#db<:6G(TD>+1&dQK>M:<^@(FO;Q[.;.9M_?Z4b+?JOeN8#?T>1.c
1+]).?RGDI.ZEC3?FH?W8RDDgSUg709PSBJ\df1/b=db<:8Y:XRKXCD&6+-&8fG4
=a&6)Sd5gPIa8BSCDQ^M/I.\da1dRDc.f#ge)5cJ&CV/=\d3dP2=?UJ6?S&f_&Zg
I.F8G^]VAM066;BI>8N,e0M#P/;P[BSf&/Z@SFOZ2^.EH@fZR3U/BWQCNEE0DAEb
6@/\G3,42ZUQ(#HD^S^N2=82,AKERGEPR+Cc,#M3J@R>EMY)dgTc9,/Z,L^V3W7F
#VB>#+:]90,><;g9=.WcCgFFB#S4=?Q[L/W\/MQ7+^7OJ)E&HP[P.fS#T4b=8,NN
Xe[XLJUB70gPdW-]NW]A)H#K:1&VG#XOUCf#WV.JJ+KSO#U6PKNC]@Sc0Ba39::;
3-7\LYAeHFVK?+3#P^8X_9f+QN&QfSWeZA0(SF](2(\Se4gCAT>.M;E>V8?GM>YH
5?ML5B]2MGZ\d=>-E>VVgKaT9)=I5+EHA\]1[JG^_R4[7bX.7_LWV3<,89V908T;
8@3<EL\^(CFNd+.HUS=M6b&MS^b9bFe=3RbO#E3GT.43=;e@:>^28H,#D6=,T:C[
Xg2_A2E,O96e.[1d]HGK279=Y:[J7#&e)R2\aLAC>;(e+[1ZZ@MT?<YU+YV8#=\Y
2.,9DLQDZ\Y6-TF76.-XW:[bVSLfIKa#4&H/236H06X<JH0:[3:@da3/;5d&1G:S
DD9(&A3]B0A]\63UAO1US24e8HGF0MU4L]Ab.R[K0JHZ4>gEgg/)WVOdIgI[[,e(
cGJ1_>BTD2H82N(-;W9QW[0^EQME+TVfL.@WK4e31Gg7@<W4&N>+)O#7JIfa>)/2
Z.ID1SCZ:Z<13f1WZHTI&?54D8>E.-D/I4H@=@M=@/PN5N2HKT@bA;=_CKW#/<dY
<8I34\[bWUg^G&-gHfRf<</3=0[fUYX+(fg9fZ@M7af8CPO([fX<</^F[77:5+;)
2^LU^5,[bXV74,2D)Df,(Pf^G#FJUBF]X:.=XbVRX6HTA1J.ZGBI.B\&75&T?(G^
dGYGY&6(>H?G?^H8f1aKDCV]eNI9H:K-TQP=:@\g09NI/K0J\HU)P6V@Z45UZ1#D
Q](ITX/RLN4+<8MF4bOd]=)V,O8:C#_(b-V2_L1_/4>V.7cWHIa?YFH=)SfGJMX[
_a]J\6BdPbfKSAeU[.7L#FBR428=>Z1f-)>+RgK+4C[7N&K3NS8&0@cC5M&KBLL.
]Fd[OSEEUWQA#1VH<RgT;KO]=1_-93,(cACPH:)V&WTN1X4#b-@=0I_H=KDVCJWG
+dUH3WLT/+BTI&2H>2bBX9W]3KYcAK9H+PT)=c@:5[6YM.XgF9RTI\DY?C@c4,a@
PB&=G>b9S&Ba>d910&I9E)??RPG57S/,N)UNP\EC9[#7QG+5+6Y&Q;D@@J-/UD_1
Mf3VG8DT90B23>Qc=-/A>OO6-f/Le4=8/;9H0#RdcMLKD.LN6[acK3]Z9K/]K@YT
N,F?BT((-#1TeZSJIEV#)a?JKGKcN<V0d5RW(3>cI90ecWSN4D\SG,X[g_CbgZc(
7-fM#f:U3a(9W96H>D/=-cBCRR(@@ST#L4VX4OC,M7?/(#(4K@X8TSf\ZSW_+WQ<
c:#\J&L;K)F[E[KY(0E=B5E?,D=QgbXQI#TG))OEBA8Z^#Z++.E06GFBQ^P=9)K,
f]8c?:1\WFI3TBZ1+T7-VHXX=N<Qec?:2agQ;HAL:TRI/OJ1)A0)Oe(@3eU^#JIb
NUN8+5c_;#7QFg<S8T0<>N]9#3f?(QN@RM?>FdXVWM&T.+OD&3>)c9BC8.U5AV3K
Q7AR[WG])<@SK>NHTF)f0C+TM&=5:/=LOHL7#)XW=9d1;J9Q-6d])4;bM3<IWC-^
EUOUP8]=@<OC=#G6O0C<CcF[KV^X1SDYcG3[&F/,e6NG1fVf5;)Y(O+J3G<\bgU>
_OA9VX3dW7B0,Xaa/X/T=#[&U9\8APWaN3\MV=045LT,OHL/b]b:-Y[EcB=L&bOC
HcI;&:665aMg/@]D<7JNadK0<I(F0dXJM8@\P]7N0SF\c+FCgIa1>Tb/H9CV(K71
6#]@R+)?V6>-2e\<A\=]R3Qd/^KVB0=;ANW=Z5>>N&S.5/KLTE>bbEG:SOI1Y0Jf
c1a)7\L[a>;<D>_G.Q<^MJ5\dE&Q#K2FMO>deTTGEH<.DZX-Z=J87/+@ZFe1;f\>
Yef.DMCU<d;QAN0;<N&JDOJ<a7Q/9&75Z0gIKZ.<AV<&=2-(8?E1c=4_S-9^P:0P
&0V.Bd=,?V(GKS9)L?1D^A1g/P-#K\dc)VL]5#K-3]D]#PBTfXg2AbQ=:2^_g[6J
)eWH<NfE)+^)GZ5&K7Def;fB1cbI0>A3EI]^<>PbT7,>0TZg3A:2]OaJP(H)I@gB
8[#(K8Z&>Wb&LO4G>J>;:W,&XX)8_=B93Xe,UbeL5^:R,ge2IXCA37[fZB_RY:?3
@#]&SD8^a6_<aIS^4KQYQQGg,b09\:-daF#NVIfVFOb=d,3K_LJLXH)cT4fC/(M-
Da^LTKGS-FgQPE^J3-FN:7:F=HF(WeM+G78V?OCBaK7.D?)?A+9HE:,..0)KA;0]
HXL/K4T^THS\:OXC;-B0NCL]/VN3]6cQ-DYC;SHYE2OI0NO=L\gH\:YW4_\(O/?M
aCX28]J+-Y8,JI8)M\FJbaNC)Q=6&)e=RV@D&Q)\dW,#3-W:B6E_VLP:Aa7T6aY+
;ff.a)-AcN.(0Xg7#WeL,>Mc>E8_\GFNe@\B?X_S.d(4VRNF6bgJ<U&LeLa<P;/I
W5@9]7:OO:\.cFC\=+b\.&eeNS4^8=CU1bdHTZ(>e]e6)RTK>6Da:CIO:aV:;:HX
ZNUR&(W)(a+;CZ:RCW<OW/+([PaFfR_?X^Q=&O+db7:<=I=+<cB[UI9\\7L.QZOO
+C>(X?bH4f31]X9117U3K-W[NG+^7\,RNd6LU)JWW03?bOZKT,K.BJTYNUXV/fMB
K-\81?/V&G@&O)A0(Xg;,>d0/C>+.>7Lb?Q@5)CD=5FT:OFAecQ7]\=b@.-Q^RG\
+@V@2dZ0M]CUT.;3_dNU-/&[1F5b>aAF9e62-)S97f@>WQZAfU&A[fOBZT<W=#^@
:aOd773:cVL@a5N9/MUA,EabWR>7[e/\_+WA)Y2>=_C4gUV[N_=@J4cW^?5RX:2U
?=,dL?NfDAWK7V3Ee4dB)[PcVCVHXK&V,2DH6(L6HT^Y=&VHE>(0PZYU;<R,a:Y.
G][Y>QRY[B8PGU-5JNV8(<bXGb.f+Xd\@fRI-+O,MJW4f;R@2.Oc.=0D\HL6)ALQ
Z;2E69#[^:G[V?D)[:d78CI>G@1=X.ZAZ:@\RUb(c@1)S8O9Q9&;;c<O\QI9(b70
JSA_Q08_+@d:32bV5,2.-be.87R1C)2IWXF\]W.M0-0ARSYeTSJ.7[b1I5]4]e9I
#0#8dFb>=4?TaQ:aLRd&SZV5,@b:>V1.6&>_G[AZ<+_HG=P^L)K2Q(OE?ST=)dg(
]L6=HHG?O#5,Mf_M9_ROaeJ;+DBKEV7:0,==Bd[\^,=[gYQ1#PHEN,4L:\).)]XN
-b/=-)Q9DIS</W3Y1T.3#BCWKbSEc9TcU9aQK]EOMF?W84.:8WFIbf73fRBeR#\J
XW/R@RV1\52:bKV1fReOEAgFeaNC3,[=DX;Te)1V@bbD]b;<JdSFA7H^;P97L75&
L?<]8>Hf;g49?#bBeWSWEN2@H0d]YJHP8M:MDUZ.:&(P[,(=-H5H?dWHKaf&?2dW
_6_SK02)0ZS8b;cEQFKA_0;[1HGB02OCbU_U9/+]KYZNS0SN1,)Kcc+1@FZ9gE19
RV8D/V:+Z&5=_SfJ,U/<(\N.\:96)L>560WIV[2N\Q]=fR#bT4#CRLT2@H/aPe3(
;(Ed0=d4CTJ+4bHcDXL;Cb4E<[S\E8#dAGTe=aT6;c4^F>U-V^eNS\B,;IMMXMf)
B[TSUQfR8B@a-\HLe6;BR5Q@O.T#K.W#&SY.V4)Q8@G])P?TW@5\9.<HBZe1U)KH
@])RU@EM__7@(5Pa=#MZ#S=R)GQP;YRNf5Qc);F\LY#JS1_W[#7_-K>IHQ[1ZW-G
I1AE-7=?@>F7DI@5HA\L2,D/=X2gC7GFHT:79W/W\GSOF]g6]@@7KX_=1c?O4<]Z
XU#XbMMNQWSAJ5S;=#7d+SKXZ3bMSG&)C._E)#E=;:XLC]+H2+Q0J)S[6gd+\]O2
Gc+WfaOfC+W>UENLJ=af[^6O70aY4S+GQ3fVN;#Qa@]b-SZ=IPV3V1;U8gE:X<\=
b7>EIOKP,7BI6J^&J>8SVW?@4.PX@-dU(a^[)7+CW3c-ONZA)M(T9+JBV4_GGQI\
,CVZ(E).D(8TVf_E8/TS,4c@3KT[L5BgS<P>e,Ie0D=QIV:GKD\QP=e(O#.DY(5X
c/F:1.9B@e5G[MJZOSI]-ECZa#g,9PZe:0FG-S:06JeWG?f0.Z7\LFLL64@K1E>D
+\#W-_ND1-VF&?@NH754_Z@S<Z)1GM_V:E=#RIXIc2@2gE)H2.L?91[W>>XD7/;4
YW?K=O^fAU/=\AY;53?>SJD(d=3dH4QHP/02]],.L]f8bXS)cag5ZR/g:,DTdFZ@
>G+CE6Y>#c\1K7\0Z_J=RPaG]b]#JM6N&-54/(5(#78)5VbNaJ+[>JFJNcX]WE;J
]ff<X6T)-M-3O2?F\U(\>NfP^2[FX>:F]Y3ODP6_Nd1M9TXTX:<,QY6WcUVPROJ/
M9,ZE[]>K^Q-cH3[2b=cYT]8U_D1^g.\;<Y+bWa14ff;BL85ZV=ZTH84(bC/,:0d
D1d)1\af.LMEcE]ND:UcU,g2ZK&2#eQ7J1X4R,G]G6G8f^G5HBV<2f1S4>V&A\]b
&A@b_FUS4&a,L97gFH:Z/HAAPQX=6TH;;21Y>UZ/P7PIFG:cY8(Z/6cG/e#HZ&UD
4bb+[C+XNQgH/:;0V@/<9E4W)@Hd-SJUIFcTHXSJ/,J2>CC2KZ/<M&]7QDLT-R2a
-Z,8@N@L>D@>N7/4I/:Ee4dRLEVD4VJ3[3FgQ7)6gF6WKI)9:W5=Cb-b\@_,/3EO
;]A.6W:/^[.ETM725Y2Q=#3;V,L3H?PO)9ZF4.IgCKb[\C)+5aWbBWH?_<N.N/Fa
W9-g/PA<;,7;L2TL.28?]VcDOMLfJP^;(a]G7QOgEAb52^7TD-1(Oe]Z0HdI)C<c
cFE0g.aQ:e84?/PXK#^=99g?bXFYb,DPOb4EM^?F/\4\)[=9Dd=:L^gM2Fg8a@OL
e.6HC8OI:?cGeJQ]^^)3?J(M&EV1RVV+/MQ#gPH#ORfM1a(<&ddZ[=2-X\a_[(UP
+>E539R0a>T.9e8H2AXgBNQ=gC@WCV318N5WGR^(VO,4YBP6X3)V?Q2)-J40?=6Q
1c086)\,bCD+,3g9XB_Eb^+7<^_-.35cK,U.M.^2]J_3TT\=??;S?e/GSEUV9AAf
,c0)3a=CNW._XCO,6#Q_>M4GIE:>SKS2U?R\C&5^HN#+-524NM2BUF])c(ZS<LB0
6[JH0:B4L4QL9eO:D24=KQOM)(G/QMgPcb8]\Jg7ONcI9bS:aF@RfK+>FC_F\X,?
8[R;X>;G\5TfS9\N9a9[X,ddSaeHG9^QVWN#CgUE=4Z1S:-&eZ.77[a)#=e.;Ag>
R88=#K514(9c+@::P#CWEg\JOT0=a6>N=0M10&EgfI.=Ta+PaL5[[]&BN;=P&7L+
/=>E(c&J++ba.TB,TdWOG8J5?4-f>5.9NQAb,G4<,EI7dc)f+WF1,<Y?_<ISQgW3
2X>9^L8M4=2Idg2:/Ig#LL))21V^_A8O/9JaJQ]#>_#TX?](B@X^1W)XS6NbKC+=
DT@?A@Y-;bT3JIDPOAAL7.Zf_(GQZeS/E+<^8&\D0STYK.YFZU<a1C,L\:BU87CB
ab5<S8)#36&Fd+;/^E,b\<c\daZ&c?c7BX27(/?1^0#[IeC\?f,5>J=M)fC@?Dg@
+Oc@O#51FBQIQ+=<I9,E?@dWaV9D<M7-MJ[,36Z,H9Y8G]4N)_=cE_=)ZJKA.S4#
fUQg:@0+^OEPaOWd\_MF(5EVcA,YOf,.XJAW8+@+T?DNKbJAWM&#YDa=&]OKKcQ@
(c)AK>R]]\#.K<G:(K9>(ZSJQ/ED&RX&BC#,6DY=&H-e(YO;.AJ6#,a59BZT.b-P
CKKHB&ada-2&/bUFC?E701D\e@f+e([JXFLd?(6^[?POX-Y\8E&@>+3,:(ZRC@@:
=_)V3CcZ##Vd>bCX;3VUC^;TZ+YNX+dJNdPH.L=L,f&<=HTSOIeF0W3.4M/VZb3/
HdY1WCJe51aKe4Q?7S[Qbc2SWfXB94T;IYKdYZ,N#A2[T(Ocfa>)VYPOG_=f\<;8
BSc:A+DdN:/Q<]+7Ke]C=OY68QbKTW9[8VCe4f4?590D[]9Cf<5^K^_-)_cGLV;_
,Y33=TW#dO\N9JOFZ.d3/KNI1c^4(G[>_UYE2DX7,#T&U64LE3_g&:DO8(\H(eI4
()LUOA_:TI)2J&U=^KPQ\GN](^)KIfL4f6^_0(CE>)Db01R;0L#OIDbD-FJ6QNVR
P)@J+-1?[/Q]aHObY05X-C^g0Q:Id.WgZY3PD\&80aPZX9]G73H_))C1#P4eE9Y-
:TP/X#>O+H2])$
`endprotected


`endif

