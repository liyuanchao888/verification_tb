


// =============================================================================
`ifndef GUARD_SVT_CHI_SCENARIO_PATTERN_SEQUENCE_COLLECTION_SV
`define GUARD_SVT_CHI_SCENARIO_PATTERN_SEQUENCE_COLLECTION_SV

// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Request Order Write followed by Request Order Read
 */

class svt_chi_req_ordered_wr_followed_by_req_ordered_rd_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
V97+F<S@:=46^>3dSQ5(+TI,ASgAI;SMgRT,E127MWe@WeZ-B;F=&):SZeb_WeM?
(E/ba3CG+]TJcC3]LA5J15+0]D_V^T&04TVf]0Y+F:X:Hg-N>2K=_.&RV\b4,Q>[
T2=QEHT2LZb_gQGc8CNS\?Fb4&RS\W6QUd.F,eDB#=T&]L6C)<3#5<L->+g-)ad@
f9&D_#G4OQ?_SU80G:2=TfaL90^4N56^)g/]9_PP>7?/bWG//KbS,=aN+DT<EXE,
.\G0R3VM<#4UgOR_Cc284d4Ed;DdG58NMd<R>]DWbCg7)HC4aN(W.LV^WRMO/d:R
JOYM0Zb[5[O0H/=\ZTL<\O8.&1GGU],DV)INMVcVO(1P\gWNbU)g.RE\./+f:_gB
63W[QF^.aQc:/WD8P<OfgK_X1]Yg^^SUIcDS34A-&B5KbHa=3U]6IEg)#;7RKE,5
P6BgUW;?[\#,OLXb4Lb>9ad/cWf(KF^#&_b##Ia,Q2Y].@gd&.KV68fa&?M\/M=^
;N-J@bZN97PPfFP;<Da4#G+aGd9fAZ5#_SH86J_JD6S<JWSb#VeO]1bcN?F.V2Lb
46YI3FTHCe<>HZ16FZ216W^7C?/\[P4^\5eAZZI]]?UbGJX8N0+,FRa0Wb/@\&OJ
M27HE@B?He?_:UFeY7QVL_Md2N/F.,eL2PF+YU(DGIMgEeIPMe^8f[Q8dF[OX2ND
OP<6Wf[^;C06g>aGIgEV\&>Y0U@QV+XURDSE668]KSJJBP4OXg7C=9S_;HJG/cdP
7+UZP)R>EYd_GF)+06#P#aLMe_-1ENW(9$
`endprotected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Write followed by Read
 */

class svt_chi_write_followed_by_read_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
+GIN(^7I\X8TK&?^f8-PAI?AdV2<B72M;a/GMW,-5/]ZA&(,L:KM5)CB8fTGJM5^
-GB]L)GHg]5L83dPH-Cf?,<,Hf>#=[S)O7K5TC<CDFJ/F:2]QLQ_HI\,--Jg<C9N
DK2Y>7ZQ/IK9bR=RDM?#>[NID@33@b-,/bE3_@T0Ae,YXQ_O>-4FSONAIYK5</<4
a\6AA64CPNUVFP)aYBa,A+5JZ:Z3gcRON/Rb/eX=&B=W33fM.H>GEQEAD7((dKD?
\EYN#dBd[4E]ZZQU]^QKGB<5;Y:I<^4^06cGDEa\<gMcZ_7[1U79[WOGE1/f-]QG
?g_\<Y>UQbP4U+ME(+e^,#BB3NR;FVN]HE=3S6C.C:;C,O>_.P8PVR?J]5YGOP,>
e7:W=Q5/AO+>>?>\P(CIW<:2IO?d<X1PUUFVV/aeMS@McDdN5(G:;B2KFYKRQS0#
J<R1BO2.5.L.fBNU7ZIRGG4MBZbcQXBO;.]P&FT#5_=?^W6^\VEY^6?_^;9[)DWeT$
`endprotected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Write followed by Write
 */

class svt_chi_write_followed_by_write_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
fU6aa^\\6;]8O=X;^B_?:W;\<OV6MR^Q,-[=HKAIZ@&a@LE,]b#-6)\;<,72BCeC
&_6VE&[J:F8NIUSDZc2Oe+g&=5W2<07=HW@-g073X2e<X&7d:cOG;dUTYa7.-?CH
XBHA9QPZW)HW#-PFU]Ya/]2[<25O2W=PEBT2caaF9=:V[@a@=XP=Gf1CGC@F++QO
?-Q?33@1_YbE_(-:]\O9^XNGAZ^8Fa97DBg98ZW6Wb>8R&E3);8B9Nd/AY\LdXeK
\U9AE2:9(A14JBT\H/-X\a5O=WfH6cSL]8T+aR2O_R49gOJe2)FeY>/OZWTEWO-G
U]0Q:,&N.<FA-/gZJ&C@4[#O&gG?A,C^/S8GP32Z5>5f+fC8+/#bAFCMQ6FZ3NfX
6cN4TXQ63>bgTBcdYGaMB]L2X(T39.3^5TS?G;.L(cD>gQ7+O#^geG00JcbZ4E[+
R40>#7XPWeGGYV1dQd:U>-P(&AdaWZX1.UbM>a]YPb(f\HS=F?FCd1\cUY.;gO.I
($
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Read followed by Read
 */

class svt_chi_read_followed_by_read_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
7GE;\/0c-N)Z4B\2Nb5IC=L1&_-P\B\E9U#S#]:PM8:/L2.2Z8.+-)CG&;=S7[Q7
>(?N7TALKMG33?CC=6Rf;d=,2L0,0FXf6,fc[&g#LBe+a1e)WBIBc0gVBJ4I@[TW
XZ3SAbJWQGC&c@@aAeJB/eRLA+d(@U?BO8>KGa+-K2aB4\8?3(bA<716:IW<f8M#
:dfJIW^9)ZYHc8P&]7ZR(&0]C2<B_WISR=4\:g/Bab8+^1;N6HVeQCJZZZ+Z@e#e
]?0ZgLPMDGf#DIdgGEe;-:>?7N)N6)H\4CP/7gW=ON8RR1.?2+>BRA##F>+UbIR+
LPL.V(&5N6be@-F^9[AWFWEOJ#I]WLYL8T&2e1(.?/B(7-I:gbMa5>_>\D<.>^[9
:cfdM49<+_^9Q@M0WS#(bM7?&Vc9@A1ZE02W6G^GLe&M91G?c]84&+T5L+A_N\T2
]bb:_[1_-fWEQIL+7\VSg9a^T8HRNS^>?17F(c0_X6XYE:2PcBQ>:IT5P$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Read followed by Write
 */

class svt_chi_read_followed_by_write_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
\8XC#[FcMT3fTSB8<;SXKE,S(]BUJGK/@e\CTPO-f_UW(>SB[gZ</)XE/F&0E6F4
N)^&X2+Y[2XdU/3952Mb3Eg=TN\WV6@B\e^Q=XRa#FGgaXA]](4AR95;\GP3UeQ2
.Ha#[U.SJ[=X3+@AE83&GCS87(,[1Y><)Ua#T=FK2-.gK,[0J+F^H9+=B9.Ra@Ec
?(XcOSS4.6.-RUY4Kc[PgB@(G@10:@e\WEJf]8A\8cSa#UCKG-RMVgS7A4ZVRMSI
&3FHdG4W:DOgP9Sgb0@UJ<EIQ?,5Z@#@D(aNMHKdAXLRK5T)HL_X_9X8(003_6<B
-H]H;HJJc+U8C@3&(/d/MDefG?Dg>F00^:U[X9-XbeOC_#gd3K[7E:F3VdT/AEK<
@HCaa)G.]X2PP29AU-]A9@[Ib4]EUB<2O<<FT274+#^DD=)2Od1(S6SDbQdCHReT
I^d]S^#]4PQK:L+,e-9/dR)V[BC2cYSSTB5ZEY&@acbd4fDQ=Ed\aS+MSQA/6K0[T$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * 'N' times Back2Back Order Type Transaction
 */

class svt_chi_back2back_order_type_pattern_sequence extends svt_pattern_sequence;
  extern function new(int  pttrn_seq_id = -1, int unsigned  n_times, svt_chi_transaction::order_type_enum  order_type, bit  match=1'b1);
endclass

`protected
15\edgE9VDWdV-?K626-RU@2A2P885_gNQ=)9ZJHKeW^:]->MZON2)US+1^aV5K:
#]<SER5<(EX4?^BFRXggJKAF8IQg=0a6#<K9ABHdH,\>bM\XF64HXfFZD<^ZO(P^
aNa5_ONK,RH=<7K5f9PdR-D(+2F_+5L0ECRQ\Fc>7-O47XZg?N^[->5ZdKAF9OF6
YX.-_[KTdTSaV4H<bU6<NJ,=_E2,4T>K1Dc4#-]9-a3WW_CeW;CJ:b=].>C1b^9L
SbLP@8(J^6CW<5&@@I0:>dc@3)?@GU<07#E<)\(&e1B]aMVZ-ICcZBYD6[^VAWR@
SM=YI4Z(:)9\2T:IQa-Y_5\Z=aH\],8C+FYAaF4_e8(UQDV/;2\O8d0I#De40BBc
.bFe#c1.I2TYa:LQ5c).:R7R7T0TLKd/V7\&e1+cR62S[b7_0Y5NV8M(]Lf;H6QY
4eL;g5;7b:eC>;U8PSFO@J+-_<2P2\EE#BLGM0ZFL<PMD;I2\+2(.+,M^(gFc(-Z
Q5g=5Z0&,G59eaaJZ+MA@gO?F/0gB89=^?T6F/d:?)d?SJWf^X\.:RKWK?WV:4#,
bbJJXDYKHXRB0P2=5eO]^?Hd+E/9NSJ2K^PJ.4_H;JfC;\AGY4e-)?g\A2JVM+_)
b4U.gGF^gbI8_^3)2cJZ[](92)Z,KQG[;GC;5]6R(0g/,1VJ>3JP?GfJOA/X.&]1
_]8K@/F.>ZJ;/FZ^2.-EIQSEIdB98D6H9\[(O6]EgZ2\?Q)T5F+N:aR1L&KZ<VcQ
:A)O.b=Ff^5P=D/44(:7,F8-JUB,@LP7B(b_QU&_Fb7,=^X6E\GKL2VST118..,G
QI/44ROUfK5gbYL&G&2,:LHI1K_/X3UZeKLIZP<aVS1H(f]J)aGF&dTT)=+CIa1R
c@E;0BC4Q<YK^c_1VSAOQe\2J)W=AfEVI=KWdeK2:.ZFDOb.J2MbWgf:g^;4)6TZ
[_R+\&VK)&FK-$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Non No-Ordering Order Write/Read followed by Non No-Ordering Order Write/Read followed by No-Ordering Read
 * with Same Address/Different-Different Address.
 *
 * i.e. '1. Request/Endpoint Order WR/RD[Same Addr]  ------->  2. Request/Endpoint Order WR/RD[Same Addr]  ------->  3. No Ordering RD[Same Addr]'
 * i.e. '1. Request/Endpoint Order WR/RD[Diff Addr]  ------->  2. Request/Endpoint Order WR/RD[Diff Addr]  ------->  3. No Ordering RD[Diff Addr]'
 */

class svt_chi_no_ordering_rd_after_two_non_no_ordering_transaction_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
CJCKH&AM_P6-+O;N5.8(_#[ePEENYY+;JE41+>@SQPGJ30.+e8BD7)I&\eN:.fF,
Z>Y#55R3C=ZIA4LI^]+fODCD@[R\#Y&3)#/\V@2a4f@S3=:GT8J2Ja6FQ3Cc;.L+
Y<MN_4ae/6II>PIXAWFG10.+FOa(@R,aRKcN@]7,+_>0:M^Bg>>)b5b6#JS>d_(K
=)<M-S7Z.QbFeY+Xf70Eb8X\16:Z</WV>#E-1.1F4C7[fXH1eDN<:;W+=eV(H1:#
9(4VG03];+N8B(g)XK?TO@OA2:=Zeg8I)M/3H)YE:L4FR@=<BeC/6YJ7?D):C,:W
3L[XU;PNA2H]UJ+17LI+]I;/g/[0,U.=KIO])<2HOOLG8OSHT4\T<)O_)O7)H(Xd
&5c_/Sc9KbTU?:I6eY[&BK84)?8(;@ZS<g^1=62_W5XJPC_/4SgGILVBQ?/:5RY+
bA-S>Gb6./b,RG/)X71C0QBT_>/F/aVX]cXAg#45[Q<9Yc]BXd]9fM0(#DX<@X7Z
P8C;Z:#gF[c0]#P^fVQ>)CRBd7M(C<[FS2/MR[(bfV+Ma8:ZbK<-#UfM7O4I-+__
1;CZU4,U6S^9]9;&dRFg?(13D0AZEV]IJ/7/3/::2L&A5/+Q0B.cKY(AEVFT8H;]
FG5=d[#V\U:@^KU;cS.L/I+NAf6D_/.ce92=3T8b9-eE[99IB;]dM2.8+L9>f]@e
(]W3B_Q<TFP?KDLd[_BLZ/e;P-fTIS_.2Md3cg09(\73H,d+I15V4@S.++:>gYIMW$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * 'N' times Back2Back CHI Transactions of Same Source-ID
 */

class svt_chi_back2back_transaction_same_src_id_pattern_sequence extends svt_pattern_sequence;
  extern function new(svt_chi_node_configuration  cfg, int  pttrn_seq_id = -1, int unsigned  n_times);
endclass

`protected
0d_,Zf.-4]IWKcG.-N.]HdP3g3b-8b;NJd93]66QG:<A=T=M&HUI-)=]V2bcCg^K
F(F0]_2cG?Dc^gSbM+0FGPCDF8BPAMST7f_J.AQeZU)H3X?PWW9-(P.AR/_@.YSf
AVee+6XCVIgdYS^Oea?BdFZN824(1+7eD954<ffOVGM:7Y]3X/YMA+EKR]]aR5cX
WP/WGQeXJ[?XM:_[NRZCF?6W81,IPM1B-WcZB9B[0W^4G0eUY4PD,40=B3SaLX>^
=Y)-Tf,M&-Q2Ca7NCU9+CH&60]fQ.<fL#8P1[I]MPP@^ANYO\UZ<O_82W?32bU42
\46G#Ag>W?bcfgdME9BB\TYO;4YTP?[UGU)=[?]W0f3Z3[8?\G@#BDG=<aY<U_O_
;+CL+Y&H;]>=7\SQ3Og<\9fYHK2+O)-94LY2P]C0,E/X4VeOD9I;S_HV[K]LQd6+
L)3WgE+RFZV(&BB0N:6f?2N:^;]D-)KMU2-\>T=/M/;P99W<G8\5E:+.1+B9#BZd
F[J2-[9RA9]2NCTaRAK1\L-P4J4V0V@V_WW\P55HY0,[/1PF_[9&[eOV6WH^C2.P
CYM)EJZ&<EW=[#UNV=7+(G]5FHSG6&Y+ET(XMC,@S(.CMS6P<#>IAFQU>e=@\:(S
DW]5eZ7EU:eAb=EZIXUQ\_b+:^U0I_Dd.9dBf7C>b6BR,F]PbD;6UL=0O(.@X/XX
0P&&?0F[G6Ib//J31MWeB-K/F=BF)g+_:RgKOM9(+VZV_J]@&)(DYK2TCZ@)56LA
&g73K+N2?#G8P7@e92-fgP3V(BDX075DDS<,WQ##:8FE5JfE@87)\L^>N.:JFZ^+
aN]/\VL.90^C-^SCOAHC-B]ZNZK^0fTM1@7\gN;cd:P(dVZU?PQ3T/cKXQUT3FeA
ae:,A1#MVLYIVU#f#AJ96&>QV?S+NXdA^+YGPXVb^=&?GH1=I4.Z,bD8EYRb?@-^
YB4[[Z.0[\6B-H)L;.2E)PG@:Hb[dNad)(MX1:)7MdX0ZX<8Ied\d?)&L:(46;A=
HcRKcDISYB_U.RVD[QRBca^4SYTFUW#c;-YaA3cFBLP\AE@f5T?SL-WR<4:YDF41
Od+7;g7[MKN+:?8a_Gf1O<VC4cB[I)O+P:.\Q(K&?F(62f)fFGBbZFTGf1MT?_2\
Nb+#01CO;gVE9(ZO]@S;1[(?C]PF7SNE+S;@E7#Ec8W6D$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * CHI-B Spec Figure 2-23::Three Read Request Order Example
 * Ordered READ#1 ---> Ordered READ#2 ---> Retry Ordered READ#2 ---> Ordered READ#3
 */

class svt_chi_three_read_request_ordering_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
[0U+a<<^NKE(Ae-6?N>>f01fU@G@ZWKT#LUOKGTDQ+8eI22<X^336)W;/F>QZ[F[
BR2WGY\1=?CB\0]c5d#&)b&-efG4SKHd<Nf)YGHPO>XXTe:NN<ef^eIURT6H6_?H
GB];]d(0UbJG>DY\KHPUGFDC15\3R3.bH@B_bRS:(X6X;S_1XRR?YIC21gLO[HY^
Q_I\R+QbJLLdY.V1WG0E3\9C(WCR<//c[JX=Y)Bd+Z^\#E2=cfH&N;,/,gfJ0X<-
f2F62ePNO)DN^XBB(G.O2=QJX4T2(S]LWV?^;V=B.b][_O(Be.<7_&#9_W<S;8.8
\]E&0e3]VDX1aO1??AO]eN-\U]M]BaSB=H2=AYMKN^W@[5g,5ZR^4_TX8IHXM&f^
EF/HK+/:e8Ff/J7f/A9E)&>_GXeR7Y/\f1?gYQ2NZ_XP64=g=529V+#d?/F/UAEe
dFaUEc>40>dDeH7;N(40DY(9^Qb\=e,((4KgCU1KJ?TV-g#-QaF0N;>dPYUT,(J7
IEe[7f0=&@BB0XA@\-6L/WK#AZ:KA0HOdJ(WA@F3[6.[&aVGfT)UMY)d^/Qd^4#-
cHFF/JgA)ZUZ-g/#b556?FF;763DF#9.GbG,dU5B?2/Af4e+7aMP31gIV[g2+4Yc
<KT.2R7e:N^gcKSJT4P05O?W&e)FcC8S7\a3#>8;4DT^#?E(0EJ1c15e&)_2XT+G
69V/Qb:G>e(5O68P(d.9(G8dd.V-ZP]>R;G858TBT;ObML5bfICe/F-<#6)=V2?A
KZRUdQF-D\C4dD+@:g9JRc(GT51]&BAK@[b6fQQC=C^LX#4TH@>DH5MSTD-RI9UQ
&4:ER_ENGd=V>WEJ=XdHbC:8dWZSed9Cf^\Scf?A6T>G9Y.bB71?GeP)1/D.gOBQ
H;U0+8cMK;;29baTSV(OZZS_>>/1LILFS8#\_bZa6Q_3@ESNf39=^0N2f:@[\9\P
dc1.[L,-2/U&2,R8?=M-[_DHU_(Za&)Y74HW?H[WTdc)>eaf\7,MK\:=W9gG9g^N
[7U_/TS)9\=ADVK1UTTIC_3-PW?_PO;4Q2cY;I]G=RWM30T;OV1AYd/7O<[D_,=)
cB.ee_:MfHF#Qc)_BAP5^&P6LOEc)8JMfD7G.1:-Z4D6-=D=TA&,JG;8WC3Ceb7a
d5R7Z)VU#O,4eA-?Fg1&VKX/11-W6fBQM2d.AD[fE@PVOg&I(1J18/cF_#,=43JT
D\ZaGMa^6=?]:#U[H#O]Xd>#N@M/g^WN9X=\L9=PCVPWP,edM]3aS4F]C4=eN]VM
2^-J+JN\9W>0&O@#]KEfMKHIOG0:.V9TO:\4=JYJG,Bf,WL;D#P-X,1K42:89^D\
2R\;C5WES&dRN9:M<D79c^&dI^-bGCW7MgG/CCd;-X,,dgJK>65<D[gA_Z,7+/6J
@FL0,8GB;N)R,$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Retried Transaction of #1 with same/different TxnID of #1 ---> Any Normal CHI Transaction#2 with same TxnID of #1
 */

class svt_chi_retry_transaction_between_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
c,+3Sf5?-gQI#CP5)#S(I=3)\TC\ZcSK/71#b#d>5SYQO=N8,B+I0)-HaEd2WE8<
T?S:C:g1B6VXa-Hf,Z;37PHBDD59ZF.X2<(#JIL;OBLe<ZJL3_VM#;gDWdbTFNQ0
8FZHgDFUY4aa2>[[F#3c<g?@g0[&[@Ua\XOS-W<NW7CE.=c&db,f2^fPGW,-WEO&
T+PV1bT<0@CgZWK)[EV>3V;Q?c+(feDe((?5LRN+NRA3#Y[W<H.gbagc:Q/PEZ5g
]]K>AK(TCFE2c/(T#C4gQ?OEXcbF-\/<+-G8(__#@Z=b:A4Q1^A0A/;6]:FWNN,Q
UWb?4K]-?JO(<B3>#Igdd.9gbgCKcg,;5Z(2dVa;&WL=IBc&]Ia38I40QSUU[b9V
V,0HTg0aJbX0bgERUC#XIc]Ae&:ScGOS;0]cRY.Q>eE-(6CMObK13OLUCeBgYc+T
KHXFBR[c/4[6G=PMD1XMHH-e/I7<KBAZ57\0:Q)QY>0((T+RdI,eR^K)gNL2KYYZ
Q@CDJLWY/bO7I5#:TBHD3K#8I6H_M)a-6/GAPdZT/e9=OW75Ea;I#.Y48HY_dHZ)
)d6Z2(>(POG+Lff.R84[7@_I(7a()_-/?HL4d5MQ+Wf=E$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Cancelled Transaction of #1 on Retry Request ---> Any Normal CHI Transaction#2 with same TxnID of #1
 */

class svt_chi_cancel_transaction_between_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
>^.?E;=A@@9KQTgF_&Q3K5M)Ad=S_[NWT;&S]EHc.Z33.)7A04bB))W[-cXD6.e)
_)@(H3?#7/\]d\+3)71_RX=fDH;C<-SJ3f)]]I^3-:aP3.(.==?gAXM)dNa;>I+Q
DTb_2H=(:F7\A>KcgV1Q\TQI+X;M[,Z4+\5_=-RFS^C:VH.0JA:@3E4D^#\3If-d
39Y3T[aW\[/eT_G;L4KBDg9f5PMSY.1_(OII,J+I4?WT,).)XKD+bR.ZMNW+@XS1
W4e8N(07@\5JfX:EJ1f_L@=4\2\4<b\NDGXO@[P#6MaZ@b9;FM\gefL[967PJ(.@
+a4d(:];?II+#V1Y4K+>2,WcAWC/-N6,@6UX>#P9=7Z&,(#70N<=+>Q_K6&E_U__
(GZYN7:bLCd?Nd)fD1ESPZNZ/KDH&W9S-2+=1+QGOFeN?,[bcN-[SA).gO3PU(#e
7:II5b,g_.]7aY-g^(2L2SY\_X55)c+KdE8cJ&FO3T]S^WVN)L>Gf?4He4J1:[^+
DO9b\>4LD&A4C9@IH;^=D[-\ge;4&?=>eN)>WQG6LP5e9U5+/+GZ_0;KUB&M?D,e
8OOZ<C#HReTYT01(^&b@G(-fFa#IM\b<bY;L2;:=VdXb&B8N@fCU?4M]W^6IbYU&
@2UIC,QcK@V;dNbO,=Q8gB-f6$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Retried Transaction of #1 with same/different TxnID of #1 ---> Any Normal CHI Transaction#2 with same TxnID of #1
 */

class svt_chi_retry_transaction_after_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
KF2IW.11d;Xed1DD[+6@<cVN:QPOKF-=K9g-_T,&cUa;R,N:<;1a2)J+><N9MSHg
aSB7NO.8_:J@/U6EePf2f,?:]@TKRX[AUaN)8_EEf@//887;.1(6gE+_U,7U#+K-
F&SODS^;V2e5/A)Y=QRN+cI7-P]/Ub.:YL^E&Zb<f/0;+59PW-5@#2/L2BZ<B(f4
Z.>bT;A<EXGS8ZS4<>^0</)c&VP]^e,@X]a0g/:.Wg85&49Z;L3G/F^WW\Nc5g6>
[=]7@<E-d>E@P+&3f]AULa&6&d+6XdF_;&>3GNHMLMGb9Fg[JI\XUX,;ZL[M.FFW
W@<JH8Mc&O5S1Fa5ZOe7ZIeP-,-fAH,(4IW,9S>bBRHEJ@].YVJSf3N2)#G.LI6g
I:SHf?XH-@3Q0,)+L>74Vd2cZ4:.XP1A9>\VRQaOD9V\><F(dP64@g[YP@M#080-
,f2B93<T7D(@G^/D54G/4A;e;4M>bUfQ>aYHe+B7EMYB#XT]B-#ZfIeRG\P8T)3#
dR>L,/\dTXC/8DES6dLI_3dL9DFRD7F154C#4M9<?]\Y+_K#>&_7=P)Xb-ZHD;b-
1+c8:\;[+UL>F=-f5C569WPY[U[>81SK@$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Any Normal CHI Transaction#2 with same TxnID of #1 ---> Cancelled Transaction of #1 on Retry Request
 */

class svt_chi_cancel_transaction_after_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
bdJ>#[\P/QQQT9KVf:8_U5:XM\619C.S]EB8#U,X8U[Ae@_?Ydb>&)R#\<d1+32B
4GSH=Z/e?LC02FTGGBJ0P]9:Ed45+:WS1f.6WW5S/0)+O,<+FP\::/5\BS1DH_6J
,M5^9e5&=L&be(fN@Eeb21bJ.ET>,=>=cM]-a>>U];?7<:3V4R,^,7>JQYe2=3A+
(#7IG&6AP8/.e7g6U\Be._(^65\3K:_Y=Na+E#3WO(+Q?VbF]He(Y:La^UC8TfO,
fE[;b((EQH;NEe^D5fWV-<C&;Q.:G0717G]50\]0;P[C9A5&3]J&fc,>GYY<)c:Y
0F-3<gg;>GX8NV4Y-;^N116IU7VgV9_2_6&Me=bI[)F9SVUQ)E+&^ARUe09+fB?U
Fe]F@bC-XVg1VEDD7:QRc?1AO=^Y3Z1&<AZ6bF-#bI5e30&U6WSO?=\,O&bLc[Q>
V[@g^.QDK./7)?9;+R;S.Q\V9Z/G[/#N;,G2_QB.I9[(RdD#D30A5VaK9gf4f_(Q
=>Ag+=BMXPS#TXZ5\JI0_.96.IPZMgd_C=5OW,]15WGU@aC2C=4dQ;/UON4/8BY<
;JRK9L@4b&3e3E\_90E4UK8@Q^Z+R?NXL>X@[(6M;ZZ=NAda5Nf)OFY+eWfL&OOG
FDZ@J))A>]?e0$
`endprotected



/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
9.-gF]Pa^RM/<eJ4OT6H6LHT)&G,G?-U)7BQK>LYFY-IQ7cQ/ZYC0)3BAB_P7bC/
PA:LTTVfa#6?0e&,(Q^[Yb0.9c.H8CeeSD17:+CI#e>\BVeeW&PN&K_1\Cb\&@HR
X\NV]NU#_?--.JH2YY83W7P6NK^G6;_1d4@C=XZE_V16-HVC#Wa__K6)aGRD@Z5D
8,40#2P4X+3VG1\Mg<fP9KaXZYg:IZ+W;0AQ^OLC?f;D^,7&&NGg<ZJefbISH_/b
_MYM4&36_GYT1@<Z89-([RJe_R:V&O+?LcKUb@=,>OT0PWN<^:e?Ic61+dLgLT^a
#_bDM,>Mg-ag,^9[O+eH)2cC@7XTg.O9[37<G9a1.#7be(=c8e(?WS8Y2g&6;8)/
U=,Dc&@?VB^1/--[6,6-Z6J9>W;EZ0R,/X45/,_U4=M5>7),NUPg)_CW-_(-SfXf
Q\M00aC#;5O1_]@BN1LOE>TM]B5<Q1@RBA;\JLWH;e+4>X8?HR=AIF-BWAPH8d:.
3NK5RAR]/R6.831_RZK?c21:V0Q?71C2Ld,I)?0We(]DUJ(8@6_XIF@_c?XONcH<
>2GdVe@D^.G;cC6Qa#eGNXA/>dddP85@,R1Q7?RMMbFE:HBgXB])7&ffde\+:Hc6
=5McBPgbH]<HF+Wd\P:3(c3;(=<ZSBE8LP\=H:2[+Y<Mc>EWCHB(;#ZN/GU<aJfW
VDWJVfWg\V2@O+6Wd^BdK[4F-\G7Y2J/8AJ\;L>UWM4]V1W[K>D=H8U,#cEdU5J1
($
`endprotected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI outstanding followed by DVMOp Sync followed by Retry DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_outstanding_followed_by_dvmop_sync_followed_by_retry_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
DSXgCJdS/VC+gf?ODX/.OFIM;KO[/C]fV\6]PC/8GKVF[U5IfQNI&)P\3F?cQJ\D
B]7W5Hc@cH35_4)Z?-84[W0ZYJ[,@;+^=2TbQEBW&a22#J#YIY&4Y[Y?<JIaF7Ve
Edd4]:UDWG.EE^;/VKU0^:=(G.V?fJ0M9+X,NBF]E7eCSf)A^^N1&cBP2bPLTJR=
G08P0T6Kd22C,cd7TbR4;-]?e=;SG3QD;Y/XZT<QFYX1/;9,23Tf1)^\ZbN,g90Z
0cJ<)PEMA,BM;&+2KIP0D>SK--FIQ-/RN^#E<6:8Q\(M,8+A7F2/d(YX,G0&7a(\
3P;F](\IL<@);FaMe(;?M]8QOa,.=;7.3Adg:UJY^eT0];VG22b15?,]WB26e<VQ
gPf0df=d&(\V61-(M=[)\@#+(Z&[CFOWb4g]c/\McL#+K&T5];8F5d<fg[,7gBR[
BfT;UXf/M_]dFSPR#36YNf_9Lf7J(CIRHcN.WB<7N8\f?5gfMWA+4;6@M#4H9@4U
S)I:AGS#6JLX](Z\2E5]Jbf1C)\Z6;OU:&fg2<+0#SNe?&KfOM)S_daT6^18<Q^\
6<X4/8N3_bSP](0&8?C6?fQ2S<&S?TRaELdM@\+6VHM0<c9cAYTc;D\=O<UXX^Eg
9>5#O6gPJ><GE:b+^-5#Z<9^8<a9E>5eK[77\UMEgM7bLH70Md1YSQN4EWAWPcB:
-7X^MOaX7e0&a:50,NBfAZd-=@5;Z_^S0TAAS(E\+W=G(_02ed/Y/8&e.MTA.BGa
ZSb+gZgUO/3J(7cL7>RQ&.aRYg]Y(6C>cB[AeH-FE.X#aDEXY0Wd7=Zce2GA;af-
XNA#C(/]3?#NMRgGbW05BK(I9EQS/UCL=X5HAWV#[&e0RFNXID3.B:0OOBKa?UeU
BgJ[f)@6Z:1JX1a6;^Q5+bB9;<[/@/deCCV4\1-L\4O[c][[CW4F;^T<b^88XI?bU$
`endprotected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI outstanding followed by DVMOp TLBI followed by Retry DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_outstanding_followed_by_dvmop_tlbi_followed_by_retry_dvmop_tlbi_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
WW219(8YE=>.IV&46fK_SQT2;.H[,L>C<@\Yc:>M.W&0K#8+SOLB.)(;-#e_#WMK
._JH&e[KY9O+35Y@>+4+A]4G@aGV#0@cX/M-OR164\)4S11K6eHUM,92F<QYC^Td
C-D4W31-Q#7BQ_^YCJ050.Z(4YX5&bNR4=+T(N2554g8cQRT[0aRB)?EBa,R@;5)
Ta=S-@cV3KJ<GI^,7PIgX\_[W9H1NOaMcdfOSc(\C:8[PE^Z&P;[,7<ZU5UV/W#Z
7S&ZCI:[)?_\/WNZged-=&?K=_M&B@TX?Z<+5&38<AO?5.c)\1J/a43)A4P)\KTH
eFE30RG;X(B>)2]Q.PWWFR\;bBg8;KKZ;JHYMBF0UIZa6/N_0:S8S\2L\fFI2Qf/
b.V<;9J::-6&aIE]dR<E)TI#=7BQP5C7+57NDXYZNW8e(9T\4I[BFPTgG,T2U6fL
T39^3L5gS4VeSF-e@V>T@]_@Z0S-<3gI>2YG47+ZN&4QP-C2914PZ=10WG8P]PB<
D>=](N4e:2)_QA1dQLI]][.g4>La>a6Pf<U<\7<@2SY^bK846DEZcS)=X_Te#X0b
22B8_,R+bdDWeYQ;2O:14KC?G1-f==)gVFC/_CLQ,<SV-M^N12^\<8(.e,U]F_TY
CMGD^LNgcL:GOTeEL.Tfa9?CLD4g(J=RUTa]DBZZ6._7MLL&GJZ?Y.U(J\=b;V@N
HMP,?bUZ(L1\.<QNfZ3:A[a.dUSg(HPC3L5(b;[ea#-;Pg],Y=IDH)D;]d@;gM?2
USP59T6N;O5WcBg.dI<-a?JYaQ&Z)8DPKBCB1X7cee&NBAN2S\)6=24[@VE8_XZ/
ZB3dQ?PV(66=KeVC.2PHJG>H[G<+g8C\TdNO/U?K2>&A;^>KJA=H-2_HYH.MIWG,
U?<6O4bSe9IYCQYDK9/3+d;ZE7Z6O>:1Hd;-G:SN#QB87-5bW1ZcXJ#S,-4NR)YC
NM?Fa)gAJNK)5].6ZS@8WHc=6&JPBCF<0KH6\FBYD[<2O0a]\-@WUcHJLL7L2Z].
YG6Yb-/T;7Y67bE]PMUF0^IZB1c>S-JH&0Pb)?Rc[OZ7(KbW]D)4JE][R#8S>7.5
RTKHHL^LbXa/^LZ4:Q5W@JIZ5$
`endprotected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by DVMOp TLBI followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_dvmop_tlbi_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
>JbHgL&gTF)4:##IDFNg9A??I-fQ&?RPNQJM-I:3g++AE4K\([W=7)_JG1<0I/VF
\JDSN]MB1>gf]6<B;Hf[UVg&S5fM&WW#GEFc.AV^H=66M#.0/L>9+\D6A-?S_Y[&
6;ZBR;=W@B2I3[^6OcQf00C1SXJ4-R_5UAe#+?;a/^YGJ5,F7beP/)ab/B:7T,aK
gdL/1MB+\g&RT>Wb/TZ0W7fWM^/UaL(.[UFe?BP5V9aaDK@:YGHSa2LW.H+9Ta5.
G)>@=JR::1;I67bY^;BRecbgb5#I2(MAPC.K.30M:L-6,JZ?:g7C7J]8?7^/R,8X
ET.24)[GPA[eH#5,Ug#0Vb1X-U-47=M9C_67S#G@.3\c?JF:=?,IM/ebM8;3#e.X
O]K3,_O:.VQM-4B#g:X_[b#S,IXOSEA<]A+Y,^#ZI-2_-B>FWc+[V^,Hc7fR9GHG
(B#</^UR1039Ce/0?3\Q-.AX8H<B1,P\dcFSZMLZfRWE9.H0.>400;_;[bTK49E-
eN=)A0eC-Oa_0=/?ENT770,cD[XGUZW-N[10a+\(L692BSDD&BYIb.8_</bdLJ2)
c/ZQO31S:S.[cVJ]A+32Od^7@eGN8@cKU:d;2T-bCUE<..^]MI&ZfX(.8XYLOU[M
?L#X3773HV&WEa3:)@]27=b+9;Fc^^eB?3&+]K?@SY,6E.VS26/QKFC(:7b_@,RE
>Y&,fA3DJ_NRPY+L7P;,(3<5S.ISNS5b+<H12d<2f0P,Y2T<bZ,F2TE5&3dX/4&]
^g-GCHJ,BW;0eg#HQ6@7A^?2N^/X),2&I_U,;CSPd@QHA2WJHZ2/BVF]]EP8=af@
[,b2eQUDC5c<98Hf&S6g@HS5XSC^9Cc1d;\RD[O[_2UT&C:/DcX7X\2JOXQ#NKQ5
SE)EI4Jb<0.?Od@FAaO4D6H(8bMEF]PMV_1dJC=FcgWR>D+AW:^RHV&[=BR5Q;)T
CU9+LK_(XL3e7E>/9fQ1+)QO;Y6aN8<)AGS-&[_;JIPV:-Me&,=0-b=GaVfMgRI>
+\A-1gY5A;7\D7=J-727aSWga[7Db<+2a.8Sa1<e5#RC[J,XFf#a]&=GO$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     CHI DVMOp TLB Invalidate Transaction#1 ---> Retried DVMOp TLB Invalidate Transaction#1 ---> CHI DVMOp Synchronization Transaction#2 ---> Retried DVMOp Synchronization Transaction#2
 */

class svt_chi_dvmop_tlbi_transaction_followed_by_retry_dvmop_tlbi_transaction_followed_by_dvmop_sync_transaction_followed_by_retry_dvmop_sync_transaction_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
#Ka1QJ#PF]_P1;:aFE<,4:Ad^=]bBgEZ\HM/,QT\4.(RTZ=/V?FA2)7Z60S/M3eH
U_CYOb=;aL#R_6Z#&#8BN?>.\(E<-Le6Baf02cXFgH/XR&+B(CQSDL[Kg\?GU6=R
I/6QZaL=9_8>\CR86]_-<]KYJSWH^<egSGI:<N;,-g4+^91&7gQ&U>\O68HE)=]A
b,DZC1K-^F<3NDMTbGQ[U=SB^KF5\@5?DDQ+F?IPOR#<OM:c1[40Q]R;2\gGc[3b
=AWH:OGX,Ne]EBA3Z>eSP^RRPdTP&ECA:ZbgVD6Q(UU^+P38,+==\.dJ7bS8Ub-\
>5V5:7H566Wde1]g5cZ,YTK6J)Q5XgO_=^&;\E3F:M)C@=C_OTaEBACbK9=bg.(V
-B2HNQJC9#.BPN7;;.BY^HKc:#4^,&]5JG1\(OYaS9;gBDBI+;->MIQP7SG5U,S1
a34>+8g/WQ-8-SW4db]@M7,/A7,Z&G[+bY@ULXdF,cG55^>L)L&&5\0X8\1O6V4c
4dZN/8cVUR\0PdQaY(8D8G5@W4R&CTDI>8W(##.GGP+>fTc1U5F/4&ZC[;F@B79M
#F/M,7_/B\[<8CA8a=,E?NBL)]B0#0D2K2=JdT+5_.^F5X?2HEEEVf[a,?Hg6^fU
S\NW+C)H[.X[N-;f(DPC)-MegM6)XNN?MPaMJNQ0V7>)AJ4F6G2aLCO69MCP<D)&
&Ae-7F?&F8fCN4WF+.N:(W&8(EP4F5Rf3/)Y#[53#9OPU].gJSGce6K6P41(F1#;
37,ZR2,E(0Eb8M@bE8AXOaB^;1FQJV43_?/_A4cf&5<U\1d,G&ZVVA&BJP#/N-AO
c[&9f#3G&?S_Y7MLL<aJ57V8,PANEN:2(CP6?NaX<<OJ0gHXR)S_;=_4CD8U=E=A
F\e=ZG7EEQR02O_=:2?M4A_7B=;.RY@D;OgKVR&+[]?B0R6(C,/CYD4VX9d:TbS8
c&;1&41?KN74f1bXXYLN>T/3RVR4,B8Ba&R2=BTKST/)N3SMKU^+8,BE@\ZD@NZ.
A8U>OQd2O/2b418]98P):bgO#+^CW^;75WG;;TWfI?T#)0_I@JC/WBgc;=AFQ@^2
SMSI13)YO.>G7CD).P#Dg[=#ZM=F0e4_^A.gPJe4[KD#Rc1MTd/J@S]@>H4-,XP7
VG)Q@8/MHL<aeRKT]03);G:(XA7Leb\/]gA<U:UaV,[<+@\\PLRa^XXY(6>FGHET
^fW[(CH:KJN:38V@LKdAJ8Ee71]4N5?,IRID.Zb1EVGLJ7dJZ.#LFD[CXd=YNOS,
Tc7d4Q:V]1:Tc+3TRVQQTeg2cf67F2:V#KSG&J:BMVDK>6J32Ce#f,AHKPG1;/BK
e;C(0#,2KLJ#9.dL,c0(XY]10,0U@[A0I)9RYLC5UA)e+3;&=g\I8CfA4^,;SO\=
G4b=I;H^Ig3,_++1RN0;7;O1T4K@\ee:)g3e<g)8bGE(a564.DP2]#Ld8O#?#\88
K[a5Jg<X<U)fPI3b=&=(VXRe9,G>PRP&O>KVVHM9X<]&P1Gb8c0FL3:H_?4MT?:N
^DdU965Q#8H62Q84cADC6;D3ObYTb)S9M;.c6#aL[;^abM56WZB8Y2Z==Tc=O@C-
N;&WH]XKeaS5O+^>6.LBfC<Z5[8KW3V=T747(N2A<-M6QXML;Y]FG+@B5#IVRLX0
a,W)G@e)NbS/.8W7faGJP\Z2/6)H<DLSbUd1-71)TJM=6,?>LY;<GT@BN$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     CHI DVMOp TLB Invalidate Transaction#1 ---> Cancelled DVMOp TLB Invalidate Transaction#1 on Retry Request ---> CHI DVMOp TLB Invalidate Transaction#2 with same TxnID of #1 --->
 *     CHI DVMOp Synchronization Transaction#3 ---> Cancelled DVMOp Synchronization Transaction#3 on Retry Request ---> CHI DVMOp Synchronization Transaction#4 with same TxnID of #3
 */

class svt_chi_dvmop_tlbi_followed_by_cancel_dvmop_tlbi_followed_by_dvmop_tlbi_of_same_txnid_followed_by_dvmop_sync_followed_by_cancel_dvmop_sync_followed_by_dvmop_sync_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
U)LTeCM(CB1>5aA&DTG489)DFgO@.H^O>:e;ZA07K#Af4Jf+ON-&&)beH=MD6I]D
g\:e@3I0-&_X@<7#4D)-O7Ib)_NMUNb<@JaWK^g;D(A4^Q+F5[HB4XVR?[VS6]^H
O9c3)>4Ye0-QIY@Z0NdI;:;)#FZT/@e94UJ<6M;Ha^]MH7FK](Q_J5cWEYMN3^-[
)BITR2OMgV&FFZ&<ePXfU)_2WF1]g5OFBTEb7.?4;M0\6X5g[S4-,1ddZVfT4UaV
[4;<_ZQ#.HN9GEJ;T^XSYLX.CC]S-61]G,K&\5)ZQIM0M:cHa/U1MO,E:X/JRCE_
3Yg,(c9d9AP.S9b==DY1-0J2P:H\/Y.L>4[AI;5e4U/2R/^^a]+]#:#Ie;W=&/E+
Mc\9db,K)+1MM7VRY3O&(N+,Va613c@78-G]=,eN6U6OB5@\.=e0(9^-E&(HfU>I
N:=9f0\WQW5O[MbV9N>;:cbO2&C_bP+&JE9IF@+gT:54@;\WB@9c&H@dJa>/.I27
;UY9WG2#U2@=XPd^E.ES+H-S?1XdS,D@Vb/VMYWg;Y5/>C;If[<V2NAbaICLK[&N
\;\d)&FJXXWcQe2SEf_Zd8b._.OZIL0+/)9N3N#.J?_MQ:57SeKOH5TB)&6@(2[,
>7/C#<d-TPE77J?d&#5.3:3)E3bQc95@K[>/39\_VTK-(bg^YcJ,S31K(H&&g7(c
&,eX&AgcC>M#V?IY7_)(2ST1/O2e@IR3/\geW<WEP?IIcQ_XJI#29bA;V1D1L<=G
DN._@McOOM856P6+]4<b;BUP#\V/,ARcFd0#VaKd[I6<T)^W.=d7J=I6VbM\QG,:
)C]0g0:4POe4,:f(9S9dG(4#J+RfOE1]gTcd&S)];&7>//PF1c(Sa0e,9H,G+Vda
4BYEH,BeA^ZD_6=QFW]BW007EP((/JUM.7b/cA6E:_E^\Y9Q@JNYg&X1R;_OQW7)
QP,>(^=2M^<6GV:+C5ObW:N=L+L/EM:E)1?3fWba)4Sd\(?\&TFD-Q+:6bg-M8gO
G@0+R=\WfFTAWL_V&5b3]->Xf2NRefE=MNa]8=;/_,X/[IEQd+Hd?[5,f4c.3&MG
U&Q>6(IXRSWJd..aCS9C+?_837UaZ;^YdIU/46&2]_TeSGS<C9c-#8S,_4(FOSHL
/]9NG9=([KW@K(?AB1NR1Q;W0]Y3?g?N<&f[7B@bP9FU2Lf3&R<3+Z2T=@&^Z5Q@
>.K[9ODH-aHE_C&I;[TWfFD?UN+H(92S.GEfKMBGMa1&K,a\VMG19>FGP#+M;?f6
8N)X2c)b3Y^Yd?1e]Q/U;EC#[LbG\S]5^&L:N<C^NT?2]4UJL3V>7ef^2abCeOIX
79A2W17),+&//#\WW/I@)PZJED:0TXPPX24:1ZQaRgS,eE:cJ(O4-/)1YNQODJ51
^^WcK[4W:Bcc(/CL\NN8JJGP6CT_OcW^2N)U<9Zb@I.5K#56Hc,(=U/[4-TTQ-M1
MNHG17a>HCE#(5[+TUY,H3TSWFH&J<RK\1?c0JQa+0;IX6-](9,1;/:YTa&RNe[&
XMNUB&I=T)4/ASF?O(Kb703]N?4I0V9@]8+@PC?ZSO&:\M9Z\?=]0>50aG0f[\[W
L(9\FOQP=)X[5(2>\/D6T7S/T#W7#,Q;fAD#aD7g]fOd-CPfSS)5H2aEAL#U^d2P
(F_@WGdA7B:RaIHY<>H;eB[fT]Ob7G^-G:2\>FT+E9\XTIe&:KQ+<MQ<#E(gCdc-
#N7.])WVefW,=6_5CAZJVB-@5MJS70a(c&DaZFJDIV^C?(^0Zb\1#E0V?;N+fU,S
[+@:6L@Cd>XF#YXXP/+^DB.(@;HfeEM/?8S>0R9P[1g.\EaQ;.f927WD5;g@/-/I
6^,07Xa7MM]feI8CYMb+\QV-@^cK3;X;@CQ^IYTF9KS=M>g16[5MIA;[=.f(?3bU
;X(D@+L4M,02[=1JMV6,SX[0?8eX;YX4/168Te)g.G(bPNGV3GE19<a.,@L(#YcL
[TS+OgEIMAcf5>0Ua+T4H3>6Z)Q)b>bG4d:9?,5?9P,SOc59\V2^KV8CVE2P+Z.f
8WFH5P0/d<82M1)QV1)BEDYOR6O?JLE,ZAK(.L0HLCO7NZZ-@=dO=?GB\MYd59&c
_E0H;\G&.<K)J&\A+GON]cJA#M..<-/G=$
`endprotected



/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by DVMOp SYNC Transaction followed by DVMOp SYNC Transaction followed by DVMOp TLBI Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_dvmop_sync_followed_by_dvmop_sync_followed_by_dvmop_tlbi_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
e3?IcWM+O24]Q5ee/D]38e&APV(BO:;:g6P_YR1TQ/?d?CVNO+bX&)I;B\d0Jfa2
[C1A?^]P\FBRZM]>3]HG_Z1Aa>^.eUB4EFG.7?_e<:6?8JXPCMI_KQUT##[:CD(D
0J^gcJb)U&g9M:ZGAM3VdJ/e5.LE.Z3USf=T[RfR.[P\0W#FAX[851/agQYXc^6<
@#a\L&#K:bU8C\9:^9CRMdSKSC;O?5R3)^X=:6/>[Vg^Sg9/[b):e55S[,+=D7^\
7RTdC/C3gM[J,,cK&eN[Vc;K8SME1E-]L0F=M?eEfKDGeL<e^,?fMb6HfB(dRZ/P
-M?F7.X>?7:Uc)81.,XCOd7+J:/Y7V.G-=U6B>S+4,R74g[79(XEEUPSL_U.UH;;
9dg+Z^aA:aB1KC=cCF>>QM([[-+0M5@51NM;]P=56&__0@/Q?547:K;dVE1=X38J
GNa]E3AMV62W8CXLU&4-1WaK7B040R,CX(_CfJ<b.@/2C_DVZS<D<[H?20<_dE]U
O@-OX:GH;]Y99;G0@FO(Aa725,9J)+&Aec74dbebd6Xdd&B6,/E<]9f:H<cF3,MX
HeEd#XYXTXIf]V^>S-ZQT^LVT-0bZLRZ]RG8g#e.8#>A[CYaZ1FBHTE?\I<;/]4S
(fKRA;51_SG74R?B(][>.JdZMR9.+>2YB3FdH?50Z7KYe+Bbb01A,DTK<6O=@JCM
eR6D#,-^_E&8_VGZ;UE\G@;9\D3&##L=[1I<X^-D3(;a=\DD/LWOW>G)7F7Y9BbS
H^@1YZA[@&A<PWQA1Z.M.+_.28@g@95(QHXLcPK;0</eVST103VND_O,>2M#2I&I
>6aDK+M8K@H1eHY=DaTcLA8<V0/ZgZ<)aF3FHZdF0?g+MHLC/J0X_N?bB&@5XEfM
4e#RW5CZW:=IJLe&VVU44adRU/:0Z;/AfH[BR[bM67.KC4Q;=/8KRae^O7>N3bb/
d6^3@BMb<FLESJYOY4ESNG&Le:M\DM@V.2VC]VAc=##=;&X1OQAe,2(Ye1?2N]23
g6IN3XNgId>J9TW-RO-eK5.A#>&Q-0GS3a,+[JCg4?:aUC&&30A1a:;F_[?=Sf9>
D5588cZg:5gWX(b:#Wb)-58=bDA=)eg/7Y=QV2-f3XQO[Kd\Lg^9D0#PF<8c/=Ef
VK:OR6N=&6e-?(5H6Y5ZCH[-]\eHZWE#0<X_48N(@@+\7b^?U#=g(C4_#^M,7[HN
fZW&HO#V^fQ1]TSHTJD7gV_QWd>B6JVQ(36bK[4@/_O.,g.CZ4Q=X@[?T8)d:1OA
LLX0?8f7V)Y:\0J3;a_AX1IdP#)?4@1X@;27[H5f^()A\f<#-S96]D2XH0CU=81T
Z[a;?^C@6^L[.G_>-A4c)_-1&RM<GM:0<$
`endprotected




// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     CHI DVMOp TLB Invalidate Transaction#1 ---> Cancelled DVMOp TLB Invalidate Transaction#1 on Retry Request ---> CHI Non DVMOp Transaction#2 with same TxnID of #1 --->
 *     CHI DVMOp Synchronization Transaction#3 ---> Cancelled DVMOp Synchronization Transaction#3 on Retry Request ---> CHI DVMOp Synchronization Transaction#4 with same TxnID of #3
 */

class svt_chi_dvmop_tlbi_followed_by_cancel_dvmop_tlbi_followed_by_non_dvmop_of_same_txnid_followed_by_dvmop_sync_followed_by_cancel_dvmop_sync_followed_by_dvmop_sync_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
8<LdL^H:O0S+IaY42M_94-(QF^&dA5bD8GW@gOU8[YfW+5K15F@?2)YNGM=E>]BF
9QfG8cL#&A,c(S-E<Vg7.dJ_^3TW+X=NTVQHRYY5(=X.61CM9PR;WQ@/LM->Z(Kd
Ad>d?H_K3[YS\+8F<795M+H?DO;2+H)(C+>d-UG^=-aCNN8F)edQ4IPaI[aZ<;-=
d)N3J;=gRVSd<KFc5LU:YV;_V6H,]S2T[cYOG;M4-J36?GD^>PQS]?XH,<FVJC-F
<N4=2A8aEZaUE+NN;^-aYb3.ZNHH_V2YV[>]]&OFd:&JZZRGFS#:_1XL4U;8eDYI
d6G8]Q,cUMA\JC3X+G[]b5;FM^NAV<27USC>6ZOHK-e=;e==eb0[E?eXT5UI3-@I
Yg.#M+-ZEC80B:d817,4J>],(_.F)g8dS1N=7-)E7&Qb]BNK,X9[79@O(WXT1P-F
CZCC].0P6+I^L9e?55+^4aR9O1I_cXR/:M6SL:0MRNDP(5E;6ZXB96PgSBe[Ka4W
KL0WMD#3XG#\#+e(&cB0CR,<)aT8TNSDYE?ZIITgG0gBc8=QIAUP[<U>LI>0c@N.
?L;:c2&7]3E=d@4#=e-bM8E&LVg=P\X_FX07C-P+6(8?fYX1CZYH-SZW>gU6M/A,
&K&Nb/))L>4)5T-gHU9XCga1?6C#bZATND3IaJ;>X5<.OcAaAGF+d#^0#IP09\[-
YK7LNIUKW4]B/=@93c=A5T>KVYbODEJ-HXMGL^Z[NA^CH30,2UKaU@ET:7B]NO?R
\bA;6dVU[J#6<[5bWW3Sg0bQ;+KKKYNdV]=,LR8gDP+L)b;TUeWcA8<3.gR:C;3/
WS@GCbRbde<4Cdb=7=25KXCBg;#6N_=6\0-7ED4X+Ye,R#51;QMYA?JU0/@?(De&
T?.:D&^U<4_f6Za9+B^P;KeNIB:M+RKcE3+A(VLN]^_0:&:PV<4(&<c3Rb+7FQ&Q
b\dgT^a)0B2K5A-.EEKaSKJW36\dX5XgVGP.7eI&7ZKOZA>XVESB6)[TT.cA?6A(
?/UYX4bAGdL,5_Y)8T:3=E1G\P:0D<^3_U7^7OfY7LDT>6S_Z&3.Zd=\D_+W(]6\
2=1MXT?JDcNgXC&AWR@:eNH)dDL#HMKA6,&1?ae,1MSD_QgI,IG?/));_#>Kb?\Z
@JJ7MHC\PX&\5?,&M]aNc1&_f6f^]46ed2U6F<\G#Y4^3YXG5Uc?FQ(DK<QV@.0@
LR@_f0g2O6aO5PB.g>>IM7<U6HH1?HU=,[a9O\We8=D8>6eBBT8/&2-S1+C[/&(3
KQPN8R:fP_Gd05JZd]&f--LMJ94;g5@<g6YE.f[F/UY/;?)K.POKE&6^T+Ua@J;#
ZQ.L/&@U;.]E&86[cd1>EA(ZUXgbKHSEV;E3TFYGLD:I\Tf44&XfI8#TcXCW^?>K
bgd0MKI2GZOeOJT@#-&:?AG--BD()]e\OZX,a2VSLI8P-W.b<D]>]HX;K-R(?,>C
D(]2bdaTN>Z#&LSD_Rgbg@XT&(:(13S&UE)B3QcTVQ.aJDU7+0<^=+@NPDHV[0)Z
8P]LKQ22P^,AYHL#WbQ7/B9K@R/K16+2Ac8)XCI:Zf[FR):OI.g=XF:SQ07M1F#0
DXd.CS,[&[<,J]/KWIFXEGI8#:LI3[PG^3N?/1F(UE9bV7aD?;@+2MT[d.-<#2f>
MR=3S_]BcN,;KH]CBS1ZW34;V43\]d.VMM,cECW6.8^K4X<]YDe@.EUWKFA7cJXG
0@EHCB?XWAe(.9YUR><Bf?.0TG8YIg&?)8]QLfaFJXTDTP.;K8D9N<GD12+PEU9f
\ff:6/O/<Q4DCG>;70EW@-]^;6O2__9]QI<&[ad]UOF,#U8)#ZZ1)T:Hb3\dJ<6[
M7Ve5=LOe[@QM_NOe&3,1LG]^&([^/eO]H+[5#eeWN?^&L^[;8W]T;VSI7U<^/_f
+[12HL&\S3;4N\c&H^^[)]aD-0OO9RZ8K1PUU(<6&VDa[aR@&>W]\e60)QF2TNQL
ASHQE0W,<VDH^XLaBabOD,XDXd3B;4Qe,dJ^bXWH1&=DB]CDV4V<e,.=8,&8)VN0S$
`endprotected



/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by CMO followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_cmo_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
)M_CY5Z3A-e2^3J^7D;bf:4X0&JOC_b?&FGUXc;/-Bg#NNH\g;\E+)06R<JI57\V
+8M;=.P4M47:294RbZELCN4f8]V5JWX&N?^U1AN@Qd?bSHWE+S2^)a:1->]TcDI7
XM#K1),G>)T^35DfN@M>LC3>TSA)SCA[E@Ee(9KK6/,9.CE.d6&6/7?RB<\8=&K9
OC7F/5fd1^_4\+37<JVD81X<()CN)d;NF,FZeJb4WIO9MDdc(Z[&NOMZY/gg_5^^
JG<aT<IJKV1?,2-g4HKf<IK&V5;.5,G,]Z1LJ+2[V-JCLa1&3H5\)(SMLaVbROOI
U7.R4P0RDJZ1Rb@\):Q?8baU^X18g,@L/30a;e1=e::ReH14T,VM)DX@0A<V<0fE
KCH6]e[TF(BT>8_:.Z.BO=g^SUb(/aaN_/\)P6<_4\TZ<VfCM6ML5aRGd>a.)0<b
+)/#]6>;ZB]<d3@4+Kd75>]GNFHQbTcCH1R6RBdORR@G3bHX4e/HBK<HHWWRN+#V
:S>Kc[J9YF):7E>e0SAEcXK&ccL]9@g4e&LJBgVAZ-Wa13#=d&RX\/WQG,3I+(_a
E\,_,cbMg<b<SfTeH8WK?H1DKQg_,..P82;D_KRaeg.MI8?P5:W4^R];3]>8TQbO
=#QAWgGg#[@HJTJNSae?1P8F\7D12@RRX:ZH=DR-?M.;b#4NSFAKQ>dgW>dC4TSP
VLQP8T08T^I2fH&WW54SY66)]X\VZ<4].N-L7:<6Aa?1M(P@e2030)P4fQ)I38@W
7GK@]Wb(Q1MM8NEVQb.73-2b0f=SZ1bbB-YF0C.GR\/K8OfQ4KKA?(4TR=Zg]&9.
QT3.b9IE+N5:1VTRNAbKZ9H&9<V\@?LQOb,5GXT1]d(4SKKW6OV]WZTZ#\3Y7E5f
=6W@-?V]>YR/0-DeZe@C9G/N:M)KYBWQ)KET;U[fTfHBIUV0?X9PWJTZI$
`endprotected



/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by CMO followed by DVMOp TLBI followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_cmo_followed_by_dvmop_tlbi_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
.-aSG126Kd<OCQ-b#WFS:-AZK_UU)K3\XXG>2:U2:g,IbM+/g.&+5)[a,bJ?bKOV
f2=:1TB[M-4[W)U<<1)Q+AWSbY1(LeEC?M<)&MXE(Cc?/N7HGF>,:BG6C/D+HMOb
?6Ob-=KdRZ@3#K/?9DPY#5U<GK91gC_eSTR\B]ebSD.LbS#CaS.3IB.N(LCFWEe/
,QIM7fP@d3QVSL]?OUBcERCJGK.ML6NB_Y\OgY+(eV>703HER2N,U@BK3f5Y>-O?
#C6J(e&_K-.KK@8]]:/&gZE.MgZ]dR/a[D8#UEe15cL(XHT1I-B4)d^#U;,NaKUD
V]T22gB;+5D8T&/3gC((LZGN:eU1)B]5T:c9]J]AN_DRC@(;B1\TY>@b?+-Q@PHd
S+-dNHG\>U7)56I_>1@OF0)EHC7+;:J&6_8UMSa42F<dJ.)gX(gQ:8UFcC@cgb1c
CF?34O1f9<H+C-D>YIU6Q5[#e.5#fC/e>M-Bc8_XNN=(&ZZH/P5S#HEbg&BJJK/U
-eT(1@6d21<FN>J:PS)(J28<F,W4CML@gP)_,)Ia[bX56MTe2CV:R:#g4(0(=KX_
CAdWA4\I,+:DYS<Q#IZ>Eg37HU]SbW.R]dHMF/4278>G?I+USEFD5_KZMZ=F?^E6
8a]@QPb-])4/O^(3UG9&bYYdeQ6dX1P_(gTaIdD;;0cHH(QO@S3?M2@,fcN:602J
LbU^>(>>/SO2fcFO.dYC2W&?CbD[RFaT1+A^2QE(M_@]Y5)]U)A#^_D7..ELU8:>
DQ=]/OR^:;YQ&,TC91^J8X^/eDHY)f(Pb+WB0KTJP06c(eX+>3DDA7H@OF4ae;Z@
@WL\P;K5XfFgM700:K8Fc1,TPI>>7@-)56B#d+A&OT@CG-P1Be5MXWeO]4?f-,^E
Vf;+3WAIcg-QO1G-\\ZCG;7V+bPHWMe>PEW97Ec[:fQ_F?/.^SD7+bFTMHegGd43
4Of-PYBP(5&f-D\)c3.FQACD?A+K7>25:0+^&PbHW+K<?)3d_U5Yba^4(TQ7c_0W
C4#?Ce+LQ6^\S(^TUDFY<:JK>^AJHH:fd-N2-).1=@g8.S)1UMc=C))9,3cM8[Y3
/4PVATFJ)>bP.<K16T/?FX93^MY+QVC+1@2bR7<P2##H+E9L4Zg///>,<--bP[]3
PNJPS[^O6[1J57DO_N^b1Jb2;H&=-QXEVP_P<H-K_L<c4G_7cf-4#:\NEO?XPAcg
FGYX@,UK&KB,]-6.IHJ.Q-b28$
`endprotected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Load followed by Store
 */
class svt_chi_load_followed_by_store_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
#3QJ]AELHZ_,R3&X0=)CK;7Q=eN];YNOERF25))YNW)AHTPSK-2G5)@(WIU(Udg7
M[+b?6c#A5A>e)D)UUWY^;^7?=;=Hb2UdegD_#7+&&eQDK2V8-H6?gd;IH1-7H>Z
J_/N/MTJK23fAB3S#a(^-;Z3R;D63b<aCg;]ggQTJHQ=g3acaRF]@?F]ZZP[]d2M
#=>\,(3&5BNREZ2]a?;M>P=e?8c]-.MaIf@)C>DdSK3\0KXUC6P+2f#BF6O9&HNB
,1eS0V^?1DA(<FVLOY:(0Qe8B7(_LI&(W&MWT?Te&^&#g8<GG)T@d;&W5YCT+;(J
LI<g,>X(,;_IdR?VeA\g-@@Q-:>O,[=Rg2^83:^,X):g+9d<cFd5Ef.K5R]Y@L5=
TZ/J9@8a?cN&++:P@HHMZFUa<ES7;J@8P(5CVRM(dRPfDJ<I-@=D8T^_\53gF:bO
Ne]?/8=N\R&63B3ZD+-9\;S_K.J5?:U;ZCg27;IB67fI\]7MG.TUcO^O#_?>(#1X
17_c5)MSP8_Y91@gU#fE_6@ac<:M(JKJ)-Q;(Oc,VT)ID$
`endprotected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Load followed by Store followed by Store
 */
class svt_chi_load_followed_by_store_followed_by_store_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`protected
8O437aUGdR^#g2?aKc.8&17O_=d]/<V5@;6cT:1c8I;L/0]]G.<c-)::KH5?CX<M
^I)J0;>A[Z64a\e[(bB4QZN?,)b-W=V>7Y@)<@L=TE:;10WO9/LBPe58M]bXPA9a
E)e0AX7UKS(aW2/R?:W)dEHQVISSK=.FDO:GeM<9><I@b8GGMB?#P]1^T_R&UC0B
0GW>/^7EQYccgX-J/Dg5C<9#O#B&(N3g?A)I#)RIVbee8>J]7HHN-@+=:>:@_aQ@
.6E/154R&.VJ?HR<_9+LBY;FeLKIIaM\=6V(:PCK+D17KUNJ>CYgBI^C18(g^NE4
3.HbZ>6Y:2acK/R=&SU2BE+Yd12_QK@Q)F11f)00OA=/GV:J;;.&;@U6X#2KC[?W
6&8/cS(->+1CHa5^O#I/7b?dc&Vfd=XWfUN_I9,-[+;@4Z2N@L1ZHOWDSXY4X559
YT&=acYe>[Ua1#eQe;(4IXLKb/a0(]V83[YQ(^fX_G[FaXSA:XLYaYCO)ZDCE)?E
KR^.CaXX+>^Pa3Q4bX>]CN-REG@=1+Z&X/UN&#]@.N1),c7#8_.I7YG<+:XD_&DH
)SGBc(&Cc0J8E3-b6(@ZQBLLVJ)P+[V;YFA=I8<MceIP2/Wb/G4KMOK1g-fJe/JE
SR8-8fM43CK<;F2-P=P[@Q/]T,L1=c5UbIOc8V7G.U=CJ)IV,?fG4J&@]3C()bMe
WW6TX[=8,G_6NML\YJRC#JKcQ8A^..WAG98>6P&UR-ECF$
`endprotected














`endif  //GUARD_SVT_CHI_SCENARIO_PATTERN_SEQUENCE_COLLECTION_SV


