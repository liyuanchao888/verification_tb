
`ifndef GUARD_SVT_AMBA_SYSTEM_CONFIGURATION_SV
`define GUARD_SVT_AMBA_SYSTEM_CONFIGURATION_SV

typedef class svt_amba_system_configuration;  

//vcs_vip_protect
`protected
L;#AbUY8A9@egLGZ9[I#DTR\D)Qg?2>4@&GS.NYEJ1=cAPK.MM;:-(V]NaI>NY4(
P#9>PN:(V\62,Cb,SM#fXS7b8#U.LS@=_Y-D]T/8FS)Pe8RW&Dd.B,R:QW6H>//d
ZbgRJDaU/,R\I-c_W;#^OFRGFX4[-4,Je:L5cf[E4_<f7fLL3<8dLJg5(d:VX6]G
V8aGS2VMc^48DOI^1Q&M>Y#^:FQbg#cf,?g:@O_86R2LH.Z^AS@43B0_eDFUN.4H
]&1?g_MP+H0Hc+[,e>(CNcIg7DHff(2XZdS+Xb[Vba#cfT?D#U-H.2]#E[d<(T6N
C?8XeW&g#Z#K^IB4Q4=D;YL7&#XF_#^N2G^=>,DSF6+.CIY_+=_+TG5TW[ONAMBH
d)3BfW>]8^;Bdg40YfL(d&4NT0F-:MFM)V:eF37K+WI3WTdBT4G.GYb.fYOAXJZW
cb=ND52=7aLZZTD6RDa/?T2BXNJPUZ:FM=Y0)_V;#,Q6C+TYPF34NM3N:8:&<</(
[?Y6@PZYeC7DYDRBgZ<,AV72P7UHKJe1,GQ0NSUHO4.55(Y+8?Qb:<G3T90P]K[_
U,[UQPF_Y+^R&D9\6:K5H1e),G4HSSE<::4U&M0D(+..25U5Q;+2bB]E-VLN2Q24
]1+_bSdR,8@9;J.UNWV,W2+;fSQ@c>fR//DZO3-1/[2-JRNd,CcZ+6#0c4^,,[&2
VfM.(KTPYHcU?g.F<0a<J9T97OLG]Wc&87fK(VNO:GSZ5]Q684EYOS1CO:F\^5UL
TaA;2?3H_9H.T=<dR7U?F3D_Cf7e9)3/MM5YUR=H1V/Bf5ZfM)+[?5C5F;G0d[2(
;=5^,7Xa:P^\7b5&A^YJH#+b+B7T7=3bP&#\ag#F<&6cE::dBV1HgG^PCXdU>#AZ
^D8@,VK.)R4PG+ZA,^JHSU4)&<E6T#/A,TJYQ>XH6Zfc;PVcN)KDTS;1J17RE&C;
O-;TZ.L_gN>OeVPf)5^U3WDL_b@J>g(HF&75[;f:ZKQR^c_LM1()LV:W:FU_305d
(LNX=aUV:SCY9>)7RR/@Y8>SSMAU70K^D6f_bLISU1Z&^36YL_(U7?IG1[Ud1.5M
T:-7Y>VDCPXS#_Q(QJG+4D5MfeOPcGFf^7NecGSEWUJ:>\0&638M:7Kd5/b@6\a2
A?N2)_>.\Ee4O/)Q&IDX(<+d^OGZ5RVI4c9#2A.X#_?3O-0NN<:;3I3CR1-JdLJ_
K0/d[72L&EDS1<?]bC(&<QMK8DK/BbZgd7EX)^2,X_?=N&-T7#-?ZP5OO(HRVB7O
056WQ5WT423QD=MGC+MVf;EA+ICJSSZE(VEd;S-6N7Yg[M(?7Y9Lb+X6#WU=b02(
gFZ>NTX+3a/^F+UP3Z#XaSWR?0ZZ1DQ/5MY>589DeHUY9?8gU]XO2K[IDAaN<FN7
KUF4g>W<;+[H2fBWFZ2016<Z4A4/34.U0.>>=K+]FZ\JQ7,b>MD?XbKXZF(.45E2
<OXMU6L.[:=.6S&._2/7edfQTNg7==&T>+@WBI7bRTA/H.Y1(Q;CA/9J03=5JP+I
1Uf4bSaWVB>F^/M8=K&+[L4W<>M>cRN=+@RC7M.;0aEfZ1]U?O0.RXD,WT9C;4(X
\RC<(7VJ&+^PB5SPOP?Ve2@MaG7[VF&L(3K>fd,B-^6d\-MA^__3a&\]=LE]Ke@d
]DX.1NZfUcU4NSBMPbQ1,W0,KQSB41],2A]W#8>_2Z#\54[\+MO0GUX.0>M5M#F,
M.P>5OZN_1PHZ04T@7YU1T>SVN3:YNg_F?=<->.JFZU;D7b?PF;4GC>\<:=WeJ+5
NHWRCRT?-VUF?AU87)dZ&cf1,=^6511baP)QSXILB574dLcM7>9DfN.\d=TR^#B^
P>aN@[@TE-^T0a^^9(#]XHIF&]=;dLC&V>?=@/VbRX(=Z=a+MYW;GIa2Z@A9N3cG
f):]IMR8H4:/&T[H0gM9KQ4^S&O.ZV-#<EC/^D9X2IVLIbN._5P9)9#SQD-NDJa;
dOW6,72U[gF?3b(b\;5Z:\b\ZCS5_T?Z+05&=+aW2H\(^;@0UM-fA9g;?aAIa8f;
gL2S)I3ZF#0cW@=BF:A+H=ZS\90RH2BBd+_P/JfHYbI/9NR4A6,CH#@Pd>F&JVLE
<]]&-YU;a;dMKg/L+\=_\V[C4gV](1Q=N2.NLI@fJYe)/3CMJZY9-.6dZK)&gDP,
6\ON6Wg&:,-^NE-d@)Q_N/e;M)=,@dL?M]D?\OE015>K-TgCB/[9[aZFH1g(W:0T
WQA/[-U&[e8YKSI--ULT9YL,OaH8a1AY3&/Y_8_aYV23B48Y_Ge=/)6HKKOd:[.Q
7:AB=I-O87.8cJb4RNFWMA[+5CQ7TNMCH_3G@74Z:5@QNXMfb[??YP[#RY2]J5M9
>G59LAN_d+RBW_cO)AM#F.Ied/JV7X1-+R8?:#E1W<VI&&Z-9?P1X@JOJE::N7]&
:X)B_L/ZD5Ye1>[E<^6LR<FLGJ1G9F-Tb/dXZB0(A<C-0L^SV^/EY;2O?6M0ZYCI
L0ND+_7g5+PLG/EDQ<f?I2P]ScV.+f1K3QVU?f?R31>Y;ECCAeVYEcSX&W47OT+.
8K#<Xd+N?cCM/DU=c2HT<S=JZ2N+IQY,.84&\@[I,Z#(2+)(GgeTW.g=9b:DW(81
/GFRN571\C_);=S9Zed>8],@PZFE+H9(Nab]J\6?d=F@:Fe2#+,<#^]AJC-LFC&.
Z2IQXP(=efZU6R96cG86N^LHI5-V&ZPLB;I[YSQRD=_U0T.>6O_X<8=Hbe4,VAVF
PJT]HfT^+HWeUd19GVG1NT\=66S:fZ:^EM8V61_169G?04MZ]69\<f=HJ$
`endprotected


`include "svt_amba_defines.svi"

`protected
N9&;E[f,3#:FIAe77^-Aa-D_.VO)Y+VVM_O6:5ABB5R8c6-7KN[]1)L9NHB>8aHZ
24[@MQK&I:5V/6\MU-X7:IPI>8Z(Sb;&8H]5+fNP,)^Hf1;c3:#V#:3Rg/3J?QH_
F@[07T7W.H,75QA@1@SSfJ;NbdHF1g5.cNC463;.5(<57()EFI/W0dG1NF#Le\HE
adV?#W5;RS?^f1d,M_3gK^S@JcgZbC4NSRG^OR=bX(JGV3?gNBU.K+PCC:[<@@73
IY_Z9,cSFL?_VaRLeJ:GfGX[DK.).<2Y-@OfIR#OSVJ]@H3+H7:Hc9F=SFe2G_6H
>@V+a7B;/;DPK.@AP(5)De)FT#NR;ZR..Rf/?-9IbZ;1;J@e>+eT6ZFN/,LdQGU,
JI5X_Mf()A@d7LPDX[1+F:@IeHe;deTBUCE_eg\O#CR@QebfM4\#e[7F[236,1NM
5NIY<<OD/(Kb][;V_:FIQVN;^=W6]:TE\ORQVM]1K99&Q_RG9:SVcc<e=V>OaYCL
JOe28e)Cg<ZH6)SI+JX;7]G)F4TZIX54YDgB2@E&e]OQ@]3c[M?L#GLTPfW].b@A
RSgcZSBFfT@T?<S-.3J291;K3,B0dO\8Cc5T3gQ5)M(/O#c=_RI<-><Z+LWTW]-Z
LYA(aJ.ee.^N]Y]#+GLM#@G8Mg3.[\+CTeIS>T\.G(90BWJ,?3cJaaOVQV8[6FbN
DAZ]P#g-8d]/OXHWAILM&U(S42Cb9ZdB._dBabb=Od-YY]@L6^ZTCB<&8^ENRHK_
>BOB&Vg-=DQGB-fE_9OH7aOS.0TcdQc7-1CgVIYV5SH@_Fa9PKL&_Q<f39859[HN
JN@\9K-fKRT<40D]DKE\KEPB^5,?+R?I(b7dYV6dLU#V:b5U95DL6?V8.8YOG<fF
9Y/R^2I+Z4@G.5Y-KE>D+YPB1$
`endprotected


  
class svt_amba_system_monitor_configuration extends svt_configuration;

  /** 
    * If set to 1, the system monitor issues an error under the following 
    * conditions:
    * 
    * -# If the AXI/AHB/APB port to which the transaction is to be routed
    * to based on the address map is not specified in the downstream ports
    * connected to the system monitor.
    *
    * -# If for any transaction received on the upstream port the transaction
    *  address does not lie in the specified address range configured for the
    *  AXI/AHB/APB slaves which are configured as downstream ports connected
    *  to the system monitor.
    * . 
    * Default value is set to 0.
    */
  bit flag_err_if_addr_not_in_range_specified_for_downstream_ports = 1'b0;

/** @cond PRIVATE */
  /**
    * Applicable only if the system does not have any master where
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    * Enables the AMBA system monitor to handle posted write
    * transactions. A posted write transaction is one where the interconnect
    * responds to a write transaction without waiting for a response from the
    * slave to which the transaction is finally destined. When this parameter is enabled,
    * the system monitor disables data_integrity_check. This is required
    * because a transaction may not have reached its final destination (slave)
    * when it completes at the master that initiated it. To enable data
    * integrity checking for such transactions, the VIP correlates transactions
    * received at the slaves to transactions initiated by masters based on
    * address and data.  If the VIP is unable to correlate a received slave
    * transaction to a master transaction, VIP will fire
    * master_slave_xact_data_integrity_check. Note that it is legal (though not
    * mandatory) to enable this parameter even if a system does not support
    * posted writes because setting this simply enables the system monitor to
    * correlate downstream transactions to upstream transactions which may be a
    * requirement even in a system with no posted writes. If a system supports
    * posted writes, it is mandatory to set this parameter to 1. Reporting of
    * orphaned transactions is not currently supported. Orphaned transactions
    * are those at the end of the simulation which could not be correlated to
    * any slave transaction, which indicates that some transactions did not
    * make it to final slave destination. 
    */ 
  bit posted_write_xacts_enable = 0;

/** @endcond */

  /** 
    * A back reference to the svt_amba_system_configuration object in which
    * this class is instantiated.
    */
  svt_amba_system_configuration amba_sys_cfg;

  /** 
    * The upstream (source) system port ids of the ports connnected to this
    * system monitor. These can be AXI/AHB master/slave configurations
    * The system port id corresponds to the value of amba_system_port_id
    * configured in the respective port configurations. This is currently
    * used only when AMBA system monitor configuration is loaded through
    * a file 
    */
  int upstream_system_port_id[];

  /** 
    * The upstream (source) port configurations of the ports connnected to this
    * system monitor. These can be CHI/AXI/AHB RN/master/slave configurations
    */
  rand svt_configuration upstream_port_cfg[];

  /** 
    * The downstream(destination) system port ids of the ports connnected to this
    * system monitor. These can be AXI/AHB/APB port configurations
    * The system port id corresponds to the value of amba_system_port_id
    * configured in the respective port configurations. This is currently
    * used only when AMBA system monitor configuration is loaded through
    * a file 
    */
  int downstream_system_port_id[];

  /** 
    * The downstream (destination) port configurations of the ports connnected to this
    * system monitor. These are CHI/AXI/AHB SN/slave configurations
    */
  rand svt_configuration downstream_port_cfg[];

  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the configuration
   */
`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_amba_system_monitor_configuration);
   extern function new (vmm_log log = null);
`else
   extern function new (string name = "svt_amba_system_monitor_configuration");
`endif

  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_amba_system_monitor_configuration)
    `svt_field_object(                      amba_sys_cfg                             ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
    `svt_field_array_object(upstream_port_cfg, `SVT_NOCOPY|`SVT_REFERENCE,`SVT_HOW_REF)
    `svt_field_array_int(upstream_system_port_id, `SVT_NOCOPY)
    `svt_field_array_object(downstream_port_cfg, `SVT_NOCOPY|`SVT_REFERENCE,`SVT_HOW_REF)
    `svt_field_array_int(downstream_system_port_id, `SVT_NOCOPY)
    `svt_field_int(flag_err_if_addr_not_in_range_specified_for_downstream_ports ,   `SVT_DEC | `SVT_ALL_ON)
    `svt_field_int(posted_write_xacts_enable,   `SVT_DEC | `SVT_ALL_ON)
  `svt_data_member_end(svt_amba_system_monitor_configuration)

  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);


  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
`endif

 `ifndef SVT_VMM_TECHNOLOGY
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   */
  extern virtual function bit do_compare(`SVT_XVM(object) rhs, `SVT_XVM(comparer) comparer);
`else
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare ( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );

   
  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();

  /** @endcond */
  
 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the APB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the APB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif


`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_amba_system_monitor_configuration)
  `vmm_class_factory(svt_amba_system_monitor_configuration)
`endif   
endclass

`protected
Sc\6?<;#6JeUIU<-e/G(9V=E9S1QffB5?8bO^M[.U>DF>G\OeBa]4)Fb#KMB(L<V
^>bXFa#/=;YO1PON@aICWfX^,H#69X#D[<;Q4I2,:C78c,E??MA:^@.<0_b>cQI-
3[66SR:/7F?56gd_aBgJUP\4-NS_[=/IaKV0g8_;_(-\9EOGZ2f?/W?BFZ(YL(GL
dILb)C@IB&A3M5CMQR.f/8F69_:&^##BE5eA^:ceJ9?VGA(7PZJ1I\,+T6V;H3,>
KRB,b]#TbJ0eaW48#AS6A[dbIZ_X^a=)O&_=YF/d3V^6,dSSHJW#\URM8cI=;GJ2
A&U?K?g,=K^>R/^1TI>WAU>d,^+McVMNX.TLEb@5.Jbe_,W[_/E+.]1T4W+eH//0
0AbG9=-?,UG^B9BW]OWFfA=5IQY/KRJ5Tg@TG]8X5;?C>03YF>HJDPeN>(<gVg09
#RA[\TT+J/VO(-R[2BOLbUMX&a.Y[_?UGeE#YG>V3PF+W_.C00GS-5N+8#@S4P1?
FeCNMU^G6X#?O3)8FST;1>(SVS66^3AEF.F)GRF2;0.f)gX97=Yc6)8Rec?5g2TV
+d2NcJM3dE<#T^Db&):W<5.^?3F=(EbS3EYR?>g]:JgC)83()3:=-2N=)bg7XW,I
W:@3G7@FV@V4[bQ4]=/@_KE.RbWP#N2K5:X18L8O0^&?#VH5e)^E4@?T^9BOJ]MJ
ZFC\SgSAb.?4,$
`endprotected


// -----------------------------------------------------------------------------
//vcs_vip_protect
`protected
R(R#E:@T&/#1cDYd?J0G6\]ZO<QK+d0&E]SP167cRcXRC0YF](7Z5(0Z0-QadKEV
\258THCS84MaZfSJ<PLT_Q.PO=@;7(Yae<,S68>;@^fG3T7fDQC9VF/X_PN2;-Pe
B-g[;=NagG/3/g2;7D3.JC/\4LETe-MLVbe2+]L8+)0V)-\JK9@FW1+cg-7b7^,R
4B;#S:5=D#2F?DJ?E?gd8)_1c^[BU7De&,ae=:+S6#Y,LG&)4\)EEC2?(VH[S:C[
@+P&3]Pc\^O8LH#290deU)=O]HOQ6;5_7gb@=(26WA:2gJ=-J(<M&?bMBV+&?^_1
Ea36B5G1fe>SL[?^7Ve52[GCP#0Q:e+2AG&=UEX=2(08Z^8KMKB<YAGYB9U#a;]H
LcCV<U^HQ?=;1JX[@O#;fS0JXD<fJ5VMf:W2VLGZ:eCNdf=ce3W:2VbQW2450b&0
TRYgVPeP-#NMT@30Q(:#JC=HPC+@,RVEU/KZdc0\LM1>0+#EV3_ANWXS8MgK6^#:
1DS@.:LSVQd15XZH0S-Sb.O,9CJQL6M^efYR4Ua+Yc4c\5X(ZEfW-?/W)3?:Naf[
.5AKJY>8/TS[(1-QeDc+G@7IRgf7K8AQJ_a/d:+#EUe-.A;#TAC=_OG+U4AX>@)#
910_X/Ta3<K:C>aNYU=_U40</69?G(\(O:ff6JL=M&>EO[@0([RfHI9eX8P^g3&M
a#@C,H/JVGF<[_8B#7]c,X[WbFa)DM.(=d3fB33?a=JIMCR<g.SW:-@B8F#0^VVU
L)(KQDLBF(;3^U8S4)f7R#6^5(.0-L[M.M?)NJEULIUUUHXD]Ud^E@/;6g73dM0A
X;H;7:,Tff-6Rg.&).Q3)WG8V?HSLD\aP&A;g_),/E)P.?XCD0aVEVN,g96BOS@P
D?cQBb+^8+<=ad>bC(EZ?^_TN[#c6.;DGARKJX?L:^QNTcbW(T=NG^8fPbbR<N?5
62;XKA9M^gS3TfCHbP9MTYKL_O@;Dg#L_dDM#RM,+f@Z@Oe6BE4b_E\O&O<ETJ_8
7(D>OCgg=HA;eHPZ0[UGT5Af&L)2^.WJ3Z6L+=/=baSTE?d+EC6eR8<BMN\-@]?\
>^R/:9_aX5.3<Z8KTfZS9^_0FaK?RGP;/<KWeG_:LNcIQQ:Jdb)5C2dXSHR,UEWV
5;bHbWT0WZI(GA:Cf6N_I@-W2aI7OR\A--(T-63;WU^^,6TEYV<LX?Q.:gE:86T<
9?cRe):P^Rc&HD_AWECAPeG4O/VOFe-EIDT<8#^N>HLZeS8EN)V5WHY8][/]1D77
BH3SVb&VQaWdCEaH:,\TH(FKcg4>/G]O;\,=Re+GD)RG4K+6=L0d4[8G?GYL=Ac=
K.8:X(?^SG7MLG<OP\[5/73Y=A6AV]3G64-)V[WU6DD,+]1d\\5]2\6J?\1534AL
)](@#1b3P2>A;RV<V-UF6+>N,L^F91>UWNE]aXQe;\]F17_G^:M:&24O9]Oa0YMT
KN986f,JO)G9X1beW4.2?cZ2S&/=(IFR.[=-D2d./OaEf0HgE_FZ<S];Lb+Z5711
@^^^CJO;^f@=]DV):^5Y]OY@JQE3Q)IWT;f8T1I5AZ1_6HD,6)dT(ZZAG:[HO\Te
#)C+_[@CCP)<[;0\Q4NTJQ-\1ZKKVJ_,H4K#+K;A9^KA0?TMB^3OQD&S<O.O7V>?
BBRR^g9#Zd^(\79@#R7dMaPOZ\J(GN@?F+#<ZK)X01Ce:fI-;FX3c\ZW^)ITe);]
VFVIBd/-eO2,GPQ7NeRR@Q[&;8X=5L@\=KI.QR_;QWQXYCgB=:>F4M-N,;AdJ?E.
3#ZG4bD]geG6F[fD<ZM#UgUbT)_RN34RDRZ>[Ng0H_;3PU-b8/HA&G=W6)&A>?IK
U5MaK\O.4Y(NZVOT=H-]+=05WbVL4K+dPeZ@>>@Z)g:QH_=8M7/\\Q#>H#cCSLJ[
g^]>_1YU\C7^^#b@,ET:]Z/Y:1T),O^[W[M(RT<3_J=LMR=:=_9HW[BUCHW@D)E?
]A#/#L6;5ZU#^;T#.<T+LHT&b)IbgON^HfJ,W=(&X3<Rf-V,7MJ:=Ie+gW?f;#Se
XKPOXPDU5e0bPV:We+87f_MT>e/AgbOaH1J9?#Y&gU.2_]&.>@V;UH:#CS/&g^9?
>7[0P0RTW]2G-AYg.@>cJ2fK.)]5]F9V+P+ZXdg[@NS[C9-.&5FR>PV34K8BKO>_
)1INfNS?UVM1J/TQ[H][[EUF;H9=@Sfb3S(#>8)QEaO+2Qb6EPO^,.+M@=Q_85A7
;/.^I>[]dX2LI7^3Ne/\H^gffT#-S;:76U7N[)(E#UNf8)_3DedfN-FWCIQ8];=f
_7&/EP5PZ(YG?Q4#0cN9M\Ec<Oc/]+X9LR>aURdWV@4I>6TRS]5:<Vf3&9\F5/=Z
2/+\B4?PN\=C)G,6(Y6RgMb8SC7]9@MJ5-eeLec#;HV7M5-6fCTdCJ-OYNe4K9,X
/-W_VQIS><--f0]9MdZK@g@W-ZMBQEZ05TF).U7YNdWg806G462G-FU7Yd1/fL4?
L4bIQW2\9VM;W[-OKI>T\F:ZgQRCJ&QSeZI.=_:_B8E<1<D4BF5+c?GVS5g>W(-C
9RKeR>Z^WaS-ZJYXeD)DH_-A[V>\c[LOC^eVA;@fJFXd(Z4FcI5^,f&+P2Z]K]?5
>Bb-J,H/&>8<R6/AIG)AHg13Qfb>a#&Y1Ac8O7d^<_QO#,PPSTe2--fe?R_A7D1b
IdNF^-L88FE:_a.&W9J?K>[#&BF>TE(R8=(LRG:78gL&?97,5\(LO.g9KB+^N[;9
EZ>C4W>T_YccJXg^HD\S5GaLZ=b.QQ4(&EM/^/b#=e7S-b:#@]ECL+07I(d3Z26K
bNO=Z.PcdfP4.gbN>XV:BbQ?g.^2)_,d-)aRDXbC#;&BC#_eB=K2Odc2ALT3MCd1
e?@[V.;6<a8E,Z_&6]TQE#Y14LJ+]0QBR^aZ)03A24OG4_>P/LHW+S6PMJ]=C-Q)
2,aOd<d9#;DLE):X[B.aQJ0/eCDH=0.fO/HTL(DaKBPc(6FDZJ(MCaD=RVe?1SM]
J=&X>LYB-G-1J2678G6E//@[FSS(FSM]1@M]X5OG388[=N@fPTdQXOP#X=YXH/_J
>3@_MB#YQORP-f0>2&A^10^c>@ZMgG6IV1-8c&HK7B=A,VJTfL0=G(52L_^VRZ:X
FFKOAP3R&4cM42],9P_14ZF@2B(TZU,bNOeI#9&e1T7IfcY-3Ba[Q@I^(5((X_Uf
d(&dK(H3Na^P.T]e=B^:HA3&bFAdGe&2:/RUPbSSQ_\a2(OAVX8^N55BV0]?.bWQ
_8]gF4AT#F?SW-XK(PZOQf3:W6_<.S,b_FQ26d<LCYG#99([Tg&T0)-I@7=>;aZN
/=FYbVK^g;eUSH2<9V@MM\70DACfJPF(_UOHTf8cG7L[dQ)5D,]#N[1]U+@^DG&8
I^JG_K2@-BAG#:HIA_>:5+If[3GMGC7(L;f3X8C7\6B6:_BXagf\eTbA7F;4/aKY
Pg@YC4.I4-<_\Cg2#929.MMGa?MNKZO#5:SRB;ZM8GW4\[7+PCcCEQA-#+<DSUV6
eW?>b.P3+\V\6Y?(@fAM8fQ8AQ&D4&DKbJ6+KU=U&QDP]S1>DDcc+&_cAHEYV/2;
0a:fP4>22^@91g2;K)5O@>d[NDWaO<16X_#f_C,J=EDDGSK;5Se&H_[^_BR:HL?7
IS\O#<^bD=,U<6DI&A8Q,(FC936\>SY>,G?c;A]S(]1R1M[\4239Qg.]eS;bGK_>
2C[?I9cP+4_Kg/.=.W/,DE0C_/<US?L(ee1\,Q8XV.9JQ@Z^W?(SO68(97VQL17B
<2=FM5B.Wg4Q9KO_cYVC8MKJK5M8B][U>5eZ:C8cCKHf.L2IJ)AdRa[?#3b0Y?[G
Q>.[G2:JP[PeVG<TcV>[=H3_Y3,+V_;5OPVe/_BBUV=.Za&g8+PD9KN,QI/5:.X@
cB6M-KPLfcRF=TaXWXRVF4:>.)30G@NX-@C0;eeH3X.ZOT6.NEg(#J\7HG[1JOCa
9eJT5P/IHXTJ=HYD[IK##VQ#N7UF&dJ,J?)OP?V98@5VF\f-HUbYg3;5Z](4=VVA
#6JYc[]#dc9,HDaf]dS_MMJ0TX>g]a?IJH&e+.MX#9ZJJaF\ZE+TbA,RJ]_&K@>X
/A#8YK,9&/DUN:>>&A+U>Bf@G2#-;dV^JS=bN/_IMIHa_NCSCSGEA)JYKDC3V\>^
66LY5_If;4S\.F@I1>/U20D(_,@\^^FI30C.1[H.f,+aD)c;g@[:<CG&e;GYJKAF
N2PLdA;J<A@Z,a8QWJWYT0ACKf=C,_&3,2-HG19e8Q;aPfA81FXQR6R=PVR8NVIP
^793FL]WR=U23OH3LG_+>8)2@F5F=gB4#QJ=W?MP_QaRHP(Ng+<D_35K.@J7R+aC
8Q/-DBff8AS7EC#SIf<[6J+YfbC^MJ65/.69D@8MaTW1NG2?]:(W+ZLB;5BOX/S@
2\O6RX5E[M\S=<7F3/P,)aT>KfUM19K19B=AcaH@/(c,CP4,=G#9T+NZH.XIOdRJ
M@3cLc@IY^;7A5]YV9P#B8742,.YbG:?B>LaEGab\-f#S]9GC3)+6g[[fN0B3U3O
</QcWK\Ke.3T@5VHPD/J;53O@?c+MEMW?ELR:0=+LRdZc=@,\3M?+1MN?]@=L,eL
LfCFfdDXBWDc(M_EO>Fed1_TTPD<V@/3)g1IYYS6Q:Fc<E6K]3gM@VCF:/g&G@&X
39J:>#6,_58[FGE\/aNE-N#W0)MOBa,eAQ]7__<L?cB+bgIT5M\+A3>1L5.541He
@ZUaR8d&9,A:KK-OZaKR9O2/B,?OY=#JF=3&T,OH@fP&O5E(>8.5RZZTGU55H8IJ
;Y=P1O>BdE;O[>--(JU0GO/ggYQMFC&]e0fNO+B-F@;/#gE0-OS_0NFLRI=,:1#b
B?a/,,c#B,.F2.E\XE@a#\&e:2A+NB4eB5fS01?3IbJH/(@E9[;;AV0/bGOKEa4g
\V#FT\Bf0ec^^XVccE-^5PFVP^dNJ8Le143@R_YT0b8gSd_UgTfCA)I9DBSZ_UPN
02;0?PQ_7<IMEI1Tb(N,-HD<ed0T(IN[Cac9Z7I(a;HM351bYD69A3M.H49128bR
+Z[L\6,U+P<3fNUO-^^A:>3b0:a>-Ue_dVSVgg<YLZ24ZFdC37c>,89_(/]OR;,W
ED]86_M@)aO=?+e5G[PXgf@cgJI.;8FF;6_//TO&V?D..K2/cWe(2)_G=>Q#VfUa
+YXBAO2DTVD:DIF/38#/]QP<5\6;2<8,HgJ)_Ufgc-Z2UB;gO4IG3-742QU+RXJO
(dfG0D5C>;-VYP\,/5A3Y8CIN8+a2F/8dIZ4F;bP\Wf]@[NaEWJ+N2RGfbTT]@e7
5DIPS=7B9_L5C..Q2:;)TbYfE3eGf9?c9QNVBS1WfDR6[c^1GH9K50AE2fAR.SZD
U@P<8]Da1\a0ITJMMC9_/Hf\^KUOg3WSNCK5:2I80d2&SGAb.N6?&==]bVS\_XMb
\4@gGFQN&H&T(+GD5HL5;K38_TE8T4]Ec3I,?_?\9fBC,Fc4\EDK6^7TN-J/Tc?:
6T0[=T5><MN\MD?<R@<9Q)^VT<QA1JVM7K]U0LV/SK<[T5G^=LR4[c\IETCFH#MF
3PNH<W[8cYDL^JFE/;52S#1\CDc=f,E[^:R-V>?D.DMc=WB8Qg[JI#Q>&?O,/.a5
J#^NK3Q2\AS.C+IUTI&b^d=2[Wb^D>.UDW7T>#Ff/Z<C4(#gO=&#Ta0^LY^MIeN+
+CM_.#Z9EG@>-66;,=Fb;G+ASAZR124c2U;60[.7PaUfT/AC+:NGH&[JE.d7,1P=
K7D:EP_ZT;FV;HYPNB(f^>+af#,5[cVVS_AgAI+9=?07R>eXVS1C9#J7?Z<J1D.>
W>+5\M\@CPAJI((Ab;1=;8/V-9X/CHf-2CD>4^W=#aDX9MC>af:^)aJ+G1#,^P0W
A6Ve:5V@C-,gg8aaM:Z[D#L2@;+D?cWAU+5BaB#eKT#f_TVS76N/0bSODI0g7LM4
4e[<6_>4.VMP@K-f17Rf8a4I;YSTKY)HLPZ-fTC\T#0GBRV=D\B<9Y4BZ;e/=N2#
3J8S,)]S,RQ^aPS25gQf^<Y9];MR;f[F9W38-FPXbQE_9-:SFdV2d+f3V?2#9gAG
aBH)DK]f?eB9aDFQcD&BW9I1P?,@AD2\,b_1gI_Za(O.fGHMZ&KXWKX@-Vdd[862
8WGWbA-J#0RU_.@eaf_P]19MB+9X,gSE,Oe7@]cQ6XId]:1;)+0EGWYISEcVV_P=
/GVc8S&<)^:[&LY@M6V\KW7GCcc??:e^<_UPGHb^P]5_@K678AA0UTO:5KX7f-(3
6UIC/2P\LRMeT<7MOWV[B<&:c<L+F&#cg8<[YL:<S&Y1FBFe#_Kf<^OA9QIVKe1<
:MEGXKaHdcVF_e4ACB20XW5V-V-1CHU0S9gN?:\Z7T1,W(@LE-EeSC\D[eZDfKE8
_Iag?=V.0>JZNKWM18BA.\MRZ(,e3ScS#\ZX/B>3eIWd@Sb&g7J@/+Ib5EdLaZ<>
-0g9(d:GLOcaP=egB4d@(92PBNc\:L57T8TWRf<()BW-0e\DMI.U8/=W4]2^8Na8
f;W@T;DO(]e@5F?MR51/N[/]U:EdZ?PV6+1DK?:WgfX7VTIISF0J/EIK;2(#Nfc=
+P85N.)0[Y^AXG(^GCL923Y0Mf.X-P+A2ZX])CU;RaXBdQe=]WG/UE^.WA0M4<MJ
a/(4SVMT7ZS@a1.W+FJ[4eIFf)@]b:E:b@6eWTH=geCDX/f3X@g^23SHK<9]XgKF
[&=P/[44I\b]:R6174@+=#)Wge6-=baI0NYE,a0e7MJPQ9GFKU(I&G4P8DfTY+Le
4JYNWD:@Sa))0[0\K@=_BXQFA,:0Tb2Q_QQCXb;4?8XKY^1IM6acLQQ6V[FQ.A_K
S>-XQ7BM;BO></2#_53:MD]&gNe&^b(8&WB/bW5K5cYN#ADf9N2W.Y5Y.>T5/YI]
8<>>8^b0<Y7EP.cc@5K_/D@OPFd5^9P]9#HWg+MTf(d<GPg@].R?JK6bQ9=2I56.
12]GIXQIC?eRPN-8\#5Dc:4c(EA@^]fYBf@)784O4]g#(RKRXD)7FH=WM_U7AV4<
H;0HfNG,]_^=)^VSU^^LK_]7/&J93[?U5>;5&6KbZ]fU])N(Tc0[+bG2dM,Je>2C
LZ>#+^cgWe)2COK3d-WZ5g&#5KZ8H6JR@aBL:PUa/L5.53R^-=RJ1T2TLGc]YY1g
D=IccKEa.<A8d\dBdC87[F5DQJ/2BN49]+?M5=EeQB\gV_b\JBM8;72<=NXVf/a4
_RNKb>S^g+4+.>DK;AH55AG4Y][1a:H,L(X>a4HZ:4A8d7.J0KJ@dF+GV.M;<=+)
_(#^<g)#ILZ\cJfa4?S[9R1+IR9F\A77M&OUSG)OHM[.X:W2O3=A>0]6&+CRQa[F
5>GCd;JRMb(1GETcN0dV/K58S&E6A,W.(VHS4+<EJDDM:1][BLU2g634/<U9MdF3
:N(XbTYLa5X0M2D8WZ1,fZU3D#FI..K5ZC.8O>.^9B8Ld-K6\DVMFNGOUYKeYb?G
H+H[YP1a46XH6:FTgRM((RDGgF0?I?d<X>98U&:&9GBUb?B338[H1Gb]B>/7YKSN
(SR;d.;e>?d6/8702+C_TLg_d/,K^S+=@X2.^4O:SDLJ,D)?NVcJEER^TL)I+DS/
2T1Z1UA3GceY#f957TagHUQ[aN]MAF<UM6.S)EK[Z-9+JK)]ZJJWTN8ZF&A6Qe5>
SIDf)73Na+8CT,Z2]1^<20M(VI9PE/QNJ;0JP&42H>gSEJ<B)9&Z1cQe]<gNIJAX
D?;1K;A.N,CS\6<AP^C^R5VTT:^,8?Yb2:+7N06B9G(_1<.2fQ)Y5-S+BL?5=f+K
W\<A73OA2I3dc-=]Q+5D@VbWDZde4<9+914\V^E&LedTBA[9HDRZ+/VE3_6=[Q_3
8[?APEgbbD0P?Z>,\--gBFS#F1-F0L12XF6]&eeF,O,<MgHO/1LL@+?F3(9cg63&
./E?L@HU5SGUKYM3\TFE2A<U8^;Sc2b2+d+B-gC_ZE_=cZdM[A[\,;Hb7?e+L.;G
bT?Rg&?6?&V;/_R6Yd9d8Hg^aX?NR(2<U?8]2(1[Vfg&?+61)W47WG5/UU/]cP?#
7dbC@[@1&RfX^2AUe]=fgg/>U=5=864>.&S2B8dD)2)K01ZV)bg=]^H#C#/CT];9
37)=aA#@_I^?K7gQ;aU71I/8.KRQ^).0&F)I7@09b2O<GKa>O+H_g#/[QDF:^eM8
_PBPVP\DUbe-=eaMS>(LNOOIbOE0I:b=\?TAUc@3YBJXO1GdD0,;4e2&6(IQS^0T
A[=C2UWO+.bXaTELQ)#B+CdOe)6)KZ;^;Mf>&><g,^f+:K@@+85:/bHc/+g1+;?e
]>/O0A<UQcQ&W-VQgC^<S_N,<P<[13,KZ(934VA1<5gIAL>:Q.P+HJ)TT,3EUV<,
DGRMLB@XC1cUIE312[9f]7gAZ8Z)e1b0M&>dYg+1+VX@J&TWPTD#VV[d.52W&bd9
TG\>a)CQE?&eL,G<9MJE,6dK(abL12<L?=D7b](f&(\Z\@L3>)g\O)RIA:VOME-Z
>Ygd:X^b6#H+45IVU_@A0GQN9QDO5@2>XIRQXWD6HcVW6b?6:0NUBSGC5gO/MFQD
>P_HF5>-/]6=FfN+;(K:2^0AR2H8.LGREK;HV\UV5aT79^)FD,:7_e<J(7gb<Q&G
:K_Y2^aB7KPbSLENXGYc@8B_GGNID@C]H<OC#1YZc^60gZ)5>[da>&D1GMNf+c-C
02+)PN=OOP>3\S&]Id7,]^,A-1E#fS3&,eXe^,A7a]6ESXAOIX@c,VbT2>KVB-D0
1/aaJ^4AaU0(T?X().K#Ka()YXLO8E[[S@^W83P,X<c[59A@]P4E_UEMg++(P&5U
5d.BZ=[9Gb\,RVND]2^YAN>db)P6WK3V/WYO6E:P^UaM)[#deM5\4dOa8NUSePIZ
),6S23SUBV5_;a]OV=]:;]?=dF^-YCQU_@/,OU,0>GJUD@D4D[e5&6[bOAXO<<IU
F,E@&dL?SL\X+/>058b9](Q5d#QI+)=e@TPYZ<T2NWb1<K+:cUJCKKI(f\^Z6M-;
843E16gXaQ\_\a\c,5dZRJS.\3JfZXK>;3\_a,N^ZS&Bf/E.c1OMJ&eR,ZFS#HRN
<9eP:.LO?AW&V+WCd2DQX9HWA./Y2?H.SV<SA8GTDTX8_FA_Ef5.0\+1;H1\.G/_
HK688W.g/+_,T0DVY[#(EMCcTD3<cF_(LPf[8g;;J]W;d/6@<^G.7D]cd4_;N0@\
f7<72#V#4@IK0OL\WR,R_#D:83a9]](d;Q39:EJ)c:NANA?:GKYP0_^bD<GCRg4V
UL0f>:8@QSe<XI.[MdM,fH(4-D-L)\\8ORWE)#/:I&G5]S03>JA]Hc;NO1(Pb@=X
O;aEeM2b8SaG,WOa#OIHWQ\0DCf,.BLAB&NC\LLNVdNW#CL;4_G5L^e3?K+H7C?B
]BRgARdD<\SKPP@a8\]6aES1UTX3W@B-OIHd\P07T959Zd6,]0c1E04+dfc-_PKQ
SV1\U_08F;LQQ9M(O+,ZKGW#)_GfH92UXYDBQ?K4MfEa&eO#AQU8d@QFM>^RgbCR
g^=&Fce,Y>C3+K;&8PgA,^G57c,=d@UL]dJC37c_4J2@]D\U<0Z^ebT;M\,[AWI(
&VcI,eB\M(XJ+OOYeI?c<7V05MJ.XS[4H=.8&KP>XTFC?9S&<>4K/:YUJ8>E,+61
YN@O6AAFVQ^XW:Zf_8V5P67[+/B:Y)&8UB7(bf:A<=3Y8S?8GYH7f@(B/Y6@(IIU
MKUUf3O5,F;8NK@GCF5SIRSA;<U3dIcD.,=7618YLQP(KGDH>OG,093W,+a6DI87
G^1=YPBFgE9+Se\:+VQ+580H(]I)@_Y>@BEH_DOEH9N/7Of6W8.-^gW<SR>SV\IN
\YY8;]PL>#.fcgAI^49OcCF1<M/K5Z:+(^)46UD]72T<O+cBJX6D^X/@,QK?6L^V
a@L>(S,K>Rc@FA,GIAL[7O7D=MP6)VY4-+W(7Z9;cVSADRG6)DS8O]#<58baL^M>
+#=0RJ,f.5YA,\LY>[eQ2?E,O^P1#DI91F.GadZ7NRKK^a[0.Q=U<NQb[<1cgQ>W
,W-OROA6e]a\e6b]0_d-e):dO]_[A?eUZ[+YEbI#38(1VMUZCZ?5+UAb<(f<fASF
^2T(<H)0+GJSK;ZeZ4-,Q#e1.CC+J8YET(E[Q.I+[>2_0PT]VcGC1^M4.5&=#c32
NaeHWPV9g7V;]QZNF:J=FLKY(Z76;?/&^CTQ.5Y&,WWOG(EEcAb]:>f>92K8[e<2
VQ+\:F-IVdN,6H0KdY9MDW2_&6]H^g9Ve_JG#Q^7[9O\d1Gff=U;#d\a)D9RIbXM
6EQ<VMHVb7bRBZD@;K<50H=3Jf4LXe/&P,:6dKaB,Jd;5C6G+0d>g7SMU8E[&>eL
6:&,91[TF<+;-[#K@>X6bTZ]a)Z3],+bC8.3U+.0-6f0S=E[\Ob9cfE&?W6S63O2
5HI9^.[3QNDe>1c)\GE4OM#6>MQ>7KQ8=,6;FYO2+/ZF.:9WIC]c^(c7B(dHI3+G
UDaUT(OaX?QAGEZ.TXTGD\8(MV/?aXL+314+W9USZIJ)M(6D:FW6Y+_1_@C;T0Bd
JO-Q,OX#.9E;&1)WdQ[[]S1c3FSTP3TZI)&YZW<.3f9Hg83OYgSX&?C6G.LaK-S=
UGY^?:5L#SJ]G]Y>1BB:;N<?Y58LbQ,>FZb9R@T>eUCQF,K/CfX3CIF_.8Hc/BV[
VLa,8XH7\&SH.]D=WF7RR1?G-YdPSG1HKCYa/T9F7(^=XV]PP<3aVa\)QGdWPZ2X
M/-O8L/[bWA27C0X)cBHCfUTDPccAXW,VME3:)DN-77-Meb,1g@B/J&TL=^=.6\_
\H,Q-I-bc57G&E2\3VP_5#0>\<GA)HKZ53&QJeHTNa_T157W#[(5+bH5b@I.A56;
gLFV,b\FL(+g7UCX^OJ8/ULggPZ[@32])B&U.HX?T&B=>.1f;c8WLF=)F2GX]>:K
V/g@_gZBSNT#VL+H&f[DaeS3:J0VK.Pg&O]FB4)]@VQZ\WVV/X,=JUQ>7I\)_E.N
cK>KJVaA;5A\Vf.O@H-XV69R9STZaN0T78I-[:#SM&8f:H<eJA78IY;0VI+QCE=_
RfRONW\@>7YM[2LLG[ULNTLV^P3/>C<bf5.LB95^AL/6Q9B>G=8-Xa<BK[D7fb]X
eD5FBW;ZHD1(I<7J<+<IKVH(=8JgN5;00)Q]1GH9fZd8VIKGN_J/IWIfW9GFDJ^f
1Pa=UZ0AF(;G76+H41g^8V7U^06e,8TR>K2@?C>.YN22],FZJZSA)e^Q.82)P+8W
V.B>9K0CGO,;Q/A#A4#N&g,==J4Cb7H&:Y;)UDe)#I,[bA1gcXO/e?,B1H5S>&bQ
QcVQgCGKBDZT]IFDGC>7-=Dc#23d9PCeDbbMK7b(ZQa4U6MAQaATEGUJgM_a_W<^
CN1XDG)N/OS7F&5P(bRO@gLWGB7:D&HBAZXWQ;S5VB+<^bUJL\&2JFZ\Q.0C.d?F
9)-UMHO14IR[D<T/OZBT#d3(W/T>C-&+=4g\EL8QYW:cR/K^]Xg:ZZeZV57fSVPO
[5?UT\S_#Q3,c8b-9?_QcF&&(J#<:VfaK0M8Z+bS2X(9bITeUULbL3XP&(+0f_O+
BD:EL-[[]ff>>672<PTPPEf^Be2Q4X>GD-<ZG_D9#+/4Da:]:BfP,R6AN[EP;0P5
dJ@YY6&>&47A@5?g#/J7N_]]:7)d?QaJL^.-\C76;09,R-0O6=HeK/M(9Re-L?_6
-/_C#D_RdRPQFWS=I9IH[6W+XA0UUG2Z3+Z=<&AKPW8QA#0AJOg@Z;=3a=,I(Ge>
PT28H@SUQJM(_41<?5,3(DASbC(5ZZL<TL-V?P]G6_31S^KNO_U.SGY)^ETA8^^V
f0e+\)K4CW1;&MZEU_=PS<^68(:Nb-95K4H^A[6+V911&7R-ZR6;9CLXW>&_BRSE
L,JH+2^M-3LL,GC+#+@_GfbPfWWX,T/>c9W1?gYgF=#7(T45b-G>0<VQ.>gY)WDB
eSBWbcNO#OGNBAGG@)@UXgD[O^^AY/6V5(1M+XA>][TI#+U=>PbED;e[1T)WV_4C
#Ha4904B9G53,0IZN/,,D0BN2Q+?-O;.QeG26fgIe<JPKgbH5HPd\f/?UfP-8cY[
a=41/?RIf2WfG9cI(a,O<#36/\?BSYc\P.(eRgRVN(H]6bJL[=-/X,-QU;WLW,S]
&P,QR>71D#0,O(.C8c)SeYGOP=5:R4+7:N-b?=:cAc[>&4Q^e/-4FS.7^<Y@3-BJ
2fY8H9_A.8[cOYcESO4cbFddEVSc_<+gJ<PZCM]a1c=G_8W(6(E?9-1bG963OGK@
b1D_HA3c[e\+?Md79_9b.Y85\O;MB-e.Cf#]EYRSR077eM>1a_WFRUH;DZ7HMQ63
NZ)@U=bcE2fN5J^8#EZ#[AJ\Z1E?_g&M9VI[,#6;7LJ\DLcU0bRQ^LSVOEfSQA=,
_)Ne\:5PHCf1:;D5CJO93Mb3g=<)FYZbI(FY(QI\U;XcPRII^T);79/;UegG#GAM
gE>Ef]Q&M1_Zf](J3+Ug5Bg7@Hg<+1H>],H6V]Xa[F)Tgd>WJK)MF]d-1N?a]O^c
0XCMDfF4J>^PfJ30+\Ca)?)5USg3O(&O:GU4+R@29&T-8VK5[]F=_\2?ZDESCY,>
1Ib>0f(K5ZL8cOb578DP1[RUe&W9X#MB^Ce(<#fS\LW<OXEMR4<86+BC,,(GFU/.
(Z+\eR2<].FG)\:L#b080^HME/62-U+]9+Ka&3fDXg=gFPW;NV^.\_<a8H-G4-ZX
9\b:SV2H7d,@JbU92OT?OXT7V?<^4X1S8Ea:UBBDFgQ]\NQ_gOIK-IK),VCBBA=K
^GeB##\=8=)g[9:,4G9N8O#R)aU&g35K-EP[<2d#KV&7,S&&Ue^_<@^GG)Q.JA3M
#A78gaVeI4QS388D\\JaLPAPW:NID+KcO-;0>:ENAHT\?Z04_ZffVN]>?1J>-:/A
e;6[d)OI>7eV=aZWCOc^>IBYS^X8A=_R+c[TD))L5FUV]VW5E<W51HU[f>cPABEG
W=UI+JRFL#H22\O<WL(c,YP(3JJdg-:ROB^T58PBLR3X=>W2]:G@XW<eTY-RTS9\
e&/>O7=4=O)<L_W=W0>Ief6)C,R/YM2RbAO4H,3NMfU#@C=WVJ=9d8D+^JE)3ACO
FR>aLS7C)PKV(Z2B=?7JK42E96FUHK7^fE@:<&Lc36U&57aG0EMPS<V:HWSFP+<<
?LZOY2a:NO+C^4N5OKYC=:Lc^=23&K;NZ?[NIR<=Z0,[-AFV+VELHPJ:B>XNCYLR
ACK(LTP[Y:,M9VQ\@:<[.PO#3?X#;HP(N(3[I=(AfW=TQV@[O9,0cabGKE\F0R/Z
;?D=M]]b]-g)?6COO:c6,Y-YZ=N:d&PB=9dSF[^1c[Y2L+Z9e:JeF\Y&J4SW.L2/
BN-YVCV#\_ID1Y1H-K1FXRV8bLP2U+^N,K5^.+.1<XXS33K)T_=X3,XS5A6KW2,G
4KSYRf;Dc8R,bTW\C;]T.K_B>01ZH78SE+&\Y2RV^S]FBNS&5P:c->@c56]&0-OB
R/]=X97b4d?;LeQ3/PCNDQ]_Rd/+W4R]#J(C4[7B=]AU]IPU-3=IZI0[fURA_ZN#
UQMH[-7.D::?NI?]V@4E04]7A<EU#E&;Pd(UJC)0)77<K2FIgJD7(1)D??5dB[9]
Qe.dD2HTQeF/ERCISKLI&f#LZ^3#E23,(MQd,TJ>_.DIBe3/^8#e5P[R?9Mc/T(?
GEeH+G/ebJ[(SSDc@=DZY<Nf_.c+3RD7&YQ[95Ab<^NEG(Z>-P:_,-5U-/K],.9c
<-eGBS2<0RQVUTW96:?L4?0L2AX969@H36d\.cW3Mc8feB84?:59\;4cg8EcUKa^
f\>DM??D&VJABbbZFW?I[d<(adOLcMEK&M,UG.?a][c=V^,<58R[(LJE[8aCCN&?
MPH5)fT06SW8.[=CB;0A;+YE_M#:=TF(#@Q&?c4a\f8.>A^)[,JGJ8;V#5;8W@9K
FJH:7^8\Dg_\9ACPAZKa:678^C]EHJV-KJILKPLg)-KJf2Y&gNXBYP#eUPN;9F5C
1K4^[H:[U1,[\f6),8YSECKdWM_C/7D6V@bQYQ:eY6V[2&]d+=2&K@AQ]IZ2^0WG
eZ3,/gJT;94)M&TE-e\15D[\)XVdUR7HB+@5B&P268H_TFBX7]b)WfEUDLS^KKb(
R1#3)WM4b0OV@[0\c\7Y?S4B66d+SeF[=Cb8>ca,WU=1[5V<(?P+\GYKfPLCL.N1
K56K<M8+CIGBZB05SQedCRDMcZ0:VZ=b/FO6QA(<U4H8DXe57gH.QTJ49WRA):BR
_ECc2=?F:FV>FeA;AQ.7PZE2GZ2bMKa-P2_?K#ZYB&#eG_cVLTBdg&CA8>bD:G]g
+.=/W683==>e\=fVR^+CPO#??Q1c/<@c-X^8SR5b\6:@/WE]4KcCFJW,9\W1gUQ(
P=Q]cR90Y3IHCeT,&[/7RB[8bF?3\XF7>]eLJ?@G8Y87EAa-F/=(e@/:LdW\41_?
V_.4PV32^ET-<W@>?EHM)9,J2/FE,BW^bW9>P2-#:6_b&R6F3V_F]XYT6.gZg>RG
0HEOH#WaCGX-7Dg\FP,)d8>;abTfOA_2MJTA3SQe?LV<QCAA_NcfOO^L3_1WD)-1
C::\KWgZ:Pf[@ARegKB>0]^bgSe_1:#.9)-?6;NY;A-F0XOJ,/KJE[Oc[YT1gHAR
5(R+^f5(A^>LA(?Ec<0ZU:V3agQD-T.)F4C=a@1)E5MI?1-R#PD9<;<9.6=Z>@bX
,R^A,-8JT&74BJ\TLBXLQ]g5aVB\c(@FPdM9-0gYGf,TJ1X\WL8-0,=g]E6]V0[W
ZCX->A_DXg<L9XEK^WA54?DXIGY:CUYAN>ASQG<WQ39QRe?9)]IRc/],\Ja#:01F
G,J\[-04K8:3fWB<9=@#6:6Q5;[^O81Ua+a6;)E\@4(II1EZ0a-@#.FZSe8-<2:3
R\B,gA57R^DEL&_+HEU84cLZ>Lf[]JKH#@U(G@g_@QI;f<KL1:gWBR>&5=7>B+?b
Pcc>Ce&Ga9<?.?D-.0G9)G,N6ATc90_V4LUKC46C)JKY?BU2LL]V[2Y4NJKQ1=K=
4RTD78OfTZ/[[7\H6LQf[/K_CP,UYcQYC:/ZXK:ZRJH<7LaP&>HTGM]B:)._X,R(
E[_Z6=):=4UT92&N#P\C=<YD>5IbVG;U^W^f<T??AOADV9-D^(^YY7BEafNSC)^S
I@K]F&PM5R<G\W5[a.(d<6LR@4>JbfcI(^5[JD)QG2HDDV(ST+OG^b,e2c?_CVW[
]72S#5A\aWUX=2[;URfGIGMVPKBVFOV7EB:<S1/X\JV.>Y7>&+DG/;#RUV-LF&?f
R)=E1L]gS<0O1#B.XBaGHZ,CH5aF1C;[[fILM^aC9UUO@agKBSH<a5O,Z.JH0U5O
g5d02FS.2EY.\/M5G.DY#@abPFUN+.HD,I-g;21<IEWVKP5O@7bEUYMP9a6SdT5#
\S0Oc@R,GXf_W.Q&ZA+9MaIPR;2@@eAYBO?Ab<#&:ZJCIeN_JJ4CN\Sdc+VabXC8
F.\&+T5E,R0:AO3)UOTTXg03b)(PB[L5IFMA2fU+134.V?^/bQLW?#I=?d[TEYFK
@&K,bdUZ,QSPId#9/=A\GSf.\+A/g\UeJ&JZFD,+#@S\T=@_;^(eTgD^@a;1c2EQ
Yab/6CA=A8eC)HSR<:O=95OI8[(&8UYN4+1SG3:UK^8gNb4DMcDCTMA5JI3fKT3]
,F?1I<+(QBS1O710.97G[_VT,6[2S8F>bUd#:ZTFOOe^9N7YPY&.-L<[Nb#?RV/d
?1?#;P;H;01CR=86P5>3EY7?\D?NaK8T8>9IeV2)ZW]W>[BW_-JPdgP?RB&9MY]T
_dODD+FU:\7W8<4N5SP?.3)I;\8QL9TP?&?6:+//_2AME&X>PKDLQXSIQIF&?VQ(
^XQ<B&g3TgM\-]V=Z_GJS(\+&PF(fQ1IV4<.AJ02cJS4gY.0dCH3;),c9,BCb:<b
c1SAS?PYNG895OQJ:KAVDg<:5Y+/89d<U&PNXM0H6P+GcRMKIW8-Q9cN?eE\DQe_
b?]\Cd)=M1]f?XY/ef,HX5:JW.FR-c:;C5-DC#GYT,;,2#](,P(QEU,,_P0?#J-2
E)FO2UNWR4E@A#?6JEa\Rf1BA=>WOU#27?IL.5?=H6daG.UZ(37M13(3O;K,?-g_
>O<;&(H^,;+T3X2<:;cRLeRb1F^BJ5WgA>1HUbZOgaFXN+9QdBSe)1bdXd&fIc0/
C[C4,53#MJH@9\:R:Z[gSR3A4f6;&T6:&3M.g<Vdb.+4/R^YD=D/d]AC_7HSO([S
g/6KIVX(V+)416V85UL4OBP1dFcT1Q5dC.KgJ?c)QJ@\R[D^Q0g01b+1NV/R>3N,
C92bK^OgdgJS7/>39P,J+(D//]b1\5Ze/ITS2CWJB&&P1W@]EH)S>8f.R\+9<NaH
\BM0I;X1Z#+#^7fNJ_YB-=2Ac</7Ma1=P]Y5AUI77Q6BL<4H4;#=>,)bEP63.VWQ
caH+O\ZFJfA8^>OUe4cWBGPNL_4#dUfgU)0#fSG2HgaRgQc>AJ\;C1=bJ?c>1]5T
?12f<N6(C.A?JKaZ;(eY5LW4OB+DFB-Oa,PU@QI1BFW3+I2A)8S#X;J^T=@M#2W9
F>(\B^H,Q#bdbYGL&^,FO,7XF1Hf&eIKO9VR?1&a^@X=1T.[JFEaR\LKEa\F^cd-
K=DfMQ73QPN&cJ]&dd@ab:[g9.76YcELM2C\\.JIWXG])gZdN[RI0(6>A0-_N2_N
#+WQ/R]eEGgL0CF\e\R+?P:XF8H;a3P;bBVd#)-:.F.T6MDXJ=\HREF,K=^<@BPA
G;#Ba0#57O+TE/UULbMHU2]_NN\,@/KNJS#T1#a]#5A@4-.ULXEHU5-?HX[Tg&f/
_d@a_P].E=()P&-VS;bM,eJFE@f+2U8A@,eX_>HLHU_1D[M7^C&JQ9FV]W(4IaE4
g;O>[1N<V<Q-QTWP=/#K=J@?UUN^TA<f=6N8[=35ON=?aM4W@a]5IPeNT^[U)4T(
-8FV4,P_AIE_fLO^WV6&_JE69>Q2Z+RM).4U[1)Z=S^ZFd&3d3Cb+b)2Y@2Fbd5_
g8P;W?gL>I9fNUeeCcR2M9WXV<HNWZAK@^2)g;G-CE\WGG#V]eE90cDa]8[#[M-5
?9WM)K2GN=GP;1D82ZUbGeO6+f19.=HKd3#J5CPL,[Z6d&I2DGaYKB]eg^3M(?FT
KU<1X(J:^Sef3\+e[[6e8[;H0^#BK>O[],J5EM:=UUWa8W;a)D7J9=]PAgfc&IF_
&dQLdU-NR,>=c@AM^[(@,]PbN]+VAQ_)c+3P0D<G1;X/2L1-+=J64O73L=A8MA<H
?=QOaDY9<XG0F7>f1@>a=)ZQ2dH6O<<O^VYgC5IA)ZJPW<KZSGB(O?53bGG&ONRc
2N_1GZ2&FcPLY6&7&C,V8d#HLcNR#\1[PA8=))7f3S2)g/NH]5S2#.CJ5J4&ce3&
6G>_ZHRB,GeFR2[:8Q&bT]b3_0Y]7YNA#6-+N:IDf;AQfbHKSR^R_FZ9Y>/(U_)E
=BUH?^)CC#67GeB(JW)\L.Bg_PBf=JZYF@;F)D3G:RH1<3U+)Ca@+0c,R[K/;A)d
C:8fP@[WP9YP#?O0T^XgJ.U06<GJEK)N]GfEQ(Y+[F#H&H&5XIY6D,)O#,2DMC#8
:\Z;VfP,=-WcEXD5gHOLE>WMG-VG[-1cXfJ5Ag4(-^)Oa:-G+=S091W=KP2<:;?S
J\f+VX3EY[U;>gW9cEHJ4)W65.cd\:W=-e1/6UX_e0Ob^LSFW<)F<_e#@H_cCa63
(GQ]H:KNA#\)7-2TIgIV9?B-)bK5?daIRdVHa-K7b^G3I(^C:OgSbC=55J,5D=UP
_g+8e.W0;a_b14]?fPdK^0H\bHKNEC/GMCZfNL??UK.^:0C9A\&5,ac+)/&?G3I>
5E0f#PRa0E2d5IU+C0#2WbUHF\CV.;T477?BKOO3d_7e+^:]e[<@b2U2?)X#aBPC
?3PAX&Y<4</#gd\Ed>EW:+S?QQ8A319SMU\0g1)\8<W5MM38]7Je\YEE)5\K,WU5
&2240FD=,9:#H70ZTZb]Q<e+@SF]R._HbS0^2bd_bUJYT)JHG;))-3A7^O1Fd8DY
JY6)6HFf;;.4eeD-/QZ+d_GX3M.WTTYg+UA[SQ>&]?D=,Ng_,SW9DgF>+L.0GV9.
OB<]0I>9H+C;?B&L,dd+c_cUL=;]D7I^ICWH8ZZ@SAQB@?f75dcTMdeQ3^KCNR1X
VWI>1>;c;+6D?>GNBI@/,6J@YOJ9G[RGgY:A97YXK(+RKHS8#LNN7.Q-1+dT1SHI
)&MKB]3/a9&Z[5JNdEO1/bHN&(,2UJT+KeZ2(+gfDXNff,(c:QLD]aa-1(2(4P?&
Q^RG5,#\N,Z.5\7TR+OHA.[WbfLVSCE<P.;;e[1,DAL\f3QEL0L8NOMI?+A8VJ:>
O>eQL4M_X((Le2A,(S58T]0C@\2Q?1FT(XVRB.G-,GfJ0-YR;d(^47KX,&B-)[\?
CZ\>e-HD2f-](?6=1.SOX;GYPFIR]<^TFSI@5]7S9D.19K>D)DICS7)[H-5g>;9D
D/)RS=]95WTS=f8;[YETa7-,]-SG4.1^;,0gR[bD/A2:&V/-f_N?1;ZD&5ULQ7)\
TZ3B:]5UQBCJW6;:,U.[00PQ.)2YJ.>HSD1#NS9FU=>.9\+cN&Y(#7?)=A5Rdgg-
<8V1A]_f-9Z;6GXb2MD&>L-PLP=1PGfX@S/QgTX2\.S1d#IT@82,?[;<;K:H4e)2
@BNg_Z=Da6fLU_d8dN9Qg#A_KY/UN=;g.V5^5f3dPP.\>2I8D:J#P\]^<]+N-G-2
>N\YJPB<MG#[=1b9HVRRR_>bK#\YUefH<RWLMLXN&=?8[],199+O;[MU_;XLVIHf
WYAMG2)cJZ5J)Tc]52<AV]W:HLJL0;;M#W\-XH&I=c9+K5c09ZZc(d3L]CR+E)f)
OZ;.K&DE-:N<b8W[eRIL--G-LNLNM.P)gE:b=\V[LYJ_:VdO/W_a<@d)Qc0O7M,B
\X0?>J=K]fRS63HdE9I_U2cS29XZZT_\<G2<3/HRZ>PTW\8,3I#<eE]\#10b<(2K
S.E.SQU\PPJ(dNZKfb[3WBVdP8C3OVU1W9c729DcZ[\;c&:9.-C4X1SR[)VO)C:c
KD0d3SgT8RUN<&1&>GK+=<U0,>VH2;L^UIAHWWU2f7FD&#B[\Wa-TS1ae</X/V#]
TZY,+K--B(34R?gFc>RIB]3(9<@H<G#C_#J_R2P#/IIALFT#U2AHHa672#(g_6&)
N/?)dX@TI?[&C,(VR/fa9I(9H>2SU:&d>_#=+A-(#=U#O^=Z_UVI>/+5b\fN.@DA
AI@/05F1KM6/E6;&c735b9,\E278L,RB;VM[I/4XDZ_7>)PH91=FVDW7ZZP7/RS+
<T?4_/G^)8f1c:Fa/JPg\e4E]6N<G/<<2]5==(6>gce8G(5JW:]LQ;gdD/]XDY2Y
0SaWV=gde0d_b:O[EJHP4J]c-@?#-e&0Z4VPZIOc@D[fca&\+O=918(J<:#La@4Y
M^LMB(F+61O[YNJLYZNK#/Q6a5daP4UM?Z(.=-9,ZJe\CUgA&@6R[;fM1gL<S#23
eEWDHO\5/N9@WgG,A,1(OZOAVdUJHfe>CRZQ.=7@cg)T:EQX-e&BabYC;B1:fdE.
CF_L1?d/XSgNFaW8<0Q71W+2&GHI8RMQ&YRFW&_M6QOY[fZV7]=)]g8U&C23?2g^
MT@4;-g[fFOb5SKg4(?>;V)\6(aD;DgTS:E5LTI++@>_EQ_2.Q41]6=\.8IEeWgE
Q<QD2?FdFP2g5;;_]ZEFUH(6OdR9BX&A8B[+;(7R;Je/^aV(;U<N7-CDX:NIXOa<
S)XS2F)e6Y.]#6aLEG?0=[+_\U\dK?^LDL)L+F@F=M\)P6]>(6>Of^\\V;7BVYL5
EI#OLdVO-d8B:[ZBZUIWJ;D?Qde-O9FYLYf2IWWb5GP=ZR+7E=feBQPK@2F:6Q6D
Z;R,D8T)>=g6P9=^T\&=?&g6G2YZdB4B\@]bHbXL]1dK+BG+gATY44gQ?OAE01A8
+NTJZS:@N/1N4-FCAbI<OHBFQN1)#dWCe2Z=I/(K2G/dA[I:2)E365F<CM^E/5X&
L,>SUadc@EM1TGa,bRHf_2P89fDD9J>OF=d)c7GP)I1aV]TLR>b4=EW#aGdKcHT3
5=fYA0QMgOGYfYO8V.0C^1d:eNIGXIB0;GbZ_H<ePRKdKFZX=bJg5>S#9^X?92GP
gbB@P+DH>E;)&bZQ?g/[)0JI4F=M.\c>[2[9Y<XGK&[:A1gW.I14bLNRO[KO1T<^
7)O@#,Tb[aJ3e.O>QT6PLZ]?NHA]J;\8F]1?-PAYcA:48(#YN==C9VWf[b6H9D]1
Y@NKfHSgQ=)ODWWR>O7CC;Kd5#<1)P_cJ&LH,EQV9OO>3cH0CIWHf5=^cXGOf9C3
LPQNUgXZgH3CD/6:&\25CaHT9.3EM/ZNG&W(_3:8[HM:-bB3J8]S:\JFO]2<5,3)
:P@W&Ze.dEPO^U1W7GB_,_,+NWUDOG1GS><aRR7-.HEX0V18[V._^2#F<a<b;BLc
^D1.:CGGFcP)3R[31.JE;DG;\fgJ<,5\B8TL3UO@:2f)^5<1(1H4,:U+J05OJJ[3
,2+@ZE=Z)2NK]&&++N#G=AaK/HV[\7cH4G^N>LaR(;8IRM@B3Ia_CPEab;6^&TT3
&FD:PG\4G[_#>)?NR\;<.Z]e()>:\.\XZH;Q>VBI2\QMOce]gG,1:@HPceE&)<V+
5C@]<5=3FSG);_4YbARRKQFH:VIbKXGH10DI<KGD/2LQGF0OOdRBPH-KO3-0KB=5
K2\LW4#)SZdNeUY@b+@6ZBRVFDC(<;[^4UbZ[8]C&PGEP<[B@E6;dR@a8#9YK-]A
d+(\[f/MU-0#?L8SUaZ/XfN.+BUe+(6+]4)E0:bE#ef609FA1S9:,Ke>1]g^7QA4
E@UIR0K08aC4B)8)8&Z&NgY8YGH3BXPXM.X=>VAVSX\PCL9?WDDdCa6WA0Y57YGc
^AdfKdJ]>dSg2P0DCA&9?3)+G/_3[X#dVRLK7FB,0Fb#=XH)8YBb8_3>2SQ]gRec
_R&.Ud7#6Ea>#^I,&0DJ#HYVf/]aV987.+EYe>_U)87T;EK+,>e>/;CC7#H)3/SK
ZDZ-XO+O)MSN5XS]B3S;E6OI)be_E=ZY+XJScKAT3+7U>9QbbBY-<aNQ2<JQC-^=
6gI2)UW_RV_Oa:E2>@T&Z^VAIO.F1;RVB2&;.d),&F\.4)@f^T[eC.0\_@=+(NHF
95.&KgLe=C55gQT>^gbe:,fe1dd\FRIcGe\Z8GXKPJ^VeQ^TfS^H#<8H;K0MY+71
JQAb.IC9L,1Z7bV?@QLPGVP6>Ed+K4(C>QKC6cIDc)IY_7TPgb?T,3bIN\eBGIH&
OIUg4L/5Rd&be1Q\7^O(8FZ\G4g8&KKL-8,AR/L_@(fR=3)P(R3]^bC+[g.AJG]A
C@bRA>W7c^Wd/;#Xc#VNSKGD6GVW:#INOA]PY:DQD=&BXR;ZE<07\3Y#</68Ge/0
I,TSW^eEcMGU/3.(2#7Ifacb<]D3Yge7W40RgX9eL>IJ>^ETS&QA#(&(eXI/(/TQ
\&]D.YUK-PPT?0<07]-@3YSZ:L1WgIX?ESfLYHf87RX?=.Jc-_SU(=Vg;MR:I;N=
/Q7:AP?\?8W)5AX:70S;WB#NY(F,c@6U]@OU#KPF@b3RLZ6/Y.6E80[dAF2B#+4_
T\Z_T&R^VKZa7)10K<Xb8T,>@4P[3e=UXIJ]M9RMA8^0bL/#,XEeaI33E;FKIK(^
;UN:gb.3E<Z6:bD&(EA3W@gEBVD/HRPYW42?J0P05T5?\@^Y46\B.9H0#_<;?.W,
GI@=J##2UAJ=EcA&)3E[9R>5LABdQFG8./QgXD.76[[/Q]00MW5?7UQ8cP?28IFT
ODFIKcDYOPcHP.2V@M_e2@e.5EB2(AK&E#KET(M9B]?5TPMOMCcQ<a;gQZX(L_.D
(A?UFHG\6I3A[<bL863^+666M>9E_PPW<&M-aU8fNDU&7@BfIW5^QI&([-U#B(+&
8,#DPAG0L5&,3S5#OgBZRR0:@NJV?d7eRM>a/TOG:MJbDEc4.?>f,?QBZ[9<//b#
MN>I,V#5#_2<eX85^EI8=A,[.BT92ac7c,f]Fbg-\)X:0I>C+^6d0SaaKXKd+@?2
R+EQ<Q6KY<EWI6JOT=#P:Qg69;b+C?\@WP8a#XP;R<\U1@8ZF5L3a]8_/K0,,K8f
egNOODZd^?J<IDL<]U1E8JX]FWBYY7OB?8UFLESL-S,[dAbY7]Qb31?BJ[gGS/C+
.2Z]g3UQXCcc0:Ge;?]]M-2H@U4;0GR/XUFaWX:Q6GXCSI^#U1P[I::fGZPV0Nag
VN3gXLNB2,+>NIWGLKQPaKXcdDF;[TZQf6:(/[8KQ0(0-=]4>HF&DIQ7JAdFO:7,
<XaZ?@AXON9[ScW35T<^ZK]Y_02@P1:.-BdL>=VM-=O>KHYK8U__/=gC5@We?N]F
PX@5\OUGA#g8FAe/7M]TSFWJB==8K^BX#BPdB04,B0V.g]=1<X_>4+X>g8_CaJC7
(X_V-Y:>Id@__^dZ8YJ=54[?SP;>MgeCW.6\;c3INYUJO[BX]Mb)<Hb7HL7TfL3H
.JFO=&^<6\[S&UgTa@338^J\&F4Y:40U[\Ma<dUaGPTbC1_9:2?U(CIE\KIQb+;#
f.K<J.dbIb)d9I9F1c.)gDRK\Z>R+bSI^S?)ZDGR2\?TX>d=aaS+Z\Pc>XNYM(<0
N3^1Bag(7I\VP&C(S7,VQ><>&DNIGR@XZV3::/-@aD4R1O-N6L>d,&T<\?T;U(ZK
J^M34-6N)Q7:Id)]0OTBLWNV-1[g:G/6B+SXb(c.a,1Ie\P7+N:9L;Vdf;a537IU
V.9RPY=0+Oc7(=BOUZIfI];^L-aF#2.W_F2M9cgHJ^77&&D3[YD@QZNUAAc\@a0g
@31^0W=5SgX@-<cgC#:\B5bC=88fXP.MTY)+J]fAc&XFT+a_YcZdA,?g#\R(.+@@
^fcdM_S1(GP#Sb:/O9gO0G,LIT^+.^]\(-KRT[aMPX)/M6;6YV_+L_B5MdBHOLUC
8\HZ-9[7LRU(@CeIZIB0X_6=J1?6KUZ>7cdVdX+C#SBN@1G_Tf[aEfU:Y:+2e1A=
#S+R(J+.N/PVZPY@IMHE:3C8J6g+_aQVHf9?0gER@EW^@Z=U.eba_+YD/\+E0Z_U
>&7SA:7,:RfA&&,S5ETg75.\7NN<82Ndgc.MBd6VYdA,LVUON(8A9:LbPXX#ZWHb
5+b]YKO2G/P+[6UNY3I=WB4KL\dJF5KJV)5-R8AO\5+<Ta4E?Q]8gRGEa]E&Oe=J
gBDdF)I38-/NT19JXKg8+Wf&X[II()ZLIYO>Tc->J<M8RD0-ZQV0#]/P9,,2;>IC
?SJbT:e@,TDeXfLQD]KTT#A6B5=->7,X1PU.?-:9Q6X(@6GT4DdHV)8e,eFC7824
a]9\^?3eZ[]=:I]G.O+dKdL2aV9):JH+]Y-8O-8FYOfE\V(]e4[fFA<M&?3,PGS=
Z^4GRU\Ug#PD-g.KZb>TF.31?,ScV+)0#J4=K)[[+0HRK5Y@Ce(c,SNA4=2aMQZ+
dgc_CT#fOJfZCTR>,9)[Z-:QEd@LRMV/YF74e7AAeaW>G<JeDdb=_W;[OT9.#E.8
XBC+3V(]c5eb_&UKXb6>:)&<-Xe[a/=@SFdAa46P-6[#_H/>2,#_G\5G-T<FgFcN
H)):(f)0]Yd+69OVTZ-^S4KPU.0A=()S<=8?C&Dae9E>_Vg@V))Z3XXdg@<a#]KL
7BMC,:+5O3[]M6OE7C5;N)Y&JE?YD:U3),BB?dG@gU>DLG:e8CTS8P\SfZT.d>D)
H2f[,f97b:5LQdd&,e(e:FC<V5D&83TO<f0b-^H[A[=;0Y::W6)(();ca6(^PeI6
#Ug\e:gaX>NBEg9ITN.e5;GFJJF9&=5QAM,#03RC_2HNF2&>>L+AfS?VKC_KSZYO
TEJNZ+^5UH_aP[M(bX>2U<7CYWZW2g-&VVGJGHTX^6AC0&J0U.(Z+-N=W0_#g>KF
-S7./M/KVY9Nc3,CBLaR#,;JYJ<>+&Fc;<^G7>BaNTW]U,ZGGC_c:eB@+b8E5Gc+
ZP-GBP.,D#aBK0Fc\D&=G<\5>3b98_Q^ddOd;.44f0\<A5Z7G1a@B5E/OZP8R^7/
BX42@#6-ZcCTHC)Se\.2(&dPZTX-[Z;0.JCKebOKEK,[)gB^V9&\4O3e#6fFTaC:
V^BZ?EH1A/K5R]^S<@8VUV;\IXf8IN?]IZFa_NHf=&\P,&_7\b2,R#bYVZ,A&I6M
&eY41gJ)E6K]B@KBQ?_DS5]eU=fg8+XgIK55OHaSbS;bN\[D.L&OKOSY@JD5<F14
MKEW=U5aR<DM,Yc]385TeZ&?bH[A<5#R2fXH^M?8LBd0bT.BgIPK/-M^eP_c=&&\
c9P(>YbUQ,PbRb^D8C)eYMY(,]A(R_P3]Ne3CF>H()>-#aeLf((6:0507]MV2LB^
F7aTb?>PV/Y4GQE&SCJgB4aHU65U6G=>c;bHU01+?K7g[Zc,46FB8@,&T0K]G+(:
B^>-QI-WYZM,G;JX7c#W@C)L.Dc;DM#^GdUcdT@CcI6^&BR<190F@=884NG-\6aG
^WFT,_AHD)2H=>fD^&CD+M9d#0\gXb:I(6-W+aMMT5e#E,D;UbMW_DPIKW\07T?V
FI>M&W@TRJ\A?c(_2eK,H4FYbTD#FRT[S1._16EFE^ZAUfRD,CYQ?CbDZ[#>F,Og
>^EH&5Nb,:9aBdWQJ2;JKcNg]G)-O:Z)EYC:)cfcA^;6_/;I^SC9&91GA:e6&U0>
HL-H^R(C?6P7SA?C?R\S==SQ=2I-IE:fI9C[/.ee7]N,G0DR,c(:COZe4.5-f(6,
dQ5c8Mc1_5@J-\8^WfLDC/\cLA6Lg:Nd\9,XbX&A:QfWJ6Q70G_P()57DLL+;-X&
K&B]ZLJ4=.Y?2S:KL0VUJNFN&+;/J072/DOf+6b4GH,4A9NW+M6L=?(deJEbF&K=
1/R<.44Y<WZX-J2GL>ZMZ+.=K\E.U><J6\:WLN]V1A6G7@g]86CG8?O(#b)0M6K[
(:0f3dC\ES9LVL?=0:KKI5dNKP4eX_5^X)K#Y#.d:&[9^S1.ET^B>8&#M0/A@,SS
[_&1C:,2.ETSHR18N1<=U/Hd84IOB]?f9@5)]7]:5U=0E#:\(C:cRQVeVc5)0QN&
[)WKY5F[^+U^ZPC^A-eAN+/>5E1<WPee@,65WgEA0WLeNOW-@WUaL<[\cR_BFF6^
U:HKL?3K4-+,1eP6[1P?G5b+a6:\(&K/9D]AGSY&1.QY^@@P6OCaMX)5-3dR]W[1
.dc-fc9O9Bc^4X3O0&\36L_6QP:BXNXWa0E4AYFO_L>#NeAF-X2Hc<T7@]A;LPV>
3@c]OTWI9JN8US?g_Z&4>EO[,9QR?[LMCIg#HKeF><2Qg/)g<bH]WL#7_.^L/L7]
(0Y6NBD)#f<EY-b607GU=8MZ&6;#INBWDFG0Y/+)6OLC9dU^(G5gM36e+YPXbC1=
ef91BVI9P1J5IS2]O4b1QG231SIV>M=4CfD\FIg:#_cBcd]3J7D]a)(b/^6.(@PX
A8Ne3b3XdGL\.70:M05+OSH@g,L:<gBbS<O_.^=X>@<HZ?RCd+AHDRf6.,DN=<+[
9/Q<bc0LIDC<V>ZN[PcUC:JI,=Z?gCNb\V9;79e1NgVT4dO,-,.J6AcNRO=WINH_
f@H5XI9UQe:DGQ/W^O<@7Q(OGJf0dU4\5HOO.0c?ba(4EWI5A/Dc@M\+3X<(fAD2
/F4-=cQ#@4Q:#<+#(&T7c7M2[(c)=a>gA1_3XKf(?)7d6O+Y=J(a;bf1(57_[D+N
553B<93aDgZJbI_aJPVL?>7OgK=I_4eMUaGa@8;[ad[PdQM))ST_G5+RHSa4H&T1
eP[Ib83<([<9\#R[[Z&AJSHP3?6&/B.EPbXIY;0GXKgU3YA25.=a@?g>)YX4@?A.
;^K+dP4dICKA;b&-g5C/YW]/#T\;IQ@,ZQ]?0ET<70+RXc,WJcK##ZHE#O=bZ-9S
>.16]-RWDM\R7[X^P?#<\8>:T.RH>=G3M8A(7HE63D2J,--;&AB6+C:d=M6@3c^W
\JZ^I-U,2B;KN@_58;&-X[A-5@?E3]),aQ,E5/KUG&WNG]4RCcRXe<=7E+gG5K]]
([F&+6IE<6Xe[KS@).P<Lb1ZA3f@5L9[@DUMR0N(,PM\/E-PS&JQ/gN4K5D.Hf97
5\08H((/7gPR:67c(:@E9D-#?2QNcaIHF-8-1c_cagZ\ZB@Z^^Y1&6QN&I2WET2G
cbHZZ1IYM4]4]:d[M(3<C/FKYg;HP(;(eRab<KTA[[N;TGIBHG<EZRX0=9=L<5P:
1MDdDSTZ&&S25]beVB4[QJDa/QX_IFQ=ZCccbLb0<<Mc98aK6b<((,?bNFf#[C=@
IARWT1ece?GO=gC)fa[KXLCMRBTI_EC(9H-T?7FB_Q,<8f^UTe1eZ,5&GCWSL[(?
?#/1;EU0KW,YQ=#D3GMe_:Q>EMD\V5(>J6U4.=M_Q(,R[=EE[b0TDJ;ENfC141;A
a&c<SC@;4_&P]Z22\#TTRSMFe;HeacD-N2Ee=XT4-PT3_7T_.+SB,O[P73U2-(#6
;W@Z,SJU8e3A6)0)\Z>VUM4I5M?)a/C2(78LWc0I\GD?,fOdR>SC6SR=L^T[acbJ
Y2K_0W4[BaJ>WaI#:aUO0U7]S<+(OT\(L4c\QET&FF/Z9Oef>D]RB]24T5A\7?CV
H:fW,-IcQ\dY-fDf5b5>@MKg.C].[c3C]D^B&Y@UNPD:C0^=1,?@TS82d@&H6B;]
f6dS)R4;XNaWJI=QLJE+8.-[AF98VI>JZ^U^8VR@=Z)PIWfF--A\@?]RRac^A.RB
&PM-VH=JdMXEKQ-N1g+E[-US=;TD72eE[-XT@URV[XD[(cKW49f.U<;2/Y0f=:VR
DL>)QPCOJ?F_2d_He_4@@fNFQgKgIZ\Z7VA85W_Q&[OE.D_=aKb\b0,_;Jd6NG:?
]LN,;>^]0R4GPfN]CV=J:N7AEASVBRH,V[,3DIbP:LWP<T7DCTJJ<K4cTW0OL<#G
-NGCN\YfQWbT,3V[0eGg@KH<YPbRLAD?fG+bK:[9F;_0Z-DgKRSI[&QaW.+b;RH2
N,Z/425Y2_ea32S?,^;]0746=W>V2=Qd_Y11C;2>NZc5\@3T,W5/I;JEgOI0G3W_
+A)D+;<K]YKF>]Ud]?-F&-\\)_/gQ]]O>fG7CYAZ-H8FSFTc\5=dYLd5CI0aNFU@
::/UAR[_?&FHdfTJ;/#FO0#<g_I\T^2LAU/VZG<&VE##/(c7872V(@+C8Z8,Z[=_
(=8:=.S:I;cB^12+5g;:GR#^>f^(Z#dLO-I&?FRBBW5H25LIQ9I]>NdfXf04X\FG
XXMC7)2OgTafcV_Y]DE_VR<=&a-GKOR9D>Y<Ic6W>?W)PH9\NT#7:GQgQ/(GY3.d
ZI.6H4f5SFD?d8L+66)>8-aFTSYbL5a7_]29==0PEeY3CJYa63P5VA2IZ/]NZV-c
=C:?gOYADLM2=5J_W?5;XN5ED\<\&602[/##Ib8cP/Y,.537T>=78ZB9XbF(,Q7,
DJNUX/0LSU+HJ@fYNPAHaX,0OL8](4[[_(=^e:BGH(6@,dDbcA.<aTZdTQE9FK9C
:G-?I#^aJ@4gJ1P#2fK)<-(5H]b&?UG]9GXBHbQ,CU/gGgB:f5(U0Bf3792Y3fP)
WYKJ[>Daf,],U7HUf/(V^R>(D]\1?UR47N1\O(#_UFX#T3U7:7X4gL^R_e[[]c7c
bV?6U&82Q=,D.)GPFE)9)NL\\SS?XRGgC8+[N17A)>=N:dU5KV67Bf<V)14b)g8Y
]QWA_c72,1\#59LRcBe=PXB5-5Nc:B=_07)<OGNVa<;]D][c#=5U0OI7DfXc4(\(
+fZ:QI4WL5\]MV4M_8)A?D;==UU<[9OW\54IGSag,-e5IggY-#TP#3@,dYB/F..=
?Q^>O7c)7@b8ac(NR-P4;UGK/.P#.2e.(]f2V0FDb+<<b5N?,YaCf1cVPM&Y6LZ-
GK,\Nb-39Y/:9#^fHE7#/7R9A60\gg>#U<Q^-RfA=B_\MeB9L5I5JOT774KC1b=?
gHYSQ3N/]GI.(]<Gb/,FTTgU=G94)T25+^3Q6OWaWZOZ=00HDeH6ADKY;H#&]/;G
WQNKW5Kd8M;.?9g\PfF>V321>+V]?#;dVZ^43367e&]c=aG@J1gKPFN@a_Y#;@[-
IDJ^eJVPPfUTRODeMPVbK=S2cQ+T_-05UHZ]5U66##fX[cSaYEKC]WbX^JcfSFP#
2CDY]b?L91F_B\Y]eF]+e[Q57[GEU2LI;DVIFUU?6\1b/D[8RAR.J5D?PObC5JeP
)Ydb7#Cc+^=\C^a^@c.Zd?2+C53@?@96_aZ3_/]=WS[#YEYCO8aTMS:#DVTA5G.-
HCb0#eW]Vc7N+5IP2#>@WMb(H?8ZTb.A@g=-O,PZ9<3DNGOBL.3,g&NX9-g9?0b1
aO;#G7e-(2]/.2Y1JV&+E].KI@E.G7IMfOX@-N(/>[_TEbY]#,Q:T_(Z8eKLA9dA
X7,Z[E=JeM5WO29d18d?_R)C9c3ce^.[e]R;=W[D>IP]3P9^#U6gU>E0=(;eH=JF
5S.?)4[KHW[eT4P\:0NI/ee@M=d-W:c;(dQ?Q,/0HZOWZT[9bLGHSd[;D=FBV:=4
P\aVQ?H_/QbI//\=@O1.Y+2.NWVQ/,fd4eYN5P]QB>K>+Kc0?_TF@E[_dH&7^2Y@
a,8e4FO^SC<D^JJF?EX3>P^7g-0+.DI/./:4a3&S(#0[U_B>gPHTaY0fUMZKcA8Q
.U/9;c7&>f)f0+<7:K&[&UVY&JWVI9GM-KH8\<&\6cNBDdN3R5F?N7J6bC#G?:YE
9PCg19f2.@(PAX(V@f;IDOO\bc+/<5X.9[5OU^UEB4[48YV+R6^>3_^]b2+\7/)6
\/(DHPU.VgSQH^Z<a8PZV4)=)g#CO@F\+O40bH\1/;+R;MHT<:BYC3PLEcNQIICU
;7cN#YB3(UQU,_Mc2X@)Ff/Qf:5NJQ:&]+CMK]cb[LAHBIBY@/(2MF=GeFXA#0dd
31?8>b/,)N>+)Z0-)W5CaICO6/5_?MLXc8U2@RO>[5R6gab+Pc=C#UXE^)5WD@O=
&IW0S=5FfGVaB.\@\QWWPVT0ad^4Ef6GSI4S]2NDUF_/(dI.YbV<=dS9Z-=KTM)D
@KFeYN5VO:SC?Ic&&<J@\17aQ_R8G^\/MX1J)F@1d8DI#X:A0/I_[^ZVa=c49dL#
9cS&#.SJ/_2[Z#=3Xg[X-Le6<(WG)_WA1+e)ETK#Hg=:]>Y=X2(Q2J7NQ>/.e0,+
XfE>T2+b#UJ_XPce#FB3af(]<XF@=;aHU4?HK,V:6=^QFKg[IbATWHFI,_.6Q+SB
E\+3Q(E:_^1a_PMJ8?FY[3=/W8-;X9;acZAa5JWWfZcBZ\>9P1ETI-C\3V/KHg?f
Y71FA1,^8L:)(9)0N7[>--=777TeGETbDZ.VH-C^;MM#GY=Q=+Y9d1#PIaQ97M7:
5_b^D#R_F)(LGJdMYVB#4PC<=A)NCg0</HfCDU9I_O3];K,c=U_Iag,Dc#59BW-A
9Oe2LUG^5CP_@F\/]\[2=GY/cM&MQd@K[B>Z>V8./eZCZ6JLg,:V5Q]?^LYd6U8K
IABaO^-#>aMOcf@)RbK(?cFLJ]-L6-YK#7?>aF-KB&2eLMa<>>+IF1)79[;JZ;0a
9R7J95H0KGfD.1/(T5g(UPHR]@;g)O7eOH-IS#DH5QV>S,:N04,V/(V>A7T@DfGK
W3]&a^\IY@f2SNFRB#DR\<E?ZTEA#.WN,/U2E;aB9+-X3GVL<-1;0aUXIM1MNg+G
f3W<KVNS[@;@IN9:5G0)ZQ@)I#JPEW-cBcR?6R_\X8IQ>INB8DJE/YJSeR\CS,:c
EV.2\7/1eQNfYP?d;6/:ZK?ORg-\db9dD(9bQdU&7,)?H\,b-:0_M?=VgN_V?@D?
FfGR1+a)T:::&+RAMf1K[9[K^5_:P@9R=GS&\NYMTG>TEGTG+I++N7d^9bD(S1)b
PO5:3\H;]SR(5Y]Eb?N3HP(4TNe9Lf^.eQHc49<5.2bE]-6Mgd#9?U0EX1X0K&MV
KEKgE3S:8MTM[4bSU\R&>=D\Z-404X]/NP0[,142c[:9YXC)KV>-?Gg-96fVO4>5
1H[L6C6M#O<M/$
`endprotected

//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
/**
 * AMBA System configuration class contains handles of AXI, AHB and APB system configuration 
 * handles.
*/
class svt_amba_system_configuration extends svt_configuration;

  typedef enum {
    CHI_INTERFACE = `SVT_AMBA_CHI_INTERFACE,
    AXI_INTERFACE = `SVT_AMBA_AXI_INTERFACE,
    AHB_INTERFACE = `SVT_AMBA_AHB_INTERFACE,
    APB_INTERFACE = `SVT_AMBA_APB_INTERFACE
  } amba_interface_type_enum; 

   /**
    @grouphdr amba_generic_sys_config Generic configuration parameters
    This group contains generic attributes which are used across all protocols
    */

  /**
    @grouphdr amba_axi_chi_sys_config Combined AXI + CHI system related configuration parameters and APIs
    This group contains attributes, APIs which are used together for AXI and CHI systems
    */

  /**
    @grouphdr amba_multi_chip_system_monitor_sys_config AMBA Multi-chip system monitor related configuration parameters and APIs
    This group contains attributes, APIs which are used to configure the AMBA Multi-chip system monitor.
    */
  
  /**
    @grouphdr amba_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable coverage and protocol checks
    */

  // ****************************************************************************
  // Type Definitions
  // ****************************************************************************
  `ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname amba_generic_sys_config
    * Controls display of summary report of transactions by the AMBA system monitors
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to UVM_HIGH or below.
    */
  bit display_summary_report = 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname amba_generic_sys_config
    * Controls display of summary report of transactions by the AMBA system monitors
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to OVM_HIGH or below.
    */
  bit display_summary_report = 0;
`else
  /**
    * @groupname amba_generic_sys_config
    * Controls display of summary report of transactions by the AMBA system monitors
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to NOTE or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to DEBUG or below. 
    */
  bit display_summary_report = 0;
`endif


  /**
   * @groupname amba_coverage_protocol_checks
   * Specifies number of AMBA System Monitors in the system. Enabling AMBA
   * System Monitors in the system also means enabling AMBA System checks.
   */
  rand int num_amba_system_monitors = 0;
  
  
  /**
   * @groupname amba_generic_sys_config
   * Enables CHI system inside the AMBA env by  constructing the  CHI  system env
   * in the AMBA env.
   */
  rand int num_chi_systems = 0;

  /**
   * @groupname amba_generic_sys_config
   * Enables AXI system inside the AMBA env by  constructing the  AXI  system env
   * in the AMBA env.
   */
  rand int num_axi_systems = 0;

  /**
   * @groupname amba_generic_sys_config
   * Enables AHB system inside the AMBA env by  constructing the  AHB system env
   * in the AMBA env.
   */
  rand int num_ahb_systems = 0; 

  /**
   * @groupname amba_generic_sys_config
   * Enables APB system inside the AMBA env by  constructing the  APB system env
   * in the AMBA env.
   */
  rand int num_apb_systems = 0;

`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
  /**
    * @groupname amba_generic_sys_config
   * Handle to the CHI system configuration object
   */
  rand svt_chi_system_configuration chi_sys_cfg[];
`endif // `ifdef SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV  

  /**
    * @groupname amba_generic_sys_config
    * Handle to the AXI system configuration object
    */
  rand svt_axi_system_configuration axi_sys_cfg[];

`ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV  
  /**
    * @groupname amba_generic_sys_config
    * Handle to the AHB system configuration object
    */
  rand svt_ahb_system_configuration ahb_sys_cfg[];
`endif // `ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV  

`ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV  
  /**
    * @groupname amba_generic_sys_config
    * Handle to the APB system configuration object
    */
  rand svt_apb_system_configuration apb_sys_cfg[];
`endif // `ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV  

  /**
    * @groupname amba_generic_sys_config
    * System Monitor Configuration
    */
  rand svt_amba_system_monitor_configuration amba_sys_mon_cfg[];

  /**
   * @groupname amba_multi_chip_system_monitor_sys_config
   * - Indicates if AMBA Multi-chip system monitor must be enabled in the AMBA system env when there
   *   are multiple CHI sub-systems that must be monitored.
   * - Can only be set to 1 when the compile time macros SVT_AMBA_MULTI_CHIP_SYSTEM_MONITOR_ENABLE and 
   *   SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV are defined, and there are more than 1 CHI sub-systems to be monitored.
   * - If set to 1:
   *   - system_monitor_enable in each of the connected CHI sub-system configurations must be set to 0.
   *   - multi_chip_system_monitor_enable in each of the connected CHI sub-system configurations must be set to 1.
   *     - multi_chip_system_monitor_enable in each of the connected CHI sub-system configurations will be set to the same value as
   *       svt_amba_system_configuration::multi_chip_system_monitor_enable in the svt_amba_system_configuration::create_sub_cfgs method. 
   *     - In case svt_amba_system_configuration::create_sub_cfgs is not called for the AMBA system configuration or if 
   *       svt_amba_system_configuration::multi_chip_system_monitor_enable is
   *       programmed only after calling create_sub_cfgs, user must explicitly program multi_chip_system_monitor_enable in each 
   *       of the connected CHI sub-system configurations to 1.
   *     .
   *   .
   * - Default value: 0
   * - Configuration type: Static
   * .
   */
  bit multi_chip_system_monitor_enable = 0;

  /** @cond PRIVATE */
  /** Internal queue where unique master_id are stored */
  bit[15:0] unique_master_id_queue[$];

  /** Internal queue where unique slave_id are stored */
  bit[15:0] unique_slave_id_queue[$];
  
  /** Internal queue to store unique id for each valid accessible master slave pair in a specific amba system */
  bit[31:0] master_slave_pair_id_queue[$];
  /** @endcond */

  /**
    * @groupname amba_coverage_protocol_checks
    * Enables AMBA system level coverage 
    * <b>type:</b> Dynamic
    */
  bit amba_system_coverage_enable = 0;

  /** @cond PRIVATE */
  /**
    * @groupname amba_coverage_protocol_checks
    * Enables AMBA system level cover group for master to slave access. Note
    * that you also need to enable AMBA System level coverage using
    * configuration member #amba_system_coverage_enable.
    * <b>type:</b> Dynamic
    */
  bit system_amba_master_to_slave_access_enable = 1;
  /** @endcond */

  /**
   * Enables complex address mapping capabilities.
   * 
   * When this feature is enabled then the get_dest_global_addr_from_master_addr()
   * method must be used to define the memory map for this AMBA system.
   * 
   * When this feature is disabled then the legacy methods must be used to define the 
   * memory map for this AMBA system.
   */
  bit enable_complex_memory_map = 0;

  /** @cond PRIVATE */  
  /**
    * @groupname amba_axi_chi_sys_config
    * System id corresponding to the AXI system of the AXI slave ports
    * specified in axi_slave_port_id queue. Should not be set
    * directly. It should be set using API set_axi_slave_to_chi_sn_map
    */
  int system_id_axi_slave_ports = -1;

  /**
    * @groupname amba_axi_chi_sys_config
    * System id corresponding to the CHI system of the SN nodes 
    * specified in chi_sn_node_idx queue. Should not be set
    * directly. It should be set using API set_axi_slave_to_chi_sn_map
    */
  int system_id_chi_sn_nodes = -1;


  /**
    * @groupname amba_axi_chi_sys_config
    * port_ids corresponding to slave ports in AXI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in chi_sn_node_idx. This array should not be directly set. It
    * should be set using API set_axi_slave_to_chi_sn_map
    */
  int axi_slave_port_id[] ;

  /**
    * @groupname amba_axi_chi_sys_config
    * node indices corresponding to SN nodes in CHI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in axi_slave_port_id. This array should not be directly
    * set. It should be set using API set_axi_slave_to_chi_sn_map
    */
  int chi_sn_node_idx[];

  /**
    * @groupname amba_generic_sys_config
    * System id corresponding to the AXI system of the ACE-LITE ports
    * specified in ace_lite_master_port_id queue. Should not be set
    * directly. It should be set using API set_ace_lite_to_rn_i_map
    */
  int system_id_ace_lite_master_ports = -1;

  /**
    * @groupname amba_generic_sys_config
    * System id corresponding to the CHI system of the RN-I nodes 
    * specified in chi_rn_i_node_idx queue. Should not be set
    * directly. It should be set using API set_ace_lite_to_rn_i_map
    */
  int system_id_rn_i_nodes = -1;


  /**
    * @groupname amba_generic_sys_config
    * port_ids corresponding to ACE-LITE ports in AXI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in chi_rn_i_node_idx. This array should not be directly set. It
    * should be set using API set_ace_lite_to_rn_i_map
    */
  int ace_lite_master_port_id[] ;

  /**
    * @groupname amba_generic_sys_config
    * node indices corresponding to RN-I nodes in CHI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in ace_lite_master_port_id. This array should not be directly
    * set. It should be set using API set_ace_lite_to_rn_i_map
    */
  int chi_rn_i_node_idx[];
  /** @endcond */
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the configuration
   */
`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_amba_system_configuration);
   extern function new (vmm_log log = null);
`else
   extern function new (string name = "svt_amba_system_configuration");
`endif

  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_amba_system_configuration)
    `svt_field_int(display_summary_report, `SVT_NOCOPY|`SVT_BIN |`SVT_ALL_ON)
    `svt_field_int(amba_system_coverage_enable, `SVT_NOCOPY|`SVT_BIN |`SVT_ALL_ON)
    `svt_field_int(num_amba_system_monitors, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_chi_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_axi_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_ahb_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
`ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV
    `svt_field_array_object(ahb_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
`endif // `ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV
    `svt_field_int(num_apb_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
`ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV
    `svt_field_array_object(apb_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
`endif // `ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV

`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
    `svt_field_array_object(chi_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
`endif // `ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV

    `svt_field_array_object(axi_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(amba_sys_mon_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int(enable_complex_memory_map, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_id_axi_slave_ports, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(system_id_chi_sn_nodes, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_int(axi_slave_port_id, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_array_int(chi_sn_node_idx, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_int(system_id_ace_lite_master_ports, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(system_id_rn_i_nodes, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_int(ace_lite_master_port_id, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_array_int(chi_rn_i_node_idx, `SVT_NOCOPY|`SVT_ALL_ON)
  `svt_data_member_end(svt_amba_system_configuration)

  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);


  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
`endif

 `ifndef SVT_VMM_TECHNOLOGY
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   */
  extern virtual function bit do_compare(`SVT_XVM(object) rhs, `SVT_XVM(comparer) comparer);
`else
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare ( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );

   
  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();

  /** @endcond */

  // ---------------------------------------------------------------------------
  /**
   * @groupname addr_map
   * Gets the global address associated with the supplied master address
   *
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a master address into a global
   * address.
   * 
   * This method is not utilized if complex memory maps are not enabled.
   *
   * @param system_idx The index of the system that is requesting this function.
   * @param master_idx The index of the master that is requesting this function.
   * @param master_addr The value of the local address at a master whose global address
   *   needs to be retrieved.
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param requester_name If called to determine the destination of a transaction from a
   *   master, this field indicates the name of the master component issuing the
   *   transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param global_addr The global address corresponding to the local address at the
   *   given master
   * @output Returns 1 if there is a global address mapping for the given master's local
   *   address, else returns 0
   */
  extern virtual function bit get_dest_global_addr_from_master_addr(
    input  int system_idx,
    input  int master_idx,
    input  svt_mem_addr_t master_addr,
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output svt_mem_addr_t global_addr);

    /** 
    * @groupname addr_map
    * Virtual function that is used by the interconnect VIP and system monitor
    * to get a translated address. The default implementation of this function
    * is empty; no translation is performed unless the user implements this
    * function in a derived class. 
    *
    * System Monitor: The system monitor uses this function to get the
    * translated address while performing AMBA level system checks to a given
    * address. 
    *
    * Note that the system address map as defined in the individual
    * slave_addr_ranges of the axi and ahb system configurations based on the
    * actual physical address, that is, the address after translation, if any.  
    * @param addr The address to be translated.  
    * @return The translated address.
    */
  extern virtual function bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] translate_address(bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] addr);

  /**
    * This method creates the sub configurations for CHI, AXI, AHB and APB
    * APB Systems are currently not supported through svt_amba_system_configuration
    * @param num_axi_systems The number of AXI Systems
    * @param num_ahb_systems The number of AHB Systems
    * @param num_apb_systems The number of APB Systems
    * @param num_apb_systems The number of CHI Systems
    */
  extern function void create_sub_cfgs(int num_axi_systems = 0, int num_ahb_systems = 0, int num_apb_systems = 0, int num_chi_systems = 0);

  // --------------------------------------------------------------------------- 
`ifndef SVT_EXCLUDE_VCAP
  /** 
   * This method indicates if any of the sub configurations uses traffic 
   * profiles for generation of transactions 
   */ 
  extern function bit uses_traffic_profile(); 
`endif
  
 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the APB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the APB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif

  // ---------------------------------------------------------------------------
  /**
   * This method will go through entire amba system hierarchy and create a unique master_id. 
   */
  extern protected function void populate_unique_master_id_queue(ref string master_str[int]); 
  
  // ---------------------------------------------------------------------------
  /**
   * This method will go through entire amba system hierarchy and create a unique slave_id. 
   */
  extern protected function void populate_unique_slave_id_queue(ref string slave_str[int]); 
  
  // ---------------------------------------------------------------------------
  /**
   * This method will go through entire amba system hierarchy and create a unique master_slave_pair_id for 
   * each association of all legally possible master and slave pair. 
   */
  extern function void populate_valid_master_slave_association(); 

  // ---------------------------------------------------------------------------
  /**
    * Gets the handle of the SVT configuration corresponding to the 
    * amba_system_port_id given. The function matches the amba_system_port_id
    * value given in the arguement to the value of amba_system_port_id of 
    * AXI/AHB/APB configurations and returns the corresponding handle
    * @param amba_system_port_id The amba_system_port_id of the AXI, AHB or APB configuration
    */
  extern function svt_configuration get_port_cfg_of_amba_system_port_id(int amba_system_port_id);

  // ---------------------------------------------------------------------------
`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
  /**
    * @groupname amba_axi_chi_sys_config
    * Sets the CHI SN configuration within the given CHI system, corresponding to the 
    * given AXI slave within the given AXI system. This
    * information is used by the CHI system monitor that receives transactions
    * from an AXI slave. When transactions from an AXI slave are
    * received, the information provided through this function is used to look
    * up the configuration of the corresponding SN node to facilitate
    * performing related checks by the CHI system monitor. <br>
    * Typically, CHI transactions are converted to AXI transactions using an internal bridge
    * in the interconnect DUT to which the AXI slave port connects. When
    * CHI transactions are sent out from a CHI based interconnect, there are two
    * options to connect the CHI system monitor to these transactions. 
    * 1) Configure SN nodes in the CHI VIP's configuration in passive
    * mode and hook up the output SN signals of the bridge in the
    * interconnect to these nodes. 
    * 2) Configure SN nodes in theCHI  VIP's configuration in passive mode and use 
    * this function to map an AXI slave port to the CHI SN node. 
    * .
    * The latter option is to be used when
    * it is not possible or is difficult to tap the internal signals of the
    * bridge within the interconnect DUT that converts CHI transactions to AXI 
    * transactions. In such situations, the VIP will use AXI
    * transactions and provide it to system monitor. It is
    * important that the SN node indices provided in array are not connected
    * physically to any SN port because this function will disable sampling
    * of any signals on the SN  node indices provided. The configuration
    * information is only to facilitate association of AXI transactions to
    * CHI transactions in the system monitor. Please note that for CHI, the
    * information to be provided is node_idx and not node_id.
    * node_idx is the array index of rn_cfg, corresponding to the SN node.
    * @param axi_system_id The system id corresponding to the system in which
    * the AXI slave ports which are being mapped reside
    * @param chi_system_id The system id corresponding to the syhstem in which
    * the SN nodes which are being mapped reside
    * @param axi_slave_port_id An array that consists of the port_ids of the AXI slave ports being mapped
    * @param chi_sn_node_idx An array that consists of the node indices of the
    * SN nodes being mapped. Mapping is done based on a 1-to-1 relationship
    * between the elements of axi_slave_port_id and chi_sn_node_idx. For
    * example, element 0 of axi_slave_port_id maps to element 0 in
    * chi_sn_node_idx.
   */
 extern virtual function void set_axi_slave_to_chi_sn_map(int axi_system_id, int chi_system_id, int axi_slave_port_id[], int chi_sn_node_idx[]);

  /**
    * @groupname amba_axi_chi_sys_config
    * Sets the RN_I configuration corresponding to a given ACE-Lite master. This
    * information is used by the CHI system monitor that receives transactions
    * from an ACE-Lite master. When transactions from an ACE-LITE master are
    * received, the information provided through this function is used to look
    * up the configuration of the corresponding RN-I node to faciliate
    * conversion of the AXI transaction to CHI transaction. Typically, ACE-Lite
    * transactions are converted to RN-I transactions using an internal bridge
    * in the interconnect DUT to which the ACE-Lite port connects. When
    * ACE-Lite transactions are sent to a CHI based interconnect, there are two
    * options to connect the CHI system monitor to these transactions. The
    * first is to configure RN-I nodes in the VIP's configuration in passive
    * mode and hook up the output RN-I signals of the bridge in the
    * interconnect to these nodes. The second option is to configure RN-I nodes
    * in the VIP's configuration in passive mode and use this function to map
    * an ACE-Lite port to the RN-I node. The latter option is to be used when
    * it is not possible or is difficult to tap the internal signals of the
    * bridge within the interconnect DUT that converts ACE-Lite transactions to
    * RN-I transactions. In such situations, the VIP will convert AXI
    * transactions to RN-I transactions and provide it to system monitor. It is
    * important that the RN-I node indices provided in array are not connected
    * physically to any RN-I port because this function will disable sampling
    * of any signals on the RN-I node indices provided. The configuration
    * information is only to facilitate conversion of ACE-Lite transactions to
    * RN-I transactions in the system monitor. Please note that for CHI, the
    * information to be provided is node_idx and not node_id.
    * node_idx is the array index of rn_cfg, corresponding to the RN_I node.
    * @param axi_system_id The system id corresponding to the system in which
    * the ACE-LITE ports which are being mapped reside
    * @param chi_system_id The system id corresponding to the syhstem in which
    * the RN-I nodes which are being mapped reside
    * @param ace_lite_master_port_id An array that consists of the port_ids of the ACE-LITE ports being mapped
    * @param chi_rn_i_node_idx An array that consists of the node indices of the
    * RN-I nodes being mapped. Mapping is done based on a 1-to-1 relationship
    * between the elements of axi_master_port_id and chi_rn_i_node_idx. For
    * example, element 0 of axi_master_port_id maps to element 0 in
    * chi_rn_i_node_idx.
    */
 extern virtual function void set_ace_lite_to_rn_i_map(int axi_system_id, int chi_system_id, int ace_lite_master_port_id[], int chi_rn_i_node_idx[]);
`endif

  /** @cond PRIVATE */
`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
  /** 
   * @groupname amba_axi_chi_sys_config
   * Returns if the mapping of AXI slave to CHI SN is valid
   * @param axi_system_id System ID of axi system mapped
   * @param chi_system_id System ID of chi system mapped
   * @param axi_slave_port_id Array of axi slave port IDs mapped
   * @param chi_sn_node_idx Array of chi sn node indices mapped
   * @param report_errors Issue errors incase of incompatible programming
   * @param perform_sn_cfg_checks Perform checks on sn node configuration
   * 
   * */
  extern function bit is_valid_axi_slave_to_chi_sn_map(int axi_system_id, int chi_system_id, int axi_slave_port_id[], int chi_sn_node_idx[], bit report_errors, bit perform_sn_cfg_checks);
`endif
  /** @endcond */

`ifdef SVT_AMBA_AXI_TO_CHI_MAP_ENABLE
  /**
   * - This method maps the AXI/Acelite transaction port_id and ID combination to CHI transaction LPID
   *   - LPID[2:1] indicates the ACE-Lite interface port ID mod 3.
   *   - LPID[0] is generated based on the OR of the AxID of the request AND'd with the programmable mask defined in por_rn[id]_s[012]_port_control register.
   *   - LPID mask in  por_rn[id]_s[012]_port_control is by default set to 11'b 0 and therefore LPID[0] will be 0 unless the registers are programmed to take value otherwise.
   *   .
   * - If the user wants to modify the mapping based on their requirement they can override the method defination. 
   * .
   * @param axi_xact AXI/Acelite transaction to be mapped to CHI transaction
   * @param chi_xact Mapped CHI transaction 
   */
  extern virtual function void map_axi_acelite_port_id_to_chi_lpid(svt_axi_transaction axi_xact, svt_chi_rn_transaction chi_xact);

`endif

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_amba_system_configuration)
  `vmm_class_factory(svt_amba_system_configuration)
`endif   
endclass

`protected
ZL(>HH@0b&J1HKW@4FRO4>BFL2B2]2K9OdPbe\3?PJ718X52,L-Y1)_->_<VNEQ0
d?f?)<_&<DeeJP-UY.+N;05BJH\<;8#9@N<]+PTV.:CPIFNX+&3?,6\LR2/7+,c4
A[fK&GEGWb::I;T:eWO^O)R[d8b77G6>?]GWZ/L4c?Z(@SQc>d?FQ]RM-]M5V^3C
<UGDYI3f3M^Q-A1U[=Y,F<,4cH9]69F,<?WA[;H(fCC=Nb3MaHU0IgE<[VE--V6d
@IaI]aCIR<fL(06Q[7HC&=f5;V#CTdcV=DLJ>/E12S8_b2Q0=cCd6ZV^B(53.A-2
/>#g3^BDVg94V;<Y,&1K.0cJ6Q\CEA/Oa@aP\fV,6OQ@&CbbOFZ0_VAO6dXgWAgO
1/#@NA0a+5?Xd4:<d_4GL8a/\V1L>.9I.3JD&=#g<U3.?S,0MK7P\a[=X3gHYB=F
BO?-H:@[f:DRbJNe:^(Y.WFacdK^T6OHOO6B3#>+N&P_/.(QO;<A]W4I.()SG=<9
5-WS0P;\gF<.<?+)FMDTQa\L(D6HFbNgRLKXYD+a0PW0[AX:0H9Id))9EM^?OS:&
_=1KfOZB+F7bR\#X)+H.<JM#CP,HW(1Pb6f9QU?8TH?-:OD4)_FH)^#2;<6BU:+P
,Bee0XVQg[T+AUcRO@UH:^9>Z9V@#D=[<$
`endprotected


// -----------------------------------------------------------------------------
//vcs_vip_protect
`protected
9Af7W_VJd^5TW5U_9L7@TT/YSHD-O^ddEbZ8&P7a4X/9>0PL[a<)1(S7Y_8Fb6cL
]e.T\_KNDU(6>.DUH3?eI0[&c^\=_6>eOeI9fUa=5d1L1<P&>:3a?>6]N^&32HR6
=Qg2a\\;DRM;Y>R0e,<STZ.AZ0B[/7e4)V.@P)VUD@LI]<.dB5d<:OCCeDT8XU0\
4JP[.fOANNXf2BEQ9G4:5V]/=M3,=3L0g4=?4a1EcaWaE^^c\@UC^GC^(_ZR6-<9
TKLZIe=(1aAPf,#=F5J)WO(I0P2d/gRXD;&d@U]eZE2^S;M9JP?Z61PJ)&0.[\9V
&Pd:dKW](4C:FaMcO5eMBXeG8@c2::e5f=,5ZZ[/IQK2:BNPI=6F8I=a]4L8S.G;
)8P&[M@&)9dHJ,eb9=R1&bE]5L[-PLb@_&61]X]?Q-7=2P9^S\0D5\M4dYdZFX_d
Lc42-a.&1=[8XY^D::&aU3#[K2O:g/^?UU\(U\I7]L?c8^c/EI9gFYLa15IA^N03
:9V&X2MOgZUKZ<LLOB.[O=FLT&9D6Y_22.1.:@b&b_?-\Z9&2g(RYN6GYfX;-HU8
9)49Ib5E8ZL9)(W\BgN,&EcB+2aK+-=TCSI,+B=@^PK1Cb&QJ@>4ED]?8.E)NGgX
K(@)Z-H>K\#c9cPd4=L=Acg?&ZE2&4e,<_If-VJdFS[9Y2g,.b7/V3ZMCK^\<VUI
[;B0g1PM?>5XE/35_:YV-00UBJN@NND=@WXf1XbL\eWfPX=#:M,9d+#?CY3MB1W3
_A+X+eM;=E2T8gEZCWRO&>?C+f7UgeE8b2^&d+0,]HJ,9?2Y(#<4fW6N&dR;REDF
.CTNKVKP2L7[^4^DN/:F^#N0/GI1,^cZ2#F+\8/3ZX)4.JX0?V68H-Y)?;8AA^BC
f9gR6R2(\#MAf#7GcWgA_bX@ZSJY1]Vbg,MO?0c<H^E]A./5C&YTR=))L#IT>)T0
EcK,FKG+R6_R3TO;]\;_;7IQg;23+,^[B(S>+^[\@/F0&/U>4WdK(.ZA[C.,Y\eC
Q&FDKgZ82PaM[^M53([IEVFI_[S)(Z13#-2C8:Qbba)7X:0HdJ;\)-aKcK_O2\fL
6.=3&c8A6b9?eV6&_J+0Q/PJHbJfSC9:;f>D^.:_#DW#TMK9<TfC:L)cb+=ANZHF
_=;?067^^C\F-.?MfCX+4U02A75NfTT76c@ETXe7L2O^\QC5QI^ZU^2C6+32I6_&
_NBF[/=2=KRK^#bbM3V(CI:7-\^?Z?5<.T>X9(Q_9>\[Z=FHK)Y2-&WZ(]14[/g[
R6g47,&OfXNRe3-3P]_GQ:GNB\9E6>O]P-X([C_IS5T.gC9\Q^,GT(CFL]=4;O,1
c<0Z6U?)R7MaH6\CV2RFbLFH732RMV;9<VDYceL)9V97cO6)5M;@YCS[PFPJ@,:6
GB_8&GBDf#PU]#ONJBTLM@21IQ^@]F<Vf3cS_X&d)RU>X91N5TS?OS)_=@=)gS@f
2c1a5d>58^NaKeEKRZF7L)@(LZ07(-R[,d^;#&=E7Y7LD<68FbG+=[+9R5M-aZ@(
6DX8Q<4^/adG2cZ&UUaVP.GZE4HB+aZe<QZ^,gZX.H;](?NA);.>@8,:9X[=<7.)
g?&-7Sg6A+C5<=G+\-@Ba[7PGGK\/2;F1AAO0T@f=,)VNR#/1aP/0?f<>0/X;\YP
]gf[_1:b^\-EZFN5e+d?8E,Ha>X-H,9b9OMeC)_OOXc>.cZKIOQA=64B^d/CRgFg
ES(A/#W7KIgOG-_R.GPYOM55Y>Y[eK-9)021b5[TOE5bN\K?]4=SG8aF)J,)PeSF
Y@<+@Ieb;\_Q/FDCFMeIN/J01J2.1bNIS59;9A[V\@T&JZ9&#6B3@OY=C=<@J@,5
T_\IP6)K0&^_.-S6\?4+b-I9K2cR2+f_SLF0\A0^.dAeJ))I[dbf/cL#LH)()Ja[
cUY0A[CUg?200C;f&=MD;FZ&+A/&OT-Ff<0f#QJ5PJM[Lf;b,V6Y&>,BBIPAN<9R
^UNaAY9V1W\C)Q>=[EPDcD5K:=/G\HaeW&2GbNWG>E=ZHLHLT>=A-LA^ZCe,)Qf+
9EI^P;g[Fe49>bG.\R6g7c:2=)3?I,M,H)=1@b0/2WRCgCN(Gc\/=FF/LNJVQQ^J
T(CK;A3K^)S/F.SUM7B/C;gP8U_K?7##Dg>Z,e=BLSgd]Fbg)Uf1)_8AcP?)g?LU
AO0BOY\:aTR<(NLLE<OA]&a@JE3V&P-VG-MF3&SfeS=gSRb-V&e8./N+_IReGE,2
AM-I9NV7,&M^]FART#2?EVU)&J\eHYGZ.e6SZS0EZB?1M0K))Bef0RDJUR3]Bb1c
.+K)/.8-Y8AV^YW9SCY9dHIDP1O6A+-_C=0W8O.>a,?R8R<7>6cKOc.aHGD]-RaB
1])6E?c6#<;[97I93B5^O]=I+_:[AJ?PF_I-WUe+IcCf)?^PEc,Z\8K+0KPB:4[C
cX@S;V[E84[&+?T5LaO/5RFMVW-,<(7>(<VQQ)eDbe]g,WGE^@68b)P(ad9[.+E4
,4C.YX_G9HcWI[Y81OKG.27P)a_cYc(Ne[2Z3=Q2QK:5^g)fY<>_Y;G:MVO9G?/5
L&1BUDO<\U,8G9Bf+e;R177@dUKV@gf/&g?e7fY9S?=N\)S4Za?8M^FYENPRg]6H
Y45PJ/X\[cTUAbP&F-?5WYD^6LEEb5Z=4d;@8b/0:[8WH_a\0T&9T7OPcFf:P[HV
K:W\^VB.\^]&dMD+/NSD-Z<0U>4AB;/JXNeJ8VO_PbK.1;(g<<a=?4WZS@=CJ[J3
T7D:Ka?>S&#T+_3:Z_,9BHX8=Q_&P>G1g>^RGcL@=M]E]?bC5=aGWQTEEaU-S]fJ
OU84>ZFA\/OZAfaf[LKI#88IP4R8^3P>I#2fa,UKZJ^K.f\1<7P-SbDQ/H68NDRR
(.>N/BITgRg8HYg(Y-,IQJgI6-R,;\9B;&GM2Kg)E&.\7L@d?K,@g;=?D=IBMR_Q
ZUV.DB(J@D,d=9XaL?a?6YI^_KeEYaf,^?]??=LEC9LGA46YK6?NA=Td37?b74<1
B\->4TE<X+_2+7@D:TXdUSU\1QM-MbY_c7aB,_X^B5^)K1=0E--g2g:A6T7e8-H_
.#Ee1/ECLP_D&4T0&#A0,U3a5cM(#>MKZZ2,gR>CDc(R^LA/T9cPVW/4ZDT&cP+a
DET1^1dX@3=<;#4&9Ia]6G<J92Q83)^b9^9U&eB=X7gRB4X.>228YL,U))=.:bS6
^(SAR.-&:TOO3J:Y;>?1S)=K/Y):_43ATUEI]S,#6f76:F@K2N-C[M0M]gJS=[NM
?8=afTcG#8G8LZ&M?RM5c1>A_aPT6c/&#>BH9^]C=C2AdIDB0>?&KP7Z/QMIZ)1W
9Qf(VPf5C021-]SZ,TMFCN1@[D?JUbG?5OIW9f726Y,_dG0-^.UVD8VC/[+Ic7:>
YUfAY)fFT:bH,J&#23W&1DJ(L3<Y]?UM?,BCITf)dO1gGPa8[^@KDZC32SDB-.&+
V4\ZZW[[,HC>ZFN9>,eL+5)TUbVUP<IP7/[<0&LLVd(?TQcGRZPU1PWLFR].:\GE
/8-Rd?g:_MO3AWU@\GME#4?CV^a?MA(7N^P5B-W9Q72T<,728(M[EPMPRC,X1H>S
<Y2?WGdTY(gTQO02B827K#gU+eUS8DIDE[I]5H?QSE\Je#BGL,0T?]E5FKR0I)[S
^B1b<W8[<98SN<0O/Yb]PCH\&:U=Y7E_S#;5AD4,P0+OS=HO7JUBbB7(Re#_:0FD
dE3T[7U.NWgf?FX0/,M<Q.VSOX6^<YY.T(:V\QD8)d/(0XJE9(?)_#D>QL#1EK[-
PP16UE1E&b,H18D6f5c?Xb8XfMESWM1L<2ZF9\U4?Z>#R4A?e.#:^T&9Y]/>=g82
L8aBGSa-#Le\71BKV3.DLPZD+=.a_#N^3I#fe<O9S5A9RCQ>>=GJ&1<ULbcbO]/.
\.44NUA#9CJ#ZdPc+?YgA&;(OOeW.5c49GOJ47R,2e-XQaO&\DE93=8)&GNadKO]
[R>fcRSReH4:YGMOPbc@c7NY2?^de:)@>J;]Ga_<2g_#.<R1WLYQ>7)Ieg,(;])M
eK<CaU=1KM>c:U&?93b,(EE>77PgQEU3G)gM/H-;O.beDXN&B)GWb_0+gLS\P3aO
_IQ(]K\2KOMIS+Sd-f=_R<\H_IL-@2cb==;-^,>&MN3O_8ULd@b?]3Yc,\?3DGIT
WG/#b\<\O-0#)e]K3\bHWF#Gef0UK=3_QJ(dQ_;U:HL/JNV^MG:gXLBLB5/>/^2Z
SB#8/4F\\Ra9#5PV]Q\=HT]JHOT7WEEAg[H>,c5G#T4[Y_SU6)6Sb52H9be\Q^8^
^HBN3L?M,bC]W(Pd]KDU&X(I:SX[B5S:Z.UW4RWL8MT_efMIE<CEe@)D/<Y6BSf<
?EZ9?E-Q/02Y?-VA[J)gbLOeUL.QQcKfeB)YS<-@@^^TRK-dNII:])4051SDQ\0)
/0?e8?B=J8_TRNA_B7<I6fGScU(S+X@Yf/gK2Q1+:JG#ReMJE=V@3MN6(9-^Kg=?
RI;e(BZbb\YZf-)Q<#(]f7D<.LG8K<_13c=ON2PT(fII?CUD5dAR9cb24;Hg1W75
5_YJXYR^Na91/+T([>KY1FPGdVXQSHYV5PIS5YFYMfe,..cTC0D13/>cZ#AJJWS)
BKGLL,>5^#XA[eNf1;@VO;\L#K2RRL2#SQ]TXAQ2--E:VeeC,HKWT7Q6PVD5.Y4/
fbL54I-O]e29YZ4OG>\XY:/Bc\3XTF8HB<YW)I91PT[\X1[Qf?cQE].,LL-1V_e0
X5#HgDcLTLQ.)D3.=P),\1(RMB5Hc,:\L9+NVdfM#MM#/@f8c+-T=FMTG5JXLGN(
GC2?ePST6=adeR7/;O&-dD\V2@=1AXEGSLYfgVDT1]IA;&C2._/,GKEg(I+YK)PM
7#]bbP_/fSf\)BbH8[@/K99+Rd)H]5XK^U;V:##X7UHO@<F(Rgd5Y3\L^0O&]SO>
C0LcB@5O()Y943H_cc[QDRSEFc^-XgS&])5HTd&T:\TDGLT<>]>-DG>1::C;LM.0
0FS<.0B^5[IfNEJ9g<S=^Y]76a=Zb1^:H3\EeRIb7fJ/9G5QK514&XEC^Ce;/U6H
_,\\TTfZ<N([0>;607d\g9@>Q7\#62,cM9=4WYK8)IJ3K+e[Ka8;_RNFU?_K+ZNN
.K2Hb\;TV/XH.d2L,KTV84,dN:X8c^bNY[aSTL>#=I-S5(J)[Z?2UQY1N>PKY(5W
R,2MHB8Y.OCc5f6>PH#02(UI6C2WGB;I>Cd;W+fHK1fC+&7GR_C:=X;=P5fe5MP+
d.?2G+JDO2Bc_(608W)C;P56SIfX,_#7I5QeN)4b1KMe9/0,aMgd#gHK0a:aa,Z2
C]Hgc=_MG3<H9Rb9QEOP6EFCVgK<]IU&bT:4W;+1N[44Y=567&PI)2bJJ@+3a#@4
+UaAC59b<73dCdCQT>8>V&EGT1cP9KeB&]3C4Jg;(3F^bF96/NC]J+X?O893SJQ4
?MLTQ(]PdI20cbWAI5+#dALAO;,^/>IOA3HFQabeEKf20(##CQOL>C.eGGEYYWaF
BCG<K9),QaBB<g4b7L#4HSa.[XXT)>JRXfD<<;]@,1@1F(2T0C.]5aTM/B7]gUF=
[IC\3ZX.3I[ZPHWbQ15K0BGGSdF&TFAFQ-RKDRbXK2>UE2E-,5]./G8=,aJR893R
QeE\Y#A<R0a_cXPD=Q,3)Ig;e:DQg[,cGZ6b91Fb[@I0aN/,K;6(&+#65&EF_g^5
48K:_.._;BD+&87E@]#\_05X]dEcaK6Sf73ZBUFU:G:;f#H@Y2M_,<I<3>Z(-0QO
OA<JU/0e.B?^V8U98WV1A@H?MVWCc6MAB^9L92PdJZ\bODg\eLE=;c5HP^WY.AZU
Hb[B:E):3CY8;@A/6)&G-8H2d/7=a=;;b0/;#.HPLQ.JR9C.YGe#Ab#A573S(=)+
8MTK>)JbW#EU//1)Z?(P^58?Ha2^1e>6,SLd7Db<@4<CO^M(8)I\_aA>YW23XL3f
DSHNWU;ORI:bE(H+FL5PK#NI:a;7&:_K3J?<Q796^UCU9S7PMcC@FC(3BQJ+dAfR
Je.f<ABTMZ&]7^2##ga<M&(G,2Xf>Ba?37d=&U916@G??GXYf=[WN9)UV)g1(JR/
[:O6H^J4(\^2T;eRG@X7AHYAI]5FSE+@3]?b1O.1VKAJI?;Xc7V;R50VT>O1JT2@
KRHE>D<XWR/3SVO:Uf])?@);eLKT_QFE8_I?^ZZJG,C]>GUM7-c[F[3:-SgFP&?,
YTF61N=Pc=->JE)&H+b(8KT:Lg^/&T.1VNdSZSbR6_;eEGDSbGQ1aLM;YX0/+XdD
PbMMgKHAMaX:H&A6Lb&;BL7DB.3>Wg;SgTCAg.F:A?GGcA?&VcOB1S8/2]<L=6>D
LS3<b_aYeZfN=6ACOgO<8MJX1^=f(C43=(6[Q;8;^,,e[c+-TBF_#d,:/S#E?[/&
.)(XJ#LPN?J5W(2bRI#+QU30If4IAT2)>81OY75L:<6_IXO<A1TU_cJ/):VD78=4
>fQ-O1C-P#H/5R_>Y<+VE\@OQGF,5HBC]5]Ec^Me.,>6U/b35TK3-GW6<NO.&<PS
20SP,@R=gEUVVK6PL?KQ\PGO>/ZS>@#dc:e?Q=Q53XLa>S_Y,1P7TIa[a+7),51?
]F^;#<M+R&/70d\/:;FQ48Za=].LO:4@8[21Y((3d6&ZIYJV6NMN>=C?N+-F:_]1
YK;/;P^RSX4dW)VJX;fbM9B5+-@W7\?/2UY829a80g9;bF>)_ZC_dA3=?fJGXJ_E
gXP/M?dALR(;EN]?,C,X_Ed;AB@)RZ]d^He5IfdNMH=;9J;dVa1NZ?436K1d1,+F
;+e&ADDI@QXLAb=WLJMKUGdA,Z&2N:\,5;[JLbFe3A6Ng4V]CKCE7J#2ff^JBN]=
VAQGRL0F[B#M-MD5FVIQ[9UV6GJMecA1IA,I/b6I(D>@1XT(5:]/Vc>Q<LIZFE8R
JNAg72;N2?A6KR/cSEQ^gA/df)8:2BN91DU>PJJ]DJ&bCX&Z<6DS4TggSc_^,:eI
=J6S/<FBE,^@V0EDKaBfE259^(cOQ^cSP5@;-IDE\^&6:SNJ.2;7<(L&e:]ZO>7#
=^8<A],.K&PIYe+[XFCGb./:eYO97LDBaOS-I^fBfY9,PU.5RX6=>CQe]X41NFT5
S\^AQAU=3:.^24MeR/JJb>Y]2V?Q8S_Fg1O/f+_=&DETGR7@9<GZ;G6F/0XMa@6L
RQ9=7[49.7BNe\S<],,;WLIF[W\7CO8E==a>M,g>F6]YJ.)UY0&+^<(W-H_FZVW&
&GK3GV6D1_#^ZYM.K]_8WLHW-e:LE2(@93CL\-e0MS_LaHUcaQZ/+,;KOb]LKdFV
G]cP#d1T)a@V9,e<YRR5UAO?K1bK0.4_\)?Z&6&HUf+@HAdHC2A:-<.V/4ed:6gE
]-Pe<#OBTPcf7eADF+/6a>Y)@\9UQQMX?4O?T(/#_3TX4WLCKR?A(X1KX844Ue,N
3(47C\;/10PVG6@.?E:Q]&\J(2agXF9@ZP]bI?O&1)/1>RPS7Qg-+DT\MaIA0#[(
#DY1\S\WVPXE.H9K,^+LN>\B9XM)g^R9H#\XNL,cbE@-D/&FF6A6.O\\4OOZ>e<\
O:EY0BC@W99F_MZEC->#RLI8NG8Z1OT-[6N.3.?BFB)=abKWV&0\Nbc-;BDJN5D/
W0.BFd544gfB7>1A/97],Aa=,.KY>V66f:+aA)bHK=U:Y(ZKa:5:@=[P=\HPPb\:
6F?O&TN-3Kg4DfY;PB9>eaM@,a:QNB,+dD,\,)-LMI<ZdE2Q6Z4ZN/5B=>^>@^+a
c01MJGd.(:]7.SZKVcP0Y4MVNQB1B9H2JScS:1VFEL3+0NeZ_8aGXSePe5P)41)Q
36cIF5JB_LG24d2--P9G.Id^\C>=FC\JY,42gGc4JCfd4].TbW^,4]L\#PQP+&X&
AJdW-UR#)GB(+6=KE/S)>2V/3@g?41Y?,#URL)?F7GYWM9<Xc_:)H3I9,bUX0a3P
8;gWO?I4MX()D+5/PdNS&A.J3b7BM.(8O@PK]G=;2V6K9;;V7]6I^]5/\dGPVd-Q
:85YZHQ-DbWG&T,V5W5F8POfff/76#.a(PO5AOcd]Zcd&B\ZVdFX9g=MT)<NOe?R
D^T[.,J1+KE\O(fT^SJCe>3/,[KY9>g@:J]^&YBY41WRX4P5B5D:WB3;(^-PZ3DC
+U2_@=I&26[dCbG[BA,aQK,4dO/dK78P4?8RWI?TYdL5?V,=OSCOF:JS/5DgY)FV
&A(C5>DN0YZKX5I=VV?IMRcS8-&D6LC?\>D&>=)3g<S-20.1VS)Q8&A1A8a.>7d2
5JO?5VcHVf6F:2+1U?WDCb.I=LZ?WV/BYc<C\?cf6CO]A&d7CY;(E-9a@K2I=g\M
Q,>8@J-aT7c>N5KP13LMQ&F1\(^e+S93:RKYECRJ-]5,/TX3J6f(C?9RHF]Nb07<
=E.W&^V/F^E^0WGHG2;e,OA#Tg@RV49D16Q:WOCC,:JIOU(b^.;&bbRSKGH.<g](
X&WV79^ATZBgQ?+S6?Y4B8\OR?.OXC5>D]I(Ad=L9LGW:CF&e7f/.T;W>)XLJ&aB
G5E\Oe.U5g[__PcZ,@6\][^NRY\I8XLI-,c=@S4739D@DN=2^#^L2Y4;,e80P/AM
dN16++6[;P@g3cLf<.B(fIP9T&8UQJ/#SRaM1YaOB,T:N[69FJO/)gYH2=XW\#XP
+bF6P4SSE1=G6.@Saf5gA[^<&8f=<Ud^#&SFV\3F()]1G3K=RJ3TO.+agSV0Cb),
C;=NSTA2\2OKb&#DJWIF^cT&a3a8,G_,<(WOY8fO16P1NW<XS_:OaRGeVTaG:YG-
\OK()=#/\LU^@8dc)eZ6#:6dQd]V00]-+g)IPR7Ada>DAT0^<Lb[YLA=##g4PPC6
W+#(QAg7:bY4<.=YE6bD-N23aNN:_I]_\7/5YI5)VC^?FYg]JKO&[VfAB/:IReW:
ePB(XQe.#+KMU&S.MY[4I;;OR<./Va+Wa#/4.P=+0G6dT=,d-9:#\9SHA>T5AgV6
>96(2XF/.eV7-R>Nf(bJVAdeDFI^?]K;d8=0>bF1BP.1NL=/:2W0f;H0(?4X.4(7
UQUNefgSa)X5bBY]]Q+?-=F]@c+-XUCQQSYU-Dgg6.5^FQGX[eEEYIN5.dZ^8[Q(
N7^4<;:c#N<9P6.e;+-b]Z]^E/^9(INL4?VQTd]C@Q,XC+YK<]\SG0)NR^G]Wcd^
.6B9a50.0g9\URU_._PaA-+B(:58WRbQVf:Ye#<2C#H;..5,+_][_]7e,ACN6e:#
.Y&@c@gSZ<^[/[7\a1c1\Ifd_b[?<fYHODd@Y9N5&@>aR9LYR_>.NOfdN>.Ld;+.
_gJH1cN8@@gU[NQ5WPJPM;6b<DB;:5aUcQSIdR58f@QQ+f]STOXbc7VOM#0f)XV.
.>@BKI\/+++MJdWYV37N&(6OHMXb7DM&&I>,b2WMIW[NQDV3TD\>V7Q(d9aZ^2BF
O?b:]?SU0e(;W[[ZXLBSOF;F>Q3-fL&>&O_6[ZFJ8NZGH./Hd1g.M?F3GMW&T^O0
GS3@WG95HgEdNU/F86=0K3bb>-Wd\&>/_ZN8a[\\e/S;=gI^Pg8RMe-O_\B_S@TO
)\_8&8a+LJAS/63bc.+:6AH?P(fJILA)5+@0(+OB=?1OZFQg-O(9bYfZ;EeH/TXG
\U5<.BJ^3^8E#3F>[V8KNG0]ZZ-e_>g0egBcUH1+ETc8B@6-<U)=L:a\5S(J#R+=
+6Y[gJ>D1.6[0(-/KMAZ:5ZA9V90&[)=UbfQ:AA9F.bO0H&cZS>&KY47DS@BC?_I
+A15Kg7:?KQAc;L]5GR.Fde(3:R>[&0Rd,KEY)/M[,DQ-@DU_GZZ[;ddTc=7O7IJ
^QBb^&;bcK>UMI@aP@KGB^=V=:+EJ1K4eG.AM4&Y-_OLf25c@8Xe1SE_FD/C8Z<I
I>@PLE7/fW&B9L31U^0WPTLH7]_WGbS[)gO]:?c\^(&APQL3Z+5b?0F)FS?X/PAU
.5\b[+1QbUAI17DS07GQ?Kc65IX@+Oa^<gY-9/H)g5.+Gc>Z9P@5VeF2VW@OQB9S
aQ0CBY)AO-0-L,3UK)_7=W>6dFYMYB7CQT)6XZYTfN5Q.>b(XVF]g93-1Y,dA0[N
=[H2BJ1R9)f:1cV6egRfV:=)O^;KNYU2:d+5YMDeU^36DHOTYNH5LL?A:RZ^dKA;
-6MA>bK#(S)13QeTYU)C56Z0(,JUgD-^BA#9.;D9)eC;9#a+_gEQ#H9+K71E.)3=
&?#Xf(A:9;G(<47eJLSQUSZK30V0SDB.>6CfSSMe2#U(1[H##27cL>:]N).ZCUF]
.L8f+SLPD,\ZC\DPX^;YbVN[g:1A+bG=>I&_?TIJH=ICZ;0.&>PJWUFff3B&VW\X
8AEA47KI+ePF\,E1(g1P&f1INf/G5<@.G;[?daTeI;M=1^XID:a?+<^L:-\/@\S#
U<+ZO6f3Y\PccW.=LFF\LNf:4V2:A,[O@G/<=^_9<f25AY\^HAQ=g#eETf@#eMEY
:5P@,H(4Y:-ML.P9E#S(6.ZV.,F]R^BZa4>=cF.>NUfT:GTQEH9PTQ_/:8@3^J1+
[C9BI0?9KbYW[H+f)DeI(Y/b9EJO3>.[#\2f@O#7H0VRU85E62]1->M=MSK)3?+.
X0\@64]JFb3T=HKUO@FC;M-0+(Z[Z_VW765Ub&7#ac-33eG2;GXBe,N..2;WUJf@
6gc1:3^Uc_<LTWT7K&d:LJO2J^L,g4/9@)3>)c3=D).c3K9T5-8Aa664DZ8JXZUM
##f</_SaB#/cRYd.B.<2]:LbYQga&\=^0LUSbOU<;9RRec.=FMG.PY,Ye;4QbE;(
9]S__Df?N3ORH>0/gI+^J:WfF,HB<7Y[,HBU@eU6PLC5_ce/Ud8=DZKbBLe012dO
<>:/g]fWZ\BRf,/Wd^bY4;7LOI@BAbC;.L;ED;d2NAacFbY]WD]><7EfYcXKWS6N
,6:d:CI/61(/;GV[&Q_0G9NJ)H5FLQ(Ag0^PBeaJfD_W?S5IeN-A-C[RPd;RbP2[
\eG)+]#g7W5@MFgJ5SeFcNSD]4a_90,4_<CCeN[bBXgG1@:C\D,+]2ff;^Z#9EaP
NSI/M[8@B0#<ge65Sa3dG5EO+Y3N\HgG=SUG=Be[0KSA@cW5O;P).)ER+@O+<aT:
de4D8/G6):]BOSR6L2>2T,?L</]/d9@P\.S-GSGLP3Pg:W5&<b6U6BU:c?559=.Q
MPN7I5BFUA>V=2\Uc5[AP>4^7F2)1)H-TR/ad:XIIN8cHCOS\TJX+FN6#\L_ZA/S
#d-F1Lf?J364;#ZD;[/fGS.XF+)AJ8E-@/HGSe\gB&HB]_X?YJgP+EQ.VKb<Oa>V
(?1A7g.</B9BU[-O_fC\48M9W40M^[a>T9CX^ZbS^LII2(>7KF=J/W<C13KTaL&#
_)K)PcQ23cUG,RAJ;aZg>GGPfVGOR2GF<2BPb#42_SbdD;4XC7fZ]BdIeTDfJAUA
/=?F4gGWH4-?I5f1T)W6]TR8_);&V2QaDI(BCYeNI(SK4?e\gX[eX#A@L;P;?[K-
M//)8J)bVM-DKZ;+ZLKEHNIUNQ7_YJ@1,C?4W^YTX556H7SI\53I,ae2J1EVNEg\
e(0])S^Y3QP&]1+QIXH(VDQ.L(.>f]SE0<;/g2LML^5-bga[7d-W17G:JY8T@/EH
2U^CJZDCU-[R8dD<b.fS2)UN=_5K:UF?@+[S[DSZ_G[G3?CeDdCHKBDC>L_+2S7F
+S7(GT7A=KSB\UEKN)<?GNR.CIV7>LE5@aS2Q+)EIfgSM.a_0^I-]Gbg-;[g/3S]
?G^ML>\HW65(-#\fV33O=7[/Q6bW#\PQ;MG2fWPY;KWXA5KVSN)+PZ5c?4dRGTES
BV18gP7JVfXU[X&-8Y.K:E@Xc/[.V&X326N4Y/J_a(/5Cg^CF/#P<WY3/1Wb0YdM
6O.F+-7c;K,+a3]50_(AQ0[-A@E,Q)Df56LYDD)G97&MER5M0Ja-JNaEE<L:8SU]
0[DbSN9JM:</^J#,WI_dDS,06gAM9XO9RFOZd\M0V?>CE0MTR?QWe,/X+1O9V3SM
(MD@C#?GOg.O9]._:DZ5<c&P]c#AUV15VPNH5;=56F8K24NDH#Z)\&7Y/F;&#V48
dCMPUTW^a04M1OR2B]+024(P/GS^(Z.SaTedg;aH&^e^_V:?fBFWZ#;(1aL;;Mca
6-(:B=;H@2@?=_6-d[Ac^DD\/JOUF:D)b(.R/#@TKT2P40HMQ,XfK0M9&gUea6)e
&O+803@QdDZcA.fPHK3I(IB\C:8Y]PB<:<g;J\fPG;Xb[>-aV).49LMR0c=H4)f^
:+RPf-6<179WZE2?BO=1\HRdS.F+;4.,^[=S=,M+XISPD]YGBFB4U2OI+c/9&f/^
VJ[fKR@@E.ZB^^#K9,Q]-a<(7^OfcGL4,R#X9BC8<0[G5Q8@4DCJ=J@NcYF4b:7a
?eQG.TQ8_5&^IYLMQecYM]WFSf+J,QJF4WfgK,=J]UEIP7fK+/=TDCC<bEa&W8#S
3@8gB4L2XPLBHM>M4WKMB\OaIaB-W7SS[(Ad=0<2_9dRbf=0_0O37?Ve.U:X:>-f
G-a4L&f&5WF0C,\S&,:D\/6)4aYV7ePIE:+RFFK^B=b(XeSC3)SU1cJcd.(4XKQ3
dB9&.<dfdL:<C[f+]5-3)f;3YMYZ0D[YD8F-TXIeT,:1.53HIf03-TI#fV2;;?G3
/A9L+-U6cIT9-J9HCSKMYS9fXPZgDAO[,\F<2Q;-,+F\2C<=dIf-OUbM-c<(RV\.
&HB:,<35I<bdRb0WZ:K+R0AA&RIK<Fa#8\LFHf9=56,T9a(.,KL4[CLgI1@594M0
e116DadcV.#^W]<g@;CXcFcJe?ZBXU+S\G?+[5Q[@QBb,<X1bWR<41+.;&bXIS\-
(5[1T8U\ZA4O_Q[dVCKX<(4PX.3HC+\YHNgdKH2+KVFNcD_K6Z8\(R<Q(/XOYX@V
NVZ87@[@@>-\V;]QCFLH]18L>YXbZG7ATRLcN[7+7P-XV3+0E\SG^R,M5\]EF)ZT
Uc\^GL(W-.S7-?6^AZf;I7B<@+EdfY5.]TDDXR_L3f/7CgE)KW8N,+:W&4)PV^P.
^@dI8V3c76=e\C<?^D7_@:K.Na];6Q.RL26/fK(2>KHZ@QPVAgD#Fd+Q_e=,+UP5
M:d1)bRGZE\81WG9OR6.FC]JX>3B#>5e-dNg7/L\Y;Zgg.3(&gC+N[@.d71e/;dQ
>Z^&6Se01;P=PFK_SeLH7F;?a@W3HD#7^XgU@UNSX9<D2[G9dDX1Z:3e5;K&4UTZ
.NJ,g@T+]UPCYH08[:?,_O3a9/=#F(T\)BG966F>&<Fd^B+[UWWG<JecR1e90J]E
c<SV2FNY0KV)KaUTC0OC3c^c(7LG@;RO(8IfGe?6UD;^G/Hd0LVR(>0d&b4M-8aE
b9^OcFS/#0cVgRZ(\OKPf>DOE7MN:X_W(a6I5W+#KS2f-T<7N^a9M@N(L+5<c_U2
1]DRD5,/;CETC6Z<DWFcR^(f506#>c?/K=;3e@F;T-LLc.>:1MaZ]4&5Yc.FSS.F
>N(12I(R@d7-;.0J@)Wc:0b?P+7D1_5N8+I,d]c.Z3/L?ER&DX@Q0DVK3fFV_M/7
;?RQ;Wd++,Z8:S=&7[B?gO5CTD;/eM?UU9f\LL7#<K9ANXK:a8Ic]AQ@R8R&)g0e
H7-5MT\;g[-N;e1ZGEP@U3N)X0cE:8L9\I7agg5bX3H<:&\[I7@NAI#E-fS+C:;S
DfgKdHX[-g>U8@);_6PG&UCV)UT5[JK;4[g@Iee4CLLHA#3T7>.YG+.V4\HEFge6
/,cQ@+d:,]92N;/M+63S4SX]9D;,X>d/4b>?HfWJM1BM0fLNc16D7\Fba<C=L]Zd
]IdYIIQX@cLWcC^]4PJ(T++3;bZc+?Y>FG(<(e7NO-,LZO#J7U+d(XMGO^=RY9#:
PI:GFJG-b:Q9aO;OCP>J]^[I&T:=^<T>eCbZ9TIV9SV+2BT#[<AS^.W:<S\N0[KB
eEODIIc;;3C[g.5^WQ0FQ\W>5:<f[^NVY@U@^fd9GA)&<B?I9P+L>L+JcL&ZVH=@
])M5^FB>7SW-CdGD.7^M@BQ6@K>PDK&Q6G6D8HPT(ETcF91_;A+;D0Q<C.Aa9F5P
AY-OJc1DYaXNK#@;KLT9]OQ^X]4\#C.aLg8J8<]8BQ;HAJHV>\819I?>dde_Fc-V
_E#2PS-6-eWA4S5WM)E&70LD34X+/Wc2XFd>^\]Pd:Ne62C>/B4KEFe3A7D&-0Z4
_bf2aK+BEO\[PD_R81XbUV.703O@TK;WQD-R8S-\A.Yg&Y=Ta/=F4Vd?:bK\PS.4
MU-<Q6SMJfgK6#edQ.RBI#>gH@6+D0be80dc__SEZ(I,f5@C,Y.3>9(R#5G.:8W>
C7VH@W=g2VNZI+OUbUEa:NX6&,L@,H5U5D6SW&G+.L.?.9:Q/ae34(O-JAcVUK&Y
\^.[&G1>W5EQ&U)?KO>GRWf5IaP9He&6Y1XQS4&#,8H<1a,)3PW#&]7aa7KL07QK
XOH&a(:Sbgd8C:IT?VN&He1I4F28#QSLWW9F3f26=CW7#>CbJ3Y<MY&WR4#)TTAJ
Y<@.4+Kd[g9I[(^XLA<94f+8Hg\#2eM?.]BHPb\VD#c&5>da?<JTMUJR>S\aZb&N
14_dUI.#fA7V>:I-FJ-WWUW.OGYX+)_6KP^XfI[^L-9N(cGD=EUVG:>.HH[8g]gO
D(X2NF:9FQCeOT&[g3?NQP,.T.@eU)[#=7:][EB;TOa]D7/C^YJKQOf<fN:-G8PK
&c74gKHBD3Y).GA.a+XNNBTO&/N+G2\gDO3AgaES1D??67Y(_46&_WHaVXe9WA\?
@GX;/b^>4Y:SL&DfJVZ94ZbL21TWZAf(Tb^;W;)cW/+I6]IF/QD_R,BaGPA#cVNF
d2DL\0)&@fb/FO>+XMeAL20(aSWfO,X0T\9Q?da9YD1SJ4_:6,M:8Y?<][F,1_\O
W#>ZCT8XV(T1db/SW3gMcO]?)a&H[,.T5@2fKW.5b\D,>(?+G2W0/+BN1@g=eX]4
e/#?O1@N-ONKcBBSG&0-9W,71\/bV^>c-TL&FeF(^LW,B(&\1bT1@<5)#b13?eF&
KPfO^c_)g8\>Q:T#SN4g_K:U5C(&W^:E./BVU8O4XYg,^R:&4V6P(/9Y?<QEVR5U
Y<@POd,SRPI)1Yd26K.@Td(/cG6V:=Y5H]ZQ#.)e-U\NN/@0X@,;VAHT38_QS\K<
R)90PM:MWfY<Pgc/B2La#?R0+bTVM/O#AcH)&gB#FETKI(_X#FLcXE(TOKCPWRQ4
083H)]Jf3K]JTDQE\eBBGUA\F/(&DF&7fc.@5/\H7IIZ=K4^TN0FBYGUHS&+UA:8
10J=EPfR9PJFZ<RBIIYZ-aUT+3D2IJHAG.d0R:3L7dJf_:dFfU?WLBFR.)#:b@S1
6@W>T;Od@Y(HHECH?+=Y:V3(d\F<G\,6cD9;>2Z5FCT<@g>g926N;d+@WHb4+W3D
FVH\#.&4I9gN+LSa5R4cCD#)X//YL^HXRX<AX@CU(/_T+8eGL<(@?fbcD/^1(\Q@
V=#N:S(8;H0KG&SWgg7#c\WO[L<I[\a-LY2>Na>XSQd+MDDMM4HTF(0TeagYG]>-
0(-<D+d2+YSNVH777#IWQOPe^M6\AR/&Z/EO\@QJ4KKda,NH6a<C;6\R0G]J_^Q9
LB8ed+;+[R81KGD<61.Z5EEZJ78P?+^)cQZ/<>&f4e>74([>Wg-_2W)K+TMUgC[U
Ff@FKQQ&eBABSYQVdU1[)IYbYc/N/YbOfUC^-0ZYT&V,SfG6I:02F6)=K1@0b&XC
]LI)0,RT>Wb\\MW3g5AWDf:AQNPcCc3B//ENX5)2<E,f=AO5ZVT(JNKU(ZF2TCbe
W>8(U7HgD_V13O-KA:PXa(g7->&8>VIS:f[^#5Z^c0D4CS?(R>77^V+_,/\S#bEC
M;UV<T(CE<P>3PUaeVcZ>c==\RU6&Oa;?GU)aIXY]d>)[DJbF:Jc5&W2>Bc#96H:
_YeAddS1WY6BCBcG2E@eAgULN&96;)gTE-++JcWZ,b?GZN9TVAEM-1f]K40AE:I:
0eBe,0ZK\\F(6>,R_6(5J;@0-caDYJBRQP.ES5RH72&MQA_LA5^WFMXC>K5g+Y-4
D]E>[c5\6#BEKF4e=U5gW-bNUUYFdR4TJ=H[L+&D?90f]&]X2^;4ca6PS[6@44I,
;T+A\2YPdbg_\,QWAAYP;=]b>3J+@<WM1,([8YFb-^+OL)1TBgNE)9PRW:NMN#XV
QT;-.OHD.GUICUE\0KWa&T&]./:@6PXg88ORG^QGe:B>BZ(+I8e#aR/-39SB0#?K
5JTZOAf<+ATU\^+fH^K-DUa0dKR7<2O#6)8L1#4R]GQY3&#LcTKYeE\X#J26=_+T
5W5;;9aJe6O#../SKJeMALVaITU;)b.[@GaPV?7\R5(dR:QE>;g+<5A]b?#1XA/@
A.N7-[aX]OWbOP8YbPR#<+>8M=L8[cE,XQTB>?CggPX.5XT4H#\DK>][T>1Yg@CE
9G/3OSBB,>V;E-f7)1c\<g&&G<#):RNMEL/LEARD5eBWOLR)-I1@Z_<>?<,fc^2\
(U>&NH;O][#1+UH4AU0=Y]-,cGeY/AN/+FC?L28O]9TcG,P?C>Rae:;Jb4(NQ\D(
-7<+9bN-)4^7BITBZ(;GC4EZK@[#7_:D2CGX\\e/2M=3CX^>5U>d)T1;4G?B?SD[
<KUe;]BZ:T&MTdO<]4\1^Q-=BIV=YP,:W4VU/?W^(K,#\aQg(d)Da58CeS5N8Y([
];00(B)>X/10aXK]d8#f(J1=^b->+]-=X/==RF<(7=8TZG7Hd>),HJ&T8\1J01/J
C;P/?KJW_f\J#IGFI:02@F/XNZ,.E&2WK>:=fNZG\52?@(RE&E0#@KPcP;T2Cff[
=DX.(+SBgdO1,5O\;gVYa([68<#N=g6P2&^L1Q;Ha)\FI/X3Dg2D+?+AKT:>8-N_
DND4PN,NAN,d4I9DD8Sg5C5)M=9Pg=a[>&0=:7&?;[W.:Y+fLPeSU>0AAM,\8JGT
fT<aVP5L2.-[cA8=DM].f_?K_;KW8b4H[\HB293>#_/AcaH\4<.<YV2cSf+Sc5f^
G)A@T(0aBB<O.1@R4)dURAR(NQ:4MF=7[ee[Kc[:fV>[e.VO2NbKg=e&_O5N@NQR
-(6BPb4DZEC^TZ:b&CD7N-?CG>W1J+]5]J@32&P&5:b9;e[68A(f50(M6^XY-9+B
@3d9_fdD@bTg71/II1ENS8TaJFJNER[.K^J7UI+Af?dYAYVI4;44?/MPC?U>H#d)
a@CE<&:g>\,QJTcWB=M45+Z.O&\W2?[0J@,Q.b-bL7f;SX3435=F2,7MA2?=U2+d
R@>4Z7Rd[MA;cZ3Ha7#L4?b(AS\BDD8>gIXaUR?_0W)gZA]b#.K\A\((QN:]OIbV
fQ6Pg,b5YC#F,.gADOQ97cRD0-\4(_Y2\I>2;_9B4&I9#C3U8eSZca8)F7c_\/\W
2421XfZFT]PSU.8\3-=C9Q+&X0.M\fHWXS62FZY(474\V>382WSf,M_@W,,(b16?
VCN,Y.Va8JKN:T:RI65GC:;T&K5SM-D^)R;>K[)UDaFSAEXX(G7SK7b(?>/.]a6;
bX/7F3dF5/d=D,_>)/Ve@aP]ZP)VV,F1,gU4Y^S7>L_)Z51:dG[Y9a2NKPAbJR[5
@@(OaVgbR6ITTaA&-H-DBEDeM<5U>/_UaPG&:V6S7U:_51,;SZ_8;ORPebJb+NXb
NAJKOG#ZP59?YPRN5B9;CW0PW.9ORJ[J)Q/AgYW<G?V<:Ne_]55E\(N^Y24F-SU.
;A,ASL;Qe[5Q:RST[8e.-(9_7dNQK[Ceg[d?HB@2d<?[a;8HJ6)YC4,4@3UGHW1=
9Reg<5#c,=ZeAE5EW:Y:AGIOSa6(A0Kd8Z>15R@EfYSM7:&D?.);1BOWP8@;CWa^
U,E)ebB?7gaDK<_gDXHVa)c1_b/:V8-PE3GQa<g([([E\P[ac)^3MUa(192;ATeX
XQ<.a86A@EU\&-f\@Q0bgFPBFXg?809fB?6Y3-1FP?4aVF)b@]GQMd;TFIJ+F\(g
7:.RS>bYU=(;>,-OOS=gH8NM9\[JACM@RJ7NO)9WIb\Ce274W8AAO+gK.\/]L4-W
[FO@NW6)f<(S9&H@&I62,S;26b.LVC^JT7GL(,c8R,-H7Vg:1@c,I(DAFa^[I0@D
YL^L[WfQT+3F>;X^T_7_SgWGgg0+HCTg34V6:BD-^QS22PS(^LX#203IMST.=S\V
bF;+_GMSb8/((AW,D73-eda]RN5&V0TZ5d\D-NJ;U##,[;27@1_[.?M7-WJ-4/;D
KS.CA</b:U\<-Y4M(:4@OVgF6&XaReJD4D=;[?+L5SX>KR47f/FE84O&>1:R\_[&
Q4NePIA@MI\,,S(0A]P6=E4_64@@,M5M:WRI@)AT?KMeNEgFBBd6S2^V4YKRO).]
UT(943X>XWYaDCb02LH]+]V1H/fZ]^GKW-OXUG_)]6d+Q2-,KT.Ma3)>^5f##CAQ
,?]b#M7.(PRQ<U,eLRgEH,dR.>@F#@.d>(0c\f1f^?H:J_Q:EX:1<#eB6+F]F&Vd
271g7.DQe?/3D+4D:)e/&gU8LL2LGC(AULDBRMKeSAS2>Aga1@#Ne+FJ.CH<da_c
1bX)+bV#4a2eb^.c(R\0eR)].9BdW8-B-CQTH@CSaTHRM]J_X2.?Ve@,4@5Kg?[9
YQeaGGVT^]eb4W9IE2U)d^3N[_M0(PVP^-.IY.CE<@b1B#Q>a0M4c;@LF_VALY/0
d5-8(A(WMaLcB6Ya3&f]O\-C<E\WUU9ggeNEKAJPddDW@CDE,50gc0PUeLD)K2F]
ZE]Y1[b1TINDUH&42;g#S.<32/YFFX92R#1]MXF#DXf[bQM]]PJ5#P?M[L8/F0U5
MJ<]9cB#6D\AaQL3@(Ub]-S5R8f)QZODZRL;DVG)##Yd]OLW/)0>]:][Ia.CG7=F
_Q;-aS9L8,Hc_=<INK6AUA_5a\\_JM0^QB;Wc3H@4T;8LVUL;MNHa[JLNe\14R8/
USTRf)dPP<NZ,KBZD.\T&\==)I\1@#9;+=;#1RB&^&[e/>ScLKf0UFPT>X@+GNDF
.,23a^f:LZ;#;(^-OB#XZ:<A4gEBZ9_a1gP_VMK^BP;fW=O/F;@IJ\OddV2C-]\7
V.40ML#Y&g95]:Z/bGMPQ68IDL(0=<XJTU[R8XE++MOPYXf>GJPIW+E+gB:V?IXa
&RK+G++g;HLJ64,KJ@[G7eI+g0ZHY5OY.VLBU2XR+)Ta346]7HD/PbP+\(e415N/
6?J)?(X3X&dWccEJGNCcWPY4XYE,Mf,dS,X+>5):K&+^6I^GVgM]bC7WX5?<G,WH
4>@8^2>ggW/I60#PX:d-@J\_C;A\SY@&fPRMf^bK+K<&:eCLLX\9B^06<0BTTYaC
MOU;J_<B,3MbLWFL55]f_8F?7FQd?4:G/fRXO^G3^+9;S;0GCJXW<4H](RPP<I:<
E@X(=5CB?G9D\B:/-)PEQ1H@?YE8?gf_^<,DK]L#X=T8dV&7I)=;FFAd)+5/Z\D2
=_KK4^fXJbWA020@R+WbY[D&PE<b#7/KYZ49Dd+RX]&9->f2f>DGg>1[9G@8+9UW
4SIQ+Y5^)VS,[9K]8F\3KdW_2EY9;BO.5_[3@X<?be)6F9UN^)(1g-QP7BM3gR)3
4+?UA_)Ma(@PC],-dWW7E\HU/_Wg)\f8]5N0I95M/Oa28E=&N0,]+B5PfH/]W514
#LMI]G2K:@E,b>Y8C_X^79F>8>FUD\.OYQCU[9,37-HEDKS<S@M[997g=(Yg8EFS
OL>^I#6WN^JJ0JfQb3/<6S&?,(Q,4Z;:L#XQ:.A_0bf\g=57.TEc,CP7?(#V:[c,
=S1;_ELL?O(bV;2Ne#@^eF[#80HZG5QQee)/FS(^=DfV8EY,/IU>IOLBK4]#9GHE
6A24+^U\TQ:F7V\gL<W\O9I_(]]CO6?FI+:W,NWAc0?C<[U7+g<AM],4L]=V][>A
Mc/E+f(9Y6:FKeQMa8F0Q]QJ-Y#QW(ZVOdcVb5]4(?JZG&MND@MA.KY:&:P4\b>\
+CS&U4Zea(bQC^SU7F66[8+Vc[<IFc0_=Z<:LZN4Z65C6])N7AS44OR2<Y11>#-M
VB_dWU#\I&FAOe0I_&@Jb\;<94VR(M6[K,+>-WVR02_8f@,gY<G_1X\3&/(.cdaJ
Ta?A/48XX=MEDKKCE3H+4VG(c?76B-7RV71DeNI8A=9)MQdU)185[MeF\?cH7).\
?V^8WT2R,ZJ9cf[@CP09P>9]Mfb8Td/(-7:0YBVb/++_9&1V,S3\W_+RQ(d(4P8Q
<J):IP[\TET]S&ZA87gRB?,B-7]TN.0#QZd80]B;&(V(B1\Na)90QR)_LO.71MRT
<;D:aV<O&dD45\6)d>2\2TXR)Mc5]cJf7fO:32N2(.]MLe54-]_33e4)-[7Yf6N9
=\[SW#L./QT:.OB6J>2^FG\ae&PYYE19R/gbO4_BbG]YO5aK&<@(=]a,.[:AeVUJ
;@Y=/N<JNB@G8[aX;7_Y4)945\;/cC,3P(J;DU8#6YIJ=,_dLN94f?>9<#O>+-4>
RQFLA)(U>A+5SfS<]Be5,Y9YJXB58b9/5(,O-..bIKGXE0PT236dZL5\?--TKDe/
(6?LeAJ?N@JL3.O^c22?<+=27K/5YW&7FK>[=P/gXXO;?^QQ]1UN(2.VdDKQ?1dG
Nc3c@gB>-6E?G<Qb5X&;/9YTR]2&_\72Y_<a23b7dUZ3@/QKXdGWP85)g_W?D)I+
WDNbTN@9cE4ITF-@T6?2_eICAJ4:X^G-<BegM@bS47</KTGR5#LbFXQ]cYGdXS;<
^4D(_1.JRTN>?ZbFEISB3L4DJ^05dDOU^]2IE2WZ[P+I==V19G^3S[6;4]X]Nf@Z
BWKH(B741<X[>JRCf-R,ZSO]_TMW;#AA92V/XR@?[+KF1);,65Xc[aI<U#K3>X)5
HO=V;WgO>9_CB2SXP?Kc^ND)OI]0Y=0U&>^JgNWKLXJ3d_5BJ_67H-.^_Ya(:A2e
Y:4Z875BN.aIXFD1PDX3\bPJX5db#B7E,=^5<=T2KJ/Xe\=D-<3NN&A@?S^-,[O9
-;R;V=4AQc081gPJK;G_X;]D/e_7;C14\fSW#&5C2F-/.F-Y5ISDO5W4UTR3\N>+
WX@DSa9>DEb+0U3-NE(UGZ3Ke#+1<4<U6-Mg7MeRP?:E+(Yc(b4Bc.=1>[5,)CgR
gP?L13?^U2<)LS1=8S8@E.R1FBMcT>]:T,d9bcCa]-F<2GG4(H]A^#+E:f(8=1JB
L-V2@fcG/C?P;5>[d/@Q6ZVcBBdg3\+2<3Q/LE=@2S:(E(T+.=5P2g+(=:W<>LZb
;KZMP#+A2(4Q;JO>c1Za5O1.REY16SeXDce\XMd_D+AE,/Y^+JCX&L6[ROQG5EG5
MY30)AL\R/gZ=M>-1#0DLKMA5Ye;#;7Z8+#7<7gAK(A<@9/c;]5WC3aE36K]KSVQ
+E,dOH&1W=S9X(BMXZ]D\17DLJ<1&gc>6:;V=S=TN&5OO:GM+dK##R^SJB-M.H+\
KMO4f:7)VfLLA&B820?f^F_9Y?MOY20\(+cP:<X1MN^8?1<T4D>@;X>7dc+Y4?2G
05XH+(];dLa=;FZE3MNS0)S@H1G;LaNd+KK#,JR8CddOOD;cUL1@G]CXS(4;AaIg
<ZZ\LTF>bK>B5T>aM&FU>>5YdWf6d#g3d0\Q+_X3Q+b@\H,)Hd:I)3IKg(,2EP[c
fQBQ_5K@ULUQ-\84>)D5^AM>0HUEcXK(^0^JD/?ADNV@6XK4feZ-_T1I-IT<8<R1
DLX#[7C1aWeAX1g7]E.ZD[Ng3R+dIXNaL5P(O<MA8@,#aET:<FO0f5^,AdG]HZea
bOdI/OD5BV8F?5Fg&17UHLfRbHKG_XD@fG&O4GD\fg>6HO5#&JK[gGe<V#9>/geF
#GPQXGb>W<W17fSY-Y]1SD2^#aEGIC]QI6._Q6L<;<bA.-GcP8<O1;,?T5M[RWda
H;8=?cOTZRJFN:U3F.S]fX9;KZQaZ\?BMB/=E.A]X[_^;Kc&ggRWQ[=_ETIT.]WK
cXDP8=Z)7G=L2EX.d/<0Be-bBQ6-c>E=&7J,5]^Rg6I0,RXf42(RfR@(3bICUa6R
S8+K?O@XS#F2+]6cP\Z+-1&UW&OUGERX]P&A:dYU5<=B>TMRW0eJ2&HTJ9CTY9?O
3J..^DU6fR&;R4d)db<=-._D_B;>G2JY/WMK@;KJGH/TSACL2e\GCLaf3f9Sa&DD
^QZaB(a02dQSM,0TW5@b9TI&VZ<#7\fg.MES6/L6]cMa1O(]R4?Z@XWX7_+2A]B+
>/3EdUNaV8>(F:K\CK+F45<+cMY35e0Ya9XXUF3Yg6K2&T1LYfW_\(CS/@cMI<;Q
ff_3]cdAdDN<,.L&&7DL;[;4P]5g@OUK/MTCTMG<_?&&GQ(P5&F-ZK=4dN\edg]^
M]HNO56DPIGWBP(IGY@7fZIeH]PWgK9SZ\3g7[bWe0(;MDAQ5F1V4/b1T?5B_N>Q
+W0IPeKG[aYS1^+EKUXQ+W&9BNFYH\B9@HW.6;Q,>0Tc?fA6IeDX)E5C36]XD@eT
MfTJH<5aO\67^VOb^e,IQDUK):aI\eaDY4;gaG\#ME<0(J^aC](&]GA?G2GK;a]W
3]^)gA^2:9+L/&f7>Bb\)1INGQ#(a)?@AQLG1DWWWX=?GB4WB[AA#>4N(MCcASfd
?(#>,Wf?H@9eC\G@((>4K4,.La22[5(/,JHGL2@;_F5H4Re/dE_JOUGUMM<:VL7]
,,7KGRN>F+1&;G4@ZN72-9THVN77F[2#JaM&BF#,EBY2C8=X6#MG[L,Ib,T79XON
A3gJb#=S@>8Qb=W2T)00+W>>XMdUA)P&GNN8f>_[Mb(T4TU#-@)LBaH1UdW^4QU1
OES_TWOMY1)RT]b7;AN]\R&#)eS(MNM7WH)2:0S,,NP.L4eKW]DCUU9V9IbK-AP\
gUL8YQ1R,1D1G[#4)8Ua_WcWPZ2AYLI+M?[<P1\YfF5S+[SC?,U<WCM+QK4CP:bZ
1KO>b[1>K^GXKdG2>/EL&4U^:S?PNF5_C;&Xg4+1_&V]#8SHMZEG\<FBD:O075+c
1b,.#^g_>P&2d\d(\BQ)dM46@1gPR8ECRb;^3,-\=fKXX+(>AZ[7W9&0UYH#ZJcB
VCK&@TN9:RdH/9KZ&dEYfEBH?9<8B4f<G0:+=T7R2>U[/b&J<FAP4Ub-SH]CdII]
7<RB9)aR+)UA99S_/S9VF?2]Af)9GUVWc>;;_>:HH1Y0<Rf,=^S+CGQgK(CZ=5R3
<[bHHHgeA7>9Kg;C/dI:.DTA&5.Q6&_f,SEMNF[6C0DJ6/C_WXM-VT:-NSM7[_HB
N/0QF#3W2\EA>9Q&FP)E??3CL6CY?/S:72g+A;<F?]/gJ&UXbaL@UI&2M8]_^=UV
Jb?IKG2[f0.FYEYYJ)].0NgZF5/4,7D#)Od-(Bd&_Wge=Vd\W?d/&-Z(8;Tg8CFI
6_EGJB/Ia0S_J=M.aVd=<[^=H>aFOQcW/E,g;?<ZUS:__-?6,(EgO_C;6::I@-I(
,4X91fVH7_T_)c,[e8G_)]@g^/.;=R?@#,UHRZOf+aS<)>D4B19A8,fe(/M=WCO?
YM0CM1OM2.W<-aW)(25P;L;BA7(=]0.+,Q6a.G7(.VA<.dKE,)]UBWe\58K7BCKR
I7/BWP3]L6N_cHP=ZK1bFLVEY73cfM1>+9HC\/#:BF-dWV:K-:)Ya_:RI4SZAP+Q
Q-6Q-:WAHf-W/(#LL30ZAFWP_<e,ZD]7\^\287_8V6\QaEa3KEHbY.(;Ya59N7?5
+0?QR/+]B+=&6+T^7;KdT?RLBG._b;FA8X)?CH):g=6P:.^X@fV5@8S4NQCX;OS^
g26HJbfOSM2K=T&T[Pf(,@a2^:LA^9\1R?,K,0\O9d_K0;ZJ,LJ>GL@/Qf6eTNSG
)+:_0#J^N]4)#C@cM[XNUg#RZ=T)D7?\O&AKD>&ZEa?9OaE8dSBYf@-_^cS(OE+U
[[N)91>7?.NK#XDASKWNb+FW_[<:+ZUVdJ=<OM>U-RNY;95a._<958]+(>K=R/SF
_?S?CRMCe5<O+\Wc_+EY96YVY&#g032+XN3cV-bK3=c8SQ6LfUEEW/EQ8Q5S@G1d
+Q+gC1b\QNE.^-:_H4bQNQbH071IT[SA[eNRM#V?MF5ARJ<>0?^VE]46OOFX(:Nb
XB?+DMga)XYGI8PZD<40-H3ZVOMG4LW&Q7869ZG]3][c(S_(-/\-(FHU_6d0bJ&,
LI03M,,XT6>FD2dS?,HZ5cTPYD\BGP4NW[Q(A>.2=VG78W8S,Q:R==LDd(Icd@H\
]@B2(GIEc^gBSECUCbQGU7_]X7SH&3LBE47X&g44KURVYM8=5=[<NTZCb:gI3FG5
dZR;RPUA8c)I(G2LN#;K6Y@49M9W#57CWbC[<B8M5EE/]NJ1@2XKOG6P,2(-/3O.
]A;\4aQCE\>GY@1-.._S-S]d4_0R(d-,O4b=F[UQ8)>J9d^ILU8b-)V=Md+8GPIT
.,?VB&VA.\/^B,bJW#?WX?4.?-8+-CY[L]cT;H2dV\:L;8G40M>(JfWPV[:eVYW1
Q<J73/L[agQ;^K9U6:fa9?M=O1,-^&,1_Z<XXS>#J/W7&]&MeJ:^La]<9@Nc[4,e
.XMR;;/OZ)_P]D3YE2_.+aBUOM]cTZ&]R)+LIASE2&#J6aHLGER<-F3HRI2/VYZ<
B4:WSCEXD3^IA/A,_)2&OYfd.@6R>790c,C_g5eEc4C<I@OW+E8W+<_NDJ0UHZ3T
BUY21PIe7)5>:.W,T6=>TFJaVD[Y_07,4G>FW]6CZc:5X14]VG.KK0]1^.K\7-f+
e]QYeJ^>=E9_W?66d=1d8R2SX?D\,b&_^_TEH_.6OK&G@L]c._<&7\<<d=_\N,Kc
/CgVN@_5BQ3TAddWUFB[Q/&RMT-QF@CC.N(5:5,4RW_PK0T-2L6bb[A;JJa;<E?Z
A^aLHE\Z9.KgCNKA95F@0-GbW6:[<ESMgR2LIPE9JMQX2]Wb-UV@&^JN7/U:JD^-
;f-VK8J_VE@N8RXQR1LNM<?0-8Kg:T&QOXB5PX@(aOGACaNY0E.82YQ@WKa[EX97
_>U6Y1A44];[K-2T3EUb1dNYL)4MgZ6#/T>c74WE#&.V#BT7^U[=?HS5GYV&E<R;
NU&56DEQ.-HeJEGLfBIM=^D9\H:_SOGa^78E]/g8#_^\].JXTdB-8acOS;]\<ceN
WfQ(?(&TF2ae0,@5D>5T<Og/K.Ad?c@/_Q[4f^RI86#f1_/MQ9XV&[<3&09_M@B<
RYN9[&P+H7=.b#0,/,U]dZR[BfG733dARZO0JBF1MCN1\\V@cBQ6-CC53gG_G(3#
P;/LaW/>4#LAXacS&]V]Z_5L2Q^5+J&@Fd]0(]U9&4VS2^)gMYBD36Q#C<@?c0OH
G)N,+[H>@?7G-O8^/4C1;SPDZCJ_IQ\5d_N(<9)0aP(]DfS@0K0AfH]cAEEGUUJ)
=APe@EX-V)W:L[F)06.a@68df@af@#W4DG5>\K=8A9aecK4)4=,),3?XCfR6&\4B
C?^.6gS=[gNR=5S]NIN^2<4+;Y32-V:=IggJc5#,f6M0V#gNDFZ#1_L4gTM:cMdK
5GbJBK\UA_W^9HHcN&QLHY;YUX\eaTH42[@NfI>V/a]=(c2=J-M<^:0aY)M^_16^
R[1G].&5ETd8)W&T5.F3LE?e?.Zg+4Q2?C_YVUCMMS-VZSa>03e+V1ZA/P:b2ef@
9&XG1MV]1HEZ_JDRIT_^efCJY<a5>;43E8PBVg0B=N_;8Pf[7eVJEe=YTSeaPD7M
V)_ZQ?(KCbJ>2T<3dD4.A#4BY2eKMb;WI[[EEV>.YgN>?f]CcP9g.B22R3O;2CG)
CZf;&[Aa=7,9.,f\L^e&K@,9b@PW]SQ/Kd.1[3a:>3C^3R(3YNYaW,E48;T)YbCQ
\,@6_,S<,cIDL&bC/<1IS3e22X46Ng=+bS/FAQ@g./?bH_BXZ[&B(5@XB.bA/S+H
_6b(bG8f,(ROff50\7528_Z3,Fc=2<6N=Jg?e,Eae8_DF,4a>M8W#M[#Vf>c6RaJ
V9;+HeK+[g=-2SXMT66#?0Pc@0YISD]&b.geC@,<:73[JH<VR9gMCNNb._;<fVE#
/E)K2F+Z8e@L21^R>=3K4?HC\<NIFXgOY^P6b(G9W9c8IdB6HD?WARZ+5g/T5R>^
9XL@4=BKg+N#E93[Y>R11)TF)H/<c2E;QK/8W9##F(EBDHReEH=K#&P>[.V[.e>5
EaY77(+;Q6D#gDKCS\#VfYP9JT+7B\8].:I&<J.[N+I/USf7b263\1eU&OgQaK>5
\U;9]MZ>@;FE/X9aA93-bcG+OOIF(;XZ#]W/[)cWG]@X@?(]_AXM/TC(<HVXS>TR
O/d7&1T(U__31+[]b(BYZ0]ZWH&M#[f-/V13V6>4RS=FF0>,]1g1ES.&fIF5BbbE
cCY5cGUX9_:CIO+<2G2=O=O48&PgHSCY2B8?S4[=+]Y6Mb)eaH&\e7a\D\?TP)QQ
:E1:A?,DMS#2eU&,:J^X=SYK4<ZfO?IUAF=?bLg=-@:\J,(7[H?M>ASQB]4Y6W5+
(FcI&>./I8;=DP)1..QZGQ28G,@OdR-K8/.&0[/QY(_#59ec;#ZU>=/Tg5K[JXX5
H)J-TbQQW5A[KA#ad<VaKeA2RdEbR:1]FR\YL0&@?;1PY[0X4FUKJFR;^Ig(:)<V
,gD)8E[3GgJUBc-PA9J5&26O+ROgB[[Y4H9SGJ1Z7\\S+Q>aQKU9PFd?@Gc=@85=
O+A(Z)aR3UM6?^+5C#@2DJ5WGWKOd1L+AL11O,GZP\]BD&/?YNX>B@=H#=R/3+-]
<KT<LEYFUeR)QF<\6=Ze?bbdcFaSIG5-N66KPTOb<URc^eHV.#?e^<_+0]WF6[Ve
@6-[[&T4#@65B_<fgA\67f-.>Sd(P)-\CcMI)73-f=JCdYXYMe@?\#7[:PUAB0g/
9>C.DAUYZP^WU6b\LDI,&T(?@1@5@g8Z5K4/e)TP595+1V6_cPD<FG>UZL@3WHYV
N9#8>\0Xca?J1[QH3bBW7SI\<4Ha-Z,>#_&SP@^ONQH5dG)A4gXAI:0(R.?,/aSH
EYVT\8_eO-2bMC#2d3Z&#(QEdZ?TbgNAde?F[>7aY;DTREL/T45-6;Tc]Rb>A?W]
0JMW?G7@,BVJ^+ZRR;GGOAB?M1b;:>CC+SB_JODO>E.,)89Y,DN,KN\YTEV61)#?
TI/.=d\W[2_(S0?4dU@R9TCK,:[5TZagAcG-D+aE:5NJ?:.=87c4U6&/J58Z:fa3
CN,T^,R<:g2V(8\7aRK&J.8+gb^8T?;c)YXgF+bbaE..6JM^5b<BY?cd&FY4^(7+
WRMH.3&IE?6eCOF&VO=/B.O\+>eUb4fY5\R5TeD@Z;=G0dM6G?LH?G^Y>+I1HQ;+
CfLQI\?4Ef_[VgP[,^/PDRPUCQ=32,<EC&Z&LaF7HEVO,:-^d3SP9+J2P(&G<61D
:e;)-9SeAYUJ#A5/N)3]V&Oe2N4JKBHZN5K;L2gB3^A8)DR\#P.c]Va+6X1\RQVX
eKZFC7e9]dJ8a0S(WgBf>#9+3Q,Vc(bOKBb_)/e^QQ,8Y?I>3B)8).9270\:CLeN
>/N)>4,e=@@/F=98F0LB?S71K<V1H9=#;8P7b(_LG3NUZTY&H0OVWb^-Nf.=&XLU
F.BF@f5KR.[A#eO>PA),<c9CZ23V?-bI;R_1#^bFFS7@8C\5UQdeaWBX&,PPeOQ6
+?R\T#)E=89MOc:&,c8#5DPc^BHc2[a#?X]+8PS[a5QaV>#1A@QX-5F_AX,daX0[
2fNaA>eHKaCdGMDeD.d^J8:-Ef8HI.@EY\/I3HP2BKYaV.f_\PN>T0JWEg#PG[\d
8OdKEHJ4XUO.[-UOCW>7O&I_L]PJKV>7YAW2>b@8,QeB<+7e9-e_O=RV^TCgO^5-
Eg>(\?;V;aPM#bF1?<R4T+bG)Ea]-NBCX4LX5?6-DeRQDW-GbRNcDGbM]^+e7.SC
7\\T_L;@];fc_UUCUKLSdf-&OK\ZU:FN&Cc],R1^&a\]]9S\8M\;0[a[Q_I?#0:#
D+26HG^&QcE.EIU2VGKB#P,e3_#KT8SYcJUC9b<YX11AE5W-1R:9C[=3gGcUR2LJ
JXJU1a,/[Z10E]87A0CB2QSS[3P=+Nc;6[e+ZYO/=(]2@2BOLJ/5RA;5fWP;9.<.
V=MCH8==H8(;S9D83#NQ8=L/ZMIFZ>b9eV1BZ;[PJNeGE(+-J:MT5RG:JbgOMcVK
0]LPTf01R4f?8F-g7+.Bf4QfF8)_5[.QXJX]5M(_JbaXZOd3IJ+,A^g/QA/L]Pd,
9BRB[R76S[3b4XA][V4c<WI1,e)6TQTcBGTg0NDd)&6]]:BG0-a<4/I2/,^ZIQ<D
&6aNWB7RL27_=96BZ0D2X2]503)K\T@gKG/M-]cega1_IaI-Kdg1VPbR-Y1N-7/A
P1f;V;73(R+G#>61,eX5S-EWS7QYb9<X71M[HE;,7PfG#;6cM0A4M[gFZ091cU)U
/[.J5Ob11/\CgNU>PJ3(1Q1A>^9+/E<2eb?HXK4Y&UDe.CeZ)[e)_J:A@90I]\K9
:/<N6KUeXG96AFPWb2fY<=D_5]6/8JE)OVDcO?EE&/\a?RUO?K/5QT;+aO62LfJ[
M-K85NAf#-0])e]<>a9f;SfRWcP:\__/_T655AaaZ>R+)Jc/X<,(^07?1G_XO1a\
0/+TXA),,M(,0WRA8A7M-g/CZIOY1-SdNWWC(DFP+^T35fa<,EUYB(E2e.,I91Nb
d;XQ0]Z+:R&>JEVC>GVbRS:&++>E1@NQ)ZH<8#U@g1D]CYD/;PT>^e-f[N@ODS#=
OeF\S>/.e1KJ\76c&#AY2N/RcQg2RAZ_EJO13&FJG7+ULc0IFB=Q1JeOQ#Q0LQMA
/ABLfa\?)9Q<GB@ME882QJNPS@/;U\fNL;^[1^^X?-aCK;18KFPcWJgQSGGQ<aJ=
L9Q1#=G:?W^K,0Y,^[+GTP<Y[f^UaB9@:.)IP=ZD#:aP<&c2UI^9T,SA<1?+3@ND
:]e8/L9;#R>JbY8?1WK2@?b^NdX1SU_KB:1Y_Qb1eSMb01WS[XGfC.R<@;-SOQ@b
6^_9AV8D#25I_Y2@=Ode+P#M__X8>RWRHMY6V2\/23@BRBaY^>LFJ>Xb_3=<80J_
+U,^C+X/XCJd:.SB.57DP\NZ.LCS<M@=IGD:&Q9ICc=?L\JYC<_d6B/OVIS.B#6Q
&6FYO&MF<W+>\@009PffYDYPH6<3a4eD-V?0OIVM-L7:_(Rb#2GcF\+J@3GAY3Zd
4S0B_bK2Y)8&Wa1/KRB8FP\3,,(6T8eB4#__.>2>ZRFU-B<AZBeE6IB@GEPQ[K^O
@<RR/Ccb(M(UNN96[b^XTce=Z:,^@3577N=+9fQ?]2RT??G#]KQ+=O6+H^XB=HS)
Q)4<^^_U+KY_Aa&YcQ5)8fe3X6FGEOcY/LT4?<\IE[aC\bL)CceKb_Z7J3eMZYJg
[5Q#E6)?M>egD)2^/GS1?>E#=/K\QLF9T#;.(@MTc:E<R,1N@@NaLES_GSeRc>Z8
\:#)^08g,b&f8Md6;dNND=U]T+KZ5a169,R5]3-L>3DXBVN0MV&:.5Ab.P_K,P0]
-@af4E2)C<S<&<3869FJb7Z^:L/H(D6M004I6?2O(GKW:/\\24O6:aXDTL-f6.P-
],IbA>,.V7O,9-DaIGW_@Q>U[_aN1_BNdf-C6gB0c6L0D2&=QM5R[(/32&6fcN^M
9>,X)+I5H]1_X?9]8c>+^XF7#;eL:G04[J:ZE]RIUYaC\ZV=a)d6<0PRJ7):72?U
Z4&VVZX<<W=5]P0d)S<WAAM)#-c,Ib<TCN)+OFC06Gf<&IgD#:4TeD_5gcJ0>4\O
768ZJ/0KO+UT?7S[FAW@L2TOW12;.W&@MHPFE2C5(+/+:YG4;E=IH:R<&W]bM6(W
6;C8&4E[f4MBT4Y5TGd]64R>,&QQ36M[B(cU36Y(d)YOD)J)B/U,e71?:7Z:1,HL
Fe7.6PLH5C-?C_56)?KC]11ga_[,DOB&[<IBa>28g,,3>E9[EVEQ;b(<MBf<,NKL
eM?Tf/INfLKF(LZQ1SE2QT&VH9ZA6U75J>&5DIU9H47S1IFWg?2>ESR=M5E:#0d-
3bP6/DVEaCW.+XKOUJY(faIcJ72,Q:/412&>H(EOdH0TZKba_D^7V.PE9(7bSb/f
#db(X?7WgEb8\O,K:g_<?8^5-6S]O(M;21SEIB)FMOa88P;0PF=VNf=,\g3S(I?2
[^0F7-bN48:U?JO;,510U)P&b>\IUB^3R+6#QU56CWG\Q(Q=LQ\gF9F?KI)D<#>J
]&#V6]=@(CG6D123M37J&AFB2Fb6UJ.-M.^YBB2OGb/,\L5NEV<QaG^J/>4Q^]d,
5BIZ31BQXG_9SNVNc=J(IG(F8#T2JF\XVS62+@C>eBQ+),E2<_f4dWCCVb5_0[L5
/OHZg9P/=NbR@gPX7(7B8#FQMARe2[.7G<PAP^1UV7/c(Xea32NN_AdBfDKf21,L
@+=D]0=e+&S&6V5HAII9/;79<G&cf0J85:NYc7cT2c+NY[J9H<=^T2B5>CGcaAS:
ff3^P8<Q3]Yg6]_e+5RO;e410PVFeGYb2+WYf&N>Lg5Oge]R+2egd_DTM-VK,d8P
@W.7X1:OLTWX0KO5aRc=5c?V8Q>IPU=f7bXT;+aR?CNb4@\=ET?0Sf6X.--]PNYA
\A?@>==KA^5(6J.S@0A3V6\7YJBEILIG2[ca#<;d&>(^feDV-?Oc&W_V_RBSI3?8
1?<T0XF,SdP(HE_S/67ZH1=;DW++>9@L4JS@RI/X7O8HRRNVb(Z5<GG60R/OaD1/
dHRBNUF^>.L^VBg43;QKe.QT9>XN6-&++W&/76_9>M^6_E/_W1<6;-W1)O_D-;PJ
IL(QW2-WF\JgONdg](T[H,5C=+N=DQ5gF?SZF#0eCe72&>YKZRP<>HaJ=]d:TP^.
Vf)OEK.J>3P/HcXK_c>]R)RT8f5KW:)2fAYHdWR#7bQe6Z/HR0U_;PD6<IAZWBJC
)eg?.1C2RJbU6+?&(\;B88SdXYNE.+^<JGN;0I/H9fE\/&EPaVfdF;bCS7527LHH
5)GJ;]Yg5gFdY<0COg6PaYK98J6IS57P@\8-G]E@NFPA.<C^6)eR#4\&=5PMa_OQ
2</B;DEO,FUT/WCa0a:a/FH.^AAaB62>N56HNI&b;fD<fEdG9BCQ48[6#L??fKC:
YX:>)^-O[<;2PeUc+KP[b.N+N_aQ^V_eR,F0:>KgX3K5)Oe#.dg\MMOP<B_<-X.c
,<fb=N<E_&DE:X9]7WP7YX\G)SXB8H)/N,>KA4cT7/C9JSBe5dPfRVLP.\>?;YNL
)E7[MH^IX@;\7;[?=3aeO9d2ZK7fWZ?F5_3T#72>fA_^[b)+SN&M:C@8SIg;[/E1
^YL<TJN&)4#R6SG)fgc&QEHO]^d^<92;]geKF=FfRTCABZfM.4]CRB)P/UeSM=Kb
T=FT([K.ON=VO^^V5Y#eQPK_J5U7R76DSgP>TI3U7:9AP3NI=J?R97KU,Q(a&?P-
350X8gQ[=KQM+WZQER0@;:;JNE6V9D]ZJL8)g5>^,,>UbZ]9(HE[L;[(8D=D&d@T
Je]a?,7HQL2R19RDf2YBT-/ZJeOEPIGcX8+;BO9-3VLZ&/aO&4F#^W;#FKNEfgKa
-=MU1#DBB-5.eJ4H[1(&WJH:<bVVN4#gN5L944^2A\PeDP.TF61UE=H.V.?.H664
Hf8;[@];Q\FD@L8F11D#CPCg[649@HXUeRf8f.JB&_f3]3ACc/D3RK9Bf?@J5EI:
B=>]LI:;EYSSWG:eB:])1;H>_,]V\;](SAf^P&RO2fKMQ<U:cI<Z)X+0cf8DNPN7
3eUAJ)WLHF,a@?,E(c#9(+;SgIUIB7@PNE^3>(b2&5.C4W@IcI5(a7OFfEYb1EHX
9L;+>?/V\-0P0Lc/4eI0^TRJG(aL\0S_.\+HG[^DBYZ1:2IW-I\bQ_+QMO7.JS#V
/Z,aQ5VPaH;^(K7YFY5#D@\MF6Z&[&UCX@SH\57JSRFFd[W,AWcG\BX9a##<G_ca
]PZ(+S0+g4;5IgHYeZEbc(@&F0>=?[CLKIWX#\c#[If[,@6NSAf:YIZ6]F@Z7ZWY
dWbE5QbU\4P2^:PO+XC=5:?6bUOZEY<Y]=aDY;Uc97#WaSZ#c,\NC1d6aOSgJ1.K
4&:Z&[9RAZ^cH?>B>I>F@b1fWUWT3e]IWM5\)O;DBaY8:-W?cbRd@ZEaF=M.?6b)
-I6.]XFTN,g5+<N^_^IYB,5e<<9@HQgEJGE;IJ?T&9E96[=#-2DEH&QV9&GPX39g
Q?ZCfa&AM+KV4?]f[fCEGKFTFZd]))_a1<GIN=^?ZMP5NdUN;;_8]?D-8dTBBTNE
&S.E\5-5MH@3f:I+_:Z:7-=TBKG&.BAJZ6=7VTAD1L.FA9Cc@HMBHHR?\a0,B1?B
bV8EH8Ee[\:\>V+I2e_;<gF-,[E:#0BWN9dfg2gX/;8LJ78\G:>f_4^DfHXc,b^[
=gZ^41@:-QT2D[1Yf5<9J^B5U^D-.REA-1AFY]_aJ+V\b+ZGZ0A;;<B)EKM5/.??
Z@=GEKeL[RFe=^+9DTbFN>WdX(-;;Ia3-[gbOd?<E/^UeFHSBfWb4JEcCJ5I^bf0
#DSDBJ;&\B=S9NeU9H(EMY4,c7-DNf1C&PP[I+gB6&?eDcV[A9=g\6aL2(9=IOL,
TXD;DI+3I5LM7bK2Ic_ESbI6YSJLa\9.g<)fO?H(fZOI&a=H:IB4AAFMB00AgO/X
CY&.VSYTCFb9>R82)+#F-I6V_2MG,4\^,7VSW;FE+=.4C\O+9f9g4I[_K4^N]>]3
<S:@MB3AaM9)BGgJdZ7;:;EU]_SEQgW)]TUd6O+26##[+E&6X/g+7>?MU@?>G=H4
&=DWe4NO\SF3:e8)@-Tc70OYMVb7<?[dAbNVM?9F/?cWPc3A-X4d1Q:925O</dXT
eB-6T#P@CfDV_HNPEg8PHPC84R#I+AFCG(fcJXXN:O,>GbbRXfD:M8,2bE&ZLbV_
+Gc@F6CW1&RWN6fQ>MBOG?6gM;P3I6[0GY[(#S;Q8a3;<A.GV@E)D-90a@>GEDS9
H^-B]]CAVE;N&+)JR1KJ=HCOP#J;N[faV31VMdRF=bE6-;74@,)g#g>?H];(LDc+
If138d]EgX9ZU2c_)b[Hfd+OK?:2,7\K/Z;FGGYYNPUdeRS&U\W]2D5+17KHfM/C
0Ke2=O2U/C8(KEdKSAA[dZdDK+47R@,;TNK[F0A^QJe>_V7;7dAI+EKAAg6-6d>B
F4NWaP\6)VKV[+Ye?.&ONK+ECV7c+IdfSWDT?[-<,Y5/7F,15]5F]fYe>6ZRBTM4
.fIeKW=P5G&UcZZ9H^BYEMV9[URbc(U9J+\BWT,)cBY0TeV7W>XW=e57B6L;A_A#
e9^\SKWb./?Hd\BAdTO]6/@d(3.VR62<&^VO<<b(8I2=CU>57?56O5?@6QMg:ab1
GTfA)DEYO59=)<M_afI+a69aOP]47);^0a0M4.G:<@(JZI7XR9(]X:42\14N;C-0
@O4@BcR=)9L[e2-Z.d:-MMV,Q\KFc:SCJ[LbJCPK1LXS+PI_UOf1a3)T[fb@<,e+
dQ(D=59],N46TN/JRfZ020(P2d?LCe&T=4K976A7K:Sg<T,Q3Z1T9&+d04+D,6dA
/YF1:1Z>ON.QWGODaId87gOeUQ^DH\2YKZ]80J1(\&^^cdYR7c_H#HPIb)UN?JBD
)NH)V?+?eTYJd=EaEODOLYb_2[MEKU\Z@-Q+;)8b#<.]Y.=6O2/FLQDQ7/cRM;_G
^gOccE;OQHV1&P:YO>VUEF\2eeJg21VcFA9K7&T>-W.ReAc3U^@_W[d1-4[0XQBP
U5c,\NP9+4^]e;39I,a&Q66F2+ZfZ6<IEI77>#07D569>#N2eP6VAE>E1gVd>QBU
7d/0UW:;+VQAfVV9YDB0/M/@L00Y[?B&^/@&d\5^7Q3ee@IE1fMQg\8;6gb^HO3a
I6Q)ID8Y>RL<K@1g753PgJW#Ta0F+@@&:B/5dL^O7FEF(e_54XE1,?RBV\5&fR):
Z&0?=5@gT6-HF(Y5+1L#<UU:AZS73Dd9FPQ(#/OC7R@\?(^[LEP)6U_04.UNGQL0
?b#&8ZcgT7/4O[80F:K[QAYA,e^[@PXU(UL;fU(D@Z)eE&\@LcA6R,,]=LY>?>)I
(f\gda=7GX\(N^(5EW-3b5X(QfF?G]Z,7cc3SI.W;SVE</cC#(fIS0-2#g\dM74:
_L;?IH:<C3,-#PJJb=@\8E^:FGC[8>BYA#_Q.Zb>6>:e)N[G^.:\9aS:;bY)1,3e
NfIS1[PO,BS^8&1,MMbT^g7K6PFa[bV6)UY54ASML^F[]a[6b=HX4LK7[^^gYU?_
ODU2?(E@NI[=]G3B0A6RTScLRT_1;:)EH]4P:ZC\RLZQIA\\6<^-1^DbM94MQHXV
Q/]=,ZeMXa&c1BMd-Ac?aeWA_L\+[VL@]@Ic/FQ@aU5K@c_)g^bbI>3?-4,&BS=B
1DF6&bY3:DgIQ?N.(<&P8YcO]<DN43VFWUT3[Z37G:aP@;a5>_4/,c<4@ZVOXJ61
0\&>-eYbV/,^b6\N(&3<[(gT<9bfJ1Ydf53,&K7RU7I4=fZ[.#PGW_@B8^d<,IU.
gE56NS-5BPPc.IeFH>9WB&#S473+TP4dOQSEW4#3Ie90+,04Y]S:95T#cf=ZX8#^
a;1?HdXY<fG^.R#6aA?,J;CE3dS,#aU#VQW0\3-S_?+I6SB7Yd2-38DJB0E2de+-
UFLM?cd0>N4FcfRGQ:PL9Sd_:L<AMQQcV3>b,f=F#0Ub&U?)b-N;Y\f7,8[4]#3g
(AX@1><.O1a7GW4/H.@F,f1/ff5f&1)_22GT=-@TGcZ62F<Fedf@=.H9.#SKG(UN
c<0);IdA7PX\HQfE\PYc4L\FPd/KO#egWH/R[8-g<1^G-,Q-[J?e8;+MEB6KRB-#
a#L><)H_(9S2+J7dKVI?AN;^BAW;?V@<&73DR+/Lb7Ng59geR\aQHF32H<ag\+dQ
]^<DP]feVAg-ENG-+VO-)XBUCfW0^<c?H>6R<\;)CBN=+<_VfR.;B9\G^efJ]e2^
/H/&NVT3(U37Sb+RMLU)DL2N2H<@DR8^;4V;deGDVTd3c;FD+9:2.a1Yd[fB7Q-A
9IO5#D_SEMQ@/=QP5=.dC#,-VY9?AUE4UJNGL_dMd.6^E@GZg+TWPEeeO/E))?I+
Z-Mb@(2)-ZGK@(?TY2<#Y\=&f>GN_C[U:]_3]8R8]Eg]dTVZX)ADN:MI/XWX4L2;
HRcFL:T&),<BEP;;;PVO^egFZPF/G?8[QRaYDHUc4daV4Eb3(-g?6-X_a01OWI1P
4RZQ@F<C9a^BMIU^=\WeB,-V>(3#6E4ACYSEfW0E[(Bd?Rb->[-&K^]-.;=6QO#F
WPJ8A?Y/4OG;=_N<K0R)afS2:gVFOUV8I>ICJS:1UHM@bW+@-FBB?H7,X<A1KUA,
(<;)R@0RH#d=ZH(JL0K2dPPP2]\K-?;5D)c47@e\f:Ld?KO5_K?A-CC^QCc;ZY<Y
3-E^N\]8KA31Gf&8e(YS)LC@\U6Z.BF1EDPA25.W2f.e@fVb8K&U,Y0AQS?:2TEK
:\72N+(VQ.=)R&3-CD/@<f8Y5R]+3JgF)YBHF_ZKaf]7?PRL6F<PU/(LbNB3E(gM
KJA_SC>afBacXf]>E4f;(B-IfaLc>V<b+afF1(B\:]M0GQf,O,&RaU51-D\Z:/15
97a())9N.cQO4Tc1<.T5dEP5+RX#;A(b2[C_2Wg>KN9#G&PbLRWNFI5dJ+0fM6<,
O\,dLcf5b7abKGRR1dL3G=4c\)fg)>I/.KO6T-E^N,Wb7_A<70W;59fF68f>N,aF
PJ2;T\f?9;39@6:]aec8Bg[,-S=.K8+2RV4\=I=9&N6ZFdSOQg@[edB/dDXMYb=P
2Ba_?K6YPK3&eDE2)CQ&Z3?X)AWUK7TI4JYe7]fV-gC1HQ=&YF[cG(<3XER1e#A,
H+G(+=T7ACDC?[C?KORKa.#WPC(M=&7a_7+]:<G^AE1R9[YXXd:gfPVT3?WDHa#[
FC3[7RXT?89.cT&#3&5a_EK_SVY.,Q?<eB,d6c^_ZI5f,P7(E]^?c(RN+c&bLQ,]
?>94QQ(d>X(-03]&.=+\()^d1I<FbB[McW0)NS^&PL3Q:c:L.DR2(e[HbGQMWNG<
OE(5]0J1(@8I2E4A1>IF>NWS?V55_F02[_.(7b\,eA/\_gS:K=A6I_DDSE@2b4A,
RgW#EY,V<ZW0PMH::?&-=WREH@?^YbX.0AQL\S;>DP(I1VU;2,/N,XEU1J9>Tb)E
O7^+KIG6Z2=EPId<DSVDd[]A+[C4M[eS=2,7_L+YH1@1eHMXIMFZTIWOY>c?GHAC
S@74PS+EQ5\A)e?=)FZF\IX]^O-^5RNB&+,S^<235(^JQ_J_G8\,g.M)5<_I]ORg
GH8g4SYc1/[<>>9F&4<7:&PH>TSee;G/V[d-ZPZSDf[V_MZBN+35#0.J8MNfG^5<
dDE#&YGWO0<]3Z)RBa;M,)\a.-Q8U@B196JY7/(Aa:R)QBGN\Z^70>KAU^&N(dU9
O&[]Mc:4?^4dP75Q,28J9/=X=^D_Q;ccDEaVgC93OB,)CZ1)9DJGS[#Y6g?dK?7)
)[K.8/aCa:N&?8YUMJIT],H6BdQ#X#98Y(6EG_D[YgTW.5G=>a/;WYgLN(IeI6G#
<5/\8f8+UN38G7e3L=EZWD;Y<Vg3>A#>XbA/3H0JDOIbQRG:3WWdC9-P=eTZg.-L
B1H(Ae.68MC(78_/TEIT.-9fY:PNbT#X)3@I=8UD9DU5[?6?J>FH>(X88.#cW;Y2
/6N4Q-BVfZO)1D9,Z..BLO<VXY_[T_F_7e+,&2Ef?X?K_S++#5Q#DD1Qc-C)[>JH
T.8GZbF<(2P)<5G,H-SV:D3(?#VR]U8V]bf]X#HQ[3NV9E)feZ7?)?04/R>_2[4V
>3#,P<4dT=(KB+=3<>MV:-A67&0OS^T(=E/P<FHH@gF/12P#\QfCG=M)VJgbLR[f
c:T#:E=T-X#KY2R,,2W@Ha2Z72J7?Jf,4+O9#dc1C6CH@[BHbIfX,>?XBe?4Jd<N
C.T-0;^]Xb42ID5,_f_TIT@b=-cJaK<]b7U73^0de0C2NF=-=,ZbEGZREL+^Y&H8
QKfZW>Eg@FW#G99[PSVa-N+?CU..I_#UP@;#^H<]0)2^LZa5D_.bNK+^>IJRa,/#
L;H2AEO29QAE]GPXGBfe^We;JdQf/1O<=009)F8Y)&LY>&L]3c@3abU:C\?+EV4B
(GfN_VOHe6LAS6b&/.B,gB8B/PBNCeJ#?d2&5J?/<,.,T[cKX4]3S5[(#IJ-(EG-
\NV];6>RA(b(X;@K5EQ5NY[eIDbQ-\d6@-ETDA0=3&L^]1UU69R8)b2I+=QZ.MH0
?Y^Xa=db58d4U7X22_,P)Q-)<JC5F]X=fWX2JGc&C#U2.L(?C89NDJI)=BL#)L??
#U?cNAaQQ(YfCTJ4KGY10G@4YGaR6A7T[JLTG3BFB8RTB+-#=V_<+/6&8cMBQO,;
S0VSZXH3]FX[=HR>TD5O9MJ[]J9Y0f.-[VQ,NZ>M,4;NA\))0?aIXBdB,NYTL=QT
ZL\[_ZA:V7K=D9\a7T[EEC(Hc;WSP9MIMeBXYRCY(>7?gZ203D0\f_IM=2[E1.Gd
F;I59FKM+<2^&IS1<=D2c;C:Z+^.g.GOZBE1eA+ZOTDPeaJ8@WUV1R/;1S//6=Ub
\7UU[U#=_PB]ccSLG)URM-5bZeX_U_:CC5c<;\dOHF.+>Wd3KOO8c4/a=g3BDZO;
eK>9W-Sed&0MFS;ea3Y/c6261IO9#LV;PV-1[CLN/M[3d;B_^3\Ncb7<;:d_AE7(
ZLBVNXHI#Ece1S90L.;A.G5RV-R:d]>X<DO>IO2&#<A+8OQ5YA-/Y92DT>1#_DO#
/Tg2gAg,?cI=P53^=#:61#78V46-#>aFZ/2L^Qe7eB,d(NYY//BcZJZ:P?<d(&L#
<?gLIDYY8SJ,4DT,F7/ESI-S2HbV7_0Q2TX(RO4Ib;c0U;H?KQaE,(487?gW4NV@
HTL6\^+(Qe?X=,>eU5U2?Y5=I4fQ&=ef]W2D^e9._Y?N],Y;f=LF^B:2,G_++eWT
3=>&2EH.IK4_(bA7dc+dGCWVF-Y6D4ZB4B<@#L2gN)VW\LE5P:AKK^ZU:P]8#G58
FY,C4<^RgGDDA^N];\PC1.&2WMEW9G5,0^F]KM4XdP.eJ]PT(NaM7cR(,8@__Nd1
TP#CLRII@C267R;4_cJN3YDK?]1Se19H9LPe]7T/.+dd8(<092I+XV0F0JH#3X?,
(N^E),L84CT.<(d6\GHK?BGAA7MD,XePE.JL)Rc#1C3,HELRR0EcYV_1;baM5;I)
-_XBN<49<RZ5[A_JR:L:T)C@dHUH8(G.;EX87V73FMIUe7#e#R,^M[cC:G[43]+.
.<]V\16R6YOTI[?QM&0:1U\b>,0^[YVXOY[0])-6:&AQN5LBg/::+90[JB(FVc^?
)X5W.(]@,B)fU.T59+0S)5^f]1F:8:80RDdeYDX3bJIQXWCV3)E(&TR;7A^UPW:5
U9Y\G]c+83A?NB4E-g[d,8a>;H<.)P.QgU)cXJY9_@^cS/dRD:O&6@d](IYD2[(A
+HKUCK=JNgKeMAR,RI[403G)-Gd@OfcZ\/K9g6#Mg=C/3050KR_cYN\HU\06+>aY
U)S<D1Z>LVQ8gAWQ/N0LQ_-CWUD-#VgFJ>Hf0g@1?:U)KCZCGDcD3O8I&@(MM,=Z
SfI+?eCNH_]fM6&\<\HE<?,Y0\Gg/0TA)&D4^f#TY<\>0KQH]G[/KGIITa[2\]:6
:[/#2TW&VCFH\fMOe\#_3.R;(XI/L\WNP39c-5@DfZ[/A9=e_b^Y,2_/2DMgRZ>?
VfeX7-;.XdR)]OZM<W\6-KGR1<_O-,WK_?:B6IC,c+?KUZGH8N094KgQ-[:&@?+-
[_K,&SVXBSH<HC[1V0OA[V_L01dGeHC?6U0^DE@18]OSDKIaLQ)K4@(ZH(@&9@M8
K<SEb>PFXM82+:\4\Kb/.#1<IN53D+VMHgGN<ZY55C#1gfbJUS@4g_]_-BgZ660E
>1X,J><NSB#@A5HOAHR6BVC]X1J>&I.\c\fW0\J<V<(?.;SR\Z,6^FGd/KOJVZ0^
AQITaC\#[JeY4RYMCWL0L30g:ABgM9?Lb#N,UceW(8;O+2Q@f#;;L5\cKTY;e&Y3
dMMM.;a\QV=3RB260],=b@VC\CQB\UY7AN(P8B+49PdVGJ6fKN?0TL:-PT:^98eJ
1Mf_S(=9::NN[8Y#Bd,+UFH.B(,g\M:#J2+=\TZ1a,FSK?<07dQLVE@;,H#&G,NV
^SIT<?A<NeBHU:V+QY_GJ\NXcT<gAQ+0FMOg\DBeON9Z;0GQ]<E]=++FJ]Q&0C6D
8Gg=R1[IEbac[1-?M3_NTLg#+8dTRQ:^\:/,>fY@d:0LU<O5,RCV\a\4<QaBB=Z(
QF9=2?KDG>9\MQbb:.RPJQ@+@V5,^<&O<5>+.CHGeG3.:RWYBZ.4NMbd<b9_G@dQ
:6MIMdLP,Y#fU(MbTPF_[:UP3A(Dc]KSE#2g8fa&gD9b?@ZWGSBd3GcIR\3gCdMX
NHBN,CR(:,6KL5Q^Pc7Y=WE0N66\@edR&^3(6J,[,:Z=LaLXbc>BfIfcTX?+RE0=
-N#,4PH,aAH41#UUB.]9F=B-cTL/:+8N.d.2=MHaZN35+[^C>#)L_,J_Y0M8b0Q;
gFO8D96S0GR&cbV.9XX=^BE(//JeR.dCCF4(5#Z.:>_(Mg[4G=8TbHVbZ<,&E:,N
H&+8RDWb4WCM5Z;HMQV]]C3XVJe7e09?acR)&L8FEQIJ44IfD>7NCE>K[-AS<L-R
Z;G/XQ#1AGd3.cYPFLR>_HFUMeGF]-fCbeEN_&daAc(REIc]24;-1M:=W?>dT0ae
S/)0KL7S]Q,PO3d(MC@752,<9dFW5ADP6ML5QgO.d0\6<.:BQB<Kb]a2UB47&4UY
E/7@89W#))If1BTT-a1]b6>J#cKJX8[^=fT_2eLU3VT+;Z)[5V)7aI^aDAgHa,N&
@P(\PU9fG/)Fd[1#945VPXRQ5ZV4[\+P3aJUL[,JRB&fP.@2gQT,U&]3<&-,>L8Y
9E]K4QF9V&T#_A76R/(DI>BIgf2aVQT@NM<I4H5;EQ>D8eeA>.e]fV?#EXHS,/_a
<]]O?S1;4GD-fQ6Vd^^.fZ-ScF#c1J9d261>JJC/9@\g4MZd#_6;F>c6V1SQDC4_
SJJU?MIJ:T)X1?6(KdeW2#22Rc#SPMF0Z7\&+d+-I0DT2VUd8b9QE_=_;X(PWc-?
_^Yf#=/V,>)SbW=G]#=c;daZ3^d&W)T&e7;ZT@IO[AMedM=71\Ub=+N(AY;0FYd;
a:55<>5-QJ-b>fEPOA6#9US1PS8Yc+;WQ#\F&f-DEd-AX><V+&LY:41b[5/E\)\/
4Ga.eTZgOQ\T2a-]WM3>;9>(LcdfJ#08A-;Gb,;0_HKcJ-dU@)?0N_4]@LQ9RVS>
KN]gHI6a0UX=K;-0NUY:UdPX6Y5R;18O7SD;#>-.=Ra?)(\KRUBcOJ7\-f1.D?K4
C6eCY(:5AO)G)O5JdOD=RHdaF[Z:g>HV0,#P#da0-SX9W:H&J3^1XaTJZ4UU,W1b
6R\QW=8Y?<N\5<TIc@PPC)Vc=#P]0_W@NYNV86BK#gb9WY,-[W<M?.5c(HgC[..\
6?&QFeUeOG)^Q0BbZTC#^e=0FHa(B>/0U9d&1+DR&Tb@Md=M>eB^Oa7.;C>DcMbB
:XVIg,\O6I1FB[>cTR;,3L\]4FdDc/I(a&,H:Q^RZ#)2e^WHc&I(+Cb[7+/McW8\
J8bOOE6+9\QWWd()GMGaAP@SK]P)^1@d-,5(MRa.SUF2^U/Zg:f5;>H[+^CKT0Fd
S>00g?HAHP0:DSg^Fa],;g+QFO1YJ\WJ[Uc2#)Y<@(6;N&S<fTOXZYMM>I9Q^8@e
KM-,]L;.J3[@SfE4CcaMfBg8c02HQ0#()>.CaF5CDUEGV/]DcC6VD7@P9ZEF]5L6
aO&[0TEZY:=7&^VHAQ8IT7Xe7YZLdBVQ65B7T\P_=7f[Q^W6_K7O0+]Cd6-6MR:g
0N]S\9?d;&D,^_P>.VY+U4fG5>+RDdS,=G)DPMUF_;f<(LEX_3+Z7:@c._Y[/&<>
(:70=KR^HIRP6[3EY0Ug<_b+JK9dW+L[aTZ6D,@W(<TL_/W-2YBAbe\G07c,V<e9
7bD;+@)(N?H]<Xe)^6TGP?W(@(L([>JFT?2+PKL;K)PYgD;,Z6TYD(.FBe?]=1#A
A+:TI@;[O,RRK@gK9_,cgRG\XU0YQ?8II60]aL[I^=TYRd8M0_E108<J091X[)D-
f?#<A#Ub=VOJP(,Rc@GHK.4bcfTF\Z\L-ZX>8)b#.#ZUV/ZWRgU7T)@EY0eFdeJZ
ZR=Z=X&QfZJXCMFb/(7/3FKQ:<:.e6Q9D,_K?dP9GT&QU85c.H.VX0<Q7Wdb#H=@
9D)\IV)CCQSbX/O)@0.\d[3/IP)P44N;BI-<[cZ3NDX_0KZOIgKLCK]5.LU?g@H0
;+L&&P-JT[V[/Hf.d&/0;/;@^Q^E9MU2.d85a=,Sb23Q,cW.@f>/;E7f.P=W2)&,
QO>M_OH8HPd2Z>V@9eM=6a-IYB7@Q&+=g\:Mcaa<E4M/E3^&dNV9Tgc5a/b-RLVU
gXb@6eVON]P2Gf[5(GZ,^8aS.,Z.QZ\\a6V+JOc#f<@Vg/WL:02PK.K8TK0PO37]
G]LL1DH^.:Z(3Ug;5;;L<D_R9+X\FWcb6P=2M?ZZcH/]/8LC8RIVX7P.U[(e>gfI
V3\^7VC\,7SI(DbED@75)()7-4Ic.BA_XPdYb]@MNcU_V3.0=2:#fG^SC.@:-+\Q
@bSOe),/,BPEMG3-@>(fbZaEK:?=0X<cX]c&AT27Y8+TR>ZCLY6L=9/PEROMWF3)
Ef:]8WR/@D)8-WWBLOHWB&DOA-,?EL+<OXg/P/c_gJU02?QX7dg\FdS)1e?:M:5O
?5Ac:LV_b?@BQGEgVaEJe,2=M11J[4(D4RCOXOe+^R_3\NU?7TC6<[G[L.4>cUJM
VU88::<NVFK:DdZWfEg.J2737,H)=LR)W(S:eI8R0]EK7T;cO)B^,VZFe,bE7fY1
&7_g2,D6\IGd()EANMV\3WD(QR^?;MW&Bb9?^5#SM)J&-2K-YK_53(+K,gY?,2::
@-af5165@/KBHa0)HY7WEO=B7<\b13bdF@/>^^?T=S]T(+VP+EPD.V-O&\N:&2Q<
[_];:Jb;MZ#cfJ7&KUdc18UG7_6c.dX<D(JQ5-A3c)L^)/>Zf@V&L<:7Q=fS-_e4
;-Of)V,&)]HcEaa0ROM17<Y80F=\]P[57\Q>F^(8:5.[XdC+cXO73FObI1((HEeb
J+3(HT,/KW2OOG;H2Z@H>]LN&d[]O;3d]d)]JZa:MKfNG&PIFAME,93@+8PL^0Yc
D[:.ZQ)6NQf2TNfQe)JD5Ig7Q+Z-F2LI7]WADeOW4\cW^&WL@;A;]EH;XAZFV^.b
K,>-\dC\)]:P\@.?QZ3L=d(X)IY\.8?0D7SQ;H+D>I/Nea62C/?Ze&GSN=A5^@C3
[(NJMZ0LP+RKVU8.&N0F+bB05N(eA-)?SGEdaaL0YK+4?1LUM(0G[(DH_,R=K-;6
+>9KY:T/;F+]R.7g]>@;MM=,;H2=W9=3/=>#0YRa&B0,:GTG+V6;>#G>+(\f5#_4
\?fd6^4+QLEa1//;U>?0HC0[,G1GLD?-92&3J:B,5UH2GF,,?E0#VEE8N[(<FH<<
4FU[<IG+O_BUU2aDN4WK.7&f]\<?BV1K#H+SP<N1??&T>6O1EN.7\BbK+^@cRY1+
HcbC>SJX3)6VJ]ZCQQ9O;I,(4(\T-&=?SS-EVRb&&5QIG,_]f_A(DRKND3#WJ,RT
]G2<@(#K_O;OWOH6NgYE<)6c-)g8@Z1O1+DH8-g:3(AGbOIJdOa>d<cSbBW3F[5a
:IR5MS<Sd5=NV42Wg(/5]6=J7fL#8a6/?aJYLH4\X/N#M4U<;/#0[9IXffLRD:0D
1VP5@d7TY5BYSOBZdF>=VIN[=:OFB<K&#O?T6?@/Fd[aMH&b3_gDXc/bY+LZW^FR
d+Q>T>Ag]VIXXKYK>.1ULH53Ga/HZCVf^TQZLc0UY+JV36KfY200aVdRC19_69EI
<YR-@[5K0gCU<(I+Y@\-7#fDK]BDP&VD]gVWb9dL=@-&.(D?DK077e84:GU&7da)
FET=)>72Cgd91_:?@(S[#eP^,(2I9<BH/-GJ[TMA[\b-C=.;e3eMcR<@,2EUba=.
:-[(A^O_U0MYKD^.9#DR2[R>E&@ecYY@5PJTEY(QFdZP=S[8C#g9gICad\06?_gC
?.[<<C#VGOYb9Wc76IRMaP#4I?Z)1I/aA>f<LN2.DXZb#YR[L0[;8VKA,+=SXWQ)
#E6MKX>=HSP,g@/1L7EVFDQF,9F);2.dP_5b[U0TOdQHYAS<>(QTZ3.K31\fb,=T
ARCU.LGb=19NFcD<fE19/=e=_5)&QS+a#>P@=AddOS7TX5P791>:;Y8@Rb]8gZbM
>B,];R(WB?]Tf]I9@._<AAENYf6dc>ZAaGeMMB[>LW\U-OSabZK=J69[aDV:?cbN
ER9&HF:D-)/HacE]-@H+8=B13XeNYS6-7434+,;L==AA0<4#a?-aRU:LOB1J79UJ
[X8[(::>OEF2:&F/(ZeU3OHNL0HRSAOGE]3MdcJH)MF1Tf6W7)Df.0Wb#dGB<dJ6
SN?-XNag^SN5RZL?T.cA@HD9PV-NWYd3a5.^>9=[dFQR6@gVZ7AO0^OZ8a[QD9+N
6E#=:79EP:3L^J[c[(=-M4.U,0#+JV5fIQ[/bY&).]L?e5Q?H42I\gTIe(1=eF3V
B6,SaMcU.+SfQAcR#+#;RgU9PVF_A2:1<K2#X\TL+U3GAAZ=@T;:VgV]6;\@YV+I
15GV13X\G7UG[EeSdObIN+C.,H^9<.>0;Q3F^.A6UP+WK:gCFAOUOZ2T:U[V4#>F
?N62Q\KDV?+XZ0K9[c.-\M5G[FPCLa(3VB+C^.]8?3Te1=&Y;8I?9=I7f[6N(C;_
LNEe2)gV@_+PQYJ=QS25Ne?SA]G&>HC9&J9eS@5./I28KZ-6CXBT&8T(D4/TC@EV
+UN_eNGX0#+^T8F:4^9S;]>MUSbWE8f]-<C9TG<Og>[,XD]V]N=;U[RW_+5;f988
BK]OL3@G8#27(^ec5B?8#b_I:4+XQRW,#P+1@:MKcMOIE8gSY^UH0QA(^\_2=#6V
]S9e-EIQ8g>\(c#WBL\f_P<FD=MH.U>MBaHG<Ff(B2K\IW:J3-L(@GYFN0(>7#=<
&d::>C:G9]:Ya^\Fc]Y)f4O.XGNOfW?PKfU:276_>][[5HeQ3a_0R1VLKQ7<-_8^
;65(cYSG=4F5S>d5I113WR?U=7&=A:5&2BQ(5b+S.G>9LI1C9WXNSC]>&c[2)U@&
:PIB[d(7&[R>BbP8P1]NBVSZ3->5=#5d\WZO.N=2[X+.d@b.+D7EI))bWObT04>I
g0YHV2?ZD_-2eFD[DNeJ&UY22]:NYc04[@+2+YYAVJ7f^^#c.15)V)\YZb\b.SS5
0UKS-W5G4X@UF-(.8J_M+/d.PQ\]=,S3C4A;BK;PWL8Z9P1AF1A>fX4W6T?DWAH_
O:\fV0/a)C;JAI-IY;eI44TSNgFGS[[2)C,#3[+WD1Y^)O^I]CQLA(9^BP+WbF&:
_]^+Z<^GTW/[SMWU3bQBDK/8f&,N:HT<,NL9Y+aXH)W:H/VY@cC5&IE#Q_7]7,;?
S@gB+>Z#HeZ-42SO9N92#\6?K^,eEf:a>B)f3g>_J@aQN6_[5(8f;28RK#7Q&@Y6
9<b.5<gP+P6EU8b1PYUZ:VBTJZ[UU,P#QbMbgJ.E^E3]NW(QL0e0DHDY+B4R\D[c
YTEd[=:(1A3#<>&1/BLAaL]BU@LeZE5I4Cc#aLJVJECfdP=2CUFM#-6MaW)\P6AU
4L2OGD6@=FeQD8AE-:,B0aOEK-]cNYIG\2I?TY(9CQ]<#LGa+b([N?JQVaA9947I
CZW@=+BPAT3RRN:<L3R++(;P9Z(J#Xgf6C_DSFf8A(01[LH@KKJfVFCYeC5/(M\G
3\:R_FOLSF8-N7G[I6b.X]C>>ULdPc.MDP5aYYB;8Z[DeN3>aMG#]KGacMNV#Y61
^LDGd:B=V158:&_.21]aZ:3?McNTfC/;S]#EIgcTC)=6)7NbcO4C]RVP&YNVH<NV
@LCY0U<2MC-L)fXU0+9R08@-8A]2eMeE#>X7ZXEMg+9-4ASNbW.DRV@?2&W?T678
-V2>.-R3/X9.YG3bPOIL79(&WH[R3IJYY,(aaY5\3@S=YBcaX@:c5,8,-408KF/I
#\YC:A9b^5c=BG]<\N_UGJCUGe0KeD05&/=0X(]27d1I>Y=9.Z6IONJ.VJKaW7_<
Hc]DKE4:_V_Qa,#Z/M0]8eb63?0cOESa;UXW[C.5f=&?B9Z^_#+][OIg3E9O903@
[]>5Qf,PDT61S;:/Ke7XLgWa?d#E]2+;fO+BG0SY+eaZcU1)aG7C[^OQ_813C1C1
,A(-N7&(PU^5M3Db?]YR;>)2L,GcJ:&_[A?7[31?P&aC.+MIBe71+f:][^7JGU@I
<A5.L8LDaEK[T1.WLBVE]IQ22;X1XHQEC3f6?YS^CL,9(OKa\Fe#W3K-\e?e<VIF
eB+/)0(A]b4F(45IYY6]ba1f^L\.2(dc7J0O;4&P^bU)71<CC=KA3[K:ZCff0^ZO
I\6T,@NPPS<8cVLJ<-g@D2A\(;0[70gLeSc+_I&Df4NH,7RNVcQH;;;>)B6R(eZ=
9\KU&?P_fV?16-G&,N(/&ZJ)e/9OXaM_+Ze&Nge,)L)#:&c]HbA-eT7>KPF5OUcU
c8f2@f-f@?8F(3[,)(DSRRUKX84@5Z_-,2aC5:J6D&A5^bLESGF7?:af(Ya8XR2a
0Gc.B?d0ac(P=GNg;=:_2/^TJ366@6,-2KgEN=:77>5..5d59859H,1OU<QcJ9CF
_JgM#CS[7(E62?1ZE#SJJ=U@P6g2DT\aF=Cdec.--OAA]dK,8e6dbe<0bcM5)/7-
41@bV[C0^=g6fW0=E#J8VeOQ[<@.<X.;;>2Vg-V/bV1Of3LH9)[RP\<5QWI0KE#8
Y02g5Z]:5U1P_2__99ZcW)-+QaQ4R-O0.+a-_KRQc1L<)F;LeU.QbW_04ZLGDXEO
d93=aQcc6,LE2(G)HOXTU54BCQ_Z]N0T:VASZ.)(e1]NYIb)[NBJIQ_.)A6MRfO)
>^WT9eL8aJ3[;Cf7?A0O.-J=d[]1eBAbH.X&d-#F8/#(K?G>L_Q,+5U0GV;0OCA8
G\I4P/a&c(X1V38VMZVA7U6ZYD^DFDW<;L273OOMT[d.M^BROP;QPJKWf,S.6f^\
[;:,6OTCSOd.^&]e022N-[OEQ=eC5@3F-?Z8?9B\cfL@:af2^#0I\-&94^;A.M2U
O9/K1JD<SaA.R6Z1F@eZV<EKXeT(?-?#aOedC(-]KP6F.8c:O-0(M8d8_AZ-b0#4
&RN&JO5+[PU\7>4H]_D81,(V<R?b,_45E3S.ISM7M6,?-C>+U^768^2[<N5,;]:D
SCN65D\]&/2af<7@JZORg+fS2YKE-/Y?XMM5QBca)MA47CR(92Rc_S_2@dd7NXT)
ZK<:bA5:)F#bWCXBU+a?=PcE\V5@=F?M]AVUEK=O#bg:^V>AcO?d7-YDC<]?#fT+
K=:aU,M7L,L)aWF)=[BaQ:E@KW&6U2ga8aY^6WI8JFc(5NX^[(a<;+MRIJ9Ha9SE
2.?EJU5@71:WZ;c-S.D6/d7RX3?Ge/S3)+JQW65\U+HN1:3#V_6I<aWXE\?/VR3Q
Dg_A[eeZ3^,R4BN2W2_]//LYCKAP0X6:_[,^7<&R9eMJX^97V]_dS_DdAOLEE9E_
KFXa\2O)78dY(K;)K#WffW+B_AV98)?<F3WFD=+0GG1WE_d-:3<X9d^NCRLeJAb.
GVMLd0NaOJYf6LLR;]R.feaWEQ:NL-cFRT0OgE;KbbM\R//7J.P>0<QVP=4e;C_G
P]PT>bT[#)5]D0+c#0N[VT_IHR#[:9#,L4Y&eZKgA7TXOE::.WYgI]YF?;.#9:2a
&YPf.e\X?g;91&de(&<f=e6f#6dLC4^6;74]>NIOV;3L2OOBc,\:LY8,T/3PK-Ka
=5D89SIMEP13HOe]MG49f.8YL^[.X#N,H4b76[UU#@GU8CMIa?<2B,S25\U:VcB>
?:LW3NNM8f6c-3?==e^X0c)Sc<1(4Pa=A.BILO?9\DB#=TfUQ6PPZRX6_43FR2Lc
&8Y3G(42MTWJUH;QMIU[3R<K+N7H>[-G3.0WK/<[N<(3\NVeP?RDJeP>\/:Ve1L-
DY?+HAD/9?PEA^31:Q@O4fG<G.CU)MKF1#Z)d+gHSAXafW0\=g;T]S85B1]A#;4U
Ob90LCAMA3[IP[C&UI@V8cX&U@\U)B;OeU(L7YP4b5+ZXXg\6O[Y:^8.+H3\c-U)
Qg6).^fKgQBb:EENJddZbABbEBaQCTgX<DZ_71AY2[bGU-d4Rcf[HVM1\3/bbWdC
LH<d#Z43<67e]g&=OU&KQ&R_&BL>KD4)6.4RX]4@-HJ^.Ea1&=QAd5WgU,=C3;V4
6S@M1(.\,2ZB<#2c(3XZIKLB&^5b&3Ue=WFeE9?gF_MEJ;_dB^gG1;cB<eTP\1M6
ccVDE7/L^55<#e^2YeOG>[DPe,3\>]&9C.7&M0^J<8CVY_+&K](66FQ>45G7d4S1
TSNeT/,IC)9BU&#]KV:/DT>O7A.N<Uf-^^BL)G[b,R[+54,&&a0\fO7FZ(-3OU:L
eUeXICb)2\/0SN5@T>]FQf;bKLOfE9<&EA0_ddX)JVK98Q(HLXTJ4S>H=,+9[S@4
C&FRW^b5B9e7UDA[G78,]?HV8>HXJQ(#40[/;/\gYGcK57&&X<V(43Y3)f0K,\>&
Tf3d137=>/Q2E\^JRMT>c0NgVaS_KQ.AVB]MM.a.487SRC@9LB.\;)(3\T<^-63I
Wf\+8^Wg4TadMJ\05#J0ES/NL63f/<@;CI<Fe^AGVeB<]?-^.77ST;<QJ;gG(^OT
NQ4[EcH:3bc26=;dN(-7AW(U\8E<ZAf3&,cK&PH.AHcB:60)LWN.3EI:6+<KO6_W
[>(@2D=AN5fO(a&N?NB2.]:A2#Jc;(;6C;UREBUcTg0X94B]B+733NLaZ=U,Q>Kb
]DMPdT,Jd67#.cK+/.8U@>7K0(<GFaFI0bf846]:D2Ica)3FJR>8VW1^[;,@M1H@
TYWRadNVUOUfYeJL3TD)0Y9A)a;HeMB>YCZ(H)9A1Uc8271?P\)&g-O^<@7N@/Z+
ISDa]=N\W)H/[;B_Be-E]]9KCE4[\Ha-(Sf6.:M<G@TKdKc]Q#4]9)&<KGBQ1J_@
5A\dTG+?cAXVX>EeL++-_CCXUa,Q;Ob)F51)72+[[]I\=T5L@U/Q8>F=C_eRA/[&
OHJX03KX@-(5GP4Od73NQM(QQ98/D4LP,+;_Z?,]AcGC=E2X)^VB6McB4f]9BJAI
I<_MWXfG39^?VFX7G240W@>S=>b;e^>BgUc^.[/Z]X3_\\])H,++VgEB:Dda@Z7?
Ig-XX>\J]^d(S[6]E89-58QQ7\@=^bcP72Y=M(P?KET]<C5NfgK+-ca._TJQJA;D
DX1<4XZFJH,X4P.<&BLV81#1V>V8IbC,D1;FV:HCDI_ZWA-CfOCN0-<XNbH&D-[I
<9C#N^F&5O98LM>gO6Re);;\21M_-AX;;ELP\YF8fP)2Y9Ceab@(=@_@-=C96P@Q
/8Y<b:)2JT\L;CXC14_ad,O2PX7Jaa6(<39<SKC2g5f5MIXaB++\9^:K_BP/D\,[
8G7J6<0.-CJ9&5&@?V>DV1@U?,;0?.#RIW92dCKQDaDD#aWY)E9X^3-.Zb;+R])c
GcYS^]aRdLMBfM(4Z?1:PXG.I[fC?9D#3)O)9900_&B1F>(0/;@SJ&3>Y1)R\R+,
1DI]_V>dRJV]=@L)IBV#O#e;X^d=;\R-],L1b=fP):f[2.IUMZd3KI7S<d\1Y<LD
@H:\f,b)O+aRA[G^<dF[RXY>aM3&-,V(E=0b4aXZ(?AI7/MgK/\>P[^,X,19=TGf
FfeB(M4XP\7Q8.IIc&Mca.&TUQP;d,\\BW_5[3,gAR&A)\_?<^UH@;YHH0G1:e_D
01&3CB;fM?4NVRO(,b-36^XWMH^dS9O5_C_[WbPFbY6BfRJK+^OAT]0MR)48Q#SV
NHTJYAV@Y4)]:_LNB-HT0G?U>7Q+e#Dd&O9a&HF=5L2)ee&<YZ65JRb5>d+4XE+-
)42DZ[-4/=>gZLL/4/@=cf8X#A3d[23N,J)1&[90448-Z?cCFS.ZW\C0Qe586&d&
/OZ>\(#8JU[(WMD#/HPd=4DX4ISeAER:ZUa&Jf(L>S8AVB8GX@&QHFY#e#3a<WT<
YcMCX+U,K?HO>_Q3X)6TNDO9_JR>cBYa>7P\1M.e(HB_BYNL#T@/:gdEfDeS#f<#
:_WI4fa=:.M.3XD1eFH@PG1B?F[@>fXDJ]-HCS+(4,&)(W.1RHEZ;+/AOJM\-FT7
L6\_#O/[c/Z)0?W_6W5(A3CLJX4N(&52?bd)/I>9g5UCgKS1a_Z<MbWWMRT8F33?
-Z:[+4#+TL)BG&I@VJ9A@::@.D5a.2I3DG.KMf#f6T16&0^(TL96S(b0#N<B-b<4
@RAc8A&8KZT/4:(G:@P(:25:R<#g25f?+0:8N@&#R64<7G21G?NMF_+NA=QIB1&E
.)S>e2DS;R]dbZ+U80Q4I1BM.YAe_KSaee^?&MFP=L4/2^gMb>FJ3JUABE66S2;5
?[B>(Z:DaG:1M=GVVG1)S8g[&Y@AH)D,BV8(8<#>]IfeH7;@7B]/&M?O@:GR<JS4
M11/)JaV>)E[-@&Q=cD1Zf6)dQ:F<;XRHACG;V,I(0U9(1-()NZ<a8<4NaY([F))
GVR?I:[_8,0^:L;[<)8/^R&IfW<+]T+\GM0O^\D@&PR,Q4a^Z>(ELYN_GRf[:M?(
#bDEF&\?7,(CWG+1-;K4MTb14_gC92C902K1X?8E;RGd>K5XW^8PI/IG#6VVg&MH
7@fe\)VHAGCB&O;(f11U/>^@LdSKcJ;6K>+_[X5BCfTYcL^F7WTc^LPDY[TQEaG@
KB.H^L0aa(,KC5MK#_d3AJDgIcA1470O0CR<D(L/LJ=2Sc#Mdb<M,M<1bKf+?Hd\
QRXcb[+J:IS/NJ2@DP\/1V3W9=[5RW/a<.?O_^.#I#[Vc\LaJ0#12DI?(TZDd;dQ
#(RL49DB7YZ>g-5E3-EKAHW2++,1EK)NOL^Y_F,RNc9dB#]8LL+X4)5d_>9]A/O>
NYFK?,KYS(7:6-?4JcQKJS>K01(/;L=+66aM^2>P:4=4g&6=GZFe-GS-(.gJOK2D
/UR1F=b^0a+Y9-7YgD85XOgPKO]VGA4;LcJJ-a9D:AF18OZa9@e,AHMTNff?,:?U
#Ma12[=89Y&:7[e^<53PQ)DMYaZR62HC)fa??F\4X7cPW<,DFH92OcgL;gAVO>XR
G;_1XT=:^Z\gEP<HcA-O_Q37&fA<F6V<:GOW1)Y:[gL>Cc7))U)7B(;JRS?T(]2C
]egTLQe)&23G]+C^L2FTPRL)TcR,Lgec,&;/GI=Hf2QPW4W/4;WJ(TbE2DEP^0@9
5J3A]0TR93PdZ??CL27GH:ZP@14-2S3QD0b(_QQVY&1JS.<@QPSZ(c=,ZHNg2)E=
/6Taf7TAF#:&UcG>Z#BfLSS#\fKH/Fd>Ze(.3:H>R31VHK)6ee_a@G]TFTCW@Q)<
2KUX72_gJWN0\ZN^/6(d>J1B8ME<Sd:C?dOG_;@]W<>0_Y=H3&@:[R_B/\RZDITO
^IQ<bJZ#Y+ab\Pc=Kg_+XJ_Lb6I70\(+CTXNCQF)@BELB(4WY(eC65_ZF,V,JR1?
\U#@:c1O_81e[C.U28V-MFOR;PRV:_S?]D#(+b/GKC6]a3L#L\\70=3#DBdE5>Q3
HP/+/BJMN2TXZ?-Y,eS3O3;9<Rd8HVLN\b_0Q?Y;-U//aLQafgG53(0MO+&CA^S#
YVfG),?4^^EGRL\<]Z5D/9N[RG)P1_dL);84gg+:?G][8DPTICS&WZ091M(<[308
cDY#<7W\(84T7a<E?W3=;cd5;gNEc,++8R-MA/V-8:P0XX6XbfZO4I+M+C/@SHK;
+)+^>5)##1XBD8\I::OQd6U?D9\ECU/R>OLb<Z=H/GJ/QgTe\.]7efPX#37@Ae=)
-cSaV8@^P778QeL=W)-Bg&M.L@EcU;UFfYE&//@J<=]b].4_7-3KJ\;8BR_#U]ZB
LT(O)L\VKBM^HYfH1X<MGHY=2^G+-UbSQ7MG@g_Ke\8e)f0[H&g^1NBMfgLP=4;b
9YXI1742a]C##f+QF:Ya@BV2IH8+1BcN#=NN#?^H^--:?Y[Z=L]TT4<?gdLN5](I
,ITGVV2\_>fBNT&&U<[Aa\^MAGQO5675XJN[N4d(T?I-B5>+W#DA\K\_8X/@0g:U
)K]g]N8+J^?ZTREa)/&7^/[Q^\BQQP8ETLUZ/7Ce_LC2-+&]YBCJ2,)0LP5a/YJO
V#4..,6K[aCF=,.>7I,IQG5Y<52H=)c.-@8PGC.SCC8MDR0-XgF_GS8<Xcd@5HM=
D,A?Me09f0;:>J+:L@Iaa9Ze6HK+]P?)(.==(-OI5HJ-1E\eFGTE102^X._XQgJJ
B/^?e<O>F@BF\@6/SS8-JRJ;5a?Y=)cKK;<A?d<T1W-0LB\K<0Z92,H8:^LJI^Pg
e,?0<d7T.-P?5XSfNX\E=,/8,&6\L/d)E##5D,^KU)(-E.?\UH(A3##c)8:<OUSf
FbPe#JYH:WN4VZU\2IFde:<X4G#dCFFQYO;3NN6b9XB=6A<F.JJ]J,R.5-C54JPM
)<E-LUMHWPKEBXB/TC5O4J-Of48DC/S.<9+;V@RW>Y7De_9V5TAH/)cfcUK17G)B
H1@/RNL_+1Z+E:8WD:T)LQ)5F.<\\JY0:IfMYPIPM4M\W<Q4W^EFAL82S(Y7eZ&B
KX8?Vf[IePTZe.4<=./6\0a6S(.^JVX#[dIbQ<JTOQ[4O-&ZQ1@-0g,N1WV>TB(2
-^K]e@7UY[4?AYR.&,.dYMIY:R6@=-^#3E,0?/fe,>VBffPc9CUGWNXY5@e62+/O
>X7UIP5F,R_b/=?&1VB<eU_HXBV1C#>fHG<9S91RGO<C4A)@M?\:DYcIfU3_V]1A
gFL[4D0dL6N19HT94:JF,O:TL2T?dM6N6R&B,baPdZgd]&<.,.WQ)[Ydb3^fLM>H
>e,@?XQB]\O:[[71;U[[NZH4LA6>:,U]5TZ:];cRbFZ-,Y0b@M6K@W6_1HE2@Mg/
+]:&#WD5R1HE8I@eB]6L2g[a1>_X:QN+]a<R?&f2X](4Y<Hb73ag3:G-FMAQ/ID3
e+fO]dOM<(LJ6T8AbdX?d.>-A#W/8D(]HE@IR&_XA:6<DV2VJZc3210#a2OT#a5S
bVOH?eaBc;U\#bLN<1\5d8V^-)W-=Y1&IREJYgD4@?Kc=MfJ#DMT3U8;\_?3(,#V
2#/X7^(>FbVKB^0-EJU-;XMZUQCWE,Xaa@_4P^WEIe3ZNMd>)]=Y,4N,/S<2O&49
0M3BKSQ.f0Q81QbYP3W=R(dUFBC:-dA;R.SE0MP[1b_JJE6[+BB0g9=WF2A_++ZZ
?DDMcI0J.,ZWC9bJR9]XfM>\TG5=3R/55NeTDK2;1<<,N.8,KZ.JIR>Te?X0V/7]
>)gGHMG,+[WU7EE@XG>X56Of?X1g>-ZL.gI^e?<Sc[#ZeA[\_e+6X[@OABV-?XLM
C2P7FBK/_C)faUNF9L8(<)CVe/I)YW=2:Z6Z724]BC#45>F3;DKBP1+T1-JFCTZf
Jc2eA,1P:3NM&89Re7-^=O?,0efDZ(M.(JLN5&GN-=KZ/B2Y7><\)]L.@5../9dY
eDgYXW\VBN,@D^3OZ;.N@N(+/<Q\4&^[Z\6M_[U-9>E<6?;&]6ZM5KH3;5G0B8d\
J/3<C9M,NA50B9N,:9K66T6&/],73P4^D5_J85L>XPU@:(9[V-4UCZUQf+-&=b1g
>\#=PG15OI3&SH04c]fUT6(NfA&NV,34(f5c&PB3GY]1Qd+5bBSC,CeQXc.+D(.F
)eS,Z_/CK8G9[;&eJ[=,RbF/]KUNYF?>X[8b-3a#<MZ5H7ODB3\)g-CN&MROOTId
&Z-LF19>A^B<G27T>AR+?0Ke5]C[R\X)EcXW@^6NaT\\LgT;9\&TBe,E89H>VBF@
e8LJN8Ld.X/TSR41TH1Vg9]gAU?.13]:OPO-YI\IH/7R,)&I<J@A)E]R-/&BUK(2
ZR9(K_<<:&1R^1a@.c,-&;,.BP3cTC,E2Z0_C:_>PB]8;#.XC]NU]=XAeA]dRR5M
8TA,aGg??4a(/KLX?&TAe#;WZ<a5\EXH8TINeJ9UTHfQ)_E3?2B;9=3?,a/:#-I-
-[,T95<.9I7@4)&VQK4H)M@aITI[a1UEP,Q&XQHDKD1GgR&fM9.V=a=T=GGB]?38
4[;X?eXH8?RIf9/))VdE=(Gb/dK1WT1Bd6KH3BaCSd6L?ee0OT2O+&gS5:Qde:FI
HR=(GM&/,cBS8fW3Pec)TCN8O^^=>c(e00(+<2\3YKR?6aV\/3d7/CY&2g(9,^ZS
?-C@[[\eZ21#D:G+S8^QeEX>YI-\)BF<>T]Jd2XR;\82;TFWTaCOGWf5d#M8P9PW
]&gb8TMSQUV;fDDQ+gVMT]VGcRd?#=1FAbb1YPcT+3g568,A\OOF9CGZ>KV]^A<T
O/:DFWZLU=D4M_d0ZN6#WN=Uf52(1N_+:BN.DZ<[;X2f8H838M[=5=AH7#PBK6<B
]VAO@Oa2[_U,GLPUV8eab^4&VNP\c?G\gD__g>&f6H>)>3U8e).F1-DW#O-X8TZ6
YQ-ZOS\BT0&a7^.NR++X79@YP2Y>2Q)<RQBB5A?Ub<bZFFYNg231IMNP=A9)EG3&
dTMM+QV\PQHa+$
`endprotected
    
`protected
\5.Y3?SLLf@VR9Zdf1I,D]Y7>F/U=(/@36fNbR4JM67f(;58ea4T1)I5^[SUF_GG
O.CAC)HLU\/B5>GC\[2_#a@66BIZ.cX=;$
`endprotected
    
//vcs_vip_protect
`protected
W2AJ[KE6_OTR_W\]R9&&U689/ECIR_:&Q+-T-Yd497SG0UK#XAfe((R+@)c-G&1=
EYZ<IN-W+G^HgWG<9?ZJXMb,5@[0-LSe+3#L246[:d=W??2G6C(/&]P00cIAN-<)
WDfW&05)E1/A[,8d:AM#_4/KM8+OB\U?3;T42H;<C0Ha(@C.fN]g678dO&HI@@)3
b+?)M10:gaeWRH<.43(^[GN,<_Ee9)QK>Ze#(QZPK2)NR6Y^^EAc6=9+:N^CO/N6
WF-P8WCLKf_2:dBCHV+aYbGdN2MW<+R>+QETX9-0(^:Ef.YJCXe_7-dfXMY1[DDO
a>#_b:S>:+3]2[gU-QH3AI-,<7VF[EVdaL57ZcX_KI@:9RVHW09T7HT[P0VK:RaU
,F3^KCBSg2B.ge)eU?[L70bN[b3.=]I+D1^3<+37V_5^&/)/GH.M.gHB60(\@PAF
>,9WW#9\Q^-5KE#]PG^LK>7G\Qe7#+Ee6G.^]KQ&D.7DZF+9,L83(>)eW&@-a#ef
]F&&KFa>]/=_]JeC6L6/V78\_O:P7g6UG\86>QN4##KP,Q&W^.e86=&R9++0\bGP
c2KCe.=1QZTD=+&Q<g6NSQOEG0AIVXA>\F?ST#/1B:g@cgH^C.#HbRNNA#Y?0g9F
Z&EOC7BZP6W_:E1N9<-8=-KKKRSED,GGZ6:\Z>;/bD<:d9Y\d6METcRHID(H(b[R
H(Z5>1f^+Z./FZFHH0D0NU=YJRLf&]OLK@-f-\\_f-6R9R[T[@gE[[H<5F]Y-1b[
W4QeOD]XgP@YXTOB=.;_aR9G\aYJVaHAX];H7G7X5IOCT,V^B[PK1L37#N5AMJ]M
IRQ-K#5a09>JT114E1NI8=[FN7AB;0c#SY8bRIU,IA/C-D:<ge7L8b;MC1c-A;:1
IDXCQS.Y7I,BZb_8PB2D0Z^g1>=2I;I+dV&OScIa--e_8;ZI].8[J_1a2eJ&BDZ=
Y=;d&6#LcZ_61E,S/_1ZS]bCRYOg[WC<=U;#f1I]PdA9\>@?(Z]W9P^=NK;P_1FH
0JGc]NIMF^D,U[:]6D@\9dcgS<f5FRFH)?#N9?(RU[&X&e[A>]YV84IX^?CWd\:8
9-[?X:6fDJcc:?+XFFP.9K71/#(I=#MY@b5.BcHV7A8;fRR13Y#>?,6&9T(J3==3
-ZHGeXE0Q+]G9\T(D5^,\Z9T&)BRS/U8BMM83Z.BYPf:T4Y+&;-P0-QKG=dVAf:X
\TW.aPCD-,81A6<Vf^/Zb0WD;1Q#:>@ZU:F&UKbRMQAC;NHLcA_&1fc8-4#F8f6&
-<#FTH]&O\aaf=dKY,1<<R]3efSQd>S:#W1]R0FWEKLJf\_c+BBbKcN1ATWSX_?+
X)?)EHLTX4HLTQ/Ef)H9BY]b5_KKBgb4#:FUNZNbI<9L6,e(=a4-cTQA>2.,J#C:
&AE&O>[R-8&8(L9KC.Y^#/<D1NBWcL9]/P24]]<D:ANbA9UdECLY3=37[>dAbca1
G9_XXJ&GaQCNC.Z&)aJQKEZbAE[B@@Ae@aI=7cOYCTW[9>)RF=\6+&4Z9g+F=W2b
T[RaW=(GAUVgX@7986JKCMDUV,dCO\5S:E8A4/N4)Y.\FWJ]g>Q)0DVZcO4-V7fc
FG?bD9;U4U+2W6>Y[P,TO>/>9E/\_NWAOeRL1ZPC?,Q_5H7c#L35]Z(@_UfdZX5f
A)[W#Z+<TaNIc6YASAWIK:@4A=-DMZeC/Q&cECZ+<CJD#6+V:28ab@WLGHc&E>UN
UT]M1A.\^<L?D4WY?&N09cg7>Af5XZ_IJg;RR=O1N]=RbaY(C^QEdC?YTf7ZD3^T
L8C9CMfUPHR.,NH/VD;U9a4<+eU]FEFE=D.#,AK3@SW@Q17@,ag8b<S]BQRa</cG
\D.0#O,M?K/,;S\)Y\Cd]Vc[#YPP[d3521IKRb(dB3.QKPE04_./Y;g<Y>gRTZYE
TK>\:BU3<#WaF@;8__]YaBeT)N^5A)6S/3)b\/-->XPQF/+U^8Sd5<&4AUJ5:X)<
4fIDRNI@(&NHJUK8cMTXU(1E>Q096<G-a5,Q(/2./5(-FWW[e3Z1F;a3HTUP0G34
-)YK7FLLcSZ4,Q9AHBY2A,g9VQU+ECgU]O5RfB6HJ<V>D4OVA?U<6;UMHUP7.JOH
=4:+MG#R2QCSJN.N[ea2X/a[\<PA5>CQ&?a?;XF>2+D;F8ZY4(,\eX+/dX21YLYc
H9<VAIR#6)aAM<IJAYQb6^@N9RJ:A,a<X]J=^1f#@0DWYbaKW<1BGV5B(OB-#XYO
/@TA)VLV:a5>)^N6H(c)/BK.4b1ILZ:Q,.KEAA4=VWg6C>Y6_A5c/P.);WaH,f0W
GGPVL/@)f;X_K1bVDPG[a\NT0WM.e_HQ^)1R\ND&J\8MJ/_P1/Zg3e:9CT4Y]2^C
7.MSRdBe^FOeMLeR^+?Tg;T.g@?=43GYDM3S<[bVAWD.P25DB_KU&@UNAK37I-RC
O7/NfO\[PF:]d=5eLHLNODeE#T#daaMYfXCebe)_9@WAJBD9BScH/2?#b77aKg:/
:P#6(01g[\\3[A=]OeE72@JfU5Z)Pg.8K4D_.VZ_fd2KDL)VT?d2K+YGQ\]CfAaL
R<g7PX0D56bI2-##Y?5X\0bU0(g=XDY-S9-P^3^];OLaPR5=]acKJ/CZ<\#B8=aS
d6\2>c+Fe,V>9b#K)8QR>?DM64E1&715g4Le71GAT9<FBJ>X+A+FM(+0_deRADG\
C^4DGeeaWY3c91dEV3Af;P\9-3(Y;\gc56VdJQNd@[)@B2QYa5]X[<&6eTR<.+0g
NU9>;&K+=+,?83Q>_?6W;7)@EC2I6U?JZGPU(;:NJMeM@YD^FF1XCIBA7f/VT,DV
T@eN;CQXYLDcLOP^dH@_&XT64_QHZZg#0=DUZ5>-TLeBOP;>M^,++EgLWg4bPF8Y
7&4)EDfK\_=#]e/&NPW\eW)#&2T>bA2ILSCM>D&S>K)Ka;_>45)7HL5De&3@Ce5[
d?M+Z(7II/TK_[gYJ@Q3&1B[2bZ<?50Ld(-DZWHgM&[aRAVLMg]OdN_N^ee<D-,-
-JT80\#If)J=U>eX47CA40LcP9Ye?dW)gH>X@O(R(_OgUd8]RS0HGUEK8RZ[=2>D
/ecGD?@dFM,[,I?T)f@3J9+L_R+C@[0G&?g4/Z4:<+N-OR50^[5I_53NOGOE)f)K
(f^N4;>W&^9F)]8PIPQR.^ZKe:Q6@+)F6d=FP6,)Q/AHGCO^4V1NU-9D[N/:G9g<
ceLM17<G)SU3YZ,9AU#ZWV-T_5L#49eGf.[E._[M=6L7&+IDOQ;0WY&3G<UT=4=R
dW[L&cTZX[aaXS6NA2?)<B+C@c+:KT1L,PgEW=-_6#M)X39E6+bOU6C+XMN,&_C/
WYgSD(71GW\E52+[SgRb9UJN\SY>Q2aY5(bQQ\EQKYKZE8T4+Ue7Je61f_(Nfd/-
bO_YYSd6M4)32:HK:54Q4L_K^G3[B-<8a-Rb5_:#@2Y@FBM9[86C.<Ee.PXg9X-c
7)\O.IDc/C8T.Z#fG9J[[f&.f#3NZ1Gb09e>-F:]Kb3b-NJ.AeSU_T^7<HZ8KeJ0
M@fEK0CFIA/51&;[/9881_9dJ:6ACCV5YSA5.^e@W<8cIL4+A+#^(D@\7C+6S#1)
8Z9Z\WI1I#bKIZVg[f\9P[O_<W&Z.c]PH+f\&)JCdc)&:>G@6Q2U[[H/6(,ZEV/N
>TT:21-9<I=YGJ6a/M1f]=g\X1:ZLYWZ#b]b&Bd=U?]d2^gF7J34,f(F7/[;>67H
Hb2#.g8,>[^b&Y6>IEgKH.[RQaQ+HHA2M@YUH_O\IK\9?NUV=f\aRJBF5>&YZ_TQ
Cg\JJIDNCH&E&3ACOG_8PDC]gZ/CXJbP>b&8MXf6=7P#,-.d?V<OaaV,XCG^;>\#
YB_LAG3E?=6329N0DK,T.ZWKU9b39T:\QO#<eJ_fX31@4-;_)78T0<+]?X(T@:X.
fPN-?I#AVS41S:ZgEBP@M13c62.<a=,.Za0)\CO3@G]R37+@A@IWC6>fZQXQ,UUC
<)LA(^Ngf&Q=W>7M34DJNL=8;.7/;0^N)LM<C;_G&^e-,V.:)J9MT+Q.9GC+5>O3
A(Y2O(1/<37AU);Z]I^6L5a7>GJ_O#VD]c5@^@R.QIg2U5Z-HV2<^O2OI^Sf3JHS
/-5b4;9LA)DZ@4Xc;fcDN(0S<g=2<.P8W_bcJ&\DWe91?H/TWQI&+Bd^AI<;NBQ\
-f?HS2A@:SQM[TT)d1JNW4HTQd_K<c->ZZPg7^=K,?/:I+8.V8MHTf0.5ACSf0/J
KTZ4^<8V9I4.;@2@1S,M6e89LV&U(5UK-5bYId[Z/PY\[c&<8\E>F^DGM+0:95TJ
gSRb0AVgX\bZZ:3VEP<;Be[KWUY5JFaH::MCQ&J\<V>1AHVe^>0eDGN^6?fL6OKP
:?,V.7VVNUP()OA1126C;)NR<cc[N+Nf?5KWd7]MK@ZA@FTJ#2;#b0#8LV1I+8EU
:YFCQU1Q;II0a;<_6)U@Wc5DDYRBT7ZdA;8K3[GKA4(a:_77_@fZB.3U@^SWXN<C
GJ24&]UJYN,1^f^gIC[)YN0L?6OLV2E_>@?R1Lf64fAbXg,992;-g]6PG_L6APD9
P0:dW#^DcE[(><TH:^STN1(J;3@XEKbQaTDCOLP04#(43bLWOHEd[c0fe:^F8@M(
7-1IUbJ)KN=1QQP>g/,3EOM.K?Y0bH+818B0?P/>[=L8=0?LI)1.;R)XJQg+?UQB
(S;ZQbJLW/3UKf3R:8UH_Afbd_-#0#AT4SIg+FZ:O6ENW<BWGgTG6a(H@(>FCed=
0,/gECeE]D:g\1GNOK0UMZKcd>3^8E+6\a09-??@fO)KITDWe2Z3RK#GRf)@cJ;a
G]\>:L.[cIb3)KP.F1.8Q/,T_)Z6:;&,gZ_:=AeRgS=U#_/IOQe5>94R0M9dTN7g
CBd-1AI-@ZT1;Q&;^F^SUU>?AWVPd6XLM,?&O9ERN+0<9&:)e#P)D&WT](XTR&+2
PT/(V#TcFMR:-0,T\(PW8=Hd7Ig[,dEUG#N&Y)fHM_<-9X260K08gc@86ZgSaJ+I
VE^7#W_\gAIM+.KNTQ-PFO(c+U#=g@=S6(#]=6_gD3R(CXG(]Y./g#0D5V\R>J.W
[15&4\e];)@4)U/D0D+V02Q?/Mg+U=K?Fc\L8-2^e>aO(+D+\&O2X3]79dXRQRR-
5S6&NP5YVYcFQD.^W6/[A&a5(+GUH^.Z?LGR@Pe4f3gT;=OFUIRG+cZ^[5Yf]IT]
f_22cI]IMDMH.MVBb7&MfND2fF;2]OWJ]]1&LVb0H6I,&>/^CZg@I=;0[)I7G+UP
/fSaIPScNVKG38I,YO?&(#d&(HUEOOM64.P76=[YfVH@0,F(Te-B34N4_7[57X).
1G>L-D26JDZL/.[OY_CH/3QXXF+4;ZXXWPc6?#N,fYXa4A9cUaGX35M2gRI/&6DU
ebH:K@SDce?#J4@IG[F;FXbb_[U1NH.)f=[CWe:,GYd3<>@H-B;.gZU#OQ1c;:-R
:V)NK@S4B9O(VJ(HbAG^^)XC,_M:>e_0?]bdgZ/c0BO=3;M2Y.XVbQTXRSF;].N)
W[5L0[L=M417@CU9LJcRK[Y?GIL&1QM+G8e.W&SO07Z-T:D8^0?7.>..Z0&BB,D&
Ad#-CMSB)9.fUUZL=^9dQT/N,bFgK\e9=X&WK70IZc]/@N_ZR=L[)YK=.,;f3/9)
;_A0LD5-J#E@Gb;&?>L5]4]:X[B\R/[CT#NG.GSZXX,&.M^gV6],DQHZNcS^4:@V
7WWCcIN)0S+[?F1=-)Fg\7KdB1A^aDKe]M99ebHbc&=#aS0[#73_>g?UGX@=5Y.f
V,=&U/_EPCA;e91?M@gRW<c-P@X;ZRd;C)#9L5:A0&N67#L\SP(fY,RA1A5gd]W7
6EYRY>?77O#ba=P9,:NO;27U3F7C/.6ZEBR_-/a9D[QLR>X;&2Q^_Z+UB#VabF99
^aT@R5D\,F<5B?:<e6NLWC</KH?()gWZ#XI^+#:&dL6=]FMQYF6V(JP]#a6DfSeA
FC19F]2-&;aD2ZVAgBM8F-4PCFI(.I^.0gG9BeJK;\^EU5G)0T8c;F&P3#[<W#)5
8[+QM-@e6V^;F:I(42B42T</bR@6]YVc5]K)L1g)YJ3g/^g(P+.T.JGIO2JZ9&Q^
QX-UZ(NZ6X-CZMILBgG1R-/&?I5<FW(<3ZQLVZIFZ_1@a0KaTN;26HA)PZ6+3eFU
-FNQ0&YbA^f=f&P5Nbb&4UTM76gc^K?@eE=D/A:ILA+c-\#gGOdB=K.4,Z.RWK&5
_M^3)g=AM_S.@eIZg(RdDTTS<VD8C..NGPNTIT<S.G4A74:EM&1\G/N(e>7UKE0G
PAE@:(USF^@,g9M&<^\ZAV^1dGU\Q58=VIYR@]EH?]^]VTT6.A)dBBWLg;+cE&F3
QGg8g68;64.4c;E#,T[d_V;\+[Vd7\:S\ES09eJRdSRH:JJ(;/I4HM3QPS4BBca/
d0\\NC?0CZ89_14b]@V2@.T4d8KD27E<(DSFDQHWaYV)GZ.XB/aNfHAL5?6&@EC]
Q0Q;TJ3ZFdWA@)^;8@C-CYC3PJ?cN/QM/)gg7Zg940-c+JE5PQP^+Y.6aNYeV^#\
bC.F5V.-\b;CK.5VQ,#9RUQfI>10b0#W&e\b30GfYE>b976\DbO):(]QXf-V_B;Q
B81WK(E8&9eHYLJc:R+YF8L-#2a<:+H4VCCg+gF[\g1,F>;FEZOU9H@MaBI<gIC>
GX2bA@?7fdHP<)CJXdb.>\P2d-K_Xd=A++WXf/\#\VH\]Ac@DZ8HRVD38B:Od\/_
H7dfLN4Z@g[B]TB9Q8f/).O/]<Dc0NN/0E^2]8Ue2V0RQI\U0L;#V#g<I]K/11-e
JO)F&0?K&K<#OVgZLg50,aR49,e2W..?F8)f7WRGTL)e2(7Z)#4@9?5_V@FIXfaD
Y60fPG;U@=ZI[8[]BI.YS3U:I8cK<,MQfS?;LTE?gF9Wb\9=Jc0PL[>G-OUGI]EM
B7H=aMaT\,?I9bUcTQMWH64Lg\<(\;=I:bUbbPYS:eA>E@6LT8/+J]Y@Ta5fQEL,
bR\XaODa>:ED<]LLUYMJ(-1W^#I;f/EC)HI)B1Z^UK<94P0XGL\CLCOYY-6D=EPX
H42?V,?;/#fTDUWJb<4)\M3<.>KV^Lf4./TTZ&RUNQ2/UDF_Z-MDA4B26NR(^/IG
fAY6Y[EN[AKMXK84aPA/F)R.U,5]NTC4F=+#:>(WN][#VBI8ENOcG,BeeT0-QdJC
L6PWe\^Y.dCEWA=P_@/B#X[^HV&I0QSd6)YJD?Gb+KP_I=FA2BLA9.&I8.74HJDN
I#,=;2..YJHJ57X&3]BUWPTg>fO+?WHZ-Yf86eBT_-0O9S#S)F,U+,Pd1LbJ^aW/
>g5Tgb\&&>U@^fZS;dDMBEEd.LS=3:f.W[^/D7N,TJW;d+5P7bbKH;]=72e.9;;,
/f>BBCCRSWUZH.HO9b8X#SRO[_>eA5?EI4>=G4f?c^\BbO0>PML@)WTB]9cd^aWa
EVS2d2(EY_LOQ@H_eWG9#-L(-7F6@F4BbP+7LI[#Kc][@N8[=\2bV@M6,[M<g1O_
NC3WQPM4ITZ69[^P/.0D0U/B<+&.9?Fe9d(4XeUU/AY>H)\-LH280-d1I:^ga;A@
Y3[^ObPZRbT:B8IYL@eHdfgCO@+^C8_I91IQ.20LO:^:cI\LO9fBGLTVdCf@/QSg
Zd+-YA0;OF.YFZX/;=e&D(NSQVI[#_UD52&].1(2>S0E3I^/0WK(GTY_45&OYYPE
BfBU)BTLU-Y_R5#,[NC1dR[&a<JG+MCBc+>-5+HLUNRg#<7P4]N[5S-XWL]]Ac]3
O\AQ,VFcN:6QL;6<7WGggCXEa(57fZbS=\#2R-QX:3.N_&7A&X#Y[1caBY+:+3Q?
0XCRD+dgL:\a8?JG7Od9Xb_6.F<1>L2Q7@=^1TK+Xbd=2DJG:&0NfK.?9+\N_1_L
c#V&UcJ^4)S//IN@Vf#])&9FbDD1^.8@0Z&7Xf&Q4;feE]\M5aLY^,2cQJNK451/
NI1;S(A10V^_K9/;f_=-OP53-N@JI2fd:W]&e2@02:Q+;4N(QQOU1N@+dRJC<RY8
9OM45X\bT,1f>gML^Tg8(Z4#b>Z)\dS;N@.f8BBUfDM<5E3FQH<4b^_K+CSY[Q2Q
OJcA<L/UMT;)=[X9>Z-Q3X.0E.c^SSPI@U0c@[(NS5#6L)DBMX94-8D]^_N^1=3a
Yce1/]]9bLP#dTR,PX?DAa]O,CV1QO>H4CdQN[d#,IINT)0G(:2Id0.):GIG7:CT
SC).K<,Ed]2<-8;Q0d)X(e/SS=^4J@#QUDa@]DCR3=0gVBY8O4P#ecDN43I(J:&B
M\4F9Xgb(<93_+[O,<c5H4-JA68D:0#U,]deM/ZO1CaGdUV>@2;AE9eORKZd4E._
G6W0@PE9&_GX=Y;&DH2HeXQ93))TE27bKf/F(>07ICVV7Q72\N]\7BOM@\Y_?2@J
G6Zc#)fP=BG8[Ze2\/T^6TaCa[BCG[QW9#5a&/-10&LbP3QTe)8SJBUZG_:6GaQT
./1QM5]e+_[d8WMS2P7D0:VCZB\d07a2bZP3,HG128cU7I7F(>\.P84)K5OeWCeB
-U5f_G\U//b\b,Ne2IT\I3.#Fc,5,W,c<V3,a&a]#.dAMb,ZK7FdX-TY?QH/<RU)
c&DGf;]#RB\MIIcJ4I6G3K]3X)#RC:2E5XMGK/U:d0b,?Ic?X8Z=gL)X;Y=XHb^7
MA.UHDGc533Zf\(\B_P=4A@C#RDN6MAa3cJ5B4.27B<a\HV8XegYB@WHJ[X8+&V]
K0_H1<fVM:]Z1NBQ2@fI<bKWOGHSXSY4RVAYb+K-VK9D33R/g>HA:-Y))NLY)?S?
-?12ROO_O&3f8S2&0d<;?Q:?IHb,,<&9Lf^7U\A4TDY&gd@4_(;XAG-Hc-YG\DGT
NSF.1aW,c5dY#A./2/EfZ&dVZI.J_J+<;6@ZC6+NWI+9[GEVY+[>[M?W?&XX,-RJ
L-)eFAZ/)]c3Naa:R0-C\/5C.\H3;EK/]e.1S2KUa&PJ2B-eT:G<SMA>d@-8T.9L
YVSE)d50X>:3VJSE3O,?Z5Rg0]\NZ>Jc@/D)/0GHFW8,1X5@+SR:Xg]WD5BgO82R
EM)ggGJ>WO^4CbI>2gJ+?@G8JJeR9NOEC=;[58FJ;I34YZHBVcKV^.2-d-4N:LgY
7WCAN53eKT)7-(P_I9EU2_@bNB8F>[_1QA_aGK&3USLWY183\PB=)N_#:TD^;R>U
ddW(<DFRd6Y)</M)\;cB?-J1\(ZOO)geKDd2;;(]7?GR-#+BF&4Le?6/5>:@D\8a
IDWK4(TO;Af9BG=Y31.<033#/T<bQ->[SBI95dFZ#+FX;c&WTaR5>Af2#&]VU;U2
V/WS5,6Y#f&5R0._-7CGTDSHVBM^:=D2-2O13eWLE;5K\X+1Y;]:(IDDE/RE.)DS
3+gP@A3O+4IAPMgf?KUH#:GXS3U1=-\VCR#2^_-=(JKQJ.-7Q)FM<W-QZVV-ZMW^
>IH,01-D?3YVN&S+?NX+DVY@S7MR+:)WU#XP^?GOdCa5?1cT6;XK>IOV(cD9_AZA
NJ>74O<Qfa]HK@MB=K5W0g]PAT=7_dQ^08P1@VdA3EGW-0Y</)9-V85U,R.I^)9[
cW+#cS]1.59S[(E93Z25(MbSQ+e(BF=W#ORG5ZM3N8[[DUU\>4J?JfV.?HL,@OW[
8P3=g3)Uf@Z<O7g.)7=V9?3dYCfGV&&Dc<,De4R\K>;fE1Ob32#T2d[^Qb4T(RU;
8d4S+TMM^.489PCTI1X5&8L0^5YaE?6?-(E>4cXF&gMJH;1g<0N\[&)HAaORN0#5
1/Zc)WX-J0G-FV-<#6a21gdcC7)f4g:.1K.?f+N:BI:Oc,)PKgd_EFe\J=:M?=dA
X>dbfJ;+T>&cAH)6UJNXI4IO/K&dU\a&NV>M0#UM)<Ta.cZU7R5e9?0RaU43MZe;
M-H/e62R,02FE>Ba:4/M.7dXKL0CR,agSJW,A/6;:K204?#)\QRdX>#N6B+eZ]5O
Wd;,#TF,\+0SdO.4M-F=K&-&b?I:PYUDS/d^2D7Pb&a34J1V],?8C&2+CBX:?(<_
-ad3[&(YSVce,8VP-T1]]/f0HB.NNcB,f92Sb)_cUb/4O>Te.\>YI5SPB1)gS0V;
eeSY]VNYc+A)LOS36T,0\Z/7.b@E([2((&#Yg=/C=cKU+b[(N\?8BgEaX^>P6e#M
J)\MF1FVKa09:8Fa;BQMP5RY3e:8=Y-DN4Z]M]HB&]VOP&&&;HABV,<3)eYFHK]N
8eXZ()<E/EE>5=fOZUTW_U0#7Y-[,b4&=4USV]OQOE&.BeV4#R-.TR^ga&?X68PC
9;bW:KD3QFCgF\X]L2=X((TeX^F==GA:^FIR7:g(g;.2FFeHN<&-52b^1(HTNJ#R
@OAaW#6e28H?8VR1NDF)4@@P)dMPE&E.UG9OU@8L[<7ZD=UF\HRO9-PI\UZE-H0g
ID#F4aIS&;P9G9eZ,Wfg.US&a]@]43F+d&gKX4Y@a\M2(<H@\DX9cdFFeCJ-f#=b
QdLe0G[CaKF;\8?@(gJO-:eYeVWCIP;Y,]aHLVZ+O.e;d)U<=bRB><-eMbgM&3UU
d1&HIUNR/2Qc2SDg6M0K/@CTL3Y(/IOaR,8MI:R:H0EGZ=K=MFU=T6;2J_/S5/[.
J313YE6dL_VCb1#OH/V5/DNIS+>^Z+>?^fXeG>J+1cNa9N+LC8JaP@BRS9D=f+&,
.4F_5OJI8H5)+3fGge6#3?K4YS;SK^WJDZ(4E.?M+g\\ILSeZ:Sc+O_TE5EL.1;:
1[.H^5.Q.(\#(WK@2;9YLI<(R^&@>2HTIWX/V^,C.CG^:/_(QORd_ed<>;,\E+Sb
b;2=2>cW@-B\aMQaS>Ae0[<RB>+&G)bUBeS@E1X&BC(@BPE9ffOKUL7VWMNHC]9c
#+3G)IJ3&Ce7,)CJbLZP.a^U3g_?A8=.3IW/J\VZPa7\4R./P,@]P6;[&:)#N=?b
_+B?@,AGP4]KU(WE;RA?:VMg/EA.^aHX?f=B6V4N84G/T<c96Oe039)+_+G]f+]:
;)Z+1fZ(/7+K35OJ36D.HEIE2?#?f/A1KEUU>6KF#@237aCN@,F+E[NL.J13=?a&
1c[UQ3T:SZ]XFeR57(-:KC?E/OKN#@&d-2KC?]U1C9gT^.-DA#=IEAG8.1-@fD:Z
TO+]d=^V>CdIW6STXb7Z>+9N8B53;BG2.DbBJ?PC@MPMMQ;(:b(4WD?G9@1:M]ZG
AHN+:d?1^/I;g)P3CJBbd]A?1#bK65U=dHK=H\OL2:,.EC];@6S6I=B/FO0T6D_F
eY2D-L0:)4:./6<48[3I#G9=T#\YJ3\Z+\S^(YSIW7T;^b8BR?<Z5B6\OM9>YY98
&5C1F.UXGV?=\4#K?.\cP-D^^U4G0BYGNA1<^4DgKc/.;b#\O<^>0>f@cHObODC)
a2CG73\+3/=^dRB7.+LAfBUG75cD4/>_G.H@a@28S[_&N<A.^J?UI81BPR\+0RCL
X\5R4&H/2d2b3@Vc\7Hd-#X9/d;bUXR+9V5L&DHaMJ.0bB361J)c.WDc:G9->^J-
G<2X0;T=S1J4Z6E1FdWY]b-^?GR=Fa^9&<JZ/3U).LD25c<1@R=,66L&I]?=H9W-
Gd+:3VK+S<I@^Sc\1R_HO,BNT?V>V2NIF7c/4]TID8bU0P-F/HgF&c=6^3MZ^(EN
aE]g5ge.D8d1;cG7AD[9SV=D5H17;@9,/QXS-\Ye[L3f8B6f(M4@GVH,@[J9:D8D
+>2ET8C6JSJaDbFT@N;?-M@]^)V:cF1_O\CIbfbcA@F0Td)@3dG;X:GUeg^QAXNS
d8J-CB#=D&T2(8R+,0C7;-c#e,V]P?]R6L;A2O/OU^&(,N0(?6HNC=)+\RTdZE_<
=9W(Jf9OSX9_5=^;Y[X1,PIZT5_SbW3c;>[I57?dPbWY/:IX3ObfFY:W?5RCgbc5
T1GGBAgV3BZe2]=\(M.c(#W@Zb09NA(LOTVJYAJ-&,YXZAP_<SS9>@IEEM5P,]]0
R?+WRK15UYN_62ET,]YKN#4T=^K?W,[INHS+.^E.KB/IF#<Va_TR2-BR&F/,N&M)
B;3TFR\88/:ZKHW=8\bFMB:WZb+J:Z8,JNF=^KaM9OZXR.T)626K8Y5JALL)Q\@]
QE4bW?^OS&b+I[GKL^0QEOJ0[9\+#1VBLHF>cQD#>6[]Xe6dESA[8R[AeXD>Me6D
-0MKCdOGV4Tf)&b\ZD/5P)R5>D/=NV1e_RFRFE&,(DP_K[H-Q+B[T]_M1&7=.?Qb
OQ,b+:)4ab)?W-6Y=VJHYE6(e/bG?5:>@3^&V>1[[?-0b#I+FUJ^YNc^<)=HcfV@
3?^/SXKZ.Q^:44GCD-T1,Z3<Wf@RXL48Iac.dL@?X55@4\[\T7;[c>Ag>#P>c]=D
G1W\&FO]5/Q,[NW?e9>^c@b(]^G>NgW\1[=XVg)K^;MHR@EF7<T:O,A6+,4L:f,H
O+6^ce5QaS/U]=/bPd>8bdK060EQ]cYc4A=\P5E4(LBLQ16TB+[S6XcB/@8V?g<X
2^JSbb.Q5X0())+c>-Ae6Q6(c,1]N9fI15a7A:Z\6)Y14,&<]e7P5B>GVFb4;3RT
W/+JKPU6OMX5T6fYF.]@&F:#RZ.0)N>J7JG]5+RSA59=,@I]9Z90;4J,Q\LDd_W8
V<D-?IF>IKcfJJB43^?5(6J<bQ34Nc@SE8BDVX5S^IbU9E#J+6,A89.6E].JbgVJ
3d=NBSA<=RBBe]W1f0T8W-7d_]eMTM7O]]cE(R/FTf_6ZX5;+gH?I](;(\F>7ETE
>F.\>CbN.7#SfH+)8:Fd/JHL]/S1-_PgO:??.#.4^-fM(KPZaa(\)84XZW>13<L(
^.I>4\fI]N5=:dIC^H3EMb.+7,/O8\@GP]YCSHg;6Eg.UD_.gaUf5\,0KK4UI=c4
Wd(PL:M#0[F>:bGGPPeV46C]SGaF(5CT5?JQBV)5M,BPFBf7bU_[TMO9c0?]D;=c
Z:R3X>2^C8f[If=cCS>2HH?\Re5\Qb-e/((-:S=]2T\UFG.Z:=#bG<6H8U>:C>]9
4C#<.:HdIZPL0QHM+##I_A=JdLJ1Z-JIK?aATPYBTdBASZFRX;V9c)8<VHc1=<#Z
)8J;8^bgK+aO&YH?I70#/2^YMZ7aI,2fK22E&6IQFB<:,E6(@e0D/ZU,9Q,A=Y-0
Jg8.FWYd1aBeJ]e+?:G[TDSS&OO=QR2,bT&(c^UU<V-7T:ZNABb-BAgA3AbSD^F+
5\@1O1-#+66.?VIef2KS/N0YT<R[c<<VJJY[ffMNGBgga>F@g9T8<&(g3?X3g:@-
fQVVLfP@2U64NPKLW/dO,)=LGZ]#E+X./[QC1&,R.c3g_G&:c<00MT#:eS,(BBIW
J\F:YLJVA]>AP)c\V&cL8a>74fCe?V1UTY4PA\>;+6U5Q-GcE)[OI@^T55T9=:KM
\\PfX,_EZVZH48@(?A9B/[[C,1#X9)d7>IDWGB06KUV?[^fD/@^3;(1)G9K/+(+T
)_9TAM762J103N@L1;5FZ1O(N4YZ]WPBD<:cbX1>.OZ^)bJcKW>9_&_R#e,:/a)f
gT7M51BB)g(ART-6(111\;b2PVgS4I_5dAgDZ1,CLKdD)e[(HCgCU4#dO4\J\BJ4
2IM3<80UFF9b,adOVB]Wf27=dL?,38>[XWRKA7aaMT&1gBaA<?SZ^0QaR/##BP:c
-^(&a>A6Xd.;<2aHa&_Q5L4/4J9gabNQfCSKTUCIF&8>9bX.)+(=2VN^e@4g?aGN
Ve_7B;YNI[>FOWL];=U:QL5#1KGgC8]K&VA6(FK4I&Q^5WKPMD-SWJ\,K5RX;GF[
U4YYWGG#&,Rf\M97DbK->YRX-D:F^Y2CV736eFMOe@(N7^WKW0Od\g[f\80:QG<a
_Je48R0_]#?T?O]>cL;bW13f>T2T1(0;R93]CE3OO@7NC[1J0N=,#CSc]WLB4;.f
ea2H4#J3ZKcEcT5a1gcB/^E)7_UO[@&=3-&e_L=b@aN>)),JSCTYfNB]8N+;#S?[
2N\+L[8-?LX[DO#:-e1R<>D+^/X>\F]d0aQ0<GVL8[W4]I1_9VMJc=ACI6feSd<5
M^Na@#KD^9=J7=F.YdBbY471g8JIUJ8))(^3(BP.K,+?0bFJ=WN5&@eMGbSL>@8=
c2K>6T+a\\b1PYaK665=aT1H&f&gMeG+6TB2IUQT9,JK+.4XV<c5@bY#W6gRSD7V
I\PGI<:SSG3aZU_YIVWa[8g;VYP<H1G;VdVG2OY-Md5.DNf.5I<BFB/,BbMR&K8+
M#1(cdB]ReM^/OBeD;Q[ZBA#BZB3A:eYV<<,U?VcQD;OG8W@LZdXK?;<GIQD3TSL
2\G=8+G)e,R7NKS^.RNQQO)GU)>BcPDdA4Ce:DTBR?c&<+2JWP<]3>#+X1[VVK_E
(<(63@,K(3VC3T@:aL48VXf=_/^8,6(bEaYCaX)C##.W;cEO-[3Sf=e9_^@a^X5a
R)@[fc2+/37=-X.USZR?<c#U6>W#@J]B30]=E:Re(8Rg+8b4)JS:e-gVS10DUGF>
SRDP1<O_&+K#V2X9@9:ICg_-X#f(49Kf[:P0Of>-7cSJW7E6U-?Ifc>TS[XZM.+A
L+9_TVGT2C,/:d,,W1e+^JS?a\BO-E1)bS32N9<NUZ^2fg#8]XFPLfg3d<cUKQe5
EQFQ&)RK>#T6Nd]TXYP@^ANe&/SJ)]33/4Q09(g0:a,SR7gTO<,Ea:1GLM09II2[
#=B:AV?dacA0[d@#;K2W++;-/:<F.BA(Rf>g5J+<_<)/\BfMW/)9ZdQfGML.,FPf
T3JJO&C9&UbEV#T]dXHO1LF669DY#?H_.85M>E5VB]f4;7O^.@AcIST?]K40+6VT
Y9-EGQX<2T&1^0Z)<W[]#^CMWgeVZQ9B,(T@:IQ9):H#LTfQ0T.Rc,97Z\b[.V._
LPMCB=/@-9:b<.P55R:A-=PA:CEc-GM[L/BQMTMdZH\Z,B>5,5OS+<eNRV7T@8#6
V3\=bZ>TJ.#D/ObM],+@L6XQF[fa&OZ\cEb+?@^2#16/-cR06c#88^Fb(2EYNJS)
YYA.VNXWdS_c\G9gO\g)7cFT@&(IbB39#.XE:=-&S?ZO7K(#gS##F?&eHC=HA-T^
(2eW.IRW&KQE;@JS9,L[4/T-ER;19dMWae[>0S+bF.OWBM#Y^XL7K(3?Y7T\]0+N
gV@09:A7]afBIHE:-#&Q\(BMaf#VXD8/8Z];>IPBIZMSIU/1?e](4I798G.L=,81
;>DGE?^?@V<6Z0]&0VKI/K3;T?T@E702f\)V1N)P]U?9]f.e,M@0>JX65BQ&9f2c
XC6FgWY7ccI+H9C[cJI5HRQS#3I+9J?NBN15CH[I@9-6Y5eN5TWe/0W2TI>cO^_>
FO74KdB.T_KbPZW&_ZPbX@9\Z?[dZO#38_ES@f@LYZNXb9<DP&a:BE<C.YL9P_PY
]@5C+O3QXWY(C7RbSSfZXY757)\L09)gC^QMOJMSg^Qd(^4K81HT.b)B]gXX:8:;
d_Ye8cF6FOZ65Y\Y:3@&_g_<8DDB&0?B01e1Ff(H)VUA_e]W9_R^(RB2TV=CMK;X
?S8LKX-CW@F9R/]D<_K5)K4FH_5I>H&82FE>G@21,)cb][1(:QgF1<?d4]<;-HQH
eg8ED?=IFgf#=]D.?.&)04L2#da?/@@?6;^=B#E(+XR>MNdE^:G\9&GWSO=EN1\U
@f_E.CF7YZO<-fZQ,6XdOPA7C]U,/d>9b2PMWT-/>/FLdD/F/e358FD8JGC<?ZB(
&2\9^78=Q)9)g>@A-d47:\0IE2OQ3>K?&Z7[I]+5?gXe@OY[I#2aT5?[ZHU/IF(6
(NH87:K&#b,4)\UcI\3b:4_8\,a>^eb0W.@E-d-8<.)J;0#NbTS\Pd9Q<Z^aZLC/
,4#;e&252d>XGP896/9KaB^&g.-#CSA3Fd5UL[fB[+bMA5F9MJAXPMc([B_9<e>#
N7-BTM9;(g]PZ>X.)T<>?VALdNZY?GAb;62=R7c)Q\0-;;V]N/4.3&d];VZV#X-6
C)2MaN&,Q,J,U3U8c-=>H@.eK3PH.D7Uf,JO8POPDF@LW@;X0\.KSJ=NMQU:c>VG
+LJSY90#eK1N_f+AW;.<+N-2L^?QX9:.+:aZ_;b2^;]RM=e>0:c6Jd?0<N459;T(
PTcXC,,_Z8V,TL]bE7MYARC.f[_fcH2K444TA1QcR@A:I?e\_W@)H>N;/&J)F6PH
bRAFd;F3fV7+.Z3K/RGWDePU4#58=SB:-+^H8J&:[P,KHdY79Iff@A9McX,-N?)2
-(20K7S<E(Cd>[I]X7:]-bX@>F/ULAW@QWLS,;Y;(EK_3>P8G2(f#I,.A:]#_SPb
(60R@HdQO2;0W],XI@-&TX_Q;D::V_dYU#Fa?-]M[L^-@ZPPdN]]M=20F-.K;+[G
b:<@=354f<XC=[_g^c9dC+J?Ga)HWaX1GcINYaR&He6=6^[E&&^6O(HY.]JB_?;-
ADPK;HM)N&dZadOMd8M+W2N&4MMb8D/c2_SADSQ+cf96XY>.@D?B1[cb:\aP(N1=
E(]S6:CTG;L?(J;^TcA:c@D1\)01.:c7&3a@9D@<)^N1<(C,Ue<:4>cD)/Bg-[Hd
Q#bPAK6\F\;J;9XN?M2S);GQ]86.\41E&LW0RV@\E:V^J/G4CYXRZC_O&WI5g00c
A3\NQAS/SCd_JE:+:c5U0;6#?86J?cO;ebcLN4)KYS\)XQc+,^S63\T7T45:)M=)
\LWH?2bZ)g08eDKR?)U8R0,XLC^@<\+4g:;MIC^eXd3[Y7=L4_(7UE\fageA_IR0
(W>J==-L)/>^R]Ge>R_>SFf.^)<NAJ=_81WK@SP9]f#5d(aYC<7:3KU9RKQJW91?
/8fT46Y^+T[&M0W3[df=V@@;UADW0^eT;,<MH[V,5LN2#VGWAc.QVBW9/@?fND=1
;Og/=a;W,f5XgO#_FOD(/1]ca2J,DE1_BI+79L:0L?2I8I@U^+)\_43NJ@U)&T(Z
-ZC)fO^(J[dEGc?25/gSXXZd:b)_/O2?+3J<4BPCJWIV,d3I0=YKO<T8YXV\^g;?
Z+XW:>5OU)/=9WD=PEWR?<8C<gebge+ECG)Xd[]R06#V0,6\a3TA5ETWb5g=5eI0
c1L&VcdJ7[@4P;f>AdMe2WeFV1&]DT<RO^;S\baR1V?H#7K0?,0L82\RWS3U<NG:
F&Z:5J,H>M4Z_Yb)T@,.:IMN[d)@,3GgH,dLBQ:bDR[1XKOINS3,1g(--U<:O^_W
e3V?-Y/:d0X)K7(Q^\_\=0L2/:)ORU<GYHT<SPI\Z9(1KXEK2DAI05C(-^b,gIc:
?:@32@Y7cOTBc)KV\>+4:K0?T^[I:&V)f&E5Uf]>.=>K107[Y/J,EeM1BFWJWORR
O>d,f8KFf^[26&<0MAeA?;b>AF#?4V8Y]]QZdI9NK_W+M9cSK(.0]<a^I>bE>RM;
<^,BVcSafSJ0gACKP;GAb5##1-?/D2,Cg92G&8?5R;]X&D>3COCM&_E&8]3Y\d\F
\KL>564N/&7I8S_EdPX/=5_@]00/<-V\ME4(T8)^;9>HR#Q=MI@aU.+Q]U;ba75R
CHgLC/He\A\N:KbF7T_,b:,<2;ed;KOOG-.)89&4U.\M5eBRXI\A=A]Scc;??9=8
9GJT&)dgGZ/W_f>_DV=d:0<YO5d3A<:UOZc^>_QSY0IZM^6EYJSdZBPfKN,BM>#)
V2<B#IYE56/gR51F]:;@NcOMb#7MD)<5JI=[0L:.N0cV+NCQQa_RR+]W?5Hc+)9D
d]O,RcXE1#)K#HfD@2I-F:RRY9)(e:5bcQ@J]d8?EL9G)T7CQK1U;(YS^,Da9B6?
e]^]_#-(&UP:fB)BMCI^eDF\JbBgQ9dgOQL<7V3g6>gW<[YS9+=AQd(?TfD=H,BW
[5_>:60([YAV_Y31MP4QAbGA[S1DT-D7g4BCR+b+ZLd0,b;2;dG?98;<=E-6B6-K
SE:8#bNcgT,-)OL:QQA1.9>LV=bN>HC+9J3^H/RcIe-+=cMVJ+IF.+QH<GD)VbSB
\P^@EVR)T;TLP)&Q^e/.6I=EF?VaY)^Y199M^2,-(OWA?0GJ]^>582.M4G;BLE2E
0.+XVNR,;VX<40dT+IV]S4A4HBf503dC.]B(5DF<_gF\AWN&>afDQ+=MG]/,:+_b
4Rb^B]QGa,)[Zd?/^bBCVLCO#FVaVHY2YY#8WWDa:O56@4\LOe]3K3d3(>(DGdUR
FQQ1;B=G3SL@b#I3cBBMf9efJV3Lg34eL)-Z]68.&A0?WY^R/[@V#^#T;W4M+0;^
?0I^ac->d2GT.e.5PIKGU9L49L_bL^<X#J/DO\+FGgD)EIaMDO=.A>Fg.60R4ZHc
19Dc6)1B]ZM1gV:443L]417,H@/HB_(HQ744>4_K?cE:NO0eJ(,5c]7/ZD=J:1)R
R=JdZ@WX\Ie#2MZ#GP(GY<KYY.Q.g?<+8UC-G8XF=0#UQNM7;RM850,?TLGZ^gW0
YaT5BDeQ-;[KOZLR_.(4:&H;XI6YbD:2CH^6#cLLN_(B6.(a,0L\Q23R:<2R7)(-
IcHfM6SG>Pa>\^^)Z>:)f67WV0(\K#NTQ92I>4H1Y4W3]-28N000,+NHV;2F7@<D
)>0W4EZBN)W&[/)0FW^;4=XAfPQ(AN;Kb#9^>5,\COU/)/FH7FD,QEGag:,<74PP
#/]/Y.H^YZ.SR(?BFOREO&I=gd)dA#dQ:ZWAP]R3#SPMF1N.U3TM):FG-]MbG;T;
=>b8BW/-GWAP,[V-??M3.95V0KT38]aab.5A5MGD)3<7W3G_?Yed)#YVYJ[S;bbN
6E;.N(PK=7C69fegJ#EN^(A/SMB=WM@AL^Y]bB/KBEA=f0)OW[)U;:&6YE9\QB8&
O0FdNXN8&G28D&e>N:</(UXf[(T#T6W,0Z.W,V>\cHSbbBHV(d)aPSW]XRf[Fc-R
Sf8V>AQ4];V\-IO6Z@HGOU6@)e&^=0I9IYcU>e-2:N3Y2.TScaZ+9U+f)cONc_W\
+Wg@;GJR[F+gNfa7G)f4c/4#&#U.gHbIYLK.MUJ_d2)Z)1;a+T&^3N?@+PbNB6FU
&MYNGT4MP-(GZN^UW>5<(^a3PI3bbg-Z5U-bA/<P@I7S7+?VHA2gb7.V-BH(:CcP
-;QFcX8,YHAgA,&]/?>BBD<\>\)BT14OM->+0K6,?ZVL=O=:a4,6acUeY5I?e-gP
G6Y=cNH1\PIU+36E+NeP+_Mf^CS_BB[F^R:L0TVPg\W7ZPC.LF[d9J3[-()Z,QQO
e9f:aaT9]9V)-9a@U-JgOR?gU6,8CcDb\/>?4F_B6N_=C/9HM_G;86M,4TLQS6V8
g.cLa)c5A2:>/E[K&:1e&Q0)[R:dbRKU#O<E_RQ/A04K_5MZE2RS-M=>[JZ):(Oe
M>L5EE+S&&Bc4A_OYN@a2?>D)EU<6C&b8&>5OWFd[(?[Z\P6X&Gg[?6-ZALXZZ?A
If/9L]8FG^:S_;5:HMG_J.;2_R=./W4Kf@.:J\R]47J=,Zge<6/IPc,:2CI.VCN;
(=fKD1;<W8cP?Q5_.P+e(4MMQF]\4.XASe;:1KC(9K^dYUabY.IfP_2U9DZ+c^;8
0abdBT69b<&UP^3]5#O>HVMTKP85[,HQf]@BdAgI/KCaYTeB9=cDf_OV(&5K0IUP
\=[AS+]?3AAU7=>(&eF)IJJMB49QC^gR^X+\B.6=</#bUMdB)O9)b,RE8C+]^8fT
gbZ1#/g947L#V7?2R^Y@=\LZ_7dNJ^IPf]?._-5_BM;#MK=:E@KV)QBELbM#1(=X
PB7ZR^-,5DX7.QMM@E[,OUSPRGW<<E,YO<(]^1+=He4LXERL_dC?(DeGa-.;5)S.
GPW9N_6LX<-AL:_VB=1RMM;FYgUI/O<#-HG+c2M[=4)WE2Y4c2C+aaY8R1-fR+[P
Aa5UPEKJP#-^8K+4?&:M9:Cb51]+eP.:K6MW&Q3O-7\(MQRIe>[?;c\H,^Q[&Q#6
KU(SS=?)J27.g+a@Qb.aX+Y/]g6SP[0<E\P8E9.J,DU1+6TAU9;I[,+]dbg8RCT0
D?YVa>]-0C56R8N.VEO3[/&+RE]LgfAdVEe(eg5c@IMAZU3B&4#G>>UYf)d1f+O1
?:ScPH3JOT:b@2WUC;.)F>OM:c@3PYTLQg,g45eJ6d12\/AJZA[Z^RMG5-8=2_R[
++QE>3=DG.OaH;3/P[<HHX++Z_:#>bBgc\7f?XN5fcefg?>[BL5\CCS6_.&C_X2R
Yb3d1-ZN.A^8CNbdRK&Y<V[=3e[/IB>PUXffcD,ATVOGIKgXFVG<#L)d+VBgDIGH
/S/_CJP>,\561cYVR+.BXTR+^-:DQ]<b_3)RV,f._M_Y2+DXF+6:K/]H01(LcCB\
BL8BXa^\U[b42>?:CJ0N+UaTK<2>gLZ6NZb^4b[C,\>QY^)fPG24><c;VC#_3X^^
\&+D;5d81c;:RfX=50EgcYSH&[6T;LR]PJ\A;V#0?X,T,<I3=QVXbT_JgQSf46JO
RZ53P]S\:J-IIgf<B7]M@)-\7A\.SKF2(38faRRfX^=Z/I.GL8)a==eMf[cae0@9
Z_FN\7-TNafcZB]=N#bE4/C]EFJ^03)BLC&9>VV+93)WcKM(/0-,\;9=gHW_^JcW
#8<&0#;_U=fL1X0L_0>&O)e8W85dCNUV1G]HQJ2.U/Pf@K7WWX\b_BXKRMV<9<X1
.FO=QcV3#_LM:c3;8^/5[I8ET([C&\G?K_B=HG<-RLH,WBJX>F_><d:IVCAFLB^G
?8.XONQ@@-2Kb6BQE#9F;K8cK=6Z,e;7W?1DX?^.JLeU/IDZY&(MSB2(;8B+Z\DL
^<9gV.9G(=:@1\M&]X3SXK7N5dGMbY8A6B2L^=[&Md\bAHfV#WF.fS,adV]J3?AW
Ie]7<?>(7[\-R;aTI1^5U0aGAK=-G.@OW^FDK):2Y_B7J6]]>9HeZ&TQ:_b620)Q
^+>dMgH7.J@H>W1^?S=QX=>Fa2aN5:fbXTG5HbZLS<O((FL<&G33;M5N@R]?-EE;
@<2_/]a=-\+.Eb@Og,@LgFK/UebHR._0R,7(<4[K+-<^[HFW/VLId5d7_.^W5J[C
.bW(6ARC26dMY[-=[&R@RX2O00gSRCPR(;6CQA-MTXLQY#)VG/<UX2:^-eICURUA
B[5,-;cY-.&H=2\O6-P(9(Ab-b6Q>Q2UBT<)ZDC=MTeB(0^W6[ZN@0^L9G[QR1T1
5QH;NfM@Bg/B2#&L)MW3K8X)A,f5<]N,4#<GDS<c,6UVGU):DF=g8#J^PdD\a=RE
.6/ZJL6I+O;F/bAcHSBG6Y=OSN:C69+GQ7fRM2TI0,:0GAR^>?QgFU.gMWc4N;>D
4T0S&4R1F]dE;LH\^-,D(JJSRN<D;F[J[>^K(S/HAgV\1+@9TAJ7W3X7::.D>?0#
EP#[Y(&1D)T5EKW2[81O#B@_.<+f4fGSHD(eTC0P<O>Q5Pa[K5>&>Q/4Jg7M=]de
]3eT#7/?3I-ZXCG?e&^C.YXE4V/eYU28@^F+X[PP@(\5(bc_=?.<JD+K\/X0L6ea
MS[b_-JdD[1Db-(EV7g1E^dABXPC(O-=5^Q4gf7a]WJ<UZCU37O>IDW)1[E))]EA
I:dLaXa9G&U\8B+KZM5>HTWN/V/ORA,?MJ)7cBA(/MW:/Z1?N0>ZU6-W4F2cG-E6
5O++Y]_=?YL;\@O&6@W^[0+XK&DB/4E&+I4EV9AFW@V#_GcK<<1N:1Q&?FK]2ZO(
AT2GRM/b3TPf(&@?g/(HRe+9G50&P/OL2d32[0E\T:#:<BD.HWEO<;eG20HbQ9d7
SZR64g#POYUc;dQ@5B4-P2_&X/&VU=]RADeN&F](LAb:KNdQd.OGDL(a[K]1JIK3
@#/JJZd&]-e)F;^,e-,R2+Z4.aWIA&1]&D0Y#655L^gL\)a>T#UZPJ32_-@Ye]NY
&,4^>Oa0BU&[Z.dX8Ng8eUc?B0f_8_X=ZcKL)YY=PcX=#F)b[Cgg_?fNB4Z1dPaT
Q2[e93[N36Y0-U(,,I>-GB;A4WW(I_ec5Hg9PcdG0&=Wg/#&VJ24BEQ26eKGO\fX
^?&<AQO<&.ZNBN7;FZ)DE-FY0[)&SV(Lb+=e&bSMf6<P<.EJFXW\H(@WL#?,@\b0
4>._TA8a\/?R?:[ACM?Y_Q7RV:7;>L<Of)?MU1Y8,#_U_^;4d352JQaZ(WPYG,)g
_#\ac\H2+&5AW2VbFOOA41:8D5+bVUBgRC?Z5ba8:>da4Y]E5^X_Z]@XED=6(>5=
V)X3/W0feHQT7EFb^-D[.Bgd65[.H0Q9g.N0BLdTK/GF:)644RV76/8@@/(3dYBH
cW)-/<YHc6a(EGVUY)RB[^V]C25;XIcESX<c,+-V[C@-Z,YDceTWWd+TPd6BL1#N
e<LQVg1bQHYcWHSY?2f+IY)PN[6GP;IAVF#FZI2f3\D0&CC^&ZE3)DZQI.3]OLf-
4>46T.&f^<5G=@\bS,cR/)+gO_[XS9ZD<eeLF?OC+[L73[dJC3?3>)E@9^#2JLNQ
^:3E]NKc_S01LMRb&bP,?8>Q94N,TRQcaRA2QJe://8TGT+1V>;+0ca=c<KDKMJ8
0e(g^Q<#;RZQ\&GDH75LFR3T2E@H;c7Z0#V+Ug0:dd<eKSfS;8KJHfTI]H4CW6K(
ab80;/A1cgDES#A];C?6.1NbWI).gc@/.8&g#_XPV-5,/J-&(Xe?SFD,#Qg=TSJI
C)/_c,[RW\GgQ8\-&(X;LAS=ION63SSaL-:gIfEDFSeQgfIg-?Xe-W)+]gd>@VEZ
.QPG)CEg\EGK::&\2L:^[aL76,-?_)KYaO<WZ97;<;[CU_7VZf(IPB?;YA]/Rg#2
->D#aPd.1f+RK?=FdH;]T#GWdG=CV#0GV6<]OdO]cV?LAQ@eV&6TZ0dUE;JS7=X_
4FUU-2gQ5Z6&\KZUX(S^Oe9?_5&06]#fX_TXZ7<@TTQMG?d:J3/V;GdU\Oc(=JRH
#9fAF4:)a.#)\80]/eE]VZP2:R9f0H0ON56RDR?c3)[+O]SMZe,KA<[91I^S7RZ9
B2AdgD5MOfa_6&eKHAF6(4LR,,XK+NG-0T]2]X[X_Re&WO21cUYbU2MNf+I0Afec
G\,]\Fd+MG9^E;:J@D6J@RN=>;Y)CE#NIY[VT[3gVcAS3d/KP?EM2cA)@=Scf];=
YV:TTJB&eZ8LD(aZ-3R#G^CGQ<BLWR^EP>,b@NYO&gObHfSRT3@IafMSG_CO\64M
>VJ#0UEKVS.F,F+ISa5Z:c=)OG4P+GJXA8d&d\TT2&NC#[3Y6e.GC(F-4HL_HcgF
0;U^a:I]LMM5>^JYeJ4-a/Hg@H:T86L&5QZ\\g=db6WU#RDf1Y&J6cTdBM/#ZYdP
[0?O[=T9+Iba,TOD_)&9b]J,XXLPG2_6.bR[H?\-IeaW5BgMe-gI:T:+/V7:b_TY
HL_PPda#]T^4(3]-;[KFY_95&VCW\.TTK&._&XBE)LcCUg(UU5B#UV5_1G\D6/E]
3Sa/?ZWHQ5#DTC5B4&.fKf^L7Hd<@8YTUL,EW:LW7Pfcfa7TF:&2+[2W\Me\M18X
-5TNNbW2,VK@MKH>,AbRP7I95?MJ_:_,c]W2a#2E;:_#MPFO88PI6N-U.GGZ3QHH
,HI(?M&Rc>=UXE[GB5)WVROFYeHWKL)U?I7bL(?Qe?cU2,)c_RJ1Q+F?W5\\:K.M
fgB_0d?1b0MX[@^?Zb@3SZ9\+\[)W\ATSe/W-+EIeg](,L+[#9?TVca702#f8MQ[
T9F7-#L>b1:J(F]<3c+SdP3U+AY&C?2a^Wc.aA-a=R[-/YN6+.@^eT+O8/.g8OEK
b?dVBOd>=e#T(7.ZJ82F<1IYa>.-[Rg3(U_KQDD:?-e#ZIYM1>g7D)T_H,<Ube@M
+F4^Fe?,>b2Pc\Fc7;dA4dC49>R?L9IfC)F\1eJ7MZ[P(1D??4B_.5f5TSF2EH1A
OIe^0TT7QU#<JU/48eCE\D(;DZa<@8d_4J2#7X[]#@=EZS8X\NFC-9Z6.)5EZgGW
,b(e>_DAI.-+]fQd1.:VUU395>@EESR=WIE6gWYc7+B.BC-+C9ICT8YC6RBa(UaK
9IG(Xf^F@-G:T]8,\Zc#S=9WT-;E:LcZAG\Z=1<0Z?.bM:#K[=B-2M:T#bX7NZ01
L-S;).;b]6VETTB1[F-/X^gZNa\)eb4Q98d1YU1<],63.aOQ6IZ<@.+4=fgT17XS
UZX7S\J/f5I5b,.MF@gKcWA:bVCVHH([c>\gF76c-C=/&cEV_MO_eb#+AaD-1K.8
P0g\^::gFHaO;VF<P5293XW53M<IBI6G9V3\(ZQ1-e_[OeRWZS]C.8KTAOe>=-c@
d#A92BH<6b<]-O2TD_HZc>3)Jf==K;b<KEPQW&#-\Z7Nc(#10D5d5_WCO[>&EScI
/f3\a09S@19-V;f&W0NPDdMDPJK2O8;T25ZZ<JYX9DY1,VgaNM[]]\Z8O1WLIU,\
L;(BY<?7bL5B2-EM^TW))BaQB)/(^HG/aD=0(-\UWJYWE&I#^/4&Lf<Lf3O9S4J8
0Y\27NH_(S.b&6f]>B3V2WX5VdU2U/1IZ/0Ya+T1^=M-V1O3?+d^c)AL6L[/WBK_
+:OMU1H7,<N-.]<-5;JSd>G#GEG\MHD53@OKJP+D(7[Nb(5)<9DK&Dc89VC]__:=
3cEeAU[Fd;LGNJC<dVH9;^X1WT(4b7e/Y@C<c[8-KVI<O_DFb5\b-A7+,<fSFR+c
4VgYT_6PD3G,D8P^9:KNgD^RYF\BA<FgF_PC..(A(N:3,F,gUYIR^\]b(12<4#RE
=(J-bc@_-g_C=-542PX:8P;GD0GFAJ2b0=WQbVdK?Kf7^LT0JMT<Pe4?(-)5b8+J
7b0JE2Tcb:>0NOA)BP.Nc_e-6@;8dFA+TX&Z0g6/?Ub[YCY6DVS8,+)07BfQ7KSW
5MLR2>QJ&6K&PF#Z.5AL[AE]@1b59fY/QReePRLJ6C_VI.1Tg=VF7K@0\d^THaOb
AdZLDB8fb-B4).S)4J:6\WT8gMf6Z@\LD7@aIZ=7eEF:,4GgU\N8)<f7gQ/;(3]A
I7P&Uc6Z>BAH[)SIcNRRR)ZE]+\W/abWARE)\KFV]W-F/S5F>9TIB27a+9&5g9LH
?b^0RgLKB)XP5O[aN:)^f@#?D\>=I&XMY4,-V[#CSDA5Z/g4I9^W0\AJ:^CZZO9X
HLSX(/f0E@ZT6_N.+eGU6]\QN)X.V8=ARO0(,=FCV9YT_V/@d@&5=9<)/6gfXW7+
XVL1(NY-2f<HXB=3cR:[AL6S\OS^8A+d8Zb.0fY3L7,SUR4Zf,f<P16(4&1SRXg8
e]_]<J3daL=/2.eO#9dUM?GM-QD+Z/#9378d_#=OSW@:&U1^,BM#G35+cG8GH7@.
)a[-2=QEX(NEHMb4/T)S_L((4PQ@3#DKSBKB,(AWC9P\fS1f<C61b[2@93<#ZI4(
g8;UW/?MWL.)14+5X[SGAI\>W,5J@V>;J1d]ZN.SIYf@\QQXgbN-de;AF:.#S&2#
V,JK[P87QS=Fa]#HN.R#==@@E20_[g7Ic5C\/eZ>^72G]D)EgZ70#\-GdJU@9;#@
QTT##K.4B?g_Gc<DgA4TLDDB;V?L4e&@^-Ag6/>9]=.G9>VPL6BSDG(WeDYZb=D[
?HHg0^K1\N/[I)L=T)\5Z=9NU76d^dPM+E.,@U\15>DP4X0@=3EVbY-JV:4B=M(I
XHF2#(1V.RY_\K]F>B(WC>ER5H^]D4H883=d0M+2QUTN4bE;SM&A>5L=38A@6FHH
1[/fYZT_HP@XO@Y#GYX221c.dTUP(FM08GX5Z\J=IWS,dD4a6F_@;D;&:YQ03G<8
F+XAOG//S:[S^1Z@G5,:SNDJ7Tb_dKUM>PK&<UT:YH<cb]@G)^+WKQa+SK/b^(0J
:YBeb=1;^M0PKQ@;6F8I1/VA8[)32?7.;V(4_9<HAVE1+KEQM8Ud1a88QMK=,3[c
@3@bVg3?-1HbMcD,4R.aC4Bg3_B_6RK3AOLEOSUAB7_K76;\L<Yb:Qg]S4fH)#3Z
?EZP^B@g^C.0VJ([2GZg.#2P?XWDK7?=IRYZ@NeeB\EcgSQ?dW5>&_;[SJ=]RFPP
RKBA/c[V(QdPH\,YO@<GBLM.]80S^;DFG(DM\YZHQGXd@=.X^,ZcX>_^=FgA2cA1
[KB0]NdL_MZ@/0B;R(,MBfM.8$
`endprotected


`endif
