
`ifndef GUARD_SVT_AMBA_GP_UTILS_SV
`define GUARD_SVT_AMBA_GP_UTILS_SV

 // =============================================================================
/**
 * Utility class with a collection of routines to assist with Generic Protocol
 * transaction conversions.
 */
class svt_axi_gp_utils;

  `SVT_XVM(report_object) reporter;

  svt_axi_port_configuration cfg;

  extern function new (`SVT_XVM(report_object) reporter, svt_axi_port_configuration cfg);

  extern function void expand_gp_streams(bit response_data_valid,
                                         uvm_tlm_generic_payload gp_req,
                                         output uvm_tlm_generic_payload gp_streams[$]);

  extern function void gp_to_axi_master_xacts(bit response_data_valid,
                                              uvm_tlm_generic_payload causal_gp_item,
                                              int sub_tlm_xact_counter,
                                              uvm_tlm_generic_payload tlm_gp_item,
                                              svt_amba_pv_extension pv_ext,
                                              ref bit[`SVT_AXI_MAX_ID_WIDTH-1:0] gp_xact_id,
                                              output `SVT_AXI_MASTER_TRANSACTION_TYPE master_xacts[$]);
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
FHx82/Dj1zsyhSlN8tA5thE8fXirAn+oSwtcoJnF28tk0AXiazETAxBgly/JWYLd
yyk2L9wzHf98Jyhn6BpimRwdl7nz7wN1qiNy8zXGlGeM/8OVeKVJhMAIIoFyUEGU
MDIgNMBlRyBCn5DbjXMyI7T1m8H62bvp9quJOazrZPE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 335       )
+r3Ve2qkuAVnypIs4NL48pWCwPDULm85g6NCBFRuvO9wuS/vMNd+tpQajPi7nY9e
TGKXHwf4CFgMnw6YBkKxdDCtBxbM+1r5LmfI5VTzQFj7OranD2WCeCekpinckapu
jDgwfFNKx1SN01q4JAJXeRvAacQZSEgs+FuByvZEtZ8hoPlzQKvu+rIRgUVf2fKf
XgdhamuwMz8x/OlI670fky9nxiy2BOr9mixBZjAzQvkDgmAuCNoD+BJrN6v8Kxfz
ToKrGV1/xTFr/ZfvQeC9DKl8aEG5ZYX3VCIXxk1+umH/lXjXv4b7DAu3WbshJK8E
FZaYNiaSqI5/r8HloQhLekvsIIU/NeBJYENXSV+h3E58/pJ4kiK8zPO7s8Zaf17v
sPkA0kO+qLZ9MH7/6h0dOIGjCzYxJrEYbrh/bFt0+7R4uoyKvOwELhNkm1nBdMtg
`pragma protect end_protected

//--------------------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
FrhLpP0zQ248FYSJhnwOwwoxSdG89Gj5slhdhTMLXakELdSrTMpznLUhd30YbRbX
I1d5duPsDE5b2GCHWL7PMcmPE3klRtIcN3Wk+z87bQ0Pk7z+V/O06PWfu8svSvFG
3cuWEUSlqEXXaCk5ILsDQWXKezsJ+6q+m7XoKQs6KSE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 12008     )
1aUEXoa6x9hbfLfR9/TorNfn5G7vAyWRXpyn3zGtP1RNkWtAWlXtcjQj/h0+VFSk
/UACM9Jr732qxn3v0ZOFUZwboSkLkvkCRXHg2gygJJjCNlXaYmXEGeFq08C+E9RA
l7bi3oa0X2ZtjvQDY/7w+mr48meNJGbxaq5pKiTFxcMctaXkjq1BrUq0OJ5mJaON
rdlPKHuch+X7INPwSjZ/IPi4FyCCg/j+Jv4IfFiSqpKzrMHq8Naz/J0p0YmPkniq
yt9kVgPfX5Je3ulYwzAEboyQuvOfmPedrSCOHwGRwnl6LE29luYXDFD0a73Rqlia
ZWR1k8rK6EYUs3PBafE89vakUOqg4Z6HEx3MgPfmBVJsKZS2zaSHhXiUqnpc0/Bc
dcstAakLeMxdWlom1Jb5vrFb0hFXV03Yk7j7/0p7cAJu5i8ZZLrhKVUNC2ZqMOnw
/PpSySEp292YGYq8ajuAfjN5hvVKLCy+3KDASzcQEYUNKlFLrQ2xTpux+z5KXbNL
1zuGpVGWgHLovAR2sKBfHDYD2o0+bvCtfmWgOSMxM38W+C1GJV0dieiQD8jc8F6j
EEp0ch7N1jitTunF35cCv1DET3EijEvSPUWNOd18LSK1/KJO8gY0AeNnp+h58Xai
MenqTnjEvWZdA9CFL0hhdpSTMMdciq5tjVo8BSv8UCPsQYYThkSPHuhPzo6zr1HT
cz7p/upA7HEnYto2k84F1hD/yRhP+OCczsTo8uLcIzLR4K0EZVIY09RHSDaM9p1B
X/h9PdpaCxlwVFJHzLhmUV8h5kUINzj8PZaMX03vblELLDfstINQSMk/XPIv2pA5
KXIPHO5lAyJX3N1WaC577NHW2PTCXXfAvF6Fuq1KmZbC+kG97+qqmdzN46x4tQvN
hk8qQD+CcbbY+ZMob8GTeSjeFXWksya3hX8My+9UknmQB/bbOXYw1N8Yx8YrZ+e+
tV7jlJrzRmtTipGLZ10XPMGmGvbOZ18Goam+48ggwRSmTadH6bBCpcve7NKfwgzM
uqLDylTlnnjBoNuJhMVlcZ6VndVCQqY7m5Ft7gpAEs0mblYw0rbwapq4EBTqM8YO
NoIZsWkccrze/b2R9T9ntICMdsSEme1j1FffqliAfz8HYIq5t7pkSD/TXV9nHOpV
eR11fYCvv92cfNy0KMcgnvdLMmgIk7xLwuyH/B34yecySaKXnyqe2Gc9W10rGg+x
bQNu/p+UQdrxuHCDLsVrzYlsv6csHGLp4l8nndjGCvsd7jEaIyaIgtGtIz+mykCL
nXcgL9XCHAPgW9bkb5BHn3Ti7PK4k55If7aXPpiofbiEFAtFCOaq9oIzUMi6xweq
7hxqw3OwFu/gsZ2B8HU8OW9tuuWDpuBU5nXaDFLemE60+Kk30My38NPkS9ijC0yS
jE6xZrn+JJnM2TNNae9yoDoMuytKSKcGKUajBnqGU8dLRQo1rQU13XMdq4wwf1jU
B1jzHL/L5EtjxSrPORy90BhBwb4dHM/BujDuyw1u/Ucf5l49aocrXmtTQK6aBpRz
lBEUZRvVYeD3gwQqCFz+TDXNq7Azf5FkAwpIHfjtl+/AmM40yOZ/3S+kPTqys6He
XSiXe+ZMga39yVHaSt6JF+0qRFN4dJNyYtZv1dQVj4uXVk9E4p50ewfslLYU3qXp
rd+uFX9AHB26c/0cHsVV3GsyA/QFW8xM2W17n/MODF8kUJVnuTHmlZFZ5/zFd5Rh
b4LegEWCXN051m61Pa1P1aMapFdg2dQKMxiudPiUVks2dRFt3CoR5cgaBjV3tUZd
YYjNjTk8hNKEeNZdfdmOYITapWzbCRHUN8C0mE6TGA9a3gknJUuZHSjVp4CbaDE2
ci7TIAMZFmKYvFWIxVoA0lOgrN/vlqm+jkDphZ/sBFdmPignyHw616MWBPkWJLXI
qZ36DjrkBMl5jDSeBgWFlkRH7R4DfmVOzBtUeybdOK/RBKggxdBxHpSRPpwn82XW
OfR4HnEVXL1GUo5ht27hey6lGTOjmCyastOUN4Lw1bXhC5mv+aXRh6IMpLWPRxax
RhU0xjHnY3FyzY057ynWTZ8o3GUKUGi47a9OkPtAabjD47D65frvDDoeKfgsKamB
p5tGAN13vU8ie7jtxP0pdGugcilH+ZA5z0KRCVMO4ExyKV2PaRnHqfXjm8iLXnFr
wAK0J+ahU5z8WGrvuoEWJbiPl84By8iYvE+Cq04geHJKA7TQUW7KN+XyfkLH/Jr0
CrbWYvJ/y0VV+MUcsSDeedPlTvIsB+ZhA15tGC3aU06XLBjBJM7sk54d+QA56u3f
l2dI/0vRd9X5GHFlhco2KGHeMvlDYXq0iFaznJOaAJMN3h1tLYFr8jjytEtjN5iB
5IcET4t4yidyLa+IwQ+s652jPy5dVLzCmG64rWBPNijvm64KC2qMwvw0zCARYvAV
lwuTO3XqEispbnb0L6k5pQXUpI+p6/iBDFoKnKphkSgU8vGOXX5q8BJ/j7FYGD35
TAu4UN+JDFw3+cnm3Ik6IJzZEfWgG7YLEPIHTG/zjs+R59yzZ0QRbwGFm6HiIvYE
b5gO1+BVP8f+bWq/wvBW8RVmRCRac2ktnvB+VVwSUzBVUzsOxZznpjWgBtsykw49
mO5steoYHsODMEeTzVxe8wX2kHhrGJc86fxpURz82TPtEhH+h3kz4kP6XndLyZpM
StQh5txDEWI2jZt1zvmoZ3tOHLXu+8YXLXTgmt55Ys5c5J5bML0oIiTq/GogZccy
1y7sGyBhzPRrxx7WL5fpgQwysosCQ4uke7mVhXUcEOF1aNOwAf3RhAahMflOSjot
kxkKRmaxxuWjvYHtGOUeDlbboJRDaCbsLGMY4pRvvSzpQZ7+Ubmhr3HMaWf1WH+q
FGWd0iHZcUvOzpE/eQS5Hs/EWXYMGSPGboFbilz73twlNiUAkpG5vEux3PC8U5UZ
MeQHEse1BstnqYKlJhUTJRRLLu+WQ925LjYWFl54tTqBi6OhEbMq2DOn/n5TTF9l
TyiAstgaXCkK5mhDNfDaaeRvEiGnXOcqgoLPeaA1w0+uMIub+Y5oA6dg+gedv3O+
xGMzV87JkA8oKchLI3InYBeCv++8OysgBmBQmqQOu7n/zcc0pUSiVL+m/JKPRQ3W
nOERidiWqbJhnO8iwjMSzQK2oNIP96023GTkfcbPvxIbAZT4K9ZRhObQ34O7l2V/
ZRwk5tNCRDXiEkJBQMVc8uY/9KF8xbhgBQAagGy6JwpLKDmEZqriAH//EDXXCXwx
JCGf0fZ266B9FWrogSYeYpQtrsuUo98siW5JS4CzPqoc3rpv3XqPNwODl46zU4Dr
tsMc4KXqmh8cxEWGSHxui62VAvERFwQZ3N10sBFIUIIzC0rjr0jrrgROmd0wSxLI
JkscwimE04D/DhRJ79dPMqCQ+/h25hYMMXcyuwYW6o3AWnqySPCRylHbp8z+b972
dWwV0FgpBfhM2AUZiJZWvL5g9FNn2eTJ2ZTYcvuguIoOi0CSoDMl74XSG7iIvars
2beSKlAhu9OcXWaluAcMBZR2BPaNkajKBjNK6GGg+olGVjf2h0llH3eX7eeVAA+Q
Y4ADtE2nVvH/+5YrCB0hQQzQIF8GKqX5xM81KCarrgb8FuJ+OumdW8AsCy5ETMDY
s4VE6bfi01m3FN0uDhskvVNK5+7e53usdLQepSRhdlFG61IGTK7VSn2UvVREyxJA
H2eTxZFZG8sNSqo+y/xMeJ8PKGw0kKaiwUdssCasS2q5BIF/Z+Tis80SARCFxvQJ
xYFSzaL2ky0vvhruPGCKh8BgGB70VE2/dEM/ugNzOBNi2t/IAOnqYNCwGBhiQRy/
eqU/trlsRyMsgDZJBcqvZhoG1Q3iMIW+XQ//X90r4/McDdHbBxZqGCen0qF5r9IP
0qNqXuf87DcKgIEwOoh625VngyHaxL2AfsRlehQgOduFGWZOAklUm4WejHzMjEsD
VleIXnrT70bTJ11dh7x0exzvlKvsbbxLOuTR0KGYlD7Hb0VvaZeo30IRi13mnpcq
pj7/JFukZuwYuhsOZSxKQ2cEAs3yUNCEUwg5l0S30SFlO3q4D23TvX25Omun4ctQ
700t8sgRGIW1uwMhCfsnoX2iEyveotPe7cRYJhSrHLYalknK31Degoa9/zpYDLTD
3HNhQlaF+VIzIlebRRjclh0i+7I7aG9pJm/paCyJcL6ZwJ1Zj8ena21/wBEohyY5
JGy65G5gh6dmIZihBOgUmi4Z73bxO37p/yI4LpVacYqLM5SOTUJzYmz7jK9BkwDK
UeMbQUAjDBqbQnnV7mndodZ/x6KBAhmsZSiOBojDz/NAQCm4709ofkvRDp6MrQk6
e3f6k8mtp64ga3WlnxLA0KTKP2S2S+lNUi+/y5JadRS5TJuk2Z1c3XXG0pkofn/3
9uJuemAqDhDJRcYyVrrMt30dl1lJCzu++6mBvYiCZutBNz8g6N+kC2ZjqxkDgdQV
jwAB/Vq3/4bcbOuFg1RQPX+baLoxOWIfDr7N7fHhm6ljpk4vEpSTsdc49ZtEkQ2d
93AiCrZSztiybFpofj6Ncx3d8pFVDidmX8u7BQ6Tnw0G0o8katySqW68irmFUbgQ
9k4YvqVBlGhsX7yuocAIhXT8zc5rxFSVoPzXLZcke75/3JHTtbacyDTSKlte05Xk
9XItgGpVgMJdCZQX+PNJyU+qTkSnAqpCA/KNKRezGp+m9LfQJPrcgAGBTmnnRXx5
/fw9ikLAHFo83GMk6OANCPXJLtX7SVjQXwK8+FX3puMeFOu+A9LUT8+jIPhqtbLw
Zs6yuflRcmM8MVO2IwkiXey+fJllM0mnWENwB2O5dBlp74ET3kgyq7RSLKK1uigP
e7MuJDrCxkqFGs7Pj6PUVFN9hX5TYqoi7ynbcU2u4KiRRc8mLWLGoH50pDXBNFsd
YytCr+kPbcVtq/ajxEtmm5J4Auq8ZQ1pNyDBZBew465UTRn93EVAdMZeDoSJSdCA
njAXq01rkqJuJ+pmynZj9F2cKouPiTKbBmWIDfibURQRFo3e48cApqnKkVSSBQCS
1eQysaL8zURxK/hbAZ4P57/mbMGnP1D4OmDXIsGGBOijV1c/yFajnrsBId+DiV01
BnG8Cd0ZW8X7NtiVEujxRFVIlCS9jd2hFBTdIfU1JkvokdWMbphL+FkXI9d/7Vmc
fCb0vtob7/LxpWCWeiZ8PJtAxTOy6wmkAGaQTddHO1H5SEFPKQZDxCnKBAP9+jdm
yluZsf38qxfVdV541c1m221w/B37oIuO6Ag8OwPQlpPxXzqk1VZOEgQExc8d57NF
Vz1u9XHMLUz4NsLCCUpEg2hoYyt21Cme4Gyxxr+Fn+sI1TMvkNIsRpoQtsptmeb2
qdHsAXmXYqIjt5Lsvbp37rjJh0eaLb2Rg8cPSPyMZfX60paoCoVmMmfUM6aHd0nB
woXbKBqw0DpZkiJcucroIUI9kcSpqeeUlGLq9ZDBqdX87F72PLWDgCDU4a0gQ1vQ
1aFWIPdHrthWlI7hwSMfuBV+etbcjOE+h0Hjis9W67RfbnnMP0hsC5fsrJHohnWL
j1be1l/0+gZa/OgqcBzS5hS5Ad84MyYV2v9iBd8BADHeHBFJIYncjgceq4DldtsO
kZHfaMULRxfIsuk4NNqoj6UIWE4+p9ktToF8iRC/NgcwUZyx6F2ydbRH1n24fTKY
/9LMZkP++RV6Ju6zgqAjVNSIq5WXAxORtg+8GA1FdnE8zoEYNeI9bl20urN0wsEg
O1ZiyDr9pb78D9AsmFlUptsTtVKHAce34GcRFhlnrj1mguVU4hxkcp7bpMovkSG2
Po5JPUr69ZwvZN9eRzcl1U6DBx3WV0NKP3L3Go239pIh2Lo98TtOQvFI53OtHz/n
SI/SiebX+V4eQq/JG+P4t+yit5edacxXYrKcNJQK9bjeF/oCfz5rZFqgBWWgOEy9
kvAKeMCm2Kp2PWQU3KRluqhvmD8KFC0jrfMBfEJNGZbduMQHslhAVGE0uNd1NAOu
lB5moHkkwdOaWzRPHCE4oOtRSL2vkrhsHoqaxJD0CYsJGMWftC3muBWfeRV2suad
g+8jQ1dSC6XnVoz88E+s6sPkgjPCvPRXftokVsuia5nmZHaw+ZhGzGbJGv1gsa4P
/R25tJuIZ8hlUzGy713o6Bnl74pBSxyVtZ9XRMHj0MA2+CJVvW6tKyi/30rKJI8i
9S2Grp2X9nGlvVn2091SSFnNUfLUSPI+BnhsG4ffnD4qDW2tyEg7kUucJ9PVDSo2
+Mh3qBLqCQ2npq+/tMCH2HPlZDJh2f3Wt3kOt/JRshJtU+4quRypIxWKZnszvqlb
5XAwsva7DXHFjlB72Odw8lkQzpfzeUvb7yQosNkNn2GuQ1lqix95xd9hWDg+nVnG
7VgbtKB3F+8gBhTBSuPkRC7X4d7ur1c2VApucfwi+jHAvGmSSOIOdaFjOVW7Ar1F
VS+bh4m2M+CinMUTS1DzZBrUR6I+H77rNs6XYRXxVyd3LxvXwRKzz+9rtDz/G8Y3
CEiOKcbE//RKPiZErvVFCvs1nVoPMRVKRUlIDQTygN2Z79ND4JrMcC8jHHfo8Dav
ENxhybSJcUp47KpYkkkdZ3h0biWm4F+iCe3QSESv2Rt5+nZaNsAJFArlRrR2H/mA
JQkOX6WskhJa+bNZTpH3veJMtFd6mcJ1N46dgkhDjIUVt1ojGctebCpEyNMxk4qt
83zKl3o3tgGG2+3iPvi/BGb9qDg652+3zzYgjZ5TfgKlhptwhV9n7SK1rSlrEu0c
1e39GXYTbzaDsEjHenb8wBPrXzB/CDldYEmgY8PHF59KnVRBEviQoxBPq35uKRDl
FEO7/vkEW1AuDnNsJdRTav9bDKWLqpfYGj7XLQxVIhWd8+SgHzmpTgPAij1J7h9b
ahLkgvOu0rsmchlmy3n8xC7tyClPYTlxEU/K8G8IPoF40SkekhmaNfbwvW6hHTnz
NnpiE3o3CqvDZNFbcw5gqWUqaxJPcNKOoj0kXGcLSFTgKr9PIl/bhX3YwtghAg2O
/tGKf8OOh+jrJE1J8boP6nJkK+JKCfppAJMpn7w6T6WzN4ZNXw0zrNlhBGo3K5Vu
2suygHuO/poWvgs+YcHdGg4W3+N6vKihzf4Rl4NYo8CPBHCEIhLmyQoUKbMY4+sR
2eFkER5hismT5ddI0nzRUyRsNQVUBDzuGoANaenGAEE7RJhpKGJnxt05ohKjCvSF
Ku33ZzKJzECrCqVjUf7IPEhg3vWEtnlI+DTSWonPRna5EdawpoAUxKHGBgUofdVG
a+KFzUd2CSBXJrOCGRQCpmsT70nH7tJOzvHY4s0j75sfUSQX1IktGQA/S+ij4njl
WWGPsUqKTJSNcrKAoNNeuR/Ly2+zfbNGrlY6UuA5GFJ3Vxtp8OU6/KioZnJKPtN0
53iezpbVXVWzdxpwnlYKjPdIdqjiBg8LzsTHHeyya95J62TblldLzZpyXJoYwqgx
PFwz+ElFG+ZZ8Cjktv57RR8fOe3dn6lS573gyO+twzsyAp5S7Y05RjKe0ebOmTXQ
nahF8Yuo6qHVyC/mspUeILQKGb2iQj5seZytoqun0+EsQQ4VHzbkU2Upf8vCu/9H
r0FD4fyub6YMPez6WUhZnvCW5TU3cOoshPru0wlkI08SEL0lyToVk+GXGeOPMdVf
Ll6pvzAGdWzr2A1gqNVb7TA4XoNTkqNbVzM+vd5i1rf6YIBHSUvyESnZSFhw5Ot6
YVdLmMEGbeszVrJ33WvmRcQ4e/MKPUUMg9Bq8EXNXR9JSU7jcbP8WnhV/9QfI77P
PrnogQOcAiWuAji5O3HV6epcLTLODo0LXovvkPH3G31A7ttWiNjK/6iRSWvqZ8Gc
fFEaK8Qqh6tNJDIe0iZlLedfTXikVdjg1oK//WRMjVoL9Wozsnlq1aBHS27zvkH+
k3uOP202bV4te9GQNFwJRAYhp+DUbIYeXSBLSlTod0XemV8l06mJJG1A5jMYd08u
BbaVvh87cI7tvUjQZn5nGHiSuvTo1ByJZBWxZlyshrQEF3U5qCHcQci3DWvuUh9i
J11lISkBRAhMt5rrh1lZNXTtzHrjLqzCRIzTpLEzR4pVVCeQDZCu38hznIvfMBq7
hIiJy1yKv1BXwLdrWUMhg+8JUtGRhBctCp+8RUPeCCC6tRKB1HJvP9BSh3v2J/3A
8cn4pDGvx9eCzhpwa7lUJds8qThE7th9zsxc1qf96EyQZos/XJNj4lP374wJR0Ol
mqC1zRPPdEZMbpegpfVUILe2tOB21hhiF0KOcX1XSDScLblawEr1e8F71WAbA4T1
v5l0oZGsZKPH7Hl3lD7JYS9oTRyWOKL4P9RBbzKn7dk/hWwbd93EKYBPjvZakQNb
tUCuI1lkGT4fRiyE2KNrmJNiDF5dhXkqZSkbmjhbZOwEnOF8TjYMSP3S8je/LvDN
+qU9+xr3Fl1cOlkRr2mCqVpeUNepYxO/u9z0Pbtpb3KrT2CnHAko2L53T5ggQ9zX
0kSfRF5JqxI2+D299UhbbeLQ6bO6iOAv/J/U/7gF96NppswnYHCEG0N+HJX61RWy
dhUd+EDviEpgtUpG/WRqQnwZO7hqMg70QxAjXP7jTQaeXHi26NWA5LN2GP1h58Vu
ndPPclV+HW7aoC81HnrrqDq0c+ltixYM3CV5MDjBp69O3u8Amxra7uE7HfJ6mMIq
1GnpR9cYINtgMAPf/9FicV6SzPfOK1OnQa87fp7EEGMtYCZWj3wjXsksqDImTlTV
BQo0dYu+zqmUoUaKxt1M8guUm7aNRRCKY+Z18I2QVfpGo50vB8d5BYqt1dy/EHJO
HrI1BofkmV+zXTfO3IIcVRMe+jfXTkJzAV7Qh3SHmwLVUIK3mLxT8RqiSe51t9dN
zpPek7UPS12/1JQqswSHfxYz2qWbN670G7+ZLZLP83cg/8SfASDwbHtou0AkbqW2
bh3U5oHq1FFpe9RPhpkzrUol0QL9NibF2lTgzW1dLgUo1J3CloMtEEt4itoDdhui
2dmAFsCH5HeyjM2aSREUTKH0yLwbZi2UzKFno6jCP1ZXgFUcQHYYzWVturuUM54i
92o9+BdHxXvAfxrvicFZY0iddmHBCeAwWmkhiAPqW/NkACVQ1eYcoi/BtTlIMgpE
6lftg8OUSkYylvuZooJI9OBfE8DYP4AGa/ZweveR+Cg6J9XLb4ZCdFNkmQSoTSGU
6n4+dYQQQ4Z9WfSRCoUCUPzSVy1m8zPuAcIT+4xbRoMyXrgm01vskdDtE47cEvW3
bvmORrTxtMUI/3ka6EpY98gZGjWVnIwjq9KSkfts9UD4mtfupHYtQ1MwETjl7blg
/Ov5DuUST49wgygjtGrYy7mNXIrqoH6WvkjH50YaeWcwuagEJg45kMrBHlwHHb9z
nJgTT+c7AYvq7jxbfqklNOSI/a/uJgZsRuOqwoG2ZNfu0bV9hJx7p1BkBgJ1z+ns
JggDIEEqG6mGlr23GvA7IA9T1r4OKuhcdUf0jlyG3xt45ZiK2uNO/PbDUQLzqC5q
ItjKCkROhwOCCqzyfNrDWnhEmmHMEj2mHAqFKdSNKY72dbPe8hURdO8Evko2Q42j
SA7RhDQfZBk832O6XcgT3GMqaeXUsWuTEZJHMmJardLvj0jKQlKobrL4iep3eplD
dzpQc7g0duYJX5W1u2lLPur9KRdGTNOdvvtFnJgJ2l3uq7FYveSQ3iEqzgVdN+kX
d+otXgC3DZloBjDcR7KOBXslfx7z4O34aO8m+J7OIUCfuyo8Kw1M2TBsq/xkR34O
1lphvkWaPgVOygSTEEj1w4IEqPM+RNPF8Mwgj6/DCaI0FSfFSzIDx/3V3/Z9lIOu
huMAjH9OsEe+OWfjLOeoM8KUAaX+P6WhTj3fBvuoaSyI8ZF4Kxz37YJtxAF5jrpt
ZkfCyFRmh/TOLrRIcvTlztrRJYI+XmSvdB5h5JYVEng6uOjLqcu9QBPElGvaGDZY
R2Jp/KYwsk20wtckuMLcaTUmBEw3BYoIZp0RAqbHIIYFYWvyH63yZjxr5csrUEPY
hBEpr+IWhdvmhWGx+jpW/mOs8UiCa0flb2sQWVka4p69//Gs5sclQXw8PHI1jUVL
YrWHYt+0S0Sy8FJ2nI7LBogU0FuUwqsxBDLYMH9h2m5CJmhZ+ziiuxfnmwRcuYTu
puGw7+5vbYLpPdiDjVr4EMhbM++h+kSrzpJPdSUhEY2PEk835+AphZLAHy6YpRVm
UZMFRzZ+IxQ6A4k3QZvp5jgkOLb/taHakIiF/ushdPGEpJ5l9gNoP+4Z1GCKagIG
tHgNiTx4/KrRvgOkM0Lxo/wUQg/EATvXArmOiZvWGC4Bs0iQoXN6rwmVbjd4Pq5Q
jF5iD7v0upe1hf1UIryvNmH7kAZ/foaflUB+GLr4fDaAkfkMZlXE7qaDtj8K2b9/
V51rfVRtaAGNiu54bSPy1o+MwTlG/xbwkd1jCznwDO7mji/kjzwDYHwRDVdxDFlA
jsn+S9D4ao4p3m9ZF3/t0EalvQgNfxD9zwHP5JojqydE2gHfL04fiZQ7WmX60+JO
JhhN+5haLpsrRAWrqYZ6XMg7qxkje5YA/ngzkzjsOYw7hDFbYCX86ZgtRKltiVt5
qsDkP1sG7rYhUYMf4j7tixSeC3jp/dw2fUVl7sODwbx1wJNQeus5ohalivfr065j
nMgX2RfkDkRlFvoOk0I/Q/6rT/PGJM5nYc0fScEboom2Zsmf/c7ye1w8DCjJBYkI
fvhL5cT9f2Louv2C7C+R0rDTDTvfkjwObcn6StiqAjCXjXvnJqC5O+q9OMmHgiYM
ry/SB7hnE1k7g3aUSB/LFp4eVHxj3LBgaaC+19ks5bO/67uI0XSztsp2AsyUa02V
D8FAksceZXlmnAyv1aUSIYk1wqjuLKqHWbGji8JXquoTSq/v/TDj0HFitqDYK+mh
O5S8CerKjHR2I8tNmWEXkHnYWfTCSSvAKIlyvgWHt6uiOJFX8NHqBnK7m2fT/0Fq
MYhI+ZFiieis1evlZqg7mK1P6l5QrGvEe97d6MJvWRtL0XuZEAvQ9xUKJVkEot7H
eLlEYk+PDeH4kWFuNcwwB7F4HH7ukyIJ7R3Hd7Gmjr30sEyfZlFpHGpqXcw6O4Jr
lS0l73IK3B35qusLk/0R880cBTGn54Mrr6tyPk0+UHmWDZh/8P7B94XoNc8AG9Od
P5wXCjzKZxg+P1N7X22qs0yGrchSST4JA5i7M9UaPOTfaXkTVVuNCgXzXKiuuv/F
OREQFxv6OBSvU8+XGvqfqHsQ0QGW60/bmGH2Zy2KpunYXmh6/q4NGjDrkUwz3wxf
IZmGceocg3uItQdZcBxgpbqVfONuG/e+pu1wUDC4vyZCxhN03M9ALxNnlc8iDPOi
yEhekUxfn6HLZPFs5L+Su6DTIBgcbrYKizyR9f+X/bJKu0g/npOt+8JHMQh+D0db
EKQGp0ruILl9U8SxgVKowDPKK69IXqMauiE9/UaATSZ94cuh/bMmIq6xc0ias2BB
M3XCcMIk5DrvplsnG8BFJV4g74/N335O8Rx227iswk35EyQkdzJNYT60pbZKd+TV
hTLfV48CJn/XmnDU4FMAOkIaVMQ4nNIkJ/bj6iH4DPkzmaQn1kASpL3y2d+rdvhX
O2CBw8koWfrYlL8MWhzBsSjMYsSyRutmYudQFEodbwb2OcWwKzqgm9B3LLAf3rCd
JvHOZQQVGdL+eW5K0/GxEHdMxjb56NPos62sAI+x0V6xjBZgnKHmdFRX++189Vqt
wGJ6F1PPNtDCOANJLz22xJvrrP2ADXBBkqO2eTfD71cBFO6IFk4Y8r6BSMMeJoER
xRlzuuftfpQIOk4ex1Km+klsFy9dC1PANRcDO+zkKGB8BwdDLx+8QfGzu/dQvD9j
6RfxAUncGaXhrZlR1jxQy5KV+TPiJdCsxazx5hAUYnDqazuxPhtHrg7GGpsavSeE
/y1hAq88w4BTag4+ZFlgLfp3bRQIUPLBq9KI3eGGx9GFCqjOlOrMlEfO6QA6En4/
oPH1YrY+mMunMRk3BM7LcqnhkD7jHSc4VpcLVEQiaeadmpbSLDgy9OzI/qFovYUa
Ry2aGQxa8pZuyLWDbEVgg/rD2/scSBOALyqFnzMLHR89Y8T1+kr5xyAE0cTTCRrF
16rSd4u5JNsG/vGuYZHt1bdtmYeGgrgbeRQS0Y4bbELIbySlbMn705NJJbcsz+Ve
IX2mveliK3llqEXAHOyqRak7CMC9oqfri9EMxgbUSs+WIJQsYyIkfmZJf1bKV8c4
76YCQCh5/UNduZZB1fgeUE8QrsrB6Sdp9hl21G1HBazVpS4pAMRmSCFPr+t4R9Fd
OyPQGtflre14m537VJUYlfM9tOkHzcndWLY1wfd1CfCXX7jbGKr4V9StxzI5ySah
oXllZxiDoV7RnZFsE2T4sbTrbwkxmt4L6vDTdFuZsNCbykaT8Uyta81DtLh2M5BV
3Ctgje67yAHvHtig0X4MS+VMUMufkGwit/6eazmpm6grsAJjpzHWXCEs1bj9yXJd
7XL/BmqR4S2DZDl2+MHgPaA9YqjEj5i8uwBzNdCSnRZf4grIfykxA7zdhlTMbBNr
EJ8Z+mdEu/m7YyETHFwj3xSmaejKUbphVfo3HQY66tuDWpk30ySmX3c6Q8GgAOen
l1layjJmD0n4vkbncKYitPonUkn1jdGeIyr/QhGsuqsVgMipSP3jETrG5MtDWrUI
0fPB134WhquWiCC4vvligC8Ch7h7k/35h7K4Mn+SHH7BrO6zo848rd44ro8rfUec
YNQ36FkdevgmGvnpoDjIOAJXFJ5HLBM4wmWkZedRQYjFFAxUWdx2Ra010HeYSrse
dVR0lFU/QI5l2nsfZVVHZBoOkrRYJ0pG9J34T9npP6fsz89UAcxc7NEB50/3IZMF
6wtUurgjYV13muQdR/JzTyMi3oGytZgb4E9ji/n2Bt6RA+zwOC/5N/4vmpIjKFXZ
lzziMJh8zSdcvot020EQU4iJ78lX4L6Su8ri8vkNq8ODR7Mn239FGlhdq8ot+WnK
UqpHQWuf+xVfbIN27LWCaQs4A8raigce4JaNnmu0dFMVTTnqpMYsiVoUv5zTzPtU
8wc77w/n+wQUcWgXQr41rcN0SWZDFVojWERhfkmevcu1fkYkr/5MekfFSSzP3MyD
q33b0u/5koZYlnOyBtRcy9iO3vCY8hLnGpx+YAYCFSsOA5z11YwYzOu/bI72nLLF
9jT5Q/zA/IXMcgUVf5cwCHQD1mVHNwE6hS6Bc4biWbuEVlnyejTOKCT8ykW9JSmT
GgV9Lz15qdZWs4FpHzuVm5urg3m02PF4JpylTNoo8BbUi+GZiPnIbp+AVvfCKbPt
2bPWjnxsua3QBmIH7Y+QoQUaEZhKVXSlBqps+tapX0qRIwW7JMl05CKI+oBmo067
iyR60gjlRZ5SSPrQx+1YPq52nB9UGji14EF17cptwrWoNI34xO2Xm3sL/HsLHGDq
0Rb/DYTnRaCExylH9EksI1PL4XJx9jnTQFcdqz/8yIaLTVO5Yp2H+YPWYgWr+0nx
UBE7ukkyBKeKeRpamtVqOp2VoCK2sMJEM2eLwl5DT0PvgogRhuz/s0TmHTu68oLR
yE+eD8T1tNXjhuG81AUfWDMnHbkr8G8iMdCMz+y/zoMQFIXJRpDTov0EV7L1Aree
FBoDUvwtTaKgjxFJHvvct2aikwNRgzfBgMifHrSYvqaLT/AzoyTxT2Fi6CRRKI64
Vw2ffadLQMwrHDxD7Ul/HlEouY+2PrUGiVoh3HS9P/UW8DZsEzf9AW4PgPgakQbd
ZJqQk8kPdAXtLqtBx4P3jsUaiajLDxY9ZQpmQ4LHlCOYMRoXRP0odnDH0oqjq/LQ
UEcwh96hdQN7jFBBJ7x6ygbQ+yFVc5UWXaLD8cimod9On++tRP8RMpVOv+wuwYFL
TxTihcNfO6dW6l3BcEkV9ZpjVqGLuxSmeO0XLS2ohUfqimBmBPU22s65DaApm/PH
zjiTx1mlbApM1mVPMBdzQDOa4zuAwkM+7Pe2rhrTP2eoZF4VcqgjoYRrICDrSiV6
aTGc4co062sSPgf149HPnzHwXi5BIWJaX8I+zTxUQ4GYrrDqCroD5hcM16t7MIS9
/tkFc7XnYsY6vnbAaZk34T1Aip5wkLKb2ehv4jyVVcgRz+l2rNYFDk4f5IwGLHiJ
ygWtipLyv/dT7NXasU8PuTxt9MeNsTBRogcrUdfNW/h8xfuHlvg3kfHGptzdGRwG
uhcovcDwEcDgwSJhxzjqiEvgit3Dt85aG82bxalgXLlQjNUvvTjPmPXFjWDNwczq
i4VXbdjxQrWBjt4xjLE27ga6mCYXuB0dPnzItN/wjb3PB9Pd6T91tiIKhCpm+MrJ
l98nMLs2rmMUGlMoTxPn7hBrpdefxE3GoUSZ61n5aqRS2FRUd3Ugp50coVsQgjbA
FvrCP0h6hAyFQx+Le+GtG3CHZxKuOOqSFQE/O6j7yzRo4opFv9sF1oMkLKATvuKf
WWJy84C4DVWJCWWiMj1ZcmjIJ0wYkATgfXdLsNaoLMwzUWA0/niW377bJWzP7Bv6
Z8FfQLMgxTsfNKElVu7YYA3wOEEdFOF9bn/EjJYno48N5n/PDBAkQV1u1o1uIzzc
T5YSpIYjk52uu0qCZDE8UcfgK5s29WlN/0n6NRWJiQspqDXOjnVbG0dS3OchMXiu
koYIFNuiGs3PhQGh5sdIpjDm2ndTpzaYgX4JR040yOpQogdY0K/yFEifi3ygDg4W
w+LjrcHau96RGv0LQ/lX5yW6p2hhenshecDMEpEsQn/GcPBlrG/aRKvFkxJYIOqQ
HFzrf35c56gsYNKqq+Dpf9d/8BV7rBPT6lAIp5WwTY1+4VDHcMjHemQaEXedFleL
OJ8oKyLPNblz+6uOHCMLz2VWVlam+RQZ1wdz/V+urF4d59TjHWLvhzcPMk+dEx0l
ZzwmKaIH7dC/9QgSUY+bJWosLMA8rhrwYc2WmK6vOCr/9+hYzXIeX3ByKwUGg01C
/uvJ3z4CE/psAiEOw+6F+lQfqkazpKcmSRBc7viYLNhUt0l3i7Qmoq61aX6hgtd4
RowdbNWzHptT3q2DwDrreMsFgk9GBLlmAt/mmxCbdMVnS4cL/+K/sVcjjf58VSPW
7YWSD4pxvOk5+eZEwOhCCS+U5CMGaHCMNs61qV7LauOVuByifyMfxXWIinwqs0wj
WlHcQ3+zJJmbxYk8Fjp4+HAIy5XYrja1qRLnNeYTFREWTbKkIZkyDBeLZT7cTy7c
UAUGEs+86DP36kGJWYoaXwnmNJhIwyqcnQocd2Kek6JIYeJbse6qA7b2XIiOaXU+
VzfKSocI59LblrQLI2nO3UYkDu7B/Sr0hHpOp07aQbA/swpfoXAAmz2IFTWA2MXW
ZfGUpbUA0DIva1BuRIBBsAGaLe0UXFQOa7WgjSJooWAUXNvryJKChAedEUgACui7
HZ1VpAzSzsQ0vcb972xNmXISP7ssnC+0eaJZgIUBncOrG25I/bDyZGIulJlCw3RF
NP9deeI/FdeBLmp7wSn46g==
`pragma protect end_protected        
      
`pragma protect begin_protected        
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RHXGidM2k36dMIe6asWaiyb6VxyqBO5CRC+WfBEILt8TlfUj0YBBiLIG6XNMyiMz
ZBFBNwwNwHO/vZsxpmbx6cKyn9C+CpXgmwc4GklIOunywyABXsRR3HWpgEzSxunf
okaT9tGUhkGX/yEvt98mOvqxbtmXPONdxEqWsAr9+Ac=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 12203     )
wBbfy+ONIXv8a69H7lqXlzIYf0W97noSvF7zCy0N39EiYVttLinz7CuYRrMebZ7u
eSXMOIAbmbvNVXq21oYEv9ny2kYZ6IXlflwLZVBVehMShy6gCs3jibJPgQ9bgWNi
1ZM79bYSzn9YmXE9IfhQ/8RQZXRWW6gccR87PAPZjgeFSWHzEN4Ij2HTaJD2etDT
wIM6d1rJTVJr1R2bNSKtzwkGr8JYA+pPxwz/TrTsjhy1mvbwJ4pN56j6SgTnfrc8
UQh1+HEqchw5KaV0DXmFsw==
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
KssqzebvG/1YEB8KOc10cWUi/io2hyB9Z3gY4/w/rHCaMxeMx16HCOw9Y0LE5xMo
BgloTzcvZ9XdY3ElWF5Grwm6h4v3MkFCbHx62wvez/F8JRnPyhFuS4LztRWPB7NT
FewazHrKIldbvrf9gMK/u+QwN1TuUe4DFssRyYi8cgs=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 19866     )
X4KGhZHoFS70NgGbgFc5k+nJ5b7FO5lgPAqmSXjhgJp+IjTEDWuzDMHdGI61rs6w
srqJ06IoHgMhLhdwtPWsH1FZRGz5Ihm2zS50iW+DsxuyAf+6AohIF8sbmXArm06G
DhoVePJnR8TbCzat4dhIMsMpNZnEmFxdwJuaaqIUDEzaKzFmy7yn2KjE0piMxVJr
Xy8JISDWQ/yUfpIPKCV00VOaEA75LfAO1YdCpR6dVszatbW4NIRQnu0nJvxqPByK
h9fyz5eCSkZsEYzZPQbB6BUD9/jERk10e5FbbeF0iGPsxEggDOzF5/appVsZe8xf
IYymMSUGp77rtIYZ5uM2AzOt00uQ8ea2V91p1ogTpU4UQHOwhapEw27+F2S/mzCY
TfGMC4L+PQRyN2yciO6B3rmZaeI/D558IiGan+CB0exSSQb00DNaIJf+Aqzf6GWf
9qfiORGgn5QIF/WWlNv+jaSkguDoaFY8L+mlPmR8vgLlh/vCp/iowCEykH4rwjh4
IjMgKpnYrasWHkJ84uRrsGKifoRiFtom9jw1TlXkQYc4p0Wl6JGq1f31NFRH62uy
eutBZkM0LvRf/NgG0GyRvqk62ZVpxUpeiknrNXlXVJRh7TBjIeaXudn+aS4/2z2c
gsr5s+jMn/vZ7Sh37JGfuItzusV8Bmcn/XOcyPUyJ+jcVIVU7/XvkofIz5gexVhN
osN8HY5CGpLAVxWA7UoTJCQ/q15Mo3bLjFamD4NegysDHggCyVVX0DVWhEWnq1U4
IGZIac4OMEgQBpY6FpSNQfsNnCi3Cd1YJm+vuR8Q06yz0oJYF8c+8qMZNtcW7B9p
rP/SLzyYMka9Ar7O6v7v5qynOqXZMQhe9qxgffoks2+1MCQiJUl8FokK7FCb/2H8
mv/LatF5quu7eB8pWZLv0a4+nmRl1wBCCfirDvnjQADghpbYwHQ0sWb1OFF40CPe
yX8UWQXk5ONSC0AH1TWUMxcSFArXFqJH6TseRMpZP2aGkgA0pV3CgIdUvUWaPLHf
Lru6NMU2nVEUmXi0HTGM3xM58v6BD6DuSoX6OGjoS2vtzVYoF1wc25KLcnpf5Xe5
BYaBbQLoZJNMar8hzADi5hfDV4ixJ6EKbIMYGDbdd7EP5dkFPDPx77C2Vgb17N0A
tr1iCThHP4umvOLfhU9D7k1diH9GPjlObg5bRuZX8RdYeL6vAUa/XKE9J0ryc8Sc
FNik/qRI1e2FdrLHBsrPfgkVp2UqCMSLygdObOmWVQpWMX/WjS8i7cA3FzTp34SS
TK8TIXLCnj7tMpr/lmnvzZUlyQJE+Xg5B529Aw8DReo40IZVe5xLsU5fwKdAqE+a
XUxXDsCWZP7WKzBFFE+VBSKhXt3N1sb26HVWp+sTugwbrmf4g2HM8K6C2kpe/FSa
FL5RY9/4ifXhHFXhLXY5nj3wDK1d1J3bg8Iy8pRcbCYaAr9p93IjnSPrSK5H1BNI
kkTgcHAyMb77vbzDWQCXxArSvsR/3LlzTqNirYutP8wCxwoHl9liyEutXJoi7b/e
2tXo8FRwV3GFK8i2qRNQmdn5yoOtr0u9EtFFUKZt0Fw1VUy2L0zUVNyvXsP4SdIo
t516mT5fHUf2GHKui+vyHeERlooGV5yZQFXfG8/wY7K0ctwZT4YEKomkwNAh4HK7
aPVi6fQeJ+8NuUn1mwMF+L0vTQRyKzJWToMbOe/BLywzNqrcLJ74QOk5w82XGNI7
wk28XIzyd3Pxx9qJCK+yHNHh7GQinUHnNcxoBkc3paTiqxZntzRWzPCxNEv+ZX8X
QI0xuNC1XddvB7zkUjAq6P9kr3+I4LM43cGxEGc0crXMReWE4IoYH4puHSJJN0ah
ymekFpJku7qwp0oWqF0Z4twtV/Ppit8bW/to3rHRVXrBQ1O62xmI4uEJJbh6TIot
dq2bX0ZOKDkCnWEavNvQ+HOAJehvodtKDYdmNClOZmhQpdTnXuK8zZSaDHBFIr+z
S873KdOCwLlPsSubw669vYITgP/2othlPDHl2QfZxpCRdXZX3u38lb2mv3xe/e08
hbRWWJkA7ilb8LL9lf97VCytr/bsVdXiv19pCfX17YU4EOAcKDn04o9UdZu5dvqk
e+mZaOZVBrooAoY3cjDRsgxWnwpi2LDWdsHKgMcUnsWJdtynvpiJ/KxdFfOQmugN
loHlBBWE47YdPKJHOGjMdxEcY4rb76LpOuZ0WxyU79C60wpCXaiV9poYWvoXdfj/
Rll8/tmcRfF6NcCiIhaYZQ0u2p2wV+43PCbVKDvrlTaEsOeH+tgFxeLThjVh9Bnb
mIN/Gh3rskaVsMEg93zEBO0haVdv/cMt9fllWYtm1R2ZVCn1bbhu/L8P8Bm7I8wx
VTGJqDmVYvhAcOa/UdkiiTqZDcDNBV9vzRqPmpjFuQJglBTLDBzArAXP7edinCn9
sMR23bF5dl1+AOpVswo47fewaQ6CeGMqkzGfa0/v3YfAXo+H8rVjRoly4YImU4LB
qfR2Ybr8nbkZtFqzZV7QdKiUcGrNCGeQciMe0YbKeoowuytOj7UMSSDpna011o0I
tDTsVCi8KvQmSWiKHFs6YGwf9vj9U2cBt4ub5glBbmgMDp3FKFnBIzuhZFk2gS0K
ICFeXUKprCHbJSEJIggnmeiLkh4aWz+KEazKfoc0wKE2Tx6JExvsAG697nevYDsj
WUhcrnCcVKqNFoWMgWfAExrmlkaw/Q7BPeQgxmqPpGUuPd2ERMbFIpdmIH5jBcyy
fn4S4TX13cXHD7wMFXAqBjl8n7jwT8Oq0bW1G9oURUltjw4tCHdu4W4NCeZv8cQn
pAhtFs2eXGHTN+oSnH2qtuRiv/tmT63IDK47IIrVQViaNb7V7TtlHwpTuoYUUvGv
adi/tYSnECH1jADA80TkxXPe8F3JDQwHeDCY2lzQaRh95P5zY7CNu3zBnd7fhe4J
MraLvnwa6HyaHmnM9gmzKrkFrzyisoq7R9ZpIaduCRaZD4ReWAiH2itUrsgwrlzr
8U4GuHcLohiLcBX5lhhbSGpf+U3vp+AtqOCD3M3nhJfHL2qeIAOwnIBGXz8rTCZB
K83voK0M/FcwiI9mM9Ob+X7HH9L/p6dSKiG08808u5lAuO3Nq0zfx4k6TwKhhLCy
QLMM+vBHFm7t6Z+Jy1nHSQ/U12Rkk9Fa/IwNqBFA0ud42CNqKUp6qSa9Ym5wUC5+
5rztzRcZrW1ueNcHIUn8MzJPN4z804cxHaZ3u0z4+w+9UkKQ8+ll0AoGoI0tuivM
bWe/V7Tl6OSD3WggXp4bE9WmCTL+U2kb+3k64dcgrVDLQzqKQBiSKb142QubraL+
aiclQt42DtoUQ74k1zBnsX9PlDeHxMgZ5/sCJXJ7jlOcPWBH8pk/9UuhyxGqd7Xd
PPaA0AYnV2r4oLUxbuuCtGW86f3uVyu/cceeIksmQHAYpj0DIwtxfRlZfRDzx+Zm
fLvSSmzNe80svIq6/zTa6OyaccX+eo6Op25SNalFESrUhz/Z+J13EF9jq5NdxIX6
amfMApLM3Ju1039dPlA/ZPesKr5BukrQYj5dMQxh/tc/zJU2HfsRK53cfiAxy+Ds
mf7G4YjITNDegJyMIq0vJNjCEsPGPGXxVP2MwxP8Db1x5YmXk8NIubI2EF5V68BB
PIkiTEQRovJj0hMA5JgG+aFsRFr+aI04bZtiZJ++I4rGk7zxSJNxoRru2YxIhV6j
RVVyc493LNCE5TvXsh53B4Ci6HHz+0mgBpUoDwfpI685cX2cWMshLmMaTVpROJIq
9LrQVI7Ind0wL+ca7d2GWBxQeRtEkwAFyXDFp3/aGnWoFIQrzruuiQjZPZI6xjSF
t1pIS+uiJsp/srS5AwKyFhYrldyrjaU0Y9n9n78Xts01TlH5acd+62CD0pxNBoze
fP1P6Ups7n7hwstVtK47FT3ro5MHKeR6PAKSEIBeMbMZcvcL/qGGaAwhQTVXvJo3
3G4MpzjSiwQzlpwdSqRnBvsncsBfYb3Xiu1jfuJsBXfbdxAiIQv3W3GA7GXsDS7A
UGrEgN7u2SaaYCK+EfDEm/2TP7iMQXgekMjyXDaPTCn+9cfPqVAuEPpwKRTmC8N+
5/6gPGSWHhHp1aRLX1rhD5551ALFwsy/ZfE+gMtFtS43K9ubdJ30liU6EQIAP7tR
lBWGotdSKExEAiqXqYnm5fyhYKw80FGB8K2jzlXydhnKfKPyRKhQh1KHNpJkhOLr
KUEUjNV7ISOwqGxzdkt8YUm49dHa6y4E4nf7cUKMdcJaw272Nvhmwx60cOFoOlTU
T9cysbvLpYcOAUMa9Sw3poegrXU9szHH6B1OC01ScltfWiwaIwmjEHEsWzGBBul8
4Nqzb1QXOf+UVCM553IQ2/0vOvuPdlIz3pAVDNDNPzPfnC+/lQ+Yn7IkzxVwTMqk
Qp+3rfB8AASUJkW1w4jOKhmDB3i2ocvTbVYYlOl5+CQ4+wL3hLXiyhYvF/oLjaQB
pp/obMxSwky/yob8K5ClwI9G9AbgW4Inky1Huh5K8M86YT8ILDdkPFC/w7RrMRjJ
U3ZuvD7Zo8RGxy2zD+PwMC0Rjq+LSLfppVnMCI7uoZASuh2OklQN6Y41PV/uGRHP
HRj7xqz6OGlZBQdUyOTnZKSNQUpRob6u+qaiWcPauJfBqk/5WUqTHFOQuaCXQvQb
d9xcmwcG9c4fP4B3nXf4sykpq9Ck7dAMrYiAoh5LXMDh5u31i+jif3yIvev9OFVf
+I+L19ohkeDAuqsWbDyMOPtad+VJOJxWhuBWBPHb+Gx9xih4+dyyKgLZI6F1VtFr
YjQTDUajsE7HWeOhU7OkdqAFBqcwq1AAPCB6A3QE2W6W2mjm9mQ8PNSNtbhciiRQ
LR/ozuHaDOEbJvPprJyzQh36iufd1FCRZweLM0CGbZmRN50q9FfHRHdv38h3zRby
ESuefIqDKy2Dd7iy1sH65vUw1jBNU5xXKsbW7nrtn4eFeVVFRjX/kuJH6Hn/lUjJ
/NZcREYgQxWGiSJB6HTeEtAzPUQUnNodgFU0Fo/wYnYiFEjlbNkrOtb/hyw6Rqgo
d3PYVnGDEDfKHmTSq8BkjkHIlqM1c84emhTmhFc9FkaMZsdUXwQQkEfzMrqlo3fr
Y0TIkdavSiz4v6yB+Vu2qYGlnATzod1rTZbo7FGA5T1nEwHqXUgbrhrwVydg/0Kc
9Q+v6iAkw1162e4l7WvgyjIWN8NdF+Ay2/YZhvPdgF2Ry6NVjr0n64dgSpcKcAHn
ErZqWz0JamC8saICbHUYyU89g96+RhmOnL517zz4LyVUdOJTWhEqZysmbI3MU1p0
8JKVRS2lnbBIWq6/Wtq/zS7pGTycFEWMJQdyfY2uE2bEgyJ/p+LKMs9t6Dd0fUpJ
u9bJrHGloJvM2+j8q6xtI9k/GxlKNMdxZTqZBiOvqiwy64PtqNaAE+y8TnetOOiz
lsKOVnSE8iX61u9kaqG3GejgYX4FVclxwaAAffMo4Y0HY3xftLl0TzRjWL+swZtX
aBfXU0IfhNXHGcAfVihB7X6dGT6l1rFFJkpwUQsQpV2ggL2DBHDE4SebQ6Oj3mlw
a4C2RvHex64HkiXLz5JXBd5Eqe8O6FisN5n6nz1t89+f0B3JQdgL7B82rQIdK4EG
0kvSnZXGTuKgwnLv6iMXuouBRDpqjD2UC8HI52AxbO1+PdKWiqJ3EgBbHPqYONee
kO5IS6Zf8BwB6M8Q6wd5B9GpdCPQKMukU6OcXAUPJUTMbaq79DXmC8SQlnIwq5TE
dwCjcuddS4j3C8PyQ0osgzJOCGOr0LetFw1xhz2s1Ri1pvuOaJabtO0ukoq9q4Zl
Ha+MOwLmxjjkKzsfMuJl+edCJxLQmb4gnHcU9hUasxw1lMtLvDuzu9oHcyp5v6G4
8d9REdwJFtZePORPZTpnDH04WOgNSrz1Nq6iKDKpwcEs8n4q3LDXVSnJy0TQXfcH
aTQp4S2sWK91dZldGZLGumZvOaT4sI6AtRbeJg3qNg2ukXeMBU2mxssR96kWfN9f
L7+Omnm1pdip+BL8PynpuGhlBDu8CMVY/ieDuL4eZf2gtTGADjYsiFyGD34xZsZW
eojqY1q2iDtdIoNjEZy2RJIZtdEziGkF9ISlcQI8qb66EhpVkUzhzfNsmzv8gnco
NVDRECFzu7w1cmP9mbHaDX2Xgh5Gq+L3bAEOGcz7Y/Jej+S8itRvZ5/4+3U20ZMB
xF1YxC6qfA1Je6CeovDYyS0zybh8F+PyDzvWu8Ii//NPA2v/dR2QE2Lh26qPfAno
Ct1UhYYXmrn6ekiIv+arLbE89B+f5zbUeGnmTt0ushwNmv58mRgSvwSODg+vJfeZ
BMttZUVJF4LLdBPs951JwfAjURF1wtH5yzlv+O9rJG1qfsHF9In4fffr2A2biP52
943+AGOH3B06/qRJO5hO0SgVEvJvdkycdy6rru4SV/zVSErCMJplVQi//C7ehVf1
Pkau1DFJnXEQY9SluIy/dd1B40mYVS7Fzx8qt8gRZ0FmchU97QOMTvG7z9HNFQdW
ZbGESD4XQy5CSCicy48r3j9Z0RCSNHA1rmQlbEhL6s8qOqatQJ9e1SjKdNwhnPQi
cg/ycuJN3g5ziE4woHRUMKtvcjGiD+Vjxs5wSNeBKL4SnUJT/xkCILwETdA2WAXJ
2dKDh1tgsp0l8H5SjUV8LC87bh+3XPhl6X2Pmjw0xWhfLQexkhXbu00Ti330tkAX
sD25KnRMwDHyISUWZ6CL83QnM2+knKVw4zEWclfLuPU9wMjkI3/wkCNs8zPxh1cx
Nx7LqWey3sLIbOzNFyuEoaWh1uzbMnEbCfaAVbXiXaVKcuVJWYslgvoCa7P6MlY0
RzQLnmEG3ai6F1t0NBZZlwM8zQ18N5ObczwJP1hVBVY9eO/ptN+1+2oP44RNJv/6
p3ZFxfUKEM8S0zmsYjbv7TwWD42oh3BNPBqiTmE+z00A4q3XE4G9JdVvs2VU63Bj
nYSRnbL4bRX5ZGaE2x8+R1iIWsPGUPX3wIPzstL0Bu4n4Wm8XdNKUxcTXZ2jxcSc
kzMVq2NSJ+s7c8UYxwmF/da3R9WdbRqUFKcP2RNs6h92nbJRw2iSs9sl1On9P2jv
DJqDxPJkYH7K0hWa+imPY2JFtj9wQXgRUlPTfDdb0RrgHPrVdvLRz1C85UWfmx4N
OiD3kAguqggFiEKUor40kSwBw/4eS+Vj9ZNWOh3opEdRL78jhGZ8xDDHr2PVaDIg
bsVgoBDAW0rb+LDAatnIFSRMfZB7eGxgdMwjmagM1Od5khTe4ex0SX01V7ZQ9kCk
iX56xO/99tZffLKuQHTOlo+d6blZV1KnTB9Y5LM5ker85QgYQPQp50QlAKbN6DC+
G8HTvwcpbAHvW22tlqPgza+PyCj61HXzDVgzWj/sh2bURKJvsgWnuA9CXNuCFOs3
I5yry2SwvoJFsm5GdhEzm4MTC95PHgjeNPKqkqaLPXPaSbta8XCdcs8qtcY4ieH4
2kKWkuDDySUYS5W3spna4l4ZiKLqk9wialoPGFUJhUCfUIlhVI+KJcgrANzj5YyO
BS/X8SsrCU8Aqw8t7jhVk0OLUAQbM5uEthzcfoamT5P8W8iMs+q4IEA6uRun9CWg
+TWUDFzrSWoL0cBZH+9U1i96VHcXDJRPFpJwynEUary/LhIgLwOwDZcKF5UI/CKt
oK7aVo26GqxYXu2R+feejPTakMnK3Xk/m8Dm1b1skNfTOTOWi5ApNPEB0g3aKyvk
Ro5dcRqnKZQZ8rPUIh3NzE9pFHh61RQTxUB0DIOJhQrO8kTzX/mcI7Hhu2Pvzbcv
xpRQ/lUfYzP4OSAUm8srXZgu4avTpWulvrHavgPrR8Yk2ppSvu/K9my+NCIzt14d
Betkrj2kpvXwbQArL5ud0qccSyioqQRn1AszFp5ULwLAvFAoJq2l/9V4oLGBKpzR
p1xNV6xc9WLXFLQ68PDbPJi8LAwYh+XPGxKJAtTLv25ycLpqTOHz2rb4gUIIHgUN
sxELnyjjEz6wkXf7qE+8kFK5/TEz8oIk9nCQPdxVV98P9SraKtMgQ8tjQq0Sy8ze
HOIzATRoAyL7f385nIEYF7wfckzCVjezuiCXx26Ti8Lch3Z5dmZsP41k58cSNbl/
0uMLt0i0qN4H2ABQ0HseGVlzhYhwyfYO37/XzyOYfy3wWev7CWj7RJdXPf7lD8C9
9xs1BiuH1V9E/p2F9axlVNJ13FkSXGz1tKcrqqrvB/l+7N681ZoiCWd3OH6wAyeA
BSTdGE8UrN1U+83ldewRFUxs+wo1Cdg+m5i7NV0m0sVgS/dvxxHFjO+BFI8OELJr
gcYpBmiXT9EWiKjvkw0VCByVaaE2pTARi9SPtPBFNKxZEifE1+xkZnVVovcBa5Nj
rKmV70+7B38hgDNrSxc977RXJH1SMjhSMHKKDZSbvb+zUmHf2iIMdVT4CWzUZEVK
R1KtRbXW38I3lkOD5zlYS6EkrSvTGp9rpkIrEsxljmJGQxYXXICfloaS/pz1G7al
IzqTwxW56p1Scd7dD7jtrNG4e28BvdBrCykdiHqn6V5bhy5PFgdQ821X92KGnfXy
J917nMjFE1NUCOcZ0gKlUWe6AkOwq0RL08r7WHdbVsZf0LT2JexiKrg7nTMiNA5D
hNA+1biTuUML1sGF26wQqprKjOrE0RRf1Rh+ig4mD0zLPQmo7Rt9r7DKYaS/eJDP
s++/62NfNftXmJAIbBcy6qgvMui56ZZ6oXiK8EAJNEVRNFQoTJXC64PUt7tptfF3
WQb+3f2/Y/7d6ZwOy8H5tuBnTUAQlK3BexsUmdOq2T9xlYM64M0Q3/EtxSSnNXnE
8IS+lxi1L+LEmyZJom7RbjhSXsH4/x6LYEnZAmAEvGKkFRaq/K36EbmkqD/FlKoP
fxaeqMZNyO36SWq+0ae4/qTbv4k2afEew1i7FcEVB8ZKxLMUI71P40sqFdqdzh1m
W7fupfOvW2lukBy67fvDemWIMxRFszlsVdVnxqODeN1STWk6/yXgaTMgH43OSM/P
s+r9hvl3Huj7HKJ10T0Lnp9TQPP3K1sBJDSeoxNojD2CGOF7Gl5sJ6D6TiR8xKYe
Y2Kr/zDcDiCj6v2V2IFZJZuNg7bZMSHZtErO7CGofxWYRhfyjBm67J81ySPHdJGR
eV2j6JKfDwCaTotREBZwDpWe1ePrOKXARuxUPcyHmJ22coZX+qgD+nX/bpgBznjy
aPAb7XOKCFK6Qw2ZM0SDkUyWRQiABFePWnbiOvk7AYPPBrZS8BMRffqkovOd0TV2
hyQsL8hN93tHgIDdeMB9hIw0CflFn5eaCx2LxOpQNdGOnRR7vEiEECcU8XD13HO8
XfobZTgEyxd1g1Jb77P0pPvt5YqBoZcmWyeWkUMeL8SLJ2qk5FdH1U/J0J0julBJ
lQhCKzoe8XuVcWMecwBcq8SVOgWkf2MvVyuJKKUlA5VGvStjHUeCp2xsKFbEeJwK
+Q3ybQj3AbTl0SB5u1Js70VsPeq3G1sj85cjD1q3PVZgFfWChNSwKLR/n2weFeKE
qF3z9GhkO/kvvvpExRXInIhpGGKel4wTKB+q483G5U0v8oM1kikDvMIB8wXfLy0Y
kFLCn2Up49rlOkLJiCwBS5jKwY3GbCrdx209VRsBbbpWVvO1Yhyf9ggCxQcqjciA
WyVD4xCORxoFnaGQXWsP6rkbk5779jhclTmwetQsVGKJbmJu11QOhYWWVVgO7OKv
FVaAwunnBog8a8rw13lZN9lfwbdWm1TomMinL8EQXb/Fo0ViG57zNwUHhJ3Wpf8z
zYAO6yuPqCNVtVkoDb95PBXoyJ3Q5hRKFSAdtwSoehJgWAkvaxSE4RCFdsBN5wwP
icCDV1T28ITt1W18V0ygIbTA/Lfwk+8nmCELPF6SzdPQFnd3kljQp5oZKS2fTRPa
g8DGwzlMkMVw7ghh43nDCTWy+202E3vFSvMP9kfNhZ/xJBH8TAzoI3v+FDbumPBF
nbCFi63UuvH8ixTALdTIsApzl1SMDWKYYNB4jvbVLEKZedYnNNDTLrTZ1cm5e7lE
0csQBnGY8lq97zZq2198vmhlSlabKeju03ipd5DaI7q13Kr9/RWQFYHonHtN4OxP
C6HxotSky2kany5B80AGuqN4heJhViMgm1/Ll78Q2UHQdhilEIqy4LTGuxSrLsuw
WOiptrY6At68eOhQG1h7H6W0eQPLH4j5XdnPS51w0eU=
`pragma protect end_protected

`endif // GUARD_SVT_AXI_GP_UTILS_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
PfCBp6iSM5+iDBj/zk1EJyLNcOgAPKNcj5HFabYBdV4SsVyaf7AkzFwbZ7YkL/hQ
w8XcbZvDSS8c9HxxxoxyTvELTijopsUURjbzQeVF3QearlGGLbIYSxSEOCPOGGrL
8XAVVfJcIi2z4+jfbvNVoMzcgMwySai/SYvJxQXwhK0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 19949     )
aslv9udMWi3QS2ZNJ0TFFnsg9HwYOCAwbMIS1MeEi2YjQlSzHGd+3QuYcTfn0fSd
pudvq9mMF1s+j5zusS7JrUEjIRQ2Ggmy5vTIQzxyGe8x+HMlC67QI/qbCXFs19os
`pragma protect end_protected
