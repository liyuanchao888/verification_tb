
`ifndef GUARD_SVT_AHB_TLM_GP_SEQUENCE_COLLECTION_SV
`define GUARD_SVT_AHB_TLM_GP_SEQUENCE_COLLECTION_SV
/** 
 * This sequence generates UVM TLM Generic Payload Transactions.
 * A WRITE transaction is followed by a READ transaction to the same address. 
 * At the end of the READ transaction we check that the contents of the READ
 * transaction are same as the WRITE transaction 
 */
class svt_ahb_tlm_generic_payload_sequence extends svt_sequence#(uvm_tlm_generic_payload);
  /** Number of Transactions in a sequence. */
  rand int unsigned sequence_length = 10;

  /** Constrain the sequence length to a reasonable value */
  constraint reasonable_sequence_length {
    sequence_length == 10;
  }

  `uvm_declare_p_sequencer(svt_ahb_tlm_generic_payload_sequencer)

  `uvm_object_utils_begin(svt_ahb_tlm_generic_payload_sequence)
    `uvm_field_int(sequence_length, `SVT_XVM_ALL_ON)
  `uvm_object_utils_end

  extern function new(string name="svt_ahb_tlm_generic_payload_sequence");

  virtual task pre_body();
    raise_phase_objection();
  endtask

  virtual task body();
    bit status;
    uvm_tlm_generic_payload write_gp_item, read_gp_item;
    `svt_xvm_note("body", {"Executing ", (is_item() ? "item " : "sequence "), get_name(), " (", get_type_name(), ")"});
    /** Gets the user provided sequence_length. */
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(m_sequencer, get_type_name(), "sequence_length", sequence_length);
`else
    status = m_sequencer.get_config_int({get_type_name(), ".sequence_length"}, sequence_length);
`endif
    `svt_xvm_debug("body", $sformatf("sequence_length is 'd%0d as a result of %0s.", sequence_length, status ? "the config DB" : "randomization"));

    for (int i=0; i < sequence_length; i++) begin
       
       `svt_xvm_debug("body", $sformatf("generating tlm generic sequence 'd%0d",i));
       `ifndef SVT_UVM_1800_2_2017_OR_HIGHER
         `uvm_do_with(req,
          { 
            req.m_length             > 0;
            req.m_length             <= 1024;
            req.m_data.size()        == req.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == req.m_length;
            req.m_command            == UVM_TLM_WRITE_COMMAND;
          })
       `else 
         `uvm_do(req,,,
          { 
            req.m_length             > 0;
            req.m_length             <= 1024;
            req.m_data.size()        == req.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == req.m_length;
            req.m_command            == UVM_TLM_WRITE_COMMAND;
          })  
       `endif     
       write_gp_item = req;
       `svt_xvm_debug("body", $sformatf("waiting for response of tlm write generic sequence 'd%0d",i));
       get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm write generic sequence 'd%0d received:\n%s",i,rsp.sprint()));
       `ifndef SVT_UVM_1800_2_2017_OR_HIGHER
         `uvm_do_with(req,
          { 
            req.m_length             == write_gp_item.m_length;
            req.m_data.size()        == write_gp_item.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == 0;
            req.m_command            == UVM_TLM_READ_COMMAND;
            req.m_address            == write_gp_item.m_address;
          })
       `else 
         `uvm_do(req,,,
          { 
            req.m_length             == write_gp_item.m_length;
            req.m_data.size()        == write_gp_item.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == 0;
            req.m_command            == UVM_TLM_READ_COMMAND;
            req.m_address            == write_gp_item.m_address;
          })
       `endif
       read_gp_item = req;
       `svt_xvm_debug("body", $sformatf("waiting for response of tlm read generic sequence 'd%0d",i));
       get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm read generic sequence 'd%0d received:\n%s",i,rsp.sprint()));
       if (
            (write_gp_item.m_response_status == UVM_TLM_OK_RESPONSE) &&
            (read_gp_item.m_response_status == UVM_TLM_OK_RESPONSE) &&
            (write_gp_item.m_streaming_width == 0)
          ) begin
         foreach (write_gp_item.m_data[j]) begin
           if (write_gp_item.m_data[j] != read_gp_item.m_data[j]) begin
             `svt_xvm_error("body", $sformatf("m_data['d%0d] does not match between WRITE and READ transactions for sequence 'd%0d with address 'h%0x. write_gp_item.m_data = 'h%0x. read_gp_item.m_data = 'h%0x\n",
                            j,i,write_gp_item.m_address,write_gp_item.m_data[j],read_gp_item.m_data[j])); 
           end 
         end
       end
    end

  endtask: body

  virtual task post_body();
    drop_phase_objection();
  endtask

  virtual function bit is_applicable(svt_configuration cfg);
    return 0;
  endfunction : is_applicable
endclass: svt_ahb_tlm_generic_payload_sequence

/** @cond PRIVATE */
/** 
 * This sequence executes the UVM TLM Generic Payload Transaction in its ~m_gp~ property
 * and returns once the response has been received.
 * 
 * The GP instance is not randomized before being sent to the sequencer.
 */
class svt_ahb_directed_tlm_generic_payload_sequence extends svt_sequence#(uvm_tlm_generic_payload);

  /** The GP transaction (optionally annotated with a svt_amba_pv_extension) to execute */
  uvm_tlm_generic_payload m_gp;

  `uvm_declare_p_sequencer(svt_ahb_tlm_generic_payload_sequencer)

  `uvm_object_utils_begin(svt_ahb_directed_tlm_generic_payload_sequence)
    `uvm_field_object(m_gp, `SVT_XVM_ALL_ON)
  `uvm_object_utils_end

  extern function new(string name="svt_ahb_directed_tlm_generic_payload_sequence");

  virtual task pre_body();
    raise_phase_objection();
  endtask

  virtual task body();
    `uvm_send(m_gp);
    get_response(rsp);
  endtask: body

  virtual task post_body();
    drop_phase_objection();
  endtask

  virtual function bit is_applicable(svt_configuration cfg);
    return 0;
  endfunction : is_applicable
endclass: svt_ahb_directed_tlm_generic_payload_sequence

/** 
 * This layering sequence converts TLM GP transactions into AHB transaction(s) and sends
 * them out on the driver. The sequence gets TLM GP transactions from the
 * tlm_gp_seq_item_port on the parent sequencer.
 */
class svt_ahb_tlm_gp_to_ahb_sequence extends svt_ahb_master_transaction_base_sequence;

  local svt_ahb_master_configuration m_cfg;
  
  `uvm_object_utils_begin(svt_ahb_tlm_gp_to_ahb_sequence)
  `uvm_object_utils_end

  extern function new(string name="svt_ahb_tlm_gp_to_ahb_sequence");

  extern virtual task pre_body();
  extern virtual task body();
  extern virtual task post_body();

  extern virtual function bit is_applicable(svt_configuration cfg);

  /**
   * Translate a TLM GP into an equivalent set of AHBtransactions
   * Return FALSE if the GP cannot be mapped
   */
  extern function bit map_tlm_gp_to_ahb_transactions(uvm_tlm_generic_payload gp,
                                                     ref svt_ahb_master_transaction ahb_tr[$]);

  /**
   * Annotate the results of the AHB transactions back to the GP
   */
  extern function void annotate_ahb_transaction_responses_to_tlm_gp(ref svt_ahb_master_transaction ahb_tr[$],
                                                                    input uvm_tlm_generic_payload gp);

endclass: svt_ahb_tlm_gp_to_ahb_sequence
/** @endcond */

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
F+nhO0ArtiM/MHOr9F+RnVL+5jAeypdUfzoAx4WA//kjJk6SQMqGcvh9p03ddW93
s04kPbtBBISvMDC/cEktWUG3PlyyQ5fdseJrpM5GIsROCrA0ieA3Yp0px1CtuV2d
0YPw7f5mgM6RBQymaQ/216cUcCw2rE0TJ5LfHNX0oaA=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 22641     )
Na8RB/snjSvacaph99FXpLM7yFkLjDmlRc+F9a6I09ewxEZnKtTBygdYQt7mbONj
bQZtS3r1vETnSuICRlrU8Q3/wC1FiSq6JHBegrFcPJwdo2NUrU/qF1B2cE4dLIoe
oeOJRGErDcwenjQJ0w7pVrSjQ4SuKPnZCUhjcwG4b1QMk2u48DP0+wYFDzwkxcfc
y3yNgqy/M9loAPWaH+LopOGKRpvPXKpfdyfuwRrwvjdy+22HF8XVofHECk4lr7Ga
CzDpDePhyaz5W1fX7/gcPX+KM+RgISzkLOA9TBf2RvmS7ZbdN5DJ5tPSubFdCxtZ
HZpbdSDNri2p6IaFDTAVG9/Vgvzeyg+EpUHmCoKZ6mKNGH3xSDvuBRpbmC8Ffls6
gk+MVZRS3lWaeuy9jk/E57U+wDJ3EeIMDheAQ5C/PP+aZP6t07Y95v9Zo9HzVSwj
tKlpJloGzcKvs6BH8r7mb6POUZ/2t06IK01vclK0f4Nh7O1S0P31Er7QP21GwwV4
2omaQVXnDmATdjcOFEKaBrkZvucdF/uCGqWxHtIVlhdJigdAgT5/EyznhsGWLGEO
u6lDOaUY9LcyvJrqqgGy5Ssb+5btyDrhwikri8b2FKF+pb84FiHu/wksdlQgOK9e
rubWfM50DEWCcmAX5gfI72mJtkTQI7by/+qq1ojy3pjXjC5DACFWVY4u131iVLAi
hTh7aL7mcqGOPf3GnuxVXF4VlsmUmwwLac2ZohrGtPvwlE77bjHIuGOt9bPtdJA9
jfzMQFBxD3Q0nUby7PnmGVkF3X4oSNGx+qoG4Ykcnaf5XYoRQ/0TeAXmDgLsTZkF
MtNkN32nXpREepzcEXYuJJ5U+Rgwgr46MlP1uQIgrh+MZtM5Wd9WohuwJYrbJPfO
2IZcXl5YzX3J4Ix5HM2MfzMZDWahlrkxSSl2gEX2IRXDSjyeNfRa4FHTUImCGMsG
JVXilWJePop8xwg5Y4b7fH/g4V5713mD7D9cjH4Q0zwrckPFR+tX/LF17KQLAUhm
p5H4XlhrQEXAgeGKbVVzDPn/BqHycGAlCM6e0N6+YAH23A3jUv7H+AB+061fu0Nh
w2ihlnv7YemL8uQrXAcTz8TdhWSJq0+lgMU0hFP+9bIhv+0oNmhnNfhSHXDx1Cq0
ZXWFZO3XFmFHYn8EPx5HbqQJTIyUatmiuoYLZy1RgZs7Hmrc9PiVrXqugwHnFD7+
zAgzz/T/mJMiVoktP4LRGGq2NoHqJTX85fudH9xjYlOs3/NKak7MMsNZY+3K7dT1
odcmVM9O1gKzUxpcrdtMk9At9PXu6kuYqaMHYwXi9h7joSYsRWwSEtss9CqfA5iR
5vQyJ+9/123FdiZRItZOxceWWSROasrBwPxMHWXz17amxR7YJyCFdLaTLf813VAS
XltTu6ZLkInw0XpW6wzMbVZu1NRs455Rqzk5WBoTSccUvCtOlE/1vrTbSOkoi3Zb
CuYA61PfK/0BQeGUep3lYdZpZq41vqMPJKLP3E+KocgCIx3JWdeiUO/WAHb/IjxP
wAICXgnaM9w+7ejV1zYzJx2kPLgwncpZLtgRxDjGkPoV7+kF0hBTu9EQ31Nfr44B
/SdvNiKjsTaa8gFV2vqiopgDCkjB0BQBQO4tdpVcVXw+BHqUxUG0eoLaayAiMFt9
cKg5IWv4eMu7NGbSjtx0+G3uxl8J0Q/uaGONuaKMSGE/pY5Qq4bNGxKLQ9zIiM78
Y68jproWz8XA6szdKxNH5ahYQtya4Y8SaJUk7lJZNpfYhOVfPWcjZFo7m7nl3bv+
Kp2h+QEvzGwEHgnVxs5DD1sryEzK6b7fsf1+B91pN3L/sYLpKIn/Ysp4mBvbb/sx
eMII/W2B4cAi45YPZY9Z0I8xd+RdDQnNmCi/E7JdDkiNPGY5YHu/pytKwxYr7zLC
+zHW08jcJUP2aIAcf1XH9tb4yv2Prekg990v80lAfjb0GhmKboBYT9tNGGaRVuy5
AZUeUuMngenVajrP1j7+ApP1gGFrkaWRchX7PVZIiWim98CAK9lkNjRL53Zo5oAm
EocxwCUi8WRQb43H31ARVjEvFdM2RSBEMD1ooDzRPuJ6d0igCupL6zOGjDWv6Bf8
6LFuWGuweueNdQjz7F6m7ovbwSH6/6JADu5OB/bkfiynYlwQcOFIxMlk3O6mIkiP
rQa3vWlY58CQI9M7Fr2ecVeMOX1iC7plppckmqVy/y2qu2MCCIAXGIaB17xiYvAR
/8NHBY+x+clFnqBBlRRtVZLCmyf571GTz8yBpTmPTgPb7nSfx66CZNZknnSiCTTF
vWAku68QUmqsWy6ZbUhtRlVg62n2EfwVbP95gwuhkFausC/4U7e5aG4k/LoVb2/1
j/gEaGu5o65KgBI9dsBcsYXXOs6cIPaQTBpDXaBKDepadnTbOmJ9MBkoh77nwjeg
hmHzZvhQp6bAGUDPgowbojjJwI/E992uNbEaLVkC5J7Kg5HXHn5cL4ia52nXZy/t
nLIfDj3vr0UEYmuBINpw1rbzmIlrSI1EXwLQ8RB4xLT5VGAtw4M8bxqhkrsXby6b
hm1h3jnx+sVb+f/R3mPMoZ/E02Y2ubaQ6vImrlD0Yv0BpLD1LWxwQM9PE6l89rIw
ShOAnzkmTvQ1VN5DYYO5SxoWl7sVFnTfACttc6Es9f2Rll5y7XzgY2ihbjpI6WCN
Or9Q3mDfhg+m0wIXHE3SyCXsaVRXKWcC4kuOxrxtbPO6odJts+oQfac6ehfNUxyN
RzO6+zK0eEi2cXfaifF/S2jcmAJr8lyG0J7zYPLAp0J4F9ESQ+TSRfyrQIfNqX+l
J+ATAzmyQmUNe661bCqbya4KsPjjd8eFHoUbaTo3dBgeNq0H8gDF3UtQDQKhLrEI
mZGg9dcbuXyKIMvgyNgwNYSHLztZF8IERwUd1yG5821nYrQJRj5Tpn1muFUM8CJv
oV+Y+yMMiH954A1pTYGeX4y5SbEqwDPoDmFjM0E57sdcuqtbaEd6vH/Y477FV/6z
z5BJGsJ/qQid153Lk5Iz6fjoK8unAmoWossA6Y1JzPpBRVxI7m8+UrVgnlIONR8N
4VDFvWgu3E2bX2Q3x8FXBVYouvFpUsdsjrWAR4liBunESpyrxRYgtdUtpxdxHy4P
iyg7PW/LGZTZrFzrVy8cqM1l6ynlYZOWMIK3uR4wC9cnY+n0qxjmn2QzvA6oSCjY
KE38HEBLTxXbJQWVoZSQogGntky0G8MJvZdJghB98N/uZHHOzohzjJSp1LKsBy6x
jLw9fUdaXDPpeRC15WrTsPXTisronwRQPg5h7xqWXauWT1OLm1fgMd2ouslDGVEP
JKhGSirzWRypVT1+AYaHmnXksShcjnWmQuFFXoFuwt9RN39kakkUyP9eQx+zT+TL
ElfxZmrWue6zH8UA5Hf5t9yCmx5PIK/rWcQ94nH3aK0j0C7n/TiPiOIUsGw543V0
InM+W/OX+rvfnuKox++4Vyam7TfITGJV2PooYAPbuBhTYoMHiorIFFaymiyk43Us
WrZMqytcdNdUEov3Db3bLShZnO86sk1GAldM8vCJpr2wNY04hQoYnF7uwYQyE0qt
l0/xMgpN4x4b1Tw2o+9yyEf1Ow6wxs4wFj3tVXBoCMf1cJVpTj2vzwMoEe/fLQsP
h6Rk0i7drLEQWORmPsK12miAuGt9brGiBoJWFodxJnw/bPKLhRSNa4p/0FYJfvrz
TAO8RTPOv6HmCqQl78VDZgAA7Tbc6s8Up71Jh7bg6/lB9ZDtF6DS+00I3jmOdSEg
d42sk1wjcNbdFhSHpaOxUvIDd2BARjReqh90tOpJcnudR0DuzABqUdwrdKrFa5vs
28bG90jKooKfHraQ1IpQvVbd+quAPdBIgaeVygA1lsFVWplGq1iV07y+nT8RNeHm
IK+lldlYq/ToCIkDURhbGPMw6tYQrYnJ8+XcauzUrnQyEYu0rQM+JMZ8Wv3UVRcG
ks2SnAEzQ7M4KvFxGeaxC2esY59S+M/s6i5PXl3GBUCgX6gyTx1CnOkdIvWoOp2s
D8j6EZLdacnszXnYu36YBV0lb0MLmmwuM8RfxzQb8HPbvtau6I5ZX9aQnTBnumG6
knSpYPNgFZM0asXHcehqX41B8fX7ZTQT3s0LcCMQPHZo1EtmC3pbhW4FlKcru0K9
MJMHSXGx7kug7Y90up3N1hT68ebnd/GNURqFrhDURAuSuKcMtaG4+lmnEt/FbR4S
kE1moA0qK4tTrNuv+/lD7V8GupslimKs20aLRnpWI/0E2YDo02DYrI8fVV/NchG1
fZOmS7B8xB+GOn0B66e0itGMJXvPhUk3NqJ/9IbrUDijG+UlSttWLjg1xlJdf81v
s6r1dW6U+DI8aQyadlyg0qknIo+RCViL2uND18UkXBovqaSyu2nlj688wcwdvJv0
rb759VRvk8Dg839a4KRHgfZRBrpsCWQJztFaEoRxIG28XTAQCklqznr7HtysYFna
FJKggoAyRqiU1qekxYT10o/6aYRkGjFGzcFauNyEerAs2dFYpYd0lzgqd3jSfAv3
MqyuBlbkPznXoUN4auYXKitHv1lz7CDxU646nQxYDxyI3VJib4QcRfVfBolXFudn
iKS4D48ZLQOOAOFeBvXZ9SpBZ62b69riv21xSRL7GNwDT22/F1IJJBDpzgDJKqP0
hI1nw0iR9wcP+MTyFUSveRX5jVyP0WUwCFfdNaX8nSoSDqNE+OytZ/H4zCLZ4eJF
pw+/XradT+GkqQqk7YJIDQDshH+sov0TjBoo09bZj8vkDW8p5dPgzb7y6pWfLyhw
JMQ+ANE0efIsqZ+eIqCg5rDedZgfD/QyiiVgeOxqlqHvIxw5o2H36loahnsaRCTi
/MINjf4USTuNNCz1C7OYo3exYfb9+ZadUYbssd4iVreBNdiGni0RUeZ/3+lNSEV5
cFkIx/ioKr9V1JF4HrMKTCI5Vc2Q9vazjNnLG+8+3phpSR7t+4QmK4pufh/49x+o
6QwTDwqOjRqpo1bTLoH+6EF7UkKU1QH6F/+fH9+nb7hbYiVU0hT5ZyvpQEU8AlGB
z7zXu2VZ2lOID+fQtZK6MYSncNfd3tBEJnRQTbTjvOW16nI2y7GJP83YrfJMA6LD
puKW4jrAt91T/TDPxxHoHmF1PCakt88csCRuoydE2XCwGiI4P8duuTt0QtWyaERw
s39X5KoOyX3aQq91onXjLajqZvp9ghVGLHa8O195lowdYsosLsRapRVvJ7aA1Jkq
nlm1cnpURJd6MGw9K2hs/scRIahYgYLZTzCwaXdCXTwbiRg+njbWZhiK99OHgvFo
wcBpR3PQzP+dbwN9Y2mjcObbmBbhxpKt1NsxbpckfzKGVyq4ydQCsrag5zsZcX+m
rkWspu6IaI+2SxyE+7nG/51FfqtcoLmWIYKaDBJWOcWM+N2iDRFAnTH3i6TSl92B
lkbt7XCx6NN+aTE7Hybl5teb1zeYWjywmUiZS63BE9gssHHZbOweomB667XJjjt1
d+bheR4ewEAZJQyBOlwYtAupJYb7rejCOXHFp6xFs9JII+NCrwiZhx5udLx2TK99
ddKjPyl00kPqx/LNVIve49B7HCqIaL6aASHLcrzhmztkPzOdloH/JmBmKmwUZlb1
tRG4kPWyilX2bUBZr1oNmOcR7pikpgv4CWBlo83yrt1GVmMtKkEvmQvyXu11BwSp
pl+CSTceAd9Zc5rMQ9k5AcE2ahmo7uBM4wnbz8sXCZMglkszEtDArphJlj/3rbBl
QYAXCnv97KJzJ5a4aWwTreDNbFJ/REEwJaTmMvaJWFWcUNIrRp0P8xqVVcjf7e+J
UCw11o0U9CiTLyq4NDtqDzPUwumSeZCsBtN6ecqlIbL+osWqxXEpTGBDcBWbhqe8
u1fkLD5zxnRHL/SeeLUaszSdPbiyNFwZTLAzVTjpevy3glluysuzKAedjFi6ZSk0
fspiiRfokqHXMxNI7kRotpgYP0ejuhNvkOpVm+XtlfXcABPRxTgsOQMxNfVYJoIu
vF2Gvx2B6hIqYR02AfGnvLjtywvWPXSJEm6GulWzZ0YOqaKzcpD5AE5sghfIIg/O
fB9w/9WnUHy3IGBolWxBnE4NyYa5bHe2vCgKuTq9RROEnlgS3U25ke+1s8wXeo6l
UE+zBtmzgYqr0m4v/AX1oTXhUnuEo6a4lGYWnKtnOtDAAnrh3OapgCyI14UUU6bD
CjPypTtvjgFk4bBPlsH07w3r2UQav+BKgBDBZwpGwOkiG0GoAOtF3nISJHyMhzgK
4RF3ekDgf1GcHY7EBQI6BVwpC1ucc7cHycxO1hKzKLLCed14SkBXaANHCoPT0FV6
STT72OlE35MDlPw2MENP5fc8iFTlNO/dsHGizLO22Kt01qvWAQIZeA5sQQF6yyU0
PEwohxIyxZVg4YmejGZEwL5Q/q7+z+5mU6h/KjKkOlfPFwgkz/qjg6YRIEBiMSL2
j0kwkezWKHwq4v39Jda4tb+a/8v/nZStI3la8szBFLY/vTMDtE26wkrxZhiZwIjq
nb+RsV0Timc54HVlAfGW7dqUUs3Eknd/tjVrFpgNh6RBrZ3o7qevWcU3DyLJECvD
CXu/99YcDVse21p8qzgbT+3wZW1iielAa5SuNaZ5PUUIwfD8posvwU8K7DtQMuCe
cFFKqYV3pUNzv+23qe84OawfB+JorlR6COomNQ/4QIEtRw9SdgG0T9DeWHGhfteN
UJA1qnHKg/Ltt15RAf3sYe9gIWD6JsXQBUgm9AbcVBINyDt8D+6+EZ3sbSQSbhg4
mffTM+EktFlnXBE99j+saTTzbkIJiUIgsK3aWC+YQ1CRMwZY9mT7vxny4AXv6mXI
kpTe/4ezqLNrymcVa7VW1lIFa979PVpIfKXeueEQF0tmU0BAd2ZHgZve/KJ+UWRw
imdgDRlBTU89xZKE5eu6d111onm8KENi00YPbQ9/SWD6Xpk1s7fyk4hlC8QOPDfI
ZNcQ4G7LSZQfFcnv7jolaF3dd1cQRunYJr/+KYYqEYJl2fRrXutwTwh15Pj7MQeZ
HiYqu0kuz83p8eKM+4ehiT44zTUDf6WI/CTwV0v1DZl/u/vwv+M0lpdSRZzHVe7x
DbZouFFrl5NZRgyIVfL4VV+izIuw2ZNvTFTnEe9KnRwXmRCCu5s0KekYi1rX3h2d
Ds/9GhbTxEmXyFpxAc+ZiOxl6qZ+PrJHC72w0Cg7FmYTiOz3I7XppxkY2ojOg+6r
Rrk3o3Bx7AMpvB99H8ZRe4OOh4s9f09/N+wCjoQ9+ldImnOGR7NyV0rN+BfiHk1s
HZTxWlIBnEeGfRXVXwfS49gYDwgKfskxK4MlrTb84s9Nw8ZRqLeD+X+D3PY7ZZ7t
p1l/jOr6ym3lE3kQ2eQdE8bq5+84NjToRuJWe1D9wmyy1vFHL6tm7pT1BDAnlhur
HYjXv0ZsEEUcualDmGT/M7CFoWjfHZJkyEiXDYYmnfOUzk6iDvEMxQHe4GCYlrIO
bWaxlO7WFowX7u3EDfkgxHHgDP457sFs8+Ic0vnTOjgsJ9EkPJdq/uZN4HN/afOc
hTR1e93Xn9xmSXD35HEiMR1c6i2er6H2kAUe+TAFsMvXOC86U7N5hpDYpOW+hOR7
yjukwsSUmyrcORSD6vrrAIHFDpdLbr32fa7lmVvD7b/W6KBXnYDZYOY41pNkksp5
yPepx5J6PMK1LpBnpedrBR4p4ZUNBP4Pz9BLaE1jNWXHPQNoLcEuK8QypzO+Q7RZ
ISVVwZhCobduIj+V4O+TbhEe54Xq5dnB1i5Agc2TeahPfeDjvuzX/TAOw6IntMZd
2S9Tr6cC1IACI/x8eAptkSTS4gPt2CXTTrUvZLA/V/WGBWAStfIIMwBjGN+8r0/c
7eX9qtjMQbP+iSIlFKmR+X6gtFrBEDRj5jvfAOr1Nw61wsBPU0PjRjRtiMaDmx8u
xBgGCP1WhGTgY+WnlZ/RtzkvkeWP+K1wtd2PM4qe6hj1r079bXhn2QG1e8zhOd9l
6ELmNun8M4sxxBJVFeLQ6+A2fp1NT2dvfy9zoDViMeD9xNISEdAISm5B3sRwtcNu
9NswwMyAeQzwWOTfjNriP13Dfd9XGxUll70bSLNt1WjHHl7AAh7xppEM0wiAsJb+
WIQzCbBoCkqvUT0EKOQcs1nlHleLnwHxvfeq/ua5BYZDFjVqIFoARZMghARFH35V
Ct3SOY17NwUbruLK3H4GVC/Vk7a/g/QM1BsaND1cB+o5Z5qOLwOxh6mteMz41yGg
cuEcIQXLF03r5hroGbtneZo9SfS6uUmkT0PbGJzNRxP2hBGUqXUzf4FGcuQd6QHG
g9VT0meBiZIJwT69kbIcEGMM54zO+uPD/X66QHdBavn3uqnklUihbxUBsaKNjitD
dYGH/tpruWdwc9FGyf7BDkqwvMyYiDjvUTR3uViGAfBh/4XtInb/l78D2FMCY9zt
sHU9mAscS1bnBB2Q/+dtlc4uPZDZSwZzuf4BIIIBCDAFxQEhA9e4Sv555+JjdiHA
VzyjG9PGd4wJBet1tV3UCBaGzEGRhJNulY+m4rONncJ0nn3uSB80tBZWY/bbo3d0
QZQBynso1VU0RVt7C8Xo0LlVsDWLKCM7VUl3QLr9sWekdxdLAn3bl9v4CJ5eBBkB
Y5Tc6Qpl8FTMryiObZraDSh1uwZR3IxnMdCGW40P8d4pB0kpDfqI/tLgraQK0hgX
drYMj3gRQvRQjOE44/HWoo+GvPdzcMDg0NC8PhR9lwp05mhs6SRJMj6Kk8lZD/my
tWFU0SL34SdwIdlsBMgRRjtUxgetqZ0sVESaK2Ltbe1t/dI4bLVeCclq0wb93QN9
TggmyTZjiPL/JvjlRvgZJGerD+q0lpq3mmcuquShczHw9laMbB3i14BnR3bvLnK3
R/2yppxmu/HK6SOFxLIc/ADy/NZ9PjBDaPRMc6y6BGvfsbBM3WmdlGI90YWToiXT
iAPcX9VZnCfc31ocqGkf/jJREr/LkXr7CAltZ2w1eniopHzpRsg92a2udza+VJ/j
nyBzcJ1EOT3rl84BfunnvF+bw/N4RMKmO35BUsunP16Vgt1eEuZpE+YXoDjafRL5
9wmSXLz2IGAfLKoI8Vrd92Y3j3cx9wjy8wJ6SN7aqhVhXqH+zQt3TGQ8CL32wNii
CQ9elwq2bTVyO7nqHF31yemxL56Ugwo+jtvUycrlru8/3dwlGBMJIJ/8JpgrEFu3
xyaqsEIMBt4I+mFoiq5c+QVBYWQv9PHlCafZjXpYyeWBv4nq7SEITaPBz/gM0FEg
b1UWAwXwj/4f1j58GPY1yFCjWBQFlv5g2rmqX7ZnX3b6Mzbcbdun1HIb54ufz+NO
UuITrWHdYodptKYNUqAMOOO7q53F4S+/oqKbVrf4mXXDBH1PSibTrgOhFFSBzfM7
B87Dk9gEpseUUgcnhXIsjnt6nbjAq8/qRMN+bxJ+zDMe+WUgLCih8ITy5UWZs7EA
WHZkTQTyA8R1JSZEH3hLrCgT4raCdrga+7lXAygcGokv6omPa2pYX88kYpzZhxa3
M26/Moh+eSzGbKaSOLmB7HpyHN+PqN6bDKOja8/fertrxK4YrP0y8c37D3Fm9Aq3
07ZaqjtkyeuDg5hxarfaCzoVJEisW0ZdvGEWfsD7i2m/vk6j3bHv5J5rYwxbLXfZ
Rm3F+YdEEPbDHoCcJLIUV0Btrz5aRcRiRnGfKe8aXCB+LZOiyd3vR0hvSpcmckrp
ihiPB26SQznBMJadN+i5mtG+O4LgrUC51UoseIalZ0kdetiahQx8JVJOj9i/GDp3
QAM4x25D/7ebfisW6fksMj5vnAwwID0jdyHb4DT+D0iE078kPSsbr46V7a+M6dFK
6244wbmBp0j7qSP2lxY/0wH1BWKT8k/2XdXLehrCHFpyA4yWYA9YWRS8closoFhx
aEhsrvXC/7wIKrzbZ5tDGaBVLbQKDHUrRuRqXcJ2qpmAtHolukM2s+MYs8j81lYD
hExa/nQxzmLmN8udiSK4HeDCuDCEi+j571TAojgXZn3jpExfnKOVCrUDg09Vdv9Y
YH+uZlmcE9K5R7/efjHVmEjkbsAdDblbzqRIzPwfTEKM7ncFf67EKzas3Yu9JCJJ
WWrQTzEqrpqdPKtVgDXDhkyi1tXuWtPoAFGTeLEiHWuDrtRysnQYepKA5+N6cI68
uz/lty9PMSZtzAuudJ15xtgrN3JL9rMsu2uZf6wg+sK7L5Tr511SJffcFTQodE2k
uVgGFV01XjqIkny2VRUxO2pCc5rvqMQLlu6XZGNBsGBY58z7kNMCXjLGUciSJRxm
4SX5xgEaVp7G6Rq5hXkKiqnQaeXy6tlF+a65pSLkeOM1gTLDsWz7Ax0U/qDnhb0Z
yxtw0XO7TvkK3GhwPE/BzujnYhz5Oq3viU6HZ0F1gXRjwua7fosCzwaJTr7pf04O
789FB2nrBUWMXeq5JbkWGuoS/KyjXHF7CssffvrNfAoz5H0sTHTaPo85py4YrSuV
VZnjEMTruOE2ZYnGwWFiYScFY1bMMLJEQ+PbrfLLbBeV0gfeSDRQBD+T8CkRevEG
g7tc9hP1mVKwCEvfMFO8GzAxLMTTc2eXjs/R/7egKEe7IbkMSYkPdTMHIVb0U0hj
6YLX+Qj/fymX/ryz59BHehNVnXsSAIc9K31SugNqoC8UQmCtpoL+jUVk52gNf0iq
+MU7lfla2q6fDY7Jn4A7svlyghS5UD2eGgV6j4Z1DZPrOtggFV8biDn5JV3iD1gh
FvSkwvGnA1xCQIkEsjZH4yt536urTdMIJj5PMcmuMD11w+Nch46jwI+hnoo42Dtl
NszQ6GRFJtc0cHTonEfSrD1EgnlZGyvxZBvd04On3pzi3U4ibQpk1wAGfH9yv62h
yQmeZgGa3ekEaai8nEDMQFdlfKiTQcbRLi2UD50GEN5UTU4ElyakY+D3yo/hnKUC
QInf2AMKx6rYYIZVULmtR7kZVccRaunqeD8GFRjfTNXxq2pgb1Q48HCJ+ARBq98b
cUYhp+NcalqnfOlUDJuW1koreSXrHgM80TFrDg5Qvpwg57XiBtKc97QveQyR43pf
HWN4qN2zfrCuA/ZkvfVY8syLbIWT8k8fdvztKNjIsYOelUqfKjYlBzM0tkj9FVkS
xhGf6H9betnfi83HzxJdmP0ZIWkSkozdBqf50nz6ApzdnAcfjnO2u7WuEipQZ1rt
qyqlKyNVNZnC6Ncf303ARtqyhfR013CfuGuXmFnDomUMbt5EQrXWG4xlHIzn8nk9
MuSf4W78wFG6yc/bAS0dk6/Vu3GbrsMjBExS/aZDyHVuZgG4RNrLhqB8enlf1iLR
BK5kvp72ovDNtvaYY+eZsxFyKGo6f+nfIrRSdpUStM4q5GTop896LVUlHYg3+sMs
ypYX8nfdpa08Ymf38RhsiwrvMT6wsD2U835/QAtbofoO9D6mOqyAf0SROMH1CVkk
+xKabpK3ojXvFxEcGvB5zTtk2VAECqLfyW8K7BLlw0EXsawWdhiYdj75wnN5VnmT
OgYcGTsCYyIkkjnuM4wqY6Oro7n8XeFb2HTVVdD7e5ZKTTH/6kxg2GbW00AxMYbA
tr5uYLnmY4fqGNn4Jn7voDR0dhaO+vsM7C/gNsCYEYCqY0j3e2nkcwndRIsEmmNE
OujcRc+0iisCZAYvOfy2bvpqlHZQyjKLP5PawMKjnyCx8OPgQNu8HjFFJYmVlQnw
vIhl1HVTFvG+N92rmPQoTzuQONJyIcruCrbdLV1djU28bWp77+VzQ1lR7qnDrJU9
0rhDXUU7X36T3g16qvWDEOJ+efcXsc2pDeBpFEiOMlL5h7dkyAsStSf4fVQbhEfa
sAJh+3DltKd4nkfd90/inu3p6wl/1iU9imA0lQOm5j9SKqxlWSrhktSJ1ctnYI2y
k48tawS0Kv1eZxlz4UPUOl7loQc20zfIsyyb7l1cG0/wEK1GdRW85HpjiwWd8IEG
ZXbSSUbM4c+wp2W5Ycj6Wu6//H9MzFHHdaGyq97dGiGRBYx0JexuoUwAnwG18qf4
dCLDjrKTwuxlz7sKDGkKWeCZ+lWlEtmwfNQBvYXBt4pgA8YWlAYS+2D3YdPMRWnx
QM2Ey82E/+oPk//PZ937ceQ5X1MZG3B7gBLzol4a8m1ebtCOk8euEteQyJDNxgZS
3KZnf8MJx8kyKfm9VTiLcpD2kr6UyXugq4GfaNO9mWPCm+LI3mxvVhbJbKOHYhGB
Ws7JbAdYnJ9i1yH5CMf3tWev1hi6t6ToHHk1TsbS7pNj1xUSPTo4sUqkGweQgTfy
gKomzs9gQdhRxsxGZ0KgyKiYNqBNgEnq2KzgepuroSqIlxn+z/miaSWrPfMJp3e6
TpEL3zZMiIxGGqfZrE6gnCYZQDK8cf5F6lj1TDeJqy/H1rcch0OjFZUhEsjmHgPf
4cPh+I3v5QRGoshwa+Skjat9Ri8f0SVJrSgFvFE2rDnyroyQYWyqfg4jp6xgdp2M
3t9w1LkEx/mCGhxHrsoF2iiizxkp+gR6GPuA5gV3BNOTsclOIv54i5TTNu0bIq6Q
lk/P7xm7/oB7XnzW1aY54pze1fSRZMC+oIIH67jaCB7q7CWjSh54m/DPOjck33qf
Iy9eG0DXZvCvHyTb2rABdelu72yqCmAm6idPW3c15tJ4fDwKrVJvK/FWLopNa1Ly
Rh+xrXX0P6tVe8ntIpo/bsmvnzoqtAX6VfeGiTNMIJhITHcWBvqu+jDs1FoqeJhe
VivfCfZy9rQ5/fXcV4fWgdbCqXOSKoOxJUXY/vAexV8nwr2M3oeHHD8nRdQqPoD7
zTvxbJOzQykQve5K9Cj1HDKmBbF4JsrtEzgHRKwG1PoO6R2dUOD8keu2Xj8TOISV
KplsApi9yoV5vjShnAhoQs3Mm/Amw683AcyO0NXPPurYSEY16ThMkcQqlnvpCUWV
R/e/N0GFXnDxGnoPOUYc9NbeTtPpNfy/Nch/QrHQ40tLp3pcvAgNjwoDCl9su5x4
JejaA/63P6F9pDLFm5DngTKqRTkJk0XJo7EZtbxEnR1eR2Ej6dCX9zXCyrP54RwR
UILmwV7txifiFX6aIi35GjzhGL+AJ9+6K/IZqAF6H9UEOxehiVqMEliNiKgfeBsf
Z63p8jJAEnowvSRpt6fqQerOocbwdlrY+M7GdDBrlNpaGIihwpKKdRg3FCWRCo31
Bge0LMx0W9lEUBLtWDY6TZwvXRve392c7k4IbEdOXTykBVSs+6uuhEQJb/MaSHt8
g7COgT1Sv6EjNH3h697uG7kiJftVZ9rAt5pD6VcpszGypHizBHCWsAJi6z/DSlNw
lcuHeduuElvNd4fIFXE+Sbv1BZUsC8Z38VO7SDexqvfiQCMGh0LbjIuQ9AwBOhNb
s1jAGHiTe6wPJzY9hDhuVReLjayymHfMmy7gMJ4SqOjhhIX7AFIE8qF2cRNT0C1q
qJ8dbC8TnrSrP8J96GBUyVvyPlWxZFYamkaG0WV8VHfZRg8qwYAZK+oC3eEbyMoe
H/OS6DPBR6GPt9s6d39rkB+jxgtu6E2twc2zu5+uBtusoYt3kaepSG2Vbyu7cLEC
foozA3FSekmouBV6LAV5vXPUXOfMHAarbLOaAqtcgQNOTPdskFMXXVZg/HLEHLg+
X6E2vbxAdIT/vRHZYXgJ35ImTBF+9o0wyBIB5pgDrDKMAECFIq2aFlX8xKQrkSuN
n/LvTN913qSigqvI4d35ldPrpkVv7lIU6p022yTJJPk1xFPS74IgNxUQesDjyeZo
YM3sXDZK3actnbX1qjZLu0KSjedKEyAN19Wx/+IzgcaYy1A0zzetzFKN8zVzFWpi
K1AJHx3UoGs71PxRkbHlngolmdikxxmlv53b5mOzTI3sSDfRQ3UcavIDW4I6cndZ
XDBM05ZJovwF1AOUJV8dAVy3JvhIUpeDU23bQra5zRNGcoHwFoeCRv3GqoS9DSa+
M7eN4ltJ6JrwXkkfDh2yh9K5W5phXa/kvviooF7QtXkzCd6ImE1miWzfnjd643RV
1jKkxcnKRfT1Kmf+xWRQGv3rlHzyY+hvxbED9PUjidop6FbDxM71V/W81vJka1dr
Td2AW/3BFq+73x/UWEAhtHlRrfU/jgxDMGdpzIpbHs09YxW1QMSOdFOB9gkjIkQv
p4BBiD8q7EDb6Ws08wqtsTp28wMJ34/m42Hvyt2Lcfv8jCqPejwYVI5iV6y3nJu8
y7CAB8I1UNj8SXAC0IjO0Yng5zB+pnBvNt0y3+IQkiJdbBHFinlggnveHS7MOZSp
JU/S3QpSo4gYBLHOFMHfvvo0Rz2YlJF0GLwY++txhfoxZQ8RFTexeeL5FDsbYYJE
zjhDVj7SZDyUP38HbhmDt+zs/C6mqbK0dcBlvxc7W4QCXpN/gyFInd3RZXppY2pe
UpGosTwEDiqP05DfpIrnziaj3cXo+sdGGyBNS3hqw2F5pCGtYZbAWp8qyfsXrQkm
0B68EgLIA93Oqss1LG01rbJqMUGFramklv1uzTlIilEFr8HVsVk251LIyS46+aXv
ixOkwsJVvTcwoNkTlDzVPiam34qn+GdCnnqE97iSageEubSaau0KnEWAK7IiI1rI
kpa8TIRMN2YWIUEfsEaHZY5mQSs+ja3JjT6UidcUisgYTddfMyS3PPFMiCtCSbNk
4Ls7qpHSkaYr9spaPyfcaJ9ghvhDRVGEP4Vr1AK0bXpU2WQ7moJh6T7c6X3RHS08
77w7LVTD8PxeJernuxKyWpEyppG6oB7625noSDC9MMztV95yHUX4lpRIiGDGCQVO
v1w6bBilFspHGAkWMJqmgwwEWGBGZkFt9dh68LUX/XIA4oJuWccYfzkK0p2F0BsD
f6xi9eQz50PwNuUHOadi1ooTmsiv9dTm+uSqMw/Nih9bUbiswFFKEr0FdaTDbn+r
zt3Izmrke96WYuHxarVdc0a/Tw7Hy3KIYJdpn7Lv/vpmy3qLuW7ci81PzqzCRBEO
CetKdd7a0rIuuBImoOVw9YzJYLpliDr7Y9App5zVfwGBUZFDD81z45MnOOXkxZVP
DmrzxKK5bFvPakKmFAjggcjXl7aseRLJXDLa7ks0JZIqLgdrPfWJzdPBpwfXuxyH
EqxajOW6EDdezovHHfieFRFfM79aj6Tl9tiH9B0IlmH0CgeTLZieYoQNznHByEKI
FzlHkycnKlOVfDRt3qRXmdIHle4A22SiaE/mKMqR9H8H6XmcRi0HCxBnQ+vWeW85
QMTMYVV44uI9N8JVC2kwjztVAhWWIqe2qgSvSJzcqTo1irE8pGpIEsbHK7FVI69v
mF9Sso/eb/hL7jChZRjweojzBwZgm3LEOqds7xvG24XKTuDDOFhy/1fW20KEHg6G
WHvuY3z/8dzFqVWIAeTpMN2Aq1kXQyuYRedBTSUeB42zAfT2j2jrGqOKenIr50yb
xxsEHiH/tnAASd9h3OOjHmIjnouDXtsBu45vgkyZBMqF43mJtrgVxNvw7nZb03FR
FkSQw0hgqkY98UbIp7q2lJpFqkA8JTpdP/0d2/SIg7xMkwqYIhmq9wBzsI66jLDw
g9saacOivwt9Bi7n6laB3qBSOx9vziT0Y8RmGm4N/EWfW3tiYgWZA51Mz8AY4mHH
1mQh3i+z4ks+glumTk3CE64+VUTE+L8k1gKfgHDNkCdGkjX2WDPPVniQHNla6hzb
K+Yx7QMttqas9FgTh+0g+zvahtSNQ9KN4NzpQURz6M8YNVKO8vW7WrmtXwiZwC9D
q6JsY760PQEecXL1lbilGjmspJycgTZouL//mkCryRLL/L1mk5XIZgeNy+jhrk0u
O+xt2D6yiiDsy1rZ0pwlF4Gz4Rep2a6lyP20OLaVDF6p9Dfye77fASXv9QhHlsZB
9uRhnAusS5a6jH+9XFSA0PJLZOhb4wG7Bsco75elu6xU2BpbZPLTxOQ8gAYfpbQi
/UqpDEif/PSZuYkADEPbgx0rpy2WpNwCqMXBCvZQXrobFJN+y75Zy68gmjryTdws
OJ30h6Vv+cRbkKzUhC+fB1bBjdhUkR/xUNKf9hirRbotCUE15PZl/6Hk8BGjsU0r
sN2dJVsyPZYid7WVptbqUdUfEoZt06aJ5WZEef9s7SK96VXD2Vs/UqI2uhqsFv5i
fpm/ILxeBpBn+5ymqzX0oNYzQyz1rwDnhzemEfXVoK+mSrI6qrqKSJsa9wrPdbzw
OH5d172B2tkhvwoYTmJkmQS/6hliZH4r+qQ0pkOSKJA8OzMFnljJi0+7jo/UB/Yp
O5H+JSUbtBKz5LhZOTv/1NPvziF0WezvasGWUynyPO7bY/ZMQKzKEx6jtJdehjDM
lgeVfgjr7ea63wnjN3hbszsYpjItATdxmNvzvdsnRPNdXQy1GiQvQOTyLdH7e20x
d8o2TY5QYqQ7NR1XpDswlLczXml03SSkhZKGr0HDm1IWSYW5my1MRYmRRp4A8Fuq
e3mMaMSUzedj8np8PhEKpCJwVmkVPmJWgGydLM8f20Kr5jW8TvNjgu7PzBm8LeGD
nyf7ipIgY6zogN8zPte3HiV5Hmowc9lWeQpl6bLikb2mYoTtfYQyxt9xDLmKRa/m
PKLx2RXM/TSFIgNuMnqVlo4fbl+9OHGp3upq96lSZaZD3Ng21xWL+EfV7af7Q+23
TJOEGl66yrFo7gnB2j7h9sOu7xKtNKD2fNBBGzTiHz32BHaubc2hReRVvGljfuS+
8EB3LtGTyEAaUK2rquh4zwPeEr2fD92X1gplMoAHpu79nAcpVcHuYepUftiN2FUi
ydmGrr/TPd3LBHVszVLkWN6cfAiGuFMqQIsZOVrCGRKmtLSBbJPvgK37zjUmBgH1
WJxVS6qTaHasCTtzywbSx6fEtRBRm5gh+n9CBSvWZx72gidkkonZ2vbCixbpcA1I
+yFPoLVjiYy0s9OBurYj94THpkbQymm5sQ3ggu6JjY5xNwSkJFwGh+t/j0ro9/rP
jQgUeQF2aYgqqcB+hWlGvhh/EKPSprpxfD6T7mYAzQxiEScfijwTzLSHPtTi0n6M
KvwfY9qYwFF8SHAWtAlponWMh2bdsbMOHvf1yn0bmOt551e4ErXANYgxVUTlqxM4
087tiQ5h5bOMMCnRGx9QQ6mybD4KT6SGtz2Dcmy2UJ22+BOPw68zbfl6k7rSLdg9
NpW/CDxPYVf53+r6kv7BaLHfnwi5y2xS3iLyrzHD9aXi1YyNHVeF8QrSgsnKtipF
hjNGQ0qxWTVeJ0y+8uR/CIzm66Kds/Xpg4AHqZgyb69XlTOoDL2Qg3zvQFIqMz0Q
T6xCieuUEytwnSiwdP2Eeps7odNyhCtF8JoPlnQ0asPFo5b9qi9rJFAymGGDD9gy
DcTVUVrUoFUMBgiPmstpHbvx8SREtr6IaeVEGgeVU+tLo7ui8Nc4QOHM+9u3ugzO
64Ry9/i5O27AAtpHv2yTXazHY/cAtA2fHQP6lMNp6bCSKfk447VgDYM9Q8X1WTch
Jqs+3a560O6MbwhgDE6d3Q6jF01ga3l6i9Szu04UbuEnrbM7OMqz2ED50PkbQFb7
xHCiY6QQOsnQKTBp3E96MdGhsgka70+F4PZqk1f8SLo+TV33rFkDtnxbSdblANwM
3xp2gVEl2qzIYgCU8ErNvGZ982P2qmz2+RV5AOxBf8fherTFuzLC6xdw74FB3KS7
deEAJemnmLs1q1kzgko9QF6HkkL0JSvDMy+iXBIUFs4ZqxmayRepivid1MXnmjxM
pTr7YswnoIOzA6Fcj56b6SLusUlzdNuFyrXjsSRBYSuT4p2Qc9NEhRh4TX4/cMhS
0Mr/bOfMP9rU8dAavcPlRms5Jvsb0HaGq47OgwQsAz4GcdmwgVBjYZYGk2f2dy6U
c5DVbwdKfxmjYKc+q2TiEctZ4K60aVVSwTYyyZmZMAvpCV6zC9CJ1femV+AKbTAe
YO+IjI5NvXAgrFcAghlR2TmgiTyOETrVxBSBOINhj4SWokdBx2UIa8hGK5Tv6rvD
B/sf2li0GkDBAkv7hsxJOwf1n+bThgQSwZT5XXINOBwcFUY87iR+Irvq1oCWM4fv
ZG+jXCAwD0JzND5iEV/0y5PlaUPvXXWr1tunWSleBRPta8CkB2kqOr1wL5+XpCzo
/xuoh+9GByT+kZoP/FT8H0z79xYW3YJmFawJ6G47hpK2INrcjoLEG+CGmVMxjeyE
lVbzGPOxTlph+SCuge68TGVhJWwH4eDtvoveAqxLE+D/qmOEkqdr3tixXg6e+5Bu
qwlVRxloFG8CBw4ZO+ORCcGNL62kiaXSjzmBhKKyPJKNMgYHJjZ1Kr0RgG6qHcqs
5DyE6Fv9ingwici4DQtQ/g9FtrOS9396ztW4gKlm9QiAjGsi+kZi7IM4zJ8RNzd4
MXp+PlvWJ5tK2N9Uy17wOO7JBccrRsPWAruy3exOzOSMo/2PzNIQz7X2mVRFaa7u
mcsqPCnlSc26w0eFMOhc0p0/n96Ti/+DyRj4FR25PouWgYpzYbtGsqFjaQ6rUjo5
VJmceqyGneIG5G0d678KhOY+mfVmKV3RlDRkRrUOh7NU4u2AlYsnyYWGCH7rIfCz
r3f77ZXXmDpqzRk+8GIOowZc9IiVUwiqQL6eSolju6wT0cQEm7VZqjjgTwSFI1C0
sy7lNyDVBc60QUqEHT7kRRuvdslcV6BKxvt39v21tNFydkll1BT2YtKkafATthgC
T0oevitBbJVRBTGawcsNlB/PzCDvAeUN+B9jN1KvTG5seeo9MDKFAo70wQb6Ksdq
JoI7v7PzDNKiVDYcVW+Gw/4cWpExGlc45rNED970dikMa7VWFSKAmMBw02mn1vJ3
qOVtLZgNVPaqloqRjSucWB3jyUxPMdoAiysnBvTwlLzna+guB18Rgra19CL8bPGI
r3FpeHnaPTsIPZg2Jbb9uyBHklP5uXyWucj7HTaf6/Af0KI1KHhY4hzwgIMkhcPA
R6pIZEvEklz1nqNEPH2qIkgFmVA7Gm75TPGSXldQwP5h44IzJSy7gONOlx7Wm5kL
UUPDT35EZ3YA54AmjJRvFxphfU/xJiDeEnavV+tSEuZixoPU5IGLvGwPQRdxjoOO
C+D0CfbLUm4NUnIxPctL7kuiAZF4NT2+70dtuOhoi3DyXn7RdOb9R7mbv0quATfC
WY0PvIROMqTLTdBjPwfhK2w3C7lGwXDJSzoGW0CdRhxeVl4p/KRKUgUQS/u4Ii09
3s+2JN7JxdFUzSU+nI7CH0zz9phpRuzBO9XywFhfl+nEpuVjv2lRo/72Ic+xOJXm
1h6tHf0xI9SsOSo+bSDxgWxTYl4XKSkuu2yCKDfxMRy9n+wobVlmNluD9VGce5uI
3KusK5NIED8fIuevRYaFZbt2l9uP1g8DGRFxZ2PCyh7C+C2MvJNIX1lzTpVfrPA3
mlOpAGuJI/2f6mpyXDuYPQ3ydSTD1mbAfg+D6eLToxuWX7mBFcn9AUBIKaeckaIF
v8QbKzP2YVRtK+X6DFxoj9xKJzRbg5BMwH7MEsY6L9Q/AUYusgKHb5I22/L/sJAk
BAcSoUIzG+LtOSKLWBjdBRzoUBWY+jPEnCz21+JplYSQ2SSqL+2qlbCYJ3gFfCkt
Bo7NMzDYYFK2youdo7diE1MNuLZInD0UrpkauvNqdrlajHyu0GQX8vjOr4SaYoVR
bdE/TVS/zohQRwyOXE+oYjOZJtheQB57QKZIRgadvrg7+ORVtT3yIjPSuQTIlOy2
J/7H1JLOSsZHLg/SGDTHypQGdcSLckLNkZtk2npv6LP8XTCGlQkfNcfAiQqyWjsP
2lzLfZCMhLbADUFLg/9rjEJRoHr6qDpYXNYfqzRhgV4+XZ404BJaDXkC2Knj6mse
unYddeB/goqlJoe2EXRHL1QwyYP9sRIWVImSx72hiA7rLHGsonqKYM7O6c2gK8HQ
1tnGVlqoH8BQzIw1u5iK5bY37DMpCaGP4JYWOQM5LM8MIWQGOp3i+R9wdyixgO4r
XHeIFd4aRmih9cv7T59svPx6gui94X4L4tUmiIg5NYFaKHhCj5oJfo7SubwRm0Fr
XThgNNRoEymOobzylC3fysebBIwJhcSPHeaG8vWBdiHdF/yXaQNa5hL8b69F1pAM
wIuWrDlwUUCpAdMFZEj2UOAMDMfs0VqnmHZvEW6BAqyLgQ4YIQtgYRochQ/TdB/R
c0gFmOESz45s9dojOoMhjLSjwK6F6ktMhnw+QKL7/Fc4IQyoSJvIt2hONFYSzHDC
Fism4mJ7LrGnWZzpQFJe+wOcqjotSTUDmLXq+sbYOi0p3IPYheqf1QDYrJx67MCv
BIltmvdIuTd5YHqgl1xs8jamRw1WJliFbQ02jQH/F5WmMh+FmVarIJmYkmAcSxYc
5fONxcGjLmnAucWYdBb6WXDsUSVBdW/bAMr53X1iBICBhZP3hpUND3oiLiU4myJB
DlB+zVGPubUA0QgUYXVV+U6/9YFsg+b0fnr+gQ+RE8vQNi8bgX9yfbhTyTBPGcdg
YlsWGMFA9Fv/RuHDoUUVY2srldJ9vKr/d3yVfEVSCcJ7XVoRAnh1knlijdYkdcy/
bnbuBAaWUztIOaXt9Q7I4z1niLTJRsJ43TjOmDeuHH/9bNESevmJU7yFBrMu13EZ
lflZMTCPd56oE6wJm262IRQAeZxf4jiICj5i0AfZm0kJbUcN1+Y95SUrTqpHWXaC
ganY1Yd3csNxGQzJE6pIfZVY4nlqLmBDDV1LtDQV79oAqgMGzvqXOCiNR8YxKz9g
4CH6B93R8ASRMdjpAO0uCecVuo5+V9x1TcMG8ATBmIJRb/d/suef79TsZkptrdx1
lUCIJVCK0LGDhSDPcT4WPGc87JU5sTUHdb8crbU+EbFPWN+iRJI+FG7q3mNM4IBF
N6uxzIU7RnFjdX71rCxP7ONM09teiqkAdzd6rW2UM2nM0s9jsY1KSs9vc2lqbpJg
7PWewCtGIFOjSFzF/StjKXyc9c8vFRiPhnW6u8Y5NeHslDxmjiKM4tlmEE2hdjlE
jX94I0q9gbaPSDnK5YZOefycPcyfLZOxX0HDdcfUnFsAw+XZcA+itmNaOFTdRvDc
VgCridgaB0Z6S05Q7HeS/UgRlezIUM7JXVW2GAvoKKaDj7B8/LL+rz0AZhOFHdqw
C4AF2QBthcZxZfT5VjyIGhG53NlMVJFHQ4LlMDQfZjHSX+PpsZirMRiEcsOKK/NU
31/MbnXsL1u2v5wk6LIwicecIMjeDvZh4cfjgkeyzM5gek78ncrnbaD+Fd+clrvA
MPkGIxTRyLWvUW4h59AgsPMzAq1W0+p/ih1XmNA4iTCD7m6Znd6U8evJe2JTppfa
JcqJTuDkoiaHvGo+z0vL9uApQ4RTWbN99vChkMxAChpfNWl/mLq5vGD7HoDZcOAd
RlicqQZBvnN9tnGYudn6xWmN2jvx1H+sqFa5czcC+yoE4YUXLILk8oCiBrvdXIez
6eydcqjCwZ1uhlYCtJw5DhPts7z1LuUarFTaw+dD8PVQSti3+RgQVJDj/JBVqzNV
O6ANVsQ5BheMbe6M4828a7uZi2Seu6PlUrohbkXCCxYxNEjpgzcdMq15MAetoG+R
kk47JsYik2/xzbxYeT6TuJnvuiwIj9XnAkw10PksK15diO+KsaF/z0zwi6DCvhDB
wTsukSJ5LjK2oe3AHbQCwjkTEYMqWw+qMdTssEFzhNR6VTNA2YaUh7rD4Kda5lY+
XUJlI9EUyQ9VbOj9HrOkuozHcddyh7SGtRk5I74KPo+wDGsIE31ieDz6cAfOp8Dn
B8apADuIBiksiygHk7zFxNgQV9rK3kam3T1RPG9s4p2O8abrvm3LG6H0D1Jy6sEY
QgdQXmtMVPBalbbFKgmLsjStueDpWJUYY3JNeZxxH25MmpSWu25XSIXvL6S8gvhh
/IPPf8poxiRKwx7bSJ7F3l0Z/sEXw8pD7Wb753Y1GKVPyK7BHaBCdsJ2NPphosdS
VTWrHs32upr0rdlRl+mf9GzlDPmHmjuy7pw3uxdpFYJI1SZTuxgWk9gi3ffQZRSN
kFyLeuAKAp7ra847y189IezIX/zB7a7hU7IyxfW+xduiX4d9+6OxShMPfHm/5sFt
PIduU3EEwvSx7FdCyyTfeutALcJM1Be1mUt0dQpR5t0Uk8uC1fIDkVqsisDLJJbX
XJrl8L3UlB6WEKVs0r1KqTG8hkHPZWezZe9yZw/68qpce9S7OMWgmnABPNnBpE1g
00kgdmNM2QYCmP8YgpPgtG9pWa2OgDtSglTaRxuo+UAGPsfYzcPGqwr5xq/tLEjP
mYUZlYzdRMQ7lYnBHLrDsYl4Fm6YxbQeRrSooIJwP/gn/sv0j645iXPAe8iSsO/j
9+EWgMV2+DgwyIOkzD3QSgsPhrY7XNqdPDtZA+e52AXzuBtgcbbtA4WwXm3gHbeL
tBQCm1Md18HqYxSLRD/zTDwqa7L/VxxSPxTEFSj46Qwa6MwWvGX7/hqRovtiS5zs
K/i+GOvWPeZ/O3SaOQePeEt8ul6A0+Giv8kTH6TXooY/d2HHFJwXxM7VeA5NSocv
14lzYWR4EY3yEqW8uz+7tRX/bNSVokelI4RAT7Vmn4ry+xcmUE6VilVqgq7dDfPa
xE3AT+NTEEj0WcAihx/N4Hs+qAzlf4khjlN0I4aK2YOiRx/2UhH1eSITvSPuYlWg
sXpLFehxV/hZQsXGYt0CUlhvnDQunxY0xnD1XatdIhJkNruw8Ac2AliHMWaOb2Gc
Bt+0VCfziO14Dw3cEHWdcPSwImycr/k9AgNWJapAgjXihpCXa2zijgWRnBXQkoaI
rarPG/NyFDrzGtZw1LkowL6ngmuA4rq9js+JpPdbDDnRrR2kQsJ2xID/SAdGpb/o
BfuVLIVlCD9PcfDjVkC/qKjbui56q459E/uh/OMvZ/okLsmEVHsj224OUSIaHwzb
RjOOOyNNZ/eyREJNJgwjL6hV98eorhdZiTWoTaxH4bqnrKp5UsPte8ybE6X1VmZD
Tq5sq/ooPyTyzI0lZVR577UTB6b6zsbp17ZQFDZkWFNkgb4UxulfHrclJLlbAlvF
X7drPkl+7THyI3u6WgdwbdY78CMm0S1MIz+GpiNmuhmgMrDnq584ffWP4BmGUZXN
83mfTLvjOhxc+PYq17laRyWNi3ZV+LjRWDDI/HUS4gz9vVWyL1coC1iZNbiYsphq
YLOz54pz15O+OBZESCp6NvfKFQDF+c2j36K+jnIn8jhCC6XNlFIvKlB+6K6oGS5f
cuslaAFZ2g4x6qPAM+AwhRSCIs7hCvpXikw15IZsX1rSTteVGJKjsYTYH4GV61Fb
Od1rqo23Xi84Vw+YeTxkjSwFRxEt1RhivD1M6ia+8/G/kJNNkgpOGMXHprfzW8d6
5fxOCld5bT4GOta+vYTzpXY7lSBpbrsWV0dk4byXbi9YQFctF7/aq0czXwd8kUml
6G5tb8obVxRJlVI+sngFmfrdJCBU+HN5z5qQX+DlKoK53gTGK2JHOsmxvkjhvjK3
Vh36fr1R1DRni8o5h8ZxYLT1nlqBtkR6YVkQrcwblVrAyv2qUdLz0F/BaUlTc73o
o8hU1lqDsCXPGQA1Tpc36Xj0y7XFnlUCU9S76838jpGR+ae8qdKR/p3yvioaqtgP
Jv7HUKsxH5v658Wygrtif9j+/EtI9w6rcD/nY5A6XYW9PRTh/UdJX/Y5OwhQp5Ju
m/rCuXHd7i3m84fPTXhDLo+LKyX/HtwpoVHhPbgoGWhB9uY2RB+PSNlatJ+ANEu0
6ftkzeG9GbhypQFuYy4J0but8kTBKNQTDbasnjHpakdKh7v+/QpCfhNZ2+O5t447
5ee6dJhCdVxHyzD2RGDfVRfsjgfiad+k7jyMCSfHqf8csYKlnvXJTa14XeJWt42X
dm9XZ1irB7dWNKO/cC1GXG4dYZpaVcooOBlUf7XSoDWQM70aqtmiOs/qdfAbV94A
BpPfC6St7IS+jNJtLP0jo2nMnwxR7Sd5fz06P67BKIqS68aWTC+X3KheRnVChA6q
Q2+Z8dy2RPF5FEUP30i968i8FBhJDbX0qBXhQ2rB5zTHiOrTXqHEI6Ew/G2WNESq
5LTIALCI6+BU4MWvI0uZQG9oNxMKS7UgXak+A5zRxq5OEF1p79WPMKTNflHSQ3ze
fOBLCZ5WvWr2nNCW/TOiLgJRFtpeYR/5gQ5dkdu7byll/2yBAR85sKVK2+rVWJEq
6kx8OdOB98A7jVITSvuQZeNXW0skFVnp9qz5Vyrr7MK6D8H7YRISAPYAUbjK6Y/f
XgzVblzHul0GPkNBFtd62RxdCsBXndBPev6+eZyh5PALZrGozKgJn3M8nPIIQi9j
NC+ahOJrrPO+6QmOMyY8yrNe7Q0F5Egs/zUwTMAKsjmKe3dPPygty9x4OeCqvNPl
qLeutJAJeSz2BAOCbcofctid83w8zzMzI6zxCFLUKs5SG+8Bjaj49uAAVGmE4QUW
VsylwNcNCo213UbPHHYgDmK0dT/g0YYK0H06B5/H+7lfdd8RijV8vMgiLW8EJ6fi
/5TkoK6MIHtQm5/hQFUfscfH9UFLZ0ijsUTLdGgKbXg/2epzi5MaWtEcEnb3hCmj
cgARZQPG47vyGhIlZQnlpR47HFMBkOv110JFEPV2MWMyPT9375OY97qxWJTrcHq5
ne/9+PlCErxXqWDXE1i0ZMMOV8GFthId6XUwQE3WoZoJ4cdix0NGbOEwM9wtcnUd
K1CJwtbVHlkrPFAwSSfGcVy/Ir07I9pWJslYibHRr23W6CkLq8zOQ/jAl3zl0YVM
IZ+r4vWQvYBNH7kx4UxMP8i7vJa/qUZCHTJ2rwy0wO66ccq+pCqBR+2m+VuRyB3+
ujYTkaSy61SO/0zzmXiye3BJV7LlRP6H7LH+O1Hib5+/q6fWVejmdsczKQ6nwNFb
8M71SwAIsYQAwOoTqS/111NWOHXDEwDiAN6FbVL+GL83d5jGe/K8hyIJIrBjBxUO
2rc8bLPIAADlWCyKJVE27zKVlO19keJodOnPDQk9Z8lGK9Dn12+Phcxd+Ee7OK4q
c/MyBN9SDuANxnBNPGH48rsbfcjdLMUqyW6GminPOjfMzegwUaVAroQbe8QTr64V
qQgCVMq/Q/YovjP5XSrNf9Ft4Zzai+cjaGGfXtoxOn5mvp0Dm6wwPFpuPMWFJyPF
yaD0bsu0pS7SHemgGhgkhqdVGvgGz77Ev+wPKS9pVlFeJ7kNRHZDSoiLPBf9fsD5
5jSTz21NiZkRNgItIUF7sODDNcuj0+xjkYRtE9cvS611tW8kNa7QuSL1Jm2BYQby
MCPy50PTKEX6GCjTEqXmUp/w6s9BWdFN1f0FmfyeMx4mhrLc8KwZ7R9BVDtENxio
G5cjJ9ecGdcH085Xt9niLFvev9WGXWV8qJkTGvQWETWH5I/GIH56oh7PvpI9FboI
4X7QA1vXEScVvxk1pKilYOUoFiQl2P0Cc5W0NBx1kO/HNcZAE/ZV25rhwelvys+r
7H8EijaJD8U62cU/SvL0AZdhZ8e/q21p280CyjT72zqLHBMOqRHOzDEwLMfqca8Y
RPLz+sQOgUWWcNnKynBdyQLXuv6k/88vE8g5GsqUe6+Ox/17vw5ZajW8onjLcNFe
4icJOOVPH/VVfOrGxzCbESM3uq225TwFAw1xoAdhZew6UWoUAkTpwuzeOJPxmt24
wTacZz0LcjxlcNThi2pRgNGFPowMsyEaFfyAKY1sKSdlSJv1thgjCqytdYZUh2vd
X4LWOmdpi3NYY0DR8EnJK3/Et0/B+hTpuMi6rM2I3NQEpjoB7ELAVmS97Ufumz3O
nyc8WHT2n7XIVcwe0+50QavPxAu1BgsJsAAWkQ/IhDnJyokn0E9LxpOGy09POBgm
eORG2KESc2hj8F+NoOsjHzRxFx+nzVn7qTI1xzxvRisvXma7JnpM2a11Nv/cIPkR
L0SVZszFtJ3VVeGYRdlJt0mp4P44zBgmLBQF4ULZBCU7tTGbdMQB+ewaDS2iehfD
Hbx2xMrn316JKOCl815Bhf2VnVbJF7aiohIIGkJ/U4C1KnqkBOW4NSkVYQBAaEea
XeO8fFVwvYXHkDJHhu2yqagP7ApLTIAztNvYyjV0FO5hVbvzxHMF0Ne7fO0LDtzX
HE2Lze/XTorjFCJ/CxY3AN9cbQ11yOGrRjQay9BdAQJv+JrIYDfPgbGjC3ro8pI+
2n+i5ldKI4i+2+AMKcsGnyEDwa4u1mSc5fIO7RGBw2kKMAuwzUUgTmvNJCbF6mCw
JESqp6frNRD7ywwqE0juFrtnjVwjCj3cV794Dd/6KIBj0MfOlMsuJUEALEOpcDJy
F6w2OiX4BAtgM2CUaXYj2g/VMek4rKLh5D6RNWTd/hDeFbxzCPdHeT+IHSBAsW7I
09BCuRAssTzI45cG8lVR3JQTRE3i5CvOguUUi2Nhhrxi94djONpqUPBmnWc7XHCG
xbEB7SWxHTPDAaHu3vESLU2BXS/WCQyKR38+LAPQsLRqncnXn7QR8esTTd5OLRfO
WhAfycXrv+rQ2VMPOOaaH585TOWabpLUrniZ8bwfemCPf0+Cv1lH0q8x5BW/86QV
iEOMAzi22EcepBx2qR6ucyW2ujgy1RecrOcuVDX1lQD/pSbr2/fxpz2A8Xt4m4UF
jBdRqGxIBCYxiOhtjosCpnOz5mEBjKDdnAs72hPVIGfUjQvfWq2r78TV6RPOEXyg
13sV0nfOEApuV/OAx5RaRMzpkykZryTqFqEGGY9RcyJgiQARYjWSLTsJ6nlqeBmw
1e5qdA3YzKj7iAz4FHSh+MRM6YxKO6TlrJWyy/cfib1FlCd564PybKslTpLOR8tQ
lHuqLrGyKTqdhkaVPTemqOvo/SlPpk8VagtdNnT8S5PzAvv2dqzRAFdFRePMJqsW
q19aFrXKH0kX/FPHiX3cHgUkKAMqgc2os/Vn4yz/T3IrNV2bEnp1enMCn3hh2wvO
1dX4fQzeT6+Rnd1JgxRQ59poL6j3S4acbs3Cwj64XTJXTU8yY2uXv2DHBrnke/Ob
KTwKxMJ6koser8NG//BYxElOArUj5jaycxw3nkUu8xybXtGhgDAfhoQCgtqzUCaf
LJWro1cDuS9MK+WDxg94RGV/UiIzT9PdRyR+AA4JDC32VvhSQOgaGxGhzF+q24QS
ECe2ewDYjtlOEvvPMQEi5l4slnhBIQtkw9m2kf4YPRIdgWKx/dOg4mXj840XqRVq
3Zc8GX9ZcqCMnOww72OIGlEIx319q0dkWs1A+GQwqrmbgYwsX6WDpOpXMTYwMyrY
hzxiD8ZxXqG3khlPH2MNASzomuBfyf0sNgIQpmEzz42Fob+1LHZL2n92CXXy5PhT
Uc4HPZIBF3tWEVACbaDYoGUY7H/qibzyLRTQUFsheRp6U8fe4rPG9/Gn9pPDAlQu
JKE62agKtu3m56pIPf8bny3FT5aCkTGRvF8yKPgjjIRH8Gm/s/ZjQZazIOHLzkJU
a2fiUuyN1N5of3fSCQAxooLdnzblZFnu9IAYQltFHEKpbimv+Q/s3qJz78rF+ix0
AwTjiXUsxzMPmjnnmD75HhjHxSp+D8Yn7HqzMuV245LlaOKOGhKC0FAoaRvKDOQt
vuRe4Cy3RwvE6lAzRWjDMkzK5Q0kZVkok1Cv8deJlWnS63HpGdx+vucTXp2rVXAK
ThFKeJNSVAcNJKrke/NChiu5FXrVgIG7HHcg7T8U0ixtzQzuYDTThOEr+WhIZLwx
hsCgjCzXG2JV348hWKP0M6dwiHk3HxJfWkCbMiz70zApmXIb6hKlCrpt3hC0CqGb
I2Z6q9aDSx2mGEaHjen1s+QZLcUI8QYVLT3nOR0lI/c6Z3vKi/hsGfwVPHMd1LY8
wVibn4xsIiXrLulrLM7MLwCaB69wTznEKBffF7tUTs/PMzm3RacItz6rQ6fbRctl
76rq7FDp7MulkSGZfGmy2WzxiHe6Pj6fiNJpj8EoB91xoj8a4+CcSkngHRsY8jEQ
J/BJq50MymF6ib6eaIQpQrqQ2zoqjPXGzkS2sxFAIVpBXphDyJ5RRq9nF4UPhDP8
HXPAhiE0D8D8q0jGgVrQ6Puy6AO2fatuhJ+iYdpYImFyqapCME44/5iTap1GXw1k
q6SD5TbyXY5+/FFWy8T6Sx1AMvWQa8d9klGIfjQfk3j0T+HM1YacNzO9dN1ANX9g
5Lq+5wlMzfXc9DBZwuxZGiBlVRg+3tGEw1S0pKDi8rVNugkZUJm4eBcCaud40yfL
DOnwYHDtVaTK5bvRx+3qUhf7DucYjdRlBKofT7H1aQx74VAgF7E500XqtZvqJ98u
eT1usz6gKQ3tr3r8ah+r7ydWYuKr0igD5WJJN5Qz33oaZ+DFBgwJm75WziV3BjMY
acmYuQ4+idzMoYTvucNZVCAFYscBzeez63m0R8cbSENBhFj8aqcBOeq8EnqjyI12
DZTPJq6cIvS+wvpFTAREMridtXYBs81ULMfEEExzgox1dY272YLTUgyzxqoW56K0
G1Ma3Pq3UNY11XgnqC5mtQPN89uuryY4nmczwOXCBHyhdgfQKY74BnIIwO7bKO0d
073aiROq3PC1wEXw8SRfFD8ZI8VsBLKFWzfVRNpy4kpvncAdTY2QAB/hks+Kwcs5
xjMEaQD4RfO2sfrepqCmf99H3F09OjZPFcdH/0CxJoR5C/4ARAUuKQFWwIT+sIPt
h50Hc4n0ZTRKZmMV+oARQMRjFCmMl3WTQdUuiP0co2Ujg/oDqoZ1vzIeaEgpuoUs
+sth6/NXJLmc09SQeuLcK9++AbcKemhHWMMbAosY6B21/xQ7qlTAYhNNr/P1KOm/
YzpYthzNLvgwUnAs1nrFzKb42c/3zT1F1NeyU5sfK4HLv6xGK7HogEvcaqD0QKh+
njGKZn8DHdXRu2ywoWClbsdekGFysMajsmqMlBEOjjmecpioT29sK565Bs89ZXjX
3GVOsVYRqdqm8xnIpBO79hanuuOrSVgkBxBOSeaC2qsIpIkubmvuDshQ3kwM+oYz
2GqlqOdC+DBWyMaIbZtWWgB8NT9HSorW+vvTTAvdz8ZzRwxbgBLRilVXf6Ww9rHr
4ulxEYzelGOHK0oFBqaaPcFKQU3EY4viQO+7Yaa7Xia6sLYGWdZWi9UvJiS2zUlT
jWkDIFxBZ1IU7OzS9CJ3XWKyQDIbiq4foiBaR24W6OQjfscSPN7Jybic1Gxsq9k+
9yh5yv/JXC/vdkSPxnf2ln6tIE7L9VVgYscuVB/eUrJtKS1wbfkJPj6JtuWYfTv5
t1cSg893P1N/RYZp7QFGa09VLF1qMzmPbkBgxSx30QKSSpGTjmhVMhY5BpZUEiSM
gn9zszOpPw9NjqYdDALvsWvJ60151P1P/Gzi45Vmu4J8sK98n1nxc9o/49scngAs
fYl1H0vZxbc+UIUyrDrOkNmnSoLuU/ntuQmfVzqd6gyFu2UfLJjHU3yh4nP4eZFb
I0y3lXXppIlH3PYjRZDmaUMUv6/49vIKhfVgQbMRzbPW5UPPEp5kZ8U9PVudpzQx
Ox8ykpvfwj8wU2lmtTwr7Mxa+1yUIDu9l8SCTYHK5zEatjAGzIm1T/O2nPCfzEQX
PHghhZMLet42mfcjPmIJUCEiIfzT5n/Uv9WQouReNjQxIe/0GlZStbYP5z3S1PZf
huGDcOJ49OdOg2rS2pEQbuUX2Asj939XHmfA77QZeq1S13OrKOMyIcVwFbRTjo1i
Eu4RDl3a2nU56rljAEXMyIT7yyOoUS82x/XYBCMU2Spa/JDP8KNBOYahUy+ITE9w
Hu29YwUu1dWDtdpRV5/uA2D8hxEDD2qSoqgaUPe/t4N1uGwMymRLxlR8rtg/yqeM
rGl/VeQnRjNvYZ7G8aSKQM8ZD+6YtBL8cdy824vJZvr6sdR0Aiyo4AhtKGn6LCV3
v63NhbbXh2IJzYkiV6IsIuRwlGj9RHoakrl0mEPsR7DFhK+9fRT2Gua/hu84gkVk
EcomV9imGS/UXeefgZN9eaoydY7dHLCrI7qzTCFbBsxygogUMfvjc1Oz4Mhjhiw6
buBxbyTT1K6OvwyJ/u6crfgxNuzuF2eU5HmbG8Weg67UKHsW9v42SM1b7jNJHKD7
3MVwUp2ux5afLMWZdA19ZXVbS1U/Yp9HhjxrwNNInF512QaXc5Nh9v29Di2jUyio
pwcUzmuuffdrwUv1KoY5dOG1kLoyrlUhZKPi96hSrHp+UtAHqxT/EHpcOEoiD2b7
`pragma protect end_protected

`endif //GUARD_SVT_AHB_TLM_GP_SEQUENCE_COLLECTION_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
j+g1OhsnylANQ2Tok9LZnrkmmjVq9V1RURg+0JCR107axewQmi4NNW4e8bcC3pcY
n9ZQd017+LBWwnvMuVWJ/AFXpuWKWePBvTpdWWrNPZiTaQeXy4sP1EMWPjNegdNx
/NhEZPQNBYcSKX+hngsM/BSGPl1mDg8KFmtq6lO3Ynk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 22724     )
wCJ2ri873ypzK35ZmV59TgPEUlwSzCWj86DoHb704D8L084vIKFHA8g79LtzyYil
zMEGb35XjyHiY0n1hXxT4FiYmuU1TkzKjMn9lq/RUzsz6Gj3TmUuOAQ5xJkgoZYm
`pragma protect end_protected
