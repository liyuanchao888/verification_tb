
`ifndef GUARD_SVT_AXI_MASTER_COMMON_SV
`define GUARD_SVT_AXI_MASTER_COMMON_SV

//vcs_lic_vip_protect
  `protected
;?.&@^.T4)EQ7_ILF-ER+_P@C;93<C2BbX(F&:;ONA2,4W:C]KD.)(d2b\)O)F_6
JOMZ.RL,1gW:.TT=TGG23V,;bZ8SebEUI]L<+U+5#9_\WTLeM.Tefb0-1]32ccQ.
19K+Ee<(LYK4J&.(.&BcCg:d)[_XO0LPQ9JKHbScMPF<A0+;D.[=\II@Yb?9U1S:
YXP.[G.HKKfF^F[3:gU?-c4V>/TA>c]?_aOM/?cG:P,;W2DK/=,QFX,JWCMc-:]Q
I/3]<D&MGaENT2Z@bX&c4N,Z?HT.P(7Bb>#5QNKDOGG:SK:RJK0gU97IWJ0FVg^J
Fg_R0,C\Y]3MS:1a[]>8+De\V;OGg-1Q46gWc/IYX^1#+Wdga(L66Oe>2ANa.fG\
]/A1I&1a1;P/7-+I7-.\g:8NEADDQO9\[<^\,SgB?VA7X-5W^E-WX3K52Q8<MGXS
1DU@H0,W<+->DAJ0]Kd.:APK-XJ9O?G=Z@JHA)Hb_WIK4Z9\WOH_CPAUTf.\HH)B
\.P<4FcGT;J9?:G(CT^G:1PZcW:MbWA:JETOR:B)RW0eg4X#WZ8;@fI_\9=T/aRU
09_fU/5R-RAO>bQTSUfg-EG&DcdJ+a0>;PAA)I[d59R=.1BW[U[eaW?f0Q_CHLNV
P:G0.=RU,1f4@3\P&3X2^B27EZDHHJ^fBNOTR4W2X3Z?McScK@@;]-<..FL/H^c9
6]XCFTP/VM\C>:g8+FW<H3McJDA7@8C&&)bb7+T#^N;QZL<[.aTK4Ub_&2HN-E;\
UW)X@\7/BS5cD;BO/cB2+[AOXPQ36]R,)TZ.98I7@#WNH=;GOEa-(DCF8&7V,KVW
cLQ]MbN.#ce\TVB3bNPa6T.:dTJd&[WCcR&g2+>5)\?P[>OFIc9.RI_FO9A#<VKW
I=USMeY3JA8\U/dR5.-#3Y##6@W]1eHBOEB.S(OVOJb(3S0?.-S.3,IXg6S]b@DW
b&gO+8+C5TNcFb/4.K)5AN^>VN7H8V?FdC+X)_<]aL//\98d7(R_<Of@5.60_MQ2
cSa&]VOQ9Q?7f-C5ZU8P#4<_9TT#EI9?-;9ZYDQL9A5((.T,&fNPH:-a,@;[-_ff
OHQE19;^-@HLf@,bF]Q<NH#g)LS@IQd5A5\E&G##JRKTPI6QQ:,\Ed)#@c)Q=^b^
(1-NAG?bBIS0T()3Q-A2Y>WS@5-8W:.Kd<83]HO]XQ_B3c9@EH5(K((8&VW/D]E9
W.NK/[I3e^O(<:2]-[/E.QD-V<?0NaDX6/eHX#&U1@YYc8.\Bb,/a8M^JN.9>)0[
d^1NB-Ed)XD-ZU)\25V(c4)]6@Eb1A-XQ:NU8^?;RA6cXDW<dc_[U.S,0TTe@5;L
N/>G,.R.S^KZ&bB9^gg0V4fZ(EJ7QLeg3>VJX=W[KL]A(/M_K#S?;B]5\0JOV7XA
^./,g(gBQB=.>V1Xeb&G\EESB-.EfB)6Dd_0H164AO(L+GBEY;O):Y:6YV/[#.Se
dA@\=+88=fYH7)4Y+eFRU1L+g;(\3RVCVB5G\F^00Sb)(He[d[;>9MTa^J)FgbM5
-90?L&f[MX>-&G6M]+Ge[d(3L^#bBLV,;8J20Kb_,b9L=d,I(E(1)aWH>1?T[&S)
cJ^15WE_[K]ePCTb?OU.M;a[]e^8[;g3e<#Wd?4J4;2LD$
`endprotected
  



/** @cond PRIVATE */
`ifndef SVT_AXI_DISABLE_DEBUG_PORTS
class svt_axi_master_common extends
svt_axi_base_master_common#(virtual `SVT_AXI_MASTER_IF.svt_axi_master_modport,
                       virtual `SVT_AXI_MASTER_IF.svt_axi_monitor_modport,
                       virtual `SVT_AXI_MASTER_IF.svt_axi_debug_modport);
`else
class svt_axi_master_common extends
svt_axi_base_master_common#(virtual `SVT_AXI_MASTER_IF.svt_axi_master_modport,
                       virtual `SVT_AXI_MASTER_IF.svt_axi_monitor_modport
                       );
`endif

  typedef bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr_t;

  /** Event indicating that cache is updated post snoop */
  local event ev_post_snoop_cache_update;

  /** Event indicating snoop has been added to queue */
  local event ev_add_to_master_snoop_active;

  /** Last acvalid assertion time */
  local realtime last_acvalid_assertion_time;

  /** Number of pending (waiting to be added to queue ) WB/WC generated to transfer snoop data */
  local int num_pending_wb_wc_for_snoop = 0;

  /** Component full name */
  string component_full_name = "master";

  /** Time at which an address was invalidated due to a coherent MAKEINVALID transaction */
  real makeinvalid_invalidate_time[addr_t];
  
  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param driver Class container for the signal interface
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter, svt_axi_master driver);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param driver Class container for the signal interface
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter, svt_axi_master driver);
`else
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_axi_master xactor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  // SNOOP PROCESSING RELATED METHODS 
  // ---------------------------------------------------------------------------
  /** Adds a new snoop transaction to the queue */
  extern virtual task add_to_master_snoop_active(svt_axi_master_snoop_transaction xact);

  /** Removes a snoop transaction from the queue */
  extern virtual task remove_snoop_xact_from_active(svt_axi_master_snoop_transaction xact);

  /** Receives snoop address */
  extern virtual task receive_snoop_addr(svt_axi_master_snoop_transaction xact);

  /** Checks the recevied snoop addr in master exclusive monitor and resets it if there is an entry */ 
  extern virtual task check_snoop_addr_in_exclusive_monitor(svt_axi_master_snoop_transaction xact);

  /** Sends snoop data */
  extern virtual task send_snoop_data(svt_axi_master_snoop_transaction xact);

  /** Sends snoop response */
  extern virtual task send_snoop_resp(svt_axi_master_snoop_transaction xact);

  /** Drives the ACREADY signal based on the delay */ 
  extern virtual task drive_acready(svt_axi_master_snoop_transaction xact, output bit wait_for_acready_end);

  /** Gets the delay associated with snoop data transfer */
  extern virtual function integer get_snoop_data_delay(svt_axi_master_snoop_transaction xact);

  /** Drives the snoop data channel signals */
  extern virtual task drive_snoop_data_chan_signals(svt_axi_master_snoop_transaction xact);

  /** Waits for the CDREADY signal */
  extern virtual task wait_for_cdready(svt_axi_master_snoop_transaction xact);

  /** Deasserts the snoop data channel signals */
  extern virtual task deassert_snoop_data_chan_signals(svt_axi_master_snoop_transaction xact);

  /** Gets access to the snoop data channel for a transaction */
  extern virtual task get_snoop_data_chan_lock(svt_axi_master_snoop_transaction xact);

  /** Assigns ownership of snoop data channel to a transaction */
  extern virtual task release_snoop_data_chan_lock(svt_axi_master_snoop_transaction xact = null);

  /** Gets the delay associated with snoop response transfer */
  extern virtual function integer get_snoop_resp_delay(svt_axi_master_snoop_transaction xact);

  /** Drives the snoop response channel signals */
  extern virtual task drive_snoop_resp_chan_signals(svt_axi_master_snoop_transaction xact);

  /** Waits for the CRREADY signal */
  extern virtual task wait_for_crready(svt_axi_master_snoop_transaction xact);

  /** Deasserts the snoop response channel signals */
  extern virtual task deassert_snoop_resp_chan_signals(svt_axi_master_snoop_transaction xact);

  /** Gets access to the snoop response channel for a transaction */
  extern virtual task get_snoop_resp_chan_lock(svt_axi_master_snoop_transaction xact);

  /** Assigns ownership of snoop response channel to a transaction */
  extern virtual task release_snoop_resp_chan_lock(svt_axi_master_snoop_transaction xact = null);

  /** Samples snoop address channel and assigns values to snoop transaction object */
  extern virtual task process_snoop_addr_channel(ref int acvalid_to_acready_delay, output svt_axi_master_snoop_transaction new_snoop_xact);

  /** 
    * Waits for a new snoop transaction. The monitor uses this task to get a 
    * handle to the new snoop transaction.
    */ 
  extern virtual task wait_for_acvalid(output svt_axi_master_snoop_transaction xact);
  
  /**
    * Tracks suspended snoop xacts and triggers events when they are ready
    * to be added to the queue
    */
  extern virtual task track_suspended_snoop_xacts();

  /** Gets access to drive WACK*/
  extern virtual task get_wack_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Gets access to drive RACK*/
  extern virtual task get_rack_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Releases lock of WACK. Decides which transaction should
    * be the next owner to drive WACK.
    */
  extern virtual task release_wack_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /** 
    * Releases lock of RACK. Decides which transaction should
    * be the next owner to drive RACK.
    */
  extern virtual task release_rack_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /** Drives debug port signals for snoop data channel */
  extern virtual task drive_snoop_data_chan_debug_port(svt_axi_master_snoop_transaction xact);

  /** Drives debug port signals for snoop response channel */
  extern virtual task drive_snoop_resp_chan_debug_port(svt_axi_master_snoop_transaction xact);
  
  /** Drives debug port signals for snoop address channel */
  extern virtual task drive_snoop_addr_chan_debug_port(svt_axi_master_snoop_transaction xact);

  /** Checks coherent transaction. If data is available in cache it is retreived */ 
  extern virtual task process_coherent_transaction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Deletes cachelines in the address range of this transaction */
  extern task delete_cache_lines_in_addr_range(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Reserves an index in cache for allocation of this transaction */ 
  extern virtual task reserve_cache_allocation(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output `SVT_AXI_MASTER_TRANSACTION_TYPE lru_xact);

  /** Writes data into cache */
  extern virtual task write_into_cache(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Updates prot_type and memory attributes in cache based on configuration */
  extern function void update_cache_prot_type_and_memory_attributes(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Gets prot_type of given address from cache */
  extern function bit get_cache_prot_type(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, output svt_axi_transaction::prot_type_enum prot_type);

  /** Gets memory attributes of address from cache */
 extern function bit get_cache_memory_attributes(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,output bit[`SVT_AXI_CACHE_WIDTH-1:0] cache_type);

  extern virtual function void get_end_cache_state_and_data(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,
                                                    output bit update_cache,
                                                    output bit update_only_status,
                                                    output int is_unique,
                                                    output int is_clean,
                                                    output bit use_cache_write_data
                                                  );

  /** Assigns initial_snoop_cache_line_state based on cache state */
  extern virtual task assign_snoop_xact_cache_line_state(svt_axi_master_snoop_transaction snoop_xact, string kind);

  /** Assigns initial and final cache line states in xact based on cache state */
  extern virtual task assign_coh_xact_cache_line_state(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, string kind);

  /**
    * Randomizes a WRITEBACK/WRITECLEAN transaction to transfer data
    * for a snoop transaction
    */
  extern virtual task get_memory_update_xact_for_snoop_data_transfer(svt_axi_master_snoop_transaction snoop_xact,output `SVT_AXI_MASTER_TRANSACTION_TYPE memory_update_xact);

  /** 
    * Updates the cache based on snoop response assigned by user after 
    * receiving a snoop transaction from the input channel 
    */
  extern virtual task post_snoop_cache_update(svt_axi_master_snoop_transaction snoop_xact);

  /** Waits for post_snoop_cache_update() method to complete if any activity
    * is observed on the SNOOP channel */
  extern virtual task is_post_snoop_cache_update_done(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit check_outstanding_queue = 0);

  /** returns the delay for RACK signal */
  extern virtual function int get_rack_delay(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** returns the delay for WACK signal */
  extern virtual function int get_wack_delay(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /**
    * Checks if a transaction can be given the lock from the
    * perspective of a barrier
    */
  extern virtual function void check_chan_lock_for_barrier(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, ref bit give_lock);

  /**
    * Checks if a transaction can be given the lock from the
    * perspective of transaction ID
    */
  extern virtual function void check_chan_lock_for_xact_id(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, ref bit give_lock);

  /*
   * Checks if a transaction can be given the lock from the
   * perspective of cache maintenance transactions
   */
  extern virtual function void check_addr_chan_lock_for_cache_maintenance (
                         `SVT_AXI_MASTER_TRANSACTION_TYPE xact, 
                         bit check_cache_maintenance,
                         bit check_memory_update,
                         ref bit cache_maintenance_in_progress,
                         ref bit memory_update_in_progress
                       );

  /** Checks that a transaction can be given the lock taking requirements 
    * for snoop filter into consideration */
  extern virtual function void check_read_addr_chan_lock_for_snoop_filter(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, ref bit snoop_filter_give_lock);

  /** Checks if there is a snoop to the same cache line addressed by xact */
  extern virtual function svt_axi_master_snoop_transaction check_snoop_to_same_cache_line(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit is_snoop_to_same_cache_line);

  /** Gets the handle of a snoop transaction to the same address as that of a WRITEUNIQUE or WRITELINEUNIQUE transaction */
  extern virtual function svt_axi_master_snoop_transaction get_snoop_to_same_addr_during_wu_wlu(`SVT_AXI_MASTER_TRANSACTION_TYPE xact); 

  /** Checks if there is a resp to the same cache line addressed by xact */
  extern virtual function `SVT_AXI_MASTER_TRANSACTION_TYPE check_resp_to_same_cache_line(svt_axi_master_snoop_transaction xact, output bit is_resp_to_same_cache_line);

  extern virtual task drive_wack(logic val);

  extern virtual task drive_rack(logic val);

  extern virtual task perform_cache_update(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task drive_rack_and_update_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task drive_wack_and_update_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task process_ace_reset();

  extern virtual task pre_process_coherent_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,
                                                ref `SVT_AXI_MASTER_TRANSACTION_TYPE memory_update_xact,
                                                ref bit drop_barrier);

  extern virtual task wait_for_xacts_to_same_cache_line_to_end(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,output bit is_xact_outstanding);

  /** This is a blocking method and it checks if there are transactions pending for the address provided in the argument -cl_addr. 
    * If any transaction found that is not yet complete and overlaps with this same cacheline address then it waits for all those
    * transactions to complete first. It keeps on waiting until no transactions found pending that overlaps with this cacheline.
    *
    * @param cl_addr Tagged Cacheline Aligned Address for which overlapped pending transactions are searched and waited for completion
    */
  extern virtual task wait_for_all_xacts_to_same_cache_line_addr_to_end(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] cl_addr);

  extern virtual task process_cache_maintenance_transactions(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,ref `SVT_AXI_MASTER_TRANSACTION_TYPE memory_update_xact);

  extern virtual task process_barrier_transactions(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,ref bit drop_barrier);

  /** Waits for barrier pair timeout */
  extern virtual task wait_for_barrier_pair_timeout(svt_axi_barrier_pair_transaction xact);

  /** Timer for DVM Complete on read channel for DVM Sync received on snoop channel */
  extern virtual task track_coherent_dvm_complete_timeout(svt_axi_master_snoop_transaction xact);

  extern virtual task pre_process_coherent_exclusive_transaction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact ,bit is_unique ,bit read_status);

  extern virtual task wait_for_write_xacts_to_same_cache_line(svt_axi_master_snoop_transaction new_snoop_xact);

  extern virtual task get_mem_update_xacts_to_same_snoop_cache_line(svt_axi_master_snoop_transaction snoop_xact,output `SVT_AXI_MASTER_TRANSACTION_TYPE coh_write_to_same_cache_line);

  extern virtual task trigger_new_snoop_addr_chan_activity_event(svt_axi_master_snoop_transaction snoop_xact);

  extern virtual task wait_for_cache_update_post_curr_snoop(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit is_snoop_to_same_cache_line);

  extern virtual task check_chan_lock_for_outstanding_snoop(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit b_has_outstanding_snoop);

  extern virtual task update_current_snoop_xact_handle(svt_axi_master_snoop_transaction snoop_xact);

  extern virtual task include_dirty_data_into_xact(svt_axi_cache axi_cache, `SVT_AXI_MASTER_TRANSACTION_TYPE parent_xact, `SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit original_txn=0);

  // This task only resolves dependency of stalling snoop response with memory update transactions
  extern virtual task check_valid_snoop_response_before_sending(svt_axi_master_snoop_transaction xact);

  // send CLEANINVALID transaction when cacheline doesn't get updated due to error response
  extern virtual task check_and_remove_cacheline_from_snoop_filter(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual function `SVT_AXI_MASTER_TRANSACTION_TYPE randomize_dvm_complete_xact();

  /** Checks if a WU/WLU transaction is received from the sequencer while
    * there is activity on the snoop channel. This is checked only when
    * snoop_response_data_transfer_mode is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC
    * Needs to be done so that the WL/WLU does not get ahead of an
    * auto-generated WRITEBACK/WRITECLEAN
    */
  extern virtual function bit is_wu_wlu_during_snoop_addr_activity(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** task to sample parity check signals and calculate respective signal parity values for parity check comparision */
  extern virtual task sample_and_check_parity_check_signal();
  
  /**
    * Waits for WRITEBACK/WRITECLEAN generated for snoops to be added
    * to queue. Applicable only when snoop_response_data_transfer_mode
    * is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC
    */
  extern virtual task wait_for_pending_wb_wc_for_snoop();

  /** Gets the time at which an address was invalidated due to a MAKEINVALID coherent transaction */
  extern virtual function real get_makeinvalid_invalidate_time(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);

  /** 
   * Adds the transaction to an internal queue of transactions
   * got from channel, but not yet added to queue. 
   * Blocks when the  number of outstanding transactions is
   * the configured max. value.
   * Checks for ongoing snoop before adding. Internally calls add_to_master_current_queue
   */
  extern virtual task add_to_master_current_queue_post_snoop_check(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

endclass
/** @endcond */
`protected
P)XCaB&5P0>QD#Nd0G(Y[3FTSO,Y08<VXA0VK(ML:5.J,XI8/=ET0)T6N#368Q>S
@]/UX=-Z\V+J&,5bSMI:@FCW_dR<A<K\O6/gFD9f#=3M>Uf?EQP9NC8?g&Y#T5c5
D8^>=XSI7F,]K>8U84QA.PW+JWGHECI\-M\OQe25IdbV,?_D#g/R?86[Z.:IS]M.
0BMbW4f4.AP)(4QBeO46B;<>@;WN8QF#2W<c+&2cd,5@N>E=e3HVFWL0:bJW0ZSN
e0bVa:BV7:3b.GVe+6PQabe3Dc&GT5)A.[Fgb<[AQJaP)TNG7)Cc1\FM=4;5H+fX
YGOJ-9(]36U]-cIA&H74d7=bc44EZa3<6CLGQBe^DcC\_Hg3T_,+I[?QLa+YU1XU
HCI8CNN00a>TVPNYQT]F1)ZR>T;3&,::O>K0)f(R^5,a+a04=?e;_R;8#Og-PK)B
SF(1A<JZD#c#GQC]IbP>C[F/,aR0/F8:Kb1GdT)0f-bb8a+=e[NB?\fNOST7Z;,Z
@aB0[M&I7Y/g_Y1C];/E+IA\]ALAabIJI48QG.@PD=S8=GE.<RC:Z]I28^bfG4?d
K=@S5d;dM]N0705aJJgJ2SN,#CWFYW5WF96S<ARII+/+#b9O::,WaKe\I-I^^N@>
F3)_YEX?WQ?P5e5IPZJ\2OTd#_N?3]OF0CJ9#^_bJ\c(;cf=[1.I;I4=]MB:G?0c
SQa+;V-5,SI,.M.(VZ3RB5=;ce#c3(=\:S8\X1f7OGSHY\F\M@3K+42:#^^&f6[b
^8IN,+AT]FIE85fWBgJ7I9OUKJ?0_9(d5TG>C7PS.[BXAVcG,<Ue\fXU;F4L?S8=
51/G:ebJ6_UECE;6A31PgNQ#VM.dccL#CW\TG6-6&cO[9_HJ;W(H_5O?8CCMJ+H_
.=>JbfL7V6Z:[b1(5N8H^=5P[-7B_O_C>V)DEN2PJH)NVAV_<&R&[A25SGdKA<be
7b@4TWVfLIE\MK44_8QbIYZC4eRBJ.>FdDPWKfS\8,P]CK:5^RVU:?8#+I9c1WF2
g9C=5#&/#^;4LGC]@7\/F:UQR2]aE[M+WQM1L+XJf)/O#XCE=AOE&]^/EFT;D+_J
bZ8&GD3gP;6J\4[KdFLYR\YJL;fD6QK.DNIGa1GE]5PV3QUCWVZX,BE0R?6.:\^(
E]9C5bO&)@Ec(Le9BQGA5?NSDS^FcgWO]Jg@a714LgGeDJ8RCe+g[e^<g6(OFYKR
(APVUZBY\a;3gYD7UM)g5J[a)+&VfaMP#URT>--?+.D4XY?-@PW-dJGIN1@&M>7c
gXJVNAQTG8)eb1I@=B065VB6RgN<NX.8g2N]cXAaR;165PY8\?WX&1eD2M0AO9e]
5E+_O=_GX\dbPHB4BYL;4S>@8E]#N.bba2DFbSaI2JI6A$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
W?3[FZV6=4f11ILV6-X0CZDJ<-Y@eTU,8bN6R07KRZ7Q6#F(UN5+1(eYEA)JCH[f
g;;/Q[5RaW1<59g_8@J?_g<>_TT,Lc,YJ7H_/-9#R]M#266dJ>>1);1-Wf-L/53L
ANPWfDQEUMQG=854?>)I#EaJg?70(c)DGY\[TQU7ZH#K.1=^gQO_aE<dRIQGDO6P
RVJI:g0K7D&9[&8W__7d6a]9AeK_A;CddW;7?R<QNHNHf#B/#Hb<H,(U&@KWRH;K
2;)Y^,2D>-QA,>5)CD,d,#-SNR.&5VS.Y@ge?8dTbb>[7068[aV^N)5E[K[&Q;4U
fRAHVBHPa#[^5R[XE@9f.a=XGU:_<.J.9gS93(V\EAO)1:XgME_07;;g/KbRb:WX
?+#<-DaYaY<B,XH1@J#RS@#R.bS3C41P1=4+ebB^:LKWP7DOf.^OOV)H@/\X^SZ.
QN1)c,2XLIQ-@DaZ>fA<43\3HZ=P87DBQ3F4.1AGFa=#DfMR^g^.&-U?PQ.f+;(Y
1[RB&7cQKbNbg?HeD+J?fX7SGg(gb^Q1JY#<eH72NA;SFI@EJAe]9_O5a.ABScdb
JdBW)b1]HHEcAUI;1CNH_=9H1D4?N5^(g?<7K\]cE2\4[-aCN0d>0FdW=E>BF.Mg
KeEL:8Kfc&68@:fBd@5H4E5a]_7W(C+:dg\YP\-Mg.7;].==LedH&I24XFQV65\5
MFN:@]eXO:gabZW+\1PN6]FSSA2SPR:X^R[:1YPeDJ;8U]P0aKf)ge#)D9TN=2:3
]?L<+X)ZC1e->d45U1CL..I9O7c?EJgeIEcY3\+-Y#SNe^4_RO2K[LE3Af+]]OHD
H.,W@)CcL0P=T1PbG?G@)._HAJ@=R#(6Q=V45L)Ke2[X861)U)4Y<f9O1RB9b/SH
KJYF7#Y8]DRE52Q5A#X>bL(^EbV.M4:D(K>N(RZOX#]e3\Sa#D,^IK<W0aa-Wa;1
c)^,H&KG,P8cC8:DgX3YP<JYT04^-0O9[MX?[(#ZPMR>.BVTGOJ-S3^>S[_>B-DR
BODM;#7Kb;J-XFBN67DF=<e]g-7/EcZL;<=>AZEAB\HU-\2PLBg6Q#SGDOOB_-f#
5afKIbL0&eB[8[\-_c<&K3J8A-:C4eVF[VB-HgXE>6]Hg9FIBQ;QJN03AT?F]@K=
f5aafNd6UXa;>]L@?^G(&IRBK6VdW=&NF+;(&^Y8P(RML5YKc6K7:\J@QGJa06@.
(C&eZ^bN:P@U0R:6c-+Sb]TSMG8G\c.X&06LYP\@Xb7O&W;=E@HFgHA4PD#:QKZK
94)bg,M3(aOI46a(N[?F=f0D:RTd[^YE;A\B;>K#fe7-9<9af?6?4bK^c[G9+Q^P
>7.fZ#:TB7;W6_\=ec3ZaNf<..;:5a:UEE5(QCE]>]PcB\g\X9Kf<2bJL]#gYZ?N
>F4^^UMbJ>Q7b74<[ERSb9ZRHa2.:B7G9Ee1(f2B^UTYXX0G=[/;6OL#+Qa?KQ[R
YU@2]H1HA)_<ZK#eb4[Z;#TTWQ0d72#F4(3G>5GScYYA>05W]Qc266XP)B&.@JW/
c9U>fbc-FALP)bb&Q-D&#eMKRTA8FeHgR6a)\A=18.Sb)U9T,2/+>K>A>&R[c40]
acJ9557g4WD&c10+(>\]Gf<O^d8/90W\[N,AfTP:B>3D6[0N+f6FHLf[5bdS7^@A
\;<]8a^M<7g+B)R?ZZGg\3#0WS&OSEdGc^J(=7[48#=EB=\&Jg(6D,gT2aXZ^2WM
=<,eIO;O>7Z13C@/KHIM.eBL1@gBE;gdE[>#c56B?.,a3Q8UOQ\We=(3<f^F5eAF
#W>Y,)P\/eN2WO&1Q63U=UBOG+P8Mcg?T_V=CG3O[XQC_96Q)IVWP7VA.1eT8XH3
\7]Z)FM([d<cgONZABL/9gSY&TbbI=>4L&@E^;Y7MNDeCSP5VS28PS8:g)5N@N9Z
Ug0GA7>1gfaJ2L((&2dBg23XI4aE99/4YLT:<4^]W7I89?b5Wd;:P?4T<B3>2c>N
X57fR=>N5K&+ZOT7KA64(AE8[\;Y<(dT+X0.705:1]e:(cL[FKgeBeUA[3/ODSQ9
Z&f>d7GDQ>6O)CC8_LDc>A2NFD9O@\F+(H[[gdJg6)--4&OZ?-.#V70?)RKS<@a\
VKee3Zb03B5M./[Yf1</[<D^JTaDX3NLJ9d7-C-^/HV^BE(Ie]2F&#XJ-98LbS9]
Wb>4-GVPS\0WSO[-dRfYM,U<YQ,S<SMR,@Q77@([LRg3Bee&185[&E5RL]1D=HWP
@]<&g/@L;adcEFGW=Q,+ZESF[:e_b2R=/DM,S(?D\Yd&_BLF39?,F]LXBS1+B]0P
UPKHCJ6>K/JdTe10I33\7^DK/@1)3]R-9Z\Q/cGR3_HTRD;BA\V<UONeY=dbOf5P
W_3FN;LNE=S^5We5YO,6OZ<ARfbGON,gLY5F+)5a<4\3E._X7=87D]4R1HO.R6F.
c\1)FPP.G#e=.O]XT@DIRf\MCB2gP[5C32E>.YdPR^S1f9Ha&#3X5\Y-M/]>dMC7
:#[DJ6L0E9UZ5;F5W2<KY=U,gOH)^PN1WeOQC3/-OTb?)]HWZ)(PN0bV@_0]RdZc
#Sbf,.<Of-7RW5:;_2;dbb;^a>A.&]g,Ae?]:JY/>E:^XDc3>6Q6U+B46g8?]U.=
K,]cK<R2>cD;2RW)42BEdH2.1BLTBI1R\?0Qfb?f0XPJ(6Tcd(02gA6C3IAdS,0.
TZ0GVJ=g0HE?@&0>TF2AJ?4Y;RLE?-7afJ0T4.^:HGPFO59H(^39EN2(0Bg8c@bQ
eaAND2eaHGg?,$
`endprotected
    

`protected
;3)XJKMeX7O+LRO995A\NSaF8=CbKK.^4<E#[]eSg[cW7bB,;T6L2)E5<8QMZ,=F
@aY<6\KA,UK+.$
`endprotected

//vcs_lic_vip_protect
  `protected
S<[[1-.\:K3C91=@S[/>4?PW@FMJV-Lf0:\P6__c^<FbA,+?=eg+7(3K/egR)<>:
a?aD[g]M&8e2?Z9E/\G_>^EaX/:Q^882<9G)_JB#THK3;)LZ1X<3Hcb+=/5\7:?;
TbWJ;J9If[U^](>;4L1:H.^ga^<cVG[TUQJ-7,1I+T9aFNF2(VSR1W-Yb?Wf;=SJ
NBYNHF:I&F)]0Y7]#f=C-,-^XC/[aFX?^V<2QcIC^-UTVb9cCPXZ=NY\_OU#\^;]
,g6?;dK&(CD\c?W8/(0)M5a6=0Hef<JfOD<8)e[OAFRfBGE1\c8>I5UA@Y-I^M;0
V6,NT\D-BR=LS;;./1Pc:.<;_-:J.aDVc<_AXf?c5S21N(^^@\>(5&TT-K3XK8c5
<49OHXH/[<W(,392^Oc8S23W?aC#0L@,B_CRe^Z_W7.QY5\ZIc4UI,&4O1S=)Q4N
^PE)@eB&0U0Db7A=Pf+4C)VUD2BYNL_:aB\N86M[JYf,TfF,R2\V<P+G)PB97&FV
gKGa:SfdO&b&CBVU#(X24[]E\b_<aA>-A&)Z7RBG7PKY)<fc5844\39:DA<L.6<E
O[8:=//_SUOBCKO7&c2C+).I.60>QV>WT96e8a)3Af.<^SW0G0O>L8Aa6ZO5@[;[
HO6VE0.B9d)38C-Fb8g[3ZDA+RDKH\>@L;Vg7/2.-\<8&D2UI5FMHcKb7>+V)1-)
_BUJ,EaG>70&\b6^(V0Q+A=eSOLP5MC@+JHY[>eU+[D<,,X>4OMZ:Q?K5@Hf+8A#
SGJ5We@d,3,65HA.7&^A+/>;HMX9&,Rb7ff8ZOMVU8YXK0c8HcZ^^L]Af4EMc7aX
[fV9;R)G#35P&TcMHH.BYZT<3ePOL0X;I+#=,)Z6=LKZPf+;cc>1PMYeALdG#>VW
=..]/VKGWPJ[P.e+X^H7U4^0->=DTN4?,F/6N&3QHT:9^S[GZedL9ccYN:FM?AGI
>3FU9TBQfS_g2Y<Da;,2F1)[MS_@ZS&FR7[Q\J4-O:OZf3=>M7<BPC>-T+K@D3:=
=?e[_gd;:&HYdaU;V4^-PHR0c6L0MLQ&_e8;HWJ?7VL8?Y48eL=We@.S[G:#B?^I
aU]CN6c7479KS.@L0U-/<^;1OL[Of>#LcKI/d>dMe>d2M_678PJYaI?^]:,Q9GHL
>E//@S0Z-Z11LdRb[HQUO?/[;=6B8\D\dEH2/:_4)G8?[7;2XWGDS8P+NBVG<U>R
02@e@1Fg>CE6/,E&g>7N]\#JS8Y;),\cY4eZWOALUaD:f(3<R=V7PG9J^+DQC&@]
\Hg2(4V90WI^L/[.]IbOGX=U@M-+\>BRJJI(H-#XS[66=9I_Sg\[T5+MG678M,<)
[).eZ-1:>eJf(&.8eSD>NLG]ON<c5=4acG+)b[9Y@W2,7c;-XHFVV0Q?&PGA?/KE
a=[>=g+DW(-A/73]gB@5B58VeNE\C=49d;@>F8(.0,,,:9_N]B[1bdd,dRK:YB33
@SHL[Z#_.VQ?:KGaK\1L=bVa<Q_&^]DG#7bDU/X^8_09BY1dadBKOd7:^d<W1>[^
MQSf^AO1>KVN3d&#RRK^1XU>=<C7105fHNL#4B6Ie/(g,/QSK00S\c>?2UJTHX-7
&</KE^V>V>Cf5)JHP#HBFe5C\O&T1#_PRY5b9/3<?;XAT5U8d6>NDd_:[FDF7>@,
B9108^CdS2A_4:TA,WE7V_>QaN_b\K_VLbbXSaTbRGF_K50&,F^6cJHFT<M<CR5_
gS@CE\V@fY?K-EZZF_,:>2X36_XZ_Q[#I0+,A)S2BFcfO#1P.PWWdB6J/=,XIWOP
MW]E#b[f2HPe]R]Te,^WUIY_&3(_.B/0KZ.OW;PB(7LU/3)PL,c(V6D;/Ug#C&ZB
-c9]CVWAC7#3.^=5.(YEKga5e-7L@X#d-P(MeDBfJ6d-0a+VXU-Q7[K+C6A]AGJ>
4,3dKIOR:J[]:(6N4;aa4)6?G/HPOL_JV?<UX6N)F[6]#=?[LH&(0QdI2K&>3()]
TYD;/ZKV6CgV@3Q:D=F3][JDcI1\B.<P^>EWS??cM3L)>CWeMcTLgUQVC-8J&0C1
]gfG#FCY7?Gf&/:+A@-#-M\7?b,FKU@EAgMLNID>/N,W;:>g(gXG>?FBNS/(HaU>
P)[:eR-d/[<ZWB2)_TX(@.:<c[?H>S1&AJVRLf@ZE7:YR5=BA?TBWCLT;P]NO?66
&@cA>L_P3;N79&94V]0J]0J+I@-]E9QX6N5D,TVa2EVHg<Qc+]KRgcg2:N1TQ=[Q
NaNR[gCO0P4a.)Q@F\YA@M,PAGdS36]<;UYW;6LE8ZBM3,U)2F[ZNW\WC?OWCSYf
\=Z@@]YbG-+.8:81aTUL19MNaLH+>3/@_Y(LF^<1//c.bHbdfF&Wf2CR<8d,H<2G
=?dOQF7128BcQ/4?g8J3@]:WX#@TK1T[P)?4\T]9<PY4OKccQ85a]CeCNX/Y8ea/
7QUcCF,<;<)_e1c/X;WA.>FO2-a>7@_TA,a&^ffXTc>Y3&dBD1W]S[Re<O9&7TO:
;ffAbDWLY;(5;TYVd6]Y@Za5C<HO(<8G3:)ERPKd8^Gc6P5a@WJEJ0_.DX1DVYI-
bLa2E(+]OD1OS0U(5Z=HI-#1/E]4PF_fUeC3#dQG;P;8<N^[6C:a?\.>N1#Y7cOK
+)3RLV&6R[)(3D#TXI)3ARd(NCT+&)):3g,>-+/H2#fMO:)=2]Z>7VUR#F4/3]DK
d_M<W8J6[/7?O47).9Xb&5JLTa65,?OAPfB7#10f4K2OA58IfCa#;=f>>K:ZF.4[
-4?CNIW4O>X2G#+RMb,V6-Cf;MKV1dOC-?(AK[WH]bW3T,XKCB>0b@gJK7);.dP[
E2HYR6W7=,SEUV+OLC\RQAF<HJROKPC-VPeR89BVI@_2CZ53E(9+[=TV\cXVA<2d
@?UCCdU_PEa7.@82?9JIF4Ra#0>c01J?OHV5\^TI<N8?a^B#fbE\8X4KaU[,e?.&
\[5P<X1#B_4[RI8EISRWB]4(&B7S##_UXbJ5?H55TTTMf0N==ULH,;c?\(+^-=UQ
G2<SN(G^BLPZYE?gf,fNb]07+#T24HWCHH4bC)Qe;-WD6C6f=1?4Y@N\YX^H^J1M
(6[^Z-,5D#QV.[;B>/ZQ&@NXFMD4;H4K374-#P^b#X7f:>FSeVRK(O?b^Cd7CA.G
O,\0]\UI+E(JZ+P.1B?VYO_HMH;5NFM2g:,1K8E?\VP#2GZ_SHJS9WbdP\ULM?=c
S3031FR>[8<dJEQKLUT>Y01MAAMb5c\&)AaKQF5-1A5<X^&&[V&gg2bAEC#1WWXR
Z)LAOM><7F>a0D[dZB1f(5UYgT_+(+XSb?;Fd\M1Je#-2@4V^:=G]-P/#RO92CR=
6^CYLbECGXNJ,>M[S8ZVHKJb+MC,&[ZZNT,I2OJYE5Y,+K7b#HWNW/O3T]FVRcIe
I+S(12a]#LD0>:Vf7^U?)ZG\Q21A7YZ5WeC.<Cb2<#2)U_.EN;Q#(T)Y#T@&-=+F
O/DNV+6I#G1OSZ[VS\HJF]1.W?KdcFKCSHIWTW.:9+,6+#^<Ee<.6U2+.g_@K[R:
DddT)&Q:c]5-5,EGD,A.>1L[C=C?R6F.V18Mb3AAbW-&H)eZJ+.M]G4QgCTLZ252
/cd0XIaLXE00,]22Y-@4eAP6YTQYU5OJYN73F#CHW)YEH],<AYI.>9S1gXR/Q?JJ
J(.]e:b6gHg+)MfB(8Q]b&e[Y#=RG(\V^<dC8L:5.Y#.^/g&.HG+a).-/W8f>dFE
:D4[LaGa+I:ZX5,^(QU;/.U-W4WV0d[+>US\J)OOFZAe;dBO[B.aPOER#b0)?+WV
,dLFA02-8c4&O(c@X)QFbcI5D^5cCISL9A4DMIAS-)GK@FR.^XKYH-GQNG92PW:4
4(5Y&9MT/Qe9Qd?<(U>a;Heb<D,=54ODfYaW^B9?GPAZ3WaKU_@LKYA/f3YN(:b.
BA\X6W2]U0WT.V.)P.BLHYPdbMaDN??)T_E[(QVV8X@4A4>Ma>WO4?7EcF78Qgg/
)eCUZ)9Ta+:U;KAJ4gb;6Kd#gG-MFSV=W@b-9PN,<EQX#cKbg;0a+e;BF<LH[KY&
>OG@_:gdX0aPHR+M[b6IX3dBE\;aE>#KU]5KcEJ4f>Z63cBgORN:5:aQgTLT,ZYH
d#<^T]0[RC8<MSFd:^(N\V\,\U3()?@c(F3^)P6C/V2.d>G(O4I77G_@<==E&5S?
>\c7LMM??I<WPe_dMg29:7\e+&?]MN1:6]TY[\6ad)LWG5,[J,TIf/eB@CULX>Zf
,c/+?<2L1/X_WcO;DUg\NU>V]VEaIN+C>f9_I>8G.Vc9OR9</MdWI6aX3@Y^+Ng,
QW_Uc96Y7\+6Ud//FO(eCP^760&cc<A=#feL)f0LT0.A,0O5Y\Z9?D1&QgLU/@=2
(&Wc(NFCaP>B,=aV2eaSPO9YH?E,1TBE^>>6;T(AG&E<cFHfT=fP&;1gb1N4Ad8J
^^7HNa9D-I;(D&:I,F&>I\,^fVe+PZ\5cH],d(75G[MPJIV;3:0Yf^>7,gKC;VIU
DE#MJ8L1b9015FA&e-YBRGR#765bB0Q/1>R87XDH+O)cCKbH[33CE.\ca8[63)H5
#M&W]KR,5J777G[.b]];Wc03;LN@2de0;]LXcT]EcKD[]5=eAS(@-.Q=MH@RFXVe
\&K#A<_2g5CbHZURHL9@,C?J,7YZF<7GZ:5,/IAd>W<bNfF\=9):Cc:Q>4W:9WZ+
N+8BOU.FSXb&M@61KUT:;(cZ9U]I2(B-bQ5S/2EFFOJW?@N8;CeSMRW.?SF-.>B<
6FJZ4=#6,#>OEdP=Ua[gXR0)baXH+&N);VVVH&DH[8T/\Jc<E.GRVD]#^5C7^XW6
fa<OBcNY,16,EH,=/VCZ4Y[;MHU4@K;Db^fLLT@QR:Z8H(E>M4^B\>+-[RO;c@6@
X-Ddd3M<^bdbNa<N0:eBG@GaP?K9JKbe1+^324cR:NNdA,e992WX]\O6ML?C:MQE
\033NQZP3QXWLRX(VcIg&BEW(gFbb:,0IHS)-&]IZ73YH?_:CX9[Q4^T7b@ZcC-.
YM^.TRIQ9M4JOB0B1[fZbEHL:@QH+-X^#XcW2a/=KF/MZC6>Y7AV4M4PN-P\W=B1
SPZV7d8ZY0gfH^XRJF737\;(@MY7e9Lc#H@#KY.)VSFM8c@]80;\ZO\#N2@2#GBb
[SOG3eQ&ZXAN)/998)W]+4a7GK-K?H(=;XJ6LA.gb^.,(/FA>aYWb6K/bZ/#@<<S
8E/PWO:b5SA:M@?)OBE:\K+V/IC^E<L)TITGD.YfM9RYb?WINeg5T)/6_a+3R4OT
N^@Z+ZO4fES#&\Lg6^O<-1[D4;93Re^^@eg/#aL)WYT43aE>BAM)B#W;)\7+cabf
bb0X:(3[RCg-=M=I2bE-aX2VB_#SQcI7+5<WK0-5,1HfY1f;ag#WRHeZAIVYTg49
AXYY2T/780\DNUdaJad,F#7D]5b[XY9\^20f@8#MgT]0KR8a\5)]?>1KBHabE(R;
2Q4YL]+6\XG_@]LWD.1<0;(INL^UeRY.(MB2C.b;LYTV#A<=JRT\[VD^YOF>28;[
3;A))-SYb#f(?e8e/X6WD1.BU\ZR>gUCQ]>Te(&#2;]\7G\0RN0,(MYH#A2S0,6X
U)5C##@??1P82V^,[ZJXM#GX4D7FRBP#.)IYFJ2UF?VCQQS(O-f9(^]YBIc:MOed
ScOgT^E,2#E2C6@Q;^1d#;N<+dY._=g35Dgg^&FM5X;aSNdGOQM9+RP;?Q[=MFFO
JV=]bGf\FU?6N+8D:KH@M&Mg0\A,I/5W63D1gK;U8X^,-BTKcA7^YdJ.;SS2DZ_L
c?OP+QZP:,dc;cALONT/2?W&64WO\SX>QEH)T-2dK0?U?&W00FNd-DA(.)g@=T?a
ESS>Na07(#4b0-;&Re]A/SZJQG==1GJM+&I+>K:VagD)Za1Q/MS3db3L2(;L/WbW
e7BCRZS/V76U:(aOZ=>XG_4\)GA86QPIg5DZFAZ0\/[c/S8F]eVK^Gc1?44Ce>X1
:I-(=_g62+\6OV5O5=-WP9H=TdGXUM@>08K8C-MS>f#:GWD.g46X#3SA93O\c1)U
6g-;I:Q)fSZ7egKR8bIM6]g:YK6-L\7;IEL3d-?,U1N;eb3&@[_KQLa\->ee]>f.
KNUC-BS_]7.#4J:8OK-M\#9[VS969^Y\_>[_LM))6]8(bD4bfU&M^TJ[TAZceT=F
[Yg[T^M._WF(KYN[@#-=5)BQfOX,-)2PdU69E]RNc1S]RD6U^PWIT2P4#c27;(Re
C/T9<,UWe)CbT2\:@Gg4[d^L)4CP8<S\2/I@2WWZ.U=]&RZCK_5-VbY<f/TT/.VD
=;g<e(:b2_gW]F0\1.CJ]PRcI-_UC-Ab40g+IEOTB=6H#V[T[?fD)e5c/dQ7Z]VX
^>D32<9YcWK56A(B3RQ<<Z-8AK17=14JQ7/H6d3\X6eD9#UO^eI5T;3I\9I0#QA9
20,:L:IZM,WT2a[U=G.U;F,Y\KD:6G@4>&>(]#,WGaX6Z<3QT^7R9c>;EUM3dKaE
@-/#gZ>8Q/58S]/H7D4&ZPUB>OWd9&9Ae0F+<c#A=1^aUSSg]?beRH/)W/[N/J_#
I0PUVg=a5cU6Y9YPb^.XFQf];]XJ_2I+1+>V.@AFeOC8TH,AGXYR>X)ZI6JF3&fJ
@<G&BJVS6Tf\(TN;,AOUD)X#76_O^W7R]ULS9?4abJXaYL@NcP7f\b1F9@>9L(Wb
X#9]Y>DgNG<eZL^U:OX=PHUNJP/<VGB[4+a[(TU0Y=g-EI#/5f5YBN;Y=0MHPA;S
<:RHT4JSLO\0L?=#+@B<UfGVHfJ2NQH]>g<7.-Y5IKJ-LM8:aU[@M>K8#V..Mbe/
ZR@1EJe76#VXRRCN1^WM5>Y(<3QN3HdcbH/,]QT+K\\0J^EA_P6RTSd4(W;H::TL
/>)\1Ac)BD;7>_>C8A8?+>-@#a60XfLA;8S=;,WBPWGX\d2P;7,X6UQ]C,A1b(G6
;[#:FSfTC6.S_>J5SN,5J4Q#a\-S[[0Mg4>C4.I^f5SX/=^cC9:NM01O2#X_V=@S
;MWSbZ=AO4_fA5FgB#8-2V^fR<aFTg?&cU,[?Pd9)1(=U3;BeASTQAW15,ZV[M62
\;Z:Va_,=/.N.ZY6PI^>FaHVO9U2(_g>LcbM6V^(NYHBUA-f9Q@O^#@dJ52<<RMK
AIL&ZRUQe:;Z)f(f:X^ON0b9LOFH52eDHAbX]gXQ7A8-+U):1X=E_@J#SQQ9,JD1
I4@Se)R(S7[02Z;Pg;<]VbPEZOMQ]2S:>:;BISY?Gc4#.>cT9;#EMJcA(3NR,P\8
,1H\26P#?@_L&NY\K<#PeCJ6CJAD6_.g7ZTKfe@5=6N8EPEO^#.]_/FA7YB?)1<>
Jb8bNc2GNKK]N1>gWNUb9<;NPKYc=Y#(-Ha\LWM8d+?#fVDK[We+C3R3JS-8,g]e
/ZHEPGc7:a&TP,-RE_K#@2?.;>/UB.Ae:\,-;7J^9HRE\4H^,_7I76@LK&4BG8FW
&A=H?-b)AFcZ1P7IgN&@ba.8M5R_.0^58)bU]&N&1c.DL/GIH1/3B/^FZX&A[X8:
^f+Cc3T)&M,T@A3-e4+#Q^.5#0D3>F&8@VT3V2ZHD8ZC+IPO>Yb0+0FbK0YBM/WI
2ZJ94@f9c/DI#(VKXYHKRE^>8#aaWN.b1WMGWXAM1d0F9>LIHRK1CS7Y[#IO,d5J
NfVP_H=PNH#\Sd4L;5@Sc^-P@Z2cX,P+ACG2IQFLdQ/?,P<?/I[<,XCfF<F<S<2&
.KT]S\<_>5ZN_)(GRLQ^\dG<8MgF)/4Q9/IdHLfKbY<L^@Q:M.N:b0VCFGO2NNDJ
&.06Y6=6W@D>VW/T&2OOc313b5L^3Y.?8F7M[d]-C00U/cT;^);#D&d+YV@&_OS=
e?&a&^1D,](8aS]@VL[fA8Z[UYKBJ9LeWV6X9I=[KEgWY6L#J+D__0T)IGCVY&>U
Q=8&W1Yaa6,?K3KcV;eI4L@D..MH(12&gEWDIXB]Kg2;.E_5aR_5)S,ZDR<AB1U(
db89>?7PI&=[ZR-PaHcD&^K1#B]T>?TJP?<(UEG=KD.EVg-Q57IE&SSK@[]824C#
P4[^Xc7\N21:]9c8b=E2e];4+fP/ELDMPZ1=-60.TC0S8]dRV\U],-Q:JS;S>b1e
XC/_JE^>VMZ512f\#LNQ;/;SIBgJ<1H5CIf_KI@T.?=&RgJUMHdSU=PEHS@@V\E\
P0B21Rb<OWQVN-P:Qa7AL4c?()B1U3^gN4S@^HEJVH>cHXX?-UR_cG&++(=)K_HC
F\-)5X0EA7GEXcT3D0X].>,JFBaNE_g#dcTB::W8A6:)e>34WP7.C24Z>#+Ia7fF
FQ(8O^/(/G[SE?f\g/@IQ=MU=EM)HL04B@^9?2c+BcQCP2IXC@\H,6OF&^3DbXU(
R](OIgK1>DOK:Kb-MX9ZXD0R.MM.0,g.#Q-P<P;;(XJQD..PA4AP#UBREa()(6>@
9GER;8GeMI+N-\/[#ZT_:a=H&6]P#>8a&M/9R/E:?B0[9C2([dF;0c-_67S+AZ_N
4FT.5T:T<WabCT_84H^G\WeJFTdQAEfb?]HIL(X+<XAdY-KRg86CJ0&,9]RSADHC
QH[DQBNeJ:&FIZVB5EZA53P/DOJ/b,]Z7ZaQ_X_1MTb<>E,&bUBJ74;C182d4Eg_
6>d[\M]7L,FE\WCH0G4WADdJ&X1Y\3/:^0XE9R&X=M,-HRdMgbCe)N?JC>>/R+aN
5V+0J\X?Y/aO14Q8ZJBOJIKWSd@8>=N.b,LAYf3T;6K[/?3W^F54<31S#NXRTN@7
&I3ZXUfV6Y\J+e((GM8NfRSW1O_(H[cbL1J1\(dIB/1^-JLE]B/A8MW[I#Y?9AOH
EC?&cHSM_RR@Q&[Q+L2T72dJ_1UMM_P=\&==T:+E0a>X-\3>30Yf;;F5b6(XO)KS
^HXc09&^T+S25+[(B+86bIGRD6SJ<D0/e([;e(ea:3<H7AUfF3Y.fb1dVF3E^I6_
E2^\)Y#IKL]0X.TOB.Q8;3_RXVC@2Q701gK@39G]8NaQeI:?):ITNXB21.6).Z&W
HM(gO?]72&6-?e9DLa)Ad6?]_<3Y8E.[KLbL](1H.&>U\R;6[40E?]b#1.e1W3T;
#QZ9/T[#Y9]XRf=CA_J#>Qg.eAM7D>7a_M&>IZ>N1^W<L&Y8/?+/gcQZ0CS\<@4g
YF(/?Y#1T/O?[dO/4IXQ&eWXXPLE;Nf(RVI5E=._>S.?X=Ug64f15F+c5H,R(^+8
XOPO3aTaeW05(Nc(GbBXZ=\NO:+8XXK8D4,H3=SSFH7F?STLebg[<Y(-I4?U8af(
QO9FR&G+QFaQD;6Q-aLg\V\ZV<2;RKYZ\b?ge(E)NAEd&EC4^LO+</.Xe0\JPE7R
G3+]UcTM^@.gXO4/gW[@X_0F(aba+?&[-f#LgF?_O55^VU3B]APU(2cbP=LM84d>
XAIJM6fc#_Z;A;P22[2gLN5PX.F8;5(#6J9J4d<L3c>)b@WX//b.(^)?TBeFMKT<
cWDQ^EC-&Hc-@e2KO4P^KX:MfBXIC4?Ie14,[S;:E;b[I>GS>=BNI4D:@f<41)A@
_F62;PMRC;<I#aDQD&fT:J6CX=g]-#@A^L1ULYMDTfBOc:3aA:T?EV_T<b0(AROP
\Jgg<>R;6RT.e](]H#N+#4DF8gI[gJUdB)XA\SaXM7A(SIc4^CQ_gJP]+4Db1?2Z
PZ;@]g:@^I\]47Dg25=I6a0G>TFd,KI&-Y.E&gc?]ec2=US:::JSSd(g&5W#d:&]
IIaC^CP>KAVQX+WeU0W#._1VC[V>2[V7#6Ob8UDE@A&dZ-VVO8Fc)H]_[8bXJ33>
R+LT<0(WNgOIJN^JNDEZUX-^+5CBC>OH<(e2GSQMbWJaVfC0AAA5gGCL0C?Cc3(I
D1@L,f\]Pc.f,67b.U45c&94,@MCNRY;ZA-Z,[.VbR.BR#-.DI-\/H;Yaa^@#<,)
eg88]Hd2W)5(&gO7V.VK0\>&LUV^SD(Z;.Xc/&DRH\b\.3Ub<>[.C-):?^.LGeXY
J<G=1(ON&>?M0<AAEPaf@ad/e#C\6YR>F<M3;1aYRdK5UgZ,H8](]47,WV6Q:d.d
d-MNd[Qc5;Y;I#P+MS(N0:0:VH4]gEHJ^0]e;4cd\@XbB+8->;\YB=bIWP#aAP_d
g<I#1O_I9HMC3@;\4<)>&J=R#Y[HIYe&K,b\>H-L;61:KZ^4;KZ9RFE]EJHK=&BS
+\_]48N5^@&O:-GJ9LFQ391ZUW[[4PDdQ+-M.#>82MX,R2>8:Y5gCPP8&[?M78E6
AH>98F/QCH/=Sc6:JaM9]DXIE2TA/&NJ)>aDEMP[BIa]H5J=^C:e.11L:&g72U,5
A1[\A^RA2<cKcNb/f2>QQ:;ORa@TZI@BG:JJ9K&CEdc=&A-d2J_gNE2KGMLTQ<3M
BcBJdG4?^D:Pa;.dC3QM]ROMgAb5g2([4L.L;3FR8TGFXF2ND.Gd(5^2?<K8Od@K
H<TCMGW>1134TSUASd3+b^N#_C=Bdf<[^4=T2eQEgG7[+]7VP>DJ_&<AX:,W1?9d
/<36-#?J10<NVWVb6JWK7_/]\2GQ@Jg+5(5WeVg9ID3,VT=DA(9Y3E&U;Y9:ed;]
F-f244Q46@)R9X5Zg#:V+dW)E&XaJa:eN_+TSTP.,[+M:H>^[IaX<@H#6(eKfOBF
D[SCLAC#99aR@)<AICWcO94=TQ?b+>>8T,_f_>g^3PJZ)4/?M2eMG\?&+8Z9Q\^&
U1-XObRc[5[fI4=::69F(J->Xa@g&Fc)(ASg][_A1\-f.\G?;8Y?7R]45eL;eG<7
LPC09]0Ec.;43G-2]:WQ[R]J0&Y#_F2/Iegbgb+L@cZCS@4cHGgf)7WS1GCEg,^/
K3S=A@QR.TXcW^4YJ1__#.TaK6[cZ\dbTHK.?e(B.^CGQ&b)T;<Gg?Og[.(V5V)Z
@>_Z#,c0LCE#8;[;;0V54G-cKaGJdL8GFHa_PS6M)GbGOWfI15@OPUHN^XJ8NO<F
^51&866Z=I>46=K,TP@S=3WP\AR;M2Q9a]cWY.0C(F^DPdG2MYeDFJAb3V>3JB=&
DMD)X3<SX08,+-Z,Z6SeMYL]09V522+5N7BPILDU>/eE81PE)YY]901a\I;+?HZ_
W7]HD3AJb\RJVNLa2I:f=73T=40DbRdXdEcYHD-=9/1ZbS&FUMN(9(U?]Z;gF>5;
=&^3gXdO]&.],?&/\5X_8RMOVbg[KO2X[,I#6NeQ,bV;4LfLdFN=X#[?LX#G5Q1+
JU3YUDWPa,+L)ZYGceT1ca-.7[WRZ6KA^03U><gDYY(+2Qbd0D<c\3U4D>=6I\A]
FcHR2VHN2e03_(/^P&=E>f[;#U2H.1&/-_S+P\deL9GTZ9b\;We;_4F-b_c-4;\H
-M#NE@C6K_gV4/:]3C_]+(Obc@HE0G@39QB6R>U2/Fc8cNc_G+IN&X_\7F5V02&Q
U\cJ&_:cgG2Y[e\+;F@dQ8<e>V3X#X>7JcLOMOCUe:3B=GUE;AGZ]4HCXV6WeZ<8
>]96VFQQc^OZ:>)EGT]3OB8-BKV>+=]MHF[+YT,)/5@:X?RFGdL(0]66-=,dDFa#
2BKJ<?#496Z][]dcJ+/3c,N9^86A@+3LM#eaK/B-CdC9YCS:_B,R+bE2S)6=&__>
[C)(.ES2M)MEAGG#&FX9bVO@LQ\dE=@^P<C,eA3M;3(:7;DfQ6[gOGb.I#S=;B47
/>#Gd/K>de9L9]]1Q-E3#]X)dLV#]BGg8gLfL-6#CY_,eFd.\<4ScKP_^;OW//(B
-N6baUWFXN@.g/08:De2:R\_B0ZU?BMKN?[a.0I?e4&OIPXGUbL;^SF.cB)GYZ;e
6e:_+>7?U&ZOBcXF5B(VYT0_6)M4afXH7X-1)EV0PE.cRD4K&987<]&ZL&d<(PY,
=d9>@\EAeHBX:=Z\W]bcL(&DU#g?IbA^#baZ=V^UgNHDfP.-TXGfOOJd_-f3N<[3
dSN<,[Lf9W>#b&e+WU19ef@A>F_F]g>#(gO8b5H+/YC,&.3e2C@&1K):WHWHQ>(L
W9;B5J:TFF7Ea45:L3Q@D\(JLDDTM;HAd2M-cXPedU6809,BLURc:Z-c\a#=4DX#
YL4-V5TT\IRH?aCR&,<.W.#0Z:bR0:ZTfM):\=;RRd:-G<H-DeJVX4g&aA2b@1_E
)&C#2AE-P@bF@&[V6ccTc1G8f(PfE5J6USB;W-EUY^d]87CJ_6Q)3.LYG20E^NIb
HKPd-[SZeG.2+8T@930U5FL]<?D&f@LQRSMLbF14HV>^=HK:QDOYI\Ff?c6P>D_-
d[Z,Df@VG1<7<N7@[S\_8LG.BM?d_]G.8DI6c++cQRM3&cUeNec3&.fGBFCeaXO4
^0??QK<22WS?YP^2WPdEDb[4,[aK1)K#[0M6+5LEXIOXNLe4Tc_CRD/<@eQB+&f+
Ge@NL3GC\V0Jf<?U&@MV\>d-&11OIJSLHD;P_Ga;F/\\]-e&QZ-;.dY?[]d7K1]-
,fFL=f]W(12@+_&9+1^N(SWd0+HO^K(^T41O6KdeG:Tb&Z<;JO.8.FI30_R;O4<,
WB_PDHV\16J-(N-D+aR:g:6:QHSBJ(X&eeCJdgZQI@a20HB>-F7Y1A+TdKb6+T31
NUbAENEc>J:]QYDE:KWeZR=&CH@\GaC19#f#I?89&ae?;^f_eU_aHaV2S/Xd;g6,
5XO[GF&21^0#7b1?=L)T)0_PJ>Y&#65;PB[V+=7+-\2e3T.c44,F[P.4-JI2IN52
:/4WY9T_6##/a3CW1[S]@,eaYL]Z0B[ggEed6KX.4K@X&;PAa[D2#I)C+/Q7dB_e
;@G4;X(41<OI3,R/-LJ->OLdGb9K25[.UDfO:9BJ]ENg_]:.Qa7#.)UPH?_P:F&2
C)V+NZT\f[^<F_^_CV.K:.J@\ea^OK2QbGA&>:2&]]]Q9[_/eY]@TW(Y26GH-EP+
GfRJc+F5DNTW\5a,&6_5K[S8700J293K^0N[<ZR14U7WRQa-8G+d0]/J5O3?[2\K
]AgF4A_,SbcY.SRcfBa?6CX.(?<7KI6&Y[Vgb5-^].T^JK^OER3fG#S&VEb^aOVb
DDW_UOR;NB#8<1c>0WM-KH(gg-LYYKK6N>Cf;\])dS(LJIZN4cMbdH=?JKQLS#23
<N(a]&5ZYQA>P52:1ZQ^<3.eT-IML&M-D1+#g,,gY>_(B)_>;K,Ldcd6F&aLGAH&
(cBA.6aJ(8_.EO-(-0D8d-(J2RG];CZ9QQ9A/=&MV>W]f:K+-9MMT(H#RW?WV4(/
^SI/KV/Z=/7S)dQ+Q9IZ8WMI95cRO>.P:Y7]_P;EIKL:DP_HaHYC?M@L0&#bE&O2
)Z>K3^/d68HPJ+GKU/c9;&+e;,^>D>c\_W0M64_g&7BS?a>eN[NBR],e\d#0)RM4
S#LMM]3Pc-@6KE6\eWKH[bU/aO?CP,Y#(,#Y.F+:HIe:\LLVcR24Y(GAZ2;L\<E(
E\8\7gLe@^9gaP>XG,#V8g/Y6IWLENHN8L8F\Q?P6P^4SA_HVfE.4)[^AE],:8/6
+f/4XZQf3X;c#]8@UWEZQ1QP4;-02LH[KTA_A#S3XP?4&AA2[.eZ^Z3cc8PZW.gT
(>A@PZ\5OC9NBV2W6^<LZZ0fDeLbE4:QgXR&ef.E.Y,^d^.KV4KH7F,[--2LPF@2
2?.6J2OT9EGY([<OBOL,]U3UMbOL7_S9250?CM/9D@Y/#P-;1-6#A1QZ#F40b7&H
C<-L8O0=\Z[0aBM2U;3e.;[S4P/W/[CVQgB[JLc7Dd50Z(VW5cN)UJS1L;:gg+](
W+<)+(WQ@2P-N18aXRUc,/1-=#B>X_D#OVZ9G<TcBWW5D_bB]O;LgCG6VMWKB7=C
U7O3,HdS_<Q;DR+\;&+d:A52Qg)&:SYa?]5GE&1eOMS>199f4KTY959A(GT3S.&2
H5/U?GSEX,:/#Q4BQR#aV<JW;Y[<N.8E)&4CaY;R47W&#KDfc+@C2H3D9.)J_Z\Y
G<c5C^\AC\;f.KL:V[B/QLV+]2KH)SUPR;SW<(f/#L,_0eYT2]e[IL=3D3)Z</#W
Od9Jb0<;/?UBgA:U?R>,)P50(Be.3?>MON97QMV@Sg=:/BP&YAZg=5#=,a;cIX6f
=B_H4g0YKXZ/1V<2g(WDF-EEc_68:(ZDYbYK5#O4R9G(-d)7G+#32:K#+J;_7FZS
PX<=>fa,5@D1UT91N#QI>NW-.MTJI((1YAGH@dHHfG0;3J2Yb#5T:bPFOT]Y4GEf
;6TH0g3b1>Xe+FQJ:76/Vc0M^:&(3#LB[B1^2eG-D7=]cIK=CEfV-?=dZ<5MH>Ab
X)(c+2Sa-.bB,QIbHD\]bQQ[f+O(gT0b=&c^=<cd>_+YR9=9<P4#X=a0>#@14X_I
KM:4>]N6#a?Nb932QY55#\bQ3]Z^LLC.NJD0d1/_9B=4@T4F]25<O.431.:1I,MU
aCI[=]0JI;U_:Xe/YFQ[W3c6F266LL3A34K,_VHg3BBZ0P-V1&]55H5.&O^YM5?L
QGK\Se_[MdK5#_B)8C)]D5,X;e&U(^9_WgWAL/O,Ue6B9AB14FD[L9>PIA>B4\e1
dO8-=@MBa=_C,e#5T8IQY/bIL02+EA=1;KKQRIFbW#+EV_fR.UNW03BG.\<OOT21
?Xd&A&SN(d[^WBID\7:g-ab/C#>=0BZfFWf470d893fVB=OgGFOW?Kc0+]6Y&Fb&
)=\cKQ.:Q0DQ4.SCS0GA-fYZ&ULPF.\-GDcfe=F7#[RTd(Rf^WO_)IG?_-FM9>G-
9b1,@_5SMU\=eW5dZT+Z7)SUO.CXbO(DbQO(DNH]&R\CS][,/YT>86A6/4:\QaKB
H27?:R3_I73A>1E5I)T<bU1/f]AD[bBR\E]#/[DaGAEQ4#.)2LX^GP6gP8b.HYXW
0fOd#?d^QbGddc1=A)]9faXf7N5I#J/)S#NSJc85Y<_c@gc/L=2\7@N+OHf9\8R&
1O[8EM9MPZX91+A@:4J\dSeF>MSIHVZNPJd&4+g:>P/>LN(YY/KH([V?(FZG.cXF
WEHGU+)F5M;8QV]9+AIODJ(L;BC3JL-O^<6H9@6/00_]gcIJEI/)3A13Rd>J\,F3
Ue[Bd:g?<3FeWBC<(C[-c9/6^#<VdK^S1<EGX5XR79d>P_\-CfGd]PJUVP8>()QJ
[8R(_\H+Wfb@&X4P=Ge60OV-dWdS68=SD_>/R)gdcOME6KG4A@@80/ea(#S8<2F0
(6:[+D7fLRbBgO/U#Cd:^g+QRJR03T^cAZ(_0CJ_1ZbBYH5Z.</>a#e/2XV_7[;-
+6:4#&&4#^LL^1K&+N[dPAcA^KM>WfG\AQO>DI5]_[c3.R-RG8<d6Z#L3NN0+7C5
P1V@AX>ZZeR)&75A-4M/W=f&T6#4JQGg7eX)E_-c(af8;A?90(BA7dS1@3J1,-E6
54S:M6;Y2c87YVP3J<\&a)(L?+MCX(3be?:G_<PFR(cTE\SK0MJU5?WI-G(<[2=5
D&VVF+J<@#A@.W353GgeHPK:LZc9(AVPBJ+MLAS[YgJ3LG0d)2]BN2df(Z:T&F-b
9W[DNDOEKg/Y9[_De4#gC0J]I,EX14RK&+P\<F(V8)H#BQ,P3#L4I5YTY@GB]PQ<
V@G07(Eb7&KU57g4&@@4-)]1VCVJ8f4^fU5&#7+R5F;d<gG(^(aR+;3Y4H(;IO.J
fNMeY:M=.U8&4Z,=\8T-0aGB.dAH/63;PKGgDe),ZI08U,g;?RBGFJD<I77/XVK-
#f30TZ6K==A/J=U<XH7eG#[J50&CHP0:[5-ZE@:;+VV1[FK9\?#<6BD<I$
`endprotected

`protected
8Fc/GJXU2?N6f0(-I,<EIPI8e@S;NO9F036EX\J[c-WSY:(AQ@X7))WOIP[c.-BD
MGP\K1<HBKQM@C.3O=#(I0I83$
`endprotected

//vcs_lic_vip_protect
  `protected
-<2?=\V&ICbMFI>/3;DQTa@WD>U=[e9+AMa][Gf7ec2Mc,[FPA=1,(E;\,XWPUP/
JYbMK[)B+]P?d[,&OP&\dQ@L9=WHJMcO9/H4C^P?bN[T=]XLQ+O7ZML^ef;\@T1e
K-JEV.O9MF^O[7c_I-U[A@7;J<YDTH8U:5cdIDLY//4ZeJ<WF(OY5JRLd+<H&,N;
Ge-N_?fO1a\4Ld7KYS49cF]YQ@=A7FDB,Q#IJD/4VGOea,)5TLV3cW=\85E&+N0O
A/^7)WV@-HDgLGFCOTcZ386A6/E>W)T;FJ,=GO+Z?b18VR7G;;:aGBL(]/<46^I?
@BDe0M-C0H5WFU^(A#KcEg;L[IMH4agO0]KEI?:gf0+M9PbI9QAZEBdIY8b?/S16
8FUURURHC<CCSVT<#@S;7JFSCC&CNY=ZUS>YEVfc(P[0-0]a+)H@6(#.]_XWb/KO
=fW6,7QLPAHMd+;IDO,K-MUD^EEM9?CAe4\;c<QXF_NX/eLVC-VC-@-#Uf8bY?&F
989XL6IT<IVD=Z+MNQSB:T0+YM:L0Z0c193#/Ce,:4<?MO1^OM@0G^OAe2R:QIag
A>CD0a:TNRM<(;8UQ++SM]K<;D,5,YBJQ<@JC.I2fX66P7C=1+M?G:&dN?,+(ASM
D[(K[NA3WCf@7faKBK7UO5O458C_5d4Z)RJSbBdK]N8-MHL>)gc(\\L+PLU3V(Q(
?HGb1ISJc+Ze5\7ZDc_Q4,Q.fAa1&M/^DWPR2\L[_)^A:\?CV=X(Bcb2c0\2B-J8
gJgGa1]:UOQT&IAATSKJ?&Q9PFbcF86O]SP:;+IJT]HH<^<P8S02:eZ_QR^d0fc(
G>HE3H67\;YM-QK120VK.fMS1Z+e47-I+9VIBPXQeC\U,DU^#8_LC4Gc;PAOU0NR
gL+3ZL&S9J;gEPL87=]SZ/MH8P2de_Me.RY[@:7#Hb2&gQ06A#>@?R9eAC\+E.VU
3POc?E/JD,fBA7bC:_E,W>+0V.L^@c)E\##XK/@M9YaKK3U2#_@VC678JQB0=YfF
@Q/U#GZ6K19\^O,D@TQZ[@EC#0,Q730B@&4,.V<2>O,;[AKD]=+=fFC[.40B88M=
Q-NgU>4[A:3U8Of0<N)^]8B[0=cO5WHMP@.ac4/5>#=+=ZB4N=+,UKYDMEXPOVaA
,ReM0_KVKD0L/#KD:]I>6g6FHTeY5Mgb(HJ8--LWRU9#Fg^8N)?A:gBF6KQQ0fa-
WD)G1;YcRLDLXP5DdG<MM=DQC5dcL;\A7[_L9GXZ:13IdVeL;3K[3ed9_3Y4,Z?0
Q_;MG7g_27d3E&>9+R<,@E:1KXb7BZFI[eg70eX]KQ_0D)_b^-P6SIf+gVMe(=\1
+JJ8g+cB_2WEMG])G88+_Z0Z.OTa,8Qc?VXQ3];/\a+-AN6EOAJDgPg[L1-geKA1
+P#4^gWT7)CZMX=XP&g1ZDUI3J#K.gW(7d\Wc3e61AfZZ@V1)\f1\,UW3=a-]U__
Y\/K98HZPRWDV_;><Y9DY:>YKV>;4#DX1J\L8+0g?,?3cC4?^X+[?+PDE;BVFb]0
BXW\#M@K0GFUKHFA-<M]Y#UAcNYa6_V+NaE=/43cXZg5CWBCMC?HIS2.A@M5/D46
B>fX6QW#^b^/T^.1^a7\a/>21a+;D3_>&Oa]:B\K(=0^FWbgW#+,AV>K\NQ<2Q1-
O70Z]MPI5M)/TUZG7P_ZN9?IL0J]A6gV/ZS)XI,YfNS-V:XTU.R<Sa;I,<><52PC
#P+;59#;H#W6HD0\2@Y?g#\#Q;:c;5,A<#DFD:7b)I/V@&52c<MA9gBbZU[UCDc&
/[57]R0cFFXUDWWeVV,8TLIOOO?Ma)e]c_V7(P1=BN)P46+-8]8[Z<R+>PPQO-XJ
D8=c5ADFUI<gPMLCc>.)N,E)BJaaAIVCB/a8[3P:)TNQ=d;R.;+fXRMQgYOOWJKI
D1W?c=/MF0d7^VDe4Ngb\@DO35.H3G@V<3#Fb<7,QRXQS9_8Wd+@f;..D4PLV>Tc
T3&6gfe)A_R(.g7&>2017)Wd3_6;=BT00a\12Qg:b@ZdD0=Qf9K:+BD.+6SGg623
CFM0ETJYZ_J6KUO[_OJ3f>T+#C,:UGaae\GG><N</8CA#.W6c4bZ1B_KcMCMD#:C
dC7cD^F8YId:^Td9UK.PQ<+FO5A(?&TQBRVa,@GG/H=(2P.>?#A?=Bdd#/7\]d9@
)H.,JLMe7L&>L6;eZ2#eQ,<^bHU;JU;ZHM[?X[83#N-4S[)YfgD7ZYI6b8C91F]P
]/4dWSN6W4Y=>XDI)g/P?=X/I39]b1RGNS8,g\&412Z6d_BbND\c.ZF8H#6O4:3T
<RGNKME.PXX)-/Q2-+G-GV?@KfKFW++TZ:D#14g<JV560;[?T=<IDNU8>;5Ne>4#
FePJFWXP(M4Reg8d@:WG+JAd,)KJeL,L<,b>\X<fG65;P.cK?D+:F/RJ:8NCNH0b
>09FW\g6+B(<gRI)8Y:D=4(3R,YY5>X0>#Hf-QTEeW=L4)?1=b1]=?R1:,0PWf<+
J.9IW3YbA=c3WO:=E#7;f#2^RB_^62_e9ZJT681dB-IffKI##E7ZQ?#8Ea9,[<U5
RI3BR9KaJZQ9FG/:&]BfPEQ29+^4^;f(H(AEHf6X^H>ZK)C@B(c-Y5XBY/.D])PT
Q2:FM(cYHM&#aPPaDK0G@\S^#;YVJOV4?(,4WeP9K_9O6@Id.HIO=W8aJMKGP:R^
aO(.2RXE#Ua(VOE7d+,/Xbcc(>H[)V4LF^Z&DQMS=[5e=M3Bd+^100(K@SBZ^(?]
[d^([:-G5_LaL)Y<:7gHX4TF=aEW7ebW-OR\1DM3.]V6T6.BT^JO+^VNNG4+0[Z6
@cccIC9gd3cO(K-\]VA(9[UJ9g;:Mf7[3K;L+Ie1RaIH_Dd[_)957EB2E3NX\XF_
B2G?+<\EQdE+(DbWR>C-1OKgFBC<7E>T#,O?cPd=0a/+CZ[XM+NS)J^_^4&DIZAX
IUeg9RPKNfCDH&-V&@L#gR5(5eXL7B8+?<a>(bcaR+9--Z0d/daX,J@:0L[#))(3
&.+4M/3KeLb.YdbZWP[+WLO-2TY3?XGObd5ML2V==QGV;eBDJ0=4HN\S:DOeZ+P^
6;WAAe#Q:=/C-^8gc>&b7><LeA[A?d#1VGM6D[?E4:NcZD,6Be4V74IWYLO:G\[)
D?X((65PN+f9JHZZ=_>.+-V&Q\R3T^G1Hf:fHKP.I8)eI1/G#>fA&Y\3De5\-aWG
a3LL.G_@,MQ@c@SUf-0Xga.]KdaE_QQfL?E]9cMaS^W7,V+EP?C3f<E=.CBfY#S_
.WJ;,)RDag>S-3[a)VGV2@]>N1OBV4YBaJT/-\5X?H,OeV2);b(70G:I[5agLRZg
6CdH0g#JaUO1:,KK+<X9=XW/&7>Se^<7^L,?130N#+H0L0ggA2H-8ZcAN1_a1LBV
1f(.RS\D@0(P9\/7c@ZUc#B.@PMX+UKXP3a>LZEH+GC>Pb#C14&#_F<a)E.\fY\A
]G.a#FTTV@#-2NQ&PXGKaCW/EKJ&Gg)#6B6C9#?_d1ZSB)^D-5PTW3;05gL7a8Z\U$
`endprotected

`protected
^L:]8;UYF>:d1QgaB#b39ad&B;=fN6;BHI@2f8-ZE>]U1;EW+,Y_/)T14&L+L5Eg
B;e=[SVW+FF>a1&.D(_@,3HYOQZK+EKWZ=a]H&?FW<,/&b7.0B\TG?)N:c2,#8>+
<Z05K9=M;_YW8^#J&Q]8OFUE<HJCU^N<;$
`endprotected

//vcs_lic_vip_protect
  `protected
XLbb??&^2FYf(XU+#I+K,93[+d?^A.GKK6I.H9UKB8V<Cf?cWV_Y.(E?&2gAWS7L
0/DffW+CDCKX4\/]\8JXAG)Y/d?Qb\FZX4Fg1NR[\a,[TD<@XTL78@JSO;C6aX_[
CG+]^gCOG.6Q2b2>,#H_feJ+gV,f9=6aB-.KWFIL_<;9H9]8?@N3HaJSN$
`endprotected
                  
`protected
[G0Y]FEGfaZb=dWO)GfI?VIO@cR=9MYY8dbX-=Mf:a_IVfIaZdL3,)1KMUOH57=(
IKH?fEgL\\OLZ^Nf-U^6bABY6&0S</NEFM@RWT^J,M+(I]@aR>.=L11KP$
`endprotected

//vcs_lic_vip_protect
  `protected
DZc#D:1a[<@;NQ-_INfaJVY7).fC2b-LZCZ33cgG@c]KDTFeF+&4-(HAJ0/>))\/
b,#XVL8bf(,QAPB4;@]6&Z:-WXVfD5WeUDI7GdJ=F2(/J;6U+_W70GRAJM?IBPZF
4FR6V@SHO-f+6AQ#,65B\SKdY(_5:UO9)gPPJQJEV7S5/T(;&D04>[L6G2aDCeP_
4^eZNC7MEa08^ZP3CASY<ZVcg/@;:@1>GN4K)S.9OWg9(,eY_HANKC014Q17DL?E
8G#\N^15g.5,fF>f3=O92cX9O&(0\-GASZ,(GX5>bK=N\9+8XfGaJLR(KY>L<(>M
a4=OL6FH@<DQ;Cg.2^Q7aTeZdOLg+/RH=IY/4A6CMR8Oe/dQQ5\DQX^#XAD3BDCd
Oe1E06KXE;<X(5&=2B@2(TK4g<G-_#,HTR?#3.=5(7c>a]-:B;V-e@I,\Q;1a9>\
Z3c=VUCb7U#[RI-[AQJ)J9S7C#T+L,-^FS(P;;Ec906KQ<QMC#.1JGVSJ3<8aUSW
@a<BfH;VD:8FM:T5SgPR_^aNR:&M(ULB7\\cM23LN^;H0S&9.gM3:Fc&b.Z6bIM;
(S#dH_Q9<L;gG=MAb93)8-WUVCb^E^+Vc?I?\H>Da3@.L^W88D^Le5,J[+]F_YZL
VZ()]b@gG,U4dTS7/N+GFYEf^@\9GXN(fW/U9D^VTA2fO<b/;SXAZe/-N@KKN_JM
^<@aeY[.8IdSg>RT8CG,[(I_+O2JfcI_[[1dVQ?EBc,0_eXQBD+[<N)CQQQ6HCeP
:(fVC0dIe@0]64/0=a>Y:\533E:0gPDcRa5L&#I^U0=Ub,cJfQW=)7K(c-d9=N3^
,-=Fe((M,IX4gY:1gdBRB<QT3OH#NBNXSKDK1_S(Z3_Yb-]b/O[T:J(,#M<Df5UC
^A:_S_Q5>8GKfAdfcD8)LQgN6N7a5Z9^g2@bM^M-[He9N/Z)=H)/UV?==NfYZZ^I
/(Z0fcMgBQO6N:feD0e0ZY&8)==J2;&M9J]]aOF5dg7OeDDI2I8>CDHe,])),7XX
5L@0Gg.JA3L]Z.f\DD5Be?+6G:D#]ZO6T#Ob/E-7O[770>dAD@bRbIO)\8R\H@UN
I<OV#S[(eDY3)+6Y7Z9_V?VL:;1Z3SGa&TQS3859?,BOc2cA0P][=Y(]]#eT;Q=E
/O/G3:c3DBR4c3,VN?/gMA7d_3XL,?/A66EW<LNOQ#>18aI]T:V@HT?P&X6GMSbB
Be6[PDYe/GXI5bJ8IC;X&Bf6^UM0\?=cK]7-)\?9R>G+Eb8DQ(3RTfPNBL8BJd3P
Sb=[a;1@T5(];WYb/4=2XB]Ja8\?Ob1_\:-Sd[g]0:a:0]F8B6+Ndb8GNa5D1>(>
G+A[WU+=e3_O0/+,],:U;IZ+^131BO.4C-X37FEQ+J>)2TC(.M=380U_1CYg\1_+
6B7#B^_?g#Ue-LQW?FF\DLI=[66,\^DC+KS2d>558H=G4)>K,QKZYd+@B_WE4R5C
B\-J(Mc14HT^(6=DVWgDVB<8ZH-6QK,f>^C+;FI69_a_WWbXKWKQ4XD=[LH;<<W<
aER734PXe8.I08N6M@JdK[T.@1AeQ#<,/0?c3/)9g@S91G;EZ&GNUd6S+P<2bR03
UVWCH))\O])9_aP0]S>127&a1X#1#2U/cUf56]V=7C[;[6[bKf:X)?A3LIO9RXGd
K7J_0UX?@^gO9-/:O^&Q^C9e3J8JG38Q3cdPRF]#6II0@;F3QKO3QZ2HTGVO\86(
VCQW#bV1TDM;VG.P=Xc?SFDVQWbd6GW+/fSfH2f^c\?1+1Z/VU+0K/=aC=e]KKCM
?&.\EBcB;U;<<ER6g:4g.S#9Dg>^J@].PgW6&QF5gg7Wf8VfM>JcEe33)FT.L@X2
Ydd&+@=BfXgPGT4PJH+9aPHgJ49>;#.138-Q8bR6DDfYE8#+//I[gK:RO43faXfR
]WgHeQ662\^6[,_)58#OFGBaMQAc78/=bfSUM+OK8ae.E:/#XbfV4[L8YP&UP@U=
:GQZNGd=cGR3B+^&7S=a,;^QZ(cS1)5YJ?;S0,K2SY0J9QeO;H1S@OeY]2-H^6^&
@A-,F?/f.DQNJ#1UV1=WE)O0L7[P\QFH,9:ZL3FGec6?G,5GW<+G@+OW9)3#N?PN
46XW7d37=?7BLQ_U_7MDfIEE/O=@2/3.[,,&MEI/cW/0MBH5A^S6Af5X+M.XR,Q,
]C3a3.D)BF;c0#QUH?,T5YVBHRc9Sd9,I.Kd?X1C8FZg]C?<H:C@VE@0697@=Ced
V4L;RQb=C9beQ)90?(35ge0@Wd6E0P15.eGf.-@=5UWfEOHN5+YNB4L(..K=N_P)
?b^52>V^AJE1.K4F12:_)>eU0DP&_:>Yf]_7X@.R^#5N1FGb8Q.,YgS2gIag.[E6
)B^b4NX4.8?VYdg1^W<gNF-L\NT_P>[^]H#954g9J1N.I,7J-eR2;a?XYga&<J6W
LN7VaQf?&F/VgdA[c)^HO27.]]f777,@Ue=40F=P6@C-(L[)21:0J24KHB=R&3Z8
1RT:(1A@XYCcN[J/(EWae1FN1[(;]f:.Kg>bN>NCd,FZ-XF\,[AaYg5\0-?)DB9Q
QR2N^DbAg@-OI14//Tfd6H.E/d)XPTXd^5/3f(-a4Y1B=U6gG-IOH-PAB&-?YHbF
?JX\0+6Fb:ad5M]dGOLGXbK?9#2LZ:=DRc++PE&-D(7M;[QG=Te4[..J9-J2X#VE
SI^]P79G>#cUGJ(eK_DB&aZ<fJ\((D]J8\4G2d4DM6PY5_UK6GX;8VM5,]:=\+X\
JKCT+FJ<>b3Z405H=g@KWBG#&gc8_9)QY-ZX5K[;JNEe,WH1A97[LNPd]W+M<L&0
27&DB64SU<Ke&LaAC.\_VK2g;I4dJgEGH?2\M=6C,<<?6-#Z(ND4?eBeHC:APVd^
H.1,3e?;Q#OFGdNBW-?c,[ZSJO^\FX6T-_))4FM:(bdWC46gYSf6TbW0/XA^>4&@
a,LcM3C]C+AH>+IMF6a/e3d76>T<-/ZVJMQ,O0Xd4U2RJZCUcMBLRNT-H[0BGN2,
@EFg01X?H=N&DbE=SJ(b;<K#F,NE1RO4CNc6#ZN/[PCHZaL4_.>(_(XS9#M)(KY+
5/b#g?:I[,UFC)Q2>bg9L:Bd=H0-T3OI,g[7K0fa]-D3:cPY13g713-gE0O+G6HK
),K#LcUdQ_@ZX+Q<[(^DcB=5)RLD;4@ITPQDV]?dCSJ.Y##8Tab/WH/<ac:=f3a-
I6O03B72eU5AAIC&&dB:Sd-5A?3PB=-g?_1bbfK0P>FP_B\HD3b1gL3K3OXUd:I]
N>\T1G_@a_cZ5g9?L[D?9aC]SU[7-[6-:XC.MEf1(NOc#SgfM27H)c1DE/Y[Q<.1
)aff(_DeDcR]eR:W9[5eC7HcC?S)M5N^@bN3?Y\I,:-Td.C7H\5.+Q?IOQX,,?&S
I/d0Xe[.G;QL7bU:LXC:NXTVHAA)]#B+@M\@?#+fL,F-O3?4Q+/^:GL9MUU(>J9#
Q.9\A<98TX4GCGE^+c7_<KeOZ=L]/L1D>e.H8,;;X&5^ZNDMX1>/+K(Q[aT9_).8
X]JLT^aXTc5^\W@>)e\]RHB5^,#.eBV;6T9,FDEMOH2.]CV.c?DFg\5:Z7<V#2_>
_LN,H]bQ/.<;#1(E3VLYf[5]H#LDYR9A7fF;CW7LE#7HF;FB-0&c.<0:OJ#COY_,
HHNbd[9:2XXa.47B)O,G9eA@90[@4Y;Y+TH-P?Wf(>cDP795d+9JE1gLS&dX:aB?
@0,,X=#DMWA>_=7YIN]7Q\BOJ;D&BO-X<0MV_FL\F162,J6)ZZLU55>B?=7VY1.M
3B>bf)1:\,]_CcA[dTXVJ>\LcGUTS^14G\e+PCIP.-GQ5(MP5RO)3K-WN.e+>Ab?
]b#8>3-_<1)T5F0aH1?Qf(]XA=cAP8RcXC)G].g7:5[ceUW0<8Z<fdc/U5>cd\&+
ecO>a4=MPA9_NcRL5(bCY4-BL41==V?,)D#@\K#&?D#+\>T-+RI,OQ=33VKA(53O
>Y,-#0dQQ+QA#KX-5B3^LR1bA7e(>4=BUG-+.?a]0>.7gJ9Q(S:&96AZV\).?_I<
QMBN#gS<YOE42M44J<+D@\3WbUV_:1/2&f@MfbZLaaP[1^TR/:@d\^]eYL7B4>49
Cd455TXgfIEU0<Z]+V9ZT093/F[e^c8=Y.FLJ954=>J=?[1K/3FHX.2PT4Dd-R^1
dIS,Y_/IUR#=&@aO6f0bJdB/G0dXC@=1=3FHf3=]&;<eX:VeBK)KWJD8-P;_3G\)
&F@PM&)Je2ZE)(MXOR?D=Ag=O239<D;D.M)eJ[@LRF:bB16HN-VZD/Ie]]:cc9HL
\2OLYNL7^#MD8U(SP#3WPUE6#;dUZNBcgSFa]WPP<LPd6G)^71>BM0P7aJ93J7;a
STA_&b_Y:WgWL3C3T)9S^T-\aQAa#;[<@Df2(OeB>1K,DOR57;PUGWE/ad-eYE\c
6b?A]O7.-_C>>B80+PI=1,B=#3SM@L8).6H9O#=4fC5GUD^4gULCGg@NR==SY2T@
Jg?3QXfN/.-TaO5+F.C-Q[#^20_dUA4.@^E<8\U(I)6JJ++>WYI,E>].8D6_TB2.
]N@6&IL+.:_GS#TDa@fD(2TbUI]WH<9Hc]+.2GaGP#K13NIfO.I=GXe?_gD_bEQM
_D6DXYT7(SR#89CN5U@#]3Ya@,1dLR5Z4gd3._^GQ<ZN^3P#4]N3cE_Jg0HP=HN]
/-ESBL0=+X5ag7M+Y37?[EF_0UB<aG;4?V6KMYg&XHVP8PgU5]ed5NfV+E,]6X(5
Z)ZM6XJ#EVX\CNEYYX3+I^_-0e0U6Ac@99Be8-bDE4OE\K.@+Z8;YBdA@,,>FE8J
VR@?Z[+]CJGSVgA3VSDA&(-W/41GcY5cfY.,28R#>Ud@@TJdgIL^U:&[#<\bFdO&
#8)?A_T#\,-ZQ5EVNZbE4K5cZM4<Pe\I;GgX[W@F53RR>#?#c0;OcN@f&ObL/<>H
U9,Qf,?_C6cLF&VWUNMZ=f?VPcR\?I/W2&LP@N_WP:d6=D0G2>@=Z)(W.SgLM)A9
T3L=Z(AJQR(V<@DCbd>>++fB;.V33_##0C]dd+L#HQRDaGTQGg0;Z/>7:QG#G^NC
#7/9.b/_U@OW&=BfAH9=ZP]PfW>a3D\-fELcZ.[8K[ML4D)1GcQ-cO8d^@e16I/_
a4RJg2LaKa0V#1I/F@EV+df7A1NbMfJ>]O+R@;5[5=XF66>HTQD_M4?K+CX_85NV
<^1]?fcHZ3JYHGUB.N&I20MA-N17D6I]>V?4fHLX1D:DZA#O/J_V5Q4G>;+gS@7S
Gb:)O2cdKI9JW_cXK8Lb7BS;HAC.1(CX#EO,D9Y+85SC@+>J@Q#.&S3=\91UV7Y3
JIEbT^_S9](_RX;IX]GD,]I\1_-OZ,VdP9G<b(0B5MeaRK9Ude0ZgBg=(S[:.+<1
GT5DKG7E,Cg_QZ#0Vc<5/^=8,P35@W9(8(XQB5aW+\Z2L+F>??>JT(SC=X_(Y;V.
QU0fb[7&E)E#[_M80\)NB?P(RE2.9)R#e]I]J9#,>:/b<6-UZT/\c-9A]RNgXc@\
ZF)XW0<#P<):DTR:[_8<;^I2aP,,aDQNNe4,V>TbgT2:@D3CY)R91P?JgS:KU<Z&
ZNgC.;ZF8?fF?U@15eHX7NMK[4,dRJ&OGY,KHERMQeM[fSDfgE6_EOe<;,eWB6?S
3]_7B.[L7R4e:#+M=fdH@9VJE]5ER[LPHY^?a6ca\KMd?V#&=F0.MUO[APOC;L4+
+1#:9&fAdf:EW\5OcTR3EWIY^0/B7P?,,O9=/>F4JZ4J8(U5ZS?5;eSBVI06eFD1
+Z_aMX)5290]7QY&22601bPJV6_N=L3R0gCR<LIIgQLCa^7X0)TX+[:geWB9YeB&
,5UbOE.:^SG+(/DL^0ZNV3TZSC0D=g0J+VKCBc8^UI)J@.d.FK\F).BSHLK87OZd
3R:/8SEES^W=9NKM)KGJJ9=MJf^KSS4P\?=BFC:+PJ&2XG,EV\?1(<JZ]:W4:]NZ
JL9e[I+b-1N5C-RVEG]Ub:LZ)eLX-;/KCWd,]3?-I0)Ma=A>F@fdcfXMB)5L.)<I
ScP4gFW#V^J_;ZKOHJb745+\)6Lfa,[,U2I?OZ..b\I67/IWF&6/0IX]+@c0g_KQ
8b1:Fc1(,W&8Hf7#&\XB4g,UbRgYM(acW5\A/8DNC;YC[FKUg^(Ug^N837/7),/?
E,&6YHGBD93Y8;TMW1KZG/1aRcVQb<ZB](d=CgWHVK3#,f=.EfGHJ7H46D.TB@&E
@@3:X)Z:9:0IUB:bLUDQ+FJUF]@9/RUAb+cK^;KJ]&P7;5#N6GgfLOO@F==,(AG/
68C(E+(\bU4V^J6_d]UDV/(V9L>-G9LO[4.G<:YM2Bc(87XA.PcO62AKbPgaUSB7
JK2Pc8OY?=JO##U0d@J:3>N2PO0:f7<aXAIXU.VJP,8]/S>ASG4,AKZg.W?R8PR2
K47T].NAV2F#.1=J:YXK]YKgH;X&QPRI4()&PKaTSWd<.[BH.:B_^>4T4,Fg\Q#B
1^&(AN/_ETUHK#3a._?CH;?<(U0b5QFP2?gX^?AHV3;+VA3UFb<;3+1YF+GIaCOI
G<2[Q=,Pa58cd\S>,)0R(#J=AA)SIA91ZQ]?+,ba99gD8\)gX)9gU;e7=c28H1/X
b#THb@9[(X,d/\47#F([#@-#X8S16F58@1Y6I<,O9,5UD1[F9U,XCH8ZP4Q(ODa^
ZL0d[&1-QLYfK-Je)/[2M1UVT?/Pc,&?e<.7M&/a?bE7gP.PV:d5dg//+&0CGf[.
DXC9<Wec7A_^/.P+^3:MRB3_^I&SG5TcDI&bAV65/OHFcF1fS>SP5+f51aP\_S,W
OW;Ee(S9UE5a/)B5BZ,P4O-D1_61SNQHaB2BB3R&3@A10UXgdDe/JX>@,3(O,&1e
P=36E0@F_+7C:0-+bM,9Fc:UXO5N6[9HBTCJ/Q3##::GGVAR2C/JL;(9T6BB2c,N
F>G)BDW=J=:BA)PC1aFc==<ebL2gA.NHVS8[C9;0#+DUU1YP.NZQ/JMBT:Y,?Yf=
MWg05W4CO;Y35U])5cb.\@I>VI/]<,8<HF&28C[KS++ACL^LEYPZ]4ACfB_?0IMV
cL>8HIYTCWAP?GV.KM,A\G69f^>KbJ9]9_)8N##YOD#80<5T39#LIT_)H/M@ORUQ
eHCU-4&L8(B=WJc?@JW9G=@=2?]B-KVC3\]P>#UFCV^(:VE#15H<IQ9WK9(RI4e-
AU,CH9GXHb:5aM,+.?b?a1;\K:G2<=/PQC0dL4ZCdBe7WUGF(AFe/6[AYW-B3Y.M
Ra\5Ac)KI,H88f64=A^f@BP@(H)U18.=1&Z5+d6H;f:=7&4B3H(G/5,f0gRN4D^T
?1J11ed,L.@FB_^^-a>g97:R=,OE-I:3_d0/2(:;I<KQT8X&A-WH@[:K5LZ=ce_>
bJ1YA7ed6JdFMX?RMOa@FK9[NKbP]J9[CZYCHZK-8-G]Ng5e7A>MWLLO1D9=S?PZ
f7;-Z4g#<T5:(1QX5\Fe_(bCK9..&Kf9><:@@R8cF27O<9RHKV_7MaL_Z/-L;e6C
;7geNa\T+I2T;:X5?]2=1<J=62Q>X3;R0B:G?&IZ6T?^[cfaUBX5+TREdf@KVZO-
8Wg(gGN@g7@B_)N?5@Y#).@&aAM/7[@gJP(O,D/ca@1X^<S1cY(FGe0PG,D>D;B;
NU2^cJg^c<W[7T?E8F_CHQI0_1CI-d:FV0EK72(5E-VTCVRL:I1G.cZNTF?C].39
]\PQ:(;\5Zgc2,K/F]FTJg@d,2,H#(EP5BRZ=d2\6TBg3aaf6&LC1#Yg(3bGT5_5
K(3Ag8HQX/[FPAIaGR5I#HaI#U+ZNY/RTC0KJ03^@c_IC&6AZAA?9_7TI9,c,9SR
(=3@#Pf8ZdaGGFPF@d&DTU>bbAbF+P4TD8TR7ULUaSEK(V2Fa.-SDA]XXgAf=Z1?
0)F@K=H[<M++EgS)/OL)X4fQ@DA^A6RI]&_/+M<,6?QT71LcC<gK[a79=fbR,/61
?81b4,+S>B)WfD,5=_+:f3+>2[Dg2_Z.6,7[FgcXe]Hd9RB?#@EOEc?-HX^):T^\
\#gVg86MSV](Z->dBX;R\ZNXJdW^P(_44JcQa0BE)=2[&[Ec,NK8Z_IGT=?<RgP&
E2DEaN/Y^g.(<QfZ/C^4#dg2<HPT577QX@M/0=+4AJVX2=S\1>.)=P)7UT]UU72C
^0,,.,GCA<P^f[0V(,-6M]:e=_<2+ZF>]M\9fG9J>KK^V=Z<.T&C&Gb(=GNdM_LQ
<XeWUD9@YaEAe7X()]7,=A>;I^]<T;W>3P4:ReZ.[^O7dVB#a38XTfZEH_<T&_J9
N3LK<cVD1O1#ZE[g8e3,CE/?6]VQ.-C^>^N9O2/L\^QXKAG6UDIZD]<SZ+dgbCQc
\=eDg>bcaYWZCM2EL>>9eFXDB[FJMCL4-<1=c#.02964#T>?WR==g&/bG^(YJGC\
E57eA@-5@8L9:MIYUOCFXJI8^GR,QU?dLG>dF,W,L4M:#Ha=b)Q10)g7U+0[O@.7
@:Zf:(_Y0SKB/273^Wa(1DMLHEb+#]agON0FH0;0/A;U:0IHMYYSD9,C<^=)J]7E
MOKb.=QNedB;F[MV#_eZ_1UMEJ^Z9;IX#ON=fJYNAQE-f=?1\fgRP_M;^IQDB0S4
Kd#<0d7X.DKV+X4f)gX;gd2Xb5A]a/_@0c<B7Z\\aa-@3R9#8SBRbVD.Y)=6[d/H
+)7:YL0ZN3BQB5aHYH@Z90.T)c&cCCNba58DT4.VQ0Rd@cANI82Z2JB_UGFYR+^a
YU6,4EJ^90AL[UEY(Lf9ZQb2H)6O4HBb2<Z02b>XPR1@b0Tb,gM6C;dTUSIO4=5A
D=/9C70\Fc@/>d53)N(Z,Ud5VEc>;W<CC<41^8aRKQg<RH4[?0&8@ZB1G6Y9FPJV
/fX\D^<STc,Tc(-Y)N/)0_;][\.L^/C)Id.EaD7\O#1.H\T^/UHS^&0#dIOY>7Vf
F^LWVfE:/ZN26V,5GD4&&4747F]:Y8;)27.+].G94d-><2Z^P2?UNbgJN9bWU;C=
A_DJQ0#L[T,CBDcF&#]_P;bKOM\F=KNd>QX6QQ6)XXEIB-]<AcMbS051-?41_[:;
J&FX8OE_K.YDF(d:FWcB69d(QU[=ZBaA8@Ocf&#_60J@]eO2&6^50>7(bF>(fA<5
57d:F1RN>L&1_I@^#8c&4_4BH>RL;e0LPV(@5a1JT>?]2/-UfNdA<U]8-5;,Pb#Y
N6f+OT<YFIY9Y]S->,(_AANJN_a5ab@?Q30M.bP^=8MBH-1@MFQf;VNDV&fQ]S2]
bQ?T&Ta(5?gX+a_(1P9c?Y;E5d&FT/ceg^W/(EN;MK+.TVPdHJGN?6#UJ\<I-TV<
\P^_,^2.1B/=JF-\S\0.N,T/D,c.38.O2ceBg@N,a;CNE@4F>HH5.=e;\-OU#-N-
D=7.H#6c?d4&6cN9\I]FC;ffJC[X.TdGeJJc=BOc(NOcEJ/]a([:WC@7E.<dbB:g
BF6Ca8+K_;_6TDZ^Wf_+N]^1N=,#/_NcD_)#LF6YFRdQ\5/5,AfS>/Q0KfeJU(.^
DbB:2KS572SJ>W;fF\TDVOd@P^F4WS+#^6cG9.+;4DUC2ZV+@dY43;C8>949fN6B
8B8=.beQ\#&I0;\D5#6cB?OI55L&_S]T?59QEAgQ,gWII3<WD?_QD.XW/)I5>I_6
\\(a\_ZGU4d(GTW,BFP-ZAD_D?Z5TS#fENQX]X115bM:K0JAdf6[5RI]YK#QN;B8
eI:\f&]CI5KU]WMN_]f/GFF/1B^KB;=UbY8V?bQb5LBIcI04W:MZD[2=GB/A&DY?
3>\X^X@]A[gL#TAWC+XQ:Q01a1#\f1&0Z5-VF-U<eHY8cd)a6^9HNVA5^1eHB\P_
JB>=bO:10[f[dR0^I=F]H^87IEd.f-SW)T4#AMDPUWDWa@T_BMa/,^M)AbDeF-FP
^Q(559e>UK38#(&PTHddW2?86FOf.Z7O7@a[R2^C=H89(>L25ZO_HL^(8a][\,O/
=cH;gS]2fTYEUJ7aHKb)&<L71I@^5&O#0]2gb>(_(c3@]=@<a-SH0YTMW/7QfO]#
\W&3;Ef?45^92PPSIB4)f6eBK).\TJZcKE<\1QI<,46>UK1[S?-ZaM4BC768gHGD
W6()3V&_@[S563a8X0U,G<8.F&H>-?JD#SgZc,e>+M)3U.a(;S\WbJ=^E&16G4\.
LB1.-((+W??J11\T9QFYJ-2>.IS=@0[f#P]2cC_?UV&4V<+3:ID:cY#12Z(+8=5,
>.&]O)<TIP?f\M(6bJR0DT-=SS7@9U81OcRe9AZB8M7aDNJA;.b-a,&O56-PFL/]
.6X[<MeH8>Ra/PXGW/Z?E9OR-,/]<XdL]3V<N-eABa00<N,NRJB[Y\_Y\^).cg\M
C>0R_0ed3d2<[(Df3H/fdD^[#6B4DR94UUAg@)eHTEX;T?U6GMb5YLb_?542#)\c
EV:-^Z8PW7aLLH8J0?YB&CXf^--E@[;,LYJ\KW,J.c;4&YC1).O+(2-E06Pba1XM
_d>e08U;HL<3Q,8fO=&2)ITcDCLWIF7#VY=[0K\L(3+;G-8H,(OeGV563:D^P6f0
B;),R&b\R=]<Y#Y6)US15f#=4OVcQQ5X[YQd\P\FH-DPDR4DFGRR4]M\THY[YaQC
g4YeOO@PY.dP-@TQ9RPf\dTI4[^/MENXL,Z+5]UC8YTESG@;(O:6>AQ].Xd5M^J4
).WQ0SB#_B=,+ISE+M./XTL7#@cDGS7I21QMSAQT?I:K+2FfN]C4:(/_6A^:Fb6+
>Me0>a>.RU5QA\9/K<dI;Ag7Ce:Y-3R<^]M=bcJJV[K3_O_5d]9XNGS+4WX97KNI
-3fD(KO/D.XP,1GPRD08?;fV3/NUKPM.&Cg7\&KPRA29G[?R4(PaFbTSMIAU[WDE
a6)b7ERd-QNO?Q/\ZU6KVS.Q4?Y=Ga6/5]:-#@1KA,e)T7,G+,)<7<5d>7<([9)I
#c=2a&cFbFX^5Y,#PP(M[4U+PTU<EZP7YES=Re<=d\-Y_NZ8/b^)4C&ZSQG<a,)e
)&HYZ+/\C:T8Sg-5f,@:88-D3(-O^#R&N,<]-T-dZ-Ua<f&4Lb+#@5S),/)-FT/[
)eEL\NYW2.+7Q@CXA(BI]LWV9]&?fcc+6g)a5(R;^^ZAf<N?MTJ/cQ9G\O/6J2^H
D_+I[I[))E>-L&4b[g[Mc60BW.[=A8[Q7:2YCEGW:RE?[;9L-9gXG6Z[a7TN7:6,
fSR[:5R.(L1M89cZ,WTP.6)HVTFKNBQVT&SAUYGII:-NX(<FXW9c+@-P5_=KE3B6
HG)DCDNLG]=@T-S1#-ZJB8=N^(X+4\41@6OH-5YV1ee]Ra[6DE#c24Z+--bG(c-E
VY1Y+O0eUWEV3S(GD;]YM>0<BAYA779K]6SB6MXB1RP@3.Oag+H-:G&]L1#RQEH@
X,S6UTJdf<5004e20eK3GaeG)]U2.\eQNO:WI><R6LBFFF225.[8d0G1E?c_GVRT
J5IG,Nb=UPMW2BAZ)U;aED1IZ/N,&E0^cF-<c,AX=a:XK5Z4?1=4]((^eX(&/>-M
)H&BC6a]_4]T_G;SR;XD@E6K.3&XQQ8>Cf).d\U\6cD6@L0U6M=(.^efXLY7Ac5F
<Z3A<)M)#g-DM6)1H+QC?KdfH(\=]a](8AQ@e<X4A=:@A#-/<4@,&9[;f9LWcLWD
=C;Ig@R+fJF(<F?De9,BG[P+gAR762ceY^F@8)-6HU7RHQee3\W\H=Z>A&#[Xd-C
bA8>ZR8J2&(90>O/#YN?&)3-IMF@E3.dO?OK4R00>4YUR/<S>ea&I];(3,U+N;dW
V]65^B0B.Z]<N8]#&0.:6#R8W\GS&(cGGR&gL&T<dFUTJOZHKbRaa_-94-g&9FA8
5&>/59>PSE51g&=>M2M-L8R#QR=X\SV3Q6L]c^0;4SL]_DLST_PNK=6\1Q/>.G7<
MFVS;Qd2H78(6^N^UN7@<E>AWbeY6-UZb&3WWa(7N5OGAL)a/W_RFF^H)0W95Nfe
8MT9GH@2.-M=;^]1):=#95KB([>:,Pc90b23RW;\daf_:g=T2OYDfgS/0BUUcSM8
>e:(7LaYc)O_50^dcEI&M6/)[.81WKL&Bb2ZH\>EaM^;@AZ:0SQ#7\W6(;?&[LQ-
4:IOFf</^Z_FHe2H,DR-N2VdTA^.Z3a^(H.aTf/=\Q]D@+A1M/8C7CB\A+ZLeF.O
UI&a^KZ/(8KYS[O-8de^3DW@3d_9aU^Sd=[-7<;=>VR[]f>P51)C8f@VLZN,-.-:
HZXVS+TIR0RXTL8F]@C;WJV,LTS5Z^\.g<))gVA4OJJGI=a.23Iaae]514O?>9+>
[)C@G:YO29K/2QcYbQa#b.0IF.R)(Hc<(5Y3a9:b3L^:D4cC;Y3@#Wd<>X_;];<D
0T02C)T2A,)g>&+9e-1RO(7Q?;b/O[1)>YB&O>HQQJD9UJF8.]0M<00-ReA3&OfO
]KdB//Z[^RA+_TY6:&bf-&M,bM6PDN(>><PCDRD64C>_RECRCATg+H>\b0O0.Ca6
IZBU2)5N7()L-95/&bGF1?EYcNDD0[^\PH&9NGbRebQP)A1O#ZK/03;)b@H_]NPE
Fg@IRcK(Sb29;0HPS@b/?M(8B.2fdE7PTHeUUdW+N/P;QdTTW1\bBW+P8Xc-):;6
\EQ5ELc025.(GW5A[&U\R_WUN&=;LE8?TY?Z0K[YBS,4fQ:)L,/^I<>fRUW+I@e6
a4N[A_>-JLU=D/:W@LOP)^0KD#9#1@TSW^-E@J0K)R2&N9I9VD1)P.CJQeLZJ0ZU
B4>?gaA.eaKg9;)1Y:Z]9\VP:CL>F+fH5JK79Ad_V:>e@G_D>SN;GYDdEXBVDMW[
&SYb_/2Q\5bJT>++RWLED0YK>I?ad)31B-6[?cC+4O-=B[GbE,Nb#^YC0c?U1=RR
BBPLB)<1&RBe8g:<.c#8fK/\gfXcY+7QH>]:[_YeaTM3TS,b\]XVB1-2HS]eR^e>
GB-g=.NZ3f#_5_fE\BfLP;f:-^];<J\>g1R(T<#==H&O<>XH0#BU0ZK<_=6V,_62
Qe]L[CGO@YI]8IP4QSX1:3B0?T^L+C_a6JMS;cKg,T-S3g>3VRYK1NY3Lde<]bg>
&H\e#T#R)KG\\bd0dH-gPD[#EcXC#RW)cT_X&T)#d27[#SUBV41G]&ES7d)=)]Nb
>)K5K:5GdTZ)gQE:(ZfS=0:EgLK5XBbCQfQZ)):C1>/FI9[[@VSTb@_L\0D_L,JU
C9CBAPVZfaX.(EG)WfE]^5U(EUZ(M2E3UHYbOZSQJZV,FNB0V>TJ=4=Zb05#::,K
MMOV9eEa>_8QT(&NO+aO4+?8./>8E,+W)OI6(?g=4)K6<9&#U?Y-&3O@1e.@BRIC
g7?D9J)Y1,b]AJ.#8;HP27<=9_/F.d?91//Q)]VJ2YV-O\??WACaO0&C92FMOXe;
bVQHAa#AB>[3<IZ4P<bZI/H>f5<+8WPNPOL9CWPTTHbZ?++)\@N6=.J&;bK3?C4b
P>AN11=N>)R9Q9X(\ReKg-]U,L(;CbK]4V/dPf<AKb>7&9VG(eD+B8g_TBONZ:(;
+&=FGGX.FS4RD?Z,),GDI&E,OUc9>2c<VL1N-YV8^bZ(9a1N55T;FLRbe-B.c_KO
[Qd)QIB--:9;WX[=810O/S2]9>Q7Z-cbBKId&6a?.#3:e@XLd:_3(G_;]Pe)6FKV
SHV9bM(^<E8N-,>EO-#E/HM#;R^V5a[6.8#X<:JA@0_+C.EF^#dW;IJJRD8H#ZL9
<##W]XG\3a:5Xd5eDb,MA4cI[UN?Y4Gf-=:0)b_dP^aP)=XGM4fG(Cg/47\)7F\]
KOESb1BbGK:THUaeDFI_.f5)/Ubg=FHXTA5J6a&\@P1D^<\9EU@\5(FV/LH--I7Z
B>ge7^eI?DR<cWQY@MX&299N@U1Wca@g)LG<_O@CRXa^.-e)?#TdKNa@6<>J&LPG
WWN<?/B@6W22JM:>@a@=b;B:R8gR:aO/4.d>^Jd\=^gF91C8+/HB,Ad0?W)H6H49
ObZcTX#N461-Ba++Y2<&O#H#]bH)9;O=Qf,0EHYN\V:4:^4ZR:UgH#AIUP?f^6ZZ
RL:B0dQbH.JM>SSR[(We&c#&Z>=GYBAA[cR+:XMN_b6CTO)g3X<&L8^,VB]JH.a@
Vc(aUD/>C]KXH2V=MKTQecW2M@K)FFJ[.^=5&6.7gUPX[_7:;]2KJ1[NfP:E&a@[
W#c7gG,T>)>PfMbAZ,4=);3-FO5@&Z\UUWY[O=/6K(C\=E9Ic>QMg54.D8,cbBOK
[ce+#dX&e+/;+@FZ9>>X6]]KDaE0C6a0@_/H[](XgN#M3>eZR.M&DFV\-.M_IOTZ
(H0NKgL1SU4^LDZb7;QgHQb,>&>.3<gJXUMfDQDS.4/@3cd@;gKI9K^FgBUXD@4T
QF]X].,EC/F8E^&fA4.3ccdX9^0>5@^@d40Ma7Kb<A(&64Qb1:AW=C0d2TTW?M.)
dRH_,]S)\HfDd&Ca.fN(,bL6<C#b?QfL98ePU6BGQ=ZUf#43STdJB(4?_NK@IWM8
[BO?90Z\V+cMMAOBGf1\SJKHHGHJU-GK=F_VS<NCc:eWHDC0afRagfDKV=@DH1H#
a24g]beQ.-4Q<D-TGdc+\PZcgHV:;B,<C9;6N?KRSCY&UAV];-<P8[DT=c[<c4gd
L)Y9F@ZNd(^ASJYfID]<P7X-ZU?@:GAH&,6\7@/d#[,RCc&PM+C9>>,>If)RY^KW
)=S^,]2&#_13M)cE2F/7UT^X(bDVL2#B5L,OUI)(ZI>g@EGJW:TIE1Q5VY(HGU5[
gCH[)U1?J<1.HF>d0&(TSVag<DZ,?76WBW<J=Y(e6V5B3C=G.Ze3V1&Q-)TLUT[K
SS\?:13J/g0f5#P(G;1F2YUC9=Yaa3@cTAgcLU5)K15Z>\S52&I)-gbbXYe&_fBU
ACGbN>:a>9)M#?W#+,U)d8SG?>2QWHec74S;/1^;PEK?f4C4E>aK^SF\(-gRX_+O
cF_LG?C.,X5N4g0/ga5]\R0HKCTU[V6CDO#ACIQ#[d0YTKQV2V)(4A;Q^]RYdggB
Sc^[d0T?TD_)K7X;X#THb^F6.1b/?NCZ2=g3VT22<)C=S4W6;H22J?d9Ce&\M7;)
8e;C-5::2.d,I0>XUF)0W#,8&7ZTC0[]FR80^gB)BD].5)#7((R@DWN]D=eaVa??
>MCM\CZMAH=J8Ld.(WdUf;#L,Ia1NZOMCNMQfB.]#]\@P9Oa49RJB.L:QVB4YeTL
IAZ15@-NX/HV[W#0C__+6PY6(NLH<QM,&]=<=D;^5T@&g)A,[T5-E<4\@Hf=V()5
a]QGffYT9FUR9,KTG&[F3ONd1@e9W#5F;/&9=WI,\/Y=:9E0/WM15^<7B,NfFVZ<
]VE[F4RDa1/;;]FT#Rd7HV]O+I^c)P^\N.6+RBV/38U7,U1-<W8TL/>,[I)9SObL
\6IQgK)fN#,NKXdA)<3D(KZ7[>1^[7g\,F6?L(6+;I.MP4AZ?LP[E&4:2X+WZ#.M
-.O;X\#?XC]U6DWWV[dROIbLf9(A&=WQ7](7F5DBF&LWYgd3F1;?6E)TA-/EK5P@
<(Y?WD8AT/=WM.c:S-I&96)3/V/NLBM?:\N?acM,41U^c^D-d&,7ggQ=@a9)VZ_2
XS-8[K5U_RQ]^dR0HZ&M=C)KB7;1]@B[4Y0BTTgM=PZ(MR0H&W&g4\6U:UVQVJ8?
^NM/GC>)W-GRM0^]KY\aYG/WM@G\84+=WKZPW+DfeC3TOJ<;De)4.-@54D/<E,Fb
2MY,U?^0S(9MHP),Q\e9EF5W.dAfSB6W(C]:N(3GI849YOR5e?&LT+7VUb5^B#_7
NaZ]/+LCR<NAc-AKI6aIbRW@.ROfMdOWYQBF;eUF=gPP2^37R8g<?Xg8g1;>[AJf
bFRf4=3VVcXGFK^\94;@]D/a?C?-HF?B,_e[_EdPbfNUe<f2/f^-g?&8c/-E90f,
4?@<c7=[>#I-A&9f\?LW4I1<cZ1;b&Z&3Hbd9_PCfNeEA.\UA&=gD_>P&3PKH/^V
RgTd3I3-3bE<]?JYR@1LT@HA9-,Y/gP#b(Jcg)Pa->S8O5b(APDQZCP0O-:(W#Rf
f#,V^86O9^D#[].:YRL(6_\2@_^9]=A[^/b;YN_6+)a0/8@@YJ6BUFV[:NSVMe>?
<W84,IcS.0)g4D8[=eM17X+(IFXXVR+4GZSJQU4G.c:RVYW-+N7\?I,GaTU_\QS7
5bN/e?,#?KbMc:LU&G+W^(/R[3eM,VK&J5-SG=13S]RF981F)S;Y/E:.\(1+Ve2Q
N.8GWS,Bb=eQ+2VJQ6+5?.M529GW?9GY.?6,#=.[N82TRObBKHLDD:?7\WXXHNEb
YCM+>6CE&\e3b6aI1@.&YGZ)TBF9d^2d^)RfDCA&JGJ)K#3KW?+3\=1O3);BJ:U)
QS#I6\27F<&(AH]T/?\(?JV^<&bR1-[UB85PIWU[N,JYg>g7ZFC=85I_JZQTMgE5
ZBGTLL#XAG7J]DNW19/9_@Z]4\)a=U[+0McbUaa>Q2(/1PJQ>_Z#a^T?.>,?,LT4
P(YH)06a>PQ>:MSB1bHTDO:@Ve_\<51VS9R_NFUL4OTZ<AM,XSOX&HXNcF?>].^\
^LP>[_Db?d1ZUBZ7L1gQY,WDUZ:USVfc1ecO?8BYONa4e=^ZIAC)4QKB9eB\[O5[
2fS;#7DC,WQ1/D<^dUB8\KS=NdI>+dCg+SSfCGNN-aX-;Zd_IHX5<)\)/c(A3\@:
SLT+g[+B,H7T^MDa-CYf,/1<4K=)Ue1EFdWQ(-H;KEU;R)/U@TQJ1<](d3^aMaE9
M@GffZAD0+GP=8d+c,Z?F6,86b9;5_^D5D_PDR1.Q\H0)_YO=3Z<>dVJA_<&/C(=
WYg15T(R6T50OJJd=:6O7?=_g&Tf0<P@ca:SI)d_M,T7e^9dJW=98Cf1[WAZZgAC
_7MOeS7;S/L#f)1^>F6eS0f8RGXCU42(&BV;G(gBOVR2YOK.]3H?:UWEY3^I;PBS
c6EQ]O(J15G1YC.85dRa7S@=YRY_A.9fF@d9(\/_B_AW+F]3Y(g&9UO5L9GREeXQ
f?IS=EeUeY8@G8@]\PN>N/A9b0N?(cE:>\]LSYWgaUbGPd1ZcOC<1b9?<?Z-4=GH
0VR_590CLWV/3S);P2b6-4eAS3[@<_g.,A7-(8<IVAL/YbP7&F?WgPUN?@eT,S)]
4CSHX>d28W]J,8_0094^Y3W1a\QT1KA(3-6<[W[)<cD[d8YUf?.R)BGW[WR>6TD?
57NdE)1N-gXH]a+D+P?&NQdGZf5J2>-:1D<OUM[XR869;b(EAQTTKaeEDdEZD=RG
<ILK4B,QL0P1>:bO>d^;(M5aE6K7@4ETV4GLaNBf?(&?S#AZdKD]W@YVNN8I^e1g
1dAJWVcDUN+Q14bGW)]]1G,1KW-/gG+EU#2V.5TT<edS5VF@M3E^?a>OP6H:0(C^T$
`endprotected

`protected
3E15+0TIV;.b3A/a8#+VMONSV3LJJF\&#^d0(5dcc:FQ#FW9A3_a,)DaV9<b,gcH
d2<#cc5-ZUIZKH8PZ&CMPE]0^J<UB1)_bZ;;T@_C/WDQA$
`endprotected

//vcs_lic_vip_protect
  `protected
8bRG-FPc+0XZB=NVM8#aN+6W;PTZU@,7d8=K(3<F/RecQ;MJ()1Y0(T0I,dgYef5
X)K=]dJ^UYH3&[f-e-9^b4e@=6#T@d<>+DLeWL61WSCYG7,A4>75a-g[#4&-abIa
STBD/bX3IN(gG2CBI&#8FKHBfe[^>>c10gU)5K&Z#WcAd>d1769Q0]D/Q/7=\6aO
^KeaGM5Lafc@f1beE=1N^FKeHE7b4@^R0E=^-U;I:^dP4)V8-cL,)JL;434Q1N^L
-FMeW3fW;7AGS?-Pb]a8\N#\+#?P=2bU>-e30:P3.V7WCEfWfA21?+D(55KR8DZg
L&/)g73CdPWTL3.S28a4,,YS+]R)ZEe+75P#D0HgC^<g?N2.A#3-XS^b&&9S:=NE
+:\ZWC=>FLIaUTSbJ-QV4a+LE\,/479S,O[]BY>]<22FKf\Q4I[DKGdU8-+7a;/E
\:YGY/Q.8A/&d;?[9B98(f..B1QQQP-4-5Ef<L1Z<W[gZL;=QDU22L2E53@XA##Y
1NTQ4O\PIE3[F?AYd=A8ATPWe&J)_PM+\(J)O?Te+@;O&+MM]b.bRWD./:7?PV[O
,BE41/;/T?-1>98dC8Q?H9CZ\JA)HI;KWI\O&Jb(KHK@,EKQ]fDV^&0[6),:B(+Z
?d1_:JZLY3OeLYR_YB5,/C9dNcVN?e@Z/C209TA-BWfe,BE=,#;@.7\:,/M>YAaL
+?>AJHJOUG@NK6=6C]a5DJK>.9+3G-1f@dC8Y5[(Y<eXK.[S1d>XP:K^7=<;4dO4
^XOXeVP;5CN]9G@3PYaF(ca]>>HMZ&22P(GW2UXLT#6@T[a<.@3E1bJeDOW9fN;-
^(O1I+8\3N9GgHd/TD0Cf0G05ZK.cR^)WZ6HKeC[=]#2PI0.2JHMR:HP1I/-U51?
c:J,GKMD/a28g->3OGA9e,5KMb3L8]]YMdBO+^L@fY6K=9P.RQWQ984b2e=+>)GQ
=:RI4H@MFB-/,4I4R+eO1__\Yd(.e_f,V_D:b;8^9)]e,;?bDS;(ZG@PgX?J[Vg5
QL\R)f\=a;=HJ/R[+<9[M+5Q?1M>De+0[9[8E_?V^,(b?1Lg(>6fF(4#17(?d/ae
D,+:9N+2CF]7;026UJU5O7b5Zbc/CTB>0a9:AFB96KddNBcE?([EZ@c\#)\JL)5<
ZOVKIF@>[G\a>?HS0Z26(g5#9c0X1Xg0_9f/58.Kc1)Pf:5J5LR&EGULdWLDRC[&
[T^&)AY1J:P]e]V((fcD0];OI^)_g7<P#cL[\fIS9,^=e455P8NZ+F_L++VSFN8Z
EgOZ=A2YZ)aI/CggDZT4F::.&UHL-f&GO(ER@0N&;Ib1F+X+8A])]0GOa4L<T\DM
ZgW\?S=A3-P?-2TW7/Q<_IC_X3ZM^R?XdFNaG+PPBJ14\9IeaGA)HS&#Ze8RVK?E
gKPa_&Zf[E/2?5\Q\b1&)Qa&?_\(E>(M5<==LJKRbX;.W][-Hf[K9/@S;_Z.1LAT
G^-AXMWQb/aXXe,@X_VL\&KTAC]?_7B+&Z[K+gB3TFW3N(BO))fXQLe9@\BIA4YR
U[^URQX+Eb]aI()HYK]#H,c=M7dC(gNfI-W<T_((LE(6L1=KcQ;a@A:/+3\PBL/N
9V1J_?)8C[[;Y(OYY@EXS[eTaEP:BF:=[gWURXPG5fDM#b.gSEMJe-Y>G6f_DKgB
:1#13V.E\]@bZ-7KRCDG/T;,I+EZ5FN;E&NHWVMC(.1fCggB9f?CYC&R=Y&aQZ+G
JdI>3_+1]<R5/@-/a4RWR&C/c+b^V-E]O3FC&?W]]]M3c[8B1M#U5]]@_LSP&EL.
5bYXJ#?@f.:[\G9F?\Q0JXT5LIWgRgU#[d)D;Vbg/#(Ze?(LR<TM+]bY->\=YH#V
OZZLd&?SB)QdM^/d;NP@6+KFQBW:7=@\1]]gA_)YOXZGO)TSfHI;VB?ZaS6be:U=
?eHMQZ^+;9G::./WLWS=1L@eG-^OPQQZcH9VY4;ND49,YfW75NBK)T0#EaZ0aSRB
/\?)<F[f/-P6O@Z_LO2HYW=)H9:HT[G3\XcSTIdWRA/5Y)bL=,]UX.NW)M5:c7TB
S5J?ASL1,-?].3VES,.Ie?ba#6/b)>c+e).W^DV@JFBc5B7&IH_^CB-P#&D2bASC
H8N/,KP;Wa<Zf_1BbOMXad<VB-D8Z3aDcV8ZXdDWKJUPJLQA81&b2SW7<A6Ubf8e
Mgb>R;cDPe=<ECUYO&&IQ<]Rb+7?Tb[6BK4a:VRL(.]WXB7AMH[)X)AeP0__bGHZ
>/(ZQ.U?O1BH&[985(^J@G\HGQ-fU@]4<ReJW6,;/f<D2B.3a3-XFe\YA\:_?L_=
&McLdL563aO\T4@b;5ZF:X9gU0\IKa94>5HY^faTUSf6L_>e_NZ+G[-Z&=BK-KSC
Q.&^UK>CDA@4O6B).>Bc/5\-3P#AUdP_@R,gUW=c,@69_g^aCKSZ5?452BT;[LGB
C5(30Z?&O.^7SOcLJENUU69G^&;7?NL2f]0,<37TXLRI^c2<Y;OI#^V_XY[<@J&Y
KG?He1K:4f[QLCVD?9W:Z+,;/;7XQA#Y;QFC>g>EMT3G&(R?9JKe5^(4#G(\-2TV
DXTFNcY]R/0Z?eDXWX+@cR/0e]+O/+:VLFQX5aR_OIAa&)ZX]MBT,Of+T/E;;A(M
WJ_-W_-V]NDBX5c^+Wa.)(-D9E@4dgGeQH&)E72[g:bLHMS-F+3\A?4.a5<cWK])
NJ^_-bWcI#(:[ZM[6_CD_PJ)(6P0#N3QC9ID7AB;1-W3VX5aSQ7e,,N&[EBJY#A/
8?+aJ]6G/C\E@)@_T=gECBbY_S@(\11-bYbL-HMJKP1+bR:-3@CPg)>M=Fa)IXBB
RN#0eI1UFZ_[c#1S@=RVa=c1GS19Ye[J77bI-e[98T6:E1f-.7SLGQ64G<g=[[;V
&)C([S4BER,GO<=dX6LOWWPOFA#J,56R,XQUX<I;R3VAQS9Hd1I1I5TJ#9]@>Bd2
OJKI+eN0)dfPe,Z^Z&5)+5I.3(.VNKEA):NG3(56QZX1aUB-L#)8]aS&G(>:VSBT
Tc/&&4=.Bc-@3IbZ9<W:b20,.)DB)eH)KE_>JHfFP+R;<9PMG_ND)@ED=CDH2N67
4EcbQGFDY]83?[]1dX-2&7UAaX1-0-2>]/d=cO;+>E<T7Hf_b24^R=;26BPF5g(.
;2B7Pc7GR99\4Z9g19N-DDZ/e?^,Ha+BgVBFc<,L.2JB;QRae3DSg)QJ(UM@dg)d
2V,&?3P@c?/T&W?gTf3]JJ0HN-W5MFeN:YH4QWbG7L:LC#_c\7^-b;^5JO9dHd5R
XcXK7UFXT<YKe_LA.,\\C_W=(UT)RCVcf6D8R&S]B198-CfPB\EeYV^4MDS^TY2=
JL8b4[6e\3T;AI+ULV&fM-b:aVB-6MK?.N,^7gKc]:W3KV5c(Mb\(9KWGTN-=8OB
A:UR3;,272NH(__EdY+6.4F]\#G+AZ)XQM@FGQWDIXT&84+8>HcA=Cb<X0cI1c,#
d:81[cN-cZ2N85bOfSADW6e0Z,NHLb@4T]CMJF)33b_d+-^\=fG4c]T_0M+A0R:A
2?SSAd13cMR2bMHGWM3Lb]KHL-_@+cIPPKeM.E]&B8=))PD#TA,<:)cQB?\CV(gJ
:BJ,S#]0.,d#Z@N>Q1J7L5e-8#-DgO0McEe.YHRDEaM_PL[6AMNPPW7<d>^BMUd.
_Y>g(g.c(E\NIYTZ_-fN0</;GR,MMPG-:eJOgJVR;WQ=7:@2\A#Q.XEKTNQ<FR?V
1Df0GL)B]N/EQe#;Z#Y6=)57fWOE5UV&OI@WbbHZbR+.XZ@#OMU;45C@Gg1J.=1J
]ZbVF8^LO(#V/DgSb#\)VULN(,Y,Y780.>@aUFT<RSV4b-Rg_e30Y55;P2DM3d<a
@-K[0_VaFDSaV<_81Z>JWD@Y3,Z?+f7/GZH:7LRZI20e4@Y>&Sg9M:]JXKSMgKe<
NC&0HV@1Q7LC&JUW.G=a3[Y2&MT>aS,3]Dg<eSK#8I<5NLMeF;(9QTB9P).PCJfV
)(RN#5EEM?\2KcfL@A]<dQBVJK)gO=+/P7GV9^8;gYL2^@D2a:Y]Bc/\/fBN28gN
3[T22677..0If6fG>ZD1/Q[:bEH4O(2HI\[V2RKc>6:1INE[4GI_X/<@S6cUb;)+
1P+0LJ&[0a^aUH,?e93SK7dJ5.NQGU(L:I[a/0?d#HDLUgUe>(A-QY):fV5G#U<g
5cfQ^G0+NR_QG1EK:2</Z]0Y>fc28J.?g1?#HED_7D5QV-6;TZ^G^d7BV8=?)EDc
:9/:_;_)_IVY&;G92aQ[g-d9bOg-1<SFMa^a4G=L1:_OH8[da\\Q/MCEX1;==Dd1
2AM\5(3MVGK.][QPSTX<G:GAeS(bZ]2#G9>Q0V:NCIVS(>MNJbI_F:O0:-_X)bIX
fU9M2[NJ]#-aRFMF9:>_Y>H,J@8YaTcU4gA3LO&=eMV[Cg>G&/D(=:R6EJWUNF_I
IJK?gP?KFe.)Q8=FKB,3O0H8Z0?BQF2T&D,?8Y-ZW9=fF:5Q>#,]ZeHTEJ=-39#[
T6SCPc7c7b/9b-&5cIXcD0<W)DCg4/c?R(.H4c_:<;7c:;aGc>Jg=_9cT8L(R>:I
Te6<B2a-W4cb/=E)9+9FEJ@^8);/]142Z4?(J.36_(L7P)C-XUT7GD.eC9X:ab?e
5JZE5:M78^;88L5>Z..NEF0(G967aa(>G:5&;E&A&D0\IQ(WOR&+fEKHT,/D)&);
\)[KD\Y9.OCA#-DO2cSJ9T=g[MFQ]=+SO2+?AY.\T\Md4;#\Q[2A=,Z5@CfQC0-R
J3YOH<DK1)E(KGgU42D0]\#E7#BdNR60,?/=TL8IAICQF6Ba,;<aJA0X3CM#BJD2
>0O(bNae#7BPX^?6XG=eV49;R1d;[fLKC2@XOG/QB;(<EMVW/6eS:a(NUcfJc7e.
-PV^CFTA)&]3^]dV^KLP7P8&L1#U-7-LZ.9,Ee9O.\0D9.G-?Q87)-Ae.COR<T(V
P3#&FS73#dEJCfN^S@V;aB)FT867,DPS[]-g#Wg\2&SBCXT?C0@Ob[S&[.+ZL8V?
9_M@AN6[7D(_N7JCY5XCM4cP]Q6]B<Sd8-6L&[a@.LBD[P7L4RNfEYF720A1\XEW
3]GMH4g456c+g?17\6T;DI&Z,f)cY4OOHLaR3:BaY<P1F#/][<[I]^1YRcV-2=;?
<UY^3>S>>L(#(P,c6<bCOJ\,H0YQeP8X7KMVS7EPOBA:4f>W:c1VP.M@Ne)S1<Ub
TO<C7E>@Hd[AK,ZcDB<PEH>Y9&\8;\c1&b8#3@[fb#a/4D=#00Jab]X#cBaP)g:?
NKJ9TV#7M5_/0SW3aC9#:c)]D&,K4\UWYKIBK-e#F,A6F]=A_3R4-#gT7J[Y@?a_
9YUA4:^8g[D-6Se[d-LG:#6I_^bC6PW_c@^E1V/f=8Z[5+0fV_<J=#4T&/1OFV::
7T52]T)2B9/c<MdXD9TfW;-N^&I&bH>RY_=>[_CMZ.)f19GZ972g_<)2TU.8S#V7
6XN:FYcJLe#@TaPQQ6]D+(SGa1bKC?=(e4+d?GM@JPfEY3+H5),WESA11,W#a<UB
5P>YIcBO]UU?L]DJ>:EGdGAT]^J787bS:N7T[2:..g3EMHeWH<YH:R/Mg@^6Rc]V
<bCB+-10N,[UQbU+Q[QUK^4IXPBS9>GQ-JSLO<.:+Z]g5@W<K\aH+LL47WYYNOC,
=d,S\FDY]>_>O-9MKD&Cf<@098^CZX5>GL?N=<CVI9RS9,X<.M>1083V/7Ja-F7I
76EAD3JENa7MP)XOUPDG6\5O;>ZP0P5@BPOJ,B7>]4VW6]I6OFMOCM&1EWGC[H+(
-fGCHO?OUV\fH\-I=;a_;NFaA@^2]eGaX72/1Z=5]I)LBeXZ]^E?Ee+?4g>H>9I)
7:?W;Ufcb,Q>@be)&TQ0<:4\V##f@9_]Pd&cKcbJH7EBc8+CRTRH,J,?a:TE#Fa.
MS0fcYYCF-)Db0+9&gVXVaQc_2.ZG2YPVZR>b2U+7d&OHPeaZ295.U(R2BS,))cC
]/05[:PH_<U&RaT-,Gd,.U/VF+&QG<HQ?X8]FKe9LAI)c54Z(1NA).&8#BG/.-P1
U0I]1,_?5)]M.?6C4,^2dN_M;#gK8]N[dgA3aacV(e>.,9K,PS4CaBF_SM5Z00#.
(B#+RT[D608]^7F0=c9.<DAA=T5OJ?RbN@VVP6,FUb3@];QHZGTd2/#1K8V+N(d#
^6,P2BgQWdYCd)>S5U=J0TLR[AQe(NH3L6MVFDQT]=3KJ:Z&G7bWe2A_O,K<MYcW
7&]5QGg>E-7C0\/[?M.?9#/AH))AHa_b(7]P8J#.QPVQ=?;K+)/Y^X@^cV3G.-6U
F-^TR0NDU)J@bFTO9JNX-_DV7eNCcH3&P?eX,T6bbTICCH(eUM/MT[.F1_c/@H8V
;F\/90be>bR5&Z8L9<eM.\HDP]RGTMEd[1S1cFU?QafC0J^)T4^P+NTV]H[J7e/e
T)\3cHQUJbZg55Fb)IM&3BD&1N^HF7e+^0<7QH[H8\Rb912N#6@>2>#RZG.;QKLF
D0?SW8FVU+\Ug@3>ZX>=DE9H18]-[,F8U9N&0)eLXD-bQ9SFL1;(3ZJO&dd:ZQfV
[]&[ea1T.E<D-PbFB:OU3:..]+&@@7:+F;1@0fN0e_1?]/ZFg>-T\8UR_a<A]2(3
)\7[[0Y80U5F([#6/:@LFL\Nc:<3)dH#8+6/YXa3EaPW2S69Jb6_O_.7E:V<8>+U
2d@2RB+;?7G75bEK56VMe@\-C[9d#54dZ&^60F=T4(Y(V^LS(E/F?A.2.1^C==N8
:+Za.=EI(KLH+5TK5/JUEAL=\3ZCXP\9,[aT8SU;3dHfJYBb:ScNgB8\1A,^bZdV
^FaVAGA\dgd)Q@WB^[I8U]Z\>2/5Z+AF+J#A#,:3Y,Ma3TBFH?4N]Q.=b2:Z[V?C
57A(<>:V_MfP3[5#^XM-/:ZEMRH_CMc[TYbdC4e?gG>[^(?e@;OVFRaKMWgNJ,TD
2,?(Y/UE.JX-@4=1?A1PRI7H-/6(X<-aJ#MI=8Zb?;f#,c7D0\^8^J=:JCdDD_)@
D+_]eCKO>Z9FF=<aPD7fUUX?8I\gFC-Ne2cR4O6ARfVcf7RVS)&ZF[A=g]BDY6I7
+_[T(QcANNf/NaTWe9Y&fd/3>.0^7@BLGWY<4I6H<^<3&@DYGU>)CD\4R#V8b^1/
TEX@O5GbJ28+Ib)//X.e7#H(0)8cO=)QT+4gc.@X]FZ#QP?Gb2S+.PS#41YL>828
6&eAG0Y.4>KF]S5I9=dW-QE)^:]0U?YE/bd[#Q4:S)G.+Ub?]>4N)V)CT=4G.UK9
gN7]/CU@?>?U)OF-C<:A?YW_L9T]aE6c8A6e(B]3EIIFREVeQaD75A\E,EIDA(^I
Xa)>5.fJVRfQI6,bU?dOT\B0-/.a)++d\XC+9E?Z)gHD7<ZJQ6;Ne@<D1U65>GAa
f(HN;IYT7-IPX8)-AYO(b-F(K#._T.[P8?>M(_JbZA^==RQ:MDGEV7:,Q-C/?_M/
E:3=]3587_G2K[,K^cN,-42FfO_ZAd;J<[?F[SVYS93?YR@d21I(2a#4#6DUY4_^
_R?#+)NHUf\Z24\Bege#O3J5,>YE8AKa3:[VaRH[V4(a\2S4LAY;\fgTdURE>HJ9
L:NG9T;?9;&^5DN(.1(NYX)NQW&f\50#^7VMcAW[MH1g^/JK=Me?MNUeS?JEX+^G
[J)4PM8KK4a(F8\&f)eD1V;5eG,)CdbR6Xa5P[7L.8_:94c5QPNUAUEO&32K&KBV
45aF4\KJ/T.Q+T]BL)^KI<#UaC?_O;Fg+UZV@1G\I=3eHJB;77^K^EgGMY=F[5d[
eD7X9,OV?@5VK#PB9I_P70\YG(8^+Y]<G@4WE[88/E:3PYX);BPM2MN3b=OXPMcb
](GcS,7Z4db#A=c9/1AMB^6Y\9_B<Xb.QP6dQRTK=aa8)IKYQ1VMNbD3#W\PY,_U
<dYOC4;M@;&[2\1[fB_((5GfLBI_^9#9Y>H@G<FPGfWK-OU3.d@^9EFXFWB9DVL#
ba08U9KCMX.]g><[N,J#.>;bFa1-cE)G6&]UB-./f=gY(&OfQ_.I.,d73[6fPVT;
HC[,L^4O_8eEYP_@6f89]1?fGJ4:<41)K4fK093;cb_41K23.]WWe;be&VcM/N9A
ffAN&7W-0F1)#d4LO3/S2C]CFB.;29[:6OWI9+7P0(H/V<YZDN@E-ef]2VV[:(?L
EJIS.g13Af>,J+A3&F[(LG.A^>,A6S#AIUOQ79P?X6cb8YZL&+BH4>7LT(0\1>0<
Of0;O5S^f[5E28d-.b;DUfG@U:LC0^IKC#Q6d9K:CgIE[aKX]4->ReV)#I)]^9eK
JP-CX)_@[,If6+8Qc1<db-NYVX?)2g,C,S4-QB?H.V>YKDSN#eH][@C=HJXFG1^K
FYOI7fB1#<)EKa0HBL59->Q@QOW5;I-?@g/BJXXd/3C34Md8W9_LL&&UW2^<V(24
L?cUc5:9DPZLB,\\2d[V:,[de)K9O9F^N;A3,1SK.[S]ZEc;_XJc&W;;#PcQ#5MJ
_UM;egbe5aWK>GZ<P<aEK)1>WEE@5<dI9-Y];H&5SLL)a:U33V.A;K&L:\W5C+Cf
KT5L/\N3Q8\(b:)U3/SVEP^?2gT>Z85c2XX3NAR<<6W52eN_<O(;>WbP.>->-49Z
[?\)c?7&[]J/(b4_@JT3,/Y2cb=0OYL&cWCK;E)N]NJ>]:f16KS=EPC9@R8P(TG/
83AA(5g=bg>NQ;YXVAVYOV@4dB<]0RIY(,:1:GA)YUF:GV\-PaE#/M:RFea8ffab
7J,^XSZ\#FG_]Z)OI]MAf#G?IFEAT12#.+6S)A(?Mg8^MU70ZJgRb11&]\RRZ.c+
&bMOZ(cf;AYgeQUQ^fY7gF<=J<W^^6\F4U:fYXgT\D;fX,F)9e?gY)E<FA=+2#O-
TZNJY-dDOTX?I)^+5?^P:HU?X&#bDV:L1KSY)PK3QIC_@5S:ba36R[MBEKfP3NZS
d@YG@R7;K?A,G1CSW#=8]#9\AC[)&Z<[R9c462^F/LLc/811c&,]EE)FcLDBNd9Z
>^^(.7Obc1A)]8ZB6G1@Id2G[&4OR\\UK9.cC6R(FO;Dd])E.MQH:UFW4<P9c5Fd
-ISb/9(P9J]Y89<.f(Y;^P2Y33@7Yc60-6<J^XRa,6S1FKYUK+H11Z7CBA\1gC1K
Pdg6Cg_Y6Sg4(fD3Kf44T;:5@,O58Ba\GbQ8T\LLaU:U<2a^ZR:5VWY?\a9de<aV
W&b0aLQK]+<I>09-Z_AO41:,F&9._DFD3(BKJ/A<HSP1cPF]F(b[Q\,&/EV?M1C^
Y>>Hc^:f=B]V?2AT@(bNeV;.G6X?4::RWH19+YAa<?V1)3.YQaF>dG7>T=MbHVZ8
437<gKW&/P7#4@NA>PH67g;)-HUDVK9fS5;(._f?#[WZR/(=/6RQN<?<I_[#Y,7_
S(a0\A9fdME3<Z\:,4G2g>.C<V1_1T#+^5(Bgb>628;C;9JXaPX1-3(F\b.0BQ:f
R<4FR1PEMETW;K(:Z/FLJDV#AE1F6b&KcJTW[F[V7fM==b2IP:A(gM_gTAY9XOV2
AND[Vf>=@=8W-/HNcc67,9,8R:9aRIM&R1,+QTS4=YAT2S&TA:LfD^)8>=VK@XeA
a.I7]G>]PT#KXPMdgLAG4fC@EHFBT@]AK=./7&HJ-J^^KK8;Y&2W+=N,O)UB6N_B
/,HD:Ea@3#<32c7>X-QdO8gHNTO[E\.2cF>VM?N-)S6Y(GF<EGGC#6HFP4J1#469
d23(AW/F,N->9b>_3c^B\+gg,g6@YPf,O(@R+(d(->]e.R\+K\/dA7ES>@,BMb3_
gb]U#193X7+W/bMJZU>H\A^,N&HFX((_)<NPa--f13Eb5=45b.HD-.O/T96K2)SB
(8IC7QM^.08-aW+dbfbgQ<5\Z.ceQGb#+Ba)UcGD^df4<_N/2:0Z\VZ-N[E;/bMa
],LVf(#H]L;8>?4d09)C\2X0\[6U50/=F21Ja;L1UDEc5J83ZPN1=/AYOD1>+#)H
C<gQX5>gEBV,<f/0Y2Ua+A^[B?J27Z<AKF\9G?^/ag/>#T\N5SeDSbE<<I2YIR6B
>R;T\ce9&M=8#V^eMgB5VJ8<(F&N9a7W3T<NEEY&8IW,1YTW499J,M/b.-2.U4FH
:8:K,aD2U;A93/^,Gf7ad^+I@#U#1V29a,2-(#8Z,W38fT@D#V..5g+Jb.a(VMG>
9B>TcgMLG32D3;_IZJA.,OH4/_b[ZM-Bb&DISdAY2,+d]V9Se/;V#,?W.fB^LG&+
[+_3YPANZMW=:U[<RT9/dV44\VBEU_Q<bDJEY\dd&GY1>OMAJ+d\_Qe=PT01ML:L
\OU6P_8cW(X[R<;^PJH/V<QQ3bfC>Ye.?QOCGbTFY;gf<&FRa9)aU/W9Xa<BV&#b
_<\RWI^<cF9P=JPQ:Oecc#D-9-97;cBKFO91=S@dZ+f5MEWMV:U^_\:N_b4]Q>:[
H+C?,1dcMTeGbR95Z549A(<N-CE0Y<,]V>00Y.78gW)V4K-2@WU.8E:8)(d(WJB-
3aL)=VME+@(O@1^N;@.JTC&JY?+g+EA]aR4.@f_7OVJNNVI7?\P<.WNW.?K4)Fg5
1FJaeHK8Y3P@?aca_4EGY^Y_HL&,B0VSZbF5@YP3-VZMMb,ceb7J7:4.:OdUVdFE
]2?U=G,O?-e5eK7>;[^1H4NKZa3&4\9+Z_:,)^_O/b9(3)BHL9Fd5KTG-.Q,b?VK
WOVRfJJF4d@8G)>;1WCKbYD23S_a2GE=MCU2Z^f&0Le3d<D1O?P#2e33Q.9YJ/E2
YT-.?M;#OU/ZJ?0YTJ?K9D/AJ(2O(R+)K=R:1e>P4&&IZ7@e;)D)JX=C@E>2OJ#D
(cH3R6TN<L+Z(9,9SA\^Y#TE7):Kbc3:8EJ<fF_6JW/<_T;b#ZcdHVbK?_3^HN.6
5F?6Tdgc:^H/TV2-ARRWJW4H68DT11ZbU9.DGG[:W;#Sg1=SX(>:Y7Ve/P=9VN[M
^\L6L+86<:A.E8c5[P:cW=HC^?,Bf/,GLYg8[._[bU\,f#^-1f/>fJY9,,c8C&K6
W.e3UL(SBA4N_4W^K_Be)78V&(@4;B(8V<,TdVJ?Oa.O[J\J>N0BK_@/bb:-(GCf
08&_&GB<+)KQc6N+_><EgFK03HQ;ZQ=FS,Wg88YMRY>]JDKf2JYALA9ZaB=D\bZK
WBceRXfV(+O#cWZL-SEIG8U0d_7^_\5++X\f?LM.g,A6LLOSCH-]=-bIJ.@_;\:2
IBX:)DQ8&ZKJ7g^3e8;?b-BVQBa[]?TdY&-fAGX+VK\W[:de<2ZY2I/eXg./I28^
;AL\AV7=L;K.6LLZb)AK=[Q<e9(Q_gBZ4@H0gF8R..+\e>I2?B?>_]:DQO3cC(QH
IO8g4gY)VHE5#T01::(Ja)d]5MC5:MAZNZA4-+\)M?M5H]6E?2F\0+GL;FM&LPL\
J+Q.P]K?#AI<-\Y>?O5)QF=<GF1bS(g5R-3[8F<RMZfGI<?,<.U-;NcMW06[3ZOD
=Ng3630+d81&4@<;V[SX;+>X?Jf5HMXadL?Y/9T>Xb=:[[K+_QeS79be:2QS(55-
a<=5[:/N&(O^Q^\+/N5PWXQHV,OC93A<eAX]PF[S1\9_DgTKL9a=ZV^0/&a=WG?W
<4Og4=65,S6?<.Fa8ES/K_+(8:cE9)KS3@NNKLOgQWDC\G:+T3/<FNXAA^eC?bFR
_26<;:C(I6UCX#.PdE&(8<I(<cgaM6cEcD<@27PQZBPAXC(<GWZ=;J-I;dEC[E2W
FXH2#3DU5PYY0Bab9Q5ZW2e3,P1M^>GCVd,c+@2a_N?PM#\G-c+RVO(BBR0c&SK2
UE\SP6_]S:X+QP=8^FY=a)C3Ed.7gZ#)7LBZ4?Lc2G/JE0)0RZGSPWX5Ua(IgHX:
J1Y3UIOR1N1B^[@GIP_=THCgWKVX(aOJM@39L]TGS,&aHVV2e.T2T_:_)aa?+K)_
@YER\-=+3[<ZUE.86@20g9EaSLCDaRF>Q&O3.BL48F.RfW<VV03]<;@E4[gE=ED=
TALZWNJSXX^]AR@;D8,Y3/QU8[1]6;_=+0f0QP3_Re_5AAQXdSQ1YOO<)HfZJ9&+
+YZX(8JNQ&FEHBH-Q#a::@_5(/.>T8UC6Q@SC&\+HK26XAX_,VXM,YW_d?TB9I.,
??<Ge2+5BI;W[Kf3X834+cZd5I.M#V<5:I5E8-0FF.M/g]@SHXU;@,@;d4/-Hb0J
0;(Q\d84V-0fG4:a;bM#BQ>X#W]gW^aDMCDQ++,5I[f.\DF.UeeW\eR&<5K0BYb9
:&IEHHWb(LNg-Q:bQ1PUVP3B#_UE4RA8+E+R_eMO]-:G6+?>PW092)2V>L5A&NaY
[Ec]dMfe7eEGNH/D(DH4BH0P5Y3GT\.G^WO>]e:B9ZUL),cV_1Y__8\/^\gg12M#
?8cP_e:dbY\HQGDJ8](;&&JM21K59VGeN]9OM@>Qc]QB:\S<:XM=Q>^Y@:#dH6C&
H?_<TadDM?Da2X]O[43Z1E6;S=9UG9.?0ZR4,)5Q9MA/X2+Tf-]d_c-=7(,3fJ5O
L+P]P@E<X0e&1aQTN@8eX;EBVXP9;)<-\f9QIO)?F\?06Ge4;>U;_C-_39AbEaV=
C98:NA=+O29XH0@>>Z)\QHU^EaM\O6bae\K-VU7C4<O9CdI>)2cY,IFNZWA^WP7Q
Q8Y0O]3Pc7.T>);SMfG6>II[233_5N8+BBXVF1<L;HTNZ#CKM9=XN=GDHe]_=B9A
0/9:5NJLWOf41@?X])@^BZ<IG4FTQO(5L=&+4[9A4G[->5OMb6IgC(B1g1FYd+-W
-N)/&aF;aaW4ZFSd_3c9g0K)a,_1/D=?#DJJHf7RIVcfgYEb0C@bYe1=,8MaQ=#1
(]ABF)B?1S)VC4H_^?LV[FCT#&<??AW+2dL.VX/Ma1J^V]T3L3MNL@F.c-.Q5]&6
9f.#GOQ:.cJ^^[:))+)WYL8HJ?6G0;&C@W=5,]P=Z\M.]A=Y=JR//;#=A3]KdK3I
X65[KgKeTZZ2Rfb^aH2BH\3+UF?.GJce5.2N^:a.=4S_Afa/dPH@86)Hgg#-2H7d
)FeLF7O>.NB].a-2TSg4f@8NK[Q6O:.7gM9.@J<-beS,W-E,d[8gSeJLH@(_]64D
EX=B?0OXR,\;R-+fT^]KX;-A/\<PKbCT<)g&#P+4XK;,^?V[Qe0O2K=.E#a:3[0M
P8\)QS21K(+gYPR_#Y@Ce(QG0:DSQb=+8EUQc0;UQU6\<4.dc&6dN@69[9CE3+dc
+#;FA,F<ea1Ob+_PVN;_.HaEISf,ZgbR+-McS-SEf1/(5Y]=/#:1/T-U+[=6O&eX
912RFI5P?P8Rb]^4a1YQ&#VI].Ze)IbEfUU[H\JR,_Rb[#R+#(B4BVY11-Q4,gNZ
GN)0)BdUC^5\H+T20[1J^TH&K2ZJ2L5A5/>Ve2dJ?d)c4SFD]+-<)1.b=9fEL1a<
CSDH;CUF<?8TNd@R2>g\L57ME)IJLQ\0gLVHE5>cZQ.VYN&RCS#1)NN^:^>V,\eD
6]bQOBggEMU/6=Y,aX[Q-B#EG<XN]6(+OF((:M:a@6WZ=ba4^?G30U#3H)&SbdYe
7/EcN[7_?3^b3HCLgM6+V=aGebC6\DWHYgF+.ZRG<He3W&/@9(]<JMV\Y&g9Ib,W
AZd)M^M)._aQI0Z+&CHSBd-GW4,(YT=V?2cg)6HI.5+XZa5OOMaFQ+f1cX3N_Oa4
V@[F6QD]_+TTOA6LK3W?GZTb0+&e7^]M4O?2_Y-HTO+(c)Q3)NG7D22^GE-Ie=KJ
EA4d2]^-a&004-B&aZBH:Y5,F)a)@-NK)g.:-2&+XJ9#=VUSVg8Bf3KA=J6-&3TE
G/1<bT\(gK>NP6#X_-5KJ,Hbe\gBJM(]d41bf:5C:FCc.:-g7]MQ@Y3Ed[RX6XW.
AR1<U4N9,f,C[?Vf<Z\6Q&8O?]Gbc[BOTH(O;A:3NIP)Y_G85J_#I;]E9(cBUNOT
.71BdU]REMN_H:@f6,8;;?U_J&KV??UcC\;d4MIGNK=E;dIG)V#e3F11g():IEMM
^Dc-7AP29;F75SY?844BW,,AYNV3,c,SFRY53<Q.Q<IX2C/#3+]\@VES8cHBS0_S
b5M>ReUdEaX45_0/K@L-]=aLI@V?Y)J^J=5bC(1Q8Z]37f1gY7Q#@)>8g&a8^cAM
+a]4I[AZE5]\^DC2K)+&CTSM59IdQ()3e9FU?0@A(G,Ie8=7P:1R,A_UE,C3-7H1
NP9A/@NL\Vc](@+#+1+V:Z;Q^#,?fN2DIRW;/2B^e3U^/7&Xac3PU]H./-PH\49?
6GaUM/>Q\LI]@g#;1[)##ZI<Q0Gf2e3<b+XPO3T_KA1B@S_cc/GaW[^)&/9M,X^V
_][9d#KDA.H/]OeV/8_eWFD5V>QFQ9P+=^#:.<CQ;0:5TMN1RBZ:RK:94J@Ed9GV
^Y43USDgd(\g]WaN-J;:<BKOaP8WC>Q23_Q1PFCG8&<-2Q6SZGI5H]+7/TPX]K]Q
#D#]&&E/^=NQd;\RKCQf8GP^6O1+<MX0SR3.ML.cdd[@?Cc#A#LecX3I>1Vf._bQ
b=<WP,#LD/1D<>O>QS>2]af+QE3,bEYd^CP+N48Fg>551c5=,@JDM^]6g&OU(#EF
:Sf]Q=K:E;:Tg-#=35>3CR[VK43,JP<gQdQ?fP#R;9-3M@fO8L>PS+;)03g6NZ@:
b5R2<3P5X2]=g7\=2Q[fTeSZURMX4Q^UL8WQ,?a@JVGWPW]5,3d-F4NI.@K@+2XH
N>aM6fd<caL,G_N0VV5R-=_.V)XJ2IRd>d3bSg93Q?([1V:gbUQE^&LF_M&+@(XL
[.4A/6E,\>3:8^437BL94g)E9&IPOE,3M3eWZ:Sc#3PU.K97,T[<B(:;D,&#8Z]<
Q2g@(4V^M=G>#B?Wg2:N0Ge?/09P+gfUYd0<,\Y-AV0fgLTf<OMVI9=E2F,_<4,?
ObSY:>\6cJebR(H[IE5=AHSJ@_I;W7Ue94.X]>,S-,3?2)>]D&@VMKfT@)X3BCT-
BgUC]&17UcL(4_DI,&)/]M?fZgQMEHaNbMVc?:5KYD&M5Z6D[40>WKCWN(C-N-P4
0X3N6T15ZW5>L^.;TaZP&0Q1_?J,M3g=1XU1W)M==IWg/+F@5]QGY.L4+,1Lb.Fg
5C[L&5<_Zcg5&1>0_:cc.4QC?69gI;@_YDA4>fOe1>1Z]CSNNEQ6XX:>_\)_D#JM
R8&fQAFKb#Y<OQ7O\c#5W2cRgS)FUHDDI:<>#,TI[Q2-JN<2,BE,_]#Y3JBM?=E)
+[9\1^S0@GW-agdbefZDZI[9(LX5.XMNLBS7EfORV/f2A3ZIVLO:@F<(^LJMa73f
219F&-G6:<5-9OJ+\gXB?;Db,NE]E/d<K2K\(.?3MH-U]_TOB/D>f9gF)LZ?:Tb3
^U,,=.;;ObI;;J+;AV-TQJb:SCbHgbKWOFG&31)I0:8B8_7F?JUEXK<TLg.O0&b3
JfFcSZcY].S+a8b+6b2=Nf&fJ89H37HGVeM)_V;NP[&?S50]DfGU3a5K&9]5F]F?
QAI2<UN=N:]Y5,Yd75NA2/&fd<0;\->eU0Wd7<fK-]S#4Z[,T<KcMHM8WA(MC-OM
4CMJRGV]]E:JJT+bPR4)IZ#53ZO[>8,I6[L5?\V:F8#gRZI/Lg?gR4)MV#Wc2@10
Hc1gC7a\\X.WPSVL;N6EKN5T28R:1a@BaJ0G4AJ\S_L+0N+B3N+J3Jd7UW1gC/1/
&0V/ZF8aX/+b\V:K=<OP(D<_N1(.5J?+_4c:\43X0L./TS_#4=eR><(3d35F-&E6
;V-EC,cbRB[^(Cg3aY(0HeBAgW6G8_U@_Yf=B@Kd2g_2;I6:?19OT#BIY([&NS\U
;W]O71AA9Y45N32H5TYO\+KT\\9d55QSO:(XWdNZU4J18a>IR@ARG&cI+7b2P&#J
[]D7EJSf9705a\D9RQJ4./\D9g,5=RBY#RKf_9#Xf=^gYW&1;AHK=Qg3AgG3L\/?
<KW6gf5Pc#&>L;4G+UF(3&eI8H]INWJ#[gN9F5Z-U=Y2KKM&/aaP,,<ZVdG;I@#,
T+3[^Z&S5bH/A5Z4_E:R]N&J5]Q,4[79gBZRFI[&dI82+gRN30TY>Zf6#T#gI&Ua
RPI#E&Y@cJ&T601+:?Md7=B^+YLVW[EQdYMaD+S7cG0F_I4YV9A2U@b),UQHVW;S
ANK-<7.Y#,LV1WUVgaBJ#7V2\P^@.7GaE2(4d.,Fd/e9<8@^P^8CC6PHffUUB4E-
JYI+XUg&J#X29>3gYd(.OQK^]KJ10AS7Mb=CFcD\K8bO]R1)ULe02NAZR&ce<B83
2Q[eH5G]O@;2)d2T7IKLCf>YCb)+bD0LfF,PFLf,Wg.97VHS+8U6J:JDV;C1d+V)
XB8LT3??ZWPCeK4TB(P-62H+[XReWc4_=b_IdQ4JCL(]3R,Y(MA35&Q&[\90IYKV
#JI)^SA51Qg8fHU_G(4Q-JSG9RGID\.TBRFJ__:4Y26b0Xc:;N<b>L>NffE_Z5Z@
&2TPb]QdR0AHLM^c7M^X[Q7GPP=L,L_VU\58&16aF#&W8-bJ]COJ^BBb5._P6G<e
=ff8;\\C@Aa)137FH]b#?#I^3\,]Z_^A_&:+-6&QTJRVV6YO:#e:bL;RJXAPb+^2
.L^e+\]#<MK1(BfR@(H7X&^UJPJV0D:1g65KcOEe@Y[5f3DDbBFF4)^O86+A)fO\
2JHdI/O_cR7g#[-cZ&S=eg;1BV?ZI,C<)JJZbfZ^C0d/G<@^0gYcPKT4[ROR#)G9
L?V/ANXA(g;/133IKY28,,;^G@F:P#ZgH1-]3VR;Yc:9H)I_4Ld&L+AL,H,fc965
_PA]QEf9-5eJ;AX@VIS:b8A1b2W\/MDcb+C<AUPBbFMRSBR2MIO3=#-H4cMNX2^A
-TH-[=(<?TW)fJS;@11O?DK39#JKQbZ8IEK06<R:ZKTD9K@^WX,.B]\PK(A=M+UY
FL6<VZ[4]&&/-G;dFT>J@RPbXBdLZ58>XI,Kf&L&.9;<#aD]c>=Y&OR\Q8LLO[>O
+(eF:,4BI#7F5<.9&)HXJ4DBCLcV=H>T4g),^6gWU;[c<VCSN:AIcb5bC(CUg__B
7B0P.4IfUSda6LWP+IP4gSD2Xg=LIS=ZC-[K)VNTFAI>RWeVC5)Q/M;0A[&<5<A?
\@>fD&Y/4:YaQTfgI_6IV@Q58QQF]:EMYf:J2:2S>8-:[cBB0]B9EeZg:\DVS3>^
[d:8f[-ZaLEZ(8g[ST/1W>.1HQeNDW4T0fP\AC6ITIAELgW.AM.NV#He7;4WaXa@
LPRS0<VcF<<S01\E+[PVY]57GZJDCIc-?O9VA61A/YUOFJ1C43M3f@?DXI57JA/T
XS?_IA,fYLK;A)W?P>;Bc1FNV@D,T76ASJAQ1D=<f<LC3Hd83c=B\KcE7,Y0(@Ye
H_][S+L(YCfRKNZPEU46g&1:CP/Q53a2.I02K1RBYeQ6:0(..WPR\,\Yaf,f:I3(
dQ^:YU?ZT-/?QS2R6<?X(,?-FD^RZ[R3:@,,:)Z/7H@O;]R>]G5JP9,55HL>6\WO
_PFRPFPW6e<_V#]cMDNF=C+0gJJ4,VKNX8cEP:-][db<W)eeC84,IBML3=3].gZV
Z57<]N2;g[;fJcU\7L9f;ELO,_bFGZZKa+2JK4c>(>:+ec98D^VbfDQ4PZN4@8Yg
RKXI2._F#a;QQW4JM;)_1R:PGFfX14b\\X<bOPNbTY/>Y-g)ME1bgRR6X:-^ZDa7
b\L4;aQQJ93??Q?EE-/ZA6HgCD_;>]1,>g.1LFJ&H4&X.Pa/H3I[a)\3.6YE42#G
40W84<0E:7VSTS/2]8\J]=M8KB^P#KQ(K6cfdQ@LQ)/.QfV28b=)f;/-4K4LfGG4
f=E3V=EfOCD8S=9+YR.4&fN?/fDa(,B=@>(8W_\ZDCOX:O2[ff+.UZe7SADc2-H1
FcbCTgc(FXgZXF,J)(#8EBB,/C&ScE5E&=KD4F6,Q5A[7e>Mg4Rde)+1gg#VZOd+
K]VIBK(0_8]W.bc(c885Qd<A3Zd[5]a/-XY6@]1LEM4WSY2Vcc(C+E?FYY?D&<,>
OX8W)5YJ<C#B7T61BA[C/(9f_dV7WU;:PH]=.N:(GGXdb2_(cP30):I&e:60EB/D
0ZX02,/G5B[MQ5:54OgZH)VG_1;fMd)7K8:R@X]#FCO0d=;;OafH>)C)M)9().<G
7.OY52XZOGYN<@^\E937]e86);EO>fQ.FY9<W^X6O@FMZGggIZ+_>&-WO=QL]X(W
aJB;2DMY9:,61CA0U.P#.K#g67eYBGS]#^.4/O<87V_3Y?d]S//GUe\T3F^-LPS+
BPVD@[f(@dUU2XV&NL[K7ad>T_.+(^F5?,H7IT<#ZfNX4ULaYO5#G=0]fWbRc(P@
<G1A[Hc<c.86OaH0H)K/_MQUaeccF/355[QfKLEdQX\B?W,^6[b,IHSb3F&N?SJf
<7=M,BQX9g57Q5]DbP\E+g_VeQ,f&2ED+bJ2K6->WXYWZ\X#Y/OTRdZGN522OXIY
3ZII_3a=-0g@B<T<]+:@(X:WN^Nd<,D=71^-5&XC_+ZS32FX35HT&gH37R#f?4+5
W19^dD1O)R1BJ2?V>Fg&U8EZ@>^HNa;g[0T[;Y#S1_IK#]BBMBHFUS)g(=R>E@J8
fD:-[b6a^Z#:f0S^R0M2M/8;0Y\TY7d><Dcd.DgUcWCSC]EO_F#MKa))c/;1@Z:K
ZQ=eQS<8eK1/#JCaeRBZ\@<C7&66JCBf]c]TAUg1TQ&7B.3G0<](a^;U3V:AeW4S
KSB0e9cQ;I(PWQ9?^6_57E>MT5/?=g#G(e79TKRWF72==Qf0LD6KN.ZN8F4\ZS>@
<gf_0ZeNETc6MUX0Y=<UWW>M4$
`endprotected

// -----------------------------------------------------------------------------
`protected
@Te+^V,C6e=9P7@MOT&J?8VS7?9)A#OU8gSQAeOOd2?,-+OFg(>3-)SX2\?ZV>OH
FS(H08+UB_)9*$
`endprotected

//vcs_lic_vip_protect
  `protected
<T6<CQ8#Ae?&?@XQ(fbd\1cUV<a0CT1[:De3O5:Y(U?Lcd0&\af0+(D.]GBg+CKb
=039U)D8=Tada5^T/+=@dH=&R,)/^72UP<]Z/4J455QKF:B26=96D7^Og78?6@37
X3bM@=dW,4_eB:NA-KAV9UO_BF+D_=;[HfZP_=)&59UW_-N8GY=e/JJU5#8UdH6-
:3SBL^UMcXIOR4X>HV=-Z-+L?[DgPQ#fSLNIb3fCU@f=8R:fWYEd<H>@LH]g&^&d
(:M1@=PPfQDc+G_F=]:Hd=dWBWQGbZ_>^4bF3UFPKEY3AKSJ)S1ge85Xa(H?=g-@
@JTPNff(g2402/eGD+23HL@-F3(a[fg>fZ_PFBdd-]/1Z]Ec2=(@IEeL-A_3>fCQ
b>^c#Y=\/Y:XH3g3]<V/[fbd\[O5<3W(6>d]LR38<0ZE,L339c/D41__dE]R;+/0
.bM<fL:IH9d;D9)W&,HBU+Y9#]T2)PGb+eMVKOg6Da&SNb@&d]XJ^=GG0B:W2>/Z
#J88gEU@_Hggb>UFa_&+9:K1Q1cGZfW(BgO58@?^&CG+Y/J51WK;0O\JR:LbOf.2
72PM]_)N]Tg9PXTIDG]88YVCYe+PcgNWY?&f/JTQ]3A91L5MF]S-f_ANIYF@/84<
V54+)+P/2P#7Y3+KKARXMEXNTH8Y9YC6H\(0(K4JZSWL&c6Ge+[J+&_&+J-d+Kb<
B[8:3[9,/_8Cd8/:c;A<1.M&2)ZJDX?L,9B^W0]g=b4,fC+P=^>EfE#7C<@CdQ?O
_-?J,C.cI9I?]<ae\Z;/O\gUZ0.O(HI)D8.GIg/D1T-:^AQ7NTbE=F:g)ZSfa+JI
Y,TRXP#1T)eMP>KK]\F(Q7\+2EPe>aXD<cMZ;2R=((US>J]3KDgMVbHAL/F:eZ43
U8I:6ZNRb-ffCZ)F6;YT&F1#OD:+#FC6(6Mg/J,9f8D8^1c_D?>065[BD1N=:\^^
HAOE-&_eKg&-U[KE:-W0A1[.66FHTFfGBH04-3I;aM[,S;e[6a2--Te>A2:ZG76M
2c]_a1=X.&4a2534DNf[8?K2H(-N&]QROdC].f<G(KE;R=B9FK)=M2WM27OP>Qbe
&;AXRM[XUR6+>FY)2?BMWO,/C8U_/Fb^?0b8O^6@a.08OJN>;;c_&[A0EEB>a=>SQ$
`endprotected

`protected
bXLULUFU@0)bZ5231f^FUT;[P70_gMe:TSETOR_6MMZSMEEdC7X2()CS=A@IP_,\
d(K40e/X<B=UbO^T1RKP5_29gX=\-@TbIfW>VLb0aH(SE$
`endprotected

//vcs_lic_vip_protect
  `protected
9cIA=&eHd4E=>G54OTZ1+Y3=:=HK<^Ve4I/=N)f@&][MC?4bJW#[((@;f0,-L:\7
BH<ZG/fc-a,N+I7K5Pcc&bdISVe,C=X@VCGEOK^<1:0#W,70B0=Y+?CAZ/=bE2-e
3BW9EgY?J/P;G/X_8/4S,F9P=dcPTYY\FAKe04.7=+1.fJAJ^0_NAZ5?3A1#)C@H
gC,d[/31LeT2C+?c5Uf/76C:gfeF5DR0\SA+LJ+:L?V@P\WRP\Wc3VYFN;<eCPPW
[8L9-WdPYd+N]R?8G3M<QB&<QE_]<c@b@ED^4G-46[,TI3Y124BcDD),S[OMSB8>
g.[2.(#HU6A=>d_3GU^NF:+/JDQ[XPK?)AM&Y6ZJNOY?P14P3(Ib<;33W9gJ,\UR
dY#PX44/?R1MIb?e3?O9:Yf11\aIUF7S4,E-\>==.H<E/(K=;:,bZ.=B&UIgdI[M
gG-?-R;Dc\.?^BfII-X)8)g_aFeSUG4XE8gb0/HIea9RR@]7gK.cL(LKW\+#S3(0
OQBH&:BA.c=?5=Q\)-EWD9)Bg_+_CN@T>@#^OEee.PMeV9aaSRf5PU]&MOPY=T56
;P4:@^>UX.O[+c0(b+0A]Ca_BA(PZ4#S)F7>g^d^(;b>QG)FP.CbK8<(0ZUa?,aC
P2?eg9#US2P1+3Z/-TE@NEGE?LAV1<1eM#/[d><+\2BOf#&[F#D:R35fT1\gfUFL
fFY[V[.U\a00d8^FI0.6TZ=:URI>3/B-f)9^-;X0RP>8XbJHI@_[V@VC8&EO(2+@
81KA5bHL?dA_RDX,eT;+<GZZ]UB/+-S#16H.;bJ&6ZQ716b[&@Z-,)Sb^Od<:LUa
NaCIF(,XX>a&B2D;C4+=1-5-ABB,(gUT2ZXCCF/>-KMbVC1Ma/:7Z;]-Ida,#)D-
KQ_e#:TBJ=8GGKafJ2d+-a\AZ;[6MU,5#ANBFf2F>0d52Ba]Ng2NCRf4,=0]]M/[
Y6:b0eL?>BY[SO[@>_:(OG>L2K(._YP\TZB#b,8Z<Y[VKS+bY13>#ICa(b@\IP<6
S0,ITc#/g>-)]caH_Y=(?RRUYSQ_FHg.HZDd74]8U4.:_9[[]B=T^UNS8-R7dSFV
PETbF8TYLKE6XTMB;0J+7E79dNJE&])4L4dO\SD]9JY)HEDa\M0ea,&FALJO12VJ
NGWcBc[d,fAff:EV]eDJ9R8MH=Z<JMP8e[]]SHNA@c3OU_LC3fSKE0\\SM/+TDad
6A]bbf80MKa628-XO9PCJNc@_F^\)Y&0P^4)S@1,>b[&>0MR+DW=JA#a)86URAMX
2?+<Zcd6&V4EG(3PY?\a47C#4LRUM1BYMG2XL6bS?A)&8IQJ2WZ_@Oe;UO@cJ/Z7
OKbbE\,<??H#)V)@(MIbA+4Ue?O2T.eTee(g@VY86fcLP[cX;]J38H2X9aM?J;2J
>aL:[@&1M-B5^68\8GeT;J1[4,]E2U-06d;O1I430CA^M6?MWN,0M0#&CNaccUOe
I2=VW[<A,S>\,>BH=[bc,dE0#cYHe^:0(/>1Z&GPN9S65e>C0\G=Ye/^QI<SG^:B
<\4VY>P-a.7,eM,cQX5gcF)99.<GE.?,Z2JXKU@?&_<C^5Ld9^8=KO]B?HCRIU3\
2POA(<Bc7(,C?W>ZP52c\HE,Q64]SC])?UF1Z//8cH4-MWEF@H?fgI;H;K[FE+6S
#/9;&cX;H-eDE/32Q(9Jg/]I567I2E.AFZAdB9C64FfHJ(PKO&@ZQG_2UP]eC;X2
^_X-IYKRSUTf4AbG/-4\DfD0K(ca&_b3&4bNJ+77V)@d(AaKKCdZE[G][QZ-A^L(
#^UF+:aCM&-Eb\]L:2-fM@,/5=dKQ<U<1CdS.AFJ7P\TXFRNEIbX]IVZCSMI3WE)
d>c65b6_G:QH0>=:/(7@c8YL-7=-VOd#JN)W7=SeQ[T-0;aCYE6,RgB0WdAg(cDe
Q-H-PMH,/[P_0d<N_Zd6\#J=^GO[(,#L)6^1FaF_V31M<CROI\T20Y,bXc52^,9e
G0HNaKVbDcTFVXKa=1>>Z,WV0\MaIaAC6,.KIa4gCO#N@M9e;E+QCVfIP_B+bGQ?
/Y4^\G+.12SO3V2Db2;[:,-@Y:7CLc\40(AF#6QM<U9VS3MV_=\+],,ZYIA3UAEg
Q1J0/>K.NVW#U]U/SDK5UHI5TWf>LR7U61@D1;/5)2?6;;AZd,\KQ,(P,eRRA16W
]HO>\BY,BTH6]=Q9=9#TAR5P,,c@MEW7W?+2)MeYMe)63Q_5CK]M7>ZN;8W[5bG-
E9)2-C0Ac9G0:DFIf6#YVB3/X=SRW&M[-f7F6ZUM1ECB2=;c@?]JGA;g)/F0b3Y<
8N)\^e-=R)=.aK)7AGaYN?FL[8;R<e8]_GRZ7A.TEcN.)0IN:fT>V^eE[29:7[\C
7Ja>4E_L1=4E_DLSFM];2+8A0]B&H4Y79@JRDSJ?3[a418V)3&d5c0ADL:fW5-c.
5+Z05G3d1^7,cf]9RgVGSX0c6D+a,6H-@S&7=@\fVD[K:PV2b:a63)8,DFVf^FC[
+Y0=26OUf@YSeF+VOD-T-Ff(3_:IZ?F8:SBT^;K9L.dNGC,2:5[C8aMc)J6E4-)=
EINUMIDg0Z-G(U68Zg8+2()P0QS(WES0OYZZ+O5RH\WSN[EIG=KKCPf0CV2BAbB<
5/+1>_.cXg/CHF7,_c=&fd@>\,[>MSdfQ;16IAdA6[]3DKO1M6DNVBd],MI;LI.1
A:F7+MS69<791fF5Y9AF7P-WP@:?UCFOJ1++DI)dHJX8FN.S+C-9eSVQ?Y34e+>:
/;D0_8T(c9]G^O#@g67QSB.7FDI4e+=2,6I#<N547L&6O8JbAgHO&))GVS-/2\)J
X]+4JT=J>=-dJS/X=f4gagQG9ZQ\QZMRMcYN4+ZO02CGS1SM.#e=fTSQQ3PFYI8H
[1@DMNM[Q<c-1\AY)g6=],AA^(\R><dX\@;\;JL)2&cYdSMAOT&fYC@9G2ZS([H@
&1^)LBPED?R#3J8MSEX@bQ#87Q]DeYXUE,BG5R,N&>T,fZHZCSKKPL/JbQK&bM,>
f=6_A-X6DVZ=\_abb38DUKA]VO^2(>.Nc(<LCSKcJ3J<J\#JdF2PDad^^JWgZ]4C
-[@F]4C#?agc[6+C70f-228-NgMA6+CReFefTDa3+Q3T,>&&9(5b2bbX>=^7@W#-
2BURH6f;D3S.;X]62;6](/JA0I1>UgY-I)>:3d^PJf[bGWQ.\+R@IT8J3dcEC6QP
XJaE/7/dQ0P0TQgT<]#>0OSbN^DaGZaC4]U\76)@OBO0Rf>=6GY@J:?,4151K;]6
T6/\dH2cBI>.@AEVLY?PK0I5+VJDcE:7/YH:CC&O2;LeU3C2H@8.A(([LK\a9/()
\,3)4/[e_cZA:eaC[BHb8/Cd<4M)3a=DYAW-ee8f^=7X2U#g=<::C7CAA:1A:QaS
6PO),_KD?P,@bC\AfT&L:+495L(fQ+C4-\_A2PRA]O2X_FgD-RLHP(<;A-\;79C\
2IeK>9=YG:.HD]Ygd+06Z8&N.98.)IB/fgJABM4D69R<Nf@B^+(9I2&Vc99ee:UA
LfC2>6@?@/T:gTT0TAA+5E=AFS))78P,c>&gg@R&IeRKZ)^VIbDb8BR4^8H1(/-_
-?J.MgXAY+^<HH4MVfcY+f2J[)GbS)\T-Z)VL?R6<\2aHTH&<\X5Re815c1PaIQP
XC_NYEXad_ab[<QZ5PP-<\gb[]KJG4ZA>CRVMW?]FI>ed^IB_@1T2ED;c8]YU1)Q
dYgG>3Y_R8/D@3Ld.9AcM:A_fD=[aV92Jg:G@/H_WH/.TUF[Ed5+dQ[V]4OfVLYd
,S\O]#7bFLgK[#15(.(RRO+e,gQ]U/)f845X)+_bO-gVg?@FIC/NIC,A4I#Z3;2Q
1VK/U^WTaWg@4N/87J;&LQ/a0M8^=^SEPZX6T5KAc,_YSP)353[WcZ_8<U+_MK>@
X3IGGB&76(;,HH67]efYMLA6d&N.WTQY2g^=?V&#-3B4OeB+]091MK1_f\NIY14&
ML]9LPECBU2VP<\P@R8MJ6-INP[UP^baR2VVbP]aU=9\LM\N7O:X_#HN&0RVGHH]
M=V7.Qa)K)O+\eEd^1K^HQQ879D/:G^/AZ-N^b/AdC&TMS3;RQO@)3eRZV(64#QR
e;]JRd[3]9aXXWNEAf@9f@?[SZeB+/K[-gdcfODgb#[:S1FWMWA9M(W=,\g\US(#
_MATG8U]O[2TY\P]R=02YS);9FP/-;fE&ge;GAc+)RZP.)+.)H66?5XDHA4VN7))
;FF^a_X8FY6^1[6];65ESLeR(aa/]^UGI9[ND-W\P4+/@GbV^eHA=)Dc=CM&&#N^
94A54#>W>YeI\TU@7XC1196g1R>&?b7#a=[:eRQ?9+]Z3U5&VSE]A/6:>.1e&<Ub
eGVGN\NTga[@[4G(25F66SU8Md,II-+d&X5N,<][IPGV.++]G&G.L/Mg/@86;bMV
T^DGCY0F2>G:.^9>,E-L>JFgG9FB(0>V8>4AA23>3a+RV;f2H+D.17T\f4bR&HNK
<0F7fUV(JY/F<JgF>=19^MeH?Tc-G3P>IM0+;F=dcF]0[[=QBU(FQ])cQ_a+(B?X
OFUV6b7\)\SHSJQH_ac^<9/JT.L.XARN[E]_YTB,)U;[SR39Z_T#-ff-gQ&&&5aa
cgA>?_O8/.G3UcZM+5eg0Q#;HT^N5OR;fQ=fRVN3c)SM=@I;DZE.DIS[X2d=>^:H
><-IIB=Gfa47e9=KJ-EKM4K(T^5UX=E,e/96BFgD<:g&fQ?<KL?\f+/c9a7:LRA]
SF[NOZ2=I7AM5X:&WBL@/U8-&BCcO=Cb-EUSA+]QBT]5@RHH7>IYP;=aNKI&ZNMR
)X/d31^H:Qd#50@DKa^4+dBJ.0K85L=T#6e#;\-/eZ=1N/aWaKGdR8acQJFeY=JO
Ze@LZ6Q,D4D1QP7HT74]]e0dUH:.H12C&[EJDHZZ@Y&WVd.WMTC^KZ4]P0FLQGd_
#dESDe,PS<W^:b9-96?LRN;=C8IHaUMP,\aL8046_[W;J^UHWU+ebQT[^M4^8;3F
@U1d[>)&eA)EO@)M[MVC,/Q/OI>eb)2d+L(AO::2b&8=XVWT-0aG_U42D#1Vc8Fc
XN3C(6=L>VS8[ME@>=V^&8S_A0a-4R-B6\H;;6BDU5E?18g_H:AN];(&M.=.5/M9
N/US7QZIFOBNGK,KM8/H;+6bd9+AYPH+f3,(FE1=[[-L&H6Q#gC0PgRTEfZe.^25
9L5D7,E\gS;aE4+1I7(TaP\Y1ESC@6F_]S.3O6O58Q[4K8X_4VD/40=R&bM9IY?@
HZ#fBL+9_[-=F:([H(g0GG&]CTVYGH7F6@7BWH=QOI[#S#O7Ab7\=I3N\Z?9GQIR
#1K9:#J;L?(I@Z<<7@,PM6/4g=GR46S\3UXMTVF4T3[8LO<B6NRZ=Uc@]Wegge?R
e=2JPeY0=^H&a9V+3ISc+&=^Pb[=-ZH&/bC3^I,-T8bR&,6F3?Y5.-CRK[ZIL:UO
DMH:B2&U8g#NLL\[<b@cB?If(E>-?DL\,N]Y@[;HTF6S(b+fa#::OaaT,AZg_&Kd
[fDg+QV^-HY2ROFQKCP#)1D/FY/5NH5[E4(6#6#2f)&6:PB#ED>?>RH,0EJFJKV(
)S.CH4U:8#)1T6#FU\d=+&b^ZLA2CZ)gd[Od^^c)9WeI4a;)2gT#1^H:6=8(VO+Y
R4S?2BSA=8/Q;<=@<6C0PXE=3[S:O;ccGO]KS1JBT0LPbGX:<;9(7eBT,=fXMb9Y
eD[JP_9HTI&::KGSOac@&63I02VgZZL4JD49aIS;/E703(XW#a(@B^bX3+RN=WY2
/G>U6JUMTFT.:+T^G+KVg3O-ZK0ZL.A?/4R:f3eMc[d\OV21f89;6fL1Y546:PFR
PK)+OM&Ma-g\SDZEJf)HXYZ#g@>/+cM4HHCIZW/DEcg#48?;Va3-F&\^F6)2A6,d
Y<Fe90[RI2M5Y]31/[#^^YORXXP-6VD-Q=:;f3L9I23(&5e_0,+4e(K4=FS3N[NB
^.Y>>TY&Y;^E)c&-5X3RK<FS)9TG-&JY-;7;9&122;?H\:@8BNUd;V/-VcRYNFVg
V.CF4X>Zae>RW#HNC,3VGV2F\UCU_V\fb\9c^[86LPRL.+T8A[/NN2L-B@If57fC
,T/1fG@Ag?O.ECU:)RCLYE9C4WX)[T.NN^GXI,]f@/@-E<U3:<M.#9Ga@<>MS456
U<41)JfE2>_.e-R(CZ97MKaSGV]7D8XBQXQ8701PXEc0733UJLN]].7#PP7]Z/X>
=NXRU]ZgUY4)_gVS9]ge^OPd;V@AU?[#O&FDH#@3KV^7I@c-[d?8]^T;1(#XMeBL
C@,,=0+G]10I2O61LOG_MP>I0>8#Z3:Q+[3I1X]E,]&WD#^LA>bg/:e2T6@:Z&.9
V79BEB0.V7&4N7SEBE&UY-1XbJK6K&gI,C_:M0XU>D5,3VXUP3Sf5<#F=P=cBW1G
O3Mf-3,8CS^RFGGfcN?1/6LQ/YC-McTE5P@CF=P7S61<1;H7c4R1-B?^[GLd55]9
Ra7+dJ_L(_-ZSJ-SRWHb1YP&+(X?3d1@MNQRBR6+eTS9MNE(@.3--?B0A^Q1A,@f
IHMP^[Z4eK7U=I]M5D7.?a9I.B,H2+RZDfL4?aEa;aV\3JOQG5_M@/U>N1GCaW-A
M-V,FR)c54<2DQSZ=^QC#+:7G/,ZP3L5=\]?Ta<O-H1K2a9D=Hc6\+>0?N9^Z:ZR
4(#LK:]SB3KN90G+-&[(;6+KKD><^+P)=)ZP0@@7@-]O(fc).5Z,#bRP;<UCZYfa
M\-f1UCL88gH>[8dcJDL+1VL97NeDAS]2,8\b4,f.NgGL;#O/;,a5P&<&;0A@N?F
^.OCd9(Jc=IdKGO,9M8Ib>=CP/NC]8^3(H5,[&:1bRX@RaV7M(<3-+Z>:Y]OfB>#
AL7\NIB?:TF:=:ZK[.TME(USYVU-G>F8IGVQ.c=J5P^IM2dcQ&aAdE3Y1=8_P.<0
4O>L?JFQ8Z2cV423?5]@0g,P,(NYD1URRZ-;)PWYc)QIfNTaS1-_C3C^=NG8/+FW
#C(Nc20aX@TO#02?CH^bW^C-;L:0b#ZD<KE(=cL@#;.N4@9[Ea_AS:VUfcQ8NN[D
Z#L5MCL=Bd=1^.K^EgR^dY?N0M8a8dIC@Q=WbV+.V\,&3B&>(6?eTF5.Mg,[>PO:
b]Q2_(V6[C+e;0<c:RUS32aVN1G)M=]I9f[]^WYO.M6JO+1\)\N5T4b(+1RZC0=,
L1ZS:DWTQ/9D&f^+9L&^PNRCRCH^>QVFH#D0W#Y89DLSTQWHfS6<I(E<f2I-DIN.
5dRHXZI,FgfI_0.30N-HT@@b6Ad#/==Q?KRP1BM970G;;.XT)L5N8(79\cLH@U2e
]@)=#5R@If54]=]d[FF/]0bAd8+\I]P14[57gEJ:H]=YS,4G&TcY7=RD44B(fO_J
70FO>8,aW.G]8?=FA(d4R[g/(GS\0Y=.77]^;g:^40=G4-b+.?1]OE#Y^S_F-#9)
)H.W;YbTDb7bUZD#VE)4OZ\)1Q@A_RUg217WgJIQK:C>b)cSgL(-NUdXcLXaF5;X
TS/gVT_6b7Vb#CI@+T#YHIK;/FV::ZWd5GOE1?W+8d]8HR1K4+JN]N[HLV(E:ZVf
1F2H<F&9B.65XgC7(ScOgZfO_^8\Y<?a?86I(Hg98DV;3OaW[?gSYF4L]NddXKgW
<[e[D(TE.KVX--_dc+5&&^2,T6LcF;@GGd+)G,76C10S]-?E8+YTb]#KQHNQ-g7P
d3E6NV2daBO#cGc\,+g>I?,H8T.&?3);^X7>Jc5T>NBaKZ66.ZJ?\=<U[)=J=J)E
GdL?<2V\OWJgTef/X:W(6B^F:IgTDD]&dDKfQ-62E,_#S&A>\fdG?A@^fa7b>feF
C)Z#5EA(&^V,Z6F18-#),8.\(5V<S7?A[V.[OdB1;N^V059aA/gM8V/4f+J5RN^R
(NJ=f?OB+2F8CWJ./5=ON=e8Y[:8N7HKI<1-Tb1N#2K6M5BD5Y&H=IS;RE?KL+.P
JbRbg8_9[NEH(_0_HZGY&7/-@&7a:J>Be9+VVPU1RHSK_=68/=P^e8-AYf1gCg4&
DI+Qf,P44fB.S@40G7fA&][)GMG_(S1S_/7]&O(K:KI]F;5(10[\+@.IO#(KXf(-
E61<]e6<US6JY4DN+e0d.UO;MAF2-E+ZefS9]LZg[G1_F_5f\2\)EUMeRNeN9)_d
VcRX505e:IN.N(&7@8REI0Y61BW@c2#60NY^MS)H[Q\=&67gJ=-WF)U4.8QG\<L<
e^[H482=,;LWQcH3E?Y-35/YaR8<I8SGa22Qc<.-]d0_6:JQFF[=6QaPG6Re]:_#
)62FKSQf<=bcN.)&U)+W7^[9Dd:9/_:dSA&cY5E:G8&<_2RXeg[:WS=cHe,G)bZ&
b9deC(8d)_YM=.aJ9.3MUTP&?8WScIRVJA&4ENTQgAW.a+,:V_3#^UXY0F,#)9?0
87S7#Yc_a68I_B<N?e+(d40DDKaR^W1VFJ^2B@Bf(d<NP@[P6Vg3#,7_QWcZNEeN
-VC\_K).US>31?:a_efR^/\X-,MN#4d#4Kb_OI^)I?Ke<B@,Yc:L94L2)PWV7DQ#
)DaRMd?NB6\H\26X97K^a7QYT8bH)G6F,L+@e01J;L\-R1d4ab?S16Y(Z=TF>1@#
bJQ1V[\.:_(>a0T1c&N5d0>:5g4Z\>.QO):-g.P/eK1M9O?W/MUfKdc6IgKfH9,e
RW[J_XDS1\?;@YE]G1]SD\D&T0\aKY;?cTZN[EXVHG;5bW_)V5/;N1B\0\UL-dO7
,ec7W&DcM6;AL=^;a178[=ScW2QY5ga;NDN(IFGGNFc.]],8e?GW):7UB&+RCD=6
3TKaPL,7PE(c;7P#:5=32M#6ZZe2#Q9B[9UJ3LW61CF:Y^1X0gFZ.[;,d,;@c-G,
1I\US\CNcH2>/e&IU+=OI+^DUb1K8bKN#KP:4]H=H-A+IV=]8W+=+]<X0T9T7OH_
<FIXdff(4MfY8e+Ba.R>>?#4Y[e[\(SLZFK9DEU5H]/=A0<LJV;_X3ZY-2.CAG:M
-/P_8)YH.(;HRfEX(57:c8;6eE?I#440PgaG+K8A2e^d])-<5546YD0[cB6PK/X_
[QVML3(3#M(=:[d5&2UDY.9Re]:g,&6fPUZI?f4#SQQF&G176#XHOFcRFb..g6KD
]QO(/26^BdB6b88aE:002[LESeY-0#^_cKKM8?X]2NXE_Y<dfb_IS/L].gA=?,cW
O6YG_-+KH\T)\-FFN-JgSM8a9\,X8\A21O=?6-@,^\-23JNFYLe:0B2,ZT^1b4_9
V#>3NC0TN.T/@1fBXCF^Q/XXAVD6A+XB&D-e+Lf51QN/XPFXE:(E154Z6+>@@06/
40@X3:4@IgbU\gIa\4bb05@dBAJaFQY.DYd0;Ug8E3;eSMb<\B)c9DO@0<O-)>#@
JcNd7;/NR:VUWSDc.@AV_dT.=C),WKcZ;)^?MTG+<ZPWJ,OdBX/Q1VC&U/EXQWF6
<NQ48)@[3QZ)P9]>?(:(K3[BRKJ#N+5]T[-X&#MW]H]&#(C7G>3H.#de9<@dJL5?
[XQ-KVOD\[P>@b-?gU[8+.8eH\3R+(IKKAPQB:W+Q);UT&DC[M0&#8COgOI1#4][
<J@PaNG)9TUGH;._^g--Y^I4TPWE-<N0YVI;,C;&IQTDJG<.K01>>T[ACZBQdR]<
)_0[a^UOG20e:Yf2DHU?g-Yd.PM(#\<)3:a?A4gM3QNOVPaLKMJST^/RAcTVd-_/
Nb8#_>M;)5:0Aa=+YcO/Q<T\,KfVD^5C<MJSW:U68=K:1@:0L98U97<bP.P/UADb
@\Uc#U943CV&c=7,UZII1A4gVC<2I^L?TD/4:2Y]6Y1#Q^F1WRQDJZaH#?Q+?/a8
G8g#<K[8<#3g,@P</+6<0SN&7b+937DE3G\,9HVO4J8T;,@gd#:.gd-<#7HVbS-)
;><EP6A<9=#cS_UW#>IEO30Ee@3g,b/:=+ZDE7b4\I&7FY)^a(a0KJWY2L/fW#]&
SX_WED+]C;8F42cD[?^OF<<S_STZ=\E]JO.^cD[aS=Df8PK5QLGSa\XY=e9b<F05
0SN#1?V\MZVW&.+e>8_I9)EDT55H\TcINDYH39YDeDHGMH#4[BXY80f)fQb+HJ9b
a1Fdg?Ec(L4X1RX+-Nc.K5;d[]Y+F:Xa5;AO(S\H8[:=B#-JQ0P@geDKO98+U@g)
<6K66?d5?4(I#/3].P(=9FFYGdF5?Q\dTZB,TLUAHKL)^7<<E(G:_QO@TE_aB)O)
Kdd0/HH=PD:UW/(AM\9b[SS?,BI@L,N4CbCP4^@3:\A;X45W8+O0FLG=[;\deXJ<
H0J?SWJT=)2V40bBO)=LOU2d4-@B>^LLJT.V)_URCN6PS4T5(YUQOBD)QX&LG[(<
34bV&\:?+M@(b0QTS)F8LX.\?#78ATe81O]A=OF;aBKQ_N7HOF^;HO/6V2=^1dHG
Z6Rad_J/1#6TI#GQ.Og>3C0,g9+Fe[LM-<HNRN11G\N&QI[#UCb,1UfGe>#^FY8#
4FICHNIYCgI(M7G5T716D:E(<S<S:<;FbWa_#R=]S4C4,a8C;&G7,SQ#?</1O7FN
);W@dQP:R7e0MR774<T#YLL9MJD0JPIe96.@J?^KO8,BA/8G</\7?M8J?[Yd3)cN
YIXZA=EFgAH.8V&D;.O<@GU<7INUUe#QT,@O=\(#K,c](fG@;D1WX\>@DDf@UC71
45gQ.,Df]^?XgUQ18-+e1Hd+(6:-9I;-5GENB,U/<BZVED.G\SO\&J0f.C1QcBM;
c7(U^GfKGY^aF+@[H)3-(_=-OF7/+TPQOFNBc,=S1RXR_FN&4Z+(?-:=fOCCT[bV
.eg2bOBQU@;_<#&MT29IU9PY/aIfd.M#Y(IU]Y5NL7)NeO?>+M=)Y9&HFEFJ.FX_
6CJ[.2RNJNUI;+.3gK@(4R4E&:ALG<V20FWH]MXb=&)[HL8]DSA02MBaHU2[0&6R
\Wf3[<YdL02JR7?Z?V?Z8K;-@L:2IPQ]<NC,:05G-5?ZJW<C:YNW@\DV+cdDZ1Ab
f4\.4OQ.YI;9@)B(>8E7;PKa1g:P4C.R[H1FL28X])@GdTL4AL8;,.@2eT:7+):#
Tc9F>.TX@feR<c;4^aB<?a55ED50dT\4L^R58?gg_7DaYfZS1CUf1:P=@AUb7<:#
A1c?;O5.,#E2UB,X?ND,BM]8L2[&->5J;3>SA#g^QTYQ&afcEVO]_PdBIbOeQDA;
.M.C5WN7?&FQ=+8C>\K-NB_GB\9V5efIG84(eUS]Ng<&4FL2K3S^.TC6;W:9_gS9
YV/8MM8SdT.Q<B7@dMGTHG-3QGOZ(O?(d1ge?3)#SKG.PQ-P?KRE6OXEZMQ/b6XB
)1_SfJJ83Ce#c1#=PNGA3[8b];#?0@R<#60W_cA=<O<SE</;0R;AE\fdgf7Z54;S
_7A7aUY?(F3]MGE81-0cHBC^^W.LB2FUMPPafa/+Ta@2W9SbHBfbP)ET--\>]/4=
U?3cXGg)?Ea_HDSAD3g99a9eXO:YJUQ]7F,b,.]&;.&9KB=:QDTRMT66O]]dT^<+
LI^=X1^APN8ROWCHg2#6XP/EPOEg9eO5)])H3RM\N(eS^3C03V2FYM_G)@2;BUQ3
.:G+,=E)KKAgdM9&Z5ge?JWPD#E7^TTBg2/JfH&gAaecYQ+]C:/W:@T-gTI[#-_A
T\#NL<V/OJW^+4K]f:LgM^d[^>_dbEL&L_@@S1U9Gd[.N=F^eWf,<KP:#,NJ_5LF
,BeaBNCY_(?9^Gf<YE4ZY:Q>9KW#ESf#/.ceYRYUga1[KEA=Db3FQR=e<MA3=LIE
5GMf6JCTJ&fV+MN\JUXX?4,g96^>MeV1&#X>?NEdEU-:;5\c:63(C#U46&c-J\E2
CGb3_-QNPC@Q<NH&^K;_::RH]Z]cXIE<AO9_\UA@J/D&EfH=OCa6[1Q8\^9f\GWD
gP0KBf=gFW-OdM\fg8+.Z1#H:)7E0]/eef65)0O]EfMD-0PUQ;Z.ed-d94VK@;aR
G1a;NI^FB[KaCX^_GHP3+?KAA6e?\bAI@QM&/0KKWG6\,))=0]B_E4HK//V>J:6G
=.+8+Dd^?1[L_YLec?7Kf;UXM[>+-15>MW-6C</bYU;fg]a,=IR>8JJ?=H#JID-d
cVgV^IMMTEaGbX1E3:Z/a+1d+M)]&eZTT(ecgQ3.P?a[UZTUSY]MVCX^@<;M;4_Y
Q_H;S/#BYRHX:1N9CIXQgMb7]9RU=7T8&f@=97_6>4bO)WN-BF5e?_37f;+7)Ae/
8Xf>>;=2S5V/VFWcGT\eK3+-deT?g^90#&:O)X<&^_Y&BH_AbZ7Q1IW53?NZB\_3
f/5@dT3+C6P2I1a2O9?L(_]9(,/[;VY1.Y^@MRe&TR\43:-+7YOD]LATS/4G^W-=
D.5L_3IVX/S/CN>V,45eg_\6_0AfXEg?WC5.7c31?P&c_<=MEF]IQCFOJcCT1XP4
(^.H71\+NMFGKbOa(f3CTZ+;@JGA]Tdf5SJ-1?<6Y2G4We7WM&FH/25S2C)3<=2[
._[V@e_IMUBX_^R2?ALHHM&(1Y4\IIdV&Na-,H1a+:LO9)KDLbc,[f@7M0K>06)Z
)8VYAWMQ13.G^&PBZ)/(I\QVaf:=,06Y1aM=(=+WJS:Z:T4ZN/d7b1Z#ZaSI#G<@
f3/a:+K+O<UOcJ_R-R4LUPXE\>]Ye&S7D:85YXOA7cPaGO#Of<V6DL0e;ZW,aLGK
CHB+N@87-8RV](4<23U]cfR6S1)@^U/.-N6JPZeV[A2S8fCd3B0cC/WLLR9@-#IA
-GaD>?G^Ea]4P2ID1:(\<f>;cYHZFA)G[-W[X&^II:gI,Eg4\XRP^/RXc>@BXW?_
a)PI(Ae28eX?V3S)PGF46IM8#::Mb<5:gMQ:2f,HefI(<)=O-A-N0M7ORI>@L^7Z
G<b<T]WF/,c3OBVLcc_6A(S)TRAN<=6Q]JT^5-Y;R#T/eNdeJWL-FD)_DO](7H37
L?KEN(6Wc4PCMUd/BU?LJQ\+_0\gTFG)0/aScIV&]eb1JXe/O/)?=#-Ob7CF?X#a
Q,6]NHdDXA6V>]04c=:YQ/=#ABD03>5@WUQ,@<_0DXGdX7,T,.POQI:C?b/]&5a\
//c\E4:3g>]S7,A3K?4^Z>0GJ2HfR:1B(]O]?gd_<U=EeHd(A<A5[J[74Q\]+WU&
O@,>]XCLQb7Va_g,@;F,/efKbNTZR?KB0AC>=dG0P(;+HWcUcS;4,XSDTf,CdH=/
9OCYO2==UK/8BQGgHe7CA#4VV3Xb3R[1WHJa+238_)7)3O]+=W(PHa9g8gY,MF(:
d1,SH>4T@_I.N2=IB7UUVI-([H=+I__QXMQ@9^,ORDI9Bbbc4(Q5AW]GOfgD\LW<
P4^8c;+)d?+S/<[dG\X/[=aTQ+AecL@:)&UH0J0O;WWB/;GJg84)#e)E^Gb46]00
-NQ@)LDC/?ZP>S&2DAg=B(S.-Afa[6V-gP6?N;c\)-7P\a@6Zg8(I3Y_><]0<@.?
@1;+&,5:)DSG10I1e<c#PMPQM<Z92Rd?CKF;R_(-U9G&Ja+ePC/EY9S>C9e&TBQ.
@^<+>[&OB896C7V\f&7T>?1BaJ93\9HMMI8A,V;,OfLS5TFR1&X8OPI6/WN_E1[V
PIa4R;+:O&LQBZf[CZS=OJPBXK:NCQ86TC0REC8_7]+YJc&^BRA@eY,_c<c[/.=;
P,8DBMa41K(SKJ2V6T95c@(gV9WL.M6>)c>P\)DBQ<@eJ#4UI\)&^b2G^J)]<(X6
6>-_.BA#+777Q]MYNU9T=eCMH<M7,eLf/MaF]P7X<6#5cMPU:DP_OJ41aMZM5f=2
7+WS:GC^KD<4H7_5=(2d3NM9^]Q(MOU,5a#begffMG?+e+^X#Y@0\K:<eRJOA4_B
:_f8Z^.d#02CG0G1CG4^KEH2gaGV[JHYC]B<A8@4-S2EOVIYELJAc0I2V1FU3EW4
C0TD]W4;G3^Y];[,KT.f=>F;G?T&<=O4CD>(DMA&DML5)5SM)Db@M^WG:KYQ?VFV
E2WGeL@LT^O<Nd+?QVDX.YM:=TVX9O#AM)OMEEd2HXW-4&bLW\=SV[@K:fb.?U)E
_7\b)E&QEN8/_?_K60]G93=)gLZbbLA5\2VZ5CZF-Y<9//<gS+E=\9#3bF_.=>/C
_+.(>RF^ZMRSEOe7<H?\@K?<V7;>&gD\LPIG0M@2GOW<0R5BeNgP,bOTcE<NMYE8
8.+LJ@<4C0)#>Va^8NV/gVT<,F)OOZA#B^#fTHDOK@1gF(1fMcX>dMJP;]^VHAJK
<M)Y?6XO>1GWP1D&YEG^+6VCPYbIA:bfY@1b57)\P68DN+(FSD;JFKRePgd]Qf@M
\>X)b[dL@XQ?JfZ@efDcZFU+)gbJgZfWH>BOD8I<VbF<TSBRL>,OL3=A/YR0OO[J
=T26OCF[\8U6)NKCE[NIODZ6BM>AR>03BI71G:e6:C3V12UQG?GL1AK-W5LP-^NQ
41W9Df9179ZV<0X6AW7J/<J3[>O5<&dDAP6\KOXL00J]^ZgH..K9ODJSSO4I0d59
#PM\E.[P?,E@e#Eg>]gROG<db>\I=:dVBI,VT<g,153D-WFT_1\Bee#T<LW234G>
G.?SZX(O+>^>cV]?D:\&F.Egf^_L/Gc:XQ?PgYN\M;1\YOC;7(RD8aXM&Q&?>g(/
=\B[U/HR@g65B:gbOfU-EAAHJ2;D\I?9AbDAN+5KA39SPVD:b^[[d^O(;<Vc13cL
3P08YgV.GS0C[F,06#:NRP7b]MJH6/U5\11<470>T)XF>;2ADb<be0[S9&@KVQeH
4gN,E_X3/64R(E=K8=GDAFUL]SZ3RL1YN_]/.#aI7:Q,<-;9(>T1(&a:DZ<=_]GJ
5LfeRVBU<<A,WD\5aS@,,91+/XV,)XUUXPARJ-L(<fX=]VDN1=YCDTG3QPWWS_/D
.TTCUG7?I1>@gg7-,<:]=Bd-W>2^E3WD+R1[2Z-7S8L6,O.9Aeg6H?;U;Ia.9DAY
&AIL2NB+c>)83ZZPC_E[=@KV5g9AcAN=b_(0dF4V0e,AKQ#2T_Lb^g8<e<KG.AP]
YFRFA<_@NV[8.]3c]Dd2g_O[S@L\C?bK(1/d0ZcQZ,A;U4dBM657&32Ff[U^HHeG
7MSJ3K8<8R:K1,KL=_dC_7JP9QR6Lc\9VWMWLbL3M&@R8OG0f1N+-1#K[#W6G;:+
Ne._gg/=^I/K#H(UG6Aa(H&^#_=7bI6)(1DD_B[T0NB+3)SXQZX[:K#D[][RW^?C
,C+@eW3b78Y7;cT5cXUUAWSC@+3e?(A5?TDX5W]#^a@NQE>+\XD=<TM1R1gDfWPB
;W_858addW<eLJeWT3-CaL,I--FB_/I5EegWb_L/#1JG29N^47JK2cR-PcDe&c?(
BR.@<A?(5e5(fPBW^RH9[cFfQVG3XDUEAHYfEHO//5QZYB5Q7]\S(Z,H;0&#V17M
Q+^QSXW;2gNWO8LgM0bI-2?+](=,#E9Ef6QH7C(J@)LXe/1TY/M-NZ)]3R@NR.?9
=,KZ;G_a[KS@b^LRCCED@ID/b906J+\Y1,-3f7V-PbQ?bS\4P[;:8&bCSP\aG9C4
XZO,.G+:V9^HM^(\PD?GLfN=A?XQL@[g3#b?e\_5]KBE[N=.F,R(@2T7@)SbFE2-
=<E7>404)@A_IbKIK09)R_BB\8-LAE=N_-#WCU:<UR.g<^OI:F;8g4/^E&5V)[06
S\60:d96S\N0:0[IQ@+[NU<MZ@JWV^BV#?bN7E1;@f2Q3E]59:60S#H4=XK?^4Vc
I_M;X3=#D\cg6\O83B4],O7=Z7/d#_7dAF7X)U[27V3DZ+KAg23?b=4\@;Fbe20?
_HYD(4=B2\DDFaQ4I&fYS-G^bQ:Mc=WKRU+W6g<=OI2PSf35R]04NCD\Y^_?3JER
72=;Udg<=\/O(H,5-/+)2Y:\_&BKU@XXT^+>]7B-Ae6V&;6F^G+GLeW@Pc)+JOF#
UdMGV2&gL8S5=#0^RB<:,=Y6>-[^+B9^eA4JL:__(f4eV2Q2?)@c);RO-],9cgD;
CX:_#N0gFJ>@6VNL.8a1eHUV1K)OO<LH+;Q+MMY+5:8a)2G28MLfI#;B,Ib2<\gK
9)e[;WP^>.gM.fU@^^V:KK6.M3,DE3@JZF:4?_eP:DM2@ZY-#_A,aG5IVJS(?[be
DbE#GFF+RMJ9>QJaVd48YSGC4-Z#T]+F_?SXWCf/)d;=Z?B0\DGZS.DY==B>=.SX
T&Y>Sf@)gf>eZG+9\(c9cT2YOFF7RVAIa,JT02Ra0LRU+=eBE3&c&QKeG7c0:(JR
_aVH(8N+=HG&3UTbddJ(W64O_D,^#TC7K+J=@V(S)Xe8,BW[3g600M83Zb[UEH/8
.>#Z[MIT7#Z7<&.8#MA2HCIO+EC3JLR.V^9X1F:+6_H,7=VY7BRgFgd4_JC50;8+
I0OYWXWM[7L5Bc+)4X0Sc=11eQD7YCgG<MK#5g8FIT>O(S?LG6@@Q;cZPTG\R>X9
/=/gQ6^FR=f6M?-B)/PUGeKL/##\ZQ;^X;3b.MY0;>RE0TV<.=;X1Yc3K)7,^2^C
KH=_L^PfMF.3A9,T18IOQc06-NVCGX,7YUK/CU4=f>N[_,,J8=U06Q,b6=3-=7ZH
J\.c#R4?Q/IH]JB>=4QQ)4\dQGJL(W4#^<H81V1V3F\N>MI]aPIN#RE0>E?ZY1;b
dUJWDFCLfRM1c8_F=AGEg;dD@[KFI9QSDO0H=^3U&KW37[C@@J1W0_H6e.@J]-PO
[W^FEQDB,U(2Z?CI\,OZ4<9=,SLNU@6eaH_OXe_W3-14aCV860058KBHZRW)&.>:
<Of][,LA.aP:/.Q2W<0FL-R44A>Q)4P>TEREd;=VP,573DBRbSPS/cQH/=(N_Z]Z
A:[CX?^[@=b/WeHPB6/E[e^@a(1[RVX6XbLcL7&KNa<D3ZLNBA?CX0[?^fW^4Xbe
J80]5;\Q6;]AFGg&>VFN,Q8J1WaIXU>QV/8aWc22N[feVLUY,>R,0)58<R9FT(EY
F-ELeOLKW<d:f8#eGf859@aE;=55CFaA[:X_F\KU,;[(8W3/DV^;FIM)MHX<+-SM
IME,N9+?a:-ge](1NZe5>8bF/)JL/)XJOC(5IVM8@8DeBM:=Y5-VOYEaR>6,X[)8
3Y73SJ&DdA1\[)]1ecRUGV=8Uc+#3aRAFMU^-;5>K(FCA1TH=BVW[/L_K.LUF:Yc
XT1TFfI5a=N6PJgMG+8NcOg/dEVBME3MG\D]+Ag&A))&A)&OYB<f(ZU5OVJYAUJW
R8&I:#4e>O)RNg/KNEC6P\X]6I_-OH_6\P8c857SEUC&VO@3M=CdT-<Lb^1<+e&C
]#fO#LPg(#)cgKDc-X+[Wd7Z91:+#NGZD8GPMcZ4TZ\V<1eg4T?f(bfMBT\BUbS^
VD-,S=dR7:F4[J1GgL8IQBS1TYP\=.P(C.7Q_a#N<5L]],]WB/1c(G7[0X;<d,>)
,.&XgOG#PdaD_\8@<,-AEILGK_MZTe)2^TU,ZCJc<,Q7?#<(FD7+V@7^SDA@3e8T
]Rd?OV4K45H]f/?8]RL7)77-d@9:#Hc;NS=CHaI<M70_U-Jc,E&L\/_^X:BSc8DG
Z;9bUTLDH+TR:4^3SHb0Sfa#Y2U#/;55#Dc&87fO<O.]9#TCZ=K>I9S2dd]fOJR8
a17baH679SWEa_D5\_[S3U2b[8I(+N,W<+OfSA,7_+AO5&caY<N?GD>0:2_H^T-G
]A,V>7#8/2+PY/e:-+f/54]U@V@]5&SS2d<&>YL@HOZ6J+O/\Rb0QE<CS+/N#6aH
&JQ1=3,JT@4RUJFc^0.VB,62de6fG02(AB^ec_6PD3BgLa]LPX@@VFWM<W:H1N:C
gI\SaP[-b1U(,C0.+SBF1c9]8H-Y2ZLeC7,+=M^&FG\V7eGTR0:Ve\^&]2[)]?/-
YZ@7dgd9@>,]f:VB9cR?_6[=N_2WP.WNZ.VdS[I)HW^Z3^0<5&-G\5Ha,70aY+93
_N@=:TgeaX[V-d<E_FbXfba[GaM#dWBQIXOP9ZR[ZAANYLD]VNU5,0H0;UA+03Wb
S)]C&&/Z+N)ObDZTX(U@YO?#H\WGeYJ>XRBP>JJU/0fd2G@ZM8eH4/fT39-I@?;V
&?HSU.ZECV]LfRf;Q,Y=0#=S_IBOCGSgQ+,1YgIbP)0Q>2[:3CXNX@+-GVLE&T;<
>L=8X#Y4GJR\4F,X2a;PF#]WcM>/<<e@BK9OZL6JFGA?@52f,2:EE?VM9KDT?Jbb
:UZAg=MQ=f:]R[15#5KC,DD+P2W\,<a^1>aCGNHg_G)FAYPYdX/cR9>9R\&eH\81
K&BbgZHg/_>H)B/H2HY(O[5IY6Y?72QCHC#TbQ2NWf]LI&+Qeg<0S6Oe<31IV&Y<
9dYZ+_P5efX>AOVf3dM6HM]4WMc1[;T\7DF?GA.d4De-?7(H\2NLGU_^P3YBL)]9
R9ZTKAgZOKJ>bY+Q/Qa6:)D[d]K;VNNb&#N3JI1D,RS4ZN//H7(^2=V5FASYCLJD
>B0Y79BABWTN=CY5:J<^N.9Sf^F#I[Id<DPW8MBF#5H<8DB16dBWcUYQA8]T&_A[
b=X86d7ga]YA9MKdH-^78CC8bEQA>11U-VT#e8VL<P)@PP#MBa3&@J+&dBW9BZ<F
7/CR9A7U_,&4DTFR,#--6PO2_?6\&7QaWXVPb]GT/6c+bM/H]De8L7R,bKMUU:J>
FFWF2AZ^L-9M.&])Db5:Kc0FMR)<HRFF,Z3GF1@(Z5UK(FQ&_PY]EB-.f8?g3J.8
Z8[O\4S+KFX\L-IVc&1SCH:0BeS\[68-_T&XB96<U-MdaHfT?.g[I6U><a85(VT#
/e)#KKMOb.UGD=I+@f5^Q5)\K(?PXf@2\\Jg)4Z9A8,)OV@Gg:NLFBC.ND._#>GG
JB>+Z2^)G.\34O>59EG6=]NJ2PQXUEZQ56JVDB9_6,)f3A84cM)RW6H2)Ff4M-F@
W=T)0bSIS;JIge9F<48N/ad^236Xfcg^&1FGcFcFPZdH;SBM;GN#[8M^6>QcUd-R
GZ_N]E](=;YRT64b3[DGa=NcRL=]Y@SX^dASdJ&;/L)].5)W^_:_(YgB(P,F1J4&
+U]7d5\PT9[IL_(;Y.<?1^Nc2$
`endprotected

// -----------------------------------------------------------------------------
`protected
Z&,^DKZE10:JEBIHXZ>/HD.5;(U.7.QEH?ZJ4D+=HRQC^PDb,f_C-);FW\,[ObI#
g++II8D3IN,J*$
`endprotected

//vcs_lic_vip_protect
  `protected
B]<YTbJf^<agT3?&0H)SGf@F5C3?2?HQ_\=TcO64DH/7RgN#5;S_6(=K>9]LecZe
.H8Jd5NIO_?4E1eTVg(C\YeaE#+R8:\/E;WU@&L#2U@a7bH\bT\?aKZA07EO^00<
<(aLef:ER=fUO1G:]K2YRZZHP_S>@O:843ZeaG3cKf^WO;49FC^QBHV<>HMGc8ED
&R)d-5J+;2#Mg_[R\@>L/>Ld-I5?E)]PV-VHgc]c>D09gU8g=X(<O\(E-KZA/]D+
_^/NELE&[SJL.A+e@f?c?+5D?J9+VgeeOMBQ<4fM&AZE78L2f=,F?9)(aL29#Z-b
a]O9,/eGGO^g90Fd46e_KPPC:>S7X.\@Ec]Pe)23R_NdQZf6b-ccH/?Ke<[#S4f]
dZAF)7@a^bS[cUNVfO@XV95\DI@&.a+R=A:@Z)^U\eD-;b&d74OHF;2FV;VgMc\:
WU]W=/PEB?JG,44OYg2ZQTQ(?01.JD#F1Pb5@IJb,4PRC+?.GbAX3Oe<:0HaOf>e
63L.IV=_c-c>#Bg/Z)BMcJL6)-9]Z6^b@ZC0>J&Y6#RRg5M9C]>eGUU>/Hg1QIQY
Pg][H-S3LYE=OZF@>a.d^CK_^#T17^3YaV/84RK=&X>a_@5WXQPP9bDTG)(?3KVV
N7eO;ebTf_;;d^)A=1bCDFa2GL=86WTJ0ZP9RO1[;+QQ&<f;:\4-(U7]1Pg[QLPb
9beTK?#J=)f];beGD-TF;L85@#-@GRcf#,Efd@7X0W?RM+Jf@QNXH.6<ge02T4#E
=<c=/c718eY?(P0-)fXH>7QM,)Je+03XRJ5<C&B,B6.?[N?8a9NQ;W\d,>7:WP5?
.\\H0@5C^-?Q^9+(?KH[AdOSKN+?GCcU;?:NB0+34B]4&5fW2[JPYQ+Za^-_+I;U
cMSc0GBPWL0YX23-T[4#f]MO7+\FBL6#^7N<GXY.,0X-RRW,RN\eN+G5Y;&JYc6M
W9#RF&)(Q<DBD+0XbQ,:RQ?UCGeKcZQ_gR4_0be_S=5YYdUe7BA.#H=RAfaQ:IgU
MH7]@T,QVM_gbG8N(0/2g[gO(/W\LWUX=UHNdN@L.C56cT4]J0+D13GM;KbfJ42/
W)\WQH[b0JE5Hd1cCM,@#N,9-<SdY<+^3]A],F?:SU@CGJU[Ne;&.7+<2..OT9/(
4MHAe8Z]:UEa@A<,_1H1EaR)DGAMT06SOBZ4IJ(EOSC,1:&57g5QGZPb=PZ/6VYR
P6\9QBg]W,X:UFP+MDOAFJOXK_Z=g>V+D/0Ve+_-P89J):Nc0(^Q[=HU\NH15XYI
/NGYV_?I#KX=8P/CB=#M3R7#]<CPHH,F-GAcMZfPQ-O_6W30[9\P?R3@(7gZcX\[
V7H80\gMf_/a:(fSJE>cNC1_d2I52>A(:[;182\5)A6gG<@DJH^0-\e?eKIUc+([
RS]3=g@SH)A=JRcG0O.F3Z7-KF,c<=>KH^\Oe]RPC\CMAg.Z8FHeOE^9I/b1K?#d
=TfC1?D7S[P>Y1eZ&^2fafPO33N06QY)@bF>LgQ<JaA-V;=U>RQ]aQM(@8g4=;S1
ULB2#UW=Y--#=9;9b-g0GE0d&T?LfOgD7]0cKP)NTQf9@L98F(&/N4Se3&C2;7#P
]gC]\=(VUW7,)QJ:TXD\HK\C8Rd-KdX#5+1d)J\W,W(e]4EO]OV#+F3).O,Ieba@
XbV64F65G\^G0&g:A#C2DecQ=]e\4+1gEJ]3IMSP:/6BfSDG:b;E^\)K<-N7W.69
GC-WRdE8:dL3g:_(cBAeg+5[>Wc/Q9(Jb_TM<VTXNT7^AQ/65^3.CJ/HF)W\0,f)
7YfdO3JFAJY33[fMPZC,eJIV95Nb9D6_^BA_KKfXR]_IE#RRE5A2gHRZ#HXQ,Bb5
?ZA>U=9Z4;#YB+R\6[Rf/[dBd@b4(KTEXY7JK)R2R@1=>#=,4#7HT[[5ZeH6,HgZ
N.UU]dPdKU8.#O^R9efZZ9?ac0VaX[E23U/#05UdEL76PV3AYH<H6B(5d+9_4F[F
>\Z#(GQ+fV1GT6@Q?(G6:cZ=KI89@]X7T;eg]_ed8a;V=&G;G5D5Z:R;YI#AB7^8
^\5[6(+R4XU@eW9TccbM<6a;/+X/fQ&^&J2<UCLe;Pd]6]:M.63K+eeE-G.:g+>7
3&?geSQ>B/888,DfCZILS.L4PRG6122]<Z83@2=ffT._<1?8O_Q8=1D<BfAXNM1,
.XQGJQBXC8H-L9((9KY/-&1\>2bKM?[fb_]O<[BD@=#QHN:)EVZaEW9\D;-C\Da8
F15)@]aH.E5QZ8e==);0678&[;];e3DYB,g643TfZR:F(#R03>.O]c;Gg3KZ+gRP
@R<A;E,Pf[.^9=48P?Ua^C=:#O+PdQfYG]1S?=GIb]OD=f@41:;]eK]+cT_.AS94
gM(Hf[L+Q0c:WV7,]W.P#,1NfBaC]N?@30M_&Zc6WeeW>Z6c&N^\_OOgXI+81C[=
7<IPOAM;W,7e#HNB:N@/T=9b9]L9]=Dde8]Y8&dL2:IL7&47LUbN_&dTSS(e&:/b
3@TbEL,JAU>>HJWc\4B\RIg2B?I.JJg#E1R/02e.5I7C&AFFD[>_S)G/L,1_4b^<
3O>@fg>MGPEM=ECXW:>cJ.=UEPe;HD7.=X=f0SJ&+\NBb3]K:Y-Ma.Md_4GKBc#0
C&KDe3b6dO3@]dYKR+F3>(2g(D;)@JN\8cM4+CV57_e[=,HN1)bB,]c.UK^=77@2
;^dFEOXKDR\Q#+O](<b_T]F2Y]UY=_cL(g>OSQ;@Q;#BGCHJHL7EJ<2IJW90WJ],
?2gZ?dA[6c);[^4;PfI0b3RWTPJRd2L;&BWCV49CcW;[>fcL_=58Ee\U??;+cQN]
],U?H<cN>@8_&:P3;@JWK,ZH8f>?[1d)BVQbP:K@aHdJ;\QI)E:2H=?S<8X/F-8:
UG2PZ7T>;7eB=G\LVSNgf>Q<Q.VU+e9fVDQ]Q^S2#6a36KDV+O7:O3<2SYe8L&ac
<f(33E_59c/He;Z0La^]^VN7H^[e:UIJ^8?g8(DEVNW3c^[-a)JA;QfeN^\,,\A9
V1D;;JL@[OK_<b]^5gYZ[QF:Q(@H-MdKRYM7JA^XgM>?ZK@FT&eUX_L39G,9=fGf
#<FWIG@CD?JBKH1IAO;J8Q7E]Dbb9-\JdX0&O5ZQ,9b?9J(:O1?#^X7ZJSca=-:M
6O;CV4G&>FX)Y\#V4V2f\/.6(eA-Qg9LJ/[?bW=RcW3S:9R@Ug;gVA5ZD/9KdH+<
Vd(.;GB3L+YXg:3H83Vac/,7:H.)62dW0=[T;gSY\8F5E-BX40@&O/<.AFYNE_1S
eVA[N9F-(.WN36_SfCOTG]753BP\<U;WT@1XMO)RT/gB85X<=CX8+7LN\Ee?a=<@
UacB6YVJ#=1@+/UUfY+>LZOQ7>F2?6FGVL6+(YUP)H1VO)_YBL[DH)0f=\I6&NKG
IG+1OT.P?7(2@@)CV>][-UCQ+L+;MLH(:54bY6O,g=/QabB_O1RXcV=Z#+C6\YM]
F^U4)RE6b0M5T]Zg:6T:a=,_Kg5U9>6(><8IDTa=K.TR?5M@U6092Q=XZ^7^894C
J+dE2QaTC0.0J;RH4f^f#E+>JQM,7a]RX)9H]I,7QFdT6bC9Q_@791C,>A#WKS.P
N_CPD0?_5810Y;)(E0a._aO6YBd9.E)fZUDN]7&IgaJP=@>EP-GU#QNA_e-@_JTK
R9RUa+Ff))33JJ/FEU9HG2K@0g:)+f28,J1=beG->+2YTVIWaUOZ(VFDFZPGK2>I
]cc>];aMZMPZIV:>@@UOB\?\e?A(=c>]WNPA;Qg+BQ4.2)cY;LCS[;>fV(8Ce/Tg
=UXXB/Z+SU0fa>8K^=>W:WB?aJBX?:\F97<cF-^Z:<8I,C6R3ZC/c;b6Z,;G#5HS
F;8Q:7RY6M/aD,d7A_a=P4(GAIZ4;4Q3-OR4CX+gbP.SM+WdK\_?KN&WJW(](H-2
N?I\-A7L2?D566R\P50WgC\.A@f^]=CDg@XLb#<b[E(-0@b]:,SaRI_:=DS;&e,T
-U&&]:cOf8L^U+G<=-=-&Jd?ARa;8[bH5.7DXTYB,0OXZK<)WXB?gXYY_AV,[[H]
MTQIRD?FT#1,3UA^KfLeA^YF.YYM7G+GQO#_S(93(ZO4I8>7QJ.c.bN>1&7QM[5C
]\&C.-W7T#O/)XN->0>K0H&dZfPL4VIBW1;U/0VER[06_cD)#>IJH@X^,P1Y);)^
-A+S2UE2K;F+W;>9TBaE+R5[gg^;(QLUN<dBGEB]_R(23H65CGfZd_:9L@CG?.O]
3NH8JCe#FS@\cZD3GP,LL>;WF)&F[_/I+R+Z@]^Qe?QE.I)XLK[e2Z0,4D8aV\ge
dWTN/>aZI:5=E#^L;P\fVTZ,2,UcF,2W-fG7B)F5-V79SA1(I845FIN,)_0=^IVf
^[#g?<TG6MLAILZb:[J(B_64cF0;-Zba+F(\])1]KP>KUPY;/Ne+Q_6=+71Y+T@&
e9Y6XcQ<[BQGQ>M-WZ?VKd6-FLX]=^ee1-L5+VLd=-8WDKTZA5\XGO,RAVO>eS9c
+fdfG29:1<91TQ&5>A7fG.Y>\AY5BK8EKF/AU>W/NDF7(COI6-DX82Y..P,2:H]@
GP/@C^4V]+Z-EC>89E>ZT&fa)\QB4>@J#=316V.EKBD^9-_FCH2?WEAS5FE-D#-)
E62Kge+\5+[;3/3G_cJV1G;6bL)PI23X#_&\)U6VV<4P3E[G)aV.:H[UM=a0YWIN
DfBB#K;D/,BM_DU=QR,]OF4,;,M.4G^aHE<Jc9?B&d:OeL(?@R9bSAWAB0eOX=2_
CZ)UV@MY0e@/KPN8CG=V+;MR_-8Q[a#MBV>1RJ,[D+HG:ZafH(K#b/>7D^-9QA)O
#^&?Yf?MNQg48)U3bP7AV-J)/,3INGHW=VLQ8eCU<6ec3:&7F0eJ8.51G3_<;[_#
C^g=5Od4CCY[C,Q8DKEGJ#:#K7@9H_\aZ]S/T8-B&_YEaQTa.;PQMPM=C5[La1J6
g.][bSC(X@KI=59<U)?a:4RU+RW+Q?M/^_U^S/b,9MAMNfBZefd/QKe@e&<TfQd^
6)-R]+-L==F]89=LM#_YYC3/d0DT_=/@)J;D3P3O4e;bT[[^EKQ4E=/RAJe?a[[;
f9?D?9g2O_@eSf<9^.B6I?U6V2^PHeF5UHfWcW8T&X2aL?Z:.H33UP9feJ<SBe3/
BNAS/<6U[_e5X/J0\T6<J1+LKZ?af\H5KO9;?J_DD:53ARMf9,);+JeT0:@8O<>_
?4B1feg<,bFQ8QHXS//cMNBI_+Mb1-#WafGX9Nc1dOE]\]Nb[]fXI]\d,00B:_BM
1?&TY\7E#=[U0RQ5SM-AfB,B4fK+F+.4P?_Y#:f,@.d0AfQ),#9OV6SLL1_:X4>Q
&@#YNB^O=.P_CPM<dS=V_OF8G.QYU]-H6#3d@Y?M7XIG2eNS?KC/NCMZ8-M#]=UR
,6U(N>?2RJD7WM77JS-#KG1VLZ5e5A#N7c.5O2_Bd&3_3.fdYJ_&:#QFI)^J@5ca
BNY:A>[cWbUQEY//=A/::f,DEC,#KBSU46T^XfSGF/QU2YB]QF6RMHXTY#=bY6bU
Cf1JZP>D+99,85VAU4(V3]JCC0[f.DE.]\,(30^G;(B2\1K&S)DIb?(AO68f\2VG
&/.QK<&.@F2HXJEAIY24?.gSa-=7TH)b_/NNZDcYALUX&V;_,fUP;TDg#]45=KL<
eNT\B]S12HS;[=?>?;GR_NaZU9)3>>aTf)ER\VJ8[2:UGa/Cb/L\\>VU#N+XRFe:
ebNZ9]6JR&?GKg5PJ=?./24NX,MM^d0Y[\L.7RNd#J?XUX6.KIIDX^1(T<TF>6LW
Ka,:;25PCT=I??77@O,QM2dX-&^?DQWX#ZUT:TA)I3JQg&9aYLI9K3<1#GGT?R-2
b6/ad,?<a6@(MQ2c?Z+[W7Y1TM^Y#fZX6I&=&NA;XSZ&7FHTBV+D<H8(3Z&C3;V@
7S:7LVI?g,NNU<a.?3?48M>W2fdg;S<R50U=;<S2Z=7NP-9>dT)HGc#HO5f79:LZ
@/XK6,2g\YX:2Ea4+3)O[363U6ZP6A#3IS)\#3NdCW=EZTDZ@3)^71=-WDL7&be]
.e:aH-c8W0=+6Q7.VbSaZ05V&OL3R4b:aBd:3W_?-4F=f6Q1d4;UR6NZd5CW,d]+
T67eT&@L_J.QUf#@KH#K3O)_?B]cH#^NfD)EVHMVSM;=)ROSH)f[geZbd(M0.DMe
=GO&=1b@M\VfK<e.DR1WR-)TZ;B,A&-#=eQ;1DB=dC1I>Cf>T;cc\fQSc-I:FS]5
5_:[6S6(J_P2I_,?.Jc#XF_)S+ZF;A^V&@2RNGcWe?=<>4Q:Ue/LNDN#W.?6;/I9
1V=EE1#BKcWV29K,d^,+LY47\=b;GTG\KZ1&?XJ&ZLQ7-DZ=9@S0X0dHGT+NBe[6
51LV#]VD5+75KF)Pe>=B=GS?:g]K.fFBTQ]R#63g)H;0CaBZfbV;P:X#3-)TG3D4
[&J2DP>5V7bb2/dfT58LH-6DZQZV0W#Ag78,#5D1S3F-\c?\gNE?@J=9A[OSE0Wc
3=f1B0HZ)_7HPZ022LH3L?-;^3ANae_bXcgW6?UZgBdG(3.+@Q;:1=VS?MMQ6]80
]^CC5aDDM.F_GB@cCIZ^VTCNIJ/DF88SM)-<3@X.4;-Sd::XIFWUO9d->eJd,V6e
68\JKb:@E>ZR1D8f#,\>GZIbEBN8-e(#Gb)&QHSHcY(CIGB^;C(B-:[)M._^,e(V
8;^GL[J7#>^dcEB:^>DNWF?GHB4O#8EZ#O,-R[NE/>T.K&I&/a=4LZ8QCg46(Yg,
gRT_aYTI]0<d./Ld9W?b#7b/W/YR+IS+?/5W3-T?bC\cVT6a=?#24f^WD\@G[C-]
>a_LdX5J^J@HBZ1#UX?\\f1IMgB3__3&1e30JD6JNBR.T0L12MT\+BB-Kg@:Z4R?
_e2G1]8a&.g<<c7_U0ICON2L?V^SDbT3REHGgLA\g8^aUR3\Ud[>&5-FI_QA#)F.
O&E-&IG/B@L\B):g8=UCc;cZN;[A/83_\,Qb9RfE,:MD,C9eZ@QYUfbb5D_B;:FM
b_HQCf^=S^-=LFb(M1X>(&DG1a7Q,:\4FHD3,;HV7;,58fXVFX&g[:I-DS;LXJUV
3/;W-7VTb/+-VYg1_<F_BIeZ2AN^&FILVa]C(=eF;)KSbR6]HUVLcSc:(UX9/FKG
dUF^e3O.d;\F4AWOPQ()b-H)?/=\EEVfL3UJ;Q-Gbg-;@TUg@fZ&A;;d67T?b_[E
H@U&1LPY0g?H2:cMP<-S>4WL2@VQO\+5500@1]M5X=E9AR8C+gP,a[J;eCR43C&g
ZELEN0A&FP-(1O9e5YM059cG+IJPU<ed:M.A^);\S/JXOd];NLQR<ATDSW_N^=3N
_a+]/ZKVcE^3N0;Ga+80HD4<YL)V5f>=Kb#2dg/5f#C^Gf6\[Gg([?4TN=4AMg[4
BWFeM.\6WIG#c-\:;N5e^dS>e:W(gBU3aC[&R@aBc&\aU&J^GDH)&9e[M+?51D1V
BAS@aW87c2=C,C9#YPdDa[YU18VR201&.I4@48OXV#C<IH9^#8aaFbJdX&H5_IN@
b_]Z_2+IP7Y\=^g5==Z1&QZ?e1Ea#]C,+#44P6XGD3\2gP?@0^.-aF:bHA.3<GVT
^R0d,edd8;L8,4I,c1),/a1)7;U2Z1O5fP\U#a^SKd@;:g-fa/MW>3_4,A:QOG54
K>f-<c#eU/4SgI91(&>_P^cUJ_a;)U>d5NM/3Yd:BPNQCD[M/X&<eH1;LY84)4/F
<T)^Q>f=AFUOg7F;f4I<G_YJI.[A_TR6AfG6Fa;\8a-]UDFbd_;/19_FLAYY-\YI
ULSNQ\/=D;EMCZ(WJQYQ(e/_FHL_JT)P:B2ZFU-\;?JYXKZ8PXA4=8K^21bU[_LG
#/&F/YK7=WN&-Fa<cX>UYBMY72SgTMNUG=.5^,RP0bL,aPD0d9<E+XY.713G:>MV
70W>AL<V8A/(E6H1@K?)T1eRCD5/7H#,G]G@b-bZES2CTX4^\051_[XMg-Z]5L\^
ITS9gCVA7^9.,S[6H(7JdW1E8,K?YH1S0;M+8a=c>g^,;+4V]I^VbD]_V@K-@PRE
(f1TZaD==7V4GOTT1ES^FM^/>69A[5+Ye\?C5c&1_\=#YAR<E3]d]]TJETEDSV0=
?;VS<+7B;@[gge7YUH5&,@DXO@<7][(>(532AMaA];WP:U#,74X[<DBHF/cQaK.J
Y>P#>E1R?/Tg7K)bUN(^b7BINGg\3:Q/TT[\;@0S[RAf+U\1.aFYK(ZK;0I[G8:N
X4A,,.GC.[+(f-BY>;4<#D(>_d68bXOM-Cf9C<eU+^_6f,9-9.e=G>d,[-3)I.#[
cAG<(MUMRF^YH(V==eR>.QO&dJ>8?<IZ<\a3]>b&0c.[c&dFfWEBBUfU^(I-@7b)
g+(6IV]5[O@C5R/TgG6-[-9f?9MS\=g7MN0b3WQb_6^UTgfA@<AaG=dVdSa-^1[+
90T(7+:NC\>Q:YN9IfX6G8#:R_:[UPR\d>I.b])=P5:U5gNXFS,T)FL.Qd_3ac<c
DDX9/]W0#HDfS9MW634<:@H8WL@<2\VDHQ<L9MP\8-,U7b?,#AeQ8O)Eb&g>-1&P
\FcKJ,(J/gR:[H=fUP]Y=/-U&8]<1M\A;)]2:6L0(1BO@H^Ve_OF:L/9DfLP9V^c
b^GGYbd??+.aMdPc<=I[IBDKI_/XeHTYNW?:HW>2TL0Fd?V]KO4/?0JC&BfJ9Se:
Y8S]5fZ(c==RLY8+5Q<+W>:Xcc1QFBN?3d1HLP@6YP-TdY@N/9QHe)UYYHM3:Z7(
FKO3[daO.@Aa]]]<)?fX1aXeNOQJ1Oe0K5OH,[>+6E<Ba^?/8de:Y&8P@f];Q,1B
(ZIa]&EQfGGfd.I&E)B<]XH=f0Vf7CG_#T;dDSH5bC.]:[,STJ@W2g6?9+F;=b3(
FC(V;g\UKLG4.94V_99b=^FE.aEWHLGI8NGP[,#I>\.a7Xb&>#ALWDQ@a8VJ=F4W
&G\+Y5X9BeKObKS9dJQ_D^(D&,CO:IM_;ScQIS@.G-EcUNP^BLdOQ\aX]E\()QNE
F0,0KAF(M6JO>],c\2O0WN?>-X5JcgHfFMY&RLLd7.8YJ-cMJKg\F7VU#(]FZKF8
,MX3Ge824e(e&LOef/4;:Y.,0bBSZ-I9F)AVG:BLSd([5JHU-7YgBA-BUGZ<[X9C
#20R8.E[PN8Q+gc#[bKZV><VUF]L8V:E^;E>]Ade-^BP4a(LZJG.RSG^.V:-1G#S
.2#N52EFXO=8V\W;C;fS[S4CELMYdL83V;K<O56/2b_5a&/ZCSX9Fb+70eW18(3:
>2XX484)U?9/Z#03WZbR0>GD/ZZ=BYe)J>TA<][2\/^(<Oc=af_Xa<CFRe4MT-2D
1^B(T.<aJ11:<X>M7LRU47=E)a3W2#\WF>&@JaZQd>:6L(Ac@X?Ab86a@WAc8Lb^
5?1](fGeg]MO<FG@Z5aeU2UTN8H3/a#;Y3D=WES[3F^YK&58XBNOMLOK<AQ?3,>,
NbZ-,./(FN]-)X3BZLG[UPGMPdeTdgMEIB&9O1&-+=?JYCd0IUGPIe5?1=[^X,F1
RMPJ3ZOU+d.g6=@-IUcE?B5d:O<AHMT.H?GVU6Xe3e[X<35W^(cO=Y2PMZ&&CF6a
TVF/AF39dB&)<<2^TPMW;Fg_dX=EA=:7>9-AP9=>BQ:VP\6,fVcE1.H=U=6Edg&9
(^&)_g42b[62YN31-=H(CJ]><GY@b??GY@3#Y#JV.(g);D6PB/>L,O761<C>S-@&
EH3I@DGaPf23BE9MG-\H.YP7+RK,H[Y1T7+8.]YY^@)O^]K:,?:N2Z<1B)YK^?8U
::>K6c(W3.gPB^;#7L7KV&c#)fZc[)Dg)#]>J??d./3-=L\ODB74X4S=3,?cU]_K
H<O-gfJZWf>J]A8-W9DAXXSQ.4Ya93fYA?dXX=(A+[U(FV&EX3JK8^5HVPIIg2b-
2^+g1ML4Ca#LSXQE+CXH2SESQQaEeOPa9e,C);X[,A612fb<:g:AC)-d@<S@YW.&
6S^4e\BX-_Q@K;X]Afe7FfFL:&KB;0Lc]3K\0ce8FcBYb>2/SD^\2+/FcEP/8/.<
=&2VAVD+)BM#>QA0J?E>^=5IcgdQR0UJ#UNV8@IP??=d^\W:97>G)HN>>X7-E[D.
55/&B<\GgUJE#CTZG(9:3X)V[@V=/DLU0SCgVSOe>4<Wf1C6H83[Z&S\gLE2aPdL
2GY=?6;-Ig7#XeSU231=DB:[N\?L-PQMdC4FT8XLMHLQQSQdGF#<N<K12WND>]Z8
@N44PN-39O@a57C@+S30AMb,XB7:M.Y&K)4.LKV.@8(aGS95[J?GFN@VdQ>G=a:A
\N;IQZ?S_0]>e_0+]8[=#KaHLQ\\6Q1T;]6cAWOgP[0.RS<MK15SbK_b+^R:?I.3
C;LO:g&/7_7SWc(W5_(9<[#7UfP/L[KH@&dV(/:KS+g[Z5AgU1BHG.>LH+N;IR+D
M\(8A;K,KS\HM-UQL\)YGR22/2<3HX.DBOHS3c>OD)g.(fX>/I8XL\@,fa#d6ESD
H6CS;MN@C1OM3M]?JX7,[:R#-4E1]3)>Ed+Z;.>ZN8ca<aTYT];QfN7MO0XM)Mf4
cDUO3W]55T=X4Q_[6)eL/b85K0W8]Z#,CgS;C5VW@N1cW:&6?V6c74;Rbdd^G(d:
YO.+e8DB..ZEAILZ_fL>B9dN<HbJ:>f.OESECNX:\He4AU1g^[OD,0dg<7?Q-M8b
NQM\.^79gG3:FQ6&g/:))SeE6HYW^Za(SbXS0E)#\<YMab]\b,SZK4:8KGSTIMUZ
fX3-M>P13K1&W,F/:\[8cQ-0NT3V6DU28g7GIJYE3H]@aM:a=c=0DP<gY1Xf.&]>
P+?G#ee/P>I]\X3>g^O.JF(aaA6(<ACVcJ?:;6Ad\8L]b:YU(_7,[\>.GPI]:HFB
.U_g6c5V]g)aY<AMe+O^=J?QgdPMAN3]/.JTSU_aPTG-Q.J]AYg8,1VL<<=M;<C[
Z+F9+A#+@dMLF4B+b&@>J<D]eB82c9Y<_e]B88/33@Y3]e.^A5K@YNZafH#Z/U@;
I_CNBY^BDVR#?.IQ=YT,c.fZ16QDYT3/0\?;)E0)&UfUX[@Dg[d5FY\B0IBGe]A7
U6,Pg>=Z/LBGE[d36=SfdBc;)?R2&@?9>EFVP@^87e-Mg;Gg+R@K6LA23O_fZC-8
/ASQ@E@ROWb2OG3ZMb0[:aOOYI)&c3IZ2OD<Ce)5-.Ra85c+P)bW]J3gEQ?Td^LC
NTRU,Lg[F?D^K&X6B?212V-?M^C86dRKL.7YZVdV&NG+GRZacJ6O#HRaM;##Ue_;
K-V?IQf=c;NIF796/XU,CKc?X\c@Td<)4C2@;TLNa[6GeG2A@2WU&&ZOI)Ig5bGS
U+.Z1\A/dd&V0VJg-/;A;[;U&eM-WL@fPAPBTf/;=ACAGE3)+15d_f[>-T4@EMM/
7#g/e_:TJDBLZAC-/Dd&///QRA5/#U#F.I8PX)SAD&Z3.7K9Wa#(&_>,99#LMQ,N
D&53d?fX:cc9WDeS(f/T)A<?==I?aZbRXag&fCe^>289#K=d@>e[&&-fMHF#4JO-
<2\+:edD^O85&7d6[KGU7RZO[G>ATX3N&6WR1L=cVBbP\_RPdRSf3g<g36(=7NJ3
<gQ/@YXH0^[9f<=#W7I;SH#RE8>gM@a(]QLHR7.?.,L7V8C\.-1K8_2L&71P2N67
P\:_,ISYag7aR<WS\AOE/<EA[8-/F55,#DZ_<^\^.^1]7]B?56?Q[Z:@65(:M]26
MEeE>/+4/J?K^b>#XM\K6Tb(8U@]EJR.>GeN_c)SK;4OI@3D>TQ[P4PW,\SfNY><
OHT^S2W.dNd-R:^ZBd=db2@2\?YGEF)>Afd\d.D;F\+VOdS4@L2FG:c=&X+X8U>:
?eZ1X17>OO(MgS_6Ic#g=BFC9_Y1[IV)J2.e+3ea]5GV=7bTb5d(T1TS^bFHCg3H
7]H1Q#,G7Oc[<3\(+Q]0^7CVN-^1^WZQE+:_ZEY,E[R1S^RA(<RJZW8Z1F,eVfU7
1G;dXTXYY^G]RQ-2^CE^K&YOH_85PT,)/?9V:JZBD;;Tad)7@#-ZUB?N9DY.NEAD
5]6PR7&eX1@OZMV1<g8e^1D#6E^8>,MR>a:TIC5:03W4A697>3JDc(Ud35,L1#+>
c9=>7Z7H=>HRKcDD>)6HBK.Gc=2IZT_]#<M6?G1A/^fKY#Pa2=,+-8=LWZ&Y(Q.e
(3+QCZ.V:J63)RC/U,F[U0Ab,J1AFDM@T3WWWK&EF\XA#>PV=,7ZFC<03M>/Ia@H
b+GdK\T)R=;@HZ\dfIfY++8^K4?31^Bg,bKJJ_g&H_=D.&;T2GM0,D8)J-DD1-4^
KL^JAL,\HC8R+N6f4K+P>RdZCNd[B1e6O-gJ61-^^K^6SO&38#NV<S?YB9[>L(ab
]:Gb/d.9f=g,M0R7IDA(OV+GaZM++ERW>-7,L#,fO,7.<[LP?.([W9[CTG=L2-R\
dO^&?V^\J\@](X72K\d[RT0O)6g]GW5/GCTHXG;g>(7]ag&R=(Ze+>(R\R=9\3<2
D)P=+32d[SB2.ITR/5^U;cKF5dH-D<FT,F48TEY_U=A+&>L-2M6/g<CE5X;1?HdF
?0OPI[H1&5dS(a)DeO5&6AZ:S?bI_KZK6XCK=,X?Ma]E&6WBf4_c@eg@F_He2\]_
_+)-5&ZL/[8M-;I)[M7^-T.L4,(9;Q;/6-5WZOWOVY4<WO8-1&:DDA5F^(A\/ICD
UNP6]6OY,SJ4C[@(QR0I_;=[TPLJ-E3,QaQ=0)WLb<9D5Df@fR?aJ,cg.L/_LZ>?
PEL.XD(N/+1PGW2J1?3<U1aMb2T<(WK2,d=0=PCH;^YUD?7W\GMNcSP:;DXSK_gV
.5VFF)A><Q[-edf^5R@M5YB<<aZ#=<#3b)Q<K.XF8eA_3U,]DaLEK>ICLOa.4e:@
L,X_FQe<0Y4[6]\@UC(7?4/BJ\Z@N+?[Tg1LXYO<PGGA5=JU&JF>;0.Cg4g^\fX#
&R\Rd2M5//VF^0TZ\ROXN\CX)GG(7:cEU;Q\6M:VMJIgM]GDRd\-MUHST[&SS1&T
\5g,3M_/@-_8D^c-UU.HXbIW\XD+:PGDOf)N\fEd2C488:QP&N9E2+RSPGf2;eR;
6IE2BXL2fb+GT(gLVGeKH9N0N\-[OEfdcXfU_[^8VKT+2];N]W._b@L6WfHeYgB1
Q-I9F<ZcfE<:VO5H@BK=(J]L^3GZ),cd4TS=;2[E8?X;?]ecC9X\0f2@=cbYcWP:
@Qec1dM7cSf#e3Z.AOS<ME2V5,f[8)^8c@IBW?+VU_AVB608)b,2#?@I7)BZZYQO
.]7A2LEYHf(EE:\;)IgGe1:O3F:1H_SH^/aM34eA5;CF/..\WDMF=b8EbeN04L\N
+Q24D/.=[PbR#+4][YdAA858PE^N(<FOQ>AP.614&MF69dX[H75XKOfd4JUR85e2
A2GbE;AD[5R>FE/UW^aDKe6Rg9U;3IRBC^MObY8-JI5,bdf#5LdY5TPD39IP8J10
:BeLL;RUY[#/g8g>A?.XG<#baL>gLaV>7\Y_TMK)DWBQ]WC1c(G=YGCDY[cR;N1:
NA>2E;U#FWR#9(:SG-.fU_Lf@LSRI>/>,NedXY5BcV/VYCJ1+[I=c6CO73B;/NZS
1>Ac.,.c>ISfcE0G=U9.eI]#bD=KO-KLEG;LR:Ua?R^^T7KeN;UgZEMA4?Y3@]7J
X.54&\ce@\:U)1OUI5&7K5fT,Q,[gf7JL30g/>8,.AL=VLfJLW1G.Gb]LRPA@4dT
-gdFM-^R&Fe^3=DC=&#KN\fE]Rce[,W6Ec,X/2)6EM@8F;2(MeVA>.DD\N3RFDdJ
G2XeM<bAfa^9&AH2/)>8]AKY7.SI1O[dPIgBV:I3b>9S+6UW=YGVHc08)X(#C1JU
NCK_BRg;)-I>H?A)TWNYE+DQP9d@9P8Z(4U#E5;;;R[9LH(Ab[PBY@A8W5(LVT0#
PSP^B]e[d#M^+N=VO89SIB#RXG5QF<JF:=<cdIS>/^#QcSd9&IU_2SQ(aWV725;=
/1?V^F+PZEC?X[[)FbM\<3&ERPaB]J^PP]AQ1UL(E>e)QQ_3K&-8bETU0dNTP7_X
AF9[&P)#EX<FSCc+8>Naa4UJ)bM=EM#T?cGZ=dR35O@@-6#,0,>1DBAL2@#BKg&C
\PD@(QOT9\,QGOK>a>]<1-YD=>VH4E@I;A:Dg&)D]0CQXAbK\<CJ2G[D<-55@8@>
M+a61)B2g#c-cWP,>_L[ZP3-b-N=^KU+8Tc-X&2#3CfgP;?;-O+^c@0D2U#6Z60;
&>=Gc#^4b2(NXc]F_IKd@;eR22gg/:N];[=7+ad(;6&RB]C.dL3Ba()1+cY=8Sg<
2CCKTOH#V@-V^c^\0#]L6_CcM],82_6bF4ZQC)DH8<FFM(H9MV,H8GfRRcD(/S+[
&A=HP0>cPK<P:CK^ab^FF^:)NY16@X:B07-a@YJ3K6C/H60=.&&V)JGDC6c@ceR<
<&<+636Y&#7I2L?;O--6@:XcNg;QaTT[JL.KH3_fP-\C8Z@AK<C8]c8AX+V<2L9]
)ZZRZ[8.(I)<^YMg[H1,9)MfcLgEVT;<B)-7b](8X^VU/[[&+>H1)P[@Jcgb2NbB
HF4[#0[+d.J[2=NeEE&3RB8eX<1?HS5(ScVFXE-\??O&X^T0efE;\IM,5[.1QAZ-
BAIJ&7d&(ceg(eFO1\:MPVE,KbX:N?TBIcA9If.OU0?,Z&J8Q.C(d[T[VK)LZW<\
+?3K+[(RRd341P^OA81)S<[55<;gK7=)YdZb7QACDA[4Z1)+LBVFOOaS,T1:;IRE
Qcf&?e]4-LA_a1@/c]aL0C<Ye_g59=0?CQfS]#XL#0Kd1R;()J:/c(>L]0O8;a3U
6D>M[]KC<fK3-ObG:Tdg)P2QP^4a1>17>3ISZ9KVYSLd=>(0D#;>QC.558:4K,LA
=0Od(]aTL,aZVUT#)]Kg@IeF</7ZJN<&C_54G6@U.?YXFD;PMd8eb^O)ESbe4@C@
JH5>e)YFI8W7-174g<(VAZfOZgNAZ9Rf(Y0K_gFIY1F4.UUT>4((YfEH7MQQ-R#4
CV__4L+6)S#ZT;TE<//?A98X3X;]CI@9J3K/^dS=/>dg;JF3(2&0?2d_,-A(PTLY
KC&611=BcZ/]+6<7d(</]8YKW(Y3CN>U)S?7HWd5f:8Y_]VgZI4[baAWG3(.]00M
Q&+7-aZY<XM[e_:ZQD<4905,\FRJC:@AP#dW?a.6>]M;/G(/Q/gQEG,I=L0Y5Q4W
(YK4SP=Qe.VHY:KFAfJN6Z3][L_NX+)@7XF_S#D4?ZJ;O]H4&UU?M/T>XdW::<^Y
a=P(OJDY<8G;9.8V=aX7=1@^DY2.GR7;T-HN[cX,b;MXNO=]>;-&(O?YATc>09SN
4b(KDB9c0<XA7ZAPI9SU+c7PS,JK90[)7^GZOAacU(<G>bCf).V7MG&5TLZK7&5.
\CO7e6bB(&EA4I=[2RePISd>JSUOffZE?NJ4/EOcc)@.gY([VUL47aIa(bYUYP@O
9#/g#K(WL;GR9V=T:^RS^3_eB?LYN54Mc[2=O\APY9B;fEdb:[KC8e[fSS^bNU@P
[4[L]\#A_SFB_,3Z]45,>O9^M#0^4#5MKb\D?L+6Jg:@5Dfa<_5a^4Rd#UFcfccR
H8?+566.-3EdQ3X>F4PEL#F/8=+5ES^0d77f68,-WcU0ER_1\UG(Hdb0O[Ab#Z3I
6SO.=A8D-:@PFU-M]9K:a\=<KT=.:0[D-A8A;QFNgVJ[<S1OEEH]5C:QNBZQ8>>\
L9Qcd7Be0^\MR#N[+D6CA.e;--#/FSIG6/SKQcP+.[\@@01/X\.Z>J_Fb-P9]9L>
01eBBNcgA.Cg5PYFfXF_;Z_YQBJY+>P>.^]-0Jf83Z^921^Z?00VS3H\Vb<8@IZe
Y(#38Aa8XHZPCIFXZ]N8]@&RJ9+GNcfb+@f(Q3T5&F/H\-3J2#@=,cc2abdU,8O)
_bEB&J94XX)^K=4T>1^;J_eQc_SO^V8>MV9G_T][NcQE?&5=b?+a_>GRV&_#_e@,
.Cd=UG0;XL5K/>)@Hf?:,F]3&a9P[+Q,(25&):(OIE\6P5P6B]aITe+dBDdZTC-R
):FI,ReQ>I<VG=<T#E@P+;P#BNS\7>.?P5g;:[bgU](+MT2C;Dd^_)#[J@BY2&X=
,f18S7=KSgHI<FEXfL-/@LLD[?@+bDbg4CH6.[Ya)H3b^NG/g0\N/+C;c,2d\e/9
28T9V^5;fg922O=KKEbTL(1C/IgC28ZTdFbXb3T4IV5)e^Bbg?BO@EHX2.ZHJBOU
([-MHF(4a>IWL_70K_gff,8IS^C,+P+,g0J,9C-(,-C/S7DM^K&?d@QG?cXF,;eC
7dCR]92_=/6FYgOdGC8^AMI?\<8;c[S^f;(#6e(SFUde1ET815T)O9,\3/G4K[<I
CAAYKXM-\M>@)-g??XGFM.=#-9N]b16/2+AOb\]:g671>;QIdNdV.N..?^77K.^(
eKf[V^2>J/XO7ER0)E1eG^FB;;.N+c46cWYW#GW^aW<g&Se^a6T:;0\OP>=f@]8N
DXTBVe:OU/?a00>:3bJEa;R#OdX[<e/KO9Y=J&g-;?g^R_0fgc_UIFIZ,RIG?\JM
Eg1Bf9V@C4E7M2#0UD<#B(66-)WVg5]#L602,c_;QO)E&FLc,3_L5bC<]F7T4(/#
GB&2Pc0^=?Ec(LE7#H2I=.J>DL/+=fKDc(FN3&\D,#GOVB]YS^G[^/<?D\3gL;?)
H<3+QW,ZM<aE85;@[0Aefd>d+0;WW(PcR\@.J^X7BEU?PJD8RCGCBCRMZ3e=_&U(
6ZKF4@0).9<BW(=N=P<\_g&>TRfF4#.&6>CR5QWX=S6V=(?2Y[)FHP:(E:(;)GgZ
UN4X=d]D&G9MEG>O9:GTKX0DR8P--P1EHMWffb+JN1X.NNb=?)IHW)/C045YZe2V
C]_NJ^^MbBP1MR7IabD9L/b12-Q-SF7T=7gF();.0g5>=/,:9LB)-5C2X8Ua_M9G
L7Q5C<aTe<=\MdFJ=&[J/AS2<Sb]1,GAe37S0OME@,UDR@(^?B@;H=&#\>7#eBTK
6FU7T(d:\U6gIb<=Q^9]5P:Gd&:Cc0?<5H#<RF9NI:NDYN@&TW.G#XCPZAfg@O@@
7bHd6PZcC,f2?D89:?9P7b?I7_XKVQ6d@>P2aOQaD#<@V_@HE@4.6,ZX\)B2-?]b
AdL<E)cBY[D9)FZ@XQ10>C@N0GG=8T+QFaIDOFP_?ST/N0;5J(E0R;NLN/DeHJM_
-?8F\X3Bf31&[]b^B.[./[_R\.BK1#bgg-YF\CABa#SacbFcdI2B-#1Y2?V8VEP&
,O2P:V0(\/H&)WGI:\MMK<90;6f&PA-JL<32fZ^(UZ3K_QEAQV=e9<9VE6[K3DTY
c/&R9(M824F_H?cDN/5=8gU;3]LGIVfM<O2=?QW5bAW)=d51GfLJPO,(.2K-_@AG
?OfOEJBJOJb?gW@&9,dUa6?JfC+Q45NJ47X,V))QR+d8dOe2L(Z1(EDTPWA>39KM
Z,I.Ec30/5(]FONM0BUG\2:G&):I_+E;B@9-[Ja/H_Z#[#ePT#X>aKP@H4Jf8IFD
WDOEGg6B;&fd/=fG]]T082IG)I9JLe<ABW2SIa+3HZZTNM#M0AdHT4bT_2\F[c.5
:@=MG4<:1L\B_P(5-:>R+]UNQP3<\M0dJ&/W3YCS\eHHA=>X;51Pe]J@@dVNf5-^
^CC5.1I#+CR\@c4O^--G8S.ac4G,\[XE234e7(M]]P6OKMSSRdYbAUH_E;K<8W,T
E_a0,0IM9Ub;aRY+.D5DKH1+WIX[V[\NO(_f9PD>C+-N+/.3(]9;X3SS:05(Oga+
L9.=4.:b42]aWTJ&W,K#+U&-077LR3X\3^#X^FMYZMa5[^Y\QK:_=^7H9E0EME2F
ea9g^6L@6N+4/T(8KJVIOb9>75KQ.(XZLVd9+f=?\^5G>+ZIIX50bQ2gfA[b6^,5
VF8&S,8SPR\]V,(QNJ.\8X&Da-B)<-^,+,K<PO?Q=6@V:P^5O>,<2X9CSO.\-T1A
AY^:2<C4.V/GS#YRP/81@dcb+d&XV@;1G=J_OBM:P=gcSC0&.aX,.]aE;]M<.:T?
DP@)NUfJHWTE17C2f9+.5EY@N):BDB1f\ZX,ZC)Ud[J<I&1Q1If9W5^cPQ)#ZO-2
PUFHBWEaGM:>JKO^cg4P:?1GD0MIOL6gFA1aCc1ETO53ZCHSYZTP/L/.L&[-Z,U.
87LN[J+UfYe;@82G_e3ZI.CNbdN8dAYVH.b]<55&#]6RAWEaCF4J<_)^?<<NbA3,
AZ]?T3_UGOJ0Z6W.9>NaINa.E:46bG1@X.-W,QPFcLbTS[.=/SKOf:T[I6>8Gb_[
O8KQ_S4\14YQ;RP\Be@\&6]Na4FcQIU.e2RbH?G2K5:P[BeQQ+XT]gYDAHQfUF1^
FWA0>+WQAR,>BO/#X\[e1BH@GgAX/Y0;3W<0.Yc>Z>XM_ZYeXJ;_D0BOPEIS82ML
^GFa4V0^&>J3cdObbM7R5D2I1c_1d<M((RQS?JaT^Y@3F(7CMIg.5=UN[<0QK+2S
GbQ,c/\.N+YU6OCc2:_Y;PX0cQH0L1SPL9=G=d<OM4Vd6W3S9V-I^g[G/Nc3E(91
\0-LJ1bIB8.P9M8_U3]BBL(fL_;\cO,RW(6b5D&=5K[2Oeb=I+gB8[G78)4B38+Z
3/#U155A.VQ>T0YX_K1gA\^@>Z\Q1a-\=(Df(B_D/)L.60L3]ID]Gg57eeFCK_5#
9KN-A4#:^+/#>]C/V^F1d@OIc6L+60JVS)=0<=&6I9Y[YAJ_dZ-KaABLH1;KY>O+
>2)[3&2_HA3-JAJU^)L+fNCT/=)9<?fP71]R/(>49(CcB>;eQ;IS,Yf76#CVg9C5
>/d)-+#75T56d9LX#ae@CJ7a:1OW7Le[g@eFfVWLPbM1D41D)G=U)\Y<+?QG2b^D
^JUP).43&:TcU@9[ee_QFbK0DX\4</F4:V,[LP+X\;b^6U5@g20@P)+O;7AU^Y=3
AS/RC1:.3KU6D_ASfTWH5IR=/3A,aUN0CWC\Q6\EY5L:DdS\6)fIX=K=9#J/ECRA
NQP\bMOFX42MDUVR)&5Y1ALe<.Y7@_^FQ<1dM-8C38Yd6/-@2egEAI\g8[ST-VeN
<F^A@P>TRV)/1UKM2^:M,eCEYNb&XTW5\.>B#T=B4Y-,NEBI=V5#K_8@c#\B1EdQ
fC.2_#a7YeNe^8,f,3M.M19fVY:;_\f[RG3/\7V<(;=BdXT/9bZD3=4(TEA)_J^E
859SIYV<J6a[?:W2FG/B#DY^7,OH1-Z^ZE,(.94d,C,/_+&^:X6\.PJ;5RTFT7Ue
#SD\U13XS=,JMc_SY^CE94_NH4R9.ec@3=ZMI5@>gMBVDe1W]Y;:aRcJ#fPOD:[e
_MT3X:#8.L9gg0N/ebRS<O+2/M18XCW>QF>Q78;.\-gSJ5R\?9@G7,OE1g>8C^d=
)A?[b.9V-1_O6\G[Y#c-Wb0F,>H.7IA0[KE1R:F,\>^Ca;fWTT[Sg&F^5&.e6TbO
B+\PD#4RD?-/1<A#ZF/;]ULXSFaY)AfN?OHEFODU#+>R/;Q#:TT+6M]@DL0XF5[1
+O<:M)c>:M&AI;8(::a+PBV/SI?IPTbW(_KM@K1^C:E4(=Y:#O&53:<b)FJRIA9-
29JaP8>LD&(8=\/@8MMIO-+ZR/^.A:d\B+/(8SB8;SD>KT]3:G],4EMEE,dWAaS:
cH]P\aHF?aG)L[[.YeV[V=R<HPS;ER^9(YH:2CK;OHgLfOG<AV[c1d_W4FD7\Y7S
N;?\b8F)/d3S3(Vb2F4ba29X6,(_9_A/D>.V88T&2+Y1SCPaOPAf4a&5DF#6YGg4
,GW1I\0ARS@\K+(JXc1JONIRR4f3\/?]R8CJBUT9A_VcIZ?</)9Gb^4AP5:bHaEe
KG](RMR26R03^7WNf;^LP^L1IKB7>N.>7K[WPLDM[eX4;@=WJ7<V0W6_9@][-JP;
7L<>/N8FZFeFeAZX>-7-/FJZ50G]==6gIWf9P2?(&#VA-B;g0e[.BG3<[5=1E)3S
-V+dKRYDF0TMM:&)fXVZI&G)dZc_UNSE1?/,NN1&(5@#4^=.Q/)JATR#=A)HJ;<M
JKVf]40IS9_FB[P[N-Z>MHfb<LbMJT9PG=#PG=7,S-VJBe#[Ad8(F\Lg0\056fNR
]aNI0JE?)43+ONE?&YN.2^)7/^HSEOYX[IXPWdAa,YP=OV+#VUGZ/02Z6IK^@=[;
I3A17?6&bZ7F7Q<GDe(L?XAUd8G73PQ]S4CO0^3M/4&SXAJT[HE)a<=NNS7X(G]>
,)AGO0efD]Yd5#54M\DMRF[G<EQVQ&d]Rf&]<7[eIC2UK:=C-.(/_b7UVO)e#1<L
PMYg&>0+6FAc#X\6E-NIGX:VEC5]#KO/U,1d,Ia9F_)E+O_SFe]M&I2KEg_T767.
:(0DJH490YJ46MB;g.c/QLFX[F/?:9Y^CAbS(&BT?G#(_Ia@J:_4,O6-/gC[(^8S
LYQSL[WPN_AGKK;fPcAY)#UdUJ[5b3@31+7,b9;-HcX=BAR.9QH+U+d@+PZ^CIR(
M,ef14H,<WJ8aM0Y[Md\(S^dB_IX.N+W(^c5\MX189J4^7_?#_ETB2-6D.e;U;[f
L=P5c^DTXDUI;:b6dWR5M&0UFT^P^+QNI)MI45ZCBOeE,UDQF:P7N#<AF[I.<H??
.5VHYBV^J1L?]>E2.0,YSO0[N\3,C?HI/W<d<.fVEA1W5?@Xb/6X;LS3=TTI<JcZ
VU6Nf\9499N+YBWW_/.\8/K^\_VaaE_(Gd6W/@a1H:USgJe8(1O0D]:b510S_G0F
R5HC.=-4D<7YI#M3QK&2RJXU^>gIQ\])[QDEc1Z8_J;6&[D@F?2W+Q1IU0bJf:7)
a^&3\1N.E]Y<\SaETMQ6+UWeYC(2NGaW]YY4(K<D9DW4T)gJ@+#H/B?A<N_[WM5C
)5,R;[<B0[eg+g.:ZKd0TQLW=+Y_PY1W\BL46TbC_26IDC[d&]BDBgW0X?&?27=F
Q\+LV47;O49dcH<)FI_,=V5\Gcf/Y:CMOUKLWM=8<><2aVE/?454:fL_1f,e(]W+
/eUJ>=fN2C.Y:9ZTG)<HBfS^NKA9gX:88SW@)S?_SG#Q^.77dFKH?Sc[Of.1UYZ,
:#(J]YLXR7]Q4B]12KRAc>VK879a^J]dVRXMF+d_#OK^8f?9VAb1YDE:Z9_f:<94
Z4c[B/GPLTO7FJ92P(GL856I3Kd-WMAY_B^I.(9Q5A]<c;DI<<W#N5K\NdA)T(^(
L&W#MQ\Q7;,_U;#3)/8FHLfO\XXZ+GAWeBfTBa..I4\XTH,LVSQ+e4QEeO;E2W-<
\HM/=<G_-_P2IU7_#D1R\UR4(>WX7_WT9T@<(\>;A0IZ-<HL(M8EVE;NGNTPL)Ga
fQSZ<9Qa3cW:-0;K218[GF4@aOGGg?2fY[B;&==>&^8WBR9VR:)#,(+&ILaMcB]E
^G.3Y&KFOeNOV+P&gE<ZHBd=e1P,08;3CK/_:T5[R^?J>J]K;F^RQPPZ1e&3L3XW
#Md1eZ<#R.T^2#BL7N/8V6S^6K>H(8M;#9a@7e<Y]Y_DTX8\]C85DYfR@]O&\>SH
KV;F9cT5AW;S55D&[S5+6#bXVAGHI=U=K2:CZUXY@H2-3#@XD1K,acJJfX[4Kd&4
b8ARR7/NZ,\Y:30FU?&RdW#JB/F5dN=IH3Z=GGCbc2df+(fd[+d/F?)0/#dNfec]
g&3+.:e)M;b\W8I:Ac>1JW]OFX-0/(O&.Q3O@;.WFQ,c9SCLWTbXV#T4J0G2_3BM
P:@Q-61((T86GR@..Rb>BCQgT@5S,3Z,b3\dC/#Y2#8AXIK(>TN@\SR@X<SM1_.P
YTUUA>a8K5/NdS-^;&[PEa65IP<JgaLA+C_AYf)T.1,[?U8?dFHCW[D?4+5^4cP?
BWZg:A,=7Ac3MV#)GO9aY@N@A]NSMK-)F9:ZPI@2CZF3cVb@/(8]SRAEL?=N.BQ1
M2^F,2dERFC[0]:/2K.LP47&-egb55^S\D]Kb8]c8.(7EBeW?cF>EbX7,cGZ>aTX
#^fAg9:X?UfG[KR-HS/PYCPD;M@9R5e;:B-PAU[WaC4K=51_^/dM1L@4=8UE8@Og
8.PY8MLODYX;FER)cHSV2E?+&-#11LT=V@U5gF5UCd.-\N:G<C9TeJAPD94KB3e7
RBIY+<TY3f^PX<fL2_[-U0+H9D:L-ZC2)FXC;9?1F@O8P(6f44Hb85aG(f>dCBEa
2gSID/H4<A^ZPKYg-G:83f7OO+cE][;O(SK\5&V6J+-QO\VKM[6c5AbYO<C.eLJd
E3UfQ:EfG@0GZ-R809\2Z73==DTAgg+>#P6XFa[ES4Z(SSU1)2RfEePT]Ac+a=)@
E;,+0[S8MagJ3T=B9c97acU]Pa_eQJ,Rga)9dO/@aX54\G<7&M/2.HG:X3]^)WF,
]#fG_INQ)/[fc-05a2IG2P(A4GF<5\2MVK6b.;&9:-7Zc.A@00^UW79b5DYN#L=A
@6:85JSLD#QDQE.E(=@NbPcS4Q-U--LaQ6&6Ve^T?]8UB\E@1=,AOE#J2b^^1NZa
7I7(f>UeFf:.H\8-S+\ff,g5;8:DP7]8.:0\3DUg)1EL&LX+.)JOD\b:6f\_=I+Q
ZNbTc;G8b,e1eQQ7.eZZ&Z(,Y\-&-?T.?;^GS@1+#[F30MgC>PMFBN/7W6I(T9_)
:H/TO?GLQ5AMUbV.Af>#2fK]XG&FAA4D0H.ZNK25ZMcCcL#PPd,A#EBPg19,JfY]
bQJbeX[(8Me2f(Rc7XCf5V24TF>:9@QaGfXf8a,E3g&d/F0P\Z8Le)H(A-9B,8[8
8YF;=(NZ7\_MX->HO90VV&1=X6+/+Y;BQX:@)He(RM;RB/N@X?ZGQXTD28]aVGJ8
9bSU&),b<\fTaf&XU+=,P(H641UD5SRSM2SW5X@2BP.M[;HSFe8>XBN_\-Ua;YeD
SM)LXM[NU]>W4gC+D3E-PNP&5YEB32gJ:eZ0?JGB+Nf7cf^(5dEB]W<S9aQF;MCA
VDKPR989^+ZE]K=a<7@TNIEZ7>MZ?Td\\1<TP55aY\ec.fO-Bb-Fg)ZegQOCG-A<
VN36CH)QI410X]J<KR8:7[VBIfLB:A/:T976[18I4+Z@E1Zc7W8T<feM1\gKVI^,
7fV],<?T[Hc_#+;;TNZG>8d][@IE]TL7S?D_,B<&I?Gd?QUQB3I]\,0U(=&@PcG(
KI^;6+Z7,.E,I5J?aY)P93QA7LOI-)2OEZ[RBYfAA@,d6;Y)2Qa>+F7]=^&?9OVE
G3#0Q?S&D7d,#PBO24T3\]R7KXAE_J6/VWeP;Nf8FaBf+7aI@/P_Q@COg/;,5DX1
GSH7U3:A&V<M\KULfECJC,+gSC2KTZ-5d_Z8V9f72S?bgWT-6OMYP,>\fZ+WI?YM
ROBLgV<61Z5LG[3/[DFQXB7H9^5Y[02\<08/62R[U^ab0HOTASGEeQB3g@6]@TaD
IUA>A9P[#NfP0]<6AFOINfA\1W091\7(L2.::9S=M;:Be<9J._DRZX^ATERSYYKE
@ZARIH?.59+:aJF;;-36Y4g(?B-EfDcVc<R;EJLMU.BM&5_\_FBRBBR/BB\TF3Y3
NJcJ8d5SW0CV>V@6HE+DPPQ&>gf1c(<XU_c6YG@94_VbaD,SDTT:R&_dNSW@IM\0
K<\Oa3M.VP<=)#S/g;V?(CM9[^&8NR+/&93b_1#W,HMX5=H6-J<Q]HBeP+,V].08
=S]X@9)QOUO2)RbO@K>&N\^D1;7EEfE\X<LZZ6M^19>S:^b#F..,=M/Ce01=fE8\
b]]AcE70.g#5a^(f0?U#D1BE(IF]3432-]OL9@XI_AJ@OLeZVT;_^,L^_4S:1aIH
QT2dc+gX^RQUX(1I?=Kc<VT&<8LGUTg7_b#5^7,gC)T7bbOX)+@b6@fROIEY(+^3
gH(R3S,_;+G=bHaN7[AgRAVDY6[61KC<8,T<f5/6fSLa@;_0F>K[@:T9B+ERXX45
&GWV8EZ3e+?0POdK@MQW>19K#35-8Bc?Zf,F&M8+L27\0L.3Nbc9M&N&Ma5d>)-A
FUgZA+=a^V&G4d\,FKA^[TeY8,g<9?TL9TPV>Wbe0<2JERbT1)G>]^c9<,8+4d;a
.c)a1PXgT(^IfU&aV#JV4Wc=7eY[HS0DC<\@)R7ccK@KX<?Sbe5(.NEM[3]NM.T@
0Q8DG\IHcBMd5/agc3^1N&&J#U_T1>B&@_LgS6J>XDG6#(:R0g\T]CeVMFbASQQ#
[I.D((/,C?b;d1::4<S5&75V+4YXDUQL]ZJV[RE#(E#L=+CJ)f[1>&G2\GY4G5]M
7G=#Xa/Q&2T4Z&K(FJ6G03,XON>J-ST(C8A?9/A>e&-W-.^RTV@216./PDSKf0H7
YPAX=R4[+2QSecUR(0TObNC5[HJ?c:.2MP-;3<a.[D6DOXM:T3SW_gE481_+@9VK
2),(eVVXD5M)+[c:K++b-Eg-MD\X[1;XA:((3_T=#]dWV,M5ND566=#8XKZ]LYU]
EDOY:Cca)&P-UFT7P9^;CWN=L_.JYD667-fX[]5+RH9\=([AOge6e\&+IW?aZ]93
>TSe;J>6:IS\OQZEJV,FY/.R5Mgf(H[If_)U)-;5d1HbZE?(H]bD4NVfS4U9IeG,
_eX3F3#:F>LNPJ5PAR/+CDag,GV?^&+9WA?Ic,M#[fSHf4#9=Fd<L,7ZSTJ)5<_7
5KU[a^CF@<>0af[8YMH>c</-O2.b)<)5YdcL]^-SR7-=O#eRVSS,O&9a>H^ZKD>6
DU\:<7#T_.M8<\W81AD-#M^N.\DRTN<2cPMgF;R&fGN/UZ=Q97C91Z,8Y#T(M>1]
_>:+;:D#[FA(3eaED2eKN6:\]D#G_\A4-Zf:5ZW^CbT]GSOUX.5L+^51N/O5V.Lb
geb0(e25ZGcW.4Ze5FDHfHEE3Y?)E=b\TcJ3X_DKE]Y)>.bCSBXMSeg0(7R#H7,0
4\H#,X+QY2D10J;;;+KU>6d^+?6GA9V+UdZX:4^<\^-#/]^PCMA_XaZ0cBR#aQ6C
K5QU6I1/R)9D^VG^fN4YMN#</\Y.&G2ZEaB^\6:W]_a8IQ+P?UXEZ^PJYegggO])
Uc_0Y(=>/4/ec_\Mf^2:0U58(4]F9g/ABc<,:4M7\Zc(A6NW^V<3TfM8IBR2.T.)
C_)R_8JRgZ_480OG,1MGH++bY;YIJ39eQ;0D^9@IG.]8ZUS6b?<?VO5Q5UBW<S[2
=4@_VbL3MEbX)B?TBD5/J[a(eLGAUZO)^[Af:+K=S.O01J,fO#UAOF-,TI3?L@^d
,4PT()C4ge]OC72(>I+N#D@3g95eK3B3&J/dC/^^E3ZCD2aTV]\><7HN&6-@U.Eg
(II,Hd&e-EaI)0QM^eC36R@Q+<S2KF/\[\3d0S5QDaV5Sc3IJ6[3]::28a6BP&<-
X;1a2Q138:2@=IHe-<c(#@GXD((EDPG_b;74LMG,K#NP2SE]N8CZIVV,R@.b^S6A
VEc(7-?E+STMdbA<aPXJZ6d@)aS##NPDWO^[4(U[JI.e]])T9+,@\6eAVNNHM)^E
JST593Y]2/IP6U43R]<>TWdBZ/0/#LHgdRGT,EgcIU9bJ^YA2>9<:#+dV]g?LX_3
YR6&#2a[#ge[8RNB#@c076#_GSa(EA2_D&,a:T5Z&PA+ceO?0=Q?241PJQS=2d/M
8=9]9)](O),=3&g53P1H6W8,3K_+N\DYG=7Za82cg>c)f=E.21M\(<6@KGMf],C9
Q[b7cBBg9S@COJVR\:@\gAOPf4cOU+dLFO58H:G-<5P-78X(AD:D2J<MT/0:7c@3
&;JbV&Iga#?UaN7SBD]N]N4;YE^2O;de#ce3.^.3FF1KJMN8:X\GN=[Q+ILK;O@W
:c(b?7./FR2CCbGUKa+-W2G:)8]&KP5D6_:<df/L/.2)=(AW]_a:7X0[8:ddc,#\
N+[IN()PBGe<5BJEf[b#]R-B,c5FF3eJU4;O,:1ZNX0^eO=aMVeUd<,?EQ&YIQ^2
Rab>SH(S#LW=ZGL+R5+-[Xd.229+WHdb@9,f0QFQ3LH_<H(IN]/9V0-LFC2^]ZMO
bT7b()E3.-QT-,XdDa-ab4?ad&fF^\JR>QQMR^DV4@dM^8L;H:1e+XSAAB6]]WT^
[d]5JY]b7<ZfC)L19?B9;8H(TOUQ&3aY4@B4.SZ)6,@T07QXKG_c-Va6H5X,#(Vd
6SFbFRB_aRX617Md:P+AfP#;5af:LadBFR=_^gdXGULJDS_KbMU=V3^b5L(b=,X4
g62ReC(DTIML#V21cSb/11>4U#7f]HJ5EeOPecdK+Y5O@FBc]c7:D-<]MA^IDXN(
+cUgU5YE3L<5BS@2=XOG29ES]VN?0=(dNGTMJe1E7Y=SeB#eRP(Pb/A76Ba[\gb;
#F10C2155U2NG=Dg-[^ZKAIaQC?7;D1(_2fUA4gXTG0,;GId.PL:X[2YY&Fe-?I4
MM)(Ebed/OYA->__C@2dMORQ5?)<&gQ]6?VA&_af\_d:Dd8#2\]#P1@Mdd5D-E<_
5BO>;,T><RbXOWLQ9C#;>C8A_/?,<8d+Jb,Ga9U3g:D4WH\=#:LJf2P.R30^SB]#
I/S#&Ed<Q&BA@:##B#XM)9-B_BED.BB1+_3Z_4N?>1I6d3A?R;0U)VUEQeXQYC&-
F>:4Y)3G-0g8^HN1FYa2bD5DXf=IK,G?Se3:PSd-PCN^3(G^8/;dDa;R?Z)V,B:E
X,BO=@e;39LHX)PX0)R]R]EcGc\YL5TDdMB&4\R12J]eQ03UIE3PPIU)D_g,\6(f
cRYFA3?C>MS5gBEeL&A3c)>WF&N116.TC^RNHYO/:=>GK7VT3>a0WTEAV)6]8<3-
]@C9YK[H5AOQ_dZK(?QdB\S(aDO#aETE-@2+&/Pa0Y#BgUQTcc@Z<4c4WB_TR.Y8
^]C>fEAQ51Ba<)[1d?.N8GEf.eWaB02?+KFbfC^?_Q,Hcb;)2=HCN]fMbBMS2X)8
I@3fXGS_R7IB#H08OD#0#8/OcR:W341GOaU?+6NHTeUPUOV(04IeY(g2VTg(-3X[
DY9J];MHAdddNOLEg<[g<g[[SVC5YS#.cM(+b>We1d]#44PD1@/HH4L((W8(666Q
/?Q:N+JO7UF_d21,e8LG7XI6KY0&@/#KE3dX3X[EXI8d<?\[5+M/HU#V.+eIL4[G
gTX+Z-aeKXE8&RFR_>-gY?950,W1c7cCLcJK.57=X2Y9Y6K&QR9W:1FS[@ROAgg)
cP)GRER32V_1(S;R88K0L-8AJ7HL)],3\#B+Qc&S2@.C^D;2#e_1O2]M#fNP\H+<
MBF<1NM[&>FYX:?;(@P-1ZK1c-.7fdL+d.N-aI@:@2JId]5g&UMGR=3T5-dX4&53
C1d2Mg<Q;<c/=9=1;6_J,g.XWI3]GPHY]<A?L)FSHVd9I[ORXUH+L&8cJ]AP&ea2
EWI]=PK&ab8/&^DZ+8RG.&>D9FgDCKd4Q:AX),S#b5)E)+8@-gVEEfD<R9YZK_,]
f79:?&@<&R1]>/?aVWBWNEJB6VfD<f8F+e7X<3&/=@d=c,WM2\#)YF8J6-7NUZS4
1a3\&Y9X+JORGIBfDBNg4]TV358V]9Y)9^B^A@YU=)R5bHRL-K@OU>afU04_14_2
#,8Za.16FCIGZ;PQBF<=?T690D)U<N&G(1./Y(UE\e-5RBP&WK+Ua/aQP,Pf4Y#S
<[Y)5:Q7N.ZXG(7W#g8U]7_Y-AITb5@J3.TUMR0-^aad7EXSeR?&7<0+6+V=;g,N
fFBgRf\99642I#ES3a)ePV7?SZbBE9XaI\/4,^3<3fT:1U,Kdf2GBL2P7FM>Q>gQ
3)Y#6e5R1NMB(g3[O#.T5.)e1CSE5g.-E3g=,Q-ECZTRUbT06^(cVA)0\^P.c3PV
TMCXF^f#&LdL\\;4@,?JK.C13eL[VT=#B(3Cd.0,R);A#4/0@?Z-R&^M&YQERI3T
e>NJgSSFIDN-QIMU9(TSZ[B8)^+&WBQ75bN6VM0UL(P)Wc=AW2c_I9c[,Q#W[RE2
PHRC@V:aX8+[Ue:aX&SPA1Z9(5#<?(?G4J_7(=H2S+(Aa6&XN)V&/YQU9<.-C9/1
;H(/NgdZ,?dUP.-#,BHP(;D3UDK)fMP<EDN#343)f.B_LN_EIL\A75_DZ=I631_Z
d.(L.2>5P=JZ.\\FU00_g?+#Cb<HA+)aQI]Hg6^fL5Gc]+V^[</KcY;XPU1V(ET4
0+?<L#9KC5M7b78Z5?VH5a9EFd0OfEM2Ze2;]XJH00<510L;3NB.QHBfU]DgPBHR
TM>QOF=64<cf>N8=0.e5\6/NN7@L+C&H6TbR6.&+4eO2XOHGJ)ZC+C//Y(^;^^OE
fDg?^0-dAfQNS3G1H6>YX?2ZE(/0?JO^+CD;-ca1g8BC]99&>&[+4ZaR/NeYCHU?
8c2<dKg@^Z5^aKY<7QC&V<eGOIMbcK?9^/KRCag>WKISdNF^Mc_(\F:V]XGgMOfS
Eed_)ORU-ePTf7[Ca;^H4H;Cf_PP+FT^QGHYT#db1;:PL_]];RIR/d1M(O9N83^1
QZHE>d2L6><aBCJc+QDe,BSN9MgUDRNPe6Jbe?#]69PWYZ;89DZ7(1b]>1=YDDfT
89]Vg<<D7&/I[0>G6c[^+FTEa.SSUd9ge>T6,NeP/S[QS^^+XL?S)CK/KQOLDGZX
D<U4T6N[gMaP?aI(Ba5P-:@d/I>&M67,L=eb9@B_8;C3],N\?JcOJ<O&2/,?ga(.
&H]-LO([8;F1QePNV(\[/QT2TgBd,];-G:GaISR5XO-(K^<+LL7[8/QQ[ORJBTf?
6FBL#0@+2:3#9MRT8<HFA(egE/aQIQ_cMHR5XfeET?O/06d-7(AgFE88\D9LGb1^
]L;/7?S>7J]/R9OE]Z>gD4,3@YDa)R7=+_7fBd.EPJR?BeF(dGP90AOWS.=FAP(?
4[4FgQ)I.#?:82eC2D]?fcOJ78K3M(<PB)+M^>1:>962f_N5AUdT,CH&?QW]PN\J
;4J\C\W<^8f5_(eN51bN>f14b?J.QJ<6:NGVWFC-+PRf\ET0++\I^T_WKdK57)+)
)OD<cC)?-WGK9>YSVW0:O<7eGaaR([Nf[=F(M3.&dWN-82O3/I#cVGT>.W;X2.ZW
;^g_>KDHN6QfO#EY=dFI11Fe.)aL&:M/ZN&CE[AST5ZLe#]03Cbf_ZVHI@4eO<./
3XV5OF&[_EH<5Y)J&a4[#I37Yf0^_@DN2DR93EPSFg_F1&GM9>IB5;[I9:Ye7S+S
U^DL>?P^K1MRCEQ=ME&E+#2a:\V:0;e;L1\U[SV)Vfg1fP0d,cV&d1FPT9^6d6JU
3;XKeU3ZI1]?9#I,XcYRT7MM9Z;,?MQ)M+d4a)LL:UFb#.AKR9e)C57PUe>7fLM?
P--]:<G8aOWO2c7#g+c0Wa_G>XJ>)>D7&g;B0A;.6#TNTT>;V2?G\_])-&UV?-^D
3]\I(WXZWe_-L.^6@_gg(>OU4C.LA2-ZI;bY0K.C;+L@0EAFbS8]ODAU])NEP^L]
bDcC#4)3U.[IfLT-]@2>X+2;E\D3(O76PRNA,X(CK.[-#<]6:^?.N8OC_Q;::+Mc
)P>LGO7=T]]>M;0LF3V[\NBV9GWCBN3>UV2Q9;3D;I7OZ#;F_+#.EVMd9L@>@0W;
:1[\Q[A6fbFV7\GJaALcI133RBfL()EAXSER9ELeLZFYed)ZM,_>6Ha5N.UJVJgL
VY\U?cTeN.XR<8F6B=OB[\GS;1TJXKP>,c.ANG2Kb8cI=T;,9^=2;7F589RDAV&+
MR)C#OR:;8(;Q07IEVSS[G0;576\_M?Z6)SLUM3Cd:#RgE9aSDddDW+ZPEGWZVf6
:L46I/;B#6?@DZJ:@FJZd7=LL3]@PAN.QBd?,Xg6]\3I#Bf5R#^2ENUB.?TETSdO
:E8N\L6UbZ^WV.0&TIXfFg4CUG_MMNS8?HOc][.)J@J+A0_KD8/Z<GR(+>aT2K3Z
b934V4MCF\([@dU#@^4\PGMV>E@>#VZ<f34fdbDP<?\;bD0<aH9#[_M2NAfGH^QD
EN#X9)5T;=-MEMX21)RR-L_@6U3OTU4)9KBV<C^+Y;PF2.4W_.C7H]GC?,H6<fP0
YC]8a4+^?a?,(3IS+C-5e4^2>L+POXV^Z=O<>BG#CWZ_L[AFDSXZ26LfU+73[QP<
(.I2XEB>BOE>&D?^GWNCcPBNS<1IRA#,<J6)F-9/8L_VA=).IZgL:O/1.AAJP4PF
Z-4L^)3S8fd=;b#/4C\M<[-.1g/M423W,2cA@W&=[01T^AHOfE/R^Q9AS2e49a;E
FFgLG_)HHT]]+f/1U??R(.0gP9M=H0^0:TACE_UVAO=ZcPCa_JL[H=:M0S5@0\@d
f21B052+Z>]K8VVF\?OM#K_-@R7bHSX6-#P/(d(7K_4B93:_(L&0C5+QFaZD?3:a
9A04S.f+@;WHL6a2(Kf6-;FZI:dY0O?B7cf#IE,)JTH2XfFZ^E@.JN9Q2K+Kd5VF
1]/CK/GGe@+B@ecTe6@/2bV9?LZ=.Y5I;5KN6,=?E?RE==>70F^:EDWY.A\YT\06
5+Z^MT^QQ3(^:Z0(8;ACV86@U,]c>P5IDXF<[-S5fT&HK2d/B:02eCbDQ,<LN,LD
<C8Z05cZ\_2>CD[F.TVP[H&X1HaH]9WQ^BdOeI_bXBB\?H=@[L6#KeQ3Y)2<=AE0
dEE<V,5)VGW1@,G.aZg\GVeA.-5(2SbLW@,=HNBN^+#/65bMM2XBecN16;L72Z/.
F^,M#Vd/WMG5;EDd<G;^Gcc>17Y<3O-I\.,BOb[=gIfQa0&fLHW,H.BY.<+H?]KK
a)K+XER:-IE3T+]F5GPX62X:,PR1/#1)Z480;ObUa[W.0-I+15?DRN>9#[I:_,dW
,RO/K6aM<d4S\;AG(\RX@cIM<XT8g_[)GJQd.E7<1c\#2YdX,9?^>PQMO29+e&<+
6C_(<Xc=:b]FUPGC]TH2N2&KG3^1RL4M0ML^PE9]ZfNd?#/0Ug:Y[WKETKFd4cB<
Dd<PdIP[PTJD;;S/;BB)RR?ScF?5XRZ-c>&4PCd]=SM>=QeY/9bXKa^TR1NVG[WL
WUc,HNZN6dNC,d?\V)KL9@)RC;d+X0fcb?L.PMUE6+g;:,I1&:A]P=HY1gf+?H+E
5]4X&:e-MBd,6-<,b&CUaeV;]/PT:35dd>5Xb@7:]]Z:)\aI:.TRf:F;fO(ba2E.
FL&3G&P#G=WW6ZL?LAHBWSPdPEAbGH2T.LO2EfgP(^<Pf\J,X1_5TBITOX6Ka4_E
/ZB1M?C8R47Q/c3_GOISB.JNP.:X7_8Hc@P&7.;Zcc_FTc)KMVD?#SdYR>BBV>.4
cXa8LG#H,2I[[D6\bB1TQ#N^Xdb(7_PM=;Vg=VJW9:=--HS^aG3S&6PWVMZ#cQ=?
AZ5RO@:O5&Vc/QEKF+-7ZGcKTdA\51Gabf-Df;=#[>#RVH5XgQUg&g08R^>Ae2KH
@8=V6-V/C@^B0CC\GD/H3L8M9#LbbZ(LXgNfaUBY-&\cU]IU-:4<[U/<gecH2g7Q
.#>H;5RLZNOK8Qa7FT,1.#=1GdZ2[W>ITV^?F>HX@1Jg_25<[X,g9?,,R.&#4Y[D
;,+V]F80VIG@HBVFK19VcT&aWAWR)MYOT/K##/eC]0TXVM?FLJ[gT)8/RWPd3KG:
_PFBeSb8:Q7_\S-<MefEZ)J#,)OO39aW3.NeM1?6_#O93;9L<>K9Zg#=?DL5XF9-
ADX?L7RGN4\1\_2>gWA^a.f<LY3D;4Q&#&GG?\)8FMF8\&AYVKT]e+Ac25eZb?7;
31<-3Y.TGCa#Ag_J^KK#MF-88>/-f7SSQXY#>e=&?8_aJQ@<a+)3<OF[bB@YD9.5
F,VPcc7O>QTG1T8T.)@<<3ZU]4GM:=BXKd46A)a2N?-5H5I[];SI?2W3():X23[,
_N)X><;D0eI?XD<4??EYCM0fYJ^.\T4GfBS/Q?ag1)<_59a<D9M0ODPDE?-LH=[5
+<0N(c57[)B/UT6W9g0FPLBg2TcY_)6d/(Sa3dM&D9VdX8XE_Gf-0F?CM)Ga=1;d
?H+(NNLL2CG.USXDdQ0U]e@6gG8]g=.G]e@S^Fg@)PR+UR_=4MSSKYQ+J&U_^TK[
5[;75(Lg)ZN5f/.0.TM(/[?EP4\)2HG(+e-=QH/K.51IM[XR59NV0&<^D,ACe(:W
RAb<9;5:^A[0;;H;<RcV0S-,gM;eUR->]X^cA4+D_8b:44S/8bF:ab(0dK(#;.UY
YY_gS\OY;I3&I\;JM@Wd:X^/<6[cOS0)XIcdQX9X\)QYXb\c?^&<UCBV:aOBI@KE
cbFB<R=WNXSa:<_;4^=&&2cAFBbK+JecM8C;I-H)=e85K(WK(E[M90a,646E5U)8
2D]cD//[d]26WZMg=>8?g0^#-C]UEcd>8+JDM.8V-+aXN&.FIZY(D(e)6+8GQRO_
;U+AZJ;@QS6LGWP>YTGQ_[>a:Lg+\=N5@6@OY82D#\,a9dLS>>[Od.6,ML8/J4b,
5^_+IIQBb0F25O56S,MLcSCVSBPL0-M&USdUa/078^W7:-PC[aC]C&-NDZ4]Y:gS
-19HK=EXV#_3(-.JQP<?=IdJ[DVQGUK-5c=/Q&/8CR2IfP<\QD-(G_4Tf-c-S,1[
;KUdJ&44ESYN5&3?1\<G7-D47Z\IDVZU24VeR8[\:>16UOT[e9H=G_bMJL4->Z5V
?Y_c&PfPE[^e;PPB5c_&+/>OT)1BQ_HOd)Odf>XgOBP#3Z#N(]>KCMKfT(<K??9E
T,eZDMFYRL8M(NNX_,.7cNg.a/HXUHE&VDe86]]5F04f70L:SP1-M3ON=AB502VB
_O_8U3^b,#9Z\VQT/cF<_9HG?]Z&?B@D\;.\>O8-NZ+a/1_F\<83bfe4X#@N&\8)
G8.;M41/@<IZOI-a&M3PLS0FZGT^NYW7^2&+DLDI+0]FUWH@5UF-I3=Z[@,;KQ=R
@)/4P,4H38\/b>)3P0O#+FHQb1?JG/Bc&ZC(e5.WE0Y@DAL\7KSH7WBbOXM9=dgB
Y<:L?SMM-.S3B9P?EC8ZFd#7D(W4?O/^5acMg2dHJXY8g\&ba1EP7=-B<\P4U16A
RZ?ded:_IR#O3\SSL8)QXOTILEUSXcM8c57g0VGFZQ0H=7M0/<#:I=><[:(EfTF\
^d#__^c3,I+[92DU?+\YMMTbU5#=b=H[Z26KE[V<(,X3[ZZb?O]f6aO?YADK8CH#
@ZP&15ZG9-E(,e;C]9gg,8Aba;JFUJPZb_?Q]d1-=((g#9J>ZI[\[U:D66&M?2]/
-37ffWOBW8D4(@[cD7[3ccVDHI78^V?AMV3J5(EGND516d9ZW.D>&U?G_O:&19K<
H^&/XI><bC;0VOb92<AZ[0LY+>4gGE@K\0JDUG16FWI6,LA\&6N\BDAZ6J2->Fe]
e?2R#7GF(#QdfK.>M+g.&Cc?g1GR.1Ab+<EI+@#(PK^,#(D<8]VMQgD4eVP321a\
TY93O7[7dOaK@^,3R1=QU#40HA2[J3W22b3K;_[)5TTIgM&P0W)R=JDZBC4Y=EEN
PcYS>&57\@N0,AXQZX#bD.8g^7E/;&SVVcTCMF^gUW&.RWBN+ESIcaW?bJ_d5>6U
]5G20<BN]Z(=LK[I>=b1;I5,=F_ea1(2YGY1HYA+LNcTF_1M^=55FWOe@#FT@N4^
7VWP98)D/MX)CVN,HPTU5@2.1L^WE4&cWN]DU^F0_#WLCO<IS1&\7c:W@bd27EUX
?gV42JJG9W_;^?7,EcIT2YI2X)^a(Z1AVW;E9MMg=Y>c2@7DJ<5T:F;FWcc4.M-G
KT&&3ggQdA:gP4_WJ&4EB6UBJ4Q6;_Q]ONgZ/TQD7=YJ10N3AELY[I@b1B);)GFV
-3)/?)\6M5:b;g61Y<7B</NSBI3M]8cbO76N6+2&b>a-IKZ((XKGOZL,SeI910(Z
7G?Cf<64.#CL#0c@Q4BA_cdUL6Eg+#)_.f1EYT)=TQFJVH@CRM[LH^_3GYA(eGME
>CCGRN77BBDQc?U-0E511d&@H]^H2RA+-1+Wa,OfWY5bR.?F@?a>.g7<Q8Y>#5gF
N11CT.?>ZEga?\&:Cd[cQ>f:<5<)f7-U<X@^G)MQaTJ15?.64\]9c?;W.M:RHBI?
0a1_2fLN]fH)6L?]]D&@_).a;bHC8V&R6WHHX9[Me5e<VI2&1(U>7dfP[=JZ_\+C
EeIY7:fXU?9<)N^.UdM1-.<,YTUO0YFJ#E>g9ZHN+28K-#RfOEE8&@U8eLHT]4^Z
L4X(d<;]QH<HV#84Q99e#.FBWdg?c1[(C2c&b>29T:Pc\7APN,.I6M4,[3YH-<4E
F<I&#8DAWef,.gKU(^-G;1F)/dJD]a+HAQRL1CG;JV#:U3&)[M:PIHZ@+RFL;WXb
1-;b4Q2a]Q]?1cZ@fS[GRMAN:&HVW-ZOg#L-U[9V:[?X)Mgd^N7Y?8GNQ8XC594L
)&\]@cL^[b,=9X,@Ac3S7O3,O<T9=QGP>e?.2I;[(G69_,]UB5eHM<9PY<Df^B3@
e(8W(TfXX;1X_9CKGg(7e/NCLSI[9G9f=3K3e8_TG(\2U^Z3=NZ.QW:&+;PF]KMJ
]71e#&LF,B?HFBTZ?OWD1R74=P87_J]85M:BSg(AF/Q-S.-M2EU4;#d;5]/g,Bc7
KKbQ[ADQQ0TegJM]Aa2aP&_I[7[KQ(N]W+GEV)f\bEf(,8e4>fBV3UU)4A29cAF#
g2VJ69.8=W>#KF?f^=^5SBd/NBJG]777#VLV/R.B,=QO#Q/2f@2.0EO14J^ZA0cc
C8?7dMC0VcLJfGB++9==N93+]IKO81)094aV^M:VAcF_>d/c9L2TP3HR4>H3J3OL
gCUPcf/MX^O&PW,MaLe#P()DTZa1,?a/T)5BZ4\K\0)_)BMa^KM)1Y?IURCdF.0f
K6)A5QCH^V/R9O>MI<N<0K.,PG_Rbg[KHa/#aB=Q&X)9OcXeGA+Y4E-8^4S2S]#1
OME@\.e]MBN<DG9WaKa;dJ6#MXIE^J:3c6(UW7d?ME]e68aH4]LC@f-<.>f+(@DD
X^3?a:f)D2Z6?7Y48F0^67J-4/]dR3<3E/&&2M.1HE/OB5/5=bPf[_\B[S@gdNa2
KSB02)LTMQ9?/g,]e?aRf=#6^YRbED,/#LYXba0VVJ;;b8=<g,#,^[1=&ea:W#-Y
T^B[,6]O3L.:c;,Lc/(-DNN<EMHea>@HD,34UIf<C<G&I^f>Jb>.N8:T.(fB-ZC<
efa0^+&cb.RZE[P;878fGDdJ&_EHV<30c:1<:PPadLIbKJfV\E1(QeHdIC^b4M<;
60>L,>S]\6:FQJI]JE\9#0#JI0f(]N31?26^:6?:#\Q,Q\bS,TQcAf=688YZJ&CF
5E&[+-BP^Ic,>AUd8=V7HZL4-a:(\:>U]M_7USLd\#,D_#?99]@J#<3=7^VO4QOV
.H_P5ga>&7fAVC+6:O;gPTf=)9#398B<UP(gYAc+Z4\J6S]FU_VJE+b)[#G5EG&8
MV7(#cd23UW;R9N\_4#;X41K&;Z[8=Q7:b<I5AFQcUGg4(b8\De--Ma@D#X3INE3
CP-S?6HGVBa8)?-XL^.5_N[&<D()OPSNPAC3gXgFF8G9#YQU^9abG20]e7a;P&Vg
H]M/I/3c3M.g84W,7L8Nb-C>X:H&I+c9CdXMQ\A@PU1PFQEbQ8RC;fV_5Ea=ac:<
.S@K(FSFL_6EKN9Z==K]V)I^g.,M25.R__)J3#S#VKDN0PVS5O0,W<a/]I[QdILA
+7J#=?aN>.BNVc-I3I]5,?T_:FdReCOSUQWMdVMS.]V16&:68;;NaDY#_Rdd)V4V
YD^,]?WbT&cN+)N(g_#_N0HcX0-gR-S@cR4[F\VXFH5[^>]JE>P:83dPDHP.D&H,
H;5Q\+4H.)PDKKJ3>KFd7,Ka>GU^K6;cHZee][2=9]3MVS?J](D^A]HDM2G(##U0
QY.1AeY0QaI3,M;#NdK^_HHK-RTc(&>.;ZQc8&V=<b>_3:VDBJb:Y1dWUX-Q[L9K
Y=HE0FS;c10E:IQEV:^FO?DcIH@f@[-R\,FLGS=Z]5?@c6M&Z)Q/+]_D4#7J6E0#
CDDKfM6JWPA:,U]6MOcVc:RP>IBLI8W;)ZPZEKJbL>KK1Y)]++9Z3PX_:L4KZK^D
4Y3gQIOfNb8L<H/Na2UDcK/RWH]CY_6M4[1dWZJ8Q\5/Rd@\,-\+_-&I?<:@6H<-
<T,07^ca\4Be,#8+c49IPbZ[)3&D)df(>LP)YcGU;:bKe8<W\R4M9GecO\caWR5V
ZT&6P#0S-M3]Y+V#X-3PMX&>18dSX,T8WVfH;J/(fK@J8^4RSMX=B7?cG>=A9KDA
37\,=R6&Y#S?=(1@7Y+V@Y2H^T-d94)ELW_ZXY&\Cd8>e<XWVW(+^;Q3>TBK0AW3
[O)(])Bd>WP)08b+[:,.cW1X[.Mbe2eM7\Q-:;.L4.#TOF\YK[ZAN.c5O>S+)fd]
2^9SG[H9V1.O(508.5GA\EJ6(5?f<^SZ7Bg.Qa1?,N.>:6M.+WVD(_5A=>IdE3Ab
H5,,2/M,7WM]4+C.f+TPC&T8&<2V_bOgO48GOXZX-&<AWKPg1_6ORO7C2JHSQ0X=
)^ORE=M_K?R=BJR0BD@JG<;(Ha&Re#O,EReV@[2AaM0bgJ?EV:Y9ePYKA^:@SMf)
HI7]=@U1dS/B6>,cLR)1=^5UZ;(cP#ZB-)037beA@:(K:OP;(a--Z:/M@EJ,^>P=
2)A3&H;SeZf/L9<C)>MFU#Fg?=L[Q\6T,HX[DN+gYB6Ec?4IaF5NeCZS\R7:N&SD
b5)@BN2Y3;.fb9Qe^Z3PFW5g1FX<#9,#aCCN/M\8BL-bO[+Ib(V3.<52_A(CY/(/
8+)J;NPU&Be9a/UdXK)TLb)H=>X(RAHf=PG/)+>6F]WFMJQ>VGJdgVWfJH/8b<1A
Y+LZW)>dCaKFYDW7^,;^&Fg[6KcR391-X[EJc1a;>_JN+N4-.E(IaUQB#Z2VCce.
_Mdf,QVTJ0[KCT,(gL+:YO[?b&3Y1+gIHZg1J>N-^>eDZaA7X9>[SPLPg)O]\5_2
:4/.^Y/<aE6c0e-ZbRUEB1a?OC&LR1#75],XQ0=CS2ScIeW&:bPUK19dP<KG:55P
ZN-5R56E4BVU7,<JOLP46?/N1YQB\[@PU3UOYCFf&_dE^L.S^)>)=V8R];<39IAa
0XYaK\>VVU)=7#=A9LIS]^;W<W[)?\[(8B9/QUULHIYTUFT?CQ98NQ9V#R#W;<61
?.(a=)/3PEd0E\3e\Hc(.>gEFT77PbB-KXT4PM;QeN.8HKK&NdbCX?Z;5V;dMd>X
55,\V=@JMVFK\VRP_?HU;f2Q25\Q/1d;NP;=-R&Df@WQH,#NZC[^8L@.]g3;8I?=
ZRODg/+I5T,_]_M.e7M)G90JE#4#M0gIcI\PC9=0V-ed>DP47()aS?7&U5<V-M:O
b9]X_#K&4E1Ee=d,AaY1HCfc^Xa^&BV5QS?#6H,IM\=@cCeg)HI(JP@643,S[c98
AQ<)QgF@M8WZPQ?:f.HeLf\W-.;+MR4<#2(P_5G\(A-6D5,Z(RD?GF7OESUQ4MDE
Q7bI2\H;(W7IQ9KXI-eRE:9KO4?\:_J^6\)#K&]9[H@9LX-FJ+FC<g+gJg3D+cQ5
9@M[g=39X,G=6YSW=OY@IS3_[-48C&eA:W(dfT+c7cJR0b]DO;Zde;9:G)@_K6CD
RX&YJY+L1eT9\DKe177M?LQGKbFI;NOZ,2S:L9G^66V8ce42XQ9T>[71Yd?@dVgB
^8J;eD\S&U>1[>TZ>NTDNNJ=e?7@WCEC.gCcd96O(YUUfERN]0L2T[/XR.HQ36gR
^C_;b@DLEN1dW&(HZUU&7(aS^L(QWFT>4;;OgYM^Y\^&Bgdd9Zc(DT3PGc0V<O0d
EU=(e(JQW-;B0X9(#:dO-[AZDg))#D77)_S4OfR+Y863#6[521+=R@G&<VGN<+[R
3IOD<fMV\V[AR8CG-(e_PbAeKFW:]O:b@HHb:aGaC3;83eRM[EON??5KW4<N9@fS
g;9S4NGL56)/S<<fK[3?KS_)K<&\J<fE]:Z38]>]CA7e8;AQ=ENef&NbVPL?C?W\
RfW,.U+JfY#G-5EcW>bLUT0E;4WIEQ\B6d\;SKXB(S<VBP)LVZ[4SU@TTeTGL/M)
SWA6gS<BDgT8G8V:&K6,UGYEXS3]@LEe.N521TIE?+c@8FafEBeP8(TC:TP<EBKF
V+;E.3U\OO_eBLPfQI,V8@>BLb4?c^;&GQG[fHL=CMb0STW=g#P0,2f[=gZb2VMB
E6,gXQMfA6ZC1UHYQ9QVWTf(JNR-?#022@HaANKFT]eHA6eCIbBCSZ\bB1f96-A2
8WfU]J/DHV?(ON9eTQ/WV]#.0[YL7LQbJc4KQJ+O>K&V2_&\)3dJ\T/;B34:6OF.
&=J&1/7GeRHQ9aEQNK>dINQ>da\TA_5GEP.WTKWYKV_.\0E@?>?RS)-e;F<?P#E1
Y4/<<ICCAT8(>JU09(><OI.Z>S9MZ925&0N^^3BNfLUF>2YR@.7CPdgZ;:)CIH>G
C8&C_dXSM6JY(<@17]Fd^<3T0)c@A-T74FM0JGV4UV#JVOIT/LDXa>HED>Uc(H0-
=BEa=e?_#gIe&+&B>NH?cGRP3PV>+?NF(3)J2Q>>5GV.);S5?8W88:=.4@HfLRgT
SJU2gcR+VRSYO5WbDG/b449If(<X_PG[20d4&.3OQHQAS8+]<S5NgLALUZWc<gAa
D,V\//SF+.;2/Qb+HTDSMJTN3ZGNOU#0cW,^^5Tb_KGA.VS09GJVP1T)OCWO\XJF
:DIKEIH(C6CcV7W@F50LXTJM#CS:^aT9HeZHbgLU;A9P)O=]4EGgY[],1YeOR7WO
C615&[)HV&M@K.bJ5SJ@VeB)ALM_[V1,/R<:eI22X1O,DNAZ1c_Q/;8A&E1_T<Q2
=Q/#IG#Z(R#W6T_FI]3d^))eDD\?[?NWfJ&CPNM,Id>G:FZ;,QCDW(FJeT;LHX[9
R=EI2Aa]CTM-BQDaE>bL;>cT</:>/V-W[&<8:E)NHQVTZFU9&8#&F)\^^WFc0IX&
4R14LI-T_Z.D):O.4(]JA3U1[bN1Le\:4+O\.W17OVI<FOgY8e/6I]<DP4O&WB1=
E<\+5[())4V#\d.6dA>cg@b(fD9;#0EW1VA=1V.&V]]bYf3HDQA1K9IT[WcE/<M+
>A\:?QP(#?>;bDfbKXI@K8=3YWE5GV-dgbD/WCW?GF>PS@_f74d<H-S,O1T.Q;RI
&H6)f3]F+<34d.G/c0@SL:XFW@6SUX2)&DcF7/]JR:g)WYc#VcbR1fMgEJ2eDM\<
eX?P0cS6;DZ6J)D/acEE<SYU[E)U^<#O2ObLb#6#S)D67c-^>]X\-79P;Ka29;5<
C=0K=eBXTT&=]T=X+4<OYYUbQ4^17FI^f(;;W=O@;,;O;ee[G@<=gECM&FC9P[W4
X<(30-08a]f/V624aQGF<f4CZLCATHe<RE^9D9)c67fU.<4+QWd+_<a3&dB8H58M
_R&e<02Y8F.4VV33V_LE[;)g7;P54-D+]bDP:J-cQ@>5T]HE,B1+gXdg1aX=+b^c
J5[-6fND\@Gd9SLC()HE=bZ;BQIeG6H8=c<H/gd8=@?cN&,NVSRf8X+UF0dc#[<.
X/-b;(>-Bc9:>.L?0;J:E@7\_V8Z@Y&LSQ)>NCeI#3&?>[07\16^B=c13M8JgW<Q
MD>9V7N(4fGAFWG,2URaVB(SY4)(6)K]QC+:EXO9[IW_C64d)[-bPFcbTa;:M>5S
P?@_?=UHH0+==83L>8]TUaYcL&S]S.K#NOV^2S214K[d[/Ra@O2^K>(KU(KGC,_P
;)dS83LX62&1MK=QW)TU9bBS_HXA:M?eGAdL/.6Ed9JbJ0>Tc;9gD,e#)FeSK[ce
GG5>ZUS2\3f<C=,,D5L+6JE\+?;N50b6KA^7=/G>[U:/LWA9e4f;B\9V)JVUNFg2
_:0fUXgYLPU5bfQJf50]]2BKQNe&50O:?NRMN/0a[@^?6(=a4dB?(2/A460#/R0d
XT;-=RgaBVPc19J91K&?9</G=[[X>9/LHdTL1ec0+ecB+.&^<c(g;3?bd;S)[X?I
4:dgRfN[:Z3G0O4HQ]2Ga->3@(4]F76A7(+WZ+AX/aJA.NRPR<WdEUUUN7SQcEGg
9cecP2Q8gJC\0DQ)1&YbL,9E0S,Z10gfB@]K5_E1H<_cV)4TDNbL#E1XgeV>2T\a
L9CT4@/]URN=f^>-AYL>U;JecGG=aNb[).bS-ILL]RFXf4Ng^=6L,3:R_e&5<e+:
df6e>[bX.VTKa_acNW7^;:fJB:e=N#6LZ]Q_ddB4QR0@8DK_AN28EJUHOZ?2@9(8
.gVKM[\G@Ag,:6U]Q&JKggeOJg&_K^b:VA6W[R9,,4J6b1]QIC4E8&4[OcSD5dST
ZV)S1@@@/Xa6#HDa]a(d#4D271,0d=f^8e.H.QGbA;e@AIMN?C/MYfdY9&Y=Jd\3
R2J0#cSTfA<3OR.?QVE<\HeW)9S]+:6YONe5?@:XH0_JD1b3U+]BC?b5f>]c,Ig/
MOW:_>X)KP_M;f6e-DbGFOW#2gV;:A+g4QRWLf0;=27eJfNC2STW64L6GF[)g^1.
C7#XHKA/.2Te(^7S<^bUT>WAXP:G]8-f2b^;cKS0#21)9^S-^_U1/T5H^R8Qg7ON
M>92>ZJK?ScTHGWEAM/69g#WeXOOb3/V/V5L737F9R/6FV6B[a4Gec/T:AVOc0;0
?-[\b/fSSW3dW7P5<ODeQTBOaO)ab(A,KED.1N\44?g?/_Wf:V2(#U9FPXZGdYcT
1\NT?D7a&#;;?RWV#BO@gNLe-#K_e>I&ebVQ+@A(-W4fM&6GbK2B6/URD&gf+Of<
B8dM.Z38UUbc/FC3PIcAbHdRa5:e1Ab(f?5=AVFWLDd]KV(S[Q]8BFRcUD6:ZV9R
&CK7cW^.dPfgQ82EaD)9O;>P;F]P@cgI(F@+Z<f,O6E(ce0IBN8N3]eMd\&]0C_R
B?AK+E;>+Fbd#Uc3Q?8GXL:LFP2S>#ff;[[Q;0V)P/IHCKPB+dFdMBd35eM/46eX
0SIAfd\DGF@D?6Hd\e>\P+_H9fgB[7?N.dd4Q,\D<#I(#EGD,Q,EFO5VTL-G23+;
gS-7aQ56XX-T&6QQ3]7g&Me=Ga^e</B6Q:\,ad6H>BDC)V>5N\0:^8=KVNI2YM9F
LR\:ea,MHR3?LMcQfLIU<Q?;+M-BV5TaC#A9-&5@VCY4\O?\_U@E:_(FeWSY5,Y6
L[F&QOP^M<__ZHQ&V0JcUbb_K<DRX25J1ARD_M_#)(=(6?;9KK>MRaLQdde\\I/>
NNTP3(3^W63;AJHJ(cK:3/&T+A5LgK,aBV:V[YcG,VWX3^RB]TPT,K;BT.+7QCOV
>K^a2FQU8ZTO\c8Z8GIRGQ_[Z/\RVMH,@FNV_CNA^e.I4g((Rf1B)I\]\C1&M_/I
X5eZ-/O9@KW\>Ud4bA/\3dM,P#-(8bHfOb#93KQ[]47ZK24Ub;BP\&JDWO/Jd_Dd
N=&?C\,+ZB#dgRFb@1_/CERV<C(08Oc5,@I#_c,GE81QG.6d]Bd\g90J+g&5H9-g
HK<\+.2:-7&V>VQSWHITH;=]&2EC5P;1e_.HMHBB5WeP]+,R+B1_+:5>:YYP&eb^
T7H=56#DeRBT17B?/0;K\_+@^N6#G5DB--PX[7IB2D452C0^eD;))OMK[ZS>&J6V
+#L+==-^4QXM4^T;X3=aEV#[2]<D+&_EdO:.4SG6/[_bXB8(QCJTRe463:EcYH93
c&T7-TU#Mg79Q[U)96SZAG=]Z@L3S)YNBgEc_bG4D(?g_3Le)X+?@N62XfLbe\9b
AQ(0[0bA)aJQ-RFQM8#Ha#FS#eF:+HO,FcL:B5P_Z.51MLOU3aG0YGe:BZ[@&X:C
+(LTJbRG9fW\KP;+,5IaPF=>2Md(CdJYM/A8=-_92=][@SN@-L.8eO]f93A=)EVI
6RER:.SID)&MCb)+/COE+FFC#)O50Dfd4;e:)B,F[FD4aYaZQ5=Xf77?4X9GdJ\V
f]W>YAg-I;3gP/Rdd][^6=SI(1RYfI#)?V3;9d7F<H[Z9\C:Y=:?B>U(EZ3?L0YJ
>aT)+KT89K&:UHL>@5,Lc>L=e5+/_W9N2bJc5Y^OHUJ>NMX6[,]FF&@/;)U)II3&
JYM-RR[[(DX&JS@e=6-^IaFdJSNBVNYc8#B\gKUE);gb;bgYaEI6B=D#92@cC.d\
3T=F6cBUXGC8G,Lc.E>]]]4C6&@\]I[e0/Ke(,MS:>=cI/>G-,6L7KR<&b9M^4ZM
R=(/?\X5:4<ff?H6U+cCYgbA3PB-gY84;2;]PM\D[M]<9/MICUV8@O6VR2S3+=M@
ZI7A\7:Y/TCZL;4c.FJJB^,.IMX_NWdT-M2N)RLIJFDI0=PHJ/3Y43ALJ,N-0SB6
WC].1Q-<=T0g(RfRgW>d^PHW=G1FJ+R-fHDVUL4N@D;&Z-S9gDc1RNe?,Tb,_3YV
HMZ)D[N_9@FP^0_+I20Y[TD2TePO14)R58WELdaOEM)9D0=BeNMf>IQ4;KC3X-:P
GN/UYUH/<KVTFFO=Qf@WBU<L><@S_+d6JXba8RY?c^6@X70>/3-WO[881Jc\QI>;
5GN;Yb&]4/2WG_:[B:CKFJf(9?&)REOaRMN2IFK&Cf-QY>c.NU-=14;Bd[Pb;>M\
ED36BeSJF3^:MKd^\W@Bc+g18(0/GgR>gCSDf[+STT:=aK6TfG[[]]#8:)F]OS#:
KCMFHXY@_<NQ=[6JCB,GJU?1=^>OdQFZ(e)Fd/JIEQ#UO;86/cJ.bYQEJPdPY>UR
W=.OZgKV_;Y=+ZACKc6?5V0TI-gd4NHa5JYE2Z)5J^H<1?eHWfD<TbgL&^XG7C3N
N?4O<-#&=\JRAMd]Ya)PD7>\-gX3LJ=J9^02XRS(e#g9&KdXdGbZ:OC[IW9W,-N6
G>/6V0EI6&I[+a.);&ba>=0B=(NfUJ(5B[BU,YQ-eSP;eC2/a7L-P7FPLC_f9V-a
H(ZH&FBf/^T7Z)S4>J..&=<K(9(3++SSW2<7<_L<),CWg2E&R?BDdNe=EIP^X0?(
MD7[(9/>7c/da5+HGf@4VNJCb9-C3)b+0Xbd\JY?@V0^S_.AQ/7XS71E+/[,ef-;
EcU970-[;]Y#2L;B^_2:O8P<E#ebUUfb+036K-H8A2b(F(LBX\RTbcK0O&>WFd>^
Yf^M,O\aQ&ZB4PX4dSZA@O6d/L.@XeF8^J?I7^1eI:_S@CTY#6HL8Z1[?^K5cRD9
aV3cQ1[::4O]>-X7+CBNV/(Q1:HK#/P0QOH+45_I-6?T&/KYdA3PdK&f]CCN<0PZ
G7cY3GL<f^,9Me:QTc+P<eZ[^/E)8H&QGOfS7dF,;:ZU;L_bfGLTW)9.V7:V;V:g
,EPVI?MSP+CY-7b#d>ba@R?]TGbbcCV(-F.fR^<;3?8\JS=ILf<g/;02L^3_;M;/
QdW)DX>[ET>e=D.FdIWD833LZ>^[4fXFg@/:QN9FOGZg/<SUa9B[[,VFcb4)bC:X
Z>Q9Q#F@>E0-0aQG<SD=+c.4#XHT;#b9TWCT=,X@U5AF23;bNO^eRX[2R7XWaB;D
LB^49BBYb?<:d\#S@406#.+C,3.#R)\8[FDf2ZPLVA<]c#cb5Q<W1[N@PIE2B;AH
bO1GDUdI)IN2<.eJ^E7L6J]L(<^NAOL/;)F2]9E48^XBXVKC\@7/EC(AOeR?U=CS
6^@,HDAFc>0=E@&7\5Lg+-PcIE5L_VFIM02gU#gf([49D<,dI2Y507RCMU.+N+U4
BT-4Q4IDA)-&(La.N.V=gVA1?c@IFDa1[J8bBXaBePgb:@P@1FXH5&FEK0<[@^1R
Z(Cd1HRP^V2J/>=[U=_9?&#V:C>V6YVRT3U=QTfZJ@PdZ07A7#85d#TbU5a5&K&Z
LMd/G,Hc]GaK[aD9J(_DbHeS[;a-=G]Y\<W_?1TfCVF.)=<Y_O]a+]8RL.@P@,_F
KQR_JQEgKCO;ddcQT=_MP-f<cgc1AJR?H1U=UX<cC#\[a-1>)2LeD.-Tga>@90)0
)b:#=#d4-6_.#E6=Wc_ePfB.X;8Md7Z?@SRC,@M&#QLBR[Y^BPILO_#Y(8)]K+_5
[1N4SK:d^&O3X&@0U/VNC1KeU;c6MN-G6),#>b>=\IgE\-9,^HU6fLg3FSeJ^33-
H;FSW,cV[K=.4X^_4>)ETf.A6fCIe1f\G#Mg<3:A8)IK>3ZXO-&TeXR7BMZY\+15
N;Q?[(ebPC\DRT[7;J2^]@PQD0@+Cd2)cgIPFWaGN21ZQ&Y&13[?FSQ/KW#ZcROf
dK5Ub7.1B,cPfD2J2;#MV3F#B>DeUFX^CPAgCV;C[;4N[]5g=->J=BJO6Z[QH\UC
V-39-NBeJ2PN4,IFXFQ<)F/_D0gD6>Ra0g_P<>M7#@>E-JTQ&:-/<T+aE>4.f1/H
LdJbTDa@8<DU1WVS-->9P8eC4>AI39.)gS9]P>>4QNg2<bcEXB+LYVG>,^JB,3(^
R7:0;GH=@9]UA(g,JYA-@YJR0)AD:HR&Xg0YKX3)eJ)Y,d+MTdFP=@cU(5,[3@@,
]cc2H38?7:1?dWC)-#d=&/BAdSg9O,0eJ&0RE9M<[5(aH(Yg?WYH/G<Mb(W6Q\:M
Zd=BHZAEX4K9D?B;S)U[[(\5Y^2bL;6P)TVU9GIfd\SR80+6gddRd,C>I]J,Gbf]
5<5TD#g>)eA1WBPN/HBP[?>@ZE&GJd=OX4d+3_,<5CV\?<7\NX#d_^T0XQbcELUL
=R?2]9c-06\BY1JM9+MJV);CI7LX(@cR^E:?:RVeT+g^YZeJSLQ9Y@cFN3aCb+)(
N^JP954gUd^0.NCJIB@)V;4(^PNRAOe=F_SE=SJUOUV_)3-UQ5H;SZcJM\BgFHUS
.>;6])NG2ZRU809##29AS6WMSe8XKJ;(?0#g-U^_dYYY:^;KX[A74BZ.NUO\_537
cW8Q;f\fd9]R@)QKa3I<WX+<3bM^/A[2V:;+6V.VHO3aBH2EcKKSVbc\c+];<@AD
=3M9UCH_HfBI(VG,8WbM8DTTAcNSQ&IAGYVc(-^c_N;7MdVg>=BLL^a:cFD_1RRK
4?DR^_<eQ2EY^XJc7528^(@-XTD8TVQg&cM\.#/XPH#BYgb>FHK]dQNS_]^U@Q#)
=Nb.Q_J]R[QXTRH#R197#+1\W;;4I)S+._YEC<EG[T[2(N4dNC.V4e@ZXEbN)5Kf
+VTO228dO^Z=#<;=[/ITeOA+>UA>2D6>((?5,^a<d[6W@0O<d:f_Q,X?fc,9J>1S
GVZH&YAT>B4[-UR;X=:0VJN0P/3HJFa^<1Ue,W<A<FZWDHBA^(06_+UX[SOQBC5;
WK92FJUfgO3U2N@)6aIM;+c@2R&-HQAfMd&CZd]R)FV[^)OZT265ZB42N_A#C2QW
DFD_YBB[f6&2R?d8&gdcWaE=Ke;MA@<1=O\aH=JPL8Qb(I8<cT.I^)2YL93N13YP
g&272=-_(P:ULX4U^Y0:I\@;?Wg8A3;T:gdg74Wc@Kb89OF3/KN#ZgKb[ED]fa=Z
Z2WQA08=]\.//Z;YH>;DSVI8/8NQ)8K/PF]fY&NWK<e,Rf36gI[&1QG0&IIdH]><
Eb#].X9GO#g9:T1UU#0J&U1NL2X55-d1<.&bW>IG]MeZ><#ddd]&5G5]bU:Lb[T/
#OW9N3[(1cDI30-[.(XQZQ/7J0OW95EB_9M8A(^.fOA,X,J20HQ_&KJ-PZ3M--c;
]Y]-E<^IF5M2@&-4U8BQUA9fa5K&MaN1Vb=AP&=K;OIHEbIT^HUN8/#-)X66-Z4\
PF\]E25]2]OA/gPI_QcSK9bS)e::JKK^HS@LLB2Z;E3I?HXCcQe/g4c7N38\/dJL
_#QQEA-[?,?3V[[)9RBOFI;<NQ;C9R]]1#.B_VX>bOAQ1\21K8,W+:g>JUYDD+VX
6WHQG<_Q&:T3_]\,Pg)E8e1M\F7+#+6>0c=5dXcQJg^?MZ@YER^;gdIZ5Hf/&/J6
cgIHC3(aVcaLX-#R#E]/JYX9E&0LS8+OPC@+RHM(^;1Fd@UA_O8IdQI/MVV_,I@]
.S0ZCd2>3E)#:S/SBHSU3NM(^B2ML0bYP/I,9F02#gWT_S=_TLAdEEACYe_Vg4?f
_L9gG9d15aY]PYD_HA826&)MdPCc^<D+^/IMJH-AE2G=8aN@WN&A/[]GVO8.Ka(9
G^]F<P.-#MKHAb?CK9dSZ=ZaO.^c]b?\)L9?c5?@)1KSPOcCG=c;X5^&F5NIDIYf
?\HIT^2CeGMR4d/Kg[=c@PJeL8c:NB[](,?)TB7,7)B^([/1FL>aeac.H0)3c55Y
-]d@A674OD2GV@O@BP@^0dg?8627.S^9aaD;I0e(dJT3HD0+4Y_g/]SHeIMUVB45
JL,:SB]VP.>Z@KQ:J.S7UKQIJK7^\;AOKe\ce/d,?:3PU#9J#EQ3&1:#UgcVIK[e
?;7eaC.3gA@4TfbYPe_W4FcUa;BZ9_ODR<<4\eF?4;Fa=CF54]&IX#90eJM=G>X&
<]R^,+;W23Y?P<bM7]TFX,9]4GaDb-OH0QB-fZ;LSN/WA[QG5g)GeW8fR7a:VS-]
[B<HZ/[35e(a<KE);7_Yd3HdQF\6FRcM\CO]202JAgEN;^_G59EeS3KOTIE6ZEe8
WgHGOE)c8:bcMYK\W7V)[0<X@AWB8[N_\J1QCN3)>PBH,GYI]P>SFO2QEb&e_d/7
gY([]RO5H6Fa:26KIC5?W_TK6f:e98OgD;DJKDN<:?BP16Q>c:9TO4V;SfMT1RDU
WXKP]^bI4,B:B==\:6O07CZ^LcYR4-ILXHaCWAa\5R&0D,A:XG[04E[C]g,]6F(Z
8RWT0=PdG-G,O7?HI#-8ML_ZSSZ0d9gP>(M=Q^BDe3LD^R?(\=\b9_Af2dT_>D+M
aZ=5UBX,/H=S]aX&-WS\WfJ13YDDY3[C:V]+Q82>>g4=E:S;1):^ZII,&3U30a,0
9\Gd=6dM-FEYRLI[f#>CCM+.5+:Ab#3P276]_?(.0[G,,5NC#eSGO-e]J]c#cMY6
<a3V==J[(#gMGGZL9?dC@#=JUSED@47#V?;>?bVOGHb6POPH;e=V)I4gF5,1:35L
G8Sd<_F;_71+^J-/QWI0dV5VR8?0N(#dPQ0(,YV9B\fB\+M:&baXJJ,6aXY6c6(Q
WREP+0,8QZZF]c\>LLDbfTA&6MRWEONY3T+_K<IBG@MJ8Q;\K>LUL]MXe/>9G78F
>;a8cJf;e?E1\;1;IBZbI720-XO#eJKF#?OgRCfCMSI6CT6b=_&45X;M8K/6N^[,
.(;.Sg=#?bADDFf?&7T8e/KZc.]?7cUJPM>#UaOfIRB?Z9P+gY1>Q5PS[U]Kf]UL
<.NRW;RPbaRSgT9=XWF[cTM](PFcV+#c8\e/I9TMML?GaW]E0X\2cN:33162@)e;
B+R[a\[fYWP>ER4e[F(<;\L4fX;_P,&gIK(KXPGL@S2O5?]R.UbD:^F+?+27?>b+
K\.:&,>#0[F(D#A2.S_BPGPCT&gPb9OIf@M54?4B78MDG#T335=Q@Mb@a><4LV3b
3P.VbHCCD///7Sfb+WaVZY)1d,;_b=-D#1RL+QW#:\<-?KEXf4&4dc\9,LQD^=.6
V=^2DV;Z^GEMQ289>?&F:OJdAKf;_f2^&g/c:TSebcG0(G9O\-)](->QcS]/fa_?
HK:<b;)H302C5a8EFC)K\Z&X2Q?8gK7OLFDH_:1,dQSdL3.Ne]fR26g3[.>KaV;+
YV(;GQP4bLJ/cOL7UYd;Q)d]CQGF:ZUY]/&)9VS^7LW5]60XSXT91(VgU_MC,-@e
1;Z2X\2_J[7S39FXRX5TGgfUQgNQ\S[.(SCeLOMEB5^/+cd+Sb[@fPWK3547XUI\
ND4fHPY)#N;F(X6G0Q2-A.6N<3/]S,_3[6Oa:4,gE>:#9fb_>ec,.aU#(VcGg8EP
e1YRe9GAa\\:U^D/<BIVD45?W0EI.6=/@J4?9G_Da/gLSFW/@CgS<K.3<^@U/DOV
V4W038e3KDKgE32)^9E>\RP-ZB.9VDWD7U6QJgK)ZC8.N<,YF.QEVQ6,K<)\]:CY
53#5Xg@B(7X]E.>VLXT1#T6+&<+LWLWQ?c6X+IQSF\X/7+A>dX4Bf.AZW4FU8A7e
1XSFA/\0/5-??&;S;N<&e+BF_KROMb2U\?9DAQ0d6Y[(O>MK4L5R70>bKW4QBC\^
DDE95;1UfST0d@Ncfd<3<O?3PL&a1VHaK+eLM^d8fP^..H]EG?Tb(SM=X)6fJ)/g
6&??WOfbA2X&S;)-D22<)AW(YR3RWLOAeBIVPQL=5QgCE92FM8H\RY1+@f.LSY(0
2T20,HZ;]Q3(eA:UMf2;I/3dfRT?=J[Y0#e)aB1U_6:]fPY\#b;-+:XZS5)3SCFF
W^aFJS3T02]Y6HIBgaeXOfU6Ga,J[0(_U<@\2;&X7UM^7Z9WM:Z,K6afa,=C\Q3G
V<(P7X]#AdE&(.Vb:^_1GD#/YFd5=Zf.L:)-R/O/.:D;^Rb>)S,=/[#YA.e.eB6F
DOKQ]B&;T4_BE.a0I9&c]M;/+Zb0M[2RDe5)?_[-&MJ5dSE46.((V_&1eHfW;LDb
RA_d&fP65Wfa7#b&7f\HM(TA@VXIM]c^<(XMB&4J47d_C>SPS&LD6PQD4gDJVGdW
e5G-BEAVO]G0Fc6Q^>a2EW2X5KG-GbV]ZG\I:_F4\-_<R;77]gg,7;2a(gLVA;D#
OCN,4dTAAOUbd)HLKfa\1FIa#U\a?&05=./^132UWO54XV86c\M2&2LYTIN2U9#4
EV=JKT65M#R6.9-ATZ1F68KC#SeX4E>aDN2?R>>,=Q1[XW?&HJVQ;a>6L_5W-GA]
5J>&SZ\HOU_^N@GQ)6SH@]45A]-(C4W?<?D127JXWf^B7A=<X.3JL0-)P[S6TNY6
PU4&e2?A)KVU4WfU\W5==@ef[Bf9P1]+c71f)9C,1_2]#TC+Q\T8dK^I?_=aNcSf
5aaeM.L5@)ZY:YS0/+4D41&Q=P_Mf//96]TR?^MDSOM(ZM=R_BJ3c0E1O&]2<aQ6
=P_4b=YS:?(Za2HQ/O:)DN87)J7G&UHe>78RVd8L89P76.VH>48[S2JPFD=]D.=5
C&)JXWEI6T-DDdAC^^Fg&9<Deb\2ZAH1_^24K,e=D2J,1#^15;3-H))\(:U,aJ?<
3dE)D(@(>ZS2U&+Hc-I94W9F6NbUXH.d1ZYb?ZM7^B(7a>DC5O^cSBeT_O<A?S,M
dXIGM/1TeO-\NC]9WGEQW=_+VY1G(.:U&f5&U<dWWfF8&D9V+J#RO9a]?Q4DK7Ze
^9#\0#,?&[W0CPf]&EXRa27ccQ-TI#8U^fA.4&TfR8c2)@L(V7/^]2MFH;18GK9V
<4,(@c8-DKA@Y6QC2U\[[Z/#>@520&G5/>RZX4@^cbZ]#3]f;?cU,0>Oa^JcXbPV
C_@Z_>=F)<d?/YRN>+.9)5Z97W\RA\[A;.\6(JI6bPH2SF0ZRa\MF2K&\UBMN)N[
.IWR0TLX98SeM8<<UG\DR]B&P<N>VD<(08,:TK-HI-=_.19S7)I55-ZOXg#55.\7
NE)44Z?=+\=<=>A2d;.M(W6++W#4W9/2<;7>I685@2+DKGYR7dQ7X</GH_,1W60(
Q_M67Mb2Z8>3\@T]/V^:5K0Ye\>&GVcKPbY8<PPAYdRG&FS[D2621b6)SeZ(BaLN
UX1Y(aTcZ6F0bRQPKSA=0(4NCB1(e\G3M)dWA16B9EV0I2;KKIS&SRM]aV=TBDZS
DHf_0IE&b4(b+4XO/>PEFS4L38Bec66dWIB/I_fY5QU[Bg3:L7KN/+47N0dX,U9]
866^aP\]\-U(+dC658+YPL]#[G:gS/eZ1F^YF6c-+A0/eY2?0?f@S(F_>E?A&<EW
3/E5B,(81+GNL[;BgLH#dJUF1_Re]C[:;K5CXYdH#PL5FF&UM1F50Q.98N[cQ_IQ
RN)@:^a9PV#Y,YPd0[9/4-Z^_MIPU?VM;>X3cF6?.7?cPBX\N:,g>.f+8U-_ZKYD
:bM[Ca,Tc&/e?N\Ef,E>7K78#.OBN4=SY==eS/C.e#2I,bC4-_CGRF:=EBe\4NH6
];H<<A7f[A+_@=EJ3>_C\c0f+HEMIYT-f]D^BJbX#W_,WQY(1=V?DR5I@+aeWZQa
H+F4S#Q/XC(#>/@L)3c94M5[M8;cM4S&8<<Cd/9=RGfO@G&BfgI>V7JCQ[YSXee)
a(ZFTF)UZe2E,,-E<Z+UEO/N7H+=,#W]7QO+2[f501HO]dH[>#HCQ21b\9ZVRX<I
WRNZPMaBO>R2^e=00:U[Ndde,4.]Z=_4ZTUXP3,LS4R3CZ7Y.DRb6WYO4IOE(6H[
(75>-=;>G.NMb#4FY\\4YWf_b+)=V@U:d-@M@];FWaA1YG&NC;-LPH^GdBC:RWF>
bG?,2]J;-e[XE,0]fU:>I:BB;B-0E)T/IS>PU(]&R]eTCS)27G+cX:IX+?\YIb[#
?gcW780P/5#^SMc.)]7KB]E55I?HBeLY-(ZQGgb.HAaRfBV+2;WH6KT@bKJYXH)>
]I7EM)],E81ZCaDD+@./]beab_T/;>CeaAQ;D>9=-0Y0CUE:e([[.R,AW9f3HGLM
D2L>aO2\8GT+B,TTG0e&2ZZTR5252_)CUPIE45d3FF0,1W>Z,]_5dJTdgULOV4cA
L,S9LEXbZY43FBNE2NS:_09-Pd;35V5&DFZ3fTG4[DBeTIA8e;GXE0K<2B+XOQ-J
-_W>9^<??]/=<-dD^T#ZOBYSe[-=GAN8R4DJFR\0L,E1TL,VW1IB2_2R28TX@YU8
9ZC0^Pe[2-gDbLW8Vc+;@-85b-3CRCg#0P8g;H4TCMRPcY[H=^gQGeD?/8D05-:(
3]94;AO8gdSC5cFU2HVAG1\a&H[^A:V4ZC,J^MRNcfODJ80#Q)1_PgNB>I.I8GLX
?a;E#]Wa+gIN9RPQ3UQ#6\6b+T;^/3F#205#9855V&+Nf\C++,)DK_Bb7.eQN8(U
^[d:POb9W)7I[b4b8VO0Q;9Bg8OR6d^TZM;9D:BgI,Dfg5,Gc1]YT?4W,8d7U.dI
L8d7=bg\@<?1Mb#Q\38D(5IS2?68W6<dY_,Q#)?]T,[[8?^+e;S44W[#F)S5(fJ<
dg?R>.2A+U+c0J6SA>Se+4IG/N4#^OW/QEYMCRQ&JI\)3B:;LQMHX-V,Z&?4,Y?2
>]9E[A2;g&TcIR0O<]29>.[B;Wbb7J(]1L?P_9ggA>c/d[7E2PMF8.\S:&E\Ve,U
#-&E=Tc@;];[)>eAWRWX?<]@?f4MML2&?IAEPY8BWdUPY\6bIULK&+g)I<Me=bLB
99c06Ve+5)K-B,8ASV5#\7fEN>))P33R+AA^0=1YECeEVCR#M#KW&:TNY39+&Rd>
dIT6,R9#5ANU-;QA21IJXGa^BgV+fT#_ad=16-ULKGA8J4W6ZJ3).4;JT4YZL@:&
a\)3N/.WC)fO]/0FW7J)LR#b/(J,IZTe&_R@Y5<A+=_YXZZ:+7:=OS1,V_#,KV?8
eI#Xa[bW-9<9?c5=NYaX=]I@U:K_\Y?(5=^>0)0gTT9P/R9BXL19K7FO]f?6^]Ja
92B_33;1+II?B-0^154CO&\UbOB\?KUDKAfeZ?ZPR\;#>B86e>U<4OE]]T08FfRb
EeFb[:AIGZQKUQSJL&6U;5efAV0HI6NO-dG+8.ST4K,eXQ?IX9b+(0EeA[6Y0YL#
O0^F(_.gD>NKRXN7W.VX\Q(HUe=SG[F)BC@c^O8EDX#;^U@gf25(Hg-6_Q<USIN[
1:>YF[a952-[@B3YB-ER,4gB97cUZW).c(X8R9efK-dJD)+O\SDI,YU0&]Ze(2F_
@A#OHbT=@U<+F9V<QI_U<CE3^4+,LJDDgP=LOJ;AJea<Q9FU&YBO3g5:g3L<]fg-
CK3K_edG53(9f1B(NW_>]<DQ&GM.]\Md+YX>#++T)T1KaTKO<8eXefB+ZJ]TVU_G
/OV2D7L.LU.),J1>b-#(FR7U\UBQ76++H_-e;_Ac/JG&)G9@P_)@M)9J.3L@(-/#
KTNCPH1B50##)-<1LeZ.KO/^EG@@QY?>0+#>dO16,7&7>Mf7Z5EY]23+#9X\0&,(
NQ5_4[T4\3:\.eH^UNNKHDL-WBPQ^#,H[/6,N85&USVL/FR+=&?5-(P73H,ITW>G
LIGcG@]?cXdW75&]TW(H+Y_@OE79MQe)g>HGA>&=<S1Y+65Qa0)SC=?RR<9aM^O\
0A7<A:b]]1E[+TJ[18X1TB8H_g]JYJW3,T@J2E;e18[0:JdA&OPSNDOF,\M\L<(E
(V;SA^:>):5F+>.&c3BbJ8K=dN=KN9:7/3?baY7;LZ[L8/Ud9H+W,H09YD?e2EB7
V_KF1?)]V83@3M2O.A8/4DJTB/:(Q5<T>&>d,QZ<->7:.b,5a<[:JP\(D>@HfYSg
J]eK=BB8<c-Z:<C]:>60P4fQDUC4GM79K&ZQ^:X:g<:^,VS>VEEYJa]@Wg=.\LL)
aI7XKgDEG77Z\40SV-AAJ6O@(_RF[a0_]_#fO\=7TDOY]cc;c]G1OZ3./JI74G,;
6_R]f@(08a#6MUZ+S/RbdS.fLK7MHMG[-a.V)@LX3,f1aIM3C@V7OgLaA\J4b3&Q
[fVDVVM\Z?95J=?ab+D.>;_8RW+6Gb\g&8+VF8]\;XK)6B:=F=,bba_S_R^:eG3A
-S#H:ZORSZ^d.;147R,;/I:C,VP9(;0eC^XD?=\(RL>+M\K\Ob@6Y:c:.]BIg#fS
I6.+VB2XV)WcXe<:2?-<YU3V2bHST>N4V+/N+eNK.<>]U5/8M<^Cb+JU)gIG_I[a
Fd=[-R4Qe.9UW_5[5,A03&=>(ANQ3\955NFIf6OO0.<=+-[cJKO[_VR]&)7d4K@V
:KDg^R6>S>6XN1?4.UUY<]_d]\M2P[>GY#803CMIE3.Ece=_-;a9Fc/3U(I:6]XI
7a98WRGI.[H&5ASH#KYXec74V++b38dUTT6^b:]g&[]?G?adEfG86XA::-EWJUZI
XRJ6U0TIVU&A^:A,GI)adG5L(@_Z>34\GXHa7#Dc[QV#VaM1B(M^ZbXKZ]9bG:O.
ba-2(9;P6SW@&O;4A>cZZ[A>66@G+\JPZEFS7MgS[1]?1FR(7)gTf)(AT<:0JASN
1WZ/L67IDO3B-3L)&I;H06c[0#.H=DIANPHSGZR\_>I;SfH=&H14@/^/##11^A,\
d)C2A@Y_)F+&5^#:4U7KM-5#E)DCQ1d4P2>8(/<7LKFBPf>NM:@61Oa)P;@29L32
ME?ZSF_cP(EY\dC73///IV59B@VdWaONCC3a/bZEQQH;;1[X=?=+)5]K6YG6A@TN
?]5GW2=G?7Vc3EE[dRGZ,.QeVG]&G)DFOGcD>1738/_9gBRFO##Zc9WW0b-_HT=M
P9UC,be=87\H[N6g>9cgNHG=R\Oe4Q]8>TMHR(Ec]T)A30gVVWW9I(5&)1aTP:JP
H_DS8&MEEcJFW=;@R#/086P_T[a<+<Ma+7UUBL->60B#\aS&>GReB4S[9KV/L=P&
?H<<D4<Z?B@b91H:0(ZDUAfSe5I_VBdBeaH&<BAN7(#OV3Q:CY9AY<\cC;Sbb@;1
#CG.<WY(P4e7cQ/ZVF_+CU]YWQ?IWC.,EB/@B/Bbc_39VVcD[#DF&CQN50_GRV@3
5EJ?B[f\@JM1,DKF5L7c+Ka@eMN;69:;38ID5&5(6L+:&B^9Z[f9b0:BH3VV(V8P
JgW4TO[WVCE=RV]Y_F&4.RKbD/S7L89e;6c4bUGBI?]Hc8=CAZ]EBS2F9S?)&g2.
3C+1LL4::#TWWA=X.9:^<UX;2#CJ-8g+b2W>JAWU9?V4(C<:<YH+R_@JIa\gccT<
-0NCDV&bdGe;d(OEXWf5WCM:?I<TZ4/N<^1EQ.UHL1=C9](DZeJ^LQ+NMPH&Lf3Z
Gg?9)1:&31?a5ga#S@6JZ3ED=;d:MXKO94X,GQ+J)fTfVX[GEB-G1#_JM/6S2;cU
E\L@)SG).VJ,OBf:E,Dc<-g4+Z<5(Q3f\bQO70?U:c7--N6bO.YL6>A_C,]d=fKV
A7DGPR4MAKNLR;>]63Y;P470I9a&OVB/.>L@KVUQ&6DCYK^4&f.1&<-ZHQHWS.fZ
b<9c(/FW,c-I3+ag2[AUHd^CQ@ERWR@E7J-SQWL;8R//.fXGD5b6?4,G_Ff.DWNP
Q^C/TaO+HFU:A<G:)GQP@[C]<RZHZ\GK:Z)AFMJR[^3NTG5[FKICKK?>L<^IUV1-
;a>WX>TS2L9]Uc@O,/B<FGH)77eB)W8P])E/&U7<9Z-HB-L92NR7(Id:gFXEV3Wb
dUB-.>J4YZAc^8bQ#=\f]ER6FXI6&@OJZG9<MO1]KKY<]-,B,]aA1=V8>U?O-2CG
LeV_##OXX])W]f+De87g,)_:UB,O:d<e5]H=7,Z>U0YX,DW/aB-.]fW^JD8;G3=8
Je?+>^0e](WF,U[)2a<;Q;3I?54&EY8<fd.RZT-2R^):HGg#1GCCHUGKNeN#+9^K
1.KdGNB6TMd5V+)=f-\PI+I2#7:>U#Cd>f\dS,,gI/Rbb^d+:C>WA)L9-A.QX=GK
RW]?\f9/ROIK[-8HVQddNW,EL5&(b&,@e:=L-HX5&edaJ5H0eW;e(HIHJ8dHWg:V
L7V^XGYW40J^^9[R0_2+e0(66:@BQ^;Q@^C[]8HL\2>V?SS[L-S4Y)9-JM6Q7aY?
De&WF4)7&g.5Eg,B)=2.eGWbK46E)XC78+:JHKGG9)_5f:P_W7]G?Ig,II.4[T5<
9+g]^S]ADW7=+WHZ02]fL19CQI2J#N+8[A5>0\=d)56+4_dHPODb+A0=(KM^C+57
IYN0FCJ1/V,EJ@Pd5U&SVH[.TN5dZJfFFW[BXG]&/GWZaKXY@\_UP3P[&/UCTAc<
FV1aT-LU]JGL7(QMcfB:L?7;G,.G=bXVHFO6b01W]PGG<_LSAK3>511e(@^I5N9b
\d.TSgP^R@)Ad_a?UQ4C<C\.0^1Se+f;:M:;+@C&@J@FHI).fD@I??<-<cVa,R[A
#4B/PXD<ZIY4,J=9=fYgYOP?X@JYS=;,=X@1;PM=R0NeD_:eN0E?;dXPY01#c;.S
&[_K>OG\d>3W8DNdI#J8eL2aP+d4&]B+MEBQ@^OSB)V?2cHP0-<[CFc;HGEH=ReY
d#7Tb9K8,UJJaR^:\GY)F:>dCCe#6N_;NR(aKXf=_XaB(^#N5DZHX;ZHU4)<K(b6
B66b.YY^.6fTeP,G96T[3JE/UR2Ke[-.N2F@IZda=XW9:JXWIJ:[a/I1&B2/5<#+
aX@XZC<^0M7b?);E\3[QHFO0Vcb^\30@U&VN0O.9aGf2W<)(B>A+D5.Vb\(8JS5f
b34D2(N(X>UR43_f3Z_HQDA]-5\TJX(]dHf&a-#Oe-a;FM+KA\#9)Z/\geH9>+^N
T4)Q>@_f^5)eZ1BX.ae5#M#B6Q(IB@Abg:WJUBLIbGX#VQA;0,b>NZ^A2NDHOO,&
G/9G-ggDZe-B=XecP2b156PU?L+QHR>&&VU]=OCcFe1+B;RC.(3EPB08AF53Y)J9
>9_HOC^,_0VO_CJ#(-N:G<R72:3-CH:2@4LE4C(L33KS:bF^.#bZL+(gdP><=0\Q
5e_P+AMH5,SVN(M_XR\\S8NGT8I&c9,^1=9gQ&P)gUNQaIK5(+F-bc7EDc8(/?-A
T@+V<-d(ee,C7)2R#S6g?0&>=O.U.H^&2G6-d;-0[)Q8;:KW7MQW;Z7;U#AP0Ybd
S.DS,&1+4f[:fbZNP2[dbfXKB5<\\=EX7B/e(dQY-UMHQ=WD05K2^BDe<cKL[QN=
+YeZ=bL;)(KH47NHL6aTcdY6J6=g-Ke:1g9NI=Nfb;,BXC.1EU)JJQEK-G+<9Vdc
_F-J?HbGE1,fB]gE))\cF.HP652(ULAXHBN=G78>[ZB#LGR&3:)\-T?W<VN<5&S>
?\2c2VP8+P&R7cW,1X?Y(Jb^dfUY+\VY(])7VE\f(G8eW^b[_A0JIJPC?R/BG64D
W8+GN0;ERJfWP=Id,A2YX@3<9QEL4U<\]M(:DRfUWA1#PI17JLOTV(=^FTQV#,5,
TaS#1fK<22\U#K.^\ZLR&M4;TKRL=0?6eXR:aI5Q1CM=e2K#:=a^>U&eMORQA-KJ
FY3ePGTBQ;T-Y--SIG+4Z],TNWIf9>@fBUY[^,1bdb9ZXWT,bO7&PgD^aRHSN\#E
TEVFI\#eb&8UK2GQU38GL+SFMG)X4I4XW?&V(Q.]K3WX>c7<2_O6B2I(5HcK)dKb
e[E)We#IE^;g<OD_7J9=6&[T8@9:]_bQ#K@MP>T/C/2J-[1e<>._2@NXRSD)5[5B
)=d<ZG3+CJU1L0D>U5ES]#0[fS9eEU5Qb=O9V39,QW^DTgM;ZB2K-&[RI1#@aXID
b]cN&^C]G.Yc]]?W?@7J;R?N(J>38>56/Y7H,C]g2VZFOg^R]OO#\,PLQVWg_44-
(&>VgMdH<+HI6V)UJ:+K?^UdYbN?AMfU8QO(XN8T9eOE6F3O8He&<I#R23H,;=U+
HTPI2,8(24[#G(8g,AZ7cBeR/[&8RR=PeX;]Y>#/SC6^5@(BM@PYXD#B(O)XaNK.
GFV&T;LDGOJ]Q=-95IMIP4c>F-WcEW01#_D\Dg+1X2;SaZ(Tf3/.Y:5S\E0A#O-f
J@(V2gWMGfUR.[eQDX#1_1fLYA,/\?ZT/DOV7:PKK0)S1gR0E6BdNObga6d<-5XA
^77;cg:?G@7g8ZD[f(cZ5UR3)4KcKT&B;eb+SaX)]C=9R/CQ/f&OQ(0JRdMP=USV
=Fg@BK/S7/+(3I9GLg6)\IXA0NXF&F6U8b)C@JDcEg/+e;^E8aKB9d)^5YVA3(?L
&OID.ER+<W\<4AJN1XU2>(5#P:@)aaW.>ULU0EQ@:.M(YSMQ,8^H3T>8gX37\Q6,
cUf8V_R^LSBY4S2;gU&I0.K?^2eL;SUDbQ]N9C^^-;035ZGE,U@Q#W_L=21VSL,5
Q3,^\<R8=e>^RcISM(^2G4>Q&[\.&W8P/QgM?\B,>X1BXTdZ7?GO#gR7A3GFY/YK
N&PBPY/S19)-7e(LL9HFA(Cf+\H#=6;HVD;C2f/;?+S84H+O<Yg:1<Re)gW)RVCD
]<S88\,B]aL]@>a.XgQ#JEPD:YWe@C#)ZeT0_&[g].5-Z,>G(W)<KE727Eg:cNb.
6R;dJ::,@-WSCYR&J\KDH&<TG@+H:8(#3]Mc<W9DOJW#7aF2e3E:6^(Yb:F<+5P4
2V#_(11&4N\1:\dZb&\=\(A,1\A/07H>G9ZfS4<Y(acYFb17G8,G>dDgC[g^DA((
)OR:\RMM+aJ6YVe^\+JUQP+?e^1&:VMJ(Z;X]-:UCbcPOZORL4U2:J=^6)ffGGO-
3#<GZB&+SEdN(gX=DKN1U+=S[CdJO<UW+B:cBQWJU)aI]96H>FF948Ea^]3@T2CX
g(DO@4I5WfG0dTZaLM;gULd4VZT8MTW^)_7V+M<IXW7OGX/))Gc4W7SZIPbA&C5O
(:RN/bLALAPd5XN>A#YgRGQ(X04JH>=gRa)7A(A^J03c#.EVGPLN:I;7Y?QRaD7\
_I#9/^8S?L#NPOO9EP3>Fb-[1XC<KgQLM2]D1&N,4Z,8Y-M;]BbOK95bS.]Q<[9Y
e>X:-^a@3.L^3)VFSgfNG&4?ODVCc?]dBdCY=-21g0?</#H==>\J.1W,e=MUbA4L
@.9H0P5RGUO9eIAY8W7#dC#L:Q1J1Q1ZLN;#8,@5d[SCBL[@C2#SWa>6&D9W3PL<
AAU.gSc7Z0>gL[<1\XK>c-45I?6<Q?ZfE,H#@#WWW-3>EN)FfYbb]H]gBW_#e[9F
Q,S#D7\9[Bc2gU13BQEPd1=0W_WYIbV3F7dFBV9Ic,gJ=HZ(A5@TM7SKcSg,ZD]<
43Y\;A?c=g=GP,;&?^TVe^^cgR4FBdbLRc3]>>-XZRV\Z1[d9(;J1dQd/\C_LcQ]
&=gN;WY-T,4825P<g0JN,bagG1+I9K8aN7aHO758(^?YFeLM841<,g47dd@:JN@E
&U]>Uc=US>02R1C9b<g>Y-)b)[8F#3Jc<:54YT]:Q4-J6WQ&CHg<CKBc8@NZR@U8
cO78A/0M(dGO7-,2d)6eE#)V&aL7KH]1\BN]>.=>GaPd^@ca6\aLBB(9(OM(,2Ta
<NJ,M5^T9Z&g_dY+ZeT3TU<e3FN?[:K9a)AG/[O,+)YO@YCCU>ef+LUY6#Bfe_=L
E;TFEMEFB.L>V0Z/5K^B3GD0K&I>XIT[P-R^?3-N(>AWI/<4[aYS1)=c&D/(:F2I
R6(5@J#.B+_14GcN<U7ZTdedUAS?SC-??D8>0F49#cFP\M_-FV<B6(T4F8bO_b3F
&5<eb)CFdLZU>IVdWc2A_F2fc,:Lgd9\T+CR#T5/M1H43PP&]>W1ADP0IWTgJQNc
HcK-\^AR4D4B]O;5REW8eJLZ-c.S/.=GP]]4\B@X>PeG8-F.F6&45@1TW2]1CS4J
(e5X&?6_[J3D[G<\R_FN<G:SX<4\a<CDICIUPbLG(Cae8B::e,]?0?GS,cVKRLAN
CbOU_/@L^HSGP0RcbId@?4_+,fHXDEFAK&.=C.9@gB_cfKD8U<NbW0>PM_6V-SJe
#Tg^>a]T5Gg@FC\cB81=;+X[QBe268]QcC/&\MGUPT9.HO>T8-I1JPbY7(9)g(>f
=aBDCe?/32LeVBU7B)RVRO(OS._T_KA2J<0G]U&3,T\bcG;.,+&/YQU]afHEF#S9
U=\_G)..?33VE=M_)=aNC8BVVWCQQ>N0C-:XQKYB4F=<_8#^8<93SKJCU04[B^5M
Y<5AV^cHIe\C]BcIOV86RXN_RA9JL6L>&OZ?V@+NZ6BKJBRTA>R1c_L9GZ\NT-A9
UNH5,c+3aV<<J4BJKWK))+E8FNPBcObOAF248X72>I\7ZS^aK[1-/E:WJc&V:SX[
@;,^78[.Y2;L6.[_??(7c]H5PG7QGUU@ORI@c2YAZE>aIW\cfVH5]+NR4X(cTZKC
8=H59c=9_>)eSQ4AH?_;Y[;BR8X3LaYQIb\5;^NJb];RIDN9<SWB9HHaDg<Ag1:g
=&Sd;G8O@I;)UPa<TAD>S4=\T(?8PJZgG1Ig_,WM]1f8Mg1C7BFRQ#@gVdcV]P+R
L5F60B?Pe4R7Q_G+:J29LR:@O^eX-PT#7(O[N];ET:+.U6>d+,WE/YMZ3&1./2Ze
?[4WEUc^8.gW#^c.S:e>CG=:U=GI_A9(f^IGG-N>U1>-Te(A(Q:OL#aN>XTZNe12
6GfS-FD]:.Zg9:J[^LOg,8B)I5Y:1;AE#dP8^b#K;c#74W)9F+0;WBb=.XI,X)V9
@YV:Lfd]U4.bN;d?QA&Z3:&.(EbDe+T_=Nf(YZMEP=UgD?SL2XW;eJ0V6W9#aNHC
PTfE6)b,F09H)[<TBNcC:.g^:KY<=0eW>)Y<2TXX)BS#7<27FLSgQY/4^.UK[C;R
0ZdE:2@e4BO6U0(P8\8.gG2G54<4PK9]:c1b/^aCHB4=ZB?Z^\5]g&G9RDHc/+gN
<F<gf4;<3eA>I@&A.-S#L2JGS>+K.M,/.<Q66eJ.\2Beb7gJXFZ\YVO9YIG,[QTc
+GO<eI1@+V+948/6AU]]Kb5-U)WW\JX9Z:U;&-eJ^\2]Ua#R&F)1\C()V/O03/I8
JG1fSXV[B]IR9^4db;aS1ePO<J=f<[2W;M1ZZ)MUDf9:6UP8\2GW<T3RW9MPQ1\^
)9^@P>KaZgLQJU0;00&?5#W_KA@;AZc@e?JW59M_LEZO>TH,g.H(C7^=#T&fH.G+
:YL1fT:e2A(^V<(S]RUCF<?P&RL)6aX[>+1@6\Z=6Ja.,JO<ND15X^B70X_ZLUGJ
O<P.>9HTWada5R@.-WXAaE:E(392J,aU5AYW2HW>DEVKd[dA_,[Z#UcfF0Z83JUS
9+fG60M\?caKVW=F(^#?QRMHNR(a8D\A+Q=6R4E_P_OPAM2.XM:64d6HD9)C;#>^
>6J953c>3DdI[&R8S)@dYZW-+6RUG&b0&\]SQ/5A?LF0)/#K][]JOdgQA;Y]A8>4
E6)2IMUICTZ([4\+/<EQ2a6K?fO]3DL]b5;W5@LFeD(2c+>Cf9@4WQcD3[C0b1fD
>B9=XA6A3B;3CU/:[-<M72M]Y1]M9e2ZR.#5KeRG+R=Ge:4[^WI8+_8UNeIUCUQ<
\U?f]D,18IQT(f=eBAME0AOI9[6?^ORV5eVUGO\&5@._G-,:B^+&0;(@bTBR=PXd
_&>F1ga9BJHf5M]#]@AeAH()<V+f^E>6#+39>1<1USTd31,>SfPVcKZC#0L,cIZa
Jf&HT_Z>?bLd8b:4FKGJ5X3WMY82?HD?dEgV]:ZeGY]=De^05VSHJ6Y@ddA[=(0P
F\M\Udc.L\KLZf__(#VcP.MAR#;.dZ@=U,ZUW,Na7^)0I_-77cEc8B=()?<?^9d]
R39/cYOb6)WcUAR^g]L:K/CK+HGM0+UT-g<;d9:Wc@@g-#P<#+MN5X::\>U0+,&2
b_L-W-6UfgAc/$
`endprotected

`protected
N;D\#ZUV:4(ee,e3,9EHDdH)U4Y3>@)G8c:<&G5-PC5JMe\HL#V?))Z/\<+L@[g-
B_<XV;N<4I&P)AE(Ib&6/9[UH)#<M&.\?$
`endprotected

//vcs_lic_vip_protect
  `protected
LO/:?(7]g;T/cVc;\[?bS,b6R^.d[g7V>.JXeP=X\TC;bBSH0dG3.(5],Z(4]R+-
UE?Y=AHW+_-;GDXH[ZOXJ[-P9&XQ&S(dTOR:L14PVRNUgY]-QA4dcW>S;68+PF8@
?cK_/L>/_b7gL5<V;/G).]G[Hgd,;QeOafK4#fb3e/2JIO?T?W9Y=b(R=K>;FTA&
T4=DU+@)ZBg4^V9TK][>W+-,+VHDYB)-DOOLZY=NL]c<@D=R5NgbEH(_d^8VD8Da
/92IY=DR]U.Gf]7),O@_@f=_I,d[X\;)SD]cN3KZ;71Q2(@FgJHA06+FOHb>0_6L
QDLAG4FR7#XXOX)#8F6+)OQbA=J,b?=X32K[B1PcWX;0O#1#F>S/5+]T1HKe@)-A
.SA#YEDNAQ(JGWZ8Ie1RD-THc9FT:_D<--fMbT1<06MKgPa#7<c9Hd7MRJ(]g4KD
VNSI&_GY4X1.PBPD&UO?5I;@A>8JSda[BQbQec]EO\W&:+\)Bb)bZ,3f;Y0/]LPB
c32741O5=bW1CB\d,C\7TeM&bJ1>M0052[O>>CS:,2K^__a9MP(aQ8OZ:Ma)O#b^
e.\77&cf^A.2[#dUeH17RbL[FLL,A1-[WLQE?2b;<3.7e@SK<(FA1BW_/FQ+WH7E
8SNa>5)8\e8M@6EHKe))>Xeg8<G=#J?QgdBX-^L999&/[=>c;-[9>4_e5C&K-UgE
H&2#.<@984Z=H.Fb&G.[5.&DX=<>3X#LgV<:#/WS:=.6/&L/#Pc(9Y2[&D?c/(BC
)2414O,ZW[+)/1)THI+C/SaA=[eQ1P5g^EO-(X9N:7^9XJ@AEbU.7YMQ>_8KTeV]
R8L#:QgIQ5>ZQa^E>_bUSfMd081]9R]a::f:,5ReKW]X?PO,N519_/2S(E:U)2JB
^=HQHMa?,WS^8W2F4P&N?TU;M#8VD5,4H>C0eO,bPDR,U[dU.(=]\G(PUUGb7Y/T
f8:DGZWR&F53a/XZ+8F5,ZCf&,-44RTeEA+H9a4L8.aES,=2K@Z1G2L:8I[9X/A1
Ef<E;R7.(JbQ3):7#4GMgA09bMREE-gT9)4CbDE<3N6^L[6gGI,F0/8bHRNf.Xg1
<fM)Sd<5<P5(\DM.N=#M^+0UWO>J]M9fPM3bg___+_E^&Zd-A,UO34R.MM1O(P@g
QZU5_5A]D\RSU@VZfS;?^0M\>(=<_@RR0bZ.O?KJH\JaVUU:.C=T(6@M6+WLa;XW
7U8)CA8HK=QBNS5S)=N)/W575QYU^ELgMK97L^ELBc(_a9=TI?1B3DaNbQS1CeNE
.\EB4)\7cLb+9beF+3CS@QVT/Y>?g7QA6#+4AF&dXA=Kc>H_WGQXBA))F:SA.([7
0O_<P5JRDa4II6ZG5:OJAO4d/1LeeYIZ4KdUR7>-HX7]?TBX/)YPHbT0a?EWFf7a
@O6fG0TSSG\[d@c<DPC=,g:Y\J4/C2]ZH7NMA+f=09:eR]YFX9V(IA?Hg_Z458OK
dba72dPY>UI.P5@6eYWG]JDN-F@\<N;ce5UeT,K>3^@T9#2eEPB2fZVfZYE7Y.G:
g6H<GZN(&Y?49#Z2=?</[S7GMJ>54XK/B?V&U1g^);RGP5QGCB;CJ1Da?GATe>@B
KaZ>V0a07S@MWc-VU&]MaM_:7Z\DINOQ(/cYQdVe#EF50&D#5@f7=-_H,e:AaDO;
Y>0?UQG_>9N[JDgVI#A?8_,IHLWHH:F]T-8a;OH97=M6<#MdO>Z;>/7,d[?W=:[9
VR-VQ&&U#A-@_S9W8HE^X-&G83g:GX?JIS.E&>WCBA,1,2b]_6>4CBE7TL_ED#TB
C3<X_bK1<4EK^I^@CDRVA-AId:S_d\^I3H+?8X4<U/NZ=O(+J@>5YPM;YaYYP?cV
2+6OV2bHfON3g<\Y_58gJ_GYOE+8GPK^/BeNBR<L68>>#cPIeb1b@e9.9RRPf>7/
)^)A;-46^C.DcLIWfPJ4U7.1eYe(<<@B>eI5E87IAHFGB]dVU@,=0[UWb-6ID(Sc
/N9aJ/Q;QcKAWSb?)=,ec]?0<cR1HD#RfI9;d8:1QR#G]RMC#Jd82\_)Y.DC+0)@
a9;/<<YeF/_[/;E9Z+YDJ>Z;-gaQLY]bcP9RMC.b=_R#2ZZT+RU-)\&P,R)8G5B-
BA@TGPCS?B&@P^LH3,aM68C+8B&:Af])LL,]XP(d/@\Hb(._8H:]M3]>:0(<<)AO
L_MDPDK#Z]2M6D]G;)NF>0LOf80GE.fYPO7LbZNAPZd8>dN]+ZZN>=@Y?ULV(U/1
cHM)&,&6_7DgF(A+)BQ+Z7RGW_DQ7@,]=5fNPG:FY]HRaV>:<;YA&YIf;0R#JFW^
f>gcE74?RbE1.L\8P&=J@e[X0^E_/O2KD@1&WI<ZfM9D4&8LN5D72g;R2bXIRN9T
c-C2EY1/^(>Y6LOOe;>S&\_CD^;G]OHf^4/9D7,,/)_7\Q:-/;;PM;OR-S;,^bZf
\BLS_KJPaKQP=;H;55YFeV(V4=8-&E6GEXD[O^;NN0J2RYCPZ<4>Vd?#C+V4X-g.
Tfg]=HKM5:-JA2E+<\\gK2R(X)<R<e;B8K20;=/E(Z=[P2RA=E1?H)793.?LTF\Z
6QBgFO#]\P:MO+P=P=9Yf7RX@QO1S3\SWV7bHa[#B=>O;&dDagC_(30CHR-T=WB7
cY-8;-(,eU^?1[[UO8cUH(PT&@DGXL>TIO_)Q#g-.U.,KN0[E/^H>N?_PRZ9SGSJ
8F8;YFO3KPD.MN,NRPTIa.Q((JRb_e(\O</L(CfAcRB23#eD?@<9?ZL@0EfeOC<0
XaGU8.GEY&a.7/g:JRALa1gPaV>NF\/Lf]XRHQHeUd7S#c;0[Uf:+#Y+YKI)R5J>
+R/19U^3d5bICNf9SU2RNU[.dD@[SCGU2[Vf&BCO_:R:4\@aMf@G1;4d=#\1P1<[
HPKR3a^b]Y.7AG45?R^PcZ,7-a5VW,9C,W>+d-BT_7W97:cafSM-KgIB9d^Wf?CA
^?WEV@86D];08EXDb<ZL@QCSYR6_ZG3\GK:+e@)P=Q]I?1(IcUCAdDe[FJ:><e_U
X+[CeI0b@/DMVB)K7SXXB;?8\Y^]3J?FV>fe0)=Uc=d?ce<\1eQDE(dTZ9M#FfV>
6/#AdQW6<NM[7.#H2K@?XM)5gf+Ecd\50PSaA1M]/=5:W\W2;(D-(]A>6:,f;C2?
D4_,d7+@ef>a_fZXT]W::^6T9:K7aY9/cSZ>V^9&9]R<IB43d,dgHU-1HH@9R?=F
OJ-S4c32AI7)fXU?;Ng4I?=(YIHF=DXWFcS37&,F0?4WS(G?-EI?(H+9Y/@[D2-&
F,3If;;,S;LEJfcOeY)Q].bHY>GREY@W>9HFe8ED\:f+4U4W3FVW2Y.eKX8KZ#3V
0<\A(9:]U(FLGLG;Ld+1If<6:JY_?,?XU[fGAY9[NGPN=[R=b=1UA1ES32e(B^Pf
<OX,,2)&MW[C.5#cLUI=P0.5LMGHB;P/7X_A[:IVEM@QLf,Z8e8D81,0a):B1N@,
aP1cGe2^S7DZ;5bR)7U0?R]U,FZ)?(7;SSSd\O)YS0)Ec\c3g#.NG@J]KY,D[f_<
#&+)cYKe/?ZAAeF^K)bE[/T^M1&4Pb6dZXG1aN(9d5)PH&,TU.^D\S;:(/3>:@bO
[@0d]+-d<O;2^Ba^=S\Y+)O#Wa=M<PPH3_5LH\FAHK>Mg<J_eRQ??)/GV[ZA#1+4
LaK.G(QOAY-&KQTR2E_?;KTAL;gG6IQGW,Ua=<;K>]]@MS8:+U#J@Z0:D2<#g,WF
F0Eb2I&@N_O>V(d__1@_HR9]RJW7J-K1d_Z4E\^JGD+M/M(Y#:+P1LL]b:2;TK[^
WH8W_S(=R:LVK(0[)@f-N#T4M=DePEYZ#4cfJE[9@g5D2[V;<=g2]Y?B1/K;QHa(
[&Gd;J+<dFc#1&d\,<^-0>@bA:MMU/_[50:1-KV(5F\+Yd:b/5be@=YdfN+,V?aT
=YbI)B(b4a]S(d7F7FG<CUP.DY6##&f+0?-cg:_2(O7UGKd[>_SZ5KZP@W:G\a2a
::>,b&?3B<O-3)4+8_KKL^WVOLGFTRNK09I;J\f-LO?H2A[dI^Lb;>[@Q#81SJ\A
35,c\([2CMb::)K#@W/8T\1GIL3:)XE>W87C0>\L<L.IM1GMBRR(&9E)T04Z^/RL
C,:E)Z;?#]+51)LRZVG<DR>V;,36;QVecZXPaS+3J+]?Z4#)Ue-P#;e8Lg80.Y2M
-eW7ag3K@A;R<W=[7,2J3@XMA_D^UcE([R5cg\L@0D4gK.7<+>#IfL^<bUA9^EE@
08;C<U^IAcXDBCM>\2<e(BT@AV&];ZgIKBV)Q_O4_12[NTB,#e+\9H4=PO^N2W\b
\O4SPT/gca7:U.e&@VE5JJ[LW@dX_fSA;/@<b0()@M.F7dB0+C(L.RMIFPb;3;=Z
3(0:L40\#WNA.[U6DL@:dBK=5S&D.Z(#A[E1d>O#R?J:4H,V6gE--55-2f+5G<PV
J,WcR=Y)RA1(&_6)6PQBLfD3;g/\dKd>DZM)f^S[),):bbAAVEXc_/\XIY;fWa+?
Ce3NX&T6?Xe^V.#Y[&.e^O6dDP=0]GKV=.U2UV.6)f6<:J7=Qc_7EaE=3bg+KG^F
AAUOZV4AaL,D.;PD#-7V[9F@7P-\U1f]I2dO(>c86_FX0cf:.J=TR0=NOO<ES=ef
8Zc(7cE(J?<T2+Z@4f\N:UWP127Z3[2V\ULZ:C^8L?SN6::JQP^O@.a0d<<HfYD3
(9V3-<GQKW?6(DfB-EQ>BWc#(V6=ca.(XWN??IF2-4T[KUY&:]aCFCX83?\W]2TT
eb4;=QK36X3=bN#6]+[aeNA@-TQ99]LXRa,18K1MG.SMf;B()X\;ULW)WOf0^LLW
8L);Q,f/E;C:c8?Yc12M<@E0OT&R=NeZX7@8/O3)<eM?.-7)5a=^\]@,A.cE1:UX
3Sd5N(De(GFA]@M:40EU9?F,6F)gV-]d]W]fgM)-f8&A,IHLaB?#bQ1,#IG3:_8Z
9W7M)V9>W&#WSDTVOXc).MD]J;R_Bde>)?)@_BIBM_H#&a)NHQ^BOX9DJHX)g-#0
(HXfCI.dCFN099;4V.AeN:_fBHJU-OEW.GS/D^U>7A+c(dP]K1Xd-/UOZ<,2_(0b
K:UV5WYX]\L&WJ6?[>P^FQ9L_+G=9E0^IJ)+\S_/NW>MDYV>QVDQc-1SgWV_H>XU
0XUE0_<V(3.1eM#>&[P;ge\])B;FR1N7a)=^IDHS#I\\W.gDcC^8g^ZLFB44[PU9
W+^[cM96c@[Te-6Tc10?4.&]A=+AT4QP7X\d/a25KJ77#-A-/C7HDE>QV@KcCcDE
DF&C1Y5b;;d/1/V&d&OV^bF9+M:(/N)9AVb,#.f.X5^Vf0a-#E(R#\/;fG?6DNC5
\76a3X=4bcF.,/fYG<&LB>P<9Y=C)ZJ-&V216ME2ccP(3U68+A#C/RTBOd02M7\6
9B&aQT(DGfWOA^)J1=;24K/&U/(VfVJAGYS#2L)BFA^Y6<_Nf3d,M]_GF#11:\e3
4ePE1d8@<P-85SS;?IIOIeGfN><0?2W_1:_(AK1>B-,C<e_8\:L[H[S>MFXMQ?13
M5J:YY(>,NU?.QYU#e<46Y-/HWP<^QVAH\T@(b+Y2D;f@PDM_Oe]/Wf\/D(aP/N:
bA.BO^@_<XMCKL7S;bD3P-1BT&OX&:KA;B8J+/&-@+\^7P\f8R+1==IUaM+JJQU(
KO:(C,R96c9:=GOV.8+]e_DR)GbM3LUN\RPU(/YCe8Igd.+d1ZU:TS/-/5(Q1W^&
QegYP7A/VAWBBF>SXB2=]LX_#4_0/c;F0bAO\3KJY-?,eSINHG\&9S83a>b2[H/Y
>4>]d+ATDEZOTE@=N3Y55OU][MRc&]Sa[J^CXL7.7UV8;CVAWb[dU6>(ZcJJ^#B]
X=]5)DRX>OO:f),AS6g>D@b[,;^D@NU<50dbFaR3U->1e&35:e35L4ZA&6XO45C.
S=7SO,27^CgcX@,YV+#[E]I)O.C9G<R_+,9BF.K_gW3>&EZ^IA24e>1MTOHNBBFE
3<F.4V2<6B[PW8[7\[MWY50LZ6SX+1Y7<TD00-OW=]9W=3PY6]2L:f-5816Z)CIb
QP#Z--TU,>_=XdQ92<)MXAd,+SBDE1C8D+Q@KbN\AP8A?>,bFH7(\WEJ=XXeAH?C
/b^,O>ENgMcA72:(:gf586JLN+<IH@AA\Jb(8TEA2f+=FL&;4afZ.<SC+f2?)gRe
]ALKM_7@6ZN[8K0:ZQ@,=?T5Cc/1eN/PDe,LDDX@P6>>1WB-,IcM;S70+HG(f)QC
eI^]IJ?&OB3/2;>\4:[@J\_B#:H^QK@Q</8^GQE>5JTAA@FGVORW5[7J/=O48XQ:
7<@W+d0>K#:IJQBdEJ?19^6\.[@I,ORC29_68gM2DA@L.65/7F8S>N8N.(/R=KVV
A3X9YUB6c7Y6Of]ONLTWUb[;eGC-[UD7@YAT3TfJX5LH4Lb(]8,2RaDA_fbPQ,.X
0XQ1SOe84NY9Dd=YD8S5gEY:\\J\@4C[T@YL)HKGKEf8=<SU4T>bTG0\AN@^AUB,
GQD66>Wb<T52_<YDYeBVXW2<<2>D825Z/Q<N)#\JMR820e#[UQ^RV)CR&);5BF1<
PdDP263&(F,QfIC7^SabaAO&_(V\#^\,a)M>/;a<0?<JfK<[UAcP37TU4ETHeKBa
(5MUHXgIc.5#C3@[@@=0;WVQT<V&YR.,E#4O^#9@-867H9.8_FE:I9GOD=GW&.TK
#gDN4)Q.JE9::Y3Sd0T&9gcf,7@.S+?SLS:.DE9I/H1OeL_O5;GV.1OH0]-9GJQ?
cg,AV_=AaB+9@KJe9AQ#&FbE37VYI^:_c-gKBL;HXO\2/[:a4R5NJP&fN];(2+[Y
OM2.E.,NX5A(Y_=fY[&e(5[Ne[4V+D<;+4GGe#d?_)+Mb]JZW&4;Qb/>EAOW_0-@
_.2?2@,L2/XbZEKe@+FS=+I-M=IfM@VY/4:=@:IM7IC8L,@00M4X0RMSY+0beb25
X>.^Uc]eS)GPTP+FD\M#fUZ@bcd#\Rg.\);7-gKa\aXYbHF(+TSLM(a?d=Q_e<bI
e9:./@KZOKR6gCZ\C?TAOX8R/5TMJ2_6cMR:[1SOUG&(O_a_>.F68dg#R]]KF<@G
THL1JOGXF(.FBAJ_FJ^D5FaD<?BQ=NNdA#)_&T1&CN)5Zf5B8](,VC.G4M1JA/A-
f,X.Wc^c@ZP[6FEbYZ:T\KGc:G>OD8X7VP/7H>-[/_U&J3XXg]>#;S=ZFP5(7gCM
^+5=HE20K>>I:JFQ/BD_\\MN@8&E+YL>TGR[=T_=EYHgMQ@^Dc\B)bU(@P:.#Nc/
;QN91?cCH1bXEDORKLa>TJT_6FCT#R5M6cgB6d2RO^8IKG)(X<dTK4c&aP/_PKT:
.NaUQ^MLRcYfW@.W#4.B(Z2B]U:(IGW6:6W_^a<K&5SXV<0De;\c58PcND.J)6LG
NIJR.Efb5#IJ.8F^QU9B3R.FdCU/O7NN_,C.48QCP1beX?F]F=2TO9):/R40DeBU
UC+D.A(W2Of46XL5<dM@_0F5Ha2=YA=-:c2C&<^(>P@aM/0;@MWK7g^_5J<6Z<G-
,[:^<EB\Kg&Kb((O=W7LA_03[Le5eOacgU^&5JEd0eZ<\ARL0WHSP,[1H9>;O,P/
YFJI&MUNCMe,1[2Q/.3I.XF?T)?]5X?0IWLL.dEJ?7[?47FGZT2<N#PT&N\V0SCH
bWA2#Y2g5^[V;b(S;CZ19d)QM=JQ8C:eE(Xf,eL[AYB..^-PaS<HGOZ61[_6#UB@
gL63d]9J_K^0Y/U)3V,-=Y8SX1<8RO[:6.ROd].F<RD=7&5:J]E+adNbA#4B]O0@
,+K[CSDUaVG4ONDZCe1P:F1FKf+HPf.W(LJP\IB5@Bec;[IQ/4(MM=K;=W1e9g2/
=WMAS@EW03]J)F(-DZ^^I-f.3K=DT\?f=3AV^N_I-\Kf/[\SGUH&#&/5^cYIT^]@
&b<2<LYGO964J__CFG=K+BE?Q?a&7A,G-DLE[b>c\2L9J2/JcTR:[^/L=8].b#0G
:)#7YL4/S.>.Y^2QcER6JgR(GV\N^VL#=)K94S1RM>4SKEY6)KWC(AT;L<WXcK;@
TVdde>#9fe4+0&48;Md#?JO>1:;,M_9c.#7WK+FM<CAJ/OZ?JXCHbYbecHEbNK3D
L9M^P.A=ZYbFWZC(3;4K(#Lc<O&?-^U\Sd,(#]6SQ41([6YT8AGX[.9D)E_9U#9b
WP+R8be;?@.[MaL?Oa(&J_\6XC)LK?ZYX/?EX6RO,-X(UW?aV:a;.W/)KeO,Kb=T
dO6Q8+K[][,2#+?+-Fe-&[2(^(DA+6)#I,.@#</XJ,FMJYE4+\637_G7bD)/:D<+
aMMV<QF<ZHg6+W3LFZABb1KKcgMWJ:^F=GEJ:cW3VY92Q;9eO14P<Aeb@gPD34Q#
6W#2^Z=.TF&+#I3R\+>,OKMRe..P<=4?^<b;CHIVdb#X??YgWLcC2_g3WM;#&#Y:
QWE^Xb4b@?2UQSPE_6c<]GVcUJ(TSRYGC//.f+R_D-^9KF;+gC1Q)=5F[JFDVB13
>bI5OV@_MW[J<8b]QB5cM0L]ZHFA^Y>gT8JYEYJ-XgQQ+>BR2#b>6,3SK]BZd3VG
<Ig@QSdP&[d+(EXUdMB8H/K,@[;BHaSc2U@F/)L\a0.^=V2JQ]EcC_0AcX(35J1C
d>4I(I0;<b55d-IX4](d1[fgIdYMJ&OS\fTWS[b#AC1Z5gNgRe9N+PX>9FF<=N:(
P3)Ca]9<D:K36QR.WJ5Ma7.1D,LHPG:AOC+8WI:d_L9C\1PaS,QKbJ:Saa9UgOD+
X2T24c7XNe.742LJ#B3)NGdL1[?RGO>#&21eU&WCNL8I7RdbI=^ZX-_WK;gZ[0ID
&W9)6DQ9\E(]17M&J64E;/YJ<C;G4<G:Z^;33@D7TWGa:BMZ[8/8S@dA:d7[E_AS
g=S0C]D&()a,c6]30\N:Oe^<KN\eYN9S.>+;N]TH^#:C)Z\A.,=>4.;&CU)(6\12
SPYENgV304HFM#OdF>ZT(#;ZA\-R4Fb/KH29?7J&@cTDQG0SQ;GfV+f=#\I[]=XT
aC+b1/3Rb84-\.ZT7Y<I;Z]@O=e[?g-b1[F+:P5B[/51aRD:cBEe@2=dgLN4KTa_
A/a&[YbSbePgEP35Y]]WaTg]R=dX>T4F<(LM3#LNR8adSD=WM94NB4R@N-1->15,
PUH:R1-+fXXI^U0,,Z@J74F-<D9T\O3,:[3F:f2_Q?.JdZDBBX&A0#NSY+M4d:^^
GVGJIRRQFS,LUDeX6)O6d)bb2?5IYUU(JATE#3c5^;0XHI.L15AY@>L<FHa)+Ba@
<SBOF:2f_KWZF/+CP)^JbJ@5QR[DCccC=L]-T^:bg5?^6b,0.f78CNTI:Hf7eI2A
#RS.0]GE0+Pa>d?a8:68,AHL[TdTW.=Y.d1)cUdWPSEQS#2M?M\HB\<MGOPNVLVG
D;#4Cg_29,W_2]WUD=+REI:_0T9:[]HAJII1._16OB<bHee).-C:F._=:Pf?S/YJ
,WTg]Ve6F]c\L8#TM))\M\bS-?XN6Q5GN2@C54\_K<V=CD?^c[@[:GPO<M]8[M4f
Y0bU_WePSgc08MIaLLA=VY&^E\<:A_R>/]d3:KCIQL2)1Q+LTDBJ#:QX7S(N8@B[
TWQ\H05BaCFJ\TZ,CWWYAC]:,SaG@]1(5HM\c(W)cF3+(fI,7f#S,P2d&]-^\Ec;
[cEG?@76Mf:,O_cC0@E/\D^>fU#7RP2]-5/?0E[:1+&Y\TIRb4g<a/[;D]ObgL6>
BZ4A#CSS@[]SbT@>aTg(X4V7Y@FAL@5)>dDfI<^],<7#GcE9?911<a8ZA0LQ&<38
CUUW:=NL4.3Vf6TZWLe&U^6TfVcR)FJ2QZ57K^0IfZ<Ub5ZX/AYNDYH1:e8W&S:N
4N^N^;+(DK?I4IJeZ/+&,6cUgE\><CY07;:911d+BIg:()EM&Z3G=0BZAW.DU3XZ
^\&gc>7cHOZg+f/RLA1(Nb,@ggWJa),3P<V9A>(GISg#OKRUA4TYO-3K@W3IM3Q5
^E-+NDCBQFJ(57AL3J-[E8G+.MfB3DX@dXM]>HCg+SH(eT3&Bg)=_9JM2E;B-+Bb
fS[F>U>?T^.^\MOGT)USe1UI:_dXU6f:1O7FUT0bf=0WN8,Oc._:2>M8:(5JVV3a
OTSW)[9^7a4Z09LIAJ6gACcF0/c.Kc^#NA3AfKMX1?_fYT<84&/UJ_GI/&4P<_S>
d(3P<+Kf)JZLF>M;,&M[_;<.-?8cXD+/-\Qaf7=X<,1#@704K#\J\Q;MQd9<&4#g
ETJ;0YX;6MR&52#\=Uc#]-(cA1-W2+P39#41UP;3J:bYF(dddZdaM#6F):_(4RP&
>V_1>I)>,OdH[E9^)<4#ZK-E62INXg[S?E?/R[Tg7#]>:9-6c4eWNR.EKLR/,SMJ
&EFP_,+,9f@[a+AN)04>CNR+;T[dL-\^N7BB?<U]cQ8&0NZ^Y2BAK_H5U0.&QT65
1Sba7]fdTbH^7cXKB.&/?B0EU590]ZNCd38N(A[E@CYVLX.6SJ[Ge19^-MH1;6M6
Y<FUV9Ig=\CY@N/YW&U(@KUeT=#>Ma,DFFGW\A1MG^27_QaaRKGEB_L+S.HL6M0\
>CBf_DK=LMg.]V##)]@<-@c][5AZS37RMW71?=9UU,B7==-G)1+cHX?6@SW6ETET
FNIcD4UK2><,-,d7J4^(:>VYCZ#+dN021S[.fT:6gAS8W5[?[Fc/P.@ea(F>U]7L
M;^@FS1B)dZ1(f>RMa1P^VD^?a&@):g=N<F[URXbQ^SPOeDV(0X(g<a:)-EcI]e5
##]<M2R1^:S@O##]<_MB^I8DFA-.daA6gY]K(:<&B:;E)9BS7^K++W[BO-a8+L;D
E>b\3X9FOfYbf1eN0g72W\/)Q8Y0-#?F]4-AR3]fH8f_EHO;5\MK18L::dHZM<BP
XN-+bK;E212^>2@D=1CC8OVZddRC_WRJ1GSOJNF1_KX22GIN/L;:cTHGO?f<3c4(
:3e\Qa:/N]O:0#([06H-Z/&Q3X23,a>>:?fUL1_L6@Y[bV,bU[g6e<HEIIfKU3T8
WLD0g1<5KP^YB-KA.#>A6Y0S+b@R1c3XdLgKBJ/JAU13M\VMF\>H^)Vc,H/OCVB1
0M4P3aA>,a[HDO_:,T:>P<LNII&1HK&TU,7a)ObKfRQ]fFSVVNA\F:eaJg6S807:
MMD<9e;FBdcJcL2MbKPL9E&)AWML&.-/I2EWFA4GgQQF:B60;I^E^@OHVG-P-,5-
@\?Q;DTWMB4(RP0GW]:>;J+b];81eCb>QTOO3Ic+_A+C6d:]a?\fE&^:5]#F/497
bX0VD):1JHGd3gE7e,.DKN<PR?;J1Fg6QJeI;:-VX+1KYd)F].XBJTg&Z;/^B/S\
,D]430QZVH1MNKX&;9D9\-J2f(-\dO1f>BO)e]]0FFA9;.T&BZ@T8;271BBU+,.1
#OfEQDZaG4I.VeB-G@Tg7<&VUU:^UJTfb_6])3ZOKWH]BC^[)T/F?#;VUBG?SddQ
/Ff(]07+\:IWbF:=^8PO/MFLgc0>IJ;Zb+;RZ.dBI@FeY.(=RZA7a;MfB]NB_HQ>
.ZaC.Vf5<#UDCHe;O)15\VDR#f(Jf_(M7OeG&@-T19Z)^<;9@<&agSWb[_3WO,YH
T#\/,_8/fUBANN^EA7[/1=N3<eK/G9DYR2)f-ZGWJ#J<W^7,:=_1Nf1+e7GWA<9/
:a,SS)6]EQT3QE#8e(@<QAYGYP9H\B61_+W.+-+(9?0]6PgUA1Y5\TfbZ<\T>F\Z
E&1;E+=H5LR;8K213g-g++LKSC62:X8T6E8WW?),;JScA55Q.EgD8b6D3ME_8#b_
Ma\Y6-+O]0a:gVDR#E>0)d<,;:,e7ZM&?=cHQF[O+D7Af:QAc65LWD#19RFe(YPM
J.KDVC5,>@AMR1>VcT810X1\aJ;dI^1Sbf#ZYGIJ;<CN:5K+@9E)B-S->B=FcIc#
YfO)N@9Wa[646666aCA#I2J.fVXY6&YDZ+<X^QQ)VXA&>;1E3Maa^A-S+RW<>CQ-
UYCE+]J)=(9CE6:fP(2#V[RdK.:]4_/:UBAV>&Rc,4E_TM0#:ZB<Q]>FZe\Q-XIX
S?K:F2NP^@D5b57</f9?66E(MfD\Mb8)RZ?OR62:+19H.X0b.,<3S)S@[c5eK2dM
@Qa=.BM;Gc9Xc?=aW?b2+YOD42@WRCCf@SbJSIYM_c5V98Q6f=b_KROG+&09C<3/
NHPT&@7EML,G=Q-#L=MIKWZQ\Pb@9S+E.IACeagC^c?/IV_3>^@KJ>-0C_If).0E
/:K\F?BL_X/DEcG]^I6+gg7]G?0K698E4^LPFN_.9],[T-D/S-3[Z;4E_>D_ZGMQ
XdF\5#W2Y\)MP:Z98APdcP7d^C]OIeKA45YQK[F,W\eD+5If_:HXXP;Jg3WC&;&^
Y=aPE;cI:>BVB:>/+;\bSORJ-PVKXJY=dQca-&#A8LHZaR1YVH2:e+&]]>>MZ/aH
YM7PLJJTN_Z0(P+&A>&gBg@1VSS(H7?HY3+d]EWP72WPNP_XJ>_D3H&WH_S6d3B@
Ib?_1Y@:fGQU[1\0^5E=<FB?_gEIA)GW]G&6WN[ZR/Dg/Q[[X5-M@,/0-cW\9[Kg
L9LD,PH>+,7KXZ8e)JE+10d_VcVOA_MIK.SG41H-c]E&S@D7LL=AS[cV1P79R30#
CRZK,X7XV;<-@WC5cUMGC7fH]@NJS0<CAY/JCDW)&SST-G2V;3(Q7[^)XZU>/E\]
M+8:P<]2Z#99JfMM@B-0QG-ZF2.eVCHXf)dE@MH7bb;2OA-;:g^):d26c<U4GF=:
?QNc34/I)S<SMMe6NV.=A:@:HC]50:a4LbY,I-4YN\GE]2X=Bd1aCg,\H=aQL<;6
\+Y+>MIAA^4R_4+_]DVR,g8f]EdDaA19Ecd?dQWU\d&KV-@ff:IeMaI=]2G5@H1V
J=^(KC3ZQJ)b#b<_b>;Mdc#S/1(a)ERd=NS)0H^W=VY3Z7,32VZX:3/=0Z)5g3/8
-4S--E,LJ@TD;KdEC:KED(f@XAMM7S.U/CYIdUcfB1L+c0R.Gec0HD/OA1<K:>A5
QG7Jd\V3SCUK(1&Ac<LHO3Z6>;])fUCXfZ,6+1g1H8d4X:#LQ3LGOCEQ@HTG2c4V
NOV9@,dP_#]f:\?AI@>;QaX28R:6Q=VC7+U3/M0E^\Vg6>;/K/C<B#d[#XL+Fa00
@B2UE(U/]WG9[>:2e21[O[8]P2WbdW2J(QO-6bW^P3L-eFT94>\6K?TZcbMECJ:K
4([ae6Q(;IEY8I:)]12IYKEJZ&APc[&WFPLe6G2:)11;BE0&+^0<?ag5YGUP2;C+
JL8H7?NA#XE&^Q8[3.HD+_faH\C]-;L_44Z-H6S:#/SBA6-+P2L2IX,PD.?=G9<0
Z3Q6J.(@PV/0@/@Xc^7C\BKbQ7GCO@a[\@;:X)d\N+#gCA=.=a6a=Fc4;^_[f(.2
+OF[J3^&ZbE3.@&+FFc[LdY)>);@B-LDa7/59VD:P3<a,VWfX+N_eFI];^]99O5,
,b4-a_X4?V1b0LXM=AK.@^LG9)UV^?7AV=7I[?>GWdPZV1C&_7<:e)U6@SaT;&F8
8?g><>?LO7<;S@-aU3;C:;UT2?IR6@:dN9U9J#C[?#UffW2;g/B@=D&FHPQ/cS+X
/K\\7@SXc83.@OGceND6PA__QMcHd-<]734)43PYD3cSe@U=0]Y\&@ZgLX_cGAS6
E7ec-V0-&^H^S\1/7I.[a+K[QX-3+##2=7CE,gU^cN>,,^a_c](XfK39)EW0,UX&
:(R8HcgIU^IU_&FaVH\DR7Q5c]:L<BdG([4B@RT@U],IAa,e\N\LF7.gP[0GOLQ_
4-VOZ[<5KI-@,GMV.(FYS@@FR[-Fd)4?4dT0>5_57;VI50ADU;UI<f@&MY9#;4BY
+>J>3BJ;B3?\Jd_Q_ZcTMACU>N\Nf-/Bb3e>&#ga]=D7>51_bD64#7SJSM-0U0=Z
0T?7b[C1NV0NaJ(QHPJ(90^,CfMBD_/ec;,KPE7g>/1OQIL32DbcF7XO5&d^\A&J
5[\/,+>T60XCDRTRLa+2B3N4e?^)>\Ec\H43ZGJ>.0HL2.LRIKODGVFAV+:NR/_4
fPAbOPN(J>O@V7>[#aHV46@E3Q:@=>>G7b43=fD=I:_bI8TW@/H)\fP,8IVVQXL7
,:OW,P3=B\dM]TK(MJ;Y9LU:acFc7@eM=Jb3f(#PA5<4(OAL]T:fKI@DX-P:UF#9
PBHbWXd1KPIC&KQ2JU/M.\^E-+J&.-P8/&MU;0LS@[_JPQ11#)#]CB@Y^cKP_:<Z
e4g.<7_.=6YTbgf@GB1TRS;g>\a]PR0)MO3MH/)(/V8@34B7b;PHT^dU,/Y(JGAg
O+5+94e/M/3Bfc2><E]J<(fJ.,[Xab3#gHDF[?]3D5#AUFHK>fR&+(AEXbE(AeB_
ZC;R,@PB88HX6[gGN6[L(]VbCHbR3d.800](F5.2RfXY(/B?9PfY)))Q3/a7K5f#
-ILBb[fJg?9ZB3O=PNa[ODA^a<ZRT3&.a9F6Q/XIDaX<ICeE[R@E;\[GZB^D6aU1
+[X]a,()([PA^9;50+PMVeZ-ON96<G^I3,5P-3P<)54/BR_Y^?Yf6NBN&9;+fY>4
?JPEN2SbQPd4(ZN+:FC+]JY\AB=09aFgU5:f2FEe;KT=@8+IK\5G.Cd)>TW8-PUE
6g0E3Y0>Db5c;8:R/?Id-Y)TU[(B#8AX5?^&OWE802edPDbI&&=?,DNgfa1-:JSb
<J5Y<C2^^:IJZCKXKZMge;04+[IYg56X;U)fVDXDRL))./BF-4U9<YNgN$
`endprotected

`protected
bGd(.Y+W,D\c&<N7K+;=/f\@HC4_L<Q+C2C)b<-,OAa,)3QZ_LR]+)Q?I,SQ]AQE
O;aI#Q+PWYfQ&V--d-)I+Ve5&a\eWP7aYRN(A@76RgcUZ0T8T1#6N07.<ONVV&;=S$
`endprotected

//vcs_lic_vip_protect
  `protected
gHg92AR=O;,SSS[X.W4V1TVH-IR]F9FFWPJ029cX^T@S)D&B,EV0-(PDH)?POV+>
;@_;)dGXR1??4?]e?fSeSUffT-@9c4dYX<Y)eGLH+Nf]JR@--R<,S8I60])\730e
HPE1\+1NQF;&DMA2ONL=NP]/+PT^YAWQ#&QF3(A;L8ZgeK?&<[X)[[D<-EfX+600
,S:Q@]LbO/IW@X-;A-a^S@#WY-:H_X@[-fT(H>&0b9GeA[@e)+ZSVTf=_.:MC7K(
&:<I15:,9I=g<g9(YXd_=<1g<d_K<6D(:XA&&@O+,+Rf.#7(e0KQ74Td2bMTeW[,
MRV9&^@Q&_ZSU?&_BR_Td6TAWY2K@+FW2&5XcC^@-9.9J7D+GA]P8#P&K)J3V^aQ
838#25#GL4QdNH1ITXI:&QQ:.Y69ZY2H?/9^8)[Wa)[>/_K_EP#[_C95-HegfOc+
<PbE+W<V)?b4^5P/M=2a_GQ3ZIHTMW\H:Q)[RVO[-g>N@gN3]0T@H;;5S6W1RU_D
H0H-S/+d+@ODE3-0]9E86f_S0W@Z<e/KYgK3MBOL?IcYRUbSd>aM][FF?TeCTZ<L
\b9PL,P?J+_B;^D2A@^W@DgfNFN_b8B/Xd0NA>OPPg]N0H3O=U[FI[EC\D(ggMP6
2,\>J,Ace<2OVW]PS(6^KERec.bdE<&1YMLdROfQe,;A<SYH-1NWAZY&bPAV-8@G
]48ZIe#f^7YM7[&KII-@IG6TH\VdNJACU/5CDQKZI?DC:L<\YU27O=W<+8:=]MUW
10BG,7N@C6M,:AR6L_CLG<eU7[=U&O,<5PC-7I#M+CAPJI1#MZdg_TWA+9/61?0)
;I]FRaCT;da,0$
`endprotected

`protected
@\+(eGeF-34f\QTbTA@NA4Ta.=9^TeIGTAI^C(7_I>[OY1APP7+<+)R<.R+Ta67A
(BH&&I<N5^?f;VGadO1QQCTa4$
`endprotected

//vcs_lic_vip_protect
  `protected
gX1<HQ(E/,.T;9acd06B2JKa+W=aP?-L9TVN5@c]cX:VDT5K/H9A&(SOU5Z^2N<@
YBEX760Q18cc,(^G1DUU2f;G<Cd^ILbJ8:NHO&]&.:Ea^:G2(W[Fc]--:J4]/I.T
BY^WH-3SS7<\c#]=c^8<JI+<0LG9=3O#6N0OCd0Y,3HTGJI2]9C4VKCVbA2GGM<4
[MZZ&6S?/BROC+S)g07^PP,P\=0G,ZRc2TAg1\g2ABR.=2X=@D_88;\XPJO\E&dU
YdNP><;:E)S74IQROV/52=NeASJF[)+O8G&dVfT668=e?J61f:-U50GH::eM+Z^P
,LKJ6d?9V0^0A44LW@NMRU1+;+GdZ4(-I=eO2Y?S=TS7GF;O(f<:;f3\,N90Z@&_
-WR>[/?gH2AbJ,8@/6RVQ1NL>OgOYY,W<S08GD-N2]7=<^]ZY>^^1U(9D==Qd6/<
/Wc7F:P10@#KEX;117,X.6SCZPN1:BWUdUZT\<RZ)Bd>2TPH\M;4.2_47DP\S/WE
X5@)<.7(:JV:.2>52XBNfGN:fEfW+\Df^2,7;AJGYb@d(P10/9cSN:a6aeHa\M\)
fWJ@L^\TZ6Pa9J.QX+HYGA<00KQ^d(<WWg+P-H3;TZ&Q;MM(:XJRc<d@OXKc[a#>
-B-F#]9FgQIHA@U4YH#MT41a]WOH?J4HY9PR37V+9KWNKBT[X-P#bUgDKG2<UL6X
2B<U>b#^UEfAZDZ>cI=Y/@3^_U/V36Lf[bQ.9M8&&a1U<7N7dga7:#M=HQ&LL?^D
AZA#W_e8>BQ@dF;A9KD\gc9b-aC=c=4-OQ99&T8\OXY5R-g;^QFGK6>=FL9;e(]_
A/eJ9XJdEB37OJWXYbfL(39:.1[@\R^HU0IQDE\88D90f8^(cP8D<R3UV4g&V]-,
a[WWAg0K,G;L7g.6T_J4/YC\CE01T\/E9&gZ&S)834ZWM8-A-fK6WSR)JF7<()8A
=dZNKSDGYAX.4ZBD\a2dK1e=J=gb__?eXHNJGeV4VFcGJdMPg^\E>5VA,J\]=SJN
e),<6>\:_\?WV-MSP]NSaXMKS1?G5ggYU:\1.1FS((59]R/>]dIU7#[6.RfNEbRW
VBPR<N>gB,4e?FSd5WfAg6\.=L-//J\?[.RM2CXQIGb)(f,+.F0IT91e.e<J((#:
Z0[6I5Y1/2g(6>TGQ_NCSV(I2#MgV5d8QR/cgRgQI1YgD/#B&(;P8>IDgc-Y1a:W
&25+F.9Y5OE,Q)I5AO>4<H5bAd.XdZBCSRGJeW[LQ/G:@_07)+-G--R3FA_bPTH(
B,9SCZb7O1(M\YGE]#\P,S5ZaA-XfKVaUg8AKVQ9CGR8PV0gNZA_>F^6eIYHT9b_
&9Q]\:DP;5G\&S6&9cc4+SgP,0SG/6&&)PGT0E14P.@=-ISQd\ZUdRC-<4?F<M,1
Bb1KB8@[0LRI3ZSBH/.YWf=.^EE3_3]gG1OL0CC>-[8.:(0.fVRe,b)ET-YdCdFT
W]94/e(AU.C/[DK#ORLJ(:7UMXaQ(_=Y6c3P)K^QM:6JU5]PU60UPOCT9gOIV@&b
f,>(1SRFBY+4(.cP((@8N6RdKD#K5GPS_ZPVN_#F5ec[I?6@8UYg.1UZFHS_Rb1]
C_]AD+63OGUB^0Y28?=@XA76cH;-V^T.:9.KU\,+-27F,0QBJ_-\3dVEK+,LX5[)
#a]&?N>&V6V8>VFQ)L9^(EE#P3GGaC:6PfKUe&=f9K(#=94-<@];4_?UBbC8fD5.
D;Y4cOdL_9QZEK=>ESU->1IRZA6A0PG69,8@RCVMQ?5)e,5ScSZ=/\&8MM<+)M5B
DUa3,O_?>\a5H@.GEF[7(\N(H[2Y)<bE-Q>/CaCBFQ?(QY]/JYC:K@12C7_A6U&I
-4JV0?aJVBZ9]]_XW+N\4:)_B40[^f,>U]<g9K<-#Ca\G)TG7&E[H0]-\,GWN0;J
&fMIR]>D=d.Wg:aIJdC^D^cbI@WGI4:]B_J)\(&8C)=1UcG]H1K<)Y0/B3Cb&AT,
>J@+9A\MKAR)/0Q-\-T#[TaG>7aY(?A8]K(Q(,FS8JA66(OXKXA[2YeE:4+dg1_5
-CGOa&JHSN#bFaM>98dNZC[\.JMHXbdSZ7QC@N66C0MbU/<>Oa;46,Rb7>;Mc/VY
^_MeOY/&665&<0F#XECC=>CfULe@GO+V/0b>.aNe<_1B,_@M^^(9TfA/;\+,AJEa
dH:eY;:V&gB(QcCEBcAeHG4\(-KS(,CB1S>YC^FTcf?3-+)eM]E]UdMMS9cDf?<b
5a@6\Sg[cN)=5\c5+Z9Sb6KT-,K4WHO2Ja+Ob#PgMB;Nb82)P>V#4/3XU4)d>>]3
K+;WN2d<+\?/M7NDJ,NK-J<X=,SWHZ]XJ68-b4@Qc0DRRT+K/,UW+d2HB\b/:Tea
=,)T@]+B8a.?</?+NL+0?HA_3(OY6/g>?4Ne)AO5A9[XU=Nc[[E:cKF8;?Z?[=TD
Z_6)_6E?A6PD-O7Gc6fNJ2=FFE8=e.>VRF)I\SB[S;4S;:Vg\e>N?BZI;Wg[>&I#
bMY=MJA+_.RLPVPE1,Q[cgTgF]HKca@T86A:LCSS<::g0D-+RNS5d2QEW1@cC8R5
<XO&68;BW[d)/BEQ\,H^59\@4a72]=[(>>41)X3SdOO&@eC,f>,f/VZD>A]X2MH\
0YY0>\S7dZ_]/<@(#QTK@dg2d0H.,XIa?$
`endprotected

`protected
)]KCU\5Q57;FgIEAF?5DEUODXK6^A:GIcaT;eV:P0/M#Mcc_&U<Y6)NN1Dd\1_QC
M\YB-<N8a\.ZKE&+5PG\O2]FKZV-HVU(;$
`endprotected

//vcs_lic_vip_protect
  `protected
H#cYE)c-,-3[fc,,DK3]V5eeW9J&:BMP/)(Lf[^6B6/<])4H686Z6([:gY>DOMKB
14VIGf1]:MN\<OW8.;Q3(#1U;]<ZXA-DNf(3eJee/(B7_Q35F=GOHcF>QB.JDTRZ
WbNF,3+F#b=M?ZEJ[/YKXKRa+EL56+6#J[E7M9BR;.f-XT@d:.)@T14Nf-\CD;bH
MVBY>CP<@f4^ZC=K.312QQ=OC&I59(74\&=@,E,L)Wc0-:N&1R_J6W)eaN,C+3AE
HOC@<GDBdS\;H;GXX4=:UgCZ+T@F]G&fK88;K@aTNR04C4596fADg0)@_QU[;eIR
I/Nc4G[B7g@_b#])MA3I+H/;#JW_]WI#MWgXR=+(D+CR,65RNY>B/,\O4[<gQ)Z+
V^OUJ_f6ZYK<&YH;W)Z2QHW\DQa#fe(Kd(e4U;IU?9M25gCHQJ5#)7\7M=>2bH,;
#e0UP[HO<ID]=ZO:dJZcc)F]C-LHX+XJ3HHY0=7;#f(<)UNFHK=6_6+VfgXOHUP)
H9T^Ue:1dKJIeEE3W8;,g7RAc6:+S7f3C^C+<c3S,7B?[9AD)SCE3Faf>I.:eF,-
F/C=1/5V1b5=@D/D9M&MaRX]MR^XULP-@e6[]>71(=g2I_=^+>=6GD:B<X_H#REa
6=\,deYB4)AaV643GED/Jd>S6RX.S2LdEARX_O<,ScAcRWM@S=36bPW?aYY&2afM
CAeYb7]2c:Ob(&5@04L1JNE4>8477<^[MN?bOegfP2F0:Y)X0K#VD/YSc0;380&J
c7/#9.f8]H=dO7562d5^Z6/@:7>.L[(FOVf7A)dMfU.1;NTG_M(G7GXN37EPV\0Q
3CdP&/AJ@HO[LR2gGJ(O6cLFeA^MJ6,^EX@d&VRY:2\,I?A8>SVT\Hc//XL(eS_=
_Sb4OQ^J@=@d@gA1daF7dQV45\.-SGf7/ED7@Y-]X_F5XC+]P=@bMD0ISgUc#>5#
>J(Fa_<.R0BFE0gO6.4;a8H\(QW7IV2Z5@ESXd0e6cS<ed@MX]F&WQ]KdS_/XUcM
H;gZ>B6SWfA[1K>HBZM^F5Q4\Ld)8#?LZ\bP_+T>UHcJ,T8\e=c.Bc3cWM>TX@YN
aDPLX[=QU4.AZbU?_--b09.aAY11]_[+8:e?^6L1,&>YWeL+XRRA+]XZ^<M3_]33
OR&]e^JKQF4bV8MPWET(BZL_YeIF^;3JO\H6e9caUL;_-9WEL,)9I2defQCOF#)G
Va;^5^7/&6;=b/TBIOL,XDORefLHb1A367B>?:7A++f;<?2&^c&SGY[9>Q=;HI/f
[AF4B5.SRSFeXUa?-3B@(5&71Ie#GBEZ6J7222P\S=2B/\e:]Q?5c=g?7.6Rg)3(
XN#J[Qg>S\\@GRAKg?LDDQZW#6PFQ3.>_CZJI)TALBNFE9:O.?QT6dXTaNBA/ZQ/
AM(ca+9L\3gPR^3./>K4VXCBQB8,[+NM>_Rg3[_7SBDf>&fZGR-8>G]TY;E?XJS;
)B9XA@<=)-b,0,1]65#E+Jg0RJEKIJ3FN&JO55)7aFW7_&-WQBg8Y.)JTSPHgA_U
9?\U0P_H34Y22HZ&Y#M,[VVbb-14OYH.I?#@1@-1OgEX,OREP5aTR^3.=Y9VO?;S
WMeP3V,a^GRF_&ML109)=:OVU=?D;,#O8G(2-:BV8E.(B/d<63::4AF^6:SSX4g&
Tf?<Y,Ke^G0G#V;QcaVAM^aLJeVBDbLF?&.-,@/C]f.I;VH?g9VgO)W?IJ6CG:Je
4CQ7O+fR^<QKcIHO5^FAe&+e392&IXN3YU2QHD=OD#e+Q.E15Aa1E#IbE4:CgR<C
XRB00)SKV,2RHWA^e.SK=0ddI1DJLB.MIN[:B^8.cS^?ILffP9VLbRHZW[3b96PP
<-PPTL;;A_/HaC>4K64b:3-cNZ6&WN1Q:NK<KDHcdJK;Q6>]Vfe2_69GeREAV00V
>&EJ4G9XFGEH-YNCBX2Tb=Fd_VD-]aRB#b_/.]PK_6HIJ\5?RH0-/^KO,7#aQL&5
C9]#LN4B>F[,C6UFcZ(7@B74c.Sc,4AgL6d&,2f>_Q@f2:0]WdQ@73ICIY+^;@V.
^B3#EL66Q\?J)2aPfcU841XX29.9OT^4@5WaWJ^\.EK/<+7+-S^MNSAeTFZ/fP66
eJ,\e6#OD^]V67^;LDZ@XYI_.c1(:A9Ef]/0)L9f:NVDX>GFMf0ERUJe_1dbJ=bP
S4_)GaP6<Z),VQ[D#)gKY:[C(G1c@>J<)B.Hb^)Z8AY-ATgGd]&VG=Y38XR+>H]=
-/]BW#AUZ=O9W[a4_:4MTf74QTcBQX&4C4NRfO^-0,/9/B-XE,bI1;ec]42E_(dC
Gd>\#.&OZGONRKBUZHZ6&WSI<\0QKf&HT2KX;d+0;M;M\c&6\]gQGE.b]VPc@3Uf
&H3,g_K\7(?bCd#CNMU#bO31-YV0QZ:I1+/Z-]V3B3I;/-0FcXC[K-P2/?TUP+Z<
L?=_=4@N)1F9BK,8R^;D&&\]7fT/d<cG#;ZgI?/V^6ZORM+,VMR7:_=B@ZNME:L0
(>[b#<9Pa1MM+)>e6c,.RVZHQZR?>Z&::?ZX(;=#YG[b5])-5fV]:C6PPdM&a)B(
EV,Y;6+CFgBW,N9]\JM3=>P]+PJTZ?+A:MCg,Ae0807):?#QYSN\@+UI(4IGMH+.
OJ9F,WS<DN<QDN2;6JQfK5^,:+BE;_PI/DNbD[&L1DOYP-^.]Ra5c,6T;>eXZFFY
4Z9Uc6J-J-V],\=_4Y/9A8=]E=g/eE9g-)bL=OH?(4;4@f>[DXgcbLF]Ec)6e2)I
&UTcfTUc=<O69YfJN3TTMY^HC:OISYKgW&X^]K4Maa:Q3]A-]V<&WXe]a5^9W<Dd
IV6268X@PEYYJ#I+^@aIbI4TKRC-]J^Fe_LH[70<6UD&#b0/+VCN<&SM<4MIe5PN
A1)3-cgb>\^T8AGGM-4Q^&.3debGRV;E)?8T=;MA:Q3b279<;_@eKc?-#O7IPYa2
,1-T??PSH_;1.,55AO147:5405PD56>FLUdY1AQCS+]AFcII?2[b_S:Z6,3EQ+.=
\\8T=.0EI,,f<9E8J3US109AgQfUdZ;ZbC4AZBWDf1g0I^W?K/.>(R(:Of215/7F
g,J]RdX-M0He/>[0R.(L0C+FbNGf92)J76/gfA]gf_^7a9SUEg)T2W8Y-P]fO<G(
0\N;IY_=]_G_a16^U0?_FY6eg_;=@c,aM\<WTU-PZBKO3<BB?UQ9;42.I+EAI(CM
DeI5ST_,[>FE)>,8/HB,LgQ7gDG)MAD+d>?/G^ef+c6R[QdPaeeY71(J/O<+FD1C
NMR,@D_._d[LaIL[\M8;a)/2(#W)IEWJ;8ZWC>5.D5JMCM6GY:A]R_^dV<D3#HB@
f0W0O/+5\8WcC1-AQ@Ua?9?ECWYC.15d>CCI2[BdYQF8VAb)@;0Y?IR,f/YJgI>W
?I36=dO:\bKFK3Tg?,PLXA5-J\V6R]6@1-2DYG4&6)NZgc\R;BFM3#MDV_6<_[K@
fIBXZQ?9HM[(3,[H/?,9[A+A#?)c?@/P3I24TSQ^+)>e/:ddeU9_af6EF>)D_ZZa
;+<L2(E+LCDXJ/6P1fIe/(US5BGFYg+ES6bLa49)#UL59g6E->D,TQG_Va)W)3,d
@;/YbST\dQO\WM-A:Q>@>+HcD;>L7;IfNd\JVOY11]@CfJN,_]_@/,M>7J-L111Y
Wc2eHSPE0MI?fRS_GSLOS^aIAB17=F-eVb.6Q@(VC1EJZc68P0cWOXcSC0H)1;GM
KR;[CN1J:^GI8DYc9KV3?fYGa\eXWKE:39=1YNNWQ\)_>@M/.X.6T9d7E\>ULG&^
&IKEdY_D4QBR,\^Sfcg=g?/dJL:-Y>A\D_[797MX@C05gMIMMa=JCHeWW5AF9-S[
Z_3@#CXcLU476C#0OII#:,;?]VT?RU35B\[?5g473c0/.#+>I;(S^YAP@)GT(#Zd
gKY5>3X\SXNIT4GIa4DT(=/H727:<DZJ]32\I)4#gb@Z_e0dKS6XE.QS)/;GI1Z@
L6eY6/N9O>?<,QY@EQY@/MG5-Ka:V+86eZ]09R@AI=<D.,221990B9F<(X_cDcM2
/6UF7?^d98Ra0_&8D/6VJ:Da[,6I^e48(^FVU3Pa@cGC[+N3/2EC5=PDH)QB9Y^:
__H^.#f7.Q1)De2?]\_27-0J,cNP+<I_84?<F+J1UY[3Zd+W2NKMV0O]FZ4@b6S/
U^;C8XOBb^e)-Dg+1G,EOZH=CT=WM/Oc59N+S8,S\#FLO4.XbKHJ=PC5gcGZ.=I?
\V=B+GPXXLD@G^NUbB\.@+>IR]XKT=@F?:)ASbGZE:eeUG,7aP^KW(WdB+<C77F9
8;6KKXX#O;[&S5I@D#8F5NDZ/8<CH;#6BNNgfDVXS?-@C6a9@f6e@c-><4\B^YE<
?Y=@./92E_<_B(XE?>.7T9VN#GNe[9MJ9AD89^+>.U_LV:^dO2_(NgJN7\_4F+&)
<;b[,7c#/GVT^WHG:@.=B9<B\EJ-\,@TR9U^II3_T[IKJAf9#A]e+IFYB0L,EU9K
]:Y><HKK?[]bMFg([UfHN-Ce(R#@1)ZbA+^6MX]H@e4T8SLR#^bcGfWS7_H9_J<@
14K,:gGG6H@[cbgSFO0L37aM/XZ/YFJ)GM&/C4=-\I?;:T\RfLKc[JE8KZ-=Eg9(
U?-ZM5JNbOR5<UUTPJ)f/5+^I;Ce\:8FVSdR\5#LZWDUXW[;>5Y4Q3[]B-/>gV/a
V(<UB5+?Hf;QTE#__:N8O4@;_O7E[#Q5^T6XR4+P?S[D[30/H+D&V7=R+Ye7_VB)
O5d0#Aa>aa,M7LRZSf95),Ubgc6I@H&4FSN/MfM9O)7P;33/cXH?^DRBU#ID?&KT
LUbGYceJRC3#d(KJO3K9-AQ_[N<NHf&WM7HS6B#_N5L00HP:#:cCCYCX=HQf+UZ5
R^LR<HXI6S:&_TU?#TRM(]\dUG+4AM172YS+#ISQ1;#2IRF.W54L]P_UW68>9=I\
GN;GZW<Xc=[A,\e^_@TgDD/.8^cVCP_cR:P+5E=NDCR:Z2a9-=&bI@S>^870#+g2
)X)[:6f<HBDbTC+MWe454+3,bK.8LRS7Q5gM1E885\c]e1)g\VfLf01c)17G_<5[
P=Ef4RQ9)PPAPI6@5S6GWG>TS^F6a45XYWTH@aUa<L+BI@gf(^TG[N5DfQe99UEL
E2Z1C]f-G14c^5[QN36OQON^(:IKedR3CT\F7@KUK.)WETKFGT5+g)F,#)Y1;bgK
.eENVb0P;3Rg>G(VB3=6fIQ\Y+<2a9gYBN/G0RdQ\@[08YbFL_9XM9#&RcT+H/+Q
CaH5AEXINNGG2Q;Y/-H8^^]T6F/JE37GO;YOM_1U#b6);EWGd[Y5Yg;d\b-95FO1
bZefV,<)4)L]LRS=\<AWeB0/MI7M+?aY.OQJOE.5BOHV:T2eV>ZYdE>T#aE\OWK+
=\,T/YBgP&1L(fK;3O^VR5>5cVH9/@_8a7(=.a+0+A<P;[O37EN5K:8_D-4[4F_I
FSL,dA+XJ5928,C17)2/&[W)@SJcC&W2RIeIf?NeRRQJX6>6>;Q@UJMY/ZBc^d0f
.Fb?/aUNR[TB74@/NaSU0Z@5#g^5SF?G2YPbO>C_^fe((9-8dV\3U<5;EB]L1;Hd
U4L9J3_4aN(5gf.?ccZ5MAWV+JFG^cUDR:X1gb@U94/NXR?CVQ3eRI?SP:FRF(@E
&I]XE3BIN>(MM,6[:^IO.JJ9=99O[A&IHcW+R5.1N&,0LV#G43=(;VD]453L?7f)
YIDd?8.NFe#?Hg1-^&IA[364<:I1QMYcJXfE-^VaaV)4gK#_^e#\U(\=2-1_ZMF0
F?>A=^EENH0S,2K)BO<&>[Z#O8X()Gc>:VfXb^dbU2dfL99_2C8=8D5\6g(+5P6E
>51.Q:EceVCbHg];eGM;75NJ=).CeB4Y3d&S=fIg^9/IJ;HWdg]>U4Y9U0]2A5&,
gVI//9bG&PL-e421[XT2C0GTOV?.]Yb&;K2<T1eS2#c6)L^-@cHfHNI0P7#E<B[0
TD=CcL#U\/OWU=K5DAH859LVc+RZ?ZTZ1:2S)3Y:K-8Q6#?B&O9Q[L>-MfBKJN8O
15A_JR,=R@f^<0C)9@4#Da03/(9HOS=CV8?O0)59)PIEFE\CQ1^Ce3LH?O9+@>:H
AXL(N57_V8@.K>L5@&ZYT&bJe/aO;X3ZY)c/<(-Ne#8C@8;eZ<MQD@d[04\U]bGE
[:4H4Z#g4&FcYA)F\+IRG1-JOEbVG0?6;gf,_>g0fVRgOT]\_PE?(WbLD?1?eGfb
R.]L,5<FU?fb7)=7cdL>4O>&QT)-V@O/VZ<YY[TTaC#bc/J>PSbKEL>VEFA66U31
([UE,W&0&RgHeI=8P>fYKJ\g&H.Y_Ag]?#O9<cf0VK+V^aDUE<2?VbE.1R?S8)Zb
QeFM>//IJcK#B82&NK=ff06&XZc<dIA>.F>GK(N?JK2B:^IIQ]F-f;,4#Q>8CF;3
;M[#6Q2?e2aeRI</2M/d#2cZc0CY(e0GA4a/L_e[MVU6)0;^=M9&27CB^O3gO8S7
=\3f;[,WE5+R@:>&V,(V;0F;2I#H1;<d]1Q_7A>EC\L9Dg\@3e39]>7^R:9cg]BN
E?;[TE[X2F?g3K:AH75T&35c9Xd)0LWY[,Dda&]/WGY6,V]4)TeKN(2&(d<H(RWH
JIa@7LM;eJMO@#f9WE7XZC23,\P516;:Pc?2KGC;PJ\:bRd>fLW-agc:H;)cZ7[Y
JEK:U@56A+\&CG+IUG&RL:ZDbHE(I]42>9YXLfS+[3HO_E<[Q6g8/eJC)W(@?].+
,9+cKF:9<X^D<\3B)WDfO\?\Q6O8g+UTC]PaEM_AVF/?J/1RVJ3F9P17,eU@M(U_
KD6>-e8e_=<bRP4S_B-,P-Zb[Q]\\Q-?/PPWg-Zf+<\bKeX+^>]QS&f[E_BZ3X?6
SJa^H;X)U2XYEgR06_:5K7ag-TRJJ/#2G;]L[[&IfO3(Q4=E5GE8S2\LYM4cLUTK
/gO2(?KZfJOe)NN4]R@1SbC4J7&OFegA@X+cXeGBAGH:QR@fR@b,W(cdG]Ae)FVN
:L5TS4YDI28S:.<RG^YO-_E:]48##N<FM65aVG>29g)8:UOS=Z#.\a@[7WUM/;F-
S7O/W70dY>Cb38J6,O+HY/46UO>N[O]/&Y+;5+XCM[9TVdfgWOV.ZZC=77,TQc01
2W4G526\0/UA.agK5]\(0eYcS/d)7XWKT18Zgc>UG,_PbffI,OBcOEGR52@7MKPc
#EeM3Hg291=1)D;gc4UUZP<H9:C>6YD^/T]+O^Q-W(acG5NBVT)[4>>_G^)5[(a3
+c3YH6B20c93dBJ^gZWY7T\SF^X>5eF)7_^_;@)_7F7XXBY_CDV(/9:]SCV>U_E.
8fHb?\?3#1:/f^0NJdcZ<(IF?W],W;E?@^YU&S@_a]<O[WaV97CbY:^44RZM2RZa
79.OJIV.&KDY/C2B4.OYd+-9.V6f4cM6[_\066F,BC.?&3a<=3RF@9A1L>gaXMR7
2<-QFX8CQc;A,F&g(0>gA?b:c8F0=GJWG6(,AUb:Z,=Y^JCH6C>6\If-RL9<NcId
QMQJB@9,(.&2.#39D-JI@Fe:Jc/)D(\^AU87[&(=#6,<:GY897?EVX],Z2QAS-1G
Adec1C=C\K2-].Q<XQf)S?f3G?Ma636+4EfE4Y=,XZa;9TdcKe3eN#(Q6fbY=1ND
A^egHMbJfdeK[A@]4N/YH7A,[L^+_+KK<1&4C\e2DfR/TOWG7,=]7C,=EHL&N]8f
PI1IW=f,gQ,\eN3:19TRMV2\S<BO.2?cWJ7bV@<RbB(da(7V>@?<0:PKBL[,);f0
FPH\=:>Y;7[ZRD1JPRM7cR=U4K^CW>,+Te_3YT?>fKO4VQU6BS>GXN+0PM<YLf,K
BI?;PO([?YJ#(8A[P4L9=^SVCN]3(CB5_Xcd&4D;JXN?_adKS5-+A2J(9b2bUeU?
_Y(#6Q7S-fdX^g,41\APEB@b]5\:DW5J,:JKd2J95BMU_;aX0SHR54ZQE-HFWEPY
]Ue&:+>GV(I\H<(18\WQ0Y0/R1ND_^N9G52[L_DUC5Y)G/FH^Q#IDCG@SS\H@Z]H
A=?)J9c0H)O_C3RW7C>(>Z>[QBJ9.bZPNFaLC7_BW\)Z3E.]-JgBBb.e?/4G4XY^
dL2&2O_^P9DX1L#:<+e[e>J[fWMLOV/T_MdV4BPDZIU=)H<A3-4d:gMS;H8A]+UV
X;H>D4(g/d3I@;B1YI)-&@a6LFVgUB\<]CLI1]V?-+CDWd,GOULe-ZK+1T??M_-f
\KR)RW+IWQI),0(;c:QCR/,QSY:GMR<Q:a[\Og+REQD5b(?9R3=XNb3fQ:<CR6[E
1[&7]VUd+3GG9cA<E&\,EY?4e8921I)QK<JAWAdMac^g,b+>?d4@_Pc.IW^,gK5.
O-._8K.S=gd]Eg:3O11;CCZ52e]Hbe5?L;_&LaSfC2FA/<+>YP+QK;QSaf<[,RDN
OP.9.@0^4.egEGB&XbU=KP]<N5]U+-C;R2gcf&6JMG#(+ED42VK>Q8[ZW22:#)=8
>>I1;)_Sc5XD20WA-F,LDD\7O,J-J3[C_DZH#F[4PF:0F)=ZA:=1a^f]fJ(J)0M4
Q76#E0+).73DeG6bR;[,\LR9#2=?g=:Va;@D\Fe7JfZ,W)Q-F7+Wggd:9\QOPXJY
W07S0+Sd-WgU8:P@-eXN1JJ3VfXL2Nc]:;g_2]D2VY<gJa<87JggB(N^2>XELXJU
#ARcT.B3N=Ua4L>41KBJ\EI>\#b&@;1R4Ef?[Y)+e2)5Y<\dT<_JeG451gfS_+,2
8TPLa3eK_N.5&AAYK2<&-M5a8ZI;2aYT^T@O+C[R>c;>F4.UgW5G<D?X\6Ce8<VZ
P&8.<Y0M=A@f59.)[(4V3EG5)4III]ZYJeKOg07Ce^O(WNMC#gZe+7FOWE2S:;fP
(@Wg.6XcXgLab46)\VK8L<BY=TXFI7Z7C+0)X#a<1CX&Y7-JA.aJXZgEKMYG=)2#
]cPNa9]DJW)K&YM23/L;X3,QTVf5b3e1>$
`endprotected

`protected
X.0Q/)E/XH>H4Y(>Pg6FGA,T[7)LOEV?.XHU&5-8ENAVE##T,a)-))0FO_.T8<FX
T_I,7.D-L9>4:Q2YLD5HWK,T5$
`endprotected

//vcs_lic_vip_protect
  `protected
)#gNUMY4C1-dTQ.&+aUPUd7Z-591USZ9H0Q?\\d]&LNX?e)#_7+f((-VCTeBf;aQ
4S,#E_+[B@<=/c,W/W0\UMDT77DZY\D@]4L63LIX(G<O=ZQ(^OA@d4DR8gE;S1B0
K8:>f+_VAVReJ&9#,L]3]7P6\H(,3e.T##NI0:#)C7]T_Wc&IMG[NJF^(^A15:E[
581.UH#8XH@5JgA@6TD<9K<B4O<d-43YV[R=.TcYJ)._843;[EVQbaO[\HeGWFA8
Gb.]&a4/bJ++dI^TT=B1GYE^S,@9RH.V7E]/aES47N93Qe4>M9g7dB-YcHO@gAAN
Mb&HJf3_c>ILO/)]1[N3(VU]]L^?6BL#WPT]e+a[I;.[J_b7Vd#:a[L]Da;.C:,U
/((1<;7b2P)ZY:4G3WS^@c&FP0XT@#9WTUd/H=,O+4PV399aQe/Aaa@#F/f2TcOF
cVA[DU)5X3NS(CKV3dJJ3\8g[9Q^ZO\.[-6a@K<bG-IQcNCB_DD9aaP[c3&c6gD2
,L8G.ZP>)N,/AZ><TU/P-\KUcNTFL)DF]SIN<&V8)I-LUbe&7_,2(0b42V:f^(Gb
+6=XWbVIDI9Yb5g;0cVeM;<#[66]WYJF:@>6D/E2_Z)5K39VHf8@b/DKCG88U\G2
X[\8GRgWS-+2HeVGW[Ug+ST8_NFH:?a@)HRC0V0<>bLF(SE<H0TcONH4-Q+7(F,&
D(4:&O0RR);0N<\E,.C@Z85C-ZbS:a>^26AB+7&f\]I./SM6c?XcI?IHNG6JS-K_
,0Y(_]<#Ub-\ICU:QQ5dY/3XH9:/J#K=CSG#[a<fKGgE)4K3WVQ:YVUB?NBR/+GS
=&6W+HTcZDC-LK(V?S=<9[S<ZT,+bHJ;c9Ie5X8@,ECOXO0QNGF_^VJN&BdS#Ad_
;cQ88#S+27+G);+4#)UQ4d.[<I.--B?G8MWS<dE&&5cbM<DN2PSAE0E.W)2Q<4;I
<gG+V9^Jb>[^<>#S224?5IY<[G:PfcO-1_U^@U>W0A/=TH:H@eJOPMS1aa+RV9OH
<ZBR_IMJ3bZG4Xf2Jg/Y<-Lb/1+:SX_0UeV6;FSaP;ad#D_O/(a<S\cYX/EJ\KO>
GD7F<A,)Pa<Ba3#\B>1H9V/UM)@b4M]@U[?Q^X(&;M7S&2S)RJJ9RW.6+H]JAZAP
P\)],21RX2=8VY@TE?CZ^]WC/_[K3S^,F5Rc7PC.9R4KL)5-80V#>7_+W(X?]-3+
>N31-Z83CM.e=T3S.Fb8^>NFU:MBRF9]RY+gD,M+Hg4a8e[VQdg>&XVDHY\++F;Y
eZN@Ad8(gaQ-5=WVKT3IL_DC@HKCg:SKJ<M^4SLI=_TIg,#(GYZ#?J@HM(+TTa+V
:.:]TR)32XE=RFGUfYaZD\_&aV8VaS8c+a,T/T8PM_KPLg95[IFZJ6;0F0dbKCge
KLUe(6X,VfUeLg6)ABDM9@P;QF_M_;16<;KXbY:7C8AA#U4AJ>1CS1EKNNG_=LX_
I27?LB0G:EX0D=D-4c\R2<,(F7^;Z14S_.B,^[.21@K@);(7XG1[(I4aK51_GeT=
S6L810O.-V.\Xa(V9@-(U]:94VBK==aIe/;L(a]];:(1KgD[YFZ+]4.NNN)PPeBL
WB):9D(T\Q:^027=Y6=9C\.bI\DFJfQaU[+&2T]:/AZV0VG\_Y3CT6Zd9e,38<Ma
a6R+@\1\SgeJ_7f)dU\N:^Rc1E)Q3Sc4DBU5RdDE5:)E[PWZQ_OT<A#cb3>?QW;(
d36.JR_6Q38HCHC=U4^8@<8^?6?NcD=9O==+F^M,;+B^MAAA.LMAF-\MJ^N^#N62
faM(VSSWZS=\_0bJ8L.3;=Q\IY_;H[gGT6[K[HIMC(J&IK;66U,.)@?T-7EQR8A^
#M4:WKYa;&=E_6_:CI]UHI5?<96T]g9TL/PP2EP<V@^eNIH6#9U[4^^5N5D5VST[
g:KZ2S.&Wb9ZeX>JZV5FBWGP[^c+YU5V2/)#O_94;&\^@MDYM:cMbN;&T#I[/7AV
(-2\M[N@?VNa<+3[BOZ0N4?>agaRX0<a2g<^ac7fdV@X>#feW4.-UO.:IG4TW^M3
3H+&1EdK/)P^-T/9Mc2Ke_7DF-HH3YZOQQWSW,XUL0&aEGY=ZEODgK77b.DBW5G2
GUGKdK24]ZIZa<3L;GbCg\-Ac2M\9LO7+RR^XV/9OB5?^V@,5aL7JBc_(9Y@DXeL
>5Y[,HQ8-L4F#LEROS5]W@:5&eNBS\^Ea@7304[N@8;=Ae(+SDJOR&AZS^\)62,V
BJE<TBJC?8bTHJA2,7IaQQKS[-AQF[9[]0YWESM\7\fRXCRY#_=XH[&S(?.<Ha=g
UKPH\2X,9La\R9+(G3.;&<;7UNM9b^fT^E.ERUGKE(5V,b>;6/<2fV?-a^Be0[7?
]H^R>]N>>dgVd+Q[=RZ9,21(Y&U6OG3b.6D#=;6BHDL>=8L0\5>UQeL=[E3I]QAO
b>egH849Q+XG+@5LA2_>10b,<@fdGeD/PD^5+K)9\a.a3;R8\.L/N.RHJR(IAE5E
);g=e3,1-&>]g@^Q:4Pf:8N/c)YF;\b7AE2L)(PT(8>X[JAZV>Wb(@WILDKX3@91
CJ,04/K/OU7:8DINPN<<SBN]IC[dX_2SfR>292Ka&04AN5HY^]A^)KIEJ7,b/3c/
0&ae6I32ON@;IL+:V]CF>HJ3-<(?eD9Gbg-[W8BU1RR.b5RV+2T7[::R/W-26+DX
C11-C4T(bFeF)DZ<-]Q=W]8d<U31ZIcb38]&K3AAJJX6Q\:\(47ZgLW<HC^).Z5/
@-eWBO[Bcef)QJ&TK5VSdB2LOQg_B#;\G7Ya6-W544X?E6KgKd98]aFB/O4cN;,O
I8:OLL),\A9.;N\];_)VO_W=E4b<M&E1XRcg?L9T?,DeYD56LDWEVXC9-Vf0e:cO
:;f&X=V_#,gG2a,caH:1=T[^R4@^2S;/(L=_[M>^C)Y7Z++GR)bDMbGFG>,.0XK/
Q/A8:Q0_V=d>EEf5V_[5g3PbGM.43F:)/;4a-[3]fEI?\LUX-.CdXPJ;K6XG.[Pc
<EKO?]B82T)ULJdf6VY^c-bR^?c\5[2MX^MZ,BK7/E64_9OcD,<10BP5+B@T0A;1
0A3C7J?0,)ZaBT9a?77@-(BL.XGSG6Q^P>-b@KSK,:=aQ;\e7155>B]=APS&/5S>
Rf3>J[7@B8:6[Z92eGH+VBKJdR&+Z6SRb[2;Y33H+b9BY^(RSP;aP/A5>d_K6/c0
CD[X4-RX1X59S&+;09>^X<RJ:LAYga/_gNS0SB?H-HGCYK;e[).G\N2@I,+#V_ES
@b&a6,d4RQHPg[,^gM/fgXNB#b1.eaP[7\RTQLU6(PT[IfFWL@MgE0#]eDYdX8cA
Yg_9aRC4H[4P.e/,;ZKRNPfN2Qb8G2c]3M24+=K/CFD?NQVW<-E1aWe,Jb^cB(&Q
L^)EY4[U3\.:L3.HP9JP1EX0[[0ZO[bBF,C&_6(8W\b3fGC(.)26[TQ?QC:.-eHL
X+:+0)&SFFQL9K&1gC/g4<P.B\D1^,Q5Bd1COF1K5;a(J]?YR4[G6WN85F@@3:(0
NSPI4-6<g9.a^C;H/-^gXf/P6BCdKgK6M.bA&I(DcV_WMOgDH.>V;<W8QF4BQObL
M0EecdSXK,dO1&Sf?ROO.@_\CBB(aTY2a\^fE;]W7PcO[>V]W5V@Z(6L7IWG=/^a
4eVd&>VfK\KEM6K4EHW5?042#&0Zg0S1H-M\&C]69BfV+a<BX\=7[AG]1SJg\J<]
D[UIOIF7?DK3g5/Q7fQe;IZ^YI+[_CbU6=0F40YP)/2RO2.\a=dGY-&fAVJ2.-HA
L/\CVF2?J=<b&?aNUd+._e81]A,O.^Wa6U.T(#g:#XR4W[cVZO]][&Gg200-gL^+
g)H&SP_0\D@^]>Q)A6FTJ@^fN4<WQeC3]1+?04(8f]@D?8])8W5ZXgJ^EIZ+D9;-
&cC;8=g?a3&FP_&.4PV]&_bbLA[A\4aGS+UgfcY#G+71(>I53\=<O&aVW6B05_+<
Z>H9]R<2:.X0TB;9B7\OQ7FK=?T3@BJ84-8MbPVV5^?#B4AM6_52Cgc1@60baWbI
W((4eA1O.7>YgI;;I5_;Z(=A^;E=13NTDfP1A>]5:X@,fa.&GaR:-00/YM,5E&Md
8b21&E+?<@WY3@<\V0V51]_J<\WM2V__T]12T<RVJ3AI+-G&;>P76DB]Kg9+R5U)
3eG;?54TO,]IA:(-Z[NQ-SV1MMJ<LPXHD.];:_J,NV;)7)-O;7;J@5ZT4GV^,Ud/
KL<_G@PL[4#413=2W=7/2?/FC74a?=D@9YJ&O2Be_O,(>S)-SP.IJU[(WA,=:_E:
>d53b_@F@/JI2<Z6:5gT97]PSPZMfc(T-K-5<>6@03a\aGR1WU&=dfLH]^dJM4cP
-&SCQT8/G&Z+b]1d1Q,/92=g0<2(3+3/BbW1e1L6;#B^-3XQD/C&NA?f86T>DC-P
GXMJ29Y4U,S=R2?a2c#2TM@;>JYG0D0<5.L[c:OR.M4&Y_aY(M-)#)GGWIS4PTdE
G)aXB@XC0[/,H^)9-:BMBf(QfdY:Q&KX@M@E2b=O/#&<]VVAVK4J^2F&:_[FQ4f;
eIQAcAY;,e.Q.\0R)8H_Ref(<\eW:O0-bZFD7EU7S,.S9JROLF-C0E[Q.AV<3[g[
6KMCCQfR^39<F9.L8&dda+EW&0UG)[AR591fWAad@T.V4)YQ57^Z23G-GB@J&#@U
A6_.3Z&.69QJLF,ZK>O9)8gN^LdQB:QY<X/3>PQD-cCP-0LE6KF^A50OSdEVN\];
<>VNMQ7EfBVPF&#+eUSOe<.E(?I-@c@7BAR(<Za3?UQCA:VXLR>00@R_2AE?/2@I
:E&FFc.3?WOW1Y^#>d/4B0\gDC08RX#)JIBee?WcH72gWYfI&9f:3(0:.7ME[@:L
4e>>WHfc,&#)5710)3QYfBSe9J[@g+-#:UT;KBXcJdce7cEHQG2/W<U,bC4Q@6Mf
N>a&&O5R-,M7Q:&Z:X<G<TLNAJNS-[72=6RWZ;AP:XB)ZRg-AFB;,IbSRCGMUb<2
TDC;:V&Md)G&eOTf_[AU5T^O?OYM\6+RfRJVA-U6Z/)S+7YM2#Qe<P3]8WVN&g>c
K?=S-=HGJ0Z<H9gK0@_T+0SOW@aX,(=ME=9LT[^:#eM57)(gS#=6b>Z,3T<[Led=
7SHQK<A_ZafP53ZZ^fK,@+FTEM768,ZM9cC6LN/C\MTcURIF;[6XdQV<5fM=^_9:
K(CXaYB?WHNUb<3?_)H=;O1[3bS=B.457T+c@&>4WL#BXTJ<:JA:J3S1[EI5WXJC
/PTf,0]>,IC&XM#Td94<SRQF&PTUVAX;DgMdXW_(AVTb3Sa/b.IG(4@K&MYG#-&U
4G0T:0R7M.E([T#B[59/,(;D37>OK9PSX?cIQU5T&225<_5(Y4J9#gY#4VBI-CTS
S+Hb;=&Fe@?)g:dc]]SPSN3TV0:&-]O;,YTTY:aV_QE7CK19gS#Wc(cD61<a4M>#
IY7U(_-OVHVCc489-6c,6OJTC7@f.E30EBPe#H-a-=\SL+WNa?cbc;4M87GS)@/-
4..af_X^)1&8V-K40#Wb@=b&+F6]=AI7e7\43aN.fLg0,1]@RUOF#/7b@6RFdbSB
+\512PY+2+-(V4BD5DXE4,b<.XO]N@Y;1dZFYKO+>@.a)A5D?M&MPSO8+7)_GPIA
+\]N&:N3H]fN][=16[C/,<(9eKKYRCNZ&0&AE>2FDc_F>^SgUQ@&21WHd(,W2&_[
8(9+dWZ)f^78A5D<P:@MR(HK?OBcJTO2Ea0Tf4=(f1QD&WC_C#e;OJ0)X.>V60dY
/5db\)N+9R]:a]F_NNX[^#M8/gQX><<a8,9ZEX3UZ.7eebN;;2&O/@I2I06Y)QfO
NLA2&#?_NV/cVb:BQ+[1EY0D+e]F&gXT\V3R<aXCa4M]06M@U4d>Z4_MF-Z<N48R
2dGATbZ4J^#I0SfAGO[1RSaK7PSdER)_TBTKP,Z75?4a^8XLKf3Sc#9FNC2=LQ[(
W:_+TW9X[L>7BY>22[dbDM3TD[ZEf^baX;<7]dYQJ&F9_>OX6HJNU10S9]CIH[Nd
/&ZEM8de>+c)7HFCQ_7WUTY&H8S-00E1-/G]FXdVccYg[706ad_Ig6L6M#W>-8c(
Add:806?V-g/<_8CY:@\LO;/EdW67+D[[=9f-NG&a0681J<cO2b&H\[EQ(J^[O\d
Xf-gDbGI:78,W.PdI4YB=M@KFIU@>[U/XB7f>:/5a>J.6=).[X,A,YK\A2:61ZWU
?bSbH_(f71SJ&NJP[GP=EBeb#?b=g+I6QK:O[^G,bYcYAE9&:#-gOc\J/FN;_F7a
Q?+Z^1N7MdQce>RD[UINL]A;F22I.64^6b8NT_2a7]>#\_S=b1I.W_@;1,Fa:NE(
2_c6gCA#?WdQ9@8>(d#;OI>JX\W6<S)</G[;9VW#>QB6TN<eMH(M+JXST?77[G#O
&^J/ReT@0N-VSH/0.:][>XSFT.-<c3-S4DD<8MUM:G6>2,G_^-L58IR?+769\EJV
<9#9GVN(+E&bgI#K#TAO5a).\WJBC0FN=<d:QG?<HN@3[[&9274F(Yd6_HL:A7f^
MEVEg9fI;b(<GK&D(A#4H\9&(R]J)[04g>0f2^@6#]<L9\91?c/1)Q8T]Od@F?6Z
XdV9+7;:A=X)^&VYBX.@3SMCBg/A2PEH6#T=&PC6_CNO,Qg3[]N_.^Zd-0V+=[0g
3[;eUW-WBb:E0N+VPd<eGBBa>1QYaU#fbDG-B^H9aL5+I,);\2V6;:@=GL3HPW+1
HY&WUI9ZAQNBWVC7;UGG1@,MVU#+W<Y@=9#Jd(eN#LfcV65<_2TX11ZZAdN8&A-0
f_7cLeX>FY>\f<T8I[<[CF^P#gb,PM(N5+[Wgd_1DF\-X/\WF]X[^b3V3^X0G,42
7<)3\J8D\,ZF_XV&CHcY(,]PHX#Q67,>3C.0N#D6RW)+Q5_2AABR@3NUZ;<K-H3\
H?(P?GD0J1dNc7@X&4ES,?_&QC^fNF8D+f,A+?,]F<.7LQ441@;#PN=_J,-5f8G<
EUgLWGH0NDC_036BRg>19&aT<b+HB>Q>O5Z+I3A^@57#UL.94CYeaO9YgO7M:@B?
.9BB^\:78BTM--OA=f>e/&2<254/CU5+RDU?25-B&]7,=[0DVa5P\=e]+8&g15bB
+YZd6VOW)NW3V0SgQ\B,#>R+N23DEH,KQPA]BRgL;,J-NI358Qg^W@gg>JU612F>
_09.dC]USDA^0CeFC[gB/5,R^S(W:a4Y4,9Ygf3c?5bD+dW_X^F:1VT-]CSGR6^@
5>Cc9GB&1\7bf_<N.=6(OR,L_12eX\:##,M5E^edgHf\4Z/2;49b>GbG8.8HTUgM
OL.[Xb<H4S9FCaVd4GU]0TI.(1Y6T86Y\V2B@/D2^0)de/#Aa,2-FIW/Yed)YJ^-
Y-AC]FgTT7&g>dQ.XUF>ECE2EdA6(G7+Oc0:7W(JB,+\,_UN\X0H/@X0)9Z/+>3A
:DL@35GgaIWbJ>(K(9eLA65)3[4:58S>?,T6Rc7#-)T#,MJCND17[fWfASc1^&5V
<#Dg_YT[PW[2Y)T&0HBB\R\ad):2+IRTY;F,0O0C>;-UD2NLgOZ>GIPTZ:HRdSFE
0SfH52)>9N2-D4PL29;.?H3g#+/U?-:[HHYQPbdSaSeH^8LGb.MV4U@c,\??e>g[
SMTES,VbNAAbg[L=[DXNV7I3@Jf\3<EV@,H;G<LdJF,-+\g@^-;ZgELRg,XPS<85
DI@@.O#UX/GDKB6SRZ,=K5]Og\CD2J/AK6N1\F[+PDcc58\),R&&G>R]O<&gISb,
33c7\e4#>-@CZNYU130Y<O<68_bD.Ba8XUfE9/5QR+[[2g9?(D2+PV?AF@c<]+(@
79-V9Y(?\,.A+S@?G9CB&MZ9J#O.V+f2L&9G23B^>.DDW=-[NOR_RKUT4CNL5=-c
[f9#K+OV4ZGTX]]gFL3OSQ2<8D4;EgYca?@g&=D)7R/9O9L7]Y+BCT_<aeH9^K;/
T5Y-fS-c7\\dYPP6V:a=NWT<>]P_/EaSS<SB9XL-]](2R+;E,f5/N.^4daOREU&c
3.OK,9<KQCX6D7NPL?=?.6YX>8Z[bd)Y[(YR,bU(4B-;]@?S@dQ_J3<,P7S<1KW#
LR8gT1)9ZJG/WL+VYGP#2\fBYDb.B-ATEVJW\]K7PDPc@]9OgKZ92Te.0NFA1-V#
Z1bV6[PH==b-=T@-dY7\@Qa+aM8E5B7.;^@F?UA_b\7HF0A0DFU31?&HORU?Y6\(
WRf-3_<AP^fRbYb?\E8V^-X4[=?)#3)IKdcTF6SM1F3CP.TL4X/g>4Y^:c^(,;3,
[-NIFU36\eb@9cP0R\<aPR+P,/CM_Z3#c/G,^?[TTKeO^7gGHg)<fb@gR9BM-GE&
.?&<Ec:1DW0B?)ZeIegbJ7&K?B;+62f_K6-3>1=(_ZK^:??)7#gCVECK>V6ZQ5ba
AF)0L7f?^@=AfbW/dKe;PD=.Xe#).8dIG<(>.:OK3>\O0R.;3bBE=cg8J?8[?g:1
4L+.V5aY<3G<&;Dc(#f&4?OASLL7)-\<b1U)A&@SP^S<bQB2G/c0BBU3#.TeJ\D,
UX,DXYD7f=MV]U],,Y17_1dSXee[L>W>[9(I9(0_H>U>GSEP37^U]+?4-eQCIF?(
C<4=M+g(FZY8-OUGBG4O>IFW^b4,,;c#I9]JVV][ad8+Y9[V.=Wd4I+E()(N[FcB
#.Wd9d-3PfBQFG#VR7B22K&1_a4aX8<cLA5,,BHA,R8H334:1L;1@QGL/f9Z+?W)
]);\R5/A0EPgR(^Y-eVX?T&:E572SgdLYH<K8TgfW<dJ?:;Z=VIEH7;W7LO-4_QG
K^21C[58@L)GXSV_LX=J1.VFPEUMB)6H8H#-):ZP:,+K4)(VL/[JLL>]13UbT_gB
&AZ2O;d0aH;D.I9(.HgK;<<\Z&Zce/+9NN/X[KFP=B?Lc8/YJ__KLVD]@fgXUL5L
3-TT#O3P02TAIY6[0,S38=I.E0b_+QQJ)[cR(Hd[]OW?dQ1_[FXT/MV1S2K1(4dL
,aH?VgTS/.^)[^I,TILDPZD+F8TbR/ULX5ZJ3Sa8/fR@W9;@?U[):DD/U;Oa9N_^
=GQ?;4;2BN2.gFKafNW48BAF9IFY(ggF=UK,I7fg?WZfe:VR2=#6L],<7/0>I:Gb
1)@5dF_G1]G2XQL.I>DSSR2SGHQ2KYZYHI,?5G>6VN/bPCXK,>FbBZ=XQAa=^SEH
GC0:5S;?QfSb_Zf;BSa?-ZR1L:@1JRDRR_XTOc#QW]OLM&N>0e.GK0#+(4Je,EQ<
R-DfIJ_DOJ[AD.T3b06^AZ_fFI3@.),&cFB9f:\0HLSKLVf]G?0(+aLGeM&WL1?N
:<Q>d1FXY@SK&3L(3(gBL;5@dUH4[Z[D486ECQ=U4^OL[>eT6cg[K(\&MJe7A&X]
1YUa)^;0:B97X##O]V@/(A^99.4E=LC(Y:SXE-RFUe_B\&cg)3GcgH#VP@_6C6Vc
IG7cT;b8cMTPV2825PEUG787?I+WA)MI_WC=Fc6Od1JI\gD/HdBO7\gV61<P2&)8
=Qe),d<TLF4&c,3GBSE)?(?@f1,=:5NJ^Q.S/#.FXB22ZYL;I?1a>K/6bR^#@\BI
DM0(?1?30fd=@2.:Cf&MC8,G&\Be/^>cJ[8SSW#(ZGEL_ZY3+P7Y?M5<D=HJYOT/
PT:7C(X78)_d19M;McD6W1LBY@4/(^@O?J3F9G(bg@MM^eUL1L;P@cD;D^?S]>1/
X[,CD=U+_Y]YAa-EA(N+&SW,BN9\K8?/>?/9S;2dMeAg:A\bI31B(YR3]>X?F(0>
)5C/e7:Q2J_H39#ZgIO,F4L6NAI?:c7+76Ab=_/QERXI#<b],7NC=bdSX_]LL^FX
(e9e1U+JC:3+D0fS<<9-500^c>\3)^K&1SIRS^Wc&OQ=A:#,YUG52#RZRDT#6M^R
Ae/d/.5Tc+e\>A<=>+^_gCGB8a<B?4=ZD53\+LIAD&N7;+3/L]J,A<8N4g:9=JL=
E[D(U&QV&WW)cg=Q8//VWG?S--\UZ0M+AOY36?3A^C\AV#VP.)W37ZX5F_eYM82,
,0^KEeQQ/NH9F:MHMTX8I8[:DRH+WG6@^+cM;g7RE=Xc:?UBHMGG\=g-T1AKTH^H
P6PaNOU&Wd0M=>OFE^LK1fM\,+Ce]fBUdJ2_gQ6GHG^ONE2KYW>@3@XS5ae)SN9N
G\.<)(QS;f8H60:-=>O+VE.g08<>NZUY39@27JGJ\:#[ACc9Q?.QIb2a6>P85Y#J
6K^YN357BU9_dQ-L7CRScROgOA?1QI.\=XNM=-BD/gAEbS09Y2Ha(#/56<&90fFD
\LJ:R\@ea^MV&Gb#4S\2>-&)_.B5=M,>>ZBc/QBCLINA,_Q4;#]dC&DFO4d]R/L_
5Cb8-ORV&/84[XX@U9R[#VT>^GOT=W_HBGQ2XO0:G&B+W]fEW7_f9[.&+ga@_EZZ
^-9I^L&EWdSDG>0M#YV?WWQ400b?g&7Q3/GB34E-QM0/IQF6RP:e<:1LL[:1_DSJ
IF0VEP\.VgJDKAXa;5J9^JOfSb9)8>WcYb2LAWMb1Z;cd/IC0P79NcZ=?A]I(c4:
>Z5EW0_BaG>-^V&U\<98S9]7QRTd@-CEa[a/gR,8KU_54c@f-EFY0fBfJYbPR9.#
9FTQ_0SbS&d5g3:SZc_Y8T5e6EgXX-6J]&c63BUU3,I[-@eJZHE^6FVNPS[gJM[K
0B/2V)QTb#c#AP<3<BQG+aDS6L/>](L3VJDN15HfZ.SH+43HAGXE@W3.VY#=EfWT
G@8(@FIG<2_DN^HPYcO8E]30Hd8E&]G9.bNdU=+.7:e(HU>B[?H(-@3e6](TPV0U
V^bL/ED5D(XXCg6=PQg_S/D9BddW<.&L;2)E-NaeAd#<L:8R-FA)<.R[IXA4(&KS
5W&Sg6Xa6/6<SI3X/Af1Y687#g7Zf=BEJY/b+cD9_XJ51B\TSJK1bB)gX4KGA-#Z
SCJQ8N2GcV:0.,SIBH+1c+S1FP-^PVQ=WODS];6Q^N:\UTK+)GUCPbM_cFc7?#6-
#,6eJI3C0RV140]dP=WJ8QF=-A5(Z/2I-^N(@V_1QQDNZ\.c:LB]K/TS/eOXgR57
6UfWg58C-bTIKc3\4O+5H6THcZN<cE,-bKdO>00B=12BVA.<dbOLO;9:+6?2S\.^
CK2fbSEX356<N>:6=\_D,TQd43YS)^?f726TXQSPA_4K<K+QPWPDX,K81O)C\4_P
_baJY?4#543([a:,86__S\fGU7O_N_JWB04GNP;8,3g;]NJ65-\ePH>6EURA#&-G
<X+bfB.AKagD.3_Se0d-/M(Y2]GSQ(g33UP]HY/0[SH3,U=O6,FfF3YXCC))[CHY
3Ad:ZL_E]DA6a._AAe6#:8U-ERc@9H@SZE^D:.1G:D7F0[S^:ZQOfUfg8cg&VVS@
657SM7=IJSJTED;/>:ASNMFQ6DQ.c;]?EUFT;QC=DJA&=fP?CY&+Z5C&:^0_W@7;
_QXSGR^Ob4-RQ&@[c?<S>^0_1@&9bBHPZOMd&e3;J[5>KJO_E5)5dT7fMIT??A4/
)\[\OD^(&gDgZ>E7J?(1^2JYD2Q#4(+Q_+2;]6=8(;@AY23^Y8&)W+geMgfccU&3
J>XH5a=18/CO1R^:fA7_OJ#9?fV-Q&7W(QSHR\3G<2#QJdO3_>8=?XL0FMbIJGT^
)fM:S#Edg7XX>IgGPfJ3LH,#ZUTHO5#/4:J6#3\A/V[I;Z&#b[W16M.>7<5de6Y+
+D4^0J8,cRNG&A6gaL./2d&J(2Z5B)=VQ)2GIC2F&IPXb95>P@[aN-]2e=R&,_C+
]#OF4J@6?DYVb3G61I^Ya7<WMXIg&@A?Dge/bA>;T8TRcaW0OaC2E1SHgDA:/DC#
Sg[]HD#O;A^H5(gX;+(SgWc=I_9QF0V6F<VA80>V_9I7_[F-#?P8&3UST_#4X51(
3-9H\B29(dY9I2:P&a=KIW7R>3OIIf^D@76V_V#;]?X(#]b=deQ=ZY8V:9N(D.L6
V@=;c;Vac)0dZ65QBLf\CQXbeT@D;WCOQ&&M4(?IQFASL@;D@g@+TcC[>+932d,:
L<F\fLO^6)F/YdOTE2H[-FZ(Y=:EOgU=Uf8,HXLK4_[\5^E)V>2X/NG&V2TQcE+M
0/QZDUeY@bWOeA]6VSdBK>C,1g7a.Fb5^G90Y\)e>NN:^@d^BdZfOLKd]J>.+XJ.
OV-=>G;=XY]B8S(bJfVeRCR\?Z/fF^MP(NEg7Q#T0fPd(]@B&N3P(N^Q/@1<IW&E
3^#-OV9),?_C__0)4C8:9D[\f)b245\U??[4DU/#V@KC?Qf/VB,AJ]TNDFH=YVZ-
f#?gPe\&@-6Z3B11>R@Y37Z-N=7+OT_KF])WA#g_+;(>#XE.=QQL0.S))ATQK3H0
7+e6E;_N@&)#>O5\7&J]RY@JSFHMbY<TC+++eT6GHX<WL?KLaVRX@fd58/T(Rb&B
9e7G;f)6UF/<W)90[_?ZXF0[5Z&a;@(G)KK3]/R\:T#eR/d+_BTQ4(daf>SMLK@A
XA)=(OF41AZQAUaKWJB^VGM]UXR28FYR=NVPT0?DI(ea#OJ3]TE?C;?1XaM)ZYT9
]FE]c^bRdI/:6QQ(\;B+AIObQZZ0[&\LMB6\_;/U=<8e5H]gIZ6>_Uf<5P/H.Id^
1XB[4VaXC^JYH,2/b[f\I\bc:L,Qc(]XLg;\/]YB^27AUaM32.&RTHD)C4:PYRE5
^NdSYO_(7f9\I+0O=U(\D4:2-21?TOV?(.[K)\;3F0\f\INSI;MWV]S=M.N)WW0E
?<7CdO;dND:6[6LRT5=VA[)[D6TSI=<,+;44e/YeQD_DR\[<?P#I=)eNA56B;,>c
GB2a(d^AP<(Q[NITBKb306DRJa9.CPeV^A4L>XS;cPcd,c?II^>0W#JMVa/M;WC4
IbU8(,=EgL)#U/]8BQWN(L?1(Dc+BaaFc)P-:?SZ4cT,,_7L(FP/_&T67,I./J&T
WA6:0^9Y.@gC:#WdYC-C0d,P32C1KbO0@e\-L?beM10d.1DCR2.>11B.&K-[4;L2
PP-0.BIQ-U7088HXYK\1;0K/Y:aRCOK5HLYQ\Edc&X.4cgB)-ETSDN.Q6#d7G.;/
LgC(OdVO,R?TeA9=86EUMNKPPCLVe//&PNf8JPee_.8gdQE2<]VDL2-5(K[d>P.d
&[4MEU3KX<?9_>@@A.4)ZL\>L;4;:Q&070.^ZG@2QM7F:b_I&a1YUN:B\],=GLMf
G.?4C?+O&.@fG&M3-E1Z=:F3FXU8@-0?ZH?[CZ=N]NO^6NUd7eY;9_ORL()6U/c1
(dgf6=>b1?ORD4,b5@9#H#0D^ZSVHUC88Y(S:#3>+?Cd5H)^W;5QE2+:W[Ce/HbN
f&IP[NNgBT)>b;;C-<7GOJW:8BPTeW#NI^.HA/XV0GfeQDVKSQ&g(GU@Y?49P0D7
FKWWFV8-H8/A-9>-LZ:caG&^FY=-Hg/86A&V[4>-3>TbCY9Z.XAC^EAX@7Y[>?T_
BW&H0+NDXU<FbURH=]C]eH#08D\c?g<aZ3bMZZ7<A(8.0DISVOW&7:U&g&<S@#b)
]T#49#dCL,^GHe+M<L8FK#NA&]5R5>OLKa8-?Yc>:0f)Db[-BGH&O+B]aU[0ROBZ
IR\TI^[D0HD1M0gXdcD^BN@2U7OSLT,;XO#9(5C3bee_5;eE@cN/ZFE_:NcOT&ML
P9W7>?:P3eJAB(\SCe\8DMUf+cFBNSEZW/8Y<R=8P<+,5\+;U;4X&^+X73RJ^GWB
J2A/6&c;EO?7Ea)S)U5bQ42bN9^]W4P=:?)6b?_5Z=^_78W&VH/=<c2d+ICDDd)O
CL44(g-:JLCN=GOVL=KN+^g5J2F](1M.W-INP5KL(.#d[7P93;,4b_g(RaS(CM4g
AE=NdIX,FF=Dec2JXTM<?(F&GME9807PHA&eQ,A<R,2\BQUU]YQ+6SFXca3eS8-G
XAe0]1V>B4PNQSEOY<5)8dUaGRR#\NeOebVW._KaX9cNIU_=1HbX\0Y.;2IQCKQE
D2;VT];FM\@f-1KfWFOT^-[]2(H,:&g>F1Z=a-J@S>ef?bC<2<+JIVd<G[.\8P,J
B6BF=Gc>?I]^,[X;;]K](e\\Q[\S?X>)<]G+LK?O)X6G@bdANbd=V@[SSS@(3]5#
;a743e+7)g9NH2@3^;5)_LP@ZUA<Ndg6:d.S;P=W>?;[Q]bDTVg\\Z#g2a#^DSfW
e6.#?JZG>7,;P/XL\]I+4H=<:;J)Ta9E,QR-LB</0UJRS3_[(Ue4(;g@#dD71GZ1
[d09]<M#>=8_9[7/b\fGc;<L8=7Gdg3+Md_I2O8/Y)BDUfg(.@&H.(I_[[2c/bPc
39Y,cRQdY82H]9]P2#/CU\N]00EJdY.D::a>9<U0dRdTNF]JYIe_&/EG^3CP)V>7
_\Nb5.?02c7\XLd+(,)fE^IT^[JeTV-L+_36G>/fPL3<aG)3ENBO,.JQdB>N./E_
](QG]g\7-KIc5WWY3.J.ScFa1^g>_W/f)Qe^PTb525POe(>_U[7.d0L9E\QLE,SX
YO85]N;(?XR3e?Z3\4U\b_,Z+<)+Id(C@E-FK6@GK&Re[+b<eMOb+E-FR2M?Q<?G
eEP@II[>[H<U>A;\Xe#_;g)UWS3=[P_5D2G^AKF-FJR,V0e>WF0<6[cLL,&&LXJO
6P39<Fg1=-#.]@1,RKPKZ4W3)46ce5g[c<=A>=7UGMc+SgO4dYd-0bN\,<OPC-_/
6@)W]UL+Vd4_>XOT:S,b/e[0O]c4<^f+e)cdZH^7/F>7c09cRFT&7>I:)3#0A\2G
AVegIYG56d+B[WYbPYa@78)^>Y@GZLA76#8]>XBO<fMX:(MO6]OL7RWef8.7>-c\
>])aZ1/>RY7gCLVSc+<[d9cN/T;7@-DTJQ=4/GK)UL+5aTQ6Ne-E.N(DWHJ(+KU_
d3Xc6[3^_9[UgYg?#_0U<)0,V82dgRVH#[WGb)19-eYS\X;I8GPHb2#PAa668XLZ
<:_4&5(dSB(La68W;TP.E=V(e([:W2JRFX]cNDN>_AQX1GKeG&fc1<AbOfD]^;WO
ZDR2DW7-,R5=,B6W28+G81&;0&>f()HCB/0)C+++TbL(&.NDbQLOC+#N4<+JD(^M
A]>Y_5BT;#A]LZ8OBG]Jc(7\J,H>gM5V:>[Z9I\E#e6U8J[U8BI06Za0?R>Ne(MY
Pf0c1XJR5A#aSM?X4B2&RX\O,.f56)UZH(E)f<&QBXTDO2de8B.;bO3600H>ZI92
,=Zc(O4R/8^3Y)UCacb1F:]VQTU>MY:cL_A[@K^TQaKO\2/.L4U]R3<O-g#WQ4MJ
91_CJ@H6B.=IAPgP;DcS\g-1AQ]:0+M0-X^K.V0e)DSU\]ag5XHJa3^KUG8\XKR5
E.F9BZ&.H57,UCd;14<PB=>?,E[-HIa^6(/V3XGN+)<d8,+W:GdYA@I]fM/F:&TQ
)Q(b6>123W[4.CfESWX561PB7-<X33IK-2X=[Edb&(LP6O].bOKbb>.=d.\#.\&F
2UA5+RH7COUX47bH;AOK#.J)eJH&PgDAMX@YHPT.Vb<0dKNV1;K:U^<CU0#d=2OD
R?\Y9O>0+>F]^)Hf</OXP<I-F=V41ZBUW7F:#:CFG^.BRMTB][?VS(;aS>7L:^O:
=4c@]45WgB@6f,BZCaZfAeV2#[?[#.U5KR)VHDG#XM9_Q(ba/R_JKN[/\90SKR;=
(27gKN1F&LAPUQHP]P7XYW7c[T@1:]9dWH0ZDN=[A7/H2+/I_J7/FL4]U887SSOc
J9]:4dRD.M:LQH-JSQ,?XUAa8(R6IXWFWdc;?TS@Gga8>\3#bNLdNP-GY+LcLWNH
8S6\FG\&K5S1XZYZY_Od\Dc1^[0-\gBHdI:fN]N?,NXC==P-BT:FN73F?6-M/6#X
0L)E#L4&45_fCe^g0O<@e;@?,5)K^T^X0eBHO?CM,Zb;G:I@c:Z/H6,Z@JaK=UDT
?&^Da&]2C>dQ+D\19E>75QGa4T+EH>0YZc9^6N^cJ?G83+-FWFMf&a>6W#83\fb=
^=^NKX-[7#9+66M>-\e)8@DZc(9V9.:@_SQWMKXbE35/3;e?A\V+7A6Z-B+++fV0
_=K5]LBd1[cG=LK^N0&+X&M_KSC4MR^15549a=_V>#F<g.e5Eg,\IMMG>.O.LdUD
_?B,KD@XK@U0HR79[fVT1AR+cJ[01]((@8=6DaC9S0:/#AK]JU_2SU3>9P:bY()U
N#Mc9-4>d[:Hf?Cg(XbPK0G7+(:<UJ;\O4&aa-NUE/U<b;)[0[7T7+?(J?\X;QTa
YW_:L8I)M64=4,/:[Q\T8Nc.SWBb..EaCQ)IK<RU@V;C85&9Q2C3MF?>6D<R.8KD
#L9eGMP+7MOf6FS\4M?Z8[eS#:3,3Z>1#)7RBX2,a-Wa63;SSH;QSe=TL#bbSY@D
c\NZURa0=&.O@CBP-3.ES>QNPY]HN3B#Q&7<8Id]a,Q9b[C28ef4d,?1BD\)_T0T
U8ENZ/b/2^/++JX54a5La5X.a1+He<B-C39RI[A\ag.HdgW4>G^V,XE^2;&ga)J4
V#g87=F=ON2NRb=1PP=cK3d6CX(\DfbR>\D8f5>AX\[<R6S.Y73>M39;5[=b1[I.
[a/C<Y?8QQbR]<CN2)d_9P7g1::1aR;8Za?AJ>>V#g7W\UECg:Z#cf5DZ29IW6^0
J7)/G(Z/c9R,@AUg26_5Hddb+dH@S5efT),-^U,d;0(=Qg_U]NaAM9RC=^?LN)T#
(AI(b9G9,gFZ&MGN^-]I^&KR>WE5A7HCb=Z=-JCVe=?H7;+CYVa1#0Ta3@6HDGPL
;DXH(Kb9AE\RG0.#&WV_6PGOKb9f?9&L15-8a9TF(V62ccG#)=ffW42c(^\:I3NN
6/=9(//;M8P225YS5=M(-C+PMS<3VHD<1,F^LNPX)SXGZ?(7K6,)LBHP30[_JOdD
S85;[RST_J\Gc&OC7+72<2@44NGHA?I,+b@7G[d^@@Se)d<ACM;B,&Sa\#-5UHb:
8E-VI@B5BJa([;XaK:1V(_/ZY_4,43b6?B^C]DUY1e&+Y=E=?X?AcR>7/[a\1[#Q
L^a#@L6:9=1.FI&FG^/Z/I+gB+P?RB3:dX+dU&P?QQJL>[KPFHF@-:a:KFV+9WU<
D1<,=Q>?@gc3&c[G56]GFI,0,aE(K:6E&5CFE[1(&U<-.KSRT\4.+</L-6<g-;7>
WRC/LY6dG4C6>&<dcE2YM47-OZ2X)10fS1V+O0^X+O(dVBHCe-?[4<?WDW1,G,?;
SS@^RX\[57#XYEe=KE+J:PM.I@d4JOIJO3fe7dASeHQ/EV)QIdB8/aS&N_+eTf&=
(H?QE4M1@XK<[I8@c.:&a\^46IL0.R5.XF,;B&&-CS4,:4P&P&B/@#b-2cAD\#d:
CcWRU0J0HTM&ZS2M4YMV064--YV2U-2N]<6\-96-g&_?;XRf\1BA>b@dU\<SL5W=
Vdf\73UZR_V8XMc,]aYBO]I4AJPdUDQW8:#]d[5g\;&G=7Z@&3b^TNV2Q\IAYQ#R
N[RMV&SKFWR:Mf-gLHEX9Q_Q&,NO:X;&fD:+1_H9>.4-EM^^TfI7+3+S?UbCV&_8
UG2S4D1M6U?2ITE:Rc5,CWG6/a].-(8ZX-@SB;7XDC^.@0[.N0>2Y]QK^e88ZUEB
c<T_NF7&7-T4@9B=I9O.Y:KRfg@DS6J2R<?KPW5E4X.0g(:VeTR\;EMLQKZ9\;S5
AX[=Ydd>Z8:XG8_;-B6<fdOg+991J\ABeHgUM=ONFA[&e8cBT[D[.&DI/ReDU4+)
O3WN7ZT4OXS;ZHYX9U7(d]J-\RTZ<-V-DILP\8661f#KVP2]DXK2O:W\5IDNU2ZH
A1BM&N;H7e/O+/fU5g2<\<4M^IQdX(\CR0?IV[c8JQ+HKg>SVXfaD9g+fdBFG#FK
KeUFSN2?[U.=Y61XJ5;7DD;0B&a&eb960d]8MfN7e@GT66_OaNO5eb#NZOS/B0,J
cEJVG,T+[?T@?UGD<?G>PYV1._QOba,58(B3BE2_N+=JKWHWR)L(L,[f:]4CR.(&
eSbW0g4f;+D>CH<c3;H1>3M(44A59Y,^O,=,4YcJ]WZ:,ccFL,?R#EP&];_Jef3(
ce8]6YgW7LZ&68VA&NHX(D09.@IUeEbFF6(-46&A>;?(eM1W<K7Z@/P/,>46^TW/
(:S;Z371=U:KQ+V&I/5)a<1eH?#^Q)&UOVgdU6Y;2>&;dC/O,_[\9\JPB\X2+8#I
W@/&DRab3Z#R:bD1bcGV9?+f.SA./e>>2Qg&+,b3HJ2VO2>](\d\2g:OZ71=(:Tc
W1QM@YD#+SgKMaT3F7Y6I6<He[8g[BgIL<<-aZV/T=T+,E_=a]b+UaQc:(G2(PP)
@)d4([\HL+\g(8_DgR=55D/gRe\2-)[R=[;#9?,,\8&?N.5([F]=a?@(.RB<NJT2
D)0#-dN:RMeX6a+K<PHaB[Z_6RACQ934-PO<?,V\eCFfSa8OIS8&2FGV&S=/A,L=
>MM^[?-D=3QOeTM19g3A#A]f6N6A;)H_(D&E\Aa=0AN_\aM_W4bdVKWUG;g-K:IB
&<-/KLZR8ULc:Z+8ON3+f.A&F&@YT6(E\@:eP?5Jd715VGTA)Te4;IBC[THEDCZg
D(\c_^^Q^@UNZ&U,aDD3AO1/c(9d3^&R#&b990K((0P3ND=IY[YU,U_KF?)T?&UZ
bZH<+SP<CH\a=^T?U](Ad@(_=-FO?5CHVBH7b@V#VVEJ/UG;Oe9#AFV@V;+:FP_E
,)@=SG.J]:_B;)F4Yd]>eH?ARaF;fKT-7CR#7UM/F^?Q8b.G5#V17cOJ.>L+++;-
DZbMSSTO:KGQ=a1J0#Yf41JOfd>1FA6(I#aeYQDQa8,=FFFELTZdeGB=b#AI9@fb
?P?;A&+]H_M4bQZ5Z<e6JW,29.([ZBNVaf_[;P.[Vc:=</DdA+0(NW&9NKNK./:e
8B>1f=H(dT+EVHB7BC>egJ-)PNa/B/9DcDSWH^YB_O6AfG/bXLb#]fO>AGG>Z5))
A@^O^\3#^SF47DGO3bAa[#C-a^<6-L_;1+8g<1g@bGc7;@&D0-87J_6@,OVEJOQ]
Y>f##B/5G&UM^>5af[dLQRBf1I_cIab2&M/P7+ZD^5S3a>5<947c7K,K)a/]cXfJ
1EZUg721F,-[>;f,P@V#>4+276]VR118[M0O6A^:UNRV[XI;EO[[XePA/KSTM:IB
2W/\P&\W^E[8&3>]/5;EW<8a,@cZU4AI1&,L(,f#0a_N?5:(O<-e;5;+E(G6-gQ@
U9GJ-297,AIHP_2FM;G0KBMD.EAbOPRE1\6BbA]L,f[LVM;YJ.a[[:Y\<M(cF9Fe
1E7CAED_1EY(E^Fa3YO<GeXKbEJZ&LOdST2Q;=ZYgQfc0eDc()3@b.>DNc\Je,2+
H[b[07SZXccJA6F>L&0^OP0<0).b8JBH]?31N]X10-01OXR6&S)FP,F8D48NWKT0
JEGA+WKHA53aZd,5CYK[C/T4;P2_@RS)@)>EM5ebIG+eE5Y[e>EB^MFR9bJB?bT<
0(1T4?dY/?IUP(dP\B>M>^^T;93V5)OAC&_>;UFFg7E4QX#a[/eF&M2Z4&#?+b>:
,2e_N3.S,49_K_P.T7TMD1^bf65Z7Cc>=C>5K]CL(^EFI27YH_J2//ca(g/I30b_
0LC:);R4C^+#M7J#c8ZUCb:4+W[IK(S5B.+H(0?J?dPRYda&RD9Bbe;gVV..08^Z
&N^8N[?P,0f/A\-ODVNc&@,11(_?UE\&+5,-YMH73;aU=CS^I?.Y+8Z(dfXKA<&+
C]g(@FS11JECR3P#cANZ0S8FG/DDC/:X#N54WbV[[Ne>IVa;N93.W.FKZ4;.?:cb
@g#FX18-21bB5HH:#4P[a<-f_c74Z&C^09cLVNMaDX226gSUHV3_L6;GQ5,X&0.T
SB+S9M#<P9P>(a1\O/ZaL4b@W.:T,F?M#->Q#WDM&KcBN6@QPK#@IKeU7R<UXW9d
EH:CcQ449CUH&>=2&Hf-b^>a77NG;<O^4_P\(S;=PJS&eEN4VDNCKOcT6SRg5FfW
)AL<]0f/.+>7ZZQ&,>&X\a-MR&/556[O87<9fCIC1VS]\ePV/GU2[;NY-4F6U<=;
LW7RbV#(>YVK?@[D,N?]8Y@fbe[&5&beG?TDD:>K1>[QB]SHP,T(0JYQ\c0833f3
64aO6;,de>0KM-,DK2E.bD24,+f8/6cgd81+T[J>\NF[Hec=:O)R@MVG\3dRg<Ea
0GM&KY)6&g+2X)-#J_<c+5CF0;F)<Ic]3.H[QWUYV1>&3+)]]+L@+HeX[<Q,W,9=
BNHF&bW:+O7RU#bTYZW/#UZS@CQD\d5R.?g@<-ZQ88__6f86,JbHaeK?D?C83WaS
7F8aXQ_[##[Nf7?TOeRaSIIW_CLI/CFN[,,4H0AM).C4I>-:ERD=Y/U?A&S]QX;X
^S<;V04cNTD^BR7A\@M6(R3;S:-]1<\ccAHcD;Xa.^f+Q+W#4JE>QM@\,C+eO_-E
8/2g;->f#:a4,N^LffW^)2P/O+-TR/#&P^FbT(W=W;O-+XSKM&>6,\W64XZWKY<D
OBQ6CK>b]cU,_#V.,gXD#\)8d8T>=Je12C?&caRe=+R60#VK&W;(G1,J8#R]@V^e
[T1&Zd[D<7P@)10U.^Y?F^KTOUf)==\XGD[,SI)]D.UL_OBg7^Q#,.XbN9>d5JOY
P9)64[.=4;Y;f.@1<B[VE5HIe<OI?6f86)(#fg-M6QGa,Oc43Nd@R7O8YaHO<&V,
JM[=Uf24:1YJa<ceeBcG44SY3V5-O#RRSZ[5VLFNO/>>SZ+B-M:\KWI8@OOaWSbE
Nd#37)Vf#>@aT#E\Qfb#X\,A^)28.;Rgd0AHVRW7KTeIG,DF=<#)W6B=SF=dN615
R79MFO/3JM4bC7aWadC_^HXLRC/<T@FA#J@Oc>fE(\AX#=^e++Qa=\/;g;OMT/&-
a\9:e5M_>0/BM?Q=&eed>48<M],HJ4@/^X6J1D[0GQ@#8a)VM]L&\9?WQKENO&Md
W1c3:Ib+R[J65gQ+S_521+:WcfPcD<a:Xb,2897I+OH_5,9R(7@DSe9R7#;_#6eW
DK0:2aE-fBPRB+&/cHSSc;NL07d224:gc+TMHQ6NDJ-g;bXD>.98-.<[;(],Ke--
-YN/@cZ8f)O<[g?T/EgcBIBf(EH.+0?TGHGaGaa+E=\.D=Z+W]YEU<-b+RYT:-78
EB3eaSHcA#ZI]:VSW-FfUAVMIg,V/O?<:QZX3W1>;bae;3G6EgYgUUMXJ\E[1_#3
,RRMd(;Eg1#bN6@E0UZ5]Z6?MK8cP(?dSVZ:c,,ICEfH=EOIW+PHU0XW_6XYAb[4
+5cN5ECG?J6/BM]IPY=R#b@=/NSeZ[9J=V?B2@c+@bL8M_LB@AQdB5=8Z<UD9d^J
(NA]eANW7VR6,gRGC3?ASg^?G+AS]&^6D^afdUUB&^Y6[9D2@F23.;f?f\ffTR4.
;RH\92UYT6L@_3g>YTB+DFW;R/;D6Ie6f@6gWOUJ\=5Hf#4LYVCcR)G+e^aE5LSd
+-]/#O]F+aFD06U8bU+bV0JfV<?Q9BcDRF<Z3fKN4IRY,g&C)WSIg:/M&/\#?5gD
QN\;>fJ7BDS31(+H<0BcRC2,G8,0:U2aR>e>;ZZZ)_.?U4YM^KS1eSF?aO:R(#e.
dM+aVY+0-&VQP=&2U&;;SSF];X:gRJ@QN,O=9#+U)YKdX<VWf8(AN6C)CO,,S.-=
H:f9[]^H8Q:O0\&TBH)H.U;<7fQ9^TVK\)(-(4LF6K@b9:E209_9eLT&V:#9bH?1
EIX2@+gEWW)B]F##;b8cNd2RDg_\OT/T@_V>,c=T:Ug.2ZfQD^KJ0I-<cDS+d,MO
DW45@DfJF/+T0J]:F7#KA8NO]B;Q2(eI7VS_b/cD>(WIU:aF<RYH(:/,I9HK]76?
]W0VC8U?<.(PgOXQ@GQ@,/=H#.&\TS);J\S:5eWDaG:a#YV_JSF98JDfa\,=U3@E
dRZ5UQ<eQ^g8H6FbYG&PSZ;EX@)E6(^-@7U&dePY:,:_29@,OF>CU?ZFeL]Xa)],
7>W3#]c#WO_c]S:;aeL1LT_B&F:eacCa)_8V)cB/>1>bNH)ORWTD73_11(>WIP@E
57M2dBWY@(Z\0^cR:f[;\D<X7)g,-?cN=&d@>S]e8eJg?ITXL5B#Hdc&FT#.K+8+
PGC0B&@AJ5b\J[5cZGDMT45;?FK;gRW9\U4J0.eFaK0bXZ#==9)[/43ceM]TPWJA
F@GFJ<GPHaMaRF7#>O.dL2A4\,;b,d&#gPQf?_#R4gC>S1f>F-8PTO(f9O,R).5a
+H,VSRDT[a2=G_.g?\C@a22I<Bg3V0<]E^dd_0#\\Q/3-,ZLHI_7\,gX4>S1#](D
-;TMb7HWAgYM</eK;2@9Pf#R\D,&cF,BZdZHXSCI3ITaF#GdXg2D.00H6&E,+Q)L
e^M,/YPXMU)[T+EGKX[+?+e[U-6(ca::<]/Q&+V1cJQ?\9<;]W?bA1REF#.KHO(F
\fW;9V8Q51bLd+[]/\_I#,758:EFL(81VQ;;IFRL3E0a8FLJH]#H@-eFN<\&D:3T
EfT?gIS1<A35KC^R;Y#57[5.44Pcg44=X9>>4TKZ=7];7I7@U]L0ERS:,#]JS?E@
g+.Q-P=).SHM[Z0;>/-aOTC\IJ&NN9SE@f2OE;78R_f;GR84SdSKCPOR??+MAUW]
86BLS+OPdgYSNda0ROVbWg_;[?+4b,[<C1@FYdX.4W(#4WAeDY(T6[+eI=fffd7a
gMN0)3S;F>(LQ2=<_PHJI;E),T:ZG,^OAFeg@G2)W09I#5bVCPZUU4@7Q-Q)>R1V
9YY3FN?U2T4Q?2IM][FOOXL4SXK[Ne2g2WY<K<@2TEZf#=HF8Y7K@4@A4DHA+d(P
U:IY2U,d92&,.4.b\V,KC]bE>QXN6AfA4APNUd3ZWG;L48G4V5J_b38<9:>IG44d
/Qg>eS7?&0_2:T2cgJDW[)9(RR</2-2]N<MY_61b_[FF/&PO7@2?HYDVL?.\?H/Q
Bc#HX8g;J^(ENb<Q[Hf]9T4X9_6VKGHCfffH0X(X114)9cGc#3E67>618;_)+KaG
RLKMaLQ;9:Odb,A9COA5T4PIKSf:>>0aS-&g+#,?:d[?gd8/LI&>__Y<W9b:T]1J
C9D=C>1f#G-Cf6eb5MS26FaLHcT.fF^GN&>.8>D.=G&F-_&1TMZM^7J=Z?P^63bU
9IdE0f,@.-;[-SJ0E=854FBM4H[STDC@^;7gZAT9#\VJ4]c07UJNEa?9DaEZ(,BG
(:6N2:REaZ,Y:_L&b.CWcJN^JI1#,<<:T)<U:Y[,]C<4)aJ?UAX]/V^QXI>,(8]I
45@g#CeJ:VU3L8,A\6bD4MVFaL3@3V\HJf;Yc_QYAHWO3\8,__Z8;Y,P40,6J96c
36DRd/4SeNY14V^5>^M7>IU8GdHRK[eHY<FGb6LTO;RT+-;1Q-FZ9IgE@NNO#<Gg
OK29B1N?1@WZ4\<Q:We@->]bDf6MM^9SE;-].5;-;#,NV/J\ZdOTL<+26cZ;E_;.
-e4GL,\O1:R+]B3O:6f;3/14U<,74@&_\1Nc181V,CR6I4T7LWbPYa^aK1#]C62e
G[,JRXLTe&O-dE)AcZUc#42+VO.+F/J5()FabFP>?cX/2;BXN]E^>;FdK)Cb+LK(
.VNdB653NB>+ZI+12d9SHeHcaX:&5LHc#9K:UPV]e<PO<R4HbI1\@D.#HKXIZ2,[
FKC,^f@VYOWECLN87YRP1De:=@-afIRa51e2fV&5<(g:<4QAfU4=(;b\TGHD56Cb
7--;5K5aBBB6UDJ/_0+>Ue/-&CNE&#WYL/3#(GXSCPFCG_#aC;9BbNJ,aK>R]H&J
@_A\fPaV6#I49]7W9_E3fBF)OA,58D51NRG=Ua1?W[f;H?RENQUMZ_&g7.G^222\
K4ZQNEN6W0cLg8P;P@3+SHE[d8H/K\4/ZLD?Ac.+TH]/]>)]PeJ[gXH&[Y#\M@/b
NQPX,,bcbX2PO6Gc9IV)+b)P&W?C(X0==9(CII[CcZ[2AE?+\ITI;-@2VL0M=2Y(
0(0I\#<7Z1D[a8cH:?\H3Y<MC-Qc+JPJV70^0L4DO=4b6LYW]L&SDB2#O?);f)FN
>QSU.P8E\7Ma]H8:+A=/)=#R3,M\I3Y(,SB\+,Z^Y6GP1a#3CRQG130<3<5bDE>Q
Xb\).?[K611e3>/F4^Tc-7/G@\?D0)B&)SLc]1#SC,TR.eX]VG.=I=-_?KECOG#4U$
`endprotected
                
`protected
cdJ:CM60FK@>B]U:OQ96@3KVB#;1\Gg6W5R2COf+K89\.R#3+UF]7)OGHF8Y_SC;
^T.+S6):1L6NG;@AcT4J-SD8>5X=.RdN]#F(D&XJM<N8[8?P=:-b0Q<7Fg/6R97G
]ObAgFO+N1A+AG)M]J/^G-(=Y&IP153e:.F1)M)G1)#()P:^7)JfLL.H8]de+#DJ
E\E;<695dNLP7a)Vb8H?-RD6K5Dde.J?RQ0,QgF?D?(M8S7@EBMRa8:39]EAIP[2
O4Q2Jb-b)dD>@M5X.=(#<+RQE>ASbdc,dSa=,2.M_E(,^S@+fB;[_^3LTY9VRY#0
TYdI=F4<6dJVOc34JOQJM6G4]cD:FZbZ>8]MC/0)bPIdB/?,&BCI+Yc_-3(4gaSO
@b?2<IdLKfg6X-051SSR2&MCc)8e;SWOEWP?^=PbWFdWP?:_]O0YZaQMCV-e;L8^
EX(&T0<5/gc#2IN4d(Y7ZA;7Tc#3)[KgN-T/1@\FAH1,=FZP1CPB\K?P6\SZFe]T
R1GfXQd,5K8d9\K>dB>4<C2]@VC(FF-A=$
`endprotected

//vcs_lic_vip_protect
  `protected
\XEK:be>+#U7XaN60d^:N-(L:g_>OY+dL9I5?)4NL<Q;A>b1O&U)3(V5,bR+E3V+
U+@4BfPbBV(6SMQY\GP=\EbGCKZcKJW_Sb\/UL+[=225Z>V>M(_WfL1cD>&G[??N
IO\,F^N>DELIOLdR:Z#S?dJCY:PeWe0,N-7O(W6O>]9BU4OcYXZG[\R/f\@HDJfI
A=/a#dWH+A3]>Z83D)U@=5=0?Y?PaQQ2-f)?Z76=3OKcgH/:d((]a3KA0bb57R.S
\RF&V<Je\>E,9G<^,XG_GCAI2((PUM^),,M@VP-/)(:PB?dP:3Sf/S_FB,K[W:TY
Be?.>)e5.?X^M6R;I2\YYG,72NaLdJA0;;1,\K7/BBAa>2;JdD@&LYdgS.FeS;E;
g;Dg;b]?>]T]TU9#&40^K?6)-ZgJ_QC.\Te6C:^1J;@&e<=.Y7QDVe+[d&-/Lb>&
1L,QJ01dJ+Yd[9TT)8[6.N-OR(P6gR)cL[>d_D;aW+B-ZdAV[&L)ABO=UEME/?M4
/:96G6,a:7;)]ZI\S.D_8,:1U0^X>:?-NSB1aRL^gH@_8AQ)bB1)8Vf:23HI-P5E
;R8YD_X:E+7.:E:Y&;-\0F8e@JW==0f3f&J>&dQ>>72=V5O6_e^F,C9TZ.(EJEMR
R_21I:ZbfQ(bKg,JAc&(GNB]K3PU6:AU>2_176;J&]GO@G.)W2WHK_RHO<T9<C.P
BV+(b4Gf5]aD<0T9[A^4SO)1=@M2@/6:HSK:ggAG+9.f>NMJ9bXZ9S]:];@.GE2I
J8a&-1KYF7__8eR]R>JBBJR52d:J[)<L9?.D:VgV])ME^<NfE7W@?)2(O;DaZH.)
g9C0\LYOVJY-[LcP5&2\J1,FdReMN^Q>X5&KVDY[@1CP^ed8JZ+-PR0XJdD0KT1Z
#Z;bcBNA2ga(KE,7cgJ<?V7La^UfgGa6O:R9;QKLKBf+aAI6+a&-O[3DTQa5G]U#
HI1NPa<BIJ5_eXaEgaQHO,gdV=)3&T3JEOWe12:X944\W8b_#TUW/<QH8J?K?2>H
N[f;93d_@LBZ000;]XbUDPS4\_C(@7&@<.eH.#IY17UcVAF(0EHCZN=<LM8S\P#^
R-3^D3;YO-e9LQX8FFNKQ&_P03d43[DS:6G]R1ObWD?V\eXHgVaaS?M]M1SQPE8[
S.M,W0]DA1S_OPY+S_F+R5\GcR&A+eVc(TTRg8HQRFVW(W@(OQI.6BWPCdHfT)P#
^9]0IFR+;J<:_B0:;#0(62dC@^#/:/.?G>5./_ZAHCI&-M9S1#P-R[D7=(43]XGR
2S:6g)R<[NUVPHP?[?FadAVI16<4J+Sa9;CBA<g)f<E8@.VU1fJ+\@TJ1_b=<ZD[
Z,Tb@192HOP\1<J#a;?RITgB.O-CW=5(DTN)&ZW(&2X.\@QC0F-TJ=G3,Lg;4N6e
1H=L7WJ7@@UUZ_aT3O&_/L__L9Qe^T/Q@4#>31RD1R4646+.2),POMV<2)WTK9\8
N1M92begX^IN(SYTD5d]E:,@eP_C@MP.,JE5O=fc.@<^Jb>&^SDQDR97Q2dFeBE<
B&@5Zb-:>&Z;W?S@JOg/a\&RA-dM9]YDeGACJ>a^fET9..)H2HOU=?5#<>7IgTPc
89NNKc.a/608E0R]Q62;gS(S<&[+LBWQPQF7;FSKJ#68^RJMV<P#/J9bE[X(;\Cf
RCaMD/<CZ.eLb5AJ[6dI(&>-^2Z25e:H2F2HdNQbK-//MJT,S)F+TgE]bOBZ9KM>
ZAWaa:AaI<X^PBG7bbG&f&8I[.9EUO_BI<HQFOSOFaF2EI3f14N7T<S9<2g9dV(K
4-5CSafcf<fGGQb?Y/2,e<AHa\^B&c\<54Pg0<CfU,4R4_2FOBc,37AL\YB@b;0&
@eG@-K5dFRgGVH(\[OKKZ(Ce6X<Kb.:A>d#=]EO6_F=e+647WA,cSBYKUWNCF,/S
6+,=DXGR7^b=&.X?Q;6>>BG/ff=.=&cC.(>=aXLa(-?,cZGW^@V\MLJ37UF6GdgO
#9MF9SSSECMA9.@IR+7=DFe15P-.OCPc^OHMZff1G;8>Xef-JEM3>?DH6@Q,TdNS
eL=g@EI?@??^>S84]YBB0CL.QJ[4KJ/6Y#=:Q@@?)A>aeOY\=0\E4_N-bdLSJ5e7
fgCc3/DPEJ3)HK9Lc+cL#XO(G>dfOb_Ga3+UO.TC;MAXGHI+YDT1ZJG5LK/K\1?,
;Q7Z:I+Q&Y8(VecO_RRHZ:DdZZ7B-4IaM>9>R#C_(7ZJ..HLC:JbZM3SI,>E?fgW
8V])G]-O_HbeBD_#C@ED+Z.+K@8PX>3cg.UR(5&R5/8\^V05d;O4,.CFA)3X=O0:
QY9BI6.Y3-^,77&@&e<_68QY96_+TDCU>(<eK<[(TfH@VA?1N<?2^4J+Q#.ZW;LM
dSFHUDI,gQNQ+_T8L#:aN)UB=]63N]=P)&eUMg?BHI3#Kc#-@^/BQCW#b;P+0#F)
9T5[c9g/3:]GK_,<6gGD^W2PdVb^>FM?X5RCZY5AOER+@/Y8(1]<dWaZ]?TcE,bY
8.NJaU;5/f#.&^<O[cQg6CL/]bH-VcReXSGMdCe#T8>_/-<V\2K17B3=1b&_cJO9
M^_Y8fZ:X_=-66LCKW&a^=EP<H7[[NXZ7PY#\]c>;\OB4O93[)XR:4VDN=AC=D>[
RQOXgHLKTAObI?.V\\DOD+.\Z?IZg1IKET75c(^3^P7YN4/.5V-UTTIKa+\[MYNB
=+:[bNPf>[@S@[[93((d+/8IN-Yc2>X2FX9If:K1VYKgY\NM-DE&8+O8fV0<^L;;
8,6LP.^5E&PIRHdgNB_LNYTB[EK&bc&f]/B(Bd#:L&M<=2D:Lf4e1Q-)V?E]d1,c
b=X4^^HKdDeNONLOgTYA#X2TM/89N;9<7@_Qc2A9dPPHFJ1gM^6].L9Ig-+a=A-7
]KZ?LcGCZ/V_>K\_(WEMH/-GLP\c,/S<;IERO<BIN?I-@VT2BcHA2P\Y-B@+@[U4
J01c4B?UPQA@YB6OEV5\D2,/87+gGPV0A=,Y^SO^(R>P<:.)<:YH@G,K>Wf?[@@N
IM7SB+,BU20@c&4b&^MDOc8/BdBV:)ZP#3MNO9>VQd&SCWU9HF(O@<DCUHN#,J6>
RW[Yd]/NRWJOLTK1a^-44]@@N.8JeC075,]dd\X2]AF+X:P5efV_8>BM1YQ9>,,@
L^[#1eS?::_23K&WXa:Z;:gEF_US0SDL>RE2g;N=]6.Q?De849P@3O,Egf,0#WN^
JYLZ3#9PP3)LA8^F>ZRHY93@YE47Rd+NYR=:f..+;/+]]U0H<.ea_6gG?&/2A0:Y
gB7aIaN#8aVRC]bOR)[cT)?JKD>2F)ECB^Y5g.DPD-U40P5DS8+OX,370\/KB45I
TO6D12e&:U[^#3G2#4_X+G?I\T45C1@U@=-6TM#7PgR8FI(P:GW>R.g(_5U,:X2Q
O&=R-g+9NL#cZT>@a>Y7@&DJ&JC98;JfDd_/@IaceZgIDT/I^MZ&2RJC7-RC9404
QR(Z-65gTJfQffVGQZIGDTG#_PXRI5,Z3JB3RF3)G8G2Rff<8QVUgDMQ=W:).R\W
OPOT\HdSR7^5_0[W(VQM_45:a<S&?\A44\5@_8cQ=3XSP^-X5dL\-T@5=@&Q2@PH
:dbT93_EFL)V7LXN.SLS8JWSgD2geg<=HB-QPVIc3<DXgZ[2[Z<=HG5&c=;&1#Y,
_V2H#ORM_DKagK#\e#(#?@3b^<.^S9F#B[D=/ODAFG#WOA/).^WNPgF8Ld7MD?[V
(5W&@XY,37?d:H^S.00.=:QaRPSFF0>K8OLdWa-2R>>474Tf<Nc/?:O6&BRVN=\D
1&Y7QZC+[eDW9^a<bVRK#f#Da+_]\>1_0IJeO-&W&d3_)O/b2ZZgZ;KE-)0,WG]#
GZ_;SfgP;XYILH(CUg]R0Y#2JE#b6Z>3=UCD+Dd=ZECT0F&)SV4SC<]cRa8V-d.Q
Z_)gQ?FP2M0a#c_c?6RBLO,JXICU_GBWD:L+Y77b5JNC-QMF@M?NgD-ET(7UL?0g
,HfN20>=KW)R+PU2O[(#VN,;Ubg4EQ[,/ZUOI#=T8aCLL6)JKa>F<#[#NUB7U+a)
VLEUe]R^3_OVZ5QN>B/-Y8;<Z0CN=EK33XPOT+<G9,&XM7ZaF\E=6-]Q05T,deQ>
CCBQgSPced3Nag6I)9FH:,Ba:J;c>eeLWf0<VE5:)a=4QU)Q0<EEUdJ+KEf#A4d\
KHZNa&FQ?MRAW50?:e5]9>+C4D1@K+c;J2GZJf97/J@CCcBR\\]RG>NQb=52A\>\
8X183>=dO17?eAMZKB2^f=3_]ad=20Sa_QBTRF:fX,._XCc5RDY[(A,.SZ:SEX.,
eTd3[&f?C/FfA>8L+(0@[?FSE&YJBAc)e7[?LM=@^H:g(X9YT6:)\O)=T+EfN>RE
ZL46Z:=WI5;&\fE3Q:bS.NSd:1+gHOK_Td5])KV1R]?.[V8HTeIgCGeC0PB12R:F
&H0II<.S>gWc0]aQ7PU/I=&YC[>U)[6YQ4<Q+4b(S4<Y-SOOBEOT^?DBJU]<NYI)
6Rg?ReWIOTb0.//R#ELOI#0LX:bZ6gf)SM/O19?W:-;3-(@6&?#SCIN<P7.<NHSA
^+ceRB:+e>[>[1<K@]U9?KN/(Q:H.[RQNFQ>5fgd9S7=[U(]8^RJ6.,@,Gf6f2K/
-4P>SB.8:aT_PTNZ+-#c6#1\fT#EGV\5gVa7\-TQG.46d+#?&&Y=dcb@[RY@YXCd
7+E(,JMb<VdNXB[8;&D;7.bB[UbUI:=:8TA(,RLMeYeI>0>M;gG)_>e0[OQ;>SM&
==Hd3g)PDcVA+SQ#@73:U3>4gDNAIg;RA2@J5SaCXP0Tf4N&)Z2X=]F]gQGY[5[#
KZPd13RO-6M_)WS]V^OHAJ4V].,W_1.NaX@3HNR34C7IZeSZ^Gc8?Z/Y[7?bMcKK
SX>P[:2,=>(Jd:ac2>5A>\ecQV=OE4DQ>4HXK75X84UHaEXAG@O/L(9WUMWHG4NU
K+Y:/MAZNCT56SZ82[3fU9K_AYMG0O]L4g:LUJYBb2D?OBCRf+5+W8RW1W(a#O4a
P>INc?bX<,6bV0G0f-A>M5&dG]3H3GF_,R-Q)@;D-bKc?[Y(6T(OXN#6H[CJdZU]
:A+,.U<E1OUP]g?SBTJaO9QKJ#E9N9-V(afa5P-Y-1H@YHGNHc@+-\0<9=WcZSBO
-G;.1#PVeM.].+KXKO3S.eO.2CA_1,V8V()60(aaP)=KVDL)(R<86c<6/Vc73+g?
BCag(?/XU8+eaB7Af2eJ[gXRXWUT?gH<=0245EX;7OD5XFIN+?D-[1/SD)7YL:@B
/?L=_BR-Gd5;KAb2d?32:&^(MD]CZ[8]cUZ)64H^G5^;@6OSL(.;?J9;O?=MXd/&
dG<94:fL>c],L6=&:ce(VUc4]BKEAJV#1YfdH3EK)@CQSLVZ-Q4+gVe4A9\5(51;
#BQKSWN&=)ab]\:Y7WQ]1FQHMceZR+gYb/eBf(3aP;W]SKe.)>f\Y6U#L)(AN.6a
IQ32D:-S6V1NNZ4IOZ;K(B]EZ#IaH2O&(=73=Fea>93EcT,)PSR-FA=Q4Y3\B1Y;
(]dY,602Y?AQeYXAH09?YKKC/E>4)VfTM^d3;U@+Z3-5-3Q<bN7E<Z\@-G6/6<[?
&BF_?g0Q]>LfPdE(D]/@WX53&Ua&UG#Vf1]TcRg]65M<_TV>H:HRB-b50WgGP=,2
Id5OZ3)]Q??/R]gcD>(fXL:B][e7LaA?W4aZ>)V?S,H^O4\VBIG=fZK-KM=1C:a(
+X?,62F=>.g2#R.O.U88=dc.44UGHG^F[D5.e4QdR2V2Ad2)-/E<^=aNObEeRa[E
)8].,?07a#&]d-[3G<HafR,e=&D+Le7?G+d[,N(;X[Q:Z2(2147#cDVe>5(B/Y1^
B9B]E6P]NWH?G:F\9@@>AHROQ3_;IA,X-Cb)K)U(ZR-=J_:Q8Z#PW>B66W7G<;f_
Y\C3QM;CS&1]S07f?Ga^;?eVV:>R8@(D1>\[MS+)>RC:IT2&30C?CZ1?UAEbe+__
@\QQN+_BAL3F\Se7.8D.H]7/2/&)Ke6aR96d:AKWJ)E1,H^=27,Fc0L??2,OF<HF
)=JQ9Gf>SWE]1D0X>UN#L+7EO@SOZ^,f_=UE8O>@;T:c@1)^ce14e,42FLOa1?)P
#@Tf;/#ZYN(8eHRS\5UCEb&6PS](AM&P+>0DH+1fFaW=R8VK2f\=F+-\V.Yc5ebQ
f@)Ga==YXTa_-9)FNQC128>A_\<8@@;OMS5-2+.XV)D)3aA)U.6<TaAAeWU9&T(S
9AXS4S:b&g)dP\88:;;\)L]cSJ9/6&]X./bC2:Jd6gLCH;AR:N-:U4:b;ZXZRWdM
H@GRDMT8@:87dNg6R4-Q?[J,[C=R<^=?GY:_@.E&;I^:L8c___1AMKPR3<gU/;EA
)_V?=_#_+f;cD.3V&[BB73^CP<\d^)>CMa#Z-0^?#1;JUdQ.D]WQ8@2Og6Pde<TY
_,]IcKZg/fMZ)F[C_1Q\J)D]E]?+0J#28BUJT@<^;dU-&X[.0(,<JMO^4T?GU1W=
IHU==(.8Z>6_aNQa:43<]SSG.DM/S>Qd-Y\OVeJ>J-MZ]c8/cM5g.6KW/cJD-@SH
gP=&W&N_W@eIbFL)CPC+UE)RL:b@6(f@PR2KX[;N:[^7CBJ.&#)d#a]S+4(+3>;:
Xa)/#-B#^<^B<H8TU]HNC+eAMX..DGT,#dW[G\&9gP=eMgLSMHU+I;UUg]@9&T-U
?JHX&E+=42FSa_#KMVa4Ug8/91OZ6UBOdcLA4J8W3-[U18bJ-^1/M&Q_N)(-\7@9
4,8:KN43Jc9F1N#8@d6b:2K+SPC1gSI.[LR0Ld3<UY;@#>R(Cg6ga-C#Dd]-WYL-
48>Na:?cK+bVKFHS7W24NBP7&<BXU:,R7eJCT,(eV?b7(f76B?PFeAACU]gJL.X&
NP/AdXD]\#)Q_gbc5Q@35/FD;)bM#fBb#+E86>2bg(\K.MC#PI[XDVT6K[cYBG]f
ac?S8L(W?(,#=0Y:6-.PPAf+A2JNW9[d9<:KAJ>#OB#0U1VICKU2R.SSe>dAOW<A
L27ZJ]Q<Sd#KYCB(O^#2(aX&P21f<]8BY:]-W)J+:,RFI9dgQKE>QML8-LaB]EDG
TEEW5D(]Jg,bO?/#G&SV,CY#^[(7ca@F;HDK.HG62,TcV[YNPM_KEJW<NA?I^f4Y
BV9?^@+_GecU5DT]PHBZ5T_b@D.SYLVZ6:.ME2>:efP[;V1,BO#Q<4[6LYgTGSJ7
G.RSPKa3[[Q12JJ8?I:K:KaeAHK\QGOEKE.:fN?/Y)VSFDg366Hbg61H^3WZOAP=
W,)[;dX^CE_VeaJ[Zc?T,^TB[:=bA<64#5\\>6UXMH-c[77@&E=+&@bOc[Q=eY]K
geII.J=JNG7((N3_4_IZ0,MgX#5SD#8?e1;38Q:7SNSS5Cd=W^7Q&+&ff:?#[9/@
SbH=P+_6,&BAcXe;<WV55c3=][BbK\:7/OXbJ/[LTAc6_N=U2M@EUT6M/IS:O.G6
(5Z24c\LF6XM/\ERYO>ZH9._fd))L?M,b?O&\W:AM(IT1+RcIbJVUJI6RHDR99;b
aN)&L]Eg.9f]@TaI63\[_B;,=]dL+X+&Y484R00-,5I?>L+.IMRCJN71c_<4SA>e
-0RXd\KSb3_[E]NOWgD=]Ac65R<K>e,DHWf0,/dFefY8FcI>RR0<KMV/b6+ac;#^
]gAKdE-4bAgdJf]H&;ADR0#W>C;(R\4]&>\Sf.1@Bbb#1-=b3>,==J\=MBG9\F:U
>U6<QQI]ZB5<S442H0dT&c.=MgLBXeaOWbE_)WD2GN@@9,X(ReL-P<S,b@,gD.-&
Q+@M/13KSF&MMaVO#,We=QV_F@7;Yf.(We-N=0=JG+(,-(K]VI+)6[0eX1>U3(YC
gE7?,BB;J9X8#PGEfJ&OAg?KJ@K6H0J=N.a7J2Y>@e=\_L??GTDg6D0<RLL(]DF&
KbE.JeEe0ZI58?D2V(fG\NQ>CJAVZ2[;040RMDY4=6.,b^9O(B<&&gbV5^5e87;Y
=>@,VH>#C>DTHG)5NR[<cMd0?/\::H8b6/GH6Z\^J@TR>S&f2dIEaM/8GgN3fFP,
He0,&fVVU5:RYNWb/TM5BINA]WbKVYe9cJ,3WQ=3W9#e-D0ZE]US4&-Y<^K\QNG>
;^QfMAHJ/?,\QbeW/N&Gd+;J9VEJ<#M8cQT9Pd)C;8P:.P=\>NUJ/bY4G&>&6c>1
?-<\#NATW0VeS)G<&[26-VaRe/G;0+1.GN;S<Jc@1B0(ANg8=NE5S&V>_>><;P17
<V&aF)2#0)YPO_HbV6S2=-WCfeNA6B-^[Oc09Wg.aXdK?0?TM3_)Z)X0(5.BK?#1
E7-@>8BMAKFWWH@QF-1._Z^>C4c_U]&G1SQcZ7&9G&ff43\6I0#f[=P)TS\A(JS)
ECgCX&Jd2+:\_:5(>e>LC.+_I1[Z^\+GJ9TT>dO8<fI>J.aG_bO4TKNMPTM2g)H@
J+1^g;We-DR#?1A7\Zb#d.E8:CXg9F7D(QUf?R>KW9O0G1MXO;4FSKVS2<[9&\XE
DNdZ(I15UE&AHO]4g\2/^T=/c;X/&[,0O-+2]..=0FRHECfEY1;R^O;\UT,JOL-6
A)E^57IE15^6KW]3>9:^AJaL@F0B@SdaC2DY+KQB9LD-gW#+bd1WeHHR6D1abU_T
IcYb/&-:7D9Q0H&/OBZT8@,NFb0Rf-+0\S,T.P1g\;01PEXM<-R7dUZfKS4Cb/S2
GL^X)dE?W632^&>,b[<#/)2,g(bd7e9S]JAaV,KTcNKW5E-ZPT7O2L=]H\N?_&KH
e)57c[<<VN@AA_GLXD=9b>9&dEG=aV4GFb5P<:V[8-=QZ2:ACW_[\:JD8HCJK>1O
RVE\PFSL\<TUJf?GX(L5@,MF2I>5LZ,ZW^A)0gL_C#12@+P/4S/#D&Ce=SB(NKcL
17ENH3]g=<[Q/;Q=&eIF7WbMK_KgZGMLGbF2[&-T:43KX2;EZX26=+772(@8L7+b
Y<VIL&70[I-OW035-ZA5N>f:>c)XBQYN\-c+dHB(BEQ<C<--3CNUI1]:bC;6E7V>
Q\\-()^gTcSP4)ZR?2SUS&?D,b9C=O6&fH.OOUM6[KgK)]]f3WGM25_b0EK,&]eN
T2R>YB\)5IcF@P#UZGT^&KQ,5bUQRE^&WE)3\4E;CKO<_W/4M(9/+M]E,:X:LJ+\
(8LaXJXc&08FcdT(I4J>9f@B<D-]\M@)Ea3GaQG=JS:.7+T?7>PO0=VGD&11Q@V<
>K0D<O,gXUeU3>7SSKZ(+fC)bfM-gee_F9#UYMO.7dH+T(b.B#PGagRYFMQ1T]7^
g=>L-@fPO@\&=+=DW])[5>C+/3NUGI<MG_.3YNb#G(N8M[:N9[4S<I8)_Q0.&R4L
e4-]^JD&TM?.gRJ?M&YK&R@Z[)gcDU([5#X/-CWS1B].IBSAf5^c4b_FJ=4@.c[3
\\/<_b,g(6\TL/G=dO7;(g_<gCE34_a5FH=#4JHKER5YP3_Da6@bgK]IXcEe)-Rf
<-[CB>TeOJ;0<fS<g2Z2eg(c7Z=.+X\gX3e8F]@FU58F2+,5&(.C1\4.KW;<ESNK
-F_6@)URZaA(6=V54FaA;B.5@H8UG]BT=0:#-K8P4JPBbZ=c\4G?cQBGfZH;fbdB
]f3_fK@.,>N27G3H+D6L+&>^TTXADM>?2#P51KWMON;SX-5.@)\938JL#@+c@dN=
#WWS#63da1A9dI32[g[)R=c8>dSVX>P.bN+6EM[[K.]+=gcR,W-91]Oc+9=GSQ8C
+Red#XVd,EODg1D_#TG(@\?.GX2I&e^H-45_\CgVM1G=X<SK4:(9W1dKDD/OXb@D
.@3D@?&\YA46IX:/bUGEYVReY#>2(>=Vde-4>c@ANL\.H@#XSOd[Ne4(GRX43:3Q
P.XOQVA0IcUb,7C>a8GaW1LDBFX),<(6Te(C@<+;0&36c32R5/a?gM/NZbfB&&LZ
.LTN+bF6fO0QZefA_-C#NQGfMEF8,@&>(9&)#CDfb7\J=]XN1\YeTEJ?eUbGP;,^
1>NC.X7:R1M0387S1,d=MO8XZSYV>;e@g@OFT#TVMOVDFH)J,M(@g5..&TfC6YIO
V7=<;PK&c<0+aPFXPRKPYg=1#H&e]L0ag.E)<c34J>Ue;ZQRHP;P9\^=G7SHKBJK
+_BZW[d+P]CaE6(5ZT+a@cTgYWP,fDJNQT2;CC&&/E.G\@5O+OJT&>WVPN\=P923
ZCFd?DT^G;GC8#4)P3ZPA)BYVUW&QQfQaSI5WH/WbLRTQ?DQ@8ac?)fO0V3WR;?F
>c(TT;MYCC)<)4?TP+VAV/DG/F+9?:3Jb4e+5^feM:9Y@c]KL:?:?eHA.>aKY#1-
5N1S&EO<@1CPT-]JOL&U1IFR7.9HWP+0KW^ffeb@AM_.2M(=.B?P7A_M:ffe5-:#
C[F>dU(@0.2636F]?b99(b6@;4?TUTdL:N7R:>6.]<2,Rbd>.;Ta&\^_BfAGeUG?
G:?ad:eMB:>-.X7e+6O(SW(eO>D0LYL3=V6JcC0XbB#f05Q8->^ZE,SUJG=G1@b[
748?baL:&IA]b^LJ#_P0=)RbEa>KFfDS[&BOZI5F&1.:-59aLbY=Lb3#?Me73QLd
/6V5)+Bb8T?P3b]cWJg<g.72>FcMZI,/<a(MRZT9UD]99/QgRL./OO0@5+16O7]^
>Od@+B26f=-W;^QeAEdXR-gH&+2Re1S.]7^2e#[M7B,:66<HXA\]D683H:H?CGee
@5GZ);VbgNQ6(M3,Y..Wac3CeM@VD.V8g-W&]N:D#0AM6?gH6[<MJ3ON6gW)UKSI
4aG(NB+>M>(]6;(VC4==P7+Ud/6bRTEP)J#FP,SP01;,KBP,dQG:f&<BXXaU<(@O
D2@g#,/GR2/#?;I][RE=cUY2af;Q_X<eQ27gYQSNKZ=0&^\KLY+2fYI<W\cEE2&9
MC,TVOTU+.C9SAU2b;4Y9<9R4S=fCOHeG_+_9_-a&_#[AD?.VTCW=9SC74CDEbSJ
U\[0\B=.]eJ.,8aSDY[+LN-7YB.>7Ef:L3-/NM[J,J.,95XbfP/<>e9[^aW3Z(CI
O?]A\E4LXEaFOZ89E2\4&bBHeC,^D_;bN0R7EB>;Sb4#gMGUZ,b8__TJbP)F;@R6
6Q/8]^TGc,L\44#eO_aTS<&-02()OEHFb:Y);D5X,/MHX7MWV9+H7bM(?]/#T<0f
+]9[Cb0H0>C0RM3#KN(2W?>d8L=.SeFJ6V?8@2SH^R&XE<NU7UXDHC\FUZegGLQQ
T?1RR02W4HIRQ9RLeLd2-cDgU@68a+_8G+(<JN0KcK/<]>8?LY5R,4(NZbLN]Z0c
6M=I#PdWE;A9c-=8-#M)0>_a_8\R=C6J/7&Z.cTJZ^335#MBe<OUDL8US\eV2:91
LPPHLF#aRREA4;8KedPOBg3CFCMd[8UB\_7;(_0VWa.UbJB0:fV[edQXC]9[DN;W
eM?#Z,XRNcHN@[B?:@.VHRZ@BdP7O9NcVOPKN6_e[>KH\C8K0COWGI-K:27@3PLB
>,-.Gdb>#0A+NB&ZRB0X4V.Vf0ESH587ecb[29g]ZD<A8N62)@@A>&T&,C3(0fe/
.LB^dC,?F1W&CZA1TNG]Pe:e#6YJ_0?1Za?YYd/b,J)EI)C\H>He+-3Y=M1cFC@F
cIP_H2M-NRDCJ[M,?-2):GS-.S<I=W2X)efc2H8B823=Pf#2-6c>a+(+@>1KYRC=
aXf+417KVD5XR@85+L6b8I,d)N#KAJ)JF0SC^P?1<<Z\LG^H&3>g[UQIa]A^Ngg6
,3B[,aY\X<dHYVZV25NQR3&E&;<@e,BWCPAQD604(I<\G$
`endprotected
    
   
`protected
9H3&Y51T44(EM5VPYZ+45Tc:,>B/0f/]N3)FP545=81-@,+f0cd;&)3Z.0e\B<PW
R&0,/HcZ+T;@GgfI^Q71UXc:3$
`endprotected

//vcs_lic_vip_protect
  `protected
A[=0dSGBK?+8;f;CW2I=)+R<3AU9]C6DO6=Ab)Q)[WCVS#+9ES3.-(A84[KYO/MB
bB-PDPH7>LPANYXfUH?M2<b-70CZ4R4EbGf(W/+#LM9cO(7^Fa[@24eS6+2;6g&G
E3>4=PIOZ9[R6T.7UT,EZ<#,&U+&@&cRXMeA(Q\UGKE@\]Z+<Wf@faSKS4N.G.KN
-Id,UPOR3F,2UdaSCW2C3IF@0D),fAeX<Pc3e\QF[Y\ePK63TK(DAH\OeS?JH;<T
[^N2?LE:,U&c2f-EWc-,HC4(9>33]H=R.@6VQa]E=ON[f3D5[5^\ZVW98(5J>IRO
_#G+cJR;>)eAFf/_2L(S3C1@,G7g8BbCROccgG10^SFW4VY:=_3KE]a?(4N3a=]^
#4=9+3CLV1)-30<Z5cc2[I43?ZO,c3+UP(VKR(b7?P,4Ja\=9\:8JXXW>5<0A?5Q
d<<_STQ7FG;J;_0Ca?UG\>?bge3;L#SRU=VgUZe.5[_//<:4ZH\<1X&dBJO)BTT1
19-T0=&LX8L[]L;Y<@06&B>]EC][-47eFF14dP?CL>6V]fGHHg0-+[Cf101YBPIN
^P81B#7PfQQeAB0@NH-Y>]dQ5J8^e6AR@.fHAffS4a\7;d[+QCX_OZ,TQM3(GEW@
T+]QdL@0bQ;O^ECKL3B[B<S,\23F7QO3(E-=Se>(Bac#AJNG_+ee_M9>#<6(\EZ\
/Z)g_VeDagQLD\UNT,Vc<&TI+[]fUeST)BTVQ4J?JdHK<]ENbY^fL52^GVG^fH2@
A(Z=N&[.X)RB+&WC&Da9<T3YI)HMC_CDP.Y_0NG_DKaBW>e@f<;9-9DVH@C2AN&3
8?C4Hd9gf,>/PL#I[F@SN#fTZ;^+SN=T^dEaCJ=-Q=8-IL:+V@XUP6@Z25abe&UK
57,:2S[TafVg8]62XL1OK^Y5@0G3Q6;=L2T94>/._A^RW9d=FNFQT<7YN?\Re@bg
CF&EgCT80QS\:&dQ;c^)XSP,]/AJYL=.\Q<BUVJg.ALY[3c2b7K,/<=2H>@XINa.
M-1]=,PX3QYH2+<KCb[e^3<Ta\]@XF?C=^UVV13CB:;#5d6/O?V[P..TXNWMf5)(
AU^:5CY5ca;>_)IUW.\E5QTcTDYUT.P,C678gNT8HK+A+_0AEYbF/\&+G4/SMeQ-
2e:ZSI-C9A4<D_<HT:>W?Z1,V2/WQ^cf#=S,_EF[YJUH>^R_-:>=9;.ESe1(?P)F
+W&D0MB96bT/3IdZF8JD0W.HTC11A^RY?C0X0>603;PI6;YcQ3J/T^2L1=>:J0S6
@2KKRMMP,/L5d&;bI77=3FLbC+ZU?c20F/GePE&fLRWQMZ[Y:;=)0&cFROa)>f^M
<X[KJ>LM,4=01c?4,=MCN&GT#7FT(X8]7XMc0UB/0gQdO&gePN&SPS+(SO0b9IQ\
MV=\,^U,HI3E[1Xg,7VOLA[CLbNI?73Qe3N3gLLN0X&I?CER7_W)R[1/[(W?dXNK
XPN)3<=/[IdQLCHZd83SLg4@KbdGfNMY\4/I0F[>BfB2bTLXWBe>]J#QGW<)&TOA
<SU#8=JLae>d7+6I9S8d+?F_VL+)H:QJg[QC\#1M-]3GOUK=T[/dd)=5\BXgb68[
?R66(J._=4SOE@-23JUfUB]7+.\ETOb_g?V6,4L+AFN15?Cb-T-UT<0G,(+1dO&S
<OGYSD#4Y_bTK_SeU#ea;.4b.:I+(Vb1:dc_,0#<UP-b<(&/;BK>QCgI\7N:>64U
++OTEe;2JLIKL[9G2eZO=AFGLUXJ>5Z@3aS6f<,#If0_?8[M@3M=364#^]XY9:6f
dJG5aC&CUGB2WaDCES7V\aeIb04QaX1TVO-<AJb_-T0)JcbEdJ]eN@[?c;-@>XCP
_-NM?CHHB7&A,Y1]^)V&@ZAB?4\SHa4=#d6@(X]bd&H+(=Z0^=H_;HFK&aPS[J24
,MZ@@,C>C3#FHfcP&I/^#aLREV(CAU)cK^P5:-SRgG8]?V@4-^8fNOKQO-;X24V9
<>e^@+JX1.Lc2LNTK2.Y63IRWceJdWJ4#]T8^TIR[1JFPNH\BcB2GOXHW/\Aac4g
2O[Q._ETDFgZ3_K13gHb^^RJRGBeK2B^_CJLED:GEW?Ff@E^dcS21_,H/2\=JCAJ
/523c8E7F3\<;MK\XB]8<>7G+EHXNTUa:AS@K0P/^1<dgZ&S@[AQ8C4dFD<.EPJ]
SB_P69S/\8Ee+3SdAYWS)W:eW?S-EV5E4NS73S@-fTfFRI>>2\VF9WYGdT,5AE6X
M6\c8fdNNQ\eR,^)CO/g<OKK]>YD^\cPcAeJ)0XWL8\b^XYD((^I=:JGW\9ULOH=
=7;I.;GR5@,8b5KebZ9W.(Mb?DgCJ-J?^b9[<JK)9bZNA1Xg6:S>2f)G]P+[8+TT
B3+3ZecfD+Q2O9]<QS6a6_FZe<?=B[&R]K2HS;DO<6R^V/Wg=.dU:W./9R>BWYE=
gE-g3(GRV28.BOb3>>D;#&eB=CEAYF?e=MP1aR0dN+O8<JC&#Q]VMM543G?Q-Q@L
R)Z&4@D1Nc66]E2Sa_Q\50[e7_9./O0&1&#[75>&=P\L4Q<D-B6;#\SAcGd5-@bU
.c4&<:+FZ+)A:?A)7UdNQM7Vd;YGU#1T)9Na].-.4A8HZ06\YHKO&M]Z.:Mg+[IR
K;\.)T-0EV;&WXEZABKCO-O1ARF&=F83c@@P2B@D&P<I^+_H6>H.+V1W@Y\?640V
7>.gAa((1.Y2GW+CFPRIK>aGW]@4dO:L&f<W._K>;?c3JG5R,#d-^ITZYVYP_d_V
DdP-/6=E?7a1#;V5<?Rc+V(F>#@fLV&7JJbJZSgBXC+e,N5S\<@H24PHbG21A#Mb
1-SP8KEYO^1_03/Zcb.U6TW>;O92])<6G?);CQOGIb1L22?b?D,PM8-\RS)KL])G
-NW7a\;M6:,(ca]6ILbHRHK>,c[5_D^6JZ<Qg/?VTgSf7.2X+9Nf8X+3.HQK6Z:8
9eP>M)^NdK(1-I0Y5@.f//4N&VgN+CbN7^NDD(S3Y\c?/G.)86]#=GTN9\)82=U5
PB1T^/#?J/Q7QGd4AUOCWAOH@?PQ+,gW[H=L#9H@D=4Q\HU.E&E9BeXeaT.[I++c
2,A]/cH=,R0#O;ZUYQ48GO-61HD>7_7NJfffF5bG><R]>KL:T<BXc.bH@HU<cS\J
I^e=b7d6gAUQSA6R:GRN^cP)U=TV-_HKU^F)1f:,BS6c@0V^P+CS5=)RPNVNVb]+
C]Df=:P?@PK,>9LW#bB=B]JNJc2a_/[HTK(WUPWJTJ\d_,Zbc;=K0Q^^B#20U-@K
cg]Ff3#\>YWd(UQ(JO:91P(?>Q-e-JX&4DJcO46LF4KP8?]7I[,G^;3X,02;6OD5
E2,3ZDf(Wb:?GS&N1b1V?gUB7D@f;O?;1Q/f1a#0A-=[?S->,M4+F+]5IU4X29C@
P?eTc]Y<E#O#&TbZG?F@^:4GOI54D\DbN.]N+EbQ/)G]Da3JAIQe?0UGNg?e:9G^
&9#K8@G5=/YGD;M=]>B0A,IXRA<_e4WJa1-FOHf1eO\A(HFG;HY/d&D\Mg1Rf\>Z
[)TPe#3SK9f;B15?(Q+8TMA#<f1_c&S4FCS(PZG#\,2>NM_3M5&CG,CddOB99&P^
fa2MI+0H,(d#+559LD_CP4LKH_K=@>^GgAJ4UdcV&++NS3MD&e#8W<X6S(]@#Z&4
+I/J]aRRE7G/;8e>:TL]B3aN\0J7X,7)-eQB((]:>7R[]QS9LWOTfY,:)4S-BZJK
VdOA=7I]PaQaBbWW\>]f]KSSV;FQcXSgI\U)\Ca/@YX&2>5eEd.HeCZKBWK>QZ(G
\.1S8N;?NEKS#BIS/&F=G?JAa]Q5bSRM+a39E@;(dWd6<,d60/[^RZ0_J_(VTdYL
R?B)-OO&#-;>/T+)HSA\C[f,4C>3^KS3PL_;1=bS^-RA<,-=^DJa;.X1-d3G@LR)
>OI-:<^G+UfHCSSGT8B)f7aU:f,D_SC,]UNH>eM9=^cWNG84b2U^Z5@[=J^9^-&\
@_NI?3YH:19V)]R/J7W>4aG8,QPFTFO7+VIEJE=D,D/6_GJEUT^O9RU7=U)=ea[f
Z6?_IIL;[-^3;U<6;C:f=SKO)0HB]bD06^WcBTfOIN-(_(63YMN=V6:,:6XX1HT:
(7RWRg[#.CYI?3_W@g46dWV=WaEb1?a]\W?A--KG5NV6+64NOfSeb[IJg@SP,Od=
\IJK_NUU@\FY#7_^fHZ?gK5TfCSH^aCdc)2TKZf)).L?0_77H1VR8#UMEM_8I]#W
,6YAA,4&:97TcSP3@;BQF<R-+>Q?Y&&R>8ge<,K/\SEIg4d1V47,:25A,JNa>W;;
KbMdF9#]0M#P?U,R\-NE&_MF0NAfUJ]Wa]D^V8O[DS\MaPBA+?(+XF.;(5-N,dOg
J\9@D2e?ME\EC.:Z]]8=E@&[U4gYCc_fZ/)dRQgB,eDdWF4->LP_e+FMFK^Dd8?-
8E2/Nf::]?WKR4RB[c9&VX?:af[4^8:?MWa=X-]&<ZbNSgO_)91<Ja8ca(RZNf9d
gFOPANJ_JS[e[HdQ#0f&MW7=T/@GE@_:17_&@X1G<6D@3#5c3_+3_48)6O?b-[OE
=#?<.U\8be1511LfSICY)XIIL(B?8LAG;45_F)gOP9AY-(gY+9(A9OWf]]@Y;YV#
bQ5&W)V.P\_d.NDeR)H-?JLe?7_E,>P0#DfeT?Y+9d;4FBX;aY.&eGVH7X[=KRNG
YNZaSE5[B,C0BE0Z1d=a;7B(5F:f6LU],=E_26ac1;f\F_<V?S[+1R>-J^1RLcgJ
:--[FdEVM?Z4[2#2@72FTc=(=\AKD6SOO&/4[JAcK.Vd2P(W\]B?4?^0aFc9=:c\
c8K#XJddT\X=_OG>W,3U7;)?W]L-JV=GL4WF#ET7?5QQeG&S3WM+=:8d6_:-VX35
d92g=4^Q\HDS\:2R5\WMF=_a2cEP4/)(T+G[2N8;gLJdX.#0>+ddO9D:/4YK#bUY
\AN+eN+/34/Y4JGOUeJP\UY40SK#X2bXA)9Gg4/]_7U(;#XP3P]Bg&F6-Z8K(.Y(
SJB)=0aDCOE;EZ<4&Na48C]QKFcMccZP^/JedY7VdcZQ+Y+0fPE?)8<2Bb;+.CI7
P<)68CLa9+=CBD3a;fMdPPMCd[/Aa#2g/@M-A0^])bHFI[+D5-;(APfEd1S.?2e_
deVeQ_a[#PLUVfH58eSVKY,dRNfc^WX@31g25RePK\fP[MYW^R_A1\4M3\de>Ne@
\.8;#0],e+,>13<,V;5c;RJ^:(d3Nc(5C8Gc),^D5V86S38=H/G_3=O5M&9I:],A
\5J^.1>\?;gJVD=5\C]=P)H08PL0gM.R6TV8&Ac91,:bc=Q?U_CdP452Xb;KcSHO
BeZ.MB4K[VA2VYgT6@9;_+Z(3QB&NUCe/A&TYfJ1,?J(SRXUDPQ>^&=2JRaHbdY4
I5EE)[I,D52-Z2K-F<1/dMIH^]^B5#4(HNSVMM)8&@X7?T?QdSg:4]-SAI/[3)/f
/b4B0c.J(_@PYM>R;VR]&@GEUHa0f4TE:K=FD:+]X/O^6+Mg#;UAGWDeDS>Ie7c:
?B-Uf;NS,f^g[HI+TPJBb8a05<#8A8?345W^S]MDIW1a]RS;f@;#M0&E]&,#GXPH
63Fb].WQ-4TKSTSTS2NdN2J^6aB2T.YHYE:gMG[:EcZ_V#82ZC0I(c2.RS-130F3
Z\8bO_D\9SGK^9B@<O8(76EQ#W0.gQGgR@W^fM7GU\aaZSA@#&.0-C=,aO5\4WNc
aB;9gK;,c,3bO/--2#U18O25VV8Y1DD4AWJ+<+,bcWYW8[d\J17?C_LfO526X9U8
W8QMX^-c>8(Se@0[QaVKNB5S^7.-fd6gK/[3S+VO=b==;+;9f65@OgHIc@;f<abe
Tg@d9dEB9g?3;1N90[PK)Ma4EK=0XL-O47)6<.7<7Y>_5@If5Y[0.C8-8]KQYFa3
F+gVLC5C?AUeF<Y:]7^eO6ScEC\P:a^EIQ(DY&WfJ#Yb_V,geVO=@L=G&NWT<@LJ
8P>(1/2^[H[,d]FgWHcYQC9LQB#g:7fT_8,-Pa7QS+=&.AG:+(8LGVd]EBHPY>H\
_EBKRHB32cAD7:54,83/<TF\M+,BR/;LEKEQHF):W+/.fSPJ#g&e?C(<446RM3e+
(eWA?O7QIOg9I=M_Z^YMT6OI#<F]_dA=AVI@:]94P9.e:fTLO0GIEUbZ):OTcC.6
D&35&e1[bg4SNV=gJELE-GYNS8Qg/]].5?9-R=W_Y^DQ@/=KC#8L8YW^Vd(QP[@b
U.g<2):J90&Y=I+feM#/\-I]R56:_2bYgg8L-?RJ&].#d4VLE2Z)bVF(5Q_,1gBY
,b(eY<:<R?8N.A-g#\;P](?^d/AZSMCS@G_gGc,dZ]9RQcE^:-QI&:E/;B6;S5QS
cfQB3GMgK42Y_7BXd>7_gYa.H8D6(U19X0^FG4deE[,H.WX/PMaIb4NJbQF(dN9U
(CM)=RU35>)L2NDPE.@cTX/M]g8.V:[beAG:&68KQ9#2Me15?a6<]4\;X[7TbY;V
Z9[Y8)faE\<f5c5CeQL;8^71OW;0+5DH>#(a\V0ac-#W=,A,2.+XU#=RO3fF=c10
;_2:@=DJZ]#F5XcK,Zga>28LIAT\OD#fAgO\]?3fScP-X#@AXVM:3V&+cL4&+d2;
,?b6X[J,QIOWCGUa-_KVEE[R/7C8@gVUE]g#()^bGI9DDg+\F7?JQ,,/R<@CVOZ2
&V.\NY+ZS,+6^R/&XI_e;-\_I0U@,R8B0)A-XVL^L5e,BAK\a4Lb6efJVL(-UaAf
fOG_0b?<4>/@eTD.W(&@NK;JfR03DOBc\P&]2BSN)0#F:Wb19GRIfN@JW1@9(O6B
JSF&K4b7_ITO0;8J(Z\0:)1S4I-dHa&270D2e>N-#IHUd[bU@O=W&[:AcZ[]REbX
d,L,&egC8?<-=RZ2_TUD_SXBMDZfSdC)c@60[YRW,FVX5aY&Pe;A&_K;Z#5@>]T(
,eF@9\-e+U2+9O)a?fRH&3@89-HIN]BFGQ<Za#NT:RO66J1XEZQe?OF8U5W?CE>)
^0A&?R,3SYHD)Z+cL],V8c+P7&HLJDM2_(2E.+K.b;Q-/9[\\?HgJKQSY>A-JCCC
(Sc=>+,#<F)BKRJfL67Q)MRgWI=aW]BPX<[WS=Y+A8<H2@:<6CCR]cb=I)[9Ida4
L+1dR^2gN_X4Ced&5NbeIXBI(e&(CC5L+ZJY#RM5DVTV-7)^>ZQTJg=]?c,#][OZ
VAQ+QN4Z50;OcULC+ORSUHOdE8S=;\R<,c\/V:=R<(ea)f;/W^]ZeF9<OLR8\#6)
&[76-=WLB#XZ91dGFNNU-(S.=I&?M@D=0,7?\N:b8_fP?8GGGC@=:]+aO/PUGLW<
FN;1QW6B.e.&0,TB:ce>,26.R/Ia.U2WSP,EKM\]\\>TVJa5WggfSM(Q3Ne,_f7H
f[X.&]F+2EcFLUGD=?,SGaE4)=FdeND3UR,b_L3Je;Dc>A&0>NZb]O+&?<3deR^G
:.c7b,:3Q66V@2<&#.0ECIaK<N.&Jfg\b#U(W15?WB2:4XIbOJ/.X#>IRX(QE1cL
06;SFP#bLbX&KG4SF6.3,N4G4^UW^]-(R&+?ReSM171e5T:#YFd3T;K[2(A[#/GJ
)-^+U\?FFRQQFH@>Q>44^;VLU9?9[QYT.P8KR=+LIVA2dNMWX(:X-1JO4IKW6_5^
&<A8_Kdc2C#@3ca&@]BY>;\>-(1=V7;ZSYU[ZS4P4X@\cK4<\.@(;83c>03[WUf:
^+d1gcI@@9-a+5F@Nf\1.gd5bfM_3#;<.;Z=67Baf]E._c;L)dM;.73PFXV95W=X
bHQb^M^Pe<RdCR#,3LA4Tc&1CO@fRg_5@CY?P=Y,>\gOP]F3[WOgPSUVN[>^.?O+
e#JQ))-J=.<7ZC5)>=DZKK<69HE<cDbLeU=?Pd+Q]G69VB]e^aEJ9=W8Z5(NSbDc
Q@=-g?\P&1ffI@K;IL^7bTO@6Ha=?)4]R-=?eGb.\.3>JP:NKeIJ\0BTBDU7;/,_
V8R1cWG0[&;.OdGY]4^)-&Z[6TOS28.2<-UUM]:)R7-5NaW.-I<0#4@)ObH,d\.W
&)#,CYQFE7=G)2E-g^\MP:D.,=2Fa3YLDH=eEa@KTVV7MNacJE0OUOBF/]Q84bQ\
E#O[S)S;:WKb(aGC+?L.P=QKJAIH78aB:FgJ)Pc@gbb23:A)96&eFGR+JfV7/:^^
@eNU6;)#6X5O-d3:5Z>6/L7M,Q(&&dfN?^5=MY,0/Wd)g]RdbOVCV6G]Ma\2/PaE
Uc6.#\-=Ne(WNcMCPK8INGZ6A\ZYMd(1KW=\0C&dKP=:@U4ca\?)7CK0B:0HR]20
U&\YUEBbRc^:#/:E5U6U>a6A>KBI0L>(_OBYdH<AU&.aWHDZ3E<EcdVHb4b[?P#^
>/0[X#>4Y/NfRQEJ/+^QZ9,M(\6[aH4<L-FcS>>bYO74LDZ[X_(83>0>F;)+5.g8
-/aA?e:_NTda-H>21_@V0<3GQ]N9)?e>0UdTb]gCA&5BLBJC]YGQD6McaTG7:\2a
S<gAECLAY\dX#d6L7TS)X_[F5c_^.>FXP;CSfRZG9GZU&U#Ig73S5bNL9=[g_PF4
S)-:L5;QISfJ8>)&\7e6>W3I4K\YS5\_5PL_A_9+-6UQ)3Tg-YN-OA-(F/1/b_5D
=>9,:(L;?L^fPX;a&d]Q,K(SdeJ0/5C^Id7>Q7fMORFJaS))c@;^)4^/^Hc,E<+F
D4(YPO33YVgE&LOJTGG9B+3>Ef1-M6[gT>UCEVOF2&?(C)15I9SO\_EH#^E;QITN
2]CN3(B5:ba9+/RXZX+H+9>BRe7eGTJI=EUcD+4W(_2Cf)U-<PGIER]V<g9B5;8)
BDZ]bd3):R9VJ#A,QTD^Ub^6[4K]8&AfKFNE&fD=4[M,/[?GG:&+1I3+BXLXcF13
P##NT2@eaN;E,T7eR3]ZMA_B7Fc.G08Wg>Z4JTcJ[_X(/YZJJOM.WG#GE.dOQ>V4
c+dP3N];<ZUDC2Da&;5?UB,9=#VM,ASG+HJ_Q(W(H.Y4LP1a-87ced,a7A8S]4&=
>,OJ#.OQH+d:g0BT8_,+T</BQdgW[46KF(&KK&K-9.VL^M:_KQT;B=RS<NXVJMCI
\/Q99ZNFDA+6-7@08ZaPDO+/2Ya3GaZGK4<I<d-\?J4@F(,cN&;A>)OO0d)O1Jd@
f4+T3e+f]Cd3CC9Y]f(a-MM&MOKJ=(gHDE_V4?HAWYD@3Ogec^@EH&P2CM\XOa0S
JL/\XPR6OQKe#?dJ?X-Y6f0?I=HNJ>BU_K\0D5(3D45.+3We=4TbM6UXG&/(H^Y4
H>]3VaJ+cL0>]G<3;O>A?&^Z1KU4S(5bBY)KM/Z/aa)JNIJQAb/+A=8JBSfVX=]6
Z))0fRN_ZYEDJCO+UQNR@X+f:JgLT&J4G]_0,^[Q57cVB<T6g/(+BZQ1bR;cHCF;
cAf3/SWgFN/YG.eA2:(FB:V1aDg<M:a-W[+/,ITMEQJOQEbCMR(FB.,QG>WTS=a>
#39gHZ(c=T=COeSTADGOV#W9FUT&11QOHV;0)(6f&-E]?3YOMR]gf?+J]W6<?;IC
N.fG[90MN6,=M43G6_aNNUO.P[#:Q5OYfBd2\#JO_3;1\ANR.M<N]].QZF^2V_9J
F)ffU)VR3).7?+E)0YK<eDAF/9[48(_IfOb7:S3J9A4\&f)&22;&+1B.X+@P,9P-
f4+&BR-P3UU/#7-LODGe>J56;9XY;2GGA52#XN#<9JRN\U-(^2>+8_DcY977WXQ,
TVED_eeH=@Z#cTe56?5X?ZdGDB[b^DM?]-R&f;,IFb=f6e1+R&/;5_W=f1#=UaYX
&ZUB#g3.,&\S+.dA18-5f::T7ZL_Y?TB\YR,-HAPIEF?Hd&Q,]YH55JP?W=-_;46
8cEb([E25A9Gf3L@>Gb?Y6[[[Qgb4<Bg=/74Z<g+H?#PR1Y3b(b:Y@:E,W<+7WY?
2Nf3V>0]\A<327[O#R2EQV\LMBEc#_],.0LHJII\\HIF<Z4&HTO+PMB/f.d+=d[Z
[@H29RIK,,Zc8R2:3JX50H-@e:]/+VC2V-gP=gBbdJ&g^6M>/PecXL)L)<aBc(+9
ZabP\E?1;a+^DE9B&T^NaeJ)FJcF2eLK9K8):d=T<5/bZ-f(g8X2GBVGdC(OQ9H^
0?>a\T]Y&4D&&QPBD>3L@UD64X-;ERNS@8XH#cPBe&97.K\(V(#31MVIUeBT\bOR
9AAZ^CL=,3>SY;[8Od+gBMR#<aI-#0JOZO&\@bZB/#XJaO\dE]KK+H^IHb?8[aJJ
B6M8f.U7RMZ_Bc-bFT))Qg-,?Q_,-Tag\c,9PI6H/9++8PM+BgHFMNS@8ITT^:]U
0SeA\&aN+HXQEBG4MebD=-V,_f(DcZELN]^1G9&e=89J]\-^:Y2=10Ub.2F-YLGg
,(c/e7/.^Q]TW1+fL.eJgW&^AN#T(^1R_:TOFK_;[b?Ba/1aE5@YD[eA&/__JWB>
.?OZF)NGM>U,bK2E4\RCQMC>_9@1JK_UZODIF4]]Wdb;5>NQ>?.dP+9UQF===ZI_
7^b8EHR/Mb][;e]]FVeNeC)bDCc/NA#O@#N>\&eBFO[K.-@e6E:2KYE(a7OT9Sa2
JONOE,;[)d(HGF>50LEYE@@4H^^=aG+/]Ze]YTS(6;3_0NTL0,P;[/-V=&dG&=LC
:T3^gS\a.,2c/0U&(0&J+a;Z0)[MZ6D.)&a]/a-dR8-M:9VH(cIG/ILe=3Te_ZM)
<CLSUR(aa>GOF??Z2d_,RC>=_9,=_R2_8b3+f1X6K(3,ZcZ5&FZK9cXDMb_g13aK
6#644D-bEW9aLCX#b=DEU<1&9.T[)79c&(;BX-,?H;V^aeDaX1HX4JYbZ[eHD)BU
^)dVS/MH.2WORNDP=JP)JcV-H=:6H(5U.>@]O/O2SKQO+0d@0-(GHWGD19IX:5>[
/#\X,AI_H[E=G[:3d<ELW+NgM6).)Mg=U)-9Jda09_FB^.bI@_FA.94(;^FSX(gB
LPX\c]O\=G0T1^7>a+#=SU(M2gK1UNb#0H39NKVLOFI])e4\S4;^S#:FH=^:FT2I
_L<-0a0c8=g5<=TEEc,]NSLY:\a@0A)XB#)LJ#?;7700A=-Ygc0[9L.F2SO^c>^c
cCbf&+fQ@T?fg+<--CGX>S])&U>C5R7baB4?>@Q9QaL/<+8_g_BgG[R=N\8:ce(g
R]dZ1M[0JCgQ7]AP.WB@Y(6JT69);#+?L)&553Re.f=8d=C.^>Df/7MZ>5=,efgT
W-X@8#Q3:VUSR;EJ)\e#V.;-F8-.]/G(>YQ_O^;@(Z+g-NY_f?V4R;9T>I-++L6_
AA#V830e@JeZI99eRa?a4PV-cQ3(.P^M3-HY+2]c>H)8IYRM;L_Hc\F)I&8K3SDd
ED#+.@D0f^3Z)8E-UYd5=7__8,06:>@f4DK)K->_a34I4V(V/94-G=dO@a<&1,W8
_K9UZAGYKTZa:>MAHA?LM,;-_/;7B[&gVHH#@cQ+43-,06bCd5O7<DX7OYR(H]RU
a7JB(]=KabfP2ZVZX/R0FVN/J]+ZcVL2(fM&83->Ec10KD)TMO4OB6SbFZL&O)c[
QO14[fCJV?=]X582?:KHL]X:SA;FI,<g9IN++DFgU4Q#@4K=#Y7I?#H2TUXS34c7
8#e6MQD/B+RGOA^(1R..9F/)<A/ZeU@+_^+K04-4-d?J^eeW^,76N2HW.M[UA>^U
2=0>-]()d2XGPZ=RON01><I?fCaXZQWe=]T(9[\D\Kc8?J<A]G^)5Z;a64.d)A7_
=M=]\OY@(BZFI^PZe.AC>K_b@)<P9/EA05CX>8e-UZ5VF7=c>UK3]-@M_,;=D:;D
Ac7F+JPS>f)5X.VPaa&#\TNKZWF1YP-_XSMFa3HgbTVRZ-FbYX8FbePI63gMG\gO
\-U@_QKC]MH#:C&BFI?^cB4.WI@^\/aM9+aK>3=c\#:6@A;Wg9TY.UG2G2<]01>J
2b+R1O:_FDY-[e&H4Ac93YWd.C;9&A?PVO&O+@WH.9f]E5,JR9_IQ.DM1FL:0M)Z
?dPT,N<5c?8.B?RJ=PdF&NYfF+dH_RMR&5CSTU]b;_FC]FWIga&Zg=DI^+3M:-LP
3He^af&)K=&I-#Eg^PB5c?a<^G&<K0#G.XPH&=e,eTIPWf=B22NgO^W8VdS_Yg[D
:1/AS\@L/I]aKJ&,,73FU2^BV3_?D?H598d-IRR0SQVT;d4a>GVYRc)[gKH3KZUY
R=NFFE?L=2T/L9+M+=8Q,]AMa)AN9bGP2XQ6Pc19XU@_Ge+?<YV8OI16Z@&KOBLH
3;M^L1HM)_DgQ_?O=2=0dADK+O^;Xe;E,M]]GKQ?Qg8BQeCfYc2@X]_A9Y2d3DeG
-F+b_<9U<4&P<g7,\;F7VgF&V+:Rb]6,-_c+U&8b5/,U0&B+]^LOMYH4S=HZ;=fG
U1^IJ=@>E#2T1JE-_2M@EOS;^4X\__H8&19&@BN[-2/Q#2/f<_-_S#_fXW(<g98-
R@0T<AL5J@]Df,:NUE)?Og-Sg1R=5)<H>QeX_AM[E9H5\QCe=B4LY1=:]TEE-Z(@
6F7]#H@SPZE\6>)e(+O6Q>NMC7H2@F&g?T&CC,<I&eaeTI?MP;5-c2VE7IV+-T5Y
\)3aLaWBd]O/_IO/IY;YJ0_YZ06(SJCRILb:KWPSO#D#Df]DI+DWD^Gc\5RBFZEW
<+bN-MGDV?S5;L>VNRX2M<9E1(JdIO.0>YEgaY[[G=TFN(E:Z#5=<_[Yd=&+L.Q>
[3F+4Q^4^&--8/DLU+&b3B?1UC65#@N9F?B34>g^DWO)>ZBVS4dg9CTHY36>4aT>
,?+Te8\+H2c?Ne4\0>3Q]2-X8]MXWNO2<V=XO@M3KG<-J=6IFGO9Q\fI\2^DUb(P
^I4;a:Ne,bX47_)>OZg>KF]0URBJ6X-_[??a=0SUW\-=R#?IT#:.G^P1ZbaZA)5g
;]:^DA>DXL;[05^9YO;[OC#F2+a&L\S:VV0<0T23^GR=aGgKHLSLQcQ#=1AH+R.V
]Gc2W\/TbYI]4-LVa4_N>RE7?K_6;_:T=9C(_MQP/,4D<R+bC3A_XCG41aKQNYTb
1FX9J:?X]=U1TZ5E[3RE/<^1<@(?bR+>.eY=3dQV-c7I<b?;C7QO^SFZgIMG#4.@
<@-TZK)>1[XFLHfSJLV\7E4K9CGUS@:^3YRO+Y9\^Aa2C&>\eV9cDS#YBFG=\5;M
b,^XRNN07G5)[SJ+T)UXaa5PV&V[(WcgOb&(e2<&@OK4&QBMb/DWNTXS4BXL(cI:
Ca8U.;^,\gQ4/DJcC[6:NSKVd=XCQZ/,/@/0,)D#;=80[HfT0(D,IJV4,Je96-Dc
A]d:L[A7?)HNZL/P=@:2<E2.I;B>Z8)/Q__(NbRNL^g)B8IF[49\;BNJ/N>VSJ+4
ZN@YV^c]Q0aTe6?;3@4R1(3V0fUOI6<OOdG-@F\bJ@GeC06Ddb6)BKL\+6@dc:/5
N)^YB,GE+T.7_Z?]DREPU-DB1^S+T?R?)fcBPK^VLLaa6g06g5,(EA-0I@e]C^#Z
H)db:\58P2@OQKMH:=^Bd<;S;ALSC1K3GAB9POKZ,D37N/IXBU5fcc-R/LNK]J0\
=D9L@^/aFJ:,P]=6\P(c681E):A1I[PNbB;82U#JY2Zc:(FX?@+XZL<P0+#d&^-=
@RHgF+aFB7U3T4DS>X[/:^:,;7a+3.E5E8P0f65\6W>=^0]MJ7G8Q,aZ+=5]MJB3
@V07[MJO(1PP&;9W8J.,NIR@GV;Va7b+6^JdF?3C)HM2M\JW.B=1GgFS[NTIZTNQ
J#Y9gLFW5I9NcK>\]]+]GTa^AL6D:=T+4=-K9=ZLfG]>A]KC[D&EWWBEMPX?,.V/
aK(62Yg=5I^M0LVSBB\KUcK=cbg/E:][=G_FI)PXLX&f3UTKLgW?\Xd2.H4/9;LU
:DfBP1AAaK&IV7_ZaX&7gaNcTbgKN]Z6T#IFJ+.^0Bb4;UJTN=)Hc8af8IfLZ+4Y
fETS(4gJ/.PAT4&\WWOaA.38D3YWEM__;AfL5dX^a3Oc3FW&(9F@HC>?<g3X)BZ:
,7c1IG?+1:Q8CcG5=b&A/]ZX]F9<bSD.XA5V/_<JASE)WT@CgXE20W8.2-gFTC6V
A(4YL4&FDcR&(39=DOeF-_\].6C>O)Z86PQ>S9WDJA0DSF@ff?Z4:+=7-D9YedK4
bQb;e@[@?<a0ODLd/1)=HCDIb9UCa?5bN,FT2Z8><0YG2#IDCT614^>,cfP;MLN7
@-&A02#SK\-P-#H)DGc;EO^/gZ^O,U0;L.(e/^:\N[.T)S54,1dV-F:T(WG#d]?8
7?-@(@<TF)9C\60;?H4F5T3O1,]PffW2e^<SC<RfS,0aGFa#fF)gK#QHNQJO9=&O
]bOM[EeLGCDM4.+2;#I:\-<dJeEOVUa/0KHCeTU\A?Nb0/:._#/ES7;CQ_f=fX<Q
.XbZ^8b]b[JWFc83E9KR6g.6&0aNP]2[OgE>QV8Q<Q9AWL(86O42&;[[cXY,cWUN
bB_NC1eJbQH?1)47^A.cCRF1\<PV<eg0Sc/KDPa+SdAcfZZNUabBFgWLB;<N)DY^
@g[V\QDP,.2\E=_M^#LY,W4T_>#53e7dJU+J4P]9(W2410\AA8#L;Y4;GL]/e[Y?
(<Q91E<WMLc^9^^L,/b-gXeA<XgJ5R?]NOX>?C)P(\3QScS&1)?]E8<2?]a2KN-O
H@c4]><PFEW8;L5E[V^?UfTfLZ0^LLAKW<fE>bWUN7fE_.\8gVf]f#HR<G-G4-XW
R;>L=XT5O?SFI^cQPXb09F0_]cbXa.ZA/,f^,=./TgZDdDOb7(MPI5(^@=N\XaNK
Aa^?M\&DLPDY)LS2_[;F86dTHa\X&R?aZ9W5[SB>PWf?SBYNc)=)2T1AT\^gdb&_
4.._/5,g=)&8XTa@B=8gL7Zb=E3VJDGS&G+_USS>I)eG@b]46&f>^]5V_FS5^2bO
?AgO[DLa1[E)_S)R4bUI;c]B=L41VW0:Q/>_Q,^X<)3T5V4F/(EeXR[aL:(?@+:>
:N_S.H78OF##6@f>:.9dKF=8GN4W<;adHAAF53#O?#12a^BQZOS81=EI_1O#XWD)
a:Je;^PDPK)GTDO@?J9U\Vf?S\eQ:#A.9WE/:Q0<e06@2-)]O35/\8UPcb_G-.1f
UMU14BJ(ON5]6L_\e]:0R02Y\4ENEWVJ/5IJH;@&G-5GL#Cg&b,D^1)93]),9Tc1
RC<d-V.&H.<JcO\UJJF6:?L4Z/bed>@Bc=V<95[]X?._G_S8D1BS3]#4U)6NZH=R
Gb6]cN5T7F_eM;#ZM01:]L]58P>M:EU[Tg(=_eR@,ePHHe^SabM<J_ZH[)6G3^9[
NIgFdXcG[55DCEW[ZAJAQg<2>^08/Wd-OTQD+X+-BM;S_2+=<)]GZF&Tf^06Ia8/
6D>0IB1;GJ[+AWMg+7R5[GZUaUN\f1^,-Gf^dTcSCBdE?G>A,-VC6O7X#A7XZ0g1
><E>40[e29,)WZ\eTZ<433)&RG=YBcdJC#3A9,bKF-=?;X,]:#K&cBICEf-9V>N^
V?8=7eU_cC.P0gKP7d@:dSJV&6-((RO+Q_29:J(<.JKPJ^eQ:63VS2KD+?PCXOOR
Nf5<(T0MM<f\B0@Y^:GQ,CL+.Wg(IN]I\:540S:#5b;UR<LR6ac(G:c5CIFT_]a6
W-VMD_AVCIC9V>Wc)+b8R&d18Aa?a[/D_3PI.RRf0;]6J=MC>Y8+@VXE3@#IF[b6
:13Y/+/>J/5YAF)7_LaT5WO\#ABMV[6RVb74:=B74eKE/JC=dg(JJB?XCQd<-BSd
OOgM1+N:S&UQQ4YH=]@HLQNWH0))1,P&E&BPV;AWP5Kd;?a,O9YT5#BVK:6)PT&&
c_YI3BDLDWH11)\^Ff0ceX2>DY(@T80G08bVYUc#/7];.=OQ4-E);F-4&Ka^f@^F
C6Z6[3J9S0I6=N&7g2G1SJ_e:,.SOUSK<Jf8Cf(@5d44DQbUZ_8#fKe58P=1,1:_
H)@,[PSJ=Z_9a62/d?JbX+ID@>\<]DSeH;.GE/MZK6K^F=C>?5_7B3JBE@M(+^7/
BDP_^Qb(dROKf&L7XPeYRSd.a,2@+P3e74,55=F7PgZC1/,Ea@JEL)#DP/)47gG6
5WB+Tg3abT2L-H8g>g1fKK\3UgVabLEV74_AB/#>5]ac-e=Y#@-,g)R?IE32^@.H
U&US2&b.]</.<1+1#HSB&#d\e8#-LK\a<aY3.P,Vb&-:\YJHCUKCAE_G/ZIKEVdS
1VabT49L@THWWaaN4.+-HAMJb>8^)3b_A;#UE=[Y.&3HQHa\6>gURRAC67DMTD(a
F8QL7+:WAB,F/9?PS]QN19_L,A\fQ;#IX-,A(9gS,I9__G0>H9.1BKZ?b)L6)g0^
J4\JSAB/U^EP4W7/:>0N?#(L7(LZ\)F5MaCeY9P=?MYQRKVcM0/=F(8VPYKEfVd8
6NWFHUYUQL.S-6C)-H8QT&eUJG_-Bdg[bcA?A-@O//3JJHEEKS?)_5fSA;^LPdD8
[YIA<YT&F5bIW+P?J#RX39>?[8D32W4IK#Z7R<YO0ITQS.)T^W52d7GgK,3K08&I
?^;^VGST;_-\;(]@<2Z@-&\A06cWCX?#^3c1UU<bRVZdfgZU:6G&66Vf6:gMe\9b
0?,\IccWD+F.c3E=_N\c<ZL25G3.1bRJac&5E8PTD2V#8I:Y,1[WPVb=1)YNI9WF
?5RV03=71E;@C83\aF)^:S9FXYg/.K-gF7Be&3ECf0cI<IGf0((S4DQB0ISV-\YA
ZZR:f&QI8?d4ZffLE+.;HHC2NM8Q0KMK5^.6\<HI[H#fecgf->RWg\27<#V]MY;]
f3eB9?(6S5;e^7@_bJLDG1T?RKMg@>B#F(T)-2dO==S.3Z:H1_P7b@<+aFC:)]#:
0=3)+/7&P>W&)G>]=-8<2Y<AFAcKK47&VcgX1XScE-)E-7-MDdSEZdaDbI@C:cFa
3;dd510AcP:1WAb,[QbGb]HOXWSdR3^^Occa2df[+.;1TN4P5?&?JC6#PVeA2OgH
&R&S+b36_EV;/c3,,0Nc]fV#QQM=[e_&:N3#5WeTZVBA3XA05>03D-B@C35(H65J
f9]1N421#E8/0KN0L:\c4J/Q>1Z0:JgJ(YFFT/0,_cD1E8)O>PHBd,2(F9F7):=E
C(/-VIQTO11<\]/25/9R@,5&-JcR>D_[bEP;]<3&D8b70R3VQMRX?2..Z69].b-<
g>0aN5Hbe=fYU0.(WN/NbI>dR;\W?GWU@]^W0<HX6;<?B-VNOS-G8cL^QR80cXPb
b>#L[HbPd(+.FT<QG:NUc^A9??EI&6B(>FT737WYdURRVb7Q&-G-@:>C3QL,1#]Z
^DK.8_4^7?RZIA7Y6+4E=5@(Za4G=gdB5e1?;E1O.WY@U5>/,OT7BdSc-J39[M4Q
(,[W?a:6_cFR:+N>ZZ-Y;<-Rd2-bZSBT;NC[1(/IU+g&c5Z3RYaee)@N4?K\JNgU
RA]&-NHXH5Y=1L:WV9K\;Z9KNb1&+7,2XZ#498VJ,3^3M[#WgCB15;BK0PSLYWD;
/DbO_fUWfJ4[05ePNR)<&[Z//ba;1F\HVe.&\BBEM048]A4IUGQ4&WQ#0VLdg,/>
c9PD@8a][Yf\C#7X(3&aGAZR@-9+--;HL]<1#)3QF+5AU:.@1()75E937A2,1bVI
5H1\>M&gE_g6,I@9#.=21QfF<9XLf9YfbG=fA7(G=e_B3I@Ob5)057a[05J2\,Ja
T/LPD=)<-.KYW57S#@SeFX9?-f&MJZBS@XC@,TD:T3O(@7,OIH<^Z10X_,6F/UVX
bR0=5PEd@O4B8(8c=eYBbSABK7f>1,3?.UPf5]=W^08b\EPSG5A:85LGJ[[+\HQ?
2I#2b1[.YB+R6YdH<V2LcdHf?DPLgIIF322c:V9D^4INE&VR<9Zab(a--_Xd48Y8
85HI5[f@f&ScLJSeRegLU94/RU&Z^e0),L>26AZ@C@JY6M:c_,5XIS&5KbSa>1.@
PWf?B)b3a(1U5?KG6<>RXKT\O066Va_KKYT8W)/641F:UFLO)b[R_/N6S,LZf=X5
;GILf+2(PA#<32B[_WLB#C11Nb_I8Cba-b7VCZb1eDSIQX]U2?fWK3gc8CaC[]SL
CZPPV=P(H\Td,H,)N8dA:@JL.Xe+#];B2PT6H:[eDTf>@eVfQ\X)I7\S\9)XZLb-
fJA#M/6^OV.\0aO4V7f.;WLV)IfAD8+E2CK17b\]ECJU_KNG9?,R03(SeXV<OLJ(
2(g6XHK?W(KgReN5eC6K+HPeM;1T-I[TL8&^3GWA218gBF<L>\^QV(CX\COQ:DW]
RT:R#7_\cQ4:_V=G-49&WKba4..<7]/[LA@QH3)##VI&TLLgUA)JX1JA00C_66^g
)\9V6d4F,VLg.,G?^G3Tf\gPT<PSJ2;gWPCF=55Q&U1?K&T4C0M]8Y57_Q:g3d9B
ca_gg)7dIHMZG<C2If4RT#T5F>^B):G4TXCC1GEE7DIQ9,3a0PdQ9PKU,-<fR.1[
Z/1_30ID^d#A7TEY8cRUNM\PCIGf[G2Kc[-]W#QLSe3b0RH8#UX5/N5HZRCIAHM;
]&OUcGVR=<3a][/J)^B:Z.P9c7QQQ=INeKD]_4W&B<9V3AA5R;++^X=JUa>DCJA0
,F?LJ]bI<[NgF^+U-(?@3N:]WHXAG#^TOA:JUTd=-4)@2,GHf#EKBY<=MWF9MP_=
Y:2&))F>9[AB)-K&(^O\_JLc:L#g^X5()&WSbbH6B>LefGCF8\^3(#5T&YbI0aF0
V7<APU()H@KDf--1&XFaLRC\Sd^UZfC1?#eSP;4T#H-UA0G1Q3?NT>]T)W,]AF3?
0=Z\Z]4WGK1Z]_:J:;/5H#F+5cSc[(B_aaL]X+\1[cH>@E3Ma:E,OQ/HH;A7+9LD
_bC_1Z?,f](&<6,AV0FUMYX(4^C+CQA9a_B_++N[.T<L,/(;,5&Z6K[IX?PgII[0
-Jd&^3-=MOB#;16Tg,E=2&>(Bf9Ga(K_Bb&[U3>/_]1TbabR6)G0Se0)[YH/3&F]
B9eCe)fR3F5392b&YZ5+<.JA,3>/1N,Ng?@UA#^.H@BdH:RS/>SA^7^gK<DVJ><c
J@-e<P>\EZ>g&cbK2DJ0c)8/79#MGPf9HQ4>.3AVQ2\+A:/_g&.7I1E0PR@X+dLQ
X>++a7_W>LOZ#W3P+?-7)[Q,Oe7^MG50Ig+fJ&L#PSeNdK4V^H8_J9\IWCgGcC<M
cV[aC45&e.;KUf]QcG[Sb61<E94WIQL@)/K+.GfX3F(AJ>82K\.F9fL):.=TAO;.
d/0XHZ&O39+e#6M<((W95FCD8P<6VW8MX7__GRP3T:(EON1F2(]d^[(<S3-(JS8:
=(A1<,g_]TK:a86FNH8^gJLVPFSdU))>dV3_K]3&a#-gACcW1Q0d&VH>HQ>N3,eV
7)0ZABAUc@)-U[/=]LJA7^.d>ILX:+?QKTQ3,SU;]U&K:Kc2S#SFWA9Yd)ADK9@J
BNOE4RTJO-P#7@3@K_g+Gb^@MSMM/1d?;g>JX<Y9b:dFN79OT7)+c(BN00DXY,;C
WP4::TB28.1[a4#^S@K82OV^;B@Yb99+A^.3_IaUL24;X^]#8GR7W#GK.)QP+[+F
5a.H09>_U\F;69@^HX/_WCHYL3d2GQ,4O<gDN\6d._RTLfC;fTZ+1/>,J@1U8\gC
39R,8UAc?3./9HgODLd7=YCO\A[A597/&:O^6K\8H\8PUZ.RN^fgWZ1JLc/#Tf,S
f0?X;c[G;I?XAe(N(QUHWZQ#:cBd[<3_FfY.J;<M9#7YTMH6AEY]S7faW(2N2H@c
/E0RTF-@Y&c\(Ge/OF+GMg>.N8L2@BS,H(bLa\8,R7([UFJDUb-KDR=X>-gdT3C6
?9Yc29?dLCM1b.+W=/NWT7D[NNU1gS1)U[.UJc^7_-X_RQ.#==U/>ae<a^1\<e=F
U9R>0:A51C.;8YCX:-Qf[I5KM]=2A4BM>gPdMIJYG^cOT[Z?TeQa3F,Be09F6IHd
N_b;fEU(.@B4WaaYa<2RXS6OdV82@e:4Q6=b+dYOZTc=4J9f7=6UH,JL?)[XBJ?f
S)MDSdgf7J)5@c[B=H\]0+YMS7C=CE6a?VR4JBK4<=&]3He^,:[=?B7K>2^fKF7L
<R58-[;8UDAcH4&(\e]1_M,e&X0+=-_aOL@1>D/UK1JW][;S<</2+LTZ5KXcE1GL
6QC^OFf,\ZV15NaC6_,ecE,)UR_ER_XT_O1JcVK\=M?8H1<F_E7\:acMQb35Af:(
1(KXW+bQOf)JB&)M8D@G&U?M#e,L?<c4&UW=:.LE,VA6JFCJfeC,O&)(APL3[V+I
<\T=NE4<V]5eYA17[]Y0@N.DEC+>1ON95Q@K,817AE\;<\OcP47aO,RCTIMZ#aGc
G0).7b9<6^E:#)N;Bd\X=Q9CHI=cgSH#)f=f+Dg=9;Uac=R7Z3eLT)-J[6YA:<Q7
@SE\CV#c-GYD1b]NBJIAX.PM<:GF3H3Q,/7U>;g[c-<>::X<4Z:,>5Rc6edeAA6O
>.Qf5CKRS54CeOe3;@O3N)E+YLA;H4X.OcJc96eD#aCPdIa-H35=&3_XT[,_:G4W
.<:gG_.[J5]#54QFZ9geMRB2F-4]##>:[?RV.abK)00\N.&)=1::f;4Bg.Q[L=8P
+:V6@?)PD2[U4;N<._]KHF6->F6ccY+0(:Rc+OAU6TL>I>aWe<dKH@0S^YP9d-MO
#-C+0R0-V.;CHJ\WG.K<]cITZggCV8<54ZCEI@^7AD52dI469^0#5-1(:Fb5<OSR
WUd7HTd:b1>7J_3,PD4N/[?3YXf3WbIJcd.MA_+:c2^E_HgEX[3g_aL\<?<(JG6f
U6TD(PKY@cAbR.TO.JRJ,PWBO=ZI4HLb_0HTND;GgV,\&W[8VE)2VB?&TJ3>?b.X
?e3c#-PJ1<\V(_#XKe:92d:(UGf/E_)87(?6L<V@dAf2Xea::+)ab#UJ^73YEUX2
,a25O2=VC<1I\V_[PO<Qc_-NdJ_;5:P2ZF>F=;)4\>[gS#[TV813CfB6VLK1e)]4
B3:<9A/YA3#,FGL#C<RL4RO381cT.KMe3ATV^?c9DM?fLReT>UVg6:eR8#I6OIT.
;C1E=VPP6T+F]A^\@NTCV;+7MK.ORJ0,6VRSV\Sf:@P_5QHI#UR)9&?^X7I]]Wa2
99)[+FFZ_gLI_T:+G[?7:e/.c4:Q8_Ee^1(T4)\;T#/UX;Xc(FIc3L43WMYPN:K?
E-3DNb\:K@)EG:eDEV&<9MG(F]][OXQ@/4c8g\BK,)X\L/+,+/S5@;QCe1)/DQGP
6VcHA+@57e0=[<AP&4_2YA,+8-N?VL-_\_@-(]Y=&0-3\g>X8dL<0.3cIAH5E7(G
3.4aB@cbIbB]::^HK<,UYEJK@TP#,gEY&RYGSfLRA2X251C#R&^LU++7HC<Y-[WR
=?ZMFK\D3#V+=C&MbKY#O^Pb6:;>[_B,2^0C81M[=URc0.fH4HbN-HI[V4IBc^1\
3d?D/8CJXOTH.+<^W@b)REC+X2&aF3]F_-PRAgX((FCK93SH\NSe9,C&]8#@U.^K
bR9Zgb+LCf<.Ta1\6Ud>J-ZPAWeX((TYUeV:X.@#7@-+e]&DQ?WY+(;aC_KY@\ZO
H@U1Jb??6/:#FV.;e9_Yb/Z-?Pe&UX>MO)2Z4COb>^=.K]W]c2]IRQQB;\8)LY38
-=:B4=GC:QV8^MX_<[W:7H,2F^H5?<8.=3NaEB>Z)4F\W=/:^XO?PVF49@]W01(M
I=Q/NGRXLM2]>/9@MSdCTd,LE#N63_Yaf+2UC&/K7]V9PK+(7-2<Ec_=NI8XfDG^
U)5TSC,1=U8DF0_Vg;IT8@gIT9;):#TRe2BUb/[+A4#PIP<dB_AJ?F+#?JSJcU)R
<F,_;:&,)[Rb9X4LIe:AY#gDJ-@EMQXQEP\UBG(aAVJDJAX&\aYW@E^)+L,c^deS
f)Bfd0B<(MLTaSA6U3DB\bL@)C92I7G7aU.e6K-MX(V)HQg<ZR:KJ+E+,A^87IGJ
[EMFg\TT8NdS/.8->KM6ALK@A<,-GLUc;;4+e?+MI?.,DD;8BEPB?)0b>VcIFIB)
\0\ca])0S=S\1CZKSD2(^P(H5=PMB1d]384:,GD?U\^NL9fBcSRVUNe03Z/5E(e9
EETfc6B9N3>H=>g=e[NIKa?O0PNTISdbc\4Q<C0R,cQH)\]2G\F01=gF.YQMeNgM
QNF9>:1(dL]1<a(eR??-KdPE,XdaOJ:QY<X7CV^>Pf_[T(X;G;KQ338?^&^b-fEY
G&)\;05J0\H3-=&[-RSBATZ&f1LBNK?PCQPO@ZN[IE\=A2C,Q4SJZ/\N.YL&\S(B
eIfYAY3S-)61I72G6a+:Wd>AB5&D[(\&W+3PB6635aa@?@B5TT@J0(G#V&<S@_@f
YH==H@,H9M3eMc6?L6WaaDB(#GB]fCG(9/XYgF=g..G^JO_-C:D=W])gHB))[X-R
5G6YQZ^1S+7N<:N:>HFC1E.GA_0V[56KNTZ3FG;VY4>E[U0eU.=<LNeb+3ZNG:6g
>&;Sb4@OY1(/QTeS.F0eN&AEfO@)(MgXFg,;#72c;FD&-WcD7>IS=W:<KGC_1gPO
\)Tc=/([f?E21,]YIZ##b>^;MH_D]X_LNH=SC6ZT86@54:;4R,=7Rd@CPMI\?fE=
>SV[1a<\2P:LC:Z.:cKMOaOeHJ1,ZHV8W[+CZ+33NPX.OEU23aR/Fe#CW(?d182c
CL94JD=\73+d:+OG]IZR4H;J][0Re/:@(W4_S?Z4#V;CWcA34c3X?JG=]/[+,fL4
TaJ\2P-4^G\]6DSZ?N66P2-^EM/YWO=@6(?VgL;?CSN/[JZC)&fO2c5Ng6XI_.Ed
O/W&J(fUOg=L6-TeAH44dWIGF]UZIC6,)56&.>#48I6d:\F3H,/2H1@VON?H+QGg
+6gR,7JH2XLgW\5OZ,VM2T-1-U9d\AebLd1gB4-aZ?#GH)C>@,b88c5bNKCG&8R6
>(]0\AY(B\1[LTW4^b>SBHY6eY06\&YP9)P0LPMAN\;Y@(cQL654DKdVQXBOd@GU
^^PS?^VEg;R<JfFO7>(gf2MCf,bY8C#C/,N-=CDKJYGR5A2[G)8UO8.g6FAK_\?6
PcW2#TZX1?SS@Sa;W+YFABG>^VA<KR2JVV@ZQ>/:aJD2,Z;?(b<bO:<],H5^K8JR
<Q\&I3NScQQG@G,Ya_I.2K@85.&7c7Q[J1b:F>CVD#+g?+1BEeQR35DI-[#^<)Ae
cTFEa^/@AdaGfbKa.6?EDe8W\;^O,>U-H-2-,:f1HJQf[<HV:&B825?g]9TH4=1Y
X8U_&[;eb)J7d)\_9=eNGD[(FaM:13UMY?\ef&PVN6I8,848.c,GR?;f-:_Ee\(+
A7ZB6d#C&LQ[SBe@U@.1+\b@E)8>Jc18;9T9c@B^>\O?YV:&B1c/\I<P5aceAQ8g
(HESL#Y2BGBNTI.-[e#D4M=WeHCN[gNW:U;D+.M>N=_ZC-MH07,]7Qg.44@8QZ^F
#KJ_ERD,8,-GL>0V\=3-04LSWLS4IJ@;fP,S+&Y6ZMd9fF4)@CK2)R+4gZ>d6]RP
JFLd;JN#C[\JSX;5Y&L6L1ZQIbLCT:Ob9/cPBJ<)UdCM0>4<64d;;MgK#P\I2df>
JT&SDJHO;K&d@;JG17,JR:Mg8IG9dde0KQ2a#YUCeDU<F0+QD/+(VgEK(>d;R8K:
&=WdIK:>L:W=EIN)&fgI<R))&I@SQL>\=Y@GE70bg::9(T3LBZ_=X(ZKO#C?2bMP
DWYQ&QK]72T\OL./L^/#VGY=0QU3O#\?=9^]AB=FH5NCcPM,/3Sc;37IEa]G#RYQ
Z,1N+(H7>bG>Z2TZ#6cZ8.-C+3P(VBTbEOS#<OU0-6EcRO+e;B/C0K-V4^XZ#SXB
;[G1_Ae8V++CfLAIZ_1[&W?0PW:Pg@CQK)B1S.e:bE38-+A.Rf:cTET:E+W</_F+
d1]a?YN)>fI?=MDSC.Ge3M<e8Lc0Q-Ye=HA)bVSQHU[b5]0d+CSMK6_XL@dPQf6S
_Q0<,TH34CI],Z338GWgQ-\e0-=.XII0+YAD+1f#Z.\\b,42RI,;H2:#3VH3f7FF
E@H?7F>#J+e7;N^?>=7(\&&[J^P0;WUHX:)=_=]F<YB6)fd1gY6OY2>&)]P0^]HD
b<a;/WZ^-+L_=J_AdbfgZ?U.7?#=(O&=NY_+/KL:9f[e<+Z^H<3U](1N-b#RbeTd
g@(fW095LVW(-AS^NW1d&bG<aCBTg]7C3JSTg8(P[_813Y6XG(gO?f+T1g.63Hcb
LUJ[,BYT.&gd&FKed4cAD;/EdfC#KD<T1W&9e+&)3QMRVfDS8D=OPWI/O#KfZg@,
&RND.,)(DcfNVJ\NFKcEX+7+b)N(29>a,UF<MR7<)_b/;7PN>I:#HaK?IB>G:#WS
^Y^/]2=-Y+W)RU.\#XgW>0?2+_+c9?>F:ad@RK63UK;N_;(@7)GPDN-Z\)W_J3.O
5e#MG]CCfUP&ED0=R8@/;.9.eb.ge<E=bb--ZS=f:;C<Y-9a=1e-E0<#Ig(05#)-
I_/WUF:)9?4AAd@Z[]BGQVM7QA>[K/&3-/:gf&>S<4MP.PIV&TV=dX[b]-3SNfVG
ceH.Jc5Lbc#QL)66aRML4a>=<2]Qd:S[;[>H:XM-+/J#E9bGb4P]>TV2G;T-\TR0
Kb>9<8<f0J3I0S\AIS:D79f;V27\_01NXQJHFAOND.ScJC.RWfQ-FCCOH9+>S?Pf
&IV,3Q=bUX8NM]3)(E73#C.<7?I4IMGb@V9((]&49I-E+,R<UT.JEQS-K2([OdeO
21?)KJ;I;5R2[=2_#NN=0NbE(]]5SWcRa\+\5<YObD6,Z;NDJ]U?::W67HebRe,/
0HfLH.-.J6cS)QE.WP\6&3OYeHRUZT(-I1;@B(3#/#I9N&Y8OKO;;.EX,:J_IIAR
P#H<#HXU&A\2<F<&D\d-?]4P\/.bWYQGR^\AEaG<?(O_-RVX6/V)#^4C0+4PBZ)1
dEC=8A8.H/6TDZgNec[TMZIU+O7I?J#-V.bdf4Fc^ZgO_OHZe5..?(F&<_,JCBQ5
LG2)87L<SC[HAFPR\)/FU=0E++3Z@;A#ETJa_#=#U_.R,O-D_Q;Vf+DQMTeAf:;R
:&DKY5G-3d=ZZJHf-E_LF;</Xa?,DK[K&9L)]M&4:FZ@d\_6F/gU7d@gWY7#MT_3
6gJa5PS]LV\-1K0fK&IV9GB_&c+f)@7V]B.DZ_C^ETR+)WgI?/K?cG[O+7^E>W+-
KVT2:Bf\-B2_H=_^8LV)PBL\&FEYL;.^eXT+Pbc60+9V/H/W3eDE/;H56(d+EeEO
_f>W7<^+eOYH@.US;PCIK[g]cH5,^.V=/<4c4a.D_)6KS.SXG)7ffM0dFLGAH9E7
^<G:bH.5=[0X;)OFTTcVGDOc&?>G:KdZ@J&_+B^O/5+@R:c(RJee5USN[S^Z#[[S
(]SXI-V(&AX6HUN/e>bE_CMbbVfRLGVZaMd;GUS0HP^X,e4.)K@@cb2^/<I2&3^.
Q+JMgB#M/W^0C^IZN_=>2S<_^0G405R2\;/W+T_HZ^,S^W>JYE9fBQ;K8@1TNAd]
2JfHD3XJU)aU4ON#F>T87Z<g<)Y3U@FRBW)R_a5Z&G)I#-/-B@E]):?46GCZcdOY
.=/0/9C@RC;^7^M>#JF3B:RC+eZF&QLLA)-0NL9I(S9TGBgCEC)d-J\Lc&d<]D)4
&eO-=3026bd<R?U4=39-).Kc7ZSaGbbRSS::+DT;ALa_Z+5WQ^RRUH+9#?;:T]eU
_5U/?+ec5J<NWd2O?2U<)FQO]A6<HDGB&]UGT@V.DN^cJNg4_KP,6aKGV&W5;>:@
\>E+Ja-:c72XN1aU#aC,HZCC2TW#Oc;C#ZV(0.W-9C-4Y+AA,D-S5LTW2d-\+HZ)
MW#0B&J(T4PG^HJ)731Y/H[cPBJ3KW&g?ZT=5L17E:,>bT9/cZ_DW<]TR+@9gO9,
>::e>R,1SK9V6_G<A.2#7?8aGg-3D6<:[N,FBB)Af^,9VD>ZIcaRYU:?R1b?ORR&
\,F82B]0;<=[ZO4/LLD,\LVG:cSNH01BPQK,:]I7JBYP__@=^C&IgK+JS73J3G\\
Eag3J5KTI7TTF=#IZK:1&^H37)9JH@aAY<).YO4Y_S:L>aF/H+Y7^/2=ZdVCd6I6
XPT[6K=>U8;GX3S6-2BO2K4V#Jc;d7>B2/74I\79?b_B_U5QggQE4V5ZC5).NcP^
?b?Df_V_<H^P+C<&c-a<O.G99SS)Z(1Z]b.9_]#J^MXT:QR6L(>L]XY.QQ,D=2\M
f[V/4K[(UO>L?gdUO&G#8ecAb5^#7/069:Hc2HGUE.;U#8Sc:H(47/R[4Y7JX5dY
N+T8C8>EPVf^_6c1bcL;Kc<@0IPcf1,7AS&E->Pf#O[LB27/[&8;+g+?VMUK(TZR
fI6XT8UM8,gT(<?>]<PTX4fe:0b#1O>1N[?-H>cFQ@?Gd?Z_SGE-:IY1bNa-RIgT
(5T3LNcW0]E(Pa(2?_6^PSLeK[A;U77gf^F53339[?]KFVR.WB.+1ZR_>M+VKgc(
^I:^2_/;&4@)\>LC[S9Vd5HA0^5Q?4CQ<dM0M:4^eO^Y)0bI:Q[?M2:U14I\.3P&
;+gb,/^X(=a7Ie9EeIe,?S=NG/&abZ]Y0g?=4VN2WM^_[gcea>^\c7X]\OM8WQN^
?P[X#<0fLS;PcY;MS]QGNN17G^Bc?Y(dFHY;AgAdNNJ[G(,WYg.6Z1G^87>)2B?&
WaKG#,fW/+?J\MeJd8>RdL(2b1Xc6+@H#Q7KJcH/[#>;BAYGQQXSdX7K9O+U;:HV
;^@ZI-Z#\=ea,FBBa;.6DWaU6b9&9Af_eMBUZdgb\II5L@RGO=RO6ROPMYbX4VSL
.PXJ.TcIIc(:CMY)J^W:NNU1R]E>ZK^-L0cMe.e\(?@U/A\-R8:^7K]R:-3^2_EG
UK\JaT@D/,TY_TT9LgE&TD<2)aG>NCQ^2I<Z9JG5-gQ5=:^(f^567)KU0/e:QO<_
6@;ZU=9:W,XO4V4OP/L0_;_OO^]?@7PF0+T>KOU=@=NefKB@2HRFF^C<(F8?b>eS
[X:S3H?,6+[Y]ZV\TIaIQ]FN\]?cV[ZZ?)gA.4ZY9cAW>M5g54>b6;fQ&a]<60^f
N+J:)#ES/>(6I_dVIFI7MbgIc(V#<LTHH.Uf8WGOZP1QXJ+@e<bEE3>09aSDA<[I
]/5(6\;R53J<#7>B?8^?F,O4#M0L9g#A&4R.&-&AA);RP^4]C4Z:57)\KN7,1P,^
Pee0f.[e,ARWVc(SXL\^V>,ca2#ZDQ<_2S_8-,WGE2)TGB4d?DO9b0>ZUC0@](fA
Y--O\\^X)2DC.R0P;aDJHQHH9XHVCHD<-YB)d]QN:#bB?.:Y4c11#;>5bb:Yf39a
QQgO(4)6K7EQO;9EO-GT/;EA_E&L/8>Q52=J_G[811=#<0IV1-+(&b1@c:PU5W[S
G>-AbXfc=\?1#4HVH&c/(E^UWI?H-,d@\&eHBB&+^(3,2)WZ79gH:&1@K$
`endprotected

`protected
DL+H.=5L^]FQ[HP98J@GHH8BcA?[5?V5BOIWJ@Q<YY)V(C#+X_?+1)?a</a8XLAH
0F\>.&DEF>Z1>Jda40ULQ8HI?=+=b6[-,Z6@SQ&8dV3V&1ScIPGg14dgcgN\O=c6
K:^\=5F&:L<1+$
`endprotected

//vcs_lic_vip_protect
  `protected
FMY:/V9<AJX.AS.V]g_YN8XGCcd=94YUE-^MG<Cde[.UVU.]H1Z=5(YQ5&XH[Y)7
SLE--LY;cC_=0W]ag4#3@OEAH82d3#\L]O;8\+:<gA7Y@(KL;Y1E=.fN]2bAZD.a
;+?34R7M14fZ9U.006I82L(^<4#8K8,D:WeS5B\M&]4Q>?J3G(@.(QU:4A3F/V=H
e)Sd1W7<1LD9]abW2^R\C_B^K^R785RCaH_=g^65-@,O>53g[KK[WFN^fLAU4Neg
T:@[_<RdE,X[cSBc^gbTZJ@AUT3^.A:A^,^@<1=\6#AO&8EQRN]GdB1=\;#F^;fP
NKUNU_@#e#M//b8Y<.CGX.99Ff5&eeB^\.I^Q2RKd)N,CSW.P.EGE2K\->U9J+#c
&=QMWQ1M0@NY+F@(+dOX2H:.K[0^S?+Cc^dK9#Bc29eHd]=a1[VE4B+#6@R^MI:D
)d)SV3]8Y4ZHOb=T8D:OMKV@PNP[Q5([KP#Q+d6S3L8-O;RW7#C-(H0PS-<OD;>N
6beYfKO;<;HWQV[Bd[7U4BaR_MRK8D_1=H5XVJ-,><CRda4,;WFWPHU(P@QV]9DB
ZFE+e.c^N994^=0b1gLO3&K8&6g@gVS2&1MOEQ3.]<=QZU/fP,=6d-@CS;&H5=ZF
;<IR5AJXP;EQZ24+e+>.Q_b]-6>CgB.6N)BL).4#/MHB.UQ&g3APEQF/)&eHM?KH
6c?M[NJ(O]5DNN9bF0-QN]S?^<T@@],9\ePY?9U?eeQcdE0B7+LKC.[J?4YONRW&
bJ\\)A;1<&8//;SHga>Y4-JCKa7=IT87[c+2aN2.#(O4c9KRC7ac+&1[XG\X^Z+B
&-,6U0DH/E2R>fAH3M5?R^e-YXZ;R-/CR2L[2+g=P[7<]_,\0WD@D89aMLE@;00Y
GJ]&;]4B\aQYR2\&YO8c(JKg6]He,].9LOW^R;H)MKVdFZJL?G_UDX3\(K.a<4##
Q&8S.VD@<Z#b2S#\T[@FAY=R5?(UCHS?DWEbH>/>(\O<QMf7GK(OI92;=#K&3Y8>
=dJZL0GT?3.>Og1>Q3-+eb@edeMB-3SYFWK-;gC-II\IZM[2/]H^/[e+]@cL[E:g
Kd>f2^\/fJ4f.80+>S0[N5D].)5d4)OXg[=G/1#J8BT8-].IH29;dca.=@IFY+)A
bG5-/S@9F9OadgHFc#&=ZeKF\X9I6;[@A(4d#M?;BSWAc3.3_TMQ80GbM&a8XSNO
JOKOULOQJDb^2+aV?+>/2:6.?N.DK93#XVeD+Y8\HVf+P#LT8617EHgOf.E&[gLe
HLH:MgI+>aKE,f9&@G/0&N1<5g=X9L.Hf&-.MDJ6<,CHBe42U<:g;,_=]=)T6:dD
I;WGOEH2AM1b_9@Q]9RP-TZg0[U#d/+EeUa[aJ,LT#7g@@Za8<Td:=+=D1#a>Te<
b#][RV]-X;+7dA6YgNYFb)/33.BT14I?g(B>]DYTfZO7,bUK.CC1K<VddVN0Qa8/
)@37BHQ2I)F_A@THQ\1IQe=^eI?N+2;2/JNA+<>QG.]c?[50d2^AA+339cP95&/R
>N]RXH]c:R#H&,UOd<77JS5[Z,A@N.\Q/_PS]5gf6MPf@(MReMWC2(=Q0I>^4O)S
NT0e9f8QWPE2PA&7X3)I9(cd_GD46_HPQ_?JOHG=V,1]-:=VJU#Ub8&e\/b@3_G^
F#T^>7>g093fbFfUZ-9^)QLU@JQ0(0XVM.)#04+_R@7(-GMP8IZRMGEX>?3\;[;V
W-@FgCTU2OH2XH4)KJ8^5=S=.2Z9R/A>#+V.=J0]][fTFXAC;g.MCEFEG9XLA0XP
8&S,+L5T4]2XXSIfZ_Z2I[R1-f]EOQ6R6@#GeE2MQU+_K@JdGZ94Z5&W\<<CfBY&
>)TBI7]>dEE9IC/7B@bTA:fSgDIQ^V<JgH:61MANSA98(>0&?]QM;Y?^Kb.#Yb]@
_f8WOQZ?=)T6T/SN/f(#XYD^P:N6FZ[FO:U/A=NT)XCOV(,HXEQ62<<f+DH;,OGP
YRT_+NfC1(ZRM17E=^#0/LJRgMTa6Qc,UaV2;3T]QgDHI9:.SYOTe+&_bGSOT&@+
@<6\&BJQ&[2>+LI-8F^O5<2WH\2;TKMaf2(I41KHMWbN598T2LT&R--_&N_:BcV3
,+[JM+I)2R^HQLI\(((2C>E#EH3a6D7H6<IT>cPKPMD&P9>Dc-4C:@]@eA#:_2gS
BfVIL/P&3ce7O7UVBd]DMgU9,#J[2N_8=C7J1W7=3=7:NYH@K6VS8VM9^@(UCg2Q
3=OL.>cBTMFKX?:@=GPMWXTgddF^_BR9aCRP@C+^0CSK@U3GdT2Ag4185\MTRN,\
LW-D3Q.EgCcdE<\W#gXfUY]L[H@EIO8Y7BMAP4STM&5#V.M+9,<@H0X+g\U[)84&
VdacQD+A<M/NdaZR,>82bCgR#7@,:E#4f_aJcB2Ea4B04[6Y9>XB07Z0K[W:5:MK
#^YT3H3[JBOW/)9<+MY&?=WM]C8e1G0.(BZgS\[LB]/d>D&dW=?<S-+]S:::W[fQ
WP:C992?/1aD0M3\/E]Q:><)6Q,a4279Gag(CDQT<^f;BPNUHLS-\]U/(KDR6Pa\
7]?\85\5AMHO]4O@898E2/YaE1I[PF:9WQbQ5d9[.4OC/F1bKd1(VW=;R[N1DO)?
[VE\AQ6AFP;#DdJ7W:@V;+8-)6A:]aS&Tf[]+E8ceXZH5aKaFB9YB;G3E<eP#>[L
c:X(:?/9_>[C^=)#Y,O1#c+E9#b,)(a;+O[dV?;PL9K@@G8e?=(Q:e8V<7--8]&D
FA]eW2IZG=F=IJ(:4YMd.:5R22X4H^]6@7(^f][aP]VKQSRG/\g9_bB<+)#8gT9c
\dDDbPLSCcg^.L+Xc_DO\Ec+LB^M2E81LR9@4SPDS4.09JFRF<Ga7=<VVE69?#HO
K)2BRa6MIJM441R2c:>cb?:FAfJ8ED[)54GNDfIBfV5O6Kd=EEVd(DAX+aAE8[E?
Y\O_R;.\^;<dg^.T]N3dD_R_A;O6B)Ib^7;A)VLf<GbT++B[dB@3aCW6Gb/#G+SF
/NN^NP40J/?4EN75+814_@L;\EO63@b4S46.?H6g^_4PI<B.@TeFV_M&XB2bKH;[
WA0.GQfYME-Jb0O^R4A)HB>Z,@Z)eYG4JLZe84Y7:]#98-(FZ/DEF67MT33BJeW4
^+,LgX/\K-P&1XR8HWZ39X(ITMM>H5Te4.1GT^0U6UI3b&_65/Z,H&CMSgYI:cA(
a9PM4-#S2).-2cG?fe\d_8(K)NXbe(OEHV#(S^RK-C5bSdR=WA2dX1+cUA:A=0(\
cb2ZVH.JacO.62-OU+)H6IE-8+23#:/cBWFJR]Ded1GObe,XX,Y&;J(WGIA:gE99
ZbENJSQ]5bD=NLF6:+X>NCcD=SL;5A2aY52@d85RfgcZC[IL_CDKS<RAg]WSBeX4
d<S2b1>,/GB/M>N5fMb:&K;VNJ;5,?FRJZ6eVd^JK((76OXC-RBIO,(=;TWX(TCI
aL-T=[,&B;K5P^_-=YJF0#T:[WM1CdK?ag;=VK:B5<A._1M^g1@GHd6V<T.g47UZ
?/g-TMc\Dc96d4&V7_B=Y)C^4V3R=]5Gc##NYIDKHUXNR-:g.B5Q@gMZVbLT8dG;
RJL_e[c,^3E>0[CEE1M:-.gQX6@?C:/4N\(MVCB1A@R90>e+,\P+8[E:E/ZL4.VP
,4-003;C(DMI[TI[OK7</B8&._22=MbL8H4:YD-C^Q/G#K?PQYD6d\^g7bDOB;-6
L0BR2:b/PcJ-;^Z2.fE6/<b[N#WFTE5F:PbBI(8+cIE6fI-NCSfPEeDWTNB#))>f
X01[IL/CO(_(\GI2GaJ9.e6GYL,/Z3=5VUABf4QOLPa(X_+MMVJd&C+5M.\<9gNW
3g&3>3JBZ:0^0CQX[X,3=<Wg&cWNdEWL(QE^&0<YdV37b?_H&C)7-0\[F7VP(4T:
^cL\/Fe)9g[HH_>33<SdW]MY]@K)Tg/0\6Y.VRcFH?D=0QeY/d0-0-XeU&QF@^4B
Ca5DE9_EP-c+DFN6L,F@G95MBR=dVA:GQBRdNbF@2\;35/JgS158C]bSQ/:IfN@^
=_P3=cA,DTc.2K=5XQ_&;5G;8M<<LFdZ(P67<T.\22f-+^^VZ?R/LH<N07f)2g7F
EfOIXMgY>R0IX:CX>:O0/8&E(LJf)e=VEcd,Q-#,[P+/)<=[YD@;GE-0L@F&6-^^
X[TP,.\YHJTgK;99;PaI&BI]:Y(e\a,f5[H89@8b@O;+34K>;XBAP&^^8^K#GG1T
dWG4D?&E0\4IY^;5UN1>#D<e12=&8F[S+#YGD2-E44V=#d8+f<Q2&O7]FD<)N\:V
T5_G)QeUgeK@SGRVXf?EK0.#b0Rf6NeRF^H=95b[+Ia#F;0PWUc(?81)?P/d^#EP
WY/.W::#:&-.^/>7A4^T[5MPVgeVS+(>5Q)Ig<HLU2N];GTB\E+gPR7HWD>8WO6Z
&CRX^VGX9,9X<R:f\#G3XEQ56JfESeRD#G0E]1bc\YO-@fLWe-W=g]R,@DKXIYPG
#_(26LFAE6]e>WfaHE9Y-f3,=.VeMC,2/Q2>,08J0\5a2]+UYfRCUX]P[NX(L[0F
@9WB9fO5?O&>_f5X4-We+ec.Q@1;AF+R]AXHF5a2>/XV@cHDBW6J.:#LbcTO&Bg\
9)(2fCKQJR:;<A0VX,ELTB\P#^aZ6-PPN/:TV9S^QOZ#,>&]fEEAQ4I+.WFJWB_a
-/5D(59&OR:A&;g7K/?Ce@ga35XG^&;5LP[#)bF@A4.GD1XJ>ZA>+&LYXIGQc1b,
V>^2Z/[5g8/<Z-<P;JC93#(aH#=[>W]D>JR?1S>?K1MHP#9)e;d_UZeS.O^GMaN_
T<HZH3GUF&.Z=H.8LCZCPAa7V5^:;EYA0MSJRDRY]23U/9V\6=dcB;2A<[=d.e9-
gHJ7H&/]Od4PHZBOI\d/Q8fba,e[Td,RBd5XU)#_DL,.R@:7.O]SS^[KPDOCZE?H
C?/CW4)^GE\,ZOEf;AWON\,[2?JT;LDf6Ed_A+G9YO^Mg2-X:A247ZXZCIE>:=WM
/EX0gAd;D;>CdEceEcR>:;JeQdNB:&Y9N+IWKGGMZT\_@7Ve,&K8)V&6DTQDEAb\
(-&ZXf\92V+&gRT&7KB<Z.eIHG&<MYW]SM7+9bS(^CYUZf<A_QY6E3e&;]GP(7)G
b>>GB(\3:aR4+<)L;UB,J/&DD2L>Ve:KYfSaW\CK;Jb/]./J(X2#UBXA7A8OdF>M
KaCcCPZ;JXYgZ,<,5A_DC3Z,HY2AL>&&_X/f6)[K=I0fcb1==6IK/7T-S>(P1[IR
Z,(U_DK@1H><#[B,Y[I9X1EZR3_^PZOJCcA0/Jg@M4+8D8(;g(?)>KE0:,[A[&X]
A-7K3cW5-XR5f\4Gd7P=M.5b>QKIX7KO+,DBPTAYd.PRWcfTJ&3_RP;QGWQ8-29-
D(?e5[GaKC1d8T,Y,DMHI4OEN2<@LLYBXRNT,K^dfG+>J@0JEM\VOa+\;6Y8BSee
.)b4B[(-(>GMNVAg8,YCR[fE]Z[:2+/Hc^-KceW(Vc_2XS0,\C(1caG,QRD#0]7d
aFN9MY##EINBK,LP.7N1)+<OST0]/QT7@OC6dN1JS&-KA(X8b.OcUDdg378TY+ON
@g_]=9@]:#O(AM\B,YQTH1C?K-\<;C.E/2W-++6&-Hea_+5ETN;45CNG15_dVJLM
>9/3B>W@MLGU(-L/dJ1UB6U+<&g5HQ51Za?a_I^2N1Ne7C-g<SK-R;RPZd-X#&YW
W\G,3BO.?07.#1V#\&^)b2OcEF@,Q)[G+#TNLS<@:BVeL/:/Gd_QXBOW;;eYX^E]
:[YXM;C\:,4JKe5B)\S&&8LDJ+>#/M.,@OVYRf_4\M.?]L3P49>KUdYY?66(X9\e
QN[O#@763g8P?KDgL,86O7C]BX/^:g.TRU,V?F[C@SULA<1NUC^#7_Ff-HWSB,?[
8e)YY=NXb<-a^]3OM3P?\81HL)-6=>C;JgI0HNNcf[NaHAJ&SJF0a=XW4[(+N6,;
=<2Q5WD<c;b\3PaVLZZOZI-bU8=?7?:^1#TWVL,AP,W,JK^P\.PV)42UeAIW-8D9
+58=0U&VLTX2X(1bG+&SAMfG6BUQO@5>,EG58;UXSNC&2g7c.UB#0BQHH#=^9OX+
@WaJ9<Gf6dK#Bdd&1[dY-_@;>85)>gFg6?;I[#6Gc&N6Qd@FfK;Z\T^SS3KSd#gM
eFHRd:?JX0)c>1^^0I@+(GMUI>NWeZ\0d<26W4YdAe^?(H8?41_2(,TP_BeL,4][
:&_TPOfD6=+E9BZ,\d><@[G#+Ea36BS&@R<Ag/;Y7d95S9,OdS_;a?N<_O\>d<F7
UW@Z#>aeT4A8Nc<J1eY&+^XF-Z2(]M2(#\0O<WdM\-A-I^:VA(J#Y9b-)1ESM,>6
8dfGI?AK^g5FE=Q&9&V0V.W#eS@YP[]:KR:\31_a&-[851#Y\6ZAIW9Pc2fB8b66
1P>I=8?7d_)^T,(]X.6,/?TGC@?5dUJM:B83PKaKO>?O8@2&5<SF9[9fPQ&;]&RS
g&:>Q/MPE\aI&S4e^/VX68^f&ZM^#IATFgF:C5a[UG)YI2VIR\&4>a+PYX9>aXI1
_21JT-6=RcgIEQeT]add,b7UDO:2da<[14+01//BMC8178dFL,XMZS(8MACIL)T8
T<XbE^2aZWNZ@g(CAY3(AICSX1XUU9K\Lf9d2+>(<8@VEC;R#(gV&>QS9/Z^6=Rc
<25\XEJ2:3A54F8)O7:XL^I2&e5A5[aNN@-C_-]3K^\J(M[/Q54d](LG(0_2.Edg
NZ_=^?eB9M@MP#Q6]2&(Y98_D)/:]PSgWKOeZWCbE2SGWVYaJL>JY6b3Ha>d#J>I
OT_F1REOc<dc0-:O8#2IH0KD\,ea]&<E??9^DKU&-Xc2MIK-MUVI2gc-XFC5+3BW
8>aMe.a2_T;9FcX#)Z+Q5VC.9DN7?YbY(+LW-?.XfD=B8S<cEcgf8GQ#]f+YFQE7
BC@-B^@\Qb_2K<)3:/-c6TXCN]#a]9]INg/?ea>HSH:D&0U);T[.#L(&/g@A-K<A
a7(.L^aWD218[D7Sb3M2g:1gNC-(X-^VWR3L8Z,V1VNDc8T-&9,6-\&=.QJ;G&9G
;J;M@JOV80ESM=c,-:b8\V<6SH(3QN#J:Z6L>Q5(\L\Yadb.I[067K-X8THH#4L+
75dQ]/2KA@N<a7)Z&XceFGGZN3XUR&)0ME]]Ob:ceJYgPV5>@ZO>IU;_dC>_J=A6
S,]BLbbdFTDc.)5+EVJKEITd3WEPV<_MQU([0g=:B8?1JWdH_b@=B[-G(32F4=c(
6aIC?TY@K(=H[T8B=].FS&[OK>H_O&MID7U2W2CK(+H0K9Y0;Yd7=Se]&X8R-&R&
CZfdFGG^V+b-[ANYA1X719Q_&]83YW9)@84JIVNX@JF,4eZ1S>//(b<K4&3R:PH0
/I#&@)WV)6NS,PHcV\&,&(E:1-f54X=A[\H6dD?SN4L=T^@7O7gX-_P96NJAN:@e
ZAOXbV;=6@9:P+0Z,0URg+[:eFD8WV^_cP70b,E4.OZ]7a/Tf;Ya0Y:YHIe:+RW.
701[eW&4Yb(3e:77&XM,X.9OE;=a\Qf:g>GN4]2+F-P=H1/OK\4XMf(#<EOVXLaf
0BZ-a:UW9dU0(Ue)d(]PT,cS0fObP(g\9.;@e[BA3Z6G>VgGB27P3K>O3#8Y-F&O
NJH>a.3]PBDKD2HB4^#R;YHC/UV?BF^O9&#OdL#C-;e-E#f)AgXP1cKLfB5eRDMK
N7=J9PE69U#;e1e#22Y_ENJ;cX(L@NM[e28gE61D)cTbG/<Sf^AO00#>V/C-#?#4
a<+(HJ:V/0&WOQ+8^L?(_B4BFL1J50B7&R;W1d&1X8X+\EBQQS&7V2.H>G0HVdDX
W4:J^&aPI&3SCRaURHDF,b=@0e5-@U-?M7e+Y_H?UGS\(_<)gUCc/\W(]#2_?>RC
)2NYB&fEdJLWa@Lecb8X8^^=dJ3d[5IbH-gT<_XG0,LCJ9AW27?&XX/Q18d(W)2F
325FB]?775IdW/W7CCN;PeSb(Kc@#d1=XbeXAKX?fW&Y)#I<17[[.PD_20Y[eP?c
C9:-PPKZ;8(X]F2C;Y1b,aR<EQaEF^@O\bf?GId9-5.0,HX2W6gXgd+,4P5&Q=<C
/]L\[>[(S,Q)a3&H^KHa^>=AC:d=f0T&Q;YdJP^A9Q=gSY>#+WO0L<S&Q.f.YF+D
P;(aEEK#R,,?W[(D7H5T;Xf@_;[Sac6UTY:)M:VfGY;M]:;0-R.W6]_)72?H_W3+
bAA[IXH<.[;C=LN>ac3GJ>P[75#bSJA_[/]g9.Y<#CT[F5&SccUO>g+-0_accVQZ
O7YC:&XT08R^DDC-.Y)F]g[S5.8\O_\JRQ:\V?f6V]>0F/8ZSY#>V,,:XVgNGLFa
A(W?7I7#geE]4(WCOD^#XEHCIFfA-1fC5>W=RceaQ^F10GC;a\Wg74ZZDL-4)P]e
Zd/7YI(TCY[dTNDLPB[^&X)?]4:?f.4;f374#1a_A&.b^BN;g6e&+O)?:U+LD&K]
CU:efbUAVd4ES58.0Ve<4.cYYD3XU5:7Y2UT,[S3\E4HC>NN80P^Gbb@ESXBdOFg
-I6c36@J:ME3@Be,3(=-BK]dLeHZ+0INaC5>g#RUHf6TgK&IOO.fgX3,<=H1>/U(
c(T^8))MZD_E+=/-L[c5.L>5A0)X\]_ED(6XXF4c#A+dQ5YKN6[;]>-P38g,d;DY
1Y\c7K\dO^U7F4:CZ=->;HM@_5(]#-8Fe.L]/70[53?7fW0_T,7MSc]8\/),#[5H
<Z/(LFF=]M2K\d6c#McUYNbdBNABN_/UPK[O01KN&2+KU0?_KK774..-Y#^M)ZL]
3Xefc#.ea=VB=I?X-:^g4EZc-.=88>71&9(-,DgSa^):C.H5K\eW^\=ObO\^5BCF
PgTT@M#S9<<=C;6K;aQH8GaC;&^?73N<DRgZR-]PV-TW+6d0^V<)=VS:4fG..a-D
UI/;UP?3e1@:T<KR&Va)T\3U3P+c:G6F([?X/fW:C<]RbbX_PW2CT+T6W6_+<QW\
a=&-,I+<K+Qd#=\>D07L<ScHTR)]4OR50)8g@eS<]HXEL[-VFCLc(FB)]KXb?-Mg
b&eOcRN;_[:0;@eU8)+I:M-B+Hg1\P2g.)DK_OQO0B]PfGc2d1@Y\T:>)M^YbKfU
_DWODd-3.fKL-@\&-7&CSYG[8INX3@D(>)(^OH-H4_+,:-8W9CW>+NONX6W)C:+E
K(cDQWe-/-^NaK#^R8Pe?;N=GBCNAA_Y]-90@HD7eI7O)b0;U=;5X.M/D@IIHI:f
dDX&6>ID/8++VPV41GLXg_#4DVZc&A^HI#EK#=KMG5+18,\dF0UZf_GJ^L6Jd6B+
d++b@eA7ec8_LC:DJKbaC]UZ=+LKPGQe>1W.Ug2R.PMC.PRI5dM]X^c44^J5W>7+
[3@^_Eff=:6O>0&cPZ@\G\Z9GE5)]=a^H_(LNB@1&D9M,]XEIGg?JJ+ANYBf;)S?
Hf=JS2PNa[LK(b=EZ=5T>Ee:VfFQS&EE)>cG44M2P0_:/+K(TUDgMT<CX/CQGE1C
D69,&A#F-V&<NQNAX,/B072_@dK5YJ;aeX\N6UBFP3fQ/@AYH&;S566#8Z##&eJA
OS5\@8]SH9Q^NBIX(+A(4I##L==#8UE3/fLfPBe&Q6\E,-WcJBK5:dfU=Na7D6DR
27eB^ZT-eHYd=1cE7=73RbVZ@fAA[8UB3ZcKA3a#\II7;I0]U,-71<?Hb#],+HG^
&O@,&eAD^>BHOS&e0M38YN=Hg3Q>6,7M-O.XQQK)^XJ2(D+91T]3HA?RK0^CeYH:
4.^VSP>Z[+#fYM65RFgO0,_=;HWJTW27&4dN^:VM28>I0>L^PVOVV/c@]5W-cUFa
&Tf+aR[9,3Z1N)/H@?aed\Ve.(-.We3FALM/c4</Q[3^1)36&d-48>=,Y/;>KT(#
QaY]g\cF@1=dA:5E/-?>]8e_#:=H3E;BX1a+C3a]2e=ZabH0QSKJYQI#U<c:F0>X
bV-?3F@)OA8&f@g+Nb?[Z6>Z;#>VVSW0AI);UAYcPXN<gFSX3L=Z92V.3R7CNRH?
K9TEWAZ#@R8185BYJQEAVfYO)=08H-0G&U[[7TPf\:CG)DMBZT1S8?&091E0D=?L
A2.M2W(&Z>V5_SH6P]?+8DLWd\=#+=e,\PEWC]SCV8A</f5(]OO>RDWKXFG?@(.@
/1Z8<eUG3TYVXU7OaS=ZEKZ1b?R(AYdH5adeLGE,Z=G;U\eB[f9c]K8V<>QFf03?
Cc-^XL+NN7QZMLQg+F0ZG@b^LJ-H1_BN<?+b+&/DI=+SZXO+VB0\42[9cgL6YcEU
>,_gS=W^-M3WTg&W>5SHZ7WL=T019McM30f:CY[T?-NI0eQ\2A2a[[@c5#9XV814
e_,?+PgJP<g1<O]._DR#P]Ue#7<G-1NE4TN=K7+ENgCT)_SLfcIUcTZA36GLBfKC
9H+G<d7W.b3fN5]CG5d:B74Rd85e<c?N,>R?:ASUZ65&KTNgg&GB([fIN:?#1?;9
7H3&Ma:G7N-5H.3UJFQ)I8UXN[]?;XR[D5:5T1HRO/Le>f\6<:D;99A0W3#RQZ^^
-M):5MC3D9Cg^KL8a[0DXJ0.QT)\RWWOUZDTQ(CCg0AZN2Q;-.Y\<Q;UEa-fVT^>
B-c&KE3)RRG[F&I3XKc]eQ0/GHgKY6-/U#[-ODF455=C/76A@=O2@]3:EB&,)ATC
)F0&b.M9f:.D6]-Z(eK((f10bKVL]5^Z3+9V/BJDW:C)-[?F/G&LO\X?M3^4QN7V
e1#8?/DFSa@BZJ-&S)K<--->eAW=gX.X[;FT-dXd74ON\@_BfF?Y2[dS)=O<>G3b
3V),.+M04.4\D_D7XJLA-#+B,Vg4N\?.N2dKEcFZ=_I/01ZRc=&9OL+U9T918Y\_
.DH,2VPWfRMMP,e7(OCU/:,5D+N0?KQSG.J67;bC=(2Gg025bN/FdMI\B>=POgS/
S5M?9[#4FKab&F5CIY:Vf4=OF<>\N?6SX:d=LB]\c(QdE=VgGA5]@KCE/?8b78MY
MC\L1\NLd^WH;J6bH>&7)W0UZ^.<]^U?:TNSC(f4?9V>9&_7^V8,3X29Q^Q&a,T8
ALYZ>RP[9=A,]:)4/W[a5,A?&Jb]1b:735+HG<430O.,(/4VcA)e>&>N]&A=@P)g
IAQgXK+_C\)-4Z8I91Y]OKHF\^@[9BgKe4E#@Y_.Z+gV1;_]29WE3=SQ):RdWWPe
#/fPJfN,/e(GTf>)<3<b[LZH>2L-(J_M75\<7J_]1[WUfP]ATGVMGMQLdGWaG=.>
[#Tg8KAC^U#>\WK(WZJT9gCI/A_HDC,I5-(M7[CUCLMg-5/N])TFNC[V/d+3IK:H
f<FOURN,8Z,K1@(?3I6_&8VWJ26-4O8K8]c]MEZTU-;FJ0BKE.QBc_I><;_[R[87
b?B6NR.4UfWGILHNa@=YOPGN7N=LXA>F,.>\7:;3^?T978F\+f?4eDWNQCKdQ<B=
61G.ga5H+,0VYDf)d2eX(=9[1g:b>L-dHMJ#g&Z1g?D]^YFA5=CMD>5MX0QN)QUY
6HEG>+7\VU;-3X]@d<8a#),MV:TM3(BYP@cEC9^68<\2H-ZgRKec=J?(ab/Y&G>D
&8X([&9>60W<-Y-XMJQM<<eD;2W9/>ACSc<g1cQgA@(Q&49&MK3RKZXN_c#0?Z39
@AL6QX@NPN-ZH7U++V,9a#OgI&,L>4C\\fR:5/;C)f2];4>bKXK:7QPLF5\FMaCR
9]+-Y^C5EXN1]bOdZAWK[X(e7^+;K?]Pf<X=RESFFTC<)MP:E;>KQfY9:^8FS4@@
:Z(<[Q=fQgSXG,IJN,[8\3fQ^9S8K;3U:g@/@N/N@MWWfSI#KG^-&FZD17EU&,:J
STVQHVD4TLW5P>8F^T\J(CfM:&S+78@<MKfac&IAc;+HX/bBBMHY5/NE>M<TN<+C
Nc@\e8H9/U.5:2WZYW1-O3-,B:8,@eE=SN2B)6OC&E^\J870bePE[P);EAR:?EXD
HQ:]CA^H_>V6<CN3IR-C?V<XTHJ<1M2B42cgf&&.V+S\E$
`endprotected

`protected
D51@LFVF,0=Z6_G5/\:N.IdXL>2^d#EP^IG@>&9@+9Oc+_\MWE2;/)9,H>-?:dN:
c5c\CgS8Ug.NAZ>=_dHDDIM8<BH2D_26H:QNKZe?K&?KBWD1>#=.MS4;9+HN?X0\
gL7T[cNG4,E@,BM/b@FZ>cA/HU<T^a])W@PUAK\g#1;+1SYFOSBN=]4;M$
`endprotected

//vcs_lic_vip_protect
  `protected
+.PV+b95b\M@MH?PW_O1:3+9VMARU3Jc=7#g>N[Mf_5g6H+P:.]X)(NfU3EMc<PO
DZ6SM-R?0c>U6.>+^=&fc2ZdD<7(#KSg#eHZA+Yad/2@SQ?-2;T[>-?aD\_..RYU
\5&;>-d2^4\H7JEK7)5.U5SR>@#?#G&]@+V9df:+dXLd+K=AX2JR,V94)P?B:fP#
038aS&4_(SW\M87(2JUA/Cg)TO]>afbU7ES<A-FFDZ_2P4Vg]_TA9Z&S&JDH25Hf
Y4Kf8R1e8;(Y6;F/?gMc]-5&^g)C8>ZKIH0OG11T(Tg\9W7QD[7H>>fW/.aX)P;f
dV31RgR.4_U1;#_Hg(4bTH[9[U+\HS=-]dgPWGb@VX#5?/Q2O>PHc)O8W&,#OK&^
5PC-bWPbTaS;7NYP>:EcgBO>[0AcSc6e]?e=BPGORQQ73\e\cGB.5TK,-^ARZY3f
ABd5T=EFH7G41,BVFH@99R77-gYY5KK):YXK7c;)#V7?;5214IGcO08VIN+0A)1.
FS,-aISAA(-Q#77#,D?5C/Q+O2PF5/,?L-S_/N^f4IZD8_bfeg0aT&V#F?2TOKJ^
,dH1Rf@]PL09c>9@@ZaU<FX4[[:e4R/[cY7(Tc6ZZ_0S7@83g=e^J\&a.4aAI.B/
.<W-:RU9.\E=_F5]59,W05&X/FQ=+g<L_5XG?#>^VFK/S7)8;>7Q13f9.;+?\Qc3
(#]]T/.38b-.[0VR.L9F,6(OebSf+A1JgK1T1gVOea(E8DEV295E#8;27O5bcH-M
#7P\ZI>(.)?0UXYUgg#];F/df2HB,KFJ]Y(e1)JTEa8fbL2eV\-?(Pd_^L=+V.J\
.3DNG_=^-.\a_BQO]?#K(ceZ96eU18DQ5=C,e?B4^L9&<GFZ1ULf<M,\+@>=K:[6
SPT.8I;W]Eb4RCMg7RY#cT7c79@G><UZ(JPb+Q]2A\eM-DX9]QYIN:+f\Z1JaO#,
T]^O1\_S,<EO@JE@:9MP]+gTafg3d;OEbeOW2?egQVAV[;ER7:@XKF>_<P/+U>W+
YP2Z]bEfGgWLR]ERaOIcfHC;ZH;3bNLKKF#X,Dc;2/M7=AZ:#M0[2_g2)NO:1Cca
&fTU0_Z[^A>4/Q0CRWeLeA4QLS\OTTCJLcQWGIb/P:.T)afE3I)4D.g^)W8+GS26
>&9^\0[8GJ&>7Cc(a0ACSFXaIG,eWSW2:fZ+P+8MWZ/53,?.T[f[<?F77C_3)c?O
e12#ZEcUTF#[d(:B]<+G@Z7ZGYeH,4;2_EHN7S&>7\NbJdIC+YJcI[]FP+UY:T#9
NPR-P2Nf,E9Z@HfL.dL@NSR0<.SYA&>d:8d&[YFPHV+3<K<Wg_UU?#[YVSBMAC@A
Rfc_N:+[8Q,959^H)eS6\JSXb<FID&)MOA/#4G.6<17/15>0<Y(TD3:dgL\g9afK
_F/YYc2]6)1&-;@Y/WZ<7d6aND3KRD],/&ER/I=ZP+GP.BZ-AH&L:^GKd3X1/Z1Z
LWCTGL6S0LWI&65</JU-aPC:[7G+J680(R?/V_3BY^Oc@FI=V_]&<E#8P<=25deb
4T0V_^_JVA\7J?Je:ITNAU4+e/8)N;#:d=gc(3ZNc(fOg6Gca?ggFC6>=2E<-g>b
\\7IL_cC:&,f#cN7IZa=H9W>+NI498a:5Qc)7+/Ld^6>aFSO@;X6(QdBNfeDMe6Y
:/\;_1AA55da))CYI6MWVR1Jf#UdW2,61RZ^P,X>^Le#f_SRNTVC6?fKf1d9H#L9
I?XT&\.QKQ?(LKe]?<2RMN&&QUQ[51W_&UH,XcI/bf,R:e]28SZ&KNNP[/#g8_4B
fCcW6G>/A\)/H);K:^f:#&@::TC?WT?]Z7:(5J4[SQbFLB79R<\\LXbSVR,KTNe;
>_O<IT3D&.]c_>?69eZ5Y@;Z08VU]G]UX/@B7>2-<SX<c17S^UX#-E_a^T786P1_
c-LS(@\\LTQ^WgSb]1e&NB)Q5J^:7;a\@J>M]^-a24EZKHJd/<&.NJLHCEX+Wf2E
CXINOHX]9Z=)>QRUOL45g<HW:3Z#ZPZ=f#[,-09UIZ@QW\5+.Te4UGZ0eL-5;EA]
4P(dUN6?N#2Z:N4R]Oda-1--\SF\_VN)WLWc]\201\A7<8UXLYW^H+_+HIV^g)(W
1>[^+W3?T,OcMLOE5&10\DTY@CFC&IDf)PeE1+9JFa#SM:A-BXV>K2)^?(EJM02,
aS?_L5E][.MBJNDWH]E#,dU_C)-e;a2+\RgL.aDOA\N1KF-#dG7e9FWM82,EZPU;
e7(GGa>4,I@bD8-7UU-a;=WZAWb(/9RBB#NfV6+-XHfM^<,^3JeRGQ3+Z33I)=T2
Q\Y(?<83_#];-9Zb9##9W9\K\W4A)=+gV1U]Z]U><a(7+HG6,_&89FX^7J48_NII
V.[6)74NEMgY/8-.,A)>VbCE-a\#<#>W\.)QEL<aMA;f?(_d_30NXLbU]fIeN0(7
I@Rc&Zbb2bQ^[H.N?,9Gb=Z;2fN](1S_b/W_5^f=HH#aO)]36:H^aGMB3ScP)[G=
#^V/5a)8@a82[+KO(-C8NcN06PKQ7-dA6g=Z^b-?E<UPe#Z3E7(AU<;.MU1E#RPU
X-]6XV3P+@KB6W?c[IGG1VZPNf1<H?.B34fV8e<gB<.9dRPC[0SN8X(aW5M&1a1?
O]A5/:T+9?BW-Ca[QTZ=X9U:e6:gb-W:L^ZC3cc\A-Y4cEGK=+gf<4QG3Og;NgXS
e]8^]JJG9VdXgSFE;I=-#\1@_,CN.<O+ZQg+JI+3(U):M#SJ]:7/bL_a5aUHb0N;
Y5(;(S8VG/=)V]bNZ;)B\5V\LA(\-1Z,TFOM\M+1Ac_V&&WBV3bUZI7aY_dc:G?Q
BPBF4??P6.:FB@JfUM3:1+N)g4#@RI>ZHGd-M4MRGV-0Sg^.)TS()1A66S]4FLTc
;DAIJX42@a>9\O\J6,g9&If>>,\.KI5=-Edd90=,+HI?NYaN-070cSSdeTa-C.Aa
YCdc<1&K0/A3AcE\\I>QYT7T1da)W-f7bJ6_9^aIBbeHaJL6O0GRQC>.4VfUb&[1
_9TSO9LR-I:?1eTYNXaZM5OQFRQ&H[FS<R)>-P5-ZZd2Y7,]3c7]798\@>2]IW.Z
_7E>ZTa=>3Q8)T&BU=9#9@W]4[23+B9=HNI=W8L215@9A64=5)MB\8,>f2O.@^NX
bV[>4g8LW-TW,1^+YYV#C0ba-N>8gH4\O>992O9>cRSYdJAZHdT^2HOMa\VWcDWH
QcN?[_Z8)EP)R[RK@(57D#U?XaLW?[MB880[.HYYE&L1Z>;MYG/eH>:D>M_#?&+M
4:_W;(c:=X)6Q5[6LaOC>5+?Z9LbcUM3YIJN4.V<]/,M-fS9cW73NU=7VEF^9eVQ
U5d,YO=(N3PHEd7?3FDEHT4P=[?95FR>-15;[6e9T-TcE;bI][^K?#&:L>&=S5)D
L\e#BI<aHQd?MI84TfMU.(H[WR_EI<f[+IT57F-#>YLg/B^[A>:01@#QWRH<d#=7
ANMIWV9cP5;D(5GC/fV+#H:=VIGbXP2SIOSZL(\05b(?Mg@0TNc.0RW7Z>FeF:(/
gWJC/DG453W,XO46d7eO#B/=c>3AW<865LD8P:c81_>OS10e((:3^>b7XYUBV-BR
LR7.B>GYC=HV#fYH\(PAL\.C:0YZZVIU466gBGQISZdV3LP)8<C]Od6/GfW#E\GS
\37)&NXL_<5&&[]]E9)ZTBJ7ZY>7?HQUd3:[Q+?=DC@cBM7,EO&Z3YXBDO^+STd\
XaVU1:1L+\f@#[1U[]<a05T6D#cRBdKa=P6(WX_L/>T=D<+;HL80,C1W[JH3WV5f
Zg_]1]EW=;),FNda?O0[3&Q8@6J[#Me)KWH@dPPS.2c/](LJ<7B6.8[W@X9&^+A[
IfaP-+bb6CE/:ABFOW4QREgNR^/722#X@50DH2>W93XVI7,>5SA/X-PZ.9fd/&G?
0ZXSQ-H&8LPWC2K\cA22N>Fb61/F#QFEW[3SgX)8];#Gb-@K9gV^e(0[AUG?4[f=
1fg])9LB4S3_F.U84ZY&.FE@ZPE86MLaQN3&(/8\^F3#]VfbQX6@TLCSWXK&6ZHU
F\56LbH;A_79#63FbfDM68RU).M)M^PH,=30RHMW#+W4g@G_MDDb_&4L)9_ZO3cV
Pg2HLU89caFdcOI6+KVUeE9E+RY9_GCgE#\X2((DN4_LaTMEWLYFW&[T>Q@<JU::
,VdA.>B-396P<EM5_]O^L^&BD3^6>@R:HI:P9<7fV8@,-&\+,UdS>56NbZW(,A-0
86Q#DK&7gcNc#@5(VK\GD(ZdZ>g0aY8QbMIH,CQ58)dO:Y]UZE\SC6]IfT&2&3cP
Ge>Z@EZ9=PMbefga8I1</GBZ/;@T+G-N)E\.#fEB=NRC(a\MFM@F[2(.eD:7:/5g
V6Q54(FgC?4gZB4Z7/@2GFeIK8.aY(^+1dB[;;S0KVIM>2LLV7>S,[c;/;CM7+d=
cgJEM27]\GCNE<5Y,g=2[J=ZK^(.K[5bd+KEHETYJ]>+B]#JF]0WQ.[@NdO7\#?H
\H^23]LU2LT,E5gIRGd.9[L_Nd&23V+P9L9SS]c+=NDcb);cXHTFe>+P3Z\0BPb?
&?gX@M#a_TAeQ4<+d&>X1fP9Ca4QW.=J818bI>#<2gE]3LL.]D<8M4C-]JTL@P3R
MdM1H@U5-Q)@B&1P4LWK]JUXI/ZcWCG.ZA(;D#\DJ9)UL5Cg>:QeEBBHFL7NA\P\
Efg+=55UfQ2IY[02_W+a.K;TCR3VMO-gA(D94B>65^6W<)VE-T+g#01:LA=0d_GB
(T4,3@:HHR>^/V.GDTZfY,,LHQ7]AH]LY+755B>J\gXZ(0#4-6OZ(\I]TJN^a]S<
DDW;L#Z@&=D.a?11fK@eFJO2&,&O[#QLO.Y1+^2K92(HDZbdWdK=\[@/-^,XZ4K4
^57G86+D^#2_JD<L37g5L4(D@>^PPfR3>3#SBY,VXK9ESLA]QF+]LHMZHF9H+M=(
^O,Q@2956dgOY5VA(4[W8/#;gS?>D@Aa9ARFJN]BGG]+[6Y5^DZ+=KQD?>4@R2_@
GCaFe+=fHH;Xe#&A]=MeE@fB.LX)@(0_)a=^7W3V,SO&(+C;G3g_Vd8eX1&X#V?a
]G(L3X.XK<OIf9OJ]5\a/G1TNfXBRS&d6T,=9Pe#e(Y2G0[RdM=Q6Y]P;IHJ@P=:
bPUKGJb=DfRfRgI_Q7?V3BV;NfB]]f6UR&K^)6?]?.5edYf,?De,&,O\@Cf2VPX7
&.SQ_:+#1P&MU\CAE\S[MX7cP(NC7YJ@@UK,2U0CDD>G@ZA(A>-aJN)7@5/7X-H0
0/fa>&aaVECQ0SM)c[W;.[b7a8NDYE=+f8N(PZRSH(WbAc]=4eE-J(KEWf(MFK30
eTGMS79.H;Q@G,3XMGaS>XQ7Gf>B0^28Q:PB.031453WVagT^_7dAb,\TdQ#_,/.
I87e/[1U?WPP:-e]6+;(cdg3:F0)81\/\A\P9HIP+LGK7Z9.,E2ZT/E;[NLO_Q_A
/R9CBO;e#VM6Z:#/(#aE/F-GB@9[M(E,[)O5K7:T2A]92SbAN&;VD3B37QOeF(+]
Q&ZJ==[2.U2\>RGcC.Ya1OS6;/Z8WE)UKN<]:P<0#dRUMLU&?f>S>bJ[M?Y74+=_
?=.eBeBgKKJa>TOa4X0&7/(_N@.F0DIX:7I5b#(J43Ba53N,X\Y),VRK6?<Hb?EU
^+^edFbe\/Q(T5c;#P)[U=]<5\4d1U)(N7RN:1Y7LC,X(+BcIZCEP0daN17R-NP:
2;e4BUU8C?[1TSZ_a+D?&T^3\ZaVe1H&MPeTITabS@B+2]KYG1E\W:@KcO959?#Q
<RVY\/KF&+d4NU-=FIU;682D@Z1W7ZG+c0>\L;Jb8eT;@?K&(OSdEVUV;NF(P?GC
NIZ-3UK?Y(F9:27[\4c]f(b+Z4RTY1=B98b&W(@e\J+dB[cg&B/BYORA^+ZE1J_:
/H+S&fPT4\0/1NVSB]K-ge:YQ.&8?bA&c[F9\LQ]8)E1<J6JAR/A9,:.)US0P.SD
PSEc1?;dW5HbQLYQ\&\c9B7-fN]C;->W).<8FL#^1]D.]H=IM^VBMES6>F/&bIK7
\aM+@MMgF)[-03AB#Q_M@=?g<<c#FIT.NK4WORH;e&KS@CPP(?&NB1NKF?_B<FW7
H5B3df7g+YPH>.#.;8c5f?SbB&V<K5e^.9[+:52V._M/2?OJ4DU6#@D3,QLab>0J
V5WOZST>\55A3,O]c(VX(?[/Y22.1:;6OJ)\@E>>.4F]><\1Pg3R3AM):60.]aE]
b\MOd-+_K@0IU0-_CR-^<>Q[)d60c?gR]V-<3KCLV1__]7#0+XD.&->Bg+#_JNY9
HS])^f0Re^c,-1bE9<=eFR39@7Z>.X13U5Z^3O4I=?<\1=(T)_>3F:GQ<A@/eB60
bD);cW(/f8^1CPPYUKOa[RS?^W7?QTaK77<+_D=.RDIF_]b4A+3N2BK;GB.<g0B4
=dG-LI&)VBFWJY)58<(X2LOKd?5/?Y;0L(##SVT,;(XBEYU^aA1NR0-[M>>]<<d4
Ec1DDZbU5,_K)Vb2<eg/7IZTIQO]_DCM^ec&(bWSR]Ae?R5S4dRH@0E,-aPTc^Z(
7f^Z>1d;A64f(@DK\DdG&8?8Jc9bag=\+.d?0XF@VW;]PfI&^,eM_KP+8CC6243<
&1a[A/R>&1Zd2M+ID&Eegc3;]7-Z+>R=HHTVa@^_B]:DRXd.2ca;9a3ZEZ)B.a;=
c<?B2F(&OSJP=R>ZIJLI+Y(\413^ZYG+H,YD3LV,WC?Y3WOU[GeebLI)2TP9[ZH5
00XN]B;5V8^&A]PYLe_,SXH#]X8&G9d#d8UB7R@;YO6MJbH#G3-=P6-NAQbW=.E)
H)aOSKOF@6:Z6fdW^-16FD[]5;+50Sd(?:Adf7S?G8XJZGOP(74FCeLIb^;_=(e>
QUMcH_Z#/-NObI.f7H22cgQGI\]>94::H@Q6_J6Z/7Y>HHT4c^QD00NND?dRdaBS
S>JSL,[dH2ROJEPB^V]gF-;AK9:ZS(:<9/[H=#P,A;KM9gd7B#g8f>;g269eLC79
d[/WMGE-]&O/Q&);JdC?UP5;,b]Y,ZRS.dK&FFXS<SaIP(gF72+(db/1SQ[HdHZ\
,H,II#2M)WO^RLME5[Ee0U>Od<6Lb3@PGB-C2Ic.TOG5X[-MHAe(K0g0A6@/;,7a
G1DY.8/:91gWb56baLTA.K:X],NJf(?+4I3S#,?Q?7XX=R89KXWW]?8DIV7HY++)
Ie&Y69dD2gD3FXf\UKG]9:G.#M?EX:A\]0&cd5)U_M\3^4</X(HPPgJ-6W)Vf[,@
HTYT<+3gB2<4_\X_H4DM[[1[:Af6fBeLUe26CE-RUgEa>[+F81KN#RVR(C>4F[g9
]7J6YeF&[fYR+R+=g@6<E+g9=/]NWg7:^Y1=F?[4Pa99XIFMA,5cY+47\S@DPA#<
IYaRL.BGg[S)^WVD&\:+/53cCVO2(3VP,2W8/SZOVSDg^7APSH]52TOcMRS-gF3a
(IGEI/OYUdVE_?fWP11_daIZI-_O@>N2;7gW31(0A?;+5.KaI_APV-CD\?Q9^P;F
a3.MECX5[gACRY_.5_K1AbV^SUM93/QeUCG5[M9?bPT;Nc-E9O7f<[[Bc]SM-YM/
O](B@O7<UH3TWb7BY=_FS@8bEIW#Q&YXg0]09\MD@MeP_<g7KCVQ#BQCY5=04dPO
5D6dZGIaf#965X_dCdDgJQ:6:H8S+G.,6E1(MY@IZ7a4ddK+0RRb\MEYUK+9IZcZ
P(GO<W2Ja26CRYGH5bCXdE+E;TM?GL^O>Be?1XL)KfVN@]BFc-4@ZAGQ\+aMHQVH
8IVR?ELY^ZYZCEQ5[5XE@^NEE?f3<G091QDddb11UQ781>UF(dO]-)96e,>2eF-5
E7=)_HWXa2NQ]0_:.<WM\)RD3H18)Af@5>,0UCZT;;&#&[3DGD>F0SE:)4J_D836
f.O#a18>(5VX?UUBH6YFP6]=gZNX&E\gf+,^#NLF)c^R5e:=C3+L+H5),Pec?K18
-WS_7#1>E=;ITe?fJS9cDW1<O&6C->^CJ^4Je6L-]):d8Bb#D9\[T093_NFSQ75#
::SHd#3YQX^RBc;6bK+V&U&\Y[12]#ZbN4Od19ZR47)g5EZ+UGRK()^/YE3;dV1H
2gMK,MMRU\b:HO:;Z;B]I]B1<bLS)IO-;2)(8;;WB[<JT)Sb5dLb#b2,^=[?;,;g
20RE@_3KfI^TES[3__SPBdYP0fXMJ\18;GC7#TRD7C7PYE>D-6DE7FZ6f0cVXK75
/7N#S(E@/J[=_1(FcdV5KaQQV?@b=bMQMYaCJA7d68Y+fON:8?d06C/)(@_1cX.\
TW.5PaR:1&R^@?cWf_Y7d_^>N<HK#:8]=c_[N&2EO7X8HA9gA4KU+@_dLTFV4>3N
#OSOF2\W5faX0][f9MZ(-5abQ<WY<USX7S[?F4?S&DV+D+PD;X77<CK-KV-)K2XV
IW;VgO+]a:ZCg.-=SAZ74JB>HP#K+?6E(V^@.YD@@,dZ3I)\C<XV>[:63)1FC41#
I=ST8BRP4Hf9[J3<\8.BUIf;&@?E/gOVc/E@c[1MMcE2UM&G1,P7fE7gJW/1&.XR
:f&fd-0,6WgSCK6B?E4f@6Z+P.K@MB3Ca)87CR9INSKNU@P@DABT1^2R33Y\>].0
VIECW0/.gEZ#M#]0Y:fWQ(;<JHc(EPI0d@RC^N_P09ZACI8L1W@g4JPIDN+TNW)[
C-B9QTDKZd0OceMa8aD18Q4SS>>G2V>]0YB>bd:B&0=aa.bV098[dI\0bLD)94FV
^VREG4B9G+e4NF3Jd5]V)+;F>UMebS:3TT,2YC<XLBMHb[BY#bFTUNCR?_G=W_RM
QN2\>];:51XS_]TSZa?eDV3M>.W_-F>/>8+E:G.FSXgf@+.a8WM.a30Z]=g>:NRS
M8,Mb+YV;VXUVTSZPe[6eWEM8,=@J2QF&NNA5]]^.S):,(P5F>8U\UTY>116:3IH
<86BWdBJc#,R@REB4_WXMFd@=;K?-Y1L5SN,^c5C2T1V.Q.[@FL8[J1^MC@@bI#B
NC0>#b9=E4TGZY+Bg,Q.&&L<2[\;,c/5EIL.,VD9JY>6]b[QCeVYA_/WW40;>c\&
&@4^QH[G-I@;6\\4J#<;S.O9^^AN9?N:3@Z0AI7a)_ZQ^Q1f?4ZXO(3&<75WY<SQ
61/(,N?J&RLU/2,dOR(IS8QGEJEZ,_2HFS84-^YgK(XVAfKU#PfJ533d0>R<15LU
A:4+<@:L5_DLPeE4SWC+QC.JKfA.[2?HA&/8@Q3373A?PBFKD=A]8C2@,MBS^DCH
^H[b]WCT=RSKgR.?F2LP(T65C6QQVE(L>:C?NdDFM1E&VG6Y1D7J;eD#>Ug#FBT6Q$
`endprotected

`protected
_g>#QL-V.2^BJ144PU+R,5=QNGIV9/+<b-6XUQI@,9V[HEC-(34P.)OV&A=X8+I.
f^(+4CXP-S@2XcJI2.22T574VReVR2/gMA_R.O&Q3<-D).J)16=6DYb\Z6]RV,C<S$
`endprotected

//vcs_lic_vip_protect
  `protected
&ZE+6>]C7Pc]OD\?X\,EMA<YU=.7,#;^=MS23>UQ-Dcg9c\>E-+A1(#S+_TVE;-+
dA[@9X]=>MNaHE;FL_ULJ2RI,,-L>2[ZgMUdH)d&MeBO6N1I,4[F72M,VZ8T_E1G
@gT/M;0b?8,e2OFXgJ-W^TIY:6@N3(3WHcdeeVO@Qg#+/7?@ZV^;C5gNgTC;VBNE
MK4HS0:5S&HW;;A+Ice+f2Vg)ZR..24PBUKUT&c##S58,)WIT=(\B84/YK:-2=E+
XB7[YQ:LP[.5d\dXJ[+P(A&),DIO58^fMg+2J@e@:]T<8_6.R_U5Ga=A5CRgQY1(
f-K?1;dSH>d3ANd[9d],P4:E:I?[N5O3,9Y31H-CM[,^;>HD<MU\(=b815495R8(
F;\Kg52RUY)a;d^A>Da[=M]aA24P/,90c@aeK_,J^)J5b,:E&+JS^6F^(Df:f>eg
,B<D&B79P(:F+JJ[6g^R0fCKOZcIZd;:DU@P/Ua99FYYSM,<QM0F&fJ[=0?.?=70
B3eP\SbAZ^TF0^H,J)7(OKAYe4aLPZUX[_E0R>-,IR4?@e63T;[1>3KX.XH]fEVa
8N+NDB-R?;T\A#+c_V6Y0V;Hf;cdb^39AXR+D3b>SC_8SXHH@3BbbNMJAGUGAIP+
&@J0V&[AfM]<d8/=.A\9Hdd5,D+H[6F:5B<:b-(,.X#F_3HCO5X)])Bfd>H(U(M[
9G&aGCLNQUZWJT(H?Z6=f(87MTaU;+93=?6g.J^/WFO:[+@PN9LUWgX478Q;N.R7
g[F/^f^AX\)86\(bB@8Q5DfRHGf=c^6QX2cAWNb9X,G[f9dQBMHXCO+K&0&?4VGJ
LG]g0/f;e=[EAUcKE:+#TKPgQdED9/6Zc#,+O14?]A&W8NC>S26:V#&UCHOQ8Nc6
6&4]RWRYK,USc572aA<[/Kda4?;KG0A/N[PaRb6B)/CC_.6ad>N#I;L_Ob1#O<CH
KUJ/=?>5C4SAE6:6WI]BC^N7,B6I/_TEY2ZeF3?/\W;Z[d#BDN0&SXW0+Ng0ZJa+
eB3RWDFPf&:L;H9f^B><F[S^YAQSKd,M46HTVf]0-Q;TFcEQKW]9IR\_=3M=(C-0
-3_;BZD_9C4]-8;J9M2PYV/(d#][>ZMJMEO:V^A7Y_Q[>Z@5];B?a#f/3Q-BZ.;^
8\]dVMKNDD2=[#4;;e^e?<EN@8SA?8S>F6[KC(<&fPHA(,3?FGB(--EX&U@-fO__
A,P5XB[Da=4]]A\Q35fed9?/J7)>2XHQ]RS#Mf:1G@,HZ0_LPFPO/ZUMNW3[EW]_
HO6R0V51X7cC8?/VYOA2=PCe0HB>D:Z9)=2S#F,HOLO+)I4FQNdOHLd7V>1-,_W(
0QMDc;RYJK[OBAG3N5EJ)Ff\X4@BF.bKMD3+S5]L>L:?[4cMB:Fgf_b-Me_=X2&\
M&gP.>>^Vc<_e^L:H/+]9XQ9N9/+PHJ4-L+,Eg>#\#19QXF-B&_HRPY_[XQ&Ye8Q
fg>]Q2QW&4)Ef+TIJH<64:cTSf:3\DSL)\IB:5+f;184H#AP]5@JeB0:8XLWY4;,
YU/>8@a;f]85GXER]=O=&NHSWO;5d:1]_@X??8H(b9@78(g.fKMOLY6^F5/6HH9C
YBXZ_ba@3&5K.,edFFP>@E:3K1_R.a_5N4-&]+OKL3S5dC,D83bUMEbTA(HX(JY;
VNL6SEID+4fL[fg0d9<]GGWSN6^<F6OcTB#VB<8]8U]-NcG&3R[&9JGXQ@dE#XPD
e6F?Y?@L6@,B;6USc,Ng:<S<QBJ0?O0/-,X_68MG^bKMY_a.HcJ;.#eEa:TW2[4Y
71H&YL+FE(aY\Q?KD[HJ4&=256C#>,-XRW3AW@X28d6Z.gN_8Q#.O>]9Wb/(TZe7
D5ZUaTQ5>FVeZ)F+=CAQOBR(,8BVPK&M&8b,d=Z+>8KKZOZ&Ng0_6M:JX6OCf)@d
P#2Z0Oag?B<f<7G3+dcTM-Oed)5FU2>6JaLDT9W?[aTTY[T8+4EO8XW:]N81;&&:
Z@K^6;+-O271g>YK;M[DLB59-U[E]54E>/HPAJFBUD5/N<3I,W\S]a4YD\dID(L1
)c.Zf:;Z\+8M&Xb7I;a<LQcGV\HKa_X^=FKaYEECg.8eF,\2\HH(2UCQJ6&ROaEd
A[]E:7?-E8Rc6MEW-[^83LF/1X]MYT0#>>&:0K],g+6[ADCB4(_U.TfM+dS&+[4+
QIK2\UQ0aC2K6#K83&(YAMU^UXV>5CT05#1>@UQ(;.f5C+0X]XGJA]U7V8A=H[G+
AbK@O&IVcA_6ZZ6gSL9V>\F?+g_e87Q=dN,dBF(AV.2Q4VQF)NH^\L7LB4f:<JIA
WRXE#<c:^PH_>@PUS-N?g@+1Tf:XSg;#J.C\/>[AW]Zg]MMFaK[AA];BeBP7K,BU
CI;J=^R</#;);P;M#H8,VG>6H^I@Y#,N4eZ46>8[bE:7Q06(XWV/#6?6B^5M474.
G>X8cB\MOfDUU<_Yd_#(<(ICJ8>&V&TX<8fa(</fT;A>(#Q\E/LA&FI&3L&HAS:I
8.@RgH[ZT])MegHS[\4T;+[EZF/H:-7X/VF[WDe==cM1H&bQ)G\g[JO4&::.?#(E
Q8<E:YL9f_Y+0XMbH?]U93KM6+L5H2.Vg>;R46N1=:Ra;G,QXM4(<+XIdKKZ9a^Y
<<J=R6&/49<?&MP:[T]C,bE&d;I0&cX<=,MI.GN8QZ/b?A9<97L.@SF=RU_,K7&Z
^]BBbXedgDR5XDa)WE;/&35IV#ED2+G)_bSaTRN0gHd9cI1LDPGUBS:IPZG-0O:L
6-]N];L\:Zc.XL\O2(0V0OP46-C]9f6#\W+07[\eLD0T3M:_A+N9M86?_,bJcMCN
C<dIT?3KLNTQ5CZ=c+aV;ObI?1:IN/QG^-Y7TH-TfDc:4;4VR,T/7(G,;N-Uc^+a
M7E.3<5A>IT9b#S79R)Mc@-CT=FV>[@Hd#]E0GaZ8CB;P6^/.AAJ^\6_5a^A7Na=
/GTY;3#[XRYVfXcS#I7G<WRcW7;5F1]0egG1O[>I<C>3d17AQ4g.U4JG<&^W<GfD
B7UJH<<F4VaA;gfA66_#(V9]=Sc_dc6Y5,e_GPP9W8X#J)85<+NULBc[;C\925#=
U=7A[-JRV]6dQ99#B2MAKb&=V634J>4IMHXEX.P+=G.^4NKF7Q)Y(#](-eC.>^N[
SKF>E&Q./LUAU(=E?3e=EAV4<;0[H@:2EE&L?/e3ZOe[@;Ug(Z9.X+2PcFFEK>:H
aS#Q:2Pb5P=7Y.Ca7eL&e0DC1#<PZL/f9-.?SAe>[(DeaQcE&K(Y#PSLIF2MNJ77
PYcC^=<#a&3b_Y-R0CX&6Ta92g=8-=;#>d&^O12SD+\\&ZU#B0BPeedWKJ)Adf;>
3?g-c9-5Wc\AT>(gD3[W8/OJ<:e0V7aNYP-bIAQT/YP^/S[<1(cX76Je>6=]1c.Y
D@1).;3/,ZTc]eBG)NDH-f<BK&^(Jb/2N4U[,I3IeGJ7GU<.b7(MUPX;:#9O+M3T
D6-a><DU53RP/O@Z7>VCJWEGBe4H8S&^-D2@UVf:SgSJJac(;5YZKQW6^HcIM5[G
6IHB>KEZ@C:\J3B\>B\,UO;X(K3N=FBI@9bK&C<cI&@>A8YJ\9]9_GBgcU>8I5=[
/-;_5(OF(CW+.0A]P17WW:Bd_7A,CL@\cG;D(NG_E^a5BRdgZ&g\eDJ#7c]#9<()
>BDb;=PRce.]OfR01:YQ@)H5SL0LF_Zd=(Tb.S;_dcJQ&6&2M];(;MF4>b#CXJB^
^\?V/<\\:b[#=:eCfW<KGb6#.6a_43((5#fNY_]2Z\LT>;aXYeb2O\:9-\PN@1_?
)d3@(VKf26X14]S(J&MRJS-Y85[N._@S]?AY<VEJQWc/cDgZeFT8VCYR);V#g5T@
+g5eR=]c=DVBdb3>W=V_K+1CeLJ[N@MXcQPP_YM8)9PM2@9R1dHA0HdL&IgI^UUD
+L)aHDNb#Ud.FJ3CDBYEAV(];(f;^.O:2)^D.D[eIVO+(5EQd38fbc@@C5_G3;Dc
-(@5a+T;@VJV,7(BQP5eGC](bCMHgg/gdVXX9e[3G.VSM7DF-DL-eY.E0>\M2_3=
3:X3<PR4+OI-73SC2,E&^<E^GR3)3B3d[1.T,_P.ZNXaPM,A90H)E/b<948-(TU@
[J(Q/4^/-]f;MT&Q<+ZZC#22d3X(N[^HMYF#U3XQ:00#RZP@UWP+A4<=-gVLG+;W
E5@XZVK/6[<^ZZYPfBUOA3c+]G;OLf:D?GdAXC-BY?<_SY7IB/O+/KDd]eUbdf]>
Z,;R@20LC@E]K6?ReXg]N^-,IL?<4Wc4?XHafB+e22bG[B.&R0.^_<4d=)T6ff9f
cBc);d53846<PS,]FP?D^UTcJX\.Vd/T3g;07OB972<MgS)GSGJ=G\37Q;,R/^NN
^d^_?ebRW&</eO)>4I&3gPE[6=a:V:U_b&2^SW,8GT9/Ba1/_A)5ON)+1F]1L6Q7
\6-6P\CH>M2g-DE6P96TZ_PFbNMY;gU/?Y=,FB1L?EagYb#.TR?S+OBKE>B#DCa3
f[#7,/Eb60BHYPXY=aeAG.dOTX/Va5K1]-58a0YId\G/ZJ>9T:K<AIE.:UR5+,=C
V++4G(ZGdWC<EUd3+4K@#5LbJ.7b#X354IcD29<d))#d8C,JN1Pg(6X>TaAeI[Xe
MRY-._LA0+\/(G_0-C<5We-<[cM[/KCA:^<W=3_T8RAYMXgIX2,T):M_a:N8J<,:
4d46,_].If2)6XVVBf.695d#MR4T5;cBgYPQ3-258##??2.5UV[E.[dbM5c2cR(B
@e5<?=#SCICe1JH=5U4^A8IF]K#:TYeHed?e@F^5\6I9&8;XQ+.L\JN?,0,d6F4I
E(&bU6@bbU^[FRV?e<E#R<I;=c8SfU@OdNQ]b]&].f#bX0_cW\V/1T1#[5M,eR:E
a4F=+DD+cV^)5Db#SQb2E(IKPE.?_&3GW9-d@LDOc08D(4-G,>8,c;MJ9:\<]W=5
KEY8U?;YYY?OC]9ZFO.3<^4B&ZYM6d1VEADM#LPXLS6E@2IWO-L,Z[5[NNQ=1O>)
ebB1&HND<([NBKY3BNZ-XZ5OcS)1B0QQAEg_>c2DQ<OI+40M.IV84IV&1cBFEYI7
-+M_C.^90/TDfYJ]=G@;H&0eGCG:dEQ7D&[,(:>P1(eQY^5ZcA9)TY;#1dO-ORB5
G2fD8QHUGFe//FW]6#^N4+dBN/2QFb3SR>b=.ROLcK8?\gT-cWS;J+T3gG37I78Y
KK#D\_:gbc3C#BS35V.geYU[Y^DZ2(SYR_fa@eDM,f,H#;0[SX(-#OH[R)SNZ=LL
c>70>S0fK^DAbN\dB>/@Z_aYQLU?9P(6>FHd1eC7+4[2d1:[]g\,]7L&b;D4daVI
]:7S4<<G,/EI?]J]a3D94+1;D)OL(6S/_e(G_FRcZ,OR&D;d(AVePMJ?YL3A\aBa
B[O;IK9_SHG+SRA/Y,QdeddffJMB\.<-1NdY&Z?K7.,,\[3B?3VOe4WI6PAY1Kb-
:4&,?eE>@<Gg4US<@IZ8:bFb=MM2OYI8>70PG[P;3T7>#5-H6Q<WR.074AH44d=-
(4BV[b&W+-99WH]HERPD@CH5)C@b+I4AbbIeHE36?81IBKCf_Pe^G)P(69?BL(KE
.^].WUK2LTD7dY)[QY@UVc4.@Yd@07e=B^&[I@QQf?EaJEEaJWXYFX<C,DJ6R=.P
ZXF-T1&4OVVQT?YD;\eU,_d;WKgfLO+?6O:[5U@4^-V6D1DGIP7X=R&V\^AJf5##
TceS>E,.]3f30NPf8@Oc.C@OC7a>cTE@#L=NV)UGaJCbgV.7;B50c8B:Z?X6OVIB
D834Q<SD;DLTJE=4:I#=K(fBIDV,)/HGNcfU4[.6VS6TNEG+HMG,G5-GSa#1-.ZU
[Ffb]&R\.)1e=^6.2;29]RU]>K[]ARO56F\(WF_WM;e2Kg>HO#f\WBEV:B/6b(8-
-e1.-R(?gE@(V[Q1Y7@-GV,ZQM+WfIP-GDZe:?Mg]_]XL2-E@,]0H.L)P1&YOg)b
WN9I_d@BI52+&RNLKD&:7R(/d=?BGW#BRT;-.&cbacMYfL#Bc8-?[g0cdC3dP7J6
36dd;U?0WIKM_+3bN-DL3=HS#ecJOb&HgY]B[J^VZM^TM9FOeH)5M89AJD2O[Sa;
[##X@:4ZX]NFDRA59\@SLcV\6#H>A4Y&C+aMAL4,F@6Z36M;/&X=OC;cX:8d=S88
GFQfbO8)Z0?O7b.S:LA/@@[.[-QB0d^DN72bD;[V^C_-90J)2[83DOYNEUX6aF_&
8LE94XI#\\[a4NY@S:UP5dgI</]_(E/:=gPN]5=Qg:XS9D^Y)\R4Qe0_C2-)B<F#
VLP99?[1TAA.V=ZA^fK-1Tc74RZVRaF5GH4.HVVa<]JIB=G#>e4ATKLOZMBQS>+/
,N5SCEbe_P]Y6U4e&7V-?M_DG_LP4=d.BaQ/&R[RbBJPNd7)Waa2NM\GHA1CcOe-
GX4=#V^]0PbfN/RS^4eZV0YB<bGD.A[RAK[7S><fIL((@aV?7G<f-7)AO3RQ>B[&
G)fRO>P2A:/TQaO7J,efKNOGBcGad9?/FH.4\1[ebBK^?<PI]gP,f:=)>SfYEQA>
UMeHZM>0Z?3_U(83M(fTN]Q&@JH@d4V:WaB89)J]U/\L=WG1++I@7DB\=V(3RIWK
^TGIIZ^0@DB91UK&_5ELgAL@Z4M_]>U6854Q:(GMaL3cHB#b(J..=(QIQ6,V,43F
<]Z@Z[K@7O=<TNWU=C#VYM1:@0WVT+N1#/@0#d]d?Z,dEcG+,_\-a@6:I][O>^HK
I[W4O0Dg&2Tc.abDCLH:&<ZK9-Odg<Jc;,C_fLW+A43D5MWIC4d]GB@(YQSI6,9R
aeS:?a=VMH3;fCEY-GANa(\BT0PS1S[M/Jg)UAY.H4]I>L_<a228KR\f<eCN)Z#T
aW8V]F][UbCfGH8NZGg9.T]@[0;CBE_Y-]J;]@X7-]QW#6NJ.8#5ZV4L-7C<c]KB
P8PeaC-aHC:+K_8)^f((/?:WH).SN,DIgLSADPTb2X)IDQ&#BK8EB(9J#]Id\Q:U
C,WP2FQ;W]J=J[X>/R]#3.YWd8+6S2C?]@BKb,^STJX:N#<W64W;([[-IQ\7N+)9
,[eb[O)T=.N]PYgX4(8.5;?_Vc/G^XMD.=(21D9_8?4L9,H8cMGQWH5;U?5,Z3@,
>19H=#J#0]_TNCA(F8ZYCGE\NS,OK402/R7=b3f5eD8E2Ag:(UcK;3dJ+F3G/+DF
TUY[,+b<8GH3DaZ?(\5]4_YO0f<:a#6b+XaNYA0CYg#L(2W-^_OW.g2aH1,\-GT3
/dD#UU:#bb,FBgE1@DbN-O1RW94?75Pa69GRcGGbbfFdS3-a2>O/>=2aJ$
`endprotected

          
`protected
b://b.<OUd</183[baO3JIPbC89>F/X6&ZOa7I#fbJF_bfa8OIEJ))MRBgE8H1g#
aQXMUgQR:f9.>J_C&1J#?Q[:+SY#^FH/J6[f,J97>P3_C$
`endprotected

//vcs_lic_vip_protect
  `protected
dGd=T1VG)UbFaGN?@E0;5]ZHSE_\fc+@dM)^g]2[4UMQR(EY<gD_((R+#I.2A\cc
XJM]XBYR<<@Nd#fG_)I:fH5RVK-a+45F963I=/SH.5?8TVXeG]DG4VRG;UZM>308
1,B&7\fB3>R9Ib3M-]F97(PAEfS>?SbE)6DCIcDc#@;2,/-EA_A7ICZ._G,d^G/?
_b6gLKB?H1RZ2fR0<fM^>I4FJgRX:-W/#;S2Q;=#:-Y9f4]\&-7T4-He9OT)3Pg7
X(9A._#<HJ#+K>+HbIG^K=9G?gf)_N\96B8M,.f,M?(0\gA>#1>#GG+e<9:EUWK;
^#d70C+,L[#F_>0JQP01/&#5ABbXR\B9;?3bVa?;3P]LWLJ2?Gd/MZ_9&La,M7&a
BSUM97,Fb,09CTP[R#_BN:\+_b][<b4g42Dd-SL;Y:)LZ9GLUbR;:8_RQ@6c<40<
[f)+N)LGaO13^3GAZc0W^J]>D.EFe(FPbPN@]F-@UQgIBY1f:^_g@dZJEf#Bd0-R
eZ>e&J3a>8QBU_MMb7->1S,9U4RJJJebJ^Y7HW+5fNOZCWE=\e2]^^Id^0/Y4?]S
^IX/CME](]-UH@>&8(e6g88KKVTYIZU1Sc0)-ALL&=X?KcJ11Y?#?]eIA:(89feZ
OM2VL&1BGQDN,9YCHX4E[9\930e-,[9#KDb@9RK6Of.\g3R_@3Qf.^<_+/9b(Xa/
DDUQ6MgB)>#/ZP16&bL=MNQ/[,Vd&2QY8cJ/-(,PKIK_Z;W0-5<H2O5].7ZWMGK0
Rd#/NfM#<C0;e_:S1cG:2GFO9UAe<[VRCb,:#F[[P5:>AZd)^7P.?eQTfSZF>f7O
M##CEe-<PG7;.$
`endprotected

// -----------------------------------------------------------------------------
`protected
SS,NG#SUT9&#0=T&V0A6V26[_Gbe(d-PLeMU=.@Pg)/5AQZI8Bc#5)M]-KU66X^C
#K0FDB188Rb#0$
`endprotected

//vcs_lic_vip_protect
  `protected
>K+,3XM;3TUe)\;>LC<&EB/[CRY,6[:QTO\>:\L4(7X<_74YT7c]3(G7H6cLI7<R
L-2R<g1J0?fdW<W5&W<aHa/YDT+eQ4&+R-cN:12gQIOVZc&J_#:TfFM>+]FO\/6-
Xe;HB6QUAE[[+W5\,3_P;5S>;g98gPK@Lb4U:=VC2X9f=3ccEXH_Qd]c#]&<c^-G
0#KF5K-UL\8C02L:)OOQOKbDC;L@4L]?S#(Y-YU>0R[M1eQ=e>K;[X5940R>+?=7
>@ZI6E9EXIMafd=NTK;>:\A<W^[8g0+322QD_8>_-A7S?>BNFGC[BOO,8aVHX2VI
+20<gJ[X<8XNET6)70.8)(.FOgJAEAI4N<f/U&B?XdW>a]E>3MQ[Y=BOaf8gGRV,
fa/S3Wb]g?#DW=S?A:B(;-cAGe#=KV/MEK6cg0Q\+;+R\=DN6a@GQ3O4Qf9;&E)9
?&C/<P)BQ=)OT^FC2Q8I(@2,6RO3D]U#(Q4M(F/EccYYOGB4YNHW=R:VK,E_K\I:
-:a),T^5#0/AEKK/[_5M,.>_I_@f#3c>\8UFC/(_aIUFa:2<.=eG4O=N9=[(WY2X
W:g:C]-_@G8HAH6AQHb6\9-WV-(-+\TIG3B7\<UW7NN:fHW.GPd6N:Nd)TYZ9Fc^
A)A(6])fI9UcD<:RJV8#RK^.Ia-82FJ5]FZA=XdHI+8A9+KT<9aH&CIPc0:J#P.J
#-\^VBS?HaP3^(2KUA(QCEI-#g=59^bIRD_?PIO2M)=Ia\b9fKZ#Fa15K/cXVACg
,,#c[^Y\S<LVWfJ;&&-WV#K^,(5?S,OJ==POE#I8W(-MW>E2Q#KU+>;F]dU6O>[b
E);PPIb7a95:AOWGRbP]c0;8>C39\V.MN8;^)A5Q6G4]+F^]YPW2RLf8_B4;AY4<
KV4XU,g7LQ^7/(F9<K;>N<#3d/722<;#2P<.U6KY3<fc4Vebe=SS4S/Ia+Y6E6^-
N0QK2YbHP9^AHXg3P,-K,S+W174a7V<-L^]dR>R(\g6UA3-@U,V10B/1;J&Z@)_c
RQ)9]ZZ-/S0#Ib(Fed@D@&YKP:PXbbPKg(8@ZaAPR,8CPI\YAS5W:0GdD5g><cBa
Q(@@aEK3#K2BJ29fN8c0J+)=HT4CT\?&:Mb[(Y(Od9bg7GQ/+g6+#/Vf3Vb_B#8>
8=GH-;1Ba;<Z5>FUB0NY\cfB6^2)&&\=+7+]/Wcb7bO(X^A7Z(7\WF9:GDgHB)2G
/ZH66>CCY#7Y-@6d\(].@>LSPRa^@M(U>E7bVAB7#JO@N&A:G,?.PQ,CLBg&30CI
GB>Ta67c#MK1W0d=S^TR=3QcTPF6V8O10R/WDV[U-G6)P\fOKeb[EPLeV[P;;K&,
463,YZgQ?.V/]-H]f<MHQ(,VQ\?W]J=+.UbQg[X>10F<.78VU4C8#):I#aXR7V\E
Q2)&8/SefPCB)261a[f9Udb;<=9ODT-@[SG70fO2]JA4_8Bg80T<282?B+gbTE(0
8X&6NHb7OZOUQMJe5^TaPO;_SI2C39,Q&)fVD//d)a3d.9K^>C@+><f03=25L6.@
7fa2&K4>4?B,(Y;ZLb5S1NcPH5L:;>@W2LA#7P?,LI5Z9W5\SP7_:e1cC.][db?c
gICfJWaA-HZI2F:_L?-cf6C&B0a5,SH,g,]4RDSOVSLD.5AXgbf06</+IcC?A3Ad
+MZBPSe:MgbH<F[CC;=g@:P6)b&Ga^QXXaL8S2P2F]4+M3_SFYO:.GQC\4[gD22Q
DbYc60gg>QEO?a:0?J47TR7cKIO+D3)[6L+L5<Wb\FGfK=[O4XJP3O_S7JFREZcO
KKS7;D.D/c8]Z&B&a[JTe0agS=;1YX6G7-[DIJZ8>2P<gI:P#<J5eF2@VQ3CW_ed
+IfePd;6]2-MddQ,D@K<II0^W;X)?)&?3g<DOaE1+:[-\WNAIg9NF1eRG&JfY77Q
\+5CS?Q((A;D9[+gg<cVX(2.cI?BRB54N;I?dYEcAYC<[fa/>)d0.,a+E)A4/gC;
J3W?#Ib<8L.c6YC@dIW9R.Y,2?7D>MP+_cdKGM:V]OUN=4MK2]E]OI>T6UYcdIJM
.6<EDb.755P_9I+\Dg,F3F.N7/SV>&1(74NIdYCgS\4abbWPWZSeW#Fc(b5B_EM4
c6OJ1b,-Z/63A2L4]QDc0A4P-UQC+8(;e=1PE1]]FgL@DRP),C:H?<U^<TA=F43+
Z46FD2af5gPfa,:H)7;6V<EA_GKSeFe^a@D0&4E\O+=/3O1ND3[7>E=;JDFCL-=@
;-;;JN?SR#f2,Y;^_LLe99]T8_@P+V)?^Mb_CC6-W/3<6=C03_Z+PVT3\[[[O0\H
>aX2bQ;:;+TfKR3EEVWYdZKONa7RKO5WRHS485Zf,Q@09V9@@&EAIW6[+\g-??32
_NZWDN&=/)S[I9EYYTeA;@2EGZVGH#5C^[KJU@^\[24#>-VXb,]+c=.AWE:QZ9I;
J(ZK4YT?#?L]:RHE[9bZ00=Y)\2\Q)Je^)7g0B=QYK5W@A>N2L3cKScc-W]d(;/I
A^QQ7LdX(9-\4GX&4)NZBBO?P,_>YW+4#+(bd9GXXVG\_-<Q+fH&S@_fM_BAabCC
)&35+S+E7bB/J/b0AGdRFg_>-[FBUV1cPPSIg\-K<E_.>>&JH-a-Q7RL)8?B<YCB
@56F[YMRG^=3LIXSNYFd#3.dcG4.9^GcJ.6?X@^S8+Nb96F0dcBS1FBfEY(H=T27
/D;fZ-TMPXaf(4d5?A+/9b2/#@^O0U@86JU0##FJK-cVeQd)L=&7WH(:c\7V#J4^
=J_;,\/ZfYeLJ_SZZ^5T&8_/(+We,ELBN&U:IC&McA>1e7;T?G\+8L)SdY[=Q\R1
0^0SS-NC;V+-ZNW#7(g@/PbcFOf:;>fG]K#MK@3_8Zd4Hb3P(SDC&=1c:Z/.&S]\
_cfS7+/aW7A4X^+E(SaV?AJcP497(K_=P<72WJ539>65U.7;Me&eOG\be\.2)-WQ
UWbc@Q1^E(b8?aT6@TIK(eD1/E9#AcMD:P4GGROFI0B_Z6TVAYVAb>Ze44U+Pg,_
.&/T@a#SbbX/TCFZ#4a9^;bLD8O/\8GG=b7K-\d)Z1b9R9>H]f+3HgeYK@)MSTgR
F]XQQ,392A\#_D,A[ac#(2U&D@5Z-FSaeW6b]706E^]>G+9##bZF+c)=2\#=^dL&
3FSZ>[O9&NMC>E(2O\ec1cB9X3IW_Z:E0[D?>61C8MWA>Y3PR\@ZIH,9fT\8eb^]
ATTX-G]RH^b-=MUDbPJE7^BQ70N;GgG(\/9+8(PQbcBU#/):2Y=(L]RWXaCc#8MY
+X6KBJ,Y7c(YbV-NG;<36GQ6fNNYJN0cMY-_+/\72I\JVF5a\]9\geNLQMRNFE4P
RNZ^X,=&a/L?@3R(Lg.6B^Y#Q[@0<(M7^RM2))D,4DQV^MJYR7W;V[5T624#7d88
0YT^QHBS);Ye;JY20GL0eH4Ud^&C#RB;eg9/=9dECD(g_EE>H)MX#5PP_f(R6RK0
6/#+6d:R3Q2EH;>-D;0f)6fA0>F\M51&ca9T6MKB,?3A\D\Q4S75c?eT\YeSITC]
_R[Nb=-ZOHBed&5GW8f\ZESW#&W]DN#Vb[J1e0cTV;W>>+Q6QW#LQR3O-gIV[d(0
_E29W0+bZF[I>DSP9.fF813?E7]0)]U-:(O3:/X3f]g@JF(gH?a2FS1LQ=_\J:,V
2K(/PD^bAO0Gd99[)QD2EH4&.74FfgG+12<&aUB5;O0(>eVa#MHb-F.?D]e0H29K
\B:ZC^X0864.Y##=H+;HF]^6gd@[&Cg+S7679b70?AZYZRD4T80^TF@bOZ>Qd^5f
c/0U5bM\+V7gdHXNMHQ^eMEUOOG^FBFILa4=;1HFM.HL5GP#\(Y5\U,(4D_CDM+(
\]3dKOY58PE/M0Y_K\P=_a]76\32304b222^BXND2f-L&cc[3>\eH>8KXA-&@9F,
EAb\APGD6/-OA]TLH3V9Hb;)7Z5(HL]<@A>/5UZNd+JCKG7ME\H@VI6X7+Q2d@Lg
,[&C4Q=3>bB>U2dL6_Z)N,7(2cH^BOT(Z^+.QGf9F.AS>ZB[9[c=_?AL9=V+Vg::
,A;=NUI_L;IE8g[A7C:GL#5GV3&UgB2/c5-8&([FE&9)25&Y9/JKFa-]6AKG-Tf4
NOQT-3XC#;A6OP8_,VWcUdFP8&aPB0TMgO9,6W-FHNBRAKO;V:6G#A4VA1e2M2@S
1K=_4L#D2HeQ8H\_dN\<K6H_(@cO.A+4caBB/NSgY3DC_dRTU<ZT9G26E(DUT(AX
X.\Z+?+cTN9CG]_8YG3PfN8_a<c1798g;@7Y51+Q]F+?85gX]SVe3HC4O]5:c-_.
Z&A;U^XMW_27-MWC>K#RAZ5/[P5e;XM(M<YgX796\3+YGGQ/c22:aO>GaI<ND=/Z
;C.8LJX[W^3Y>C6N3MEg]L#I[BADQ(MAL12K-:2.fF6\B.\H>d.K-2AH@]8WQJM^
Dg_YGZ9GVX+QTLGI;@CHU7;B.FXdI\b.C;6;K&+LO]ORI9KK]IZeIKPSTAf18aW\
B+IJOJ_;JUSJdG;B4Z0JG^&>@6G:&]-+PDDTeNY@&3UMVgRER.2SVRd)PA3+R_LY
E7?Vc#F7)=NM=F?ag,dFJAG6c-g5cKZ2LC#U6T7BI+S8HdRJB.NL7S^+07+U<(,6
T=78cU_MYUTWI/M)M8F5PWTS7eXOAADGc56F(M3YV#Y?.Z^,JG/-XXHR,(@TW\,W
TN_Oe736K&)1&GT^>NJ/4c,0W8GVV5ND&KF]-BW&LL<L2BH]7223Y\OO7XPbUaEC
&Q;d#N=&9^XCE8c,MaA2+Ze#P3]P/R3gBW&R@eNSDA>U,E]fQ<VA]#g\>aQ;B3&O
#d]H94]f(5;U8dGbTf>5.\;LPPA:cEGO]T_6>,U\6=FI@LH(Dcg;_e9UIG]YV4>#
eAA:]FHG[7RY;(_R3_[]6<,QCD\)16g)>M\7?7A>#4AZ?;3[HRTD_F7c4?[f5@Db
50JAf+47XYAY06SK<g>]H5&fNBR^Z917NH.fC<\-H@5>U.^98-?_:AES\E3Z8b)8
].)?8XNNT7O<C8Cc?9>1K^_XWHI<[<U:J8&YE:6#f>Y1,=TR+U+;Z5)<L&I4AW(C
VPJ>\g9[Z-XUQbZLF5(Z(+^QG00KAgC:HNL)FP3fI\2=cEFdHPC.TX;ZLU&]<_],
U7d6>LHGL(N+cdUXfe0KSVfa(38EH-bFgS=E75.4a(.\<MbXgAaTKKJLI#>]OGf@
TY8-CQ&Z0E47.[,5^XeS&\(+;(AYU6OB&50cGfYe(P^NCB>U,#HHTc8H0C(4IP^?
/0.^W525/77=IdQOIgT.N(AR)G9e(/ZX7>M&S2?LbO1X-Q1/F3g9E#b9e4<8J:X>
9NfIf@/\]+I:eOgDS8<a-N;5aD.Q22-T]^T5<fT]a-\Z[Z?]:CL.?0#J7RKYQ;<L
dNE=28SL2&P0Hd6ZV5P,N@MX?@V;L1>U>P:Y@^6_N@(FB3CeO?e,ZTKW4X-^:8;/
ZHcYK56ZHU;fbeXT[5CfKFCb.6.B.a;,?7DgI-M1eQbBI3,gHE#RAB-HYUaXZ+A2
7[fUEBXIcHQ4:R@61I]HA3Qd\F6>N(PS\:JbQe[&fH5e@Y[C90+X2PS6X9FEgIK_
Y?7YERec,,OQ3_d3e+\S1HYdg<AA-)N-PMe8V9JLTM2S?\037f?:Nd00TJJH1ge?
K@BNZe)-b9N88N]?JT2_4QBC.-F7,WB+:FFgELS=FRO?aFH/S(E.;I<MVQ:29&D,
[J?ER:VF;ff/Z+&L89(=7.5C+0-Y(+]Y)K<W];;Z0]HG7N&dDRC<W68?)5e9/))0
_^GZ:<C8.L3I6d.GQb2D6bSKMFF@bCc_LTA-TO8bK>.:f;cWJdaLRE<2WOM9-IV?
XJ9LSb;#bZfI=\0aQ=JD2fVgBWb-=eE4;4V>g5#GPKQJ6N;4290<KcA:,,3fe/gH
L:&Q.YQJE+)M;9WCb=IZH_Y97_];AeX@GEQ9[f,TH+T=F23+E_C90P)@+7QMAFU1
FX[7QKD:8Jd-4HOM814[HZfAW\4[@e@81]V#FD65_CAUIDSKN6fYcQ=SaSPA4HMZ
3H4A]VOT5d7B:,#,D3XPaE5JU1]Y@e5a.\YS1\HI,b[,G)E,5>RN,X1P68+1#LV3
2.cYe2b)aG,J([dcA3IeQ\]5eF=#5M,IFQTAL1=056AWd4YGASB:F/C\7+G8_J7B
f6Z24:,O6[H\OIKb;;0OP;/&Hb)>58bUD/PaU\2),TJ6/TWS,KP2)d8LN<N315&J
<Rf4US?13N:HbfRE6=BD14\67E0R@G?;aVbb(8:<g?+/)ZU#DI.,2@,.6+M?g9(5
ZUGP31MK=EUK1BY^]\D,+e(82\B?,?_d-J4ga3aR5c7bFfTR6O<4B0+?9If-5W=T
A[+@P@Gg/G)R-\=&#\@\TW;:6W?1Eae#/J:b52VS<<Q-/Q.g4<G=ZO54-(DgOO.]
MGEU4JWJ8cAHR4ZTQ(S@&4D9WNa&P(c?_ZI^TD-[<WA>\_NZYK\8Y.IR+LEe(49_
ZMQ,L/4/6I8=J^@dM=IA<85<KB68V29<+:&6cR;RF;&A##.V?9fYPF\B&,)YR-_)
C2<]);OQ[FH>=KH+A:WDf_:=Eeb79eYY>ZN:g3I?RIA,;?C?B,c:B+XBN]P=X\@<
],b)];_N1cMB2E;3-]Z;QGJB@0N5=94:3bE3;KGYg+bIa2SdU^8ARV3C@,XF?U=@
D6N(g1e4NWCP<Fe?18;?e/#a<#,5+d.(8,d,^dE#(@K4\@6Z9[ec8gd3IcCHf,#:
fF0GBa\H7aVND[=LMAO9RQ(@]Y]08&Ab04f)=a[QE[2Q24XP>W7GB.;>_9c9??/8
c=]f=CWQX-UcGa\PBb;+I>X.R,(.&RP_Y52FMI_O0@4&QeSNGdbbB0Cf((.?>I(S
])#KH3I+F.AF:P&IMbEM7+cBJ]MY&b1\.TG=\VPNc]YBHa\<XU,GOGa0I>C>JC:2
Hd-?6(4875>0R9-KMVLa\_=Y(bH\&LdcP&bCKc-E8gPY-=Sf1-H(>]95;dY6_3]-
_1Ba[EZ\(?3KQ5,_ZB,^NXJN]YPf\c7DM1_+^:T@2[,0(E^#U]ULf8G[+bB+BgO>
.RLf#CdR0cR23M7KX.UB;)2[48L\B;d8M=aMITP:.K,QaY?&>:e32P4QX)HNM6fR
-9(&b.b)<:\Q/&JV(L,J_S=?57-X]BW]=M\WJKUD])e=1,#?Pd#X4H0/WK7J1A-L
K;b.&_B,:FTYCJ>D4=>(6@[J^>5E^ffBS3H9\?EQ]JLTPZ:SC5,KUBRW_26@eYPN
I39fdJQ(4QX95DI4U2^=(XWV#U5I7<)5=Eb-FDeTf_#,HW.)I]:PDG3XCeCaG:A#
X=)>7)^=6gJZaT3K[L5G_KefMNf)@e^#QX9TNVJ+CGC6&[+_fE&_N-X94.adPHd1
_^D=Y;MXfV18\</G@&V\KCeCOdSA,S,BfU[3c7P5N@5Q)928+e-4=H6PFP,<?IK=
[(7\>YW7PcQ7BVdIfb>GFAa3Y^F-SB<K,c6<RB6CW=QRKKU_2K#5OT=9=7aQ2S]b
<c+AbYA_8[/+@SA5D(O(61A+XZADF_)CgORbD=@Q1gLcD@NH<UT)&\&Y_?HHGa0;
DS4#)&4]E3I/&U]JTSLLY&V=@_08Y@6E#[&UO;?g_8.3B^Gb67@3e38T.+^Z-Ce]
gT:A6,2>,(T\CMd5RIVL;gAeVG.\<7[V:TQbK]c&[U@8QZ;8#Jad3eM]E.MI3d9_
.L;B_FZXTJ8+:28=EO.=H?6.>.aC>+fI;R6^d96Sb3/H14DBcfP>P[C9Z()(OY>)
GD>cK0OV7C\@]K/S?N-\;9(;L[W3g[HGGF(.JR(1Q76T;[VZG5G];^^H_aX@;6#R
-##Sa7R)_OaV_7^6+fd=BTbAPBU-];V-;;\5=/-@K.F+\LG)#GB>;K9bXUM_P?[?
?&VDPV?LWS\^GEC>dVO@Y<_eV4d\f(=FA6/4Y<EC0#BHOW8fN(+TN-80^e8NRCGb
];++&&R]SQZ]HO3&=+SK=XVaDCV4EJU6J&a-Fff+DA4@0O4R-RP57WbTHR,V8D<c
)K=MA\EIe]2Z:MT/UVaI]--1MS>,gS)b.:[7@3&6:Hg2O.T_DHZ^NSU3<^&/bO9@
gS62)_P_COXY+CNDS5S98042)[B0J)GLHIH@F??,F_OZ(#H/G7TEV\4I_K)(&SGE
[a@)U9GM6:+;J:Y1G:c(G6<Mg<;NS4D44\[0NfO6S>D\OOF8BY0+#.&-0<G7aLQ&
CL?#+)Ma:d@U;MZ3a?@@;F^YGa6\7XHLTX;RI=Ca?O@c>U&eGcec=JAO[RNDD\P4
N+UA-J9A,V:g^,ZWO5&IDS_[6#]OL((YA(9@\6eAU(@f?4.GO\Z\&P.(=bV#Vd(f
(TB?a861_NGI_Va3X1c.bTFcZNP-T:[->_7)(?[#/RCVB8f4g\,SR-))ZaK#S4<G
LW8EeTWP+Wd8\;]L+H[T0[5(;\2cKI7XH1>V<IVZQ]NCI4350O)>=F+F0?G^>J/>
^J)&X1\^:c+2?J847K:8M?M:]T]@7_N\?G-PLFVY4[NBE<0MV@aNe-MP1TX33PTJ
VSTA[#R(Z/2LU4e]PWgR:dIR6\W,#CWHef)cQUI[K_gL<g9G9#W3D.])ag?.K3XC
cR=\V>X_(Y/3JaNOBN+_6_A<Z\SM-IbA4K60c@_&4\&V7UD0N:9ZYag<f57;9:]?
85RCRJd;YM=&JQ1\K\4^B3Y=,:Oee&K20?05AY;F@,54.aE1aWDK75NE+:bYWV85
39()UY\\P[\M<&Za1ca4<\W2@TgNKWY?C7MH^QAGKG^Y?_f3QgQ.fV(:a]>_<@^M
ef=[D?3T>MLY;c]bSC-\2OA+b+@@C]<e=1d;eCdXf-HBQP23RT2^56LCD]f@b5-.
7ccN,/)@Zg@;MN2ab?_ZGQW7WR1^5]R]Mb,A7g[B/?NS\1#-9eCJfN>T6\1&bM0-
RF)9R=7g;G7a<Yac9V;XW,F]51[QF>OMZ[@4/.OU&Wf.UN?\=8M6>DZE32+:D8MG
;LOG1L_P6QF]3+@0bd4/;gSAAOaVN&e?D1V?LZFVC)(]?\1]8/9Z^b#aUTbWeA.O
35/^&)Q;S/bC.Zc4:2L1Lf)d<?Y#a\Y[EL3MA4^AI-[32-NA/d_A&S,F(Tdc[XL^
)Y<5c(=TG=Y;)CLVFC^I+S2/0OR&:N-Z+3#UU9SCaTfc_Y^7]R.#]<@X=L>eI:]\
0H+F7Zg>3@0CLc8K5#X&I:G:a7WQN^]0-fA\CO2];W^UN-#I5)?T/&JV9DfV9-dM
I1DO2QEG;5RICfLP3:&RX;;=^G2@dg^4@=9A(.4F643C6LNS^S=d#]]?Ha70+cE&
_&ZHNgB@\ND.QKU9),-0NZWf:BM+eD-WQUT<1SR0KT/5GfS2e1/.aO]TX()L2Jd9
T,IPaJH0KQ2F:IAVaJJ/bL@?,KU>[GYV[/3C,3cTLRAQLdYO:1LKf+8GCC3/YTb;
4g&YV-JZ?cEEUIKS.MJO)SP&YW3]<=e2Ifc[]#;&IG9NII0J\Q2-.I?LgJ@<M\??
IVPE5A&6DER@d4)6KLKUg;,41IE>;YY#D1F^ePAJH>gXaUd1eRcBPW_Y#21a474\
606IR2e[GaFNH>^,<H+9<g5WBK-(SVYR7>;9aIZA.)HLWO\V_g)5.:,dMWJ)PNE2
/&UX?JfZ91E5@gSR>J;XRP7W:G<#_M:C^f)F(5CFC/IS/#[8.@ZO0)^f,5?P1JCO
L2)_<b1Q]H#181Q);#KH6dddP>Q4B2>.?GSW[L+1Z?&+F\.d<NQ4\[?&;X?b+A76
cW[K6T86\Q)0;G[be2PSMJP]-0T-UU8Q=S,5VH7Ud8dL:XgY./1Y+[8Z@EFYg=C\
;MX6I:K4bG[W9fX>[b>QNH>CG?S466WI)QNZ(WS/XZJK^5f&K,74:(>?ZLKf?Y:\
#UU^TC5\P2BMS.ISPB=)2:Fb9g5cO6,T/.9<E&&PBbS/#@ESKY24FAZbA<f44e/P
D<^)1I<gN^RcLCDcSf&SXI[-fg,N:K-/C;bE/N2BMFJBNN]Q\6f;V=+6UGd6ZggR
UC:6RSM0V//5R;3ZcbH6?a4S^T5G06A724g^(>^B0\;\^;F]Ba)/7C;>gMIP_53H
-NfQ5,Te6UW<.MPJ-@L?7YgI</&=L,7[ZQ:65)>G7R\G7[V_C[2L5-TUEUb?>Y>&
.>STC7M^)8EO6/,0M]UaRJ^VdSG/UHBNGHI,TKMK@[>SWJG;@](c+>_>&R(/GB&/
FC=YTE@\;aNZCC6E4Ld+B@.bRZO)W_YCLZ@G?:5G5P2.4eg#5OC>L&KK40HO>[D&
gN(eQSUJ>P8VV(O.LV9ObB0Y&@0>B,-;@Yg0BOg1fIIOTM-IKP2X13.C4V3FQcW:
L(COI;N+d3N50M_P4+UQE2]L;8:_=b\g8NgANMPS,+7<Gg:-][J.\Dg]ZS5(;H]1
XWC&WU7?T)B@Y][L?6F<b]aWb,G>PKA0c:/BZZ5N?GFe/EF-b+7,MfL_D1_6+=b9
86FaVG&.C[A]0e?B2O77G#S..:/HLFA#:329H=.B=W5>CEKRbgGI6XL/OJQ[OG-[
Ub_U>@8@f_8Y)M9.b2D7L=C)1LdQ\gJN+N_,ZBa)=Q<Ra\_G;Y@f0Y^YZQ^8H:7W
V4LC>EaEcK^1ZGEG2OK,3/.58>gI21K2VHcfdggT]4C;^?#3<^^/f,W:e499D+]/
/7JdCS>D4T0eN1\9ABFbZ:KKf8@VJ[B:K35BBg)R5W:Z8SP29((Y>>g.>:25Y,TM
Ie2G6@@Q6gHCK76Sf.^1^LMQ5PaGf9P+a3O(LVWgJG.&Df2Le32db8J7gDL9DU]^
BKGV/N]YQAP0?&&<M#^gH([CXFZ_#e(G./]EgM_1Z=+40)QLWE7WN(?([@40XN+?
6S&_J:\N#KVX4B)f9C+BegK<>H-6eG6V)_g6O4d2/IN;<dC.,.M9M(A-=71]]\/V
Y.X:IUJ3HRSC&Rfg<KYYYBL6G[4FA&W]6.M9bW&b)AIF;I^cX\;WQaD.HG64(eAV
bC-OL83?:3N3UV6\Lg7d8Q.M&-AL:TBCZ]cJ:#QEDg6:c^+]-.OBJUGA4=N]A>Pf
YY?.(:S#N[<ZETO-K](Xd2YbFdXeYOZ7OZ?XR9.CB[^,AIe\\f=\D2?8;?gB[dRM
R-JYfO]6@)P?].)])[BRTLWDc&6eQ)g,0gHH[1XK(Ag(Y\HTY0W/d@R>JPJYZIVK
NZ<aa\FgbR?e]Y8TXbY8R[Q3?a^6^-Z@Q[BK9Gc5NfAN\OQ1;V1U6;W#.DbR[>0R
A\&=N9Pf,H>Q,POHTSFC186PY:[Pe[<2Ob9;&N&X/7TB/0AY(cHZa:\GP;+/C(-U
[fO([\#(:@6^&&VL3A-FU#-KQD,IWca/].IZ5Q4<G0K.:9M_&?-D&&?RPMAL[EJM
=B>P=+P4+P4G6X^042gIB<IED[MUYZ,GA@ecU?#JX[#=.5P+]\8aD&c^4#N2(e\<
\^I?3JfJVB/(#.PeeGZf:&G5a5KNb.#O+\OTge4GQd(]SbGfT(eeL_;Ra,?g<bT1
5MHD,D\+;(a:>\7-LaZX/Y[)Ad,N)Y07OD#ENEV9Y<bT84YVaO^CIO6CT]^_Q7GC
MMEXW=HA5K5)0-L0V8+:b&e,0B6=R/c\\efZ2B]abMLT\M_bcgd?I0:=EaX#55FG
@YPJ;#6XQZ\8(CNZIQU1H\fdK5B=S5NaXV\+7>?a&::4-g;7g+LH#0==6&@<H/D8
,<CRP2KND4^:b-);=O)JV.<]>T_b9]]A/JPHV=F7Q24RGfOfILUMZ0U),CAe];5Y
GVQ>>TJE#8\3eULM+6f@F<@KOZbdEfdAZCbWagSBI7c0016)A//P)a/&,ITSbc-7
Y]bF#Uc_8KZV=VTOUZR2&U7)gFf0R-YS6I0B4KIeNSMN\W,5b/J+E<FDe.fQXE[Z
<C6V;#OU6dfEH88:.T:cI5@bAWgaVMA>N1<E(L^<,?L6g):@[#U?H120DI=K=R6G
.F31_CL36b=+Mb.cM(-c7PXIM=(^a.=#abb&PS?W@Z5CN1O4^VEC]BRJbJR=(P<;
0/+d?QMU/[fJA\-E)JG-K3XBH;MUFI&Edc0W7;GBHcIC,F8[(NI1+S<K+QLH=Xc&
XGG<.fWJ5.;N^Q1@.2b4Qea8AHXO_L2OV:8&]#AQ9@L<W;JZWM17dXdD-@gBC9[]
eKR,>cU+KYZ2:^@I-[_W?@Sa+VQ5c1c>/RTZ1;\\O14fCF8]/a#2.OS_,&B7\N?g
gG6Y?)]IR_PgLdDLa5_GK-d-RW@Y@IY/0RZ.(f:.YB6^6N4.;?,)E[CKY@aQ6V-A
OOHPQ6(HGM1BUcUBaL>L)Y<QeI\[E;YaA^F_\GF^)7d_&<RK1#.(1J<H/f(KU(cR
eG6;ef^KTGCH2Q5G#@/,J8;]]LV2PW+-P9S/-M&:b0H[;X;ACH0dR+aPV[PK_SFG
/PDHW#CV_?0J.@f@43(MJ3G>L_@KQ]DBT^QYS&3+e&[,M^#YQ5Z(-b,^6Za-)+F#
W:-WCa1eYLKb-PA]))<H0(2>S,ISIEZ4c^(DL9,ddJ<QN+X#@Y5aB?.[VPIf\aQH
aX+3eOU_TJe@bH8\SW+[e;f]C)52+MROK&5O;<HSB@=C-Y#=?RG1CeIAXfJA1-;Y
&I;.gX]^4;+=GUWQL^E<85]]Ra?E^(;2g5))c_bY-8JTX2C6&@8TbAb,9TeRQX/E
R,Df-F2geFPP]25LZU>XA#.D_/-5J#:[<;;)RfLUd>0K?g3?N_T9\Xe7]DcQ0MdP
^KQHGR^/T(+fYE/1d6fLHZ8HBf&dPI4FE\Z)WCQ:X&\6]HD(X@P,NUeJg<)RR>B]
QW-&TgfQ(fL+@fQIW@NDWQ8;J:;K(H(\YcSF^B&@XQUM-(b\D;Y+8I:1S4T/-Z#:
^=d4;F6=#X><g._7H)WZ:f,-7<]AZCUS)04NPccT;,N-)\6CF((\BGQA#cISFN]_
MB?&cP_aYID-aXd6J0Rb9,]faUe#COAfPIbH?+NIP8+I4J50&;XJf#(KI,[+9TH#
;>PA;27M\_FQ@g?=eCZTQ9.Yf/Gg.Q+^F_Yc\?D]5W57L4>[f)#LFH/W2Z];gL9G
6VYHEC0fT73K<bXQVMTaH_.5GJ+ZKAQ+2OLe[[]bDdT]5e>Jf4>^ET3_M@JD-DYG
[&g@V[YTO.^f]=M+O^B[FMK<2a#Q(6(?ZPKUYBI2L(0L4K]D1S-AMTM?KDgDZV?7
O0C)5/3P-WZINFV#>,L=,T[,&Q(7[V:[bAVCWM@,?GJ)[08J+SSU+T1/H5[J&8Tc
LA,^NHe_+,3g?3>_f7=8I;=IT^T0->]^f&E8_0M4HWQR,U@A8+H@@2CMC#7Nf+IH
dG^KU0]QC-aY?)GTN(=f1VdD>A-J(c^&SJN3;,WcV7><[1K=1Q10<dg[W;_EIC,e
JS#eQH-V1L6#S-^((#SC\NE0PB48_F2)Ne+aW[GQcE6;];S;TSbMaaY61;O:@Rg@
30UJ2bgW5Xg,^E@5F>HN6QAL&g=5,KgRU[d2PX&&^A]R]eP(_)-7R3PQUHEEI(QN
aGag\:X4@6I(^S1L7\A0>&[Ka]/fDdC@d7LR,3:EdHQcE7U.K;S=[I@&)ca,Rf-(
O?[5GM@9_4;<NQ5\3ZOGP;:Y219K5<KJ;HLQd#IPX7#N66BfKIU?E7>@_^M1H_,>
3:]A?LA>fV;eA:V#,dI2?N2\UA:dONd=B7Z2NH6fPJB-S3SgFaNTf1OBIbZ\afEb
J?_3Yaf_=7\?Je]c0?#(Bf4^]c6PbeI<Y?6EF8+QcM7B2YK@>(&VLW=EKC9E0[9G
]ZCI[#URG]g:IJQ,5V[J0[\?gV@8-/X?f\W[LH@E73DX6&>DJ;)aT5^8Z&/0XK=M
9@eBLL\&GN#-5?]Y)f1>C8V\VUTGPS/_e)GQUAPfUY]6B)Y\TKXXBL,<^&H<[E?H
4\U?BR,_(bT9OHUD=6,>D&aUBYW?gIW9VRNOc^A<42T6&+NaVKDLIeN)515GJAWM
#bT\<<H2FaJEYJ3VdDD&Qb0AV<?Z&3;\B3@M=1>\JYa^?KfCTG2^\Rb5NMPFg+d1
[:O@=A[7A1,WV^_Sf?HQ9PE:MC-V6>(5a^B<Vg5KGI+e(6QOMI0\U9,ZIG(Taf<)
9+JZ_87J/UVaJ+e1/f[&JNFXOg3f=L^QZ-V,e/EJe9g5R<VNCJ<DV<-J@a3I<G;K
21@^P,&e_[<[-K0+39&]c]41/.^YcVHabM\?#@ASI[SB[RW#IHA0XPUHf1X8KT0[
WVMA_T#RFKE7MPP>\]XB8ePFIKI=<g:Ld5eZQN8GSBF7Pb@Id96XSXG>&K.Y;MGV
PXdA-@^3-@(D.YR90)bV,E1e^-Bb&0:.B],BGRM,eKIFDORKY&?4G.MdaBII/@]J
2-(0.M#GeCg#59T7GFD28B08+FIIc;._-FdcS.L]D[.OE9a>SP@8WV+c9<+VI\:d
UTU4:;(T?P3Nd:]ccR2fU,^]d4@#eI,D+02=efT5c.NDS5109#LW7cK@D1,7Kf)+
^X\B+I=e<_\UMMFA/32J9(]#,=\>eLXG8[R7+VQ#VJCBfPZaM=1e]aES/a)=K_1F
6_ND29=@LTUe]6IdF?X:8Ia:NI30=UK\gWg\O/1U@JXHLPD.C-Gb.3K4.Zg1PUe-
C(Q-V(PR[+4=W80SVXA,DA,2,Mg,15L>Q;4J4#Vf7BgZ-,+@7Y8T2K@K#2EQeW9@
Md57>9BH1]ZSTXHM?4;Wb6;X)8U2>+UK[_A5580XD2QCe(/,+Q7S0g]CT&^H7:UE
bB2e_&MfS,f4S&WU^/\H\;6aMd;Fb4O7BZf]-AFfbb)WA9DfK^.da@]a>RcI99cW
<3HLb/_(O)3+M1PZQ,(./-BL=_)M_0@\_ZQ7fc]1Aa3#7YP4//M#=KM^>AI\K5YB
W:F:9R6#eb4]=NIIQda=)+=KY,#IHYB\X9DaI0G<ZBF27Me/P6b-TCZG@b=O/(+-
b+;DE4C]W5>W,[JM>HM.^E2Q44G3S2X&E]4JNIcQ-9a.Y1T8g39@2IV?Fe[YUG\F
L;WTX1&gfX^GT5ZL?[7;HUbBg,bP\^R<:egc9MC?b>[-L:BFAR,efJ)N1CQ@^V8?
VWC9MF79[VeW#R_PH#NY=Ca4eF(#FC4bIDQg,dgHPDg-OgNeV6TFLK9a.(YG.(5+
U/<BJSK>RQ99D83924BCXS=cZA0X^f7_caa#NgODRg-]?1R7052fWR\dV+GXHZ+[
DU]KE1,R?KK>8WC16@?U0g=EP)16K.]EM]9M2,a\?aJbP-DJ,A0<+ZP&-IE1R.B@
09<R1,LC@JU[CYER<2>QWKIVDcD1e7I8Ld5Z72;C/F](K9ZUA7YKA36<5R1dT6N1
a#AY/_VTFS3ZA^M7_Yb\_-=P9AeC3Ga@3CT9W.Zg)Z#V.U:GYXZfYc_A#BHJaT]/
GV(-a>D[ULDWdBB75WFM_7/JF=VFXU,7c8bBH\M3<QLdL,#II\<-WYL(XO>L[g+0
V9CG+\:LXY&F_O=<X,)#T-b:&H:(9<9TV#X7bQ=TN(@@O=)3-JI2@>]<O\I/EN/+
R.aV(Z/.@ZVD0^=a]S+OW].5_B\-aGUI2O-.[W_2PBQ17YQ,HO-<TH\UgZH>N67S
M5LJLLM):PPA&+1SWI\.RdP^TY3BaGMOQB[<bD#0D=SFL<IK-G>f?1-7ME:1/dX(
0)#EEDH.<b5GFVM;5(@2:?CITX([1TZ6dLK-1M57ObNc=,B\32GQH=[_?K[EO#PE
DC&F(g78O.?]+46:DF>B?dES1G9EQW[/)1URbcOD(OZ<YK6>43,fI;:5/L&VdcJG
8@GFN8\_#M[[M>AL-dT[6?>/c^#J6?XaZB-=\=-PE2OF\D)TAVZ(]+QTSOP[[?5R
_YC#Y=YeU//LV+(d8L-F1S,.11/eX46[@GL.A:AOTMUGB;=-OA-O?QW7/6]:1RX#
8JN^QBOO,\BZ14G24;_2)a#H>+KY[[Q@]&-g+6;,L1NSf#<NDDAE<W_35[6Ab-G,
0eZUU,AONWX=V2G)-JF>,d6B?N?I2(bJ,>7[gN6&Ae]Y22VO]&E)2.F+HECfCZU\
R0)Q:OPFR:5J/<24aR;LPW6.M1Ze59GVe2S1E@2[WcECBLR:b84ILg6S[-U9=>[,
;W_eUbM1LA#:@0S^:D-R1SRV504.+)Sc0,(GbS>]C66:d/;O.6XSJRXN8DO:^,/G
CHU.&ULEC?OB.aO_WG&Q@?&?f?WO#(8gAcJeLc-ff@[@-?^FF<2afJa,&83gBEdV
[X2V<Z2)OWGM9?+E&G+TH_GE>[H7-Z/aUKgeU7U39>Xb#b(4g\A+F3(T4IF=Y?SL
;8a)YQG9)Sa79MN9BC7:A9@+G;YEa-1DMCN&?&1/5LYaA761L(:<f/E=8F/^R32,
J@]1[bPQQd1-CeT;6NL(2<ed;#T#f\&+Y\F>JN0J#c&@b<C&L&H<;VZ_W1]C11@C
7/P://7C6)8_+GYV[DYOX5=ggTB3Z2Y)AaC/0QDd_gP@[M.(Dg)ccP,<Z-e7W?e;
4d)^CH;T<:+5Q&KbbeKGWKB;]7M:Z[fHIEL:g/\aP8F5(LDOWF6\cP8UW#/D5GO<
/EW56O?OUL8H#L/@IcFUe>]B=dS@,>/)5ddD<c+FG#.EEL#d.,J#9f7f#H.=,d0;
V7.AQ/f]B?fO3HDZ_aF1<c@#-\fU(CT?#e;^d\NH)Y;U>aLDU.?Adc=4T-\-OD79
+ad@Ug<.2.T3Pd66TeU:]&-(\PJ=WZQF_Wbe<gL#3/1J+,+P6:C#5Ld?9[B?N#^Z
UA>59bZXN1(MX<<N.XUSWPYP,@W@A45K6MJa:fFV5fPA)<YFDaE:^(3&Z1(aR]#L
TC+f9LD(eB8KM>OW^/V4Z6Q]Sf>5AHZMO_VfB6cDf7Y(LY;W4O:06P0d@3H_\[:@
&(cX\EPA561bE]Be5FK.TI9-E^BA90Kg99U0,1(YSD67LH)Gc^I)8dRNMP^FF>VH
QU7VQ+FAOJe/X<IaO8Sf1W:I,6Z2EDH,Y]4.VfVNKbRbE;Ne#S^P=]A/#YMT7?C2
\:TF>9&\GO8>M=H+dY>]>;(+_G(NIRfAfB=<Q+TH?23]:<<GI]4g1;I@40RN>aQ>
:.>)^e8b-9AKJ,KP<DA/F+)[_T;(J2S4MZV-TCT&1;:0e7TVJYgA/4F;5XKEf#IN
]I9Z.Ka2bV4#W1UbECd+P6cNZZ,(gMZ7_:82<XTE;[@D(7bFGDgJXV-fbU69PMI&
AJ\^)CHcY0a_ZQ#TPa@Qb(O6Y(J+TVbFJN)B.J57c9+P0da]>6TT0WJb\a\9HMOK
ZC5#eQGPW[B0\@91IMN=_;>g;e,KR2PBfUZ6&9Y(R;3X^cVG<#=cEe;e9Z,BfJHT
.ZQU[OdIaL&Se^_Rb&R?0W\>92XT9:PVf/L#9?c3PG90>7aX7Y.CJE4V@,/7NKQe
2]5#2A:@G46efO77Jb1-5^^<&6GKGW2bN8;Qf@WZ]PA45V]KfY4ZIEG\H#+)gGXf
SYLG0=c\5:W/_DE^11X7bgIL)GI]=,aOF=?^cZ:b05Qce3_&<FLP:W(965K>ED(-
33LOE^RNB&6^SXgFPSABQGKgZ,O747J(-US[V8UMP0Z\+YQE>IJFM7OJ]c677/c/
PT?&5Zfg[@cf@;G)B3cEC3MIF5a;]c(UR>XRBVJGNe\R[O^&CY[J@B=X_S7D,KU\
Ja<\X;VY;ZdI4PcBL[(5V(O4SA6(K9779IXC7?eIZ;QR(0<P7;RN]#g[1XL>N-41
IAYf<cNU<RN56dZDc#]P.FLNGDQ77<D,K.T#.\WO^F6JP_?CcZaG:?]5>dIc58D3
E(?CC-U.LJX]TfFP;^8MW6cF)[)-;^[=3A8a27e_=_4&TXa#+^We-218EHYN/GQM
9f)7a-0P/g<77<N7cdMC,3_7(1G^.&,M09PQH,)^>RD/5N=]@[^IN8ZGVIUL]P^b
Y(-NGA/A:=U,fT@-d&5;=/@OMO^\SA+00>)[EJ_WYQA_f.ABCS(P1XZf8aRSUFPL
ed7&O&OI\55aHS?d\03W+.D7cO,]::IAVX>_(7GSP\8=Le=BUKAAZ#M5b]H@H3Ta
6c6[J&gc6[1X8BL7&D>V2H)2-gTNSXb\D8SRBW\Z95fI=3V1A11EFG(<c2VVcAJf
L8D^4cZ-23d[O3U-\[<e(@UVOMC.\REVP2J_B.>Q+L3/W-UF^1(]A53P:1#8/]c9
MO;+Na\BC2KGcHbbLSI>e_M,/)@#a>aWa9KI1&T6C@EZ:AP?RgX<@Mdf08Z42NL:
36<4U&=4J0R<agHPce9c@T_fO7D3feE@\Tc#=:E77UD5/7@+C,@[LBKCe6Y9fZW_
<]dS7Mg;F:VY>daHD)]cUV8#LKFU.N_H1b?@CK5._]+5KW)SBON)CI3:0T<U/3O+
AS:;AI&g6\_a#FJ->BMRbJUUN/)4),d->b<KI1>J883VEaM<<MdF\BeNHAGDIKWf
QIG=H=_XGDW<90HBd?Kg>21<cS=<6YF#eM:X=YQB#HW)d^XUaF#;9aEg,aS.D1/H
4^?9TQV11)a2YGf9;<fQQ=_ICN=))?\ZYaF8-3+1S\E3aNLA.fUFC>NHR2C2@I3(
?B3@=YCJOVe2Dg^X/<aU34\DY=@1:_&H>.^RdRDUE?SGS3QK93XCL;A\R]M@K.fA
?CF:=J7<JV8U3[,N@KL]25gc&3b?B7LH=feg<V#/45I\0P/@QQA916LMYN.W7/VH
HN>G,7(XcE^/#HYYYfP#WUb\S-(de[UVQ0-2b;JKBa?fC^S]PQ;XFLc<bE82MRGL
@KOA57\E[)01(:B9FC>&R1T96DC&(cU5J0GM:;LT:=1_fbB=d#69PZ^e4.STQV]N
Z1.>(3EfIRS8&]@>\Lff1e]W#]JPJ3UdQe(4I:AV>CWf[;?a#Yd;Y]gfZEF8D&\-
T@+:M5_(aMTA\,Z3Z4<.RR/9;GMP(Lb-gg5GLZB:0fc+HR@_c6&?K]AAO3d^dg1F
HcU#c]J5.<\0FF^)WP2?bRDM3_f67:d&UR/,OT2cK&V,f0BPg1Xe66@\G&)dP8\g
_&.0I^+]Y>09e?3?IW#4;AaT0X-_bQ41C.F_<X)5PCM&9dAZSA:/\YK8]aea28Ra
D9Xa4HDD:0eP4[F_MBbNK?VKIGSNFRQd1,0P>126U#KM5N4&B?4H/a9#MZ]IBFDV
(DHUMQYJ&eg.@Y)#?)>5g<\MU;g>QS\?XP.81^5-G-e(=:3ZX7V<BIC>6Z2>\R2I
>:+@-#CTg(YgS1SQa2\X^XbRN]MFD3Xf+fFYG6P8X8TNb6&K4ZS+@FPY,Q:,A<Z^
_-DP3Me+3;L:gMcTUf@W:,8ZC@PC&,I_V<I1_]Ca+,]U#5L(N;=DDY[=OAC;+))c
e\@F25+7_HfALF,;ERCd8P]HJC)5F6.c/AD;X7C0NR>TR\db;dXf49;HPR_Cf0J[
G+8IU2e[=V<9G8=Db-@7R^37a--8PY&8N>OC0d>7AV#@5R(X6)ZM>C/V]B0:c?E3
8JQ?Qf^:L6RD69NcL06H@_^#FY&d)GKC7.:gXW=XKc8aG3+??>38\N6O/_U9&(4N
)=[f;WHK[NP?L13I6,,@275_X,b:.VdV+X1#JPDHREGRQU=XCJBUFf-#8)BKAW,7
:.dQdEL.&A5KA:e&^L8U^DP5ScFZ_ZPeTJTRAH\O9F4=2;(GYE408L\/EPO[He,C
CSPA?K>Ce]&</B<523;J#T(_U/I.V+@AM=I3&@C>Bb5CV9;gK0deZeV<e;aDXYR4
3UP<C?GJ-V^3SJ8gOJ8#.1KB[]@VF0ZJ:J>33:;[J+^GegU@YL@g?9VYCPSa9R-K
8_R><OV8fE88dO)cL1LHgX7D7Vc]6P72OPa+(NFP&4R3Mdg)BbcU5T2^22Q^3[4c
,P1P89b?fE\J9+GMJ3)M\UcO)-ff(=<K7U8Y;ddM\XNASO_)N4Y2UQgDOURWTB=3
,\AePb#S3;e^U@+M&N.;-B+Wg.FKV[8W8#&D^(Zd,FLGQ_EE<,+GZTebF+&P(P.4
NFc/,H#+>EbgL@09VI[<H]Z2RR6gMBKJ.f4?#8gFEU1DgVfF(]U4?L=-TEa74@E)
IHZ-;AHL6cJ]Z(A@1e>NSOgXN2V.8G/#Te&1J0DWPN=].6BT=G2(R=5:S,@1Yc37
_KBE#WS^b1NVJGd)-OA#W-E.Y.#E#FJ+,WJ[Q#R&-?d?gPO6()2,S=>+d3d.:@VX
Y2d3O2\&AG+:KMDcJ[Y-.GX?f0=X1OBVI+KD/)b?B[C5>_bgP6_L)S\T#UYJ/JHP
T)SH#(URW]Hf?P)1E^PM\bf8.Z\GCBQf=;NJKCHHOPN\P6KE(&\e]^0(4E]1HA_]
X8f2]_3MgN.(?d\[PX)4;+S.<JZD@GK(;21S&Fc=ZS@5X3K(E#0(40WQST^0?IID
_K[O&6TBLUg6X[[gS_UdF[.<&TBCMbKcAU/fV9O#H:;ZQR3]NPa>08S>2a9&a>7#
?GLWOa98#>V2821N8<#c:/Tb><Ha2U0_F0;X(.Q(cfW6Pa]A5,69d[JHZT><&/SO
aceLVccRg6BO,+?2Y>?P@9>@-?,bZgHQcG\fccAZ@;@ZMg.TQ1(1K^W2Z(_>13.U
+RR36_)72BMT;)^L_N-;Q\KH@H==91SCf>(WedMSR5f[VM71NJ1VSM\F+P-PVg5@
9=&>Z+2\A]^5:D:D3+EKcC([\&DcV,3/VCG;L(^EQ+HR\E_c=dQc4+Y>-@bXTZD\
PVIY+Uc+/Z=7=\SS42aIcR)bdL@[9b]SY6MJA^U/VV2.MSUUD:.&06(I3,=KT<Xf
U^E@V9EY<\-:VbII=_fB7dbQA<@KQ:=3^cTW6\66(4+dRT^[61MS5A_4d0>gAH1/
D,J^F)\HL;A9/Y?;1.eJX_LUaKWX<c1MF#A/7BYWCHA@E]^LS2AA]75M]3+R&91c
f)eJ&&<.2G1NJR&?QVW1dL@M[c_OJZ?f37^:C.CfW,&Q@/7-eLHb4,=W7Da612=-
g)3-gHGCgXSE5E<9TR;GB8NS]8Z[+SGU_5M;(4E@I<O2efA.3&4;eE0RPC.5VU1&
cY#&#[@CCR<M.=DgP6BN63\1cHgG_9Z__0QacY5/+K<P.TIdJfCB)CX=4F350:30
AUYEBg=dXT\W:_.X<G&c>/F.]170J7S?LaM2;HGc7:=TK+G2>D@2]-YADBdKC,d-
FVJg[P/5K?9dROP[8[BPKJaY)]\M2BRT4?-6,6NT)\BN[\&aG)EIW9a8+#-P_:bA
-,0<\+JPR?f)L@FVB3-]RO<./&E0Ic<Z=aAf?+8,R6G5,BfXf+AFUR7.7C_fY6WI
#cFG-<\YR5H7GcV#+AScL,HD;D<J))?F5==-VT4]=GB]e(a5c^EA,P:D/4c?;?f\
0/87X\K+cU\Eab&VMB=/R/E,?=TYMG-<@&63T#>A/Ta7/8;aKLf7dT(a+@VIfRaE
1B<GNH_QJT0W1?@.PGYHHX\,e-QUX)5(FGP\91=;E\B0;EE)O/#]f6KD#H\_?)4g
IeJD.]@6,QUMH.#&(@O2H&b;VbSSW?Z,MEMY=8(CWXQTU:3T+JTc;b.BW04I?+^5
Y/>,YLVC8b[S7;RK(R=3;V4)4aGA,U.ITC80&,EK01YdTPH0;ZYG<OSTe9&b_aV\
E/65D32UZZM:b[7:S]Ad0CU_^AR8Q8ME^4Q++Q11@PP9P3IMHJbS@X=YW5N1E5KU
4J-KeZfE>\\KILZ0NDSUI_dH^SHZS2GIe3(.4,-<[SK#KbF9&-F73P@-[-,X=Q52
/(F\SSM-_2,]T969UI,GdLcSTDZXWA;]\CM?S.[Bb32@(2c3MKbP?MXdWgPO3RZ>
J]dCgf[^LU,G0ZeM,Pd5938EeBL6f#\SB2A6X1KfSU4=7TE^/UDg.IQO2L9YBJb8
NcDWAO5OEKbC\;cI<SLXF3DLD<(#Me[W?$
`endprotected
              
`protected
R3;NBU.)SM&IV-1-L8@3eXbX9J^EOGWdfVd^I941bcR1Cfe/_^>@6)-;gQ=SE\.N
(5=3.0MZT;DdZ<CMPH[:YO<V6B5J,,J<RUY8b#PT/+f[O.4KDCKWVM-;M$
`endprotected

//vcs_lic_vip_protect
  `protected
)VBJ2R&gd&8.^Y.9La)Ggg>Yf[B[3ff#[9O62dB<VIUY)T1F((;K-(Rd8ELd#cJ;
&ZWN854Y5Z8b[cE7cO40G?AEGX:X\MQT[)7@V(d\OLS49Xc9#gNH<HF\WH01C?0H
DRgBC>666HLA4=_^KbU(=@NdE:=8YR+b<e=T(+UeJI.]AB_\X1+_6KTd9L>[\+\e
(bS;>aB9P7PY>)542d]V#b5cW7gcY]eBJUW=TIC9/Tf]@2IgNQ)LMVD3G5QU-5fK
6Nc[AfSQfROEGX#6g;9<5gZ.@a/-#&7+_Y=Uf_D.B=4=0&FZYGQ\f0VG83F^P\?W
&Sc7=#NEKaRSYFH=e&DMS-EU3RPO8fN^:Y,7R7=N5+[@7g)&HHSR<5dD_I#GCg12
cgQV(8SV@LLJ&JJAR_JSK83c?F44LV#f77;:]-1_DVSP/6aDQIA_<dH1GIQCT>WF
P-eI+g(+?;WXXF0D-/LR:OK38@,746=GLRD#ELIL;QLe+>TNfB-VG@1,:gbHC\/4
<E4L+G&SUOMZSG<@O=+ZHa:(g,EYF[GXb+7QKEXHP_3KDSBJ:,d1eFWM8Bg7@PJA
U#^Y.<O]Y0(-:JcRf8]b^NAbN?,N_f;55T6C#_)#QC-T@@MBJ2>U92IM+N=V-R+7
+>)RaR1QR.BN30[)Z4X:OR&:2=;LEN:[@P1RGVL+]3_g9TU4>UCQ=a@UZ5_f4-E?
N;P_9,1K2Q\D,J;V@NQ/aGGPJK?=001a3N=Tg/N.V<d6LZQ;cQL(U10^/bZaFPZ_
];gfW/L8&Ke0Q.&L7J>_C>?SL:1/RX4?K=[B6=UM9/]@RS,>4^DbgD9[RVZaa@(1
)5<+G9M<6LQAa7:72RZLVTNTa[)R@K[d#)?Y6/SV=.KTFH@Bb9aD>c9Na^07VB&/
S.Fb)[33X;#.b2WDZH[DaA&3@8CA96dO5MKML+cg\eB8AVYDT?d2[3]Z5g@YgIVL
5E,2)1eF0SALU514ZG>C(<?SC1OT[946)PFQ;O5[(S?)1eKcXR7,\OX?3+O3dB=6
\[=d8\LXbMTWL8ZA4Z+@B;X9MG/dJMIRR8[MA50@83_]J;JY9g83#5[2CDXHZ(F(
@+S_)>Z<-U_e/&,(Z4R1>WW6V39.SWOVX+Lb7BNFEA[H&P:CP302[M(5db6E2/@4
6M2P32a0OCFP@2N(7D7@^UKZ3NNZ41I4)N8+:f51=@(?4@L:Agg^_G[(J)7L,0Gb
LgI^-bDAT8;ZcH6cL<=6/DC@MYG#,&O=V\LOAe1T^=2K^;QD6DBTS)Z1\(IQDUV1
WD)>-#VTf06HN0_UD.gROBA>G&b:P:B63[IK@3KL/PA0QKc,E?]<)TM)ZE-WQJTY
1+1W9dMUWD5M+U[Y\<;7_WT_+c8@):[fXD0Q>K(I]eQY-9@a<<?S7AUK15f;U+CC
1(a=H2A5WSJGAa;SM.#19<e:WgfN>V->,^UVeQ?BYB71FMfI(I4,RP6=(M/dU0))
:&>&(7X?GMg7W7eW^+N+9@16X1R</d:/>4C8KBNb@:P>@E(/>E&1E;W;:UQ/;ac8
(#R4<-Y/d1V4;bb9Sf=&<8e0RU8d5P8R6ce=QU:M<bJB3_^4fXJYCR[1EHKRL4UE
)&9EF#8\F2TOJY]TX3ZM4NaddC<[d:3K@T9ST4P:DG.63Q-VcPLDg326350QZbae
V:;H58:(DXZ^C>=VOH53)&OY\G>2K+Z<fb:^J8BW]44c<R8AdS63).C#<fI=aEE\
NXe+;MP.gS)b:.39+<Z[I8VQ;K4:R[G^@;3X=5XHE-V-f&2\c5HZ@E^B]8DLM@g<
QW(e\]We.(7M7H522MR=NYWCe5].-[#AF&BDDJ?EM)Y3Q9(d>bfb1aMR3?ZLgO@4
[NKMPY&^ILGdY67CC].Gd5aWZ?:\c_W567=FUC&/24F4EBeB</SYHAG.KZF/7AV5
[-M>J,L\Iag<\85V9Bf9Xeb>/3L:])JJ-6U;;V:;YFbSQY+YSXUfZUDeTJ=R0PSJ
.7_8^g]9@f&<0?gc1WW0(7KJB56:7.UVF2H.-NPZR/^aaLEZg@VG6[d\aHcAYJ6\
H(MKU10UXQ+[cD7LJ[[=\ba5FN0FN3Ze)P:^.L=d@TfV86Y8&L348RJCcI]GQE[:
2[:RDIH@e>S5#&OF&OSZb-,-2gF^5N&1HYH@PG]\LVGLP]6a<cIO<K2W)EW54bHZ
g(+-M18NNbG2f.-HFB>E<LaN&\Z/D@@#_:6^H7#Y\aJ4.AW,,;]59A0&-(5+,5af
]?CDac[a)_=MHMd([cNbA(YAE/a/RfCcZY0;HTaQg,H#2PPREeg4FAeH)\I<A^f=
=S3>cRP4,D?E((\Lbd+LbScEbL;<0\&G^SO7fF_EaBWZ:5<T#?K).3\8(<71/B[b
AL7;d/=b13KWB5@KOZ)V/,69Cc,PUd+WKQNCaO=b13\=^VIB+I?WQNdP@HXIR+P9
[?8V1XUS:LM]UKB2S8AK@BCMQCTbO;D\9?8O1T<8>H[/;WDB;MW/;NB+T0U#>&I=
&cP?@@Eb\0c/Id8e_(2UVM<9O+]CGGIIXAab,GL#)Oe9R,ZX@[)>?g(^K[F@O5O\
b_=&-Qf#;QSXMG#A>,e:\D6/[JY-J9b.@bFHC3V.-[]_5g4H?ZeeJ.:fPKg.YFaS
(FE<3[:8QSc/W0+^K=(4M.LIHW)2M?DK=1)?YFXXF3K1(;ac:[T^LL2bg;)-5G1^
:UZ<,(f]\KV4W,bb[<-&&ORF]AA2^_RM7c:[L)^C6]#52<5e2-[B;?3NI(763#Y\
;C=COgaNMGGYIa/Y+SNGFL)B(=2B:.-Q\MA.]6a>Fd@,4.[0<9A14SW-/OH;Cec7
=CQaM&bLe60C]/\A=0<)A[L&/^bac.+e3=D2H.F?XQC:N=6N0Vd.+3RM8(J,S?Tf
0bU14H-d?Gb@IC#^)[WG+9gZVa3(ZJ/I#8,:XK9/HJWK+B=Q<&ARKD\0B9,#UJ1O
0bSE^5[BGZ84#aWPE1&9>T\5Lb:49gZ-08U]fP^U;;BA,8K7aXWHf(H\W=Jc:FKX
,g\U@S_-_P@QcTO2]G<P>_)c.5&N>/1-YA478:a2)GZ;XL^-Q)\O(:0WHO_LU#f7
W^O^<T-)5J0]KV2/HGC.:JaB,?^=Z&\.<Pc03VX3N76ZQJ)HZ&=^V?b4:NI]J755
g^.2\XbaGQ#-:E\#>]E?Z/S1&ITB084a@&7Lc4V6I,BcUEPZD3;XC(DaSdF#GOf2
3D4ITQ;>[L]WDX(#K?E0&&Bag?X0OD,fdgbB5dV71._PJE-VMIALPK+_?ZSU(U#[
V7Pd-g9[E@dZ#dG6#BFgCcdT3[DfPQ90T4CNR9:X&A=+3#(TR6[N\HF[_SfIQI8@
WCcC(.=<fG0CBgAL:[1d3=4+34f2[P19#)a9d^;PW/fNVVM]C=J^_BH2<E\5E@\B
W,;6A_<+1#f=g?fLS+VLJX4bF(:FY4)>B9_#C&dbIXC+\/4c0/5#b/&J46WS-?4f
f=e+b<a<:MTOI_<XKPS3D&6c[<NJP_NbJf\I4M0,CgVEF#91QR3eG)9MT.8J?/(&
\M,1GNIZM4MA:7b/TR&bK/Ae3b?Wc1C0GgFZ\[bCgJcQEC-3UJ3N\R?-92[fDKCD
SFX+4>:+T-S\]C0<#6HU3B4ggCZ3FFRRY;JdH^I]UTBadM=C0,#,5]d6@O<O(T;F
Cg&EbC:]T>E1]CL6?4SSEg(fDgbcTGP0LV]a>8TK2/]SOE@UfTGeBF+6J-K3gN]g
BF3)_OSB5LeU&e<\RB6-aaY@Wf+V(]J4R0,#QR=&X:BRdF<;)ZPC5#K5>5b&D7_#
?dC15?C7NCF+_-+JQ;NFD381F-Pe7VIN+??.30-eV,SE=g6ZT3I57b>4b:E>fA-F
L@E,fH\/@LbW-49ZO:)_3>YfE#/(BKCJFABLN?PQ@2BP?@5O0BeI,W>G14NR_;R&
VO;92S]GfIT[=IE)a-7QU:L[IBXY(dHE6,64^P9IX6b1\U>X+fHM.)g2RU,/eS3g
f4@,[E)3Ce#U_1OM[#BM9-Of]D86XA5PZ,O558:YW02P_Yb(DZ-R3<gM;c9-?d?C
Jd[UJBa-Yg-a6Gc=.a?aW4CN3_&V)16e.^cdN3_XGV1.JJ9MGRZ6#VJMSb9B+DDF
71(e,ZS\afaJEg6G#H54E=U8>e2Z2UN_b+9VR/cg\.[6K:Q.XRGV/:48#BFI,f3P
?WBZI.K+GPZNg.X:]K?W^Q=8A>M)=ZV<G@+5UE]X<U1df7fCWRcJ\f1L_KV2QY&R
WLdB-2cB>I&=SbQWS<L(O:)RHC:7EM@d7[D^d.5/K@WBd>G+[)C1TFD[PgeSg+Y=
)26Q6S01^OCK)R3d[+)e5Y45[/Q.QXf2U7B0aQ4IT.P=3=^]@#O:gRGC=@P-P<Y^
g?([C4:W\9BeWc/>)g=Z1Ca5Qb,53-VNI;@[g[+YeP++)7@Bbg]#RUfN?2DVbK7T
\K,@-L87/53IH5ZMPN[^:LDO]H,Zcf/EV1V=e(b)_BGKM9MMUELeSe\;EKS>;,:Q
E>]fcQNFcR@MdPLFAVUaWV7@eB7IFGM@,Y[9G9,#[+4>BBd5VAbK^-/fT[+QJcLS
><@SHa0>QfWD9B#gfH;^2I//(0PEO-_4[CXg5OOKca9>M)?,QW)PJ^dfI;fA,7f/
B:)e3)db&R;)#<ad0Tc1DTA9Z7^9@@(?,HcRD97<c6BA;ZDIEGZK-T7[&.5J>RgK
a=-4Waea[[Sc-F2AJ3G_:05Ma;]S<[=I]-L<+WQ-4-@?\N[:?.A8>CcNCEb(>C9e
MYVQJ.7#(@bJRbT>2N5N>\cF=d67.TCcbN(0#LHC:R^>2KD\5O(ZQ<>HI9W.<;8]
1I3QTDdRY>-V/_;]#QO)5FC2C5RD\78YF:;MXL\g2=5?&7aJZ/YcQ/YL7RIRUZe.
\3F?^8W<?B=A4\IPeJ^^9:d4T>E9d9Q\;PT=1QG:#)-Q,C13JL,4Q3;9JQBA+-R&
SOSAV\\IbJ=E_,fLdNH>]N8;,A8QI.#IRU.)eZZA2RH]1OCEWW;2,cP4.QO7/1BG
)8]X7@MSC[?bM&\c<(7cKDcJ--Zb.?8-O<QYJ)P=OYgF8DC])QE3g)I&D_1:2NZ&
+21EB9?F:+E@91gdaQ/8Id1fS,gIP6RaIc@Q)(2_1[=]:#C,K,@V48Sb0W??XW&O
DgT(B&If&0\XF;@=EVcg6\RQ?J7Lg,7N9/KKaJcg8UA@a(I^d?HLSf70WV3]b55^
GfY84,WN)aK[8cgB=3I]:\D4V7;]_<VF.R=RKbPO82K-B0WS]N;\F&fX@W(8e-7,
N=&S]A5M=@LYHY77;b+:G-&RPc7&PY2[g[FZERSZ4A+&UE2:AG7D9#5W3fKHSONV
<[P3d+&S>G_eI;P)[L00E:3A[aY)fI+X;A,J4O1<,;H@>IBbUISS+69.?4fdg>g2
YV#aFV8R^f<)N=QHQI;12U,+;?,c@<7Q4O>G0[-F^S1@JTF@UPg(.(Na986BEZ[>
=)X:-UW5BD4,-]e>>2cEZAWZKWc_0NW.6<156SM59J:^E_;_Q3N3T3f6a13BR4<e
M\HE[f?XT3B\<:6+fe1e30W\IO7+]IU#6S4V4K#;3RU-W]B1gAQ348^bZ3LC0aTd
P=8eaY+R,QGaBP0>:cAU[@]bMZd7<&BMdS2>./b[Ja+:&gSDP]MgC]DYe5[)0W,D
<GJC=W1:8IeP847,eWRMA.JP=_;d7L3C[49XP_e,;SX;g037&9L]E_2@I,Ed.R4V
=F:X[@+<.Z4P.>E&)gJPR&US6>ZWYZ_4WLP:K0(Sd=9EBW)[/>G=-b:X:B;.PfVY
IMEfJOXZ2MV=63_dA-TdC0.1/5)S<4HAJO.eD2\M5c3#(/6&acS2,@USK:e:X?,X
f7BU>&J5gdDDZ//H?F:IaL1,SDDU?egJ)7G6X#gSL=+]C2BP/L?4MbG9dI^0gCJO
/TX<F(3eH<cP0DV^f,A4EScM3YCM43Yd#4/C-51Y-f=N-/.LBgR1g-ZZc@I3U6@O
-Y:4:U^a\O,&G92PEOP_2+5S=9O-M=QaA.Gg)94K8c7K+8.3\4FVW^GGZCB#Pd_0
6R=KJb;<Ud-c^I]?9W&:53B?/)0((L.&Vf6_(P(G0RD6Gf1.-#3#CS2]:ZIQLNJ)
a3F^3+QM?DXU2]0R9a>NBJ:2YJ-XHe#EI=(/4J__VY&/(<^d\C^K,Gc,e/8Je^.P
?]BDX24Z7+^J0S51=7M+[H[?7^=(,IS\;_M(1d_FPc\]MYJ;FJZE8[;9>W_=LJ^J
CHJLfIE5<;g&?D\<^7_8<KTUWgG-.+NZ^)V1A]>=3@(4X7/Z;UECXW2Jfd6ZQQ\F
HHXc:@C,S9W6>RQa\.>I.gU(I\W5Z_GW,M9GRfO.C[:IVUgBbE,Uc;I^\_OW,Ra8
Cg[U-6UO6</O=CYG^EP</0][O6E/bXR[J=.H+gb#,OBG&S(XYK>6EUHOegC#SdV=
>D6c[;K4?1@/XX?S[FZQWTa5Z5NA#EPABafa6\QQ?<5<6W5X8C15DF.1XK^,:H)X
aLL=SU(?ZL=7J6_5gf:9_4a+ZGJHLZ08.N\-]aSZ>P,(JM\=)RW\\RXV4(\-7Z/Q
)gVO/2B>(SV+](W+7BMYJ31GA2fFR_gUOD<W=KI.g>ZGeR\MVe^=YJ_6WFZ7Lb2^
[>[M#IK^>8O2CSW=)Z-US@U[198A&L76KL+&aO&8G6\&PKb#BR#VU)IUZc/73&:]
d&SLMe9Rb6R3c=,TUTU>9-J_<BP3bGRUFBKD05M_I,8A<(NBEAQa-4Z)<E)HTR2F
C@11<,\S.6,@&)f@4@f6I4WJgG3N&\72??2>AW96acU3ZC3d;4I<DU7TPRH1A=T/
EQD1=&.C_38?[8A:P;&J?d<#D9J<NPZ/7X#PN#]3,&LQb6HWH#1M\,3gD8CdOHUO
<c;&Y-c7e+//&#4BdWJ^;Ta28^1c@L6J)_H6SF))>Y=[,T+J5;@LgV/A9,FG#XRY
EX>QM>N1,aX1CIRGI&Z^-R0OFB6G=+_YEF_[F,TJ1>JA2O-.(IINQ)7H)^_8-(J7
(QB]7_dP#7P-MP\Oa+-9N/g;&AL8f;NFg.YA+,]):ZWb(3c1dcAJ-ETBSfX[N+00
=8M&;8JNA./5->672MTS3]bMU0?MDZ33RWbVTCM=EXP&0[Mg#?E9:ZE#8OeN;aSP
DTAUUYe;gSWTS-O;MS<X;W<,]Wd]YIIX5L.ZcTV?Lg81K4U3[.TJ-)(2H;V#?/.:
P7@UG=b6A=69ACI>g8@NNWOU24\O1>.fM\T^/D+/CNHK.M+OP=\_D^;;29Y1,-Ff
D8?O;A:6HOTS]b?OXCe&Z=>41HA8ARO@E^^+V=S.V-YQ.5<D02BCNCKCMD0O:Ubd
JEN;E-#(,45\_aOPE=LAFJa(0SOFH,3:F(bXB>1[0^N@6b&ZRK.E;a4(fZ)BIWO[
cR3C]7F-KZB-JDN(E_QKL\gQZ,ZJ4RK9QT?cbRB+^XLUE1+?_2)4:TaBZ#>IG1(/
GU(E1.C-B(-aZD&de:P.;HH@NaKO+A1?0650I)^dB>K20?Ig/;-GF^_-eY,d5A?X
.-(NFD\D#Z(<PP9XLO\Y?\^8ge@=S]8=]T+Rcb2[XdgUKc]KZf=UL_.IgM2A^dUI
F424)a7b@5]F_cZ2VI>Z,89&^?)>;\J,;=VI=>AC0Z??cCf\=_PMZG_)K70SEf>D
WIMN059V]b&:HV.SQ/G7K5d+9;+OYD#@3>[[9&[U]EP21f;X[FD#6F;)e18+Ta5]
5F\G)g39Yc9?Pe#X(c(Ja>ILGbV<H^H2P,UU.9_[K>8:[=^2:VB^\HOQ2a-KDDHT
/eRAD<T:,7->+/A];:]5fZ.K6)VD+JYM3EB(6Sf2:cV[?fXZ.PCa(@B2+]]:IW3Z
B5V-?ScRI>0HX<Je\2+9;FIJPeF6<DIQKC[gCK0XO):5R#>OgJ<&U.aWgF>IF1[R
aTX>=JIb7^TL]W?1_#9f@D@0++U94-J@QEDd]JRH0G9+Z+JUc5ge,IBH&/Ce/J64
V;-T<aVNRHY;JNYO@1TLEIK2R97gJGF-X#&=UHYX^6ggZ@X6P[d1,GC_He483C0&
<R->e0_B,LM1DaV9QRS4(ZI=>Sc>/P+P;#+:Q8K#YRK3F;+Z&>X65C>X5/ELe&G.
fMNX)ge9OE#?AUBg/G[8U+]+CD=&W56^6KV9gE:AaR7KY(C>SC_O=-gU4[Q,0OeD
8@2M/@28DAG4]EeS5;^)=X1FL0B\T0QCOBa5[Q+@T#5/:4[WJ5G05_P6;LUOKV=#
W1\Q4cFWFY.ZR&QK2@C_gRb@/ZCBT3>]SU3aNQd+G?LTC,DE3c6MI/ZQa3Y26_G+
F(<S^bX6Y]SEc/OF_4e5:RYT[1PQI99J6GBb2GTPFMbXB]aF.4W?K>@bQBeAg\V8
c.M>>8gKRBRAB)fc@./a:-F_]3M?[73+4/g[)YZOZaJXD$
`endprotected


`protected
H0)9:Q9QW<:8gNGQYa)OR]eK0^&DfS5-8ORQ)KN21^WZI(PR9Gd40)X^(.R^ETF[
&P5cTP57Z[OaW:&WA\d]B_eK3$
`endprotected

//vcs_lic_vip_protect
  `protected
;g4_^?U5C_]S#?19&IgJ5)G<P[SF51.6Mf3#C\^>gN=0AW-d=<f>-(]B0?=@K#>_
:EBT/Ka+-dF^Y=QVU)ETTcDRAfQ)E81gfCSDT)\)]PGd]3aH-90<>?)OK>IT;J80
ORX9S-0K:PeB4d#AP;Ae:VWL06g6NcAUHEROR)8;eE]fFJLB791@>8]@TFaa0:X6
<AaCZ6LQHK86@X\N50YG3I9Z0?+JcA\e.N4B+=#5@>V/ESeNMM#K1)#,G;6)RR0)
aO8\YWVVG/HX9Tb,3g9-O@B#\[dO)NF/\gO.CAc+ZPaDfR>_L95K.;P[dU+>^_\a
HeTYJJF,.)HHFJR<-;75K8R&7P0N1bDZ=<LQ2__L/KYCOB3YGCF3/?AaP,4Z/L(D
C:0/YW(I(6YbVH-G=/4:g@L7YR=Zf]UfHG<Hgd;[G]b\V+eRT0eX>SfEBYNdV].U
?(8X<A))Tdbd>R]QS9e2c-efc@-J<C-;6a94a/L\g9)HfLYQ@Y,5-4)UY1Q7N=dN
?4HgWT/1YM(N8bd#FH+=->I&D496SD-C1a#;@ON\JV?aG,\60&5L=fE0fWV^4CJM
G:LD?DD-MGU#>c=I7F1,ON@=C0_:V#56(OAHDB1&F,5Jd7@CWB2^4bPWH,+RF2Z+
8f1BH9Hb7(+QSKACI;2Fefc,9aJ:Z<#LJ+2TSM0U,[3995Z_J4,+OO98T9(2W))K
5Db1FVE]3E6++<Db;2&/16:06>Z,KABI?I[:bR2:d_M1Y,g+e)ZPQ^e+;.c960ag
6gBS(Sgf(DaMPKC]#@BDXTIWFN+<8-O]#^?=N(fg_Qf,A<a=:YHb0;/]R247E?2b
73>:_Y4GL]\^4Q\V28A(Q4C9U>@T-=U]eS+^8LV7/.Zb7>3a>,3P<<;/UgV+GF^5
XMf)cC0D-&31]AU(-NPf2MS52gZ0LPPdG@D,ad:1W>2LHfZU8#GOQCGE\Na7H@_W
bT\W&<I[=)7XIH6P/G;D#-6TD^O)A/1S>Y^8[E=#FE4KH)?Pc_?5_9a3_N4K1J8I
+H-6:)<>FQZ5?P8-[4(H=]&RZA77g6\#:>X^L,eZ+C(DPb>JRAR&,)4HH,G4AJ\e
H4e05[L>HGP43>1N\\32[\G=ELIEV-)TEg]=e,DMHC4(-)Da=Ufg<X]CH(I5MWDC
Md5;Z5Z:UMW.L^=1D&M,OGG6[Y3/FOO/6)I1<gAU8dB-Y]Ug9QV?<AG;MI-J+./1
]>3bS[\VY\AbVMA8,QYFTO(WC(<FM#>G)<.CC0M4cI<2<[?9[5CTKX-/:<O6KXd;
M1T;Y4[R\5OG#\84.a_(&gfFF86OIcC_0/NO)[4b-=:Z+@1.C_X#20E57+&#@\.(
Ya2Z4_:a]DRSd7YJ93[W?(EA[R0Jf;^2/Q+d,H7^a&8;F>L#aYP47H<Fe>6W&_(2
Va[:HPc;-Og6F<UV\P;2fR3\-48PY4cW)[,(HAC\CAD.(@CCNVUQISeKU?OOQGTF
U:9S&TG&A1dTIQ#^(B+)d^CQ9@EN)07S:8?0,cSGg;?#10\28I)Y0Y3bg\TNVJ/+
H7=ZcaG?M0e77WM18OEf=FTBN9g[TVLcD&]N>+KLMAYV(G@^@F^Ec-Q<U588X-RU
gV#XO?;ISR>7IdR:e;K<K6U(7EA[O?MV864f.-V?Lf23T2;<#=;/79bM;02M1Sgd
FX&P]cX8C<f9PAT?YdE1U+Y?1OBda?aT49U>@eBA+@Y:(PVDFM9=&Q2PUDfS0a.M
(2R=DM;K9/OG?M15?M1,9]-cDOO._85DeP_C:.cDK80US2^Gb(B@JZ.72]A/+5IZ
^TEA#ABCX7_^Bb5]L6+8:9&(X@#0B@=(1QLb(&)HNGX86]DCE)MY:=FNIeGQZ-:F
a,V13]&]_eK.AR;I)2fRa4->g+J,P9>-(XAVX7bI>ZC;--[18SGR-b<Uf6?aR>FL
ELY&EPNHU7O88D/O;P_Z,Q/BGH?5M:FUQ=W4KU^.V?(f+]4X5W2];>38<^V0[FBQ
UF\X&CT^.7TBL0@Q+If<ZBbYCgM=@ggC2OPXL#CI8RBTRdI<+:4Q36&#&7(Z99\3
:>2+1A-\EQY@?)L48&1B];V<3FOMDD\aMWS6A/E#BOd5.8-=XRUeE6UDH7/E+Q2M
OfR3--@26T9T2>\[^FL5[)E8:_1<:49;((9,LU\LV6K,f.JfDTdR+<6JTL,IY/G9
.M5+9:UA=a;EP@E#Rb[)cANHA?(943X.SP[UgJ?gZRKD?a6[P@S1H2RPP7EM,[K<
C,/3Y0J2C+-6:<S4OG5#RJNST3bLX<M:F?e;6fcBP.A+FC/EM_cAPQ0F83ZC_&_/
MX^L;L0OIKS2FQcCK9KHJg>Z[eR-CG5H.8^EW,e_4UHe;0GAP_JN/.QD7_-.0/UT
U)Y03T@S\cI6YJMHLZXe0N@6#I^X/NG-J0_5)@NCb)a8SMH-K@VFV#G<Z_JVaV:-
T\cIJ<TDKgDWIZ9?\@,;68EWU&W?2DdH7\;48C;J0M_?B8>3c(-Y=YA,QB&BD@dQ
9:g]I0c)5U.--@LbF^2Qa,c&13YRYM(TA97R@2)^/)A_,I;0T#;d6<_A[F0dN(S_
EV@6NXP4+Z1WCR.BDeCa;&c++d(Y2C42E3OF?BAF6a(FaD>;8E1J84b>CP#S)GWW
W9(G=R0AVDd8B7Y80^&Y(S08U(N7961YPEALcK7/H@G^SAafeT=ZW9C<4HV(0OdD
^WB0@UVd#-,>aI@>dcK?-d7)2B9M._)Na3G)2cA\GRP[]^P#JK4M;YSP-,C6eP9Q
;=a&OW+=(D;Ac-9,-^2ZE?G(GaP/X=Z^VYE5B=eO]PCUDCT)_[MZYf;G6FJDZQeL
Rg)+B-ZG6_1F?;eS:F3?;/2T/8,X:9Eb+^a:>6SUa/GU/XJ:THB9XAF-V;C<[^0T
U=8#(dD)WMZ<EP?\K-BdScX+/S\9^+GT:\PGec+@)/(\JT>C.d-7D15XL=K:J@L?
9PH3]eL4CD;7M_7&BG=aWXKE,X+b-C?]?-JO_D3=?TK].@.fZI]M=4+8^+dG_AaK
7Y,[BCG;].<=@XCcfVD]^X^F0Ea,;O>;C9+G05g.b35S2F5#>3Y)F6Y3L.N>I::S
d)^<.CVc/64RQ70[3J9e2?Jg27W287@WO@b>]QYdbMf5GUL]aHA8COI1^FAJ)8PV
G2bKY&\<;?X)RYX@O5;YdNRRG@&.KAO^M^]B[OL9&C5[0IaUA:L)-9cN(O-BXE&f
#SW)IFd/E_W^M</^Z^.]be2[Ld#V))b7aA^NO)dVWHcc/f\(-PJ>8061DZ26][2c
c(E.S7P<]7E_bKT<L^IPJ,H8e+^^S-<O#BJA9P]e_]235)9)L)]d,V@_(@FBd[EQ
CW7/9I;MMD/K]a.80Q4;Q&>-][5KJG.(/L,J/aXKT,M<4YfT@C_Y#_N4K07\D4fd
+gH:Y55eQ=FTBTSAD3:aJYN@4+1Bge:5cL4<V8=PCKC_?ILIcH3RHa:=:INc>849
K3><(\G?>C\&aGM.5T9I/#W&8\[b4fcg@K-b5,5F.Ae&eC#[FSN7)VQ.V?3bKfJC
17XE>U4U9(cW2&1,)_,]I2gfaR1c+3D<9-8@@W1bbgg;0TC,L9-@JX79NFC>A=Z3
f<5Lf)X?,]^W3W/(BK()@=d[-MFf><)eJfG<)V6Y,0&;bP4A#9D9/<8\W)_MV0VC
H^[+W;DP27H4^M<IQHY@3KQ#)#0bZGJf[^8W6@:3+HUCV2F_gg=Q]\8^5&24Y6Z&
5O;M#XP2gHdQLOR6)-B[ZIGdSg8B/3B&,6[Rd,RN@T+KDeE;XaNTCC<gG&_HZ#+(
L398Y>U(gF]#S0M&?=\8^.Q)#Ud/]ZF(TTA2JXSR1\CQB:IBF@:<\<.-N0+ZB86R
8<KQBPX0Z\RGP-@c;6,&1]IT?](\9_&.PJ-;PY9:d2>VXcD;SWWY4H;7&0KJFIcT
JQ:[R=[7=NG?#4R5Q4P@&2Z=WDQL@N#YZcg:GJLRg-c^-KVDB_CSK9c.H=?dU3]M
#S\M(@Rb;;UE)]AWH^9NRY2?=?AY5BYXaWW2QS?S)XB:RdDTc75CHSK3KRD/S\=+
.CedYaKLG:8HS<MB2(LWa1X9H0(<eEAe5ZX=3E(4YTE9:PT1c^.7e3;3)(>4GT8#
5BWV2:#&HD)Z15^2F#H4N=a[P>If@-^16@XD;Ld-2XRTHgf-N-TeKT_Y:<3QKH\,
Q#N=1YBg.FD,c#GE@03]eP->X]K:23IZ?70HI(M^SU/YRTc<M04MOb2[SH_Ye>2a
(GFf):?@I>?Y=KC1[H#W_#D2OG5U2EV6AEYJYc_<O^_:#_86+GE[/^>V;@?7]SHC
)FE\4BT(;T-)_P#X^,#V(T]=)V_^ZM4=@IW220ed[2:6bQd=fZN+e?c?YY4<1g/c
TI:-QDR:Gf-=>SV3+dK/4R>KO3J(OP+O/3Ig1ZR1e^9ADRf[[f96:D&U,.bV1.3Q
8e1[(FD^gD;a5Nb@?PKE6@E2:/O3WT>BT[.f=V>ZBP5aI(YR?9UQc?eOX/&gCc1]
/L_)5<7:6BGA@=,FZM<^eJX:H\?7:C0-S4B/;P_BWE,E77,e8F#^Mf<#_<(#,#,8
F^OZDP-/1JK@N7^b(0J>#b:a8+Y81_c92K^UU[GIN-\SU2>5V@../X]2K5PWH)\Q
GDYEaGO=YKJ.1=NcYF.>MQF^cK.)I43I>W5(;1+Ub=/3&9M#H7#M#O>JH6QW)X_@
/=;Bb_g<Pea:)4IWIC-2XDCb@;[FfQ?8Z?RJ.8BIYY.V_DH0&YBGc=Bb:8aC)(S+
4>I,FY:;^793cAgb]2aB(BTD;@\/@DYA&58gZ^12[T_/8NZGGbU3G-N[);e<0/YB
=Q+^Y0F@GB9)RT_::?XVUd]@][AJ9B.N?[9d9I^99aBLaO=O=T>5):5V<GPXX@e@
A<Z9_EMLOCCKf@8cVM9RL<&+D&=_R(b-Z^6#Fb?]8UHDM[XTFg+EKc#ESb55IcRD
YI>3F?X_M77\g(W/;FN]76:_cT5HX?>3C2C[>P_8].LE6DW?STLc.,RKd88d6(JL
#M&\SM?f-eSN54D7Q;C-N+Kf]ZC?<;\185EQ,MUR=NfWQO7J:T1?QA2T.VYc-)aW
1JBF-GV2VDYI^?N/)c7MKV/3e-M#8db@[@Qe?:d.Q[2GcZ1L#5\;@MB/X)+4@P:K
^Ib</QN##]SeSWU@Z#84E=<&AAbW/_916d;](P\S6YTJ<5=I-XQYQ.#.KaA2f50Z
_&8[eN4JYUD7g9DH6^IdD-fgB_?BPK,OR2L,P,?WG3#57Q&Wb#Y?8\XdQa]W^]GN
&3#<Q_]0]f]4PM=WV8=eKO137DIT;,M#6b<8#f]]cM=?bE?+cW_b,X#2[R?a-G_4
TH.91&A]YNZZPHF&^G&d<QE2Pc+0M.b?02CFNCG[\,6FZGJLf0fKWf\gZ>6[NfM7
[N:M_7T3g&BbIabSFM9_>P0f[^IK#WcZ3aF7UZgO-8aA8OG7:_&IPe8<Q#X9Z[U/
LBZ]B:g>(2N@CAL5<QCGUXK\XH3)4P:DdZZ=(:05_AUf<@BK>gLUfbZgDTTGM._(
&a+b:8OP]b0L>G;0N<S4>[a@eTC]f0/Q,I:d91EP^HV3)(7NY+;\PSXTL&>0S[aA
7NTbfDUW>HV=XJ_WS3L^d<8gI1:0fMNM,L3_TD/X419>TJg2#W:FbJ^+:(LRTeeS
Sebb(IO#7:EdWe<)H+RX)6;&3Y5^A6YZgM)]&R>5QF+AGN(E.TeCU@.6G+d)2IK=
fVTaO]cTTdYP&W[F6B>>T>bA\cGE#7:DA6T0g5X(R\J(HHPSDO(N,?EFV=E[2U#H
\D\N^FaR:Y57c)\[I8TYLe/FYYfR_Q\IG+\#2/8SAFJ@EBJV0W=bEPaK^GJg)f2E
EAHSO6a/<5CdP<CN,dIX\D/F5$
`endprotected

`protected
OT,^/)VA,-F\9W+R>-PVNW&E,AEcfQJWg+a,YCYBE:Ue[5?-:^,K.)5+Cb9SNP(U
=P)>QJPV\\6\0$
`endprotected

//vcs_lic_vip_protect
  `protected
H9f5^J=+17QMFZG>;3Z::TMa:F&?[G:K9J3\#5[\da_e?dHCC,#=&(=W=PHHVb3-
R[;&-OCc2HVA[f+I1M0K+<(8@a;ZK+8AO-B^I1Oe5e30<>@Y&WD)RTUCXOIB1OND
Z[4=@eWHNTD=[6S,H]=cAbdA;A;\MZ.)?69?.&1Q,\>T&XG;S/d?]5<_KC\8ZQI_
V;&8(YP/2R@5T&R9Tbeb7e@A-?>>/[e_HC12]ff_H6XH3f.g_27G[0M3@@gEbQ?4
BGac0M6&b7]^C7<cU1^.SOCL_&MIXdL=9#F18RaJP4HAg8OMc(ER@DOcU]7e]TE-
9>R@]D@+K6F.#BEM^A^eV]0&F5cG@Be+NTa^Z#?eK(KW:21EX)?aKa-MNJXUUH7W
&Z]<bf:0FP_@1,OCC8OYL4_1<#82LU6/?XfSY)<6gB4;2T;6#@1>Ca2)4Z#M]>0Y
@AMBaF3ZO=0I@,P6U(:5aO5:JY>VC=]0(4:6[/1(_O_\fQO1^YSW48,I4C]2cfJX
H:LD372@F:1e\Z\K]d4<Y^QP-VM8-(QD.9?Mc+A-67CH?7<.(5-&6CC3I:FA88_\
2f1^;]I-e90aF0^<cSe3\H,TZV-6E7P[=bc<H3-W+])<Rgb.O?W2AL.=/ISC&b7B
f@c;aY^]?.RTG4F2BJVVc20)(90bCEb-f3#?a3LPOeKZ:ePK2QA@-63])T51A4B=
E,=9?6KXY+PL-,4+gWWL<JEP[U;T/1KQKVD[L<:\fS/^<3<ABXI42dYeg<9,@HC[
<TI5F@-NCM<D.MA7?BB13XfX3?OfZ@7bIV9#f:<a6D8-F^/afAg,\,V-=U[?^S1=
<:?M<.F..0d>UT9BYIVJ,YP@@S&(Ua=_e\\+9a4O+D4YMYePG>0K#]+//.N4(=/V
,bR3YSDE;DAeNSg<S(P,K8SP0-<>8JW:3)RYBH9C]M(f2[WN.0BPY1g;G4Jb&?MM
G2M-8]HU>_IS:b3I-6bRFC[@UgeFfD[Y8((^Md>6cg>cP,S4-MC?c5N85KXUZ2[U
F;AgN@Q@RI;J8]KPZCQG#P3+Nc?&<B8A8EL_AQ-fL[?][>GeN3GN@L>K,[b8@AM8
-C;K=d.+[N-4e[E,HC<7W4V9dZ-M3bW[c>e/AZFf^QB_J7+LNQ.X2]4bGGGBGRL6
?SS^f0+OV-Db9_;Y;68Jf,DdAMdY1Q.7bYBe+db7)YMI#;g-L4-f>S+I2)J:3gM2
+(fb#KH-]9=8aO.BTWJe(5Ba?L11,N40a)O19;8G7+Df9AK7\AIc@E@6d;XL?5;S
-RC50/)R9HD[F&UeBJ&4?7F_O,6EQA<I[1Yb\;g1@QdN-1MLcbaSZd+/Hd)V)@7P
=g&_B]B^R&aA10K)U(1BP,=K-R=G0R=c87V5D&]4KJJ?\(+KHJ8f7(,1+(FX^Ob3
6#IX:GfDGcPO8^L8-AFaBdT(/9H7W,0I,W<R(38Ua&O/A5CQ;Ra=Q#SF8[9.<(O#
BcMOP?NJAIQ2R3Wa4JDc/:\;5Y4&5ZK1ONNSQ6CK5EP.ARCK1)T+ZD;c;.@U)D,[
_F/50Z,TD3_g;#fT2QeDeC&g_NQ?JaU^#2L#HQQ?:7gG?:DfX/-I[PNCWE]&2/1X
,[^(H>^\6/XbV,XB<9+9fEK@D\db5,&R=_3A<QCD<&N+Y^Xb;Dc3R#Y+7@H/?8M;
D4F[9eIFBgS-_<#150eIf-BK^c28,;J&72]I&1/64NVLK]a\]6&5#OcJ:^-;V\.[
,G?ILDBH=fN8b6D?\Z8QN9?+65P#+X:gb<gI&IS7c&SKY,E7B#\P>LU659.+NFGR
\acB.abR)84YS4a+WGZ5a#Z3cf5@.LD:T&EfD,)4CIYEQ?MScII]WD<fXI/\f=S-
VS[6Tb:]Of>0G9T;W^J(&?ALBc2Yb^.-A?gZg(>ZYX<CKO4;^PZ(\NN>B8PT64HC
<JbN#D?]ISJ1;8SOVWY0\H+N]e24>1\<7<b\I]=A562(fXHF?)-gMGbf?^4+W77L
0&MC^a9ObcML&@9EC9N^;AU</WZ/)<.g^\b#/]d[Y]-B?W\Ka@Y+_A^<RKH-^-VD
g4GY(VaB<,LU,[H.e#C_3(]#Tc.AH198LQ0HS7)A0OP4\TAdN8@M<3fCJQ5I8Ta4
gDSM1HJ^=Y,T7C\NMZ.WKf<aI._FU:B?K,)72RA;W@CEQ?:?6(?S7TXQ6NHQ_2f7
K:IA:S0cHDV6Ug118E]ESScSR_?2P-[7TPDI5I,U&F9YHTJFUQL-U2J-GTUS06TF
BBX8KJ.7H1D2Od+R9HE=:21D9C/7&W19K9MM[P)S-;\JMe/KMa7e>VJWX7YW9KD5
MbQ[S7;F,C]CbPaV_cAdIKbX.A;T;NF@27;P054&FY:GO\B=WW8b,0>KJ@[=BR+>
5J3>&<EU&.<6)WPMVCV^g\BL8<=-bUC^cAQ>#:6b?dN9PZdFZLAFRSNIVdA^F2I9
4@XOT(MS&Rd).#,Ae9#b#c\g-ZLET+C5#M28acf]8]A/8IPdI/cRD<#=ONZAK-=g
T#[aKA@84TS4FdJG7HBK;9Yc<E.)ebRX.e(]LHdNe4b@NV^GTc_-2?]YGQVe\72d
g?WH@3Y_F@a7H\ZCQ0RCQ5N?7O29#XRK__eaJ/>IZB_L<ABd3ASY536:(^G8@Da,
gN/+19]Y5IN)W^Z)F=(,XO#N\H5IVg#f75V-RG?0WU1&C7+(=Q,8R,b3P?NWB6E;
A=HE8_:fcF>4D1W6&[N&<WBSb1@RCQK=C:0GdF/1S&BOI/LY#.gLV+.+AO4\O>E;
/aAX7::.bXEPbZS)Uf0E?RLYgg#N@9.KgJS;R=DCRDFY3_bEPdK\S3\bVcEK9b0P
;Q_/g_P(]daeA<ACJQBST4E@+4PgRg=8>S6/58JBLdHVH7VP/EBO@JV]AcJ>;eSL
_e5DM8(ZZ=D/N:d=35bS]2HJRMG#ffd]>\@2OXL[>#HWP(=U^]A_YX5d-H.6XX56
f453fT+WNS7@?eA^G&I3CDT1=NJ(494HB^,\G,AF#];N6<,@SI[7fc9LNGKWTWV-
H02Feb:/F:0b@<,)Y_<=AV_VaPdIW]e]-A0Z,d][3E=,eR#48WHU8EWaPD(=IcgT
DMVQQ\N5.[Y9=KV,#?P6aPKdZ:51R;PF/3Y-RK2-Ye0VOK5K=CYdc;L^WU3E9AKG
#\9aHe+WQGY[A_-^0FbJ;N@Q+:UaU@9?/0?#;[[;a?5G=INJCKF7L#aaW@GY3<+&
<&EbE/aR;WP1)QUJ?e#fDTI)L9@KYe@L#:CL5MaSUa^gYN.-DE&5:La6b4Z;N[J5
5#=+4\Cb7#@\;eUGU=&@9M>J/d910Ke>3&;]]V;1<4WcUC[R43?H0f+L2aaWFXZA
2.<K\3U(eZe[:gO,J:2JKD=+0_J;=H@f9Cb8T_4PS,C8&#FJMEF<A+H1U;dH)5ES
].>KRJ8^LXH[P9>\7dNP;4b5:M<_U2/PaD&ULbI#Q:A]O+&UWK/79HRN@M#;b579
CZI1f\]71(;O)Rf[:G4[Q8/FD+#<,,f^MZ47ccTP0\STcC7V;M(G85,Z5K97+<U_
CU@SGPK/>cKUd4e7c?0^GTSE)V,3\DU,6,T9KeH.>H(AaY03Z>0;_H]37S#P>Z(]
eI(f:)aI8=@IQaN#NWP3=95]TWV(_PJ^UEYR8a.GdKR7>6<D&[RCR(eCSGfceMR8
,]B=/A0(16<@5<CP^_WR&O@E+MFD;9+ZcPMOdEE&LSA,ESgDf,]M(<[.JT0<dA1c
g6&9.+Z]@_:+Y44e3g]BBQ[15Eg(dVT<+[/A^fJ5bf=aH@F[-5;c^M?JeCYVZ)b4
g9Q<@AXFF?Vf&V-P.X/^A\AHbbf,LfFfESg0;NEN0#+g6<BB0&QS9UT]AbU<CDUJ
SI^J2/^=/7._CN]8U<\WWN2W?]f>M_74I^4(G3.Z#0OfNI9]NAbaf93Ada0\0cce
fPO,I&TR2O=VNA4WN7bQ?/aTdMcN<FJ]be;C&[5?3d@@7-F)31PIUA7\V-W36XZb
b0(dEbWYSO2b:d?)Ha@/?EJ,UKU08IQJ(ed)J:0Q0T>AbY/X-YQ<3O?b:B17Ua[A
#[c\<Jb=Y@CGKO9LIIGZTaMfSE_/+JaB_9U+88VO)7FF;d4>4=E6-)_[1bTL,g.E
P5<dVa9J/U2.2UHQ-)IcKY()1(IF,4.8f82cA<?TgaX_4^H);\K9?).PfPV.4dHf
gQF6\DN5Q>5KYI<d?7,724A9FQVL9,.eE3g&L;1X@ALMLXH>B&&8gQ3,;P,0>MWa
&1K=_O4P\VAcT0b@C<dF2D2T1@^9?c8>ESAA572b^H;\7f:d9_2[fM264P)7\Ya_
9dbY^HE80&^H1NJZf;Q4?_F(f^)31/UdUP;)8Z>>d,J[^;U6d.2JJCg>?R]/N,@0
dee<O1&RM4T80IK8@Sc\_JF,CUM3=V29I(5JH3.00Tc6=Qgd>+>A;McZG?__\gPL
;/LRMWTG<Z(a>+N@W?:/UQN8f]\DKJ7;78ROSYJDRCPK;XGH+U;+(XSM;B8M1H^[
[1MLAbF=YB484;>NNZ2-5E[\O4<0)6;c)gV+ge7#[RZdAbUcLOHU9KWd\S7AP;Ud
JGW>WX,geX/CX>Dc)D)dg/He-(c-VT;=JY[SVEGC=-)U3)(V+#OBPED5D8NHdRS2
,:)f<GcMb=(&4V8S-0L((BgD\2ALbgR)=^9SEVg>?-/]D+?;VKWMIbV4<J7D8CK8
.4V<NB3:b=>GCCT:_b]0H4-((I0AO[V0)7JQYJePbf8R;I2P/.?\UK:8?XJ(;a-B
ST,)1d)ZY0O,<c9@<OP_P4H.Q;N8d&?BN=?MO/)3U1_3Jfc^cZSF:9NV.26PF4g-
,#Q#T0Hcb6@:_UFXIQ_&WG\?d;Z=:A0/?]>+ZdfL[#I6TAC&(Ie285c>M]<660E=
]a+)3DO\40#S^Z1G6&VV;2^/Gd<-+?3]T<?EK.V:\CC4WJRL^;RT/06\=8@_CQ\W
J06DY6DHQg4MU2f4H[J03F_8_8_,[I,F@eA]g5^S+&?6@gH>MC3@O>eZ;U1->S?8
2)O8T70H-XVcaSI_^_IKf=;#2H:CY3gOb;1UQ+Jf+0YUD2C9];G=DM(gXCE&(7/&
?C5e_)PE/#LH7=)4B\0#g2JXC5?FH=C)2fI2N,,X#C7)FbJfT&Z172C:JP4_PZVX
9dI;B#P6LQ5P;J)^OgIK9ac4F;IQ+cc]8Sb0]Ug)XSNZ0YV^7M]Vb/NN^PZ>.CcM
MH(:abW5T;YJPTG2eS)UIK7?.8KQ4B2P9/J_M[(^Bf<4cSdH^O844gVN=&I#gW()
GWH^<0MeK3f?eH0NeXT&+;L8+2RV&6XW[#/NSPT9-OAJH+N?[N[+c4EcLZf30DAR
6<c&;79d@NCe9ObO:3QbA+D67YVQA<L/<X>J_7X4OKXS\Z9MX[0#B^G^E.-EKZD;
48F5>E)aTUXZ2gV:/5a5&\9^;N^VV:\TF(V&.:UGe\;W>f0KfAYB.#V@A_Mg,#^7
?4O]cR_579U^<5UbN[;&)H+[P9\QWH@MM<>FZ3^VW(f\O6M5.T;48=JKV>g+M)_+
WL6D+E@C9HB90TE&FfT7d+RdV=-a4(B<,VT_ZL]4ZEMTIS84gaW7(UWB=0;2QAHJ
6\/@3SCW+GW?0Uf3CRd0(PMNF<MGGMTJ[c2YI-#g@IP6P;3C^cca<X:)L,;.IT+.
2CCQ41PLd5_(S+b,]2=4UNeaGWTgE#J<?a?V3O[R-:ZNMS:OT7:.M5e(.CQYAMPY
<ee.GE.9^a<#KIUVF#<C0T0N<S)##D=fRe&/[SUBPAFQa?/D,Me^O(0V3YJ45Ob^
1&&CbVOCD3.bZ4]@JGC/gU1BDdge@S;2[S,3^C(A]bSa)LW;A>E459:#..7:e8?H
-CD:#5=B32@+;g6O3<X+Q7O@49@-=fQQ@M8FbTc./<:C-6Q4V[_=V2FL[T:>cUZ#
1]DP57f]dg>O31TLR\AXJRS@U8;fSEOYJ>(-JL\0K]He^e[UO6^Xg,Mgd-:.6?0-
E\MfQVgF=?A69@?<#^=0=EEI<:5#I5NgK4&Se92?WZ;.U+AN)J:_Q(JD-T9W+(:[
c-eePV560bPYHcCcHGKW0VR+B<V:AR73V97LJ>eg^,P.VT/):):#HT/Od+Y]<)U[
;0Mg?[<)P#]T4DO>MHB(972#4O#bJ#1-61+A#92W6b&2>fIb8L5GYY=Y(T4a-/LE
9QI<;Y51bGM.]Fe[MGD+K/E>(:J+2Me<,,ecMF0SE\5H0C8aCMF)F(TaI&+gY1BN
)UA\NPMeF^O>;=2=27eC-g/4;cEgfJ)U5;2#6g0UMML\f^6&P61MVD^:FLXBd+X+
UAB=G=K?-3^c/<(cg?@OYZRdf;FN,#.Hcbg#:Ecc8AHS&1\.A5UF.[03I4#ST?]+
X[df43,#Y[-EcbK2)_SN-bDN:BF.>SX8]7SJ)=aV<._Z>aI2T<JDNK[V>[51GTA+
bN4b(4.BKG?(&VB1\8K7NU2R0A:IUL]9-Ec?dI+FSK,Cg96=;QSFeQXSJ;6?N2T;
Vfd[,>#c?#BASQ(gXNJLB].N[D54GK/54.Dd;2XDQ8=4DCTJ\^>#3IY>L;553Y&F
S).X&7:c(g83VAXLL\9W@c:7/I-JA20<D3dVO=-,T]Y36P[,38BdQ]1>9F6b<7aM
4A/GX]F\JEXGWdOD:+PO0\1QI-HTJT3C^fGVB15T7T:5BB3ST0311M1,e..9;W?-
EWJfW_2A@L+eZ&J5B6K]ZG2<]1AZQ@C93f#7^;^#D2AbeWH[5/@.@@=;Q4;b#d_[
X:F(e=C7#(Y1,aTON^LEF@H5HGZP<U\TaKLG749RO;Q;>0dUKd0Ib[SJ2CQB1E+X
^RSLOR;R1g7MO(./WR^+Be4;/XEZW(7g\/ODF8,70\7Z:C(Q2/:<#Cb_VF<3e/#@
CC^.SGc7>Kab1.ZQ27TXY\BF_=fH?H]Re#W,e35VK@2F5Za&H;T=b4+c,,c^HDOH
;b_):NBAI+L<#5QdW@CKU6NJH.+?)fc=a=G>P7P,PLKOc4;:G5SN:2c6@#_O0NZ2
66;F5g@RIPXM9PPU0DY^Ne;9QZG3<IS3W<[eS=>KVe7gf#:e-HJaA4UBbU>3I+9.
dX4?/8GDR3KW8\O)NHCcU29RWcUXIAc&Z6R)6MAR.UN,22[L5<+Ga7PHSQIfA/e+
[gL>C2c-RD4<U&4I.-_PI(eFG4FRS;ZYTEde2<U/b7,73_d<.I@S?#V7#AHY^DRC
>[)SEe15#d]B@.O6gfA5ERT:[SS]])6@_OSY\b<&9]L:O4#_:?VO?6RSK&Y\aLd4
@>2ICa?d)RUCYIV^6Y&>dXF2<)-(-&[Ef7B&GS];IV3,bUE6/M<ZB/[\K<_OYU[f
EY.[0=R\GA\<6KDU9+OOK+9L-AZDg43R??MA+BCJC:Kda=>4e57>LYUK3,_=O_Af
c)-1UJPACQgQ-/J.P^Y0&_F6MT9&fd@FXLe/G(IeYWB@\;TQ+0RgNN=.G)S7V\K0
AY1O[+Qe;T,g0[W4+WAF7EF8G\dDG^GW/e&@.Re\\_2Z3K7D/VfB>_E\0adCf7-=
MWAe^RLG49GL8TK9PS-2,JX^;7fD0GaJR6,R0XS5Q>6S(C\G,0&Y2L:[Y,_PUVCb
/fSB&VAg/HS.@GJa:aM>UXWWXBaF@f;e3#)Za^3Z-TE&H0\6WFE;D-A,\+B60ONV
-Cb5RH2D[O9_RQHD&Ed-1KJ5a]93)VB-dI^Q\L=H6T-f00b(Z^5=baQgP@XMWH[0
&R:L9e)#&Y98[=f8U^2/5c9ETF;LJ>P9F_4?Z=EeeTAMXbb7?D[.#5:]Q31>YGPb
dQZKb/UX&e-I5=?0)Ac^,;-R->5)]+bBJ<DE6EBMX5.HE/<6><X=,(8&R6KLI..S
-BP7)baG\H63g4&>eTQL-1-M@A;(3E):dX?-G+>4CUA9ZH[f@8TLB=]P4XU/A=YL
BN[cAGV>.f88W[)3>8E=AbJE#EdPMfK4E(N&<fXIA_I>4bPT;bVE63?>aA6HC0<L
)&;V)WZPIdKZbOFX_c)6Y>Ha\KNb^T;@B<AY686=A=)fN12(F05S5/EHc?0Ae@JY
Z?DC;69@dO?6_B,MA;FdC<,M0TU-E_W@T\>:ADaN]G>2EUgOg&]/SQC,_/6?^#B<
LI=ZOT+LXGB[6/T+Y>6K]L+,<T:FJ/f]LE2D5Z#;T(DEXc#/0cZZ=-]2/XS)^2fQ
>:X;N5_e6^YK6K=ZK,&N07A.d:Q^ASI:G9W9S=ae[PTN5)Ld;5@(\W+<=F>SXJD#
R=3AN;5;XSC,5<U,VQ0bICSB]^-]7]X+\>[Z,&8CGCG;TFY5/4;O5FL(JQ67B&A;
Fg^b1]e=Yb&S&g3[P_/e-=OZHH@GgeUJg,0R^[)e]UT=aE/K]884?<C>V-2R<SY)
=_A;S=a<73U7;1-gP89ZEP)^N:Y+\\-b2K&bIN[BOFT]ARO9CY7FgBc,3W\YY2/_
<BM3L4&JU_[9VCf&]T&eQJV[,;&I>EJTH8#)K[B0L4;8?5^&SI=b5.T5TW&8X[@O
&5J.2576,;6bAV2(/d\ZJMC&V:Q?ZS](4:2PVXF^f+2?fbY\T]&IEQ3ICAT@ZG-#
WR@W:/CI&7,Y<.3O]?R;IgT,NNK]BXK6\M?19;]M9J-26\+d_1SfD=GdQDHC8e_=
:7BA:d?5UQ(\8UXZe^IY[42=gfW&L.d0:aIdEU=H(Lc.E+I<WCcScg0Y.\N403SS
Hg/4T-QX[,6ELVN8?L62Z;T<R(Q&WX]O#a?+_5S42Fe,1TS1\Yf,,,NRa?4K2ed7
bB[9O5C&KbVM]P1SH(7,3>^P1[64BV8H0aH?/<G]2D0&&K&)fI/-eX1?D?_8/?=E
Q?D;28.AGdZ_JS:Df=TKSPDQdAVG4<.0H4?#F-[.^(+S(7C/:^+N\I7bOYfKS0U6
5,cRR-BO,U6(>/f@RXSV(B4X6M\0E21P:XYe@Y;+gV#8V<A4E<_G<_4YZ43&QM^3
R3CW<HQaa3gCT^_34>I+O5VeQT-F4B]=bPYg+c]A?2_MKeFQ\2F0TP7c\KCW4Fb=
dG;X4/Z>7I/]ULd5(2Q4Ab/S>HfLA56ZCL<gXT8dP91bJaD-TgL7W.ZB-aK<g>2_
[9@9bI:Od^f#/P2P/J:Sa3Mf7[>FGBJY4cYK.84b)g>7]);DKeA0fHSC=XJg,5CT
EB3M#[6/>].E@[R:;ebX()C<^2>HRN/[3BO>:N3QI<9IcE2<_?E96V_G9DP-R8YQ
b5g6Tb#G6)?@MSDB\OI[;DSO\G:P&#;:S,72b(7(DMB)YE5g5;:4Bb^[7](K5GTd
gF:^PX7Kg@PO[0VLM^AUa^E[\HV\TJLO/MBef8IJ+35+>D^:PJLTKN?eKZF\+/2X
OA74f:=X):.MMG<aLEAQ#Q#Jgdc60Z\fcOGDW,L.]S1@2N.V?]W+1fU,_9bg@421
5(d(ZR^W)bW^YJc=M#V/66=J&a.XX7O<>[J4H10A,[#=W6;3bZ?I)gGV=aU>3deG
MX#)gb5^DbSO4P557)MVD&)NHa#Qad47WMIG5I+2I@WJT\N9+A^&#3K@)/R++eE3
c0f8:V-)EKABH_AYF_56dD\=KHP,BKV+44<K6:8[S>A^Gb)NSO3?S(PF&D6AGL.+
)#DS6O6.-4_LA2J_4R;BTbJ78ZR-#5bV6OFL._cgP?WgH_83dJb\)+M]MgVZPZ_=
N3e<E\>,Z<<[6d7XQOF=a(TK\G-L4JbQH.a#P:]]cX4CdB(a[,G(1DcP+M;QTO+c
BQLNL?JeM.g(<,B<--(d:bbQdXaYV55RB<#M8XdFY6T@H-VEK:1?-C2a8V00CR#9
9\2Q1C[4\Pb9N.dRA>7,f5Q(8WE1<V6:.G9)):IaFf=8(^^YebafI^)3^X,a1C>A
I0=eINKG^5^)cWF&.#7,#,VL]U28e#.MH]gE8fR<;M]?)2WGYLeR#2LQ5K5>Bf#S
<]EaQ0G-Y<f.fKRJ,.Z;&c<IW6bG#<=W+aDE8,GHES,<;E40?g:52Ua,cZV1+3L?
93HW2_;6?0e/gLA58+EO#@QXJ3F_\N)]E]:Rb(+\YSQ462VM>=)cA9CBdZX+1O&f
/6[W[_g?&&.O^]cKfL0)>=0VM^RJT9Y:^FWH[7eV(Y:F:Z]DIef(FI]=Q7NGgJA1
D2-V[0=MadZY@6J4ZFV<.M_#a(-&#XDRG3K.W61?N\>[WI]gUAH+eFLCLY],f@5b
.TV66V^Me]CP\T5\.<_[0#f><+d,&LQ0_@M[6TNP.NN5XU<a&AP\,@)BeI_<dEg1
WU1RS>MACW@^VNO4?.:OX-E(@5V&@ADeEd2eM8G8;-=HB9O_DHe@2eS]Ycb]OKM_
3cP\F7/25IT49,7VE7)@IWF>)aZ4)E@=Fe.HX<bVV94P4B4=;NB8W1_f#X_4GRX+
aGH<36S2[4M,GN&(cIB=_C.bc?@9E6+E6AaIL3L,I(JC[RL>Y<<bO]YY)HNd]A?J
AHR^+7OWbQZdZ)c\D-AQ<L.XcJ49R>eb&d@ER91O=^=<N:HFSC92S#7a?6-6P&]c
J1bZa_3;I,c912?Ne58(WPZ]AH8/7B3_QO#S:J\FHBHN40GKF6N5@)7eeK^>S<R+
/4[&Ud3P8SH)[7Md[:692LS99(R@E802_TSL_>_\[N6gYfW_A&O\(bZT)OT2GA3>
4@&-9f3cg=U)?WN6SfGYbXE[EQ/NE[gU66JT&3OWBb0=JO8EWJA+M0&&V)PC]Wbf
NHSW>3ZDNM.M,E@X=PdYKG##IdW1_B1@S5R+eV1/(9TYTO.3CM/4U4PXOJF5K,d;
CDE1.d>G&GeV.O4)<9ZB0,1+UHR]Q:L:.Mf2bY,f(NYTE;9],<,aL(EHBK,;D5f_
A)aG([#C+@c&)U.V+R<RAZW-WfKb9Ka7:;deEa<TR;:aCKDBT#SOAX@Td#dM#BXd
OA3/5>e6)Ca@_OZNc;<A15G2JN+>[RZb@c9U=dE-;1BUgAYgEIP\2<1<UbQ1Y7O)
gg>d\T.c3>V:ZZF.Kcb;0Kg)UI\ba@KP)(=C)\EC\_>bDPG1J0+a154;g2I.1[T(
V?PB[&@E0?L,4]FMb2W3G4)C#<H[<ITYL=Q?IE(:d3W[;O(W8WBA8K^>5Xab#Y\;
g#9:@=#Aa0;W0P/79IB8+Q1VDgM]?Q3S##].MT7>@+C]E@>-bD7D71DGB8/+CJ(_
KO0#>eB4U&)Acf=3BcTgM()IBP&d9P#UQ#4ZD95KGZA.+G;.(0XEcZ5Ce9_@a6dJ
A9Vg9(&ZBW\T<\XW17_\L501>Ha^N+.fL6]9KdJ@FYKdbA)VfM/8b]RbH6Z+E8>a
S21a0789W--@V2BK>ga01EYZ\OYb@[Za-_9Kd(WcMF\)::=adf<C:3.5S02D@H5#
P1Sd2B>FX^COd-HG(=99U[^WVOHc-V.0F&=F7c()W+;9_>g\BDKaRJ)L-<f-;a?=
Og377>RNLDQPd[A9C_T8HZ:e:\ab:CNBKf>DU.EWYc3IaaY,&:FZW@:c^g#S^).6
XQB5&^L5C1NB5.0,f1A/WX6;CLG5a,6eJ:Q5Pg?[HLZ-e>KRcTJG_d-J]NG<0PNP
d;DX/-73g,(C?FW93&,:8fCdfcAC0+LKN)-X8-^)de+3_fNG?08P<?@X6SC(YYTU
W2\5<)eJ(1f,Y0Dc-aINL7eL9Lf7Jf:N(C>06,8GDF^^ZZ.[Sd.3PJWdN\QDF+@Y
=WDMVV[\FV).(\3Ef9H.\fCII7Q0)DFDc_XF;B23D/=AV@V,O.,7KfOG4CS3PMQ4
5TO_+M2]PB/(a.K9-eN17F6?MeTMQCR1I50>D5B4_IXV;H3]GVI00((B-A&b^8;S
d_@K<A1Z8G@YFd3U@4;Y)GBMa2A/FO,f42<.Y;S=Q;NI?XY2T63AH)EL>Deg(B5[
5N^ON/e-^=KA\aOb>d=X2&[@12YTJa>CFId;M[AN/5]686g\c/DEN,8^=JgLDVW=
_I8]O7EJHUe[F&RcPcMDT75C0;;A6WcFW&2Ve7(?7L4H[5,53P0MKPMFeP6LY=RX
I#FQ].(GKgH,?B[?#PJ.-_IHMIL7N,9(XY@ZK0:e.Ef(LDX:V_d1gN3c3<VTP0LO
&/K/J]TeedJ^#7&#>PQK=A\NSL2Y?FgGa4H.A.R#dcR7G2HB[3DPbJR2H<Q1)C]^
C]d^DM=GQ?W3W18F@@IIeDTVDVbT1BO2Z1DV&RAbcIR;[M9255[^e\a1+IYSQ=#R
4MM_++9KXBK\IXd=2;:IX;2ZOgMP[KO[AV\>NF#.EdZ-e13_g[7D?dWMa:cNCUe^
bc;OE=bA\1@4Q;I-/,&MOYNc4,R7,NJJ/LNYJ7I68=@&c5ZTa]RUT3bYC(NHSWIQ
BMdTAAEYSN#VIAI_D,-;NJ)BQ-M9e_<J4PB9-A8TTSPN)^>;,5;@J=bUb/^#[R]B
]EQ&OY<b2bL\@]Q=ALH-)&f0#XM.E-2c0\4AQ]WQ@7fPBg&4EUb(ZZ;63(,ged+U
GFD2+VT8]3AC9J_I.&dMMGE>DC>Y)#BD]13&5?6/^>@.6+_ZFPTL)HQGQ?J?DQ2a
>N/aA[3)U<3YKSML,;6C-:d+DI.]QaJ&0GJ8GDD&.68cg2J/R)Uc?>YAN9cT=9gT
4SF/TY6PG3:DAM4+4DV+ae?.?&4OTOUBebGIL+bHR,fMb3,_<<Z6RVS1NJ6UfI>Y
\S+]?@@bH??;HCWU(_-\2aV;e4F72Y.,@cSJP.S&U3EQB7PH>IgZZ[J^IO)/PgRE
)_cHa3,N/B?../1I\(d,EE5T2N,;eL6SGfg23?.J:TXf&7US<Z1BeD>4\c4-TF5X
@+GFK>>JC>[6H84<)\OG-aC6HOASU2K5-E2Ld;f6E\)U[-R&+3JAV60YQ8[[STT1
bUQ=e4Da4&DMgLH3Yf2APEFZS(AI:R>+<^-eHeX,1bIRUA[@9CH1ZMB9/b/cH=UE
,,\Z<2#V<1,&aQ)I?P47/WdbY2VPWa#OKMZ59095Zc2R96H98/5B-(d)+)51@9aN
QXDZJN(5VER,+D&;]]4^g,a-e&fCaQST]-dS[:RGbE,d37dQXY\YXP?cUgW?gRFY
>3K?:\c>1C5-c#TPa\.(ZAb3HSb=2-^[G0WX\:Xb=TCOO;L>aZT2E;5(8QJccIBB
2]3fAAK&]AcUfb<FcE-8L2Y??d+?C8]S/.OL:AaJ>;6H1WTaeD6dA5Vd3/VG1a?#
A1O-;+9US>=3#;36819&#8S(0507B(aRVB,d9YBK,7#6_,@[8IX8-&PC<74B\R,1
F>\E9ccQG1#(Xf=;@]+E/BFZ\,AWEX\dbM#de7YB1I8>.4IT:C+62E31b&fN-K7e
^+&(\\e1I\M9PQM[Yc)D+fH?7G#?[_deg;LTFTaAYTAB2S\EW.YNAC0b?>N884J9
F0PV=ABL<DTg[g<VQ&Y[7e4H2-CeGJMPLUCAQ+T7-d@N=M9=e5O:7I#PGN)b>5#8
^0QJXMgCUZK>H[FcXK4;DcY5L<VcL.0,\R#R3&1;GPILH:Z0R3g@R<UGKPY.ZOfe
/\dNg-cEGIOXN.2-:04W0Z[Z.GJ.=(A\W&bZLMef2>]7=6;/#W95+/K^YA.IUJ&E
b<7\PYG/[H12N(4#b4bIT7:EG\,^NV&bRI)YQHDC4KCa=bPJ\L+BfX2,KMN;D#W:
OeWZd&4;HHL05)7Ub]a;UPW@cR5<@WGB)Ec;SC=B;1(Z79Nb;]&d,_g>RQK?\Va+
(;JY#8gd=G5F3:d70NA9\W]U(OZJ.c7G4[.b3ZB/2.@0g6YSd9.05;.b,FKIgOfG
G2GUg0>S&@Y)e,&5HCWA87JedM],US+<;bH4([N<1bMfJ)L.Q/DfAC^WP0]VVD0W
XVH,>8>D05d;/TF\@e+&9RbD?bAF(U1>f=Y;])<cQD2TM^a@cH)+e+J9-#.(W[@E
Db/TH=8a_63>6#&9;),@LGS.8N\U8NO#]5caQ5FJ>/cJ88Q[3@+26@W>UbMf]E=N
L2f8LJVKS@GOT\Ta9;Tb>BR9GFXEGNF8W.[dDIgF7ba)X[c]1WDaIRETd=\3>N/T
g<OE1-.7R;]2/>3(C[0gbD6EgJF<+EX)fcK\K5:+A+:QP#/34-2)YI(CH#[ePBLU
)A6aIT8-[PMeMg?daZO?KdQ(U,ZSd([4eF;aS=\@_J:U7a#7>H+QbbL6CHVIEaQb
@^;#M=_2dBKO,Z>\O)\9>,A?EE/X-5].Q@V/30NA7EKH5HPTT[#1ZP917O/4F6+D
_YYZO1gEGW2.d6+YU?^-)5<[L49=]DHA/R3DKfd)ZK#aXLZY0+Z,g7/9(:_Pd=?4
+g_\S)(2RT:I?PEIOO:Aa=NO-IUQICH\Q);#a+MGAa-TCbYQ=5Rfcg,J<6??82T&
O^R)U=Z#985<4ET.E+/E50F/11Xd]M\DLc5AgVWB35L@K4PXd5de0(X19NT4fRP6
#/XW<T7XJWS-fF7ZgJG&IJDW/df.^]a[3g7+AMG_)#U)VTKQ9FK&INTNWK>gJL-_
@T7NBA\JV>aECGNBP3K3XQ\Re,3FH&aeeZJbK+AV>gB]01e,@GR;+1;Xg?>ANM8T
FbYR3R0UE&.<0QbDF0)bH8;@26Y@9HS\/d_DbQ/H@(-OAG,^WJFJ(6I2QUc8b6FZ
,KV[KA[L]E(FN35#)15/Z6ZLOHK85EEF-&M@D;M3FTR[9QdCMLg9V.08NQQ?AS6K
#b95QaD1S45edUHPSXZC<?FM\c;+cN&FRG@VF^6<Q52S&A?Jb\XO8g+><]NZ?>A(
aHWW>3>E]V\)@]U@GLBQFHYLY3=UJ3[MAF=&BG/d+5OC2;_Z^:@ab8MX.3?04SgJ
1[2(\J?\?Z(=#9;9>F?BSFI]8(<M;4T]ALW9+g[8>9E3B3Aa9?aFD)S>SG^APdPX
N>c(=/Q1BW4g+OBA,0HYN26ef5da6/<MNZ6EaaK-N>)Y710@38HYZVcY6I814dfD
XR1,G2MLJK;e]Z.8_Q[Gb\IDf.]f)ATDG32L#H4b@37/&=Hg9#ReN<D-0cB=bU&Y
>=)#+7gG3MJHYfW+//JVdD:^S2AQM(8ZaOIJ<fMdVK-OQ^aRRP=[#8A&QJSL-8L9
,ZE=X=:]?^M#(d\:@<ID+N.O9Z2_74:@S6\^MU)X5/)H2eZTcQK4d>LWI745M9(b
PWW)=C/cE]O?ANPR.L[>1_.=_.Tg:1E05c5GFE=+N&fY&^<#[\6L[])W6c&C,05H
1@-P?IeE^g83GF;,D#R=TWb1=]ZfTcfI[7e683,UT9dLC0#E2Y.NQYS=)0\G((+Y
030VG&&?[500MV@R6D7F@Q&9^IK1UIfPA.E,RE)aGUFeP8f-,EcZQ):)1c<5D_Z_
A5IYL-eG?e.=?4Lc1eKK.>Z3Y@@4-a6)I>egWWa9d(EPN^dDU07?ZWF@6EY3EM>(
EGBB5DdAAfWH56^V]V2^X<a8=[9III9572?C/Hb_Y/=SBNZJG&MS=TPK+ZD.]:4T
V07B6_JQJF@MW=XeFIZ-5d^(Y\8bc:1f3DR:dQ]:XS9CI)I^6^<NEN_CHFe8_A>W
^_dUU5DbLVJ+>VJJT=T[-;.M>d/:eOM(2<^0RaA(Q26,e52S\H.b4=S;4NCBGP@Z
Ie5cN3a85W?;[.bBWEM]^#P(c7GEZ1O=DN;.E]<\b3fR]@H)g=B_Z;.a0>Y4S>cb
O?W0(XOZb;,UVCELX>Ue@fe=NAHF8b(C\M9[DeGXLIdbB(+ZJW3EeKXP^P,RY#/Z
2)\>?]&WM61c2,YDPb<U.V+NXgM?=UR,<6BJ_B9ONJI;Q4GZ5Y\(e72<:VH>LMIG
]4_SCNae+E#Fg5LM\QVJQ,,2OPEPVbZ(IY)CR]])REWY3<L,.<GHPF611;3+@^b8
RN5ZcNdR-&>a3@MSM+;JeCI\WIa[SDM?UU:<>7LS8b+Jb8X8CM4_^aaLK&J.CW&C
-@e2EKIN\U@[95(+MJURgY-GUKce]DJMZ]+[d&S0^O-4[@7N^&-N-+<UR.0EOJAf
d--JWdU>J92Rb)ZD@M3Y2Y4FII3@bB4:Y0W;T>R4PZ8d/d81b)L_L4R7<Q1;B>Y<
@B6Ge9TgY;eK2^?[(Ud9Q>RRA.542b&QUb0D7?2C-/D91OJM5CM6+(1:e-VP<0SH
:OWP(eJPJ_BLWCTX90(4ZE:-=cK6Hc)<1NL(I&2M_BS(^J@NP?O^0S>T,Lc34988
TG1gGV#Xd/W1@>28DfW@0.FBH9D9e_6AY9eY?bD0YAc<d@UKVNYX[eD^P>N)KLK)
UI208I;HOIS,-.[YX5@(MWfRV6e;T/T^A8PHTH311FKQI^8KQT3?a+DYRQ83(\bL
e=_;GHfA(:(71:T1<R#F_V=9&a+T<<N4Q&>30eZ&1e_E)[bZ)fL+W]7)9,,a8(g>
X^g1K+LZ&cf).,]MG+^fgJa(B/dG20-+c/-KLS:Jf&Z5ER7TLFJ:+]](d+)(EXJM
ZY+HIU>L1aQUd<=J#A^VeM\Aa:BBPN40207&59Q:]E^^IAC>G,@N2PbW6B2X2aLb
Q>&T59=RD7.6]1EY5J;H5WL++BCfgV+O5)3.453H,Pb(2eDW=b3INd9cX)QI4<d8
R,5[KTHT-B>\.Y1CL&C7?.@IC<dP,0W]g/2?Q?WgTFRY25b@31SR+2M;DSdaRT<7
,2aZWZC@;ES.Y/WMU\R6-OSe-:N#CCUa[:2+JB(IJF4ELLZ#6cCXLMUO5BUJ6<W:
eW&UW8IA+dDWeRdSC&,c0;_8RWfSL\J,cTeD^9YY#d?c];FF1U[S8RMcO.,B\_^9
_We]aZ)R@A::L@^R0#N(gQ;6FHOGHb(OE]Y/]4=)/E0FK;^IZeTYgD+(:UJBaLHB
6?1M:,)[-5V5ZC8,YX(4\_<T&Ub3?,^#FTK1dZeT_M(2eB8(U,&BP+Q2ZH)bERIX
@P2SG[aS?.C8K+4[/EUV@<)f]R2CU.X8Kc7TL>3fNDcI5<538=U]>aZ-6\LfP_Ra
]a=;)+Xg#BGN84KO8:6>C\)B[5eVg>=ZIfcA;U3?^ef<\b#fD<5)DdK]a^WMJ^8G
Kbbe9F]+14)BLgNL&P;fCMN#6SD/U.M(O420f^RJ<\BKeCX0YUV+beSC5OZP3B\g
/&V4B7PB?YGCWC\a?Va(#ZLX9@<bEa_BQ=6#K=@EK2[M,O250ZWU_Ug1adST,ZN;
+#Xc9SO?/aCKU1QT\I7IdF;N]a]F8,50G?[FS.7+J6:++bd\6@H,/&-XX&D6NJgX
6^&FQ2?78G8V6Y;,F(Y1DLR_3VIQU+QC<-;DLbH5E[T8#b.a5HP7Z>]5fO7<[UFA
WfXRF\7N]Z_LcBcb+8LW=N:ZW->&&L1R@P0(4(Y1(K).[ZG?HUDGfAHFd)=?Z#1^
.);QZ;^ceCGA#ND4=B,MaS-KHVOMcTYIg:Hfd;gXKS1)+W]dS>(FQE[Qb9K:f8Yb
:cKZ>-B3?GC6)0e<9.JPPU;UM_X3,fBHbR7-(1WJX@=]cW0J7<fMTYD.92YB7.O)
E#/e6H;THYR4gX@C6eX_G]<Q+cUaO4,Ue>f+3<+L]7HZ-?C^C0^QPZ]/AM+D3R]3
T#5B4S^<L-14V&,RfUGEUV_0fLFV)&S@OGg#g36cZG_QW909>T8?(2^GQ)ZJ4P:/
2^ZO5MS;8>4M5RL#YD#D(74FS(,>0@5SQI&F1c899/\eLA6B&7(]=S)+?8[UfCL9
TPO8=Zf)8\P=DZ-P#:O:8J#1:DC7LXgKc4/Fb]:Wac4J#BFEG:fa1X-PdSV]2/@(
+3GH,5IcIX<2g_K=;2BYS99>c3Dc7T6O6,XIMDJQ^_#/WR(L#Tf;XZ>=SV80cEX:
T>KT=f1-#(JJfE=\85FL\SH2CN61?Ge]FEfdSLdK@1b_gd4FC9F6]^,6UbA\ANRR
F4K@]aT22?LS9Z:Y-6,O&)M,7IXLRI_C8\BET3V4I.<<C8MD>W,DZ02@CWd2MM<^
4W0eLf#,6Z6g(#6]UQ/E-C.&(U6O9)5fA<I#?\?X?=E\N\WWOXNK/FQcFJ(>H.>a
ObNgA3PgMNFX4@T<29W&(\\aV-(cB(;#695&,da_TQcgY20R+_F?;</,TPE_g70_
:;c2(Ca1,J#GG]_bK9A,d_66(:K@B1_BWFCeGW1Z.^-Q+gYcKOa=9MM]^<Z?(WPO
7I]0gPMT.gB[CWG]77H4XY/L74MF<>1__?PD_YQ>^[A==,C)B&KZgd/Y3QC>8@)\
GHA7#X6\TCd+C?DX=?4T3Q6LV\]O=#4cBH7?&.eLeXW3S;SGbfXA<b?7CV/&>+&E
<==bI4OWJI(a]QVN-Y)gPbN@9gFX2g+Yd)Y.NW34I#;;.,c:aO+ZAS5-A.&f_f,K
BCXReKE?TXGP:5+LE)V/LKHIZ.&F5c9.H&P>ddY\Ze<IJ9F0T0H?8J)_6bc[KURZ
3?Q(6KRRHZE-QTS4T-6:?+WNI<+0]IE-_C8H67a0M7.b^J8Z?(Q1bULE<;>D]0+4
+LO@aNJ]2VT?HfNd)C./Tg(V6A8Nf]]<AVL]/MB&7T^&\UPfF?T-_8&_??W0M1Z3
QaKX(AKbVgRa/RZT_37C8Y-IX?UB;@K31+O;WbLZNaecBELC(ASW)f_FJAGP(^Xa
cAc0AJ>MX1#][)F3Z<?\WUK^-DF7@,2KSZ=e#aPe-SV_)dR92HEQNZ6KQL/D=A-8
NPV5_-Ff/]J<6bVD)06&GMegQOg&S6dG_G5a7#MQV-.Ye-fbe3cGKb0LU7gAB0eR
[H:,J[/_?E\^0<N-D=11@HG@^5-XXV0WS,]Y&:,14@<4BY^;U;<MF.>8eZ.KBb/1
1<E_ZSYUPb4(3-+O;_O^E0SKSRa+0dJ6f([8f371UUIS,6;S^DRf-@9X3=B\a->\
^A#[N1LL:28IV09:de?+_e:E_2af1c5O-aH.>2I)ND:;Z4/R0R_:H\1,<7c8)XN0
_VfS71-GO3,<Uf6_R_AaHAX7eGY@J8REXL,_W:K+P21>5O;\=?8)KIU\W,KCS(C>
CFJ;.\7]AO]0=BJVS3WU(>WbQTZ>YHgNV,dd,C<#)N3>e\BQ-^03Q&A0?a;GdM\;
bV0Ad+8K^d@VFQacB?+VdY>2&S_Jb++JM(J:2=0?_B-5\8J^+_AJ(CI074&A#VL-
f#X14;gG]UBDgTU+)CC7.UASD8#02G6ZZ_Xb(]\XK2CcaHa<T1J.SdGfdDGeIedT
;^+3ZL]_C-2&8OP(4fH?b<.#(A]CDGD#6>0L3g+FCaMWKC<[/YU1CUJUXL?O3@P8
]_M>673PRU-HbY)0dg]V(C[\\0-,7+]aE(9FQ(<@\\#\g+\E8BQ8[^_O)d5PR.8Q
Z23F[>,9,X=E5>>[C5&LfXDdIaCBKYSY+Td+ZJaLc>U&DJ\FIWJ764e?B47,3PP/
6?ea1IUA@e?G.^BEM<\MM)WJQF/P)NRg70I><7V5Z2S.(J\0T=81ca&Jd/4KMdbe
EcIFF_5a]=aON1VB&L@@.^1@731T8DX+@J.6SU_1_]F2/YfX5Y(PUZ0Z_R31&+_;
4b0=G,Q2<9F4c7I.1RK;6>+Z6_5@_IfWO&P&2T.-.fd<d-V[N=VC\(J@GG0?-3L.
ZJC/E3G0K5QSdTK<Z.abF()Q85T:VS#g;KTcQR=N#))WZWLE9NdOB);H6VHK(ANQ
T0]aVHD,/fS)Z+.DV[O@G1T7XU>U3YcKTZ-S:BNZ=^[P_[X1SIgBHCcL/D+OC6:&
B,3CbUT1>5FEOTWP,XBDH&[3[YgD(cNcb8#7-c8#.TW89A)H1+<bLP:(XZ&GNGFP
?3a5:I\f@_Y[687IA/SN#?D:VLY(bN85UHW[#bYTK]4WQKM;H;JAU22c?#Od(E1H
DD]9;.M=CdQ1eSWbN)7[\OaegST]QGU6eWNQ/Q-51<,.KT>-H3dd1T#4b271N(Dd
d=e2PB/ccWLCHQ-1?B,32VK-P-:[X_\6#[I;AMJK+W/J.;:^OE[T7Z<I_fB)Pb.]
b#JbfFATaWIYgB6,#S,.8b@6LV0DS?A/KOOa[eB[+.?2fb0,:V,+[C@_W_WW.B+:
#Gf[F2:<E7][Gg(/(@,=D0MNa((YMDg5E?91)4]K&CJK^:[b6,bT19>D2F&/9<N:
7T7C4T>OT3TOM#=J6c\<EHIc\.&.+X?B[ZWX(.-K)GS.J2HQ>P(#->T:=EL)G-S6
R,f6#[+,aJ:BGefARaX==A6<_YR1JMBD2XI?<FY+(4:P:=XQW]Q+c:5N-JDD^b2;
f/P3BYfV+#OO[H6dM3^XAfNBL1NW:_IJ8791[A6UX;N]0-=O/6-_aL:1_W>90&8?
3/A;f@=B\#K1Lc#\VH@KA3,eR.;91X;-7.(^</.Q/1;]dTRMYO7(]f9H1_U489.\
WI.GI=89fe-P53]IXR4(K&g?cbNR_H2W)(R&DIPY=(==#LX)A8VLW2b)>O/]gfS8
(+VAHSC><]QBFRgFP)+[JAQ91BA=;#\0VaBBGdUGQJ8UF#[OYN-TAYR/T?[5]d>E
I1C/0+S7].I(22?b#P1G=J+J0g:KMf<5gG4PB:I)-9.1Z&BM+?J&1LFaOF>4R?@X
TGQ\[UC;,Ed6))8c(4@\?Vg&gAfB,2Z@B=#VGR(4GAbg3-1A\f4=dD==<.P6]Z[T
[U>MFS1^3J_Q[bg\0V<W)ERcg3H#L;Dg:g?R6^?3L0F-81=&>G21)I7:S+@:_;LA
I/6ae-HQOA^YVd(:+Z<@e)Nf(/(;VE5[E5g]:<H0K2e4e;L\GEWDg=V]J,9_FH87
\2XA9TL^,S/[;8\1KXK-MM^WKM3gf-MSXf0Q:XQ@\K1XO)TY)MMI?c]=#\82B6Q\
V2VKPN0D2f[B1e>8&<ADE_B0,S_dB\@b(J,>M[UZ/c4F20MQ#18#ce]1J[N(dX9E
c^TTPDXN1>0;70&]\^SR^9W3cX\O]X85O7:(]5]AS2e)#VB6=(_7e@5N.cX+?cMY
E]47+M@UgRTVY9fZ?Fb_WdS;XdU5dLd-9dO->e\Yfb=-VX&AF@N:=#7@TFN?9g^0
]EIET@8NMT[5)&UNNY9#@XO2YeP85(O1M?e5OV\&PP6I/_5(BUeZ)E@<VFD3&>Wd
eV>aWec8Dd:Mf^,&2;JO55I4N>PDM<?1C&;a8c]#\T0b3VbW(bBIBJ]1<9CILN)I
7g,EfMO6b&#2W=G0[eC)02TU2MBW;Y(7#f@U?UfL1^SfdCUU<.PXV8?[c/B3UT,,
48M9Wc+d.)R72MAVe>54QH17&EF^eU2HQPQ#C5)O0>5]aK)5b>4_V\Q87R_c2bgM
G9Z81.VGK2-3L>ZP6VABYQY7<SC,V78ZM:WcD?a#-Bb7R:,?cc@1<@(8=cJA+:O&
9bTX_GA=/e[L4)3T51L8=9GL<@I\feLd6H13Y1b5=W&#V<9?);-fXU?HZPZ4IDJ1
b0LY.G?DBZ15J7IM,8bI&,Z/36b_3UNVWM^(J3ID=F/_>[DV&K>V@N>,6MXe9^:T
2Fd\dBSBB:Q9W57]L:Q#P<<WI0L:5>6K.P/+^I06]WYJB9#7/dI2),7RS#16UbI/
bZ_;8;?[4-YK)H=Y7?Ae:e.^bgNTY,;VH5&&V@?2&V^UBV#/XILA=e]H;98S#AT3
YG\,RCNEEXP#gZNe4H7Z4bK0YS5.]85K_Kb1Q9A\US^SH+HK2DF0L/VVJ;H^J4X=
ccQPeE?_;bVQ6-D:McR8C#fe#&LAg\2Ud9[+?6+16@c/,fQgN>#QAT?a_)e;;+Z,
Eg&HO?9Kc(JQXd6ZY<gUUPgIGf,2LP3)913Gb\.?;\_BSg/IAI-f-g.F&6bA5#^-
]\EJ>RF-bKgR31]C(=;=HTW+KI70/e5E\T.)FF8I7.C[EOB=CO\CS)agE\UPW42I
.KN@8W/]1&659BYTPe&G-a8][aS4UV>=XZC(DH&U:U<[T@50e)6QU#J1R)(;ZWKF
Q/KVdL]BSSNGcf6[7;QC7N:5<B>J<MCaA,17>eE-ESbHMPVXFNU5[gF&d^>?V+59
9XT9gc&/,5)SYL1O]R@_)QN2X89;KCO)g))2EEb:,57^<DJN1fM<W6X6N3])4A>1
X[#VE8:X;JX+RR5GZ4G..S4aMBaM20[a[5YEAU7V/@BaWZA:F11<>_96R#S4<f0\
,_NJ\1;^=8Q@IQRc?_T3<?5L&KX.,AeCV@#caG4J=S.,^.;&?9\#6X]11Y6<MF4<
-7.C4]9ebIe?dFW/[7L);//?agd=<O^d1,SS+\]XPdMd6ITZ0^eUBRQ2L]FbgFKY
TfUI>Z#85:X_eV59b-Sg[bJ(I3ZdPDYK6,UUPD1:<;8Z>SS);5LNdPSA=-PR9]cG
H7U([^+3R.L<DQ_G7Ec<:8@MI)[1Vc@UDc6g:6Z??Va)>YSS8+1-&gH\5N=RMc1E
-A;41:BRGB=]6?[4f;/#U\Z2TcUgc#9HRe(3Y>S8U3O\,EO^=F==EKeGLUJRAPWX
D^@S,KaQ18(L31Lc5JHWUB/=8X;bL05ME)C,Z<&6OYN0]e(SJ6Qc0AN/KDUAG_@R
]+T^cab-(PQbf<Q\&P=(J=\C;66Za[f==;3D8>TF\]8>D1<=(.D5SfGA@aa(,@e=
A1-3H^1cebW^V@253A]P:#VLC3C4FS#A5:&fYC[41D57)/:8bPZD03f3@\BC&:>S
L@DQf98CW?5PR.9)Kg[R[9a]2.2Y6RfT[L4_E)L75-(1(,HaQLJd@T>LAWa?;90a
C,&CEF&9.NI<)ZNeNHDcLa>P,AFeM8AHST7-7;VI0V5A7YZ;5(Y=V)Z,HQY,W:Jb
WYMa.P(e=J@>P?^8(DK#DUP:5Q,ga;IUPaI,T;2.3c?db7H+-^P<]9,AcG(@PfI^
^/<3NKbJVR-NLX&5Y,6^-WBU+^CfI\.X0Q:7Pa2U+LR9#9ZAJbO^(K0I^0SYE)6C
CO4?AAEWRcd(+]O+JZa_a+I7<,Ye<WG]M(Z+ABf/T.78,1)R_W+26R:K+e/=>@AO
SN?e)d/XP2)6B28EW7:_a_#BacXLV+ZU0VgAJXZO[?BNd)HKTJKB:-AN4FeBSX^9
)GV9)HF^2#UE;T,gC?Z3&PU0Y(>E6265M&SB1J91O#)<CggLOWM[;97g40NN\d-\
=-MF,6:D+2.?:aJIX,f;H3TB[:)ee7T(G37V?=\d08gK=RW]\EB,E2[?5Y@LbN^8
-D&F:g9<B?dT_Y1SE9S9BZG^E]OAcUV1We<,=F@@+O]H4YD-c;=c83g?G,2]@XaV
1CZ-VT.ZSbFaOY)L.E(?#8XJ4(FPOeTgOS/4WQ=5UV)JI=L/(#/LCR\57_-]SbGC
7e@TV3W/gG1KCc0&S?f6KJ?J;L-=N7S)8VgKRfUEgC0IfeCbOVPdR:WO-.;[XbMV
37?3(M(\6,H0IGa5\Q(c6,#__-GP\@UTg_.b=U?g5C2(RN<@DcD^=L9Z6/B]R22F
Bb4W5af]8E4[W6>4+KWAY1)d2gQA0;N4Rgf@5WTCcWCCED#c_LG<?)QKYGAfF@<^
R=I6cX5^VX_H^<gL1Y.]=)/84Ba2S>\cHS.DN]&\:-UII_;.XKFfc\=E>BB_eH)W
gZ\[g?6,S[-62a&LN,=TQ<Tb=J(eLW2a4Q#XV1[A=O_NNLY3G<>W97V7943SPB#3
d@&K,E(Z4Wb<,9MOW&Z97IRZK&WKVKM@PH=LY>^#L.c;fCK]D12]W5d/8T<2>1_)
7I.<:&d<>1FREcM;V5F9.I^RDda=6X63^YZ)c]M[-TY(E)>LLR32E:d2<V()c^.T
H12TI/5/bRNIA,8b;VX_CHbYPcMDA[&aPfX)ZW-5_(C#Ub70B0=^?Z_a\(3#]))O
[G2LUD1OPc=J@<9b#S^51_=V\Aag&6Jgb8EgJTdZCa_40CKC7YQ\9=f_C@[^D0XF
D[;L0D.+V#HEMa6S+g[_4YJ.d#^LLP;A[:MJ]GQd_DX69OZ0O#f.;PF8;G.DGIY;
T,D5&S7FA<4]+4>,3=OPT=fDMdIXgcM-@1e-X+HTMcH[A:O7Eb\U?OU0/W+TPH83
Q4X6.fL>^/B#[S[#]CT?0f_P3N1/Z_F<E0OC5QadeQIN?dK&;X<]LgP+AW6;KOYP
1&bIR<28c;Ac+E.6._eg?N>3I&J^U/)O8NX#d_+1#fP\@_7LRWY]2@QT\(dI/.L)
a2>XH42MA-IY5@\1FCgEaU-U,7=F^P00G:H;0GUJfNOS<:)[:HbO@.>6H+P0:d_A
e+afSR]2QaV1GFD=:_5I@U)X#f39S\&f5CeI(67CB[3JR)d_>dYXGfd_TC=\.LG@
-J,A\cY81@a?4?):L)DgOgF9)+/2F=76R4bHJ/I4WY+6K,<P;=ND[Z4:f207S2AG
DS=HH=3^cT]>FB+EB(eCgCG4DEf^C>7NA);_K\9T=0KfPKU=#P9_)YO]):+Qc615
^efT;O9ggFV73^EEbTHO4gHCK#;A__TY,)]Vg>FD[Q=4MTM;/DY<AQ]R?PaWa65^
IT=EcIX-(=H:XE[b0OY5W->3+,VDd[dd3]#;gA&B3eK3C?V4HE1_0PbV)fg&I\\N
NDPEcB,d#6>RR/ZZQF9L#R#edO=I9I&8DPaX#P6eU@161G<>#=7,&G.@0>HeNV[c
)G<0140MCGQDX_TQbC;e(F@9dVO&T\>Q,UJITNO6aUg;Y_E>VE8)/ZP0,9RCa&5P
7=3&DL0^BDOc;RCGV7JRL,8^;FR4T;E]@P8FQ^BXCWFSJTR<gT6>O5NIZ]g70#?F
(HVZ-X9K(C&(XNQ=BPZdO5e[1W-OHHBY?I0]/AV0.P=c);\=S5cE<M\PW4Z6[Eb1
g>Lg@4Ca+G#4AM[T32e5ZQ39XEe=-B1CO)[4/d6_/+0\D>Z(X2Y.@]K94MGggEVb
#M1GE2I\2USS5W[2JW)]aYS)?8^D^Sb2?aRd@Xc](_L4ba;)?L:Y1BC\U23\fWLS
Z>E[YU+57T.a0_8&-b(^BFO/H0NZ,66dfJP2ff_5=XRUQ(A>D11GZE8=R^HVM=:N
;DIJQ;(](>8754O)LORHOY>7D8<R,dEP5gIe^FLKO:[_G<b&70fd7_VU1P66/cR^
729/8U09FG;MF^.KDb7Wg&cX#XAFCG)UUUe]WSIX)HH+)@UW7PLK,4IO6MDMDB\C
LAKR82=9@TC:7<)c4]Mb5S4T(?II4<X2?.3fFQHfg[BUEFd88]<15PS4\+[^\GL7
c/:)HK_TI#bG3ec0[Vf,>b.<8E2CaG_CFX:Y^CN2L8#1)Y\e.HJVHW.\_&@A;[]H
Wf:_a@XO2aVEJed.@USRFOT&,g]FQJ0DR05Ce0N_-HX1@2\^2RMM(D:9G2@g?fH+
JVGY@D?I6<[V^@SF.-dX/;_7-[b#\7IQI.FNcg\RU]VWOCd0.A7U]R\5ZS+T:P^D
J:LGZ&Z=+N(LJLO73U#+A-g[d/O?6+;.MM5DZ)2WX=/6AE-gfC0]a8DYH[c6eWaY
7;@P8cJCN<//Z;;\PZO&0[#=gS)9CH,-K_cBKaYSB459NYDT^YSRA?DYM$
`endprotected
          
`protected
[b,A;?OSDgeKYH_=I<Y43G[)cRIMOb\agPDA:0>L?4>YMLVdQ.1&/)I^dF\O)S;B
gX@g]CP84ELK,$
`endprotected

//vcs_lic_vip_protect
  `protected
UfXaNg3.C#037KNHC/ZQ1<+e=QSd7P\E5F;9_,eK,Fe&,O0Q?4[g&(LDM[R6UEe8
25.)ZgV_0/S]LQ7O<bUR;4I&7WeTe)4ZD8=U5@L3=H<Ug0-]50DQQdD+GA5#.W-_
ELca,.@_T&f@\eQQ\Z<3KWWYJg.G11\d.,3NaBCg0gQE=2ZVHXL3?TI:9;G8E+c;
N-(+<Fef@ZRWe^f863c_@F.D-EfX-1NH?UB4c;8MbFN,I=BR&\gM/b?]DDI?N2:X
5;=EM\BEJ6Z.c)/,-g\^([9SF5NAFe<PMXP5<,4La-/:MG.^UNP#B&[,BV8Z\7?1
+Q+9Z4[O&9;PUfJB(W^5\1F]3=8Q3V13Hb91e9HXP5RgD[BDM01_Gc]dDC,FT:_;
:<;I\dWO(T+Z5Z,DfA00]6H11SeHe\c##]AT,Z3Z-;PQ@aI<0\Z+<f+Q@8Wb;=#1
9#)PeB2]T1P3K;fRN:E:T??I5MZ/.Q>XA;;\.e-Fbf,TWLfB8c,]7IE6RS-+B\M?
\FIWN;V6,SE75FZ3T:VYa)2E;GV(#2+--<;]e<=fbX\[5@T9;L:=J63/cNd0F@D2
.85,OV,UfIYda&=#DXT,g;YEe[8;N2S?&?(bMM1V/&BQ:XJ8>W^A8PET89cX6-+\
g^&DPK&CXR1[/4)^3JTb45WWIGBV<51Z<2:KDBP.O&Bb6E/Z?^8M@W-W4Q;DaPO^
HRagWdV<\b@]B7V8=0]L<eQ-J:J\[VY#fN7;1eOKVg5G<CcfNA<gPSJc^aKZ[.V)
gN:J:96,)V-_3+GL6(YM&R6FXY^SD8(_;:_1d=+ZU-]=a35cP_b1T-#g<1-(FJ=0
&IC<8cfH0(9Bb,g-Ce65>GgRZ.1QJ,1&EQO2MNK6XR<aG[cX-N9Fe+C+BZNLC)I7
23HcGFE3/XeCJC5gG#RV=WP4+)M<N+FHN+P,M_4d08&]/g;:LMY0_gTZ]:[D\+L?
/RY7DYgX9aCT^Id[_/+bC38B>24SS]36[FSRYPK^P.-=T14#VID3^0#LAT[3[ZT2
T[G?4G6DW<_MMRcO7UYBCU.-R0H.U4ZP&U]1f5_(U2gCI:9ZU/&]K2E2cZQX-eEE
&2HU=T@P_AN5\&V3S??Eg30I;B)W/>.I^J<OSQ&(NN-;U>X/?\LBN0a[<Af_ZVHF
JJOP-XEY0R4_C]#3YA2+.-\FWQR_SZX/1>Cc#DJ+HROaPI77@IEfL4?>Ff/./;+(
A)Z17^I2)R>BBLE:a5[_;&2@b-DKAN/#fa+XdWg?Mb#\4ZFO@GEY@EO,3\/ADPW2
f;dT_9Vgd\1D;GZHO29L^M,<OFX[F)H5-;SV<1CTP;f0fX97Y#^f88Q/b:aPM&Q)
TV6>BKRDP1Jf3&R-3,)c+&>e::B43&Z<.:81&Jf;;cO5)/#,);M=O:IWRW0dL&XM
+gFCDK51CM=;Eg7Q<M2K76KY7;0^6bB+:]K-ZL7;Z;?MOc#MHFgU9OP0NKJ98U/b
,gUS\\NQ5XT<<J:+-IO[(WC\gP)IRd>bFHD(WVRaXAX8QNXTKE58T-D;^:UOAC3&
b(,dG(UBBcc#^52g#,Rg_W8a(7Lc3Z>WGYVA#fKV(PX0+@?.\Ba6R?/2BHZ9+-2Y
BWTACdb-OCc7\ZO@,Vg/B/QV7[-0_>R0>HWZE:cR)&1<,aTNQ7IUR>9cS((VfEIa
@3V(&Q[]QH)Y-aWfCA,<N[PI>2JCb+0,J&3JRgE9eY=AA6OgZ^](H2HE>a21P;6/
-<4>NYU>#;fGFE?GFEE(&c,DGU&L3@CZ-b-Q2JY&e<RO-0&VNc:PcUM,^HMOd](&
4OH+g)MbL^fP>SZ?M@1bD&BRZT39N_>F/_R/g6M3^9PKQ(g],;L/Ud49O-]S,&/9
B0YFGIaBOWgUF/M(Xc0fQ<3&W@22=+gHW5C97aXO(JFN:dA(P<,[)cICE-5/D(NY
9E1N-fbQ^MHQ.MIO\b2;G+RNO65DJBO+SK^f_(eQ8Mb9&J?JSV#(I,#P64[[MX])
1U,X#/6L1,FI;>Lbf\g[X7P1]0-/A]D_[8]+Wf9GJ37]Q,+^ST#TD@.baPHNY+5N
IC2?g9TO#,TR+@EP0f>/(8e5A+.P,_OKW7a@Wac&&V1NA?D7K/>DYU]JGe-WW\Fd
Y]3.+-cK)&]CXE)GRe^N^MZ@Q\:6922N:?\\E9WEW:4X#92Sg>9,BZ?LK3IBI6[I
bd,If?(_7304S8PCYSDO[Q934TF\S4MJ#L0bKLgG9>;PLg:8AHN@VK+466WEB1&E
;TM63\OFZcaBcdP@JXT^&IPf,8(VO08R(fQ&2MS]P2e?d=(-M3Ue)_+7G>G:CHER
V_M(Y?YD)R:PJ9OLKX9UHHf\6RKM2(/L#cRDdQ#/<D;?W#YJ^B=S967841f1S2F,
#:Te;8[Vb&DIZ:H6=AO(^@4;85EaR_MAJ5,;VDS9F6Ia><IDG.g13[=8:\K]N@[I
B-7JDJ,)&,Dbf-cF8D.;cC2g4C>1d@#1_;5e+XT7>AP^[B@Me0DI?D4@HAZHNWe&
-@R/a#N0VO0E=3W7F^gV6#;/CM7+(b3[.;KDXCPWK7RE0C1FJT-^(R3b->RF_QG/
S:-FWPY^((bOC#3K[)Z@7EdAZ,f51[W&Df?4KYFERD3aM6Y^97D.RVNgNXYS7(BH
<QI+?D]F9IA&,:A^BBM^1=RT.^(;,;3f5I[5YgBH_6_2K)e+T:WaI([4Y3641)NQ
6-4&?N?LFWU0VKO7<O^]\CUcHD<AaWV1F-?G2T8YHd=T#]@@B]cTB>30KS=?(N<4
8-4g[;OQ_UV3RQ7DWPS+KJd\^XL])+J&Q7VI??R(\C&B-aO[74(H88BgRU/\aPV;
)@^ZfRa><a_cB#@,/K1;Z;R60?>f9b.V=5K_291cf_F8\0>ed3,GII2V,F^a\6OU
5\3I;<\F-SX^c51>CE>KA+033a8[GOZEScg/4),PeQHg^C@N-T0QB&?Wc86=#8f)
<^.J?;[OTXa0)-7ZcUBM)R03TNePWVI6f_5]bC^5,&_XaNQ<eO8c9UZSH@+<X(T7
I^)Z/<)P_BbMXTc0GR6(\TMSRe#Vb>U_-b@DL(U^67@e)([7W8S&DGU3]N^Y8QX[
V.99OaEd;-1bLR-5T#YEJXL7FSdGd;Y.PdVTNQ3L-f=C)3gT2V^^(^)1b-I9]9<?
_N^FGdV,[]O7]N?WM980>L[7#O]RKTCADgZeY3&T5T6]d.]#K7WH\;V^:Eb)5FX[
078ffW/S[BXaA81?+07<2#4X;&[Ig0U],53GK5;^>7b65;DQ:A<4/O8Z,7cLD_W,
HR?<<,1)e#UB&<E4T4TcZd0;3>1UeI39[K0A_@=&99aUXfS+Lc4HS\H81:HFC4XS
@B<4UU<ZRZ\;.fIF5\MZ@>)J5[_&SeJJJH:3;+CfV;/_XIee^=A6VbefH.F<JL@R
6S.Lf3#+e0a\B,]:X69A8F\LVX^#gTN,?C]S_M=7^aJ<e^#\37+&b7;/^f^7ZFeE
SSEYK,TO,QLLMb)RLe#af[Q1F+\.(/4DaMP0[_Vf#SZNc7cLWZZ)/\EW8U?da+_-
<b].E#1FeARE_).JPc0A0LE-Y=#E;d;/10>_LdaU#(#KYFO7YVUKG.<,KeLF=5.O
C,Y52O99#.E6:9CGVK.YVS4J,:Df/gPA77SURaOM[dT=_EDWI#8B?agV464(G4&X
7>?H(V_\UL=I&e8fH#\A_E_N5I-+&e=M6^,LZ2?fMT:SM>g(Z(5;UOZb6B#eGfT5
#UZ&>FJHL/-&]/\[>IPE-\c4b+B<<W,;1/027EU8#[K5T#6Kge\<XV,2VG5ZY(<@
F>8R#[.XB[<U-e0+>][Q=c0@VJ>299LbM2.G;@MR:QYB:5HG3?=6\0U7dK4E-P+D
IK><S0Hg\b](Be9b-eL.\dV9Vd?U7HCS,JNZYe@C0ZLW13EG7RI7I_Gb;,d:VKO-
P&A/[0HI:fZL.8;CbB0_Z[RbMVRQd)E<&HTK1:^Rb^d8CO(R_<IJ^e]f<<VH1A\T
Y3B1S7)2T0O+VL_f,G(>=7/GQ;FMMQQOVX/0W(:M)3cVL32>8[>OFZKB?Cb:P1\#
&_0QDSD+g3K+68O<e?VF.^K8D6M;OI6Y1>/RQ^M-TA&30]>20ce=-bb@A\5((70Q
8D-e)6Q_X0#R-_9:A2-+GC053We(UaU;dEXH?d2>KRa(53PM/LC/+RC_fRaZAX7,
K80dU@;3]=bQ0bKX_PAQ@,BW&5[T(UPAN/VC)DA,\Jd[@).(19@WJ4:\1bWX#eZ3
5-Sc>WA>dW?e)2A^:N\Jff,bRHIGF=I0<0-bJY#&]F=U_V5+:@Y&/</&aRRL^3a/
J1]JgFdWH,#b]_DRQE+<?J2J8b0XX+T8cA?SLJgE@-ef3K&WG/?MX3E:dOI^TVeN
G=6Mg#9_0[-7U-SQDI23FM9WSO1aKTLBPZEM79=@,a4]b#M1:QO6BIBVXD3TQ+dU
NKaJ&@Y3G>c4JMc++]eaCN)JdQT[8OY0O7B>:A9FBdXX2O6c<KU@GM>7PROd7AW\
Q4X2a9_\L/fNbW\RH3\,_-GXbM<:^J\UeJ-H43XeF2:^c/\(0VT4G-]KY4f/1Q>+
b4A/E#RQU[RR<4S(<NYId,]4)EJU+752(U,O/T2Q148H4/)&<XTQ9c>>OWe2G<J-
0.SdO8C^=:):@Q2[?F<Wd5R3D>cK+Pa;5;ZE#EfGXJ:T:d?CM#M3H<bcUA>1M+JI
TAca<819GZRQGG/H<H3b:IaK(;L\1BYK5Z&R#K5KeMHeA\K5E5cQ.+>9-W1K7XW_
KR2SV6A(05f&>fL.5dVY;?X.7b&V):g^FM=fH;\@^eMYZ?6(V=d@8Q4M:UI@8P-R
J;&MAR?.Wf.?g<GNVJ<TY7bQ@g_T(S#4Y>V&)JV_UD/^8NI?SWF4X8X]?c[E900T
KRX[]5(=Y81U46P29J9##F=ZIW3/bRPe2;WLT/a)>?Z3AE^43/V84)#d;@cU5\JI
1]I4EF6deBGL[H22O-FNH;7Ob16F_XfUEeZ4K0ZEfRd/I?&]4CQD6Q8;+;5L7.dK
JV+>Og1EbF,<\/WHV,ab&X1+bM,?TMFJ/[&GPHPM7c3X7^NX-KgBY#<?;EYdKF#)
:3F2+JJ.TG(/5N0=Z[TW(FaV).&>Q3Y:XU/?FBC6;S22\fMce<W#^=(5Ng&,Y#.W
W:OT)Q8FIRU9_R:TX.3BB8LJE;...aO.(F-9?N0eLUEQfP;TXbSXFeD02)g2U+US
.gZ?K5YT/U?^+5I[/>=Cd,\(QE0bF0K7,>+@1;P&ON^CC>aIfcWZ#b>N<8T5GN/J
#7g(:5#cKRVBb2\(KT918PN5=VG@)cd_C#W7[)<0D-Z+J]WL>aV?aO.)W8GK2JO?
59:(T+5\aF\:/2T??<@GTZA)Y5\W=NL_DIP-6-0SW;-DM32b1CXP_)CY[YB5(Ib:
cCXf-He[-263>9WA7-VQDg]U69bR-[)fPQ3OWFRXe87J&,Y(_=4)?VaZd7SNd(<V
]25#eS89H6;\#Q/N4??b+EbFbT_C;=ICK<c[FFI#V;L=65ZTeES@U12^Wa+a0F70
K[FFGMK54E/AT@C.W#N(K,@6c)Q-RH:U_ca)3A\:URB1f9A0@E(cc;OgQc-C.81X
(B71Y[E8Q2C;L_f=GVCePaU3BcJ=c)+AF1IE?F(]#O;8c@g8Tf,IHGB:KRBJ\HTR
]S2+/[DP_H29Q2,&/^D,3)]g97:4<XHHPa97gZfc>6PZ)8R&=FJGbYa91PE^PN7:
=9Fc09O/0g[V:#eCIaTKI]^:_a3^>=R>AQKed/T-C6CID_YZ>V@bEeX2_fGSCC=?
XR\W3+6@V9GZ]I@>B<KG;S4VZU>?+V<b]^0.X.HQ2:FJ5[3(RN_U[_+B(]J\IHJd
V2,-ZZa]_H0),:>V5Z6+^:YLb-W<d+-D5eaFVM/[?0BI:-c:TaC@T1.YES_Q284Q
WWgGJa)_9P(#+5JT:=7<5FC.ec[[b]E;0Y<ZHP3SA7Dfc1I&8OPFceZb1VW(Y8HU
4^5;KE/^E3;g;fg=/BX?;UP(Q3R4;Z+;IQ)_F&>_e:^(MXJY#0[U11NOg<B#Z/^P
bLJNDc,+)d\f>BI+:ZETQ3aL8d+_7dTKJZX3B)9cU=]Cg/B1WfbP4NW4QNg.gA9X
N(\bd?VRG0Y0GB64L=HM7^S_E,L&9_^KY1Y;=YFA^8YdI&W7aHQ#N;e9Q&6KC+d/
SIZ];e1DCU>2N6DbODG@aBb+7dF[?#2T6W<[2;L#+1&g<C#eaD\Y]#2MOXaNY5G;
6B/-?-9fA=_C5X?H7A:>1<4:UVJ\^YTaU-gYd2&1:7GUY2TR/FZX;H4CdS.G1a&&
_FgO)D]<#fFD@(\a,N#SN7L1dJ30[-<F@)Z^>P25(J<WSI;&\Y#/;-W_1OU:_6cT
2R,aff+EYE2HTRCDYc:LO#DPGcSDQ_)G7Z^V2B3ZM@BUb=KDC:L+N9.I9DGCE1WP
Y]g,AVIY+(W1[?(deDWdTZeQXaJf25:a&W.HUZ7_?9CgOC[Z=ER&GRLV-)cf]cM=
Y?SWce=AF-BZ]GI;00.]XODR6SGH:?#)f1MA\_5K3A7M=69>,88^B06Y3Ha1-332
X1..@@F7a4V0-/(F.XL89_8KT</]]M>S+V2&:NUe_@8>OZ>H=5fW9.VNaI?8)BFG
E/cCA?E6bSZDF+E@\#<0Odc#L[5bcUHb&L.+:V1S\@HZHHUO^O9A8gT[>7=9@C0G
5931W(KPdB)&2P#_>#AbI#Zg&T])]d5[Y^[;gND=K8.YJ-=[]T=LIB71>[@J4?cX
cW.&+K,>>R\-H=NX+]e)a&#]LVW9FT//IHQ0<K=A_TUXXf@?7[)UH7Sa(6T?T[Y;
=GcWaWa+0<S<g7G:f?:5cZ.C<J+DS?T(-;0fS@C\gYaY<I#K>IaUKf&8>^Qg]+,T
&)Td6@#P?-PP6B&]e[acQ1a>-L8acDED<JbHd8)D5S@a.FdbLgf=^a@eMX.GOR0[
IV@D[<0E/9TL1Ac48@5O69PEaG\.cU;Z>=V]#)2:B;S#B=YVfbO/6ANId#fRCX5I
\-U,T234-QACae?dGa9_6_;S&U30aG/R(A]SX@.(Zd]X.0EBB2O0QM<._UF8>g,0
[<)I]gSTK:WDc?5D()5NUG7>:;:KgSEY:#U>ZDO\/VNbWY+/C>EY3\4:__5EQ=)<
3BRALW[bAfZd5d+X#R:=GW8,Lc]IYM]MPD>Pfb/HE:(<;Q_;Zg1@SG2T3D_FO=d[
RY.._/O?6d+94LA0Y3+Y/bMeXd\78-;K<)W48<VB)9L^K5f4<ZSJB+8K?6c9?BG^
B7_XH&d95b2(b?KU=7#0HeFU=I#QE@T=NgA2/PW-LA\S1&.bVGY[1f#d[-KJ,f;G
[2:&G(.XQAZ#ZaS6@TQF&\94(Z9@HY[&U0O\7PNcb#Hd+bdaI.Pe\b030(.^R7L;
gQYE?\A:Y3Ee?d3UT.)QDf<QdH&(KA/->X;8Bg9:+1TJK0+AgG/)b8FV<.>S-\3T
dL(?W^2I,ZQfM^VI4A5E&CUE,(]MfU:g<TRZ2e6M+-O>@fd8U0CZ)RK/3L2ROIgg
?(+OGVV<eHF?^cN-?<-(:XU?@Rc7B^>cC38XS.]&SJ+4=DIX4+/=SU4IY>O=A4UA
C<_UG+<NgRJ\[9cGa]M<Q5cJX_R1D_FXdV<f?H8cVG&<?L,&bEfY)A?^O>?8?X.L
TA3\cL[XC14(-;&RW])Nb#I+&J([LG>3e]<fBDV1McZYeJVXOUJ5BSY1F2UHFTD3
^W&S(?Lf[+IN;<aQg9RA5WKJ^;7M;6E&^>S9cOGG1<]X()=^VL9:e<<1G[Ld@,E;
f:<RUS:fJcTQI8DX]+07SOMaL)Ae0g1,f#b3WV[A@\]T8g5]VMSR>:RR:A-74N\8
M]GY=EcaEEEBQ:&4VQeNDG7eA(A_ZRW4D)&)/)0;-FYUI8/RT/:6gbZaMB]S^+Pd
+NB<O?YNbTK8FL@B.@[[=KZ9,HF^CL\HNPX[G9bASJ]4a)b72e8NOc=KDUBcKD2<
:Q>Q^f/8FA0cDFWUTJHTB+.S60=(8W>SO0NZ65:37Ja5aG9/0,28-#O=P23M-SV5
#+GZ[],0#/G\Ae/+ZU.22JL/V=XTIIUO/a2BC0M7K\W?=:YK:Q3bca0=4[I&LM@+
7D@_-0@YW/B+^8G54cLUBAfD?RA0cOFL@0W/]f3SJHO6Y]cgE4SYWa?7FL@B[7#e
3.SECdTfeQXG6:R/Q&A:>TJ4TFEIG-\bBQ<C\50ZSTOJ#]?MRJ6;ce.P\GFCV,PR
CFR\\N5-#_]6RKI<-MG@.^=c.7EOcV[_A][&=T=gg/_M7VFY/D.aA?H.MgR?EU:(
2O.fI#3YPaaXB_N9J6gE]91>J#;_T.g-I_JMFc(I1R7MVa8=SOW>-0FNNV)H<#D<
gJZ#ZWE(ZB.7=).^(G<@]bgHcRE:T7?@N7N\b5@B955CJ49BAI/H</YcVAX>aBUe
)P-HRdAGQgB26CJ/\Lf(I)[;g[^1VTGX3?N9J:_NAa<^3dcGE2FY_[V41Sc]U6[S
.+/T1UIaePOS8d@7E.IcNJ^8BF#NA5U#\(QP.KP[)#F5QW/cHJM5<KKU,D_#Wf>9
2;1^d&)>0gVL+;]7XJG#8C@:6L(1T6FK)5A>6a#P(Z.@8IY.J3RXIb8L&_EKY_TH
XFddD.BP]>#&]G6)-@-=c8:(NC\_GbfgX/c4)AaMX/,Z?FRe(4RN_-^cW2OFC\K(
[<fUfPaYKd>g,^&J7G5I623.[1dLZ];0[/aQg\agE_8fT_#f^>6?:6ZOX>A6A8Re
B_)S=UC#/f2GKN/PgbZ6.AMB:2,D0:ED.I1P=d[aZ0TV3IVTP/e4=8(SRK@K,XD9
H6g=@U=aV)P;d?MD]0aTedEBE(T=</g[bX#Jb3&AQ/&YX#.,:9[bc0[N]Y10QT5P
=)B2RE^HX-0DX^ZXI9cTe4EB5$
`endprotected

// -----------------------------------------------------------------------------
`protected
gf]c;X)d,]I+_+VgIN3O2/KG2ESI_:f-BVYV6c6TK28@&5bD3+FI2)Z^_[A(ECFL
1aYcZKdH1HAD0E?A1bbHdc::+<LYZfC/c@=O:>B;c6]Z-X5E>a(7QBdC-G9OSW4d
=MZ__O=.@PEf0ZEKO7LXFF_8bf&gS1TMaI^MWB1MHE,UKFAP3P.[IO?HAC(HN/CT
U#2.f&)Z]S0=&\YAcN.g_ISQI81,+ed8;A1<d<&f;9b,(7?[I/@=[P.,65,O]VQ^
BEa](AD?e]S=.$
`endprotected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
-V.NK,Cab=eeN6]3Mbg[E3+WYQ_GRZS9aOGQMPb0V3@NY[]/:B2E/(d(:W^gBI)+
c=4KM>g:YE^#Q_;VdS:@Eg(bf,R:R;^+3(;(ABULSOCDV&(]Rg6244H^JA#-LVdA
eTPC(UF_0OR-]eQ/F=.E&F:]BCV?)/QbHMVQP)_^W7GfEaf/@8+NK^A.-ER3/C(N
Yf[O+-Ed>O_T<M:;]YcHWRSJ\1TJH_fNDd58(VLEfW#A2<MZccW7X@X<^2]2.0>C
ZJR[ae.3DAU[CWg_,GLb\<518SE(C,]:>UYAF-M[1#08PC6ZUXe7[FNOZE_5K=6O
A9DefO.V#^a^-Ja0R&];Z4U4YPSU;9>P&2@M8D2IMd9]T7>1+[NVZMUKd+,6D4P>
Z-VbW/;XPA22Gg.AV7PDaH/91J5DeFHE(S8Le^(e:<HSJac=AY:EXWPF7bSY^T3g
BW>P,=bD\R&N?5]-ELbT-aD/9UaW+;-8._/M94<11aS;TZdA8DU+J8/&.UX\[=>G
IKE9J0KV.NG_e(1#.;Uag9@YZ7GC4MJ;c_b^IAVdI\T&f[6aYH@Bg>C>I#/O?-JE
e])(W0#<#/K,(KJWc4#BY&eB@0EK\g7SV_f[DXS-DTFHRHV9:M0^G[\1f]/,(X)?
aEI1b88,;0PV_JRc(PbIZ6UcX)ZX8ETTUV.0T1)1Ze93J^Pf976#Q?:_1JY87;Gd
SJ=P#QP:HH=;K)ZJQSMfHQ^EgggHBc&<USF8\4e.0?GgN7?:#I3.S7-S::\:QF(V
?<L,BbLT.2C37Gf4X<MRc144g3T7/412b^f8;,J-P5^Z-36EeICU-#[Q5:dAYXa^
^K(0YbeeP&7UbIXG?@L0>1:]:/H2<:+O&Vg_]]+Y8=D6@<3I7V53#3ZJC.fBWI.B
[4;[Ub?^W3#PGU(ZI6T6X8,H0(ESM1:&#3PE9P(\25e91-:+_R1Ie9D([SDZS(31
cK)QRaX4K_cED\GW+YQQG6J)FO<Y#?:bfd2:XXcQJ)<gUR#8):K&bg4VgGZA;LER
^[\(PNf]HGL,EZ(;BYTX4,18ADLE/e;K^A_6[@)4?DDR^@Vf_XdHFC&:V:+;YQaR
ORMSb&O[^F>2[e&.VagOK[:^MD5B69O9gP#MDS>1YcV]+DSJP^/@=9D4HO^.FZUS
@g5.=g=gT7(MA=P5eaDb-C+I[O)([AaQ=441.fKgBP-5MOST4EEC5I@G:ec@&LPd
>0<,g;-X2IFA)?a[FMgR-\;d-P<+0V635&<fP_=\7=)V,=T^N:6^;TB)+&IM;Z53
B</=,D+8&g\[@-Y6<LBUIeE=I<&c0H7g9PHC_gb6XSPd^LP;-a.aC8D\6I#2D2[#
(Qf1UGE<+^QAP]3cYSd\51JE\f9e?bB;3^8UJ](>NcZV22)KTIc\-M5Vag]U&^(c
-5FUHX-?85O3>)1E:6LI0^JZ=a9<X-?+F\TcYF0+\7d9C#(;8^5I-B8D=[EK#Y,,
,]eeX9<:[ZE2NV>N=\4SNd^T7-0[3.5.ZdNC,UG,16L<OZ:7WG3TGZCfa-=T)>C3
e)P?33V/e3=KE]<Q,ZM]^:6N5CbYZ4_XX9LMOB7[dc0+N(@[Z4.X71#D9]N?Q&Wa
L:X\bIG1WN/9XVc;)0,=,JO5bF>c]C-ME&<;-\OM>5VPSP/@,VBG+;#I;@&+,>a)
IH@AE<49LRDUBS(BB799c8EK7O/O.>PAL;MU))2X)1X#V_]:/#:E,B6[0A<361D2
OOd/efJQbH#SLKMW>dE92+FDEJYW=V6(BM<6A40@.@(Q@DYM=+<RWRIcL<5=cFM2
M=CHcC[^g\cC8,#H1d#FVFWR/0[(9AN^L9RGg.8A;#JGZ5F-D01Q/;=?NTeHD=6N
bYgXXc2=gK5XOV:a_fVL9(T.1?Mf3C)@5NW1MMc8(:BPe_?Y(A6LUH2(@5Z?,C^(
?6[#U]-AU6/f0]H5O83DP13?be5=?0>)PfN#DYL.U,]?)D,&EIY-fK&TJUU0FX4;
OP6H--YNJ+cW<C+5:D<XD=]9B7)0EMK1GOBeg>>S_bHU]c[O,4]GJ6]HWC:,a=/W
3V^Aa;L\^_VN,1BTU6,;dNXgWbbQI_+[.Z]ZFD1K>[3(1b5WHK\@c<9PbQ1[K#eE
?^4G;M>9fO/8g,#Ag+X;=7dfM(>SKD&07T]c+_H]1<gOWPZTVUF-6GPN++-bQZa\
T>NRM(-Je3)K.Z\8f;L&#bcV=W[BT_Nf+D(C9FGCD4[Z)_51F.+=J9]//+d09D0:
J#]cdSLG8VNXa^D,-Wf-#,B5W/XGB59#5-G<[c.aB7ecADaAHL(.T#/P0Pf<Wb0I
R\GK>,=IIKc^@N,1]E8:\/</TdRaD;VfDO1LLO3gZ[]=gX=<@KWO3bOSUS-<Y;T)
4-f5?+92GFb3E:@Z?#g=VaXSVV2?ZN[:I#48HRP)F3^#0>H?JG0Q5[3[NFG=G7F=
=JM=QGc/Z8(XD7Y1/TFVC)bD?aMg.>.Jf]7Y<._4ML4-D0>L_@+X7+XZ>9[?#gK.
]/_eAHSSK/.BXb;3eY2E+9JZEIB+S544<4975U-8VX8U#T9<bXFH;M0e66#2aUML
?K<B6K<Aea,QQD>/+Q,Z+Ha#:9PIc<]S#\bX&&9J=O:/9?d&^K@N3a]WD3?C#ERd
LRJ)ScK9TIZf10I;1Z#Q?5)V[@P9OQQd]TCH?AG]W\^N5@P5>DBOc9NDc0D[)Bg8
2\8_?)C./OG:dI20P@b,g/P6M\<CR@NTg.+QAM\SN]C+HM\M9S^Y<8&S_>Tg;>FS
.9Q5.gZ.VVK0<B0Y@/\J+V).JI.c+IN4gX;RMgRS[:fNFG>bCGEAeU)QZAO8N\K3
].IQ4JZ=:-RB/A]e7cJ_D.]X?8.6-&;&\._RFgN5V&Y+5.5YE2_e^7XCbDGf6WIO
+Gg:gMCQPC>AJA[@/-5,>OgJEfKWb[P.[f_FBA@8/_G+LY@_S-694\=^AaM7?-EH
@1\J5cE?f@f_4L7H2+fY)5QF=U^Qc=:L5MAWT8SD.AJ+[^XSbBCT<eY079(<faHb
b37JH3]8UPFJc8[I86S\?F3;DaH66#g/DPA26OP[<,dV+YL?g:<[DEDWg(M4HK5\
:5N7@NAM&8SA:HM_#NUYUU<(C:U(1O8dZSQ:d]E[Q<gd+<#O/<c]7Z:VCC(M];>_
[+BX&T26_Te5KT+C,YFd?5?:U8PT\Ee<7Q>G#DB16J[Vd.bHSD<D6RE,#5PX>I_(
>eT0d>N;_^N@6W/4WWV/L.UBR2gC2<CZZNfaP9PG3DCgUCVc/O23BN5Z2I7C.CVL
OW:47K6CNV,NV/;32+@PB<M>]_cH0^T5dS9W=d(WEfT)egT\:deK]T]L.\.:P#37
PF&f+H4MZ+GA/cS20(->0I;:a<&HYLXX\E12)\dN+I?U/W5HGa2+(D8-GWI@b)<g
2Xd&KgaNQ>ASY>83V0-#UIdGa_^KQKMX&-CN<c&c/\#F/>?MO_,YTM</fBW0UO27
PZ-1Q<Zg[a))B063X1P;K>J_/c]-89>W]IGeLc^(OXeW]fc0VFTV+GQT3Qe]WPR;
&DBJT;E<I)0/@287H&H]0#HPNg4dZ_._a]=&^U+^6>0B(NGE]Z8MAPZ?@II<;SF.
)&FLP^e1X(9=#S/MY\g-((;QQT7DXL2<]2/aNH2ETM[Cb0DdP[]V/;):MXa?K+EV
F0../W]Nd8.a2Y4J^C.RW?BML]#.JV:P0_1R,a>BbHZ-3_&,8N;_<WERZ:SB7YAY
a<OA<UYNHQ[Zec8?g?EBfET7S]I6>F&GI7dW6e]>VbB^Q4]+E2(FX94:_Cd9W6H(
b]JQG;/-Gf(?ST@/:IXR:_8Ca[(ab^W=MUbW#^NfE2Zb,].J\>V4157Z-R//@H;J
VCAZOV34KZgO1cD2=C)0EU-1cCcTB=5?XdEL?M[V@W,<b9#fU18_WFd<N[SZ=9Rf
Zaf?VTcWNcAR28=(NVgTLK2@KQ^[K]\<@[K6])BUX+,g(V@dL9gd9Cf?=dR&)X5-
OPf#?IVgIg:8(\3#9X<0;YV>([/g[D.VQD0@7(+aIIX/\@8-@ROOdI>Z^N]ZRO6\
7-F4?K(eI3eQ3]ffR-MP4@JORTF;Q8V]-=X[3C-O8TG1I\X@+;/Ja\^/Z59a\#LU
[2SeRX8>=dK]P3&/>,JRK/f;F:GCa3F(.=TICc(f_A5\HH1_:c-Kd-XZ6ac6-&Q\
/R,/aT2R[.A2Ga\UBJ<EG:\fIQ>(Y0]]<d#6DAWV^5#&#FY,UF)QC(I_KRgeP..D
O0.@/I[5eE5\JT(A?M9d@19<<6FdQd[g,2MB2_.e\\gTNLWMI3LKS=T>V=.Ba6LG
9IZ+OA_0g8;O^e-df&H.Dg+dXGYDG8+RX+:&]_7,WBeYWDU=d\N]I/fgERS7eT#[
CKgPE&G21.R--U&_.DB?,e:]QFTd2P]6XR5C&a.=9ZaV77-g\ceB4<UB\K26SCaC
=WAEfOA3dbYg.4\c3BH9C;PeXG[+@W76&#;OX-^A[S=>(.48H?LH[7NEQXE^K701
a,LRRVe+O5ef,I;ff(T1FHJb?c)S:A;WN[Gd9J+4e1@]^+8(,P>]\]fWa9>=d\N[
0f[1\Ia.3#CQ#1g#^F;4)LS4\AUAW+FDXY.SJZMGf3DF?OcXU+)KQ&Pg9aAd7O30
#N;eNC6-I3YRFNM5SaLL_:c>2fN>#9ZIBKOB7)([aU<W^:#CSB[H3UEAQOY+O8^2
g_f3c=XLM)79:1RUY0+bW8/EGIS_WM+QgK37)7C1>8/&;U@V0[Ff5S9A)6#PUYCe
V>eG6Y)FU,.(Y6JM+&):3#f5c6(LF1WSA;22T/f=W5208eQL<=D7f71F)bbDTS[[
-3^3UgDV:>gI,N2.U8M;1Rc+_Vb7G#N=NWV/bgJ>9GU@-a1gIdg3d^6.GNYJC.5;
d90gdX1f&3]Mb-3H;\Q),=A0[A\6YL<Ag>6:K^&f.+94DT)U)LdJADDB?CT<IWFQ
RJ7&B#,QU&##-7L(ZB@Vg3E^I^<HN@NM\B,?AdC.6c=0G3<CG/@1KV1Z3M_&(V\c
-.cG^4-_b^<AV9D5bM6[0YaKE@BEY2Kbb=EIcGRF;(7K)Wd_30DE[RT,dN>g^9:&
^TX+MS7,CY2D-HQ@g@QPD6f0CVMXT941_&5X5TcS2GX^X1:-=4;:G9.LXe)HGA]d
;[YMU1KVPa6IKKc)SOA&WMFNX=OX2(#V(Bc5I_)[BYM8^I@ge6F\DQVP?3@&/PF2
T_[[)47>Kd@a#,HY=aKEI_EST@(:_4PIa\_K5_K<HXg).(d&^gcfGAF9E<OD(T3-
:P[Q-[MYX-N_@bTQ-dR-;W&RdL7H0#R[09:EW9]cf22-4D^>H?^<YE#D:,P_PY)&
(=C#G=QL3PQBO^OI+UUD7--S.Q1E[O>V^#/[11fPHfL0aQMYGS7dMH3Y0adFbd:d
c/WQ)M864<G;dc,B)a95e9><g<#[BZ4>H[ga_MD3@1?,Zf5H.@9\Q)D+?)XdYVW@
9<^.I188RMGb/9B+bQ8+eH8B^XgLEU5B/Q[b#R/.aG<2f[cB12eWee6JA;FB9=]H
]0HOD2D>KC<&b,^[6?OH<2LI,CT_eAT;C-[cPIBc).<e-E,G)A_\C#GOHZR0&1G]
aU;aUG&e+K5gEBRbV=_[fU:6dAg]Y?@0\=@.FadO,<2f(MS8FVF1>(T34=UHcV_5
P]K.cT28P1G-23G-14])GS=9J(;&G20_&H51U+7e=7C[JV\)]_3TKY;C1Sg@D&\b
0gaHSW6GFfY0)+HOC7^,O[D.Kb@d9O4N+)L5Q.PQO?]<<B)5JTUO\4-PH_@3E>dG
KR>:d4AM_H@V:2.5B:eV<?FDI7fe(<@?[=XUC6Q+=E=-IJ+7<a_4U3](=O]@g-b/
HPgDD_+SU;[.KbU-.<]g/PMSP3c_3Y]eW>4Qc^<\Q:.,GE2QU#dI4IK/_+HE#c0Z
:7ELFa_1gQSg(UUXK?E&SAS5LXRR>3Y.8a_f)9>c[NAVVW0);W:CJT;X,d-8^I\Y
_,UC9_EJAAdGf<ZdIGcYR/G:1=2cC8G@b.cGOHA@V+fO)5.Na0Y_U=fGe;O^OJg#
RUbde_D7=D6LC,J>MXgg-Q85)@eVP&&/1@,:>DUJ;/Qa#+#0]0JDMfPVX^\/=\fe
Yd3+6FOQQf3P4YFb)M,O>g@c;e&\V(ZL>]<.;SXS#(b?28N@&(PS>,OZ)18+3\33
:EKNV\3YFNF.7[KdR+Aa_f8aDRQXKYOHIK51)bTKS677J67fOQ;JdH=:?0bUFU;(
8UT2GLJa;e@21N;IZR:fLaAY3^_,[]MMSfU=64g6=KE=0/[>_H1)O_aLbE#=?C?M
6;92;Z?R-;T6GQ6O5DM9EcKBb[.2P6U?3RNe3JE=9@NGCa712Z1f;#.b41@/B#UU
89_c,P0O->.Ag?Y6DbKQU:JcV85JN1W4>,\f[Na-e]8,ID[)[P@cQ29g@;\8M)E6
W;-MMf<,T^BC/JRY_-0bFIKPMI_0G24O[eWHR_R:^G5ZY@D4T-?\(bSU;95cXWg_
_(2.HQb;0420Q2[K[@#XB?K[PK3LeSHg-L#&HHEeE@//BQC42M<#Me=bPU<SR&7(
U0,:F3=GZ?B3E>@R(3,e6<JN;T&/H,NGO?U&5>KSC1]g\g+BT)Q@^Q(G_([eBJXE
2JdW628=d.X47RBAPQ.U_e7-@+IfNKN=O(1d]SRVZ#8Z?BZM>7ae9W<BO,4M^Z:/
;JTM5:G61cW_H4Y=27Y>)(?_+b2I2HSBd2[V0dZc_fN#c[(F+6FHHL&:;;1Y-c?;
1964?6:27I[7:7#]8X+;BHd2.@#.YG7_78ffMS=eXHP1GN6\H2S-Z#g#7ILTRAMg
17[#K24L,OB7ag-ZUL11YW#W62-48/G^X89XR@V&+#OP8&B,N>:VN#J)gFEE^@/J
Q@R10UXNd:)SD0D.TWW2Q;.fg0N#][6&IVA@GeDbF2PRNEE+]g-.A]D;(Z[5G-DX
GgD:[.JZOgE37eIg:,BK]?g3EN:V@DZO67[Q2^??3G#T@FLI^;,I\JH,f?D&0T?@
XL)gG?>C52P<=O1;\_>D8g>W<VJI\eN>7/VL8I\M?6/4:Q6X&94E\Q_7?E5JY[/P
ZKf<9e4YP^YWF[T\9/9ZQ97A&S;GJ/;>cc)#R#):X=XD::Z]KI\WfRQDQ/+CB5Xf
bOD/=@gZ_HcYZc?_E0;<UVU3^P9R6K1753<S39RA6J0Pd\N;@UA47?N>83c(9J;D
e6O3O<R6&;aZ_X9FE8-[F3S3#dP#3L+?M@53G[XD]\V-0HgJ/S-?CNMPU<0=CRT5
X6P?KgG_CBS&,_K8GgB8\=]U0L<KdG,@.6XcM8gR&VOWaW#,+N^.ZR4=Fgf7_<VQ
V[32JbVYBRN<F_Y=6TS2#\YA0gC(eQP=Q4=NA@J5.3X/cX=:TeMTY3N^CQ4C3YZ_
;\4?8N7L4a3T?/^a;+6K1Z+V/=YgYM+@HAOF;G10>J>:5P;S7R9BDTI\8JEC#\g&
.;U)GPYZ9@+R;E/gHK_-eDg+f,782T7OUG(0T5H(;b&C2(?FOQd5K_5.3^=&PJ5d
(+1F;I0ZBA9<A=Y?)cOL[GWSO\PA2Q/\J,b[[3__&;1a>CcMSN:eM/Q-AffV/OJG
(?eITH3Z_ZNON:D)9++:A@^S\&a8#2<=]9)5Ab(^LQKJQ.g+B<B=KL08He250GK<
-.CR<8/Ibc8SOE6O>5(Q96@L0W4Z4HP.CDd&=cdVF5;>(69]1Q1GD[X0]]CCPfOB
K,1@#D8[AbQ3Y2@H>I?387JFJPV^.PQW,EK4e@.TEL+a6g+_?,\3dE=4;)J?#8TO
c&Mc3#>:VH&G(-2,K61J9D[#E9PHXf#WROfU<<9;dZ]Q=[R^4\G3JM&/\KA[:JN2
d,P,e?6,4+Xb[?]A;&G@0.(cA[M=/T7^IeC?]AaJdfRfCXff\2\bPX0BLPdI963c
?^9b3b:c;XQP&:NQ(HXCG8;6HK5M3VQW8QX-E+,b0()4?&6^f[&5Pa[#<)[<)f(d
?bF4S1f(2SPH:S9L@NM-U(/Ha1YIS<e^Ye:5;WMS)R(1[6Z<2X@K06:[.98FfN^=
<E>e6V[8L/3\NZ:-b#OGH#0+Y)EF+E_cW2QBbVFZJ&N^QR\,TGX0F=?7bgg^Le^)
^HYcL0N=WQ_3^,MJ6D/T.^Y4]-(7C.7T\Q=>)C[2e/KF;H#/HDHa?5dC[R<8[3G)
U:a0_g=,I[gM5MNR3d>@Q/ECF^#F81cGPe^?F\8,^3C.:(a/X.NVfIaX3]S87.5U
@TBTF,8HUFT?b=<_C&>c,GEa=YLLUJe5EY5-d45)+/c#,.WO_Td(\GK@R@CB3ZM#
.Q.4b[+;Z4BW<?6b5F+]b6H25Dg-9e3(TZf\7CZR]TRJ\U:6>?^V<5B2_FJUT]SZ
;e.^7)=+,0?UT:R&Ng>7&E,:7NK0Z82:57@,>1/BF8AGNAKS_RO/OK:\58T42[XY
D6P-O]9cXX[A2-HSaFg#FL=NNF9JI<eeGNN0_]1]0,X7\7:)>=>S<bA[C=;GKX=_
-3e_\C7(9Q:8/Y\/EPY#F/OH682C=BXV^KPH00;OR/O=cK9XbXVd6g<1AE<Xc->=
W4QV3OUgX^_SaSY)P7&B]ac^K=b^PIB.]NcGC__/&NHLTd_QV.H<#77XGgaQK5T\
e]XNLY?:661Rb4d=RL:+5D(W.;:.Y?,M_]<+3[eb,BSgdHD#<SMID24g4-XZ8LI&
S2?d.UH9?-KI)Qb>TU&8<4aY/\]aa=c\0LIP@/]c[gPGUZ9QA:P87e#QI>#/LAHQ
GM=eX)WBVd#1_8G>^4VG-J76TP.aE]/d-f<UC:X(c]<_RUP#73b2A16?H21TMW5Q
U&0-e3B^;B+Q+CaHDc&[GPRZ?J,HQN/dFJc)33K=YK70PWLYEFW&JH9fP2CF5-@4
eCOC8/Og23^\N@Y64^BYRQ[HI+f]7>K8[))C-Xf442K((A_GB5+];:g]Jd_UgE,f
<:3:&L>=;AVC50W^B>G[R<ef5<9QY02XPUIK2gSH:;3G=dC>3[>=:23)ZU5#bBgR
aI/))X7egJWH_?E;:d-#PO2>dcZccN.0X7W9(H\X3RI6:2)B&[;@RN#PY]ZgaVTA
58N0ab)f).0EPNY3]&dN8R4X81Y-T_-N73.edS0:?A_,L3KGKY4O(d0L(R0.GVYg
V784=OVUC#.+_]P=e8[a<@OfTa[VTN+<QUN=5[ZU\O]XMJf,JNV(GLHJ)P\E8C?@
8N3I>O-&WLRb(G@7Ie#/KUXV-[X;=K5H\B9Z0SB[=X]c@6,,<@_#3S+@f)^_GPI8
A1:8N?MEdW:T7W\g5/EGV+ITTY]4N+):V#+aLU=QP7f][Ee)DN_:9dW[X5IV+QVD
30Q6EU(LP^Pd]5P0#K0(;J19>X:5;cLYO/@?9fdKT=L<[6GM1:dKP:L6?SP/<(Y4
JQVKC]4@>c]_7X[e?IHINIY7O_+/e1RS:JIYC&;9Ie)FW0Og#<8,Rc9TUYRSI2]-
fB?V[S[#VI,-,ALC;QXBR&1M8;<IMXb@3Q4(5ceM]Kg+f_g>Xd^LMfgGb5YVI3gT
>.([L0WbQcKfF[8:[O)6ZLGQ)<E<cX[ef0[/H&._1gPYJLYO56e]Q4J[^c:XS/@\
4MgSbJ<3H5S0Ad)_[ebS,M:-+<8[M\])UNJbR/CYMHL##dO&46V;XP&\;#f4?[AS
2G2N+/LMD>;-Q#,,fgY[0?BH3@5Q-Hed-@E-,G;/7HLTLXYDg7]5#dMUMA60gFGY
OACN<^_^9]EIP=RU:Y_BT0Q9-?I7\@g;5^_H7\WELXU&Yf_V^@-E\=[EDTV>cHNe
fBA9dZ0f;Q+_#PR7KZf8]PFC69-R+6EE-OG#WYTLIg7:=0I0&U/gf293/.A4QB;g
_8V>.ZFF+0INegII<;Ef6X+2-@)PV17MN?PC5MU[?RM\L>1SLa)&\f-=2\O+96XA
SC4a<[Z4.YaO.97I)2;2N#MXE>@X:\).Jb77Y02TFYfZJ6I7TSY:U33@BAAK.J@8
J#_:O,6N4U&cI),Nd1(=\Q9W-6I^Q,EW\3?F#+@:VK&9#a&L37#H&G,C;9WQ&R4-
UE1Hg2>U5BIa)L-,65@E==;R9SU\^c-KJ)93_76+[\2]JUg4JZCRZdF/>.2EdT9E
I<NC7B3?W:.<_J[;gWNK07c)I1JZ7?SFaS@F/.#_E^#3010g.eVZ4ON)1YGFE[71
4\IX&Z<XDgSP+7ERSHOFDZ<CD(F-PBF;7GPJa;RHF,G22a6U=ZNW?cK07GDc[#UI
c/V&;8309#eCZ6350K/@,@5HNP87aAcKRJbL0/[JS\NO_1:AZLGIXOBfF?VK&4[I
d=\5@.4Ugc?g,)(,/,_O(fMdaf;/2<MVP:Gd0<ESD#e-E4fRc^dXC_JK(=4?7bWW
N@@Y-91c3K?P4fHK0]_=HSFKG1eH(&O018cB/T,H[8W/RBb8/#(-Nf&[U.UFZ42[
TA(_:GJd2Y?W;AWGH\<?Od3d-gO/B4?R3?Z_bI?L]G@Qf+AR:Ag8/>6;T0C?:06@
8,5/?N/;J+<G)dW9?G&:)_0ag2WC(VggUQUW23@.86SeTdGT_977A37BBD<4\CZ,
X<a-\?7:;S>ALaC.XFPYWNBbX6-1X@1#?d#aF)RKDeMb<YQR=eW_S?\)C=NFUD4>
+aN=K0/YD3?a<L,5D45Z[Sb1gYA;WdYCZf0T\<9;5fFU@MHPL38Q4;NPU(9\,E74
a@TUOAW^X]fQa9ZMSSb2OVcF[RYdZcb@H+]2_AE-Xca\>,eO+gAfQfbPgD4bafee
_5YbAd<WGH#YV==/gB6??CB+;K#V_2JFQPUY>,)[64?>db0f[5;P-Y9X;L;H.FW^
18YV@Zbe#-UNWIVF&,4C-9)a9#HB=[^\:a@7YO6UF@FD4e[[//6H##5.d>&<0aM7
N?aEP+K\K-^d&d8NB]R/Q4W@?]@(_Ge\YXN5W@O@,VY+E.Z,gH+M2H&^32D(.c78
Xb;2G0_>cgND/D-/231JeNGO]9FX9FR;H#?M..=^(-T)K71KP_M6J9-4bH?BP7J&
CY]C7/D^g+=XdQV]U#9C_G>&@9@\RMgLLJ^FN=7\0Q[e/ADdS,T\]K:V?bKUO9B.
RG3;CD56:UDM-E3@W(VH9f:O7VN:N_ES]7XJ2GH3S^+]-EO:aEUa=a&HWb5Y#@(G
Y-@(CO-J?<VA;])DA#^70,4C6_/Za(1HF9Ka>A)fO&Q:8XeRZ_^dN9/=^C)DbMa9
MJ+d2XfAeW]D8_cYG(5S+/31[aG<7cHd0S?76f?2Z\&;+@.Ce>YSRRD3dERH;,C(
g(^U6BHD/;E>#0@d.II(d2f2[JV]6ZbT4F.g^[0YNDc:gM?[JRWP)V)aD1TeIS[S
Q3fRF]L@G0UFP0(MRHT5?9,J\F_3C<OBLDZ98F0&S&GZIKQ\O.G;?V.PD=AG[?cD
IUGc]Egac0CYQcH,6IDcg/Se=&4R:(B-f3a>T48\&1L>AK[,J-BGWL5/]\7^&MEV
Q+B:(1Z[JM(RPZ]eLG-)X]7[45JOWX/4eS6V3g?4c+;73LG67;JY.RE+3J5Z@4>,
f:?_L?Z8(YDYA^EXOT?.WYK92Q69Z\#Ae]A:(B&J?)JGQ\fWP&V5D_LFYD.a1#=f
>^79<]WNKH>[;O7=X4B</AD;O_d-Pd/?-ReR7W/J^3?NG45G,e/]#63FgT9H+N0&
<ObAIe88G[9IO3L);E0g&#>X)1fTD(F&Q:K+>/X9\I:,+F9)fdZ#AS20,H@4Z^Lc
M\F^71;73)[QJ7da2cY70JbQd,Y3)_6NO/@9.C47K/3e0TWf+JEbE-BdLKYgZD3V
aOO4UN[XUcB,/1M[eAQ6/ZgO/.b3]YQ]M@-aXT0V76#WTDV]Z0+R2TeLZg?.QH-&
f&f=QII5.6eE,/V98&J6?2\LJRTV2UN;;YWX^KMBJHeX0QA?,@FV>X</:E::T^7f
?(d=/?JK,.dd;XE5d2D>F-5WI05ZaADUfJCVf\\P;_U&-T\T7O7Q6&[JR,XJNdQG
2ES2(BX5^,af6GCL3WY@g]AAY2fa1,RKP>(V.]4:cOSX)?_@FI@3)Jf[>ZE:G)F?
M,/(Q#W-XQQaQO&OL17<,^C>RcT64>XJRL:L2W,^G/b5W@W7DXQP:(]>0FH\?+aI
BCe2<d:+66,a)SN<-YZ[Y,@42c6LC.fdcCC&]=<E.;II>3G-^)E?@O-J0]H>eCT5
0V0]EEGf?ST#Q51AQ(N\:I#IH)PVL=^>RaA\[Y<Y5LXV:U4L8(Wf?dTO;.><J[FA
T]DK_g.QY>,?Wc#f&>+832P<^7M,Fa0bXVW7.4@88HA+U^C=:1CQQ\<Ye6cM+6N,
\8R4Qd)6M9e,=Jd#>)aA5<D+(;#5I6A4>/5I[[W9QAMYbeFL?3&^03W#J3>5D35?
I7AN>UXT&4CS<RJ@]8<0]@c<9&cfYG/HEFIC@TgcX>]AR[GJFA^@fN^H[H]/_3Z[
8>CZc_8aV\Qfd71O5HS\YBVQ0Z#a<Y+2JL2;)O.5Me_OS2KF\_7<XAc0[7a)&>Cd
]@7<SJa@+aF-T-EUP<W)?+66Z5WOc6Q:2K879:a=fS?eObU#U@/@ED[:e)^LV_Ob
[_-^G+Q^IcCK2MTR1Y;_[,22HG)U7.P_K+Xg_fNc6-28Ca(M&6b:b6/d.^I\a6YX
6:Z]?,QMHFaP<_K\/06;VR29#-E<-0?7e?Fd,.A1?dOB0XIG8BB@L57,H+OO6NQ8
S5+R56E(M.e@-GFS>]dd^aNASO(^:-7E.V+Ka4H_OGR)\(0PB#c[\gGMN#AR>\aY
be7NS]@Z\ZAae>KJdC2.U(9[U_SJ]^5??D@:V3(.+=TQ5gf=M\+Z_L;Q&WY5FGNF
.IZKOF:YKD>^0\T480(6YW0gS):-)STAQF5ZIH;I71JH:R;=-LI#3#ge?K1>[aeP
8)T6_\Ce:BNQf096D^2+_Y>(0/?O60D64TVXKbS5OfHP&#a<5<.R^Y5@\YF=//]A
^gC:Ue]LL34H7aDB>gA?d,H<IJ=P\9,ATQLZOL8A@@_-5aDHCd;ef0BWY.>SW1+.
AF0)&A2?5M>#-N]aIECHZ<F3;57_4<@)3#9^cQ[eI>I:/4=eLG))g@54)+_O41?Z
b,H)TJNZdE\+Z+LKS=P/[,ZE009Pg^&6.@b53U>0DX==T4X9UZ/Z>bRP.MG1OE68
M[QVCJ8,3ZAcF.UF.O;A27f419G6QUYTXHcYG&^AHa^JJDH)09/FXIb6g5M8M>cg
[O7@VPU&UQ)[Q=Gd6ZN@B8?9.+M5;CQ^:5(>ZV)@VFKa84<_Pcc<S/E_/gW4cJ^8
<VK9=FZaH:(JX/=+PZebJQ?J@^A4^>DE(d.4T3g45GO(U[O:W3^?e1.T#17@gTLS
?H^,dZBO/FRFY>5XTLT23:1^1AGIPY.KFGC:L;0>Je?\&<4/a>FRTU&g@O:E;W]_
,MCLJ)WC7/U#_3@f1^,3XF]24b8C-9>BT;)6\8F0QB4FM[#[9322ID0.20:_UN50
:QN(VH7W)LK>MW]2-;J@<aZ.A[+>VK]EY88XJ9D4^\7XW7:#&]H:Y,51Jg)A0>bC
eV[859JWU]AJ8VD-dCB8)3O(SI4GM.9YOcMIYA,U\3b?R6AONb@M6^-<>K0Me#<2
KdC6SHSJY?;RZR4\=R5ZE5U2:5J@=/QAYfa@daZ.e-I7A?QI19@:2O9^:ME3f2@H
,IK_>QCBO4BXQSYC\MIZ79:.\AP#0@1C^)=7@Ba\;=WAP1+:K5b;/RWLJ5)9V+Sc
:9^\e@(8-QK+_ZQ7TCCGG711W[g53CYB=0CNTK@:Oa,W)Y0.E-RNMK+S^>>=ARNQ
6gPID3E5=QT&+H[_U_<,=NJ:ZF2+Lf1gRB:1H0LH2#NJXP.LWNcXM;8Fg+2gQg1^
O>TF.b2G.#L&QPYPcEHJ<<DFVfgI[/e@Z#ILJ&Z2_f6e5#F<YS=+T+HK<e0I_+/<
#V0LNR>KRZaOHBBJD3UIL3)O5=YfT0WL(ICb.T9(N;/G]^J6QRGMB;##0\ed(>>W
2a#ZFE-7SUBG<e<d57+?HL#2fOc],/J1V1:V:?>]RIJQ#RR?YO,]bTW^JYg1_fM+
50.fH&(^N)(7+d_.Fd[@L+J97HK.X(D?QJNa?/<Q3+#e@0DaGYAYWUQS]cH>+g+C
@@I;d2/<O9,e63HD1gU>TW<968NWP7e+6R0KW>,=_.CJf#Q-FH#2#AWV.?+5K0fc
g:L>TL]<+F^O)?_&3YMCQR\;T=E;&74&)INA.[](RW/cU^7bM1cdYE9/Jb(E7(OZ
b@;Gb(M:HCgIT1I&(a^SH4KeHMV-P8g/AULd;^>WWJSZ^@H1<&EG8@2P@fK.BG+J
WWZcXCK7BZ85@/\2SG(eG.V5G[H:TBJ\>)cV5g9bf#Lfa<PGE:YQ.aM>)5HM/O_+
cI2f:#J\VXL4gZZIL9DOO?.J.&JO>L,K(T<V(UUEA_OD4U(Yf1X:^:=.VEUUee=W
BZL9:RaKV+,MWR)cU.#^Y6A-dZYDRO\FAJ58M6g95=[@4WI_B^2\SNI9aB-#OAX6
aPE_4LBZFgJ6gOO519TQ>))XZN(=P5^_^<58f@&C8ST8Q-V2>_##/(D4CL.&-_Sg
:8RB&O>/(V\DA[@@4,fXS5(<SKNJ7]F(S7SP0VdN_LY8^B;[(BBb1X2Ng7]3>ObG
BeWB[]L.\C#@TZ4LCTP7UCGJ)U^I+^I4#2WO8dI3XO))0&aAZ7BbX@]5ZS-1fT3Q
QPTNF^U[&E4ZNdU,<;./&ZHVdI,8_e[B<.1#c7)K144I)=A4]4<fVb0O2fY.V6d0
.Z;R6#H+/#DCJcc/9-W5WBP(]UAD#+\K038&;B:=(ER?c+6,PR1\>5>//O&U2HB1
LBO)N)c<+E)F4UPe;^).WLN&5D.RD[,CbcUDZcfYE;Y?5XX(ARL5/_0([H[5W<fF
;HRO)HW8=U+H^GW&4L9B?;bFg)QL-=(BA46GAc+EYbP:4[2f;Ka&)TJPZH\<aGL?
a#^d:1M\M&VP@=:K#1<].=cS9(.<B;PPKaBYYf[>4Y-/FHeT=#/4Z,#ZFW;D9AUL
YY-@fTF\#ABdAM91[J<0PEc<O..RQFQDTMV@\P,=aYS^3aE-7aE7LMH/aCJE</XR
GI8KCA<26G4D0cP+2a^JJC/P:]NW<[R0,G=Na[&ZLD5=K&Q;c3-E]?5Vg46;K)<d
P#B2;ANb?e?1PUgZZ=WNaJ<PIZ6BL#M:Gg&)_1M)&I1V^CR@#<UQVQ;W>TIYH^ZB
L:=d[S@>>AgQAUX)JO_5G>BNZ;b\GG-V+WLQgU<QUfg]F[A#J?8Q)(,:H^2I9&gV
Q[=/N]UFYY-W#87TRB4;Z;#WUG5J#\e8Z2bMM)P]SMN.EC)Hdcg?7^KSF2=0J;dg
MZMbdIGQD84K9TH1NP:^2F))JDML15JgQ:Yc.H(E)94^9JSWM#J&7d_HUB)Xa2IY
Z;K/R8XG&VN;[2,0#XNGc^7:ME[#)Oa/AXQ6F_^&E?NNd^?2ZQ8WTH6(5Y23>Q38
.JOP;(\eLJXGLES[T.c3;EbB0V-g3)>&::C9#^J)Te5I_P&&5/1>;(_:3Hg0,9Mb
NN:BcPY?3_JP[DUDTKH<)aWV,bM_0[2?I,^</RFK:T?aQFTO-PTEYg-\.2RYY&7?
+aR0?_<0E><[74(e_V2=a2+bBF2beUHN/\1gS[PDWFcaV=EEV^9ObZI)b_0E)b#d
+X&7D7:;e+FLXd.P7<>Yad#\D:gd3Iff7I<:./DJN=P=64P3+aO&DRcU>/EV-<JP
40HT[X1A.8+^Q/]]&=U15?,Rc3@B.W/MefRg+1U@&]PF561J&P9G<J,D/C1-#=NJ
H-.-0X/9;-bPF,2I>_Y1[2_0?UEN::=3ZP-<E_5C@<cT#YgC?/_,9K_B<-@O&O-?
eHS86,8cWc\cF=[O[XFU)JBeXRP_(D]KeQ[bB8)e]^F;-7AVK=Q:=g>P^#0e=cM6
Y9C52MCSBU]fZTZ&f[APKDIR,@<5[T@L\99084TALbV^aWG8d[f-,Yf(/KPX_@__
;.eM9=Na@8TgEA5H.2<BU][S5g<NaGX(Ze1+HUF48<H]G#/-^]U@^fJ42XTI)8X;
Zaa@.9@T[F;5H@?D?2#E\cT_@7CSC&86,Gc;0\<bYF54Sgf.dZ@>5e_1M4A?33?S
QIY4G.FAY3cWVY>5X5UA]=&f;T8PZG[;O^-K.:cH2CO3X5MeF0-2NB.^6/WBF,D,
Da+2CMQ>e;2OV>55]CTV&3O-@MZ3_da.N6)9Y&d>>(.B9;S0T3T(Q?RL:K,D))EZ
6#5Z(NH53(R8U0cN]JV-#4E9/YTF5P,K4KcFNQ3(>:a9R((g0&Q-EG1Gd.A#f?[M
g+/2@:4.1CL?Y=KRDX1IQ^,C>NVXcYd\D8^K1^T2J8SVQ_<gO2/&R5#18/=EWMa3
,BILUW+;A8=A8Z)#dLVgg1.1O]RWE?C;,TNgSC)\a16T2+-ZEC<UU<]IW1NT8>fL
87D?T;]?Q<QCLV4M\P_NT_.57.229M\&Ra7b&Y9,,>_5RHK]G[C::39VWC6KYOQc
K@gRVfMWKgV&<Ob1B8MK86V<G\SWYZOEU#aaBUX:G1WT3&QGfbK5L;M(GE6&F\U1
K@ZJK5J&.JYaKVL(M&Za(W)bT]/<F/d\>WJ&F_5\b8KA(#:0T+LV(\Re0@aLXeGZ
/_&,[4;eK63O<?a/^:E.C9HJB1[#M]_?2L<//<ZRgN@?KKZYX<TM<9).J\8TJ<e=
AZJaA8@JN3S7G21ZJZd^<gB[G&^<UG5S3:2E^A^]&gWf<BPcZ06@4([#d8Q06b.K
_#_S:;:,G/>XMda_^bT>PNCN#_1>CC#8GdZ^gAH97aCbbfL7/+2;8ESVfKD<CZ_E
?fd.Y+Z#VgE?3_B48RF;1&6#JBdU:[N)])6O5YRE+JP8K-W-J@P-NMI6-EOLR-4b
cEfOCS>SZZA^\&1Y5>c_D0^cV0F=OLE#b+7[Z\F1GYTe+O24:F@>V9P;dJ>V.(\P
+.WV?>RZ;YT5OF_Z2PS:Se]H2<bG01[e9,X95^M14-R8>C&@OYJY>MM88C#b=Z--
=G]H2?3U2VH9Y1KGFX9^c2JK9LJ_Q01ZP35G9QDPBDf^d9/20;gK?YCL8Z-Ib8ZK
XS=V/ECdK6&>X4X(B.GU0(5:3bR<CCN(7)35MSZ@6eOPK4F^@DCd_UJfNE:.e+_5
C+ag=\31OROT_4MFG;@&g(ca^2(.eK2_2BL#-\147?9;^H1<Ceae.2MdWR#J[<M5
](3B>QJL+d73&<N8RGH5LM4JI8?C2VWY)aT1U]@0VJ]dQ&-,Z(d#I/fH8Pe/5W=A
P5C?S+8&EcH+X4DS&I:8AcX321PS&;J=D5ecgT)63+6M<O#A(]Y>+>(?L^3YFdbC
LB?YL137+0AU1Y+=cY+fLR981Y5bTC_^e7ROVa1C=9XT^XM]X3(O&Y7-MK4fB.Z^
T8](VD_6&\KgS<X:I2.=\)5V_/GY>D)fNU85H^CY;7Q.[IVG2N)._2VIW:FPcW>;
fO@cJQUBX2#7G+OX#W>)b6CY?)Kd56V#0:fJC-;.M^UKH_7,=1eXN[aTXeJZL(;D
N96,YMeY:2X.;OZI=(1OWV5H2>;BJg=^4THg:V+6c#@DZ=D^O@@a=G.G4\)0<I)G
DA65ZT1+H<S0f(DZ+aQ2NeAEAf\SYH<0cPMK#F<?SQ-5(MX5C9;M<#VJ8@Z(b_]+
(]Mg3VIERc@gK\QO_9U4cHN0;=AH9D],306P@dHG-22bCKbc?N(3S;-.T,,@PL8E
ebG]4Q8LW-bR^;#A7I[YP>5<5@V:8DXN:M9B6;43DI;/XW(L+ED2\7I?@WPHAc8>
bQ(^#_Ic3O2Wb9#R7eJ,W/[I5DC>/NE\ZSZ)T^E\,N,LZd.SG4U/1OUZD?V=-<YG
HH:PX<9K=aB(Tf>a=J9XA&F;7C>cf@T/);Q&GFI=YMGN05F7P^-fRVSWcRPCSR5e
H)2U+^7C4=?3PfR=L[MA>J+Q1XL0:A4YS)ZSZM@LR\>0>UYI\RTIeE#cfNS<^6@g
+#RDQ()HIB2Ng\P]NBWXH<PUCbBWAN)4L0<Q1a@B#WK7OW#]RgTSDIc>Y)9:B95D
#2]G-U77e/8<WB_SYT0V>gJ:gKU#\g]QKIeJO/WEGe7.&7;NaeJ7H<6ANFKPM)O&
#;XH3\8AJTXR^W?:D>EN]cJWPO0aJN?R[QT1a;FcJCJX.6YQU]9a[KLUL6.U(\LX
_GY]S##+F>I_]ZWLU?.IH(g)I7UC_D\)RL/3T3KL1Q?bScKX;1C,_Xc.=U.Ob6df
?@-++?Zg7.PEC(SP3NA^PA0<96V\0)HSFN+1T.8&G)U5K=^X=QQECZYE.a1?Z&1J
AU>M_JS6LD7OcR.=W/.<(=g]W9ENb4^^bR?3H&)5]L;c?,W1,.NU#QLdK<f_.,:]
/fR7=I,3O7F+Zg_.(LQgYH)P5H<c?\TeJ[SX>Be9C;PBg18Z?O2);Df3Q(c0c[0-
_>fMB]PRe@c.QQR)I3/QafXQCZH]=-/+A5:USR.a5=M<^ZQ<QO;>I;7+d2C>TJ(_
PBAKc2S^6V;L@VbY]&eF@W78Q.]bK?80J(bA56U/ZR_c7,-8OJ^d9MA7Q-S1/-CU
f8-T5CYQcNUU[6K^f?,0b;U9dCb#N@S9WRW^KPJE/HVM+K9GK4deF[QRE-C-HJRN
Z+S>d3GOMV7_1A]Z;/XS>0dXEJ>A-cFN3:R#=Ug/g+16Bf,GTg:=&&P0NM@,#I=.
HXQIb?/7W0Yd&FIa-TgG@@7>df#KIJXE)cHg:6T?A/U[8?LSAOe5A5b7BA;<;[;Y
\H>X?^OZG2fKO78;J9gO8e.GG3M6&2f#;NYO\V[fI9PG([\6EFaXLUKJYRa7TZME
/TAB5R])NT5&T),8Eg9^[eKMf^XO9,eOe0MIPP^Wa5Ye3AHID]400SBU#,0EUI8>
9>&FSJRXZ3V,ZA-e2K>aU6^JQ8EW7Icf:\G&GJHFW[S(X0=(S@)E3H?[<-VMUWN3
<2ZOC#I[WU]5c5)2HcO[C=^8^7#,7Z:c]5AMSN3PGJ._?GM3AE3ce<2YX,3V6Ub^
V\(V[2.,77F3<YK9^a<\)]0YJd9IZ@DVNPD?B>/Sa2R_Z_[\Lg:9HE:Bb-Ab0BNF
(>BDFb8db4/8)Z_-cZHaS=aRg]Cf7/:bLQ<<^4CWM\6=68/f5Y.=Dd>;W>35bNSK
=[N=057]f,RSPB:]5EdD?H86dF&Xc]dT-1T5_J<3Z<-IcA7b+3#ZG:2.9Hb]Eb[J
SgSA>QVSONd\ga\3?,5N.J,8O6OfQ.cfUIJRJYFe.0K+6HLEBf.@JBb:_S\M+ga1
MeP<WHE7^02]MFGC@T_;ScMK]B^eU^<a):b)b)55?C79d_TWK5TU2;(IPCeI<GJ9
gJTIQb4&I6B^\K4F)Z?X??#,Q1(I1I74N)=WLe\JNcbV:c:_IJW0a>TFVH<2H6NW
:VV,_]2B_cG((IAPd3\M=J&cOB78aM;4P0W)?K2/3=:)ZVORHO]-_c_F7L2BQTDL
AeQ9KJgbR-5c>Z_\X9S^\SLXN4Df;9XaIa+]eM\Z(@=]0^)4AAF1BVP_G27b>TDN
R91M\>5gC&1O<4SNF7RGM)J5Q9UfG5a.ZX<C8e<D1H#10E#2E#]QYOF@g8bN9L:2
fY:F^-YY0,KZA]B[S=N>=I4eBa@=75;LPELcDE6>eN#M6O_cYOZ[\&WXH@,9OP7S
g8fOGY&2)gW@-?GQ:/DQ7VM-Ga;>Z(?-E[^TU=^D]-3,.>KMFNG^>Za>_;,MD][]
ELTe\B.9]XA<J-g76?3>Y\,-1+V/?Ya^:[S6Z-V^2]@&VF1#4@HF-[dBD,R;:-Eg
f>@N&P#T?ESeM)E?I#DMH(G03_[]V^RCMJ.,0@1bcE0[=D)/S^aWW>g/c(U/5BD&
4FZPT,32Nc2=C&1@XeB^<P&I<S9H[C7WPC12J<&W0KT:8b4B.4]Y?-C1b[8458YG
AW5ZO:?F9_7c0F0P,]N-3DCO]6R)7SJaBc,A]DV;&^7P3?S97]@gC7ZADAP,/3?<
NZCc/D5&D#U<QGG]R+a-eaP+@7H)7YEaULHU>WDeW^FG4b4<c(CN(@A)fVLF,6(e
_C08CaIBb3/V-c]P96R1X^SO9.PQJcEa1[N?2JQ_K6aCZ7,,+G^cI#.e8;gD+3bb
3A)2.9>X1gHX)@U4[a1YIEJ[.Gf)/A@fQ+6KK7KPDYc#FA),9B\NY-K(M#(LQ;b4
#00=(MdSb.:4Mf8S3Y.;8WY<>3f(RYVXc#?.[CLU:FHg/?0S-1X8&4aI\QEDCeK+
,?=S0;4GJ4I0:S7?M;T/U5L5Z?;XgY[X:5DM1)=E#.>#-&TGcDD\@+5aZ<.,P_@X
fET&I3/)I(Od>-Uc9TK_cP[c(LMZ,HY5X?-6c,YWB?#ff.N26I]-N^P;]>B+LNZG
?UO7_34@U_aA\[[CXdHL0^A2+Xe>dJOZ6Cg_&<MPSCVU5.GJ/4cX3Z#39SZZ1P8R
E<Y(3Y(H?BbNZFQ.FIeKbQeGS;R7SO/PDaCILUU\T8LDKSWaG2XB,=&bOU813GG1
\_+A@_-K?UYT?@=9G_-L9Z[.b,R-_Tg[-O,F^?VV-^V+#;N?eJ=<.G:?9[d_D1OW
Q(77RP_Y,YK-g2FV4E(^AHg,<3Q8(E,?9(+;M5EEc[GR:,WUfHSN-B\MU?cf\P;a
E>2PFF.IJ+<C6/d@f&dEJ-g^[CG,NO\XF/dP=69PI7Dd5;7S:C1&eT0&ITH9(LR\
Z[5])bMMPHG6,27CZ6eIaQ7^<aQ=M+7E.?OGH==>Z-I@bCe?R6IaKg>NTO@@(<C/
#=fdFc8We7#fcSB>CJK1_#HacJJ^3\J#6I5M@>W#]a[[N<YMAIVZ]3HegE=E?]6a
N#cC?dL4VZRe+O@,=?7:O5[IE+^(R-;.Q@)._-]W-ZA6dFSR3/^LQ9cVeTfQ\OBJ
VTV47(V=,#aBBAQ:gO4>E0#OJ>=8@.+I63&I[N,JEM]YV;8@T4-\_6=?e[D@7e\=
0H7c)R1dX0SC^BVE^#P^W+N55TS^D76?Q65/)AL9&cYNCCE\21W\6\U])C?1L5>X
#bX.BLV2<SEVW&MZERU35Red+@ffe?19(V\@SLKSS_X8\6cIZQNCJBDB5P9NBc9I
43>@8WW2JPQ-3UU9Z5JF3V)WZ@NL/2<._V8G-g.^G8&O5W/J:gUS^J380BR[(C2@
IBK&aYF^&]K3K-JZ@1.VaT(_=eLYW,gfZ=L7&7G5J[2&9U,Fc\\5TY#F&a@5K^U9
^LfS-R_2-(gb.L#BE]C@B)+ZUb=1MMFb5Va4&2CTB_S-FEU1aW.bQV-VMFaN)K,N
FR8+]&O\-FCKFOU/4e[XJ]BU4ODUR-(U&f.1_#Sb^B\IQC.45+\_W@[HPb26VJ(e
cCJ4F0d?P6\M053A92gS.8[VH2NaVc,eBRN2BMUXL(.,6M9[QCFB^A1AIPU^b1ZG
0E_eWRM?_@<5gaK+=bI689V=RD-50TM]@e.#G]<7_B/M79.VMM=\)?8Fc+6EZ97B
/9WP.#+W8PQW#b4AWWf[;;g_BD=R+VMf)CcC7M:1V4fg1FNB/G&-45PYXNF8TaE4
&=VKBeVUH[ReZF.eHT1N<F[B0FQKEDAZ4([U_I@],Z<EONY<]a&-=;3E:CeXRZL6
(9\U@f/Q>\S9[SgOP#PO_.]Xaa_W_C[KKJF6d)2+]d^)M3DC)9[A_;>+Z)V1K\Y\
a2/(N;CaC,6fW/L>2;WH>+:BKJ_^]S6?NN7+2Z1<bY??,NX#^><P.>Ob-@-4JTaf
bJT-cF/6f+b11L<56/cSK.72Y_]b]Z94M:G+12SNVb.#f=2S3fDR&daRX]R4C87G
_A2@a:<;cMfP;(bWWb3+#@<0QSF2K4^A)9:Rg>\>QLRaM)B]:@P[<a[V7E6Q=>DV
B2:a\N)+gN00cc2:K;6]<:_Z\3BQ#/JT<US2SZ4G:ddY3?aE4A+Ed,e0_G\XJ/FV
X1.NMH[Df+W6<6Tc1L/O29WHU[^5ZJ#6?gUA.;WZ-8\XZ_Z3Y?C4KaSVbde,LX2c
D#]3:G27]^EKGXQH@g9GS<?IbO.04VE/D[aQTSGHB-NU+1X///_;Z&8K?0VQM3/Y
c_,Y6.TS/&-+(YK4)LMM+/VTPZ+J_bYWUcb+^]bUf2ccP)LbgPP7I]AZ05V/=/@+
fg3E4:.<OZV?DgfF[00_)Q#<RDB\0?8_L.--(6;e1FL:[O(eQaN)+(J//C[.FU>7
(CZZ:SBF1[eIG+(f.KWDOF&4L@C38-a]8JCTK^7BHVX#DF4P[BcF?f+eG:bT<IKI
482H=P+C:#;5N2(TAaB(40T@0)OKC@.dTJcLRa_-8<G9<URf^C[ff?G3.<e2\.0[
Y[3\3<]_L.(A(.dOdKg<[CM@Zc^cPSWd0Q6;S[\WP0g0<T1CcGE>.TCN:>+VFaNN
e,6EQ7)J>X0Ua\^e=YY-SY>1<BcSe1J\b#M?H)RFOfDSU)+fHO]9S3F_OLRG@I(2
gfH\PNI.&.(9<(US<CJHfY_4.3KW<C6+XYY&WP_-#&=]]fdb<.YQ/2-LL2DbBWN0
.Cd0E>2KKTcIfd12_7[-V?SbR[gSXF&]71^BX^J-JZ3F1>01PBR1e6-M\0[RR;M)
NF54/U\:\0Sg/LJf&c,KX3MY>SYVd]8U8./?L@P9)N#T1;0D6<98[>DWZO3V=FY9
2N3D/D,-BN2ER@<B<6D3D=M]>g\_?L_5YC]HMCHaIUD2F)1=6W5:/\:NI(Zc];CC
>#M8?)@Rac-b]Zg0B#WXT[G&@1c0_e2.NIf[=aB<(?Pf?0fe_cB0#&-\8Z93SGaF
[AYC]O]ZgI1A.60G]JbAeg1cb,QXSc;57@:J7QAa:I>7fFeacgcEUV/43N)Kd-\>
b8)/B=8)#LAD?;f1STZ4e&Jf2/H:L+IWd:gA8VQ1+:I2dZRM/8[.S/1,(>Y]&\-?
\)AEG>?\aWb;LbYdU)57],Kf6Lg#X[]L<K>AVaB@\U?^J_HE3e4[FKAS^eOKQ5N/
YbVeN>\)Z@2PdCJ6.7SRAIDJLVDYaIV1&^;EcH)MGa,1f=5+CTTDU?W:2,G3a=6_
=L0_Z[cP\WfC6&LH&X^#9\(]7511CMZJ9eNCcL47PHRNA.<)B<]#VT0=QgV+5,GX
M[0Q8_FaLDP_P.36)UW0&FQP^N#-BedBFQM7^B3A=g7]VXG@U_M+AEJ&g?-#;+-Q
+,e.^>Y=D>DX4I,=);3,N7bg@3d7b9[f5R#MBVb3P8^_SK\N@GZ&,SWXSd9UB(MO
=\b8/?>>#7RL&Zf)bPIPO=/ccJVT^CXR<KeS1/NAT8>\g:?F9<>Z.b_>^=FgZKRS
)#84TaQ7H>^<dESGZGC&DHD1BCd=b#aV+d?/f?^DCH1U:bSUS#QBT3T\T1JT^c1G
7]O.8bf)?eQZX9PS:T\-a2c,\X(@+?JN2A[LLD5Oc(KAeKN75g)W6SE3<]D1e5[X
OT:;S@dX0eFcb^RAVET_0M7AIcZ<XJ:b4Ha7XgS)B<-,#7gHZ;HM?YZfXHb<;W>+
\NHI^O2E:8B]ZV4<7KB&].SK=A1EF>_X22;A_93:JZ_0B&5P_S=g5.KJb>#22[K>
XbeX0)OQI&K7.Q.=#S4PfA/S9D-W=.HW[FcW#(DU4d5#V:W:d<[_cEXe=1fG?a&^
Z)c7ENO<M6WW)]60OcZC#)e2bgdID#^F5_RFVVXM:U6>b>XWd(g7dS^]3TWX4L_S
F?Q@7AZOK)ZG+DdSf<aFN_EE8#Z1]QOQS/PL[_D#FM)P-,2V\L3)ZfAH)L)(5<D3
J(TQI=1ZNd0?YJP)IA^J:4IRUYB/CRWd222Y11/ZLJ-;I4f6PPUaH7bFSRFJe&,=
8QH<8)9^2dYceYZHLS4RAf&9g8^<X.M(T>3,e9@3K+DM;A)0DN=8_21XB+7@@+.@
8bf;8KQ;Y2@Cc#/&><DUQe?K\SY)(6@c/8D5H6eMN\(J9@bN,<W]J,B&AOA:5MAF
@O-IZ&gZ=[FJ441ZU;\#5Pc+(IB74Gg=UVcEF=U9U5T91XX_c11-LIK[QLI<3D=f
JV9d:.>OaOAgGV&W77bJOQQePWM;,f4^YGK^UP>W,/?1^>/=>3:]+RXK;d,PaG;K
^@a_NQV:Y(d@J3W\@YP#IHMOE0ZM3S[dCCc#?U^_<2^+I2dRC-26_>75PNfE0f__
Q[>A9fK?IZ=RGd)a=D]UUOM]gM&0UV3L.(W6+]630PS-Y:e\9?L4\VMbDQ;=6G44
OV\4VDa\fcJeU>4M5\D.W8eGgWaF#6-/FbV:ID,<+3X-4aJO2c:6UK<\6FN\>R&)
SQ(P;SfdM5^<a[MMR.V^>15(=/9Gg(()b&bZ#25;WV+_=7PV2f?e01cE8+8HN;G1
2H8R_KF)F<)>cW,g&5]b88fK;,0Z=W;5/4#T6M:H-;.>Sb4Qc_d:SfS;)DC72LC/
8<9Ze,6XO#34A_[N_1Xa?U8O164LUL[gM+&-E54eN?PQ<YDF6?9EEX&_<+Q/BcWM
LUEX=UQ;9e#K@R<#,&..AD>>,bADY#VE#RKZLeePF,,8.<PFbF2#OZZUac^NdEJC
EA)([c82>4Q+[=4_;DF3XS:-0L2MEI8:SMRG3FUB0X?KDKA5U9GT_NU7eWHA4Fbf
RJgG6aJB_e_/>>+R4H;)4LWd@R;2c)2QcU?X(S0RgL=.Z/<W;/3=cg#aJ:e9STLN
]@PVZ<2+B0SI=eHZ(=T9;DV94bb\c4/>0K2WG064D[5Sa^-Q#eJEc1D@)UL[Zf2^
0E-WNA@^fKM>GSN_?5&,^8+4b.TP^1Q&2IZP6d=0)20SI[aHYf4#49L#b4>f_9Bd
31L?\T#2>2dcgBa)6N<&Ed,>6LESP>0<U-2/aUE:2_A.K9>5YZ7QGE6;5&f8fFB<
08E2Lc-[NAgETFBM6@4[f2E.<9e42<:I6CU@TLG&fQ0SFTPMc&JH^GSZF6C77DJV
Ha\9[I<X4Y_,,f(:+2NX+87(+adFOP.G5]4FH,/8@<gaYVYDE:EY\(-;5MILZN_B
H>/+Q3+-T(7E8SCYRY<<cP0-E9Bb[C&BSc:2JJ]/JMGOWX5?DS+=<IcXW?4_-VAb
\VQ7:52YOQ;+W>JBW<<7?-#.O@+f5;_8SNH12FM#(5N<E-:&TC_;]=/@4c2QY_2/
1d>K#SMgAI\[D[c[1X9N(\IATS.A/KR;5TA(0Y]e[F@JO0,7B_gC+I9@LEIN.6QL
De[[N?ca]@2Lc5dXfW=GZd7I0b#d=AfZ#eP]Ud<;Dggd<>:=G-XbHBO[[d4>_]bX
+-Ob?;XgUWU6&<0+;bN#POTPLSSI=3^ZME0,OKS\?RGVE9_[RDd.XT,L9Y<#a#Y;
NJ9N6@@IX-;S-+BYT0Z7:c+T/P[U<-ZG(X^BD0T2CHGLad7#PB7G4<K2If5dZaXA
#P<O9d#;K.BHI?-Z7(,\g)25[[Q>f@N^A\6[A\d6YKCM.VD.CW[)/))C;P6023a1
DW<ce4@2JbgTf?[\EBFJ2N,e[cMadPC&Sf:8)V7g(IaFH2U+3R,:YF.e-fJD(ZXM
<Y[3Ve5MWM/Sef-8S4+X8BNabK4S@+PRc-_N3_P+4UC:XQg,5S.[e[.d\05O=DT;
-W]6JZG2&_cU3V_[2_]X0NZ+4MZE:_:4PH&2De&MI;2VA>JXILe@Vb93BVQa6ULF
#=/Y&YPM15OY6aX1:[<XOBENFf@.Q58+70E/8+^g(&S2\0WS]=>@IUcAS_f]]D.Z
DZJ3O[#R>=DX#9YU<KRZJIQ@Q+:Ac&O,W7MdGKI./AEAI(L/9gB6BeFILUYe6>7Q
,HV&.XdKHBXS=(H3/8LPC/UF9,)-9d\6SY;L4W?#M7a.[+K)eR]c3(fD9:[?^N1a
\fGH_-?@7T#G=1&=,g+A\bI=3aW,6-d5bY_.da,3>V+Wg_GYg>W6TC8eb=VVYF7>
0RW3Q3QLb@E,^U&J<:WAaNT+;&d-H/XL2@2Q)gV+7^DKMB+I<X_:@#RbKfRRcRg/
<XbZQ&)873e44-L@?;]UbI9,QBD[Dg<PEVP^B2UJ?bEIbc66CTJ9&#bF@b?\1ATA
T>0@>D0DD#?G0F^a@6^W9=^BWdFd(H;X<1/2\ZXOP[M.JR4a6?00DcA88WD1.C]9
g1=:3)CNeIUZNMMY:,=.AJB(WI-RM3RLd:I\ETQ]3]V0?ZF)KS8BM.GITWQa,=gR
e0Hg^1.\:+--<.4WD4O+&1F:#>=MDD5]1>Z>8ggQKM>T,#.KR&?&e<,\Y+9BMcFD
(NDF>d\5DOHV2)/[d4Oa0ZO42IG<f+f0YU0>^MOC=/WO/YeD=R0VZKRaZ^Sc9/BU
bcX+HeHSTb)LB47\.Cd[Z3:BI?YD\UULX>Z[cF#))<1FeSUF:+W)DKL(d<ad27O.
<,R7d7<Q>&R_TcRYDS^Vae&P5@.cg)LS2IR)73L&D\cDL_2/J]a?Mbf8MY(N#JW&
0cGRM2NH2[Cc.&CD)5bK0-Z>gYQUI-5Lc&<]]56[T0f^.;@,aJ-4X]b:9+6e[Y_W
7R3\2-;b:IJa]^_O_^/23@;/:,Dc^BI33K^17A>Q78W[Vfa.YE=O_V3),TGS1Y+c
,<(e<a<c0MXYKc/_fM@P,eD<:123\CMB,3]O#):JGW+W8/W)H0^-+E=eCg8R8e\H
.<0R+BA_e;THRUO<8HU7;D6d1ZD;C,FLdRK&57e9eGbKDHd?QE\dFV0;b7,&R:72
ZNUOF/d0)0NQNSJ9AF9T[>YFO1GHJK=9V4bf0)f&SQfM3KG.eAe9,4=4A?@K1aAR
9-K.Cce[aB^4+HLD+Ya38SU(a:cIAde:Dg\D2=,)7=V[Ed4301a:+QZW=(#NN5e5
0C+CH1-(((_fF#O_KHG7SU7Z0^ET-c5K9,D:)AA=:@\a)\e8IbKWgY^(LM@Ve/PE
:ac).4RaZ(^&E@(NCM()0dU&JH[URW.0;YgTOWD#OEgNeHCP:R9VR<Q-^dZg5a(7
6]1CC)@=XdALHZ,75AQ_]TfW@gQQg+#UcLVd7+?30DM<9EbXbGZP,9+7NCWd?eK:
V;>a,D0A[&=_aU(5LY&Y=KLH6e,bX-Z39aQ(PgGXBICJ1.c+H>ad]]Y;eDZ?Y#;E
Q)X9XXJd?gL[/=SZ0625f.,86_=D<N<33a5+a;^I<@eXS>gIR7X&0GI\)DdGfF2S
0+QeHK=M7)2aE6:<3H6<HA^WC^d0PD3:fSFf^(V)0L2.-]84c=[cZR/gA_@H)_Cb
+e0U4QT-1YW2:T\LGFe35fFT6X_Xg^F/\Nd1M7Q84_#gS@Of(D@6BH(b&a#AE2c]
>F,3GAHS=bD^BNEGGgB_V?MN#JgX=Q#I6[=1<E/)UA)[-^6TY0/\c3E-dAWA\=<,
_?)BLIAR/(J=JA2;3LGGC6^)5&Q?@CFc=,==1GF1>@+=dCG@NG6;N\2>AHTT0Y1T
FLaBIMf]IWR^)f5?WBY/S80AZFA9L0^ZdDRT@fN9HYT/]M8P/RV^3K-1MI68g0,W
86@W:\VMRX@GdG8]4J0Wb<BL@DS0G50VHb7?,0B=c=^8eM=6D@F_d+,g(2PUZ#U2
bH#_8P/<ZbA0b+dY-0<ZC139JT)XJEb^/)H,I:+<Z#EFfIYP--E@:NQNf+SC@O8;
E]+:3(eXC+^/>U0baZJ)c\QCT81PZ_;Y+b=:AZd;-Pf#9KM;c.[+]JOKd/IEL1Y:
TRc;QXge,DGQ>#BAEbK;XYPL#f_7da04OGMV.)O:^,f)d+&#c>T8M^&f.d1)03+E
=AY#01gb-[CAGf.A[WN(S;K;5[VVcXT><dNM9^9@>W]Ud;>4F/M\B7Y:SfH9aA8A
NbX3TYA>[;<M,W:8PQJWGQKfOg1S&9J]LW>W9,J5G?Z1[TG>-c01E>G2J/N76=.+
W2b0>_S0<ISg<ZV-L8Z>WOR)(LCL:>/G_EfVL,)WSVRQ)Zf(/JWVaU][Sg+]U:H;
H<V@FcGO=\c;?XFWKV3FcMdH#E-fS@U:.CA><c;d51H]_Y[Z6YFf91,+U=S&?)UY
#9YTO.RB65>Q_/?>Y9PNQ.+bW7RQ.:E#P,9XZEX4XHJQ\acbe+MP:,P\(W:5b86b
Q+H#;<?IUJF[f^RE]T(SA-,_MfZ@8+RAK3B3Y.DR\[@EC[?eXM]L3[1]Me7bReBU
Z6;]BW4cbZOFC+3cC#W?f#W<QEdP)be;GfDW0[D#FCF&#C/)]8T&-=EF,O4<S8(/
eI<;(/f=R2]EZ6_]F&&QcA\CR-&,BF,e55/HT\\fb1DB;1R.S3N)EaOa;GS<.JCf
f0538-e(X7I_f[_cMb^.2&E<4XaUgKO>\=2DG.#Ib-C[HGZK5)D#aCY/.gWaQ=P&
K1>,J+>\NbDd\If4e.g&TN7WH)E=QO7Y)PJNQB+J\4F4B]_R-eO]A[9J6M\FG7_F
[gHG@LA.[7D#G,cMX4;I1K3K5A,cV8\CR;5<AG/:EAdP+dMccS+U#G+SI4:cL?=7
]d3Q];&eWR9^FKfb,RK,G#&2[J,MC>BQM.9XceVMPFI;,d4+\X?H<cT&?LG3F4b^
=2-@PTJ686ZONN(b/#;15\_2,S;B3H-0-]^3d5;\N10?8g>SJ.1ebAA130BdV8UC
[>2JM<>DF?DCYHX]#\ZfD&4bT:T.9##)f]gN62&4++EP#E6P<A-F=b<BZb<K73\=
=T=525,#1NJX356YY6fDWVOf^6D(ZW(Z@<)JO;aS4BO7gZ2HS_\PJd@V^a2c2J>:
F\9g8g=JaT280/IB:V.ZQL4A73RG3S5PON0Og(bLA1ad<^:=^PFbP:>&:WecX1A6
/We1<BIWfFTUESGM_=+>gbE\4-:W0Ke-;_V)cO&9>S&2VXdN9<S-eMc.\@NCb1TR
T3?#(8L0LF0E6QP9;B;Ja5KDP/+TAD8RLcJ6&/TVTgO3/LK.TQ15L=,A.+/)@45C
G.Rd7L<&&UNA-J/EI70GCO9/NA90H5+BNE=G&J/GK+Q42AGQSMY4GG2H<Z<gYP4R
QX0?R?YC,aBf8:<9)MMR1>S8+)=bHBGQ<=+a?cg5-;7Ng(g,BM896/K_\gecc[6.
G)/8,C(.TIV)Q2TTObM]&,7\3,ZGWg:>fF:M^4F5XRBILa;6I/Z^&)&3S?H,.aHX
=AQD^1[3[<e[;5[(4X0LTM)4<f[(N&J2\EJO.Y(5d=L7^5?2)L93QFbBM3;N?@C<
>9A/86]4X94=UUU#-S(#>K1JC(eV.+B)\I-(A15LA/]+_K0bNBOUNLD,/RESLMCK
EBQ(a^9(_N];WJJ-eNF\R)7EHFU<C@37@LFc5G3,@)GVY)Q6\K;d6a9X,bR]?\9\
eWD-eg^f9#H.?DG<_5SBL_]ZW^LGQ?<)_)=<,9(.,e^&>O5)dY193aYgb:W&VRdJ
NB0>d3Z#97C@7GZ>La]Y=XZ-LJC3S51NZH21V50?UB63:_A.5?,=IIYE85\=3@YM
SV675W952]Tb]8^YL//e=6e7])f7B>@b#@He(^4W1-Bg;XNS/5QY\b51#0&>-g7I
HD],BGg6M+L=fWaf7g63_W0U=@@VPa:DIPd;IF+PN0[RA6WcHLF@&dg_RUPe^I>?
ed?I(DZ,O^2JLdeYPKcY09[C6J]<C]aT14b)bF:gN6cFf45&2R:SIcY5=>,9>E52
Xe./F2O)G.\8+PL.W1M7[=?X/^><J]CQgK?56cR:5W^1IX.6=9X)]#=)gU+5W)VA
DO<gJAFaMMTV,[bUe+,5J&\/#/BTRD.-A3>b5O<_>8L#^M#,<aP7/P&-\d8D.LCH
GM_a_\7((#gN=ASKWQY7f)=F?H;d\=b_<73@A@dZSX7#<fQLL]#aH2,-c&\<Q:<R
6SEK.D11^a8+WZce5AP.U&A64@b0?cU,Y\>K,-c1d>..H03W:-S):>LDdP#5<&O.
dQMJEW^I[c-X#1>G8WZ]ce4J31W64Z2eU9GXS)\Y:Hb-&WL7<2RE@233=,4O]D#.
gJ#X0_#4KN[U3I,[gC:81H4>C)S)[N4eT;#:]@K<#<U7V7<Ye<S^QWNE^,8,eE>-
3TQ\SLS/3;+&E_LSebT5+7Q-6]+R-WN#83TNTE_(45Q/BG#69@R^4\JIT2,a0)<>
YA:]S-_?>MNU93aCHAaV&Z;JB^W2?3ZeFQP3?O3#,[-G,)K1YbbeNcQVIU)K4[H^
&9Y1Dcf<cUab1X@0A)RK=8;ZM6<b5BT5b8&.<.6+H0H6XQe924UUJ,S3#,T378b8
?UR\,LC4bE/&cRWE[HZ#S(KA9#.,ZbC?WSd64,;/cA-LeETgf_dZX3/KGV&aS+(O
.8L?]E#O+FGZQ.@D82@)?QVQ(;@#8-c-)WVgW-[R[fDI#F>G0U-I.76Q-I6.7,0/
e\]L=_\V:?.WL9_a?6/PA@.MS5/;\M\Y]ZQ)>LJU0^Ne_E6Xc?d2Qd:+4e23Nf/T
L5X8dVKZJOd,+UUOVA8LB.TB)SH]U100\M.0c;cLD8&V0Z,@T&5C8.R6F187)?W,
dP(O&WU0<)9I,X>S^dW<)GeBFB2,)]W)3>aDE;G+PaDQa+F220SKPR:G2BY5A2D;
Y2gDQONBPYOgE1\GI^L/1;B)A2/J.>>U<R..?G-G(g;ETI+a1&Yd,)8998ZNFBCC
KQ7?2MA&b3cTON.-09ePBJVKY@D_>>Fd?E#eML#)@^B0U<4+UPHBQf-Fg]YLEEWG
[RRGD(IaR-=/E?1D;=db9b5ZJXf/1JPYD>f#8>=IC2[BOKCEDX/L(f2[HZ3a?ZG)
MV9I(,aMG]&[b9E<4B@aU86FY@[I_1[[b[/IX+e,<.2f^A)^B&:YIGS?UWE\Ne9Y
a^/6IVJAVHGKDcFM5+;I<5c.VZNgI(5YH14CQ,>e0AO.?1>6W\&Q2YHWNE]H6O5N
0NWX7#U;L;@f#I#TT1(,XKe3K\?/V>\0?MR[(Ic\N625c7UcLX8<JR?.]FKZ^6Bf
<g^;W5(6Wg0e-KE_E\8LR(@+)5G<+/,+^.O&^#VFMBWY=S?e2d6+_bGb9Z)@7Ve#
05/C^B8H6WFZY8RZeW)A=g:3;DbcLA;H]+1I,,<Ba.8OU7=^07eU_K.[RULZXMR;
I-;#64CI#=Fd:2C?Gd0LMd/=)<<^=^Y8<g/K10gPXeUdYRabTL3QN<-3Xa[,JPX-
LDP)_VOLWO>fE11,+\[&5V?+(?2:XX/L:+gfGQTBHVf,f(JGd8TY_L.][OO&OWCa
.1Z4I[(A3ET/O/D<,0?Hg>29]f5K.M]91d]C;H_FQ2dR,ZI(M\)G5S^I]Y)-;#;&
V75JZfNb[<,Ad9[,d7&Yc)Q,5Vbd7?A(dcSc&XNW80cRV@N#YHPMA]SMJG+a73B=
?K-7fe?98N8/4[_]95>O?9E\#]SYLa:cVM0#RKT\.0O>IA)JT;\\(ZDTE[7P7RQ^
6&S9ODe^BXA0,Z//_)8LMD_P^b#7U65K,EcW?@/M<_K;I\G_KH[&K_JN2+JQ6+I+
g#MS(G_:8[<[-:#-OWFR+=eYU>bU_g\FgHU.5DMB:PMLHOda#ZF6&E>JVcd&RR0H
:ce.H(O&A[,#c_9bYgN<WKLM192E>P3BE8T[M\1NJ.;]=_H8>fWA4OWe,XF6ZRKV
/59,UC-_EZQ390fI-f4LHdG6DNJS:C^D.YM8f=A03IGC<WPNeW/P=/7>HF\NZKKZ
HBRW9X4PY_b,bfY5YcAH1LW@e,[,QT>Lg<_63\X4[@^=f9f,OW1_Ia2_gM2^\H=1
;RJfM(BX[aaD8O@B/WRWf@5IYCdBKT#YffEdWJAX-+eJAY_YbUgM:E0W:9f(5,T6
M+)>XY-260>B(fD,6,XaDSNOFaR#]4GfGFa3P@Q8A?Z24e,#:UC>H+^FYMF@++79
33:Z96?3MRd0=6.K,7N8OU#EG_b)ISe@OMWE(5-FM1#]VZ?O6S5O_bP+/<68dG=N
ZI>WKFDTPgAg@/.EaTRI,+B9,@Z:#G8(4^ET(<GGRWbVUWRA]&d2[c9aM:UGMYE-
X?.cQQGH#IF?+Q:GJ<L8OgXN5dZ]UH4O[TURebd6G;TY=PM+]=UcKP_DN,G])\FM
7R96M7WRG(g)J\g<<>TS(4GEI6U5A.=[YFH+-B1T0?dV2NA[X&AGZcV)IEc#ab]H
+6#BIALGK^G2T]V-DP0&>YQY4R&AbBOQR)0)1,2@-[LgccDQc\E\NEg<-;66fQ;?
6QTR?\.<OOK)c<9=R^#COK\NJ/Z3+g\AZ_8L&;D[-cVNWU]BQBSU;QE;-)#@/E]2
[SB<9PLUJaGKHNA2a/A.JWg9S\cH)MX,0]/LN5,M_M_)6-IZ-H2MeT,=O+Kd#T8>
d7^/0,E\4bbO^cY4eZ^4VdU_N=I^W:>F/05<,-\3?,>WJU>&E=PHO/TX]6&/b+5T
?I]0WLS1-@8;E@e[KY;^Q7cF\)?Tg^-YME.SfL:?LPD?#d#C844A)+NgI)H6Gcfd
6S)1TH+0WT>6#[[U9d+Y=<HXC\TgY9&OMR?/)YBHX)EUJgD77?+LA-?UC;89?A<[
Z[M4f?T3T[5I]IfVaAN3K_Q7=_.5P7HRdHH)dO#Ue<)OI]O\ZGE6=S#UXG0QP15E
2_QOfb]-<UgaQ63T?6:VCAH/DCbSgdI^7>6E/H/:bR0dAWZ8Q2f-+T:@fDCDJI9_
19A+Q2RcGQ=GAM;MJ]M2FVDC]7H@D+ZUO?WJVfA)c)X7XGT3P2G[<7,&K];S[>5e
-P_U<ae.D8g1P__b7g)M&3IR=bgdE9H3@KK6EB+XH+?,S/155=,T8a\O[)(^A[1K
_[:E<:BH>;abTDJc8T8JH;I31C]2P,:VebI5E+>5MZ#+\7&&MYVIA;Ief5,_82M:
^83ZS/PZ[/RcQ,bKGAfQAac<#)3;L:M?TG@99ZM1]eDc.M@GB^Q9?WG74VWf=EDG
ePa8Z;a_1H.+OL266eeb;ZXY_M=M<-e35-=2?3TPE,,@\CF;XBF@>dW05[1>[eQW
Zf>L.V?bW@^eX[.Fa:7=&@ALL<EF-;_=cfX\._K)gg;,H_(QeR<L#MDI_a/6&V9/
8W@?HF\N0K[Q>,3GaGI88bcT0dHB::VRRa]/b]T8#9@@,@\IR_LU>(YU\eI:UGdd
AcO-A/O^YEV1e^BDN.?3RXA.YW]O(J&/&L<+/g7<[,3_C-):<.eC2Y-Z&W<+?K5F
+e<SS7>#:T=b7[5PFMRb>7.P1XCPJ3T\.((-=.B77O5L<)__1BF0T&@6FEE\O1fE
Kb93()M(XdV@8dH5gf,Pc;Y@b-)c[b8K0>MM#QR,LYT8;_(da,f/C+2Cf@<#.54Z
75Q]afB[?O>)G>)T]I(Qf<(IR9^Bc#:dU1&P+UOD388&)^3?UZdc#d;?@@@VIRC+
SSN5.VK1660:XG0EGM;3^GKa#ZQ[UdT,#&+Sdc1/;\JS^2?QC:H]Ba)dG=CX<><-
N[R(3OYX2a&/G(1Y=350=34.g;16O]ESgM=[7/1Se,^0:e#P7d,XfX?+gW@VXZOf
)(R2-eKDO6[8+1W?2D\?BOcD/QGD8H2X7A#\3.@dfT<5N\35TE<.#\fD_/S8B_O[
53/^<E,&dUJ46Db<S86M<5&^S>?R?a&J<ELN\MMS&X6L=<K8M]PB_5:X-(-O@=9=
V8?C2&SfIO(L.IZ1U[I>6bZCg(DXHb:I0:WS=dN9A6+H[C@D._;QJ&EL&&]<=46T
U-93?b8U[RO4JCYQ[RU(Xd^@D5?Z=H=gQ/Q,M#2KY&TV-/1O8OgK]-PC]\O>KfEC
E8>&<::e.0,aG[8)aD7PPJd(E.9f#OfACGH.X4[g2\QXeO^CJGV#D7b>=_25&7ge
A2O>#BJ-LE_\cBDg8^Q5Zc8U1fCI9/]=/9@W\E[V[fJDF<0QPLZ@_Q4aDMf\?fFg
aYC+fP.Z&T@-aSS;BM)I^E:[^5cL;?QHIY9\AH1AaQNDB8Pb:Y+6.g/[9F^fE/E\
I@/?WFS>DVg[aE0?PC>68[D]P//VASLLg^VTf;CV(M(-[732JeX;LFHRHRR2e3B4
&&.2d,=1#30a&Kc.K#68fSX.+c[eS=UD2g<;g:CRd/MVW9S,Z9X<3^3&/_8RO#.)
+O24(=K<H(:D:Ncf3VRE:\FM;?a-E6>SebVOgU<.MPU]IQ=QDQ#:.dCe5@4X,e,0
C81R6EPV>+6AB>U4>?9X_b5S5U;H0=W08-W3+ZP]X8>7A_+(68>UN&3(\X]=e^f@
27_G/OACP;aE+W(O1FeO(2TF,b<4f7Y,c_K915^+)((B?,=3\E+]FA]S@6\cO&33
KF>?aba18(DKN^VF:]=C0>3#K[]+]&D18MF78^OUJDCedG>_5:1ECYE5-eQ(>@U=
IB<#8+OIR;?\?dXE&-A@_\)gbgLYMFT7=T,4ebaLc&>INZ;eK]Fc/0?GP)cA4C08
XV9IaB0]b8eY1>_ATZLGGe7F3D1-J=Y_#[4=-,1>feQ&gGb_3S/O>fE\+/BPcUK/
ca12]LE)[P_)Be50K#P1_J.)^_Me74\</c5H(9GEWLge(5@a8/gE0,DY#F]Q)G2R
d)D],^I\D@beA-Jb#E0+7&<Ef))dWf/gMHK//?Oc3F@NL^/+W9HCPbOA6O:Y>:Sc
f(,J/#_B+?STUEeYPc1Y/#K3(PPZ:Q/8IY44b#1PDM;:C--2BC-=3&&/P1g/bI^d
?)/VgeE(B<?AO0ENL9G0=Kac,-\N:VE&cLH;U;gf(07267I//6d,aXSR>H/,Jb;I
E6/5&&775c470GHQ3Pe5bJf#IDUaA,J-Q/B:e&.JC1],(ORg//0<B3RLPYg)Q,7C
08^[Ne9AeNBc.A]BVTfV,c0+XADQ:Te54=-1,;DfEF#a[+b5;R7/JTMg4SKg6&AC
K2&HW8O6ZMS/J;<NZKaY?.(Q)\#3NPOU5<IA]LB9)JOZSF[0fI:+1JKa\b:fG2S5
OM&8ONPY30WX+,gaBX5aXdU=E#_@133(b4:DIOH8>UT0&V<?<\F>:089M3Z.EEUN
U6,L.Y:4>URVP_Hde/M_SS47S0N5==?]g:?@:6/e)V+^VQE3gWW^ZMUKfT_\>f]=
d^2c5K:SS==B38HIQ#07J;C,P@V94SV(C-c<8d=0M9EXL:+6O/JL(L//RD0cU-@4
LNSc1U3U8fX[B[5GP7d;AeAAS]2b+ZN,X5&G[6X^40@1RGPVGHeG>7g9Ga>c/#aG
R+0Te&UC=1S&=6Q#Pe8UD&>9V.^&KRB,_T)4S47JK3P\649Ng+(A[28aVf3/=&>H
NW6;d./AdNXX)I8W#B^MY][,,,)+.@>F6@<:A3B;2#T;/#.PRUf-\G#7E-)dH0DS
8K8_+I0&=XPVL;P1B>0L2>S7+>2DF4M#70egN8IEN2DX<V):dWXQD\RN_1;JTU>_
Aa:^7[#C0dJaBMG&EVGUfWH&E-D2^53LX00SLCW4Y9M7T:KZcIS;>2[??AD7(H>J
G]:B(SgI(AT.b6&2EK=PN,&6M9>gC4H9ZFL3KGe6bacKRMSGOTcT<:W+JA(/&G-c
Xa(UBJg=/D.14SZ2KBT]W:&28@XH\:1AWNc14XMLO_5VB&78/M?-JZ<6<0^;+1R4
DDa_5U;5EbaUc6ge\aO5:8;b]TK=QH@ddKKb91OA9_gP[T)7gCe[IJ38V[_O)@2T
>;B-A^#>3(2F@#&VT9&Rg@=Gggb8Sc@fDX@d]a.K>a&Uc980HF9,R@P(8]]F3IY/
NHP+5<\X\8QSf5>.E4ICN(HPeK7;PY&^&MQL5U/F4^#(1C?G12X+&gb=K+2H(;/K
XcX+A=T?>?P]fMSM3::L,afRZB:.[^(fY2dG<&36OLIK-&N-=V0fXZA)R[TRH;.(
HJ6_8X.?=JOPa3BbYH5:baGFPeEA;2;c\L&B@;GNE\+,?M<DV.8/E/A)f7/V06]f
I((4CLU.YYF+/N8KR^QUY\BK^\PKb,b\C2WXg\VI[<(EC9B0@b5-B/\(=>YZgSB[
9WAXRNFH7UX6+^Z;=F861KLD5<g.5BT^=-?c/8[cW>PIH3Z.>J:>@bdT:c0@CKdc
Wd8S8>(942#//831=UV2;P9Q8T3>D4f#;BRGA]=CZZ4OIKZ;P[>cA.>X_E6DeY78
)7)b+D\;]eF/C@:7MJPQ]HICM2O^8=8L6DQ,a-SX^Z0Y\Q&</ef)T.b1e[ZEFZ-I
4@Z;89Z3C>-VYE=[T..4AQ=:f)N]#&b1\:-9PGWQ<O3W5BC)\Og/JC0&f3A:LAA4
P6NGF6b,OcbI&Ug:0aRIR5f)@#NcV9;-Z:POPP4(\;T5R6Z(_383?43T_3H.7c;L
Q70f\[F#(KTL:&a>bOVdRU?Cde]Z,RLF<.Q[gIIa-=.9>\S0(QR0YD?C5IAL\Za3
-]b;c-Cg-SU.CH6eM@a[Q?g=2NeNWfWDH9F&2(:9AW,-2HI2<6R(3JSR(B\X^]Fg
V1[2W<gC]G3#gX.aA^MgF=+(GT^0f<V8>FB29N[Z06PU#^[4/)W\?KMI&+N8UTP]
QZ8GBH-ZZ;Z=L_HTU^^RX1+OMNI]>4BXM1Y4^<YP,FEXSM#KH)f9=9W74>@?2CE;
P55X1e#]P)(BUXAS^?W(RECP=WEdRMNAOd)NGGY?KK_,g)OLA7,E]eCR[JCcSDcM
CB:47Q7dQ>C?fWAJY?gOSJZ[Z+G(bNaZ0D)5CG<9IB5D_M>^cOc?a1+bb(b=L<([
+<<H@;CF^=WVCg@]M1G[&C?6T>,XE<]VS>B.T^-)W2=4G^3>fG[:IDKU/N7B./]C
>J=GBR[=F552e7DOV.I]SgWb(93C#GUDP9cKE.CMLdX-)2NR\WGd:-4M8;ZP#PQ#
effUe@^&3P_AJ:dM+_OQd.YZ-egFV0+4cP5Wa:XJJM6cCH#Y0A:f4[?P;ON9X?d)
<:J_YPL,?<^S3UW69G(a#>ICT:H]H<a8O[<6Ac<bV89:E@b?U.c?dZCa88LJ4[N:
O@VgLNKRR.A)X\7?K\]9K.X3I^LFY8VA8eAF^6Ea4G4W>>b^@FA0+d:LT=0G7ceY
7_fEM-.g<9b51-2[Xc?b#[TII3<,37LNKW+&S:_L1(5<^D8gf7gIILF991a7CS7P
\W,a^E+R;>5H\6d8WQa>8R]?5V#=SeA<PG_N>O+)FJcf^6<H:RW0OGYFV1EbMQM#
AMbMG1VW7OW3EedEHN8F?J#O3],9f?Y\THW:7Z4>U[6c:E)4/BMG8)QBdG_(Dd=;
=T0;M_BWX6cZ6D\a+L-E#QG>)^.;a:aL(#]&Ic&;@EK8Z3>YTICF-A.L^f731Ob/
a1:O7_^5D9KeI6#BRWL,gY^^+2<GdE4=.LB)#aRHG/.5cgD9=Uf5#Q9>GeJ+,b=Y
>f&:KS/^S6Pd.9fJ6IaZURP]@)@^DO;dA:aO8W2OW2KK,&gLYZV=7CU/;+SOG3@;
RQ8fQ6C56e2ddD#GZYdPcEDbJ#+]N7][]IRN7E#PQ&6d,GaV<_+-Qg85e-Q\).cg
<C^5^_2RH0GE)PY0cSMFZ-OPUa/4aJA;V3HYGNX)MO7ZJGKOg;MZdQgP;Y7d]Z7\
fg=_BJ,.Ja:=:Vb=Gg/+9Ja8CQ@]18DCd49XNDOa.]EI7JVM4=S6:.-J7fIEELXM
c5[c\]7UN5Ige&gX3e@WDK,=0U@XfXT_cdd(==@)@AD.@^R#GS.+&U6e\Ag6=FRd
@35b8DU0Y9Q&I/NW@[FTX),V>4P];Z\)BD=Ya&4:B+dU.BOS6Zd-LL-2b860d9Q1
66+c0<PS9fVE)_]^+BM>_X-J9c<)RF0d6a:ER?=:59b><MJ<HSPA9a2ZbHLYcDHD
#0,8@Z+8M</&LdT?dJd:U@aRCZX;be,]L+R/f)3c<2;Y@6D[2DIdUd>?DE[\8<CV
L7ZU==C+97Md[UM(3+5RC1]]ID\.QISTF/KHYd])dIF[U\0@R\?=HBA;/P:R]]dM
eA2;d07/e,UZ4;Nd,_LOC7C/M[J[C7F#4[S?N0FV^fcSe(G]S]IWeD2M-(Z^Y-XU
Td+PRC^VS6b6\P3+e::AS36F\7RfK&-T@8/:L&28@80JL]63<NYZU/QTYQ=^1O52
B4J(DG)0cZC9R<E\-V7A+Q\;1Ld&H<(7.6Nd6V><1(cQK5M8)<70WK\[4A44VS.@
.JaHU1V+:bOQ:b.HQaQ3Z><SgT-+#)VBTNMLJ./I@KbLGgNe@/@J\#BQ?A1#fK2;
,JG?\@T9<+^U8K\dc83Vg,.K^&&aHD8U=,MZ2C&)dW\Q(TIO-ZUO57ZDG0SVFagK
:XaWS.#MQCN9;Pd?Q7]Q7@M1I=,WY8-0&c.LAE(@D\CULP1Og[0d49?X3d0_YTIS
20:#][Y-a81T2:(GG<S;]J?+ZF9S)CS8g?e:dg-L)dYfL@L-1;d:2ZbOU)MG>[CG
2N]22b2Tb_/:91.Z+FRTP4WCDf\Df@?NcA/A4^HaU\Y#fW8PLA(L/N+@B)B;U\^d
.)X]0YFTZR\B.UBBW\4?+(CIfB5>;Qg@9ZFO/_Z&AaBW(]NcaG+c2&.3#6f+03M.
T#9_Ge:4XH)9Qg91KW)6da[cL52L9?:QK/?-Y&@89;23L?Y7/SKdg.46aYId.K>1
5_<CD:a>gfPbFgJ7H2PQ^@I5Yd4M<MQLW[A)_>T=c^bN3AAK=@1M(aFc1Z[94fQ=
7&A,BMd.?5WT@e:b=ZD+VH+#TYd=5.(ZdDY>WE)C4W;ZIRB5]\6gN\VU]5gZL=GD
>ON_84EW-UOYNJ[ZCc>0@YJK>0P?H_<7AV7dN3O+5<EU?7<1/YOUIg)2JU\995O8
4,+Ddb^E/G1aCM0Gb?EMCJ#=YUL([:aC=da;TIQVZT6J-3HVfH&/dLN:YMJ8Q+DB
V,SM&U5g>>4:6E#A<+SJ_Y&bBB/GBQA@F=)1V#?Q.S9-TcK^_GBKZ6Y5eMZ+_5WP
/7G6;e-N2N.cZE)@FEZS3>QgHRaVUQ4bW5(X/,ZM_2DG6_REZfEH>3QcU(>0F]KC
<,Uf.O[Y<BZ>VNPg/;BY8GFZIU.WTbPE[GeeIeAN:4SMFgOJN)T+-.B8O)M/:f7T
1&.e5SAe_cO5DN).FH>6BEW@c4_\J)/Ya0J[(2JEW=c4;I1fd<3=FW\J50;bTNDa
/;bSA_(Q9c^(P4IWWgUb1R)=64a?>ePa#W?\)4C=/D;X(Pb2geD4cI:QI?L=V+7&
04KR]+275ZJVV/3F>]ITU&C&&XB1Q_HKS;>9\bEQH[KAg9e58:.>aSSF<YLC.a9>
fY99Q(VH^1PZRC1+=C+4Kbd&Ld@bE[PO=_IS:)N-YBA69/NZII6Lf\TKV).CG:#=
ANM/7aLDI+K6Y,J-0GKN\eZ=RP#F/)[ZT[?YFO.eURdB@9)c2^d6ZPD\\LU8PX#a
X_ZXg,UYdbXI&fU5R&W))VM/D^W>g.<02EK]Ba8X7D<-#GV=768Q8ECS2eMeXZda
1P4=T]JKdT2f^Bg[HS(O>NTg]?2^UHH^K(1T&=R6:a0B0];)JWNUg1D^865a[ZL:
\>O09+dFZ,SEY<YMcVa?:H[CN7e4+^KCf^F.VM/WTV),&S@;5VE44e&0KZ<0=>-\
60;7@;cE[^fgfbG;B.L=BP<?(Yd\ZSVU\))JJF^2\3AcG5a9KN,1D91g]\FAYaCX
g/(Qc,<G];+f)HYcb#e27C+CS+=HeJeOSQ5<(b(YZWN84KYbPV26WMP33TWeE^V4
0>V.T?;H#+[6b[-8Ta]EeD7_J3aF>9;EfB@;CW7/0<4P-TabJ5)g13M>2M2Y=(FS
QZ:0)(^UfXI;&A/&^HTKR0CEc[A-OGW6-+&?6P\GS&=;E5X,;IVZ2@#faA2:ZG@;
CDT5H9Ya0T6(^TV\Y[V,_;G>;_LVV=1,eI)SQUOML\--&0P(\Ja(KHOe-9B1PF&X
N90Xf^@VPP&575TfK^?g;X9839b_&4TC_+W(C.A]RZ0g_]dFBNIIPcTDPV@9d(Rd
HUdSYB2f3W_K4Xf:H/6,2GLH)X<Sc3Y4C,aCJ3)M2\&.DF3cZY]R&a\:7B]K0Xdc
a:8gT#Qe1]ee.&FK;-U=ES;MKAR3I849-RE-\&b^;9.CMW=2(/bEITJTBWC8.,,#
WX&23<0+)P4Sc#7\/)WdAC:6QVGM0@]D03L:[:S<FEP2LPXBC?,A.5e_7f_I,BPK
dDX:DI)7.@.e7C(+GP37Q=C^9_b3@g\NH@PR-e[A];2_29KUY:KNJG3W8Nc@]/OR
9Occ6X=M6:9,d>e-C,0_QY3OB._>\8NdWJcaJ17Z72Y/[LdQ,(@dDSf2CfY]Jc#\
fgQ_+MSW=OQ.[G#6VfJ/.4C#+7g2,QOgdQKeT)f?NOKNaE#7CWe,VF@,A<-D-gM[
NFH^DTA^C:C^81-SP3Ha)8H>R.e[1+cd6fAHLQeL&]\J08aA/K39F;0F6(K7PE:(
/a)bF(D<T4#dT5[Q+5_b;M:&&YN9H],bRJ\d[M-1UEY8a0):V_UMHYgCfeGeP<<f
)M\S>E@:/D=Q_2)9K_@3H7B:MFH=(,cLON4VVcF4IcM=+ac8T[?2>?IaI,Yb)G&f
/[1-YNL.-COPK&1V.\ZMEAEW&_IE[#T/=.eL8_R?D4ZX#M]TG;M(=-=+Kd]/LX_W
SX)P^fd/(EY-[F_A/)XKT1Mg93CQL#@;>Z?LB&eGL:d-NR-0>0dX=?_e,b,L5[&R
;6MQ]JHeW:#a/)^e6SJKPQ),I@1E<RH<77[P<M[5JT;N&K_7?3YP;#KDaW,H[#O@
f5#eP_..BK8LD]d#4T?FU-LF?DVN:aYBR@4+\)>F0[&\5#[&#T&Oef/KEG7Z=A=I
O>NIL8-JU7RT=/##\NAg1:.(;Z(JXdbB=22g5IY?8K@]c@A:R8W6:H^294/=40?+
?#0V0EFH4=KD87N0H;KM0+dFYFD9S3HM-<,-\O#EPF6-1O5LA]SB]O=F>QPO[NTK
N238/.-\E(E:T&f&I7=e_f:\55E)_#3716)dH[70Z,I_E(^K\J8ENA[D=UC,C1Ig
F]L17OBG/BS-a6g9Ig2b31Hb0>;_5\;8BC3D3b@+#)>F=H:_MP,gO;8#4O+?.IS<U$
`endprotected

`protected
P>\a/>gO,&@+QPReCX]W7[7f]&]U/5@P\5/G04OHQ6@(VG[&BX@)+)3:,Rb/+AT>
.;I--4AadL]Z5cV3KdMXgc7f4$
`endprotected

//vcs_lic_vip_protect
  `protected
MOfTC\FA?(^Q.2<8.QJ.0ZPS>?:5Dff?Z7P9d>(e-T).?deVP&H-5(7),:#JK@Q1
4A/1)RN@T:<M1>fPS1?YH:cC.+/5]TNX(\S<L<OCE)ZbJ(c0WY9Q/aO5DM3(JCH7
J4Q5dOY:IIFW\F#eZ@3D8Q@NfNb6YW4M&HA:M<VCUQ]3I=L@25LV@N]]5A(J@=+R
K;1CR3fe0U8T)(0MSaDLL@X.F.Jg:1=eXV+97R+Z\GCBaCXb?/Uc9aIME_5^9:BI
dM[.E;f5LZN0N-cA)07Kf[R3De>?Y\01F_J=ZR.gH9gc+^<RaP.7aMR=P923R892
)9:[IQ]dDQF9fJ3K?[-T3_P\PY-\SC>FBUF,5HKE[CSKB])Z3)FV<.PT<fZ\8@U<
G;M+)@e4b=Og?+6^cL)g&/bf12UF1Fa^E\;>4==H<WPTYL7>>B/[.VY@^,E;O>9Q
ZSQ)a8T6_cbTG&/6gK,NSXJ;Wa/D4CYd;A_bHLffF(:cMK:BUXeR:/7dBHF&=g;9
OZ5__&3e@11Mc11E3H0PBd9B/5c9BO>CCB#<-Tb>;/J6FBOe8MbfdO&TG/+GIQ,X
Ma1@aZR[2[C:..4QdK3FAOVB)Z/.P#3cbD<;C33&#R:56B-L7)P(PESFd5)OaOSP
JEI\#U,Y6W_4;Y\?8\<-cQ[a-<&-b0GJIU,L,7\H52\&NET.394WM^MfEIZd5FV>
>9dg,e&[dC1_]efNW^/;=R1SCQL>F:e@O\2G4SJ286(]?5NS^0_A1T(=0W4UDG3)
ZZ_4/XGd^@(R.(K].DR/[T36/^=0B6N@VF283fKK4E_)B80.OK4(E[=R+fF\,M>K
E>4-F>EXb)FOH[\4HWGO)_.2;/I1N5fE>=O2,X]TJ7[JGVa(e152Adf@fKB,_7V5
2(DLK#BTH5QEJdccK(GY8L7eTfJ)^Z8]3UBQgDHTP@1=?C4L<B#/>][7gfRX\[M#
1TXWH[-K7M\GJK-MNK#46AHeDN^XIgS(2Vg1:J&f?NdL7gTHL5QaX^9P29B(fFEe
,^255;ZUaX)KfD2<N4/D-fc7C4,U@=2=31UH<aFXJQE6I2<agN_bD^1R/H?VdV_C
PD-L]O-d4BSEF2,0g-###9?AZ5e-HCS?Cb[FXOQV@>SfX5,c0FZ+=.@GF\5b1YP8
S=V)D3MA9UXFUPKF4=KIb1b<JSAE?1e>N5TA9<c/Pe9&Wb<_\2)D>=.]e\<J=ORF
7SC&,0.3[eJ&d[THM[(@SaJ9eW0<L:TL)abG8NaWUIgLaX<5?@M2H9NZQVAg5N+V
gJ4_?HfGfReC_].X-g:@2V,ZZ=B6;@:?9_H;7JN9f)K@gU1,bQ@0eJ1GR)a3HT:,
eMg\4/I2geOEa/W0_H:?:R=>G?RUUb,DLPIZ1-X>[T==?5Xf@/T&TBN^NJ=52KS/
JBC8P/RCDWPKB>I+\35:IK=@bKYBJO]b>OXCeU=E@?EF>B8d:O.(^B6WO84.-EQg
YEK+^<>-\?)67>UJ4.5(3NPJRe)^0&B_U8UQbDI-S>&_KL\7?[4Y-f@I:;V9:RB?
?b:dYeB,Q/g)K1KcK]1P7EAQS^c5Z8:=VTf&+69DV\/:1(/0V]C),2+bWMJ)RdL@
V/F:]K[JNE+A1FVH0[QJ(0LYe/LO<Ff1f191R@Q0_T\RX?39TbPBcV0-14gV(<@,
W9M0>OU84[M&AE\MH@_XP[Z3HTI+T4]-V6^^)>)&GR[UG+QVI;Y=E-.,\9N6GG)c
g[ed:Ue,e>PG--fQWJ&:WP[<B5aOFW,HQZ8fD,T:e6EJM?a1[\8:/2\;[M[0Vc3G
IB(1W?d/X]8/>>;.==8G]>YeT6+d9X68C\1J+=)<+ST)gV_5Q)]ITOT)0G-@=B7U
JUONA<gKX@T,^:C54b74eDgD&>g#WW26@>X7@<]5A;BRR8YMZ:P=F3.fLF3,3PC0
YNN@GP^<>ae@7>ET23RaaIM_77c8)KO2bR=XEg<XF8M);adZ<ZLYBd3fY5A&\Yc:
QD1WXE&:93D@cCb50I=(6Y^+A,gY2GY/eWgU.1895/YV=R+]Ca\I,B8J[X3>^)8P
@OU#g0:g/YdORJD6:#JDg.TS,7(,(c76.:)#7AK>+8NVF\_HL)6-@0,-_XX<3a1U
JDFMEM@\Q#+BHFZO2[I]V<b5T.:440@3dd9H1HWT8bKd/UgYB]FVaIK&D5aa9dP)
G\NB<]+XQg7;IS,J88J/1/c/6(7W5Q<EADg8ge]4fC7-\ER1LSbIF54ILUTa/<LV
?@)5&Z^#CZNB:FIXYAI&1BV+IO^>,3Rg?+<.cRYCG]1]5:aZM8TB8^[Fg5:S6#;J
9;I=a-,;e6DHaYgHS3[17VNL7:#.]&G<ISJR+DI3<NK?,4Yb7:]XP-OQY(#;MG7&
Zc+ZN3J\G=-XeGaH[c_+I-)Cb-?<?1(K[#AGIO@BD3-K+1#)2F2&NL7-d,^><X??
cR:79YZV(MIG#>&V-g+>1BAQ[^LE.J,?=#S7B-,2BP_W,NYQCG+_@_GD^g#^c>WL
L:[3Q/WG=46RCeGd6+F1W_\T^aZgE^/]KN3.:-ba/XH47bdL@#7N7HaCQAIKH@-1
:9aV>e(@AF;KE?==63-KAbfW]?.0?a3@Z,GaBMD.aK5W4=8@b\VCBFO8,@4V491M
T_c,0VB22Z;SA0IE2Y]YXgN:F)a[S3_,C&b7f5cA\VaS?f&Ca&8b<13_O?M8=,cN
)Y6,FU&K\Q)F-H?\.I)@UgGJK1EO[67+LH5c1cY9M9MW#9&N&G.U-gA_OGaDWZ8d
A1c/-M((],QH;ITTSJ(+S\LfQNO.ZBeJ&5#?5cW<8Z/REALR)@+8gU<GbF99Qd+&
)9HA+;aZbg0/+C]:SUf.a_:AJ[@[7LN.BR9MRVB&R^-7>+K5BX+[)CRWgZKf0g<^
V2.=4);3^(Yf1WFgb>H#/?LVT._(@(Z&cQT]4KaF7T[\N5LXN6FF=,S(;6/B(&2S
S1H2gEU-[H_-J[LNa7FeC_I<ZN/Q.Pb7?J-TD[Uc^-A67C[=eFW^FR^\_E?d]gT\
7d,.eS=P]UJ>6RUU6@VcR&M9U2>_2B@d--0;2.dZQGNT.91HaPf1#P_>?1K>&_^,
H#2S6VZ:2TcS;>-gI7STIZ)\R#eVRRR3:&W5E.5_[UZ3a8KJ1eT&>PB@R<e[SV6b
(80UgD@1J;RL].b.\/AV?LDQ=DB>e&HARbB.DQBaB0ZT[Q;AHN?ZC0KSQEg]JI,(
4c53&FE=JNH[,2[,;J<CZACD7V.M;=N#=GK#b)?e]+6f6X22ZXgQBD7,>)#+.\.Y
_EVV8Bb;]H=9LA_aEDN9C54G)WT6ABG\?,J]4K.8K#M)?\&1J@EGd8b^Z0aDT]RN
].gH_?TfTF##23;-Rf(g]NEY[D1FF]aZ:31WW3A0&/.USR_76R3ARG:<-D-R=LN4
Q2E+>Q>XebT#0LJRUI#7fJ(7?],0MSQ3E-:bc6PH;A+d)3<FF,=ccZYY(&L-@TDK
QN3C@Q5e\+=A]JW=\?O0N3N._YK.d#N8&Ee=<TB2+fT5(D[3VR>g05HB5aYIZ:)N
@f;(fGd#Ac9)Tg.KX2YL^<KgJ7)(,W]BSEb-f^#B[U&P<=TY8dg9REe3Ja+NJ)12
,E4Y[Of1[G@DHgWa2,T]\B,b&?P/KL4HYd&QZ@@=.&)#d.cdDDE2<,).Id/CgO=P
UB\,:<?g8eR-<-BLeFOH1MJEb5<;LW;L<dKIU)2F;R8\6<8UL0#U)d_bHc6OI^SX
\#?AgX=6M/[U0VE+Z0=c]5XZ=AdV0YMf.OXJFOUQ&MG?X9LDF0Pb?f_f-97XU+cQ
9+GFR:.SV[G,8Z]FNL6WSP:MM?fMg>T.O:(H9)?^;E=[-3>6e+0E57FHK(SZb6DW
e^(-c[=Y3+O_3)HD^)I^B#g=RcI/g-\0GLZYHYC0>+WbASg?]IR4C\3\JQH?K/@4
RZ61(Be7I[[U>S8MFcc6-D+(&R;I/&O0P#?DC]PM^7Q4<96bOfT(O=A1bcS9<W\/
G45)O]WV20EY;(4.>Y\eeDAD^)a2LB<]XB:KfN7_M)4OgfSP<1,LQ98I;fJ-J@.\
4gM1BIWe\[B);RVA9X:EXY^F#=.SOQIgU2BLW:E).[<;-1@]#[5GHc-=70ITCV=P
d.X@A0Y(/^d4GZ?@?4[gTHR=OPgc</K/.2\_Vd@WKda4+VF4(,S0)bD0/\e6(W+_
@0#3Z,:[:G,HAMC28H[^H>O<VbLEfI;;G&I>3K^G(US<Ia.02d4b[@-5Z@:1H>,E
MW]1bOR1fAKdT1)N48QTbNF_LI^#He+41d)0C2_P:EAdN<\bCd52<4S/R-QaITEf
JSHa)Y(GI-W@4;24@#;7g-KRX02E_Q3Rb&<J5S\H=/0gYadFdA^Z.g;.I46c/X&.
NGE=ZTL#^YFN[9I?^YKP6\e0]S8D3[:SAg;/LIO\J-YG>([33-:0:DY\gcKJ20IP
4OScN7I\E&S#H7eIE<d,B=c_(^YT/O)K,;R@-6@7)][g4cD4;-Ed?^-LL=/8+4+.
<?,fU2AdMK;ILDH+6,Z9-:?3&RLO][ZUX3?S^e?b>TLJ5+(P2_f@T5gg=eUd0-/U
^C4g_/.AKQ6Y;7:gQ0R]BI5Rb\<^W)bU309+NRHV>9PQ52+WKcgZ&[g#\fDG311B
YISI:d0,RN&V-Xa0M,,PX.<IJZAN9<=4JFS\6[fXG5([3VX-d@SLb,P->07S^1JS
g?3_&B6#J/.U/.:LT<.>=)X-TWgLd>S,2T/5Hc;P[.^E]IIOb0.)\_Yc;A7/g/[P
a\V8/a2#NOK9;[T16K:P[ELH]&&KX=CYVPTNC>+3S8?,T+JBDS=Ga>FcW2eJ=aNV
L>[BG=FE;IDDc_/#ALb9X]^QaI)SKGG>COWJ_;ef<^QTZ1U+gfMF_Yc>.9TRC);)
TW:bFCHHVaY-KdZ]VaQHIU##Z?7AVJ8V9GWW0.C]6=Z^5K;0Ad>e#OG@WAM_.c(.
@JF_KXQ0X)Lc]1/HIE.7.)+7b&a\GbP^6?BSGKM^SdJ.+<Vf7N;?K0d=@+\8^(Y\
de3NI[[aGg;?UP^HE)Pb[,8,V>Ub/H#1@8RA/af,&MG9SQN=W?LH/QY&EX7FT&1>
eX8f0FZ=WdUXPgZ@8BB83dLK,E&#[QDT&?21ETFPOD^.^NSLCS7CD.HH#QW/@9;.
b?:FOGPLC>_]/586\,-FY7SU\9H>GNSN0L/#<W0F<G#]4@/DP2CN;@^_Y/;NHPHO
S.-GB:PbO@V.U)>,cF;8e?;_\MKXM1VB.3cH9fW-T.<GAO-?Ee7@-NCW4;&(]9?K
QWBXMY#U]TP/B@cdIX8OJEWD[VAX]J<Y@FRGPCLLOPgQ8J#3:1&BR([7?_IZ4B2D
gE7P0321:fI?6@V/#1>4@Ue<K&MW\OOF,Ob-Df7?1Qd7N>1PBg:04dF0.0WO([;T
P7/_;I9#=V&EeXH1X@Y:cMa]\)DOF+KBYSAN-I)AUL;g[QV^TN^=57YAcK2_&W#)
^F.FH,&8#ANQ13=#O?A,:DI)dK3W(M]N0&-::^R_G.F^73NQ:-A61D8[DA&:Qb_L
-ZUg>HF4?9J<Z?WO1&b)HFH@.bdfI90M.QMGH/Dd+)CXYPbP4PC(.L#+W^<NdaA2
)L\8geXb()bN)Fe.YC8B>7S]CcC-CQDdH]1+W+J)b3<PQ?+e@R=(a,=IWaI^NNe+
9f77a]S,G[IX#+g22VMPV2caB::39WU-9M88b#BQ]ZeTc7;CAH^;M[Jfe6-73F_1
PL4T9_L5Z]]-GYAL+52b1T>N_RY9[G8(/I@MN3SI0Lf&S);Wd6\-EV,WJ/01EYC=
4XG0YDdG];Yg?L:S>G0&,\aC/a,/S<Q>SU&5[,8dICXKbPe>_/H\DeAQG-MXRB<d
&J>M-Y,#;8Ce+TDdNC:CR2B^=M:^gQ.E<JJV(U?[CZQ>]^#]2XJR_(Z_HZZ#RTTH
,(<.=5<NeIME6V6EA3>g]7g6-J=]@EDFG>6\)F7#I>]Y\4BVI07ZX]>)#ZN/AHR[
T9N(?7G_?KK,NC=A?ND<0E1:I=S_WWOZ(G<&fF@7<3dCJcRW5Df[WJ_cI)=;;6Ca
OED.RURQ?c/6Pf+O?T]1.gL-D9KBBUBGgBRG0OPW^bcU=e4=<L.PE2+;/6K?&]WK
B?3DZU;E/SGKJEc[K;:YJ?<;+(U070)SRBf43Z=:1H80+KHUW-Nf+WE#?X20==T1
Ee5[/)H&>Z-8(Z-08gd+Oe>RCHgf<T=8P>B/\Y)O8LK6b1fBEfcOQ2/2X&eBa:^1
DJ4=;@Hc\>;KMRST)L#IM?BFae,]Y)\W=E0g(_J<@H,PKZ)F;D75R[I:bCB6NN,g
J<REQEA)b5#3e>Zd6(/\>-dc=J)22]bcG\>g)8BeZETF@B4O3=dO:..MH;,42V>/
X=I\W6Q;b2P:RgX\#[4;TH9NVYe2e,\f<0YQe<Na\A&)/TY7+?-P,R-B+ZB;.9XX
Oc]>&FPJ8<R1[:eG#S^X-4_MQVN-)6C>^U/YJ+]ff0:NN=NULZLT6\DBPa@HLA.Y
c/2c-9gd9:45E/UEAM_@(2AB&Gd^)M&@>&2>_=5@>g=Q\B)2E<PRRFCX.RXZ5<CZ
OD1f0DJ4UV2).Rd5DKX[Y1V;.XbcNF#T&;O=(A=8[LPASG9N4,UXU]XLDO/\+c\7
\HPdO(d+JQ]T4H7QfJ-WGHIf+cK<HZOb4@/HK2cKg;-TWT@W1P^bM7OdFG-bgV)-
MZ,FYd4\H4>=KJU&]@R;->E>5[a<U9VB@S4H>X>5C]2^U96N0BY](H;:6A?VVXK?
XY0H1cSgXK_L<EDf7A7&G/;..DJ5T59_aAe@?:/_gG0-)9U[<AGO4->4?F+7.HRM
8AYH<Y;+fff;WcGC216:QJJ+PR52LO,09XGX4eP-7<>U)MBD=gA;>#DB/a0Dd[C1
;c)^d;H1NI\QX<7J??2X0cMGAQYEZ@E:RWcZ)bE<cZZ)^OK6Y\dRb89d-TM()dMe
IN@=;-GRPF,,Va]E6^.B16dT\#a481I+=OCON:X^B5-<LKT64g54C,:9G&&eR1@d
&80JcaT<Y@:S#)H543K]B#Ng7.C0NJ5M)a_Pg9_;=<Z+T@5/V>@4BL6>V;5c1119
UP[<g30aH,gZ+PNb@46aP[WeN28)b65]>S7@@22a:9C+6YB?P9;gV<6JfaW+gK(N
^X;<#4S6BZdSNM6ZUK0,G15_(FZL3:#Od<9D4.OIJH06Q47#Q[&e?Pbe5;HO[PF&
d(@4LV+BK^L3G)6O2T?B9UAE6A3)]<D:3Y^,(ag?XN6#?1DFX181J37a3/PUN0AF
@+QN((9DgS_UI]_/]2X?6-c(B4EB7,Q_5C-&,0F:/f(-8=QN,c>JAMEG1J#GI=YP
b=<Y0AN5XTb[9H)IM-\dWJO^)GNU/UL[71,e8G6;1]N(<^I-?]71:EDcf.(@Y,SA
bV]Jb4;+\6T/-9^Xf1N4-Vb&YfWg6Z6G\>6G],eHORRL_GW(4(8Z+IX/W\#1V<:(
:I9S.+8KE]YeQD)7P^R&d\cD(HZOR.I7TI0Z>I=18L>WSQ_S99DSS:[9>:/OQGUK
S^N+)W?SQE@E7,b;c5VeXYWPA]<44A+B?K5;[3V9Gg?39Eg&)KRHSRQ]+.H1>:8)
[8c?+M(_@EVP]F+NFQa?dZTK89-ZV?gDaYV+,SfX3;3V8E)MAG.RL;#4XLND-XV_
(4HU]Kf-+P_Q+G=I<^Sc:9W+SYKD8GJWJ#;9U<QJ@JePHA5)[=G0f2WG/],7a_GS
^.0_>ePTBN5D/Y=dPNPH1K,ZZ)g?VQ2EO42[e@USP3GaRH0F9KK7,1g<T#4.5IG2
@W_W])#IZ:ADJRR8?/&)UJgbJ_73]&H>G2E.]XWHC<(H=7.G:@+M10&1.4&(/aEf
\WbP9a5IR=N#_/IJ6[N=.\X\c4BN4T+Tb]cX@b4f[;Y9L14;FQY<7U6.L_S>UXCe
M[6P).34-BK+>M-A;Q_/T9W]/+aeP(&@R3\:7ZN3M^JPC,8X6_S\ZRVY6-GUFF-J
_gPRgg^8R,9Pg59<EZL:S^-Y;KMB:G[H.@d@ULW/&dIPR<eL9H6D&HHXD<0;#1TW
]ZSP3._<UNH99V=\g_)L[E1N8)RIDMc.dED<BP2ZcQ^5S+&WA=K2OS<AGgCM\IAf
C>>&@DW^dfGI=4DE]gHI9-Wa3E@c+gbD-]GO0[X\0,)N4^,^K5Y7^7(7.>9G<,NA
(F96A1VB[++&+,ge/:IJX-IH9(IUbF7GS[.L?T3d3=NH6LK1)RR65^gaf=9d/VgE
3]4GW4e0-RP);UA>b)b,+f-2HCN[>-4Eb:9.B6aC0^/98VIAO<?HaOg\E259L[V+
;;2Y&5)0/(J:F&C34f^<MF._B??TINf41R@5ZHGD8.KVMM/-46KGVg3QE;:N,J03
deAIMMgec_a>,O((URINJ=C?3R:EIGQ[aBE/cfE]2R3F29H:&?DBSY=5G\G7B+5B
OPE_1,&0I&)8R4GBRG)-^95??2c+B(5)AVTZ@;384IJP2d4L6c-MaB;TXaeAV(U<
WF,a(W?-BRA)7W=7U3D9B[O425T4D/8+aMb1<F/<@(M(SN,F+;)X-,0\HNBQRJU^
KS\2<cM(aCGC+\450^Y9Ra/Z&&Z0X?E(8?M)f@bg;4^-?cWK0dRT\2E?L>06C#/B
-5&05Be)_K.HS-1@1H(e/=Q#[+HG=XP/ON/+R8IEefZR,+Q,74ACOUS]O=+S47/.
?8-GD9aWY&^IGf2P9+.S;fX7DXEeW@+TL^YST/EN#gcCVa9DWH4=L1&)2g<c/1&a
YUfbP,ReIGR;T8W81LQ(=LPHNC^96;3WdRG/IFVFc0cf@fF0/C2gK?_-RI/TJ9bP
NF<[Fd4:&J[TSXM+OYa4R>3P?];J-;YWdCL02EN&-6ZZ&B=2gMJ.I_J2IT<JD</U
aKR9;QaGf27W1(#<12cB8.B=0/B>B5:Q0@[]/E?QM]0dU6XLS/HP&UdT2cJ)SWB(
Cc6I:?J5^SdIe>;#a]?6bX<5.VgQe^Ce.WUcS5+J=gS#E3VYc8g_0,85R\]e:CWT
+UKKA)C?O#Je[L=?>CGDAIQ,6C+aOM^SY#Y/(APT.b2.?.SC8T:85G.ggM/RV<F:
AP?:18#Qe548TB\DWf[:A#6Kb-;+A[9IO3a>:78HB/)Z>_D56D],U;+U):L]G8,Y
U;CSCA_5+bT8><_:Y387@1I77]6J6+b@7F.-5M/gfJKB]1a,4D]IX(6C41/Z9?)d
&^CH&5R.BJNVW?[C57D/dc#SaY/)+-@NVCIY,A+PSdd/GI[I(CP>G-De(CH-\a6M
-S2??ZZ:>-Pc5L2H,57NJS]a19_<=;a0J7I;KPHH=,6bBcR2IRW_f7AB0OaSWXG-
_@BT[:8RTaXbG/A\<WCUDMW;-S:^;Qf<./3E=TN.K[Q7XK^.L=d0)4.fNa&C:eY#
_>YT<F4IN17=IeAC+4J3.[EW#IE):[\CU(Y\KG;[Ud7:G3d4OUE_S0D:48NR_=V>
Yb6fY1^b[FE6bM1[dF:]ISH3XCcU?V\WO]fZYRTGN9Z\+9b=BLKQFC(]>HZ\TDSO
0fMLd>19JJ9R:@ES1(EgYXePd?+Zcg^Lb0N?.,aPM<7[f\S19&LDHS#O<4)#^W#.
fGBAC>=S7RFZQ7DV?d&g^6eJHBG0\4a(2_0fGU&N1d)4AMN0baE6)U/MAgA5ZL8Z
=19VWYW[26JBeS//&[Q5[Xa\UM4U5\#.d15N7S5A80da@&[P4<RNb<aNAKKU4fW7
aaTH;4QYbQTOM+M?9P)4Y1;,R-bRaL(_KM/QAc1CeadHJ)BT[@V)01J1aK=TU+2?
>#3[DbW7-HWge@(9R8g^AfNVcE0cYJ?+;3)Md(=J))f@]0=)F\,[ee+OVED)O7DV
Z:PfV_=&<5:J6_;_>)9FQ=S4;/)/DZb6Rb]27]1a<&ABV#IGG0DH^G1.+S3Wc(K2
=\X-4@+EL^#baN9W(B1?(6T\ARaPM7Z_5c\7gH(ESV:0J.:1dI3c-@065YWU/YNN
Bfb7K;@Ed(^<NQ^6XdWf1U]HdN1M65(MdITHbE2Z[?1P3S4fP?c+@/YJ+;A8M1\5
.g5P;R/T@VPIMI64&TQKb/C)S8#;<=deJ7&fVY1,dSbfZF;d@:8[5HfJ,PF>[0J#
URdLJYG+97I;_6;:@QI7cM4>I3^OVW-<[FX,9UWX[2aNASLU0N54L#PVTMTX3HEX
DV]\&ZZDV.NZ<AN88)NNCIca\W6DP.O1;0CK,O:+84,_777dB&&b&f3+AC4O506L
(6)2eR75KCcI;L_&5&9&.?XMC)Z5;<;cIGX\0++VcLXOfWQQdd-4\9\2=XW-T/>1
89RIO#=[+f-J]U?(Q@7E=c=f-<W=PgSZUbEUJX^Nf=<NXX@::ZS(\808?Z10-Yd-
(Z^\_>HT;<B-#=dA)O1XPUWVaQWA,A?B&e)THH])8#Q0Q:Qb)&NG_K2652F<U7BO
8Q8K:,d\df&#=ZZA14+#8(M=(N.GMJ]OE6VIF5YMQCQM]XV33_Q:ESDQO:@4[X4J
If\;eE=R27;C35/.@WTg0YgWO@bD?>WULf14AIe:HZZQ\aL5YRCB1#QKZ/UOYC>\
+3DKF5E\PK9:10.2>P(@dG,fGc,)\=KE(H_1)K,I.U(HE8Q9(FG7YK]M4KKXg//g
=794-ag[\,R1F,>7Be-V:3)]\H?gE1RJF9UNC)U+Fa7S?6Fd;>>DE4,(Ac^EGeVf
@ZR5/3Ae_IFKF.IebB6d.=SMb/D;)\gQgLWZ0I.1\(R-3VL(7/]EL,g;0TEDM&)C
<[H\W;4f00&UQeV=IX:gP[YH4A[IFcF=8&(@?,+/8;Wc^Wf1+e/M@N0HR&\X]&6H
8WT)@T;D_IOOIEP]^O^=R^&=PVCDQa@Z=JRKJ@Z7[\<0)SH6^aZ3,E[&db(@>O=6
IU2H8>1:ATe-b[0L=N-=I,1)MUN8_KPDO)5H)T8:4G7,d-(Q,=g[g?bWICJQF\,=
0f?gI(Ug+6(2BQ<9@b-8E5<T_1K(e1C?[(@8639K=XWM6>CW,DcK_;4:8)E4/5_:
7D]Gg-<QcObHU8^1FIQG5Q,?FfME(;.-SGG_9gc9C=P;g<SS3?R07Id><\6Q(562
T^GC^(95;YJ#Y,V]5K+1]448@g\]U:G_gU@KTIHbEEaI>O[U^aRV[:M]ICX@I-<M
_25U&Q2P.FH9bBX7)Ye?3.J<8Q8KWM:Q+CWU50\Za8I2/#5)5>&5ZN.IDd8\3?c-
,1B9/@0bN(G+6aDH-]#IG]B]P]BK0;0Q5c;.CA5JZG8NM6K^XB(7+]gA=>=bVGB8
4<M(2ADS0BZHH/@)6M,<F0\P34GDCQ>dXX2;K8dL,1B=0dV.RMU\#UA)(Z80G:S2
KSW(-HeJPM4[;V#S9F]UCM-K0QKU8SZ&=[0:E1(F83]##M4,D5H0&Bg/FR4aPdQ@
M(g.H85=FP(:Z]gDa@RV498APA&Ze^UVHJKPEE@N/2M-FHA[11AL3YTYXCMQ4CGV
f=eS/SGT-&CcG@TII6b>CVOO(HW[+&Y#c#K:FfaQg-b;#JEYPGINBdV[W>f3JVDH
S:I@0.@>QC^>caa8B9ad:4XX)ZZCTY@#WP@5QFO,LD5geB@4cJ#6O/A)e:gCM.A&
.LG[@4&]O>A6O+/[8KDP#\c><6\f&f5a2&L&+aD\e9PT2AgG1^>7@PVQ1=,]F+@O
)5L3RL=-L9>DR7_dJ3)DV@;^MUY0dT_PIKPQ5,aL=#(TQ:Y]JeWIOO;-=:0IFdBF
HW4]F6E&P78:OVJX@G5SYD@8Z[MZcQ]<(GWFSZ\&MN4e;\b>X4/<][NEB7QfRF8_
\1:=FWK@ZTdNOF(VHE&2=1(2?S2ZDf66-N(NUDS@K:e7Rd4_-5O>XbUU.LDO\Z[7
]9e=X#F7[L8U^f0>RH>ee+dJbQ(6Hc85K(;AL^dA6ILK=eM.\DW&Y6Tg.0AXcWY1
D]@HXS\R2c7>)NNf?CZFCRdVIVUcFILXR]J]69ZI6Z.cU6O/a(f4Ta?25=LFYSIE
bQ0M-fdROR[9?@e[C([IgSQP\\3:J_&bAV136A/DaK0/YPJeH).8eLdV]THPNE3#
=Z@,+81e43d53TeN\&e@IHV=.[()LJBc(NX<PHOJUKD888=)]14RYDcV/;\EJCGH
V8=[0>WI\.U2R_DQGM3gI#c@_;f6O9KN2.2(+X&@4-?CdEe/GFedgc9E?X(/)+5f
K&<9Bd.TA5CAJM.7f-E<C7.X6&fM:4ZLG_@>]ED/1cTH#;6OSN&7]F]M4.R.4aZ6
:EUJH2K_WCEVOfNIHMgER0((,C^.7F&gRAR9bO-OeCHf3K<88U#T#(EQZ6WQQA>\
@fc+R753c^T1[GcG^D+;P_TJ_/N\TBO?cM)a+GB^J_98g0X&fOFOHMF8SGP7R[_X
WZ6gH\LVb?Gc,<B.ET?8.,^cYFDT8Z)HBE(O;F3Y/JNe2UXF8c.O\RCU_5;MI915
,Z>+3UdKGU].YRK-I6YUASI,@0?M\-.b_1SVe>.5)-QV[Bg9@0a=LMgc/E5KL__]
@_FS4ff,AF],V(O_Q4\C.A^LRMQ1E5,Nd:A)@8VB,cS2]aQ7+=LW=&5RW,B,2A&H
R]C#ccJ3?N.Q)Ec0#=05<?+PY5QdB<eb\7f0MO7]C-WNH.EP<=eTUS5BL7WBJNSg
;Ygda(9fP_[4(:6R6c@2VGZ]JHXDdE,-EQ=3.d?Z#c#5>,e1-:6=-XA?\7#4UU,#
/C+Z+[^\R#JePN-(TS_Z+B?Y\Cb_&8TCf[P99]UR6MKd>/SSf)F7V9\^N-C8^GO&
))@\3#cbJ),0Qc[^)]A1]5Uf93HX04]?\?=(I0TeB7,ce/f,95+-9,^8)d#<>TH6
)4a/49TLC8-dQ3<V5LQUE\EI:aY+B)CT>bS&g/C1IF>_/C-[cfI,=GT-Nb7S4\@K
?bW01S-Sc\SLVY>IdC)T-9b@;Sc>&99+OKT/4O[9g=K/9O,FVVf<-Q(65R5NRY-#
R4K,N.I&ggGN_+A=@)b4\Y[f<dKIccJ8B.#)N5+gLB0,@ENFNV)d+<0a6e:0GH#1
8Ha,4G_Ac5IIE-LUVK[O]Kaf8gbR]2(39==&#TKV)[MbZH0OS\P[Tb@C12S\@_.M
LdN,ZUc5Wc#VA6b..a62bYcd;,0e:fff6_FNHVae2/dSA(U4UJL501S^4:/<S,XI
#8]2,I@N@Tc0Z]WZ7G?R,V2d+VW#=E5TM[=_?^D.SN>Z>#1:cO]4_>(0:bA?f1&-
\1FNAQ=.-_;+bU=\\1KHIM).eF9dUF_KbP/-E]#0=GEF)S=#gUNW9Y^Y7-7\</GO
Dd1e)?VdXR3[P<K-)Cb/AM?=7.>Z-8@TeK7+))?MGdEJ(+aOUNW_;KCL)&R>=\M5
4B3Bg,V#W;?@:0\5Ne,PZ1N9W0?<G)MKfU]+P351?/2f(K[Cd6M=:WL3d]d/_(O:
FY40=[C&+F.\EQ::_\cO&M@BU^7H@d2bJ<;d36f2bL7Cgf2J,(_>E<A_;27eC.R@
+W1Pc#L=a<PP);)>A.Q7.4P.d8HHRTSFHd+5,0.-f+.,)WL^&>df?^/aZ?cI70a;
9FZ>M#?S#+/@-=GYgKV99RRIP0e9DKO:OQW2B^,B34(T1MMeEL2>#H+/;WEc4STY
1Q\cca.N2=Q)D@H3Z[&O90XEGb)/N,GA32/BOQa\1T\B24-SL84M8eYLdZ9S72<@
c<:&E>ZATL8(8LO&2_Ke5^]?FY,<JNH7<14dOA[(_LF9_XgC^XJ\ADG&XXb3\aV^
;5+&6E?.7=WU\?>6OgRBF,Mb0\;TN[4e8DJ_BYI]Jb9-71C&@:EGb2DVAK3c/M[H
.b&Nb.=BM[c[6[,PI_484)&D?R+_#4R42A[L/&H1eW0=MJ1.=?4BQgeg;c?=P?X3
Z.W4[\W?84.N3AdSZE1,e#C)G64\&^OO^SG)J6_bgC>4?L>#[M157)AB\;ZG.@Ca
cJT3WA+^e(]AR^5Pe54IT#:6M.(7UXfLAEU98UOW6CTb8Cd3FB2]R<-N[Z\^X\/3
+.gZ5RCBDLbdF+)(9LWK:9.bZ\e;MO:O:LI]CD-4a.Lf&_5fA^C1eAXD(?HYO072
WbgA7.=Z_(f]),/#J0-Ve;Cd[5g8Af+R,,D?be1?]G&?=FZFXgT31gDE@37SVVS_
FcJ@^8UFCBCeB?4VOC((gK(E3Z]e>_U#Y>_b56_GBS972d.\4aI]A,EW\.VK0PbO
g:CRc8IgURW#ICB+T3U8e,f4_fX==#Y&<,dWZ:WeU+XDa;Z8R^?+A)Y,NZ91c;N4
G]VTP(6ZZd_^J-1af&gQ]QOJ8<MGR3&NH@8+BW,4N+]=a,=FP[VNL9>VX)A.7#gD
PCJ>1?PT14aXSdZZgE33dN+3b[[C).7Q[=;Wc9D<>04[<M(^<)]A5;Bc;Y7e8);,
7^=d1S/K=/D;.1HK^+83A=<_(8=)3dN(/U.L1],(Jb7F=QWY6O40=M-PX8bAbF6I
GM4RQWT_?0#F&/(c\7]IR3YOY:U&SF1)[(fLWV[/Y93++>Q]JCDF#cFNIV4bK.),
]U5L)S)<OIc/B61/+TSEK6,L52UXC9B]&[P)5gFLc4[[]HOB3b=:+VDNE8>d2\8>
M=C7:d77N.\@bR/?)9:dI65gXE5Z2Q6UHbI:6(>_Y.3eHB21+O4GMc8N,9N0SD6K
E<D;eIEZC>=&c,\XKb(_5Bg0a7a5[9#:^(PgN4LS2FHBF^;3QUKNFZTK4>S28T<>
BYL=a?C05G#fe9LO,1@8T^1e\I[<:\<QC_[-@dSE?=,GQ)T?aOK(F?8YYO2<1?DV
efOBT>OdFY-VM9JCd+PU#(d4L7G,&a-@Id=+-)L=]A2DC)aH/aCT,+QD\C.SAe/?
eB\HgSWZR]&=VI<32:1-5cY;_1,f9VeXHP>Pf1_(g0GWA&7Jd7b(U]\g/NFcI8,A
D@DI^Od[WB>=d9ZBZ&^6G3T_PJ4<^^.3+8U9a?e0<O+>JP(dR8;HW?bAT+ACF74^
c&0HO.M\dc>b,U/55[8_,ALEeGK,I^1P.<=CMG5RNE;7+fZ1cU>&\Kg[=21)gW6@
+Z[Peb37^=&VPUcYN0a-AVf<@9685.Zc5N<#L0&68PCg0.[R(6^Q;,A?<,@.+6:C
gL)XU@WSRYB+)DW3N;UP>G5;D_91g7X4J@7-?:MRA?d#:SbN-F4=gW=X.Z3@U[3/
-SaKO24>Qge\YH4^dEe8)<<f@X(Tc:N8G8DDe#X8?8HRP418KWXZ[S.:[8PT_RD(
=(SQF@&3KaPXc;Uc2L7)B/Ga>VDD[@0I+g1@:R:RbFY>,>8P#UD<7&L-F_eIRD@O
Yd[a\I:1V/3.OGTLAXDgLQRdgML_R-BMX<B8:f88.@,__0NKf,72V7B7?D>;Re_=
R-S;+@]=L1)Sb>gJ<(OSQ5>YXH>@ZJ?4(e;H=B4J\\cZT/dL\,2gYCX?eYe&(2e:
ceFQ;dHGU6X:.H_9#P\#[dE)(HG<9[g/S&_W].=+:>/LZEH\^#PA.X#W,5@B+d14
\>aa2=aJ2Q<D(FQBPAeXFX[M.gK;_Uc/XQO7/SJ>X7Efb5C0>ABI@g+40Ge2,=>4
aSZV+5ONeAff>;ADE?a6Y^_Y+QYH,E)6c.RZJZGMD#_db>Z@?dCc<E^WE9/:CZ^F
O&RA-K5(GYLQXVLgLU:/,?Cgd/L;UDY,XZH(24>Q?4a\Q2YOdd:6-RA=T][GKZ-d
:K>58D[_K/4(f8NP7f8]/a?g;gO>LO51?Wf_-S[#4E+9EY\C,EI8a5LIL9E?AU,5
1g#9]>a=V>2BH51C>,9Y,5RO/))MR=1JAcbLX)CZB2I2d;JQS5+SL39DcY,HNcKX
>eATfZd3LSO5G=ZGRV7F4CG^B:4(0H]BKBL12LL>d2DN_6cfaA88Q=e1>&+c5#b@
43)3)W:f(Jc,ZcdIEf7M5FYUTWRFS_/_U[))0#>/dFcP+RU&,W=FNY&<>>0e@Y)H
W@J+Ke_#;&E+K)>&CU?Mc/Zf,>7)<\L,e5;PdM;K=+\?+I6<d8L2&b>d9F]C;C?g
302WL@Y&Nf8HZ\_c]2O6eCg:LR5.4<OEgQdGAI.BcJ)(KD(W_cOPY?]Q@F85//9e
4=,LW?.aXd;@fB4;^<b)A.@cF@95bDgHU]KH?IQ.TR5W.P0Hb>ReW)0C3B#35M_&
UXKN)0JE&(<].e&(MZQK(YgW2[Na(;QS.VY.Ab.6Ha&?W[:RG7ecc2J]H1:X=.[Z
^LJEL9R__g_:TOc.>7C);eM:(#f/7<KZ#;@HWV]TF73+U<[fag=/7ZeA+M;3dDP4
PGPBN&dPf09_e(H4_=Aef1A]:V,=&a<JcCgdQ9>N3&99:-<XNf0aK>173E,51(_)
>W[K_QH6;.]&4],8&WFD0#eE5Q.)gaZS1+Kg.LHF8]JdAf39\AYX)/JEa50<S=3V
Jee<T5>e0Y\P@XMGQA]8],9XY_418O3B0]Sf(9Je#@aYG7Nd1:\EB-.A8O]=\[]P
MLHb^FaG-I<.)G=MZ:]4U+a[PD2;_KgE[(UFa;E3;=@DVS:7_f92JbO=&YI<JJNA
+Z;ZVcbJNd+J^W1c3bFbZ6<TV(^[YZ?1g00[\Z;g;>5E^\<KRI02\-,:@C_5OAT.
<aPGX57LODc4XGX6Z_>(S>,7#SA_,ef=B_=Xe\<@W/=<3:VYQ[@N,I@.CXPED>6P
fRg9Q#U?RfgfZPg;:]P]KN<U>=gSF6=-=HcT[T<,Q3R4&_NYFHD\Y+IZ<5U#fHP?
/MS_>#3KE\?S=GOCbAEO^eUbG4F;:DDb706/&?\ec<Mf=,bPWf^=B@WAD=-6(8EI
a2..._cdGUV=7e8?-RW]CQW.2#30+2W^aeSC=N]M\7?C#^a\KU?Y34a]WSgf>[D.
.-NADf2.[#TcSD=XCLc6:<W.6)g#3Ab)5ZT200I^Y+:d_(9QM/,Wc2-.+&Z3=Y(P
9?7<>(3_W05^4F6@Z-?Q-@X8CbEN13(3NG43SeZN_31<,QGDIUUgILAJV[DJeVNM
fB(QBL[^2^W4eNKg=EeAPHgAd@JJ<bQ9X;eXEg>3K2;-e8b(aC>/FK/L+cWG@FaJ
^67gFDNQT^DcX:5L.GIKIQP#?:,T[]>@.5,cE0bDNXfE]@:Q?gT/S[A<JM):JUV1
&1)#(&@bY63=ZOEM^]PDU=6_QD=??#HfdZF#Cg8W27Q_C6acV?:YJEUD;)+]/MHc
BC;/VaS/#56-R+K\:/HW)ZD/QV3+F=#K+WA&&dGT=R#YA+Z0=aJY)X0bDbP)]9^R
bAgR<XT573.6UG57R02B@OJ@[40dJJI9T\=;D-@Ug-+c38L>PeNa?gOdEY/4ec2G
_fFZ&Oe9,RAZ2.]QS5fbL7=fgdDM2bY1M/7Hbf4O2eeRDE<GOP>ZUGP3bYHIQSER
f-MVIXIU,2K><e6HQKd6Y.0\a/49(AW#19cYO]Ba;V?3ge)^>1Z&5;@SRT2>\U&J
&URP//G]5c7@O_8Dg7c[e(AK<-,+M\?-aQcb&cgY5O2&c#>N^IddO@AICOb5W,8M
:N+Se=SX/]PQ=XDcM;+K^TTc+5UM].E.-@;,.aOcGI:EK7ea_\-S]c^OXH1T,4U&
2TQ\5934B-5<,6KC#ZG95BMXLMD38A(bG25]/T?Kc^L]44f#)KX?GLfI,Ic)XgNT
)0XUI;;dN591?6ROa)T8@GZL.L\TIIJD\J8bRK00J2/MS8ZdTKB4I)47-;=2Y3<b
3X>28ZF/3)]NF:fDZNbf(W&OELE3,F6M#(K/A_F@8,ZeO?\Xfb=M8_<aU]0ZYTg+
B,^4Se11gXKUgb8cQX8QA_@Q\43-CW06H320:M@HHW@3A0Y)P-0OCO3M]3/I_AJ@
gS3@VF\IV>-M[3>KXJc6]RS[cP8]L6.bO8dRSQUXV,Y;gRB\8/,/B6a;d(WEW.^J
1^&Xd3O19:I+P[X38<b:;E2LAD)T+MY[)OWFO1VBf(-WD==S,/f-R91e-\9ST=3>
W1(@A&FWU\UO>=UU[TCG.NBCa2MeG+I>bM3J=f3-@/;DC4Q[c&/(L,S;9g@/#5A.
?20<FbO^Oe/W^4+B1e+39QYAEVP<,e+VK/:a98,0==7P+\P\bF&MOAGOVaMQ8EYB
&UZYNK5df;f8;dD-HFC<La9AAPPcH.Y@W3e4c2C]49K.H0g^7QJcf@W,>b7W:XQH
;a:MGY.66\d\NB48]f,4T=c^WYZ[\6eQ1\T>UKS1e<IB7&e,DMfM#@GGLg?Pgf=N
]4Ed\GXG6:\AHS;T87d:U7&ReDf]6^JJG>3VQ?ONg02;(@),Z-,Tf#)6[#VeORO)
@#ZQDI9e)FH.d:<<1UNUYX-g(:gS0>HJ7CaJ1EL0H,:&7/e(RAd-Vd]NLWO)XK.<
Y)(A3Bf48VV3Z1/):97?TUg>:ZKAg42>FNgP]@<E-4VR=\F[.?W+VP<C6S@N.Y0C
LaI2&]Y_50D+,CP_2X5D6KT)R]e;,WNQWKH>P7J:E<7<C_\H8R/^6GTTaFY-X):P
S]IG&Y:W+W7BZ[I38>#HE.Q3:DU>V_5<]a:3\1AU:FfT1I_@JZHS<b0[:NXNZg4I
f3^N#[W,X+E<>ZP@W3_-5T[ceBb.#:0\gdF=4\KMgbW]TM&9M.I(6AF((@D^d:\0
=9P5-<MZ]OF?f;YH=#0B#<6GNV:]UOE0C\MV)M#_gYM#(dPeNQc&&&33JUcFL;0(
3-+:H-E-7UF>.W:D?L/6Eg(XN#M-IDS;_L=3f.R/I4OT868@/BUcDB&f(MXMOKd+
MNWJM_>U99KWVV;I[J[BRc/fZM^E=LaIJe>(XP9Zg++(2^]Q8+5dgf>LNNYId5fG
TD,#57;95PS5ETRY1G\3-R6Bb?6-:VBM1-W.]DFgITEQV.;1)c[G_(OKTP+3<?.]
Q.]2-g3JN]2bN^)XM]GBaV+;Rc44+9WCE58O=@P.1.b>XE7/T<CF<cMf)F>Q]3E1
18DU2(_[V(TNd-M):AE_4GDa?6aD8a\<CT@GN;P1g-CeK5,_3DAKYSZ-2\EJAS_3
b^2AH)8[F//]G,2f)T=B5>d-^:X3SE:)+-+V65b<@&/OYRZFc>b2^fF]eFO?/A8[
9YU_\:G_B)PG/?VXC\SF;95E.N7U)6:e0EV-X7/AR]aHE/X[V10)M6@?]099[HKO
+3ASG/(&3Xe.POD75b=T4&:[[FFGg?T].2g-KTfKKM/dY)6T]2Rf.W\42E&0L2La
=>/ERC=0TJJYCV=aE)UP<;He7gAO..<]8d@)4TKI8&f4=aFF:-P2/3D8Q?-4gVYD
M^=,AaCgV\LAcM9^2-GL]V7I[28:GD#L3TQ,>A>(Z:]/Q/P,A;SL^SCRG+0_21XY
/SggH4TI[<VIQ[EeR:1R=-5V27b8.^CG1A7g=R3HM\Q_0QA7Z,PDWM=YJHE80)]A
NN+1-e&2)b?QbR<SVPU6b5R,130&9\6A_a:.MG92Z#D1K_.V):N8=QPPD-#>8^.F
1NeSW1[12bW<Nc=+:AXd2FKc:?f>:5)ZI&_RKgSKA>G\3Pg>I-WWUe6D#7/g9<Y3
QA^AG?3.JVfVZ2/>15HB.AWeb0870KM5)+&e-)YS/AH)2_Q=Q_UOOf5BG=CT1/a3
#X)A@:.2J&9/dN<(XEK]K@4b;:1O6#\82a<U4Q1S-MC1L1MD11#OK1@XD[Bb,Q1O
g9=4[+SZN=b\(7\5?Q:g56[F:B-ef9NW_AS1#&I,Q=VV_Y<ZaR-R8;6Kg\f@RFZC
f.(2E4,g<TbYf,XDK[6^)2bRZ/PI_M=H8eJEF_KFN1V+81E@FgA)<NdO.Vc;Z+U(
X>A]E/XMX,RAL3#&-O(dD4T(G-WLCe9B3_LC/=I93>E?3[WB5[C_RNfW0FG)D6CI
TJ<PF6Gd>b-d.YKb&7\#.(QTOMLH/V-T;7OP+a\A5@7W)KM[C4_M/R?<OQ.I7\W:
;#F<?GKLZ)BWHRMce(QfJSTPI0fU-,X<KWO3dXV=?]=H.ge.NETJQ741\7@#d790
BdM^;GdKfASL8]E91S..c6\_NR\ac5?8)HKaC>]?fMd?S@W62JVJMSG:@b)R\fJ7
EJ-Ndf^PZgQ]_TbP6-4Sd[c)]g^JJ7HW?Z3(K+?DA^ceMbRc:4HZBI9B<MYN4&?W
JX;,^/2P/dF,YIa1FP<KdPg)QBYYUTNP@+gO5.4MTMXB@I8=eRIUN8R9>6eZ5P^B
#86A^I7^B\0+5<FHRQ/=X(LJE5WU;\\KA0LK48>V(M5>:^6Y8B\3OSY6B3=<FOZ,
^R2C1Le0E[O6]Jc]>,60<;D9C.I/G>TbCA,3I.?Te7A\eUAEOg4A<PW8H=>-YFQ5
W;9RR+9ad.\;NaH/QXD]2B(NM>3V^-2GNeW-IH@Z8g>\J#/7dU(#NBR(D22)+4=:
MZ.X(ND.]b[,(46>]+Ib<TZG#,,[O>66@V6(:5GK4f6b<Sc4U(,Pca]4(8A@FDQX
A\)Re]W4:@cDA1/D#)YF2)d:d^.ZH,XU,]fWZIC;K>b-F^c:>^O,19:X8PSQ>O30
8YCWW[a#PGegT7LEXSH&7d<gXLJI.8(;^_&N7?VJXOYaK07J[BU;_=^e-+L0AISa
I^8DLE@?MI5[:g>ASaLBY]VMV[37NK;IfO(Y7bW;\/3BB<L?V#:NC><13=A4[;WQ
2A)_DANeV;VE1(\3B8FT[a#,9&C0Z,HN]K)d3(0TZ<_LdeKGU9bUXQ;ZeAGbdb\/
F]5OJGY:)WOLN+N&7ad)XZ98/6P/O+dA:?FJ,N]6QbI]e5\N-KR^;-5C>H&2L.)1
DCS]298?3\[-7#2?b.fd9\1G<AT2ea9bZ.B_f+eN(PLAa758Y][39K@M8(<Q\V8b
^/3R#PJeYTTeL5M3(_88IV>[e,^YIL<UB7FF0^KT/_ME41b@(JWeg3R?\R8F;73N
VQ:M2[5OA</SQB,G:OZ++=)7V[AG3U:Z(ZE/9(BO7NfVU),GMBSSGWgL;=K#\FD;
VATN6ZV=D-<[XBF9_@EMP7R?eKAS-OEbXR+2,G-bH\YNcA@@Y^97W4?UA)Sb1;#_
1N[W#T)ZPdgM4#VE(GLVP(]Q@0L0X;8,Cg_F\(16<:_S+SDU+<RF)VUYAT,Eb1<a
A@ABa\+JTVYg3Z4e);b#/WT,H1Sf(17=b.KN=C-]PJ#eNeYb<3?Q/R/d9M;Z>D@O
[INL8(ZIQ6]?@2_SLMYXc7@Y&JY[fC#84g36-7&2#,,10[U3=(/?<5PbQJGMBZ_&
WH2\1>&&Q5T/N7R:)-bUM@(=;Q:b4#I[1JIBP-OEX#_>^_FE6#8.DH)K=V^A8VPP
^J<VTOPCK-V9LNKX_B+dI3B=\RVNNC\5OJR?Y//1EAVJ3e]PdM;=]\Tfb7?3cG^(
&&;VA1J^;ddE&bTM=WV-FN1XFNc7W2(;MQ>KgR;20K:D)]>L@52&[D>#D)++1Q5P
NF04Ya^G=@L16&2WBI_gccZQ00\]LL[aQUZ[L7B+X3MEFW8a7LAK&#W1@B_aXPB6
dH5Y7\?f1I?)E&O@OZYCE0-8-A6&6H_G@Q43R5P333?W0WdEY]c99QG9R^I\a,EU
CeBeC+MZVO)80Y?H,+bXA,2>-;c@WTA<IRWT4Q]NFHDKe#J#9ZfAcBON5/CGR/41
eM;c/D1UKB6CGH@4#SN2bGZ\B/_<MUG(_=fX\;TMZ,&\TW5eNUfG8MLVP[4.)I(/
P>VBON#8>Vc.gbTH=E<7d\W>3gVF7P(S<AJ=S)&d#&T/-I<3)S.ZH:1:3Y-()ccP
VQC=7GT4(X.^+3UOG)BJ2#c>AOCcMSSF@MS0ZDO8;d9)>+c1b9[B8ECJ(&OLOCW^
QOA<P.HJI)TM#;O9DNGf:L<F2=4YL9ec6+R?9N6>fd]?#T&1RMD,3[[aA#XVO?N+
/d0,9eW(_C>5e<Zc]<V15;T)KVfJZXaBN/26^8)B/J1>(GELZSNMW+LYX0#CH..5
7[CaQY;U,BRWRWUG]f.],c/]4PMBcG?YcIeQ.0/=-5>[D0/1a#g_La.T,9\&:K1L
0;,bX]D2UBBbU4\CM0RRZ#\-_SNe+80.D^D2cf8]P4IV.<>eC@b4K\?C0]DGBHLS
0Z-T(UL1,O]eIC#&;76^LRfI1AKbWF]C(^9>J7@>P4<dF+U&_aA0)@THd9?W1[P+
ETA:XW#c,>Ic\T<X7d4C_=R.)8;(8JK(7HESC?K?W6LLU3/OR^7SO+E__^AW6T9O
Rc&\;R>0K7P2W88:@/\7HJE@27#N5;I/0;ReE@W=6JNbb_:HIX5#4dPQ_KNWI)^T
E5-J/USY7X395QZ/XU^0C-@P\6JA\g;FXbaQ3GS5<P<9gPYYbD/FZ7]U^52[CgS#
WOc/=J2HETIeC9>-B[HWbZgB;2/\C5&(e683UL],e_G6_3b:1F8S(KO?\L,a=^TS
Og<JE0F>H3_ZW:OKJ?V:WeM@&84L#)6)I>GQYH-D.CfGDRJTL9/,C_S?Y)Ub(SE2
SZ1IeE.#[;#1TR3__D@bfN<@LOQ1ffN_J/0Q&?-A1GBQ96[0\MBNc(L^Z#ORf/QZ
GgafCE9[d>7NIG3NZJ\D)f,T+aM#ZM\dFA.<L=.<+UL]W:&&D2]0J7aA.<aYJH:1
H,eT4\G]QNQF#0I6e.ged[Zg<D\>1Rg#91JL79=J4]@FL2]RF^@G<eNK?6^),5X8
E,&CW4S)V^VR.HgTVcMaY]g#PQ&Xg^?.UFVd&UYCeFbKK@&(/H/=,J+b-cKCNC/1
P_T;Z;JXG10ITV).,5fZ-B579.T52V7XOP3B-^(0]52W;Vg/;a(A:@;W_=]EQb6J
Xf[_c6R?2XN(1R;^7=75(302,W++V(e42NAP8eM[eMM&DWJB&G4/7cAI&=^KW+eg
G6\CW\S6L+5C]_IfXD3AZ26&0?G?44gYdR&N)4P<:@#H5dN/@^b;gF^E^0fJ)VSX
@)e;Q_b^e@eZ9422]cR]fDM]R#34>AcZ+ILb+-J=5=bQXL:RgRR7FB1:+18QUI[Q
aF91[63]OBT]7@9V(C\-1Y7X:^EE4)[&/1@@b1OAKUIHD^RRCW3ecH=X[4d7:=MZ
]Z.a0+Q><GX7/1TYHX\(JB\J/H+1+[FDAR:;cFYRW@K8T?aIFdBfPH6UGKQ(KEDH
O.;QP=_9eD<NX/cY@+R^886\SV\C[(1H:@cRd(aTOYVQ.U_^+e>SKRJ4WIT\X_]R
O9]-81f/=1JZ6,T5[)FA0f]N5^a9V]C]91DC_M8RKb2MAaAD8KPP1PDad<gDNbDf
OIGN8<22U?O@8\e3W.85T86(TDcQBE]F1_X8fTEc24;g42CF##@/QD6<-gXg&UFg
+]L1<g\R#ccY2Qf^,QB;@QH,W\Qg<TF\Y@C]F,e@8513OZAPE@_?->FXX:JW\0IK
B1f4.Id5b@I-@;Q[]UE>=807\/CA(bV&]:8/KgI1UI.53=af2WPWE2#B\SeeS8Mf
LBJQS8U4d-fTU.?KUHE<b/e^Gc;G3R4DOAU)d-d#5e6PIVJO)YR3[c/?7P>aeX\J
3R8\R\W-PE#/28/9G#)H(>HOgBPgfUQM[cDd1fUHZE,=]L2HK.)>Nb/:WBGSO.<>
B.,VS2=gg1HbAT\SbV&\^R([5b5,Qc8Sb^TAP8RNW]J;<?e)OZPR5MPX78X?fO\=
>,Yd(#XGg&Y;cTA@WIc82L3gY<L/3;^a._E?88=-EBK19=8,FZ[3I#aCG1FV4+g9
R</G6GHTA5IdeJ@HX.+ZFb-#+I=ZA8PRJ-=WFV(;VUJb=VXIKdL4WE@D+R=H(b\S
fQLXdA(]0QK?cDE_c)aB?#+.&9X7QU+Qg:C9^DK(0.W_J2Y5dQ_TC):CQSI([FHW
1)1-,5AJ:5aC-F^.L47Wf]+02XYe6X0_0a0KN4c>QRIW;?f5?\\b5cT:2f#3:[#6
-b1-.<RAPf\6??ag-b0.egP0#&bc=7G,VR@aW2:2M^eNF3=Q9=#W85Y8,F.bbKAH
5NN,/.Ng@E9C<Y_Z/WV26-==:d+(&VDS9B.ORAF6B7^K\N6;CIWW\(Pb?g3-;IZ8
\WNb+O46&?Y+KY@JI70BS090\]U1^]^bg+9LV2=J7A9B@+&R9TGG.F>\EOX/TfM0
;]=#9JYA_T7]4gH)Xg-5NF0&9OF5:4>.ZYfHHY<=;=TP1e9AYXG73e+CgaA[^Dc8
K+?VfT:]e[&LNZO\(4WVN@ZQGC>YZbFG=-8:OSER&#F,I68VQA-,:-ZF\6eZH533
KQX:\I\+080MI\fUXF+RXW.P,VI;58eG-D9;VD_H)ERb)EF/P8b4@(2:]H,JggMH
+>MGa/Y&M1N/QMN;c>ZBMe^0E>ES@OVE\g;1P2K>CN.b5+Ub[GHY-&MWQ+,7;V)^
^JTdfE-_E98aT_Y5(;;UWfTU[JYYCcV,K2Fe\HbZ7aDA?HLJKGDYQA/ab,GB6K<]
[(LN+YO\3gIL+\g]W3C09>d@;f?LZ[-R6N35PB@aT09D]F)1TLOXONZeS(fPIcTJ
b_NA^J,TPZP>7SJJ1I2G182.3A.F/N;]SI.@e;dZO]c.W+34A+NDSH3P;1J0_3@T
/ZgK^KYZ#PgZR&SZgeeB[FU^O/d.E81)Ned;[82]7WJ4XMF[bK7607,fI5.\39R_
?gTT_8G<\,eYB1f?X^40@O#FHf_f[2d_P;\?5WRWXdN&-FS(X??A1B+U/--#4+8O
J8U7/8C6aRIQ?YY3SBGUeK]?Q(:&g0bb&;,5\5V.IWP,1g[+[AQKRKW?<P:VdMX(
MbfU]2ZQ)[--#D8)aQB;VP>QXR<A#T+>NDeBLe;1E;ZeR/dXKT=;8+g)4C@DZZE@
JW60G;25f^c:=.QW0/N#Ke5UMeR:[4>ILASPE]2ed&AQY&:RA@M-b9U0F.)0=A[:
;?4+c+aOgU=ef9:05b)D/D/0IE/XfSZGc4+NBV1D.#XN(^V,1:Y2-Z,AZ/DHBQ(_
d\4J_\F,bHa+CM-a(KP7+\_S(_cX_P+W(cFTIcM4d)WfUc32?YYW62<bN6)MO9IS
^Ya6D9dBP^CL7MGZ/R^0:YJIa)1VK,ddI6[),B64AE2YZN^cGcW3O>Z_6YZ>U?8N
3&ZW@VVMa]KNM&>TFTGAA,(-9HF=/T;#[8L7cK3KM<0@LFfcd15JBf(6.,0+<>IX
J0/D?>H-1EZ8bNGW73-?J1E-6,+#V#I(NSeMC(8@-LQT,+-9<JAY6=I(WL]egOSE
SIIR54G=:KQQa7?b.]\T#TS9dgA3Q_4@FHGM\A&^bFS29-7&8F#b,1],\@))-F/A
ND1SSNIK#;W0+^BG#/WNR45;EBfGSd(<d7,2JEVPQB-faP\HD(HL#?OW&>VJV?4#
)b.?HSS_:4.J]1-7F:]PD^:^/XMKg6T1S#Kc<UJ5V=L@5bXdIQPDB^>/R:-UJgTH
PO#4HR-JL.@[b>=9:?cY2Aa?]^3^008,5))BG^Mc8R9);FVHR4VC3,TUU?<,Q-Y3
LceIWe1T];C(Mb<Y)8C^(0/Q7DU7?PI\.^:65J8a;aRgGSC4^BN)VF@b0J(6aFZS
_bYY>Fa7/\67^/d.,;\5NI&SXcN0>1S@7<>dVF9dQBXeEN=IFZ0:ggOGZ[bM:&IK
[VK20>HT,0SJWDB8]ZK<QbD::T80aS2VYIU/3a]9..?+CL=/_N3bMWHcL^2c53VG
XB([7_a=MUCY\(F@fMBTA@1.DaFCKSa@+LU<5FZ?c;M+,&>(Q_6JKC=;<9]4cTbV
8+^If9JX_Y_#M)]&]AV&HCc=+&@XgZ328W0M6XfKO;3T/MUHIdZUd-9@&UL17>#Q
&?5QbC[3IGTTQN^+)fX]:,K<f@0&T),.ea2F6O98cZf+<QM[:VKPL)@WXFQDU:5g
C#\J:2_/S;dVGN6M;2@VZ,:FLWg5L7de?E(E+[;Udbc76g=(MfL3-<Z,,:-P0E=5
bBBG4SJ4326G<IO4LA,5@+FK3Z+1f^OJOg61(4/J5/A(5D0-X8HJ&(5DYM80-8A<
@TQMf.9T]9aQ=37eIZ#JbL^4aECaT<HeK;:2b0>/#,B<dZ.b]CO<.C1[T?EVA4FO
6QgZ)MY)BQSB;DU#M6]S<8IX:WQTPR\TKa_ITU\3?+PZ_:a<H/2=dc#BUVc>/FA5
<8WK)MJHC-U<(<+Q37VD4;=4HO]@-YfK<RA(Lg^ZaC<E&]DL<LF?I7)FNa\4_PVE
)QdQ\>F0TRMZ8(N2#)W:f5-C;?/;XEZ8H,g6>;;RR,K8WAb>/^O\85Pe-A)@N5OR
TV8V@DX3+D&0VEH[WQ/gGaKUFY]]61+&RVLaef8&2597e5;H<]cEOMQQEHd-I/G#
SKE5RK[1AJA_(fN)I6a&E-0L(W.M0CG^C+;^bW;W;3aWPY:UIGM5(6cP.U?IUTQD
6[+^/>J8G4PN,7-eU;-dHcGK17H&?L)Y)/MI9[DY#MR<L)B]:cA9\<7&F&-C(a?3
aKN5RaTdW=UNb[/&XXD++^T+^<dWe==VWdYM_N.I0d2^:=:e##0WeUN?25V)19CA
5KSE]SR@UN8SH>9ZP,0\MP)^:2=/H&4A)Xd-=T8(c@Ff&E^>S[MJX9&(aSMTRE#X
^8D7#U^b1;6>DbdU\#cE0A?HOS&V=V^O]-N[?L@P7/2_>UH@7#?3.d3QdZcQ_T;2
=.cb0[_\H<DMa.agcI:REO<(02P.1WZO/AJ9K7G/^)M/?SHQ5]eT2RHBc8/bM2dJ
QgME;E1PW.&4a>8(RQU?U<ZgaQZd69].)>D=A4N.c8.3A6H-:A/_ABQ.&Z9_2#RN
N]&^>&MZT,B;Y[HU=L9=A4TT.Sc^MM5fT5:+E&_=?M]Hd0K^2V8OC^&4-6\KG\JX
BS.FV]WLb7YfVT=\/f&C;X5,-[M^e/C/@/,VJ>U=L[#HFR@).[cG&QN\VO+TV1Md
bQ,g4_+FXD?H(+9;_E&DS2Q6V5A&VGa@E&,/8OK]I0G7N-463L?P5\E78IRQC</I
Z:g4X#9._UbM<E<G4E7QE_FS0b^g21Y];V>C9/+^0c(Z?I+-1dI=d2][70AAVLAN
+_3c[AWD_A6[39-0-9<WbXV7/35Mea=7/=_8[c&f]4Y=R(\[<WHK):GHTQI98R+K
dg-0XV(V/DA/1US7C8@bX..#5S[5F-?;(/bS6\PGC0S)Ud=Q4NQGI#\LK)6,I&\7
\(eN&N8<.aNQ@,.Tg^E):SQ])>IK+OHLTAR/>U@C]L2#Wg)RcQWH_8LI2JJB9ESJ
Y\fcGgCQ+S3:IUAdWIDGTg+X1M=L&^KL>J9<BX&PQZ6Qd-D^#L?VA4Q=7\X\<Kb2
A@ada832YPe3>):9J2[Gb2(0,JDM6_E)S@(7+^A(-_J@;Pgb3DUaY(5JC\+MZ=YR
SRDUIF:ILee4;?+Z4R280SI,I8G[d<(4[V1ZB]-dVS]A9&YL^P__9:O[3\X=T-#4
(.aI2T?bE0B/)FR8H]5]<;.QXZb6-)<WI+M\JHSGU9;(>F=HZPdc[V,(K_:;R\,-
YNJI,1UVX6#BU&c\f909KP(Z.+H8@J#15L(LSU77CY7]XOV3CDN8J/)IDc0CX2=f
b#V?H1>Dg]ZQDaS)SE]H57fC/W..NL@24@G>G&fW>H;KfZ8VEeDKL6K,eI04M^M/
:SfP>HZL7PO-Kd)IcBX;(^Z5A?A#4TUPN+6WL).Ke9Y\BQ>-R(8eM)0?bcN9:FDC
aJTJ]7F)JNA2dEaRF&+675Ke+I,(=V9@H8f(.&2WOR1eAOT/.T8H.XS?[FSfKSF#
_?a)3I3>>9GAceS/Me:M/W<O3Y1Z@?a3R^I,DD2:V:=8:.bS&K2ZH^^09@PCBEHJ
7GA\bHWeFd?/eG9ESG]AZN=])6_1G+dT23Paa<NKceU_XENHY3(#E+R5b1(U(/S)
&MM&QYT@[0;&D;\#)J:;<QdC6DCQZg@?NZbY^_HD^]0_6IdR\LW?SFEUGMd&_Abb
>_&B48)2J8Jd-47GCAP>aCY6_Y[L[VQ3aO+7.^Ub6gJ3e2;G?H[\<WCZD^?&08;:
eS8XQ>5S8[]cG@aA9W5.6U]IQYd1ZG8e&3^[25\T07]c0NOP,07/[CM9[aS9JBM^
18b_4A(I7K6;XL?U,;\aR=VMdKE@,=fLc_-D3(IIf>B1/?.dLaFMD6P?(:5FEb(V
RK)VQ(JA+S=\3Z&9Cb->FUMVAa;-Q;>-H>^2)4dVS[D4YKTKKcM<\;I_A?G<>3VC
RXSN&Q(?7Va>L37234=),2WVaI\aB@&F7J1V=DHbS7IE#9Y7^#9TYFR>H^[BgNN-
]P\H)WJL+G6T@&[aSWO[L==.L/<-@GI1I<a+IbGQ4XK,5&BMF72JbN;Cfd(QgCe_
97U)aLIV(U+Ga5LdMM[S-U3Ia#e1Q2+FaQ>cU00&8VI+/(V5W&4eeXU[LLe?)).f
S6Cb39(_V+Y=HO9)OWgb<UI=Xc7EdUP=L4aF?E[X,f,4bg;V_+KETSdOF+0.C-^H
EKd+DIMDA@76SPMF16:C<eR\Nb:YKU+8B5>Ia]OW?OUS^:@9-=_d4-WfPSO3.\R=
.F^OLZH9;+BWF@b/VX7>5D\GHL1.&6M&[2VW_MKZLKK)K/0,1]_/d7GH2^.MN0@?
RBS/RD6=&:X5/JGaRZ69Db[6+]72B.f\QA:R-<\51Ab7[;D^a?,aMHQ:\g+6,Kd2
4fE\HR5WOZ2.7(aG(@IEBY7XcS.9&?17[Yg]MHXD&)PTKB.;\VaGI4[8O3CK&fS(
G#RU-Y10XK[XfYISMe@1]WcaTE-Ba/HAVLM(ceOaLP]E-c0POI4T)T>\Y0#A@@_<
XAeSVJA?\U(-LJd,^C9\NJbHQ(a&IJQ.==HP^BQ0QVSV>-.WWL2Ad.LWTTDc>OO&
6Xa4<YR<9;TRSC:E,Z3A-I/QU9cI^)BHGC=T9JOV?7Fd<,Ig2)QTU>)_B>;[#/6.
62O\;O8.J<4:).#BPH3B4T.QYKe(RgP++JC.H03T2V2LIA?K?&/>4f0EfV:0^1Xc
)QXV;FYLB&bY/HTRdf_<1f(4EOgfT]NPU#++G/(K681?,1PY[&AT_L-MO[]M?KD7
8.[+P.]cP1#6>NR^EQG]3_0AOYTQ(O_.gCI(;4>^Re]O48III]5;A;OO>:TND@9Z
b_#TV[/JIX7?8IB,@)WCe7,4@2^.MHd=R/F>.a+e5KId&@<4XWV&ac4TIR,deOe7
Xa]=c8_g:YPaLfPg+<UW:A]OXYEYY)#,?B;3_)X0[^)UJ7.2[^ZUa.GL:GVAOF6S
&6D.OS\@]BJFN#O5=N9RJP6IFY:=OMgEK;_LZ[>RMV.X^334A4Y6-D(HH;,NT8HN
&-gc>(\g+b_EBc\8HV3T52ETZaI<(JKZdT<3)eJX=HFG_Pa1;=A@7K/(9-)G+CR4
4\H..dZNK@FaGZ8Ge4RBIQ5P-EC<D2A+16<GfQ[UMC1baB2R,>W?AKQ]/7#?<Y-H
4RD[H->)f-D<]2Y/b[5N=RH[J^P<8=/@@c(IFH^U3a2F5a(SGc=DgB5RTGI4_ON\
DU,NfEY+4I&G(YT+1M+8N<1b\?MTT]A[3ICb#316&WS/A]1F?[MM?EDNC:/\g=Be
9()</8_=PS/_\/Wd,Rb:?3B[g5@M)]--QLX&E&S60=gOEAgP7@&?-SWWOb#Sa-6/
R(#DU#KX2]U>#R\bR6/0_];8R-#L-=7a&:.A<KQ.1bA_#dAC)&C,1O>-L430B,VY
@4B0/#B41./L<gJ-U1MS=,8^TIM#G/HX4T/6V0PJJ>1P6OP?,+D1JN#2Lb;P>EPO
O8TUN;12fCCg7Q,1QJKMA2EU2RGfFFCQ<J0Bg.MG;:@1ISF=>89\^UbME2OP/d@(
4@JPJ86AGJ70fYM4BY@J_]gG_Lc#f_:cG#+<6eBKJ_#EYK\5eT1VWN;_bKRD;8:&
_D2[FLZ(_J&\,DGX<H/F0Vg3<T@I)bILL/adG0_ZCf#_[6;<9g8N=4MJT&>H:7ag
^U7e6+1C++f_]L;f7O?f+90-F3Ca9Y=Ib4TWQ9D.a]4:OGR+f5ODC,J37-6G89eI
>PG;[M=3+]TC2\DOTd,VG]+3C5gHAN?]A72LBKMLX:aBJd<>\6[3@B>(bLc339GO
&][),_6XYE)Y9[YUa&LCF\T,U4bbT5Be8Y<a#M+QgYK9>=&7VXXKRIIFgT]VX(G3
W#Ug]WgL02JSce5Y1/cSXgfE:?B=H#GCRCEV-fXfHf4?25Z@aN/<DZ&XO5+DggFC
(@3M/UfYL6ZN;<4W?QHP:>NTK\X,ZY4/RaaST^Q^UX-@KZ(gZ;/W:Z73YBC=ZLH+
X8ZAHf1.AT8/7]A5:6<Sa@LS40TH20c503ef(HfL)d2]6EZN_DEK:RIE<WDBaK11
bf+3dJL-X)(3FC)dGCBJ_-(FddMA;I@3:-MZbS8AIa5LVegYT#LLT3CTS7TGEM6D
.8WUI?C#gf(CN3B3-+5?(gT]Z[H7gN7\TdY(010SF-X(N5bI_9H2ee;JP;RW+/D4
LP98G>\DNC6DgW,V95fMCDDd<=/>RNH_D=8.1#8>9>E_@WOU1>USUbO2XVP?BM.X
?CTJZVWIR[G7(<BTdeP_GC[R&a3aT<1-I@Xc;ASbd@C4F0[8_+b>PD?+LO7R[0IV
7Hed7[C_,AcNBP^^/>0KMVS[.102A5]DS.0>,>CCWYH:AbSdWWVIE\AUASXG65&6
BKI()E@.3T-LH1#JW4W7-A/^MF6>73HBCES1\;eJ,NdOf?]T4(BW;_[_(-eOZ/@J
+AgBU)MR8.>)L\/SI6.FX,-=NdMcg^=00PI_L1\\<+UV2PM@c_[RJ?.]SL3fF@.8
7;2(U>^dQG1=L3OXNG??9=SR.P_R_8OC368cB8_dX+08aT8;HVC<)B4D??d_)]P+
M0(P\&WH+97MH,bET0V9-^X?Rf9@eceI=_O7aP6ff;?VY@5F>8dcM99JTOLaP@,\
^HJ<R/&?H6,79_&6:\:GPL^KW_,;^]I&\G_12HHLcCK<aW#HCeTX?ac_7\3I3F>>
17BW__SMcW@]B0,S:TM3EbH.+@Mdb/_L38,TaD18M:]U3/dYOeU+NKU<7>3Sb_7-
&91cZD8LZB=(&9DNOGY_bIK,P[:)Ke\OSg0=E:;Pb2PbgfO]:^T6b76-@Sa=UESW
M>FIBY.K86L7&W#AGfUdDXE_#G7#R[7/\,dE>TgFIAc3A5[AT+NJ_0:8?KA35e77
V?J,YXZ-F[1L[]@J,(@QL4f+HPCP252a4@2F@bg5c-aDD5^TAgJ&Re+R\b(CZ)E-
JEY;)8Kc))O]C8UB)V\fa.1I5?QdJ:b[4T\BA?#\H-dX).41A?C_+IT:CFDaT_gc
LV/GcV>(W=H9NR/.H=9e(cW0EH7:?3P:0b</Y+U?A2V)JL@<R-\HEI7FIX6BS8+P
GY8/;+W4;EE)+e#B9<?Y5=5,\@AWW,<N<^-2<=;HZQNf849[T4+>2WBOXRKQaG4T
@<W&,+a<(Z3aJ2K@L(J,,XOe5^A#LSf+H:C&=.K^]+UF#LPJeJ:We&2(AOLg^NVM
>+.Cf(U:10R[:<Fc4[<&:5c+>I5ZCS+5G.DOD:G75X\U#]&6)7eZ,6&\HT17G5(Q
OMZ9EEXcYI[CA#(K\ZefMgN;^[gFK/TIL<Lc#.)SNE(]Q0;B3_(5R6-NQXQ;gg/B
a<&:WYO\&LZY_6YWI8H(JT791]=&DV/9-.5(;74cXcFE>DRJ./BbKf1Y&(<Te2I&
G([N&LgF=&=WOg(T41JGa,I\Le3PU>Q1M^00:c7>&^V7F^BB^Ee7bbOK\9D039UC
a,(.bN/^;\ZGAH;,VUS6ZW72D2>Ab[NM4\A&YQ^UI^b<@Z_,\3:8H=H3b]2013a0
;ET@O0<-2SUc32V#XV7?1L/AaD1A6IR+2_fL9B,7R1WA+TAVb+8]3C)-7?,Xf4M5
RR@PG-cB+@3AC<&g-+&G;^TTbW\IB<+_27#/5;ZU?/2FW=8LO;dHSMIX,OXM<d_L
MPQV4A>HSHM\#ML\:GBee<g#>IQ6f7O)RE?4cXC\C.7.E_;a,D2D7RCN+(08SdO9
f5-T=IeZY/::^,&dN//64QUUH7,SE999CNS_I:)X5FXW)J9B/07I<J.[3W>#=C<c
AD5eRdB1S0=)1_GB[Jc+;c36,RQL^^UNG+/^WHOQ@\DAB\E0,c0bLe@a7>[81JD_
;3\cRcL61J3SYP\T8+#Q&.5WYTQeT#05B,325<I9&\@d,D:S:0ADf@)&[V.Q.+J>
94:?E1T5]51JEE.bJ(26,3GGbPH^R&1CO43KSGcNYdAS26WTH3.>7A-7Zd1CN,=U
GL8:;T9C@>d_<.CZ^/<<#^Z?\5#Dd_3Z(S_&UT(MG8/D85eG(ICJ0GJ33gAG)b>7
f64ReJP.a5Qe1^T)/G?82c]NCXN4)e3fH_U4W<@X(]NcI6Ffc.JNbR>K88>?@[H:
1fV6/a),gV33Cf,dF@A_g.L27)XLg@>#N7gEFeE8_:6&+?f?fRTb\A<7fLG4:Za.
I?KfLW<=dDT52W(XO]&CWN;<Y.27P[W),3J#ceTGbYT]#QR25E7,])MD)#A#]R_D
\e)O+9EX60,dN<#4:9YBF_)2RR,A_g+^:.BC31SeJ^[I@.&:L/BMe+UB_FgT=PIY
&@6.V<<QXX][f4BIZN_Q&U4EUPbTg>XdI_QIP8.?W#K^9I4gOJ1DaJJZ=&g=?dcA
.?Oe6B@)LVf)_5(1UB@Z+dZP5Fc:1I5#,NP]6(=EG:g0-DY-<;3cFXTWX8cfRO3&
\GZT9ZXRU[UF.F=\DEF^Y/3=f)QT=@ITFg.bY=6_dC[^Mb?\c90Ha=U()fA2]JN4
72(7:?)eY88U@E;,DgfA36d2A\cgeWT&H:2_/AM1BdU0N(KRD,,3+WQabb^2U3ZM
98e>f9(WC\X=8BYf/)5d\:.-][9gdUe)B[H#aeSa7Pa&.:H]gZfgP3&Z/dI3a_-8
-g2Ig7ZC(DA[P#JVB6/-1d]8SUQ#&7EW>-&Nb9&a[+b2N=Ge7;(\:9G0Z?PE)18D
gHL27M:Nb)_0FWTH9FGM@?_25LY/,KQ5F6##;LLLAS20,43@7R-MC1YTCGfI:e&R
7G#[?=UeSRLO(G9;[->[UEdgRc.cT]G7;7HfI[<N-T^/Bb6N4ZdDY@DbPR.NON[Y
A=D\0(3RTQI;P1X-@O=3e&?::6.0C@YL[ba64P-/IJBN[TLQ8JW?A9da0-9YSYPN
>_a_90g:VGNFS[adF]_<+^D:5MG#/V61[NP)d29]298HG\-b.FHebYN,L9-RR\I+
8SP9Q@?.AOg7@4;[C]FPTc@9#&)-4RVMUfC,2O[PfR0bB>Sg)_Q77)EEcSJ.MQN>
VR6/TfP]ZIA/Y78Pb#GIEBaO:ALGX(/V&d+=JM]W_He(V.G>0S+.@?/^8a6ROKM3
?M@3Tf.(H851YC>7OANV-S/M<<;O3\E-55#ZA<N_\Ed<_V<3dX?L\A[[SacP&#Ng
8Q/40+8E;3CJ8:?MXB(9P/>bE>L=IZZ/PZNH^LYaYXaSbGb;88>?1b_=#BW,N,N5
KOUNDfWFb3.3][PGT@M((-_Q\bF?^XDXgJK1egJ(E@8+]g8^?,ESYCNC5.D/^UbT
XgZN9C2FYKedBGX)G98XMK<=##U)M-AbJ]I=,U=BE0TRS=g.+AR,c7^C3W=\Od6X
D[a3HEF.@?,c7.K,ROZTI8^Q+V=4HHB?.<I:)63[eP950.1+4&e1<>Vb9VGD86AB
c5\WI<d>+K,I(H;SSA/,G@IX+:e]L:JTQ0dJ0E(-d-]B:MfQ[5Ce]g)O,=G0S-7:
K4+W?<U7Ob&>4;]#A+C?JS;c6D@dGDAOa,[Sg<dZJ1f3WYQ3M31B.Z,]9M5L)G)(
5T3ZD<>\-JC9gCW:d5U7Zb]X@-#72[JTO,:UF@IMX_#US8HeX#f7]:,TE<>([RgM
DP&?>3\Y\\HDCg1]46USX=f,X)I0I)XU:g\5bY/,F?Zb_G[3>,2GB\g6M,eUT,+.
4RPZddd;LI8=LM./P))ZGBWUH/<-B;A5IFXZ0Nd0/HbUHZU,KR2-LLUH)<UI9^>=
aZUeG?fEK(DW3PNIQH4(1/DR)+9.=^(I+gAU\AW6gR8e.D;FM5H/EDgUR)8TeZ>H
52P65O96N8Q,U4^=cW1@Rf<:KC@.N2_g5F.9@F,^ScI4RT02I6#9,c4CS]>N3\9E
X5]B08d&.QT1_;OEOVK8eYE&]F06XW]=0PFffI(dZN13_4^)_RK<&_b#@:=)H)Ig
I\FdVKG\eV[XL&BV.<+.HbX9HBN12NM[>=\0G9TJ6,T2g6gXU47aNADLZ>TZ[PX,
A6UYE6:3B2#J&V&B]?4Rd6VeKKH>87AK4;)S-106_)_7_VVVe8b:_B]-E#R+B.=H
?B-V+a@:&R-?MeL#JCJX6g_/7T4I6bULecT7US6\dAC+6H#QJLGCUFVRXYbX]5.(
LFLGHUU33S/PZ,I:a/E8OYFU^\EZ-5)gVXYFS&S?UL4EF=4c8XR.0WL>IH^>#U]A
aHaH#fPA.XI]H9RWIYSU?b@TW/=RXM[bPGaU,.bK:>]fg\\A1;@Z@C@NZC(G#fUN
PM+FOe8BJ[N9b-.:P_UIVf)aW+0A2dH-DLMZ6MaM36_#K261V>dD:IV(NLQe31TV
MU[8?TL,c:+^;,B1,a0H[4b14)Y-\cBDQ[GUIK:<QPWND<@#&?M:c[2K3M6S+Aa^
8#C8GW.:&@XK#C2/FJ3d4SJL1LbBRFM4D4,,<AXX42MGC5[>D:X&\\B=,O#I:g(R
)HOCF_B]Og3Ye3@F,SU13]R.eG:I)F5[H8W^gd9C9LA,.MW3\2H1;5Z,[(&L=TNX
[LD/L(;N16DdFEJ3:,#COeb@.?AJD[:HO4R-2H82L)<HNg0OHR-&+VbM1c?]KBEg
576/+^26WZ9QZR)YEHJKAK-2/6:_(QaKeZ&BbVATFeYSL,SJ9^4@+9B3fV2DQ8T+
H#daZ<IdBDDE-Xd[dbaB?-<Y6ZKW>&UMRPIgcW6F-dU0=9KNe2\T7P6PR06P8];K
[G_#b2WY[#NSG@37)7.:^6U<F[RZ0SCe1>8S)K<R;3Xc/<^Rg.XB[]d?aCR/[@JJ
#]GJaVE(5-(3=UbcW)7.[]L5dC3R84Og>J;4ZU^Oa>RBDP&CCAQYIG,2PS<WSS:(
H^Z>ef5@MR-Ff::.gFC,FdbE,aE:gLbV^=G2PACA^DJ:540&NGPcQQDK@^545##]
Jg9+;0SXIHP5IfWC?\)LTRJ/)NMHYALW36_39C/I82_D5KG4)1R7N=5MY=?T:X_S
:^aC:6\cac8/2WB##7\9B-dcXSAbI]2J0:b7e7RV4XV5T>[Fe+33g-,d:F18Z&c<
SB0gE6#B317@)1F3]eNNUe,YeC4E&S^-?A&ZXRd,SDU0I4Hb78X9K&4McaQC7AP=
/bT6d)7,.#,7F=ZLBI/OR,H.D:_N5/-MPCQg@#-&JC7PgT?(Q2?H^/_Ob@0^)]Ng
DBM_d^-)33OAWN@XE8O?S#KPK9YHT]WHA<Y:4<G+XX[QAH3[8AF>/1+[YJM\ZbX3
\Q/X\D?cd>H8V3(&ceL)=6Q,\fR573e]]QB?3@H1J[8AJZc?g/OaY;,]\L6I9eA5
:JXV;#NZOP;9L3+/Jg)HOeb/bUI1BM446KL@66_X5W@\>Z<Q>YEITV6>]UeU+8-)
?1H#8FgO:<5NF>VfM(]U7#5VUXE@+dg.P?I?aG)8N[)72,4ZGRIM6E(1)N\FREbd
Dg(AEc&,6-7R?#<]50=.2[B-+;gbb6-:<5G@a\CeHSS]K<IdV/IZH@^#Q0(2:J;=
+V.e5c9&29MC&=](,E2(I.B,WFa=+),]9;C?=CDb^S8f[F#Y_f&Td5J;33U=b^f6
C<B0b0fK&>57bR)T7S6YLXWY^J@HFR\)Xd-L-WF-.A0MN4ed->,CB6&[C6,70;>c
f8EQ&He[#ZHSF[[_IQ?<-QHE8=>dVSJ,EffgQgZ8Y+b(#7<-GMOL0Fc5TI[BNVZP
g.+;YTLX?JTZ@6)\cU6P_O3GA#A^?XG6?=\WfY97..I;5-BJ86GG=IDYQG[./LDH
VSWZ&cS7&VVOP(?aDB_R[6T+f9/GAI5&e&^IU;]M,10VcMX2[83?_E,3KLcf/\5]
dDF>fKX,(ZXF),Ab@=^\6RU9;fJC-WC3Q:STfb-DHe.(2gX,f,6AEZ&c\DYZ:Dg-
^[Z;;33EEC+>fDDN+(aS&1.RXTV56ZY0\SfY)A]XJ;[c#768NGS_VdT#XXS2M@H_
f)AgO64)4YRQ@HP^VA=(/Ac?2OFJeGcI1<SBe7eOCe<1/:ZN6<dUUF3<g=VCGNP:
&/^V#(.[@A3M7\CA<\?aNU/,((d#&QeR9T2GVLR7K@AFaPD^+N5-LgXNX(GVBX\W
-\0GLPQ9QZ\d5=bA?G+.?JL5,8-cC<LEHZUbb6R?ffbRSHJgC1V4P1#_e:XHW]T\
#&)9.M6B^/NN69aQ7&Pe#X&MMb\Q]48GR#fdf3fH\V^[>V^g/>D:_>\bdT]dVUV6
a9H&CMRI;4;VNb_&43/I10MZ9O5.ZA#KLGe?X32N>EGT/_SK9fe1YX+J&KcBcWA=
1K75Zg^U:4,TbLQI99<PX(?#<gY@3f-F3I/Y7.3TWK69__acV<L5/.Ce?(c0X.AA
-37L;=f6&7A>[G28Z-bTb_bRQ>&<ROfEbS>b?eB<0C5E#.FKX7\&T#4GB3_M>;a:
LY-e#PW7;EDd_,]R(95d6XM418ZZJUG\[aC=4Mba=]f?@KcEc^cZGBG@WfGU1Y53
0(ae>KA=&A@+E)3X#JFY:eCHNK4CTV@1)RM8ED=>=MSb48KH>5E=Fd)aZRTA+DZE
K(3HP]Y)36&(952WK>FafG&>)F?A#3VYZO.0BaTK]NH\KG5B9C,S_e[<>(ZC?+[5
bF,BFB5Z)Ma,eTQFT.f[=C_VVW1I]]NT+2<5.aM<+I/Z4XUb6/HPQe1R7EPL-b^c
XV>TQOG)_8_D:.=LfV>;@,_L_,6b:BPYCD0BDM_6]>C@3D:ALc-BAS@+MV>A;/f_
>@,;@6=XJL]M^0Xd_a<<AE+35P]\M0=.dAPL6Z<7\a]L][QIfN[c\Pfec:]2:H;,
JK^&M\)2HJVH]+\OZ7^[ZD:N=Y]DRFgS(1^G=^<H?c1A<.53d(^O;TRb:]gN)34L
L1Ue</XDZ#7AK8>3.]#/\-Vd5#N^Q.[f^D^O_L-.ZL9cD<E5bHT^E+@<OY\,&LG[
,;6Z&K,LOKR,(>J1=I(K.R]f;(?;c#Y8TV4@6-egIV^UCJSaXL)1@IF?M/?H25_P
c[29J-gOZf8cWWUQ+F0e]U\B)FQSKQ62TSVJ\V^WT[^6S@RZY2XfbVM2/@bc@_<_
\_/5T,FT>ae=KY@Da0&5OCPJ^aRZFA#,7#/F/@Z7e7S2_&X+N3K\1OFea\3)NFFR
O3?N@,(6SQJ+]OVU4HaBV/#LVe53.BB8<R:KTDMZ-c)S^@4b^JDT;gCGFOW?WDdO
H8TcJBQDPeAM#.V-ZH).W\UD]_eRIH_/2BVXM123HBb-9ZGFf.=EBOBU2SH_Pf)e
X#P5dQ22NQJ<(<Ue-#D74c+:cE)3.65g5Cd@Q?Mdb\(EDZ>cHV4FX)+6A[O+Wd@+
O/(0:4>a^U9a\4&&fS:f9eU/JRU3b?:b22^@+5:JIAaP4W2O(BGOF>:^,]Q=AYW(
2E08/F:?MUAH<H8C[LE+JT/4ZE-]+;&O4>b_02\GN\7g5V<LZ_BGc[/#HQ6IO:3^
H^#V&Bg2KUP==4ZC6?#g;H;HSfNHBfF\3[0fe,?;D4>PKYM2a00UB6>(Q6[<d(^0
d&];BM_N[O(e4+PcdJK;L)?\F&MPa8([Y6DgMQ)BRB+.512:?ZdRfO9WCP145)b2
]&]47DHE;U-)e\=RPU3F6Q8ET7EV8-LEg&^8fG?;<B)CI)3SMP1Oc8b3=O49OUX(
:X;\T@dS(c\S23553G)[Of(Ad8>Ee&KE7S^;_GXNF8e+/Y><9_N:QXGBb[<:V#0?
\R-)U,WGXRU6c]IMI,1M,#(K8/?XHU[g[=4eJ_/^_Z1MFBf[I)]B>1d/L=-g.I;;
(A@?EfTXVB&BOPHSBg>:_3T144Rb()FI5LdcI3(),UeC.Q7.U..FLXW&>YY)]F56
0I,fS?HN0BT(D7F)B&B0??V+Y3(e707?B+0@,.#b.-)/(>6T_VO9]Sb4O_dKM[<5
1CD1GCIIBXQ3Y1DZ37Lg7HR09I^EYF+EU<UQaHT(3)2;^:D8g/SSZAS8H_52eGf7
#S?-aP8b+T;GV=7=T#/QF+WGU_H&CO,?(^^R<HLA-Z75LgGaRX6BY6L7:H6Q_4B]
Yd:T6A6-=Q)LE@F4Z85b<SM3-cTF_Qb.CF1AGAYf5fQbFFWeQdcJI^DQ4O9;E&55
HSJX3[c8O_UE2#D98f46H>[Z=.DIa2KC>cL0.cb-9cd6)<)JJcO48)Q0>Bc(N#G@
2]d2FSc7.NB7<]FEY4=QYAP-J(cN6]cM9=HYLJC);WEDX:;K-W6W6I8-E_gDEP(#
C:RcJ3)Y;LG6H>D7G_MfN#([@0A?WGJ5U1OW8_Mc0eE9;,[U,e],OBL@7]55Q;\E
YC+L(?)\N>a(@,?&FF?+X+AVS\RJJX\:/LI/]UPdG50Z7AaELB+bW(-/4W0cdJ]G
d3W0g./WLLCGRZDSb)#><QN8,O3.dd+)D)e31KGL_A/EZDA,=#c29bFdO-+.I9Ic
ZA3A8I/c3/a9:Q=1g=ABKT@+#^AEH.\]4E]#NX;dFHL+DS+:J^[L;AE9>d?E+8ZM
Z=>_Y?@AVc(^3BI<G0dY2GdNVQ:5ZJ3XACCK?b@;+=HUe5^NRKg^g@;Q3VO1E>UV
C(HMZ_Q+?HQe(7ZE4#M2T1Fe?5@</Z?Gd^J=8TB6)VD^=T8/ATWZ9FHSF8&1?BU0
b=D_F&;\A]fP(&R;TTWPXPb]#gNf]2eaU40dVE_Z,aP>._DC,V,P#FU_K75bd+/E
#?P\16a18,K]UBH]gAO5eXC2LO1c;TZ+?^A\CRYY^/E2ebRUEO)V44T-NHg+2.A^
39fbQW#Z,UIU-HGVbaW[D(O81gH)WP5^:(e0,?X@fRY-B^.)ea60&AZ>fS.TAHV9
Yde5U#g)6bE1ObQ5V+-eH6)WB&f^#OBTS?F_:d#fKGA(^d-_c.ODX_U]0P:,YAQ,
c?0cPg.Peb6_JC+fNf^.gC:T\0K+4A<)^U4(&<,Le=7;W_RBQc0Ldc6(fJ3[/427
<d;.>2DB)WgY8(,;(@9VQ]c#V;6XRAJgV]APTI/7PHBC6eWR]8dFf?:Yd+MQT-VC
YDI/.LQ#Q0<D)^&R^b<,\8W-FY66UfX[_Z5EBR/D);9?W,)FS&gDUSLH_./H?6VW
19T<4.21H-U)69&IL]-f56B>O811IHA]V^&YDW9\);5)P]0=&V4X1Y;=2O1,GaKG
?fg)OOF(-#^C&EV7MI1Ma(:IRBPE7NgF1ZDQ#I&FEMBJ>06D<cM<4>feS&gZXT_7
I84P9g4T;BQ.]bReg4cJ?LaY^DXRW,/f9(1BXHad<c(2#^1f_/C=C^+3V^QaLF0)
/_CAX#X(U=9DBcY?Y6@8)H20M9O0?2+.48V2dHcL6[dXJ,(<>d=X@@+S,LV#@4ZB
H6&;UC(&LK)P4)Z.@.UH6bNA@E9&IA+8:=1b=IeGYNCNU7M_D2J5HE_4TPO\=c<4
aBB^b:(>TOK7E+[1)?^ce8HQeJ9D>#Q<=0b#2_/Va.G6RG)@CHUNX]BR:WYE2UY]
<b.F/>MLBJ;URNN<Pg(]#BV@Y/H3\XZSfY5XYWDG[=M?g+5@];U5._115<6OBVIS
a?FKK[P4DR(@0G_5\#A>HLA.>L=fWV\N663;Vc]UAf1B.(&;@bK(;?T6CP3R]ELR
J;c+QR7X#d<F-8:L#Z9PbL:N[901Y]ASMZV9OH(16K@+9.IN_Rd8B&b]^9G/Y>2[
?6:F8e)@Nd=1N[M,#E2+1@gHRabIF[_4YWMLS>-3D6A,S=MP&b/9PWcdH/H;GK-6
,O1NE3(+A17<):?#1-=+M/cY3FY]T.?6YBa=B7d.g,:,\T\fNE+)=Q(H\WR08d)]
IH3>.)F7CK49(,gG_Y:Y8W<=>f((M4TVHY+J).FN.ASXUMR#-(TG[V&O3]H\GXT^
b:8e4Se:F:,ZQ3[IOX7]KCKSD-_C1fNO)R^N935GRL(ZO8?>^.,:HH^>b\GWggVR
c1QFL5O]G\>b\Ebe-(<)gYNCU.:A&EW-9WJc1KRQ4:D)6UOFKaUWQO[Q@68I,3-^
HNX,516Ib&:;Z0XTF93Kc-H(]A/W-b7A:3,H5O+EQ;;+A6L^OKG?KZ?M10.=&DP#
IgcP-7Z6-ag^MN==\_J_Q;G3F8?-LBJ1+Z;^^S5WQ,-]Ld^3W[g4_CL)/a33VX,E
,@EPPVP[^e[-A4Uag2_]3^#^77)\9c#\71H9XW=(O2+6Z+;)+UNe(aePe.WL^6F^
:^<B+^bRNMP,C;4BETc_15F=<Jc+ebT?1@T/K>F[56;]84)@b>d-Q(dQ2]/cEB\C
U2E(G@GI/L>M?GW__Ba-(0>fB+9G;1KXZVR:YX<=IU>E#/H0_0?JHgM.(Td/V7>X
-D,C6D70F]TOO#EOIB(&gOAYa7gHNHN0JF9:d/=][R>g4e<WP8NW;3A?Z4.^Z:S:
>WM1DE.[QOCe=_Q/Y;,Xa8^/7RDQ6<8fRJF7g/8DCXXMX1<P,3297cT&&J[N8AQ5
+a=)/<(c==9N6-LD\dJD5Ta:+EVOV7_HAc2]KUDX@dQ3TefDT:CVT4\YKE]>Ia:U
DUbXOYVPH=X;,HYG1Z7-D]N]RV0aGO(=Q1Wf@b3L^2&/e5TFHK.e)J[:aJ^V2QI,
T<P][JKaM3GM1/+d4<)UE@g0DD[_3aA)fT/XbJ8ZfZU98.W.?XB#3PbET?^\2PN)
>VC#EG?d)d7ZF?I4fQ+;gL7>Z9C/gCB@cfK9F<+F1-+_S&/fe,8:>>/FEP_&B>cK
N5[MJIP_<LcI]Yc1BDDD^5.X>NCcS1HFaBP?P@<fJ5e@+?UJVKGeC#a6@]7+G-Ke
8[>PZM-cB.b_OeG6)SeL_R9B(29H8)B]O782\;JH-YC9EU5ZI&XLdZC@7;LHa9AB
C[bTcUTXC?F(TeMG-fCX-L&5XaFZ9N]4+UTUg@S&>Bd;dWKIQC8-U.&-00/)HQC;
=PX(YPD3R63(-YZ6>fM\);#@AC:NgYSM28@IH#T_,LP.[McO(@7EA&MQ--MYW,AO
52\TFe,WC0#=.5-Sg#:L,E;XN0O#;a/:4TM>N.Ff<A^(F;^R>D7E.,P##[+(bM,U
[^W3.MCJ[2C#UM_ea3AbX3e(G2_=:L+D,)a(.=M#_cE<GK8Q\dS/PgOb=-D_dAJ#
9[@LA@O.=BZ4G-6Z,1-L_2g(&=6d)4Bc>3A1K6YbOA<L00b2R+8:8LNE/)2VK@D#
^KZ)LDg(ODeT7]E.6^V&7^2.#4GYN?g6>HX[/:DfRI0cBET(PAN7>#aLGPdUCVB>
YUg60g[VK_?ORRAeZcRWB_]SP(+fIWNB?:(.]67:ELCC5eC)3>YWHMg318J6IY_e
X:J0AAY\0eR1ZZ(#g:>J>2UYGDEDXgd+&]-Zf6UJ/GD[fL60ODbU3P+^M[V2KcN-
W(d^OVfP8I>2M?_AIf+gHXBcJ#(9@B8;cM<A7EcIHL[/L#fG3X.Q<<GgW^/-E?Hc
EVAb([:\24@^)22M+gV[,)/)>c;&+9S3N+C(P-W@SW(/?]LB.?b?#&C)\_P<CAAE
)(LFKNQ0RgbN:aD9JX_I9@Q\FFg#Uee&W.>Fa&F#ORE?:,8;bVf<45?@8Z:1Q0<d
](f/-LH1UYSZX[NC_e<aTT2TS>QPUePcLCe<+3QXVeFRV0@bdD03[J-C]=8.P2dC
gW\G(J>TKe8K&cH]BEgg^O\5bf^7-2gMX\3E7.BT=D]/_(R(__0Yg>JMLI;QQ2LM
QEZC@HZ#L[9]E4(#dQf>Ha:dDV9SI6GdYgXJ0Xg4EDMTb6c0eF-)X[T\]N^4AHgC
6-SWe#K(<3\,SR=1A7Fc^+(OC8-NMNUPM3U5:+H\J.GT,EOT7=cJ?7\ST3X4#]ec
N078b:4.0;bOFQL;:[N8b+U<&d@+&A@gA_,O\K@:K][eUaE-+BS9LF@Id@91ZYQH
U@P<(]__2>8S7YX33=WV^>c-eNb&#0K6KOM.;@V;dB3_a]@6F42bZ#4H)SW\ZYMW
P+/+>,VU6N<&F0];MYP-=K+=^E&^CMMWg[0eU>=e##E3Le7=b;FdVfKc?CZ@V0HP
gHB^_W\OLZHES+K\EUHL[+0+d,?GE,CI4><cCNM?Y3T5Ac/;WGX+bXR^gS>3eE6M
R)9RKWCF0#BeNWY0D36Z7c<OBaXeI1J1):BAd4cE1246f#dB_^</;Y;31J1f8&f?
J^E))#[7g=OI)OQOa9M?L5ZFCg9O3@Y2TNg6Z(g:SPVLE^Y_)bEUf<NOf/3BX#B-
VXfV.>5Be;UHSa1d>g&,11:-4KRIV6B\UA_K/DA(1YC]g_)TS9S68;XdIP)c5U1b
W8JL16H,=7VCagRKdF)Q=HdCI6RaDFe&DFV\<dgN#]59>_)A6VL(:CEJS14249<7
E^\F+K;WR9MKK^3_b[C,@MOD48?M<\9A>I?EXJG[9Y<.7TJ:6cbUQU/LJC6?V\5W
UW[]E83.=J[e0R,W>HUP)[bX_DB1BFUJ@@1=]b>,J3Z:b2Z)H>@acXcVPIALTD<M
=&A#B)D]ENK0Q030QgGDWPDGE/>@e,Cc:]2+60Ue:UY_.E@REAf3^3ILPI4]?9TV
JXR^W5#Y^]IBRCU[b7<b\/bW?2O[D@=(@\4E?,X;F-T9(d][YKb#GIR_+bEO=d<b
58Q/DN/S0]]UK[20PIJ1W+g]F>X\6\-CFGQOMD/RTPG/R2,&fRCR4N#J6cN_VIe]
QA:6:,Rf8(c9#c@B5=511Z&4@^P7K]VMcQ)?TP/#@WP@)B0#e8-d^DS;X6O[HNW2
c&E-5;W.MD,M?K@.2.?+VRWCGKc<fLR0674K8(WZf&6NX-+U8d-AeFO;dQeGA9=R
VUfTJRY_)B#;?Cd--?0\CUCK:2X><)4&Cf<Df#K_ACA3ON2d-4RQMZ6g<>??c:7f
-_5M)TZ/OC\c.UM#UcI#V3;aK6F5TY00McU[>&^ZL:Qc&#@H+9a5;f6,?DM3W^>1
\(7#>Sa9YK[6Dbf.4eJD6d[3SU9C;L7AU3Y5;Q7#fXLR-\Q58#,=P?a2N>Veg34#
XY1&+[J[[Q.^V<Q<VcH5B4@QU4gRbf?L_R]B.-K+c+7TK]4.T&-/G[QaE4PQ:J2^
^MTf?G9HX(<@9].M>W2\VX^S4DN(-CcBa8_fC]c0#BQLARP/R^O(VFI^D+@<SV8]
-f+;@T,).+NG[E.0(&>gHg/0\@B#T(:#RDfD8M@Y:KZ-_NcI]/10\+8,.((fT-d8
N3SND<>V8+JHT,SC6\Ga2=H@bTaa:-8GN?^9bROc(#T=d/+R^VGF.EZKbR2U<06?
UAUT^c>bU1&#M,(_5\[(DQK6?g/cOSQM59SZFZF/@COS/[[\7-3>FA/:a@<ef9]@
5>JLQFGRU72+<G#6Z>H2N3WKB0SP-844AR0A2)81(1W/^M5[7&>3L1RgK5QU<H\(
RB/([V=S\&ZcM<(UR7cO.C>9J01I2>/Q.C/?BA#2O-/HS7g\&_/[-^D2U)31>44)
MLgY82H8RSBS\,2PY\WNQB=@c1bVUe^<)Y.;G:FQ.D&I]OEXKMbLJA^1WQHKg_a1
B_0IDIF5DSKYCOVc-0ONTW1UAO7(2e#6#XYg;:eNEB^K1(U.AI0eP(&0>RJ:>DR7
2[aZ3.#g\<MI)B6aD6\e6eIV<fTTcgV]^35^#eEI?J]S;@DJDR@B,4=YWd23\;,,
@C&<2#V4-aT;dCG:I@:#cbDEGT5K&VZ=c^)_4XPe#@7YTGMDGYNa7I&64PERB[LM
>La>b6F5CC\0+4aYHeCU@<ST\Fe@D6OLcceS_a>d?=:Zg9Mg=ZITF@ARDIH-1@fA
ZX(ag^;4S<a[])L2LQ(/T>dN[].YcP)2DBQJIU#(3RM/DU-6e]8=eBR/Q[78CT(J
YKV[90][fXCB0L3?gd>d,)XN8E,XCT;,S;gU9YAeGBH9@,NW_<(:35,0LUJTKFS/
\TH]Dd_IbAU[ZZQ79d^UC0,-?bDDUJ69a?COE0-.=J]g:(FRT8HM2[-UVXe[-EV9
ELCbQBYEe:bL@R.>=2b?7WMaCY=;cQ-Z-V?[NJ.1/fXd#LAg1aU&-0KP<^d#^_Zd
YXgG8-.VQd<1[ef1-95;XJb4UG4E_V]e7J\6R;gE9E1]Z=_ZX7=Bfage;DH+:QTY
H=M?J[g0O?04SPM0K;Y0aI+MJICLg/S9./U0&Le(7:R1C5HL/C;Y^/H3K/@UWF>I
?O\\^]&Tc5K=&9>gM[[[eIe.JRJKQFDS>fWEG[_c@2]?a:C];_Q3Y&/VO=L1>CR[
.YIW0689O4>6CWO@T3<H+X=fKS7>K_<:fJga/G+2/e2RdS\7B/765>-QE3MHQM9^
(8R/?<8W8O3B>=\NYR.(<C1D?JLL?@PE1,56MCdQ7&0B?4I,RGX-#/WJUQ6;U(BT
H&=P6Y2+=+(\7A:GGA;.U&VgXN.0YWE05[]8W3,5<8JJ\I>0g/I4NNHY,5JZLX,/
e6<#[0Bc/fNdVAM4#TU<S?AB/:F.YG#X4dI8.a5TAX6P^@ST5fC71HbV9f,CQ.TC
N-Ac.OVNf^W\:DdW8V.OR;]MHb1>deC?C(+b/cCPJ(>EHW#E5KQg^G&A:g/M[12[
1D?X:5A:RFG;e(U9eS_Z9Rg1TJY^Ce_&J#HAN#IHM?@3.NaFH+94#VKL(E@]KWFO
P.=-eb;169PZg\\C_\#7)75<4;_IO8AT0aDbFJe;c2gV:^S+F1(>32c-^bE99\0e
V@,Y^/384E_RZ+8cG?]PUc-GBB9XUIY@H)0??-L)e\HI>PP?6Q/Ue7]d.\Kcfc#W
],94=GL.1YA([(,HVGBfFQcVKLee.1,[RAER8@L^V2+0@19@=Z#I90C1X@;T^CTE
&;:WF&&C-&Z/aBD;cVQEN]I1a)db/Vd&A-P,DY#<#Q2PJ77]Fg)HF>>g:GCbRAdZ
Ufb^71EOGA=\AeLJU/Wf.-1=P)/,MGO8L5PPN]1ADW&?L,-1-EL&7B3#B1G(TaA4
VMCIP,)=6K+c5fNb/MCC7KS_O^+<\gUD]L.GVLD/,\:\[29S6MH(C1Af=P?&V,#?
ca(ebDRLPOgcDMTC+;dIaT=H-NC,[W\I>\>3OG:AI?<#:0GFN^B]X[g?ZZ]C&R5O
>6_c]D&1XH1HEb<?\T^.P#FG]Mf(>P&=)?GB/Ud@cZ<7dKd#S6=90eHg.GB[Rc<F
<P<Y[QV42EUeZe@XOaWdXObIOGZBPEBg5J+5-_>IcgE)bHGQ[fa@9>U<5;&R[g9C
Feg015<NA@[G\,4H,@_dS/BCg:Ea#Ub(=DM_:+XT]\EagE7=S_\ZO#Q73WSA0T4e
EY+;RWHH41Ea&3.L^HX?EN)C#/E?:_;<FfBDD&]DfC\>@JRb>8Aa6TcEL[HAc9VG
:dgJQ@]FI-NK=M.Ja>#Z1C[21SGM^=?2c0.Wf(759dJA,FCN<E3QfX7?):d.?F:L
0W:1FLWP)gUW\WOHS&2X;L0JAYJMBEc-CcYY0gCfM09b+QFe=XCBCHW]cD5+R?<N
8A;DGE)>98&eXZ7f)Q8Pc:6W2M2JcWFEa31Bb+U]D&X;A3a6gd@6dUO#3I,^?0IF
g^5(KeSG)9W;+\eF=(]eJ,^6JG^MEcE&GgRbI7+W4H8-KW1RegA@2ZZ@?^/_Q,JE
DC#4U(I89c9dHP>aMLG?Y1\.b3U.c3gX5B\A^:W9ab(I[ZBXd.E(T:D/78FOY6aV
(#d5Y4XE^0/dQa2dacNX37^E?Lf,W<SH)58>_2ZgKe<--TcXD)=f,OaSW7__.?b0
&QKFM3\CNOP.6W=(I65+=.K&I&/-+:ZbZ^0_A3DL\5J_S(A]17<Dd&Ya^UJbBIc]
<g@^59D[L.dZa@O]NYHdB>LIQMMWe)[b_?LD;I-?&110C:d9,(UCQ8KW_=/4&BM8
O13W3Ng:)U^]]=Q8I#<)Q1Ya^AL;;WR-NaA]g.67#4b)GF6)&RD4V(MEJJ(1D_?S
c<EM0E:0PQ<#?Lf7Tdf>OI00\G@/QQ8/g.E9J^:T<U:dfc->[?R&_4C[ELN/7UXV
J2/GF],F>I[W(^G99R=0bP)E^D=@N_?;0F=P\1PCf(.-g=[X/5#JA5M>1EgIB>@K
+dg2Ab2A92)7W#bZG\V@21/GAT>8Z3bO9958Fa7e3\TN2GG4R2Z]]RE1XYS--;KW
7J&90ZHI@&EbOD/fGVd]6#];bO@UECg-Z?:9]E#/82H.b<fF#.4Q].YYd4)T,36.
<Tb&VQ6OFIaG&.#FMcd?e@\b[>e=E.]^B/NZ.V282.WUf<IHYA;G;]9X>VDPGbd\
BaXAQGa8G?^AWKcYL[cQC[ASd4Z2W71X0)bLZUT;BgXNa-E8T79C?3LaORAI0bR[
J;Wb#b8Fe\L?2)5Ee+a)MLSR3^HCLSLDBLcIOS=QAgR-.=Q/#Lg&+<O2T.aED&8C
S0-:]&2:U(c)1N+#QTMP8W3KgAK]\EWCLE/@G;?a1d:<K9fPH5-MWfF5gYP<PbNJ
aE2L)Q.gZQ7F\U&@5SRX95Md^:EM:EM)/(@_(F#W2K&KaT@+;0(9:eEOX\BU9X[+
@&69ABJQ-2gV4405M/3LS<&Z;08ZMc960OAEJa=61=g&S&db=UdN\8UDU):-GQ9D
&-S,gD29S>DF955EC]RQVH;/Ta+6=SSC[.=RBJ]U^C]Y/1PFZ84/bf#N92XeM.U1
;:EJc#=AW0H)RKb1M^A<DAN;ebU>+1LE<feQV<<7-0@S_DW@>-G(K(eXH&3@BQDS
g7_&^<D2..f]EWI5Ge=V/;&gf6MWN<JbP1eX&[_[_7(ga;6ON\>d8\/;R6-=dNeb
f,7#DNa[cf[gZ5&XPT3E8]+S:dI++TWEK37,dd+PSO,5)D9.0#d(G\=b;@CN##-S
SR))))Y+KcNQ/Ua9ZK^.-T.?<#5=8P.^ZF83e4LE9D=.[D)UJQ4493]SMNH5)UKX
)UR(SL.T50J<.59Q?38bFXCZ.#7La@GF@F.0>/8W5d.5RQ9&Gf.JBZFP#WP0e,N2
Gf_LDJXZQaA56NQDP(;9@])ZP>J-R0R6#B,G0BQg:eMR;QdO0=5fHOB-:6#Q6Y4H
JS#YaMgg79-?\S>Y(UJJ&OFZ0EcAS;N4X&,,FR)^ERbZ;@NH]LNCLM1B[7&b3S(B
,8)UdL\)\a+.?7R((Y/9>@QO<N[#-FWP-,JF(D3=BQ2A:3Gf.(W>ISW[H/(Y-bdN
Rc_7aaE5\fbbYR17+YgfW#4-Ge?1D=/8I\LFF0)Y9?BUGaAf<<><HR/+I=F:OI;f
2[?)Q7#2+Z]WC/+>=Xc4,]g8,c_L8&+C0_X//<,_V9<HJ=DMVbRaIc6e3A=6\Z=-
BE+8_Ib,@[E/f70T[FZ_g9SbI9.7g12(YD3R3FN@C3;]FQ:.F[QP/5N\J(UFdTY6
F@#ZA)F&Z^;6D9dM>:OKD7JUFZUd7=d@KS;JeOPJ:;7;&DdT.9O)TA?8e3=5fO^P
B_RPDD?a8P.XdK@Xg@1OG(JL]Hc5Igc<[HGLEWQ>?.<(K^H\cgf20eG@^-aNP\-W
ZGL[&g<IF48.6KX2_\.)QJg+OFT2#;0_-1^_?\MMPa6QH?V-C4;JM4M43Q#K@b,2
0R@ba3B\:TPZ9]PZ7KDLDPR5/1WAc[<5;gHDG@7&2\WD_-0?./(78_4eNSL+6aH^
c<a>5@#,aCTE15JE6&SG+,O2&Q,d,)5f7Ia;ZLd0,-M1?V-e_7[C.2Cf9Nc/GAe=
D4W^a@eZe@^;:H=7YB5fV[D?OW[ZEY8cdYQI]b0KLBQKT?+e95I:MSC=^--9_?S3
1<>b9L=/]aR6/;S6Y1&U^V-D-J5-SA2(1VMDF&U,@AI#b+0d3QSHZK2c4#cE0((/
#_02AIK:fGQ:LZdO6QeQVf2H3ER[(E,#3B?Z\)?8C>:fSY#C;e(ZS=\Z:@66gR77
B#8>2)O/DXF.DJ0GSU=LDSI/PQ]<&T?6O(7XW+Q>U?:\,^[(7TXc,1J/X8V(GfO0
a+MH[5:ZZ7B9CbODFTBKc(X9&@J5UE\(;X>M=bSD.;<,+C@?S[bB3^6^O^N_VKRB
)2GW(egB#BWO8L2P4Y:2OC>g#)VUb5J9F3]^+0MFW#f#HK3?bN0=cU^TQOF^ACT(
)Vc;G4+UcbOMf\M>O>ZW9/(OCbU0H/R.c(I@/f#?)3:aBZ^MNOG<(I(\0OGc^ZE=
,ZA=0&7a1]+[\]SG[AO)GBRPgSQ/A_#]+8\ad2X#..fb-(DM/B6ES\645P8dW=Y:
A)&U?W;+-B6:\[<SNb(,^[7Ge/=#e5U^.LIT>>^<7:<gd@@0Fa;Uf_A3gE=@UJ-B
A8HR2+d;d6/=C,33Z=&^79QA_.MVbd.T^E]E55E]^H8_0=0-:D@Ae76Ja5aZBf(\
W8LY6Ia-;#8FI1Y0_\DBIdW1af5JHRMWL^0Y]]B\\cgO_K3HdA[314Z,>-D<2XWJ
D#aeg0V?Q-UEI>R+;0DYQOC?WJD+g_[H,32YfEY0U@E,99TKLP;E)UDM57?>\Z82
EM#e2M-Wc5B2_.W0O+VeM91FU_^NOX-ZgOW(g>(LVJTQ+a^]+@]T)@<1=FJ@3DW/
=[)1\@0J)]/F_KM.[QITJH#=B-RTREN0@F6RZ6[#7,JE6WGe)RfG1VYG.+f?]COW
JI=RXb-)c\V.3QA8_e2Q.#)6Z>U;I8J&-LIR]d<9b.4(]8-e6P+O]US8cA0VF:SX
Kb-A?gZPBAa)XHO.U^)G+8cLGN>K/_-KHQ@U9J7C5@JXK+b_UJWC6V)#RdS05^8c
HL.O#-MZ2\IR;HKf7._^#M3].&YZ9;@dgb\@C?H./D9>;)=C^E\K<EWNIQWKEf^H
I_F4AE]Z/OD+e00_<P+2^+g?5Hb9])O]5;-_F^9--7UPeS45YTfFO/?XB(IRa)]U
D6=Q#YT-<J)S]<FUX>:JZX-aLPSIZ5dg+A>Y#NZ.aBe1fB89gdZU/NB7@=)<#cef
@]\Y2ab#-(]]c^,J-ED.=+TOT55Z:G-4NIOc30[/_KIX(g<_;@_JVC(G)>G^ZO:a
ZFS#>6(Q9d-X,BU<]0#).S0S7P&dJTBg&U0BeZgI=CUSMLfZ@T8+PUE-TTA(ZbK8
@KDD<WB[V]R)-(ANE&.eI=Y91D2D1g2)0M-96fD+)F4;+E2RYB5<I[bXQ+<DdfBX
-[IAFT11YV##X4H?H+G2eS\G956T]L?TC;.2L]-ebYV3PPJ&.PED8<bfQJ7I9dD#
LPZIIYA,A,3L(-)^Mb)3R^6PC2:-NRQ@V/0RO285=4\@-a+:_2e?aVIMU;1c#+S>
Q@V8dP8Ee)=3=9dcKV4)3:9PQUc37f]&Y^0Jg:T#ZD6-W;WfU\R));16O+4RZYgP
N]IQ@Y.36F-KY24Z-3Xa^]N]MIP5X)^Q(CVZ^]JBELaXXM4\+g^[FVd,>0Y6/bOM
(f404QC9b3AJ8e/\CZYYe)VTA.afg1^/369\F)Mgb;f(=EX=HV;7KZOU7A+cd&/f
CO+QQ8AQMX(T3Z8geDI8.c,SG9XC3\7bad2FFGS;bW.3F2@5?;AKA3,fWc-9Kf?I
)UIaBKMJb142eFH:XaK>OGZXG[bZaE1A0eG0e1)KNU;#4.3MTcMA4JZS&2c1\3]&
6d+:&J4Yd1+787^5dTXO_>PN:;4:2GT,:[OBG8KG#IRCL.,XEeQa)))&527_eDL<
Y576&Z>]NY8EN9YZ0S=78@L1f-/L]5-bI+_9);d8eG0;2[3SN19PU&X[,+HXI>.A
@3&c+U(CGQ312753;LLJAW\FV&P>-O[BfJI)V7b_084U=)&C_]K&0I(9/g)].X0N
A&&XL=2GZYeb/T(JVE:Jb[ASAXK>0((7B[(XZ8T&&QXc3J2#2CHE<e(fY[57,&IR
DW4-PAWH7,VFM];^4acW[IWT)C1J+EXP_FAbA1Pb1eTI12F-7+a:#^M),3U2e#/e
-&+98214H:/2S<?JFNg+Q?AO9/cZE8Y\Q@ZU#7OCDc:UVd7EI2?G,d3CCY)L?Pc1
:&)D>L4RC5BZ;<Q2SRJ0ZIb:]2Z_;O)6G,1;NX2ZKN^B>COe]GF([@SXUeJF4<U:
+B]YgF,ScLO;.,W8)2@Qg;B:C0Q[gc^L6?\P2;=R)dO_,\BP=.4TBMBVBQ\KD)YC
/EWNOP.PDQ(]73:]&BB+EKa:IMga(T50geIW8K?@BOS4;5Z5HR7Y2><UT=+dK>DG
g^V4dP>(+H7^^a95@2OF[/4Y.B&QIf;,ce>OUD+NAHH8@=@E&\M<c\N34[KS5G##
1R4bTE4TFFNZPV[:@(_V6Wc6LD)9RdOBXRTP5VULXSQG8If/K[)15B:fFe#X^TB)
:NKERD(>QAY720RD8]Fc[+Y@+VbRZ2R(67(:aL.@HG7N06c-:,T)@JEW4c+,WZ9e
DN&6\<e&fb/0&^^>:D5?R:\SQ(7V&Nb8FeP0G3P:0;#^;:2[[B7D,-NX)TMOTcFU
^]67/R3RZ?_cT87@3?Q>RIILN31:O#CLRQT^KbedHA?Q]g:dg#<,@-Z;]P<;[7B&
G@0NRHKBJdReL>U0?R0/]U=JW2XHC/2&531Y>EWfa<9Ia,2H7LC[3CB_N9R<4RGT
2@Pg/2O#+EJMFT,58I,0PB)VF>OVMd2_Z0VDLTc-K2eM?;=)M&4A:)=e?#RCZTa:
CV]5ZP2H>-BI<5,+\,c.5]aUgNbHRU^QA,-/#;Q))&Y=4;1N8IB[K2Ye@YGM-8d(
W3ePBVVNFM0eX+&b_DYg^+\<QC:XRCd@&/B/NAK0U-BVZL,N=eDOg(AFDdJ8TaC9
K[B>93f;>?#aY\Q>Q@RS+^S7N3dfFA?N2e^RDFY\H-UeX2=2?[YNDbKTNGW9>)@R
?)O^^M56eP:S.O=&Hc#2b2Md,-?9RFf7CW(gS:>[(dXXRPWZa-]04Kb):FH#HZ=[
5DG;5;9D=dQ2E\-=N8C+D3YV4][eZb&DX.:HbOB\P8^_b+1bE08IU04J]H,:2@6,
5_Y><0-3X<,/[9T)L2ETIeBC>c..QPVUFFc-9613[g8P0Z56?EWG-.O0VY+=;/AK
R@L^@GD@V<GGRPX=JYV-SY9X&45K<f(?EXdEBPTEcA-&^A.89?<IVYS2IbB.ZcS(
:+TK[77<.+5QZS8F-.7(<@48-(Ze;f9T?+,?VR,/.\K7cO3Daf<JREZ>2+Id48a&
@c.8-V9eY3C]FTRHW#N@L#2-XL_7XT>O/6eE,ZHDB1RYI)Kd^@@-OA8/;EIVY=QR
6Z@c8W08)Ec1.BIMN:\[WQZ)EVESb0W:WYQ=PCDV+3HP/EX1J@VNaDQPfB&,TDVK
6NY#5HH=+,7@c@9(HaB=MPM6\5SR1RPG/,c2=J@GRW0LRG)_O0\^F(<]_DQ&0_Pa
^(3-]=aG)[4W5(J+e@>Vb4Ka)B5-Zf@ZVW/OOHXH6F&7AaAE_FDX7:?ec<]5cGd#
EAVO1^OS658BFUM8gL9c_@#F^JUZMcRc;SZbJ:R2Yd2#S,dGEX/E[S)N+NY,HZcd
UAXD3^>>/cDGf?f+Y+GG_L6DXTL-UFEZIIF\S6>UV;<Vc2IdC)TK4c<f50ZUI^0Y
9\2_X?[d0UC9FCO?[=:@P4C)ND@c>bW(M#fHZZe4CeYG,+8cTVX=P:V]4/E//)NM
@DW&,VdZB\ZPS?U0f<FK(U&gce<G(e+@:F<[BVf0R=V0H#+L-#Uc&&5bG+M-ZU&g
HKOc490?8d(PVA96]g4aT(\=I]^@Vf3FE_HPPYX=Y[_g]7<Vf7/;+e@<VXRXZ7WU
X\>Q/F@ULMJfXeP[e-]_cCYP&?(.UVU,J#6BS1_#Q5)Rgd6(]V1+1ZPIAKZ<1MUK
3EZ9T6^1\4a@P\CFb0FNZ.G[U:C35#L50/KIJC=\L3B@>=WL-2DM^W&B4?2\<WQJ
?E?,AVP>UfRP]?H^1eFIDd2cBJ;e9R64@>JIXL>bGC2NIebYH62Q/OY[K4WX5NZV
N9(bPPVRO)P8RNUYJMPX,PD43YZ5aMV.e<&W4d6RZDe6aSG/f;I&6BJd5E/aIA=.
&]bX2I&aI:aYCc0L_DOT((+09JLZGacJ<;LD+aDX:7[3L3DW37:9.cd7&K\X]FeT
[3e:IATDdSFC?,DAc-WRS7:]1Uf9]VT/0Kbc<F<,.3@5eR#06)_Z\ZN,3dGNFLIW
51810F1\IEc?0P2;b.\+&4L3=7SA7ZFe+F,eG@8>47S#?3a(@Y.Cg[5(\WWPcDAg
S>RY-84=9Y4M:aM-&R[.38ZYOg\9)).gbH<<9:f3eL:?:P#]RVRX]&+SHUJXGB[R
2BV,G<IDD[4]^G^Q/ANX:@S.UQ3YJ0_Y0<V<.SC/#]8(TTXPL?W)fQ&U_#6d]&NU
E7=3_:/^]H]CERWDBX,;-g&P8>[3L0LgLE[/0M;1#O;P7A#0FEeH^1LW?UY?7Q8I
_.Q?2fE#7LE;;>,T586>?6-SGPC4-,=./WJEfa;WF^0>+QW6dC/U@Nf.T;G2](VM
VaZ\FE0+.5F>^Z(77?VIIL#W^2M;f0[[-]D2)_aCC+ISXO^,JJGQGAeTZ,f5d,;f
B1J^=7&&@f+F4^6-ZUb;1(f+0N8Vg?<Pe_?ZEGP4F76VX8RPQVDPVN:PeGLK&SIR
N]854-#X<86WFQMV^d[;?6:7Z_Hff<=#:3^95<7,(d6>@IY33]aN+17QEH:YU\=(
IUYJD[NNKFPfIES^[0fM41cK1?:,.7?Z?Y;2\R@,Tcd:\CQZN_M#Wc4PCH6L/[D4
FHX#N\Rb3_e)?DeIQ/>LAK#P17^^1PU?(XQY4KVUb.[SgX0Z@+/DMAO6>Q-4NJdA
EJ^,RCX1G8#:)Q1SDg\.F:9FaBG]MG3F;&(#T8;R5_JgbZF2^^YH2X+2_Kce.?(8
LH3[Q1D-;=2>_2g?).UEYOC4Sb<[631DDQS71?GHa5VcD[6VL6YUBCAB-UWUSa&,
V)Q_[_WR,MZBPZM5ZL5QA::5;,I,P9O38-:?1OQ7<F<FICF=YX2,])5R+\BSTW)X
+H08@=^9Nf:IOHSPGD:034EH?2XP]d(>73<4X^I9C\3PV9H>UY@Sd,IDTZR];_V8
PB&1Rf#V0]TMI/YREI\N:5Gg0aMP+agZbD=9b1@/eLBWXD]82\+W\97:DdWP\Z=O
IaKKc7RMV12JY3\<.[<;09<JSaaF>VE@W/ddT=T8d<M.+^dc.>_@UWc,I2B]S#D?
Td[Z3F]:K_Q=F46gUS#Gc4HNK)b+_gJEESd,?^F]fS[Cf<RRg)HA#+N-/[?Z:7(2
9)d1<F5PB0^3<P?>6Cge\[G?dMO&0:)4YSS;H-[\2gQ)&,C;J=V,XHG0V(@4</=H
@O&Y-X_50ENd:3F>eMa=fe20aWUDDg;.(9R>N60Fb6OW^8\6P(?1]UdG\]d>\Z?7
S4bbQPQ,<#G]LBee12Da-CNc@4<7+Se[:N)2BD,[1aeROXGS?+7f_8QM+0DC0:1Q
4E91#0UQ&4KQFH_g01[A^D7LM=-&7Z<0g&(PFQF9f@UHZ>Z]PPPUZQDSXI84K[b3
WW84b+;=LTg<Uc7:,6g#KQL1Hc=b_(C\g/fc>#RH8,NL;O:b<W^[MYXDTaGGY+/Z
d1BdWVZ>N;E1JT\KK[@FPM<[J,b5fJ)MJaE?AXg_a^H5AMgZ-CVSA?Ne:+FXX+;5
d<RAA)PYAT@)T<,V)cFYTdV)4[dQX>IX5FW;L_U)KY0d-5YX):d6gDXEKd,CV<_&
NFg@5)_OW-TfUZQ(K]=9WBP<fTa(;g.-(=4)L\4:1:EfgARMH[,SL(Q-SJNG=^ZH
g@,Z-419LH=6EAQX63+Bb@2B<8-I#b@G:\SWU=Uc8ZaNZZLdAU)37^ABe0=N(]O;
PLLZ/E>5YAf(W\a>))[)XV?[9g(@7F1b01NXA9WB;(->9-[gf,5NfLJLSd)b:BX.
DTJ,@XUgCH#;O_R00WbD#]a8=LWRD5BV7)414I=Fc,0d2a8#_38?>_B_=-)AM_Mf
Ye[O:NZF_S,JVF2D<g:]#-:_52H=(._77RNY(U@=>/U]HY]N[8Jb2bPR[?\-(2:6
/b(f9^dOD4>e)D+);?L])(f&APQGO[#eCc3cJB<=2cOT?-GK3F5@F2)PPM5P&b5X
b=X^B&UR<A-T/<4f:Q)8WRQ#2KE.8W1XVd\:_XJ@P>W0=]fY_6A:VG5gO/3Y.g;,
e(9G39(&FI5TSD;L1/,^.=BW,J,7+-+Q_4VR[MFDNI/5@462+/>;8L<bNcV^5)+J
c@??fE-+OB&3#TN45+TM>)O>Z6]^FDD-Bf?Ef2[.2:89.a#T_aI@9)G/Y+GBBP+G
R1XJLHRBAFd(POQSG&+#:<[69cebNAR,[Jf7RY<I8C7gL#YY1]F\[e2]5RH@fc<T
]Z[L+5770?T64W4E2bKR.0X7]F]EOZ=3CVcPQ5AC+M,L8K6[&JVQSNX)HQ>-U+>H
T,.1.]DT,]bbP\f9)<?3+T(-V##D,W<V96X3G<<=2;c<7D#<WY)S9-4fWU76U^eN
I]3-@4Dc9_33_)e\5CL8PUNcLA7eMURW8.,C^gO;R1b[3J+WKd^YOHe1D_,fH&>?
W2B3+NM6HSDJPcf>IGPH[TSC<:OF3X2N]:H(DfOHbQ;7=ZYdg+UV2:Z]g84gOGaQ
/X^^02:B##N?MO7^1a^6eW1?&_^Y8174G5@)#PE(=c5[^Q]HRWZZ,B>24AH?4[AT
=M99\Z5OP\AYDX0b0@BS#,5gSMD^Q7&N^UBdVe4TI-5+MJF^[UKN;\S_K<<@QW+J
,fS<G^P=<VH?4:_69<Oc<eF&JA>5cA<X_2K:3(7\DH,JDNL\E1:T\3PW<I(Yf>ge
fNKU/#KEU0eSN,G>W;62)@GNIZE1.:4E^4V@BCMZf#_&cc7H214M,;e<[&49HaYF
ZAMH/[551gdP-_g_N0\TJTS56Z)OA<TSRPV5C=ZFRP.5&\gf(R,UN#INdE:f?E.8
34<aYJ-JW\I_R2I>YgP17A6d6dD)a9Gg-+>OE/BT840GN\9#2EK\&IX697[EP301
b#,285>V>-6f]_OGO5C,<<J^;I#:0>EP^[;UG<2L]>C^2-27;.SX72ZL]fI>Kf//
B8dW,+BH2^/Ng87M7c>fE),2&]&+@=B_^SPHQ3IbA1K&F9_3dU]+Efd@,AG^DgR+
HJVcb(1(a^S[YAYLGX/>SMPd=OR^b#b(eDKa=&R_<C6)-fHEABU2M-W-QN7+J3I0
O0DRL?c&Z[VDAPCJ&L(&f(L4;6b:#UKHOQELJR_=),QTW7H4]Y=)OD21K_3=]-AX
5].;d>OZOCS[JE8\CEIH(MJfQG\XDZM2J0e0+.@A1T1(=8@XF\RRV62dX.d@V4@A
HB0K4XgXY0:;eb2T47Z>;T0A;L/G/T77E])#e1J,MNXL_LfPPaHKT_7N;7aY/D=>
]SP[0L?5LaAB?-H:HL1Y-S[M1/P#Oe9)I05,])EUc;N]a-DgV;U\-:\E&5YfbP2<
RdNgHZb/;75-eSO:b37f?(XCX26G]#+QINQBZ[P>J\D8]H043dRJ_Pa/^PM+Q#R2
E>F)e7IMfeI0H1\KB^-eLS6KRI.?;^a1,_LP@3JZ]3-/O,4)9eLEPdBD3YL15-e6
=eOR4Dd/7TBY[?GSLLbXNLW:6\S#FJ5AWA4^J_:[9Me&f<IH;XNT]cJcDO<I0\B1
cY;00Q/RbV03X957Q:]HNX_(d507P8a+GUgM==X+5L;:WY/7/P(,A9KO=PWa1,(O
H@8?U-CF&56QR0=:PHV^(/G2+b\f&LQa3;IVLFJ2X<48Z>,6]H;1TX(T,SeKTR)e
C5[U-@L?,fKdZe[eT\Z)-_QgMgJ_YX,[]Ud4)9c=C/5X=:&C-MI;UGY+3LF&/[eg
8c#3-PVNA06Oc0KMUO[Y>AU9/;16Z/_-eMdYDUB^&5@b][/3Z\1SG4KTH/VBA.c3
O19NED4b50^5J)Dc.\M+OHe3+=BJ19BFUGD_)2S]dYLd^H(6\:)12:S?D=b3I\R2
Z[B>dZ6GAC?/E4Y4+B]C&5EY3McC9g6V:0@bWaRAS_XX[/CJL(EREB,#(c^KJ(U/
Of3@5&bOM4X/MZ^X2CN5E.g-Qa-X&@RC3UE&:_#OS\24<Z0+^gX5(]W9C-H=6O.]
cBLL?[<f-4A=11^>0?H/T(V;<(^L(^bJ[<HO>;(GHX[>93WV9gG<7-7e;/L]F5/N
gUGe18MLOgggPcfPD:]G:M62gPB.9#Y8R0G(?)JVZ:EC^C76EfKSCOZEP5RRLIf(
,KINJ[Z45QXAQ^4U6OX8Y]Y0<V#S>/1X0F3R?;9gT]HJXF3fC?ILO8:a)d_FBP1N
fPZ<OZ9#F?QAVeC5&cbcM>]5cI6(HE\d5Y4HW.1,PB.a>V4LdZM=:R=X?U;fH1U#
7MR7dC</GaJH_f(6FH=1+I@2MCT94bABf;gV>B3;^eBQNFS5Q0E(eB\:;Y3?T66/
NJ&e8Y#9D47JNW8HV])@c]e0cF,[B-B2\PSK07&0(#PFHFOB/VdE6@La-JJ=@_dA
I(-2C42<Fa)TRfK<<eSK+cHfT=0WgP9V_M_bA?;5B^W>;);&;:=ZF3O4V>W1BMP5
7Lg-15c<@[;ZbU<[6J1G>H>CAGHX[JA[[9IPK=cYQMWf6RU2+]\ZgN/-9gRNIW)H
RHE7^\J9]Yc0Y#7^^&ddEc=B^HBL\gH;D:TZX]Y,KV&?R+\_?FN1X,(,NMVJfL-@
_7E1D8);W_=NF+]UHM7P[0^B04LIb7U;T#CYIfSO5fXL0g^@YGeAcW=aZbbIR#6Z
:WZ\F(5W8:O\H=W^B[W?=fFA>]NPH,II(Q(Yb=(=.UNg-CX#42Eg@Kbg?54[>[@]
/4]<I]#W=O#Se[D1A]QHI:IeZP9<#:?fP4I(6/X9IK;09aGA4685O_V(bbc6T+5<
GD)+(+Rf4&8bJ]ZD7MKZ_N^J@QYXRQ6<GObQS7OP>Ub;/KY;cRb@WR5U)TPVE^X=
/bM/cd)aL84><JE+Y+NYLEBBM>8_QYgfCGaJS9([;OI3dfIf_aSI)?^41NgTWVB_
f^+9&YQ9FFWbO?@bK;V=YcGA[VS-e<a+?0JT7KS1<UOfdYbH5+GS\8?G-f?]3cMX
CCW&]EcR<L69+9;1KXU?W]=CH\feGOJ_))33QZ@TM5NIS@EPG+0?#JB#=Q4gG]>@
eOI.J3JdGL33+P0LH.Q6:Y?;D7N)0_gVg=UD[;JB(RS2<6I5F9#/DT^:5PC3eU-G
)b7&X]J.8[dbXc4\9.GFCcPVFA8)+YQdaS(V(#/B0,OR6MM\C7]GY0V:G\48DIa[
:_Q.Vfd:UCG#SIRB#@49gB-JQPH(-,6;TBFG>GLL8R/SLDT,;R?(QJ,a/JdFVcTS
2-RU\LF3eTA6C&&9X90Y46dX+d[V\^X=IP8,MK8UK>K:OQZU(Z:G(e&aaTC[:_0D
Y0)3d&(KW^<>W9<WQ4X3(ROLg;_QCdY;G-HERb3?V<b10;[AV+0C[/49SRdU&_J.
3D]b<OEdQ^3+Z5a\_8B,e>JJ8D^M<\dFDeJ-Y5KI+]6L4E]-8=bI4U+7\IYCV53[
>fJLQaZ1CFAM[]I/+/>#R82gGIPZC3.eX@)G=YD>LCePI_9d0HdSPS.[4LOFe;Z#
5&UOKN#A<QR(27bQ&#KgX789696W9#L5N<&7I+)5C]>@YfIN2ZB;-a=aR,/\EE\Z
>9:/K7/W]VZ;F]L>56(cdS5@aP=4&dO9X]G4Rc#G(<1]W/0WKKGE+;3(9DX4Oa=2
.P-EP6YXRDNQC6SA:#B&Q>H(##0WK@L[.Z^1PXR0R\/X>#JN=F3#-+1+N8:KW4.4
R-d>CKH+b=Fb8,de\3P.A&,O\97NZegTaRGHT.)P9DL7E73O=R/+N&:dLGYKWf(Q
)T70/Y_7UUOJ^RdND?H_?C+#;BP_[9R&gbBQfNGRfb22JfGb;J+(gg0f9683<\4/
_U>-E1a6FI@4?+D@K7gfJ,M6O1eF1MUXW-:9JJ\/&\SZ@TU7WGVZ3Z9gXKW7H82N
Z(,?Qgg.\63MR>CJO/)O?,7?:S_JcGGA9=+==Z5^>:0RDL-G#Ea+d70+,L#Pf5R+
(.c?OP>;[GOUD&61TX9#_GeS)OY7d<>G.cR3E9QbbD@XZ=D2f^H#</(-f9b]G<YQ
/8b/,,d&MW>/2IPI):0?8H/+KY/#:2\Q52^9P59fHM7>VaVf_IAIL7WZB.0B_.1A
J\K2f-+UL74,B^-+0JM80f2#\W?@,Ie>X@;7C?8/5_3SI:Z?GY8OMFK;=Xe6=Sgf
]V<,;5Q-e5UP^)c^;P-Sg2<9)SY0;:6S-P6A8-:S-08FQfEZJR\-NO,dA5_/<T/2
_<>[;ZI?WXITbe@Y>0U:;279Y/ST>DPf;K0I7#YaWUHTg1[[8bR=TU5H-dZ1(@d?
\@RKb]?)P\A?@O\e@fYd4OHE[+2@>+IJ[6(_=>LHADCXMO^CI9MID+]9\:VE./9)
T-Z-95AD/,B>Vg3.7PRA_NCR0?KA,5V=87QHI@FLTU85GQ0ebPUJ+T&&KVAWg)/Z
C\B9M:D09J;3:VI^@Ba4^HXR/:W]-6,NYO3Bea/)2I&b]^-B6]MPg#&T3VIT_g.:
dd-;V8_).ZU29[(1,4>#C_LeSf(dfdgBR:T=bU]Z-20U=RVKfdg@I;H]NWLFHM]Y
HcH\6KOO32M.GOH;JfFT,V,+5bg/NU9V5FFHe-aY:=C.KCX@#JW,CB=5B04,HW_2
BH<^+?2RM_PKZ5=?9B)a@NYOUBI#FCF9:Tf=\S<Ja,FB)Re,97)WH,:KE0e?>G2P
Aff/#NT?4AWF?XQG\\Mc(^_c-dCT)gAGOZf6SgASKNGC2;O::@IDCd1b5JXX;WN;
+e:XMJB=PHQ&f8C+R^ag,ZCA+#=0IDdDA:6,a9SN-IYNDX^^LYX#V&cSWNaJP3b7
;3UG7-U3BHcI#FY5IOS_(O\>&<gDDG^/+cEH-RdP&AMP;b^c,20+D65d=I,K?eS?
RG9ZU,/I<TbdU5-dJ4GNU&P9BA5]\cY/6RM7RFe7_?8VbX\Q^A=T8RAf&X?F;&:O
/OJ#cgFQgHAEMJX\K8EFePH+0PdPDfB.^MW0(D5_Sb7VE$
`endprotected


`endif
