
`ifndef GUARD_SVT_AXI_CACHE_SV
`define GUARD_SVT_AXI_CACHE_SV

`include "svt_axi_common_defines.svi"

`ifndef DESIGNWARE_INCDIR
  `include "svt_data.sv"
`endif

/** Add some customized logic to copy the actual memory elements */
`define SVT_AXI_CACHE_SHORTHAND_CUST_COPY \
`ifdef SVT_UVM_TECHNOLOGY \
`elsif SVT_OVM_TECHNOLOGY \
`else \
  if (do_what == DO_COPY) begin \
    svt_axi_cache_copy_hook(this.__vmm_rhs); \
  end \
`endif

/** Add some customized logic to compare the actual memory elements */
`define SVT_AXI_CACHE_SHORTHAND_CUST_COMPARE \
`ifdef SVT_UVM_TECHNOLOGY \
`elsif SVT_OVM_TECHNOLOGY \
`else \
  if (do_what == DO_COMPARE) begin \
    if (!svt_axi_cache_compare_hook(this.__vmm_rhs, this.__vmm_image)) begin \
      this.__vmm_status = 0; \
    end \
  end \
`endif

//`define _SVT_AXI_CACHE_DEBUG \
    //`ifdef SVT_AXI_TEMP_CACHE_DEBUG \
        //`svt_amba_debug(cache_name,$sformatf \
    //`endif
// ======================================================================
/**
 * This class is used to model a single cache. 
 *
 * Internally, the cache is modeled with a sparse array of svt_axi_cache_line objects,
 * each of which represents a full cache line.
 */
class svt_axi_cache extends `SVT_DATA_TYPE;

  /**
   * Convenience typedef for address properties
   */
  typedef bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr_t;
  
  /**
   * Convenience typedef for data properties
   */

  typedef bit [7:0] data_t;

  /**
    * Enum to represent the different cache structures
    * DIRECT_MAPPED: An entry corresponding to a main memory address
    * is stored in a cache line with a unique index. For example,
    * consider an 8 KB cache where the cache line size is 16 bytes
    * and there are 512 such lines. Then addresses 0, 8K, 16K, 24K etc
    * are always mapped to index 0 of the cache and so on.
    * FULLY_ASSOCIATIVE: In such a cache structure, a given main
    * memory address can be stored in a cache line with any index. 
    * TWO_WAY_ASSOCIATIVE: An entry corresponding to a main memory
    * address can be stored in any one of two cache line indices.
    * For example, consider an 8 KB cache where the cache line size
    * is 16 bytes and there are 512 such lines. These 512 lines are
    * divided into 256 sets with "2 ways" for each set. So any given
    * main memory address can be stored in only a unique set, but within
    * this set, it can be stored in one of the two ways. 
    * NOTE: Currently only FULLY_ASSOCIATIVE is supported 
    */
  typedef enum {
    FULLY_ASSOCIATIVE   = `SVT_CACHE_FULLY_ASSOCIATIVE,
    DIRECT_MAPPED       = `SVT_CACHE_DIRECT_MAPPED,
    TWO_WAY_ASSOCIATIVE = `SVT_CACHE_TWO_WAY_ASSOCIATIVE
  } cache_structure_enum;

  /** @cond PRIVATE */
  /** 
    * The minimum address in the shared region of memory
    * that the component where this cache resides in will access
    */ 
  addr_t shared_start_addr;

  /** 
    * The maximum address in the shared region of memory
    * that the component where this cache resides in will access
    */ 
  addr_t shared_end_addr;

  /** 
    * The width of each cache line in bits
    */
  int cache_line_size = 32;

  /**
    * The number of cache lines in this cache
    * The cache_line_width*num_cache_lines defaults to a 1 KB cache memory
    */
  int num_cache_lines = 256;


  /**
    * Flag to indicate CHI ICN Full-Slave mode. Set when CHI Interconnect is
    * used in Full-Slave mode.
    * Default value is 0.
    */
  bit is_chi_icn_full_slave = 0;

  /**
   * Indicates whether the cache supports storing poison fields
   */
  local bit poison_enable;

  /**
   * Indicates whether the cache supports storing data_check(parity) fields
   */
  local bit data_check_enable;

  /**
   * Poison granularity: number of data bytes corresponding to a poison bit
   */
  local int num_bytes_per_poison_bit = 8;
  
  /**
    * The structure of the cache
    */
  cache_structure_enum cache_structure = FULLY_ASSOCIATIVE;

  /**
   * Indicates whether the cache supports storing Tag value
   */
  local bit tag_enable;

  /**
   * Indicates whether the cache supports partial cache states: UCE, UDP
   */
  local bit partial_cache_states_enable =0;
  /** @endcond */

/** @cond PRIVATE */


  /**
   * Sparse array of svt_axi_cache_line objects, used to model the physical
   * storage of this cache.
   *
   * The array is to be indexed only by an expression that evaluates to an 
   * address within the bounds of the maximum number of cache lines in the cache.
   */
  local svt_axi_cache_line cache_lines [addr_t];

  /**
    * Array of addresses mapped to each index of the cache.
    * Whenever a cache line is updated, this is also updated to
    * reflect the updated contents and may be used by the various
    * cache access methods depending on the structure of the cache 
    */
  local addr_t addr_mapped_to_indices [int];

  /**
   * Sparse array used to store the number of reservations for 
   * addresses for which cache lines are reserved.
   *
   * The array is to be indexed only by an expression that evaluates to an 
   * address within the bounds of the maximum number of cache lines in the cache.
   */
  //local bit reserved_cache_lines [addr_t];
  local int reserved_cache_lines [addr_t];

  /**
    * Array of addresses mapped to a reserved index of the cache.
    */
  local addr_t addr_mapped_to_reserved_indices [int];

  /** 
    * log_base_2 of cache_line_size used for aligning
    * addresses
    */
  local int log_base_2_cache_line_size = 2;

  /**
    * Semaphore to regulate cache access. Components using this
    * cache model can use this to first get the semaphore before
    * accessing the cache. This is useful when multiple processes
    * are accessing the same cache. 
    */
  semaphore cache_access_sema;
  
  /**
    * PA writer handle which is used to write the cache data inside
    * FSDB. The data will written out only into FSDB and not for XML.
    * This means the handle is instanciated only when FSDB is enabled.
    */
  svt_xml_writer pa_writer;

  /**
    * Transaction UID
    * To support cache operation to transaction relationship 
    */
  string transaction_uid;

  /**
    * Transaction type
    * To support cache operation to transaction relationship 
    */
  string transaction_type = "";

`ifdef SVT_VMM_TECHNOLOGY
  /** Shared log object if user does not pass log object */
  local static vmm_log shared_log = new ( "svt_axi_cache", "class" );
`endif
  
  local int dbg_indx;
  local string cache_name = "";
/** @endcond */

`ifdef SVT_UVM_TECHNOLOGY
  // --------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new instance of this class.
   *
   * When this object is created, the cache is assigned an instance name, 
   * cache line size, number of cache lines, the cache structure and 
   * the minimum and maximum shared address.  
   *
   * @param name Intance name for this memory object
   * 
   * @param suite_name Name of the suite in which the memory is used.
   * 
   * @param cache_line_size The width of each cache line in bits.
   * 
   * @param num_cache_lines The number of cache lines in this cache.
   * 
   * @param cache_structure The structure of this cache.
   * 
   * @param shared_start_addr The minimum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   * 
   * @param shared_end_addr The maximum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   *        
   * @param is_chi_icn_full_slave (Optional) Applicable only in case of CHI
   * ICN Full Slave mode where it is passed as 1. Default value is 0.
   */
  extern function new(string name = "svt_transaction_inst",
                      string suite_name = "",
                      int cache_line_size = 32,
                      int num_cache_lines = 256,
                      cache_structure_enum cache_structure = FULLY_ASSOCIATIVE,
                      addr_t shared_start_addr = 0, 
                      addr_t shared_end_addr = ((1<<`SVT_AXI_MAX_ADDR_WIDTH)-1),
                      bit is_chi_icn_full_slave = 0);
`elsif SVT_OVM_TECHNOLOGY
  // --------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new instance of this class.
   *
   * When this object is created, the cache is assigned an instance name, 
   * cache line size, number of cache lines, the cache structure and 
   * the minimum and maximum shared address.  
   *
   * @param name Intance name for this memory object
   * 
   * @param suite_name Name of the suite in which the memory is used.
   * 
   * @param cache_line_size The width of each cache line in bits.
   * 
   * @param num_cache_lines The number of cache lines in this cache.
   * 
   * @param cache_structure The structure of this cache.
   * 
   * @param shared_start_addr The minimum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   * 
   * @param shared_end_addr The maximum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   *        
   * @param is_chi_icn_full_slave (Optional) Applicable only in case of CHI
   * ICN Full Slave mode where it is passed as 1. Default value is 0.
   */
  extern function new(string name = "svt_transaction_inst",
                      string suite_name = "",
                      int cache_line_size = 32,
                      int num_cache_lines = 256,
                      cache_structure_enum cache_structure = FULLY_ASSOCIATIVE,
                      addr_t shared_start_addr = 0, 
                      addr_t shared_end_addr = ((1<<`SVT_AXI_MAX_ADDR_WIDTH)-1),
                      bit is_chi_icn_full_slave = 0);
`else
  // --------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new instance of this class.
   *
   * When this object is created, the cache is assigned an instance name, 
   * cache line size, number of cache lines, the cache structure and 
   * the minimum and maximum shared address.  
   *
   * @param log The log object.
   *
   * @param suite_name Name of the suite in which the memory is used.
   * 
   * @param cache_line_size The width of each cache line in bits.
   * 
   * @param num_cache_lines The number of cache lines in this cache.
   * 
   * @param cache_structure The structure of this cache.
   * 
   * @param shared_start_addr The minimum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   * 
   * @param shared_end_addr The maximum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   *        
   * @param is_chi_icn_full_slave (Optional) Applicable only in case of CHI
   * ICN Full Slave mode where it is passed as 1. Default value is 0.
   */
`ifndef __SVDOC__
`svt_vmm_data_new(svt_axi_cache)
`endif
   extern function new(vmm_log log = null,
                      string suite_name = "",
                      int cache_line_size = 32,
                      int num_cache_lines = 256,
                      cache_structure_enum cache_structure = FULLY_ASSOCIATIVE,
                      addr_t shared_start_addr = 0, 
                      addr_t shared_end_addr = ((1<<`SVT_AXI_MAX_ADDR_WIDTH)-1),
                      bit is_chi_icn_full_slave = 0);
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
`ifndef __SVDOC__
  `svt_data_member_begin(svt_axi_cache)
    `SVT_AXI_CACHE_SHORTHAND_CUST_COPY
    `SVT_AXI_CACHE_SHORTHAND_CUST_COMPARE
  `svt_data_member_end(svt_axi_cache)
`endif

  // ---------------------------------------------------------------------------
  
  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given index.
   * If the index does not exist this function returns 0, else it returns 1.
   *
   * @param index The index of the cache line to be read.
   *
   * @param addr Assigned with the address stored in the given index. Please
   * note that if the address specified is unaligned to cache line size, an
   * aligned address is computed internally, before doing the operation.
   *
   * @param data Assigned with the data stored in the given index.
   * 
   * @param is_unique Returns 1 if the cache line at the given index is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line at the given index is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line at given index.
   * 
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   *
   * @return If the read is successful, that is, if the given index
   * has an entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_by_index(input int index,
                                            output addr_t addr, 
                                            output bit [7:0] data[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0);

  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given index.
   * If the index does not exist this function returns 0, else it returns 1.
   *
   * @param index The index of the cache line to be read.
   *
   * @param addr Assigned with the address stored in the given index. Please
   * note that if the address specified is unaligned to cache line size, an
   * aligned address is computed internally, before doing the operation.
   *
   * @param data Assigned with the data stored in the given index.
   * 
   * @param dirty_byte_flag Returns dirty flag associated with each byte in the
   * cache line associated with the given address. '1' indicates data byte is dirty
   * '0' indicates data byte id clean
   * 
   * @param is_unique Returns 1 if the cache line at the given index is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line at the given index is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line at given index.
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   * 
   * @return If the read is successful, that is, if the given index
   * has an entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_line_by_index(input int index,
                                            output addr_t addr, 
                                            output bit [7:0] data[],
                                            output bit       dirty_byte_flag[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0);

  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given address.
   * If there is no entry corresponding to this address
   * returns 0, else it returns 1.
   *
   * @param addr The address associated with the cache line that needs
   * needs to be read. Please note that if the address specified is unaligned to
   * cache line size, an aligned address is computed internally, before doing
   * the operation.
   *
   * @param index Assigned with the index of the cache line associated
   * with the given address.
   *
   * @param data Assigned with the data stored in the cache line associated
   * with the given address.
   * 
   * @param is_unique Returns 1 if the cache line for given address is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line for the given address is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line associated with
   * the given address 
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   *
   * @return If the read is successful, that is, if the given address 
   * has an associated entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_by_addr(
                                            input addr_t addr, 
                                            output int index,
                                            output bit [7:0] data[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0 );

  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given address.
   * If there is no entry corresponding to this address
   * returns 0, else it returns 1.
   *
   * @param addr The address associated with the cache line that needs
   * needs to be read. Please note that if the address specified is unaligned to
   * cache line size, an aligned address is computed internally, before doing
   * the operation.
   *
   * @param index Assigned with the index of the cache line associated
   * with the given address.
   *
   * @param data Assigned with the data stored in the cache line associated
   * with the given address.
   * 
   * @param dirty_byte_flag Returns dirty flag associated with each byte in the
   * cache line associated with the given address. '1' indicates data byte is dirty
   * '0' indicates data byte id clean
   * 
   * @param is_unique Returns 1 if the cache line for given address is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line for the given address is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line associated with
   * the given address 
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   * 
   * @return If the read is successful, that is, if the given address 
   * has an associated entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_line_by_addr(
                                            input addr_t addr, 
                                            output int index,
                                            output bit [7:0] data[],
                                            output bit       dirty_byte_flag[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0);
  // ---------------------------------------------------------------------------
  /**
   * Writes cache line information into a cache line.  If the index is a
   * positive value, the addr, data, status and age information is written in
   * the particular index. Any existing information will be overwritten. If the
   * value of index is passed as -1, the data will be written into any available
   * index based on the cache structure. If there is no available index, data is
   * not written and a failed status (0) is returned.
   *
   * @param index The index to which the cache line information needs to be
   * written. The range of index is between 0 to
   * (svt_axi_port_configuration::num_cache_lines - 1).
   * 
   * @param addr The main memory address to which the cache line is to be
   * associated. Please note that if the address specified is unaligned to cache
   * line size, an aligned address is computed internally, before doing the
   * operation. 
   * 
   * @param data The data to be written into this cache line. 
   *
   * @param byteen (Optional) The byte-enables to be applied to this write. A 1 in a
   * given bit position enables the byte in the data corresponding to that bit
   * position.
   * 
   * @param is_unique (Optional) The shared status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param is_clean (Optional) The clean status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param age (Optional) The age to be stored in the cache line. If not passed, the
   * age information is not changed/updated. Typically, current simulation clock
   * cycle can be specified as the age.
   *
   * @param retain_reservation (Optional) ensure that no existing reservation
   * which was made for some other transaction is deleted. The cache keeps
   * track of the number of reservations on each address. If this bit is 0,
   * with each write, the number of reservations on the given address is
   * decremented by 1. If there is only one reservation on this address, this
   * write will result in all reservations being deleted. If this bit is 1, no
   * reservations are decremented or deleted.
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   *
   * @return 1 if the write was successful, or 0 if it was not successful.
   */
   extern virtual function bit write(
                                     int index, 
                                     addr_t addr = 0,
                                     bit [7:0] data[],
                                     bit byteen[],
                                     int is_unique = -1,
                                     int is_clean = -1,
                                     longint age = -1,
                                     bit retain_reservation = 0,
                                     bit record_to_fsdb = 1
                               );
  // ---------------------------------------------------------------------------
  /**
   * This function writes into the cache via backdoor. Backdoor accesses are
   * direct accesses to the cache in the VIP by the user in the testbench. For
   * example, if users want to preload the cache from the testbench, this
   * function must be used. This function does not delete any existing
   * reservation made to this address by some other transaction. Reservations
   * may have been made by the master VIP for transactions to the same address
   * as what  is requested in the backdoor write. Using this function for
   * backdoor writes (as opposed to using the write() function) makes sure that
   * those reservations are not deleted.
   * 
   * If the index is a positive value, the addr, data, status and age information is written in
   * the particular index. Any existing information will be overwritten. If the
   * value of index is passed as -1, the data will be written into any available
   * index based on the cache structure. If there is no available index, data is
   * not written and a failed status (0) is returned.
   *
   * @param index The index to which the cache line information needs to be
   * written. The range of index is between 0 to
   * (svt_axi_port_configuration::num_cache_lines - 1).
   * 
   * @param addr The main memory address to which the cache line is to be
   * associated. Please note that if the address specified is unaligned to cache
   * line size, an aligned address is computed internally, before doing the
   * operation. 
   * 
   * @param data The data to be written into this cache line. 
   *
   * @param byteen (Optional) The byte-enables to be applied to this write. A 1 in a
   * given bit position enables the byte in the data corresponding to that bit
   * position.
   * 
   * @param is_unique (Optional) The shared status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param is_clean (Optional) The clean status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param age (Optional) The age to be stored in the cache line. If not passed, the
   * age information is not changed/updated. Typically, current simulation clock
   * cycle can be specified as the age.
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   *
   * @return 1 if the backdoor write was successful, or 0 if it was not successful.
   */
   extern virtual function bit backdoor_write(
                                     int index, 
                                     addr_t addr = 0,
                                     bit [7:0] data[],
                                     bit byteen[],
                                     int is_unique = -1,
                                     int is_clean = -1,
                                     longint age = -1,
                                     bit record_to_fsdb = 1
                               );
   
  // ---------------------------------------------------------------------------
  /**
   * Gets the index of a cache line corresponding to the given address
   * If there is no corresponding entry returns -1.
   *
   * @param addr The address whose index is required. 
   *
   * @return Returns the index corresponding to the given address. If
   * there is no such entry, returns -1.
   */
  extern virtual function int get_index_for_addr(
                                            input addr_t addr 
                              );
  // ---------------------------------------------------------------------------
  /**
   * Gets the address stored in the cache line at given index. 
   * If there is no corresponding entry returns -1.
   *
   * @param index The index of the cache line
   *
   * @param addr Assigned with the address stored at given index. 
   *
   * @return Returns 1 if there is a cache line at given index, else
   * returns 0. 
   */
  extern virtual function bit get_addr_at_index( input int index, 
                                            output addr_t addr 
                              );
  // ---------------------------------------------------------------------------
  /**
   * Returns the index corresponding to the least recently used cache line 
   * between the given set of indices. The least recently used cache line
   * is the cache line with the least age. 
   * @param low_index The first index at which the operation is to be done
   * @param high_index The last index at which the operation is to be done.
   * @param is_not_reserved Indicates that the entry returned should not be
   * a reserved index.
   * @return Returns the index corresponding to the least recently 
   * used cache line
   */
  extern virtual function int get_least_recently_used(
                                int low_index,
                                int high_index,
                                bit is_not_reserved = 1
                              );
  // ---------------------------------------------------------------------------
  /**
    * Invalidates the cache line entry for a given addr. This method removes the
    * cache line from the cache for the given address.
    *
    * @param addr The address that needs to be invalidated.
    *
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, if
    * there is a corresponding entry. Else, returns 0.
    */
  extern virtual function bit invalidate_addr(
                                addr_t addr,
                                bit record_to_fsdb = 1 
                              );
  // ---------------------------------------------------------------------------
  /**
    * Invalidates the cache line entry at the given index. This method removes the
    * cache line from the cache for the given index.
    *
    * @param index The index that needs to be invalidated.
    *
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, if
    * there is a corresponding entry. Else, returns 0.
    */
  extern virtual function bit invalidate_index(
                                int index,
                                bit record_to_fsdb = 1 
                              );
  // ---------------------------------------------------------------------------
  /**
   * Updates the status of the cache line for the given address.
    * Reserves the given index of the cache for future use. The get_any_index
    * function takes into account the reserved indices as well so that a user
    * is always given an index that is neither currently in use nor reserved
    * for future use. When a cache line is written into an index, the corresponding 
    * index is deleted from the set of reserved indices (if present).
    *
    * @param index The index that needs to be reserved.
    *
    * @return Returns 1 if the operation is successful, else returns 0.
    */
  extern virtual function bit reserve_index(
                                int index,
                                addr_t addr
                              );
  // ---------------------------------------------------------------------------
  /**
    * Gets the reserved index for the given addr.
    * @param addr Address for which the index needs to be found
    * @return Returns the index.
    */
  extern virtual function int get_reserved_index(addr_t addr);
  // ---------------------------------------------------------------------------
  /**
    * Deletes all reservations made in this cache for future updates in cache.
    */
  extern function void delete_reservations();
  // ---------------------------------------------------------------------------
  /**
    * Delete or decrement reserved_cache_lines corresponding to address
    */
  extern function int delete_reservation_for_addr(addr_t addr);
   
  // ---------------------------------------------------------------------------
  /**
   * Updates the status of the cache line for the given address
   *
   * @param addr The address that needs to be updated.
   *
   * @param is_unique The shared status to which the cache line associated
   * with the addres needs to be updated. 
   * A value of 1 indicates that  the corresponding cache line is not shared 
   * with other caches 
   * A value of 0 indicates that  the corresponding cache line is shared 
   * with other caches 
   * A value of -1 indicates that the current status need not be changed.
   * @param is_clean The clean status to which the cache line associated
   * with the addres needs to be updated. 
   * A value of 1 indicates that  the corresponding cache line is updated
   * relative to main memory. 
   * A value of 0 indicates that  the corresponding cache line is not 
   * updated with respect to main memory. 
   * A value of -1 indicates that the current status need not be changed.
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
   extern virtual function bit update_status(
                                addr_t addr, 
                                int is_unique,
                                int is_clean,
                                bit record_to_fsdb = 1
                           );
  // ---------------------------------------------------------------------------
  /**
   * Updates the status of the Tag held in the cache line for the given address
   *
   * @param addr The address that needs to be updated.
   *
   * @param is_invalid This specifies if the Tag is held in the cache line. 
   * A value of 1 indicates that the corresponding cache line should not contain Tags and the Tag state
   * must be considered Invalid
   * A value of 0 indicates that the corresponding cache line contains Tags
   * @param is_clean Specifies the state of the Tag held in the cache line. 
   * A value of 1 indicates that  the Tag is held in clean state. 
   * A value of 0 indicates that  the Tag is held in dirty state. 
   * . 
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
   extern virtual function bit update_tag_status(
                                addr_t addr, 
                                bit is_invalid,
                                bit is_clean,
                                bit record_to_fsdb = 1
                           );
  // ---------------------------------------------------------------------------
  /**
   * Gets the status of the cache line for the given address
   *
   * @param addr The address whose status is required.
   *
   * @param is_unique The shared status of the cache line associated
   * with the address. 
   * A value of 1 indicates that  the corresponding cache line is not shared 
   * with other caches 
   * A value of 0 indicates that  the corresponding cache line is shared 
   * with other caches 
   * @param is_clean The clean status of the cache line associated
   * with the address. 
   * A value of 1 indicates that  the corresponding cache line is updated
   * relative to main memory. 
   * A value of 0 indicates that  the corresponding cache line is not 
   * updated with respect to main memory. 
   *
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
   extern virtual function bit get_status(
                                addr_t addr, 
                                output bit is_unique,
                                output bit is_clean
                           );
  // ---------------------------------------------------------------------------
  /**
   * Updates the age of the cache line associated with the given address
   *
   * @param addr The address that needs to be updated.
   *
   * @param age  The age to which the associated cache line is to be updated.
   *
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
  extern virtual function bit update_age(
                                addr_t addr,
                                longint age
                              );
  // ---------------------------------------------------------------------------
  /**
   * Gets the age of the cache line associated with the given address
   *
   * @param addr The address whose age is required.
   *
   * @param age  Assigned with the age associated with the cache line of the address.
   *
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
  extern virtual function bit get_age(
                                addr_t addr, 
                                output longint age
                              );
  // ---------------------------------------------------------------------------
  /**
    * Sets the protection type of this address.
    * For is_privileged, is_secure and is_instruction arguments, a value of -1 indicates that the existing value
    * should not be modified. Definitions of priveleged, secure and instruction access
    * are as per AXI definitions for access permissions of AxPROT signal.
    * @param addr The address that needs to be updated.
    * @param is_privileged Indicates if the address corresponding to this line is privileged
    * @param is_secure Indicates if the address corresponding to this line is secure
    * @param is_instruction Indicates if the address corresponding to this line is an instruction
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_prot_type( addr_t addr,
                                     int is_privileged = -1,
                                     int is_secure = -1,
                                     int is_instruction = -1,
                                     bit record_to_fsdb = 1 );

  
  // ---------------------------------------------------------------------------
  /**
    * Gets the protection type of this cache line.
    * Definitions of priveleged, secure and instruction access
    * are as per AXI definitions for access permissions of AxPROT signal.
    * @param addr The address whose information needs to be retreived.
    * @param is_privileged Indicates if the address corresponding to this line is privileged
    * @param is_secure Indicates if the address corresponding to this line is secure
    * @param is_instruction Indicates if the address corresponding to this line is an instruction
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_prot_type(addr_t addr,
                                     output bit is_privileged,
                                     output bit is_secure,
                                     output bit is_instruction);

  // ---------------------------------------------------------------------------
  /**
    * Sets the memory attribute of this address 
    * Definition of memory attribute is as per AXI definition of memory attribute for AxCACHE signalling.
    * @param addr The address that needs to be updated.
    * @param cache_type Memory attribute of this cache line
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_cache_type(addr_t addr, 
                                     bit[3:0] cache_type, 
                                     bit record_to_fsdb = 1);
  // --------------------------------------------------------------------
  /**
    * Gets the memory attribute of this cache line.
    * Definition of memory attribute is as per AXI definition of memory attribute for AxCACHE signalling.
    * @param addr The address whose information needs to be retreived.
    * @param cache_type Returns the memory attribute of this cache line
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_cache_type(addr_t addr, output bit[3:0] cache_type);

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
K1LVRDZCn8LJE9mhRq5T3kaAWbh3LMi0h2Xd6P9jLu7rPDAW71gJiIn6MuNFpXSo
pfvggpBMvsxFOv27beWdh4Ycm2MGIFc82DQi7guro69inZXFP1ma6SV3CtrkSSFD
lmksJGXbLfpTBf6JELDGJjpo6Fa924g4jq3m4Y7D4EcfyXSd5O+ZzQ==
//pragma protect end_key_block
//pragma protect digest_block
8bIbfRLRGATGYt/K83Z+MtPKSbg=
//pragma protect end_digest_block
//pragma protect data_block
FmHUj3sy1DLLfGk/Ckgz0Jz4wc7fCi/+dtQETj+P+JGrnzshJkW/iFKuriYs9CiX
02CAsspeZWlYPmqrw/cQiBHlRNqOAzK627rZHushOjyge4vpCJ9/+rfZZ7a8qM8b
de/LwhO0RULvjLyMNT04mtcW46B5sizr0NvjxLhPhZc3Q7q21f5V21XD3S5DBNxx
V+rtBPOBwdf3FJyxPGXQP3hHm379kyQYuZcJzK8cAqI5JuJq0SiSQtfIelAV7+On
K4rYOhiTL9VqZPxczNIOqrF3wRO/yKJScosQ8QJX/SR2kZM2zy2UwX5p5z9Zad0E
cES+ChLWybClwFUOvPZwkEeTFl5ZDODzSsAnzyR3GDN17eYJr4XHmieYFgHPMDeI
u8iCU8SAE9gjC8WlsTXbP6b8tpSUB4XvhRuA1l9LhukZJlpduv99tOC2vbrtHYDE
pxPjvfCFGYUS65qxsDtWx3gykKN5cCNpuzxC1zJCUSmblokMjr+JyJz+h1xE5j+U
Hr31Nds7wHqWfKJcV/q3c1WbBbOKTf6iJwNAVec2pKUTDs45MeYtr1xWLoUHJ179
U/YkHUJ8P+yz7MJ9qwbNfCkjBN/TA46ptx0+ftGNtT0vJQSwDgIOmzLX9ZRu8SDW
0T7ugtxmtHLSNWueunaOQqS2XpATROamdllGj3Fa0dk/2xgp7ifwumZzqD445Ssw
y+0XZIvrIOr5zy/vgiPhtH5XmW6snYrpnT1iPLh/95W647EjcO3O9dkYLuf89+CB
9aL2mCEHWZ2Qebk9YNWIBdiFweO14yozTCS4blt23S5XCmzqzyqBF30xdNrrgSJy
XQaJ4FnwOUnTNs0u3SCiPzU9OzEJ8E+nyrZaXJ2JYkmYfq9/yL26p84Zx3eutKDN
T4AqHkh+aAy6QVBv/7PI2dMbTmp2LjSOoQJfksehwaiiC39BOKzoNlK7APgdjnOm
6+HdVRW42yNxg6BiL/+A6Mmlf8W/a0SdqYqcDO+ZovFJEG8pONpZRLOao7PL4h4T
NXyZlgXb4RtkJcVGCusEsp0cpQ1anW1lvQ0ohVLtj1IaDzWgMXyJixP8pO1801wI
3SVPTgDT1Z4lucMVFJlAou4vDBKn7tCIyQDkgX/SbAlZogVPwteNvi/rq7MR2oW7
KL0MM2mRvFL36RJ0+SALjez4wI90w20gUh+N4FZrMywEW5fPDsiOTy+AhnSl7vBi
fncIU7tjMJMRZmVLdPTvGYrGSylKV5YPvfKaN6Fxa1R8wZa3EJTFmGlAC1EZsDrN
vgUKzh88pKPhetLjXQbPeA==
//pragma protect end_data_block
//pragma protect digest_block
r2wsPZ5B8+rTF+Ghr0vqZIDDWQU=
//pragma protect end_digest_block
//pragma protect end_protected

  // ---------------------------------------------------------------------------
  /**
    * Sets the Tag field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store Tag settings.
    * This method must be called only when the cacheline corresponding to this address exists in the cache.
    * @param addr The address that needs to be updated.
    * @param tag Tag settings corresponding to the address.
    * @param tag_update TagUpdate settings to indicate which entries in the 'tag' array are valid.
    * @param is_invalid Tag State setting, which when set indicates that Tags must be invalidated from the cacheline correpsonding to this address.
    * If is_invalid is set to 1, tag, tag_update and is_clean values passed to the API will be ignored.
    * @param is_clean Tag State setting, which when set to 1 indicates that Tag state must be set to clean, and 
    * when set to 0, indicates that Tag state must be set to dirty. 
    * This setting is applicable only when is_invalid is set to zero.
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing Tags
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_tag( addr_t addr,
                               bit[(`SVT_AXI_NUM_BITS_IN_TAG-1):0] tag[],
                               bit tag_update[],
                               bit is_invalid,
                               bit is_clean,
                               bit record_to_fsdb = 1);
  
  
  // ---------------------------------------------------------------------------
  /**
    * Gets the Tag filed corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store Tag settings.
    * This method must be called only when the cacheline corresponding to this address exists in the cache.
    * @param addr The address whose information needs to be retreived.
    * @param tag Tag setting corresponding to this cacheline.
    * @param tag_update TagUpdate settings to indicate which entries in the 'tag' array are valid.
    * @param is_invalid Tag State setting, which when set indicates that Tags are not present in the cacheline, and the Tag state is Invalid.
    * If is_invalid is set to 1, tag, tag_update and is_clean values returned by the API must be ignored.
    * @param is_clean Tag State setting, which when set to 1 indicates that Tag state is clean, 
    * and when set to 0, indicates that Tag state is dirty. 
    * This setting is applicable only when is_invalid is set to zero.
    * @param tag_str Tag setting corresponding to this cacheline as string.
    * 
    * @return Returns 1 if the operation is successful, that is, storing Tags 
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_tag( addr_t addr,
                               output bit[(`SVT_AXI_NUM_BITS_IN_TAG-1):0] tag[],
                               output bit tag_update[],
                               output bit is_invalid,
                               output bit is_clean,
                               output string tag_str); 


  
  // ---------------------------------------------------------------------------
  /**
    * API to get poison_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_poison_enabled();
  
  // ---------------------------------------------------------------------------
  /**
    * API to get tag_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_tag_enabled();

  // ---------------------------------------------------------------------------
  /**
    * API to get partial_cache_states_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_partial_cache_states_enabled();
  
  // ---------------------------------------------------------------------------
  /**
    * Sets the poison field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store poison settings.
    * @param addr The address that needs to be updated.
    * @param poison poison settings corresponding to the address.
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing poison
   *  is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_poison( addr_t addr,
                                  bit poison[],
                                  bit record_to_fsdb = 1);
  
  // ---------------------------------------------------------------------------
  /**
    * Gets the poison filed corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store poison settings.
    * @param addr The address whose information needs to be retreived.
    * @param poison Poison setting corresponding to this address.
    * @param poison_str Poison setting corresponding to this address as string.
    * 
    *
    * @return Returns 1 if the operation is successful, that is, storing poison 
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_poison( addr_t addr,
                                  output bit poison[],
                                  output string poison_str);

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
dUJFLcbsEuvlW3LXrQs0pHc/Rk3WZMRnH2ggQTYr10vxQlSGbxTL89J6GTXosJPg
6i4PBrEvsZ/1z3pWdxGk6p+B+HkVCD0arFkM49dIahEQtOXAq0P6p8nrmn22R3c7
MWZa+2SOJYFZK4iiVPy0soWzFOSfQmpgHikt14wZr/RAnjStAMoM2Q==
//pragma protect end_key_block
//pragma protect digest_block
bNGzfxuzIUENuw36fEO/obNbigY=
//pragma protect end_digest_block
//pragma protect data_block
v69xU5lHOwJPGOhztFCK6s+I5BVaLMuzd47XtZ9rqczgdQ+QHEUKVVsXGqeHx7BB
0TEfDl1wIyK1mQQ23yy0g2sw5fovX4RoY5iBWhoUK55E4XrfLEPV5jbADEHzVtf5
UG6iCPNXB5f7plPtd5KqbMOueRFb2eM0UmLWL3kieP+yolsY4nbuoBEu+hEJtzPQ
iinUBF80EI7AxzzTJTmo287/jaxVi1h3oojsvDeMVSVii8jasKt/TvpkemljCZbW
VeegxodQhtlRja1ndaSEOhp7fNIGUIaV4li/xZe7IS0M7wiiOzvvr0qMCaDUUpw8
ULSBSj9pb2dLyOJM+SUtorBqENcz+mwvPYVk8SNE5zPqJGcVv65Hl44TX/P9+cPH
ryPipNTwavjI0JR8iYjQdZb2KiFQ+/RTMF/BiwljiKcASQeArIvLIZk9JghVWife
n5Bs/3OyVviIiAj3Ye5dONcl/v6ZFdlCVR7rDa4HxPDLtIHZxeFa52cuskt0DZbD
71RIztWpMQooPwNEQ/nYau9NYpleceHiZpAkJCHJTa9k6uhl47+yfjQrQIB79IhP
wiV0U63xdcmM3ueMOJfMbc/v7zzcnIclCJKHY/Nz3jSm1/lMyHPOUUxSruBLQRHx
IsGb+E0Ea9bI15LiRs7CZJcgJSxeZ7pDhPFxPLWaTUbdLEheFH5AUtMK6y/6j/lV
59X/PbVkL2jeVMuDFm0P6KOsGvEvw1l6mu/SujvHdWbFdgY018pJ95WtHaEZvRGP
A4aVe8SCm1fsec86JY0upA==
//pragma protect end_data_block
//pragma protect digest_block
0O0PQpWzHrA6FZt1Ii26foCVvig=
//pragma protect end_digest_block
//pragma protect end_protected
  
  // ---------------------------------------------------------------------------
  /**
    * API to get data_check_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_data_check_enabled();
  
  // ---------------------------------------------------------------------------
  /**
    * Sets the data_check field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings.
    * @param addr The address that needs to be updated.
    * @param data_check data_check settings corresponding to the address.
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing data_check
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_data_check( addr_t addr,
                                      bit data_check[],
                                      bit record_to_fsdb = 1);

  // ---------------------------------------------------------------------------
  /**
    * Sets the data_check_passed field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings. 
    * @param addr The address that needs to be updated.
    * @param data_check_passed data_check_passed settings corresponding to the address.
    *        For each of the data bytes and corresponding data_check value, 
    *        this field indicates whether the parity check has passed or not.
    * 
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing data_check
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    * 
    */
  extern function bit set_data_check_passed( addr_t addr,
                                             bit data_check_passed[],
                                             bit record_to_fsdb = 1);
  
  // ---------------------------------------------------------------------------
  /**
    * Gets the data_check filed corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings.
    * @param addr The address whose information needs to be retreived.
    * @param data_check Data_check setting corresponding to this address.
    * @param data_check Data_check setting corresponding to this address as string.
    *
    * @return Returns 1 if the operation is successful, that is, storing data_check 
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_data_check( addr_t addr,
                                      output bit data_check[],
                                      output string data_check_str);

  
  // ---------------------------------------------------------------------------
  /**
    * Gets the data_check_passed field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings. 
    * @param addr The address that needs to be updated.
    * @param data_check_passed data_check_passed settings corresponding to the address.
    *        For each of the data bytes and corresponding data_check value, 
    *        this field indicates whether the parity check has passed or not.
    * @param data_check_passed_str data_check_passed settings corresponding to the address as string.   
    * @return Returns 1 if the operation is successful, that is, storing data_check
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    * 
    */
  extern function bit get_data_check_passed( addr_t addr,
                                             output bit data_check_passed[],
                                             output string data_check_passed_str);

  // ---------------------------------------------------------------------------
  /**
   * This method allows the user to get an index in the cache which may either
   * be allocated for a cache line, or not allocated. If user specifies the
   * values of arguments is_unique and is_clean as -1, then an index is returned
   * where no cache line has been allocated. If user specifies the values of
   * arguments is_unique and is_clean as 0 or 1, index is returned where a cache
   * line is allocated, and the cache line state is as specified. The returned
   * index is between values specified by low_index and high_index.
   *
   * @param is_unique The shared status of the cache line which needs to be 
   * retreived.
   * A value of 1 indicates that  the cache line must not be shared 
   * with other caches. 
   * A value of 0 indicates that the cache line could be shared. 
   * A value of -1 indicates that the shared status of the cache line could 
   * be in any state.
   *
   * @param is_clean The clean status of the cache line that needs to be
   * retreived. 
   * A value of 1 indicates that the cache line must be updated
   * relative to main memory. 
   * A value of 0 indicates that the cache line must not be
   * updated with respect to main memory. 
   * A value of -1 indicates that the clean status of the cache line could 
   * be in any state.
   * 
   * @param low_index The first index at which the operation is to be done. 
   *
   * @param high_index The last index at which the operation is to be done. 
   *
   * @return Returns a positive integer if the operation is successful, 
   * that is, a cache line satisfying the requirements is found, 
   * otherwise returns -1.
   */
  extern virtual function int get_any_index(
                                int is_unique,
                                int is_clean,
                                int low_index,
                                int high_index        
                              );
  // ---------------------------------------------------------------------------
  /** @cond PRIVATE */
  /**
    * Loads the cache based on the contents of the file.
    * Each line of the file represents a cache line.
    * Each line should have the following format:
    * <index> <addr> <data> <shared status> <clean status> <age> 
    *
    * @param filename The full path to the file.
    *
    * @return Returns 1 if the cache was successfully loaded, else returns 0.
    */
  extern virtual function bit load_cache(string filename);
  // ---------------------------------------------------------------------------
  /**
    * Dumps the contents of the into a file.
    * Each line of the file represents a cache line.
    * Each line has the following format:
    * <index> <addr> <data> <shared status> <clean status> <age> 
    *
    * @param filename The full path to the file into which the contents of the
    * cache are to be dumped.
    *
    * @return Returns 1 if the cache was successfully saved, else returns 0.
    */
  extern virtual function bit save_cache(string filename);

  /** @endcond */
  // ---------------------------------------------------------------------------
  /** 
   * Get matched tagged address of cache lines with is_unique, is_clean settings
   * @param is_unique is_unique setting that is required to match for the cache lines.
   * - When set to a value >= 1: considered as 1
   * - When set to a value <= -1: considered as don't care
   * .
   * @param is_clean is_clean setting that is required to match for the cache lines
   * - When set to a value >= 1: considered as 1
   * - When set to a value <= -1: considered as don't care
   * .
   * @param matched_tagged_addr queue of tagged addresses with matched is_uquie, is_clean settings
   * @return Returns 1 if there are any cache lines found with matching input arguments
   */
  extern virtual function bit get_tagged_addresses_for_matched_cache_state(input int is_unique,
                                                                           input int is_clean,
                                                                           output    addr_t matched_tagged_addr[$]);
  
  // ---------------------------------------------------------------------------
  /**
   * Clears the contents of the cache.
   */
  extern virtual function void invalidate_all();

  // ---------------------------------------------------------------------------
  /**
   * Returns the class name for the object.
   */
  extern virtual function string get_mcd_class_name();

  // ---------------------------------------------------------------------------
  /**
   * Returns the cacheline stored in the specified address. 
   * If there is no such cacheline a null is returned
   */
  extern virtual function svt_axi_cache_line get_cache_line(addr_t addr);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM display routine to display the memory contents */
  extern virtual function void do_print(uvm_printer printer);

  /** Extend the UVM copy routine to compare the memory contents */
  extern virtual function void do_copy(uvm_object  rhs);

  /** Extend the UVM compare routine to compare the memory contents */
  extern virtual function bit do_compare(uvm_object rhs, uvm_comparer comparer);

`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the OVM display routine to display the memory contents */
  extern virtual function void do_print(ovm_printer printer);

  /** Extend the OVM copy routine to compare the memory contents */
  extern virtual function void do_copy(ovm_object  rhs);

  /** Extend the OVM compare routine to compare the memory contents */
  extern virtual function bit do_compare(ovm_object rhs, ovm_comparer comparer);

`else
  // ---------------------------------------------------------------------------
  /** Override the default VMM allocate implementation */
  extern virtual function vmm_data do_allocate();

  // ---------------------------------------------------------------------------
  /** Enable the VMM compare hook method */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  // ---------------------------------------------------------------------------
  /**
   * Hook called by the VMM shorthand macro after performing the automated 'copy'
   * routine.
   * 
   * @param to Destination class for teh copy operation
   */
  extern function void svt_axi_cache_copy_hook(vmm_data to = null);

  // ---------------------------------------------------------------------------
  /**
   * Hook called by the VMM shorthand macro after performing the automated
   * 'compare' routine.
   *
   * @param to vmm_data object to be compared against.
   * 
   * @param diff String indicating the differences between this and to.
   */
  extern virtual function bit svt_axi_cache_compare_hook(vmm_data to, output string diff);

  // ---------------------------------------------------------------------------
  /**
   * Hook called after the automated display routine finishes.  This is extended by
   * this class to format a display of the memory contents.
   *
   * @param prefix Prefix appended to the display
   */
  extern virtual function string svt_shorthand_psdisplay_hook(string prefix);
`endif

  /** Added to support the svt_shorthand_psdisplay method */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);

  /** Added t support the svt_shorthand_psdisplay_method*/
  extern virtual function svt_pattern allocate_pattern();
 
  /** @cond PRIVATE */
  /** Gets the address aligned to cache line size */
  extern function addr_t get_aligned_addr(addr_t addr);
  /** @endcond */
  
  //----------------------------------------------------------------------------
  /**
   * Sets the 'pa_writer' required for writing the cache data into FSDB.
   * Also this function records the meta data required for cache visualization
   * in Protocol Analyzer. 
   *
   * @param pa_writer handle to 'SVT_XML_WRITER'
   */
   extern function void set_pa_writer(svt_xml_writer pa_writer);

  //----------------------------------------------------------------------------
  /**
   * Sets the transaction uid for cache operation
   * To support cache operation to transaction relationship 
   */
   extern function void set_transaction_uid(string uid);
  
  //----------------------------------------------------------------------------
  /**
   * Sets the transaction type for cache operation
   * To support cache operation to transaction relationship 
   */
   extern function void set_transaction_type(string xact_type);

  //----------------------------------------------------------------------------
   /** Indicates if the cache line is in partial dirty state 
   *  @param addr Input address
   *  @param is_aligned_addr Indicates if the input address passed is already aligned to cache line size 
   */
  extern virtual function bit is_partial_dirty_line(input addr_t addr, input bit is_aligned_addr = 1);

  //--------------------------------------------------------------------------------
   /** Indicates if the cache line is in empty state
    * This API will return a value 1, when the cache line is in UCE state  i.e. both when is_unique and is_clean are set to 1
    * but none of the data bytes are valid.
    * @param addr Input address
    */
  extern function bit is_line_empty(input addr_t addr);
// ======================================================================
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
tKv7KLTQf+a6koTHdoT21xeJdLKqbKJUK+FI/btFlwMCheNSnhifVQ5O7viXynKK
7OkWpVxjhTFRAkoZ4MDNkFCXW+/e/Pyd0G0cZY/7frvJMuRSooTYEzao216b5Wgo
CFRlilhM0kDeOeA9/76ZkhlQrEyutsymtVEH6eF0JlE+ytdOlJKNEg==
//pragma protect end_key_block
//pragma protect digest_block
jLp/Eac0b5ARN3rEgMFksAO6wQA=
//pragma protect end_digest_block
//pragma protect data_block
As7RZNZ0ATvRMTdKYAVaAfNtic0oQCfPHvdBKmexZ4JRi+y9/mP/aq1mcaU8A0uv
9cbKxgK0J1FFVm476TNb9CoLB4hw0+2dI182J74GkYLVP5QiIcMH/gBjVgeGQLNR
TsRj/o8il1c5+ay9XaH0jlJQswOj/M3zP4WrDgx4M0dweQoGW7TF/7D/6lCRzCO6
JvM6RTzyYK+uOni20jBNvHZeeYZ0vyJfXkZcQqOVWk947EUTw5idE2IoTrOKmBqS
yYFskYKEQQDpK9VbNQKAjZ2CsorVEIR0p0m2tMqxVmBY7NU3iFZ2jPzwt1kpYW/c
BvZMBo08Ns391GOYOL4go7A6EKUPpyNpkJg90bMqdyM5hOZlapz1ih5ALj/vSFga
98bUETh7j+Sx+5Ta3KZxBf7Em0FKwpfAgq4G7QeNL8o9nIleokm4Lg2oNIhJGCGz
KrnZfU8/2cV72gHgAhrudr+YLSq7UD3gXc9424IVW/rZYJBR4/YufVHlqrIpZVut
Xd2rx2KInZTTe3Fy/fJOJaHHlns6RkBzUA+OhUUIgH56X6d2Wdj9Wiw6KrMr/s0e
ihhUZSBlSzINGfXhgR24UnJLyvc4/hs0ehH4qNDprMhlHChcYvKaMEXefYBEp/i3
OxoSJXJthwPOo/xFNH1AIubJHm/xqhhGZjrVFT0dNWAaI6ZM6Gr1LBu9aLfXt6XV
tbWkznPrwZoxhODYU9wpHfdg51xXm5hvp4YmW9iCw3ue6JNqT4SWF3Yz+boGcM7t
gud8y9dVb5gA60uR3UKcKs5lFq+Q1LhXAp6yHvzQFi6o/thcaytwF759zLC5Z5Ar
PUAXk/0nPy8lg//LLIHOCzdCLMQwMGw1ywMoX4SO8LJ73I/87+25l84pm7fhkQ6J
qRPVeCups21oyeu8sTe6em4PQgOgNqDeH1udWt2vgFczuLKUcLxCfozlOBWdpxAZ
n7SvOrtc8UQScMEBSAmluuJ0Ng/33564BUFiwvl52dADJuB5u+pnvrUwF9Vd2wOZ
lXU+b5c/Xl1N788enrZNwhBAvdZqtTWfS5mqmACJ9ybQcLkqNKlSLSBW12cgzC1D
jJyH1bB7AtQ+UTY4Iqr11cvUzrfpEQRFtj+TF5M+KR2Ni/KsWiRWBZqrxXfiq4q7
6/uabhMhNS5aoSaS2h5rkBJY52wSLCu1eIZH/0ll7yCLDw4r7h7FliMi9svWl3v1
vLlsglqhFomn16JhHlA1lBFMougK+Ozb1+C0xHWY7k54PbgY0BWehDKU8K/aBooz
pgIeaiH0oPhsRjRDpOG84RJ7nCcoGEkmaj4Cl5hazs48JE9mkQqg7vfyqEKMIILv
6mqI59thO0Pchkm3TNBW1zd5l35H8yohg2fTekOhCXMX1kxxcst3LFT6TyIAs8md
y4kwHDKxvVagXZEuee2I8CGnwu4ucbGakO6AmdZC1flrxTIRjcRoHgVeeoJm1oec
dWc4/tlYz08CKmMtQtVbpCp3L6QKk+xvMioxMS0xC1fIQuNyw3/0794XUss/lu+z
HbfXtRFuNH/xzv+ddpiuDIeRkOdIUWLUP210ugWSQjUg+vGlpQ1z2NWJpxqIyDAR
D/78keaWOc73fxBbdVWjFCdMx6XTwkVJbMeCgXMCpP8dG8W6Vd5V1Q70Mo9kgcNA
enTKTzHTttJguirHUoyRvIiIhj0TB950h7oEVxAeRM7rCUSFkavDsQXE226gVUB3
CasKOpfxSNzAFBwhyqoTysOW2vTkeAUwmSfZDT3m+adD8+jMcq6jt+b5cXBtZHJO
j4iWykISeqtr2I9mFR3/gAr4rWtQVUfYeEm4hX573zhiFMZPtOgf0U/E4iRGqjoe
HjjSzeRXnkFZoCa0jkGBly87M0FBIDuZnioPGtyK/J6e2sJ/IUicKUted1JuR8C4
3g1SUIcHZ2Dtq5b5osD3Tesox0jNIDxzQ5jGkt/kXAyEiLLEnasXlNTUgHd5Hw2F
LLDCLzIJh9klZwbq4XEz6JeDknPZX6R1gtbz29Dhhb5gYsSz5tUuzwN8tZbjaaXo
i0X1Di7xdjVJgfl8L0Jric8mNFfq9UQOo17bXNfsp2SHfRpd9ExN1BN7G2HLCVVN
MypowdAsuDSyDOCQlOnupGlEcQHFHRF1VoMW/plAmCLii8d/SKC52eHQgVl0kK25
TYe5VmiSaoo7bcuPP3sKCgKhyVhdeNi1fz9YNzMtRnuRB0A4TpDB5vq+WIFaHHAA
aE1Kjr1wgGit15MTEDE+WZGBIkIoFrfIwknHz7SlsaNrmJn0AuaX9UvDF3vv0emh
nrP1xAJHuJd3ash1sIpp7iQZ/pnP1xdGJqSUpB1HLIChD9Kzmx82IRwMHuJ7uhF0
kUInqNPY4WkMZh8/CZMVIvfJevDopljPBeNA2dgNUh7yG0zZVb21JGv9Q+2+KJr4
pb5W4u4yKySoeRRbdnHVoSWNGbXJZCrqJb+WhrvYPxQgSl4tHn2UemxxGWqls0W9
ufzClhDxOXSm9goQxXRH4xoe7RHVkqj09tXzHvalwrn5tRfeL2ET32IMuTvAuPwG
3W42OzcOyi7ZqPUzjGUB6lbqaYb2z1HcjpLfiSwQ4mbUzjQ6MOMILwHGwYrRXUAe
1Uz2WM/KHmxusrdRbmvA7Xm9LeGzHgsh3P9uwqMboMU+hae9pLIUifYYPOZZQniY
sIDB4WG1utt8JmOBHRR3NHxAjCXfEE+taeIXmM/5YABKNMqaUYL5XtyigowIzVvu
Bx9IMYsKbP42xXx/2bBF7+zvDrnJvBKqh0sy7Tt3z7zUCKwP6rx2tUvnRvu3EyPS
zXAOgJlSQSplsdrP41jKuhvDlPVaA1wYpXzVkE605rP+1BC75834j6YpnZAv1cpP
TNiw7BrwhSTfNN3v9QdbKA3KKRIOVgwm7rLz9afQW1cPCH4PxZDXpYl4nFGopPw0
8lN3USsaYeAASVeKDFjTZX0SYZfhPtGnTI4bQUHbc4kTZRMRvQ6Pbj67bZ44x64t
SrlEwS/Hq6FWwwPsYTuHseMdTKcH5jZinH2+B3OTKKdW6QnQYQ87BiVwj1HV0IWh
y+IAS4DJ8EPNTDA4GS1P0/C6ed2QG4IApUkeetSTavU0phkM0103cZvBhoIT6eso
o3YEXrTAihGqkd0llQOj93YOwenSaCS8EB06lMRMnr0AbcCleWB5qac32OPmUBOl
racmLF8Qg08JLmO5UjNgvc4HJJDfPXF5T5EB2J2oKDpHUZ6UkSH6Go1AY+RfpTkW
XQ3/R6m91lInPnzCE5rBUNFWIvusUbXvXHHetdQZfQqiwPKH6RWMGLfFjWHhcBJB
kuiRKTpXijweZZfpOSVdc6fny5ZiKErUO9BbOIfHXnW4Ny47B+7gZjihc61Mwxir
YzjWXM6MJ2MH7eaGAaj3QnERgx6dyBlFKbtH6/H915PsYYdkyEJEOwe60wgZl85T
5p3ej9jzsRthchUEuKvS8vaHXEUJGpUAy6kkMySezRSgRyuanr6JE84p4Pj3gRVs
a4L02us4NgXOm7mFIpw7No74P6Sdvgp6RE91NaAJCITSRvNsrv26Of69VQYusAHw
9+OxZEVTZeG2+UbOvY1iFcz9t2D4QrT8Yzstc+35Mx2NvljxmWU1KJVcOYbnVH8w
pt5MLrX8t+W6OVv35hgpRTeOOO1vm7yEbCmf0bv44uMM8Nu4b5T+A7ed5WcjCZl4
uJChHDeucATkvIbnbHnwBqiiBDbNv+arSCLUBnwn4fqQCqqPp5Smsd/MS2YOPzNj
QguhLu4FPfq+typiTgGkV9CxWCeqDBDVfvHpFoWi+onHEeTS0HgTczbx1mmSsEaE
li1Da4F9A4Wrzrh/CYLKLjF4HM7dypz3WKi4q9NigaAE0XziuX45rop5uoeLJG29
+PP7WK+ZYbx2tpO2YQPn9uH90ZCvTgzUkZO91q+RYdgYefF2AtZmp4FS6nHeBlw7
YqyVK5VQOEasbYVyuX6USdcnVEAZk583T7EdFUZ+dLXXpD9mE4BZ2NEoFnX3pD7x
DqjxOK45ztAxAv2rPyxsNJMKFXpQYQC5aVhQpbuVbhV1/rHlu1W3cUZTER79WjEk
jLrz7zYDKRW/ZX61RuaEJdvu2D/iK3UDc9TTB2dlh4mesv83l6SQO/hqQLD18lrm
YEWfal1Ivn0KcMLO+/4WtkUkC8AIEeCz1Lu7NAsOCoA=
//pragma protect end_data_block
//pragma protect digest_block
kysWUoxjVIDz4uzi53rKPkxu/mU=
//pragma protect end_digest_block
//pragma protect end_protected

// ----------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
o1XaS3zqe8k/anuOJLCq0WcFBP2b4dbsRxSxwq3PfFh3h8KLxVj3EFct8XG+H+4c
L9Vxd56HGkCjU1e14cdQo9VLE0S5bIbV9qselxNVHwQsxcr4uZoo1HVAL9db4/9G
XdoI5ZFiUPE7NRs1YN7PE11S4+L1HsFHrG8uA2/Uc9EyG/yR5BjUCw==
//pragma protect end_key_block
//pragma protect digest_block
G/cG2sn0NwA6ZXfsMQTjpw5BGhc=
//pragma protect end_digest_block
//pragma protect data_block
8U6DGD4KnUcinFRk60nSnjA0FexGy60DGlYHte+38LLt/k4Tyhc/i6CzCtATSTDf
RvQB/zGNol2YuS8ZPS8OFfZ+5j2uCLc0KCnEEtzrl6tFHlRH4THbVbmbK43jUhB4
UwyhNeE7ROZdsKiZbZDTtj2ilfBGrOieqSQT5kE4xwONGbZAVgiDOmJ1btf6nHHo
9fwcnQZzfx6/GiLu0bJIrmp4fXolWbSuXByfWKlH3ki1rTiVMv42d6FMFzt9n+lC
TnKjDYl22BSwB1l+autuUHJMO0jKOWI8zE3kSf3la4M2vmlW0PzFzCDJiswSwCmB
C71Zf3eKTVFPjf/WOGxSYOvgugNnorQebycjyteqs2LQDFWnmq1QT40DDuNkaK7W
n6K3ks/Bi42JOOZY5rHmdReMxuaNUl4D94tMyuOr8oz2s8fiNnMb0IGoWBn5cYEZ
UkvmHh2QO6Yd0oU7dqpyA2+kdlmXytQwJYilwFT7kpQ0rPBPD2qZPXRAgDPgzuOO
a/cyF6ox7TngS9j2u3lbMg==
//pragma protect end_data_block
//pragma protect digest_block
LvMpkg9h12DwiAoLlkeey5wDLXA=
//pragma protect end_digest_block
//pragma protect end_protected

`ifdef SVT_UVM_TECHNOLOGY
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
HUA/Pqy57jbA/BlIaHMWKLN9pJbIG67NBNsuIPRijhaQaDYLVYEl17RhNM2YAVub
/QQkejR1BspO8WoXR5CBEtL9/DxLCaESxmzAat2gSnEaP9dYmLeMuezsJnN8r1AS
AsOXcJnbZLiHKcD7MJdu917a2ROU4npNNoEyLhGOYNpiCm2kCEntpw==
//pragma protect end_key_block
//pragma protect digest_block
ans50ARoZfLtxUemNu1o8rVbUw4=
//pragma protect end_digest_block
//pragma protect data_block
Dcd908AIWe7LOi/hFKNSCauTBFZVH4z6MOZrvo8/vxY1QpJahvoxcMQUEIJeAiDG
dKeLU62fvpFGyfPbvjgW5izDdq7mjG4+gC2Eg/VzgvCjSWURbGp8wIkilIR4mWwx
Ia6ajSb8dgdDJrHyGRi/7eVMNgPdZKshld6LRq/4cgbqd+39+Ii0n1TMh1efQMmb
akcdxL4AUmHCBcIwSRzHcJcYYDrqrCZmlYwIoZzCFOh4Du3z0JMJkrz8i5Q4hFta
GDbuWIjCxlmHVgTLTZFbWsub/nbc0XIDdy8VbsguXsNM5WY7swtGMQCnWy/n8YJW
1+DkDYHEL+w2dXVeqLTMKaaFl7gSMXqJYWZafFTIqGZ7rCDTEdbUjJrp/In6X9nD
zsgrVa8X12/8YnMfArpcgTjMMUQECs/fYgCHqvSohoxh429o5Dqc6PA5UcsXhh/r
EONO9RNzsdS0hJxTXLuId/0SAMDEruAkgOWG6DGD8wyat9NByGEbbwZLjujX+QqE
fqWNmL8BMJcF34vxpoTpQUDHhnF+1rxIfftcyNDleeVogqIZ1si18EBdTVi6ZSaE
1hq4QJ+UaPMK4LKaGneKITsJv5gdnF2BVycdL/HYuRYv9ymFOKWvaoXB6WavXMSy
GSPkMevdNFE+86NgH88B4AGPxK2VJFXs4qyTXBCA08AsC//FiyYBZPKxSrgEqrK7
kYUBdSHVa/9A4K0fOJeobduOhFrXxmnZUnjz20ITxAS0jjqqxQDItvGhEb1l5Thj
b3/kVdRN/IriO96uyAVO48CEHQeabIdg6/2Cl3TgjKVGZ9YF+8O5yQ6EqVqKxo77
1j3tevNb/CLlqafGIXT9zPRBfxOiwBZe964NzuWaQeU1zbeQg4fMRtLfD56+rlmL
8HEnwwMWcZPPFc0JOCc/EXPVFPl1lxk3DU7hsDwITSxsR3ZiXXp9bxlhUJnLEBmk
NZxLS4/R/84sr4u8IBpgULnU4dD45EGvHBUo7yBh7/k9HRJU3LNtgwNSFRSmKLCK
BXQTy5KLwuaRR1VDq1RWLxGYvzZF08wNV/NSvxJ7zV8eAd4hAe1qj0nMkooGFj1Z
x4GcnPqh+z/VBh+4Ewbr694KP+89T4PmyyWJ7Wanw+NhIgOa+2XE4y8nuiS98qj4
oiwsaeJEuWBvto+4VLUoLEXq4mUpAYILo8J2zzndycoY5iNYUTHnnAKs5JifHYpZ
XYy0GpuUz7XkrI4IgQ7A7bPK/Onm0PrvBCkwOdzXcZSSy8qzlhvHbYPIIWbn7KhG
tsrlGbvhRuXf3cc3CTk4oe3dRx5jkqxu3458r1iuLTL46TWnsw3WtXqdKsZmgtAu
l776tKzGaBMCS+4CvEYFcQ914SiVGZ7tZAt1wTX8A0hblC0WgBDdL8uQGCLJ9PNZ
RdpcxzkqQKLtNAO/r6ECd7THL4GFXUbGdD69aj9uz0WodorBc+SQY76TD0zmRpp/
Fd9eAj8DpJ1zO0GT7FkoiiHJgBEC6FYVMDFqmxl7FpWdXTi21lQ1xYf408sljbjq
vk5m4uNspHY9JBBn5X+GTMSoh7V7bN7b6ogd7qlJ0Vg7KG42z/1Rw5L2gMspcJ7F
BW7bSFmbF6499oZ2jXicEbmDnZ+a4jFmpk6mU8dJaK3kAiwuNK9Dco9+WcHKJMMa
K5uwL1tnKn0yjBl1YxfshWdOU5qYZ/zuukT/fQiYOKyNYUAhrvQOLL8XMWrEnT9V
fCqruFBpN3OyXIJLRoPZUHjl1ekrU63L7cyYo9qoNE3tyLGZjk+jfvC/Qmy8UfKi
l3HxBDuXOiG1RKyuxwO/FoGLVP7UZ3VJlykuhZdJOzoSSx5F4LlqNqET08YpBoNU
bztLF18MGSqM9Bjpfp7j1VaEKhhPgeLuGyiFdeRegtDPA93ZVaFUPgWiJNFvqOGy
i42L9SJi27OUXhvRkbmHW8Chk/wK8dTdJtPP9KyCTojg2/pid+t3OHvmft7V2XCj
vjXJTmQ2rpv5Hj//765x6fM8vXG8DZYC0m0jE99dgvX6ZXZD/qvCUKng2YfgNFPe
fWMGj1l6vxX62pSsWbWZbXKAoKRumrbCVQtCNb6k0AOFK2GT4RtVDpYJQWfcwEYj
vwoadSszXPfrGAZxt9WDdzDIZcrshlgBFsfvVGBfSCQB6bfsn57mR3+JB0NM+2zp
vWPTd5gq1NgHbr+wPIOLYizSfpvb1JWJLeiigDEdeIA95vGbKKRWEW2QgFIHh5GW
O5bIIohWGT4G1m0v33XZARb+L5xH1Jhfm7JdxTU625m923Wf7vlJdCXiqHALWA6j
dJcqkbbqOt/4F0bJ+C9HgNNnvYKdiTn3D3C/9W9jtBgPbkQWg3X1RhBpk9N4wbS3
yilxwKcwRFJ77nbwsUWazPtmGAriTkhCbG3zIhu5vzq35jTHaWgUv1hECurw0VmO
AoSmwsMQRPWB6MT8O3LWy+xxku8DEd/sgNZp1WfYWZbvuYy7/js3UiJ4UiL1ZiwK
+gcf5fWzLCV3VWI4KSqSPw5nhJssWesTT5b4wc+kmg0w/pV1s1ydvki7DH4bVDzQ
xapDfebiEhjCNHkIEOgITiSxOVJk0kB2AWkvCj+xz4sH0GMmhcegIi2JVuo/ZXzw
phTE6trOSexTdTAvzaNUQDxV351PhDcFBjMZeqoaRxUeIG3kqcmPFvLIPyx3Uuwd
CwNlKfBiM4gzvrMVT4LCQRRO52u9OFROQuRna1vZwjHerY/zT3NP/aiXDru91vS9
Yvc7kVizIz4JkHwMWMolV9pKVHGnO/2ITbKCZycZplIeJwMGaw3eMgOLX5dJnbjh
uK+MFN7X8r6Mq78marahjwBr1o8R1ROVoo1DPBu9Src1E1IwBQ+LWQ+pw79Zcpfg
4UOEMQOJfS5LE74qAqX4CDLKJnbUWkV3Q9tdCu/nfBzwiuXPYwK65Lelm7LZfWER
um+Knm+2I3yE0Gxoyi9weCTLSRgJi5Be/Q9pwCRLLoLcPm+YiTMOGYm4UNfVD7IN
kqMTqhl8NPPk8yRTW0w5tA4Pxus5hTgSHb9tq2X5h/jiSDzTRLRqEB0CapcNtOlD
mdv/Hg16U7DNfES5dDLwQ6sF66mXZ+YERoV66kgwaWqfQ9TnTpr0ouiomCZ8/8R9
0PovB36kUZOJhUuzgMoDkR7/gjEiTXACeFYW9EZ+xu8=
//pragma protect end_data_block
//pragma protect digest_block
m3x33iieTbt2QKfgz5KdE3xrS3E=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8ECCcltaRL7FvXyamKuguJX5Yy9p9/mjXuALrcbLagcqS6Vtr2GmAzkAZtluRXt0
UxRks1cEXdSUaKNurga+CwKmzZrL9MMZqEQwNFr9GMk8/Ky1HewysrkxobgRf1D4
sxJ9i5quShdoPzgxbKR3UfmTdQbPlzepe4Jk3V9uXmJWhztGC4Fk7Q==
//pragma protect end_key_block
//pragma protect digest_block
4SgX4GPk5a4O/Ix7C94v/qJiIqM=
//pragma protect end_digest_block
//pragma protect data_block
xuE1ViOcYPG4Ds61TggCRbADmej6uSylVLNi188zPGq37pL0RFusadth3C22/TYo
y5/6hnaDU45dRBhBJwwKA2rBHaZFYHy70xsLuFK/+X1Lvm3ioskATNERuXERHx5U
46wE8mY4/ms2LxXmlxrmPX//S8DX8qmAMtxpu5XYJVrKoFqJ23ONAduTExq7Q7iL
9MzxSZa6+0XSQzcgBoqwCmWL4rKKPXlhsmKPrG+az7obpOC376dnKeXA4TtEVGw3
+39yOm5FdFsWGeiNK6Ml1/q7yG0PN0o+xhqKhjvY4w7YXo1CiWpADk7FfuMUWuQi
22lFFwnBc3XWhim4/x2d21XZ87A8Rnq4z7ijzcKiAXqBqxJDRZD01v638fDygY83
Htw7GyDz9v+qmEAlPUaFwsBuwuTxSPBmSB7Pq8/4KHhbO7a2yxS7AO0hcQRYPF2w
mhQu9RJvKz4ukM7rebTEoBCdHBvV2RrgXuRLEZjuAdWBzCzcUVBwqapV2ycuxI9J

//pragma protect end_data_block
//pragma protect digest_block
qM4tpuz7dv+mR4U7Z8siFUbKG0c=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
gSPSJjOAhQoDNai4fw2umiJnOi5J9EWOXuEjMmzLTCIKR+iqy47hFz8IATs/prqm
ntYch8QqQXNS98qQJJ0Mi6fKzBhTsythrDndMlHoonyZF8RKu+U7jDGsrfPuxASA
5P6yM5HPizSKAmHgq33ei6O/RxPASV4hxy1f4ckpXV7uDXfS6y7vsA==
//pragma protect end_key_block
//pragma protect digest_block
fETUpkDvz6G8LeTQxayC80+cp1M=
//pragma protect end_digest_block
//pragma protect data_block
Gmq+AvYgneoWDVVqDEUNX/Mo3QdxlsbmXpnnBjCPN7tuIiWMJaSIaa9VSEc2U0uD
UfE2SvUBLVpfoaIViChOGjMzEeA0QNqtYRjHM5rHUuV6O05A4qFRNu1bSwZwxQMG
uvYceUFZSAC72HXbrNYU/GeoIcnYahudNwGq/4Uk0xUE2z91lyIS4l7+TzZOaVoz
WkFcu7rG3HUf6KeiC4OfYSv5L/zu640oZwypmhkLhFNK8Ks5CnN/yCmZmIDQ5JAq
nHFAQdyJ1JBc0YybTSvUwaXVF9ruTkWLHBen9aT3yK6tpCc9IBvPzhVRpGfDUJlh
xWsJT2U+lGAhD1OWslJbiIC9RvA6EYuQ0XKXIAHBAGB2QQvz/7oB7WODdzr1O/Ro
FgK/p0AKmBdUfKRBGy84BuPvt9IfZGcb/+by8pqSZArZnEez0oBsOliWrnEtKBcE
4mJPZVnOsaBSR5GdbIfVsvm/y6drzhkDtsLCXKm2V/TRTMur1+QK8umGrhA8IUI8
MkYPD9k07zJvc6Jdl4bvIoGKXP47T4zlKhqwTkgrR6Qk794HnEMKW0c4I+9EvuuJ
EQo2055eXzrdtPqGm+L9/uUmzQ4hIda+Rz4la/UtRbDckLvGaTA7ABqyu5EHdCx9
7/DxaaRrNs2uOaebQ8VwOByjv6Mci6129+4khrEaxqFsfsym9GE5pQC5MJBEzE7c
eUtD1lkszGbPR6RHbBAPnTV1kt+ex3DoFqUQjImoeXazugLUbpVXBzS5LJoGAAEE
Ai1ZrOcgR12K9R86dWqga0Zxt1tHD7JpEHvkHGnMUkbCfgWV+pqm7/vBFdrpR2eK
oYvfRxsQ9eEIMwcR5Tn6wRjNgpfrmkN68nUEWs0WOLPjj33Q59eJ9jLlCnnoE7hs

//pragma protect end_data_block
//pragma protect digest_block
5in+s6cBuMxE/9o8BnOSE4JJ2qE=
//pragma protect end_digest_block
//pragma protect end_protected

`elsif SVT_OVM_TECHNOLOGY
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
CY3a7vU/eTTIQzjm9223YUEwbhc8N4NSUFjesaW9r3cBoS8wrTD89LhO4vYAGDTK
mIuJPQ4tGtGwUYVQg67OV3ZgXbnHGLYhISi1/4F/dz9tLbA6AviLKp1rdX3baDqr
b5YMFpZtBslFbEoSQpRMXKXWaCnSDjnBjKNkeaatWcYahCv+c6tbwA==
//pragma protect end_key_block
//pragma protect digest_block
E1Y0cPmB4t6BXJ5D1wuGkiGxkp0=
//pragma protect end_digest_block
//pragma protect data_block
H2P93b+SHhH3UZ53ELRBI4EZNrXPGbajXedrUWCoJztdTmC6O2Nv4qmGS4emNAAY
5XYr4tg1YFRzMIcbIrAWpVTHEcCCjUdxe5hBiVzqdOIvkoAYnmYjob61PauvhU/Z
gXaiAAr9mTI62VVdKLxr9ACUFJwTqW0aDxvbly+JpZbuGOzgmh9UAR3hj0TkDtmC
Oeh+hzo2xiObhSbyGv6Kb/zKVfvm/vI/duz984NlkjDivhNMaHtjK8o/r7Zgnljb
a/jIp9hm9PJ3Zz2gZC8XIu+/9znA8zPEjMFiGxER3x6Mj0OQZxHmQnwngoRK10Zj
a/Sw9thdB1n/wGZdYNgIv/0IvWtUYVJlBkKOSsdKyS5sfEvSm8eWpj3+SlcRVbof
8A6BcN3CnCza/qPeFBOBEDy3pQOguIzoZRFZsejSykb835H4zpwAfI8Npmbr92Pu
0ErT4m20GYFEu6PjplcfaUmdSrYQ+ps8pUWZF0vMdp6jjIw1BpvqS993tO29UFNh
uMkKr6iNy9EY+pbMLlnajavOyVbgv54mtBzUj+COPlFlm+S+KFjLkwXH9V1wL89D
/DB/ZULUV8QQ1v9hQzZyMWDPdsNawCCkU2fGilrBojczWhK+G6rqNHFRkKqUgcT9
saJ3E+fSvBYtlFTV11/wzqwv+EBi2x0eWmBVZ2wdVVcTjo7YJa4r3MN+XmPaUnXl
4qsZpxG0IezIi7fBIAxNZbjojAJFjh+St/d0L/li9ToUikj1A5q8UQ7+vQtGbMWf
rZY0JMwMY3LxkJ+lYQpSO3Zs468CUEiJRvqVbdSgOzYsmYc1rK+KGbEUoMk3xKJD
OdCZ1NrbwfFtcuLXuIApPbR0jo1PwfDGpD/68BOQBd8ZrK8gEQQBl57wX6S5hUir
t4Rznh6oMiDbhVJYLnMY1kd95s61jrRQJwS88xaG7sZDz9RoUeYQM83YioRNHb3R
7vlf/COy81JvdUpZ8o/L9LyqMZ2wR3kR2D9k4iqPvW68miZVyp1Nywvpv0p3k23B
vqn49lQG9MEw1glpgM/eRBc2TJInqDt09BaTl4/iVaNH83LZ/NyuOjLLB4X+0ieI
VkR3kUzpyq78Clrq62jq27h4JX1bVdrMxnuyK7SUN8CSmjx05vM8vslm/vGtkIKD
t0QnPuybcdLi21cFQGPqPlFWGe/GQNqpsfjqB+SqX6PtjdG0ZdLG0h3p6eOxAI7H
7s6jXFID+c3ucpylmUpfS4J474aiKAsVX8kiVNLb3a6TLmzMs7OwNLyn8NaKI2Oo
CCMRwnZokQQAZVvZHKCr4mo12MXp2dQS0Vk1QTt5KNnm66GsCkThXnxXS2xKJxcL
URnCc1oURRAcxu5T3Wr7YqQwA1wGSAZAmiiTGiYDNpJdKh8sIbdB33duknONB4SW
719OOrHxrU06k8LlI60bRqD8IXpX+qUjY3yifzxcY/gYe23wTQPNYYYMlu3Rt6Kx
UHz6lXOt0J/fRLREeGEKMgzILb69MbOnOPMDzn5lnJ+zjlQr0vkECeTMAoyiFQsJ
Nlh1ITC9cgD6Yx+ZOGlQX3wRzw9P9Fe67qaZZn/21j+hfkLphEsbf3Eydor9QB/P
v/cNN1SxRELrfOUwjEuiuy4nforin0l1/8zQlDwpBmXrad+MkHKXh7TWo1ZCTglY
/F4idLq6KgG4xYbxB5RkgPQQrU22b6RsDWiUQ6jNkOONDwiKf6gRDRfoPOTFBG4J
ERShF2HTxBGppwCOY5utXEzx+8gz8k+UcowbHp3enDssFfVo3xSJ9MEBApr+hoEi
V7ZtDUcmuHe0RzdxaZqFDZ/bfFmvCghg83q4JdHE3PSnqEU2CCY5Q0G0ejQA1Ecg
lacVShnyh6Tdyh5kMyydaLNSro0zTOmBv1ro4vIuU6+ziNAfz1o3wbWkJn0bkd+M
SuqTWUAYHGOjmVphx50vosJzWtjAPHdziLPILdkPVXu2GMA2bjl+TYKkr4b4OOml
FpvJUGlHdMCEZqflMdQZ+0dKLMpnNmM/pqFNAfZe3+CMywz2nyL4ayCR5nzWo0Td
PSLYHiiq08dMK87LSyswtlH5qUoqWD2hNLBAjBI4HUX2WYUFUKfLZWFdEwTZptwj
Nh4uuLU528StDvMXrfYqjkTgJKbBLWG59SWdvAvlLbCN0sMJ89QD1lDcrNlX3LVY
z9r3IgoW410ZiSVtkGYi9nNbwJeDm3OUYGXfWv3lWvW6aEUC/tpVYoV2yAaF/lOk
wodOp9f7kJjXJ0DLK+ffTgbD6q+8QsYBXuOIN2mkFQVmKAWFqYtSOjHdDViWMbIz
B1OYlK7xaUbbaSyIBiJ7M0/WrM6lcDxRcI/isfusUAlE9Rmpvb8Anh/clxJUyswV
7g2/GVauOBI8XrXumsz/2OxoIpDLnHhI/eAz/xltOSmsddL2vI+RlzXhvKaGle+4
tofJCXtBlK60l9hEoCLOPQOwP20keSHZrMmSkIEc4Fx3BQ6kO/f+5b5DJDBIxUzo
5udyRImsr/F1PAuO2mrs4sA8NVf9OTqWCGQgXeptxKRHRDk7GahiVY+4ABAUhz6k
aY6Cj4hxAcJp1yVfBRr/BhR4tF6hWSXRSdstYhI9gRPbZUEdeIVDvx5Fmp2Er6di
KN7BeIzHiMnOKV16jaOx2VAnQ05W5vmphuVJ56ZmNTMIiqZB/7NeIHvaiolw/vN9
E+to7+RZ52YA0XVenMkl1y4DyxYP6RvKh3dLf/w9BQfDCcJWvqkIPvE9DmqAVlSW
WJpsUtLiugsZSDeA6j4PdXMeIjo8UovGcVqD+VjacGOvxHyiAMwB9T8GpnjOt3d5
FXTI3RDXZCX4mlJOlBIHhoOeEP6JGcicxpLBq/G5lunbyiodaR5S0ldGJqAUnu7C
qmW7BUR93DLPMy8MxOQnIFTqv8cAJjZCoDYQCatLYVqgiZ90NE6Pd3bXqN4M3YNz
ixbzD0Vuv1bgnWzoqRShqJXLdFkL+4vfwZhM0dYpi6DU/wTeoPim63X5xr0gadUt
h2mp17UGKp88HZryMoWVQB6/gVvxdVWOZdvbPkGtZsfb8ioA0eryzRu+EdhX7+cm
jBXzJY0dIPA11r2M/Futj2Yrn7zOf4V5hm8i9cK00GaFaFf6VY/yz0YgK1LOPehI
7FYpacUxnirRUKf/MMJ7encth/qI8iQQVv/s9JlzBPHRHDbEV9jQmnZprQeIIuOD
NJThcAYz0G7oW8YlbVrG0WrLGXs4vBzyrh+Hr1EGKXhWpmd5+0R4mQ38kVI1nvUS
EZ6+o+pkd9hsLooB/g/1PzBmJW45wssseB4XXmZ3uR7CSQMOgE8JQGkhVvdlE/g6
X2qja7kwdr3nj+W0UQZBQ76TVlOXMEJTBfR6mJ7he2OOykmf3NP69jxzBVR9whOv
+90AlbVjIBxDTbupSy9TrlFuu9ncYWVu7nAv33dAdWj84HzGJWgstyv0WJlwyMQy
IEdcOTGk2oSROwgHotbvcrhIASsRJqDCZPSbxgCz8jdqMNOAmNrdRwwJAHw7H/0D
p6r/1fETQ0zqr9hZNnYqPcxWT3qxC8d/f915HylhXyJwLm4XWO8yqSzy0KCjGECo
rfUd+Z3pS8DgA9q2xtSS9mOA/l474mkZHmDaE6NcYCV0sDy9z+sylxxecPuX+x8x
019Url3q/eys9DbahKkDqZga4b3yOKao+dKt6giq0AvM9Z0CgOPYjOPA+yZFITEb
4oQ9YQaIFPY3G5iAQbAFRg==
//pragma protect end_data_block
//pragma protect digest_block
pdkggpLM4j14ULNvfiPc+1PWPpI=
//pragma protect end_digest_block
//pragma protect end_protected

`else
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/nB0G/O+MgVO6QSMsBG+MInwrvHoOT/nQQ1t28QGFVJmCico/t5Ws/vJMDxEmWIy
kwp5Vy2SilJl56Tbem7L2FAcZ3Vntg50hlA5du0xYCyjW671jf/F7rePva24S739
35tts30S5uVaIXahx5NL4xJqZMumWogbiJZ92dUp6dkFzGGnYsNqxQ==
//pragma protect end_key_block
//pragma protect digest_block
mfFeL0sgCNbej7dpOmf651DKyBY=
//pragma protect end_digest_block
//pragma protect data_block
ziAh4yXqAx6tu3MnRRln2Av5nFnZlplhZQ0qjhltvvroIB6Ro11v/3dxtAw2B8IE
tVDnHd40rCFOOJ8aWf4SjXSByfPKC9UetuqYPaY6dnNLkML4KEK9xCbRnN2riRFX
XrP4Jn6O7WWUygKUYQlSpQ/Gt2V3ej+qEkw9H228DTNSL9Vqnw+z3MckcH8Jxvs/
o4CINVdzND/1Lk2XD1jW/SALgerfREUxPDDDeR8c1IEUuYxgcZKDS30zDJOoDTpe
T5g/ZX+P4OH9YDOXMWCOgkQV/E3FaPl5tdMYAvKbfh18i0S8i7xJvGDEebbFTG5s
Alo2HBKA9rID5x34D2a21nuPg/9qKWPO/HwoXTtn/sOdnTVxGpArh0ydBHn08uLx
RjuiMnLDOlvgz1tdlTJoc/Ir3e5bIGa3fT0Y7xYXhgnV4xl0t2sYOjkJvQRZ+cOI
Y+ozL9tgZzLOvCKVgQjL3zqMGHq0rX6XBc49tUE/6mwhkaRsdTmf0nL/vFN6SrN7
xjtod3KxQezk/JLRCOUoV48KEypBudN5geC6nCDnADC7xx/XPUBAo5E/hSaUe+MB
pVyrDgAE2SrN49/4w30hN5SkjPmtPI1VVClTs1pXfbRBF+S+IvNpwz+JLKjfDgVs
XQpkVMRoRIr6+mxZdyKIsL2i7DqOiQz3IXSZrIabDBDQ6DMhIFMM9SX2gSNUn5Az
P6tXZoXSBg+LO+y3NLWRjZg8Fz5yS7RPTLTxKCDbhNSw3AC6lJs0nxLveej+4TJt
ARft49gB8+N4VRUfZ0eoPJY0BcF+bS0kKElzxuPe87oGKIHyX7K7E8EvT8LqnicK
JVsKpRhzDPQLgP3BGyiFqtxsavqalhEH1IU1pkAp6pRcajPlWyAGG3I/3aWW/tjb
62IJOWpYbdn3TERTux1Y8jTir2AKi2kqKJx3QuDfID44QxgZxxvI/GUMsPFD/SAz
0WLqDmnFE00o77Oom9PkGfu5PMRwUP/6hYotpbYk/XTb1oVb0hwHC0Fvcr46xInl
VeP208O0/4yjEaIow5w7mGDaCHLRTPFtFm92Jw/f0eKqs2RnXAjNsPhiiu916Wce
QZzTdrNGvbQHwTowqV2dIe+0l8E9BnragmYpDwFLVW7ATxhHBOeMAyr27TcaPRFZ
9XeTvLTC6g3qiX9gKWZXfuip8MrRyfbo/hEVFVVilsIN9xfA9S4iSoSUoOdHxDxN
98oXuAD+pCKyQlPVuCHn6+EwVyxQyIep2eXHaHeRaVB+NVJn+/yDmOuWLOlWWGUM
tAOGVAK21vxx088bEoE5eL8EmpOWFhjvlb3gAVKVEKbqlRG+N0sTCTIhRsd4mSTV
XvrST8SHEQ6obmvtB9rKsrT4RoII31M9eDcpABUlRdMdnk4+4T9l1AJ7X7VnvSG+
lfafviBg27jcawg72ouvjJT0SJP/yy4WLlhaNE7GwnSwxHbI/wDqw/N9daj6xDs0
0v0GT4zGV4lQf8fEPCqJpoyAdG6YkeKpuQiwBi3qs3J/xmNy4Dfx1HZmYlEgbsfX
LdKADYzxvoqwlyD1MvhfAqm+kqR4MHhkUesXmVc0r0dQBCzvR/wfNNaoNc8KD+kz
DywfRhHkTkg6tbV1qApb0VbWUocrb0uFtse+zN3DFFc6cJNC06XzKb+PPtQtEuBW
a69UPEk0mI8UkcWWxgqYDy9sf54ohsrm1TVq/JZecOXzofeTu5KpXVYn+aPLQswB
XqT9o82F/FbI+UWJnoW61IIAH0oWW7oPEmv9Zs5cljOBT71zDleWKwS+xk6F6Acp
ZrDtlSXVnXX2FibuvwhPaxjZ9MywCnSv7Oi+J+0b+a2SbQcfy2QycUXPh5S2hQQP
KEkwn3O8nu7pZM3JO6H1GS70owwr81SJpp07YhhiQIg5wLOLNyOeY2uw4HOdHZ4p
8T0U/VGjRWV+BRJb/Bd1lYhhUu0NzPj7NG27h6F3anYI0xytC4a5qbWNaI7MLg82
6JfqfLFWWP56/O7YSTRXlfa2zzGpmJ17bNfXlNcO5g55mdw0blmG102uq2Ri4/hw
ccych7viqhmfTjESHplr0VAXgwvqa9+MYf7j6/aDhBYMJk2pNFUi2ZWHrDx8r4eD
aJ3UQzDmHdN7vmVQW6NhBsgFl68CmSwxEFhYSdptr6mrmoLePWAQx14lgKOJhLNr
9rxMmc1ExeLcVm+kaG9hUFlC2/en2uSaF9f0NnCWrY6u+zgEhFH/OWxyBzPCJohM
BDwJf/Qbeau7bLNH09YgZD+egqQ7DQWf8pv6PK8CeHS74Re5EhhTKwD0oQ/9azh/
djd4aui0kofAfBh9nawjGwVxiTe3vGODEstBbmEDue/wCR4nKSQhDzw3XglFzSZG
hsmrcftZeb6eRpSXCEct39kMC++30li4RRK+iU47B+gs4mGAi6unot/WuTk7fTyG
RVDZOJ/nqjrKF3DbH1Z7Aifcfeu2DsW0sJ7QPawMOtEWXAYXzGKC81qCyTw4Fvda
8buTAJp9cFvkvtjWSRbxLeLU1dVh7gaGI6egfpuaHBKJYcMWcgEtThNlgu1Nuj7c
xF9W/9Xle8iQVmSc8Pv1xcS//o/5Cfe0Xrj4kL1AdqeZBtd4/dKz4nA3/ezon6Dz
rxGdRZT2MbGeSfly+iemgPI9HQ+lQHwIkTyVY9hOYQjhd+VjixXjiLTi3Lz8iVme
6CvsYcAoQP+gQysz6AWXVRYm35fgnK7nXFYByJN+AYBk9MKSJ8V36qbtpEN94W5Y
mOroBGNX9BiRUeBFT4S0xFacxhnKYt/gi81BtX5vCMfD0AHfUpTF8JU0MpdOuUDh
oMzyeOYEY40z+egvrmZ94GVZfZ4G2WYI2330boS2Ly0XmiKUVEFo2OjJtdoRbUDA
80IhLQ5Wt4XEYE0+GzQuJcbh0YDJDMyI529z2W6AXfEchsNr4eNuraBNL9d0fYAG
/xcN0OIJ6zh/d7B9KqAl8o7Uw6cm2TvhOVNfJlLS2A66sBK3LoCjwFTqAJV2ukYy
RIGptn31j1Wjarfs//zRFNDpH9UylpOriqh+68MkJU6RGm3UCrJvY6LYzFPW747C
Lyg/oobc18VISAI0WX/SG2ac2KpuIInmt6GX66lIizh3jCrpyu52aXUaZNh0OVEO
9JPbQJ5feUq7bqsLzFQW/USoio0E2TKJjV5y+NytlXTaJdUdHKbm9tacvrGDoVd8
9viFZB/cQISkGw+4RNTq/FzOpWuj/GHg7QBdJcrYm1nbBy5/NOZsq9FUaQAHPWYx
b4edT7CCcqbOXoOANVDwC6UkEr0dAkLKac56jeEItnyr7/GUXMS2mjo4SeKRAKs3
Osxa4m6Q/fz+dWJBcwYFF9CYe0rd7pcLY9sBGbrEI0HKwnIOHSe7K8ZuUI/FqGF3
z8otVTbgjpMvNW60ZhxulxE5WVOLTGqO+Ex/5iSBZUvljWviKszNdKQA63nAM1Bv
bXsRFsOQJBcHsa+PL/9gtvF2A3AY7irWRGMd+RddR33yOSArSsFibCo+Heg4k8HL
Qp/K50bDyh+zF9VdwuL0R+KFFlBBY4vYzLRv0+aR6T8JQ2ha5mvEczFEstqEk7Qw
sqAdwtA6QjWj+kjms0R+4O3KJLW9kY8BHzaH8nmeSWoOQd6xv3xEUEBnYNW6T+FM
BirywBwq6DaKS33GWZiV1kmIugI/B4GY1GqR9UPNJZLQ9DpvDzTuPhmD/Lw6QXoC
qV+sUrBxnRKMWMtZXw//o7roOg0wifW1hPx1o5xYIQ8UxwMhXVg2q1pTw1aErri2
67QsG17FPVNx3gdM+/jPwZMGQcAuixJHHZyFnEXwiN/DmJ8sz2KeNlf9RDw11DPH
36AzuWEI/nn1Kc1+3Jk2itlMuKjNvlYxuoqwmGmLkwx6o41pyyUY9fJBVPBvjTpV
3l//E39Dt4WqqyIep3LB1AebOy1emAy+VevO1MEst3OrUOe4ZAjhjXxg3/mFkIi0
/edCvKZp9fsYbJwrEAgO1pjpGUYYtToDtZ+vjWu1cc9GPJoh3L7+o23wdLs36L0U
bhMitBeAsw+6rHBJGrB75Unv1box12xtadY4w17LgzNT3h0SAKiBWbHSlBDTFLID
EhQWWdbG4i5Jmh6gHgG5F28riEWmq8wi+JNVD7+gRuSNkTvYpLiqkveO5uoZBXnG
QY7YQl+kkA7QkxBxSUBY67feb5/TXfnbjxhDdWog4ClrLZCv82hwNIJeauooK/DC
wetg69+srDhutFmMFS8Shvfx7uXmmP7rRWYbQDa7aJOgXjqe8NUsxvBKXwL3XzT3
GDA4z9MKYhP/hyIrmHfgU+4wHS5HK1EV8fBor5X+MtVsGXpkpbkSd84YTzv6RC9D
3f3DYpgXLJsJCXiWf88dp/UPPu1ETt4Y8E/85jeXo5R78KSNwERZPl95l5js+8Sv
+AuDUEdbnguNU9LWw87XOAu4OMcThCDH2tsowNU80iW49f7fzFJoxxofCukiYCVS
fyMzMS91N/s/Lldw/O1V8G/L81GCYQU2PPFDE51u9Z5JVcRF8pgykBIgquMa5TeT
QpSafLhFsY1V6I6m2hq/kj8aWkTRD0wqdpo/+Bz5ySufcHjXFKEJwDCIMhCTMyjs
QEb4sYXw4ZitaSlTUKAtDsLgNm4cbbTHYut8XljIlgiRIm8FscsgfH9xsUPmZYfe
JElUt3Y/ykHbCb1+XUvItFtcELNuqsuzW5c7y+mY6ob7gZ83l0CC5OUTrcV//csj
u+JhTDWTAURJcfIrqGxOl6U+b11qRStGDM2GOa59qgYDzOyvp8niat7H+Ad7fWlE
w1cvWAHUC2O8w95pXCneQ8PcKgGRmPvmlkrSkMBNh66FO8cdZz/lyCYFKcAtdQDV
y8MGCAH0WiKpkxY/EDwY89Wjh1nykz9FIW+hVyLufBJQaGRjTHk/Ubn6GcU9xjbj
raukZDzUhK4/1tNHB/yjM6vY4+bn9a+lagcD4U9JOem8AK9XM1y21UGNyGQjU1DJ
tb6+XqzTI/1zlmu3VBJR1ymtFxZtNEfl8eSYYM5a3XkewiCkwsM++B2bGnHYQkPO
zzADHZSTm9Xpe+hZyTKXxK2dLgNqGNkifSbDwmbfihg4wCedUF7PF2ANAINhHqxZ
CUTFjccGIVVoXHLXTFOGWp5XZyQalNXXsAw6MGA1/+2cukg7LON3tOC5jhmAvU9e
a+HYQO73FFOlsl0+UGqGbUuo42E4ktz/X1RbWV/waStKkeOKWR95OO6tPbPkQBed
kPGoKNCJTPBpaKNFFMYmf3kPYMZsxv7YNZh6sMC3sOaWrmz0pKI7rdKDtTDqk/db
vtf+lctxj4l9pdJibTtI30lvH+aKwctClk7mRpF1mHkta1m0eTV2W/Eux312VzRP
XfWzEHxO5gvsDDjR9HZDSjNNgELYSSeAaIuRE4yR2Fa1J7fU6l3rtENKReUqhJcz
zx1uS82I0fd4KzX10l77+Sx4/sGrv5218C9Np7dGDnwZos2YQ6ErBCk+Z84X+SQo
X+iuE3OWqMWSf6AaJWcYhmImM+4cI5Sb+TQqzuklLOEUTVzcHT+qVRqWuyypomif
jX4S1NbllxKDnLErOyIbNez3iwwyCo1pBSDQyXSegbekVh5CZCm2l6qMksiXpNrP
QPBNrDQXYK30mV6ndK1JCIzhSc4mt2rtY0EEXETJellWYbNRofTY6ksBTvrrkTQT
Jvl49sKgKJuJARNGhevArVSoaqyPAicA1mCrMBoBS0Rz0jvbY/D6xsj4LWei/62m
C9FZpd3Ge7CohtLRXYdHGtnsD3Le9/9KdyJQKVY5Dw23FEmgKQjln+8yOIIpxo5U
zHB0G+/AFjKhhvGxaqLc7689EHsc3KJoEfMdy+ge51WwwXw3mzTnoDm84YFrouHP
Se910FS0UVE7fUXAGNi9UlwmdrTDtMvHi7TGvAGOouq+kneVRMIA9ld7azjDHLU6
lBNCMKT43BHP5bQKreUvt+1GF5OI8LB+MWmUJNyh8F0SKLRQE76YuuFpdqKlhYDe
rmDM7PM8R8/ocXUgP9ifOY8xr7R7Ibvlb/igjdK43zvy9A7pBHmQlxwGW1XwcNXf
16xaGdayin5NLtCbnrhY9G24SiKhTlHiEGj17gEs7uE48cUV5HzxQL3QFzRr8fxT
XH3Sg+SNO/6eEPJZDoAfYmN1RrdmsjiHIF+WfsAXcXgABejslqWEmhI0zvBiuv8E
OshdCjoyXwsrfDcTtW65n33nXuS+pZsSrtLdQjuQT4SKvq/AFsBUnin20Ps5S8XJ
oQ5edcjtzMvSOqPjyGAiflrd99Rj4DK9B4Ltog/d3yDM92RxZ19ArXxijR2eRROe
457y0eY1V0XlLM+uzp/fBJLRwPTG3w3FfL2hqxy7KnLYF+ptDDE/dSF0EOpoM5P0
7VATzEIuYlPWe0Nv3eVUcOzGE9rHiW/BPe9ld1ryPiQo2iLxalp6yJ7tXUwA6FVp
cAbyFBQCBpk8gkh4pU2aLbB+3Jb3WGTn9WHld4TSs7cNwkXLhQiv+hnDmu01629K
sYAyEnIjRbG2b2TBYI6TldxBy8J50JBVIroeJYtFA7zjI5a2YjP+XQV05EAMlj8G
2JuFU9E8l37hpoutI3KtNXILTMB8Z0gpBmydX4rjJB77GOFy7qT+fgMMgMnhWale
JZZJxtaodsUnV2MaLHFMsyS8FTsHUGTPgk2osbvBHbiaovfKr40uVX551sXNCaYm
yrjS1SMzteb/OAO0uPkRl1Oyb/v/rRP2M6nI6SWGWkZP4wON+vKrBx/7+sXHDZzZ
asJOf6T7oyFKnoEQQF9S7v3fTEMdWTKnARckL1nx4rQOjPUpPgstocWznhUW3yhS
F/eJK64zOgJtAfpME2kOgB0gwYKKbdS6gVlUQTMIxqlODLlSjmzBToAsJBEMootw
Ye8j8nrhRzHzEM4JjkfqIngjstxskCKhN9JCJol9PZqtWwNKgiyXXSmO5Xmg8Wyn
+uNBLRTvPH40wB6S93vOyIwVSyHZp+1scCJ7Y3LqRC3MKaUsLrN5+kbH7NYNm9jp
2+J0CxnOH4pqv4d9t21qx3NwRcPCoqcWX0cWM4KhY2Wzqz6iK8tDd30LUv4KZf1t
l0h8Ih4rLEr9b3MtCZqUQA==
//pragma protect end_data_block
//pragma protect digest_block
s3guskFruWhm3TC+sGSNYLEftWo=
//pragma protect end_digest_block
//pragma protect end_protected
`endif

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
jJs3Q1oY1hPccNzkZU0WWE5iwhAhBm9oF9Gl6ZOzyek2Kh5kvu1rt8AhBrYIlhy/
q7aZC5Q/Ae46wXmGbXFjQKvoOMUjbOiX97XTztmGOITkiOOGBo7D6TgtkSSmDBUK
SyVzOS8VHatJqyUPJjttkJmNRqrYDOipbJxp90goUSxHU7WjE90J+g==
//pragma protect end_key_block
//pragma protect digest_block
xGck0ZjPku8nsYN35ZO3rGqaciU=
//pragma protect end_digest_block
//pragma protect data_block
xv3RRNj2+LAE97qU7Yyu5qsbBzP2mTCRDfMqtWD/Fw9dMZyndX3DOE5QLJF1M24z
KU3j7ZZtqFD/ykLHOuFjOM5IqMq2hVv3fGM9mI48FfgoSfJvKiabfV2UnMXA9ipS
Frl2nt2JblynfFNdCcM6x2Z1x6iWTe2Xd5wPhIbo3yCVS0+c+T0FMN3/3e5bVCEx
s5ze0keGR2rYCZ5k0XH4qz1XgAExPGWrWYVWHKgyLjNjtQ2Yn+mktMNg35oqLZso
R6anlbqkysJyAPeTx0u93t8+FI8V7Wta1lxDw2dm36ba4oR2lSpo3M/jGiSWUF/N
3qS34+vJs6nxxLlufYPECcfLvoQKzIFUmA4XUp1mnLECzbfM7lCWU9T2KPoi8Q0j
ZZeeXog5eePwZ6WXlqqrYhAnswsQKPFQDR5kTIFbdWMjWLPwZxqFicxIW7dvawdn
f2cDI1eFkMNU8rvBTQSx2vm25zJjA0RKT/gvcqhOgCPSBtm5kYnVOQKkkZi2/TAU
PY47vdt17KIW/Q1sCqg4phF3GeXoBXjbTtowzJKbzm6hjDu22TdmglRg2uKS90nb
vny2N0cipKQhjfqtHGsvYEeg4AmQhLJVC6c0p/uPCTbbtTu/GbD6zhVBWQfcCoSm
PQq3DI05OANDom4YzbacJfbO2exnmEq3DcY7mpH8n0mWTjWXcDO0WSUM6SuZgirm
zVbG8Jpza1Dtq5mLmZW/sBISwYDjU60TRPFb7k5umkd0qSdEjkb1hJ4HlNHVEYdU
XvaC0t/CbGfmaPiOkP1GVngDM3EnjtOUAbs8BoqHx+2SPEdvY33PzZ2B31drc2rq
1VbuMM0nxjf1lA/0jd5OQil6t8V6Ax7d65Zw8+mf1XIp2QhJYMvFCEv3N4HuwSzP
DzCpjOvg0L0VC3m0ebbbnlF8TgwP4pDzwBGqdJPaAaJL0T1pgJuqlnJtzvg85vG0
fAZfJs5zDgVHh9oujhZr0dcarDNQoi8p6VV+LYSZvt85PrQoLb9h0l4DArEHx5pG
Gl78h0simHN96KjkKIvplRIkjeItUJkuvvtzy0AMGDE/rJ1ag8fT1hsaIp7s9FFX
W+tZ3tydqIDUcn/Ou2yI4IcRKKpImzEhRLAw7FuDDrPVey7C0kSLjv9sXHn9kygm
B8LwqTMVN4calnJkkSUpp4VTCvWvT+4IggvzNkzvJgYCdTRTZ4I8U+FfZ6r1KEMc
C8vOZWnFGjJsfB0kiD4hCOnch/di6H70bhrRDSYPhpAnm32rDCdkRcOfLV1hkKhZ
T31+/V5W9yqf+q3vpiCYsIi3TaU/rW6G8RoS7fOKyXRjKGJWGPMN171LMv8dIm2G
X/E2ZcdwULhTlbGC7Q0Mr4tAhENxT3/C3BxwETJfJJRibJ68m7EVid0WK9pgmZt8
bhFeIWglWAtmCCr6iMa7obHPnyhO6mLXYxTz7HbiurpM5YrC9bHh1j/vtyszJJhQ
UsMyF1ee/693UDTMtP8znCDAZWj04C56mlZtG9C15v51+T7LPjSlncqo6LtO66Uq
THKkwbo6xWAspFf7yukwrIrG7bTu73ihVw0VqSAiKX3dwcjpGit/UhPlcMp4pxnM
knqj9gz+isGU92fZk8P66vNrrjhiYo3JV83dlzQZYV1WVEtill0MMajayzrhuOvN
VV61x0QBnW0NaThHFvq3aMEbk+RtMiHtq0TerDGlGA6MpVj4Zwpu4xd+1zekf6n1
2Vwc1QMjCr5qCAc6Ximnit2fAjsp12YTorS3bGrasTD7uZUS/yz78EmqsV45ozoz
JX385FSe+elXkeZruiYyY89GsdWLCUpPkl68b7jq7lOKaRhtu5elpscMl10ZWLeM
eJgDPdkJE27jp68dIOfjZPvASCsh8JDn+psvWo7vEFP7DXrTM9vf6H9lsauPHkzm
MllG781dfVa0ztzE8WUaebIOkGIAvuTGvI+tHFIjV6YP2VHLqauiOU/UL032I1aw
QnczAbxU0Fa9u52/+1STBSp9hAuYGSyIWO4CPc6eQMVhkN2FHJgFCwYsUNNTphQo
Dc1wuOT0DsIHcbGmUYMe8spw5eOyzy22gTKpgZUDxWCUBsUhhpxRScZgKjz+6RfQ
0zj5VHyngAejrnD6pg67tfAa/hnTax3aAwU+MwVvN+RfUT6KhStr0oylMRsfnSyb
p5E6dfw1GwQTpkL7VaL1Lt9klZAVx/0Y8926Asuo612q5L6LfhZZJhog2EU1TTee
WWdkeeCdBgWkgsjXQR+ViCgM34GwhtM3dqvLVzHEESwTpLFL52BmLCXeItWA1VKa
yEMOqlSMO0mHE9RiZFh3lskVDpOF9hnbwM0gJukwS5FNZqG/zh1iyUF820IqZmZx
D+IuewAGSW0fZfEJuH+smEyQJvXkcbrVgxNU+KppYj5HqXhOi0X8eYnYRC0qJx2e
2CAg2rmdOchFjjfEZndcKNsZ9IdgX8Ic2mbA+1u1I65l9BcdFS24SzkoqhmWn6ax
NrR3OROGwK4CEA+kEiZXFMe+ZOySY+GiJ5G06R2GAvV0l6hxqMhTuavoCw6hN7eg
KjNTLrbQPyhsXawWsAFmkI7xJ+g6M65EQ5nICLJvHC4uF8bXVPNmoi8mULL8U9aF
K3HWBal04El7mpCe9O8wbqRzirwih24jQ8Zvun4B7gb8HheZSAqElyY4a9UBv1Q4
owq5xz+MeHLCK/M/DSg3tohowENlgIw1A4O/aKPPd1CSoGvfvnEmYIj7jAB116Wr
MorcrGghfWPSSnELfcSirKdlJygfoctUT+49s2zBKFzPLIvBhqaEcsFwWWN4bKOx
HTydYLU8NmgDrqALmvTTS7Vfb8Dgk4+C7/UGAc5YxMA9m1gKVSAWcuqc1llsEzmZ
Q6vxX7XdphLT2IVEuKtkAAxJydY7lh1EBG6Xl2WaMQDpS22oKZU2VS310joz4dsh
Lr2rTFyAztpLUCWD+9L365BvX3D0AaT1W26E0rg0UGumiAofhTj2fLV0FuIUi+h7
+3bJbvuwUeIkaXYeRYTZhsh9Q55lQTVxlDNO9iHuOEnp0WdH2FifWNc4LHf0/6mu
MJx3rrCql/CV0BHnBV9SpeJTDOMfTeyjoDCJy6X1zHVfmxJ4wKhpFEKspb9GMCc/
Avgjdh4Y6kE1gpCyVCqPoVRWM9hBbjEZDHVHtXnQGFojg2UW1rNmk/tF52Wz6gUn
JkrD1xhB/rGwNgEFizJkZEEdL0alSkiWahtn+0ZaEiReY2Ma1UADU+GbKcISvujP
zqOSR0t/k4gXLDdpW67nJGIrjwmEJqvv5x9ZFU4LDHcqwhS+CQvE5YzkOZAiAKWU
2K779Lyb01FaAALl9ArNbd2VyR+2C+t9Yo1V390iTYbgx7PcR0PtdEZp1YLGj2A6
Tc4vNoESFHuWlbaRvjrEyV8s0koVC7LPZV3sKfkiaoT/N5/p05ua1KhnjPYem6oS
NsCMRh/o/UmcbcIpZdEj4v72lRfZGXi/Yytmt4DmlYDaNPxzObxiui9YZMx15e8P
NaT7x4ShxvTm4QGFefIpQXSBJbgAUiLn+ZpJDz9M/e7XkvzViu0LAwniXHQ5DbFG
jo/fLA28ttihO77ztuOKOWcMJOx6XHEqnQeXZe/yjxf+HUAYUgUzN4L2u94NEnnm
r1RqLWc8qE616rPU74yWC7CVgOb+oh7UViwva6PKhB41uIEnDYOKRlzDkWJ20gdF
hjufp4ddGJl83XkHXpdziM8BGN16LuuwbZI4InWemKQb8k9b3FC6yOIDkEKImupR
0jOVjIdtgbac0cIyvU/9ddNAQm5TTPCfL2h7BIvCvJacZMr4wMfsQDIa7iU/Zh/l
qXzsAzKoNbxIaP5HdvAq9FVHX69biGd2WaT4dVC5/vPY2ND9aXKXLKiLgEipdv4B
Qdm8kWV4gwVXrImwBDwcJoSBJNdaZJniwBPInYnPZE5le/aylr+wDkIKI4kZCxFd
pWM4VoRXnii8xAnUMTgKUQNbNBocfJIeDEechWhQo/IvvU8BwOWZJo/NGzo2oE4L
QSo+AvkGvBxGoikuPa2sUgdlSNxzCQezWSmtj7X5CWYtR1ucSo4DoLsMLZVTu5JH
gESSao9PzMtfZ2Uz1RV6IONBhWNdWbLIqyiIh2xdGC/ipd9yCySus4W4jXuzrev+
cLmI82d8AA97gEcadYM74nPNdm38HvonJU2jo1dTLciffs4jQ04T1AAEisUKE8a5
xpCQpHV0JjuCUZ7axBcayyRGpKnFloAIqLxHugt09aTGRpBaktIGi3z0QYM80NM0
E9jrWpL4qZWJ7e3OvfTRrHvgQCH3/+DaZe/cgUSyWGUdPc5DysZtBQA4nbL6K+KB
nrm6Toy7i3a91e25YFv1Ll9NxvODylMVSV9hbIgWUWennotc0n6lC6RaKvIpeYQ4
22Qmw2QyPHPY+HusHQKTZbmZy+Y9Ngsm9GHaH1B8PzyG/itcUk+RYGk4kvuBkQ0c
pjxF5VNp2J3NbUFN+ZEPtZCVyvTu97byWJ7bokn2JG+F52nDrg2yAwHLTdQt0xcX
RWn3ayVOlOFGsihp1MqERDX1WjakRA3phoQkAjkiGWmcsIYT6d56jTTUO2dr1SqP
49Yxe0J+i8nBq5KDuUdoRR25y3fBsydJM18niChfwxefKt6QbQWmTRnNlJSaWOwE
ubQWJ2LJwhBPCU2L3f+NEB/dCh8F1rCVDUZlpSgnxjmRrinTBvtDp+8FhtEDQjh6
TVwhusWrBdHOKl9TB7IC6Yi2K6nLbEzQI+4usFfhLTc5J64KbEUIPGvwgdeyGVbs
dHk5Qgpt/EXxvkbFwUzXJnfNlkFVAuYi1ahWAmEdMaOqzsGttU+BN3KuXpy3H8hW
nobJArZb+11DKULJUSu39/OTq83Aojp7PBZDe31PH90iF9N6gMjhEt9xGbc2AQzf
YtF+8LNqKK6I/M7S7MN7NLNIfqF3yy6lIyuB+vOVs9AptSlFybYdBTGiu+/O3k1p
cmGU6vOq6gdvfJ99qXxAq0XY6KxSQQE1nyLtUbgbMyI7vusLYZcd2/mbOzbIZc6t
YikYM/LQCWIz75J2UldobBY/I2Y7jLNlXChYYAE9QNGW5sqHkLZVOGs2Uu4nx7ln
tNILjJGOlExIhwvnYcqnHA4Z1afJU9MJ4v+cdKmSt/5cCIB+al4qFwi9VLCjCgZP
WSTMb9scDjnzNwm+BefITh1hxUVKCo+E6WeIWMBONQdgKwvMRLUiBXpb6kPm0Pnd
iqi/rT+HPzuZ44BQYYtMCVQgZz4izxTgmgB1+5DCKavfq1qpn+kpRYJ+DihCd4cG
80YuWVpx035+SiSyJ7oqL4YArizp4nru/M4+qYNK2uEQdhfOOU379AQzzYUGshpL
bFtHMY5N1Nidnqm+FJ+zc5JqMBHb+6TyXMmUQ13uFUXqjeSZlZZQl5zP/mBZjEBT
ABhH88MGITqjQKsJMDuY5qvhHaBuzdClMiNIrLWhu5Hz8cN0ky6+koN51NBP3OjO
k5uddZzWsVJsDHbOEufwbPQCNvAGAEPyPu06LrDsRdij25IyeKSkpA6K3i+RlFtv
xn7zGgY06C9ZQ9Azlc72bPFvofuZiXYd6hFVR8Rno7VHUBOJ0Rzxc2bluXIB7La5
kyKGXxQoprI/ck7Po19k/2AadZwRoqKGiNPL8f/9T0MsmmcXGZ9OHLhcLidIyzQg
VhNkTxkMuqzbMBiKNw9YBQ1xvshhF4oIB1ptDgYwWKBVBEtVL8Ft5NEQCGlY69Af
PVedSb33yu7al9p3s5PF23wygztmf0k3a7S6LWPrb08TZTDPS9DbTulvgNK+HGwo
+c9zpOG6nNqwX0mjkxosVznjcpPUKa0KCjQp4uPjO2iTCNUICo2J0TPx7fRjTEtA
GZGCbMSLvC0ah0a27qOqJWlvUWXZ7DOe/IbbPMMtCtrHXfr/RcSoENEVGCHY326/
d/4Tdg/KYuAYTiImwbeiT5vIljAk7Kuv78+LZH6/SEsU1m0ftM/EDwtamLQ2JEF4
gLmtt9LvQRSWtN1UL2sGlOvZn86o/T0qO6qjqqi4KmOfwRCNgBsrwtgffO79QhqO
G8DEVoqLr6JG/oWC/TeLHnmTesOTg6DPqwHKr6dfc5YS77zx1Y70RA7tpSkQWtKB
EWvCLFrg6YW/Mio+EEwcsK3RvAiRgEg+1O2/eEfnVPOHarEwzqTuwu/btwt1ZHHp
pDXiBRFzyTWDcLtUt2dyFE7PpYR9j/ikF+TTvK4OQWk+kgtlV/xeks7AHeewIijX
WxvDr/IPzPfH0twFV6Jzfk+AhQOV5dm/vCC6B3Q2H87JrCv0D5j49FtS0JqWCbcm
3AtNTPjpHC2ck3t/uk4KTdWG7jm6AitQJGZfZXQ/cOF0TAcpsEUp13onQzCn2Djc
RydvSPVjvv5p7ymfFxFMiXtCtpf4ElRtLGIvTVkdua2kjd5S+fHLYwM229FwN0TL
xG4eaxTHBlaPJpyp6o1O6ziB20jYEnfnSCtD78SFv3uxZGRvK5j2yqTVj83WpNo/
Ubl6mr7FhCArceTSUcI6DOKDn62GEVqxD7+RD584fP0A01jw74Io+F6928haOXOP
f1akBQR83/bJO4PZcKGSF4evMbDtGs8s3hBE2uYZ7VvR3PeruQ08wjzost/F0iTA
SspCuY2mOopQnZI/XnCKJJqAm7tUob3+F2eCrYKGq0sKCeW/mFi+9ojzrvvtvlS7
0j3mDR9xJuSLJgnuzib15qabmcCIGbF404F0nJ0TnwA+fls1q4mSVSUFSVm35HFb
OicfZ+X5WmFr0q5FK95ThilOxA1tMQZxt2OShqMydtIg5V9Kt8zeljBQ9US93/vH
og6pY5MUrZIfWzOzGy0vzikgB9ah/p3RffvlzSAffjlB50psivRfZU1tUgUZG1nc
sFIFkOHGCe2vZIALyTXGqRktZt3GyPpXjY5zY8qdPIlHoeFmgk84rO4dyicelFC7
wziVI9p/rwgOtQNSDhhZv2C+VG8hP7Gt5tVO7Yzfop6vZExi1lWAmd8Bp0huAIc0
pckEzS1boaPzq5UU15H7Jw3Q+9Vqda3OmsXYZC294W6oDMT7bVqmFX6+6NuDM4fp
RlPnrvXcPTFyRx0E5NvHIq6N3ZgcMlCyJSR7YFuspLbg+dC6VQOsc/j7Nqv/VZYD
vjBNa7CY4sZhlmQb70Jc5KQLap/BGt+xJMMaVCcfF2ckVNpnZI4qqFjuis25b+NO
sYFYSqh5Qm5P1V6jpkPEFGQs9i6Ruj+ifnogvsnVPtXuHuqxdsWUnQwDE+mnyDxW
4ZMfhzMY7oXGdeoV+gLdeIFmIY/xeOtzOX5Yrc+qtGKVc5XShibtVcPuDLQxvEam
9JjVBzAqa+mQvfVpUHK+hRpDM8PbNigVX4bgXLmRFx8q6ZYcDWRCldg22DSWJfFH
o3d0Cu2OqlvqzDRWPE6ZNwdv4dY9Wcurls6nvuhNMzMR92zThX1fj9IL2kAiS+1F
Tez6ddDZLB5c/+gdS6tezoZnht/hJansW+UKLMsL6cQaxLu0ueiVG1qIG/p4d7Fb
eBX53dmTGyvYmsOu6l3Ej7JN7wQh6glGaDlS3bdBMt2Y2QW+hFERPtnlYTn9HlRK
U3bifibbK6wia9zclR2QDSuhbNW6N7BOZ3+GubaWZ95dflEKft0SCmuHU66iGZ8K
XpU/wEkfdRoQKeSt3XjiP+3ZTTijKQgESKY8vIAVF38dW8LBY/ldX6HL0MoYum4T
fUg1nE1YpdPyOSMR8sExVfW3ETrWOiseDQjKUSUeIihnZYoHBR8/4ny1l71Snauc
r/S+Rll0UBGn31e60ugq9xyveeobCUpcIXrYy/Tsg4ycQdrU0kARDDPSc4agymLB
IKqBRSSWtUvKyli31saGTF7mvsuzHOePgMVD8VOrWDdteI3JKZ9ATPr6hrrZunk5
K52IpiaBlEZVGdUj6+8QzLJVN3G23tLhf+UIL2Wq4hHiyLEqYFdDM/iW+0jHPMVJ
xoQwv93/zwC37uFU0gMImAdDK9ukkSY+PmLH1dj/oZHfrMmtKADucQRDmyN1pmYN
mUCk+yQm8d9TwXDbh/tSGFkTTnRLYB4pe6AL/RSoLGxEa35PpK4oIsasPLNrbNmj
hwDdpDJQTJBRZ78MO6xu3RkZhGSWFvAIHhSPvIskwIPceKahmr2gMCEmH9AZhV5+
Zyf2rJGBpCYxVmMxECqltBwcy91W3w2KFL4ffdZt3cZaM0beVib9z2q1aTZRiN4U
CxG77NTmD4gE86LmaokbWJ5TuYHyKynOmY+PuFnKBkhsf5gpSl1w2fVH8KwFBcsP
2RWgOLkmvhKo9u810/ZrIHUGkfMYdzni8zS+BpdxX1LX9UvZI+l5rFk+liimAMRn
d1U65DdpxJXwNEh6XNQgUgANoOcU/iQPFYv9Q2oIc+buSml+D4jXzTrlAy59Q4v5
81fRk4biXsGXGf0JALKt/HBvVIGvzm6Lhtb4P72+hs1VeH1xa0N4hVqbeWXJSpzj
GfmLNqpbajrlwhJCFMSY13ttzcvfDxA0z2ICvdJRo3or+fI9ThSXuWOGwkTVe/53
0yKX+bBAutuelSC2yn6hbra17tPg8nFwmULmqqGZhijbHsoYg7ADUrQk8D4R2NBZ
GRN4zsyP1kWJiSHJsMkD1A0A1ARlEa+ySIqs7lEo2Ysz3A4xTCUEDSgNZKkpLt0B
/Dt+ExZo0+KBt1mlxNQok3EzAvfuKcHDg7Pg58G27pjjUQOzsJgYx2sj2j2gbxUS
/5GUO/h3/oiR8Js3NeIOuj+ClY6UrRnd5GcBlJOZtzxzabnZvc7TfPGKPqK/epAC
keRfGUMoQwOEGAFl4WDzofprpvlM3pUWPoISR0fJ/CazVhKByJ6VBhCa0JLcPVdK
jhgkYmRFAJwM0gjFowbgbZqxK0ZVSgJcK23sBiYK6lEjZgFa5g6ua7z57ydz5YjX
tZNkugCVVgLiE+e48pq9upjmNycdyD/KetFaF1NOdUg0A3M5ZEHFJvWipn5i9AFa
wx9m4Mmf24UdMrdYsxuyDr/MNmwdFZEPOjZH9NWYKGkIaxWl0owktzwVOGkG9Tn4
jtjpGWu/O1dy5BJggRbgWnjctmZyWAyz2fJTp4DxyLN3It1LBnln9Qa05o0pnoLk
aWMp0zjUt5l7YXxKg1CgK1re3aqICHQ0rcrtyhZB//NF9FHfOPGSAcR0CCMg4dun
+Bi4pA9i/g4l0Rzc61WVW5ufQ3PNGomtwMBBZw4PUu3CrDLgj760rSRXI8KbCTYZ
7Oox61uI/XN8sJWMNHHgiQZWAvaKmiH74/osy4FfObYAW5BaRgS4S0G5xaAZHvb0
oVtAjA6Lj8XyMSQUyPCqO5idWMjxNpHvTYgq2ggTbMahWvW28sycm8tc8t+iu5pf
Qp4ClWvfKmcy8JnVTsz0n/JK1YM5BfpihfuhGz53lMKillbE4CJmcYKzIkM2CP+K
MGCxM9061iLXxdPzswIFs/i4x+Oh43ds+x0LrC0jg5NMYkoH1TKowVC8n9LOF7Ly
preT9A+VwXYmvTjafixaLGNJpMxkpKM5v5kg1ZjMw1zHLiF/Jf2j7jEkNnPk/NKk
4Tr/iLInrNUnzQ3SixY1XqQ9b+eBEJ7YVsAstT2B93BxCznuoiwECx6gB6IXGmqu
1h/jrz67ugksFpmXz84WJGDO8AY5PIjGXw/eRG+UVEvY4wi/5NNpCUAAsCJreMMA
9QZwTXka8lfjwj2l1gPDboNX5YNmxM65XIcW1I5+b8w/N7bBM+rlTKogtYiYiLpp
XSg1vDlcud08jHqlHb1OuwD5v81EwHTm9eybPLMyswHwACqU7T+ObZ7FZhWq0hAg
ARb7ZE4CXkrCd+tqPN8ldeDK4CsDUymjOEOpasy5MmiH/ggBkWaNJ2nmLT608y1s
jKybdEjy3AVsAvF2q2CH71Op9t5+L+7x+c5A3K3/RKQRl2p4BTcVMZzD98SGwgCZ
0fM2FgB/GAYvfOOo0RluBLy3XSzBGA0AqIEM7P+A5WXhxEZaPSmBSGXyT+NHtYOa
PKs9/BmeZr3qkZRMxLO+xz/VBW5fvPUrMaGT5HNAYYN1OJP/GIyxdPq0v3idVJys
a3rgskFVkcaXBnpuE/pxCumCBDgPe67yLlCI+d6FtLBpx/pBt1wRbfNRyosjKVk3
ZCoWN+XeLu+MWAflNusvLXoloANyFAcc+tWny04d9n7MSoZZlsFpKjH7I7MnUWIg
Y+KFlxz/NN8tejwoC4B/GO7o6mB77Q+bwyE1VMgdsFWAQ3yEQKHKOVm+oN8Ns/wN
qQAtet0+GlEjGB4NfTCSnWhsQ289Dj3FcnRZwQ2o5CrC3G4IHtYqEhtDd6U6c1Xr
4nYOE0Hw5SV3r/QzvmJs0wYTQYxFTUvfumHoWrl3+vC7NZlfSpy01a669kIxeEcW
vs1IE3/jZVC5Q2EXsT7M8iD+TENQZiQxXH5UnXxGfDUsdk5q1SD/E5gN6vnJLrxP
8Bco0vWCrXICufqOAXulPSaqRwKPGq2+4CWRdy8eqrTZr7zDjj3rlKif74KkucfY
SoFVXX3m/+Mber0dlMSpXXL6RsdNdUDO2wZtRnkFpa8mRwE+er2B5CeYcll+JzAI
jNTAK8i3Bhx0sB09aIpWTkNYU2MSkZzaOX2JC8raSmtOyzoqV/IFkQXvmFmwA+Mc
SYiHZe9fre0g3KiEuMBdOSsFacIpiiiwKNtFV1cSDzMwNHyCd/Li4LU4idfsD3hq
O47IrosZDhHbZKazHcLiT7QEWfMm6gJ0CuXO+RTHN9iEowLy8L684a3hyVjRul44
MD40jb9PrVKsYXAB4XiSKvSyXw2lnfwyv4fONffLwfqKFvCLG4wwxpc1HreBDTvm
3eiPsYfV4AVhaNRbR9niSaqqzyCwpQSGIu3ly7YzRqVAXO74i1g9RkeyaAWJFXic
H4Y718HJ9PsM0wnjgd49QkP8Vvjob2R0PIyIx4Dhhi1gJN4MQT8GigvMgWRFIT0a
6+hJ2Ign2bUn1kN6yUtyk1uJ5nqRs9rZNd+WXikYkqRBzOT1LGWMsMtxJclFRkzw
fiaLFh4vluw7QVPT7e/EY1/TFy/54AhBhOnI12nPW4Wrraj+EBpOEULoW3dAURi+
vRdAZgqPYbBIB5EFJrvhuYLZt9wj3N+unIhRCcmjlsKVuT73qyfm2wQjK5rU+dEZ
7c8GAVbyrAM6Y5kUXV2fKcMkuu/YjAfM5YI84EdubAS3bUqv6ANZHeWBa3OxMb3e
b36u2s/1D2rxsTvZFwQjiV9W2O7Oxbua5GSyyG82dxA0gcK1mBkdAIbTMlLF5As2
C/7lueyPTsKHy9jFe4h4G3xHaH3udoTdZxdOQTuhyZ3uk6ZvEnMNW5NVaG/rk5FK
u2lnBWJySy1ulxCCaTa8gKED+8+sISop7glOqdt6enHOqScWZsBF18bz34zPQu02
JjDJgU32u6GEeXeIEVEAorZwaoPYjkbOQ2TeYpiQ8t9fT7TUG9HVbXiGyFScgtoG
4ayF3XPAnibjKaZ+KKaxrzeO0BRrqYpAX/oFE+Us47YQsQWL5ClozF/DLXx4B6d8
+GCetLfMN64KhOBHQcRkBISC7htcKrDD9fboleK2HwV0wLjzonNSGTYqbgorzypm
tr4u+cqQ2+DyuEzNvTI1v0PhxBGP0FMNdfE5gA++p/Ohx3ldO5n/0MLC4SBNZSN/
okfVI+zj56eZP4WbBZwMOJiZdVJaqPvKLJTYscLv/Q7jdviUoJ+FYUc537Rp0NAg
0iYFihwk/pWJg5f4S6CWoTJ88GTrBV/02IZN2R0e7MMUyVRvSLw5sfqO6VRvSG6K
GsJlDsjODTTo+DPGbd2cUgVa3NeAUX/x+QXC50TUo6JC9N0g+jqdY9e3WwCkcILF
gJq/DZHDOYSG7PHD8d6yb4W3Z2qqSvKNGPNPvlkHdqZZhlLcz4eyy1p6ZhgBTmLR
vsD6yaCvFh1WBameqcae5uE2I7yiBa9e5dvoe1yYzdPBuAs66SHf8dZeiEKocIK6
VH0zQp4Sc8kLET6IW/jj2fFOP0nprSAm8yJejdxMKAGK8Qw5602oWLKBP9NqyF5q
SLfT11ZIaC0GRfUEd3F5H3wsn4DZ44kSvvbT7HoBLR5eUzWpeSIWNc9HRNdL8FJ4
jFQQV+JJBq1vtihOUSE6f8dDBuiAZbAe2XgL4OXoPesDMURafsOyB6r/yvbnN8bE
IKPfTtGpkHw1AbAA3U12pl13t2NH0rYRwpKkrxTwv+5k4Rc5kZ/kbBnN5OMLX1DY
uHdPbDYKBWWmBvOYxRAZSBEkGYXGzrIhOYPBeWaS8JtFONcP8Ax7TxV2RE8FkcyE
eFMRjN3uVP0doOA3GEzU0YtRgwR7ckGxWugHsXMVabSPRWyGkjdgNyPBnTUcE64v
sXGTSVLDLh5mIRFwzO82kBuY63s3pdFAA/P6BhYMaDi2WX7jA3YLBFtvQE3f/AbN
nK0cv4iJYsUmbef5pI1wB4Zit5wj4IiPGCSCI4NxlaBVQone6HIt0WslSS9SppFo
R1Oi+im+WNQzlWa59vGbROto6QFiuTXGvWmCePF7ITmUy/gOy1khs2pBfiSqnviB
8HZUvb0yRPNZ1O1xZdL0KjlgjxzkIcHhGDLReUK6fb4LM0bbi/ghhFgNTTImlgxJ
68v4FgQYYQrcWiKTMyAcLHrCcoSevZosuiSKTZlU0I/dZZ1HwObosNTb0pG+CYQk
RUQshBkqzpMSQvcxKxjdFBzo6HgRH/uKFFt5kmupwACxuBxGIhyKiwdX1K11gHXE
My7CMC3i/dMakLvOtrG/mpAJWwa+j/DV5Y9G2S98cVu7w6Y7iVdo0iqmywCcmvZr
BKlNJ2xtmQzvcmrO3g2vumSb6cNxuCHZAGfmu+wDZBwVESODGK7Pdg7kVcJuZBVl
mZ4yxo9jMGyV41T0IO3rKFwBs9MnDD7ayUhbZmfoA+7PtUrKI1Al4RF1/m0I2v2f
XY00M2bgdax3TCpiSq16lxxtSWcCDK631uMOxf3bV6f9ZWHBqYO60QFNiTGLl3uA
VqRsWIp5nNaZh0G46N1mb+/clVEVco0jYggvPF41xGXFmP1qcDcDQDaOwlM/CF9C
SJaqbBSSGoLixWLcQo4fN9ltMuYzUnjGTwcg/KtKSv2wROt7IaL4DJbiWGn+F7jU
0K6R/qxeaOlzkNngjYBu7fPg8h6zy0TVRuQmLIxc00498HOgjnFuXRtsoDFDG8ln
oMgBNMc0EGhwLsShAbGNRaLQQWnZ/tSSWhowooSVlZxx/FlDUB94gCHYFYAdW2Uz
9RHSt3oaPgUVz9VWmTbQ14F8umI+S+m3h8A4X77t/yGkr+0+MaS7XIy/NMiYmvjl
bfH9pW7T+MD0GNYqdm39zhuSCl4absaEoKWK9bAxPxXiuVULtSVeA0n8/944SElU
n9a5b5V++31iIwVq9hA7/RUqIIl/b2/mgpH+xsRarjqtssti07hO0disof/wzAFh
5M35Vou7KptckI3RrRTux99xaAONC8Dyn/1rlt5B/u7/5eHEFOhLnjW+UqYMMIar
1H6WjdOJiWrOXIhvJmkFghklVuZ/Ejf4d+F884YrcFaHlOoGwvyyk/CZZ6hCmCO4
pZqvtWcJf3vAdr2YUhan7wh5PVqX9nDczlFzi97IukqXiGLFg8DHpZfr2RKbfTnv
i5gb7D8kJVdrdQx5k0P6LRLwdVZX0SPltlYE7ucZRWdVEEyDXGCLzaCeQXdajZTc
3oryLzPpqMJIhWMzobCkBcmsZdM2KpwmtSxIUr435lTg5CTMKtyNd3I7xgxTjs/I
u6SpZJ3s9VMuBBvXE1ZKNS6Z0+U1l4MgnRrf2t7AU1n9HmA+c9G2Il7qotA0wlFL
siG1Aci/SQhYrpDQFLD8fWv0YxSUoaBseaZ9LTibtl03MvZaRnCA0LLRdGGjtsj2
dcQAMwUG9fdrpSUJlfkQBfXTmgshlp6yOoGbwG6ALvgCoq2dbOHZedmhRLHEnnk0
XQJGOq1PqhtftiQkJB/aUvlRvQjagXVQU32O0b/et1T2vyc+vPszvFiGVyDGH94Y
p+J5CX85U713lIz23vPgkIyp5N2gPKyAdWOUgypfJim+hQtEL3RaHN4IYyHinEn8
uGEPl8JmYfMAril0nfL5b8jvH8yOtql+zPCAEkZHjnaduBzRkYgNZh4AhTWnHzS5
Q7eLF8Zcn+tmEW8MKUGJ6tEpV0hkRZ29ddFg8fFKdNIWLzwPEC4QwJP8I1LBHa9e
MvUgwiS4jizKiO3J0iYBWRKmDcq5KY1tkVFvf15cf/uYiFNo9bfi4rusS8ZcfSug
yVMHyyEoiPjiF2o9QqSJjMDD/3PK06DXX2rJ6YNk9/Z5BAmuve5Py/HjNDZNT6ik
oa+4RzmJyc09zwKRIRb7Bz6gee8lxq9zCIDcomtFJbyJ+isOfdFqtlZg3PhxqLxv
x646x8TGEmcLy0IEJNqGTfvCiEFQJJIf7NpyBXB78cbVG1glN/db3gDfkA/kdoka
2uqi1eJ9ri0Y3RcPT6UIKEaJTCuMCDdQFR+zpJ+fRb7QqZHSN1zOZUMgIdfv7rxw
SIauZluulBmhj4SKN2fQyA0Trmiypsh5y7292pEeb7R9XfPgdLAAOFIqc77mqy/b
qMdmrjgQKv7kOgvspcc0AAlzes6ZuBmSO3CtTthobxwDhlUiPIZPT97zBLrTyojo
xhy5LR5CtIOwsEhqvAMy4RgqeSym5MznfSgstvMfg7VcLPTrCd0XVt7GvloQP+W/
IYxmDYkm2KZA0vluH2apePBszqns8fvD7Cb8Rkziniqb1W1vP+gT6WaXZ4kbFF+U
6dL9vtIfm+OAiRmU69CaAKrcE2r644uBAAVNb78k4euX82Amp/x09q8nnTFz1yRE
igy+rSTms1/sy2TTxBF4kbFyW2ENBN9CYmK6fB59MEQ3Lt0mKXzv53vLwCM+JN74
pv+YZjO9f1Fx/47yTEIfdgV8aTvOWLXw/G0M4i3n/pDPzmGVV56VngNx+F//tv7T
ybJMbVMDmLuUwMTlA4L7iuLdMoeZjJop5PF4gCrSuD/EM4SQm2PvOtVwu7KtC6BR
FRw4J/j1tERjorGyCvNunurxU2s0NFGKSD3RWjyP8q2zHdPvkRpoK6GF/Ni0M3MA
r3NFLGntm26/HARKGbe2yzKIqwh0Kd0lhmNLoydcC1yjQh/iRfl5zYKl1GkAknmu
wnPRend+TYQWkOpP837HR6Zl0EYrebEaXRm0QG4daUU6AzWyZDwiAGvZkBmKCGKI
FoYeJci5ha9NBlIwNaZRgMcrrNPjg767RylquxV5uYr0jt5oH4L69Q8Hk3oEjq/s
GLZyVnxpFH8fzGZ+7wgrXDhZOZlPiwZDM6R++AdZ3IrXfAQr1RZt5nlCLdEtL0Ve
E1eNqTZvvoPbwq4h59vp7M784CKLAVE/xZiXSfZAwaQ/p84nUWnzTXmiskHNtHii
4+VY7dl0xeWnWz3JTrBn+WTP/rweSHJ+HoJBD8HcrNrN4OFpvaljAkwG6yODwsPl
7j3Ca1hiA80z4sQMNLTCLzsuS16kZK2niCo2eulj26GNKUZ0LactOMTopkPObN+Y
U/RZO2mFNqiFeEaU12bNPX8GFEkW1u+taTZ7oNEBrQ5PCU4jPFZt6t6GaBBhT2kA
umpshThrf1KbERjmuzdJTbaylRuBi8StHHw4+xanZAfGgwFTCfhaU69Sf06wZjTN
eTPdVXa8+UG/Pes+PnIl29nW/ZSuu0v65zY9IOk5+zwAUK+L7/bgYzBMaCCiP156
cadSevS/kmmteJycAUM7l+HbQhPv3+/Jd9cWKH3DgbmJHwe/0rfUbZKhs0IExuFw
cEa3/I1ZBlyM8ILedRmYQLPFHyST31nFB0U0nz1u9aQzHcqJwG3wnKYo531DgPN9
0iHvjz5a37Gk1JK6hEyTS9HjCKvLezOIjsdTwvIDvLYsyrll5A+JYQE/HKiRYR7O
JXONyMQct8byKbOgUH8YsIzLYp8U/XDXSuq2FZPfBEh8mpzx7WM8MWHMQlMgMYj3
oXNOrQUZ1t7aOXn54jaM1vjryAdS0os/v0xgu09/7hT+9DfpitzzNeSdCSOo9v/X
fdjjs2zem7E/g9CC5hMjb2galjiHcn0sUpHzk+FCUADzxKVDY6U+grx0GEQdMPxP
xm1x/a7QEWRpxAoQCiSjB/tkxvrRd1VZ2HbF8Lpy/dhDEYb1B7kA/i/gJh94QN8u
cmxVB6LOqPzMPOY0dmivD7dt8I1yhalD0FJyGjUp7SsH7GylmqZ6wPlkCZUiSJCo
9gNHpu1z0pL1yHJshgW4nkZZO5o636OOuIqabhzNZc1DQwSdHQQswuTObXSuQdgG
d6wboY9DKHwyWa9N5nAypsz8VdIxegzV6Qt2TpcZYNUFlFb4apfoucw76Mn3sier
eJ/JAPZi4bkpUXQiu3phbxkMRApqE+B7+QxG2EoJURzT7AoQhuLsD9L/A0JNGH98
5yL9ClGp259L7ayGZdWky5/0bczUoQDZHrqseybgmvGkxx7rHJkpisoZzLz1tVmL
/ugVS79XSvTsMg6CpdIbKczNIM+uci0yggOyftquhvLNbpKA2/jHIJrXPJBgXASE
eQ3a64pRmakwgjz+/jX4Mgk05HhZvR7l22A+CX72STjy2v9DwV01hC7dDUjScAKG
MMq7/SpoSkEIHrKLmh5FBWBcAvwh7vBchGy6fq1BOM9Zh8QrlbdMRIcoHL/1kZ6n
YGMi8SbUA4IDEsXTsT8IgGcY9ktZbZ9EX/96If/XdrvA8puqw6tW5A/tlODWa7uq
e02ZXZBQPYx/I+p9/2H403NWuNWIPQVsH3Gic8cWym3ym6sOvypja5ouPnIBQxaO
CrIvjwlXoQvMkdxwBytdCQYkeku41Qda/c7BxFX4x5F5ePwkynNOG6kM4umLq2an
E/bkvlb3Gph5KBme9mFmn+Ly/AeFK54YAslCPWMrgsaNKZGGnuUGKcod2QOx0AoB
yzaz9h3ikTbTGrHYe1P+H734nXa+PzCXkbWoC1A2C+75V886YozuiJM5FE2IQQF3
U+R0hbEHST8yJli06BAQrT2xsT3f9NXALC20HyLzADCIteq9yaehqVC1rcoAICIl
CIIcoQb4VluyugP2wbN2mDIbaUXxKr0r3zTlFYxJzVgmMpX9a6p1kamtQKQFsThK
pBsqVUMgc9LDDCOOFN8mwKDTkgjp4oX9SmJRNmiVROi0lvbeoPNxhhRJd+8NhQys
k4J8F3GWGIbVJdwDJVjYS+2QoMVC5WcazruM0RvY+vaargBhzuNv7yV0g0RWxytl
zJE/a4Su7KaP1x3jsCtzI8GQhjYVbmC9t/tAU+9V4zcvz835/Nnx5ezwNVlRtCNb
m819zDojdBmFbqsp1SqYvDQ1GCIn7EsylOcFwuu8Y0FKkUYlMF9cxad8Pv+QGzzi
DNbC3tBmCgiuyGagJfFOACiFeK0JJCOw60dYjmySWFeiSK65VG2g3GMijVB+dL6f
tp3wE3ZZ57XmkAbvrzarbX73k1weFLBK7Ocuvtx/U280Tm/iSQptGJUIviWZSHrV
pWNXGfsTLnMxnQtZNEJd9Q4QaZwwmKSC0AVIo5TzgXeu3/hWTy6odSpYspa/w6Aj
1HrzQnWwZkdzb7k+ppQt04CVzlyq7KerHmNfZWyHjPuP4Knbw7n5nBNiB3AOb5A5
HX4xILnuM2lx9hUFsmFk++hNOuh+iTTMAKnovxT040wAh+u/0PTw0omrRQzVDply
YteseI0Eh4keENWWVSsn0Js2xlvvoP86Hl/LaozFdKq2XzCSNo8dDGWliSAJoKhF
9lJnXxU4A/rWXt4OnSnV9ZDGpHc/W4mhej8aWXyDbVdE8n1lR4F5436UC7+WzcJI
wXXeiulwXQ/gF++rxWJVfOZZhABPpUvyQy5NCsrk1QU+PHM2X3DjL1qV+K9DxtzL
lXAa+1X8x8PQujuHIG0vkpfHAnXUAqOf7bp1SS77O2H2HJXnwYk0Q6qScRd3z4SC
owaoQ2ERllantyxekUa233i+QcXQmF0F9fXZqCe2TAH3OGg0BbfWBApBB50XeIFu
lHezRWBPJsfxiqBRCCKPbsGWh3xogC424hYrzC7NY5wpHWCrJ2VVJrNVgjR98lh9
Xbl/Q0h0/H61Xjezw+0l1WsZLzzxrDwV5ZSDHpGUE6N8Ml8j5Y8y9O/h5aZtXM8H
u4a9MQ+4fkx66RIIFUSrP9QqXoUqKEd6DwP5xNTEyg5ylIlFrX9fnNp7F9D31JLU
WPSclrVe4eVNsEhCEY/ea/ygN3J4roXBLsTZcxe4DXVIRf1FBrI8ADNU9OpR4CFY
gQTBfHRcIM9rVBQe1gC6/M8rZqFRukF8xSLHK0MpEVNYaH8FkFBBzVYNwiFQPZ1H
4x7sy2knB8/csU/VFpQTdXX4curVJMoDtKU77YaqXAn4eHqDVBR0lFkskBqqYLcT
h0IyMT4VrUHruqdIcn/nb+NKVyOBrEjH0g9KKqgCQcnBmpySA86xqMgqftJHN2vE
qHkqgI7SIxr1b4lqJBoNc0nD+wLBRsPvDV5pfFC/2tVrZ/bYtRWm7gCyE4NYoCTu
H+Njdkfs2NfRDCLkepcGirTma7kp/Q7s3MUM16pwuv1rNLD4bfyLU8aVDXDm35df
CLMod4yrMFSiGpOj4v+Uk1PRPEOgDY1Kp4YT/ftrlbOhMceac6EyjcWqUVFtxZFP
hziJixy8IXLmCpXxY5sKHjdtmm/oEjcVKeTqA9ocvMYJfDx8Pr01Qv7ex2WDZpRj
UNgHN7bGXrAEWl5t6RLV4dslRiMnFkpIHKFKVLGsRtgiSoJWmdbelBS1h4T/rRY/
m+D1L7gc5mfYrC85Mh/+TAW4/LbfZ/d3O0MZ7OFS1ZcFnDR6vTLcUR0WLI/JWN9S
EIAuMXX3m8Rq3BU7u4et3vUniT7QrvgRxzSrd5Qff/8RydFkpBJGxDG0wGgckAy1
1/qy/i5QxNiZxR4Z/7Mmk3rBbrYGSEyZrdFtM+oKc6DXp73YOFPLZCmk451ddblJ
hX6TPLWoiAXaAM/GGG9u1cwjJF4v+k8vpeFTXYn6X5eBkzdaUCZKoOhjj1K+U+lM
/qdKWCTcx5Mp4zlyNx1T6SQPHtVmhQ3oXyhQ5KgDt8LXPS8V5Exz4+u7/5eo6LkH
FpDTugkiJ6/xm5BLkOTZmZeCI00z1b8DJfYDKJmRiuG3gAb8k2J3LsJ3o3iilH27
4jauiUgmRvVY7eYlN3t57iKTLPbZ2Pze1cvRusME+Ig+NgFMV7dF4VKKvSumC+P/
UtN3IFy6jVk0tcwS8G9iU5WJ2w5NU0HLwLASLEUcq7FN3RmxXIXO/vjgpL22uwe8
J50g5f2eYvrjfn9fawY/wqm6SUhLKkixvcQ7D+PCbh0N/UyDnv519S/cxnjHm4U/
pKRZZvlpvyVLvHn6q1AlLY21OWcAZVIqmb5yoMzCSdVZrXxiHN29EvTSSAbY7DXQ
9STF0D8xgeVd0489C81F3v4GMCim9/ra8La+sRdEy9Z7hAqGdxVENx10jAA/fVdl
3qRkoKgdjH3cMOUrEuER6eRqUH772i0qb2lowvE40qAmB/Gmzt62B1iJq0kAFcM9
+vOEUYo4yr1uQ9YMdK50tFlRo3zoREQAlSRRgrstHkooP9nMVGtSTs2USy9KARNv
jwYwmrt+fISA08yo0DMIgqcejb3VNGNo2PvXQ58Ql0n7YSjApNqf/HiVhjLLogpj
f8aSA2mzFfoBIKiIU5i4dh9/ZJUyu9E462iUXFhSi2Coe1DPENyhBmoDCIdwDvbr
0PsSo7xoVJj6HCG7/xnPLBLP+QIpMnsulTwinhHdPXiJQ5wRhMP1IsXPd11iKYpN
bjTr4hsJWytzPnIyIyZABf5nqVflF2KriuIjWY6wS0+6TXs5FRoKG/bivps4WQFI
N9sqtlI5RahmArqDEer5VFeYv1I1BfAsgapfljmL6omGIxWVM1hlQdYiUn/u6ta7
ubnUe2eIpbpeWBKvwh7eLxhPFTRyS2YVOBH9hdBeCxdjEFiAeueygzWdxDP6nH+r
8HZCQZdaAQBKDY0miU4Slmp0+X4SyveJKdlQOB9UxaR2rJbOctNOCaeb4EUezEgn
szcdqrOL9/VxdjlG9lKh+LDFGKfItYHCZ8fLlZunjVQUdZbM8B1U1fXKmMksqjTY
pf9Lf7dWK8TgrBAZRmvc/nrZrOXs6vSg15L12N67A3QiFmbhQ+x33CcOVA6BGse2
gV1yqMEo3ocC64ECNOZcediC7Zcf3EtZsAF2jl2nNwqnlYNldxFmya6+E5q/yJeW
rEiehh7pbyjILSOWWzS0EoTSx+D020kFBDk0BbjFo2KLu72PTAulfZl/+pqgEIGS
hGwIpU9ABrOSs/3bpRe1NGPdPdZ2oLc+oSWzEm9iZXXvHSB3ySFNr1sJGKfx8fn/
HjczFJjzTlfpdxul7vYGm4Dy83tJ4YtYWyauXtrMCcMZLZrWDp7Egn9YZlHUyAtm
4bWsZdMeFAuunJs16qAOhd+lMjzl6KpxeByeLY90FIoLG5RAmHdZDtGzhBWEW4ij
OiwDml/Kw0SVhHvxIaYu3rvKxdEuQmVKbPZ9fiRhFOb2pgjw7ef3cOBKtdc3HfA7
XYAnf3aowPCW/0ANCLBo/hCNO2hdwX3jxz37hjoNiYljlpBom2YAAobSufSpRdIq
k6rfdKra6XnWOaq6oCT+NyFxcO8ZpR4NTtSM/IVf8RtMQDsNSB5MRMrdWkFCc1QA
g2F+2IgUsppKr3vElBZGw0ndqHhUjqHFHfMX+OoFRap0qjJjaW9Rbo9L9E+tpEB7
S6fkvlgyQWH8Sdruj0UOsfB0cta1ZkEANGVmr8WisvoKp7ShIqaZNGtIHYMvIiL1
SyXXU3qBqQsLf6tcLY3/SrBCvVd9QPbvhYiNgWZjiaypRZpbTSQ2+dFge+9CJvX6
SlBSP9evUKSMYG52IAnCx4foQ1799+rTYhUBqqEAQtIClkBJVAV4RP6HCLKxs1/8
SiyYbOVX/50vWVXhN7moe1mYDR+C9I1eA6BIZRlZEy0nyXZXdnUl9GwN2uCeGML2
EKp62K7G9iIapclXJbof2Tfbwk0K2BMZI2qjBl6DGwylxgqTQiC5HNLMcYIK4E4P
ah1YiVnsl66eWTcdgZfMeVg/uf4+dyfjxgoxJ0ENIWEb94IByVSGJOOt4zrt/0mM
5bC9IsTV/TsbK8TBlcxGEwfhcJ9SRFbwXtWT4Crt5/KyxXanIH7D+7JGlxRx9axF
rKaiUhcQ1sDO7Gyt0SmEPHmryYGzVkpxb43PpJu4lRUUPOT4WW3aQ2xUzlnUgkr/
fX65qZHs3ZKn/Ld/HVLX8VFYG8ehfTXO2bS2lHc9wQwezScyN/IS87VCocZ+Vz8k
HYZ5tUF6QcfxmxTVQA1oPAm5sPi8CmcC5X4lpq532M/PfXBd8DOGzWWTiT3bnZWh
1L/VXx3O2YRUCTy9ZQ//c0P1ViLzyJXo3WFlgavkiGKRokwDzvF6bhMxIsgn1+Da
9yJlWQYyCa46Xttl4LrM0TqEA08EACN1ayPq1LwxWFr15YtgxnBUfGtPLiekArun
OfgmYQefo5UtwBaN8k4kC0InMXPAn9DjcLB418ImjYX1gNZoIEJYjqG9tj13aMOC
J75o5cBu/8Q14BaNKIuTEGe1r8SaK1xGQ7M/weVxOX+Muu9epQmRbzGDn8EQ1OsC
F5IoGcK7SGgevGfVA+iYMhNKbM1XWKIwY+wG9XKFLV4l9TV0023uOuOsmSrUq2Ku
9n62KUGXgY3V4WFgjAYaXCtWEt3ObLvV40yj/x4ENx+MRHlwTMnIOKbgFs6AY34h
hqDOgZG0q28VEcaKAAHTCbZEhBxgw+Suf1wV7N9P00icLhrrOHUcahTIiOBXiQIu
QrH0jhxNJh/bAheXE1Wit88n9RxEA89nRqTK87fTFmXYr3B6mOHAV7fnDf9n70D5
x3Gb/2KPMRzEQhPY279OHxZTyH+7reDbSvR5Mc/fKbWc5RB3c9JFbqU9JKKN+4qe
/nGi00BPltr80MAK5y+YYvf5Mc3hJkElyUDtAtLd2Ytpb0lh8lORRQm8t6p6fWEE
Hyjw/rz0YG17IrrBJHqujFZJ9EC+VIVEvxNpVxVRAWywQOw8R9yBUr64V8JoAOdQ
ngGZGSypjSYHkes4zbWfn70SJ5dG/Q36jQfn87UkDNbOD9xhCKaJTLbuq6erzjLL
FeqkBHLGuOYExh6KHDoNwJQAA+V2buVnymkn7TEZCYgkK2CZwq2CJT9KfWeceOWf
Rq/AVx3tkoCj5NET4BZasOtCu2byNHCyDq0xRtbVtTo4rAFxaxaGO8iN8KOQ3GkA
aOKfZnq45pRhb+RG2B3hMN1hy9n+MUK87ZAAey/peCW76Otv70Ish99meF6qI5iS
+7Jotrm1cD72xluOiokTT9RwipOfSePXrY0/zhI7QgrJVXETzaw5nWLG7tquhfh8
GvUbmdGtRxmVN8vL2/ehSJGsDpHmmoxZqrMGAlAeH/+WAkqmZvyazAcf12vtcIlH
9I05XJHPDFSe3zjcXmYhF1sk5alJV/0hDxWqCZtw8kXrmR4fjjCjRA6H3Xbvy8IK
CeNOEDcJufWSbRdnNJg/8j9ITeKRWBpFuLWPPet6AKe74V/Uht6KbkJY+8LETtYT
iEROm/btQfcDwXgvPM/N26/Ys5DgUNPu1WXVWw9xJjJVedL97roOx7m0DHfgHFoX
MAa08+sHoXKUfTr/e+ALrQOEGQRJtC6+yrLuGFUwqow5Nd43aiP/9mdO1OLi4Hg8
P53S6r0rWJAYWrc6DN9p/Ewv7+wyfWEWPM4Ws3GLczfAFO/Q+DaRgcWLOmPxfVo5
0YN2ig/Hs53x3eZ1+Op/KeFfgCr5BDZTQ5KuqgAi68Cfdvd+zbAj3k+7wY5jf4i/
rnxjEZ0Ba6ZrFDi8meQiGaqnzS1N+Yu7u+R6k7qsOFcaz8khN7Hx1nvFvWqnLQi7
WydXrzLyUfRC9HTMS88OujyPW/vSY6ObuONGBRxCzyg0+iYZOywAwpW35f7u9yu/
PjZr7nDt7qb1KpWRvBO+j+LGtVkGw74xQEar4CmWHP5Fn/ZJG2ue+EZJhTc97SeS
Fr2gxy9FlUA6XhbIOtuvKBGcAZWRtz+1MBQwRFZBJPYN0hN/dF2w+lGwCIpzwVrA
KSlhwoA1jR9kL8nxzHaH8Af07iZ9n/suUTend/ZLnAyM6aJY89EYkjhDyLzREGTu
xtMYJkXDGCf8EntBcvwULPDlSbgTYDgNkiI9q8sZAqsJ/ArYMMKKBeqQe271KUWX
8gtBzyCr8TKUIuLdLC5tNuLYMJiTANfEiseYZBUgIlOTz0CKECzzl4HRIEHq6lEN
hbr9y4kfZb3+w36dVcUj9j0Zcabbm8yB+rSHFTn5KhUan7XQcu80Q+13867XpBSU
3skVlh7vGYDxD6Ph7DiOt9zLrlKOntHD0pkUJjqi+9w0ZMda2Y6yz/3Bv3EvRuQA
vCZSU9rjgir4OZ3pvBuCixS4EBMIK1w89Yc7z0DgwsAYgyBNx05eHa/CETWgbChr
z0h7rdKT7mOoTdH0cHJ8zpvzu+J5eiEFFl7Dm1hD1Tef5TmvVLWpvfGaScLQ/rPl
LuJAMxaTpMUB5Tlm8NZEroo9ViE/2PfOwOERT22EV9OucdhK/2NXG3h259Nd0pcu
NuuR145s9FAzRNKKIKHfS64RLYjF1ASPHRUrui58tTvjVyFe25Btk48ZGBleLcTH
j2Q6pPNvs/HZz9GCvOZbRHBaTC4kQnhGu4Q6WUiNUFazT/ZslQJWaU7rPy2JQQ7T
9KyNLmgD67YMm8imDrzvmpuVGYBOgI8LURVL6tfrtmK+cOmm+FqAqt/T3ZEY9Mcp
OvkApJ2OuUARdWDn0vrnsM7yVpHZxbW01YEMVq1nyXMZ9oLMdXaTOcHaCrdpGIGJ
7XoEyWUUYBHp8gROYRQY1Q6Knf1ZI3UJe2ULWa5xdvmW/WwFLNpUdwHcwgYqnimU
9a1/5UB/s2AISPXFzhX8NcPJ0z71VF7ovv20zTIzSZK6bI+K9LAivnON8hnUE01X
cS4BwHEAqumQ6ZDZZ/j7AKPLo8JojCB+FgoVKDT8syXlYYx2OMpB50CutEZ0C3Si
gbCeV2Ja+nRYNV4tq94vTfGRxxPhIWONPrvRel3ryH54U185z7I0N58fUJZFQSfu
iY5GG9MXt5IGE5TsrGSqDeAe9MIVpLRlz0BaY9oOPRzQvQgbbuY/brhelxGOAcGS
X9HcSMifMe0/TTj/pCjSSHpgBH8SNM7BBKZcCgHU0Z0MSk3dAxkTdrtUkMSU1bni
XRI4URyLTQIBubEADBOJz3JM+3aU/tH622YPrYdqovDo4wk08v4W6ANjUjxKiSm4
qkU+ZM43E0XPyi+WYmuSqYrQD/fP+5KiU8w4CjcPdESItQfUNPvOYQp6GP6gvs5V
dRdlz0KrDkvjqDX+jmXqMcEjV5cTu2hP4c8xZlr8rBDac2ItyL5lgkZRYjNAnQ7N
MtTK6Jx1Q4GmKTUqMqWoNImMfpEK2IQU7r0W3MqGsR/lGbI5XVa8276tAcVkBhF7
kzZ137+Oz4r1vVdGxEiYDBlAnt/YHSde5JUN1mHeb9yRPD9ev2GysNG1d/tQVthM
pSxJstMtAYbfAJo7ZpYOR5r0mjk52TOmujCKxro18J+/ZHJhi6pHnMa5binBjz2R
0j3Mb7i1FlE+SBnm9FxAKxxr9kCBzby2wIAslDA0iBGONYfOcpUbspi4bddzOfNc
ZHxzC39KwITOeDjdfxpkOvhBfupGUf/j20Rr67B+T/FrmUSFPv4pzFEp3Peuts4d
ltvn2A8UFc41Eg6WLK9gULUfylb+7PVBxhAF5XsovLsRCC+O6Xc6Pdn/OY7TVcML
9bD91OEvFvH/OQusVI1AJ8SSY3hJoZRnGflbpcroPtL+6QNIaUPRR7luEMCUFg5r
LLTXlypAIsGGqcSfnw9criCKbCjSqjLMhIIQoVmL0/05uLEMvTUXSKYESRo/Jviw
WmvyKMbdh8g7Qc0HdMaqV/yirsBOazy/mj3zI493usI2xE0UmmDjOCH5hf90lqEk
XWLwcBW/8ZFbBmZdGV8De2fjjEwFRu4QXJkgM8Nb97uV7+6ZyoIIsvHaIn2BORfA
oKc+9QB9Eur9yohvUIl7lt3mvxhP+J4GADgWovUY2YXP/FmCt/UJ088xLEnc6zUt
jTD6pt4nGRcuTW+a/dyN6GAR5QQE7dbyXM2pM/bggsF+bbQp69HPi8dsghweszh9
ZMF2pK+nI6DCI0QRXuc1aa631tBtgEmhfKVFvZ/erZudiA9JMrUTOMVntzQ92Z60
34y+JvIaervchvmU6M3+/YP2VgalaQa8FT7Dh8dwn5XYViEZKqTFjmW93HqjJU/x
vuGkIYACPkVePaItSTcp7zYZWX1vjcab/dGGrJRQY92F9pAjF7tsTyyBmHB7zFHS
tVwLkSDeL/n+w+2KCk9B3WMbYYcvF9AK3m+25lXw9AZw4mj9pYmzUECA4PIWoZfL
tFR2bb0yOBstD4YaCXMJ38OHNi8u6Hmxda94VBGv8DWvywYBPiCTNgg0Qx48J8PM
A42na642q0Yl0PFwEdmUIofrApEi58CrFqkv3u72EiuU0/UnK/illlBTJZUEmUk6
6MoxBlJhe+cM6VH/SMcKgA/3oxCzIaFJbu8nFFhMx4xrMgiW8hUeaA5kr/znCxZE
K8p835jrj6Box7W0m2K/7nQP7SOJrwAg9ixUblJscBvJcwKRqRxqQCoT9KCJnhN/
W9eTkauhIOho0f63rrFJndssrSjMRW4/nJYYT0m+Lgi48b7ADMsHtdeosTDfhQ3V
jd5YEdlwHwbklV6vrTSUs/89nh3VZPH64+745l+11LYgwb7VnJJBFnyXrB1n9BFR
pkA1Hbg+5vXTkwcN+TPFzOCjbjjzEUgBg//jYFSqZuzsDehyz2Oqo7Lbk24jIRHl
KOw9W2uDClNMWUUxjaVAEs5FUxfgPtB0e45eFVht/KHExS7s5LnSmVo4AJkVM90K
AU7DxrUgp61J+3f4PqVDHhmYUVa98pf7AuXH5x6IE17Ok/6a3+wiaJY23BFAecqh
sqPz1RPxJ39iEVdLGCJ1aNDC+WhYiEFNQA4I3HAo/K2S6K/0XMqV883NezL5xQr7
YbnkY3WYmo7ncRf/SfLdtf2iDugXXB1OXqpTy7aSe9kzZvRMy6KjDDTMPoZhxGgE
BDp2aUA0m5k4aD8ijT99ezmNtpeZeCk/ecS8IB0qfz/bDd6SX+C8P0bl4MhCzxx1
hg/a8le/rNSOPYQrliD76IhxE676q3r95b8624/u5B5D26zTrhCKnzW/E9itmrH3
lzZm7UIZp9oKZa8tryg62k5S9tU9bJ5UTayhfa69IbdiAHGaLDtBsCtKX7YDvpeL
DAg11+lrgqSSQ1zH3m9DiZzmmYFmu1GPnKjn+LEGVonfemtfkKkTg3LiYQPknL5W
FZ5ETSgVCD79z1D1L68a+fN7FpVwVwi/FDqveTCITW5m7831zCux4D1XKwSMUZZ7
UnR+kYcZBWGmw5e5TAv8/gU29xHpgWDBbZf9LrDzTww9oblxSKw5X0pO0e/EoUwZ
rrK4nHU6HHPz7cV2kaSB9JEk2LtuN9r8bRdGEcRazgo820CfhUFswTOlu7PY30Kf
YHuqC2CvnqazrVpm+LXEvvWjEpJWPt3aLY24lUm2qjmBNCprxpQ8JXBulAzQDxfO
lKPnCvR7yabr15VDDkI2Yc6LM5ih2lwah93CtBtNOu69tvR90OkbE1+4oglOSYEe
PvkjoMWYgWjvrUNXadbvVdB3iA7Yv0XWrqivRwiHqPlxuYjSjyhDdiFioxFILmad
65Mi85ybHlrhO5cQE9MweWXqvttp+mNUvAVy1oSOLfgcOZ5IWcdpK5inL4XlYOVR
BZK/HjEK/0DjAXP6XSa3pZuZ3IaaBRTrISBMUd9VItHbujDlQ5qPvBMqZiy/MdTg
aASQsTeINNmdIg4QrE8lTK6rIRuAebsk3VlXbQYrdTyGxanbj9HS/XvcTExHdBC+
84rFiBCRLwNq8sptiOv8+xD9c9QwvCtFlbyuEMXq0FGZynO/orJJCTvLlys0Mm8Z
5qVzOp1nqcy2qUXAPLyFztIZRccxTIOKui7mShMeT1p/P1ahA079FnUVNakocAP/
1lLJc/u/HV3ScCXLsQnrGd1+9BuuYCBgO1Uf6V5DMUutj3ppuRCN9Cfp8m0JxHkO
0c9H6KXYfMW5AJO/IBNN6aZlEdGUZnWZMOxo4CkOr+9kxHa96yrw2GgBcE33BV0h
HXqbL7kuG5rhFe3xWC3x/YR4tuOurRTC12PVhoYDqzVb+y9V3Va8nQ4Og1EF7NLQ
JsafKwYz0YmgzQqrTvEllbkukPANw3RydgwaPQWWPneUYM3a5ET9yuxeuuVZdd8R
0vPG327H/vT/Uh05HGXTd+1ByFqFHYT3NwPmFSKCaAr4gk+LxrYfA7bheidXpXk/
EJpJnOiCVQYOeAPS6wtDXeIbmtvfC0J+c6gAS3wrm5tKw/7Ktfh4bizhBdypAZqt
38U3EOFpNZQqI1c+3w8ULO0AlnCJst0eg3Kf/m47fGrKkFnHgKjUpvGIUN53Ahoq
WcyAPZ3VTyCpjGasKfxhmSzYchepeWdzz3GJtN/csTpcQYNhFSVX6MYPmadAQFHl
4SI1mOsazvVqdggsT3ucVVZEMLeqQQJm7BPTrhZIowiuZ/cGR7uwNf5ElxppFx8z
Z8XezXY2hQgKficG6O8HTHOpLRqHIvbZ14BT/jKMqhTEx7aTtAS+y9wLChamrQis
atslB/KhOEgmpXKF6cRb301tt3lRD9uoWm2prNczQTM5M9cDoRyBzpFtEiLLWpLH
8wMaPDLVHv4019L8aNnqeaAEW0qhYYnIB3YgSSqnK4HXK9JQZdIwsBSOJUruoFxJ
AAWuYJ5VXlruUKSBbQyQQkkl/qlN3rPPvtoNUQiw/h3aZ/yLSROkIomCDoF4sbgM
nAKUFRJSKyxHXo+nosLOZCSzVk8XOzDBcBnX/dwwAwdhvejRqGQsIj3/xlZ9huct
yXTHYEXU7Kfxm9up0TYhQ7z7enwDyMi8/v3GpFmdMwF4RpIYKzdo5DlNVxkUenJO
SKIwFmKirm/ux5HnYsWcjCk+rx+li1Bcr5DBhkcfRL0SjB1KZcmco8HKbLN6WKYH
Qq2kTuzVy+VX2Z5xd8ADoH8NMr/Ay+hSJs9szP8c5xN/XQhUh+j4DhdVajJX9SUt
aEJTlfAWYwkHHTI3HehzT+FCwJy1RUZxoP9faONbFqHMbx9sl/pNEpaOJH5mwNfR
AMt/mhKZWMngJBrgC05lCJ/Q875dwofa6e4IZiGOp8B/W05gu9avaYPozinLQrut
7KYFoLTgm9PkeK2KkziXXAxp3F6TlDh1Ao3/mhrMeAN84QxnQmuPoDjonEqa/fmm
s0FYL0TWqYhMM603R7imTo7SN/udauiA8yVULcrj6jOlI1NF1fxIRZqeHXhwoNPB
rCszSospFDul00/gWiF/WiLJ2l+lKSRUmjQJwZyCNa28OcnPR+lsNIzmYW7BQ4VB
Ho0tmyQlM65ZyPSZTfuJD9tOCY7aaY3AsrDKdAYioxiQjsf9iCiOmOk2tZ57dGQp
kdS0vuRSqUpqK3hbVcIbhqNEzANfQPce15X3B/TUfmBUSpeycj2jZmprd9UGXNTS
lubN33Pyoe8gV+uQsDmZ390XSkxNAjlKU/KBoiFMaepn/Kn8KTUIvCMbpOz888iZ
q46H8+9p2sM5RuJketFUCOJul30BUjhDMhByjSczFrNW1bJRwvxAHYZLnrlDpULx
ZdVA4oZyIPrgrvHjKw4wDcAybwCR9SsVyR8Ci4eJhy6xi1yGIO1rStsF78O46S/x
fCNvr+3wOhLB/Jewf37G/LzlIfP2CFq3qburkHsya2KSNwBeBYcIQjYSdmHK5QJ7
u/fv0CD1RkHevZ0XnoSLDiC8zh+R+LBCmBjg/1IJAROFF69gUCl0/2Y/YkrQhvUe
U05xu3w0WXPhopLyWemC6ThmqAIwEyoaSavyQpgFaKXQ0jsrRdpRBEWvWPOx80UY
IC3zFOZoqRcEO9/QztdN6ds1n5d062rohZg0X6T3XLaKCO3z71UGyLne2apvzmBY
Wja2Om5Pf1AxpmjjTQWdKHuOj3471TI7wn8OlhoJSgev+K8tiUuni6g+dPrOa5sU
BEq3ezma75TDEDrQc2fmuBGuFCSbg041Dh9kkI0oQMGMOe6zafZDQ9epZLYSxzZJ
mksFBPV2jXiXKIOb2dL+p3S++ALUpiJKvwTk8B9JMh0KE4fuMNABzcPWTRQ/yNz1
mjXo6L5mUH5XK0+MYdiF4cleMTqc5qU6jrqx6wTwOtJF3rv+QCdcBzEyyzcDLa+k
nhXkVecivKEA+/rj56FSlKU8u7wwjEZrac8Ea6fv17ZPukyC3dYqNwCOdIfuN1Ef
M3nzroqQmp8ejPkRKsBo6J11QQw+wtGO1+6wObWpfIZJ/Pe8rDIFAAYDWQRAHwaB
2sfoN2RidA2DMrppcEoax+oML82doIXOULvP5u1pJcH8NarogdAPikGiLQiI3eOi
FQtag0pKHWx0r9GGJ47jp8cayRZta1wKWvdKt8+ELE+uvJIBHmEKRrJl5STyqd/c
QdNcg9Hdzf80ayFbKGmSmJoNskVSQS6vaT1Zr4XoFxf9wbSd8Gj7gsQWGNC9+DPv
ZSc+zapCia4ZoATedLiJ/4STvuWxkFkqRaN4Xw6Xso8IhuX9lZmrDPIPlTj1C3E7
stFVrISic2yfY6qQwJ7zrFK7qx7LI+79kwaK/9dz0qte2qoiNBnUKvtXRziuWYbe
jfz4xdzDighvEBOqG7UjnB2ReiGlX74UBwq+xmDEOH95ls+nnfvess0ImSkN6R27
UqTGoz6lfkgq1Lr5RvvOtXAU/Fe6MJIghy8lGVIsGNvbuXd39+073pwFI1vCXOdK
PhLShlnWkXfogxMqaXdemmNOwBne9a9HJ59jDotOYjyFa6BvzrBZyJHsurYA/x8S
SURfJ9rrpXWLaUXE8Y2ljJPw7UDPEHqYCkhZuW/rwKjtB1NegoWjU9j1FlIk/lDL
i8Lv0F1tZTQeqrL81TBhQOLLSKaKPwOFGExitJMMeuM7GwDWWlJweb9QoikgMLFy
HAnbljbL/B9VlrrFMesfk5SrIujhEyQG+NOwUdFqSb/Sc2lIlTmGa62bT8dO/jaq
58XgK7695/nQOfZv145zDZa5EVrtEOFYnpVuenNAbrg/hEwuAeM+r1Xfs8PveXJh
eEpavA5u3kur7J4GbutmZINMViPvZ4Dw4sfr+g7CZi4jX6xEuhfsDsNUyoHPPsUU
D8schiir0eHeYh+Doehheb6EEGvl38RxMzS4JW5Psn5IrZJzUeXnLxQZHRqEeTvm
KO/mQdgo3KuuW+JNyUsB0Ayps3PP9NRmyPJjAW+wwff+vC2QLAkhZDtUoGIH1WxS
SMjeMiysuiUDYN35jCIDihh5bPGhBtniWBsOvvbNdWw7EhFwSiwSbOmKnpDMlhcH
lCl46rGoewQW2mRJG/XQDDCuCyBPYNDiwPpdsGCcgA38WiqQTl8nrx2VOQj9O97x
nS1DcacZmRzkkn6ccxV2vdrfhoPUz/VheErcCttbYEgsoOEiiRFXGLl/CvUy7iQE
fN8chmq89zndNDQcXU0RhE0WadGkdiKhGZsf/CvRLtiC0G85eji2K7P4+fkjCA1x
VMQEBZkhwfGU45YEQq5u+xvrJh2Rkzh7sT5Cb5bU98QXyPNIxEee3TP6zSBeDGMW
SQyA5U0P8Pcb+PjjSqueCIoCajF25OV6v53St35AOtnyiaAmQU6ZnHfnzhBUeqcs
sbFJ3OM+OBc2gDx9e2+FVcx2k3iAQbEKjKe4QJgfm6cBamupfQzJprhMf9BXjXPe
MtUPkCvlx9ZfjEKN/tYnuk83DZZES73/Ue9Aygpb/CdGXWG2qY0mL9asH1w961/j
SnsEhZ07PCVDWU9PAgVq2vP8jCgMIeBnlwUXP8s2Hh2QMScaAz9Ytoglsh9PWp1L
14cg7BWWRb+BAkbDvabyFZiQAHrRdAW7M2nyGFEqh1WWUC6u9vFoG0guqpZlk5EW
Xa6wTsPwDETA5kSzptM9m0NIfmEIuK+2RKSJoTY/9QJFGQ46oTVVl7JS7a3ToXOy
WdUosJCG2Rvwe2sXRGD82DvRzY/g37bFK1itvJkJkX07J2GaD5iEBkoKaKi9956W
7K2U+9XnrA7pyDvEjQNflaK5ZaNp7B4qaQ+IeOngIchP+Kl2d0kFml7IqrtvnlRt
R2kMLCvDIJ2FtjCQG6tcsIe25CNKuaoaaf9D99GuFpdM5yYueWGwsYNhAtSkCkYi
8NXxMgri/hNmzoIp9eWdmFyp56sgnCW1Pqsmmpu/o4328Zo5YlZ2lMBt012I5bkC
RGy6GaP2ur5wYL1zBiXyQR+Gu4C0J6dUVuunPRS6mCTx32VA4/CiolLkM6O4hPVY
Hpgwxzuy0+GLfwNNcrUZh2yJIDAqvWv4++qGD6OGfT+d90kLiFbab0zzsaOrGrp2
D4vAxjBzJsf6ux3zYUhHs/QNL2AYTj4A4zzTrf4LNgCip5JZOvdl/ZJG0fSjw1zg
KhqQZd8fUcGjboLa3FGgHGCCzjwCBhZnLGpEgdGw5/aivlMrjPCYI0Y8bACgVLnd
XwbH7pBK5/StxjXE8aNhpGWWtWpMrMT09RpBzoynhGgEljqGLCMQuV7bpL4PezcS
OCBr/Ysu6XoZXBYRka7L1sZSTD3NRzatyJ4VxbmTxfTPXFcCsPFMkvftwD5578/O
vhf121yIoBT53JB/tN1N88wNjoT87+PYWsbqj47liL5Lc4VV/9mX3hGGB13593x/
5O6FcIPkpJrov18pFGqTmVUUwrbqcU+povmgfJiP08B87dq7/Z7eEkVdSvT+8/Or
Wk7JiD/t+DMcOlNaM1J4LO2lep70uBj8XuoyxJmJO9I+/DGd5RxQ6lwSLnHqaihx
fStOpDI7C6w49V99n9qYhXdTIZrcRs5saa2LDmc26lIWAJE5gMVcWz7zteSiTM/I
SIG6yLh29ka+bm5k4NNcygHPSERoXBv4QQNy8mCNwBXBAsXI29NUHMpK7h+WGPki
doNOSufg3balQq0mZe/H93HDBc1hX/RP1tX/3/FaIBTBuyrtZbMuL8tHEk+9fsA8
KYm6D0BIy3OG8h8Sy5o6sq2Xuc+1wHGmix19VC8SY8ss5wfDDqbGGuYH+Myx5oSK
9sL+33UliAlqDztJb2VbMzSGvlvLzSbh76wgHp30szVDWG1BpLbyBx/mmICO4OWz
N3VA7FIS9uPeqLkbmcxOmXmHE5OdIao0ZCy/TaW9l8KdN2uI+UcmGa78NFNOWuXK
Njv7xshoHLyDmjAeEMO3QvhwBpUeValdJs8tbRLo9zXe1OIQ7Jhh57VCobkpV/KZ
98ESxwbykFloss6XRvVAu3SFuJEFabGLxlHs9S2hl+X5+4Q8t4/Dap74nhr/It7U
b3nUqsjo02W5jRXxv07QdbLIWVsTA94GOta9zur7YuDMj/ge61wmevHBr1RHBpok
o6rsI7vnG9sLe2xQKwrN8rpy7P4IfznQyei9pE5gR7uM05aE8z3s3hY+7GRM3DBh
WB37CKXF0nnIC2vWFyW0q21iWr+75ryAHV4f8ZMewSobBFGHYifLhkVurdyqqdoK
oZ4oiv1MzS+JW1jiGiNDSZVQNRZ86eOOZGaH9CH8eRp33OaEr0c3j3qC0hjCWtTM
UhzjSFRcVeRTdeLvNLpFmkh/5q7eKzfcDw06Iwf4yyDuGelxPpHH2oInO8g6mJh/
jMY7K3T6JnvQop45ObioRWuoIcph68ceB8rYN4vQdownO+hh+0MH4eSkS9rWpsN6
B4QseZ85ZYsVfrkMMvU+Dol1HsSn673YUEp72p6o5pRORnydBfss+bMiKRHpTgI2
I8jBCPxxFSbvDdykPGjD9A9IrZHMrbuPniih5g8W5HPeKerFsW9zMhEtascavBCG
Tll6dkQO2cbkvyPy0FAne8I4zEwSa1nza9T5+SdbA0QLadssMShVvlk2WCb0x2Hy
q/tbHz8ROvOSDotwrLqoeE+3BkxWqx8dU8UWQj2OurEyB9UJEg6vFouqrieiSgjX
luZHPm1JF+sA5qy3N1C6HblGlxOj9YOvFrubmHO4LRCfj6lOlAs2EcHCzdlQN2Yy
xQs33lZxkkEMLcQWauQqtWFeSs29s+oCrJeuSkCz4z8oqeKi6vp7kUj9vfzhm3LV
eFEhH8WsNrxGaIllFYziUaBkATrVqe/ukgFvXeCmvCVzzNYRXxyn6t0m3WaYbB8B
zlHVPBpDeMEqM8025wO7ffn7KTyotiR3QX0wRCltq9hfqVYv+ieHI8v2UTD9Fklc
1yuro2/5HNHAvafQhHkUqUD2a3bB+n3785G83YrPFItu1/x2ZEOSLSw+zEoO8V3j
GzRlleQhy6X1X58MUQjxCcyDUu7/kzP5Sr60t893EU6RC+BTeHyOdOXTprq8EcJ5
VU05nCHrSwfqfE1XMHv6Cc7s3GetRBoQo4KCR77xXZ9a4a2aPbx6BbiYzcM2Kr7v
gXPcURRjrRzk5F0EICEwPMwZL/uKd3J1H5Y4YPFmCkqYpesgsnu8Q+0mGG7pzNIU
VZUHw1xHt4H05+XV0QtO0nejqy2LAk/wurxZE4zqqYi9Rqo0szoMNasb/rHGqcGH
VXfrLWXg33tegOT1edq9t9ydA9QZFMAYGVOnTgd6byiLTPnpH47la/M4gim3KVqn
q/noH1BqZ5vkhVP/KdUE6FdwRZMEL//riYR4SSu+kF50aiapLWLGorqcPQwElwgp
fp6LnxLQwZTj2qksAdcpw8BkONa3VtZDaDPFTzZmuw4Cp4sbEKV5CEI0Baa8wVFX
rF7MIm8xC67WxKMLxRIZEZZdkz/wvJ8A+m2Y6mOoU8se+X/PwE03ci1Hu2I8YB63
ClVNOKCoQ/97H+Q3x17/uOOEolRZj1MBMAIa8rpJNS1VtsFDvlOVKcTVlANibghU
WA8cJP3rcEup25bQLeX+aIpaEOfQgWF23dzz0dXwbuyKGEQjaSX3d/kSCo1zkFx1
wH5jlvWRuH9Q4O+1KY5kHq4EuhIy6LvMB01C+FVuioTslqtTlLiFygtb2Z/ipdAc
iSuM0qzjS1AIhYq1IKQyp/yfPkNtBRVSbVD0lYmevn64vI5seYn7pwzch43Knv1+
yEF0rWCLGpfjDTY/1+wP6buCiErFWLMc7e0Pizd39DSkMaOZ0qzWjTIqbNM7K7V2
usQTiZMZgOyqShvktYkxXxlnhiTVC0BsDhPF79yT2AT8alU+LHjewrk9StcRudyW
HzG75AnHI14moC+TwciNXssD5JsXgZM4bdMA+sCZuZarmpKfNHV5zdBaBzo1lEwh
BaWtQRwb6ix75h8kQhAcOksJGtVGFFjf42AupePi920pQBaN3OwD13tyP6kcQ2PB
/DKeSTFfDPOPn4t3m+w2G7RzlkfBF9+TexE68PKEqCZkL3jGLME9S3tLd8ybWbyV
0Bxh8uR1Or4G/uimTlvDN4FOJiz2z4gfUzac/p8/JxqdfjfiKXYZv2SPqEhi5NSa
q3XmUqW5sp+Sfhujd4Jvirfm5+qc7zY/XJxoMEffr1UlkRrJT2KUrsjX1GwZZv9m
JAZ0l9FABgoW11ORQwe28s0feWZVSqqq6CC7SmR0R/OxligySH9fxsRi0ePqkN/x
nwqKFp9ZuPSWiDW8LIxX+OSaMLfxYePSWIxCECT2yJ3o3DCvZSEueBBmZu9kPwMl
bSBkDK38uiLZLkrpA6eHrPlj/Ms9AeDkz6B7mbu/3icBf9tRgIHyNd4ki+Ve/bo9
SWqdTFr/C7nczxEIC0+KmDu1kLwbsHqClEfmOSGtxMMpZpTcWucFDp1pUcTTensi
FZNYuL3A0R8m52aI87r7FDr2hTkh5aUGWAdKI6qIZBYOvVTUpgo4IoC3HwCQnOAH
LBrhrGINOh2LMMgCVFhKIf3f189whvL0Jk6g9QocVhZtcddSPfb0X0orQbNeRRGg
WEmA4xWXC7gypgK8d43qgJOt+CyWlqcn8MMV8MbC2Jf7kqzAkoNOAb89zbQ1Ru77
zI9TAAFZ0cHHkceBKkoxTEaFNGHQNVPzka5QvLb/dM4Nj37Jt+3MS6QxL1AaOXV9
edTx+OnxS13dNlfOmW4a6UtQi6kaKo1rSrtxKB5zveMiZADptPrqa2juFNkbSS2I
dIN0VmJiWuEpdPk3ys2CBG4WyR1Vp5lkkBgoJ6BMg+REQN0SlBXRnm6/fVXmCGGR
+mZpdBcGJEz5X959n/q2Murv+IHlh4iIzDZ7ObpSKTrWvViYRk9YvBXsROMuWpaG
rC7cA8m+pIJADOwA0U7qXk1sKBTbWlvPCVoFSKkbADBAuN14HMwDtIpsCNMpbPmH
bJc+NY6UAP3+njf3fmfD15LaR0aSJfyYO0StNp3g6jHqTHYgRua+jo7T6REnChPv
b83tmtIAnuDrzAkTh90g+oxGIeWrRFD6FH9WjxCzY6M7HK4r/KRT+1Wre1r8Ehuh
8lS7lLzqqThEt+KknoB+0yhQm8izkGfv4gC8QeRDXn+t+yvDSqXLPxPHcsG9yFg+
pwgt4kxas0WE+9RjqsPyhU5IRm0GY/7StUSlX0ZyJ5EQuut4FU41b5j/JAqE/FOH
MJmbQeoAYidD1N6qC/QM2ytRJMV1knpbwx500wiq5JiR/CFGmr1GwGIjMe9BJ1qt
4/KJjPzLtY5QC1WKBowS2y4aLWrzVYVLj0L2YaRSgXU3BqBKHBgBDK6TEromkepN
uuKiTpH8Z7nUKa5vtWqvGrWITE6Q4EC/gSiVnPNP9jGHKjaa/229YQE++idcvRDZ
JolGuMgH5sDZ3Q2MbxQfHsTNsjIAMX1SlnmDHOWp0RsVicCc62L6wblJ3I8EVQFo
J0zBlj7yvpYajgMZ+fnNnMa8KeC1vgAbbPi4670W+K1G47ua8Nq7hGjrPNGJpdZB
HwbY7M+Ynyy7CgcqFu0h4/tj2zqwwqOfnsmiC7oFGkMrxsNB8AXIWoHa9TjYHH0G
v8NA6nHMhSBTFKu/FrwBZtdglxt9Al1PfGW6aJT733TH+Jlp32ugcN15+FwHzvzS
iDa6qQ9JbCsJpAs+8Je6ZQussvyOtbRdR81Dbi9L0GmnkQHqHSFKJ3yXWnMuddUf
GV60lKcJ5T+aQhPrqVPjMDdJ4AOn2blce2tIfiJrfj0mu/PBr0SzPYuj1jS1DjpM
N5luu/m2E+oHvGbmPIJTCjtGKKDn5RiPSsaKUdStbNnh5455nWcMdEkzXYi2dGsh
2B4rAm67+w/KIxXHOwYQUFQoMwA4IqAmxbM22dp+U+VlLTesEXqH8m84KtBn+3Rj
qQCOrssUemTaQiL6XPjgqzp5QfGxJSlhSJ+LiUOfJQwTiTxMIXm+1yfgA92y7KmV
qRRsVnllp76VmgSeqOuLBEhfJK+RnS2UN5d1T9xS/zFl+n7KRDFdQsIS5EpvgXUI
5Hgf1n55yuGjmvVzEK58QK/utkDBNDpit5mg8MB2tJP9GSqgYYP+zJxxpjDyYBiW
kVtaLg2pF8Ce3f1P4VIvndGccL68q5bzNtIpayMSLWyTXb4v9My1NiIWb/3+C5u6
lcj7PyIsoDNihqYibo/Fff9cXFicr1RaTUvKuGFXVfnzNJU4Mm8cC7HUExq/YBdQ
yzmtRFVMAeiQPG9f7KKq83NtwZna5hpihVsZKyX9VtOXjpsOKop+pGgEvlRJT2J8
ZE8UGDLCrHfRGHNPK//sUL746qpGVWxsOg9cRiIkZbSk6rhjddDoR948eO0ihvvO
XXgZfmIhfUc/lxBJs9r3obcnofYqBN/j6GiLZ/wzN2ODsIqWURXEP04N3F+SESGS
zElT5nnOnnN0Ulu4ZmiR1p+h1M1JnivOHxwzrMZXLxl8yWeX9EG5EBz0htMRmu1M
m381k0Nv0FsTJxSTgXRmX0NErPGEKWbBex39CB7EzY7Ty4abCAvEnSHvXax+tyk/
WN0SXs4zuWf7WgQXFAfkDRHTZ0sg+B7dLsPe1H3SXezxZ38b65tykR7v5nCTcwdK
ZJ8CsbDt5rBsyUVcdgG3tdRCzQSw6hFEWlXyNc+0moCSAmmu17mNr5IEAbbXQ3Ax
mbH/30k5Jcyc6TDY7jQDqItTx4RwF8lqC0xJtPHuq4rYZOkgXlJQ+pHIqq37R7Mc
Ig4U00vkWQyKfY8lqfM6p750Kj6v30U8UXG2KpZAr5LTC7XoScC7Jj2zh5/F8Rh0
Z+3F/l984Br8zTTkD8A/7dogHho3UEZhiLpr0z7bt/TjyhPLctMVASbCyFrCuEnP
/Su56NXibdDdq34OzyDz29ArGqpXo0FeAHBJpCWuZVU74vJryK4gkflY/nZ9vLEg
w6N4GkyBQOfgd49b4cJl6UVrHeDaJZgr2LDRzzBAO1VzXKmou92lMoX3EiYBbGwN
PBLSDQ9oZ1AS6paQgEvLWp0gQZyuZgklDrXI0+EOSVmN90KEK2CM+Lu32Hy8UZ0z
YzoJZMGhNSTGzK02QDJjR6ub+RlJ4rmt/aiKj5z63CBsht34O850sbo6rlamq+Qd
8kc0ne1eFQQcM4fz9nft/M3+/wWsGWXUZcDROnVs+gqhuahLz8OnBOnyVxGombQy
QrFgCZvoa+pY9eA1vJdnzeqcG/vwNOxwJEKLGvOTlXD8f+ANLOsXZQKyR1QZqR8S
rwdl1kergflOJ/1QM5D25cPYb0kjOsa+jvI3wjG5EKibqyHdTsEKCm8qqIHyUr4y
+0L5MhzkHagH0mdEb4EORFtKpn0kkIVtfnUVNs3WJmb8OB7souUZ+ri4jbFC90Vh
gKUP0/18Jtznr5oJV/7L1mJidtcrsjESpEspYBxq9UlKt+V2dJDx5eU061p1DzOB
enNtws8psdhiKDRHtPF/H5THQeC2JfZg/cRp3PEV1JtbPVGZci12vCbIIEWyse4A
uMW5/d0fwqaSQIeKhon2iydhk+221uekbcRquR2R9dC8SvGou4rtwg02WZcOEB8E
xXgEn6VNF9xpDfimbtR/NEb+TC4kQIywAaamH74JmeYrmTLXcQIuFi94+p7Owobm
CqsDRQKnaT0t/AQywmJTU2qTY+kxXAr0X73xN79dcliQ9dWRK3ZpkGbQHaV67Z4v
hby7dRJ4iIAVRAOm3Y6FC3iJKiEyv9YXZkf5+tWSUkWuv/o1TQxzyeV9UgbkISw4
rFiJO2ccP+gGxQPeN1hHTVqEFPN1BXUJJTQ06l2sm/Ut0oXtTpQS3NJ7k9GyxG2v
NBr7fjhchcpjEGFdqIjNR5v/A1uPPU6s26Rl4QOLbDPPe+ugHw3T9suMfw2ZE322
KZRuwKhS0dxHpTs0sOWSc/17dDp4kdOmA/+ZUjCgGCAvBQKLP8WkIvmG+iMUapiv
S+EOAWHZNfi59Kbe5QFGenkbijDcyraexN3JFp4/NxzNvk/hc3I5Oe1ewv3cMdB1
gfmEo3aca9g/1s/246PNBVsLR1rQx8lKU//IOl2D3aYBZfG7AsCWws2NkPzdCpTu
ZcMiq8EeDvUQfjDYVDFPInbn8CBYkU6wxviyK1eSaTb8bBDHGqzX5livUETIXp9p
xragHMyxgVmNs00BaZ1KSKmcBnFuo21K6KNn93ihFOairdF87rl0AWJrxSmTH6mk
Zu5c0zUau6L06RcgE8F+MnfZ1NfGi1Wl50E+mBQfXUyowyvKzNdRcOCOK0am9rA+
+/H9Re5qKxF1uPc/R34B+wBSVPSxdej4Ywky1sRHTiLuhrw9QcwOJKh6GKRYPt5P
yVEOBlloKMaR1JE3Pd6ObAYXAeriP+ODs+GSyoheibG7cINo0REBL0NWehStZxcN
oH5shPiISNb1JhZpY17vr+axoFy/oYIRkgMxkeUl6/a5oyL0dhiRzf1bbxDOobWw
scgs4cyzq/MvBqm0m0U6YsSvve+UoAbo9FIfohKm/TckNhkBighYzjbigllAs7RG
ks3otWr2txlHzUYjl/rMfUgf8G0xJ4htk+RnDfeBm3479J3ycas/viCxy5BkZpJr
lLfIqtdYxB1RL3dIMmtYWq5+NB7C9JTjuBblfyhFMkLJudTd2dv3AMJAscJmV0HN
yNm1Ofjy2+r15vL8R/wZ0gUF/R2iPsc9TP4ac/dtrUBeTdboum8MgeLzdXNR1bDj
NlB8+MDBSSSq42SIAjzBzQwMQBof+Ut4VMOEw4Vu6U6T/vBGhus5rFk0x2btt0pr
4oSBrxGhPdm0qImnW0omSWBHr1Tqtzui1ygKM/Gfwot2MmZdHEBdt8QtP/HRLIpP
WMUB2+7oq9ArdGpeKiXU+ccz+f5E1cLcw8jpwEXHX1vzIsIf8+ri/QmOHQTKTtBD
KoQ3NkUFjrPwJU0vPWqs5mMRXKQZD0gzlSa9RvpU+VrcTHu7ajOkkkm82U64wK8g
+eCCQFv8tQc9U8nZCIir7KH26MLQzILkLvKkrolCIli+c0qNQdj09WHl3i/e73F3
LGD9PTIVSAnmmgjXsRMbQ5D9MmziBxQVFFLdA3Bhlm82ur7wdGMdygAHxa865HZo
FuuME3Yg49fnIVck6OHCopulPlcmGgU2u5dpb2XTOGnQBXyLgXTHYx2hG4jT7LH/
iRqHEYJ3ua3e7EHQN+5tRPHkoN4HuFsXGec26i+m+v32IcLxpD9td+kferc5mU6s
IZziQ0s/J4KhVGCL1GVpkosgmFOe3mXH6WmsRuzn9rbm/duHM4ujFRWAx7gbGDz0
MXye7Wh+xsq7mUi1kKIVEaMCVqWvK1lXmsFg/IlUZig2MqlPypJNmwt6BQljy8Tq
lv1Wt0LPOwSDNV46brM6YK0EvUHappB7MuUfD3w5m8hoZnoSMY1ATqxI1P2AB4VZ
YKMdNiNIG0NZHCtsZfeFEjyvK1pA/0MnH/pe8v3Exls2XAs0Tr8vYKBhBjuyizIN
FSI6v3ibC/5NO2/Rcqpbnd//6/V8F0xfvnP5CHXPyOlahVYeq7qcwTR2B+/9t5Xm
lAeimgrYXAFdzswk2UTYrJswfdJTujGdEmVGE7ZQrveG8DR0OCy+1i43Qm+w5YIG
TLy6rSYZlH1uNCkLfpPk2dqYgLfwtbmvPxtaZS7t1yyPHsHl3PgR5FzlCfAF89Oq
n1I4B/NNqblV0a3+WPSp2jl2UBeZzuX6w5IbMHxkJ09PPQnb/xJA6vDfOUprntG2
nq2K9Sb9CE4HLqw4dGifOdSocP+GBryOAQ1ULEZw5kFghIgGVxHPAPMc7/ybjEjI
xG0f7R32+BwjhsPly3MDy1urqKPvlIu/uv2AxOKc4UPgPOkr/na5e/4bTKkrqy/F
sUCTNjD57Dw6Z590HhmViQ81zQoxcRKpkui7V9HJ31KmKGJwUOqhXKmmAkRpvvW/
1DE4ASwT36au4I3tJhVUYpkvKjdl+zORJED9QK8FdursVW24P1tvY/t205Z4w3Yc
ncj2iiYhvyHD2PVOfA+qSw2ii/qhAVXPNSu+neTOfZ7yAPc9ANqQcIOYDlIdodzb
EzJQzSnWT+ETVxywz2WBRulC9N+bydywBdZcvmOn2VLO8KN2EaZeeGeJEByBc3CR
PGFtKsuCpPqWNsqepIqaGM5zZTUrUBJnNNZYQ8fOh1uGGBpge0FBKmoNueKh0r9a
5om1mOs0afSutUdvGBgLSdln9kO9+Npf6ZrQfgi0/zZ6CO5K2K4E9cIy17BByhuX
+I56RmT4yYLzUH60gKKdRJJ2NPP7tMVr9DPUOtm2RWfbq7UZ/lv2fsLyMsAVsDyh
jW425akmifIGEMiJ2biKhoeOebwgpzROpZ5WZ6SOqDtG456i3BVEIKevNRQafJyE
gfsb7GJweU4vibNyutWf4MYAGpJteqqOAUMcwzCfze4UqH2uWfi6xka3CmhdsYLb
WupPwn/67oS601pqHxUkOMmjj62mkYcic635huoSTQ7akvV4WED0vpaFYYu25pXp
L5slR+cBvQTDhfbvN7Pmg+4Wyn5v6FdpdkzwstnFdi25vdAhCCl95+bmmdx/FACv
fKcvaImC12oA8drkZfpF9RzreGNquq/PcculedpO7kaW1jRn1e10qoYpAALu+T4Y
w6fHVKpQIbtIYB+HMoktNY/1IG39IqjDUzr8Q9BvoeYSJO+LJL9886iwohcroqRs
fLqrwVpOySeFoGruTX5PyGvvTqx9teRzlCEgRSkf/aOvKLectWUw3ZHylQ+QVRqf
iGmoEEhzXv6UVVUlMr1L6h+iTuR8dOlaeUR0IM1k1lXnPiS+8j+3IT8H7QRHud1p
z+gLqgS+pL9QqgUW/RJTgyY4YK++of3SCUEUOqG2JdWvxNTbSlNB2j0RQBxvGpdO
E8ZQcncafeKfFb8IQXO3LjjLUr2jHl31/jHLI/9diDc8lTgz+aNP0x1td2h/7fQ/
Ka8igxiNU148xWQJhkvGZJdDnyBUr/+DiQGQCFmev3aC88YtFwlD4Yk6oLjz9D0R
ZB+yma/mlSyrdqnp0LvAKtONIZRZ7AUGjkSKsOoYolPCOTsiHvJAD1OgW1dtwPEx
fdHszkgmRxEfF45RHWI6ynUbsyz8wI/Pn9yCrFyUPqWR25LODXedpABRa3kUuCPW
kRjtuxuo+ei9ZpIln5kVQlyLxa5FtSvKxCDG410C/o4S/6/mV9lNqMELDA69/y90
Zf2pVhZW1X998lMAHblnWKK5uV6f11gJ9o5S6OUwyKlWovL+OvUS1KR/i/CFz9VT
adEa7NLQ6KeGs/nurC+xgW9Ip2sM9/968hY6NPTs9M21aJ7ITnO3j87BAsfJVfln
XI6EqO1CwuuM6MUwJFbPjdvGc6c0XDlqXc5j/95w25ZORBoEvmZxOTp2jnVRX+NJ
oEQJP4Cr7Ts/6NBmuPnVinfb74F7BgpLLDC5v1L4uFQ7ZSLXJMo31bFOrqPmHsh1
nR/C8kb0k5+/+KYwoRyM/tRd/NEXAHT/6AXzWejVZZahAeNqzkyjRv4OucX+wNeH
jBvVhEFKtgb57rDschQcqNTCzRZvrKFZ4YtAp3mnQKUqfQMtZwhUaJDwEeiO8tJ3
0yEhJ8j4n91ifNit7yxGNO1sJzmiSzKBd1vXXUbNOMEshbMVseq0eIaWsg1YRYse
7QdnzGAgpmI+pfmxTW9cK5BHKOZqBy8FI7nOd5/PIOTNyR/xgIlCVpPY6wSwQz8Z
jpN809vPX672JEBjTCJYGGINTVawitaNbWhtyR9ob/nNHM3lw6OLlVF7DA+tVaT3
kS2U8YXuqBwKfwwIdddJif3Zu0OfTGbx3IvoziCF1gH3yBCvTfbn6tZZKMW9iiUo
1lidqNJ2G+LSKIEwPY6Yn0cYBt4EZ1MU5kQp9EYLfdNRuSD+yyWVTyOPOUfn75s3
PmM3WvQw+CtcV/bro2D9EFw5yw8wZVFHlby5cvAbScsK6GB1Zr3REGN4dqh6gC5I
O6GbdDdq2fXpKEPFZS7S39N1uQ7Bivnr/S4fFXb3cEbIS7osfUxY8jyqyanqhnSJ
kCb2hTbmyIchgDZVeKIdCJA3gHGmtBDVTPcGVqrm9HYenUVCT479Sky+EWtI93O/
PDb3Wx6EqvJfoAmrMhNOsDkoxZyKEeYp29YwMlqWewQrhnj3hVg71OPh1Sc0rCFD
TLBz04i08rK2YVqo8XTWRaJehPIrMuzDkYaxp6Clt80jPnD8jizAqLU5WiDF19WT
+6/FaQtrFHGha5weWXYmBrl1ILvCfoo5g9rN9r+ANeo754etkPaHb1eiCQ/MeA02
pn0CFpquEeK2pXVRRrT312broZ95Ix0ORENIpilk3jy1RJKPPFRfzWwrtYR29SCF
m49dMrowlZ/UEcsDBt+SfBPf+vzEilUR7FVAhJ0Yeoz9FsaQ8jSz3EbDAywJ48db
u89mjp7tYp3Mj8ftPeFJqU6OZWKC7WPxiBHIZm++yydPfeKw22SqyN3T57Nm/A+o
bYseAf1UegsajMMVDuWb7ZQoV9q1nXTh7ESxdt1skD0BIhsKumQS+gskU0e2sxK3
mCHWH0WfySfgZ0K+nw/3IIBEo/OIAFjA/8848LNvrLR+xWXn49VIB7gcX/MVIXIc
MWe3gp7JGf34Dt2Itv7e6+hDL6Yvb5ueVQDJHP+ZSD6O0xgxFAbw7lRcDaCEOdCm
eTsior0lz1aCoeDJkXCrWOOhrsDcjKcSCehmUYbDCnGxE8BFz9AA4vaqRzcOMs2d
44WQdqzR4aGzveEUXUATS6pKIkZddaklVaOAyEf8vI4nz4NuXN6vclgOFQPTm6ie
j2mWzn0vjbEW2ViXDK+WgLdROEIh+EPTdf0nEAp6uyhm1Fg12Ni4zqp5PZrW5tPK
3wep4rl3M3a/OSyj/l1yG9XbMROkpjYcKArL9jOoP/5tupqWSkWv6DgMeoAPb2kM
y6Pjwi0U14nGmcByQIFrjg3VNOcNpVcl4uCEWT03VfjU9yMim5ZADDWlDunaxFAm
sz75YxOfWgX/LSeF1DLj9qcuOfiTYDHMWY8Nst0Zoo9oX44SjtBVAcN/5XTSf+ac
WFzQkgOl20g7nRyp0ppEu9iExAuXtKhN+Y966HoiGfjGHptbrz7J6Fv0X8L8/Pwm
P+tULz5BOqCgYpxPHCW4QjUCVicpeILdh2OeAxJQur5HdMZqm2utszOMwScqBiak
wxotzaLY6BpRig8DcjgpPpVizCvpFnBhvCBzsEuDnQRP27vzXWVWErJFnU0kYKWg
4tisrHkOWsknf0gH4+HxfMkv6cH6XruCwG/CSIWySXxSfng5r1DFByesvWv8zvkn
UtgWhNjRevWnquWF5PSiPRn8SAPgiBbDgZRiZh26Qbg4R4d9dSsQqaavw+8onCEf
dLLsK61595zW+4pZMTI9YcJWjFrwj0fBp/9FAUesGUcJoxmcqEkdrnI1QxNOkjVq
IRQjaH47jUZm4xmN4q61u9Qsb2/7cGPmHtnHlLYbvrRIXrEQWFKtR2IBD37LRpZg
5Dt+DecgaPire3EMpMkdpQHr/bjnQdBGimuV2eUica7IyoiqBIc+/3N2qUdexMz9
7XWDORrOFfIeP1DwJyiEqHZAIBIucAxATmoydy8GWcw8KEyuGGUQIkZzBNR9K4P6
5EK5xm84duUEou3u7eDmoiV536F3op64Bx/yfn71wmAyFaCiWLxoJreEivufRjt8
BvjDGoeIFlNoUgbYuarkxneYpusrYTBj7xQnpmBJdGAEdop54rQqzrFIx0w8WxBP
ig7KNzns5ctx0h7Y9EisN6eHDb3w8mP7VyvddjNXrV/0nMgpJ/LtjSL5s3UTtHQV
J2r5Ucz3UPrHR3Z/faa8nUC64pUVcTA5a/fAcEiQBun6N0gKhf4U7ynilL+iEdAQ
16Vlid4GwCOCcbXp72G8nd02w6+Q71KdRuSDd4NMAc6U5V3cCf3BNMOgWDm0ayx9
vyJ/x8+1iRcGKgqkN3R4KY0r0lyLn3F8NPCocHZQFE28dbRPmxHikUc94sTRwnqG
BkzImX0Ckm97I7Qx4oW6Zpn+Ue+y/nbetoQO7/aVqppwtBylHxaVYEgJna04SOFu
ehvoxti4r5Dua5bSjRP3sbVKnn3uvpXWIyOtpiQCFsCalnlwzKs4Fo/tHDchEVvY
fZTatb3R5LQjeF6KcmEkKs4soA+vI/wb21qEPWHcswSoebXqE6Z4l20Nz9aQN1A3
XFIotFvo0DGiK1yY+3bQ/Ws+I67izZuyye43u1UbEXzzdxhgkAFvtNdzY4x9Mios
WLsxWFiQZR8wDdMbnUPtbBm45ffnE/fX9opm4awNCCYIQKWeRH+KAWXhlDJIq7IA
uVJOUJviUsQlGKcu1oN77ou71PwOc6jUlseun8ML80Usx/XLdPrDLbf2H48LbDp3
c1lF7yAHOpttQ7R24NRe3Al5ZngVcWNZigL8qCsyhrTRUZVcpriW3Bqx4Zt6KQFU
/dK4V+j9MlK/ehOGNRH7b+iPKtADhZFRXSwX3kGemOn4bsymoRMyj+O1cv8MTR1z
teZDe5k8tQBMZjhwchO7+J2sMh9Hxi0INf65+q5AtNM4HFc/S4ngDFFimJhvcsDc
mXuK4vEu8wHgVdBSoSAtuVK3AxGapjD0fEaNmmgaKhZr+v/M5FBvzF/mwIPQPmMI
Z97rCzeglz5AxzkBQUtTzwCRJL2LjIiqAXn8aW2z0YyCI3RPNVz8/wY6OrziJDGP
vcyrodvhNZiT9VZtW6rn5IePTvSFMtaz9hicpl+mtwcIadiOBCWSty+RwQf3GEBZ
DW6VgI87rA6j1PganV8yUzhtfeVFN2LjRsVYsmmvxHQHBTb+7Z/l1/pX3vUpq8VT
gO9Kj/i4+qYyIvAKk9Ua4W76XE5KxC1Dfpl4ArpdB5dXX+/OROMBSZebAk+zVUtk
OtNNUdTZlCuJ6rqJ0+FuWUW/3QwBp1kpYf9veWY/3AkVInWcoUav036WSYojeSYS
wdPkvdKIfgB8Eou4nr06TmzC7ndUKzSAV0TPpiS17bW70U/eAfizsmFTDAQDjHe+
7vtqP26D2KeSNpMiMK5zmgwO0sx4rJsWSb213AOhqSqaRQ+w3SABiJoA5fNUJmMe
aK2t+GWEtD08vINeNGn01IMpqf8bdtwVZ7ZBAtoDL6DcP5ZYxccnCFDucFxgudnW
o0g9FvOmyZatij5m9CU23JM1AjbW8lGYBGnQgn0aC0dxqiMOJDLRHnNp4AbhtTV2
ICMTx73xUzRZilhOjisBGVzA/zoG0v3HKbtgJBHvAol1H/65LJoGxXi16l0s209R
aCd0qHgZRuztpqCc2rHGpYFCEaXxVkYDleqLqpFxYPO+C6DgVMt+BtNk8nz5qOOg
L//8xWtE7GJFfyGxZQYBRvW1vXaSf5Jy1RvhNVv/T6m0gyBW7q48vt3kr/y1AcLu
mGClrFBRGbi/UMl/R0WVQw2xmjvsTtuwY7ggTffGT+kvcaOUADP0WJbAjZ1VSLDV
2Z050Vk04H5dF0lkTH7GjwQrwO+wdbFE/NdvC3/wlSW8YV/CcX5MRkckfaSpFByg
LZ2tdhbzxMXylm5cWoTiIekyNiap/H4mp5uJWerScrctj7YRQpmT62MN68G/JJhL
hA6QeLnYhcjDX/+8bSV9zPFayRzkGPqKAPvH+oGsKyWDvKas2b5JfDfWOyDCK5+T
ZQ9pfk3D0WUhdYCP0Mu8R6VlEa82xi7ELxezxYXLwb/HxybeUhZTw3bVU47EPVTA
gug79Xr0XRlOVd+o1UnYq7pL2A8G5OKxEQXW8eQG+7z6Vy/34teCXFwhuOOe2gH7
quONBsy29RBbz20PFtEyfuq5YiBcpHH3Hqhd+DcO78oln0/JrKtTP8LOvXdPQK8g
2JI0Fpfbf/1QNfD4gWZgYfIolXB95FpvbwW55+QpZt8j8+CjQ65IVhqSfo45z+5s
J2DUG+9iejWAA8jEyrCzJaRjm91Nlm0XLO08CNTGoxs/uMi2dAKEO2O20Fe5JnGV
NdyS53oSapbdXrhy/wWuEXtSUIKsFtDt4qg5DEN+xfFThRBxq4ObnHHWNTbB6479
ym+UmYwi2zJMdzV65T5AC5lN7Ky399kFc6n5RjQ1SkzvBUYgLWCOqxENgC5UIxrF
xo2RWYkcJtoe6Zqo32nKbdcSu5xERCDzYAI//iqLTPtjmy722U1HFAKmXZqtM5Qv
wSx5pyJcXTWFvcuIknDVl1riRN37CteDth71P/jv9tn6zXTo4GqDteqBv02SdYws
D3hCMEIB4j1Ji4xlLBZrorx2GN3vordlElDyA2RIT3kY64FcwipBgz/gPnamQSei
qk6LG+Xwefetc5E7enlfTCjE7vLqLnxJeZxZ1y61H6KXJlqJCCM+wYOa1ts7i2Wa
k84U314EFJYZ6X/cPQF86M/dn7c9Hq9A/5QwzkuHHKkPzA7eXn1f2DEVqnaw4/lf
hz4z8BEw2X4WrkdmuWsOHmWJDq2QICtM35KbyXa692lc6IGybSrhveVHbZA2pd8M
aTo+mabxeTQTZ34KcNh12fgW9z1SFM6P14vyaviWrndP32PpkFUaGM3f1h4hL4hC
osEgEMxPdtSPHJPVZvPzir3V7KCgFPYWZhyOTOcJGgDvlfUzohT8cAn6TYjoZofT
Opv9gWpEQaRrQobD01T3nbR9/Kgnc9SAS3D/TAK7YigbbgJA/FOiOsSw9sU7Sz2i
hw3VPFZVEECTBekYEA2UIsN944hcrVbbC7AJzZ5iCNLJ2mlI7kOVgbLHua7Xj15p
notIS4Hr7mYWT8xDcZSR8T5t5CpYMRjyKQEEO641VsO+eiDXp42maEgCETxPmAH/
aM8VtRd4lmKXU80K4b+I61SQh4WqmePjL/egZ+rBH8JUkvxCR8UjgdfeWZcuxYUH
R2oQ6zaIju17fi279Cy6/NxL/44GU7WmpS3ICod0XR+8ixkmL+UryOW+u5Db2i6j
9PS6KpZpYNLhFSWBTuxN3oKv8k4Wss0Ev89s8Lp9WzHagIJU6un0h9qoHlyQBk5y
Of1glhGl+pUf7YsNpDz/umPx7eKJ1g4NaLFBGz7XypK29N8y1j8xo+LFUxLNHf5Z
3AVBwulYTDZeb1OgISZR0+spfoesUX2G/0Mu0W7FNfJzk2FYsQ/Hr0nuwErAXptM
XWPV/XIsj/ywNlJ1nTmFwIX/IN9e2pS/OE2vfnvcISk+vh94KCgDuXX3jT6l3/3w
/tCUda9FdVF5OeXUPXvpeNetE8d+ATdlP01Fo59mTVoNDdoRyaJV5umCYPtAO9Y5
+teeogX4LoiC1VaGUN1ZrVguhG9tywlnOvDTmRfnezYBuzzIBrcY8B8PLaODYq6b
K2mAYm3EwycD7va0FxvnZaD1wYVVEYb5QauTB5Xs9eZ9sRJ21izg27FU8K6cab2E
tbJSPLDXgp5onHhsE4SdSbmtX89nkWur/kJigMS5CdkB01/I/75HeontL0PFRZed
5MO8gvTgZXqETtFsbozDa/n0650eOPzbgVjZbk8TUfYZqewMDT4+xzUMoJaqCjvd
+YMbxZjgR8jc/oYYOxv+8lVvgkAfCXnAnfAoNhVxvOKX8ThEG6h6QC2ELlJE8gUd
kAHGZBaAw5SFuq4Da8LDUrNKVU7WqGaVGHWRIqY2rT/eM9H/1RETqj9rkawFXRtc
fa6jash2nUNZ78h9+DrmwPLZiLxscTw57WFBQfw4RMnQMiPMB2G+TddgWZQnX3A0
VRUhWojeIg2LtzRnaeuoAGNp1qfwCIMSb6buWX59Wn3+R5R4HCJPUuV0pWkqC8SP
7wOIuyS7HPzmrsfzhhVPyEouLkw5kY/h02HKGZNCSwZTPIDwXer1mjcAtW51HKXn
OuavZS7ppUG4fwyUKP7+a1eikHPov811laefw9u7QtnXR3PRj5+Z6GVhYSpWLLce
YqMgChqTPsqx5hPoTfXKKmADyUOR+lCFLXOSg1PhXcnJ+jmxLApbBohns5KBoRHI
Gq7cKe0Gz0+WHkcowhiu3LzGhPim0X5ehw42YzSdMUsTJMFwjknRuMwXjjGaWEOF
HLf9QV70rhGuRBKPbt/3UYPSvIp9ptpcvxO1Fhd8Ac1JRi8Z5JLd2nsQXkGNw4m+
bMbvqwYcDlRSEYux6dgC6DADEqvHdJ1SpUjpziCkd2iqVAwXocy3IWs4i5/Gyv7p
aAat5cth8nLpybRYdhwN54saBEOTuT+ELYo9+nvQ4MeP5jzRQbVjVCnHqajju50c
bFvv5xheesqtZpPyxUbPnSkRSBDkerJV5L5iUU/woIHXniayUjpieSAVHIUNhgr6
zevjoiPbt1dmdRQVNv8sCLZ78GCGjiXdFdQy00Yf5/kGDkA/dMMomdHMV9vL6zJD
0ODlj0paLuAiSa/xStMt/AA0YeiV/dUH2RqwMFaYs79SLrEo4SPCKTvTlllE7Y2X
G66/KBGVc2LPI3g6pcHBfqDBHhQIMauX925ClDoEmnjoy/CE1wzvILSTFb3FL4dH
SVtCJX01qPCU80WetBYp7PUwbSdR3uvlwS068bZUSAOQif9QKlxVDZEADw8381q8
bdkUs1qlJA/5iz0AKKZx1h5pNI/0ulhtNEiovj4uH+whT60I2JCXfVwWtbeWYiJt
CjnAbv9itze3sy8BmpgCeoSzGzLUS6NZKByLch4n/ZIisJ7F7HijCtzhPhbHSoFs
g3WlzQ3qi+zSjCb4CzAV7oTWkFHFShj1OFi4TEM7OcgBjZMgR3xvw5i8bZ4UKn5T
+CSgBSIEgiEuN29LARxBUbUGLl2GMAwyZAgcM1VZ1mabsi1OcU6CkHByFZoCLTs/
GtX3oJoT2QpAycssfMtxNn4dagX7r8t6D3lYujO14trjTnKrp2KnGMf0q/mzDhWt
Bcuim584vwkwpFZGqmEqoFB6AinhjIuiXN9yd2ACsrY/JUEN4FaUsZnIQe9fdaga
i3W25PE2NwM2lhOCx+xZGzJim3rhX4MD1Vwe9AQGBzO0DCV8RcAVxLJ5u+GFavJs
cSLE5N40bh8MJEYlu7TpkDsxoeq5nhsl0NaKR3evpiKUW2Ha/YHY05edgS497G5A
o0HM3Em2G38dZyo9M4jCxxNYKetVg3blsCCzG9F2qyMvLqrjOEE7gYag67yrsIdf
3Ov2WFZDRNUlYfCosRMrO24pCP+Ji5kAVFXEJ/DB2GwffOB9xUEqcC+0EG1fPrVu
4KD2M2VA2gBY1xGJk8U0iVNIitlOklBtmTnL2pEf8CPCQuPLnLZe2qY59LKak+i5
IoCWBSYlUQOO1ZQ0O/3DJoKqYj9AOATqkrSUtm6qL3hralkba3G2SKHLvgGGxowD
hDEOGbLAaRly5ONuWM+BrEi90lFybHfBW3OS/xGnqsUFtyIn1ISYOw2WNUzv9Db3
WlCg9GozuZoMivbquKnLvWW9PDIX3tX6t6zctQ8m93oBv0ctJXDufTu0dIhrAimZ
jN7QobJoyCjB4MuvwkjPY5olNhaF6HUAWLY1vTqvRkO3HGVpWMjfTBpfm+rXH+EE
G/LNUjyjX/u/xSPZz3+UcrTjSQ6fNl8PqC5FyiGObKzBZUAUbKaSSbfqApcMBw5A
cOurb/mlB9YBziyqP3BmOrpCzJ6zdgzwlsTcByn9nVnI3sdTBUVeqBMyOoeLaioz
zAPBgTIF6yyPu1dD/3dl4OhlvxVe7r6Ynvf10fueGVEfi/D6AYDxKlnPs8mzBwuR
Aqbl0gYrk5/pDAd37P6zdFuMvG5U/n5bRrKo7VYXMhrcSPEIMypW6mhbI+WKLAFQ
+3mZH0Obf560ZVNF3Zke3VQ076qoZq0QMpSC5L16OwLwAqhml2cOFI7qC6/6lGYO
fl3rj6/iKNED8boyhBoD2UxDF/OIaAt2aR3pxu04WbYq4ToNVm7ZwQJ0AIrBNf25
xafNcl9nRnXz9tVVUOlgsxh2KCOnZGppiBQllQk7fXhd2s01j6QgwE7fVGbiXlEf
bkMQwtoQqGxMQ7yvoyDgItxyxiRAPEGwHRb2XbjX2duzlfo8E8Rn6KyS46Rpv4hK
njqm/t19jF7L1tth9wNmjQBLLR+jgluF0W9BiMUHhNsNlbytFpD9WnIdbCHLJdDB
tOjE2YMsEaGS/jbHYaRGNm8RqEWChtFZ4DFvRtUSjT9GZuV8TzwJ5f64R1+BEpwu
aYHJk1cFGYJkiFbIcSe989lfnn25aDC8i8kZvA8OpAVJ9CS8WpUJ7NkgJgJBI33W
964jDsUttYxCrxq2B4Lpl3FBoTTyNOptfsJ9+q3vDx6amOSQ+LH70nlgpiHNdaMA
ENdgt6XotUtgISA2DuYZS/IUkDjnHW/1VBklTf/lEvRbenBDutVkH5X1/a0hT9NT
leFEAEJ/JZHHR+cxo+lKEMSZg31aNe9qCoR0/MqRHeuDkS8RoaPDy/WiN0FA0zuq
2LCBz3HsAgsBmJRWa9d74Bc36ram2Sva9mtc8m2FfUAW/35h7bWaJh+Z3q64YsIE
AaWvvrSQ4aCTkVA/C8EEfHajbIVBp4oUWWstGvWQnbqugklf3ifo0+uDf/ypx2Y6
9G34Q0T6tHO8hR/tFPKhiBWxffA8C3lj7SyANcdZwjhKq4ZNmOAulWMCEPbYqyVS
NZ8BN21T8i+0SUobbxvOLHQKGYzTMGg2xXGsQN/nylqAueb2xLsvw55jllFLUiJV
Ffsf8NuVQQx9lv/C4ALu7IQqXO2cjOd0tM+61KEwxZxiPE/8+C0SpiXvvW12o3TA
apNad2T8n2Jvh0LB17Q8rjM6BJfAiqfrl0+WO9S5S/JKGiR1kDZRhu3zdTs7JveF
MneDXv8689RdIJwdCq8wmdlQohnG157mQuj79f454y9xVYhX5XFiAe4UhmsEw+6Q
s4Ffp+dGMFoSgD1MSFtWtoZXN+et7UxGDXuibu1VzGmFP4V3IRvv3yGFq/lu3lZQ
Rpd4bF1ZZt8bbtfUnY2l85tI76sXNjVmJY1vn1pnbImm5NJza75klyOb8V8HPEJK
5zJWJrZJK0XR2xSMyDiPET2YA+geFsux1cv0iDCbhkrxewwSPo9NDUC9euOD0OFu
PpP+su0A4aGbRHZSRmDV7gNLCFd4GUN9ChHnOPscPE9BCVOI2IEGoZdLchm1rVdq
xuu7D8EHZ+Q06Pdj1N2qxNL1Kpf4CBqw+wlAmFXewYvjEFBhUH7lJziQH5ad1cRF
5hbQIfUGVbgAHE3kFHknz1SXGpEbcmf1uO2l/08b1EpmWd/p3KgPz4EiRS/S1F3K
dhGxXc+sSZ/ibAZqR/6lzbrakpABt1TC9qlaMgo8a9ixhb/5lZyOBcRdaDyfCOpK
SBczOhMAtEOuRsRFUAFS84PYTBCclOPeAbnAw0xoWnlzkEZfyKOD3YUx0jJMYrFA
26mbiYaRlsmg7NTNA16xfal1vsVq1frg5znpqcjh3KBbOtZvb83D6bZwFkGT+Mtk
sB6thSM5aOwUBUbi9UTxlsini77xDoLK+ZdyfBOs8G2UuU8iTnbFFa/v9/h+ZC5f
nqx2k6m/ghQOY9G1sjEGuN4brnINr4V9LrD/nmqv9BMSL6yyqLJxDWX1WIsQIaQ5
OcYhc5+w5ufHVlunkivMHkoR2e6+0l2JGtLHjTEBe6+vIEfz9xGsVqeU2WzkivnE
BJVVGz3XDRQwwx0dOhcYwLF9j9lLqzyU22JIi1UcwCEVIuwaUAcPcLfeyc0isqeu
XTNXCsDB/wXcF/qRehlhDCzZxIrVpKBLhdGN+bscgv+utIGdM3yLYQD9x6xs/C+b
QTayEwBNFqF5bnYJt/IxVDrwyCNOTHCyiGVgj4LPtHv6mcnZQnQG634uZmugLEWH
uZGj0Id3Kli0uYKTf9F/OU+W+5ap244wGZWkyAcOevGAQEYJWPmXHaagu9TvYo5z
owoZPk5/lMHmgMvtKhuO025O9DH4pm32M4X2RwrW8tslfp7wp8oNWu1ysGt0tta1
y3tFNexddsWogkOxq+PszvLZQghxSad6oJ0I0gNnhLBC52NXkvYEbNVIAlu92wWk
jpMkrw7i2zyR+c0VOmJVkcIWFqbI/GUkgw8nGaceurAYhMMl/uoDYomgJbcD4l4O
lxy58V8a/qagyRwq5MAM6Lk1jWf/u2KdODEDg9M/ut01C//VZIPF8hWIa2E2Zm7m
dPo6DHYAtAn6MBH6fXAv44uZ1z1f0waVrSOExgOE+ccWuD0nDX/vzRxYhJWWcbK2
MrbW7EYi/LH9hQhpWb4mUsdkiL9KC0986254AMPlw7CtGiQcc/JbFYAkDtbDTc/k
/yA5io3ooZqcOzTIKvAWcNWxpED9QTKmFN7OrYJXGn3EGXHez1Lr5rFe3ALIjnT5
KzWCbs9bRGjjT3hNuvFBEpXBfOOwhvpcuUhq+1hTylJ6CIjN0/rDDRtd5PxiWgdr
wH2pwXn12LWT27F6qDgySRUJYJ1/lhrTCVmtGungb5zyAN0+36TG0aUElHNZg0Dw
7ddx6E4dj3fogfPiOFVLOXc/QiFJAfntIA0gwZzAvJfV5EkbGavjlQ85Do+L1NK6
JBfiftJ3kx4Lv0UPaCgLFVU3UJ8xiv8zDHSoROo+fw0/EENq7c8n15/rIrtCE2UX
2FkBvb5lFhfQMWxyvip1ZknX0/mjdSHwt4YFUMhgtjhkeTJ1oACc1EfgvyZ4yuF7
dED+Lxg3SepL3AgZXJM1at7baq/SWkbyyWX+5ViqpLWTAqpXJSAwbvMJUvFYml4i
jOYk81tRzWTWxclhc0w8zqBR+OBC+swovJtr79ngaaxTDfCcgz43cnFZXRtU/Rx5
Cva1/lKlLBdvhlwDNcJ2aYeO6lBYWTd7PwRkYhLck5TcaR2LBS/emK6nlctF83Ej
3OuEYO+BG3ZOT17jJ+2aD9yuB3UwqLOMWccLxWT9ZL4ItURBwhlTlYfFHRybJOlD
k+5/zzkAoPfP0RL7mYZTRvqxygRU8agGHMrvlIEC3n9Qn+COgqbAkJuysKR0u25s
ly+XXCXzWerlr+ZCXHuT60LGoZexx5HTUsvHS1ZQV3CJTUcAthGceQzBxevclL7M
jn7uTbAqbFQERQDC57bJaLyYtKgw8pzqtqYB8Tb8urBPIweilMh5pg8bb/fxU27N
+D+FCqMSSt7uq45B+v7YTeVtlTpU4IZ9Ms+4JP3lPiVyPVSlkuCe1IwALenbUkbF
Ttfl7U67DpKq+pk6gestDSgS2iGeIcekd6pp9jOGLoL2bQbN4f3PfCpgeaEn85g9
CZKFucLCNZ1AMgDHmnr6oYHJ+2i6D3z5xNzkZygJGj+5zzabkmXaZrYpIsyHgT4+
+bKm/vTnm4kbuyccxT8SaAn1iZGMcU14nt4y5D6F3yvWWYcdNA/EyS8vkosv/1Pm
KX5kbJiEhJLfZZdmEM1gtGFoKNzM2WMLUqDcz2yjxJiPw32djqV9a4ijRGZDMXno
BVpFWSQfJG/gu6fvm9qdtiGr3nZgm80dGaatP1CTjDEXTDIYhDBo/KDcuyUohaEa
vlKHgPnSyDfYRRTvsTG96u8WDxWO/zUylEcmBdNmQTTWNCQ0aNcHAlu/XddxWR5l
OfRQl3Yh5EAIwlxm39ri0So+nB+qPKbgDBXi7yQH1yZp+j9NZ8d9cQijxaXvEjv7
VKdclNCiVB+AQi+cqDJ/U5FNL8sPWFVuxK6G1PHcXpnipHQCTUQubSptV9yzwMAV
COr2XTFGZtANCvb5Wa3S6M7qV2itcNMCgr20P7HxbBM8jd6AZz0M4HcQZWeXxtjJ
13rUOceEXLMDpEDQtdcH5szun4JYg89o6iaZi6GZwxZuHmxK8WKTJpoGNs6/xA1z
ady1CtG48hbdbw8n1iPxA8sKPch9esmwWz0WwrhCWIoqQqS69Jf8bhAtmrboj89f
FHxRYWZRFh6s8aJkK3G7qO5lYF4pquwqiPJV3/5yUmXMRkqN5rMc0kul2jEeBZ1f
KwLDrDWIFHZFUHPwDWS2DNyHnlQyWVB79TM5iggeB/vvN9s6Kroo6eLee6nO8EoD
rPIvZzRe1pkh2f7Etb3nhaoG9qw5F7l7WQ/wrwoCCsW8UXW8/IKnrdNs1FlTxNsa
Anx++DIAPMVFKsjuLuO5sOrIJwCpSBaD3KucIPA98QU+CQOR2NJ4t17Vut1xgqSW
1CkNH1B8UNzawq+OE4u1VghLi3T8tvze9ai1espyx29lI6Z0unv4+hM+dCwn4oSZ
/7WbAn/MRH8kZX2r/nfm/E3Do7NP6ZbA+xC9ZGdJTkmEf3g1+voPtYxL1joRGIP7
ifw4sZ+CMAwFFr+6lG5w789aCEwLczSfy+99at+SrVB/7uB9L+XctznP5X4mGeTi
ZBBK5D0q+Ja+/dHRxs5y6UbtXcPy5oJYIAk6y741Tzo6PbeSanWzvrFyYTzbamfn
7E1jFHWfPe5UC3DdDui36/Gxd5TpbzA61apyNj1XmS+ReNHx1i3YXyxHIsCvZaDU
OqIiOhGDsJ/eWdJFcPH82KJl5PwPFti+/WB25/5Xky7crVaDkwP5DrHqUsVgJjuy
b5DyZPzy3jZd/Xj791E/9Lc3B+4/ZYsj+wYuGH+1+i27wy9z01mhmOE/fNzdYc1f
5OLGTnL6uY1T/CRFNS9vmAGqe4HHYNuG1jA8aAlcc+FnFeuQconF6QzcXU4VUOh7
tnDP4qEsNrFVhehQGSs4/Hty3QzdlCk8CNJjP3CbtS83qYJvsqsmU8INJgGXXxTA
slTfySl9SjArE4Aj4GF2Ex4WSuPDxGOn19rAyYGlov93Spr9qP+504U8DRGZBB8K
twQmFojMg5uwcDjVNYniJoATtY6QaDcZ9bB8jUpQImNBmSkRlCqGcYwdptK7dIhu
2hUNXh3bnsL1IXojNjPtS9yeZndh8SkFdmZ0F5BueVtBnjm+wEA7oxMPPOH503Vq
6DoJerDMAnLtBXd4nunskSAKMj9VuXBAvm6qBOVL/1dFpwYJjdpH5nlH3eODMVj9
BzZA1ANACdcsoWTljo+0GQJPOY+Pt6zb/Jz0Dsu/jT8IZWO+pTuFXBelQBl1N0Y5
/5llIkNwSgetVNEsnfSnVTQQ398yunN2MSkBW7Erk6O8PT9f7vcMHtdMjDfxFKb2
6QOaiW4sbmnsfEqN17YaxVQ+VoNAncGLHGdEDYUS7GkaDZ4WTf5tulF3fkugXel+
zM9VQBwgf4pVmgAs4SUxvf8VTrMZcMBrVCuw+ErcKdTP/o4qj7R4qy6tDmeRhoRV
lpdpU9tW54cShzlYUT9ppEw4hsub22LCRtHUI5k1ywmSFS7lWnuKtZErIs2COOQ+
9ELuHKdqtwEnWpruFKFxf3AiNQttyGX3Aw4B27afRaCXTtt+fVBXa9cBhTDdMkXc
LeDF5F3RLnZXP56PYY28uTlMT90mGP6MLm+BnYrxWD71UVXf1lFouTTMl+yuZ1Nn
rxybqgOBW64pRfiLgbvWF/CdoABlUkWnhvCu3Xns73ZWEXcqEpk8UC5LrTUXxTNS
szfjhUZltBP2XneeCrql/e53bGp8UKcJPU7L/6XMoR81zF0DR51WN0+jXBcF8LKZ
hBcEVvdkDcW6XqoH/lamHPD9+BP96NojGauDU86JGfAc2JMt5c7Pgy8IrjaFVtNi
jSkzgBancGHohnuoDi09+1TAltsgVIB8Q2gP6/sZgR12dvirBt7BLW+tF+rnvAyZ
XlO1bZG9ZMHJGxFBOR+UyuGMFmqFdTjHGnXThDn2hqUuJhY08TXht/0JtdSGoyK1
k5H78eSzM7mLMWEhU9c3JarXtzulPF7qYGLCMP3kCNU0ArrcTGl4hwofyxPDQNhW
6TSS4S3rwAYEbqGW7ObmEJggeRnYgsoOLtKe6e6BAoUL/XLgTr2IzGj9hKSEEYOm
EVekNhP/VUDTuGf88sX6Jr5L8fQUpGC9Mospmdm6cNesEwufYAk2EU/cT8fbG3B8
ZkE1PEXDOg43BkgPfwFfzIQvBkxZ4/lrplETYh5G7LH2ST2THh35fVCyai36SD1I
vcPO2FVp7DXEvOGi1mrJnt6dgIG3w5OA/+yOs1a3TqfKUcGWPi7DpGW/KNeXHteJ
MoB/B/YduYuNznAxh7F/XoN3XfWcTwUPH54S6wW4sp4q5iUHEPsNFGxzQ62vcylZ
S1BFQI1IfqxzfpXtqcV33kxtP7dmaXLdN5QOrLOUYMIbS5C1BvmWYtQ+dTRLcmF7
fJFyMORDn5FDxhRpdqADzo17GzcNvqtQVGd1099687yqH/EZJqlaHrUaLwYLIL/U
4875nb11F0J2uGxACNJLAivKaaVPwKLu2JUQywxL2Vsx8EWY5e4NvBKk3BQpmX8p
Lskm+K6+pJA+yc03DQZwxrOmEfswkA1lP3m3giF15OffoR01/4q7pS4Naa6vFADs
duEtHkbT+VSIG8xHoTm1hbUxGp0DRD6pyWVuCzZs+iacjqGVPqfOr5K9t1TZy+BP
4QKV84XEtbR6x+ywd6H4XylOm9xLhFKHvJMtZMuU+bpCfKGgPUTLh8Jmw5WjJgkv
JNNrfGIMXHhpwwzyX6OsXTxF/8YmIqEQQIQF2QwYUhOZPS2WQEDHWmQBnu5XwyvP
c3g6FmDQqhTx14YGy4uk+knxQ/aBfKADDnKi1l4IpwNkOup97UYANwvcuLGeTkZP
Met0HFh0rAfEJxojyLbHYIBIDDYbS4jK97bk2D8fSzXVHWEQHES6riPQsGHf4RmJ
7dJGj2lbpFhPPiGo02rdYKUrnpueMzAwp6Yfd9ta45NQ52U68RtHhTvP5AH3zfnf
GviDrYn+Kuiwmn7jgwXpiioSQnZn/deEMM2dsUSwkMEALhtbWg37RjnBlxsVSZz4
4d0P25ujNXRWEVyuvOTyjRh6/MbaYasj6CTTUCgbu6ijZe2e11aeJwKHUGqpfx6d
4bsKPYK0qivfdghYXNIXHznQOFBRg59qImRkQiGE7f0TYCOImBhu4UQeiDw42ues
2C67zY2SUYexTcQyFajsonzpwKdR3pc8K7XgODgmON6G0NOk7rZvXF09FYjOjVyH
B/8pyF0rszo5VW2hi0SJxFBtxUZZcKDD2tgMM8fkuXpI4bk9gt5i1eM03BHdqnOF
NSaE+bsNJ/Mf6/SYLfeK585XvpaxllPSNPTVl6RCKeS9koONhvjX2TUvX7N3kzu0
67cVRGe+4CU/I3Iu33wI7x8w+P8iyQ3I4TUFTJKkLlyhkl6Kg2ZrnSny7/JDynLl
n3/IVeqZzPzY6V9ssOXsvooNLYNDLJgXfTkdwbgzYFQ9cBI+aPdu4O5yM87UwqRi
GnxEg/K3NgEHGBxbZTs61vPUMSUegPAJS+LJ0ag/JOeFwRWmDAYkuNmGsOw9w7rw
tYCDOJC4uvFyAA645YVgscUSjmVEvT+ozj04BD3aaSiygNC9dLVztozGorZJMafg
izjTnBsHS1sl4scz8QMme0CFZQfOdvpvuqlpF+UAjiNFNDK1kRe587y/4PUMiKkR
H0Zz+yRK/fAj2jX+46FxkgYzTTug2eHlmdgXLnM+ak6ThVj66WgKjNOLwuOFfBsc
2F+QCAFVM05IX031/tupBJOLYxyRLhM8T7Rj9IiRe/V0NihdoYepxm4jzaqz4iAH
tlxCjpWKihCGsw9yU18GNgdQgi8OwccsM/TnO+RjEMqoeDNszx1QwvdBAVngxr7d
CuVXHUTZWPVMjM3gPTgOf/Gw0AycePz67jUlRXDe5CtManvXvALycBr9+P32+qal
3+UGhg1NA0mnHB/CaYChTqcKOSgJoANp/gTlsTWA/f9uULTIvCGkNqppftDjRZ1f
qVeaEUnitr8JgKJhTzIQysoRYceo/1oV8PpaEUKGQPUJpeLX+zPtZ53lsrxoHgka
xIFHgSlyftX1hGwJIFQ/DF2OyKbuPY1i9m8xjMFFUoY5/p7vg7EzctV2vWOo2RD3
kaYIauixVS5jCk4jktFG45nMwnYh537rG98k1jrSOiQJDXZvXyXFI9c6qswy6B8M
heXpIYuW+/NqjJfIIoSA+wAIRl7Fa9Stu/TtODBnRQ7/83BB5wKmnTwt3z8EKuWI
Dve9Lpj6VzFOFWd4N8LpJP+L4i83nFbs+iSlfPgGnjb754MQmK2mLPuYyAaKT9jZ
j21OcFxLoQE5Ig92YsD5ZM6eqECloTg4NQ9mh+zeUCnK/pgQhoUM/0BASUKmGXcP
q37/zQm2B3o4vzRrrlZSLKsWZr1OATwfOteC/2Qtsy5Jy1WRpjYGFtZA/Zm0Lm0I
EAlRLhXMe+rsz6S19w2DbKGsFOpC4r7vnA+0VEw17QbYvJkexiA1QRGu1kApwtlQ
3fuh29JCYokSHEhXvUroSi/DfE6TMXt55/k1Y+8kK4D1mgtAZRYaRk113gfXi6NL
rApW7ox03Ph6OSdtqm0Aqcd8YgmG70mkBih7DJtMWSvLAF7JNW8QOMjUkOckScwM
sKT5Z+6sXbvS2auuKmTjJpTGSAFk4sYrbOrZOR12iV5MNqn6x0/JgUxFnpAbEHWZ
pVs1pcnUgGrYqe4WC6gTOeCB2mobmmcqnN00c8VeoPJhKolaGI5Gj103Xlc90OEg
okWRJQ0TGRRc1YZKvTDgobFMeTNT+kZ72B1ADJfFt5XVsewSvNZHhjXxAKlTE90b
qDFrg8ItPwOyDosf07lcKId0Ges8/Wrj7FiBjl4ucjixIRlyNGm6kTr5T5cB/EdE
W/3ml4kS6AQhO0iVIRPMbJkxm6/faMN9fgSz2gz+KpcKpuznE87qafaVzR201CUt
iq8TVrwqE8bqucoJDOHKFSfsc2x/Pio9JSu/RauFqiNSMcmqTR/BtwYriXvPcNAj
7Lg21iyLjHnXrKlbs3tKGu/T3ejBCA384oGculDrQoBk9gBc0H1rVcx/eDMVEbmj
n8iBzy/pQy+crOM8kVrhTCNqJMPmYpxCDNxCupTmO513KXZ7vtx8/4uyboEQyzUl
dXEceabcvJ4jPVW/qfcLZZye9vu6Bia/gplOtZCsEkd54eKYuQD56xCt1OmQj6EF
ESkqfV2fojIvA+4+gjWbQuFfZ76iMY8Ij9PRbQ8u0uLDUavIuYTfrP+wDwzE6O25
r0ZvvZteMVFRV1QVMaKFsM0LRE3C/0UWQq9cLyjAUdQeru1HjAleSivFYJKdlMz1
YUqK4tpnmlSHPXvNgJxuACTDzASm/zlo5anisC5akOpZmo3PXfv5d87SqxPbw97u
3FGx0gVcTEOT2pASaYYI87Q4GEFpLyFlrrHJ0y+hQohQTbI48iwPpWpcT9tFNSkz
XP49SCoS6u2dbOXFQHp0GS3pI3pASlslDHcLTCl60l5AM4DyRGzxTh2PdJa4K33c
dc5HVqZ6cHYJ3kNh2yOXDTJlFVBf/AF2WrFUjlKOdSDXWtvLquAPIk61LlTlXaGL
bBa3Z2+DbA6CnskJLcUqRfcnQInLp7WKozl2X1k2hOqFznnJ17c5UaAVktJBtbcH
hC+E+UBjMJ70yypXY6abOmXcNIe8/qzqPh+CwOnE7lRw/bdguQyMlGXrNtTdx1j5
FKUml0VjMswP0jG+DHNwW3Av/6yjPoV6p97ZpWd5kyOuYpVRqb28vwQldf8f7wzb
MoDxz1u1DpJWxsmEq9Bq5m8z8anpZewoyQYT6wHbFTM77+s2bBaIeZZ+mmz/umWG
TG/PDPgJjRvCfw+fZg9dw9KQKg9X77SMjVaW9XyMGVA/0uFuOYRZBOcfjQ70nx6g
6TdjUAJzhoGBl0lRs7+1incst7t5MQ1RyG1GGOb5v/ELO9QgU4Ny05Fi4q4MQM6r
9SWf4P+4mFTqfDC1wo1br/OQn2yAN1WV9/KHJmBVsn5ZtuZatw7rSn0/jdRqQtp2
hWlgHP2GXNQoAaaC8nUe+VHfqr0xO5A3p+tLHrGCL07xeVeScEybT/XhCNYHdysK
pyNOecMziV+u+bAXh2WOLxL1r2RpUnjBAaeVYl2oCTZGO+QzWk+NB756PAbN0fLt
nI681SQPKthrWlhUg6J3ek5iqAD/HFtOFALTrlc8v1Hk2fg5BNLd+JjNw3dg4YnY
nXedLKdkbin67eWkQDzNRsimMxqBhRjh2jRgXSVLGFbsn5JKxHahqqdnkhlZSdrG
vAxcNCI8SBhiZHdHXaTVJRP6jBykmfsM7sBqau7A8bDfyRh54YTMv7pHYf2ilyG/
MxXtzZnCXuToeMwV/jc151HuMIhVQXk2PslP4aXv9hxqCQ+3kGAp3zwWe/9/QCaC
wn762hPFhBflxXKokviK97AcEPIY3idXM3GMk1x626Xk+wp4tJ05XAZM4LhSE0iD
dJOzPL4T6UcqTqfTZe8JPXg7qjbeA9c2IOVXRkPFDsw8U25V28pxEu5nlNNyFdpd
sAVNwavEnbWrn0fDcknGAskgQLU7dps2MyzrL2VwHCTTDz77jkefze0OLCUwCdZo
/kvazGtu0RMb9bpRTFxtTiiDEzeRp3f93DdagCYp2q+fMk09RwZdWKZbMVe5OfyT
RadwN9eqpZCnaTEDdnx9Jfpi5kd9Dgqe/TdAChvJEsQTi6Vv+PYan9xLvnytDNYh
t7xN6gzjEIODhKAKcswPY5v6GOu5QLWRtlmlXrJgpIXa84meueRfN+hq0I8UXZCo
1T6GkNxB1m/+ASjPtiMsMeStv0owtBqpNeoJtAjlbA7cEztBW/yIeltAfOVz8K6p
+lVHDPt+lVOirl3FKhFOB2WJJ2c+uyaMUBjZ7YWHfxQmBMlz/hhAgD39NMSz6fGz
oaM+bML5MUiDuLkQjGaNgsGpXo+iY4mU/MI0sw5bpT+nH7TbbkR9ZVZql+10hSsP
rRPjUmsaqB+OWD7pc5CdAQESjItEjfpiPq+K9PIaah389A9O5DDcbESaodvpcavv
ID6aoJQaVALkSEmD4p/s+BraluO5qEvXgoomvfc4vb1NKMG/IIj8V5/6ZTa/H4W+
7x4SKUidPtGVX7/fYe263V/BxjSmf5FPD+M5ihA6TPeVyrllAyEWoL3Ff0G4pSAN
6jp8w0to9cYkP+46QCiqPug/HZIK9dMeTm3lLebtRcy2NVx65WmKsujAcdADTl71
SvZZSRh+rEByHYi1u4NYNla2tmr1EsfyCB/DZldJvIzwSUS/LJGQnP8rZ5E5WN+j
zkhC82LpO+QPUPp9ba0k1I3otckO5z7mA8jPU9ugYcqr1IY1gX2ZSXk0JlETnYEC
FaDxd/WccAAUsnu7heqrP97/mnOBJzk2IDSWEPN55yyFqcjRSMA96bg+zoY3PHPb
aDSB5q2qojnqATr0TItCmkSUKUUY7qjxnNRwRsuBdCFOvQC8vZocHLY8mX7/lMZZ
udDztQhSroSmbE44SoCbLrV1CnwpWxNYGks+3EwGH+2HAJzgdmp3oeRrTTFqX8+n
YZToNiKEFz6lMp0+6aapt03oy3X7z18wCA9hIKHGEUU+7GSatUib01F50ozEXuxD
ZVVP6BIplbVfd+dhFHyHJAA2MpyunieozaYHNLfBW45v5EZ8UZDliwYywXDFNjMe
5GNuxMaCBqG4U23M54Xs5jV+ARETAje9CZO1KIVf+gTh+Erq7pcEekr8FoSvW8EW
LrDKSREc2/m57+deCXXtw2NJMiNTDORH9tWFaAGCRRtWGUSCOWpiP0fvrS22LjC9
Y0VAVsMs3JhcZfyAlrnVrqO7i2bIfRnAZgl1gz4Z9UVrEiu3VmpHOD9A3uiU7t9u
sftO2Txix5cWVB9WT6RwSn3bJ8hKCYirJEev/Ysdfj0AZsoqV17K8qW9j4TzlzWv
lj0ZJY0osqWQwWq56+QTEXaO2aq0xZ/wHW+FSL5lADSjikQAjJ9eWdE4bQE1l7Qy
/mDUd9HKjf8PRysRaD6ICM5UQBUrt8b1dCxwbdcovEvHFtgQQbb1TTAhb5MKzzMG
u8RCLcyppwfnQcv5DbkxvGwlXaFku+WVp8eVMZmkvQPysPeERt4E4z4AsBimxAyh
udo4kyCGxXQ4OiVnvWdaOt1ZgByY6daoU+7xzHThWWBJRzcLf+OdQnoSZ5814CoL
gsJg5Y7KvEzCA6YXqLItpPeCYYLZSo8PG8UHDpoYz8Z30gmLEk1i10ZrUA9aDpOT
3oDwBi1RLqa8VrtIBB96A/ovPNHidjwZn780fiOfe9zNC8yRtOs2bBnMIGA77NoS
g7a7aX+L4b+moEXyxyWUGD3R2e2K57GFAcdxDmOnJiYOkLaPfVUsqeAkVouQ9eIq
XKmQqxnjXta7+3H4A7WcXJ/Gm1SqO8QsP6MGOPuHUFOB9+jevBKS6WYQ1NMNAShk
ObuHCNpnGJHgKIHv+QtI3pQQNQ1MZ1Vf9tGIjEaPUjz0mvVdxxcly8AoMbI6Mj26
cij8z445Y7IH5mDEPiGwmRxyeoENRJPpsYViZOHk01h/hLpZtLbpRIVwNOKSNaf7
qsmDkNHNeyLZZ1ZnBUNYuADuBX80O5cLjiPg1IJIGlFqQp2Folr5glb7XfwOoPSf
FavCKGrtiZzV24MTHecuH+SaL9HrZ7ic26gsVK8w2kCrz/34uoHfjB2PLcOWCzv9
jMw+93eFfEU/OV4xmAl6Ga+Ir9NxhbU8WRznbyQCRXEYyjLcMusMaEGrajqv73Fm
w0XMV/Q6RMV9U7nXCp/I0sGTGTfrKZv0V7fFkaoILkDoJKelUn5LfjyIUQpyZOgY
ms647+WYCH5gRznMI95hBZKuGoEn5R23ZyTLIV2fm9E26zqCWK//kmdRBOjMI3Md
l7X8NSDs5roYgPw+/Vd/pTY8ld/7BsdPcMMYEmuCRhF1VQKxITuNrhdclxQzg0oz
UKM9qtWLezf4NImEpApSulPDXSc5vByhadSnAePPxoJuFF9Drp5WfmhNo7Lmv3PD
H0WGuhOGUBbgiA2GwMZzSAmACxSt8b7YMvYT+Vhv0rr4BD3Ws+zD7+hD/ZQsPBGh
y5bAjd3N283s7JgdfnKe03+4G7h20KgUkVIwQ2PbdQvLuovUnl450yg2vud+g+T1
YTBr4A3bF97720iPwRoGPBKXkpI3724EwmNmm7i1kjzGxto0PnxqeNX6FT3Vm+Df
sEjSpQGqJ/OAtNKkn7ulsvTc8cMdaikR5OzqZs76hQnt/rvzE94eRkFwilZJxa7i
Ni6m8ntrpRYa9cXhjYG+N+Vb8E2Ix7npPYaHdykMLrdgnFixbRc+36T6I6lXVWuL
Kbvy8FQYTuDn6Y+v4I8448bxz+liIl1V1z44kkxcE6BGLlnmYROyEyQrtAkpu0PY
yrKEUgtgKcavIwlwFmbZRLb9FUrxk0ag5QSxBAqZkIwq8kJjXDADZvemz3m8lX0s
HWifz1K/4vsbFgi1IT+qT1kmMQaXLbCoYHBiMMTD770VoDOz/JeMpbTyILgykEyB
yZ35ty1RUaMfdRcb9//tSUa7b/c92pz5AdayNhEsEbtRzsfXRy3M90O5zRO+rui9
iTAxMHbIaP+kPN8jQLjPiqZ8oaIUFacYd663pU+YexCzDf1KKrK3exd02BtXBIIU
WuNde4jey/n91SfC+mofFE/3WihiTq/NEBZenH1Q97BeK2yBDkdd00dnp5ZD4leW
cdiTBxaz/95BlUNvJBGaj6RrC0GyDlZF41OYlRYwQeeK+Tg9FiVE9ModZCrW0Apf
bqwjfJh7daGWudgUW23w4RPdb1vzquQvQxhpntAUkMTSf6JyGDqo2RrL17giOOqx
caX9KG9O4X6FrbKLIGaRzIGE8hBpi3q8W0jFuUg39k3t/D1T+jOM0A2FGjiT0yyX
VjGAroPA5rRuVzojI/42rg9RwewfZprVCT7TRDoLt4lwpcegRAV1E5ZNHNul6GVW
P7qqAJa+KgTMifcd8Cc2LF4z/3akTz+d0EwvqJsl6VZenWuBCmP5tXqbyVYMmIaT
TMy+YBJb48x0Og3WlJWCjqMwgSEBl+J94ATfqyQ8Hg1oNDssIfWezgK2fEg+w9rg
qtWUop60vrOrFHeb1vRPrjdCu1t5oLNdnwwJ6hHNStVtoGKMxDQXlZcEktqPx5l1
TU4kkAX5Llln6NFGewHyn9ij6oCFfjX4B2iLQKC1Z8bOTC3Tjfip8fDceJJ1OWfg
X1JkyKHbiHePf8gTGX1e6b5saonbMX56mMrgJAoHnis3k/Qg8fc8Bii8zWXes/54
NF+V+I3u4Gzd67aHllghb1DJl3hnlwSbSJLzEuxJ0ZQ9TixWz779rDRZaGz6A8cv
IMoE4Y0iSRr5bdClFCtc/GBVb7IsEam3Qp1bpZnjAY+VdnmYDCEEDEgqyjRd/mns
gcKqId/hasuuw3kMY+qUXaw+IwrKMZlwvsahIkkomd2rUtHhmlBUPRXu9QcGpvj2
7XItgkEdzbaXsO5Usr+tf6VP9L8tDaQ6oZ6wEqxzxVVk0BQbcrETa5daVIgK+2lU
B6UEa5EPzNrNsgtJLD8ZGtzdkF5Vi9UhEIwG9X+YVGK2KmUYx0bx6jAxuMEy/dSz
0g6ECGj1iq9lh5h9CUFvNdIFHK90WVI168TtbBA5SfffLLVlnCGE59BbbsQgx43P
f/C6PZIdkOtIy+d3q0GiNUbtw5G1J+QoO/ZatFglFi8kZcO7GSNWpejzFm00c11B
Nwi6tHqo+Rdw0eoskGlVuP9HssDxiZt1FxHHPphs8OlumeOTOAkiQNpN0RRPfKpR
Us3N52ja1gvub9DgWGLFvcuYWNdclvrc3L1xGEBRKvx+SK7N85X5GYx2b74yjvrp
BZ5Io1S+gxgJVhR2/F1VcmOlFwFGZhYxd8oJN9hplPZEEbqOcPZFf/ca20tO5/fh
jrarAU0YQwAwrc1Efk2LumKzsIYMCc/I6fP74bgFSxB4Kyi4QJFRv+ILTGKjrOf2
N5XuSxKp+gEJ5jHoRJGEN8kPHGCdgyTQ7GV9WURkKRTLB5WqAhQUe/EpvgPHIpTc
hXOjAPWCpNmv2PIU8iYtE/YHbvgSVPX7WMQAbUeUGcadLK2rL1Fqj5cNGhRbfRJS
XxU5b1maO/OcDSTXMSAIQlCtg3vIxoulvKZIlUmvXjomDydigjTOCmXzZ8JSbt26
VNZwQ0WPG2e32ke1nb8nf0m30MTDwI3As44Q8qYbuEcD1MNyc3lfG2uhyhyOhEgH
5eJXisrfNFUxbaNJoOJEMA1K9fxpWFSnKWY1s9undd8KqmCdKvxr8WyKNHwmVtw0
JULeRmcFLncAEYUuo7gerHEt9wio6aTXpGt4tpp2sOS3s2eo+Qt3qQHTiZeQxkQm
K71TdvHjpbIH/SYWSPWH/kILGVhdnBQWw7p6oY/1WizMCRDXmFjtmsdKTHtztEaP
AXbiLkyb7+mOYZR+m9s4ZkJO7qh07vNVs6xFVHcaY7BjF55jbHkLMQ4iLR8YrYti
IsASwgbDYpCsk7H9xi6glVamkjBCNxSMzheENTESYVru3VUqQCN3wTp8Q1TBMQM5
ydf3OeXt4qW07Tje3hBM3yrMUfKQZxaZ2HNKfa4TiuAh1rPTEJmNxMU9TzQhf2fB
e2nULgbiLt1oi6mXDY5NQIvxU5x0HYestNZYhrLEpIjBHZO5vDY4uCYzo2SjArJV
GQIWv33tfmJY1qj1aBR0+SfeYrl0vEkc8x0RAITQ0PIJBaZQUopAOTc0FfTa1E9D
vHZ3U2HCk1cMT2uXYVF/FbpTVH08LD6ThaDfjvoDN7cblhLJUzymHqsIsceV3Fdg
6XalbtPUPm/5kkO9Eqy3TFkSo/wgtOMNOpjmAIrlP2e72Sqy1phCQT5caGAGpT+q
rPkMT6OT157y4rXguk2RVWfiZ+GCk8yXnRylK7pih+Au3APDeP1KbT34UELDuMrE
6nIgJbV+tBI+uOcyGt5Yeei4jgF0q+xQOJub7ZOhhsKfwoOyf0eoMpf5un5I0wnO
UsPA3+L8uJ6FUD569GS6k5+88AiSHOwjmiHTrUUcV6EPgy12z1jGZ7cMl1CZPE5W
hcD3lyqHbQerXpbhpv335eGfSEko7/qPK2xRZx3mobITWAUNsY7L3LOnJr0cUZgn
PU+0a61T8hIgFrhdUJrl40M79fYL3c+f30j/jY0j8vK8CxUebaSXx831VDbzXr9D
2VdttLvEBFc4G4JOISRPeksbfX+yQNVwuJwNBA96bluGcj35byYNAC0GCGHNdRzM
d388MuOj6pZHJMpyOJNkEgYL4zgK6RNbSIrZA1vTnjDyAWS3KLjWl35Ckp4eAHPX
/VXyIZNHTHeBmFIV2hv25Ko6rZ7I0f20cdNi4EgOclAzWt5Hgg9SIKrwypT8oQMG
f/jfhSNXzD3TQDwYAzqlH579PUHjZImnlNekU1fC/4UmP35WzFhh/69KUHieq3Ly
HuDO3jFtqVuQ271rZnJXxLNy+W0EB72SCfbFCSjuI9No1F2Ejtve2kROduah1sRV
bO1SpuLAnTDkHd/IW50CD8yQqc9juJBZnOvBKkRK8hOT4KXESzgl9sLWmjxqKtHq
ZZlicm0Ka+DbvGD/gz682A8GbzKn2J8nY1UzWr82jt9kCeUGMXJbIILxMRZmQrrl
zpRuYod0GjT+N5OsO71XezPdt9B/msVeoki6zN1n9OfQv2+5y+hRyPP9VTn0uuSw
cCqvu8vfPXOf8LoqKkpF0A+snUiZqZztQi1xOfpafmEhG6xGsNAjx/OaEbaSMVtW
iWuphhcodw7CIv63VHI6QEH6PZa4BRc8rWHMTwBEQAiheRS7kX3TsZK+flGLFTIF
/elFu/Gea2kFIYfAKngf4wDpWWx/idLOepdZT3pn4xShLG3usnuAEHkYFbeLPXUP
fdh/NlCoy1fekNMPZJQZa1+ZXhaD/mjNenm0GHcupT91nAInFuM4cH5k5jXcfliT
/Si0eFucz8fZd7MrgJJH1PGQPvklsntmOmYD2IeX8guydhL8gqwbl/lGisHdwKrx
sh8MOYrBHggKqC7IaX7rwiv0FvGpxvkzQrFYIrbH/eIxtBdEqtxyPiFkD3MSWUK5
NrjqOovvN9HzJu3k6R3ufbiz7Y0vm5/zPqUh+JYnM/FL0jbEAKTndjUEYVb65lHk
eV0uLz1zds8YTb2tnxfyOBoM1E5ZaK4YWyET/+Uu/Utrcj4iuhbgJgLe5CHMca1S
T0YKIaUAehd02QUZhUpazKKeiFBUxyx267ilOu0Y/fosJiazguG4p5tZDL71qqZG
JKeqtejikasYgwNtQYQ5ThnzBt+zQ6PwzzXOyGgSQLfrciN9hLgyd0gje1FMrAqd
Rye9iTCuTT1VbnoIi52UMHSxlTKIbNBwyvrTI0OLLOgCppykh6JjTsmG90Xgkb81
iDjZDIXIDnJ8WORVCezaVOdUZFcGS132X6lHV0V9Q9KdNB0lyiMsBEEe1KKOkAeZ
WyKIlN9I8zrEgX2IP3mfq59CaGQyAAlCb6cla6mhbl7N9OiZAORHYMhHlchv2tKg
IK7Imc/EvvIKSyR8WprZ1AKcUogBB16N9yzJoGmWAhmuiBGePQ674HMYxamrlU+V
w2EBv2xGdx9Y9fVmEvUWWywU6Bnu63Cj/Jb0JUON8PtNgk19sQA5HZe8UEqbT2MT
4w0w5o9CuYS053umQeMFilI+OrU0LRAr6/A73m/LjaLWuyAmf/KNVXU1cPFDUmcb
MBbhfxP1bXerQl/PXx4fdSNzF/QODYnwu6MsyOSOx6E8tNixKc3Ryv/JBfjRqLR3
UNDTJk9zZ+BuBLrB4I2gOCxKbFQQ4AEsQxbIFgbsuh0GcFsvx6R/DKEbXljhGIP9
QeLNEjU04OvpTQZRI+WwjY+Q1XnUiv3q9x/zWmx21qiczruoN3Aicu1GQwdHhs8j
SPeMeiIqA11LB5iu1HAK2RBf99fmAOFh+YqeEGb7Kpi/voKUmv8LrfB8x3+o8i7Q
PRmNloX0gBoiLyrh+hfLVJSSIPZQmlaXSBh5ZFhZZL3bw9J1pUoWA562EQaX8WFI
+AFvEPUlXV+wk0RLY3xh4VqUTk4hkGZFcQ+FWszx0cQUfhZQrDq3tj/5WkBIIbvM
+ECCETXkhth+d1tvOf4mPMDMu/5PsqmlMeVVAcIdf/Fp6ecoe3MEyz59fdkhtzGf
NFdNIt3iQDWr87lld4U7lyKUKmtTVIZaWH58uhqLwUHHSlZ6CtAnNn4sHjV3cX9m
FW2oUpjRaTlvBoNXwFCEdIgnqQQSIxQPFDf1+EGExMZ0PI99ll7lcbeFkHfiM6ux
cVr2LlQv/5YZqZXixBAiBC34gOkfAJDugmJ4uiUsfQzP4JBj746deA9d00ii8e4M
RGyYxYJPSSm1XVZ2YlIQWLBbjOhNxwdwA9i8k4t+3F5QO9YSRB3Ten/wEoJ7t0nm
3p7Jr4o1ss088Jg/a3Fj8o01RvOKbyacYTGZHKPQYQTESWpcSOKs7cmL/7XEaziB
xg8Vk0u9Jq/+9kL3TTP+X4ee0Wo3b7KxYNNRjfELx38GRhN7xRSKJlMBrhZsaI4U
P9uqXs4aFHkd/n+x7VEc+35cRLzF0lI4YnPLwHLw51Ae8GyCY+GO5cDA8DCh3YJB
zpLCMUG5myi1faxOjc/RLHUa/+ZD/wEBbuKSrsNjy6Dy4MnvdLW0w5vk4OGtYilp
IKvF5hPS+CWxx4uBMUp9QXKkeODmpFXnO55TbNwIMy49kKmDjyF7yrqOBKlWZdqU
xRfQHFIhK61WNfSjbENdifMhgmtUM+qxSdYgZDAzyVv/U3cswZE5edMf8Ru7LA6i
Azhuf+5OJfCUi/+z5BOlxG3c/ed3lJrLny4zml7lDsFEWBKYTI9yehEpMKaUqFIm
22mHaJZQvFVn1tb8H9Hdx6uFHT/qMoVNZan2QGU6Mfa+JpEdQc2IvcO4yEfGEP9Q
jrKcjJL2GGOtftnqAZCDQHKsSepkFD8AbMf5NvVYAULITv3G+dGAn/4jYj1eLoEP
wc/OzS2ldntkzOvjRey994D6xvmJu0lhk/PWgSjwQlPwrAhffiLU01q1VFvuZASX
JdK0v0K0nLUVR0jdOIyCNVWrZQ1MP1mwvaVFSD8ZX0mDFKysZlM3sNLpZMzbI32V
3RFanUx7IWsytCbZdJKhk7meaJtn5gP1iFMUqyvg2k969N1T100ScrsIYpFMcqhb
5MMcj2MbyfUnYWtDWVbSnb6ps/2G2QvVZ2jLha4GL+h/gLtlLhpnuoJy41Ay/Pm2
bJnFCOh3LUlO/OGS4goQoJ8eRPoCqFMwiFVKUL1ZfmRBjQA+kqBk+t9Qio6XlBwf
5WRC0jWBaMevjKO3APo6zD9z9mEn4w5QCCiWf8O/1njD4YnRsfLOzhuZNVidWcDU
V8RUdQDUU5ySO7bI17n7iylQnnHaCWCsa0AuR2h7BcaFZg/Xdf/uKn3OYrSdQw5t
RSSNllsBccr4vJckQ5kkeKciIx2Kb6m3Of/mj4ElloUuqLkN7nqgknSOrwQ54Ytq
zUO733jN9EvtUlUbaRiIvyUe57MRIF8sGG243Kozw2Mb9GdrZ3p5Nm70aw099HnP
NkP/zVI3g5/UqzWoOMXQPAbhCWE2Fp6ndxjaFF2A90/LOnnluTNA7SiXCuWqjmjk
OA7GGKkf/XPXzI+HEYUFqmn9MvisDJ12y0u9tOzxTr50kyC9JVGN/shx+tTvaWZS
dU3AhbpU0TqaOjtbmdyBZ3Z4LiHRg1OPOUAiiasaH2Q11d0hQU515t48kl4VxQxN
aKdYfWM6h3GzXfQlXfKl9tE6V8fl/fV3ukHss/RPtadSXWQwSPk9ihzz9on+4+OU
NAUC9h1OowQ9M0h0dwi9+FzWCm3vaIoDf87vfMU/qUmoubbyo8p6NCU3igOKu2dG
SNHHgubdCgbifxJC3nw3sjNUsLL60uveEDDDhGU7sS3rV7caQApzWQBn5aOPgI+U
gVy9k6z3A0LCUm5R9mg+koLsFLLODjZq5kP9AJ4Oi7oLGOe6MlZXU7Ga5+Nkca1F
LIps+nPQyApMAQUXwfSYUMV/BOtN3foLY64WKT7EUVZoERtjdN6fJ+llseyWpbYa
z1Eif33ASgj4a5WEe1w1qzpOD/UZo9cZo1xq2URLXE4bZ09N2o5ErweVD4rcHErV
DLykuhgbxgL8dsN0upj/n4YBhYZoTgc2+EJGuFfpApQZobFq+ysK45uOdchixMEK
HtV9V+M6V6vxrOk4/M5qJXlLnKm845XgLImFrmvxyZHidhNjyhEy0fhWtL9T+AMm
zhWmNKnlsfyGDOTZBkATW4shRRZsW7r4krWZaLqOxSehW1swligeAnIZlysWihpL
jVB3j3DIbqE+FfTpc3JYTLLHC3eKxH4M/PWAWnduKxJP1Ab/lalMF8adlVkKdH1k
hvG8/cpfMiM2Y+5ohMlcHtB6wjEs+Gz4WfCFjQZKQ9GadS+HIr3MyrAFCKsJxoC1
WS+u9Y2e98/eXe2eeXHS0mKDB/Ec2w+ai3WDO15aqL3RH++tpKd3YVM8ttgQlo4c
7Ck2cP3v2uKLcl96UeolIOwDKfYB5Iy5KOUYtcY0ae/ktPx+zGO104Ti1w9vsXL0
Dd1jNhqMy5/M5KFq9KzxdprTmkatRVcrSLnTIwnvRgletCrXAYYqmir5XqaovjRY
TBnG1UIRR6RsLUL0Z21ZfHUIEmwR+lIBrI49h1sYKHeeJ4qbMc+16hqkSFy4JNOF
I/RzHKUGNnhmN27pK0jmmYMYSVlY45ug7hS+ODt+kKIckjUefyQxEJ2kaVkX1tsr
rVdl0Vdmkv4BbhGv9G6Y4H3icART41YhXSFGUISVywG/0/pfMZQNK79ibOv4nbiu
j+uJg7/S7ntN3Qk0QD3tu2L7xLdCyVcE4ugUbV3gp3ah1GMj3NvZx+sj5PWhYlTQ
q84eKHKUdQ2ElUv18lQhCbLdFjf0fFXKqrYusWm1j9WD9pi5HBP3naC0AkAEj1zi
rc1va4hpFIGzv8xJFobGkH4co0d8rtFOrtdDMWv92dSuJ1fuycuAnSh+t4zhg5UE
aW8SYrLsenk/o+JcUYKG3m30RvKcPRjvjex/mqJhoUe/Tm8U2nJQrUZ7QzwqGN6z
lrykg85d+y9l4Kpg1PZSg6zKbLkhmVXm+OtD7p/69qV7sf7uTE9ito0BfjEu6Mkh
mqdl22aXc5axbep7ka0ZIu1hdRUCiriZOAMPA3j5FNGCk219VzuxiyyCEvhBgTiP
6ppIKrxqsOAPRPR1UWaV2W+f3nyGF8sY0u/+uAwDpV2H9RZQhXL1QOolltzPI1yf
AkBTgbp1JUIc/QbROFhiMKlga0l0ZgJU9Ntr3gq96iB7wZ36EGE10rU/CLbKhuqK
P8uLdGQANyZUeQ1qc3RgIxng8zBvuO+ZaWfl5aVcguQl5tucHuobWsmjfhzpH3S3
tuG9I9xK2xBAc0eZhMTxOPw1Hy9BFOksEFUbBcKl2UVYqor3BX7xpqBUR8CvU1Xn
i93/yMnQPqXn/n9uDWl6LJg+TM30+/Ms/ppGuRRzCwMo2DpQPubqP4CYnCZNrxtw
6faEvqf214f7JvWW0sZI8QOi+7aLb4CiuTFDvqyjgW894mzDDWecEsIiTsDrB4Ym
+EEdJgvKgoI+Ii7WMKExgf4gXlzRxlPGxouoGE3lS+XaMeboC2moaWjSbfGfU6jU
S5niYRnSivhnLlCeoJvRhiv98qqd3/QsH8pUMdUnNFe/W7qVW+j0o+sKcvkjWYzQ
YlUIcmvw4Nw1w2QEg6gtFbev4G5OUzmuEXOivoUoSBa9ej27Ga8kIRn3S/HZ1mPB
5ow8KBdVDQvR/dyJ3HQ0KGXGlLfAZmuaZ9ItXdgLBV5jcN42RQEL4DAWBglsNMCZ
id7zHX9Jv3XbXAoyfe02daW9Zq6adKHOLymOlNG9s2Dyw3RecbBh2LKMv+WXFgAn
4a/W8E9YW2INzajE5O3p+b91YLCyQUGJphogHhyT69ECGuZKlF4cYnwVlxS0qQVG
lBA2BzsaNo6EqBv4myDRM1aSsR2ZR3MVSo9JccWxnKNxnaMVQ7ZBsDsyHeI6li6O
jOhDKlO78G5ADhOEDnBKtT5cFpXC0FVvXBmw2M+BEWW/s7NW75WQodShVTwCp5mk
tNamvFeVT5ds6gPohRfmYP8qdIMM/MkPLgqd+dZYmhvHFtRJcLz/r0CO9MO2pQji
aa9MNecS7PJH1OOqsmJH10dXPoVD+aPpiq8oVCDtfxUQIi54vIxclAugMHMtyRVN
r+e+CtAUI3LH5Mh5u4Q5Kqgk7mRBTFMmeJQUN4QbMl7Z/nO6Lm8WX1rVzHIrYNQ5
3s1Ir29WQn1tbqP48WbwVOICsUbsWR0GXDErCHL7bR1Cqg/05HeHRZ8KILgotUTn
it7bdNIlHagvm+OUxCs0GaMrZXrDcSUi1px+Ho5JHhNAQ4LMTa8ivUS9aAXaGZp9
GbdQBWJkQh+W+qjbL/TvM1tlxekcP8+u/yjQnzc+8Zt1FBbrABTACffegPZVbYFx
P5nuHXxheK4mzuUGz5NFnUPan1LaGARu+KZvHMlQftlLMIAfVbt0QJrnoHOzSwLm
1t668WubTPG5K6VGni79q+3ooRIuCty01D5fDxx7Hg+ozzG8wd7bcMmNVrsT5azc
sTZcwS2w4cDWwgA4TIct/d4eZawHWRIlnCxsJojMYkl2B/qPR6e+6WrCoqKG2+PS
QV9yocexK/cYE2OtL4rvCCc+4FSCCbErBfnz5RnYAe6ntLmxBAQlEu9e6wQg89Nk
8jaV8PWwjRfjuRKRe95w9hMvjzc/MvqkU7mhpx7XplatZa9wK9Iuvre86oJ4PENg
aodA6a5kYwdlZT8gBvRsoi0qMAxu4AZ5zPC1C+VYMILVU24kovmBIIxInPfM4bcB
difh5WD7tAj5YR6sJ7jdNX1n2uB/aDF/5DoCaTT83hKbJD/8TQL9+XAPkLdNa93P
U5z9zrSUZJGaDW4YIutz9XA/07qBNOm2+RfI+TCuBMNJHayexTxZTnYZZ51zevTI
CqGw6vueMfLszflBUtBz2hmqaR7+fAFjnEaSkJmsU8PHfZ/AA0H6wsTKCtqd2JKb
PbPTHhPoHgGk4nIXgjVh1j5o09Cq7hTr2taZmlsSht5QaaEtv5slZk1GGu+DtkLu
tyCzB3pPWBRvaHb8Ft8F6315K5kPGQGQD/4BHzKMjZfyzWzUQDQfKWOB3BBBXMGi
EmMuqH/Ei1KI/84VO0kW+Rcq4Lvl9po7SP5cDZs0uBrKmId3FrtJYkMx2ET9joTA
32FKwN2b8P5cvhAJBEn/CswDaVp2Ynfhxox5UQaLYeDsbfsHeXwjxDdfuwySa0iH
yUoTgCvL/gzDTaWVMkgEnh/EUwIOT7xk0GPuaXhxiYkPZiEdOHu+4eWzNhKnPf+B
SOwd/JqHQWrKoRFB2WQ/PI5epf1Z8wKONNjHEPyx77/ThAspV8EAHXnsmVUk521U
BDI/X8DGniScxiHiVciIoID1bS36VG+JOXAsr2YqlOJd34Gk9TDc9NJr14a/C8cM
lM0Ad7rgwLAXQtcv3fTRFhMhnKWKUDj/mPtTWVROs8hInHQyuLcbq+ehQyHWZr0b
LmQqHEOaCuUMkpWpDdV5htd+MWzfMh45ywsi3HRB96NQacDdt/yc6KkDrKr4Fwu4
1ZbmK3hy5aXwO1LX3ZKZ9Oks1hMPt0lEFh1b1yv1o9N90/hQS9rE+OOiYbO2ptx2
XjgitGl7m5aMx/xRpKVAqOFPpGyCiWUkS6s0uoOc5vbcGmKXRryQXuu3MTz0Gfin
29Z1GNPDA0b9Gb8tAz1AaEIuO6uhAciRUeHlN+rG6wJ4VE00iet5lJMT/j47g+ZD
Q+8++TEXJNZ3DlL7cZpZDY9xS0lEP6Bmz5G2W4OVcrE9VguGaOo2KUoNiEBr64pV
QBT5OctcHIhe4HAbXn8Qo3cnNZ6Ne/N6kyz91bzYt7VfnGbM0uAR9Syiky/0T8i5
xJOOiNaM5zt53qxq2ZOHHjgZplUnUUfdbwKXPWi4RK4VJ+uVHQ4g0FkGiaDhR1/j
v3Tr2JsN68ClxkSmFwabZ+j4CpXIDd10YcyETjQq7T+F7coo4XfzPdVFrzF+ZXf8
vR1+/bT+Jlouhb1dJGd0qLSsG8IsOAAJcnX2xXwAz1wzz+H3RZbG/qepAyXJa/SZ
JhRv81GQJ9CYSEFcEE0Q7riplUxnnPNn77E3nYcR2KNIhbVyPGVm4StuzqYz8v0E
ZGw3puVy8KnyCgZV4Kxe8r6IAnY50gRZMTppYaWJIRLPCiQcR9vhfpB7y6YKE2Cd
0nlFG1REml7V6AeTjzuFmX+G05TQ3QG50aKbq1x6vOoT8sjwMC1+jRHqvZ9wNnPI
A1AwGxnS6aoOZKXB9CuUpuJG9oMUnIR/ywqLZ1pthO80JeEwGsQAM8J6TV7vd7ef
6vE1OaXpF/AlyYSrXodVUnMIgrrPiaywG/1CNiW7LormGTG1e0gfsk1RKIaQFq5E
aPp66Zuq8bVGeEmYiJqf9WAUugiiqmTLIKOpVHxKqDRhh7tIUpYed8JkcpGSSXQ0
yR7f6HwzoIgLxqkCP879uw8OiXRVauUDSv1wb2WAm34R3k0KPtiq3pQtlykHrfAx
7fc76nej6Z2y2EjJ0ZZQafZxaqpZ4pGD1poJIlFrE/zvG/nLZqweOL0Ac+pH2UKA
hk0hxaj1136py5Isx7/wftyFGCnTEdMdZMZ0JiGtxnlJfXvral6gTdIFEs1u49LH
FO4LCUjnC7hn6Tngn5TApl+ih7NRoVbd2e3MdyoUNo6j8zA4Zbgl602DTK0b7kSJ
eNaFNK4JnwugrZnrxeFINeDvI9+AtCGQb6bDe8lMzsNRZ8Ua7DXwe14g6GLun/6z
ZGgOmoHaZ+Jsv3ziB0RAZkEci7UXSgWrucq04t+LsyNflefZxu28dKJz8R4c2tJ6
217YnJsa2p2umtZAoEAbq6BLrZJhd2PoyGqgefsF+1TucwI//JDsmaOY3KNu2MNu
AK+8Y9Mn1rr1R4VPxKCjjXhEmb7Ns+5WQKd1m38VBm+NbuiF3bqxcQ+YOAb1hLDb
OaAU9apFAZjzL30KeDbraiFPGBFp0TxijZ9M9qHe55Z2PHyhWnRi1bCRcwZR20MM
s4/se9NTTpA72M9ZKbdx868YdN5JDGAXNH+o5TlpgbSOVIPEcvt42VgmwpYxgX/r
2fCg8BLLop51aTHl8dptX/Y25LdCZyrSbjVlB8VBGoVliomVCEkbeduXKYEkWEoL
audULcar8lV7OigJQvEXv0DyiyFanVlnTzDdCjkVws1EWE0dg87KNvzHWkpIkFev
dwreT3fJxHmrW0uiSv3XZVmUQNOEY2SvyQWIfcbr7wHSqdmDA14/5a2CZyoAegjm
C/EO6/C3f1Ff1ED2yhvgdQttAZDbecOx2KyMeAZQUXO+KiCwLLduyr2zRXcmClNS
I74nfmiA89fuCGMcO40TtzyTk2vbnmWYbJRdMJzTX31FCN+zhnqvBgGtSQLMvGsB
4W+nt6CQ4+Mc87zDORSfaqtwdbLBhVV52p8gtKW1jICc5oCiSzvz7fKFF4hnpj9A
48k3E38Chj7sYiH3IYy4rgkcKXw+M4k2N+1aBmXiqFSnwt3dd1NIDIM1qyiWV1gB
p5C+qF/vlHsRfKxRjuS9YyLWkPziQPWuo3Cr2QziRTFdXjayR7bvSnnXbSBNJB43
VoJcOe9J37uWp9Ew8ZIDmeYPiJnVurS+ir1Axyo7V0Ie/TRO2KwYi9RZGbEqf8gF
6E5p+cXNvUmgoRmIgKVeO5+mWoe4sMGROMXip7WdQmBeYKj9xXackFUUU8udWAuZ
pAQQB0JAEWTJ8kUAPVO95gTr1KSW2rrNCJplnstm4KYdoFxMdimv2wEImRK2xo5B
C55cOtkwt/GA9XHNef22cuDyTaARAweTb/enzEIgQ71kL9nyXrgixc7x3pHy1tKv
Ay9J/9fvuP2C8cBZVKSGkySLRvIbTLz92YyvzrXHEl7p+TgvZ3GeXni63VlStCa8
0n+uC4j8R0B38u5ZwLT+blRH5DesVcw0ZUnuwwHE4VR1L5W1D55ZDMbWcYyg90ZT
vmVtKtc/wizoDkYkC0SwMn1xsaDUw/UZ4E6sE+Vn1K8LKQQPGgrMi1PD0dCoU0Ey
s+kjwu/CpMNgxP/uVpIux37GW+f8wRvNP9KHcU/vI6ZvpzcyNMpM+uWFlxj5UxlI
M/cEgEgqyu9PCrZqFcdNLGasdWT/3eGO3x5QqLSIj5HVeo5QmhIhJMMVmKWgzyrA
tJl61swh9YJ9T1IM4vO9OUVY6FdJGuG+eQUvVJrmHemdYI1K5d/Uk9MR/7TSMBR8
gCME5bXfeUndc6BiO/edfFOdm7A+UounyMdd2uDyf7nIPmoiURcSZ3rpwklXhZtU
Z8khVmzzd/WR1OEfyBfZ+AqSy1lMfFC9m1Dx1DzJTkvtyrZgnR3qcATIKPoY4QlO
Jo/Te21eqmOxwgJUsTjGwqYh9gXe2jAmkb+XUmIVixZmS0STUz558rHhluaGD3xk
NAzLCwXMPXxQ2FIAVk6R5Vp9S+2D8/DWeLDY59xmcmOvmML3Ldf5hsFICbgeFMKI
oNKTmsM9FfwFzB+jOkH5HnKvDQxY5rsBXgtlwXD+RrlmCKPa9FeH6pVoXCsJW0R9
xfPinvmWw9gTi4GqB2jJ3HNQBIquRWvIH5Srw9xBhJQ1uvk31bBn08cbP/DJHX5B
Pz25gn+JXhIxqJ9BxTDXSxXIpBn07ChQr8wSFhs5CVwwvwQKFDwhfQV5dPk5m2Me
kPlvBnzVOGRWnYo8+UNmaUtgY+FQYz/Wk2z8/VNw1DJ5PgrJmySHSJp1iT4wsXRp
iWPzlrLJlIaEyQALAI8qMLcatPja2Dux3ChEshuC0Xpfi4gHf6AuVEqBGPj272KJ
5onYl/ibaos4odnb77kyFQgln5dLUfFnou/IjG1O1+byqR53i+dPOa2Qy+dS5rOf
CCehpq6wEL25PJeVg+HW+2pj24edc36NzqWuXUz7XLlAB24M8uRSv6Qd9lU9WWEO
pyIA4BCovIEO/9nLK3W5WHVZDRsu4UNDZFDe9htTK1sEOdxEvFahFoBHJLejFOy4
E2z5lsyCBouCouZsU0FbD21ETr4bXhXZLuzS+EoN5kaz/0vRZ1ofyM5heUS4AvHn
Z0NyAlGBLkp8QWV4BtHFloLtUHc1EkbgGiIJQjQ9NnJErBshXSe9qJdiW4odd10H
ce4kJ1VlUItSw3LhKN92/l8DTsiYs47txdAOxsm9naQeRzOoa9dWFMpZ8aIIDrC9
DxlHtm724ts2MEFgu8hYfPZz3Yh53CKc9witdCX3OQqWYS6ex14dw0pOGybaZKK2
NCeDfSDmLEHjtlc5ctfNi5RbOLxW++Lw3VUPhq2BLPGh/9IAMz/0KHNN8FAObntk
o3mil4ru94srY8oEOsCEtK1dPr8rIKFPuEVM7s/SyWoKMJ0eEFQjP7CSeOIs8RZ1
AoB1PdXsLnxAkegEQ3/DGTd20qjDRqiU3QVnb3kx0MuBJ1svjLA7mA9WZcMY4KjP
5A0HIxWWeqaAzGltpnvHIclQobPf11eReQDV6/TEITLFjeJ8YL0GrFo9ykd9/8AO
NwbSRGwfHQRhSzVOkdaOJJKageWkmRb2+3muNEh6NlbCmKbidzsuaA7LWCR1R9v1
XdIVHMvO4T8ZQye2PtX5ilqT0VryGx7zqIujLhwlLJgXgVNJA3c6cMhgALU8Zr4l
ycSC1Bl0dHHf2WtgZMi6SDGzyCX1C3yEPwGadgfFH6II/rufYsCt0wsf9YzThmvj
RvgzqKeZc2g+tiVM3FeTxHBwcst+9ANbhf6402BWeQesqsVednONWMI4FPpX5Qjv
LXkAaTB3NnOeZ+1A8cC+wXgMRm4yZd4Fsu2QNathLv65U4MebQ/rdkrbol6WPQqT
jtTE3Z5n2lKupbJho0wbn7b4Ctr8aQK5YsWISu6gTOGwtTAr1P8cDPDAQ6BvPM7N
QHDeTHabALirc0w/MKRV5A3EBZYqKHgSYuJnmPRWBe55RK+RaiqBKKwu6B9xtWRx
9KkOusuK/Mv0LqaPqw2C2Xr0XnAHEuTVTj67NNUZoiLBpKcPsg8oNUSoCvC+Z2q6
9JVePWCE7ihq2lyKMMhHunS7ZFuGuoB9/ktGroSOsQBhbHINfd6myR/fSUjcscCw
8mcgkYjRrBok2FTadsfjcntiCOeOn/l1IV1gyfoZq5qTP0DIaqAcPvjz0j3BO9GJ
O7bFf3cE5I7aSCRcapUs2cxBx78LrPttdbKMOZgOjDH0b/1VqvJi59cpOW3DtKIw
q37h+ib3IktFSBMI+jWLprm527NI5CBd7dHv5Y/QuGgTHujPJqaACT5SlwT6Fs0f
lMGSHp8sPrK9W6xfC0FNU9SkLiN7Y9O8m9vMYZAbw0yJTWeb4GjO+RNMpzJ77DEr
orAAOW48BCCLbF/OKbAvdV+1MEPdGf9Ph8wR9Jic0A4M4wS3E9e28Ks45QCMrvsN
Yv6J4D5NzecOlRocsGyxpzPK+jbuDHH/xMVb8Ae6xiFzGMwAvWv/YkQiMNSerbN5
AR06svRfFTrwk6qhYhey5nSHWws//8rrCyhHbbfEYs1Ji9TXMEJvlhuUzOOM8DSa
RoOtCaqXzUyxbwz4dYdbWq6JdmRc8Juuun4WHHPRuC+K7qGu0whgxuEe5HtQnZrx
yUYCjsp4uT5H/yv920/f9Z+TCQAKYK1VEKwwW/UBWKZ2sqo5paz/fnUAeum7H8HI
pYaBxujrdfQzzj2+4ddD+kPMj1l3JWNntHt5Ay5KDkYv8VZK5OFjc215ztPQvjmX
0Y7hWmxuk7rnDsArqV3F4U51jo0omJj6rE0Hc75gfMTsYDWqoWeWrwog8GvcKbXD
P3emexMY22DBh7RrkEMDf7X/dzpdbKpk5Ojg1YbptKoI1L5OFQs8f2Qc5yy3CToM
yRFDocLeGKLjvziyTsIeyNZ9p0OwJILCPHmb+QLNvyDsAU6jVFKq6rlZggktQWBw
ZrftrCr1R083T97dOhtYfxNErLRDZHTJ0SpOnXO09gJ875xtWK/ECbFWzQGgLZLM
7Opi1OnLhQoxBNY8eYPSmOzQHaNqkGW6PaKixPijPW/dk+v8arlvXTnJEoDak4xB
yvfODok61oK7Zup9ofHfFBnXGGdnExnNOp8en1R2eGUfSipapRfqvjVh4o1agqxg
e6kh3jY1d4L+S+p4wDdqueHnFF78d66CRGR8WQzTkP+l5EqJp09d3ZmmDG/neDao
bYsG0NmR2wdRxWjgXlkLUyMLdw59XgEhvfBuDtCszL3m8q5XXM9emgXcEV//ps3U
0BQ7U3T/HtgfbFF4dB4DFJDsM1Ubuxj632Tky0W8ubJ7bCGnHA1obtBMZnmCQDYp
knKwbTSzNg+Ye3rOdeaz+MyS7hBTU4nJHamUlqiG07KqCh/yH3+lIDcFMIqnmBls
whmsIMpxqeT/cwoqDxg6WwP1T3GkYAsiGm9pyHapXP1BNMPmjkEK8hYaNoTpoC1l
Xi4IGGUATtEtYZPby2pr+SgF8wXBcOHrYExGXjTP/NMqlhvkOz8Ywl3OzY+D04np
5HnBK5FD2Rhdb1qTMt/0zyHBRY8aGZp2o3d+WYxcNv+BztsxHE4rHN9tdNQXsn3q
SFxTvHL4dSelDAVT3Vt4mgnDKgygFeWb0S2sYCAVlDuD9ZeIVErrZdByhc5XQ010
KKwFpZwyBsIOPELTnQS7eGnFwh1pfnxTng2wxMNvKcreMYYgwmS6F8egOPLb9Jh9
SIgsAXDcu3ecr4kirQSfw+ZMz8GxsjXn0S2Dq7msbjPTZ06rQYCgH0C+IDnWkfkM
Hr01FzGIOf4Py6BENPC4kTkbSDbo/EI+g1FuB6KMnoa4rTRUhTdkU7l+bvUbtdNM
y+AaX84ltVb5vM5QyQ2lMVMGuwdsZmuNtPemi96G/SeKK8mKU3Jy0yvSyWWC8Wd/
mHR3B0ZgYjhV7GVZK3ppTcb0JBFBX9mGedCEYDloXBQWxuMWXxYgEr9IpoR4gfCS
+14MGInUhprMzeqGRjw+jz/+Ysxzak/xV6bzIr0g9cN9BDNlkrDR85v1xO/6l1T+
iyQlXXh0hKecSBSQBtwPtrpar35+6BuXHBKYrREXQPU7XNrxifLxCq24l81ulRS1
J4KcO1iTsphJqvG4IgqDc0kU7Ms7rIgjstfX4DAFrlI2XtRwtKsEjpEFywofBtM7
rLNuFPmSIxuXZvLkjS6/+4GvmAiS57PGVYctB7aiFvKq87/i6OT+uNAMG3zDE/er
sItY0ObVyUYN5XfP7C7/8FmmLc9Q8IDTeGvqNGm2qVOfoK1sA9178BJyxxSK0kDT
OqtyeS7NlwfoJEkSnz8seYm+3PqMRMWNV+Z0kmbf3CuLui756HNxJqmMXV224qWf
oyd1cq4dQ8+lwaLVeu3MDBdhB1rut0M2DGGJA9z3cQDuLfG6IADHqGegVkfIrtLc
Oa35zhtWIZM6irbtKo782GvP1mT3uUdEsdcum52yloUwge5WGdVYGpiQZhBgE3xh
bMK8m6T9KIaqEKj3bz/sq+m2cosZ3kMb4LlaTb76nalXRf0DtFgqbyBSUFC4n+0s
yXsOd9JdoCSIxGiJpuwPaGqQonSn+Wz1YvBbqDcLThtPrXBarQ4Y8Dq2Lb6ltNHo
B+CbQz56fWq9MHOJ+MPutfxXmZpjW1H6k6NTyC1MynCt8M33XX5cDHSMZTKaCFnT
5HXNnkmJRqXh9cDDh9PzEkM+o3+UZ3gcm1qMvv66M7IsKjpTK5i2F0yFNA+IFhuL
jAs1t52/IDbP+dXYCHt1VW1u3XuEYUUHJuyZ/r6I9suqkl9EkWfCct94FsCD/CqN
GuQaIuW/1iH0SLApZigP6vMSpC2sRE8ThEwHbvHiHhtnN0kaLjOGnueHdEw5zDVA
fhaZrkRETiIZT+w9CJVzln5NzoQ6XPeeghCl1zq2uaLmRsl9jQ0nZCc949quDrH/
1T/l7yly+4X5+0BLyq2avA0ldXhMdjN7L0Spqhy+93zLVKqiw9JasuLCDM0MQHq0
LJtWNBYPkzzHBEBwQ2G6gi+Y8MN6ryVp8ddR2oaTeAiN2IIgpO3GyOkLO8QS6kaO
5LzFirTcHlhi+MCGK288Ow11x7jDRwozsPYfwkvL/kIA1NzZ/BYbTt2Re969UAUA
HAgyydSuxuy2aXGFO9PBcoCysWT7FHNcE0f85aILTV+GBD3G7AaiU8jju9YCUYbf
OdzhqQcT3FbJEE9jbW0eSIlIj0QeTmncj3L/y5rEDcPNBdPfVgAh06xm9JnU+pxD
+YcYJGBVv8vV5mGEAITQvnhNOA0EONEUxcp67dYZViIi2p6NpeSj5pl4FMDDBBxC
AmENXMVTHu9Xz5fdRsxc4qqomhKcfQ+bi7IvsppdbyJFqeCLapUHx8yX5XKzJSbW
nitnc4XfQvAUxVPC2Dwk1uff34E4n2DB4r49PFLRHpw0G1kSTYh/sum8IzI6Fsxj
9eHyBLQ+yBtAyXHZIOg1eXloxnhetLKQOh/EAY8c+aN/zRiPzfr8CqkuTd8XY/JD
0d4bxtlmSfHvT8H0aCNQza1/2jcHfkQ0ZyXliCeK0NwK3Bb9hqPAS3KlogSBENjS
z6d8A8iYobW2BMCmDLonTEX5+j8cO5ReEQCTO/PJzqYEV+b/syMZordj0rWai9RA
cmRuuzdbo2A6wcoeWAoPHs+6JBjDqTDbCR1RoDhLIpFRaApPzN+4sa/bq404dTg6
H+N+ANFWYPL1r3/zRBYyO23dIcuc/Aj1mBHJjV69emKHYYDafRmNsy1WWnQjKJUK
kgg5LdA6x8E4vHynD+0I0LKJTHGFOop+HHGD/hVT4mbJ5FNN+7X2njUCuNZO2Ak7
maW0OJYpM6WFQL7gA7eIPPEc+B184luX2mJYPDrGYNNv7JYK42yTC+Xazg7cmgS9
x2fUM9pt4J0dyXZuxFyJ2Z/NT6BkDZpgV5yChO7KnX2yXddJlCXyoctdba7h61J6
c3ogfVOZxciXHreucRfTC9GmwSrJi8+clUeztE6U1OrHInLUtnc2qRcu7Uok9p/2
bl1wefEDELMHrtJ5P6/YS3sX2RxC1zv5yjoo7zXVgG5HmRq445hAfd9oemR62UnS
Sv+uWWJe5BGSKifmqgA91NT+Ga2oGlVZkwjgbfNNXZ962v2FJaZOlIPZ6OGGGOcn
4fORADXT1Jex9IT5h56B2WimqR+CcCTd8T+3cY9bOC8HpiuZNYmn7mtQCdA5cSAa
haSBRtWUagBvEfV4dv32sVt2OVywQWUhXHJIN8bJfSDZg9DBGybqL4zspDmO3PAy
rb8H8ur0TZM+kJrnMO+DfFovwrikaWfStK5hjnOqzCGslvKmgWgTI7Xou2Yt3SGd
RpB+7Kp8KLMGOYOJiOfhsmPGmmCre2Xi0a4xHasiMUerRg4xLenJ+SoLNaoXK4Pj
fhgQSHdl+7C1S4sMUTTAsr+KQyX5rNo2m40qNGURIGhtkaFye5Cs6nijNJVJtXg5
fBKTtXlX+vIokns+VwuqMs1kGbVcc0KdMNnXl4rcWcHgsz2UJxLnIbKDQo8nzRBS
7Tyx+bG3Q1bx+axodq4zouUI7TSi/wA49pY/DPwCRJ9OrmSujehMe1TMeQasOlUF
mLP674Fcw2wFk7ePsmXnOLmsrMMn8r8p9Qbq7Ep0qTz5VRK+PrZS2uzGt4pjdj3V
jNDCmc0coqMg6LlRkJJLqory3whAxzoNlIM9rPmtYz2IUHA03Fq1Xef3k0LQtLgK
KX+oeO4rsYjCyVhFoRpsfzF2FZYmXkT0U5IJM4WMNOWiUVtQpWVotFOSLuGvEc96
R0ED3idnLl4rE79eHtovsFbOorrs0Z1ueZQkxaJ46eCJx+XI7uvXgbtxDWtTlkGM
UTLBZlfCPtc/EOZY0kKq5hPFanD6tlBBuL/ly4XtAs3EUaxHerH+KYUXRoM+QJNc
7iNLmWxGs4fMCLkvTLsh5MaUAOxcMXhuezBHi9hlbO7DTrgv9/MkH99cC5ezEuxp
0nh9GfDeUUjft0uNkU6+PrCxWzKH2StC1Fnl2KkwgLdbcvuW6NHBYBX4Xo3IgQQg
+F57CXtxLwUBRmRdbht2SkoN/TuKoDszoWAt1i509JVIr3mjO9xmahikDLCnL1nk
ol7IagS1O+7L8IAph2io/RVx56yu2OGRlM9zIy4ArQO3cRSotx1kurk/Uv76ZP4Z
i8WPefgXcIoACutbnobAj2iuKgb60EfZgTNoae0jN88vHSKjn5+Fdi7VLjA+Mo+n
L6w18TASpUrBHLrGFtLUMZm+FUEJxjwmzUi6wBeKEd3S2wMBe2XydOn6WpePwkhi
0g9BUzKCugKsT4I+d3XP6LKGt2W67nENd5s0Bsg4Mh19xht3HdgioiDAcaGBx9cy
X/WQY+tA0C1CcvRDnsKsS+1LT06jrHTPbwD9lisgWID5dNgKsM6OoR2r8ZBBNvaS
gD0Yvl5fb4HRYFzRriNzlOXYnNbdyVJ3rT93Rq/tyV0Dtc4611ndPF270FEXIkg+
GwHlp5hCsnOq/VaiMW6wtjx0IMidH/1VQ9D+NW6+eoIOPeLc5uAuITZKem4R1C59
oPYDf2kgPeX2JBXkbBctSH5iEXWmO3cNiNJ/933Kn4pIiMPZ/152BheOn4gjYe/b
7HkusrEBKWM0Qphe1wa4viW63IBShqhPzVGrhgVKPVvgwQn/CgGuVWAtZ5FS2bAc
o/YeAmCXrryRo0NcKjG3+M8/w6uKRQ26NidhjQ4q/xU/2IZdhsa7PMaMX36Vvzn1
4G72mdRT0WEAFgfnELRKR0UqNfTAZhrNMOiKZdwoGF6QxCtHVUcP6V3k4D5MaoTS
0pa5/3I5lC/XJmmd5wsPlfo/tXxko5IWa7s4+DT1jLUq983frPNSBmIhKMO6Ss1Z
NypxIBOOVp00kULHuol/ShPLYQAlIHuLS3924Z26+rexDb0y2vKVmaWn7RFxaV85
+NXalfXFvaNVNz9VPblqQfj6yPVjdMCIOsTamddJ+hndCw7f7PVZcBeZaL1WRrWb
Kpm+KLgBkeL/y++dDCG6cd8T8he1D55ab8+6Yd3KQmE22UgNG8HXrVS8um5NQDsP
emhkpzeQ4E339CcmHC+vJ93KMRWDMw18+qCsCJ/89uUnDXloWlH3TTZTPaDlZtsx
PODVQv8G3ps1EwuXgFUdzAbUcotp41vry+/ioyjX+E+8iGZe6CTOXfwWdUu1RrLc
1xqoLf9oXXFrsmVFgFtRdZ2BM4BTGb97qq93Z5bEyB+u8tlGBK3pS0kmguij5yv+
YFIxG2Uo3L7BIMzIRwCaIgfs6iCryKTML2MBSrKgNytXI49h6JXXZS0qEU7p9EdC
K55o0Omf39qsbjSV6tU8RizRMu+p6ZwH9RWDbwwSBvfmKE97n0KSzvHl8IauH9hv
7R9Anq3Mm3zbTtE8OpY5Tq9+LbT42VSwRbEcGFWRZZMDG6HghxfAo4WVystblsd7
FiW1JyGmEMssQ+IG8MnCgV42VmkuQOZUjSHuxzXG67zj2s/lVGUuLuYr9IYx1/MA
2RXTUA8dQimi53VAFXZQmLu9m3b/QWLrsRQh8uZM7PobtO6SJQ20xtzMcZz37bqQ
BvM/WBK09j5u5UQuVu4d+/poTDU4myO90mQjB30S/8wq+nLsKDUhtOOB6ETdC4vd
XTBGne4BHl9rKBClSmMppL+9cqvsbpqHA1aZm4s0dHCp+rZOMr7zUNtzuQO8gMKe
1FIJSHje56S+IWCuRUMHkohqDO42u0v7TOdyinpaj6XpfAL941bxa8Ijl8ChqGYS
KUUaTF0kP8GNA11q1YHOFnnL2UFNNzZr27tPOiVrtOlcA7awkmN7YAj2BQh5EbEk
QN0V3wmhzi3t7wpE64FPaQth3DoxLvDWSNUrWDnAfuy6dhPbEB0x4AbvEOwRXU5i
g2slH0N7dnuW6VaAlxcXAUyr5frHR/oW7MmJwriRVYxbbe41V63r/AUWpoMnWzlB
QAtKBXooFjcH3A4FQ8m50tCbbQbnQ1/H32UccxGNYXZtUZe4LVOpNjXJVgiKR0C4
j/ItAH2ryYodFGCDmAT6E208w89SHx1A15JlwaEO1hEuUsWGYPT/vtgt8hYZJgFB
vSLyMryTKOecm8gCDOsMYCXgB/v8Z57MwRs94OVZ7NFm79b2VNlq1wHJ+/VnFmfn
N02fLR1Vr98kDxe1W0prGQ08AfwSwFeZZc+2jrTjMHWQn84wlITe5EyW4ivASjMr
IAHsdFqaXKCTQr79bwxfZ6JW2aDy8lecda+8u/4ILh96A8AI58PtiVvz9ywv1eQe
cBbVysBB9UqXmujh+vXluZD+jiEQNTpTD0douJcKxfXj18WycZb9gBSHZONKQeWS
5PPfnR3nkpRZrXbI5pz57/y2F4Z1yF4l/5gYBtqbJ2Wq/vEEDLZ8vk0eo+K6lcQ4
tvQQlb08MT6vyGhtm80RvJLwE1o7wLjyibAQNo6RpZt9v7NipS/Af6VJ/aqWMfXa
hKC9iSPtdmQG3yaItTYJNvYiuGQ6BgqOmnXMEjxY3zH89Ys9HWAcqks7WIWmBOrz
IncGkEws4RJzLiBkiUhRvq2slGlm1NF0xMEukoT2VsK5+1NCxAxpiiQVKgkgS2A3
dNPzV/zHm+N6BrovN2yiRcuFwr/ueLZaxHBEkpVuhc9SKGUyXV4YWd+KQkxrw7Nh
mG+jz4kcoff5nI08m9at1LYtl0ptaQrUhqzzmaCGu0pJF0lEd+N0cPFpm+2k4X+j
cdDjgB0taAY+i/8CZZnoAomN+sUj4UkmaWYqrpgIgUJd8BTTVBTKN8SMeuNR9wfM
4YAdw4zBqKTGFjAA5jlousOjkK20fn7XziTBpyc48GvhVi0epUjlhxWVTqo//n8J
Y1bHlFfcaENFP/CBUmV2hS96HbGAa7Dbc1De2aqzAoSAOKsLu+KpaKFdJ3i1gK/H
TgEFD7RmDWGaKKmFzEYK32zwBGe7q8ASd5AKQM2SkujcuhdvinP/Fa/qmK0NlRN5
+fy4CNYE4U6NGA9T8FlZyBKj/1Ne5yAwLRUylGYJ65wHEMOTx69cAZjjQf8pt2m2
MSW6G0s6BwV625SNGiuEr2ZyoN2mNkVcjXw+b5+R41NrtiqPn1ALwATK+UkDOeIp
aHAa293V/5yMvjYV6+S1Rg5tDhEwmB9G4SPg1ZIATGUly7E5xtVqX4ye9lGYwqDb
PUXHDzJ9U/v2H7IIEq2o5O/ED7gcvehhbsysbN5Tuj4n+d37jDu1t3om5Esbn/IF
s7K2KlKun+h/cIAIL3FFhQxBHLORagYAZ/lgNo2tfAsnF8aWipoPuYeFQgKoqvw4
wBnK1dwZy7/A+xp6/5dcIooElFHQ7THkAzPd4YiO4dP3Y55emyV6RL1bmCHm8U6b
9yaNInPUqDO448M/HMt3Ao4V+aMineJKPTe8EJLlM2LETwnyN9T2DdRQf+v4y4M5
EGba55utdX7qw3SpnjbGVhoXeZQLutULvC1eT54MXMputCu1xTj1RzzkvikDPYd/
fdWIPn7x6Z9q6idj03feC09aoHRGynLY0VAbgUbg8mjrUn+l6d8U69pQkIGyIkqM
BRQ2q1bLCbY9gQQeKbv8cfZow1bJ7AZa7cwRZmEueC/SgRyhE2DSKJ7rUHhVFMap
jFjwWcQyaU+oKmD5LzO3XsFigIqVvMLCsOQlQUKRdsvf99QWv69zR8KUSl/cHqYr
7fOJFnbcRMNRDqTk2VHPJeeyz2UF095zOJo/m//hyjrd3xjAzwhvISRuu9f8QbxY
7VrOEYp/WZnSTnQidR7K1V+rz+N5jpP+1mgrvd84DW4vXkQXMMJ9moS3J2pI0PDk
U4zJVEG2DZen3/19a91dKaopsh/ChRiASyrvGWViNtjW/w63tM8k0VIHOtXk/9q9
A+9ZQpXEwIDWWqMM6vjjpsTfgLi34desajeJlpxE4EyWtnXVi+dTHyyumIQQ7j6f
hIM7O79Ih78UecY0XJaWcFY6JoyjvqXfL3ZUyMQM2nVB4CzEFTu2bNXCqj1bwXNp
6aDHnupebV9tyq4XuLyBQ5mwcDBlotoXgeQRW7riNUI4hZNaIdZKWDhbMzjvQCIT
4wFkW8XoaxZxLpNMmRz7Cowh129s5dwjBQ1MVeVKPW2jsGCKJvlT9VBs76dmT4zc
5dGg/hdaXTK3Y4QDuB1pdKqkdQYuspvoyupfy63ICq6PO72Ud3smQu9Q3PCqU9p2
K3R9VwRZZ1cJD3rrLl9Dyc7XI2edMXsNTA4siGYbOVcjGok45jeKFYUNWNZskKLn
rPqE0VgyA/ZNugusbEnmeGvR+6gjZueo3i0hMIlY+M8rf3n+vXgW9P/5UovcRTP9
38H30UYDBffbOyoqry0eO5Mbv7RbuvAaFjd0g3kYOK71S0JuThTlM6yXmDWQ7jL9
uswgH4OOsiZ25QMzKaonqQ/3Mym551Au+eN/n7fqfRoae7e3XYP48YyUzlOKk7T9
m+6T9lX2yWjJ/h8s95V3o9B+EmW220nDvD0cOZKHWPa9wqLkXnyv8zAKIhxr905+
0N0wEXonWFp07SmpgHc5uLEYo9f+7pGx9o98gLd0PZVuPkiJun2nLEl8LIsec4fT
Ctv9f3cVTcBNcBb9y4OIyUvLptbxksg/A37DjUi6Z7hwmv7wB3vUkJZFzPN65TWr
+UOJqoi5jLg8ll3LPXfPSPxGJ+MY4M2BQ323fr7YIrp1UU1lW4JNw2+iEgp4jiRo
pi6b/MzhBKFfumB3fJ/Z+FeX/Cmxe8SW2zaGNTbHMFD6xpfcYKrPphDwyGE7V6cb
y8X7TDPVi9fooCBkb+p69n8EBhUnMhz7vnLMD8nOucWtKML9bHgPel+F/ANhnRLa
NfTr9ImjMydTLpVECtRQGNQ6lbsbsCUAv+ndpq1rpZ5oGqNBICznXpiwe7z0PQhX
he3lzbac/XWLdwY9YR8qu+9hEggJlH5BoRc199dyyAsxWKJnrX2B8HxLUtJurIhn
IPbW64wpUwUzd2nBzonqHo5QWrh3u2j9HdlL5O11G8aKY9nelHFLlKyHiWVI3DRA
aiJKB0rx0YdSqubti8bOLLhKi2SYddR0fVBAEh6zIz5kY+n2sG2jZlT0LiS/HiPr
AkUsvmzj0RkoBFxOwJRDWlV0yQAgJhTF2c/loPiGH4iM3/aTr0ilhyUzSWrVCEmG
m9KPtfez3HVd0pGSQcDZF0HC8eTaGRbHbl+V4hGFK4rr8fBsIl3FgjFGAMiPU/J2
1AxUFU9BE9KlJHR6UTKIFvxOnLhoVsI9OGWQkp8y9cKEudYRL/rxghh7rDX6qL6d
VW6bznA1LK1Xvgral5GXW4KlsEaKAWpo1jEO0e8TJu1w3kGsK3vivvc3rCbpT2pj
a/qd8POqyOkx2dTLLCnboKm7rrESPyvxfq7HlINzuU2oK/IniMweectDuMLvYdbK
CRpc5ValgRSdtTeTEKZSI866740IX8UBdyVRJSbSAr0roAabVXNUuMiqScOQ4dWv
C+tUtQ4DyAlWentJFQd/RvTD6C0MT2kwOx6PA8bmWhtisdfWZDR8j13ktXPIsIkv
+CNMqwfgdwFggpnLxRrmIJ3lhlJmlg9K0Vg2JXDzBrAy4ok6gLPMRZmL7ZjlzDQZ
E7liD2yB+9rBNoKH/npq+VB2C+wmUclfyR2R9Iks3KtOuzFdURIfh2crABWFRqXe
POtMhWrAa0zHtJsRLNf9vpyjykTrArD+DjeGawUqy0DJOhY4smSma1XDA7Gp4D5R
xwMj0kRPOy8HrC6DRxwXVkV5FE85TtWfm5I8tsRBO2mhO+tF3VNy2z0Wgf3qF+rY
3If3F8T79Kw18FffE54vHaOTc2OIf+tTEIeoopPDgavsOR4sVLMAd88MfO2pUXn6
N/5rFAvm4c6dJDjaP/qA6y4vTPCHKMEaGRU/CB14PBCB4eqMfTOjdGZSepamo7Sc
swBpA7HLnkx8DGC5nZS/VUnswHq5v4XXkqj+QQuiwvgagy7p9EBjXpUgDC/orzTL
lzdL8wuntMitK7nvRRwtGiL/VYoAFnvp4ssfs1rK/U953ZSTgEOyEdbBYymuVbLP
ffSOrBKX9A6b/t8HJhuDnbHQvip4CW0+9CAuxhkWHxtRGvilTligiFEVgU1ghKDj
BAzTdrpP9V+0ioOFBJ84gyBiy+bQS6tbGZhJ0XnFK9gplfnwePZDD4KYYC+i0LFp
Pgk4LhMcw/utH4MVcpy/VxnU/LSKijOv1SJTQnyXlwjcnmzbaZTiinnJZC7Z2iyK
p5PLF4Tv0q755bMsI/FLvCIohtKY6QVd0ur8DbBDO5gxYT5XvR5F3cRvAKhB60Je
v8cgO52m5r7sorHbeomKmfFMr2MiciXkfaPFQXDZIjB46G6D2YET3HaWnmxKQPrn
dpwzjNa3L18JlVp0a3M6nmhAuD+FWzcN5uWU3ukiQLH1Ph2K37yecerMkrhVV5Ie
RJiWIQSfnuTSn46sYavoieRWys+ihoFBqSqJCKA7qFA+qNI5lfLOINbveLLDaVVw
6V1Cv+Ch83YrQFB1uZrv/8QRFD97AR70TLviZlg+q0RE5kQoL+b7G0v2IDTYNDA6
1mpxrwBk28OPcZuMgrrC6FYp32+FsTU/7AIak1O9gBz8CCTwVy5kTFM/MMdr1Ag8
h4Wys1cB7FK8yS1qzQTcolu+zHjWpNqdv+Cn2MPuRWZH7pdRVZBsAWv0+rE+hAeW
tRYJMRoily4BHmj6Fl7p3a7o/dKd9iH2ICN2iT79GhStxiZsHCM1ty0kJGo/4cOy
xYt2m2uYJz5egmEOMwychW09sQZzsLrsVc/LfPk+6J8uPVkqSOSZVsIIg0s+BtDw
QKGKjtJ7kUWc0inye74efUqTCFURCRoA0DK3Kv1Kvz7pSf+3jYzOyBURvv3X+Q9Z
PNBE9VkR1g09r92w1YTzdhW4F/V7CLnjt3bMFW4DdeM0Dy4AD7WM1mB2aceMV/no
76HEO3ohSyEMk3YMN/W9WUaXM13y/xBqHv4/zLqJDk6J3m7UMcez9tlKqX3U8RCP
UyyIgiyMn+koFVmue3Vv9fWhBvX30aRQR7iAhjGVXMhCES/Nr5vysMDBnkH2ysOC
RvTqcQ9OXxfwAyN2BPdG7PhyIr2Lu7cCPQO2UTFwyK14IBGCXPAvY4/oIOQXSDDs
MvTG2ky7AFYnj3At6oyP6JBVSqWDZKR1KdXN+Iu4t8vlNd8kBrrwMTGSa6MoB879
bSIKYN4m/dSq7zcmZWk32GxB52sRCTUCOa0ZGLtgs6oI9pgSFSyv5vJZcilqsl/c
KwAfEx9zbTsCjxKaaJrpQdwrkg9NcfFsy7Qs4IjyLbVkokhBywfbAR3oWJNKQOrP
d8usPXDl333A6oTKWrYDJo8IIcdnpJP5nB5MkAbhKJe/Xb6IlXA/S4NJxknvhcSf
/BCDf7aHTAcrDGJBy9Rbu7+W73qa1QA7K9OvJ5bgufcVUCzRa2ouI4JNg5eWuKin
bQ87w2b53BnjcBGOeN59j2ZTgb1tHdk9DZRYXoh3SIiJNZWr8yTsKZd+Ttl+/cOa
R2k4utqt5M5U+pX1quJNRStjT6Kf1VVKIF/Jua3SswUhZDTmiMRobwlOR988uecU
SMHckF1ZQ970jkOepi1T2MEEH2N5EUEBsiMUJe8roYGiKRkWnq9ObLWiklsS1pse
3AUKKLiMcy6ctWai8+IbXXwGGBSMP3YQDovs5yTXMKIW0TGjEcXi3X3UR8fhVzyB
49LIYUuUSxzl2ECQYIRq6i/oM/chhA65cxZhAapC4KLELk90yXy2E/vQ6DDKW7rN
T1RDVvVR8rHZlYRhfDv4RWs5ai6ceH64qUIGSSftqH3+Ng+mskbj4DSXZddFNcrD
6nkMvwjsZdHctuOvljQ4MtfmD0qOLyjWOMh8ggyAejcoSSqRLcLfZZD8oLpqcR01
JSepdsS6T+nDLUvREvcn1n5EicdEnsAtaD6dhOSAvn+gt0LqCP90oCsUgBewWPz0
1ijvtoL9coQ9mG5SvHjn9DJtdSfNJWfGeQUXxjz3939wtYBq1tvApqw2D7pZSaqU
bLH3CDKXSY8cMSxko1H7gasbzn7W+ogb546My4wKXSS4R3ky0aBkTaCia2hW5lbk
ofycm2WHJKt+oNGVJqeJT0RT2ahyOKbNipT/mkkmQPRHYEIwNTe/oB4NmfwP3SJx
0izfBVS1wLPyv6o+9ve8YB1bVUdAvNOwrrwEtquBXfV/1dGqhqBOUF3A8kLPw5BA
j8bjUVv7qXibEEbLbQW2BnfUaCR3c/KZ50R/ZqOBwg2FraPJkV+WRYuM6rugHOMC
QsNLsmtOgW8VbeyBVpylCIZMZzmG3W1GfRQxXBqo1UdY/lMcR/Cnpmvw7tIdmtSR
ZvoyvAV1N9zhqrN8GwvtMYF61O2MKwZxDdMpZzOZ9aG3nU1yBMnwV1ur0TksGOux
f2re3/WLeUPrO9qu3VWTi52xJXTrjLAaBQ00minmEE496EzcQFn7iPUl9X6t8WQY
0p2gFz2v+H+ZvC4GBdVVznOpkOuCb1+jO6kRGJ4ATjC8j/3YIsTNu2PtlnbOdyVc
aT3Xjs+z09dk1J7avuk7nrKo4+rjHrOKQQqvYuEPV8hUVncMOD21vufQP/yuOezn
w9EBLmSL7HPEyGzCShj0tRmr4OPramjLr8dqnJV/NceUfuE1D+B/4yPzmxW34+kT
Uve4943JNpPbJzcWhcx4lmHM/WY4Br/F5HVVs8PILZTKgDCgX6KCCOf8azLUpFD8
PZSeK4L7fKXXdq+Tp6ZRIhTlEWviUwmFXuXH0fgBdCZkJhFvLJdQhx7X4PK6xMS6
PC1KQodYa506WTkUsO/f25Qoj8mGdan7+I5fZ6jx9q1/MHUTR11PZKUf0Wiz2q3k
ILw8n4mbLHvg88m5fkjpVIQ2pN5yVzsvaERQh20eyI5u52zR9hZUK34F2lY62uPn
LS8QdbSxNc8/WZfA0Lxp1DGWPKPv882mGbhDurg/7lV+fJVv3Nbi9/XPfoQoU5T+
s0Zw2bvTLtDkWwXozKozOsgDm21DCJOLVcX8J56KCINuHgFyXbw7yX8cHd743pvF
qLT1IyVTm8ur4ID8Y0smNVFKN4aLZSJjMnaLveQC4zoi94SAjovCB6FgUx1kyVKw
Od/TU6cQ4I9MKKpqDIkdTy3hfQyKdqu1Q5R4lyua8d4xZObJX0meJtvQqjdOt+mN
NOhZOusrj8fh+r1CWPhv/DN7Su6VY7cVFhRMXLUKMF2OaEl92sFWy96xsld2dNeU
QWSfmOANaxo1/NmKrwP5NFsdaOOeBPfBrb/T2T5WfIqn5uSt3Scy3soUT2fgddd0
DHLsW1HnLcF0Hj6N2QDpNxc0FfhqEq+TdRPZUB1DiKhiS4M2m+XPfEe4oJxPhBlF
v8ASsNGtOTDh8NeKt/7AoK+9hgRT4m2K8vYB2YYI42k8q2mK4NwV2GsFNHnwFDdz
al8JqrIthEVFmF9g/5HQsBFOi4h4tQJL8vnn4mnomCe9DYMevnLhZClsqGNMR4ZR
ulGYoBfSW4byFJArZxv9zFXOjfBTP1IXSO/+uQLsdO8rj2o8hbfB6HPXxXA6zm/N
DEN+0gPEnk6pa/Jxe69E5bbB03eez0VfMR7o4BArQxwqOVaCDtpEym4btfGMUKJx
J4BSZmX6OJFEsCAFmM9IQE8Ronq6F2o4neHZSzgg5BcfjMGb0QANC/D7g/bvMZAU
v/Thoq7uZUlLaSiYwE3BHRAGm3y3+4ErAguxGrRPH2sqkVLSgjaQoxthl21Ta1Jo
/wWS9xT+HyUFS3rBPErNrPtG9dTLBSXF26dAaMYn+NQie9uTTPi65BOQOKG5HOhl
6b0yIOHHwn3is9aks3BP+XVZooE7SIUsSi/t/RgPEUpqDPUEdarSK7bMmF6emVsO
XuvckNLcWoN7kcp14sRWGi+aT9Kc+LMh66AlMPBEcwCo9KThLbV1yuFuR+uU+MO+
mVIerFbT39QqWLiHt+38qSwxTFd11EIY8V14PcW1f+XrnBWmy22gOS3x/MLEj8M9
FC3OmpTOU1/ra6MxM3gsbkeeRNVegCV/vMSfgtkk/s9oOptCQ5dUjmoB7s9ISTvp
S0OKqO+ypkKZ0NNq7g4uUQutOVKRKMLJtNbUoUx+NeX46yRUwI+DxT7m55RyIuTw
A9+N3BtzcziS9tqjJ/kBgHh3OBso+RxxgdwBfquomcMHevrsbAildReDKhgpl1Kc
8sxNubxjxKQyr6+HiVqMH2YGNlvx/d7KCYEiZI2Aov79lFqYdJTXgwtKsU1Xv6JJ
bdO52TBETCA4SjZ64jh5tINFMpMnpbMp19lbNn4mMwrVKo9S2m/H+9yK5i/szDY7
+v7a4I6JK0VDfquJGn0e4UK9CPVlDo05pBwLOPU7LFybmxidLp2D8k6TiFnI4V8s
zGtJjnSe+YfxoJYysnGVKRwzYswFDr5Eqh71hhUhjtGSGlf0oGOxYxWnNq0++eRY
rZmIlhcU1gttVKiIAvCEiUhRK+Tq3EXQpaxo530tMuaQLRoO5l8aUUQ5Zr2yOKOq
qszhxrnQhbHEtlkKALPYkuqWnSYjxZZmwJhlDpiOTHV/z2Wx9p/iNt4f+IHbDXV/
k/G4x46HYeuHMph0bVWJhIhb2ywCIKeCjPpgxTYe1PtxZBnjQF5MRPd3Wrgehn99
32rOxs6NMRQ4HyrBly3lameNxoK6dFqpEO65jxmKVw1LZzd3knzXvdgeWN1X1Pvx
mBFjoUZZ5gUlTJqgOQbGSqYAz9Kl7qx3GoTn3NOeppr//ZXJ6qOAprrXTuFwSZeW
pXuCYoI9pC1whE9Iz+lDgz76ahoKnAoBt/Qq7/Rb8HjSVpdxtH4HdVho/F0Ou9r3
4bsSQkNK038+pfHTXKhkxueb0/JAzQj+xl4bjkXaTQIGl2wXTdW3huiFKlfaUZNW
UhMUJjVkAanqNsD+YtTxk6a0HSaxwEPDdmKmpRaplyVEFspoD9JTgYMMYF6iKT/n
RJ0VG/01PR7fDGklEWB/mCV0Av/lDqyVsdR/SRXBzF8gIAlxp6/nbIiCimEIJfKZ
N5XTymL6HyHv6vo6e/P+bHuSldBN6WFOHFLoNKJpCY/Vdk7WCLsqIHBxM9Ftaupl
TVF9SBBXMsbYmPTFvqJzAzehiia0qHjafYs0AsCzdsldp3xid6qtnXqpzSgwqU51
9yiwDNBPKx/g/jU41TUoMCYhWprXTJvDFfCocNFn4b0FJM6dy1Rtog1X77B0K/N8
ALcuq1IC8z2Qx894h2YmgTQqWD5WmYuVS/k13csvqTC47aumh9k4KvazuFsraMZL
tbgwLgiI6QCEOrKryZEsUUkGdNogSWr+4rxtaJJIUXF0NOZ9VSLUSXvZjo0WlO/8
m74k9ZvrCf6M4wZLs4dl6ivnC1QXxemA+OxdVeufDgCStI6PG2E0nbDSweHVC0CC
SddpVJnpdcFbBSAFdUz6ubDeh2i/Vu440II/qC48FMGIToEDdCFdkX5b+NqMQkrA
TDmOSG6fjhzNEGmMr/hAKb7FD2X3hJnjIU4EPIwA5Yqo9LOqu4wK6GMQo9bXS3aF
nhpaNknbwo/3BsByxU49cS55rOye7uZw1+XKCQfsn20PWo3QuPFBAR50JNjw0FG8
i7qYLVqwA7oYrkbAor7F6nmXSvIitfY2rjUwJbJFq9w9cGx2XQlyoLpricNNlu/6
OnSUvtcE/yxopxKZR5rCX0Mh+10ZnDJBXIofvzVITE41S8Zre6rPl8O3ys82BPPi
n3QB9wE6vtstsuLOrD1Nxl/bzo+PFVm5kFEqtTcd+yHx3/Wi4HwoTIDp4k0jIOIz
5vTpaR6uS0uqKDYgGK3Ahp14ikb8grYrCkGw1szD1dbC2H2S6jEeWQg5B6SIWZrI
KUmkw2cBAcbep00Hh1dZwJltHqlXsBBKoAUzYhSdiHjOhHpPanKk6QpU0tP8B6dZ
r7KT2cUDy/kvaBb0qtl+iqur5NBAU1eCCW7wx/KzfvZNerBvqkJrZFIt2GvLqncu
g7QQYQCSN6g5KRIsvmL0B2PnYOugXW1aDofx1ONnrGEQr1v5xoGZzznwdMOm8RJ6
0U6KsQ3AtfVpysyHjDYTeycH/4BeY1rzRpg75WfZoZSpUs4SgZzv0DkEabzF38xK
Llg4fJlcIGS74EAGVQOyMcImfoWq2ar6+Vo+H4BjJo5R9oXTM4L1q7tuU2KuAHsx
oq78wZs+2dEBd1IdDR92ctlSW2woi88pu5KK1ICmZeglGt+B44/kIfR5rmLaZtRs
nkQbpsx8PORp/4jUFjsDiq2dXyRozhPDeCSJntTukJ0vb65Gpnyk3981Cr01TVku
SnYSM0j2jirNRBnqsYdiGqDaE1yvlLYuz0PDyrFe5U0nnnVZ4ZLqgsgt7QOtKlS3
L0UTRHxISzfy8Qo1ckDUFdFUb5r/edKU+W/DbnGna/C9vDvLGa9x0uzhHDp1y66n
zAaSEI99GVQV2m0sunRZMx+kGdYfW0NoreJNrJsL78u1PEKXA4lLTNuZ75Y08s8H
VdFIRIGNkK3eKMGhaOJTUKIVwcMVkpnsZdxg+B8k/6qP9eaoVCM6uhxTz+MbkYDl
Iq7quKGom3WDeZ85x9q8pJE4go4a7JW3XOp4mp3nMT8+jDtptiNwXpzq6SXk0X8E
mpx/+ZIolz9k/R8BNB8Gg99swKVMScu2WyRmN63BXzilRsUIF1UL7a1YzCdnx795
TxcSZuantI9o/dBxD3AP/PMoYcl9SVRBp9//A4NEofCeYTQawU4/C9QPTDmj6qzp
A1q0eawpAAtTeeneFBD9dL1SzkSQeCc6Cbv125XaX+3nEbzCyGSl6uQR2dPQPzTI
ciF3fBu7fVCjQhbQxeEZe6ZkAxvol2kLGVsUg8d92cXhDTzfVCgqK6ulZ6LVQVS9
CVESppL7uO/5JmeIByjnhrST+tTNtiUQp8GDrJbNJIxocR+0YVMR452pqdOUiwmu
ItLPkBIbp17CCkwMWjSxR/M6AE601+rEAprN2zpqQqSCYaZ4qgDCcXCOzPOCEQAK
lODiK3eg5zugpClZmCWxnmAbZXdTfGfVH3ZlXFNFvxAT5I31kf2WpAbIpx6mUai8
D0ayH06haFEHiHDAzQagtysu0Yr/URzlbrEuUxUPjQNQ1dYqqXQfaYGJd+NeDz0b
S0SVNWahGE5L6A5DNG9wgSjHOHKjgHkXBeAKbVZWlsrS6kRRApKDaPlK23BQEbbK
hEzXOxEn8qMWZsEMgk8HZZId4V0wXoi6ILJ7OHXMs4q+H7JYGCRqkmpzSNk1t04L
Ul/2E/5H0o0Ghrh5YZ772Jn0AYq7IDJB3JZ6fe9J1fWjBwLhpgEAzUA0XQyOuC3a
OLBWNHApdQBTbeKXpmc/0XeSdgzQDwVIWS4aDgzLakz6w6R1yYpcRZCjBKx9lbM7
yej2YW8PdBuTkdvCJu/pREMIY7U4l3cFfeWRPbQOgHIBR7VkufXj32W5UbdQX5YY
fA33QhReLlbrDqxX1wqiTr0zQIKIWI3gkrwvr1/5zpQ9fBb7/h2gNmxYdHFdImgA
rIUvJhvMp7zf9VkZ4eoqYvBjRwYvcSNszgffW6wHKDBGpBouxGYhCvG+pEJ/gJZK
zRTHJE/Qpfn6tQZ/2+Qn1bdb4ft0lUn4YqIqEWwn05tCeV5TNcBb6fd08faaMJQA
qZGlYMzYhnYbNdlnxTCgfIjFy1NxYV5tZ8fMZMYvbsS0bsv3G1cNF3Ef6Mo77Hra
W1ChBkIx6ip/L+s6B19hsMdciAogGMdlbqzgVqHIcrR/DnLGmxdqGNN+wRdXt52j
8F/Z0kPh9u0jpwKp8D5MAN56QG4Qjt1psC+UeF0bxMfgLxM+TfSyQYzTXwNKQDYU
Pn5DzRxPq5y+tLcqTaBdn1G8X7M6p0nw5439Wx6TJ0LVVkzN0EHQ82ykX3i+QqRD
WXh2hkrRHQoMc2irUNGCY3ELEH3gmCb1MM7ON/+N7/ggUZ1e9LR3gtwMxOUN92U/
bRAsvDYqtRbGWvYQURcCmyj8OpQIulH97Dy+Y/ATW7euHy0ISMEwr5TJPkyLUbgq
s/R1tzXBEYMXGDX5aQWW3voLhkL2/SgIquZ/XSn3ob8ePddN2ZGW9Xc9FtbFiX3b
BdjvBXDLSCE9XHq/qyqjJXV13gryosOg7w1qqDaPFBg+HLySMyzBBnlBjk+kdnTK
DX5aq+pNUGcJtZWkYT/RaU+0EC8R35Zuq2UFexlQm1bDECmjrTlAPVGhji5thh+4
qgYLbVw1JcP1SYSFxrE9l4H2b8kTLJVN2fpr/ipa1+yyIwybE92TzOgJJZo7DG/B
uxSFidJZSk1dGA4M331CVHlW+fUuidclyHBtSrJ6gdS5qAWDQHit5Ze+Y/TEk6Pr
n5qNP8Y4/J9tl75fqm6HVhDwfw2Td+LdT5G3zQGsvLH3675HJR8tpvBu8aXQ0vld
ko/BuBxhcw52VLzLNg25VYEvzKrje7FQzU5RJ2aX4e0TC3oX50vtN4k/h8lEIseo
UzhRM6sHDpOBSlwke47QPTjrSgjC6zXmn7jnlJoqmqcmcK6BBqS2Pi0bfKryE+WA
zCI7xM42fioxupDXZMq7Mgne++PKDHwFn5LOOYwqxnBIx3BUiu+LzCGJSM8IAZhi
iZUNimCTCl103P6Hjd6K7r4cDJAa0ceK9wNuyaBmofn9pMExJyuFjJEJitA1mVEF
zfsiHHRmh3DXIas5seX6YGP/RgKTCDgcapZpnJtRRAPt9Vso7dX78OK7xPJho8aT
ZcgqhAIEDdCfCnKJVqKwyKqJg5+zpft2OeJc6vpiaKi2Ge4P7ThnFQAqfZ9+sq/a
LIgbZnZJy29kxH2KV7y7wCvDn/R3yYYgOgRkWb938pTTkD8tibDr/0UKcYefWYTS
zLc+Q1DdxKkk9mxH9yA8e8CMeVeOxzPa3/6GdocrSc1qCds8Vi5sDL0oUQPXCkf/
zYTaarVBA666TYhSrp4B9OWZRqrJJDPPHs4mwmPSmt0TmDgkIvzPRc0Rq2zNFzF6
Cp+ZMFgKUB4Y7nAnlVYTP1IMNriniXKIEJeo3DCYNk3Ku3p7u8L/PXMCZywFKkrS
n9BC8orSzmKJYcPMKVTLxYAGxSvrxR3VH1VgLyj7sCenBBlQpbRR/RbUMG+32wjM
eEZG3fo9u04gLqdmh7exutrztGNEdoaavTtphGS9ZFplr9Q3FvIHwFLQ4Fx/z6GV
7FtbYD1D0Uw4UQ8lv/40IuN6R4x3ZFLRHgZzceYB3fCMnWr69eNrttD/tHnujxrR
kjSw4w03Xsyo6t9lo8erqYbdgOl/Q7t84OOHcHorBv5Mr6prkX/ZsHhyVKr7ofM5
HrSGrqAF4kPrhtWHn1VX94WjBS2xru/RmPfED71uipVnYim0kB1v4QoPMyxkau9p
pRQTBshJ4Ou3b6XO5o64TScUWyNf6vq6fI2Kf8BiZuRCslkTDJZViTDpZqqMELSz
sk+3Hgf2KqpHrHv1j4aGqv14RTsFs1uBeGuNwNDXG0xr4uJScefpsDRi+XRQ/S28
vIMGRqLpsfshILL9kFMixWmvHwW62rHlGC/Qt6l6DdiVw9zrSxCT92sHeysc6gwX
sWwctcqAMGuPxMLZNVZP5p1p3AeZE65N4bLs5dT4SwBuLV4SXw7QHYG5w7pihsiQ
Tmvhg2jPfvMODJJ4aIzBf/sams0fIFsIcK9DoVoxnkIVn+AJ1VMJQqLcxSFcdlN8
b9cSZhACIEtGg8tr8Wf6etoPC/GV/0pGdLBd03skc/zizk/r9Es5vTBy1kuZKN49
asA7C42iaSG9qtuS9ZxmwdPY9I3Xc5d6aPSEtPkaxoPzuCv1/PA4ETXXXPOhY/dY
E7N7J8lHUkgarUrzwsSTYFsnxBjbkhG0ErgtVWhuKJxg2YUsLdDpmEh8eG9KATOS
/Ah1WzWEy+UkHDIeeClJGtOE8TYLacWbLnGHxYHKdrPSzggAOvz5BPsLeNc3sOKa
KokHlCY3V+TpCnzmhqbaLfW9Var7Z2hYueME8+ueglSUPdltbJ5UjynTnlX7XIDq
RQSf/GPuHLLbLU4vfSg56s7WYYdEsf1UsxkulafurWR5WGNHVjiaA7PsJOF1YQsF
SxJAyHv+nB6kyeepGsxYfmWRngmspqQj0OK/EG3FIB0MG/55nzZaS/FMXtQTOuv9
ONn5NME7JL9C1w+R6uQl8is4ZfOo4ybmavDOaO+jriSvsvn3psHx6QSOUAmnYZNQ
3d78TkrXeH32rJF8wPoEynGgyJhJFQ5ECoeXHRd5WnsnigsdPVrzgNA0Z2Sr6WDG
evcNFah0tcEhbMHrP6ivlnn1Mz0jUjTVHt41gl4JCgbhrLwpWqSm01ekDf68Im4+
crKrKggpXvSY+GzGogGd91gONva3mZ5xMqikhTR27TtmYjIcoBqPap4MCz6x3fxn
/CZhZOXo07NL8cp9Vszlj4Pg4yb+uXp3OUZT0bScY/JXEbijfP1+xhRBl4SLeP6Q
WY8ce2P+nUNbegcy6/eH9X1WsL2RG+uM7H4Pc6JSsTdfmytC8clzZOeXeAYyf27T
LVmaeFA/JYWHeDE9jVsqvOGmrAZ3kOn3UDtbJtxlwa32ovJxGJUM4TvipuNitQ8w
tONsryHYGyboebODhlkGNb8+XFxqFYQPSOOd2PMwoZnJAb4piF4djZN7wxjVY1Ek
/zlv/+VcmHniXYLictuGzm5XCuYacTp5Pl93OE6J1SFUpyF7jWEXDyeylacLhEPO
Dl8JW92YOlBvmt+iF9JKnrAPkk5b0Qo6d0gh+1hPqoDRPx4Wo9kU9ntBf9Bj7tz7
qFAcJy4Fek3tv4igHX3kF5Pdsf8rtUBcuU7vKx3Jf7sJVX0OpZ8k2mrlzCayM1re
kuiSsXJtXqb3WwmreAqPwjAyHYdiQsdcni4zX7+lAR3iBpffDyXD3Yo4oEgGnGF4
5i1+ug8gyRuLPXnrwT8BS9Sj9PlfCsaWvuBSGqYuWt2quVwNLrfhe0ASltYXyYsh
o5h+44sTopTmA6ADUC9evZA5lfJRTpxABbehIfqCO5zrqiIQrDTy6DLDJq2RhDnh
9uuJp0UcxwzvyXpGJddGVxSynK/LDjQJLe7U/hMC6s9owCeJkt3gYc0ZH2siCGcm
AFpvGBpKY/YbubzZMOG53PujyQEt0/lGXc53fOQZyV1DIkaI/v/r4T0c1kFzsXf2
qP3zSPhX0aFGgfHXUX2OSX8Ukz+jyxagn7UX//vHwa3B/lALWAvkc2Z9FCzzJVVK
/5V2pQWLRq3S5VLXGTXz/V3slQziFoU+2kKhlz97T+dUzG7FPZWXprdys2Dt+rVn
6/G/XCd9MMHLji7/Ulkb5nwQ21kDRcwDI0tlObZzEFJtVVEG6/vi0tJXFRP2IsDX
3nPat+LbKZJ9JrjRE7K/GjOWpd3mgGBXNx5Unpqd8/LFxti+nIRY8AmctPSkcfnW
kpUeQX63vCVqqFKqboKV+bCN68wX27l6kKU6JZZYUhQj3XOyvfKGUAvy715crOcw
X2Jl6siOYiFgj9x07jSNESeZSaJvJh8PHvaYUetFNZlaSSngBUkOemreI8DwHYhP
S/1Y/GKqrsZdPzVnMn6gHdYnh1RQQL2O/wP77KfcZ5XL50Aa2RPtSYycrfcpu/pZ
DYyX9KNDvxA/3cf2q3Y/gInB/966c3+PLSzQkJl+7lPf/jRbUTkM2w1EBDjYFt6e
wwMl/xFVM9nykxW5uQbpKlMgfVtG2o5Rdpux+JPYP959+ASsPPaL9eUsg5TqEwnz
Zmtnrt2SZ1KLTYkwPAsb7XR9B1a7XAAw7waAan/Kxh8NlW7/wEgEjKOnIttlBurY
RQuF7So4TFQwBjzABmuessJsLcroKJnwPB+cWovz5htXVOlai2oH5IUe0s8cs1Ky
9PgtJr30uRndBTNor8fIme2DqF91lHILHz00HTTWQvTZPwn8KqQ0KMV7/XPgDByi
/EOTSRZO6pim2FDV6NoD9U2R/TkMb25A3/63QwwoWQEUf3p1ay2XGehJ4eDneb1w
RAj9lbw4FATYQXjVdr9MuD7Th434/z0kXN0suw4hAhPoxIFIN52exVkSSk3YlHRg
OyawaLvqkTySWyAjI/8veJn68sIqW8Dhw0c6amer8GDJrSCX98lJAFQ9PAhjc7K6
4rGdUcyinzi2VeJHzngdnOijBS9pF/4DHp/Cic8cuLawLCIbsyNoULB5Q1szUqNa
EzyIS538OM/cSaGbF2kgyXMZkE0i7zTA6/+34jvYV2JSiVmt/i7s2jXz+v9/9kjq
aZ/CL7GAGlA7XJq+8liZjcz5iHIAoIDYuaIVLN/Xq5+Q7I3fs2H4EOU0tEvkSf0C
6ZXbhL3g9W/brJP61NOXwGSUAn1C3ndSWgLN0+0qlKx3Xxvin2qKwGfnHBaILK6w
65JdR8yqbuSob9908DkvikkHG52ZPvJFfOb/fYXgDZo7YRSmenZfUGOlxRL4EVVz
qDp0fuc0LtaXEqmjr/v2ca6HpnzGw2Bz8GGM5b2SBj8TDBFM3aqiJrlpg/aznjYn
UVJs7OiYHduB0qdKyQSUDgO2OgMFaiYn9o3LvPOY2NBSVElg3eshmqb4IB0HUHT7
Ua2x/QJHqkCheqd4PKGwCVm4aE1/zP3lS9bBkE74L+HGRNNDCdLjTlLSiQ3nGqVD
MGr4UoIBUkv1fPoR+ljoNSoFqFmqn4AIJY33upYAbSpygHZbaXLwcuTdq4XQRxXQ
ypLMifTPf3He1+ScjPEc0EAEYBpHvVpZLFFuxcjI3eFyjqcTYk1jac5ApFfNBfPZ
6HEgs3FU2JBLuniISDhuqDXt4dvu6JBfx3dvuG0822himCXSM9nMoLPBJpw9fMKj
JnNvR6m87OogLw4NZwNqqLFTyKSascvN5v2C39wN2agLGstdghbwwmdT/Rl4YH3n
HSYDy65rPdNZ2IRGwQ9976x/u0cuthd7IzRJ7iDOqgyRlfYp79x/leIBhdgNA1Je
3UT9Dfj0bCmQNZpd1TdlpEYoBC4V66OeMyI5VQVaXCeG+W7e6XZhXbP5DTqS4vZG
bpJj6tVmSjPgnB+gbJt3hty+vyWJ7BvAQkzaRlLu/AwdJ4UX7YyqoFO8T73dnFIW
YKxqT5/arCAfmQ9E7oqbmcGzpophAc5Iw5NL2Q7Tmb8ZohMa4OP57kiWu9O2yeob
rSv+qXlMltn+4tHt2As20Ub0hMW83+JOwbT1uDcfsBWf6wgjruHAv7VjgYs1YnoM
eXtuEmGRgAaJKiyNjAPKKfjwUFlrp21PXg9hkxqt2Q1dnvylt152tMduZZnNNhMk
PJEXfmDOThGRjmbmWiL2neVDyqNy06b+xcsLZpjpM6/bMXkR4S8UKkBNuxRCRR69
h7HfNKA7Yv2X7V7lEI2FmTBtfGOEFOdP7YzICS1suH3oNVVJMwLr3WqtiydLIIR6
JxOeHx3HVGaRTOxlUiKnMLs6nRwciMWIx1nKFKsF5rz7hpTDPSG0g75dmwwLC7bn
rL02HOwvEr5omPHqxRSHKMwCJBN2ujX8ICS+ymnSkdOx9Lmb0uXKijKdaiAa+E+R
4R4bL1szpkkVeAae1WyywkEpEzvnsvDZ4Ty3Hm5OoUbwiR0ZzQcWo8RvXDH0zzzF
zTvLzv28RuDWm/oQuqPhHXJMo3owas8K03HHD7lff7Cz5WFX2BV9EGiGDKrxstbn
2Jr1CSe4yjjPJAFdtS2fA322ClDZNoTP6wyTi0DBoaISXrCQzwwAztPDBPOi5rED
bixnONMM/mKoxd5vAxeTUYy/vg+OKsbOzzRtdVm2+iRrRxiYVYmfOLxShTuTdUpe
Nkq9dBeklW4R+pBeG9AZPJhtIPMyPITBc/AazAtre9dISZE9uH3MLfISzGXbZ6Ii
Sw4/nGqvkMgyqJ7F+Qnuww4Lr+E3pgr+5qdYjey41qoO4DqK3FvDZ22Q7MnLtdZP
tXa90fPhZOmhhfFMv1+6l1ddP1c14bbkrhUm1gV+okhT1IWTcO/iNHEF5djaKmPn
WCQRntYoahOI0QXCqQEeF4l0cE8f1XWM0ntpqD+Yh76awMMZwCZXNTxBrGEPcMJI
MZoGb7fitFyMVV79L6BDY74zCDsoJXYgGiKbQ2byC22EYbffo+oQeqzQVqbyHMwp
skToAFF+f0Y8YwhD7fCJfV8EzLSPrOLXmDxI7xKTIcNVYlM/6ps3s5WaLlZ7BvwF
NHAcIq4blxHlMr7QWa9PO8qMVVQQbDP/2DYzO8bpvuGh8ZipAeRtBOZdxCjtiCj6
zcn77Efld1+zhwXmvmQu0xetRv4U7MrsHzQTOfPMN3E5uzan8j4oXthuNNezYWjL
H5oYbi1Gh73hTC5HgoTpNu+PxXUitw1LyTmjyIItvTlUuiCrELbi7LUX7IULYxyb
h24f1p2vCKgwzUOvGI4rwxPpZJcGQe5Kl0mdFWKWKCnKtf1Wa9xtpOb/ZP8Rd66a
KrRTK3pCU6aUR7+M3o13bxq4gIbcRzn17caNjPrr6krL7d/nyVAYidAxsuhb71gx
FddXOQPHMtEnx8ZCdguQ/y5NWJltQKUggxcI2vaPXuXK972kO2cUjYGPhjURIheG
DGVLeJSgpE1dn/rIidHP4A9Adv0cnF+SwPcWKbWF51BhuHQvFPIsvxxmLxf8kdRb
TpWdwGiMiB9BiFoZeYWDpehZPdqroc487P3u6kB8Tlj2Xul8RiMk155jKmSBjxxp
+7GY5Q2OQQClKwX+WSEx/wwF5jtjX9XnkyS3lLaiB6+CAahk0cO8D5TW7/dL9fjQ
+IX9W3csDu3OQLZGMfW7Zjo/bUpQh+L6f/jNAM/fwAt25HyZSnTamp3+57yq207j
j3rknJ+MpIyDAcPaG0gxVIsjdxTbQfYMNM+EtvJmLXAB+QZoOnswHK+siPceM2x5
oIqcGHvr4vdOBXxN7brTcFMU6sMOi4jbfFF/7SfZHAa2Va27TCweZzm7A7sR8DbG
0aXp9lh698UltlOIpFMfi8ywsfDzt9r1qBxEPVPd72Bu+bqRCkWddKVyMkKgblZ8
6DKiW0Z++AOA6GV7nUdIIgzSoBNMWFL94QjaXNXPFLaY5YkBUidkvZsALgfMCTox
VDJcxSvsJjjvGAAeTliTk23/74y7cgYdYDM9rnOUylIbRPJFHeCReYt8qJC96IPy
+1c1ZtRx79CbtFicAcXFLAjrJfHDzmnEL8ubHN7jgLn+CXUlbS3ap6UIfVBhDBbV
AGOOGFiA62+YIeEv0qn8eRvPereQRdcYd39rPEtuLgDXQCtYjE89xiE0f/60Wt7t
NUyMtkDnrZy+QsBYE3gn31phzT9JvQ6VA/LOhsrUPypq8gQ04xFlt8qs3GNk0hr0
13ssq1qHZlTahQ4ZC+JWcBzsAMC+6TsxAQ313gY4Q2zSVg1+XyqbMbhw2MNtp1Kh
LYwpayKNm36uUaMPSy5LVKcgVjTc66i/Hn+b9c7+HDrxZAVAZfhjIAz3yVC4QrSb
KYJWtGX+ruKOPscGFIYk6i0HuK7JEdMbUFv39LIzcGiwrt7NPpS+UeizjLqqVmWN
jMZmrxeM9IpyGOH4oLh0XIjQL4tFPCJZO54OCy4XuTaV2+peFlFEZBFlcW4os6wP
jMgwdHbGHone2GYrPzFQLRjHqdwry9Z5muVsCadlOJtEmB+OB5wIs5iNaJ0F3L8O
dMH74MmInu1zYDWFg6x+O7uHUSGm2C6aGz2VUEJnfqy1IHxhawgHVwYGt012G0Sz
kHwNHLnEEgr1RFTQDwCk2Pnl0BPL/6Av3wWPRmUwLqJM6ifX8i1TsvY0KdZfv1Fg
7iOq6uyGbh+qgxZjxbd5oVxp47N6metNm+XijSctUMEiaxCkIljutxOOHtpaK3Tc
ybG8Fyo7+cbymSSlNlofvITg/09Tw/DmWKY3BDrOj0OYHctcnAm44lU8E6dykU7J
zTAFtUeUBldN2lcI4Rgge7aWe1Z2cf3Gf3dG49a5eXzR+VdHSVb016cYD6sdyPXF
pN3cjJLt91UuGj7l9zo7wHh5GfxGl77K+Lbap2Tl3rHQTRJ/WxUpkKBmAplDMuaR
e3NnR09oAExYEOTxgcSydSIjxrcuY7xLd5euvq00jFpV0rHWtzSYaiVJg79xVgSk
tMKwty42XZVMpFqWFbW4wIWjlHnKdhOxHzUWNDOhEDkeSq5hBpqA0k9SY7Xmx/8F
LJ9gV2nK+Gxk+G8DhUIjMAJQVniQ+8lKqsD6QXFZ/ZV4N9CI60LaR+q8vopjYcHm
5Rtwaq/Z49Q1HPnKkuaUqwTfFRk9Biv1eP5v46h37G+YYGIrGFyXuOQQ1An/j5Fk
+PUi+mXcbL+q6ISi5sGS1mL6ZI1yP9txlV9fkbcHMVHoWU6tL/usOArjN29M26vC
W2xLvZ7+r0DoUXnc82O/O2jg/AJjxfifVIIONK1geiCofddMtpv45OOcY+ykbCjB
pk3jZ238nLTNGhYqOp5ROJRFcmOPGIT2YJZCPf/dVmck/e8i+aghRiHuS43E9djR
WNTcaLHQ1SDplOGgGHE8hEeKyahcyiFiZwQCJdom95KGxkpc+P8htK2pULD14zlN
qugu+JzX8fVVnAI9HGHAC3Jz7CSJkKg0/veu85uLWngNBxzovKTjKg7FiashpyWd
IoccJxSyf5xftlPPypZonls3uLIkw9tHGw1oChi0Q1LKbqxlAce+8ChbCjKPTlY7
qE469OQtOiviBuUejkh66nfEweIava15h+x7AT5NhTk0/Xhl/O7bvxBwpQUT5AL5
pNQnOxaj9mgsTOE/aZSQda8gOgF4geE2L1WB3Q3jgRueR40dEWYudxvN3lKDcrjA
2BdTM0v9zy6kZ1eZnSSA5RseRPTf8OAoo8TRdpFxRR6gZ2rVTIGHqh5Y5gPuKlQj
XAY5ZUMjBu9zvGY78OTAInEzWBBeYGookccL0jvzHx7NN+UxQF1I5KkpoRX4Vfo0
yENiLxWB8lsDhtcGE7/PDhnk9fgjn1gpMg1WzMQfvGAdb7b3i9OxiRlGdmQniw2c
PHrvhMMM2ZlWqHXBtzRVhZ8AMdp3oTeHzNg+bkLo/qXmb22GyKyVBFLOx48kdyN1
aNPvZnE4Y/DkM2EP8j4+2Fnj9B0rJZOHSZO1js5LrSkbXxbTPz7ThY2WXy5fVZxt
FLumgE+ka1qzGhOdWxV3aXJcss71k8b4oPkrt2b4kFxB8LxP6FkZvgK+mHA0UVNM
w/zOrpTOLsrxT9AeHH0pW+oCSuthud1oOHYFf77znd7ilHICfIkwjNjDOfdl8Qtr
3bbMwOvgTnUbvJqE5NGjANm24CT9uziYE0bUNt0bUt7w8vFAV4a7D3LIJOHpv2lG
fBIL4NX/KeYmAd8u9Ok+17NYYbdl/YwWJE3pghBJ26PQ7DKg+4LZcCTDWi9qFSsn
xtCAZFMkWdiDpsyV4mJpKcsx6yOeGL5Rpy7Hh6OdjUqKvLifdsuz4Sc8XnZl2Rvm
afofRiDXs/NWfGLp0D/PsskTzd1tIpQuW4ZkVHUW9OIz/VbaPKpw3q+NTgsPcSsD
Jd/W6e3p4mVGDern4YV4W6fMKJbiaiYikkTChP4WY+TubxYimMDsquI1jYjrzJHQ
UGfUEu0ct77zLZ2rNVa6+HQsVHmaA80Oc+pJItAmpXma73ZGjRgjQmXyS3tRavfZ
aWdd5aWZ2YMekNgnOPTtnammhSGEpL3QPnxRiAm1PIlTNCKZbzwNjA8OznGaZ+Ab
ZMvBKkewdIAExuOXa1Wb2hfe3ToqP8SHWjnMaU8dfcr6BByGjGvZge6xEXWwH7BC
SPWv9CA2eVCFAdbl8XnoF2Kb7j2QSqFm7gtceWTZOy++V3wEBCM90EqOmKkLfkoM
uJD5nPQJG+Ov9ajKM8BHAtCPWDk2KK3u3ahbGLn9J/R4/LJn7DnQUYi/3266Z71v
AFzeicE4O+xaPGr8l9XvXmeqU8XwflV/Rry7ewmGa46dlMDOio7jm9xKf2zIIjdm
WKSk5QNuEu2jmVZCHXugzDnfElRANyavmwqepcBbatas1mIPP8SZaElroHZpwMbS
1sr56CUyKlYywKRVkshrH4zINgh5t4upK7CK3UGJWulRFCg2NYQ9P8qpixAZpKok
BKk0Z3OWYAqzvTSqVJaf5t9P4m37E4nA8zWAqxoHIqN9Qey9f1ykxG1Ttlbh0hh8
bPCMTWGEy8+Xr4qo48eJTARMExgZujXS27d9zUU6NmZsm4rBlSkfRAe9vFN3zUI8
TMcxPJXocqzuLW9CtOYBbV1rWtsXUC5etYyYaLoa1k553exznMr+3nyrvzKFjZKe
QJi4pByX3ZgLVP7NGZ83/i/c7WKt52C+wDVwuyRcKok8BwRbMqqUx7RUbvrF81WY
MzDoig43thz+/1JAlvh1txS0wxVwxcpg6YvaRqh+Sj05vHpLardNRR3lHb1i5LL/
UtP43hOSm13rTtDCvDARg3PsXzEweWdwAWjjMg1q+hk8ZLZolrwicEUhBAUWop2K
PC4Jt6L5baZtPBCC+W80JPcf2zCSYAt5tjtkEoYi3DpkPwGPtTdTtSSu8fi7QZY3
XaatRAaqtUM5JvFmKl9cPtKhPW5uLu+eIXdH15sr/cX8HLgt0zVATjwUu/jR6cuQ
G9UwwFlilnlcEqTYoVVgilLS+6ocjX6bpV3uxGdV7ggs7jmtsQGhGsmAONynYqDp
FaF+o4+BhCLwIVMBLJW/+/pFbihIbrxrw1CRyylgnMBuWOUlpqBj6Zl29TtSsS/8
YA9thU7V2D1yP5yivFRhs0d/beH5ooyqv72UNtvyW+mIC2/o9rI4hTYpSrsNM6Rp
6qFo9zamhThsLSxCoqKGPZlYMYmAshqdEwuCWMQDcrNFXm37pg3/zROZey5jVOej
ngakTJHnH3AbHSCvsP4n6Uu+bHyENqL8cnz7gT+syIlsyBjvLwCnuyjLHGATGNul
lTeI4p7h/H8uN29H5iWFg6jmOz6efNasKKhYh8Q1DzAmFd583QWQ+SBB51HYSoBO
RjEM4Rqjke1c9XgKvV+zzltSqAW09NUWg8T+l41Ic5svk+/xw+u6+euhmKj8uvIo
lXYxHZFO+IifbKasQ8VKEXPiz/D81yAMJG2GydbvQRXUgMsXq7ULx10iXoaadEIt
s9IhcU1jrU7cTTsEhUwhqZKh7JPPnzuM+3ozaSS8Sl4RdIU/LVwZSn48B2MilwnG
xdIItYCAatOloqw3WmJ/VXpCMruO8qS6GKq28Z3uciOL0zzfUNp7WkutjAdnARLf
zo56NFlEy9gBeyRSwRas6poOCxxriE3QgP89tV6eA2QL7P86bKyeA+zIGnJLjh+r
BgvW7vMGPI5GOPvMlbqeqCW48zVhATnzbOfuJ/hNEP0tYtPcs/etyWPTbVzY2yUp
VbDgEGiSaVQ1YxME2+/gr7KgJ3getdeGEp2ozKp6pvnY7PocKjyiDL5tSEZDlyhv
DzYkFLJerllMgpBTNOvorcV5vYneq3qdRchCieC79vIkZTCU1e5fFYmJe9kBdzVX
O81FLmnYjYIcPuQEuTX10bpTJ0krfs1nqrNZyupb3JGTS6jW8NaQmYHWYQ8XdSot
Y+36FoLluhSrrWltkmrrk1GPvxCz8c6tzyokpAh2GPfhd3OEd4IvjMsTMEonbzmV
qOdtT4q9/mWLvf5DwxEvJrqB2wbA+hI3CxR54xSEojPis4gJAYpIp/n24crGpUQM
Awe32zKNl3R+5BQLWxbdXHBJXC23fOrd8Sp47zYjWZgq1hdqndxqqjoCDL3+5odh
TCH84HnW8FNR/ogA416wkrpk83geCxMz+6cjeUe/pURdmJOxUpf6NHmA3cLOghQv
ETmecW8RNhNOHwY3hg8L99uwIbsE+iSz8xcCVZmRN+9a33XBDfTB/IQGf5JPMnIg
67dQaG9bhclQksCPc0qOXuVKNem9l7+AxHXz6hwlU81FOSHWvte+bthlQVXs9Mf2
ItmvjjIK2v2Xh0LXE9imjL9MoQI0fpld/liNa7yv0RQd66uZ+Xf18+xPbg2D4vEr
4IVH1ieXgSWdFoqammuy3NOGhfqhg2bfNsgFbJZQA3/IMHYLCt8p1SyH8FLLJjWF
FcWHkS1Z04UsXJeys5pGKrDPoVz7HUPanQbpYrrxwEYopMqgcgPJJ4aAojWAcN/Z
L2W6bGCHM/IvU183CbtJIvJxHOoSib8oV5EgcHmbSNCYv68Gn7LXxGUQxX1tQgGI
sr+oyGMS7HZOdjRRUJlU3276L8WLX1XXZ6t5SLVwoEq4WoGIIVJ8p+OGMhabxRun
DwnWlIHYDdlB/sWNKQ1DyXJKrIB4RoGSOGBDWAgBA4vLZZQsIloT4D3l1XcmZ7hu
fALa4FyWykxZfJn05RqALnQsxWbGrVThOvAkdD/mtIhjCGfvymm9W2ioK/2l10v+
5/EEL7LpPg3JZRNR0F9QGfYbumYDd/+88XOew4mObNLMViAyBhV6YS0wGcnBI8SR
T2L+OyYTUpc5YYeUY5SzYMTswoXKTMKkmZsWyRWUEYEZO3HiiSY7SemLKobrqBCA
2zk2QiBtlRaOIHAeAP5oEZQ2BFiP0cnumDwHrCi9O/LGwSDQxo4B8hplsmh30XVO
JxvuKlNyFeBbSnx2IdxdihvniWYuJTNZaGYKCo++4urxDJNHoJEth0MCe9vkWwM0
qa40fOp5C7iGW1xurnevR1hmV1zwrOlQTXmduM2VVjQ4ihqSOuk7lAfPbus+pIHw
wwn3hzaZKe92rYaQyUiEB8VEImCh0moVrE5IZANeXM1bOSqYeZJUcEFhI+p0qiL9
qgo/iWXQ+oOqVqPmEYCqMNiW01NsYiZPw8ILjftAeuzNRrf2ozi5QEh02zFIMnxa
YBrJzr9YYVLUhF7a+H+qxt+k7Z75OwmqxDxbAYJbPwNVotftfbhuhh1ws3Zaj+rr
vcaxnkSZImo89z5MXpeik18DYk7mIr7IoMV+cN0ZnGYX61DSMibFj1WL8VKBC3E/
6oMsDxJ4a0bODDfWEtMLiY3+BYBckC9HOcJex+Z4IB3qepxassw93Bao+n8MNmYr
JZVTtHiYbpvt0wal5nVHkUJkwzI1yyMIZrQ0xihxq/YlAZRJknUcJzdMA0c4pRaY
dXqNEsFmguJFqpxIbBukQOo/Y6dr7GxvsF3MUhJN4S0uZdGVzWMiWkUbVQZt5okd
Kvubmr5vF2eP49YThfWOkWb3O0uQqsCrjnYMeu/3E1plp/DF6UYvOxGD6UqqWXN3
U/41+dHGVUnYG/5pu5O/1YI1KtH5XyQJM6kFtWojDm4TCKqxqiJwUYTNDrjHZw8s
OVa+Fe5daNEsF4t9F1a0JAf88dIy+tUGYNXpGoPNx0ZE0xBS/avmI4fmocKhHKGd
wwigjabNVj2/NjJQVt4UmsbjAeCQSNliHViO7paIJUDNbmLF14JUPkJB9bLT5wBb
2AtCNR242QrqT8JKJSgMI63uF4IOlEHBzCe0a3kA14J1QBUMwzk9+SiFUICcLofO
pPsk9smQ+lA0SS2N5t9qQs3pPRDQpAgQrbSY5RWs1a9ntY6dpBYRiK8UvrBR0xn3
AqvJkrMGbGTtOdqwtzJjv32Qz4F6SwWmxjF+HUNbAVskY+PG5lMapKbXC3IFmJKL
ELrhyIU3to7HFIbilRVS14hV3tbhCA4XRu8Z1cqNn35DkZ572d4phm5oWbBe2kg+
JMsOeRElhwdCMTw3u13SHJyxq0A6A5AQqK0O0bXRVdEqwPnYwk3ToeoL215jcfJt
JXNmBeM/Ya7v2j/PwMXtxvj2wHnEy8JBse6J3x8OoZHDWk7D8ygr8X1ivlvpaLmo
yeJvSpgrJ8TaqKfBdKiptY9MoHEnYBLuw1FQ6I08IxmN4TxqBL8OocU0G5XWb+u6
C3KwtbxQ37YJHH/dfxoyXRWTx9HFP6vgDPYlwOSa7J1W9n2+LNQDbiP3MguLPGp/
FB5fX2MiwYJ3BthbaYyFtTPo/1jM3fhvLz5Fa0OPpZ6UazMIuBjOx1370KA1ohkw
gI7b2SO1jtxNxPxH7VPY1U6e1xxQYfxsVag+Jm8ZmnwT7B7t8yU+5hctf/TSbBZI
64OmfppUKq4eA7EKDdQf2A/CK6/Kx8dfpz67eVI6hCVEgzClAwwPcjmzpgwFDdXx
D0vk8iCwrsnoaLOCRkLCbuWuKdgA55OwadAnPG5gwnuXGbkZr3MeCmZYSyaDyI9g
pNfTGsLS+ct2g2UIsKF3kwCwafiRq5KD7XxKdzfEaGR2mnjTaIEln8/IYvMWCbCn
eT9CajhXBfKXyZmGWpamatI4h3B7SV7vM310wzmqLt9sjjaoQWUCBR7ZWOJq7/b3
Wy83A+vwj2iZOspk9S+cK1N8a+McwXXRGsY/+wv4rJ4TMUg8tFofxHEaVflm0Njy
vFLoZyxA6GXDLcTFD6eWNs5bjIPV9NhSsHU+WAMmGlEeijWrpgtn0jhtPrdYCWTK
f9Gh4P/BspJiUyCAeKCk7DpUyuuUGPRa6TVqur85d2o7+QamTWHd16a5Tj35za1d
fRgDo8umfJP8tYET73w8xKVUt9zsyTL73p6AEuBTVgRKRiTSPLhrtRYaVu+bC81a
yE7n7q9feao0WQY/neNACmgOFHzv/WyRCqkFaPKedNO6dlfz9oVYgJY67dkwadbp
KY/cu/M5vBhd2i9CxNe3R0InVPI74bTICHXG6z1TLAf282WuLcfqNUVCzL1EAivq
TsThc37Tbc6k98vkIVRJdooM5j2MH7ITAGuTJYuYRRuH6iVVwpHorBvPLxovcs1s
F3fEZsCiXG4Tly6qGh5UheTay8ijGI8tlqenI1YNwlUPi0vb5A+wRzy1cnIjjPVE
2MONtREeAtx0FxgGvJCtFiG5I7S+f9T/DqKG/rVnwIuuhnBTzgc2eAOJTeno08M3
R5t0ssNGqmexH3scQCovVXn82E0XH5JIM9XSglbOET3AQ/uqwRXTEQn/zWZ3J0yG
CrT7TyHOsIr/4swQwB8ICqTSfX4uoYV37bjcOUqF76mc4U39teXdsiDbqfB73XKe
rVV+CJxtpU42mqriWRtzhzYZE7/D+QIosXdcFjTA/b0rmGYBn/DzOeV1nmQPDUJu
AINRBbktgLd4skL5mLziniHMraf8anLDLRi+wjg6YwWprRpdneT6f76Nwef8DwzH
WhP4T30KWQt4l/AgBebcJYY94AmGxpRyyZDFXl2AWsn51w3s9yRxpR3ZmD29CYsW
B7K3vOlU9PpCIfp72l49HeI4R6jVr/hqtj2OSq1OucxeWpyUVcw1IhgLxOsqqp7x
TmoJlNH0lB/zujn64MjFOr+3xi7+K61AV3P68IStcj8jIzjwHlcXfasSoWHrgfyf
8OFq7/dkjOd1U3+Xd+iajdzEr2geMTemuAoPVm66NJnIE0UOoBxx9bKNa9aD0R1+
/6A2oEPF2bvFM/Q2aEJx8L70mfThKRphjqiqRK29EVZoLqqjD4h1f6s8kEjI+K47
tOl+0P3ralU81V+aCdPcEHVZwiqGLt42d/YEDnQS5C62bXRWYv1QYVISB8/CJeoC
X5ySnE4yhE/B6CkKTuIMFRNeQlkIYsq3IFjgpX7oYyLiQLbF/Ad0LfaPWMsl3kYg
itndkO7sxkOhq2nHV8DeRZ42BrtNlAoBg8Av7D9OS6DCEREQMBJy1Hb+XeYyEG27
r8E1F3G8j050wDCZadjc86GHgLFwmCPxUJWZz18N20Zg0nrEi7wQBBoOBhbKf0iR
OLOrUOOvoPhec/4Poj5uN+2o004gViISv167FVROcBYSp9RPEC+6HFj/vA3+D48n
y2JYJeAGL2cwXtFh34Q1KffBK9gru6L2hOzK/My1OOExztjBRPZTCypwxvBdrod1
iYBxGfBtzR8A1EbtxPXFU5Ihq0igz9QLoq6UoGaPk8bSusvqzUeTR3ZnS5t7ZqDV
ceisJ2iN6w9wayApmImVL13I/DcpEKGcxX3xxEnAxzLm4pcdNDmW+l2G8EfAmUcG
1M9TYCg8OvNy1AAfB34rk9KpLHtLLWFIM4I5CDPgtQOh+IxIrmYkxpBVYVzS9FVH
2PMVqzYaFojX3R/8IiH2eXe5ikw0ZdsmHQcw9i3x+GGs+AY6I93VylSDo8NW094e
cwYjPoP/wbzE7mr4dLF93DfGLZ9OZyyIhI6U/ZnGz6d3KP4hWtE1UoC38PREaww7
h7ICUpT54gqI19jSU06cE8H1wzc1GRrs3OdMsrL8MfhQJkAj1WzyTHPUTOijUn9L
TPEsqnpj9+23HrHkA5fjo+lYVUaQbeyDnGgoVCobbxEidNTS3wiLagOFz/OBFSLV
h35IgTQEOD+h8CqUjMDYO2got9VI/IhpgWP7Hf1jNT01qr+38Z95Puvez7PgKLFF
PI7XTxf7sH0KLZq4Z9pp7SsiTdVcaUTQIGbLNW4d2KsIIb/5UocsYROmyjX16QKB
HBYZAp4FlxZEFgJsw78gQsyCkF8Be/uy4yWCkkxU5t/ZMiSYYWc3TbbKLfp/RdIT
myjCNuM7WDyvBNykF/gWMo9n6Ypa/OYpd/wAOB1jJcyUnBFdlmJilOKEo68AoasM
eW6eb0NbrOP7LvoGkrBthIH9NOTCKi3FmpTrjaYFL5Ka7L9vnCcC81eWSn2geyJx
zEtE/dw1uCfbo8q1RtyAptN8pWULucWiFRZwwNmJWv39ujuKxXqxaIaPRp/aWzcQ
RwfIn437zxgPR47Op0IjuVR0jprVZhcKcDQMdeN0QYHZDMmKTy5xd63T7pr7EYQV
Bkvsthv7SL+hQtVfS0AE6Y68ZVRoyf/QQKjuIimX6JZHw+NBf3ZI0W+gIokcoLYe
g+oWkvEIDr1fSTlqwIkLtwtMz6W9WBt/HkZgAAmR5+O5725whN6Z6FXGV17ruVIM
EHpsqo1W99dHSSU7hZXSCaS+oH95y1pGi3CTY1I9iS9boKzc7IFUWHLrOgqsK7BF
2vtCJPiAZC60XCUoRIencVmjWuBna5E9jiJ47mX8SC2DufeeY63FRJ2jWuzK3XEO
kH6t6H3gjj6T6U7TGaJRsF93mGieHXBdwqukm6wkMbKn6grao7lNKQGS9PSy3FQX
+5xXigEY7RsWmaGRz7Rbdtvxzhevy4uE23oTDZ48XVza3/mucSCcsRPJCmc6kBrD
KFoy/J+Oj+DRJsy5mKAwETaLxCLEGyqTR4Qild0m5PfctksBNArybHY33JfYGPOp
04Usjtskv5kM4fxC9Y6Th4g/Z3wJ5yIgRVMG9Y/P3CterhhysaUK8nM0OzlfUByc
4UyBP2G+mCZeA/5EWMRmhp9Kg8lyvAT40eV3twxYHlWaRPeeCRL8hH9WPMLA1XSH
uOzn7rOGphT9J/N5xPdAPUoJ3k5ZAWFfIlF09vGjatfIADZpm+6GKanHOF/RWw/z
kGMxsu4MOJH5Lo4QfMf/R6cj0ogVpmmVahuFl2tjKVkmQajwHdpJ+E1KEtkMDHNb
AjfNHzD/3gzMRW4JVAIKJgcZfREzLE2VzygaGlkVo5J2izkTE1A31/oOssUt3bZS
Wn+j743B/O29s/IhR6OpsIM9gL7JAb5+7wsRzZUAoKohrWDHsAMPKyvdZrS5vCuH
IrkSP7lISJ1sIgGMKlLDWpDPMDXTRU+T4m6Oj+k2G1C/HKs8yzGD1+BycWT289tG
wrwRlRduwMtRpkDXXIFAn13Y/cdDKzr6WIA39ti6OkyMsxg2KndKhUwd5RIa/qJ6
nhUpFKCs94aD5OOKol9lpp1hrUjwHnCbI/APm761A4HlwM1HLGLNORgXB4wUd0ne
LmbNxk4iHZ3/VfExXOHrUd2vkiUBClIa+yBAB1xF+3P2GC1CBANWUw5DJUR9qmay
kHETbohQ0Pws1UVa4V9am4E2KQD+8eHQCOr1wJqjhPlD32MQ6nPbsIc1oylT1Aax
xweMpEXTqAy3YsXN71Cr9NeJrbNLOA4DPRKw7e2EDLCUtqpHmKfLB9N+UMODZxOu
mzp5g51gn23Gv54kZszWXqlgjG0JSNBvPJR2M0dsUVt0uQ2nS0kGSvd/HAEUzRkH
NnkYUiQSW29Rd9aDCsQvmdxw/nbaZAYxiW/eL+3oY1qPL9m/xYk6k7vSiX1LdlZe
9oCfUGA6gONvrQ5ASulj6XNsQLNiosM9nStnlz5yjduYInuAH+Df3oHm01ngf+jS
3XxjKUr1whc+dIaUQlY/fD3XH0Wwn8yyEky0u/FIR3zcwbh9cUFI6zYWzUJ3hApQ
LJKTlwFHC/WII5f2zMZHBbTA0AbpedSjX7tnASTOJWjWDCdwwvPbYS9lM85sjtlj
qLJVtyu5fKYI2gLqsfK8NvQR9SEU9B1lUoMTd+gBD+spqy0QZhsW6j7gLsb/Y8lw
JGotHe9Q6q8ihBw5/1azvXikAuzrCDd3zDQIgzahGUG4vT/x+Xu9imckmyOmRWip
gXMzcL2ylJEJqJEh9XNmx2Cpg5DyXrN0e5f3RRZY1D+iny+Zk7haGBNQU2IfIanB
13zqkH9zgd0gjjM1eJMEiGf9f32ysaM+4cVG/0v3b8AT0jECFPWtYOb36cTEV236
nHQ1ybl19pevb/9HDqFY+XWBcJLLGnKDvM3Ux42l3KsuyErC5RtdW0gST7NslB/l
sN8Lxids590LmmFvSmzFTXAMaYtIcHKtKoZ32CYsrFLmPcMgL1MGccQXGPstG4HH
K+5M+lx07+ruIWsDDwptdEQgfPpRm4bSEoMlKQkP8KOurmneSs4UbDraxjxwg7fI
TsFYXhHz2PNE208N8mscNpSh2ut0bE2D4C0depdsls24GyiFs1eJOgsJK1dUPNl8
giQmJSYpnv342b1oB19yuamR7ELIYPTz8PBxoqvKdboLdGZInukmABLvYeIKjp6s
8Yn5/6koDuGLIB8OeZ2gOVDACi+zJmBjwk3B8kvaEoFKNE3aoge7C9Hc/yEmjb5J
kvvKEFuly3ktORp0La97Dvbb3n75U+Jm423nCUCQZdjiPbGoiskV1EcfRK/AL3OZ
RbqP8aSBP5y72t/+aaAG0T7dfOC/+hwcJPdy8DOHE/RgZySp3pgkXNpeWNrzAQm0
t8VbatSdcF1Kj3kFycbGYLG9oRkv3XZaDc3qXCICfgQh30eMzag1Y5Fv0ltky8lU
MdcPz47zAxDNVZ/wKdpnq1ZAR9b/4Akdic9VE3xXHf3zXesMcTu1lpf0Ywb685ST
ZuZxYTSeFG/KLNJnte6so53EIzGuBuKJWAxnyYG1+UELXcR+Cv8zqzYUTwQYKyX8
2nsnyKhgnau0rENfCJemd+531qYIu1YKPOnx8kZMTEQKoA4IQhFoN91u7xCQJDGz
blJgPAaF6GZMfx24gXbu2PN/ql5sxKiHWNNOtxIq1nOqSBxGxj2eiyaAraGRKKLc
8cd33m4Spb9DhQmDQl6xd1aVUcEVEtfSmZU+DotgjQmSiComYS0kEB8pSqjazPht
agHtZX4/wuVk48xPaMJFHKfFlpiX1SsHjqCAQB/yV2IQIw01QSSl1MatRxx8AGpZ
t43EBB83v2cUMtLO+nCDhYQWN97AYwn5J3qN7RiIx3jOCh+e9g0eQYxJeQb8tNuz
fq6iBGKPQiCupfd911IRv7lPDmxPNW7cQgr1dCy4EFZ83Hh6X8SRIqfm7fPuI4mW
UNT8nbKqqlYgEM5OjpCVdGqT9P3VHzg/1jezQ93dPQ+8zcAh5isZZrxRp1DnpDtr
EUXgnAMIPq1grG24wO550j6NxazKmyhCjRRcjtf59f/rnrnfG5frn9JBpTiACvy4
1T3xNTeUoXkBM3gl9Q8ZAg08Bxr+sWI7Kx++diwAW4cFgkinx5rrJ+hT/bLvrAKw
zDlCO2dWNvAx6MbMtc9tZgnYnBsRNmetyzzrTZkOx8sOpti43D/fWoAe+U49DLBk
lSNdVzQLQYLmUn05o09hNUhHSud1+lyF3zaHVEXfB4azAd8sAji73ylkARR1o9/v
fK4Emf12pgTAcPNpYWkf5KywMW3es/8fPghFFSW1/MrCdV3TXnEirCsWSdwNPUvt
kIxNZkKvDKvZeLxGF4dD2Soe1wQI8n+sc99W2/nUOX5H8BSq0ZWQWY4Ijkrkg3wn
mMEUGB/E2n3zRhA7t2nd5+OrPURBSHUGN5N2rjmCZqsWS/CJuBoQkfjRzfnmyizZ
/wp6OHdR21fM0iD1oAGUz6g/5kWkbrObANAzmbpYAS4Zvb+bQ4KJlVnF6LO/rUB6
68Cl3oxCRh63Tot7h/JPeIy3jnKDMMTTpqJQndOpwLhlKp+F/ig4qgvNx+2l3ICQ
vavlF+3ZQgBYBF9wYCf/E3XHtr6gk3caB2RVZ9YKdiCGJd0k8iS3F9Urjd0wFeap
8uzjc6nwh4+1DYfxK+aEwkIQZcwNn0+4EU2gBYoAzbmm/qHbHZ4g2tPp2H6l3hib
Q/02y1/HPRmMoSNanqtD7/mO8eQbDzw2dH7Lh/X/vLsx+g7jWWRHWamqE3Pum098
/hKIybQvZCW1S9ZAc4/s+bG7KT9dKrU5noI+be2nBvtz3ej1IoftdOLraX2nYh9S
r9Bt+kAE6x5jjZVmcgbeTNP5z5Biyk2Nfa+SaBXoBpn332FmzQ5tRfmOreRdjzhj
gWQBmhFDrg3zx+3rc59CJkQsaiKObJxlVPeM8Z9z757OX2dRwlD3l5N1EfRtPgGy
ne3r7rZGU0hPA0pDf7rxXmR1A0Eu9HFnbj+JPNs8XJY3ZWYWdrGhA1sND9o9w7At
XpPRSiGXle6ZUFX40355kuDxDm3jGNTI8wGFYIUaE46R/Ggehnp9cnqxWj4aaN/Z
pVPvL0CnnLBV9vrudLJlDLvrAaMeKexRRLtNhXs+gZ5ZlutCNZp2KgiOm0NO8iYi
EVA9Ar3x1wvkTEU/bqf7fRev1FrsIl1Uy1jR+DvAZT35N203Y7OsAbqpRQ2C8FAv
GDca+MK4DdhL4y8hJ4/2XOskk3C/3bbx1oufIU1y9BQdrPwF4nFW6nfk1ZnEj98H
reHxGzWXL+7RaxbdBkBGgv3OfpKGzS+kD/ilRjCjMRooPxzvKDye6EHhHDqEwBkF
su6VOrQfZ1EPWP+pyAUyz1MmtARzbw+jgQ5iJbuM9ThAla/ngwuLghvpyzcvRFuU
WFE17cvM8KHnDtKPOO9lsG6Y8cZhAV3seuJrINLyIpdj16BfghXH9ld7EU8an5OR
5TW7imd9whCcf92kALppsombYHMj+irgsaAlFeDzVz6TjtAZpd01+7h2695h5g1+
DABp5xOPlWZDDeW572a4k1UCkedTReyNe/poGv3vVIC4GcdvMWX1IMHrl1lciOg3
YzR0WZgkl/iNoIOT+x5qP6qybh/tSdCSb0TtEjlwKNOkPQyXqRJ4k8/BCM+bGr3u
Z17sKH3Z8HRp0yN4rQlzuS2AUAatLd26DpDIHW4xKVwlWi0c7SSHIJENJMHnfVEp
mZasxpmsP5kOB9q8DLBquSGKDvAvL6zkTAUQY0FaqYcNoBrD7S82NRC2M/bWXJhQ
TKaTUgSt7gyG9fNQ46O6/8wF63kiH2NJNO/NqWiwrj4qXb8M+dI/icSMR32YYHok
aPbwk4jSltGa8qSNXCC/a0JJzGSCMHO88PerR62QLlL0cXQN3y8Q1Ad24PkpX3CV
E78pHq+8Ls11xAj8K8WOLCItdbd5nJckrZjzjkrWJrj+rXMLoduxwD0BHaXlaT5F
/GqpBIhQkNJwWdYePmS33gwSM/ajatYldPZcly7r23GfUmGdZkthvpB9riWZf7Kg
WOMkAgd6t2BIo/atcXpY57inpf3lUsHDOq060AJQACV3WzTqjmbxI6R55Z8jhUld
O33VJ+KWvFPNZR34NpZ6gDPAjyVudfng4GTrQoEZg8noR7aV/14tfGB/cUpaJmen

//pragma protect end_data_block
//pragma protect digest_block
HzbZiq5GR8DaC4mU+F/4Ti4BFj8=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AXI_CACHE_SV
