
`ifndef GUARD_SVT_AHB_TLM_GP_SEQUENCE_COLLECTION_SV
`define GUARD_SVT_AHB_TLM_GP_SEQUENCE_COLLECTION_SV
/** 
 * This sequence generates UVM TLM Generic Payload Transactions.
 * A WRITE transaction is followed by a READ transaction to the same address. 
 * At the end of the READ transaction we check that the contents of the READ
 * transaction are same as the WRITE transaction 
 */
class svt_ahb_tlm_generic_payload_sequence extends svt_sequence#(uvm_tlm_generic_payload);
  /** Number of Transactions in a sequence. */
  rand int unsigned sequence_length = 10;

  /** Constrain the sequence length to a reasonable value */
  constraint reasonable_sequence_length {
    sequence_length == 10;
  }

  `uvm_declare_p_sequencer(svt_ahb_tlm_generic_payload_sequencer)

  `uvm_object_utils_begin(svt_ahb_tlm_generic_payload_sequence)
    `uvm_field_int(sequence_length, `SVT_XVM_ALL_ON)
  `uvm_object_utils_end

  extern function new(string name="svt_ahb_tlm_generic_payload_sequence");

  virtual task pre_body();
    raise_phase_objection();
  endtask

  virtual task body();
    bit status;
    uvm_tlm_generic_payload write_gp_item, read_gp_item;
    `svt_xvm_note("body", {"Executing ", (is_item() ? "item " : "sequence "), get_name(), " (", get_type_name(), ")"});
    /** Gets the user provided sequence_length. */
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(m_sequencer, get_type_name(), "sequence_length", sequence_length);
`else
    status = m_sequencer.get_config_int({get_type_name(), ".sequence_length"}, sequence_length);
`endif
    `svt_xvm_debug("body", $sformatf("sequence_length is 'd%0d as a result of %0s.", sequence_length, status ? "the config DB" : "randomization"));

    for (int i=0; i < sequence_length; i++) begin
       
       `svt_xvm_debug("body", $sformatf("generating tlm generic sequence 'd%0d",i));
       `ifndef SVT_UVM_1800_2_2017_OR_HIGHER
         `uvm_do_with(req,
          { 
            req.m_length             > 0;
            req.m_length             <= 1024;
            req.m_data.size()        == req.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == req.m_length;
            req.m_command            == UVM_TLM_WRITE_COMMAND;
          })
       `else 
         `uvm_do(req,,,
          { 
            req.m_length             > 0;
            req.m_length             <= 1024;
            req.m_data.size()        == req.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == req.m_length;
            req.m_command            == UVM_TLM_WRITE_COMMAND;
          })  
       `endif     
       write_gp_item = req;
       `svt_xvm_debug("body", $sformatf("waiting for response of tlm write generic sequence 'd%0d",i));
       get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm write generic sequence 'd%0d received:\n%s",i,rsp.sprint()));
       `ifndef SVT_UVM_1800_2_2017_OR_HIGHER
         `uvm_do_with(req,
          { 
            req.m_length             == write_gp_item.m_length;
            req.m_data.size()        == write_gp_item.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == 0;
            req.m_command            == UVM_TLM_READ_COMMAND;
            req.m_address            == write_gp_item.m_address;
          })
       `else 
         `uvm_do(req,,,
          { 
            req.m_length             == write_gp_item.m_length;
            req.m_data.size()        == write_gp_item.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == 0;
            req.m_command            == UVM_TLM_READ_COMMAND;
            req.m_address            == write_gp_item.m_address;
          })
       `endif
       read_gp_item = req;
       `svt_xvm_debug("body", $sformatf("waiting for response of tlm read generic sequence 'd%0d",i));
       get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm read generic sequence 'd%0d received:\n%s",i,rsp.sprint()));
       if (
            (write_gp_item.m_response_status == UVM_TLM_OK_RESPONSE) &&
            (read_gp_item.m_response_status == UVM_TLM_OK_RESPONSE) &&
            (write_gp_item.m_streaming_width == 0)
          ) begin
         foreach (write_gp_item.m_data[j]) begin
           if (write_gp_item.m_data[j] != read_gp_item.m_data[j]) begin
             `svt_xvm_error("body", $sformatf("m_data['d%0d] does not match between WRITE and READ transactions for sequence 'd%0d with address 'h%0x. write_gp_item.m_data = 'h%0x. read_gp_item.m_data = 'h%0x\n",
                            j,i,write_gp_item.m_address,write_gp_item.m_data[j],read_gp_item.m_data[j])); 
           end 
         end
       end
    end

  endtask: body

  virtual task post_body();
    drop_phase_objection();
  endtask

  virtual function bit is_applicable(svt_configuration cfg);
    return 0;
  endfunction : is_applicable
endclass: svt_ahb_tlm_generic_payload_sequence

/** @cond PRIVATE */
/** 
 * This sequence executes the UVM TLM Generic Payload Transaction in its ~m_gp~ property
 * and returns once the response has been received.
 * 
 * The GP instance is not randomized before being sent to the sequencer.
 */
class svt_ahb_directed_tlm_generic_payload_sequence extends svt_sequence#(uvm_tlm_generic_payload);

  /** The GP transaction (optionally annotated with a svt_amba_pv_extension) to execute */
  uvm_tlm_generic_payload m_gp;

  `uvm_declare_p_sequencer(svt_ahb_tlm_generic_payload_sequencer)

  `uvm_object_utils_begin(svt_ahb_directed_tlm_generic_payload_sequence)
    `uvm_field_object(m_gp, `SVT_XVM_ALL_ON)
  `uvm_object_utils_end

  extern function new(string name="svt_ahb_directed_tlm_generic_payload_sequence");

  virtual task pre_body();
    raise_phase_objection();
  endtask

  virtual task body();
    `uvm_send(m_gp);
    get_response(rsp);
  endtask: body

  virtual task post_body();
    drop_phase_objection();
  endtask

  virtual function bit is_applicable(svt_configuration cfg);
    return 0;
  endfunction : is_applicable
endclass: svt_ahb_directed_tlm_generic_payload_sequence

/** 
 * This layering sequence converts TLM GP transactions into AHB transaction(s) and sends
 * them out on the driver. The sequence gets TLM GP transactions from the
 * tlm_gp_seq_item_port on the parent sequencer.
 */
class svt_ahb_tlm_gp_to_ahb_sequence extends svt_ahb_master_transaction_base_sequence;

  local svt_ahb_master_configuration m_cfg;
  
  `uvm_object_utils_begin(svt_ahb_tlm_gp_to_ahb_sequence)
  `uvm_object_utils_end

  extern function new(string name="svt_ahb_tlm_gp_to_ahb_sequence");

  extern virtual task pre_body();
  extern virtual task body();
  extern virtual task post_body();

  extern virtual function bit is_applicable(svt_configuration cfg);

  /**
   * Translate a TLM GP into an equivalent set of AHBtransactions
   * Return FALSE if the GP cannot be mapped
   */
  extern function bit map_tlm_gp_to_ahb_transactions(uvm_tlm_generic_payload gp,
                                                     ref svt_ahb_master_transaction ahb_tr[$]);

  /**
   * Annotate the results of the AHB transactions back to the GP
   */
  extern function void annotate_ahb_transaction_responses_to_tlm_gp(ref svt_ahb_master_transaction ahb_tr[$],
                                                                    input uvm_tlm_generic_payload gp);

endclass: svt_ahb_tlm_gp_to_ahb_sequence
/** @endcond */

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
6N7i71JU5+6LAhUFmPgUpjQ587d5n+QfnVnMknwXWOhGOsXRfvAKv+Nio0/aU5mG
J0XN8nBCSiNcNvCANZSmfGZqpONrww5iJDZKMVFlneEjpiGPIf2p5MFeP7eSAiFH
a0AjRVPX38Q5lwSx8sAtczBfat9z5ETIZrKnhvD7ydYFLJLJbq4Xzw==
//pragma protect end_key_block
//pragma protect digest_block
MeyvlVtrVNJ9OgMNJQVqds5jO9c=
//pragma protect end_digest_block
//pragma protect data_block
4aWyw519be8aVaVPt7Wmrv4JMTUAFsPsHfyrdCj8/5u7kUIPiEbXCzN23DIyuGuW
hb8p3Wb5XszVH07HdCvmb3m73q7JXoAdmCezvsRnkIbPWVzFzEa1OVzRYxD38gbV
Xa0kgHsn+r6xqsKjystPngjrgiUWGUf+lwI+yL6MAtwkzgcPFHFl2XWipZvSUqjQ
UAghmDluBNR+aR/IqNf9SnBoJOTsf2WMFfsYLuRuk5IpHePEVVs1Mn0pSxfBrxZJ
1seNmkq0Zpz8ggqHP5pLxRZIsh79DKkGupEcscOopRWY4Uyh2kFdf/xpIRQg7vc5
qmg4jf7Uam2cUJXzCam/XbdmSdSqXNX5DbRGeldorHQJ737M++uLC8yRXW2qTNVu
OruJ7oFu/UEk7Zbvgz9E4VQM7HmkXFigGK2AaIK8mTC/9aZtnD7Oxc/e8Y+FXfeG
cmbaYq3EnLVGXQTrxUSPw4yjWbDMaVNuot2uTnBv/jNdG0mpBLHrtMcrMCR5kxfx
PKrFxnbtTPMOL59yow8fx2Hqf4TgiRB2aJAo97FzBBf7v9LfJnhSjc5ecTUYONPb
9UBWfZGvyxBTGRra5Q93Z4Ys74nvN02lJ7VJIscOZT0EB/YlCJj5zsezEnABwpCN
Xc/bTy3fqLJW7OZbj65SshYk3y90pK9sn+PA588I7r8bJzuRdc+Ezn/sGKfOYKoT
zXaXOXiAfSv4jtf1pA6E1FTgAPYndxi5ygJoZZYQtEYxJ+WkxapaGbeKX80MKh6u
IY6p/SbCUH907nv5ebJLvtezZ8PcILQiIIeujL5xsx/T7vXt3lDmL+RcR+kYv0sp
NJUUDm22vLyhmxgUzRXBoywji/4EhffJ5uVk1sOk9GIvbwcLb4L0o3v4NZsDdVUO
/ahkEhAqH0t0L8DC64IpjOKlbM6BgeZMhPoNsvEJla4nF6Rn/J+2skwCX9/z9yE5
+f3mYSLDGOK/uWgLzMCc6VQ5MRgd4OHCnZtpclnheWdeILROepMNA0XIJaekY8Xo
8N/cWELIACcCqLYDLXeQ78IRnknNB/TaIv5fZ2koNHs2lTHYHZLAfR2nAvGQvjQd
8wBUZnHQ6C0myqZsq8BPk42RQak3Es1Lz78C8kfKCFalJW4K8piKV1ByUuKSXazj
2k15OAxZyxMWz7aMt3q62Kk/f5LouMQgjBQ+gFtky7u5rC3iwmxQrEbk0caE9VWC
ivcIqxphoDlvoa6JTMdD6omiP1Co1NhRAqwV0/PP3HMb1Ja4PaHpx1spEt+8/h2x
pEYM+Otti1OZRm+4YKL/W0C4Q8sHnLYwrVFRkX7BMGdJ00iVNqE1q+VsSiV6qCbd
yZVOeo2Nb+wc835+TLcH9nRd0QW1yNfHJO5B6NI981HECwcWlKXLsErTKz9nDUVj
nUTlwSUkQkH2uw/vvCmE04ZNCiERzknI59sBlduudmrGW8P9YOUUvGY3ggh8NKK6
tjCfXMFT+jMw/CRJpaUeRSzX10F8JXo8ilhFlyV3dbbG7ZPlpP+buWlz1VPsAYbV
mv0agGVQXuM+QtuOtwK3YlOaPGBL08W/KvTKY3kXJs3+unSAX9uDazsMNlqKjGPa
LrNGiZwjrS0B9BxMlt7XAO/6sVB3GxPNibnRaYsdX8zn+d1C2DcnfUW04l9CjW6G
Rlk/Gta8+wlVaKPNT1rP1iDZRyz4ZxbEahr45J8gXOpCkZxmaIFbo4lbZrDaDzXU
aIq3x8n3nFcZQbpefoWoumX2IJrObzt5T1IfEmM/zdBn1W04atK8BaYLb/UCcarC
v9yWVUpZ/KPHoopoBY3jgAb0YqxvvDzQWvLbDZqrsNNnyuP+jfzK1sCPzdfUXInM
IcFmhZBFU1glSahWHhhKMTU9MH1bb2q/ipnBT+7ZCSQ5pgb7Id8pK0pKlS8XvhNK
AnCfNahS3VscpCiLfRxCMUefhWK7jJm8sSMyJ+HIku26aItxw/AqCNteIl8xPt1m
CB3zmfpBZ9gKdmh4aK7jIgXT+4VdqyGSBWC0MRFA4nYURLUJLi3jOBxQQi8p3ERE
SpChFix6hPruf1vnmppxouOAm0UExAAPs7+UCXDXSPsCjEI02K+nYK3/sS2mEerY
HG/lrXweKRdq2n8+jTxobirlBVyVwpGb6w90uVBOFnZ220dA+reEUNIaSifgC1ay
LezwdZqs3P2UaGwHEaY57ltr68mRxgXbL1NO5F0+e9q17YipNMS7jXCNdiu5FMB+
X3uXO4SIRzvhmuNa4lhnb3jwq/bxhhjZWv1RXgkQrqpHgytI819MD0sF170crefP
YaYAvDZbJcXnhymr+W5JuiMTcZAhl8WIOMQQADobT9L6yA3DhvxQc1qFgCjcs143
su7cOdgLmogxv0oEgu5g8e06I79hc1TCYMOJlIFcPuDxNoLCpjaeX68xurVpxcqT
1qSpC1fvt1lC5ii2DjAt5p2PYStXsTr7/TCtFCtWLybhDjPxJ+sqGiZiBvJfX0S5
cI7dJ/U4W+eLcBidCzSmL09bocJvTiUnZGL4csumc/+rvObmeAw6usiXP+8YvGz5
K0kPHCp+geDu/MwTEBS5NOAnYtVHge+z4f88h/SUcvoaTm9FLyNDmOltmGnCS+yi
qIASwA82o2qIfR3W1CK3qhEvD28xWqww9ubTo8OLAJvu0sXtPCki7mIqOHBaqRa/
NdgME4OWg0bU+FHNKvV8FoW/6eJXi/6oYgcYeM4HV/9zlvAXmP1vOVtE2dAFA3Am
UTx6cQ49mmDdWdLSE5yLku2lgEBeCcE1aj9z2nb13Csw3BsVrdJC2ND063bZyWP1
8CSMAk23Ekb4rbTXttv53SGpOuPvSidHoLjrRfHSpBGB/tQiwZ141KJD3eRUaUeb
fPqk/RHBELJ2f0gQGB5AiAJcSNLF/fRqjK5qiul6D1P9aD+kYj0iN2PT0ICBikOr
1XMukdyKJjJOMGqOdtHGqCOuJZvUjLDrWSpkdNrKu+M14BSkzW44ygKAjh6xlMBL
3nHzO5PETAACxGihoER4woq48taHVIp0QWv3lIF0CBmQfogkqFlGVvu8cWF6cy9G
DPK6t3DtATQFXLWVkHGpIZvkeJZXm3SjOzX7hxSXc6UvilTkyXaPs8sluBpngRmd
xY5QhXZPJi4I3zcqQ1H6Y/yFmoqVBb3JVx78ORYeJP9fdgKzOEFTftUFPCeQWyfR
q1FtmTgjj61yFudrPwIoxbbx/3kGljFIOzdnx0J2GmxIOt+nyNSGfUlhmyTrw9Px
WyPbaHVbjDuDovVAHcy4DLamlYlUwMC36cNBG3Yn0d3qrf3IR/DGq/VWvxDwuFLv
1ICP5sBbLoCrlviYhrJyedDtSI20Z+3Es0lG0/GY+nWIh1poNsPShi9vYNJByjID
1aAa/NkvB9wjeFMGLk/08GVo9CwynCPjx6/56wDPkxwJCHb9kWu7RsRH5tyY1aGH
APEejT2paf4Cc/mrSdWFGh5BJeUXrqlnK/BzyawNWlDAMuZPo9GUqcSFPrH64sBR
kTvvqy9wAXdPD4HJaz8hxHSg52q41EqOUZMDZ4w1Gp+0oPvalacHj48Z/0/t6+b9
AMOVZtT+V7LuFK+Is/Al/x+WM+sqE7/y0CRQTRRKHwis0J9jpOEfoyV+ZahlYrCe
6OJMcnvhkNyfGy4Q7r3oN36/0ateluokAKCDugfWDJnJkjdiK0n9//Fwg+NgAwS3
Ch/BToc/DC8IRVtjTXR+LbgejmGoSjJ0Om0x6Sf0UTcGuVZWOfAOCkWiPCmzDxnk
pbiBcVQZU0YkyS551MICOHwI45K20hOs19fc1iHV2aInlTWbjh6yfZzC6G/OnL9I
NrKgBmC7c9j4a1LZ9AsgAnshlzpkacW3DNHsuoK1xxDYHBvw6b7KQwlOR12l2P16
RlE3v7b+pdzaWg52D6uQ1gapWQ9olBtCNUvVgz2gOmERPVIh0H4583iLJb24EUsz
XogBjENbF1fMEOK1k6SPQhPN5DdhLXQ6P+fOFTfqZjiUcvGw2jJpMCbAVugGdKe3
N1oheRNyFblRByFQjnYObli8rKjn4+xYx+1INBMobmZ/OBBMvs4AsrwXwsfphjL+
/o0u99nYYDz2+Fk4o5fGtSoPTPJZ5fcn8/7p64Wbf7trENVz4rkGfR1CpU0onF5T
thBWHsAtX9aZbtsy7yhrHxp8je4Xu45bsSro5o0JhyqoVNzGiPv7yGY6SnZQvopV
uX4mJ8OTxBhGa2I9OT08HI19sIX0NuE+GNFBlgXoaxZ+Z8//jPJrMgjvS5GOTr9m
uxui9EXsCwI1Dnd/xn1bwIcj7lxf53MQkmRboxAhikIGWNPLwhHOFuFYthoB77cj
+VfVr5/k44BSOD0l3ecIVwFDSTkqV+03f0UAv7/qWytkxtaChZATzYH0Pbwnor7y
grudMmo7MKTvK7quRTn48w9KUuRM2yvp9p77lfS54ZTlxxeA1J6uF/aNt3GJg0KT
QBSybN+h3y++s543LR3+YR+hpiN3FsvUgZv35wYzUoWxgbvuYjgWRb9gx57QXwrS
axy1/VSJtnjSZ4T5tknLeTczf6Ex48/nBEUYKHtMQZEbXZDhPePl+spliL3qiuWf
C3L8MEPzvbjNp1CVZCgUwt2l5+LLMv3SUnBuvueP2b7j7TbBATRJKG0XNcVMOI1A
8bm5DdTcfXhg20K+Djeunh8qlg0+NDnydPNxQSoQyLyPYkbu4g4lv3GOIr6OCa9c
bUTn/6TZ48CWRwP+shCuFCSz+LqOhCkYEhKDNWSTXn+uxV2FlSd4Nw+7nngvraCJ
7ytMsUGs2vB7UCnAvpKzpVuEwtUvPKvqeVAAnbKYxB3e2I27quoKvVg8eP3BfYyl
blwHq6ElmKyQQNcTqJc1cxHKuL3m4d8jaVP41Lh9EQk08s3BXJVdQtkVFd2MiWBH
FfCAlu544Y6dyjkcAA3dhR7trnFFX/tmbXolk+pMGMUzI3xArZXjhV+6BDaIxGa9
vgAzqsHCbJukUh4YmKTFpr1rFX+CvrnJW4WxjDVavpU0A96SDWYokj4rU638NkDh
a2EVlcCYBwFiR+N5ecE9zi/UXyEvwTQ4NojcUennASSZ/M1MqLSEmrepPhFD3OlS
+/hBLfc1cH1DxGhppUSX9hGddXNmgH/ok5qzdWb8yTv9EXJ3hlIwH8kZ2tycRS3e
+LxPabcolmWGfpElhmvFWYeEqK05+7xvgc1a3i8oyPuvVBNSYCHfCSDV5S7Ut4+H
pMTuIFJiUHWg0Ny91+Lqh90MNquDQl1DJePPzX2EtLDwDWnlonKL1xzGZ6oThkKM
e82tI2mFSE0T+dXGFg/X1edmqyiCK49cykdiX34Xk06odY2ap35eeohXIjx3CRxh
ajpYVwqvRqodRVtn6TzfAcfzozH1VKKJQIGo/NaEpDNN15TihpU+G0VemIl/fnWp
aY08uH6YJE8gsz/eqhiWYvIUscWblAKUJys1f8VbEK1UuOhFVuT7mta6TxtyERgX
1FN+Wr3YenWTGxHtVs8mrD5hv5g7zKZYWyyKYgCElTQnpw5ql0Sm1z3GTswZJvbS
8MMmajpDWLJncB9+2DG6xBZFzuKcnamrt747WW4ab6EEGRrzpCvWlxXPQ7DIAcKy
vLbeS6RkQW5ednEJzyQCY5i9rpdIqi0oehPFC9i0/0v6GCeNJOv4KbxwmmDm2En9
6aDa/cPyqTYCAa6XNnYcvq2D1X2DSr0azNxKpnkI1hGKFeP0trOtbKjwYoORKvGJ
i+lF79Hg+ZGCylY/mD57XqgLWHKoBE5JCjzs2U3yeRqf7AJjC/NzqRqb3bw5Z1cN
jyBi3Gzr/oZo/liyik9Z+OHWqS3Z3E5i1/Hr+EDfARGQWzz6p8L9z6+tRyFqoZDd
+NwZX78rDR9ZeKudfPqi9UGH1b7y8nSeEptxfWUjM4ZP+ZGef2dGcfJ1pmJciegN
1/eFmf5tPFcl5o8BwQqYZolelDEJ5m/Z8wdGGOyM6dKIQbf/Ue4rIVwWQjwtsq68
fgFI1plQR4iHVBTEB+5qz6lz0VryaBkH+zcO2Rao8r/uXiNT9Up1ZweorNmlnjt/
HY342EFWboGaq5UHaG40ANCwqmQ2Yk8bPpHzKcxvNlrO4SzwswsNNXVB6tYI6fcg
d5yZiLbAPvCSBrB1bdwh4NtiNq50eg9YyqguFqalZh6REa3Cga7lEg+jMrs8jCDh
+W+GDdv8p25uuRQPyqt1YPTMp99S3NLpJ8siGS6xM8x9zt1aigKJ6WhsuPyc1hKi
VVh0wT9zcXc+VUwh/FKQwhmHv3tYYzgNY5rOH3ATpGiKyaUC+LCli24dYAuFcPC+
M1c0xl66Y4t9tBNMKVbwEv0X4qc068q97wS7mVKWzqFNgqROlFc1IW7FvarBD8DJ
2ISrm2NuIjrzepoItb6OjWqg3US+yT+6TCeK5raNQrMveEZUCV8CuxgmENnl3h5X
rPmxKM3ACAT4TPf4hb7UIl2svGWXMFJepDc25yeMAZURq4X5H56N9ugfQRYA+ImM
pu935SngV1/VyeS4LLxeD2eBOToyS/18MMyIUV7+peji6h/y6jScxYsAZkgHTEFW
NOwxoZnNqlIeN3yWl7TyiUikOKn9jIWzk7nxWaS0Zx6dqa/oVASnsw3M03NRs5AH
/V6JV6PkAo34bKGb4oYl8rPDLXNFHA6VPjXfqCBY191FgbVO6TMoC6JeYO9KH3Ox
DUT/zFeqaozqT6LNItjOKw5jhwlxoG802R2z2mpyruplkSKAQFlpk1UMaKTLuNyi
CJ03VMFWLtfGO0QdEZOdaqedVZHYr4LMiLhLiYJIJ4rtqQDWjYTniXpdOI4qy33Q
YimYiUauWzAeQ+cOqd/xXc8QjZgJF0UcTKSWiBPT6u2d/l9NUfadnBQpQcOsSGEM
kY15toeR4dg33QKLErf2+ssl4FV2qSn0dMeLtyTyM/fJoQ2YbiMtG9GQwKZB6CuM
Wok+8xOgaM5/SCbuJIwIO3l957Dxt3tyIZo2qBz6Uu6U2rEgGYOjC3WU69zFFUjX
lZGHhn0v+uBQ+CJ0V5rlSeT+akeuMI/Lv1PrydAMZaNnVHEVuOmzJbcqINJGWN2S
2TdV21G3khucae2gKcf4CwVrYYsVPKE2W4j9kwSHHSQc/OeJ5vEabVXU4YSlCXzf
gdVccfObt2nyWJq0AQBqc4y2tHEKXm+aBpk2eotu0W0guGfBZ0ngw6CX5ttvJxhz
p9s8tSWS3UQ6m2zuIU0Sa4waKeMrSTjYFNMtzkMSg4rYGlGuQwUZ46Y7oTVzp/Wo
b1r7ql8tM0lclH6G9eO6FQJh7/ik3vsMm384ycITayXLnN0epfk8WjFRPbBZTB4t
i41ZPm8yOqt6NY19YUkCOKx8KYtysRdIUsomRR77ah2gtbYJJ7WmE390vby/mkKF
pe/b9keW/1K8JQLp5Lgp7ySew5jijfKnMRa3S3YQtdc5Ht1DZFUfscml9TyZOhKb
alGf2178b6VY1mMNby8DxtMV3WX1D06tbil9LEZAnv0jCg/1Y0caAu05ooXi1ZTf
VCHh/2cftXf2FgDsd3HveNqxSi1GotrKau9clreVT78PcLkLAFlwy2YVsog7snb3
9NHhV+rOkzxNK/G4IRBEiyuvTBepigosvs9TGDifxuc3JtDwdlNnjsmkQdf+owf9
+hjrcTnCMeF+8YaYdFCE4SnoW7S3D+vUqYU6v4PhUi58PXEtt8qZ9xz+DJ2pYXFh
wVuZ4+lxjkMR+FZn1FaZcOs+2PVZ4E8DLn6yFHgok8LRmsxN7+Ek54Sha+zxEXjR
3wyjJaKb/gB6/5a5wjOthxcRqKZwtT0WGAj8x73m25mdxSyUOimnqTwT2eWf4n4Z
eg2ze/JPQqkf6sZLnxVQkTweokW5pbkIQNb1RVU+Y0oA0NK4uIpFGRRv0QbvRuJy
OyDypDHZQcjvFBfWZO84X6iR/1W55MokvCjPPROHCGe0oKo21XePtahK2We8e9iL
qzo4+l7XNVS5Ss+DTq4k/oolyJ3gs12AOPpc7eYGnNWHbfyyfyb+OS81U61LMj8W
vCZLb7a+fTYTf7OUdKA1Ca1Kk4DX/4QZEU0Bfk8hy1pbiuqu7Kv6cTcGZSxfTsAj
cFe//Msj05nqG8HLTWJcu4tQOCdxR6vcRE+uiJabFVZZBEXPv/XSnGyjSWfcVrTf
iUDzpq40a29AM9W1XOZoOWTmsF2BAPKoZpluteSp4RlYhV6V9EliiNGdAtTJ7Wtf
J6kQzic6W/TKqSJ+dpcpGOVLCpheAW1noUWAZbODntQpgUloZNOBJmDheLM5VOo/
0eQgPLqU1MksU6jXFFUatWavlZE7v604I8TvHF7XMWWL/1wLTl5zDaCwtjmpE6gV
XX7Zg6A1mmFMQ0H68KOQ+0WvIhAsyMTI/X4vngIAfVvzOIXl175vE1xed0M9XRqJ
bwv4/eO0pj9dE66ZlCBVSZt/Q2GF+Vxg2pqtIV0cKm/UBDz/iHI/EKyqP4+AZI26
TpegYBPBKCyn9I478XFm+Icug/aByZqEIguU1lMY9T9J37IB7M4GktbAZWoQMPrU
447epde5vcAjCk94dB6uMiLfawjZl09ZS7dEDHoyss/z1oMGiXW3EOckvIs7AUWl
2huZQ5iGMpAz+UI5Ad0QABCeJn4nzZ/LO9vsete3OMQbnMoBEBuDm7J4aIuAZze7
3tul1HflFD0n+Zcfl06gEoIaDYVkzdm+Ea+NYM1mQ6XTdAg7IMH9bN/c7cvb5Mo1
cCl7jEiuJQI3HWOp5F9AnRIXt51fdeMHiMqmdDdw5x+Yv0xYesB5Dp8QB3xVqHaw
/uCHTT2a323nHgcrW10lZ4DOl1npVk2/G+dXlcN5P5c/qHYhsyrxNo2LqJf0siRW
96CWvp6A+RJbwbzNdkBeta6pajYeZJQY8jZFv/AFlPsg8D+hwpP+E1f5KJy2NMAf
RyNN5EcT4kBwI6MQk3fZ8rFPWniHw/g8zSApAgKmu9k6NgNz4uoMT42BDePVeQLu
PL8RJVoKA7BPLK+9ar57wJ9KfklPBa/WcceszLLzWqVMky2kd8fIYBjQsB+kvgv+
5CC251W1438SZBHppVdBuUi49fH/TVthE+/Mc4SFE+LKY88CFNMQy2hf1CTQpAFJ
OnJxvH/iz1X8QbOtcb6MCpShL5xYTczd4F+F2ftxB00ZuzwdFu2ARY3T+cc+LXo+
J28E+Yhme5OMtrY18mv4gQpcu010Rhv2sjGYWeLdNpiBWdux2kHbJ6gIhhBpCAQI
kHbzJRcbYS+WkU7ytpZmT7lDKGOkAec9OTDhCq4JhGyRcfpwzS2sUOZBtk9lZBJB
arKWXqJAmMzw/FRja5AXeGxjizlBl+8rSXwgcWSPnOJ3YOxCFpYXyxTbLBezVAGf
Xhc76RCcNGOjXAzrmk5R6YyvoMIYJ5VQxLzB8+lhiRv1IryrLZvEVNKLjhjNpseI
MFyRWfnq89h9KqQti8gKSoYevoikj3qc1mK+bWvPRosb0dWwrqaX95qtVz0QfUfa
WrbYyzC1TIjtmICE1poNfsb3xYl/m/iGCk+jjCCj4ip5LfbwLgqHEHKxFZVru6zr
jkMe9Ci3HXVI24KOtI2X+95veiWdTykc1XKDi1k8UsMg46yyB76SyuEH2EuDheet
aT+gS59LcE2/syNeKEso8+pWSxtoywWtJWMu7sPKgcUxfGZf1r/aXOgJBXfGrtS4
tluWLzRZPMc4OJ47MzOgXW395f0pT2uYXUSEose8p402THvYVlNc3sgSk+867/16
R8nkStc7ldzSj8b3V8rnPG6jSfu+HhxACO/h5jxr4pUPihb2+Vly6sytNAQrfgvp
Xgr/Y+xAoa3AT9ewzu4vqgZyZJk1IpJeTzkra6DbIqHRPUN4CD34lyhwSjUoW202
qmbs5y+v34dS7zaI0qM2TJf0su+kDpLk3IPw+F5z6ANEFV+1WN1t+eKqybVRKhXU
wwLOS8IkZgBOTjGEV1d+TtP5Kf+ggvxNDKZgpFfeZ5XbV2ooI3Wo2n9Mb98PjufD
edd8Ye6idIwoUOrHT2hr2SkOpFbGiXdtLKzYaACm0eeeoV/iIbnwO4x0mgpIvnHw
FL8D98ONdl2EB0BppiePILAU6t3H7QFZSF5ubeB/A16lUFEOvNbpZqKPtKj5myn3
uIB/qeFwq9R8jougKKbcS+OO+B3TcBdWFwciRCp91YRNmRY/B0KC1G9UA5Cku2vg
DuazjfqJvAj4SzChUfJwmXra37q8yrrHrbs5fkUMB5Y/COVlo2uu43q8kSIFAdOT
Wjwmn0bw2MDVpMheDbUTPz9ATCTMEv0FwwgWoyRQcbm2QEN5mfNVvYHJ9wXjlEcw
WypYBmu4G2OAzrZwW+XDaY/Ap7b8Nco97LbGw861kmFPqnpVkqUbUTTeLFMgbc32
HB6ml1rtOzF6ZG8rZ+Yj8VNLRqZSFp/4VGRxJLEke0dv9Zpl5TZP3a9+ASMtEFVV
RocbQJZipBXShmUKnoyL9n3UiRWSB4rAnfOgHPvUc3EKQQbBSjdiEaSYVzyQGmtO
PkDovoLOTA5NKrqF5azwbK9U5kEGOlAo9SyDix6RjqF/Y5fJc0nryHfvK1ZDQ/Ke
BngGSNqgT5W65aftY6R2MSCq9VM94fPETN7uGw9xhDlzylOUxxqI2b/1qWkzTZlj
B5AhZ13cay7C5fOtaSVq5UwB83lGTJ1xG0Q7sFh/AnyDPqgLg/4VVGWi36xNymuL
GA+FnUKquKENwYUqMjEY/PEcCbogY0keDDWeem8eqqmivOqYqOZ8VbB45N46pUao
gL+E9J0pYkFBcE/eN+2fzJJLNGswhLY9ggl2zIUDiOs/eBh4BLmgeypkOjPhdzEK
cm8qflzweuUYYPUF8XZIshxPzBEyW5yLAfdFy0DmL1xzSz97M0ssgWwYmLIZz1/g
MNvKe/e010f354yqE2C0kGtHiYGVGgn0F0LVouMK4F51wWCYpmjMPpv8q7O2J2XV
i5r4D8ErhsLW0CR3o62zU6UkVgBn7HBFCWtOz9o1AxrQsZSDY9K0YCQNQDarKyf1
JxFFdgnK7vhLDPqPflKJ50osWDviK27+G4/wTYyjZPEAU06gFby7VK/r3p2EbNiN
zW2a6AEF0NS0wC4gpssEJUuxheZuiT2Vlp7TeEauD6wfS8b/x+WKZKcSQwxrn+QK
H0tkPx0VcFM/BTG7aCPdWp2N2LvKgU9J38ED2eI/WUPaJ7ftoVgsZGYjlqd0pn8p
y6rITZ/9OJ44vM3JB3/xsKRnK1rpZzJcfB23yLO71DJZQsT/yY+Gl9ys32sgd/Sq
M0aD+HOs/CGjbYqn/7Zoc2Z14CbGcIFZx8GPovVSBOQHqb/XUNi3ViBNMJZFh6Hy
kRAMVKBdlOXKdYnsdvjkjIQhkIRMK542ewhYGefdoe6vYyJu+XYWeHAcayiJC9MB
Xj3Y44GKeh+OQnECH817JsSWIPlJjBXWeE3veZmXBYesXtmSbpP+J3h3SLvB9S3w
2OokDubMzJ55xzRNFGJaKqLhJdJWb92yaI1X/bD+EgXYSINzVbMmYJqUR9iRpu35
DSe2004azM0u1HKBYQk5Pbbfo09iaL/BrAhfUIdcTJUOn+4akCP8I3AoXnaTUqk6
GJ1GlIDcdAnnZthZU9B/7Ci5TtRovLhTPxttMRxA7JjUXD7W5hl8motBVmFKWaok
VHlBfhInEfcFTAfCr+/CetEJKHvZkNkTg5a8Aep+6OmjYAmhFduQNO9jxUenSwYE
PQNpLAmjUQwhKhGp4rGicS9c7+FLRrK9G6m/9HTR2wPMJTxGySg1EoQOTPAjH74H
alzAnoaVU9VlBu6kGfHSWyR4ljEldq713szmDaDPc3Ge6awX0o+Lp4Ud2cCtvM+J
kwfQ49Qhf3k2xCbCZ6Y/1SLbX9uylecuxLMjjwmMfDgLZgIChAo4HAOFPgSd8A5b
uzj/8Or0yY/e3mWeVComky05DuenmeYNIW74owboajlTm9k7w9m7DeC6dtMKe5ZN
AjS59G5IBc6T8zCc9Bivj02Ob0IunaVpyP7gdrVckYsZ4Sp5YTojUql58L5RGrLx
nbGZPCRjvX7La0WKmkGcGeXzj8ieihQd+BaVlihPJA8cC7a2w8pjWkGGk7MV6VbE
xJi3bzDIz1aSLmDRFaAf2GLC5lrP0Pw0NqDDuqd2i/zV+fVmKWyMLUX+Co5phpMX
hWzdYTxqEfth2x/Xhbyrc0zmFuAB8bZPaCdXVRmXSO8pC7ah3nGHWMcwVZGOCfeu
LbBrUEsIbADgiOCorPMQ/cQ4wuzAlsj4tDBf7y8A/aUbVUY78MBJrue4JPQFxAH1
nMfquBXlYpC8WVAJsYqPCCcI4FByh9sxxjJnpP8Nk5/EF8XtQBhuwk00T6lkjaGQ
pp+KPG7QBBIOVNd7nOJBXibm2GOSXIDaBafE6eh3nyynrOYkd/ln1ptfz0Lq//f5
gMufj+63s7BhxOnGeuHtkVRl5MrIFkRS5UcfMIwoernd2rL1eJJxkyFtntj7Jmzd
2EeQ4mnMev0r62+d7+s8pAbauxe64xW4H6waUwwJJMWuw5+IlcVKj948KnxZkzT9
NbVhZAEipbVV/XpfwLomsnqsf7s0o2e33OBv/IvwPJLpfJCHYvyL2huZDOrRiAHg
EwKCs5pHhMn/BlPpBIqPYB/8c2ey4S7l3tsvXsPjMpyz92jjYjxFgDmGBtvTvq5Z
LvcDvZsbsFJHVgLrnOwGVYy7OAjCYZudn0KUp9C8mf1fsOjz/CBY0IK1hP8qXnDa
tqrnE12Tgyl10iWn9zcyUnoAj3yMflbQCzGNdAV0H7AoSbG556rYliTtQOT8Vjgf
uA58HgfUc9bLRig3BYDvr/sOwgXWXN7gfkMBsefL9iBDNGulQE0pNm/gyXQIUoI7
RpcviyhH6/oJisrvI8m7MD3yJLg3LbJ/KnGpUhCmom7zH4Ygv5LiHcTR2HxgbSdx
EBrf6KOxs66Y/NlKwznRnoTWCJQ8RLNYWFIF1omzDVZnPsIaKBgYzUV34m3hS5pq
pJXtu/Hq07/u9qfSnyz8p4lWDZ7gyzRZLS6eMcT5L/FbhgwigzKwBlv2RuX2XWW4
/6EcD4Hb34YAO47DOJNQbGrv5v1QKS56HjzN3DWDNqMD8wZilY/x4foFpREgVkZM
RiEKKAsTc3hnhFnwNqh5ntcfiNwPs9d0Ocq9R1UyUkWjW9IoaIHhyLOSLxNcZHYO
BjRj3T4YCymBR4mTwNNDOnbqoLLm4fTH63udFCaw+53k0lAU5yD3dxlYjvCxZhE9
aDcwFv3XuIAblRHW5iXSlsfPi/gN8BGookAeff5C0BF6mEyEZKKltJVsHFz4MQqb
nKr6QWEgAQTTqHReu2INPnsEf+KwT+3GxF+khoVW2naFo0/A12zZQF/6vr96CedI
f5JJsEIKYmvQwCyhsQFZ6jdBUiZ36O0Xezt2knWsVJzYIZGS8PkAiXanwDHfcDeU
7wXu00h9JOPJHKcnhVQ7CmtsHzDs6AZxFsSfXtMMh9cGf5ASnCvgpnwhRxKxyioz
UIzqhP89iglG9VLOrmdUbvDjlY3s+pIb4LnvxCUE4lA/r5W284kfVREF6+nbeZS2
JXoJ+aPl4AUQUFurvWSnB+DOblY12y61oxpLdAbAUsqe2bIp3x17ZeaRQ1di6JxW
XYQl+lvjQgeWZlJFmbs3Ed0Ho4cADCo6wAu7ke4wtbFypEscNpg5rILfdjvh6jQT
uNGUW5LGRh4lBv35hNF5pCtSwRZhfXPf4VUaxmTntBxKxCmNg2HXdAFk6fAQh9GR
b1IB9v+4QmiZKSzzn7Necv9A/KdJ8D4kCCdJBRjLtLafLam3vgHvfRuidn9bLiZ/
y+jdZx5e/z1HTYOpV2pf417r16zw5ecPWRutDzh1Kk2//RNASwoZcVwcWG7bE/fh
rsSgBQgHCp06EjFCaexikwGkdVk9u6qbUMsrq+pLlkNriWVOy0FUQCkZ15LRQGty
4XJb91rbTfjRSLIfIPU1tIcpWTflmOH5POIwgRYMVf1QySjZXYMAdw/A1levrOEz
alxan2n58HMEsPvX75/fKUvA2FFwDF8TNctKVgJY5ih1tVtRq22p9OA3j+cW+RSP
CFqn3CQ57grpQ4uBr4nMn8rTZ6sOJufz6mRH6iBVcRM10FYEYWPFIaQLlxh1511q
0zUYYwv+Vub58H+YAeWnHxitnCOAe+shpCBXbjak34BZ+4DtNN3+Z5qH6yRwDHZa
lapmqYKGnA7mXvbyEg0rOFoHgC2+ekbmR07evkQMYYt/klngu3avMqfSW8jawOvs
m+Ha2yXzHi+GYvG+bThPpV6BNsKxfL4ixzl1e+fj+oNOoRYGWOXI8fijwz8e6zTo
kgtmgu9c0gKa/CYLT6jhZyO/GuMdWNdupAJxKM9ZuTdAansFCv/KrmCMEpjr8BEQ
kf/KBFPh34pC3kyXS/XgVeH6TUNUJCvDhBnlYJf4EATFymVRQcjsteWENo3uRusN
FZbWRbrdIulelcAJzupd6Y+8eZtXDi746vj9qdzHfqIzwF5Gb5XlTlnKLNAm5NcI
XiiKSBUtqPyHgZjGzz/SSJRXES0w/Tl2ojTEFCHnNV+5l3WjxQBQRSAJHv6FcVeo
HaW+5vwt8WsOiByZKZH3C5zc6b8lyRK89OlqmN+Qts273v3gAM4C+jr56sq0MXTR
MPi/KAIRoKCbnpHRLrHV6PyUzm8MpZZHG+RCIvk+b04TwJ4W1/mBDMeSD9X3wUNU
KY8jic9YCpUUsj1DmHKRW77FqbCkj3fqKAdS4DiQG1+VE8SNYyx7GAzPJWSwVozF
CjVOdJGY7/4x9bLrZznV0iAseXR58fD6ru3/or7dNCTnC1qDTAcTosmJ/lZEUVDH
I5jntALpUNamyUOjNYNvgTEp4Fi3wTWA8s0dpwW+GwckXe//XOpKETGm9wgac+qC
PxOKA2G4mImaYrgziAVgVy5mZVyi5C/673iIzXCoo9W1Q8autnz3k1Rwp+rqjjOk
XRy7ZeJmh1E3VosBVeJhEUHyz8CQ3JKlQq3HuyYhEdsTvb6rRvcksFxkoGSrsRxQ
FRhMGGmuukDxg1WQFeSFlpz3fvlKhTy7LS7Vm5XD7RLCP5hea4r76rFdR+eLrZTU
nCM+3Y9T++LPLoHftiNSxdRRL3H0yTWIEBQUSkB17SvdfAhR4sEj3Soy/rOYiWCq
lZ5HV+LF98C/4P1tl7U0oRnocugrtxYcjnCMMr5fJK1YJvsnazYj4vgwYrlXxuT5
Ua462ODzbWpRx2XSxQPfDsQz2wHI6jrFVOt5Dg8cnDC1k0zS76aND4qLcUmXRAb/
cvOYcna9mjxUdQsPozQYNhp+Xc1p3xO0OSj705ofh90qL3geMtW6dn2C+Xo2H70m
cYOODbt6vGHWqtRJ0jqhxgZ2A/XK6A4dCuy8XZe6Rl2eI7ucw1rBJvHiUpamNcFA
Kyq/sfop7LUz6PjVlmjdJwniIvtQrJyZd+Cnpxz9b8DpTi+oT7NLm2BQ/inA4wnz
DROErmFSCBhp9mStMFwOZxShQR507BkMoGL20jQJf7ojIlxfh1AuciLE0C66SCYS
4DQ0U+TEVd5M/L368pRBLjBhUrQ/F0A8/afu214S5L10pC11WpKP7PpdZZMdtpTx
OX7I4uTumcVXHW+j3TxxSylF0eRRfEIKqUPn4+fhScMRgcjOhg5SJ+jQvrNqqRgV
TOL2H9+DHRmkaAUOVysNg6qx7q55WYqKJ4j8TeFGvxsVjUpbjFbu4VxSUBsRlbRz
b/PSkTxvlmhkVevj2odpx0/whABqQpAk3xouLVzoCC2hv9lrbsAjHe169uQbhId5
XzMgPMcsPvAgs2xksE1WGTUo9uB6JDBBrcri8e8TpLgo94NoEcHbe1ZGZvqjyLv1
hXGAUhB4yo0TTK1CH/6M2S2d7iPvtx60fqBb49eJh//SVt52Fv1WH4LnNoKXyJ5/
4QCbLMZsllSv/0OmsKp+ezfLt3ZQe2dXuJoaCPVDIf0MrkHnPvavPiVsydDxBZ52
rcXynwmT1tXwQFBrFQlMpQx3iehtJ6Chy2ZdWcfsiMcp94mYQDrnf7DlqlQjgjh2
0yqbJ+LnDb9kS5nHx0TrrJHPxjpLlUntn+uPlaosBGBjXC7e96FSrmNqbEvbSmTS
T30xI8nCzsWvGLKTtPsu8HuVKjIYsSb8OetqfK0kXrIrl9OmXnKGuEKXxoNxGn+G
MM2Q7PQujtyxDC0S3XS31P/mujDX7QRx2vPMCm06z3by5vNWBTxV/WE95ZTsQA+5
UbVDo/cG71ZBtk4Auw9Dfx2zGuUu+nFDs76Q8DKxr/TCLrwYrbwNuUvkCup1ErpA
oCFZSOYwPafmTCIBjMfdYFt3+jzlKmdCGTdzdEBi4xZlUxKSddo/oLkeVYXNPTVU
FEUVj92rrG2X8nbIY4/pakaUmxztif+dLOVNBMRNYTSUyZuUYZVudi3rmObPRm+R
IxAuthyvWggluXEsleyH5W1EY/JIFz7bwYLxCuCWpNAoUg18o7KeJhuolUzGbPlu
XaRclMRHCuXa2jOhQ/shT6GCSwebRYHQejZLt9zVwyl8ltrW6hdK+FT/ymM2y6el
VG5jlqXY0iUl13JNfe7KG791LzmEZL4FOWr1hJfhFh/S6eeXiQSbhbVsNr8jISDk
bRwZD7BniZQCI0q/Lq47LiWaowS//e4d6Q4zxR0Glc7jJkDLw6dbEh+uG7QwbOoK
GYyFmf8yD+1gMswMXK9EnO4cqnmEyLcj/QDRXSg9xzsx71022WISA3DVE8yhZWmX
xdWv6ttw+qtcs2oUuMaZjEiajMxHR8zl8OYDpCgixUXA+kX91xPV/2dEknRmpHCP
zmR4wz4eQq6IW9RuzwJfF/xvQ/8lX+qFE6fBQsogHDrK6BgJf0MUelZE0dLCblhi
qARrnYb3Z2vhHwnI86mWb50B5d5/WQXLU1q0J+Tfx3TsHkfllWLUcUlVg0nKW+W0
Alt+D1LwQa85qSblCXaEsRTLAYTBGzg9+isP0kqVMJ8UlONvoAZ+92deExnUqPpr
XpAfTdO40tL8zarp9arpFFMQXk6LVy/lNxqOrpFn7M/GBsNkNco7v8DVu8obw47J
IcGG/JGahl0kHbdUU6e3MStc/RE71u6pKLNjZuXI4yVnN6eaZ37jA4C//C0q7Ya2
gqUWAOzH6+ccAQuZrQzS0BG8OaxN2NAS3e8AEtM4m8SQi0wP7lc8TBb9XeQ/BUMD
meOzGFfUk53DvZyLDKZ0VcsmX0Qn5anL3ac3qE/aIWxOdrOI/9vY4jYk9tzd0o/T
fs4FI+yfdN2d2HjvJgAQnQBJLUZzGEEcoGf3j1juplwhaL3faEIVyjUxgsmf9cOQ
NlE2mx54qIleFNo3rRGRJnT3W5awzJiz+yXb9tDVb63lI20DMZBt0COpEzasF71V
KuKM8CIc/YONogLtiJGf1G5wFt9npHq7ugkYDsQF7x24n4pYmXHogRdGqrDG6Q/d
VqVuNHIhev9d0eL7NF+LIRUP/x24avg48ax4LVj3G4wYPbR8SNFyzr7L2M6wBpHm
q8N1eWbJw1p3/ymZ7eEeekEFWVpRoHI8tTfktNYPqxbmmN+WK+mAKxpJ0K8MemiK
61J9lL0znZvW7yOIjsdxu3S82zP4fSAv2HqhGEXGxdBSF8bKJKhkKpMW2u3gvdKD
iLiNIQYtTNS6LIi08ixzIaEBinq0YYx8SaElYgxukEgxWjwJgcG+Ohwt4AXyFHsQ
gzr2vihl9CZBqDVyHDgzExPF2U/mU+F1t0PynIkJ7KE4f5O2ZPzJLDg8sbcDS0Wr
bVbch39aekeWhL9Rg5gWSvXRihpAX3rYWhdUgR66yxzaPX/IE+FGN1nssu0OTM/A
Mrkd3kP1UOm3IkbohvVkesG+pyj3rgWIk/bkzJ+l6hiHU6aqptw7qLRfGHoVSzmW
91lKwZWN98mz14egSIqqpnBc/TcaSbpaTGlE0gntHV02RXxdUM4+2apEDJJ0MwWb
6ZOuU1KgutbGkfYdt+LU5D/Aaz+571RvwxIYxJuIAjkBLJ3D17m5DN66x67z9C2E
HdXBm0dPOoVlYZUjaw9y5gR0GgP702JyoG17I2jzh7RXfufGv/qWOnjQHWcLVGbe
m267vgnl6e2oJHTAHIjFDrrAd4o/CmKPeJ1FKgGu7aQc1IUwKEnLcoO0UYmyV3FW
KsQ39mSNAM4vHAjugtuMyBeUA3Ojdst1T3XlbJFLik0gvqZXgLnD+KV7rF1WoMb1
bkbLHFieej6VsTQ+8dFYLR8eljYEjkJlUD7jgLnWg9XGdXSNYndF4zJImunFylvY
DnRAd/Oaah3VW4B1vuQmQVUdTprCCcGRKqIBvwZfqIVXnUuw4ulyCUKZ6xiFhaLu
o6xvqfWnlgD6z1BYN0iVsABM+lrAB71vWuc/c9JMCFNVtkVMgt4NQpGxbDsG4VBA
VhRk993DaEF/nqBdNgFXooFLwU2vNcrASOZwd+7JKMC3r8hLaqV0ZcKNweiPCc9C
rlInBtWuSTGaI5yGOsKmHFp9wSn15Y2KS829KShc/NU8eeUjpGkLkeYJxA5aSKNx
5HHEJ3r2DfzOjguBrC9hL7LoS7cLNGkfTqthS2R6VdlwqGL+kB2P6VnvIGn4T9f/
8HCwN2YSd7YDMD/9BNAL5uk89r65S5CkykC7C0CT3AoaqJjZE3NniB2YmmLoalqG
ZW6QxkTu3dwBzmG45l4sDIIySzv+8tLvaj6ZOiWjhCHXdacv/1DeCCBejRSaEhCc
fxzxO5szNPdL+uEe3JxWqENOvPUol8BQjF4a7Iyys8+M5mVBcXmpDc/OVmFCAX4v
kRPpDpO1ehpZQ/5xtnCnxo02SgLEJ56Cq5ePXI0lm8EoiqCOlIziHYUFgqvbAG9R
Eft8ajrcwXeTa8G0R+4KkEtzEPqSAhNmjucST8ho/NFN/fBEnmKZ541fycNeUnNh
r29d9bMt0sficl5JHXDm6JfIJ3A32r4+r0ApZ55TKMdUSBu+w9rGFbdWr9lMhpd2
wnTyNU55HZMUyIn1Z37Y9q5IWpdKrAkKFEURf2rYbh7bgS8IzrPH6pZsomoZ4We9
jpt0tNPrbcnbZ6MGj+cZ2rzSLCHxZ9jyHHygKhEBwEqISz9j7IGyCdJc9YlREpyW
xh9pbfwr3Nm1UqHY6myFFY62905Cost1OA270VuPGzlYyZxsnRYBD6abQZErq+dK
DMlv05ILt4aUvvG1t+WJKg8kHW6u4msm4sbqpHZqa8hUyh/fgE0DXdO1GNle8NRA
OXz1K1g9SOVV6m2tTQgfosv7kCrX5YNCa9toeb4dOMz9mHNOzOiMNA71+Rh+0K1K
ino0CJQRH/N8LMkZ+X3Ikfln1VdYeaxqUIwQ0OIgQOFBrzwaonAteDfo+T0joUqQ
tCMbgI/PgrrSPOeGc/fZLArfniR4ftDyx5kPwagUR3/K8mn+cAo9aOrdJsrkelDk
kEXh/m9o9+7JD49c9wS7RMZOIGckKxSFLi3Y8mGybqSv0tLCqyFnTy9dRbH1NO1M
PL+z3KQ38Cab5A/szaeRLBnWoj1rFRLtjlNUAomNVaO+oFVDzkjBVN10FHn6FumI
12qo6nO/9L5Z+HGHxWGXcqDJOsDOXFCLkuCnqT5JJCrSeB3eZ0bCqtq+ck01jma8
p7pzo8/WmVMvrHNsx9vJuKNIZiLYkF6vG/E3zCqPch4Bj0GRhXZjugx0w+BJNCCU
nmGh9ZwKfZ1sno5mgfzn2cmAC82ZF4WxpcNMd6/NFtBCpSlc5DBV67Al61HhoZMn
oAGXzDFPMExLvY3AMPQeqnATNjxaH92zrXYY050P/kvvGb2OQt/f3oxLZWWGErRV
tUBpEZMRkFTq6rjMltfdkRBL2La6cpftP8nDwuqfL0gqe0tYSnYt3Z4bx4H4hQhM
X2TMuo+EObeNxopl73YldsrdhZUVT5iXrPhw6n3IA0FuFcbXgbb3EqYHIJAfB4b9
0kB6xVF68nH2RCx2KqItTr1ZO2N1pwhFGS3whuKhIonDEiN49EvtcXlHFTZ6SLju
5qAVlpFo6sr3qtUhEOvvP7f286uBTYk2wSILVj2tiRmuG9OBmj6fJSxivE5wHqXd
tUFugrivx5rdkzWKsOFzl6kFsegM7hX0U80c2qHSsxW7qY9E6hnppAZLVHoiIXhq
+D5fdjBqHYDluei/8qrWDwEYpJWK6Jr+oya4l40mKOElJ+OzeJFI6GGDjkYFhHYE
nKwewZNQIwC4xyi03Z2YUbY4AjZ1LwHMbRvkTIWVMWpXJDNslq1VczaKxIVuqHHI
NRU/LqNTB6oR9QjvjAmWKOZLzS9JPEJ8CNfb26M+w2M4s3hexKmk5zMrXDijE5cv
O3ssFd2sORyel8azLiGHTgRK0ADBOboDXQqCfH2u5T/fL78o0v1pqEUzHSOrXLiQ
UjvylbPYy6tWrY6W+WzeG8phMZpaPwwCT9OAu6D0OVy4FbB+QT6BHOY9cawrf2cA
+CUABRajNH7WmmrCl/X2LVELkvcEGF1FJ/KnQKosfWOsOPcSevDIrLzwMntMevEq
wxBvxYtwxUeA55vdedknB6GvWX5A77xJY9uLCEXQAljLLTaepCCM9gwgHogS0FOs
36uJV7FiA9ZzKfmD8CLtOLZ3BnqjDjZlCyzOT/y5i8IoIsKk0DQ/DiuTf321mXQk
VQlj1nwhXeFsDMhfa3Va56bPF7JGQKW9yAl3prvZmkVLpgRa+zNAYPe5G3IPkAw+
9Xvvvi6vYbLyHuVAktKRXqt9wL2zyo9xZLqATWoQt1Dp4FWyWGpsytxYhjlFElhc
sOiBfeRWeUn5JEXgiygIRSrQjENLma3F2Syn3Rj9IX1w1gKX4Xj0rDNBTyTSnSJz
kLRcxaj12KJImCG+OyLgiBGzhQzZ8dgTEVKeJJh7dfgLFjrfA4gLY+bcoqgqNP/X
+Znmo4sfCgXW2HTpb8fmD9lZFMmjl6CIpnuZU8aC/Mrv8NHbbPf4Cz0pGAK/ygRq
Jjt7V1u1glrb9VsenGZnAeSj85LVSSYi5QTzas02wcW0lpXbgsXdB/kSjyOLeL2c
py+LGrCtXeqpvSwuFDFVHOJ+FRI7rpnkqfH53yA8RusEDD3+Igp6/6LunBM2jcli
bpFYe0wC+4rntDyno+mFQmjVf8X8WPnG0YnRr65LVncjB0vj51uHJFgPihSUrTbc
iKgGCW5T0Ggd0u5rK1poqN+oSnLy5Yoti030O+k5INZlMdRo2cUY1OKvuLdEQQfX
8p9l3exZbNgJBKWAhTq0SKSGh08BTyCXXVEJBA0IQjZF6VYevA19uwT5YwwQwtuM
tU+D351VOatCzLKSxbfZnoRNozrDFgm94/ZrRr5Obkzkeycw8Nvej4YuGUsTPtI1
pM/WpIAD5piVFtxGbt6pyqeBxzE+y50/21RGIEIm7VjvS1LECF30in7THQtTkJVE
neMPCrXad59aR0WW9bhMmpRFvabG0P4mDcPhuVlOopngzVKPwKy0TQHy58wwCoXR
f+obNHhNgtcdZxpN9/5XzWFUql05cYDCnk/K9MiqwbDAoi8FCouL8xSjNfkK7UtI
cCQfVxVZwXuY2m9eqp5IIRinwVdqCg8mY9FoZrGqbZ5PlUjrMwxWiTJcWR5ujGwX
2ZhXpK5pFb2KHuY7j5nIFDhYZdDYsZK5kqsWctzNQeymNyXXDjPlEcXRmeg7L9tH
oqp9z1Rj++HEuxMdXQcTbNK+Frm1YtIrnrDx6vLrazTLeu1uPPznF5rGqMX0uD/7
JitVRX46H+36b1m9njP581mfNnl4kPdtWGGOHEiLNMFuiwT/bvGZHcCCl0crjNGb
KQCliMUxIK0KUpxSYqWJZx1c9i64jrwKbW0oRm1XAV6QfmX4wsSo/0W5AW7noRku
SQ6zERAyCJbQry3bzYviZKN7Z5nx6vErOaWnPyk4DEAUFUU/Tn86orwfuvpZGuHb
M2JTGgaCTEtBE8yfSh1MGmt1n5FUfe62qEAN14WQPIJhpkbwTeL2tNndHf9Uez6M
j25337081MoR+Smriy0XWGoPcXINeSK78LmZyyxi20+36fzJ6vdlN0lY7pmJy9xu
STEuaeydZniLkWXHiG9FwTMagzsWqfQZC4oDxK4IyLsdKEFlGV0cQBncR0o2RG1f
9ffhcngz1szHxHekJUsqMo1TMMgYJCmMkS1ShG41WPJ86+E5sYuyUdil/8dxnVCK
ErOz1tKRUVpVehaZvmNO/x+DrmIaGrovYv4Vh7YNLH2yzkmq7LKdm2fUzwNvC0/J
HTcTCLFT/xpnLjN2hGzu7RMqZyQQVfDkFh2e1mT26VW0scsbOdN8rCu8d/Oa205n
zGtuzGAmXFKG4aOIu7mjK91Hca8vb4SxCZNaP3bTC/vPyJ/rJLsLJiENruWks9qg
HD8chCKk2kq5gw6l6wrC1QCdhpXtolSF5NttJu6smWdMkc0JubWGsHPIQKPu95WT
A4BhZeo46y18DGTbwm39zncayVSBUO4VtMQHKmRY0BtTPnZs5xvupY2zqNw3ZOvw
ivgCPZtzZUj4UspS8efX2OyPuPw0PFhGTej1062tq8PdngtcbBR53iuWoStcQ9uv
UtRPOPXrZOdzrmZuOS6owWTWBlPxIPRPbfTkHBNHf7OiG3Zbh9GzjIlfMugV0kIK
3Cl/fkgzXammoN67E2G8HEZ92r+7cYdZ+9FlZRGZ3tOsxVb/xg28/2eaHmd46ZTd
QKWmv+8It40EOt/4kRdMUoq3TOAZhwfN13GuXwdSGWBHh1gqCLb2EphRE/uf9UkT
S/HUS/eylq0tZdNvMGM++dO8Bdv1VbK6aMwHEtHKKMFIhjs4hpg0SF0Q0QTGB1Hx
8lBOv2ERiOBULR4thbrSYnYl6aIz92yk1Ank9+HvnoxCKhw2DF4tipk2KsjL59tz
oc6uKKodtu9H0noHnfjCzb052VbEQLLAS6PI1etxuXc0ryPFOuqylXXBhcMYFXQU
P73FuCO09OgxzjGBRYqeROeff4gmBjc2Jv0ziu/ShI4SlwM9pI9jSvHpVdT3asqF
RNBQ5mkDch2TrT8ug1BBadDxAJ9nVKN1eKhwFI+KsJAqGFU/xVII3ivoLCWOpCut
7rQRxZnt/5zGtpS+RztK03kM4zv+WnErhs2FtxX8Fg8R0zQft3de+w6HF4DFdqj7
2BJaX1dco9GmiS9stjWdwc0/W9HBqHz0JSzcPc8MGlcyGUgwNGS1uBkItNNt3FeR
WPzrowu6jo6dcj0B7e0HjXYYaIPH8GTJvznYmqbFoby7sVWNYnLUV3ZB7pyvA9kV
gGIZp9KuFqXlwaMZgibQJ/FYZDhSw2/sFAvD6byeMkmF02XSlArN5J3Uxsl/onO3
Qzy5eNWnE9TFhJEX9OVS4eXB9rWJYdGfkRoGMy6KhirjHMeFoNtUBPZB23udtrOJ
kKfe5AgxHLo72QtSIu+vHLDFjuiz+smgNGPEWywQaN8jG95B2H21PBb5ShIL2V8D
bHWhynj+odKUhbZN8l/IEghzzh7N9BMDGnBkdf0UevdqUjPrsN4NmAMQ1Ztbjem+
lbfNu+dL32xTaK1uPKBCCoSuFfTC4S73WnopTqLY7xE7gjhoKg0E9BgatH65s0ZD
Uu9lki8JYHs5KJC/9jXMdiZhNwECEHoyJ8uI+YhytILO7sihjVGl6YILQ6RXc36P
+CkPe5wSDLIHx0DMNagZESxznP4hzUL7l0dgvAWBs3gAdq6QgfrBQpFqd+Km8lnj
gIZv+zG+NPV4Ap+/60pbFR16PaFHsqoAG3uYE+knAVhhUuoD1jPM1BIYDKI9TCnH
bV9xfS5Y1YqA8QD09UmvK1XVjoPEsUJ/31FsVFSoINPuxmxkNvCweYm6DVSzeZX/
rpN7rF5CvzrTlkdFPj7eOLwnOHwp3AVu/7SNgFEZEW9EX0xiWAS0Ak9dIR4IJ/aj
gog13iewxKcIpe+OzbbCus29iIe6NemdKVCm0ErieYKE+ybkoSUo5LZY4L89iXvu
snLHewQrRn1/C91RAmC/5us+q7NIw1Au7aNi31dloVFT5qj9cMa6WCOlRsk6Ce55
WwW11w1ZqbB0h61uhju4zB7MVbe/VU5bqsDBP6pGakvGtLKBPSyAQGYeceomIBHv
yc0Trfga1MxnWBHvDJ2DoO59bvDMJ5eBD9Wurrg/NAm5DIHYojskixkcHSwYwc7K
uoHKNunUT4xhCEURQGL6kzAyOXF0qHshm+Ec77LjCBCpiND8UH25sqkNcFZtcyjT
9zF02U7IoFeEfFpXZWsroGTxs1jjEjQap2lzNCTQb60krfDItTS1FvKyFkFTkBab
e3oYD47mQp4Z7weXQvLcRH/ALdm0xB9WEhk0foliP6f6PQ1nt61d5DhZ29FnTSSV
VEc3vmJcQxxWz6ok6ghVcQwKmAdW0Z/ryzJ0tX47y3n2ZyKFmqPpYCvliPCsjqWz
BniNIUTfmultMbHJQB+v2IsFCrdvMatHXoUnsuLS2ELWt0wxY/dhIJ+eoDCFVQDx
hCHxKSjtaHd6crRrvaUyZzuKMLnXF+LJB9nzC3zGO8pmTN8T/bmRzrgtbBm52g1x
GQhujB5GdoRTrs06pOkBRYTDax85ZuZOpyOwkZSaVBasQ+2rGRLnAw6BWO0rId+S
CiRgddCeMkLx7m/kIkog12u8hIRA3GLF8UrSvicaxQwmwrFeq0kGQ5jhOUPCcFUK
+ks0sPLzu3xU9sBtHfkxAKkxYRQjC2pd79lZV6VwkrLPYK1q2ytLj0W9oLMavqPq
4lJj6ygUvS3++fKySlIF6b+Jx7YXxBWimFzlCuXA/hTzw+axkiIeC49gmI5X45OP
mvfJARwCFuFK+s8kP/kulgRv9yY6b0GWHpzuH9lNgcoqMceeekdnqDGl9ux5Aqdz
RnZ1b26VpcrYDcBsxi8N7sEK+0OuDCCF+kzKx4Amdxxtnbw07AThZ8wDCH1fyTHX
XXypvj7o+tsUTwHIwxdAQ1EQaRRFFM/EsPFuN+fDFuXJsxkiuyJFHKnCI3bDioR5
vgZX09UoZ2gYCMnktRIfHpbVq1AGlBm2rKzxEuEi9fhI2sn+v4bdna+OUcL0LwCv
jXMFM6SQe/RrMAEK3a9OM/w4k9popE1W03+LjQfA8bsdqaFZfVLDxlk5+xJCpWu1
f/Q7Xqu1REpQZHrMyXTr7uUksGApkG+VRWS6YDr7TAhg4nIt5y2z4Z+z2eX0B6sg
1YE2DS0jnreBDLJrDogtLeGp8KCap9RJO/kwpXUuCsytIMLBAYW0cRBFBWZfNKi+
pWM+4goeyj1zAewuqQDDyhTQ6dLK4Cd8k3PMK0y4NFGp74RrLSdlwxDl3zw8Gky7
IoMdleS1TlUpnk+kfcaUhoSZeSWR6K0NGN6x8Tr7dya/yLTOpIBWsWH8/WH/axBi
snNmB7csYJfKakiDIisLxxrav6fHW8EwT0Lw8EVosXvAEspCXYq9gQB4a//OPDMp
7K3oiGFqjQmRzS/buo5Kd2mIwHm4nDKSjUJRWyajo7eA7QjVP9DjUh9SezaL9Bnh
wj57Slnyt6Zx5EgaZnZgyzfkr/6T8ldU1zrNAkwFdzbAxthvFwI+T0TFtP4Le97i
HMJCJYCstZibVyLU3V07BuGv8wLHbFenrryXogKWQbFwcSxS7Jq+kB3TJ3AkQB+b
++9LBt71z5WBNETT1x2XkY8tEFr71hglxmGQKnA1LMDksVfskVDuvdPeGf+IHkmP
+6YhVzetUnVznKYaB8dTLs7Gn5iehzvo4soxH/ic6Z5KQwR8WX5YlmT/Cz4pYQ8n
nUjzqbs9mVP5yfv4CCMkmSxE2UnieSX5HmdGlytjfKMZjmUidijYuXZyxzkw9lW9
TXqY9TeF92cpNqMtIXoFEZY1ncmegRQSXp0+hnxsUQfy5hLeiZ+9aAK8Ti27tfjK
v8ZaPq2ypsKQp7hvyfbUYrcgqpHte/lVmc769kO8OnF4eL6WMIgbWArHTbIncdvC
pofFEw6yQ/bZJuX7YZ5iA/9I+Bpr35QA/YUrU5VV+QkeXNa5VRYVTAWJN11aURt+
AoQIM6OdI+jhJwoYkNcx2jdiN+QFufSLBhSIoY6Sqk5mCyHMxaGa6ZqumCV15MOF
wyb317ZR70bKzFBhXwOcLjVpBl5i4PLpH04SvqwxFxF+wGS7oQWWxMXSCCjukzp0
mIS0YHUgAEW9MY7yDJGiEjTAP7vK2KayisBo9rsSNF19AKPGSeHA1jkXwsmdY+cC
gRY2qfcqcanKBYdl/dTPWyBAvKYGoim7pfqxQbmOYVkcmIFYtdKE3BooXqhhy0Nh
qrU+/XXScXzM4/DNWhvk65MmgkC+eP/jmJm2UMk47qS+OTx++C0p28SNVOMDPN6t
fT63cMQyxdeeN+NOnZVbHZG5JBRGOjfXZ61DaBhux80eW8fF7eitGbSRigdBp7a/
ubr/Dh74U9rIWtwNKOEZ6f0hKzn+ZYzFl0k1mzj52yj3ffVxhCO4WwjGbaYrLE6e
ig5Y0z9+2Bzn0TICjQvZKNHdHVYKZA7T3z4B9AdbTr2GnJraSv45WCFUFi9hAe2i
PXY1VZCWJrZvIb7rldFuOG9nQAH3eax/24TyDM8xpsiO308Vo/C3fpkx2ka3Vs4r
p7F132z7G2YNGLCceU5Wbq1uqPTelXOQJ4n8izCbTE456bI6x+b3Z/KtdTduzjHU
Agf4YP2XLAotuXyDFRX5no3piPqSpF4Rpj1d0f9khh98bMxB8SeH17cT1D8Qqldz
hN/p9Hthv5TYQVHX+f58K0926u9gTFfAVt6v7aq+0cNekWzIqYIRjAmO5oW75IvY
Qtn6QTxb1F4K00YKMvD3a9I6XVIVzB4xh+K7wtstjqRiaqGLwIvdP0K4OVg56Vqt
3NIR4+00nqRz0GY/Mzs1q5Dziexk+CyLn7UqZ2NZqHWCrujvGzvycM5xJA0l2M/u
EWCYhz1HVWXhS8a6WkApHwPuCcszmPXnhu4r3LHNed6Rt9PBHVOAjtBZSnACXnoO
bzjjkIyciMdvUPJfUHI85kbQA/vqOseZ1zWOtvsfO8DYgzC7XnhrGr8WkzFS0nu+
G9AaLoxujitR5RWGrdSj4M+MVVQiiLDy/e3H+ym4NK9sNnR8U/pWzH7aiJvJpx8C
0UjqND/DOuoUIHcbBHjRkuM3sv4MPp/nBRodHEVhfe7tysJzwARBsLp2zauM+c0C
7xv2HL4zroFjX+mqpufG6TAdMqIYncbSaukn8Ijgx8m5qEWqjge2YZzrrecAV/Bm
+kFf38QHe8ZQUHY0xdN37uq5ibA/W9l+kNTsk1oM1+hq2WciCoOZ6j/GkcoOjgKQ
kpE85RVppIPk1e8aDEkNuBk5z6dKkR0lABZweSmyI10mL00I4q46KO/4mH79WiGP
yHyAk1vKsklLJIWWLzZMCK7jA7tKVpMVxfZkcM9Hx7fVFAuxqgHsxRFwCcIkG/yV
vIVLTDJVoqY0eVTeXX1jyVg1jw5wl0NiyNjLMDsXx/FJTTpNGQJ23S3YBrR4Lh4b
5l6LgIYDROsgGJ4NFuF7+3v9d2MxOuI+y2scrMZNutA8ocExV9uUnwSbE3WXG7lU
hTZ5PoHMwB96+8RG6i9CFjR+lQqApOjOs6T63W9uBA/CfTeOYr8HaPy4fCkE0F1e
RckNoHBIF3Oa7arTMoRF2acDnRaDOrXdoOno75gbGF+TACsinb16N/VWRg6tYF9H
8eItSdZpnD0Asg4LGU6MLcwailGw4SOdpehhZnpWnSZAZRYutoT5B9bHeN+BmvrN
wtufn+MdY7iPj+WgV49TOKFxIHJmvB88E7T0S+hsclLT39s8PS7QBt20ukZfTCls
zZx+xURsZzGk9RZeowmoCwOceTAi+RhfvxLcslWWGbEvQJtQpcjnz+RdGjMLt1td
LASqdpuCWg8m7djKaxHwxxZApeJxrtR42MXHDSAb2Ht9mStpuxhjHszetdWr41TK
bXlPpdscee3dMcBRl43Fk2E1BdeUQVPwki+tbhzno08PM8jGlJtq8i1txCBXwcuy
E0R/Ey2MmO7khDob3OjaHLV2d+kyUSl1BsPX2gpilCVBp7AFYAjtutgZtxCIx9an
YUFhCOxAy8ieglXKRupQD7Euh6C8dAE6CBuso2WzgTuveBhtRUq/LNJMW3XlyoCW
qFEDD2do9fxgxNrUDOgnrPgxJPCyZ1YP+vIQc3bY4nqQKmokEcFqqTeIoZHkS0re
8nqpIABEOEi7H0KJPscwT+rUN6+L8BWoIK6v0reTx4g5bhi3mQTnqVwGrk02F46S
gFCArx/Y3V/IOOosGA1soW1VFwjK0A7w4xPBjmFq9IkiO6b1UwNOhfNPaQuz3Acc
/Gg6x3X78iX1dFoUJkpYaDXTAynnhdDCxYn+lrxHxOU4sXc7JNm2IiX2z3D3Fdou
kRHbXC8y+W2giDgngvL2ku3ZP7KHGJ0Ul5/0MboArCiXqJ7UwPiBEJdymrmGJjal
OsJqOvsw/5PVjr2JvPNi0tFXd+2HmnC+fgE8iK1iIj9GAlqiyR9COxInnIedvH66
d4/DSq8QRK+PIrCy3KZdfaqILS8fv6QXpe+G0BtzT19QJaY5938xA3K7hR2Qmyor
Mnt5M2mcBJARZ5rGhGB2pJ6D6SAuHOC0fSW11SwP/5fwovANy8oA2oYTGXkQcjOZ
jP/ELmvgvLQIrQeimDoagGi1ZIIAEYHhekJlbPMptfF+hxVryNfGkZAOmMjPGVIG
sufklYqdNDsV/Frm2+1HzwE2kHjt/VramyzEUvScQyvYx4L90fDF9lslKVI9L+3L
7LLcBvdpeREUwnOkhRhEO07MsQF7b6vhYxd6gH6zbtTaH8L00LtKVqtcKMQOhmMO
JZNPhzDChEQhd+uO+L5yiYzaSUstS/md7TPoKyjhSadhUqHL3YFfusOxe9qOa02P
K8YNW9uRqjS0EbTVnhGegscIrTN2l2oSYBH2JurllaQH94BkAQdpic4s404HGE49
3PlrdXPl9+ptqmBywCH9/kFSkZOHQg9SFiJz8w682y826Ciy6tDcEhCJR+ldyuGW
//NWVqHRrM3+UeKqDj34UoG4FBMfva5FDwuKZ1YUyqfqJuLLdTkhFuBHrV/DEwy8
WkbPWjkyV0URX60y0K6wr61/AzaVzBCuDzMzzM2dD6/HOy0qC0U2OUDuUCn2KMgd
9ByEGm5YRAZzYKmWrofVy252JHNo3Mgy0NOXoPvd8HoJoGyVOOCF2U/OiKaSensE
+9b8KnpzZls6xzJtZP8jjDIpP6reXhKiFXZAeZhU5mt0vW3TyBTxyjPg6Urmu8oL
1X1F60ina2fdVtgs1lKhWrKq4kJnQuAkewQXGv8HNzYkZhPmaywGl18nfAtSCn1r
vBPxo33LQEgSHmJZJslnRDQMlcUeYL5KR6wLdpcf0OeI4ZV41QpnLsMqpeIhJ2Kb
xDO84JQoZdMEOYY6YLZeYgysnp8urwhZLcufA1sa8HeGbrObNhiLNjKPyWmXeCT6
sfs4DnYFe46zZQ0xSNkgRe8gCdfXcOPJTlSUVBLW1l6V8nQ2RRKfndbIA89Dq4d4
rfEcI3IIWFY8OZL0UhT09Uelc/2e/TltpZkwFnJQYpef6bTEohc/s4Ea+lbv3+JE
OP/AVeM1g0GLe97C+PhkeJY9DPslDHNLH6D9vqMhGFxfgw52ZWLgDV7OH9GPejiU
C5LkoDEyVQecmfu8/VmMOVR8SxWdvWKJdBzKu5Y5xy8hcmM3o4q9xJSI8lL0W8f7
c7oC4Qf85giRWrzzn2fJx40m+FjZEva7BhsI75WyoCVCpeF9+0Z9ULge80lNv3rs
jWTTLVqCT13k4loAuTEQtFZqjD2KU4ftaiSU18gpXuL9JR+JpLCKuohVmEXyAOBX
8q65wJ/kW/oLKa98Z7b7gKQdmIJaHjyyJlFb2JAeYrYM84RQSbuTfta8H8n/NUU1
e7MPZAw7pf7KTUCvQUtDL7ePDlD4cRVISWSLEtF2PiLPSX3q0xFEiqh4POxDXRoQ
PG78VWltxXDtytmTwoM4gR96GzbEk4hZuEwBZ4vO9ZCPhMQRVImLfYdK5ms9BdWx
RoAww6prkOc9fhJNN3EKV1LMWzWpNgmA2HjeKT6RPg39GFmoD+9bKO40UjPaKdk5
ys7X93vNV7h0UKMGHSZl6l+2tcNvET5h6VdkZ20FDr/BYI6SQFzARk146sTlbKrs
ckNwrNtgGoGBalkcIhSXqqKgWx81lhZJPgMwlVGZXIo+KfMi2SOJ/cWrQsxbII8E
ulvC71XgKzwcKXyr3vqAFBWqttR5Qxp100giAZNbytQ+muAKtSX374IcknMA9BJY
/XsXNRq86Ov+8yzRSACTpQ==
//pragma protect end_data_block
//pragma protect digest_block
ViMZ8tSb2U79D5ovJNkh3SSZ7EM=
//pragma protect end_digest_block
//pragma protect end_protected

`endif //GUARD_SVT_AHB_TLM_GP_SEQUENCE_COLLECTION_SV
