
`ifndef GUARD_SVT_AHB_SLAVE_PASSIVE_COMMON_SV
`define GUARD_SVT_AHB_SLAVE_PASSIVE_COMMON_SV

/** @cond PRIVATE */
/**
 * Defines the AHB slave active common code, implemented as a shell assistant
 * which basically just converts requests into VIP Model requests.
 */
class svt_ahb_slave_passive_common#(type MONITOR_MP = virtual svt_ahb_slave_if.svt_ahb_monitor_modport,
                                    type DEBUG_MP = virtual svt_ahb_slave_if.svt_ahb_debug_modport)
  extends svt_ahb_slave_common#(MONITOR_MP, DEBUG_MP);

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************
  //vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
YZaeoFh36OF21BovYfGaDv1G1pw9ADMuc3mgEA+lTks5Mi0rHeF/kvIHHwff8rdx
rxef+L+/inhqdh7ZWitYcRlmyUE4br1a+VIDi5zolTMjihtkp3eie4IuoO9eNux2
sxpjVKMYafAx0vQeeK+8BAd/X9ExiWeD2QksXUgxehA=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 253       )
WNM28dMIp611N/hK9bR49MVK8CYYtwKGvU7hq+Vwi69aFylA8iH/+PaFTc1qvBME
XB3UeyxxzhUhnLGDnptRKIsTd5FnBbAE18Nld3WO/eW5VukYeX1IBcE5EnXZyjSb
ROsn5TBEEVYQDKFwHiqqq4LIe+u+4Qj0dBtdoINP/wGyZo6Zkndfksk/owKYmOo7
qoMyHSyfW7f65UwnowvgodsI8J/uUB7kEHNTPaJk6ayF/0gZ5TGj+XVuCeZ/cjss
NudHGWL2sylcncR9W90HAo0FYhYANKB4Sivmr8twjE8MzoSoCFS/9Z+nNnCAYpXe
MEuvmHwtXcheC9Ni9DTo4A==
`pragma protect end_protected
  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // protected Data Properties
  // ****************************************************************************
  
  // ****************************************************************************
  // EVENTS 
  // ****************************************************************************

  /** Event that is triggered after every sample. Other processes synchronize with
    * this event to ensure that all signals are sampled. Note that if a reset is in
    * progress, the reset_received event is triggered prior to this event. This will
    * ensure that processes that are synchronized with this event will be terminated
    * at reset.
    */
  protected event is_sampled;

  // ****************************************************************************
  // SEMAPHORES
  // ****************************************************************************


  
  // ****************************************************************************
  // TIMERS 
  // ****************************************************************************


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param monitor transactor instance
   */
  extern function new (svt_ahb_slave_configuration cfg, svt_ahb_slave_monitor monitor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (svt_ahb_slave_configuration cfg, `SVT_XVM(report_object) reporter);
`endif
 
  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the signals which the slave drives to complete a request */
  extern virtual task sample_passive_common_phase_signals();

  /** This method runs forever to check that an active transaction with trans_type
   *  IDLE/BUSY receives zero wait cycle okay response.
   */
  extern virtual task perform_zero_wait_cycle_okay_check();

  /** This method runs forever and performs hsplit related checks.
   */
  extern virtual task perform_hsplit_related_checks();
  
  /** Update the component when reset is applied. */
  extern virtual task update_on_reset();  
  // ****************************************************************************
  // Configuration Methods
  // ****************************************************************************
     
  //----------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);
  
endclass
/** @endcond */
//----------------------------------------------------------------------------

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
iCbFawE0L0JkNsMR0ti+LHREmRHuoskL+5cMDU7kPAqgzX7TH+B6B1u8oloVHwPG
8SUyDAAOhD26gbaZ+KREkYPXM3kQb5RKgY2GU3cY/Quvrv98YyjakOZzJqfzZ1kX
8OlnDfpF7fKKAZzJrEKtKYDhi9p6rtDTdE9y22rAZfQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1059      )
Uymahc/lVvjbyuMavo7DSMObJ8oBSwGnhGuSoR22DAjkW55MHJjgeHRhjOOcSdZL
C9vIKt667BqvQCrB6VVLiZPwl+ONLBTX9SsKw9pxAWMah3RwtQYwhC2dRZhNjYf2
SpTS3WCzmR1lHqDdS8Fw/EoPI5yWb+EImwWBDrl0i0PrVxNqQkoASlhFVbwysDwH
htkNvI6Q8uNJ2dDxYJui6EcQtBEMbAW61gi0NRKWpntZ9FYx7s+xgo8fq8cTA8zP
R5DQQSko8PxRFd0zXFeVff9tH2PCmLYUPT3oWaPafMzB+AqsSmRamw4W2HeqHUV5
dvMnre/vOSrdb4jFJaDYkM7ejlQssrdydlOgrWcrCfjGhGcIMtQL975OZ2XO/3se
6i2n6Bdj5t948ZKGC/mBqrdZXLD4kusDQDKLEhXmi+UIlSNqYMKE7vLgWctelOx2
WEehkcl39Fa688h0VQmSzZBWax90hVmwc5SJhKo+CDTZffaPaspGvxfXsBsBN6PO
02DG7iPj4aQ1A7JGP821mNvKI/zOjqK51Nx/ZY57gka/Kdi2JWB/RwZin0OFJU6W
kmzW3JVqp/ooKKcFT0njdyUYINsrGojm/ffx3uSDbwpqYMBgiZNPmKN5LtIQUvtP
z6dp7BDutAuyv6OKzZJuwdve9PYAs2hAMUDcixiHjKF3vJ/AFOUWIDJsBD1fLRX/
HqjZZnr1KIYJQAEajrEQZb9s1X24QtVI7kWlvn2BR4j+rSDfXeLyVR788fiyLhzC
1qyBGCy+O8Dzn3Gj4sCQGI6klbChUdEbuqHE/QiYw+04Py2q1XnEBLl5rnDhRYeK
XEGgSnX9P3YURPOcLKL2Img8Dn9bZ6rDDFUd6e9K3pVZCrenm7d+VGxLYeX4r8C1
GZzpmfxuYsobWJEkiYX3a1UbToA+sebzgsNQujpjfzhfsg62bZzv5D/rBZSGpPdS
9b3It2r86gX4dW1rYyXuHtIrepuwGum62ky9uj9ViEcX0WB2R7vtlvNyLgXHJJNu
AzTDo0iNduU7oUZAlX2hxuL3OLOocFAmv3XNNjflSi0M5fYDpRKDvf5wnhDiDco7
`pragma protect end_protected  

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Ox+wuDxKiQCl5qCDoelh79qX+QoTl3Jxdh4qS/xBueUnH3s4rG6HIScRZDNgpV06
h+o4zwMKSCKgXEqP6uN9CPYcb761fjDvHH//yxCzSrpQymFHDG/o1k12iQZLuZMk
up0yY281aoSOx9lxtRRVq5FQStwwtLhst7qxw1zsXfw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 2702      )
m03gm1Be3Cavi4gKOoP+A4VwmDEQiWOedsi21OenZGn4FDYQOOxilIKT2CJtOTeW
llO5sQZQWg0cvK1+18QfKcs9nh10VvINlQ6OLdP8TuAS4fZfuvf1PJjUtBnR3LfW
0f/OI0mVKrl0bPX58ZeMhMaeGrYsiOpRSZkX7MfPtv/+FuYN5zWOsgKtN2LKGDHj
RnL+03DvvaV6Bewu2QaQnsSLOIFRlMIHEZYLlzXyKGqecna3Syysnzgo3vm/w/GJ
D4ucLZ+HmSk49yw+yBwyrqwGppPL9NU7a3xj9PDVdogF+Gs3Tb0/ikxrW9f3N+7/
CzDfdTYTsmREt/UUn/gzq0nfO0nNigJoLILX7XCyVryTnl24FqPFTJ3CzmCc+h4B
k0Tvjcy3V3/HT/qhR75/lGeoaSx+6z27fFOnE/Y5OjPDVoQo18AR0osTN9mqYjKo
7AtWB4MP1E6vZJEDYrZZzOJDAAAIZP+CpuZdiGqOIeyet+8yBFW9vmLKnPakyOmh
cs5VNPtfwC/CPqG6Wuru7Y7dDVY48nSjS9hFPp+S71uQLcgkphyL2DhivLQSoBa/
104wO7rgmRuFlalxH805aDGLT9jrS8z11QVab1Ry+iOf1f0+0GWncNAo46tRZ68G
59zkeNz8pm0XJo8hR3NkS6ARbGg9m6iQYP91rJSRnyRs/CYobWwIRnp5S33URfGn
wMdt907SaDVMrViyYdgBWEPBVm/PMPYuzIYNhQxYWVfj35OaYv/J1PsxwfrhGONS
qeIzCToNFYslGkRiejoB6hFnzI/l2aN60O7iT+Oxlo0vLKPwH2aJXVrLyCC5yxxO
QPA/qKlw5JDNZjjL5Om0kcaLR6yVGXIJgw0GkwiM0ejIubg0G/SOy0pj8FFjR424
ELH4OTKEmA4nj4J6x/jETqxgiJnZwNmjvqK9w/wflXg2VwXAi0yxmjNeETwDNwBN
UYmf9iUpnrgiNqlMJY0OkForqBzuOkeQ095xezS/71v6UJ2otIXxFDaCmmAnd5l2
mj3ssUZgcYKoyvevVqOPe8MCMCDOcHAq4zx8VRm5uATeyqAizJ1Vqg+tQNa4CZEI
ngQKTwJYmUvlOWwsz3eoAqkZ+9hPELAlTPJOGx56GupKzRvHVvWNZFGyqtxgrgGd
GpzTjJxmsV5yXvRxexa0afbEg6YAJN2Axy+lavAFcr5K01F0C/78PsOEZto2XNuf
kIFW93wNg/z1hS92HwWawDoUkrcZOuarl11nIslsPNPh+ahwEDpBl8l68/hMTZ28
oHkvvndOq9FnQgKnM25QWOsTcI5IRlLqYFOVjtAWy3e6ZraeIjYKpq9HXBO3EIA5
AuEI72xRgGeq/AUosXwvOQ+16gmepmBNakd9P8+J7LHr1bVo0QlYH5WSNaCGP7JZ
umCUoSs/CIxIj5aOfQc1+BzhSiZzNZZANmjKYTLAi04A/6c1avMYj4QDoUMV+HnA
yE7DuED53PuhOc0m2949N/TjK9WT1Rv/8BH46V8xhUPHUF98a1NWW2z4i+q60/OX
zZNCkleWGeR4/utHCrFiC48ne2N0t4gWpAFjqbptkIcNi38yXaYrLd9wu2ZgPqNV
s69M2CgOWV6rD950hBCzkz+DXEFah/QOtQrqL34O2PqgYPV42BDMsrOazo+OCULP
VSRyQL/VLon9AsnTRMzb28Mph3KoMtgrrnSsNVByntrlUbaZDPHsZ4z39u95ZngF
X4KlHBCKYEZzF2V+IP3+n5mNMN+zc29lp17CMEhjodGrVtuc1+U1OC51bKDrQxPP
mNblxgH2eP6QEs94ln2EfkuvURLthvHlnWNOJPO9FT9UbafTqITMmRP/ARTq54bI
ooqv+lwW6ukEA/Kyn364ncSZVpzT4wBI9u7GuutGtIQXx/8uIZFvY7GHKIhj1FX3
LQuWvDB4yVHVt626FvcWtR45+4WsGy6fIE/kiMyu8bwYiZQ1n6Lok3ZoJA/NDZBg
APDFfylvBdyBGTe//A84sxPxw9ddJ8bIBuSq0DgggM44lP46eIS5SzVNSg14HOyx
hG9cYCqwkGbiqiZ/F401wjKwVhKy9UiEle/aSpvaaMf1f4WjBwBJ1HZGyddDu3ps
Vxi+OCGdOo2vc4UFvMbMS0SPeb5tUKi9ngskyGr8cTF4LzRltanl/I6o/GgXYItL
tN186u6c6nuAJ9BCyvr1yA==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
K3N1+p80dqQJ5eUl9eq8GbvKavbvdzmdmDSIa9NC9EShK1z6qTT6yTS/ZoTOM9qq
tCD9jsWG/d++BY2o89+pjM+a53kdVyyGbeffA03GPVO2yaE4yYm52ZpTVu5rU6Rf
k3Y/Q0GW3R3ugK2FqfX2YtPgCR3XQNcJ6imkewNMlwE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 2980      )
UQ5TXpRqbOBEIYTV+oCkfLhjNVyIf3A1F2jZA1hTLhHfmuONTQSC3J4D23X/+mxu
hd3/8C9onnnEX2gCvyIOdlURwNLRbpvki9R9CVQ03lOpaEL7s6sYicpmSutnITXv
NRxGdt766Uqb/YDD3uAq8HkGpplhZqkHEGOinmhrmN7faz6XHTJjfiT0x8/lBsLJ
6eEbYHvaTQty0Qnmtw9A+7YVgWKfsW1OMguTFKrJf88hrxRN2FmBrsfFO+W6a2Q4
uxE5oxmhOZjujPTrxQMp5g0uylHHwb45dOmCa/n/53kTU3H9bAVIvKIrFMRgm80h
SUPnkEeUP4df/x8HNONt7f8ApWDU9UvFfwOsMRQ8fd9gODiGX49nEvjczYewuBIP
`pragma protect end_protected        
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
WFjsy5/HbsaW3sX23mBw6qsHw8r7aIsVchXkZg6NZ78YU6apca5wlZX5SJX7wvEY
g/SH6V0J6wNgQbeByAM3M0tkcOa5hmzNE45uz9NuJP5CgD0+xhW204FvMtDIL5zn
va0LUxc4MarTkVMrVsSChQdjiWrlav1RVVUi65oSHqI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 7747      )
e68GxyRESltAELqyU56jX1WyZbZUu4Yne0K+84mldfc0C2dLCDj8KBfwbyumNjHK
CWUcrtWIVnL36lNpuIwIbUZGc1khHk/c4EteU6rrmuTDr/dGFiNvjCQUMzjhOwd3
cjWlRbSV/YQmTC1ggdza9I3B4zWS6HzH028qAS9WIRlH++st9MYHe3306v65JLz/
kraDXbLU/t5OgJDA4Cbzsea5g3xdU3TKylww2fI2sqTyvdTrmNuThxqlwv6JbgKy
NXeauPdYUKTZjMLii0pbr5aJAJ47sbbcvJGp2n5MKaynldUIPOodNDH6yprqcMZ5
MD1xz/Q/XYSYxU1jWvZBDeXjzfhO9CN/kjge+3PuUUqVmbELEEnUihq2hmUv2ebi
nS90riHaICGCH+7II7ZgRQPYlyLfptQzFOuKHrFXx2v6KWL3Ee8Kmm3Y+YJPYhON
7OStkgofp0KRDEe2dpHizSbBolvbtzwDDpewnC2XZPi5sd1jgCl57e0/E4a5U/kr
82Nk3k/xTzhTorTR01i7ZwnUI/xGpZ8DLXk0DuPVrhdj5wnNan1wFhZTKVsEiteb
hvduvBzCBleB05x/qBHF2yNA70J9nHlDY00AVSVAyLA6dViJWhfVht9f1ueZwod3
hidZSMoPmtveNOPp6vGFfjnRKMPiWoy0kRmV/WEpzJ5UoCF+EuM5GNf0jhfo8fhY
RLettWgHDYj8yfKvuFfYQkwsY6Apsm+do6WLGy3O57KQbpB9HNezb0ryLHFYj1np
hmVF970OeSnqbwZOqee9BIYJ2jBVw2937tbmG7SREYK8/w1Thh8XO55t+zYF4PzT
Y9RGO1OX8UjHdJihJgj1AjaWrtpWknWl4ANZkdUgerJrGZu1rXNoH6EsNKRnvDIZ
xCCR3Oj/SpbP9twQxreKpgg1AZvke5M3DxaCzv1X/lh/WGDR8mmGFOvZDEhGhs1k
ezCa3Kn3xyrqK9OhY4nJ93/zStVJshi4GzKnQJwLag23p3KwOQek+kQvIAiH8RLh
DvEUAN7CGAVIScaKLVCqFbFQrFH0qzugHlD8/3Hj/MRjgmIxlBOYP5MnqtMeE5v5
TW5LaKkZvFQx6zkMSCNoRoPKXzKEu0x/Mtbd/eNln4ACMcfM68b8HNCnlV3fmVTE
ugJ3n9wLT0f/rCIEw8HD+xYXaPxscCNamuYxai/ISALcHKuPAMkP/e8AmYeaZu28
Fe+eL8MGi7iPITxyFBtv0JrhWkIfHjCdqRmu1TI6jWVYbxKkiEqctGmoWCura/kV
aUQBAYaACt0L25I/Krta8lR3JkjMWcW8ij5uNKlDJOoucw2a6z9kXxy67vKTyE6E
Z/ECY2Y3dJxGoIkS2GNTuoOpX6uKyN0NK5E/DpGFgz3BoL0QVPYjR3A9uFJT/08D
4AGlANhFCEa8f6mly9lw/w2NLpsegaIhx4swl6VTK/umYTNtQc8qKutOV/tU8S2r
8J/6rFieL7zywJbcCNpNsqEXAFa7nbKg+1aGFmBjJzc2iBApyzf9nqlT7ZD8nR3y
1V+HT/LKJuIh0gGIUph+nWKo8OS1SKAz1McZ4RBeO/9Ia1GRpJCmEa0JXwa8bMrS
ckfIlOYqONeS0ShVt1AU1beE3BFT3H5UpgCuXR06HLNgYCTmjzC+PwQPUONT71uJ
nVZdQq8uV8SJFcTC1ddO2XIaiU7O+m2+sTqP21tnRnkCHTkSYWIzREdehHwZyZgk
vIEa0IPb5FRs9wegBrFAlXSnDjcNM99K8v01JoRRaaAV5WkSTAoadEnjZixXj5np
KFbw1Ud+gw2o1cYL010Rawalaudg/3bqMU+f8mqe56SGkUIcWWGjVP8UKrig34nt
NEIp+qnq2a/iXgUV5FSrV21CIVLVUnth66HOTt/rGu90jGK5oMbmwxQ/rJGJZBjT
HARU2IwSVlnlhdXffrXEr/PZeBAOz1JkpwVELlkR9zMLhGesT9rUFYhMDoWRaPVN
ClMMhKLzGzjw1AWofBoUzQ6cC08s5y8GhZZhJX0IXqBdvn8vf3tTQ8f0WJ0bPRua
JsWujKHb7XFrZ0DSTtczMZMTtk2kgWMwNUmt2F9cfsMRVny+b9dqkdEJMyxEH1Pq
2nIzb8AGIGXgvv1mWxhMPNnsZcG+dgRzmf9hiTy3gX7fkx9SVQExC7mA8V/1BnO/
8xMPTopNAHHmXpqTXarAMQ+1cCpQj2Hp6qoy3QS1IYORRCI/7eSRvb06fgqH7dPt
csjqtz6g30ywTBhQhzRbtH89k1sZN7H6ySW/LtSA0O6EHOMndQ8EPBKG7I40FLk8
WyCAxgsnNkHXEBkyPexJc923vy648SrlQEnrGlQWpQO5pVBZ250h2iPCHq78xjsa
18EnscqT/lMDQIYmhgtEZr+XfcmB9DkisOPDACu02AKJbbiow3O4smHUbgw0dX9l
OEtVWx5lSnEGwlUX9cQ9C7vHBK5yIwNyUkiFjZXIgm/D+FXHZ9tdHDkl6DPluGjK
35eIduSjuhk43wpWIP4qyYVGioPfLO84LDAnW6XPKKs+LLh1UhQDgIzk1w9DDscl
Lv5nlcacSwRP+2WSOYHwU9/ZYHod6UocOKMsj77t3f1olkPjiOwwI+owX2oQuauB
W94mzK4SZdzHHHuCk9RJcG8r2A2GyFdBG3z/mcBgdpw9PdcnG+peYAcuPeEXj6xG
/gzOtzniyBFLuyVizQ5ejHxLoMxH6m9XNox6CPb8A3YAaRpfY/TgKJCraqJTQwR6
0ygxBnhFHbk4ZM4Tp6VGdRalgit3mUofwovBAWc/hHoeN7LncenYRihwlpMW1IM6
FtyjrWtqJTxfzMylOg+cXV1Jt5lbD3a0UoBFYjM9n+t/wFn1GnSJH0LamWnknNh6
sxvvuZGcoxsFh/nGdfTMhbklSo/Xu4lQ8DtvAa189YCuVL3PY+jKCZkUiBIBx+QI
paaFE3nsepfsIaZY7KdO7J0+hwoW/Hp+MAt48q/er+ZuiZhp4UGoEGcEE9oZidHk
mPasAENIYh/pLRC/WfRTtP6dGUeX70EgVJVJyoSkHVTCv5FzchXJaeAMZzrj1sTc
CtWT33Y92Vg4NG0ZMDP6t5HHg30q6M5Nemn+eyjWBQh1+cRrFFIPpywTt6Ltpvmr
Q0xYs2qHhOMskuDocU6dEAWgjhgOt+Q9ycU39qBXcDUOeGCsBiprxEzE4tphK3gx
0RG2aDneLCKe1O/TR/YRTZO46YdI0hdItykTm6TD+UloURvdm/9L51sVennVcplB
+wNCIMPvSdL4UMrcLQ+pUcMRuo/rkyN/VGkO6X1m2aCkGqhWTnfsEII7hahRqFbn
cZNpCyQSh+j0VlRRxeGZUFfeZ3ELs2jGDDdEC2jD6L7dph7HgdLigvUvJ+J4vgWj
61OqwZlfThrEz1EdERfYaU/1IEi5/qhgGDzayRFAL1bi3P/r2K6mZELDL7F/Z1ae
bzCSoq+GKa6ui2gW1X/TUmD0dUHNHdDIeUKpbHCMn27eZ17w2YmmCekScKL64X/U
iIsWRuuWI1l3WKDnKsTVV/2iUQ6kC7SHlxnd5Y+CXQmMUHMn4dZhrmjIOuUXmcr5
SFjLEEprANg4IZggEpnwWoA9k2ySW9fBCEU9vPBKCSCr4wK3QyrDej+pJWuUGvUx
Ng+iEhAFezAF/L06oniIAKPE6Vew8G7cmpYmHXnmI7QXIjKkjHnVsS1rG7wfayyz
kN1OVBrBlbkO6579DUELeS2AQUNuocI4Qe6mAhA238HsjGS2mlp9tFY4x2pgbBnU
I+xvGOm8bNpym4W/GMyahYDze9JQwrUywKLLy6m7WNWCuaAvGJXkfQcGws7dFcUs
lHVP2tp2dcqPlRufmHi778fvNRtrk7x1WIYQRPKNis9NqLjsiphSl/jMEV4Lv+pV
nfUVv8jiqjuTkuYeLNInHRThEyerAd0rBNM1zNInfZ3g++LHkK104U6crQEU+83B
4PiujCkXMLk9soubXeR6adQtymfcoK09PqTvY/YAfUdNEN7APAUuciwm9dWcnrOb
4Pkac1/UQ+kN1kqhdBD23K+CmyrBQfdezVn6HL/TJbAOi9qYnFBWjIGWbQ1Rm+2M
b0sB/R2nDy6oI0p40KF1cwrMGQS9DjTISZ8OawxjxZavOX1+juY1B1q9ZfNTS48M
sdiOMUjpdL3/bptomZt0Gw8gqhNcTXqOVPUAXl9MQTQbTBPHZT5iC6ZbBpjH+28y
dhjT2pFr+QkkA6PjmpaIBWsxXM4Fp5KzQHTL14fpwuOfFCPgKcqyIlI5Y5+JgXne
HymZ989QxjKqk5UUqCiw2lmef0QXluD7QAGNgJvYiQWV+R5DbUyJbpQwi6h/QIjP
1/gXfkeoQBTwUb48ABzMxJXaFwRyn/w/rYf1/5zr7yIEltP2Z1MRbSzfmalZwPY3
ipggW7IR0DdxXYKinl/8j9BkX9mUcSHmmjJ/5txVslWqljuU8mw2lyCXqKuDK75B
Aer46Cm3xV0m9T0MfS6tCmYPRNVhLUEiyd2k1mTXfLlcknj0rAZR69qHWSAo8rRd
p8umOvXd03Tf1MywZntiTGvOzs/l6omKiSeDh3NG4KydUimL+x62iPxzGGijx9Nm
Uf8dE3fOOTBDYPoagYRQ+BbFur7AUVVhqVUy/vjeByijlSgch+SC9Y690kbe/VxA
nXvKHa7U/6lsGeLHwt8KMmVHqMBR/4ZWO2J1ja0b6xa4551o2jiTBK7isfRR/wx7
mTDA51uyzRydJUDgKMxfr2aj+q3Rc63cGUaJuqSCn2AxNNP2MorScIDCnruW8fGd
DYTgJx1bPjE+IN0hU/wQwjuVeOjftqw/UeyK2aYYv/XFfTDFtOsPGYbUp7ttkpB+
iLW0pHDAxRiHdwtNWrTyFSYaaiHvaBkQKCugldhkXk8b7zh1M9uxsoHKhZFJsvOg
gVhhdZQJ29GwuNnl3Vj2EK1kJ2d7pos2TP5B5BNzT0+Wf4IADVmuTY7Bj9e6cHTS
WB9tbVWDID4lNvzSVT+mueHdOvetmtikFTkywfTBdWtWs5mWhbq0EMZTgPEfvJOx
s+Xk8FoYji4LLacvRBMhhU39L1UG3d2V9hi/i8ZwxrLpd33iiZA0j9FdUGAREnIK
VvLD+RDVOQnixlrv/AGO32UKNkw2mbNAogdrMVjpUxf9wAIdxqsQr5nlnB3gVFDm
sBPOU/IOO/aSRjQgXOfxwPqsreJxU5q4I3anMGPAmNDS6pTBFQr//aTO7c9LW44p
mEFPfdlg1b7ixeaoidcn3QABk06M0URQwRf2xpbSnm8nGlYxxFgAt8kEADYF9R8c
jgC/mXe7GwpkCHB/3JB0985JXeVHRu9KRudAnvr6zywsZLGBvlIFDZt0Xl/2VSyZ
fW2MtI1KdX6gGca5Bc7uap2bFkrZoMUthNXSnZwPfMMH1gTNdhwVqzgvOA76u9xi
Jc+SIm4OCXJto05a4mOA5oNwl3ptwzeQRrA0PCbO/bg8XcU/m/wALpHw+oQv2uTH
thBEqNVSZ/0QoEO5aKTpZsmyuUxMdvTIGGKLFqvrpfPMGuM2CGSYUrRr14EnsKV5
FqWxhrvoTM3ux9llrTL7N2rS5hZKjoLOHS22yyOoua/OcEYId7SsPo/qwXcBJ8D0
M+3vpNrqSIX29JessRKV3zII+6aC2gRljk089rGNygyEbZsmqvE7H9/UIET9uAXT
Je26Li2uSb2k/yhtdcTW9AL32QH10bpavTCCGR8Kovlhr7jDcgDezNIHwDYXTFuw
vyVKF7DrmiDP+vaEpc55moubvafYgxBS1+bSnmaAVTKX1tesefbDT4oXGLfRmXEW
h4IWd3HJH6QFvD2iJwUT8KIaNCNDp+FUHCkeod7WGUMmvJmp+6G0CgGzuQW25kXG
u/1Dcfdl0kSsNGUMbkCb8TfVcP1THTC97SGqnxb8w1J0gQYBMV821RnNjStt5bSM
rCZF5n6WnjGwg36/GEPX6SYXcFGzOxKvxMe+zDy2U7J89FCKJWrNlOZs03c1e2Tx
Db0ePw61zbBMgOj2M6bijHg7Q1R71MfsebCRCZg1O+5OkCj46QvDm2x3bxrsbjwY
43wxzaBGpWLmryIlJorLozUKffuL5n/9l+6e7gfIF9hJ+fDc/3+o15F//99O+oSo
UdT7PUpVOyx0miSyUbO/GRX3WCnnIWtptAXhZv02NqvCUlvgy5G5zTeOQs/hHoMQ
d4uC2FPFWTKPa3wZZPCCzwXrxxKnHu3TNsewl8fxj8wIozZcfTL99tjvLVHINLkG
0JC4ed5H2gWeJqic+RywJZ2Sek2dC60erLZ+IF5FWs5Lh1eHuIM5iKnhtL8uNmbz
nWr8BFFa4B0lOvTuzgFhIA==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
nFrDJUrznN/FybudGrn+gyAHglt3tFLCvmEs4aPoEsubLbRcyelhrDHlLD9LXmCf
Kn3LwJPzA1WBfoYNP2/etgWulHmY2vAFJcy33ehIS8leaCJTBcO7QogGTZc4Qx8T
Gct5eET3TX401qFTW/k08dA8ihZH/kNLqMitwMPZDmA=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 7866      )
G6389iB2rpTBP9lVxM39DLSgI2xHUwSXEEppLGX3uUtRIC4Qjd5JU+qYnhE47CU4
JrTW7VNfM26ioM6gi+So84Upmi0P6aWu2KeyViKTODTU5+0k/gEEy/6YFdOz+HRk
zIdAQot5wf85cFVYCbJtHBEU57VbSs8bXASq+DkyDJM=
`pragma protect end_protected  
  
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
M8StqxhIzwQFuLuuA9tkziF6KUJm2lVzaF170jQpDe1JrGvPzcMYnchUGOhbcGqo
5qRxj+WnhzrsxT3jUG2BW4Mv/NEyWc8WKrjsJCBNCjNP5Hh8eBnevtVh74KxB4yJ
GTJRrcZ/URQXViLsqF/dk7skzOKZCwIeJbMCBE/Bp0o=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 50621     )
olcK8A94mqOI6hs7vxH46/YCaaEyrxN3HBHj78Wbl6VRHDqKMlPZ8o5Q1THhT3Ki
ESE/jwEliHx6PJvJF2i8n1Ylvw8JwXsxbD7LaURqF6W/sJ/OjPBx9cvhLEwMLaXv
p4SphiZH/6+cpsxL+LTMlQLuk0i6xWwpLpNiNyX1g22xChAVtIBXXmsSevLCDVIr
rK+Xp99N4MwBQtE+wWtVVGOd0WcguDTAtsNe+/LkEoPzMw1S55r5loiFLw6FLJr1
zjXzMtzyz1o77sEW+4xwKFVXq03ownwvxKKioliHruNmwcLMcKuS5VpnFE4vvMd2
K/Zlg/y2OxOUDXm1zlSPb+TsH/cUGnyhsABneK2WkWST5ll2uGm66nMMwSRFDtCr
UUQQDzDLU1hYlWZqvt0luAF2RizheonPTDFUXaY+C9xQCRZ3svr2cIStaKwTZbwl
3SEihIejFvVayL+gAQh/ef2NJHO9IsvEqO7Ox8AsjUFBSiWhhuey+oAJjrB2muAH
iI0AF+dsaXTC6VFJVC6sWYKMxZwInlAZ12rk8hJPnhD5TMqI8WQMXKzhJTBRxMcT
l8am8O3I79DbUTfnslPS7tEXB6DQenL7Q1x/zV8MDkl6qlkG26jD7eP3qnQhKqaX
jCoEVHEvRP2+UdgLme8LM+rEERp6DlCjD4FYAbH2H4UyGLvBXw22FYcqK3iPniHv
iarRXvgsAd0XVyNRBl57/PgeDhZx9fb4UowHXXR+1thpUVTUpfHEj2JX2OFHQlS3
uoLNqZ15bu2bokpO2Q9v5RaS7c/rexL7AG9csWqHdz7HYwCqN6HdbIKVdFIEpq5S
nYwl7stMLrPQlt/p9CKO5vg4ZW6GZJLw0TBGEZaUtt2ddpw6w5xS4teK5PTFKtb6
sFwv0KMlzVSpG60fzLDPYjwWdbKbMXH9ZOxA+lqN/PK9faObdfamBwn8pcX9No6Z
PPyf4G4KwXfxj0NAzyrzPxoyC5NmH7r6xAKVjOtndmxS5Kyq8FfpjncmUf9+OybM
X0F8k9JSheRnR5ADJZHT/g2WRAVnSX7Vg9Zmb4A49V7AJdGjF6HE83ca0XTGX0VT
yymuS+223O27x/F8YUyJTOjHe8BlkumCbgEWfAYBaXyaEluHZZaUT6kGSTLJRKVQ
gPyqB5uaqEL6HlzIPLGoyOpD2/Rq/BvAwWmhWbo1vLhsCcAmfNOuhvX6emgVSK6a
2EUDDR6HJjQ2oTK4lPG5a/2cNTzuEwJ0uaCNoXiVGaphPIf3fdxqXfcAXMzNjtrg
4Zoy+cbJQcaG3/9+ZRoaVzX7wkPzaXh+dxtYsfTbs2TyfcYx1F0OjJYPLINLCOZm
9Vx3xayEcGXy28DLqUc40nznith5XEYCuuYISRTZZe1a/c/CXKIZSW+GPYnYenzm
D+TXDESf6/LN2wXsKNNuCtDNmDS/AZUmWmIJiFf7KO8Mx/pf1+uu6RU0g3rKR0Gv
A0fnsLh093JfC9c+QBqui+K0lqlp26tCRVdcOs7RzBTREcfFJy2V4JEJnGCxcKIx
s68lwUCv5+PhYf8zJB5g/pW0Tv2TBCsDA+FSdKsMQ42tg7ZDYOsFYZkg3uRmf3xm
eL1mC8QGceh9JWLBxOX5ud28sbQkvmdC7K4PUiQL+62knwRB6xzZwdMoFZLycpnw
quD1+IHF0DF9TP3p/LsjwZlmVUH51fN7BwkuneR5C9IQRyMJuXBzdcUxv/rXzd0n
I/z0ku/8c+WJiPrKGdMb6c9j5V+4Uh4gAsxQBz8ySD4AqTTOD5hhws3Kdg47gyzx
8Ni2UNdKeu54ds9Ie7XWTZh7s61hg98QOd5YkzxKdxsuXTsgfjbrRYYiwAC/gq6+
DDD2OtNckOZDF2XhJ0Y/8h+4iSWrNwpv4yYNkjceacGF8k/BTdKw7qL1vqphGg1S
lbps7x9Rxae5Z9fpf3EP/kN4s3J1I9G4YnOS+p6FAY6DZCemNhBznbb5VV03YAEy
nbQquz4/D1+cy6p04ZbnmP2J5mfqkkcmG4QVjuL9T4spxrEHO29EuHDQ40ZT4DPp
6w1xrEZvMDROQRQSte+3btaA2g0PdrqifPvxEnpJ/ELIrqvuZxCaQqWT+eHFrJUR
rmbVNSVnQSrynERvDmoelmwQYoNTDHS60/LpFXQIvm2D2Kjd/QwUTj4qSl7mmfz8
R1l1g7kp9jQ9hpuXlPQsaWvnN4vmvszfEP84BRNZX/vRsm1JEpTPrp661SWPVm1x
5h7oK7OMtt1hF/yAdoQJlJzBID0XUCYvm7GMbbhq8ZgTXmMawMTo/p083l/bGJIm
w4SabWlvCVjj8qRAMx93D3B/9LTmZVUrSsug8aYXt2EWJv1ffJbvNVY240NyL6g5
gm6prJH+XW6d39ZI2R4arMjHr9W36w7k9TK+Yo1z7N9zpWAq9nZTJS15ZGbBLIf+
CvxCKKiZ3j+InA6j2dSev9l1mK2mGcgUB5vDtm8i1qFIy3Q9blSOHLnSTJWdFzts
8PKzaa93smQi7PW+t0zEn3DsQd7iOKuR1IKhuAV82hZCWxNyjCLaSLPvBDsG6BZN
IgmYRqru5BFVnRA+gygQ2jAwB7e4k+4ZLAFl+164MlgsXv30mCu2Awfw9Ur6+qP1
QZ9URmxnKibrpGN2JT3mNJs2/k4KKqlw3yBrM/SJz4dviZ6ukKSDenoEMrFq/hKz
wTqQ8oil+cHw8nfpMH4xtllHp18ttRRQz+bumSZn8uJMi9C1i5qvf92kRTeTthZl
2uiiL+7V6sP5hYvd2g7K/Dn54iHTbNBguZdRAZ46UKdO8MwymJHIZug9qKq9bG/d
AQj2aPmr32jK16nSBHVSTT+xrbUM9+FXQNzEVj4Y12UP2BWOqv7Q5Y3P7ANQBBgW
n8QOEY3pv5eVq7NqrkPsJHHaGWkpe8xt5c0+9DDTu8T/zEOQs8jJgkDCKeqy8JGe
3N//qXgYzvbMlelCggXprqO0G1luwzNjmrgKqaIrZvSBYGZb9ki94N0Oo+w+BPlz
le3WLjN6p2KkJl4gXUTh15/IIrAait+qPbO6r1ajQqfrK2NFq8Iu9jTdr71ZpRQx
krn4wBK9e3MmrNpQR0bWtqaxfMNfSMrokJbneJBB8fcQVDIaXWIt7kq03liFj1si
ccwxL+vW6xujKKffcPvdvItLG0LdFmlb8xhDBFz9yIkcyD+X+UBsmiRbM7gmu6jw
8Y6QV7gCNHktscwTO1NlKEjB8pNiY20HAxzDg8flaiCilkouTFg2k3QkES7vEmke
LDGDlRgIrV+bpCcUFtNYk0LvRDbvu3aPA4gV84zb3XXYaQw9oUKy/oWCE7zlUV9K
BydypwP+beILtQjkI4SSEZtyYjr39RWPoeLcKwbB+sRGVmyla3442gNx6IutTrUl
gnSuwbutyUUjGqlhUx16xiUTAM+pWRG6WX2jC0JRyOm6rF80USQIQymaf9GHspBI
wtrBlx6QCDkaqDlIUYvUz3843YMA/J8k/3pRJwO3pu3qr7XiAq2R6CFsLVWQwnF/
h6F6NfOCjk8Ew1lST4XXw5LBK5ca/4sJ+J9uwXfyYjt7mg1p+nYq1lI/ibYgDYFI
5HNRAHmxuVDgXqaiHJhoL3cYaF3A9BqFDaHxE18DebGbpw4pB3AjUdZHbGUkLu5t
SqdykXVsA91S3254/NzGB2AQXk5MTt9GkuG74XRrpejQOliGRZTIHYnkQkx8zrzq
P4102SvjG0nQEozvEuh/LoSbZmwcOe5MfZ+GShturhZUPxQRP7vagHTCKHN0F8cb
5z4JjvTZVc8m7spnyDSZgagCDiT5nOFTQiTq3DrJryDEMYvMn46M5TN96BV5rTG6
COuxKB2Os+EBocWI5VePM6foPYI9kIuIypkDS2dR09ie1+RstSBCKwwuHTjW2TuO
cSfvn+x2SnKBcGGBH4hTxPm6Ky6T/yCl/NLXMB2TN9HSNgVGLIaQudxeY5utpgDw
gGOqHx9/tQGvFXxXEGFHRB3VwIhxxd+d+WAQE5VJIXpCLvy4jrvfaNuw5Ozl/2HN
tzLYQxVCR+IrQA9JZvS2uhdYBPIa8lWj9qygBT0fv4p9Pt2gEI4GFyG+FwfJRMoq
LIfNbfWd8J+jUWduPt4k8WuNYMaDgYgo0J4B3EVnhfQ6NnjE94quebSBG32cjswd
V4xxhkC63pPklbi+GXPcvr/Z9JoDI/RlEKzIYxdlSojhlGKeQSeND/8XRl6RKBJQ
rrmnYteoqPNdVppkbdqWazUzl9gHIxvEscJN0ZtYzL8NjP2OgVCYWpgcx92bIjnN
Bc2o+5d846imXM0usS+dNMcthQtG1NCGxW6RJa1vVq7ODODM/Wv3R8BRTp2Uiscb
EGZfb0it/Vgn4g1wO09sttqcU51FAI6pi3+TSP/Ne6ZC7Nbj6w8eoIa1MsMkBvqa
iREtTEzxobbnTdK9i6BI+lQ6Vs5rTYelFz0k5X/wa9liKr4P+SItD6XvdW4Crfti
z4xJz4JhfFX5XJPTVLdOr0NB58iLyNbdcyAIfGdnaZ0oKF2+RBKrG29Kt3uTkUsn
NP3ChELkywRASc6Yl8Mp2XgfKw+yLCDR98bf79nv/xD0OlRmx54iIVKyYV3mVJd/
YlW6lbqPzWSfPJyXQqUBhVsM6xw5mKwdyuAkmRl8ihgAA4qxwSdvAfrADQmIIoPR
a5ssYejBgGvWZLxNH05TWiCqcVtkxo63X/zxK7UKMhSjWCMzCwp2nQW4Qk35vRMe
uY+20Ur52zVJJ3PYa8OkvZZoVxrev2ucNorUI8AecM9rGITurSCmOWF0UFdiyvJL
Bx/+VzmSP2xfo80ChFIV2imWlQU/R4Sx6LTJ3P4ecH8rndEms7hauQsOLM447rWj
CwtHNoetsXCuTs6Ju6IwfgaqhJtSwKxx87A6FIclD+ULpxSrMYWCycMDYETqXFtE
KkNRwQR8wMrdiFfkkhkpPYf6TJ6occdx9PVC9u1TXHDcrDySxFBjCAW4qkQCgci7
egneQzLWtxdwkknDjFocm6uE2cBrsrP9tiM21q/+7RzemlEMsl6ZvzF1wlUrZsU0
PoNOhmGE0KjUuIw3CX1wtSzvL71dPmScf5E5E2ZEstZI3zgS+sE7UFtSUFrUbo9m
qXrcp3QP3xHPHzSp2VKBrh/JwZRtbiRqrgo+7IccQCKl6T52xzv7bwjfHZkkuEkS
k9XOvP09FU5V1Nnwt2jmfY9DniOt3g8xLpRW927AiLZRFjTdEIK4xk0PyrJhgZai
A2TnlFevPyJdXLSk21MquMZ/FcZxJyKzAnuK1mLjGxdiR80b7mzEmzhsGxk1nY/1
kyvfc9H0qzE8ToGUZXUs/KvFJ7CvV46/pD1zbyGyOPVeUv/T3SEookxkq7O61+eF
5nPNFvAKAwP+ZdjCIdDq61mkw58a+JIMK2fmYJcqp95go4kxHohNnEp/GnEUDRlK
Gmns8y2/krybF7NBx6hfu2YUAzT+L+0u5glJLotJMqFZgr+tltsFTV98nunxhNuZ
wk2wdDz9GlXhJRD8i/g91hxwBQWktreCy9MTuFrBHjB8rhTg3DXbG90Ss9xvj+/3
KkllqHQYXef5H/mDvxjyPYdxBYhgLB0OY2cPDprAL78k6CBzhBNFlsAGiKsWjR6B
2mfEee2Z5dpsjMGKBKoNd0qesYrmGPTyM+kaAyG9tgljSseY4c5wkkn6rRk0bQZW
8EZms199HexFeOqZ3xFkjEJjqOPB8RFROjUtPVLBTyZ3ldcKF7sbGTcuis4cy3gp
qkwL876oiadn7QkYmL8wXf6Iz5frM8jMXzzGMTyeV9/Lt3BnwVGa41FdeSKDJ9i2
RgXT74lJ67kuL2S/q2D76M3QS3rs5pkkJyxEI7rBSvmFpOpeXTtSivUB66/WomYi
acLTW2l3PwpoLq4FIR763FHi5pfXP5s+ZJe7xwyGhfVYqEdne48X78l+UKNBVE9O
NlcyWhrchUiORG/zfoT//w6hef7GVNTTMN5uf1Y7cbsk6FkuYBiCJA6344XrsZb0
uGRT+zxmc6pxiz+GFQS0/nrIFexdslEVvS4AU78vKvs9SX8i4zJelWfhizj8VhF5
lUFuwm2GE9ITgzkbswxLufPErc/vvGKPmaKuC7ULHwH+znc0N/Kta0Rxq9wRSd6J
37PZGZr7ilZ8WnYUUyAiPTB29NbhWDTTz5bQsr/mB4lewEOkTadoqyGU5zohC6xg
mirVmPD0JgPn8G3DAJoD2yOCJ0Zhb2xiv8ogcGnZ0sxsiweBskI7+QkGY3bH5dyS
/o13IBl2MQvaP7y4RQVaAImdgTFUxtj0EAfKkPvtSWkHcnfZg7+bgM2KioYoX/0/
H0VBhNtQFBmaVpl+z7AIX9Z/kf3RN6kIKd+4MK2RMH085eAfV0+erhQdeLiFwYCd
40vScLGnYcGZffw1sR0W7deIV87+rBimynDYurgRgww3+kOiaKzSM9IypRdSdBHB
EHP3Kgr+e21m/mtI3vfjE2aQ+RzkYUxmU+v47jSmWhuFEs1NpeS3Ec/r4rTNM7v0
dVqvmRaQqNFmnZ20U/kW3vn6fHk5i3TGmnK30r1p7SZzXeJaDVIDhoLhkkQe2/2k
fKPhjRrBwfD85fVp/DHE+TpXtdo7l0bj6T5ViZf/j4zNEoOcXkyad82QPfzhueRa
8WPMw0iBAO9Nrp4rS//n8tZ7/e37gYpa/D1MFgI18Hs17mAdqBW8VZCi3cgGAcCk
BpsgMfkHQNpaJBazZf46qvliwczGox2aT0imGfp/CD975TBVyxRkv0/bMQjv61d4
29cd8wH1IrYX7qnyGlVg2v3C9k4znfvld1vGNImMwvWe9kR9bLBS8fy1DWd6wic0
/730s4BVKOfSBy8dieJOYY+sbiUPYoswBJQEfhL4NCF3oHWwqqo4d9Yog6LmozOt
pL17PdLGaN3TuQF8PveqKwiZyIGhCNIWrg5EtDHrV5JqrKJzNXR43S1PSFqm4e0Y
UYUypIRm+CqeT5HuRLm+LlSUHEbXvif/X6ulVKJnwBrcM7drOa32CnXrl9cjyWQC
QqNhYlfzRNlYVsKkbOpBtSDj6pqM7afJ8Opxh3d/OCd60XdqKFa7agZJtSe7a/at
e4EAz4wlCuxO41TF56uPQNR8vJj9YbBCTgX/j1w2ZGOD1qxJazos+lnOZxIMYxzB
yNhUL9JcTMrFyzXk+TNTDrPq0wRjJIsDU4IGoQEBmNm0jLq8OTR+/dbSdpGJa+sN
8d4kre7fsNuKZoHss68Ot2K/tR9h7ExiuimUAEGkIvyPBNHtB4Z0svGImdHWDl4Y
u9PBlPVkKgdg9y8z716n7WVFJ3bxxlymnEL4137l/gd6H18oeGl91W0AM2aF5rtC
c8GNtapcyyZmxx8lDZv7jq5j4ikAIbOGnxPY9bCuFKGxgac42Ef5dKalE0xKdF3z
mzaHRjmTzNOJuq90rZzFJsABSvsqnNWZTC3+0RTJ/OJ/hr3tBl30MaeSNo+RRNlF
D45M0LkHGfwkWHtFBsVioFqvaVC+r0jQ4DVfVRlVa1veWtG7U+Aq0ODmeCJN/+Mz
PhTGxXta/2LFFjttCX6o7gql17wxwi4i8lAQyHN8YlNE4MDrlpuNt3p69b5VIIsG
0wsMU/cBvSJ5eAoxGxBTxCUBjffu6qfq+5HNTdOXfbfDGLOlmOTEUh+eKyotS+DE
pugHKTf6isLW1Uk+oxBZa2l4JvHLNLCCU2Ta4sQ5MyuHffYWrNQEorOHnHf0ZwKF
7v61HYvag/0ud3zWosbhOBP0vk5S9x04xOGZ8m1PSymduAq9qKrhGTtpagtTczrn
3zN56Kc0bfOXhZeW8Vxqd3xSitBZUD1fXtEqsNEZB9iHHu2rRU24YR4lPoC6+KnO
JicRMDMgfQl0T1z0W9JyloOvPtilA/04FIflST2nfep8vVzJyec37vxQct3MFwIe
Rvk4RV91p8Puhth2USYuNyGUinKMhUgJzr9yp3T/AEntSJ8fPho5t1pmg8t6mio6
7q0za5YJPDwkNiFXvX11iP1+cEJn+9UAjGTyQrpZOrQJq3QMbQXWZQVPqoASgOXr
lv4xQJ4Imp1jtRSo+DAM0cMdLMI8OhTVEeLjzMfdQfCJOJjDq3ncLck3mABcgXFY
2y+JWvnk0FdLQDN2hbVdpp2+Jno+BFqW/s95xEykeAH4/+D7QhzZHJ87w1hOETzm
bxJvi1LyN2hPZBqINcqVybod3H8rx8e1f3dcW8XIlAxYxHM0jcjPD/c+5Z4QqpCQ
QP+t93BovLAo5tNfpgoe5331Na9oYECHcRWdmT+qMHCWzso9dCj0U+z15RtHf+ol
Ia9b+MoW4sEEncfrBDuLK8YWlh+bE87TSq2pzPQg8GxJPWAXLLBfT1jM+fA6WqhX
L5A8WOpmxsSDBSm/1cuDpzJIB/rdjCtK6bcnFeK5ydvudkeMXuaiogAbX3yvaxRv
XKyO+QB5g6FXvxstIOMsfBtK1AdvJepsBy0BdpZITpotxQonVQIfsUWcmBhlEhqp
Zalg/yG7DE+UVdKhF6aADgnbW5ohUGAceqku6fnEvAa7v4omeSlk0CQHana0dxjb
n3Sew5qrmDv00xNO+zILl4CxziFtmcQltAXEmrg87CybQq5OBrkFDVxj4mpvp6C+
hU8VsSgVcI7+Bf69a8UnVqm7l78W0pp06AH5jXJdR2xYIOK0mIz8VtQW2HP34w7L
pN8wXXxMLdirpPXzrKVlUXGDO6nhW8vTLoT739ICMOXnSI0U4GVIrIRViISk2WkG
QApPuAsVnOHzxD28Fau1NamEYRpbmJ3+tyorYBbd80H92f5L+FsI73mPYgYdsrI7
kTywHjWW3ilXw9/S5VZofJsSRbGsUWiIgPma7554U+z3syUVInP069qbjwLnloC7
IqEezvEOmP5TU63rSdIfnRswIrOlVhoDbOopTyKWepzBOf4yuP9gsJJfjB+lTH2y
I1Y6aL57ndf8zHh4Z3hB6XHy38e/shkFTCDMIWC7lEFBmTkz1q8uJrFr7QIAMblq
EOVzU+3T5bj/C2XmiQjO1tVqGby7oUS0UV8gEhPPvLiu/xwEi4F33LgiTgg+eKTv
CG5KCKRz2dX6TW4RHu8I65bLUO78zZ7x5BPrjSxNGlJcXcoeC3KYDd/OGvLflo9a
PewHHlfWk7C3+v+680VivDC01uQ4shyffJHDhVyJvBs6yCks76+NrysDT3HB896d
ZwhedaTb5ZerHIKiImiSGabfqxqMht+qzxVqGiz2b92NAAtedT3Y3ajzYYi9Qpdy
zgX0GMBNr6dhlRXlauqDnHXZlIAtGnsrYmUtOa07/UxahB2xAemuhym/fRpRILsW
YeSyW9tDOLpkaWiQ1EAu4H32mPpQobExm8aeUyjoxFwCQzjWlsbFO8RSZNAO47GM
YgQRvcJ87pEE/tgnCaQD1cJ1xIc5KVqtVgaTuy4IF0D0Fmru60VkQwjtSOk5+WDP
vyOFcSK9M9S7Shio8TqT+vFK9k2vcKWgqZPWLg5zdYe0Jw2HZVnB/mkRbnYg40O4
NH3iS1/YjAt22d6oalTtiW/bJAmBwXiOIKihffZZqa/rBWP8Dg+iPXUtm4Qpdfsy
lACabMtQYqEyOjdudPc8cHXZ9aZ4cdvZg3QvB/PPITUuagGa8OB5avzFVbPZX5uK
GQf07CJ1GY1TEcxF3RHZD/TKCSSF20wr1UH0hkgebcPYC+XbNasQqVL94Mv9JNs3
96+GfFCY3hLIj6gIZS3kiuHqNGFqUuveawjDzJot0nY/QPUC7SB/ELVx5kwnQOtU
l35YRIPHw4qt7ReaUhZYUPJTsE8JsP29/nKLAcRIzyLtAhIQolUhGWXJB++FAkPX
gVkPXIVhmxBb2ZJsM9EtGxY1Ea7hPUyLb4WGmk9FpPf9pAws9QN5K7MtTXFHIJLS
MqMRAqvImcaVHPu4Czvy5a9NTgw3m0loGNimx6qZB7v3WEIM9No1SMM1lg5FFsMw
fBU+l54R+eupdH6Vjt7FjOcQ09SC+0bEqHQ71zWhJJ4PoTyD8iOHc52Mo87QGssG
1wj8xpQdc9BydKOO9iJVgNAyM0PoDIeP3tIcF4TJW5a34rX7GWSKF5VX0Vp+u5cG
R04ye11YXidmpHq6wQhtuq8bU7pw81igoaV+PUYOfoG7YWM9lqgIVRZlKs5Mi2e9
hRBpIvXd9I4me2k0eAgRlEXCYHyVQ3dafBHpZFAEKrjueGffkhxTZOnKmJUxQ6+N
99HCRFtracuMUHd9fZetSWpiLRBbqnDEXerb4WGWJO64J1o/JEtilkyO1dumoWy/
7Zly5nuxhBNQRZPJ43RY8XFNMrF40ZOyEbi04CnUJqv5gNW7PI28R9Dk34QwPZS9
0YXxwobegsqnNgHSXfFroepfLKaS2QhxjcXtJUg8xkBzYr6456IECs2lDxU4iKMQ
z/ac2px4Ijr5H+nC0q+neRu6mhFtN2TQ7UyWq4pB373nAhQGbe7NtCXZDZ8rIqvl
i5IFoGCzAbHTXd8ydLxXmYlfbbYUr/HTVWFa/1a9FM+A6URqWonH7eev12+QuaO4
O9T1xG5FWq4WHKW0+muc8fXcmfarBkhz0R5lISHIPNyd6357iOVXLCrtZYB4QNle
3HUAMNWMaYYZdQTWo7RCwbgoCiuM3feADNPmhl8QZx2xyij8BjGSJKIIhcc6WbPc
DGlkQbBqkHJ+sg5F0vvi6KIu+snJq5bDx0A9JWE+n5XkdL8d4S5arIXj5rNCjlB+
6+tvTznSiq29iZh9DEGi5d02JZNne8+mDS3FG3gSjVGmDtgo41v09lLOn/SIAzay
wl/GdkISVL3/eC4O5B/TxhPtz49l0lmpMvZZ0kLdZImaEVPhtatyPt5z/K8pNZ3j
sYHdyiBWE8qPeeJrMiRI3RXLc8DUQkb+QoHq3PrTl8QvaEr8gj2k/pgdTSN6nTCw
K/2IVGRKlCqAiggF5wRI3spUDco7MFs+vOEf61IVqo8m1aonYxm5gMeaUyJ39Xnv
c9iUruWqCADRsWIVfs1Fmak89Qp5FaQ82ayscIuvK2TZQEJcahER1RUU61K+lQpP
ocUGwCMXaKooFaf7UtJm6AtU87qrRzU4BimcCg5+ypljgl4t5K8AY7z3+VZWEZQb
yqy3xSk9+KB/iPTAXXmqQtB7h1RKzsYZsfOOebmyQgidXl/esHdloWgZJpzNwM7s
zOjQ5IBJKproMmycUDaqD8YnmaLdXaK7r4D68utBVogXvhSXMxJ9Xzo/Baxvg2C3
ibGG0qO+bwKGz41VpJECA9s71Vn/eZ3PfrtlOgNpaELRmjdPrTcyAX8AEWfvwvBl
VNTYfnRDlhpYNJZZveIYOQI7HaDtNCnnOU/Zq4+MZoHE+NXyWY6KU/b6mraHnZSX
NgIzUJHZBznzKNdbAHCXSzNygy2pR0Fr0R17oI9G78xekVRE4djDVPTOfe793/Jr
xLPxpOt6k4tJNSDmRTmclIGNi7I4pBshOOqf5HYce1iNfnc1FKm3TrYtvvdIoyw/
Itfzrl+hCTcDToFwCABy8+F/EJVf32+odiZ9hH3n8XdRq19wNiTBkytnlW8YgfnT
tGs13Ah6y1GpDqC0KpkOTPfd73/c3DEZIzngrqYhzLbRi80j5c+J/VUwvuXVLRgF
nvaqReKBFRBut1MaR7jBENUPjKolLqgnBQpubEtz5jW4xLoZQA9/ycH2QfG+NIlB
bnCfq1MJUkDxNiES/HQDR5YrI3beTx/O2g485vWX0Srr2bJZHEsQkifneBJo9lkH
6BMrFbqt+XNZLcDTsds8LxCarDK5FvAm6ZwVH5NSSdLE6LdCeO1FSKfbd+4/BNy2
i4sJUJ7QCoOiJ1PWePWvhxNyu0Y+GLAv5ZyHCcA4YxoplZArDoMfXdaSvSG7gevK
wfn/HfiqECE0JF3V/3ifPTzVryKiFg0wAeXF94e4dob0ernnSP9hexr3NWE1zNrE
5urfqHknEDGz//qqLQyhFFdmXB7qKlMSmUAjM0jhZ8qRtW6nmP2QJpf5q7nBqkri
KSikWviGQ6DKt2UKDumj2mJisyd0OjOMbXjr37ZS6wsmbKBxWXddhM/fv9rNment
Oki3WuUY5iOpf6BcVFdh4Y4BgGiGo1/RaRPxCXs9XBzGjC0HcKEEQJaCenlqe4eG
HrZPGTZgSbmXvZ2qgrw/ZLR/hzrmd7h41GXNX6OSjlNm41MiTnaj/N0Ycw3wFUfA
cKl14U9A6qpL3JE6y2qqESrVOLWhKLfEct+kZxmvl1jWSKoN+ap6E+bdfR+2fj14
4IXv3gLjNOPVoQxYILXvfbcuKHEJFcxcBAwxMzB4tg8MNcusEzNqztf/EiZp/xxm
/UwH06fp9+Fg3tEUVAqdO+iTQlioa4HiNYYWqyGQziiLrW1hcQdJuY+LczxWbe1R
1Z2eMf+gEY28lPDH9GF18Ps3z6tcXMFSdgYpIgB3zAByMHKYQGfxTwVDKoe4InLi
jD5OzsaXbGg455XdQT/Q/uUwSx98ELNtYE5smQlbhb+4S0SUqo3oc8A0AkGFUgUq
8OhjDyMNp6tn5Gb4LqsbzgEkQjJZWaxBp+Mi+RKgVcR98kCP0sC+4Z5OOjBzMZFC
fh57VMmo5R0ZDNZ/Gx1/WsclQCBVBz+/IYZ7c1qtJ1OUSDrtB/oqakDjx8YdfGK8
8HQZAZRTJQX3yioraTvBlsqaJMiLpgKo0QH0Mg8qaSEKW9Wwe1kXD1dPYLus0qsd
uQjCKGZsdjruTLKXkTTm4FmiVsoxMmYTFI7+bqLm6PLZ+DY+iwEjKt7E6kovNcNb
p0ynGpF2nC5QArSvxSwlro4aspW5msnsGjjpzA3EEFZmWAZiTrXmITkFwZqPQ3Es
YB4rTIL54sWzm3Te8MBuPq2kDIkZcEeeqrDYC4EcqzzD6W+/2QatM9thEY4XpQup
auDajRUoRIkE7CFwb68+XzhePa7x3daj98ZcfCKLSsovVc2hNdIRRtkltW6vRXkc
FvSmushiGfPGmlK3no3kc00+IaDBcfhvEDQRftq5LVYBnSTpDkVfWuFB52tJ0Rdi
+Rvi3jVmyTi6DS7SsLKz+uw43xiMTEA0GlbT5KtPyPQ90KZGuEZRqRDnoo896ZXB
uJN6cALR/Ke7NAPz9FoJx9h5QnceBzoiZA2/WQthU1KeM2v4n2pHTI+jQ4KARh0S
anxkOGiMFeE9nTqg3BIMcARrR2n+ZBOFZfJxKsHjXICFMG+ZXP1cAUVT3H+6cXc8
Pn2NV7eC6qXki2uriJG0LmVNBYzCljBSbiMINjgDS7I4JFysQiL+cE+bWukTGNyX
4I+D6R5fw1VDS34WXuSVuMJdvDh2cQqz8wwAEEfAqIdhOIvs0394+71NLpr2UnI3
CFQ49hsSn0m41otKGNFtGIU+PxiN+meKtcMcKigkicAhz0dCcBF/kOCO9abZuNZk
T5+w5o1nAU6pDAHAjrv5b1jM3oB3eSrwXRRn38ktzv1b1x745ySp8+4Pj+W4cdBP
mYBKyw73GfqyLr7boUtTyk3Pi1pyGM2X5cMlCEhMwbMFCsxi6+ReuUorafK1hrbE
0e99Tz1HbEQ9G9NzHZaxcT3rty3pJDE8FtZkN71uc5zyoHJTaNSNPP8aPMhtq3d2
Y5Pe+PD+uzouj0STpQmkFrO4WT6LJMKbScne8+xE4NCff0FUbs5K9mglLXR9TNbH
V2cDP4lnS9OB5lYYhsrlSkjA4Ht3DYuT+W8uCqGJ840Qdn3niHwieb/meExRGeuL
PkdTaY0syEj5TLN1T+VIn2h3SSQjiYLubELXRpE7qHcJLTfHYbZX5LqPMxToCU8r
mGPPNcbZn6NNE4QXsCwXidG1nCCl/qzKohzPhUhwZiqDjccDAoMI9Ls3309XiqFK
LtfURvksR5oYV+PkX5wgGTEhSXVgNHg78EDKD5dLYTfc2o4JEu4CY9eXFbuL9nrh
kLj+Tl2/F8b1/IRgF8xH6l1GPMaJfsQWpxbxim4vtnFCPdwL0H/30OowrmwxPjb1
KhY+wqfQOU7Elp6jtM+1KLp47wnI8wPjeZaUVjScAhIW339EZb7IjfW4JhCBYt+j
qVySDtRGjT5SsbBKpnM+cKMOkJLd8iHQbl2YoBH9dV3LHNqR4GZ/1pKYO+mwNF04
0FSmcbaFBKeWQ618dV7+KJFHBDlzoO9GM9dgdb3Lk9Hv4rmeM6xeg10L6QHVAvEL
/85NkDqHAPEXRU3MViqZF7MVoshM0y87TpKDi4y3/X3kSSkznpz9rx3N4JmMgvfh
YVIj4vUMIJXw2hwKw7Cig/YLlzobGOt/pI0may9EHB1pmHJyLn1UEySSacM+w64g
e0+7D8GNUFttzmT4nFT1aK/lZTdCihghX0SsiFUd0Z7L04vtWKiXVc/U93AaWHYF
2WViOTEkPSvxbdNERrDa8LeLQ2Kmqw4o34FfOORuxIjODxdQLk3YYlRejhrguONy
QFYmm/BPX49TCEclT4l/wazavOywdYxe/ikgmgBfXL7CXTuEJbICxl/GdSReTJCE
HUyuuLr2DG3NqKFq9GTfJhqW7PdJOHSaHYPREAQ8SyO8vGPDHqkCN/pr/fmZOqq+
lVaIIz5pxm/y6zyevXXE5Ks+V8SAZa6Mb4bf/IHedrDf8oRmDwFLGnFaayicJw4M
V1bqKu4W5nEOMtFrSekE+bXijXLE+MlbMiHPi2jddWeJryTdEyq18hkWc097Udfo
05EVT4BCjzSWtI7sXeSpofRIb2HG7g2OQp5ywPbl7WtZZ3hSWAGjmxeauNRx812f
ffQLjlyaFOFf+N3Iq3rTgR1mi+Ibaj27/92tzS55xGO0s5tVc11snhD7ESNVUrI6
5HjU+7ci3MgVNkvXPJMMYKy25qqqOKZhkEppjnjVLV4gvuGqkPn4eV0oXIx4SdgJ
/xPUwGeo2I/bvTSp8+AYfHLs+GZZR4EBordK4ZQj2XUDgo13GHGyn3GRccQkEQDQ
f/leuBhC29sGuBRCR0Ws/JwGIsYxdtNyK4/6JLGcGNvrfM5jjwzG7yMFdl//MnFy
AHh8va6+oUU+7vXmTe40wW7j2iw5AToIXE1d3PFjQVKsfpqUb6GCBGcOCS9W4Mnt
oQG+Wl8eADynEQIfo3wAtvpCjHMUF+5bqz49sItXCn1O0AW1Qptljr6mFBq9Y5Iw
znM90o2Lp2Q2nH9p+Cc0DqxJeK7/fUOXF+4iPKnMfGDYnAZCXUvmO+CjGEUI326I
24QZESiy4MMxAhzwrICYr5PjA/MNVrrxmSo8ZFtjHjsa0du7XVcVodL0D+PZ2cF1
aQc5ezZnfHm+I2TDJ8CFhCBsmvgq73KyshLpuahtr1kH1dez8NbiW83Gx1K6sZkt
lP75IB0AerW+159h7oHMhsT4aOkEIhkujD2Plf7agofpzX9EPCCJnixWpF6Tgxrm
Hn9NeWg+dX+d4kK8q1Fqk02hd+4poJRt+Eu1ipsqOPp/4OC04r/ip6uaHZjjdWd9
0qTeoe7YSEjLREL6jpSx32KIFtmSPp458my0NOCBxjyyr4/mmkUFvZbC7LFtM7a8
RH3RZ77oQJsEaCCQUMawuCAbKlT1/VhMuD8cwMD5i3GDmdxljq0nRrYhjnIDdKnU
7zj3JsnOS96j3YQTPJNKoD8qtUBg41cOJY1PlJdUuh6fzFgZK51QY1b+bq1RukTP
ZYCsISI8sGAPaARLdX/fDEiUmVaSy0u/NCIgQ32kuafTQaP/TMhqL7KUGOfpChel
tK8PSnRNFK0kUvUvzkHWzLFVXHrRkvnnk7g6vO8RYXH0+w/Rb99xiXrEGz8O506/
SB8jvavFrLkVd7VEoKPXVmrMKdu8q44Igfv2J4aPNmh7CxFxtP1IdcJ2ssJVAgKF
vIUn1/Hh1S+ZlNV4c6vB9MWLNF8v7chzCRukPcdo0tNFytKrKznZWDeMyR93E3VS
7ynoBe7K7iBn7IP8T9pC1BX2tIyxPlFSCCzsuXW/SFm8OzxHcelYaKlEa94hVRGh
N6ivPHJFm+t5CFNXxn5Vn4oRN6VLAA0kJpkXMoSk4REyNolhgRcFqQLUNyf9Dh5z
rOmrbneWTTckiUxo7NAW88isNQKEAFACSTr7Ye6ksC0ppEBFZoOMgjJYc/c04dum
uJ14kO6gQdGIOgM575Q3t87JJGlZjPDVibkLIjyiNOYoUSHrtsdbNreDwBnd/rg6
mh98g5N8kNuky+NpmoL0otwP6o/SwA6gJ2IdcGCeg8NNcrfDDk9GSS/0wd17uika
KrGftDqEETid2gb3MiJKIsV74oQMOIWNVXwyJDhISD/ERZXP2XOlYZ2ROzjANL0g
fmBCQ+TK29HM1NaEIlP/cj8WB2cMQbRPSZrqROS0gCKou5NOa+SqG+0IhDQ57sAk
zrHDwXbFfntxgLMGzNSugcWq9GoKR1L2S2p7tNBccd3PyfPmamwjrbP2VLnibyiS
bpUBO0dHMTtfhOkYtwlZfk8KhaXvEkgbpJgD42M5sulE5Ns9KZSl45EbssVsZwuL
tao9RrRbDGgn9knajweoMMY5q8fkaroQJXd3fyNV6trkJ9Jpj6VuJldXpzWkI8Mh
L+4m516paYegRUD9tNNBZE6n3z2RL6bnMvbvi8OvlS7FjgFuuLsqgjeri9FZhTHx
00WAgC9ftGpb9iNclGDd8edbSbwIaWOPmOWvN/009XQwvnAzsbDdV+ETN86G5iTm
4H3NwU40o6is55VpmJPgFUvnCk3I2iRILqCUC4Fq1xfKbIKkkfVIAmulycxCkyPG
3spsvDe7JPHzDPuHVXGL0xB7LE+qPxLtvOAB/8+KmioAAdQmKdkvZDO1f22jNPEM
Utlv4HMrzb9uBFzRorQytC/n7yIMOqIfCkO9ye4tkCPeUtpAAHT4UiQStBtCtXmS
OCRhmAx/HUfeQwC8qB2o01WEdKIPfSfgg7r0Ulehgut9AEmKeBXnqSEvon/4hzXd
8y/+AkhXbZ2wXSSzrH0rT2rNl5HnSDjCTcFHSZa6pipvFi9lzicF9lUSzxoBPbHF
GTTLiMW/fN+o767BjcO8bPJU6QnnIFS99YVo2njV1QthW2F/DuBTpUhwtuX/fTsB
LeK0azsFffOlCocNvGsdKyqa+zSvCuT/QYuR9FUXBMqkDnpyxuR9pr4Vnj8Amxpx
3zu4u+VFn+vX8b+FS2Gp4uUVs4Y8jSZ8aaGGT2lHwyv3730/sOwGJBhydYFksRWA
9bE4j5xULuM47fx+JtAWweRsQ22HOCy8W5/7/aJYn8UdpoY8kAAmlPM4rRjDDrM7
YwF9Xd2q6PdG2y/0bvmJ82clzWUhZw8AiJ4NPgpzqUbHdtVUtbFTD1bNa+Ozqz9i
GO0DyeTxor72BiWWdAVjxha0ISFVxQA9tVGxWd4EsP/Bake3ab3yBOmAd1uGgzmz
y2VYXn+6VZ6XiZN1kDJZ0Zul8yH9JR+jY43oqmWIdb5BmUALmC1PUn0DdPgDxKs2
d+P705Vvax0IQzcil2se8h1/meGCM3WVlf0Rhl5AjlaxJSdU1oVfnSbpKAXKrIq2
yzyEzPzbApWWo+zM4HFYjgkrxss7wSYJiNY7rmK4/S2W/Q38Uf3jSJKkeWMgG3p0
KhACjmto4biuvLIHrcNRpJOwpFcQjrZF5ru/5gAqT4g9ILbDMgSkW5XYHBb/x7Hr
LN9lpPQ7NjUi4z8Cqp0cf+WJsY3yctlzu0p7djhG8yit9gFe0Y3SUv+VCYv/LNXp
Ht3IAMTGn5oy9QTzmVuhhl0nzRyCDmbVUkdNPYQuZddfGFJ/rL3PTdE2Xd1wiegr
v+fDGTt//Az32hX/PUVzUGT35NKZ5xU8RX5e8h/G2tTuouT9W4Zhr5lmwvrG9kTZ
EvJUYCmpFjVL5QSxFJgkn0yMIBxfO3XPOO1QgwPCzRtv356DX8I+/NvEpqJCMJLt
wCsSgmLB0hJmT7ka3TCUIHHt/9zY83IxnQ0iTXOW/GdjIkTvt86MBPO1JxVsHlQB
5hO6nCfKqBveeG4HCTd5nlaGXNWpnjGO9Um3SQDQMhoMoMcuKSJFe0juO/gMBih/
g10pyuU/GgAxI1M25kWTutMDawUGVmbwVom7qgPfq/vP+O9Out0eNDkJCl9rXvq0
my7LHhA1GZhYa9/I6mNtdAXuiJIXF1VtndR0znq2SG4+GuKUtn5FAL2tJk7NS0bI
GmUqdDQjBC2IJrTHeQNv6k5WQH1lyp/gG4cnIvKmZW252RlHiURyTmp05Ye46LRL
I7F4hLWaW2IVnESoeqhpcnsYKG3lYBxcwbB+TNC8/20liMIhy7iXRdVoWJ6SCP6L
ov5EPngGiDFOW169V7cyfidfDQjZix/1E/gtHUfBuUx7pM37tOqUSFJY2S7tq7KT
A+N6zmrYLWz0/W+6BuZzq8f0GbIyHHjLifZJkBcumkNIRiUKIiODg6obtUhAWzE4
RzX+E+SYzd93dSxRjKakj2RxiSzS3S+AIGowo7NR5Q9E8bDMleWMFFEFhywEaNQR
BXQJu0W0xLXD5NcVZnu9f9m8mbx+5gJHsBjwJRkkW4ZfUtb7Z2IrpSnl0F78Ep2Q
jkQeq3wEJhozcPXvJpLTOrwfZXMXK0i3qMgK8T1QaNH4JDSBn7vP/iozgEdVFtbf
HQ+58JwHBJ5z/MoQH0NYPDdBSF97hgLGB7BPphDNl/UJNwssW3YhyCf5EkFSuOHN
WXdUzHUCrc7KEmxpSo4i8Gu5nXLuCleIeL7QC6UeWY7ECSC+Q8/acfgnmhJ1GF9z
s1bMTYxTV0on99LnxPCtFuC69mQv4YMCysypYDp7uistOWllEte7vdY4hTWVOalT
Lewc5ozjLoSHaYWYKua2EZ7Ol/NdumrABEFcTvuOB0YTCXWTZTMb7hUFWNV1Cxj1
hNTEt7qt+PadklOKDfnnXEIf//92fBQY7EjmvvPuPtlcNSsfYUosfWNN10jDTT5y
XzZ6AfvuR7NyC+qgzIAqMZW52HaEnIypUBd6HjN1GWqZpB+1B6pUKJStnRYa4bnc
cDwhQMgzDTEFQ6qCZJzhjJNd/ikWqW/qX/Z05X7od3+22yuuzEO/9WnCWJNXh4U+
24n9XVwloZ5/f9YjqGu9Tdld9Yo1z4iNPiXuZ0R4BfXtUxvlXIQqCtDniP2B/8T/
rsw18r8ePdVbIuhG/DKZdV+h8A9RXjXsZdlYjLgNUGyq7W9Q0Ncwih2haHxSem6R
NW/ow99J7V/oA5cdks00GMU5MyTTbNyE3O3yLqBgJr+uloRmr0lhuf2jsXG5GgXg
XsC8fen81inTuIuPUWhvwWEFF4MCOwTWg0wfjqW7UWyBKNmU+l0+/l060ibmgckH
FXnWRwTX5x+oSLAClp4YcALG02yXI0+qpooLTGN6fEB6p28ajSbIq1SVnxXPm5CB
LZBCfbuP6pXNOQ5rUne+gng+zao+a/uKoe2IjOPaDIviXjCTkUJ4SpHs6LHkezAC
E7sf4qTNHJTaukaQ8XxFFwrxepqJMs46UhdCCrwjDyMSvpvKD0POsaBXwCBW6NYn
/m4GdVZSukg/+DKEqX9hd8nx75ztKSz55QI45whooqRRO8cOmQX0hb73Wo5Hb6I5
pbqxiyhu/nnEvnXTnukPRLZ75xP5QVVGkwYqf0M735ziP4Ivu013W1/rQUVTBqSi
bsAFL4TI6dNZmtLRtwZuIz/ZOxBlsyx0HY3t/3NDsBQ8GyzDoc/BwN/j39Ewr9G4
5s9J7nWnrVBlZvrKkhY+CUOE/+DhGUD6JQi9bpH3diFcc7DbLKRZZi2U8Ggqk5ld
4Yx2Wr9Cfa9/Ce0FcIiTSidYUz5TesZ4oUa+E5xAyFOShtCY005FoTWNrkDEZjDV
VIDPbYkTkA/FEXXME80ZjxSoDwVofcMtBIGkMTUrxqVCGyrsuCyUmoV2ejc1qQGR
59SzzpYj/CNPclGl9W+PrBm0mIF5SAf/X5BBK7p65gEDxL2DmRfBHHy1vmslRV+K
7UH69QpyY9dKGXHDgXs9aZnHRPucdsh5CiyXHPXHNyCmXCkAM9bQdeIgZ7R8Ygya
IKEMG2o12XEXnGHY/KD4pRebdiUcF2Zn9rcNuTGKLwgZ8L+QWZIrzSrx3leXE3rf
ftGvoaBdDIf6ct+N0oaUe+xmNFPWTs+9BYO2ie3hekVe3bVlwIztYGovoTcfSgyf
dABzESTdJJghBfEuMk8cXDlnvhLtsR+ZJ23jaB6L14J44cUMOKtZyXlQV0KXdA4H
7wujMNNJT4Z3DRdnHNwJJ4mFeIPYHnZWxszSYLc5NgL6zInaNVOwq3EaCwDkva8F
kaq5q/AqiHYLLuJTrr6QEhBqc239hLgqPTB6qqPi/KoctGp19t58mLjcHAYuTM+R
A4quF0rsj+MOeoRr2BWvK9nFN+RydOEAvgQWMETyCq4tFXBP6Bkq9x47iRAcF/rn
s0BYC9+wTLzz5QbE74uw5tdkAoRvmlCMF0Cvc1jd2MU9kpnHWXpXU3gIYuNpFjPU
kxZdo0OAEy4PDbV4jpzj6qSP5eIpI+AzN7sMlclrobAini34QRsOAPUgiOH1uGHQ
itxHKfYfwXfWFiw74uuv6/FH1SKa2JyWOkXyrGhjNYrBsrw4VvcBx0xpWw1lfjIe
a5oP6Op2BuXRC05AN/rKUfV2bFgKR2GhY72RiODLn7RskImen72bUCsAQNrWfNZU
y315ehA0vCUt936995wCdTFj1smAs2X0PrR2GJKhYJ5w9Cmg3cn4vk1MyjvWhZPu
12I7bgw9QhQkJ+3QeZLa47IGce/T9VXZscQVdLjUGWhKK6oiL1MZhRAWzX8lPSOR
32jZzN42CVgC3yrW6hCEjjirXWey7tBaZb8735oWrQbxqvzkXW11oSIGoEv/TyKV
AmS0tRAoqmIGTBcAybbz/F1QSmcnPQXcrM5m9cQCu92y+aEiYpunm1DrEYGkMebc
FAX+GPeJBa5fomqW4h0LlAqVWXVGDp3d82KpJ8PPcaHLVOU0R4iDHKb5RuDQnB+t
78xHWYcgWwZl//VwHErTQONYwOvJHxyf4iJFZMQurFoM1DISpO0DzJx3RY34UkLw
nrzUnqYGMFwDEeWXlc6HNSCxMEhQfGKpOnZSJ/p4IP1GXn5vAfevY5zGJHRJAML8
aaCuROt7Cflnokjp5QnuiS0PoKndMMLHpvj3Mxqz2KfKZyBCjfo0SxYf2B+U9bmj
HGn1oxM3zXPwd4RZbBHfucjR7fSz9JNdEw2hcWSZJNigQENlfubSj2P8Y7oVfQXG
r75DIa0bHothLR41jlUsAVSKpG6ZRDzeLmNVuIS5jkWavx808xDyg0aGFRBuJwyO
42te9s+kGDixdw/sdWBBBxtRfJrJMj+WPQMYVXoiktuiXzkZaynbQR0U9atdkTt7
/V+zlro93NoJWn20U3yqZpgDxone+1hQAq8+0VWOtUkFYoKpwGuXShDrU/UQr1oA
ymC1W9Kp2eir6OGR5QelBy6gdEOSzlPG5dRtChfw07JW/AihF+8tGwWktBxorGlv
Yl93IZKaX/6x/6208d+04BFYN05vtvQBIEHrAyPBPQhZQbtXy3bwfmbIy7FxSzku
1XbPmfmpIA2ZXzYQNa++g2xY8s3EWBSZFPxdZrdkmJmNnpDLkUE+6lZRBz9Bfau2
rzXEpFmNfDPb2wALAYoE/yIqZVIReBrXhruphDAPicXkl8nyl5UjTx/rLjD0xewR
WCMxSl3P5WJ38MnZd2+2ZyrSzk8f+ZYko9hQgGLZmG5zIWFTszCuzHBCTZbSkMoq
Yw+iw7GN5iODpEk1BM1UAPTiqhfBF4usJejpkqiyQJ+Lstu3mxEAFT346m6xDa+7
AlOnxVbO2umH071s1l+JeZ1Uz6qLjVgOW5tNzgiiN0gQayDQ0JL0acKVizniQnDh
qFl4nEBu6k1WP7d8iuHnBjjf47IAdEcFPoTbMZUVdlOKPYSCK/mZU1R3yFVbGK+i
IEQiHg5P+Y70BR+H7v+4YVoMyq0HJFUNNzAaHrwL30IY+N5L0LU0fJu1EtyBfLki
IpVjZJkL1rkMtoDVbxlb+QnFgjIcKisEY+rp7SKjBE4khqP8nQG3KtAvMtRo4WiE
XB6PkUyG1iLyJdy8Ddk7v5mhnVBIGqeC2SOTlpdIDlyMKrS5Gs0byrkqN71YgNtO
gmFNqbIgpU4dNvkjTuFmyE62vvabN1iRRfkeYU2erkYggmdPR7Y1rH326XOlr5cD
o2Jc0ci6JTamMERgSnRefvigK/Of6QjMjCnQkZB9VyhHicnKtwnOcYkPrYKQ9Vw/
HGstlrtqU95xn8vfCvAZR+8AkfQxEkteSpty8AArzOAXHjxbbaGB9F2f2y3bQEaK
9TqqJbYqNlOULnnIJRZzwu1kp5+PqXXn3WQd7SbTW1wfWztfOrjY7T7mBZQBn9z7
yvN91WrBwXUlEG6FYZgBq+Hu532NbPExmBqoewhPg//ht7ucDcygbUyy9UcD6ggV
KF17iAskkM8+p8qruJx4PHzFldQnCCMtkOa5qwlI8kvwig1NMyNF1O1omDIKUk5l
i9/MMd673SrrR/kYyw0t+XJi3jccZE3dIdUdNIEMF57zxwzHbd+HecV9oYXu491x
ZVjiifsAclQTsihqdCxHisxQRQ2iOmdLxb8/5F4H3YEUHQ9XQSLTR7vS1kHY2Vdb
ao8aZsWvPFYTORK7Hz9AZTFf/vv8/xeIWIQMVdQn16pNdq62gVf/lQEst7sqXtvQ
T4KtFRdTICaKZottgXyavg5VhV5RxwTpdFFO7DJwYY4OMieeM2u83m6PZPgTPAfX
T9npyrtIS2PDJV+Iy66xhmcGJXFf+xoqhsfCezrvq4Oih3fvmIuMld+/YIFGO6mO
2Q6il1TERX1tAwLUvsMvC5OqeQFTrhI/9SPKaxL9spqaYZHQnkkQ/QRS2ArUF+Pd
EWMaK4h1D7TgF/oWdbh0HpjT34mfVeFT6p1/z0Oe6pShzQEeP6/wWGXkjaqnRcAK
yzAiXKAAMwPKg+nNWTz5dv9tDp5OUujZUpstPekxrAvvX2Vlalpzl6N3+moz50iD
B2Rmhw2dgu07/pPd9DHW+s0wkTlf8jvul8ByG9JAhxzibzYEG/ACiuaDmlOAJken
r5A5xGjoAvvZJws05nX36dkoKFEM8rzpKtq/Y0s/J9afIum680kwNnuK+Y7o7IdY
qF7KFRoI5IPKkHf8uy0JwLSO4fwyp4XYk+bE/oAvLGAkbV+uyzegBtZqQWBAetZl
vBVDxdxAJ2Df/Cbsjgx1dmNtdfl+CexaRbsZjEvKrkH0ly0stS+aarzpFtLCn7vF
RPAGbh8OoQK+Y30yVzEL8dZapCRli67Bc09YyW1DTkPD/xNd/bNK0uUkHzQ9+nm5
4wJJfUsrtL083fco+BU2VTYB+R4/GVAtj1MjW0DYVMfAiQ0gAkIVAZ5KTpuz3D2g
izkMxod2LrBmDy1xMq2C2MLucFDP30sb7/lHtgD4ZzCgnu7TCsymEpJkECw2Cs5o
4g6czYHHDDv0sWH9LO1FTPpylbSHRJfRjkBWwk4ov9CLYf9bxBn81sksI1DpKvqD
mBxEByh5SbetZKJBxWJC3At94vBydv90tt/F8mpCkEIspff11YF7otStfL+n42QK
gXwVLlAllfPGiPJST0xvDRDwyCHknZ1MVvxsX8x/Pcy8YqzbP8dSPm/PiGb70Gyn
7KmRF7Oqb75Kmn6IoR5sFZUj44bewyRB+tHt5JkcQvHJ+ML6EvoTxMTlB34H22Fw
uaLuBTptiTPRMCzW9ROZxLGKHTxYJMdpza2DF3YRGGB/erML3j+XSMULYNnhEmL5
9OVwPSRaffU1I28yCWTTiDPbohJSHd8dNj3H0Nht60oG2o2VZa5iYITWg71PUThf
0IekOTqSmVESGc3svAXj9M3JtUdUg+E3JPnaqlrLj9RAgiQTjvN/Yndq657y662w
FXq/BYRyxr0AmirYSIWU5EdgXyHOK7tXgDizgEp7685/m7GtxOLFVxW4Y8iXBpjZ
j+NVIR8/7zhvKl05NjBhDy4/qIHvrcaWvAnamFuNOpURltjdYzhRtYqUM65Kmv20
F9t3yy/rR+y172UgY5IbaxcMpNpQPoAdXetMqwMmyeF7wkIYL3DUPVK2DNDH0MzO
c8dNnsFwFHjRkCaMEWZ49o8laVVDDA5qQOJOo/qT4Nos0hnIDWP+naaqcU6eUdZ3
+/sjyCwlt/mwnYgqMYftZ4Fdo3MC0XXVPOr1BJc4lvskGP639kl7T1x4AeUw75VK
EJXmfL/JebD7HJz5lcCuZTlzxhsJyziKy1LSohLkmej7nzqJmnC2GzJ8o73mm2zz
u7oLlJMeTfDGoBC6MlAnWEkq6rDnRU2wgAAjHOxyXdLrhVgoh1VHJ4hYMm7GlZun
70yw70AwTmlHPihjuzJvmmQUgMkzFK60XM0AvCRq9DmII+LliMEoyp03eH1+n6Q3
lX0xLt0+WAy7cFi1gtXby4d/dc/zfLPWvdLbl7s6NuLft14oaUb18RnQTSlS7uXg
J+TSB8gGB1YPoUWxePwDaIPdyPcx9Dz8f+3M221nDJYsilEEa/R8VqD3B+wTHQmT
Y8TobTX1Mb7lA40oQKO4Mn7WRLS0zUtbkOjyRqWqMe4NaV4JaNcJ3+imTz0kZJY3
seQGKqf14HVuyxRmzqInCavSG17B3aRpbN4eixDsDu6aAeaNRyfqVSgPOcfGX79b
lo95rY1eCeEgzQ7XEf0le/w0k3Ub9T/2SAdJHYFcCS3peUBD3o8JZ1aXTiFoJMIn
QLqvfie6YL7DV77rrmfn2yVwg18pwFkNQQbk/OjiUPX5plajxmW5QWZiv8ThacfD
UYQv5SF3pf608qYxcEZ7O7NFF9pkMTWw3xBR6GqxmrDsBieRcRE87pqV28TJ9DRj
XDj4uiW0SUUhHBlf6JIcNykGZuR3oiSPXd2xPqjXyy9Vwrl8V3Fhxw/sw6Wc7qu2
JsCPD012xTvj780mHQsQZ09UHYTOUbbG8NtmeDXSAXsRM6SH3gcZI1depQe7lsCt
0aYInHUg3/bXIIcPYpDES/YLVnAn/6/T4S/4PAw6Y7ZQD3l96qYW9ZfZmQ3fwlCC
KL/OQdO1zCy0c5i0yzv9W2A9cgsG1WI9k9lf91o+x36J6fUs70tEJopHSEVgdOhb
0jMN7KDI5d8h8fVtG6+2hSyMnepAEM+rj7mA6tGfMr9muNvNRot55oxB7N7wGK4o
m0KxXF23Vv1Y5dOr6M/ad3kesZOuHksjdc26YzafawT6uVQ4e1gAtsrnHMLDylI2
fCAaqsWQ7Jlr6unNk7ycQMBAKPlJ0u+xHF5RCcRcCvXVo19dEUEMjgMvS75EdonO
MEEgvCAGNTdBOeeQK0Z9AwuCsdIsPFa/rD7qSuweeBKFPoB5hy7Ecj4yGHV/9MMA
97lbd8WS1QmjqfcBzY/d5p2HceF/+zc075q0cx1kdiE75SYPbHGqjAAY/F9/1mxJ
svPFOzeBR4OtP51ykjrF8LPmnQo3A0//yH5wulrfw3Xk0H2g4dJ1DiCp9tdRqdRO
da0oK0AJxIZXALuQrQMqc3Gu7o4fYtnWqlcuZWHVHE3IKL3mpiDrHJcXXc+Ue2fR
5tfFmUrKLlN5xg/hzcQv8ZDq++/qLrooofhL9XhOKaOv5lQ140WRQuqsRJfFKBMJ
iL7Zn1zzj9XROoou7SnXPRi8+Jtc9RJnkGr3w6SbAVrIrrxkyxq5BE+6txhsAZ+K
faDrKg7wcYSF0fxMS+4RC0FYd8tqtqpI0HKpN9e8egefcG4O+yQE2IDvSEJENtvQ
cQ4yYEG6RofNLrHkoXOYBG804jJWFrOdqn9DS9I12wIF9y8E7ztXm3UVld5DV0Al
xbsp6cYYLlJPObhM0UsqtigT5YoIcshTP4Hixtowep1PWtKBv+SAyfLF6GKQO6xS
8GMhLeXjQgbspTZRKxosFkdbQD7hi26iFmSsD6PlS452t8GF4fSPw7t8Z45po87w
oK2UM7n9kSzu8HQ9ZpYhV2m92kGVochvs8CpI3lrlQ9QFWZhikq6f/BftqDBxqC2
2D4yE5ZjtNwPL95EjA5md9MlwVIZVjRcPumSOFgAfCjBMdSFGH7PSFNYxQH7NE5v
8zYnQrGTOpm8k4ORJNlGwH42STk53F8uKxZMGzqG8WghiSMQBFndQK8bwzSAGNzM
qUyRAy7gRVn/KEZFE3xmrO4+IAGWQ0AXgxWQ1pW3w6Ggs62oAldVWoWGoqniMyyt
HwnvtsU7PHO80orIg+7nJ261VD0j/+45KfgXwB1ktOwgCB+ebFSX0E8abaEXWXOm
g+ehzM9fU/aq2OXJVSnlOE929g3Jeo9DYDszkO2tJRXIb+CaWX0zGNPZBGgFo39V
+xge9CW9/DK3WzpQExr6ahhBcvGrviGZgMeghpD03AnWJNszj2DvtP44bn+W29EF
td8n0R4YIKoZCTfvP32C8UxINobyXTzOYncRlU5RnoHU5cRl02n9t4TPRtuft8Hs
U6fP3q4cT+YwPXZzRxLFxbx67giV2FeP6ScdNv2AwLvc/E7e54COX1zkXzwThfE7
BDG5nENwSjcYExjx4YmBCQ/b8NJXgivplwRumkwgnHC7Vrob5Jm666VNk9Tx+cre
SCd1PHCtpLh/lSfKF1wfzC2TjV7tMFi73Q0CkLJx6ojfagp+9VuIF2QH3mZfOPmp
IOYFEzQjhZ88/oPLVXCzquIwkN+WJ05KdmqoNA+uEmMG4ZtTrHhyz0OufGaheSNu
IsPv0RYPOMJoqMf2PRETZUirCkhiRIasZes2yclLaa+gGLpUw3Bo1QUfEw7un25t
Iufh1C9oBNpzhc4Ib/jZCbWatwjBFpMZsHo2tFv8W0lL3Shhjj+IUasYo4U+pCDd
aFE5CKOBEFgi32lxVnIT0FW1f7HPwCFbk1V0ZMZSHxw3F5BACIfXbOS5zw+ssD0w
8T4GfSJVaZjke+aZrJhI8N7jJtN9dLGd9+OjRi6Ag2zwPvYSjocCruqKrwTwxEn/
+JHpWzPlMjmW7IENGhlTVi/z/3zrYXmb2pWTuhsL92QutV3ZkU2L7vZGf6mOPSb1
wVcRLs9E7rTR4NQKJI5YNHZGhG7eM0rpSjso9A5qjLX4GOZtHGDrirYncxFKyHko
m30Mz2VD8TxjfBmujINjIp8bUSG80GQubmlglNijmY/HnxbyPXCxPnOG9EEJVXp1
4gUoto4UlbWOxiqIFzGyb9UYo539oplXn28I5vCK9OE+NLmKFBrUbU5owlnygHpw
akNJNFMhFEP2tTs5WR4RjFtQO5CgxJm07mHhcUrrTnlDd1cq5/aFynEks0KAMnWI
6mMwZ8mwlAcQwgGFqddZYZOgArwWm0Ix6UEkSQtEMqcWAj/hJsrWhmIDXbORkTJi
G1IBEmgQT59fpgLZE69wv7i8oH7GKZZtdfSTM6y4jfBQqN8vw9mfq6LyHlRM+Kmi
KXTaIMlUuYThCewGGJkKynLPuGvcbciDHsKx0mXSCU/2GZ/puwUKFwhpUbINZ9R9
m4FS2arXWh6KRFJmW4lVmVRXWy96Uqm0NsuGUUN+hE+7rbJxWjQ2qFnckOS5Dj6Q
aTKrZ5p0Qx+kNY9TEbDejwUOlFD8dbCN4BOEEcyM7qk8bhdRYUxRGwq8p2MYuIVQ
4XpGfHcqnOPDjyIbB46ZPQIMxX9Wx4UzYv7QKVzZrAFTvgZB0UNGfwMZTdFUmIib
EkBskU6LXkqplKxpYZ58KcRk4ghX1+dnrGUCgk9o+1bOtLzhUwcA160QswA1NTFd
vVMb1puwHEKXKyRR2TxdKN1genWyW26dLhf2dqACfCTmI04VLl1go+jTtzmSoeEs
774y6G/6eAM6/3P7EJxEHeo1qCzNVw7yMjexOVwXTOKDm4JeYHYiI9IKioNaWz37
6ktHEf7AOA9ULu9w5+eyUxpvrjTxjstu5KF2/HJXBudVeKgXTfrNSB7jKpuVftV/
t4LiI5KVH6/vsQGBzaEWr0+zvlS27wyj9i6Tn3nGjgKo2y/U1bGVjujXnqmNZMGJ
kvVZm+7lwQxmp+5K41lFnre+fN3e8DOrkXBawQRbKfoSiQLGaDDLWMl+xKC9gFpp
FLGosFQwl2B/zIGpkU+6uUCKKic4JZDtuePazs9W5f8QIry9bWrVMbIfcuAQn7EI
dI8xjVAOwdul4RCVh3CvOIfrNAuuz1y5p4Qq87TAKb0PZPpLbBdvMhW1XvVx3f7c
BvlpPO1CzpI+T2lUZlK1GAxFb7cOBv2f6TTJrTCD+n5VqzRWW5/DPUAawvH9t3xg
C45EAwJbI48f3mhhAzQ5JTNau/0T058hPsBWOmPQG2CTaLkKTyjz1lz+LSeiBlRe
hEdmDLhg6auHdOU78CESX4GHg7Bn/yfBRqH2kcqEFj2jmig+nRhSoaJifGylkkeN
lnykIglCgVMbRd2nkUJGySIJVj6aw1hw02tZxrXxmlsoU3F+VYCkBR7gFdE8twbS
YfJ7ysfrIAgB5p6Iyi1QwGesBqx2JhRQo/Vdidwuf6vWJO1tNmMo3HKmNPUq6xMg
6K1+1htGdikwEo8oc2mOHDHxrwukAV2jd2MCMNMN+59lxe9YryE9EB3O1lDIqCRW
pdFmIqMjFfAZ0e3gRMrfd59nRJfpJk3QQKtqr315BcAiBs5StfpKZuOgxhBfNj/5
hYkRYtUJtNa+mwQE0DDLRcMP0VLwPChOAYKetP+F5w5SPw5L3aqD+CAmFZAVzXxk
QTFNk/6QMjcJc49rP3ye0WJXNzJZMwCNaQKlI8obXYIESBA1t5FvAJfDtwxKkFOt
zjPuELL31TRQb6hASSLxN0f0yXpKu+Lgv6qDF9cntnWr5doB6nxRmktNdsOfdkK+
NI5dHoqwipziZ8a9r/cMcmTQCRn7qA6rBfX0Amv+w6FYq/yBchrtVKh4fgR4v+/S
QEvNpsY9B+BtcSNAbYN0kd6OcgqhO0ToJQrRfhZmmVrNPM7t5Gfh4ON7AfHVh3Nb
YG6Z7bLq35oFpsy5l409XkGid9EYJ86S6tolDwPLz9QjIpUyd5AptFiy4J+WjxW2
rB/COgnUlUhfL94e8VKTYzhENFd5oZn6VI7Wp1dxNvRfx3yQOomdwxI7FyPMqrs9
C78kiSfTrBC52/CQAfI8e2Eiie332+W45nMaI/cYlkwGnJfhiW9tgAN6WAN512TO
B4+Bs/V44L2qp4jI9NAzIuKVMcBMC8GrPtbGbj+EFTMbG8mOjVvJwxdgybbCup7E
wfnD42E4uMhTAzo5IRSbhK2NMfx/mVC8JowRxoK1HUnaRtlIBV7tDtZfzKsRJ9hw
WJagQjHRPgkCbuaIIsKpem/1MXY/lJhUbOWrKi7Mk5+2wMJ3p+DgBMMmdkzVprpO
xFGndkHKYyR1JXFTkFQmnDa8xE6kCloWK1yTbndJiqMlg3e0hHe79hbqexx0Kt1k
X0dKHgEguNpY+PDhpPbJTAUzbfVTArZJmrquEM4GEYIDgebC5oNWZwW4Yi5QEJkW
g3q0XvdTPU3YG0XPRYInFdIeOLwFjCUxwyqDG7q8K7gZpLl1O227WjIeOt+jyIA0
5mfIPxuaxut2O0Yo6mjGXLuuITfA2EN9nAgvozXPiQhO8GPfHvG/ufuEhL15ue2H
NfWWpfwc8PXgmw414/7oP06jtkdi2qYJrRmdF1zS89xjn3l3WZ/Vl4io32ZzJ7bU
Tw3iV0RtYSAfK0p3p29IXDNytmuKpVyExDhlqRTbjPiN5+Y+1NiCQWQlfAixP7nJ
sYyXxTAR8ABuBjQ6JNWWD+OG5OyjWmxx9K1zo6MdUKKn075RHlTIY1jMbuUOzFdd
cqcObOv3j6C2QVRjMWoUr3zK/+9hGjQ8C7Uil2A6ixBYxofRkn3LVhSEpsA8CPhW
MWPNm4it9EY3Buqby0MfaRiKzXdOQtkoSTe773u4HX+Hl3ghtZWzO+q2GXEBRK3T
HRjy1ZSRWkySTnsAVxIGLHHBUufQ/PUFviADUlheizyhOyW8aW3B6l/zOYQEhqTW
vJhk9vdySI0sk6jtXsZy8FwKbT7vB6KnQIVas4Z4HxkbjP1GH6peE3uEUJxEfyxb
j1hWQ8X/7nDhtQPtURHmoLKCZoBXjkwSuzdIGN/eaJ5+I4/5QCNiB6xhRe0HU546
ISfcV0iFTXIqtUthCf0EG/a8pr7MYh6bVeRp+uvJbr4+ET7yrKwC0Kfib8JqGyCE
/fl6c+bGDeuE2Wg61RY7eMqSL1FrJOuy+TNh3y5jObDWqyudacYwXJHLd2uhymdU
LRpfTIqM7uDk/5TDX1YaW8k35Sug+aT6D4mKaQf8q1IEV6flalEgWYS+l4fqf40P
cCPwaAw4pwvefh+2MnO8cT0mwDPVAZGLl6G6m3xd3p7olSsXtgqHHQ5fBbdORj5r
UkyfA1+xhWQLNf8UQkfv4Ox9NAoxNg7M7XW3T6LHFZMleS6XSQ0He5hJwNvCSpZa
vcofwr7qvaDaulgO5FFjAS3SjLcwoBnltB466VtCd7aaDlKQjJkwSLRyfN6g+N35
nrxyJl/s4PFXQcrR+gqlQnTzxrd+t4X6Osgs5YYSyEY/cYJA3EE+nwGn3UwTwTIL
s8zc2cq6OQd4eKVzyrdQMKE7LI4dswfR2eXrQJGdmjkGtSYX75fjaQ18/cjTM/Aw
2klTBF9hWYzLDRjbB5LmugLO0xQwGHK4yKXlFINc+8/yf+oeRTfq1rOiP+thvsLp
buMEv1LacSwTHqZY3YJ6YKI2KpqPmMkFjLabUCcG+1MY/HA8Dma6RWyyUAHcvInw
Mu2RrJCfaL/ssNrXdybADlGH/EH5Xly27BMRN//qa5sleVfvfkecnJbTITfKPBn/
F3wf5CODTVYQVraRpC5HEv2jr++4bW3kY50iGDPKTFBXZ2uEEKiIQxt2AUFQs7kp
ZgtS+xiXBXs48bj9jqmugn8GEVCwkQXy/JsepKrM68ZHkj/4smBMHtqVOA3jKGQu
rrC7nBw38CB3DzY1pOAdYWOw93wBoRZ3cR7KPi8lFd3Bmbtu5OnHYJRQVpzdkkd0
lNn5Kg1O5uPrvefI0z24YBbqFLvTDZX60f78sWFUei1CHRQ3IKENVomMQUslsSLh
hOrWG5Kio8INfOHHsTDEpTSoIM65j05Qx/8XJtL+i3qSf1uAcGUai1lzZRuWw+Ov
3DhjpsSx/4XIYkNFGe5b+QXRp6pOm4EBHnyB2G85n1BnVp/dkcXVizhn6UZSuul5
s6Fpt+uZrvnQlUHAtwC6rqjh0JRWST31TD0Ef6dsux/oyMlxQcewgvpRpSvFVNz3
c7LYPz9omvthrku8hpqmFe6U3SXTEYXQx/SOb50qo0jKZwvwTMFf3iayQYy/2ep2
gffEMpPFZFHGPxtQRXRUf3X6k7B0TNlSumKq221JCN8XyAz+VqQKlDG6iBQNmI3X
ZaR0+QK60HpQBZjdFsUZdYOKwusIdqt2K5eBMQDre/WrG2P/1rbIXJNvsMF3bCEk
PBbtR5yPgmR87J5Bkv40USHiyE0rvN4U6QJLouTROIdvuhJGacqGHN/c1EzMZsD6
DcsrEjaz5qgbZideJTkxDRllVyLsQ8wFAbHds5MYRL8QiGRGsOW8TdNTCrQrJSqJ
EdHGojQgR5WZaG+yJfRDYYS+AxF3B1twxBIwRj2bc8nzbHg9/fUCBTUa4A710gD8
QLGz2RoE7FX2LZg6eifvocPBOni5MsGpAqUDSXAEve1/tTRxvj2BNElW73urfz3h
RP7Iid9To61JNfJnnheGJi1eMG4GBpeP9evB3GG8mu/Ayi8D1/XF88iPfkRShwAW
aFQ3W93FxhwQuIs2HrPV3uesRBUCdNrn9Yr+r58s9r3rohqdKjVb9Ec8srey2atx
co67dxobB7XNwih5ViCTZ/bQeafZoPaIFDnkDNPdjb+HdRyk6B8AOuJ/uEdvHTLz
i3L0kHRkqkMhvYg/xQqGXpvz2lH+8zUtiLOmPxof9WrCpOCiK1diQayBBYode1eE
ehIVwwKgKi0pkNVMLCQa3xUfh+rI3DkjaZrk9GkrZhnrR8ud7PrWQ1HarZE6/B8U
obkD1h20mgYjYLCsZxew67ABm2WKwjE+WWJxcerDh15dBktsw1vZdc5ZtJZnzjeA
Zo6lTdNl2OQNWB5myqYlAEvY3QtMs7amlf+RKA02DZAr5h1otb11Iisz0HkXJv+8
Dk65yP40jAJPtK6YCp3/V2FIkCPDBZa+MqMiOw59NqqQ35xS+py6PMbjRUGQWudW
+DqtgwQomIExBsW3dBLKv3NSuuFFgikub//BrwZu6rHVcuk/t7iyEf6roj2kkCx9
CXJddhtSJvgURAOCi8/0CLlppHDx2ugEjHnoiSzNcMi6hA295sc/8qCR07QdseV+
US+GAhMu4A5ccYIZb029TNodfIaThIGDpSpuXfvvLISYSpucTHFdx1veuSK1ByQJ
VYQPqLK9RQQDy5W/AqKFtra5fCmuV91NFtaqPQ69YbbOJjp2TIFG68OvdLqK63mN
4yiOkXNmRNk5ilGZ3NALYAXE69vzq+4vT8J0wzWGMgJEXgBmohqLVA+wjHxlKRi3
sMYCyYrQQP2696TnVd2GFrtOID0+qkT+kYnYqg1IndXyN2iXESlukjNE9iNUjIgL
F9DtSsuzt4WvO4yJATk9GazZQKZdZLVtf4ZAC6yKvvHmb41WbFuw2cv0V0BEB7ki
nfro1R8THgw8u0X7Rn8TkkizOEByErNpc5Cnz+ABmRvmBE/ZtG7wn/rBvcpjyzHo
lHYrNDmERCC+XW78S6QrmGlkf2Jtv//lwWHFISlkIzbcdqe+zZWPvlwI7sQ8KBpi
tksirrjT9T4i+5MNIjLwhY5EIYfj+urICEafh/gR8TI+QEQr0j/YZLNPz9SjgbgK
GeKYsBj5KFpcn8oi8Zj8RCqU1fKXGFV/Y57HUSy+hcZ7YZbqeLZdoxkqB95TSyf2
wkWLHfYM/iGooISLcAr+ooVo7qVGC8Ppi6e4hj4dvMBpg+gl5N4r6lnrTFJ6uX/E
EXrPHRl1Sf81bxOvoudy0UWH0qyy9b5fr3vSAfSiNWghtLy9rMWZoA54J6/4S/MZ
IRQEayg4z0MkmY13O33EYlfLSC9cEuMac848Wm0lvjOOB6Uyx65vY6NBMWxfnCTY
2/8BaLnrX1lVKkHgj1qmKM961UlFiI8/DdhY7qSO/TqC7QKM/LnNEDtJwzlBzIeT
ta73e6CAICZCJUXcf4tlCgw4nnoSQolol71PycH6LKXb8anFymvb/k/gg9aGVFv7
Em/WzldZamstiQKZnqGSvn6/R1Bsi/GffyxlPCnG3/N2t4iTxoLG5kArEmfYd+51
iU9yjV3BLnmqDUsBxeiJSBlkdJHtiif+/nSeIH0YLwZ8ZTdsoPH7VWlaZK5rUebI
OrSH4i+wF/LHUSRvKtEn10NsqTG853wqjVYSAKEh2c/6BxAGYOkYJey2z6lEHZ5Y
fWvtum4c1F9XOMYx9EHMAq7mXxzR/KrX2b0CXJAowW1HyJkUWx0f50N/QwBN5AEM
GjhEJnMadBxhrUZoB7aOe0J51qP6MCLQ6tWU6AiJJO20jpKQfqbRaPnkiufmyOFJ
QJpfJElmatgw1Uj1628L5CNc6n9QydAFOEu90NZ4KiW4zNjVNEXPNvLj3UZXhvLQ
gZtmGicW70sWyiV6GFoBryt4oqFAgXRHC2cU4RnHhnz514kHx/1D1aY28DSnHTnE
9KWRQAsQxHSrEfwUC0+c5dVccxNtten8EbFY4Y3eUiwwK9pbrRBOInlh2yeMnCmO
TL8U7SpEbbqwGdvIum2PzqX/xV/oKU2Zkkvbw3UpGQZlsqom9mNKlNBGJiOWCbL6
ZFrONCXjlMD+mQ52CytOVFJgOwmUw2dpx/MHoSq4vktbXG6gKabQlDLIXzzrLD+h
jHourJ3juazLKab4l4zdTZHvaYirTzGfg12S+zhtex/GRNBFD4yqof1bc7wU69LU
Bu/zETOlQsuq17b0LTdIoFsOHVIiGSbVxfqR+1mh69veIolKgILhFC9poOBVPEIx
AAv5byvwRIyz+1HcmbYDW7BhTE+yR7R9kCf2nFJ1qItO+PSPRFGhaBNarGaSWJOY
8Fr0bnA4JsMk2TZM4XxdU6WuwBI2ZZEqgzLB3LSB5+HETnIyGBMnqjCvAcdCsVly
StDNI05dsNOgSMQN1CNTgQVqc2yhybq5/e6rNi6wzcF0ImD3Nau0+JDa+ppSdJl9
DbaX8CHoYkGyazhTiA3etHl8B29eHmK10aYcomgoB346A0j07WTQxprcKRFIwuSI
s4VZJtzi2aJ6fbAptDiBe7LcdSbNFQFn6CN0gRzwz8nLG5xJ6BbTjkfxq9iXwMcq
UxDx6iciPb6ng2LNW6Rvd1kuyn9jxHKOhm/l00xJkNe9qlQcksc1MPXTEHQPH86a
A8BZscNgivvFH5ZiOE6GrXAdHG9uVpHCMV29s/+tiW1dyB5+lgJKS3hGpyu9FG7U
4jzXEYmKqJ5WINo+5ouCWNhDsNOh9NdG/Hp/TKvri3LKRR2q4EfGtaxuNMvGvEMC
GHv0cvkNcHxKC2JLiEqb02LDwgMr2iJq8U2eybo3R3YmiCirK/vcqemHnhmY5sT4
g+mX1gF20HLgJi3ZhpMxAxWigV7wwi167cEeyIjQTv1MPoDii4LTt68oFG5Gx/Lt
wuEsAdCevZnmUOYvL5C7jyVpz6x7nt2ZUmQm4plcd4/4GZbtctJouXhEvIrDW7Ud
fYczqq2cxX3dHchyiQTHRkSt1ixBS3QGjN81tVQcUJ/MAHJ7Q75hWvVgCmHn19oB
7uTDV6pfG3gHmmyAAE+rgXoeN1w05Cpgv6bFncFa+HKWwbGvBsrsQsmJ3u5e5IGX
ZkiuRZwdcfo1Ax/ovigObfC2Lbcptc0EldAq+/tO/HXBEaYlujfG8xfT7YtEXBEy
3tACiyLWtjQTaqtqAWia7j7lSKtHSWAYq9yAfpdv2zd0wkjv/yD+D3fJkim+/bLa
xKcKbGRu3qiJ59Cetf67Awi5sNK77HPu2wIhh6uvRDqCe137u+hMhMcgMg903i3H
4uexmBIEKDU9AjToJyWujQ0nq/RVPhMuSXBV4fqLtdvINJZNx6FUk0rE2eO7s67u
AKmxYG3Tbcr/pvoisbUmx8G6AnloEohMBp/Ga24OP2md+3YPCGHJukgZ6PEuH5kR
/DSMymecGgLBt8t8j6LYgacItf05uxA9lk7oIh8svWZ1ipOg++jPCLERDNiZGGfn
m1lRclnySy9bS8KS24Zm7ehB8AvsL84U9AdyMVaN2NrpN89zWOuwBoBeb3TL5KAI
8ievDqxbGl2XKK/d75ZGjQ8eqAVLmlxm2EpdEx2dFTuYgQ8Cg/rdymKMMx8bqRoR
laOwBJzGnyaU/jCkHeZggY0vfaPUhdXvAw/atI+XnA62qzmyRX954KGL2zEcZAYY
ZPtsegIeMwt5l8NBRpJW/IRlMBrL+mM3Eqv4ClOsqw0PUX8lMY6k0mZWjcXj0vJW
rs4qHOGNrXN8E+4XnXGUooN3tlJeZKeZw11ySHB/G1AZpZCR1+8fJd3ZUqe3cycO
7eZ+E7haBiP9VBxF8O2PvKFKh/TGIT6LjKRVAnVsZORwJ0S/6cSMmx+jU73qXvQn
8H34TtXaT7j34+u/V5jMVB2+0dqojXQ7RJX+YLSCd/2gooNyo7GXOcUm3ZakQlSr
eCSyujKn4f0/68r28+gMbXC08sNVEOyufX4yyYh3M92FTd8eosPumce3f4T3HhIQ
wuV8OTMdk+pYLABNUIWxzjYf45wnpy+/sLp8QF9fpWoLJr0wvtS3PLk5Dr69njlE
ILV1rtMRwgRbDTL/GrCSy8+TFcPWzfZ1k9yxY/qJa19ZjNMek2BL7+fpE3sM7sSG
oua82Z/EVzhcdVzLIimwNIYJ2zwBJuNSEk2NZx/HMiHehgS0XQPqJorr+7Ugew50
utZxLKV+N1AyfZrStrGGpKPyA+os3oz6ExxJQmU13fwJORwORuSdstouuErrBLFv
ggmQ05OgYW4qZjZ2fQjVJXn9skDOYBcKwP3EDB9p6a0bKq8WDeHLW9fMBWJYE2W0
gcCFGCPS0kiJCdhrAlOfF06RSZhe9JnzTxiFfk0kRB93CERTho+M7izeHksOWR+H
OpnTYTrppHMfWHFrKwA9OuSfGrVrPAJ8qdMD4d6w2RTHYCj2ZsMzQmyXWVaKA+mk
JM22OoHd5k7S+x72AIv+pZoyDQvH8dmelmCG4iy1P2GGq/0DtRuJNQP4mZ2Y0HUq
rPNx5yDFQCOmduLMPuY+VxYFSIGLam+SP7NQWLNwHe+tVlFwb9JsHYBEFP75Gj8c
O6iDkrxOH13NoFbdypNjTXu4qyUzfKjnMEVfKp6stVy56xO1+AbXFEwkF+Sr5qul
Slt60o0+8YxgrN7KmmNcdfdirSY/oYfPVnsGwsh+n8ntVeM+I192XAMeop4NgUBo
BGbT/9h7uM2ItbUV9lo81gH0tL1eicXsOSeOlIB68Q/ZbJV3+hu/78QFQwEMvHP5
4Yrao1UQMahFV/62iY/QvqT4abypOxNrIZoLMYhd0HR2b6ag5k0jX3BvnDNeSInB
9Fa8U042W1ALnYzGdj0HgC6N6yOAw7rABnBfyYS3tenq8WrgnnKDPze8dsAMKKm2
opgqrw/yv5FWHgJfZwD8EZauIxBIRXFcECPKsARPJhm41UaJASeq8E/1tGdLWRg4
gE/xfjCUJPs0FAbSE5xSz1iGn9aOV6Qn2Cn79vQNfUW+vB9Ml+N05M8+h+VEArik
BWrGKT/fYauQL1xMgOxVeTJyW6FsIQPrastMgaOcGSW6MW1jMcfHAUEx7yYIxKTd
MxeoKNAtuB4sGum0R5eQc156qyRRlprriePQgw5UL4kmMC3oJUY6sH1bPYvKrudm
efZY+zkGyGgKax0kwtrPnz8HGPV6uM51raE59D7Pe+ymHni1B5QiuHcdrTrY2GnN
LX9O4IQXi9yy4fR020H9twH+jeIcLVQ3ZiLdSvWnCHvwUfqd38mBuhQzZy4zn1Jp
+EwRtQ/HfvN1fTaOFdklskov6IS08E0D93pg2mgCO2h1jEml1xGmapAIK3JmdXb+
F1fY1B8ydj1KRnqyCLY1g5eEeazv3XZlxevnd5sLmR1mwNCmNav1XMvgR6Url94L
KYSvmsffSbLT2b7fF4lWduEyRuKNRA7ZczM5+ZRWGxZN1aSFK3U3cYU7j4F/8X99
IsyLRln1MdxRM1JlUcyl9sksjnnYb3m2zc2vJxe4Aa8xMmhE9pWr2DabYhOpNpv0
fN9uQ4a2Dylgv9EInRUJ3PRGsV+0VaeK5f0oRBquYbW4GZrb0E+02Ra32CJiE8kP
xiCv+ROGxlJvjpQMSW7NKap5NtiBn0JfGmjWbOFCGd/L7v+5l7xaAMy+DgkkJw1O
UIv8/toW+zMJCrkEFHldhxGcmyYXwCzQfUiAi1mJ5uHTKKlDDORkgiGZAnuMnBqf
Q3DYbUP9Qv21wgGe6ljQpj+Jd+8VII+zYdh5bhA9tyuZ+kks5k666FuAh1gT8lvB
IeJHjQlGi6/nheyCUAk/m0EFKixGDKtAxBkorTb5oCI1BpNGTHr5znoN6XDSijFU
7Wd/jkUs7mWB4yB9dNT/gSUhM2lz5Jz4USwpOYUDEi4o/l61g0cAaTIMAf5Q/j+C
9Ls5AfFYoxDZWdT7yfjjf87pRrCWYqbDAxbm8LsNnfIr9tZbKC0jgQPOmOkkBLE6
VpmN9aXSFbgAze8bPbCvSXDjkillIkqGZEbk1VkUKLaluKd0u5kMl703xKIKDhZU
bokYYkWGgiiGvcPuaNX7/6LvMk6gTvguMGqXno0Jhc6l5IdWzthgajOfRm1h+nKZ
OaJcUF/7O4o5Q5Cy05eE9gT+RMgeCkr/n6hZeKJAiZ8cvSo4DGawQP7g2fpJ1Xbp
FmjGLoMqETjK7YccK1TTbDvAJwj6qVo+CZb/KXG5i+dPICAQKHOkjt3NHqHVdvQ9
F7boEzpGnUg44sm54qWFM45KJz61eRJZTFUZzdvn8Fem5DeRgMHO0YnWh8kR3L7W
wgu9dAaQ6aBqWEWLCMK/xhFoCi0GhDbdBUiRzJA1oJ7czCF2gf8rLHBKbmZPaKoT
mn9+g6OdJsWgdQ28R7ffunLp9GRyRixI5xBpwt5R+Ps4vnVm5dmevhA5Jw+qqnNv
zdVTaeMHX54GyLSu0FAyUCRG860hqJIYv2UHkgxNc8uRB+NtwPAVKUAUUUmbTWhe
9GNjQpP0L8v3TyRTBu7hvgTCz3a/usZ1bUwb5mk6NN4HXn3Ex/VXAovBKUHjhXxB
zEEYCqFqAKk5n9N8z0niJJHRxBDslTz83VByu86fDVOeDH/cl/hAdiU6jj2Y12WZ
fnWrwbFvDYGlA8EAK3EwMWBaoEYbEx66IhgAOoS51TtKjytQwLo+pQCMrVkOOH89
5KDMf1aLgkV5NldM7KxUDYKDWoNkQ1ycbB7V7nA2RsXzAW07M+AJeV8GWp37V9by
QK7fUtTumLdAeCYNner3I3UvldPPaDYGTi4Pa/i2t3vX5IxaoMqw6ztpiYzavdTw
zr79ilZ98UPItruJz4PTLF41zIvbEzoKeozS/zEIrx3K7pTsCyS3v7TFX0zLhJXN
38L/2Tkzeq4LFt85I1yf0i57XkBtb9oCynDMv+dN5KX1gtnNDeqVqJYXsjv1GeTD
Gz3UKiOrGQos/TKIWQDQ4Fwq7jhaory846+WZ92r8O5bGK6z8YUwu6y+ZzPqeT6I
3QWEyZx/SmvRwex+Frz0868ZjlgAZp5i7hwdOHXLE1N+PkQAkOpo6Dus98neE7aT
uHdKpCtT1t5E9e+JtgSm8XgdoIJC+wV29HLE3pwDw4Mb7V5TwRd+UEMj4N6soU8t
ciMEHIk/Qgu0WvqEmtLj0XhjVuBaJQBxa735l/hIG9fqkPxfgiOE6ZBg+d4c1AHy
IV1LKUmtfaXYZThhxFxH0AMzTkN21/GbvgNbbKs77UmV/B9euEtr+MnjJ97wgdeP
hvy87s79E7agDNzXbw0KgLsvC0/STxOUnPMl8iQOvI9MJ1ywAVu6jGLAAT1LQYRV
tuR6Zqfsabmq73M34gxntoxX2EgxCTH0TLZuyZGfHJrlb7grjqRf6bgzfumZC6xf
/oICq06K6irW8U4W1jlGeTY91yalegVg+2HqXYV4vyzs9PqnvHZq97g1PTWzYElr
1HK3NnmX86sP5/fFgXxbAaFZixSmp7D4JQtVC0Tz7XWHfrsj5tywhN6BylnaYD19
1HWnhGImkNOQx9otrej4czOOPTk9Onzxwqg3vB9g+5QjAAFwavKa6FrVuPWpasS/
/gJh0lRtgeJ6mBUsy9H/WYRLFGBjBnWoqFwj7UPQx+hSbvyKCspLEqEE7KxBCz6v
UMUhdHqfzu5OB8TowricLPts+IYZ1f4zFKsj3DxLhlPeOwK9Z+zeEbTWYYTni2/G
PRzL0pjzuFtmzOKoYYIi7sbAsM3acsQrY2sPdbe51rsiQWqx6FHSeDmdXFtU97g9
grHdD8x2yMqJDgA5crBMmW2YLyVx7YpcltYa58zZFo4F1XW7j+svR0uHDBGuCnNL
r08GJMXYpFVW1RkmBMFWvZ20jwdgifQifXUEvOkG//CNGMkTmIjsqnn++oWWHj4s
ZrVYuemdvGPiNdy/Qwt/2BFtP5/u/0M3NmtnjGarQpgrW4gMTDlkkuZs8eOQ1CKP
izgDnfg//H1EETUwZYmaqc5G66nWQdjBH/i5il5TwQHgOuw7FQt2te1jv1q4M8Cy
+yplAcXg6jBUA808aLdbz/KEVXrptW/cpH1DRD0m7dPudiMUe7brcDUshRg864Hk
kpx28goG61pvkz4zM0Y5Qq0hK6X3ITXS/T6P0PcofkZ7QNB21xkQ+2ELCDpYe0sX
ZuqBsO1fycEinGNtZGFaoVEnAl+Y83oOM6v3qzw5qFrGuBjet0iFyK1b7sFOUadM
Ytnl8Mu/yzVACTK2xbUNMacrX3H2XDJg1WV+DOnaL7AwCVzBEHcyQG9GB+9HsNQJ
YCGqe8k4ZKnvxJZSJjcGsBTJScYs3gJ0jHxAQFbvvnV3Cp5i5Laj5eDlYaoK2SQ0
vh17+goAXEy5s8HSs5yGwmNkoVQJH3gxRlQ1rwPunaVA/jDF2gvq5sSl2cHJZaZ3
8Oj/OFrpdGs9Mi1GHL4YDZUwzroeNJF7qeKdhkqgHP3MHQ13FgYUqEaYr5wscbCs
MenqLBOgSb5huqvuraLK+odUuWUdenPXuE8Gfe+yMRXpvcibBaKPOB9NlAQdhSdl
ydlN+1HurhtFLUNH8qGO5BbtVAtNvpUSAxWN5k0m6qwuxHHugoNnk66/d4p9yNRL
EYiiRiVnJyuQUncr57S50A81EgkPBj72fTXQl207hAvxYctFR4Fh4j2fEfs24sbt
ChTFaS7Gm1oQ5+NYX/axr+7vWEzRkgCXk2HaQmvvcNohaNKjW7GICMVYX8X61zYI
UE1za/XozC0W/wQKJ9oYGER7f4lh8o0rc7Xl5h2MpvyoDustK4Kb3pd693+KGs1u
5rttxbNp6pz2hdoQYyHIC5XsIleTWqAWRq4J5Dd/Z8NTBSJniiQ20xETrBWb9HvM
6kme27cm6Ig1BlSSYJurlSHsuTOJZ8v+jmPlYBEHQYYfpis+25JJnefxosmjPxO2
2KsVW+VxzHf2rlFHjbNYyyVApjmYUkCotDZMqMp9xZJBck0nQFuWIYGLfH0mY03p
QxULuC0UsdWjTlaoiQjz7M6b+IHPneWHhiqXT4QZjrIREwXG6F8BWoxm2el5gCA8
+BrgRDAd3PT4+pLDgAFDAABHwQ8r1ERs+kZL/lJCaX1JyD1UH1ebiv0x6BlEC00B
XSHALuLCiEjplO/oCwJ4CfvfK/PoTY1JWt610TnKoWi3qglQDJb6K9QHQGGtRuih
N9HRNQITYeI6W7H5oCeXCGk6yTRzjdR53dHnXcI67LtQK9lD67QLwuygDRFP0nn2
dB722EgE0pRZren+dv7qDjxpBHmd8wZ5puZ2L+pEBJBilN4gjYHPkwwEIaZ/PQPG
KXo4fskdGGMPFGMDobxLgMTqfYai6QKjjX9F3xfktZFqEgRmNzsejJOct4v5SQ0Q
SSMZf1oJO7UGYqbfkeapFESdl6hKF/1i30fIBQBnw7GnesuavwYuhYGKa5ZEfUto
5As3o+YGuKSVTq8nb/WWHi3HAbxndOlYqZseVacIrqtTLbDVeAteRHVY1ZR87LA/
6ZLlfYGFLJZ619c0Y6ylAcAuREN6rLh+4BOv45OpnatCTCu3MNvQjFgtTx867l3F
TMIg3vK0kSplLmEWaxOvMCnKxAzP8dTkWhmoT4jwTuo++KhS//d9vqmuJuWlTJZI
dR/O/X6K0SyQ/QTlpoCvgOpUlTDiLRr7kbUW1cNrIV2mUMAnkaYR2ANYoUWFfZep
qAx9M2Q0lgkBiWs990SOZOwsrEaYsDfG/DAXxIFoQwkADz2zt//e7JDWZxYa87iC
M5+hQ7rHCO218bUXwsBU0rhjeZt5w5qjId+CMyjQ2Av16+dd8S0/6nwwpcxLc6H5
byhLoWN13reSm76ivxWCTDZcubXTk9nihQPINbj0uL/OzccJoDAsh8J2ECp2Ovap
dz0qFX8nFz8ZIt1LluPvFsVztv/B57vI/x0PeFJcOp6NYnWByBcwRdYURdgp35L+
T2Rz0t5R/bMjzh3Dvt+Y+A7aI8ZAqr4OB4XOlFlcXT6Jjc/Q9aIT9uF4I9qvvi+a
zMErbNmfm+ySW6CVHUvbaAOCbpl5tnMkwQs0TEHwCLicnCqnWrzO7YVaRFAAccgA
L2KKClvy+e8XYNZCBYvo577a86sL/XmnJuOVYAshWu721GDHn287rcxrSKYFpD1e
BMQh0mc9rP18QKa+APd0kETT+Cr1tq8EzkW7DJW1/iG9p43+fXtjw1B8mUxaZokO
mzKonPho8J431AnVeIbaRSWNe1KgjzteJBa+9pIqJP90YGMhPbLY8uTuwpFXoOif
UwR3vfBH2s7E+6V63sKsa/Oyf/cycZFoTDqKIENeF6/0x5cb46sEsQj5/N0l20D/
oMbY3QB6zJEj6gpdCDYJ+m8v61fxSwW/yw3iVeyF6375aWMechLKfmIzZgzfzHAU
MonAFOWhphLscnqWGq7r68Fky1F/HLkxPTwQyaqUXOyTaYiAsiHlWWy1B5T403+x
Gia6+o5BEYvvdqxwDmW9F4pwCF79bT49dE6B76yY5kyMacB1dt3bQ9VsxboZrPu7
vd4cUtYGtTTCDkeInh27d3CC+ErRKbWRzZgTcK4yiD7AU6pGwUydU4BRyaKVCWqB
JVudPQVHKN2EqSGDPkPVtU85ytpN+YBN/vV4mYhOyWE/phh4sZGcZH1uCamvDhqM
MVQaqS048KGyWXs1WrlG7c/jWeuujLDNSCQtF71aC4u32Dg7mHGi7A3TSXxzW1Cd
cRlPKtKP7nAs1c7xpJudk+BvICqylEQhTFVW0jMnWeA3ZImkEU5pB49vglsuSlXJ
X/0IiQtTodP56SXY4Eu98vrqhp0FtoYFUKqLnd8qCvAuZXOjUVAaPgSBF2gTwdBw
WPrSqeVkk8GCHKzX5Qp19cUEJVRKuirPqyOU4b0vkGN9Xd8J3owTetFT3SgzUaCJ
eXlDE4mAri0WzocKKWU6KMbW/1Q25X3NoP8DYp1tz4nLiTWPYFNQl5uCYBLcV5lI
wMiaKL0ZJ0fiVN9r6Ig184IMedCSBlestoDgCM5RRKqNfmemYT2A42co1pneUmym
wiMe8f3vdQ7MrsMiz7A/tiUgUL+WYa0TrGC2zrfRJrD6JOfaywOAjYzrpUPzL5h0
9bnK0sk3qB8EeRuIMJQz7nxPKTv8sevAdfy12Zv1IYBv9fb6M9jHWNNKLwbpcucc
3vap3PZB+JGYNNhOCsLuw5JFUnONOyv7I5sfL/QtAirRRmeTy4dOkIOVeXxWFh5c
BNYgLumHQNWfK5WKMRsMeiuwyk30/UQ0g8FmcisC/MPY56CHJ1v6bPXf+qZDu/Hy
iya7EURObvYg1SxQVzhK0WBKKm+3rTM8R3wJEMVgziMyQYv5FVIBflmP1KJXqPBd
RVuaMOCmaMRLGSRhc5laPmkqeId8Jf8jnuoCReEJ3ft2k0OdtqfFsyfEHu7TATNq
ggOp6mu9aldU98KPcUThwggy4Zb4tOF1DwwZNJEQAOVED9gX5glajpGwMzJvTD70
jwV1j/8Mx0wNIJMRSzY/whrSPgQmhm6aDX+vsCW2TCkuDBN8lG1l2O1WS42kZBw8
e4nR+O9Gvvts5pnmTzMUhul1fydS8yPvaizhN8wdiIvUCqohihvZ5u4vL5eg8yQN
HM8f4sruO+/vwl9otc6P/SeaKbHsjjPfagOn8mJZykJ0FiBZB+mrd+55gwYBn5sJ
kCxWubInLscEIM/f0DCX4/MEA3EQuZcKiw3ZSD4WklT7w6pugyX+y2Da2ROCbwMx
IzzRs6yLB5W7mfNbRX5bRcdQz9jRCF18TEk7sxRyX2zy2Bkl6FQ3Oi8LJ2xNeLFq
AXuC9oz/LFh8t4rYywKaXzjy/CmcalESPW3vt+MRXdbsg6ZYyB5MTstvp4fIkigv
vthJbHiperF/EWEXxezXl1dvuSbYIXZzGlbLszSX4Mqk3iVkezPJxC05hlOTcOv7
0Sdc+xzvEeUlNnnUui7wJsaoyUO20sDXCS+7m97K7HpUyge4YfmzLanUfubAXC15
+/hIWjBrWiVd7ucWVNOyVVDdEEXMAo84ffN9C3DjAJF3vSWH2YUlJRcYTlv5PCxd
LKHJLxOLw11zcqqTHBJjFEXj52LHGTirRCm/Y/IaWS/HUrZ0UGDkTLDE9Ma5jTis
qKP3d4L+N+8yXa9rZsjAYuPxU/eqK7KnvCmiaKLdGnc594WPaCjyvpejsasDr2a2
8EtYQ1K7DdygaTOsgjjY1Y9zMOQncOQhXh41UMfbM9wWK8VuG+PDAdtQTCDLP7RO
gzWRdKDbnKWuxAzFFx2COJqwgP5nu293dpGp57emnz5ssfxL5QMq0w+HwMoFJIVB
LaHc/maqQ+UUO3oijN9QXsMfdWEUrh9X+tfvx9ndHqMTKoxR9hRDdMsaX62aYQHT
gMDUlLnOHd6VmS165B2EanD0zbHhuNAnofUUkA9XDQNR2lms7N6fcOrS8MT8/y8L
dnrLDJh8pFyKguBgIIyjBrgvjSCwmxu4Rql0Vep5iW9tbh7cgR2FgHWIiApKIJTJ
Dbrh28ZEvp6vm8sMjgvZxobSZgbma6a9R7h7lNAZtOZzc4Z1lx9o9PPsQJ2itZXQ
O+MjMLhr9OhgL4DLpdyiR5sSLYnPLqkWXRxeVTzew2IVtC+owgrdi/fRkVqx1JFH
ez9NqhCXhHkRi5fa8SJq9ds0JbqxCaZbHt0WHa6jCkMqUSc2rqtK5Xb3uk1IQCN8
EMtp7A3uRAHSww/sfe1GZFXy04NkbsaJtp6InSc94MrtCFQHN3HooeRwExhvyLBz
A8+3P84Y7vBrZ0RZ7XLAWa/sX7SvhkJjN78iEYo624+/Nj546nrX5pn6k2M+qMlp
C3MMnh/etkjucHaUDZugereN+z1t20L6w92Lb94UewVkI27ppGG8XPZPpS/M4aol
+NTgyz5TVQPzdFkES8gA+jgV5pc3jYrHLlw0xBEkgw+9+DgkOhS65eYdAQrod1HH
szMAAxJXEPEecPM0y0rcVI+HUPL9YeSsi84nAVZ/D5jyvNj084h0VrPbIR7nxc/8
zcvDHRSif9Goi+plUn3THd9cAZVPUT0cQzbTFQRZL2A822SleQdcCex6lnHDe8Fv
J+Wlt7ed1QdYvan5yfkxtXV5JO3Otkb/t337shAxdHFD+nGqaLMoxsyvQnrQV2WW
uELwpYWAN+z6KjZX1pAaBNlV0foLr59WPNJNvKX9SaiIvQdJ0BHy6WOIKW3r2diW
H4VlwbmxNVysSkHFiqUc62ibxfR3zduZPAe8Y9hg68RaLDcrhUNtOnDPzhgsYdw6
+VZq7cUNN6PD9i7XeohwidsI55sv0r3zKuWixakyMw3x5FjA3LHwX42urC8bNSbz
b50KdRxnnF6VDz8M5K+QoOduQ9zhDIlA1Az1L1Hd2LeUPEI8sCpcAwZJocOfrS/3
tKvWIQimkcUwldFJUvnXZQh1XSuXusn7Toim8qJzEKfQ2tHuB8m6NR2jo6SpKKef
jjyqdcY6SPvo7NYvWFnazdUyaCi+pWTIcd/HG7XbTCR3NlbJLI+/gNt6zEJL1Fiv
e++ITQPgKLf/K1RMSsP5xgegBvj+pH2Xigqqpy2DMmxohcaMQ3jZGSxPAii/D2ND
LQcSjnwS2zwy7azHnNTtE52Ud3QW6+Ra0TYJQR7oL0smjRZBL4XWGHihQHckQXMv
KbU/aKXCQGIzSpAgE4fgIfLwLtTQ1LUCwk1bpgy1Wd+eJNRqN1s2oEvFtYsnlIZF
Mm9P6MKr//qRxrDkc5F2xujXYXoJCGSBZaXeR6NAyk0nUDxEWH2GMh97oDoGI8CB
ZjvVUztPzD/V7G9h7Ehf+Q7/+xV0cqKkVydk9DBbj5dmpRttCBwIkBX17zPhSMwE
dKsom/1zPoYfU6uR0oqyyWXsoW2MCQr63Kba3IhmQTTVLnVG+J5QqTrAR+m414dR
e0exEa58MCciyqb4Et6mWpEk8/MZw67HbLD060o57wzJQ5AZut0fL7n6KPcj2bQI
rcU07R+bu9i7DxG51A8JaP3FW7SLqBo4CFgasH8g1wNAIKP7s0uJzTwqwBfE1OjE
aKvzDd8UiTqbl0YpkYZvWf/QM7g7vstZWpqfjb3l582u8erBtu2szcxwmW5YIhtq
lJAYEb/F2wVxuVo9jF/ZXIYh6AyVEDEnHFzzznlqaezldLGcDnTuunImdd5fiN/Q
U/e7LO3a3zipM8BSJeRFxIbRBTKKTI3T+uTpgnDzvDuGw5XH08jYnDhoaO6xgaPn
M3phOY1gLI1hGUY+2AZzAyITptCXS3ZqRSWM3pkd6hbIrnr6G/j5dZJSrqxuMPa1
HqgCvRrh4+dQO0Dn+VuSG+EZhTUDx8tQ3dZS9gij+nAV1W8X0ZyZrsUh8uRHIbqh
BjF5FBGBoyCN+snY7I89udtexNMFna3ggK/JlMxh9tUVcKssdnZXs8FEgm7a5pgU
+rexTHdfHBagswS7/uicVEhQgN8zFyWzlsZsFZ7eKJFVuvde5ZQnBFXa4Nv8gsw2
upIzKQhO52I69z+Lahk1ASxi9sYfBGn0+748IUpmRHB1afjoeQ/4w6lyQi8N3FiD
/nANlmZS6DM6IHQLOAPEyzMz2NLHFqOE1S00uURFMPQf81fM4s4LKN/nwCylXI96
nM/DPedB6dXfodbKFiBGxUvTP5ugO+OBiNXl2fg063LvbjWhWqPn6xpUTbpkfOwK
ByNoDOcEBnEArE7AbPtjPI3oUrRanhsV0yB5HbV+RYABYS8lx1ZBa8GKX3wDQkd9
kqVUfrGep5z/GQnG8Z24kh2J0q+nEYVxvqDgW4qacq4zQxUVnv1CymIbZoxqzByS
nruyjC5v5JyA3h/SKdIgmkfihFaO6/oJtCwUnOSMIbVclfC8TFbHrRvPEWNDldAv
iik4Yy04fZhkdn9lu14tZSRSKsR2uxw3BoZDt1EXrw7JiQG9OTiUJvT2BLEQLo7F
L4iNUO+o8eue6LChPcqTPOVWWC8XmvE+1JMLaSToNoLSsAC4Bm9OR1OtmQRF78rL
Qjdy8C2SZOxysU2N0meg9Jlw2ZNNqX/Q+hCeFlg2hhQOC7bVlphv5ApLwjQmhr1z
XDnh6aIVItOVXAFnk8EWYBVUHak0QsbmlgNApUE9peoa44BOTqsTsQhozc/R/UXA
3MsRLVTYhuOEelN8T6gXbms5esKDeSm6ZcZyfJYUrsC0jZcCXh3IelOgrK4vK9TZ
WzgPyNiRUfpwjVvrwd3u2sd0xHts6Kc7yS2nmrJ6cK5KIomrW7tFEsgfEZIrKpXS
E8vwqvLdJDS15Vr/F4apJWqpHyV3PGvcVtxzweCySWtMIKIDfBjamHiF6IbAcNMI
asjxKWihMLkfPewNXGl12xC/TDVIsRQzMg+RbMlxixqGvG1hKo7B5rZfFsPE/S2Q
fGJLbUA8GmnTFnBT4lgP0zWram3Ta9qkc/e6yjRYWkYCjuoi3kTbOEEGVBI9CmGY
xLEH8ssSklO+HhNfbva53Lzbq4Wa7kWkp7uzjCSBglsD8JJ5vulr6YIK+u3ZgO6C
zleh85m7z+RPCMLIkE6xVH4wyITfJexjUs8LG18sxz894G1H+RG9wKNQpr5FlvkJ
j+TEMWo7jQI4pSF1wTDT0LrTRUOqJzZymiGHX/9QHSImPJ/MXcTlXY8ybv84rpBA
pNEqZ2MfCbwEeeTUdqqQk3p39bSlrH3W8f0bMO4etD5aic1/4cFKskupFvWu9XHY
Uxdktu2Tmlh+Zvj1g5NdgDW2HNQyde4OYUva8UuXj0Cwn4JIqCe/OUGGhw+rI4Br
dbRtaXG1h5Jd1iM8lY06UADzE91j+jV0XJopkFz+j10zAdWgZK52xkfR+SJKl61W
5Cn8RNAgORUfOAWanpkxQfBN1k42AQZjPkJHWjRYVl1wbHNST9TlvGeypfiVZGEH
9PxijCVujjU7OXyPsKYJ6UAXj8E9gEAdq40l0IUJnRUTOhFcVuZ4zb45wzFb8rCT
rrryttWmH0ZywP6F550kUi13aBsMCjU9sLoyaU0CuS5JlbwovpG5NecdwvzDU0fL
TsJgTCgvY8ZNFsNOfcigmGG3wulIdVsIgCf10SVN3uefr6JloXaau1eTunPzTSkP
nIDLUOdn3uRR+6iO2VcvM4y9WaxjKQydM18VPRZmdW9MJrtGnbxwriz1vOX95nll
1SdDQs57k8Zq/R67fVcSba357pOWwK5J4t8ZljHFNF+HylaTTAyv5cBtb+KiNdwA
mqvnyT/qMlJCn1DXgkHeTWe2rwwGYVceri5dBcLmMvUrMp2m49Apmfav3dy3P6BV
AsNJH6dOO9XOJjYpJGcdfNuP83yh6oVoH7UdubUC16mQ5UbM8ysX3PmYMPl14YE1
5T1rezCICcVnHhU1vgr6pjiS3outx59krnAmUS0YE/psHkMKd33xYKvu/vfItXrl
w3SimQAWsevtndZ42oyivO005o5xIsHX/AWzxSQxOMXXADsZ1LmwkpuDe/fQ7pzR
Ohby/YeR9dn5bsYW+IJP1pvyTa+8pIvxiS1mOTOdyfKNy7HAqacbV8wby0nmpPD0
pLDP0V8bUCw4LDo/LIUjTFycHPifYh2MjvpJfPqtZWUlrJGoPolnpbXobGBxVUiq
BrnhwpfUdYPmDmZ2nvEgl8P3wg/vuJLfUZdARH5sKQIy7GG7166b3Cpbn1gEC9XR
ef5r9mid7UBJoCiJCqxgNa2AdZSohOVEl4D3x4NB/4H7PX7lIscRJAgc+ZGo+k6c
UMuWbrtfnjuVCQ1ApZQlnp06AilFBQbg1KT+h2tq9ls2vaL2iCLmBRfaR8WRlfpB
mSmJe7qMuq0DJ9KO0/pe1k/GSlBi2pJvMxBJkVrxXgrFUBp7DIUL/N0Rnorq4u2h
+CN6z2qZF0nqjkrUGRZn0/r5qaXuI4tUg9SB0+VypbXfA3yQgZC7s28qEAWzenla
ENufJS5b6IbYhnv84sOIoR/0dFzpHs2JZdyF0mVRlc+sjkA6osdTOSRGxHZfUo3c
x5HUleiM8qvWeQArbvUfoTyF/HkSEOBA+xZMhR9Az5MjvaPGQNj2x95fzUmaLK/i
I549JJr+4wgeOizrlkHCxTR7Rd63wYhMjn/5FkNnlgkASNqQeWelqdlfy3NRT97c
VwLXqCJ/CGZV75C4zhxAxwUiTFLXt5x3Dp8UAZnIzlOSHfRe5cNwyOlmhslA9ao3
DA4puQHKRWw3wJmcL8Bi8eXdorQiVpqq1gEkR8zJTmIa4KfZu/8uf9yEgiOBXqCq
2AsKVNGtE7PlJFv8rbKueP6FMm1qYFmtHAD5EGaFhLHjPLlSHRENcBUc9RNSMtS1
FvIe+V6BtJg88neLH2ZgPY2htUHJ7+xN7oo5nl1MLUWgfqXkYhPpfvDb1U6a3Tu/
gtSNqGvwQYbF5djnK+M86lpsqnV/GXc4GV+5lwcrecLq6syw86cXjvbLxg6Wmq2X
Qv56L+s9a0ODlSD3QSUb1uXNZsG0elESo43uUOOLmkC9R1YmqiuQmexfJVBZ/t2e
Ie/lnkTXAyDrAcN8PYCt68w9J2QeQpNFkigRfWxjbFSj4ByaqO0u7nJ3r53GRwCB
On8Rv/pyyxsCW+OmQVodYsWxkunfrjz1Sqi0kDwA5r6Q6ZkKc/PyZH/Dt+rCp6ki
EjL+C2XXGxRNVbFFVJqZWQrdeF6yy2Ng8uVOHIlwKGDjZB4PveYgwpXiQabwFKrC
Nx3G5ZqqsusWTy7bvw1mYaKEbkOB+uMG5CXzJEojBMHdN879ORn010S3mxGAE0fg
i3QQBJbdzObHq/svA74EjLD3WUDBt59OSkM/dEdqr7vx7+2vObLI+s46GtwqMl9n
SvYlEIqnH3Km1N8mJMLjH3BjyUKYjHJCVZGR4gxrUouT70BqXxNj1Wa1NW24ufgt
VonFbv3/3Hkz/Fz8LTLhDALweib31CvRhVPiuj7FSreiiveekSiTn9cFBDXuhzO4
xzzYkCOOIK/YXo+p2ptlMDPMlO+bHd1ju7bIEa69wZ91Jq52FHkK8aBy5vqyL5zG
duJIh1FSY5ZbzjqWQx5ZDTR6Ch0i5i3xZE9Y61b+Llx8ePiKYWWMEx45vfeThFhE
Xqnclys+QDVwU0ObiCNim/u5uN3Nx1EomD9PKaoLkCgwzFCy8q17C74E1Kp2OzG6
UXC0CmeGCS6tvvE+7rwFdlSGtTD9bl+Hz/9noGyDmPtdw7o+61SlolkHQ9O+vOqB
lftcP6z4FjasV7n+7X5MXs789dZyJF52cMTT9ogo1uU7tniqRhx8a+VmBDqj27JC
Qmz+6vgodR9vzibXOJtFYIViesGFCXtr5bs9Vxlhp+5Wariv8gNhNaGM+g6xAHix
szQbLkmSr8O558niVaZz4ntRamQjtFzxHhrO4SuNq9lIP6kjEh8AAyZBDi+wbrr+
zNZB6ZEgNJRKdj7xWXPUH+AIvGAA4w8AizwqKb8g1VP9tnWUyR4JTAKry+VOpAno
oFWvud5DmfQ5v+2J3cnpoPo+hvMwb8YKC7qsBV06X9QXlX/XOP9WaG5eL4hD1MU6
nNNcWBotDW3gSCVc3FN/HliRB5TmU3jbVCA4/1KZoL0wOg08gyPCDYybEb0rLM7Q
FKpsTRR6vlT2FiJyRBh7KAXd2sZ6zjdX8gxti+KXcgGNhb+GH4L9xmLp4b4S/KR5
cBf3zhb3fnmJWpExfXAtvsWveKejYXLt/1+pYjaA9McDl9E2SWgM728dRAPm4+/s
+oDZTLdcWBZYEifxej29UkbDlH6NBUzu84rr1IVNBcbBiNkzfTcumyuLlLnpdtFi
j70BlDPEQhQfqeBaAgYL4odY/VYUyp0K6QFgNSR3eC+e13zLbwdTzox3LnE81SPW
ZdsqByjU+xKvYM+3uWWC2C/mSFm5/gPx+8SqnZLit4xG0RyqP+NJBBIgEY9IEWe4
nw/j4fcdZQlbkQeKscEiUEi0Je/5RKXsW8O2ahEPqxg16w+fiPa9/qIiESPqcPPa
iTVtCkr79ehzhgCOl97rNhvKP/KaKjvVBKfMoLxGg/iLEEs7QqMhr6i261jW8Kv2
xhPzrNYs8tiWweMLXfUIXXK0MgwnowBWZ7rNgO6xo8p73KjofKtVgPbGI/RYdS8g
bHrAH6EFMEKFaDbOx4LPXy0vJNKqvdzScgt0uxz5oxaeyZBD2lY9qn4ahxMKoRp0
pefa5E/n3B86jaUFgLHZI5bXY01EhF6fkXgZIbYBrARZ1UcecX7e/8+gqIFXg5rz
/QU66+BHjlPtksNxzNqs8thCti164j0n/o0cyuO2O0jUPmXk29ZaNhYw/VzL4AOE
FHulwEWuhEvCa7OED4+5fz8Br47ah8Oj6bfH3yGW5cZ0USfuKNz8aZQFzFlXfX8Z
O37qKxdBs8TtN8LAHgOpn90g51sidZvI2pe5VzmCY1jBS71+mT5tvPz6QGi8j2P8
SgJV9zbHl0fImvmXixQsWFtwDJtPeinluo6pec3FH5w/i6mZcQZcZ12hmyPNi9aO
l1++rFIfEt5BOpcrEXwlVybm3QVx8JG/Duhg3qcqtMXoObBj1hYNyAM0t2eF6q6r
OoOgCMUY92N72q+rFnZ5qqwO9hMaAG2hx1FmHQQj2tEllkbvNgPCurDaQhTrw2gx
94p8PcE/wnCDzbP8FHksqN/XV2rEtANTNZEAToQS4NFNZ1nxbfdxPMLoJZjgJK+O
tmrUYva/Cs9GsaecLFleQaNQ/Pnf4D+feCyzd6ekEvvw7Gzx0RdP7c0gxvPwdXRU
14qUK4ERFksDG866QRJHjhKKhDoWHfDBRkP/IMBkxpe3DHAyzva0GjU3VOLX5ahd
HAmpRkhLtR6HWQ8Krjvp6M67+gv+oXPSdoQYpSNX464kD5ov9pGHYsq4F3yvFp1r
t8B4ZoU9UQabVxAr3oObH5HHbpm8TWl0VBnWkLjddpYmLmVyfUMA2bm5PLJpj9k2
ECL+Z/3inf99XVpiFty5XnLqtRygU12Xl3aCHS/Q/9CcN0ayb4pFVQmVwHesqnto
bsbUyMX6h9HXq3rCLZ2UnFWzPyKtrKRDTsdmYGmSRFaKEE/Z7KGB/LCXnbrF51jR
6faRvb5M39OFkUsyx70b3gAI3TsYd54PaD0zq6Y3lWHhoEGltd6xVNa2qM6bDM56
GXRVoHtR2+/2aR894rvN/ujHrgukKmswmbnkVCSsBGbx8Q15xBg1LAS3Ew+WKmdj
d7jzBMHPZfH4GmSjZ2Jkwf+Jr9tl91Ju1w9yPlobcf0j14zKTwbXbAvvlew3D8qu
p4U9Lqewwv2pUmMDeRoGkdZ16xKCvyxvL+H/LrGSF+3gkKAo+cbm4txGrhZ5pPL2
CCJn27c6V0SRnWbyKxvB0OYSLLE6RfShl88P+rHEM+PF+PNz9FwD+VnzzZYvu/OK
ZaoIeA0X7iMpH7G79R4kVGorVixkvNIHFXnsJyc99YbjmYzEVtik0+aDTXKUhm9V
Igc9/459P1CXPygwgjxqTHk4qEFJld0pVaB7M3ZGFEHXRziEJbJEAvjEbl8QKx+Z
vFi3CXKEHifgXz+jpUYzVX/UWrvMvYwRnYUvT5E0TaNek1gumVkdWQwkpyd4Eq9M
0Q6I84cIuAku7w6YrpNXnNQdtIxuF6m5u2Uf+cOfNar6LOnb5iF1/j66z6mHLX7S
lra8aUoLgpXwaVUJI2uW0huJws50QjrBvUI0FpXcXe7nc/kkhRYojKkY9/muJ0Dn
jOrhixkmUfm7OmIxXv2lgtHlESGkgK6fmgKbkK7Ppo7V20LNt7xZs5slISnQtcul
1zok//+p4CdjU+7IxW+3R2Rx5uW3E331uaQLlYv8OPc7zwOyYJCBGSoQ1HQPZYJW
klkplumY/nYHgI0Lrhgk6rwxd2h1GZKqFyiiBGGM+35Otha5ZW7/WY/VdIMPQIDZ
j3LIlaldKcISTpW5LYFQ1Xb74YHALCEUGel8LK2uK6r6TbEI3anypb8quroe4IjL
kLCYP4khOmh+HQMo4+PUrJD8kuw0ro2vBPhOmzwtkW9in8K9ryh2q9GkytUsCcEP
yBAXTlsQ03xJuSrLqIOLSB9uG9OjTLb9PurcbNDHyoGNfUJh9ow8RIs8pbokBbdR
TxE2NL3Dh0Pkp7LUdP25NYkT34Awru61/e5R7MiO6iw2foQL+wFB1LvgW621TAAs
jVa8LxdGhpB6iCNjHGWiYpeJjgBr3iS+knVWePzLefPgYO61O/+tCdrWtNuswPFY
BGXn2CTD4M6DJtx3qou2WQtgd3iR7zKLrstegCJVGL2wydboBPewzwt7P72nwwC8
QZZMdUsz3B0eRYY5SBIpI7k/l1BrnP93KJggpMRsWTPp5y4iD+dlqJIOdZgqEAyd
g3UtPWo/0gSwD6GDhP+/9EhEote9koMOjAycRwyz++qeHGKoBJ6OpVDR71x3Q+CM
npXsLEyaw+junelsZN5RnsnE2vTsoYCQulbya8hAbjb3HTlEKk/OZDXgthhHDJob
J0107ewxEdy63s1xqcGPjCiaQzj3uq8wCT5Ra9nUa1gDeXThi2Sa16T33iM4na1f
yWvmpBmUkJSLT3V5tQXk1uyjsBT+J3SXkNessPeG48ncA0YHYLXpLAW+NWK2azs8
DlTb45J+1iWvmqz/sLtj1BYsV1ISdQgk27uLjEiymGFm3B7HgZWI4wKaxT0QXb/7
DhPPGXjCMMzaC+QJWCPyCYQdfH/rMvab4Pbr5vM50MRwXw/A6amwLJLKGV57VtkT
HwXvBjmCWrpbTlmGwYBTvM0X8WwedYLIoaEj1FOPbg3aFVjckbI7dnRi5ak7k1gx
ecZhbVL814UNbch168XSwQe33UK3gvu2QdrFjn6U/BtEqjdqm/T8g7bjsYNvnvvz
hqrsSSBKXNKbTjv0B3YSe8m7mICjELqFWsPY90NvqeP9GSV7YbCCKJXNNFE8Owxg
jZfzSAFkCOVMuyweKI3vINT1mLirFTJnsjePO7Tl/ju2NopSeiRN4MtCpt96AVPN
/knS8J6/U2usFs3WJ8kb5pDb3y43kxQUpvZxl7uFXQsBe86743+3/1x7m5qSqDaX
MIQH+lkxcPqP2LLEoDTK9DDLxgH0ERvWQW/Z8hX/tObyMUbnFKIys07DLiTahrUv
NA2206IUZtuNzDGota/t08hTx/gZwWQouBVBlMFJigvdLcMYZ2I8ymeC9hqCY6t0
kf2ghqo4tJZ1maWomX5w4CRFoHnic8VNyz7kt2NWaCN0nD8HUAw6d79kAGokefZI
iHrQwlLSO+p5jm5ZMRJdRUCW14AuLWKJX4RSby7Utlj/NpIIzVdlHKIz0KqocauK
eqTLO5pFpwu0tWpDemh/1tl1KVCoBvPzIjbKdwg/8XbiSwG7GVEVEHvRMOgQAvHK
65052COb5aLHbz/xSky1S4FnKEqHeIkI0HwM58t8LuPZQ59L69AAxfl18c3Q8aE9
ClVnKuE21jjR1itYJtpiOYr9Zsko3rk3NbfCGThtUSSaRRKINmTLDWy3mWD9O/68
7JtljFbwnjcP/nmsTKvd4+x8v4mFO3ns7XV10KdvL+Q61a7JLk0bdMNlXB0hUVeH
4SXEo6TnFadMMyxexJpzCZX45xMm6AVgPp7UfFtL4KBTX3beNM5tcYUCG19hAQjS
rWXg1WSsvepvAfbG1e/0yXrugR7/0EZdYXVvjfvByaUmF/vLYIBj49FpH4g2gvF1
h6FhtMHqFxBdRJqN1K1ass1IzMHzTD+OlhZYYxvunQsX1i3g125Vr1IKsD/WEkwf
zvmyXDzstSocSEnsru9C1yYWaq2mHukygwZIUzy5KFCdf0kHJEbFWBR/90owLycV
8aq/DWtoHW3wsrYWuMo2r9B3IGShJQaVteN9Vll//9EjDroZ9MmMJ1v7vi21Hkhq
o589DQCkfhh55Xy2LqD3sblNkWX7d+ugj7BOWi4Yt8TtC+HHArrYTuxo5s6Ypz9d
RRLs8EzRIvn7B/4mV34t2RaRqJyZ66kjSo5fqmCYpzQtyDXk2mdWfuCgfHCN/gpU
7txuARRsVeGzs1fAwujJTFY55E8eFc3YDUVDmjv5qppI+5Zx8NbMp1Q8bBBUEkL2
Z5IP3i7reA7yObyjQYm/LdTkcWP1xf7iALBVbI/X+3yIsg5t3L7XODuJ03B7SdHI
1sxsawaP9cj8DIZINXkzmFxKtUM9A26COxzn5rBxoEWXY/u3vLOhgZk+8p0NcCur
QMp8Rp9RWVbWPACPfSHIF+6v3N8W3KQUvKcHXKuT7HBbtlhR/w8g3h8ozs1b+oi+
+fKKwtqVH+4CcwzYyRQS2IYWjlDPI+gxAceuZ1sRpol/O/U62AdF5tPLONpPLJYM
tDPzpxtRBpzJa8DHzpauQEzKqdg2ao++Gop3ZUVB1cUil9/faDULu/CL2GrkF75P
+fuBDM7N/Dxt4RHDXc5SaJqoPiM9DPZGfU0m+wU+CvwfGubc9IKaaSrG+IidqZWU
GXwkH8FqiXZFkcY11iA+ezrsNsMXKhCglhAcs4L3aBVMb2K+otayPYdjkHN3CVPy
2P+y/I4mZfvIHLp1q2gYy2UIqq3+pa0ABzv+s7YxHf54z19SmPvoQP/WLsCen2G3
9+8Hn1es+KZf82pVa/9g0yjOFLY/0CUU+O2FyxPBJYUaWRn9tsTndnDoInxdWLMd
nxyyP4zbMSOT5H+nCLJAtgBFbi+Q7vRmnlyT78R2YUo6AoKNPXklsyI5NG/2w4aH
S3+0mSO11V0hVDAbRAoz8o/dRuUh5bO+S5gYQ+xZgWmXQB/k2tHQKVqHdJmXOLqZ
3KEUxnBSXh7cmIv7dtARgHP5M8b6uMoNsD0s6DiNgcpAEF49ByizkwxaJPrnZrmr
bTLvwek76IsFuNKpjXBpLZd15yr2xwEIPBjnlXaaQ1rQ9e+/UH6Q/Glh3qy3RVtc
aAzevKpBa4FY3wkAPeOls4o/GGfRlfQVmh/hPcTl4wMOcA4DY2IVL+1PuZg48kTM
/kNr5GyQZCEagW1HM4SVFvEjix28pxTB3KSOoGz2wAH9ozUMhYZHLhlpPgFbJprN
Bu1TQ52HSBt1ux+AL80+jz1bsnSgP2cqv4hS7jeCCw2wa3zj3pSkOCVySUC+V8b7
pvHalSGfLtExHetpmbjBwRrkyNshClyLbAuOzXEmgkHtsGre0+XedEiuOAfqWsgx
0f4kGnt5qEt6buZ7QhmvhB9WW/lNQecqIsuUeUbiqo6R9O3/GPrJZsUaSSaJjSKH
xdANT6Oc/qrIGbNG8DaMfoqoKPYVSB6gQaPfljWiUPfWOmpvHKR4XJLGQR9sl9HG
1dPE3UPoSdhY5IKIneb43mqGP0Jqjjcg31EUjWTayOD9gMcjmnZTFolut8VUIpMw
5YWUAOh6ex4utDBF7Hse1lbX0h+ur/mvmSNBolYsW1wmHRyud6RRWTjyiL+ayewR
+gHC8IophYGCteHmsBdPQXxH3BWg7b6dLli13iossgkfq24dPGxwdOj846hLB3m7
nsRpFr88BhYbtzJan1kPWtpWjwdOmQS62CRbG+ju0UgJRUcbJDrF4kPEjKtrwKu3
P2Nd2qgTDK6+bcnL07+uIIWDyaW47FWuw8L6QvJ8Nxs56slYc2mrbnAu2tGv5N8H
6Jom02IAunoCVIH+DbZo3mDOey1dxXu8cUs8NWiHs0budnrnekjes7FKkWlS47tX
ecKYcsm1PO612ERJjcukL5NITCPj15SSNoZzGBqDx9QvOyE/Nm6Vo6pSUxvw5hQS
8U1s97uwueAHXl6/0xFuUhzWTKx/1+sADcEPXjO1K01OaSQv95LIcwYrqLEDcdQh
JLZNuw4i0pVeTOzI4xyC+ulAmzrUb0/gq0q/yCYcbUs1QCionrGCQJB29cSUhyQc
G/kn5bERGdD9JgIVLhNzhVBI9QWmsqkVL4bD8giKCzoOUMUtpKS9Y2mNw05zzxmC
ta2XbaLWjT1rXkpPOB3z0nqI5C8tzg3BFd/WlUdhTsq2tgEnSivtFtJq/Wn6V95V
eRQIwKwVDoGrY6M1+PcI5hxApPwAhwh3wqfVYMQdgvUGyCykQx+4wr8J1kDwvV/e
EZzWnSA5amnsBz8Ay4ftjBlqnD96yMt7wnHUqYr0CHty4CdxUsJFnwmNAbnpiaQJ
rTPnC3K2Jq1m9C4HXPEpYa3h3MHpzZRDs6VwuVQQ3OSudH5bVtu5PpbEO1RFIofy
SW3HlffZPWbt/5U1Xsqs28vcO7APLABBGT4n9++Kk7eTuwPhRy0yojr5/t8Aze0O
`pragma protect end_protected

`endif

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Z3pj/uCVl1QVtWPsimFXr+d3/unvAJYD5c02ryt1qxyEWQWZhIU5v/dRBmHoWhbV
ARUyZsCob7aCYXIJYg7sABIWVOe1U2IhnbZvsp0jA6rF+6e3RzC9rpiVNfW4n8hJ
0/NGxvC8sqJqdt0QMxH8g3/LT/n27d/6y0Fo0mNX8SI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 50704     )
RyLpR6JAnNnXKjUyT0tQlJoYYbHKOSFzsDL3fwrA2LGwl+i4DBeMuw/6qIbvS6BE
w0fBqSJIB0SgFTjHaCzZC5fwxxTTa1lFeFm3XiXlGIqfkaEpsyDWH34xfIxGZqEA
`pragma protect end_protected
