//===============================================================
//Copyright (c): ALL rights reserved. 
//                                                                 
//  Create by:
//      Email:
//       Date:
//   Filename:
//Description: import package , include file and  declare object
//    Version:
//Last Change:
//                                                                 
//===============================================================
                                                                 
`ifndef CR_DEMO_DECLARE__SV
`define CR_DEMO_DECLARE__SV
//import *.pkg
//`includ "***.sv"
// cr_cpu_subenv             m_cpu_subenv    ;
// cr_pcie_subenv            m_pcie_subenv   ;
// cr_ddr_subenv             m_ddr_subenv    ;
// cr_dec_subenv             m_dec_subenv    ;
// cr_gmac_subenv            m_gmac_subenv   ;
// cr_etop_subenv            m_etop_subenv   ;
// rand ral_block_pcie_rgm   m_pcie_rgm      ;
// rand ral_lpddr_ctl_top    m_ctl_regmodel0 ;
// rand ral_lpddr_ctl_top    m_ctl_regmodel1 ;


`endif
