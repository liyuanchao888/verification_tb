`ifndef DUT_IF_SV
`define DUT_IF_SV
`timescale 1ns / 1ps
interface dut_if();
 
  logic                 clk  ;
  logic                 rst_n;
  logic         [11:0]  paddr;
  logic         [ 2:0]  pprot;
  logic                 psel;
  logic                 penable;
  logic                 pwrite;
  logic         [31:0]  pwdata;
  logic         [ 3:0]  pstrb;
  logic                 pready;
  logic         [31:0]  prdata;
  logic                 pslverr;
  logic                 reg_sys_rst_ext;
  logic         [15:0]  reg_lines_num_ext ;
  logic         [15:0]  reg_rows_num_ext;
  logic         [15:0]  reg_channels_num_ext ;
  logic         [15:0]  reg_filters_num_ext;
  logic         [ 7:0]  reg_layers_num_ext ;
  logic         [ 3:0]  reg_kh_ext;
  logic         [ 3:0]  reg_kw_ext;
  logic         [ 3:0]  reg_stride_h_ext;
  logic         [ 3:0]  reg_stride_w_ext;
  logic         [15:0]  reg_dilate_rate_ext;
  logic         [ 0:0]  reg_bias_en_ext;
  logic         [ 0:0]  reg_relu_a_en_ext;
  logic         [ 0:0]  reg_lrelu_a_en_ext ;
  logic         [ 0:0]  reg_relu_b_en_ext;
  logic         [ 0:0]  reg_lrelu_b_en_ext ;
  logic         [ 0:0]  reg_pool_a_en_ext;
  logic         [ 0:0]  reg_avg_pool_a_en_ext;
  logic         [ 0:0]  reg_pool_b_en_ext;
  logic         [ 0:0]  reg_avg_pool_b_en_ext;
  logic         [ 0:0]  reg_gap_en_ext;
  logic         [ 0:0]  reg_sc_en_ext;
  logic         [ 0:0]  reg_sc_add_en_ext;
  logic         [ 0:0]  reg_scut_mult;
  logic         [ 0:0]  reg_scut_add;
  logic         [ 0:0]  reg_scut_sub0;
  logic         [ 0:0]  reg_scut_sub1;
  logic         [ 0:0]  reg_in_bypass_en_ext;
  logic         [ 0:0]  reg_upsam_en_ext;
  logic         [31:0]  reg_upsam_input_size_ext ;
  logic                 reg_upsam_table_rw_ext;
  logic                 reg_upsam_table_rr_ext;
  logic         [ 3:0]  reg_op_ext;
  logic         [ 3:0]  reg_op_next_ext;
  logic         [15:0]  db_size_input_ext;
  logic         [31:0]  reg_relu_a_ratio;
  logic         [31:0]  reg_relu_a_A ;
  logic         [31:0]  reg_relu_a_B ;
  logic         [31:0]  reg_relu_a_C ;
  logic         [31:0]  reg_relu_a_D ;
  logic         [31:0]  reg_relu_b_ratio;
  logic         [31:0]  reg_relu_b_A ;
  logic         [31:0]  reg_relu_b_B ;
  logic         [31:0]  reg_relu_b_C ;
  logic         [31:0]  reg_relu_b_D ;
  logic         [7:0]   relu_a_zp;
  logic         [7:0]   relu_b_zp;
  logic         [15:0]  reg_gap_ratio;
  logic         [ 3:0]  pool_a_kernel;
  logic         [ 3:0]  pool_a_stride;
  logic         [23:0]  pool_a_ratio;
  logic         [ 3:0]  pool_a_div_nomal;
  logic         [ 3:0]  pool_a_div_pixel;
  logic         [ 3:0]  pool_a_div_line;
  logic         [ 3:0]  pool_a_div_last;
  logic         [ 2:0]  pool_a_pad_up;
  logic         [ 2:0]  pool_a_pad_down;
  logic         [ 2:0]  pool_a_pad_left;
  logic         [ 2:0]  pool_a_pad_right;
  logic                 pool_a_start_ext;
  logic                 pool_a_data_type_ext;
  logic         [2:0]   pool_a_cut_down_ext;
  logic         [2:0]   pool_a_cut_right_ext;
  logic         [8:0]   pool_a_result_line_ext;
  logic         [8:0]   pool_a_result_row_ext;
  logic                 pool_b_start_ext;
  logic                 pool_b_data_type_ext;
  logic         [2:0]   pool_b_cut_down_ext;
  logic         [2:0]   pool_b_cut_right_ext;
  logic         [8:0]   pool_b_result_line_ext;
  logic         [8:0]   pool_b_result_row_ext;
  logic         [ 3:0]  pool_b_kernel;
  logic         [ 3:0]  pool_b_stride;
  logic         [23:0]  pool_b_ratio;
  logic         [ 3:0]  pool_b_div_nomal;
  logic         [ 3:0]  pool_b_div_pixel;
  logic         [ 3:0]  pool_b_div_line;
  logic         [ 3:0]  pool_b_div_last;
  logic         [ 2:0]  pool_b_pad_up;
  logic         [ 2:0]  pool_b_pad_down;
  logic         [ 2:0]  pool_b_pad_left;
  logic         [ 2:0]  pool_b_pad_right;
  logic         [15:0]  reg_width_wrb_ext;
  logic         [15:0]  reg_height_wrb_ext;
  logic         [15:0]  db_group_ext;
  logic         [3:0]   db_pad_wra_left;
  logic         [3:0]   db_pad_wra_right;
  logic         [3:0]   db_pad_wra_up;
  logic         [3:0]   db_pad_wra_down;
  logic         [1:0]   db_rd_ram_sel;
  logic         [1:0]   db_wr_start_wra_ext;
  logic         [15:0]  db_addr_initial_wra_ext;
  logic         [0:0]   db_wr_finish_wra_ext;
  logic         [31:0]  db_i_cnt;
  logic         [31:0]  db_o_cnt;
  logic         [31:0]  db_sys_st;
  logic         [31:0]  db_width_wra_cnt;
  logic         [31:0]  db_height_wra_cnt;
  logic         [31:0]  db_channels_wra_cnt;
  logic         [31:0]  db_filters_wra_cnt;
  logic         [31:0]  coef_i_cnt;
  logic         [31:0]  coef_o_cnt;
  logic         [31:0]  coef_sys_st;
  logic                 cb_mux_en;
  logic                 cb_rd_mode;
  logic                 cb_update_coef;
  logic         [31:0]  cb_in_line_cnt ;
  logic         [31:0]  cb_in_row_cnt ;
  logic         [31:0]  cb_in_channel_cnt ;
  logic         [31:0]  cb_in_filter_cnt ;
  logic         [31:0]  cb_in_kw_cnt ;
  logic         [31:0]  cb_in_kh_cnt ;
  logic         [31:0]  cb_out_line_cnt ;
  logic         [31:0]  cb_out_row_cnt ;
  logic         [31:0]  cb_out_channel_cnt ;
  logic         [31:0]  cb_out_filter_cnt ;
  logic         [31:0]  cb_out_kh_cnt ;
  logic         [31:0]  cb_out_kw_cnt       ;
  logic         [31:0]  kn_i_cnt;
  logic         [31:0]  kn_o_cnt;
  logic         [31:0]  kn_sys_st;
  logic         [31:0]  quan_a_i_cnt;
  logic         [31:0]  quan_a_o_cnt;
  logic         [31:0]  quan_a_sys_st;
  logic         [31:0]  quan_a_m_val ;
  logic         [31:0]  quan_b_m_val ;
  logic         [7:0]   kn_zp_out;
  logic         [7:0]   quan_a_zp_out;
  logic         [7:0]   quan_b_zp_out;
  logic         [31:0]  relu_a_i_cnt;
  logic         [31:0]  relu_a_o_cnt;
  logic         [31:0]  relu_a_sys_st;
  logic         [31:0]  relu_b_i_cnt;
  logic         [31:0]  relu_b_o_cnt;
  logic         [31:0]  relu_b_sys_st;
  logic         [31:0]  upsam_i_cnt ;
  logic         [31:0]  upsam_o_cnt ;
  logic         [31:0]  upsam_sys_st ;
  logic         [31:0]  pool_a_i_cnt;
  logic         [31:0]  pool_a_o_cnt;
  logic         [31:0]  pool_a_sys_st;
  logic         [31:0]  gap_i_cnt;
  logic         [31:0]  gap_o_cnt;
  logic         [31:0]  gap_sys_st;
  logic         [31:0]  sc_i_cnt;
  logic         [31:0]  sc_i_curr_cnt;
  logic         [31:0]  sc_o_curr_cnt;
  logic         [31:0]  sc_sys_st;
  logic         [31:0]  quan_b_i_cnt;
  logic         [31:0]  quan_b_o_cnt;
  logic         [31:0]  quan_b_sys_st;
  logic         [31:0]  pool_b_i_cnt;
  logic         [31:0]  pool_b_o_cnt;
  logic         [31:0]  pool_b_sys_st;
  logic         [15:0]  reg_channel_wrb_ext;
  logic         [15:0]  reg_filter_wrb_ext;
  logic         [15:0]  reg_db_width_out_ext;
  logic         [15:0]  reg_db_height_out_ext;
  logic         [15:0]  reg_db_channel_num_ext;
  logic         [15:0]  reg_db_filter_num_ext;
  logic         [15:0]  reg_group_channel_ext;
  logic         [3:0]   db_pad_wrb_left;
  logic         [3:0]   db_pad_wrb_right;
  logic         [3:0]   db_pad_wrb_up;
  logic         [3:0]   db_pad_wrb_down         ;
  logic         [0:0]   db_wr_ram_sel;
  logic         [1:0]   db_wr_start_wrb_ext;
  logic         [15:0]  db_addr_initial_wrb_ext;
  logic         [0:0]   db_wr_finish_wrb_ext;
  logic         [7:0]   reg_data_zp_ext;
  logic                 reg_para_vld;
  logic         [31:0]  sif_0_debug;
  logic         [31:0]  sif_1_debug;
  logic         [31:0]  csr_r_baddr;
  logic         [31:0]  csr_r_len;
  logic         [31:0]  csr_r_loop ;
  logic         [31:0]  csr_r_stride;
  logic         [3:0]   csr_r_chnl;
  logic         [0:0]   csr_r_run;
  logic         [0:0]   csr_r_irq_clr;
  logic         [0:0]   csr_r_ready;
  logic         [0:0]   csr_r_done;
  logic         [2:0]   csr_r_error;
  logic                 csr_req_strb;
  logic         [9:0]   csr_r_auto_ptr;
  logic         [0:0]   csr_r_auto_req;
  logic         [0:0]   csr_r_auto_ack;
  logic         [31:0]  csr_w_baddr;
  logic         [31:0]  csr_w_len;
  logic         [31:0]  csr_w_loop ;
  logic         [31:0]  csr_w_stride;
  logic         [3:0]   csr_w_chnl;
  logic         [0:0]   csr_w_run;
  logic         [0:0]   csr_w_irq_clr;
  logic         [0:0]   csr_w_ready;
  logic         [0:0]   csr_w_done;
  logic         [2:0]   csr_w_error;
  logic         [9:0]   csr_w_auto_ptr;
  logic         [0:0]   csr_w_auto_req;
  logic         [0:0]   csr_w_auto_ack;
 
endinterface
`endif // DUT_IF_SV
