
`ifndef GUARD_SVT_AHB_MASTER_CALLBACK_UVM_SV
`define GUARD_SVT_AHB_MASTER_CALLBACK_UVM_SV

/**
  *  Master callback class contains the callback methods called by the master component.
  */
`ifdef SVT_VMM_TECHNOLOGY
class svt_ahb_master_callback extends svt_xactor_callbacks;
`else
class svt_ahb_master_callback extends svt_callback;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_ahb_master_callback");
`endif

  //----------------------------------------------------------------------------
//vcs_vip_protect
  `protected
e8C=8cV[=[R\JJAILbgWeRTPf-,Q5e5ae1d]H/C^GX_:?2FfER2(((TA>\N@NJ8-
1BHH[5G&7ggUR:Kea(84C[S?FK4WVAC]TJVFAKX3KaXZL)OI-6\0^cfRM;/Y?6.b
;@C5FPbZ8/+W:3IQ/K=gL1[a9/dY,W-gGJ+_C[?[d;a9)MN#Q=5G8,Of]&gRNS]<
,S8CbNCRPe;FKg:MD8e4?5A:D6RE-@9J+,/X(]g-YGBg/TC3&K0FX4Y>QN870O8_
F23W[+B@^,B9CX#P1LV<BQB46U1\BJ3#XO\fY1HdgZ;RTUa_cD8<75YH/O#>TY;K
O_8d]R:]JQ=a78<aP\bQKM7)(;9eF@P-@U30;QS<;YL1=8?A-=Me@M#C821J&8]=
b./2=(F.e&(AN_O9cHWKY/K0.>cGag4;^+1TI4XXS\]J=OK+[70_7A2f+#=7GT&D
E(,T&RcaST3+YY:<LAT38KIR5,K?a>a5@0LdCWKRT(GNf/d,&+Ab4=bJ8E/fB\V?
gIG8e[FJ9aAPRKQ7BG]>_<.c;ELZCf_X0TFE^XYXcHd<4eF+BN#?T8_XF^)&>JNK
a^0VHC1[=:]+\dQN[^GX.N6c/ec5d3J(_e;G246SQXe4LF/_PFU^14eH:LAC-0WS
BV/)K<RJdBC)d+.\2LObc1B<&>PgXL6?&DX:^8-+\MQ5KVV]K@.XY).1QFGPG6^>
bN-4K)6M^<S8U2acZBH7Q]aP</cGZCUc=gNEE#CYD^Q/[fFQ_8L(L/A0AV,E/XP)
8#NZHIMBVF28(Z+_+U+[f-&C+J][W.+gP?@Pf@KPA:UCMf->D0\gHC-DX_bEeV[?
_dQ0O@].+E\.IU8JeL,ELQ20MJ-,0ENFWRYVbb+&c]OKf>\+X)0&#/RVa57e-PR+
a;f.3G>;[3<dMDf/B.I/Mg5O#PP\REBE&I(I5B6Y>cWA3L^4C5E/7L9<C4C(P32]
TAg&:PX/:UA4P=5#a[N+1S;:eW))CG?R)NaL\U=[.]Ff&RQU&<I)6DZaJRQEI19W
aCYXA0aYQ-4@P)Z;C&;L,LU8b0R>_DJTPdE^eZW)UOC-d?/e<8(HB?5ID>Z\_^X<
e:UU5>0\C6AJ+]Z]:I5/&43:D)bf:.)G[#AabD+fIf9?WC>F-,9FMfggNXbJ#(ad
];XF8df:?@NF)Z2#PKERTeVD5fS?OIb^EdcbbdDf6Db7.[TDg4A5e:g5]D43KI,4
TE=GL52g-Ob&?4G3JGX]@aFBH]\?TQ22eUQgHUX.>;N/K:,FZSCX0-X9MHM;(3bB
-HWg#XY_BY-^eg@WLJ,[f1;bK5b2365B@1KX/1_cOMMD1>P8PeIgQd6IaJ75[:=H
G;+=F]8ff@:,Dd-X<T=,aTL]c:+U&&8PC,VSR4Q:WJXQIS=^ZgV#2-GgN4>c=,1g
=?:4?6P2L6C=1)K<a3V.F,FDI5LBWB>RSNSNb58O8]:?^2,)\D(;b0O_@B@UGS[>
+M6]0;Q](9VI:G/[ZZ(V]RaB#;S2BNL6AMJaEPd&f3a69Z/U0NR,?^E)70?:;.g>
:T[cOE>>Zdb=5DF;L+L#I5,S-53G<Gd@MbbYfg[3dD]A6A-gPfR^&ZS+4Z7V./T2
]<,<DKJ+:F+^[[K<bU)I+]BKWPXZ>HSg56,^<E/:T]27e/dgGE):0d025T3+_)I.
?Sfe.8V9B]_>2I9&=;IU4?QRIJC-.2Ba4<aCX,YC-HM^DIaH9^Mb5eXe[UA_.,70
5NZ)&N>4\2CT,=_8c_LYX-RQF@ddgJ\[_#eg]c&93_Z42E3&D?EKCQCMEeZ6,<Z3
^F#A)d&&Xc=Xb[SOLLRS3[69.b_M_OfCKV@5^8A5Z?GX_7Y][+XBJU_)1<g595Id
+9@dWM+LeF1fKOcQA:]C(,ZZC&)(4C=XNaBU@G.X;#ULeYK0VX@R>:<?R;U0NSE.
(Kg08[.0SPaR[BJ6T_U0E3d[WF+c:QO1gM-T;><>V=,H<BL7.QaJ0QENS:S8(/9.
2[EGGXUT_-6&MH<,80&AI@A,Jb,RC^aT;.M9]ID,BPKI;E]:T488MDPXAb:)<e^a
_W&f?.1QA,4^ZL[>Z]PQFPT-&R-L+>:.?Zc8&W\Zf>H7C+^E8ZJ\Q?4@V22e5.b?
K)]MIHSRFbFR?51&6+2K40)MLH.0ZHH;O#eg775.gdf;UHT+P=SQ4MG8ZN#QCWB\
\G2P/c/51^+XB:4<AXQ\f\97f6eU88IeW3UggD/8M\I3&GU)O[Ff7gG_X;9_aPF0
:4TTQ2-X[c50AWNV+P8;,HBWOY/6a]K,2;KXTB]0@MF4,(^]8)C\N5V.DAH8LKFg
6R1.fD2L/GC&<H2SbU)e\LBW4$
`endprotected

endclass

`protected
\G9>#@1b23);RHIVX>:81@3H?NQQbNd=YfYbU?:1MC9N,PY329b[-)AQ1cWbf2.,
_RV1^gb3X.VaH;<45=(WZY,[bT?=1d)6QT1Z;gDTQE,^W0dFC14:c\c23#6&,?YD
Td^gf_NID-e?=9_5e7&dV..cC1:/S6N&)1=NA35?c()/&ZLRTU4;[^48V\b1GAA9
).C5P2Z>-\O<D:.6?(R-Z8C78]CP7VdOCeBX]b6YFQgcb94)&Q1EYRCdNbPB#Y5N
PSRb)BW1VI9e7+gVLI.BfRJ<:E.c25R-T@BC<OM>LS<U5eK]?8PW2#CT07ZCN_IO
#EU6U-b#<S([DZ8,QN,+.2T+I0f.aN,R@$
`endprotected


`endif // GUARD_SVT_AHB_MASTER_CALLBACK_UVM_SV
