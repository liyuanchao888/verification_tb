`ifndef TB_DEFINE__SVH
`define TB_DEFINE__SVH

    import uvm_pkg :: *;
    `include "uvm_macros.svh"
    `define DMA_WIDTH 64


`endif 
