
`ifndef GUARD_SVT_AXI_SYSTEM_COMMON_SV
`define GUARD_SVT_AXI_SYSTEM_COMMON_SV


`include "svt_axi_defines.svi"

`ifndef SVT_AMBA_MAX_ADDR_WIDTH
  `define SVT_AMBA_MAX_ADDR_WIDTH `SVT_AXI_MAX_ADDR_WIDTH
 `endif

//`define _SVT_AXI_TEMP_DEBUG_MSASSOC
//`define _SVT_AXI_TEMP_DEBUG_MSASSOC_L1
//vcs_lic_vip_protect
  `protected
5WSXT^SB.8<W?=dS_.3[>(aSN0N@K)Q2YT&H?QNQ:6E5B8;P,G782(49GO9DaA9=
9IS=bXeLJb.KNL;Q@:VK#]=[ZC)4REJ=@ebEa./AcZg.^4]GDNR0(N^(S<^-U/C;
5&c]T9KX>X#@:?Y_@)DZDc4U-N:#^PV=DN(Uf4BaGfAF+IGd7P@ZcC2)7PJ&C-XW
_g&4#AEZ]bWXAcBX)5DdMT+JZ1^/_WHYAO,Cba&6/DH(YCQ+I3b)L3(6>bcH:P(4
f[.3X])a4\+bP:2[bR>d#gQG/I_^QDVb:5JLgT:\VadDR4#9^=HP@J,_X/9-<E2P
.U+=bC-&-a9Yf6ECY#Ea<W+Ld1=#8>a<IXA-f-[UfMTSG9<3fR?-W/S5E8.QS.a>
2IV)1Nc8=Ub1;?YCc9a#I>SeFV;J27:-=P9>6Oag,1_:(MXGODc7HBP,P1&>Ze0B
6GYJ(dD?S.-PV5)0F36,aR3^cK,_fP/ecf:1\+:MB?b&HP-.Q[HM9/aITFR,_52F
J<U=(TVc#:Q0URE@GANS)T.d@[\a8]eEUL3\A3,JfW4)TZBc;@WPbaDeE2(#6D<W
UX^,Tb1eOQWcZ4\L<+O+:0a=CT3T1>aQCVQECf7fb&KNTCBF7;72Z\4E;SBGg]4?
aW>LSA3e#=1=^,\;e)C\cSU-g:B3.:[0?@@H(T)a[[L&IWe@AF1PMg88NE=V_A5;
=<d/H>LW7A^RJPILI(+I4\+;/U()1H=dSPBS6<f.Vd\:SZ#:5gG[+/=Fd?7Z70[N
+K[V@90&.L5?eH&B/dU2]6VU3&?02]<B\;.9J<XM;Q9F1[/dJ@E+],(-0\[RP>=P
9[a9A?eZ.6L1MX\S94fa<gUY;V5U^9U0ESdc)?F0GHZ0\_Q?Q?KRaOc^f7f@[>4[
?YW6c7cIE?7;0Y)+?BFB[U^:[TXYK?EAY=[aE>[CNdEJPU:DN;K-<^9R^8P^P.YO
bIM)IZA04[F.4&S.aH+b_A#bZE1]UU<.+43X0Rdd\K_BHKaHN.(?DG]=Y>^0155F
?aM--N-G]WDTVdH8&(T0@:54;\I2#a95=)^c&ff04;cUH8Q6VKbg3TBJF73GcFcN
fVC1W=;L]d,](>H(/].PI);Z2HF5HOM--\[5.M_=2K7=S8g[2XN;OIBd,gFTAM^U
-;cJ&I7)Z31FQ8C?FSga#&LQd51>O5HX3UQ)N3@\GJ^eS@]<OPJ@g[5d(.egQ-G5
3QJ9IPB(9ZN.D75AM#>4-9^GC:BKJDZ/:XY0eX3@NYb)MgV05a808c[&6A#E0=@P
XbM(3Z,.,X?1bU,^(.O>Q+79g^R?]SO1Rg#V9W[-RI0E):^&?76W+(c..I-KbT.7
(._c3#6EX-G2;(7(gJ.3[-1F[86c,N(RF+Z=[S=POBP7@LaTc8_4N:U3\Gb+a:1>
bQPGH7]YRN@8L/>3_W?5H,+CTK_e0PI)^1gYS0fKAgBN2M&9FCCR\&&Ue;<6gZ97
[:B0_a8J9(e0U[HZQKZ.ZR^&EagE@/^>N/4M9+8_6-BZ9S8#/22I]+dB<4VO8?Kc
5fA95V)>7TT0K1(USE:f:??G,U,&8aVTW+9:\ffN5V?+ERcgfJaI_OA2-LY9[O16
gG-I;8A=FFE)bV/33:]>RFB#-?Md;dOB7bWE6G=(L-QaWf,0XXHC]&?ZA75ZgGQF
C^Y3Q<_EXTQKZS@T]ZeMQ4:)J+;OgS/#aSR86Y@U1J&5TPaM^BCH/99E9KVL[1L7
#8I;]X3GA6;>7]Z.1F4dUOB,VRU0FCAF[E?PHTV_X=[306;590S7KfQOcE)(8K3@
?@JHeX^KB+LC1WM,H;E1F[MF6_dPD7OHcVc1A3\99c3bQCX[aI[M_f7_D4X-D(aM
AKR<&MSP.eYf(04.</c&NDa+;P0)G:d&-9[,5:Tc[W^7#VOS_SfZ]+^?ZGcIa,I@
dB=R(98SA_4[3\Q[OaHJ9,6;P0=\Z..;PQb5T:V[+^d.).Ye=LVA[0_9gP>9WJgQ
H.NE\9=:;B4R=dIJR[E7[S:.5>H[BT_3AG.b]+B])XTHB_K#D54;WYT2M9Tc_]dd
VYJeJ9TR1>g3G[_G1M(N=B[;>HX\HIR1P;Y:/[)U,0W_X,,:5=1c_ggfg5YM55e5
4K6W9,FFIB\,^5SHIZ(^Z:++a][_\8IZ-g,ETU73N^<9Yc.9Z])2BI[TA>RPAf;Z
-,N[:(-C,b7(f(2PJ^;+1DP+8\?ZCL2\<CX:(a?6EQ)aAb_F]IXADGU7dXeWK>&V
#B/_dU:SJO>]Q=3e>#]e1L9H)<6&A8@b>b(H3S3=WD0^P\C1\[d(57EY<L&A,F9b
MR@K(\G:PME2_N?H(g]/b-)<-PXVYM[07&1D@1/=D</4/MW?YRDZI7g)2<fd\.\O
,H9(47C+?HS5FeY<K]HRPgFM&\b6?WgcgU-DL2CJ:-.M<6f0_>:+W8KKUK@N,cDA
>UW:fG?BO#DSG&-@OBf?/-Z/Y8BOPNA\5:914BIUZM:8AY.K8H3@aVWZ+He^9UAF
c[RYYV=.AN.0d=W3BILIQ&Eg:8,OIM#X4bRg4VJd+23,Zff[7?TO&/Me<AO28+9R
KgK6;OBCB^#2__P[)bI+WcLcX9ObHP@dfeQ,Gg_-QF@3@CL3(\S&+:fcH8JMJE<Q
WA8G\=T@5&1;5aSaAb?^;7+HLX5/CY;9;(B5b^f(;__>M:,,-PK;:=?dbWBaRDS(
_9b1):QQ0]&aI[<)O8F2E>83a9>:-5?L\033NCU;&/dF&a3RK2,#DP:VU)V27FJ<
AdIXbCY]F6PN0,N^;1YH](BLV&&QDL7.P^4,Z&,VE>f-.H1?@Q1&O3:d-(:LeId9
;CbWaX3S,SE@E]Ob@Q;X=bZ>:(HD0UB8(8+(fN)d&YAb]YBEg)=&_VNCSP?O0(9(
cJ^H/]2CKN0_CP5MJ#1_HRd8/X5MKHIbYVMQ970C7\-4@>TP-+]a:G&<]P>@BG]R
R]AfL#N9f?+<2L?V2[\+g0<[,8V9P:?.06I5DFYB@(KKd^Ke5@7M1T,=#\Sb?>-D
_R@f1#^S?.e852TCa@D])1>NRQ^TL\O=_)dA0ML5/0Q&gc4N(=>d6PbGg>QUHOQD
\/M&GQDG5[Z^ZEP-S.N0+&<febcG0,)g/)f:Gf:X@&L?Q^2GgOH.+8/A?CM&fVNJ
OHW)cQ.MTTWM+WEIS=GF[eGg6V\WBb1TSQLG5Cf^Da>2L1?G\M]7=(bJ,BgbIbEU
Df0>OM]gcBUL@SfPd7cfb#K)UQZ\Ne++U?-O3WMH##bX7F^3U4HA5a9UQ.4#eRLa
8&N/N9@Z\VVJ(NdKY1M.5ZL8A)@L)Z]=;4JbO^Df3Q:3Q;_<Ce9fK@:TeQ14:[EZ
bd7&OX<2ZW^L6[_S<3YGE>CN7eFcSO=.D[9Q&B>(A2&Y9]FBZ5e3FW#RU;J/XL-P
B7)4\S+Z?&BQ1d[c82f;4aS[7c\]CR\<f(Y75f.S8e:^dXe7\/4,<8:V70(TOZRX
^9.;^]A2/e(6dg@KYLB9[I.bfg:g3Z#=I[7K<PCGeSI=RR613/-bg\ZZNRFL[;e+
.JRJ+BAJg[,/(FOa59]\97[YcX3CIUfQdGS0(PHJcKTEVP>2?=U-Y-N-+VLV5De-
Xf0=JJbBYd1CbZ_TNI6gI.91-?OWIM,M=g&6X/:=0:+=YU(^(DONP0#8fTP@KZ0;
dZ3A=;7g=5NDU2=I^8dX_I+,8QdH8H16f^.=MW+0>?e_N^T7d1>V.GL+Bg0]--gE
H;QJ/^&./V/dG(#<@#a4V3CfcQC:D.B7\#5B#3dB.N=#^M=,N-P?O8M)AKA9J]eX
aL8X/0^0?JLA#?(TNIB)0/6>5=-UKGMAb>^dX=UPNeZNC0+@>Y77d,1IGAZ?<WVZ
(9NGJZ4O(HB,SS^(BV,YDYFJWJ--eP54]Pf@\7&2UU&6PM,3O5JYLE<N[MFR)A8Y
&PgZ#A(+WfD49McZWS#gV<4C+;S<-\g,1?VLIa<;#9\@?VTE./_B,;ZZa/H_YA(#
ggJ3\E]5-2(2_f)QF4[X6WQcFOOCc_K@f-?AX0X.?gGQ54.FS_@&RffQLWcKLZZB
=c\_+6HW-=VU(Ia:@U5KLX71>\Y8^Xaf.Ue9[2JbcZG^;ED&IRTacTc0VXN&OYfS
8/g?@X[1IdW^((;#^;Z.8O[(\_MH\#0d&KVZ?d1T;DMX6L\1<Y(OLg7ADeJBb->V
Y>d<H9U@U3YcK8^0eT0LCWN=e9c83eKVdbV9IaZ7\fgO4V\S@)TadI_aFNS<(6(,
9[M)J:(TPO.3e.-;E,^=)c[)1gfW;6^WUA+E(Cg/b>Og+VK8B.aUNG0;@4OJDRaZ
f-(#HKMJ^;LXHP/+P^N[K>,>545e?SV</W8[>Eef@TG=2:Q7c;A6GOV;B2b]dJ98
8_9P4V#?)T8H>-[Gg4f@1=<Qb\9fG)0aU6J@_1I\8.H>0(/X7Xd8,T+)CK@FR[Hg
#\e>_TFeaYBI5=+)]^d\JCK2M6IE69EaQb^&W3YL6D+O:</I/-<<#V36/^ad[B])
6,I:=KNPdVCQVZXW;Y_0PC6Fd-N/A[,\]a@:-OE:LX.eg=3+IQDaMa-9BG1=<Wc)
Y/f/Ug\JcA;-_f.-J_,KRR0>L5:N6W^LEG]K/7B3,7K4961J<0KN&#Jd?Y]+QA8-
G#0H5TZHUF+V\\:YW8Ge<,10Qe_QaJ8>EF=F@;FQb,ATdV(JB9JLQJ2J-YCI=7aN
TM^XV[)cH)R1(<^4U/X:R0\:A.@?Z>NMX1B;_2?PQGU]C+dIHUBgV#))NNU,b@<J
LJ]IQL_-+0WRXW?[)#Mb6B^.d5<Z9EHV@<MNd=UOA-Dd+=/WOdTO5#_@H9,)Y8C>
FT0#C60a)@B_)J3a-DaB&6FLfeR9+;+]YE+:/W4S1T2\ZK3gY39cCF#E9/0e^FMM
X)(LK8YFD-P3XZ811^]9O&ge.3aYb+N\,Y9U[_51E?^Q_EF4aFS5P8BOZdbe@4KP
R_S]MHKO&[C0(E[A-Y27KE]9^>3>GE]PUCUBZ6(WJF&UA\];e_-V+2CFGBfcG,_.
S,TX#YSF:@F[_P\M/3<#E(C,L>/1aRcG5]TL)WM4A(N-\_>HEVNH(6MIR00H65;&
)0BOefAZUU1c5eWL(L2^[#JX,.OQAUD?7JB8CP)4W1Y\0PCHP\7;3W6ERLFMPQf)
<GcK4_X\DR>F?6OfB/JDdK<>aC->cA.&9+>+9(J+.M,_NH8LB0.5\e.5&1>53OXG
N>,@)C&U^]/YM/QV]>A49=#DH=G[7:2+W\EaL4ATW.LP[:LA)ggZ^LfaMIO3(TcL
UCMaD:GM\Z@bFBcL#DV1&EFT4Z1D\8ObREa,+ZaBDacJd@XCK/ZfVNcH>>43<DDA
HF.I<E>BOZ)b@?,Z(DN5N6I9W5e(N^QQc?^e&;4U0<.)6F=:6[VdC&GG1X]\HO/#
gR\<HJ[3NeT;0Ld+8MB]0e>f4327_9c)A.>CBNUL_=J]ZLACZ26[\MeKD9&Y(+1P
<0=4K4JC9MGb;K\Z[af6G=[]-_C)U^Q:4MXeWg2>B>#bAfXDZG@)ZeHHY)e8@MM9
e71[_2,UBY?VaIa^:/>@a>704+eII:#gS&0\WKOVZ-e2VU)U)T_JH3,4XMZ1VF1)
IA4X3=T;21[UP\3O5?C--d=J:I(K?V#aN7D:./XXX708#;f.._D.@4CEH@K[,16+
/dHB/^4;G?VW3?KH>If6:[VDB?,?EY/Bd^:8d/MDc&R6Nf;#PL3W=A_^D6QNY,,F
].JMM3cPBTdA6^ZU[D6<(=#4P[,c7EM@FSL\62HKY.CDN/:^XM22#b>?e,d3X4\&
5X8,Tf899W4<-,C[bF\57]JWcO)ZLKZf2I[^g5?8()W_O8T18?EH6S5<Z41(0#Vd
:d,N?F<7b+fY8-B\eUFHa5A[^5Df@IgDNa-EK:[Y0B[VQ&O=MA_>VY[ARQJ(SO/_
>FF:[(A:F[4\2_=>YMcXN_]\3L_5H@R&J+/DQ,\2&__W?L)f9GJ9455>Q_gcV0)O
A-I0Ie(-6&a.A4WVLU5\a]W&N8a,;g+]5gT(706X?,25EIBG-6ATZY\=-15f]\_b
3>MHM(\@RG.4U78M=^d2,\G[Ya@U(7(_UN9,44J+OBILSU+b?d_=M&g(a^4ge)1#
B\SUb-K.KQ6\NI&#-6<C)9P+C\OB+X[8JTVJ&NLU3<JS/GbA0@U9O07+dKIe>&]C
E3\\2e0?+:aPTO@[UA[:eLEM7M^bb@?4Y<X]IL?DXBg6:A0O.)OJ1D;-L_,NE8JE
ISSGL/cH-#;6eQCEBNcH7aUX2(#@#3.UJfBX>0Lb9=4CWSFDYGJ</W:)W6ZI1<[Z
D4@\B,/&M?A@L/:0ELT?[R6J6Dd^-#\N0MMQ/5OLUW3#ZadT:(I.13=F@.U\fa]P
-481[fCVR?(C7[;7S?A98HTD1;?CbP)UGY9LG#7W\OZ8QYe.GRO=4D?_]ZA.6K@&
9)AT&@S3I^)O6bRVaBX-YN7(#W>6g@6P+SX.Ab>(^F?^gc-[E#S7g=9]@e&3D>Wd
6(X>#cS^aCZM;LS8+dF>MH27Ud]e@g(^K1-G)N4.22GWV8IGM?<UAP6FI_cL6JW;
:P-dAgCU:,c?3K^;OMF2]5&:#f^CAaNBRgS6C?D8bWMWLB3YW_5A?R+&a1?dLRO4
/H]>,MM&g-EMP^GgB5dXbYIAL,A9ZQNXC7R;aJ2eZ68P\A4,NK2fK3:@O<[MFBKL
3D0<Z_6@b6[V_.FbWIICAY:E/O8,>WTa5VRcN5)e&DC0[(c#a_^Y;JR8^TK=>)T6
P\&9b>FRff&UKZK3BX&ZdU_S(a00\65;_9DRUFX+EDNBb1>82?^bW]9LK[S77(H=
Zb9,&#<G@f<_M)c=KZa4++M_:a]4NXE)[d^aB_Y.XU_T2WgZBT1dDXbI?EE1Pc>?
eVSI@G])ZUC<QccXP@R?bHRX(@^=D>;+@:O1<>]_SC.K3I^Y4:)PE\6M+3ObXfO@
5N1,816(>GRU45V8g8SF,PJTc)a]>Q?DY7@+d2<8E;QY&+4[I#)&eC1I]AfG)KJ.
2Ja(^?W.N=BP/CMBE>=N-..CN4c,L:CT2)Q\M]1Z-Eb.@E/aG4;3--XL=ca3N]\B
b<?\E4G--VSQFNG_cDJD.9X,WX),O#:S+_9e+T1\Q;/Q+^38DXS:KK8.,4XX8BQd
H;ZLF[(&DcV<;L+8dGHH>0?J[Dd.UA@OC4,W?[R,XGDUM;O[cSGXRe6&=<IBfB(5
^EbeUF/3BS?T]RV8K3Nd)-@P_MSHCFCN=(;&RIe-3Edcf9/fPe0C.1).;/aLf<UT
0XUS_\-8IA?85JAD/-AQCRGHQb>#&Fa\^)PE]LT>8L(H&a23S.+MIFQ\UcOH5J7P
=X)4,@RfTTI>=B?TBUI@@cC8b7CB[AK+EC+I3-6?B-4CIA7USMY]1MLD;PRSIcNX
4.PEN>9UeFK6[Oc6AV-eB<UEU(,Z8cd+D3+A#R.gXY;OO+.A53L0TY^AdVa/5c(W
MHN-[NFcQK(NRLDHGMdT)>>IPLB>3SVCJSJHEHD=LcPZBMe5##ATac35>&UV.MaK
gGgY<M8OHRZU\8b:N0RTO^I5FN/1P9Rd9.)a\MM[&/[M&/GMD\=AV&X(V7S-_M>X
.MAFeM>a<Z\XQ#5d@^f)eTQ&NU_BHV?adKO.Z<I0(<LO0&53;R]Ef:3A\GL6P;;-
HTF8-?=+;D5=QFK-Kg7XKeANf)GRe6TP-(<=/7EF:H-(c@\S/6^,A\W]Y@@Ab3WR
/gVD^U/W46THUV&I\PQfQ[a6R&U8/NaE\LJ<f2f)4IXJ5-67YH;A(T3LM/?cW=3(
TUf/]NAVN5KceE-SV;;BW79WXI2H&/bB+->7?QEg[P#c29/+UfW3\BCaHWJHF(0>
\9gN>AJa#/\da+.JEEG=AOXRPSI)>J2dDJ9>.5K[WA#e0<f]Z#T[DT1?(W:gO:/U
+,ed#5+\#59VJaE)6+Wc<E+;M#cQeNU>eE18e>0:22;eX)DNKNQO+OQS\^PEg]AC
C@^WJdfM;?[30a5#eYI4,Dc8b_gCDgENf^A2V1gUXDF04)/GaV[_A0#+6Gc(92//
9aYO=T/G16_5U=Q:NUd,g7eB(?VIWcTUN;e>cY?S,Za)K?L@BGWX2Q2daUe[@c+Z
41J4=@U/fT^H:=0?SL=(YgD[=T^SF+V0a4PJa,<M][Z/>9EYNBF_K83Kf1S@G;fa
=#PD(YLOSZe(7B_K7YOWeMZ7R00YeQEfEV0I/G51=>AACfR[=Bg9=FS+;_#N1DJI
Hg\6g[<:UP1IZVf2BX5?YN3Ka64IIQ85;(H8^[EWadK?MA<D<aR5Ta1de_HI5X<(
\1ONV<S0?L]Z1#)&6D,YN9C.L;(++Y,JUAL)d0<+R&WQ]bE=MMGJ^/U[PIJ2C\Va
DQ>TZJ?L:4=-I=4dSV2=E.,fWa8Q+b:X9P_A@XT__RX))eMXXEfOBDD]FYGg,=QA
A1AB=-B(OP7UACZeR;8XeTdXbLCYF]H)LTD_3RfQHOf\8]2>.AdLa.=,/0^g3I;<
AWY>f?YbE/Nb0MNORF4E2I]+?(#>.EaCWMDgVcANZQS/NcfY0T[I7_#L2IFA@OPg
2Q:D7[3GD5H8V=EC)O=^]N1<7.8TZ+Yf9],L)KAHVRYg-T-&dfS7Y+;+_UJRMaFb
.aK<0JFg@/dALc8&?N#DZ,C,B<RME?cX)\CY-13+M,.f<CM=IRC@90/)b6[2I<SJ
:<(RO3A5:?VD,_ae4Y0TUM&>LG.(YH9D^7:K+Q-UX7Bc?&K5eKQP6P:a9Q.UbNBS
]3);X332\U3<ZPaYZL[^5Oec3YKXR)@Z44M5b6=.Q2-+_;(N,9TL4>T>9>TNIg&+
(9/@9LGZd37&<@9WGY>,GBYGa=[6LKC4RF>4[M(9K==bfOKUcLXLY-I+IUL5T.>0
ROKaZ@S?e:[^e:9BC69>0E]J2XH<.(R.T&JWa3;B\>U6#=9U1H(Q0bKR-)[6\PeD
.R&V1D(FDK3[UV&@4f<;fOCWF#Wc&O3;H155Z9Kf/-VM@5A?3LVRYJf\KIUKJCML
:IgcMH=59WKR,\X4_6(Cfa\_be,;D5HC?\4J9eLYB;-2LRS+-TaZdfGc))\aY+eP
4#WZc95eC@=]]([-a7?(1UO9\8G]_H?I0aOAaKTA29^AFW\@,CYZO)0DdQ]UBXFc
XY)H#=D:Pf^6I\AS-Y8?<U:4bBG8Y6b.NN,,^GUHcB89\&J+TGScDY.ZbT<K&cM+
Ib)fDSD9;bKG-\b:5Q]MSbA8(a?V5QHa2XJIdKVWDPWCdUC&IBSI=;Z2D<fbg#7L
UF=6=04QC+R.eOS=d+?bGB@Z>M])Y9L_95G;@+d6ccSTYEaZ]1_aAGLV3QZM,W&#
)^d)S7_^?03>^TcWO:?ba4[CP^Y:C,JFA>WQdO6RbQLK8-R+0bH344ALe<&519?e
LUb+A&/aa05T3\CG?MLgFQgV/aRcRS[/_]^A&+SGW8F<###b9X,LR&A=#D\N34g+
.QR,=AY9<-W+3>4?Yg41ZZ.U)96V+.7&]@PX5U+,=5JL-#PJ/bA_W20&:Zg:ZP#0
QKE8ASYA]JV-1/<],JCQL/GV6R[U[YL_R=Da[AJ^ABf<]CAK9)[b:S].MJU7L@2C
[Je+EeJ8BKX@YW9W:cYF@C-b:<dEIBTG=f^O2EWN0IeFCBW9^/\J:?LCPYL8(E2=
g+J)#_f_38F4]e]F2-QfeM(EXE8dU?FaYT]a_3=Q]GCD2^Pgd0:1]e,bS>a-\FB=
Gd98CGL947?IY5D--@dX(0gN+4+bT-F[RY/01H^3=07#94,7CaQ2+aNN(GeTG2<#
@2TBYQA4OO06PVFCgP;1_H#LLH826,aAb_T)@_:c6(JTEe\MHGe4B,1<J\]VFBg)
\WW1A85DU]GJ<caJDO.d<7-3e[=>11N;PXY&:XVCY_K,MO0O3.>@a)[RUZROGI)^
)e+>(N(R^:Q.JEKCZU43I/XQ5aS80eQ:B;Nd-@)[9T@H=643+_W,\+-NZ?V?7D<-
@4FLaQeV_[(A00-RcWfc<gFA5,MG<gaZJO<@D_,V,6fd@e^\1ZE,YB]\LWLLDM6K
gS6Z^>Z(AYIH^Q5<:)@NV0GEcDdP7WV4fV-<B<Zdgc,<Gd8DP9T_;\b\(ad[[eAE
6BJP5GNZfOINfbBU-1eP0HI<<KIa/2F;FNY/f?[/C(<.GCTc8=J9/Qd_.c\(5W37
4]QGGLg[6AEV.T=A<7+/XGA.FSP&#QA?-8DGfT.XDBNB+1:Y(3Y/E3[2YEMZ<V(6
9-.4V;EPI.#7886/#6fdb)2^J+_gd?)\UQ/=I;B0IA<Dce5IK&>T]IJ#7FRVI?-Y
B&Eg@8XY_.H1ELX:(I;@dAdD@EH@RdPcVQQ9+#Hc:V<&U/]OgL8cP7.4-5S-HE2T
->JF6772NL3:7]EK:&PaR>^).?P,YI-#)RdHT1CKc^](c/V1g26N@d)88VNWNEU_
2,N9&8(/UM-fR614L5-VWWLDZR)ZTMX(\)73RYOD-bS-;+VN)T72c5][IfG9HKfT
;+,f&H+0(a?4EZBVWPK)JO&&F;<T7U^Kf3a[K)g:VWQ2dGa7<d;V.>@(L[eb:O3f
Z<G((a#H/b6IV?E7:K(Se8<g3V33O/fGSR2^1=+@TH8IQ0\5a9<WYK485<SYXY3]
A9OgXg]d:I[(Qg;N[^C#QHVd_4e+N#70E5_\ZV23Bc#DS&SbKJ_Y-UQO<YZVA;fS
T6_A6Tg_JONXTR2+9TY8QHM+CI4UbcS3-Q.9bO5\/CB3(8ee.fG67R8PD3aJd2^K
5U,PgUGY<+PTDe)Ya.b1PSG0@PA_eA5)X^:]#0(1<F:0>?:bE0U[92&VBV<?ZJ<E
=-deM<_XMAQ7&EEB94GUN2@eFD_],OZ@8^I:eM_P.GL+T+e?QEaTUQ&W>-gT?.15
;J19(3H+8]7.+A>[C9FLEeVN>/f1LE[1)LMT>XZ?6TgV?2cSEHNMCXecZY8&&Me^
C4>SBE7^CYcRKK+SPQUU(fRW\]dd@00Y-DS\)FY-74>0BU3Kb.VQM5],)AOS-V\[
aaD7&>@Y2A<3.=8<:R6U&2_G-(/R-LEgd?Kd,::NXT[LEZ^\@74V:8X4IWV)>DJO
GfWfT)+[(DVc?NGG5C?g8(XGJ<7=AO195X(A^@U\f4^+R1c@;KM9;gQCR4e@?,\6
(OTZd0e\CF,_/\5-V_9b6YSH]&=BT5@R<80H?bO&WP^4:9V?]SYQ9UVQ#],P9E[\
(1MG4C>:,f,0ZS0?-^\HU-.F;6&>6HBW>MT38EMTA^\C2;IbKTMF@2JdS&.d?]_^
2Z_/)>HP^;BcdR^O9&BGfb_b(<^->G+;cX<7.(9JA#gB)NUJCS(daF-RIZ46@9fO
RYg/M/f40g7Y-[==(2KZPF/]XI>U:YY#QQWBRF.)UZ>,SJ<TWM(f[4]H1SGYWK)b
R#Ufa(Cg(R604:=6LFR1ZI-e9C8&g,Q7EO4MK-^#X9#\4PZJL_Ld9-X/NL<ID.D,
M?PG2fW8^OQe4NfOG0U(#@V?gS;fR6Cf\<S](2adVV;N)X&S4]0/<@daKI83V+LC
XXgHfOcdJ8\(J&7/NQbY;.@#^[YfeSBd+2cQ@DK0JF1K?Mfa8V?ZFceSRg^64\DK
741d;e:9-eYV+()V57ec1dWI,MI_OfO0&?/:W6.7-5Ia=@+Z<bE&Ba]5T:4_K/1M
F/\W0fZc(/^Q^K^,A83L^.^(>ICBP7-S7&/a0<?/LH\g15XK8U4;.5PQSBM]:cHc
\?B3Lgfg7Je5&5S5\b.EcFEL,#I4a/W2O:Xg\YA/62VX>LE9>ZBE8RG;4.28YS58
J&B)70_>A^>F3W0QcCNOAGMNWM1KYA7=>3<YI]HWC_#)8##/Q;)Me/T9OB#/Sc&_
FI2dP9AQ@IB@g<W(2^<DYOW8A]0[U16?Ae#a@+2gc#<c6;bQ@F1Wa;b(8DEfSL,g
>RNH0I=H-.#Z;2?:.YMd5,#&Z&U4LfD>B?RKH+ZIGCND18K5^IOZ;JF-.3D]ZIWX
8\2S9C9<;3JOY)&J/,V#+1QE7E)A8_D9</F@a=b<0T6>TAHG1F4:YMHFeJbK=T7d
3_A#1L+T4f8-bA4&.1V2V^>CHKPR4e=8,L\&RJa</LPZb6>U8B8M>:-+.E/DdM@>
b2H#FY@K5/+RUCc@WV\PBL3K(=a6U+CQXe&1#(?P3.7PEDIb0OU80cdX##Y#RSHQ
L6:(3FKdU4>DB&=1+_Ud>-4cBIb#?ce(G8K6#45c22dHVgPG[@=McgDB](F@&ZLB
T5.?DSgR;6T/-=H_Q_/LW=ZOGH8RVU5GI]@Z=L=#3\<,KI_3J)e\H09\9/H=]Va9
e_/,]>=\FOAb]ALY#8TWO]S<;H22N[Sa6aT#BZ^5/g^HBX3J5-8dA2/3HW2C9fN8
]=dS\&SD^63c(Q>Y00(.4>M+8^OF548XRTZGb&\-60]K=SZ?bEQ5C1Q;-@B>Y/1)
fZG8+3eX?._)6A&&)1cS3.COSMHJF(72E[?AWOD,cTI;Q_N3/Q6XKScWe^#X_4QT
SUD]PDXW&?D?RH_7H[3S=d=6(@I8K>>L#0GFHOZXY80U4W@34_AH@gFBCgO>Q=<@
U.:a5FWB9CS&S,]bc.bW;,N^G<^4g>gLOA9^/d57H7]ETaUC6Y#GQKN2ZB=QfY]U
a,)cM@RL9F>fWJ#^Ma/(gA48dF-AC;?+R21:7?9>GeGAQ+9#LP921eE9Ob.B=19S
#=f,\Z8E5F[C2KU?(@,4VaYSNgJeK,V7c57TRGBCA2gFR@^(U@MZ+@TGFRR^P;)_
?G-X(c)25,8]cFTLN[@GX/eTYU.+AaH-SR57:H5Be@_Ce6MT8B-VaGZWJ_V&6a=^
X0AD@6d-&;YAaU_1A?cG((D&]S^QaX7E[(N\)QZ-@66/3?3GM4(fG:LQP<;B->gH
UL;8eTcc@AKKXWY1_d_Td=g;^<)AOIU6LEKH2]V\X&CG:O^_FTKY]PfY^bdP<;b2
V/>b+,8#N:Ta+9?;;Ta12,\O(EWdRbDDI5dg:7<39HDG;RdI\ZM/VNGNL)Zc-UE)
EgGV.<56Q?HK9&9JUE6G9D4;J.4B4\We\LDI<>GC?6Kd83DG@SW34W8\D;3VLH0^
MeX0<P62Oc@E,aQ?YQD6ORYe:g7/FP44W/Q0)V0I1<,)&A08C7;<.0aI[afU<]b:
D/UNE;Q2LF/GUK)9:T7A:9H(NP_5aW.LZVG,W46D:Y@G6Taa2WZ4</Q?<ZPEV8-B
]-d^W>:]<1)-(ZX/.fV]18KMEfN;M+<f#Q][ZZW\#VM+]>GeZ#4_Z#^U<@2Dg>]4
d=&[NBc#U_P1e^=J+:#U@f8>78]\1037^A8IgA-55[If/;W])Z@#OZ^acg\83D9B
N+^WFQI;6Y7@d0Za9#C:Q^U?c;^8Vf<:&.cDVP&1M3]@R8TaP)fBc#BWD:-0.5]_
<W<_-P#<<da&:]Nf@?[^5\I]1cC[:8-D\>T\[7NVTLF_ZCVT^>T\eJNT+2A8d#.,
CA^EDU(YGV\)31G+#VHO:Z>aHI#@G(9-+G3-J&X3_g=/U+UQ#bBfOZ:;a5E7EN/.
UM#5e-2=GIMf1\6Z,a</[SaUgVXdM2B<2)bJ=V)ROZS.S#-L\g2(YIe,B]S8+VLH
@JAb3C1:0g9eVB:LXU-E]aXAN:=>O&:]3[>WGU2FOSJQA5#OHC>OL_4C]U+]6C<c
-]BX+A:KCRQ@FRG/FfB&B96QQaPf5ZE<9MN:K-Xc>DJ[J8RA^cY0gI_<X,a7D.JL
dJc9/08SbMGIRb29C3K1_H1J^K?ZfM><bgY7Aa6L\;Z>EV7O[AHX1,YfDR_X>JL]
IfQW#Y)U^5bOBd#PY34C@I>;GUL&-X0GU8I2fB^0dO(H)cSe?<A8,\Zf/:7L5A;)
3.T4DO+XeUC@TWWHLMAb4J6D@HYN9B_L_#J45MC&&D4C&_4?3M?X3-8R69d169a+
@dH)5S:Q4IdU_9P-V))BEHQ8SF^^;RQE?N@CUD[SZ/D>=eI/aIBRD3^gPWF/8G9K
:Z9_H[K^^&N.gRVDSV)71fED7(-ZG\19IEMFf).>,a=X1XB4H)N&).,4cDPNIKOI
>.3T;b0_#DXOZ5Q]OEe4>C:8c=&?IX_4\)T1H^M-U0R7cdR9D/d?a0DVd-=0T&Z3
K5dU(,g;Y@JMH5Q/cCU-W;d6BKHQ-acQ<&?b0N^-Q)R.3VLOJO[<RTSNI=C&#\C,
VP+_DB>@5&Y/F5+Q.G5_;D@@I=[Lg7eSQDEC>d;#@TQ8+UFNZb#>D]A^F1df)c7R
Nge7E,<AE[5]./:EQ93a7+#b+:129GXODgNKZR6dU]]aKLYE9M[7Y@I?E:MJWAZeV$
`endprotected
      

/** @cond PRIVATE */
class svt_axi_system_common;

  /** Report/log object */
`ifdef SVT_UVM_TECHNOLOGY
  protected uvm_report_object reporter; 
`elsif SVT_OVM_TECHNOLOGY
  protected ovm_report_object reporter; 
`else
  protected vmm_log log;
`endif

  protected svt_axi_system_configuration axi_sys_common_cfg;

  protected `SVT_AXI_MASTER_TRANSACTION_TYPE active_master_xact_queue[$];

  /** Internal queue where coherent transactions to slaves are stored */
  protected svt_axi_transaction active_slave_xact_queue[$];

  /** Internal queue of slave transactions that got an error response */
  protected svt_axi_transaction slave_xact_err_queue[$];

  protected semaphore sys_xact_assoc_queue_sema;

  protected semaphore slave_xact_queue_sema;

  /** Semaphore to control access to active_xact_queue */
  protected semaphore active_xact_queue_sema;


  /** A list of system transactions used for mapping master transactions to slave transactions */
  svt_axi_system_transaction sys_xact_assoc_queue[$];

   /** Internal queue where snoop transactions are stored */
  svt_axi_snoop_transaction active_snoop_xact_queue[$];

  /** Internal queue of snoop transactions to be deleted */
  svt_axi_snoop_transaction delete_snoop_xact_queue[$];

  /** Queue of transactions that were a result of back-invalidation */
  svt_axi_snoop_transaction back_invalidation_snoop_xacts[$];

  /** Reads which have an overlapping write during its life time */
  svt_axi_transaction reads_with_overlapping_writes_at_slave[$];

  protected int log_base_2_cache_line_sizes[];

  protected int log_base_2_slave_data_widths[];

  protected int log_base_2_snoop_aligned_sizes[];

  protected bit is_amba_system_monitor;

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param axi_sys_common_cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter UVM report object used for messaging
   */
  extern function new (svt_axi_system_configuration axi_sys_common_cfg, uvm_report_object reporter);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param axi_sys_common_cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter OVM report object used for messaging
   */
  extern function new (svt_axi_system_configuration axi_sys_common_cfg, ovm_report_object reporter);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param axi_sys_common_cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param axi_group transactor instance
   */
  extern function new (svt_axi_system_configuration axi_sys_common_cfg, svt_group axi_group, svt_xactor axi_system_monitor = null);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE
    /**
    * Checks if the address of the given transaction overlaps with any previous 
    * transaction. If there is an overlap the transaction is suspended. It is resumed
    * only after all the previous transactions to overlapping address is complete
    */
  extern task check_addr_overlap(`SVT_AXI_MASTER_TRANSACTION_TYPE master_xact, string master_requester_name="");
`endif

  /**
    * Waits for all transctions in overlapping_xacts to complete. Once complete,
    * the suspended transaction is resumed
    */
  extern task track_suspended_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE suspended_xact,
                                   `SVT_AXI_MASTER_TRANSACTION_TYPE overlapping_xacts[$]);

  /** Indicates if there are any full AXI_ACE master ports */
  extern virtual function bit has_ace_ports();

  /** Gets list of system transactions where master xact is not fully mapped to a slave transaction */
  extern function void get_unmapped_system_transactions(output svt_axi_system_transaction unmapped_xacts[$]);

  /** Gets the list of aborted system transactions where master xact is not mapped to a slave transaction */
  extern function void get_unmapped_aborted_system_transactions(output svt_axi_system_transaction unmapped_xacts[$]);

  /** Checks read transaction timing relative to the last posted write transaction */
  extern virtual task check_read_timing_wrt_last_posted_write(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  extern virtual task do_master_slave_xact_association(svt_axi_transaction slave_xact); 

  /** Deletes transactions from sys_xact_assoc_queue */
  extern virtual task delete_from_sys_xact_assoc_queue(svt_axi_system_transaction sys_xact_map_queue[$]);

  /** Checks protocol restrictions for non modifiable transactions */
  extern virtual task check_non_modifiable_transaction_properties(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Checks data consistency between master transaction and slave transaction */
  extern virtual function bit check_master_slave_xact_data_consistency(svt_axi_system_transaction sys_xact, svt_axi_transaction xact, svt_axi_transaction slave_xact, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id, bit check_one_to_one_mapping, output bit is_resp_mismatch, output bit is_dirty_data_match,
                                             ref string master_data_str, ref string slave_data_str, 
                                             ref string master_wstrb_str, ref string slave_wstrb_str);

  /** Checks data consistency between dirty data of snoop and slave transaction */
  extern virtual function bit check_master_slave_xact_dirty_data_consistency(
                                  svt_axi_transaction xact,
                                  svt_axi_transaction slave_xact,
                                  svt_axi_snoop_transaction snoop_xacts[$], 
                                  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] snoop_slave_addr[$],
                                  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_effective_min_addr,
                                  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_effective_max_addr,
                                  bit[7:0] slave_xact_data[],
                                  bit slave_xact_wstrb[]
         );
 
  /** Checks if the given slave transaction could be a duplicate speculative read transaction
    * This behaviour is seen in CCI-400 where two transactions are sent for speculative reads
    * one before the snoop starts and one after the snoop ends (if the snoop does not return data)
    */
  extern function bit is_duplicate_speculative_read(svt_axi_transaction slave_xact);

  /**
    * Checks if a duplicate read is expected 
    */
  extern function bit is_duplicate_read_due_to_overlapping_write_expected(svt_axi_transaction curr_slave_xact);

  /** Gets reads with overlapping writes at slave */
  extern function bit get_reads_with_overlapping_writes_at_slave(svt_axi_transaction slave_xact, output svt_axi_transaction xact_reads_with_overlapping_writes_at_slave[$]);
  
  /** In case of WRITE transaction, gets the number of bytes written into slave memory based on WSTRB */
  extern function int get_effective_write_bytes_using_wstrb (svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact, bit slave_xact_wstrb[]);

  /** Updates the number of expected dirty data bytes for the transaction */
  extern task update_expected_num_dirty_data_bytes(svt_axi_system_transaction sys_xact);

  /** Gets the associated snoop transactions' data as a byte stream */
  extern virtual function void get_associated_snoop_data_as_byte_stream(svt_axi_transaction xact, svt_axi_system_transaction sys_xact, bit use_dirty_data_only, 
                                             output bit[7:0] snoop_data_as_byte_stream[], output bit is_snoop_has_data[]);

  /** Waits for all the conditions before a master-slave xact data integrity check can be done */
  extern virtual task wait_for_pre_master_slave_xact_data_integrity_conditions(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact, output skip_data_integrity);

  /** Waits for slave transactions with overlapping address and which have started earlier to be correlated first */
  extern virtual task wait_for_other_slave_xact_correlation(svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact);

 /** Waits for slave transactions with overlapping address and which have started just after this transaction to be correlated first */
  extern virtual task wait_for_later_slave_xact_correlation(svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact);

  /** Waits for transaction to be accepted */
  extern virtual task wait_for_transaction_accept(`SVT_TRANSACTION_TYPE xact);

  /** Waits for the address related control information of 
    * transactions in the system transaction queue
    * which were started before xact to be received
    */
  extern virtual task wait_for_master_xacts_addr(svt_axi_transaction xact);

  /** Executes the master_slave_xact_data_integrity_check */
  extern virtual task execute_master_slave_xact_data_integrity_check(svt_axi_transaction xact, bit is_pass = 1,string desc);

  /** Executes the interconnect_generated_write_xact_to_update_main_memory_check*/
  extern virtual function void execute_interconnect_generated_write_xact_to_update_main_memory_check(svt_axi_transaction xact, bit is_pass = 1,string desc);

  /** Checks if CMOs were forwarded to the correct slaves */ 
  extern virtual function void check_cmo_forwarding_to_slaves(svt_axi_system_transaction sys_xact);

  /** Executes the interconnect_generated_dirty_data_write_detected callback */
  extern virtual task interconnect_generated_dirty_data_write_detected_cb_exec(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Executes the master_xact_fully_associated_to_slave_xacts callback */
  extern virtual task master_xact_fully_associated_to_slave_xacts_cb_exec(svt_axi_system_transaction sys_xact);

  /** Gets a string with short xact display based on provided transaction 
    * An extended class can append context information (ie, the source
    *  of a particular transaction
    */
  extern virtual function string get_xact_context_str(svt_axi_transaction xact);

  /**
   * Returns the requester name for the supplied master transaction
   * 
   * Note: This method must be implemented by extended classes
   * 
   * @param xact Transaction for which to return the requester ID
   * @return The component name that generated the request
   */
  extern virtual function string get_master_xact_requester_name(svt_axi_transaction xact);

  /** Indicates if a given transaction generates a snoop or not */
  extern virtual function bit has_snoop(svt_axi_transaction xact, svt_axi_system_transaction sys_xact=null);
 
  extern function void print_debug_info(svt_axi_transaction slave_xact, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_xact_id);

  /** Gets split transactions, which are split at cacheline boundary */
  extern function void get_split_xacts(svt_axi_transaction xact, output svt_axi_transaction split_xacts[$]);

  /** Populate resp and data in split transactions after transaction completion */
  extern function bit populate_resp_in_split_xacts(svt_axi_transaction xact, svt_axi_transaction split_xacts[$]);

  /**
   * If complex address mapping is enabled, this method translates the supplied master
   * address in the transaction to a global address, and then uses that global address to
   * determine the slave address and active slave port ids.
   * 
   * If complex address mapping is not enabled then the address is converted to a slave
   * address and then the port ids are obtained using the legacy methods.
   * 
   * @param master_addr Master address to be converted (can be tagged or non-tagged)
   * @param system_id AXI System ID
   * @param is_ic_port Determines if the address originated from a port on the interconnect
   * @param xact_type Transaction type (read or write)
   * @param is_tagged_addr Determines if address tags are present within the address
   * @param is_register_addr_space Returns 1 if this address targets the register address
   *   space of a component
   * @param slave_addr Local slave address
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @return Returns 1 if a matching slave address was found, otherwise returns 0
   */
  extern virtual function bit get_slave_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] master_addr,
                                             int system_id,
                                             bit is_ic_port,
                                             bit master_port_id,
                                             svt_axi_transaction::xact_type_enum xact_type,
                                             bit is_tagged_addr,
                                             output bit is_register_addr_space,
                                             output bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr,
                                             output int slave_port_ids[$],
                                             input svt_axi_transaction xact);

  /** Gets number of snoop transactions that returned passdirty */
  extern function int get_num_snoop_with_data_xacts(svt_axi_system_transaction sys_xact, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr, bit is_pass_dirty, output svt_axi_snoop_transaction snoop_xacts[$], output bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] snoop_slave_addr[$]);

  /** Gets the number of slave transactions associated with a dirty data write by interconnect */
  extern virtual function int get_num_slave_dirty_data_xacts(svt_axi_system_transaction sys_xact, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr);

  /** Sets a variable indicating if id based correlation matched */
  extern function void set_id_based_correlation_match(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_xact_id);

  /** Sets parameters used for sorting transactions */
  extern function void set_sorting_params(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Sets parameters used for sorting transactions where both master and slave xacts have slverr response*/
  extern function void set_sorting_params_slverr(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  extern virtual function string get_ms_assoc_dbg_str(string dbg_str[string][$]);
  extern virtual function void set_ms_assoc_dbg_str(string key_str, string desc_str);

  /** Utility methods needed for correlations  */ 
  /**
   * Gets the minimum byte address which is addressed by transaction
   * 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Minimum byte address addressed by this transaction
   */
   extern virtual function bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] get_amba_min_byte_address(`SVT_TRANSACTION_TYPE xact,bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = ""); 

  /** Gets the max_byte_address for the given transaction */
   extern virtual function bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] get_amba_max_byte_address(`SVT_TRANSACTION_TYPE xact,bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");  


  /** 
   * Checks if the given address range overlaps with the address range of this transaction
   * 
   * @param min_addr The minimum address of the address range be checked 
   * @param max_addr The maximum address of the address range be checked 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Returns 1 if there is an address overlap, else returns 0.
   */
 extern virtual function bit is_amba_address_overlap(`SVT_TRANSACTION_TYPE xact,bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] min_addr, bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] max_addr, bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

endclass
/** @endcond */
`protected
7>W6YU(7_^WLe.V2IWdNa=)>DE55^[1A+-WRaH/cL]7<7Ie,,#S&6);KAg&G=M@G
7HDO30W3TQbMV>R2dWF^Sg8\AWRORc[XZSc,@X\F75K]1RYY(_dgY6UBPY2=C]^4
@Q)>g26bVZC3,a3PY)7KAG,)S,U-O&X6McANH#5BM#U<)FM([^IEA)S(cCe?H[ca
S0#Y;?Xa\:WZXd@;d(+&G;aK178e;d<Y97CAaAESd6D,8Qc=54WRB+A(RMP#T4#:
.K1YM2Qb@O&a-N.E0f8@V1,N)1GW06DMZKL\ZFVIO:0,O,77X#3H<B2HJ^P_g,T+
UPX,-NF:HJ1NR/1S&W>;YEaSEC1#PL8d2,b(8f-GQ.bP751VD7K7(60RD-MJRBNS
[<@3aP86(/1V[e:)c<?SI<6P12;TCJ]Bd-aWTUV:+1EBERTDgOG>GfSEf^B5c0J;
BYA_IHA-8RdN:cKa28+bN\Mf4II;-S)/@UfU[L7e6f1,#O&6-NJ-GP&M7N\A?8eG
c@_BJ3035NGDIK743HfJU/W,9YOU&8WKGL(c?V<HNBgCRfH&bfBc-dfF#N4#e32d
gEL6aQ573aC^d8De871GPO42T2^;95ZK:QZ19-J([BU,O]G5&-H&ZP^N7YZBL0N8
(T_CVc<dU5COedOeOZ>aK@2R<#(.X\R)dfQ4:+</bSROZE?c:C[F-R.FZ#PBT@E:
A-QDDb^d,YO.KJ_C@=.;eB8=4FGSa)Z9=)HbX@g1AY3d#DV03:LJHL@/gS1X(1I,
<gf67Q]JK-:F)[@H6ALH77IcJDWeE[\<cI]=I>\GOV)2P8GWa/c<g5KK<GY/bV/.
EgJ]XJ/H/g9N.5&SNg;Qgc<d^4&H6TPW\afAd[c\MB@=+8SdQ,FeEIZALa2LTRIU
fKdQF=C(&d.9dI9EaU.Q6.b./)+20d30AcR)fW@U#DRLAV,gQY9G=::NVV1DMFLZ
MIY1/45^&FEE-CXa>QR73&HH;7U>_1,YBJUU?a=2?+_8Pf-JWd\]N>d-YW#8E0>J
11R/0OEZa4)_5+YU[9?bb<2D<gTE?-W8C.[PH8:&I1VDcH<P5/?;30TfL=(8_gYb
G,.HW0(S.08b=[P;&c#;@&bGM:A\c-Z;=\;2)2ERB./8DSED\G/4G&P7I3)T=LLa
>fU7cT@b22\>L;20AB9c::-B+)c@CO(-55,YQR(2#3[I(->dFe3(63J_(.+#0,A>
g;>(?[HLQH/>f]^#>6f10M5-[.Ka:JS:)\.2\(92e(5CQ@cJH.cT?PdKFEWN8d\G
^\/R#5c=UNS>/$
`endprotected


//vcs_lic_vip_protect
  `protected
LRfWD2GD0W.K@23Rb,g][@WDS/(QRd]dZF]f0eA>ODMe/ZE^S#,[6()N+2.MTfF<
eXY,X4_0\(O\2(0a]f(+R]:DUO80I7Pde?317g<-4W?]LgO:Ba44US_7Fb5EG8(@
,#dA\4Z/NGG3F5dRE4#D^I56?Ya5;CUa9B,dg7IZ82#H7P0^[QgZBUZ9)R7;_3Cd
?HKagg)7C\6ZREFMT0O=Oa_66B==76Y;\8GFBRMYgH[Le+,e1L@S]\HX8I90cRL5
gTYWE<:?e2DbD/^ERFJFbZ9B28dO<eIEZB:g+01A[-F34N5_cSd]C<<S64^E.<d)
MKc)gS:X]d]f329M7XNT=;G@>d\M\e@9c+H.0>Bc^eWA18,cZ0[4XQd&__U[+Q,F
2MC\?;_Ka_A@Me:7cbVBN=P-N:KV)7>;>GK0Deg,YJcfC4adPbKC_d8+(6GP?VMa
H<H;B+\3OI-+M+B60ec\61^CNZ+C6>#/&K8HgI1&\(>DJe=Fe;OIE=^-_=_&e8\F
+aDC]BO5P0YUcZ5_d7TGBTZ(/0=gWcPa0W/F.0B1:0FER4f2fA7Zc##10,9S^Z.D
1fX[Wb=NFfcR^.R_=Jd>d]Wd/XDL:?4Q97(Y<UK^?BMVU5YHMD.+2MLLDV<)\eTW
(I[<;@DIdMd?HYA7Ic1?5C)fQ3@\M>3ZJ0OUM2E5M8++72=fWeI<Jg=4?;5&1J^K
.We4bIKLP_Z?^/T^cFS_V.U-V>.)a9OI/XQgB/7AR:-0C>T,IfW_G\^U&gIP^M8P
dcKV)QY=g.0Z[<3H)8@P0T[9SAK>_T8LN#R][4aX07BG:ABXQ+XBUC&<.Fg6OA3,
;5g0J6fWIdVV5a,O2]3;AK7K.?(1C5@+,U3[D;IH6JdQ^>H;:,E:,.R9=Z5F;+KM
I&>@2:5F.QV?7[MUK=2;0)CaYQVJ9:Wf4AT-2aJfHP?>0.=\7IBf7F/9(.8e&OU7
cWDY7]5(a):AX\O?D<;JOaZOC;CCaO6DFE+CCC_&-bI-.6/[C@+4\TM?e^;+3U^U
LE.PGF=g.^X[Q5ED3)\22WR[>cVQe+I=O>4c;MU_BW(0]\?(g/_c83SAY\DW_=-:
OD,Wc)P(NE1)H)K-^Y>SC16+:?N189\d9)4N4/#+(LKM53e=J(V+N/>#N;=P:+0d
L:#<e1f#c@#^<f\^-4&BP:RAe6JNVN+M(?O.KZDc,5H>B-4.=&7d<3124cGTWIFG
C1cGXHQ4dH_&Ob_7(J.g\VN1#W(aG[a5-afB@.ag+O1(>7?WR_>3T>N2,A9I#;Sb
)5##F[<FQNN^2fgd_>Cb]-C(XN6W^S#O9RLK^Yg4bXD&b<dbZ][>e=<]0KL:QF&T
gWDORAB-/?^6a#9MJ6E^7[T@9M/1I<&W:E<:LB_1XSL+:;0e4G>VQ;(B+VI9#8QL
-7A,([2X-=/\&8Z6bT6B2CaM_LI2)B^(4887KS;3UF,g-[^GI_f?bF#NKSBGBH,L
#>M4#e(^>(ZDeaeHL.bLd&OI<Qe5:=G;5_JC#b7c-),TU>JBN6d1e-;Y2+]dG^4G
2(^fMJ2U5=7N<=WD3#9B<:U=.(aOP@=K<bb><I+M\[-.FC4E=VDXf0c+c3+fO7V<
AO9;d<.:1(F/D27e\\a&&)62g0P9JEK]c=?ZGU(T<aJbP/<A^#W+f:4b:XV:EL+E
B?e>C;>b-<_:W\0[=+ME&98OZGHGfIg3?JC/\;H(F;FH?Y3Ff[^g)XWU8e-<A^-M
&c>5/RA;Xd4@W16>MKRC.9Xe;CJeR_:KJQ+1#?HI]]B)5/8=5#D+B2eeL&-/#CNR
d13b\F7(cXCf\6ID?#Z?H48]F8\;c8FVJQQfN</fYUK-./ILTM<06EUC:PP?2.SY
Mf4-1&;A[<:(K^g#Q^GHRFLM&5dIW7bc51P^fZ5_9HZR]cHJcA?XIH1SZ(ee4SLd
8&2HBE+Ue4B=71VgBK?Hc&2bLZJ6XU@.MC.QL)&DB9#TW+9R&(^#)V>-L<dR,]ZQ
6d8fTI25_[A82606HB/##/NI+4caND(_b._1]BR(/=f/1FSE96CeX=ST@)S4N__9
S=E1F,=V)?4e.=G+ZfHD-+1/5MRfYTBZ9^->C#]^g04_Q81B14DK6O?D4+&b3=M?
4IMIe9-Qb(<f.>3&dXBQM.I#BACTLVK2gF,gC9g&W>#/AN/;;Y\=^XdMQYU>-2/?
_R>.>6M9,\^<,N;5cXCc(UJZVV>:^/X#FZ:ee&+fYb4DfCN-:6F9Aed=FH9Vd/^N
Q[[[><d&Lc(+cbe8T9aYbOd:aGF@/1)gN@7.944?f\;VNW&5J(RbFGBHaK16H<HN
TJeLD-ENf29#WNf+/8>?)->dF.KS-R5]C5X[F]Rb:8:B0E-dNdF_ATOK#VJPU-H2
F.>\]f>5)22I;HT(gG)6SC<TTSf4ZFdcOVFE&R@/3<CTW:gcTb.WOR_Y)U;>cE\9
M/4c_0O5geT8c?.CJJK@]4M-)@27U6>^Z0ABZ<c?UAF(4eQ8ZHD#,^-g-e4XS_CV
PTSQbb^AO]IO69E4_9=>YXRTQWD&.d#G.<3X0>Re9b,)KW5@VIU09X\4ITQ]5/SK
c89(;BeQa_8/BPDBC.f0AGR5B./F+K4Z?\:^REG?K+JNB59?0abD/S?gA\-f,H[I
_PC[];CG/.@7?3e2\DV;d5CV)361\M1@LZ>17b&VBD9CdQB7:bL;F4&_0fbC^,g8
S0]80VD&b)be9RV3]L\8XM>/V4)92/WG;\a9I;^JHBYKbB]/,YU]fP&354/K(.1\
-BaQQEPKe>Jd276M41;)\V/f.I_Ac55f2;d]UG&U=>:8UN;DcHV+#:5OL9;B[U7g
^C,[CDH<Y>c#R?M/9P,;NL=,H3F<N9=d6)L#gIV1P3(K+X?UIf>=Bc/(d<d?L#B_
]4J&WAR7HB:TQL@\[b45&W0OD@e.<-+?@=,W^M2+/)-/8+ZF<0-;O2NB<&[4&(^b
D?;=P#dE;aPEe<#?Y8ZKI?7.cdWOUU=A\4FNR39<3:X@D4fPYWC8AJZ+PJC89@SE
6?MB5W2a[6I:E;/R10#]E2TO#PJAUeX3(VJb[XWU;DH:[.ZBg.R?-&5&=MMSRHCf
WW#FO6QgX&P5=:0C)NJD6S@3,P)AbO<LeeJCA=.^2^(c>U<\Xe&G0BWR2>&M4:3T
HbWb^E[#ae=G>EXGfCDfSK#]6)^4\;_V5c_6-&7ZS-^J;ObgK.8E[_TbJ:J8XG64
L1L9HB:OfUM0[-(NG.3N+Y4;BeNDg>8\;b9F-W4M]^7^XaQESA<8cUPYUObZV6RQ
CCaLAMRB13DQ>g6V,@M\B<K:6;9<.5C&[[/IJfZ(]&XAGA0X8R8/gE57\(U]206f
,I9,-?V&5O@5XDb;fW96R]f]EP0eW_X74JdH,.L>9F32eAf>Sb_SA/#H,[Z2]L1_
4e[A4.C@3EN8Y\5+,c-=:X[K_RK6=5JVT+fC&&HaFSX1B<_a@(R2d#U+AP6:H(;d
L=9b88I[9aY58/9,?\]df=T.IP7&[A=+^V7Q_:B5dD3;^[eY--GI(6B6^-fDYLD.
^9FO(6FbRSLUE3e549S2(.F+eM0<\QNC?@g)#EIVfURZ0X7gF55/<D/g@1?e(#5F
;.+L0R9C/7?@0#.#D()QIU0R:@<S,f\-J/<OU2aeI(WK0_WRUG]W1V2:QN17:,/N
N]ET+XMgY?2e9A/-]@2>E&W])3Y#KLW>D5LY,gW/BV=-5U+0J+]BK\ce>dJMT@.&
AB1Xb,FFOOe6/>C=VYdYG-LY)V6]MTDcd+gc/EY@P+6O3/XF6GF8-3?);]:H/RSf
_BCP5CB>FB]3,H.Y/02Z9bbN3U6W+@W,^9+P[/]?b;R=]3Ice[B2-TCC)M@NI:H4
1T@UfFK>-Jge\+Wa)d.U>1g>HeA..1@NA>0gcgDPA?===0H0=?KX\10b.45XLaL0
1=2WgG4GD^g7K11)Gg5fcWRZcef&=WW&736#R/6IQN:PP^XU<[T?#GbPD]eb6YNH
/@224.]ZJ3.L=)_9L181d9f@>gDT12;IEgJX.YEQXG.;(31cbPeFQL\:&dNOHD+Z
Ab@^e-N;X^J:aG0-9]a4H@E[d@(ITQ+]Q=+DP[R4dYeG[c<2Ba/1)+&fXaTf[79W
AJP7A4FLU82d0);W\#IOZ,O(F)<U8NQObJ=ZEX(A4UFG6VF<^24J+aKK2I9(:(E7
6O5@H2^<N&8RI\L?RKe-7<9d&<75/D)9P.]MP+4#AFE[\C-O9M&;Uf[dCKVQ=?+g
8abL?B8J8<WTe,6-R1\C57]PGdD5CJ46dZ>JZ&H]]IB2SLOG5/,Sc0Z>aD9XX8>A
60N)EU9@Td1K_B31RZ[17fCKECYNXR\9GQb0-Pc).KKL)TR60TG<W8gJ+>><]MWc
bV5FOT2:G/\63ef=JE+L3JK2K=4/@&TSLU;MM&L)e2D.\fXG/;5\RBa_H?bBK)EX
CFQgEAMR;eS85QLDFJSN924>VgWL6A]H08^Q/=SLOWOX&#]P>6Ia5;4a#)253/d_
c.)b?CF@9T(5#Mgg_K]d)IOX)A]>UH<,(D1/[b;f,@+_d5ME>WG@LJ.&:8OW(VIP
9ae:HJI.YZMMQ:O<e.^#(M@cNW&_a2Q<9Q-K@bc8MBW5UcB6F/O@04,)J6]Ug#eM
OTR-]##4.@cQA5JV@<5Ba<;UU]=G/;DNP:3OHH[eCbWE5</3;]ZM_<DJZ>g(V)e3
a3FAC\LGVA-9K@#cW1SAaVXfbgFO1>f1c79Y>D_BE3_gI_W2H&<FcLL&OUg,dX8M
ZaF?R/d=WL/_Eb<YR1U\F7fcFU7A^];LCK4L3H,DA<5/X_V.YWNN7#Z;D82Ya_\R
eSeAXe\<DZbbc\aX5#X<B;ZeBLI9L0]aENDF>ITgYK@eY9CXb<REGcTfB#Z:4Y5,
3NJQf5Z/QS^7&DYWT-M.QJL]S<;4<f&3Tb9ASd1TMWOS)_DF,4381(7]2gN.<VUf
7&U;af8-UZ(V0Yb&^g1AR^Bda&_U)@M;7Q:H]d_?\IdK#SDE\)7I^90<[,eX47W4
@ZDV<dMN([X<OP5eY=L4_MMHR8\cICBEAS,7>U)9c5&19<EV/A_IGO#XcWL[C[EE
OHXYgS-W@UJX(PKI;O221:/cIREL8dQ7gaCQ<[C;9Y?#,=:>C0<UY)XcRB)9E3_A
E?L>E5HIHDKW(f(E<(3RX;HX4LD5XLI#B9DCbU>X-Af9V7-D]H,AW/4DSeB>^UYc
TTXgESOA?QZ0dd\.eXOU+#HN9c/_V-YSF<LI&NZ;-)3U>7e(E-H>=-0\0Z&,Ng.^
3aaS7+17,@;Te4d^(R[FOD;?-?GU4eM(Zc9@L<P_GNQHd&4&K=,)/[86-)[KCHM@
30T]b;,6dX9?>d[IMNCQV4)[=M[2KfF,RNGSVAB34Kda3(9e32T2\Q4.X?.DgYIS
PKV4I)A^)eM[WO^gR;#S>1Cf^+FaO^A]^dg->3Y71F[B(3#Y2LEY329]6\_9JH.3
,5Tea4J<KOYTX<.8=4RX0,K?;R,WVTd6PXf9KJ,/+G^D7YC>8.4+g5XPLaJ58,1[
,D3FF=9ZfTZgNO@?X[/IDQ.aTSB;EULA(085]Ne8T<IVMFRHe6WKg6(54R\@M+0X
I..MCa>gSFUH]_B^(_7-G0PBZ:c;D\eRSb&EN4fW@ZVBYVOQ8]M;::KZbc=;B49.
</?WX=b)[@>g]D.FaT)=O0G:a3##MSR3eVLX>e)5,_AX)1D6YJ?-<7_9#\;1S]B=
;_FYVRNBIA2:&gNU?eU]G[+ZgPIEc]QD,OJ:>EX38T?KgWQE9e[12E7a:bT3?Ib/
]^UN;IN1&01^0NJ>OPM8Z_>3(O;/^W,ObKOO2XU,LORV6[07WZFA)CWb4.^]P)Lb
&UJ?A3+7_F[B<MRKCFX[.Mf-c6_B>2/>RQ(c3PS3[_&\2d4UfF\5OFc_)SUB)<8:
fGdC<g:C3V:#Fe76^f9JZ&g0aT)XH?V8U],9F4)GR=8)e]L&-1Tc9)FU]=WbP\_>
777B)>d#-Z?\NXXWPcI65CZ+0XJ:8=E27.1?8RC#+&fVAN=F2d@??==556)-4bJg
I&15Z,\[AZ,bbK=9AH(N:?-4e7bC>U+9RCHSe_JF(([FJE;)_/]#&0M-F:]2B4VR
WWG01OF9:Q5&__+R4f&bNJ.6/T#BY[1^DPT+0BeWC=bL2;AR-<K1Id-cc3O;T2bM
K>\]VBW^C2Ic>IW;fN>ZJ@;K:fYU&]II9:R?g)0V;<5K8eJa3\-eV-#O,?bJZA(S
ZCgGg[+eO>?O:>E8><G/a\Q-9<PGG.^#Wf#O_B,Oa\OAebR0YfP88>_\[VF7J6aA
&R_+AN<+a3LSGUBW>@X@VAJ;4Y<C2HXbH2QAI]^b_,-bL2f<<0E69<AM=5-(P9:J
R-F<cA;c8FQ&U4,5e)05X.9Y>(&\4;V+c>?Fg+Z&,9VM-:P56[C(F6Bed>WTLQV>
]Rc)6KY]A6><L>N-9\a0D/:6QR4>I]U;5]OYd56V^bK9K:V)6aYVYV7:C#d)K\?]
X56<4DJ)>2T,2?JWBJXUg2N(0^1f2c8-=gGOTZ(JH5/GXI<@fTEdcFZ.4_H#^^F0
PXN=[PP4/(J@#/Wg^PA)(#Xg=(@4HKSPTG8/0^-Na_S^A3H#c3Y(+]>-b[U5SZJ)
HHQT.T],8+P-TEFb>5d^XOca>bdKbH-G).c4Yd+6KV[B(L>D_Ra^6QOY.XR?P)7b
G)X7&>A#J3A/POX=/Y]O;HKG?:X^24^/f[/S,NS<f4VH9\a)GQ9Z7]&AT7b+\2.0
HVWfC3g3XXGVENL2=.^6.c=453N##HVAL,feJ,F9Y,1QL3a(e6eM9GP,/?X4?ES<
21,a-8Eb&fQUdSWXfYcWTC39@2W<.OZ_IZO7GM&>TB^O&FRQ8aK1PdZWNE0^DL3+
WH^7MO]LP->,>X^O-0\SCV/U-X.1R=2(2,XC/<;61T>d1.J/A-P(3^K8;)FI<>_N
G[<LLcXfJgKZOQ58G6F@gg0S\W#(GZPS?KR0fL)Y;C;I/K[YF01bA59c_bF/6#G=
H)GL8(<@(/@EPJYfD7KL],QO6bS)P6I-</2X5OD;gQ<J8V1H6X.#RG7-I(_GS7YR
PZPDOdI=QE^_PV\Ga_6LY\D74>^)D=b.[WLIR8NHaU&7:0b3RQ9_HAQb=[,)fP-8
_5R>I=05A+H^0dO>3.@,,E(;DI=aIJT&)/#eD3YFXM0FI]HA7XVVY\9)fI1bD..L
#]FQ\@6d0Q2?A<J-/WB1@QWIR(UF=2c-?^4(+UU77ZeIJ@,3M9OHa<_Q5YN3Lg@;
QbHN_3f_AL=\,:[[#L)76\7^J>XL&g)K)SGH(c)-)]4).]g:Eg+BDacZQ)+8>>>H
g^OQWfUbY?\L.fYcPOfQ^(5,?1I6^D33,^MOPXVJFT89OEHZ.]04.4KaM>a1D<CB
/]0NYFY,3XL#-+GXXSW>KAZ2=85H@#gc)@b1X(5ccBbN[N7Q:Ec0]4Y2-I/=H^98
b2VUU(X:4E8K#T#I[+e.M?=DA;1=<IY:ZGR)dJV][JE]b_He7]ZS5Q/VVH.3]>Xg
6@c)+=Z;3HWXA2@U/23##f>b2cN&Ra&2U]4BNE;N]DD9PAM07Ue?02UT1A[:\bDX
Pb;M(45P0&GaT4/d-Bf[9@<)TDN=\CE0MOaVT&ODafddW>AA4P+.8,a15BdS.[=>
\3CaBQ=RcBJ]V3T(/)NU<<RW,,L)d78f\I=P54gV(W?73.0J#)^HK>NBEKf;8#PM
ed-JH5:/620//=P+0^UWSOba;S+;9g#\.(<d6QYC+C6G20=7g1QL?T^<X_]5AOI#
FP<D:9^\>C>+4b8_&XSGYDI^]V6K;D>_/d;fR4.J:Xe0F&aT--B9E;_MWZS^S8WC
Vfb#;<T<S,9__Y4;AUPPeA.dKc2f8A.\?PLPY/01+0:?b3T(Mg?(X[W82EIAE#,Q
#Of=1_-faABXPE7LY.g1W34O;]B51V3bE]]7?=cdW+0YdP6A,[6bc.YXL+d2-(;-
b<X#b#8I,/DS8>e(8P5T^&aC&V760I@(+GS52HIg+b=\]\+8f8?GfT4:Xe2g&B;1
ELRC2Y.A)L,(6R_NJ(DF@?^1L83,ZggUQcBZ;Pf)UXb5QeT7L/]Yb&I6IV6N[;(P
C#YbZ2\(NF6aQ>/Yb1Fd5M_RK&3eb?JM4HLGPbAgJ1&>(-0AT(g&&N6ETP\4\;b-
d[40=12ZIYg.XC#a><+cZR^XA\NeQLG]TSaHf9Efdg1,HT#gOdK+a1E8@061a0fW
QAN/H+bGL_ROI\f#1</eJ/8]@42@,(P#Gg-\N@S^<Vd;Y).b6\#?J0=7U0+WOSA\
Tb7]S<Q)EI+&d\(,&^;C8/TWY.&dVLLPS:>6^TN])N^=]XO)M85V^Xf\S)@AG>UZ
+@CR7RWC4fN.cfFO5CcD/g+E.P[7=[AM<\6W[HVMfWX,(33ZQA=R@eOIUd-Eea).
T5cD4^,Z8923D@L<-3IQ,_dWWN8#=77Z=PA-Z3^DN2g8V:&>B.8N;(27=)R2Cd-H
a#YdGKW]1Td-V8<2g5a^;8MH;ZEQ7K-)HbQ^0e^B+/dbdJXX9&KB147=8GG[JN?D
2WV_R&A2V]>LNAZJ>-2=1U@/36g.^[,=X-V_XZ[RKUTQNU5=U1=d4f?F,2X1gTTd
.WOa:VeCXJg@=(YHQ48F[0^,HW,EdH;]I@:KQ&0?X+UH/;X0#D;caWb03NR.a+EQ
f+-^#Y8P#M9#Q.[T,_\)W/SP?RWbN=@G<&6ONXT2.^4^QdBPB+dI]X4V;XLC.@<[
eUYA==XCf=<V;\4]WJPB2Y9IFaV;<[,S^LB[@_eb\c026TdT]g3T@F6O66:S8MV_
N9EFU<c>c@N62G=e[fd6T/^8OX1Wb_H,dR^f4VTRdG@SJS8ZN<4M5,XVee61L&.=
@\@O\5[8[,VPe<E==R#[?O<3TH7C>3/aQIW\VKg/AQa8055U?C1#<YTEf]TG.6PB
,d6?YU),,:^]O1^0L2=L?CY.)KNBEE,2g\5BGdGZP5)8,2TK7XC.\:6HK5QE2HOH
MDNSZ84f3LgO0W(YC9NOB]&:.@#eC;MeTIe>XTeT@3@YTb#9UGOb>OVT:Z><?3g^
VGF]MY5)>DQ_KEA8RY#A=#3GXY+,KdSXID>+[E\).F8J>:.#ET@#NVbe_8=Ic4gL
b/;..^Q(R9?JAIZ=dJ#EMg65&1egf<7=2079X23OM1I1Q=\.>5>M3WeZ0C,D8g,Z
_QdW&1HZ18c4\ZXQ#=437dIS+LI_1?UY10^-M2+U_S=M)90BNf)Rb3e]gcE]#-g)
2L-2BKf2VNKbA]AaGMS+N_T[;OR:c[=8f&OI=83HKS29#aM:AUa>;Sc7&T(3,.5[
@-L@)^+D/RRYeX@&R[dBC2O:5>,Kf6cTJcRRB[c.O[M6@gN,\.(5X\3-UPIT8C3,
.6He/\>6Q)#fLFS#4;8,=T&FIE]82NN?0V?0A=?4Y6+1UPgI<@H>T1NX2-W#fg66
4]M4WNU8;aH?.LSdA2dO64OVA->TfU<<:?\([=EW39KO9CMfIV+_O&aT)aDEG23^
;(Ee8-:MJ6&LNAPFK+IRH9Q1<+\LT89Y5V3O#TM<=@UDA4Q]\d4+^[fKHLf-JDAU
87EWe&1I7Bc/E+&d-;cYMZWYWWd\)E=CR,,A#4RM)FfIFd\@LT(>CaQ<4,:g=K?\
E<2]5c,)[eDRabd0^)@-.BL23fL1;eH3BYIE(CM3Z&_\;OHbE7e9YY5EQNK=g5\[
]<NCL.S##aPU?<:<OF)ZJ2/<Ca#55^<;[VDF3,NNT:ON?MbBWWa/V1(1d/O3^TR;
=e7S,\V5Ng;Le6,gcM]#E(:,YT_Q&#2NgPDP5H@?f#>B:.M/[.Zg3I<+BU&[4(^M
eK7Y.P6;E2=YbC71VeG73bJV[)G/\C,2,<dQ_SHQ./N3BA?c(&+]QA5]V:QDTDP>
B=@,,.Q9P/3>O-B0K0S,.CBLdY).7#(+=LL7a5ef(8Cd;/?TPK<fFE::6307K)_<
<J#]P<1T>1K6ef,&830&S9G@09_b-/92:HL#@-1(#HFd4T1cSNUHgQ0;QgU//01]
\_\_:b?ggAS^\W<c7+cbU/MLLGafIWbd#N9[[Tf2fUABFBWK.M<gb+,KaCJa^Nee
IS7X^WLLY5?1#bEN9G2F(1a_@>U1N:X0g2_]De:De1O5bU3U\6-XMNf)JVVT<E,V
M=OTO\?e4KfO4Z#K[_Q#CJ\<KFfYd/JN#<@_H)M4=IKAS5<4Ne\==]7^.>6[#2+-
])Ja>T(0(O9dA7f5b?f<@SHY[aJH0cBZ,#+E[KEf2@K<MS&EW=J3;DV_2I(Q=g+O
\IU041cM>N83R/F@;=PLQA(E,O32)LK@B5F22YW;:J6Q45\Og/J,dJ)PQQPbPK)S
gdGU/TI[/1>XXbe[#H8<BDD1),7O.4@S?.cIYeA4\Y,:H[A,^H77E)1e.1e:92Q(
:^(Gf8Q1OY+1M#g4)gJF8JWML7M_(MEAWND&R?VABA;:7:1eV<:CQfMXL3_BSWSW
_+F-VDEBX9R<7VW@]MYYB;bDBRY0]#8Z.e&K5Z#SEHIN\W^/B2SS+7XVB>YBe52Z
WLZ9eD@NX.<cbZY,KKdI6(Qb&f>]-]a-HL:+TIV9I.RYB<&g0GYMBHdE1B_+cGX3
a2Q^A/Q0\d7>?,@-c(3=+V6,O0<5=0RMDMD#dG)UGc^_FB)/7Ob6IdIKJA(9f:d=
N&KPX-fW3d/1J\fBVSN)=aAJL3U^&)8,g\BG+c.SKJa;WbG](4aK=2O+]KDT&bT6
C/6da+f<Z5TBbFg,A63;,9&1XGZNY)0Z281DIJW?>#3FH]:R6FgNPG5/252gc8XC
+[00ZN;>gH,Yg\FU;0KH_K\ATN,\a[<JR.TB2VRRT][9fH68:T^?(\[GZ@ZXMb^+
N)gb+7X(13,K81BJI)]QRNT2S_ACG-=5f>,=T;,ZHOM7]A)@8>Qc3QEO^V7LE(@F
BUAO/-f5gdY)E=F#DU[0^.GZID-.+QcaMNDe:R:De0\b8X>RPX>#QBU&.]2DTC5D
/2#bEK&]aBg]0&+2R)QcV+f=\3:?Y5PT[7=]G\U9)LeHFO9\+L9]6=GfcP0:6=@/
X5[:+Y^LWDIDe[Vb728:].#acOR-eS[01NZF[R/5T3c/JYR:(I]&</L&:cac@e?E
D[9_Ig,B/6S6_IVb-QASY8/AC6F(1VKc?]W\^bVZBbAU7cMNNW2_dUJF@(\d@:<e
67Cf7E2?E_36e=/82IVFRNgb1W0+37:97c+>N@5AUIX1NFM.\WB8LV-5R=X9B@]M
G9+V?5+TVf[dVG6,R^T9/4\J3HMD^S0LR89_E-,YRbG6F?2[\O9eRO4;N\?e&L7(
5[1JX41#;.dA6F:d:MQ9X#[TJS\<L?]6F3+b0bMBgf?3Lf.9E@JV_9GSf0OCFD_-
^:&K7V);^OA)8gH\@Ca#-WSC?X;@(0c1(_X]6H4SRHU^AVFNF<Y^P+/3R,KM4VZ=
fT@]#][@@T@M<U1eO+O;R4NX_CM;L::39[+9Pa]2aY9YVaCG)-&-2aDN.WQb500@
,7J/<E2ZVDA_Y5E1Tg_QJ1LIYUUJWPHLdf8@=^)0?E1^VN1MJV4GWIP8K2^8UHDH
WH(J@6Q#DP-R0WH&]N=g_aEN_Ye_IUfN4F&@R:a@3;/6_.75[,cC\,:N\O84G^X8
WE3A.DNW.74[aPL\&cET\@TY_EO&#IW/#4G.H8@NT)?@?NEG4<Q9a+^)g&5J0MA@
V]Ne^_f30RTIJ7Lg=+dMYVVY_>BLS=gdFX+R?(7@/^GJP82IR.eH:N?2D1aQ]0&N
9))2C=fD]IJY?&/G\LZ+6ZWT6^>7@MH_[94IaC)8W-[B^<]DK&MDT3\H#D876G=,
^G?DFHHBBPE0&ORSH&g7RA,)[V^D+D^IU6DM#QRYG\g[-&GI=+Y0(Sc<dg[WEU06
A^:GAcTXCKc+#/0=ce+?<X.EJWc?RWYI1=.RUU\KI.2.OeB32^WT82+Z0d;-d1/f
CS^Z<?fNQK<DHQV^49]B?F)56YG4&Na:g>2+JU7JLK[7&c0(03Q+B^EP^g,RY.WW
0UP2Oc#>3F+QdKb8\3<GESd+B6g5BeV,E>CdUW=,@URgXgBQ.SadCS@)QgQ_[O6.
WT:-)RaDJUR;Rb(2,UWc^XF8G,+NKK8#eQ]&G<F2@;FIb8bSE0<R]C8;eG7RNg;(
2g/;YNS/fGEg0+D2@67]gP>V.);4=1b=L5D+d([21O(A;d1QASANH5(aH8B2H:9X
#\B-8fTJK#3aDV/J@/a>0:S,;.FSGZH^\55bZEBD2KPd+:fG4)LeF@.3D05>/.M#
@842CR62\RR><P^5<1D?VfCUV:56e+L>=A&E>8UZLD-&M-XRTe\@;3QY^FR4I-QY
APfbA5IPZB;2bWFa//05TE8#?[UD9(^NV5d_LAc()P)8I<;L^S48P=?c?OBQ^BYT
e;>#3EU)L#GU/)9=9g7[(O#+KIG@+637U2NQGO;N1gcT;A3#IKg7V&MPK#I=^&C8
Z>16(?]e6@T?#?C]4<feBA7A5XJEX04WLUCKRA[NPG&_F7Zg-1EQd[=E?SF<OY1^
g;7?gGPU(:W=WD4M35Y.#6f#e_)+c0^P=>Wg^RBXJ<5#X@\7Yc5M_P3WTRP17^9)
7dbI^__(&KD1L?&G@f3>^B>F\7c99/XgZDgJ7_52-E07UQ.OYNT@KIWc:DgWYZ8A
2-WZT@/L?Pd8&WY&9_VFJNc.<WH.be?S?CW__D4N/(J)K(^1P+1\6/dd(\?ePVG]
^,_/K9P7[2?DWH_].?f0.;eR/M>\;8KX1I]6ZN([W6[fA<8A@#Y/aLN.+X:DS+85
SYY3BCRG,.D;:JVS/JUaG0NaO,;5B8Pbe9D?e+@XQ6MRZO=I[V@F9c?KSP:6WZ/&
A_d@WE6@IZ/^(88P)@F/<2f_8(HS6<EWLd=\Xa5XJZ5DG@af9.TN3;BRc;^-]?1P
;#09^@(S_eYYHNO+X[2Q)X]^VBc,1.T87^d\1U/CPf3=f)K]X_-B)ICJQ&IAK/DD
]_<WD-E8aacK,4[ZLNR#D]&+Q2^7DgcFACW\QHG-I1,)VK7)/E)-6fWMLJBWfITP
#SUgP@:A.@\/1aZdUKZT=U2TXF)Z,Z#672A@/-.4;<PWaW^3)BaYS[B8c<9_[5\F
)G=71^\La(;NK9WB\,382T&D19Ed]g]OUf^JD=?F(7H.gJKEBUBMA5NK==(_TW.B
^/:6#T&-Ff/CX@S.^I172Nf_eTD6UN3/W>+2;bINLR)P\W;;DKP8_]AIFLL&7XB@
_))R92aQ&YZ7V(](AUZ7XGBgGJD+_(XV5_-QF_8@Z1/[/B\<:#0X,gAJGE8_O7B_
5/K4[8@B&A=^J,4+ZX+1ZCaMB-d8Z/OV)58(U7=?IadL8efZ.CUXFT9KcX)M@Sf9
;T1MZ[<@->B_@:a9F2Z[9RaG_C&MfIA42XFR2CWOF56deT\[b](g@-,&:1/e)cQ^
7QW9R2Q:Z3e<SD;7dFFI8H&9XD8VFF>V?7JT^S35+F9^W_&f[_36H4_O4VU9-3Z<
-=7Pb--6H&.cBI2Of;,&K9.-_FO0BNGK;VaTX3]bH2,S2CJ>NMNR-VIee@Jb4#FP
8#6B(\W:)=3BB1\Tg;;UC>.5f3Y<9=9cafGVafP4Y-T/@WFJEA1TAHVD8e.)E=O0
<+TW45X=[Y#YEH(SD@?>fc8\(LGWVg>5+3T>Q\VAAe\GQC^;b59F:;R-=GGd]-K^
+Id/-VEdXVIF7OKFOa3WEWL+c.MP1P:&]+]4b);WY\+Pb,^LP\7KJ8]..)7>BMN9
57#P4))7.)aJPM]0Y71C;9+Y[@.:,[DX;EMMB@H-#)C,UO<>ddaL,M.Ga+GYa1.^
BYT8,-G9K/;[GLFG4\H)TeII9CIQag:R>WC>9SLa@L^M1G6Rd8)BffWUIQQAC0/f
45(.3;PUJPIW[7<@.@\BG/Q\5YffSCEPR+TYYaNH)1\X(//_a.@0Q/GMU^+B6OO/
M<DdYg;GZHAS);TCS@&((]gea,/7OGKVaLL@CGEI4I[224.[>JO&;TM)/D9R+a0,
U_[4<O=K_BM<E3Rd1c:fP(WcfgaS00),P:+2W)XA=@T?Y/aa#\F9fH(&/UAXVKe]
G7fg<9+fPEHeJC<SBM(;gQ(5UFDBbFC:X\_H03:#50MU-6YO8DUSZ&J10U[db&XM
a9^+_#J3gV;<:#-SI&QeBP9,[S3BQ,U3e,BMH5.B-^1^=^Z0N?I[C^_VR-R@+L:K
N2cJQEF?/<)T.RC+_O1/-:UT-a/1S-cC9QT5,8?C<3]6cMA[-F3f>RFIbd0\RO/_
ESbCAATC,WNBH_G/ECSUM23-I-9M1YAaV&)DgL=LML9gWa)9&N,_8ISA/4398>S_
Z)JOGN\+VXKg(bZeZGbY=fO<FW?J(gBG6_94PD.AAI;Z;-9J,U,Ha6BF,+E^;b2d
,VTA#Q^gL()QXGV6/;D#>D<,bBRf#a8L6]\M+4Oa855O7,W74Be_-Z>\2R=;;7^7
Q,71>IYF&.+\U4,c7#DA;2U<EcH7?0;_>6/0]1O7?YGRf:.0Fd?WJ>6g5Jf#3>,N
&gaK34IQcSdN3?ANLQ@:Xg:5^dA?]92/H;Bf7+TLN,-8Pg8W(EV0H#W260+JGLKW
a<FE4TA>e(X]D==/\<0g2EHZE+CF3FF7:e@C=Q@RFMaUWQ8ZK=Z--#)7AO@40\_]
B/)R:)d?I2JZcO^X_bC]4_=LFJDU2F3BG349,/Q/(H<1WZ<BBL=abVHe6cfS8fSU
J5-HF_f?<cW[5H/:5-;P[5BBF5MZaSAG?>(DK21d]FL0#dBUNSgg/b6M/d[Z[:G]
?W>CTRCWD)N?ZHSVT?1YK5&<b2Pc/DS&G^D-<20BY?:U6W&[\cWG]QSS@U4@^\Lg
9FCA&(?9FCSMZ/S\:XQBR+M#.Pe[=S&ASG;Mb@]f<J[7=M]61YHc^_gL3^b)&\_R
8.TPYH8A\></-#A1:3HZ4XMJ[R,@08N@Q1g(f6Y8a0/AFO_8XPSbQJ_L+.+dE1c_
eV>X#/-5SYHJC6[e&9b#NNK<4?M2FMW-V<)H7f#Q\6YNI:YGc)H4EFT2&C=(R/1L
dKH;42S]b7H7ON5)3O.YM0cYLGb?8A-E0E0W?e7E[X[3fL?@L]/c/@:a+FWX+8),
+eA9YaR04OE(]g3M6f@:VTdCX3R84RcE6fMA.70HJ2Y)f)3cW&;A^7U\D(M7HPfe
4I3<.R(/UcOV+A9aW?((We;I]I,L@-[@>ZV<I:=.PYM2+6@8B0d44ZWEcW4)=H\P
8>&U\TX.C0:E[:TR/cI=a-7DV,NO)EUQbENU01Tf.Y4U3,1D<A;,WASc92^2APUC
D,G/0DT9X>Q)A?T704W-@)L(B2?JX3S9J_]GNBG9@c<T?[W@1O?3c?^^YN?NbJP)
,7)EQ+GY_fgAGaDc(381B_Jf#:OTXc@fZ;^UZB(cUANb[3+:fS?V.QZ?M5:5DSV<
;Y&.^SNLf@RBa+HdTX^LINc<:B.F89QE+Fd,YF+3d/D+dNa;6,eR\g]QccN3/G+b
K_>DGe&SSO,9)S[e9[eW9CbT>OJC472HH=S)bPOM^2Ha4=LL0HY&>>RWBd0F/Fc6
W5,8M^fN?6SW/<-Yc0=gLZRf\gPCe4Xg_=XW<)b7a.V5+\S2C60_OL-&5IQ@19,A
IXfS<&@3.Kd+&D52ME3K1<)<(A)<EQOf3+LIC[[/JDS8=b9C_?8&f[,ZM?XFdbTg
?[V:(M_]B^4Y#aZ#KTTW8Y&2FE:_W_cPQJf(7[G)<F@9]aH0J>g-:#33g>^eEX8M
6O\W(K#F.+OY&\bF=_HDK);-9P18#WI6T<Q=)O+Y_fD?F4[CIWMG.\&K@D]3,FD3
T?0P#3KC9S?43b9H\.A<2a[2H13EA026&J@:&/e_W_GgVLgFXcARZ7+&T,[:@J48
O5,,R+N[=#SUU[LKM2D:=_#1,>^]EYEdE(a1[E-;f1(Ic+OR(\RfKRKb^><Y/4[g
O[KR2aI:GB9Xa^60#@CB>9WPBH5Q^2=5H#9NR^_:-+2,8IFGVTdX9e.dE/bF9Z2F
5.Db-@M)\,DNdW8APNL:DB5(9a-gN<1XCa6-HG[U0Z3]BB/BD;]C#WL6bHbW=fSP
LB4&B>.9<>&F]S&>a,L/6WPG^XNQ<a[V91RU(If5<:Hd5e5c[&LJKJ=aI=gPb0(c
C7)O]f.fV=AF]WJ196Hf:DT:,2b#N+=D)/IVQR:LJNLfI.F<9aX+_,I;FKEFGa9X
4U]c32e@87?cMSJM#CF6^D.G6.DDaeFEc:3Ef3?c(\E,GH(_Z09^Vc1KM=f0:U6H
#=E]7a]a_Z,8f1]I0K#IBBgga=fJ^RQ8E_TM0Y75W(eT^BV1bAHV\=X61S^8\F5,
#)]1gc<ZdFK=-&-_<8>IPUa,Q@#dTHP7>K_\&\@PEQ>5U9(DQT<<DcbK?WR/5I^7
JN7O55(S_gd,GG^&\4TS#+9W/DE(42d#=E,CRQM#T@4=Cd/.XGGL1U^21:HS/U+<
eH(fQ4(GgPbB#gS>@TU5cIfA56XFIReAD./>C:a_5I-TfB>?_)1Z?+(E(D<a3]-b
fdf(@>[P<D2aN>#KSTKKJ5[8)TC2C92N8TUB?##>L9<R;fTGF(bCWd:#b.><^SOb
VOT8G3?GFN.\d>94:aZOd.#_F=\:J:aZO6--X,/][1bdP,eL<S/T6W?KO:bA=QS1
6::f\4L7UOXeb\ceT++X+,4QK8(fc^a^X/>]L()e001_O<9:#<MRI+f&E([g@D/+
I>Zg\80B>Zd]bbTNE,DLKO8)^G5R\?DP0WF51-0+N)EZKeBBI=QJ1HA&U#V6OZU^
,9KO&;SFM&03U)^;F_eODYHfAL8G0/e2??,-6Q.7M7\_?#F,H]SZ\^1OYR09;0f#
HOd<:OH5]Jd,H3#&=H^C@cP/a?W9AM86]::EKAaAdARDQIHTCDC=@]4,fGTF8]Ad
2aU>Z04CVd4PO,Kc7a5@XMdc3J?^d2M(V1g:?b^.94dL,GZ8Q-d6Eg3.]JD4[97N
UVe@f0CK\S5>]4dTV+b<eX=bPM=VDDMTL:97Xd[WO#8A<\-I]E_Ab=2DW71gY=6G
/^4H[4fQ?URD+>K\Bf?J@Q9WJBW.L)SBLDWO?]+19d0J5)=G#8c)e:J[bM4O,@B=
H8=WJ3=:TIK>ZN:YG1F:Se8EMAaX2^?aT2B?_La6YO/bXM6PQR+&FO=B58JEC.OG
CC9>be@D3;Q#.Hb^,RB/&5B26ZF-]=TQD7)HDbA7&1U4QQcBJ9Xc,L0+eX5AQ31>
R9P0]3+GNPDA1JObYKc9M1abUGX37[4?Y+#;;S-f&#OB[_Z<X/KDOJLH9?P[T+Xg
5^B]+,EW@-KSQOHN&C?aKHd_g2BY)3A\LPLaN[VZb]U[-P\\f>5KK@bg((@77BcZ
EGCga,AHL3ONUCIT4GIG]OSV+BH]?N(FZe^F^8_.UO_P64^H2QE9A+?]LOM/ANFN
M(SHZKIe_dV]6L?EV;F0@^LfdG\W^g2HLgK/W&#M@6@?@<LQE_JSO<#J5.Y4),D7
I;9A^g2e1NYZ0YNO.0UUUGYT8H?P\W&E^JVJb_74YW)agdFBQ:_D;+7]G5J+4Y7R
dA559X#8-40OPF/T=VDS>/3N=/8,IB2b]#:d?@<?aWT@4+P,;B,2;]NO)+7HU).;
b[@CaX08f3DYK2[c4G8I;\)P,R;&g/[Lg2@.,ULRESEN6gM?f2X@_6_V4U,@K=78
1_ME8P6CJV9aL8aDFUNQ<c<F-+Z>J07UJ>G,\2Z1FNWO\d7eYVRg^>UO?8)C;O7b
Sg,2dX?]^a)^>c<b+gfF>TF&4C8(e[bcNX@O.Ye>TWX/E6e91^AT/JQ)SOegXcP/
TP-N)AE@5N#6=4(RTYL1d,Id\W[8VQF?D7DeYL4TO)\C:dQ9D6Q#BP]?e9G?V,Lg
Ta3?4Lg1WO(-8/NNE\NYR^^(<A4=D8J-9ZB(,A[S^F&aO9Z294/FMJDD\D&:X^@=
1aAXfA?\B.X.,CDWdIN,(Y6.ZaLIWA>./IRR/M=:Z4\03XgeXD-?/0dOTdR]B6gQ
)<MK/\NRSPHW0I9_#dH^R,:]3NeRg4Ya(=]J:g=T3\+b78V5[VB8@HB+5E_6aHDG
H0EeA,M;UC?23((\T8Ca/<C,[eF33YXNLWD86M?WaD_G8:7Sc+LKP4(V#4bNWgA-
&N131>LB,[&?=T=Ka9X:4c)>9Y(A-ABQ(?C,&<I6:H@Z&@MI@\3O<H]B8K5eA&WQ
=+=XJe(]\[U#]gYZ[6;+Pa+XcVFQI<Q>f\2<@/^X&R>CRR]VO6L:OCA\H<ec9Pf7
S[--Ofa&GPJZDd)3Uf@V,TB\><BU41[Q(Y9.;IIW&fBW39I2<#T&C2NMUAI]4B[a
bfEV,Z]=MH)Kc_B9\>Jb7CPDa.2Sa_SS17c^\@0,bd1=eL5e582-2J#.##,OX2-7
<#11+\_@?A4[YT=#GH3S#L=]ESU&A<+ICUVN\0VdJWQc9[gKN^-d&E\a+ff7UG0d
#.XFKa(M(]a7+\+S3E3e4E-3M<+P4ZG1L/J9ccF)G?6fV^54O81<P>Q14-AUPA,+
]M+&2Y=1SIg(ES4X=&6VgPSfY0CE;dV),8C/F-a2N&R2(B-+\&OAZ_\.c&a_6b;f
/@2D46aTY1,^?]ZLFCD@FOB]d+19<N\^7/)1AM6,)(3S<2e@V(4Z=]56&FBTNO+d
2RAIbJ=Y)@cQO+(Xa7YL&Q\?+.;K>2:UP7=@K(#b;B]_N)E&Q7M]6EJ/R]\5X=6g
CC6CY8?3&<b(QZUK.6&2D^U8)^02QAFZdWQQXYg7Ke)_e<8#RXL8(+c;Rc+[bg&^
\&7<_d-;24abLWXNU4=EHIM4b,FS47G3G2BWBD8/+2PCC<Y8[dR6RdY]+:<@R0^_
9(U0fK?f+V@f/L:3-8)TPV?eBcX9YR#<a><LM+_RIY<\01bb:N=9+J)?34KT9]/+
:C.B\7##Hbce:f_P:g#(E+-0R9OK?@EPJAbH_1Z8T1<V;fPWd)BF(8Z6::2KP9U0
F-:HB-Q-d/7>>9M\:J9dMAK5+>5:P.(OP:;M<L.&G=NSS>Z.YE5,(P(VQ&@>dBI5
f]YcWa))HVKAaO8cJ;VX9JGK;W2f[YAKbaF)TTdGLTc&\4g[UQ])W@F&Sd+=R/Mg
8SQ?c=UNAZ+<2Cd,8[Y([ESB]:g[4J=<)_8@1,4[#0L#&HO.6P@-P.39X?Y\J]_M
@.CZ;G0f/_LRN=/Q2/ECW+Y\O&&X66^54[DbCHNObU^TC0R2W54fL[,-95d3Z=;]
++RJf7JKCE<6fWgO>)D^AA][c,#>P\2)NC:YU)AHMa+&O_M-.R\)SRO=aC]Zd^4+
E+DQ[5)O836-_GdQT2_b6(g.1Q62bP=A?HVR/E&CO/QP4DUL@1>[6#E7T]:][7@(
Q=H3[XL-L5B4aBeZf?G@?S#4CSUYI5D,@5/7FU\-<(LO[Wf;c5cb3dgXL3+A2EfL
A;QfW+1.:S3NK3J/b?-2H/D.c1,2g=6,bDWPAg&G&#CR3A;6#=7DY#-FK)Sb:g9e
)(EAU]]PAgaMdR[Q2MZAEB:XQ[13+03H^,4cL1RPeTQU.eYLc///H/67:bGNH6Sf
1A&UgP:abfO2-Nc6JaGR2DeO,7161ggNB0KQD_UUB^bbBH1,+UaMNEWF9B(FfG6O
\VVO/,>6f6de5/;bQ<)>K8K0=)-]YV[dN69=]YR9@;2EN/]T<Kae1<;dLE_c>#92
)2-WE=S+Y/TC4&,GDZWRa[)_6V:M[1C0-caLAP-PUF7_E?0MHP?cF]JWY/CDH#+5
ATA;gL7/-HUC+>,I4S>753G>[,3LW-,)-0ZMP^>dSb2^^\Y/;>I]:fN)c5BI\5A<
8OH3G<4E0OK2,#T;3B(E)82Nd^ZX>]Y6]]#M3+\_-b;).Q=&PCc]X+(g79#>#_L0
gV0S?DQd4#TZN<K<#V>1:=-ATeVIB6C5Ia3+^3,VY].:R+0Hb/gUed>YNOW=:B;\
?TFQ?gG/A.)D\,KKKV4UZf9LQd+V4E0e=IJ;\&8WBb0^R3QRSHOEYg/E+\+37)+W
UQgP5ZbH5X;DKD34=B-UCUf5=W^GB<]2PcAM\I<?E3;WQS_8:#]XBg+&XIO<]DJF
TP(0;NA\aFXNZP_CG(=^;C:]d_<1DPJ^>7USN[S<W_+\?,F89:SWcaNg+YC&c+g]
\Qda&;#(de,;0>OM..]^N<cDKIdZ5CNTW#(2WT>,1+DURKeYT@PAN?7eHXc-8XJ1
<=_I^VX[2bTN[FC,552#I2@#;+D4JQ+HOKD,g;UB#,@HScVbZ.>]AY1DV]MW#_7P
T-CC[KcS?]61CNT9T\Z91U]THBRS4#+,FTG_d\9.f@WAM&TI(D]<&Ad3>E(&[XaP
Z;4:5#Q9#a4eA4VPH?+=XAG].P?\U025_8:GU(OLa)\10M[SG#D5-RB6K_A6Q;SM
8#7<KE9S6OH(6?a6VN5FXPQKH540AD5IAX<;bD_;WEK2D63]H7KZT4g]gFNS>?fC
:6^8#<+:6?&4-Z8KUQ>aH8(e,FHUFR_SO)F>=Qd\34^KL.0EIOE3:;KBNTbLDM6L
;)5X+e5AReZ2XU\eW,3J.g[B)AF08MDA/R,[R,M]NXZT)<&e#&TBd3SgaOa:cF,e
TeD_4cFbG6ZYaWI^RIP:@P4aOH5eKAYde.CE=\f_<egd);e6?>W.^@==7,D?0W,+
dI2WcQ=a-):ECbgL)5G#dV#]/4]=I_MPGZaKOYSEB5IT/<Y72DTB0T5OUS(TDI5I
S&a(f<^3&Z;P)=:eE.SZ]cD3gS;:B@:a)P_O63512X(NZ_)RSLM@RG8F/WAN12>B
9A[\[3@gd)O:=BVDH/KG3=b+XFCI:L#;;aOcSS,WfN0-[WT(+468LLYGd[87f]N6
1e2&1VA-e?g14YH9=)b;)Id4-M2WYG+DXQS22Dd.BGCd,BKcC\=4][I,H\PI>gJG
[4_.NBTgJd]#N-Q<RG,O.8g=4K\C14EG>f:&2eNKYS3D3TR9F_KD_MSK+RL^Uc[V
(g(Tc,UUPLa=\8445C:U]MACV)Zbf/(>g,;J78R6Ze+c0U_UY2D[?#?5<9ReI88a
^AB1/H3(0ZL,Sb@PB8/Z[ER#;([>2.YYM(AFLgOS)11-IGN5[b-A)S4a/;J.P_6\
;Gc9gEdUY/]SV]1;X@RG+#f0.-Yeb,bNTZ9O>C=/cNOI)DY(GT^D,d&7T8972/?[
b@9),RSAJ:J(L4UcV3:=D)&FUGL3M4Q@AK^-9G:X8/]#BR-EC_1ge->(XEV+Y#U5
<-g0#)\PN[51D:+d-5A6f?TJ;/2#RBNW,\QabGK_&PP\_E)+0VLcT-RTWJa9>8HC
^)5)Sa8+MbBac)T,/&aG.]\d-e\7/LW)3P1AS.c<Ud)a[V66[d9D)XT7OKFZ6-\/
]A[&GcAO\^GgW0<-5-^be^&@U0L1-b3.(^JM7g_\]Y\8[;(Kb1fHR(>P_2UL9Yfe
LP&9Ab7#BB).F&&VLS=-6AM,5;d=]H^fOTH70Ja-dPUZd3A-,dOHY;9P&_fVZ2RR
Y#KVS2RB&BQY^WIc23YgV?FgfWJbZ)0B2>;T8V[1D84+4:YUWa8[^bRHZ9CZ3YCD
&V>(g)99AKFg4^I[aNROK.0Z:Fed=X,+dSa4O:JV)7:7=P@C))(55bdA#AF2R)aO
bU(&#QA.80<V-OS92O1eAY@[?8?HLS4@T),1S]TVd7K5D,UJ04.18Z[DAFX0SR3B
5W6@T:T[0OfJ9@[0dY4a0?J<d/[V3./[,K-5S\dU(Ia/5,&1BS]./IO+D_:Q44aB
)Q)XC[)7ZPY;:WP-YFQS]/GO;0H=>QZP+U<;7>&H09^BXJK]#D(U)2-ZZI:6M-C4
NY;((Q&g,K<;CHVQEee_a8,7gcRZ5ZZ;^?F(Z5[0)/W26QZX]Fcf9S/-(7PI9)7A
5&;;b?35IA_KEf+9SfUVdCaL@8^O2F:18cK)TNR),gf3P6@g.X^?gVA_7XJW\VIT
R/42LHD602X]c?;LA-ARH,AHHX]0A:\@A6K[-[>+E</;82_(RBI4bL>:-4dNccN5
2516/XD+CV\8UcL,dN=P(AY=BR3.GdB)-9)b(;+/.342P:9caE2eZBK:R,+M:+WZ
-Me17B4aX&+?=FOb@4OV/L#96PU;Q?Kg<S?1MR2M5QQRTRU>,F]bN>X2.SH@C&5]
XXaMZTF;g9GL:&=]e5C1_?)g>#AL<gB3/<g8?\-88d/>133E/IZQDL=G_P5@e^2c
^fC3I@6S7T@M#WWR=W1R395F\UC^IXNAPg^D^-fQ&(PC-^4Q;BZQ<\?P<7>W?-SC
<?a9@:DRO71H38e,+d2YIg6L9_CUg_9I<DHTd4_J@T<97WCN[/d_6.RGU_I^e;DN
(D?2e51Pc3,JfaFcK[@BHX6g_PUVJ7H<1eNR=[BV?UPJ3.K0Y()1#\OG7<5:(8>N
e_^9WFDEDbVBN[U]RMRTdgTI;9MK:>4RYgeT84CZ^bBO@U.=VgTF7.#;)8#1,H]I
FFL#fY:(FFg3BE3I2-\.bbdIR]c4&+,N3KO?GGf]CZa8=H&a(2\62;.B&f?RT19_
\-YV;A=;6CQ2B327;A59;U?+)dE:L+^PRIBTXJbAaUQ^0&@X\[bbV/UL/&-N^dSD
N4X,V6d7(YR@/#V6-J/WA\^E>)Z<S=A&J0]X]+<FdDZDW^f03YM0)/:PDADEg6#A
#R]F3H&WHJPe8P5J#UDU(6CA.JPFBMPYf)7JbP.5^ee9dMI,T@>M.L4c8X(=P>\2
g_(98-H(+Q2AGQU09,:KK_)5,\(<9>.OPTB1Z+bNg^V=O45/ISM1BW<A9Ke]8XAQ
c<G50_7VNd)-3bOfL8U.F+H4C\5)/W7c3ZQ)+F?S:YC1,X(LH<.-P#9Dg&J#UR8F
@AR<6^XdJ1LXUKD29HQ1+L^&CT^F.1Ag=>C/F]((AQN+,8R2+&AMcU0=BcS;=DF2
@NZ?<d\>A\#/[XV2@bQNG-c41BE=^5b;2(&gZ&:gY-aAY(&A^QP7P4D7[GZ9L]Q4
^S@8ZdEGGaXC=4##HB?82HY206aPc]aUI[04)Q?D2AOKD&-d2,<\\B>XX7QF8,R8
N3GS\4&4\Q-HX9N[8=JSPd.4eDY:d=gFb<5e]+,Z]G(>QIDS4^Ig7#:I-<_;&DEK
X6=00ffg<d7U40XY09Y@V3RZ,OHC5I(1QMeCWE9,5NRXeY=^Ub#a->WK/(2DH:/S
#dgYWIDQ?K_&)/XQ6,b<3GSG3RO>FW>bGdKW.R=c0YZ2\8YfKB:cF/)K&aD_&RHH
J/]05D#dS.8)[+1IO6\J;R[8cT94c&Gd8N1MIHEJ;S[SX?g>dEI]>^\RTdRA50H+
-?V#F0feW#^9c/:R5LeR39Xfc:S@&d,Q:@J:KE(ab[Z,MBKfDEfc&YBS:T<0=-EI
PPW16Qf^2baH\:0DeW>b1FG>V-NO(0MK#HH:_2?P[.cATIZ61NG]BCKUVWa64e9P
Be/K9HO]S.dFQ0Q,)V[\=6[R=G,gL69G826Q>fJYR+.RXLJ8[M-aZ.F([)<g&OHU
bC^8OB+NUR9>B9C3:DB8HAcYY]d;71?;L(D_Q>Je,bZZS-9:TND_TX=89@J5?Q6Y
4I.cBRRX1[=.>5cg2ZVYJ+[P.;LeI^N2OX9ZJXYebE&Jd:<ES67,d&1Sf>O2TS_5
bP+a:THT@1\MC7(-ZH9Be1eSdbEBR8EK&[;5>MJ;1+0/U[Zg0;3TRD,F<&J5RRE3
U.N2QTOF5GcP,^-LIBf3cQ&Y.:.g2Je6[1eFcN=5F+-[;Ff/J/7gEB/WJ(K8#)+G
L^8JD:.IM(IV#:XW<[V\JUg<KIWM<V5QY]:;E13+@-MN^NRV@gd1_MCCCL96T[TS
f^ea&)dE>&:87Kg0dL.UWSg[ca/gEDNMHS=7AJ;?#_3cHD#:MT#1:05]f^+&:..5
Q>&gY##60?Xfd:GfONE@9EH_/K.19^CA,\-H2D6HB_@NNT.YA8BID&V[FL9L(0FH
]/a+5X14YR,)MVNDT.6E_VeM@R&5L[b&YaKP7W(G/Kg(YV:3,&9I?6+(U>D?FGeN
OcWEO,R-NPVccTF;3cf3XV/(<MgADD++FPbfI<g3M+ag=:AHDf.1f^B+b\55U?VF
3G)^bNVgTF4VDeKK3Z(I@^&@0=7)C3D#UO6a737<^6S9g1O]CG(K?:CRR?]<C.IN
^@<c4B_f9<N4I;cH()HT0=VLZ+a>J+KW5ZECPK>^4P7-BfWJ25eF95QLXLLfC-)7
2L<.D[?ZfEL72;DG]1L-<6R+Hf4BD<e^W8P13[91^SZ;F@I26?_<4/J0d-.2@8&6
6.IR382A[YdY;?.5W;NEY#P-RNaL263b1XE?,V2SAE-2-REAf]I7aIf-EYX?TT>W
\Zed=VH29M#2T36OBYCM=UM<@6<Y^egO?I1Q6a;[Y9<&P&7LScRBIX6JZ#f)I^18
2]EMCC]87\1DVaSY[)<096W&V2dFUdG.OS]8,,.KCL+TZ/2E;&ON7;-\Da6.A3O^
_+Y3<A5LKY^e^H^OG@:[X=^8gU^+eCF6<^R52)Bc;?@HbXV.=-@NO3J])>_W5.(T
VF+a@4Y3O]N:(aW#?)822+W40XE&4W<D&DN7.NdE:#0H:,(9NGe??IW:P?A35Hb8
87ATC7]2>fab^ZPN1d73,5WBRJ/#0PQMaLXEZ=:HIX1SDYEbRWE,D_/T_13AO3M<
fe>7CJ:QB3e/(1,A(N33).eHVU=5AJ:eSZO>f/+^C0@[.JbJ2.#;Fc?0)(^0)c&8
9IGN54S]^?TbL,7[Z+VV?)X1I:0gdK4<<8N02&?QaW^abO#BVPX7Q<f5/?O1cQRP
d<=E3=DF(=]Pgf2I9O]J]95M;(ZBIS=(N82W8>L)>0[:E5\]ALA#MeHg>E0#EV?f
9:&PYF8P:1RM;LLe0UE_IC:OJCa4LO?.4WZFB[-:L+/#Z2#IP_1-WT#TOTVb&1Jb
d^(,OHEDCB<(:b-]5=g_<b@/42JAc56YX82c,/cW(ZRQLT2EETJ95LVd94SXf6UZ
?D4N)cE(IE<<]7/P7])Q#M+[_-<\dDMc8_OAIM:YPdC-(8,-GAZICZ>OJfg-XD)L
=27Q::+GRae=DNY&9W)5Z<g;LKA#X]C)+Q?BfK2K0C6?RIc3P#TISKb)3e+[>?&;
E,AN4V1RY8E0#I:=#+M]1))Fg-C32NS,7]99I8P1NW@D@NCGOPda&<.E2(_<3+\F
A.(9D3T&,UR\^D\PeYNM2AN0_D8A,:G]._EX-c:JF]:DNDGRe)+.;QVa@S8&]Y,E
@d3e)Ie][?ZXJG+&Q+VSV&GCR@>b(O>dDCf?5D->#f[,_K]aT6_RF;5SP?<7&/-Q
T-(c)fD[c\TJ[_1F:CWVg:7GW/@EJ-C)6-_>.JI#+LL8>[[35DZ,=3FP.fa2KCA:
ZO<aeH.E^E];C_2@R)&Fb1?]GB1QZOVDZFA86DB-V[78,gBR(]gcZ+d3/.QC[Y&L
JTd[U\OdcR4)0J[;4BC7JJfYg4167J3ZS3ZQ]BCg3C8<(-.8a([QGZ&]&FAO.3WP
aYMYNB-4/=F#<VZG&4P?@,XR7EENO;RQM\+6FP2Z#8OJ1DFGBXNT):UN5K)@6F8e
@Ka?Ad)f_7W:]f6J1(0Lg/A+]6<3TS\\)&@(T^I-.f=#;6-fZ5W+.d/FP/RVfMQ+
L;5/B:?H]]\7\)ea>eCH:584Y5SMVY8_#X1P0^cP>C:H&aC^?#S2H\ZDf@cC58NM
8S7O(=2bTaSg@+;@/G7:_W9Zg(]^[D2\aaI0@OL4_0FG[G?F<3_]e6MLe7GG^J-M
Kc0/fW1=EYQ&S#&VKG?\SL(-(#-Bc?JF>)T98EXRT#/BJgJN-V9S\1B.MIXHU35R
QaBYJcSP/^CZ8e/DSgO;O>3:HLQJC9J^Q@WU7N#D[Re-=,XVR//#eDOSFB(C@0Fg
dL0T9dWdZ?TeA;T1/;:Xbd94_ea.#X9WcU(F@,G=8-_Za1VOa5&P^Ld3dV>J.??[
BVbefc[<I8Z2DQ7AZ3N5C&ZY&cP:9H00R,>)_aD75TEgd0J?Z014Z.\+F&F66UB<
?@L<V<FZ=I020$
`endprotected
          
`protected
ZYYeZC45gD)eXed>U:@O[CIg]4E#ZOeaN5.f@[+D6/YBB8Ff-aI#7)CC\\V[EC1;
9.L@g_<9ZM=9a/g8],1\=]&L81^g1]ZSJ;ZL\[:R+NbC:g.#GU_+#]N^3-_O-+[c
DcFCZeA71X<^=RR,JJ)^\5b5.DU0(PP^dRL(_f7(Z<a@<-7^gf1G+9b/(#7-9<LC
?8.gZI-X(fO(Z2.#<+)68Mc5OAaC&GIO;VZeKEO1E>.d5[D:3S76/2,@R6g[0;9E
AESWBP(8>9Ng:g2A9(9:(e[TKf<W#0Kdb(\UNRBS2QFAL1SIZYa@^]@(&PQ4&=dJ
P_AQ<3a;0_#?bO?B/\,LXg[T6$
`endprotected
          
//  vcs_lic_vip_protect
    `protected
b?N_AO9?#\DZ>1d\;M&9YMCYM.e8TLCS>g7A)YRJR,?=1W]R;MCU+(T]+.8^>>]9
6I-RO4JLSPUOBEb=##4M@5S5B,L/e3T_d(I-RVg47=gVVJRX(WI53Z6JQH9YY_2P
K>[MTV_E?0_UZUWIV=M<M2Y,fOW6N?KIf7G1M@g32DS?X,;)4RK6>>[Af^6+YHUa
Be;X<(LKcM72YXLVH^8P#+RAF:J5O[6D:aS6J2ZLH)b:XSA+L:0QWeDJB:<GWb\e
.Ug90RZN1NR:Ef&A?L\[aP3X5TBG(2BED#+6>\-88)QRe-QQR\G;[/&a4N@[Z=]R
>;=S>NEQRbdc:-_24_4,OY.9A4O7WfQC^B<EC0b1W?\X39\VY.EF[fC<PPOSA40@
W#5PAa,TH-2>d/VaS-Hf\AN4&S3_>+AZIf;D[g@c=MC\^GD/c0EZT:OcVcVH^_MM
R?9[a<D/S2P@g+B:OZAVJ0?#R&H4X/U+badLS#\_?^.YOBV6_04Z+_BKE#K;46e8
#WC3KX7OdSVZ9QUJK7E+)SOTV&P1&)3@,Q:+U8#LV4Z&COAQGH9AN0<B:)(&FQ<@
;^c5QBEX=TOXAM=XeL@UHHAC\74=(<SN5]3:GBgB=]M6BL7@WB(K9R)F=]:3dWA<
a-bJfY+9I/V\6SRW^Wc6KVJ(U)I)[F_=OQ&:,@:5,f_P&=ZgEVH-d#K[L9>+3W)1
UV>/RWLG,^SIb/g1..3Td_W7@9=,0Q<Z6JcGO]:GUIT=HV]D=P]a@OeP-94NP&bO
C5F7V4P<&(Q[VZ0T]Z..c<^EbRMcR<EZNHZ[(<X#QW8FAUR^9BS.R)Ie)1V2VGBH
bS^Q&3EG>UG@)0NgG:D6].GM-H4/0Ob#<Df3daZ4b/JDaW2X#ZYJSeC0f)^>D.=J
50e:M;\)8bPFC-D7U+,NcIE/^(0(fbbJTZbQ):_J]V4b.6-O=^U@)U1=WO&:;?D(
1XFO8\Y5+Z(NM(gZ01NO:8Y2N,IK[IMBJR#HcOW7g+aQKOd(C,(HIC7[EUD)PA.F
<.VA(]cZ9(XFV851LXSQ#XN]]1JG?7^[)U1LC?5FdR95WQ6fb7[UU1MgTL?VLL\?
RGUgXd?)LE3)0cB>/Q0==5cM>V#=5\H>eO5BZ&?cd\VPZ1Y/SH(WQTI2PS[S=PBa
:;K8P)A5LeBK#?(FMIe<98DPVNN?OT8^M2;)TKa/PC^f.\EdK7IPABOZF0(;)gL.
cUFc-_-)S7@3aC9eO&(c66@9<SIf09)LZX&</A113JP:]A)JG\><I3Y:/[QMF^;)
^NL^E;QH(dH<RHZaC\4PUeWN,DgQ82K8JE[eJ,SEVY.#&B59g3-I,2T#97&7#N8+
9IaGXBNBTR-HFN(dR?B3^-eHK+T<BCAT_:;WW@0gYb3]4a:Q)N9\NfS[&e=>2Jfc
T4gF2e8;04Tg&JK><N-;N2C^&fdGE?;,:G)BLGKe#LTW-\beCg)_+GQWKGS52f^Y
Q.-+ge[fN910+FHZ,06^0WWSUZe1J;30X[,;JHV@A)L:dBI2Hd/&N_b_^a:M(XUV
991QNYf3[UVQb00gN.B[eOB(XO99F:V9HOfdKN6R=X;6f1B:?V9/&#6R>\3IWMJN
<,)2OC3@Y46G(YF6&0@K4>8\(?TN,^PXdISVKXdK-Hb^Uc?AXeF)W_e1?<fJ>[+3
AKJSNM>H5F_[5]>0@TMg53KSbZN2CYRVD,+HXC08TP&-+Ic=P[bIGKTYW?K7.#;Z
JS\8\f3OJfUMJ_B854Y#MacP;f<:I;gSbcRIHQ<e./KO)&7_5H#7BCF_948;(<.U
1dGcdJC2;I@W6XEeaaML[;FK0B4C0bS>a/@/fYAN19.#+?.Z,SIH?#&&;^.;AMgS
8UKB?cb@8O3>O3b7T#:gZ(84FA)R6E@ZWV_[=.f/K,8)94W?)ZQB8bM:)1(Hc97I
VW)2aBJ,=-5c3IB8==^RT)05FH+LFgYW]<CA@UYa#GMWS4X=AD@+:6LH?B6S;[;J
@Y@Q6Aa2@O+SR2eWF_MO_6GdE2ZbLR@\\]4P;>P8OCbdcO7KMEJW7?DX]5GHb[@?
<B566H5VQ9..6X7]R8Z7:W^H^KRS?Bb[FO]g@gdgC523CTP>\/GRZ-@T/G5R#S3E
T22ATN/-3UC0)DBQ[^Y96)L@16M=#X62S@egBA=?0Z7B8-b_]M_?52FcANF=F2FP
5Yg2LWbBNd=TE4CG.>bNK7Mcb_W.#@R:WK;ZF.V:G]]XW;dF^,S;08ZW1e-6fWV<
b,QE6]M5a+E1TMGH;QD3>71=NSR6#BO?/_L6]V,>H<1EB(R<bCLd=HZ,8YSGQS1O
W=D)B)HWX&/T0eNWG;O4PRVGe=bUD?R(2KbQ9J:RX&.?]=RBc7PNYVReA4,<31>J
Y)6.S4IGLCcdg,-aN>O&9Z5Y4B?b:a52,&L)?Pg3^7\UTdTC-VaN,aI.0Z6ceL[J
F6E3635JB[Q;&EfP4:_.Q6L)=++8&57:KNP-A/=1<=9F(W==)B283aKJ6_g]LKcM
W\EY.X?.@a;8Z-[M?KTKP+?fgM)L:1<>H<MP>_DJ/d,0./KgO>P]3]UW=2V(]#_N
B;V?c7&@H8D2@IR^XSa]db22g4]T@ZA,G-R@f>ZGYg4Xd#I_#2Rce_;e1\H0V=V.
+5_8P<D[8V<A-RLJbC]g84@8=ddO:\HN24M3RX5\82+Mg;aAHP1>./XO),OGD,X>
<KQ2N6G)PAc=3I>PXY;TLLKPbN:S&TX?=I7NG\-H&H22N(=TW-Gd;IF@aKM.97Q&
3SZ+)d9UR:DbD?S15df::>:b312D18fRX3@SGZ\JY^,UT,&a^Fad>1<[AcV9,DV-
>HCfR-\3c1/=@?;0+a=I@L,]9>2E@YV#5Q@IVAHE<9(Q^:E69/Z9;&e3@M@0e)17
T&QCDO,7SAT.RZN[&2EVFI:f:6N_F(:F,=,J4fMP4X<02+M;>7e>,8GNO2]3#H66
(fHgDZ4g]_Pf)GC2>6Jd>]\bf_&V@LX?-)(WCgGWU4G[E52A#[S[M(]Q>U<5Z.?F
9N;Ug019PF03DVX9;2W3IeQ+CE5O@>\D9>;[.\,\>E1>IM=GH+ac].58&P<EN<\7
:H1S2J@B-+8PGd14S9:?H2>Ud&,RZb8/7-M#,eRO]39.bAU##^aE+<Ve[>UM0?=J
U_^_T5R6=/FQ\_\D)AKe6\V<C(?b/T)&2YPNJTV@ZPPY\[NQ1ITJQefYLHIX\gVU
TfE3@8/U,Ma/?W_V6(O\I-C93WXDb7Hb3aB2gLeY4.?TH2c-XJ4>#27(daa0:/3(
_15:A]LSAP(>V[3DFOUK^LK-=W\D^:/,;1919^2@60NMK95CfdH;8aaGNSWZ:]-[
dTXe#dVW4D>;G[baSbVB<cR._[69dfdf5Z:1=Q]HU=..XH>Y9=XT_ZWI[0RUR1/+
CB-><(J#1bb+HT@3b4MO#N\3)-2:K.):X<J_<YD0/446g;G<G6[3fLX5ZUY_Q\4Y
I;AFA,;UJAQ>;4+Ge4[LI.(SQfXX]Je?=:c#P[-a/EM2N9N;_S:X1_T_:MV>6ccI
2?+VKe+X80NQPUX@7MKYPa-#2/B::09<N3^@=TM7R0HdL)^)Q@2OZ>U;9VXK=+C8
d(,Z^U[9:O92TG7V4G-#V,bA=)^\##Y<::3Oc<C00d)5^U25U/DAYV2.C[bUTO^e
I0WVYGROfE]RbaKEW:gEQdH(<dZJ0ZH+T+ba)P&W3_6](gQC9Z@9IG+A5335YHT/
<JO<9.M[ZY:60->J)[K1QRH_R5/>V)1.R8Y5F]Ze(.NId/D2JUAd/4/?X1@)N3,F
]gV]EP0bE&TGE3/_cC^g7PB3R(](>T.USMO.V-1AD+6+N>UR5_eE+[1Ofc\0K\eH
TJ+#+5_ZLITJG<Ug4[,FDGSZI#()e&dFaIZAce[A(_57NZW]MULP6)>+\SL-[e(7
aZ/bXPZgc+;S.2YaUDC&LUXCHY&Q(G;S,65HJ5E,,6>3DGN2.(<3R7J4W+-7?=]Z
J4?ZcY6dAR>;:gNXA[^F6L^:.TaV_?5/NWPRDNWXZJ)S6:/4g;Gd6?<PMQDcdD1U
05OZDO[Q-gOPcXG1-DFYC.)+EEZLLEZ&XJ5?J]_d,<BXK+dd;P87c3<M4fB_B+]A
FFPYY9;c2<XYQ]&]5XNNA>>[&6K1O&d4JZfKWCf1)QN]QBW_gFAS3?79M;CG2^N<
gY?68McDHUN5Pb7ON\Z,_PD6;RZ\EBI?QZa7@32=_XFccGD-^gdG;JMaH;:<HDc<
K<1B;2KQ;dY-4IGS?BRJ,UXBU(MUD_&_g;3bCE_&#6)6^7+F,IKIMMa1bd7VVRO]
,G-W2.)6C#;=7&;<Q;DO:Z)?0JI/E/LKO7Y^C/[Z]:0Wg8Gf)IC?3@=3IW7>PH<.
M,0G+d?eX6GgZ;bCa=I69[CE+QQNb34Z?7d].C5KBYG732W+WPSBVJQ(_KF(Q]K?
28-cE,;.F-3<D67BANLb^K_H?T_HA6+MN[c@82BPH9X8@)6^V5.LG(UeSMHHOd4b
=<-cK\Bg;=+GWJTM;VAB^:5g6,6V@ALPIPJQRTVd;WJAI8VCIeR)a.]8YGPR8A,f
f@(BUdTN-A-X_bWG(ELTaS66TJ>\^L(Q2IO)AB2?-CWS_74,06V+d-f?:P82=a)-
O;IZ/)M)+3BNV69GRAHR>,4>QgTRIJB0@4X[-QB,(dUE_1)-0T0d#@D[?914H@(_
)6S0Y(_2Q]T;c#M?3O>@,&?f_BUgP_,Tb.L^RX-<_IGM-IC?(^XFeB(c]TK-,BMc
ESFaLQfg9I89f2#2&bKOPgKRN(W/C,U:-A\B5]GgPI@Mf(bDRKA.B08LNWfcUD\2
_TPF\V<ROIW\(@Z5WZ3MB#=6fRM)P&E.ABdUHVW1ce\9+KKSY(GHe#YN^,6g9P58
?Sb35(X\;c8JD+7]^I)LF1OFcGXGf>.3c?PN>F/+.@#(S5BPNSD>@MIVA?\SE(E-
]A++_]IgBe,I<2B-Y/M-c#52NMc7f)Y7Y.1D#?=<?WQ,YYZ((6:0c@[SRed<(_F4
DbYW[ce&19V#\](DdHG^#;J&5Y30IG=.@eU[f).cLO<&eE-WH+^Bb;J.dAL5;TXB
-B13AKG9KY&4\]7_2,_7\aNZ_H_XR.9N4^L^agH_2WQ@a19<T#+#g#UUYHR(]YRe
=SO7DX\.MA[R+(H98_[XQ+]3Y2[&0F_]1WO1K-Kc[EJ6KbZM:#\.AN17>@4@Rd8P
52MIZ61BN0AG/-IcSQ?>f]&8c]7<M)28@AWBa9(bHRA^^[RG=;cAA53/f9//EOd8
BJ889e#L.4LW#A=9B2L43VaL0):1<SeP;=NM?@Vb-H^11G&dT#>I.bJ6^3=K(JLV
A[T.N[?d;Hg;B7H4EZK)Zg2)b7/9:A7RD:fPc7[.L7DWgTOU7/JFWd#3bL=E[17I
[ZWbOeC_:]-IF>V9D3^C\:./9J2De9VL.Qf:N9ZWPZ@bJ7;(X@CB<V@.61(2EJK^
_\agBfB)QS,8F[A4^42R/57^G_M&<@fMRMJcc&]ED(YF50885MYg-VJM&XR.g(7C
(CL#b1WV[.2<K6=7>XaJcO]MYa?<81BVgLaVdSE9aQ,S:/&Iea/[4Ug_5[Z5AWIY
@=C8[A)F5TOSf:WdI?10GIF2SEF4LK#dMYc@/J^d:>B5S0_P(09(-A;YM9#T-/gP
J9BUA.?cdbI;7#K6OXVFMTLHgf4SU;.T^QaW1O&RMaN&X0CK,.cB).;=87M96O#Z
#A6TRdS(UW@Y5)Ja(d-JD63O#;B#&>1f[@+M=^e6)CcgVR:L:P0B\##BT8Cf?a)3
<-EMfa,OY<4VdU4=(DKMMK>J4]<.TR?[(=Y?AYg+7Mg2SF;E?2OF75XJ=DUFIefJ
Qb)TOfSa(fSD#;;IgJ_eaac:L);3QKSD3LERb)acFS5TO)^#+H/(FV:U/6&FIUC?
e2>_FeJ3>VQN9)dB)^9ZW<3ZV\f](WFFZTgA54@=708Cd=,^VUONB]Z9<-(MfORE
dXN7CcC@?eS&afNO_,]fI.68KM[V;^5I\EJ\c>440KVaYP<>NQeO6fH2;W=2\XIc
;d?f;=G70VA+>/Q+I53+VJ(H0df2d&7&<\f;PP(:WP;b<G3<CU<OM5DE0A/B_PP]
/_:-D:JVJ&)1@_b&,1:aXS0^_X:#@.e6D.aLS#YB(fCV.]-./#,1K1b?5PI<cO<@
1)A1>O-GU5[C\L?AW==8=[6e/cb]O1EM^C[e0d4.\.#MA/OV9aAOPODJ\-f\2H:R
C=BQ,,\a@L,7[W-b&9AXf;6TgL6A\?[Kd^QS,_;f=b\Rd3E,6e#^b8Z?6YG[LQ9C
V19G_DMJ#d(BCXcgYC;WCA:3Z@\=:)SZbC7EVVNc+P>=3XAOM3&aC=g@WYNHI1f]
AD11Y[<He\+<Xc@-)H2>JH1]NNA+Y;0G6Yb.>,de.6-0_[e8;&20^;9eO])LA)-/
](bA..3J([_H#M4a422+Sa?ZaIDX9JZI(_WJD36,@(-9,#5PB_HH:Rc?YA?d25\Y
:7R&<:UGI3>)aH2LIeJ:+8THdG2gI7dIbXZE]FEeC-PKG+U[H?8:fR2HJ]d(\S33
S2BDK?Gc3AQ\&.KcJUF.7:ae&HYHNL,aaA-UFL@D_?F7]\HeY#FScQ;OT++U2+3?
/-ORJ+KO^.6d4e;P;\Qb.G^YZVHD);PZ7d;O3a-F#/+IgH:\?G&H&+JJD-(KC7[6
,GEF6P[PB8QIbYPT;RaRNS<8fS)-XD8CJSD2aNa\0U,BIa49<E06?@7>NVE3QYea
VJT4>]df27e([W&U1UR/NQW[c)9bSOc=QTfZ^f6=760JfO-D_Z_dSR\>:=H<<Z,W
\e+<:Y84UVB/&9(QOSW<U2R@F#FI2-V0ZFA;A&4?+(Vd(+6O-RNR&F+;67=LUU)g
Zf?3N(;OP<:R7=EJ;Wa3H#ZTNaaU)573aU/=^AM\ZaUK_HN5<FUQgXJP^&(]4A7_
1=D]VSMTKF@Zb#N)5R,SbQK/A[[TcQ..TE.BKaCf5N<aD9gP57a06B;/JL1SNW1T
<(_TR3_[,YY_4gOBLE6GPe:74>Xbd#EZfQ_J9I)JM>>^bS[TEb>g+?L[\<<6ARMM
Q&IdD+3<gP(GB^BMBRPBW4.9S2cJH4U_Z@</EP0#HR44SVYEDaIY2gYd#1S^g4/L
EAf]gQ#GXUHBF[gS]B@&SX[FQU<>U:#DE=(7QG>eQ-8P-B934P/2HZCSYaB&gR<7
2TKdI7eB6\#9<^9>Q-VIZeV)]3SeC1&X[B=SUFO=FZ2]W:JRS4.IQ&58SaBOP[bI
2X3.G3+fP,dU4dQ\UEM:&)\&g.SV&=cGf[Y5&/bA3=XdBXDHBE1J9SF#f87;]_9A
QB\I:6^N<Df43Vd+e[B?)_3EV[OfG9gL?#FSP&=6-YA)DE?[c>deJRg.4AdY:&OZ
<>F-I&+L>G]V]L-)<gZ.4O\H8gc/c88R7HRK,fX(SNBLN@T49[GA24+85a7#Z;N:
19-.@LL8@N8fTU(_M#]2&2V/D.7RgcMa^&gW[I30J-#QBJT:4gT7Y4bH=Q&[.-8a
S#[acX-0/>TEI=&1dH0:]P;eV2ff45]M<(4B_HP-X2/G_H+=KcF\)Q\^-;>5<&CF
D4VM4a0Cd;BKW#,FG0KE2ETSdMGg3]#B,SER,IG?Y>GVA\Q/AV[\A&g.e,AMg^7?
).#Q4C0RV;J.V(R+\EF<IH/X#c]-Q?e\\/:L?,93&SOg.-(X8U7OG+VGWN<MB7.f
d5f:53]:6c#>L)?A9RBb961H2PVE=Z<ScWU\Df\G?:TPEP74>\MN[VReZ.6+Uf3B
Y-F6C-a<eHXP,EBZJTce,>6^TdE(]3O9CWg.G):EN#CQ_T\MV6(I>d1=49[PC:@I
Vd27LG-,3K]9D4.=Q]LBb+V:B^3OJ&G>e>aFO?L,V0[_E:4]KgTQ+@LDK2XPVQ^U
Pde?3?GK=5SA?>LN5IECN&X4eD]EU05<[5T.aC(MAF77,HcUPSUbMW=W,5<#,Idg
ReL>L9P<g..6aX7b)-7IS[TJ@X<Q@A-(fSd^c+-T@;-5MW@+B?cb7dA;YC-3[K4d
>bVC@E[;-dLA]X;f6V9=)O_/2XaO@?>ARO/-\Y0+KUA[D/:JL0NdC]OK\MbH]MY[
=;,@TS,:;e;eTIJ8R7CQQIKHL+B\R>:M,6+:76T?+G16Gb13Mb_4UOTD7De9cN7a
.,IGE5UIHSL<1(Od)(:>a5#1H:^^YOPIO_\]9TcY:J5c0D/;0F#e)cY/67bAS8XX
7Z[QEF2/9[2C>.O6<fGY.BF-,]7A2eZ7c(,=;9Y0:)J9@8CCKG&\^^]X#G>f<2OJ
S3Kd28fK4P,YDUAGB&OK(&<H1@P,,1ERH1f=dHQ@6P80NdI]T1RWSM)I99-8/dP2
3d9L9;gH+Q-8D,cN6d,1@O=JY8Z6KT0g3?O1BdXD+T/J?^/5aI/H@:,2@^\0gd^+
RL1)1\/ZH8f>(,ISD4&ZH6@:a(g0P50[(?1SCbIZfMZG,\Q5==3;WHKEW84ZSSZ,
+^V\\15(dW=V1#G]V4:3d[DUJR]=5V>RK^C<\N8:O6P/e,=:M/a&G3b8Q4VgS,@H
FdRL)c:,H&9RE,L7PK[.635N?EOX&9<./YC12R\:P6b#FfCJf=6?9QHG?C0^=T:#
c9,aOF^P6)TL[2EbGMOO8J9UXP]G:E)0#:QD2E,2[ZeKgA7;_UEE3M]KT5GDJ(aE
[K0Y<L@W,:3?^<8T2TRF]./@PRc^Q2+M<IF,T0N3MV(aZ5I[&aL]Af)BYbBgIUd_
Gd5V9@Og+VKB4/2_YGHCJT1>],f4_+FY9Xec6NM/3<\\SBB.^:O4BFK7S3M6I#\f
L^;GdV\HV=H]fYc/^HG/BKRZ9\dA<)1Z0JLfdQ8be.1^SA0JEEV//R(WVJVJAORN
fbF1eF\SDb5Z6\A[R5_5+3(?9P@;^gO)BXT(^.TQbf_bF)8FAP(gRe(&ROe.N@GY
H,+b^77W<L[7.dY12BNFU7IL],U.e8JKW=,:?<H5d^Y_f2bQ&<d#;?[&.NJeJU4P
JW-,=&)J;g2W=S8^WeJU9b1K28Tg.Y+SB+3V.Cd_cAA^[A.#?VSeKC-],I_+4X57
de7STXD96B3PM0.]a8045/\0>[3G,^M3#gK<#H0CV&GGI<ccO9UQAd4g].^GIXQO
6UObb4d@G5,eDO,2)-U#T_A/cD_XC+C.E@+1B[A>F0:J&OMcdgM8RcF=H4W#WG77
-W5UG?&e&BG^;;VPA66=EdfFK7&=UCZ4Q@M8#U7#\]2/JT0^N]WAT5N:^/622-eN
\((?4(RPL<a;]6b@KLbFM^#S5X=#d+ePN&<M;Z/^()Z]_XDNZ-(O?HAM-X>YF<I6
H#(JXD4QCb+BXTXBX_\J.eL=TYJGcgfX.W3+X0?HKK/)e-=5WAXZA34=d>)gQL&;
4C#TA&1>^O#KOe34A/LK;Z4=S[V.@=9f/3@f(@V#?N[d;VJ4\2.\9A0^Xb+EO-14
G^S8&B2<:dH)4f6H@T7(HTVNM^9TSe7fG(@A.TFV0WU[c1Qad.A:HJEAcd/5+e;\
0)MU,99ceEG]F\IfTJ.]TJWf[4a]C=J=4@3M[HM9Z3:ND:&A8=F;U(fIcW@8>R5K
.6gDeOUI?DV.HYZ?H1e=Jga5e9fKL26Q5F+U[gHdC,#4YO85E]Kb4V,0VcBHF10Y
38XLK_=YIJ32;:U^N\)[(B-LW-/TV)(-bBd^60=JGUQRdF@=Y^ZJ=CLe4?85_V&/
BA<f\710aQ[ECZ_;4EH-M;M)8Hb&Ib^F#RI\:XMNW_4Y:7JNJQ5CbDH(.FG=]#2^
YO[W&c/;B-Se5)Td[?VZbTQNLaUe88U7Z0&YNQNFR/F64\aL^Aed8<^R/SYPR]8e
96SNW?N[Y@E[Z6&BI0QT8J/-(XgC\GSHL-(9cI\P:\UUJ28\DLMO(2a[^CA/QMTL
2?\U+&8MS=PMU^G^b6/2NgO=R:EX0WKKOKC335Z@<[BJK49HaX?BQ/Q[X1].6V0:
=T\+0/@0DR&b(>0;33#)3=4L&;#Z].E,]3SL.fZ-^H/]7.]Q9<H/.=_36/C/>b4U
F#0;W0NGcDK>Pa[F0dg?L+BBWUWfAMcG@2^gJL4-4FaSd-^Q/S)(KfLaW;8?^c6d
a/-PAQN#QOf#=ba<7VIZKW<ELS2+W,gF2D-CWS7#31).Z,/URcOX>D)X=JGfF?Q:
&g)2)J+Q46?<IZCYD4_K)H@NLDLaAU7NOfCJd4b<2);,UC7#S>EgY1AgIID#KTW9
1b)6Y66=<<QdV#[bFE3G89^V@X^^HU3E=f]KGNKVNYU0c=CTBU;].M;.99.M06fM
,1BfAN1ZQ+-^gO=HQGU[beEO9J)7D#[YX8.Ze+0,4[W3[O.MbPc9@1L1J=RVDQ_[
d#;0;<ZA3dd7d4dPB0(](\b3270Ge0J#Jc?af1I]\2FPf<A[EDf1X_VG@Y3)-IM3
D-_GP:5_CAJ^;QRP_I@70V4U76PJWVcT:N>33;R-/G)Vcd+[g),/HXfZA_B=L7H]
^f=12MWET2XaU=_(JK2dBJ5.)77\@b8:^^b9DXaS_?]8gP3QeFc4HHBOO\_gT.^6
ETC?WFeD2WQ)=cCM9N/(BfE7BF9RD<SDU[>JHIVO.QQ9-4])H^-T8;;WW2Va8HPH
,O(HbATCL7)<,W4=a91OCb)SMJU,((SQ,QP?gY3B1#\W:&JZG@6&7ga@a@:U#KNO
8G99\S<)gD4TO[NO+=EeV8d1HSX,\V&WEeC6a1M1cKKcTR488B^R]5JM4&[\,:H5
]N(,Na)g(fDZH#@b[OU.8Ngc::B-05#N1#U<5K,P\W^DD:3TA5E]Mf,?FC,5KV7C
dD&F+<RY+[VYZO?bZT[8B&](>PHW3IC&.WQZcA:]/DALYeO.14d_U^(D<BW2ATOV
(#Ca?7d&MP4]B>B/49:SbAX.@WC6/?aN19MLaI/d-T]M@IC[VC/Sf6^)e2H=ZG2:
V&2KV1dPKaC+KE0PR<E9a\AG]L2>U>0L=_>g/G]f\9NOP#EAMI;A.<8G=);/PLGS
)0f]QP.Z>fZ0XJURQ//BX#,-/a1fMN]UL0^\f(LbB9-E[5YWDIH0GcObG.#cX9?(
/IY+H/e?A-ScOAgEHBgO2VGOUVY#6&b]RM?SYZ4d/3HX?fda_:bgB]=1<T_J&+bV
]O9d2ICU[?G0=6?FW44D[),_>L0)H;3HHJXTIY4Pb?G#>:G#g=(I>S,]G.I0:eaZ
FK-30AS,JLeE@4A14Q6A>D-6Oc7Q(7+2P;/+Za5Q<V82NaG)B?N726,@gP)[@GOC
;6<-OVZ[J=dQE.-AgPPaWU^e[R6cN8XRA8)@5#0fR=G4OOE;U^YO=c.B@?V/a0BH
WBH>O@S_(UX&0=D#K2d[E+8@#/VE@HaQ-\A9HE[AbZXa]]9V.EHd6GJYaHJ=DG.P
K7\U/O^(>1b/NGR0eY9^^gF]@>7J(dd-T&94bD[Je>]9;#;g(cY4^Tg,1)9(^(<T
5=K7I//>G0B\[N8FY15W?c&GCN^;5B0^@;?FP7U41S#=U76@N175FKC-6EOU-Z+G
M1^\I\JaQ]0^S=#bYKI[3WaZA,GF+QM>6ac/L#H;).#)\8GXZY7>77G+GaDGR#^H
?+g+\a5,AgBe_L)cd&W#Z@eFG#>,#S@&U&8CS+\AeX]RG<;&9;<6g=O?+GeBJ(9d
G,:?cd=af+&A3:/La4Z-;#]]#_+=bH:H=S/FX.F5RTRJX79IV?P2M1OcP_Og1.RM
E@_6.ES-)f^UXLR(U=B^M4SAY<\>-+9R\bEVM\=B+6Q,40TN^#?(DX/7C#=F.]a1
I+16;c0PfRY/.cW@AGcdB1(KbgJ@#?:5MX\,Z1bgP/URHT&GM#&e60W0e(@fN0#T
6EZ+\MO@0FZP2T4MU+1^4;D3P;B&L(EH;94P<OcY2-&U4DBf[&CUCJI8>PM^LD2Q
YO8JY>1bN-P/-+?JUJ\PH,e#N_=J.=N8>,e6.D2:ba44O;ZF0V:DGWQZS.W(+0G\
NV@1eLK==(Z>;U76K-6.NFa_4d:ZTbY=&Z,ZDZ8H?)0bJ6H]3SZ.+EZJAUK\LA(D
GK#AW^+84X^V>&:([SZ8)9U5+eSdaUY@Y)5GfNYAN1#OKaeF^)M(&=C,F^TB>T^N
Q)JKad5e0[42OPKQME10,FJBL1RT\8RLYFATf_Z<:P=]#RE7C(4(\9<e>8FTR6/O
^-:/#;KUQ5RE5M/facLb6eT(TL?g=)EWJO9G_PBFc6?aIX_D&XE.),?TQ6V5UMTR
B;SSS.0:B89]XRdBVCSQg8^#@/HX./WEO-HJW-QAU4(D\WYV8:5(M1bf1E=<DcY#
N(0>4<@gB>FP0145cFN+XUfDUXJUfN2^C;aW7TCdRAQ?)ZOBb6QTUFe@=/d:ZT+6
Xc7P:ZT,EbHSXX4M0I^_f\H1f23JKX?OIV^?\+^.ZX90b,S]?>_>^/0?4\DQE]Le
>KecU3eQ[]&<ZN9N-5e,^C@gN]g\f@LT&+FH?X1[#01O<:\POd-<ge3Q(,\g-T43
=9CRVFGeJ6/0[bZ)8bN&aL\DCcJ^edI,V/(G#FTcW_9+MMA,^1KSRH-;TB7<U1G#
#QA[C/X9#HNGa68[O8[C[;50871-1J(;_UNIgDB13X[Xb&;J9T?=Z=LgHYgB6D5<
Vd9cDaXI&[\5R,CQJU+<K.bYKSbb/g8c)RL,MZg_PIc)PP_+\]&.6NGN603?GZ)g
bYB2f1Z<5FSddBfFf60PV&L25_9gf+3-4K5GSVd+2);]ada:<Tg(C1M-&:eN8;gb
O<d.;3/A7[SP.:#dMT3:ffe5dGSDG?XYS/MOeC]E>.SJK;c9@F=7JOgP.Y@SPVad
UE-Z9:_O1+E[P=8#fU[+:EEES6(;BQb/9cg11RO(D+3W&]bS,PGbd<gZgZBa1]YL
QR=df::2OcBF^YS,@3S//A4FXDe&T=VUEWBM?1Bf>-<X59c)e@#N8[;2eUQ+4<0>
U]OA(V&7c6,8O2MGCRKM_c/VEBK/@6<\<D8HQK^1<I?_90:f:,.B\7:F80ZI^,J/
4bP:YPYBH2C8)bQ\V=bI<cP:=R&;R[EFG=)H68J;2C>D].(e?D)+OP=IUIaG9/X+
[M+C;F58>I4.\T\E@7KY331YUL<6J(>]EDa)/f>DI7U.5fLc_4;A,+_>&9g_WQ:,
P.)3]R#MJJ\2M)C\S6&0F#)@&84243K?#&CB0W#)(:,N&V=_21gg<]@a+c<C9--e
AJZ1[_4K&fe.76<M9g?]-+@3G1RWO8?WRNT_<@SDE^.]K2fXLFW1+OHP?<<HO0#g
[X>\b3EDY/O>NAQ:RGY\95?7dJ5[5^NNdRW&/b>LL1?R_)QYYHBTC+,GB?T?g]@3
,:E;&cXgZVXfa=0TUEE3D:+f76<MDOFJJ,>NG4@GXY?H3GVbPHT,TL\bZ?>KXJ#5
a6MU53[P#6[NU8BOP0,dZ8FOf<VATW^Q\2+\ZPb(YW[9^D+)X?<P4XR6LEL_;X,4
^5GVEV:.6Q5FI?KE322VBDAgR[);72SC0cYR#UHLdg<\HN1Z[FIYXY)1+ID,^#5\
@(>2MU9@Wfd0G3FPg?;E0DXf4K>>YQ/5KeK1.cAP4fF@MK:CP/#G6_GUSF.TfPUd
BNI[SFdYQ9=\IE@,CR(E(a=.N1_@BWR]0M>WNG7\ACVKGW1O8^OgS=?\E2N[Cdce
CO<AUZc64C@X\6919=DTRf5LdXL>P7]0,=V29TFf7UAYf(/WB+SfS]9WP0PNA/cd
#IO59QY[V8\F;F#OY@:@BV(Y&HQ-\P/^6(57##)=WE:84[30,5bf;&+g2(K&d4NH
<<[O@WJ)O6H_U:AbX11CAHL8K\G/_69F^?&CHQRgD_EAGD)D(@06Ff:20&8_f,Uc
E/^)_^=WV7D[].LcWV72H,3U3H/KD)a7OR;XJI247]48bD1]OUC4TZ&ZeS@A;5;9
=#Ad1)/WAP<QX9Z1e2T4^SQTQLO]HD^^#;1OZbeI_?f+d(/;ZdcBRCK/,8;O]>Cg
a\Q8YGM5^4E07Xb3EZNP_?cSC\C<gY^=Yg-C&(D>Q#T8O4Ze:G.]e&bN<6e+EQQ(
H_3GTMV,HFTRdVHQA(>@DcWb(K1fT7:OZ#g-g38K_.+V3g6J1ddKERHfV)J58c94
UN,c.E7ZU,aVg+VbX;5AMH+]W:#4dT46d-_Pe5?Y=JV>F6KW9QYSL5X,)f4TdE9#
>QB2GRA2AVN<a5JP9CdT.CJ1dHJ:)fg;IgHA:=PX4?TLN>_K/EL<;HKL(9UZ4bWY
^;[K9[F?TBb@]K8NW.)]S7B/e&5HG;>RBD.:3-6[?eH0G^U.5-@AMJJLAN+:dJc5
LZQOCLHRS?cYJSG-DgOUf415<feQ5:^1W7&Ec^_L&76/U^FO>_g991K5GM.CAW(U
<Tg5+GRFQ6cBZG4G>=6.57&cG;,#1(Gd1I_7HaP(&e(DM_[C?7K,2]V8\1Q+UQ(b
2:\5>7P=65G<NQD^Kb<bY8=d?UG)2+4TV)S6WC;f^fIU5L=](ZLTB7@Z?MUf[Z4&
,FB(&1@NXULZ#3578g1[,<e/P=U?f1c6EBWFF2FD&c(]K;b:E\JV6O3\b:/YbGGb
[L7WF/c-N=.5[Mf]8Ed\4?S@c8E35>[J.:0(8)JFe^<ecMFHD\e18^:KNfPT/We0
>D/a\=ZA=7W?X;ZUa[0ReET1Me98=M>NcJLdcJe;(7fPN.gC7^C\4C#\:.^QVBA9
T@,g0\\ZSXZ1&Q:dOCge7+KZ>E9bI;dEfU=>Qf^Lb13MX?dZ?NVa8@(RJ<;MVU-2
06=1>:3B)OcBgZ56/<SeaEN](#a5N<d8SH0_2N\e.GG)RZ3L[]XACI#FEgFd53OZ
g=>9&Vg?^HSW4TO\N?D^T9M0bG2\#:L+@N39MbdccQ?QffQB#4N,SbIOGN.^,DfV
W)eENgZ#Z]b5=gNG-[DHA5VMXKefd2;>SQ#a/D=+J#\Lg9OCGE:8)W4MK6R1+.d4
_9H<8&8Z[/K\OT;NLNQ+Y#5/3CB&gSVVJK+FL]^PUdPH^..H&0U_8K>8?<,TP^L>
aPfIb)3;F#@_76c/HH2MVDfY@8e.JH;/)cAdN#XW8OUCF8O25/#WKZ=RM?D&(8>=
)4aW@;#U5/OIEIb;9HQ8HJ1g,PGCRCZOBKEgFCcOG^5++^-eY>@:+V\=(J1(D&G;
:5>#(^Lc.NKATN(1BHb(J+\/0d,G6a[9W0AbWW<64gb[[3,#=VC:HJd+cU10B?@S
2K6Tc0,[>2\#c(@T7?]d;5FIJIF:EYe]OdE[PJYH]+&H0:.9ZUbge?aaU2I@Q/0=
]@12-0=#b4:6UeP.9[X9W2]M7ZfKaKZXfXA9K2DN6?>1=,[<c45UR(bB-\;1a;f=
)UcYF?/:c#L4f=)V6ePR<RWIGXB=.AL_VBEf)V6,g=dM0aN38O_)TK3A=<)+D=b+
JXbQ:C#B:M.J1^faaIYIW,1VUP?2^/V3,fZa5XUI^;JT(?7QJ[Y,f90g_.=FU)G&
f)Wg5^Ke(33GaSC<S4Q6Vd6)]\.Y0<-X]Fg6C/#O>Q,PUJ@e(0>0d8)->_4SMG6V
5DKV8c997N+&#_?0H><);gH+d09)R,6V02._=UB>JJ-LC;2eB(1SJO:+b5JaESO=
UC#W&PZO353DIB6)?96NS\\0(N-_eX3]7bPZRg2(,&AYZPedW6VDL3f2ScJ4=eC3
A]6IY[<YX>,U#8YMI83\eWH8><J+0fEPL0f=J2GB@LN[-MZZZ^^e0\?/VMFNgK51
WE7c)?3gBH6I:0f,&IU)5,WDEOeTN^8UbA/c0Y+cF-AFK&6KFaRR<@2JR=^A3Egc
Xd]MXBVR<f-5#Of9FRUD9Q^/.Jf8@\(\Z3U6)QJA.-\Pa_9R;LQY:1GYB.N=AcGB
QODPQ:.+[Z&d?<cSYfN-We0+Xa6=(7e1)(:#ZK^#.VOD\>-XT..0I7EI?)+\KV-,
A[B[L=&F-(=877b=8Oa3UA@.c70#MJ(^4BDN\XL?[B8&I(Z9-+Eg_C(\fdK]gQ<4
X3)3(.WJZK+0,0I]T.<#b4<B3WPP>B<N8-bQbg=RQOQ).;.QYE7eFB9V#OL5Ng_b
adJN?/--B6<a,.(TARCZS4HZ)?4UB,/HM8FDBY8bfF#T2STe+.1=UPRUXT#Q(M98
4((F/-]H@A8<.=FQ.<LVd-+M7V[U+J[TT_0.?@;=5>1\;6C0H5=9=c0BYMFR\Y=g
X/_-D0WdL^HXS^fQW-2cK0W/2Z67W:I17MGcI&5/GU@78-4UccK?e(O@JMMQLIdH
2)D7a9(AQJ@NdE_@//D7.R+8>.F5UY/Q4?SJX;>IA/4]eL+QTO@YFDf]#F1PXV7N
+dHI3XN.Rf[>cC#OV0Z=IC<9aXg<?.NEC<0RQ1H2ZNWL.T3G2Y>T.R59PEcEeRND
I:-TH0-@84?8-J1GRA.-BQK>IO4\5dG-HcTETJYf\4Bcg6eY8:?0).\A>]QI/[U)
f.8M>1=.Y\8C4M/3FaLQ/7-W5V/&3.33\(U,a_\?J@K21-1[g,S^D-GaBGO44<^<
W=5T^;PK)dU64=d+;E7DC8RS-Q5-CHbf0LW[)0KTgbRLV/(EgUT3&IT=WWG;SS7L
Z/-_F.S)8/Y4e=Q#O>S6TL/#-g<34e(MQ#b\AB]]4[@NNJa9YXd.ObUXW,1@;7cB
4Z3-WW[&3:(UHFXQ/TN5U^6aO0MbGdL&&HL^&A;PK#LSFH<15\S\:#4PSPeW@4HB
KefHZ:-RX5\fIMF_#=16\;#4E2>beeeVG]<0JEf9d.[GXNC8V1)8WXL=BR=;A5(:
gCD(0Y;2_9CI^/g7J#\)QHYWOCA2eX[O6=;VW1ULR4+UGGH01-I20DQd\NKY_8Bg
)8g.DXQH?TX6.M>8X7FG8?f2C)B>LFf]\,R/H:&dIAc.aJK/4W<4_WXLaM=c5\ME
RM0R@_aG@C9^DR,XdH\T;ZgA^A;f-3ZbAZ7H\JM52G.dd0aGY2U/I2)=)#+QCH.(
-RUaI?1.NCNc6&@NCOQaceb0#E.bFQ#;>&#EHHU8-A#c8-SS-GOG/cfg)590Oa,B
L\I54>\8UFf-QP)QT.,C;4SKMZ6MS->;bd5WDCUKOG:8aRSRVN;]=/aGG/7cZT.+
dQCT6[QF2S8e&ZQM926VO4dQ7G/0R_VZdI##_K&:0&g#&/YYK_KRO9B7DV+F1=FQ
-M6]88JV-bL)cCRK^CGZH9R;1+7Q1a\b]^&V?dX;C2P<Q<eQa<^e)BfXJ=d91\_D
a5716a2W:?->_7+2\f8KYC)QVZ,O6&H2\\^g:\CV=&D,J+Zb)H5U#C50W#DIMTS-
bIe/JOXScW_CeRe([,gdG8C@IdgO)#C177XI<WJ7F1OBZ[DXHEGX_+/MbYEH.2H2
Kf;<MGYQ14,/V=]2KOdQ\GT=5_M(4DO&:;6;W-A9ZVO?-Yee0O1PdLSQR5/<-[eJ
.&Kc26B=D=81ICTfD0&OXHI??;#^aF[U64>&M#cR:DU-H_fG\0@YN==WPe1\]V=d
T)+ONEM/&RYQbUPfNg_eC_W>4gO,4.W/[2aW]=g0OZ)DW?(RK&TC-;=M0JEZ<fS:
L_PPa03XA/RWHA,6-He.Vc]5146<_M^YFAH?<4A[USIc[aKF?V0BN&^J[OKVXgb6
]KHa?/0A<0N2<:(aX<EKB(L__]D91b8)Y?M/TO@:]=/V96L.L>,F+Z?<Q>U@DfM3
eOLL/4:&UBe-6)YQSO_+G=>a&^Ea<0[XQ@MV6?,CN=\E#;3R,G)Gba#Z.QPF5U^\
dC\7:G4X,PRgV:Qc5,[G2aT-3)B4F((Y8C.O4)26E9;)@-a?6-?9?S^DN;:UAY;@
C+X:WJaD-?9;;Hg_b-[(VOJ5)@gXg/L>VYP;0WKc_0=E[e#C,@fW;4fc6SQ:+c&:
.Y+D_OY@J((VW>eWU[<[5J&DHcc.S#V[]F&Q_@<=BYFSLS,c0agGD1BK2L8T_B@=
2CRAXQ2XGc/L(SE.Ga?KC\://T)B+(1YK6D]RORZCPH8XC,?1Ka+3K-EN>JB?AO8
ZAIX-MBWW;cP=8/Cg\(^[UI8/A,E3bPF;D.2.K0da-YXZb3QKE:YVd=370gFM4f\
3&F_P.a^B37+;PK/607Lc3+TLB^:SHb4J4f+V.[JE@\^63:(TX8(Y8J/I^+A6>,(
Kg]1@Kg6Wc8V)bHYS@<A\@>38_VHKY_OD(XQ/,VW7aPB]^BN1#P@NM7)&Z7@e6=K
5:N&fU]C32.,SZ4J\8^4P(#0M0=4OUP/?2[FZ;2:73+7OW?50Hf9U75Sb#1EKB4>
447\JZH5b:Z:?PT;D6c<8_ZbEgH)c><g-W^;3]O8S80g-/;cH>PTeHQaFNWb/:5-
/[;T?@g+^Z?3SH\0]4d(/+I[\G.4A+B@9IIGe#6)<fQEWf)A)#;d,,^TX3Ha-#7B
M0.X\QCL9/Q#2[EXa8XA_VA8g17KWg/N&LB-b]H54NF2I[._dN#_)N+?_JE0b_]+
Qdf5I/<4A>69CZ7LN)TBGe8P2MP>Q8E9fXc#BN7CK7DB&96g19OM//+1aF,]?4g[
6dD@a<2;OFF8dRdBKH)+MLfKH0WKeK3Q&QDGK62Wf#[Seb#_EW#HL_]HYXQ:I3#-
G9I1MMNH\-b]M]7G2Z^QU968WM2-@^WGH8LE6H]VGCZf>2=,XD([/g6@T_Zb:C9e
CO09HLZ+5F:H2]6^6&dES;@e6??+B2(2AM):2S?A^N(g=Sa(f6&2P^.Ec8U>bfWG
g(&fc3TB.-cWbNQI\JK/1-LA?b3a[+F+G.V>4Z.A\[J5Z@[R:ScMEd)V-(XS,b0\
&=L/\D3_[Q.UTeLJAWQPE3JZe7;+&>,Z_SPAeV@@710U,[.#A:DVdMPA?cdY)dF/
D6a11Ca#H<HWD.W^b#dS[0O:2Yb]8IQVRIFaU8O_OB@)I]JCfP_)\AIJcVU+I5@:
bWF>UCD<.\M?[B8U/b4F(J)3<_(FZP2a8FGP,2XFdB&5DL0,F2AT;]+)HRX,B]&M
:a=\[CaFG5bcS1MFVd)^-Y6^=/_C5W#8?AC9(bKa6J-^=:,W[YT]Q4<G[YFK>,MU
SN+d?=DfE[D>VQID_(/d8B-ZE7L[VL_PFPKH;]?I+QRC=c;fFA)#JD4eTA2E?NGW
;8<A3+bY>[=DcaVNeA]U<WT6N7DfH<Jb01WHTAEb<>gQOH:)H7KUO-F14<+6BW[;
gRQP5NV+H+/+bG9A)6DFI0E)IEZKcB+8/UQ4C=UP6J#K5A:;31>NTfT9YJSH6S?N
0^?-D^GU6JX]3f#.b8[QPGIZ?^Qe5V(a_Ja<eSAMS0<:/g+Z>-0(KS=Md/[L^FW/
Ke=[K[D?]^F:@\86H9SZHZL9P#Z.Y10FHRXaJ2Z+e<.JaPM\A0Fcd,9OJA9G4TU8
5XW,d=<3VFH=6WIHf0:I9@D59_.d8APUEX+Ze3^IcI:1289+CgG[9IbEOZS1\E_2
):&E+,4UUHeIPd?(F+;^8LSYW.RC=^Fb5M>C,7fIV:YQ[8GI0,f[,NGS=H4/PeZ)
;a=gTL)1^E>:O@J:G_/e(d)ZFN-;)O:40YaPBOeH.48</8747/FG.Yd[+#.3G32N
EBWPLO@G??DN)HMG+F[L5/X#GN^JXRK(H?6QA?Icg6HSW1>\UZD;47-;B[gc5C(@
ge&62#&dMFA79aGU8D&LR6PeF-K^QNcGTD]#DR?VL/Ye;YV@1ET2faV@d#bKa)MU
6)YbcY@AQaK#;C]:OW#Q^Y_f7&#-HL/+[2^2?-@cUGf01J9LQ:(1ASLYgeU7/0+<
X<F<-FgLKD2UY8]#BWcgb^_[D?>OJ0(=afMeD-b/8@H^72=C?eaDA+YRHDaHOf^8
2V>)<4SSN^gHUM\bYUIc29N_b)0-NBSJH(H(P/dUG-=J;MOJg,5>G.Q>KXSP=OF\
&^J0V)ad2eT]6bW5VdL9U0H#ZbdK.)EAWR,ELbe(BP?SfAZ.ga)E_M1CZR@+\(3X
-CgC;18&^PNY?00a9&7Fb:^=(N_,I]b,AJI;=^8(e:ORHTeR>QBBF3XIa1@b4LS@
HfR(A8P+8+?F2E]L72P-BHN<H&SJ,_HKP<<5]\^[a0TEH2-\9W\=cKML^d:(P[:@
EMPIA>SY5UW9e3&JbO^Y\I&QHW<81W32E0J,9e@.F+HLG:J(ADRD9c^(E<4(<JSO
g4PZe-W4GEI,O-G@]a4)ZU@e8QPb_\<A0C_a5R(QHV>.B4DS))PQQJ,,==OD/e(]
)XS:ID9YeZHfQG0K0BM/0QV^UQHBM27P[(deKTC[PNNG_+BSN8HSafCV>&:#S<aa
&;XF\a_5LUI(<U/9<]_af0.N=cZ;Q/f2A@^K+\<&Q/dYe^DMdN=N;c[S2/DL-;1.
KSL3ARA(Be\YF<P-BY)(O<)#DYJT34J)SdE?7B2.(/L11SK\;)8gU&B,QB(P_&GW
39c_4+D]XZ#JVU\U@_&>26NcAJ0&#X49bGX53#2d7(@<B1U#V_QWCGT1S;:Q54GL
=:F6V4#5Vc3WBDQdE++<GE9JbF(]2[#J-;b1Ra>JBX2&a(&^)(?HN+eXWP.5SA#4
>M;3&CN&2d#6.Q=L)SO,e?ATSOgTfFagN-?1]PP:YFA<:LC;>3BFc@2E9_a6dF-#
YPJRf@3LBZ2&FF1Z]IbAc@+IMLB+Q3N,0[bHLB9++<0)-P1@J_E_.G41A6JG3<TC
Y<:/7EDLB1:0K/TB>g#S=eBL0a0\SA_8]=B1A&YeD2gUCg2\aD8eA&=Na<6\AS(0
#59bEFNF(H.a)a5QUdRW^,^OAY?0Ud4c/)GITBUBUL3;+PAGUKe7]7f@G^^[E9Y-
bP234;WJbY8[[b1eK<c,@84Mg>=W32YO=,Y2_1(8a3S@PG0c@)W[NDX8+9.Y4g3(
dT&@FC2O=X30CG62Fe27HX(b,9G6<cEb6K&e5]IK6D6e?:F47FVPK:_,eIC>\^Z4
\8\g&JfPUZD;7X)F=M;,KTFW^ZeWJ_:,(_?GbJ3KY7Yd55:)A?0?:.7b=95=L6I\
Y)K7MK]FX(:@Y7-F<gEI#HP^D0-&3TKf#;bdVGaL+B];L(_3ccGEDWdKf43NJ=gJ
<T^R1OS=Wg,:H[H1SZCDXY+4B.(<&YSeb&dH>5;KcF7,)IQ1fDXa@AFWG&]UM80a
R\<R@@+(8OIH@4>W7O+g8e_+-<<X@]MGfc-U:+1C&.Q]C73@F?\BMed<LR#HV\JM
8.)_YgXf05\f24BD4DG/0JDd4P?HRXF\36]8&NLY4P#g&DYcKFAGHd:;@;=H&f?Y
;)A):;ga//RA=OKfHDV9\R;;Z[f./O05<?C[T8)dgT:NUCPQ?BS]_b)R2-NRb3[X
)3]a4G9W/_7#@+#)ZKd]/44,1OIb./DS/[C&?131+E<.DR4#73>c9Abd?4;U?MUM
Ib9+T1X-(>Vf-4-8T1]/U/_?&5Y(](31=cgW@KIcR-U,.YNS,S&6G2_gBS7&C/.1
,I,EZFF\8H6\X,(2ZLZ6LZ@BaR8((EUJFDV5McD)7L-\HIAcJa-c8b3B1TdMH3<b
ZcMaE>+AR@76;^)aKF:EH>_-6_#7,Ve:IA<VKQ&U,&Sg9=eN9BXS7O7QIYa1@2c8
N8XBeJYbFL1#6>FL28f=g^NP/[^72)Mb4[<H>cE@2\1<Z)L@fF;IA+J#68G\=7[R
IUC-9Z/V(f/A;R#]D+S8Mc1Jb4._9_-]Q1E3WBETR38d[?XQ/1,\40D2Q<B::#Z0
Q=AA9de[\<9d[4<AUNUaZ]6(25]:V/GPG+]_V,/IQ_/H5-E76EP_8#R;&N?+@gW]
+ge^ERXM#@JgD\L6]Gg6f8/=T,R64Z[5[ZNUQ0b,G;L#e^06bCT_C)]J^/=00edI
@&2Z<W/VR@4\NHSD4:;K(c:cK?;<@#.gB8]dS(Y#Fa(EJ8UG2P?=#2?JF)EJ5E])
?N^TITA745>7I9GV_Q.Na1S.c#,:?T3-E0g-^Y@g/.A];#0@D76;(>:]_R5]]70&
X@@CB>9V>;:N]ELI=YG,]CH3f&GO&]cOe\>TRKFG:1\a7Xc>Mc=ab[AGPZC\N&g0
Y3d/]5//KM;_1QbR_3JB8F?/0,MLEC1_8e4.Y_E9KKZObdKYH98BSb,M5gZ5A=c&
VaKPCR_G^DH)gK(#66[[d^DKbUbQH;f+dQ0V?/.NWPb748O(PbaL\R47LcGM2-NB
66=0a.S.RD1E9UA.cDBfZ.YO(dBJXQHY+QfW#C,B)EVR^g52M#Q0QH4;6@@54WgQ
RS7C:<bd;2ABEJ-6Zg.P_(@GYJ23<DgcJZ6S81=&33JM7g(@Q7FCPKV-JLeVG0)4
b6Y^7]FS#&KV,WR98#_EJ6<9QYHXU8]TE43T,I9P1J6OM8==N-/FUUc9C^8J9W.S
_9H@S&I\T;Fa/^ADc;2cU6<33)+@TZ6N/4aD@SC/=58f6cAPDUTRU&J]S/EbJJP)
G:I#=bXGTZ0Q3-9H,05e0_c8,R0PR0+V>S#M8R<L+^DITWHLC30S4LZYU?]T?IN\
fZYga+\#\5M2:\E17-^FMP(YLJ<&?^>e7&5U2,KKR.>XIIL#Z8))I8>P)NT]C,H_
__SF+#6.09Bbc8b^3cgEPRgaR\JGA77WJ:GK,Z.@M>>H45W@ZAc4e(aUXbHc&PYE
2)Q4@;591UK>C?-7<AK:4_>LD:S[0FUNFUB,D4(e&^H:_2BfPL^1Z1NDZgNKF:@X
YL60D5QSKYfDTV]2dRM37+YBFM([>>TB1(6LB41)e>fD-E:JI6JS+Je)IMUI:KGB
_?YGc(R;,+aAZ;\?3G5@eR&_\=G824(I?M<_K7LEaD.-+gI_Q+QZSY#O/Oa.cZe=
A17BBOBNJaNX>[c8A]=dZ5LPSYL]d9JSW->+X-fV=]GGg#1WT&J&D#Z#_NTSca[:
6^Z,-EFO1XZH,W)NY459AMg_gOO]@W+:UQ9L^YO]AMRQLCU7J7C;>c&E_eI_A#Z@
^e3dE;.Pa@@#EXg&,2G^4?[0:;QY?Qb,]8IP3+06Z^,<3TS7/3Q&6LBCNEc-6RZ-
a)aXQGQ?TK(2?PGT.XacCY)C:BR5W0]-4GGVXg-AfU4T=>3XQ3A&C-D4/71G4^@A
/:(S^?#@f,cE=0V0FB-P,P6O?L2_fXV66/P\c:MEXZS(U2=ER+W-LT+gI<;AKO4G
QU^cW4W_.,AScbf5Fg0:OUH7<)ad5CDaYWb&Y]X.Rc&WX;\]&LR;Be++XKe/JLIM
c4PJB;A_@D,:^VK?F[eD+U6UVF1(.7T=>JKTEMKYAA,ML@ZPTW6BJM9=LOW6J0gC
Td0^-U[a1=:/3YT)U?b8+Ec4]QJ8;FFI:G[caC2I[TeRM90\AV-;X5GH+.9(S8^a
B6dTV<b5V/WcVB?&OLa&H?\Q([,cSG2Nbg_P/eF]dQc=,cD[/(?M+=e<FJffFdbT
c:@W;NH/f\#X,D4@^/5d1ZQ/Y@)7&]5>O0J5b^9[_CbK/,bO7)/F2/H<7YZgPM.?
>g^H3S?XCdK,N\X^(\S.R?>^6BV--;MK67WJY-gSR+AaO37(GP:&ffcPeF_MV0]K
_bP.c@I2gI@Rg&B=MdfNd.W0E4CTMEXX&f9:]7S&#L[8OgUV?[EZMRHK=/_D9KdY
;a:CFbB]7C^c3/CCd@1:[Ng0\>R/Qaf_2P_eWT5R.VLKC(.6ccgNM=:Vb#AcV_Ba
c#YMR[[8#e:4I;+&&Ka[XPJ(9@aKV-JY39aeF_9U/3C5^KBb\51G=b^(GTR+H728
HM@PDBNU3<J6#>J^?ZFMB3^B)6>,4G1:O\Wf\QXYQ2#5@#P+ZO,e5Y1Y45XQ5d5P
:/F^dK7FcYO,JfKbPWV0H?.=4WH<1VAgc93:\]b=GdHS1&<)NeTU79AC@K28OH/J
-\A(<e&Re9D-;AF,@N=d0O^44WQ39-AFA?Xee@]]XSfCJFOFfSU7G[OJ<J,&=77#
=&T#4aS\4Ef;e[&SIRMD2cc&XU41\?&YeXO2]:@HNJ2MO+MF=(@I7+8K:E_c<CWC
4>-0QdA9L)G-d=GCU70F2OVgCS8^J88TO^:O:0)<]#](;bXT58fB3f/&G6\;-#Da
#M5LK[J93.fBT_D4S^,f6>b:U[ZA0/dTWd=)2VW+^/DG^#aKQ&+P+Lag8-T2O.0U
SSb:7Z?UJO;KQ9FJ9A8DW@;Hgb,c>K6D,Fg/@AHN/SbYeK&BDJU4QLH7WUBcA(M<
&?(>5d3&#=<GY26dO,cCO0a1(@TB@a.Y.FMO)X-20SE899G+8T_GM).BTEI#A&,A
D078fKS8J;_/#XG,]-WdHQ_YGNV(H+W>M/B+X^3F8gM5_W?SHV)##,4GA,[[@+.6
4^VKX[aGS#&H-g]=27UPYYP-#/N+)acY.U\F&-88:XRLDeBTP_^@-Na(eJEMOTK,
;1.d2eY:OfPB3A9@C<4@FX\F6J7+\Z30IH.g&2\:JF@:.7(:7:,7g5S#.g,=T#;6
fXXY#?RI0N#2Q3c6+gS]M@&Yg+&<[:f1@[.0W;IQ\Z@^Zc/>+>\3B6WX.K#___4-
/KRJ7]XYS4[,B+S)<;E5_F\YIMY;H=LS[<[/WKgERKYL+GTN596]^@K5b6],^\gQ
FRJdJ<MM+UO<Y-PH]DGY2Kf+&6CLNIU7Cc^>==VPg.9d5J:&Y:XV<FBX.55O/,>N
#+U@;2O>76XNYfc&Mf;bPG:;G>[b+[C:XG=T7Mca09T<QC:\XE1R_GKP)VW?J:NA
QIF1)U5UZKeR3K?7,c:??Y4I#MGDA)c@AH(HVU6Z22DUGE4AHUT#a1#C]da@^8Pd
_HWY#fF<&ce3X1,C<7HdM?+_)Q)b4AS4NJSe/]CAR4Z[=)V#+?G,bVSIa/#M?4c(
9A?(,29BI;L<<,-8UW9B+_@OJ_25NKaDcG\_AgU;_HN[JMB,eNI5)UcY83<B^:N4
CgYYJ8&a5BdQ>]8J&RX75Z<+P]Tf/dN(>6AJ\01J@M\[AK8\=QA2MMG5[/AR,E>_
UM<T_DWI27HH)1<bX#</75#eV-^S#6U2_Re\Q_T8d:=ME@VZ-;/;G?VU_;Y]fQP[
KC976D5\WMfA+9VPdWW[Z8V>Y),(,RKgc9GWO(/;P;4WUPA2\X[DL,D:c/G(WC6I
;_g943=UHX6<eEPPa[LQDT[,S;Y:AD1JL.^;QEK0JTUQSYKQ^8aW&=A16TIIg9K-
c&F6>f@WN:9[4db+1UO3:KUKa0Y\#NAWfeg#Z,V>)1\7&F-J1HZab&2__R_T(U1/
EAW1XRX4ZeQ@_1gWK>,gRY14-8V7NG(Ua_;RQY=];7WF?XQJJ(77N+g=SKePI-3)
7R(A_d,+Le<a8KBgg[X19,A.[&C;FGPN#b;8AF&GbQ\dR_QMW-@&AD8H/CU6CdWP
46e2d-cLE1\^d9fd,JWI:6FTRM+0SL=<SK6cP/BDdcb-+:aQU6:G8>T[8?Y0^_X4
;@=.U:]5I>a<#+1D5UJY3R9c(8cTI4,OYJg0MAYNg8NQBQK>#NPSA-IYK)Q+9>O_
2<B^EBeG(@HNKO-I^ECW?@8E<E/QW6G(PYXE?)b6[^_H:+QF0K81cB@Oc))A@\2:
=PH_VOVPFTY/;P.<0KIaIF\Bb.b#[-_Q(DXJfMM>R+YU4Vc#&@79gG7cT:/Q>Y^?
A+A9&,<Q&.fIE<Y[CPcD];B0BeWb1/X)PZ6TE_:c9C(-R8#EH7(8#3L)FZVVCS^5
M3)<??,^GWagIcC1g:4[(K1WQR7#a[S^:gdF_O;+R2Y>ZULC4;Q4Xa_+PUP.@0K&
LWT;IH/AS\O;fEZ\BNOP?K>TW:7SQb0TM[RJ/ee)T2DCY<5fUVUaJ9L+VAd+4>WX
Y\NV;g.+/b60e&U<Z32=;:cZJ5=X)J]gY?J\>W(\HZ^N\-T:_4/dLW0&B4eQ)+LD
5<@C7D.+fDaXW6X[WgZXD<_?Bg[9OW427NBQdQES.F=deDH1P#JI-=>F(\EKQXC:
M)8VVHL3+KK>A0b8=8(Z2Z#>W056;[EL)bDRH+(0KB,caB7E)+[SAH5;eXC1+.H4
]@DXJ^GX3e]D4[6P4JFRC#\WF8#KF:2#60I4S;LF<e<IT@)SPLF9FG\X5Ve)>d#7
KQS+]<d?YCC4TB90Y:f--4E89>(d<;0b[H8\A/EX5/:#Z)B&+.2K)4XWRFD@98Ec
Hg.]\M;4RL=5cZ5UROK1>Y8(cS?bNJ-Y5M:]&dIFWO;fF+47OH@S)W5Y,#^;MK)I
0BVfd^>O>\X9#-D6,c):^--_JD#.TA.J4J>R(AJ3&6CORa\f(c3d2O(RL[WD)&(@
65@-^6AN<-9]ce^KV9N0U>GFW>O6>ROM;0&@6R4(#+Va_fNc4V#C;WQ4cbXg6HE3
,2&G;0Yg>0131ZX3#Ze7E]\9LD1CW4(Rc#^1JcdP>?OXdIUNP-KJ/,W#^3e=c2N9
5-]J7G/A(=E+_M]c\YS]TURV1I?eB[FJ;1:GL.8;O&)>?/L4YL^YN?Q0Hb2.>G8&
a>C>H]fFYA)5_30_cGI]\W2T.(0cTc7W#a/2&L_0<Z67A?0O0BRT(\/6L@PJbVW)
V:Y+M(Na_ENIB5NMgMRIN(.eLAgU\RB/GF8+NUHV&QVBe_FVUN-H(Y9B,)8g5-AF
10/B3<=W<SV2&IHD4LPLM>G&4E.MT;20+1=B0_M\1FFG7);]g]C@/KY)Md;QQ<(.
YP@(N0EA7D_V5>.UB:??#_gTNH^,/ED1PUXG7/?)O:KS^HIc=)MT,fY2OdVGQYF5
6AAY]>/T-Fc/8QbP.f[99EPPBU-:CXZCeG77+)<CIF4e;VXMM,VD.8+P_B#^aBY#
)+#++<PYWM@M_;WN:g.9W:B(<d3GS54I<S,4]C@f,ZC@f[OPcZ[ZHA;YQS]#E(D3
N3-EcA&=R2g8]W8cAZgceB#,@+)UNbFa,5d0P-ZM?E>/d#e;ECE56O-=#ZS&01MX
;T@04B8PUW.4D2(<5C=ETJQH@7MJc91@;+H]?#<:EbKgWgL1gB\4IFX24>KY,D@+
U?8L8>df3ZR-X;Eb[JHgAFUX<S&E7#C:,3L30Y[T.S[#_(dA>TTDcd^EA&:GL/0d
/bZY5@Y?YMX[>]e?MH-bDU?O=BJ?ZCJQ7F80&_E)J^X774H8bE5T::^Ne;OO023g
E.W/#<D\1//PR:7,^\G8IBZa-H5Y&O0LJ.OC;Y9^=fAX#6(8?<=\<BQBCM#7KRB[
3cLWDee)3<6E:>[)URdTa5efT_3Lg5E^];[fHRS(Ne0d[1W#Ef<?F>/fTSe;dKF3
V1Q#DQF[NE;,_L7\&7+;4bVc@1@SNERF4<?SOVI+g<G83OZ[>^ef82fS_9(#@E-B
[^0403OaY(C<@B:)6G[LbN=(=XBATU#M@cXY)c:.2LgZ4f#IO+g^CdaeCe>bMPH7
5MK7^VeM\[BYK7g0aL0/N=:.0bY\SBY@L,_VP1?ICd#EG5/UOKR&@1eY:CW&79G(
;3:<58VXg/N1.;<<6D<4[V5MCbTS<aP7+EXe6<,0J-RYGfKHg4Hf:,g,SbgQWHA\
3]L1W.B(7PH5^e3Y<WS;COJ)M8HG-640UPc[)^IH_D?DWR3JfTf:JNY=0f2Z)H5F
OeS8PAc0\\>.BG.CCU,G9H_@=U;H>g;6?[R#5:.S,)<-dX9IR)&.M]Ub=I3,DD_7
=cY11A]<.RZZ/^M_I)Z<LH4LTaJ&Y7#MF=NUS;KPc#(dI?6\N0W,:LPQCf;]A&5b
VGX@TfP+>&.J-O;ES,6FbT1]-DM-&YYb&OUVE]D/TXg[F-CMP_bc=-(56Vd=:AUX
7Z3g.U<7/ENN>IDSJ=OT^FSGK;d[V73U^&L]/.-^-CC#SJG6?K]OLQI@8(b9>2:E
=X5/FB#I&L5ZKe-PNV?aY(30/W#.ENSH/)XK000HJETcF/_@1Tf5+)26B(SFJ#SO
RRR(f4C,bV47159\ULL^K,.PfEG71^V.@gNN(F54-KdDbEJa-?4NW?aSc\F-T-Z#
\_b-]IO)PdVB=aSQT]@(N^XF0FUVX;0N@Xb@I.AZeON9@,AVJ;B_]=\ce1(LDA,2
6I:C<BBF>&fEZBLW8g>BREJPI[0=5gXdY74N/MOed5JHR:;1N2NW;[GC8T^R9ce)
H_:3SR)[3H[;>&EGe.TKf2@[V[MDZ?HY4^<_L]&4c7PP:X4dX1cS+JW]JD5BFJ7J
1P&9&MAH>[aQ;(UdZH9UV(XW]Z[/H@#JI+?<MVMCTb?U-T8YEb1\VO0@WCa2/<?=
f2Y(9;.E.(B+5]?](;SQK>dIF(IQV4eZcff4caM>I+QIGQd;)RFTc95<,c>,M;:A
RBX5bYg7BY]C?:Fc.=_15#S+60-I]]XHR(10G6_5S=\FXFHAT@L__U]Ba.d4)+#<
;1I7OUGad.Yd=9OVB+WPF5Sd4WSIa94R)DB/ObfH6XGU@WPAWO#&X>E7&21R+8)O
([B&.VL64,e5\5@9e@OOG58f(=YO(HC]27CBCUY>)e&Cf,I:g\PDL-:^>HWPDHW8
,W,d/1PIbXG-I=BV.b<L6\b)BY19V7<&F;+>=V=5&C7)\->[cKZ\ZJ?Z.BQ.C;\Q
Z<gdH(c8_XU&I5BQ/S7Q]G(/>RLD69e(=9gH?EVeTHLT&:?H92K5-B&=7X&TEUEe
V(eXN(?#(DE?T^N[=7Dd04MSJGHYcXI_E,Q65b.^.SQSY,:CT@RTdMgg@XSW6IH[
5)A^5SJ\@Ie;BWJBO_LD6+JCLQR#(d@[MaVV5/c5[.S\+Y;CY3dA]_TDWO^6af,6
&;H?U8K_B^@90PX\a?/T0&W1)2Y=Z<(A^(N&]E[c\Ffca?F+c./79F/495.@GJ?#
W0_;>]7K[bN=-Jc1;<E2K>S#J(/KVa0IQ]Cg/J=[K>-.3)VPT[#2X\;9C8NPA3Y[
_M;1.5Q9aDHF@Y[fTQIe(346dXUMdcJK4</K^Y/e^fEEA.+(:/]Y3EZ2e+-[6e-I
&;:8UV,?N36L0d].),[^]0BCVSgJ.bH>YCdN4dJ^44W3GK:Q[HG5PfI^S<FJ=Zc^
LTM/I#EQ]^#,QVa2bNL9#&>gM\Q+TLSRQE3c4GR.D/e>Se3.A++O[AH)7N1e<346
CF89?Ld].[X:.9/;,S)\XF>WB]?DG^9JR^4/@S5YXIPMF3GR)B6[-(&6gPUL#6P+
_F6T-D&2WX4XGO@<YaY3V)1W?]/^G4NgbIH46Y0JW912[7\SN.S0OaF)HHZ-aRQD
EL)b-O6H/,@G:M=J3<^CVa.TD3cPa[7]:fDdU0MaZ.4;-/?.N-U.86;^U9H[O1Z/
CF15^_HI4\]c@Ug]J,f:6VQ)4YfDCG[^^5]0&VaD7D\I=Z.1RG9H)XH[a6-Q/[LI
(cSJ>SV2Cc/B#_TD@Nd<-ZSC\+0B[Z,0&b,3?[WWF@LJcF5.L54]+H;Ue0/-,]FJ
A1Z2-;JXW13+eC=:^<>GP(ZTReHK+<2<]3bM9T@EA@(-G#VA>_gQ.75NPY4Z4gFd
f39ffXKU)bE(8E&S&eJ5aB<\T[Q8.PYRa^ae?@EE9\g<,D@^I]RcLaO1\=B17X[S
-;1/?Q8P<4S\J_52)Yd9V<<WI,&L>bKcS:J9&2[@JUB-d3/fBAF>6CZZ5D^5-)9e
Y,1Z#c:RRTe(;.52H0Q[^^5,04f)__OI(?ZbK,4@IdQ+Z)e#H.0Q:^7<CAMF>QLS
De,I1cD1,:-U:BF2R-?+_D@W&e0S=J?VafU2If/J60D20gZWF+UR8+(A>5DG.]GJ
^ABd^d[X\C#(3/eQHXX0V_(2D3#bW^0b>E=SQUIb+f[])O.;3dN]e4B]0YcLDd^0
9FEENgHWZT^Q0RF]^YAT\R(+_\=E3.54a(SA=O6D(5X;.4V\1KNbU3P55gdWLY^+
<U@e<d\V(B2>HgKDT/UdIT_U.[2(IQQE(<X_CAD7LYJW+9.F^G9SN;J\fF[=_0c,
9.7Q:/5X2g8[8^MW&U5[TJ1+9XL?-#36MZN::eRWb@HdISN2JPQKNC@(-MI5S>[-
;/f[KPCACUD:?LX<M:?-QD<(V^>_gd7##_PPafaa@Lb[+9:+f>EabQA.22L&4R+d
bPVCWOS\=L[&Wd5HW&a-/?XG3PQ3GQ.<>PUQb>U+a4d/c:@eQ,AU-=P6F)8U4bPV
?Tb@fTReCMeUZf(//.A:fNR:I31-aG]\SLT(7.f;])WXeDK_8(@L/+Q)CTV(eM[,
+@NN&2-O.#>Y;@Y<J7+?Va5RSOb:EVU58>W9\.H.[6MVT=+NCA.-R.=L\/;3\@8:
LCF8(b<3aRZ<Wg::-Ba=FJ^_=/(6(G.3X1?X86^g8BNePVW+_8e2]gKHIYTS@dd<
b[VP@#_V_RFO5\,dNW>[(-I6I=E9aFT\Df1_EMFBY.BDT#.X])9DHXB,4K0@/[,Q
bgaH+(Q#,8=K\@3V6M@?aX<>F>RDL+X@2(V)7C4P[(/bb:^=d0SALg-AU\LaY?/1
bY<VL/)(OH9)K#8G,/D)76W+&<F^&=O5UXVG:fFfd\4KL@E\[7b-)LYeF5C&/0GG
.^88,_^HXHCV6CNd:55)_3[CT9Z3=H8g2Q\EC^5gA2-3GBSG3f1F98NEW4eS2>]T
GEFEW4]VgfJVU9IBLa1]N)P]J=fLaZg1?2F)#2X,BH)Ed=ETZFVKS[]=A:^/Fba0
7,GZVTbG=(GMYf7-@f6)20ZReRaTYgHd6;(#fKH^J[P-@RQMB#Q?GK9Xa?fIHKS,
MZ<UH7PY]G\SJ^+@^K7+OQ(?]^G@2;/O^,ZF5H=5I.KLS+O]S>;3fLYH^,[ITe7g
R(\F&VYcaZ^J8fgM0&)BEA_TAKc2V^=D>3O)YXK6E.O0P7N&E]deY4gKBX4+eQF4
bA_QdSeLFbL-1\+F3cGK<.50;11WCE_+Dc3)1&@@IB=Q<PV4=6efdP[JeX#QaK:-
S<b;>c8AYZ_5-:?-<0/H;L<FLLP7,geT:d-5XX1.R[cNJ^Y,@Pf+]WE\T[N.-KeT
5E&?P0;K)^2FfS?AN:HGP=,NB^1)YTW?:.)bgB;GfKX158f?5L9.OTfb)MS,IaJ/
3&TCJ@TVf;<P\GdE95>XBMP,CM^:RK)]3NG(#gV3TOgZOLT_WV=gL@+[<ELYK4D#
+>NDV[^bJIU)R)F+-(SUaGFe>1a(c&B+[+[O)0_@60=^V2)?>2B4P[;Q4=?C[Mae
:BN4@RCAS[e2TE=TN)O(b3JE8eQ;XY](]RL@EUVI>D+[(6IT-Y=dWbO-Ca<XB@/4
.R:]BZ8\4,[8/<W->F/>JY[Z2<WPDeCIGU#-R&;-U@>c[\NZPN#0B=__:ZVBd)+F
7T/T&>MSaXKO_fPKNLJTZRQ=L#5>#Bda7F(<B1Pfd6//N]c3a&RLce<IV;c&O_U]
4&b).@2V,=1L]dG?#Ic99V<\1LL?5JI_R649./BaZIE)XW,NX_ReF[:O)2Y9D,g2
H;T41+_AX6_E^.(#COV)3b2+>g.<,A[@22a]^SV0(^+g&Jc@T36eRFZaFgM0)X55
[b_8X?H_gFFZcP7MF.[+]fE81O\AA>+d#a;H;LL:^L,/2TO>61F2.TS^Y?\Ub6S1
1T7DE/0<L+d0Ye3P,QKZ1&@#,.>+&J7dH,V9;UY2GX7SOg\>LEWQbCEC54eg6A.H
\dZe-JL,?7VaZWZ9T]3FZJS=e1U,I(Bbfe_2TTgHY_GDP7NF?P0R>cZTBI]O6Lc<
ZF(L;E/Eg@_-)8aX/1W^I27cAIRJ8(^E,3d+,[3SaI6LP;=9M?KbYB.cNXeTU.6d
#PF@X;PLRMA]RWVSPV)F>RJ?Fg:R]L)dCH\:GT)g&+;9f(WaMedVOK06MWVYU]Y&
b,4]_N9ASH/Wf(8BKXJKVHZ28BZ>aA&0c?]K><_KM@N[fN]f_Z-J45[N1XXH_<WR
EKXXffX6;<P=Q;7,BLIa@3+XcCW/R+18A8a-5N;f7EAC.-NHDP\S(&WJ3Rd)KVD0
>.29.NdAVOG_-fK.L9GW=Z\9W?GcN9I,_8MTQ40=;YNI0#,1O>3YJf,<BAF,\VHe
2A?2>KH/,.bE99a,SM.W0)+_bF/H\]D7.JYJC4,Y@;SST-#IR/&>F+>IKeH.@/aN
X)=E3QWV?=CK-cEF>6?>8-;:S\D;>fe2<5O9&31GT+4@/:7?F_48]B+=HR:T)EY)
W^-X>0T6.Y^W=V2.5_Y.N.?5.Nd^(dA&d)62I(^L59gTVRVFHEg/T7H5J0V5>.Ia
R)LI(XU>6(2\?eE\1PM-Db4_/KKM\N^S66&C<Z<7;^WZM#IfC@_S[0(Tg1OMHV44
3T4GCM[Z8cAKA]REg2-^E;eI-UU@F6K,QNOdWOJZ8KcXRB/3f[.;Q)Z&(<6e5C2C
K+V09XY[P9,6ba(L>IF8:VXA)b=??\be-F0&MMZ)[=MDG^R3_6;Ye6RODUV7BN(L
DBTC515N8Pbc/a_LE=MEP_8^/TW-=0]GW=3TTe17cAMKB6(W?c,:93/Q_Y#.cR_7
X:KP#-\(B0T4ZEMO&HX[9I(EdcVOK)(WT[Y@OY[2OUV+GDOT:C=:/]PVKY3/\LRK
A0(9;Ybb\(=\1:,G9HKTL37[0Sa55cFNdRYOZ+=YXA(TH#2a(=>]OURdZ_PE/T.f
-).9UVW#IUgCc^/5L>\SM#W,Z+H0?I#M0RI&[eN2Ue&U]05ACO,<3K:>P3fF2XF:
BLIc2-d<)^CF_A@4XP5GIO.:>#HZI,6ET_bAd[?&PPfBB[^UgJ)DPH^^R2#a,U.]
FYQL.aGDR>dLZTOLc3BOe7P_-1M?RIeSIDHK?9JD=SGJQ+4JMe;+Mb.gYU1)VLZK
G]Z#.QGAX3VC(@Fd^#ZHCV3a@UUFaB6]bK@:_B#T\U-;@(@3ZQ6eTcL#c#6fC(((
E+D[.dR+(UEDdaP,K(R9Y;UaVL6(5W5RC7Rd-0:P:X<HYA)Uc[XWMIH<HPKY_1+K
9P:SQOaY2/]X/7N?INGUeGF\.ST1+Q?^WPTV5Zf1TY[I>Ye7P>#fbZKJW[PAP-5;
R[DHTP)SB+O](6dJ\M;K5:Y/P=A_3\fOf;\fT^>[O9,e0/GB2A+]#SFOZR=Y?dK5
WBSf:^5g<[F5aa#MeXMPD.AAGCPdV\+TX:C-aY,LML7(DEMO\#P[;D3>-+1K7F<,
E9\d+QVBO/(W]NA9Gb[34P_ga;B@ZO0G)P-S11OcK1JRY65D:Y.662KXT4E@CVMU
_CaI<EE3O0[O.4RF=@/44TY&:LLg(9KHMZ;QNT(C)X37bc3#ZXD9#1;+P[75_gNS
)eQNPNg#SIQ7O43Ff3AVcIHaP)Lb@,0@^A^[=L]\XK[ReT:VJ)PI;PaZ?2HUE?5B
SKHM_3NYDWO0^I/<@1DEGQ/cb<f_+YXGP59G3@N<e4&14;T_Q7#K8GRd8ZV[2&E;
>JKc\e;+\b.=.b3;@9Xc(H_17.OL&a+;&SdS1c@P&D0H3Oa<@]3)A:0c2:e=dY@/
TN,aSdQ[:-X)gGN:4G8J:Q^7<.NU_NeN\8O(]@KY@4PMT-42G_9b:;ZOQ,JHdN/]
1^SQ=EH:M+N=3eW^_01V_QL7BW-9bBVWGT\,GGR0-cV^P#_JYST>Ye/Sea]7MD.1
ac;,8GK9fMDZ\FcYa<9\<=fKe;#V:,P(0ZbfR6?D6=d1Zf2Kc3+P)9#Y\\(3./O<
FT@,4X;T5Cg:a^WagRCUD(?J+DWPWJ/+W<D(-P0d+-JMLKZOI]L+^cVH9^#<8:PA
YBF?58@D,W7>37bU0C^T()ECZaZ+-M(KEAO5PP/YR/K\CE0XB(JRc5H_C0=GP4@\
9P,^V7;0d\+:;N^0e3+)0(<cC.7U.MK<IFSNcNe]GMC\OHZL.\X7(T&PcYE@f\2Z
B(;2QFD]-8,MRM3:(Mb]bCE@S0DPbMGX<5KAdaT[c+\cN96,_c0cc.N@6(Q:JWIF
8^PJI[RTfEY+=\KEX+Ja+]-GdH_.9WW5)=GJ+QFXO(g>L8EN(O/F&R8d5d4_17&)
3#YA]K;<F,V5Wg54O;a(W]H:gA>H<eH4L3=U[EfU?a,O#1.;(;_NVKO-E5YYR.U(
SLN5@ce]VeB?ddXTB/e2C/JC<f#da0E]/2F7^.dWN70JE\\J0ec@6>aGW8+Y@P6K
B,H8e@[a<_fOI4G=U06IFfRd.7K<-/bH&d==5(C&7:0KXY7YY:4;J642]BTe_0#W
A>7Z]ZZG?V?KSTM6[X#DU-OH1QMcG\X9L@Y.6:+,@26\-G3TLQZ]cf57a265M6WB
WU)JbRV_.C7gf.BGR@47g>.3eSXUb:I)[8;<YdAUF&Ja^@d/e4YPb#c12O5Z?Y=^
aF7Aace1;+NVHDR#.:4]D\0NZ/H-<B(V+0Fb=9==?-51ZGZ&;WdXTZ10?U4_WJV:
;X_;Sg4</OIR=YDP0Cc2LXL#Lg)K]MK7S.5X#?(7Ve6WYS7].e.<RJHAG/e:M>5)
#.+_&e-8P=ZF+FR8GYWU\K/&Z1N+LR\.C+VFILOC](I6-@3[2X15gU+c(T&2->7X
5BJ19.RN?>/::82ARMQ>d(<Ea_/1@Hc;&8;gA<e1UYLQ.)\^[RENQRCdb-(7_ceH
1<5U-0BM#Z??EaKe&=PQVNZ&&/<XEf<fVVT6T=-9GGV&?M3WgbQ11O>;?0-GQe7Z
0NdZ#:bICHSGIM2_E>fd/GWMI[#aUJ[37IRV40:?9V<d64=??daCQ[#dc\M_(13V
g9N;O8gJ^FH+;S[e[^6g.Cd8CbORXB.UQD8U/R<J5g#9UNf]KVANYHN5Le3HKJf+
cV+[E.ED8[VFG)L4/RV#4)6#Gg_c/QSQ1RVJI^R5_C9K?6>A>V:8-UT,_N&TX4C?
GM)QQ-(bGBE>@XDPU?+(U+&6^FUUWIZ>D22/CHDb707<5Of#R/e[PQ1?8XL&;][.
\KL/@M)6fbUFRDH8HeQVQRIf+eeZMD74B.;;M7B+#Y1^SJ<@gTQcD@4fEfLT?[@^
PA9.(I=YJ@W[@/I1^0G.ZDL:>]S(+OMZ52]Ua(J>W^S:bC04K7=0B6=,Tfb0aOQ^
,9)Za=Y^<I9fU)>@5aQZTSD-IeOV.8fU:I_8ZaRPM>;G)7G&gdfELDd06DK^0&LD
O_W0M1)ARZXdgY6V5,dX=MFQ[b?D#?aL#\_bA.4:NAQ[b&-?]#;]eXT.FQd]0>C3
8:KMf#__&^K[=T0(-+_CG-WJgg]1Y&J<37+/_0+MDc:QaXANCD,Ef1Z;B)#W1OI_
U0XTC+7;T-;1;dFd6BeTab^eDTX.e:#c<1.S(VV[M/TAL0+,a\6e&ZU^?dK^G0TL
PJY.(=5A0X8]W838Y)66bP]bA.f5Jd[4Q=BV1E1F<EZ3>\b:2+1f63d](.<S@-eR
X]9-[82++3^MA;,VZHc5GH?;=Cc-FFcWAMQ@R2E)X;8HZ8+)W\[Kg8Iaf0@\]1C/
dF9N7W_a)?XCeNT-f0U)O1#]MK+FURAaVOg^WL.JbAYa44(,LXB]P8=c7Jf4M.bF
dKL3:/1]H<O2T^EJT&_eJUg)XR2U@)g\.Z)WX@g7Q+eYRA6N,NHQH&GU]AYWCU<;
C:6c74VeO9/-3M6)]Ha.NbT2+1Q4JgC[.;BK8@?LO?9,CH;L/fV4X8-]JZ^K2A[N
B0=[P5?;T10J8Uf0B?ea.;VgN2^bG:E\W&GY[M_,Ma9d8a^Q.:7MI_W6/L[G5f]O
5VUJ(cX8,@W-B=9MEPDX8U;fN?cg17MJAG2W7M<OROTdf??J@d4Xa.]<@8;<-5#;
32AX3P_&94fL\dK_(16L<BL:23X\2+&dU<Lb<.D+/BN5@aa&-_g-#2JDeDI@;c@D
d/8WHB0c77&9:VMbOR;,=L=.7-AD-90#H:PFI7OFPbWSeJUAfXa<JINU8]?Wa>[:
+JCO/,2,TH4O5fS#3QC9_.+)2=P/?V.SXGRNXWf+.0U&Kf2^E0?S[#JMJE@G1MB1
(36PL7b)YA(/=HOF(fgW6cB,aQ:3d.I_\a4M87,O6)Q-K[IbcbaA86=<?Ta_4,10
]9F=>L.2.W#IK1[UY+9BG@T3S_dD,SFEO]VJ-g0/eJT_?23f714^6dUWDe()I6U:
&TI0Y@EQWRc]a/c?F]@Lf<X3LK[L<&3<[IJ(IGAG9\/O.GY[5b9V,YXY_d^EUH_&
:4/Q?12H07@C86#Yc(<;d(6=[dP6W51::PR]9R+:F;GVNJcWD+L(6)@[J0GM,>;]
(\,LYD#)9V2GS,c61K#F#ba0Ic50?H;@(:AA@9MNVSWP-S\?&+c6Icb9@U^X9^9f
ccg;G@><N=KdOTdf?[b]EDd-^-FI(aFX)Z_Y&@545cSEW<AaK:XZBA?8JE;(gU<f
6c89C<K7/_2eO=(eW/82&3.QPD/Pd2L3IH.02H6_/caE/7R9T+V[B4aC]f/.PC:\
@7M<<J2EcZ>+L=+aNKS=g@ORY(XQ<9dfNW>GBP05WS>LaTJLd>cMG+I-J=(B#T@#
1D)26PNVLff3K.AbUUN^;E]7OaDOVMSQEVg.PdG/7EYK[K38O/QZ.+U>S<@0N5^C
9)>U>cVR(,(-MW/#/@4FG-NLP)6RC_b779QCXZ0\YXMcZbWFPb1]dcW[5eUX\a@X
3Q]fEN[9@Y>a[?W&NGO&3TO\G:7=BQH/2^Bd(S\.I7-d[K\(+YXXKZ@LDTQ8363T
M032b+@+\KC#T0C?bS21IRdZ^JQ7/B]IR]9bZK-Z?\,OAJ_XVN/0aV)T.+&-cHVa
:I5ISO;\__(6M0R15EC.0__<]g5Q-R3/X>7f?R/<3OLJ<)(DE+H@)LW9+:>G88[R
J&BB71:VR^N,/Vc=B?L&BJ\#5=^2:4.JXD=Fd=]@]6L&_KG4Je#:BbIEI;C10QI]
O7SDb]2K]dWQ(F2JU3bHVF>X9V4ZHZANJR)@SP2HWY4:LDIMOdO0L0cK4b]>;9f^
[)FGE=/6IG4cHG)(DB+=U2DV7O#TfS,4)U0=Mg:5bJZ]C4:BRWKO74=PPNcG@+YH
5.9Xa5/HgEB@GbL:W<3S/.W,Vd6OOgL-K:OB]PUdRcgLWcGSUXe<(G+D9V@e)DUU
DJRQ6?M#X-f-5=A?__4dP#(@>b?)Y-8cV53=,QceU(^b?ZfYFS3,6fK9KH_LX22R
-J1Xg#H1)fg&JF\\<<-5]IZUC(EbBS_^,10O_D^[=,2XeAPLe<:KI(P\T^MXC?Rc
CK0IL08>RL=)L&.NY^2?ISReOARYJ-C.>Z8d]eB1ZSf#FFY3dOaG^)9Q&@2+PGQP
]7COeIWKO^3T-=I/AgeGU>AgOD@Ta?D)Y#-e6>;BN@g]I8MQ9>6AJK)SO58[G#7(
7UR3#9S.W7Qf^_8=d:1E-I:8>5TO+_5NH:2NL[M&#2XXT@>[+#[G&CWXY1d9+9D;
Z.H4D8I:N5.LJE;_2)QT<2b,e)ZSe5<ZAA8G?V9AJK8B55.[ROZ_HHfD=FV?K#e3
;-68R?5d>8/g[VNe<bTWB&&QC^PcDcaN4F](X#]&I^<M:FdA05XF/E&PAVS)[L0f
ZM-HSL8E0?]LU;PFTSM?(IYM70d95F1c3UX@K(4QRQFZXUN_NN]W?B^)fGZf_EXd
ae1VYHMHNOT9-SG7Tg(8PK3J7[&@6W[,C2T@:8)@67e>cb[3X[Q.UQZ2REcA1QQ;
.Yb/^ZGELX,]L+1DfQL(f9JBYE+b2VeO,Ced([DWH^Bb6T.dMcGQN]QBXN-(F\6V
W)c,.b7B(FH^/M]5#5e6a30[=K-Q)DTgU0Oa1=SANOCWWSVIM;@3JJF@0OTc4]J8
#4=(NdY-M=a8Bd<fO,\2=PY&(/H.eecEXK3,cP2B#?TC3UMYBe[/410+^@egT3d1
AZ.)Y+K_c3+TW?GD7f#I^(9D8QFDH(9XDN[INB]Zb(.@KDZT8b3<=HOADI8FECSL
HJFTETB>-XFaM<a^X=5PC:d2,aM)^NR.&T\[T630[K.L&7LZNd-;]FUF<Ff09L(+
?+U.#(JVVeK\YD\<R.gA[]eY^Me=81<F-4a5<,DETbU32N^bfS?-UaZ,T(UZZaRU
DK#L&J(eFZ9+1gaT[36KM\,NDb5GE3_93P4a6QS=.=>1U.]8P3/+A6I6B6G6;ScD
-/3I[@fe23(S&5QXXfDe^DFaZec3d1M18T8f4OgJQOJDaKLNb#0LAHXPT<KFSb9,
XLcb&Z:=H6L+eD/Jg+c-5,(UC6c[8#KVc7(HL_,;1OF\f)I<@gd>@A3PO?gB\@T)
+8/58?Q/gQ>#eC-Q5//([AQDP6..D8NYNJ2N9F6bX>W]HTZa2A;V&(/eFgK&aODK
+efY@cX-\UeU4FZ1[T#/@P5K4;XM[47&\=YRW(GK^ZHcDTJ[&dcL-d\VEUSP6<H@
BH]V]f9KZSEQ6a\PYaNFM+YIfZg+aMV2QPY2X5QNKL@8M_5<H9/aFCF#Q4RCV?#O
3TO86N],E-9?5bWD9A9W#6ab425_>9#:8JFCHIQ&8+8YY45D]ASeXH@+Z8B4AH;J
OWD.YHZ,(c&YfYfPK\.bLXf^P<8P)e#E+.B^1K+<a/eZ/g4]([>B[BE1?@7EYF_]
Q7F2AD_;b+b6+)?dEKP,U+NG>XS3VS>J?e=cVZc^_GIf//H29[MEd53Pe19B2dKJ
=#3;U7L]0:S,:J1QVD;OR1:^&MMd3#0N2JCCYDQ#/M,Qb(39YVQ2FQUg+DBd<CNF
6\,K?#.OG=G@PC;36UfB@S<=YL4Pa90RgWN5&M3@NYe)f>+>Q^\:>,Q&0d0e@\df
fd@G_bNQ/U<[.P.V26d13gJ,WVYMK+c2]fP:U/,.e[(gJ11Ra8C](fOF]@<;g.?8
S<,WA:44+.8[.&MJR??8a:V;X2G7cb5,-1=RT]V3?b:WAaNfGd8X.J</^c4U5U>1
2fNaE@b([KfN[8GT6UTT)PD7);B7DP49gD2MBOIRI]&M#EY[&7Td&,d4^&AK8UH1
6[^[4HR4:P.+<)aY=VGMG@=g7\KT3AeYB/G+,J[/64_+/F:S<X0J:+d/2J??fDWV
/ZR^OM(@<7E:e)FQND?_Ke/WBaI/8SYNOZ8/9Z#6A+bFHVO3=C)[dV>0?RB,]KF>
-3fdeX5VK4B^.8SWPP.<aTO>fa]7@<+<]2]J7Ke#Y5IURL^KWc_0V+,SJ;8EA8dc
?\+.Z/H9=;gQP2f<HM<VaLG1Z50@XMJ7-0U+L;>Ag11e-TaI9;KIbJ;><cabcZZY
C]Ja2N3]S,Pg8,E5+G=69P,a)c6>cD.a0-F,G,=g/-be/JD\K,\02\[;K?P_3Z)K
=[[f6IY=Rb#R?d92eD)64??b_=O_HNCD8Cb7^@<B[0@:EKDF43Z3Y^U98JD<:NUE
+7<=V9Y9ML.aD#9_e;9MdV;f)F]9_<GYaCK-77.\9,5+-\H?G\[U8R@BKX][GQ1<
D>?YT<WRG,+[?b-f.8PXDPU=7b0H6N:+^;WXJS3@S7&F5P_8+<,@7,-1.e&4>Na.
>>3>X?e.H)50Q(T+_+::]9Q\MM;0MDdfFCO?&F/S:T\_SGfF8fP7ZL[(FH_<[IGB
=MR2?9;U;4SJR<[1Vc3cJ]6:OeUeK^Y0HWX7@2FNfa]89I5/]>IAHB4]O+OBVU_)
JW0Me+)?T7&8<WF/Y+M9_C7[OZ_I4Ga;Z?NJTSC3_FE[^<NS?a<Ag8ZQScBN@AN3
3)Gc@17cW2gE=F7]:72(KJ/SCP]SGc3(H84>/(AO_[)FL^_])g&]fQBE1b93QEJ6
O6\=4GF@3B1Kc10GA]#H#1gT06[XRcI>B;J]>#90?8BNYLbF\&4SJfWEWB-UYG=A
_\R#>[[&9__?6g:1MgKd(/_2gdM<5c./f;)8c)&PDPW7eC1T4/BEN4JJ3fLX;N)_
#XRe0V.;BK+(:\:M5\5H.5e3gegN)7K-JG.:5-42)Pa8RU^HM&8^=G<5>G9IWIG>
W3>W+g:V]F/QDH2LRK>SL4M^N-[:dS9ZKC_&-S?-M^TOf=;a<.DR;3,I&;Kcb)\a
ND_-BEaXMf<T@00VZHKbCL3G+dD+AZbHeMZ>.-1IGOVGNP4EQ]1aQ+H[c=OfS3K<
V0Qe,A,8V<gf9EeG_#/9I^5].FKY>=DX^Z++a=f^F_#da]a_84DJ=W_\FXVH:_3[
2IQg_M8XR=(3\X@3NHacSRVP]A7->--.0=ZEeL_YYbTZKSG7B5J9/WF33KdJKBC?
\=b+X7.B0(YaW0_5T-f]D(C>1HAJ\5>=7V=(_^>EIce<CYXHA,PgW5D4^&gL;)&@
>Ib\NXde01@FWBCAd1Z8[2>fWUD&IINVGN2N[@d1)#W@E)?c5&_[2G2WIQ^9M1FJ
S3<G=Vd\KZ#R&T2UVF-.D(a>Cf(H)C6GJeNXFbIJC/7.(ZedZbbD+X-H3JC8fe^[
JV22TAd9:=VB(;OS?G2]F.(QAA<>e:/12R;\:O0&BQK<18fZ>Bc^LL(&aYgSa5>:
F#E5H/ESaTC](.bf-)ZBT\a39c/@bRN;MNfN,5NX<_-R[-1DW70^D5Q;E0>=\LTa
(Wd+69RO8bTA,FE^>><U886\Fg80;#0J+/V0TZYKMTV5W#-]@gES-]#F?J8ZHOgb
-GEY_U=2B0;M[e(cLKY33L,H@U37c3BS92F>ag0c@@Pg3-<Q7RO9?SR.UO>J/&E:
]=7B_[b7FgRT+Sgd(\O/A@MFgg160b(5JX;)X-<aC5HFWOJd8B>@5O82.+3?f[[M
[F+8-R)L[ZDMZ([3VC7FIMfDeD2R+O9073dOG9\]WBeI2g@@4^0LfDVBd@_:^6I:
AHW2.^KA[eJSf=@O8=I=RCT(d-]D6K>N.#VHLKWD2RBL>K_eM.J(_4f5S(d045&H
_GaT+B44-;#a2XLcaVUEf9ffC):8/23D/^5gg@PVa_YHDSD]QWdJ];)b9+PeAdPK
@C(C-;ZC#d3HPeEBa:OO;\N@1.<):ZX[H\?DFKT;3BJT=S[&J-X9E4S(>E/b,e^?
04bOcLL:00dIMg0-aNHaT:.=Z_CC.;Q[()ZO&dC^Kcf2AC<=12J\TQ3;NS>Xd3c5
^RT7YgUeN9XPUII2>Nf@5[+??B=R\c\f#+WSe<ZLB-&AF\PB7JNO0HT#&\M-WB,)
Nf:A716]bg0P&@MGG<[1JSQ?44U;NG.9<--]#.cP;A[<9)2eH\D;2,=&I\411CF2
a>.,N:.+3RXO61:X/B.=S\UfAI>\Hfe)/.3E;8/IgaJ?a>>c#I(=)0S[WW7;XGZZ
^>G<<R.WU&BZQ;K<F4&E)IK2BI<?\Nb86-4X:E-00a40V-YZ-NK:X:,d:SVAbK/>
40][,gA0BOc&/P[gP);E0>Oe&#LR^._D5b>[#cae/2ad5NH_(5&G?.K+BdC+3);:
2@P?T1_(TC+BBQ7RO4/VaUWPe5Dc9L#E+88eb72S85JP]J<\/.6HP8W?VX],GMR@
RfZ/11^I32ZB3W?T[I(9&\G/8=W1gF>.1>L^UYdP8Z250PXEfF_MJG4TOQ+4[:27
e==QE6aN6b<KBV;C3c6:HG);X=R7]Ka+ML_?+_?ZbL/H9_,&YCbANZ]T[aCZ#<?:
N>DB<0R/5e0Q3:VRKRb^<HN/M30g507TP?c3<6+6\[5ZYC^d[P-+QKD<LL=BAa4)
>?^DD-.6X:CK&?9IRgK3F/aU2DT&C-X]Z.S[NZeGF1/^TES#S+T:dJD\#[-H09NZ
ccGH=[K9,&>N[<O3K?O:L?ZQ=S(=&MbN0_5EMP1DYUFO0;[X5cKHBEbg/b+K>7,X
JLI;f4.QdL99:Z&(7UAS61LZc?I5/HUeX0+RU,e8V007C4Tb&5\)J=JSd1I5?T1(
6-?--4EQ[ESAWD1Y>&>0#+KE04S9+@H(gC;+_:YVD7_G7],2TQ2cA[:bP;6_T)1C
>bW^UXJAA:]4=^,@0>0M/QVBcPJ[=a4C7_Z3-A1HD[f-:L]?SbGdO[(^.9:8KR,1
fS,=/]Q[6[dUU1BYOfEV><(#I<6_C_6Zc^;P?f;X(a67I5gP14G2OEEO7+-(VV;>
)LZMC#2<B>S5beAO5B_#LCZUdc=,T?7R8N@=X=6I,Qg,YAfdCZMACA-U(=U8?Y0X
A,?F-d;__AFL4]32/G,2SbKQC:F7\I.<HCJ,Ad4S+Z(7?Q)\c(d5U7W[-(=AQ0)3
XTBV0>;A3e90H2:A<g-=:XXJUA?TNPcd^RII5O)AEf:-fK;4JPGU[O?M(WFc2>L[
TOa>VU3.08/5USUW04<.+e]CW[J:SZRRK^,TN&F)4JbK:R39;[cWG:)>ATZK<KR2
]c/EM3C=E.<BRBLKfOIJ)&RE[A;fVU.HDTUPR+Re[#U9:ZO;fO2UKL-QNLZ4G7/]
8=PO>9236D]\+aCI)@<D^]-:+M:(Q^bUIU).Q?U:<D9_<QG.GI2eE^G.QT5VIM4S
e<#0S^4-GUd=C/\)6\;Ef.+L[I(OX^D#b6JDFQD[)E@6V2)5UTY^7>]_77A,4c;B
N=dL&>/5K)32a:cg-=#@7)b7eR2W/0@>8._;]C#LAZeN_e:X#.CX#F;D3JR;0B^.
cJ(7L=1)7TY(0/-JP[V-V&->.6HO8VKVP/ec9I0dZMS<GgBLJN&YB>CLd\RX-C,+
VC=E5A\2UgI/-,HD?HOEDQGG&GGS=9[.ZbM0QVJ)?G:R:UM-PQW8#2VK]/d-]O#P
K)MR6:M2<,KCbHe5S[B72]?UP9REQ0LF;SYSEU4H:+,Ne-@5R_^..#;HH=55YSRD
?R;:D8=^SO^[:8YJ_cU?6B]R,g=X]XJT-b>PWg.T4a0MHEH<CVdbLb5G]O0-(7Ce
\^:(X)K:J,g/K-.5R]>8Zf+HAVK=\gK9_;HW4.,]c?\R^&IAOF7KYH>_.8>,6NBY
,6>W25a,(Bc9\8JQHCPgN/_G1PI-)e(9\#c2d+3J]S;OcRGTdZFX0F[Me6@OFR:.
)74bS1++D=XQWc[8J/^QNF)E^D6-L.aM&fS24]XQaKP.4=CR&NAUUY<:MXgdY2:U
UM_ZaHEF/.dD457T349TMHKCQgdG94dEK=(90,:,[2d_91MSg+N?BY^>\ZIZIU2N
+81eA(:afE@=J;LBA571L>Q2F#\K?PZM<87=58NMU@a^Y9_ZQOfD6MaTM3F5RGbF
(Se7A7_7cSS>f1I<#7A.(/48K?.e<D,<VNVT8S\86#d+6>NF0O^7;JMU)[51:SYK
:9QE=]6_07W=7XY4P>K@P-1FCHURP<+E42V[V)QU97MA9C4MR9TK8LF[[[5TN=TV
,@-+#IW414-[dBA+NI.V3\1Ma);A9]9>/L4N-e5,ME+ML#7LQ2EaK-\10NWI3/_W
WVG971[aL]/^SWI/6B,U<>\2_G/ZS4(3>V.QfW,,fbS@PH,a4PM,(AgCQc[AaG_J
M_Y+P,dWKJ?d98R<>S@IW_:S;0NK/-\V@=A\DUO2WeRU#M\-Ac.6CW_fCX_QH05U
5D@MR:@?cb3d_B?\1[2AP<feZXJYU(2dJR]V4LZ)0TcN3@83ad5e94&B<V,57c47
JO<N7]]Q<2,ARO@U4E29E/P(<9K&^bWD.#BD67/3,DYB#QEN>+13X^-&7;GIC:H\
[UF9.SaD(#&=B5E]dOK02/N.1&abOJPdLd57WbS,DD[-Z+e;bD1NKW5#U?6W-+@5
>.YTVI=fCS-JV_W;LD[3/W/E^3d/SRYGO6^]^+<IM1VWQ6+:UGe.H=DNSO?DW_f[
^LO->Y0EDG,ZO7fVA=A-:3X7+G=V;7Ug3)2B=\GD.+[6T(Ue>f0UWR9P4C52E9F1
KIc@KHM@e]g(=CA>HZ6/C8bKP^P;=4..)^9U=cC.(J.<IYaJ6UHE>20;IbIISPX?
QO+WI.6NL-J17Ab^e+.VZ2d5,W)@@g;#6AUO_Y)f,E4+O?ZO/-5NB_[=DfS4^dU8
^7MJ3(<=&F@^/CQ4d@NBX9X?[021TS^.2f^e^#8SEWPZ/cDbY.#50>2E^8IS,2?P
+-=&NR(;1VT<?3QT@8O2a3^;H,e&MJ=f-AX/Kd_O9fLa8UY9@8?SB0YKM+eKeBDR
<#3C.UEcMW&A7WA)a:6eHM+bNMF<SU4ecS7ZD.\Pd5UA7&0;FBVV/?YQ^Q6_44TM
4P]DG0N+C?eW.(bg&6H-JD?X_BUb-6ZE&bX80+Xb<V(G_=F/6--S;57L-=PVDN;1
+gH+_))\/=bc7@&&Z413N2ZGgLH0;GSV5F-eNBCCg<KD7ROF-C:KX?\J,GGJfUI6
]2WS+6C:Q#OE.T@f+=EbIZJ3gBc#SOW@KJ1BSdL(D&;^>fVWTcHBYGYc?/Ce9RP7
<[dcLT@dL?4UI9g8[QY;.eB-@G3&1[KB:D22X4<\Y0GbABg7UBDF-GSa(Z+5=gG=
B(MPS1W(H[GVMcVXYD,_3S;@RRcJ/J,7a9bJFH-d+d,d=GbHYZH6>?G-_;5L?8(@
?3I1H[B=99>OKRZd?#66QgDVQ,X1=(#K:UDO@DX(@a0Df#8ZO?Z@+D&?QT#@LF,?
ZKMHH++EU+SP#H;EI)K0T>^@Ya\TH[I4[f)XER3L>CG,#V#g1IEd7/+R#N^-cKGU
JfHDF5GJ,F4\DS]MeI4F>RRNcVG+LdH9,CA2@IF09(KZdBg6(aMeKIMM>SJ.B&4=
>UW]L/L/W7-MK&-URRc#.9[09_.b5a.]FI;7c.>QG8K[VC[F]_)2LX^_BJFB@51=
WITb:1afQDHWZeU9/Ub;1N]>,KcIRJg>Y4).LR=4g8#02Z?<fNS/-Y=K&P/++D)J
(#<L+.MGOa2MKFB<M;K<T1OT0>^a.Ib1Q5IW-cYX,]WX11T[?3bI1eO;B__Cd0I)
L68,G?EdcGP,AaK9T3(OP:M0e-Z63ZR5g<Db.X+,88>OSQT/?:gf_[fGWB;E\X?[
U6X91TGK\VG3?A>DOQJ/4gV6V+XeD;dJ)(4FVDGHA:BYO]E9aYG0Fc+W0^V9;<LM
?A#.@R=YI5bJf^&#g1N(eCCHY#^<F,B3<J-8,,e+I]58#CB#ed3^OC/]3P4cE(4T
I<#81K+\Pf9O42YeEYA;R9]R9B.EUL\]#bV/20QY&S]^@OAIdfE>&a;e/D#@7D+.
daOg.N6HYDVX:?(H^HN/^J@PZJ7,\R34&Bg7[Jf+bf=&?1c.DPa)Mc>0/\V(ZZX]
/Zd;H#G_#?YMG,;_Y,6c5OEE49I0A7PTN1B5CdE^:R2)RR>CD#HPA>Y@4(ZGf#f9
fb;gZ<^3MTPBLS9VLO.>>K4TMU.NAX2+33#aA(I@O,a[WTH#a6,5?Ba+71_R=O/f
2<2.HWID;F/d=B6F:&NBCbQZB?/GW(:C.1Xf9V=3-6R_;60/H0JQY6.Te.R1,(.N
Ydc-);:LQb4=,cS;Z(LRcbUfV,QHM-L^>ZEEb;B6AE,I]>[M#/1J>K^9b\^ZOG[H
)8gLNZ0#RaMBcaFgab7,SK[RWOA[7<52(DgYLZ_P,=9P6ZLI3LJI,D;P7ZP\ZJ(J
3RbY6Q3ZYQ#:8-BIcJWSN;>8f4);a,0KOUW1\TB6,LEYM&6]I[5LK6.;:75\<b@,
[5-+P?=AcJ7X#+]7#?eEN;<[gI9?>X0;9Q=(9E7Q7e8,fM:E:A6G+b\5afQD58DK
][VRfB/;>,I2gUDTePVFd\^2?#g9,T+&a\4:69H]3()Z41(,2Z_G?^Z.#)[6AT<a
\2C<PR9?\)?]D;H1DHdGC/YGFJ6VXEP^S^B^70MMf=RYSSMP<SQ,6#TA(8TC]4Z/
Ig82BTMZ4MPfYFXf?6D>R)[+CVP;0P<Va+f,(cP:.P:_Y&bQ-+Yg06(3BBRBG-/T
JU>VN@(?c:3768CB@-FXKJc81<8d2B:7Ze/b::Q.^dL[UA8N41YB1[U[]#Qde#S)
I,P-2-e6\CL#DT3d>9KZNGf>aM[9#=\8df&+JD5YG;]C>A?eLg/N(g2^Q4._/=eg
53<W2efQ4C]\S0=4:B=/@dETR-3<L[VXIPOfX_N&-#28DN-WQ0H733dfDbS8CI_H
D[+0,\0P[.NFe11:RADYGTC;e\R^6XggFR)V[=HJ?dM7(a98a<8##88-I1\EHe=Q
eA:CEBKe<KKCO.<?+99\#Md])4SU9b^N2aBF><:508S-Z#U_3Hc7>9\H=EG)+9FE
b[6bR;G;Vc9@T:1b,HCPBLb9dR<90GADVC.bYUWP83Q3O]Y.[A[5,JPDRV=A.KOB
<,34:5?CW,aTd^5Q^YM<fC,,E<LAA379:8bQeDEN6)PgFM1>&C6Z=/ZUNQKBD(03
bX-V<8YJa1JVUF&_NAA=1^KJ,QK2cG+Og,GW\]H&RH?\[]3[e9,O_(W?L64ZaT=E
dP:_XaIDPOfE4VKW48F8eAb,29;D5^0Z:JIc.+G6fgS2025GgA4[<08;VKHW40fO
S[X9F)8(7@,V,^O]2JG6eg@dM54g6LQ4Wg(BLXYC<4#^56HD09JeEP-.g=(E@:^T
RT5gXaSLHf;\QX6Z-7,Z,C(04GTA^N3^F--d1RgXME?=;EMBMEdbfIC3U,Z_-83I
I7UdL&D+MR9?A7YXS,QF.BUP2=GSb8dI6A2&eR&.Ac35;.Yg16H;L_We\G47X,-I
,ZVT1#AK(NSB^[7&2YC+-)]3Aa/O/EL7]&1>,X4_L[514D-9_78c<(KSKX>L_d]>
BI34F?fBA=5,9.;UWS23WS?T45L@1O:B94=X&7CQ)W8>39_YbMM>J=X)[>dX;+UD
BdP2a+d7,<b<BW(<>AOEEe850@^Q,>_aW?&#V(9@T8L9a^8T@_1A8:C<2/BFEC1^
.7L=cNaJFFXN#c&J@/YY8TYC?TQ.Gf4^<Keg(<7>\:QUB/4]HZJ^QaNJQUYaYS8)
\a(eM,>8B,,e5BZCY6.HQ2^5ZYfR1_cd#c:T,d@H7cJfg5b7LBMEH><Z7A7c&]>7
,<7d]B3H6ENeG8P2G\BI_H4TUHY6>QSL<SEJ]R\?Db-@;:Q]NJ[32=M7]:0C3:F^
g-b^K2(Z?<bB2QTab7HPTY?<eg\OLYB[NEf[9HOd<>[N>GZ<aR:9?H@2UVJC(8T6
7.7U_AZ6aW#>f.CcJ@7<I_H4NS:,Z/P^6&_ZRW)^(6d<c/Q(eF5Q(OcHc_B.<@QE
.G+FF>5Q_Y7I5bRK/>/Gg+=Q&LFV-Z9f]T^c@/T6L,F8U1BOCI?VdUcU=)dSe@^B
).RACJdL-)_<d3T5)3P/?Z9<N#BW;YPWDR2YE=5@[>IAJQ9Dg25B)5/[AM:OR/AU
CW]PcLV5X_L)@JgbEOT@@((=GS<4;DRSb4D8-2T#7cDCgWEXKB6IGd?]D)?9XbaG
/J<8^8E&6_]Ie9)c#UY6:Fd=#8^J@R<&L7;>?AU30,Mb\:/<7Cd@Z#:f,),TcNGP
c/.,W.a73M8)H](BQSe&9I;_U2/]SfE4AHET&(YbWa0;A(9>N0&8NH)8N31fW7+U
5>3fd0R22<29I+fPQJgYH:S^J5E2G4T6_e5,Q1,4dI)SQ[MZ&b<Q?b.Bgf9;I/:.
&KDAL:JG5[e<Ne?gGU0PXK_BaCcMYWRTX\/]dfE64[Y^MY#6;;3TbfO4#;BJ(>eb
@MRZ?[J&>C03Oa#;)GVdSXA18<\>85#OD1\1[32HX;5Y,2W6+^Hd+56X?=>D@V#X
7OH32JN]1ZAI]3L;_6-D\2=Ze^IUIW?1#E<WM&Ke>b5OB,c4+K.bS5ZYbc^0AR3W
M(GXG=->5OLJL</<I1./3bdg#0&:aA0\#(OEO0A]VGKN]OTY1We^_HfF:;JS764]
4&_e#d(cNU\TP_G=Q+b.,@V1AfX:gdM4.ORVN<@&+B29eT&H/80:9.06.;8TbNd1
)_g<)TVbSNA3E]=F\VRC?>O:LdF0=O^6bg2WaP00;C7B//A/X0U-HSa>9QfNFWVB
9FK5TO=QF-@300e<(a+Kd)441ce?F944.]^Ec)Xb5\aHaC7APM.RcL-GXCWW-V3C
cY9AXE7<Fa&G&&?XGcDLXF(\?V[JRX-((JDH4WQ^I-1T8[4<Hge.M\,YNB8(1^AD
L(IZbNFM\AD\<b5<P#3P6^[_CPLaK.?RYE6,C[@V/S^d=DAB69#/D@g=fWZUT&Ef
^I,e8]U:VDAWbgJ)JDXY0/BKc8X+=fU:-6M-JcVSK4AZ-4<@H?8X\<4>G//NFI5R
LRd.d0aIKfDP\gS8SL(/QGLM]1=3BcgdL7D:_3P1DcWC.L&>,,V38=@c(Gg(@5JI
NLL2R_WU@:(]L1WWX)aI6V-DI@SG87JK5C)gQK4[6^Lg(f-e>Y2\.25>IP#Y9bdV
02JfN\8/D9HSH:37<;,MQ?#^4NH_OM&:NL3Vc@,aV8<@[>\C7H]I(<3.e7<RT>ND
#OD>2[D:dJR6P\<Scb4/?M?<G2(0#C73=7[\Q#IUPA:6@-G#(]B\2ZbC0PFKeEAH
[=HVNe-;LJ?4)XE3>9>H7G<&9/D0a[@-0L9Pa])_>Q=PROLE:C(3R.\HK(PUSDXH
Z&QD_)NI.GZE9982V>]\U83+#0?B:H>;1,=R[/Q&ZC>e0PJ0Q:+P0Mc)UJ#[GPH\
b,(]MW_@^IZN^>d@GY3Ce>#/C@M<&L15f[5<+T,LG)+8#7Z>SHFEEUS]a;8EW2C8
c\#7P>R8Sb/VM[>)?Q,B)/FT?G2KMT7H3L,XZADBOTZ7/XJCA1TL[BX9&T-]MQbC
4>6Y8#.W4adS;R0_QL3JB\(.H:ZYQ#LbML1_>XTR7PeG+fM&II/-R7WQ/?d#[V,H
7dcZ;<AW1=(EW_OHS(QK\1L@J(Z]F^N]Y0GRT+Ab\/C0H1I#SFbgG#Q0G@5:@WUI
)]>]Ud1=)J&<J<3<@<>Se6_J0EH<eBC[2W9^E:V&2@Pga8)JF;2=^5H2+aV)AEX)
U+6B4e7D1K,#5X3e]..@dGX>-W_IWGff+d/F=bN[ce()-Y3U8P,@Oa_,XB5T-C(;
CfE9-A[-U^(HZc&N#(,D=5:+(MPTE^X)18a_Aa2g?_=4LB[1Ie=I053GB@(0,)0L
51G\bE&Ha7:>C=,c3<&YFL3-[]44B=S;ge15RL;DR1[C@P1#W1R7+M3VdXH-Q];-
>dK&?_;>#5;+&?Qa_4ARS;R.PFAK/4^HdZ>2e]0<<<6[QY\9O+g/dB-=#6gVR@88
WC>H=KCaY)OMVIcL9\TQMK[Kg,]XTL0B69(aI;Cb-OT[KE,3JLa:0<U6V.=JcY.\
7L_f]A1=1+HfNa@G09+1\GRG2YP5/f569gO?SY^ZXY:=(;FC,YX^9?VK0.M5eT#M
OYHE_Nc.0:]Q>@Qb8>aWW8M#G/F05O]OR:[5d23C(;c65M_\8G-+4&R1J)WGbL&2
WH?>JQN](KcX7@E?#F56V0+X?NL;FZ[;/7d2>_PR]MP]9)@-,E(.^/;JGAVMC;1&
2@]_:8Ua/DU-Q>c^P86FZ+G)-C<C3MV1YK)Q(H_;cHW1#JXI?TN=[#VcRa,>M6+c
6]HOa:2gfJgUP\:e[F#MdZaZ,?R;VQKQ]baMW;1ZJI?E@3K)4BAGC2_&Og0]M#DK
IO#5BDC=;<^.5Wbb+3D&FDFBD.[N3;gV9S1E\PQd>N:+Vb0_Q;Z+a\Y:KL]/GNaT
g,;)?&&#1OK&cg7)2^;9:/fb[IBIbV18f::d&Y2N^cO#D.>;G_DUFO,KY&-E5DKc
-@c,8TfJK,C>WI40_GU>0TIVXH0R:HHG73N>@6@BE/.b=0]5PK=IV.M+g[#X<8.O
KJ;+_A^1f7K3&D2Qc9)#,K=5f&1H<)^F^>8)3)1Vf.d,S>eA(QM,R;gT:M?f/1>P
DNPP,BKY0F(JZgVf098WF)VYafN8UM>X9H9>^4B0(gLOV@GSA^T^-/[>#Y@8fXL[
LIB?4<+86L3G=TUM&+\HI<+>\SIW16;CG[PX6&>S55XaID#SC5P\BA^IR-9M_^WV
N]f+WdfJ>C2TGIQQ5>+^:M]8\Q#?-3<9/Qf=R3:^W:a4RgVH^:H=YY[.2R=b<#YW
1D3@GXUSDIR>#I(5(6.V2IJ6LJdUV=.A\f5TLe-6f;NG6[3RS32c[8GZUA>[HJ7e
Y,R5Y-g6TZXC6/.8g6g,,92D=(9SI\\8[1N;1\dT8gb3ZPgbO)ED=C5?Za/ZC6b>
WO^F@?gbeIO8X<J^d^CVd)NZ/+gYZZ]H8D[DA]3Q8_B@9_,c#,(/f0>,P/R<U1bN
gXH.-Pe5=7BU;E@94,>W/2V/R).#,7^B?P7fO?JM_TfH)g)08T,c@U^Ed;NU)@.>
5[K:\XUJ8Z:M[6>P2-745UJ1cfR05G?IMQODBSKS4Q#PKX8\XLbSWRTA;@T?-2bE
GW2R7R2&>0ZZNH5O)C,M>e2MS47.<J&9=1Qe-@c]550QZba6&V[0SC[+f]IN/X8c
<#TBR52]F;dNJf<W,Jb#>^X:0R8;<U2Z6,6S^2.N.HJ32M>>OTaagI,BLXR>Y@(_
Q<ZKA@(D2RSG+GLQ\(B<EHM2dG0<8[ad/1HFf(BaNOB5V\;_Q/]cc5g_06a/cF<O
]GJRfW\a=U6+ILeVWD]WUI=C+E]Y5T9I69+gNIZ)G@?,NDC7_e48)Vd.[bSd/@M;
5_11g)gLOG5.5#TRgV(3e-Dg6N^BLLDVH=4):8TTWQM8(_PGFMK3#2M2VZP\QXD)
I\eYLF7C]>3&W2U=BB@BN?DgOa?08^,]@M[JUR&^,8H<M07WRUfg(ag_N<d>ZB8<
Vf#B+I,1,\;=&C71R;&]YOM#1\7;;=;TIBXC:+T[3_c=8UFI^,N2WD1(>La[e.d/
8BJK-)O)dGE5>;::OC)7D>?_GdR-JP2?/XYYZeP)Q#]5NY;B)IZI];dT?&?JJ?KV
g[Z.>CQLbDWH09)Y;WQ:PJYcXWa?6/TI+GH3.4)?^-Q<Fb2UN-d&M8_BJe3H).9:
8,3LUe]N6FVFZ66W>R#Wf;#SL7=KcUIY&VP^6@9>4df2=Jd^cH5])e()fU#JR&dA
UGXEGCWZETUHEBb7VeV@79H8F>LG,)&EW(QJ&a4^U_L(X:EKO[8Of0\L^Pd=dR7=
/=WUAY?R#La0<7M]_Ke(17TITOA1^Nb=WSX&<6N0\LPW<>4)OAa2UCAS5VWJIZ)[
AU<(cZ6[7.W(,6EZ4F^9NB>#CgKXO)aY/OFM>Wb3D-2(MHX19:L(PbDPDU/gFZAe
=(&S^^AJ[(PMO8EaBC-4XN/15ULe;g>\ME=JC#-;[e7[KKc5,[E^RPO,PE(P?eH:
W=O86G<[^M:]K.5G\9UH1Z:<O>(5@6HAJ\YQ.Z@2/TM(93_JL_<P@#0E:,8W:=_Q
;/Z^B:gU/3][8]BUGBg4(R;[X9-WIa:&QAZ^FHT#A?\XPf]1K>VVGM+YY>G?<5Z\
c&C#MMIc+JXgTc#[:E?_OTT3E>ZW90W?EKLZLZ?[SLR:4O>HB96>@#ga);cF(1PN
EHIESTI)+W^&]O(^ZN+4?XP;__#g2GSJH2N#[geL;=LV+eKY]eH;V4Vf3gCZbJFY
S7OZca&(N3bR#G=Ub:];P2cM,KX??G5:EAC+&@WEH-COK+/,XX4H=eZ[-1P;<D^N
L,[-:>E:Y>VIRNUgU,@&&GL+Y:gTgfBKO)#S9K]7X@;VN2c^DbYP>?A&D2&ZXX7S
./J/NS0Vb<W7G6REH>XT5E__K;U/f-<g:43EQ&F9=.O_+Z<Y9WX.?FU[&K<UAB5=
2a,YFKP49cDa5[>ZTX]e6.?)HHJ)R#W4a1;&_35#I,g2#HR>C3#d(Pa9QR,&?(OL
.ZEMcf@gH3UR#F&:Z6]AecC&DYF[87PJ_&FU8<3CDQM;Y+Fg2=8/I2:ZZPVSX2?U
D7cV+]J]2CGWGL>1TXbU5V4feI4V1b4X+@^7FHM4d-X1G&<@LZA+-9S3I5TF9>5=
_TF?g6@JDG?OE<QNOMJ]_1<V?)C0,?V+6W\YeG]J^Q8C]&TE,14&J7/EUgS6/f-5
[gEfX/aZ12eUSScH+S4=bR^b2-:)07[:U5fNO\f[L^G@@,7>Mea+1)K<>\)JB_A+
#O5/6CMcD>ACTY-5]CVA]9XJL=gQ^UJMFggRdg5GN<(CcIgV,==V)R0fKKdg8L,U
0+\Q@3M+KM1T>(XfbcZ2+e>?bJM6>#Q)Ug.e\MP?^[7fXS9.Xe,RZ,8XbI]B^>3@
MT25]fPH@IH4T<7P/_F2]X/P=J[Mb09ZP#K-c.;_CcX7W.>_V-N8T0PSPW]3-GDZ
];V7Z/NWS?NdaQP?5X6,U(QHH/3?)Mc.WM0^ZC4I&/+d+-[4cAcS4:U[VT.PF[e)
Db\2VUg+DEO+2CM+23EUK:e(Oee,.Gd=ZN5T7P@X#9;GZ#Dc&M)-)R3;CL)1e2a_
\e[c9(e^B[7#5McR9FS7Qc\d9aQ0R09I]cZ-g/ae\Mgg4]EY(C.#MOIP7Ca]E2E0
N1eR#KN6]ZPe;GE;Xac>Idb:1LFLV2CEJeeb&<]Ec)GA[;&#5gaFEW;,fbcV3YRb
1^d(E;N&(A=LPS#?9P:>.+Xd#ZZX=dO.a@.If8;b[f5R3UC1FUL<I6\<b9LFW)BW
[++/N:7BTH<R=>WM@EAZ:MH5SP+[X9)U2P35U)+B@.Dd1Y54KeN.UO1[VS94IE.T
L-,[RPcb-a7#SeT^F?f3=R-V)T?L#>]>GeEFDG_U+_P^)80dTZ>7>d;SLDG(<J[R
=3B54GO3+3KM_8-LS/JIgVIH3CO72#7-\H_DB-:(7f>IeaSPSSQ5@EESe@MF[8dS
=+B,2+C[6H>L1J6-B4M22EN+OCKF:M25L^KQT)(=W>_=gH0V[DfMSG,0]RLX>dIC
6OW]>0#?2#71MF6=PbSLQX)<>gC^0@c6O2.@)1>:a/.5B\a0V[9^,(,X)K=(bPQV
0Y,\U5?80:[KF])0^8WCRTg,]FZO[:_T[YY79=6TScU;IO73K=g]3)9,)?eg=WBc
8[bG6@Q\MAT2VfU<bCP,A\eJg<GC93YaEd(a+Q?7#aFM.:8FY8M/4>H+=;g>;R5K
&551gN4A7+cR7JU14+[QN/HVa#A6N+AC\VU;J@07AOU0d=aL.RUVXX4M5,R6fRU?
7AO&^.<L5fD=/0-ZX&(S+\A(3=<e-+-2/-4JQ:_BVX@I(0e@c5G8JP&XKbDN0IR8
K9IKg4.B\-QWEe/]OLg&24dIP)^fNa_B8\d9^dTT]fG]YMEE?R?GIe-2(FA+C<Ne
E0gJ]4>X3P:K<g?ZH@9RRD#VE-1^RMc[@aF[N#C#S^]7K8QR6+=33/UM+c\6JZQP
&JZ)c-Y6WJP@e9&#eTcJ0c(QEa5:0fb:7Y/S1&W6O>A/SA9?&Z#cX;29SIAR1ZcM
9MU=-LQV2JI9Y>^bd8W^BD+NL7]XJ+P?fTYZ(<L922=9XHLJ3JPT,\V;STF,F8Q/
ETLafUTKfEJ;ddC>CY3P>DO&IWU\@.gC#eAA@eN2AZ1(R[.,:?VQJ;ZO#K2[(&6\
R>JDSCAK;c>&@W=N/8F)QfWB;f6AH/9OJFQQU&N5TZMaeA-/X>eD[S\IBdC5L58M
g>c2.BUS4TW=4:Cd5e]fY-H1[JWEI&V/C@KI.b((F,+f,&UX-\#>.8YV,.._CQ8W
Q)\&[M5+KWQa#[O_<^,0G#CYR3[53_YCb/)L?+4]+7bf,T8V8eZ_AH?5\V;&dc5J
RR:_QW-<eSWSL^A33E8^.[^V:3d&OI[;AXZ@#?Ea#5\aP[-YYWC.:[/&bN1e?;<1
aMbaO?M(>6Dd@NBgJa+-Q1JW1:\./f,KbQ&,Z+FR#:QAXAReQH[4D@6])5^JLS.d
]V1BOX7_e-6BA^c4GG]KHTC\;ZM^J?)gYV]Z\&FVLd]?OWF0Hf1)W#U8&7LY0FY#
G.f/SR:.(3GAW\Yg3D;,MN114]-ZRb&4dR(C6cVg3bXDH(DIbB,1gKDCUa)d;fI0
^Xed&A+75<;PCAA4J8_)_C/cPV=[c\QPSIbGO-dA?U^eD^T>8E&UPI.6_RcIEH[#
G9;O/E,?BPD678L2VF>g:;,bU#F.JA/@&;#D41X]7@Ag(P16/4,S27IcEU[I+O-6
dQe9&<WIBM4)e1Y0bVKUPTa]G^+@\(-fP8HAPF_<85+]6gF67PG5YGf5-F4d,;P1
5\8c=YZ[?0P.02T@a\^=->)O_XLXbP_a.UV5SG31YPUgcaQCQWad<#C-&_95A#40
THa<<R)O5O0(:VV?.5K6S4I==P37J+8TQ(_b\]W(gLNL))43^2Od909+TQDecVV\
>;._I7,bX,6E9M/,34/f;-BA,cMdHA6Xgbf^XSdKW=XA:9+@U2cdVYc[RO[I:68X
GUd)V[90+#^@#__Hgeg63X,e8S/):Y)1Xc?EJ>+[M@8MOO5[AI4VD09d)P:3G4;\
EBd.1XdJR/SNX).CZEOF2e6<F?2:TKX](-R(2S53I+aT]df&Y:>L@;83/Pf:N@TK
TV2;>17F3LNHIaJGU84fe<\.<<Qe_ZT-#4B-gFM/GN+?AgBQ^R=[IA5dKa=59[cg
<3MegB]Hg(\,H;3U[+3&ETDL8f3fId+@Q2UP0R@b&A/KbKFEHLI;6d/2:^L+&;S>
0)]BbD3?L(J@98\+<RL=?EF+Y2FcD^;0CNaFGf/)6E;=EE@>9Oe>@;7:SP?/;:2+
JM2U4R&8=GS@&C[,,:0gTNN-=P0<96<_S0V\ZARJaa@1<JFSC_.D;056/UEH,b8:
_DbZ3Sg+3b05WS,:-,Z4QVC:A><GCNXf6KR;5c6P)=O5++UFD52eY;cf?(:7V=c9
=MJ\_Hg@&S(YSJ;.:OJR[c7L7VB:U(#a253c;1Y/d13Ib4gHdG]BQ.G#b,1T7J-E
4(UW<K,K9#@f;.[gcN=CP1Y1L8QAKOFF@g._LMe_><Wb#(TfZCTO\@\RY(BI]L\H
=D2a.[DXY-B]DBdBN;[e4_K[=(I-Q659CfK_0K/ED?f(>G<d##G3#S:&g-(,1&_Y
@UV>B)^Q:/;W)Wc0Mc_aG)^XB8NZYFOW3<HB&Q^9?BS,X&@WL>d8E5HU8DK:D-TU
R033RB5-C1G5K.:b<K2-&:V;?NaC>a)bd\-H<0_B&A7FHa(UK[_MR2Ne+[;AOVI;
DU:f:?ZOMIQKW8K_[&[ff8V4@QHIaf>&_CXUda3Bd\-cB3bV.=^B=?DT;5>U95-Z
=6dbB#\OJ8HE10(.QN>-ffb5>Hc#&Z:Yg;NY16_P<91dfW^[fWP]A.6AA-P,/JEV
:4U+KJaeGb;;I:8EIdCS=dASR<KO.B;;6^XaCa]ccW^VA2;^Y;FQ],+/TPR;g/7L
F=H,X=FRB122Gc+S69O0e6fWU6g8BgJR3dER[HN.@=YAD-RU3Z9d)FC&_MTFFV&J
6?@=\IcCI@4-f+L0OaP)8=BG\GQ2YR(U/<>^N__\b&O0#@D=LOfg+M+4:J]MFU6U
X+=VGZ21/B.0e9?AXeK1P;4-PJ\6^a=+6_:2#@]L.<L4@1/S242P(2OAYE?7]>M;
fHE-0[bP/H]ZKWFFGKX.:__1)EEL039W)<U\3+Bf/N<E_X;B]IVQG0@C6gEL2H->
TMUU^5:dOgJT/^D&W8ECRf43Fa@+:/<3fR?V4347-C4a1XG;[,0Of\LC(1M,;W<F
;d0X0X_H3a,gA^=OO<N;9DXFcGXbK[JW9FMQe<J<T+(8P0?0P@=TH]6>e@PJTG>9
=;QDWQ1,-#V2^7Jd);f:&;0T&9K/2c\R?5UO:&Y=[68PZ;WUZ=>_AEYO3([?\XA^
c6QLL4aK1a9.F3Q#L^=fQG,+/HARRa@6;5SK+a(g26;7ZLgOb@VJ\A@R)7OHA#L3
?)3^V?A14HQ1&E31c=JJ5/OV1DS>2G0X<E3T>2aO@LZbNfbL83;P;1(TG^@Uf(Nb
cO&;6#Id1=QIPI8LZMH_(Z/O2NX?T[5J0&dB=IAD0BJ8^;,K&JT.B3[a]DfaKPfV
5?XfZSP)Z^X4^DP8=0L[#2->1V)_g5b6fEdH9@>dWR[FU4MXIYM4XX+AV:#?H#[M
_H->GE9fI<QNcT^Qe^UFG@3W1da:M^N)S\g2^NF<C5-Df-OeXaLF]HFNK;>5W-Z:
W=5:)XTY@geDRdTf^2gcIQRKPS9^UD-XGH)(0,]E5.5;QR-PB#4REV]?)MGVW\/U
.-+&d?)DY[eOD]=->3J9-SJ<39B3:Zc/C#E3^c>(SMK^.+2&.BAKBT&<(URGb4CW
f;3]VDB=DM44TYUg#;gCYO&cILD>U]d)c3O1#2-YJgUEVDNEJGD8_6LU[E@dY>.,
@N2UbffA(-6),e&7#:<\Q+XD7QC1a5D(KQ=2gLHRRPgJ_U/PVa7a?QW@0DQRQBTF
PR]YUM(?.]?7]QUb>\O@B\4AW5D7NTHCLKWO8\PbHG+&?91fZ^GfZ&L#bS7:G;=Y
WgFM.#(4TZNAUPEV(.H#Y+USSJ.]bAgc(0,WM\ARVF76Q50E<7J^_+\cWV49:2ed
5Y9S[6c/>5#=PF=L)8_D4/P;#4.&eZf<,gGFA^SVe9:G,dV(0V)L7DP^BcGLQX=Q
<ESPDEA+FbG^=^XORA_dE[b\)-XdR4G1IT7f>@B]V,K7ML?:@YbDO7#/T6?>;B77
Ta(9-5.INLWLLJ+F,E;F]=R))dbKN-GDaYf#DZAGb-M&;>B65VTCOOOG:BDXRXb(
CM_c&O<<e_9A[X88,-/MDMAZa4)?fO5GM>@0Ba61TTEFTM)Q1>+)_U-^;4\:&cbJ
-CL,beRaW/7;If<2,gA#[Q.>X/_1&I9a3;GW#SBS6CKZ-3GS]da/.5fK7.,/Ef]:
>9CM;>]TIN<BL0OaAJJMXT9S2CUP7KKC0)HF<@LJ5(L:-BWVP(@[#4=VDYK[/#bE
[D1IL=+c>a1bT;L.\^ZK8\=0&MI[L@1T6>#A^H1)_VLW6Gf^eN7J<)Da&g\4Z.G9
:NXJJ\B@R[[RB+aG</^e9J(-CH]1_[R9FP=VAcR:ZCI)S6YdAa:gV?Be1D(AGN-=
Y7eG_TU\)Y^7LBHTWO#(dbA.;.8>DL5TBSG:MGa#)+G9,KgA(X9&OX+bMf\P],=+
gW)Jf\3?[Bf\8/6XEHEZ[@,ba,7a(f^O?<fWE,M<)def4Bb2(^+A8Qg=,+:/&/]U
f7SGT47Gb>b#H\7ZCCNVEMTZUM&gVJV0?Y2+9M,11((S.@K/MH-A=OfP-<F92T.U
G<4>XTb3A;J/T#CCNTQUa&)\<V/D>R6=05G#N0\U#)>DO/d9[b:0PgBf\IUD;S-_
H28V;=3;T-Za1AUM(&T3R6\3H.TZXTM4X#/6]69OJ1)YT81HAf(-4JDd[GGddeAS
.U+Y?3g3E54FIPf+g6]:d7V0:E2f3^<S<WC>>e]4HBKGc^SZ9Q8d]f)RRQS;YB(V
XH\ANdU>GXGP7=#_d;e9<eY&@,X4dH^J641YC+P(Ub+]&d4Td@[UGVN7g>V_&-L#
B_G/:&O<8Z)+WEMcN6]I,QdcRBW/,D:SQC1T+R<VW613C,26>BW\c\K#[MAF.CA]
G2g/bO(Sg)VPW792UM&94U1.A33.eVOM.SG31^e60A[8.FdWB(WLWGeEDTD[-<gG
\Ka&=D]gW>f,>]>_J>fMYHXZ83YXO.B\63W:d_1(@V<P?E3F3PVf34@69,+EgQD,
f9&NI;WTQ38cV(^fT11B.^fHRH^_UJWcNO6+HTE.R)fc?[RR6E]0\OHMK-c&G6UY
9LUYURf-EBd<(g8]TSFY2Z>dRaC<[8ORf_-&E/;]AUGS6gV]BY:T2^VD>Q4g8VH.
?,,cX#&S)DWR&=8E51+V-M6MZ0FcWScQ]5:DUS>Ua=HH3dAJCLc&6d\eN#6_M[P>
FQec#b]GW21</e0JY#8ODXgI+[52:YM>=1/L(f;C9cOFTHYW<KOR#A]GYC,McK2Q
M)A7=4e2]NGTdW:f^e(.XYYObW\2HOe2F&77(MR&TKbB7D/UA]=\&OBUZRcD[&>_
LW>fMcG=;?,E6CYecTD,VYXa\e:Q;Y0:S-[L_b[H+&;-3,\_(NAR@Db7K[3@SU?:
ddA=R+5:^.&3Ca#Z)M-@:NLY_PNP).E3<GO-#G0AF,BH6K?5@+Lg,IUKMPE^Q>DZ
;^6N.Kb:J4].,1=(#-1TP8O+IbeES0QFE8Z.KGaPf>)?BKF,U_(:a-NWEdd[6A&6
NJ^4;bA@UWL[N6e#OdUUb:QXR_b,.5ad8A)I;>/VE\>f/^,OXEDVE5>(=B=CAT6H
S[TAZ<O\A-E29,[0,XO5Y8V)a=JWPYc[M.e9:A5REZ87f>20TS4UbBD/LUfJR<<I
A,Sb607L@CgR7+FXBLgZH0FQE970SQ6[JG>,OK_MY[3;1\Ld\/cZ]M:-CW7NRPNI
&A(E-PV^)F6KQV<)6ZK]F].GTQE^^.g9\,4U-6a1>.;](UH_M?NF@0Eb(2--bQ0/
A<?2<&HDM:K<OUfXa4]<ScN6XD+SG0+3aE(bW<>H?-5e&O?138_XP9E@8YFB(:4-
>2=3;/XH,)22B9URMRQ[U^>\TQGE8:]X4g+OIgP8&dQ-/N)ZCD(2ZA;/>EZ9:KRV
7b<9K/5fE[BTA\A1:;1F#G\NV:]J7;ZETIL0)92VX0X=Z1gK+:Q33d^5<eO:E2YI
Y)[MT<U0NE4S+NZ/):a5;DK#)c<5EZ;_T01-M-]C8[(U+BdVX;4g2N)UZ0]P[<([
KbH0dX.^]8gcJ)5DE29\0[I]YdAe9ga^Ka,>aCARC]0RXAL]85(24Uf,f#<;eG.L
AP3;KFQDQ#UK)Ud6N<\Sb2DJL=3G^(;f?4:406\C9X+>GSE^0S:HBcLOcJ(4TA[=
<]</]L9A12XUC<[EBLX:dSdA1gaJ];d8S^(RH.c0-ZC9.2Q;8G6^KO^-8R,L6]^c
C\6/cT&)RSM=#;X7c^2a,:@>.S2ZLTR<f/;4C]?)>#<KTHS5T,QLNIaJ-eOO2g^?
TGI.A86<e\B4+_R5RGHOF0(4A3MDTeE=+I:Zb)H^BXZ8:Fe-??FRWSQ&LCf[&9G-
HDYPW/W08HQJ,8=^[/XG7IE(>69_@?9\,=bbS4RRRY07Gc@20CZJ8E=L?E2^E-5/
F56#6[YOW3XMe\K=5L/J_e7E/:EbQaV2^>&aSSeV=BgKFE5OL?\H+(--=bSMA.OJ
&)Z-70cX>@^GX8[KgR/8\,0.c0G/eI=@:E<T+I&_9MIJTM_I<AaXKK)(91.eGR6-
EMO<a)(AW(WT1-IbI?(-61BC^0IRf\OMAD/S,RXRGT/,XbF@d>08,GUU2c?,dA^e
##42aWUG7_b5/JA+C/JMbX_.FK..cQ^,fQ@UTL[I,&]TO?_[F1CSUH#Y=U1)M<99
W6L[gfNgM)A&09Yd4eDAg^?7WMOGD[Q?^If=&2Fd/e)9@@Hd_f6fWD;=4/&S2BFe
DB<?@6dN^N&agdMb#30Xb^+@E<c1)P^K+=\/V#(&P#fF8UY)>;P0>0\26WM.W<e_
D8f>V<F/\O[#VK_RCVR8X7U(9fD?NB-dbOd,FXPH^c9XHEWf2I98.467HRCDEGb6
V(\b^1?LKbQL2#C;_R;G-738XfXQRL6cNGG-2/R9g-L&<dH]=LQZg5_dFeIE3gaT
W7P=,V;K)fP-3gA)O3]=O+E._dW.cNe\<)4A;/6AP8//3:U>MbW;=ILfJfNAM:K_
O4K2/[2Y&H.USJI>XT?AYBefD.1g,AXG/N?;ZG-,MGW(-a7A]b&L,?cQ<=2^MRe0
JcN.EAO(b,WGN&Pag:]]ReGbB49VU)bV9FBROCMg9c+_b;4A:1YR/^[:0-8U/HgN
Y@UgYML_84>#B_/HVN6Ba2+L@TCc\A6bUe>A,A:Z>O&=FWgWQ&3/(AW]8Oe1RdY;
&;;YZ\#PgcY=LOV_g0+FNZF99<7KNFV4#[FGFFcZLUW)U/7#]MA[#A<()OVKT6[8
+2?S_S;g=?X(H,=.b\FX>9DV>f2+cK=C_0AG@,\9=e;3PVc\)[X<;IMPW^3#^,42
(;JY(]/RbB;<N)7Q+_<W#5&fVIa[:\JW&8b\>7H\Xa>(3;4YKRALWVOS49(MKbeG
)^/-C&([0M/,7cfL3QaWC3(#Z?P&a)^Tb51c&)GB[#^2MN(AM;KOZD2dgT3GJA;#
2dL#D7AUH\SBIV;]/JWR?.L80-@UgJE;UCW5Od@VER/S-Q?C^Af(eIR1g0\=KTYP
V.^V/#>X=\A>KbV0#@&8WaL6C)GdgfHDIQ2^^JF#W5_Z6GY/^;&+WL4;K:<LSLE<
Gb.U,C[<E1I:+UP3R5:10,[1.32E\]J^,e8+af-gDY<X1Y^#(WaI^TLALZXaG/5<
14b5495N?KecQPN4F_AHEGEAW-AbDEdA_M)f-B?Cd@IMJ&g8&IXNX>B-9/B0g]+>
)P)?K5ffM<4TVGA[Y8)F/e#9V@ZH\d(&(>S,I/WK9M5V18=0b2LKT/+ET;BW]EB9
2PPRT7_f6KW2<0R3C=9]ObZM3GUVJO1fX\LHHU\HGB1<GGZfN\Y^FHc1]U0B5a=-
/CK0T\1)>HQ8J)=SMG#fGHZ;6If,b;MQC.>0/&\N^@+Z[fV:2Y<=fGJR]#gGM:UI
O;Mg9g#aKcV-BgOaF2N?S7:S0d@\ECUAW?-9JTYc]^)V67X4G/fQd8@YFbYKT?[<
BZY;UW,<b<#C/QIYD#,5U&NgI2#gMMH=[b+8/7=@P]]^@CGD:>9)[:FaYaOF>@OM
c7Z5YC-R::YT:5@>J,</)^?OB7a.1O)A=XDd3,GVMX>G?55LCdZ<FUC:Ccc[X/OU
AacKX-C>PZ3C081d/YX:L[I[[f-27aOTN0HWSXLA>S&LCP\0ND92\2CG<,KbC_W=
(:_UBTM;GSa64cK=+IT23+g>,RgCfSEJ49gWQA6T^_cNYe5BS1(C]DA8-+/<8>&<
1MG7/-4FET]\Xb.G4.<]H-Y_/QaWYd2BB<AVe+@,(cefC6]VSWXS:V7Q4W-170&1
>Cf2[(UO@\KBZAPM@DX,bXHeH/08BL[cN]Fd@cgDa7QKK8.O0?A_R==UH\RX#VFc
6PE,PY1Qg@:]c@D)2<W:Mb+/R-EQ90b+,#XP3YO\/TN.L(#O8B:VME)D7OOR<AG4
H]aH9LN??;Y1YZN+2FB/QXdUV<fe5W4):I?H1P>/V]YVDANNbM9&(CFAS#;.NHd-
D,7MD2ZS1B2FePg#2GMREPgKbe&E.;6;KWEL],\O#VC-,cR(3MHgEJbIUF6R=T9V
-#DO:K,I)g/AA1NCXf8P^Ld#2(FQ=:7=Zb_5aY4/5_+D[YKORR3(b9_O]/TYgC:.
=1g?M.-R<OB2Tce9)6_YX6-+G5V<[X9>DBG-/(:g^:<&\(0G7a\f:H6Yb6d]:9#P
PB#XS>+Q-<8^)c#MG,#\I.F(TO]9f-6gQAa537\fXLQS/0N?aHa&6NLLcAF5-/?6
&L;.M3&bGK8gMC00^#gC@V_f44A^5a4b/U-U0Y_I?@dIRb)gNJc9Id+WWcHT4a-E
IOWL9S4,c><K.ZcY=J9d;N1[]AeFCG,XJeLT96T_aS:ER+CRM>?IMA[1RV5JR9I2
C)M>(.DA/FK:QL/fa.>3WGf<NTWE5Qa:^H06FSIQdCRg/f6?F,4657L8d5-ZZAQQ
JQGZb/.)fB-+)K#(@C[_b)^]^Q1D^?e4799b\9NN7<Q>:Q8I+M[C5<@FZf:]Pd=L
R/#18N0A@A_1:9-+#]5>L-U7#??2GbJA.@c/N+4]LOS-HN-B@PQKXVf&VZbc(F81
NBUDEY#\6=(/e5BRNLPI?0]HB3cYGF9M9ITM&^U>A5E.K0I.[gXA1+cXO#IYB&9&
->?H:=,Tb+f608V_1R03Z>+I\WY;6RPcINJDcTF[_(8@?CIef(PKGLVWV^QV+Q_6
[C1FWcC_VD1>8.1?\/S,WA8a6U\T]I&1-+>Y5909>2fDe4C[<aIcS5V9(9W9fR?@
eBMQ/OW_;Y<gZ[V=3WgN+X+Z8E8c/.D?E4.M=X1cWRR<N&ANE#SCYVJN0(3QDZ1)
:<X=N0N3Z,S)PUSDfS.;2,cN?X(&eb_6UTL>aU].&)KR97.YIVA+<J#],NM8[Je7
U.KT8ag73&@<R88;1I^&]GW7N^YFB)G\8CIa7?Z^X.]S[=)O0fVHEN=@C1]D3Q(B
=G.J6./VJ9bU3>\K2F0d3B[UZ,7A\1:7FDHPGB_WTAUVBCIF)[+X:#cd)cB73KXE
+:eH2c_WJ5+)c)Cf5].f,bGXd<:7Eed3G=BFQAF-C)Rf1^&I2\[ATM9Ed?D#0AI3
Ac\SD^>M=)ZE/2THWCTd>P-ZY[(+)0(;DWZe4M^1J=&Sd2c8=WM>H[J\SBO94U.)
.4PLSd?EC7D^6-QI1S;M?M@DTQ@7DU^@P5+&0WI2BZALCS+CcULSRc\J.86]9cef
c7+(<ISD7QSbC1)Z47)Z:bI0,F?8WF=:DZB[@Q]c9)1>OQD.EK5,Y@]:K6e>GMRM
9?+NI#(2J0(WKYW[b,eT_]Xg(-:WYMY<AWWg3C>21NQU1LA)9>V+CGK?X@O>8Idf
M4>9Ng.B_I#afZJ01fPcac(_R@g6V8/#54ERc.P<806JVH=?^9C]<2#1FNQ:@IQ,
1T-^.HONB,I7-54;@E=FA]=>PW.@Y[QSeFGJO_;(<Qf0OB;QZC([)\a5Wd,CgU0g
C==@P_?K17\[2CfQ?ZWD<HGI@@g,Q4b=Y0-[)(\:0U6Z[SCWJA6A=B+=X3VDQR5-
X=X90]:^K2I2Zb+0AbJ4EFd.4&E\fN1H#CI,,FSG6D/a6DY=F+Fc/Vb\D<NS[>Z@
5AV-P>\<]LH2G?/8#0MVL;+4^W3=MDD+R<^O=ccXBL3MWed6:(B-?_WU9eV5F2+F
\BJTb#?Y3+81+:fZX4fH_bCZa+Fea888PaFX^E9AS6V@W&Bc8RB72/_C=N6UTIU_
8_Y[KQ--([VH6JGS^#X+4#P?W>,4]a])?dZOc)2c<\;8];XTCE=eF_J<L/7OD681
aJ_E+_19(]RW<\cBfd/4BTdK2J1C<8>429gO\)P;JEDX1[J/cd_[1?>OK]?TJ5dY
(__\MY.<IN;T-)4DWN@;-4<3E&U+1>9eQKK2g6YYQNYB(B^[>;BE^2N_-g>,)8F]
-],[G,2_734F6EL\XRJ=ZX.ASe&=UFGY(;1]Q1H.gHYNF6M&Y_QS79BY-MR<[WJG
I9[+2,QUGTLa,T?d]U84JQ-O0F]38,M@Pb\bC?..79YR.VX;:S#]bC=V8\XVGMD<
>U1KF4;TegJL460A:I)KP(/)&>911#88)=T5L/OMPEfV?:^<?@2EgRM><J3/a1d:
=3BbOdIL6;-.R2ZHA#RV\)_D<4HJP[Z8W0fVOU[5f)QYA424S8LaACd?YMYeK@L+
DOBf_Bc)RLWYLEP^];2bEeXME+e1fac-d?cW(P7+U5;BL?<KD1gQcZ>TU+>IE#H1
#IE\NKD>9:_.c8524Q^aNOT.3L2SV^6#=f4+\R[559FNB,F.dG;[6OQOX&UT(;UT
MS@MFZcB:e+gTL#\QW;LU:8U/)A6VDgU&(8:/;+Kb^fT,O?=G=(_,e3KdP#MfAU/
)McgZLaR/^JZa\6T_d\6#Va^#3^B::(DNP\U8FWH+/4=:;:T-CgC>7PgM=9AQQbW
_K,fQ3TbN2P#_dg4-VAf.,54^@A^=1;R64GUM6c]I.+-dMfEU=eb.-MKPXZ[L;)J
<L?ePK@M@@G:g;gKFWg<_2;8X5&]3YJ-3AQY;W?@GERd#CYN+OE;\IOE(\/9g#1H
EB=#VWERV9DN[^Hf5aLOCAb&]],)ZccHf-a(J9G:_XFP1G].YdSS@K-5XF7G:<0]
Pb)=0_fN#A@d5RJ?fK_,g>[5D4AI=(:=b-7<2D@BaDI7]KE/I2)6A8Kf7R#bGBd[
<,dUfEf+;g(:IgS[,CG=LB]@(71dC164ORQg@FFYD\[ZJQIVa0Mg5PU:1(RY<#HZ
0@_QQb/K?L7@@0A20QOBMD]d77b;@8,E#XVGQ?A;GZ0G)F:fBcgH>F.\Z-g,.CQe
\1I/2G_N7.dM]RVWRVE86(Z:dcUX7RJO7]W8NF_.)?#?.7X^VC2b2geBf=,bDVT:
,-N,#c](ZF@/dJTb;XHZVHb0>g<6V>(-dD1@bbg2.@N7J(N4HG2=-9@IHG#<;<7;
\3e#\IIK@O#[gJ?J+SG6LS(#g7YTHBUCJ-_8dI;90_WBJ\43=)2TYEg3_5:6cM93
/)HM9P.:,,b&GMNBeXJXEY&e/;]>\292bGH(B)aTVQA8UXac<OAA0TEY6fWYT^g^
b4a2N-@K5/7VU#R^;#Y^ddJ3/cI>]B2<?IY0NB/LP1L_<a(Eg;=IMDY_0f4P2392
LX;f:/8KLN.6&Z0:-J+1##)O+-)d0I1O9N@\c34U&UDbZ>Oa@]TWKDEF&7V:.C;B
+@cZQSO^^Ve?&-+@BJ&J/e0V@F[M&Q)?5L,db4g2NRDXQ\CF)12\SH=^a.8ZWeb,
.cE:R<aIF)D9d,0JOLbP-9:O(Ea7(I?[LJg.:M8@L(&[,ZBSW/U:V[NBH#FR8,@&
SE38JMRE4M?@1eEQYV-2.1.MDT]-RgdDd<0X,;QaPRYaCf/WfS4=V&QJ.Pa]S>08
@+0eP?UP:8_:2X>NLE-c@NeBP3M-?e)5I0(5(R+F\HJWU59PSE.P@HP_J.9ET?G@
9L/GBQ@OH<,29UY&4c44Dg\I\Y2UJB>+8#DO]L@f]PWREKO?Z:0U3[e6d@^I,VT7
GMX8EK-8;Zc&a?TL:D4(5g29J-/N67gRg3-#<IeKA#6U:aC\#IR/]72A=@F_.f<H
H74U_5:(+BL<cRTMS2a[7;7ZNa5^5a,Z>BOQ9P5:AM4G(<F)>KCR\:?MK]W-7_;N
GE:4D5EP/&H3F(EYFK1H?Q<3RWC-Mg1U&6ag25+QXYMQd#D4-/4U0EJC^(M0;P4-
_?:L8.)-13[68(c:L:f5IGd8C8Qf>QGVgC?8F6F_YZ80X3Y5XX./7&Z;<f-Pf]7e
e\g4Y.GgPMQ^)=;d8P8.<:^;4g&0ZN@)cfQBPZ7BTfI.DYFXALKF9d:G0UH0#M7#
X0S/e:\E:@F>WLPa6()J54?R0BQ\EOL<8OMGd7V&fa:10\HZ>4EM>HOMI89S8K[<
I>(5T1>((2d:N1)c1OTbIV+N&&)-cB[_7A&&(Y;fJ>He[-TVWDG-/)1@,<FX9VAS
A(PbRN>2_A)BX<0=:?dT)>eb3:bA1<+[JBP3\F?bHCKMD06XSI895N59X@UWJAbB
KHfBTTB_d7UVg5->;AL+IG<FRPP;6DS)3)JSV?R)cC+ZaZYH@+f727T0Jg&0/U-[
JQ=[0TSR.F,.]fgScWB?=<d9GHH10dJ>_BbU,eVIW>O#1aF/O]B;<aa,4LYM&TZC
2)?c&TZ<FO[06a,\ffBC94N]]OEW5=eKc\HAV@XDP(_;T?B\@&RedRR0=21[9ab8
VQ0#[H1>=/9a(e@aF;38M0EUa.J<?V.,&:/N@\^KE&_=,gSBZ7&X;3WY6?.D=eYT
Q(M]5:8M:X9+8TA7[)V?.+<^V1bCK/Q;DLTWC.(+EQc^2I-+,/W?D\I2)SVYcNfU
bb9YgJ\/8NN(4c[(#-AAYTfV)\BYSN\]3KG;c[_K\JdAVG:IG:C(<48&OB[4=UJ0
:8-\8C(ZI3fYWVM.f58)2@O?4Q9G1[VVWT^b(#XA9RL]_M#NU\^S/3F^KcO0=7)4
W<\70SP=g0M=9fDZc6/)#\;LB\B(EQQ8<QfWB<:J&&6L=MPEbN<FJK?RKRW3V[U.
7b9f2d4RQ;gbK9DN<P:gRUCB4(#O&9NDS,\a\WW^SY.YPf\@Kf#I-d9ZHYNT-^aJ
^OQK(g-ISL<KS:,I_.7D:Z,Cb83KgH,(3QO[E]PS1EgI(eU&R2aFIG#c_.7FJ@^I
GGe9#P\[7].14^2H2(Y506+_/Hgec=OP6[>G4)83Qb=<>GaXCPKdc^PLIAOZ_A:6
(Oe#QP0?Ie>>9@]D4T[1]YIXJXLYCd9;&-c.-ISgD,OfB[6FF58.<ZHPb_T1aRe6
TP:Ub>6C[]HQ]bX0#=&OY;6O7OBe][.Z?>XZY13MG1>-Tc]gb1f1[V7I1U_R=R=3
cJ.H7K0?Efdd1K]f5WR\KY+eDE\)\cZ[dYAL7N5@,N)QQ3K?=T@C&ga[VGY7?_e;
G]cVSY(d(\8;&,MIRRAYB07&F=ZSZ=#?^N@b=CM&5d^VeXF@MY^?.(W\a[N]>+>a
Lg3,\b&);+d:_[=@AF\7P23<GEB<9IH#]M?0^7I4<3FeUUGbXH_BYafMUB)A3TQ)
H8<a,02:Y,SQ)D#OTa_]<#+#FP0W,?]R#-7PX;IN6J8V-2:fO&dIU9gAPIQ;N_H+
Y48@+)-N8LG)_3O-^:BRa#GX]7Z_=7@PMUM+^6M>d+I:eaK^CfZ_#B9Ig#5F(>JG
?2JO9b_PXS0aAX:Ec.NPdDJ\7@2:C:HD6c<?e7J@K#P]\Y9H9UJ7;J4[_F\_RIHF
?TBL#?+2ZHW7f(U23EUKBbL.<BHUG_9256QG/\g<M;P0SN<G5aVAL+]0C4JL;2E<
6E7b?BIZR()5M8XUJT;8U&a8Pc^]=T82D>[>=/MXXN32WMEQJGU8:Ec[fe1Yd3@\
>cP^b]]?CFX(0;e^DcP@b9]QK[=\NgGObOa);;aK/\QP.O&22XWc66F<HFX;eGZC
RJUM7?WdBP1X;AZPVF90@P0W^,::f&Z1IE::CX&]dO)\8UIBZ?9LW/D1@R]gP+ZA
JT4V0<M/.AgZJD,[;Vd3RU<BT;?N9+<VAg/50[]3\;.P5:bIBA3L((W=EK/+-_f=
I.Ia2I[)^5(UG8:)DEdQHC<Y,T[))3-PgD7<RB-3f#EgQG]YG:e-:=Z/6f1Z/aV#
[^2@+V3\)Z7D(50LK@:e&C6XHR=5<9DEE+4bQD3a<7=.XFI?CcUY]<AcZdS]:J^V
PG.3EKV:fEJJZ)Kf]O]<M::UJ#Bd^I^VYNZOdWF;5OT\5Z;WR/-H-dW[ALc<C@OM
B<-PKFHdZ46+&BC?W.+]FI+;PO?&8X0U3eCIHA2N[H2<=8BJR=JN^.I/Y_PLF?[6
.EI+f4F@LK[+OPK96=3P>1_JR8#H5@-V6PY;C1fU]/NCZ1?[XebZH/E#Y,0C2@OO
Q3]XSfM@00?TXHUC.:Q,G([;e+KJ9.QCLNEL04_C?eQI]FXLf5@V/@&J&+63=[V>
dCe.N,E6+dcfgN,LF#4(0.LSH.:D7a0YT3DPH2;8\(B\V-]OZ).@OY.9@-<C5C<e
[=4[YJ7^/&LJ9PfV.Bd3@WZg3G^-7R9>REXX,HMZ7[<G-7]/XQNA(RNXBM]7)fDK
Z@_/<a2ZdFH^N7.1:C(+EEb.A(SWa=XY4A,#M<RKK67#.I+A:]6\G2A7[=\U_A]2
bb]fR;;^X)b+V]ZG394R5C5+UEV18)])db^/LC.c-?c(=KP70<YS:IS91/MWE_a_
98[_ZW[Lc0>2OQB7M3=FT7/N.BZf#NWM?^9Sc&<D.6a:ZK=\X[0^?-c7,9Y@I6O+
/NC#3>&c+RQTbC#cLYZ8KZMg:K(3f;9Z0_V@U2<]2ecb</8FJZ>W]+(((-2+DPT>
HTT-]=gf&G;6Z2U>-C;ZZeOVL:IYZF-RA?>)V:3#QXB1^Z+MOP^OTMV\aWWd?PGc
S5)D=>:\SE[CB;N6R>GO?N_:Kb/KJ0_2d-/7bL]OYMR_,)D^PaQK@gJIDbVd@9R:
O1:X3QUgQ;6#cSG&@7\M6+6H^ANaa)JS3/dR[Q^<[J3/2V?YS3-ENc2@>fMK/<a/
P.eFa9b[0aOUV9gS=<T058c+fD2Te^FaLPW()NWJLZ[BX75]@FMJA?ZX35_Y(@W(
><;Y1AMI>7b3HDNDM?e6C#=OP&F4_G:<(W)2BeBJFBPV>ENQC#@gMgWLC,3QB66<
CIK]g^E^NgC.DAgH>XWB2GY5XMAL7S92&R-17EXLX+cZ<-8;(AGaSYV:9S5=W^ed
P^.]#ZK3_e+\gRZ5Fa]XV/]bEB7&BR@f6<=QMg=a;_0\..+XC,[2cF2MQQ^Ee)Ke
500aLgfH5:cQ=/BP0O2QHD-;TTa#\60GFWKG>fe9-6K,bP?:WB(K4f;TR>g\Y1T1
Lg;098dJ?E_-?/c+YE)cCI7a:R_=<_>A#YXOX&E8@]K^>4>ag^[I>HRf@Y+TEBKE
F:AXTD?TJ<#.\<_.4g6DQ2/?LEOY8N0C0VFDa4Y0TT;E5QE_:Z)ebYDXHTW^8OQC
E&4-I,2B9RgHUP8QO-DgRZ9F^9@PKO2/68EPVDSEQ@C[)^GPRE#7efb#L.SU[MbW
X_Laf\MC][E>\#+CfLF9@8];P;(IYgJX,K5REJCKNLFEAIAE>W]KZV<KO(KZ2Bg5
2LQ2C3I^XagG26@Bf2;bD&6&.0^<=E+D,8J<2[J&PN.IM;aIUQJTE[HEcQ9&1-T>
@@G3+N;U;D/U6]LR(@5Yc?9[A<)>=A]>3E5a9QM?R^&+FD(D>A/N,\=ET\>4JL([
ROFBXW=L1FRNS5E8c\Q&GM<<MZ+<=fD&T<AE=3e(NTRDbZI9bP4X)N8[\8ZO-6d^
R(6EXEE>;QG0JEEg7[8I[\=I4])DR3_@T59DIFE1b>X^eLGe5aBW/ZNTfZ,TGA8F
a>3G:F2N\9S^9A2VF069(5]4,N54dJ&39<#VdRM.L_;[^+<]LW;cL<X/cZ4e9a/5
KM1131gV_=>DgfC&N]67b92EB:655a</7Rg#+Wc0JVAM,5<DU9QGB:@/7H\RM__M
?1g+6f(>M&fZH;]eWT6J&?G:8>a7K9d_)XeCD8,D>I7P\1ReF\8:JYZc=M2cL9]9
D5,d6O;d-S?:/B[3\,9P4>-Ub;@EYWW2TKCU54cPH92/K=@OTIJIfH6W.PXF)RJY
RB</MKPb92g[ZeVN2f38c-I)M\N?Z4<eR\5BZZJ+[\(9DbHN=(-1I@UG[WONC2+R
0S60M96+dPb5(CU26SJ(Z)-_M?KF,P>aSQYAQAT<]QW+Q@5GEPSM6M,2H6L^TW2#
b&E4A9HRU/:>3FgY6eOZ8@1cPS_D0EL(MSZ@\RadD,QJCd]5:#J#&U,/?RMf2VSQ
=9NU>PUUI\f#^YAH/C_(UL^5++EATL2GA4DbR)R7PZT/fR1g8+2bU4(LT)Cf,Z>5
[7#(fd&E-6cEfR7V2cY,L^41cF134.1<&,IQ?(&J2a3eCY^O8V]ATM6+);\&:AG#
E-aVVX<aTM^>X:Da.@LE;)AdeU&V(QY@84dHYJ]B24ODQCCFH+a53e,X6H^>AVRO
9[eMPN)Z,eIaAgd7L+5/<IOLGOe=Yf>?:bOdC/F@W#J-&g[^7B5^V0C0BF&2YAb4
eC+e7Z=fB^/L2<J7Z+d5)Y6CUIPA9LOD2(HDf&MbNCVB#<W=[VWQQV3(+3VP^A,3
TQ>eS2CK/,ZJ,-G@#[be+@[<cBU0U]&;ZO.\R>OL+BNe.PFS^E[MR(44,M88?-S9
4(J\5-Oc6//.2fLW9WNL3S6Z-.W13^gN+/\^8528OF3)64S487^ZA6J=#5ZR5J(Q
QV:)?;+>73b@cg+XYcA&J:GKR3SM9,?&DYA.IYMT<E@Z2:OXgLBTa68DQg9OY?Cc
<\,a&e(IK9=4@ITI]1NIa>a.\Ka1<(.WV0^I<RKgd-#=e8X,@X9KG@9\T0ZK&&]E
4e.bY2=3\-RA8[/X4[.FW16f(9DKEeT>TZ0^W,&^(#+@H7&;.bf\8))A@g.^3b0g
6G^gZd4@7:>.J)?0Nd_95Ra09P1.V6/AS-7<Hb+YQ54cQF6K+V\0(2aaS\Q;76dS
DWF5\.M[/g,?J<B9/RP_(4(X@#2Tc<Z[eB>0IfFX9A2b[;-=S,,-(V-3CK1IaE#\
4\)d]@F68EbIF2A(X?T5_801VXQG6P\MZddB.UUEUE3U@?a3[g?]35T-NC]D;REI
1)c[dPS+^RQ1QJ4V,OEN7L+L\Ra<J_[_A#?6abAYG>,AfPW]B7aUQFKAEV+VCTJ]
>g_6f?I_74T#dEP>PV.89BFU\K4<BPUM5PU.SCF2X[H6aFC)V\KPP,)DWfT3VWDW
&AE-a]V_UC,B./4^_OC^WOeC82IYg>G],(gV6c;N,,&7_(?Mg0Q22[1?@aIGN^.;
^7+IP[P8PY#6&2Z^E#DU>ANZe\3@I>FF+(:^:34WEKXA@e)_\78.Y/aEYaBJLDZ+
+6,EU.<OBKL]](G@LGMK/N?:d-<PE[3e\KF(;/1JB8XY.B]E:2.>\QA900M#f_9<
#D&G-;Cb9Bbf?)X<KfT;K,cU.PaHXAZQC[1ZN4A9431ASA+95>JP^YAA)b07QIQ7
&O@5CNf,6BF@F+@g51XD1G=&./b[)\LD=4<_aBCHGS5eF4+ZL?Ef5gLIe9L]4S#]
E83Zge_I2LU:R90d7TPfF3fUPg/<INK4H1;/BU;YAc_/-8QW59Ca@=<g;&7J[YMa
g?.Ke)ZB_3De>50L;W<C[_SXKW.LG6_]c,)8VVeg1?Qa3#7HW/Q],M1V/NeXGQTA
faEV;OA>OeGM2BbaJX8XPNfQfEB>N[X/e(Wg_JVfMCWbI5T9[/4S#ZJfDZefa4SX
SGOL;UZQf.cA3M3U@@FDE0cBU0c1J9gYCZ]W2Sf1=6?f8Q:]LB.J;8#DY():W-aF
/#,E_JEB8EaD21?7]FKG;f2W)dJ(.XYISJ>C??>/d?P]79MNMYA9<YN:YB+^YB4Y
1Q<2<M&YU,^VQf7@V)b1E.W=>=4=K7&<+MR7G;&0H+aL+F4S4GDBdM2YFESG##LN
6HFSVV=CabS\?BUZ22;-I.VIB4V6><b;c9)?]L@4\;/3e(:[AA_D6QEFe4@P,gLZ
&KX9C/1&(@R)<_b]?BJJ/a._E<@A>76Q-,8?;2-/E(N)CN.DW@+9U_?.Z+4(C3&W
7A<gI_bNaS#64X?WeS6\/=b3:A\X9f^W(a<;@Y@#b0+AA<X[C-[T.Y^dfI/(ZV;+
K9Ia-STPF4X\QS?b39C22RYe&EH7^2g^/[X3);5Cc09[AZ,161^^:AeX6H[45Cb0
cJ6XH)Z/#..1>a_fLWAQ./d:8;KdD<a#MPeT:[8Gg#6N4^JgL6?0VJgUN3@(LJ#&
Q6b#SG(14W=gaI)#5,&.GTFBB(gVV14\+c1&EN3)-SXLaW?H8&,g]Pb+M0=/&:O;
6,<R-]-QB(CD_/AcQPb>88=PL0<@7GNLV+A<?:eLggQCICR]S(GZ@X@a.Y-a7WeZ
DE>:YI3[T.U6.Q2FJ:G5@2CgHR1a^66IEB:-HMZ[ADK()dHYe>GFW@FKZS6LA(4S
1.B21QBOZ-M(AT-GDT^,?/?C=.=ZJ^Gc^SNKL_O+X,5>:TA#Z&WS_Fgd=)cC/fRK
]NX9E1Y#U)Q3C:A(e\]gT^3EE2^K.QZR;/L[:>#eJf5+FG07SDOR>S#>^X0355_a
)44f<>=JQ:bH[VK7+G&eD#DD;7DD6?#LeP.J=[[7e^>D3-JV^?U)I,?/AM^U#-H-
UY<I?/QdVTGT5[(Ec3?R8Fe&E+?^LC74VM:Z5.CY#R/>Y:&c_-+V@P.cDC8FfL@c
6U+CI-Q,QE6G+]E95eSfL,WK4<]G,8dQ73XWJ2b9<L4;=>LKcO?XfY6,LQRKUR5d
)L3BI,),bVM\A>_g/&4H03FI/)02S#f@W55UfGKY5FL&)b=MIM.1./EV80]RT+1a
:ReYP6>)^O1MF33Nd^X.F5dCLA<@N69_RL9^WF#0\6e]=3d7FEUeVgX25<eBRRDb
5L<+b_X&07VQ-NVICU@==F60Q#&5BG\OV^-F:VA&E&25Lb&4P/[&Mf48YH5f@6)7
M&Rf0.]2cMbD=]AAA[HU5D#CM<a7:V.6&@JJE80T0W@(/,fKW,4A-IUB>^1?S/VX
.gf=3LcD[P93^I4ZQI^Cc;OABFY_/Y?Y(F[<#B?TE]G5_O[?dK#1/(.>2SLE>3OJ
N[G63b-@S7K]6&ZfEO5Z#4FZ>EWOO00:?VFYQ2\)f(<HA2X1(Q^@()LID\@YQK\O
P_BeYKHcdfJ434egPP?1<g[QWAP[EGVNgcGJ-TC\@#@@M@Y2+@CeB#&2U5d\-]K7
>f>daeC]HSE@[8[W\-]^?#HS<F65PILN;-93D]/UQ)#FX::L6B\)\C=L:D)5f+@a
(&7G/7PUa4b5PA:X9SC?+]5#>.;-BeZ(5..L&#Y6.b9M)M:&#-[B1VT58&UWYb31
7aA2<?PK_=W.YUeE=\38Y/eTgXJfcbY@I/VbE\-9\dDd0==Z+MH)LbTaO32McIDb
D-\:=,9&[R?#^W(G#8JC>TQ=[J@:(4QHG;Pa+RNeO&)/a=Ka;e[52#cVUI0PN5R[
++#f,4\_cT^2VJL0US,[>^AV]7C)U_7817CIgb?GWHBL7GNSP8SZZS]5#8:^GU;8
VHGDYWD@C?2I61R62./Oc1aEBLPYOX0-S2NYNf^DQ/<E-<\GBdIT9,)A^PLY2)([
ITa,[#\NQe3fXH.2=D2>VA]<@P^5C9HM?8B5O+:BKRV]JC0ATS\C&JH?[JAP.UYN
<,QV=eX)fG0#BU]2S1>YdeA.)LeD@A3(eMA9,M5EGaL5IO2W:E<&UY44MZE8(MJS
:]3eT[3?If?A=<;#>]d67a#N[4aD1NV3,Y&#:=SPg8J.Z\I[32+]SCL_(+6V>@\5
R1de(;YfIX],@:GFPMA&Z<&>\^Nf3LN-,8[:V,MP3MF:8)^1Ga=@=8O&_>+O,SQL
-7H>=f^g+/M6>7E]fgXM.;GRVGJ]GHK27=L&970GXRc-(_B7T4VeBQeW5^U[I4C]
H0Vc@#B]B+cb;Na.BV?KVbEfKLe7Y[bP119^MHP3@)aWVJWBKc8>CeZ_1Zg=Ke[;
=\eR_gARN.//H>7LRJMaEX[5DN60aNI5gO7>7IGV)HT0f1F3FHg(b,@[\Kf/[4F>
WNKSe2R&98P>4KfMgO[E@NMY7D)UA.K56&b/(RYN3AbL+(;+AHe)Z5<WW^3Y+FS:
I.#5YY)&SRN(KS/CG-W)ED4E;;:3cMb70S]7F]a-[Q4cKL@(VJ:gZG>HFMd3>0B6
7@TPTOE,G\_=AID\:><B@.P)\#>aI\\-AKEacQbB4Qf]=U6>1]OZ1BWEcO.WbDcg
):gI1fM/+NZF&\2<LFD)_N,Z17I2;U7P6c)eK[e(;H9A&97K,X,ZWQ3K+<U0O3R:
.BFU7A>T9W;Uf<MR?d-IE?(@>)].e=SOdRg\&/-A>WH:AOS3)Z>Z)PagA-M)<VU=
bZ[X_[e+#@GX7YZ=fZQ44I#OS:_J83]8_(AJLJM?8BgZ0a7Va#)FA)&eIJO;gF&O
&5&-:>dV28#42eg\\e#T-?/85-g0LX,?[_(7E\P?2?Z#Z-S^M^cWcJFG,UR][#KN
9\d6BgbOJ(+QR2^183e7NIfA;O2H2MY])#/<(-1:Z:_NK1E@V0,AY:#IHO15V(26
RFf7<+_&Q&JAVU#K\\0fICXZ)7cW><bA^FWR2g9;W\5QJ0ZVL.IRF=bERJY+WLf6
2JQ67bG_L[g>,BDF5,d;6WIg;=@QS>dJR0+;,a1[[Jd1.6;)AIA7?&YD8G]\;#EV
@GVA1,&)FX@>W=c[D5..2.)9EQ[QAHa2A[I9,]><MTN(?Q3-aKK;FS8b(2g[9g=A
6FU=65JM:8EcLYOUQ;E.S5d\bEOR-9:7P.<\TDT^+JKP<dTBafOP[?#e:-6D>M>.
PUO.S8F4Y8-ZI@IM_ag_d]MI[C([A#[E2V6QdHa\+2_)=&-,e7893O=HfV\^bKf5
U(]Se6c^ZB2.RE-a5SSYGK62T\g2:>0L8H9gETQ\D0HXBO2K9<bYOJ[g5D^4UY?)
aY\4fJ2dC5aF8]RR=<&[7+F0&,#7eJL8N2dbHBM>SD(4AXW[>Y3aO<-3?M?.-+<9
VZA=,#F]f9Vf;9HgdPISI>;;+;LAN/6Q[HQ8X8U\]fZ<4;<_g>Og@/H/P7\UgA9X
R_1(RV6CeBJ,S<?TdY>&W>OXf(W?TQD65fY:KG@)ZX4b26YcDJ4+4/b-8bYH^WZJ
3?7AE,]MRGJX9AfWJP],B7bXPA2Z\C7ZJXZ.cH)1cYA91I6K9YW00G0cb&>KdNBK
P,.-I:EOD/G\[VONH5K4d-/AG-6fI(++2.48WeE=S0@#Y#3#+W7_[8b^X5K1NL]d
WfGP&cLAAY:]O8:b8^24;+_.-QF>K&5J/XF]X&06Q2[#<7MKHDg2ZW:ZBYG.fHXQ
5fQI-DUdKY@X4)-8ZbNEASR:e/#0KVOWP2C9daK6,g5<P^/_6_.I5\Y_WMRDeZC+
gV?<[?J1DB=QY(+,cJg/&?W#_RA:_L6\<X[;(]fX[X;EO^H1-IT8\6E1Z/0E7?O;
E_12)-fRH.+&68/We0FI=RTRA)dZ##VgGCNODDRIFe?@4_MX^VBM4<I6gK2<EK)L
4LN\DAIX\@.FSO8\_30&g&e18EJ72Ed>I,W.PTC4G_d_Z7M@Y,HT^JHSf4V:&/S0
JYdLd=^X_F417R>UVF[E;Df8MVF]WG9AOdV/I>EM,CQ@[La.>B>UBJ6I>eg0Gc49
@6+RLQ1M+0(<T235:ce?K?J.VW#T.<IK=S74-XM3]#78e^>8V+2JWaIcES)VZR)]
2U1MTH4@a:\g0LG18A3[H0[f#T\#?g<+:_3>B?.HHSB#L8,M/^LNVa-T@0F51479
&1DaV+GETKPI3MPd@BR2EG)CMJ4VXcP?1CVY#JDOWMaIbOc[g)44])IHb(b((L[F
N18V/>cD,Q?#d:8GK#J_Mc(^e^,6CSFU9]Z1HM<gWX+]bYZ6M+>B2d9EOgDF.89O
BELU^3MQ;H:0a\L]7)IZ[G]1T(IPX-g)IdB2#;/+a:,NaLZd6G-[=gS\_/IT>5FH
MbFJXS62-TZ+D(#_dVC_Z?SE>51H/dU7?006-/63aebG3]3cXM\+H@VCKE^,>EJD
H/fce@#Jf;)@FVVC2>QPF,35K?EMObKJG:D)UH_Icd68g@g[9Z8+BSF>.G4YNR)A
2[R-H)cYaVG03/d_OH5Zb9cR:^8HW4H=,.(cgCSS/TRV1OTI1a+6A[AU;KT1>WQ<
VG^<5C)XO[1>RWNa/)\1AT<;6M8Zg^FSfg0R&)-+ED()ARK^)7@)OF(@gA;;Eb?-
V<RaE/H1&=;8I[>E0GV&JNf+I=AQA?0Ja69.-)1:2g)ER;]#P9TW+3M8-Q\L-4,_
dQ-C4DL]1Y7_15C08:0N-)gP@eE1_X>++C0fS0LJX<a=f&Be--7K(I.d^5E,@76R
(:.c)UN:\0b/L:dE)_f6K&CDI6F-N1BeFb316..^^[71c)4R32_5>QS=)6(HQ.eE
gM?,Zf=UDGDfTUZN[A>==R)FY.M@P8JJVCg7=@)M-7d=7^-]HY7MaaU5Z]BVW9AL
3WDA4TVgZcLcAW)afU<J81M0LAD5F>f.]ZY^)^UW^#VN&WeV(eZ^DC>9#5T.-^,4
9?IW;UZV:4&<M8=OXMI9bTgHee--;6;7(]##,SYVg45GaS8?DA[b]XAHO-1Q]P\g
b)@U_U5M+T.V/EabZgSJXDdCO=EGcSNgGaD]2aX/GJO/8Pd#_0bYNe&._]aXILed
G(>faLXX5-&bf@F0UO5YYD2-QTTf4eOgg[SQDV?a;__FHd:>RA.eKY?W&cb<#QI^
\#_3XAXZ@?I#N1U=2[d=84a@ZN@0[\EB^G+FG#XAF5:Gb<(2dHU5_TI?eaGg7aCV
\3MW27[N/7cXTPdJeI]RNF#@)YcWS7A]&F=5?\(5RV/,@=fWT<B-/CBR>/H7c<@F
LNa2R89G3,>A#c<ea7^H+6Y7E+e-JEA&>Wd07G73&CG+B?Z6S_HUF-FPD8HJU7(e
SQ.<;MGA:<CH@(&MPc9S@G2YFFL@T\]+:9I97-/=T]8PFD\S?dF,NQEFMXM,2(?V
:9#f3Mb[f9L(b1Y:[Qe/>S;6871cPfHTK[V+d04:+c[#Q/K.3)b?(Z1;A5.7&;YB
VVT\/27+-1+A6fdQKfGHUQ.DZE.g2C(WN#VV7(@EJ/Z3R2G4+;O)IEF>W-/A>eCf
]cILdA_:D:>Z<fS/MYYYI=\Q^-J/MP10;_L)S4B1-S-01K@\7^^_DQ@Fb#d)(NF;
4E3(cDLS0T51[?W3UI7Nd.e.Y=3a)[WeNTE;a#02HCKRNN6-AW&WK/24.4\1@G-P
0a00GRZd(dBIdAS2LU-<V=Ef@L4:M<[&BGZ_GHB#J\&:#FFTcTQO+Aa<7ND0][EC
Q1?W/:7@?bT3e:gOG^Dd)27\)4:]]I=/<4?Ha<<S+D,R)dBXdW^I+KNQ>MD,1(^-
0+:XS@]:Y8KCKEc:dM#;14)./PbMVL-3L]TAaZ0Ec@a+fI?Y95D1dY<(-W;4e>1f
TXP<V(IS(EaeRgE(d+Cd6_J;fg]Q_eSHEM4.[^YfID)cRZ6PKZG<DN[62)c5c+8&
@c_LDBgL\2;)4LGHDPIaHQFAS>X-U:aaYDP+K.;ORF>/aQV,<aRMc-N1M@QUJ9L:
(CE>WbK;/L:/AJ<<H9<@_&3/;(8cd2:G/X5HL<(JN@E+>b##^@X6CIZ4_Ne5<fd_
9X-Z2YZ(^bC3->UKXCI1-<_QY+=Y)FAf]4Pb[N<>?H=MLV7DUR.;EKIW83SQB2NH
\-M>c._[4?@&@>c9V>4TFOHCYeF799AJAg/]MU+P989f>]c>?D(ZWH;+AC[(^-+[
Xg00]RSEPIL\7,\U3#6YSDX3]Q(XOTCc@W.[]M,<^JcKK;T7e-:G+_Qa0A_+4Yb6
P=Vf]UaaW+]>P].J(U-:4I2dTF-Oe36=@W,aRJ-WY]_DG;C#f9Y,+;EI\\R\N1@e
QO9Z[_LZdAe=W9X_P+_PR=6.:-;M563T\WQ\9821RC.:G64f)B=D,+TUa;KG/bff
P/&_,>NKM5BN;W\3VJVgOYN^M)_F&CN6FXLM[AU\O@dZ:_=cU3Ug:.>+3[a1fL^g
+9[/AYLObaGRc_=#FO#>IAE#c73-)5LPQ5T,CNAY.01W\5OD16VA4Ic?ZBfB&S05
GY]@]d6T_&<T)7B<Y1//gf)W3W>6F@8Ga8;/TXIK.U5N9.7e]4BKOFfU5)1P6Q,T
9+#cS-L#IYLB/;ZQ-[4&\3=]JJR5BWDg=V]ES@(#5OG]eS;:VGcN31&QOg&a97Af
9g_DJ9Y(;HfPOC5R+7MA?KM26gV>AG#HK-c-aO/gIFFdW>MZ@E.g0?9Y6+aTHP-8
#4?4G&[H]7^b7Z]^[I-+TMBX(FWb8c>IV97-1EgF&C@cSDLa>6?#XJIQ/;9ZZA\M
5MTLg>:^4Y4.EYdW.b>+bD+cO_[F8ag461-;JP70F/OFcR,<NTM6UO>OEWB:N=Ze
+N:/JM_g@ZO]8N[<gAdJODOeB/3TXgMIb.S3E4UAGHSd>L5.3=@B/.BFQGd07gZ1
->Hg4;.>&@c135bNI]X;O2HdG-O/cFa7RDe)6(d:@g-fg&HZBZ2U#KD>bYI6J#Le
&LCX6ROEHF/#AQaTDZ892^@]+_a.:eNF@1LE8[Q6YD,QPK:[(:5KETZQ;Vg1\O1@
>DULW=8.If#4:R7Bc2Y_IWHdFeNY_ZG)L:9ZX5W;;;1AME77M09>X5Y+K5R1,[JI
^J9a/?;b=a4P@WH.(O,SEY-YLc#Yf/3;@3QPAAO;_\_5H.7g?>O>IBG6O>F7_3>b
=;gKI\O4cA)7CaS;YacIT:FdK0VT]@aNJ;G2YVaVNA6@6(+QY/6+PSKO]b[TQ(Ld
g6I>1ENT=BGMcfd;Lcb/fC=GY?6K_Z>Q4P6U(VO[(3MRJ7XE(>,I/eB=.HF@a55G
M?;A7aS[d(ZI+7.6.Xg[A0^=fb6EYgP4F[_gg&2g.:HN:HA^8+F\cBN-b8>I]2SP
XSWA&6Q0E\,[;Y;@S)VQJHKe>8X+XbcP61J7BdEe(X^?PV(_;ZE&Og3]9D^ZD.6c
+J0d=>\>8QXVCI;>AC\J<B2_K4+P5S](X+Nc#/_&[0FbSNXeJDXW(QRJXYBB1Q:U
,NJKECV,<Q>)Rbf\DJPd>O4\-&9PXeF:>JXBQT.+];//W/I)]&ON:&Cca,FG)IB(
a3L7_UN/+3[-2EcV&aP-[GP]Pf6J?=M0M;Bd,GM=/FU#D0PI2[V(7_=F(2??:2b2
2B[SC?c>4,#@/gJ=MV?70/M[[MQA^X+)bbfH>8d1+MI1O,+X5\2J9D&9O]C8P2C)
#@[eC17;^U^E+LScZN60YYg]L?.7YOe\AYF<a#([6BO\4.Rf^.BFIa8Yb=&)?PVL
/:VQ5_:6bF+UGR8U)0+6XHc+=bGUI:22\8g3O;@RE2E>R&f3;,D&-<D\PQI3L\H@
+84CYQEP;N5AR+=K+-dU+X<42>Z-b3RPf\c6KTM=f-:BONBO1F^cU-I1Q9][SYYa
.HbE8HL906e^X8JUP&ZE&Ub5R&;)K,GFVBd1Pe7O^Q/BYe;]e86O,^Ia9a^V-?=^
,@U=>/b0[.D5FNF].+D4BUdPHDgB1I4TeJXc9W#e8S/<ZGYQ6)9<@(TVT?,3DfKH
XH-R,8.\5Z#D(B2@^_P#-I\-CG]g[NHa()=&K4=/e4\S=6DERaGFOK]DQWa:@\FK
;4N[FAd&Q_@&5)\NV;BO.6]Ee[.fCf?B^O]c;?;dH01062b@a5(W=&X##?eTH^ED
B8\((9OCe9=Le?R\D#B_;<7W_K:((?NMFLbRNcR+=dW?)b.D;G),[7ZDd6\I]W0d
B&Ka0M=cf9ILWMRG_[S0aT=gMI-;T0S)c,SR+6,9eZ@Je=&BWRf/+OXCBO+Xgg9]
84#@ZAL0RGQDe])Dg[L_D>eL)?I6B62\Z9S42]#PF1gD87T@8#)=UdUKB?9gGE1R
A07L5HJRZ;D7;JeB/XN0573P+SP08]=O3eg0?]F]77QU.bc^>EZ_3dV#04VFGVEe
ZGQ0c#&E6H1+O,OL_0AY#1,,eRC?SFSdHWG2<8BI=YGe=O+NCM5W(6&M<;FLa\9]
>T#\g?;F,[ZcDeXR70#B1^(8OQ\5[/Sgf@;\?5A9OJOGJdgS1I_Z1XS651gPX9Zd
24XI1?8>C2#(^@/a0CDZ]A?,J:X:ONO>M1G<WN?Y;#;+;PeH^4+_AESRa6B?f/J_
E<K?cL\-0\A8#5LdF>Ke(UO[5LD\TfI[]4<O<6AY=#)#/[/?Jb)CMSXEJD4B2)_U
?PWUJg-Zg?M__T2Z<[K(-XS^VfVM&O=(]]@eU[a.EeH@MHNGJ52R3Q,gVM(EIN;1
@,bC9gAP.3<W&FKec_C29d>@;gTFbA)Z5RF>P[4f.[+IP+-6?dB=3(.C[#1PPNV+
IHK3d1+cBPN2c[])Z7;#>9C]E8dRW<PZ;E3B&C&.@@2#45VD:00#eU682^N532c0
;E4-K=_NAdQNHODQfbNL:d\,NFNDA0N#,:H_C]]QFY5T:UeMFC?W)NQ3T1]B=eN.
;/&0\]5LU5g_C>_PHaVO;\NE?)=gZc#&MG=G/@ZQaPY,(2dV0?96RPbNGgDRAed<
]/6)N.bM2gBF(V+.Z>cXFU[&O+[U.++E;-JP1[-M.S<IcB?)]L_<gc9_0S9)\E+5
bA;c/6GLGVRe[A6b/WN@?6C;30dUf\^?F]<SIdL_6eS@9US_FE\Ud(SdUK_H1+6Y
Wba,YDfEHPJHSZMKeJ)\ZHQb&U/;V#./0_>5JCMf3fg&^7\E8[\&8LIJ]cWHO^R<
>/IC?4)>(PH@@a2ICEZ(f9;(2BJ(83HY?7.(]KNY-X0<.R_\_U9(_/dO24+O#Hg2
(b?DCcJ#Q#]?/EIXI4\;K-U.J>LZ++2B:\:OZ5#[eKGYA-Z#)eR29g)W=I&:^,+K
BN@L:BEf&ZMJUd)<(FG6BXD2^]OJ2FHdEM^/UML_0:g@a79MQb+-[&G,:UaZQ8QH
c-5VB(R7MC(09WXC:;>>CX5^#4+;/N?+8ZT)K>WG(Z0AOS+&R@N9LQZ>:B\0ZY7S
d2Z&V\;Ob:9HbgAVJIIGRQFW-#6Y+;ROAOg>O_fdFMJJL188agUQ;:U(YdO16Xe-
ROA3ZO/_AZEVF[CB9/VO65JC/SW\<_40/^?e(L6O9>&FTgJ)beO2H;-CW>[.<7\O
d4I5Fg_0PU2=Re1F#P-SMA0>1T2<;.8Ac5?;B)U9@B2]d??XWbc)UP8@./S<,@)D
c=:;(?Ae,g#H9CX55ce20b4MUO0[YCJ89bP/W07<E]P65C(DW@A7#L75a^D)75E#
]U._?8CM;<IF3TbA;c0&E_OR7fLF2WNW>:F.U7X@L2?a;W4@c61YLJdaTZI11AAf
=5NDL+fVG,U8V.&eVADd#VA9TFMN5JVO#[,b;229E<V/4N0TGNbCD7Ef^/4(HK@.
MR+7)(MT<[b,W4S\U/PW4gW[K1&cHeeRf-^F:./QFS^7Yg\\KC>e(&dXG5&=]JS,
)U&D/WMc[Z-=PEg]bQJ&A:OOf:cB6M3LX&_6Lf&L<Pa1^#/eWF+2M>XgNBWGB8_Z
/]TQOH85I;0&T<L.bE[gHJ#HB+J4E#7eBIOD&+fZ]H8&aV[)QeBU8S^LNH5cGg+)
75G]R^H]5@<HWK&F3=N\FSPb2L?0JF@(]<KR/VNbEA@5B_+GL^E<6__5^N.SaIW:
Qe=-,J1Hc>_4U_;J[5CC?-dJ9W[]H8gZ]\;B1>3OR0b?KX7^IgPZK1Ue_4_Y:Sd_
J9\R0G5?eI\DIH;X_RI33Z2-V.b6.>2[Sg0_X(E[(56<f2O66EF?1BXH4ZH>JQF0
5T+^faI&He>aU?N(CVT@3]6+c_,,N7Wde7e5aNeBRgYa>0FXcP+bP##&d&AOZ_J2
#FU=Og3>QM2_-0DIC,9K\PF,\T1_Q.7_T=328,I2(@Uf]YXd95J\Xe0RR6T0#@KJ
.LJVF5K1037eG6M^GNb<-;?J:b6Q5G-ff/@+##[b;eGc=Z2@.?/[?LKeaB[b9fZQ
E>ANP:H?4(NJ9P<B+cDPIgLBcM;5)30P,9ZgIS#A:>HN>;M9=2OW;K-c<,+;#JO>
(-F3M^V1b0Kg])4<E.L>5X5>XNOQOeb.\IE-J3TC/VDceb[e>4,C(MH0^6.fPCc0
=aZQP0bdd;3(B+_QfCbGbOaKI0I-S+baH>AQ92R2N.G-7KDU_WbNFLQ;\+31J^7J
LU^Pda)bg<,?TLaUE&g.YK?087I9B=5I,Wg(JRE4ONVd()N=NOOTN?-7UDf3.B>2
@XV1]6:QTG+PO_52?#.FT(5MJ;<-d:bDRY<;&c#DR?VVa_4Sb.<0&AdJ:a/@^3PY
5W>Y2_5<0Jeg>(b&d#\Cg0R84/-2&O5Q=Z89&7N.gC=[I6WT#=?)#=8)DBLXGBNX
0XS&8X5#b3N0a+)KDRULc:OC&\J[ca9O1J:?MaM&&aX&L8gZX_(8T/U6EYO07<N?
A:=P[&fd\^6#[-C]>=+7LIUd5:<M9)YWYMAKCM_/P59O<7=B(g\@H>ZT6N2Z56.T
9B[M]0RC.;c7W@?aLYY_AUIG5[Z2IL&Na;@^;J47>SOGgEU9_T&H^RW/:F@X2806
)R;DL9<C-:,:OA.NHXUeT]9E:6H@RM.Ca]M=23fF:Cg.P-IO:LR:/XF)\#EcY^@O
PcN<CRH5^V_+Q#P,D]2&Rd-2IaP0OO,5]MQQZB]5d>C7J<.IAPX9X@O8J7^1.&;O
N-Q39L<^7:BQa8K@.NDQ>]7,T9CQJ=W(#0J(WdL>O6D<]f@T;?<JE+eSJPX50VQL
9;_..H(g2R^NL##)[RJ9:3<N/<1T.C55TZ9g\0J-/O9+NAV9)JTQJZ@U=F.?9YWL
<>]NOR_bI#Z,)QK7+TEIc&OW&;P]A[SUO(aEc]YUNMbYM:5aeZA[LDF>BAP__a6,
RJ#<bfM/VE=\9KW>fCAN9:c]4=DLTc9cG)/\4+gWK7daE^>Bf&XP=V8:;0/QZ7YM
2dV\CFb&4:Z)<g[ScJI6VY.E)^Fbb1bbf<+^ebG=-FB)bH/J,/EYb50T&MdIaAZ#
;A>,;BC,#4FSPIgQ[[6?EKKP7.NN,a65ZM8^^Hfe+LA=E_9VT0.M=W5AFNgE^08V
-RSM=Y8+Q^18;a+cY1/V@:-)2U+;D7NUY;,^O.57#Pf968Y;:9(_L_W_:8_S7;PI
UD^KRY)P#(QTMM9A?cN6dAO<)UQfR0H]FZD:/OI3V)7a<cR3)F&ZS\d7BR;72gE@
d_538N1R<[?g_Kfe\^:MD(d6XXM9R1ERCZMXM#@5XD&W7J69IH8HS]5f[Mc4HL=&
,<[;04/a(Cc56S>I\)7MQ]I/BYXOQKO\X_#SKa+XTCB=dB>4A7=d<LJ44A5ECNS2
\,7#@+CA(Q0V[b5=DSdY/KJHC^Fb4O:f7Y85G4??VORM\@Bg.Z\de++CJ22BDYB)
Y@9<KVFM3N#cCMd^>;(?EECRH8=\O<Ib&g5=MBd/<KVH2a_:D5]_WZ,gUV8[8dQ,
f5OJ7)d:OPHb.47:HF-e1(3[;>@;A/Se&c&E<1Q;a^;?,Qd+<DbH87MRFDH)4.J9
IQJWRI?TR5Mg@9/6V&/>5F:\:DQfKAS_6c0(7F4SPN1R7ZD^PS;:WbO_B=/fWCWb
Pg<-KU2YDM?.3DcR[D<HS19IGdXAbU2N,3P5@U/W<?f4B+NL&aV]9^XQFS+B;aI)
MV^ZO:=T@ZXR2ga39/P@\\/a><RVV+3\-b#I0<._YQC]OBX]3#Ib#LU51gP;.dEI
_I5:X6.0A+#PQRHKDY-FSI^O@;7EMc3F43GV:9R1WMR0^Fe-JKA?)6+-C13?9.Z9
10RZJJL:BHfN;=Md&3[:12[d<2<#A/EDA(9:2?XBe[Eg<V,W9c#2Y\<JJ=MC<M\/
I8<g]Q.)3BF5N_bSH7+YI\+TA5^Z&GbO99EVGGF7&:>LBY5aU5KGE>?dc7X)?3RG
E>.0&fTWHBY#P4>_a4A4LI?K;0<geCZ9YC.8][VaQbL,5eU#MdFJ>8,eLH<./Ld4
YEN4C>27Y9/A0g@]O#<--Q#gAG\\Wc,eALLFB(]4Y2<034-LYQ52K+/.S5Ze_Yfa
,7R)RdM0<(&QU5HKJTTf.)ZPD,[_/Fg0e22FPOVX?WR:;SK#E5<3H-8L3):SfdaG
W=]>=7\/O,d=1E-K-<Z4U=-D&(^gdFbWb([>/e79VRN4ScS4&8:7+(<T9b=dc^/V
DBI6a4G<MR75.cg\GYCJX2A4VTD9P)0(.gM6+3IY[Ee=Zd=abQQ+=-H?<ZQ3f@?4
<g+<P]dKDEbIWKg-PX04(5CW_#P-8CgE-1)RS0/)X2JA^-Q/<Y;1#<\&]-<gI??P
cLPA5GV:<GF21WV2CC1Y/JNB)-V&O=<#()UT2S(M\[f@AZIGG:9Effa8QKU8D&eL
T5L[QEebU<;fBQ9@QJeA>Ygc+OG<[-g++eWE.#J2)PO#^/XdF,9gSQYG08+0.6LQ
6&U(gZZ67\b]Qc3DRS8Rfc)X.J(Y?;H)Ya(OMA81&4PTXSPWJ@)193++.:)Cbe(N
UX,<2KYZRL(0;+Ia.fKAW@](EY/dI=Z5[&(V?]ZL4BWN7Y]&=-:;;;PEf61BW]c#
]U^XW(4b4Tf)@Q1H_A2]2;]H-0#)BMAI&g^5=Wab0L]EcGUeS+UP#_94+F2X#Dcb
EHg:&R)1188C?-cL\F2UJC@5X4?]H[QVQR+dBQ8S\IW&P#c8a)g7bRI;MaW/Ndd@
LCX@:_7CAc?JdeIJL,)79g2dMWSB1eQRXdW)>0(44UCG\@GX(\WfeSe/7aJWZaCH
bL#ddb..\JQ.fKfg-F)f=R2?@@^V0GJM)8A>W5C+ESCRAb<C^437#Q^E)[N9AQ5Y
=#[FDV#WKb(ZEK_bF-ZM^:L=RGHBMfDe.K>Q(X;7ZX8UHPbX<>8WU=f&&:cR:9;/
/XC.^?H-H._+a[]g;CLCYLD)&MH5NLI@3>0)P>cP[9F@:BA&F]DS]N2FCK0Hcb9G
b5IWfX(4+;YK76K2(7ga./K@CWY;E7B07(,_<6eML=+[e6a?&]2LHM^+?+Y#H8#?
_X#<#XgQa+HLUPg#P<,313>)5M8e9^Y(?=\;H8RE;^#F<,ZfZ^B0B1-:c@U=L67H
)83_LODDeH+92T]^>50(:B<JcO?cCDHNU3EL7\D)/K>X:4d#d1\1R>GOd#HJDaY7
^S4f^AYFH3WZeSeAPgR=3Z8=62c,_8(V(,D0<H=XbP=</35>9/WgA/8U:ce#W/D/
;INEZGKKRW@+A8SdWZ(g.[@N.d;WU+aE_4dOAYCg01\GP0WLcM^RAN-N]bT13C5#
=40>40;:Bc/&cKLf0aWG^1FE<@;_/M?2.EV6/\5ESg)-PD(L,1AYA1PQ5Sd+7L4^
)HJMTc/G?7f1Je06)fYG0NaZ4MN.UKI.)&2.Y2QL63E9(KKQT-?7U:f_2]/+BIf@
NZBM6bO:AWS,J44B5F6W+P84MXXggQF+eS2P#2=FF(ACPFDX^GH8=R(.3bOTZTe>
4H_RSAfSH@4:U;d,;F/#-BO)@H<KI][Q_BEW+756)GT,:<[.5:8d<:.KF,N/bLWA
)VJ@T&VNTfU<.dD3UF5O-.HJ3RJEf#00>3(##Q7X005:.fBG8Y46D6XNGHBL76VU
W:EP@c,>.>&Ra<F>31RXYZ^@A@4QeS1UL50)I<^MS[L,>IU#dC;(0I.EJU;#])40
_5XPAUT2C@88&&[&,;bGH[JR^b,B;+T>Ob&R\,V--/EH/:gIT;=PM_,Ld>174J?L
Z-/PAfN-aU@Cc>[&WA5Q3f\EREVdadcCHD/G6Q-VgOd5gEF;^WIVfXC]T^.W73+,
)N\T4I.9O]5<OYe;+<#Y)SW:aR8bgVPR\9<E/TVP4-@fc7;W^00GB5H:W_HSAd6g
GY&=L14+]NS[g@:Y@\ZW/@d1&>\5H(b6Te^EK<5-2->D+0<g31=aQdb]:&LK4e87
D(a/G-Q&ZQ?dGO)5QV/WPZd>7EefS,#282C;=R0&9ZW4#aTEEY=(,e=ZY\J-WcVg
fLN@2Ga;Z#)+e9a+D,e_534RJZ&I#.V4_UMa3>](8I5+AEUd>IS]X3&15])._-EY
540V96P@R)fM98</.f[-B1?+@KQ13A;Vb=?Xa?FDO)Y/QOOB=:Yg/-aC.1I\[+c?
U;8;65O=CE)YP1I6K0N<\NW#_>d]:6MDG-C<[(TJf><ICS]PGfQ,6)Q7+WY\RLH3
XgQ72;fGT91.)Ge&gH0STA5.B@g9MN);\MA,+.MJZKB8FgYA:<<AbNDHfgBQ01bV
\;#[F=:ga82GbH^JQ0\R:I)J6,eU8YIZ72ea&0PY2\_e<g@&D-@JJUf=+\G\e4EG
+_PQTbV3U<0Rg9bLWgS3RJZ1>.<CIYTcX>_e9(4)b,JK\4\ZL_IYLPcG4Geg7fL(
;=?2;U=&Q,.0L-FdXg>dYM#AIbAa2Y[L#X9AV\Jce\,VL+Dd=CJX3D97,d4^XU>c
9T2^UUcW35@f9LYCU^L97dW8F^Sg4.^K(OV[KGS(UR_MIEg4+&@b+S_77eRD>dTL
B@IXBU0;5TeGHMLgeX:GB4M/[42]JBUD,&OURS5/L?H1.\ObQ;2\U.<:fG5B&c13
fd>CTAIdZ)?d_R\NF=:X;8G9GEg#,RST&)gJJC8]9/(K<((]XD1NL1f)bAb?eUV&
Q<7#R_6b<\JG2@),@-?48.;-.;E:5570M3@KeYDaAJ]MH10.\FCHGbJR,<+c[+4O
F0^.4S=f6]N]1FbSG2-66GZLXO0D/[.@M]-MHF#c8F,Z2/H=dHTVJ=3E];\B<bN/
I0[[52C5IEP@6N7DO2H_YET.3.468L8>#/M,6A0PJ:Q5Y813P+@2_6H-C)8=:DZ9
ReE=?TU,]+0970W0F]XDS1ALYL>Pc7^MJ9K&K\PP2bU[1#H3P==9([(:&):LeSE-
3P<.c/H=++8[K2OL+^&6-G5@ag4,Y#FB]QEe(X;7-T)\MQQW]:DW4e2&b_/d3BP5
3TIKRLD^)[.Q:W9YcIEWOTB@8?Q_A:S0DeXK#^0@/MZ#:EVE^6QP2JR5NR(e/3/P
-f@K^+c^F+GD)bTTEXJM;B1=;V;BF5fKD^eFXa]IWQd7a,4EC>Pc[^^IK;IE=57^
&>SD@D+&:2IYY_FZN)MeIR9ZS(_6(c0Q;:N@aD];O>\>ST?B<UGeDH>H,[HV6=O/
.>&2+3=M@d]AF&W</d(#X/INXd(V[b43Y+3E7D8>dW(9E=-,e,f=XWF(X4YY15(D
/&Kb=FG\[eJ]eH,P+8d/[?.9OcH:3-<#3[VQ>[A:ZYeX>8X6X,V0dFL1BPcN3Gc2
gO,gW>3)H]GCXZO1:CCKAG[5RG\g6S,B4NE]U820?cM)aA#R,Y9;VO)^99^8MDe6
W?@Uc70/c<3XXPMKCdC?g(AA-f+@04O,A1+0,K[Ibe2@<cNJ+U&(V>I]+;+K5:RO
XG60MN4J5WR-=(fOaae+66:Hb?8e,MWW0_(01O5JPgAH3]U-Ea4::&\2c8:g0IGZ
S&T3P.H;KT_N[5H^DFF(e:aZV,b#6@&abGc?AWFF:QfU7D6K3PB-7a97MWB-+a3W
_M>c@/7?Kc@,X.^2QSf=..S+bU+&)XBUS_9F>1?U^&_9DOAL/YY62;,()&3(]baU
b,FF=b+]8^78IXMd@[O;YC6=V?+&&+NNA>)BY/]TafR7;SN#9-/3;LH1a\V/JQ7S
?+Y>Q4XK9M4WTNMBBV&Ad]V3fEf/N)V_PZ67H^dJII]J@gN1=d#1AN_H]f^)E??S
,c(_S:C8T.dEVIGAM7E^Q=1dE8GYUf247EU56+aVUgY=NE>GgH9O)7F0QfJ13=0(
D1L7]=D0g)8E.V.@N(&9P\fK2;E-1>V11]1EZ1c&G7:WXKObdATb\G+=[3<V-SJ?
UWQ6VD)@ED^^KdT_6T34Q[PcPc?]S=>MeYSag)1a?]+:@9\fbDSHB7.:g@4fHI,8
1ZO>B(Z<ISH-[?LA_;L.3.&gOM7a(<3A>T1-4=]13NfEL\2Bb)[DK&G=S4@Qc(9[
3)Z9I&U:>8IfKaBLL[GJX2Ag(V.2:8+E^OW<=GY3Pb3VZO;BX//WEc0If\\ea=d<
_S9[618QH;P#8M_=cbFL>?[X^KcP\KU-.7HF@gcY32O\Dfdc1ZL&=^SK8X]5c9AA
(C+0Ee,@6g0aZEF;VbM9BQ>bXOJF)g<ZE6G=O,L7@ZX_3++P<fJ&>,/^_eH,(H,#
\[gb2P:SL?DBR1,^]GH:7K:-:FfJF,e:==(:DV[6NP,@eJ;Z2O_-g=baAU8F8#F>
QB4)17K#:]/efP86UDU&aWI:PB5aF#UF0RGQ7BJNT<^05PV,&)=RYO<V)Oc1=9ZM
WXQIe9>>62>/SDHe3eVK=OLV[MY:@f:6@b4<Z:A.=E1,B.CG([A0[5&O>)cf#9Y]
d8g^Tbgb=A,FgcQ]#FGM&1(\c/VU-^5N=bKG#e=4bUZI4Y&]WfVL1>b])0LXIZL_
=JP.AGfeg/fS]K\J#d=]g./e&;+ER+@A9[P6?;;:TK0O>V-0f4.[N0]X>GQ^X_fF
J]c6PbL2-3AbS?Q@(J]9#OAF)&_XN5A7;AS)--B.S(Z>J[1X88\2.ZQgA@@dI.+e
2JN,F[1d?e\<ZM6Z.54])/,6MQ2Rc><N<V_b+K-&a+6AK-<=Te-0VK)L=Rg/J>NO
;>b4M5ES@JKX7FKc>\I:S(deH2IYBMW0SPC-@\)X2SJ2e<Cc6NPD<G-)E?G>=H1c
J:4gJSG#E36KG):T6K4QQ0_YRYI5&^LD#-T4W?X4D,U?)?4XaOd_HZ^#TOMQ]XM^
9=66<@dB>OJ68_LeU,L/3g(#:9+WN8YD]SU[E=WdXDB)#/GWI^DR<+5R(FBD0_WX
;)B9D:&X2,UaHETO-?HKM2@R\5VCH#B4?\bCD;.a2d/U(8@EU\)8WC-LW]gd?e0+
b;_>988356&.3_^W?F8T/C)U+GLaHZD=g<7I_).I^YW><.IK]FPSA+65>ZX1\PML
<)&]^;PYJJRVN?7:HK31;JDWHA#JEd,SB4A(4+eC;aNd1+dM1.e^3O=ZIHA+9PM:
;JGbbDDNGEda36M3LUe>.=KC3P0:+f7H565W7S)WW:3,^5RQZG8adB@H::;W1J@c
)e<4^)TH];/_3.WR=KR/KC&.aIEN&Z-?1PA/dL<>VXU]WJEb@cV,(WJ#dHX]>77^
M[(TGCMT3=J-82?=7681C)@2]9:C=7NeU)[W49a0(I4e-KZd;G6][DN@&H)bg=NV
6=\b\VS7+cJgBWW:&<B(;EdI9E1C7Gcf_D,#0IdHOQ15,eK0BHHF=BP<#F[eW?OH
?JMK_RFQQ+Y@Od4A2)GD:)Y-,E>[0S-R;\gBcWSNK?)0P4AfSMNB1QT&CA:U<b.F
a=6,3YB-BO_B7=5T:e<(<QPE,QWFI8.>36FTIUfX-0\D]TYXEAFB2PdDSAdN6&..
gX&fU6:KLdBab1L:\>HV;M-P9L=8PDbND=/#0N2);]E6TRU9,(F7DE;.FZD;R]NY
-W2T=-Kda3@g9][@)/1Rgfc@J6_(IXVa[4_0;Fa4V@_8ZLX7/98]aH]FE66[cDAb
+;4:R[Z]2<K=+Kf6.F7TW6DPDBF)@7_OA[5@UAeUB.MVR=Q;8J(6FG(S<+a=(+ZY
D#H)EZ3UQ.65Ye>-C/_)5edPH@,Je8E+0&_^7+^B&[^@RFF9GaJZQVLG[#>T^<g4
;9SA#T0gAd_OTe[(/D9&Ba?3B74b,/_O^8ac,\)J\Z+2OO?YV3C=[4&<aM7#Rb?g
_G^T+Vb)Ic.c?RP6/QZ+A4-J9[/A4Kf@3KD.J.A(EN^a<:1[1YR+/9N<&<YUa2dK
)2WI9aVdc.]#3-;OILR)C]>IHJH@gXWQa;7gMa\D/-WRW8c,=#901CcTgN2U;T=6
T=RT#_Q;/AGTc;L@a]&?RT_RWG2X8K]\86/gY?e9)\=KR0V]J_Y#^N0\@-AB[c#K
N,>;V-V4Rd24)<f@VJdOFOg_ePfN9:NCO7Pag2_?W98CR4^bOf5<QcBgCS8(EP/S
NDZ[ZRZGD:6,UO=XY<&1,ODH-Q.5QgV[<-+PU8E4-g<UbGfCA7XSD89M0b:_N.0?
7VUU.+\e?4<@Ta932WD_@#S6@6:e[;>9MT=^5_XfCVcJ\ZBb/OaG6&b98C7<)F45
6)26RQ(cRRG80P-c\9YbDLZKWMLS,&<\/UG2V[_1HH:8bcA]84g\OHd<WWLb2==7
QJHU6\adN^V<7=Y_C0fE@D:QgUb2A,D\=]PO9F.O#6M#QS<(g&Va\GSJX_]H+:T#
[MAET:]Z^(2GA4G]0&JY3YSZN0KXNeMKQHNNC;T@S2cd^aOe1TFQ^_M@bXS_J7KO
2+VbSWRXOOI&.9^K@2N:SedL3Q0_OO8YdEI71P-B2S(WNH=:Nc5052PFd9TF7E-U
XDTGKIQ1(XcIaUJU[#9P]VZ-C/:;)=KJNG-Rac>cC?.3V9DFdYg2RSgYXcYLU,MY
N1=MF6-&+be-H0KWH6=>67L0BY2QJ2b:dUC5Q^c\>3ECYgIb+.,#;=<,7??Y:55B
5&_M&FD(ING#(8QZ_AN^V)G&()BI@\Z2J3N8>8E?VSS=\PeX5II&3F^)b8L#T]Mb
\I>T8<&A._YUDfY>O7g:f<6S])UU=6FC3ZVL:3FR6IVKUH9-#YLI#EL.N&bGgKWI
6LLT\QdO]C0-(.<#2V9=5bZ<F\Wa>g@/]@4a8=^O8a-.[?B9YE;Ig2OMRY,Z__,/
Pg30/R8UD7C8aJ_C[MaW^5M\O8NM4M.TdK[S2\LUa0RA5YN#@]Sb:CX@^a0^HY,E
#(,=7:5DEZC#5S9#5.cH+MRfN9,^X3>W>>NWSLKNV@21:XBPb#Wa4W<<DD@Y>,\2
4N^^CT3ZNRN68[19RI7?&NQ81Q/#RCE#O&.4DPEYTZY1\,=a[g@\-0.W,#2\8?O\
@;_+B>E(EE)/5Hg)0;MM8R.GT(IbBF&9C)5FLB-5)c):2UHf6K_<_1J8AaY;P-?S
\>.)E]cegJMJ=7ND;L#/]XHV-&A(=5F\TSI]Qc25.EPP+>eLY-Wg/)H>>RcWcJEa
D&(VZ_0POER58U\/bK5f5MfJfS)KD=5[bD8A5#8(9P05e4F&cH]<#U+#>/)gK0UN
,<&24K]-MR4d1Y5B]@+XfYfWEZffH7JA3/6QKOABVFCUZG=]?-OMKf[8<-EBH0BO
HPI/A_5AYKZID.X/fR?O9DJKE\>8Z/g?F9De)^,JY#OQ4_._9)=?X-)>AQE9eW=g
F6#LS:_HT<(X]bG)-3FZM<g;d1_HfI9^.\KZ1B3MM[P#8/Q00e8(>-\=;0<,8OLb
BG(9,<<\/9V-F&3,92HA1?W7O7SC-SKOJVGUY##SbW,V(C=c_)VG2@]77H&[d?cD
9<Y#>#>?4(+9<:@.7@\^HPM-:gFQU/YYN)R<H#7_KEM2QeSa6Y)/eO>)^T7Z0]--
3DegG3EZAa0[_PLUDW+;<c1G_Y;+;)4ES\g(DE@FdA,W^B70O7&=F\X?JKc;E/N3
#@.ADZ)0005<VW4827a:E/cfK7c.L4JE[WL;T^1WN)b(VZ[>,f>3A3fS+Q[#.2;9
IZ@C?g@,1eO&()Qe@-<G-=;@=TL.=C>]bZcVEg1I1Y+>>K4,]O3<(5ZP-H&D&J8#
WRfdBNMPa#47cWdFYX3Rf/Q0#Y&cbc(01TNY#4)eLHE/Pf55<fIb<9&R;;&bJBHO
373>PSGbRJd485]8]YWXMXbTP,b,]/9+O/:K-J?5FgU+X-#3UE-A2d-:,=T62156
&AC6KBWQJB6+6T)L)/RNgC,7B=SWdf5;d4KUM)6(Q4GJOHgb6bd@>+RS?fF&PUf+
Q9&_VJL3VU;D,G9N&PE:F[-1ZQ9SI[Z_#c_OK5BI/NB.,fG0.4R(@RA2X)dIEV[B
/[8,@R9;9RJQKV5b1bS:?>?/NLR?bNM0>-b_O:WKGP6Y=Q>5a[VZPbLKM/34#M&]
E52e:fSaaLbM4,W(Qdd]@aN0C=CL)EMH9XB7E^^6HC)S/V=TYWaULeS5225^c:FF
:+Lb5)dE/@@Q#0L8YHbD+g,(a9&-]TSP;U=,DYD&Q#)->#7:gZcF<c]RKJXHXgaF
TGP6QI1Dgf?58]g5#[8IQC7cDM.^161[fM.FS)bLRPLY0dJ6QA^b&]+8M&V9LIf1
OX=;d\-P75HGd]a,3+/R,gUgY0S^^O[1+4PQO?202=IIaC:HLOge?.2ND=J=T=(N
eW0HgF0EbS)FCC\c6]L_>\FE::b3V2-YTRgK#CYZW;2C1F&INFO9@&Q^=<2f[]R0
5@NK\ZF_g9I.e//?:G]\?b]ea?9-9^O?4Ff;ZAS0Ab,.KJg_a/Ec1Pb3ZWV@/fae
OfF]ZV13-W<G3XAa(7[2>8Fe=eMQ5EH8?@N^[M5I,LEaQX,RF0PM3dYfNKS[UM1O
<S&+40\bNQ,eD#NUf:5]<-<b]C?=6Z,e?W[1G^HdRU99X3#-5Gf#_N1+9ZGK3N>=
VA\P5#2J3-7Y6B_I?=(J0JD3()K+XK2Sf)1JD,G9Ocgb2+LLgLQ6_Pd+X#>5NPO^
FdeZ5)PF<B5HA#FA/1>gT]K9#B]_,<(N-@.SX;?E3UZ4YY//87LOQUF6gFRg][K4
e2d2RD87GUKJ,6+Xb5b?B(BQQEQ>Jf1[@>F83@/)[,@HV[:ITdM/d,X=KA?:_Rc+
C3W2ZJ67Z]K(G?((<D<LdWfNLSA:P0X+TX2_V..6#^WJ(ATPa(7+7TG>XM@0CX=G
#-G2.2@SEEOGFb\5IdE[02V9aGA9G?TG[QJ00?M_&&RUf\G#H6Y<0BVE\>9._+B4
./f88_gYOd:#FTEb+4QHSQ:[C7;@YP/-M0-Q9?_^+,\4ZS7D?H@fPJSTUR3aP)OV
;D.cI35aZZ?#@_DH6Q]Y#2XTZeVbd)g#9E:]2)Nd,3T1B6Dc&4I+SNSDQ&2d&B6B
aeA]6RF7->SP+1c#CgG_/M0MIFMNI;0^IV50dEE.P]1:a?&8BH^]c8Ge0(>TS8;c
=J),8#K-g5e>VQY[MEDKN+1;g5Q&<[5&[^S)E_A0HRg3,=;?(<R7Ce(8,-VGO,<&
)I543?YA:#V.=I:Cf47MIMFFG1C=/PK1@^:+_P:P/>0G&#F94)FFQ@WBfcUC)QKJ
4<>WV6dfR?5_41OW/AdV_J?NQ;Y\&84VEB=YeM9>d@M+L/UV[Rc:B4f(W+L+\I7)
9bN6<YQgY64H5Kc<^+cHe9c.=?f,-d\3f0_A,A@&]c&>gM/\dE6f@RD+YZ\Q2f3E
CX@a(W]/C&D-.CH8&3A,PPM8;Tg)d8CD2Y3Xe(;/@B:+QACDN1#BdTFBK2=.Z;<V
Ueb>Qf/W\OB7,ZPNfWfEg&AV[NIaL5>&#_[1T1Rc__OO<S^@cO5L/^eXT:>g\Y1_
;IDQ[)LN3+D9^bQP6+b;8<0Q/DgHT;;ZZ(6cLX<,e77BYX7AN\W3F(VQRX2>;=d?
ANR^YS,^DA5E+O+O(^cVKC?HTF<9Q^5GWDSLcUJA_(<VZ;HCdOTQ?9P^gZ[.e=0U
_K/+GLU9-K?A_AYO&T_P;dHY#[=6V;>>7KF69RSN3HE=FX,=#a\+RDH3BG18e-Td
.G:gCS#7ZfW,LRPR-L<Z\[e,R09/G@?WM&cUS?A?>\f1&.B&1LDKJP^fS)ZbAO+N
g#<(5XeC^.]f]F=,Le:E,Nd+S>c[+LV-g^.R[W:L8K4>3\Z>?-8f5LC,YT^cBK;)
Y]=2-A<fNB@YR,VH(SP9C0M>N^5-eZ8^,,YX&M7aMMf2)HOdJNL;ED;7<#F0-K=9
g&f4dGF.3Bf/E)WD<7E;&)>=5e3&&W-=@d4YK&-<AN\e-aYP\KTXF5=CZB5BC>6(
Ig6+[+LZ[HGH=ZfV826:eZG(/J@.332aK?YPdGY15,Lff3G5B>5WV,HdFN,>5DN=
3e\2<B<F7M2NJ6JX)&PYa9-A+&Q,TUE=8;./T9<.OI3XTg;<F-;865RFD\5b=J=+
BG_./.+9GQa/+SMSBRVT\T?DLRZ[D4GJ?=R>2&ZCZ-T(]a9B8^A(XE8WK,,H?d>(
AXV2@2Vd5>2.0+I.];/45_E)^QH3\H8gR?#23e>\BJH@=GbfH]M,TGMLK4b=R<(W
8D)(.WPV1cV\U-OFNK.=1^3C3UDb7ROWV8FKUSF-^RD53,M&dU1X<#0DUY9>8PU^
0_(3[5b=.-,_Q9G@T6RW/d\G96ZS8]VT1P_9-(/,,]64.G]gNJg73)YbV:a./B8:
Q2[8c[A716=G2B[eGY3:a<9D7[D,.LU9PQS?BSF\aBR:ZeW:X1eV#1+BHeH\Z6_P
),57_T.X(27ZBRK#:Mf2aPQ&81.Sgcc(4a&Q_IfCUY6N4.6?c.JU\+\LOF#)HHE9
AFVN@6K9M54)S0:VX@QXS;)/RS)7geMYM,DYI/67R^G+6J<df9fC@1=a4,+,f5#D
NaX7/\5V0]eG;:<3/TE:TC81T]M:JcM0]37[eg6)>[_IaZGMD;/+4/Ee?P7WY.R/
;8OL^)R^VQRVAI)T07Xd(&?ZPREP,E[b;CV5@WYP;A7RN4d(VXU@2gPFUWa:3_1c
,Aa@db[GbOSFL.dgTNMJ1<Q;\.AMg7AQ4U_,J>(\Y<J(&KMH(UJ&bAJ[TdKILU?V
(#(0RL@a2d1W:F8908VD04f3>L/.4L>cXO8AIKTOI;QC#UYQZ,Ag2a]Z+g):#c^a
8XcEC^g<PN]0IK)e>O5HF2C3:699DPcOdW(9X?],GY@]C3)Q#;G=Z/W1Z0V1C6\\
N694.93RPcL[ZW+B+;</35#<L+Q4=S<Uc2@Ue,@[;eW]Nb[A)gW_4,K@DCOd7Pe?
)K+8/]_\R^fHG@5[4AW4>RfA)S];(@.8\eK-?QZ4EXa+&D?#bXgO<c[>+cWD2_g0
+^A7;PBT(7Y1=c(PRPMY-E42e-Z&&..J7g)?_Q)Ud6,Fe6HIP=>;bB9c>3>7@8g6
M^gYELQB&<Ig53#5E&Od@8CT\&#N\:LW^#OD?Jf-\C5>_=A=P=b_=-;gBc#Y[Uc-
^_<4>1AB69:@bF(URgJQYfS(4+Wc2/SV/?/+QH85=A-ObI&^eA<<3<)fJ1(Of]8b
P7<1K&-&-A#K]f2DGG?P7KJK0?T91&Hb[6/X:eA6Pff4RM;X8/:WKfbHIM0#^ZOH
d;b9RUTXNE8c0gE-bO+IaCS4<)H.=Y)?]J#N;U[)Ec],.4.C;V3K@;LO,9O7E#F-
>9H6+2_f1R)Z7baE^=4QVJe&TEf#>5QU)IO5bE6B+F\K.X(O))\1\ZB^0H?H2D,<
:&:8A#cbCF51=F@\N?/+A9W/B[2fLWW;gRZV-=;gAXeW?/ZY3[&fXSPAKC\d\U8a
?cd<b=9.VQ0[ggf+830f6LW4[@4c-JIY<(V4?Tc8a:S.g(S8.6/]^0cT71-9ZBYH
/&SB?EZb@@CZZL3PJ+XQeH5]2g]S9c(J\EeUPS#;6T4@JI=.]&bP><7e76b>8&Mg
MHU<V&XeE(Fg<0fTHb1ea1,e;S_E:d.b/J^e+)?DZN1B-V^3WYeBTRRU,?cbN;#/
8PQcKDfR]?R+/5bAODNA,VXPBHCE+#26NO>)Y:9_(4U7f2[E:+Ud:JVH9(@1L@&B
2ZB0FT6:@MbTg)M6(+E=L/c;D0Q=5CcM57)_IR#1H+\=?QCIOZA9?YCFOf6T[c)3
XbJAHe5/0fGMe(,LWVW<--69MCZYD^L8<J;_]+Z+MN]CH[:<+YOEbe51;U3#+f+L
BQcHVC0TF<]XICL,5DI:N:=Nd0fG?N<P#_53/DPcKVK#aS7J4b;IGJY)P6Ma+[RB
2X[O[BQK&3&@8@2M1A]I4H7#)#J[IR[#<=e68Gg9K)8+ZaI^D+0-/Z5gATNV@ZG?
Ic.O,#b<Lc3(K,BU4DI9A&RN3C2L98OHa8JT[I[S/O.[[.A^80C8LHY.c)OEG_GR
))T_=gG7ZO\c_-+ZON=FA;08?[Qb-T@g4PW>/[2?3RePFSeG.JC#EgR/CD>-_Z&]
Q<aM6@.HDQH.a)Y&F+4^DbR=\4G(Md?3N@6Zd>K#EWcbQ,f/^[D3V)0f?a@T/ND/
a94dE7_..V_=5:F:-V<DTYZ(1Q=0F8TYbe8-gX44?35@X9?/(WZ:g\\,(bUT7R_:
NJ2BCbKB0DNP.5a,UVWS07G(-e)UP,K+VXI-g=(V^BSOLRa\9V1V.c+GX6@AAM1f
@8D#19PD9R2J_Od]_\?)0I#S8eF5F@eY0M0\;L-K>,:=[WF3M[-KeY=SaA6f=.&=
^V8HO,8/F_#&;Ya\]>,FE(GVgdN_>4,\BHXb0I4SL7f;81(T-0M_+[=O&1O[=:3g
<<2Db.0H^MFf.RWJ<W8dNWIf@8L2eEYTG85GVHI\V#c.ARGBQ0D-^E,d&.2_S=SE
&L90:g44UE(CMCc52U/TLWe8ad+dG4B3=;\W7AeM8#KPRNNf@e^2a^TfKeVS<Z&R
aL6I756eP^_39JME7W=1:HV5CbYE<4[dJZ4L)^X.1XL3]=>L4H/dR.2+>d-XaDVf
?<HK?[BI];@8:0,-(VN:M;cJ02K4G;YE=cE8[X47@KM9]&bOS65AMg])fLD[(H-B
/V.2VR_gHFRBZ6;X#_E#4@\]aZ]gW(E&)XU0D1W/Q(1^2(?8_H];Xf,YcR]b)@BG
CbBE?-ZT^E3NOg_+Y9<P3FV5NXed_3Q3KeZ#ZY=N,QJR4(AW548b9GE0.&BVZ?Tf
4E(V9-0LH,<-dKe?1D6cLY>ERb@CN)^FT@V,6;-2(:eMc=3BR[EN9165FBeYLfBP
(_R2Bd:ZR@c;K)</DCcA_<18]a8VW)U_efJ[?+fJTWgWX]WK5HgK(Z:?V:gIM:8;
5E^41H82G@NeKE-ffD+X/Tdf8+;5G#c_cPecW_-;/D\=T]D8QVS=6f]5;abdb\]U
5XZTVWCb:E]eT1._J4/5EO/?<T7Oc/ENNKS<&=c<R\M@\XfO.a&\c<R)9@S@Q1-@
<7S[LY.0?F:4F<2=ZbLZ^FHY5(TcB@CP.=GV8@;VK(58=0YWHE7g_;Y]SGT6.UYK
RbSaWO?XC(7A(+YE?FJ/\gRNJ+fb._?UPVTQ4Df3d1]<7GFO[1[KeHWPEUFM&ZS8
&;=_33FTM-4^Y_WOC(B#M7A;26;;1GW[3SQTYPYJU)&C,2/3?2V@aU33GeIG\3gW
-6LBF<)Q^S,343TLa3S?:;&b=Q\Wf&;YbBb+PWBEU]/4?CKcBR.gd3@YL^-MdX.Y
@#E31&20acf=7[&5:1A[RXcBO;=81,^/RDVA7STLK]c>+106Y/A9_3WA/T//M3B)
b+6ILDYaf=OLC4[2KZ<fT=cPf1eL]C4L3T[#d>J/K^5-J,?Q@_E2?@,V;]g@DBH(
;KY6NT2^:?WYCS_L^,EEOT9H];Mb.\>-0+.QgeMaP(<R4:49K1[GSaG:(bC89P)+
,D6;E3UR8@31T\13NG0K/(f5eX-@Q?gE+e9R6&FQ,DM8WceWLfJ#O)]?:[>TF-(.
+bMFc=I^P.G=9+J)U-ZN8aFY0:CVA89V>c<0Vg.#J/X4S:V@(@4b33K9ZK2?;8[8
(V+OE2[b#cAg)O_6A&1&,]2>>aPX0TG)S=R3K+L0=CGdNC0_&B_HL\>5DTF)E@1V
3QCA-87A7)=GET>E)@S87JZCPN)\C>=+N3/;IWVMbI9[\HD<+__Fa.(-T<0Ycd<V
dB<Ne4OcPG>(aa__F21d?=N:DfgMR]f7K(R4a1.N^<H0[I]D_DZMCe,NZ9#427Ka
I<9\E#QIHdc9C(eF9LYJL]]?535/<)7P&^AH8OV:MQ&6Q;P,B+=V1^(]32@>SFXd
FYL5]^QF5e,&5;BYOY0DbGf-^YCH9aX/TScc&Z[__:>(U/9Gd+=AD)b\<F(:e7IP
V]/#e38Q&0;OD)V+3L<8MZQ@@SDX4FZOb/d2W>I<Ie9aYID9.((_FCIQDAb/+JH#
26:WOMBN\MH7M7bR(&)/>^[PI+81?^Z>(g5CJ3P>:)-I@O8;J3C//G^[LMSX-YY)
&E>C85:2P)NV#4N57KAgE(?;.>:@Z3-_RUXM7dCaSfO0LV+c>(+-,dSW:(C[=a\I
fcA95Oe/1XTOC@VLVTe#<[?f:O5VgVU1a^Pe+C&F3JgJa=5@eF/,Hc_X6bX?De3B
-9\D1g=S56&\eIK(J9/+1-6+>#S.=T,[fB(g>GLHb^HKbWb2FVf9:5EH3PQOM89#
9H&0d_D/0Z#1Z7b=1@.0cB&eP(]c-(U2PI4/(b#>;A/(KNJSH_^0.S3;d+Q5MX#d
.67ZL?.+IS0Df@a;Y-DCZBJ0f++4Y@^IfVEHP(O1>D/.ARb_BWRZd\f-OQ7TP17U
_IC_;[W^_89GMUT,b2cDF&)E61S-58:;?T:cV;FIRgM@^b1U[QWCS:[LX&f]R\HG
RfVZSJ)&e2Pg2=96BD_B,d+)L4B5<<#UIV,-;G&U5B\VZX?+HHSQYHJQQ[1fULV=
](?U@/0ZEA_.[CH][Y[M>((a>gV<b,cOBQ33^1c,E:2QD@OZ?E3M31K7I17J9ZMB
5TH],?_VM-_-U_\g6ef549C(C2[_LR2eK95<N;/&L5T>;IIT=_fU48/^3BFK+H(M
+SU^V3TX24dK]/,D>8eQ/P:03W@@ZR_#+ANW6[#gCW<63bQ@E\XNg1M7E=B7;(+S
&C+M-J+=L&&e#B<:4b2HKE;X<O,N1F0R(4aR#M)::O.VcO>]Vc;>Y?fNQV<^2-QB
1)KM.7D:BHRUS)^^c@2)9NMOfB>K&c;_:76JBc:-?V]@D--a9#URCBLQN2X)(]PK
>1.Q+FRFE9]QBJ>BP#,(VcLN:7O:)#,BfO+3CS+#[(/EB#4::6>><LUBGM9J\Y#-
8gIeSR8J>W]MYLJXbA5+aZB,KYNcBZEOV;CVCQ213>][?=)5IEF@46/LKAB)L@dZ
P&Y6)#15c8/?#]f]9-+b2[2135L_\7<I@X1HCVPNgHf>.ZH1)YM8QY,H@5Kc0.f:
7IE)?ZWY8bMW/=&;O0Ob@@@G]E&GPV]fFe/@H9bYS<fM0Z&K4_7)_B<F(]7LBAbQ
bcSC+9NULPLdG]/<ZP?g<[Da9UZDdb/)?PIfMcJGU5L-D,E]282-gJZJWJ<OPGDE
GYe8M-+8&UO7I^VZKSHZ^3Wfd+7_UW_\3JLdS^(^U7SW1M3N8/+#QdHAL3acH0GQ
Ld#N(PSM=aM@S0KJZ?V?][_#FQDIY11M/Z)N.-I7O0+e7=?TVMB@8TgY.A92LD\d
A(HMN)(YNJW=G#)7@7KW[SMR;]dgPfg)S+,4YOC5a#g_0a#[2E:G,A#3B=;eQf8S
B5f?aZS2J\=V&8BCR+OfZbF^TQU>P/+ZW[aQK>J2RU3dWWWF<_KB=CP273-,d[OC
_3Wd)=_6^-3f&N9#.XIF(U^5NZC645R+N#Xf^WbV](NB^]IY7Y1V#;WV7VWY&;PB
gA_9d8Y/[NC(YX.2(6]3Nc@_DVJU1REUAU;;A>+(;:#C]9#E.:aRE3WSbJ4\6S7W
egOE_a57&N<L<C=U.Z55AfY\&#V+S3_?Q.O)0PL_Ag:fQVFb>BELCd7D,UA5,L+B
cNL8c4(\4R2V0QC(DTcT\E\<#LZb9Xc-a=Z&_C/UWf6ISLA.C?5>MXB7RXCMG+<R
;G&D&:<^]096]SVW<U(gTQYc9#&LYSJB+J4<gM/N))3..f4]2=_N@LPVLRKWa:cT
4<N>++\IA2X>VU\2fSD]5^FOdd&CO6R<=LY91NWX(+C+T6L3BA.=9#4LC<PU:WZH
>9Dc?@(2))aBQbK?(5@T=D;0SS33>)_?->fE;Id>ZW\f6NdO:1BQ?bWK9X+YK>d^
RLNINDW#gNbfJ]DDU[G]Z]9VKIK(R5]\B>&=d3SVH8_Y_^W+gFfLCcaQ0O5:=X[.
b2&[W2)2#:(^AKA9Z+&7g[XFI1B1.eB73fa13Q=1>ET#6<Qa]S2b1B6B19gW#Bb@
QN>FA-;]d_-.<]NRI9(aX@Y61?][VJG_6VeG_U56c^:>/E+/GO4GS-NU1L]U+d7<
GXbQ9U16@WfK9Z3/G;a5dURUId\ga12Q,#CZ:fVOdPR&<OG#MTdK?;gZeTY^I@<S
JB1AcR=1^KC;SM:fG2VRdU^PL=M[-,78(@bDa&Q__O3RJYOLFM5CFDXL)A[&,W>d
.@K/abe/&\=CT1T-\XYIc,<bKUBXdJ:C&(0e0X_4=dLKc2;(dMDD96)]UWfQgG>/
R7UV_?BV#7V4@9f>)\4+UDD_;ZdgC&DX]KZ]\1KJ\QZ:B]/L7[-B8f=f0F;W)OM<
6DVDY3YYb2-[HXQGBf.3bVB\LH./QA4),T;7_@T1WfgC+beX:DgNS^T9W-(,YefR
J;T57&W=,fg#W^SX4#KBG/VVPEX]/]4Ec7KAFYXG5E<0Ffa,=Z_?[Uf9d8OOW212
[_cT+BQ#H):MT&,G7U3.fBLRB:L29f&GSRYO](Q8>^J3XU6BFIHCd<MZ5T.d:UP3
\+LD.+-BKRHHS[cg3PP(Q0<EMFUE_:W+;[a>JDUBIPEJ9\&?[[R.;_X<CGN/-2KD
+f5HcW.bQ^JT2))N#Y03^^8bZc3]&2@4,MTQ4KQ>,Ab;e(YP]^[W?Z(@OZ>@0d=@
A62KUE<Z3)_7aNL=g5ECDK@U8c8)MQ/G_U,NRGHGP&;>0-]_A&.BeCd6RSDJZENR
G0CP,@7[((W5&TNGeVD]=-ES3e_Sc#VY(61U.b@AW,ge5eXH6M>2++-VBdX/WIW\
F+@WdUDV>,/Z]C;_/;RSdd[H\A)f[4]^=S>.J>,YgeB\YJB-I5T.01H#D\Gc9@3U
F]aT;fc#AU#3VO(8M[7ad?N5Oe=aUO]V@68(5+2./;I\BAeDcL(CB4/@X/:QY@#2
cUEffd>=[QNW4fY=KVd@3C4QeEb]-U/gff]Pe53J2SPQA\@&Yd#U9a7(4TX<?^,5
AO(D)6OQ(A9E/Za^=fe6#e=U)O)BeDQe4,H2&L6T5[A8@68W:]RU<OKG.b9Qg@Dc
b6Qd-6\;1HO@FZ)K(K9Z_^Q,SQC-.<Z)45RcX^HG39:-1@8K();I8(P17NC9+bE.
=SV2[UJSSVeJ+50a#_LU?\EAC1<?KM4S5^Gf?f?2T[?VP]-&M-(U/F7FaYHT)25#
e?XL(d3)7IM^@b_6aL-,=9[QMY?IPISKgQcfP0K:RP\S]-R:9WU._2^6=DELG4DH
1<H[\@a^P&O2^fKb8D)6B_HCEMC9@7P<V597S?-b;B6/[=:2Gf-=1KLH?6TT)3+<
^2==/Q&66S?R6G^+2(0Y7GH9N&558agNYY3)Kf4H2KY0BOdI;K8_21RA0f.V8fW^
NdG?2Gd?C<M3[f22>bTM=F9VAeNSaHa[3BZRg(EO\dB6O3g0<+.?cCbS]Y+6?[IY
Yf[T,][8(TS>5)SF2-;,+)ZX_V<J<G8.0VVDJ43R<XD2B]DSQ2-O56YDT]SU8cTd
RW0.I=W.;+,DD4D.V^fLP<e-8CRX:1TJd:JN=@ZQQP4GMd:Y.Oa9.ACM=QK^1XU#
6]:I=>MC^HW2<Y_AUSUZb102Gc?XPY[03<.DPI8FMYaQHfT6I#JJ#H:L#8>=Ce.&
]g,>9eRT>?RS]Tac7.g#&HNI\4U;Ja6#gYY(]E:6:CaVCI_U_FQC()4c_X)5;:&-
0LeGI_4FEI&8[X<b_([I)OcaMRE-#^OS=FFd,&(8_9bCS-#c<QXX=^)VKKP:>88a
0ZB9XM[MB][Df[bC=g9c\CUa4H+cEXb=7+QDO5Y7<X,O@GXZCJfI7Z-H9Y.290@D
.=Ob5?I-UQA8dHP-Z?(?M)Ca>2J7Ff3aL&Da(VOEgLdNa:47S/[43Dd(D_9W&d9]
Q1\a7&_c:\QDe#>HBCW=#G]E5@3gFXSCQ+#E),IG)1e&H]5R/69+W+.Z>96+b1:7
/SQ[^A8?7\c_eKG.43T9=.PZJPHDcaObfJ3CZ4O9J5Gc;]?4DV^EZY#VTQ@_@)E+
Xg.3H+Kg:7EU(gYB=#KdB]UG:g8=)H+&CM74,L5DZf\I3e/T#D8eZOP1=5aVG-fU
->d;-C,HHS38Z^SWY1agR&N9IO@#0M#EA/Q-2K)U/\_BaS1>TEIL>^[N;,.CF3J=
>6SdggMeN&Zd\5OJY=HS+S0UDQ,@/WH0<2ST)X1W[44+<aABDRBSOB3\--cG-M+e
]@\cCB(,fVcXQ),d/-3<6(e^P8[4U^^>D1G7XgH;7Ha2D8Ba[_@ZHAN^WdXNf#1C
9I[6a)ga.@2Sc;f7&5C-J0&6EGFb(NHg9([.>FV?20\8H8[S+[L08X39ROgUC]_4
8\YJg]RdgL5UUeONK#8LC892bQ)5/-.aW4_,^=IX8BLbf3YCbEEAP:.64Y.&6FJE
e>W1[J3c8Y9=GBgZ3DK98ONa>FD,M.0#DPRY3c:6&@C/23)J@BGT8/gbcS4>SXM/
&<CD<([@ZZFM5[E@cTVOJ_Q7LOBG7Fd[==^[0:#O[dPI(dZ;+(OU^@[XfcE)SU0T
L)F^H7),TT-bRLAf6+5bgBE.)W3K).]GPKI>A23=3]?(Tec8P9+U0&X0&d9BE67Z
_;W@LJBXG\ZR-;R,Z=]@/WQ327/_?,:\_1,P[6WN](fW.I-6,HY.^&H7[GE:5N=;
XF+5eEO=S)Aa;?K934]F/g;O(N<5(aL4?OQDCg7#/1,^X;_gb=[=4>4-6H&+_]A)
?RAFA3c=^((/@^KKbTOW1#KUa7INXD:3&C2<8?1g7c[:fAK2D&O;^JL7-g8R8Z@1
M\&4RP2?LUEHD[,9\7d&4CFBJ<;?6&H@CHND37EHJF&3P,a5]R2/RLT)e:U/Pbd3
IHY+ZVH2CP.U?Jc1NUDTdeG-9aD>]1A-R<Z6#N@f(e:R&6O/B)2gLHe8-HQ&dL,)
9@#S-?8KUHX)2cHSg5IZP>UJAD&8H51:a4L?)ded/6WcXV4S-8I/K.50^e(W>We<
M?4Z=R6ZT6?9Gc+7;VdLL.VV^Sa(bZ0Cd@4U5J+XfVIg/@L+=^6VdD[E&GV?D)NY
5PFK=^,[WS[2=K[#Fd3;)D\4.Ja\fO9?&-(Vc4CTf0_d,_a@d/d?2ZK77=,TBAAQ
8F21&S(YM:KDPJ[N18K8S2#@E,^(gCGYI]8A)U;=DG^O8_d]&4Ie<I4J1dL\a1W9
)?aT@[g2LV?9PE=:UG/6.b3F&78&0C2f5@MYY-,//T4)J+Jb+@_e+/NLA#+KCHPf
W_DUg=49L\PZI&0Wa-U6TPQ?)UQbJX?O+/UB\Z?<&,VBY]L[,;41d0;I](b\EKeQ
36OE#6C3,2>Y7eCK/I&_N<#N^FM&\c^W,41^TR[6]+fB^@UFV?4H2JG=W5E-6/aI
3bB=8,_[@S)5HB]BUW8c>:JMNM16<AdV=.B9Uc7a8\G#NWWc6a/=]YT-NQW[2GWO
d[T\=^<:B-@?TN+.UV;YH(Q^9L;3=GXSE@;C079C0HM59Z5RWT7T1A,(:;N>:RF<
KX+/gSB:JbYWVHFa(:YJEF.c1dD;/>7\D+dE;HOB+H(Fd0F1I)d(VK+(/c:e#6e>
QZM+\YFMJ2V]TDL4,&3K[>IF>WB^6[AK5^abc_;QFMYM8VA18LL?FQ9bYV]4c_14
fBa.YW#K@:P>+=8MJ#T4KdbAbQ8SSJ\4aUZ(+>.2F2X&<U13Td+0A5^VRMB\#&75
C/3D8:<:0<S+FKGGP^)7][7FBB(/VB];:<]42L>Z#.?::EI?YN58.K&Y>W-ORZ&7
2917JbBE?Hg3fc;V3e],691>HIPZJ:_.HDJN\XLW5IEOV]8XD@B:)GEe/Za/PQY[
7=26AdOT1NH/,_F3XH3>3N6O)RD9)gdV-Q#J#d;EF=,B4-cA3OUSD-EA@f\O-8??
dIW4):3L^82Pc:=6b/IJ@3R6&W(S6C32X81HVA<<I^f9f=>#=gFP3WF1Q;3.eCPb
CR0)cRb54.UW95DJQS/8Z2COG^dK006G(>(cM(/ee-?Sa.GI&6KNX^3;@T:HMD;B
c+B6aR@=/dgSb.G^.3,>6\g\^@B];/ggECC_30_f@YY.@a6fZ/d-Z6)>?:@1b/90
3]_0VcG5=OOD_1WZdYI;+?ESTGZ.IS_3FE:EQO-VP(G3/U)LG=);6Z>0)3P(LX^1
]WQ&]07[.E_&\LggL6>^dJ@W_af[&JEDB5[MEUMGI1[LLPR=@079UZTLc05\;Z^V
-[]<NM:-d^/4dI[SM@8\.-KXD[3=ERM78ZE]?^Z]E/c15H<NMg)b+=M]VeRM]3]A
()WE3\5>,EAc7WGEGM](dVeY>^QPaZV/McP2TY/D-OL\MPT>Y;f#N[3B^)R];1FG
cCcd=S@8/6UZRT,0S]6;9I<OFABAE:[LK[afBdQP/;.L.+:I9FW8,5Q#QaV[).@a
Z<Z=9MC5YCb1:[AB6M\bc8Oc8IN6]DFa#CG?+/].d<Ja\4@+-<Z4/2MG4M+0-#,D
SVVT^3?KT=9+L)04M#S]MY2=^5:C[c[f,ARO.XA1)e<5RK=-,e16bPUYcgJ>cR\T
C9d_2[#,T9-O):VL^;=JF9H416@JSWad7\#BH_-+XN[/a]O>Qa[dE.@&WQbW4>IB
bIB?X@FYF;VYZ3@Q@fPV_L9f&G)N67b>.2f8b5((MQ4ZW#WgWVUaR#=@#276CC_K
#XE;c&D9c<baKS<0\2a4c=_aN]-G7F.ONS([9X,U/+7OC3Y)J40T?3NT;:+2e3?W
DQe@<<FD_fF7CN\d?3PLYGT?^.G_&(]aEeg;7OT.QB3PCTJXSUZaAL->ST;I5e(a
YQP1[;b-cE[#8[AMIZR[E7a,IZZ7Y)5cYb6[[dSHNT;c/A=/VW[KEQ,Ue]\^O2=g
0L#3U-3\28F[2KGL8U9ZJ]+7F&M4f(W3JC1-H6I/,RLVWP7B@-&F:@6fb;b]Bc]/
^9=[f-CL^[O,gdVQWJ9Z#.WV-6fYJY#Ie9&;LQJ01,Kd-#TSOGS3BS9Y3^(4gJB&
0O-gK+ND6CS?Y;V3bP:Q>bC@2g[_DPK@a)S4O,XCRX(d0L=a:@=HRJH);MMQYb/K
Z&6X?A/8Z\]:I<9X>(Y[49T^4U6O5YLD4\Ge^acKZ6AdRB2N,BSV;L]ED\/Q,(Fc
R=.+8N)LEZ;?,#UFZD^g9DbBY-TQ0P/+#1f=_\/LJ=Z?33/\#dS8d2NJW)-_Y6\(
F)RIgGD8QSeO;d^AeWBC_YLBAMa>6AB@+#e<3E>U7N]R@)A(3_QZNCedbZ(MUI<9
b+OH#H4US&bceFJ_bO9d+1/?AWLE>d@c\K-OTc0P5OLNP<<LKa(/75?JN_?SE.aU
)f>K[&9-Z<H>TVJ=(23A/Z=L8EYb_KLA0[PU_#_GTa52N.&;Vd&+?NLS^7bW(Y>^
-NPe/L-(;GZDU3=Z9LYANSIX_^&]R/ce^OHQ:I5VP-&Z-].::Yd72B;NUV.&.I2_
;?dO31F&bWURD7H;GXATE=;?If#2W63P3^1X>0]L=&KDI=]S860O_c>T@IXYXCTO
MR/V<.SK_]b(30)9a7E)<VY7I:N-fY7C08/8T-3bY)D^R[C-#Ff.P]CS/>KXMWZf
aScC?W8^(5[K?-a?@ST-]:1/5DCe/:K5)fa3B^fHV?#D-b[YKD(5B+9PW#]_\_6C
aET<YIGH-;A_S+08EOd.#_O#W;P&49Ib:#3I#dg(Yd1::b:TQU\\Z4-4/Yc[6\IP
+DEV9RGLIH]cDWW)0=8Ta_]5M]fU2-[P@R+1F=8822&6I-V:eb]5OEd[3\7U2/AU
/Md5]XEG=/H;(E#M&O:bC[eB)DdfFbeTH9Uc.TIT&4_d1FAf+4)HbN\2^9bY4TN7
5B9T05^NFd=R<=DfObIYeK+FM;dT:;[>Hgb(8W>EUCD/5S;6B:Db7Q;Y-d]<>F3A
X/Z7AN<2&^M,#E)5<gNE<#eMAN[;dD,cSLXW8NOT>VPKM>cL4E1g53PLG=-dG:5G
E0PGUJ,N75X;faPCR^dR,5_PA<OHWVUN1^((_X&36TZe299O,#F.^M2gURYW8Z)T
PU\)/Y1gY#eObI\J2UEX,4:a/R^a@c(^Oa,b+6Ra,V5HaIK7_=.N+VR3Q+S^PEgJ
1#a&_=CH58S?JV6M+4X]#OW>bbS/XFTCcZFK&5EJSc&?)c)/P+Z1,agVdW+8BIG[
5HRE4U[]N7)H]H9^Z+a&bVSW.1?=9O3S=6&LLO#NGGDX,P&(6W.3+@e7^4+,Q2cF
@H+3P.4:AOFL\1LQ(/GE7M?+=TBODD/^c^bV.ILC/@5T\1;3CP;MZWKYJTB+g#6D
+e70fB\#<c].1+P;5W\?f[eAMT9Q^9PF(_LBG+)Ce9XT-,2G45BH,cQ1eW@.:.\E
0R?3^b;[P38<K:Y/]E=\KKScH[+(^(E#JgB(]g=&N:M5<#M^a]1VP=URJ@S25Sc:
d:)CJ>+?YT=bF@6,-<PVf&K&9gMR=?A4A8\\5g0YR99D[1:-Y;)RR_c>4L0gc;c.
#gYQ,?Z-W&8ZHP5&+QfZ7X[<??<+3&ZV9+E[Bg<+6#eT/C=5SeQ2QbV&UQVb&O^F
N9W[6ECFP&db9<1,Of.\WJ[76eM=DgN)PR3aY:Ge?f,;(Y;20?QD/4.CcHW39?aL
[4V]JVN3N/eJH^V[]QQJYPKDU-CZeQCG0L;.W??7RTOV[@=.@ZHWH1dQ^KEY\E67
A23N-YZ2#5E0E5=d-:O2f/QG)EW^A36ENF=VY0e[A;_P>d5H#<2J37>&AI>TgfA1
a-S\68.64^HOQ:4[>.P:e4_XKE@[V#W,bQe,4/]KKcAG:G.B4G0@J(D5:LD76XDT
PX#-/PF)FJOV?_^8+(9NV_9;:1\U(;WL2f[6UOAH;FZ@/PTF]XR^<Mf&^;O<>e<2
BS;8)0=?G@DBT0gRX35RP)#?a4,EF)^^Y/\X(,0.^ObUMNO[3cD,8NFRHcGb-^c3
[79N-5c5676[S^P9<+F?Yb_5g/R)9G\I;E15ZGS-7=7J6b.KfBN=6ecJ6b85ZU19
]LW5MPOa3-\5EeTOdZ8C#^95Xc>CPTGJN_=P<R#P:&f+M87Qg7:<e=]]\7H@4?a7
WUE1_;S,^0ROW2I)a44QW+KTT3CdE063RIE_Y;S-PB+[D@2PD2P;\<aCIbWFF2Ua
>:L;gI<2>=6WD@,Lcdg)CMS2E:MTTg;VQMKL2;&AA:Xa8&ICb_4ILE/3>bb\OWgd
ca,20G:7R?8<OKDW+gZ\dfSN8)]P4\I[L.K/N1C\(/G)+LJ)7fFFKFF+0692WLH9
IPdgM=R048#4?D_6?a=9WB+eZ-TBf<6X(6cfIV)bO.Hb/f^WeQ>O4@4KH7,0CFOK
F:4@#<Ce[9.:e=AUddXAP4AX9DTS@VP#.?G,]aFAT]0Z?G0R&JF&bSA.69_3NNeO
B\,EF?(CK20.TdAPaY.\c<)EQ_WG,PX,8=:5YBb9S<R,6\KW?RH5f6+fSSAITPH>
:6D(KB?)MAYJ&NCQSB,5X-2CTZVf[-:3YX8OHXN/cO[]898abbL6)agHfV^0P=S#
#Hg.0TQ&<K,HcO>WHA==COU.[I3GcG-4ae@RIS4=Y;A/N?#OGAL)b1&/1Eb9U&a(
LP7,,g@Q6,Y7e1Pe]9Tc_LZ+HZZ1XSeH6.f?.d9WVYc\d,==<)E695Yc[LRFV\0d
B5CI+<7H9^cd29GQP5-d@Y]TD62X757<=L14VbO?cEMY?Vd<&1M67IYN6KDE^K.V
=@7X_,X<0JSc?.&C&EY3@3F;>Uaa>[_8MOM&KGMDRO&9A9X7DE5^L/_[/).246CS
29FSXX>6<^@g),&[B;QAfFa=0SeZ^:^)Z\>\DX+f43+96_MY,N,TY.JOX6+S?Zd3
O]82P)_]2aaPBZCR\-?Y2d,;M[<3c&-@GW91/.0fD&eQ:AX/RT_V?4a\U]\SCUV-
&XC9BNVI:bHUYX)L3;GVaAeP2ePN(LZBdE]#Ib4(22.:\U5E@G3CWI@<)2K1\\D3
J7P]XZ0575Q-6.@,U.c/F7X[VJcg:H@DB@^;S6e>:La(MEOcIZ.W;F8MI/Ta?+BY
8_ZFfgGbS0P6<dYUT.a#f78UVVL8OY0H<<[HID]\;?XZWdZ2/I[9>+EP0H;#PZI.
e>KZX+ZfNP7T^&OEgK2PF:[Wab0C<M3eL/ENgM9GXc@:C:NKHK1:Wb97?c&(,OUT
cdScSI?=?3G1W#.?c9GS=1Xe^OFW([50WUX\_C+Y1L8fU;7M-5U./5TU.aO@(Qc+
.40;ZFc/(ggeBW<2PdX+J)0]\99c3IAJ)ON7,J5ce8;?0,XCU0[IGBD:Cf<ef<QQ
Q.(@HY&aI[4NP_CE#S5&(T5Id+d8]9VHSEE(_<2&cNV&JZS/0CF#-g3Gc)^4fJgV
^:PWdGQ)cg_H7@5a0]d5V&c8VSCXY5D^)QP,.A7><?C7#&fV>HAX\NG0:(LcLFLL
RZ&&2#E&.371X:LY#A0<3afC#O).MD6P(eDgHOO\P+7OX[?QHV3R#a?17a0^aOW0
X<,.W[/.UQM1F(;SD6(eLQC3cM.40R3OOM?65(&E#L7)dZU7RRICA7[A\ZO-c=X(
aRdCHKN0QLg&5Q23V;++[9dL2&=Y+JD+BD>FO;N-]TKNg1/+C_@V[DM9(;PUeV8W
)2@g^..QVQS4aEPVdLRO./fJW#N9],WeC=Zda<bRAJWcA^dWYFZO#c<Qa)O8B91J
QQ1[e8+P=(IFNMfN(e.XP<+E3cdaS/=DYHJ0@[)/,A3KgCI3GJV\I-d.SCAFD6,[
=VHeYPY&fQ\M;L-Z3/b=G)bS,G(Hcc]388J//fGIHL5bUHPY,XQBJEe^UIFOXbA\
/GKRgD>.=/FOf>-P]e\CNg04FPYRE^bKXb/J\V6GZgWa]U^E9J7@OX9T^9^ICENW
^eYeb98PG3YI1-=HPZebag&PA.5^R71XRW3ggZ_WJc8WCg:(AAKY[;SZ2e<&b_,3
PeSW5:]@PFA1;HYX_8[_V2/<YGQ)^A?fW#5RJcQB-,\2fSC,VRE2-YY77;C0[=31
e3-Q4PK&dWf3?UUcW;73Z=:[3QLP3#AZXRA7/8]^=NRYe#c1/TD=0dQ0](35GBf-
[a(&L2cA&Mf,ea@=.TU\g+L[U4ZI&YWI1M;/M:KfcTZ\#44K8db(g=[J\b,CI43#
_I23)b1VfaK2Pf.Qb>9C^,R&8:0#H)d,C5/(]L[58g_PJ##P]CZ;Rg7Q]]^8Pc_<
<S+Db???M]E6a8WcUeSO&3[X+W#^c6U=<VP1_=OEMfbS/I,FGaa5X/O(c2#7A=:6
>D4-W/;YXX)V+R?8-g6JFY./gN;VQ10.AF.QD.,\-fS=]a2U))E>f7>O,(5e,4LL
AV6^bQ/[KQWg:TXQ0WBE;7V-E+@W<]gb\F]ET_fW.U-ZR#/9G(VbF=0W0ZYd3Ae,
a2R#+ENMQ(fW[GW>>dG:gB;T1#\<V)/aOfXZQ0/R:?/=G_GVWLQ>HT_JFf7(f_6A
#PV(,/,_I;L=R-cJN^3=7^\>IPHIAD[@[cO]g1g:8&d+<f>DU-]SAOIZHZG1:717
CA_21)=+4^2E^PI(D99=\6C2\)RF-R:(I^E1,L556F=I_G^-2DF5MS-fBY#>)U2>
J+;1I)0B(NK0UX?>f61K(^1X25T+JN<BYSW_/H0A;DFaRQB@bC@Q;R0T5BgIDPTU
;f,SZ/g0/^TI^\T^,9#<f72gR/#&QD.=POB<22UXF/LEc&:C52HCCU?<ffUQU=Q\
_\3K4@GDb>>8#KB_17CDQ+[LOEe5LL#VFM@7,g(AN@<57P+(2eP)H.W-KTLCN@\4
1?,CDE<P5^)NTG,WL5E^7DR8&F,FE=ZE11GHXSWH-(bY3PQ3[fEaI6f_Ne+4W<[e
dB=YTAXB#9\L+4]\.QRMFFO8#[adL)eaLAJ9@AdMgNNB_RVETF@Ba26BVCG-.1)4
aT,F:ZOU.X)\PPOJUb3>JD4A(NMOE,T0fZb+38,B=T@W5--#\)=AH4D7LC^Z,Y:e
6g&QYXZ)C^-A8NG+\=WD+a6N9H2e6-:M)\8#17.4c&B,]DSKVd;e9>PPY3K3(c/c
eB5gG=08:E,dOY.JYM[]^(]c6g>MW2M+@\>(_c7U6#>/2Y.29H,[-DCIe>G^6gCg
K-4^3QX8^78+84.P1)]LeU.2J^+R^(,5&L@dG62Nc.:WgeRT.YL,G&>/(fb:2dJA
3+KaBIe;B1YeJAZ;g+TQ38SW-6,M0GU\bg;bQ1NATTFV?D=T-O4)eb,,S4#S7_)e
65-CbV&-BN?d[>.[6E>0c;C>ZVG4WgIe\5ZI)9I>)@P#99(#JT&9DN[aA],S#,01
9]=[Q5fc1aR<2<59<X<b4)#E?ER;Y?DJUYa4+HAOC6RAd7]F&P44dR0GFF7FN3N4
C3VSBcP6Bb&b:@,8)8c6XX654<aHYTJBBc.6:F(]2]Q\b=e&JFc(QU\02G47be9G
YC+a#_4Z\?R=10(Q)7F5?-4R_BBUI7R<3Dgd(EBX#Z6Z2c@S/M61Pc50f+_UHbRK
1Je[<QG5X[H&D/5XE6cX790?O6,=0f&^.b0X84e&:d&D0G&T^U#8I5,?^:UAAMIg
Eg>OVd:(MbJ>^(4Z<85ca6Rd?3_0dR8OAL,A4.04-Q1=-;bD92a9=5eMEF:QLDcQ
d)4ZQLP(6@<(([2X2bI<>7,U(;WR&#3UP]:;>0@4gQLJ4FR7+Y<g(AH75V>@\APd
HfLOFD3gH:9^b3WY[=dBA8>=)A0)<TLBZfY5PD^J_5c#Z#.AUXW(^4;6P<:5b4P/
YAe+&3D?@1EG+OaObVU:K5I#E<EUASMITLHD7;Q5fOZYIHQ9;bO_07Fb:WFe(K-c
>W>;8HcSf-,4[gK^()<ZW<;4g^Y.5^W+AeN8)C+K)CdW9U5O)8DaSE?4#1Bb-H69
:[8?&72^Ua:)ST0XXbg#A.HaBcMTYZN+IQW^-V;N24)L7LIXPLTG]\+&68D+WfFD
c_0WgA06BFR6[(VU;BaCb)^\gR>+)DaJPKaRU8LXb+88Y)a.g-9/XdYPAU9f2L\A
If?9/>P(,^B[V.S^@S(TG38V]\XfMFa-E6c]L2F0@,4EYgNGaB2>OX49,-WB>&<W
UF51+R]Q5Qe@;S&O>62f;;=A,OJ@^Qbb<-/2HJg=<@1>]N,-=e;]0ZVHUBH1GI23
[#JD^KbPCg,QBdPAPf+IQ=L5VSB&@G?#cT1:)\Nd<Y(_IETTR(48>QX+6f&@BW,?
S?P3e:;RT@dWU.S9]-Q@HQ6f942S[W_e7VBZC=[CdeWS;WH;3\#8V0Mb6PSE6/\U
[I;E2[.+7.+T<Me_4C2.B;\2:162S_HABA5b2>E,;a6,fMHaZ@,O[\0Hc\>6GW@e
5L1U@;8V7L,[2&]6Ue-SP<1PN=V<;F-26eJOTV8e=Z>L?=3Ug&SeH)(7R_AFdcNY
?B2]TX:;cEggAc#2dDW.+XNbE7^gSR\DK0a]Y]-;1S@0U8K0K(,BYe&FgLHF)7K;
>cS(PM;>G06JTdY-8K1bA#?6Rb\&gf48NEc^6(/Qf_XNZ-].NEEA&K^X+0:X,9(+
7U&5Hd+@RQB8L>1A8eEO8N(MZ&9;3)>Mc0PY5REY=<MJ2ERX([NFA5#L/[;fZ5]-
_P(6-LaP9YQ,b=?@RMNZ?cJZ=K<CfCcE>F6ZJfA1Xc)G<U9IP4T6OU&2IPLcaf:(
E>>/\Z2U=_SP(8]^]@<f5]H;WRC?&d.baA_/@dgZ5FQXTEW&E+GBU>.;JUC&A,Cg
OA4WTZP&HeY;(#68bQ/M3G4b;M=AU&-I=&XG65QgfZ/O7d[(U:P=KINUH0I+_\-#
MYc8J\UPKYNRa;:Q;&H9Q>5#c0N<:&T^5OAYV8G;SJEX68:&V+ggSA7]gHFWJ^KW
&1Q1/>+X+#bdP.;:GGC=HaI96bW-V]LT#&^-<5ZSN&ef2GKVf=8E2JXH1+fG-?7#
D8T+08b+G&+3g+9YP9RIN6;VgJ6a5Qf71JIdCD2Z=,0XB__C4K(JNS:_RZ[#L?SC
CfZ6B(@AHY&39CcBZFFg\:YQ6^T-@+/\?ePMbTU:A]#NPdQRe5FB)Y0gEXM-E)&b
-PT?a</4T:N9CM:86.E@6;0ND#OC^K.ZR2O@NIH&+45(0TOK2T4I^Bc@GOW=N1:Q
YGD05]cUXVb7+^VJ?&(?6IH;EXKY6M)7F=7c4ZddgB0:^2V9\])A]ZKL9[;7AT6&
R_@98RBLC=V>WbUW\G(5ZBM,KBMf#e_:.^=4KeTN)/cd33]T<2NVBTIfI_G&6Q,b
F\[78d?L1;5cX=_EJZ\US]3;-L9O4,Kf_eZPX7)\D6IaO_2aWbTN55;GP4,13/..
A)^^\;/eI&\-c:?+#-_ZB=QN5K6,XdU.fEZ1(0Q\Q]&/HZ5gd7Mg:b(bH4@(IA0F
W((\c.0,ZAKCFe]aD(G5=RNb;^[dM<eP5<3MAAK?425?<];)T[+HW#f(Z<ET<;TK
.?F)K:3K#O;g40E@HZB:bC:(9I#@M7W6^U?c-U3/.L#@Pf/f#aTHdC+Q5+9?.H@>
8+);7fXWZX;5N.6fAJDA1GK<\T1T:\ee\TBfM]+\-GWRI]\=S3Bg,U^3^)\5+4-S
,F#?0-Xa0:(d+c&K^=X0eZQ7#V^+gSOM<(@2&K]QCB@dVP+I;R5)8;a^CKA389(Z
H[F/,(b;FaZVdJKV,W6+YfJaCL#/=OI4+OFeDMdQOW\N>?.8:9U]&&fXZ?HU2Q>W
Q7CN4\RA/SCJ>WWAM@f;22KLYWF:<D:c)aYf:;Y4YTYfa^[6T3@/M+KD>6SOK<M]
fYVB@52OWM=_-AQGG;VbG+?\VdS0f-[HYY#:P\U<0M(BQD=]+<>QLdSTTRH-LadF
-,QCCYT>QWCJR?g3@/G)\1gP3ba>:.d-07OB:b56UFaH/=@)-edAN)PUY7bb;X9c
&^2@GQ@>ET_dMD9TD29CO4)g,6-3:GCPPYD3UHHY/((#PQ^9aR-DV,TVG#WXb@CW
bYb&bLUF7#J^b=0<DD_3KO+T.H9E<;T:?e:NG2G2,4TRf(/R21gP95:R&C>M^E/^
G#SFdZWSEfUYa:E-;_,.2M6LPdOe8\AdR22EL51ENE>_+9EMAc=E9BH\dL-#=YYX
NZ<8-YM27>6ag?/Wa)7Z6E+E6H/HT5_F^=CUQ,/&[^?7^(.\63U9>Ud6@[RR@VBE
#HD\bMPXS]eG,<3B2B&7)KU[TIcDg+T8#-)(DR1-+5APSMVM5X9X&f.^H:_#1e.V
gb)6./eIZ_0FXP2I+<Y9Q_,MQ1:#.JCPD(cHUCb)1W(DKNP6_E6ec.-,W#I&f,]6
9d>]6U-BeKP66P^aLC5fV>O<QK;S2)TO817=g&9bdVI=UT/]59>Db4N0LJHX3]EI
a:G#,+]AT_66P(#.LM9TG6Y_XGgdd0A&MD3WG+Y;2:^G/,N6O2D:Tb>XfN?Y9\YS
_T9Q6,L0JPe(@X)[?^af6a3_[^Y^9KK.f4cCV26<Q&gW0]2=e[[0gA7MY8;#C)Q2
MZ]1Ae[NbEGO0QB#UVZfR;^cV^\&5J@P9^Y<FD^Z#eV-Y#FN\K@NB.M@K>F+60W2
@HH1E[fOf04O&g87a?#-EO@Ka.>>E4G,;,<Wg3>H[N&:A62e99U]&+2C>>/0ge_0
K[>cKZf:U6T28^GT83Ibdg;BOBBC+6>?[6;+Y9WB6ca5CT1=LGZE3W08,/+\KgA.
.@BH&0>NFMA1TY\)58@(a5R;=U)N79Z&\:=SIOFEAU-gY6a<?EgAUBI;4KG8\<M@
NJEB1H,,5K1#T,Z1V6cIO6K[/4?aJbH=cT.e8;^;3HLVGN8)-)><gU<<1\UT>&02
Z(g:VQd4^cbUgV3H[+K_60^QWWL(9UMFL6b/&<6.47HWOA#_/GDdDS,=P-L\8Ddc
RTOXEP2=:A#J-M?.dCB-Sf5cD/YMU)<Q0IFF>-YRY&U;c=TKgH^35g,-O-_eY\Ea
b6<,.:TRTL[19<M;#C+?T;@=QSS0,Q7392?81EP;SNX[J(2_])C7SYQgVXK0gg9g
\f8[J3-VR@^Y,Y4J[MFfd8\-cKA0d)K4#]NWA6?EHB6]=R#U&G83V^3Ad4@A+A&S
V4aA[8Xb[(1-UF96Zc<Qb9J-SBI6;bC5R0J=G4d75Ud/b<f6Sg13VbR8QG;,T,8B
5NGTCd7a:\,OTRY9?,PZbe9aN&)aW9Y#aH221@FUOA6R>-,8M[=IKG>57LUUE3S<
g33/7V8MXeOLK?1KcYM[X_+SN_Ad3<9QP&\bF/MTT4)ZP7X/ES/H5cZ>IH[RA-X+
<;LdWg22.ZDSCFe]RRTSCdDVI<RX@,NN]EZ][2Q_Z.J_79(Z;KFJNR;cJG(N)cLJ
;W#=<]4T6@c>=g\-WSGZ3dO>Cb,@B4ADIFR?[_FBYVVO?gT]a_Y^\/Y8)]/_S&Lb
;4S-I,R_dCT8C:,bBEXSL[F7;dW.&3/[+Q(bc];Ja6:QXHA8/13aOLJIJ7\DbY;F
,QPT&#)L3^W/7YW:bQ]XW7T<AX,P.R<+_G>W?<S0D7VNR5gQDHdU4J#(dRWEFa.=
&/2T>\cR]=:?S(9G4.@R?;6VbUL(R=]-&MSH0CdeK1N4K]KA[g-?,5^QZ.H-bB+O
O).P,P6?NaR.cZ7;UW1(&Dd0PdK<C#\)TJL38K<-fe/CA2M05ePR&(ODQDf3b;CT
]Z>-/:7IKQF&@S+QXXP.eWC1L#X0gd_dWE]\C2b-cdXBIZPZg/75ZO42(X[P1]:M
GB/6NdCEa\gYg=_XZ9/ZY#9C6<f6>DB,C2#()_b=R+aF1):b)aXY/XM1-;Y@^Y0/
Ge0AJZ&Y(5Q]Ed5.CPXX)BML/AWW@>bA@,73gEYE5HW+X33AAOG(C[L/[1RAE]S>
KYZg(K4RTH[=E)F7QXgX7DQ2U2:0V@JVA1?.G+9;cgb^796-eV<CDZK/J(35e5.Y
Y[E22bD]^V34M;d:gY6#f8/g@OELV<DJZTb)ZA0DJ5_UZ=gIO[)KO)48a;N[L?FU
gee@3E+2BZIBK.@EQX3++HC)MR.+F@PX53[g8T2E1_^>=-_Wf/6CFgTf_>QT]dN]
UF0#[XJ(5Taag4aZA9fa=WZd\?I97=</P?F)S,^FLJ,CHNN2PSMegJ<5<O&\)5JC
>F0A.aLQ7[:M-]MX5PE^6bcgfV2-4VbF?BTJ545e8\D,4(@&,9IbYb:=GYH7DM>L
Z5f#V&-dH:eU?_F=4[ELgM+0<S\ebDaP>,fT29B/97OH,IYQG]+-,H]64\NP8Y.D
Vd,(PA(5-E3a^7W);Z+B<H0\WO>CF9J-gF/72@NX99bEaZ3(X)cU6GN+c1>2MKZ]
TK9[Jf=GKBdG:06<)C&FEgb42?:d,Ia<aO,I(K)\E=V?:,HFU/?Cc@g+ZY_<9JC4
ZVXGTHK1MFbSHWQXR3JSXY9M6b@Kf\@#X=Z;;^^LO63[IP@&FA<=4ZBWW<fJdQb8
NB<QNgMaVfHE6^[gGW19P<2OW76YINfE<<U&31=L#+/GBg]dC90O9,+J2.[Xb(-3
F9DdW03QB1N>a^X(8ZI_=3#E[-RKD\[-0(-X[PdO4:JRW8L9a#3T9REL:AI)FV+=
QFXIc0;a))AMYP;fKN95ZA:3#DET_7+A)#?ZEV5;,/(515O_?[X;/e2(/WAY-4\)
M?8T&M&W;3+EPe?g2QN?[KS8-J3R\E:1a[,ET\P5(6#EdFHSHT;@(9;7JTf/GJ@O
?8[\_B<&[6/VbC]H8^]O?QL9A^J)CHS(68F?_L3[E&Ldf._EL?U(G-.2M#(Zg982
(+?T_E#a)7](5cB49I/]-UEE?,70J9<>BK0JXDW:cD(7>eGDUd(6NA:9@@@dX>\N
2OF.E,.bP1J_(^TK<_+.P?QZAdgGBPI<7gScBO^AP_?A:S=QCYOB)/82Q13CIS<;
I2b>Tg+()L38g7KgF3H,cN5dOTP]70d(X+&,+4M&cK8R@e0^;8G<X2K;0ZAYNf7>
W3;/dc_/1QFc]-gWgQbZ>YX&W?1)YXPY+a\AJ#L6:P[S2M@bXW7^UI9P^.K\)K+4
XFBfKGIJ@E1TJ-Dag(I#M+/f^JJJQ6K9/fMYJNAg5-KP/b[A^YQW/F^GM1-bLFN[
Ea9Jg1:GcBXF<TT7fBgJ.+2JbP>2F4deg^JS4J,@/W/AgcWQA;23f],.B0.C[Q_J
?f:2OX^68[C>_9<F<V8#&^Y6Z[X_1P>XW3:c^>PVeU:)X>BS:UG,\6M#+U<F<5(T
<544D;M<eN&U/>+,K3W-Z,N52dMZL]c42@g3+6<OMg@\ZXdDb[N2U6LKX,;N./QC
-3_YY[L)&^H-P#D+T;Z))PH3JcA&C0JO((]eae#GHL>&U1T8->71<TT=X7,BW5AE
.M(2(WK8PC7d<g6A=Of&TL=P.\.IB5GD7.;6HR_@cR);\LP\#c(E^<S<aNg08#NS
]@]c[T:?bN]?SZ\RPc#8].[:U5<D365;W(^BBZI>2@MfYE8-87(>IF)5+L81\Q&g
Y\5-da+\8g&dF?WDe_6Z?><\\7K[2-]c9cbKB;/7^:1S,DU<Q=H\g051U31=_5f^
LaVY=NJ#9=7f-TO=P:R(cUe^B7BJ@=);d@#K/dYWS:e;@MTUCb^a(C).8CUc+&M+
7YVb\\(C/I4<KWbbNbBO-cXc1^b)X()4>[K95Pec_ZJ?(>XeB9.3^U+0I<9S<T3>
(5T,cOLM+=6(GQe#,233?a:.Cd)1Q-)Gf6#[Y97,B,S6)c)a[Z/G/H._Z=AIOM^O
&/)->G@VCK@L^@DK@XT-feed])TK7U_d^P)_Z3)BO1aG)_?;U_:M.HLJPTRV(N/_
ZfZFUB_@2K[,1415<Q_dUMfE_DZ60?e[aIN:]a4Z2,f.>PfO+8f?/5Y=VdbY>)=a
+<7AQ^_?<T?,J04IST&[/RG@QV6Ke9@/Oc[VB?-dJ32+fZ5/66+<]d=cC,[FS_\9
P2M1P1&ZS,(^-A,E(G80?af2KKX]IOeO:gBD7AW[g:]=d#dCM@UF/TGTg.BV3a-5
H5L6>N^aX_B)LGeZXR=2E.XM4H&94^92XZNJFV5:-K0HZQ/I.(#3OXS=L;]V-1SG
^Y&CX\dNbeE76IfP8X7W7KG2Z9G<-VU?G8A8gZIP3H)aH+f9+fUH+Z0V#-gZZC;^
,[E<(N&G+f&R/^_D(J7J^SaOE+-ZYgHZM#YRd@YZ-ae,ZT?@(KV(Xe-ER[1?U[3O
E<XN;H:/4^^T[Yb46Jc\fR9R)CV8(O\]c[W6c&a@-\FFY+B9+fJJ1Xd#[[MUGcKA
\+A24H-CJGKUKJ[FMG:Bde?QP^Q4c+CZ?SD2RBf;0KRL[7-c8b]4YC;aYQM_Nf/9
OT[F.W;4&VM1fe+^cGEW[G2V\,GH4_2c>VAXJ01B89B[_#]6QO(4fJBW9OaC/J^@
S>Y4cH,dN@6)L8.#HA\^4P]^=I,.:Ngf,d^(7/aNB.H?D/?P@PSd_5e@VF;WK-d+
2?-[ZF;eXS+SRKY_eea,B3QXS=Oga<RTcM3P\[8d2b8[99MCeX,+S/J&_1?R+Q),
M]L:F06(P^:e](_S\Ac9Bb#AbI22SMT4,VO/;_LZPK@C2ZVe);^=ZTcZ8c(fAgaI
TP0EgHQ0G=NPRQKYbcJ_gQZ(b#6Y58H\]3MZLIWJKK3:CR,+WS=]gI<#)A;,4GEP
RI>E]U5K-)dR+b08c92E@,^7@bB?SEI6d6+<7N2?U^M6bA>?)OTH8,P@_0+.Va>+
fE-@-+Qf.G.,7]?#aNf&>:5Z,#Ld8A1f)X7Y^QgH0RJ<N.Z&CP>d=VBeeJL-?@;c
D>RE4g456OJQAQ?X0IcMZ0A_-UEXW_[)8>6ZWY179gU<O1#Ha4I.0ZCSBJQ\WCTS
f564N[@^Q82?2&P_#/F+/JM#<.A6.6^SGS##EMK\Y[IIcM5L;(;&0d/>1W+0fNF=
]]E.Zf\a@ZAcM:3g5FIaFJQG9c3A@LU(Y5+.5F&W<0f<SQAgJJ9cVZZV:,?P\3L2
6dMM5<Q5SQgcX(PeJO)JXRKSdC8XS+?^c4Xg+O:[.-eLLYY1)]dLf/V0X;3UL=_c
e2??GPN\A?VdJIKE7GF)L^/OJZ&&J?OH7E@J<#Fg<@Z.#JA9XGcU^71U/Kde@dIB
#1DYU>U?U2VC:a[dG#\G#QQ90.WT)4W7);VKF?-Pe/YXQVfdT-1aa[48&>)g<R@I
VE;RL-47Sb5^(1[X3IC)f#5=?UZ^@:O_HHT-dCMTD5R1BUW?IY\Y.6JWH+AE0Ua#
U_B>BCFb^_M9?B4Ce,7&-_(JdT)>O]f#4.@,aMTM7fI5d])G\Q5=Q14>>,B0=71;
J?VO9\0FLVJ)K+Nd22Xc-U)M)MX;6FRO1^78MLC-.O;bS+6V(9J0:93Ud:c^-FHc
+f4C5M<7,bYN_>QQI5H6\9?dG#&=AKb7C0f,LV9[UGD5I[[1<A42TBe+]]T;.:eN
FX3Z/Y/e=bRGb=)B>W0H/SX\ISe->WT1HBbR_C)Kg,0<CF1Ca>LK671,c6==DS>:
E/c2OS924OTD_V;@Lg52:-]9V;E(;82H&&Qb^cFGU(&e#WXOL?gQBOB+A1Z\:<bB
UMPf^K.4G:[a\gMOH)##U+bH]1[<_1(\Gf;>c6BZgS=bQC&Y2Bd#82+_2IC;7@+T
997#Z&Qec_>NHMgB4S,<4IWWE6G=XN6gACZf_C4#5S3V\)b;+WY_O<IU(B3aZ/<R
g0bddZ\c+BW<B.E:XT04+)VdJ?VPgG-QJKaJ6UBHR^;^dN]6(N5U&Bf=X5DP:_=L
M;RG6[HA=/C>bP0;.gU&KJXd(7aMAXDJKG5K:VT@3^GY0199=-\OCeY4e+?8[\JB
fbR4gE6/(-:X7,J?.agIIU=3eZDH5BTURIM(PHG&L#a[9<37^^)Y&UDQF0])X2L(
DALAEceW/T0N(gDWf3]IYJbC);D3bg2H9a2b3AD\-8c-3>WT2e<+#&UFb)B[L\e>
GQ/WP8A-BcRU\WA32;b3ICN?L\/E=@d9BX_2[Y8&;)@.;6.0M(BARN\\5LQeW4)g
\^7^eK>K+P[D28S/;8P_R-Q_>S[U9@,@2#)AGd:cb/0)b,1GSg>T3PM1(=8<L:/g
#IbCY0E29Yg3fGdV:DXA=,[\Aa#?=GbJO8Zfe?\P;\Z,NK+K<<FQV(4M=>&cW@+A
=_N6B6b>IH43+I7+XE@X7Y^;BOee<_G<7cH4d\<a3-GgWKV^8]1La#Y&Ba:IW(MU
G^.>b]eO-<<Pbf^dSPaB_5<eR/,W@=]ccJ7\A&Jb7IL>[&e.U8c.(-bT[b96F/>7
_Z1]_.(f_]612;BW4G8]^<ZaO[\.,4VL>#,OD7FOe.B-&)baM84;]&)W,SL[0NAg
ZE3XLK(@=AH([[H#4bZ(4d1]EeJCOU5US(TTSUA2:]Jd6EN]U\#_g+30RS@[Q,Hc
bFCA(RK]E7RSeEY_?>-Kc#7;7fGa@59O>TP8).),?TY\JA#dJWO=N4F/4HP_7B2J
&[Ae/5NC+/A/BWWZg5e)ZKR3g3^GDJV-6f?8CJ91//NQLR=S+UJeaT[3Ib.b<I>A
2G_Y(@]KBC)?4/NXS:W:.7.H&b(]U;;(eJKeS#,O(:B7G>Ed@gLOZWQ.6QE8X(W<
?F;_Q)?9,##82,K>M[,,34H#c[6:)BV18ML2daN3\DP)::L8X=BPYS8WST0#Q<L#
&FAC2Eg#OJ6a>F3@OePG5<MO2)W[V]gFJ=0PRC)F^M07PM^?X_N(TR:]>2WVc//B
LSM,cE_ZGZGS;c7MJ^G?=(dA+2O1^L;W:FPX(_bKW4VFMca.M+4:/]ADUcgJ8_+9
+HbZ,I,UJg6EFKRN/NJR9ad4A9^=7a,?LdXKbN:#,f+RO4d^>WX=:\&UIAR&[G5W
FJ&9DP9;e0YIMee.XPUO^3H6I[0_/Tb+HE]QPNCLE4GK?g4CKFPA;?O4BQCe7T,E
^)+XO(M1##MVNa0Z^QA7+^/YLb][>@CD(SIB8BXA#0aC_EcXF2-JWbG6O8I+<4D;
ETc9H7N)cY1aTI&2]aDLSTI9]E?\6>Ngfc@/-G=e-TZ3ZfdMSZ=3;fA5RG,SC^.)
H=g\U6J_DWGZ.JedC+)GZ?-)Z?(N@=/,a@4J(Ne;cAXJ:3Pe#&;2-D:EFW+7+XQT
a,,KY0<S^ASIQ??71@PaHBOF(O\J^=Ne51]O?L64U,4582afbdc=b>Z>76143)TL
_RB..gO?\XZ=d#dQP<a]\).@4)7K;91(6G7c_OSZ6-ILRO;bB.,X0VBX=9FL5RO[
B<RK#5,bVG,Q]3ZSdK:/0EE0(VQ\,Z.FLeL9.51P2N@bLVB^8XZ<:4FIF^@bQc0Q
]H2e61E#LY:B2U7_B:?1KKa^QQ&;1P-[,6,H[H#d#]&(0>&YF-#dEcJP50\=Ef)U
5=GT\M;-Q[?\dD^#f;6XV[.#=b)&A@?[Of\+O5I+V6&Z#:)WZ&(UNIA[Ld\Q3W;_
ADb33NM7FHC+2ae(X7M>g2;4M(^fTD(\C;fD<c:[<>@2)HP2]0<N6O&_/N4FEQF=
7=1ZF)(<TP4]G/_.Ob5b4^#JGc?:/04/M)g6BUL/YDLXQ<N^9Y[&(3NPZO6X8C]X
4&-W1>]W3-Va4[LI6gEUEbB[M:+[;R\^g0H4BZ5KP9Sg7B>PWB@+#:d?0_+JTcFX
=FMIG_;AJR1U]U^/d\eVY#,]4Q8B=)-bVg\CQ1DN,<3b1DX-Y9^BaTefH_2C9#<3
<ff&>WFEL];QeVdF_G#I3]_Da?OY@YPdCY9TC&JE@D_WHHHbT+B3;(H8I5S3&,L>
NYH<<P:/a@IeYZ,:YKMKZcCegNJ=cL[g_7]gD^:HAXK3W)]g[N&HVfAUJb0<]Ee;
bZLICeAD3KNJ.Gc[SaJ>1bVfY2@GGRA\0;Y_4B-.#0P7RgJ#;1^a(#;+.AfH940O
0]Q,X()A6bG_\A=VOfM;gPAP5P[8\?\ZP0Q)3C;,=C&Q4e<(7Y1+BBf<X-:^VK[-
[LV2>(4b[&.-aF\M-Y[fLeRO<7EC.&]^^6?SWcC)AgJ3?8)aRD&HKM@#U,MgT;#D
5LY+\<0LaQFCA=H1Uc&Z2^8\^?]>IIc\>O22^^[O/Y<SS:I=3e1^MMb#<:9Oe?c5
CZZ_/:g8E[V32Bc_.+,0WV<9N>#V_g(7E<<?\[;=91,,8:K^b6#QH-eY5QVM&^Q+
CIf-OL7:E=6U6V;OZbDI>bC^6SYL(=<4-c3@-1SfW\604:8JTd4BgLX4gb_:PS_?
#\\<3JC,<]bC;>cK6,<YNg((XU\.9;FX\+)&6.<75=/1-?T+aVV=79e+P>#4V-K0
VKa,YP;1OJ:>+T3+V(PY+S]0<0H7&a\Dd?\KC\/4Z86S^eMZXH5f>4&AVC7MW6VP
4QI5.<87+@-1#8b4UAC_>B)QCe9XEA)G[/ZFU_RJe5@1&7^Ee?;C76N,&U\8YcT1
V^R>#HQGPe<Qa/6c(29X(JSRN^gM@d1aD-F8R[D6>JYWDfX=O;.[Ie>^[g.;Q06&
ICX2Me=8?^\R;5A^GP)/L7.BeOOg,7^(Y\7#.e03]S-)e/KVR6\O(P?AU4&1UIR\
YXRG\dX&,OLT0YM-4ec@?L]7ST9;+=0B#+^AeGB=4)V)McVQ\I,&K(KXYWB;WL0,
UT&NVQ:2(fUN.B\/L:NI[MUg-RFZ9OO;)C=/IAKD)U9dXK21#&^/UJ#,#@]3O;J[
J]e;@5K-S0V[7I?]W^R-??>>?&H)/<;S5G5&CANOE@-)H8dSfX^I6aNMRS?M+80;
fYZMJ8D#aN=S#e:U8EASYUJK61\&4e[,02TC?GB=4AP@R+@B_#^FQ2M5I0Z5T/PY
+#Z)DKHWI-9WMT+,[A/EH;a/6G-OZ>[KK+9bVK9]]VQ@H>H4#6]34Zd@R:^Q2)eR
(8(:VLN#+cTE724=a,V#VZHJN[aI;3+)L[S-a=@BRY3J>41&,JYfIDAR:3eBC2cK
X06ZJJ;]RgC>3,=-)Vd?g4T08(PKM_,BJ2dBX)[VDa3Y\0cXQg))ACZATcC\QL=[
X1FQf;d[@MW)[ECX)^A:GG8Y<e9>;8WcYEGDd=5A9DV_:.,>#;J&>F^E.ec7Nf)[
9R7+>WISN0X?N4MA@7A<AJd.@]]N(G[XUZ0AX81J])]4(D9bQ(BB_+a+G(\:Wg,f
0Pfg#a;]R5A7bZLbE\DSTPG,c<O:cG8<I+;SK)Rd_)(3I26@bTQ[KY^3>(_NQ<H<
B._GMXR5cfTDMJ=?_bU5RD71IgDS.LeG9D[H50^9e^-/Y?&/M1Mba9I;gU+#c2/Z
UN3],XdB4-]3=/F26KD_RZ8I,0:?SHEeK169.H0JVFBLC75Id6/L@bZ#)1e7>WZ@
:-&OMacPMF7#/c#4\#FB.Q<S4YXfMHZ0O[C]e6GaVf]>&,/-gX>DLZG>^Kd:P4U?
I0@TU_7<dM#IPDf>fV8[9U.TNCZ)BTS]A-5\0gZ^7cSHB[[#Bc(>G8^&QM0]E<#5
7I2E2E[,d9IBW5WQKJ5a6M[-IVR0Rg^ZG-B^44;:3H/f)]C.WMGA-4]&].W+Ma\(
Dd[?[N</GS6:JDBEV3\K1T0WW]KS@c3X/\(25dJA>3.d7TKfd5/,FN>:#U(:7]WP
]E/<Zd+R_5=,+>;EG6U4<U-agEXCH,70QSRK/QIXBd<=[\=JO+KDL6UEa.Y3R[6)
89QLb^7RaEO9WHWVFXV:N8]),79HbYBR+\ERO@efT-NPPcBbYD12//DX48+fDg.,
V?2]N/WF[=fLMQ0,3^E19#4Q:BKHLZ6NF/>Vf(>U.]5C/\X=8F;?a53d#A3E4D7D
/e6K3_\#K6dTI=LAOU&:\1<-S\+g[F:IZ(c]a3VNfCCZc9Q1BA&-Y:5;J10+6)^O
Z/J]2ADY8C7Y562WfgFHVLY:UZGM=16K,S2G2YSBF]T[VeRE61-ZTCCXgLMDJ\Ec
bY@G1\eFeTBTM0OJQ]gTIIWU8X0K?V>6LGH)<Z<@I\QZF72F@dI88A)RU4GVL?Qd
5BR3FU-cENICIBY-7]A73)+1]8KDe:7c<0KMaL[)R:^EaHE2a)9P.ZG+OVO:LJgS
3,^GFLG:(^7#.KD:S\cEdURWMCZF]C2IJ-GVAR#W74WeP,+Y0ELS4(Ia_ZIZG;gG
,JVVOSU^[<;J+cF7Lc30CS/.HR^SK^]Yc+45gKWH6^.4d^G@]@JY73g^J\FZ3F<#
a[[@E:>HYV/b7MDf6()FXE9(@D5-7[XJ]<LW2URWTA>@IQa_5H]&c&S2FMRC@KAZ
3EUAQ@g^B&5(;PSB)&@AWRdZ6>+Jf?_RJI?W:DXWgX;14:[FY7[K0VYWQcCWV=dD
E6JM26?Zd18L[ZdRc12+^Nf&F(&=cPK]39eQ6E<&LJ-9DJ60RPV3?7-B_A.W)3@<
D:bd-fLfXb.dUES.e#(02G_UWG2\[5?4#\SSeB&&KP=Ae+VW9^TQEXe[ROZB;6<c
G#W=f81A]b#6N)A>SD+0UC0R@35,>YYI^-:g6NPM^31P5N5-=^@/2EP8;gPYEab_
BMCTP#S>-IJ85G\@9K;^77[W_6?ODYT=S=#BKO.-I2e7RHIf;:D/N,.(DVSKD/RA
bJ5c+/7H/3HIGA_@Vf92FE)8Qa(>SfDV,)gO0ULI4QdbV7KgFg:7aPP>KQgEIBL-
IJ<JUT3V/-2#CX#=G7)#GI[baf)ADVT?MYOAF?AK-9ESX(+eZK@@#U:CP:QGdZaM
#V:H7,2J_?YaCHI)W.JJO;[D+9#6MX\c?@6L2P+,V&?LNG^VUIZWXO,\BK@\9I/]
8KW@FCN^7)=ZZaI,dZKP:c_>@8-Q)]gC=?;1_MJH5WZU;;9V?1W:V8/++[g1<EFe
T>;HBU&(b7>-:G&a)=PK]UF)KFX:J.GY);&S[1B@G^:eK0[)-/10_^f@SM,D?0?D
LJVB(HV4K?98GJ5KB^<Tb[&KTH&11BT,/[U4\\<+-4H[IL>^Xe,X[?FNIOXL.3/6
9L(@#_ZS:?NdcOL+&3CN=S>ZK<:GTFN+FY/3[IVM9L&B92eRG\ga^gdY-df2/K5M
:WIIN7?QR/LBBWC5+(6W12OHC&QZ)a37QEQSBfSLebDL4\,?Tc+TB5_MD4PM6b2e
:^fX=[PE(_I3(2XOLIdA5]HF=fQ&(FBM8N2PZYRe(Z#Tc:7(RcRFIdJ[VS6GIVRC
:#Y21SHL1SJVD1eMbB,S\@gGY:H8T[#S.,1\RBO#c91JKKcN6[3-_JV>a52GdH1?
NbYY5#+5@0&80d_Rf:b4fGT2T&a1Y_DF.O@RJ,[)B=AVgMa.[11:WK^,R@G2g4a(
G[a&ZDJIc4AP8dO0PLA8=Kc46Id3I1UGdN@N21FF7.fNQK@a-NZ:I#QdX(,MX99X
OWA9@DKb8WLW4eGMYIE[OOI>gYU1N<f#\1V#^Lf1C5ULWB,=:T;?E<NDa2@\<4M4
,D?(N/:@&X([eb17@^Q>(PSeggf2HO:&J@Z-OX?,Pe#J,3G?)H8-@-=53)JC:aG+
7cWBM4K(Z+C.L+CJS]@X<&K1SRMafAFW(f[8c]B7XgUXC6f@<]R:3<+a<^K+(:ZZ
:X?<eL#.#AMdSV^_B0UYe]3.:_GEP#8X^X8FIG.65W6QQL+O_UJW240RXV+=H>;]
;^eRVM(fKK_RA;@_<XRHE,O6)QQ+B;-TKTa&D25]27cXcMX98Bb5\#JK;?)?F^,.
RPa&(:af@?<a>ADd+IY84K@:\Y3I+S]#D;??BSXEV=OZ>0&R>fNY/@_];GgH=P6(
IY)[NG.O^:M_^7@#T<>,2eG>cSK77?X46fUV/)\e\NO.T\YX=U_LA/&1,3+ebdDe
4VJ5Z1N3D9[?Q;b>I6PYYMD+68d_AYc+V2,&2A3D/&-3O\9<b.=LH)NNJgKF#J<5
\3W+C)\1@0B6P042WQ?(Hag<#VV)FV+\+JL:fHBPQ8Yf4U[eY:baZYE9.1(a#?(+
gg&c@NCXGU<RRO)MR.#,MSAI/J(5Q;VCGX(4J1f);c2PS[e^2IG(RMVHP.]/&6Ue
F,KWB?]ID5,Bf7NDDVK5DgGRUNQP5acQ#/+M&>?CIIdR:3cbaU-.H(;?_Ge?TJ#3
_T./2GF5JJbP=-.LP<K-BaK.9HI272Se099=.b#50aPRP@HN&d;a\UUO-=1,T]Z>
.M578&V-WO3a:DDdDV2F(J77D/c+RPda;LT-L,]:(L_:D#A._QYE#42W-=GVE8a@
3g.a3BY^7.,K?.A.V[\O/K<0-;&0IJe.VEYVgf;;5M)AZ\NZTef:f;05W+@H7N/>
Q6Fc(/0fd<SSD-B-fYdG/NV0E3_40CKKVBH@aG&-^7F6P/SE4LdM52PdKcV3&V+D
DV#-1eY^5\e.&9VBXDK@D92^A84BGF&HV]c,S]4Rg8bN/3_fKZ7aLZ,JZS0?.:J:
TYM?,/0#(9FNL-&47&\]A:Wd]\)I\I@S2AcR-UP&:_H:-Lg,g4b^E63/EVYQ+_f0
5?8N<4&8aAW3(EgN/R70?H]?a(OVRd>/9dE017>a_N:fMfc4e2NO@J2Aac-ccUP9
FB?RA-.<#.,f1,,3NV5&]IQ[1N(00:Y6eHa0MfR3QCO8-Q;K,5/ZW(_>L@9&^YJ_
T+W<PTXHLY2-?BN[XXF^Gc+W3EM=#=6TB8(M:I^dQ3212e(8;C6(>8dX1+If<;Q[
6I9;_>7E);._Y+].7X,FBU6_W-^M8c:57DgJZ=GU/(PE8P.:VA;EJU(X6f].B/:5
X#^]5?6Y3&+DSQ?_?dfX^Y,Vge2KT(8e-UI^g[ST8Y(KeA.;S-UWZ7d.0XNSe[3;
ESB^WfS(3M#O</R>4W_R2IWA,\[J6DPU5&fU<+N[f)AB,c2E2D)=>-2RWS5#9eG#
OJ;Wb>O8R3c7ZG2@>&HSNTC-L4D][GPU^^C6Ja&d?ZXg[]W1K,#-)F2^dNf\1X0<
K[g1A2e(&;6dBRZOPe50R<M3E:7c4/De_2W8)N?^9I/B;;B<b]#0T,fc_E-XK1J]
;J#,I[147X26bA:I<a538(/6V+I3a@JA/6-7R_=\FD#=K]6444;/(E)7#^3)eO]?
B/>]f0PAXV8J;&eLfdYK6&58PL1]1+LgHC(.EQI;FAHd?C^FK4K(b##WdII9b/X(
AA@aBY_bFcW.b6+0Ca?BQTPfCfJaOCZc6/1a:c;X_]#ccd7(6<4bKWT(e(9^NHe2
?O3X<6S#88TP+U?GQD>^7]VeH=M0Z74E47B8SIY8-A(&#,5O4M75N=KL+W_?+_4V
00^W^YACd@P2/MTKJ5#3O)O;4WTDW,a006ZO]N-CJCLeLN6-,USS:)F_S]OR]g^)
d?@XD:8<b\QEVI/N.)6V7ZO1H5#V(P8-bDV&(:\\7\HYe;/D>G^D&-@\+[C&#WP/
8-#gU+1Fe6F;c7F8.>X]b:B_06]Ob>QTa)0(;QH58dH)E&ZY;A31cg0:D#EAAf5S
\P9Q^36D=YPaF@-b5P.L7NVMIU)Pb,ZZ?<CKH8H837/^,6I^CSDC0XAC]\]GZ@:F
W123dBd+/9#NTH&:(DD\\^QQ[?bX]@1NP,NG9^\D@;F@NI[.<I&Sc>e.Fc]O#W=M
4(&fLL_WfS&I\I?BIF:4AM&)cZ5aI(9N7Z4,\EfDVV?:H-CEMg4egaaa,)&ZN6[/
b?ASJdda->,T(?(8KfIG<HN1909\d2V@,cY0T7L2H=g)5YbXL^DFHII1EF;I08Y3
(.RCdcGZ:aPTWb\_9K[BeXT#OOcW_37B/d8+E(-^@P7aa?I)SF[X>0O&+&AAL<+)
Z+]7RP-?6;OTR.XLE;85^[^QCVGgLHV9cDXHN)NR6,H6(+-U_a\F9EDfA_3:aZ&,
I2BZ0<1=?+;fZ-a@\[]JOKB5/e0Vd><CP[Z;J4T:((3NO:Y?/..5N2;[LR&M2>K5
BK_1a]71AZLS+9Ab;NMW2DfK^9:L\X)+f@cRf6<c5<D<M[8ZT0WX#NGPW(g&d.XJ
W/dQfOKCR>g=)PU,@(,S1BA2b/7]^SJ((:&TJ[FUF)&VK)(5+XUgg3H:g2[2XL)9
1_@F1FW,5e5aQ/P1eGC.B.IaL#97(8g/WaP89=SG:3>31SJSZ<]e1b\R[T@gU/^5
44dL3/3<7Jc5BOUM<cQ3H7T<JXT>)UVb6R?[6:62-8Z\e;O)XDH+EW#Y>+ZbANLO
89(8_dcFU_A,P.+#W2GR92>52;VJf[/[99+&+=9Z6M62&MNDa[S.DYB>CE#&5Yf1
93e0HD7IO>0=FOfb5(f#)g[]J>P6SO@M/S.EbH=]c39GRTdb&X&]^bcPJYF&X&>H
dXQ/3RSU.e-NTLLNF,X5^C]?[QMOOfUcc<eTA=BJbf=F21:,UNX<27SAg^\Dg5/b
XW?g)O/B4+/812RN]_QKA.,X\VDG6W+6dGVI(8,VU6LG5C-\1OHVD+R@L=^#7\5B
_&9E?13Q3L-4f#g<H.X/[VTI_(HI5^bU.B]0U@:7P46Sa3[6RV^cXXWf?(F:9P2Z
a(&X3IH^T>@[PM[F#\1&a,/PbW&SH,Q,BG.7SEPZ-:GLJgf@,C[CDFH.4>#>X(b4
8_6PEL:9BgMd.07[B5DK+=I,?g4QeT]B78Z&P?W]X9XV3cN>+@/=U;H1?:FP;IJ^
(/f6Hc@OG?UKXd.KRT:bLDGcNM_R[g6T+EZ48.OY--Y-g5N/Z1O?b2(ZIX46WTHZ
(7cUV>Y\)GB:cDfGUD7fUQ1&Ob7P+3(M<N)EYN^@dd;]REWFM#YL^eA5QB(e-@.E
CX7F^G^B6He4CD/28/.ON2UUF/?(8OVW@#9Ufc56D1ZcdD4:01K&@DBQ7W#2a?T>
0UUGGN_3F^fEK7GP7JAW\;P=8F1]@D?=eLND4.U_MWGf&aW;J1cWEaU:U)&P?#9C
K=:SCI3McN2[/_d6CUf@JR3=Ja@9cbCgb#/L)RD7/6=@5D+H.A;LNMJ\d8.>S+((
XZG1>=Df#agOQH@c^R02dZU\ZXO5Z6Fc[8\A+YEC<[\:0):D6<[;M&39+(b)ad0_
Dg2:AF?4Q6\[RP^IN3E]f^fN4/]A)EG(QJ8TYO^QW/G7/;U(+H10H]=(=P@-249<
d]Q4WV@#PAPT3U0@e]P?+BGV3C(DN8Aa;Td9X1>D9=J7,FRRYX@[?L[MGJaBG@Fd
N@_?Nd\PC-HJP1.+JWf>N,);P+aI)3>/F=\dZIaMaENYFN?]^9<#X?4N6@&A#:/f
ZW]cSG2OX8591N>]>1a9MaD6K)=fJ-]/O_>6&O3>191)VEaEY6R)VJcGOB7WaT>1
5gZYP@;a(+ZdBN#-NHOH^;G,(fU?6>G;9gH2ZA9cEZZ]/^<@O9#L?WE.2fdU<2Y9
,/5RS)^[A[d7#-U+8L3)+,#]M/TZ:+>F6-Rga).G48e^SgcS46U[A(7XbFJ&:V.S
gF,9JE)L6RBc5YPP]3KACZ;6Qb7e7YVW?\F4ZA(aR3NRZ3McF0G8O>=a>:Za.eb=
+PRV9T?SDaY;LOB8D8OCV0J7/3L2ZJTSeT?9cF<-Cf?<H(4Y-RdZA#NI9CN8Y2PJ
C47#LWEBOB9YW7IBL,+&;[WE0K)PaPeVbMQPE8a_cBc]QR^@MARbgZT/;_I228:[
@#Q[[EM=/-2/aY?;)?c1OP<B]D:GY@]LYY.1,e1=SSafOO&7,H#[VUX^:[\#0B<+
_)JC^M4N\LK^#KXF93H>ZPE-cYO\,:U-7K#adB@JAf0OU5Q:I^:488LH>&Vg3g:Z
.;<#W#gYF:U)f[JeLgQ&A0A,APXD_edH2PD6>TbP&5(<D<Z418cF70+Pg23;0\]4
9CAc;5Q[C9g;],LT;#4?-N5Z9+e7SgVNcKgNEW=\bZ)K=G\/.dT^R++d2eSgG#;g
(bHL;Ja+=:/OBEAcX[R?=g&/>\\,062ON4TENYQW_5UcUNT#BN6G-YdC+IRWTc9W
]S:(^JgUNQ-+=V\9;,fKa,6XaMK]gM=OH6AQcfO8<5/+&K<1.LLQR=5H^4^YK2@I
86P0[Bb2NG/:dT7ZBdA]gG^?.]DLWRZ8,PN#?3B94EA0Sd>O]ceDI7D;8#;Hb+H/
9BFR9+<,,dP&C]ZTMCSVg,PECLe7,5^&E-EJ[^KX[X@f+1,]C:E@G;/&g1@FaZQL
-=D>CHD/ZRbe&EA=KVF=fW>af:HI5S-8_Y_HPL:J2-V_O.dK:[=HE4I-9+,O\/@a
aT>P/+@[Hed,L6VRK;Be00MGT+cf,DG;>KS-U7OS/]#6F63UKNJVbb6@@\f:;db&
A:/P..2A=(,7GN#]W#g,VWHRS;:N&&;[&/^ZT\Q8);U:WN8_&a>#GWg,?=<S=\7\
d_?)@_fXaD?(=VYYIY^eLbX6_a:P;-NOC(BIE.c9g?B,;WLITdVLJ?,6e_Y8\96]
H<,8^,[L351@VXUWT[Ha;9?K@K6XgRDV)));_.I&0),b0@GfUNf.4PH5+;A#6^TC
,g9B5eS)bd]3[bBTIC@JB&)WF;a8@,gP0<PCNd//9RW7B/e[\73H;3eb13D=>(J/
P:=4E19c]IH8^26Ea)HVR?83\(:>_ea7ZS<WUIO&e@eMIXP^9G#D/5C,.N/(7:J#
#53BIba(EI0MAR<I[Y<Lf&4=>;dV7_#EAc//G^U3YN5[?5.2BbIW/K/-bYe7/F&-
E@\=WA?)+/PT()D=>aL@bK4,RL11VJ^>e5_E][bYLB&.]=&.F@0L^I+R0H79TN=K
A&5^1/M6cgL))<+J]GRU[A2c3H:=.E\DM#eED2:_I;80#M=CT0[OPMUbYd9=#]N4
2T&Ga(I)-]RXA\CX0XN.Gc?Q.3ZCdA\E45T#3D]RQQd#M/e^;()N:A8R:Z>6LecS
J-GI;4QaM>6XM/F(b3UXa#<Cce]<eFRe-&Mbg=9D[7\dVOH-5+gY0]_-1#TY-0R)
IF;^1XcZ030K[G924.)MZIP+f_+8DLJ)&B4DTddZQ,=5&KgU.^^1g[CMHa[R:7&9
XVLbA)L-NHC)dcEVO=1AF9]#=\J+MeeAR,99G8f:A,(;aNa).-GQ>,^5dP-+)<9&
#1_-C=cV6&_]BJD7]?8/4B+H8/+XRf,2@O0,POaT876B1^\)a2,36(d<H-_>E3)1
^R&(JOg0#AJ1NJ?CMB79DI#<G4UHUP?I5d?+6<Z=be?eK->>UAb/ef\G^7KB:&T4
a320gf[Yf1AHZ\e=5S5@:_c]##EHSG@NB9B]HTfM4Jc)KZEab1@>LW7^?E:YBO;;
&KIHB#30[?A+eN3;MDg2aLKPG3-3P3TZ.9I):(ag3ggX9YRg5WKaY@;931029TE1
5Xf]Y^GM>LKXY#485&HB87BJ448_aW?D>/eN@1=cI0]WY(J?\22IgT^/TJNF<MGf
UbM8&0VIS?Da0HK4B#6^?b>&,OJX<51JC^K9SALNMTM3A891a\a3Ae@eWNF[FB-M
7^][/A3BS+)?ZO&JYPRI@#JK.X>^FaM;]&6]N@b4]1S1T&PK:-7.G+HK#-f,.YWA
83WWZ0W^baedW6FFb)EfXUKC#Y=7^T=^.]F]2O1B<ARD]X7AT:\R3WLX4?E:9K1W
?B1L\OF-SN;9/J>f5]=OO8VSaMdVP6d_d8#Y4Ta.bG+5AJRgN\R?_T)8>f8NMDM.
D<>--HL41<<<3+T3(I>,KY4Y_=6_IG&B^ZSC9Je_W=b._YLMQ.WMSYHTX7BM00D]
41Bd@X<=W]>+L?MgT4-RUW.:8,;K:(652JKD1OIgM_4eaR2^Y&cMfL^SVa=<RgL/
)X&]e;KX;4gG8d-XVVX&_C^R^)?R))(()c=[GMI/W#1-L>^/4g3SKU6+YZ3?[&dd
-)N+FWAYD;&<f?X3K9WDDbX.J)2:6SL5#F]S;A[P.cEH>D:[2a>)[d/@f2bA^25f
BWL5b+-ag5399B;FYYP.db0>./+)I:0EdCVNO3N5Z+-O/d3UY9W5BW&0=fSG.gJ_
)U<DLW^V4c/<NUD]R5)CO6ZB.?^Z>#OO>YEg0:;-WYH[DS-JEa<JZ?Y8D,DBT.S#
8-FB)0GOQ.#9<\+cbDLB;Bd>QDeL5[GT3,XU_IL(&#_J4-+.&7a\49)=aWJB<AO(
IRO([HFO,;BK;AQ;Nca&JJ6G0V7Xg7=8(E)8JN[\4,#TX2<JD2IbB[C4@ggIJ@+&
-AXS30SK=FHafF?>&A<BaMRL<BcC4Z)JGa5X,+&7E@R,g;_4A1Q7GWBY>H,+<ZbO
8JHFXY@#ZS&7E@:T(K]Md36:Uc8C)cgLfJLLM1@=[Q&F.7;+_C6fbfJ<Ze,\]8cX
E=^eg^#6GU7,)O.1#L^5P<d<6<QdNQT\bT>g?<QdP&0+-HBAAY?b(H[^:1+TQV-K
)F-C3A&/^>PI@Za+;9e25[@YgUY@;\HgTNdYWQ^6V&8+AFVM:G?23KMPJ,#/P97[
7NFdA;7?TU[+L4a>X7CZ)ge<D6++V2V=Ra()==RYQNYaEYb[JTBCJS2X3],4NM_Q
O:^KaN:1^E8G_^Nb?CT522Y9M4HKWB,+W?>OFLZXA&QE,G\5XbgAgge,CdKE[Q0e
7+_UED0dPV#WbJXD7.bX0297ZBQB?.[+PIEeH2b_X0Z.DGC\VfD(WXGS\S@cgNK.
9\R9,V:6T)JU(7,G/IcLVaDTLO>[R,#O738D2f/bgL(gNF8V7M[c[3,=)<M3C#[8
IP0)Le1E(9bbe)B^[\YH?PB.df0b&&3gL;9eePc3GfdRC]4>[Y+67H8>a9dPTX9:
CfgB_e27CgcU(]FZ6QC^UA0X)G,HLF(#f0^6I,Bga^U6)KN6;YF/Mb)g]-S/)PNI
4,3SHT#JZ5QQ<X1S50CgBT_[Y6V36,e^f(J((KGQE+-L2IG8<UCJLT;&[,@P_c]-
[4d)V<M=ZgV8M3M18#2dH,)E_2L7WUf;BNFea,8T[SK202Q[[4\@+31\geXO#=_7
/(Q9((#QFdc^)@:5VVK=aNa9##WXCFO=?/^<7,)C^KYBeC[A@YX?cG(2Z;(R1WP)
1H+CJ>Y9b_I)>J.H[Q)]N.#Ged1d[c<XZ#_g1?5dAF;=G007/;L8WY/bUZ90daXA
fV\c>J:FG>8N,-BJ&?S9OC>1_5HU0.+3WL\<dFQ^#7?cdDG2;VZK=ab_<>d.HDKO
dWL(,-CcMW;UIO?O,3a/0U8DWLd/F_Y2,S(YYI0D5RPWJD41]O?ZMGOf+ZY9014E
=FK;/7UK6NC<3XNce^WC9LVMZ?,1]F93G-PaE8:OL&0I<d6fM-+N:R\&EG.>(a1#
<TFRU<O[LZP7,.9>]AZcU;Ub1g3\VNKTd3PU,7)U:3;Y3gZcSbQS+^.]VBD46+c&
8B<HEY.0aa3@YH<UX;YD=X/4E-Gg6TV;/725@U^<9[EbG&4#L^0YVF@)[9.))_dU
^4H.V31D&T6X_L]S7D]?=WeBgR\C-(YC]@^Wd6#LbIK4S5R<fDINF+2MCK(/5Za9
V>:#L[&_E8T6V?Fa9@Ta,K1e9H^gA#bF-#N1g#\H^D1R107fIL[Cb_0Q/)X2bX?g
\Ve9JB_?1?CD,&N>ZN+KPLC^0NE1a/OG-F.gR,HM)7N6RH\F9CF=EE[T)@b\4B0Z
?e:]/L4-/,MBc5=C2B+AJcIP-T(][:XdcHdGM=M/Y=\D>ZUb7Ia]7Q^PYSP,R40S
=b)S>FU/RG,bN,OK[<+O0NG==1S<U6C[&::bV@JM^7XH+=X:9^;]Ze-J]>bFc)DI
PCCG0c1)T+_9K3L@&:#Zf&\6,_W+CL4S<,,C<S^H7J\K[G9KL?/HMBCZFg7[5.SZ
Z4K]-b&T<Z>60BU:/;F4>dK3BXGNMb355IL+F8D4a8O2XA.++G7(23+E;(KA(W]3
M2Z[VIYc3.SfGQ1_0,I^GY@[<.2D>W(<&YD@TT__Z&WRB4\^RQ^C2E_@:@40b)&b
@5\?.CF<33GNcdA28X4E7UU(/6UaFQ::L>a?HT9:]K.>_8HbKKT1JP.P;]6AI02W
?2_U^V8;<&MZNB39aFFB-cV95L<Gdb35?XNZ4=^U)b=28?Pe=g0a>5&;b-]_cNd9
+8=4Q\LG;<N20719VCOJF<L^Od&88A_TL\TSX8J+6ZXIdI#+Z7Nd6U63CPX8__4d
PD>;FTB@VbQG/^18EbVII5.+bed0G37.)8g763b&?-8,G/5_7MKg9O-[UDAfF)#8
0_;.VJ9XR/O(#7[,9TZ=@.41]?@)#fNHKI0V^NV2AUaJ@]G<d#J^H&9X82<UT+R3
JF#M(Z;=b^C?:,QJ],IAM8UAa3IHF-@?HaJ.2MfadJM.B=(\c-B<[YU^HP_Yd]56
3I.V],0F_HLPc31O6aYWS15@A@@F1g:^,0?cc5[?LX#XG]^<00\J)904>g;VdHcS
_;45<J^;7EKID6dAa<_[H+WWI_:?<&U5NTbRbH;OEYWg1??=ODGCMKLTRIJ\DHE2
VM<T7L^R4S?^&6^g&2S3U00UX+dG.M^a@LVecW2L28MN-e[fb:9]6DLZc[MFIYcc
MFa(P4cPf(K]5EQ&T?3-U=E3SeBg5(&UHg0[d>3)g^;)B/aAF@?K[8C9\?T\;0H8
(&(TL0-PHa[\#,>U03O;O0&DH:G?./a&0f\HbfK0dSZ(DN-0C.U>J3?>3:^;H4Te
=SeF:@N9BfC#H;SM8F&L\L0N3IK^V\2I+NI;d;V,[Mc>L)^3TP43BD\SQ3@R?bCS
Ng[QD5Q?>-UKGcSe4@IGS2._&I[^(\Jg5RJRg[K=U_OMIX,7,3g3aT@e?<\,G@T1
#U2Vdf7PT^T<V+>8b,A<6)S93)d^RAG5>d_4J_7V_c()5J>O2\Q[.AdW<EF@+)=g
M@D]@ZE078-&X+?<c?S(&fB:4V+ITS0D\<#V6./7M7R\Mg^cEHZa3J8ZFXN/UL_F
:81M0?=P=g_0-U@R^<T<ES((1JDGVN1ffc#+FdcET0[IN<N_gDJ>NLJCd+e>Z3M/
/_TgP.M,O[2Z)TbJ037=0/IQ10JHVbW#S<[BQeL5XR#7D=92QT;G@Lc,5SM&GYZ.
E@A^aDX9d=SfD@H3Uf=U4@O&_J26B/@KB\-fJ.;b(9eNbFJQ.Ic17R[#RE55S@&(
G?6:g;5c@J:]>KfK?PGMcL[f4gQ_@+e3>.;b;LGgGg[-F2<Q3@R65GCdECd[QfY(
Y_LVWR-//#6T.W6BaM/&@Z?a-[NM8B_&R_@[;U=J?94WAC=g]9(Xe0S7C;#Q3Y8;
f]DK1d/W6:g_>X06/3(UE4MKVBC15bO=W/L6J0ST&EU&P3??1KJ]8AcA(?0.X;O5
bA352/>S_BF;KVT&;^-8>,PEJGePOB<0,73_FT>70J/+>.gf6ILSE4-I,4+WZL+1
2^/I,gO+>48]@8EH/401<R_T=3BM&aRNPXL8;4.NC(M3^DFOZ^0W3bJ+;f(@9/ba
5O?YeJDAVbeP<>7(NdTLbR(=QC5D_[&L2BP;WDLL;Jd#a#;PIeKNdJWbSX8e)7G=
<4FA#HS..53cMf0@3ONU8=<V:N_ZKR_6)IS.IH8GU;Z-JTOFcKVT(6Fdf1-NfG-W
:6>I/YTaW3A94HN92<58S5ZBea2#7>JYe5:V)2<_c@f2HB^4A>E_?Y??IgG5QOC,
#C.MF_T:[Ja\B0(;C=V3eX#TRWf],J3Q&>4=4MPf\(&R3&c(e<0:\31WdAU<<fSF
,/Y@e@3ED4++9B/W;7SP=24N(5LM+.g=):B@=V<+,OI]N4[b^6;1aIcAL5I1<2QZ
K[\YdB[JS.Ab/@MJKE^<U+3\=aK14[0BH8H&GWSE:1H-KaX/4fRQJDfLQabGJC;I
<9Y@1]X<G/KL\Fd2GWBC(R](B1)a]HO.VK0f<.<&KZd?eX11@6<T0#U?<-8RbN8Y
;VV&Hd,_d1JP;ELQ0(69?21S#O_0cB<+SZ1bgTV_A1,+[Z:-H9J);+A6>6#]3eB1
f=AaeEH_TKSS6cVA>VF5)-I/cXQ(DVMO>A9LT(M7KDDPO0Z,0</,/<Z=BSc\5PFY
b(f.K>H6WZ6H-#?.DNS/ad2[?3CcFV_P)Z2S#66?Xd:,;fCaTg>&debAQ9gZ)P8#
J@Q_eV;I3bf/g^^d36/f;9FB@<@LVOaSE(]D>97L6a8a;c^<5C>CI14b#>^=,LQ7
0cF#VE2FTU.^>]_.(Z_]3S\1eQ97beY,UEWXB_daVCWH7V^J-eO=fH>22ad[dX4=
QD2_]82-9K1945e0&XdO@c)I[]]H\OE5/_\;S[Q]N(3eJ9M0XW2beQIC(Wa0(I1>
37@:B(P&LT.#YRZ&[Eb=S&;0-b-bF[4fHY]YeC4X0K[a92BEH95g/(+272T.=>Ve
@A(&#[8+XK34a81VB5V/e)F;g][TB//<c>Pbd0N9T5C7>7.G(fVYP@#:20[e1S(H
2^:(bQQSERDF&AQf#IY&R6&.,FU67YL\gO&e:U2VaX#+6L^dT.K58Tb?A=\#O(<1
SG;UfZSe?5E4-@D\fD]fJgZeK[e+0g\?;Z9>^2Ob@I<]P6GUBCZd1E10+\A[cOS7
#?7&dW/>J,P9W>?QHLKLLZf0(AQ(e6Sbb7Z=6\5-dY\E8U.JNVa/22gVEIcP>F\d
:dW.HOJ;RW+)gP>-JKbPcZX?&RI5DP=RP<da8HX.-.K7Q?M0QRFg+>U5J]ASKG@L
WSL\TXa[.=0L<\@),c^(^3RfQKQ&Y&>.G^QE\gCF47e1X3bF#bgXa5-_aK=20DF9
.\/&O?UTW7d_U2Fe+ZOE+JgVI4ZC??)bWU8EgGKf_bT;McL99U)/LKHLYC;/TU_g
G2G+,KBE2>6?JbCYYQeC74M=B0EBX725+2HE#&(d@T>V.[O3bd+,9,;X:9=?6E;&
8=H-O#Q\@]U^LMW&T@V<Qg.>1f7D:7cb_WXD/_caKSQ;N#c#U1#O+OfaT=M4_c6:
\-:J)E<C12U\YWSWUPCYCZCJ/Kg48YQ43O1f3.NSDK&TbT,c/7Jg_UWHSa5\KcDa
#cIHfJefN1Wf@E&d(06J;0/MQR#>g)ZaW>Z:W^\+5<bE.SW2Z/8d06U-JEEAYHf^
N790_9UE7#0EE5@BZ9E&/P=:#d[=F)JPP/EXa#aP[#CCC9PR1&+C5C767P5\?<\,
JKDT[>;\[)\XEUB0\V<PY\X/)&YOFQ)_^+,8/e&O557V-I6FQg2=A,cB6/Mcg\Z2
^[f,@?9NC&RQH>aIW^;44EKHUA8H6?eO:+S>UQSI-)R\4M#09OP_P4F]8Ob(d_/L
\YAXa/2RJ?XY:J2D)gDW7JG31&.9JaE^#,\2[AXG3->R;cAAC)/c_T,CfH(-3gY,
CX//]?\fKX<SVfPCgLERaQ,(P]DXQ89M)A[A:1/a\3Z:b-@Vda,.RA.EC[[7/\Xe
&V96B<a;4,F+]-CM7>/-WE#Qb50A+(fR=W1.QT8S\NBMS?N/HFEb.@cUF,&TS]8T
0P?a73:EG^H\@USTb\4&A[X\9eG/MD8)(BWQcET--&XU9^4KZf]Fd_dZ#B314d_I
47WV?S]>fIa^ggJZVf,0Na0MCO[f\GV@6cA.(C-00@<[-59He2:M=<ecIVLOe?M2
dIfH]-9L7@M-&AZMB^BQ]N.Ma@<YeAPR&I.]a9=RL?8(Kf3LAKA1ZfJ2:2TaNHB?
OPI)0;7^gd[6U,0ZK/_f8?-4MG8:21HOJTVWS)c[=X?L?OP-3NXU,QAMT-\Fa/)I
EOP=5-f&R26D.;SVa4SEYecIKbR7OQ@#88>UJWTe2JW\88gEYA@OTfK6eS1T)CU^
S1UM2#d92\3O[@8@.HHY?LUNG=F;_F>1IE]B)U_6E-EK9dJ-@+1\UBS.=gP5bb85
@L)HdW=N#(H_FM]R?4e2(SX+fOCY;HK/\?/FHN0B0RZ6.:WTdN>Yf4>dd=5>2V>_
Kf-2_D+)@b.;4LK(F[.NLT\Q-B;d)M[\AV<1\XICTZ3[cW_KS9T:Ge@=G;OceAD-
X3@#Igd+1<YMX;8WQQ>ZBc<IY6@R7.8+XV.HB@ZT]=(O1KBB&@#GPBC3+;7;,^_,
L95VJf?&>35+E8QV>[TW?Ge4b4gC@^JfN>[ZdEeC3-0GV\fN64^5_<1+UC03(\&5
9:M)XM6M5>]fEG)@7G-?VVN]-M18>.M]6aaQf0R3FEVd[Sc8:]YV=[7KQ]H,I/W5
KX?NQAcID@BYSgL@a;\7KO18F(7S:>>OA]DGc(()7AK&W-g)6U<4U?3KPDTNJ459
F)Y_@EIVdOA2IJNAd79BLIbSMOS.PX;SAWLR_WC\AQ4A3+f(5>G+V<I9B[F\.32-
Q9..&[<0dH-B8-F]-537Kc]FDA?&Y@g>:#bN_bN+G>9+);(,:&?58>03BN\^/W6a
FeeRdN;-.B:CE3:I8RZ)d.:#[U>cc7+2/F:6J00\\X-JS1[CY65BY3CfS6XV8/BS
O(V4Qg8D+ZZ74&3E1H[IT0(bc3NeIPQe2GCY-?)QI;]a&YOZO>eU;=U&R-<Rf2EJ
I(a,Ab,-/Db3I>&8<)e99EOL50;Y2_Q,8Wc4^27G@O>XR<b1cG^^6-a9S]A>M:ef
\HePe(fd<#=dX+:PD4=S:AUg#9ZZ32f]-UQ_,DTEU]NF1=L?IN&ODWdZ.?;D50L8
1&\1O,NB8,aGCS=fC+[g<;(BU1.g2VQYRZ(+]Q]\EP7LL0aQ^abZ8+0fQ@4MbNQN
g=@75<1e=>_V20B5Y?\W)8TMJBF/;ZH:6_PCND(>>]1C4_dUN1<>3R=>>ScZCcSQ
gB@;DW(OB1@\>AHLFDU.OWAfe69+dWTKC+#(QKHQ:TFH/L^g5TZ.KKDgQ>\W;02>
[B/.\#-A1[8Y3&38LJLO(<Q?#J:8IV>(P8@SX;9Q(ABEOeP.eL,B<&[5@43Z-8F^
D)@7[6NeY=6Z0(Z;Y_bQ3IaTC)(K]A,N3:@KLZ?@T^c8EQ7L+3Z(e</>1X,IK/EI
Q)[:(W3J?E7H)_AJcC?6B8?5MMHX?b\YYOK18-:A0.4:?C_?S1/(,IL[4@V.-YTC
C[def#M(4BT#54(B6<c@&WK<7K)WdJBOTMcO(\EbGP/(Ld8.aJ48>L/_DPGGb_#F
D[;@J>-62Jg&YMYY5#]\ZP(S^2<N\MEQ?B#bS,)ETFG(BOW^^O>[W]-Jc]T=41N6
6OC1Uc0X0cGS3[7@+NN<X,#-R[_M:V2=R:9LS\3^9EFZ[D+V<@Bd@-[1_RH22F0+
B=+-K-[1W5CF0Q#d1#WE_:N2bfO9/LSP#/7U^d>125:U#V1T#<3[96H-E8OSESM>
O3c\:eZfIL=8#0_JM(9:;R:;_f@5fS8>=C09d?1_QVeZKfZ[].97@Wf<R+XY^QDb
b?R7)+EcaF5_cSO8C#6FZCg>?.^OHY]_5>P)e9^MVJX(Y[+DQ#IAJV+T7,dbHY6T
T)d?I/fD+D,S,YB&&\UM54[Y\g/=2JNO:<QS:64)g.=RF/R/+-,gO2(Y,IMYZDe.
U_=:#.5I6^a,\LE4B]MY)f8+4^#J)c?@GcF#cHPEZ+<#DXGB]5UFg6#]U+8TVTd?
85P1D?R2(XK,(BK_1^DDT]d6HH&Ce=Y&0Z??\F_&A8?dA)\=OB<=(D\4,F/7N/8O
?[?V)-URD?FeP[:TEBFbMY9<[eHIPP#8RURFOJ&L=YG>(SA;AK(1#PWP[\c9dSC4
1gB)0\GV??W>^@T&:XI@fF6D;+[HX]E\F4XR[?bE?:^\0BYI,,gNbdE0#[WP@@,G
e=E7a&BV,3#_<PcSDGQNS?T@Pa+(04]OX+\\gf3f.0\U#89H0>(NL/LJ6U/Sg(-X
Yg^bAG0&^I5Xbg;e,2G0]IA-b&G_:gNO@(b-EQ,A/gLAB.f83ddXW@+0&;Y&QNHY
fARK=;S85H<?YH^KWMYc434);SOBB:M)RT:<f#B+I)gQLBT6XT8-YePY[2+)1@<8
H2ag<>AV4[1cW1(Z:U4_-c#/_QZO:1:,;YS(AZOg(JaAGb3VB6<7ZP0-FZF0:Je/
Fg\,B]8Hd@2=K//4W=4Oa=]T+.ER6[N04D&.ZGU?W=fU.:L9B^R#T#d]Zc3,KXPK
-Z6<,=W>OWW9(g&X,be49.P2^<C2UX5)5[2cc:Ff)^;@C<RG826;[0.3HC\QWE.[
2R4:c8bM?7B^<&K.Z8M16G:Og/3BA0.gTC7fG^]#S+8^GX;]I9<L?d0=5/=LL.Vg
HWYNYCb2,M_Cc>Z2B4RX<acfce-W)Fb^e+AJU^Z9_c,4:YbZ7;0V?28+6ZFCC]#H
\E27UFC_f1/D?N.M+9_R(-L2LYYb+LT6?QQc,0\5I,2-H&]OPKZHc;=\aWSf8E+d
B,c<SRW[b0]2Bd=M)@GRLZ[VN-E26[N6@EQbCXXA1@G079O/^)1acCEGA@6>I;D>
(RR5c?e(1^DYRaI\;/G1(9da-T[;,9UJ/RUL:4La6eLI<UCJe#1SU>T3Ke=HLI.R
C]0>A+cQCJ&TN:WLNF#VKWbNA+g/RN&8R49b^CQ1Ig+#L>Ke[4]W^[]W-U#77X/-
(H4TbRGH1b+68T=;:g>e<4S>Nf?U#4DT&I#b:DJH[f]Z4B/ec\g_NK9D>T8.GXHH
X8HHd6>b(E?.>M\gF+M^\GaXHF@eF2Vf0[6^DWUGC>C(,N.QI5\D9\SfeVc[AX#;
)U[+fE\YPHbXcVDQ;H:9A8:\d<5_FIJ^P7OXOIN-cH0+97A/(CW^)+U0WQ39O1(@
A7K-SL0.07S?SPMgX#EJX,V(T/JX10#DE]QR_d]RN9M?\Qa#VWQ?2E6>93Ec+F.a
9_UKM&+aQQb5O<Q5Wc6FITCYA6L&GeJ5GMUIFe[/+2N]R66G4)QY/cgM,(-4QS^[
(fXbC[NHSBCLB)H&5C7Xb[5XYJ0P]c_SI/R4FS1gQ;Lf@=GJe[:2)&</1>:E6Z2<
((TW]BG@g.S3BW1^-Y#2eRdM<^HA:96YD.74,BA-=ZEDH>.+CVO3L91b\F<Ba:[.
B320K5>/SfDSAXaCM[K96&fRFcI^=d#8.TBbg^#>;GJXE2)PIaLW@eDKEf<FC,;A
+MSU:Q)M/g5JC=L:YK/IT2@c=W5-_1?TDT<.g:Z.Y(\__bB10X/+H8T:/5K(PR]W
FaDe1=#0O7;Cc:g;(J_J=FIY?X?.]W:V?SDIEY1)PM8N.Pd6/<0Q]b_B15ScLg&8
8cZ_UDM8e?e^8YQ..=Uc19:^XYPN7)-QdF=D)@+[F,eO-UM&VEA;8aG4G]1Hg@KR
U(@+SUEea7:WXVCYFAG<07>d90WWSWJY0eD#8cKXV^[#fNe,P#b,Z_P(QfVa=-)M
([54H&E&dC]@aT4\7(R^g=GN>I5eWAI-QW@+>^E7dT)FUH,9&Y6W/O0@L;&5I2<\
J&9CYa;F6M2NP6R>&5OM7@UM=#=>;R:-a)B]QZ-2X<dY6&IOHaF4AX]Y,]Bg&K/4
>?TYDe/X5_)bF@dL=6DAOU,RP\bJ.P9.L0(.<9G1/PW^CK0X_.42B=Y<XY.>6Q0R
c?H^[:aA60fdJZXOa1Z@+\8#B;L>ZcNXQ=;^f@0MbP#SVMI0U;)<9LZ1H@Z[4c-9
YTEX&LFKN65;M.WS?Bd&XENV59.G^f\5VC>[9)e-+(MQ6:TI-S)c;V[K;#A;I^.W
W(4->Y_\aT1#D1P>QXCJ.b^-Z3e07S3IO(PPPGaJONA(CNg.<^_)d<5bBQPeL1b+
--#39(V(OS_Y8LZ#(c01cXW]]AEd<N(:PQYU@7/XV)&O=><;]<G)JTDU.Q2cg1FF
O/dL6?J]8[0)b87+RCbD3@DY+_#W_#VK+D(a/Pa3[cM/<BQ#F0?XfH\.>F?CS5@9
2\GLNL,O:Pd[RZ=19_b\IWA&aX7N@QG:;C^/c0H=O[a5g78M^RJ&6.2)Pd[1OMUP
GBfC6X5\^3LbO+3Vd&,fV5[]+;2;,O\@T+JV=K](e+T@7S2.X?gQ>8[S<bQ<7?@F
G7D=?IHPH<cDGPbRUTd4WO<@H&W810U+S^e[,PH+=g-e2bcK)2C(GgaMCb6-^ea/
[N)X:IT.1SL(NU=ESMU7P^XDINadaNaY/+RUU8::Q(DJ\1\>7e33HQ;34b);<7JY
ERB?7\?TVeEY??5GcGV;:6JOaaM2f_;A77&NZ#<^\S]EAZ/#d7Y8a#\BM_f</.Jb
g/OS?MU=;J04&G3:#bQCf[;Sc;@[cfF+>0/JN#]A1(+^WXH6BT2cR2HaUEfHG7CY
/)e>Q4[A2OE#H(ff6G&4N)MPHg#,AY;eE8UM:=@W168BRA0X.-+7XWaEQ:c&SLSG
6;1+S@WccPg</;S^+^:40,U=\+2a\O?<H[,.]PB7c<G8I\&8J0&M#D\)/)#T+S:d
Y9g6\)a+@J&0YK/-_:]H:<=>N8?(&a8B])Q)J;ZX#JcBK)H[]@+3/gQ,R)5Q2<,S
RKFbSWW_:EDY&?,)(12^U16I[Hb1?,BHR+ZU=\^ce1b,(BJW?XP,eG5F_SEcV+.8
0X#0VDI5-4B58=>&]DZH2Y[A=Qgc#T0HB-FZ\5WA?8.NY;0),BM=dW5]WSL5Y)\L
ec9<ge>P@9e263XP:dc<MIYL2ZF#OV_F+Q@<NWRX/6O,g[M@JAPfV02N/@_e^O^,
c?3DBOV#>G-LY1_T8^5]fO&39;U\58UW/EEH4@aA[J@\2NAgA\;?K0Tg4-fVV\RO
15()GETOV_?dQ72:Q<9ZXbdLgagZK:&QD;H=:O&^C.d7/0TTf^QYESP.PK=SfF^Q
:LGc&3SGB^(E+IY@egXZA)e(^P[HGDQZ?^8K66UK(#)BKW#5b;MEPEfHXd]d5-Zf
.K9_/eEFL@OVFWD1VZ[<M9[VY>PY]A7B\_PQ68NX]gB,3\\F\Tgd\L5Z&JF_N&\T
+,L@<2Td4e+VZ.08&\<.cOMUO1R/^;)@@3MWS?3=[:gT_PE7)T:)1IN6d8KdR4af
,]6:)C/X6]f/I-DUgXMPT7;==eUE^bDe]F3-/f_dR>#9g3GY85<[VA0L2<^,^QUA
Y_O73O;6ULfe(,V^&##CW.UM=8D]#)#Z?2VHZQ76MMB/Lb)AS,^)0gg,Ab-BZLUB
Ea:>g?3XT.ZNZ;BX\5<5/(+Hc1LTT7UPF2e-KbJWd<3BMUIa)K2+e7/Bg@=gF);G
]KURg#Yg-9^gF_#VBRXT3Bfc:X:,YOa4:(HE3c,[=MQ[>@=b-7^;,g4K@,ETJY1D
UH9N;eW1SF.UT-DXHK/Q.@?gf37J6:-Q@HL-YHW4:PMb&,6N-Q=M()c(X@gD.4a2
Vf@/1/4(7^V\P5J8>-30R#FP<4Y.9+6;TTT.BJHGJD5O=eAZYYb@XJAG^,[/NBO6
8B?/3Hd]LV^aQBGce9CKA?<0FS>34V:E?:-/P^=33H?C[>Z;J0SUf\U\KO4+3H<C
J,\CcHM=>3gA6UOPA(AXP:;.d^aXQKS,6S<XR:).WX(eHX=K,63bMaWZQa&Kg/#I
(EDAVM0ZeHLcUPRMc&N#48L7IdBP([;:gXF-URY\/&[R=Ae_O2:O8CNZ=FEPXQ(c
I,@,fAOP7QF6,Ib]f3AG^M:0?1c/,-e_9c^6OV?@a]^N,4Tc\#L;JC07C,GU(EEd
VD:KTDDbCc9?\@&IaZIE>Xc7CaQCMH>ZBR8DIC&1NSPO7;-VP:Gd?9Z0>:UFNK@1
]eYFJ:V[B1GERZ<e@3ag>fO+PVBW70JOENE>JXba4RW/^T[>#7O[#RgM\QP@;?Z]
R[L]^/IMR1f1@cb?c6><@[;6)<cZANW#fB(b=Z7^^G1J#2.OGF;YLd8.6PPO:<7U
\IAWcdHPeY(a_+b@J\O_TbJY9;BgG9DS@_-JGOeX.Y?Ob@(<SC.TTNCTOfB0#PBN
/D1ZE4LKg5eD0d6-UWFV]L^E+cdF@MQ#FXIg>6?.GDZgNKU_;VGM#SfJ+<)2<NN/
X1\<:5[.MGJ)Y9LQ-KA?>??:KL/=Q:GN,=>APWN<2PDP7_MCWGGIc&NFD1g-SZ74
eA\e:cL@EVWYbIa:OQ+[gS_9#\.DD;EWXZUVV?2&EX9E1H-^AB[Re=A)XP1UaP9&
3ZA#KU2HZ\UUPI=6#IgAO/bCaS=0+B[,L;/fMLU&(7df4<HCOJ#TR(Q[=OS;LObE
RTKHAD3K2?a)PX1/2baD\;G>@e[GZ&SG5:9g[A&f8<b7RDKL37(K^=;X>A6W7f/C
3f[-a1ST7S)=f.R=83BC((&Sd502#L/EJ_ZY?a#)Q_a2<3>)V1#d<d@9ZN:VK0R<
YMD9@c],bWU>\CY[Qb=@UE@#fHTIcY^_F)ebbFdO6JCX,WNd+2[_>S]fTDNR==dd
?558@&/+N?+a;:SU9U>BJI1dNfe8eG4/97HJB5Z6K7UT8#L.T#__X?^/QF4cE#&1
5=_EYfY.F?gPYBdd_TPA5HfSP-1T/adOf.6#F0.ST0?[4EK)76;64KB>UGXO0g[d
&S7RP_?7[3T=#1bf]LY0DL60VZ=0O\ZaQ70FDE++F^)DcR3:fGP09ce\1HA=VVED
3dUYGVGYad,E@b5c)a_TNCfK0F--^2IU:L>;>U/-CZ)0Z5R\J/CQ#YZb]0VWP:]D
0WR)LbUJ7UW-ZF#>1__6Y_\0/,L[]#_E6e6Tg:NAW)3(W[FC29aHcV9W=MCgLSdA
ZXXb0>#=-/[3e=6[Sf>PG7gNY[^)4L&>[[B2VL[g4,U:#VFGNdbI_BZbAUX^(OI]
+cga01e?]cH9T_<g:1;4EWIR<5>(@ER[Tb_@YeDT9K5[H>XQK^+\XW<J<(FOC3GQ
f[7)A-bW:_3L0Y53F^0^2>&L:62?&>XO[He;B[LW^81]>cb57.1e5/\F0c(0ZeU@
f]KNbY::Z4+,ZJ)JE]-\O1[MF.Zfg)5E7gHc[Z:[;21+2T4bNK[VP1/^0LURd,.#
4M&@/d_C03)8eMAKfP7aP=I5#..]H>0P&f@?fV2^[HeELc]7ad74_7PR>00V-8MZ
MM1(C+<.#c]3RMH6KJ?^P;&7..IN74?g=L26e6J0<YWO5#(FSKMT-CRcSWG6a.UH
f:H)UCI22#ESA.=GdCb#eR:gL^c\2.)EQF,[B#[eU,8<S<0,<+YFfDU>;72,7\+8
\6aKNZC8X3E(/BT9[#II1])AG?TMJ6C42;g^8d+\dC6_0\Q>Y=;+:T3cS1<Q5YPO
R?\fL7,Af6dU>DM#E[#dCS-4AMRgaBd5G;RDZUYJ<NGgXIK8T0a[S&M/9H/GHga/
)[:IY+NNPfT2<I60HO-defBWbO(N7//X\c,2<1[ND3TUcX+T>>e86EV1ab&V/-E5
DZJ]FffWFN6Ld#^)^,#I2c.<1<TGYYUB-I4-Ned6I8X&Rfg\\&,O-><I?W:+;V;/
;Y(.8b0Z#,AH_@^O&V.A.cK3;^+4/.dG&g_2WTeagV=/D1e]ABY<T&N5J,fL//Ld
]3J/P24&g>c2OU2bX6W8C0KH;10GGSB08]/L2)1E)G#-(KRFD2>=6.[<C))<H?[M
2ELR/7ZXGR+g6RQO8KAE^P6XLC+:Ud,dI9=9YgXd1Qe;4).\A.O-a3#cCA,f8W^&
KE.II.@/,c2cN=DHP\>9.M#YJ>).aX99,]cGT/?N?U7\cL&X;MC9WN5[F.RTBI2A
EcGSX2;CK6IYEMb;59:=87W=HR&F.M@6-KKg:?6B1H)eZ\&2IJ3OO+].V-+O,=<_
cBDEFBR+PQbAfZ)^^>@(e9-?,CVJFSR8b7E;6/a?:O3gSCUeJ^MgL2;V;0<M&S_=
O8(_BF.eB)Wf3A?ag>eQJ]S4UP.;b&N)CWRYCEPJgFBc@+3=2Pb:)K<I;.DZ<A8,
bO4WIKU<X&H-<UOC2F6,4#D0e#GOO1eU5R8QC5SMNbC8LVbBE_6d>\@,RG]_#9/=
<O>;dYXS[76bN&bEcK^c;c5L^?9&fRTF+ELKYARQRR@@\:>YC^<C5/5S=>+ZHgUF
2bLGb)_^+2+7WX0<Vc.5S?XA88^NA>XFf<3#?J\&Z#Od22>_3JIV1SUI1T9gURG&
LGaL<&A0);e9,Tbf+M5B@B=(CIEeGb7gcbFcV#=Wac,60H<2P4+Y3<;,Vfb)9g8)
e>EZ>3YM&fVV3_>Q:^B0B5SKHLUZU15VeSL4#Y)N1GCQ^DMO3PZSGUEe5N<eeX:e
<[_X_XT(I@SI7MbXV[aGC+OVAR0FV5A^K61-Af;\;f=LJg83H@JQ0J32U/I#E]\c
e8:PSc;MX&^76)VUaHLK5(>BUH9b[S(&gJKe1M<IZDc(SgMT0fcbdP4/J3?Ef/J5
Q<M334/]T(_I&7K^2HE&^/.:VJ0UCJd,U/6JSd4WV&/UbI<dCC?cbb_X]K[6JYc+
PSf,ab+WdYE#L_6OE68=A@B4<,NK3fa95^R?;@fU]AV+Ze=X,,^f88W7Zf=:^9J4
2P^9aG>.FLT;:dSd](Ve)F]-XBZ/JcdN2MSCaQ3@T\^70IbFWF63;cN1@EM/6X]E
=GIgd[Bf&SSF(af1_d?:4c(Fd82WV8U8b;OY0&0d;/a.Hd39?#NP\cR4:CGb(efR
NFQBEJ=]>79:e,8Z913LfN.\b=d/(R;d_JF26Y8=WZ(CFOQFcR2[3d6D(BNIL[PA
U&TZ=?Fg_+J?O_^UQTWPP#J(O=H3KX6eaV560QC9#+U^)\IJR]ZC=UaE8RbM(@VZ
5/_-8R?E?8&WVfR#+=AN_S/:?e2gd;0d3RObU.a[5Gc>,;W?-E=_I?cJ(V8fUfY\
U6DHIQK1;H,/3A=D.2:fKEJY;/eQ,BQJ4E33cYI>G5OS9)ca+YEg[],3@6,M6#X4
1e3Oc,@Q4R1[RcVG;W^M>5)]JDY;7f6535Y<6HV:?X8IC/cO&JJKdPRFYMPf3W<(
TI7THdNJ_)XU7RNWY-_>73YdT])^1-MKVgKb9?4W_^+#/PHG5OQINfN_.PDR+4/E
_GG\\TOdd8Xc>5gH=@(2g/MJS5C/;SG;5YIQJV/?;#A83K_>_WE\R[_cH2S@2LY\
EA^L\afXgX,#ZHYO5>&dS&Bff&/TX9&f)P-QW4+OLU4gB;6\&2;Z0P>6:=3Z9<(@
;7,e\-L1<MZG6X./X1Q@MSO[g2QT&LFDBed@C5CQegMWC\0f2(&LR8\DZF:=+7W)
/MUSgK<N]cG[OLDH1ad80_0Da6Q;))cU\cTg1M-E)=,0b6;eJgZV6I,^YT8c<TAQ
(OKYD>ROEaLO0F<UM,A5V.>)WMY0/]+1MCRF<R5X1+bKZV4:^-:9fFC8KI3ECT>U
<]MJgPD&M93.VS1K_d3)6+@=R;PfUTR)E^)YYD^-AefBJSJ7g@f&7EW?e^G33W8[
)]7SHA[I1fKY:3L]E:.9_(][QY:UVRQ+#,/a__L>WB]eN;^RZe.MUaeYFP#F.^JC
F)RW7ZZ6BY<WeVf3VON37FS</N=)<f<QTI,OWZe_bI36bK0cf<6OR@I1(,e(dLS?
_YfFE66YBP(HgKG>:dMB<G_<SYbV6]&0IJ61^d??g?L]B\V)+U)9J?NRbM,^PPEN
N[f=7@H/gFLB.+=QO[74QB1[_0:F2T-B2X\L2T6agV/ZCWMT2LTYD:S)Mf^[7&dC
-:+E9,U)LYeGGE7#GD7PA5(g,_4M=C>4_<fa,8@6UT#BP:d\1gZgXUd,;NSEO=L)
JfdP+)0+QN7ME&I9MB@A23IW^S78.U.]OP@VA_PUJAA;TLg#U)L22<4TCUIPX?#d
8>B4GU34J6CIIDZb<P[_H0C\PV9-_==GA^0B.2BePTLD21Xe((cF:XJ)_HbVB]_d
^LL1:Y^7B,cEQU_6QPRBWV51<OC64AN_?MO#V<,gH>fOX4LFLO,O;SN]..2db0+I
bN4JIFAI^4P])_,U5_W\2#X/dFX9>DL8^Q\Rg0QP;ZVV@UK.0@Z2D6XfePe5O:)8
;VM700fb(Od=@-^QLYM_>D2^\3AI-7+;H-99YNeTVO+-7:;(55bS>[QJ;ed72B08
cL=#:D#^G)JISRg&95Pd#,0SUH4d8PV347;a-6OF@G54LJ#dAL:[4\R[f63g#Mb]
9dN<Q3Fc5D#[^51L6eM.I-M/\6,M+_[/Z#-ITfHCaf<Y.AWg7>egN5a-&W_/B_c\
g?K:UA0J:U:fO)Q>JL-GRV\PeTI04X]PcdG_ZH]e?G;+=5#aEVcXQE3\R)_+8)-,
.,Q2N^9+4;PD/R\g@OZ.:IOBGJ.MAcL1=4PF&US36,WG2gMO27D4;>+?A[=e-./;
(5=F+2Pa.CJKZW]0JPVXGC#N&@5b9KNE&f;fBGB8bNb2VP-g@Y??aRXaRZQEIY9g
g^&9=WSJfdGgLHP.OF<JcJDO\R_LU<?=V5_P=eX>.QOL1ZB[IP^:MW.VP)]YcP.4
=1<[N>@F\adH1G(2PBBQ?>TPeeH<4cF3VB2HH3Q8Z4<W1#AFH:L5[N-;#AZ49(68
::W)5fbJFeaMFW5=O[P0CfYG^(R@341DI?X^EDHZRRBdEX-A\a86@,CO\?,Xe]b5
L3(WLRPV#YC16f#S^gC,gT?G&UM+b^Z/-?bVXV_d+]BSV\#OVfB)BF):U;\R_Q-C
185OXW-(>Z0\XcC;21<KT27_T6:8.W:F:cSNC;^#XRYLTc)0DCQB<eI1aSV8KAa2
M<E8?VPLMR?CV32_<EG8UeJ(NVOR^N<HfWU)SV:20fDMZU@8d^\W^g+O?a-4H4J<
Yc8G(=PL0eNSK5Y4g60-=3A1;<>ZRV61KU2)N@W/143(GFLdC4QB^L@a=-(:AQV>
CIU1Xb-AZ2M18H5.(RFYW,]#@d?]P1UM7Od2,@e(&H_JZ?9W;7a9GIga,DP4,1^,
](Q]gH(W9XH>RO+S6PPY-0PdS-B8c81d+BTH_,9OX2dG;G9B]6U:RQ,F3e:&&WX8
0b?Qf5VT3-VV=d1b#>[KJA+)1LDJRM5A2[T6@e7NB:^<YBLGIM1K_F,R2a/5.=+b
-f?J=)[;0#N)WOf@7C.KKG-e^IPA1BYNb>,@7:)W6B^B+OeeQXG@d,JWYPBVE5BH
2?XabG9#4gLE=C398#e[98Y:M9CQ2X[Kg<H-U7VGDC=#JFL6SPDGH5L)U?TZEgDI
E7G&Sa],JEUR.,aW4]BCM]UcDe=W3YK:R2K4N^b1+b7;F+F>/V?9)O#QTP9=?dcV
aA\\d1G<^_KHV]e^B,^fbAXKW\>A17J9Y03-]FH+U^dPcET&RO,f.d(F^+G0=^::
[3AU9SW9f.Y8f9fVY4Y-0/39V4gc657G?F2+A=82[#33g9(g>?eBGbWcZXaYWP9a
[/&OfAaGVdFgULG.a(^1>\RWX;SG_+1VBg?[b/S9d@?RH(eT^OLNE&SeOS1,=0V7
G5WL1/W3E4FD8/4B=MC5_):JK01@,[)2X)g5.bHFD^a;./QW=f[SD<^LI0B6Y_5W
UF1TONV_]?O.W&,&=f/?J.P8f9D(#b[I9dKCHYfT;L^.c+_[KXQ.[>U[=].X@TFM
aDN<M-D/CD>E<cJ-FU9@75R-<1_J9(W?DPdSg\bb^Ob=Fg[7/;TDA>d<_a3Fa:]D
VK@8MPbB]&/BJ3]LDeJV3(aD,2^\Dg6L)TXT3OYO0/A7IB,EVEE0bM3OEP[3:Q[@
Y<:cUG26DF=T,#Q#5BD9=ED,&YU9a+g7WUR:01FDb;ULV?=TV[^/cO,0\?/E^-a5
Wd6&=]2O9Y[;J2&F&K,QC1.8Re&.[_/LQRERJgFV]MAI\O4IcVg<4f3Q,=S[aR[B
2V6AS\5=SLfZ4J2,3&I\N@g^^STQ_C1LG]4fBV]>Ec@Df<B_L7R#=_N?IY;F/I6P
Da]E/DNRcFe9QB3YRZY+f,YSTdFQO>d;OR8EJH#7Lg:CP@:g]:EOPW6\AXVVf/Ma
QfDa8UE5DdBM_dZ]L@+fg\GAT10AX50F:J43=99.d:5[_6YGW;/;TFAB=AIMONTX
bIV-R#:;_3_V]O6KU0_C1#VJ,F=4A)0_Q\?QdaLUPQ):QJdXP[_e0:T.\P?9G=OC
KZ]53d9IaRXIc,?1IHB1<YL]JVLJ1WWEU],YW+^OO>_.4[9I2?3>)B1YB<S[#,YA
>VZ(4-/cNJ,2ebK3/])LC;I_6QUF8gCS<#-Z2g=1\#I<:QZOFI2YV>&63[8_(IS;
E^BFg#ef<B?=3Y9c2B_#5/TeM]/1C0gRN55gWIbIR\O;]F0R^<AXMS<+IOPY6,Nc
&Y6QUf-6@1PN=1/7)R;7:\NFAe,#P[W\_5CDHD]&e+;Q9L4XSUWOP3a1P3L#X)JO
VW[B\TSG=<ZKcTEL+,Rd\FbKZL:cZ4@]cHa22_9PPR\^SP1g7Pd(J&PYg=bE&6F^
Z5HaVAK8F3Tf^B(O-S0+P75.W(U.CC[0(KaDD;1BCC/?=BbE[/\bRA.@1F+/F.M^
V3L/8;2C2IdHD4Pe9>;#bI88WQf/0L16DGLJd(+(AHPR-IcC+)GfW92^WHHf&1&c
TQ+^3W4AJFQVeb+bGCX@R?,?WH(ef;>V9D[a7O:L9LPB5cOfU_Z4DKKe9>4=a4MS
G,Y]@eS&BJS]-T@IKRU8S#=>C=\/b[(M4b_WHI1:=D7b9AbVC,D1RgI5aC1b2(;c
D#:G6SJ,_WB=XXUKM)Lcc8eJW9aFQRG?V/,QaO5QS++1X>+:Gf8_fCeG]323OZ@6
,=9SAac<W5BQ3V>BfTKeTbcXGaAWG1&T(LC^WV.gLZ3_&#=(68L13W:VI_7>ZZ;_
N9V35fe5-1VEPF(A7<2J?bIY]ILAUAYHX-SJ1daJ=<U62eIDF#?NUL?@3?]X_F4M
EAE.J/29d?cY4=cRbA4D<N&EPQOe95LA\:HKd=Z6e?:C=OQMMI&SS1UMA_HYR]J-
D(9cV;(N&eYd:N/TWYV-<]a>.?&RRZ]B2bbgS\cS?1ag^94_:R#f4c/).P0[;WW-
-3M[PFBT9/]]2BT#;:259INV2KR49:)4PINCICR.?5PP@6Vgf4/LSXgD\cT#<cHe
NU?b4XQ<KA?aXO.7cO57bBgO+g.e9;Vg[fH?E]M7?,U3.]RG>g-+/[H)Y[5_(\d3
-:K0eAUW-)#&E-_&Re2B.HSBBP?(Z^#bX6Hf9J3X,eZX1K>.+MR1Ib-cW7bEH2b7
QG@.O3Q8[(K\9Z02NV100;K19HB(G8=EfN76a)APZR&aZBG@9=6S=TIOOX;,698J
27Z=1=Y;[dG3>#>5gJDI\<)13)9S1H\(_d.GK;XD(B^3.15MD1F)A0L?A3I)NA6T
):3,1]&-17_6DJ@[\QV[)2^A;H^U___K1G.1D7L\a<(G->\C]U;N4-/\b.db0V7M
QM/,S7egS7dW&]b<F.J@(DNGM>[/+.SA6/<L9Q<;9U/g82f;>0JWUC)_VG)^NF#U
)c-D,UNY@RL0Yc@?VC\N;-7?eSK?(J?4[8Pf+WT]Z-J@RYXIZED+2H@eNRCS8gI8
0CMI?@+/OX<R<Je/F0<ELVE0?c#SZYAN?9JQ/C4J)2>D:A3TWKPW9)UAMgXc3gC5
AO?&+CNeYc3K)N7QYQ]JaMC&DbN5M/5b\Ic^BM1Tc093)N9WbAS[1CCXXT(^,QbK
KCWMP2dYG,BYL>aUQe5(HY_YO0@_(a>[.7TK7VC>9WPG@QT90g2+6D2&\dX3C/DX
?P5Ef)c2dAZ)Q7KHX=FTY=_:W5D8dT-&b+ff@AZ3^.D&V_>0,Q@]\EN@_;f07JA/
7UB2G=&C\c3;bEd/WS-197:.(&#H4@E8Yc_+-ZXL#19<T.ESMc\&Yf;&c;BU15bA
:2J#.,VDO8/4[Ld)]6c=D/=N)RS_9ZEMe54BAAPTeFGL\7DUYS#]9W[H_-[T7QYZ
V\aPaQHSeGD60F9NG7<?]#OC^7+ZU<a_,B?N):^/+-P6#_#4c.GR&WX36)[dM@IH
#VVY>PO_7E5:@<P];ZdF<3IFLY+9K,??N\IgK#;\DU[DKEG\A9Mf4Y.9].C)-44^
C[Q9XR^I?26b/2#ERQ\#e1C8T]J?-DNc.^Ubd;35KN/g;<8SAdf^SLI]H[]Z&cc\
F+)f:;GW_CJF,c<gE4@Hc:NDgLLW^cQ(2G6O?],VGS.K7L9WJ/_K5D#eFXV/K9\b
I.9Q8)=4U_,cggH]=g7?LR,027e(PO;M@G)S@<T(ZC,1V)8KM6>_PLOH^B6f(F?e
B\R0Ac1dQ[?/[PKa>faLD1d\K8MF<KI1Q1XD83YZKcYXOQIfdMO:^bS.OZcAG+V-
B-Kf9,S:GS94/CdMRM5&[HfcY.<W</PR])@(F+OD=a7M0Ba4<C.3c7V=Pe\X+C99
_&G9=Hf?W@]G)e,])cD;c>ZHQ23OL.I2EM:8]^(CFU\(dI@\\TWgPNZL<A^Wd/G]
5XZ<M-SL3N1Z2(V])e)-IScMMZS/TT7B-IHPb(FP[)C:(<E[8)bEI_Ce.QFVN3,]
@&5J(T.S]([G+1P_BN9eW)g@eDHf()(eHST7VB8I:fGg0)B<M(cLMRX9W6_A9VdW
)FD?:ab31&H(]F#6@12a9eM;\FF63J#\W+[B>f\QCT[M<Y_?aEFAYRB/Q[Gf4O,Z
WD_2^1b4YHO&BD-aW-\ZL]>1@PSJ4ORZaG5GQ5<BSXNVYSb>bD=<.Q_2<]SDPN7C
dHVe;(BYOSL8@J=cGG&BgZ-cL4/8D#H;6;-cdN^,3R2Q<b4>.40CT2-1^?dW@C/f
/7NWc7I7T@NB;=?,--McQW<Pa0>.ZW.X?\^:L_/IL,<B>&,89+_Lg2cV4Q(W0;9H
BM_Wgd.OI+<8LgZNV3Xe@V^-FIgM7G&BPLWee^JBT\Z_#F5Ae_3=^fe&>P^J9Q9,
\:.\PORXL56)?7g>M96OEMA+14F#.W=<N@,X+V&T2]c-T1cJ=K4Q/_KR3MT9=)F2
@-3^&1,8QR;@@g&9Q7+Nc27194(OVdg>(cB[KV:@]0BS.X2#H#LK)&PO^f@;^0KH
6UQ):>:^bKbP)_Fd49F/#C^7;J@=UDTeT\TfTHW0aL0ER#4Wa6.(AVM)VL40+^:A
\?8I^E=D[g7Y8;KU]Y&64Re&]5WW+S5S3+@9>N:/,33Y=?>8C)eGYCN/=8S-1(0@
M.0?<&U._Ab)R7ITe7(@f(14IdR,O#Pg_\ZOR0(>UY[X4@O3V]L08W\/AJP/U)T?
Z_cNdd4VBTG,T,e&[B<S^+<EQRMLb2AJH<NGdV(PBP80b0(M(:@@J_.:S[WKT<;=
COdb>[)/K)^TZK\Ra&d0DW.9e?g3A1&]ObMfMU@F2.1Q2RG9X)#KdMC&CZW3)M[^
H2^Wb[:7\M_FR+)GEG@0ZLFT;&2>M)@W+NN-7N=dBRe_22XQ+f)KSVb/a=-3==)P
>PeXOg2R^#4<2<ZT.[U8_Q-ZKTfLF9#+P/Vg;87:bW<8>_(AD4;WSK@&aDOeadKH
AfAK01c=Ia31?[]N?MKc2CTcR6]3B2)(C&WWOLCO]G@KIbE_L<(9f5(3;\]63K;_
(I;M.8U5CMa2/ZfE6AY9TU04Pf)4#Aa]/U(@&6dY7\@X)5>NZE;T?R&ZSBUI3ALb
IE39VFJ/IV93:XVb9;e0DNgUg3QIcA;:&N89OSM4MUa>Z\;/<;A4N[1KCCS-943@
XY8I_d^FA32TN=S;]-L@VH/AR^?KFN&gZOOgAW=XDU0a#_:L,T,B#HM.7g3ODAG&
&])O,:E(@8-HK4EFB9)cF.@+d5[KUST7O#N?A-Ngg5<R-Y0?(?I]4cL#cB3:&<&b
?@(V&:\7dYSF/e857K/&T)H1.a<&_#_D-&fcQXC[C/A+a5a=F-/LgEOSeaeG(MaI
e#f.XZQ6I0aWK2aYLQ,Z::aAMN3#_4BI=S87I&L_VgOUMO-832=cGc^YCO?b<[aG
E@=\Ke^gEY^6@HR\\#5gTA@CLR^:Z>1A/A_;bU4]H/Q\;/@+H>6PXU9F\NVPgV.F
8&_)5\?NAR-02P4NA73HDMIGR)<R,;e78=\:4Ofe#)gTf(UF1?GL&6[aZ3I1W#JP
OPA\:C-DQ?7gcb/-FZ.@CT,?5f=;24\Y)>8G#ee:Yd^IG^ceLVSSQ\dVFE=^KgSa
[8#+Q?Vcg<)<K8JFKFIRGR[]@-ZR(S0T:X_KSgWd\.N0UK2@)gaMH&a0g[V6)Z#E
1C2OST,I:[I1V,#Y=BUH&G(]7(BbL/DPR55BJ77J;9P8#?9T^U&4f]AO:[+?e5<1
X.A,Tbg08=_<^?QUN4)CJHB>R9?>2B3\K=#UEF&^)/N=>dP3>36MN?b2,E(C75)V
7/#]3=T?RG;EV3-c3T)LTAWB79@XZBBIV;_eEA42]65C?ZXDN[<FC0OTe>+]]b3:
_9:,D4.[/Nc+5Y?a>#XOAMFd(=R0A#@^BAHOYbJ;=NSA2+O8&F5.X9f)U5D]=()_
a#J?9Wf^2<Q:EF><]HaK)@-V-KPE:aIJ15>MW;RB1>P@(Y;GY8d(_BP<bHFS;,:@
F+cY?=RY3W.a2;]9W:a1aJEE0<H7bLASPDFS-H3LBSg\YaL7\^d\,8E<+DFB7L4a
S:#(ObL-Z66c70NfRL;1Ad9ILG@[Qg-5<2bU62^:YJ_b/?^\H?&g[c?-8Q/;2VNE
gc=,OZBD#f=1Y,96XMX[-A:2Z^6^FHQELd[,/eA]NL?OA_LDZ_dOa95HTHEPcD6,
eT[7#ZI+IaZZG-a\O/LLdKc71A@6RD::>(g0MIVYV.CE\XgbDF1KB2^M8B5_8d=0
?W3dSI^T2&6cQ/>_IYPRc)&D3UB/#&ACNf[>4_\KY?/Cf,LZB/3\gU-5LQTUL&OL
C]QBLGCDT[>#8^3H&a6I-WVL[,EI8C@>DS]N&7O6d)gN&[D7HW2\<X19/d6U3QfJ
a[F,[dWf+?RDRIQY(P>/W+253PTfQ7E2FF.UX\.C=+]?@&BV?cdcO/O:3,BN_@J,
81@C688fS?e=UKA(RWMc@[RIDO)-5ACB\C8M]ZSDC@0YT08MH_0:aVVC_e:),#bV
G+^4D(>>4\+1EN?g(99IVT7A166>5VA@(Qf/bJF#JS84JF]..K0ZBScI(d[8)Qd?
f.U4O49<>V;Y_CU@.V^^+1bEX[1G_#L&c_A_\UP@IX3GSMT(TACKbR/>#]?P<N2<
HKZ-9#;#15/07Y2OF?Rg.SY=+bFI/[[_V&>H,PYC:TCc4-BgcB14F[QLC63)@P4#
J@-N6P\AeaI4<&a&)WaKcUf;fB?\DQOeg8&Ndf>gbg?0=@OD9gFV/[@/ZBa;^T(Q
?B-e^):H]Ab[VM+SJ45\N8<,@a<VT+J2:I,edf?1>+,-<b&&W+]J)EGQAC3_A5,Q
HfBdHbA+4PMXGV^/\S_^dT+5,&,CaDb>dKL4>Y;&Z+27d_1TUA#A)6#XW=4@D(S<
^^_<X<^(gLaV;]_;JFd_@?ON=#6B9#dWI/A(+Eb7?gBVXdg?_L1FH?^47JBE&)DU
bT-_S9f07MORLa/g/4]5MYcR]#Bg/c6aCBM5\S>c]@#<QN>C:HA\OQTBAM5gZb.W
1(A[#NceBZ=8LE?I^=R+f]c4<\0-bZ<30;U8.QTP)^E6(I(7/N_8_a->)972@+/#
/:c8B:A9&EE]AML1Ud2bT\bFR#NZJQJT]cGVR6:28YfaD:b[9>]\c&DTV;[a,032
)E?eU]]7RN((eDb6>e-^:GE0\c8@LXZXP4?;^e6L]6V]YFFbC575ZfL6=a0cQWTH
Z?C@)C\^I#H<4>WGX9UcW1789Q7FV4dTN<M6/ICBQRBF^^NDIY(SaDMDM<dCLTD>
a[=1XWS52NG)/F-T#M-:cVa&[&R.OR8.]gNHd53ERggT)RFT_-I9>)D0(PXg@5Q1
eTE?I_[2_ZEfJM>C<V3:F^=H1E^=C4>e0D8F7KSF7ab34#?)E7_O?H1SH);7_.E&
5Q2RdQ[g&]9a3fgCOEUg:9M2cQ&^]OPdOCaV9/QCMEgS.?^d/[OUdQb:bVUI\.Y)
1F>>LS#^/8T_AYAb4fBE(?;W3Z:3.BC->,YWOJW?M=+ISRbf1Pc)#U-L2B\K-<;X
gc_&Y/5a(?LF#YE@R(A8GKQ--_>YZH8].=)[&JD-BP)UGB-G=[f-TO5.V;1-7]/4
8^7ePZ4;:6La3PI7S(WM7UCHc/[K=Y.5H2,e=AIRDC:d).NWb,e783AKTV)-;(]M
0KK+.FX+59.JWf:aIKa=4BBV]HERRH5QDI4M<E<gca_d8KG+ZI5[9:MLag0IYU>E
]IGQP719/T#><IZ2ILV,f-G)<\I#KH:d//?ba][:caZMB)CZLcE1F&R[>B>-<9?a
<<#U3a?SS2+(XH5#LV&_RHSJB2-#\PJ)b;)4F,eHdba-a(<[U4OV#1F=.)O(^[<Y
0PYHFO5ccQdJZ:K>ILL(8OK\cCd.\C1Hed/G0=KIcT\]#D[1F^XS[CG.(SFI;4LI
4^M0GE51GO\ZPSR:B9L5JVG\L:Q1^>9QSNZC)D_:aH9>9A6d3Jgg[1I3e1ag3KA&
&9gdT+L2@;40?52gae:;.[WIM?.0UE/Sb.AF9Dg,VE[OBQ/&b@44,G.0J?1ee&L5
cKTe])YTI\59>3O8LV+_Pg.OV3VZ-9b\[aO[I[JB\>IBRL>&_0\WI>RB:E-)Y)BD
fNND>+eBN2HJ37G7]4a:e[->,=P1LS>LM&-5>N1?BG5L.QJ2dPK_MF9D@gITIP9T
RQMB0S#dFBP&d&E2dX]a]T4V)(1[@=OAeg;fX_Xbf02WX8<Rg7UA;&ebMa,&eW,?
IQJMS[IgVLEaL:,5^)^7KQQ]Q\6?4FJ_FMB0D0FU3a9_e]_/(9.0G?TAWO1HRFG^
HR<[DaRMNQ,aJgV)D246f\@UM?g-\\FXOGS^,eG=e+b,GTNa[VT7LNF@EC<<KZ87
T1f;K@8c)a>SYOObD.BM8b#:Y(DYQD\K&6191d_W@-b8C:Z>eKGM?=4X[TUJ05@/
HFg_+CE^B(T-6V3;LDN/c?aE]_,.,56dJ+.P@#Ocega^Z<+c<NY4?8,bL(BcK@JN
SV425Q3gONG5^BP-Y:6)E8Ed^,\?<H=P0Y?3-9?GYR##B8D^e+E8/;1[N3)BW#3U
b_Yg=]O37;A=KU0:1bV.0E4;&;4cec6XAA&_K<Z\FW,-0g>A^ZXc?+5XCE&WZ#ad
XXW^LeA24bYV0B&gaCc1U9KB:SWTY@0cc1Ha]HY4_?X5_PO@DVW/\cOQP(ZFNZ2W
];\8eV>dIW8T;W?Y&G)XB1PM]8=R1/#efA,Z76>:OEQ3gSK1]fS6g3BVA(H](JgV
?EfAfVgE(XB:0Y(aI)R>>#-1YI5WU=FB:0,>cH5;]<:^ZORKGUYL]YMN\VYP]Q)<
(&>bYBNH\e#b)F-fIEV.-RG@8()>)<VB0gE.\Z2-1e[7AKC8]/P2\&^0JI.+]#I1
Re&]/,Z<)57JB5R^F&67S?H=IZ1CU,=Q(FNJ_:2/7MGaMHgI.0G0G:SK^1_^5YBP
52ePd=0Q?^A^\A/d[GFMSJ3F_H3PX&5I2TYOSA+G:ANdS@HR(MBB0AYgEZJJ;U>#
FdP.UXaMDSF&P5I^^3Z(0P=P?H5Y>GM27\\Qf+D=#^\C4;KO[6Xg_U5[-N4.X>D=
5K/cdAW2WA=0Ucd>:LIBXfg\K)MB8SEg/4.33b>^cYOZ:C[M>:&>B7>A@YKOY,0b
/<OX#HAI<R;;Da3>_:G//ZcV(2B-De@-82LQTQ-#eXZ)JZP<#MA0KMGbUa2bJT+7
BY8,W>M:MfVVfRIO#C8J>/H^+SCSfeF?1T9)M,R)S7Q,&ECA2:[U]?-TaJFZ#YI9
_Jdg&X[Qg63RJ\[EecW^Y(;Nb(2EYKYS-bKf:SB.T?NJ.9<^C9?d6TLag(>IaHU9
G&D_1Ja@b\IS?[R8DBYA>g6fU7E,DN>FP-M7_DFJ)cb63?2]+#(<KIcO63+X_EU2
CNI+HM([J:0g3]0=RbGVV,fIM[[#@]5^fU(M#g72]b9=?aHeRVbH=>Q.C?FJ4SN@
^9BK5\e(g>7PEK2fG2_f<fW-G9&))e4&b(;DT40;[PI.LaI^Lg6L;9D:^36\NTZS
\E4fWY3I>X9>AL_K?d18><9CO^AO>WF=<LF1V3J[<N?72\2CD;C^9JU_)QX5S9>8
e<:803CYZbT8-FQ5aR2a4G76+aRXT;?YWW[>BL7-);WK-a9c[9>U+:J8H>+OG_MV
dQNYF&QUf[:KdJ>:4W)IT^)35.T\E(B1ZQ.U:V[NbY.<<WF2Y\Q1]?=[TW)Fa?DA
6WC]b&:<&Cf;IYa=(Y6BWT5-eHXRDd@@?Y_(.;XSOITMc_AKP3\BNMcbC;>=03AE
)fK&YTE_Y.dPXS0RL57ERC.)G>Q:TXgTXeQNM/3BbLZ6(/_[2BKge0^BH>Y=+QGY
bRK--KW5cWbWgWVN4@/-<b]X-9[F?H\UTf<dRX3eV:?\I#]bGXV(3B#?.?/Wc9,^
A9#_#Z1Bc_=#-Xb<^0]VUWd<8fOMWNaGP#,(,EH-QF9=\-[A_b,>CCYQ@G[c2FD<
+:YIO7J@,cH.JKdHY)?d=1B;)eMEHVG^R@DO[2KJ3HR@[f:WSX=@=LbB]IIc/3Vd
0QE@\gHV\1[Ra1&EcY3&L1291M/<.FH,KSN7X,Y[[I/d,RK+_O4@BVN_3__#SONS
I-R/RN:>-g8,,cR9?>TZLL\6Hb-7:TbF5gTMYWG+0G7G0[F8594WB87M_WCAaZ>>
T/31H9AWg4OBWDBS?[R^WgC7+PCbR7T_93T=AE04Y---e?&?:G]F+C/WRgLE@d&b
>UEfQN<&_F,T;NSeU&_4:NCF/+U<b8:[,QeGe?XEWI1+PM4847g-2Q7ZZL#3NN@N
>XbPgFUU\Y7W-NMge<X#TS1?G=(TOEL_W>Yd#N.1UXcIYSegd,EK5@JX.NUE,34d
0F\)BS)GGEgc@:N=KJ=D[b/6fg=FXYK>P&=>B+#;[]c]]G#YOB1ZH<EdJU6<SJ=I
dMgDZ9R[dI6=.FCeJ?6?^Z4BLT,R@:dO:fbBgK>72W7=@Z-2:MAJ]08XWFb-1gAK
)g2&1W/7R]X&;[H@^5g_84;U670bS08f,W-]GN8YbQ^U=Wgb]1g,[Ica3Z)_6f#R
-/QBV\N(6K:KHUE6KK(53VCW2.X>;^[?S?:\,P\Gg7>&+a;UB[0c+cQ]9:Y/D_cL
.4:6e(4&Ef[T14LH\2&+a+3a#OU[CW97f3GL.XeAAQg89IBg-T1?1#X_ZD+ROOQf
OTJe.a7,4^DRad7cC?#?M62G6d6WYSE1KT&E48.00V4XA+C[<1Yg4,6_F1TfOHF+
&_\+XW<SKPKY^?JYB0)T+9gd6=3,:a2VU[,bD/&X.1b+#>d&WMcXT-5NSYSTfRFA
9:](BafR:)f7N8&JFR5Sf/JY:H7U\P8@4O#(W0eNWB@NIM9a/bAfG\6R67WOPD-T
XB>/Gf9bg)TZfebN;\]])K,6Teg,7c]e\B47IHEJB<@@eaH1#>CBLLSG<GQDBWQH
e4=-8AOLP[M?eb>2.,dK5AAgG56;Ef6TbL=/gT(BME^_/+,HWQSWQ,B2BbaeYQET
R^,@TR.+eeW[cE>UY;I_-EE(L2a:./@<6NYK9PaS+;fR^Rc/()ZHR9#1CeCPdKKU
c]JN(4]fP0&X1g^(CPOE\NC0_+/=J:C(HF=X^TYRN\HF-N5/bIVXH=D8F^E@1:26
&UJS9RI.EaFgT&+[3SV&8LK_HCK&+(HE8T8JO4/B>C10E:dY(a@YP[JFLYM3KFS]
:a^gKI3?4KM1C@FeAPHB=<Gd3B+W-N^W.1<V-RE6MGY/EbFZF>b.5gKS]9f]Vf;V
<?4B/1<bXJgOQ>GFUI1(Z;\D9&=+ZFO<AG)=&(NZfUZ5VIGW&MEa?U4f5-(aG4\9
5<bOG1DbZ,Ff+)0W,+U2-eZfQG4_&7P;Nd^ECKT#;VVK9J2JB(=8>X#Z5c<F=70T
ERG.T-df80Q]CfWdeF;If/QZ=LgF1#a[aZKD7Aa3XUHa1&,Z&UNg<L,8S+27R;<X
He+<a57IA.L_OK;CLT1XH4K&#&^X+>EEQ-QYAPdMg92Z/QLT19DON1cY(5CSC:0_
.NC=LN,&F/J(Af(O?De55Z)P^3bMT4P8I\1IGIeDT&c.VIRC?aB-E(2\H/?edV/,
DX?7:_cR6ged3IdMG(]-cR+c9@&.M>?Q84RZ,\JS<M_V^@de/7ZTV>(8+F-Aa>aD
D3\K3)d5+g[K?Jb5DG@JEUPS5,V1H45-5QSd\G+D;=T(dggMMT0^E<g)V0^W1fGX
(Yd5M<-/47@Gb^)7Z#(Y676UaCHLVA]3:@6NAA;Y2RaECQ8#)ZM0YKN1PQ6.T);K
1\<b\V\gJ#R;5)^.1INX@17H#1&+E20)F<c]S(2J0?O>g.eJBG(LA+=R^5c_W(9?
0<+Z41bP,6U[J\.eQBXc<_3RQQc1JY-A+cZf>Rg;0?4deK2>:6Wc55ZPE+J+Z.Y;
U&K9LHI_PKa7b^UXCT)bOO&&NK<#B8gJ3YKHINT2?8dG3[OM[&0g->ZAUJNV]66b
HN#e189<+2+]7g&@N;Ub&X=DJ6BADKf+5D6cAW&6>0<]Va,O6@?)D@M(/H/87^R_
4cfYKb-R+=;Ec()cX#7@T1>GFe(@NIa9]-acIZ\A9+-J0eWC[_5KJ\/9c+SJJL>.
e6+GME/=D2I8#H:7ZCWM8?JFE^:fQ6B9N-?)2)W]_K\M)U?)L<Td8=(#VPaEFf@U
IH5T7,.)ReZ.:2,5YGg>GIffGdR;4J3@(\NCfJ[LZ:g#X@)5VXUP<5.;]K<8+YJ<
ZEV<^2[:K]>X)c/5<Ig^?;//.K6WF/]7e8T)B.S&a@E0+^:-S^ULZ_==eZ:.Q&1-
1MdXaL#5b1CPF8/@UX#Yca34;bVO<=95MH.^H[7^>\>Gg].D\:O8@2,06_YN)Pfe
R]PgGC>&K91TO;9O1==;e4J2IE/e=KdX@e4+2EG@<Xc3IEY_a&Ad(RV03:RbE.[4
U&W440Yc\-@].V9.[N9c=_]:EGW(?HY::GO@g)C-M&9^9P\9_E=5Y4/P_cRUgdb,
3JKFVQ.<QeAV16E<_=-1<=-ca-R6-QB\I743K-CQZB:-;__@SC#WL8=)^R0,WOJ:
ZF9\f<f:B7@E.QR>I<^XTAJ)Q?P[;E<0Zd3I7=?Y,N]?UX95c-)e@I3I8PJV-I0b
+AJDHNSY^5bM^3<\L=Q;b2e8J#JW?V[0XfCR1NAYICMNBde=FE#S>][\]^8Y7\Q8
=gSaAB:M?+TJGAEZ>O6AaATV156_^SVd(,^[a],Z)R6aFA7JM]NUc0)aZEX56bL;
1)b):5CB0/K5Wg699?d@VI<GPQc[>/)SN3:bE,KD>Tfe9d++5eSVOAdN5X6&#K)_
,BZI.fHB>2Y9T;5T[->6N@RY:58aF:->d80(N):Z(\Y6S_Ef\+UXZAg_c=XXa2fX
H:-VWA4TdP34OdD,fP+?S>UP_+J)c3YC>]3cE@I[)MbRPdXXW?F>aLFQQ(,K+b_S
]&d;=WTUY^dcI?YaYT??.Na7NeMc;g6Ka:cS+f:BX&/6\@-M-)f5#I(dL9#(R6S?
b[J=6KS0IS.N-V.5DV?^F,6F9g9g&JY=UT8,.=Td5;;a\<I0Ic.26URK5U-]b/+F
J#=>4@@6.b1(J&)8HJ+2XASWB,33NIVA;/3Ugg.EY+HU8J]&K7\cX<eg;VQ3&:M+
A+3eS?&(Q6Ef9YUDMDQBV-5bX3[6UG68WVLB&H\BVFd]@&7AZU5E?D/\)8-#TSS3
+.@Y;68a=@@T]HI1K@737G^8dMW./CM?aJfB2>g+52M:7)/[,[^ZCDMD9LXRMeEM
+2HY^>6O8ZC8?#J#PY:+@=E(_#=WD\@gHHUH,M_FQ]>@)B9g1RZAH2]7<T6,9T6C
-fU<feR7MZ=/)PR.fOYUgBcZ4&1EEO.#&,VgBPG;g#cSR7ABQ;E(7&(Zgee\A-P5
(/Q0RVSB8W-7@,Q@+dA#;,gX.>d<:eA0G9(b:A\ST[H&;dA#JQb8/,)8B+M]b6c3
U)bN-gT[fd&L-aIdKY&T-PZ-10e:C:>@.B?4568):;YWA(M8aCCSbHAY+01f7M3I
\48K4QDC>A;^#NENSN49GZN4N\RAc^@e(5Efg>\8786)D7V>-VK@858A\P?;Zf#7
\3b@#KK4LURKA+e:41=^AWB.YKK7EA8(?e&S<Y2E2]Z0MWUTPX2)4TSb5>DRX)f4
2O>_]-@CKP9K_CGcNfSQ5M[(29UAP&IHK2DMY=ZJ;&egMGRYCH++H]VBD2?OFI?\
]cB;4^00;F9SX1S0#YaEF+f^_U@\W\@4&;0I]<Y^BU]91KT1C0Q,:(I:=OJPbEYS
]AgB&?c#GQe(_F.AOa>\1I22V:H_S=\Z;_#M)WP/GQbAQQM]>S[IgY8E0B,B1L:;
A=#\]8.8AY.PP5QXWHXD(,CCL)97H,(E6RQ:\Za&&7UMa2b;ZXFF3+)#B,/DAa,T
>P[:F:</YaQGYcAc20Y?6O7:Xfe3BM9bP.Z?/4^=@R6O0TgYH8B;;D.d-]e4eYHL
A\^.;XXK-eFY249ZIR>O0H(\]fSb&e&>+L[e/=^3\a6SKVg;]AYKW=4b_g5Qc5UA
+5R)I+9]8MIW(<8CJXZb1<MU3Q3J41)He0cXUcWOI76U)QH\O=W;.,U-0BSBbEb(
8YZ)O-^_dd(Xe7Q\f7C4&HV89_<O8Tgg9MLZ_VC-\N4c?Z5/-#.BQ[XE/AQS#HI?
bV;\ff1&aA-c)QK4BKac#bH+M(7JHD/c<98gT,].Ib@=\H]:dS7>_XV8^fG[/>2,
b&TEcEKVPa&(Cd=#M3SGWU;G:(.gIc^-@H-ggOP?(4)X?g,17AcHSg_?N5N),EC#
4-;dC5^8IK3^P]/V,3@+)5PN:GHN,.RM#4\2[VU5Q)]GeJT54GWTX4[M+Z\(&b^R
^V5fcU(0VU,),89eUMQfe4VgG1/=-ONcdNIcK@[6#A:Jd5;X/P]WUPbE:UJbeIQT
f)LY)&fQUa^ODg2?OF81AET\0TcD[8:bV+38c7W6K]0JZ0L(F3d;-5N\e8g]cNXG
Q+25=.C6-TNNB_df9,TDfYYZ@31]Tg2M7@gf0?&EQ682ZV>#7NP8ALGX+:e9H11H
>RK5YVU[_K,=/V(6<=2W6bMPZMgL^WJY<gN_\<AVV]FYR7/126G2A:+>CZ@/R7Z^
<bG,L&d2R6N?U<H1P[11@\BS^b.4e^&XLZ(JfNN&/_=YaV?;552/_>Z=#dUM5IS@
P>^E08;Ad:<@.R>K9X_T8TEIFLU.LMZSLL6e8Y>Qb0aM7T=-a_\IT]6_1eNe.6VL
Ag.550fXQEH&<XLWMA2C-?cU5A:E(I[0&IKW_.S6Gee.D;GC8SCP2Ud=,KP>H)0N
=FC[^CZFcPc[CD5;EEPD=YD-<.74Pa(V2a(:Q&Y&5KbTUV@M#:::3H_Y_I3BdTT7
;@A;CYb<^O>2C&^FbfR\5f&PJ:&D\49RET]/>]AI_B.UK)g3;D3#0#;2XXXPbPN_
8Y3>K=-](X57La-J(2BJ7YG\aUW3YPW<-J@3ZRPcCPYb@faPT(c[M]]BYAcZ:AWC
E8TN]B:/b<V:)CG\&4GXAB#ERTc:F:>SS(B6c]YgP^S[/O;=H4/GWZ]S0810U?R0
#OV.@ZCc+=I:G/D]V6KFW?QBg@HO/T0ZBVPRa=L0MC5[^T/JWS4O,gW.CcZ]6OgA
Q8&6@PTMM62&6GCOa8CIX/Y[7Ub==BUNTgU]c(N<1f-2g8WT:#<BML.QD^eV79G?
DEEJ(c;KKaOE[aY;2GQ[MVI],bL/7>;Wae^92;EF(?<R<(cRaHcPf-)SQ1HgM(2Z
IZ_gG><VCLIE7T;B,/DH_^TOf=Aa,97d&G5+/Q3E4Ya3C\ZSPVLfU.QWXJ?07b.J
8(gY0FL+\D+GCJ=RYO,,22P[&5ADBRbU0U_BFbY[0\B4)a+1@:#&5cc)>/E;g(Be
WcaO-a)Q#gG+YL8_#J8.@]+bT4R.c?g4(&>d54U2PN5Pdg8G4;?Q::_4>XEM3J,f
VG)6B--FYN-G>^LaA(0C0Ba3WOY9SB,Y@Q;[;8=+d(U2-^(A/Tb5O,GI+Ac=HTgY
fA#I&\GCK8XQ:E/+>_OecL_>D3Z(bF+VTDQ#(F+M<IQG_c=9Jd4fP8b4KL.(VT0a
fK,ZAE2UY\eYQ+c;FgeE=T/NK2Kb:4,8Y;A@AK./,A=L-.TIddPPZNdf<>POeU57
SXN+Q.&&7CBNZX+9ECY2\71HYReS2^Y9DbP(HF)Y)0>;0T?=H5._0KZ:<M:XO9.9
Tc0@OWFS&4T[[ge2>b\.;Y.0]VCX^Mda8C&G7/=Z@:/9ROg<E3a1BO3X)6@^5M?V
WW#=PGZ\Q6+Q2(@F3J@4OW]Y/4LPca,@<]OcN-FY7+3S_/OK-Sg_O2:R>;E/AL11
2e)^C5c6?XGGJ?PK<,<#>DKZg0SWMG=c9MD8UbZ9aeLbPd]a]/TN44NJ+ZQZF(.[
\R^0=NFT69ABA)ZFA;Y#VSENNR>dcCV:W9.#g5:J5FJY]Z9=A^90Y]L^&0d5&W#L
D>;#dJN>41eX+If1SSKWe\L-B.@@Ug&6;#IfFGKaDcCbGA:VJ&a+>QY#LF/E6,B_
1f;LBC:4QTXcRE:V>P]74NUeO1bL+WeO<;.1d&;_-:g1D^BO#GRQBC)[<H6I+17O
\6],a=g_.#<U:5_g(ZV\HC.O4<HcfX=9#e.KMfe(I.WCL):DQc_dgO8Hb2;L@30I
J2^^I7DMGF>XA6JXZXf>f?OUNSB=4UEE>1M#6@S,=EZ)R60)-6;7eDKZ=44LXV#V
ONT]?G2G_]NH0+:Of7_?<P&0JDfFWW-fg0I6.?=5AJcMAXB^^e7;9K2))4L=/La7
FS^UAPZ59(JA(?6/28<_<FFTRM@UcXAFNN=;@gI4BLaR:PY1d[V)Q&JT#MDX70TC
D\4N^-<V\Ue+&8R?a+.bS;#.A\9=a2&\/T&b)/V\C.7CS)USM/TT0dU#)DJ]\5:(
gI3GRIL/QaZg(-bX=c3[ORRU([[U5[G];DMQcI)MLAHE#R1HIfCD^:_OIRDD7RQL
Z+)Ud>8.?BZ#8.U3a\9]R1g-.K@VIcT/C:5=(f4.b69#C&aIeT^/7P+2_OC=_Vga
g]Q5)N]4d@TdK2a=:+3)L,UUVXEO4RgYOS]T^bNLL]-X.Q4I)YON+TR8WdV.>:Q\
]GWIIcc:S#7QH]5ZWb]E8_806fJ(bZ[8L@>SbB+-g#g-2=Z,.fM@E^)^7Y/=0?D6
[aY=,f&K;3-+HO2ZA)^^2R#?1C:LfA\&fUQYI1,@1D,AQ/aEFZ,9d&.fA5=,:;.)
8UMMdCERedKS>:<2Q\1;JLV;0\+X^9UTGRGN3f.Af@;D97f6::ZF_YAB_+MH&HJ4
#Cd/:a?VPVa;<83=0U:&(HNT+H<[-U:O]QdcH/KA7#PZ2O^3gONW=.]BOR3=aDDK
9f;VUV]4?GU&F(A7/@5M@ZP/I^+;9N;\O>gA55=)[-]d]+:UT0()XJE\282IR12V
1>Yf[df#MXT^LX1dc2IY]#fR#,-)gR]OOd2J3dKIJJMH/0#Og&=AecNA1>d@AVg&
I3?X2YBgL/\&VVM(-Ne)R&?2-4?_3d7g)I7@SF[XECVL&+6[abbfK:)fRRN.A\NN
O^\,?b2]3;,I(He;ZWUKSY0H_#YKK=AGA_R]+]O&I698##&B74@A\Q@>?a]YW#):
8-=^/[YSSS#g.X5H1C?f:>dLX5d=Nd,,PE(1G2D.edCg<cGK:D2ISLUX9cADMFT0
e=a,dJOISZacUZU3eH@8A?#VEZ:6F7:-gOPc^]LJ=a:HP;@c<3D(<G/ce&Hf^:M>
&D3Ge2b(?DDLQ4agbMN6U.eaA1V;C8#F+2)ITW).ScMHSH<b=MLQGPBA>Y-d>9V?
GX9RA&>L01d#V(bPbC,<Y+Qd,(CM]613d.cUA\JDH>BB7OBe+N;d.(A?Y26;OX&X
D#FM83LO.Y1.YbF^5,(Tf/UdX>DQG]=aDY>.9:XbeTOGG7V]^;>H.0.U/#Y\,,a8
VT]/^+0\Y7UQ:J-e0..f#,O<.J^O0ME:J5L1CDGC-9&Re]>YBO,\g<&5D;V/2)b)
W2WS,B^&<UG?A<Pg-^N),ad@cc@2@L>Sf3]EI+V2?G^^V^TeA#5]H<&)U8N?7ZFZ
2^<[;eN_<OdW)AHGMY4KCT>HO#AWe[]IgU)PEXY-FBG_)8<Rc^]cMUb@QbD/eDQ_
b+b80:fMN03RZQ/SM:2eL/8LY[f=VUDWcFBdg_Y@Ga/:<G8_3?:,B4f>W,Df54eB
RAMYG/T3#=;cMcV[.36?S#YQ?/A388[cHS(9]C^d7+(.+7\FHYSA_WP[.&J9&e_W
=)>:1R<&c/M1LTUU_?W>K&(+[b6EX[/)H^O?c9MGMIH<Da2/8N2.8W)&fZQS^DKa
(B:REPJbCDSPGEJ:P^;1(BbE-b_<1Wb)API@dO@[6KcAEK/g8+Ad/GM2D9;KgV^\
D72T[Y9-W[AC,N&]S#g=<7O&>.4NC?)4c,/(.#[Wgc+CAE]Y_#d,A31/;\UVL?\5
Qc\^;4FMSW)#4<G]cG/-_c=FJS]/O2V#6^G7\3S=?3+?R#e0d?Y:eI.>NU;,XKSM
KI))L?BQ;C2/_KB=gT^#@U^WR6;T?R7XCfPKOHUTJ/3&ff:?5Z:JRY)MUH(JRGUe
7XOD9\Ff?R,f.RUIT>0K>3YKD<3;>_85Ag]]=5@5(DHFS9.cIF,OOHG.A\F=Q4&^
Y-RU;&JHG1HB,e=RTZR3g0]BX5Cc)e#&/KXM-Peg7ULCO^S=73FU;(]T9RVe<b4U
#W_)Iaa+^E;1fK&(E1:.MS?0[g63^2D.=7E26HG/RH94O+9#4?aQ]_1XKWgN5@ZS
5eaJ+?O,RPE4;5#3aEAbWBO]AF?Q^):Y^aAgb_aTG7X,[#YN,1I14C9R@g,STM(5
ca&G&9JGe+dV_2E,bVV19SY=Y/F?\-IZ,^UF,4MZd<TgMIW?)#OLc\,YbR(dV+bU
.g8&2/49S?G=&&D2T<b-bO:D=V-A#(-1VZH.]9Za#:A?07cM1JbfQD.,fA?05VG1
2PfYaS^MXIHNG1?_S>V>-,S/@&dK/BOY;&-LXI]<H+XdCJMK8<4^SFTH(W[\FYKS
OXEAU(:)@)-U^N\.V7VaP\(O,bFF4B=QL96TT8#/R/864/,RF_N0<#YW[KXf^-DG
XQNg:F<P0T2O+J)C[T]K.3ESUBe\@f2Wa60K,ccfN\CCaB6VP@<0.c[GPQ]3FH])
YCgLP/-E_@=GZ@Mb_+7/D0c15>ZU_-)3P8V,Q>>39LCHQ;C:/2,CVIe78#F]JYb]
Z]O/@F>KQP;3UOUde\3.KB5,::JeH)aL[<+2I5FP+WM&_4@4D>?M_RD?&8X3BY[7
A<U[&I:YEbQ5I##e/5cI>/#SP:A)6Z7feY-T+-Cb>SAK?Z#&[YV=CSRW4<?bQ9I?
.C7B;7ITV4>X=6NL,]Be;U&LEV^?YD&XB+B,]000VR;eBKSX[dSAY.FGEC7d.#5?
&[/-U2K-W].6S+>J((2ZXKV=VEE#,2G_0;d(KC_7R3KL1F,2@W,e.aO6WEZ_2/:b
=dVH+PBG]J/U#IecCC?C_/V_D<6VeTJ-DE)V84fTa,&Z,WI<T7d>5J4@-Q?TL;V)
d?KUWggO]d75a0U9Xa50P8Y>cgf17.C^a8CefTI#U<)&c-XP37a_>QIEa3YbQbVI
JI_<JA3YZHEW)<##CFIWE=P5DA^5<LCPG+F-UcEP6//:#c?:;6M=>XB2(;D-4-0=
=BRNB[PW@:E]@WfcY3cc8=_Z=\#e(])-ILG@6/V[;NL8,<VS_])18M#,7^ZF(BE5
:H&Z1=BZD1:bF30?f18]RBELfR(693_DQ;Ue)UKe<X,<IK._dGY=ccO7E.3R2RVZ
^PAZM]3-e(0Yc_&-]d:^?W.T0#bB:\&[>&3#8=)V>&?C.B0:TH,[040(b[.fSGfV
=QbK^a7&._<\-bfeIQBJSUY[E54Q10<#(B\]cOZ;c#UPIJ[3/7U?e3F15:R@E(bZ
GXI.LYb6RW1XgT=+Q0>0?R4Wg0/.I143,BK&&Ia.W/GHP>]MUINIT9[<6X)C9W,U
4WFE398^eQ#6JVJ??OOQ(c/6eC[(DV@8[5[=UMZT0^#^]/g#=95QRWfB_?A^1A/d
I(Z@@P6Z[f\)eW-0CI7B_P9C=B98IRV89?OWd@f2;?<(AEWD:TT04:>7Q],&A+Z;
9M_d#eS28:]\EUL=>X1bcB5;:b\Vf=OA)\&aPD88(g.,UM\PU@^QW9b2@^KEU&PL
:-QEC<@)@G_L=YbHQF+g7#(N>>GG-0W(82ddL:cN+25#W1OOKHYYFQ+E_843H_Ea
5&ObRXR7>D3;8QgO\3\M;(@?;-[D&8@T,^LJ)-[YVRI+H7bbOC/XabX;NX-+[:)>
[61=JbGe2).O)RU]?;cK;09U8-0>.S2.eP@S#fbE_(bTWQN.[_P.Jee::)IfG=&K
CFcSd?KeH=HeZO43:.(8RB:<62P69#SF+])U:CA2gM>JE.GQ<<\<2KA375,Ed,4c
T3..#R4XIWFH6WVPG,Q#N]>D7DA@<(0AWd?[T@-FdOLA&TbQ77a_H:BX1\\&K2QQ
<;c&M0R^:B3_RU=&K94I=\TbZ2[GLMPY@(Y@_U\A<D7f2b42C)eODE:6g@6-O5.Y
Z&=1a,S^IE#P\68eHRXX;cM;[/g,/c4=e&ZZY;f1K?AebV#=fGK@AWRP3\-:O\[g
?<499N3[;1@7Ne-a-D59HO[^@KXa7B8RODe:/GD,_287L2P6;(2SYgV;0V74KGH>
3KV4B.a@QXJZXVII1ITac#+J=U+[AS7fL8XHa\TE-Pa65&OBU<DM>ZY1e0S3WAUP
28:?McLcW0/6WPWa(R@K=d@(_Q7H4&a->;0d=e+VBdZFX&IXLU)\E99IR]]aY-X&
a@\WZ@V?<]^S<IFX+d;Ze8Ac]8A^:F@N(>J40&<JF/Ccc1[eID?#0,dAa8/+Y&<?
D&RENOFJ7\R1-:=(.^4[Z^N7;7[?[a(><HWN@_L_6,CDdR:H<cOcTA<<6+EX];C<
Af.\4(g?Z/ZKH8E<R1Z@QI-F#fBIeB[FSEC/7EL/.[0Q>\>5KS_N;J/-6Q/=WVSF
)eT_Y1<0K(R\9816;)Z_+0.J)(Mc0H8TP)O2,_/KfdA04>QB5N-_0#S/>+=^DO67
;D-ZZ4U7J2U;2V/ON?0_MJ?]RL@PJHM&]59,A+cY0V,\PGFJX[_e0T4R_@EF-eWA
)1O]V5V(=PVQHD6CP/_R,B5:YJ-c-^:3L,;N<AWKOBe&5[(_LI;.=9)?I8NNRLP4
H3#PA?Sf0[T--Z5b,MX>TI;[8/M#L:L[^+bMb>)BKWNA+KRY0FcOW_?@E?(D,V\1
6FZe<#SAKO[8d.S2gcIDD[PHA.U<NGZ-:]b9[,.Aa.0K=<Pf22Z?^T8]<;AN7HZ]
^>&?d\FV2NFNb(E//C=A8@MV?6]]d+Y5YXUY@^_8IE?44QO+eF7CBE(DI&f<J#.4
[#,3P6-C</.C(FCa&g+P+(ESY7EP86\V>+7DZAWHBIIZc?U:c><W<QR:\2TAW^gO
#[e</[N:c>PY4&)c&2SS=(\-/W-D^P[C010MG\H?Nd+[]<T=Q4KC_&OFPJ;>78MI
f=\cJ#V=Gg?>+LQ3d#A,&1[5;--UJMD#-@1_:#P1@c4+X&W[6]7Q\c0\e7d;_IVD
3;ZF]OSAYUb\SCcJLe:78VaC7cUOVc4,T0O>?CNEAc]G4V_0_8\U)PVBBY;5/]Tb
./+X(g6_8Hd0N&D[eD0e6V)IV[@R60(;a#>(@F1:JcJ.UGKXV;?1466EM7F@\aHF
6?W):ITZ9,=eVbA0\]f?EU)7NLLYWgVcAM]N>X2Na8W1W&E#B>2\+CTJ&V@5B=\[
B[+WTMYX#B3gT.MSL6eXE=XMP3Q]XL&EDZ>46]&2Ee_V9CH[J-7?-7(69CYCW5>C
=>NUOgE=K6)FEEQ^OYAF&RgILG<=1\U^^D&JFG+fa1R4.E&W,YM>@Ag:(P3&7QB:
5f>_HEHA(8+5Q#B>;cFd6Fc>NWM2,[8H_1T56-O:?G)^YYQ_&W,IO/X1c1(6+,+A
PB#:?,T_6e.]M9JJ7IBa(3)>QUVcFcLc[D4,<S05EUb+cO?D=(WMb#2[e9&ZLXW[
F79C6>5TWW[VYJc;@1c^g^8Cf^C-U5;?&J3[1F6J1G[<>MQ6[RGQU<,=]##?7JRL
9:SScQ-#2J-:RGKc>;GgIXf4-Z(U:eITE5-X\(gBHFR+X<Haf_g[4&IH=CdO);Tc
eHL9/&=4?DFa?L<.2JW8R6E=3Y@bg2<DLNT-GR[Ce/bc<8ZU>M9<,S)a1RSJ=)>E
ObB2D/edZ^I3LB(=@T.Wc=Q/@(P]O2;?^R?d]4^\/H7;NF=d=?MBdeEUIXYD1(dA
96E]P7DB]@/;d1S?/K16E=.U8H0LHH1J?D^3f^bV0:)L<aCbX0];HF^HDaZ-[5UC
Qf2&#V1bZ+NW8YKN^b89?6_U1gH]a+4da^Y8-c4OTeUK^Z]@?M;TVYGBKQFE3;HK
5BeS8Z#MJ;dbRO+gC+OaJ^JB15ZQf,0d=F-,LPa@7M8dYVGBg;(c<L(WXaeD<;S;
/7)B//,:eUSRAa5R+:(^.[(H,E&A+bL3&PKF\(1[6\9WHK&P<D^ec?Y(4S.CMCS?
B2DUfIPJ\UIXbdQGe]Q?YGg91&)F3_B0eF\O_;0>7Ja^=CWTH1\W[>f)Y(&IHT[3
Ne&JZ&Q^S]+X3)?@aVK0GL1#SQO-#W82=/991=gIeMAV3S020^_Z5:QB;F&L&^QI
AH+(NPQYCaT)O,L_KNAKL9NR/]N1;F::5O1AC9H?H9TfS:4LUZ3.2LK3C?:8)1<b
X(\Wa1F<T_^]NRa-BG-Db<,:-F/cacR\XFH+^6WP.-,PgF=F[K&b[2&b+<AA9ZeT
:47b@a=V6B)[+H4#WS-4eP[67:XHKdS6^<ANUe8dIP>+:8f.ALPLK92I5QH+QY9f
_::6KVR^W[VgG]>#[&9G/&+acV\CCYbWJe4dFB-1R.c\&SOM(e[2&JbKMeH79gYU
T7c+Ya/?<J8SLO2)+7MZZ.Q)H-#S/#4N39D__C\H:eZBED)Y:H8LQe9WgH,:fZ9N
.Bb_J?LDH4@FVWF.?B^3_.O\HF,5BRH,+G(,BG8\\8>TaE^BG0/11;8:gc[NR+g1
4VC]./9WWFg^@_Qg=N+)]KGS.R=1H?O^g^6D@V7&Oe:cGHe.5&YeO4>-@R]Q0aS,
#^9Ke(7XO#Lf1;c/2:5a_H#KE6EbWSeW\\c]^?:Mg&eO?(eKH9M>ZR:H^Ca#f2&Q
TH0?gPaD:,gM/\\^=-1aV8M7G0(3f(,2??O;,b-O(^>]#.4PI(5TG>ZBA=cA6B^@
cRYFQ:a/FY;@]V[8;4W86UN#b2g6Y7=[W]HHNVOQMa1fKaO3X7PH@Gc_SN5Bf;]f
1=5,LU)?Nc/g<:9JFKH&/aRQO\B-&.(2\aX(OYFR&X>95E=P4(EBKW,EZO#A7:]A
7dQEUBE.,6G.7_7+E8\Vb4NdF8_AcbE:Y#]3.gV.>5ge\9KgN065;O.K(Mc>dWd:
BK)Td0B66P9?P460007L4-ga/?ENO+6+24NUM;(99_YVH0-P/8<O^#cN3S:J<3NC
4#J>,-2?<J-8b@NLZ2g0#dYU\O9e]YDUJ=)7H(c\2N-bTADZ:83XVK,fC1I4C.Y/
\FK\V,MZ@>e_CTQC.YYaH>Y5fHG4XYf0;W4;VY[0N:25=IN,HY?#<1]?^W-P3VHR
G<<-H0=;de>.L@S#B6[UJ7UGWa/TcS[3@2DFLQVTK)a-BUg4DM+S/=[9L>[PW,C&
A)AF<=#A:PR&g1+?Cf/TeH)c.+?#8L934J9+HP[L5ed25=V8\UXS]/,cO5@1-KZ.
>X;J>/cf<52a\@;fY(<\[Ig3ERa0NB,_8/^;D:5)c)L=<(#GR821Y6B3OBIe]1_?
J/1fR95>23A8-F\S8SOD>X(2aR,X(A_fJWg\5:2f?5E[BH,Q3R;AJ>gPG>ZDRbJA
<>#GTL<(+L0F0)>X7Z38(cg,gCT3CR3Q#D>>EAFS:I8EZc<>C.(a@?9/]A331+aC
BZV?U6>XZ205BQc<RZKNGJ9VgC=R9QL9(^>I9ND?^FE^0e7;dc7[MHd+I7RV[O@I
J&ad_21g;\>\/&=RF_+.<;bSAb1Jf86-WbMAd<D<XQg3L/+Q9@cK&9:NB>WTKJ)g
GA@L[9?]@#NaK+.^1A3#H;c_KP(YeEJ^[\\T>fa+G,FW+.@0+26)B:S0_O(E_U3.
DI+/C8&d.JXQVb7ff0[D.JCX6OM_MF6[A0dcUOc73[Fd.HC7BB?A27^EARFR(T]/
+T/#Gf@KT2@PU.G>)E0U_dJQ=XR&@G=?;C(\AVI;O=dTc(KPB?)B@J0#,BEE]1D-
XX[6V6I068NZN-:6VC3F6J.[^C2?=_/E7>[C,L,J&\/R9bPA(+9&K8;7/)@+<Ige
T09UVGc>Zd>R3I6dKf)Sa0OR&__fD@=:T/N5K-4(PY9-KE;cb?S-:Qa/0F]I<28.
,R.9N5O-CD(/(I(YKdVJccWD.>U>C#ZS])V+4(^c=U/&6a/X7RQ:=RL79.-L#L@6
4f\8CWY/VGMP\T#Q)R0:F_E8d<]K5>F+OFCT#fD/CDHDQdFD-Q[gOSK[:>&<4S-)
N2=]ag+O6LEH+=eHdHLG.F#\d6&60OA?d\Jc/\;GN2I1-TJLON8+KD1.HP+EGBcT
(Z+2&;d>f+FFb/U?<7C-SS184BT#&:ABN#27G-/_cd0]BOM7fK7EU]Z6Q/>G7-J1
(CH,]dYWa)(H9U=(Z4V<f5bIdXYK>+ZCf/-QNAN2L[e.\RXYA9/M2_WCL@U>0O:O
C:6beN[NP)@MQG=_\LR6cfV>^-+HE?/c0LC/MAMB\M2,;N4LGZ#^fY8S>2G2=:[S
;\P/9-V;Z,Y4J209?fHM.bJ9/<\R@d<e-[DIeaRJb0718.ZE5[Eb4O0I[Q7Wfd?>
GSKIEd:cICZ0^<Ud^7PXTdX58#Qc2-GSQdN-BPS89__UHT4?XT<a787C90Dd/ZJd
AF9DGc>^/J;I=?,AD^OAAXJ=2Q>(=1IV@JB+abQ(+?FG>AT;=e;;+4d3UJ26_C@;
5^R<;NWWQ=8=P:JY;NFPINUZD#\SD<Z?^1M<YV[dM,5KGY<&9(1RD/dWM+96,/Pg
X0OKc[Dd;[@37(Fe-afT_)FNP3R8X=1f#fCR>g,4Od2<:>bJ4KTQR(WM7;R(c:_0
<#9^8;8F\MPX#e>-Kdd>R[-=T1_Q_<&75g0BB?W=cKg@g#_Z3)gc4?aC.C[RRF5C
,3#7bD;HVEI<25SF:/V90TJ+U^Wd+J&(@.X8Sc9f_TSMKU_WIEde]@;/#OI>T56/
51I/6VL[1]0#,1IP;)>ZFfcdcZF\#[UVJfC9D)O1^5F0aZH&YD;UaU<L.7;WGF6f
EISUED@GJGU#]&g8PQP=^V0G^L^;/^RMEbZ7]S5<8(;NOW_0(Z-T2BGT8FN1MY];
OA+IGY_7A=eL&4IH-R4^Ua-GS8WSN]65ZCL(=R9?Eg3/FcEXd:KNE<+<TcJ8bW.3
b>+TFgD3F(5V<TU8a>DNS.d=HTSdd89A6KK_]P43Dd3#W@>NSNZQQYV#Z#]7,:OR
De,6X0X(@D.@4Yd;O(NN--KK5+cQ>3I?AHaC7a>MT-e25C,O7fYI.PgZF+VOGc1S
[d4XWfH\F)f;:A,NPN)V8>9,2SZ23;XV,PG(7Q0deT,ZNV,(ABa=&4V6(-e;M-XC
913-L_V9W+4(UdYd1-TBX&g.NA,L0bL=M2eDgJ4L#13V35DHWFCW=DVIP3ATA(R=
:73_[#WK&?9GcW]+TW47(4UZ?)\d233D\0_[W:<5;KWFKOSRS3#)[=S:R1e:(XC&
bP(KV>WD9c1-fb2);#NTAPW+c#=PG&CV=F??O6&IGW.WDZ]2XSI2Pec5:P_6,M5:
HJb:QJL^XgA(.;C<E=H6B>81&G>gP289;g]]B,SKYGWC.0TAZBLPW&__UWGe(PN0
Ic(dXYE;^aQ33f0K45TCUNA5,/#;F.UN6(77OcR^G2IBH-3?#fR)M;/AX]KeXV^Y
ZFgAMB?H&CY=>;-/Nc=EHH34^);11LH9EP1KfMWe9+^b_(,7^/TLFMP@XNV]NOg2
,@fTIb8E3^49gXMRF>,J30@^=/CI6ILSQBIIATdd-9=:?4(Qf&.Bg5M88be6T0RR
F:#IZ2ZG]G:OMVGP>?[/@6>4(LQS2D?(c.KJ+=CW#&P-MB;TJ9^:Y)G>f,Ad.(4S
(6<Y2BcY&.#V3[O/0OPX0DRbZDPYST-(6V<W;_6Sc&Q_#O7E542KOM0OE/Cc]a(K
=DLKOI6=0\T+e6ZPA.WPI:O>EaDcdK/9S=W85@eI/6O))[UCWR:dG@db9f+&cNRQ
6PT6D45IG\J?g67#Ig&_QXBQ&7AeC5_1aDR@TPaPTY@0B]WZ]baa=UCCV?\+R/Y3
T-d^eF8ffA,;(<KEIKcc&JMRYJ8P;]V#G><J++b5@:]WJWXDJ(=f/:6f2D_dL55Y
JL-;;4<9AcP97NHcQB4YXKbO?(+65#(?&P<QfJ6#0_dMA-K\ZOIMVX0V\JE1gK0I
+9N[W5>E@KB.Mga61XVV9O1bFUC5B10AJaGB64[Z[?]I=c3#6G8MVB?6-ZA@HXf6
I++59/>Y/T-d?K08&@cB>M4d,EZT7<6VgC_W]W[^c\D_U#)A6;AU\@VbD9:FU_)>
_4bN)#E:^;<>H3#GS)@SgCgIG?d8GJdW^4>2QN2Hea0QBZ7\&OA&a(+T^IW9(S6G
HNPA66aU]&NBdYg+(8&UD)<6)f2H\5-J:N2T2b\L;7TJ<d@IIP_N)O=17e3DM0>0
B1CX0X7#H88,)/^:eg:eB2#bXC:fJBC14fXGLDOg_:.?J-N2X23#H(&J.3\Uf.fL
b\WRA7/LGg;C(=)1/:?0D475S_/A)OD9)a_54TIO?X1MG42[B3LAFg0;+I[>Z)@-
Y5N,[6EOG40&D8/JCU,g^:Z=,+&[9E/dE_D(ee,J3F9b1^9:<d6TVF3,cM9LA>V7
S(E?K4[A+OGMF&M>.,B-ZWOad4QJ6RSYeR7(W/.Y3>@HJJL2ePZ4:AHV_@7]Z.+/
I?V8SG@-+eg;-[eDM_JJYC)5>>UeO-GFB@:;BVOH,&1FRa4[FW\:,10<TKKLZ)UT
UbVgSa?9,GZ&Y91[/?3L7]SS_M+_P:F]]S,1b#eU16KKdf[B;2KJ?I]\bEa4<Y8/
=1?A(gZ07XdVAS=f36.H3gV^W/RD6HgIHf=H&a1UGBPEG[.,B)cTF=9L52O^CQ0(
F\LKZ+3FS9S.\80>>-&dV#E;4We8D3//F3BScOXGLePF)EZ-/;PMM]UMGP=/MX,Q
3#11)AEE7,2e/g7,(8MGX7L[DAMX=UNVB/RL4POV\Z<af4Z4@6[B4FJ\Ge8?:BV?
TWQ9&;I0b,g19R7ZMCCa71#\86Pc^^>f\^6F<Z8J+0>.[)+N5c]P<##+ZP<UY)5(
,J5ZfAUK8]6?gAGP2MZAB4._-I=-0PgW@N-Z;VbgF@Ma+,B=g^d,d<=C_Dc\-W:^
)JNdCT]ASU-O]LCP:HVE20T5]NcV96L8NW=O^7Q45[C2H6>(\M>g-D:bA<D+C@O^
1N9@dK(HVE_H+KJN/^(-KTa;;6K#Kg1.JYbXX.=XJ.:8M[eeUS,5?P&L,Y;@TFb4
CL^ccO=#(45[.29;C(LP53D266ff<[X]?TRcM+VA5)5/Q6P#gWD:)ddESH[VMSM8
0[FP8NeWFY69c6J5VdYJ<WBD2+1BM5#0P3Zf+,U1\;WaUR+X\R@H.D)=>&PH.CC>
Q:fY\ADN0[N5R9U-b?O,]^1,bPTd_GAOE.SK/89WHKTcP0:b7^818=UFR-PVR\YC
a89e&c:8H.38?MV?OK(d(bRgWJR:>JB(4T_YSFOHR1QQF+JJD_C:&?T88E=4LJ7Z
,Of-U57<cZ3X0(@]7R<9#_=7\=#<15>LF&YL<K4<??gCLS<V(76G-fEP.(>Z6BT+
?5L-L++gdS/3,C[5WdJbEFF8?DKbQMAO..bWV5Va,TX_Y+JC7K9C#[T_F&K8dZ]&
I^QYfE4,>W.YHEb[^]A,9H68MQSZFe[\dQHUF+-IeH>8SUCPET<bI^SbU,U,Me7F
?/_,[^<07+V0Xe&,f<N5\V-NF(/3&_^H^>9D6[PW5JR3ZDb.5W1X.F=OM-f,&L.)
fWdg^G?GJPYIU8@AJS7N+Z/bGRe<)Y1QW9#Hg[VP/&6[HLN:DHV&f==ARY5HD]K;
(_,28.5ZIW0/ID^NWc6dM_AYdd=]D,K92AR[;Q]gA\R/Q4]]Hf@]+cPK9e3c3G_L
T<#Md>c,-cGLZU6NO,5be.DZA>@JTX&DN\Wb3(O\7/Y:Y@GCga<6V=FL//XBM.)6
6FeRU?^HB&=1119)^@TP+fM^T;[GZTM=#?dUR?IFN><fPKZCB<@C0C&/g1O&((a<
/g?U72E56NKTCd5Ccf)7\89;1e.RSDR)W7D89&f1)QRV/1-fPONDeVM);7JC#]/0
TPBJAH1WcP,_+\>bIZ8+M\?XH4TbWJ<.YX0+eM#F0\ES;-B/gZZ1OF2aV7dUH3MO
S@KK[UJ;/2:ccDTUR3_[dS>b@[FU=U@6\UI(g-#_5@[beUK@G[0fY_IgHM1N(K;+
A1TZC^T:CU:OO=&WLW1=8I/F:Nde>:eMTP5&8/F8LIKM.#YVC?.@?0+=WCZ/_QQd
b_6e@+1(cE9de88aVI_Hd6+<7QO^H?Y13U6fZ8/9fJ8Q9Zcg8:Z\L?9JECS:I+dO
K;eSE;QG+eL-,-BX;X8RF0L=;+?gB_ag>PS#LZKK?TA(OaU#;0g?_+[fE?)a?5<)
#62,&4Y;]:UO82;JM463#>3f9Z1.]1g.X?4aY9Z5feVFL0WWD+_dD8HJ[9/g9G@@
_@-PcH-RD6B@YR&C/g.=-A5CIP[^8df:U;+ZS_D)7Zg1:7g?UW8,I7.3?/T-fC07
BeI4RMQX9eS4aQea-+UK_>R;D8V/8=DbT60^[E@&[CbHT[e0Kd/7[NT>G^=2NDdF
RS.7+^73;UaM//a;0?I:#d(-d;L.SU0XVQYP0X\E^M@TA;fJ\(1J0LM66_ZJYHC)
e_>MSN9O95:=&Qc/c98]6L#ePALOL^g1Dg6_UT3e(0e:QMd9a8N?>]I]Vb?,.@)G
7EE0(CLd:MfY^IF5[@b@0e8;6CGS(f[a-L[/DB<>L^b56_K))AJKL^D2S>R?UD1/
9C.8>e5&e^&FNJA,PAgf.G2;[+F=aQ<gH\>,G<>f83=XD9RQ;PVIdLVOb7H@T.FL
W9A@BU]AXF3YI3gP@MM_++52[<#V_?B=LVOcKQ(DY[N2+KY/_^=1)(P;d&I_QZ,U
LO/9)>J1W8bUWbLG#G@4W?I)/G>.0BXL(?NJ1\c.g&@V,@I+R6?fU;/7G]HQ_(+;
0@Ka6WfOM@:?#OK8=c]:;QTDHb)ec03]\)W\#F)JT7G-#=UE[ZPBX7[=GI,:15\0
47XO0YX:KCM:F+MfHNFNX,<\=\MaJBQMWZYDNK#H,A8@EU]&]03#Z3^CS)_?ZDI>
GFAJd0:KEPDCX&BFG[-OcfEEL1J)3?A.VbbdE@5fE2D:N0DQ&gP49R#O/;;A>J(]
9JUeP:P\D[Md5V&<;1d834)DO5S)>PG0L1Z[1_:)/5(<38[)<(<^eNRM6<6;:RA^
[@PFCXFKK4c:)<YCV;He@R57BPaAEQWHC88QAY0D\]8X+#1:FO-Ra_7Q208ZH0G@
6@d_A[a>BS<RI(KJ#e[&eIcJV)D=dT?@S[B9TG:/cQR)1e3KgNX97GeA-IHAP\9K
,2-)3>+Tb3\#1=)J=I9d:@0U(B1Fa\ML2dT&MPN/&;=JMPVW]]TY>2^V_Q)XfQ0e
3C=Y5-K4)N<@=8M38ND<[UMP];[-O?JC;GK,GC/WH6X2>d6/]DbR:<<bE7YF.F44
cDRW1+CV[S]L=I\_b#07Fcf&(OVP/b@TBg9-bKdd^KONN>JKD;E@B-[/<P5X\@=H
TWgF(Q-fR13cX,,]-0\dJg/ag/,,J>96FH.S8Q71&/fR\&S)ZJ+f0[MM0Bb\5Gd0
B_)N#<1[U#&-W&FQ+a@cJ7\<GP-T:4Tf@T0QE-P+[IT05/L=VOTW#T-PUZ0^cH2,
C1,Ig&WCLH>b-8-9@^Se#fY[F:[\)8?6U1N1?E^Nc@3/dRU<FeOO+&L>d>I;HI0E
/DZ>6<03PP0A0?fJ-8_<>-)DdFCU/X&2e[N6NN>SdFH9+=>dMPI?a<(^NXV6YHLK
Y+&X>.3W+c]SBPc5aX5eWLBaMLS5g^C,7-[-:FgP\_AVV#=EHeV7e^KB.N:[@Ld/
ZNKD97VQgbgc?DFG#G<GXCGEAQ1>K@BCMfKEUMfQ(:e91M)IfVd8]0LR(cH^=YPd
YMKa/EQ)6Ia8(2.#;HeJd_ab016U#;gOXcb\N]RVX)gE>]S=.Z8Ab2e<OD542fKT
(9BQLZF-^CPG]2+.+[+#DgFIZ)Ce8f-#Bd13VH<d80T#\@W/Ad<#dLOfH)C@=6OU
F5K_@FgTNG3aS32d4Q0T2=)@Gg^@IgL>=9G.;FG&dbQNOU#/\#)WEPLB<;TC_HHd
?Z?JO0413LY07bQ^1.,;#C^#TCK64C+1TXC&cYDgc#S1V[=e+3YgF:NS:A0#NaN:
THC&,2/3^B(V(..c2I+A09FAeZ)#_9G5SXBgVZRfJY0-59bZ:JPKG;FZVa,R/\AJ
;V;3KIQSI;51\N=)93;DVcOF)Y,\1XNV:8]H@],_9B4]JA/<eaBX3b&Fb7Z7JVOE
,,ZJF0J-MR5T>1[UE:,WfW[dFY_GL&A^]_Z^WYA=Nf:MG7MUeV<01,fZ<NR3:eV<
3e=]f_PZ4@ZA;?e&=HPV[PMGPe-N[f_E4e@9+F=/d_-8b77[CNA_B;e/SMA;CXFd
JG)ELZg-?VfF(69KQNZ6IQ.2XHZ<PXdY,&eSbZa(/_60##,-YcWe7QT>B9CPLW0)
4JEO_+<J/](_>#RY,Z.J>=Tb#bZ=;7W@=,\ZH&?ZbaXABF^OK-(KCP[GC:PY83^,
?PgGJB_I.R;ZW6[A(CC(QUHZ&[(6>>,e0ZRY:RE:UDP>cY,[[X#Q-J8I)I;c77XK
a8<K#6B\C#OD;1TO(P2M08P)M]g?>HVQ&4?3H=@>[8-<;=[4YK=G[3;)BQ4c3(0&
66(O8U4/H<dD3bYFOIUSd@,LWgTSMX=)1bXRYR85>UFUY=H&JFfNYd-N&<53X9BF
D-LWgQCd6LEA?JR6(MQ.H<e7eV7AQGRJ9LMCW(5;DJ=AJ1BQf0eIfY=^?[Xfb+5X
.OWKEf<#)Y-+1]5V73D/IfM=0Xcg>@Q8=-OUYP8PG)Y7D1GX[IZ#+Y(-e<)TYJ^.
C][:e5Y_J#Og:3)YfbCfL7I3\P/8b7^>\2ILJ\C-9(,-:5+X]#eFMg7DQ/7;>.A0
&V-TVO:3NTbSKc+;.<XP/a;PNYY.FE7C0&V6d<VD7G&BLS[S;a3^(S#J&Pe:5M.a
1<Z7O..(&CGWdE4XdP\94605S2BgM1U(2@20QPEJC=AJ@MXV/.9UgbQd_77U+^P0
gZEb&#d/#7E@(7d<X=BL:NeAPUFU6Bdb1:1Dbfg9FR,S4:==HZb(:JU\Z[6b=KZM
(fYP&c1D10<##NLc[4S0)HHK;8=g#C\4Q?#M;XA;=:R#Ye+<&TK8&-RGB+&)AaL1
S?K)3,&5fG,-H/,=P]90>?)9]5_gPcMPB1R.GZSL22.aTF/I-YgZ#;2eT\2/+1IZ
J-Q/\Z\L@-G9b(</RP4ePH[^5f&VJ7YP>4/G2AJWZd#2U^L(J-dI7K.d3SHVcUEL
,6eb+-+CdM5^4)V1/,@:\U&-b=D]YS5@Og=DLD&T=[d#]?(CQb#0B)UN(30P<a.@
-KPO>eQfIfe=A.(OSS_Mae5H>QJ<>Q)72?HcKG[F?CBC&XYKJeY#[WQe8bL@3fB6
M@/2#O\MJH#INM/baVUP#R#+e+.Nfc4-@?(T_4b/_HK&a+>/(X21)]fEOa>/3N@W
.b;RE<AaLWG;_^LI[FRB9fWEIF+)LSVTP>#b_1E#8BKI8@P.HECKFa03FTOTOM2K
P=P>gaHbBRS2&(.QHHH[BHXDUU?84:.<OMT7Mb:gReUSTcG[IOAJ+S5&HZA=N.#-
\@ZTL_X8Y_@;2fBIBOZe@7(C[-Q,2.FF:[M>#I0]A8-25LCL@W3^)LP+@c<F4KU^
,&C5]#F@KQa1+c@2IXQfL;#D0G^,c/@^LZ,CZ];J,JMe0-JQ:_<]RGOCW1_R,?^C
S9fD6IO)H1:g[T2A(F@KNS5[9YU7FC=b#+BZ@?4M<3,8)TSOg#F9;2?O/NN79T[>
SgDeF75&G=4/Q)H@2^,S>P)AS4#HS0_@;HUK]DFJTV>[<99E24&F=CV#?Be#7b;K
_:;1MUQg1[4[8FF)KKA#GZ]UV4#J+D/g&66:VfPZX5)J+d>?1DZ5EfD4g8&,@=G?
3FCG+L(cI-\(d^HXA[O==]5P#_7g^HL-e,EC&.,[d1JODXbUObbPK[L?V+2\N-X3
^@2F;dTU-\&)6B>5d-EX3bgEQSI@MFgAOF9BdO+7N_?\6,)D#U)<2>KDE@Xf,,N1
]HA_e9^RQUI)L@>&>O[Q0^P?>XVMG@Ac;TB5.)be1[B&;<1_YNKTWgR]UKMf?-U)
fR^Df+K]?Wc=/Y:&YL4#D+aJ[(\GH;A@M=&?Y9TKb6a6EF<>f\J6=.c0g_f\@/U2
Gf\/Q\<B@[[@X6PgTHUa&0/U_Q;a0^^EFX)@0ZHRaH-cc6G55)]dIPN)X7P-E]C&
Y:gO2fJ,4G?-ELL@G+7a>>U(L5RfF]GBZ#OJ?aFYLP9e>[fBfD#?]E,cG?aRgE8#
6R/O9=]JWZIM>@<1:E]3:H^U,+]K8gOEKZ.Q#[4N^=EcBbO^Kf6M;1_L&)-7:AQ8
3Oc?f1eDA,^O1<&ZXRSA#6eP[=U3@-D#BQ&C-.:E+.A:HN_O+KP3[.fM0e)ACK]4
OaGd=dB3T]Q:e]NQH3Edbg3AX_dO:=XA,0cdUH17^E3>;-fcX[2PJ,>>g0T;7Zc_
N\DNbaCTO[U2]b;aJ_]7^+[/C?-0J\DHdWeR2R<gPY&\J-d<78-ge;V@C:Y.f4[[
28G#0XUXfcIX_/VA]>RPcW4A3.EU<#B#UKL6#7MZ2O1==SWLZ?F&J71-+R1XUAKK
.;B.K9J9MW@#X=H)fJb9+4ZL_6E^FS#IWEM>RP]52O<GY(Qd^\Xf)O6,8WW<^>1M
+:[IHcbb1c>;6d=,(W&G^P0Dd]>,2?,AcZOB.9FCHX_J,16?JG+OMPaOIFDXaUB&
X9#.^HSd_S?@(QYUfASK:7<X+BWedH59/db=QV8aRa03e49A0S=KPG;-+eJL/1NU
b\9ADacCWYXe9cDIEaZ64,=d323S^X3C)9L>,OQ9XH:AHG5B2g+#dLL?,EA^6f__
9Q?a&WM,ZbaH[AC@5;PO&4V1[a3Z-FFaa;J[NXWgKD=_b)(FJ4L-4GGO-[;UX]=I
K/?abQ)Ne<]GdO/6P>FWGX/YRE-?=E]4^A\?[-PU/I^2M\b25D>I0<A9D:bLSOX>
F47DGN/-5Vd?=0)[dd>@aOV_bZ.8VCE)>PQG]\U5R?@VE83O^_N/BI>UI5dX+CY9
>ZRTA@&#[S:C0^a74Q=PX.DP(MCYJLN\26]^=:8B?#5NY7.WK4LV?&8Ud;ZOAf[=
_)UEOHSYg3#A#:fde;&J=XWUIFZ>cc,1G>;W=aWJ[L8OC5X5c^,MJOacN+_6P0HL
.I]=b\Z-87NJS[V)C:B]-M(Y+^:R1X<8&R^;Q6MV5\VVTf)G(Y8+@8.QI4g:fHP#
6(gSY-7b-SSNdaRJZ++HZDI+H/3f,Na\N?;SF8VBZ(V<#=.YMX_U1-:DB,fX:fRg
TF/9.^c?eHR><\ZG<E6[]P8gT(RO-9SM?WG;YK7@d\I];LVLfK1.B_e+=<#CX919
0)M.I?L_/770LT^&0F8GB?[3=_;ZeAcBKH?<NdXGBC35SOE;)A2\KbF27PCcbSEV
4(<5,SYe9K4&W\865]F@ECM.N.8DM3.-N:B@=YO<+ag<?V7[JDGVT2f2R/OD7#][
\A-2+?2UbO8C6.VdfgO,N70aK]&J+gUg#<[>OF80TH6(94R><6fUWY^1[CV]HDgZ
M/AD:g5#734/GQ-R\#\RJC=K@M1F;5W&Z[6b>dWRK\gD8C-?R-;6,VPITR36aca2
gT[X\9)OT1ZaJ8G\(7HHa^JRO2(Sb,#6D4U&deHZ57;]gZIYNa]XXecJZB7L:87/
e\7Y0@Ug^gWZ.fBW;]HF)N]P&gI9Ua=+NQb./+(3IM2BUcE&J4>I_2f=gF5b,W@0
3HK&&R>T&L16eE82Y9;+>SSX18>O+.81:c\=:#U,4O+X<\Tc=>RQ++8dD0V9;0>U
a=a2AgJ#g=G)OPM(YXag==OXTYBI_I.fLBKb.A?E;LIb8WNSf0gC@]=N?T,dJ>g]
D\N?9@9B_W?b=aR+fAJEQ/KGGC9,=_CY3WBV:]6KO-dVE<g.b+G<;<6Rb=a#783C
TGS_<<NXCW\XUOGeJ/b4[G:(?]?TVb-HUJZ4W0>S6=Nb[X)>L+Vc.J^UU7,99g.[
eGZeX8ZYe\,.RYc@7^gJ8VLH]\.bH,1:1X+aRd0-cg=LB9._2RANM3+FP32/eN4-
b-#A+CS/>f12dJ1A?2gK=ZR,&+06d[2cSb&&+@9O/?cNFdU[13EF;<SIBHX0B;GX
aLWWJ0GXJ.Z78,^8M,:7e@F_A>WbC\B0E6EQdfc(:#XQWcINL)\1[1;WT)K8I+=P
VRJa#+G[H66He)TVFOR=-9g2HN6N^0S)-W\O&,aYaDKN0GVGD3Q_C;2U2<T(/VZL
JHBeZHf#\23)GNE)2<gNc15+NSS3aB5<LFU@#9_;2,5;bT0;4G8IWXfV4Z7G.f;<
KA4+,3OM4+MD@>bPQ,QJOYO,?BXXE51gLb/aTJ)1>B(+>37@8PC;XFVCgM5L76I,
>-),TOPG9H[DY?PI@HP(XP.PC/;aS5M\Z1BYQR.=EO^-=]2QIFNU>=?bVe[]_7E-
G<gLKQ&C9&S4N/3Q2K<J/[83U<UKOY?0gQdU<R,BL\Ja2H1PG^?I9V9<_A,#H0&;
?GZH6SPZD47X=A_e.O9RDTQ&7@Ya=(M>4a+5Bedf^W+9#D>;:]X]9-WX74C\d3Qf
\QDOaSM(6W(5+^Hc5:^.0KR@.K6fdDT6;XKGRJ5M-bL.PB_PQ721^VW/.Ye44L^=
_C@FYW[1IECRML9_(9UF,,fX=0.0QSTX_96X5fM#e+cTTJL#/-MG.7K9CT=O:/_H
)FCRBY-,B=-;:f19(>EB??ZfU<T9[L)AK(@R2Y-]4GIH25,,2A)+;a>23WZ3T@S\
:;7fEXTb8EbKKZG)Ia]a<&>Ya4,G8;OPXZ:\+fVZMF7T@-_KL)IS;G_b6:Y?a0PJ
OXbJAgO6]V=_d3NO6g4(5_#T6A>BgTDQFL7@6K&KBR.D.Le2Z38^a.RA5_SW&7[Y
9L9P]<cJS9]=WJA[<<NF.9K14?f>D48NgaLMfN0:?U2<2aS)La+3+5F+[VT#1JZS
?#FJA8G<^cFMJJ@Og=T-COFGHL=VY58#7Pg,P4;W5S?^N&#+Y&C8S-+\.]=KVJV&
3.[SDZGRLbA+b=IeSXg8<\0+8EccT)C3Vg#\W+\3D5C]edO4&=-(6G8Q(M>DY&EV
0bH&)R/-RW9UK9RG_DCDaB^BS1(L-bO/+L(8Ie.80\GZa-=?;@Oe6c.e^L#1>([N
LR>@59U@&\+<7f<W?25FTOU^D9:Ga\?HME81)=RR?(aDMH6GaYRb]Z>fLUAIHE:W
]?cJf\ZbfO_#H?E.DbX,9X#>W?G/4KfUBO2d0e,3N)cfTa#,Qe09-33L&cRH];LK
#>XYSeKbE@UbdeT<d:bI^A=G8Xg;(IA:34?[8;.ZM.@IDbGaTWX5&G(UOSbFMOV1
LY=c:7P2^dKgSY8(B((1&DJT111ILC4ADP]DKRU6aSTZ.HJY8D9>1b+G+a1ca?L1
1<Mf#GXMZDQ(C)+M>>]GEPfg=2YaKRc;>2E2Sg8):V\S,D_JGePEgU>aWR-d.T[g
NG(#d,IL0a3b:b]d@,U?-#551#g/3bW1RWFXA],>C3?ZCC/95L5e@[;H#S/g=FAJ
-VDM7dC-K,BaZA^YKI]f2:MMcO/SMcgF&(D+TK8.L08???NXG.QXB-177[/8&.;K
G5(?dE)=9>Z^^38Ta?)^A=B:+#W7/Jc0NOaQ6LEZ0_dDH?:A(@C.&bfO3XWE2d[C
8)<Oc3-5T;7T:MXdd9HZSK(>VIe#:0YFEDfM,Qb<-d9Eb#:TJf.ePSUXaP.0@P3N
@6ZXd.b3_HW&H?X>fJ3A/NJJ7RbA?(1U,4GVMQF7#?01-)]B59^0]Zb#.5](Q+XW
W43?(]8^-_ZF?(e#N?>[P87\gQgOY\bQG5_W^AF#:VI@PUJQ<T1]^(5K1+EP4;d&
aMWI4G2aK+FDU&bOAGI)4>dX:XC5a1\-5[\_G>L3C2;gSHLE67.^[@,6423.-,R/
,aR4eZ.Ic++J_(\E)OSXg&a5OK63Ff]]acf[-Tf79+V&9E45D^UD]cE=QP[C]I9;
&7F7GWe_&LNR=54F+=EDCQMI\c7a(Bd^bXLIX\:A/e\E[XFf0b<VV78>GeH.TB0?
7ad_0(aA7#4V1<\Q&VcU.PHd4\1/OC:6JaW-:KA<1SO6]KdQTN-LE#O]==JIAS/]
K3^/>OJA#MQbc.X(0#S//^4,WHN(&CZLB>6_<e8H4+NZ\<Lc8a]?+J9<6&[3-eO5
[?.DHR0ENTgG,DD>#5Mb:[YR;19HY&A[A/3K<ER&?9eF3\/ZGW&OT0=IJ3LLfT#:
A76+UfU#GG[^?CKT_JRBDacLRCV6:FO[A8S9:?g5LF_RAOBd2\GHQC86^#O>\[EP
<[?E>ZYRcf]fLVHZ\(dOW5_6M&0[@4&@b-JH4Ga;7dD+WW=JGSg4MVP#f:P?7V)T
/_/0&V35UX\6BM,:/PB>[R\(\2Yf=KS;VPIca6^)TLL8&B-O.7NXVOaVGF)W,M#=
5RA:V<^8Z=RFPe,NNCc>J?MEUG.>BHL#Z.eXceWGS--GT]a1OBA5/Q(8@E/4I_G]
KD+ZFYf)XRHbUR5/E=LaK^?D],a;N+ee]M/)b6>McY-])8CFCP<A5TcT=+?.NRDc
FN#d@VJ<OR]05>7\>3Y2V-Hc:QP-:R7OXe8+SU2c.^VI:/[TI=g5;NC;8/7JSI1X
N7H2W#ZMb6=PBWN&IQ]4=5E:T_=-2R(&+T.&E5QN#]1/6W^:JNTM>&dR8>PC_8G+
\3)DNfX>6ef0cY<M[\S#(N@gM+/[eecQ.?JcDgRHVY<:^6B]J;9EVO.JE_A>)A>.
ZfBCCeA[,@R-35S-b_/?b>;&WQc>Y]a^UF0Xd^5RP2Hde5X+Md<X^-&ZB^Ye#1(6
?+MRGgLE/4Y#)gXT]U&NN21>U:T5V71SZU6HS([H7Q,T)F-X>W6G<>+?(UQ-+YLO
E8f_SG)OP(VO0?S.VbUSGKD5fc./1:91T_III1.e.cJ#PfH@4@G4+B9X_G61]d./
W5(I682/:ZKc4_WA3:)Y.<\BK(C+WeD.>aa^=V@;P=?e?T)(I@55&WIZ[UPL1TBc
Z9+RF7CPS1&/S_(=GCT3?BbDC8dRC<)#\6S@\M<>F(A3EaaPHG36dfT7Vbg^\E]I
Z^,RWTHI(9>#^O(T.K&^^,KPR0\U/MXJ.dFRU]gE#<JX?CabdN@\gO,AC^W,)d4#
^2NG,Z+,;cI<+GcZ6L+8_S#SVY@V3[+_L/CDLX#PI5P23,<Z2C-=Y#0ag?7f4+7C
cIVdCc+;P?:gOM^\#M^Y,e7AUaRd=Og=_=\U@[:G9dX>N8\]KX&;T)Y^H47PDO93
Hg\^2#W;]gUSFS+W_e)(#,+/FS-46@K>?0Y1[d2SZ)HGHc#TeLdGU&LL[;KFc&:+
C8;2R?,^]HKAL1\5BULAPEOB3R)E[+7aNXZc#g@FR^5G^GKUb]CM[+L)\R:2&dPa
8TLYT/N)>6c^L(gU]M0SLeNP9:UM]=\KbWf+SFJQXa)>+11ALa9^8RA82=I:<gf:
^4+EYNLN7aJ@K2YZ>@JV#/>ZQ&X_HA?\FF=4/PX0Pa:g=/XHO8:HdC=dG>SU2DQd
-D1/2Q^bV9e9VdH_UEVZcH39(9<7T0PSfRS6<89g[8RPOJ1DB].7We_IJ;6-R_Q&
;b(&BIEENW):(1,@6V1,aP7C]TXKgO[717^WCF7f+^HGX.[bZ@#F<)1c)828VO7d
S0d@0YT?A7-7VMO:MXQT<\e58Og:Y)CFZ;10KE9A+G-e[gXLJaU1/VA6(,>,JP);
1Z794e?,EKOE-3:0d+\724/]\993><@a;KE)eZ-V.,&:PE,<YVNbPNTP;dXdA.W+
6^D[WKFVd#cRL&8SZX2acU8[;d7-<J@Y-0D_]#J1cIFUbfVX?F8b25JX\F4d6C^A
OSbg2)Za0bQLK@)[BX1;_FRDEL9_YJJU:f0V36X7\FBODL,-;RQ@a@U-X#@Q:OQd
@#@_:91L>#)#3UO[P:cTGV<RHJGaN3/2>)Gc1&eN4M=c^aMIK^4,O7MbW=+S6f/I
d0_-+2DD3<F/J6Me(_E8TfIYZI,1P&^32VbVA?]@9[M1^Kf]9-YL.Tg,@:dX_@__
15#2V^RG+IIb^YRggB(E4c@FTH=Z;)D3\99e<L;SW2(4J\R/LR^Ie1G+M.+7M1d;
\=G@CX4T>AUQ&6e,\JQa\L]ddY]J:#=)_FN@)AK1/Sfg&]9U1XL<1RQe4f?0gd4?
>AQEd38eUBMSE\Dg/4T<FXU0.)>69>A=UL(aDG7g5IN\T^-9eV(EA\]-UPD6O6/e
\8b=W4H.:R3ER>0F:A8/IXAB#PC9H47D=.dH,RgTUMM0aMe[<,W6WEDCEDWR@R^C
dCe,b3QTG80BW&UP.L(\38S#CZ#,O3H;#+<,YgTN]aLe/gHB;ZUaUF3;Pa<)+2TK
6S1#GdD\e-6cXLVHY[MUTd#E]8+]gO&dSb+8f@14E(8ZUQ5N1^E]&O@c:+3;]0]M
9=P<a#@I537K)@I@?_OPd92e-Ib/I@=f?)cLRC[^E1S/HG<<Lb\<<[X8K;<BETZ8
=U+c)M2\LH7+gWafgQ:+O2#IXMc7Y<:HHN(,3a@LdYIB/,QR\+02GFXZQ084IT4T
GP=aJg[_5-WaVC>SD?RATYEM7SJc&+(fHa#-A)<.\9N=JL@6@MbQ[N1,QfJ=4UH)
W++16@GQdIXM2A@_IG56YXJHV&53bKb5Ba[R=6e#;HLC+gKg5-M?/=H/H0>\D>MT
-N@31#SM)QJULTYLa(6g4#;3+TFXfK9\GN7c<CDN),D)J@g-,WVbC9.;QY52?^50
L:#?A4.],1\-ZcK^J][@?[@MFHU@CM/MgYbd+c1^KV-L429FOMPIcLJV#=Q.0/[<
)8Y(?:\;AaP1K:(L&T7XL#7)DWVf@=+7((V_HVdd21be>GJd&F0KAf6ZO,S86c6e
@DQR^D]L8JT9/f&ZacKQPVH<J9F8K-XF;b#G,EWb\_/XS:FO2;d/;7a.U\F+CG@-
>>1Lb_.4YW./8_,US],[RFJ,8R2)+V/cH]3?22)+4\VKbRT>B/Z1[_CZ#cRC\G0^
U@C9a[P/@1J_KCdTeI44;af=\6JP8^?S=IYVQ)_6,L>B9fLK3-X6E1-(#&O8-TAF
XgP4D0@0]?WL(IU-8@S\65J&S=:b_)f(OTQd3)He58(c2^C6&NCBNIE84.24CR),
&/N?:dbX(M^T>Z/gOgCQS.E8ga?FTfgdX9FB2LUO2G([LSc47/@W::-W(559WdM0
MRRG=Z[AFDfJ<&G3=(8+d)(#CIe+6K^ES\/=[C(A&KUc<WOIAgE[d=)713aOSM7.
FSD1I9AWFI5Nb.aD1Le3B&SUW)XgGTe43K[R0-4KJ=N/ROJ@30YL1J@<?=,U7^7K
_L_/bLTP,VWD=\QU-+_aOfJ<XI)RV4R:g/ff.bdQ7e668=>0WRXNaf31NJ<V^5C4
S8+I63V_CKVXZYTFI^KaAS[&dIWAI34_I[3)>B5)Qb+8W;@NANaTMFeK_+>;;=+I
N.J6&(Z\@&\S-=NPWEKNRTbG/^:W533\03>\:fGKKFF:_:D;WdA8G.W)I)LHWK80
-P=4]17e)\YMT#fHOV1\AaVXBDVc4=7O<G]PF0U<BEFSgR?V+F/;DZY,N??aWWC[
E8=eI;1=_NK<W^WQVHZ].[=#c\W:I&PRQ[7L9(/BURga@:K;\F6,9.#G+]D?K,:&
aa8d;PPQ<[+LWYCfgSM75c^^ZDL=.]ZOdZKA/Z>GEJR5<U<fLO0?V77e?BUT:SNZ
+(T18Q?cE()bMJ15I.TK:31M1Md2ebYd&K^XB=OeKdF:92:<>ea#IdVLF)Iaf37;
9CXC@\9AIJC.Gf#CX9832@:?2;NHYe2?U\KD?C=U,\ZGPM/R9(7dU3J@b:<5a5Y1
F#(;GH?-[Lc0]+EbH4[Z>PLaPF8JFM9/;E;0?O4N8GOe@b:G+6=2]Xd&O#2ZBHEN
:FVf(SZ<c-SZ+N_b5d/_T^FLHB&2,-@I=g6cWC6;L=+[S^C>^7AT68>UY(9CIA8>
fX-AVS,A@_UN@O/?D4HGYd(c&cYbZ1R1/=I9]XD&[YIV=6X^CBR02G=3,,>AC8,f
#3)@Nb_X)TPO4:0e=K;Cf<1NIOC;VK,1--1+P+GC=NC4NH@DHcFRf#R.(V<M3(Tb
daC]LV=cP@gOCU11YWQZ&=1N0(0(.82C<T&bAZ=R2\fO=bW<Z]]XDQ_-V#_Ya#g0
2+PBNS1FB3)L+D-I4Jf6B(+73T0QXD&S=9<E8d2,bOLX48,R/YKBBAB1S\42.E@3
P&?ST^S@SY\?)29I43)AQ/6O2T_BI)0(S4R>3C2Pb&0#QaW#FCPT0fGc:6#OD,V(
KXd/:J8OeS\3G3@DN]b.bN&S?4_++d9]P;L\X)<V0B#_-ZM?0Oe(W>I.HNGGKU12
UV(VcPcKK)bHX#@)65H4YEc[IM@5JC(;J88@;NR,8(W/YMZYD)M;_HUMa??EY((.
+#(_-G6@S+fZJ7/_Kf]]M-YeJ=5^AXNgG<3S[YW57SBF;7(GLEdYDfB;ZBX^ZKZG
6[ML>LNMPQ.bFQ3JOfQ)([LJVFT.4K^:M+G[1\>(dfLf>1B;DCGTdP^3e(Z;aNWd
C@>/G#?P0OX78We8M3W-X:_^4+7@2G?Mf8EI1F44A=?OaL86J4[CY\dVc(5/Z9,W
I#E&M-:UX69>/T4\fN=F8\K-F#-IVBT-L,AUB;253L/WSXS]KN=3?gP7DEeR/)MD
g?)+=d2E=.T:YG.O.#FHQ>]?#b1KSNNcGJX]WQ^BZU^XSe#KSgZ>YJ^)(M9]YG=L
@T)d3>(RQG#5CU0LR^)K<B1V39B1:G]feGTKQa1&G(1NLb9LYfcER>)2[\P/;D^Y
1#Q:\4ec;:gQP)Z7+K<d?ZVHB4[5>,UZGWDTHI]GO>9BK=5Q;.23KcMK,:;XO4<H
H(5(Hc1R4c[7YCU#\Dg^)?JY4S<ObK8c/2IL7(RZOKe6IYT#]A&#ATde^##LA></
EHKLc\B&4>Gg(e,2eM.X?@+GFL>4:5cbaPHQBU)1]a6SBJbN9O4<dO\S/Y5GUc/9
)@?_Pa-F[53OdVDB=E9\\07^g=@M;a:H8CgR8[MbW,H/:0XQ+/WEL.6TXH@_Y+&@
W>Y3<\aT6M=VKRIS&SV-TN<5fg[RDP2?ND_8F=]N5L)&^aWW\RT\&OC;<D)VN6H1
]DX:@4XOf45M1+QdZI=Z,0gY;V@MFIW.&>?ZB?(RW:\W^7bg8QJ;W,-<.OYUOUa(
SIF4UIg-N/A=e+IYA#87c?&_.\5=FK<a_f6Vg1CS\d1U[gGAS7]7+\KK@45.TNGX
A_N/QZZ@<cJV:<>J/cfUG(fIFHe&fc(6b\WWI=Z&<[9#@QT7.B-MV(A_d7OCWA+)
c0HW;^gJ/FOTJ>)^JfS/fO/U&-^_\<;P)+KU<S^cJAC82_0HL92C/F9WAfHfIXQO
e=(]2c87E6O<.e=PE9.;Edeg4T]PZ]V)(,,9FP3.agcP];RcG1fML8/&^5#TgUO[
&FI=A0JO+O)QMOFZ;LQ+[0I(>N?dUf)TG_X(]AfFE)D+AP_#M@B9.7#KcAP:0.BD
<ITMb0)b=U,;/XL0O3a0KXZ-Xf+NQ=Ra_Y<AYdV98BGR9@_]YCg;&QS8&WP[.TBe
eA)W/e:?/YaGgYK>g<.T[)Sdf_]).8)EgG;^G+M#W4C\fBI,gVEE7E_f2Nb>^1f(
XR[3bC2W+E03DN;P]=7=#KY<Q9>3QIZ/=Z@P-g4cb=g2^KH=)4@K9H_H.=gc&Ac=
_>@[BN:PdbcKD0,4/bg]-HO)DS1:1^df]Y5QcW7PGeP;Nd_WI)-08DU4CQ39IR6;
8\LEQ,7Ac.1ZS=K,4++7@1B6/A;QF,a;QZ\SJSdTFKPcW.1<bcM]/3,gO7ca;PYF
0JZX#7>PU)/).I+6cNQ/]dBbe[#RB;6\L_ZAK=2Q8GI;ecG4VV.VY?7cf+gNU5-3
V=U6X\;28C.g92eR8V<8PTc+D>gKN52S6S);d<ZF49[bYFfG?JSc8g@R@.72(I&6
JJF)OROU8PZ:a\aL(1=Y)#6YaeK;1KAeXX]Gcd?>/aS>[FQ=VZg4WH(_(,#.NPO#
>&9eVQPP7=L-61<82N<(6UeM\10OWeHPS?DKWc,cLW)R(He]66f/F3E_XVcRGAg5
F@V23:UeAa^f+E\:J3.9eP=I+ZKc?cIeK7DVcSON-[gXS[\;L_LOX0^F2@5=?L\f
L#Y:aE[c/(IE7Je87gN4LF+J/Qb?9ZPgC.+2,D1=Y]^gdg@NV7++:I;,B<JQF>09
a-(VP5@2PXR];I6HG\RJ?;Fg7YD)-><RUBYS0<7YVMb+O3[H,eBdT:If\NOE[EC/
0C&1VcX&L^<V8eSbY3T1eVXYeLM_)5-L;7[aJ2#K<]2e)\9X_1VAC[3CY<bC?Z<:
4U:EQ3gfZ3daI&92f.<#aI&7MLb?)TGLM&eJJ[V)):]+)<R^g^MD;aYB&003M^:a
U]O<@MA/<5^,WbQ]V7EeJB//>a+X-J9BU8=B:Y_Fg:)4cV)=]DefJ1U:\/dTE=Qc
=SdDTf&LTUM?6Wf,F>-H]JB5]feG07Ab>E)R_8ggC8e)MY1R8[LHgH(J\[><&#ba
9GgfU?=GKT]RF-EDJ854&Pd\#]1e94a=d(dDg=B]5JWP/74VG4)Xb9fFPYVTbNLB
=4bEeeL?,4Gd.VEQ_b_<)18gNg)O]b\Q.X],H8a7A#9W)4;e2L3??#VScJfV(KAe
-QITNLF(6-<<E2aEb^]63(;[C^a,9:MU2-MGM[GA59FD2&<agU;J>,Q1>VK4Z(+V
Y]6B-)93)21g16b+4:YPJ>.)EK=Z\.[M_=1=;L95Cd9=LRA[L,_)Xb,>E[eLPHZI
M/SDb+9ZT=bK(R7g7P7J:PM7f5I>^BS,f;I@f5X+UOdL(=VcB9\L6T(N:-?U)S73
VbTLB;PTB3/K@?#bf:4:@?CMI:O]U&N)_?SHc68E:U74e<b,AX),@=7^I&VSST##
;<:dF<8U1&d(JV<_6A+22_)[I12)0]KZF#e.c,AA6A6-U5b+a\/<ga>[2V[ZS<2>
K7eN&g^Q5E\2I(1U@U(1,\=+JL8O7V@2466;K@^TJA8NBC,,0Y#M+b(Y#0+03aU\
,^]OE[8)0?cDB:g8H:DLeH(a-L6]LJ6UZc[\)d6@DKB&X85bI[PJeF_9-G19M032
=C-.((>;C&/^/ca]),@eA?8bUaN.gTb^A]Lc54Gg.fV=<<Y]^LYYG9a\U[<1=69A
W6BM2<L=ee4+J@[I;[A[[GF9e00[(bN0DTNO?E0>TN0b#P3fecT5V:\;C1+]d0[N
5\4SVLWB56eC+3)1UP-4EP,1EKW#+bUg<E-21237T6JaCZR0U0(dLU+HH^EUPJQ9
P]G(>:FCe+KAZZLS8C#(/_;MF[\^^C2J_^6J&ENV<-CPTN@RP??TMAbIWaPX]C#_
\+9e0:&7\Ba>a=bJTa[J\Z7@ce]RV#UdK4Gf6>([Q7#dY5Vag9SLQ?CLV/Qd9BI_
;XAYG<Ta,WBDZTS1\^<.-9?CAK60caHd29cY]<Ng9Zeec)0bW:ZgD>RVO#P2gOa_
Z>Y=NZHF<ceAg391#JZ;8DZ:1?a#fZN?[GB:#f#1W71VB:IK+LGO.J[b^BbgT+NJ
BQ>b_:/2)P0,<YRW\R:UaTKDEA/7N;f.-d+Y0N_X+MT_M#[LNZbfgAe@D/2A_=T-
566:9@+)#J.FVa,1;geSAg>N=bFNf=7Qf[Z#I13K(&7/&X#)L\9<NL1MQE+\?]]D
.+fLYEPE>cF?OGZ[D0_Ee:@c5\B-)^,TKF@@]1b^fLHYf0C1;?AU+a@ONDLK,DN:
A8&H;8QI:)#\[@=M1TISDAb<fd,#e+@f]Df<I?b[NU@JP7.K-a/HaS=IBSVZD7(T
NGB-OaFEWSHT^P\&GYfSDZ]YLNV;PEBK++L/RV8L8=.;4FK\\S7[JZSbaU9J[N40
V^g1(OI;B\ZQf\#f]U18LPfbB;L#>:@c7WQSZ+J8K-=N:RZAD]>+=JY(FfR&LRW6
,Q_+T8#-)d[FSYO@3L&Wg9BP2>0HU0SbYa/1D?+8XX&P[6O.5W7)bUe&DA1;g9-g
C2RB[W[cFe?TX@WO4W\FCA,e5T;BH_+IWbQ-YO#/_AAPEfZaC,I]LWb58D/S)W>?
2KC&,RBEXBI:3FP0QK\(5-G5P?6+^(/IX(R>39VXA04bJ235Ud2(FOBR6&=A)5_.
IR)3>N5dI)]+1-GT@cZe58AReMFSNOB8H_\V/CR0e@HG#Y5M-+25bE4ef3UaY\)2
8A:L94RIOTcH55&a<5DSUcf.MF&_+(+MLU9V;<&[cBIC&ZaYWVUeF>WG#A/<SdDf
GM2,132009W)GfI)>3PEN6@\&H\//NJeWK@)-RDFRG<[Meg5-I+R\Xa5dK.BMc==
WPZT<\eIaQf+ZeF&F:Lc(VL<6>JX8bgI-PCV:ZSR=6Cc]V.MgWMA&=4E?7aY/d+>
.1/_3g5LWFcLYbUP?.]DbOC^OY=KMC<<Y>PLccI1JCY1eFP77TO9GZ7Z,:c(MC(,
[B&-NHQ)c/91--<SWVc>5dN>N@Zd,7S8(J-NSK>&R-RSfIV=3F4E_L3IZKOY9C@=
(RfEQgI&SPT]Md]g7V3c=bUI?:4LG8.4?cLVg0SGV[\:#(X^cFQ+TTEUZ=Y\DBMT
O>-(Fe^#d9.A4:Fa]N24DAZ\c3U)aXbC^e+E>RAaeT[,\_fEE5S.G]_&GQ7Lab91
V<2^Qg:I^VS1#.AEVOa@+CcL,D9+IKRG\O2bJ_RVT6KBXUa(bWKR@3R4R<F[_WY;
a]D#AedGU10JN=067IU;a=:M^cL.I==4K]>WW[P#g+&V3-U^M:XQE&(F3_.FEZW.
#=]2W/g7c5[<\[J_SP,/e.IR+B7Q7TN.28DHZE<1I?f/LNP0#3IZXZ?],Te,148E
0T+I95L;Y?dRfOWZ4K7_8K<K@;AC/;aQH/G6^-?Q9=9SE;b:e>BE6[)e1,&BU-=A
3Y,T/gb7OcGgg5HR>aP)WW@QbKZB&[bg5JH9=X#E]L:4(=Sgc6T/N70OJ.4@\_KY
+Q6)V(EcAN_Y>W6<QOa#4S9,D1D2?&CEO-?Y<C=>N6]RAKHI_L^c23E?@_5#WfF1
TOaIQ(a9L5eX@f/TMP1Z@U18:/f6GSNC2W@.;g3VA7e3/#D:14^a/]]600a)Y6SB
ORgZV#\OWYbVDMgQM&&#,<WFQX&c7dFQT#55M2_+e3=@/-Q]B<BBRdV.PN1O]V&f
KcM]d>&-Y1P>61]0b7LaM+fC9BK_6V\.67XACGc(6C4[/g=]eX@8X>5?4CQV+;V6
<9^4CQXD4^5JI8bA&)aV@g.3YO[/0S_6=I_VV,-&?G>U^,0L/b]L^Z94[/9/H-VU
GaeCde1X6V&Q2eIdQK/;#D3_4]2&,AF)_CQ^D]._(T)^#]F-A+aL1]+IF^7[=+Of
&DfAQeIH>;CP<a-2RL\))OI+-5+.R@1U_.4g\bfPO:5;]Q1A\_ME,^PCg]U=(4(I
1>R1RZ1VEc\#LY[Yc:cDc^](GALK4Hf57EZCYK@=XV;[H_DcH?<.>=7@d_O99,OV
OZ?0.#BU<8M/9>F1aa##6gV0FO>V<\3038.#1R9,.AXfTV#Q#M-:;9J9fDYWgV7f
WM,1g_ZEZ(e>4D0[W00E,<ZS\O3DKI+LK(0fN,ZB\DDeO8\NM<RSATfb_IC&\3>0
LKJ2;AO&PKPHY<3?/,LB[:>?f[A9W_Rg1MA/b):]LA8BYY2=bA3+V=[YAB8YDfcN
d15PZH/M[caEUXJKTJ3b_P343H_L@XGM)@Q7^aTX8WeN)S>#HARSEY2XI8P=+TP8
3DE>a-@/_F@5c3WD&JEBR\I_Bgg9[@[W&V1-Gd^HX+X,@gd<PbO_M,YB+Ce8[P6)
@S2QeNb;9D8>f#ICdaf<<L:<,+@KJMD;GQ\Y17VOTB4U>>./>CNJS5_D7&d8+F@P
P6V,Na+3#LY-HT#OEd3BRafgXMF,aF03+,b0]#?=[H73Oa)[5=]O)+JeMWg0_YY^
&>V,UBH4UPNe(44.;8Eb^M-f/F;bX(?Z\2HP;\I8g=MJ,=,5QO=BgV-^A\>V/YV\
I-/HeEA<#X=41eZ@H^7NG>CH<2e^?0f\<H]B;D;cSND<][EK#N<.e]QaJ^gVP4Z=
:dNO(]9<UggZ8V:IZeD+8=>HT8&3?JE69;RN=U_-G^T]6.<g>gGVc-7Y?gFDI?f)
-5g?/:8QbN4H/9ZY^TDQ,^H\b?cXF6YSHQ+/=LVIKRX]_&5=cf-1c+QPLF2,K#T8
EeB;K2_>=6[>5/=cbGBQYSMXU.eC<-#YJN-2HJc>1#F_-84E/SIdFZ\cfL:>Bf+C
bT,61,=PK&O6CQ(3EMUX<H/1]PTQ15-CTb6^:@H@I/\B[XK4A/6Q>)U@cJ[^\;Df
B0f375FceW#A2DMFPXa[CcJ,^-3Sf.8@]<6f;LIJWM?5(IZ1dGO7_D]/?=?Y:K_A
GO<6LREC2+N(#1c/OCJ_[R+4BL;RC7U5<9.5eWK95-F_1(N-ZFa+FRY_GQ+VS.b5
7FKYfaUUb8:Qee^R>4&_N7e^SS#M-(K0-)6Xca0PWR6L-cg9a;J>&P7/-RNIdKA^
feAJ8g,D0bORZcPHX(5(b6[(W--\A4#DQ]:.c_a[2M\De76)]K99G&R=0d[9+A+G
JZ]XG8;A2Y1f\M^,67AK(c5Y,=-X@;WZ7d=_;H6(DSJ5MLLR-]NMKR_1d.-UJI^E
[9bceC3>VJD2R,eaE3W[LQ7QUcUZ;++:1:(9O1QJ^5B[OT<.Q2#@ON28Y]OYSM?K
:_fE4PNXE15b]La\6ec=I?3Z(SUI[.@1RT;g2A9,Pe11e#@),cWc8:1.QU=?H:](
BRRWaNG8f59]IYOH7H/4N0FRP.X:R(LN4MO)MI/U#O#Qdc2b(8]MNN9YQ=)g7VY9
[7N_.M,6Z6O7QX4))DgBF^U(2;)3RgS_M3+(UAIBEYO/_J\YR01a?WN9&?I8]_N/
7f2#<VXX@:3J-36-/YZ6F+_g(?+N2#e]Z--[X4e,f5e32B)WCP8&=]EBJ8I:8Cb1
[-OC(9,A?>fLMaZT,LF1cM9W(+TL\\g0.@AM;cVce>^N66be3MUW(,<3;#JLa[(0
eV:/XL;B_F6==b50MG+a7+.A2:d-=/.S6DI.9<(9dg<cE,,&B\:I,M2Bgf&35Rb6
3N#3Z191L<0g0\g:W.f81-S)(5GI0Q-(Ge=/Ze@E@VYJ8;LAW&M;L\gSMDcXH?g?
D4D78_LeD.E9.\MWSS=Fb.-,bacOE2a^0].cg5?C-[@D#)]MXdR8_MFLO3eb10)@
=f,_A_.<f<RW7T3WGR-&X)&@H9[[cAGgBD<,?b>c?<J^#d)?=JVgbYS,5/8W#[c9
1-d7:TLWMJ\/7(WdDS]ILWXQV:d3cFC+2PC&M0^GNU?Le&e_,FaUQDP9#91:JE(S
N6Zg/@<g2OA&[-6A>73:,dc==dg.Vg]1K7]FGe>ED/6FQJCS(8#>B6Vf+PU,1Ya/
fN;cGLPB>&C8G_LTF;-\[_//Y=X&?cNa?GFE6I(F6O1..O/]/,.(73bCIS(2>_GE
(N+VLT.d+B?[f#6A=[?RgT/].ZG9f_6UPL\R5&I5@<0D@bfc19]^@d>US2OG,=:S
7IIfQL3-TW7@XMWI?5Q,+B\(J@?C2)RDEKc[YY(gN#WB8&JJ.,-_=VV/3>T?IXO7
1DA#Fcbd48G?RbF/a#f,E1;8W21Pb=#^N0dE,I^,1GZ^fDGZP7<>8T-ELCJLWZWC
D/N<O28eXF9d9QQ:\/)]TI^c_cWc&FEV[4O4>=/M1S_1d5_/ZQTg(YPA9f2BGQ@=
OBN+(d8<bN<4X<->0R7YK;a+aCG,THP<4OYW9\>RM&)GA<aS+JOV,D+,7K+?6Ze)
=NaQMJ@Gb,SF.g52eY(&(I8@e5IgWfJaTg7BT8cG.KZ4eDX#[-RNS_(EN@54Y1eS
ReDN#f0c6f7>.AL9L)@c3W9:+P:B^D\dJ\8+P@+]SLS-XYfS/T2cDSXG,b@W<LZ[
^_7+3f6g]X/1d3+4Z_W,f-M4CZf,P[_1X#Ra.]#YSX@\DW>I)c;_AJBf\5>Y1[e^
#;B/RR?XH-a/^#\F0&d;1GNbSVD3A?&]0SQ5>ML?#A.eW00FT2Jeb8(c08LT<fT+
gTb#1T((@8g&1[W^.<^0@02P[G::J.M0_cbgX:TB?g/6,6Aa:Q4<fE[;c/D<F>Wa
AQ=O>OE3.BYV3K]5F/N9Z:_aPD3Ie8CS[=:+&2CV<<4DC\/H_X5+J46,[>MY13\+
B@d4QU<d5]__N6RD)TIXQK4RV?eb0#+UPX;DE+(-dF,+\.C-ba,TZ;KPZ^GL[M(K
81.=gW;(<+VcLf0^d(TE7K-TBT:#+S0BB,3KUQN84A3&H+d64FaBWU=c@BJ51De-
+&A?[J>(T5O?]P2V,^0T/6KUU-B99[P#7^^4[E[@L,PcO;K\5P)b3M:IB5#1#M2H
_:+J6)0)fMEd3&=)A)99B(+9CMD102A+-a^Q^ZBPXV3LB6Sf8<agUO\]\OX\#4]N
C&,7FCa;_1L04[V3GC[1&9Nc/,0f_eA2P=^/bgO<H)C?+PM;7_+>(05=OF_OX/88
;]XQP8QgbNJ]g0.PL(/RIHR6KYN5c\3/@Q-M5L\1EP24M9EO/C7e1f_T^1J.6]:=
CRRFI3+a@<HDe\D+1Y@3VI)1b;MbK[&[BYVU0>ATD1CN;[&-dP&>](/ME#P8#?fV
McQ9AF^5f>dG]_B,4Z74&DIaFM>-H8.HZ3Z7Ka)9I:K87U-6&#4fe9OT]Y^L>#41
W4\H[,I6RcMR\7&cJSQLSERHa#YBOJ[.RXd8ZHCTN^K3Nf_K6LPU\CKcLb&0:1D/
ML=\Q1+V-)OFg&EL#Bc^Qga#d9Z8(d;.a]3(Z:H>cdXCHCMG7E1)EVQW;bB]B7U<
a5Y)WbaJLQB[\Ee._aALPO;B@#7[HbAa/)_,dN[<8CE]B>LEU4Ea#Q]I).5[PQ8(
A/MD-,)<0:Wc6IRTbBM=N1EBM^b_JdCM&#L@3U/;1(;SBKeeUMIAGS&JX?KBS6b?
MP_14+1^bG;<6?O6b\1?8C=\M,\XLcJ)2d=]8Kb@-eU5#8+?OaW#:,#g\GY_U\?Y
1CK5-a4>,]@6)H3:J\dSZZ:C1-46+D^^+4&WM2R:W5<40:,[&eL(c9?a\-S>OPgK
5--dgKQe;8?,GY^O&#XKZFE?5DRZA.VL.-;Fa2\KdfDOf^.ca24OC)LcLG_:BfI3
V@N?HfbJeT]FXF+EI:)Da>_V^Z11-cdgN3->M3?+C+^95R?B-@6<:40e6gJ(/WT(
GTPS3e0+CC2:6IQO[-PJWKa)e(fRN@O0X?_M-gO_aK/3FA9531c6#TT]IIWWUD\f
,98<g=](J7C@JW(9<YDC@X3SK[^c<1DCg:&3UcHP/?Lf7A:c[,[#0MQX&fdM6fdD
\R>RCRNdaMO]13H-N;EE(V6YT[MG>gT7c<@?[+NKT:,9L:8N-T<=TCdYF\N+RITG
e&BdDWS:#J3Q++I=eZ@)P3:Yf<^e<M3Q39A=GRK6AU7PBZ,9B,<H?LZNIWZYC[Ve
9Z&a_U&.^EZ#TPN/9#E^A0SJ\;E=5WG,3T;5H5:\#HP9J^+e5ZZ55A^>-KI@f5e6
]LP.(3GLWCO9.?3#,;M2MQU1X4bd)X^;C?_5_E(-Va?bM84CVN-4>>HE@/8eRI4;
Qb1WL.X2=)PTIRS=T^OH^#>_U^B@NL<XbIW<N)bQeY4eXceQY8T:U8d)74_a_@Jf
XD)Z&daRU+-<0-Je]YXFeI7WBf3]/E2?=BI+TbXA_,Z#[;JQ3JA0545Ga4E7@2_/
_R-?WTZ2FE,](0K]b3_+c7FZTJSO(e>,A^LEDGJT4N#GHcJEZ@<g+HgAa(BX?4OR
H9:f/XeY7^PN.(Q;P#(J-T_T>FVG?G3@^8_07UF-aZa9-eCF&C=+cFHEb&C?4CH/
d(N;D8<HQB7>>NK7L8NFX)#-gEAT(T3BXdJ;O6#)YV]?Ob,L7D.]^)]QB:;cG^XW
SSRb[7P+[SQ@;([dEg&0=2&6S#G)XfP?b1,0:3Q51]\,cOBeJ\_-<7]X-a>=MHDN
WUQ5,?=HTLgSeKKR1^:fK&J;:XTCJ[U)f9RJ_Gc8>X]f)QS@,f187>gE&gVPe.94
J[aJ<N/7cA#)^0Bag@Xdd-_S,VQ>FG=8:GSPHg+,S;A^?W>6<QB-H1cHPeA3E,gF
bQf8[_F7TGT766?+HeeGZ]\&1MB/.1gC.d2:1+,a2]d:475=-KAHL+EdR/.8;7[#
Q)^=KUca89R[<=(\3]^TDY,a&]cY;UGPO((5?e9Y^bHR)CND:PWF<H-@&2O>RSO#
;UH@,2U^<c]=X0WF1FYYf8aeJJ#8RVg>H<^VWFAcGK85+Q+BDY@@1eL<bHOIcg+E
SLC<[\[3&V&<V<VP[\EA2PF4E_IZ7cI;/KaIKK4\6>2-5Q<0U1A>e8f/P4:S@L+>
bJWG8CP\Pg25/)gPfEVRaeVXP&1Oe>gd;;O_5=#D)/fgJ6_@ZXO6ad;b&F1[@L,W
_Ac,ZaT)FgN?gaR114fB\DP+B@g0FEKbA>fc8<2fI3gQ@T&E:J2F2c9QZ-T&7b7[
[Q2cBXS0FX9E26]=MEGTC,[^bfdb_OML+I=#d7MHLZ\:)FV&&PF:/^P88^34B>Mf
U2S&NK^1OP=C\0#e_M:JK-MH]RO&e<Ca<VA]-DT6A9Gdb8^4-T0H,)R\;CCX^QSZ
/W/W<[IS61)Pg;fZa7Q]a;g0g)3K@HGc3WM.EQ^LR)@>8(2KY&C7#9g5O&.EH&fb
(ABP0Neb8L5-V://)N]8XWGD8T>&TV\R+Wd50U.b@&0gN4(8FTf@[HO[b[ED3#d4
g[K@?/6FX.e?Q-SZ6_@4)c/KHGBMO)W(]YLH@I7a3e4PK7D1X\Q:>WDXC10;B]Of
Sf_&B0Z?YagZ@/B0K.\3F75@CQW/,/CGRd^-F@)]B.VA86GPJc8VEd)X6&fI;f?L
B6N++A8()Y(ZMRUR2?d#K.40eY;aMXQ^KRN#(W;_9G5DHPV_HO[1BODESd)JH&R]
2V4<1GQa=4+OQ+.PX[a>DJeZI&[8&-/C.?L1:W43#Z7G0Y3^C92e...>H_:[JE(E
W5Q9U7+b>X<M>P_1)(]KdY,LK0=&HGK1AL>K8A.MRR:e=I2/;OF7FR1G^@/fM_0#
+dA)F_X>?[)VfHNC(6eS/^>>Y,Q#3L:N[0O]FY6>&=87Y:=>KOL2,CS5.CT(J4c&
4>RV_30I,2g^U>12N0YJM;RggPZX6\Y@dGW=^g(@9T+-E8VEX#<be=e;dHX/U6W?
X(,6)Oce;[QO5;H)AL.9=99SOR/KVL/MVRcYZ>V.#Y2aTJI6^-4]N&0Pe9Z_EI)J
;^2+fT/V4:)_RU1T<]/7_5/]->U]_&gV55VS#XXUIG[]D&N=_(R.aJC86)GVG9>e
XdE=g([?ICA?&,<F3/S@a\_SCOUVJ3^N]f1e\5(@8&0&fBOK&:D_;/_cJ:0,(.G7
RU?CU+M_N6NbGDg,7-T22?+)2B1SBGb)4dZCYQCQ?;);aZCG?U^K_MKQ;L7K8RCa
8>/QUB[:N3C<-P9<CC;;<VS>ID@QYBD9FSfe1PE]DI[4;-TgX7,cIE0>YGA1U\L^
JM.:_V9>.?QE=+FUaaQ-:^d8dQ=IAdB7M7N],#J8T(A>;B;7P_e]WSQH7#VCXE3S
KAb..QRHN+&-DSJIFLaJSLf<45;E/d4F>>;8JPG3=+,aIMF[J:DG.?Z.DaAOY&G[
dXYPX1^6Y6ETC8Qb?67f/PcdPL#a\:4-)dKFVTc5A/;6^dgegP)_F3Q3=/<^CNR,
d?5YM.CL(3:J@4PGZ9_\:dZeYA7e6,(I=RIGF7/M[d@W:XfO8-NG[4Gc1c8WYSJW
]>H2E\Ub?A0e.6aVR&X(MTIcg=D=<YFI?cGe,[]X4X&9@L3bL\gW>(JJFbQ=CCT6
4BR#,/3^f;+0F]57,]7NH6?ed>@KYdQ_4bA#F58=O..V&c[6e/BZ2dS50E\@Q#58
H)><[>B/\A-LPA.5&@I\RU>Z+Z9C(;SbBYI,@(-;@((R5NUeXLC]\&9]A;2-STc9
3TLW-?2?:TbH8ILEG?47.2.N#&F[^HVSA-N;G3J()g1;UAc5Q21FM77>VXd)BOUQ
HD;eYee@^6cMK2,FOfL>U2Sf?U_4:L5PG05F=]#8BbMRKeI495IOE3IcNMR,=403
A1O5Ue_3<KNF3@3B-cHa]3<6;bPaTL^KAcQ=U993,a3eM#P(Z66E<2g\COLN<EFN
g4cLP0DeK#15\b?J\Q@_-S34ZL/@a#3T^YabYPaZOSM3c2fC),&;:[\#bZRZ8RCa
b91F,2Wa^5?Y@_N?9f-PcTD:Tbb]_8?0dCEga-BLA\VSGgZ+1>ZZ)eM5H)1U892c
F_U8BgV3^];]?:J[Yf1;3@_Ce?0b,cdJ]a8NW62cJEd873ML9?Z)c_YWbe/HFQKA
(Z#fXdT7WQQR&)I[\(P#Y=0UQDdW>dV0VR-?JdM4c?HBg2PP.e?PgND]:@cD8fX9
01WW5)7>0dR<eYPX\BK,??.6REGAFMbE+^CWL/GETfXbg)D(d1Ibaa_Sg0b3VETQ
)@b5D3;ST@J7PUC,9>1/JR/A:Zd>:H=?f>T35=)+=?8e_K,Gc&f?87eETV)5Qa?W
8a#C;eYRP[RE)FAU]0GGWaJNT9JZSRM&D_I?4=a1RR=7c6INbf5?A:8F=c;>c8]X
QGO[ZQMIeIH=?@P#?=RCGdB=g.>,;aaP0>V#7FePO2;[c5+QD17V(a8F@a\6;gX?
H1,R5W;<L,fQMZ)&\++C6]Z(\?3eBZTCV,I6)_[J/XN^2=>PKaVaOLQe-&dRL\DQ
7L[VG0JJ(_^0[V;0-f7,MLT4(>^P#GA1fLKLbaAQ2FYC[BQ^8DJ7=@:P7&?=a=^.
E2:0&Z01,9UXOU0eR?T:\VY/0PUV3c#5#ZL>A(E[?A>>Fg/Y>f[FI]8KW?O?,4c0
9+6376bP-Xc?E0YQ6+^N_GIU7(I+BI+MF(IGYDLJH49?Yc1#-+4+/g3\8?2C;F3.
[SJ\#E=dH;^>fIY8]6SAOGVB\W=I;EEWD(a,Nd;38E7_/2YdI451]gFb&d#egN?&
R2g,6:E#_]cH0II-bXQP5VQJB/aQ[9LCB7[.GM5QGHgKJ-+FJJg:c9OB5Rg^#Q=2
WI2cDV](<U/-;UC4>_bGS51/-&O8#ccd;R3LFS1EWUV3-JR>5=MD3:Z96U45XcG^
/VGJ4TXKG2,WI1EI?,N6:)];GB/J/?Db]d_D@cJ],3HN/6ZHJ_NLgQdWQ3_LTc-K
)a++F]TOEVWX;RfCO@N@B@[5Oa,aLM0YE\;7(NXg.1E7(:L_/&_NZH4HJXaJ8>cQ
ZUN^I_VVQ@?:A__);&OQZNSS=G3M3]b85bC39YRF;8JH\a4/FDKD;7PN7]=NI2?,
HR5OM(9cS)8=V3&L^4U3BU3O[-cZQa4J4Z96[N-1\4S,eT_ZVOAKTYfU-C-]TE1E
=A4)a;B#bL?KP,QS=3WKbA20X9g^/?0T^(^EFW)D(WeZAU8]5@#-a@cUggVY45[D
+Wb_?]bLAdXSUB\BASF-WMbJSY=&)c)56?5OSFeGRDPE&NIgXYVMNY:^^ROVUUd6
GX+c=;P\R#AT?7cE>+K,J:25;9.;+5+:aeJVb=K4&+Y=U0(b(N3-DGD-D_6C@&DC
:R][\R-/=eVeXRHF5Y8UK7EMH;?GULF12H(21JEfA0E7.J9XTU)V;a9,IG/HYIgF
XP1D-XAQfCg3(c?,PSTG)Nf9<[9eOHSFSX#^70,:b1^^F/UP.KGRXM4JBWLMbH>/
S:EJIF?L58#]Q/TZ19ZSb=AbZNZ?(L3If\SQc=<RJ9NT=N)RJ@3+AV_0cQ3&9XF6
<7BL-b);=c;5>f5RGNU95ZOFAUaC[:baI&>)<E-6-ecYC1FQ\\&A[O+_P#A^E=f[
H>(c5/9gT)Bg&/)-N.NC_d?]I4=\)WUF+Z7&;4gTbeJZKaUa(V=:T7]4AR.3.4WN
IgM<#/S;ZdTI6OWg+0^gR17T<a\>eg#a>ecROOUGaA,&e;AA=YARbNVUb(R9H8^6
S556SWKL-[D7)SIN4M8:/4,J)7I-<G7Y)2^JBHgBUCHJUIX\G\&ZCH&O[SOX[4c^
1f0MATUA_;FFOg..2dAKS<D+a/6]6V[W-X2/bLY@8]\0eUY4(\]],\,T^[D,Lc),
#?>K-e:V9_@4-Q34C1_NNQ+EdV&&BL3b/,aFDR9+Z;T))N0^<YS,?2<LMR_PDOf/
FA<-U^1KI^_4a<HJAf,SO,f#CG64<#0X[g1b=4DKG@3&efL3d@:;5EV/X,GeOD?2
6dTR4(1O(cX:N1H;O(#02/Z+SLT\.JJF;:KVYeUMXeX7#^3LS?#9B^g<;\A5Q#&X
1?S(ZJ,b]FD[P4T;_]U.8MF>Y)Le#QWg[,#FdJ;P3b(6_CaKa>eN\^3KL#S)aRfg
1YPVN4Zc,c3b(@46LcU,Ne[f+67@)<\:DK#S81D_.03&6b<O?f543TCH,MK\]4AU
=^IUGI0P/ZZ(Xg)/Z[JSA,NMQD:ZK2DJIGDG9a4=+U^+<0Z64TE^e)L-GD/M(0G3
T9RLY7KSW&0HM[2S@aM:]&B3Gc+3,[M1.Rb8V4I:W-M\EcQ+FZZ_H8[3].GbbGTV
+X48:@WA]CUZg4JJ\(HS7(2;B\<<Q#NN4BSB19Qcd/E6V=c?#&VOeddO0;67TD?Y
bdT#I.ZWCGCNDeD[S[Lg.&/PU0M3)#RC_Y)8BILU.SRgUK8@aI4A8/I.[QE)0b(K
c,.KNYF&Ac8BeBJ&e8)0CQ>OCYHg\P2KF&R9DZg^NSMUFb+3RM>/299G6\CJPVXJ
9CY-B0C#Z&COcZ7&KI4)\\N<:]Pa;d2a>L(2(d&#]J?a]c@_[.Q(MZ.e;;<:0KC>
&.aPB5a_XA,aMFGU[_&NR+LNJH3Zb;e&BaYMNUG@KH4,?TCf;dXK.fJ?D)INJ^bb
bRC#USALW+Z:YK@+1JG=D\D&:2_Y5KO03SO,C&<GALM]T6b9.I.D9BS:X]8WI#&[
R6W=<TM2;GCNQOeWg&D1O3g28d<g4-1b-I;MF.>+BJO;f9c2\^)T2RE6S6]X]B0f
_Lf)Xc_L0>EV=NYR:f,NJVL&/P+R:=KgM;0YKB^)=NUS9gVE(Y.^LCdg9=M[/D>O
Z4&\5G8Ted;2B>;MD0^69&GC-S:g=Q->7;F.X]S^E4VAV:0B8GP62_H12IN+85X/
HOdS40U.KHBVLbUP]3?QR+7DcDL]^C<QF[+),F]LK&FW?P9GPKOXb)(Q@a;MEcY7
;SeWD,f2<K9/NPCRMD^,eYBIaP#gP5<^_NN]X.?UE7\+G6=bJC/HH9cc#4O_(L?f
Cdf3S@4F5KG<AVALKC/e\CW01X+P]H-Q7(E8bd&GVVTJHJc-8[(,+<:Q54VA95A1
:JZL7N;29H,g0;G4TJeZ7aYM^PaFTd^gD#f=J:6NFY\a.?ZVQ04X[#XPJ.4;NINg
YgI4@INf(LV;XFf+-XP0S3#Uc(OaQO.#LF4HgI/68]JXSe,J(VdcaYK;NZYTIXND
VF<0SF<ORDCCG9KP9Y<-e1Rfb[IeX5PM.B&Q>LN+<53MdW-e?T/E^&<)\&;b5Nc(
@/M.SAEK0Zf8_)DdWVJgZ9B8NT0:?=&g=,Y#O66[Q\Ad^b=TOfA)A;<BPQa,.HAW
-T+6f2RgV^+Y482#R2/7,SKJB:b^9UTT]KBaWVBfEXcR^YE+CP=,IJ]A/EO\J\/a
/RME.)/K[1a.)&Rd<&Q@e=H9_.\?f84ZB.+1\.>OZTL&C03+UW<87,(3?AfN@I&b
WbAGD2\SdTJVbKWCS\1TX=_]LOL=A^&#efDBK<8W3SXaX+J:#GE.<<(:D;^)H,W=
F@@ZL[b<_GWK)Id#<L)H?-G]a.J_X-6:1GEJ+PO?Z_^._Hb;WT0-_BL9^1LZg\B4
=6b_TI,.WdH+],OVSM>[AEQG4-RDJaNY/Ta3R?@IJ]K((CJ0gN:0VT;.)SUY:U-E
c@-^fDU.MS)H(Z2d1VN]P4CWcI785F1]?TUCIZ.76Z)F.AS50(bMcDEM1:Y2[;R[
=14DF+S=WgL:SF3,d-CgT\_LdH,A9/>?,)B)UN9/?16+g0+9-4U1+HU2+,97f>EJ
7MJGBNf()J0WI_@V+5>&5AK^S-9d80g_+gA,KN9<X^;#F.Z)I@:E98TMEd^=Q@7>
=ZNcB)aXGaV/V[JfEcg+=2c,0\=#K@J7eRZ,^:,Ra301?O#L>K=c-H<2Y.PW=&>>
62GcTI.U^CP59>:dW(>,e2B]>U4@Pd9DHS6:(WYdCd/?IT-._[753UBe6<I]18[#
HE#Z783-;HD7)g/Ra4>J2C?41c/1SbCK.PO_.>=^4a/^f_+)9QLMHb1,;7L)#aE2
77RBD1^,&_>\ZW>CAGPBF2KZGSQHbg5AbPGHRUb@:+daJa\QYc3?>+[9U/ZV)BeR
7BWS<UQ6[SH1f1Ne^S)1@779G_bTOH,QT#SMB-H8CX+E8(?9.9GVE<g<\=T3&-OK
OC)(&b#7=cF,c9RS/\d-0eGSdXFTL#cOBZM.HQb^RG1NL2QWJa?E98/-^0+3D@;5
QXc?-QOGH\&J(U]S+a1P;NJGO5\WDRcLXP2c>^)SUW18V(@).1&^0I2A/LJbEDC]
)#.fbQVcP;K^:K+.bH;CeZE<SQ/#Y-M.;g1PDe\7M/Xg53&E+UJ>/f_HJNc78Z&&
I6-/XdOPCXEY-=b:WW4:3dA7]V<EUTgU7ReHX-+&D;2SGLH^]X4NZc_(G^4?0=QX
[/&R075(W^Ee/L8B?[GN>J&IC1D[XI7E5AIVVY;D\US+dT.0G?-AV4[NU2CR.V=&
V^I.9AUCC9P.DVFFFL]=BPA5Q;Fa/5f+@6K7V?H5b@-8OJaI^3dXI]Ud\cPR^7@>
aVgD@C+c\2<46,fHT^G1JOgYb8gO9/#3HBDV;Q[19[^RSB-LSc7A7CccReS6MdS6
VX:<3&^Ob8F[HfGcEa)88KR?5&1\Wf0Y8GYg#7CQU>Be#AC>b@_;(3a@4@:A>;A?
MCYcSAHf[Md##^?fWeQ<WHC+,^DX\BMOfV)N(-Y4MV4I])aX/_F)(#OQ]P+3:?KQ
d>Ff&47/\_?LRSd++RS=PG\g2=gNB,Z1<I[P_/#S_#Y=&^E)=2@@=[?F[dO2e8IC
[H8<SVMK=?RYJ2_.OR^KVTY=(Z3P8JKMSaO<Z>f9+HRaP[0^^XgM/Q/[ZWHcZf0C
c,WGK8SN8f56^+J#,_YD-UV2YQ+M_EfU549BKYO0RWHJW57HATY+FR,VIJ1)+Ze-
MgRFKMgR5O9)^-S2IIJ#[@]7:6MF/9(\L]21:cIU_G97daK5ReaCFf-?:b?c,9C?
U87Q2>UBATKX6He3,+2K^9ST_F+>CG05YdR=U=K=[/[G3e[b2fD;#CV06&P]]:WR
(PZ#U\QKH:]V4GX=[#;[:I]-?,I7VZ5JCaZU688[QI+Q&c,UXeSC>2W0PC3\W+NK
f0#1HO,Q3)f)2F?E)\GC0#-:>2,X4PX>1aGTRTREJ>Q@B4(31+f<b5.=W)8-/HDd
fN/^,[Pg=LD:_#]VTFPJ-af84G1JX,b_XPc<<5S<N3H4;S[1^/Ba=AGN^1=NUEN3
67@cNS5KIA[B.1aJg;0f0&6Sed2N6-<-,0XC(,O-b\/7]_2@9_3FA,VG;cV/RXFg
^Q#EU@.=)JMQ(\>>A<(6/bfb,M]aa?@WWD1,RS):a9=.L<([,>G^-=XQQg74G1_V
gRd/Y=HRc?^84#B:Jf_U[]0CbXXF8+C^Ue0FTF5IKF,=,]c76E]D(P5Hb=/NM24+
H;/^/ZR&3Y+b)cZ\+Ca3Kf3.A\+;1TYGT^.?Ub.d23-9;59WQA(M[,g^eb2MU,>^
\+AdKB?>4]K0<HDF8b0IJ6BP3IC_:>@?daS\1T?SfK\8fad)H>Nb=(<\Jf4;MGVY
,-:T:0_AN;U#.O8d[[a-Q#XQ>FE&TUVaD?4VZA_FUb+?a6N25f\aGEAF&?<9CFN-
W8T/.<TY-eN3=He8@@:IK2@KU)W^KC=6#+(L)D_SY\CH7G?4/_S]f_g5Y#9I@N]b
I0c[[K1c2&=Wc;VD_2^aCfCX,B8K2B;:(2V5+P?_/1Y<^:_abSa_B9MZ30e1]R7G
QEU.4H<<Bb>b.))XV./dO37HEO955Oeb0>[ZNGC+&R3e+JILM;c+6R7B27\gIcMY
H5&a[_\#)ObA([MD=G4G)SQ:)VW4LeW&B276\7dcQL&R66:/RU=9W5+LUc5](4c,
g#F?YZ-72^C+FFB3YXb6Z&a]c@RO/aHAXU8;_]LFI:bK3?H@\JfQ+g^NYFP_&?13
#(;HHM+=H0(_]?_>F\4+7HSV>F2FcY,S7YJ>c1RAd8Bd3F[L/BIc[1@ZJ,ge)U/:
G=bU+Q<7W0181#D9T&QK14@C6()[;a&Eg91E2-6bdcgBRD1b7QXBID+[(9c39>(5
16d+(IV#\^&\aO=6#Ig;:4HBJ7U+4,56]XBE8,GfLIRHZ5)4KSF<]aZ\KVL4d0\A
W[GE&1&9HM4(a^XdBR0QgL4LA=#[L_5T.QW7)JUYRAGeEI\<]ZD#>a4-:A&<H.IA
LEP:d402FM\5eBZ]CPFTJeAef=g@+R#01UW\CG,Ub5BJ^]/cG#EXS&3GUfaYKB3^
MY+S6d2VaV4W663>C<3Z0QB#aPD:MU\R3=PDOT@/TW=UL1Y#SDYCAC,(^-13FO5(
9\+<:VXKH_]HVG4&Q4LDX?5Aa;4+P+VQ\)^?:F9L&dI_(P7bN6IUQE8S],=9ScG0
DZS[b-c_CPCf,A>+_g^)@?bY7J[E).C5fDQ\]<SF,#g>O]a/c,^YK\ZcWMf4+PD=
\.>):<YH\L,De-)XOBZ5)0]?2\FV>3?g3WZG[\T(N<Q5/-dc9.P9CLF^7)@T:)bA
824b(b&:Q_7&abHLYY,dd/QZN@f<-AJH.TeS)E;9YL+a9-S:JABF@X\^I.1O1BQ(
0F_R#7):A&f(S_aP\(>:ISKfcMfa,3/_ES84Yg02gGRTA-TC3JbE(U);J_aZD>UX
gc+,We+PHKBQ9M^^PCM&7fU2JSJf=:DICb>YY(3@_fL>?L:Q@,a,3W(UD>.WP?Ye
e\gJc)NFD,-9e=G1,NHC1K9UUY-J_MIBH.)/GP_B);D5<>50(ADTB++IdCQ&X6^E
+Q.F5=c=N+GILPF^(?V?./S5JU?8&YKM,4YQG>aLd?O\#dca[eMB)#2Ig\\P?0Ef
LF>BMAJW)5JH[d@:/&K9]a[6-g]>K^8>V&[K7S:I<7#P1A1EReTU=O6aFN[,O-XB
.)SD43Od3U;U,=/FQHILWdR_J_\AR+:954e[0;b(_>IC_?S#\;@gCMV:3ad9;ddB
V,SPM\[dBU_<A.X(bf&F3\H1=(VC/9c-JK0Sb[cZCEOSX76GaBAP_)SVL&>2=Efa
Q9Yf7=@98B0NJ4#0Q#G=2_:fb/A?\DFN(c(XDAT0c(f4PJEAG[VAAf.6T#1_?:Oa
/:P-?]#6P/Q<K9&MI;g.EOOW?[+3185\PY02cI<.PRSLYbOL(F7S2C^>FOSY(7B]
ZCC6@bJ4S=^aWSD?Z,EYH]Pf9VFU>B;[,B7a4Ug)K([Nb;&U;0/7d9VT1c^7^Pf-
XY>QWb35FWS0R@f].c6RDAEH^\:](e<&>[M#W9=,g]@c4\+<,OS5=0YfcZK:ge_D
;W)]d]AF;gPZ::YAc4O\^dA^2-+7)4@>32O@@\0<aDB5(4YXg/>R9b.H-=OF9#_[
M3>>=X\PaMNB\eZF_(BVZ2=f36[IXV&_JGI<LZT6QF.3NS[BLJ>db7V?09-f-1?(
39[)A-IXIUCWL:@M7;9+6V_Z:E7ZLaJaVT66+gc:PG&.2]gG^3N<PSb-ZgO&Y?EF
]YTZd2g7;HM@#bP[TfGEYLbPW:(6;<@^a.(+3?V#]\7a,eeG+X\_O(D]^#M.K=FT
bIU3;S8HO?a6)dN8a-?FccXMMg9_3E.f9[0?Hd=.B?](7:4L^&(9NKC1C,ON5=02
e-1>1CG=@FSH1UJad?W&]()c.-&bH<E+RMCCd:EYaEN#ST@]8);g8G:6&27]AQUc
b8BMAE_<Q/R?6gJMABeBF(^D@eH86FHH?MYS,&Nc=CI9?/YI=[9_EQO3@(/_Z&?S
E_\^_^FT4^.b0A@fV@_Y8,LK:?H92b+d64W-gU17&;f8f/RD3O/bRW4.0+0D+&V[
QG)RB;H:=:NIJ6:Lf/fW2<JSU)_#F8LA#T._eUT5H17ZF(/cD:K;TV;UD]&^7A1G
O,DaY^Q#UF6:U?)7Q7?70&;QSW7K:^-Ra;KUKU\7>8eHZ[-R.g1d66baP1+Fd5L.
,G=g;C&7)Gcd[/J4((CII;&?5S4AQ92=G98BO/1MTS+4<4<SKGe.MGY9TS3af5,&
b5SP6NVGgG^HaJ-=\SJNDg9&;\1f[f1fTJCHMI_B3-KN>EE6/[[a]FR4^+:e7d>X
K2?>R@6a>XXEZE:0>+?H/UH2M+a,&3=57-LbGX[_Ff[_^.N;;;L.XCb>;.6\N-R.
T[0^(^8VdN+FUbNCb9UL[M02>&&aQdJNeM\NQ+/[AHA5#3-86[\:TVB_IN[P2+9^
QQT9&F=,=^B467]2d@fdS2g>Od2[PR@&/[VIKM91d8_R37J@UT^JH=5<B.]ANEfU
4df:YH&L+V>OS/Qba:G5MHL>5][=&bNS8Z\W/?_caB#>V:McGD>RP=&+G,YT5S]#
V/R,PVTD-<d4K-X]-4R8dNYe?b1@=D>5+W=P,b[cK0DG9]Q@W>BN?J>3XVNUQ<<0
S=H4\SZd,aMFMYD4]N\K_X1<&:<::<E7e<cP]J5;^2g7;C5=4-T_#T5_Y6C\33EV
D15dMP:-e4Y[eO=aE=a\ESN.=+72d6D_K;3A6d_Zffg(Q8D&U_8f;WLS95D@V:.P
QFeCE1^?J:TfA9CKIA?Yf2&4)KNGV17U@TP;T,,44D3_G2>5PIHZTCIAON76OWRW
^ZBHW8Ad;A\P?7?Og+?CX_E&(de.:M=^AGPfP32ZgLA52W-9CPH0C((9EC6JPIG6
[_Sg<EPQA+>3Q[^KE]I;_UZJWS[[.=E8c^Q#WY9AM0.\cZBTfFe4.RIIZ2--cCfV
&\eV;\Nb1BbJ1DCQIQd9K]UO#ZSR_)+;=Za>Ff_@XE:4RQ\,0E:]-V9S4G-U004=
bGdJV00FQD[Y2Q-DV_0]g/KX]T^/-31-2W5eVH,]^K#F_QP:@WdL5+g1W-MJSO0]
<Z-T=2;-=bMR>UGN8OBedESR20#/@2Ab29fF+/b(a<9?-7/geN;I]UX4-1JU3GH9
ZH0c\Tf3d]7_#<.UJWENYS8VNdaV0AADZ&&B(#H^^>\9F5+8-)gGLN3H)]ADST2R
M3A>\=7DXWbZ7EcN3CeOIc088\.U6M]1M&TF7]=BH(K+eGab5?K-LdaE1_aA6cRW
]I&/XLPZH?.[1[egN/@U7[Jf,BJQ.+J3S98FAgI6ZB6>^QK_J\d\RH3?UT;TR5&>
>JMGaBG,\WGG@_?fI;SZ4?7&e\^5=Q;-bE.,f.ZKVU;YNKW/PE6cU?SY3)/K0EX2
EO)NDS-/3-;B0]a,MWd&bCD33^BfY[Q#Z;V/Q;UM<2CQ&;ZE@OFA[B7dBW]<=fT#
IDV@A)e810QaV(SL;Q(GAW9QV3d\aHV2BO.=_<D9SR&4dRf(4b-[-eB1+M&DU#OA
6#;U6A8SSDEU9(T-TZ]O]M>Z@:6.Ub]H_)R-Zf/KHIYJ9L,2(@C6L@;U3HNK\8)g
gQNWPF@e:EAF8:GS?9)F@eceM9NI;978>MeX.cTXHX-d=cKC(AB48V(EL-QTGQ-B
FfK9-)B=<S6FV??M;/@Tf2)M4bK^<MBO:\QIg^C2K1#4;L-?GB8>E/#.R,&V+N>a
LXJ[UB22?)I^>S^<BHVO2C&3-AU3Z2^?5FfQe/U6_I4E:O.KQO#BcZMd81ZUMg_[
[A//&NDOOCXcUZZa14O(8ZbY_7+/HJB;IQL6ZbOMXRSc+OM4#3bQdN(Q#0#:c7,:
EIZFX3Y_9^?d:Tg2cT9-K5,[H.GPL[]BKN.]CR^7b46+)6=-_EP[CdY8V.)NNG-=
K1.4g<_/XA0X>TN[6Hdd8]g:?LeX,KDc3]a_H?bPc/&XZOKHOge_W,YM7Y,VU_&R
][@J1N4]Va_O,,HQ_(I4\S6Z\Xb:c##Te/#RFaO<BEP[6M#K/d-]9/6AY]1?,X@P
E&.V2;_FH\0EH+IFVFOTH1:H4-J3E>]R]U^Q\J=LLf\+f4<4#UG?=Sb,HQ)ZH-L\
]TNdO#aY)A(C(0RZ[#::aXg=IeVePOKX+BT_A@GPX6ABeXaEKN+fU+aV)XSV@AW0
U6:;>_5=BK1M58,QDeA6-]b8f699H+34IX<cN]D?+J(dEN5]C3F3N#GF^=dV3]ES
AJKUIKaV7(J0g/FI\BQ1V#DX+Ff&X;<^X_L4X_BfH?TM.a.5bPd@.6a2NUb2ZR&0
1P55>[LIU:.9Y0<3Tb42K(O)UF]^)+T;Cd48POR+QY(N7[-gR_\a:&DMYb^bc3:O
(S2WHR?YWROe1T&IW#2[BO2cA9AE;_+b^KbXAd^W#9)0(,+)7_9I+_@+8c83.Q(1
385S?G+H>GU:Z+CVVHK+V=?Sc9IMd#IZDVXf(>()T+V]S+WL_;0>-?-#H==T9gR_
<afgK^UcOT.:W_KWFcFK8OaO>5,T(c9c20CY.;aZ,S.fQ&;d[/=\dW#8>I.@J:/1
6Ha8a?d_1YBc_R2RIWQ/#KK&\WCI#fb[Y/=;Y:Yf67UJT5E7(aSF)Pg#87,=DN<>
38F>TUV-0YRXZa?M#\g;e;KYd)BT3\Sa2@I9b;W-A]11G@ScGdVDO6Te#\a]gg</
W(3dYe(S0X4Nd,QH>](#_fW?R8O0C@TZGMbRC9-0>#_1EX2TN4:@;.+H\>8Q(7a(
O\WJf;<W9#&@E=/DO)YBQFWR1We6dcAS((]R;ddPUZ.5_aO82)EG2.Z]/,4^UE?)
(^(eQD8TP_@QN_&I-(A@>&T0V)8+5O\3L]:aQA58FV16JN]V#L&_687GKP)d&_;b
2dQ)N^5LMFLO#5]9IG-Y#S?FGA@GOBV&3I[&\OWAE:Q?G)RN6PX_?)/712&g85d:
DNVVbM)5DPRP;+H[HBCM15>Xb\;-PINK;b]4]Q<H#;PLDDEgO2e5>W=^7?2gCX>(
+VC[SKc)[N2\dQ)bUWWF&bcQ;8M=H9-AGYF^)A_F,K(QIIa3fM7UaSUHR^6,W-G[
)Tg\_,,VK]H+)M##H3J?Z[F9YRTWeJZ6TE,cIS^D67VG@]ZUDE&]L/AHW@=/K8aB
[0ecDdZ_L#SE9L_fC4E]6NXPM1^N7=S=R-AP&Z?&:XbVJ)Zf.Y6=YFMEI,;ABdXZ
]=e#.<PH:;]FXf16[#Z6&gL(:TU:0^.BSf[f/<d=.,YE;[]1eIVBRd1]D-aD3R2Y
#//V)Q.)Q]-)#9:#&WDd.GU/PA2+?F42IW^7Z1SDZaa@GIVcF+4Tf7BK\^\7A#^(
GPDQFEMXZ+I<&@1gaPb>E68KQQK>J3+I0>:=H,]?Ia&,16@_T^[?&>)M:I2.8;fB
cMMfR[+4]8.KI66fBcZLSaV67D9M5^7+2F_3K1_3^C<-)]&1<A1<?P-f+]ND3Tbb
&cI?BMfc-4GANaH.V0&X#-6=Q^9JDfO#(LYRadFL,VY.[DKb#WMH[g3R76?RPJH3
O,59K]EOL]?TgETH<<;8?L6-V0,3_?YWbBNIXE47C8dR\??XFD,R75;G<NJc?C#.
a&L1GE#.dfX3<f=?Qg#&UDMS;1Y3b#P5:U\a6=_a+S<ASUK4Q2Z-ZQ=@JMI30>7;
;W\NW9\WLY?B5.:.V7I0bCT3O;4DF(8[Cc[)HMUQY]_3(C?><SZZ6NYSNXgTMY_Y
DV/FX<g?#5bP+QC=DcGI=K-FEOI5[g?,f:>[XKb\aAWU7XFV]>M&@_R5fSQA81G,
?^H0g7\g5.F-7cZLM_]cXU?2N&_[/bgf))D)KP1Y:/DGaG:BN]2(I>f?@N2G\L^6
daPXg/aKES84R2cV(_aX6MD#_LYe>(@P=W=]:e.:Pg@.XFcR@&Y5g=Z70+AbYE#&
<A-82X&B/Q/g9ZAf;X:S??^Z)Ve6DV^AH\XT)7<2bQE?FN9@MCebB8c+CE.=S>UG
=Q02CV/U<fGLD?>PIT^?4-b?eOAOO290NGJ_g62L9=\\/CK^>[&P)3<P#-+=,>DB
N>7_6a>QYXg_26;U+WD9?CPFgc_Y/@5ITVgI&7)TP80J(H;<JfbJ7,N4T,7T=?-L
R>;73LU;I;&G:bQE:?3#7PgETU0Z<&SZM0(HeIL5K(EM4&E68)]5Zd5=;aD+dJ\1
0XU[&\-\@;0(1(R9+F&VA^CGL#Q8I[1,fgU;2OQ39Q@)5Ra<EHg8E>2BS2I-HYOW
:]OUCQLRU9a79=B8,9-;+C_#9:-F5)7Z]Y)N](SSAe+_Q1:c7HAW6ZF=.RZI/eIf
@XAME:TRbPdW.I>8J2AY5,I(aVa^FgLB#D4_KL.\5IZ<1=)a:54e,ZXBb-A++?+c
XQMD-(/\J3&7c+F,^[4V[VVLbN282BX-PWC(>D1)OF9CL4=XUa8C:K2@5f6Xgd+\
_Gd1V_bSU]G.3g=#:.,]N6O/.8OHA1)g@WA/@dgOY4c>M9-1N.)bO8ZP7T;#V/.b
XM)&cO5c^4eY<.4/8WC#M<FTM\UY+.@K<.K61C.U4O<Jf0)<YGP&\.6S_,Z=&-f1
OaMdL=ZT6HZC>aV^P7IH2:.D16JAGX=PV[N1(3H00TBD^)GUZ-6a,XD(d.f71X_^
-KfIcWH6;6R+#P(41+aZ7W0GQCeN<f[&\DMLaD,BM)C2/b(T)O3gC<I##SOD<FFe
C^0fL-J.f8F:Z+=+3Ca&f1gCU]89E(7+NY#:#N\7:ZTI8PLT.UJ]A6Y?^aLDg,E<
>.?^Y;HYP?_I18CDgfYZ>SP/;d>&=MA(]\VA9>?]A)]1983C.IT\aR5Cb0JFBPZK
F/8RI>Jc12c5QRPO(_E:G5[#CGK&[3P#XDPQcB9)<&[M(:;AM/Z7V>:f?+,F-G)b
cC[9,>>.g5Je<IM1(6VSI5^?dO&5K-QGCb(BIPA7Hd(e44VS:+&@:Z];>L)92\c4
e+4=&RV0V[GG]\;TA>0Z6DUT#C[bg?SN&0Z=ZT-2]MHIfb_)@2bETC7c<2/CQ5:5
HNO@\S\8_8bXKBPcd9+R/J6,&/1(G99b\ZHb)NJ00;WTW0W,Z369D4:;5d06IM;C
FU&2E6MG<#A8C3dP[-fQ&?)457W,4^-][S3J-aW,dPO,?\()4=AaQ.@<;?FdOV,1
6YPX,LLA)U)>>X8O@c6O,:PaB:+d8CE]3M2<V3Q(9g9OUIHcO,-8.L;aGE60eBg]
Ag<@^]ga:[1R-_NU7_93OD6bVN5M.g7J&]bQHTT0Daa49TE:)f;OdWA\I3;M@139
_VGaed;Z4+EeI1)EW?d7GgAZEaC0Ke2?4F[RJU=F:\G#)MB7W_S8SW3SVV1I2bg[
1BI:)bg3Z;&@gB_@Z+G>[+aL]f]cL#b+<S)(64[BLcNY,7^<2TKG&OA8dE@51agc
@g]03_5GPHL>BI)3C;L8,_bg\0e.J4#MGc?)V24/2O(I1Nb&a)<WF-f/XW9Q^Z&W
JX[OY^f+B+Tgd,85@5FXNX1&=c1B1)UJVbEd92Y)+AO<]B79+X\T1F5Z?5Q7?JD<
QALOCSBc>;2&S2F\AXI11<RZ(QA;;_+POabC^4>@LG7aT::NNC^32A6:6MVg.0JK
TW&&Q,@MR?5LPb,+6SYU<B>OW\Q;-LT[Q/FXE&OY&5&EfVR(,G4O\N/K6WN\^Y.4
ZEWc>3R.JfYE6A6c.QT)UQ<V_N:>b,I1#^+dcebdgIJV8)WGB^TWgE/<+C;I7+=O
O-QRG3a@+IJ2g.E:>TQG9f(R80#H4F]((aD2H_H&7\HYMW>+?14Q\^;5IRa2geH#
D==?Fd@QK:ZT90/UAW\2L]_JN3cNX:+:&7[T&2D<_DWLT^fG423^-_,3NTHfVXE:
]^G\;<+(7:f,GCg/Y-(T=0MPW^\@@A;NWR9.P^VBKVCAb?J,M+&53gVcFP+E;CTc
@eKUMMHO>A]=f?7-CM2DMSX^4.2TNZ_W^)g,>B6=LE?JJE#A:)XGe&6.Z+f5<[cZ
)MH_B5^N#^U)YBcd3Y,H14Xcf:]eNG1]B25E46@6TR+12/Q.3XTL)6+:XbY[3[4S
cdS/QY4d1(-2@:1?W7/ZUg8XBP3T@/eYS\M\M0<]\M>H3.,N2)=C.C/B?Y#F8/Og
K4g9WF8>M8UHc,-(T<S7=]fd^O>LS\:@UKJe6YPO/LXLK/,6U)dN^34=P7.fPEJQ
,_-0IOF[fG6g;NT5d5S728NTV(a]R3H6_MdSH(11(R[Y#P+f&d[I/T::0)=7<M#J
L5EFG./Aa8f\L9H(0_>cJQWgX5V\Y[9(1\6+0c1/^?\I/[\7:XXf;ICdWBC8YKM+
KSTB-_0WYe8[0^JS\:G4Z)>+]K\:>13L6OM.G2cC;d?M9XgCXZGJ_a1Ag6#LSISH
WY-U#+^NL?J:4a5-Y#//bK=AMe[14GaZC1\+8F-LaeDc7-fPIgP)?CEV@g)]&RfU
BD._=;N+G+ce^SFT\0MKN5\3)VMe1PU_?5VFSBH>d\ee360M,7ND_?SVYAOfU@:7
fe?_VHBU6Nc[c;(#ebGQ=/4PA2W3)^YY-,g;BGcb89H\gML5\PE/LRH<f\F?7fY_
#dG;JZ-1HBKPPKg+dUOPHF7YL\_X[<eU4#d_Q@9O.TQ=c7GUeIA;@bX.,(W)I_[<
/?YE&K\[6Lb9Dg:d],(#U)[8e](3A<PD4\TYS0@];L52SVE\d7Kc?)NV5Q@S<+LX
&-7J<D6A;<[d)+\2(9U&]GS<Q_UORca#;])\ZNY]HWO;NJa\KOVFA1fJQ43:>5]P
)R<Y&f8Y((O)/HNMA2,-6(d+L-GPWQDL=NSJ4gDG>(3DS3^4ZI&&g&OM-F-<SI<@
CR\E[UVg#JFI3.ER#2ZbK&54YN\WS<)NEcNRFF@/=1eYZ5YGHH</A)X_32.82We>
_<&&=0,/Qg@Rd[@)DBJb&_.G1Q\1JM492d80GY<g#7#dV[EZcKJ#-O,3eY;PTJKH
MA:;,YW&>cD9M,Ba&]gO>gSMN,)J<#ES1.(40[O6.9Z5Q9U3=a^6\3DS(a91/@Wf
/((_/DQgd-3Y7e<Hd?c>@e,Vb[;VA+E\8NQ)<;ccU2Rc:Y1MRB6&BP1dO(4N,D?3
1VcD;aO]b;))GQHR2)bY&?-f2+6NgbN@0Y(IdM].EZ(cU=J.U\+d]ed+HW+-:IC1
]&S.#AUK^K-1XfFbTBC2##]8[<M[1V[(B>@B4]3]6BK]/+dMV4#>9.g,/HTSL&7F
3D:5Q6L8J+C@gd2-N:5PUQ^U4KV,0NC?<S9C7,X0L8OH9X7a^2E-B/VR>>RHJZYW
VM][AG[[ICFBAQ1=\GKQ3E_Mc5&H<O(5^S)G<_d=9O8(Mf;@]X;(,5A+SAbN(E+[
eeM97L6f8#D@_=HOK9c?#470H^PQPZXfRU8T)&+Q8Ye+,4V#)XQ@ge;IDUF981#0
JB]7Cf8VR=Pb7EDU6afNaJ?@O]\\1?#5_:B1_?HR4@c]YKfP/KIYabe<d6^\7KOA
RI3bEH5?E2gTfU#G?;.(aGb0YIDaf7Hb43<D]ffIWX4GR0)A(DXIR\8]W?BCcGC#
(Y(KNK#Ra49c@gG,4KVM[C268^/@BM6=BT-=BQcSI[MB9G^f;9G#U)^GbMa=2eA[
=e2I,]TJT;:<P@QBZFVLb;<N40eFFFP+aD?)SFT1W#,[:3.M=D^3F&PGT[f9ZK+7
d<fMNKM,.0Y7@.3)]YW_#>Y_1FAaN.R^)c7eN:_8^]eYQ34Tb+WXg),R+[-?[111
Id3HYI?[ad/YTZ\6Rb&7K=Y?3S:G?1gEO@N>LC>-7>gX3L)0e)QOFMM2-&ISV)/B
:X2:/.I@eM8=?:TQb+P[RZO;d[&_.JT6ZQ+Pg^).0/7BF2Mfg,Pd4>?\JCCI:?SA
,-;UAF+W.#X2WZb4gDX6>T7R/K\5SUTYPddZZ-)8?[43Rb^\S;/[Y&WB-:K&N^[W
(Y.-3@DSZ#Jg-@,DI?M&#UGQ05fY\0W/b8WJB#],BM-JB&);=fd3<K@Q6\JGR64e
/.M9@5aNE.g,2=6/LITbY_^+RP0M@9#U=Q/IFIgQ173>/EOaO:KL0_D=&^B=8O#M
e_T;JFd3.<b0YC.^>-D;^4M:-fRaA3Wbf.))0cB:=/AVB6_[/XUWS\C,dKGYF,CQ
&@CFbVHD1aS85@6GSHV20f-KbO27;E.VOZX4BdU,KFCNc8gG_Ief\/aF6L[=#RdU
^L1X:cC#T9&W@#e4Zg<>/(N:?0^T:@CZ8EBW&Qa)2I[bW0[X95744cT<aLYAGY9,
Y^C)66ReFXaMda9XM63,NBfZEI@Tf8La]Q)b(+#^OCOG-.K,>.AL].bXGD[,WD[,
>XGL5/KPF&&ZYg6BQD73^S#JC8+6E2O-@YbEa<6FPXd4-<a2GMTLEK(N\/bNTdS>
@_L+f/,aQO<(0BLgJ-D(C5:-2+U?4Z6@&32c;/&G^D_5D35ZSUa&EFA.^MC_7,-8
V=)d)d+9VZ@YdOO(5V&+[e_D]aEG4K\bWf]T0T,=IYNM;3f5&,4D+[+6U3OC<E6.
;;Ud:U5d61#LSR#b2)Vc5R/Z0T@[UM5JJfI(dW-7JTAP5MM,R\0Y_<BY0EA-bRL-
[Q1VeBJE+Ua6^Qa3c4Xc<Uc4-NNCTLDfKd(cF&_E7OeKPNM;G,45NER8E2=Dc;K1
2f0,R5XP]CA(T<C+>9f9GW)6_XO.=5_f#gT?C[1JX-7d0cc[-3c8RSg?^J>#-fUe
7fHHTa[+.aFIK=UacMcFYeIQ5A<P);dDb:7+XgM5YE>(W[a8/W0C/TE?0.5eZ+1C
RV=I@R;Q,SKX+=17/ZZIV0T2(K59PQ9B8g,?2>Wd6@-VJ;9+MFP_,X+fW3#a]H8E
2FBK1W>A^U[Q)a5\3W13(#/,(Q#3c5@<,#<>c)^:K(T<3[FF&M(;9PB]W96^U:HY
/=,[<S.GLKBc26;[CB.?EU=J&b-gW2aWA_#De6PBA?)^=3?\58KIVNYSOGKD#\c1
N(#d6Og,1g0]Dc1S>[Cbde.JMBHA,YZPY86YD[#U=^1G@XJDQD_QE=BURaQ.IgD6
U3[P.R4Qf:+Xe26P1U-XP5=L=d#M.,IU=SAA>WS+3BQgaBAS(gc8Hd+N594/P)L<
NUM-WQ4.#feTF+bZ??:_Q5G^NTbSeW<[V>b:MJ>S_[3E[f)(V,)77(OU2YO@BWK3
OR4g>,@-9&&<\LdgE10S?7Tg>eTS?QX9<SI/=HJAD&9EXYaQEK<UBH-5QM&6^BT5
/)Y16=b/_@;4//2.E3X8&H7@;&D)f5SX>_aZbQ#H>YKZ#^K.?>K?1J-9f<B&E)bI
+]+>([<VaQR9cGJ4/39d@TD\>UIIQHY1ZVPIa(KeZJ^\]S33FP:7-K9?3@FQU]=M
\TXOK(0^ZA^<I4+3H6;^6(R,=1IS>3)9=5fVPT5\KWZ/,FD_UG,+\@a)O+R1_:74
<b4CV8aP3gIX2c-/^^c=a)=cJL\>?YeUSN,PcDY_#.LXU\SP9I8KIZ)e3I+1A+I#
WMSTJOC[KCH<0cN+g@YHRc/.H3O:).4V,0#/_UHe&Wc19#C0WHgWI&,\U/;/MOb+
IWe;C\F/BN&OYRIcJ(U5SGgfC,V0->;:@>R8(^84a_LReXe29GRH+-8TCQEM=5/=
VQZNTc87W=FER7=?6,,=Q?c)fgI#R//=_gTFYeHA1M\B9_gb+2QBB3Dc,9K([A0G
1S<]F6f_5H7TR;PNSSCg97@2<O0e<>X--<-X<c[H,e)KH(0?R9F;;YP_#G+c#VCF
Y-X_Z@&OQ_CRO22)QdKWJ@#1N;^VD)XF&R/</K(&^(Ddb5;32fCfT969HI;HDW=U
A(-P)V^U027-f2Q;<g5+f/1V4<#^CF3\JRdR1.B5&N,eL89K0\2WeeL3Q0_@N,_9
T32WTTH(A,..eV]\:Y4+5H;4Ac8;Y1LbL^K/LBN@:#003f&R5DBa^&g#RgCa_g?e
+&?\^bA]3,1(#5Z/(&LK/]SbY5\:6Q&cfaPSUb^,9(RQg\>D@2&=:B/g8D,6,aON
S4(PT2PSKA)5Y#cOHe\M^e)Q99USS]^.F\KC6Md286-dFG:]]]7&^=->/EFELe6G
EZDcJe,-(W]NfI>W8@LJ\-eBRd[fDeH=6^-=#)Q;0DIU8@^P18R@.\/fQ5Y,=#aL
EF)).YMVE+Fe&86d69a7/8P0>+ADP/2/&WG6LYN\EZa#\P&aUWLY[?>K/TNDbMD9
<bW^cHH=WA4RKXXDe4ISaY=&N[M=CF)I>>5P\P^RXVD;S&gU/\KYB5Y?GI\+aa/<
O0D=4N2A=/.H@=eF6-9a8ROH=6+IZID3]be/AfFVf4MR63J-;2^GXCGXXH6?F1X]
4Z0WZAeT.]I1Sd/C[3d_?E9G=]gMM7(&W6;g;\_=7C(8U-TS],b4Ta0Y@DR\-JOQ
5ff]37/]b(MSZL92LJRg6_BI1.\J4K71K49Oeb3\=L2QMWRRg<[2O+0f/-;@fb1]
fbUd^(99<d4FeZgMJc^c8:GTd?H(L<PK.9BD3P1)MePBNaT+<EF53?#gE[VB#dU;
\)>P/I-?P:S<@MPBD]b>bA8gPd9NT5=;&3+e-IPOeTT6@=AH=.2EL=-gZ&PbcF4g
gFeE?Z1ae0fWWOUJ)33C1-4#c-<V3<AdYe=1=F,)DeYdgTY?I=MUIP[E0b5b6Q>&
8F_KGPMKCH&X+.SX7^LFb[^_NEMBC1HXWbX\S1#14-JfTO5N:E(L?<K-cdB6F]7+
.eM12DI&dUdQEegG?&27OYTW:)>#g>=1&04KXT[:AIMaG[B[XYS#\/0WDDP^#cEC
[,f(;M2T+@#&&HeBV4FbCIZdAa3:E5eP4.&3@M(?b9Z)_35Q/ST-3D2W<IgWK^g#
Ma7LCC??9YV]K(30a1Z6DR:WJP2DMc)&Z5aNDCX+US)gHgO8QMB7ObDcO,.E4?FN
BCDKV414SVe?@c[V(+88R-YES(ALNOE#[=J+(IDab>5SSHUSF-^^Id3_ZZEI?DIX
89PKX0(Zg+&<^<,&),=R^[VL8FWaTB1Ja6>=&N\NbY/JH+.+=7G]e+HZ+SK&_NQ7
;XMffT[\Q=R-d\a4=,)=d9??[])L?Z,TZ430DR##2S\,c_Ra.=TW5&??B[WYf4I>
DR\JLaRXFcON<cREgUVHedZcXdg+VY4.f6L5)>+#A=E#=U,efZD0P,J,>(X)e?)&
M(.43^\Q?Q=9\f]7K(SH/7[P>QaHRXScd#D\Bc[9I7Q[S3=cea4\BP)^)0]_FS-=
Z0LHdGHJeE#,D4=6f5K\PIV&^UJNHVOc8>H<c6_D@/>1@(dCUa#PAZ#;;g0@WUT=
/^5T&QC[5J=X/4<6bX:]f;6NOR2_:[+0[M0CbTcgC/2NgM,6DZ#=YC]/\VL3?1;)
[8_BX\@4K[JU;7IHHEfaM4RN1?O]d8.>X=8(1SUGP)QVS3K>JB40Pc)D9^DcE#VM
@-cbcZ:RMBXdKe#4KOSG72?<e7-4MI]IR5T)8aZD<&>Z\WO=6U/>M4?\bG4>fDVE
\QedX2U8Cd;7XN1;.1C[(3BA&\.^=QO7(Rd[E2>+9WAeg_IVNY,K3YA:b;0Ie0FO
Id;_CIdX.2@.9d-6^D(Y021L_X=.J/,VS5AaW/Q)L/U;H;<\&&R)V><8)B3+61&D
Na8FZZ3#d[b[H@_3\-7UbSS83Jedb;/f8.K6=YUDGUSPDQ^I^ODFU/SHW,&TJ?1=
@2&\_+:J_A,b-AZ9#\ODD3J48P@E<H=KcV_-#G,;^b^K10\SR,.1HFD8]DUbKEYf
d1]>E28WEYb=44:SLYf,b@eHEGE8.VE-;g1I<.SQMPQ)WLC:/>_;aIM1)=\<#c[D
KGZ,;EC;(/HB;BN/U4KICBJ&V6.;W?&SW)OK0Qf-b/YR&f_b\+S]5#c]O=EI7I?=
28V8R;S/1b>O;BG>Re&W-:U\\B&?)50\NJN@(O.?Bg>RUC^M1[@HN=;&O/0]COO\
8(F.Na0ZEDW]0MHf8ag(f[[Ac5(D2>AJc622:VQ@\[KK7W_0V=(e.?U#)IK.SNH1
OfWJT5(1J)9Z:Ic-D\IYX)@PJb\=X0LAdM-FQKJ4TDDF+5&UHTG\PP>LC7X&0QUe
Udf+eLJMReEEEL00Q&<N,<&8-[5E.\K=gOLeBO9WH?TBE8>a(63Ec<D::M1Je6S?
C_8@b&KB/(AFJJ4faF-,IKD,)IZP;b>Te>aBTbbH1MU@=SV]WgVe1=AM7Ue+&L&?
I@H4XOD[2#;+VIJc5GO]DcRIg3Z]M7+I2bSg8e<804Te7L+E=X#:89-QH-46<Icf
XgIaMV@2CJcE#^.EVd._SF:48O0W^A,e+EY[,X@Z?._d_.<LHS\9(=5#@8LG:]NB
8U.=87TgF/9()Q8eCH_51W7YG8+T&\W+\,JEacDZSA_,Rd=T.Yd+3PPWT.Q7[:SF
(Edd[5AMEQB1+YJ]eAIaF#&\/@OWJI<#,#IY&]2@_9b-SX\f^6V\P&cMP:Ifff+c
C]Y_1@0=@&BKW7E;fC2XL3B^EI_GF\P:#M+LeXP.?+_U9IR<TGcI^+6_)<J)U/3.
S[RZ1A2ET\<4U#+HG-<-7/#;BU,D#9g[T8cLSA+de?B.>,dCR.]#NVE&(O)/+agb
aGgB35/XQXgB=F=,b@WNP735[)8H)OZP#Acb@\g,4cWdY?KN=PR4;)c7#d417f_Y
gaWN^4c?0G2(I/5XYRZBd4@EG.V31>;3-H]Od+CN&eC6CA4]M,=Y53]G7fd64J>G
:D]6N:E),@CQ:LJa7>XCK:UMf@MTF]2?+4O8ECZ\+_IZHPM@\N&SRJQMBI.@2dC0
eWF2JG^H+;VC:P99JQ60_R]V#ZSQ6+E_8OT^b(U[?]#Q#Wa(ERdL?--QcR;d1f&G
RRgP<[G>I\@:<4S1S/2F6_6AGW_1;4faTAG?L5GfHS2.D>7<((+ZgIVE#,=2VX-B
7_4H9:c:aA1,KJ@IQ,+U13G?:MP3NV+2A22g84&O:>.J9gdcY?[TGZ:5O3TdRe[\
4f(YQ].L#NGgK;<d+:9\.W9D_EEYWS#.>fQ8B/S1#-KQVcZ,8R<^/6OK5f3d+\2E
A\<8JT\Q/:](Y9R29M>d_dZ=KfVK1bOQf.8gYFV2I;0M,X]gTG-O>AA3U,@cE//>
&9JU1f/Kd((&,@WU2\CK3>2g-U>WYQ0Y1C]KeVD;8.TQ;A?L-DE\@LI=I,Z>a=VP
EN??K;)Y2#;WC&2Ya,/4W)TeREH>5(V&dMN5dg:\+-RR19T3Ig&AA<QIH@Z97[MK
,=N5=H/\GV^[Bf8(V.XbBL23M&/:VeE-PH=:8T^VL#9C9;eJ2960Of(H0]cb5L@4
.1Y(C^fC+MM3ZKegJB]K&_bV;ODJ#XS1\ZH8B/9B);6.)@>M5I^3dLU3:/5#PcGG
U/7c6=I,C=^]@d_3A=K<P)LgCXXXWNW)&TY]2M86.a@U0.Fag<4(Z6I(:9FL(6=g
5]9Lf\VEdC@Q,3c9](aTa(0P6<>:b3DEg.J2W4TXQfQ/Ma@gARJ8OG/dL+</7,P?
KXC6@Xgd/dTMaI)(?B@05])KKEJYQd>@ZLSeE7_=/Ea_-^CX;W/4OFZgGLJAXA:>
B[:KT@\6a0(C[-EAI-Y4G7C.^:dM[]C?7+&b\U[@/>fd?O+^ASCbX,EIBgMc1L@1
=Od.7Z4G31VQ-aBKT,c^-gLJB4LGaH)D.WPC8^FV]?ZF1UDEV&gOR8RHAE[Fc,?A
W;U8QCL8-F9H^.L^9FF70?(XR8]UUNDYLgW#(1^WP_L@CF8B[d<4eEA(N]Xg,cf1
d\fEOD92]R-5CR1;SU;f:]EV3HBC2X3D/;\JN\^f#,d>V-E.cZ_8O?HIKFdfeBM]
M[,ZdS0/S3#;#<cQ9@#2a?R5>(d&_6/B>I==#<:d^(O66KX:b=cL6O7@]/Ib#]cQ
8N/1LDN&g(DLRBK^54O@JTJD5>J<8=Z#aD0^UUYF/TGYcYKfeMJE\IRJZf\W=VEC
QEPbIZ2V0gEL#PB4RI(2::T\<G)[>Mb19L73F;U^-d>H3FU;+L)4a#5UN_;Q./E_
#gC0R+]Y2_/:2\SM&QQ9_VCQ:g;VAW,5-MZD19Oa1X/V-AQ^ZX)X-?<Xba[2^EOV
4=bcMNQM]IT0MdI;#Eb0\V?&47[Q>&WB_L4/^1>)(:1DXZL0OY3V=G7OfUR=:NDR
DQ\/&YSYD)SM2WC#DIN_#9W.NKg&];[EC_FK2PULg8GEY39\4@M4-#T(W<:W(1=b
OAUEZe.EcSEV+ZbbN5K]#R:bfKNN>BX3D]C8IBaN#USW>-)COM\]MTXD19e^_[cC
^eFP>.753eCD+8gf?DTGEGD9b67Y;CV0TLB&IYA0;.Ba#BKN65N2>LZD&85J<J,7
7&@1EeaZ7TQOV7D/Pg:aQR;R?D@@.Sgda@QfX,=X2625C^gRf)[7a9D@EO0-8@(5
A@=^BXb&48(]^D;5XZRRT)=FW,GAEg&9[&KG\=X,MNf=6BQeSWLK>M?F_IdJHb2d
_BW;]:Q2O,J&e2U0&)4bPZPWQH9DIGI,&(M8:YU5+SMZL2@cFM\@+1ef9RN+dUeL
(Ra_e1?#D0O)F3,2WBNA00Yd96^0e=[Ye+<bUY9Ac3-#;c1M#cP_FEFJNfZfS[\7
7c2C6D[5&aUNV#+3Tcd?7fU_Vd/(^4aP&1\/)&<2BR_BW][)f#4\,__fN</JOW@(
DT^_-O^J/?6]bgXE-.062[ODAa82(fU/6X)?J/f+G-/0O@WYJBg204JBc:2I-.Sc
RCRWLEZ7?P+]TM@OC.:N_1.+FE7aP2OTJ9H#QVIcGd)L4+a:S?>5Wc(GG;X^XX;3
NL)db/2fN:d\4;6BW6<_AKBKIG+LN:\#e:,Me24?HPAF@C<f(+51:8@TAF-59D24
M(GeFD0#+H2-2ESJORg3>6dMH36(JOXX.[c@cc]/8S>HK=HF1M?Z[e9D#NS&;3DJ
6,fZ^c55=P(;MV1cW(XQ2#[>#XU\>3VJ0OP)GVc_B3eKH>]GEK#0XEWO\4&PEO4A
P5/J#EW0;KX/[@K>DcSMI3?Z@Ye?Y&NUWPE;GU69=9[]J?WVY\J4&ED0]R@Jac7f
SUDUIIKG+aJR]0]eW+XRgTdbg(BZ[eYCDY&E<+E9B22&C@@f]S:DW2DAA6b/\Ze,
:#Gb2/dIcMY=,W?>PPS-2@H.K2ZPM/B\ZaK,ecfFR:&PM@L:K8G3e3I]C/V;U0O)
a1R.0=7C3H=S+/RLKM[cG<&1-:76cOOT::KDP8:G<F23Qe(BDBd\8aUU5MG7fPQe
5MYN/BK:;W9VVV#<7a=0,8=N_<gEGV;dB^QBB[#-])T;?<KE;KeOKG2_J&<;f\.[
[<eEcZdLI&6=Z=DY[>EP26M_ae[OZ,K=?Je#d5(NVCcg@X@E4f;BE.G5=,VQd152
b0P#TGKDO\PTDFQ^/eRcX(=9gf.B,X;4PKd(_aD@-F?)2f+C)2W/Uf;N0b3KWIO)
Y/RC2GfM/C)[8a+B;4=[_]P6ZM<99()Ed.P#GRgBb8O4YEAME@6@0+[1=W&7WHP>
8B[a:PL@IcIP8N@9H\aNC,>+ZePCWaY_ZIOG0dDcT#?c^cQ.K-@5AA&N.4FfYTXg
A+-P@cSeHL5J<1FW[S\?eO,_Z6Gb?&RKYTf/W3eN0/#&Z4RK5MAb8c(C86W>Z3ZJ
OO]?GE9]c836.c.SQe)FHe##Y@DRKB,R0:g-^46[aNd+cECQZNU&P(bG4/VWBYS@
Ef0QR;Yg4_(_7f0fT_gDReR_J:9P.-A1(F\Ac1B1NC4IW_>e^R]G2bL8G29B]M3B
d2JU^R@QdQFW#b#E_ESJLLCU36Sf&.?@[g3,Cd7DXY1QDYDgWZC?:+2[(=2gZJG1
+CP]BI8</<Vc4\LJ#.K,\ePNOG=D+_3)OLQXf,L&++QCKH-.fg-L(MKC5S9HGVN>
C[A#&>XBN1KUSV4ZE?G)4OL\8AM>(8<(II1AT()gV+UEDcA[/;+&)(GVVd[4G;+0
0<MS<L2UU8/V7.>H;_WO?)SHaCAQMdP-YZABWPR),A-+R5@\XKCSW3LeIOPbU3O-
4M3+0g+AV8b<@aA/c]b:ICW1E9I3VA\O4&3Z<R,U_?6/@;A:6H]W;Mb7d-SR\Z=)
&EH5:Z@ZW1\95[bS]ReJC)-P\^0<N6TFW<,1dVS_<>U7I(K^9b:;XVN]Rb1<_[SL
7&01@HX9L[SE/Y=0X;^BR]0.XZR-9cG&,TN6&S2=+[=eNBVD?/QPO@;S:.0e1L/4
,CE.;]+^YPF>EaX^+YWX/Q^U@P;4K>(L0CJVO9?J&bCUOgbF=F7g3D#cK>VG<9b3
S\EFD;0FE2;7UX]e9N5^FQ/K7P2CCI3&>eXQgL@fdH0\,8,-4XN0C42TgD<KM-18
cN[[cGVY,R]e.NPRO9KI>ZeA?QU@RZ)7?-=&R;9]I60HbN-f()#CSTB^BSF_I(9F
0&>/3((2SOSEV4=0)GL,RbWcYRNO>0VVI33CfN3M85dIKb^g+TL1Z#[R;IXf4_/T
b5ZVLbM:WD&EgB[U_MX=:+2T+^&.RHa[0P;C1]8_H,D01_E&50:09>J][0dN07P8
(Ld#M)OI3FY15g#/TRIU7OKVL3=X^+8G@P]CV;.5TQ801]^gg3YbAP5F#<HdQQg#
PG//E^.W6<<MQ]dZ#2GM_K[SJ+;@gDVf)\GZ.cd>eFIDacJJ#Deb,3e@_B+)>J1<
Y]@>0Z6=YP<Wf39^Xf=313OC.BX5EEGWFI#+>]QOO;(S4+DI\#H2>C,2f+OeF21B
;(c;K+&>O0?bAR-GTe(bW4\ZJ)W^1O;#1MY4BE],T.A>Re&;>H=-WIRB=JP,@:&/
eH@Cc,_X3C3aUd^BB-T;-BeB93f4A:;P73PCWVH#DP?C?7Q.:D6Y,W.7e;X8>W6D
AZAE>a[A-+DVH5D(B8(H)]U@7b)HYMSFPOUN0.41;d=W1-aD19OdT+2KB+/#gdNQ
>6bH/;b3[F+]\;#H9BT_W4MNQD<1.._c1]0LU-XeAA:9&ZPIR#EbW5CVUKSD.(AG
J<3Y7\CLK0)T::?Dd)Jg[3BV(ZW9gF(Sc;Y1?gI)(#[>PM[T4?ZGK5gYJ?8=-36:
dK2:1GPGTO+9L5QXbgD3aI<3FSI<=G2Edf]d4;WA81T7^282#F/KU00CEIN>g5b>
Q2:#MeN8(e14g8F&UT:XLS]Y/##O-[;]9;_@JF6OD5.C@B1>McaM&Z+80Mf1a+5\
^G-C&^E:QJ-Fg1Cd@AO0&,AS^PK:9ffH.9IgPaL6CD>OHK#RCLKD>A0Y<6c6)#)2
LJGcPHRJQ@@V89FHP4^fTYXD)GD2Ra.d18A<WTUa:U8@=AEWL;&KVD6MBCF6?F+E
#NEf<a^[RV:C?K2R_9a[?CE99#@8QdNCN+;C1c9,L+\AVSITRQ9W&Df]ICX5A#62
fPW=\3Z?C_]CEU-@VBeE+17+2_2_3.BPGf7E/=Zg-?c6P+cS6:be&_WI\E;cLY@D
^c?1H#ga2C.Y#W=#<_F=R,a1&U3P.g<f97<(O07_gf7]-I1ER;6R_#,E]K>^\LC=
?UFI5N1R.X39e)OUO]QLA.b5cW4GO4fM6e<W1&7JOSY6FG,<M,O:-2U)O=Sg/1;L
c@)b]21YN((QNO;@0:.M3;R6T,H-Q\@)Y\#LY&@N\#YUK>U&=g,QIK/+E,3+K&&:
1N7IW)D?@&OUD=UQ7T>-HPUG&56/R9E70#HUW1#4HKUI]+<J\&d\<g\I6@=e=AQZ
bSRRVGSZ/_EN/dRYZ?30<ag4;7J<Wg)-D1:-958ERgb,>Z]NX^#cdMDV(;F3af7^
cHgSAL/LA9H+FWT58Q7;8VE)=If;^ZgI#INMBO94@#XI0/^SM@V106\C\F13)gGI
H)EF(ZIWe&VdAT=VK)#,1IEQOFDO=[JT(GNd:Rf_E2c+E^?gLcN;D?YNWT@VWd^5
,(7^gU),g<JEe4-+Q1?;b;)H#49],>7,FI/,SDAU=O-+EC,CN+[fA5=.X?#@BJT6
\V^DggJ<Ja<)B]_D(0bObQ7(VfV^6FXL^@aI09DW5EB+g8ELPMX_=G;2?\6)AH6\
gC:cBXM;[3GKc9923+fOda^LN-a1FEIAEE/W<@06G[ddJ#NcMg@Y[Q33+2?67Zc2
OL-F@Wc/>7Ia^R(-4M@0&g1[56,Kf;:[9dcZIIa>b_NEF:ZBFK-H:J6+<Yg9>,G_
06SJf7?B2@Z7dQc<?L:ZI1]DbOS/_3.8OAacH],V)ND,G1TT.g6;ZXB.E>\g35DL
/39CcOCU(3L6JYd1HB?4I[6SFFQg[>+c:<J7YQd9@Z9BQ_d86?=^1[QF#<Q>9Y.d
5JW86<6/>]8/,153.Y#:\BVY7O]HVfHGZW9Z[e7E@)2aa?#;7E;;Z><MD8CT8=,b
:\H2]DM,\fJfOgR>IfON439)9;RNQ1I\3/YR,(fd;:=)W3>AE2&_McODR7C[8\(M
GLR,\H,/a^191\]UBFdEBWMQ?_1>=Je\IgAHTRGI3-eUSg?804N<2Q_2R,/E];IU
6LA4aN+@dUU=b6c?N.5f=&3X\Y0MHV^7ffZ,=PORTe:<[eZG8JGAV0W==6M0U.0g
,M0:XJ(5dT0GeWa1NYd&A(,b\).94E-cKW,;)MUK+ag4GDL32.?3I)WS@,Y?#7K-
<QeX18^@HaTf5.DB>-HGdd0^2McdFZ3D,c+^YBcLQ\V3G.&@-4>BIZ_:S^(;VZ8N
,A1\6++SR(M3[&G-fa_CR,;g]/@=.ZMIIKQf/:F-LCM5MQ>BE/DT]A)c3bAG@cEg
9a;GL4Nb?d.#d1c4#IQ1D9\HTH>Y@O:Id^L/?:&SRg-AdY/e2e_^HC;#F/2N+;GI
H:L@OQ70MgYWCRF\/5P\C#RRU&<UeP;QS[2,?<U@<SW7=+;eQHGcZ_^7W8BM&C6,
e-Ee,AQ-C@>@5(Z7+\FC\f197.fbKf@CLG0IC@Wf0J58A\7H?4#==Rbd)>Y;59dU
+7Adg-#HY6QUd0CcE/-YDF(UB=XUD2F,VU_de98.4#6;MM4B7/^.;b@9<7Ng80?G
93=ORf1+fNeG)3[XR)#1BA9[.,UfCD5f#gT1.b5WBA&;+07=&b/Z2R3>BF+Q;4YR
eaO/1e+@.18cC:6>?ACNL&U-W-DLWaH3CUGT;G\-7e(M9.-S:(?6c8e:6FSTd<Af
Q6,.\60IW]@A-Q#R@V5UE_C0&#YMcZ;VGBLW[&6@\=+MgebW^>.EK85]gYH4O/8Y
bRHW(\=WYC#5&J#+:D<#U@eN0E7&-.JG0WSK>db_KF+J9(gUIdA_3KW9&BD[PON&
^P6\g@<P2+WV^J(\84#P&c8O<Q?/G#g1D^9cY\fKY^8LL6X\P+/#/9-U/4O4E/O2
BS5DX()Xf+WQ9NV3W4C:7dbMCAI4#S)fR)]OXB7J3ISbQ)BH<[H4/A8f1E8g<LY-
RGUH<)B0FdBQSIJ9];]G@A4/I[2V8YT5<4I-C(_([]c2(d#?1M336<PKPJ[U;9dV
=J]a[a\HV+5)JOU6<LXYJA+?DU=4-cDA\fMQZUP49=TUg_EJ_MRIO<N^N2VAZ?.X
WXL.a950X]HgDW>3VK1C)[e6@ddPQ.A<L]Q)6(Q.PfU_RG_J_eM6F(,>9GHF3[4E
_:,,U8gb+6XIL)5W4a[=W_;YK;ASCbHGC8(cZLGT@X^4>8&-f5SIE^..f+^>KA:,
\K.;@,U[;D@_MJ62GAYA?#S/9V2Y;A&aIUE,8D^Zaa_:?0a2Ob2Pe(T?F0R/d4d/
NUaT3e3-[B5+S9,]gE-V199S7Ha@_]J8SR-KDB/Z4=AYL.aIMb?6:ddd4@,?T6cR
1CcI)(,c4VRf?DM3+:4abPKW4<V?]9#I#YdU(96\-5D3//1D9;F1[D6QGU/H;b\/
X6+EeX9P06V@721,,S^,3.@#KZE+.C+Yf0F).O52;OJA/.DXb;G;UZ@^54=ObKO1
25>LJ>Y;f:BcE/O)D2#4G>HT]Q@P3Z>;NZeeQa2UH[M?@&2(b.M+F@WMf2?)U;PH
S_L.^a&T<CRMTTS8+#;a8aO3YeXR+:+.L2W#V;Xd.V(0QPOLaR4/^X)U)c6\,(,-
@#NS51I(#^KE,BC@-/Q;d\.5aD/5f2ELI4J1MS]IT3&fG8UO@1?G\P5L).U4e;K\
^V.2PS8DbJRQ3;;?.<#IRNS6G;B>3=?3-cP8:QVX4)Z6Q^7ZCfa3^#:>#P9Q)V7a
@S<1C[e+<e__Db9=)TA4)bOM>gN+0TJa.U.)[/f4Zc#WG.3CD6W;\5ZUT)C7GCEe
2A94ODJ2cSa\G/)_[EW51WZ:5BPA5/7IS8;OLLCT311\::O)^7IeMXKY=\Uf./NW
W^eV+=_Q<?=EZ]8bIVW<>BYL@6C1JG/6e\0F4X#=S=+_X<F83E,cH;JU]Vb))I@I
;PbDX(\2]=?SY_M;0=B7^9Y.Q4-=aMgVb(#Rf]S8A;UYFWIY21/T13gU,Y5g(aJS
4^>H&aYfDN?Q#?;T@L)7#Q/Obb&5]I?a?LM6:2f)FA/3.B=:;Yd+_X7d0:gZ3[4F
1+L>]/86XC99@+ROWK#Zc0WQ@^)#K1OY066XbQMKe2.,]LGT_;d,XOAQ]bQ6A>(4
f5JW(NgCC#KDD,>9NOG?L&6ZP_e+?a^>W7OJF[N]?N27R_71QO4.F]F(LD/E(g7(
)414E=NJ8MaX9@OHX7^&I=C\L7OXbSbLL-K?HGPc#01;LFcf>)UZ>)@D[2C]]g_7
.E5F4g_/P>U(1QK9C[7+7d+,[)QcId3:G7Mbe<56QNK3D3Y.#3<;#&6W(5)W_@M1
V53W;Y+=d7?2&0[HG8,b8DGI&.PL/f0^He7+g5Y#ODE@3U7[/XMXW6R?dQ1KbgL^
BdRH=2)/c;NM8?)H)((g^6.7@J?@]0^ADf;WEG<)Kf[MG9dQ5a@]FTM&;#X9.>J1
SC]gK\d2KUYHRdKAF&L2D@Y;e9M&^K9Q[2H9W]68d7P\^YeF96Ybg=SZGI1\dO0,
#0[#.,U84/g(2H7g,Bb&>Ya:<66^79Jcc[f8^e51DIJG)-Ub@[(@.^-JS:;BC:H(
1DWV:e2M7</A,RfZTfag#<)^[:37>7P4T5;,c2PX@CFW1=ZX+K6NP1#9/I?ZZF=U
JXg4&Zc760TdK;.dI>:7B#WOB\\Q/gX;1aWE+EJ-J,&X#B#&-:+;=dQ/;<)Hb;V?
5Rf.-+>8;KZaFEfY5]?2;\d8a44G.HK@G:cSRY(U<M5:6eeOQ+Pa2@@4RE3CV7:6
e4HH[_1eA<27\KXG<B5b-gdVeN-,=,2c:/P/;6#AVMb.5[HJbO>F13IG=IZ96bGQ
PL8^_4./BM\+cSgI?M9a:QJQH)M&-]DNf_?@32[?<1G2;Z9E:^GL20<0a<Z#J^8Q
;bHAS8#bH8M_,V3:[gCa?OH9FXO:C(gB&Mg9XL5N.Ufb)^]_UUI5[Kf#WM-77SCa
LIZYfK,/176E_Y-@H0I-Q1Y/0f\aeC]MG;^,NN(,1Ic(D3Ha2A<_VY+DK,=8SdHM
0^/K7G(3GQ<_81?Pc+Y5dYOU@.KWc9)_K.^K+\DAGL_<MSR:La,ZM+8D2IV[fOMa
\1CP9/V2_V=U-&N))BZJKDICSfT4XOD@FS<HXB:VXUA5gFX[DW7S4)Z6B0b^IfGB
2&DNE)RE9W;TX>QT+]#MDLfYd1(TJM#?8:TO&aXAFYS8Y\MPWM<,#<cP20TS31H4
.eDW&cJ3EJ)(295EQ+g1:30NM4J_34d&@]M0XNJ<R,BD[ZfXfZ8RN&93XE28II-;
Q@Z9dZXDSF^aNcH.-+LNW?TLDe4/8U6P&6O4[X#=)bfO&&C@V:>3WUHOR,?VU9?I
/PgF0=X@NA/HR=M]YbGJ)6<?ND2J?0#M(T41EC89afge_(#9VXgb3#>@,PUJ;R-f
WPdd-)^O=W-a6BUVb\Y@9WBER6e7L60;(1cL7Q+^TA_FI(Rg^d?g[MZD5O4UcYRC
];1EAOIF>J-:UNf:G?+?G)^O(X71\+&eFK4?-(F&W.DU>J.PWd515F?G+dSKS[Q:
dSK-C=C^NO2XG3ST3cNLNVOf&A+>/#Ze1#PNHee^g<#\Y)e/F@=9(dg(P8@cZ1D8
0\0+A:OgN=7Sb>AJV796,4U/#?8+28FCF6EDPM&Nb[^6-V\>FS#Q,.[9)e-/4G6K
(/Of\4b5N=5(1L5P0fIV2BM6TZ;]@F/<TKe>@PbN-6#2;:(TV(D)N0>QgYM&GZg)
cZ9(O\UTBJJVgJ@96F^^Rb@QR&/6YaLV.dOLb/3)aZWc@;g^([\[W1RAZcO]1DEX
<c8(d?+W4#Ab7A[=BW22G\g:I,=cA(6NL0gOWTQdbNdB^N,EV><&2eYG3[G^3?93
]&(P]d5J:dQ&(f<P4c+.IET\cMK,F8I\gBN9[,S+.;WMWMbdS8CdO=Ra[f;Jda0S
&e?IKb4W7c]S2-,2CD^g0,,FZc0eLWXW<1QQb)E-^>]Nd^,4TgIN:98CWOGGX=\,
&N7<#c&-W5:6aPg80?NZI4FgY\1GAFRF#M(69JB2,dZ^e<K?TP-[6R[EPJ9H&a2/
<G08P\F@#N.FXADE03Y_R[T[NC\+DaT#[A=U0D?Sb3[6Hd\:M/AQ?8MZXJSHU77&
.]7CA)8VO]85D2RCf_39I&4;F-a16:CSWaBQd-1=))OgQ7&F1S+G-#4JS3];R356
F\2^GX2Z<_[PL99EdQ+G6#4K3\G;;YVYHZZM.-)76W(@N<7V_L_L0)N&4aV2cITc
NZAUcH#5[H1,4]dX;OY^_;OW<37,5.Y7c0[OV6CaK3E(JD<Y5&.W<5E/1L<]>83>
,CA;B84)0,F@?:a<EU0b&/[#BO\W_JX;YETPF>Q,=,g&3gD[b>>.2D>P17:5[R=6
e?4:J#c=aRY2EHU4X_FHJ\&C)ge@YX.L7&);c&>Je,J^IJGBTBF@QG&AMK/P06cS
\)J:S;<SV=dZbIJdUY[B,]BTYGB&McF96gO,Z9.Da4R8YMeGU_fb7KJHP7G)@0PU
_J>]IeG>:LDXQ[9AfC@a>aD917:-:VbBHBd>S8AGS5=36Y6=[(9T70A=\gIFV;>M
H.gBYSY/CFAba.bP&bM\Q/;X\->7AI;=#>5^5dXH0M@aa,Y8@2#A9:VTe@JZQ]T7
(4-d8_,MLH]:If)gU,[#8+T6]7_Ag_3?g3F\B6O,HO;QMJ67RKZEWMSH&F1=^#(a
+J;B-Nf\Z^N6HGJTKUPE\e&e>g7D?@cMMC=4YCVR1Y1BNM+0.UU=?3e/XP&JaL14
^eXTa6KNZ=Z12-M^/S(c:Ig64_0+/\\fPT^VYM<_,8e4=5]=bG7&AXE@Ae>#^Oe/
^)ZF0+-.Zg3Z1UWGLV@WG2W<+,&YC3&XF^9G5MGOTAaSA).;c_bCE((]>Ig3/M-:
SW\][;4)>ZX@Zc>4YVS4_QKASgQTK7^F87&O(Q>fF:IX&04BBWFDJ1gfKDPPQ<NG
O0?#(1Y86KWdJ&5;,&8QC.HdA_bC;TDUWTb>Ic[8[=C-/H_<?FD<\,&?GWLWa_R4
D;25IIVSg-U0gcNDV&I&3GZ_.HZ=0GG8E9V?bVEO,+46[UGa5M.L]d);9;ga5:,c
T[2F0Ta5B6FZU=>N6P7Z=X:78]g@W@:88-0311COe?QFNO2CT:dXef-V+(?@S<e6
&J\NPeD\4C61,YBAYF[XBE9^gd8[(416fUaRE=JK:^G?T2BU5\(fB/Q.QeV))D:>
Y]2+><N(B>UNP[(&LJW]Z1TVQC@4?a&D#8CcJMDe0/6Z2/T[ecMc>b\/_A#Ia(4^
Df?=:&O1YT1OND+C2Z+.I+aC<Q::bD?I8<WOII\e^N#>0S6JeA.+SNgK]H[2Lc/4
&TD6Ub/V[._gNS(\+0ZLc-+<N?@#S/9_>,BMP4Z>dAI;K:H[;]F@;2S[.:[)RN_X
W[S@_M\X^&;eaX[MU,N@Jd,:>>CRIX_3+.;gTgA:WIbMgCZ-^.1R+7\G9e+K1#WG
/JOI63c;P^:_M@]d8J=5cWE9,/6].>c7dF5)5WA>g#:B_PK7Gc,?ZY^?)8.;\/TC
I0G__L5107@H,-HC;4T@#8cR+F@U@?8.(7KbS9b\:,6C=f9f;[H7J=C6PIWU/3Sa
-@\;)X>WaW8QZ9.;Pe:NOR?0f(QV[>Y1<PA89>c+]W6;)\D+d.Q9gcL7,WQRU;:N
W]&T<R)(#e0\\[SR>MZ5>:NY^()>]4Rf6C<HH=Sa-_E,3\9AB&?OLVU(\cVfe?1_
f^QC^,dK92X2g)g?D@1CG>UL5:9F_+F,=1b:6H]b-KQ]<(bBFX5/_gSFG?R>fB:f
69S+;+/=.N>P.<A]/Hf:YaR;1G[;M2JEe<cfS,7,/3Y:A]T;-3;eM&E+Ac_-;^J<
&\:2d@JA]DYIWaCAHNB9Abb4:g;<4L2?YX;&4WDP6-0EBcTd&7c/_5Q6]eA7H@+G
^F3V(TYE;<];7;Q0+H4bDJg(R&:[=^fRQ/4)1fUfg2SN,RB+9#fdABUBGJXQU_1d
Df];0bNa01b+c457Y85XVG2=(,+L[>RW5:EE=\MT^9YT50][=^:=R1c1@S98S:b>
24UY^G)gW>QX.>RO?]1E-/3EER(1ag?Y>:eT&b&^]4]Qe_)VMR<F<gd-)LYMH[VI
78>b&R3B@6V3XTbFK;R-B.cEgGND/dGMTTM/VBB6401SAB-V^X=g\FCScb=+?N;R
bf2]9@>0C62eZN[3;Y:RT=e8Zc[E8)MPKU5LP>O)WI(R)cQ[UgPR24-D_7MT:>6?
eS+6/OLa&H]C,Zg&a_X9>eK6<P[@8TJJVK-OR[QSXM/IW<LGf/.H9T9L9/#R6[=A
6XGJN160^?<1YcB^VXHARCe]ZS@QUY:7G<2d.C<36ZeR34Jc[d>8SJR>^/[W9ZDS
Z8FaW4:EXA_ZS\?MP[(M[2c(VbfN9]X@&-?J)c^\],b(:H>#0K\W&#^a-c8R&9Pd
)]^g(NMVAf8FV\&eT90+O^R]#e2Z/a.QcWU@5Wbc(dUgPLGGQ-VR=IB;E,Te+DId
-?G>ag82eV4g[P.E;Y;+_;<UF;)9&<:X-[_6fG7V?+(GEcdHO#3b:3,4?TfYO+S(
Z_<FUE,:2[RNG4GKZR(gT5^_<O897,[BF.DDUQNZ@<;b[CSV<MR^.LeZEfP/#<CW
C^]>4IKA?A(6QGgKR5W6(]c1Se#e#[E<4Y6[\,c7MC8W4I\AM=PKSeYJ<GAL_1>^
A\OWV8DDd#E]4.9GY9.;e6\4AI+VYQ^H)Y6Hg7,E0.C2Te39GZc#d4K>N<DfO>Ze
Y_bOPDV#dGG@43B=9FbI9OD(RUS.Pd=acab_J+EGYT,>5HWb/SK,Y4_:Lf:0g_8b
7]@gD#RT_8=dWaULG3D23[QP@CL&9_M=_Kf+:.b(HQ4E7;?B#Y0?-Q(Z6#H+=[PT
B&Ga;#e@66+cVc<)7-YRfTcQQ6_R;7@&0[c4ECBBB&_]5=[+)CT9=R4F-VM@QB/H
:Z78V?#>d-,@F56Fg]gcYILZN&0WUG;]M#RdSC>S>B_HOD1X-(;,I+8CK<_a662F
10VS8KG;^;AG@1DKSNOW:HCWD;55cMcECY2)WL1f0_A:Ob_DO\1S&L]]ff7K[Vc#
+SRNA]GGfb21_a6?ZZWBRG;LI,DNa#;T+C\>INW?)>KP\E=L>S+1C6dSTADOT>f9
SK]MG6]eRfEf^,@:@11ULPa_R.0K:b9,b-[=E<+BfD)DBC:6b@5A>@LW@/>EI@X-
=cae,F_^KK7NCL-,=M&]gQ6Gg4J/)]c(U1\I=)AJYd8:N,,cUM);VZI1R5ZC>dOE
aT0_I90=6fXWCPdEWd;4K:IdLX-W/JOQ>G5WOK92=\V-VH;PSP/cNaU8_7K[9RB3
#+BRU41/X:\PE-.HBT;Nf4Q-FQ_UAVBDMEc4K,>=U)g7-H75#PDNE/9b&]PcY>V>
MZb#JScg&@-aPY_1G55b(MG5]?a4gZ7d?Vg/;L,FY>71[4eE0D:/(3ffR9ABcFH]
3B/YaTSKe4+.BDUYbK]aQJA^&HTFE(RZcKW4aK^d05=@[fWaAQ8:ZGI070DS(.;O
f4IQ6d45\DLPC5A#UcfXa/0ZRLc2=]bebg.51;X<&1R#;V<N#U>BDG,T@AXQ26.g
H1Z0=cOcY]HLF^1[PVA#GM?Bb2IAd9EfZeL8CY[cU?V[0\87LJE]>\33#7a+)Y:I
eN-N;VEJSf?A;)N=E\#[PP:H04G[?QSDSb/4HDJ?]85V:BaHY,RKTQA-8,Y-e<#^
SB9Y/R(K).CeAc?IGe(/P3>HEX<JR4;T<9>^g(e;#.2XT[c_7-+A&5-<2XL[N29N
B@Q.;K6fFgG8DUTQ0>.^G=4LfI\T]Z=XXRO=84HQBNbJ9:<WbA;GNX,ee(X+P\#+
La^@fe.+gCOOKaG,FC+)Oe2+c>4XT<S#J=aGO[6HJQ/&]9DSM[DI\-;HN#K3N>>e
-3I/bW._ZZ=Ng_R)Z?LK[?[7+KRebX[(DZb[?9S:V>TWJ_YXQ/>f8_Ee2./\b(.Z
Bf^83@Mf(SKOD^N_9W]YZ6L:^KBGQ;8G>XPK\(cO@7OZ66V8=_?7?2L7_)RW2I)(
-HXV-J#I.5@.:NI#UXY4PSfL#KZ65BJB>a>0V.4agIM/^87/2-99O0FT>2WDV<[J
=Ug0BL(+&IXNVR\5(143252K]d.K.\6OGb?V0L7_C)L2Yc3c+&Aeg5TIJ)WWS3N?
f6-5.ESEO0]X;T\2b?:DOf>c]X@43\gJf(=+BZ-?O;&.UcT?CSbeEX-+\e,3^42,
LE2JAeN+3T,IUbOD+1A_eaZ#g5:9=I>UF:Y79^a/VYfU#)d]N5)ceKOUGEE4A>/Q
S8I,>Q4L7&dgU#WE&^TU@03fHD=MF_a_7N&gCR/\]12>1bc?0>RJ>N44L\#JR8UR
<YJNXKKf&89=K@8FYP,OeFSf+2Wee1(Q8/\0S&8VT&>EIcKH_&4H=X#aWJeN9c3e
A->J-K<-&/N^.ZO:[F\cRaB7Ad,:R-O?7N/T0A0<;>.6[-ON6/7-JT8_L(\:K;-+
=H144ZG;6^3O3P1/c_BYYF8<E-gBV+d6W[,A8M9gdNZSJGcgWWfG(C^]^&bV,5:[
XV@gP_a>H1BWWS4)8eHbT<82:&@KEe,9WO8Rc:dTW=[,2VKTHZ6SU4T3GgS1,/He
XS^(VYO+V0ad@H9Y5W7H>RROULb@KU.6UVQ_77HP,G^#)H](AG&^.DL@-T_].@[X
DZ8S;Na,#4NXDedVB3GaYL?R9O^R5+8/^6AS2LR.eXXfY_A0S??5U2Y66PA8-1@Q
=W]@0,@P&@KQWb<QGPPD)0,T9>TFe9A-L6-^ga79</@HXL4WP[)NWNDODa74F8(\
6gJS93K)1SA8RIG<7FHOK7TS,5/&)Q04>M2[@EV;2]FOc.cUMFF@;?Z8\):e?cc=
?Tc_P?<IZS+R\K9V@Gc4Zc9PV=]]3FcC(R]+[GQ2U>#O_(UbUYPc3UbaKS-b_-d7
2caDD9L5_S1-fKMfUc+=21,g8\<>]Y:)U6UeMP^cC3])]g</Bb6Q5(V+L4R])<V_
+I11ae5[,(:W[3NdaZACMG4:1D/5PT,4+1bK\50)KKE(#1CU3:X+B/2L,ReTd#D.
5Q@dKA(:eQUE4:9?F;\)\(?J+#LN^5bP)\@7aO-,ae+AeZ@Z_#F<aX6)d7@:AEXd
7&IK89dOJ,\FJfSKD-W=HB=BK8-6QB6:;IK&>A3]4-SD6_MA+&6H,O:8?6a>](33
,+4LVS>f[3AeCCRTaHaRS2TZ8#g&E6,bVZ&7U)C0\GYfS-),b+G,T=.8D&]=SLCf
ZJ<Z]<4N^>N26U_0PGc&D3A&2<117P8<C8?)9@U#ML>MAb&<P:[A(QO>0BQgd#a/
Q428<f)\XUKBaXJ^DU#6ACLDGf?WF\0E9H&@B3_:1UCX_RdY[2_b(8#2_-Wd<c\S
\ME;XDGE#C=ePTW\,7IXcd(UNBI?[1<)c4[77@P+:5&@S4H<LM2D#=<Le0SXHAX;
fP0Of=3eJ-K.;=Q=UFCYTE<,CD\e[FX_:WTU]<f3N-UfOS<V/]?c:2gBM;^DXGN9
=-+b8I9J6JT2I-W6c^I>]F?QST6UT+fK89VfH2<.R(BJO?KX_22IEfe2)K[3H7:d
PeRLAK.,3UF]DcC(._(OA@U0ZJ48UFI+:@Pa?8]8-.)28BPVSagB;I[14NT7,YMQ
:#P84Vf2(CXN+>&=HE>CMee?U.U70T)AP18DYbI1R)RfJB-V>]5V#g[NPG?7W=Ff
0.P4U]b\[+Td1=f=R;_J28;#.BC,]T,:B8a:T\WJcObD&E^A6NQ>FNDMRKNIRE2B
:?8^N[C;G-fK(daS#QX_ULM,98A\d@MWb)5\RVOf8WeP?B]^f)PU-7EUQfb>STE=
>c=6#@YTFC&Q^TBNKP1&,E2,)-M73&Y0?(45Se>+MEW2#+>-5H;@<f=R4ffH,74:
@^Ja,2_Y<JYcXB&=U([4BZY<75QV[fUBC<W[+P0XU@_P]G)4XXDSG)4A.QL@?eRQ
+EL@>(\6PYA[9N)LB4Z(M1f^8D8G\<Y.-0#37NBY=U?.Z9I\WW/C1#@=d\8A90)c
6,3-_J/Kcf<NDJP0bHQP:H\SXJHHcMd(PL]^0;RX\Z08bZ?D<-S.dff/WN@)g)9>
X+YE3S+2Ibb\2bMeHS8(IEbV&DQ/cJOV1YP2VUJ(A;:_[K?5O)0+YK]/dS-M\R4H
aV;R?Z7dF&(ES(.[1+H;B#X-7;83GP0cKVID/?-D55O36Ca8HUfCB@=#HaXX&NAg
3eeQK:be/[aF0H(>?X(acTcXVVQ(1<8>>=#YAEIee(gHSIMgKNU95^eK,D>G^1_^
V:@(;\f=5f17[IEbRZ@a-@f>YE]T,>D&,GUP_b\EgHfK:GMED(-YTTQ_,b#9.;1F
EG&Cd&/Fg4,A9-I6@ZO/ZI7<d#J\;Ae9LK/;5\E32_d#=;YSOG:KU[70(]c)D_H>
3VF\/fd+XN9@a9[G==4SV[F>b:W7XRcff^6ZRCJegPP7RCI5WfG)<be&g2db0-]P
=4-XVBDY0@:21.&LH&1;#^^K;)<4Q:VF,;d6>^(XE?cfR\PT28Y&(=(W/Q;.21E=
4FCabed0;3CdAW5M^^?Of4@/c@/IS/F1;\L3=:9R-FgY_CUX0#N_EAIfKIfEN/<.
,3:?U2NX3cdP.C(fT4V.O:4/L3\_P_M:]?]O6R@V):#\=)@1gF45ELFWWfL\3O7P
ILQ/ZK/1^g<;KV)_T.>OLb@B9=?S&B#;E][X<,G_U)8P/ZCTIJ+^IL52D&f7bc)]
H^^96O-]Zcc[\WP,fX\ZHI+Tg]D<:c_^a5HV5-KECAa5A46:Z@SXcLC//8496;6(
(E-6LJN>(aaP9EZbV<gK3?8ZUB/&YSEH:?F:Z\Mg8<M)2;]ZQ_B\XL/bV]R/1H\V
N7ERIXQ._>5=&FYD5(ddQEUH,K?0/^M&83J)CNH=/aWg/<&CZ@.@5c1:BJ5-LF+A
^1EcGS6bD#LaM0XQFGPXTc7^KXC0CFg(;RH8O[?bc1;</>D8=[\T/([e)ceL\#XH
U,Q]DEG1Ec:Z@Tb&ZN_MRQ_46;4M9C7+AP<1L4CN+KSK;NL85K\.RFb7<OgSbPG/
eR^Z5I;H\V1:JPc==)(/-3@0K3[\V/f<ZT4+,76G+,V&^CNO+QCI;LO>9IeB^;(+
:22ET67&[f,L6X.@8V1NNO6V->Pfe_H1:92@V7^=fe-R^PK_]1PfMb(=[??cR,7S
\H(bUYBPMF10/4<5JT4g//Y3P<]70B6Y<]&IQ=0\e+e_gEI6eP.\;g5?>ID(C\:=
@-d2V^CA;6(d&a@5?>TP87>PgP[B6cXI3EQ]2<8=<@^f(MCLHF-cB25,Q,ATNK?^
J?XcVGT+3>X\\fc0;1)@=bPO^)YAfH6G]PDabf89\955>d=fN/:M7=^1WLf1UF/^
UGW<L#,O0)ZR:Y[PCI86NL25=7PB&27@2C8+6MZ5QP?I2fS0H\(_+W=W0VPI#=&G
[<N\&#2S=EeE5;b+(M^_L0fa_8Dd-_QG&,+3<^SL<DOY9f;EN/N4,YaX8ZGQFE=>
M6a^1B)E_E4K];SUI7L0:.S-RT2[)E7MLaI(,Ae=?Z?A5-gC\^S5OH324&_A[fV(
=/<:7_N9=R2(39:G/(\Y,)ODF<VK?@/>Y(K-#:(\6\^FSESIR.?BW=_aI^#=X.V-
&^FO^TL:T-HP[W2GLFP)M(E3];J2#)6c6\6)8d#K&L84T-#8IgINLI2-^Y&)]aI/
;)L8ZTd.DAbUPF2d&UK64dOe]_.dZS\3.7CW3D0aB93a#<BSPQ2;ZB4>Y5B6Z:SM
?GEANEP3,e/QeE-HE#BdCR#Je)L\].eL#@1<W<8KD)B7#>+Ba/C2>@KAW5KS\K.^
9MRf-W[,2cY?Sb>4f7G)3=_&E\E^eLSA_GTDM(d;?Vc3SQ85_<2Za]=\X2ba2^+.
ag+T5;S@RQ5gUB7?O?4a>.Cc8(<[5I>W?CDJ,TGYM+E1d<J:@US)=NAK<[F>2P5@
Q#JK(ZHABT?X]:@KF_JZW<7]?\6E-=gMZ?STNW[4?Z82:P,^Oe^;-OJHI\=/29>b
39gaGVTeS:b?;R^JQ[@&L5-TfdJ1,cJYSeL)AN[5P6LP?4FAYa8<ddJ_HfZS\4fC
Z(gGB:b,Uc\0GNgg&FYK09BS:aX\KYAV8)_I=V3(YD8H,)AUT<-1gBAeP/e?I-;+
f/V=f:@C93)3+)X.(,@BW@f]O<T0F2#VD.3-P5ed7g+)U<?cEbR.d7&?dDW/AWeZ
>;#<aJVEDP^+K8cLJeVf+Bbeb>#1RHE^.1EQ]^HDa/MMgHV]M[S)&e>&H]L-JNc@
ZF&JB:7aQ=)A<X5RK-\QRaP_J@&K6:,B5VZ#;5g1>c=N1T:4d^6^+9O#E/gC:FJI
#V?O?GMH/eR(5^?=ZT&fd:NUMN^[UcUV.^];BN=-K\45H&&K(F:W_EJ<7/=P54e2
>:C<P\fRV)9A0F,RF#<aU43W;?F^dd2/KgI6VR;RL:>g,MIV,fY=U_bPdH^AJ7R8
>B=TK2O-M2VI&dfHFG:;dP,C&aHM>37Y#EK/#9PU[FFe24TN+R8)7G[M95L6\1d?
W\ZJ]Y9G4F(43W^&_bHSIXZ5;#6PUJb;]X&/c=]K\dc2N8^VQHNdd2cRE.13O#Z0
?PYg)>7#CG&>3-RPM2\<8ER]B_P[Ua\AGO>H,ET&O(2Eb-^d-^T\1c3T(ge(:XM>
Ng7a7G<1]<0[7RdYFA&\>PL7L9MD9YcSU_VA\QOg/;(8\TY.K2(B\K@-[)aaBc+;
)50M13U0&BKTN,[d?])=;f;L:c(ZPI1b=eEQ,gd5IFW5PKb0VLB=4357PLZ5NPQS
IDSWBLJK7Bbc.ag8:.#5F;N17cK7=/=MQ=4[a2-e190^BdW.Y]4:VCKGZbB,c(./
aGQ+Y+8M7eD+3W/;Wg;:gB4gN0//N(eaH.?;7,^Mf\>MG/&Nd._JQ>cde10[KfKK
RS?J/\@gGM<_.e&g>US>[N+3fJ&0FQ]^+43&^dZ2GGD6_1S&-e0[Bb=;K)^dQ-&[
H#+\MM4NKY>K+U&A5&ZO9CEXd#[K(?>O0Z2KV<\3b3??/EKW6gP80SK^cZIH@T6a
.S0UAfI\=+@D_FM3)E:S#6:Cf&EQ^Z(Xe4>3V(A]#3D]:EgR4IUCB<c=P[/KM-\/
3Y#OLc4OYb^JPCE9;UbbZ=J-G?)\V[?BHTSa\NW<4NMCMgcMdgcX+),d?I_Y)I0^
_D-eBN:I,AgH0+C[:=@4EN&g-(AK=</\E#g4b/d?/HTBLHG:-?@a><^XF_-@EdaY
+3Ed?VZ,PBBN3E]].J+ZKa@f:-U^^OQ66BP37^Z-9A<bLS.8SJBC^+(YX-)63QG^
a/YRQJ,-a.HT(a]1K0/DT;UQK1W4JDI::BK30JGPa7AJUZ1b8dIVS3Pa0K;5UJS)
ERQ7BTOUP8))9cQ&I_Z[.9aZ:H08039A&C=fc/QT9FLCPO[;3<GS<#aLg9aB>CS4
]IgX)12JE7eR(U,A(g1^0Wf,Y=_R6]_UQMCF/,0O6CDM6:0HO3cGNCY&19R=J1f]
cc,6-[dH&dg?Nc0?;8)M4/Z5g(X\<dbZUYL]2DUZ>AWQ3JD6+Qa286<FdWW4G=Y,
.>=ET?-[TSH2.A7#@c<Q7A6@[M@SS<_FMFQ7^a0A^LS_X?=9734::RUN,8bdEede
]XV\5GGWO4OY.d5(59(MHPV9c0U_0(6^FX3WbPO6WZ[XPc])BKcOLMC^fORK@6&E
O0UIZ3@:I[M=Z^PUL<6gU;.Da)NJfH22-@-XbTZ)d,=;3S_&0)C,;?8:UG-[Ma:3
Y]=O&Q<<6X.2;XUX;RT-UO/Y/D7_V,;^)BVJ8bFNRag(dgV/1]3P?L3.0>:>Hf/5
Z\G[OS=_O7]b7@C38]5,MW:5(C>F6gGFH7-)0=\]dO,G3Y/B71fHP)H#2ObD@P]R
.[Ia@YR^8WL?IOQE)fT9a@2b4Q8BQ&OdIIa86I+XGCG?c:0aJR-S;M[WRY3e&K(T
fM#7B6bB4(+faf2_0Rg8[eYU9QfabaT;0UQL0(X/]LJZBf_)P,PW8T(,+/R?HQS(
9ADZ@?7+W_@8#>A;;fC1:RO8gC1M7.#2HP]\YYP4OS_N5UaZ/#2gBGYH6<aH+Gag
NJ5cR=M667]MeI8._R8NU<S1@DF(bYcK\Xc,G@6N[NfBZaCD8bMFM]ARbHg_eYe0
G9R-=/R&\3bEBHSWg6XG-c_>aA4+dS;.R&\VP<9DGW&_7FND@#PM[04S[THJ7&ST
X>VDA/E[7UB^;<eU6V3a9#U<=UR..OM<FRX;a^[W?N?7fML^I?gN9#\c9L1VP?AA
SH+b;2.9&ES8TI;+&UdAXb9gLZH&dYGdQ04:2IPZdL2UON\FV8IR^)\F,Cb).Ad^
T)+e6YMX_JE5D6YJ?+UG8Ya]SZEX2g;<;eK1bS/&4de^YE;FZD:WOMZ)A4fNPY0A
WcEcgTa_3M0@cfVBW[O9aK#=a)Z73E#PL&YfS97UN+53:f;VK\g_8Hc5<V85KZBN
9fUc\6E/MS]GL+9+O98_B9TXM(cK@F8DESXPZENeMdE3^:XLX@EEFG6D(SX;]9Ce
W0@a\PN7VPc\82/9\GDB2WJ>f>6T[TE@BE-eL5-Ra7-_WZL<TY@M-)]0@Y+^0cB;
+PQ(M+SG2_,W[/\dNAY3/0]7d_?XQT9FZGQBR7Xc9)3V)C::XLEFV7]M\;9RcMVQ
(Yac@SXg/EgZ5b:]((GK)THX8,GS(fG,7ad)6Faa?##.PW5,?UF05-IJR)L&2.T/
4?U)-@-QY_fc46PcKdO)Gc,BQBa?2#aeL>+d8+G>F+1NR.NE^0(-H<REL&a\_P+2
L&)HbMd=6S;-Q6&/[e,9,79e>,9:GR4&</4U>#E26e;)Y;/H,SBN=?->5#PUN+[G
C;;(D]??69\.&W24AKH&7R>-e];@:+[]6N9I+_:I3&M-aI:-)>T/AIPV5)ARQ3WT
R9U7CT-5?:a62-ZaJ39;c,;K;>bWKZ+AZ2VB=&>CK\\_(&ag,dG^O#,U18HR.9ZH
RJU^2,9(]^^_KNGLOSXP]X;.N9[AZgPF;03QA<&bTgde&@?<-GF[)/DOcKaS\690
T6/O#@3G/TGLWT)#L,&DJ2L&DV:I>6[9Q&RbZA9H[aAg9NfadSHE^NW8A-XL1e[3
]OX26=J8d#/0@57+L?OW&Y_d+2IT+M5O0;_^@L(&3?>\@Z^X=O#2?6e_3<:A.W>3
d+Ma3#dWFCZ&&G]B#0Egb17dB9Mc<^GC_/^,YD.+_KBQCL]?)Na?I0[_e(W^TPf+
aZ1#Q9IHT-LEOXQ139A6?+=ET\X(cQg>+S0(R:V&L+],1-.GQXUg6MVX7M_P,)O7
+<7IHgWKSQ.Yd<g+dc7=9HA4@]/cFB9NN(cPO7T]<c,>.(FAIdV+(IG1BIV:f6U6
-+5RZc\A20+-M)FB,FW?H7IgY8LCQTYaH8:/TD<>M_I;)5=9XQA.N[PPU],B#-[6
JQf/fY(#I_YJ0fA2M,b?32<CXBM[S]1<.Ra0g:;6@WA?]C>URe<5#N7>9H<T6>cc
0Z-bd24e[6ZV51,Pf&)g4-.9JGbN]I3MPIFG_fWV7.[GWYK.d-_8KF5TcBB?V/:L
]a@aIXQ+/a^>E6acZK2O(AHRVNfe<.V?B<cd<UcQOU];9ae.BA1RMQad,ARY+7]/
XN.J3#=#3G;P_B7Q@_YJKIYKXQK7TI98]]bJI9^)TA[dN&/NM-aEFV^P4PB0+AEG
;#0I+g.1X1CU3<XE,6C_2Ca27_5b>5gc6[SbFcD3U8,Y+B?:?9(B2DU[(:+:7LF]
W(<36KA&XQ-J(QJ7XU[&CAV8.PGX0c<RCf5C@,.C-U>DIIRPD?3OdK3\<FMY=.YD
@.B0M]Ca)D,I(U3#VWB:^;6=M:U)?d72Qe_T]cfFRCWX7]APabXA(B&c+Nb,eFNJ
RbQ>1WL_A2RU4g2(UKW]PfedX4(\3/L:UI/2#(JM#(^QHSf0f&2Z^FZ(dd->6cFc
-TeZTgf_&631cL6GA;?M>U&6L=f,a8J]??2#)UH1JUN>&.a?8?4[=X9AFF/-&Vb9
ROUMf\F:K,aN>4SHD\(E@9Og869X4>7915PEbU#]\A.-^T6G3a-\#CQ/L=)8Z6&U
,b-IEQReWf-/1E^,TB@6Y]C4/_f9=[#W1YS&J3+&dX7aMe+I\dKH(eZUQV]C;A0b
FT1U+7U#X+7K[a,dJ@,B#3EFH/d&NU53a,<Q=WP&E-8U#RM1(FdS#a3K<.Y,UI[=
YZ.aH\T(R=+SSR5IY:g:;_AYc@0ZJ7DU(JM5L4a#(H9IMQL]LQ:(#:5eV:XI@Z/Z
c=dHW/1b>gIdO&-IdQ\dJNTM(e6XMfKYM-cE]CEB=NRC=>;:AS3Dc6PWZL6RE23F
@:E1<G2AW_8b+#QWZK_)g@KUfMDf,(@^2F-7[^6bDHcA,ZEDPb@V5]C4P16@d^XT
91O<b<+R5b8#+G7a\0W=O95D50+I;Q2MR4M09M\_85#O1eCdRNcN@2(Ycd,J.N?<
g=b/.G8SWFD(5==2:>bF09O5A:dSMd2PCM=NfY;X8>cOcQXKQ;#E/bO)T-@Y,LX7
)E4Ua<3aI6a(Z@L2gZ>9+R;^(QTRW^,1=78NYJ<-O=QEYfIAgG>;XZQf/(>;--GW
EM)VO(8272+\d\V-(dQWL2#2;M;CSTAbC^8,ET</dU^&b[NN^>P#:B^-]=A.VO?H
09TdV,M^YWS:OJV-_HVQU_2,f=\4bV5QAXe;/8Ge(+f3XJb(OX@>+;_M331YXI+f
FRO]Q++H?4&L?40AUQ9a\JbV63#gK>P2LML8LU?@L]#);;Hab&784^9+?IZHS6AD
)4cDC@S23[YF/R\;.R__AM1ceT1,7T=-_-5QU\)#DM6bBCF3=-1JYC744E,]/=><
R#[7T1IX:L-F[XZ-4Y[0a&W_<>d=\H0Y+Z(G^R<>G(cGR;d?<Wf3=b0XLE.9.DM#
LRA_HN6HS,A?Y]0A6[L(/b4.GH=&RWcO0fAYR-W0fYTfeM<7>/@FNE4\\)(_Gf7U
#e^cc\Ka^8Z@3C9<P8ScQbbKc:W-D&9BfQa/+7+M(^R7?_2#JT1d8^3C)Vd0f4@Z
<C41AF(^^ICFVJ&C,fKgEA.#3>d&6?0:^F8>e1S+<?7OC(//U41/N0QEHeI_0JWT
6f1>eV@8.c5H[1I4#DaC(V\e#)OLc:5I5[<\L9<<H?Md[2SMeW494KLP/^45=a?3
6^9M@1</R,0X&ff.4&/B[KU@X7I6_>?GY\[2O+@OFAYNXZ]bM.O2#[8;P+RbR&@E
,N[>?MEMUNA+N_P478>&8R2g)A2H7ga)c?_bF?>OBJH7W5ZDFKX?9L>OCb7&3,16
E]^^>DTO31HE3K-Rf_[f#G[f2U\]\Ga>bY]N33c\3?GM6VSfdYXNBORgU5.5_V,)
VQ#4B\U?/.>P6\X:U-V5U,BA.SO5YB\\5J^AKQ5f=f[Z<d_N7Ea2IXPUaf12H&/>
FId<J8);NPVTHR\+\C>cGf3RNW2/T-[@S01+>#/JX7(O8D/[g<Pe[NCHY-a;-d98
[V3_?R):E)2QWK6#-@Y.9O@T>)8#\XIKGOE(9#^&:EX/H:N[PLBPAE7V9(GU]aP?
ccOA&F,S24RBP#.cKd2DD3ITR(3Q32K^,ATB]#]1+8CB^02]6/+(N,J3DHd-\C]6
)C8O=ICXb+P_bPJ<#H-<TWP^CJ.)SC8TIcG[Q2K</7&\FNg@S1FR[8#@+=\LH=G<
VCUeb65)BQ>&1b:+>V^H<&KT>4@Ud/dIL3f-ZX7XGaRIFgQ00DLNTbXEcTVV;aN4
D5/N_<7Q^DG-EY;G<O)S1UQ<,GG\_,0Y1f=2R_,17bZ//dgfJKB<8MD:IbC8g][]
IePYMd,RCB5gMT\.+KTg<[e8Q\&g&:EF@K?/QPIe4XOf(D(VDR_^LT_3S-)4g-.d
QXd-&]\7R(:D,9A,SC-X;QXJJfP0EJX0VVK3RU:2LM(GV@NRMQ<=N8JF[f(N5Ua&
XYOJR/M:bPGb0RB.e5CaDOLd9Mf8Cb/N0KMJDPScN)OH96V3TIC+=Q22G6[Og4GQ
C3-N#YebNg_X\=:SWA_a2.V#2b(07G<S-6H4ZD&-^9AHA$
`endprotected

`endif
       
