
`ifndef GUARD_SVT_AHB_MASTER_PASSIVE_COMMON_SV
`define GUARD_SVT_AHB_MASTER_PASSIVE_COMMON_SV

/** @cond PRIVATE */
class svt_ahb_master_passive_common#(type MONITOR_MP = virtual svt_ahb_master_if.svt_ahb_monitor_modport,
                                     type DEBUG_MP = virtual svt_ahb_master_if.svt_ahb_debug_modport)
  extends svt_ahb_master_common#(MONITOR_MP, DEBUG_MP);

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Tracking number for address phase transactions */
  local int addr_phase_xact_num = 0;

  /** Tracking number for data phase transactions */
  local int data_phase_xact_num = 0;

  /** Track the previous HLOCK value */
  local bit last_hlock;
  
  /** To track if the hunalign value is changed in middle of a transfer */
  local bit initial_hunalign_value;
  
  /** This flag is used to disable the EBT due to loss of grant check
   under the genuine conditions of the grant getting changed to 
   other master after the bus samples penultimate beat address. */
  local bit   bypass_ebt_check_flag;
  
  /** This flag is used to indicate that EBT occured during address phase */
  local bit   ebt_address_phase_flag;
  
  /** This flag is used to indicate that EBT occured during data phase */
  local bit   ebt_data_phase_flag;
  
  /** This flag is set once the data for the beat for which the EBT occured
   * is fetched */
  local bit   updated_data_for_ebt;
  
  /** This flag is set when complete transaction method is called for the
   * original transaction for which EBT occured */
  local bit   triggered_complete_transaction_for_ebt_xact;

  /** Track whether write data got sampled for current_data_beat_num */
  local bit is_wdata_sampled[];

  /** This member is used to track if htrans is driven to SEQ for current_data_beat_num. */
  local bit updated_htrans_to_seq[];

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new passive common instance
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param monitor transactor instance
   */
  extern function new (svt_ahb_master_configuration cfg, svt_ahb_master_monitor monitor);
`else
  /**
   * CONSTRUCTOR: Create a new passive common instance
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (svt_ahb_master_configuration cfg, `SVT_XVM(report_object) reporter);
`endif
 
  // ---------------------------------------------------------------------------
  /** Initializes signals to default values */
  extern virtual task initialize_signals();

  // ---------------------------------------------------------------------------
  /** Update flags and drive initial signal values when reset is detected */
  extern virtual task update_on_reset();

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the address phase signals */
  extern virtual task sample_passive();

  /**
   * Creates a new transaction and updates with information from the first cycle of the
   * address phase.
   */
  extern virtual function void start_addr_phase();

  /** Terminates the current address phase in preparation for a new transaction */
  extern virtual function void end_addr_phase();

  /** Moves the current address phase transaction to the data phase. */
  extern virtual function void start_data_phase();

  /**
   * Terminates the current data phase in preparation for a new transaction
   * 
   * This method is a task because is calls complete_transaction() which is a task.  The
   * implementation of complete_transaction() is a task in the svt_ahb_master_common, but
   * it doesn't consume time.
   */
  extern virtual task end_data_phase();

  /** Abort the transaction for which the ERROR response is for. */
  extern virtual task process_error_response();
  
  /** Update the trace arrays for SPLIT response. */
  extern virtual task process_split_response();
  
  /** Update the trace arrays for RETRY response. */
  extern virtual task process_retry_response();
  
  /** Update the trace arrays for EBT conditions due to loss of grant. */
  extern virtual task process_ebt_due_to_loss_of_grant();

  /** 
   * Abort any transaction currently in progress. The argument indicates whether this method 
   * should wait for reset de-assertion or not 
   */
  extern virtual task process_reset(bit wait_for_reset_deassertion = 1);

  /**
   * Utility which can be used to determine if the common file is used in a passive
   * context.
   */
  extern virtual function bit is_passive_mode();

  /** handling of rebuild_tracking_xact on active reset: called from update_on_reset() */
  extern virtual task complete_rebuild_track_xact_on_active_reset();
endclass
/** @endcond */
//----------------------------------------------------------------------------

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
qsJGtaEqMXEg4eNYu5EXlHAIrokT5CmE5KY0EdWkrtEUzNF4hfT/KwTKJCMAF326
ES0OnMV2DPmqaswWJY8oDKyQ99NOr5T6Q393peOSS/EMJUE1OWmYwbb+XTeTYh/5
2WF9VKst87KyRlzggnGebjBxdWidUNvLYb94WfOMNIuaBV52FZlyWQ==
//pragma protect end_key_block
//pragma protect digest_block
kGVWvRKuIUt6gw6BIOJjwCn+7I8=
//pragma protect end_digest_block
//pragma protect data_block
2wx0U0kRCMkxQl0AJIPtNEO4JYDkNl04YW7bfe1+QWIsHSOAX+SvYlxF+BauXFxa
TRFP6ZanHSeUWw4qRWOp6efFyqtMtXktLKcDMEG5ZL5WgFkP6AimdSDdBTNnEX8U
4Wuwdrn95HVE6lO5z58flIepsIIV0EEHF1ffue/BPlcUGO9vod1N7AZitDROmUR1
b7GliMXIF3cq+je0cnicF6KmDE4B7Od1zc+QiRaLwfHhGaxvhJZ6B6nMTd+QMBkh
sNMw7mLplMgNuR+fnWF5VlE8gNbRktJzHEVrR8p65QI5JiQohXRVmqvQTVKOJ5ea
91MFKY2jzAocngyS4Eb2uC8bPmJR6NO/FVtGN/2NO5mYC6X4HdIHLs7/9jEisfzp
PiF44Un+ZDiUdCPh6bNnGKVB9gfsa3NIH5zHn/auBJQ5THN1C7seVEw79S66IkMQ
j8ZI+NB6QtshVykZLKxYUwFriwD8c1xznjJPTR2gQ3O3kMfkIouxr/Y2IMvKFGsm
RWaXtdKyJWCT4lXQVEcOnXRjS0KJA55khozUaU+AVKDlpyylAmWvVsHbJGYGPCUk
NpzsQ0APQIijCMtpHzqPvL8VwV/bTW7TWEJWj+JkMV8sKgzTew86TyUz77op9O8L
wUY/RDb0IgyRHoID4N6LTURiEUp5nTaGNjMrX7PkEn7ywIIsHMHiZN2R1udTJhJ1
u+sIjcwpYRzmexxFkwO6QNBzqpr/elOCpLM+5Z6ZYYwd5Kzses6BxWoUGIIRMgqi
UV9+880EN9/8NY9INsoNZUYHoh1Wd5Owr7L/O1msKQk=
//pragma protect end_data_block
//pragma protect digest_block
xlVb3Yd3kW2Ak6krqko2JLLnric=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3ZZGZ39LM1Gg6i3/cK6W/qAtQB8KrbSWKRtOh+wBVgCu2MnmJrAVG9KtISONBgv/
ks41B/MJbI2adi6lJby7D4eCBE1Tvyw3MlxPnrlHDEG6BJlyb1gCdds4/vhhcDJ4
oI6dd8Xh1hYW26XDVzGfPd5qoi3NGjaNVMUMFol0X5SkdfdWu1djkQ==
//pragma protect end_key_block
//pragma protect digest_block
Bz5iqkwlOwtr3ZZB1mutyEUnH70=
//pragma protect end_digest_block
//pragma protect data_block
vXkg0vedieqeu4NCx7NtL7GNm1QPBz8ZlaLOUBvjO+MTvhcM20D6gfjXd/5IgG60
6zG/MFDvIGXKietfzVC/mdQ5wAsrNy819HCKwfCHEDn/yoDwqCPmilYalUfY51Um
YgVPEmhty0Tu0gYDWoJlLzEC+xATOUzXFij5YVMqKGMFH6MX80yVGW1d8Hru0Qs6
QT2NkP5MggPQqmff1h0/klWNUUaKYknLMq9WCW8mTkB86J0k5v9RqVNXJHFZ7j0Q
4icV0U3aCsZrvqNMgKJum/GtjoRC7uImLmHZo7//EuUTxtltalYx1ir6g8Pnma8w
aTlLdKqGZyBEdvvTHqbaZbSXWQuzkxtjIylptU7pmvmyRXH6M/cSmqWED5KQtjYj
lJDnygscSDTqtT9HLcnfTSALA0HHNGfZxy0uP4RRv7zlUGLuU1OYHWrH7K3Vhylh
k9x5zVbHGlo2OAzwKITTIgFbBzVbeaLK7RgQW707HktJkcN1QNlqaOKMI8bi+i3D
/2LhmahCTz88+aieMzTqpummp/CmUWvzhl5o0+6PRyr449yAWaUqoG/dpXsaAdP4
AfTBwHWsb74TTJg/1ese+6CysCv/a44K7IoKB4z7MJeqnl1Gt1soHhJ5gKp24pwq
L7vH0ePAN8fA7Nv4XJsaT2ElzsqKXwD5gaKm9TaC8HrV0FWGVfcbdF2RacZiJ0dw
SO1FRVasP5/NdGVPvczcTLQR3qQb+i+4UIzXUkjHcTxztlQ/M5ODqHm+iufH9zir
84bUQ3qk5KHqd5G0FQ6SdKz0FFjsxFNlljLAnusAsNMQSSLdvG81lknp12gB6SoB
A3+awdClA34lUUkIza2JasnQEFGqGa4L0dXYlGw4fbw2K3mB18zfwwiDQtOOrlB9
gLnHhbuLLWzT7jnhm90yNHLSOgz/fcDri0bK1illXx118eKkEd1vKMcyPzlkJi0u
2SdXqJAGfm/C0BczHfhnLkv3HFgIMJTLtcecdtSOP+Ne0SMIZ4qjnWlTzRnoA+Eg
FoTr3Ev5W3gM9jBHgHTwqbqpcskuL/yIIaMoizbMz7sSNLvdK0pfk1pm5kjQiJ7H
lo+MAYqq9/VoD4lGkU3LB/j6kGhUvgMgUnK+Pt40+MIikUXO1Ll2H5Q7JjEVqkVt
RfgFSK8uokjkWtLbI+U8nUx8Z+/VhwCSSrVO95BJAgTby/ZGZ4e9Eowh4hTnhV9k
XDbKLZaA1kbEmqiqcRTLCzhu5jftEhupK9D41Kf9CtkUzkEBr9ImRAlYKRj2DeSg
xSWb7Jn3S7Lo7QwYJbIpmUftHd7oRj82QkkrrGz2HUOe+9oPLq21SvZ/pRt+Y4P5
pEI74J78XSFog4+H8kbatRM4TgLmob/2x7le+oj0w6J0+PHIFt6l18/2lMV9otk7
kLQxJhXrI6pZOrIesEcms1OFnPfdDzVXdksmDIhBxfIk1hsGMiY2WqyiIby8A9gN
1/egnsmBDUkTxqIiPKxc4CE07sflpNRSw1wwCQUf7bkgfvmMhjCdsg/sy16Zwa1u
Ztqphe2eaGGSqdHYYMF0Ti6S/47np8skmwjJCnM3Wifq8JyLvURN4ga1TU4qkVUh
4zwNgHNla5F7Ju4vJzFzswjXxajv/hUOf4uwUBfkKnOMr6ZlhcW7MgJ95R6JYGTS
jzMU9QP17oPAP2FmFAbEVvJ2SDbXsFB+lg7ivdFK89esxZ6OGsXhCUrB0tV+VzUi
JwnWtc7hyn1DyoB9pEizg43Jexvy/ZCKqTlF16DfOqWzkoVAN74An15KhlmzphhP
Zvbgan5HI8Hv3rjZwC6e7O9J10wzmdqyiA63xDaV15f2Eq4sAt35U+mXtpp61uQn
27WEqUpPE2whjGdyCrDV+pyK/rzSRPCu/0Bh9bNwN6TWZyh4dTqTlOFtrUZUDxcr
Hehwv6dhFbTjtGx4Gmc9Yw+J7+01HIHf7U+ECF7RjVuvwskBrANeKhzyOPFynCTT
rG87ksImO0ElrbvUW5M73bj1cKvIbXAT29JlrzJ15FbM7CySXmpJ9By6MsXlwv5f
YRRwE6t+WvOVG6jRYB8a5RwiYbrTiaIwoPsY0TVFRO+5mTI9NMjaAW5PP4kD1KXI
jcVLWzVtnclN9vP2hn9gUSMWOdMAeWWhkwAxFfcivwZvLiJyAEQSVDaaBUePg6DN
Bto0FIZEpa3c/dxiqIthvNDmCtZEKUYJXBdkCtt76KThCSloo46Uv216BqDDAweC
w31HngbnfIwaM/c1mQ+tAtViuluLf9IF3kTQE+da62iag/Tip0WxAi9BNuiSWaPb
ZUiybPZ2XvKJ0sRnisdZFPrMWlVC0EeHbbV8H+jmPu1vLf6fHJy9EZiu98d8tUMh
2q4ApUEiTGW3S88h/IP3IuhimrbRFDtYx0xmsFl7TESka11fIE1zZSAKH5RBxU6c
WZBUhKoVzoD9XVV/ZkrYW5HOtvhN2J7rC5AuUiH0oiIRhjA8vF063ww3y3dDQMxw
E2pQItNQ+0oJMcbsmqZmJr3D/LAt8NfRDkQqP//JniI5IP8YDonWh0yKIwwWLEqY
bbVSKCAJKNOJ/tsRgyn2CyWmWo2WcG93+0toMR2PqUWFtqyGenU31bGoNMj7utH5
HjiyoxChisAkm6A2HWxJCcSFm3gGX/BI+2ZLcIcNQJzjIROeOofo2nC4NV8xgxoh
yfn5yUk7eUr8NYt0nhWqSRb6fF+JeTLxFpfNCqJ4P+Mxc3JLcuFHB5TaYwoV7Or6
bFBjrN07qP59NqVAvwOPQHr+AY2dpHANYnL59BHp+nosjwDURZCG5JIib/PbDUYi
nV3CthlL04tMTaXa1HO9kIh0WYAi2RVdChp1IBhVZ5KRmD2YfVb+YJgz+NHAli6t
fy6Os6D40tF1w2fayifThdhq2MzdioWOLwXxmU1Hvi3oWMU7xAKX/ywQVvF47woP
/BFwbVm4y+HzAui7R3RG/6WJTGEK9ROT1yYOsY0bxWmREA6lAydF6M4vDMtZs+6f
vdsGS0E/48zrba0rScAihHTR2geAtTIHXhlYbAd9Hvd2K7x6YfHk5i4HwLtOpBUd
G5ovMxMmxYi3nISlab/naKPysGkNxX01dByi4fzbAN2eWiJB48WJvh1YfTA8fsmF
avB9P5yh1Ily4oC3tMuT+HH+8VLDvLIhpmYMKjc8d974alXOpfE2eJY7/Zgfn0ls
ihiMHDAUja6Kf1/bv2xDRAyRoXpVj7p9m/5mrwDN0RgzjnK+MTZOtksubv3NHCrJ
NXwNPmcvJviGY4EgT8QqU1gj4XlFIGljL1cDDRUHSV4rZQS+Ds+I7YFx9rt2owi6
C7Q8xExqZVSCPOD5CwjPw/T8PqWVHT5N13NVcxJyRSOQRYj3ekUpkjf3S7F/eH9T
zTOD/XSVxUaatQTtpC4ex4BldcDHo13fqTMqf/D44iPEhPemrGNmY/ujs15nxfgB
j7au5bBcQ4iKIC5Wp1fI6qR8MPK6wuLrZ3939FFb2pHBAH4tQuvsN1geFPgs3tLn
8zdLVTYi5b3tQS586xqMBDjomnqSPPWVnxFMhEDYG1i/88AIPW/5oGC0EzDCeNpw
VjtvfWx8nKRrQVd/Ap2tdCIV6XfVfz8oASYeNSVxF1THd5wLgBIJ+jT+ILey6DlC
Bwu6uIznER0CarxHkCvceiAobC3yztuZCUnJ95J141LLDOgFFxgFEX4IKBGJ7dBV
ArirQ4tfbBOZoh1v1vR7nDayZXRyKxw+6BDyvAxRMBA0cRiXeplQ/7FH+X7WowLw
5ZGBYU60Pa9qcIHby3jkiRnd9DKSl0gj8QgfsPvMPksDZzYqaQDZZeOx8rTLDi3u
38Q80tv2O1NVeXzBwIvwglIJ4xivhDEqlA/hSaORkzsNZeTtiYpvebaaQWtyGIp0
cFjq7JaL7EZTbuqH4XsHl7E/2wPUCMxaDpjiVPIcMxZ6J+kHE0R6KtgV0c9hlVqs
sqRAJv7cwu4OKMy3hhdN1g2O8As2KTNVOjZpU9eRvkhhun4WjkMUFFhz6RjgHWD6
wHzD/ybXM/j0UXMgIZ6Q8YLkwxubXm0GxEQyzG9pD6EfisQ+rLr88+c65yP92gRH
5HZq4BmNpdbMqTDBIar/mdSbS9yHPC2a86O+Zr4lfa6YYDMSjFas6cXFi+DaqEWq
doUme8Rkw7+/ZIIE6/VYZwexPJUr+tUIUgZraChc2yDL2QBQc4jPDvPUEWWStcmf
KlrwyE2SK6D0HUwK3picH23yZC1i03RjLuODzd/XqbZ17FjZlySiiZW97NQzY9Fm
j4Jm2HmNrmWleGF+hXGJXh5E5k0RRylFi3k/K8P2pz2egrjkjw0NU1f8Rn7Izfjl
zQbiQanS7LqNbn/RoDlS9D4nLxZQb851MH06mqWmh5zRUZWjXC14KIgELujqjNHR
ClTnNoJKfL/8eT8F5PrN0RVe4twsFUn3iwOL1YAix+g+9fZdQRemtBxh1vQZQQyg
KlHgSlWtUXNH0JPEjY9yQa7ZV9YkD7Af0trTQsAYf6fSCBOKpd0EGSEIWSCS8CGF
o0QshAwidPeTw3g789NlXkEoyqgaZ67gMZdsagrfPTkNltMLzWPNTLSOUbX15Qgx
A/0cvWlQGs2eAy57Mh6WafahcHMwWyoB+xgpEt7MM1ffcozyiQJsGAorYIR2Efr+
WW5NtxJwZ6cF3Mdw7pyjSBiixM0sriUzZ/qymskm6biqW5EZMnPMz08qtYgLxr7v
d4dBnRPlaRv+EYSveB6qfcagPDa+7MPw+M5od1X/U6He4GEk0DGNQo7jh/i5L6rk
a4I5d9eJyGYLGPZrm2QgJTS5VQiNk2tMAp6db55SeVp/4zdTmKXM14cabVsOu4gr
kFJyovfu+XhwKtVHDalSqjZgrNSxmbzC0tvxCrESGboGwPYZz5gbO/oBeqD9XM+Y
o5YyDOfsNGge7QzI+qIXWHSNwWbcf6/NjlmD5s6lHzxfEk7a8AQlXdrkzIhWIPv7

//pragma protect end_data_block
//pragma protect digest_block
8QvFuBKEh14npNFk56jKzMVox8k=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
IRNwy/cL0+sKCjb+NB92vExZ97ZC9Hrl+V1vQ0fH91ay8nu01tC2YasMVmVXWQ75
pPcLQbAVuffP4tcRHlm7HfQlvUubeMy7Fg2eV9Sf3dTY1f5WKaX/h2TAa9KvlJsm
dYs+ZBETjiRCv7P9b5steVTHssJaDJEjObaNR+5Qj3QfoJXuX2C0LA==
//pragma protect end_key_block
//pragma protect digest_block
tlo4kWkZLOSvoFuZLCnVWXAZbOE=
//pragma protect end_digest_block
//pragma protect data_block
QDP1sd05vcUeoR59GN9pMK4OgYbcuuThUJt19sE7dnb/wPMOZ1PZ7KLFMO2dIclu
QU51gF5pfwokxZ0sU0J7J3iBVvHjNLQF9P454INNnC4QJtNUUBo5Cvb15cC7mn2R
ZjkhxC7WaXdMMxaSq8/YVPWJ3tzHuNIXnPiCUEVPb9alp/aHQHyOZZo52YMlvVRB
krsHV0sxasGd2YDFceUVKSp1AXQO7FmImusmIEjKf/HJ5Pu+i5pgryR8S/Jw9VKD
iZP0hLrfVcqrHHUwt+MuHqlac6BilYeB98WOssxn+lwjYQHklMusUWi47bUP4FIl
1/74f7Ny4C+xbPfdHtxqRncRNuTMVWC83Nux54aikx2X9+1SB+99vCS30JfA04uA
hWWmuaUyXOQaYXVYMuq3BQNyIDGpg4AnC8OydMoGp/+PVC4nsDK9fPMnNesjxky4
N6Oe+SdwuVV0Z8CH+/9L2+gfj30pYyGHDf1Qrz2IJ14Zv5FLM7JJ94WqP4sxgf7k
Ob6GHDdJUVJg3VjAGIwFTRc1tPjfM5q8MO3RUJlRSi+7ohM+MZwztPbsJyCqnrax
MAHxZOG6W0pNp/GmIUQV0rxW2ZvpjBXo+xPSNIubwzc=
//pragma protect end_data_block
//pragma protect digest_block
toQKq8s6nqvuSZlxVtvFkyjI5Ng=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
1zFx+guma1rjwq9pWIln2n3nTxWBmHBvvJHl+i5q4T7zfGbZjyCCd0xnbVteBGoL
urAJP6M9RG73tp3ziJP3S9eFvS/t70tFcgwk77aum3uCcb/kSqgDlgq3PxQTXLCv
VDNiTJT1NNFqK18U57pJHCcvtSYMfUH0ZQ9X738SNyJUDvak8UhQww==
//pragma protect end_key_block
//pragma protect digest_block
+ymVj/USrajRk+YsFrum8fO+Lfo=
//pragma protect end_digest_block
//pragma protect data_block
NS2Ko1GJJpXNb/QtMo2Rrir+DIMB1GCeydcskIEGz7kxo6XNPl40dwkQURv7F58v
Zq2UesNgyI3Z8Kr1ghg/vLX4M+B+Z0AXh6kh36CVFOWsRxfnVvW+IDibMlaevECP
4PFjyH4yzbIFw4RfvlkI8Sl18B3yZAt+VFL0TkSX2LCZb7uUs6doy9vPBX+DguOz
CLgxB9RhjWztD83t3eY8/T7V/m+t7yJL+Vol7QO+SbJiY77grr4RYR5dVNii3bb9
npouTVZsL62g8yMn0mKJwvtZSUl/u9OUSUmVZqg/kfCAuX9Rajf4amWoAkOuelMm
clBGhwswU7JZUCFzTXqMB6cUGBqYjxjLV4SwCaBeqBAglQzcBwMcVIDDH1eI+WUs
TEJy3fi7BmqXHY4MGwRaDdCb5qYQHlu5/BRNnctfyPv9n82i3aZjmm/g2ARqcZl2
bfBNezeU+ifHPBQfOhJrgk4ICPFDRaMciC2EO3KKKys+wZDptvTwS9zUwk9+KfQB
i0YDaPVlZHmiFRMTueHue4uZXMpFFOj/fZ0q00fAgmgMxkix1Eq7Udxd1iiUfVVY
atqzxSvAZxHUuxkO5JDWH1dgfWPZOKniJE+Kr4PDBUvvKXg1eCQQ8Tx30JGscXLX
REaeg55DNfyk35SiyP8ufj7tNbL91R8X8slYIdKtQCY1H92j8CGJ4rbJrDfLJN40
vYuWl/Xjhr6iytkKeqQ+T0sWaKLrna8PM2Jot0BmP9JBK4ca1g6PSxFNV/y6jhgg
2Mub6mgdeoS33FLKernCGaOchjDNvobmS67Rrlv448zVzDMjQraCBCJsIycctT8i
P5v1BE+S3ml4vOGlCpxhT9sm06jtdN2E5izz9ZrZkzLM47e3Z2trmRnHTAkpmSL7
EF/8CJGt62JEq6+mOLybVwfsi8vlmrumVAWfy5h5kb/ZGIJwYfDKCzmZphl29KFh
xoAJ3NiMlIexQShcI7zTo3O+vBfCCScnswN/8AjcRnpalQ/4kyocQGV1ltr/7tzP
LAWSKUar4umyiSUIVa+Z2+Kc67fqrxF9ZvTTPIj4xsyyrAWnlzxAmx1JPs0I3+GC
RseEfiArly6r3ebg5Fcst8kqV5nCC0+0+wdqLJwtFc77zGw1Eg0iKI2RLUFTX+ce
CmChRqHRu0ITq4RxbzD3QMShZLjOL8s76PuIvvvqYQfGpMqci2oG4c8XMRjd+6Za
LbZ711nqXoMMabrDnXt6i/1NPbb7//rbtlQ2HiwxL8rpYCARh1Ib2tSJQDJvOegz
Z9S1vaPEG7o8aYTt97MNeBTM2Kcmsu9hJdokdxnldWCYQfM9dBXB+XBXxQkvpiGF
3Y4DxLSmPhOcrPxOOhvn+vo8VFX8G5bj6b64tK3UtJDfi/LYRPqBXLIqV/50CL9u
YJ66ZrsnI8b1dl7QuJyMn83YVhzlHgXobT4B3CHZIvle3u+evS923xl4jX4we/NO
p2u+TtgzwwsNh2QXXY81MHhxtO3RCPLM3meqLpOMofy9F8oeurNBHT6sNqQdVXAK
viEcJdDJbbiyl1jg3pGNiOlm9y+Smxbb/nY3aDOv0DFr9gKgo/6QbzoY8ZAl8Zrb
o+3SSSCmT9qKvxwBGS+LkNDKPfO//zNF5o2ZsXglnv5VifH87bAbB2M18+pmnXH4
Vi+TNTFljoJAF3VQfulGnkOtZoi5Qoh7ZkexoJr+IPR3uk5hPIOx1ZQ5owyjE9SV
1y5YFr/FSUThgHyxpK7kT4UAViLjYvH1WCJTDKVOaL6psDPy1xhG2wc6ko7kIW6/
hMIu1hkzMAfclzyL2LPF4C+1mKuVDMHdoEEN7JaKwaLOFf0egw4EsTLnPbyv/9IR
y/qhsU4wB3IiJGbTjPoslP1ICjrgUlidN4TwZizhvz+vVLu6PLjAwdmpQqOt1t5m
/nFZReNNpesHSvig0mFsaF3VmnQQ8uW/5z2n1MyNJ4CMfyoqI9cSLpbceSba8l+2
VWDxcrkI5lZzQoYdYVFDNGQc6bvvnbxfPDB5sobHCPkBYlQT9p7RMsawnK6E3RmB
walhVnH3YEeJgD2e6Bn+yiJFikYdbOisufXapYZAGCYuZl3dqWJyazDO2phUvZU3
/EszwOguhFe9ZsD50IgS9+jF0Nb3RxvHjLtOEJmO+Z1wRAhwZEzhxcEcK61JMlm7
JWMXaBvJEllf5pbC71Iyz+KVP/IArE2UnHFqIMmxMeADl6UI5Y8xn1+dJ+OdFBaZ
Do26m5eTTBPAnLDTLLnzzFwl/d62B67rZAqAPweGYsTVwH2lOBZ39p8lEEB+dwUy
TRyXl5GOVZl2GsJxLef1PJygMC28lEGqRTEg6gbwj8VlLIRARuC7V3IQLrCTG2Uo
tcuODblrLtzCJqA9D8sK6jz+1dqKSWU0KvZ9dVmlN9VFOE18kURwDxwqQNr6sp01
MCY1wNKal+xidb6wFhnOaXD5zbo61TgUHyEXL4NE1Bh92ngtvdKLcsxAAmY1rkGv
exSmKA7EmTpgMpWTiVhbmEGhT+P89XmhUfy0Bx11ek6YfjjcoWMkxFkKOuJRyJ7+
sJjzNMsjZfyrgkYUXkUDIZZ5tt5M/ya+BkyKrKknpEFXx6tS3lSNszWXA0dP55Zn
6wf2FR8fsTeJfwBRqbThfRGDDpi54kdoGHIRy2bVrnO/dBgImxVDM3jqt7XS2Zbp
3ABx+VutO1M59YXF8OhYsmSNMU5KccL2CsW3vdWboHrPX2FQCbFgrm1UokRzL33l
1wRTe4zknqbFGZEzeiLDqNt5JjkUjogkR1pzU6B327EzAi8Fs+shMMP6oAv9W7c1
qQOSerkZkZcPUrKnAcCha8Ajl41JlY35HhNN6haOD70hBmILzg6UD3NH+N3Bhz+t
C4OpooQW8eTszor/M5zYQXgzsxsqcY2iF5igbSFHobfxDzwZrQzlwbMy3VTo20l0
/uFbpV+ysLG2VL5icouStmk/2+zvCjnJCsc7rIW4fBkBgbEqlnarFSmfbQbdbfnI
S+OIOjfDNxa5YFxRJfumeIbNxdyJAG2WOdUe1uOMG4qGNiJY2O30D32fot20WEDS
Ske1/0qSA0cIXwdjRKPAlx55LBHrnp/C36kvuTvJ/dqrYlDzKq0/25XCT3B9+oVc
oxNtHoqwVzj3HhBujsqKVKumUWbAZ3+SpTHQrzpBxMQqETsz/cFqjhJ7FssJ+KsF
7XrIyDSqCP8LIQoFGG5zyDlJjcy7CT4hKFJphD+gK7CUbz29ASAczwIruqRsaPta
kHrY2laNawvuhJtWhW2omaNZfPrqxZRR831ozCzubTvIEF1U71kKxQYx3JuS341W
8t3548a/Xt1jFqfRQLHdxBS1o/RanUyvK/RrZnhLN5Y0EHibg7sQ+gtVLaqGt6x8
RD3XN6Qs+NObBdhPkuP3rQ+SEkVBiRT70EjEArQOFxbUPpEdzdMdjJIr2g1ZUuMV
5XSHsV5QtFYY/uLMi2M9AuTPVftxa0SKU2ZFqIdYxYjipUGugFXnq9JfSF61FE9w
To41mhg9bVwBXZJnl21KSsU6cZpbgYTZsoCSxvXSZ2/iGpV7/vrAAnUl915OZPvw
J4YV2BGUpMj0n1e5KmkaC7kCYzXOy7xd9Ck02k2Cljv5kT6+ilEQlmqfc3pNt89G
TKgFt+WPGdAvAxT+BNqxTrrrJQiKjS5MKqSnm8VxgCsem0ZTcwXKrck0RqaYMp7e
UvVjDjKQLdUdjizze/axVtv7FuC515DwlSMieRFuirHu4yGMBi3kzvs+AVyryVoS
e/R2LM+61k2Ahq8VI3K/uan18aXLUukFUblHj1GTKG/wEZyh+9mrZyumj7Eml2qq
4bT5iVhFF9GH4rJIy6GaIHXfPL78fcR52+0YuGcxLTZAfK11z3nBFkfGnD5WGuZA
fDIZOlVIqRiODb+PKCGMQ421t4oiYzJj4UghRUUvRuSl2BOlFMYXwR7McK/hvrIP
hm06WkbU0O3vaw8rlan4COAKYuStN2FNVIIKAw5kZEYV0b8hS0FQ3cNIwu/0h+Sv
87JaZH6GvBhG8oAHxNtstsFR/58uTRr5Vi8JLufpy1hVB+bzSlzBgEmnpMBYaFSD
HoKqk+VzzKdResj9YggfzcBlCf0+mNtIw8IJMHaTam+vjQz2MxoKSzoTD7vECEca
0O7AJGT/eLmypV0lDaJc3/jd+hSlB9IozIfP8GisOrSJOs3UqVjuJCHJx02ZbL7I
VqNO+fCPQwFGuuMGZYh/+UlDrQJZnYbGGTnh28KpXUEs5SszNi67C0t9FIkbQlK9
5H1u9t4BB7QSLdTdZA720/jUVUfxKTbAMHx1rwhECJ8qPH6eDMfIziqe/DHztkXq
C/mxVYJRprXaHnY7xRnnOBvG/6t/654NHMc/R+SF5KePbaNkx1mSkaQS+dhdRPWy
YVryFfF/bNOfzShNytCA+g65T4EAwS8RwHvD3VGpyanbTWzHXpbiBph5QbZ6wr84
rbLRkwjaAHyZg2kGSX697BEz4ev6y9zcgTl5xa8Ow/jwD3v/IEGqaN07sd9AFdtr
ca8PWrgt4ijzNHNvbdEoIhEgNQYOQTHqm3bLjSe9UO0Tf4JA8m0Fkh8ByRd9d44H
U6Z7g/rqE+IuyMyO7sakJbE3x90sy3FKdKfnpeD/fACzkdbVZLaUcWlcJIwiBoCh
B9uFU4n2166679RZIqrpB/BnrklH11d/KI38udTeDS5Jun++EKreiDGIdrFyDNjx
7k0Wmc1Cb8kX7cOiMyIWbU3Lg8Vq/FQRLgczraazbo4n4Jlo68O6l2djzgAwq+iF
obQXDTbJoGIa/zrxm9/Ci3MUvejqcrmyfTPIUy39h1PaK0ptDcoBexsIReoydoFt
ZPQEKmCEh0u/z+tLp+HOhVXuk91cgjw7L05aYjCDucW1UZyAoZqEWP3q4E324XMB
Oh57o6SN2ZIiU085fcZeB9/6XDPVWMJ45seYSuLU1HUnmtZY2+J6gMJPYTKRqQRD
V81w9F/w3pkX7BVYD1yOFUfXP/Tkg/hGsVrkrjVQPtL2R8XCLqUDekSAymVAJsU/
4muaEbUpTQkr/PPoH97hSsxLhq7fGumFqG7eEJzZcwiKK7YRj3RVnbMWibGuNi4n
2aJHyDKO7ej/J2pOAYorkDwpoZCVOHTF562HHeQgsnn1JEn7nCp3URExrJVd86Vz
kglXwCaAzv8H+NW6sE/FyaO6UOOORX6aDcywQ8KrUQbVk/DBN8yUzIM6JbkHylOP
u1qM1z9x+EI1brtfNPL4spY5OLJ10oXlWwfSurzGv80LJKgj4PHbhT7DF0jSIQ5F
6MXC+zv/NmozIgVVQ77GjCNOuXXvNikft+QBXDZmioydHr55VnbMaWU6b1mS1TXM
xQo6f6Va2ARgLvEMpV8dklVHTtzjlombNTthIhrrV8ZEKYDKEgc2zIUebmAPEKmY
PvP4aTpWWd4ik9mEq83tpF2rP3216PtJe48mlfN1WqHHKClhHRB6dpgPpA90PV3r
PF5DRxCFogm0SJWIOCHwN4uduXQVsJzzHt3Zap/4gij70sU+YSJGDr9XWOySU5Sp
dzwX+6ROENoHt5sCEXpmmZv8rmj3tWzVHFQWRIqczRxm9qMDM6BPL0V/TZwc42RR
yrMRsvK4CUYd/Ow0c2NzN5SiTi1JYlifYqTto3bAQ982Tna95ySsrvLGjWQPoh8x
YwtYO1P1DxaVt3VRZ2yA1sVGZTbe+nsAJHljhvFOHIXeY+GnJsGf0LyINsSS81oH
Z1Zm5ifuIxojSZay3gj+aUi/qLbLHkvTjNw58sUcVS7lbCNcu2NkBmW2Fcv1mij4
IB8HAUzJ3iLyC6citWQj1BGnIeTiXj+rgceVP+5kYaHQPv3srBvCLkIM4suMB70e
+MMa9RwpHQHu1ne/M02O95hcBG9NGll5KXTMpR99xldDtV43MMlnut00OzCsXjCB
Cb2D+MXXHrCPtvMso9otoRkx9SRpHxGtVMSWgBG1hu43C8bEhem/XstY9RL7y7rv
2O7nVcGlWhLnlW1WS/+u8CgDZf30Yey2fFgmHvGUdoeoJRQ4AX3tWY8Hwa/n4D6I
cJZV+incoL8sbDiD3rYo1bMg1sEc1vWnZNg5sHmaKYUf5JBuX+LPorxJhaK9o4I3
U760qZuL6y1LvKkDWgGx4r+eMijXvl9lFuKTfbMkStQr7uoFqqaM/mqtsq0Empui
lHhfkenp6jZsOX75fC1rJvIN/tlz878PU9iAWkdWuaptX1byhDeZ47ydmmdeIudW
wD7pnfJU8EuUvQM7MeWcIUJ7G/gFVVngmF1f0Pz1I9pCUhby8wb4/Qp3lyeB2lJM
GZNzdpbhLd+hQOTw3d+dmbvFedK5Xh3gRNHIXUGSZbNTcQwsAHCX8lMUyamMLM3b
Tp5uKukatUc3ybj6dDoBS7ysoLGnqIffmjnSEoul3s0cJMPwoozCSThGXXYihFNF
+vQy/Yycc9qVnnsPb5OQ0dtkf3QeFYqjk/zkb4Gx9AfW2DFDTPC55rQDI1njobBB
VJ+8V4BLwRpDR/oKcIxZzgZ/C0Y5QQecHVPJF6DSi2koSp+Ty5zB/WJpV09wouw6
HKj7EQiF5YA96nsMnc6l8CLQ2hsy1rHfn0KIDh6zCF/WbAfBZudHFNLFOLsmiv84
NGaYO6T6VCQ+8U7h2/wFMXqzzkMHtlu7Ss9cbFDGi9ZQb7cWmRZNQQn7teeTrmlt
0iUCDPm6dfV2MP3c8/F1e7FOVTRczifdvgkLv7VfTAT/bF/lVzZpCB+Uoj04IrA0
3ldGcEV3LviBax9YnjRgDLTzvWDrWm74GTOmmhdWwuT2V7VpEBXJfeY94bKlwuWQ
rYjTM0krT5PdilDg4f39NI7VAP8Nm2XQfLH0c76L+/V0z3R5I1z1KV6AJiiV38Q4
CjaB/r6JDukzAoNxMP2KQS0hQ2kI2ULOInnDNIMv4RYqY60afXF1GrssDwzQK3Xl
PJ6aqkazk0vwdksNNOGGiC2hNlozUcdbdvFko9lMOp6XKr/C6kHEtbpdze0GHzvk
zuJsWG8/lg/HjpjJVw9Nc/30ayPUmdRL90/nIOomCNofEjekVP2NYbJOpnX6ApeD
XO1XV1xS6xHPncXI8Zs138kWIijuYfvBkpVFCIcae9tWKaX6yca3yAmDjaoXHtS+
HvgoFz+2icz6Eay/8/hjNHPz7YD6C23N+ZzSTUBhW184K8ZnCSxkkVEpx0cDgbLv
CwkuuuuzQRkwAjRteoABTGpZyCaqf8kE/NNbIw9729LA2nZIogZxhBN+4hpmA55Y
81vQudFSq8UepGYmXBr/vX53ajcjdjnGl3BWLBTrvrRcPly54yqM3iYg/U5zjVGP
OA+d++6QFbcMWxxXre5BB0qZgNZ/x4tgaSRwtlr/BuckARzAl7cEy8tjkilE9YiV
55Kkh9c2DiZN2yOgyA5hHwKgaeXp4DrjJcTIO8+lEDfyojS0clr0qVLKRfc6clmv
pMWB3wOLSXyghuSjYusQhKWgig8355KiqeKLOzNTzqCMsqhdtAZMefO4VNmF5NuR
axzjxS7MWgSl8hrPEvVoEkGwDfJaC2+1nmUsXTFStOOjPQgPDzLV4YIVasSBMIv1
vyQqK84fWj08dadQf6Z1xhzPzQWKUrQm4Rcnv3xzdlmhr30XB9m6JoTQyI33k0ZX
/xVng51RqDB/CDY8ou8f7om8TzUVSXUaCFs7bPqj0MoWI4kFubr8N7UUNqKSqsvQ
JlkIi5R02ITOrKCTssWnLgss7MVphnTiEuf9HpWAnejdovQsFo8mv9+zL4g+T/kr
WTnMhWM9P84Ge0BMciwvUc2cJAZhj0Lc94k4mB7RnuJn6EaX4rakp2Slztb7pydG
kmMBiGUxq4BKa5ZnPqpJFQNkcmU/UpS70fVD0+HM9C3Yb9QWDJPYPabrAN8bUxn/
PLX4/WeMHr+veo4DsSzYvKhA78Y3zFK9s20n4LFU1S9JmxQwU+aoSOkfFFDYL+hz
SG5yCDN24TOcKnNdHeCoWSXJznUk4XZ22bOVctfKcaRGGUlFPrefFdOuOFQ3Ip+9
16xlkZNKGg8b8buCiO2+3I0uuAlQ0vrt0k6vUNu7WnhstVMUWVA/XbJkkU7KYWNj
DP4UGJVH8HloAxgT0b/W04Mg+hSaC2d0oCyTxv+4OrghfzoPsiMe/MapvrTkctw9
FoBFEZjKz7VbLeQWSu9mk751dypiUU4uBPSyQa8hl11skKb/mpkNc+XWx7b9sItx
PbCz4lF6uU7Aq+wdIX+rMVJqlyn5R+O6QmYQrujXVIhdJqYvA3txdzajSITc27Hp
sJ2UIWVIC6SuM1ID7OUnn3EweW1t8Sb1AukidOF8FymRky03YES1Guf769vomw5N
p66eO+u5/BGWRF6bwQsPsQvRPToRoCgxXBNPf+arjekC8g343Tl5uKoZfLGpo0N4
no+vR+HTINGSUV1l33KPuMq0dbSijb+ZEZE5C3oPQuOhGE0jJ68aTDc/Qtui62Ft
2kY6XPAd1oACurk+sSdl5repCi3D4kVS1Slx2gRjwRj/c2R8OLN0wX2Q/7qjJi1f
8Gl9dGoFEpckksyZhLo/W1ZbS85I5AhjABV7nD8z639ggCA4Je9pRSjsNyx3giMz
hj39qg7HGKLEeHo6S5FWHLid4ngH0FNYy5JYweJ+AmLvhGP/IdbIMHKeWyulJTAn
d9C/KxOK9/bfr+BkjEbrysMFyF77ezgjES5NA+nWabOY5ADKThse78271f1nHSi5
s4Q3/R7YdCAf8kfxtaO48o2NjSH0JdrqKVCVU4fIIVza5BoRdeEsdjrn+dGA4N51
iQvZchQXyjPFr1j4sqewLP8AdJOnvY2xUtg91IGjfOgGUqnFa/RX/V/mH8VDIqdc
54k/ZcNtP+pEAi+Ut2yfbFLvFfuFAf5xL5za9KO62rtqEVZxr5GASipG8PsfzPf/
5GDVX4r3tshDUGVjVFcDVOSbGX1inpDjcWife2nrNRmMDBA6RzviJIvCpNAOFAnr
wEu15Hdnohe1mULQJYKArVlc+pIpCDSfzL8O27OUyN/wGiL90QJhnO9aCdznOUVe
8U/7jna+Xt9nNXrtJzGW5cP/PZW7iiT7OCCdSbnOdF6FwLq1Myblub+EG7/msk7u
O/zHJiiW3m052rbQVjtC56qgHiBScT3a+UB1xK/gxWHBRitfFFrQrh1KKZhu3+Vb
Y4gpYDVk0xjZAN1hKZMAB68OIBNCytPvi/g7AObaTx98hr+q6eSA0pev8zew21JX
2NY9NjbCpu4B6lVWivjR87kAUQJ3pgGiKkBF195HDOWRPaLZjT+oZytVG5Ns8JGQ
JOcEC3QeaeSUyxnBXDYLB7wQmojFNl5fvCRLn1nXF6XD80i6l/C6UEVsOB6bv+7/
hd1XIh7DzR3dh2W/upwe4gMXlSUIyEFBZ1o8s4vdFtU76XLXGoVv2w/TWUYk0eDM
jEBwj/mdmrZvykJ1necPnYBwRk7LiJLNhPdDyCRfoL1ItyRJdFJQco36lQ1MI19K
VJ5rRBhXt/m59o44C4jGusIu8vvbHdjierdHGpT/keujqiQsaGXBTvKnwhbfr+il
XkB88DZLa8c4o3O9BDnPl4tCbWF8rY5Oye8rG2pC+5yIhccVaGoxhTDgZl9vWRa6
hyI1rMlDFsZ995h40gMa7C9As1t1rkKEQKs1rCzma1D6GrwUYEdIP7yn+YIGwMTe
WKKhF5Af9O5Q/fPdGwzYttFxaT1Gce+Xt5uTWAJuHwGlNkpiDZf6MSFv0dlDEcDz
Bt2r6PVTjUzvKUPvImdFMSLDvHJl9rZaLRhCq2Mmn9B7irg8aQ+GOEFWUe0N8vJd
WahI8ZWefyZeVt5p/KeXoapRTEiQym3cl0MN2rZeoae0go3nH4HoulXFV6xXSihN
KTIsjNIuuHnn2kUgt9ZNCrSyFJlIQL+F/AzDrQrb7jOv2u51MQW+biH7k1h8/m/D
si983DG4rKqBMW9gnChP4ZH93S1Sx6rM02k3G/6TIGGAcqHN5lYCW05UQxhl0odG
0KzoW5TbeJdRcYr1An9WEeplScvKsBwaA/9va/pkriQuE0kteSrvbKzX50tWNL7b
9EwLb7snC5COOlsXtgVtRkxRGDJ8MPfU2XXoWDl3vECYK/VXTuhJnvLYWo9Nfq9W
eJMaRtlqCR3sogYkM1mLMu0UoGUKa1xnEN/5sdQtOjLVNusaG4m+Fw4ajbZub+nB
VbN8xlNIO9ebtqT1dU7D2ZsvApydy1kpfSaPY79KQMz2AQvbLoIZ8Z/61zgHefVD
cdO/C3Uz8DF5yKwiNiutsYcZJZjurQ4iqX6WDfor5I/T6wOL0xf21yfmW9QpTzrE
xiG9lL29aCUfIw/enNMNgd8iRjikwR7aXaarh6OjgxgDnKf2r1i5Qj4K8S0n2FVK
Dc0+z4UZY7Cww+HNspJ8xX9iiPqyIg0+yYUV2JoaY2KmXS4oGCIxJC+IcOPoRlwy
vEKzRfuT1xaoVhvbSr4fn6+yMPDtEYTbAnTxmxOu3dMUemrz8naJo/Vva+x7cn1m
LwPo77RgbeMEpV70kp+3vimrjEVqZjbUDgJYPD/x+mDFMX92Ns3YVBoTzzveD0eG
eY+OvqhCBNxgWrGSdM6YL1+wF09RwODBu+O3t90rfr+Qj9ZG96bJI+GSWxxA9RhV
7lcuZyS2VzkW6i4a6bCAh1KXgT/bPhMYFJjga4UWBdUXv7eUg6akyO6+fd4detzc
X0TtrPqNohjEdpUiEpOg0LNDl/6HLGIQ6WjAy/xYRjqaMeR4TmhW1DbKQzM+lLFv
vLpiV5gfoQdHREd6DH9HM0uQpngHZ+DuBqPxHX1HIRwENS7qaSpSTWxTDzCyGMNu
ZpmWr21tw+9EsBTIMbf2/LzVb9DR3pwlbYNy7hcLbgeinjilXh3glRW5LbvEtYAX
Rc7t9XsYbl/j7y5tz4Uz1APHbF/mRKm4UCvssYbMBRE3nEXdA2yz8mnXM74w1r8o
B7qixZ9IHz5W5VSzQ0Y9U7EpzUkQXdy3A2wcKK9FCVfwSNHcTTATRnpKAs2ygzg6
KF5v6HJ13mlDn1NujQtt5LfrRdz9Hxa93ipcxzJl0uhWtki/RlKZpR4HZHRAJVu6
nH5Th+C7IqFG/cGe9OyEC6mh6RQA5zYNgI5yGiNSF1uQOSZUU3hT5Iq1hmmW+uF7
pEuDcW2hj/AXOVkdfkEMSddwRiqYwDz4i+iEgK8xVNKnkdxYf1ER9tnktlAoKqk9
14dzx0yFpiUe6G/jsFZFEUT0iOlyTTaY+kAIhS+/KlwRuNHTQCvsv9Hrmuck/UYk
cnugTLw6qUzKwTWRBXIZ7j2sIRPt/yRQIDvW09DKDcHj1YkA6Ya+mOAU90XK1njy
zS9eQZBehAAar8KSyzK39mAm2dCUODXAq9z0nSYyIMrBGAeUi8h27yq+Ft+F9BTp
1aOsBr3IQRtyI6Et6CbpZlz40d/bG4Rsrp3Y7sz4TKV/fDO95y6ZwCoIbakJHKql
gLIoPrZQgabIIPgCaCm6puE3G1Qw/M5+LYFi+XPyIYY1gCIAie9teImRyK/muBbY
wPBufIFr7bEU8d5TJunXLfUAyo09eMRaOa664no2jQaYvOxDJjn4dYMWw0IZtu59
cc9po9Nn+v8u6ZoQuo4DkvecBZjaAQdTIFzCfXhQQr0cfYdqme5ypFacFRP/o/pc
ulHXxmxciuBTj0hSLDLkrMpt4Y0raax+Ob1MHXf3EutGB5OD32q/kSUp1jDBQIU0
xcokhDSRKopNr3J95OZdepje7OxarBWMH+dptl3Opn4aOiVZsp8QutwkLP7mdQ2N
aA24LvHMu3nLtw42Zbk2dvqthBwAoA6sNQYzXzajnK1Eg5+pJl79QktS92lD2tba
9+gXLOe50cStuQvucsvurrZXk7aXyDwdN+Dihv/X/RQZTGO4cU7sk5ydDZ07Usen
xjpaEdsnqW2KVfHTudTtqrXkfw4+aF2K5BP5t3BP/vM8rONqzWElOJ+ni1HcZ+sp
EsNSF2mGgLle5Bk0fMcYhaPDm/ZyYfzWO/Mkf2bsVjwbQQvoIG2zvIJxydk7gb10
qHwyVzOtG6/TYmmOPj3to5Cy398zF4QHIDAIdyBjqg7cPgabv4y5F9RikfHvBliE
wZU6UE89/E5yPKC7GHcP87avH0oA7myJ0h/sRj32FVZ+UdDOj6K6ATKzZ38Ls5Ln
Jn69x2cHgFKPQ1k07vc6hq8EKOKh64lLeAUr8m3CIvFFpkoPbmPTQPPpctPihmhc
Ogsex/FNLrnr2K3Sjyq/xkz+bV2+x7BOC0n7bWaWm/qRytb2qHxA1hnrjfV9HSjE
rp/WyWFaXPz9WmkKp9DsH5aslHAy2wPafOEjwRx7fTz2vj/X5MTcV8dS0u5Y5HiU
ytD+/6luoC9JJPkavde9DJwqhDWBTk5SRCW+Y8YFIjFShzSgJ3bDkhMyJMYPcbf/
F+gGuv5w4+tZ0sz52aq1JSyqS9pHxo//le0R5xQGq2FPiCD2C3sL97j/jMXq0sX3
jEeyrDviV0yam4rngmgbTwPfFPQOmCgdXET70PvZOWuXAtf69GUDI9M2n4Qg1Zs9
C/ClCR+gM2bQ/Nduky0yitSdP4gf4YmQiiSYWjPv3drZLmh9aRtgnCnewovuNZOS
0H+8qLqw+vDIBfd0G0OjXh9cL3DfjRqAzC0pfp2M4k7tPm/M+PtGh+sAQavNsjIw
RUbWJBm45WNOZXQ8YYW+0e/HHWZvXyaR5FKtB+YHwcfr6KMKtClhF/7L+70l5VX4
nnF3Go1FUu56pazvZsBQskThelGFZILm++vashqJs/mLDJpHjnaP4Olkl3yxkOgB
12kjQrcdXF5ym50KdZTOBUVJ4IgytjONi+hV91e9KKhIbJ/tXrkLxRPYSGd5/rQL
2W/nfN7JIaapU499IKk9At7K9sJVW4v3uKrYGha7dGTnCtI0hlxT8OPPsjqnfgle
H5AX455z0dkZbwEQitb5vEjFGAFPB9H+rTJk8gossXvIXCGTYzcK9/mpKCaaQzXZ
H34kdPnqAPKT/Nm/IIiQDNRz9SvIgjaOOhi/wCPuaq18ceLRNDxQ9EN25nYNhm+b
c1nFTa+UUE915bjRGQMmFRCFBc6wCKjFK68ZHB1DZbPrCLNNrcfMyuJcxwUSnk6n
Du/dDlDUlIC9Z/pS8YJPMI11uP6tV47yQe+F4OUCKsxFQDVDjIQ83twKjUU6iimL
JGs3DpmZj/CALgH/kcCPvJ7/0lV+JHVhDMNgb76sJARbKn5Zv0wn+oGmmep+b56a
N04rCuNLo6CeZq15qnneKy0hEsJZncKqZ46Ew6DOUKwr4UeITYjsKEmulf3Uu9U+
m0Zf+z8yjxuocRYuAPjpdlXjQffC3xIVbzzqjEyK5oqheu8Qkvw0eB+qgo1mz31p
LpvDlnK9KCfyZe0XRyAEU9kWoL6IuK6RUC4yCkpXupi/cdAwj6X3DMoBZtVTo8jJ
0yoTxdQzqkqZC3mmirlP3dlCDPGwVLFDKGBhGVfSZWKEnaR4cjmxmeGVukK+Agcm
BoqX+9KVqvk0O8bZ7IlRkPVqxiWVkc9olZkGTqgs7yjJ6uWQ68/P7Qfb0UsboJ2O
nXvqGKbn2e8FMdujS6uQkb30ST8YpIbYDsxH7wrvjdWguGCVVXKdQoa1h9Ym6wcP
+UDIIDkExDT3eRkNRbxvkiEXFEtP3rs1HmqGlgekMG5nF/LMF5YlO3nsjpBIn+0O
PbV9DKw2S5VvmNbq8pd3fWkjBMenh93xlIoGAgSCIwR1qBnQPgnK2x9czEVL9eox
hhc6OCBRgnMOiMqOfByzHvS4WwkCj0nwWSKcm0P0IvaqDrh6vMZGbTVDeWvfwn/R
0AGa+8jasMCgqqXWnF1Wsq02cGnv+ohlhtlJ7GvPfio68o1Vo70VjuyRpckrCyIN
xeE5bPI24/SxwfNubkrcFCIgVb7Roc0xx9UikywE1F4dth6t8+DQMCiKi1wV5xXg
JYnnG/we7LkiwewJfhBSLf1hyto0qrG9/u95q6ThAqnGoMr9G+g9ohIjkxLU9V57
gRyqCbCWNoEEBVtCJ/iwwXtM1fE26zSR9xZKhx0IJLInJuJ0BlIKr8/s0tz8ypaR
mKtmB1HJAy1xaVMElnFcYU8OiEB11viVr08SfXsyMbEi5OaPxZMv+yWfx2A/drRE
mJRHaqRdg3/LpI4aG4Fqt6FRbEEUAvCOv+3YR+pSuHgIPQeE/s1N3RfZX4IcVt0A
18i1gjt372I3ccwgTF1/nKRfADEcO2FJnKhVVR2skB0fg/jyEaVfNhqJQE9ecFjM
vLqApf0mtxvQOKHWiW3URyVC/wCGl3c/tmek+X/2MhWaVbq4algSaQAVDtcuqaog
KliV/UM96qL2WekchgTlsfEB8LpgP1LZk1YGnoCaNLLe2CXkJd31gP4VYLRcHohN
kyEgUVQCKIuEhVewIdCjL2B6Tm50xCA8SlIQQlZh7XmQp1A5NJfOi58VMGBiX1Xo
kwFTQm66uYUbx/CWuSVp6uLV0+Mf0JVGO8jZHfovUW8rChxpZireVMYMX96SjXeR
9en9W2QyW8/F1fI58Fxx6YGPKZY+g1HfUDRot5BCno2DKrQE6n4i18Qhz6liCRqx
Kr9CZICS3kuTNkPYWtOEhKW44wBX6FJemBKw2KFGv41uUhHMFjH76Ni1Qo3O0LvF
w9aHySs7fIub+5pGAxoMB7J0Y9IDiyrk8wEX3qVAbzPspb5QlKB7uaWdll56HMD8
66YArUxhn3uDcNqNhlznku41CcS7a2tyz7ypW7uvjRE4C4jpcxzmKDYkJgAXdwpd
g/lA5L7pYE2P6wvGK07w6NbNEVwRZlBV7TBi9xpc21kf+sHvk+6feVEpPlnRn1KR
wX6OFxPfQqI4w4CWL1Z1b7kyBaSKh0kktc2AMSAeO79o+S605l/2wyh/AOGlsrjR
bR+FtkhGM9r8q+oonXoolpmCFhjPoCujCjNEsChWKyNJb4kN/atW8a2RXTgHtlPT
x7y6Rfnh2VCzTT4HY9jPDwMoF/AZvvlGDdomIKmsOuV2x9fuLCj1wIxPBVsmQfHT
872OzW5gu+MVkAQGW+SLjB1dj35n0WD4Z264p4coXWeLot90bv+sc6HyKe77JPK9
tlJPvmdubwYgwzVeSroPl7N/r6M2wEX93eIiILS+eOvzQFhh4fNaGOmp2G5dWe6U
gSw1ocj/1BAEcHsCnEqLFYxf6+Vbo6csJVbkia8vptADD2fX0C1Pd0zWyi+p1/K+
wBOONeq5bsi2GLb+e9ql8r07WaH05Jzmz6MrI4fw+0xYl1D8j7dDQMVMqf9b404x
rnEy4efMRSkUKzEWbtr+d3mCCad+7V7EZz1WvXrPP5XpLJfI6BioBvMdn0Oaeuwd
kKRougCTuFdFjrHr5HunXSzo0oJ960RNBdmhndrvywv+i4mrt1VT/G97+CKf9Yvw
eO64Q+r8jA83qS5IrAVuhEAz53fT55AVRvGPKWHYWAAKdZ0nuXKAk6+ld46kx3+P
vUR5+UQEBgFVo7GQyHOZjAlQfQoIcDbA9IS6gVdYcwXphaeK/DGRzzTtfiyaOkqw
rAbHrp7rfGShdSLZDmODTzUpas1a89eoGt0Dabmbye32nizZlYXKAc/+/WFRU9aC
0BN86HaPyM7FdLhpC8icrgCU/0A3an0ko2ji/SneJIaEomyer9e1CqlXDSXNLXfS
tx36jX+tseee/pxms3uzvDaye52sZAcY7c1R8o2cwI1voFFYyywgilm9Wfm2fIPz
CPSfMGd55uozfB+/fj/eDcLGWy/08vRK6HW9H11iAjYB2F1VXIQHtqRwlxXh9idi
exmRlbafBlXCSDE7/K1T3gs+wTnDWntG64Vl2HBLYcvARwulH09RNT2D7oQ7zX5U
JDrdUNyHW+sll39KBmz1wbe16o2BgAKZb18HsC4tC9k/lDoFIZmfbGI6emaAHf7K
VX9pOdZ9Zrwqcaduy+2CRA9bvF3Jkn+FCrs3IGgvjaP9/AgcyCAl0T+JikItYo42
gEKp5tQed38oKcLJ8kZddO8fKM+JeqMpFB7d2GeOFplG/qbmxDaFX+8QQjCnJLaK
aze7RptQ9kzKzZueIv8BmGWQ2tnwM4xGzm80w+rY5f5pG4Kxtpp/eJSU0+1btqLI
wDVZ8vgSPpIxSryIW3rW+t/joO+Vz26QCffhQvRxg/Kjsy6Hyc+lCIdewgKrCDxa
boy4smO8HbJw4ImhXyTBoxzSuAfVx2dxc11vgegTnVAJ99QGgkDj84X6b+A+CpyR
UiKvzJI1j4rSZ6l7aEo47c6DuOWgAWEUcOU3953Q8aRDabo9ZeIqIlrkW2lKpBlm
q3oSQl0W4U8cTckyluXI3qBFsBNe9Zrb7l1KN9/fbUBvaPA5A/ZJoJ9cKHAimtgX
aZr52qwMq12ZbPN8yqrnxsgdDDeiFhRwHyvMqp/bzUOGudus2Vc1fiImWvkqiVdm
MRmwIIdLN+R6e3s9A2zPw8RjHvN5cskvU3R5Ij22kqnDIBw+Y136Rx3Ne0buHWgp
2/0kD1ntldcgnL8c9rtSiXt5ZmbtBh6N3ki621oNneCUImiGyYvuWxco9UmHYusm
lt/HrUWbkGmnQYWSh/6qTLaMbel/5g4Roxiqz6xO8MGd0KAxX+WYBAgSe63keQeN
/IoCJvWYWrC1pKgqr6wRq7Y8YfMw0mhE1ikO11N1ie4uvKTmr0E3+KhOxTqki5GC
6bjj+anEzacgLR/PlZVBG3fXinynFhwKjDkGr1dSKm2leWRoqmH6BG45uIJI6Ybi
on4s2D7oE4EAjWA7h7tguqGe6yqkNkiEzsjStGy8HT46TF4xvLfQ45iviVLy6DWz
+ZBqhtVb7+DiAz/+mbLsauJyHQ+dSUTJYyBR0sHpnDvCqMLLUh4qv/7V6mQZ7A4F
pxNedZ2qjv7iELM/bDxo8j3fDzS8MYULxVMAfYm/Gh5dQAtTpuIQZghVrTiVKVbk
e2WKNjXdO3zTbJcsOI2ReLne78lHgTi+xTIJwo37BAxVtgTm20de50KVET/cMdS8
dxRffccOoth0mntlbLTENAVvnDmInDPFPniNQFImteuvqCXjargzvDa27SmRkP6m
DbyN1KkGyOvO8CE26H0ARuZHqpE86ZASLuvsJVE4UKQEG+pLlH74H1vg/QKXqkho
Vu1vipjCDDUbDz6xPvoGOvEZio493MbvkMoDy6TVtcoee8WO2+fbQrmtAU3MHsWM
5YnhHC1v+D7aq4ACUKK/Jao47huJKgj2xPnT+NZR0gA5Zm0tgBXd47ER/8Tltdoq
PxhXPBZAquR+7EkIQz2qNeGEpcV5HL9Nwcfl2GIcwVNUGdHdMJezM/ylzOO/uRoA
7sGDwPAv6qrhlWXnPperJzjwlHg3mTQdkChpVJm/TiDlOPvDtEY9UB5mpx0Xplt9
HuKzWD0epKX+JfbzYMJ0mWz7aMxlmmmqaXaShloMYus6/PTYKZknkFrWdjnZ59c2
v+YJzjqi/KBIbNgBANYBsyg5e8N50FvcY1aJBxpCotcBdwGl5FiKleqLBEGy0jLW
l//qySuwAvr+6ZV/9arEUmpbdlbUSvrE0Z9Gyg/Wx+WXL1GLiZTgws7JXAw7M4hj
b+Tht2OlmmVChdAbnT2OeWr2rRuQ8y/AX5BqcxmIjgRgN1RJLV2CZb8Cpq9MFVDj
/6bMk/5po22vP0r+JkM8jUI7kdAOU+W2kG5cd/JUOfwJ+tUKq6V2dM3zuh3UrppM
ik1tW21RAW53f0xm9lrr8g/647M/VO1tsQUio5KmvXcLmAvDypHUIYTpK2V1xioS
5A8EeCizhs7BTnFiu8YVO2BBTVXqxYGqNxkwqx2AqI5yV+nSThog0cjAlBNYgkQU
iQQLCLsz+pTHRlW3jWWzD+xh/fPDfXxtlTV0wN/L8mn82MTaPqBAToa05xm2GzZr
EsSCJEmUM/2Cik4b6orCZC/u2wt9mRSI8zmZbuiJeOhjU8z/QJsciBx+/Lanmnr/
xI9YBNWCwNO3bWw2CLx67ogZE0az/BBI+D6ajBYVvvQM8CdZn3RMtqphUgrRj7Dj
GhS1SaHZrTRtQrMLclzdncB7Y7hk4Wn0ahBnf6C1Fz4Q2YcGPpTZ2UWMPiPHQ6DC
v8RHQxt6aOPHQARyPugNe3pUnz6V/WGdfWmniNVUfW+0PKyYtZfjVowFyoB7x2bP
piWsJ/FqKmGsNFDR+MNGFSsR7hSpGPiNLtDxWgSUDFpv3BQHerwXhqnxm6Aqfvym
dY/wHmzOWouLZWrIQ5f64+SQV3RRjOdNXONGumVZXumFyJpQr/CodmQGFYVlnFcS
H6E5uJ0LBII4A5sEGZWKu9+2M/S9h+ad0WOiSCSqhWkO2fNcqEElMo6BGbtywLyd
hKV9z9Bi1P6dvUHSTCNIL1+TTJ+qWsEJo5t+HSfSrFZNAuss4Ibnkykt1MXEwnDx
pbPaF7WqiNRlYlShQHSpP7l0r8GXei/WozVZ1T/QfyB9BGf8UgY7PzJUZXwueY8P
3VznesLf7q8jhB0Uw4ORGstWsuMBqRiter9pDDgnjBtxZKU+lcn+WF0GeTky9j0F
c9gxUNxim3qlbuSEnSwlqgTy11HuhkwJzsOx3AbX7bbpHqF8JwaSVooymjgKuvhC
YZAdRnxlm31uaYfTPqG4F3iCzUYJlGV5NEG0Y49Dd2Yx8TTwsbvAMsK9F5GXed9f
uYW3wc1sGv5pRFUa7QREeZCFYtJ6uYxGI0BJp1B/p/ssOxYsgJgWfrbCYQYtDNbt
+Cr2YTw2RuRwE3rvdi/SayjFT+iASLHqpUfvJcy9ySNro2QU42P1hleHSbwOKK3v
VK4ScDN9iod2VgFVabg7OrNClXpvzuUplTCDt6UjQWSJnH3d0CKl7uKITArwmeDX
IgWInvWN8qt/EWJUYyO+41FQKZY0D1iIC5104Hny2YAJaNxwz68wPNKIHVif4ZsQ
hfBiBingqzLRH/Wy3DDOMRV4lSwZdtilY65M2be7tW2w8ScrRExdRidIm1STZbtE
IsWn6lnQozr1H0YOc1To27W55ew+y0wSvD3p1Hp8MNKFwfW9OTwLiMBK0nWP+7DW
Kh3fQJdsUN9rBU5aT9e1jOcyhLzHxYwzdFa5t7tW2p/4skfqfFzs9XoAphGHEN+p
qx9TYVEsZ0Ieq8pRyAx3qXaePRNy28Wlc2332UCB07dDLEOxsa02Re04pQex6m8H
szsXH8EumRp+aisR7mhRSJaHI/igvROoejPlLbIqzjg3P8Zi2LEs+29CjntskUKJ
Rs5HWN5FdNTLljlWCnox6leTAtYsjEBms0lGbXwqkO7XRgzETTFCv5/qyzrIsNHb
lH3sBXhQV96Y1hpgP2gI+hkBt6oRw6uWsu7Vrw3L83XE5e2u6K+CGsJ/ufcoHus5
ETlET8mdWTkkFI9BOQYWY/ou1QpWRNCG1z6RCoMQE3lpqRQWSRgMLHJJ5/LYYao6
SIP5yEGiItCNurQ+5hedgI3n5jx91szypgz9Yr4XLJESaYG20vY0ZppY+pwsqehx
gW6aiK2ZmR0oHTE00bBVTzKBsSQ9PQ6cEq9tNAvnxn01TFrqJ1TBeVG7R0/NHi+p
JV2aytiyrS8yR6lhgp+PXLwLQlOF/NosrvjzyPIiznft003A/J4DVmCY/SaPT/Vb
zDXw3IXZG/bHvsvdVMSS7+0CRpYRXikwkMJZSzVtqoeCbLQlwjViYDG53lVKyE8F
WySnKVKLqzwWCkERXdC3L7PhLYqI0/q8Z/Z9ZbJNhzuctsFKf+65Q1lrFMLV5Z8M
taGzF3hhZeu+hGbAWtYLy/U+eeB1UTR8OPAA/Tq5z+UvVfQF0nUhKr2K7dNX92nD
QBIYs2rmjBOjzL43qCOJ7nQ569dHuVIwwoLlP6Vkv4kIBnm3OjbEUulIXQO5WX1K
zjtDFIwFaMQXEi+GD2BjhgtwfOuuCm91jJI0seB0q9zewakD3qfqT/HtKSRmtxlE
XGOjjL4yYGfzoJuvYvpmWkbBXCi/guP0sRn6gOKSPOLhFUgC4oRbZ5Dl5FAbbSuh
Ye7CO9Frqh5wSqLSW4LAWMhZbrM8Xo06oEkhIU7bK1h1BwOfxihl5ufgtYj3ZvH4
TTCF7Fvv4PvrAeqEWmBw0JOJB93eNx/M25/AvzfL+hWi5gIeabzF678kUIbdhKn9
vQdjba9M5x1azGrcdxBZz+KtFywmtVY/jNJp4UgSRKkZOn05GQChorEaDCrGNwW3
jv1dc7FL7aBZVYI1VTZW1RnIqVsCa7Wb36MlaG5dHV15zc3N7PG1Yl4cjDntlJvB
Fhtnmh6aJwyOu/ssD0xOw8LwB8BoMe8pnOf+kf8FDplCxjWIH+Z2hrDoo4HL7F9h
CT1YhL2hbfUzh0sYraV2FUqLB2cfFqpxYMidqogzutoi5vJQFjdoaxYS9L8o4h6R
GClu0BftxIWZeeTVL4GYRfpWiFx3l9PV57GYVpHf12xmYhb/Xn81PqFLgU2xHRo5
P1sxGVBW2WwJJQep8+PcTMErOAoMY0bDzxyV9gzFp69MgiShdd0ixUz8PHrpdN9C
7/v6GCZnGalNyeD3oLdpkhYiFOZwrqe7hd6wEzjg1pRpsAF3nia9huHqJv6oeQvM
Pj/ySahiZMV7x4sbXuJRFfLRpDnB7I1sxac0iz80igXY/ExyllTeQB06qsQ+IoL2
VdEJQXaNiMoAxkeqpIJ81+zH37vywWrtOsbF0oS2XaF9BRmRF7jVMaH6wVnGIQD8
qMraUN2i9OjefGC82oS2vNrpCWcWgcDid1fLbZUsb/M1m0nevEMnmvb25kR9zytQ
Wcu9c2I1/2SWtemrM0qTigE5BtdGrNa8jK/oJ7K00T797bb4icnrLk4GyaPqjrFY
BVWN/29NG4KkMuUjcRvbrylTdyq74R3Fpnqpa+rHBCdXUPMYbdlZsSdLYhy/rO3M
8P83URdDYsDEbhrIEpZj4USaoNDCISxrb1Y1jVEyUMUP4aVRUIct0a4yv8Im8PMy
HJL16PnzYUU0EVNiK/up0LnDE+89RYPCJKwD8JHCtM1D3Do4miaJMhzZ3I2K1wO6
NwngK/kegidQgO7CjYsTovHHR8nzjIvMkXrHMBEQEE61yWQTBsJrLC9pvRp8gBdm
soG8imvGlHZx0M73a6HkqLbIQIex/TDEIxfvp7GyXnVJ+jpsgaJs2jlxcW40/tyE
cJmy0MS2sN71yRFHPXT9TzeluD6kvZSyStXqkZqO6+7IwMfEShWyEgmaXAhJrRCQ
Ikrn7bhQCI3OsXJ5iN2vdcmfqsIb5fNQUpWMxp9YEX1IdEb1rDqpu02uk7rqX/sV
5Ta3msqxrcsKA2qmb50ayRbFWHhgg/Ymwl7iQKhuDIUYnEmbLNgBD19gdtGZc5jc
OHkIzMUJkQlPJB5vxsF68sPz+6dvfm8q5z7CB/xsw9Eus6/YmWwAiKLLwuB3Ur2p
PTf5G6EiRzaiJnbfjTiecqg6z9EuaZQNHL5xh125PgCnhIz6iklUhnpypit8106X
I/FGJqpkpeJFlxvGsmMNHM/zrcGW60C8zzjeFDmytEN51WTiA5NNAikDeeXKttjv
m6WcM4svwD8BNXGZx/Xecy/pTwkq1t9OB/vi21kyHrrCHQuCbg5AXjNIEe3JTpUa
+MeTIbHTCzbvAOVabdxWNW4+xwF4aS3KA3OVtoyxl/6syFbw19zLtZBBDwJQgeVO
Uod/g3LOFb7DN/xNtKgJi+2uZs5csGExZrleR6Kd46cQpryEFfc21KQwjX+i43mN
kozxiT9AasIbUmgsxW0xoiel+uIBQ2OpCjLSb1ZWjDC7n6EKQBXO7lELf0upwzjt
D/7cKmR6l5BmuZHWbxiSNQOTu5uaTpmjlStyz/Jr1l2D9KG0Jv0rZPwcHTshIcy7
JAmoznitlq38wUiRKfeqDHrl+QsScSusgC4zrXmrhUJSSTtgfbUZrNFpAO52B+J4
pz15+Xj6pDyIl0uXCPFg4uuhG0T9UUGtX93V7ubyGbPfR5OV+rDlj9KvvGTZXC32
TVwWnw1vpv6OWidX/mNZkE3dSOPzbnyIkyyQlmoXoD1QC6qvJ8RK2oiA4m7r80wJ
YD2WQjIkGIMApjERSf3hLPfE/MyAxznEfQiiYGrmVY+OBranoLbOGSczvy6spWlH
mbSh7P4v8yM18Svd8GFh7y+vQhCkkV6m61k2FAbd6qc/h7b7k9CaPBN28j/KUjN2
e8JOY4XmfXU5HFykkzJNmoitDaAqzU8YTJ2nAhbQMZW5QJwiPiM4aX+S3+QFtJPX
MBU32s5JyHG2sL78gtuWx9HiIz2h6bDCKFGpPcyJlQ1j82lcSjdv4y8a+NP2Rm3L
1SmKTJ//Y+EXm0L1tbgrF2cIrEo7Rmbs6uP8cZkMdWXXzUE9dlk8BKVAGadCDMBW
6PEtaV3x8yIZ+xtPiVSH+FfMptrKj7QiOo01S5IiB6dCGuSkWKzDDzfOygRV2NcS
BLZvN7MyDjT9kAmy/JT1EFsbWwT5HsyJQnQkcuVhZkhVVjtUnI531iSAY1+/G9E0
PXaHsvfDHOBaOD4cLS9zOtbPpQRyU9LTR+gb0xy+k80ABGk7ZLnfQv9j58hLIBgc
tbZB6FskA4s1UKhpylEeM+kvJZf0JmNOiA38IQL1wJpXAMgzp+DDliwShccU0+8d
FirGT8yPx4vT4A+IgPxHthcJeyDVuqGMgjD5/gqev2E5oEGO7v+2XB01wGODwCUi
fYxYzgjTdRr9QW5KpxtiT6oUcYL2OZU+cot6JMT01bJZxY3M0gv+ozyKZAZEjMk4
p46VCxw6vcVrXuCgKW6yVKJQDNXLwqFGl4qah9sCUOT2qMdxfujRFitEiWTCBhUb
aWJKsL9fJ+3kmxPOsTf5/F37Lp2motsj1eZvm768DtS5LDZxIIhYei+cy4gQS/qY
vT1nmt/2gIfwDNwqWbJbiSc6lCqOGOmv5qpUQ5ZGTWb/0ru0BqoooD01CtmN5gxH
pdBnathaCZIV94yNIpnj2QiSC0byin6Fs16RERCtMfxrnak+Xbf1yfqXffaRjljg
2YH6oHSZwaRmNFaTpTKKKPHiAv6aPBlBsMcm0sI5PdoEtk6rHGwMhNyA9jHKdJ8J
ymbjLTJ+OGBTt3YKhwID3z+heTySK4R5ubyNbTyRJ2DTEmNQPDod2oKEZYBFHPit
VBNPCMbz3P8dDkiaNizzaq3SDvq+IsRO/hgDUXib69KEk0sbwWgy8lgPimo4yPyZ
1YQyqfoGxjLo9QoosLJcBemxZDM8CwkxpNIv5QMDmZGdFKnYaW5uvHbJWtSXeODU
ecsdmZP0BxqpBGAYNpnDXLyYMSV20TQI8o7aZd8SVLsJ/YSIQR0tNmw1KNMxA9df
fktpVpcVU/FjIFPbkc9K1Gl4ReyGlrjlsueExCZAZUzpBAs56NEuTZqBQTvhLOdU
9AcNGdmBIMbwufsrckzrynOjwIobPIm5FShbfnIE4Vg7yXUXggVkgH3XMR/1YrZ0
3b5oiRFpVbXDjx39lehQ0iZebC45i3N7nDXjuFqo45NZB6y45S1ifqFYvx668rMk
cuIdtUK/+CFLkSqAhS8yhRbhSpf5d4m+DMgP1LYUJ1X3eo7LKs0n00MZ2Pnuio3C
WO0rUQ3fA81G4KBd+cHb4s/avOuxB/RsKFvUKhXrCsZSNd/h27wIsyMgCthF5GKm
8aUBDld1zQjSL5AVfqSj9IoP9j4Ph52eqOH+Dtg162E02chHfC35KTM76dzmNvna
Yp5rsodMHLZCmsxeczAhr8xqcSt3LbC4KuVJmrye+OtGVzd17BvAYwfSa18iiuMT
/HtSL9Y3q450jfoL3Q4CAdt3CJ5FzNOzIAcYjUGlX+OVZaiYrFrf4RlJ9UeA93hv
1R+VBe06ebjWUcf7LyGNOKOQUTAbTDc7j4jqYA1QGtAbBqR3br6azc8Jy8ACRaFh
Zz95MpwDUd9+NtV9r2Gxi/FLjG+TLJ9APR6+xertna5PTdOvCR7kc8tw+hqqqbVA
eubK7Yn5wboGWHcRavfF10vfpXvWBaMKn0+Banbk2XUBxgwZJkVQVEUMfNa8G0Gk
iYvtT3gRqvFWWUxKczUf6R21FGYj98j38VVx8o4ZQHZz71LHrVVV0eMSNUPJWjcJ
5cdAf0PYUhI8TOnMgdljWfrDBHwcBCtsOiOhvS4HqubejZwfRoC1Ty/au+w1gHkx
ng3v5lqdydYaorzOIi9IY3oOekOHsxR6uXF89pib+3TjG5withTbp+/b/J/YN+yn
I4yRwguQlD5G0iKcBPsPb74GBCwxEJxoYwkN2LwND4pX6CgQ8tQd7rAab4KSidhB
+bsXln1sCXNipr97vSmgOg04j9m9rIHMYEZd1A0W4RE4vf5Z3eaUuvtXFU+qAHjE
u8fW2EvTAXVSKwrfxqkfq5FztMXXAfGX7PmFW0V2e82IeY1Zto2VOW4L3VGQ/8GX
gtQfElpRvSFdDqMVm6qctesPE37K64GFrH/JWgV5Rowud6lUoQcQhM6uxqWMMcdN
5EGlUqPlo47LQMv2PqOlz8AdvbzUGp8xkLw0mRky9K4fwpqdTjHXv0yaVddoKyS4
r/A5uQH6qt3D+XVrLt3lJNSH5MB3G/JWhBQzxivG6JYkaH/kR0Dw+/RRMXhxVhU2
Mru5tMXtO6YvB04pAQNt/QSTK9hgR5XDXUjmz8OCdgdJ2J+5tbltOjFtIv67EOIw
t8GKxcnjrmxqAE2uLLYre4A5PIEtUjajSF/U9Jl4uwyHfKiJX6SKj0OZYv3XSDvL
C/mnafobMYh3cfn9Q2HKrd+rTd24KfPWwhrJ2Zq1ApjBiQrLheDffeboOkc6JJTR
1oyitsuEllDmmm4XrzNzlJiDAfVyJ3m+UdXqRPT+mo43jjRhUL3io2H+zkzYpcvg
cgo/gIexMlyY6qcGFhV1FjJTCcpOX222YnBBo87aZEZMENunPy6UhLoT3OLdbMDT
qDiJgRC/MFtYu+8YoSDG0wuj2dsacYA56IBj4unygeBrcT7DrM4U3eF0tm1323/g
dYvWmI+GXOnRtqLTNM1ygltk2zKC4fl0rSAlQ0LNrrPHx4PsXdWtF1V8z7szMa8Z
5wc3vGnrjxNe17oqNJUABRb9q3EIRW+nzHN0wYDuU7BXaKZG7DbUDUm/5sv3LVd6
GdBSqwAIpA4OS3oOdZyi8iGmFKr7U8OO5KZnzwKBqb7JLYxsbSqxAGe55kV9/zE1
gToJxSAi6Qm3gSGl7vsvuW5l82aMYtbKAOjg3+sMXPVzcmGuAilXLp2dLXyTjquZ
d1rtzFrvPPlyEAJfCa7X5WB4lILRvfkY3L+7qFoSeStWOqb+9ACsiRGx0A+GR4d7
obDBhesKcl3WG8INYPqXyWaongdt82r9dvH3XFF1/TEd952nTfeW7G1mi2QItAbE
4n9Iu8fna5ov9zabsthIcpRl6DU6lonZABHJI6TkLbqaaa93+eEoHYi6hJTI0z8n
l6dfWKCS6hfAG6pQiNw/+VjbQWhQ0pEN009Qa4LVq8wwlS012jDFRxh6Q6mk7Wrx
en4WmzVlx98ypegsK8aBt1paqRSeOU02m35w5m8nNog/mGDUow0MNmfXKJrlAQbv
Uxvc+PGYccklSMyGL2HeIA89/tdo8Yx8W8Tm0MIvw+0wpjah4OMuhzaNt7yp51Nt
IdHLpaU6osnLZV/oJTBcAsv+/APi/zSDplFyvtCgfl2TjYyrwGHHYYhSYJUF6waG
GwGZGZqyGTt3F4m5/O+XHu3iSTDVL72yFs/d7p/tamoujg6IsPdeb6EXwQmlwOo9
kiC4nfZprsGt8wQ5i6+jll0FWX+fQkdk6XIu/QJxuqXfxRzSl7CzsOFVKdpZY7pm
0pUGlmSPcanvCpJa4IRaOXUjBzr0s2xKJBmzG45+1kmqJi63uie894ZUE/fELsAW
XqHuDNND0PHzYTiF2FgTJhrYg7WRfNHYV3HEWTfiinnqafPM8OMBP5ha8ZLqRW3H
GfYpW5UBBObnYzf/nCs0Eux+mpVKeQRFPacaFn9aXa01kaHSjMNjECGmb/p1yGiE
jQIXsEa66+/1cPnSVokt0zTnsxUOGxr2E2PYfDbn3SYB5R3agOLtrbVJk+Ymjdj3
bzXf2hoaK1/yBMsXz/Dh60HL+HJWjbwzsBjo6Y9GMGGj2QmHk464eiPHqQqM7Tuj
WMGbuFJa8HTABC2hCTdKlri4vpWP3K/qx8D/MTriMI+4K2T69aV6eJwCED2LPGCL
4Ml77khczIBnE8gr3300/JwC8ZOt95oEDI9iEVRjIUkwy2IendyxHxB3mKuegKQL
7qCqQUtUi6NIitpnfI1SyAi9Ltab2HqeUrwolXlPz5JTKGvcSG3vYgaZfGMzkR83
lzncqSTfbVI1E6r16gZD9jWvNGR3ynRyPiQzsrqfRC6VHZdr0h0wf/T3X8CUr4is
nHhEAlB29Yd6YOPKBGCmduyt6jgHdgsWmoHH4+gnNYzKkWsjpKdy6qc4RcpFpHcm
AP2vuPx9boDDGXPpGTycM2yvzp7aChXZE4VDIIIM77aB2Gyks2SAfZrdLgi5ln/b
wC4jV5eloyLAvt2JtL55V0+dxKfJLPslwMaIZkWy7Zak11YdlFMyHKKIilRvAjoP
FvyEk2NqfI5O69eSgsPEAe5Hmp3icDbH0shEnxY+psYOrD/5f2axjt8DgxoszefK
MFvkTJKQ+vqq2QGHrNjPKTy50wBQNWsZkOuCLoCOUZZEs3aPeY4n7qB4rKJzq0DV
453Zpwo/oZzxltyc3eG3I/4elWRgUHvDKAMWehFiPIEM4OpH5vFqek7/tc0CP9C9
IPsseffShKXNtI/z+vJx8jBTGgNUZglC0bFHmOSuyV25k6ZcqgGC6pks+6ysA6RY
0Ngyz1GWPwdkk7z0vN859HYVd5URK2wcWXJoB7i7eKJLa5qWUHicIY5ympJy5H5m
lEXhlTAxc6UzGAJoBG+PhuVLncQQgrzW+IA0p3wf0a2KEPzjWDIxFOcHXHs55o6T
+rx4ZpuQR7h9dS2K1+cbRw6ZiheyDmDDEPRBUxYkKQ1sG5IqIq7l8YDfyDgoiTMy
5t2UOzS87hpTxxOCMX4qt4Pe7CFGHuy8nGO28zaU3IWgXoNA72s1ugpZInNYh6v3
YasLIDlUKkpB6ESo+MKd/YKhuMeGgrKIVbjg0W/FsEtRs3Mj7b4IKxKo+OYVSYSj
aMLcdavNLJmO2Mgt9FQc97rD/EQMkY8fVtorcGZoMcCgescmReJRlE/dpqky3mO3
O4LK2nqGw5WKfP6NL/WuZTGym8JVHTtEmuw5LA98HVwZrSXArBKxY7y4wRcNhqyA
RjPBXdY/WUFC/CzkWlqUe+nOgI9HrKZC6y2NucwMk4o2u+dyYanGXYtgiIJJhbKl
BFnruFEE07UU1K6PodLJu22p911DwXrjmAtaQBc1KY+swkOR2qoGEz0pkdZ6a+17
2dVUnp2BYUbYlfiXlJqDDj1NavBCSz5onbQlhPmRAEIXxKldZ9m+F3xJAk4S3pu0
sqGQ60s2syjOiRGsuK5TaBd1JZ+xsZx1C6SoDOyoqiEmQKEQLZP7L0FFDzisT2BK
IOqECbXByA5i0F8bKmHRtCjhc9GuWO+syf3RpZ68Ev19XKN2ylmEwxSk9pGUB0zx
tFMcreiNJIbCbznYkSF50MynuPlIPDgdcomw8u+QUNdsl4FjUNRHZbDBvhIRb+D/
x/VY1xP9NPDl+Q7st51oqu2dtlp+f4sJoBpig1v/sjjqv4HtPVh9xY5OZrJIwWp5
0tUQY5gsjrKXZVtuKrMzjF2Om+f7nUBGn07XsXlMPT4HvGeve7sA/J/VpE9CdEQz
8sBIkwMuLF6rPCU65yoDYapKbsBpAp4F0HsRMVZlADwOGVReOcKz0mr70acbKbD3
chIOaw8P/GPo/EksVPGNsu8MFf0lHtKTtd6+Ti+IDxp3t1e/VhIFwJ6IQEqpt+Et
nKTmkYsUHbLzbMt0Z9F8o7sgd2R0QEocpLxCgGcxsBNILrYfKTi1zTdtRo6X603D
NWX4pUR/cF3lNaxV6aSPYEolOBYsItSpnfJ+qTwodkQMKtvUOhzky4h2KhVkV1/g
JQMUuvpa8KrjDP4yNjcehPwEceOPHEmStgKZ/S8DVjwhjCm5BwGCf1zWCmplcwXP
LoMKUg7g2QLE+8A9cGFcFc7yLim5psrK+t6stdHEI6iSMYQC1GGOxg+o13v1eQpa
FWmGWfihvG85nqfNRRuxTPe8Ttc2vw40Tw6XGHLv4eq1h/PvBZbj+EH9hD0xDv4q
kF1HUUOWBv+0QMUiGiPhLEbXwDm9aapa9JeTou6VPQNP4SIKJh/hzQGVWte2G70c
IyffJ98S7jfu6JBAf4vwEoGszEwO4sOHNbexH9JhFX+EHVV/Ro0SuI28f9yXXdJ3
9yq7hjfZtN/KwFwyRHXjg0Gw9fvXunO8SWQNMw8EcJs2T2zalWfjcky6QY6yf6P+
3mEZx+0B7aTK8qCtA7AVpXjuoVc3of+QOaa5kLZpifKP+53WDo9/PQ8n1t4W7gKU
Aob/R51b9hfhUihBnoolFe8FX+6a5gGwHKrASSwtxzkzT690wLdS+xfgB9Vxib11
3FzX9lXEPoeWeZO06Y5u6gr18faWPHbD2DkiumCSPqywkBcUqyZD0fC2NCjL8b+c
C0e3AydBeuvNdSBsNJRz/A3vRSy8NUwcX3FLrUXka51YS+BEJ6BsImZnJZJpZ2K5
GegGV4GbN3gkJCjP624DcNu6b/0zcGoPjh14lcAAJtfHe89vjezqIYs6UuU9zz3K
f9F7p45tT8lPWyavKQj5aWj03+WF5nmAlqZfFz/ZPt//Jued4pJ8pdCXbWJwEYjO
Ee6I9WZjJwxsYVtT9LykYhhYsVrIFCA1buoOnlTR0fyIG5+rra3PiHaYw6WAXhZD
xIWlxJvINTaP3pCiZkyVYpgy/7xtZb9HfEtZZdulMVSHvAzZ6IDO8zddVPAKlylP
J4vVefirdadS8vzEsMupNQQb6pgnXy78Qp8EOVgxIWvB63bZH+VE+SqRjxAqx2jx
7S5XPUABB+hCUvUw5NIrEWmtCIeUwjKH0xg0Ibe6viEJboqRuVrOULCRE8GP+yZu
hrRN2AS8U4f8br4FU5yKBRo2zJK8NTktlLSk+rHZ4yHzZ9QwpTXR3ngP7sMHzigP
9McrxsF+qRMHcIQEMeqg8SGokaRlyzEqfMIU1J8F6Vh27bc+3h6cZDfyhP11tDns
vFjhMGZw5XnzR0qyjxTGbM92Nqu1cPYOmpMMXnUdBADsCnQogYJAyYwgmoG3ZZdD
80WGgw4kK07L4hMkJDTOdVTPFdJ6aoSrhN28Flt77lyZgSiQniqSw2vUHuuek/18
+QG2TrPKC9F04z0xWRqt1oHSIJuliUq40s9Cd6ZhPqYR6zXr6zlM1xhxrQsYweyz
8curaUsvFNmGGCpkbdaDZDiVCHbDkrnEC9//rqPYzLwg0ezUulT0duKxanGOboYi
ras3l3gkE3x+dB7v0ny70i9IxSELfEOt7vMm11V9ObhyRbBKcGyojHeR6QuwZp6i
S5zCkLxbc7eYCNQA1quPMCBxiQYhuYarvskegai6VmRno81OCtpUeSkuF+hutUQQ
CDORPxGuKj0ADfAFlFgq0guNhBocG3TVI80kCfcQeN4zLf5c0lKccC4hFTFv51tO
p6zB2cOoTPe3roovUv401XiwEz3I2o15Py/xPQAJD2f2YEy8bVoPUHs/OQHoGs4y
nXvd1m+/W+JDnJhAg5R4kzURsmIeJfcx9OeVIGMc/Yl6c6ihsvHonzvZ8D/S9qj4
uGsbqQ35cqHbALqWOMYdG4r3btQoQfW1ffoKjlMA/0Uh2iciNh0OoeuWlX3zdNM6
UtYaUm3XqQQqGk73giXMzcsMKyEVbn/zFDxmjVYvBlVRPKx8OjMRgBCM0jv51z9t
0W8gwGBGXBcDzs0RY032nkA1Q1jcdkHH8GSWFdptT3bPERyv+pP9TZUzBWzY2DS8
djjGjf6+u35VAYuw8lXHxHyLeuEj008dk9P7Ka4k8yVVYWwK0YeO+55KeL5uIQfm
lAVlsCQebNftl1U1r2ifAbueJ7hUOy+JKkrYk2gx82jpFgG0aJlw6B+1Zf5OWL8z
cbl4FSq2QlA7d6o2+inlOTrL2XN9BJJrD2wqyDWtYU5cKKJMIp3NvVbww72UF37d
Wo7m6xjlawapumViqfYRoq8ikJ7sDFCFD9AzsiBpmdUoVW9FDARvCQvMQ8xLdjai
hM4EPaSPUoUD/31TfnjAtQi/bCtzAvWLcX6W/+4IvQOEojpWmxlb2mJzvtUw/dGL
+P7u7C01H6UPklcyZ8NcXLN+zX4NJeaklAm13RUGDt/BwRRJfa4baA5nT7ge6/Hr
kKifYb118LH4lAIvi7iLSFomy/V5+QwkbDWu/SxuCqzVFRmoBIxKCFiTq1HTfy5w
YuH/5prwjrsycMyIHpVTthhXt0N6C24Lz8b1HLhFY4cyl98dIWJ2ZXjBIyqZCb2m
g+n089h8OA5sntoM1Ba3e5aTF+8L+OzwVsYRfuMIm2BWsY5FjqTWEAJ5pXhRF0wh
aDF/nFUIMqJYP4G2edxfCIVjFfi1CQEeUN3CXaU4pjSq0+tVvmgjVra7sQ10q98w
YrOfq0jE12f2VoJgLuadf2cGLhUY4yruX0SuMP5ZpWYcIlWCgqhvfoSW1vJwSGKw
5BeNmSQQk8oN70Rvkwa3+v1Dknne4X8b3rNv6nIGIUG0Q+YCjdQCnyXdkPWAADrs
7OQAsOLZlEZR2g4a78uArjhWXpW10o54TVnweSyBEFDx9w1dJDxUnugRxLSUVkdJ
O9/PtLioJYT6RCdKq7+014kctDxlPszT23aZSmR1cAz4JPxbrsOt4zDaho92H51v
Ka6X3OaYYqNG8bvALrcyN8JHWDoL/0DTbEKK0sptbQHAERVODfsw56YCbpaqWoPP
ZnlcG7x+O9sYPhyt4wRCUlFBYsUH2S0zJ5cdthrVxixzSmwR78rN2YIxoPO15Esr
dZHqW0uNHHa3hVb73UJQKViRe2eowHi2F4HN5VazmI+X5FJXUq8+Ur0+qLn5SS3W
Ldt2RGpbfEfm4AqDMwAb8Po5ACO1B1fMF5DuyiwErU5Ez3oW/jxBndYg/0mkZabX
jhkdTTkvdzt2ArEGxZT4na5B7jhV6yFX8wc97BqbS5bvyHGPGIUKJTfjTbsv0E98
uJ/0m1KoJU9gUvHI7UsFhnGcOq/wqCvTO9DlUdGz01xuNkZ2n9ZZBYZ8nU1Edc6F
FWguXtvFczRcIfSUpQ/9J47Ggy5a6C1jCCDNbWbf0bjav0qWC5IZAwi+eR+eTpIE
0ZFs4ooYjlB0qCE4HZfv/F3+pbl1yzpFxCi7y4IjvJh44Dw25hJjn26lN/ZOTFvu
Ah6hWP2PEni869jmXfeWB5hSRKM5pjpXPqiQ6m0x7fa/aSiQ5Qi9GWP6z1/4jIAE
xCWJ4NUA0sz3/ZefsxaYCvDhJ5U2mCtGexmbb9n7moP6sb9BaYCPHHHyd7HO0l8F
AWbXZ2Usi0Z83K3UUsvQYQZXRE/XC/uCDcrJ3R3i7EzCjF0R1w5xgdVXCQDD1vyd
WWBQs+p7K3h9mIgbGqwhqcvyX2UqG6HgMnEZtOC7eg3AiY4w0vCtD5nUTDrFAX9u
HOn1RmMF854/t2EqMWBY2eYBUB4CmjQ06CN9D3JOHETptKOgQ4RNIR6rQW3NmkHv
BesIwdc0iFoS84+IFySyzQds/NPEQDB7OjeGaYczB2QEgRfIjm76v4LPQpOolT3A
VHKitda194GHWOgNyXmeV/mlE+XEdlO6Ijr5PB6bZAnvDHnnVP22m9P9chuzu99e
k3wO8/DAxobOu1BmWHd3BSzux5ZoLSUJeLf3POjDoOOoAer+W6e0PQoAi4dZ9NIz
VSftBAECYJBqmRIw+Vkv8GePWq4EclogH3gV79KxgC9rGADS5yfJmmV7zvnKXH6u
OwGwai84hLGeBuLDKK1osh/6znXFgMlqJqfWoFjpzNfsZafwo9V8e3RXzLVcm1Mk
mvQabORDwa36slbBomnSsVHTr+7VvBPtzYyNbnA3fj1oA1u0usncpM3NMD2iyX0l
77JmiZ4isBCgBcTQ9qE5bdG9LKd//CDtpfGDwRq5jXdaezRaOdx6m64m3ujOtjtR
jKAMAtrBhAXXyAORJPlh4kyvJqW0BJq1zA2R64F5OMVmfjXr9WXf1ikURCeuaRyr
Ifxv12ixfuLHwZu010ANgI6bDB+XM1Sq9xn93QjZ7DDeikCLOBI6mf+E5GginE9I
nAN8Z3ebJYC4d/3oFLS5GsPMl/0TGNLDZJQs6tsre5CZUAXu+zg5uXGnkWRo/wiC
5a94n2rC9PAPiAotvWchhQb8yDyOUZQrIDjtlCD0/b7vxZa6drMWPaG5S3IJjBnV
tmtA86qhZ18EDMrE1kjcHCoEJYlJFqLMAnYpYha4RUOgp5TI7Jt/9evXANz0AeTA
Xg0YyDHwVMwz2Ksi7EnBCRwbZc5nlV5X5lhNtgeD6VZ/YQeJVTIGqhIDYPweuTZz
ubIWhfASRwj0Lgek8pYTvLrcq4wXcqlWCvIYVibUmB8/WoPlxL/HqY/1Xy5Lp1rW
lVjdJ76JefTKjMZO2NfiFOEAjF4tXajqreNBv26SonS5E7fcc66rrH4F9krQDtyE
nDmrLoCde37V9BSv3/oNwSE1hC0LKwC1ojkaI/I0qOR3HEZm1vkoadVfTpDfSkQh
3624hdjDAPxtSXZR4XR4eU811gx37ETIpbsnAkvhgrlYfyUt86jfLqrZqDBeoF4e
A19FVrrys543qZcnUAyF7IU5MTDriN9WZTYilH9IxsKklAheIN8lEecERCzgLfYx
NbTOkoiuy9Gq0AqIPyDRGE3tma30xevwj/oo+noOF5PbMnjVf2nzZr+zIjifMBHV
vyjT3X8g2GTtmWVqVirg8F0L+4zao1ClkYQAOdAowk2DbQWhZ9mfR8TxbaGNJ+Bh
Ddy+6XSQ1awK3wQLvvopOLfLClfBwG/5GbxxPIhOWP77V2UVDiEZO/utzEf1BCf0
WaoWZtWM21iq07TwSEq93sHiKctBTqdGI8N+4KO1ilEwSRATI0nKuzEvRzCTPXPd
HwyoThAmSuPIzdaavdM3dRcKloOzMQIwUiLvHW+5u/YOurGQdjxpxj8pJ1PEvo93
H/LromjSwePQTTxOq4oWkyC3UzXg+mcr3y0vvhiUW9neUer507ikXBUPpwXHk0eg
rLKh0ZO+d5GOLNRQU/co6swhayaPEDuJ7mPL1PSyZSWYS03lRl1Nq7OIoP9tuPLx
zkFez49IPpjicwFp2oX0c1DI9D6hlDXgZKC/okYg3yg0b9eNGfTRyE2ZsiGSqhEn
yZlN37iD7YyzJylBQiWg0v4Jf5PjLI4shwUZ838zQBVQzYblWfqePZUo+b9sCmav
xnJDoyfDwtXg/bf94k7QruvG+rgtUhtr2Kh3rTHV+XgIcYN2Z8ZqnNs4KmWKXFzU
Pr+BpRSukn/Fym/v+XnNTE/XQdSsa8J8zZmoDlotXgdWaYX/bbob3mv0KNiS0lue
nFVMxc37QpMZfu+kbKGZo4r2gkkLxasbCt2dpdREVpOOoxI+o41Ggwd6dk5Oi71/
bLuTQq0z72Iy6uwkl90fusnpJTTB+ZFK5OiRS6kIkurjocntg0Ypswsl5npKfRYr
5QX3Sg0UOMntrUIJ03A0hExRRsiEyUSr37Bur9sYQYjku4oiHIjNIRMtGTvzcQE4
rr2w+BfowxwJ3+H7cx9n51z1r6iBxK+/t/oSTzCZaDQdxIGSdw9OBt4sRPQy4m4P
77myx8FIn6OUWz+5IUxo7JSsKDwqTqoWCrGtxfvvKiAT/NIbyZCwYNlpmWB5Qag+
wYgvHpffkhalj1QKPtXWzYYTrXfgcbjl/GmpG4uqi3lI4Zw8RRS3Aaxqbn6MLItD
/VYqSSuNSzkexqbRYDPcXRnhM+LCplpEObgWqDvuqFnx5l4006DCc/UJId3oHA32
Wkr11tkXWRBe6CvPBZaW8HfrQcBYzeRA3aHcbcrjJks8+nTQaef+U8rf4CkJaoP/
JusdBu73goHQxGiSh/egpZtFTPpvH2Ihfy9+Y/u2CYmJA42nuE1fVE6m0uDVFnB4
BPd9d3iXVwevJ4AeWDhEmFCNAUZB5W9SgSueY7ZZ/ZbtEkAWXHeu32oiwrfWgJcA
ooUD4CknK51hhavrCOr6ufFJeH/+Qny7hqZo0Qa2c4ABZL1lkfd02j8q5yEfG/vL
TGuK86mncNagRsZHsLGmo6GfgKLDF1lcFHAtmfXcGhXz519EbwwpIDyVwpFod3H0
kDAZrzU/icdVotth8WqnA+UEbsB3a3xd42ju2ARg6quiZ0DdZvKozJnazM8iYOQY
13LuwiCvAiOL1mrgCs7gVyRiuULT1veKJ2Eu/8f1QqtouhshoUAa39gwDMxL6+Ad
VoaxqN7T+dZ2nfx18ZKPTAOUQI0V8r/EMKhwOeqHgz0TtG0tzUqw6XUgZ/9q81aF
WQEjJmUBt0+9igENw5t+JAKgRT3uHOO2aCCNHaXOso0lzi7oQImfdqcHYQcHgx1l
UyFomC7/9f8/EnM48IXTuGn9ZZpdTsLmAJQysY45M+V1FZEaj+XMWQCum45pELTn
qquZYLGFxFC4ah1GcABld4/HswryrYPGN/sUh9iET8d2Njl6CCu0VZ6FG3nDe/hD
CYqmfXbH4hj34TiGU+EDjbyEU8ZTJwpHEc67zP8YFdNxvdaRfmqUFyL0FgfY2ke0
lQoPYFZMU+q9XUGa/VvwXRSV89PWKIadlOpd/8sEm64CeeOBf9DPT5Vsx54QkmQg
gcmLe3vFSdH6a9tqH+syGdwRM6SRzfIvygXiRH5ntr0qXJp77Yy3xGwLAT78yQUg
Y8aIhZGXo3kAX1IsTuCPIn37Kj3CIP41LPJNU+YSP0pPP5gTNNGub2RnZGaAGJq+
6Yt1ckd5ZD82gKC8WWMvF256O3JEbPhSVFRAsiaJgntQkM6c2tUeHwep7VnXeP7I
LsnMKooqU49FRTl3Im1GTVu9+pl4v1nZ/FAVmpE0ylmVmgBEK9rYGZ0z0f9x1HmJ
tJOFBY3vxy2qyW6pueu0/KJYgfaYv4sxZpkshKJ4/SjjMomNtDzA7C/FkHA5ue0p
2mscqae4jA1jzB4p3lxZ3WDDi2bve1mjw3+wUZydgAwTyU6dEGWDEzfXyQAaZihO
4o/KBcnoHg48bLlUexdq9W3hz4CQXxtlFLBhD3yEYn/8b7gNwEJDyzBTyqnwej6v
RjPGkukmqfuH3DSlRtaDwerW8sfZkN8Iu30MKUpWyfjKqtoso+qXKqbYIx/a3aYk
qXDKcIw4b/Sm/D7MeEpNq50Q70Y04EyIO4WIozwQCxt+EAO16fV4ttjypFKklx2C
XZVySwjcTq0k2WMwo1JcIrKrHJD2Mt5S20UTiHN65iNPY1TYt+vA8YokRmZBy+Ns
TWlNcq+FVV/qrcE/kFD6xkErrXm0vfw7jj8WEczXGEKu6BFpdfxYGoDtGwMg4bHi
d14Yn55rChp/c5TlHxzeGrG24reX7Qk61hdYm39T3nbvFAAibC4hVFz1kCbNnnD0
jDJXPmnxOKkXXbKCrubKaoYbcoCNUHoP7FSDRJJMUwA+RWI2wwdahFYw+OKEm79h
bIzbVoMK665lpdcYYC2iZ3zsSWbDIDBcIEKo4T9X1nAA8eAzQTim8MJqszjJO5Jn
3FQtAqQVmcGzcIjGzu/UeHqvGaQTOxctYNxU60CdWPc/kMnRPUmoV7C0Tel0EL28
SjfyOfM3/zh9wqzhuaHb/aAoOs6NEObxQtLfjY2+RwAhxyhuiIw2oHuK7aDstegm
nJkvHS7qV9UAYqVvtPvNu0SsLy1Rpa5uQfnXVkPPCoaMP8SAvTY9JeqN9BLpK82v
IPos8unOa8d+rWflBm/rFaA1NuhFFr7KpptipHH+rC4HmQEluHmMmNLQvdcP8zXe
xyfmCGmoJEfl+0QJLW2e3uEmxrpcnf4eDHjyy81dElg4ZiQuSdtvbuAe81vOw7kG
Y6+WNcyGGetI0zCTafQxM6YuibUOsgJp//oEKfb2PAECGW9s/1FnCVaFzAjQ7X5l
SU4zmFoG87u0Jte2V7uicpG5Iv92mWNNt8LVUlftf70ea9cULZHIPqKHBit/AY0m
FgJ5YIRH8R8/wTE3teR1vzPQb5cBRWfaLZCM8bzCnhXeotEKzFwCB38qm8JRhc+o
x5VOg+U++mW/6f8ZaqJzSmwLbEoZvOeYbjf9NEHTBotgwD8/lS3jv2JmQv3myoOx
EGPuzRlPFVKUlLl5PPFNlgjkJaKaNfrVBFJtGwseNN595OpyRj3VuXnzwqBfGezj
i68d2VEprfnyN9xJ2iVE9iu2Si5/5p8AgLgVa3LGzi0t96qkdOD51qxI0Y22ZgaX
TwtBAPACKT8vBuNe9TTNdQBjOLhcGYXNRrLiHiWEaRxSEGvCrw29P3MgyNFi6uoJ
A9u4JqZr9BwM66oKvp9v7yut+3bBBpNrB3/Bfly6AQg3VPCRwnhKAfek1sgHqUGG
erIO/0EIJu4N8R2gUqVsXV4J+R5EVQEG1wKNAYVhqWtOXMqqzGbcOQ08YCyqwfmU
mPU4xKF2B3+HtFApXIMFpiN7/WGdfEZ81UEYaeyMLOo61g/ka88UYQ5B95e50SvC
VRpB8lJLT8Etm4T5BheOW7iA8gIajfvPc4bi1Cwjh2eQv/Ee4wMU2ng9xP/8ioZl
zyvGKgkn2vy/JIFQZXomriUcTWLMEvqtHbkk0vv/fgvtZrD8IlGlZrsUNHGSsjGq
MOstYp9OJYiI6wsYaONGn5LxJ3iivj/UfO6xKPEdS9XymYrvxm+IEg1VL/87RggP
qOvEX0tNM1YyT4g/xCb9ElzxF6+9nnP0R9iK2IjT/jCKlnYL8Dz1O102P2ATO5EG
R4eQjM51JnkhxYEICVTnNNADI+cvp+acWg0QiXQAhnQPPIEM0gLtIBQm0em12+5n
lwjtPz8/tQemq7mQBhsBioDOYaS5eB57UE7rcFvDL/ACI9PtbYMbewQeaz4SG+wr
bTsR4lOPckR2Xn7ManrJqhv/tSMOdS7GNlWYWkyjBflU+7VC5Qn68b9GAPmND+vK
MuWDpshl/jt1ZnxdLSnwQFjTBheEnpXDBOn1puqzREVAx4bx98hygPKcD1VIEGvT
+F4QWfHD0du4McK9onaq+pCbdxcnLXk3EgJVjyj4Hl2eTAgL1vxlkhVHIplExPOn
AZOUU+5jFWAhPcPLefQRpFDbNsGSx1N/SZ0cOuUCRnusUcx4wu7N/LGCkjK2pdiQ
IRC4jqIRzDg02U0aVsOLrkQLDn3DgDKIRILoA9v1bnUSpq97uh0uEp9fV6AB9TZU
cdpkwKt5TraX4TInq4Osg5JhUdwyD4jUg9AUUPp/SVcwRnGsfMK/Ks4Z2i4URzso
e04WSqLTeZSIMpd7QHkAc4LAAHOtMJBHg2XNYhHtjRKifhAqvdahFFqOx1jPIQ4r
7gbQDbKNqxdRvQSBaGZEqNuq4WMWZ9VPtbYItp3xM1FmKoVSSnqQfZhjRrNQydlJ
/GwPKZYPSBcQ/8r0zD41mPAJBap+wCgY2+LUlRNdxI9mYXMeRyeWO8Kfc2TowaLb
zhcClBIb+hrBMMeqhqsqj7lDijn36IdU3dGRJeCgTIF74oxGBJULnee/XNBl7GxG
nXYB5m2IGkio+4pmdbKLRGGBsgua/b7DP+52DKxKBNkeJjs8qcZqaKE9ar3SAt5a
ysK0Ef5aEQa3BoSIN5tCCdNmXtHpsBcwbfxHK64Yz+sgCPwVHfndsGwUDbgFXm9z
uHXtc4yBsPokroPFw19FEl6neg7AE8TUv9SQYWEGUNCX8oJUCcJaMVw1NVD1alU0
lFDGznwkiF4GQySkP4Iir9CBXNdukYgP2O3nw9+ImsRCcsmBxOXT2AgEOJc8cDlj
YsXcj8jKrOTmINSsxYLx08h8IOKQTTviXQu3nePKLrW8AwZr0ep13skBWtJzkC/L
Qk7iDobFJlrA4R7hKdaS91EnjGsiygXHqNbjXFcBoQV/LkM1Dajk5i7ylx9MQ92b
QXCunYK53iZUumeCw5pgFxxL0MV/MfECF+YWICZfHlqitV6h/7QDaBCkm6ZUDYxP
MTp3c4Ax4Elxe6ORwvvEvZYxpTl+0WdRh57+hDyHVOwBchqc5NCjYKHwUwKHkiE4
r7B2BYkh7sWoO6LSQ35GaGuupj/3bc97PpiGTeMeNRAFcVzFxveC0hlZXsk4lA0g
N3eOaWzKZBJPgeFOY+CkF/ldpgwNvf1ufijGl1KkMkYKvwdBIWS1dxvHrDpBWe+z
h1nnpU0XvZDOz1diE0eW5JoNVzDqTy+W8WpjwpydF2h+LoG3qXm4kDbkWVs4QD/U
xz0cHhlo/hlSVAi7ZBdo3pFV2lChB+a3O/KSwXBaJ0oM4pRfFNL3x/SVfQymLYo1
eZkPbX2BhCCnYE0z32Ht8eHqcsUV3GAEg4cRXSH+/Ou/616dAEZfktMrmuUl0m9f
8q0dufJThV1aP8XsDNt36vAku4fmKpfNEmy8kroIpayJ8u9LrkeyJN/DIuFIDzF5
56ygbUitSoZbgoImcW8X0T6Ke7rf2DnsWtqHiUYAP0PNjNBLgC+F1CSsNoqB7RWx
xlQWCpHHv0Uzq1O8uat0DE+tav1lyqgAK3k0yiaCxkdlznPxf63B0I7m0v2HK/6B
7onJReTtF1cLpRvGRPGjzDFdYw0dZiza7mpAxJ3qAHlAk7uB87/wd2iyf2ZiCo+S
OP9kR3nHsg0eJGii4T4JguzVmiRsqmHvlRCQQET39AFFUc4pIr/LjB2S0arIwc4K
hPyrdrIExri/UwTbgnouaVAjxnCV/pipRqvaHXLCkVAiK3uQf84UlXzNT5AAk5a9
yhZ4zk86bXI5qChMVy/7TmZnjQubIOMRR0CyjYddN77rTn5jYpIc1/FW9bXm8AB5
M7Iw4j902BJ3YF6t7xSyCEGLTbUIyIVAnSycjCFShPix1ZdYWK1KKK4p8wlhraEi
m4JO1n2Xewhea50UlOQbFj0zQIyfjsh7RWg3nCTn1Nkl1YK5sfyfGhsaFaTffNqa
RCJ2xcHJq48pWC3UN6q50ZXqdxbnjuNyKsA4EZvh+j6CNDcTKgdSaCvAqa83vF1t
M3Yco1XRJodCxFeGO313o1PqP4Il6ZfEfy8FIrsFDowzEzWsxkHeOQ3xFzuNEm6O
H9bWVQ+qXWKGF89xYTrbJZO5hVCUw+GtQqpsuA6HRBG4uJMRALfNSGlS867Fp3O0
0MRRdc42HJNrOgcpKHL7BAHnBWkX1qaiNk5T78bFPxo5mh2ySli22JIHS2b4cD/b
V+dHXy9+eVgSjUPkl9hGctDSvghjMYtyNZOo73UZ37MokPp/VACZxi8HhM1x3VU9
9h1mKCWxAimReocDz2TyVc8B0vQGcmGacZp2TQW5Ngm5h9mRRLfkMMwTNoexexdP
fS9hDV3Ygs3tuGuIQJOmAI+p/+KaqdytiQJnSYf8x0UIvKz8XubyllnWCMy9J1tJ
lqCk536VahZ+QQ5VYbgWG2UR5xLgtSp+rmiqBE2EXK6ttAW/KIdA1a8ebhqNX6bV
AEVExZmoCI6gzxxTyk8+eYiSTpzhyeUrsLfpN960zZdWV6b2u1qjVwsOIeSH/Czx
nWy5izxUm1jD7wnf3xDgZCF7vimjJ1bkD+wIwd7LzBJXmCTfYYCE9bnT5CFIr18d
qmJbSvk1wHZYYi9KFdqjmh02JWxaKwYEWjw1kCBD6kvLn7ydYrDqAi4KS9Q7tEMV
6gqeo3xtWFds14A32FElSpESMDiDBjrkJYeeXGyWEud2JPa6fX83ylRxsIl1PgqV
j4ANMWMqcozOUTyLKcYRvoOPjC2lQ4/RXZ2kEfUmxqQfPyXHdtqd2n4KTUIg7pxd
dzgLIPEXmeiD2x0+bl0LPhCw09PDyDNvOMjd/UuYnRQ7k+/CYCmf0aYqbY+8sVsU
7WE4XQbaTpJJY/8m5oLCeDJ3H6sxHuJVaNUmvt5HMIsl6ufpGn/fWytJwm/awUuK
xmfAwn1LuO41uhDB5cF5O16+RAW3pd6/qCN+6WqbAbraDNZWqrbh27T87/eAPDgt
R9Q7cWB5SRqemQ/DCwelCH9Usm3YIilULlllhPTpV5HIRTCFt7JXc92GZisw8HYc
+4aEwLZFk5cBmPxyrK8fYXDoZ7nSScpRPIjZqUQbt6ThrwfduLfPzVo1Y+TR5h0l
0iiCaJsE/iMiKxPSGbAPn2vnb3hZdjvWTaHkLHgYAdfz0ribZYfZMKkEh1YjlA3k
NnW0t9Z684HmDsRI3cCceWzij+wrACtVDscyVGT2lhwF7Zwoq+/X/EZxZ31F1yHg
7vop46fT2kOSMkzRz62eEc06YfEZ81c/wbGIuWthpaRiYuWGz5OhQErALI5cYxtz
rBn3JtQWla6f1q8fwB17XM82z4cYY8Lpw28nZtAmTepnr2YrIhrnt0a9PDv7cGDW
123zRxOHHBdBYy9E0BC4GN5zChJ4GO+JYeNfgONgP39FACKgvZ13H+KLfKoTLLEo
gayYv4tblCUZ7PjLfxPZBBZFlOKGtCBFpQu4PFHZur0USzxiTwSbyb1gEyW5RorH
TuordCm0xdcGH3ZCIIxsSabaqaTDkynVP3Bz7A50Wbbuh4H/SWwrj5H1JpVLzRWM
xEHfUGo3gD5oDxq/1mtY7GMfVJqL3QBbJbiq11qNiHXyWeJpSCGqRLL/E9s0hrQL
qfus/7joYIGYQ18hdqHaKaunC5lT4oV7QeBQeQvoaz6l0ro50bMl2+//5jGK2x+F
E/B6EDGDV/xNSAPhZEElEuZZA02mPV6eEbQ/Sn711j3Van2ncw1HBp7/dSyWUYIH
n0cyyy5soZbZ1cleselpnRCo9Xl6ih1iH3j3/PySa3YfUZqmg8xYGmQeaYMTfRhy
FvjuLc//e87Hn9iWc2DIeMc9qK70lVsR3q9zQlOmPSjKBHk4L5r8dYQHzEsp1lDg
vUuRGW3Iz3AW7+dYUjSoc8kKKc9kONmraOSck6p8yuHGW44mteeVkXtHaXsmDbtN
4iD8/k6FHGNGifldCdSx2JqGbsiBRLKdfDwPjUsg8rNeMAzhbCakpxGoPLtOrZp0
dOLNVTGqKB+w8t3FgN7yvwxznazEM5reccffkYbH4SVXOLKja6FFu7PRGV1j2YmL
mzzVKeLcCGf+PIxvegbFa2WkoBYdji4ZU1a3IPsKCfr5I5ZbTyH/iATAXWIwYRgb
e+TlsT9sbIYEbRAotXYNqSmmikDv0KckoCaoShThWNhNicC7UijCXd2X9IOM9L3G
ZJZnerV1d1fe8IDUeIibNW0/Y6FHxhCmEA2+Tvu7kt7oXZJkKXsmhvXm7/Gzp3ia
xG138XcwZXVoKY8einKPcE429dYBwegGr6VeXet2+kw22jIfz3Px3+aR1U1WzPfj
PO2xkldo0p1NR3Td4yOdDIL/3MC5CaiWKTLoih8/bM9d+gFrVKJr2Z78dkXlkU9V
JLLczwk6kqnHFDQzqCdPVl5myhAYU+c8RQ1QUii0uV0Kcu1OmnSwVFJpGU3vxJ7V
L/1zACS0W8Gv99hHhZw3voBnGgLr1GYbxaPOkDgXJnd1Cest0KVmEtIFOyjICDNE
Co8JlTZvoGcomiuT5smPYs+Waag6I58+dJEXI36bCrEBAoGna5zJXU/hinyN0las
uUjDCyPwIBH6XU2wa9DTgwRZItlCrKzjYC9oRrNvEMuouD0R+5poivqASb3+l8rV
l/NQHZhpSyz4dx2L7h54YOYSNdS9eZXlDDB5fVLvGgtcE8T1XyGdhlLsjp5ISLRC
WbXA1Z877EXTlIlMQ6VeLYGrlQ6ziin2gqtmErjNomw2VJqa/H3WZfHkryWRUCW/
bJqPSoMHUx70LubFwzx3hjbN3xvSKJ/+8maqjFA+2MalwEGXsHkg4riOSeP70IAh
PiH8hb13UsyouhDTMXOLrcONFdqg+Lz8+r/mKcIzBGGxDccCYUag2qAfn2dyXnSr
uec59KuMixr1fLewpex5/J0h2fqpUbRfY5dYal2DwKWrMuFC5Rqn9ppozJOHWV+U
m8uP4gnQLNuSFbTmsUf0Z5MFxyR4sX6C4gnsE8SU6UXD93vF4xtcInosNYb3hNwO
vlfJNtIekx0AL6rJUgwcT2uYPpD0KOIdVIaILdBCMNVd1VaDeXdXsX0D9tuL+QST
T0fTZkgGL4vKrxTdo/izM/ojYY/I7sUu8JI+823XfFwYzT069ye/qBSkisdSuaYo
mfZOIJiIiKFl/NYCjQKL28Q+MOIgQ/3pDn6EL1QST4KozFz2l7lZzRJnt5fElObg
CF/TpqR+cs4NjbWa4mt8gF1Qp3Y0NQP650Cd/OCBGhrkbE3xhx/qYDAPe98cYKMK
V7kWL2Z/7k+t7+3IHhNC8KZrPmZ95kFEds6w4BOOwzAbEudFrqe4bayYzZPTYmX6
uo6SkTP0zsOMBkgjVMU+YOwFzYizkbzWKzk8HCuxfY1EKTU8kLP+cMn5sfgkZcgC
QlasROqbHlsk6OJ4m6ygeNxQkq3a7ErPRj31O9PdEoPofrl5mKDlABn7Sbf79yKq
np6LeoJosVumzxRgljqhHSRPrr0dDbLk4n0G7+cLthM5zq+Uxt5bmdjSV2yPuY3Z
Z3bvbD0cE+4p8x/bdewW1onvvUKMPxb/hwuHddb3y0SyE4lk5VonhKETSph39JDb
G+58S7YK1sRP2709W0EvbFwHrZC86LZfJVDmTbh1Dbehqw1xMEEoM92T5/LP6d1K
j2rDfOp9hbuJRk9SmjvUnpONv00N/HPcbVzy6dtg36x6VtDaGlcLOinKdph2wSod
ktIbTl+TQtjlYYZWvhq2+U/230AoKEZpI5q8HCen6TlHqJo5uLZHggJqIFLggHp7
j2qigo8fT/3VmTKYzWmVQcPErS7remYe028LAP/3y3FFNlEuZ4wjea5yO1TEbmV4
c/p3RvXBotKjTU8hsn2DALlZDPY+ndTN989iI2MEqZywFX32cODxkYsx8A4eJ7Je
YaItb5n3dv8FUKp5iPzkmUGjr3r27ug/wSsEgSvpzW0Cji9tLHG1sbs2ZdGRtIYS
NIgw7y0VfjpqzlINzLH7673Rd7CrAEDiCdG1tt5PpIz4T8/IZ0Gd6S5rJ8nYgzOE
G3Di24vVj1FDug+rDaaW2GNzOK4JYUliOIHgDkHdk40geQvzLhE3h5Ku1pkjP93P
zD4hqWOYfPL3WXLRI2RlL0EXcuB20mmx7/8xCg/nVaJCFrE9czTmwkkyKrGvxtp2
NJTKClwPn2QogjU/NTe/I8P1wXAmPf+Eg4nBiHI8XQuDHgDMgtEfJRpj+DXKmMBh
Inqx2zhjA2NbSmWR7ya/dn5DWS/oIzCcCu2ewwGw3vKd4XnGIwCcQO+epDgWl9Qc
gk4w1Kq5hKJb+e3BiCk2/H06hXlplqoLdLzkezwux7ERo44Y1AyWv3b5brSAQC2k
W0/jRUViq9OXOD9KikH6vcNkTcI1Pkjxn2+g4siSsJzHWuVlrbj6uaZ+5vu7ln8d
oVfX+7I5fMssc09d5ZP1ICkj+0aNQwON8fBl6DB4gh/ETeg2KvGW+sCeZt9QyMLy
OPPlBcnAUh7nDJ9QdnLLHhkUp5aSt9dFMlsLbqwL6U4bZSneB+id2xEyeUvxxR3c
YoMXkx303uXraIhnC69cUgmlWxn6annmiaAZ6q7Jf53vr6INSuDljhe5yMbL84vA
Xlg5sZj7y7aY0q0NHlMero1DhIn4mHjiEKOTXkPvHXrwcduWNnwT+J7ptfdTb+Nn
mR8E4hHnZP4Tw2XtS6weC6zHd5LyQSmTeWcpsnpQNn/GlBsIallOxhjzPTjCaMKn
6KMZHkg6bABNOmJG0vzU2ZcXMFFpLXQpDFURDnnrQMNoij90Zo/XDqBtIAa6Yb43
YSjwuXi/OUwmwAwuXGLNMwLY4qgs1fxRviQZ7ZSlRiIpGauCaVcrk2gLvrb3icM+
uiltO1y6ox9b2yN3lj52PEdgYv+Dwp/DDXPuXeHLdZnKLeAVMqtBIDf514k0Ucsv
VZSga3F0qd86yj71cGAsSA3NEcqNDHdOcaLdhf+y712v0uOmntGrRqtQfwBT2I6p
ClYB+8XlctT4qPxY5B1dn4nIOnpbpMqQx6ip41BUL+7Zt5dx7se2pelz2Hmiv+Rj
7x64SdC5kguH5CybMcZ//srgb0cz69GEOcoST6RoRUC/d2sscOTYyWLwXIYyUb0p
UPe/9PqtSMfJ1RGKV8SfChm8AZpG1DmD0zRUMlxDVdjxpzSyVfcY4yabISFVXgIs
uSZt3Bmou5+CZb/xqEmj9Slua8/SvUUZzB4rKFEBhhtVfxy0WM8BT7QGpBXzJ/0X
PsvuUg6KeOp09ppaOCaFA0ae84lwgdqa/CZdxtc/GnuynqaGT+/An2uNXTyMp0st
8gAJSrQcb+ylFfs3+lW91UqWWEprPq8RABL08/gy5fLwjKUJ6CAWIlzgxHsEZg3l
tRmfDZuyybraxjSrdM8+eIgsyWQNUi5xBA0KF46oy99XpbvVgaZZbcV8z055XKZw
ijQpnTydDW+r2iH+zjx63KViJq7WIJH20pnYD2ChEW3Filu9Rgsd4Opv66KsL8C7
iJofPUFbMMkeNsaY8C5F/O+xaD15ulZECde+sA3acsqG8fjN6YcGSSH9AXN+Yq40
L8x1mulmAN8kU+DT27reDFukQspMxoP8LM+4iYv/C27NEGTY8hut1c2FVBZ3/idC
Ed8BW8ZgaKYqtX2xwDQ1w183bmRhVk6pbPTuhdURXWJYNiBLDPWfp1UUjJyb3efL
vJbScxYfB9VOESks/e9HnJxguy90HAFqGRqrlXrzE02iEu9vr3Cnu+mt3nmrqv2T
1XE/OqvjkJBXU24ZmSS1JhDKvmLmHN7ehoo4GpVF405Ym34jioxfhC/KbL5kZpsd
F9z3GhJZWONz9foPZz9dBm4ch+zVT0g4hF2zCsUr6VcPZzPRCsA9tJGEoPjMQblZ
oAPZZmMO7GUeUQqCib4nqWaxCnk+ZwRv2aAciVFI62s07bNhn2xVs+dG4dVbC6lM
qB1xPSN7TRjVlbdDvokH4FrAqq59pjNH9Pu3mEAA8d+qb/cprgaB8lZWfjitMW7a
NIz+AyHV7twWf0yNZJ0kQUWXQ7O4BZ0waRMnlEC6j/G36aJl6Vr57Dqf5yTT2+Zc
sQdnuJ1xsW2KTcXynlZXMe/40fwaO0oD1tHSwURF0mCv6kJCFXObXJojEfvy8YC3
3pkqm4sn4xxOBPeKbKBxCh1orEqSfQP11HEvkincxUckh+/1Yfg0uzS9KiM6mbqN
JVy0ht7sIXR5oxYTtAWL6vyDQW+x6FnPGHSaKdcWgIe93xLd/qNzPyoJ+yLtFYgI
GrboVRERBZgelYWiRQV9tHxQ5ohtUpJ6Umbd61Ziq62dZokwUm2+o191QWJ+lQX/
Dk5lpDCykVWvVFeY7nL0c62J284X5c1sWkh1ecuKC1Uy6C9DddC+2ry3Gl4uWe2Q
4IKhAvEy12769rrkzpU7+f77/LNzjly63QZ6KcW4Kzf4npmf6g/cxdV1XrIjY1Jq
7smTFnYmAWiIGLDUTp6hiO8SIyvAoUjea4Pdscn6XDhKUujXynIEVHheOSdhHSLu
aeEpjU2ZzSMD0d2WUFIHB4vngpq1M9Q+PjVi2dUSILuBlEGaYBTYgM/vTodN/4Dn
58+utrR2/PWjtadD9JVShDvRCv1f83Cvio8o28ULhqp1+GWzt1qLFPoaWK39Sucl
A2uj5yf8IIqTI9ajKz35xT+JhcBELZKrPm8wY/BTaIqBwU0EKuJ+GzEup4Ayiftx
Cb0vIayY1jNGEIrfEu5hihYFpW0GmndidkPLq6q6goN+04HUt5aizGi57H+TnA88
UI1gd8bhx/appCx3/376LIyFvTCugVXnOfXSY+RAP0A/7t/ZWi5IgNuaHtF/W6uS
PkrrM4XJ5m9eipXG5Ek1Vbs8nH2Pq+639PFI6qqiB83EUz7Y5jkbyv0RKBF4D3cK
OnRXrnDNBZ7ijh3mDWtCU/7DbKwfbJTnaOxTpKWyQnFGoj6Q9Al5+iPl4ADk4vch
WES5hcfBJ7cDPU1YS5FGpvQ2fg8ltNKtWLRQAuCNnCAFZm57WnhPGEISP3horhB8
NC+gb46uc7jm+qWiCNtQdPVshPaE6sbQxFI1xJ9FzcXSM0CPCuUOSEBYW3UzDC3u
L2/lF1VB4YYkit7OlZQ7uXFvB8ZBYBoLE4UBTGXE3sNIx9N3pXvYsLSHuNtk3c5k
wIBrXi55b4Cbj8ITPXJ4p0kNt8MvYx3aIroU0Zcg8iXJWF3pORHrtGJDzjWGHEiO
GI5xgJkUxDq2MtGj8VUGoKTKDAwmh1hn92HWrsxD4Q7XIbIVT/jLqb2GD2Hwc93T
5SNvdlzeRhsXye2NSWLNVGQ3BXQJTRaTxEUMNQgi7Egb2DCzX48kh02FAxPXifmc
JdIhylfA5+KwYZKPGwDiaNlYAlG3oMO6TK7ltO+U5PzjbUd4rgdMTxspedV5SN6k
grOg2MOgef9YMfeWJz174abs8vtAV6Aw3LNG+u3mEmFIEK4Gvji5vEToPkMFtz0Y
rg+jvQ0l1HRAcqY4S+lztlSDqvhc0C/G5IEQqL2NhkRjYhknPOKDVWlmkOjXXeHv
qaz7KKS+Dmt4PtSqaLL1w/BDY/N8d8255+VmZ1biZhpU/NFxqtL2lAWEuI/+l+Fr
337qYiWJM5olVrlX8Rnm8vC9Z2EmkqcrfEgFLD3EBCKHRW41Atnx1erCXBQSWCcG
e9lNzGxKLwTqhIpfn5xUy5dOeiUqpY/qXp7bTJmgBe3q1QOhzEm8AcHbfqINIgQb
xD3ti7XymNyn9a/AxIlJgXBw1VljO29dUPcZcV6s15s7lU21gPsgQlD7clmbDTNM
2dhEk8VKoaAtM57m+ANwgOcV7oOSgdA5WQgBOI8mzEwEBWwurz19ZkkEh+XFeXqT
bs42gqxZZkTVK6oWTUnDNNP6jePE7v9Wtbr0wotBpiOxIKi9ndGRkNzJOntaHoRK
Ju0KC7hSMO7lLntzncbyDxFTyKMoFd+4MotVTNCjBCLA6MNA1KGjvUsykdaw5G4e
YmvjCnJ1IYV+ffM5+G868bcIP/rgZwWeUEUm4o/18BFS3/u4J4meInY5/D0sAJkh
cdsiOa8Lw8xJoANJdYOBlgbUVhP/tuf7X1ecIqmsga8EBQMGXbeojDIVyy24n/5x
+yK6MW7Z5oe9czd6+ZrxWTYSWfQ0e+t/J6o0EdXmNlroZoTzY9u0MznQ4XbmQNjZ
EHjm/S9TkU3ti4Ua6N57xZ1Ah8+iVawAyh3hHHhcnKywg6vW+iFkyd+10l5Vwphj
dYXa08D/JuD1AiDL2i8+3271LZgPvjzZGdGdLvGUKZOFavEy7O74x3AKA9+k5g7m
PxmNMXNXDZBrc/ob4D6G6D61lyay+gq+f77erQyl6h5OxxAXbhF5KYxAKzmVch9r
cPIYPwrEH65rkoPTiqwQmH08RrudiCw1fPbw5HvR4+HTlbZANjrmBRHkFGeM8rq/
tPcRXapWK7WtgB3ZteBCzCqhKxeP0GxgujGVCeqJPUp30waK5LLuqlMgimMTMD3m
iGd6ocwlXbTi8q89bw/6FsTa593qLsVZ4lzFzn2EgeJW9AGaAl8gFdaI183rzMrJ
25m5qdPRQO/U0MqxIVp8EE35BtojvEWNq4mTSQJcZls8pzE8xpKRoks2ULONXqlX
JG8YmPBV0vtTYpVUBto/XAC9VDisOudSgAUvvJ9ofAAgKTJ7rdIGGTCPp4zrwvR2
aI9U5K/+PkRDW62Et6VdEmPpbi4yG5Jj2jtDsxAn0B+9p08/Bcj57KMSJjHdHElH
mejCHMoeHfF4L6WV6xSxeYoAHq75GPErRmoq+66EUailho9iHa98d51HS8xo2Fgb
su3EdtKUMUhoPNUhBxfeKm8rHfGCQLSL8nz+N84C4C8+Oo0WFcVy1AwydauPN4E9
jgAMHTzUiEOzwA3Hu1Yr7gqvrMBzN5aFwkP1yB5jYwQZ8m0S8S7DRkIx4ns0uJa7
isSeYQ4UCXDaiFymPV5K0p+aVdwmZscaegtkLLBSVkqabf5hHiuV1PU7Vl1V1P8y
pSxV4l9Xp9DX4zR//ljc7oRrfxyGw+YFSasc0AdDKF5MIYjEK1KdDuzfIgZTeQgr
1qZZLJSoRxHCX1/F+5DIcTwgA9oyw/4NbkkF6C1YCWRK80IST2xeT0lszk3XYHKb
ObUk6C/I5sUftW8zIHTH8UsR3RfqCPODM3m0g16ZFWSZYc69E1yYhe+Bi4X/I/y/
zDLp939u/0P6+6fCcjjoaBNeLAxkmXdFhY0rNxV2K2vTkNXWz16GEj0ZRBoiAvp2
lnoVTvfL/2YRWb7wtFGeZNBkpD+r92UfyinXYWbYRz6brhZXaqygBJPRePl/9lwD
XNMeQeAZmoucp8mRfL3XwNprwnrIAHJGYtVUiQZ07WVbBauyI0pAnAczACuxVeN5
nnH0ymOS9N7Vj9gdsH6X5RFyCgQ6BGn4dPii0trokbDJdRphH+9vdUkt+Honzpq5
vW9vs6Ry1gfNsK+XgjPCwGhNs+oMSSQWQeTy0EdXx++C8Toglc3o7cEAwJ9LXhCv
KEMhEmPzFFja18mxpbaCToGR4LFCGVzimdO2msX0CYA+70Ws5OxntjvG9/q/vviR
n5yHq1IGNgVwTqYkPEuq/o9zC8NTx71HkX0H1sEVLiMeZ8m87GBk6i8FvcGQGshR
Ts0kQ5/814mk2bnEEixL8J7DUqg3/boNR2PXEknsVw3qs480/QMUcisgFwQbU9eS
VIUWacqtfWug0dPU1awf46YubQRndst3nd+VN6tkqRzUC9/ElHJvlMOZLoz8YTiS
WtFpGmbzVHU6yMgLk0MeZwA9pVpa6L3A0YsZRqnmEUydviwQlEIivA2KlZcgrPnp
B1czLwhAvNZKfE13+h1teNWe+/H4DfnfivR2JJgUnkbYL2mLrbP70k4qUOOXGQoF
RJFbRlQW8Z/gQ1RrZ8nJt1Ro6mR+sJ4Vsmflej7Kw4BEm/1p6LDC/F36JiswvBs4
i/Mv7dUtG/2DRNYzX5HakDw2KxH0GR1Bz6zuV0rqSmFR3ysFEf5x5ISqsii0KP7W
wI3D1aFROquhcZZGApAear4WJWuIV8bMs/GTZQSEG7Oc66/5FIbz/Bz1V9r3O3l/
mzEnf16NSYBQx52i5RJjiZgdUdox3nyCoYDP4AKrYnme5peTkZHN4yyxteYm5k8X
CN021fwWLZYghKUw36bZvdypL9emRVoZWH3s3fUx4e/imGTGttQVTtogfFfUIJdd
ZKBJqxxYe1/nbSb+kpHUBgZWZ+fPKUvmmjtaUNvO5TjV9hrFr+vuNttWSeK3kGN+
5wAETP2q1BsBSzAoiBeUhAptxkND2t5TwqngNjiUhhepXIi0+mFW4iMIyHBlObZt
+PTPols4vBJyv4TrvwWqd22bk8C7Af2z+nGyvMN3L7TscCgQAYbH0weGkMaucOy2
0jRlYiDDm+sc/CMTUgDBxZ8jzaU1pQHZV0d9nD6ENCBtuxuuC9dYAefOCwPFNssd
UVHeyPUdEUcEKY9ooQfpZzisc0pKZ16B3/BwAoufWjGtkDLSHuDPTh56kYCDQtoY
SwtmBcmZf6hFZk8Wz7oIvijq/NVz8Gn+uJkj41eB2wiKGBFEYPlHspmTM6cPpuiM
8X2it5aMXkgM7qLfmS3WshCofHKKBu4iI/U+6i7XYPS5zk/Smd5AOzzLthwvwwrO
a5AdPmWHxoWzgVvblGwzR/W2tsVTlqbIPmsoPIIGGCurEAdJNfQj6gE74Q7l6IKI
YScdUlkWrYOG1lX4el2UbJcvJOSjjeXOKzgkwIVR2TWK5rLGtO/ERgOyMuzdwcbF
CYPM3C9Fdyb2T74Yoq0m7K8ipb0yN4dKQFqyO/l+CEEKvIXA+te12eYnYC9KZ2dX
rw3723j7mVKInTk8exWChtv9gDCA8Cg+3Y8b3f2jMYaMAUjDKVIHhQH1pEzZXvDV
vVv9zJ6tbGt4HoZfzg05c5/BF3iY2p5aDZWmC75cznJjA+LqCd+SvCY+h5dS6yYw
I+QK3qTBBL5861Z8jkTeFDBJ3RwAvvv7Y7T3Uvb/0Au1BCFzZ3pJSvusM0PSk4UJ
eQBuTJv5W9273jFnXz9anyddviUHFnkKI+xYkRZgQovqv1zwClLeCGJpUJvdJdpp
nAfbRwPYehB750gNZrZQoKyL4so3UJRWfEB9qT30T++Y/G4P2TIjy5ZzQyg+K9Mt
kgQCKeZ9LE/dz/bZOQVAIxmkG0AjJp0HhOqFobs36MMIWViXudkO/QJYbHSdW6Fy
pvJX1aeWNwLG3DMyRxf3XCqr13jqIqpxRyeSxv8T/nnJwvhjTvau+EsrA+EucrOJ
qnt9HAlv7fB3ZpfYoT+GBxQ5IUcGlfjWsrzB5spLJIn7/KNOwjNhXbfFunYyYD1V
+GATH9oqo3yJ2totz0UCO6xgHcseCz8EVhmx8z8Wmb2x9+kQibh/I9YQCIHbzUiG
U/2BDoBvC6+8yje06r3OjBJIfh/kRhiVTNYM6QcXPuWhwNeppE931J69IFWYVS/X
k8iiCOMNhRCX85dsBaGAm7NKjPUBF0+ZpBuJl5N3R+lTcZyAoZDfoIjXBtM0pGo3
oFWvwJnESUfOKEMaQPDUTbtEJo3SsrkKBl9CHFkp4gc7Qa8d9tWvVPQTx7MYtg4A
c4J3aB2dkpisVmX8BhKB/2ed4nmc4EJts5I+vxkMKTl4s6tmQE2vpCu7XUlfSBdT
6mGDbJ5alOExBy4MNwJ+yCnbBrbkyXk5NbNcGzZkdgvYkvDkmazuiWMvhh0RcKpg
fj+l+uOB0JJ2qmx7qTg3YkU42LovQCxcpq5dxSXK2AgjvpDLNbiPYxuMyG33r17J
KBD2L6Mk6uLAlUcaRsy8u1GPLfHns1KnpSSl41SDG8JpAUNXK5nWBJKf0F9SlAkB
X4NKvofX6GJeU/dicSLAeh6qFrb+Y8BCzVs0ub4YrCoq0lLDLOfA4xoT4XlezX5q
5EiyXb0krt5Tzm9cYW77S9fmfSAa7tiIWfVTtMIxjWTjpVEREFE3AXudjt9xaYOB
e4Kg5TZcHrOEy+hxC3O5+iAgqKD9Xc4waDL8N+eCC62Nj2MBVtakUYnbM/C8YIlp
MPHbVGlYvN6VVbeNIjq+KyjYCBJM2Pw7ikYTp/dF+FXnEPA092BR13Q6Q/nA/kiV
80XQWdRkeLHH2CSkglntrf0YebemAw1Z1hMVhRGAh5DB6UEdLUqnmBzm+rj9KvqD
QzC3xzqaw1TINd5jRqt+Vrj/i0t83CZROtoKn0smmv/2Ds7bFtvwyEAzR0BsFmVy
cnQB97v1kWah5DjU+4Ujxge3fEqVB50h6pd1vVYl+bMnHg4b1OgMnaVLunR/hYpL
o6RDi3vpA/sW8b29MfD/cw+odI0SSOik7XytsuxHQXAqs5fJNZHCLZiAqJ6/BLBb
WCFvOBrQkCtWqTCHRHTHck8rqtM5mUe+g9CBRjIYHKzbM6WPwLlucsT7g5WMmlpL
pgxqTtZYZgKVJHyAjRJNi537vWnYgzsHt7+5RTplJiGdi8e3i4NhGmz6XVEN4/of
nmSFLHyZBuLxPAyha/mFyW6BTObgH82gWv4nfhfl2VjsSpogzfIdSSRsAfDrV+0k
jc/xQhZs/ADYbM7zb9RuMDw1Ubm6BYwp7Zk8PnKYYTvAxlzY+pKyT2L6dr+zs+/R
0Hslf+ngJBxrc9P4/b8/VmpFnHQBn4dScQkvFN4jP7MnIsOBg0AL9SzAewJUayKT
sNcRXck+SgOUgx6NHomcpHaNW7Gt4Tc6E+2USwpzhiq09bGlgPDHbrhOpJI49aib
eoMHBxH500ok1dlHCMNCw6GeUZyOi8WMXhqmuabA3rqsTcD1MvmqL0M9Qp5X4QLn
AYcqJnUMhDbNFA/jWI5T70gXdL6OLBel8j9eLOJ8zCid3Ds3dtKc4mJPimNAZ3kS
Xf3CzA2tPNBPG4eoTldnECpkXfsBnnL72husjl93kIBvqWdnC1TkN2B1V7G9F2lu
jZWE9M08u1xM8w43hVIv0KlgPKaSrQ6tSn/YmO/Z1HvizzlV56NDb1Dy0+0MWRkw
fyP8uPmo78bOBAVhesNH282ll9ylUZiFGwsNttvLf+GGsJM9XDACx3vZE1M+v2Ct
QS/KsMJ7hzPpiLfCbiG4Ubgeoe8yqfc10HPbYImQHowdLC09P8Q611u/j2aBOX4C
0fvxUsjj03Ouq+6w0JtD0fJj4QKyVU0v/16OjpUmTkyThB0dL1jgZBK3vns4piq7
D7AYpU0Y9DmSuVeLIu4XQj5jK+2ZKOQbtxoQzinEAY394jXeeYpqC/mOcm/mjiZ7
LMImOn+Li/SucBCMjB+4MkrfkBYAU/HXQFF8VUq4PFxhXrrGUTu2pBbgWpZIzk8s
CG56P5EDepCWM/YRBTZj0izC6q4CAP7x9F1bZZLH5qdpCmuP7j+W1Hd90vJY/t+U
KtGzw3505HlLYUWC4qYMRGMwHiI6KnvMMmmvU4qjKeuAw5GMHdCCoPWjbTrkSKgP
Do5WEaYAlisT+Ojqu60gU5KmSZ+e+iPbAvxYaG57zUidfXAn8w2/i1shKweMA9PB
CFsyBaUXKAJnf4RX4HtONN9iQCmlJMFvMHF6Z6YYTUVrKuVNrdOt4YqoaYqf/ujA
Nu2ZmpBPHkrNnKij/ixzj7kTfW2WLm+pcLCpBiX4RfnCIulX2XlOTPf1XzAGSCYK
h8fWW4m6Qn2fJKxTuDtwNh2itX25OIzf262GgrKPwp+ibnB/Ta1NcrPEJUaSogaj
mCpNxkY+AC5eS0sRees+vDrJGJReYr9wk58kextsuUU5mpAlM56B679ENJvDjAhS
GtokPrmcxMgMzF5hiOBAfBDNM1qqqAAHZNQ5unk6Dma5sgIIeAjDbNWNaJukygSk
5cqA0Cckt7xMRSIRapZMBE4AtliJcHxUNb8kZPObUggDGqUTHCtpOFqQ5ly4aDWV
3pK8DIvLZl3EC3lPYRE0LQR0NjJli9THa/PZKtCaTDAgor8hHgx7OBjgog/iB85p
MmpfRqtJBBQVN2Yx0yiTqDaSe60BtROplD0gT2mP/gVI+lHDaYgdFPreqTzP2mrU
vAxhG0S5hg8OG2mf9fi1MgucLBLlRDRNn2nb/UfdYPWLDtX8KJtOCDwDsgBejv98
l41IBWBKhMQJ2XuhmJBl03dKkInkXEND7DLbvMJSM8zYnVrh/Al+JqvVlhUihjYI
4Z8nutYXUZNyPzkpU/ZAnV+zq8x6z66EydSpN9cRDHoYh43GbrNFmoRPrNUh4t5D
z2v6R9pbvp+W7zio5If3LElEX4e+smlHqiKQ866nAFtbTY+2wG79fftUs/f8y9ZI
LjWlZiBbMxpa090eRp1VHT5t2ugAFLzO7TfNc3LSrRuCZCAcAoXIOmEVlckEsal7
CWHLcCQroz2J6zcuIqS2b9Z3YiTNye+nxiLHM+kGPsw5QWxN7Uk+/0mCPNOlyc0e
1Rc0rLi+To5vTdgRItbqzSb2Q8VqB9fFJ07E6lGMJTIDnS9lMos7UsFZ8qixv0D/
Vkc7F6v0rmCNiW0IG+jHButGeCfqa/0ygPZ7QF3xhC3Fb2crVcD8AHHnwFJIH/8V
r16k2x25eJ5ug+mpi+pdONnPza2kqduBQoD/R9xL6A0lntxCdOKxvxOpMAcraEIK
qZUf6blE1pefIXUYuYqiGz43MNEsItRW3WuMi1C1oqPx721FoEQTnzDlRfCZ5fAF
z7iV4AB8jmU2G8TLZAH5STEeWBInk3A5c/b9boWTBTNJKBisIERWJ6mNp8T8XPqe
n7malb4a4pJBX768JVlTamY0mZbYWjFzsJ94uztZb/U3ZhAny5VD0OFn2MoIyOjB
qLlUSI9M/bB+BTXgGuvZHDG/6Gm9Z1v5NkZBY8GSnD0Ytz5y4YtXnPJFhTkuOpqT
zMdIJdw9bo0EmhrvsuMt2o+8kODIjEQtmbepzyCm3UM0lgn9PpnOlN09PAGayX99
2ZivHaammhS+2YSi6W68CPcdtP2eHHBX/hOz5Ls1Ow+A0hwyaBQpDJGI3y9SnIXT
oygY3f4gr/H7tZv33RoVV+c7k8gp7F2bSJRXJkVUfZxtFFJN1QSt9O8tPsCm7CMU
RJGS6sfTga2Ruye9cwhkW3+vduKEZYS/4gk1q3H+GabkN2cZyqhdxKtO7PAzWCQH
l6TyYvCDE8Zp7FcPLFwl8e9tv6uf6pQX9ZdUUVC8ZiNHulWesXUnkUBnWeU9Tj5x
w5VSVzRNe2beo34INKVvbPWod1FR5pB5vK0LQLht9UcCXEO+9vyqtaPzVIs79tHg
Zi2WrDyKWWcv5ZI56ckqTOqyIVhbWwzD6j9BXqtN367jZIDJGRNsZcOoUGJKeLhn
xR81k9+1mI5SSHw3ScsIo2X2kTCyxfVeA3mTfM0xFheZjk/oavWsCBBC13SCZsty
COdD111QeLDomRueC2u7PNsc4NKLwHbmYGUKhDnny7lkYt1XoHvOm7ELAQ+FuG/+
CAx2HaUJrvDMTLTOpGy0zafTKDgi6C3MIfNy2zHLUpGnCjkIXRbi40hS6adFfNSd
v+ikwRqjIacpXjiRFQo5S+4Om0ZlZHYLkw2Zw/QSsIjdlIKkTCcTQbEoaVc/u77b
YmVxoeHfJB64GHvlN+wQO3rAIDN0GHmStHa/cQKnHx7tkL5dd/wEJ25jJNrdCIVF
JZQKK2uA7xxxa5jhxz6EM4rdVmJx2LGvtfvLjs1jr3dd46zhxElFyNscnHvRgkCq
txDh7uOinKxUPAuAB/6JPVO+1px5ITvsMJul9R2/mN4iiRQ11BauSHw4nYWyh0Ca
awgFIw+RkV4KsNXpzXSSvNtqyynIs71F891+ORI/keMAvxVWxzYrjwfsC8uL4tnn
AePVg3xKsntqo2/Wrd9fIrxC0eHK7RUBW3znD2/4zOfDNSl9aSK6dgNJ4lBxgR75
wxuSfFJZnQewMc8wGSvC6AFc8vAfnFz0YPlHgBXfMLUyk4zueYNrz72gCDjdUFHO
TBO6655a287zuQF8i3z6PrY5HEzm28zswoGhks6GiojLi6ZwbIFKDlNDwnAi3+t0
vXzBEvHwq8S5bGdnd6FKVoMZRCey8YewOFY4LljVsQs4ISf3qbVd4YAnuUrNirBI
UHQ2pLR4s9PNh+BNSEyT0kPavaCvWrDYmuNK1tPxxXu5Zv8n6iFIpnGEykD1qDVk
TOLAxT/rBcxEiaFeSDMnLl3kIzj4bXM4iQVh2icV0zBk0aPCUyho8bFEG+1f4xWz
bn5akQ6BQbvg7JIG1mpxRsgsaCzKraGmDcTg33HAAjAsRh/qN6n6u21dXhcavDo9
I/qNqot9246eXiX+35Byvn87z+LuvllimSDqomOL86bgVzidEaK1b+OAHpEoK0Uk
VpmKzv/QI3sC+fcZfctOcR3NsbKA0JybTNO6KVDloacwFhr7fL9kli80RAZ3qQFk
WzvK+T7KFnQLO9aqMvgeCPtqeo5ik3RREVihzuhvLXrztQD4A0XNcI2deqHZqVdL
ti0Hn3+lMpFWP6FLmsy0SxZ99f0KGY7PRSH6oInwkOT5ceEO++UUuYchcyy3msZs
dzkESVA0M7KMxFrDyOcg14Hbb7Hlw7I85WbUBEBIxVHWjQGPuQyxmhc0CKb77Roy
JS1nelXNPc2Sf/mnWIpFlC6nQJ6Pi1lE6JJtsz7hgKC+UM2wM2n5YJfwp4yvyZZJ
Pn8fovcfwEYjPlNzO86uqJK4EHQ91eDe5N4zHfGbpl/LqFdqS0DLvtc0XWqKjGgY
5YXSiHl5Xoas5JFulnLV0cZI0d/pZU+Gb+Ifyj0UxQk1sk2k8rHwLlAh5VQESLU1
8MJjVNKhLaIH1RpPbTwMAbkFGrI39hvOXF7HhakYxWjr3Rs+K4GYpvOeCuh1JOXm
lW8XBVN1bnqxsrSaUkcJ9b6OFD+tQcpIAXLYcl95KgZwTtjOtW2CjXi7FtCZ3K/K
XlqE28rvgYz4mWRpj2NTUM3l5kq+iz9GSxsHF7XOgCX63H6EVXyIrdZ3vNIioNWy
yAqfYnYQTTY2U7QvPvj3dkcZrLGqvXSJF0fA0QiniJTtYk3lSNtaRNfG8n5RZoQt
Dn9yWJvlJ+Sal+CIgfFdFnVW0nnyRBWBrZZXQCXb3q0pyeW7yI6lWxfeYWCDjfNh
CpWxbi/ED6pKSPpZgafiraZhgMHHtBxKT5E6loxKtdRh1DT9ux2e7IBg7ymWXFqt
ktVvIQKxHpFcvtug0dcsw/mMGd5bB/8cB9rvgmAf7fkPR2gQiSAfduaoL85tJsrB
fmXyXwZPVkxiWq5hb3tQE2sLi7YbFNexhGCxHKCycOc65OSVkg74Uq0nLQftgrKc
SpdPJUW5OC/sKtdu261C5vCEa945x7iUOsPLsFvbUC01GhpHlEjquria9EFxdam1
V6h01LLYd4dBho+ULljEyoKJ4e+PBCPnvArVXfb2AjoYPifyUpIOI0h86BQK2cbp
koh6vQsAaSFkZUbWl3c6MUX2cp0ro0TTv6jCGTOcvSzYP+4rdhGyeKxYj2W8Z/j+
R6g7MaBDjDxEZlyySfNpJyh8yWD+wlZMhbh9cheu4C3m+HT2zz4PjDhED1vOExDl
5gIMJvHneQYNZHNPpJODJLXDSSYTFMF2M1dNDIkolx6s9ApUGC9jg4DEqDAg1Zfc
zmJ4KhMIue58GUgrmW3WQh27PO2BFlQcmYrXXcbx3UePEOC4zTN8abK5Yew5+M+v
2iytZJj67S+lRuzdN1UnTmPssRg8SOkjITLgu7imeI8gOYVua/eE2s/6sh7fNcuu
kbrBh5BFCdekGf8MUYio6Q5UlDiJ2OUJLbQ7WCFonz+VrlIEONWi/Gv7tlwAzQ0i
U0fsRJ+QcgzftHXGPH25OVpRTYeadzsgrb2/PFiduBnoUtXhdoqk2NwblHWzF8Jj
B2ELZPtMpZmDGaZX3wiCoL1EQw9YX0fj7UEUzK2CbaRYqOAgzg1AbjFpLo6zrAI5
45rwPk+k4f4UuLE4inTTnbze/9Xyja273rALUdNYObxeH+Umgs1K3WdZ+LvYKXFk
8bWebWmiYiXVR7cjnXki6b4r1m8rb2V2ZQKuLzXY/wwdtykhlM5lo0xPy+ybxbqo
rVdS9y6TGo0DCN7sxXwlXrOZexRpxfu+BK3dTUmIwesQzaea37kXcsVEP/HuzZSh
SHG5Y61ZjUzzyjTf/DJYWbGG67txa0uZ/+mysnIbc1dTNXgMNOQ5cgXQPUe5AoD0
GPdqdiooWiQSA4tDBJiWO64DuNxJBGp4GIupdWPWPJMB1BKkONKjA32QxBAGuShz
VbczQeevk2tmX8RvU5YwOPtKNung1KsQzgKQlnrtdZqAaUwLyxOKcsYC+oWIoeDF
cHKpxYdbN59AI8qpg0aVH/ZeO39nH5bprBhvjcQmv2FOk4VDmLmDmTeeVdk3ZOoC
C16Fl51OUdJRDyE8H10f7rwMmkc1BzCwEXg3PzW7rSiNvFhVHLHzq80iv8yC6e6l
9f4QyBGp62lw5BVxR64NK/b4F/rPSkOQ9C6YiuAOXP6r6UeVmlWrlhyM/BuEvWpp
Rd1BkEtM7bJH8z7zDz0LoLWdmVQZbaPEAjdCRxztBx1MYkd2XFVhO1Ub0qyptiGA
dJAlOHFp+qdRbsMd6F6W5i724P/JaVUyzvko2mUYfUZpzhorZKbrx6tVcGSHyyx3
7vAVuZcHij2NEiG8gBta9ey8GcQFiyjvZ/JZqHWHAHOCxTfm3HH/qL6nB4BOREAk
S/qS8pA7kZRk1XvW4In155HRK2dJI6erWJlbTXxr39QYA5OnO3nZkxZlwdaHHnia
xQp/MUyQsl7H61Pq5IXauLxiKxNNGMCVf5n440JugfytUY2UEQLYlmo2km21IkBn
TgBew2LkCtl00biBWyWi9NIm4wAlOPXuxUQ/G3ZO9HlyhtU6E/k70xhRpsk46gd+
6r4rLDvv537AFFGilQ6cYLL0QibY1bSZYA5BVpfFuo6KXhMg6y1eHmyYQdBg6Tev
8IQt1VELe+KuG489brv02jMvhAqdnCCGWKw0vgFWNAUbD706jwoup48X4eXDtKhL
dZ6tV1g6wGEiALEoPMzOStLvbxDR+FUgC8t4/4yb+zGTSZXBbAJfvrgZXMfWslqK
S9SFjZw4+TLrLs1UPCzhxIfDOhPM3HCR5/QihRRgCTOtDgCTdigy6SLNd9WwUx9G
l64NQVjFFA4px9DCvyRj0QFsJpFbLvctBymhw27ojsATJjlmPVawxNXtbo+z2PXe
VFnuP3IXuMNHUlz5OlA6A26SDPdvPwzpgEX5/+LPkdV29NDh1/B7SCNZivDaMQHg
YcD4risZLz9eNnyfb8PgfIv8MxzmmWL6aMOH1uJOhYrE17JA1wd2WBWpSpEtyHWd
Y55RQLlIk0DCaBvN33GHp2cbzAyfAiFaYCK50K4y60/Ia4iGDQlL5A6fLe8uLnMl
jx6x5ZQgL8DeOB2uX5IdP5+RQYfbtXOSrs885hM6TWKSt5nq/q39/EOkm3kIJtUb
RbJQsBClrzXpTLP4C/umZGhSiwbxr2srxY0UXK7hJvvRhcufLFh8LhiHxdG4KXlg
0zUUnP9ofYIArMdEw6jE0f5jYxFqhPBRnNtqflu3F5YIFPz+maunznDzZJV7RmzJ
Vq3BXJyNMRJzGi3r/lvGtCS+wfX4kxCHZT2bPtcfvMmVGYxJ/SfqV/dz4NRB5mCN
TweTjDQaRK/2QGyI0SdaWIorZdJpcqKGY3xqwE1n0A8dXgHW/xXHnmLLgvt8Mzov
9R23U7otECGLGrk6yuZ4/rSAgQWBnBb4WsWGVmb40hzz5rcmLYEjHkI1BuLrK6NP
dWV+3Xk8myhfNzhKMlEquJi9HkkwvvviKQXvIl8x778CKkOgJVFKzbe0YG3v8tOe
8onpcE6nCfaNIYKYgccdzeyjeesDPihd7NDxxqcahilDnWufnr6KBDcpTxLNrrP1
38iFmQznRC3fL9c69rZIpr8MZvbpLbmDBgY/fo+BobEAMhnQSEURblYP1aELMivb
k5uXZhZ/N6h7YIPGtKvuFmhO/blluZxKlGVh2cwPHL2rpBY+SWIE7DTcetYbcgh0
Qggub7Jsg9IDl6n+Ikc2Uth/cXgi+5OnrDpWdFIsxsd5KOgW5d37ysHFQNXX6D0N
tY1ijkNbwyjebR4sdj032Lz1dWm9BB25IzP2xf05YLD1+uyBLEn1Ji1QLmo+JE7P
h5sYi4s9yYxHq6rAZympN3r4M3fO1/4dq+tRyIBPBl37tc7TCp4oquy2pBXFBfto
w2DlKDmpczK+FavsZiFtJPx6W010M2e5Og3fq5ED4nJ45zkEeYkx2O12YgkhvyA6
Tnz0IXCIptT+RmQqTAQiBE9NIU4DSVz0rmXo6cFPG13BfeBCa+l5oWRwaktwMiBj
cWiMNW5L1L7TCo7HzBzM/5XsR6RjnSNEYMbfcXxVJoQcOmMR2jYLZ67LE57lXczC
vUjlISI4GfFe8lGc68F85S5X3mPAwmGhSh9leLDXzmZXtlRIjrdFziBtFRxj0F7R
IibMpKyk9XCfEfJe+n1YOxf4ZylXaWfNLsa8WI8hlGZmMB9/+GXJu6IOuN5KNpga
qU5AlB2A6yza5cuv5BP0nK4IjVaQ1/XWbwFKHz+EBZSgqg6DOgwdoyI6yH0lnJj4
MTIibx0OdQk6d3Ht7m9LOGTFmKevSMN0oajG2QwiUQ33NNekZ5u5OB3LtgCWg0Xa
IZjBtDpYumDaND1jZqOHgeP05WwzDW/vC6MA5QQmyAaqFvKiMq1JFdzy0TJyQxcQ
GTgp/IugP4ju2lYUdmJbo90+zh0Jm/esge/WdXj/G+oXaSFLXiTjNrEe/Wau/+qM
lxPuc8d6xeeTGtRszML58fHntB9L96sTEUzKkBf4HP5GmgY1TmlmdZgT0fHqSlI8
64QNYNO81MhNtb1yYU7NDonF6c7hNckQ2cwgtHhqafHtO1eZo67KmTaPaZ2sJS6k
Kchk36Igw2T8vTIHCIr17XKtOdgYasZNB99plO0h+4EP8YJpWBUZg4VEaTY++d2O
faBZzFdWG6OE7Neh8mAgZLWeoc+x0V9pIYOIpBSJ6P7IN2ZGWk/1qWKmvqx6mKTS
+D8EOjYrB0W8Z4G1VGKdWEED07LVRrbTnbgbgcxIeZ171IngG9rj3eUX/Xa2FGLn
skAKAFRK2PZFHRlPIjImKOLoiV67vtYYeACmGiIQJMNNZedFZ2h6eRsv8xauJPc1
xhShhJNkgzZkRuAhu2tI2aGCo6k3ncMnLPwqvp+cE0wWoouxv0ARpwLtahv2+5LE
sOOz4WwKw3flUN1/DRGjYUjIH8lO6k1QBqAa5TDwIpEcZx1Qv6CvThE6E+mntbAI
RoiysNbAmvALyG251RM3yFgFBhEgqU6NTyWHLajg+rVIw4xPTh4QtZeZc9N+F3Rl
218SUQNs+UE7GD7PNa9Ro7bdZQMp7Z+DWYjEqXimPuQrMr7SqQ6Usw1AVWSuin2g
L/m+ad2pShQ0S9q9uNuE45S3D4ys2NeS2CC3GL6hS/uiw482P3uZ7VFSrcZarfl8
uy7rFHdCQnywZ0ViFLReSOzaB220ydbBzDSIULXCb6bICjY2YijoqDh43KQ50MmN
5majFY/kw3ENLQD/zZT0md359DlXQW9YBha7XcVsVpXLat8EWt1KI94ZxVNrVq9q
PLIB7pBxd37MfT5/rqfQqiXthmvPvJHkr04LQlRTyKDdA0bN/b/lLXZ7Sd9rlHGB
M898fzU+mbIb8/wLTqeuxrXjK81dseE4Kd3XIKbzDmZHKFzdq1pX2118zQuiOPWU
lT9D4O9cRwUFt1jV+2G28qtHQdh5m/d4aLNBcZDuyVw9eADVhCsaBqaQWW9b9ePr
p0c0/P+G4Q231bgsEUqzOBp6s1Ft7s5MwIbxm1I8XEF4rT8ZVdbDTtHjI04HWX9G
AT7p7capcFw8ULOI3+8URUfAOBDTHPWm91M2WgIrUX/A4g5px8AIDm8V11RnWssg
p/1mA5+3VLuRZn6er34vhHBE7IUXQnnIpMdhuXDpOuapUJtgffOgA9ozWaYIB8l7
kCAnk9yl6hHLhrkmgJVvdGccaS/augChHNLArFv0z7RHMBVLRNrWhWqSyHRt6v8C
NkJbCDAPMHRytKnSmjHpzM/0jmLqmWvyXY81Z+nHxxSjPfSV8LuHXQUgnSF6iHpH
4046vS1fJmK088yDfdpaGUcyrPUKKwm85dX8TSJnbKdYAKrg8Y9D8BXaHGvV8RVP
nXpGdYGzPylETUJpXFRfGW1Ua7VaAfw00r2pq87xtkKNpDaCa2cs2WppXkjZKI6A
C3iBJXnUAaCyUOpxvpy7R9wLCPae0LoJwLTLWE07On7x8cKbQSiTC+maSF/Ga/lr
EMQtJq0k4FZqu2mDqod5lhHB/u71CzgPyEEPX3wawyX9R/M7bmgcHBH6doECa9WM
x7eTNOj+n7HS7ihS3doJ4mQulyk8WXO6fv4ZPrPzqe9d9uHHlwADnkAmt+MYxtMG
kl2k1yFCsyUObw3lVo8RlzunzKRuSBqIwIeGIV6O/Nnz2D7v5357iVX30iUg3tY5
k/+BusWG2wdzf9DevvJnX0PQwwQj7PVsgb7LMzIUJeXKVsNmDrZauKK0AfvpyL0L
D3ONGGSfBWfv+5F/5AeDWQHN3Fwc0pYojLUHNnD6G0HQemjep5UTMWOQRPdp8ihS
9PH7/sR3rGe4FZ1vOKJSM7JB4wdrhkdfXgtuEPIAzkFMLg7np+L5YlkG0ImerxIf
5Lo/xPNUpNBgNmLT+zH9SPGcmoRJTQBGcjWCP8UEmAiV/oVvtooGeHzvtM5bKeuO
DYsdTKdwQkCJquq+WxgoA+/mTtQ8DOr8oJSy8d/d1D5cU5GrUmnRE87Il5tvNYxb
C/N3rhRrjB9PgUu5uJv8z7MZE2dwfysjrcWLB7vxG3VWOmZbIkbuYg32nJMuDp7M
q6LU6WeVTjw7xSJr7l6aZBchQW87/Yf4mpLfyCtSkmvJ1wE2JS8l0BTwSP94KiP5
j+O6YeWuTdVI1MkKNAgxcaCNaUIWfTawEnlM5FQQqYPqkv3L7SpN6bDsoDfqnvBj
5vKXjfT9e8J3kV/Gz5gx5Gr++FZF6rljA6VnfFbIUBV/XncvwjziEsFCgZ3S29Hk
dRBwe7CaZfgyyeQM/MSDpw9E0oNBLDKgo8dB5rz8pKWcOL++jY78QPlv8RpG8ENy
HAmEQRgzTEEYdPoq+USODArnh2Apr01H0wCQeO3LmA3SIfoinN+tAokPSPexZfa8
CKeGsg4kWJ68r9/Df0BGab8lRfx40N5UQfOJ9qRG8y240I6MH5NvWXLr3g+/7EiA
QZgKkYmq9T1LevCQxfx+56vQySUQzI1EMvjiF+q9wc48zjVYux61bmgUxqjxJrdn
5zT5BezLBG3boboleA13HSivHWVdntC607HkZLRzMEcAWFrGFLxCTGVzYnK+WPWf
Bj7xcL1zGeqR7CoUKgajgfxr/H+hZw/qZsxRoJNxBIvvnXFgHofRH49FZuqDvvg4
VrALCQkZlXfvuBq6UlnsbqFdMKi/OAzjnBPiLwMQh5Y+aoWP2u2N/8W28/WdIKwX
ry3uc0HdJCBLdpMF50CwhIJ1g0ISQWGQd6z+XWOKj8EhtcYBVNriS1TdpSYUbsXq
NY8cLJcQtV5GCeifRMH9Dlxirw/NdKbaYRi2Ph/5DzOPkAAPAzsOeofQyF36Q6SY
EG94pV5gCgEmZhhABmIFoTjCxCgy8bkk0OhZDX4xqXlKPwu6pJeWmbhW6N2JQfoZ
BP3pAjumK3Bmbm/OSO4nPliveHDQcIE7IH8hKxe3mZw11VdL4AGpPLTjNq8dwD4N
a3Xla9u6QcfPk+j+aiz+pgAdiVA2BbwG2VM0rlXB4PuvD8rMGY1O61RK2P8lBRtI
YgoFp9LyyTRp0ATFcCJX7A1/PaLVPCgPbvM4DRe6C3WeX2tFqfVpY/OWmshcYfUf
NDtR0Lt8SQMpHuo/03PPj0JGM3BlIVwmTJib923laIxd6hp+jDj4ZW0rFbnXVOcs
V6+jV8r+3RMj082SEnvTg1FnrqFpE0DnFpJp16b0FONwSCMs4wMKvEOptX/S14nL
8PfaGIlH6uLChSjkPGwNR+hgUtL2JTAaUlX0WLxbUQBFfZaGrtQQm61M4A0obKaK
MfaV39gRlD6p+P4e7tkiV+jbjEyQG/YZWyxppMaOeTA8dmMxVnMOYPlFazLkqC2A
CUR57iQwJKU20UaHtqPFPjN3D0PUAswFCfI8+tB9NfXMoIpebpzzvaqtldRm81+W
cOeoBb9QZEe8TPdX8NKq6BURsHXaX0QNh9ifGDM3ajTzHGM/eouspeZz0QlARdCs
+MUc7e5CfiTOe2Pq+H/fNenUl0jJioh4HcmX5tQy0kpB58peT5pKbd6inVQmtVMr
NFlz2AjUQWlTYNs9r2jFfwreu0fDa1QjGijAe4btaHVog3G6rXj/h1ZzVNp2hecn
i59yRUpdIRWwQ5J/QJOYMiCzoxl+cCdCeqSfDE7yeo+4zvXSQ9WJzADpHgXpohj/
Juqw5Xmr2Au5+XJzxWreMHK/oupcHCkugusRytQNFXvC7NvcCULWeUdEKLl2djGG
zWVJs42fqdtuPh8voG4Lz8Y8MEYXHDET8Yo2BH5pq2ph3KbvjeJGxdPSDLP4LTLv
Ak3t74xIuvAlh8ubD/9G7JIOJwq76yJS2+Lw9kvZ/OuTuL/ytrF5AA1O6SuicBjy
sBdpI7x4tw2Ge+yreSisG0jAet1vy8BtwSgQWWv4ke+VqGrHE+heE/kon3S4iekl
QrTK3EdShbq++dp2V4EeP6IRVXPl/eR3J9jsYcwn3o79IqvyAPuK9KBtC8kcKd/e
BMp89TlTsqLLIC3dzCXSIWXhZsvk1KNF2pMMPs3y9yBmsYTitZB9W3xAW5GlWsrh
lZnVE8DsjRz+QR1SybYPpSH5sOW1OOChuVCnG+rh317oLPA4G1O2UD1Ma1uvBQ2K
mxXRf1kVRr1bblmEUzEUm/suER5Ftm5iHvyshD87xIRtUPq4AUw/3eMXN19Hkwj+
HAMu3OlreitLQcEmcaVjeq1up66cPbk81jtAs1a7K0/dQXIxhhj7usiaVdU4LdXL
+kSC+wgemb4Rq0lj+gNzWkY+YnymoBghz3+GrNftIEqyJm2thM/qF8oXpWAqWqu4
Z3uepnH6fsZItc4hZiBxyQmMe0mjntRryH+Yoa0UCv4TrekM2veIQRvOoo+U+54w
t6Hxy0rwrrdPWPI/QiDT6+czl7xTETDgyvZ0n431LUcMhVqIWG4GlVo7yABPFoka
Y66kHZMpVYAAHKT47Hof10BjzbfDmzIX3e6a7Rwl3pCQq3FPqqfrowCSXv/1yXcH
iC41EnGJVs8VdueUjnDWLMx9s5zZuHBX4yFYJFoGUiXj3pRxGDHraqmEQT0P1MIu
+qy4/v8qIrQoSp5tqAkZ1sVkjcUE8PvzpnnXDiv/Y9NvIO9oWFW7B/KiHQ2DMh68
8fL9R4ErBUgXeXSeEW2sDJRcUbxEqV9jCziRMB3KKUyWa5bXQjNvy6WnFqQ5zeyf
8WuQa/uEF7/mIIsJSVsQAdZZj6JU+N4j40buMYM2mV+zZkknSuMbBpvrQyMLJeWd
mYzfAfmlPuYX60IpLR7MFr17v9yVqCyXQB2sPvp8qm1f5H74Ucd1jknnAwoVxHXF
lgn4CT0m0dNt3sq5nIGlmQhwR/ofXGRUg8aY7pCrNCy15x2yphf/SX4Sxa2pwL7l
hQ3mRgHZCxhNH7pqz2YdaxJDPz8UjSF5Smy1IW5p5CA+xpPl6c28k41E5n0n+6Ih
PIe67zHx/i1mOEoMgr/cO3ZcpdN2Dipp1filS+BbmQ84yOz9+P7oN4ZBD5sHnmpB
qe5KpXCAnXPDq1Nl6aCLwhQdtJ9EUippUy+E8gwR3PcCYurY8HwWBsSww7GBtnWT
Mc1sdMZXqMBwsQg2Wn5xD9hNHZ7q1c9UHgo3Wz29DpGXo1mUfrojn9IHVvFlK0eG
zmXd+jTDgovibA2sjbbLgAY2rYmuG+E3hphquFE+3/m4daoPi2PB1eMYhKQWZsHN
om2li9rS1VsltgurOZWYeT/xB0kFwDo7GrcGwcvVugb5EYhlQilpO9kieuVRjlll
1J1D644xkeFfy+THiHnnPWG7oXXGah0Ge5m4jqKpGAt5K///1cenNZq681ggYnyU
3hmAPSMxwUKTfFMLLdBQoyil9ol0RPJ+UVMIhS4gZ0uXLeXjD4BqnDBAda1jMdxJ
Z3R5wJJj9WG/pEXNWhfNoc1tXRUka6ZOTeKr7wklCEpoV617Ze9lW+VrUG7yyRLv
RTMqg4SDSMPNdG3FbLrSEQCw/6gAFVa5JpVMX71rzKW9jsWd9ArPm/ndRnrfGSgU
GGBrLkIz78J3Kw262rqYcTArIAVLSaK8rQEOv54y65bGy+apBrf/MmHe8Lnf8A1x
I5ahqdEFZ3izXFVzvt3lGGtuPOm4Z/yB4OkMb7SQGvvyUDNUcphQiR/n3eAiIs9U
bjSBtXOfw6tQQi5iZoM4H/LwoygsiHGuJL+5vijBLhNuYNQ1yAXfvChg13xD7iEx
PsL2DiBSyd4kVj4rCdOcZdkDMBH/iX0WzPxmJbWzxoBKnTKn5l6q8C/slFFQiS2Z
Y0tkJCgNpH/HRR9/YSy/fE8hPnvhp5lsHsxcFwMly/Bx9+px2cri20rTDhHkyUbq
FDZ6fHbHvNl2/KF5KUU4zC5Fi8fijk8yo27vjHvFUbrzOVjK9TocYUXmt1gbZvMY
y33SBXha77Fg44tQIEsRHYKYE+yxSPndwtYkjb5jKKGKjAflJ5CG3vthKUgJNfGv
GHzKJ6CejriG+hoNrgMQ/RO2MFWmpSw4YoBysWFTtzInP2EwrdLmM2YMY4O9hJCN
yIVrZzgVI/+gX4G+FQOjc7ofRswRsuGHyhB8MnOiGQ27oTVqPHSyVMB30gZqoeAR
1eQakfaqJ0tOdTMRHvK/4orI/lkGXoWq7CjFni9s+vqdEBZbQY/pHCpS/4kw5Zcp
hbBL1ZbNkoUdkQnxIjiPT6BzaFF8wmYfSj4qW+vOIkcVvYFNo2XwiC1y7JllS94L
x9CG1OMWbQyHBVZiwLSZHPgfg3yJKYQcoGsvH5ek4fuhC4kKzGgsWWgs8JbdOoTC
5R9DpoIjK8iA3X/gjnnse4jnG56SMA0Fp14mitjNoPXhlyQ6usBjLEcthSEbV535
jVXXuE9YcL1yl1mHFgckZrMjwkr5aGbDuarlIfkaXll3UjJVuxYDVv55KgmPRSPs
Wra5jZv6TvNmS3GFfF4aeD08dDyeETKE41Y4VpLF1a3ddC/khSDn70wZYmF/w3EH
e6dSTRvACM4gNOxfQQ9WLUoz3SDO3KRXkQVqLGgh9mlvJhGJeh8VM07UMTkxR2n0
g0FgPM7AQttC5fozf54FkwTrJeDbKwV9dzsnr7k6Hizs71xbIwsbq5KmnkkQC+DA
2Tfp5rHnHqFxO1lW7qq6YTueLO9nKwP16MPutZBlYiVHbhj6bqeJcsRbj6Hbpnzl
vgj4YTa6+Jhw9o2tOBl0o4XaMUElndsh09E8xLMUncZwGvF2gMJe/p+Wvk9iaufh
qCAaQi358sTwqk4dtQBd2LIKJpGf4I5AacA9hQRYgdeP3F003NSlkFpnO2PoEsn/
x9nbkwjwEW+tWhPnDjC0CIzxG54mb4/Nb0bNNlaXauzOxiKfsHCcc8pznjwN5yOF
On8GojuFTn8N2D/trTy8+YmD91EEK68jY1nhZHIByTDU3IzHg1pwWmqde0PXo9EP
iXaLIAGVXISDxY7ecGx4yG2aS7ZvXMfG0Z2Ms1MUvW8KRXNyBAlbfSS+nwRZB65g
bDCuYegiNUhuW+UK1Tp790hB0etVNqHnhiTg/AXfe2iqO/6O8n5llv068/l8mq7P
uh51+e3Fvda1dKI5QJwxRSohQeMX0Uf82zxe+NPDCq1ZZwnI4FRsZ1BnJzmFIYpb
eqU6WAFPt4iKXZAE8Lwls3f2ew4c7D7Dku3AyM+SupAmkLqxp9zPW9G448R8AROA
PK3YoKG+eryGby/u+k/DOxR/bhFKQCA+zGkTSqyIk6Wp7OD+QLYAPd5DEKoPywya
8hTpD7CE0Eneb8qHO+Ri2ThnlBoKOsOysd9MI8KZ0emq7jFT6uUN3cEOK+MMgd5u
hKqvUSpDnNFd2z6PaUWdq+I6iH3/knm4byYhuv4mvzg3fcQU9gxOg9lyhdA37Utp
RAz6n0PPIuliedRlTUQwLDjBTeeuY2xkJ8VZsT+Rn+Cv11kXBnflKDkF+5fjQDH4
BOPeqHgqX1z7k/W7YelEfX0lEVT2wuYhxuvjCpH+/0KavokoZios5YkErVfN+OkN
M20wXrjGTx4+V49oVNHQK/T5w91PrifiOAEqYfBpx4l7ctn4x2sbu0ef+WMih+G2
tqXmpzZx5h1QgtAs3vD9NzTP1QYi3izlk+GwGCv1Mv75DGcYrpx6har6f0XFK5Mr
B0yZL4nQrU4TQu3pcrGgE6YlrCTY9lmIEzHzBrHldKkOYHEX6OhG5JRZeiH9aLpI
pZtUvEiN3XfEECHngMBl/+tFprlD1iQbLbE5Zn+0zw6iS1I3KLYU4esYRiY//eRT
uq2GsmOJ+naCLqqSMi6R4XH/oHVMMEAPbRO2y0qs5JXyeEBaLURu6CSgbuj0HSS6
kYwUgwHJ0kWvVuOaA+lIDCSQHRQJpxi4kA+DZN2YHIXipvBdeXo6fH8Mvv14YiiZ
O83TPLyzMwLG4a0B7woj43BjOp3Xr7g4ikmhN5H7BT4vFcDFpiQlPB9Myr4PiK/2
PjWIiV028nVjQJFB1eXuEe8M+hUxDXeNQnFzNtPnz0Pp8RqtiNkfaMaoSRgKh7U2
1kF+EBLdv0bk09Mhm8APLXvCknN9trdtBmX1W72Iv6cAEyrVIpRi7rBzZ4bCEi4w
LktzQHRPamjy9sVKAGw2OiHrO5GsoUcuv3fpkk8kTDDR1th51gZJMDxqx1vWZ9Qt
uHDKg4EE1fA1KgCYYyUsNsuzqdv71FunJNfczs9X0eeBkOdqS8HmpEVNuJRqBrbJ
rKq6rD472laOo7jpjGwf/j4KLBCfivFnuFO+738xSeiEFYWwjhKCZlLvSfFfMLOy
tF0lcA6MllIbwLy6uFoVQ4iKPMMN7o5/wZMsFg68WYo9Z3lto1wPc6Q51nmifB3b
dB5vtbKDRpxy6fymSFtr8KI+O4zHyZrOZzbeSkXknxoZPGQjKxNDclb4RWAicn1M
zU37wz9XG8nlunMwhFqrqydp1ctxNhJRnvZJNbxD1SbRKtRGJqvi55Een/kqWd8y
s+3g23Z5IogbOvoRsAN+kXWfguSDh3IOtjCVMyLHHPZzHsqOSSbWuT9/VK38X+YH
MfUZDk53MX7y/oUwDhVq+qQGSN+cApaje9E0yqQHiTHhTTRC5XKqbOTOFD1b0ywQ
KkO2/V8kJ8FhthmOK3erPPbRWRl4dZRSQAgQAAtaOlb/rCBq9zq3B//tUNEIHZF7
hIE1+5gVGLhxeuYHZuSi1BjbN6VAJG2CFLoTTwp1y0HPpCaenCNciIvOCiD6w/qJ
qsDRCm14wK7cc/DCnWSHNg9c16d8dRLmtwwsKpaCe/xoFJ/ZJv92Gnff5/LR0L2/
soH3MOeHlOhysByuwREYjt9xJNBZZJLmk717qvMvQqGRkeNwgCppMdkxy8bof+PD
2aQjgnEMK+QwK2/BQKyx0H87+34vvCbQZv6eKJ8cJi7DT79AKVfdPQ8AdxzlZH9K
q3omaZJOEcP+iQOKDtYphG7cHrL3p+gcMErYWq8MDt/U3RxzSEAv12TBLPAZ/70f
5Bt/k4/bovf/OYwaZ/b+MDdAknitixd/RzT1zeNVWbUOp7e75QkA7/jQhHCilFUF
RDwt0LS00wqYLv1B5zWHnmVVjovd72IiR+DC5YMSxpZbop2hGmKl7ovoKK3DCnSs
YLEL7T0bVDzdVyg4CowXIpnxKw6iN/wUo5oOv5k+5iApdT7vyTc+jzAJ+CW0yOWO
vfLv1MX51oAPkViggXk8sJCFwdzqfnVWc76XawU6rPfnm2QEfuXQ7ffKj0RNLm7w
/QnIxMAHBSAvNRApPRkMugDcA3gPLf6nWK6t9gPZnf8MGMZNXStvjX4gwevSytr2
mDF86X7xlh3hRqSh77VIlnai2NHajyu55rU5U1HggOjjCGeW9KP79ACZYG2sN72c
7fibmRXxz4bUir+RmA+kR/eP1SxYCp8Aw/OuoB1YsPoalLBJhd7RhlduRzkctDS0
+xVSFMvT1Y0ifwPyYvN0ehP7Db4UsXRgMk89Jr5gBUv5CtQ4c6dYPmhnsP34jcod
Qn5xiR3qo/SXfpgIYWsyxbNv5HR7qhbpoxArC5qe+qQK+nkNDQ1N76kg9zNXJDOv
yO7+BsbAYhttMAWLr6q5v0o9Vg0omb6bwxggA20C24yq5oXBLkYXkgMu8miAkUs0
L2mEltUn/ZshihsV2nYX4U+/qwiUMR7TNjw00k0Do6CUyBYKLOvrqEYhQ2IPaA07
ysHPuPR8qODhRKuiSEqXbRliSUpi8LrqVRWWt1+XXG3v6y78V+dFCijZgd47cm85
nKmSXXu1L+SevXSG7kUG835WGFQZoHzSMLRXIAmeaR3aIeRUyOdvhv2BPJMB2J0h
OR5+m5bWTLSnAWbXTbE21UmAAS8zEJfDuQbvONKpYMhdSC9m1ecxY1SSvwLItIWQ
VucgYETs/0fQCpz+ItoGaTkPcjLmjm1PYnYDPMYz4IjbV0Rcz2aB1BHZE7D4TDr1
Sz/MmPQMhDy8dvldYJbX1t9DLtbm/c/4Uo2zydkSI3Rwt5EhAzjHsVaNXfV6oIit
sWZhRw/4B5/euqdAkOcBaiRFy4h7fQ6nFd6Z1QF/Tkg4vxGEPV//Nr9T6MRSvYVf
wrKogeI/XgrflCx2qS+CKd+IM7UTI6FYTHhN+q0RFFiXERt2e5okzl6DVcPs4uvI
AK/LNkV930NK1ikheJ+xy8dyR+W9Oj2qt9bR1sD+GEz1Kria4NgqSGVKDWkPNqz/
aJvPTZNkZOoyoQAeT6t14cehZ5P0fTuf1K1RzvaV07C8PFdSI5zpDCNidFOle+Nr
pR3sZqW5vS3tdK83I/tgBu/ruTAvktNEn4QccNNa2Cs5cIrnoe702nSytMCFfDYQ
dRhi6pdF5o27JU2FMUvtd0B0/CSM0D3Hq0Bp9/1uKN/fudob0VBxq1dwW82E6lTe
3X//bx+lwhetfbSrq6My0mm9ZXyIwNh+CDr0VTakUOJ5BoL7I3Zjyjh+MLcE+x9F
2fP3q7C8FTAlLjw70HwTBmLivZE2lqLlQFUxw+ehnbH8bsp3dU2Qt9sCaslhk9wt
A6x6nVrpDdkRcnF0dNdBPJV8Q8X+l0omlkPBEieJS74Q9VLqGm8Tb6MtLQmdNPqa
C1bhe5NHd9WbAAzIL950xR/idaU5mxqxDSDKx2haW5p5Z+mQgcwVF3v/FM0yoIbY
eRxHd4fyGgi4camiN+DZ6XLUu0zG3rga+PxmE+WtY8qsoC0XbFFLasLxPyOjxBWb
jgZVXZ4S4Y6S/qnEvXYKQyH7o027TIGGaVjPOQSFH3z4xO9TpxMtnWOjV5jHte2S
LmEAfSKSn0EgJ+we6O4NwqdQkZWP7Hs3/Gr7rBcf36P/EqYhK0b71EKil+53GPle
kZVBT+NHzUeRwZBrYU1vx08xgZDrkwWo+BfzlvKCLCdZaFopOL4SR9rUQIUW067G
pslEHEJd/wjMYf0hMJOqAIWV46XgGiSVhC/JUYAC38EFhny0SZQ1OG775aE8ZEZS
tS2LgMqd+HOhBC9VOQUAY1DbGBLmDBuaNUsZdKOAr4qfBOn4K16wAlMdCIaGeHtv
yJpMJxtjYtRCsl9ZXHx/IAr9cigUIzrVChzP4XBtGJKCPlmQg+lIFnzXYxl5EHzg
rJujNIbv5BIlrMr0TCDxrhBOLgecWMoq4ra6VjhRQZTduX0y84+vMf4AEoVNVIzx
7+44j0moOfxmC1yHTsHtXb8uut5ljeNWHpRwlsN1jK9nH5fX2Cz8BeDPDq46qU+t
9Aga80J2DypWWfHTtvI5z02MgheSfi3ZbviV54lJew38CORFPOhkrE1IB+R9hhmk
rJBno735kjt12H+o/GNI60EyYRLV8MF+WTSUU2SKVJvhstGJfGuCTZS6T8e3SlNn
ENZ6HOIkhBaJz0b6lsZiBaiRxK1hFF52hw61BVUIcAraKd3m4XFyvcvoO0AqxXam
IORgM9Rmxaa51cb6/cIyM1c/SO61Tq4m4gQoEGisGRTC5lUMtiohiMLf3CpZvmve
24aYC+mCAblQ8Op05+U23P/XnYegozGfnHfTCukF/PKd50G2BojFcj+XSWXljLcU
Xa6xq+FALglm+RLlkl90vTXEV5LIovNoHVg6cPaFCfqw9xNEoqdiSck69ZAUc3+w
hpFzyw0krY5y3OIqG62VXpBahA75Awl1veCh7Fhq3FoDZT7qViMw93eKi3LyaTxt
b6lFSjz49y6LVQrQOET8D2iaK/iTZW0bt1PV2FnYvHnaKCDhqsGnNnQlwbjZIxrj
sy+lgbs5iECsJmv45atA1JHi7FgiIdgK901l566qaArDpPgIVUBTQlBC4y68apQ4
tvATBymCAUhtDpNfgNrafX6ZNQ1+DOrBLxZ4D785eUlvr7O1AvbXnWTehJAKMNE0
blBx1WswzlvdJw+Ou3yEvdV4yfwyr2hk5nAfJiejN5YY1Q81cdO3lftgcioj6WqU
IE5SsqgiEBqb3V+OGf3jb67zJ4mKlM61WmVVznHNB1ErljHh+IHt6QKaRI88VG70
GzrI4Tc7gfI8s2pb6xiPfwu1FEp/zPSHxt58Rcsy+duSjx9LcUdTJKXOblL3NAYk
i9iTWubpcIXE4G3+hUCwl1dtFudK9yAutQPl+fIPzrv2E1YYHnwSPHAwuygesEwm
j8UbFlvJ5hmu4UmvHzL1sBTKE5G4ST/UBtCD051YxKXLYXjpPnx2j4HfaOQEfKoc
AxaqPx5aTalwLSU105uH31ILpD/7dQlBhn/zsvdsuFDjROU3f0bgUTHT8ifSwZOW
s85JT7oVAOAaYTb7PIywL5mv78zqSK1q+NYzdKtrbwbVGtaWF1cNA/NuvJNDT+Zk
xe7PPMg8od0MTqwquHyC34Pef7g8G+gf9Tv/NqYd3RR97eXrJrgtW0S6ZyJGw9Jk
848sG8w93gIpeZPVl806DtfKog0y18GdtluFzOOTMF16yK4VBO/MkJy5e1jyToAX
XqEItRLpHQGOJkpXrE87o9uNyo6VTzJBxcjQVlvBFtP3v6mpgp7PYDPYinnX9Pc6
KRmkC+HPjt9ZDPJmRDTHwxNRh17GLDQn0S/XPPchTkJDd3t8Hrh9uiGO/zquc8pp
6UI/k9ShKIfA5sSqolYO6bl5vNnYeBTEbBWuwU/SrNUhiptZJo4MJ2aWhiYYRn5D
ep83NOKJPmxVerrIdm1GG8U9QX12CiotjaxmQrzD26WuO3YAvyONU00AgZVDzdQB
s+PlP8LY+3J0yi0kA673t9TEvoQRmB5VIkyFaB7BYfXKfgjvumOQGd6jQ1bIMbY6
cRUVHLVo4ooL+iyT91kdAdTDTOKsIBXnJ/sZuPkEtN44fM3S7yg6kxWKXW9T3g0D
LiWKRRviTreFB8jFOKGrC3GiZ9bvX/wAocFW8jTX1ps6a23MG6xIEw1U5xr70zsI
BpIPDo6JmBM/+vYGiobJJ1z54T62MeoWiP82O80SsfxCXTIAHRYJ6xmM6a84mKFi
1kxACZIfM1wgjC8HmnXI9wrVraofQJePeMNtRVBt5dr7inyxMsgj20F/xeQ3/cyl
A4Th3AGI2Tbxe4dBHs+r6sKvzUjUU9DxpiQ3JeYDsdOfKtzbQwckjHnkspbsxZoX
audD04CrY988cjPDljFGgY4kEoxHcsRQv37J605MSQ7Qz4CKe7KvWrfaih0TYMy1
HfW+Wrpb/dRNx8n+2olnh85k53XRwNhsgC7UfzMY6dmG+Dtp4iSJO/2uuhA99TFW
10SIY9gS4AAxCiV6dZcU3/3w9WpNG3Qnuw8/80auOgbhd522Ral2DEimB9bAHY05
rou8nxvItt1+iXU50xyEv5pUG+obgsSyVov21ITfcadPHIV294PcgcAjsujy7YdC
qgyxaUN9hYLKGRrv/KHShcywrRHcUKs4pomSLgT4wmC2QXa1jk9gnNq36bCyxVXv
z416ZTpdZbwZyVfFRs+CW2Fz8Vx/RSyYyLtWZDwAbx74qSo9twaWtJA0PSpQrChs
ej5aALFUABvPtmucXMu1UyWW35Fq06RbUiEkFd/4mBsG8OxKY2euXUj5v5I8cWnS
JJb3PPJMyVz6SmKk1VvkVJrdk/ANc0wIMLWU7BfxOY4Dejp93EKEWg1PwZVxtGnD
fqYeDaT9TO9jsYy0YkmzoxqmUcG54x1pHaxfjtZe2GHgvyD7GlBkzZSBl3qzSXlD
tfPhS7pTIHqlO7TOeH6fqVFE/Q5WXsx299iihfyWzK4U1R8A6QBzU8929kvPzXnN
aEdg7dCGt7iNdj1/fcQBNhS/QOicY7N74F5GmT/Bhi7aI1AsLzmBPFpC+MPZrZsp
l7uUtHyAIZw7pcK6rPe/IButz3mhZPZFctwWE9w/n7fSGTX1rTXmwTCMFNGRBzL4
ke15a0N6/5M0Z/rW2lNwwmcq9lLd5tkJ+RRcvG0kK9RyRZt0Ey+MV9bNJoexLlN/
IeBA7oFujZKN0qlf2zt6h2g9pdttQbG2iLUI+mydRi4Ede8pXDFrus826/3uDguJ
QjCfcYnpOUCfzwVhjkpjyxvB3j3sEgT37/h4Y99M5P15ns1Li8mSYs3OVS0pJ4lw
rkZk2IlO3ItdwZ8qAV9lPYD2oyJMKkaGPtRigv/hmv47qmsU17UtIaSpW3xyWYkW
SVSIEaWiaoTs3WBhRRifC/s1whQNERlk7GNyLPomYFXu45nFdLBehDuQOOD6sgUZ
dM+Ud7EvLols5RqLqFHc/XMqimzry4TIX5X7vbZY9eIWeO+S2z+8mDapKsDTV6SU
Ov7wM7pI4yV3aNSCo2NTYxTcoXdXEB/jJpChtUxVLLBnyjIkMdssMxKRbHxNjJ5J
xq7D7eqOkUOrGuGAVZ70eIafsJHrmprS/+84ppm1pi97swp/0nmbjdaa3vCylq1G
Nc22Eagjmdv58HEuPURC1ocWh87EmHwzESNEMKoNtK/kcenPwdkcqLDCQRfcmquH
ePm/tz8voHYjv35idXBRNgEs2DqU8LBPLcw3Ii9lngVDVkJDSI6kFMWDJACd8zaB
coovU9GFxbsEKnzu75fJoxrmmYnLutv6Z9DkH4X+eUQch3Evs345dEOE+3UWQ4vp
nqIrgWJ9tWW3fW7UeuOlvQWDj+VFVDMlez0vdbQAu6zgmuj1nRfNKep/sOVeqlGo
FOJBsXZlU/s+zKTKa/74IsTM1LQmfHKdCOGPjLtzuZ33arSzptguD8xFZcNv76u8
ihSyEsRx10TazBWzxD0DunOegHp1KumKTX1RwjRU6K04Q771t8aFcDQ1EAruTPqz
GWmyFn0+ywo+Pjy8uvmSr9QD7vl+JCyfohu/XnG24Oq4XzTFbf9QuuvGJi9Fby9N
D1eh71HhmkpzDnjboYAliAuAg/QcXAPbRpNeno2cSRfU1zOiZlZJ60+FbuMIouQT
8LBVhopb1oRpnQNQmHaUSW1uxZtzwOW9QI9szdn5M6q1ji/2vtBx/Uz9+rNW01st
2FZ5gDI03pRq+QJKlrrKoUu7zZrjLo3fUp3MHOhU0C6gnGFJOtOqaPoY1hhmxA1w
gHaL4f2Zkr+pTC+UjkY/ifpWxJZ4KxbKRS4pP2vAB1ITYW4dkcjQz2VkOwkRnh3O
T2Yc80ysLNQnDonFkjgHk5PH7Qd38c2TllW/o37rqyLhYp5lpdtaoLNusPoy7CMj
/TpY8jB+bll2kWMQ1I3kouNJffjLh0nAf6g3hq76iUujoWEFGVxfvurUKbakLa+t
N1FaQb132grmc3nFSK7R/glcogqx8LxF6ScySZmyZ5pdzOSdNVYDtq9m9Dg56GVz
yM777n9ZkhJkfZY1ji9hKdiVVqZZHYCRmKZHBi7RnVTB4AV8pzajhdJDIVg6yF6F
Ep6+r/CE2svSPYy1GVpjS/IyHd720Wr52ZozFox4Vxt5Rexuc3CE+Gf7GFiB/PV/
3OwHXflX50IIE0+F/QeRyOHgf+x2SOiZeiVx22rlJZ5Pjr5iNX48jZlaGZ38PBT5
SxSaUWVpblrY+T6W2zrhagL3fQztpevXuluMetTryBqQHhvZMikiQjpCLUR9BZT2
z5cM8ifqUJNIprYDfSW+jdeQN+sWlK9zl4RhzicGEmU/ORwWGPdiP3dEwOZ9yq+t
gYWr6PxeTGGj+x3ptQS5G1LAl1lnWpRnqn3RA/W/+CwzWS1yrqHZFfBeHRH9preY
pB2h0UD2prcMq3tt5buhiJOKYcoTUBBVT/oTS+RnE/tIDl/gIIrVaPSHxBxvmkmH
NZze/MIh8EbpBKmPHwSi6Kzv+Ym4GLGI0RAISrwHRMd64Mk+Ru4UQ2dBjmBeM8Qn
4qWYYGoVENYLXQZ0TPHv04fdJK43Wv87mml707jFhTMx5w9Ci2E+xNLAkGdCXq1m
ZufiPymkcAEqUGYNffT3X64ViJAsI8Xr1u1Viokk6GMzhdFg//rlCcx7vmumdr79
B9fUwSc82BdxeAjwnoW9l9l1wAmRNThjF6NU+5zt/FDyUVF537AnjZim+jEaS5Qp
51NLA2Wovy4sTn1SSunLuORgpqKlvniZwVbLfmOw8XK/x4bMoICaXx+uSUwCEHfc
YYwnj1D8Q1nKHiCQj5ZagNHN3eBlvm3M6yl1Ymy2Gai9EhMuBKU8uctx14YSRduC
kaduVvd2pJuON6fPwKlsXQVIwbLiSYIq8wz/Gts2iDFE6FD7p1nQC3xOF/geUgr8
N1BHDOlPMlzVlThjHBf38+ojtsIv9NEr9KEm2qyNcG1jhqj/YGDjQKrMWhJLFnfZ
Z57ohjrv9pZDTq2V7/vfxUkEYFPhjKj6DBzIpaE+9PlEyvIzFKO0kCw2VNozByQM
3EXnag4hhiqGffr8jRiUn+1uhb+V6ZZ0qjrsLSjzGo1slo3VweYqQ1VZaNQ5cVza
5OaOeb4T1KtNWGqCUCVK+88XvqjlB0N1FNxh24aTgqI7Mjtktd9GNUnIS87c2LNs
4Q6ThEC4awzQnCOIdo1CZkayDIrDaICXV30a3QEpx/3jj6rgHTSvwoeL79NX/i8Y
LorUY3N713hcfkFa/6gQYiXdeekQnpaUJID/9t5oUz0kuwuU+9+Hpz96Umvyvr+R
7/sOV6sh6q0SSreab3VppLvbdlnUSd4zE8aMgl1FPDszmjaog8Y1+y0nbGMm6s57
ZBqUtBC4WfL5SCCeUvVEyRl0ZPSmVdMXhdwr235pbbD/jSxVORec8FhSVmIQeroy
o9U011f8YlJzBl71hjEhGbyeM5WtY698iG1rBHEeinokPd7uJFkowpB76kG8HgyU
vqOXxB/Mff4GuRlMYMgnVezYO8D21hx9xV8PhJwFgfZ6stYMiPDxmeVpo7UYv2E9
wc2mV/n09o7k5QlCc5QNHQtdXqeHlHG3AnN9xr9snFdxuR0BZeZ/uJeYH5iT1xui
xnmIsPiN03vdsIU9ifDXlKJ40kKeFWv7fsBCICVbfQMUWDNq1Dz7mUM3cTY4AhVu
Tbmdiobc+iZRagLk10Op/Wi6Pj4+7mDkoZXa8IHToFGTpb6kmVwe64NwJhLhiRYr
GA9WqBVfjv4W/lE03OtbDO7JvlEeUhE19TGRx4PlPBJZavtld2EjraFveLMqtJVr
JXqHkVEx2wNP0AI58P3dwtqYVmVG0U/0WAXPJ4u64nhsPTc4ywWURfgMi9jKij0v
hNP82TCMuNpj6mgtiVnTJWRyVz1sFitwuUl8tpGeA/LG3jJo6ZARslFD2t5eWH5k
d6sc7xXxF8pDtL0XixuT3mXcnra3XCaScIMWs+kgrLEY2zIHDBupAJk5J8xoo3xM
kQKROSJyVjNkB6mUPZiOYlwONTpPbHI2vLVwJXi6ASG7vrT2E7M/ZaQULp5RHkhP
Of8QhzUEdCYHRhFZI5G/jKI0OpeeXMpxd3DPC31Rd+8OWovtysPGiG3Ve2FoBhPd
D3hZQ75KYteBAXbXCm11EcGX28syXa0u0HlrgiBmnFZXGImIuWAEyIW3HAySm4CV
rw7XOWqSw0GGCT0LuKf0eBl04trNpZFHNTb8uR6mjM2pEfJ9rboSBPOkhSYjDJVQ
Ye/u04v2TsBqMRnhW0n3DxsWFtTzw1v03O2yxWruMEo3bvohWiLC/CfUKCpgFqTf
Fg+d4L7QD3aIcspHwJirSprgQakuLI8AeDPJ1Cpnyp7sryhrPBo/PPJcTpmWTliV
JKu3X+UjlcE12tKlq4eSyODS3BPgscRXh24As2uKrIpmoISiLC1bgT+Giwrdik/H
OTi3JZ49Xr4L/auNlZeQwXKBOS1YRVkr6kMYPJCpFT85vT/oE/LA8fGI5u7b73Dj
kQKvDIr3453Qwth2yM8yzTwh/g8amkq3vCM5Fj/B+sw4CWC/0JcM1KiUGft2jQ2A
Wz4SZ43DbukxF/7M86tBGNYKOrJZLhqUzJRDbJdtp9Tn6ym2GbDCMRhUeGLUzQeM
Efyo5hOEUfxP5QSZH7WlmaDhKpo9GnYn9T2QlOK60x7qZZ4V9LjJM/ipV/MS0ART
Ub4IBRpTXNqKlE8YsAS6RAdoAvbzGxqVlPQ4HTM/PF3DdxOC1Y6Ec/uUZM8vG9gJ
vcZ1VKtdOQKGYsGev03dUWItfl5nwMwe8Ibqn04iwvH7qW7KZ+GSqeGKAuF8MMDz
v89OMIIFaHgAiBcnn2LXXeDPY9qZfx+TUIIJkc3f74xoahbcXCoIDUdugiLYPnvi
k8QHYq8ldf9p67U2/cdXT+UGepD/H2ezMSXDy8jh0szMhJh1wQMNldbVhHxjGMVg
RUTszLqZqKIK4pyQAXTOt4rr4Zf1spM5OZd8n3rdg85CWfxMul4r/+K76JArTRQr
lxV4UiFm+7F50ZocTIjgj7qChZGtFmQz7lx0FhukuOaAfZCNpdupnbg3GZRuzGRb
67FYXtwp1KkGkCn/24CUYTv8YVM6PcY6Ik7mSNXm7pLEjVWURyGnvE2XDpny/VLo
bCf11MwTEDvVxmt74/hJpQ74sHWz65dhRaiK6QtHDrAW5jFmt/1MGwJ5qnvvhziT
Pa3ozJsgkTi5gb6w9QcJWlFgOG2FzImm7JZ2dVfS0qaUR9TusLMZ0fHsjM8xa0P6
FeXKFTBQEX0r6gWQocv5ztsT+CTtYuxOdnlihStvNZZ774T3i1QDZ+Uv9ygtiFF7
rUFiyUOm9IsxM3EW+Mr3Sz7r2Uv9goAqxJOysh6NPmJvQ4OobSReIbMoPdem48NG
2H11WStzL0GQMqqxdoNB3aDrhF6Hgd6oI9o0eS2efhkgzY8bLZ/b86fb43OQ2p+d
iAezE07NxXOcBw5kX0huu4CQLTDJE1Kn5nNO9W0wmP51Rp1EqPdNJWAVuDwX0Uu+
34AQPtxxmocZJmrwFMUHGCgrtClAmdoKQMmvyNL3uk59iv0cNau/5P3QkIfJ3Sqh
niaEobhRl2BLq8GmyTUr5SFy3BYBPxFbxTuqVnd8v9aCu1vFsJomWtwMYVITqtmM
pJmIkO1s3sZs/IVp2XG9HXhtT0/jw/v1MZhz8HzWvOu0TfcM0rb50wd+mREf7k1B
y+00+WT70VQ+x5gDAnYL5b9d9Nu0nUHq1nQF9QKRuGZNbtsvi4cwKJIWl9xW5qeH
XLLu8bNuqViQV0MtucyOd6QaihvCkhq6Nu66KaCnTXcLX2+UGtOlKx5JLDKw6RB8
HAvHsVY9j6Ct7L5Beddh6bRe4nJI5GoiLFXAi56LlzIOb2TYvaVnu9SI+UUDDbdC
T/+sOmHCnBUQyopbvrsL+9XFxF4N2oVthiBFDxu/Bq1YWEkER1DdBuuInRAXwGU7
GwJW3izHAtjZ6FiZp3vKuo9rpr9z173psqer2pWDzzJ7+fXcg5RPUxtoZkoNhUx8
Z77dd8R1OKx4o0R8Y9FLk/2GZVa7WeWWhxQKaNBzQn5CYPR69mDZ0UtzhFzn/ULy
xyAgIhbW5XPSaullAM/8DKYj0IlwT8UEVyjT5TnAHecMUcDZwowq7QX30orLEV0d
K6s++hm4lHgHgHpcetFUUUNhSzpKfVNwU888ZEUFiKNuguk8gX4A9K+0Prkvgs0/
FjqJpMvhcOnxse8JCPjNpda5SCtq7BMInYPOAzGt+xMpvnmX7JXE6ccb2o4jo+I1
2kVQBj0y5v+9ZefFoMw457NrNY8QxnI0lkE4kifmol28NIoZHDVcomYOl4yUtne0
ZojMBsQg/lqBEITwL4vjiNK19Adua9tgbpTohj297Ov8yE1reueD1FIaj0QwWWMa
m8OuLTeLqYLgZu/ZKuTVIT/HFZa+vp9W4ohvLr5sAlykd6ZSVoszHRdnrx8Jv7A3
4DNPJfd1BIW27REH9ZcN4E41Xppcat/fIGKjSCps7mrH6gfF3dCSxgdh4DELu6vG
w55DHhAf5r5hCVU5MPRB7w9B0k8T8l2VP9dnZyVUaMgWwAbAoW0ukp+unXEr5Xig
ydoeGWGyeenXWc6YNxc/co1ICyqGfQna+W3Y630BijAOTCLKpj0jUhGul0fZvWNY
TZ6ckWXiZiIizpXywrCDDSbLE7lMcZ88RMybh+KX5ou6ltagqDIpjktpxocQLuBg
lLMZDyybZHrW5c0hNwb84sqZVwR8/oYRG0SSh0q9FR6FFmbrpLdLyXLHPL1f8Kt0
dtuvEiE7ltszE6vd9EJkY5HMv2pLXPU/pAAHV/Ae17xcZZxFQjuu2/+nWvQb7Hw3
m4ffwee9F385KCLoSCTidZOHZy+HRVzoEpsxChWkhzMiA17jHy3ZZhaII0V5bNsu
I4xBS18/xI3qgBIYqZ5v+7Lq9WJSChGGantfilH+9W4XTS1B7GdBtzy0ImEbVvz7
UmMdsdQPZ1ISdq0DurhHfuouZ+rnmWPVrR1fOJDoa9kZBcxEk9aejAZ1Wo/jQuRk
FxPGhp9IlIr0RymvgZrN68ico551ZgHwBTf1Oo8GsSgz21IlqEXeymwVZcGtsTP4
FcPmIm4WXyf1Oaha1YaY2/0r1MdglccwWRhUcbgam0Hp7iIUmRc3qEMwK4+EixcB
Ab/wT2TiVkem7iVmBCZD0giJ4zKEUdT8jajlM2henhPdF3DoWofPOUCSPAb2SDDy
1ZlFLoAzEzTsKC8T6jm4JpP5FFBCbBDLJ7GZb6a9kXnhQHknADVrQZgBcYZuSM9L
166xgqm1GEdb/J+19k/0tOdykUTTR/X+gzLG0sa+y0iOxHSvjBfgGf1X6J6QG3Ur
AIZGgwhJW/8kFXn33rTJHYHhvA1mn0k58X3uMOKhIPlfrn6hueMjAdlYlMq+iVJy
vmqTSKNuRjDzwQ1GHqNewq0teWtDftbH6ixQKdj4D2IyR90OYLNkH9AeG7sPDV9D
oogZhpcRJ267yQp18SHd6AIG3BTZw6q1+fdxFhFB15AFqTP00Z1N6mQnxiW8mYOG
85otohTT8UA0fmoC2AAUnkV8Di8YF5rdd5RJ84chLjUaRU+jDTiP8iOhB+4Lti4L
GqB4JXZ1bw7UtW5JNyUGPF1jOWLzXaHLpB+tfzcmkZfWz9ey5Pe7BOOi3/mbPt2w
1PLh7HZJIYe2WWfm5NwM2xeDTkxbascl0K8k9CxfPhl6ervmF8nv1GLQHj61dXsB
6eVGoZ31DE7PwkpHJxs8I8nlGdBDQxTcW7+h7PFxHrB69jCyAaAREpc0bUx+dCiv
ytLQL/4fIOlewBrpK51ZM17kSL1ItylEvqRgoLcIzXPr7+D+2Zxfv+NII8DrJ0gb
3AZ0/f3/gGEvDOhsk3IRak+kFVA+sigSKZ2sp5LbFIB70o8INIyy4r2+nfvzrr7j
i4MnskDwouG4PCPALltR+2js13I7lploPLoJumTmYQXoAXUVeWw/EJh1NepSF67F
8tN4YkG6Xkb5j0f1A1aWdaac2I6MqsRy8thyytPKTGg/GXmQnXSEqQ5d3rwYYjL4
XZTFrX+MirekqsxaeAZX2kwid1F/Hr0+bnSpT7iY3ozUgDH1nspbRYwSl3UVIz14
ac6sLzbX30fi+zw+xsoYctmRwQqwR9zUzdYEDwXGkWm2YsMuXzAI8yHTh3hQ4B+B
MCwCraYcagc2z28CbbSWRN6Gso543w9hEB3cB+M/X6jmZmZsaLxqazvAqhIC0py/
bAvvt3KxT3TE2IowPzHElOk5EphbrpdDWZxLx3vZbuniOz6y+ANqctWoMukOzb5F
GUJAgJGv7hCL6OfeIHIpVS5LP/wFNkmaVXlwmOx37ObADoVH1dIEa+2idjLzklHm
9nkFlNzK07kHh3DxSqfqCsqATS9QtqBAjigebR7MxKqbVSaWBS6dxLXVNGOQAc6j
oVSQauTOepwGY7iH6FJmzk2rYPj/okHuo4HT+mfyUxS2wX5gz7efa0MWcv0jTpts
qpJ72u1VZ3KyC3X//bzxRM2UhY/gfD9jwCR7WW1lpbtKOTsVLGl8E4MCqnN5sJ3F
4jFGNrlbtd3ibSGcZzQDEVxbL0Pp5TF+WP0kTPA2zlx42cMVDQ/g8u8wq3rpXt2i
p2FhYDLX86K1wSomWpD+hIzVZ60XjcvO88sdyOM72uIiYoVyvzOP7d3I8i8w/Ped
PATf5QW36UQ0OU7lpXf6zPl5iKehSEsUDe5pBvEDnYp0i6nwrB0Xw/p1sJjzGYCp
eeh0g2F4Tw+A8fYitmfwNGCnGAS8bssdOcRGX3SETafAQHXOioXRgwrRBgOcbgqC
lz9laIadlArR837xUj0SNsEqfmRP3zXTmV/OiWlnGYRj2ogTdXinxb7FvyzDnD9x
PbNoHk8UohW21ainHgM9SIT9V/4otqODi5eozWfCzO7/abdjO8dCIT1v/kZmoCMY
DXFNMIv/O47ldY+o8bsd/4ArPWMsSFpa8AK6HCfTk2SHPybWQtveVWjmACpd/3OU
paJ7cb+awRECJ/AN3rRKi7p9fzJsf2R6ihymQvKI8rwk8tc37a8xLyT7kdmQ174J
wekDtTFD+gBEQDotG36bMnUF4VnLvnuG/RemOutG1I2KN2IibfJij1LH7Noaw548
rb5BJiRK7TRbxVlIfkZein72da6YiTOVJ+iHR7bQCOzdSZoqlUoKS+xjCPZwVqZ5
IJtjSZR8dydGuGOxPYcKqJ34vFuiDIMZgWP0FyaehXQ3LaK/QTAgkTLZgSYJQMRW
KdAubfCCpNayZHY9vie+McglDJeCTqCVp0/vLfqpApwbpPJmImAWaZogbU7cuRxH
Vl6zUWW2z6VSMuXwzN+rIenxjE9I6T2WPLVQfWChUk2hSjpJFUO1Ut09VcZoj/89
ncczDH5LY2dwMw6OmUrmOB+BCFnAtkuy36+9u+EbpBbeK0sh8iJ4zgKRvi2873ow
+DdGpQA31OSYKJ1kM+tPxa0LLcWYC8fzKwJ5WZ2iTmSdUlVQ7GWtTMrCtNoQLpXQ
8gjHNnwvM/BQt7DBCQCe+f67z6GzMVmcfAGDRwdoMgbcFGUb1jqODZNutD1gAK/B
+V/Y3FoqmXFXhxj6niAOtjv+fFnlnqf006JRV82AD35VMAbnjx0pDQUGafIAvkqI
GFCAXNnMfJ/p4DdeHCo6sBz7f9to4BHfeaOV7fxR24y8xewPUaMtONCd5hhCkCKJ
fh65bInQzJkr6VKaKTZq3JZwJq1xWKLUNG3cWs/6PcA/Wg2Rc544/g6G1nj/brzS
mflIOaDwRsfMIXd3BsVm4UDQd5fK+9t6u19KnU/ELpnGdbRi/M8+4zzKzhP/0b+K
5VJ4g7uCBIcXf69zrQipwNas/T5+CKl7efPAVTU1JppfZSrFu4SI/SRg79DpoqPZ
5yrqeS2MTBsom5XyBdzUn2gn9bpDw2UF5EM29FOen6pDCBYvRHoKdaItdiyCVZ8E
DGftHI8aC2yTBflWFtHGbR0/zbFVv6gVK9wmISL5MOU81NjSsmxKR+WgKlHTDtTc
nhKXD2Ows78mv2FogDRKf34Cz/m85mutYENiw+yx+1t3tbH5ev6R6GSfKpAcG2RO
sfVug2D3raOjOO2keysIeGORS4c6DE9Rcn6JblIyn32KBhxq9ODTwo1kIPKVrodT
jf0wxw+5ZPagO73pSKrMY+hZedmE0G+1bjGYmSip8A30INFSD4fzLEI6wokyUtJP
ahk0MOG43JFQ+iKyyRmXJvDEsKOtR2F7E//tXqh/k8NVv6QC/7nh+V7H7Usj+K4H
VenleG13FvdpYjBHcVCwzy3+8b9i7IuGHuIKavTwgOfnUE/Z0zlEAevYxm70r3cL
LxECJ/M2yJmTsjjZF60Kgc3jjKg24nVmKYLSL0F6C4diz+bwrFpkA0j/c1pr+NGI
FlpYSld2yK6yVCI084i6u+tgJ/IyE3OQWS3c4zm3H005R3UDkKpfKsQYSUv4/i3g
TeWppANkPqmR5JQb8mvBBLegZxx6oStTjecxdRXlOKX4/ufbFgEHW7hP0SRJbGHL
jSI/qsVC/9aK9QOUEyPZzM7/eahbV2mpzhiE91xnkeCGyyoBbVszrfJM09uKmDmI
UaNuEc/Y5YzmWGg5OAFd2pL4YQsIrywhhNq7QfmAQnCoCiqxa3xXzBUPEzle75DN
BMrEVNiXvjv3EB+AbrvfKXvir9PZtG5Zh5dgn0Oj6KwBKKxDmG37s97zn13Jkx2o
RtY4N45HAvUVneUuDNcGHrFL9b04MHJSkZSrh3m0QclCV6yN0tE7+noJ6UYk8Iqu
rW5jxXKCCDnSteM5q9kvAwkVV4Vs2dFHPheT/U4GlnNU5ch0XsSJ80a/ZAElBTOL
Ct539j8UYT70O5vGmbqrj+ld+hF5hi2abr8U35GYRB0nZHboMUAGwE55Cqu5exwE
qJgCb8kUj0X+n5MBMdJSG5rg/ikqmvRgh3A85ckZct6A4OOSDgFuBS4LbFNoctl0
IX4OGSUg4uF27Vbgs44wDODLPrfrYlihKpr31BiAAfC0ATieDLmUojvb94TI4DYj
Pc1t5rCmQU+572//lXgnU99Y31YmhAdfyweMW3fEDSV6Hw2hQ0txG99rBjpykNO5
Go2mujOPueKJqQDGQY9W8jfX3xC7but7EENfHtk+2MMP6j9shtEzv6sgympfg2hX
qdwAkLDUBoYKhpDZF+sTxm2JLpx3O+EQaioSSYIfH2aNgMjA94hfezZKZEVyRCTQ
RyK8A6fmojt7Ui3WvfXZquGJijtrTbZ7khI9WqHeWWWC0BgHz2pE9bwvLwfZMboH
/uoTxvgcgLO0nmxJYjiV5bfOSnAo+2XjYg8QlAffI3DvvN6RWxUOGiW/leyk7UKr
XCzTDl+hrFzRMmqlEfieQVuoomoebCKjOiHKdrxpRYdIAyWWQmSrX0uwfqnDtAAg
nAQnpQ0WHbCGGrSzDyHWGhdZtOEPbJsgPPRhm9zg+8qqNBYwPI3UXJA1/jrkkvg5
arf8BCJIxvqJPgg67W76RcE994qHfTzfaXMjd/aznD7Uy9WV4J6dubWRVAYvOms5
RYocYsuDa6WdlsuGwoC96Mk4mYSIyETazoOuEKtsGMty7Yt9xXCRiO5zgO+otb0j
YRkxr6n8t9RjQ5WE5Og3fSGLbsBBS1jjf046TCk6eUa+Fsyjs9I9QLJo47ZMt4Zf
e723xbZjRpat45RC3H8lV0IIZ8dgGAdkPFslAojQBGAuFV3eWfJmTDW9gTquAdXz
4iygEM3fZ95ls1ls/qZNX4EPhwX+GqQITAhFh19PaCnat1a9rY1JXyQZNdZGh0yl
jt+seeIVCnSQTo8B8B2ZUzMIE2dryH6SzzXxStiFcbIGNuo12RnWrKByZxQGW2O2
sBd8Mt/whPrUMGC2ZJHsIBnOzojP2oBB6DDYyWflbdVS4sgpsaakz9CW19o0x8Gj
y5Z4ro0eOnxeq+oNO2EY8+pBLvYCXFfZNyVQtAr5GRq+51000IvRgWWgFKgdbJVa
jbeMDIGxVBoU/VOfb1zDEEKVSFV3l9AcrPojTLz2hKMrQm9xoTIzaNRRTBFbr0sj
kZdkrwCwn7yaC8w/UGhKqdYKG0esYVRz3FZZmFf/wBLv9y6Ks0Ze1Ugya/nVtFd6
B+oujnNwLBIeOAJkF3nwslprUmCyGViD9NrX41QKYFHQrXW70rFD6DNQzfQCjQxm
Evgj5FtYiLjpJxRM0tRGIg9VBLP1aZ2ayDPAuDYUm+xJEeMXjSoPc7IBA93+US+B
T9E0TV7EryvAVHLNriqwS0XKVzDN6jzLY3gmU6fEgW/7IS4TlQ7NfECwuSnEjHNy
9tFfsOdQP/l7AaDFqXpYHY0CsAWE+WN+KZcTHTnA/qCjDSPeEshGny8y/gt4f48M
sEB7CaJaTvisACXsUwH6+JPQ2fph8H7cqVRd3CckLWcj3DL3kBwJuIRDawM7RW8e
CSIoLgHwcwT4fi4bf7/csfwZ26Hm7i4Bm53w0swQ8bxRFhWNh/D2pf0Bch0eXb5A
6Sm8uggFQ2WbG/ScDNItt7p0bAfJBeF1K/+qS3pgSLZK+7vP/zp1nRc2jv1yKwZ7
5xV2k4wN2DrWthAPSseUVjAV6ku/ENNFSweXYUS64ul7r9L9k31dsmAqe1LeiBnJ
Upg0397gObqxzHWsOJM4bF8wHhJ+zQIkhyHIHM6JXXa5/p7mDJGmaQnPwngCBio+
IS6TRM1gqCwqq9qGsefXjcaGSJUl8EDsvCQaLSyt/LUnVYEb7S5yIoZ2rru0mi9+
XaG6nVNDh+vimcW1xzvfv4/zDDizglBOi9rOEaaVtaICvXEvd9HyLQO3F0Ghltle
us80p6B8nnNZCoVLyQpiy4foGOIEmGmo7ib629wkf4sLWoniCgszuJDSAeY/Q1Ca
i6pbbxIOT2eavSt895mJIyjMrfh0cWWll2eypl075cZ4CvYKjtmeUY9ZSV++vbE+
U7m5fo740Kv86fp4pdGT9lSe5Hcg7o35lpIPQMHfJ5JdQXJYPNhrZt1h1Z1oCT/S
DkMOws3LGwwjAPq1KreLsPIWxaiC/zECaCLpgvOROePF8UQpz6pycU5fKbdmDVuu
OX+z0qaTm7rEbETP3ABZ6pG49Fj+jtwSpXrLNEk9GwZXcMA0vPtIabck9rgchPSr
YluO+OTXdUMkB3aOf29rjaGDj1LEl0t5qoLelqTCkIYATYL6KGh/u4CNN+yGUvSk
H0BLmUmu84WRpMAWtbZc/OYgI0+jpvMdA7iEr6j202TogC7ldiN/qq1qJmLA0tfQ
xu8T3Og3IHIhg3uUYnscSz7CC4eowsXR+lhgtLLegWeVctKjwhuaWR7/uLbRASk8
99EJK60p+6K8AknHPYjInYcA2xjR+WmH7HcVCkzsaH9tq+0IXkXNMyapqzDZC9Ie
F5UrdNIFbU3xrpNP9vuM+CtuOB2T6ZDD4ZB8FFWZCno+x3MUfAeeJZtQLRlHfLmV
bAHlLgwrzxMT0UJ12qv0zw3ZFs0MDCU5oi/c5KC0+Ql4XQz7rNfTEtyRabVogaRd
Mo4Q0rBJ++eq8M7LFMJ6F5CeXFRVya41qZWCnPQIO9avm52jfEf968f59QQTgpH1
FmQ7fig0AedfOwWnkcVkVlz+Ag0GeF4kFj138woSbE9AOfhXNFWVYMKApOXhiX/P
O/OrTXruh4ekt9QPoha7UDd+vqWw1ZndQO9eHKVzILi8pqyhvdFRalDKxOGhs1PF
fUoDtzpPemiLdGNigejzuJbor+aAzdm4Hua5TqkLv1JMnfLRSUCULJFOv4kSOguu
dfuk4/UQrAmVs84oBsg1+zXhUZT98wGPW1JWxq+/fCMllfkavgyOjVDmbn4vTIl+
bxMq8MM5gg/VNWnj1I1lM67gg02lhrPWs32nOgjtBRyrwv0rPkAIPHznguTnWGgt
lLYpB6OKD6guz1IKY6LrWEdQJ/aCITcLq5x3iaDrSYylal+oGq5klvXVxjekXbOJ
qDwdYCF8d5Re+kNf1HrGnP1DpeRBgOowSu1teDHXg2QYgspnFuzUQZgzeNUEmnjB
H4JQMHp1u4zUhCQF/SxZQoaC4X2WAI29f9RkMUkKevdAJf47YhosUU3eNKojCeb6
SWtLUjpJ3BNvrnoUA+QVFcUg5zRTVWpuIYYy/MBOcO+p6oE7V3UbgsdfEIdKlvle
kHsE/8fUKRvvlCQoMJxuukBs6la90Q3BzTFaImrSDo5tivFDzp9aZyMZGdckpLwt
QVBpDeWhrO0sIJQmFeyaWI+aB+jhr75PUrofDAfkxBw0hCTr/Ju2398kCdoUGCUM
JIclbgVZKxf2pmrOwEoHYAH6vCsEmXiv6p/0sYmy9fHT6D1l0AUZhWcLa5dDYS7K
3qEXFZdz66nA6sK31ds77xNzy2Wcl+B31WCmYZQ4anYJIiiiJENcYelgO1fgSSzn
3cqXhJQjEoSSnQopWQUyqaqbDII56HE3xN1lPXzeb9zJa75vrQJ2rdKGzI88DE6z
5mjXzpAGQp1mcq/MC2JApF5IKAY9lkLmHVF1AXHg6E7FtZtgcUN45A8njrRixrg9
8F78r4Yate/jGl0GhM+5xvAF6quvdCmnBCSYxEy511OHrjv1DCIHjVWSxI+P+izQ
4+mAmHjSjWz0fJvBrMVFVS9evAAb8PljWTClYRkv0cZEJ6s/XUT4OgPktvNN9Aq/
hNrXRhi2y3gNkbVVXDyteVCZlxncyxhNtiyU4jiRAkeXdHpcdj1R3+pY9L1CsHC5
UGl3QzGsIgMR10NFsIqjK3kAcTkNDsYg9l38dz3hdgCWH/EFiUMoReYqZd4oC0Da
/drnYywzfhHUWGYTtXWBWLyH5ZNcAw65F3QX972D1/dWLylBz60ndvwm7GjhmPdc
OkrvuoTmJohbS0Yd+V6LadLjEZJhZ8/Jx0xNK8DOpDLLJW1wg1VjGg1F+6ejLenG
5brMQXB4nXCkAHUNfISbnhwgrTw6IC9mKgXEoHF88WthUBnU7NxL1QnMCD6HdIAV
Vw3p2akKU+k595eOHfF6CxxmwhDPAoM11pZJsRsakuz90XRX/ryph/lDC7d2zJ8a
uI+MF3pmNf5BQV3Rt1XXCpJh1FdoDRyY+iC0qX61qRiBi4loO6lS72P+z+NfHi3O
S5wA2A9Tlxd5CPokDPKWm7acTaac+zy2JeOL2pvfOX7E51AZy7Ge/AfVZxtCsPIe
fuAaSWaS2QlmhuMlx0+X+7Xq6GvpxhWU7OTSd+kGPuaAbFKsM9J4zhkZTADSFqT6
t+FhBi25GeOVggOogDuqG2Lk7xfTOm30LCvmatBDmEz213gYx0dRnt7tBYUixoxK
Ll/ogrsOYqn+6v5hLvnri07aRuQNRnnkb8iRiVadHzUWFBuWK6GHfr8MeALPyiko
CRt1I7PEhOkmNnvs8JqODB2OC2vYOg+rSngAoQnWePwJ+uMiqYoi2HBgOOUr7BHi
eEpAH16PZnKFDuykPtNdii2vVYpBCMVWWbln7VfYXqWsZd7jM0srhVjWTofd9jsE
kmTEkyktw1TEDIlBWcotFKntK3MBlcQPs08+uHgZTKr9QSrQk/q5YqiUVCqy/j25
fAv1IOgZSWuLWIJr6ySIB3z1y/mIJBXnLCBkr4VjYStEmD1oM7TED0po3CYVsWGf
JoPLY7JdboTOtVScHMwEOh4aduZItMPbTrQ8wDgDvZvONuB7dbj99/4F7D35elxN
zvD0WAITx5P/TkQmj14dT+MUDmk17SjkJIKyoy2JvhDP0oV5STufHM/Cnd5aBwaF
qQKSd7NZvoOgkx1u/kYzf3LV5EW+GKCIaljAnLO19UK7j3OfRi5ez0l6h4fLP6mH
7kO/OnE1Y0c6EhnMDFj2HgCILrXrM4nscdYm6eqKHwQy47nmjv4PiJmsMGl5lpRm
ERXXhVdyw+g/OZYvn8PJO8uSe0vgHNWvO3FjzQCU3rNjxlBjGr5pzxAjkFtBZ1F/
Xnob4Iwk1lb5xmuaSAP/355lPT+SMbrodv81X6ZQvj//gmfu79Ridm5P3jeYhD/t
WMXnzGNSmjEkDmvYDwK9jsEza9smnsExNUGMHjcxZoUe4QR8reIO6GfA6EAdV4qj
Xcm3hDRhY0fjgr3LA2beOPbOUwUJ/Srtmm9OhLyXCccC3ORgMSiRgn6nFZXG6uP/
LuNl1g3lmHa7xuD+rPnGC7ceDFlKOpUfE5P89QfbS06/G3q9QzZSwl7osny7brm5
ZUPLm/YMqRpgsqnTGTHnJ4ElvHcalLVdtA8x7cBJExTztQM//H3sohBhUiQ6nZ2q
MOS/OzqVf0R5XNwf2ydQdO4egp6qddXIK0FvROUhIH+bu20E8EDvX5RXn9g2Uu3m
CBN0QLeEs2toX/BiFN5884r8CWTsX6fBmr5iPgIHhIvDMzyV5Xdh/KUoGDvU7FTK
v2xtxoIR7HW0ay3Smz1dnb4tCBS43LDYduUMTp/Jgq+3Bzm2bcHQkX9RxcRHRHs7
Scu4csnozS6I1OpReNaye5MmsNzwi0Gv8uERS1SBx07VAX72zTJqwi/qa8PPzPZm
o+//tqIIRaYSHNAtaICLQLsi1kg00sCn06P94SHy0pBWD/7E7A4wHgMtje/lUkyO
FGtsF5fd9/ZAFxrtBWVekiLP80yDmJHMV40MCmXzdDlerfPxxcw+p3KPp+HWyOpV
uDhN4xmuOibEGqFCPZGCkE7rNRgHyQkZ0o2gR7pWnB33GsUSle8Tz/xMuPgSB79j
8IBhs/H1fkToQExyETYRK5CW4fI4SqGcMs0wXHRhchBtHJdesKyG9x4Vm1Of7ufi
ou2YOelIvEirZEmbcohKMRZ4OMvoiZDnItvvc7rWSUXZ/G0gGg2a8vn0E79Olezf
895kVEAYuYCSyWSod0RdSVzfyGhmAfAlhmgIZiuhU+A0KqCM7hbLfGL4gTHcwafP
ugqbz5DeMsFAw2yCjOkZeUzc2PM4SzUdJHATEWRvGWl8/Qe1+IKW0pTr3JW1HFVc
WgNelNhOwQ23JC5Oo73sX+z8ArCAQpOwG7frLVpNXzgWw4cyG/pq5b8Q5gflUl6e
sHfHGDgWHyuKFc1+LpiK0cqQEIvIzbJ2omOWLXHA0nSWnGXRZ1sw6orwQPFidIG6
tuGDj5btuUPJRycu0HjOyJnqLIFwqjfMCRBX9f51G3sTMpM4ptHexDGD32s0wF6x
EEvyKVSccYhd+mVYH99AxPoQ6/jQujNYxuo2vh5OG2UIIjZna+fLbmMw3P8mU5L9
/jpRkeSMPnahXNVsbHGnfwdDmctGAXNCPQtPRyMjlB7cq+tvuUdHYa8jUUDaMy1k
fCwpgULhRhAaOGIBy/6xAP1o+dd4ckNH743nVxsesZBZ5jkVTI1DGknq8nh5W9r8
DGyDbWzEVrYnrv23bq3PHbREKq9w7oOMPmK7EU3XHoFErUx0nQ2g5VlqARex+iY3
5CzCn3LixZTwl6RghdCDfigIdDY5u8FEd07qJpznw43mYowmfNiQio/Of+kYIGR6
gKfR9he0osWL7Seydq14bT0McG5TYTiccWHLM6w1F8cY/U2oSopQOWoXpBEhDcFB
7jyNzvTEOxzfX+3lfdFKVp+/55hbe1456bD3zdjvxZcoEA9WuO50NJIKR2srr20C
JLGC5073IQupiJ7gXvgeQMw7A4F5xcDoaGc32cTtAXFw8UcVhm+IYS7nnCQrvimc
yB0qlqWpNpdsNgYM5v3FTUbWhl1vamW6m6XM7MHmBsO9xmeL4qtVmYv5SAS/rYF7
zs7FUgM7DnpueWfS/YiScruw0WQsDPCUiJNiKUMguz3LXUDMx8DXTgWU/H1S6Kv/
tny34n9C3clYA0l7zOCKBwYEqNy3vFsIzNjO0oxmhF+59DPeHI3k/8goPeXwhURs
dAYR8M8r4NR3rLup+IG+gN1DJg02qybO5wNFByWaWFjXapvl5iptB+r9jtEWJ8sy
xa7I9TJqAWSCf5R0yD9bsMH/RjDK7bxJwuyt5UhQjSo6hCwTgfoMqRKUyFGx2Rg2
Ey0NxAFUioSfaHXLFvk4eQDKlTanQcaZitGchIvEfTnayEM6f8p88XRCZP6+V/1N
unGIxrxNJlEjA12h4XfY24INmnuI3g7vn+BOWF9gRTxPWxrVq2On6w1RB3HU6SFd
JVkFfMZ8hr5YrPKoFtR27IW3VYCi+haLXZaJYpzpbx/5LSjc9JtXjThHSOOoyX97
+l4uJaMM7qau3zgZNlup3s5E82SoWPx6rS1qjUe/1v86MDJrc9jsVgqZTEw68qYH
kz1nZFvG27OjStERSjqxlnVlx5p83grpKQiP9dmeuGcTE5JWWN9h7ofUs3RvjQB9
mHt7hDnfuK7xYLLMEiNQew0XNUfHCwAgoFX8ZCGo8+ZKIUxQvP1e68Bg8uOU48cg
l2tvLJBVgmSH61LSlPtZ9bgfDpbiSEwYBzL3mxLbYQgBJwwcWQPM6xFW78L582QT
aiqUM3WfybU6Zzpz0iVbt1XUEQbt98CqoOsx3b2g1Y5y2poaM38T8r3U4BsfT7Oa
FNDW/Ds6fItR624ThjyiTo73D+3SBcfrzcr4bdbj63BwLPSflxDInnQ+Xjp++NT3
65zcOXY0AR6u5aZHa34IG/pdB2+1xhD7GrCgLMGFtI32Zml3E2k3cha2I8rRKi3X
OPW2ALCWdqhjVYuLWciYOC0ssM/ksLyhZi4IpV/hY6mCd63n5gFiq/1c/9MNZSRB
IUP88jNmFC8BYfa/F6yFk/Rz4Z+sotF0WO7+nWtP61oE09j078T87ZjaiooGoYPN
HvYdKVKPi1K14ae/6q/93wB6R6R2ywKMumpRz1UTuDawF+ix0001yGqM8EOraR6g
kONHHdesfmcXEDK3zu1XahyxBYqM6i0VL6yAH0M9XpuqMs/HHlDEBNX3kQnu9rDh
Euc5H9q02x3EtfZUMFPPFFB8G7PfIdZaL3ybSelORsmZ1x/yCITYgHnZl8Fv6XW0
8GEy7f4y9Rpw8W91LEoz2Qgl4MI+GFw98S5zrnC4wNj8sLv5t2uA5aD9Uh76rn+6
IJL15M9bq4/VrQ56o08eyIcKV3yyXSvJq4esaUxMHglarwsMuuNkiWbBIUcU3rR0
P6V+H/Td7GQjxYv8fOGrxqXsjnByyETYf86g6Vap4pCvFXwdJuTclQoQynkJJ/ih
aWe4+4j6j1WxupR9PNgQPiWQ6Ycj1+k8PnfcMnYfMKH9XT+9RrLJFm1t93U0zH8l
h9FN+9c9Qc22Zsm8O+R+NUWNKW6qYr0kHBO/ZCzsNW64Hq2sP1LNkMvW9MzNQvcN
yl15X9cVmZkl8X79hlXS5l7+MC5TRfd8dTDXvBT/o9M9AbAP3tWH+y3+p3t3mI0S
BWm67kW3QXlNEehKxRzA99HnOg68rueTVVDfOOOS/C2PF7P20ij8qkn39a6F7sK1
UPll7IDrChcZ76IY+eGSE5iLNZa/O4rMu/i8fGaeYpvtOFjUw9XKRO1DUw155u+C
BDUCxnUQxRYIlqNbc9Jw+sVpwsWHv9wd9YW+pVV+ococakQZasw6yceWiEeTEfMz
tm2Os6OoiPDokglbjTI1Mc5nuyjyGoIvTnw3J0R9ApN+GO53UT7NV3/o1fWsbZXz
KJMTS8GduWgfUTLcwHi98csDsqXySm0zE5AEfA6ESLO07FDFp1iYJwWqsFWnn27o
5VM/rwxcjRMw+FvYrdSN1FoHtjqxu/jlDPeZVFhTIHjhwC2kUjQgynJf/afib525
SKNdHv8ofEbo+YrFOyIxZy/Q2iw9M0TqLPzJszlABsbWXENDK2Mwx16UVPmaIFH8
4OSZZFV48Jnw7oCPlsztDzRPIoi3A/PT3gN9CyUE7mqe9OSUFT2/aFIhRA9pb1DE
U6gP8O45F+roBOAWAbNFd3iPApM902sPZp40YDRuvTqUCkxV6FHINx1pOBvwNVUp
LYWiq1bqYICsMHJOSCR0StxMqdyEHVhYkjYxEfbwJzNOwSQC3iX1MmWDTVA+J/Ad
X4hfvFmH72csw1yWQKemgxUEn2trAqMkShiOymdq4xNgomuShgCVJRNcGnWU8Ssz
hfZVMnu5V+F404+npQo1wSxia/+lqHhT1usArRjW2cNi38YLNgpYE6qgBrncCusD
G556qT37CGx2Kj2vfB5ItuhC4yQ8+RmMCO0ZknR+lpD4vwlEH1acHAXSzJvgBJuA
afC5bSScUw/W906juxtl5R9JbQfIIelPqrGGAgYgVCaN9Q6mPPeIh42qJYNfcnM0
W6AVwVMYw12VUFm7FTLZSrH3tAdk20Ov15yOdy4bARgxP9+4AQtXgSq0FqPo4HIg
WfN60zWcFc/8Wccf3KGaYgXahpYdb52kgm6w6gQLDi43jzsV5QTgJboVDu9dBPL3
fOhfrwvEHN5A+Uf8x2sGlFHstXz8YqgvC/B6vKLwc1lIO0DKBzHbS1nKDJIqF/Dk
+Grvhs8uwhAv7f0mOJJc+AU5Qa+bXmNTimyf8rWUq9995J+O0u+HBUFpMtm9yA08
+HUGSMSSrmJH+wjU0H8Mly4Z61x5vsGjS2D6Nbj2/KM5HDFfwpIhgB4EcjtoeqpC
gJgFisLVTnQB+RTfuPXkpXmc0ciOAa6zl2LkceywOVOACjki1HUehXK3kD4oHPEe
rsV7rMZUxlV4yp8b1Ptsqikcxu+2RSx34Rttx+gF2YXWXIx3jEPgkMgLq4H2KYTr
IlRzzGFDUqydfm+2xMTytlGtw6giPEUT1DwGRoMgmNY9o0k4wAG2tbxeZHcfAozz
tEjBfPhFDanZtgiT3/gV6wal7/I0WmVmyPuF21LvyggyU5RTmcBl7PZj9SFOi5Q6
GuKGgtT29yrXK6bQIx1ZzcCG3i3dzIC/ouAIzoKhsBZKRxVDJDgSf5XQKZLrUQ8v
m6GM2ZJDlr8fB0IBm/SthaT2+C0ijBmwY+5lDrFbJvEx+Px3LKeZ36bS+8VhRcY/
928W2vqLAIp1T1QABtQPOUZrpTqZmxvdOWYxZ9C1GAa4WqWhf8k3bE9JjbCxxG5A
ORLtkNP4GgLX3LQeyO3vWT4gzL0qyFEI6r31m1MKxTKK5QWUbJ9pvqHaHFdwxYPB
9hcXigg1VBFUJ2+r0bRqvTC4ATimrXLGSVYqiHSmFCF2eog0ENw7jemEKRhd1aay
/JXcLGQQkBuUSB48eYU/uFClUlzTAfoH3jCRLfsnzQCar85vqOlCcNy7ndswojon
x+Z4aBasLFaHJl2cGw58JwgNxszqtpjriLw5jW6hcEn8YL4p7F0Rc2oFzntiy55c
qv+Sce0R0Ik58vZwv2wIAKj1ISVfi/YvvaUOhQ8zSdLw28JNXOZzutJwrWrixErf
0S1gHQE8rq3WGtTXyQCD+ku4C6aTiotamFH/VogF+2rowTSVBir2wIDIxgmtEpRq
FfjPie8TmWTFB6LEJ9dQlOJvhUUXZ/4qsgYfU2Y1sHN+r8C3epayHU2VJKi/8dL7
piOPCFoDxpBm8chFlKnH6WsuAdVqANwh4IlfSGecZlOb6xdeAhnK6kKKXZSLyLPp
rknyvGIEan5bKHABu1gDN3LwyTSHs9kCQb3UrxxTzi068wB73STN0IkiJGRVsI/o
Lw+2LRHCI4pgP71gfNt8xJuUpdzfOi4To+UiRffVZ8tqbtDOz/8OdTx8KppiLwMc
e6CyMA9BrzJz1AdIx8cv34wP6CxmtqGSDDCZ2Qxp1CafwkxFoaH+CrATUMWs6Cy5
v1ymay3pxbnMJ+5Cihy9eRRUiUNtzjIreAqvnNqEiI/W1uxnUlKfoDlTYdlrlrVt
WmmhKcyHYb+JGe+nbbKtO4vy0GgM5EjJZxdqDCLY0SJAk41xSIb3eLXZtIbomEZd
c/zpsG/Kcazc2zSw8vc+KBNE27VbX/nptBmMX+1odaAe2l/dGVa68tu7zc09BFsA
U9nKx/v/wSq60QOa4ehiL4QC0Vbzz7vwowIB6tGbpaeqbL4uYfC+6mA0ow7CP9u6
+zS8ldK32nmL06b7n+FSjSExlJdVMFhzra8oqrAGtCVByUiEU8o/iCP2ul1c2+eo
4UaJZgWls8llCblioynEpN2ZFnWmzK2NRfXfA9JdrlCqCFBhutOzES6Zgnk4Q+z9
bZHk9gtx4MyCzXsUGNuymTzgArxlYNSa2JYb4TnBq42nlqbLIyEC4YyTZNACIIBF
m879UsxydhzHMVn3qQYXJsB9W1wVZo4DMftkZMxaF686IBrmOTa0pFPZ8rKnic+U
srxqfvoUaR/gQUykwRbtIw7Kc7Fh8MobQ6N2VQDExm5LL82OCjYg/ieYdWo2+JZR
rZ30nLPXZJf6aWURigWWWZc3Bv0P/3d7Zq/zXvRgm1VCI8D9gzDTPw1wFZw9jriv
KnbmqQFRcDh5DEasyu5kjTVFIb2KEGCh8GcVvF8VDuzc9UUUdnQdP5LN5WIKl5Fa
arpxCmbjKl7zxy3ls0qqjzadCSVigkQiu0YHstM6ojZfPPeHUwVoMXkHGQ3hiFza
wzDcHNxRi4JznTCZPIsAG/AMo441kP5AoLBjuCPpApiRT5oX9oid3MvYwfkzf/h2
2r10eCliAkyg0+5BgaClVmf2fSEPnNM/VS9hr8otD12biMwPwST0qhtp/Eg2F5O1
RmV+FkPKNyxRquQ+N1SONuE0KsEikHIzLB/FfDoDAF43dKbnK2YgGIecNCZiwgYH
qLM9jMyIuX8yK59OIkLJaDbxmz9jre4FvQvZMSRdJ+V3BSkuG5srQoMjaatpIUek
O9bKNuNreT/YJwlT+6w1tSCSTTiuRvNAaNxNb0IDcU+FLtnH0/klnoH6chATVjPg
Worwg1cq6+OnFm4sjSnFb5/YRib0GXzJBX8xhS6JCN22mnxBNr/oAJqWtV8sRJ5B
xJaTEzuGVmE7W2iHbdwQmSQdth0cfM2thb9CkFPJ/UkEvJuFriVTQu6lBQnisXMh
mAIDnN0XhX+3oUil03de2vDJfBjN2sLQXXWwkD4E6QsGHYQIbGJYCK9J8jKo7wEe
6DMb0JQ8VgMjcBilUEMXkiZC2nDErK3KrJ2aAywTmvEqqLBzPAJVGdVqedTi1A8+
YmduVPxNRGQfG78646Dkw4/1/a5JObGbG+Trlg4NgJ5ShlLImPd5qvsoFqL7wR2E
NJNFPONmcodHaSvPT9ZJoH/w47DwV6XjyN2TIrbT0UIQAvwRM1XZgVUmCcMJtLdg
NYoJDd8sW/jaZndHRTXLAgqx4hBozSRVCr150g72v+pmCJUdb3TGNkQ1tMa6Lozh
WniKuhNpbUITRofXpvnLJtfTT3N8GgJcEOq7Qlm8tj41GC2LCt8Q6co1FQy2qXhN
ASChWGdQTmgdOx8WE+Vo9WTshNEXbCHJEPWBiJJdLoy9QZspIknfUZ7r+9r+COeW
C8zSIqkiQSQxJ5gaWMv3nPKxAkZfynbGCD+J99iu0NrkvFR4leH2VpOwmF4GtUS0
YNSOq9P1YcimfWpm4sma8aBiWd5u1rxiatQWSvuOi6IJWzClZLpl6BbUwXfYOsVR
CNtxdfYzQk9TMITuNd6CalISebeP5kDKd8/Ml2wBi/hFn4GE6Zo+qsRKv9CvsbHE
K7ar6rr6KmlDS/Mx9O0FqDb4HpdIQHGIdYDRCWNwA8s412FSyZgMWSesVtwC0kl3
oP6XGCLgj+0IlUE7KBZyNWW2E9AqSBfFm7orlwiigTXErXO062R5cTLdR7RERMiw
EfDtLiOXVWOlRStdn+PPtShzBj4OHIxcDXjtcEdhpm4eJfkX+gnrcGzOR0hyEccr
4rAwCIKtP7wdRr4mINHvngHJwhyW84qr3MZRea+3JuQZWG4LzPX3BsGMZ5tk34O+
zKmfqYQKFgTx77o9KC3GSgty0Zh/wdkDi8b/h0wXlSpy/Y8SR7H0yg/fkF9z8jkA
9gc4SHXcElhmT2jKX7ywfiy848DQawv70k2pXh+QgrV+EEsSQUVDk+jBDiMvZLxv
vUgYJ+v7Yz+iU3k1LT1uqlscsmO40Cr9uv+nJRxfnLqTMwFT30LJoF1S7nKn7Tb1
ipcwz1v21kbIext/CBZfhU+4HQgerAgbicHta+fmP24JjdmVpFywYCqaBJo17DAZ
ZXxClSkt35jQwj2Yq54zLelVBJRz0OCdPBjBU4AfMyvbx1Y1Grs/56Q6QPS0ELTy
YqfAN1kf+LK7/xw6mCg3dj5GpdntCloJjUzSheOvHcO2eq5K2TGRM6VgPZCX4/Ol
VMu6GeawlmA7gp0UK4up5EARFDB15jKawx3P58I1/ECgx2zX0xcBX3z/epbByBi7
hwuwnZY+m21DfCNh4sgEJu/cvfSmMkgWBHmpZ0mS+70qxI5dEa+mw2InyWB/w/Ac
HqhF9xHpnlbQQULsktN78IkxGrZ/8iQvzjUmdSnrPx9BkHIJBeMlQbPvQoigxSW4
3J9FQ97cVdLTZ4jW772/XpDeDOy173aN2zg/nQRjsTjmQU+g68JhcoIxL4olgns9
o1sGrNzqpQZ9Ti1RJm7Y6Dui1zHbgB6VwzQVHNMwWfqCPCc+KqftyT2fXRCfws55
h8rhZ3Mqdxyvi7FN76/WpR0SNWexEik2lrGp6t3fJmL4JNWRj6XBBH7ukrgGF12N
H4riXipm4cvi4MHw3ZTARRcjktHYZJ+s1HlqgxrKHUPsPhT/zFWwcDX5XH334oQr
DRyEn7imT45s6/IIShiiHGFe2gvJVmykz5pZv6xMass98bKXvEF//uWt/lvsJgn+
wKgZtDmf2cjkED7wiQFFRfFyj3a2gHAMp6riSZrufeixpZNx6V0YSdJap0G4mF0F
31hoce8wa228bNQxJmqIAAJC3P/taw5G2X0f2lpERPSax9X/1xsKg/LWJXmefg7Z
SS870lNQgn56eKhcofMICSyLRjzk96gYlwnEfLpOZ2blF1iqC3dHgviSBz1y+ZwQ
ZcRmONtRpKcYw6mPwQeapZ7SreNnyBtXGyBi8h6+MC62G2EhvF/pTCUMH7XUVQm+
dTTBulThnRMORM2zdc+7cIkC74Zi8BATHdSA6MQ99vAE1Us2IyOy9sekl6gMrPwZ
27qZzVxEcBuV/2kZw5229zGceiNTTNxcbqIEQL8D/XpPPCCpinTWf7Bz8MrmWaQN
/unERhHBkfEUSfOpToKm2RVdouEWaerFsZX65nhCiqlSlzywtvWyGv2r6ja4maoL
LY3ko5qcxxEXUJhzhH7s8Ak+TyqIXHsuZF8GfSbbaYffGlYZU8SFXmkyuUg+8Idu
MagBNXe3sqEmom/qWql4Z6saNH69ctOathAG8SLojSWWxg6/i7EohcPpdhlfb0jM
2zRb4lfrhbztVgqP6E9sw67Q4rIhKVUZtPwo1x3yr+v7TkiHPkpKZmFjxW+pHzE6
MVrH8XHro9t3R37UpLlIOSKdqL379aSkQeGHfZLX3a0GZtidZpdNgFDEpgv+qfFS
MikbWNZQzE0QFJs0Ivps8CmSA9C/NrRLfqx5xeExjwmEhpcFkhnF7tduxIh29+K1
dKK7fDKHr72vKfvCcY7nzGkeanPD9Xc69JySjCsElcHhMR9slZe+tZTjaGEXF5im
Ch2ruQwBXgPR01tNWc7EiMiKpzuXwDQMZ6eJUFsgiEpreaRZfLtwvyaMKDALRDsC
9fnlto1hU51iQuGysTLStp5qBF9wVAwKQO2bnp8RBf5df3BCOWIBEVPt6cEIcWRA
YfSSg3Ar32y20MsjPzikAKiEhci0tRECGVezSkjQTLWQWx2hZadxC40aLEuyFS68
9g4uniFpwg3A9Hg2FQOzZcNcEHvH4RfIQSPS8T6E0akT7kFsiJIivNNxN1pLJ64h
3kIxdYKI23WHVYi75TnbrnKcY7rYKucxDqJfw/R04DlzR5aElMcgnNPDF7cpI8+A
nQme1WlhvuIP7CQKK3bYL9figwWSwCq3wLuffp8/2yGFq6I4+9pKAQHGGVOH0DJ9
6X5tZR5Niw39iFS8s7scCZWqSaXz0lP9fXEQJmbs7XtI06JFI1lGNcmFKCElUBVT
I+Og5uJovLYnTW75Mc9gtisWv3CsM90Mfh25KxOZj5F7z+iG7w09kJDCASUOT9S/
8GhvdB2Eo6rk43caao6y7J9dcRWPHiRSB4cEFXACpF3Lpt9MU/v1yqjlV1MtEhZn
v3yS45NhkRcXTXFlvq8aUmyEpoGRKvy5hQBZl7atekilkws7qK8Kp+v+ntIk3t6l
i0t7/pa1gFtICZk286udBF6oHw/m2nP/fMjdRCchCHGNveEhKn8YiqM/VmTeDIPc
gBa/njkvOawKHlehPazjPEsM6wZPbbbmohTMCucaoW0pqubcYoAEa693g1T4FZ4E
R9A9eXiCWsVBhdqq96O2MjMbekVlyu867qDXMAJ1Tle8PiIMlqwWut84LpefUs6p
4Le8Rw9oDHDC1SowHTiJNxsYCBGbexIMZE674iIlFAJUo7mywiUNBuJ4x4Wc+mly
d8+HM/XhzldCmw4Wk9fGMfK/5Oe/qRdy14Dsqqtoor6S+sIK+Q/GyVaNnzcZm0X5
PulsFoBbda4Zlf0DjG+0kshzQXN3xphEmYPpaFHuEOuH/Vo+cpeIzyZXIjdfzIAF
ADEYm+owkCXndc1/4pr4cAPY3yxLa3JRWgqtmRpibza8tpktYrN0q3o2/MGqscdJ
YHtg9PROaKKS3LD1g49vY2y6g1IjyuolZQTwWRDPYm+k3gzl0gIjOzqJYas644cP
glJB7IQs9xW43b+YZjS8MNtHzhqyuzBIpkPvbYxCL80G94lqr6EmHpnVUonG3Rba
jBKE2/ejfd2OMhN+Rf8d0VmZNM1A8IMVlzqIEK83gIUFpz4feIsJEOH96akzn+Hn
+U43aO5VJKyMbad6J6CwySqm30QCTbbookXzTSwOcHFU887IT/biTZ+EJbnarvda
7kolQ9DiJtH1OT37peZblGOsRL6Da7Y1ptawNnhickYSTEP3iSkmxP53cG+AYiFP
286oXyi28zUBOs5IIR+brtHc0LRAY6UTLcfJ5UnK8f4CskXQadOZkiKpQ6lZZS0c
dB7nhgxjfiHYFYWE2FmZFjVihRi6It24TY7BsELAiB9G8GbdxAFPWU+ZRJEHb7Nx
D1m3yV0Jn+RwhStMcTILKZwXmuo91TM+r/g8I6vliO56o/muLe7GQXNMUorbq379
IiCtnYl0Gngo3lb7cvkVxaVrHEx7lSpL27evth8JFdjF1SFN3tfTHq8m9TAoyqmn
9SCywPfIFMlWzYEV6766bx5vlGy16+Oqjs+JqnGIowGXae+egtBjoLHSOC2fT4MP
xg/eq+PbMwXPhBfXDU5+9LIkTg2Gi0nFLxv/Ndoc5p9OILvPDkT1+0TkxiBTgkQ4
Jkx5I/W6V7KNJVmY658PCeZZwI/NSW4Siyy2xwYm7zweDF9Y0HHGjrP4QoBYMgtf
kylVA0negUHWuqEsaLmUVwfAGwdGFSvQAFEDvQSOJVuIDCoorczESetf04ivbkwD
FqiPVG7Sywqjr8olQCB4Bt/8CfyNShxv+yUsRwCo2L36iO2gZm2aK2BVyPvcHHCr
JvRDDGaaxVpYkOCMynhEJc0UkJ24ARsYT+aFCLSJTeHIDnfrGcTYh7bWn3p55d7T
MKMGbtZc5lWIkaN+mimpflZXIWGrmURYKU44KB9pbregBKXEN6e5USDK6Sv2dnxf
emH7j6Yq8tii6uKoCxFkbEja1ZQ6cj6RtKNHEmUZwX9gI+iOdNNDTUR6ky3metX7
PqIeJp6KYybYnu8Pn1E4efLk6dy2Oee2MlxXv8vALOMLKgczPJNP1o27zAnilZTg
mK4S+mxKPB/RB2HdbStEsBUiuccGQnJWOY7cFWAUtB0woz7llO3xiE881LsV1Dut
F1/CT1LX/yeW+ZkEJS9LUted8pQ7TZ+U+hyksL6qxckmLC0y2jIWPPM9BizCOx5W
PS/Pf5vvuyXcD1CHu+8IFpy6ou++4i5lYILBsjKjf2HwcIBrJkz1+TwPYqKTdHwe
LJz5844D1kgX93l+JjmJvayjc+4hi2/1dBa9u5KHOPkGPKKStDevIg/Cijc/D/KY
U5mx3K7OA2CQdpj5zyTH+JP2q2e1GQ/ZokQzNEcTn3xXCiIl+huipI5cANVJ9JpR
zY1E+Of0SH45wpdITwWwm5fld0FdndfC8Dr6Kbm50iMk3814sY8fQzZukmNByOEf
z00fXHjN+xi59Hcfegeekh8TOeQucOV4ORTipm2iHvdU6zXn7vQXia0hruO5frpU
eoWlxsO+BHt1pbNQjqQeoup1xY50QXgkYMnecQaxOIbJUghcdA6ktADkoaP9oruO
31utCF7Z8zxxfm3BKUXHTUDjZkIDU9+5gp+X1sZ6UR2UV6R3WqdPrYUjXr2mXToE
tUs7F275cBbHKw0SQphTRQjmAzarzFqbnfu9ighTjucfl4DECDl0gSkYj2T0pE+k
fgvdIxrfFWwFYAyAR/o/o3aEIOaGxEqVBJ4z599O+tDn5igsWsMUikaxze7PboZx
6RD/yZxFs/R4VtY3KszDzvFNWUVsJOHkrk7khQEjVs4uX95L/YQovfFSkq6gk2U5
VE6VCeYpT83WDx50tWjZ4x3gwa/qm7qybxJRLX78VE+V2a1Iu+3TvWtwG8dTeFDp
Hna74StTN8RBdo6hNjW2Zun5K/uE6wQhcgWElP3QlTb3VVINbWlMm6CnDKCO+af4
3iyB3icZsBOVDF29Vo+zBCLTqurd8ANi+Kl0UAF5Vb67cBYPH86Z/0wdxwY7IYpE
XXqk5qXxF+MYh2AKnlu0ugjOxc1jJ5fRwg8gNX3rCbaJWFvgS9aGSi7bA0ho0tvM
Cy8rYOVAsjLkhl0NdyNUuajU3qqP2E+Xir/SDu/KGgSwYhaGsVZMVq5DN+CuNIU+
Ro1wpN0tr5rlcdyB/DMjkOd0uyWIuLU7bAhNxXwXBMKrTBJLSmKugfOCEShh/jqq
pWeM122r3Mw6QOY6s3RejkxZrVQMo6J0KhJfQNZFFe4MKoNCDD5tPYSv7sAJHFsx
f40H9/RmrFtLFfuUkn85+mE5dCeWcNx5tuZ0CtTcvOIbc5/aGGNgPBhiaBaeUuXn
8vqFdqxKgXP2JdKr3tNTFvpBcx6Iha7+QSFxvtoFDuwfS6g3f2Kd+a1xplJO5cKI
7+z8LMK06U9lGGdDWUUSCbHuUui1ueQcf5Q3TG+oG53i/6CKy7y41ILSBhqc4Jd5
dTgd6W+9tPoLj8AFuTFMQUst1aotKBhmOgp6AhlWdUhFkX49i6t91zW0lYsxDnnK
hnIQCn+LEshUafLRVK1B+/iO/jB4IDfOHAkY3RQZTB41Ht7jdbVIY++v8NrSm8Ov
NM0eR6WzEKhevwzVzPuqiHkwikIM8A8Loi0/6cN3p/GeiJIjWgj1BjMYC+md9n/H
i7K8IDslohC9r36fcbJZ7VFpZylJ4zyrC00Y47s64Hqku75jcBwn96z36AqMVkZk
rqaEWwA/wTMtxofl7cADE6BDfaZgBhNRy6Ff7Hb7pyO4cDwwoW08CdE+VWHITjUE
jsu658GKolI0sOM4Qnwebsv3U/A6E0P8GcjMAhNRdXQU38a+fvrIltdkc5Hk1nHU
IGY4zILJKq6+u+htZCOEGSkNDsjNlk7J4tfEcd36hfuS7UeEjQSu71MGy869Lkwf
h5UtK++xo7B3MAQrS+wUdXn/rE7IF4Bv5D7xwtXEVsHmw72RYsRPt/F+NtVzwrz8
/TiR2Mt0ev343viei63z4AjAvrVwuml57P0gHo99BAeAno/Tbsaca5keBSXeHOhH
g44k//qkVBR2cTdFZx2mDWlGYLWmCi0ZKApv1Xn4gt7NwhxWwkt71hNBzbgL1tR/
bpmLiYAcbM3sXcc5HBsGXcZSCn9280QicnP5/65/U7AZdf3tcVZcQEScoh7Yktzv
t4y81LmVuTLX7oQdUTTvw6Y1jA8cH6ho80oNbK8OwcfrftVk8pUMAotSg/tqq063
tEUwJ9qwOSJ88U/HmzlRWqglLwg2nsZHZFA3S7nJEWk+zXSIPS26IvWL99gBgtiH
nVq4L2APDWcnv+V7BXmMcPC3Moa3fezB5DjhRSKKLZBcACkid0SQhgy9qU0/TODv
8u81CUBxiasALdCqU9Gp62PHekXbszURZ3ZWLa9i8AzM5QA/xRk6SZPi99xGXmVJ
1gTO7EKBcYlB3eeCEnCLfn3mF44A40knulwyb76z4ACxaQUb4sLsW5Ki46RFSH59
iHZomQ9HLmsP1n9stxYFbVxqktAfiOHkxxnqSPEi0lYBzhwZxs/RQdrECwAm6OJc
2mKkYZjxbzNFb7DqEtPXKtDbQkQmlysU4PN8BaCylesynmY3Z+aDdRvswB0QYSoC
XNNjSHd40prN46k7hzYMN8N+JMwnd2ou/Ouz2mg1FWn2oms8sH4BusYdEFcezz/6
M1NWptBUKhhGLIRbB5lye73tcKnH4c6t+9JlHqT7exw6uIk+w/g64RvMOu/dcJVr
EzV2N0BdaVEHo5IcFTqy+cu/90xjzKLz7QYBljIYK4RNlD2Quxvyq9PMhd8VJmEr
FnPezhPD60Z27WUqRwt1KvwcqNeEYjusMJpPWiIWiMlKdBtbBvEFhzejJ+fdpbeD
2SEUN+n+x7pHgBYTY9hpJsjwbNxmWn24rKsXVQzQfAOFhgupVUHutQNdSa4uloYk
w2GS8d40fsbNeE84BDKRb4kaYel2f5qcF4xwUPnVr/yV52X3AtC2kZ4Px1qUfXAi
5OPMAuJG+Zyqv+pipG+iOi3d9PAKGx5cUKMUAb+UnUaNxizqJtAmfPpl4rAY1SZm
cAdtChhtPzpyCTxcMkM8UvViUMWKXlHTNoN3mkiS5Gp9ncrXKu93cfOdVh6rkLmt
pWNTuRGvcY5hMItTS2DOIga8GZMYxYncyqCYmlURRpJWZkqXr3JlGi+6efcbKU/c
LeiLKle65zlsIkiGy+2u3FZUOn+t0QVHoa4DBMzRVYv6K2vCOzNfrwHbhNDk4tgj
EAb4SfwQfR66vLZBeGgx54rkXoHj5fXX6WTRGFcLmbRDIQ+T+QPJaHQ65soTWLw8
FSoIgSs6LMC8/LyE66C19WtEImdkIWFuLYDHEJ6veysBrV+qQNzjJxqXelc7qXOT
ypxAGXpJDYnCihTij2OA0kPBkIgo9XWbaNezGsNqfRNQ5POcjiIvx51+m0S0mH1z
D1pg5KP0+ClTChZnABS4fK1vqL/peEsjOsoHIVGpGKzAQUOPUnp1OZE/cMgQLbAt
hz0PqbBIweETt3ngyflSiGK1sDE+vTq+0tgHv1kjkp9CyDonpcvugAx9M7h0rho6
qlo7I8FkKP4DJ9H+A/pF0/CXvm1shRyKXD3JDBEVsP/nRPXyompzA7YlkkdvlKmp
GSnMLoig3DT9AX5JLX7FA5YmUhhZUQiJaWVXU1w/onNQOlAmlTFyhofayohc/+kQ
olf1v6ZBTLPw0uwy5gBJVc+JsTUTZ2I1hxGUwS6bNiKCmFXEtL6M73IA6kQSjz22
omPPqzxjSZK1DXZwU6ZSvQK0ZhD1rtmRxp20UlJMctzEhEWyyeB0SxFZ+XZ/6iej
xh8tEAaES43HfdVkWLpHQbjSzm/1Q/iVLCSQGEWtPkiFHUSaGgInxG8Kqyr4M7o3
eIPIMxNWXuTx7AynBgbypDkgS81EbSEwghsu/c05mYksV61V59X0zwKS7RwGkWQz
IVDpAd4nMYOVRMEp74QhpTGI0DjXRuk+O63aeUwY3LbzH28cuEX+sGpduWNfm1sX
0IJc3a+5t1qllQ8PLXw3tf0smU9EVeoBhBYSs4NEfmw80itUH2IGqUA0uQWi/Xeo
MmLXRweyaq5bpjjnOvi3V4xHyqnH7i/aFs1HxkeWcKUeYO8btD852QvYBTWCJWjp
GaiCcpyMd7JL6XQ24FyzF6kwznkUl82LsZ0vTrJskBCEZNyYZ1IcgGfBLVPhTXh9
bBw58sa/xMzAwPT+4rm0c1R/50x1M/eyBcYbVWwHVSBey26gTayEUHFz2rz4kqY2
2POND/98KQeJ6w1NORoIImt3YkGd4sDbWp+iz4BO/VHBAEfIOGraW+84JIWLM58o
3fSBkJvY9QQt57IR7G0i2iPjk+q4lZcsO5eXq2sWfH5cCv7qCb0z2mXecQfrg0FE
Dlu1FoBcaSgL0FW0cGnwwwTRNjVe1QTG9vLk2lEORKzwnTZ7Ts9zKjDG9Kz+aNEI
IFieUi31sRVydQn17MV1oWhq9BHmZgKZ8FSVRFmuiGToSO+U86ZDAxNXAobOSSf4
df1kMAYdlwSw6NAMzBO4Q8Myr3vkFsVrfYpDMk1JpziSReishMtDoJ3Mq+Rb4bOg
QjO9n/v8ktC45gKY2lTCdC8abgz1c4Fyx+lx3qw0Gpo+5v2ItJ9tEQPQfFVbdQs6
AaDLzk1A814dMHLU0wP5HXieCR5b04hSnWFMWdZ9WWnxoQY7HxrDnfFcZ3cDyc1W
9vAZ9WcVqkH/JEzt6pxTyj4CpOJqFgrbcuQngI3jzd12ShaSiMvPauY35ItIV77H
cQrJcXKRz879xCj6wgxK7Xf2ItgLOBeFQ4IBUecgpQvuCG279ubmDyz5oUcRmrUC
/hAwG8uPVJhtQyCLBE/20WdYLVpOH8Ijmcl/lwAKJ9VHVmsvIvrhSu4CxzepGObG
iHVXHF22cKYJf/dKF89FKlh4sqa6qjinNjaNUfrGbesuf3ar64n+1W9VKI3FBAyS
LvkgdpkdYhajkp7kFN44uFnPJ4MjMlMLz9PTbMMwDKQ8Hbb7Z0jMJsCBUPM9VHKO
ayrhBRRDE9pnTJjYfxVVo8LSlRfWX3c5qoieZqDA0TMDzn/3vxMOZJSi2Gv0414M
IT8DdHLwnADZ53lYeeTXae/JWXl91hlnJb9i2KBQkCFoG0pQ9VmAWdbT0wRmJkGH
G5ZRcV/g48K/rYpxG/UmMRtcza+MaW1spfe422bbKL22juRgxxI83b317j5IlBsX
1wriwGszOLAc0DkdwuwD/h8GV1dDD9EpnoKKRP8PjJfWSrpbVBFUO0qGLv+L3gia
WYnQMimPhpk0sqXip1Bi8g9oimY0/Y68vUPxZ2Qxk+m/zGGRGM3/zkDO0MPbQfru
iNcJD3/doz4Kg9lzrPCzsgGobBgIbed7edTenviO04PtPd40BGYnRbG8/XU2EsDp
EOuCNchKOUjb4KWWPRaUCI3VMo5D5HJyp2MvFPZwUibd4FngR/YHWpkb3lBmpodr
pT8oTtwYHIai0Pydvs/zEvm0FTqvq64/TeE9dDk8lOgdUfIxg3p+4tiw8e9DcdYf
XWEJ8dRi2Y/CNnGGNfxj0ztch9Zu/AfmELkBw8rfDV2TSkz6WhBVOinitQLVQMO6
t/D0ScAntwbk8xsbSzn1qONN082dk8VJY3+9GpILXphbDQj0qVWTnlfRbgCyA+Pj
esniBmvBAZ3hjs/bSTpLM6pSeYDCd6757WHNMacEpRWAGkptxCLpDKwQElTJLIGU
FkfHsjbn5Wj+MA4sahn0U2fexQx37WIxSygFLRroun2s7DUlyRYYQsG1FP8YpJXZ
3VdObUMAw1cjii7S2JXClUsm3AjxjNXOB5DbvHSRJOyPhTwkDQK15wU+mQTSBG36
igRwVG7yopGnZ5LudAXPZbG1Q9oT600nfkbo7J0n0jfwsErJsSNy72bdzV1AEBf4
n7FdWbXS8GuOWOAUtdVTEQIkfgRhtwB6iUx3zgivwY6+TrrLT1qO7kyJ/Q6+xax+
Pcf6ajg8iWWYPDqd5kV9M0H/eUT7jC5lUwy36bsxYdcl/HpBc9pzsjk/INpqL7OD
RFd5Ll1vjTcFiQrrmW8dh9vvvA7b7ZzmetMsHwHXCOTL0/I0IwSsMHbxvS8uMnGB
Q6qqThlgj1+cLlZDXjVkpquDYMPf0WW/MFstUxf6GXGBmDC1GBlzI7mHaiUTbY2/
aB6SQ6A8ZVojvpEUsOhV6e5izDF+Sf+3gIAcOaFAp5G9VW32JRtaRtD0e470qH0/
IDK15rEP2IfEuH00AbmQ0Y0NTnuFlBzmXX0wS+aT5LK/s4yBl3FHyD6hchChbLWo
xTed63/9dczHokdlKM0jaefqlS62YKKs4iU3njVOc8rRNAD32PR3Kya8o1EL5LuS
UZzHqDl6ZaD3Qu9MWpCPFRJjNEeBnNMtcGyDe2lBngnE7yvclaTjX2DA/1VjxNk7
2H2ozO9v1drtPvynmytXpd6VZzXa/m1bEDRWVget78QHtXoSVTEi81/VMn05nnag
HopJXRQ4FOV/Jtj0c7K4kJdVRKXo72VmtY35FrUY6ObOatd0MtUbU0NjDR4CpCEA
BlcRoIEhfKDeLDzDKXF7Pq3yGm+KrnDMM17tEbRut71QHHhcFAd0khgPybreNw3X
xT8WTQltKL9oydJwwY/mfYrQln7OSP8CMWaMSxz3ba2CMOb0GhVYilzeKDB7aofy
WuD0sbPYBkRyLOGzj7r2FT05NkwAfgSuHyORH72cTs6zsQXq3nC02aVCNOlTYd32
YLZlLKa50RCXlA8EXUELN5w1aQhuITvcfbA8UQg8WsQkZvW3qVINTsILEG9/Z2qu
hCT6oB/oVoGPYQN0pOc9c95C5FBFUNwRU03IbT/6NC0p++teQFFkVk3bxwDxTscZ
3ldoViRfOpjz/Rt3cWjkIcMJxpaRgBD1lj1LH5u7DqddqbkClAZIKloSbNo++Wls
JYp72HW0Jn8ar7DnI9RxjUOl0TaM6XK2Wp5phZ7FxRLD+yGtWeBQ82Bb59Gdgefq
aEihJFGZUzQE15LbfFZ3hLt587Q54qFJ1Z2Ym58nzjOWAOH5RM4A/PXOfGesAS2c
TPZoH2iPgWnMRX0mvsXPidFUNrTOiVui9uZYb9H8N42ylC0fxBw0FKWYcaSvMR+i
0QAKX3k2fuOjn4zp5GVFTw2i5/46IuU2t0NOpKDOw9UCytAwUNKF/T3qscebK5KL
8KExhSOvUadZcJpPlwoRy9M+IOkt5lAtBS8ADP6dw7B5oyu3wktOfEYm0+XbpLfC
1YUfEScMVESukFslwGCiBs1WZZpMW7ZTIgLWfmUdkx0tK+c0q/Aro6ZM0K2RT/US
MaR81CMcGUzuaIOYLwTKrWi68R7kkdFEG8TMQJW2CVvedLSl3eRrKU3USyEQuK+r
mi/+pF3WKO8KDMaEz8ziG24TvjqyjKwoznAgEjZX3IJAJPwlwlpE9F9DJ6piBCDG
6vMPHJLPWEP+YKYVGQcTmCWmf0Rw1I/ODOlLqLbhfb3PxqbS0lSDZTAqe1unj564
fzNO1XdqzVSgbOW9KhLd/U9aeZoVWr+KAOseFl/3RV51sRB4OsznioC/g5v/LrLF
T01oexFfCNxIN3wUl7Bmw3dQ4g3Emv0U2uOpn1C0QCVvwi8pT6oZcPsLLqbpaI8D
/x47Lt6M6YyDwgcXlOJL2gVQKzL1FvIOSxXrnAAqbouMXnlQ/dLpU0Fr2slbO5pb
h7A7FX6BsXylsnjUZLHQdh+sEw4bg9vdEjD/bo52qCWgkUGNB838+cr4fXpTj0eS
r8oweSO5dCxH/g+zTfSdXko9wDu+y/ppV5GTSAEGxg74KpZ3C4SVI/x7fE5KmlUV
vL36QK0hjyxoGQD9N83jQy79KA/uJrTK/LBeY555vXDR3zUyD/IIe+y/hEp/QpYE
RxjQpGQ3awzg2N/BMIja/+jkcldeZiC+qgLRMik6Is+W4pN2typ5gwq74rVyOCNq
ytcvlyR3KI07Af1UP+qSkPxcIaE0TylDd7eNG/nwB2iKW+5lf3v1TFDwZIu33/EQ
h6uSLCd9Tyu6epMMHbgsWh3NAbsQg9WqqXexUaUh0ZHOU5m7gKdphTr934z+GfoP
APM521cfCTxFddNNPf31ffjwuh0NNvYdrCm1WWXUasQr/rqc+uPBswWDx0ZjBLAd
NKYcYp0C81A9a7uo7kwLanNRVlCv8V3nRDWrVXSCFfqkDGBFZc5U0MZU1zmn+KXw
U0wynWbDYZGDPSks8aZPmza16Q46YPs0jLEMjUqFlcXI47jzSFj4O04bD/P83dhF
+GB5Ebzj+bymKuRwKPyFttJMvrlz//N0/2V8i6alJTD9kTD/bceGxv7MHZhfziGP
o2eDS/9jrd4QtT59wsrc/c4eODP3nM/F14W2S6wtb2awmaSuL27lmid4OrIkTZAP
+zVB8Ro5AER6vqAfMhnZdkeFSTGny8nDuBMpmerwltYVzIu9iNvHTiGHj1aAw99n
ortgzYa53HvryTpbJt1FJwSHG9y1c90H03549yWRMMRzb2fTYrD6H5b2Pz6ULF5R
G3I2SqXGF3Alp2747HjRol7EqjRwXikJ9dLxbeWYzjUDlFQ7ifvD6eD3ppCQgOAA
tdCnqUtack7TuBu6UXkk/o948fl6pCH2Ayt26hf/wSNoGuLIRUYMMvjzKHgxmNF7
ch8NYgHAAZG8POeM8uvd5+ZwKS84w2BHaVDbz7IubZiiAetnP7FGJsALLRhCnP93
zLyMOCDUpS4o9jZJOd6jw7a0qFLrLU/yXrJn/ZEq76tcK5mjwgiMQquBC67mV99K
pKip4VKNOQv37K9RDmM5LgNEdNYvU+ept7fs/kjFwpzYvCFIWUHcPsfaIX/zUGGw
mnutynOdiwT1cWZmeYDMrtocr+GvCxraDh9xLR1ghQVWcTJL8bmwSCHflkGdqrYr
bUUBFfY4Y4OqfLYR8Jj4mGJtOXYeodzGziOq1xf+PJoKDJ8TDjqTLO9gEizsFC3A
wmrdYUuacMKgIRKVv+8GpkShq8627Mw0tG/iL/1TkBWO83+TTjM9LrSxs9dnyc1M
mjr/6L3jraj2QyU72xuKFMhgvm4MB9qsqtOnr83slVw5SsOQGnhGjzbPyPIVbIOm
o91MPO0lT6OuiF+qFyzrYHufXjqD1z4sxv4dWsmNufUzZI/zVYtcwpOPl15YUY3Z
IQzI15JH+gXvo+wFxoVlJEyLU2+SCdUWXUDZ3kKWDUYd7nOCbrxFEdc+Vdpojdbl
0y0nZ//X475Vfdzm1eRKTpv+cpxqx9ZK0WWH9AS6HufaY6ZLUwjnIS6XUOtv0NJw
aq8Z6xCIm/PbYDVTngrmUjzUKqYqeibAQgquQAdLY12LOJLr/IF/ISGK3b0OHZPF
hZdwM0ilZpKDh+0xN7aG4ssdRQvKellDriD39egw7pHo7uafxN7QU6l4rFkNoPUC
ofYCD6sPYaNsJmlN0jbwwp8s3CBDhqDf8AjvRphFsQI+HWLRXB2DzW6mNlJ10k1n
JDQ72Zac6ZBqMvf6Hr5ZE3QZEzQZoCvIKTHsWwjid1Fqz4U0FUj+WfwCDLPJxi+2
Co2TpqqRbAQbc1WUEDYQdRNW9qqeBZ2TD0YeMUOogNnhePYQjdr9NxXBCNxI8DRr
xiqRhxZmamv1TvjRbRoH2O0ff7Ydlw+NCOblAjAfA5IYWu6friPpHQUouLTUOkqZ
w1COmbzhBsmOz8wESYYJW2E36PWI5abkmQOM3grAzRtqvM6uuC3gIWCXXDQjTttI
wbNbU4MEUiWyZusZ4vemxHkBReWDFLLCo4PdAFkAaYFfuLC6V558LzHZaoh35mDf
xsoXXz+RnUBz6EIx+xGp9gvnIuZpro/P5RJtAW63OThGFNQw5hwEsGU+/OnLaNce
plMbHM9tTmPiBTqGvo4Rr2RlXIX1o9CpamYfmmaEJ3anSgU4F+h5Op5JOzIQS+Y5
FgunV/UT99d+OZ0mhUBLua+oClq+gambMKir4kribnqKmV9sG//EzFVExs+Aoiv/
HJf8zNe3cEEny/rP0gkMuoB/JKvCd+V67VcpY/5AaoDrBcnV1K+M8flCJyVMzIm+
l+3Z1xTl61oJqn0l/fEGTFxEiEkMOFWk+uDly1vxRUwxfaWtoV0HmbOvteIVNors
+gbwCAbiSFtwCHIfyoSWVj3cNt0xqqc7Fi7aTvBjWds+dRRSOrkqhxM0VPczhNwo
toB9PP35SjrQo1U4Bx8GqMGfEr1dd1V2KWIkVccYaL+dot6Nu3ELMWzhEGAPffTd
5Dw0xP/3N6wy/Ge77uSOU/W1mvJtXAe9H8Y5rzSxn+jUt0lcORJUPlfgmb16H5h+
FWaw/zkNsIMwGymtathnTc9cZblZXw4303XAHBF0wua8fkBH9LV7ucKlo5mJ07on
H4nPNUy6v09CmJ7BeAA0kWxWA83ySstKZuImNzCShewQA+5PKNuzAKfmTqk3h62e
754gBqVyXa2p+tNkFXGVtELc0K+rQlCUGRVIa7vvj9w+Uq7Ln9uN3sJqGOwE0J82
Jd07nM3CN3E2a+t3KPIo58d/VPmnfkQ89MCnXJFXKYE5SlBZYTVFAWAhPAZLUfcG
9ID2QHpfJuRfkhTfJ6zCWt26AFlYZdfZIHTB6JpOEEESpPfxFPrmx+St3lSsyqZk
GypIp3+AMRR71mLKi8M4k7usTMdaCCvkvBSqIEbl8ir0yzjGOzIrFG312qK+13zp
d4ow3FrjSygyi403uOqANgMvPcEgaRTybMbVfCZWsw6ZSBs7nh8v7XfTl77fuIXL
hzGvFVVdVcGPTsCziIEvJA68vUTDvXz3RA7G3ghTP+9RPrkMgn3vWZr7n5Kh/tJF
J7eLGLP9vD39WcwuOqBUpJvyTWne2UyHwMetpFVabvLnmWOeoseG/R/8Kt8WxRx0
WVY8oyxfgTNrNsYlw3JyEGDEpCUTOOwb9jol1cvifmcQrYT8GosiQsSI08UEan/P
8eD+Bferxug4LRAHUXR30PEtgsx04nQkH6qYK0kdyV7M3Je6w82WA+FsEE2Cw8mA
cNYruxpEdz/C2T9V9pQYUEtkEespTEe5fN+r1ncN1+NVdtCWiSy6DCJPOl4jNVL4
SY9qWV9jhzWPlKlEl/vsk8MX+xq0fwFbEf4ZbhKmiUoZ6F+riQGhDIifKdkWun5v
rHce0W3F7lKoe3VVLc8wWKd4Ydz1KG2UL8e5SwSjO30DuQqDg+QZQ1wIbNZN8hTV
Sb8XBnWJWfeAiaaN8vfjviJGmIuz7zj1wK/1cXJzN94VySsU81Assmeb3ZrnFBgO
WChi0u2sofHIXcDX0ORKKqc5DrM8fdiNpqVZ2HbiJLoVmidBMmwNdUM7xWymM7tr
HM0Nt85eVWF5RRdiJjHi4IIdWGUGsAfzDhxrm6JC2/eyvi5vU+0jXq3PSk0F73Dh
moKxhwIjdgqFktWGJRJJ4kOWHZfCz0KkDCA82xjh4BLe2MSxGsdGAXlIdrEUBjDG
VhP5hmvaInNf77hv+UVYAswImrEnEB18sxJkQJM/WT803t6kcxTMct9Qr2lRcHVx
17s0uQGCXy+32bA7C6iA38mIgWDLgqRuKzeA+p38boq1m3cCvRsi4pZoBizSGKco
4IXEBW6H+LRP0b1WWsDDF8Ry0/kpqTA44/siDVaA59fhE1C1mw4tl77Q+16ZOk0o
oyCVRIqHOecALhffuQ4BTXD5Gelru1G0OHEnsQnDJDA84cakthk5ZT3kj9+Y2p3V
qUGPzsw8XTmHXp+7MAuBaJDsh77yDZ6QbqZ5SUukPXHdKfS0+lSVXIgYdbnvGa52
eBpy1j9LaoffMpXCG15oQKAs/sQv64IwdRhumvesA6kr6eUsFj+KfcyrISfkGjOD
0GCKwVOsNFpCF9IVJaW3oz33Pem1Wkc7BV2RwlQ01Tedxa4ntqxsCRIzQ+QZc4SF
WmtWgjqd1pOx8TFjbDt71gX7pZLLsFnYsAXSAAX92gnhwtxVvXzVCMkQ1kvSnEPB
YrhAxZtpNipGnlD2zs96mv1EU5Emu/E1ynMaw5/yBkjug+1KCKoigxGnMjetmch4
al14Eht7CGYCcMLx3fOc0/Ae8W/3lnCpF9UbAqllxpOd3BFNd2spiz3YTLpqsEgv
hoyKytOHd1cpUFmA2x0cJ+LSmrbvdBj/MWf30UtU9ZeC5hjHxRGRqS4/+UxoSY7N
qJmmpC3zxjxsVKjcxgzFNl/6LXbGDgpbnZ8jRAzviCYhlfFnQLuS35T1f/pfC0XU
MyTvNujOXq2ES1VLcZNiySFImFipMhkiQJzSJr/DzwynAQeEBC/fDaQRT3UlzOr2
KLcXCJE97xQ49cmA4PpwWtT4WYAXFGIUGBqlzv8D4Pp3TGUJ+f85NJn6HtuHuCKm
LdEYnaEiTq+U4rkBtQGkyCfAu6F4nGJv04UywgydMVSkvAjdAjoTA1i7Ot2eEBdL
kj2oJ2RBpOsZelnAdXC7MM76bWnW8Jw8vUCRDMn7iAYjLYmVfUrqJ9z9M+B0B87d
d89wk4dnY+LqZjQZ6/CxUohiu9RHZ8zZxyyx/90U3zR8hrHCY2JQr+OIiawbl9/I
oW4UdhDuwuGw4ZsXG520MgDeMAC8Fk+qWpCi+XEHRwvu4AFl2x6bCPmrxouFM6D4
2QuYGOx/ZlJ1FAIbtoq5aPJWMtC3w8oj+bSIxOjJ5uhg7q8LSFxVwxunwIgXdkwU
xiznSfdBx/Tjamdji3e2xJyFGqgRAt33//ZLckhS8CgRlbx7tPkBU1DilMZkW/vI
FpqS4hz+2DIox9Zs8v81whGoRZKMTO0ZY9+y+XQMacq/tsJIRKUbaTz42rU4HDsf
JRtRzlCvX1XjEMoijVV92mfUXCz6zp0cS+LcuMpYccC8ZUhZSI5RfSkW/mjnfp35
z1r7LpIxi5KGTIJ0rALIEEuPfo4qIIjloz8sFUZHvW6Z35RWilfLxH8I5NgcuyZu
5ektiOtGGbCJ89k6UDtkm7hVXeT6vVfBulDOWZxuOFaOOetfZwqb+XgArdiV2auH
mT7s55nPNtEtNBtzlp4eKzkVpkyVH3lV/fQ2V9zCm39eBr++/BuDO+S1JShYcK/P
+Y+gfKTOkOdHJcu7kLZazRI9sYi1rjtmXkePJcaXj6HtZJdqQsp1ZR1CpB15urrD
VkegObFBrEzfcBF96FIzta1cxd+2mvWzQzAUa7HuXIGdVWQTe0JSRfsEWADTABbJ
8ERMQ+8JEvvS8kkZl7Q2hj7cYqA7Yiw4wYWawE2ETI2S9TOx7lgvdIlASm8sezkl
+Z2p1DNpPPTdl4qktKryXsPBEXzAXSmI0RabFn6oJwZQ5hbbBnw6anSt7uQ9vFRD
EtBjBmGw0JJit+uhLAjNKmihgnriUvMbGITsHl0ezE25cgc8UUpK5jlpib8FbNC0
5peD2RdaSYe5XYWrpL3RRlKZ9ScD6sm3bRrJgdlvU8XAn/ohrHBjiqsVkOT6tTn5
qZ0ft0vtrKIirghSf39Z9wt2XcdlrYs6GGqkPi4mpFNvu1c4X0h1aHy79U5/d4W6
hCm4oeCO3Zp8lpmaKAsJbO0D1V7HH56D998sanFdG5QxPPkGNyc1blJmwM8ao4AT
pqjKox94ERURwlXgF5dtqg6tX/CV079cQ+vgCnvYEnZlO2tir8zGDnfB/OFfRszg
E5fSbABhqa1SiOwu1FVyJSS9KWgoYnTJENcFgMaewVeh972LvnoFll/C7DotLx2y
iFtpFNcZRtdlvdAXNj1q1t6Pm5phYqTMCKoyUV52dQM8DEImrUs7zsj/C4ObTSDj
2citG7EWNtUA7BLZJrezwABJAtUmVtkj4ZMRoYpYYS1MdbCnmo8rnPmIwCpLbaOl
EGPSU9ruzmOvirciAbQwiOJXgaZM7xTmF+ZTYkLlmUB/0Xs6v5EuVt4uoF91Pn2S
ThKgEYBcuDW2auRzapIy3nQNad7u5wj6jMgf6PWB/KSYgVSeI3Aj/SvDdgvVvLaM
8a6p33EoB2KyrQ3KQbVbVjvAlPqAJW+4uPwSmdB6AV5cxMju+lnCwHQEdVmmFBek
3PhGd9DPZvgdWXW1esjo/+tYFwmvuo4yhVC1cQGY1IrUF3l9wnJLXRkbeeqNuexW
eI7vkYTMHMz++O9h4++F6TtyCq7IjVd57GlS+YmL84dd7cyDekJofEW5YH6Bhx2f
jTUG24wnV3NMb+P9v5Svr3O/nk4lgnXOIpg2NyFBcUEPMEHX1GuZu8Oa6zNIXYHe
whYWNTloLmAEA8CNMWRJ5qEik6F5XxKxk6HB9h0mP1YVovyFPATgFQc5fduzPn53
4SvyKnxi0g/uY97pv7pGofMkOZe3YV8OYzi2oeyZwjIQAiU7Ah+sV5OAq/5qvxy+
2egEFXjPjVWGroab3HW0du2463Myo7JO10siP5VmKdLMaf4mjDXHJhcWi90Gje3r
gc1xrnKO8lJ4NjHAApAGzePPhtKYi+/cic9lg9mvMJzPZUGHQwGmC1q8AsFDJoJ3
Scm0eR1Yfgzlzidu240LfopV1CYWHiSg1EAo0+Rdqd/NZQrnjnZKUKRaxrIy24ya
va6i9EgSM2LXRpKM+pl/aqa9CClggNp47371bj0KFPw9NWRdm7mKE5T7+3OYE8+f
K4ZnTsqBDP8TZYS528FGanyU4JUzork7dLEr+LOqWTJ6PuktuJ7JsoGmEfg+mmyT
mJt1fCOcFvoyJLDAV3ZoW5qOGXhVDlMXSKF9XT/5OT89m+BlbtbCizLbj7/tEb1P
kg6gkJywiP2lYtJ+TOyCMkCqA7VkYmfJk2H6TTHGcRTr2O7ZeFXnNa9qfLw0xous
Ob3JiQ//1MKlWMSZRyrh6mrX9XAmeYWnRM5Swa4sAyoW5R+LoYy16CPc5va6e0Mj
jp5QbF0NLDF2ErVnKxynbDqslvVUnhtLMsI7R4le1utVUtTI52tK6/WJW/mvkVI2
jowr1ddcbBls9Dv2RzUdpYY6iG53AIZdyhpcQ6LEhdnBtB0t3jrsuCGQdqw23+n5
+D1TIHgqEp/qAbwrCiwA3H/fUuD0NfkoOlD30BMRiZmLNZPYn8q/XCqXVXcLqZ11
pYoMFZX4syiw44oUO79uBOVjkrZoF51sZSMyxl4fHRvMYIjAj5/5/q80FL3FFbbA
C5/X7uKvA+55o/GH8ExU9+dZtSkCmt7RKMFN3gukA9QvbBCvRhaju+0EIbtZSgxh
8/a3lwzZfGXvrUNqb2SCSLjpQDctuqtqrtGcuvACGoPZEYfZXsOJpo0DEBdsxeAr
M4smSGVob/APhB/R/10mnNH7u7IEkCx3BEuzxtEG1VlSeGfHlJvphxgPHJC+pJ4H
Awjl6jZqKRXQCizUzN+xwMGJEyShM1kq+d2Kub3OHxCIkjpLIED96NM6X+H7WESO
WgQQKcl9BEbEwNwMg49kd+sRJKnd4Q6Zag6YvfXiN4Uu7YLyBdy6ZMd6w5nMs2v8
0y1o+1vg3GG6d0qB3AL2jkQ+9blDqHG7Gi0Sx0eLpwV8jZBuxV/tI1hBKxUjpAx6
Q4SyOI3a0/eVaFFrir4CxmUrqvLgBAlkyqmy4SS3YWHoiFtWbVyTR6nw53JvgM4Q
rzuW+gb1YyJmnA4B+62LoA/a5dEUSf7BVhk4+gLy5tV+uHD2t8GHVtatSQf9JB4z
Z3P3+9u7cGDg9m6NdtXXUPF48G/lseQVQVCH4tjjbTxC67kTstm9Sunw6Obl9lYI
kwDawxNPdfFItgwg0jxOXJgvKotFiW3hzBcmGX0hLYyq/YxtAf9xg39g+CqobT8A
0JuWFxo5lowXKin9A9ufuolI7MTGlYPkD2xzmMVyv3ebUX6iM6Jqp7JadHpS8kb2
2HSDlae4oRky2RSnPGr/Hv6IX6c8gzAEL2jlf1CtD+yGUL4aoXXpS6LATD1ozkT9
fLeSEs17adiyp59P7zxdVDIrgwwQwEoXWnmDTb1SSf0WVNH1jK5cT2yqP48BVx/N
pNFFtYNK7gLkgJ800+Cpj8mzB3kkeKRwsCkAYWpvyhUVWfLXvSsAfnElYaf7p8ty
0E+9E38gzxcJ3L4XDHw3Jz218xSJ5qmqN/aJjnfxgVC3x64rDG8vavZb4L+vgSwK
J+I54yzuxdkTRtTI9D0XzMS2I6+9+i1LJrWug6Dr5WhyE7REW2Pc+WYYfIg/mHEG
sCLxze84DQJKKPGe+QwOICQPqq81VFcaxodOgKF1cqUVwPCUOY9Zn5yFMT868PKR
JBmHFECUkrKwKkrvieTG6To+Ciy1HYJo+Zm6bPKTx7v6qTlXfqLT/qnC6SbiVsvM
Rybocm/Gr5VMO4r32r3zXU6WiAY4mMAiT/c/t5pqHn/0m6cGwmcpOV0WF6sobUvf
/3xqhQCqqvxZ6wd84UNCvyT99aDimDq1jaG5OBmRWpeSJyELVZgXiKFRNIrASYlw
MvlQOIoaBVNPQG9i3Ynbphi9UuSmEXUO2U1U4XmyQuHIQLCbWuAlNCyyySa/l8Vg
euT2moEDuU3ZFCZOSuarHPGZy2zf7c34yfWQkskT8xK2Pw7LPoMAIR3GgGABTWRR
JI9zvn4qZz8vTximufN+IPCVMHlHFimYplZdg1N7S+J1zIkjoCv4+E+5VIU2Vwqi
EIIOJ5dyqjno/nhP/ITWSF7uPe7LG6nAOXiBJmgnwRGyIS6RsRgz27e0kh7cuprK
accE7CUDVHXL3fESNKlYgiMc2XTpclTFJtGZHlSU5DBL+JGNTorizfnn0ZqpMYN2
kpWvEbr96V2vHEiuXdpeqofJ2nqhGVY4O/EyC9RAqw6UIHGfn3QMQTZ6bqvblRxZ
lwNwj7rEMUn6ERnR1UcvGTzOdXw9alglk0G+9dtOMPjYlm6LK+LEkfN5CKcng/tk
4nnJPskaDJrlzPY/SuDg9HKFRae27v8WjBp2ks6rbxhlZFzAF2wllnqh6psZnGo6
7Q+JZi3OqeMKZiEn7e7Iot5HQIgo66RXRcd025Uqvs+lj9z87gcBtd9hOG63su+U
T954Zmcxms6rZsJlgGG3M60mCE2H1WDVCVCYcYU4uX0pOq7yagfvr8QorwO004VW
xU/QyxcNpa9JJHAOleToG4HIShElpZ/khjQAtedMO+JOcwlPWKcqnsfZQxgWvNZG
ISEoQMOCRzTexLvzfVc0pBlsr4Sl7/pjhDa4CiM2qHksttkpySGVgH12vBjzWuBN
XySQH++RySWm+bKp6dqM0ir4rd8NDLg27FkPzmWhX9Gzs3tIwryfmEXFJXZtvOjc
WRuDnAbL4sDoiAfJoVFW6EtOmseCbXADEG3Dz3GejxmLgo59ql2a7ivS2lC7/Yn7
lWo/0PNDyDoztv/q6fUO0K6FHHF98ne1FRdLq4gf0rr8LIY11QzsLfuL8amyH7qI
UtPOvHYm9RiocXezCzqwMtaQrQmRfQRhs88A03njTbUCYaXxq8UqJUvwh3VQYwBz
YY+uRavOezERFz2dblZhd8+btMypGuVyqAlu+X7R8CzKd4XGjCqU4xM+GX8gWvGR
szfGnvr+IlfM7bOj+U2hpvswGmq5/KjKxGOdeesbITYYpSvQgPetcvY6gq1H6Eap
n+K/dox75aJ+ZhRorHIMUch0zCjuOXfADb+hauA/3Ih/jlK4mqnH/1riCViewOFr
C7Oh5CfCwM0BHT8Q7zQQ6PdactBlqnSHmo79N3+DKULWRDhz3MxruypdCZJhVsGm
1Xs5RJS7UBEwKvnUYEO8Fpqcf6g50fSAjcJAzndaFbemT9Bd/C4pGXM8ZiGL6Dnd
W/LA7VgJyHMry4LXGTMnmg5P5xR96aTCcOGCcF87Crnk/MyeS7bODudEXBa2LKTh
QNtakq3yywaAnRNuliprVli4c+H5zxD/1XLJ7f7scvQaz8LvPwdrrK0hsYA8bsxg
eaJoP5PtWNxooExTryZfsLJNC41n6tQDg/20I1Sc+hBl2uM6UMH9QG6RPjnRN/VY
zEatjp/j0vBDnyjBr8wJihOBjZrAewaZkT+AvZBFtL2oAZmQ8yHIm4D6uewRI3UK
2EadHPYswOvWGY8Uzdeqxwhkf1rpS08Nr+AZEYlwjP5JlGle1LC94VujWn3+glmB
zeODgKzcIakUySKb0POCgp5d3MNgQq73x7gJDx3xvJq0b2zgx7xp93DcM6QKVpyW
e7zSZ9zReKrqBAfSVxAoCKfGlOyetfQqGOx7oX1IfwfgADLPjmJaLTgIAkiCnwW2
hOBYhWwyQShPZs/fRKwUCxOo/e/tYKw7H5R/nuuF+2yj6fsrF9oZPwMRNEObtwom
9LHKgPAtbczDyD94l+qSnESrVKFkWs8tAGukWiXqtZDZZjbyGkbkXDF9dRSFDLft
Ogo0m17Xyh5j7M19Nsjz+BHEZa5dP+BjAuthknw4rVnJ+JnskXZc+q9V591hwD+F
so6zPkLA+N2fQ7L0JvBUi0SasPqgDXmcR0g2Hib9ZC1ISdhTrMoI3BiuBemtHzQG
45p4JqVTej71Ndo8mPSw/RKVYNUzj3oy+rfw3156CgOZpSwxV96wzaqeqXH3AnPS
KZe05VEBXkSfPGZUVXhU562Dt3SOBg9LQdkRNsTdA9rrzjeoBgYsuaqpB6Rfv2tj
MW9K17dmAhWExEuFwxPG2TljVOajivd0xdIpEsZ8/PZ27F3FlAKKZNwzgAPfVaZz
WrBLg1E9LZ5OPkwlxqYeWTwn5IPN0qlyOd80BRVFDoDRudAoinmFqv5LBZVpAfgZ
83FNoe1LFwM/8e8JvM4EPIV3A2Ts6eBL+TMVoyiBrXikVNCm07d+lBtcIsHWpJ/J
nVT/Rk4T3p+YTlY8TGszNcqGEtypIgTJt2LD3hrxuS6ggSV1gs9JOX7RD9do0R1K
FsfMfMMnrGQXdHfGAa2dRTI2etE6clMlT8eBpAY9bLyS+dj4yF9+NU73xWxazAba
ySS3NZf5PaMq9GhIzf5xK2Ab4tQIfvm36l8wqK97XiCLvxe1Do/uOz/vomT/VXfC
WTMb/NjpDe/rPSSviTC6b6HTZlwhqSp0Li+wuI3kmMF1BGKwofbKCLFyOMzJgqHS
C8/huEtwvr61AdaLKVcFZuggLZD4FSB8AeHYE6UBRo0a+KK2dFAp0p0oOMsAS4AJ
JlfHHAHf6sLBgg9qN2y4lRK1IMTCGAUdQZ67DPKZxH1LC1Nj6t7w82OK345Q6nwD
GeLMoY2LlV3wu3xSqkFyUWSQdcUHLeJVLsZwFmgJzvM5nTSVPShjgBwlt8ilZgn5
AeGI7X/qA/oE3CCSUJeXMQYa/bb/YNf15UBPVgGZ4DgJ99PX/EvyOdmmJ6ZeRggs
i4kzfxfbNJ1EQhOpx4DhcP6K451ssYDS107dXkyZCzQAe9fp1carF4yJuBioJ8Zo
OLqti2fI6OGuDEcoeski4HJddT355dYGdRc5+3OS29PA3H98Rjrh98DUtOoFmBo1
xwSFVH+dOhBT8ndccHphUEUif7XgDjhmBoyU51NxB1JW6BPnu6U9xyo2DilChLBT
4nDYlfECPAAq+B/jGNi/1oxWoP63322qdWaHCtmMh2RcsdK50Ls552MD/wu2mREk
rly9XzAl1MPgHFdycf+0/ev+f4d5TtILI+m4el2mO+PgxZhrYKCHjRapo+LnZOUR
InAfU8GaXXtUg3L82HJyTm7qdkoyWpT83YlkSXm18lKoMZqDVEeSuGQKNdICKYJZ
AjaSO3HjA5qAXA7AWdZ/bbmx1yGRqn6UoOGWch9qOYizNg/la5jRrVbEfl/a1+ez
1maOTxd2JMdpeU6DuBmISvYMqqnsfFOwkTwNIVexv695hJmGlh0xLbRVYS3w3pZ/
J2t2B1Z+j54vIoni7D5paVh+f3CRGqO4t7gwMK0/mp0sVYw8iClwvNCApbj2JBlB
SRH2WkIHAfgzF9jaCab4bmDKrWoeswn/Ek+F1+2KmIcYqq9cwriX2Ecl0irRVBZK
Ooi+H2aKxlwmRuV6z7qZWU9NuzBF362oykSH1jqv8x1Nsk5inHail0I014UTF1EM
1wAHW6eInI2fBqNa6t/+6QWiuo2tfDalUGFBvfKyx/NRodZ00p/kcMxhBLq6eFYP
r0a/ybC0fwIJbyDbaLwgZuxzmlhwNgkEGElASFHJ0WSDLeXZKvkVNvan34CT9F5H
b9RQQnrlhOBoBCWH5zH6QIYZzxl/lkMajI+wi43z/AIsjOVIf7OWgEXGYrwPLFOw
9y3/HMqg8x6dNIM2rzfyTQI4esXHQ1Mf07ALbNnV51oamWHit0q6NTn0D1BfBoqr
qkfpfSMbi7Q0CPiGoro/qvjgajBS6yCqVogh/F+WzDDYfYh9sAHnwi3POliUNbqt
K0sbcS5k/0A7nbYXVvVmwrGgSegvNKzpYGPL/V1cRTYooeEeOuC1J00zopkoSWcc
IJhIq3vRC7JezokMJ7iGIpSCDQnJk5qaSIK4SHMTUVG5YyUDUebijCcT6IVLiGRq
aDkvUdGcGzAqBXvJNtTcxC+eZiKtMIy16gL8TTkL/hfU7srcZ+QtWyAoPW4qZ/il
exymcmmhMQjcOHFLpJZzq7qB0e6H8k+d0uD29yH3yFtIjHVJnXZFX1wZmBoUn+jB
V/5QHq72ZMTux1dgEc0t45BN9gXGam+Qs2TIBrLBM//jiGq2gcHLvRVlahXYSn7B
cdffLgZ6phKREIBgS7srD3ZaXmRy9i2+5M14O7YgUKaNuAqCtwz7zjqvqTdyNnWZ
Zr1SVPiSZOirMKANQmbkNi9vu9w7V6BFI/HY34omJ/1xIuS58JfOC1jxcyG8MX6J
X3+5c8ZfuFlgpkhm+B9Io4qJtN27avz2nwy72ZzffE6CgtIPp/DT016uxONfp7V0
fpOUyQMqynxHFxLHp5l0H1SxFSm0A1tYTbwpxRYQGTn2f2hjC86DHqSo+Cdn7G/f
ao4fDCPzkXbGtWD5SAWkiEBri39+zrBwWPo5QUcv2v12LVmmsSpuBXc6BJ1WGC4C
hId1FNGo4KrCspnfxV4/w783+aetOasiKDALlrnrfRbckww7EeQkxtv2Vh1NwSV9
7LujZ+9jN2A6zfQ8zN9XIRoiGgzR7Xz+QTGXJsTQhWgVk4CMwA3Bg3sK59qfNAw4
DPoqDnr5HhXTDkyq1agGiOMs4OucnZeJOyy6gvrPCU+Y6+y+3cvd8Y1odgH/yVLV
2Wul4YrhsXbWjqtfOFpedEUdF3SAl44Eleaz+Vp+iz/Q0Dl2v9REbWA0E0HNNIGc
GdnH+F2/ylyH6diWFznT2vtCxhVr1r7VYDkJ5yQKkxF4G7Wh7Jg8P4aDMYaf3qVe
5EI1lj2/IKqwiDEcuvDdgHWPPm+oeEiiRWauDgQwa0kDrg5+u/s9tPlhhQqqWI1B
jlpPoq5iXOHs95dqqrO4xccqsAnEUgauMLO3ShIRBPe/2DrUTNgU7ZjzrQdMh/38
PT2s5FrwLucIpqCOosJG43QovOqQgo0004s0TLr1vfZd3ASC12Sn/uC6qiZk67g6
n4tgerpcdrzAJPSWGupOtqKXK3AyUpg/RhZNz80rquxPvHalE734LJQK7gFMcwiz
dzlC+oc6+XRMe6DM5HhQFhs0j7q5ziPtQgvECa8SdAPQuPLF1GsdcJtwLd3uiaad
vQ+fTailaj3q4HhtLl3IHhLTzXo+9u4iORaAv8Hms/i8nRpXn7e080/AizOCnvlF
yCqMWjMGtbiDavVIB+8laAI1Xrw0+d+DavI18IvNR+4E63jJqPuWkqDK+VYf8U8w
wgZUyWD8l9ZcEIGrlp2Qbg8wHYWN85bPACliH91QCmvBvoU/cz04TFlmBVqODlbR
nsNApH74PjASPk8VaAUTJ5Ng2C0z3FoJLAJKqnH239+7DnPhgrOlavj346R0nF+c
QZ2MGJ7bm8d1umEf1EjAgWzmA99m5NQ7yRMxGnOz86GuGyaF/q9dpM99dd3Ao2y5
IxRzAWzbReGp0SirhnwBjro7XDeB2x/fqZYh6JGuoLHyziv63BtIWGQdQceQJaX+
WnNHkOKeynxUopsM42DM/mWBMxKFW2zix8SpCJu3lkP2tny0F41QJLcw/wrKzqo8
7zHH3uODkDQA5NSXyb8NIVHJ53STkPRfuoqXHEt5z6LeHvzaxpn2XiWFSuuRo2LR
ebv2s1FxqOScC7CiCPLIth2GEyVE9DS+bhT/avrpynLPHufxY8+gi6DsIb6ZBgKa
nQsaEJmI16zNubibP+YcS22GK+rVp79s7g7iIkxLA9ktHgIAz53JQDmryOSRTsQV
yUuWo70v0E7CQjc5QsQWlj+LZLw38t9VlS2zs5PJ7qQmfgCzZ3tsRck1WdVv2x6C
JCzWPoyghBeOT780eek+UOTwiQZ4Ydbye8ahaHBIYnWDIv8DqoBQtWZYKcE+aPnU
JlUi3ktaY+dz00FKQ9+WmCiEPxBO5t2p4oaJC3G7vdV73MJ8K59QAOLf8P5UE1i9
1hYaA/Rx+1inN5SjjTFSIic7j5VFw3mkuo7vZjLJfKonAO+zxMThCWoiyiH0kzcy
yYGTuwAgyU4omOedx1wf+QVpQ5SEYXXZBS/gtZYYgBOYFoyGBBndH5NWua/0BsY4
w4trIa7KWgL/4ASxScrXtXWeqhef6kGEfkOSOwPIxkDqdMi7dKdCfYw7zperWvvs
SFwNj+O024zBaiyVSVvV9i7OGH/8A7oe3CK0T6GMTAXYH4uRkWhrt9UTvzZN2CZu
+tZVYcJmuYY7lT2qQvtF1jRvdi+/IY3RMAz397/5wkCizB9HL3NLgO1bV4L/O/SG
AlKFjRiNsvQS/gUln3yKO3yW4bKedXN+eZTn3SdBNaJGuaT0oDE3Fh6EJQY8EtH2
aHwVtKxB8CA/5v/tjD5L6Wrd0bV96brRGNcP3gt2zsVcB4bVdyIsvPoH05QeBaXl
h0j/Pm8d7+hQdfgM3c65rAQMO7s58180BLfngjPQlOibL49ewIi+8hNl77cQ/0uC
Nsvy4orh2VVymv1+eKYc4+lFe7Ddue3zVrvF7WU7h4biRriEPihAMYu0WYn/3Crp
p98qxTRQ6xHiNjKciTMbA8CyFWLEVazwG1vAO24TfciLfSxArVMVptp1+eGyPK8R
ZB6HqcoKsF8qJi8lK2cAq76c7kVC00LNvL345MuUZNbjrDMFgCX9yG+NabrZPFA0
r3QyDYjzyqE2SbRyvQX18g4o7Np1PeTVsLtl38zR76ZFUmrydvr/XvOu+7+W5xXE
vYz6RKpmx8dXWH6ZXXtn7rG5f4UNw9j3wHHivoJPlS5NqH0IOoDSfdB0CVQJxWSV
5mGXKPqGjkV9HvWq3p7rdYusfzKeMPDS8MfgBNESuJyBNpjIykHoipCSd7xndUg6
T4zLess2QjzObd6ERHZLo7C/byHBDEdi2qXxaKTP3CMYfKVWwVZrW/M5W8JREMTH
EjW5O7UEKB/+rPWFdlJ4kCUX4s7HkqB3T65XqtukYShwwSuPxyInsYYiPFcgQuou
3khhw1vDFN4H8eO14RB3pqcDL0ZlyZef1zVAYVCOaTtF8GYvIgu0otuqSkRePyxk
ALiIVqKFht0wgNnfB6Te6nF9V58GCmOMQFSYcJq9wHMRLdwxJ6qCgBvU0GAY35aS
/TwnhgW/9vpIUCSudOqmXVwNDp4X54gb2Tq3Uuj1rW5D1wSq+ioqQRxNzLQNDXe3
DhU9RqdLhjZOeMs4oHV0vXc1R2echqTDKQBaJZsH05bkcAOYH4GrMHsS9Rxa1yO+
CTZSqxxvunPqUCAIT0GzjtuvrK1ZekZrt4HlnZv0deVHdpFVDU4Gy/TL9NzonQbz
QnSOUadNowhdhDKhZWuQCuc/ys/yk0h4SYpT8qwHxQZ2V519MWEvn7Fq0VpBJqa7
m2bzd9rZjLuVpMEzY6lYmZ2zTG/Euo1w6X3T2t2xUeQPvVGc2wNFW60HgrX0NYnM
ziOAfzKVvSeE/dN48HmUfLbWXvyKISQScc/3hM6ZnLouNksU1vd/tMNJ9RIB6GZn
lzpQg+QuJ1EQgiEmKjsBuNeGD40eGpJAbwrcj70BuHCXqHom55/dsP+FiRynkNHr
nhcxgLsWu9gN46N+KDzRUTV7sjTftDUU147dXOjdR40vo8WtpUyzOaUK9djczJSi
UG32q23TyIwRVm9Uny6OZZlEMuus9Am/4ryIHI90M2mNqcP0xaOPHphU42yxeVDY
doHspSaxeTsdTCe1B407QlLKJk9pEIHH4s7FOk3P7+rndAjP5Zc/pHIV0lxHQwCf
RC1TDnqDbz/KEb8Tb30iBfs2nS5Y0+864haVuVCBwZHs2umTxT1+oB7TaPKJzzkM
Ozsp20YoPeJ4unTQrFxG0WX/r0VoVGBpIYNwZCazfZ1+j25Ysv8puJLhdSIECPH+
CLdWg8B3BfFyzu8hySWHY/hQSuAOVgEtx1hFcDP966JqcbaEmUQQj19QHeFvk4vg
TP1AETG/AXEAXb8y6HXTOB27z8gE6SMuQULM838Dd4YnOe0VsNoiCAl238TYJz8C
tzfd6y2QxU0htVtoCDlVcyOauRhTTBB7Hg90uqyp3zsuvCEp8qEL0qrYyLDttJdN
GPvbOYBmtD1Tfjz1NyP2EMIiupifDPCjP1Fr/nfRW+RcS1fw1O/yS5drWt1Q9NCT
yii3kTj5oPoDRbfeX9bGH8Q+0BOyIIl3OlxONp8SRvOxycLfxcYpIRlnBg0kI9ka
uuKEQkco3M3d/Gno7YY/k7tALtjeovFnzZuMuoI+AyhDEymvC40XA4J0DQh3HNf6
Vt3/HTWUb9uGU4oP5gMej6Kp0PWgm4Jmtqb4spOmjl/3pb0p5/OHjVToYy14Dc3j
P73Nrecs3NS/qbLIZ1cy9tH6y4X+DCtyCS/yOsBWejpuYqUpThTHVLSpTUUbPS77
KGIJTLls53oYW6UGiNrJqx6AEv7+qGGls1cl6584AoTx/Dy7nwz4hycKBfU7okxr
8Z+pQ/2/pU4A9KO6YsjPdGxObHPzC1SdnPbD7tvyutteVzu5jSW3xyIU07skdAE+
MvRjxlBpbHu/DfbJ5r31bI/7Hk9lbJaM/CwSKyqKrC3QueWcYi2ZyYAl/wWN6QI+
egH7HNuJi6bbvDm1kBAQXnGSqGVwDc212Qt+kBIthCauSlEixbcfzJiDMOXSBVX6
dJe+3BUDQp47BCWzGTd6I0EhWTkAkuovMGHL8oVp4Fw7B2J2kOouUWgeOc3jlY47
CfSd2mkAawAd19UX/r5AfDOOuB9lvs7k34UvsJH6sT5pXyldSzPCX1xXL4JyafSX
Qo+xBFHLgS8Nx//z9LTZ9dEyTYw+Ru1guCdrEs4ejMUgJ7lZZbrj6pDEEsOTk9JD
jtHgjWCsVLXQnS9TpsqUeaqFl+HacL2mmlGQV0wICF5ACNdxwG84OEtmlEUnMaJO
mWbjchp0Yjy6mJDYlK1udSpB0/qEmqGgq+HOYXh9gaGEOzDqoW65rFDpL87k1d8Y
PkT700dctzDuOt1J2I12a18A+fqVY1e0Z/+pmK/jwDkd3Zr6pDcS4LxUKugc19J/
4j7OwTrZW9aEiMmUy1b++WP3yrK9PBr/wn0xwC3MNbNrLOhdqkAHHc0NYhmpaNbN
mqELLlwo10muCO+TNK1lekkphGiHDUaFtBYL5Jaf5AWfOeMbfzWOReUBUkUqkfEv
CkhAu3TkQrb9YSSzi7mDRiHm/t4vA84vgKMBOlmA2pO+SWB9c53EeLwTV9lB9hbh
mZsUHafQWvy32QrvSo+2D/eVwFz6v/YBm+GeB06erafYfkEjlyk7+Kt5gDZTjCR4
+vNmxhKnno1BaMmFRd4caNz0pm1tg6FcjllRBrreMyALY8jFzB+8i0JUZ7BvNgo4
i095j+UKWeZiAXPoVXG8C9t4ea2W8xyq9T3jY+LHBR3pxI4JpPGP+La6BJJUrvzc
PiHzLyzkwwwpMQmrogzc0ghpZNiBikENOyQ4gJT4tuPuCm7u4mPs/0VGxsr0xfdF
Z415fOItnD4N1EG5XxUhfr5aKGJfys0tnEzpkinY+b7dwbUjehGQsGcn0dQl94vW
G+GeyIjxZ05UXxKANdhQuGdgzssPLsM6hk2iB2KJ5bl7l2hExaR2DRZMWpQ4pQc1
M25iL7DV1z2C/PnCG0BNtd7jUjQ1cvv2J4vcKXiuLNqgAlMnKjEUu8Ww7PiguiDT
+PDAIFb8LRwAKl6EJAUVAywiXOhJ33r8XrrgylbCRRMgzzDIuAidRuoPNncqiQSw
ddUdRHPXianff/V+M4gVbiIreIuu1OuBiqbnz4XYpT+knv7M0ADL3T3sVz/HCUO2
20m2sSUktHRLcHWh0fcUYpNuS8gfN+XSZ+k9O6qG1Zr09tZVWAFImrwGBzsd5HCz
3FnPevrnqAIyibVM2HlIgPZE7JAEGIC4zpFdjuVzo4xXTQfML1OVTy/EbgNw2lk4
ZFECm1JiBXyzKAEnoYtfweB8Q1oZBaxU0Y3wFMKR+U81pUeD7w5mK6ELDs6yz8Z8
W+C0VZOdQzfqM1rmZpCQ63wlCWjvrxHwdz5D0N/jnhFNFrq1/JrAbYRbOedY+IVH
HjdGkI7fn+4xNPFlMhqPiNv1EskuNnarSOBSpb0VJe88jokXftNmYkPKdba+2Cwa
0QylaphpfoPP1WgUhbNsQQ/55D+s9OnFFNZcYkBxX9/3IW04plHaLsTUekQzpzqN
8aH7bax0qCvM0aII4BMf5rvisJXGtrC/soFQS/cIu0rw9w0HVb5g3F5gqXbMjF0c
nHtr/yzne8UI7WXBBA3YDc+56Z9+/BNZ9WJ7EyTPn11uvtAjE8fZQM2bNp6doLz4
zZrs0ALtGGyLDv4y2wTwvpn5NscqO2XX+Hy00qGGdrArpQzPVyeV4WSsrVTVMGB2
cCQPs3+4pwy9eDN8NV+dVtWwk+87fAM7UXsclGz5PiH2tGYcADz9gegaPhBRcTzd
1w0TiiTg6SsOfpnCaW81j0+veAELKZwA967hv0a5uVGA7KHalvCPou38rHD66uwo
NpS/8j4BLbLdAZXDJ6+HmMTYDL89EEniBur6Cs6T4RxfJz/ZInWTQQp0AA8ir4OQ
SglKIGYSJkjbg7HZUa6cN5TnXE9IH1/cSa5NAF8dXQrcEITqOoK6xIOxm6XEl8gA
+NR6FF6JcWGtfNVi7SbQXhylAWWwhH8p6rTbuuo+HHffzReeqxajSZDgJXypnvLy
DrK51GNOjTOcMgV63kNH23lZJ79hYhyZnd5QHfyGjc/nlFkmVO7vkDmiSGq2e9gO
RlW5pMWS8tDKoeZ4/NjjOtDCBTaumUhw/P0jaRpvFwKJNTdcCpBdm/IVpaD9udk2
axoxivOfqA01jdqmNHdZc/BVpRSIMhl0ZI26RK2UE3uPRZn5FfbgdXcAQ2b4YMVW
d3eUNwOqGEwPzf1hq/5TeA+Of1SMrfaX9gYB9Jpc5ZlgRgCcq/YX4JQPkdnmtTwr
7uhHWyYNdWA3jyQxLBLHHjy3KmP0K6N+ly6IFGjm2Jg+YcV6/alyKAeg/PLrd/fq
y0O6CExpel3e3hJmigjCfxIj1HvR4Eya+PgbgEIV9jayecaoL5eyzFoKRqbgqwKt
ao51FLzEq7XmMQG0jT8HzBrS4hEmkFPy31rKThK0+B8rQsxl8CB292lsZF3cAwGy
D4mubQJIVZHXQRWq/qYWM535qc4X/rW14JjRkcR4AG7fWK97m0OiSNrClHso8CmT
K/mVtBFd/xT1Qux7wBhoHTbxixKoWOiMGFFWRgB5gvi3EL+tf4DuuugBoZyERdgp
ArynvHi558/eUa/Bcdz3UOLW+7duTTdjrNKnWl9VwzJXoXeqxVxb1SSlpJ1uLW66
MbcpMsww4w1i9m+wRRFn420+OBwFEScoxbntmD3bP+qKLzVPoac3PnQSUYGzR/UV
3k5m0ngxytKZSHBRGK0JSuPj5gY7gcXeqd+9N5w/j68cTedAVKBYPY1lk1k72nlz
9a56tNQeXJ2ECPZ1B78fXXkWHPqStH18xC1vU2WMC6ng9h5oaqQVlkWCEWIwn0s7
vLNjf3Ia05K14NF2/fE+8a5CPKBZLxxyrNfM1x3EVEmy8DHuoGqkDDfbmriINsm7
11ad+rGtZPG+H6tk/z4t2uIUeS3WqM2paDh/jhtVgVPNmzKdc1L/74qRIZWJKp6T
lsuEu6DcxUz0b8vR6K56ydKeHvto0FO28k72LjLE/bffjgQq0AsBcWb8GTGhLwZN
E+NrGGdzrVKmvDqw3MFxF6m57a+ozR1MEOYO6S/eSTLavH60fMaW1uip/u1JjYAC
tzWBi17JCoDVQFUQyhZVJPy4hetfRjBU0Ay00KKCMMJQUu4DofuxkE0gH94ROQej
ET+SIOUaU5qLBDjRfds28DO8zCbAIfYQclW5aK3yaanhDOvGlscZbjn7qOBu2qa5
PufW1CZCP9UfmlHHIoWgirQv1BxP53B0ajdYxBjMZJTsU7hfLbgNTUvFy5+IuPvf
IMosKL4mLhJfWA7al0qEyeUZJFq0/kYcqkVeY1QNuZyE6tPad5xg3ekBDUQ3M7vH
x/c/dXat6iw5ZDR+zAjPIhlNcL9d/dMsGegC1TKFRgP/HSf3CAx0JFzfy0oly3Hi
/Hze+4gov6V01M4DF1BQUM+UbtjA6jmqpbOaWJoWxrPwzN2kU2POab8yJAXKVzi9
+nkk4QTIRJe7JgLkzEWolScWNoTNZR4URW2Z03afms3lhqUbdynQvGzOcxKGQ47f
OTcH5IK/+C/ET3zXP0+6iXWGlxXdVtCdY9/oGHSi+m0tCGTe3IAXfwHa3i23izRU
s//Tshui9Fy3RytIUZIL2hSN5FKuUWn3JobcW52ovLQW1lPTL9Flbx1RsZxSaHiE
gZGQp6OTpma8EKa99KRJxiyzN/xDey0lTx86W5913lRSEb7A980Du1iYPSMWcKt4
oF1L/siFBL99DrOBbxTD1NvBFsPAZpeQXlOdOwGzyjhp5l8F9rTTZzxqGqAUMC30
xBT2QTGb33uYol5UF4erdQtfwsc1RKfZgAuNNkBdCSt4X5NXliJBOPquSm21Yctc
uoAXVCqy51f8mFy2Se8OXiorBORHfw6AZ/qlPohoM1/65Qwc/VmJOp3bCr6ssLJG
yUPKKdbX9YI7y3Q2vHqOJogrGZXncNwbClgrrJWgIvHbHGKkte6ihhcWZvSEYPd+
KmFmaWEd9URkn71ozcG50pmbkZ0dakILozDKMBHj/E9q9vp03K5eJvpZd5KysvQU
WYL89lAisktoYEIswh3jedHwvYAyJopSOvM0le1uax0LqbW88JcWxxcv+EOQbzR1
XsBIx9cKf4l6jIXZSRnx3wLzP+z9yChB/RWlufOrYJgjOuj6QU0j8DkkkXm4IIc/
4uu8d+AG5wlssh5cqXcMfBOC13VBAIBPGIJ/4ZvgHBXGtwBXt9lGFsqv+rEyAyQT
LZAGrb0HH5IHmkHkyHLEpPXcIMEn2APu7hSK7djmgbTC5U0m4fJkGh0NvF3I7944
pQVrP1PRUbhOuz5O5ngKxTJ22snOt32cDkYaM/+ObmLQNa1LVF6zujWS/kl2Qor3
DoAemsjh43kkAsqtuJ09ouSx30juyrrq9EJmmNlwVP5T6oPrdggkSd4FOr1rhHmZ
SkJPEvFEhKMTBx99iznfTeNHQ7/edLBZWdFQVcYJnpLEc1Nz4sPU7nJLuN9bPYGC
WD4zByPWgKNn9R3udjrtYggbSv2/8ppnFTQq60xwMFNunPRmXKQ0uA9LScdlYsaQ
nG2Z7eatEEQ+wNi3D1P/6EEDGdZADV/88kfTgQYXJPf0blQqos1rlyk4m0BssB6C
9AfqgpVdx2R0i5DRWn6eO2OT/Cy+2h3H1Z2JyY9WICwL4c1gwHfyw1/eQzDsCqPI
nlmEdpCP6qcaQ72w7nyW6snP4C0x1vLtaLApMv/Sddme0gGri7ae9Q4F18GRNB2b
IyETRlGnE58NGzWkuCNPGa+DHZuZKXT4cDDtWdEZzZbJnCToNdVF+dnUXydw0CqS
0D91PmMy+Id+umwV95br8t77DVYkZtxNmazR5nAo8zVXiFJgiVxU7edBYBlYnmTR
bsfoH09CPQNE1lW4JW0aXb6G8N12PbLJ/m4n6FodPV2wuz3j797ly6TJ+fF48Dc4
AO3a/skoQmhwJPmu1aczJtwKwetxTXmnnSTPSEf+aAvhubIzIpGNBeHieDwTaKu7
+izQj2AAbEFesxj8yySdOPOKioq8HLYrbYKtPrguXawSRJ+v4okYQzdlIoM3HR6q
Qk8EpFqPMmhx7l+Y89x5tsD87xlsTA3DyS22ozwedX90bzplaUTAviw1sPJlgjtD
vcPuEPYIoQa+rX87e5jRhB9dR8W6XnNAqscDC9ANo14U4A6QoJlVu5ED3wTNg/+g
hv8jslYou15Ug8VaQ7YoYARcpUPjnkoeT3ESt6DsG75MT/n7yILv8Fn7aKREWzpo
kWJYrqlx3jQoPuxEWZe75Ro5XXnXRemojClg+DS36brtZUyF924DDzuQY6+4sobo
YQKq25lVXX7HcjgXlzWsAxWhkAHiZtSxUEMN58UcRVR+0PCPB9wBA5Nx760vKobG
O6ChNzpNB0qP3TMuxbIL3v823MI+7+5WvaxxePGbIOAccMVRa/nm+YI2Uyzbozoy
zjLwUDyPIxZySqdfky9lSBdRlxMTrffvaNjHJwhuBshR8u0Uush6xNp25Or5cc9x
AaMsI10sxf+dDGHJov97aXuZLbEGHTlvhvB3O/aWxy1Gfsw8ioBv+eYiu72qkVxk
iGUqBal4R6k6T1c1DVF6hVefrhKt7nYQUXtdgEgzVF/4/cSMun6nHm4imTW5Z330
IdCwgWCZ/f60UWTHZ1O6/BEbP6mv8sroPUfHaXwAVUWZNfjdJcEVZfCwRBFuxC7c
tw+KQpHuDClo316LEBOU2GBPeAPGFuGCbj8s7ubYKnAqFgsiFccEi4iLq5qsXadk
QIXwU0IWWetlSPXlqJ3Wx2MS7nebXdqpC0IGXaFwn8ALFYq8LGmoaZWiaFsSQJzN
w+TSec6UPTgU0htEuVsg09E061c9uHd915YJYu0Z7xlJMTsC8wnc+5OXEHOnPvRT
pf4wDvMPVo3MelA1vyxNVxfZxt838RDZ3rhkTfKahmtz0aDGjFvJTyVorwehvPlY
WXEiB+R0zObDeoosKsbiIK/WXKU4M6XL22QEFS1BR/BUtSNV/5uK2Gep9OkLYL6C
ZhIJ36dRSlH45LIG0AV4qWUsHPG5RpKjkS/ytirIiblkEP+0WXKP3BIlF7gZDE1b
vExd8DJxt09VoQu/sQt24sYAVBQgXY1Ljn7FLRlVHIvRpJB3p9x+BztRBN4iours
hmqIrjGlasql3vEjRZl5qInokLYIF0EgQasePtRQ+tL+PxGxwlrR3OQY2c1yqdoE
dh8/+qnQqzxU4TRFr1zGR45M+dkzIgoV1fMxTSxPfTS8AQ68SNpftYlMmhMXgnHz
Z2oIgh1Yhl8Aafr9GH556dem6/EVzH/fmDLSyEdowWtLj49gcuG3Yh9sc7pjS0+B
R8Aki4YL7F8KhkF4X6i72UohAbBdsH7vMh1iwcXdA7vr6TYL5ztP+8057GcjFg8t
XAyKRORjYj44ibrFacz1rN/92TIL3NgudNwHgyIb0PY7uAGg8sCvNXSstUqJ6Ujx
W3kS2OYEe5FN3IWFKRatZjt0E1IxQWtTUzLDHlrlUoMzN1YvnmkJylVmjrgq3qkc
DXKZHvlo1hP2jWNFzwGGVjMAn6nFfgAjdHM/SzSUnHHHHEMV8VjJp20lbh+LaE7/
US4ZlVfBPCt36Ye4NPs1VoAbwJpwS+G7qcEs5Q5GsuE/NAbvCVLPhimaPD9eB5/+
tgalDEBp1wJ4sdwI9PtPExwAWnch73zs+gU9NvDP1KyDtLxjN9UqIgAC7we07x8j
h+AiPSFyKMgiK3EHaHr/qTOugwncUVznVXQn9h2RiElHk6VvYjVIKMpipAiZl9mv
/P3xA28EVRYkL8S2eUW9QI4BIovOCoV7KcqchB8vKbt43XpqLYrGyt1Ko2UnqeFi
NlWQnQ9KuCfKoHpjQjKDmN9ePRPqp6G9lxizlESryaXifuM6obMGqyeMad18k+T0
QA8mzWpjSF8OhX1TxgkyaIYBf3imq0kh/1PhDhAKCGOqbA0cUEkbe12qyF9xJBmi
Tsq2H8sZmjNmMAiwHndI1JtTW5I+mNRNa2aM8U154Qt83DjTjP3W7vLbREL2lwqY
8m03y2PIyh1q886kZ+rS0xSPCDlnTMCEgjZdG0uiL8yP+vVl5VygQ1vLw9maOAKZ
rMBvB+Ak8dBz1ZMtc3Tb2rogfxo4kLQM5FG6WdcJzFN/8K0xIlIrRvVitYOcF+eA
gbRlq3s1MRwlZlXonZvD28pbLy0QxAciW08DxpO+l0FD9ptbHDfg9QuOtY5lK1Fd
skOgHlba4KWt3ZGw0r+1itMkjaaETc7jFSAeAcrwc/IKCzexIKpDEzTfPOA+6WSg
sHeSsXA3rAGZkbf2NwNGaYK94BbBkV+bCYvKsyhCyrXAmwrHBkJ+LifeO2ExVaKS
YV/qEPqWnA72pWUFTGoYgF41Yr7ZmIVND+qEXabcUDLtTCDYxYSXtQNGFbfdDNz4
QWLvbGcIvZMHnY2L33JIwNQpPWuyeS4W2szTw/EwrfxGLav2dOa3FIzBBZHxVIbX
ZpaV1QEg7MZ6PAd1jUUHXR2WaQ9jOYdsCI+fYGknZpWb1D6UzsStW4oe4tWCh9lm
jznS/C6zyMjoiKXlmoCU/0kIyk9bP0E8K1MhP2kB6k4znAqhGHcShIUCH//Np313
Iefh1IQUusYmS2rLNkZ5yik2/FezZUvi8myNjHnGSdDOOb5c9OvClSOl6P2UM4Hg
41E5/g5OmzBnIYXjRU4cAWp43o+5oFk3ZJJ2QguVsPwexF11P/f5VHbW0f+nRr5G
5PuqftF72I0of3zIGEVAbLz6F7DqPxg3OLpPmQB25LHdSLlzgcsotWbAeeX4bm85
q3YrG0Kjwv/It/x7LCZS91W1eTKRm0HnWBWJHWU0M7l5YENFLFaNfUdv8kBWu4EM
0sadybz9fMliDnoanfGEynGfFCD7RbVf5xW+FKdmODe2Nh56cEeU3/Uxg1XJM2mt
jtz0RCyjTy2IY02hYfWJdoEgcz+zLaCLBLb1dQ0jz0jbT8Y5eFMfA86z89VAzzBC
IjZXp0Mwl+e/tjGS9nAaGocTyuBtG0kYGkZCS7+ZxGsCcthJGF0+E7eXR3mDDQUb
F1WA5yM51u/kVgszDp6UFpxhXCINQ/DosiFcMa3OAeNKHdxfuoLuPrKEENx6JEH2
hMtrsKIRwUApFj5GeOsBq2nQzlTcbR3EEkbF8mZZBbtLej/3wpxxOybD3IkQukRb
tcygW+2/6FGKsZb959dQNZSu/tOgicSr7RzxOAqa2smpQw9NG8ylJvvFMHnibsTN
cNPE6l25cWLZhjco+trZULQtWgxCoUfzkTlQ2Ix02niLQJJ7iCqLu12LjEohyW6i
en/tgc3EMG+EI7jun1r0+a8/8hSu7IcvyeR4olKSpxjve2HbqZvPymoO9i6Zh78c
MbaWHUqemiLzBRUQVtsOZVr5MFB2mhKjuqMdStQHPUEZ9+GQALOFPdm6z+4RT8/0
PKUCEfpHldk1So+A1Wv8sPtgNCm4sXVcuS8o6YsKJ48CqkJF06oxBwAzJveSZfts
VwOb7l1p4kK7/1a5Iqe6m/gsOElBae7xJMIAVWUza9OBVX7vchOwzXeeSOiS7+I2
njuvKnYueC+YLAWinwWid/bGBG336SMnb1rBXlpX3oWtHs0ibNNDyrgEWYmB665Y
/jpQshGqoMp/M9B9GQ4ZgwXIZa7MRVvWqOTDnlcSMh2AQe0mGbcBPZ1JdsH9I29K
J2nZiw5LckctpRyNs1S5Gt2kV+N3ioIz5ycdUGfkS/mwusD7sGZKNueSx8TGrfwi
nYAeslFUGBKvxyKIRHt2P4/UDd0yywUWisdpt741vrI25qW+pmIm+CaW1QulbTMa
nywYi4JIYEbtqP9A3ucwgGy0n/r3KdJx0ogMnikDkYSnz+qEikk9LHKgd1/ML1Jr
7k93fPvK/Xi1BuaX2IpYRPHKf0I1JHVHOuqTNNDRSm19Fa7DX0fcjvLWL7m/jJ+4
G0yLP5yj4R1qWfBB9i80rg5m5q6R+pBpIPtp1JdfHW+scifNl/SrpGeVXed7Ui4L
M8nLCIv9opcAFEU9FQbrBMcBE4KfRWNN90eO7c8x3sW65b+H0cKml2nJvbQfienB
fSzU8H10Ia+L9ToD2YNf4Me1+ZHfkf8uy5kdQsOhKMHrh6EVmJ8IBZQXYlW2a51W
VJdEqvJnka3XQHBkKvGESpaF2ILWeGHAicSQg9sMAbz33sHHdkXm0wwdLrReeH1V
hOBZpBLxbn+T7saAlT3sQICpJb5H4b6BJojxbVQZfa2CP8LGQJr7PwRazOR4bLH1
DscKXx+DmodcWysZC0kAYCiFhNZxzaqpPreplk6UW3852FPkrQPo6dPW9M63DnQ8
Gn/1sKnlgKhOt28gRKcMfRY9/M/QpJ3EnOBa+wc0vCaWREpAHopNuuANnu7CbVRm
X5kltKwXiG1jB6SKcabVPzyYuK7wOvzE6V341sydcrRyFuBjmIvzFgOb4jKTrvhV
qovFNYQkppsgBRjgdTZlmxZ2+srN+vJ5rkKUeISU3gERzIA0r+rbivOSC9kSzG4h
Y7FdaVrvT5ST1ciSR9MLCs96F1AYTxd5x99EGyyAd/HvtPXwyTiKH64EBN0dfH1D
RGbMQyrJAAQpye8rqzMt8ZfSFCAnGqPrBv0fjprsAJWG6y6RXocnkGtkBDdVn/J5
bjr//l2D6ifxh0lU0vxZnFYtmqBDpm9OESPVPQl8gQbWfcxGLT/H+Tq/7Jxjm3nq
xT6T0pjJQGW8YwiidGHV2gmwLbl4dTXYgCfoxhX33lJTkb79DurEWt/y2xexNRS5
1aFLbq/ML91xnwekTlKdXUZ2o6YRbifnZNBt1CPNquhkR1ECyTMLSmrwurftBla2
ckzwyUm3R0cv5YV/4fwZGHf+dOjfzyqjE+JXXzB7m6E1OxwpUnIe8E0aZsFEdlWO
FEwAV3ml8cLpDQ9qEjHSbHWIu4c2uh0wCPJBh5OjZN0y7NRr7aXCZlnVsbbXxE40
9QnMkXqbYp8I2NeSUDBIixXK3uZN3iMkHVII1v6m2kmYAyMyLDUPLpdUQBXIJ+d5
fCQOw5amARovi7V+wk0+YGQ9b1tDUwfB9ybEbgJl2yKYkAyT5rkwAPKN5VmJ/mE+
uJb8522vM2zJ09p2TZtmm85tVLOQkyEGWSagff7MhdFBdlkkr3kAKwF0V8On6QX4
R6HNE3XdidkZPnbmVeI8Ja31i5Xb9d75qqq5DjAt8HWfhpeYJpI+uGZNqQqgtRBB
ELAG7zyTVsJbD50RoRvKR5s3vj6xBJV7FIGZnWCn5/B27iSCEjvAWYhefNDseD87
Nr3mkniV5MvDWqWefAU1qWl7LBfQ/iJtlT23xwouEqakRgPEydBQQJkG63y74/tl
TknKHtNrOuidFCeowe3rASBEsnZ3z61snr10jwfleXVUq2dd6O0AwPvx/k2CCpHJ
Gq2/2j0iqcnf0VgMh+bI5s2Vgojx12+fHOBNOFYEUaoy/qV2SxrtxzLRefHsRgYZ
Nxpiwf+nDRjLXcg5cloVT3aCzbK+kDpF3a82S4BfUs/RlzzoSqPt2Rlr89sHzS1F
ijD65ObJKTxgWE32qzR2eKGihVWroDMFTzxOs6HVSOMRyWnhDB1gKOHyF7FToFK8
oEtu9K3oSmdyhI0SKftaqwWj2pTYycPFIbkcuZh3MdG/argWFBt1pO35IDjHpOoq
yTJRXfoOGPj0fSZ+SeEMRBHHZpoXzfVdAzlX8j9rlN0QDBcYUN1XRxKUXmWzX4Bv
VLufT5c1KIjo1oWSb4EKxKy5RC4GhKYTTYgxqbwRAu5Q7MIitzvES/n1iNL+tM+e
6uwffCHO+Yis7JMJenY1geIOl/QhbmTmIGHTtdxRC5ZJCBWAMQPGIdlkXoWTcuYz
IuoDjOwZ6mdQeWH+2mdVuH1vnieOiBoeP0RP5fy6RnXRVXaiv8HHR3yshRRmvBMY
ncZIxIFwlU2vIrXaCbTvuh8qUC36tM30Nl6QZmSeHVCUI2Sg7HoTW49MD41T6WRb
X6II1hpiCfuk4XY27TQxJJn2U10y7PxpUbPWAyxWhywXHkd/wSZKxllfFs8v5FTu
9Nmd1y6gNNkdCeHcYOSWvP3zJSzXn16mqoPCsNBUe/spvJ+unzvYHZH5wNa1IRtp
++lK45Xc5W4zbORNsXfr+EszzaSC1ZN+c+nP3AcpCF1C8O5A4tgfWranamUbmV6G
tllDZKxUwdoeli0s/7MBto2J4hqe7dj3nEwUilX/KSPNmKR0tWFfk+Pq2joF1XsJ
mNa06/mF77rVO8MXexTgVxxsFqIYbhgYLHk0EJVfekQgYr2dGHjkDhLul5GHHOmv
9Rc3v28uF63dwxpaF0eGfvcrO90enfxNDr6Zc/SxRfhhRU7Us7ySuGXtwAeUVkur
ja6tqbRDJCe7NDIa3N1BjirpCGsZi5TNXdsMAD4M9sXVgrj2i2CO9Nt16fYOjd97
HJucqSqptKVvdbg/0Hjhd/7K5hN1ktdrYp/P2DtFwUPfOCYDa7xeu0Jd3FDx2mDi
+aO3g/zZ53kKFC5Ed76kzKVfiTt1Lkja6JeVIS+JLOt8yWbQ3yCPRUXWbIaqCCY+
ACRj9wyf+Ig/OnzAgPKwLJmjJ1CwighS3OVt7lDKWMLDU032fgZ+SHCgcJFLbb5k
TaoWpGsTEu8quF6TCu3zejiBe5MGBm5bpXGbBhElEmQXBiHepaTkUvfBlvxi+ZYQ
cALnVYSfHOQBWxjtvEL22QH61c6bT/ZcTrX/ak7SzWDk5QjpX4KKGS/3iLX0FPE0
eHLJvb1ZIlZSG4LUK7VxQq5AYnijcHhQHiFqtoV1WQuOS6LNeIHTpr14J+m6qYCc
IsMwVDGlA6HITEP8Ww5abZFQGMpTTqK7stZcW2oObjezUdMTBfWonkgxKWjLLtMo
tWul1OxTkgD7pb0/d7iiF1DLxKEgYUtELMiqm7djYC4BZWoiSz/+f36KreEZ8AXu
w3JWtezvGf/JI9vxwf8kO+CD6Zudz6x8zDYZNWf+XV37fdHJCdTEZSbfJfbvuMCW
4ECiRwxBuc3FwB1eSHiqiF3h5nncOeorH657EcZLwkI3YzI4FVoqxf2e1dHyhggR
TwzqCnK9Xb6NTlcFQDz2XqdZPTB7fSXLmHQ3D30O3mbLw8UBuiz8VFngTN3YkF/W
1yjud734a1RKR3dwz8/xzd4u4+0qicdaZMCEixcWqf6vDdIsmDGO043S139oHiwJ
Psz4ZhlJ2czeHd9VtRNunRWuilpXLXx0arHZ4iOmRi+dBbEstH3ZFIWSWctHC04+
G+NvkaT2B0gCGfa1GVnsfmJDrG9xqzNlqI/p2nHCAgsZP+LS/COkSKrjCnR+OBJ2
6ua4q+m3FWGA4nL4kdzwgxF/6VyNuX0b1vpaFIsKKa9YJpYky7ml4ub7ls74C3cm
7KG6W4sQHHe1eHBR2wl9BxuWrmAbNW0xuwwEVhwPbBkSKZU1xTqbgB92CXYsrIHx
xwtTQNsCQAmxGV1+GbcPYnMo5EWod0CR8KljbhCftze1Wtj/VoiDwYiOTb5ka01G
gJXuqZMRXwlhT8eKe9QCfMZvtkoxUaINQiqTk3F5QgA+zgX6sUlUgJatVzMOwdUO
WVl0WvOAGg3jK4YxLgwbEhHQq2yGrfshvwCb7vxPYo7gCcBZ6O4VuV9271/dBvzZ
RUn30SVi7YTTqTREihph+IsYHp4manZXA3StV4ojvtv91yA6u2xrKXfPnY9/tqdn
Zv5pNUAtqXpmh7AfvbuYe9Ox1ZoK2v94qaTrerAELJxWQ6YuXlGSKNl3mVO5n1+J
W/7/D57DUbTzCoNrCkptHQ6BtAeslg9i0DAYMXHd9HponPwc4Z2uYKTAoBz0qK9K
btEFeSkN/BteZKYjIeAsBfLMBF6VWTUh1mF565YqvQhahnc3ZY0//okAP58zRguw
lfwqyoJZuE7w/Ej21i9ptznchKK4yEicRmwtzTyUEVea6n3QFL4atWdBpPei9gfb
s8zQg9eVqsRovqEpiZUuzayE4n1YTd7bAk+3TTk8udnmRjCp+Pvy9TgSfbbECpP0
bcp0kUtAAXcoqeb/EaxHfez4rWB5NZgZHgEn2STjGXw8bkAp7tv061DiShFxZJtp
mnI+IMpaWe+EUVHvfOuO3WEV269XZVuGzpcse8piDWXI5n7Phc2MBiycSibszFVx
pwIqf8KB8Vd5VWDt7O8f6+XMDO3mn3zu9M8SwKhF2Tbcy5CIqEweFMrplWYHRfYD
y97G443JtGpiKIJ1aqxGJ602xPKDCIUcfnoHxDdsUQBZLB64Uk2foPyJXCt+9UTG
zvszyzocKY5NDXY3gNNeG/KkSzjz9pECzh0hI8uFJ6CDo+sjtrhalim64Qs9jqak
xiE0ryiaiyQLe5FhMWW8JX+yzS20jXbJO9qcH6i/ArsSe5DPn6gdosboT+fG0qJE
te6g6NPWGzNv0AGQ8aYQUx/pJWeEEEx8krfBh7LAiYz7kKfbLPNCjN1tlUWiLH9S
QeLqXfvMHOZWmcoa+iSpnnMPYYC8LIVg4fTlHk/lfHOTpriqVhlWmDXCJz606q4Q
P8ZHB/qkx3cimWbHp/WpCYTnqOZgINZg13FKhWnqpCIlygXp8uZa9go3AUD950v0
sMlNy4UOKslbd9lvk38zcisXthAxzjQ0MEhzJOlFw5vo6JnhicmVTlsM/Vi+5JcW
V1LzVKbh85mAjA0nAl6GaKxlLznmyS2FtnAhvWWFptiXgaqBMP1JZJUknA16fjHa
U30dpsggnBR2WzZ0WqwpoEcgQC7bgao+cjy9P0s1kuDbgHywt83DCMdWuZvBDq6L
j0bfgeaLSODRi/1HLaqxUyt+z8+9sFPYucMJNPA0MWd1a2XPEyaaX6VKH375lM5l
x1zJ1NBtx0+gQVJnGDSEOdZH3jj6w9+jZHPmS+jTHGJgJrOVwIUHIbLSTXC0uWaw
7d16btmm/2MAWotGFBasZetrUI9e03ko89OzcAQ1B6ZOw+3dXZFsdpyMxNOp4axV
Cm2MQ6KYHsMpmaM5EhQ4bdcDd2/fUtpJfx2Lus7vb/+4tm+pQm84ZjCdRiqUA1E8
SGyGKzyj+C3U7rKGcyLjzDKpmgO+fz+anY/PmZqYdByk7xTlkbEBF1kt7fc1u/yG
tKQb5Ekr4wqJYFFsQKefYZPrCrUHB/vtaAbuGydEAKASBliTXCfcVarzUcXY0LxQ
UGPsCaN+3W2jVYzpaknqLznzV/cXujqbEP3zstYRaMzzGMWIqIfqC9h/+ODkmN2H
dcGoXd6knmfTnALMsDhhlHdKo6yIwDhDjzSC/RBui0wogukr33MOn0DpBUsiG/Ja
fqCeGUxP81s6m84iWWXYQqH4AqmokTwrcSDe44VnRz80ZSeXKbI/EKG0WsFxrfsU
pW2P9Ad1Qy8DMtT99A/QkPhGuJhe9T3+Udt8Mwtw8uQFn/DcayujXI7VacuYGk2V
8JthbHvGxE20UqDzQHpywpQD80CXTAQopRzhiNq/kqa2AcqJSzmXCQ+LJZp/FfjL
D5yzSGB0gKaDeFYGupinG6qo8DJywagrUKMQ7pyccpLgZmc+SbqtAWkl/XKdBrQL
i6hyii0h7MqoYM7wlL29Am/cfoHWNyEBWjYyO2uam0Wh9KDrGnebN5tsIdo1brZZ
0Nqe1TaKQTSUTE7NQ4eUzKN2Y86U8MYfuwyILTHmRlSAd7+/gI2EfTI2553oJ6yU
WTwpMg6a3BO7oK2ihpUqHsE59nBhPp4jMz93+VlKSHzN7A8MMAIT3XW9cjywSZaX
yQdKa/yVEFAHuvap18JKRxkYJlrgLevBlzn5ckJdQ4vopFQBlDLn3buHafMZWtX6
IOSaePCDwqElPgNINKUFq+f2jKy2No1vmanPbY/fWa6J4vtykyANAs4uvyK92B3+
2fQeXgNX1KmGyioH/Ur28taJQpv2OZWREmmfV/XAjqnlDu+JBcn7VB7mz17Y/QHr
9J4CXY21aMIHo1yFzo8y6s6oAxZ9f+zenZWTYyPfxW4KQ8h3Wx68NKrhDNZoZIH/
kzmwqnc9bQNC3vot5SjySsPghhIYaM/bSOJmhwZkoNYpeFxhj5NSm5cjnoj/z0on
neixa3m0twwLP4WMTWxoZriy3TYWOg1fiIGS2RUYSyFNS+93mfQVEZFSw4McJJlv
qcCqVLS6Abe1QnvZOyjjJSNLQPaXi4CVuvppaHIpQNZZ4Ul7IKm5PtcJsBd6wZHv
hrrkS32DzGqF3b3/paTA74oCO6GYyx1DYQVOhcqM5Y/WO1jnLQjdP+1Uqy7oxXEE
+x3RLYek0L/wnF0BUnnrdZzhE8a2ali9Txa92U1fsibeFzDYCxP8N215KpeDpQ/u
I0j0LHszLkxUKOReEag3nQVnKLMnxEAsT6FwzxSreBVfpje/rIk60RpQCzGHrD4c
cXbGRf3mlNcwe2xPGw8ZMjhOKKSc7IFbBqRdFavodMIUJS7udrSg29ul0L35zNe1
OAYgWYzZULya3OFEovE9tmUNOqDE9XzWmS5xeQGIKuMBZu7H+D3XksgnHptsH4cZ
CfgrQu7H7r3mAHYaUfmVdlTm7pPmigGiPnr8F3pXRvvpgv1I38LxpBnnPAS3ztG5
q4EFP11ROOof2A2HoDHKt5f1K+Q5rMseOyGg6zUQXS2BirvGOKN7b2vjEGMbFx9C
YsdCzaMW3x9opT3RvdlFL50v7mN8TxiOU05Io4xl91SQX3H71aY5JcjfyLtzgEsB
zGH9ItVpSMoUhc4FEHNSlWvuM1o9dl7JHxmAEO6DCasRGqI2fc9TA7Cud/dtiUcr
/ca02aF/XzJnrWL3TLIHKvlZ3wRGGS0LBwfHWn4fZ5IPpJBLpWDPjh8dthyrjjOE
inziCs4DkShtbuIGj6yjMpBUF5d/vnzwU2MXHZOQ86W1vqtpPUmmUIH0kZxczOLm
ZuHv65NBBpvqSjKpQqE+R0zaZY4XXMG/pR+87qoCfFGxtoi06mxCSHQl4aaancMW
cTr3jeLBqXsi9rLqnhrsW/f1NfNN3ghBAnhFYegaOwgJRxBx2UrB+GwH5q6eFUBj
RwLoQI9Da0inHZcpLZfyTY/W8Kge2YmkIozTfpM2a/yOvWjsmgg5yZNoZvEuIe3U
ATCr3kiAEl2n5889ijaJ+Ki64uBaOm3dkn07DZ629EQfWkgUnA+fKrAnaWmfjDkS
FzS10efkj4QZLW2wbrQednxJW5bol+PjFndYqwPsSNSQMCNMcVy2mmeZebvrGD5g
o5iuXTnV0D4gzz11sCLqPPpVkW3s5eYpUZTo5lbkrfOU5Ty+5TKKX/XUVY1W//Zj
+HcpSKo+XS8Ic5CE5cBP4Dllsi85bZtD/v78ocKT0C+/2kOrSJM2TK7t5BoLw2TB
7e5/CIp0lXnqgFQ+jDJkf/PzIUUUBK+J5kiZdQBZ+ZFG4W6JCDnKkOuU2ooNbwia
iISVxE9WUfp4r2lNP9fwz4i1gYaWnkmbSKtRdCojjF0muqJ/UwizD29h5apjYBKg
hCD6iW23uYDTmgcEHMCpn1i5E08GmPWUBXASUQEUjJHqcV8na70dw87uyea2+JL7
/Eyi5iEzKxcn1ju4dnqbl6K8SgeZOUbvGwX5Xsi2aI0snq796XK6NWaoBQxRkgzF
rzzgWCkQTOt5LGIZWQer6gmRkXcTGnanlHqmJjcGjN4+vykVCvouumAKOCg4wbE4
X9HFiLZFYMOROD86PEujPzmIHW4hy8pg6plheBPKigUGkoSMFxJKBqItUddyAsBs
tlK3spMx0n8Ud1pRnXD221PS2Uu51hBAN5lXKjMIaO3VrHkSg40Z2hM0i/u+IB/y
aQJO0a7KP1xnOF61P9h0OZ0YOfINcYycbvbddum/NqNo2C6sxzr7YDOKC/EC57Eq
ntXgV0VhOBcEaC1tUuYlNVaFG8uhkH02j2398JzzPr+oCoUi7rhrWr4O719rRPLh
WG3ayhauU3NLxFDbainDl/P7RsPeR6yQz7fwPMXsLbugCPJCflSIz5ywotQILVPI
7MVs+UXy31CcO1Er9as5IuC6QUFgrMz68DjHlnGZTBN4+AvsC2ZtSTZtVA525wqt
GzCGHFW//bpo1w+2vx4s/z/ozzx2Q+a/wZwURcMIhN0Vds0vsXfDb43DvKGwyD72
8J7bnA/SQ4r0GGQFI1aUSdmBpaL3jzd5BtP4+9HevaksPZ6u/Bb/3G1qyp6TCXrx
WV2/wMAfOxnyNhCxsf8yZhZe/8J913usB73V1OREoR5BpEt0wE0a8Y3x9Qkvaf9w
rJMwuJjgyGhk0x2TReaZaWRebT/Eh5iYuqCVd/SUixUXtOKCT7QvaS+WkS+bBtC3
vRDECzkd/XPiAtwj4Rqo7+2BbsWj8lRk5Sce6bOXJI8xS3eKscxv5MRkXRNpIscW
H0DmQ1R2gj3vhEcvXhBIIVJwOAbp37nSI+nlaqakdD4deffOjmZNNyGCKpY4/cdM
OpYeR4hMIbKIQtPnNq07DgfX2uHXthujLe7+uPWed+Zdalf4ZANGEKbIDl3+tpB+
eIbWtlRk1yOlwJhuq8GfTKZL4uOoJz2GTLA1dTU8ayM/yOt8zoqeGNtP6oIow5l9
PXZVbJf6O4QU58FQ5YCQHaPiQ9tPjQ9GFD42v4s0j7EPtuDPTtPUCT0L4aV/jU/4
MFoubFJEzhqgaiJkeS/vClZ/q+aj3B0bVrFAG4lIiJGPlaZ+bpiwFgcbgU0kyYbd
n8Na0K8jNwVYv1V4akRDWlHwc+0xtA4bAyeuHocnPnsQbcdNIowC8HQYtAJ5rsf1
aYqjltpAhCS1MpoUlg14BVlBZXNEh3seG4c6EQpvKg4d4P8hHaMy/GGsYtlGuopk
c1ICHTLDaWI0jYxwauHrhscrVw6smZ/i84YmjTPo5J1r1pQ2C1/Z66ZRJkwF9E4u
O4+LDE6EL59Z1bWqyJwoTR9QDXfUOfsGU3HnX5Nr4KFUQfHALB3hcCa0VeLQsGhd
2PWyRk7LUqsYZIW8TgSQjzZu9SCng7ajJLsGD/auLjJRY4STSIhFuYF6lMWA6zsz
mx+K/cynk+3KedxFhjNZJ3FvwrGiSabmvbyHaZH29DmuqmvSubD1onP/d3p4VKeS
mFTFdExiPrv+Yo+yXw2cwzcyBKDPtQOYERQP2m3LpCSc/VHv4r9/L0TuodaWRxCK
7oNl8ty4kI7u/uVFncu9fkQXw8XsLD7vo5O5bn7DPl1QqLCv+ZpwkxdysSdAQ9mm
ClppbvCjtmXUxEozmA/+EOeHYdh3xQTHtbXqNX6CfOWSWssmsWOGGBC5hObmYHNd
nKML78vLhvz9/NhdQFx3MWBKHeoSRWh+I20QI2wgC/JMliOClygikUfW/s7Pbn/6
iEk+5CX4SvaW7FG1pscJ+9SykJ5Rz/iwDmSrpNPZh/end2nXgRKzyHnbCTocQpz0
14agxJUu2lAL2yZZpqLDoDoeIiS7PUCnUBjm2+7zHfhRoLlC4UF3S2RghHnUqVlW
BH9sx2kCEgtAJOqE7EB7ZzCffU75U7t1s0/WK7lcfQatgaLi09wTo9GQf8MF0gPv
q5DlE8vZSb5MvZyZKmRCyvxSMvaKRD/9B/6+8jAc/2WvDYdQdCcnUNYgJq1oMP1L
+gvrilzTIZGVx6cZm7UUt9QSVqZ4taWkHUJN1yisOxpJQZ7K6b2V+jyS5u2MPnsn
EE0xIBzUXHGsieT8uQyrWXIML09yxIJqFycIBlC6xdfIvFO1oqwCscvWV5u7+wP/
H80uwqIXtqcCXtjHtjrdbse3GXSljqhVfi729Tl5WO2jx2ADee4cC0TJPuIQv06n
2sInHeMEIUvaLjzBqpHV8ttm8rFGh8i0LZ9k1tB8k4bvCPBzFG+YvlNyUGRMWkxP

//pragma protect end_data_block
//pragma protect digest_block
lNed3KW8TCjC0o5WYFD2+prr9VE=
//pragma protect end_digest_block
//pragma protect end_protected

`endif










