
`ifndef GUARD_SVT_AXI_PORT_MONITOR_PA_WRITER_CALLBACKS_SV
`define GUARD_SVT_AXI_PORT_MONITOR_PA_WRITER_CALLBACKS_SV

// =====================================================================================================================
/**
* The svt_axi_port_monitor_pa_writer_callbacks class is extended from the
* #svt_axi_port_monitor_callback class in order to write out protocol object 
* information (using the svt_xml_writer class).
  */
 class svt_axi_port_monitor_pa_writer_callbacks extends svt_axi_port_monitor_callback;

 // ****************************************************************************
 // Data
 // ****************************************************************************


 /** Writer used to generate PA output for transactions. */
 protected svt_xml_writer xml_writer = null;

 // The following are required for storing start and end timing info of the transaction.
 protected real xact_start_time =0;
 protected real xact_end_time =0; 
 string channel;
 protected real write_address_phase_start_time = 0;
 protected real write_address_phase_end_time = 0;
 protected real write_data_phase_start_time = 0;
 protected real write_data_phase_end_time = 0;
 protected real read_address_phase_start_time = 0;
 protected real read_address_phase_end_time = 0;
 protected real read_data_phase_start_time = 0;
 protected real read_data_phase_end_time = 0;
 protected real write_resp_phase_start_time = 0;
 protected real write_resp_phase_end_time = 0;
 protected real snoop_resp_phase_end_time = 0;
 protected real snoop_data_phase_end_time = 0;
 protected real snoop_address_phase_end_time = 0;
 protected real snoop_resp_phase_start_time = 0;
 protected real snoop_data_phase_start_time = 0;
 protected real snoop_address_phase_start_time = 0;
 protected real stream_transfer_start_time = 0;
 protected real stream_transfer_end_time = 0;
 protected real snoop_xact_start_time =0;
 protected real snoop_xact_end_time ;
 
 // These arrays are used to check or associate each started callback  with the ended callback
 protected bit  xact_started_cb[svt_axi_transaction];
 protected bit snoop_xact_started_cb[svt_axi_snoop_transaction];
 protected bit  write_addr_phase_cb[svt_axi_transaction];
 protected bit  read_addr_phase_cb[svt_axi_transaction];
 protected bit  write_resp_phase_cb[svt_axi_transaction];
 protected bit  snoop_addr_phase_cb[svt_axi_snoop_transaction];
 protected bit  snoop_resp_phase_cb[svt_axi_snoop_transaction];
 protected bit stream_xact_started_cb[svt_axi_transaction];
 protected bit [7:0] write_data_phase_cb[svt_axi_transaction];
 protected bit [7:0] read_data_phase_cb[svt_axi_transaction];
 protected bit [7:0] snoop_data_phase_cb[svt_axi_snoop_transaction];
 
 //string to store the parent child relationship of transactions
 string parent_uid, transaction_uid;

 //string to store the object_type of string
 string object_type ;

 //counter to count the no ace_bus_data object type 
 int pa_start_count =0;
 int end_count =0;

 // ****************************************************************************
 // Methods
 // ****************************************************************************

 //----------------------------------------------------------------------------
 /** CONSTRUCTOR: Create a new callback instance */
 `ifdef SVT_VMM_TECHNOLOGY
   extern function new(svt_xml_writer xml_writer);
 `else
   extern function new(svt_xml_writer xml_writer,string name = "svt_axi_port_monitor_pa_writer_callbacks");
 `endif

 //----------------------------------------------------------------------------

 /** Called when a new transaction is observed on the port */
 extern virtual function void new_transaction_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);

 /** Called when a transaction ends */
 extern  virtual function void transaction_ended(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);


 /** Called before putting a snoop transaction to the analysis port */
 extern  virtual function void pre_snoop_output_port_put(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);


 /** Called when a new snoop transaction is observed on the port */
 extern   virtual function void new_snoop_transaction_started(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);


 /** Called when ACVALID is asserted */
 extern   virtual function void snoop_address_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);


 /** Called when snoop address handshake is complete, that is, when ACVALID 
 * and ACREADY are asserted */
extern  virtual function void snoop_address_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);


/** Called when CDVALID is asserted */
extern virtual function void snoop_data_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);


/** Called when snoop data handshake is complete, that is, when CDVALID 
* and CDREADY are asserted */
  extern virtual function void snoop_data_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);


  /** Called when CRVALID is asserted */
  extern   virtual function void snoop_resp_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);


  /** Called when snoop response handshake is complete, that is, when CRVALID 
  * and CRREADY are asserted */
 extern   virtual function void snoop_resp_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);


 /** Called when AWVALID is asserted */
 extern  virtual function void write_address_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);

 /** 
 * Called when write address handshake is complete, that is, when AWVALID 
 * and AWREADY are asserted. Extension of this method in the default coverage 
 * callback class is used for signal coverage of write address channel signals.
   */
  extern   virtual function void write_address_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);


  /** Called when ARVALID is asserted */
  extern  virtual function void read_address_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);


  /** 
  * Called when read address handshake is complete, that is, when ARVALID 
  * and ARREADY are asserted. Extension of this method in the default coverage 
  * callback class is used for signal coverage of read address channel signals.
    */
   extern   virtual function void read_address_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);


   /** Called when WVALID is asserted */
   extern virtual function void write_data_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);


   /** 
   * Called when write data handshake is complete, that is, when WVALID 
   * and WREADY are asserted. Extension of this method in the default coverage 
   * callback class is used for signal coverage of write data channel signals.
     */ 
    extern  virtual function void write_data_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);


    /** Called when RVALID is asserted */
    extern  virtual function void read_data_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);


    /** 
    * Called when read data handshake is complete, that is, when RVALID 
    * and RREADY are asserted. Extension of this method in the default coverage 
    * callback class is used for signal coverage of read data channel signals.
      */ 
     extern  virtual function void read_data_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);

     /** Called when BVALID is asserted */
     extern   virtual function void write_resp_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);


     /** 
     * Called when write response handshake is complete, that is, when BVALID 
     * and BREADY are asserted. Extension of this method in the default coverage 
     * callback class is used for signal coverage of write response channel signals.
       */
      extern   virtual function void write_resp_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);


      /** Called when TVALID is asserted */
      extern virtual function void stream_transfer_started(svt_axi_port_monitor axi_monitor,svt_axi_transaction item);


      /** Called when stream handshake is complete, that is, when TVALID and TREADY are asserted */
      extern virtual  function void stream_transfer_ended(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);

      //==================================================================================
      `ifndef SVT_VMM_TECHNOLOGY
      /** Returns this class name as a string. */
      virtual function string get_type_name();
      get_type_name = "svt_axi_port_monitor_pa_writer_callbacks";
    endfunction  
  `endif

  endclass : svt_axi_port_monitor_pa_writer_callbacks

  //================================================================================

  `protected
-b5#A424ZCc2)\CL?KYJQ^,>1H=^,3IA=(5X+0DW\PJW4d(6AXIP+)?HUga9QIW<
R1V8,3e_bO.HK:/#?P6R>[U8YD#,:g9K_/U.55IO=<(LR>Eg1Q+V0W=PTN&OR1I(
FAE9BSA^dGGDG1SS+EH^cOMZd0BH;<=g92J\\e;A@79R[\&+Q)WYga<B2,gTHg3T
5[@_^FF=(+d2c+L<0LWTOS&Q2ZggB_#1.=^SFF[R/@[C,]C/.#32L,d2GcY6QOaX
G)63L]^2+<A(6Q#T1Xb<f^^X,\+6F6;&+9<=fRI3;GT[L3Ac_G/>A#BG-+;,Qe-B
]d4:H/[bgXa(LC^Z6E&TK]Fa)H0;^2P8;,?CI@AHbdV3HC#/PSae4Y,4[NZ1VSL)
R?>#GXbQ=>_U-5]Q)M-a-(:2=?W&_>5V;T&VO7MTMDV?HTBE0TKR^^-8S-C)WI@?
QALgHZ99DU5B=NLeCbBU-U:#;#W=B6Y/)C6Yea5P[f@IFH5UXY\+WdE5I#46IMJf
f9g#fUXYeD?4Y[dY5Y:,gNN6K8&.d?-)E<?EWGHg6.B#3;?V:Z/#HJ@DODJU<D7?
cQGE.__KHc@++_/aYG(U\XZ(N+-fNcSYV+>?9)XEUGe.8KGGR=/8#I7M7LBN2R4e
e2Mc:fZ[X7G&M4@K_633f^&IC)6@_R+\6I9ULE:9[d/F.+6a2.L#B@MVSVa<P7.7
)R?\d+;.3R/d7X\YWa)/DG)ETgN\)Z/AL&Z(fM<7Z=:2U=80d[-2UW.4N(G^aT0P
RVgV-81A77_g&581_2:I@L75Jc_5J,XEEMN2U,f9ffZMY/bJ6T306#/VOVF4b8XD
>NE12:4_L>1DR5JS2221cW2C]>F-]36GZESZ.F0Ig<G_<.UYbWD\)bF>dgQU2F0Z
L?b_?;T8SPIW,Y0UbOe+.MT-cG=3Va[#NGf(N+b\E#:d5Vf0ZB))M))^Pb+\1G:F
^2JWK;HI,(f&QT>e-OJc;TN+4X+V#VRd2-DNd88DME4<GKcRP8\T;B=;+Z-GU2K9
8A>,I)BW;O\a-BV2dMP&PFB4\T?2EHB<MY43/c7B9G(,^HG1e9TT35==CJDX/W[>
]SLJ\Ma+--T/.NMHC2RL#HW[b_/Ld2NR8HW:>]WMcGf8fVf)JN#KO?RU[1eDd@B@
\gKC>M?#P7GO;CK+[O]JKfZ=+OH^gCPH#+[+@=e<)L1ZD#EQA[DFbAZZ2.5]\9WP
@09[?;O3T5.;/J+F)G4B63W&H44Kg80cV[D7d-^#QW/\O)PH[?\3\QHV.[9.0AWG
W;9C_94-[aUOc>I,P3Sf,6)62VD]@@F:3:VR1VbH6>3XA\9,g=:e72-SLY/;J+M5
fW4B8BHVa/KYX[=&7;3W?RB[QEMZ0V1.BOcW^_(2ADKH6b=bULU/IX\DKYX#]gf<
K>Kd/>)-g_P4>\=AJB[-[VJ3JDdN)KIee.gL,N@3]APPJC5YDW8(eOHL?)Cg#<P]
2c+[I^O-2,^WYD...RHX.8V<JI6SI=]NKQdLgcT)]YTZ8WJDT-adV&G-2SVFG40W
O;G6I&2TK]\GO#ZFQa<Yb?GS\A^XJ[[EN5B/9&8XK;DX[1@PY]6US=aY&2c<Vf5O
B\I/Q.VOXAUOZDS57,O^F824\@b^FO;+U4_1PEeHGVRM:#GK2-QC>Jf4)UI-Xbb5
]F9Q^e:aJ)#;Yd<S/a7-6(cEJ:9BKCG_IOHc>cZCHEgZI^Z2+07&cDcbMWJ3ZE#G
cY,QXVQBI#7TAV?0G#IVd/gfND[X/3G((YR&SQ=#AV:cg:I#DF7UFP\-EZ;HL9_Y
>.@fd\#U0^WKFDd^/7e2@5Ob=K0aC[QM^=6H^-]Z#b?XbSaF<_<LO0?WE-033\AW
&c.@4=a3)G<[dQTCXUEN<).aXI-g7?)X2;>&Ne&1DJ5Ng@Q:W577F4?C,fLWT_/E
8ebRf_LB>Z<,D4KI,YgHV[fGVRLddW9g77Z+(dadO2ZaN)bAMZeA:0\,98/NXfW^
Rdfe3)T>P&)&I\7B&fKK40V225eb_,02D9T>5@:Z:1=MEd+/I:3MHYW=\^EUc]<1
;dP).4J(BdE^,f:S-ID9LZMZ6g[TS2@a]]b87Gc6d54+\F;B\FfA\]M,CW76MZAE
e3L</gCNB1aK+X\Q4,-F[LU_DXdBa&6<C>16cM0+0C3;\9B,FIOX)+0UII?KRW9Q
+&^.A^d,B?S,^3R]B9Xg-Z8[Y&?D0EgF7,YY=P#dcTQU7X:9faDHLU/58g?.3;/>
-/)2/b]+R5UdGKDV/X,M.SXDOJ2.V(cO94PJa4>2<_RS<K;<ALeDG/+;[SE#5A:4
D_[-2C4IG[Xgg5-IYVUe=MV-845)PMQV:BPKA:>E/1+#;A5B>^9]@ABG(^5./cH;
:\W2A]@K\R2[,;@+MOP,J>YId<cX2_:5aef17c@a]JXBO;CbcCMa&:gKaX@dKe<\
DN<1@?#D2U2XRb..,ODF4BS#Q[\CDd7;EGPS_YF\,7LG#?f(fS548L?P89RN)L?E
4?I3)Nb0DZ8c2>Fea2N>KT/gOI-?OZX;?U+BXMO)Cb83-BM;V0bYGccTQ0K?b#[e
@=OE=b,GI0J9f6>=\B7ESRa.@#8gZ/U(Pg@LQbZ^.9B_?HQ+/O.XMbf#CD95I&2I
gJTIZX4Ub3^C[2f_=Ne(D@gG6YG-P8./fC^9<3_5TJIG-fW)9,F9Ig1J)De9PIS]
?[Sa2AO<(cHD1#:HJGW6[G#U\KbC+3MaDS4YY),1Q6L1.Ng6gD;MZ@G:_365-cb?
\MOdf0JWDF#T?K[EGS#.L<0JG02D:.KHQXTJC,VfY]:EUNdURP7++KdIMO4e\SU2
:CGK_.J,c+f=.?U=/,]aG?&R;YH^01+[7^=ZH/_Od9O^E5]&Aa]&:90>(5BU^eF(
3g?X2:PEL3bUgb8C?,XSN(=Z0GFZ2;6U7#e/Lf/_C_GL:fA9;(1VZ?g2_7_D,(=G
R-CPU08U,8g+fPHKI@O4X1U_9\>A/,dVBTcf.UB)aJOXULGYB)OFNL4-.8eWE>&0
NT0>WFTE#2/C7]bdV2W\4(_7B<>gXI\T:/^X^(?.A\A0CHH,W34&7<(DQ2]Y+X.#
ed>MVOAY?YSJJI2?3WK_Q-F]FCgC78EB:BA3VQ@:;VI?@@dLATAYb>MU^fTL?9:^
S-D:5G(I]cZ#EA.<ZXRY4NIPGTQW\ZFL2.8POGAeYXMO)-(324/JfJSR/\4f+BJY
MU,#EXV?Xa8]8KUCdeeT>&UT/b0a>[e?.S,J>9e)BRcbS/G(,C?BO&@(_bP6I/RP
57UCTF(g>]U&,:E27^N_a3#3PeN>7dW,+K)ZDg-f(LIS9[3E)#N:RPc(Y-0K(5;V
2?EbZQN<.Y2++gd826_C68]4F\,HH&\A#d)9L(2\B+>S[D#UIfQ^bE^=08?KLC&=
(9+<4&VOI#EIY0UgX+XU4-S@&\gPd6TX:(9,Z@Z-f1cX70G+28WW6;;^.8Vc@.@a
X\(2+dQ&fN+C(O47(,.T>RRaEK<-dPf<H)NVc]D^[1dI;V,8[fg3J[W+b6baEL?=
II,UZ/Mc+)T4aTTV(;(@Hb=A0g[3AQ+L>?;J7?9[K-3@c-OIJ?M.;KIZ2<U0A9a7
5QD-8HJ?Y.R=Ie=O)d\84GIT\^PJ=c^+#<)Z=1gb8gc<(Le5e?<5cVY_+EL3H]OX
O[JO][,]EY#6&(E0]-dH#\8C&bC5G;S\6_U9EU[UE=faWNTNC8]cg_FW\Z(2)N2@
)[FJA3,G1(I6S\f64F8d,QM,c?]ZdfIVH/45\M_cJ&85F_Z=PR0ICF4V^GBI.O0Y
SREA)dRH&8I=?SZaAQb(\.:#(eN@<a5@d;YGR9CQZ;HCXSU4f:O]4OTUUCe4^O:N
2][0ff>;N5b@-RZ/,gBDL>AMC>/AN>+DXZQ7Pf?S2fgX@?M_NS.,K+T2<QC7-?=&
8Ude/SPALUUV-b;\BOKC84]8254W(JX]bBb2SXVH<MY7Z3)R#(UX3D]AGWH#PQ;L
+[T<9M1b,:.5>TBLE-6PSH<J@6L79dR5][U7\-E4&7.bG-N;gF-T#7>fO#BeJPJ]
bZ(C5L36BA5V,I8XX-EZ/Z5>H=DgT<BO;Gd#7M8OFW+^H4#H6.<Wec7U;-Z_VLbV
^]UQZ<f>[U.G\\NBCSJZ=LTCc[G0#7dA2c0B-C5O)G1_T1,gHXZ_3]UdH@YU[808
UTPcR[I[Tg.5?I^,3X\>B?)Ad=(1P<IZDHAQG(YOX47gfX20#IFEO#8a8#-H<NKc
Jg/NO]1,G&M+;,HVg&)gF01D>4O]aAc];C&OV:4JRa;>EfJ)eOI@\VF(TL5C6MP7
?+5AB4ZP0Wa;1:TQZUUYX3:39[\I;UfKR,B<ZZ9=0U-C4/M0/-_Bae77a1dage2N
;2YPY8+NX;)PL.KY3SQf3K(]dd=dHdQLY9_D18=6HMN6gCK#dS5IfP\>b-5IbXV&
?_(U1]<Y6EdWM6eW0Xf6&@#.#.=JLeH,U#eM&AF2#fI/RO#ada&>^-d)XS[Ad_@_
CB.JB.U8(YH\[)/RBAT4?+UL/]7W:DS6SW31RKB+WYD]Ae^GU1X,L4Y9W9?>;fF<
T,?L)&__J#/50bL^_NLI^0N>Lg>>?C+>PV71]ZB]:g[d()\g=gR@A0CPD@_[RbY9
,D@+eP@4+@FC56]/C:UdfLGS#eW:P\Ga>-e=Gf9TWIcN\>>Pa&dVGCS+AC>;5\c:
-U@e[d7@db3OZ)MaS08@6.1WT+/VZ]b9/F-Y5S\/K<9^)VXX]=F_/;]MMR=Bg8JY
.+PFYb,Ke];?D7SaA/>)7cCV045,WXd:[32VVOE>9feD/EV[RS0/)[;UaW#4CX^L
eGC#^Y_@bHO;AVEG^@>-5]EFMK>T(g2P1@/TY+TY/YT9HTJMS/EUU,]G//61<Ld4
87F/BC;Q=I=0_&WC9^05>AZS6,fDJ4R-UA80??dS,#LLFQ-Cd[fU0Ia.+QND9d&D
#.=U<QXUC8C2JUAbDe]aWEP3K:2B0b/^84L7e9B:>IX\).Ua(:T4C?[)SLE2XI7?
#K2K.g5O>W2TB_bY&U:,#O//1V&4F9W/?8fK2]QDZI4MNW.(f#</(+R,23K0:/IK
Q6HN#U;e.c;0)6T5[FgdIaQ@C;4I;JYR@L668-)BUIEZg&.6:>QgJ@6&06&)J57P
6R@9ObX(]>S?_g^OV08D?aA1\e<\B/&BJA8IaHI:0E\;_)@;43CKB3c3-++W]b1,
RFQU[5Ue.Q,a_:;L-&XDC,gC,=e2d(E>8Y]+Q\bg[\f](ET=TK0IRF=>+6OJM@ea
3V;]Lf5R=ZM[O<\(T5PbL.VX#9/SX/CJ+VeaK1Q(Z4WEM\Ma700ad6Cf.E>?J8WE
<OVCQO]P7&BJ1X=/F0VaS(d.&_P1>]HT)L8+S/7PT&/-e)<4d]YG21V[,I2I>ZG9
.MYU\?#AI1D1\eC^3-[CFE>ST;DK.9a84c[3T<,RDG\];Id)H:K(MHC-&Ra\&@-1
Q&S/7NEFEL\WXLDAR]896Ia?(IYWS)MKZIEbQdfXbB[^bI;+N-\VJ.SCRKL-I?2G
2JeLB.^TV6c_B5FSI.[4WgTLf60e_HC4Ga6&,<(WM]Ga(g/,,,P&Y8KaB:?H;?EY
)-.@=ZQ>@]bdT1#e^BQ:&#[WX,.>^/E\FcSR6@R,8]?\6dA<=A[9/M1]EE#[#9;&
]-/#HJf_eX3@]f8)c9[WYDLCbKYQ\&d9MYZ#aN^AX-H<_,:5(f=b15(Q#GU17TYR
=fP@S13;<aB>F9MJ/8NO<,g5CR^=]d;W?B6RZXM_N/50eI\.@OT/)WN3\caaL:3\
&V76a1=CV/9M,^(&:YMFCKA+)7DEKQ09f&FDeL5/bV:c5VU0=:@_;K47:75H^>[=
.?14b&X_(.cSXAO>OO+[R-+cdO733)1bF#[cR>K3RU2\/b+(PIg_;),Vf\YSU+3Q
IQ:IbL@[KIAb:<Df^>D0bJS,+V33B=\AEGQGIY-?MK_Ze9f4(-4fK65@aG[><;[.
dbTA;57_-f-Pe2I[H&@eS5PKN_[[YJZ6&4U6>@_SEX8FG/FE]KFA3H3[+V_f]8UR
ADEQ;V5fD8>;c</+d.2,Df4W/RS=&eA;4GE+X<]e43bEP78?H0RI>.f<0LbdB[&A
U:;2WQb0S=19,=cE3M&?>#edbD;ZdLX.bA=]2SeLV,+P>5B9OdVB[O)M@LN-9C:2
CPGg^M@;27,96T(?O+HeG7RWAWGK)EZ59XEDSHGT;aZH#R_B4.Wf4HQcZYYYH_8@
3f(.J9\YW;a/eU(@9>PK1BU5>;Q>.VT,VbUO3;8OeBXc)_8E(@;ffB7ZA7g=7)H,
P__><\^aL5KcRZ:#WO_c2@b090V0.K+dUARMJ8g@FTc/[BbR793TS9#4;WT]2-JC
g\903N7MA;LC#&KOc?UXTBH_X?ZINIaQd/QY7/83c9A1SIQ:U_<KGedCgc;,WPd5
JX9beMZgK.M2LN#5E]G8d9377(00U:e+ZU(J+_&IZ:Z#F)^EHRg\Ia[M0\L\^J2Y
5BOORX8bVBFQKCeK(NMW/K>N[IdJg;H9)7J&T53cb;?,RA.>AD&T?/b@,<F^;-:a
@[6d6G#VC@Z7aDKCd+^Q21<>/(XTX.[69)d^TSS;:T??_?&\Ie5442ZY.Oa0G1ZZ
5F<L#>4::U8^G.M;AHV6[S@QC>WF.7+736;JU@9)aMYYX/5QfLB,9EQH/[8KcV14
[B>fOfCRKOJ\6ZEO[R-X;;6V_c=O6\@;UQ<PK.N1_@5R:<2+J/H1:+c,-@?R<WU9
IH+0GS-_ZbI/)g@f6D@6/E3OT0c)W9EF^YZBc1d@DD^;+RE3371R>abIYCfZ,E;T
5IdT0KU8,0LKU32.1=(1\/TV#d9X3=N68]CY=;EF9gOa2XHSJ4]]:MaQJ2=;=;2_
CON^Ba4_.PPC2T&G^702dN08K_FQQEIZ=>(g:eFd.T1.Wg9B::&<TA\TZ74Zg>X4
1?5.JNV>ZaC4>7749CT8)E/5<,1.7C+c/S,7Ee65<[WP785=UDYH/135JPecVX5?
A[Z#Y=c7=dMLISC7Q04-D7LM@]C^169U)E(U?N=/NLYMB5T1/QMT]\DB^NJ?dB:D
Rc5-bIR[45#I#F(ZDb3<A#8FM/fg;O,MDS;ATg^F24#@JbZb][e2RPG<M3gXDZO-
(1@G&fb2]X-4[Z[3>/g=X@]LRbH]S]MPd<gg;Dd6,A8f0#V1a/JGbdd&UDL7XGM5
BF;=&]184HXegCXN_9UYH7&=P0_J]:R6/QY.QGDG.H<+;[)]=_=db^6=(_XW>[XB
^W4OP\\N9M&L:PV6S-/Q&WeUU,@+S)(\T_([bYBD4AP+A@#\GPUVJ;#N)P822++(
J/3JK(_MgWZ+\g?Q3BeQc:a?<E:=]YPNbOL+G8dEIdX,6EL3^C=Z=CaQ9\,OJQZ>
2g^B\W@b7Q:KDRB;/FEN[GX:VP3:Mc=f(J1RMeU.UW.2MN4VDN5SI8E?@OE7.QH/
^LWEM8@_WSO@3<dK2SAR-2bHCdJ9Y\Y:=a[A7(PS3DOgH1E\@JIYeZ-:<;a7a4Z6
4M@^<3>Q[;+9\\-G10<+_1VLOUZ-.W<-9.S\O)_R&&5d(3B\BM:J;(HX8/.3\;bd
)3U/JI3Z:<Q(W+ZEJKMf&#I0:W>7YVFH2a/V=f+SO6>g_#EaAF9[D(>Ig4]VVdUP
-P6E5S:L+ALE\9GU(:7S>FMdJK:A:-d?&GgHS/GWdedJ)RT[-99g1bBYBA:g^.?V
a6)6Id)(DGD_cd3QE673Xd+.J3g>A^F\A4LBN+^8=+ZQJ.bWG898L>De^<;c\VY_
00^;2E86AO&36<BW8S>N##MKB)-.e;UH)LSCLNIMR(H^LQ-R]J9E#cN8f4^3:?S2
LId&2GA0:]I2b\OA>O(&(\O(^D6e\eSRe.D1Of2<;T9cN:E()6SI#O-R#V(Z?:=/
YD-;G9?4/,Eff1e_XaZSB)V][:a-#C@99U;f04S5TJ&.?B-f+S^SF:BK.6d/CG=7
(73CYAN+M;[1&02LXcL+Z^549L1NZ1J5[4977+4ACXKQY/5+Q[N3O;Q+<#.&OWE8
1OXJ>4JTMD(-8>TSH_[fP?N9cR_V<V_g4(3WD)9SeU_MJNQf6_=R)/Gc/IX&/W/+
TR@H7SF;82B.,DYWX_cV0=cS,VaK?]AG7Ecc.:[1DS>+G-A(5g1(_.,aY;C(-X[9
>YTI-_B4;])WId)7EfN&XaD?QPDA-X108.#JQd(2U,]5D5<.fRMP9;E4-S_,?0E?
)R?3a@]f/CA;+(gV:-UQBT:&.HI?6E(W=_\:eI7NXKZ:.=^g&+;Ve]\7=0MIQ.7[
&TgN4^>.,=&=-dB](AaMHc+JDLgDZPEO^BV1^F.78_D<9g/Se+=b?O9F3\Q<XOWX
Ld#db_e;R,6MXaYH:&c6,_dY15d)\<JXTT#RWe9/;2:J<.-feES(6>HU#4?=5Ag)
>.-UJB-(JETANRGa0-:X>R4GFA0a17eX(Ve:U+3B:RPHS=WC#R4OTFM5(3HK+X.b
>(9dP<.YOF13+g[0W?c33bZc&()2F,27TG5K5--SQ&B4A,_@G-X9I\,)9,_S^RcG
0]FbK?f#Y-]90SQ:283+KO,DM7<VG0[+_=b00,<&.6@IGZYeGBcD2,ID57F&GEK8
NYc0(/A[GCb>6R4U9H.MQHR)e(UEcS:0c5=0>JGZHC:0[=V0<\1eg9?2S4^_\NeA
G;Y\=J3U62=8/N<&49PY8ABUHAJcH4J]/;<L^.<K0T6@bV.E;IFJM1T=2^GT[V3R
IFV)=fK^)Mf7#S2G38J1E65J=181+bNSEG),7[UG1ZZK-RPC4DgSLRWBMN;:Y+IY
=SeL3gM&I\Qa:<6<_)1c&8?HUFPe#JD4@A&=RKT0g]#3ZfSYWMBbZ==-WIc,9LBc
#A&_0QY\H#ReRO&VY6+8G]]+M+/2><KFA2b3.4=>E=Ka^f:IYaGP_Q44K]1/UNL8
JSI(?fF_I]=(E[=A-E42bZb2RJS:97;V7#@MG_^4;7/[^06(-5?<UR34NZMD8A2(
9WLcJX3@F;9bIR<U\fAb_EDXT35dN2TQRNMfQBbCNR8?A]);^SMARN,N1[=)>/C)
PG3b(eM0+O&<7_b9+I#g(fG8M_LE4eJ)^EH.6Ia4(:<70?E3GT4SH_[14ZAH[D<:
UJPg3bD9J2K_MV),87>34/9XAMX_SJ&:Hf\.b\/L6:X7PaNY@SH4a8M\;74^1J61
S8[>W^4F5EMXD\XfFFHaIO1a;UE<-F>I7@O;^E98W9Zg2e9aJ5Id81&d=6>//+I(
N8@ebc;LcFbgag4+SdM5,I_Mf8b;NE>_M2W<W/@2H^b(Z>581<a\#U=4BdT<@<SP
_[\>K^KSgd>W^E#U94^g&E1K3\N)2a(b:MC83>_)bE\LV.0(+;_J12AFYa,C^Q5d
BX.e2&B9[T9_W?6c]f8JZWB8[)9M,D=VS+eJ7;&QCX1[-7c>M2DJ+/1U)#R[21F2
LR&X5NRa[geP28aeQI(N7beQR(KZ\3CM&.BBDeKABO5P,#CW+W>FaB1Y8eP5CV./
0df3D1T<I?B0JgASbeUA@&CHeSV+e@H@B@XYYP+.#=?aFZH_JdG;EXQ6B&aC71;^
KIAKfg#6-R72>@_S^<W9Uc#]<8cGgc\AM_8[K[W4K)JR\:94ZA2\?c5W^3Q<5ST^
Db^65KLfUG6@&b0TO4372/bgW6H_BLg5RF?AHZLCMML3[a49_)1eL^8?/IP]2369
4GPf=VD1BG#IOATVLLGKcEO2ME7QD&^8d\P<c-0A7>1UVLb:aLBTdC1a05,27d7H
Z<LANXQdK#3;>/T6FOXL9)-YC;Z46][,=<b<4Z__8B8/Z+)[WR+,dIV@Q9&afOd<
:_fJ1M7c6T62UJ5MRMHGPE>K]8+c=6CBJ+I?P4NIWgLJV-gC#UI?N2Je+&<2_M)X
f.cC_9)d3Kgg@@&fL\MOdYF(g.UC.]]MD1#6GMLX5d/SE3:^?F[_#VfMTM@?#7QQ
W=Oa@VG__Z^NM2bEQOY?KG45X]Qb)T3IN[VdK_c749R.F^929#0=2VU6P=P(AQdg
&5?c/A6:c>J:8;WO:G0Ge_J59c0F\f]5E]H2X9L0/f9BZNJ#4NEL)/ED?RMddg9d
LJIWG9#9W)/4?HMJFG3NCZ1O-C;IP@Mg/_.=E[a/6>]F.#6#/H9Cg+9_Zf7R+N_Z
_..cR799X5<R:[e[<K7D&/QZdMR4,^O(>CGLG]D69/9;&f>&c#WUMDAX.0O^&3F#
]=EWB7.WTEW<9L92eSdddc&ZQbb(aR\S+T,@O-&4O5fLH-3]:)HN5=.:8<=DVd.7
:<W./4b6_R)W;0DCOXOUGd<T)ODEC#B8#RK[55,BCOb9Q^M^fB?@D=U9#_OHVL/W
cE#+FSL;6/GU<4QL)dZ:&SS,O&KOJMZR/9JB?cQ?L0S(^L_.-OA[.K4#5RD82Y5-
b\OBAeZV(3SCgQ/UHMPV8#^O4\>dYN/]fK2cPMH&A4^.G.-=LgbC)KU(f(7+ON-V
UfD0a[9?3/FcD[V#(0N6WJSGeDa-OZPcG9Cc/#<IO.[-Xc-e(gA=J?RFO)]&68U5
EA_&5>L4O.0D0XAg8Xg^W_g[R>3/>dHW;Q&(X?PGK9^L#Q9^a<3MV.MMV@g/JB1B
&DW8\DOIL5BIa6fND\6MXV=R+T7E30cD#^[JET+E)-f72Se,6_AHR9:EXXLbDe:F
T?__bVNPcF-7SBNM^164b)OAeHNC.?:E>KM\QeH5Z7M]gggM2TI\NG7b&J8NJ[^-
<Y\;D]ASZ\R59-fbT=KLT]OQ;c:3O>;_B>SdKRV;YHNe-f4e+=.55Y=7.=9;]d5A
N0+AH1(Kb^V=#E[3(R/BeZ,\\-L][Hf(c[c=4;@-:9_<4U1GZHFc+P6g-W^F7\=.
gg/H0K:>8PL4MN@B-,U&d.R<79e.01>GUaD&EG\ec#8(5R6S721[5=:;2]+Ge6O\
D^<6D3QVY/N6U#b<R9@4#=#5c,6LFM_]D7E=N2^:6RA)RB:6Gd2<=:=@853JS1PJ
^L@.dgDK3>>J_V4QU.)I>])<FbcW-<4,CgJ8I^C3J6^-0>]3g#O<_?RQIBDeJJ8>
TK>FB^bRLGQ8K,#]efQ7bd=#g,cX\3UY&f:>YLcSTREf>6J=2S<@Ic.;FJN].HTT
^[?P^\SDc\-N2W28?2[?5K+bLCCaV_B>e;/g+YVXV]gc;8VHge1A;Q(Q<<U1]1#0
Wf;;Nd4U>-KC=.XZZf-g=W]F@V(eSf,A(3IdJ;Y:NLGUR.PRCc1<8:;XPCTKU:CH
+Jf&9SB:.)#,R\dXXKbYC.e3e-a#_ZH4V0<EZ<W#JfJKH/@N2DZC^C+eITTW,#GD
+E)LTe6EG]gYe8D0=3TQ22;AbWb;MX^g]._b=IB,_PLBGJ791a&XY\H;E4P##)4c
ZAQBYY0Pe::>gPa^]M2,](\,N+3AHIFZBRSa#30U9\2I=&b=A;(5)0A1S.A;ZKWe
0(<5O-<;b][9ZEB_,H?45)0T.#(:<0O>QVf/[:Q=[,\EGJN>KZZ(B5IC1#3)e[Zg
#FC:SM5_L0Tf8bL/I#7--[>g+GRHCa2FOJV.21,8YWd6>Q5;QEN0HfT7,;(-\QYI
Tg?P:U8E-H\:JggM5#D1DXY1OAH89I]_(XK=M2[<_??IMEH<1[/PaL?X0R@3;D(B
HOIC6[B-510gc?1>?<&.Z2bKO^&N^8OGV3:O,#V?gOf6IBCG(@Y9;7^,fTea[cO:
aa6-BR^>:MC.T:\&EHLN>TdWV(,?F^AW3-Y>)OFW&NZ@c-d^=TN[d[69L,Hdc[AK
F>^3/\P\Q>,Y&(KHNcW1-R[X&?S(_56RB)W(<bX?VH8BB=:4A6PTf(PNX6E<1[O+
Rg#^[E;DV2&gB(NFb;&>b]_FKEY&8-Qg,ZF5Rd;\RV[+U61Y5eacF6O3,@Z-/&?D
AX\d-EWGd]H?a:@JC\8#^L]\Le/V1>AbO6B[,.I&A_,<;S,F^FcC=8<[cFV^L)I-
0Q[GW\cM]a\@4T<HO=0A_?Nb0Hd^ULM](GRa>MS6(23LY;KP[<WF[S6G#,Y#6-f.
8I83d8^ALP//?<KFKEX=3,^,6D)W3J&N3I1MQGfN+W3SRE0bY36CX@T\>J:gQU9e
^N6<)eA[7A=&abYI9DC23Q_]A?G:0YgdAIO[=QdB#.+Y<GfU[fMT51JJ9gX>CA9<
_XV_-&ID92KDg^7&P@?DfSU4YAYVR4]4UZLd+;B^=aB9fEO<;#K[CF>DS0Z?>Z=c
D599_Mg;dD85d7K5@J;dfKI<I8CK:cXHZc/Uc?V:S=+8?GeKB9(dIAI0fGKZ].(U
QEb]#B1;ADGD_aFN^FKd)<?(T81a5c[]9A:3:#X+FW]J&K4++M.V^:12^LNWGKS^
+\ILX1(D)E#7/4HMT&4ZD<RT#<(CPTG\Y?4@BW+<bWfC/OaBeL@EF4\3HN2X^g9;
9-Ad-U,U;Te3.^R-CGQ-c&CRC0YD8D6/A#P9&UFfP>QHb?-DF0PK:&O_,ZU7?[M\
[NR4GbdG9Obb8&f1UA-_..^S<AS8J<,7.UYSS6?FgMP7&?]/3?fMVL?HPdT7=>EQ
eW1,/dZ=A?O@RRRM]6:Kc8JU]a7B20W]IcfC/;HZYYSZK:ZS=;@_UTM_,TZ+=LFd
L^BY#+^8E6-;4IH:;F-T,OW73I&Y5>DW3d4O>fGYb>gU-/P&cbId[-(@^#IW\P^3
UG/a[Q8BP\3#9^1E-(HU=T0;Xa50UBJ[df)c9@</g3eWB187aKRdFW?73Y]M>T97
;\V84e80E[UFYGYPEN9(bN[b8c>C[-.=Q2WdaRTK:\D>45&K3?Z(N,O@L^+O@1)F
F&^K6D:9H8KfR:a_<#/LEB;IQ?V7a7?\T-Z&V+-(>26.e^_G)WdfJGCdFg10E#L9
0X31<E;FWW]O.HXcCf(HIGJNCG8a3eYFQ7a+a+UWd?.]f#&&gC34Nb-79.AL<YIQ
\-fdN;gA5^/HWZZ6N^]=;\2GC/Z4HI2(E]7<2G)ZT4DXS#[&#TB=b#cP<8UP2f@V
W;FP1dI4,;ZLCK@[^e8aaO+NBf^;IE2?ZZ2,cUW]BbRb@fg5PCE=(.CZ<S+M^(V7
MHX7e1aYf/6H8e[b^^IZ.NfEe;cP:e9U29K&4P^R+I=J_?((,aX>SIQG<4XD#>_@
3BJB6>T6S3@4L?N0AG^gL<WRLdf2/[24a&)N=.D?W/\UQZCVa7Hg:[\Q1O/0RL8&
-.5^O<#H&R&>?YVe]]US+GZ;HA3/e,F?\,CTJ^[bee@WJF1D@-XSAP?/JL;5_\+7
c53#[dHe(DS&?:8f^4^FdVLcZaJ_HbI9>.QF66.SI[[H.M;:6L7UDPbV;F@fM0GB
JG^D=52ZURFFb?U(eY7Q2A?D@L_N1FT]#E+7H^16?/_<31XWNO,&2G&TV<c[_GFU
GY]R260Q47Z/0U,O.X\I7+C/#/D54^^R<@W6eZ0#?YSg,1,^:NZ&=(30=<4g)E+?
GR<\EgRaIC&S:1WS^\.LWe>B&5<>S^EOQQS7,5,HA.V2Q&fM;E#P_B[6VN/JA/QH
1#g6O-6H2=N+CgH0,SQ#,ECab1@fY/T;\f:^(Y2G/.Fb0,d_b/S;OGQP772H;IJa
)6N.T:b,9M:XSIEP\5.+@NQ]a;-JJ\,fX^0#9\)PTVf/>ZTV]X9fL9^M).&#dZbM
,cD==N&>&._\>WKRF<=GI.WZd#_QWaLVPRf\HM4BN@aM:JDZF]E\QYO(P/+0U7^<
M04SU.5_[J_VA#.P\U=ZX)^[H7#]6H[d)YZCZ\S1NYI240RL)c>ZdM<3DGfST0S0
XV;d<Ub32=f\JP_;55a+7D06eg&.I\N+VLYHP&()CC4=G&YJ&a[ON6Yc-TZ?->9]
XO2^G;EHLS\0&ON;WH-6WQL:8Z]H:(I?c?&V]SVXJ1R9#/KK=FJB@)e4OS.2OE2d
,9fE?feB;L6V5PGYbLf2MZUdR>N?7a<gWDN;;22RB^TIO+AWMPR>KJ0:6?EYCB?Q
?3a^/X#C7V]gRV[@BYdAV>^-XYFQRZ8)WTZ3SXO38#W/E\W52A-d,d&)(LZ@N:5I
#7K(@e]QVOUdcGQ</PPcFC<9UH:A[+06M/G=AY2;@Td0,XTbce<Y4K;]e7G5US&+
?LH@M=f-\f#,Tg?;M\c#[g+0(,A=_Kbg#YI)]F,FV;DKb?=\A]6D1U4UP-A/#O7D
Za8^FbXKSIW[6XTdUCXAHPXE/.5;H_IX&KK[P^/f8^4:X+_^YeZ^\>>K)Z,c5N\Z
/4Rc>N3<44EPc-J8LZ7.3.a8OP-KDV,H<&IW,Y\73O_gV_?CQL>-6Y^A<^aaA@>(
84WA&J7SI1,d798/14W[=f5-/9OebWU;K&Q:eE7AWU:RF=/1D:/N;G.)G9[IKT]]
\c5=ZPU6@(LcKOePQ+[9E)M:/c22g3Z]T/#^BC=R?AaT/UX/HbLDE#LHNL3\1DJH
S+BD@1L#YA-_V_W?19TaL;cGg\FDf;V-O:fIZKGAH(XY,B5gVEa_Sf&(b48-P#P9
^O-cNAIb0XO6H72NO5YQ(6O]_X;=<P@#O35OQZMOPIaU;3=S^7.K&#]fJK7;Id=R
@QIg,S>.2<fgPTBWSNVM./CV\894VbbR,6O^#X-e@9g6B61VPHJ^YFBa3Fg=<L=.
eK0B/YP\/])aY:/@5-]->[[9FPUL7J332V^6MEfNHR+K;-0;ODG>:BA+S]C>c82,
@#B,3JN9.G(Za18^:/5#KLVSF;UJAZFdSb4eKL<=FG,3&4B^G17Ug.._=>WSH:F(
8]5;P_+E/VgWa.P)#XT0OF)4E[=:_WbG/R8\6S[_d/&edPN.M?1M=Q=/Q,GgbA<K
#0OWR<OHSaT8CA&3PIE5:U_X]XQMZ=9d7C7-5WaRU3O+MC0:C#Nd+c@gPe)YP8;^
df6(X<QMLeB)&^@.:d&9S7+@)&_9[BU4(Pe-GV;:7)N/&Nf+4c)QHCZ]&BP2<LVV
>QLNJFKa3&G90G@9=MdHKRV6<)8VQD;.Q)(P6-W=#-g6T08\]E)_V]S6.4;Fd=Q2
].T&D.1,BUU3;\[JF03&EUV(NFE[;#-cNWdK0Y7\adY1gGHZ&:?cZN(;DQ#UX.R4
\Td-Kc?dPR_eG9)Ac.MdHH#QS#=1P]>=KFE18E53PFbT0:?X<bR\8a>a-L=(;fWA
LRa,1P5<E]Q?KK4D7_E,UYL#EECFE345?G6^TWQ3e8f>BJ9#ZW&Zf67D3eNG9d\W
718gQ=FX-=OB;4C9ZR?I5F(;:36MF3-TIUg4\:JD/C74:AM29))E8&\:(U<4(F6g
#5.250^g0I+;B?)XCGb^,X8:]FfYM3]N4]IXEV:cID^EI,^Y(R1LI@@2=)95=\0\
PWaG/7L#/OdUI2KbC6X)O;c;#]V>5_Wa+MWQbSXJL1]f&(/G8E)efV,:FQc@g[6a
S+C1(a.CCcbP8(P:A#E1/#LM8)d5-gU1IL^_fYaS=?OJ>SN_g\IMR:g=06aV+60e
?BGZTKd92Lg5c+TDK9GV,Qg)O0YcU#c/OVC7FE1U#F<b1UWGb.EMX6F=A&<>TRKF
J0E2C@6^5MW8>,.,gNd\^ab)Sd@ggBbW05=fM;UFDQfRN?5:H3B+08-7YV9C3\#&
g17c;O6/dE=8Df.;NHK2^.XH4)B)9Ga<^:)cFG>FH2/S:E\TNAX9OHd8beOgX0GM
/,79[LERQ#0a8]DZ0-/ON21E@Jbg-]5:5?a^&-MMZ=56]>94DGSb[?VLMIU-])D@
HIV5bBdS?Z/R]R35V>aI[]+&=H@]NPg@^.,]G#_5Ud+4[)eD)9G&:341eG>LXI+A
GL)9[4)+a@\.eDS3K-)5BEXf9cFMgWG(#._;W-_c7f0M6Z.DFbeABf:9GaP^@980
e+TQFCVF:+R#_KK[>Z\\AOIQ8:][^2?#+d/[d_DbVJ-RX&F]\F#PD_(4?E=7dJ[+
OMTJ2fRc>+]=-IC&b1XcadUO4-:d^,@BB<=>B@MYb3HR@dbJ1O<CIP2RADCTM[1:
TMP,<>dDAK>,9VOSU9c<Ie[RMLH[#)Mg,XG)I(G=0RYTBbbb3]\7fKd9?#URJDb)
9eKa0(&8<e1]Gd7^fDNDb3/;0L;2Q<N7WAY3PcARU?3RV;9#-N3[AG.9?cIV&Kbc
bJbK2g5OB7BV:/^)cWc+D(SR#_&/UI^_4YGR,VT-SNXQ&,W6VU..AUfO4_VaK527
T6AL(5=YJJQ9_L6>EPHFR589,=e54704Yc(ZK5(=6GR:3S5IOCR#MD(3ZcKHc+GZ
>(Z=7F3a02AVGXFT+<J2[>(:_ZM4+\<JAVA#QQ72<2_QHN9T/;ET^CHaf=e26BEd
[7G>RK&:Ed,LacQ0IfGfdD^dH5._Q5bQJG\eJWK60WX07:D9_M=_fU[Z1WEJa7?X
Z++ZK#=E<ZRCQS;MW\O_WKKdO5KTULV=;IWIbUUB3(aB^)JK+#47a\)BII/_HY\3
bCRF&WG@5f4WST>-dKEOUF<1WCWe&fIWDT^Rga3XcQ+G4QP4EZ?GE&4b_U68)UN/
Ib^^>?fV[<&ZMF+<<5PX[N8F(^agHKQA)F;_];Z^ARXYF8Vc(B,59a2gNXeOUH6L
gZ5D>Q/<g>(8VXOC>c/HaG+;Y>/b)-AV4UR10gFCQbR.7Gcda>VE;N;0b8Ae0J?f
:(Q0,M]:fJf4>&I<ZG.eTW\7OQOe3<<+/RTDG&aVeb/KF(4?>0gV=Q_d99OUg_X;
dY.>8I<R&JR6e4)9gSQF&d1C]0S@@gB:Fb3#EeB7M1\9,Ag)U[Qd]9GTT+20)S_c
a^[bT-37:S&egL+DIab)D7<[09M<.f6,,1NP#Bg/Y_P/1#U2d3\=,DZ?P]M76=8G
cF_fI9W\BABQ_5GE2G:F16I(+],+2U[;+D+c8>?\/GULZ8fA1f=.NV)AXQOQE,QQ
,#YYX3d6YS0b:022aN14C->c:9P94PX))OX-RdZJ3OaH;@MQ-GeE3#C^gBSZ+4g6
)&d^KIa)G&QAb=ce^Kf2eEUY)OI7fg6@1ZTKMbaf03_X5ZZ;PQ,@EV8\+K@UJ?],
65Na^^W(HHA5/M_<[c^.8++&56>7J.HGP/_&ESGQT5B<]&+W&^Va_HAcDgM)H(@:
^\B87>SE(+T\)2R(]dMR4<WH9T#2)A.&3[>I#EFUc__Y3_G/7e\7IYg/E#Q+da\]
HM^+LZ42QRASC-acbb<b<JUeGJ7>d.)AVf_-IFLZNZa\,^>97+Xga6a_,:PU,36@
c5d3\_@TRNQ.,P(<06YID,0(N&7KRDCV2;?L.M;dM/,3_c/8Aca=T7FLU<f.JCCe
I=Q]##61OaNe)/TD).Y79P6eO>S3b/I^3H?K]PV:;ace8ffU;2UEIbB07U-7H247
YNc,d\<15AUXbS=d]\GHKI:IgKSC.[)0X.f\,Z.V[/MGKB]S)X[[+;95Zd@YQ@_I
eb>N;OWf?SYU2aAKH+P9UcdA1--dc,bF>?G42>BD1BJ#QPL3+eAgJ\5\KARMC@[@
,f)-4OPdGBaF+J?_FY_DY_4g<=XgU)FW+K.=?N2/W+RTB04FSK_I+32Q0L(A:VB\
ZDd]:5ga<DJdcd?WO=bHd<ePBPLPQ_&G5>0:3,W>PSYAK\Za1d(AbX1W9J[UfGd+
YFJ3XX@e4-NNYA]XWX+^(G\:,^dO,D1J&H;6A&MNSd#f,VMICBXOU)FNV9(8LK+<
>L#(LG_S)7U@YVcG>-H>.31&bU5E>FX6eK5MB+0GMJEgLGM+E_-#?e;c/_1VeD[A
.4ZBS0:N1>_#^gM2K+O3^&[/4Z-()T@5&&W<RKW#a5QN[gZ&L1E>60>8edB/+-P2
4:PJ>Q&#7B_[98Jbe79<gFa<P[)CO&]b^?gVR1_N],_WI9FBL9b7XUKIf1?FQ]gQ
7AVJHK#4E\B2d:-CRXGKSg(6K#(ggKYG0H1dUW,>Q@=(LAab>Ug)Q;L=MSN:U,5L
\,S8d8)F#5feeLPZTT5Y-&Bbe@F+P)I3Ua5<]#aGKY<8((O]#a2bRJZc0R)c.(d0
2Q5bf\=Pd?W5EOLf6.MI+Q=T;US<]NbFN/>cIWOTc2cT--\632KY+7XVeGNdZHUP
98Q=fHWDN<8(M2,/=TG7UfQCcB&]QYQJdFV5adYMN(W5T-d8VUUR9LM=FN0eRa\.
c-@JQ/IV@9.AOQC6&\fH_BOHA9eY8O<IQ>HgfN1U-X54>9NcIZ<_@NP-KK:#91S2
L5\F/=H,Vc2RX]DT72:XJGU4GH&-431-,@1<>FTF:[C7U:^)3EXT7AQ+F/=79\_K
\,HEN4;&+HJ\JEaZgS>cGDGAJ/=JMU/8@?CC[JEB.=@#OBOOTPc:N>;K:A=bQ?_a
WJAd>BBg:<Y<Z>Scc)_cR+:UZ?9,bbM/,URKT.2V#4M7C0HO<QP5#7(D_G+9Q^Z#
bKGMNF#P]=ER8\IF1RAT(-)PUJ1W=[;HHBRgY_@\W[<#Y<eZ\&)0GedTg:La?M?D
0CCQE_4+554^aL9f3DgdCF-TSJCNcSDLI:)W2K4J=??^@bHKJfX/@7#)0N_GIa?U
GJ2Of4,4M8<#[BZI7@We_Y7YX80]V3>Eg3gEAO?DI\M4ZW]fQK1=@(V@M278T_(M
dae1LC+,d<2N0+e1CU)Ea9UIc,2f26d;KfKd,Hcf96;)P/X#>=[f;^Xb#-2UZc-F
]P#;XKbM;I3KAEgT@?(F5FS,D-QB>cRL+5L0a:c&+(GG5YQV+fTX\P0Y_QPaWeYf
6WOMeM(f;K^5R:f\,3SYD-D#>2_d/T6/@F+7B]P(Ea:A>@^NH:^(a[.F#.BV_OaE
B>V?X#KDFBQ]@aLM,4?;.g7I:NNXWF?.3OWII5=VHgbVMBa1;KDA5EXI5RaP&g^c
:b?50Rd_.25IL-TDV0H#@I,?+9E,A?_]YU_3]QMQ227/GV81()@Zf0G,9FPM#C=2
)9Uf1V?JdbB0@<@g8(,-9e82F@_DEfU^C42+.Z0>2]:G^:2gQ]TcgO470+\?QDU[
(V3&d4=EW,X<&I47AeL8c:&aZ>cJd?Q6J-QX5GF.TRU6Bd07g?/7.<JcQSQH-=V5
23AfEYY96K27)Q(e,&ORY7)74J8g=.6dg_?+\b><Id82Za,,?>Z:eN<#W+R0005K
]C+E55Q4eJ9<R4P#a+bTU[^g?2?ZP1V.O7IWPH&)9f9:231fNMISNU:K7c)DGe:^
->B^#YMH5SG.G7V(?Ba5Tc&@0Z<^dMdWK4[?_XH6?\\5N]PXID>I1D&FRa81.TV@
X?Q5Mf4c>\@#7W&,Da^8OV&&f/73+ab4J)(MQP>gH(?7e0McNU>XNPT5:EG-#2Wb
EI9&ED5?c+;;04<,();+R60YaU4D;e&5OVRD:11[cHKI2M[[0\.fe571(7:eB2S6
U+CHc,74;?E:a<.^:^I0c8OR5QVE-_Q=3H=<SD]?IaPU:02XCC9a=\Zb.XIA+2&:
+FBEL[ZL>P^WGfCIS8H4EfPM4dB(L24=;^VOYTF:YIPOH6066.(#RY&aMc6:<EFc
;MRS4-];&DHT.Ka#H1/b7,M9fX)II2.6dX.=MDG,9I5CeFUS4@F+37JdI;LH7@NT
4L#A6[2+2/b=M2Q)dM;CX4c/&Ja4YF7:6P0LM#HE>?N)9aKS1YgCRR]YJNcQ,^6X
aZYUW]-(M5>DfLGaFP@AUPT9QMK2USKOC-aYd&g98VU2KYc(;B-=&N<.LB^RV>K,
;E\(&a,RX2X&GP9ZZRW)U1KK@&#XST&B(>P>\^=1RVC06&+/IS6#0]V?T:0g,?)N
0=R.+-e8[OFT.^dJ3[YfDBBCaFGAB84([8L?BJ]6X8_>(KM;HLd&@A^G4??e5OP+
C6B>HSK\d&4U5>>:C@WL&I+G>V7LD(;a#CTO.F\<,RRF,)6b#,,IR@MgOb=;P6P>
Q+f46._H@DSIK=ZQdgce.(BEaD\BD@KZ++=<\3CTN5TND=7IE,=?\c/;.P<W@AJ,
+G+O>.2N]^Ac7Y[cXFg_L+-C-J\7>AI>Nd(f<@]&dNW]F+0<1<gMLA.,&OFEN9[C
#@C&2bK4@MSHCV4AUE.L4<R<OE<PcJ++U(a<DX4SK&N.H&<]NF19.>\2/EVPKg<F
\P,.5-Z_A:?8L4BAbOXDOGF;&aD2W)<bWbP[Y;5\QJ+V3EJ1af,A[Z7FXO#\2:\T
CYKKgg1&?1X?VX]f@N1QXM>(^;d(&)EY?(D:0,9D#P9d#F6E@@:b#b&CaW4\)\L\
[V[N)eF->GeCK#5B7_@UUaa/GX4FCSV[#2I@#Q,c^L\B0H-=+:[FG;:5,HddRGgd
&-=>.5TA0K@19TeeO]5-1#)[UfX6]PZ9R5L;>5/TBMe_[>]XE[a2U&)=,GO:,GU[
Y,EZ5PIE)/Kd-0N^Pe9GUF_/M0DNVY4VQLY/YNA;C\gG_MY.C^B+?QcRDZTDSOG9
YQ.JS8/G+.+8II@J8VNGJPe[SV)UJEFY;?5F#9[#479=QVe)c:b/8Q.=#eHZ/;K0
@2AG>SCMCcZ2;d0RZ<Z4FYg(IV9Y4#TA(U#C=#+dc]/4]2\:GP>c,_UA_^-B&M:b
V8YK/&W9dJOLYJGZN\1b7F3&J[/P_d_).0PT2)V8K5NC.M>^L3g).-THa^-(ZM^=
+>90Y]Jf9C#=@1>&Pe3MFSM:(^E_6@AC#I9GJZJZRPUS[53>-<(&YcXSV9B(,_M=
(.,EMML)UC1UM4<87]HGKV=)/)L5Zd.P44_Z-W&RUQ7T.K2</B2ESeb428Ra)-W9
cD@@a[Veg>-9S&8+FSP;KIEPE3ORMbDPUX8KK[?P9N4MdW[TbgfK>,a29[W:LS+\
D20>U&R4b:<>Ka@PU074+#dbP&>Dgb;1-H/UU@(c:1_>3V=8N^Y?8O-6f-?E)Y:c
b;>]@>IJcP0f+GDJ5)d@.)C(;D;M^^EdGd>J.][_YWa#)FU1P193f:N)a+1(YHU\
c><-:6c,6>Y&OBNX_=4cO9-ggB:[RK70+XZ1YIV>2LB7@Ac,G+@/Me&[RB.&?f89
afUf>OcGbbCaMUHDDR?7gU3G-P]=\[K3JKLA#NeS1J/./b_N9f(;>;-K1C)/.RVf
1(0E8N_)];L>#]7Hf.05C?D7@c@?[8+J_A7BY8N8:A&UD^&QSYE4)NQ&,cG-5fW&
aV6CQb#SSYLKC\(ZNdWX[U<)6=^/8W:41NfP2+Y(Y<I1a4BKXPN)CC[.?LB&O],B
&f?K9E?+11cTF:QC^BS<89EaP:a\SG7NJFeHQD08UD\#K3OI&5XHWPWTV3QB,-#K
53.?\8_5XG:<_D+LC<7EN3^UMV2V=ZH8T:0O>3)dF#6X/CRZdNaKR_8&YOARdFXJ
OZ&<P,69W3LM@CFM)bJ=Y-2D1MDRTRB-&AXgf/)Nd;AYJOBG+&+d^c=ZB?WG(@W7
?/<R2]/BUg(:D#/Y2GcMg]dgcS]be3U1GDEY)5cb5_eX_96<H,[D-,QRO#2eV]2J
,2_ZHBP(6W_11?AG5\?1c/T#O7OJ,-g\N6V<Q6\H=RO.g6W>IA:_F:.?d1dWW>>B
H\aXSRGHEGD9GV?3-d2=@97F5]cH6=Za=&XXdCUA<<_XS3+.AF#U9@eaNBIL>ggC
B6E]:?cgKMbQGSM?0X6PfZM(Rb@,f=MUN9_f)PXG;XU0)0fGc[LgQGa,W)SV#792
P=L&-XQY5@C-GOAR4?7BB+&IS5SC;a5K#)bT3/NXCgHdRO2>HU\WF]8]A(-@Y^Y+
g/6E3EMa6OX+.G:6bM=EA)=eTB5<G;TIYY46R6M;NYU@RV&dGOE35[?L:Y>;E;U]
B5>&8H(U0__C+0-1)TL,UecS^4.<SeV6Cd.55\U62?^OIDRQQa.UT.>cfT(;7f48
&\KX]BMH0/4:-_.cT+X;2<&2MG<O9Ie-C&b9cIR(]-HBT>GQHOA;E(V[?ASa_-H7
,2FT2O?3AE(da-Q.ae,TPB@Z+V]UZS)QX6UB>T?aK9^A4L[Jf9f2#M4X]a>:cfG)
@F91--c,D5f54/N=E55B0f_MK(RAa93[W_J+@X[Pe49]\-.:ZJ^,)XS5M/eY2WK.
0W:L[JV#VEI66,@e4;PZY^AbYT6M74,,?\DR.Vc9&>V3;d^]3^L9)_.\>a@:Ve?7
OLFEcUPYYUg^Z-U-A?GF>Y;2@b/<(X<Ca?32Q<-\KcW]P+#9#JE8=RZ2_aegJG6V
a69TE#=[:0/?@J/[g:/)70H3KH4\@5]GES[cc3WW9BQF>gC4#KdLK<D8L1D[_RFB
J>E;7K5]9Q0ZfgD=Off:AY,5C^@d40#&8,B[7EU@(47#>B-Vc-OG#>^#:,Xg#.4L
M]Y^]#a>_BfNIE2c3N:N1N2eeEX/&1e-bHOZ\8]#f0C1U)C)cOJ?#:eD:dF>RdEL
U+;U0-/ML>J<cL;)SKS,[=4bOGbA\-KLPe0X#58AaS_2CEcb=NLTVeHQaSL?]L0@
HPc820NK5=gQK(>=6S8^A<.cgRPLeE/+W0WOV#^Fg0-FeT_QJ\IcG]S4MK=-G)P)
U2-L8P(O>2O:JC7LPWK5#[-RB&,)dLBbZe[\8B?cP,A,V^8AN92M1b8b=O-[VM3M
B?SDUaZU&L>8aZIC4:)@B7dbIG2^d89c.KB8&X33.;>UQS)0TcYO=NBDU-gcLCW=
#6IQ5c;E.f-eG1bP0BH\/CD]E6>eY0ebe-&:E,3f-EIfR&T;4@,3-[46>g?dM84(
a.-+1[)H3[Cg)3H0EFC2Yg^Ma+8^5<X+RP<7NMG6TUJR/1C6CF+56-E)eaM>GA#-
2\N0L_A?3761UZ7Kc4dU;YL+[PRSbeAdN&RXdXW<PKebA2]8=^0^H+XWHC-JX^7X
Bf08ALX=f-.K>CeLKKbMX9GbR(9DLSg_>MBV+[=U<_TEfbOS+-R4M#<AedT)VgKX
AZDG=)43>U?\GQ&1S1Y[c])AB[GTR;VQH=[_=NXSMeWIILdNP8R@I4<NPS6AKP6(
9[E^X/TXeRF\BW4Y:1O_2:f(S:g/gG;Abf36K9F;IJ[Mbb+NJ@:DG[3^(@(62@)L
0@a?Q:F\#C3eTa32TJ?=2.Y>+_S1PS\@FX;6[FF&Cd=MGP+65;-MLQ88/0VddF3g
1,-cGSWGV_>-F]7044>-b6RDJ;NQP&6-@f8W?1)GQUgH&[@<c=Ece1UA.aVMZ,gX
HK7d#@@cX8dYI,bV1=DMeJ\6fHVcU6.;2>c=PT&M)^]LgWAIO]U/L9DTJ3.@\75X
B#9P60R>GWVXIc7PF88S(d2AM-)7+,gE7F:(@VI_H+NCH2]WJEG+90Be4(\5SRe.
@HF83eX&PEB<9d=<3(^2.d0NFND\@2Vd&J:Sd0.4OU+=MeHbRMAT]3;Z-dK,:#OS
=eTA=>&W2_V;FR>8DDUYLf)Xd25dfW#c57f<.(FNgA7T^W7\?YS^#+TD(-PGDW=)
[FG=9J81>-L_bG>EJ@:52E:7@PFfGLE@JLG0/]@aC-;4&@(BB6:4W5,#IUHfJP\O
@8[/NL?O,6(?H808I>FeG6Pe(+PC?7]fXcN30+4CSX6YF=.S(WS3IR_0.HRXXge>
cO(0/P?L-BSf;VOVH4eGMC,@^?1aX3bXT0:6AW8dRSTe22P<:K_:(d=3TddfQEU4
=29gE#1PCISOBZB?49c>##dMAP_@U(I]HQ>/W,e2HM_gH4DeRHb8]+KE=0HfbOfQ
b@>-Z,7ae32)G0UM&:H&eMP:A/N):c_)MTU:]UGGJ-:(Rf_H/H=KV9E13U;52Qa_
.AOSZDa2C@Ed?#L_g4:eS058_90C@9_KNc:afKf_3>G65CI/?9b-&,dU8B#1eFZ>
UIbc7DZdf2IG.S)c,&TABGT968.9K^,HW&U@<#M3_7Ha7@<e)G<d85USHE8?:@-V
LE^9KMWB;)(@C(Ig1]O9[3.^g>a]2]_b)Oc.bNR/W1a,W8N/5(,)(Ic(Kd6[(19\
BSY#&cTW<^ag/<+JH?D9Q,?[R??EUGQ<7ZLU=W4\S7(GIM=3bKQf3>8MOg_P>5W5
B73.@3AWI[Y9fM202R>-H@8WDJfPLf7=T-VXR?;ZV3fK^A(0T\73UdKbZ56F2feG
Z06JHaHS6I-T=Se<MFE]eX^;6(H3V;)KTgB?]Z)&D;MbXJ(UDLT]-.Y#?<FXT,&a
>-A3M5[[[W7[fWBGfOTTN6KQ@bO:EOY:DS<c6FMC6>LT3W_)1OJ\EEXFgY,N_:R;
VQAX6G2]6<5.DB;cU1dY>Y&CYIJNL[?e(290I;f]W8J@5?^Ld[9.OZ@>.6):U_1D
A9]>\+NI(DJM;.KC+32&;C\3Oa5?J\1KZeZZO)WQ.Rc4L7eN\agW+;bd3E8a33#R
SES;DP]I,C>H@KJ=ba3^IRU#+F<1NOY:LSFXM&eM\GbQY&c5F=Q#/^6Ia?BGN[EN
I[ZI4e8/_B,AT>PWba&8>7_1Q-W<9WBAMPE84V+7eSDKTWXeg3<__#JUeW6DE_Zd
;6^+]If9RS_;]eD96L?&X2)V<HCFYHHB4@S:?M/MJe7W.?+LX<baabYFaCALB.3+
VgQUYV+-#4;XHb@^@:)/EFd9AE:VZAY\Z8X5DbVIaNV:\VGZ>Wc5(3&Z23cK1<dK
#P47/;FCV8S=G(3AIaQP))D@FX;[<8d)#>/U3+\(D2B^@@MfBCK:Ad.?]>6+K5W;
:4[@32J6/JUVU.4[##c(0LZ3\YQ@+ESZaIDM@BD)7]cg(e+19A,-Vd-)L7Me9(Te
&JQ,M8K8c8S/8ZD]-):.ZHf1GRJMPVRJ<ZFg\VEc8<6YV_a3+=Q^+:-6c9SM7Y3^
#0N/8VV_?5=,WHD7Yc._2BX@aUJcK2K1+^KK+e:Q:=7EC4QKMB)+4_A[8eTEA<(B
G=Xb)7,\.M4@YV5U@B0:5SH2Qa?S_YU9OCbbNP^#-a-;FGR3[Me+F=RefL#0^TPP
,4AET/QC\H]84g7c]D/U8,f4ZS>#O?SL,X^<@MA<?+gb)0gT?4:V7<UQKS0N72+Z
Y)>/ZFISRJd96Y0O@YB?>8R(>.K7(95KCd>9F)4Y^fVd;?\89b<HIeE1Gf.+<]Ug
<P/]O]ZN\]GX86KPY1gQESBELb]39ES7E#BKYCN1+_YW:S9d0\Ga0PZfMeIc#aY;
E4IY<c[;;?LM_PbdUS2UgLfNCT28NIa:2:?QE>>POfECd(H(]G;10H#EK_QF[f?.
9#K]H;??UMY=K0V664@A_W4aHO/RfKXe:V:E6E\2[7)95IXeV=H0C9J:U]S;aff:
0LNCX=<A7a3M@:Q@,dcHgKHPP6Cg]E8\.)ITbaX6(37P3G[.VZN;cLJ=Cg?7.WcL
4?NL;b8U>^3,3PG<:Tc+B4[8,U6YB>7OXZ@dREP2;:#H)NUKVR4Le-?_5#c0H)FC
T>3?)B.=#1C0(8RJ,6A6H2@0aA9>LZB+T)H&JC/fWfV&WP>.,5CVG_A_55\I6>SN
AUT(1(]PBI8T/?(Q.(;HSN97Q]d^e]72VO>,>_N&/W(]-5Aed[CA;6KDb[)O9-W5
I+58Wa[U;R]K>)\F:^4_+Y@+a;.8c<6C7@J37CT>9T_W=Ad.B@N6PgB7:YI^a,bc
&;MSR;G/Yg:#[N8+A3g<eGVR5R;V^HF3a@E\L=O,c7Lb3NMeZ]?[R.3g=K+/GKS?
=#)MM]F)dM7?A[>OA&F6ORAeGf-=fT-GI&51GYHZ>I6F6Za]I;T97Z4g^.XUc:(Z
HZ6JR@_>Y/@H+4>SO9,2P3E/@[(_=AWLN;(BJ)6PS#X_(Q1Z(OYeC,X.7)bJ?OH@
IKVFbP9&]a_@FQ7,CSWX#WbN>FfJ/c(7,OeNA1S/CJ8YQC.c41eY;Bb+c84R^A]d
=WBI5841DXJ5NHG)a=PQe\A^GG6:HL#e_4X@:dT7(L1YMVL(gOU,9SCcLU61,^Sg
dJ.IFBaSe(=^d9\Z:L_6[CBTLR#S>T>1CBcNOBZF,fK1[PUNV4KIMEI#=[\0U?Z4
J1E<dgAB#<<+#<bF]D3NH[(]WL7c+B/>?a?72WS8>\E4c64=K#eOJE;7,Z+g02bW
P34_K(B3J/4ISJ[+Q,Y.63QQ8M<G4@/L4.E4Q]&/e@?EV6-GLLP@EZCTOP1EDT:d
LG/gF&V/<bB>;Q,H\1/]_aKN#9A4-;_BbFKH?289MU@fWEc#SW@\C8EQE/_PIQJ\
H(M/;\^^XcD^ecR0=&>6-5f2APe5\[[VXY](:>AYH&JM]Bf;1@g)XRA_F#>NSIf=
dFIUe?,0+6)AId78(PUf/:6(O@4Y+-e^Y2b&e++2BKg91UQZYd#\Agb/5g3cQ3\^
?[?5[;U53<1#,\B-ZC#cK8TWPgPb]\\Ze\Oa\8eB4#We9ZD?/<(\-)8KJ8G18VLC
;C[ZAPHK4[)>WA;H\N:>ITUGZU@Q/C4.59,PF4E7a+A74=?fH?RVU-\eJ4>ZGP?B
MI+LB<Gg+?D<UVSVG52QH<NT8Y+U\7.>3Q(U/5.#JdgNSUVEIT7(QKI&7cbe&..;
QMRO,3J<(=^PW/976\YF/.PLdX3.?Ac#_PJ/S:I_ZL@_<XCY\P=c1S5O_3<HIL8T
,@U?:8\--.83/3B4926X1UTGY)b#O04A3ZCQPR\LZaO2g.L8e0_Pa/N-4^ZITNba
99),4-0</((Ua[1W,K#cT2(9A=J(4X]Peb1(D>UIfSD#I0aL:++&e:3+-3JOBD16
2#CFU-K+/83ee2,:)fY_MYCXWN(>Z=I0-cUcD<gP61P8+_L7P7efSU]_].L4X3UH
PbP.5eS9GKaQL;H#5(@J70JEY^1)Z.O5eW3^4C>[bbNO,BEH?-L\3_QJaF\=A>5;
Zg0&<QQ:.1:B/J)]4RW-QFG5g2gR3<TO\a1_DVT_GAT-;<]227MNA-aL=\WUGA/1
T/\E,4;[>72#G_ZIZ.#B)a6-;OH>&b3Aa:JN>g5RXb7Fd42JHMbNY9c>;L4BcTA:
W5,YHR2\?RE,/E<Z\472VI95a#=(e7Y,^D1K4]/5^c&9T=TUFb8PP[GS)3/IP0Y+
7KB^4g[R8dNPC8.2;F>SLb.32eT61TW@?aFfF@>eG57G8#2eAL9):Sf9/CTS[fG(
[&7WKNQfeJPf&d5A,&/3[,0A=<^>/E\Oe_G[B/_&9W.C#\05/25SOJ0JK5PC])@9
>\K)MHBOC/3XC\G^&E]J_-(>MBMg,(Fg7ee?O6[OA3Y;CL2=CeDB0aQ-2=ca-aD/
@2NV[WAFUC^D.#=H4)D;6f#\]\<L,+G8XXH[#\V2KBHg[+8b4@^aR(gR4Z5]KJQK
=01XBEGXW-+OX#PJO&.35Q23\-fO7Q[6B/KSIBf.6&)E5;EX>f1dd2cGTE,B>]=f
a/83@QYZ,6_f&+3[Q;,A][7.9:88cPT>SbC&2OXHHVW&OSKObV7b9cL@4TgXAIQ]
HI0Pg3AT:;e4C9Jc[c&L\gd,NW3#.F4TDS(?b8ODP>;Mc]F&Nf\6A3F=>4PP[/RV
IVC_2F4W.A+,@fGO6=[Vb#PNeN+0GQO9e9,g@M(L_AJNgEUL>L(>W:/>N1bM=<\U
MT^beQ7:+f,>T0-W45>#4WePI03OZNYdGQ>eK1cKD-a6/OHTY;B+?cP#HEf.P>Re
3#.g@P3Cb=cTa[4L7#7H?;VDI>[SENA4&@6[OOVc]Q_(9TTB&Gd(>^/FSP6:24;]
(_S(GKFe0QO^(=L(6Rd3(>;7Hd.bVWGbUJ=+[8Uf1_;=0]Ka@6&CHFE5QdMge>R&
BA^XV4faQYZ[)E&8OLe^be3Pf8KS)&7-&FO0dg77)>;8-9/H2?M@@6bY)9Ge9?0[
#>>KH.X:=9N>U:deMQg7R9B^U\M]5#^O53(\V66e3(3R,.KF1Yd\SLLNa5P[.>?[
^968LAB@O.PT6^Q_Y[4A#Z:TXBU=6a-\,bP((OQLMIWJ/F1V0EdG@408/-L.b^U\
f>6^7KH6f?JF1(?+H>1#9VDN/5F>:+\5HYa1[9#]Pe+daZbP?aU#&5\60Sg[Ig)-
K.aM<PeM4Za)_Na_Z3TEYHI)2IP99CKR2#F0+.VS);c(4Sd1CB-G].@&aIB]#-\8
XDA1I]VJc(+#>4a<).Ra<X&ZGAB9QW&WCZW<-;BT28H5eeZHD[J\JEA&\.gCJA(H
RIB1KLeEOO+XAM#SO^cJSc&YCHcW18e\>&dDQ4+I^@Rd^8EBU=AW&.TGWQVJ@X(X
3MZSM7+&VO&N]Vgcd(1?P)0eJ0I[Q^VJ1<1/H?(TBGbM\X/SFe<X5^\:FA=17e#9
^XR&QI<QY]=/Z]568cL71L+@e)P]I..P1gS]ZR]39_VYf/Id2&-6[G2/JgMgQS1Q
O09eP;;K[PgP0XC87/]1.>E#[KXX2bWEN>VE[6O+dP[UADfQ2X_XB1a89KD_&0W/
[@+<e:A8A._?;aa86N9Ng(c+\b^1HeP7&.-,L:H,Fd<H(U4I)d?bb<>ED<?<9b(T
C4L3(?JW/L9^9)Q.?RBIa,geV74W0R-IC>#OD==(((:&XYg]>Tb?0T3Z;U&XX3&[
(F_fUCc0dTfY200=[6.=a+=]J;Z34DEU]=GQ:OTBa;JTXS)_1U2,2]b?S)GQOORc
?-U0_OSM3ASS^8PR:AbX\U,M5J4]GgX]F]+bS]_>g\E-Of:20bG]D@#/2N@gYbY;
^J2M]HI107=^)NOFQ_cUc=7/PPaEFJIK[@H8L1SWB+219(b8g7(>HM<HQ;fODWYL
-J5DR3L5@@JcC0YWd^W<6B]/D61KMR)CL;3>>4eV;@VU/HX5eGMeSJZNO;=X<;0)
Y1>.](&b.I,KNeD[U)3a:\gdHfg7HNZd;.5U[(A40XQV/DC4FC5IIB10]@V,UBg3
K1g1ITA+HWR.^1Od5[SP#G&R&K?M.\<:M>5+(CL<-GBWfB(3>[<EcC#_F+-F47eT
:SI^c5c3D^0P\-C>C1(]QP);F..&UBfAgNTNa4f\EP7]Q,70.aI^WC9&G+K)^\]e
LSdA.)UWe0U5+TH5ZJP&,:_:B#:Y2^ST/=BKJeFW<VX&S[GU[]e#:19?G(.7/)_8
F_L.=<g.XcH#<54LFSBg7/GBTQ=79Q5Y,_YD3gbP8-#98+3C6@#.F&a]Y@):T8(B
Jf@EYa6?G&M-eRc0LW@:&PG>7ZU>-3,QZUX:_+@&3S\=NcCC/b;7&Ad,E83.S^P,
>=?2V[:ZgI)6EEHMU:Jc+.HH;Q#N?=LESbEALI5)b>BgEA_bLKDf>e?KY./K8dVf
H6a6e/STH/(X^VTG9SG,SE+5#^@(5#gDWL&L3[4]:^O4QJ.38.>UU3TF.=W8Q6SV
U2OZ\PG\C/WeAF_C&6]0JN#U><2Y)WHF@dS4(8d0L9D(0;b^.]PZE5EcPH\[,[,U
6M(F=?AL9Z9fb/4e#RC->9#I7Q?OPWU(e8UDcYA7>dYA/bT.OXO8[gc;MIcM.G].
E3GS#W;UgB]Id.:+QaZg9WFZ=M\-5Qg#PBH3QDa3O:KEJc2>,658Ub)U2.L7_QJO
O?&A(1<KQ^49>J,?,2>W=\J?[?RP:.S+EK/GeOa(E38J9fdU.9_1TOX+aZF[?[5@
U]R4)P;8g56g^?/ECAeOA8)8\-7K^8J(-,-?M5]N&Y(\/V/L[7aK]Mg[Ob;UB,LM
20IWMf,T?Ec7KU5,SRe-M+K1Y,NZ5F89GUOfNg]K5A>AL1@#Y#O9(#W8:0&<[=bW
dDFgc/1cFBd9N?OO34fWZ=b[CNHNH=;=CL(?ZPH^WaO?f)R\:Wd70BE<W8dPCQa/
Q:CK=/[N,/CZ>XbVU9a,,TaV]+(F;c6^O-\)+AVWf_G_3dH.2&L<)VIL.H4L>)L)
4,geOW-FE;_:PVcccdX)Eg?g47EfT3J:X)gUO3>KM,].(4KVWMB3?X7?W_6DTdMW
Xe7E0&A>VI\+&GF6F=:_QdNg]XNA?C4BNeW@)F[b55-KV4a)RCUPVX,B3981DV\T
.68bZTP4=86)DQYB.+EGSeg5U9K6PNc1/,Oe)#J]8VD<1Nbg&.&>)I_=WE,44R\#
H2B27[VPe1R_d]HHEUa?^,8U50F_,R\;2,FN=;10+1Z^4:?3H4@X=X0VAB.IPTJ7
<V_+FCa-Xcc9A-59/@O+[SBTF=@7D.E[BG#(J-d3=^C,f_@PRY5VDQc/ffc.;+Ug
-e(#ID=1ET9(0606aLV-Z3(,Q&4I)3X&&+3<S9Z8X/Y<Zb5X=7K2CG8TOAIg@.8A
(>)b<BS)2VgA#N?a(4La_U)5f5Sdg_Bg=777Pa\]T,fJG&1<[G+^NX;JdXOHE9GE
6?4gB<JEGNFfdGT1:;aV0KLU_25Q9dNC_X,SJXMLH2^NG.4dVUOEO;_=.V;Ha[L(
?=0_7]JBKR-1]+#I8\G42LU6>)33])F)6b3?B.cCZ7c:2#SD\gW>+dg\@ZIYa317
C\5cAAFAVPKF.e&RQ^5_c2#ZPfJ1PON;3+J[STUZ[E;=^VN8/He?>&D&1(>HfSK7
YU;)4&;#68EC0E-R)?&F=R<gXTH5)>6;\HQ]HSR2cd>:)WKZ3YMDKKb(IP2_JMB>
NVRU2(L8I?9U=PF=[b?M1>GG/,d2aQ()TGK(2DP2BH8XF)\N[7[Q9I#]NJ_>H9Yb
5]gCIUcZ.Ta;e:OD@dF^T6E<:5A]C&^WG)\C<cLcBY3aP)ZTOD?BKe)(RWA2TIbR
(1G)3^RIeD3-Sc;6.4=V9.>P@5-NHE<Y/(V@WYY)R<_Ee:e_S[I[Hg<],<]D_f5L
S_O7Q&;#U2cc)S;#f_\aT,d?QBT1F-3_F3OGKcg3KT-S=_Ka,9C;32BKf;I@geF:
/1+.CQ&P4B3c/5RORIZ24]g1YEOZWIVB\3[GJgLD)_0b2\@-N,P-F?b[L9bS<?6B
\aMgGg2\TGec[QZICW\:\W-8_,Y3J:5(O1M@U:G)61L]B&HdNO.^H8W([\H+aW=#
)d]Q#;E?>+976?9ZE+C]L0)3D/9:\V3/B&Q_E2C]aE&<.3W#IPSeB2Nb\0PQ=K,4
UW,LOWe]29#4dE[>WXfJ/6g&1-.^WFL5_2gS6?fF(aY>E:SNNYL1BSBg&=T,5DZE
D_ZLH8-OUF+E#/U9S_QY27+L^5TN5gKY@:.,3-gJPXHLX)gaEM_cI_RQ.D;Mb[,<
1=N@^K0OTG[(/a89JV@c&M>4.;,O9.FM@4XJW6<WG-f4?LSQUgDFY0[7LE]XH8Db
\DBH?S?[YQa:_H^#O8_d?\+5_NM\@V(Gb@2-cVF+gS(Q_R;9^VWO2a4(4JF;-#5L
cD\Z@\(W2JVOU,3bX@Q7_IV9XKI2_Z9([W[#:NPUJ0C?K3\<2D<=JaG\E&L]a05;
+:/3#\HWJ-]bA/Y?\4PPP?a;dcMK5:0\<M_(.:^Ye-9e0gg6ZY1:QJ?_Ne;.:e/F
#;(Za-b0^\-BERQYF#/@bP&FHdecHd,LgYb<:9SPN<0K#\0_G>?g#)9eV[@91[N\
#)AE[W;XSH3L9__&-Wd=c)-AQWF@;4JOZgb4,#V_)F1[A<0B+]M\Mb9BcW]GV<E;
E6DOVK02E<\IdN+9ZZK8]#EOX1.W#QYQ(Q)ad,93G(4dd-123#U5JKSC/f8(V[5:
:aBVF7JUGCGeW)K20gSfHDPcT(cgg?.1SQRK+RMY3A,S2[I4B=W_TRd<(UK]NBKX
^?5dS^&:(Y&=Q^6g?)QSUCVFZG[=]N^TdGNPK14Wa)^43Y]T&3RYOM_EC=;FMU9M
>)0\cac2L_^:XUSaS1TFP&cdTL7L2g6,QCd^YbS=,gJ^H3/?SAT#/8_EI$
`endprotected

`endif // GUARD_svt_axi_port_monitor_pa_writer_callbacks_SV
