
`ifndef GUARD_SVT_AHB_MASTER_MONITOR_DEF_TOGGLE_COV_CALLBACK_SV
`define GUARD_SVT_AHB_MASTER_MONITOR_DEF_TOGGLE_COV_CALLBACK_SV

`include "svt_ahb_defines.svi"
`include `SVT_SOURCE_MAP_SUITE_SRC_SVI(amba_svt,R-2020.12,svt_ahb_common_monitor_def_cov_util)
 
/** Toggle coverage is a signal level coverage. Toggle coverage provides
 * baseline information that a system is connected properly, and that higher
 * level coverage or compliance failures are not simply the result of
 * connectivity issues. Toggle coverage answers the question: Did a bit change
 * from a value of 0 to 1 and back from 1 to 0? This type of coverage does not
 * indicate that every value of a multi-bit vector was seen but measures that
 * all the individual bits of a multi-bit vector did toggle. This Coverage
 * Callback class consists covergroup definition and declaration.
 */
class svt_ahb_master_monitor_def_toggle_cov_callback#(type MONITOR_MP=virtual svt_ahb_master_if.svt_ahb_monitor_modport) extends svt_ahb_master_monitor_def_toggle_cov_data_callbacks#(MONITOR_MP);

  /**
    * CONSTUCTOR: Create a new svt_ahb_master_monitor_def_toggle_cov_callback instance.
    */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new(svt_ahb_master_configuration cfg, MONITOR_MP monitor_mp, string name = "svt_ahb_master_monitor_def_toggle_cov_callback");
`elsif SVT_OVM_TECHNOLOGY
  extern function new(svt_ahb_master_configuration cfg, MONITOR_MP monitor_mp, string name = "svt_ahb_master_monitor_def_toggle_cov_callback");
`else
  extern function new(svt_ahb_master_configuration cfg, MONITOR_MP monitor_mp);
`endif

endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
b++dmB4WKAAKfezI+5Pt3PBUyOCcfbJCh85ZGMSP/FZ6Bn53XyUI00Nspb00+vQ0
SscByOAda5aSe5gbcNecVWW2vSvmpTs3N44/FUqtBP9s/aMpJXDPNjxya2fsMyT3
NxwmTCtlFaO2tAKgB6jTuKzchAugpaZcZuiGm1ngZeLszF175OP1zA==
//pragma protect end_key_block
//pragma protect digest_block
VuUZow6Gig6SzSJuoTWTUIrXBXY=
//pragma protect end_digest_block
//pragma protect data_block
AFa6Y8spgv7fXgo0KJMaKJ86qQDVecd51QFa6PFRgZfe7E5NjQT3m/P+vosRit1k
TAewmmleVoHgTCC63ayK8o+6JFU2n4L3KFwhXE/cMqnjDe/9y9TcpVmUH9TsyK29
1d9K///A2EXq7yvy3hLtPos24iiSMdymmwrzKPMmB0eZbEOJPQ8a0H24uxuVNiZO
meJOQj9vDWg9NUxVI9wu+MiSk/rc7+zjxKceIkUE+as/uiL0XxFkuHdCXNbf+wzU
EjJtRmV+TcFChMbw3Bha1Oq6xN34Fn3oaCi61w9BLJ/sTV8hLsnWlF0xAojwmFSX
hj6h8RvnirPoIFuyYhh898k6CNUa4AmZQwEAO1pq5cwTXasXdemCkBOtWf9lWm6F
lp9RlQAJPRN1OzyBveMf54BdIuKgs5KJSGzqPobR3rfPdi8Ufn7IrQ4UCpt1S6nZ
5auXulvK2KRPi2P9ocyHYkLIoXPjyMV78y46P4+Mb4dlw4NlNMh8XRF+UrFowprP
KTd0FgLIxvW6hnYc+vhtH10z7rNocySRUjXkXtqU8Rh7L/p3hqJG0d+B3ASwHWGE
h6Le9GddABHyx2X1ClKtYL/doSP9lg6H1ClHc/FXvXHLNdP+plzPuMozDCpMvH7L
ZHQUP0xYsPClytrVnCi/Ks90gi+7c/6mQULZL5AHlKsxT1dZn/FBhHEuDAbywbhW
WwElHZ37QDOvsuNSDsOkn8CdPLM1UgwkYboIub9GvONIK3mnPgBfzcSgz+gmiSIK
4RKmDx8LaW4+FApTt3v0ZWzcEzg98EOD5A/6i2KxN0SZjTguG+dENUIh4WAM9ovL
Jh5xY2GJvQ6r3X1cfOCbbSeYSYbx/pX0HlE3W/YjgCSHD9dFy+6cyj+RodP3IBY/
rPis2ccsC+u8QvMrDX8UYVv49PGOXC6P0axUy92QBKpD9QqU/Y/oGS6AN7MP5Yow
FhiMv1nFOnIFp8SaUqOFyoULO+29/880EL6cve5RJrTB2pvA5Rp/p0RTR4sfJ8e6
V31SZz1CYd0sdaviYo1jsVuYSci1VGbxspq2EJQiHt2rG54A2846veDBmUJWmv5/
MozyvkeJ2JU2yFYfi8qyedFU1eJXjfTHF0ZjYAmtd2AEXj9u/Hrc8i8+QJ4dcdAa
kRxOEcwp/3vm0pOYNWdBJeot1ficvVvimPW2Fzl4RDkaecTP6+PlAjBBvY7WCGta
PWHDefUZAqUObOeXyZZGR6Upzf59wj1crd0fqD3No+LcotiRHENXhch9/jl1va0g
fx3K/b/SXn2UvjaviyZZhJur7Pafoya/hEE9Ksh7m4xYPMvfG3LGAhgLDUEUONVF
Bvy7MiIu5UkqQtw7iMF5WWonV9OqZQXZx/jL4iR1NA1RwvzA1PDL3jQHwQb+7J2p
8fTc3zglHcmEnp7tmqIouuSmrsC1Dk2PjWetNJMN/AdECcsc5lQhcJdc+IUnhSsN
s/bNgVvdvgnWvNxYs6bhQ6e0n1mAb5wmmH/KWL5JeH1ttkUMGoomlH76w4H4JLBs
IqJskCQKiXGuvtfYee+oYop6/rWS66fpD+d8ovNoJbjlGT70yGJtFb8SzTl7zNl1
ukjvSV6dOjOuPVUrActTyi5wCIaxnQIwzts0ewXFREbLM3wcRkTokeT4+jihnwQG
HLxhjrQuT3LsKMiGa0W+c/Uibmy+PIRxSE4ceHOWNTKvLoIzpc3wpG/MvBSl+pQm
XJS7ZiS9alvLfIHqcvWeilosYNpHW5A33u5zzhCI3JzPjZVY1DfPt/y9eS2HIHOo
3jw+V/wRmv3qZx+oOB/EvUcdvUTHJThA7KPIkBP+8wg4YpfahsimegWCOkap5x07
jmqITNwZAajlB5fJ17Hte6m1Y6VcHN6U3Y0hPnTeWwwWQLfuebFQsqQmtmV4rL+B
tqmt63gbchUBHo65Bvw+RnR59a6gjQB8uoqPPIHxhocxUWN16TVHnOa+RmMmZ4bR
0YtFTTJjaLQnziXRG2fmG0RLkZqIbpSvEkLbwKZtVNTh2t68BYip+2oHx9I+vGgd
GEqK80SGd+3G83ZiDPrMOGeTzCHl0wG5WOjJAkj/65gj5vP7h9FBCYdPFqox/c5w
KxSgNe26bChYfxFTtg6GSTeNGf9P/EBv3h6rkwuSsCuOZe4wEOLiNzjTWCYbKdf+
KNeIf1AMspWc3nckvfPyfXHO+wV5L7aFVKXKR4aMNxJgAwbC1kVsqzxdXwCGesBk
gPbOVn2mCkvElKp7tz06zIwrGlPkSrks2oKHH8KV5PGxzdbKi8dWHSEl0bUmASRU
xAbKbUU/pInvLKXGzsk8Qi7eQgLeE4xav6G2plnLuOLuOooU0LY8AZTxMbYF5hHG
iV5KwxpwMp4wQv2FAnJwbzoKEPqqWKIIDW4dCo6NOlCbDuWpVNlhNcCliSMm8eQW
t5Ws1g4nYU+VewXcYL4MYL/qxdWi/mg2DA+oYz5emdY4lw+ITutz85KD2j3pHEmC
jSP20FfeZY32aN5Ds0+kX5Ar72DlKuYmb7v/aC47SSp82Ie6llNBTR4XSKnfrJ18
rPIqjbKrDWZOEpj+3o5HbIh+iK1cd4gXQLVsuQ9gBY3KfuYrGlZPCBvB0wvSfVHI
a2/+/EcCiV/kzD7sDQ9Wpx1+G7grl7Ypds5ckrcg1ko1yZa5qtxst4HAQOH7ZSrV
tJ6aQ6L5+r9x6KdFx/7y6BXbxvsAzGQUrjEuFZTYGkBB9MoZyMg8prWX1isr1nxU
B2orZeEHHpQwK7T38Dx2S5Gwdaw/8W5KuKmJWCvyFiNfyc32xKGJnakloWf8SpJU
stTIHkCCd6w6EybrD5kvQYPsUZFeVg21gDqQSNRxl2F7WawV+QFXrimCmOZaI9zQ
k6FuQ5LJh4s6kXlQsx5lRgXk1UJDIl5kVt9CxYtfFo2OHmHX9Lk7S3oxsxibjnzA
luFRARvnZlhPjJieABtw036tOiaxo4S3bI8lANXf9/+DgYBq5QM1EbZ664oOxYmy
+49E+GzdHEpoUz0/XQsDvovcRlL1kgORtxqbJYTjNIKMPZ6+kmKPWM73JMsixhvK
/tpU1cLmGdYtMJa68sexbtzgzYMgkNWDnnl7LGSVVGR718ApsY46fIrh8ge602nm
lPv79af3zn7/wJ4LjpWxffp2/mw7PzdzUVL3f8ZD/m1m7MurQUh2T09gk/novG1r
XpLLO8LaVU4bcbTmeDUDH36gj4RW77AU70toqsBBp5g=
//pragma protect end_data_block
//pragma protect digest_block
FhPZCAjQEVTy1XXiHr3ElWgbnJM=
//pragma protect end_digest_block
//pragma protect end_protected

`endif
