

`ifndef GUARD_SVT_AXI_PORT_CONFIGURATION_SV
`define GUARD_SVT_AXI_PORT_CONFIGURATION_SV

`include "svt_axi_defines.svi"

typedef class svt_axi_system_configuration;
typedef class svt_axi_system_domain_item;
typedef class svt_axi_slave_addr_range;
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RcsFmdXhjPUVOPCL2RirC+i/vGu8afqocHlfNMpvA2J6exZ8ASvELYr8la0vTVww
6mpFlUvmDLdc7J7jeY6ff5NuESapAFWswASKFuI/M4YeBLqegKUiFRYaBxL77Qky
ljQFUX464WA3g+qYviva7AfN66SmxSMm6CHwJ2AhS9A=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1006      )
9DKCZWzEHu9B6KbAVVRfCCNB6Yw7wSGEs2HpHmycZibfaukKuYWBQnZ6NgNXJ3N9
GvsbKI+st2xERrdu0sMZLceSjiW8CytbO/5EdP57xBlyLtOdsLTKOPsuXL9/CBxq
X6TTExa4utfhaHu9T08qfC2NTSIHik8bJlD/TfFxIGYB9qJklcXuMVKKErd+ZU0f
t1Kt0YAtOycsrzeBq07qBGGCfGDzoSXty0G1S5iEQtq/jwBW1yWBf8A7bYWpsG5K
QTMGQaE3RjC/zp+3WWIrlE527DsdgCRioS9phv0LGonjnBjmtuVeyyzEJpIBMlJZ
bGryBMAAbrc/JVToU8Sr5GSy+meUB/y3XFSL9ukOngrDQms6MS6pEKW5EZGC/ict
BtGdlXTzLDVu132agdNImV+GxsZh01BdHJv5I7zr/79lxs+jDGpKtlNS/yIyoUwq
stkgxTn1Y4bWnTuXxiVx7shSGEqLkPR+97hr0HBldueNuMnmoilGWwIiYH/Jw/Xh
cakgdmpn5BNj16So6AVprbiASmYVBXPEscFOaMeQ56daS5ZtXNahWvE1RXdgUxwx
bFpqi0iEx/yf8Lr8S0/bgCiGmtliW7k4m05Ifv3uPxYFPhfwHyL/ddrK7l181gOm
ZlsoY5FNMZ/PZotAAYkFXcEuc83xIPKhfY7U/8PUjOZCglEZ2RGiJXt3NUA4wTjI
dg1yYUgVDH7DsldZmn+2VDKS//ROvpkEqwtUUSknEXiPA3H5915hOhz+QCdibwrE
w0SwQ8lPEm5yW+5p65B2KOMybxYivAVL8NnbkssOO5wSw6DBQMymHMISpyiRAnpK
EPLsDKZFw0kY26BWYTOo7Hhj47ClxBGRBDUFeV9VVrDsPn4VNRx76W1qANef//+/
7uWGGbgQBc5saPsKOFkJ4XmZ/qGGzB5QUvSCr7sR2uMQ+ZO7vpiLiirNVQ7F3um8
IHmzJp1/4y4RzyStAhDC2mdElcfrmgzAU/2qm+6ZKP0dsPfSKA4ZBcgf/miqtoxM
+m/V/GHLrRl4cDc/1jbTTaG3bt6woVKDlgVC9f+fd+AIdUHiM5yv1SoOrvG9PHe7
H9aywUrN1NzMSs2tn8Y8vETtt8vN6w51sHiCDE8GAvNv1coc5P6OiPUu/wSnxhDr
/+cN7tsSTImtCRd80cHJWepAO8DvHjqP6cuHkhlNUFe+xGDS/7i4X4XkdUh/pw2s
+dxrsK/Iew+3zWsuCuUPA1ByBUDLrb+MaVGIgTjXGa+Z9pD2Muh7FqGjEUVIgJeE
iteO/RdxfroIxZDAUIJohaXENf30+yFuH5ZX1OUSqQm2qR+sS58LIUknayo8kbEB
`pragma protect end_protected

/**
    Port configuration class contains configuration information which is
    applicable to individual AXI master or slave components in the system component.
    Some of the important information provided by port configuration class is:
    - Active/Passive mode of the master/slave component 
    - Enable/disable protocol checks 
    - Enable/disable port level coverage 
    - Interface type (AXI3/AXI4/AXI4 Lite/AXI_ACE) 
    - Port configuration contains the virtual interface for the port
    .

  */
class svt_axi_port_configuration extends svt_configuration;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  /** Custom type definition for virtual AXI interface */
`ifndef __SVDOC__
`ifdef SVT_AXI_SVC_SINGLE_INTERFACE
  typedef virtual svt_axi_port_if AXI_MASTER_IF;
  typedef virtual svt_axi_port_if AXI_SLAVE_IF;
`else
  typedef virtual svt_axi_master_if AXI_MASTER_IF;
  typedef virtual svt_axi_slave_if AXI_SLAVE_IF;
`endif // __SVDOC__
  typedef virtual svt_axi_stream_if AXI_PORT_STREAM_IF;
`endif
  
  /**
    @grouphdr axi_generic_config Generic configuration parameters
    This group contains generic attributes which are used across all protocols
    */

  /**
    @grouphdr axi3_4_config AXI3 and AXI4 configuration parameters
    This group contains attributes which are specific to AXI3 and AXI4 protocol
    */

  /**
    @grouphdr axi3_4_timeout_config Timeout values for AXI3 and AXI4
    This group contains attributes which are used to configure timeout values for AXI3 and AXI4 signals and transactions
    */

  /**
    @grouphdr ace_config ACE configuration parameters
    This group contains attributes which are specific to ACE protocol
    */
  
   /**
    @grouphdr ace5_config ACE5 configuration parameters
    This group contains attributes which are specific to ACE5 protocol 
    ARM-EPM-033524 Version 2.0
    */

  /**
    @grouphdr axi_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable coverage and protocol checks
    */

  /**
    @grouphdr axi_signal_idle_value Signal idle value configuration parameters
    This group contains attributes which are used to configure idle values of signals (except "Ready" signals) when "Valid" is low.
    */

  /**
    @grouphdr default_ready Default "Ready" signal value configuration parameters
    This group contains attributes which are specific to ACE protocol
    */

  /**
    @grouphdr axi3_signal_width AXI3 signal width configuration parameters
    This group contains attributes which are used to configure signal width of AXI3 signals
    */

  /**
    @grouphdr axi4_signal_width AXI4 signal width configuration parameters
    This group contains attributes which are used to configure signal width of AXI4 signals
    */

  /**
    @grouphdr ace_signal_width ACE signal width configuration parameters
    This group contains attributes which are used to configure signal width of ACE signals
    */

  /**
    @grouphdr axi4_stream_signal_width AXI4 Stream signal width configuration parameters
    This group contains attributes which are used to configure signal width of AXI4 Stream signals
    */

  /**
    @grouphdr master_slave_xact_association Configuration parameters required for master and slave transactions association
    This group contains attributes which are used to associate master transactions to slave transactions 
    */

  `ifdef SVT_VMM_TECHNOLOGY
  /**
    @grouphdr axi3_4_generator AXI3 and AXI4 generator configuration parameters
    This group contains attributes which are used to configure stimulus and response generators for AXI3 and AXI4
    */

  /**
    @grouphdr ace_generator ACE generator configuration parameters
    This group contains attributes which are used to configure stimulus and response generators for ACE
    */
  `endif

  /**
    @grouphdr protocol_analyzer Protocol Analyzer configuration parameters
    This group contains attributes which are used to enable and disable XML file generation for Protocol Analyzer
    */

  /**
    @grouphdr axi_performance_analysis Performance Analysis configuration parameters
    This group contains attributes which are used to monitor performance of a
    system based on measurement of latencies, throughput etc. The user sets the
    performance constraints through performance analysis configuration
    parameters and the VIP reports any violations on these constraints. The time
    unit for all these parameters is the simulation time unit. Performance
    metrics that involve aggregation of values over a time period are measured
    over time intervals specified using configuration parameter
    perf_recording_interval. Measurement of other performance parameters that do
    not require aggregation of values over a time period are not affected by
    this configuration parameter. VIP reports statistics for each performance
    metric for each time interval. Each performance parameter can be enabled or
    disabled at any time.  Monitoring of a performance parameter is disabled by
    passing a value of -1 to the parameter. Passing any other value enables the
    performance parameter for measurement. If a value other than -1 is supplied,
    it will take effect at the next time interval. If the performance
    configuration parameter values are changed during simulation, the new
    configuration will need to be passed to the VIP using the #reconfigure()
    method of the top level VIP component, for eg. #reconfigure() method of AXI
    System Env will need to be called if AXI system Env is used as top level
    component.
    */

  /**
    @grouphdr axi_qvn_config AXI QVN Configuration parameters
    This group contains attributes which are used to configure QVN features in a
    system.
    */

  /**
    @grouphdr axi_tlm_generic_payload TLM Generic Payload parameters
    This group contains attributes which are used to support TLM Generic Payload feature.
    */

  /**
    @grouphdr axi_traffic_profile Traffic profile related parameters
    This group contains attributes which are used to support traffic profiles.
    */

  /**
    * Enumerated type to specify idle state of signals. 
    */
  typedef enum {
    INACTIVE_CHAN_LOW_VAL  = `SVT_AXI_INACTIVE_CHAN_LOW_VAL,    /**< Signal is
    driven to 0. For multi-bit signals each bit is driven to 0. */ 
    INACTIVE_CHAN_HIGH_VAL = `SVT_AXI_INACTIVE_CHAN_HIGH_VAL,   /**< Signal is
    driven to 1. For multi-bit signals each bit is driven to 1. */
    INACTIVE_CHAN_PREV_VAL = `SVT_AXI_INACTIVE_CHAN_PREV_VAL,   /**< Signal is
    driven to the previous value, ie, the value that it was driven to when the
    corresponding VALID signal was asserted. */
    INACTIVE_CHAN_X_VAL    = `SVT_AXI_INACTIVE_CHAN_X_VAL,      /**< Signal is
    driven to X. For multi-bit signals each bit is driven to X. */
    INACTIVE_CHAN_Z_VAL    = `SVT_AXI_INACTIVE_CHAN_Z_VAL,      /**< Signal is
    driven to Z. For multi-bit signals each bit is driven to Z. */
    INACTIVE_CHAN_RAND_VAL = `SVT_AXI_INACTIVE_CHAN_RAND_VAL    /**< Signal is
    driven to a random value. */
  } idle_val_enum;

  /**
    * Enumerated type to specify inactive wdata bytes of signals. 
    */
  typedef enum {
    INACTIVE_WDATA_BYTE_LOW_VAL  = `SVT_AXI_INACTIVE_WDATA_BYTE_LOW_VAL,    /**< Signal is
    driven to 0. For multi-bit signals each bit is driven to 0. */ 
    INACTIVE_WDATA_BYTE_HIGH_VAL = `SVT_AXI_INACTIVE_WDATA_BYTE_HIGH_VAL,   /**< Signal is
    driven to 1. For multi-bit signals each bit is driven to 1. */
    INACTIVE_WDATA_BYTE_X_VAL    = `SVT_AXI_INACTIVE_WDATA_BYTE_X_VAL,      /**< Signal is
    driven to X. For multi-bit signals each bit is driven to X. */
    INACTIVE_WDATA_BYTE_Z_VAL    = `SVT_AXI_INACTIVE_WDATA_BYTE_Z_VAL,      /**< Signal is
    driven to Z. For multi-bit signals each bit is driven to Z. */
    INACTIVE_WDATA_BYTE_RAND_VAL = `SVT_AXI_INACTIVE_WDATA_BYTE_RAND_VAL,   /**< Signal is
    driven to a random value. */
    INACTIVE_WDATA_BYTE_UNCHANGED_VAL = `SVT_AXI_INACTIVE_WDATA_BYTE_UNCHANGED_VAL  /**<Signal is
    driven to initial value. */
  } wdata_val_enum;


  /** Enumerated types that identify the type of the AXI interface. */
  typedef enum {
    AXI3        = `SVT_AXI_INTERFACE_AXI3,
    AXI4        = `SVT_AXI_INTERFACE_AXI4,
    AXI4_LITE   = `SVT_AXI_INTERFACE_AXI4_LITE,
    AXI4_STREAM = `SVT_AXI_INTERFACE_AXI4_STREAM,
    AXI_ACE     = `SVT_AXI_INTERFACE_ACE,
    ACE_LITE    = `SVT_AXI_INTERFACE_ACE_LITE
  } axi_interface_type_enum;

  /** Enumerated types that identify the AXI interface category. */
  typedef enum {
     AXI_READ_WRITE = `SVT_AXI_READ_WRITE,
     AXI_READ_ONLY  = `SVT_AXI_READ_ONLY,
     AXI_WRITE_ONLY = `SVT_AXI_WRITE_ONLY
  } axi_interface_category_enum;

`ifdef SVT_ACE5_ENABLE

typedef enum {
  STANDARD = 0,
  BASIC = 1,
  NOT_SUPPORTED = 2 
 } mte_support_type_enum;

typedef enum {
  MPAM_9_1 = 0,
  MPAM_FALSE = 1
 } mpam_support_type_enum;

`endif
  /**
    * Enumerated typed for the port kind
    */
  typedef enum {
    AXI_MASTER = `SVT_AXI_MASTER,
    AXI_SLAVE  = `SVT_AXI_SLAVE,
    GP_MASTER = `SVT_AMBA_GP_MASTER,
    GP_SLAVE = `SVT_AMBA_GP_SLAVE
  } axi_port_kind_enum;

  /** @cond PRIVATE */
  /**
    * Enumerated type for the kind of inactivity period for throughput calculation
    */
  typedef enum {
    EXCLUDE_ALL = 0,
    EXCLUDE_BEGIN_END = 1
  } perf_inactivity_algorithm_type_enum;
  /** @endcond */

  /**
    * Enumerated type for enabling a particular version of ACE spec  
    */
  typedef enum {
     ACE_VERSION_1_0 = 0,
     ACE_VERSION_2_0 = 1
   } ace_version_enum;

  typedef enum {
    ALL_INTERFACE_TYPES = 0, /**< svt_axi_transaction::force_xact_to_cache_line_size 
    will be applicable for the agents that have the svt_axi_port_configuration::axi_interface_type set to AXI_ACE or ACE_LITE interface types. */
    AXI_ACE_ONLY = 1,        /**< svt_axi_transaction::force_xact_to_cache_line_size 
    will be applicable only for the agents that have the svt_axi_port_configuration::axi_interface_type set to AXI_ACE interface type. */ 
    ACE_LITE_ONLY = 2        /**< svt_axi_transaction::force_xact_to_cache_line_size 
    will be applicable only for the agents that have the svt_axi_port_configuration::axi_interface_type set to ACE_LITE interface type. */ 
  } force_xact_to_cache_line_size_interface_type_enum; 

  /** @cond PRIVATE */
  /**
    * Enumerated typed for the memory kind
    */
  typedef enum {
    SV_BASED_SVT_MEM = `SVT_SV_BASED_SVT_MEM,
    C_BASED_SVT_MEM = `SVT_C_BASED_SVT_MEM
  } mem_type_enum;
  /** @endcond */

  typedef enum {
    RECOMMENDED_CACHE_LINE_STATE_CHANGE = `SVT_AXI_RECOMMENDED_CACHE_LINE_STATE_CHANGE,
    LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE = `SVT_AXI_LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE,
    LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE = `SVT_AXI_LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE
  } axi_cache_line_state_change_type_enum;

  /**
   * Enumerated type that indicates the reordering algorithm 
   * used for ordering the transactions or responses.
   */
  typedef enum {
    ROUND_ROBIN     = `SVT_AXI_REORDERING_ROUND_ROBIN, /**< Transactions will be 
    processed in the order they are received. */
    RANDOM      = `SVT_AXI_REORDERING_RANDOM, /**< Transactions will be 
    processed in any random order, irrespective of the order they are received. */
    PRIORITIZED = `SVT_AXI_REORDERING_PRIORITIZED /**< Transactions will be
    processed in a prioritized order. The priority of a transaction is known from
    the svt_axi_transaction::reordering_priority attribute of that transaction. */
  } reordering_algorithm_enum;

  /**
   * Enumerated type that indicates how the reordering depth 
   * of transactions moves.
   * 
   * Example:
   * Consider the read data reordering depth of 2; R1, R2, R3 and R4 are the read
   * transactions to be responded. The behavior for different types reordering depth
   * is as follows:
   * - STATIC:
   *   Once both R1 and R2 are complete, then only the reordering depth moves:
   *   {R1, R2} -- to --> {R3, R4}
   * - MOVING:
   *   If any of the R1 or R2 is complete, then the reordering depth moves. Suppose
   *   that R2 is complete before R1. Then the reordering depth window moves as:
   *   {R1, R2} -- to --> {R1, R3}
   * .
   */
  typedef enum {
    STATIC         = `SVT_REORDERING_WINDOW_STATIC, /**< The reordering depth moves
    when all transactions within the current reordering depth are complete. */
    MOVING         = `SVT_REORDERING_WINDOW_MOVING /**< A new transaction is considered
    for access to send read data as part of the given reordering depth when any transaction
    within the current reordering depth is complete. */
  } reordering_window_enum;
  
 /**
  * Name of the master as used in path coverage
  * This field can also be used to specify master specific
  * slave address mapping. Refer to the documentation of
  * svt_amba_addr_mapper for more details
  */
  string source_requester_name; 

  /**
   * This queue will hold the names of all the slaves, including non-AXI slaves, 
   * to which an AXI master can communicate.
   */
   svt_amba_addr_mapper::path_cov_dest_names_enum path_cov_slave_names[$];

  /**
   * Enumerated types that tells ERROR response handling policy for AXI Master and Slave.
   */
  typedef enum {
    NO_ERROR = 0,/**< When set to NO_ERROR,vip should not report an error on receiving decerr or slverr response. */
    ERROR_ON_SLVERR = 1,/**< When set to ERROR_ON_SLVERR,vip should report an error only on receiving slverr response. */
    ERROR_ON_DECERR = 2,/**< When set to ERROR_ON_DECERR,vip should report an error only on receiving decerr response. */
    ERROR_ON_BOTH = 3 /**< When set to ERROR_ON_BOTH,vip should report an error on receiving decerr or slverr response. */
  } error_response_policy_enum;

  /**
   * Enumerated type that defines the behaviour of the VIP during reset
   */
  typedef enum { 
    EXCLUDE_UNSTARTED_XACT = `SVT_AXI_EXCLUDE_UNSTARTED_XACT, /**< Only those transactions which have gone out on the interface are ABORTED. */
    RESET_ALL_XACT = `SVT_AXI_RESET_ALL_XACT /**< All transactions which have already started along with the ones which have not yet started but are present in the internal queue are ABORTED. */
  } reset_type_enum;

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * Enumerated type that defines the generator source for slave responses
   */
  typedef enum { 
    NO_SOURCE    = `SVT_AXI_NO_SOURCE,           /**< No internal source. This generator_type is used by master component. This specifies that no internal source should be used, and user is expected to drive the master driver input channel. */
    ATOMIC_GEN   = `SVT_AXI_ATOMIC_GEN_SOURCE,   /**< Create an atomic generator. This generator_type is used by master component. This specifies the master component to use atomic generator. */
    SCENARIO_GEN = `SVT_AXI_SCENARIO_GEN_SOURCE,  /**< Create a scenario generator. This generator_type is used by master component. This specifies the master component to use scenario generator. */
    SIMPLE_RESPONSE_GEN = `SVT_AXI_SIMPLE_RESPONSE_GEN_SOURCE, /**< This generator_type is used by slave component. When this generator_type is specified, a callback of type svt_axi_slave_response_gen_simple_callback is automatically registered with the slave response generator. This callback generates random response. */
    MEMORY_RESPONSE_GEN = `SVT_AXI_MEMORY_RESPONSE_GEN_SOURCE, /**< This generator_type is used by slave component. When this generator_type is specified, a callback of type svt_axi_slave_response_gen_memory_callback is automatically registered with the slave response generator. This callback generates random response. In addition, this callback also reads data from slave built-in memory for read transactions, and writes data into slave built-in memory for write transactions. */
    USER_RESPONSE_GEN = `SVT_AXI_USER_RESPONSE_GEN_SOURCE /**< This generator_type is used by slave component. When this generator_type is specified, slave response callback is not automatically registered with the slave component. The user is expected to extend from svt_axi_slave_response_gen_callback, implement the generate_response callback method, and register the callback with the slave response generator. */
  } generator_type_enum;

  /**
   * Enumerated type that defines the generator source for snoop responses
   */
  typedef enum { 
    CACHE_SNOOP_RESPONSE_GEN = `SVT_AXI_CACHE_SNOOP_RESPONSE_GEN_SOURCE, /**< This generator_type is used by master component, when the #axi_interface_type is AXI_ACE. When this generator_type is specified, a callback of type #svt_axi_master_snoop_response_gen_cache_callback is automatically registered with the master component. This callback generates random snoop response based on the cache line status. */
    USER_SNOOP_RESPONSE_GEN = `SVT_AXI_USER_SNOOP_RESPONSE_GEN_SOURCE /**< This generator_type is used by master component. When this generator_type is specified, snoop response callback is not automatically registered with the master component. The user is expected to extend from #svt_axi_master_snoop_response_gen_callback, implement the generate_snoop_response callback method, and register the callback with the snoop response generator. */
  } snoop_response_generator_type_enum;

  /**
   * Enumerated type that defines the barrier transaction association approach
   */
  typedef enum { 
    RANDOM_ASSOCIATION = `SVT_AXI_RANDOM_BARRIER_XACT_ASSOCIATION, /**< This approach type is used by master component, when the #axi_interface_type is AXI_ACE. When this approach is specified, a callback of type #associate_xact_with_barrier_pair_xact() is automatically registered with the master component. This callback associates barrier transaction with normal coherent transaction in a random manner. */
    USER_DEFINED_ASSOCIATION = `SVT_AXI_USER_DEFINED_BARRIER_XACT_ASSOCIATION /**< This approach type is used by master component. When this approach is specified, the callback is not automatically registered with the master component. The user is expected to extend from
#associate_xact_with_barrier_pair_xact, implement the association of barrier transaction with normal coherent transaction */
  } barrier_association_type_enum;

  /**
   * Enumerated type that defines the generator source for DVM complete transactions
   */
  typedef enum { 
    AUTO_DVM_COMPLETE_GEN = `SVT_AXI_AUTO_DVM_COMPLETE_GEN_SOURCE, /**< This generator_type is used by master component, when the #axi_interface_type is AXI_ACE. When this generator_type is specified, master automatically generates a DVM Complete transaction, after receiving a DVM Sync transaction. The delay between reception of DVM Sync and transmission of DVM Complete is determined by random member dvm_complete_delay*/
    USER_DVM_COMPLETE_GEN = `SVT_AXI_USER_DVM_COMPLETE_GEN_SOURCE /**< This generator_type is used by master component. When this generator_type is specified, user will need implement callback method svt_axi_master_snoop_response_gen_callback::dvm_complete_gen. The user can program the delay  dvm_complete_delay in the callback method. */
  } dvm_complete_generator_type_enum;

`endif

  /**
   * Enumerated type that defines the snoop response mode during memory update transactions
   */
  typedef enum { 
    SUSPEND_SNOOP_DURING_MEM_UPDATE = 0, /**< Master suspends incoming snoop request if memory update transaction is found in the buffer, or is active at the time of receiving snoop request and provides response to that snoop request only after the current ongoing memory update transaction is complete */
    SUSPEND_SNOOP_DURING_MEM_UPDATE_IN_PROGRESS = 1, /**< Master suspends incoming snoop request if memory update transaction is found to be active (addres/data phase started or about to start in current clock) at the time of receiving snoop request and provides response to that snoop request only after the current ongoing memory update transaction is complete */
    RESPOND_SNOOP_DURING_MEM_UPDATE = 2, /**< Master doesn't suspend incoming snoop request even if memory update transaction is found to be active at the time of receiving snoop request. Instead it responds to the snoop request with allowed snoop response while memory update transaction is in progress.*/ 
    EITHER_RESPOND_OR_SUSPEND_SNOOP_DURING_MEM_UPDATE = 3  /**< Master either suspends incoming snoop request or respond to the snoop request while memory update transaction is in progress in a random manner.*/ 
  } snoop_response_mode_during_mem_update_type_enum;

  /**
    * 
    */
  typedef enum {
    SNOOP_RESP_DATA_TRANSFER_USING_CDDATA = `SVT_AXI_SNOOP_RESP_DATA_TRANSFER_USING_CDDATA, /**<Transfers cache data of dirty line using CDDATA channel */
    SNOOP_RESP_DATA_TRANSFER_USING_WB_WC = `SVT_AXI_SNOOP_RESP_DATA_TRANSFER_USING_WB_WC /**<Transfers cache data of dirty line using WRITEBACK or WRITECLEAN */
  } snoop_response_data_transfer_mode_enum;

  /** enum description for various address randomization mode for nonshareable transaction with domain type SYSTEMSHAREABLE */
  typedef enum {
    NONSHAREABLE_XACT_FULL_ADDRESS_SPACE = 0, /**<allows full address sapce to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
    NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE = 1, /**<allows only address sapce outside inner, outer or nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
    NONSHAREABLE_XACT_ADDR_WITHIN_NON_SHAREABLE_ADDR_RANGE = 2, /**<allows only nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
    NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_ADDR_RANGE = 3 /**<allows only address sapce outside inner or outer address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
  } nonshareable_xact_address_range_in_systemshareable_mode_enum;
  typedef enum {
    STATIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES = 0,
    DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES = 1,
    CUSTOM_SOURCE_MASTER_ID_XMIT_TO_SLAVES = 2 
  } source_master_id_xmit_to_slaves_type_enum;

  typedef enum {
    FALSE = 0,
    ODD_PARITY_BYTE_DATA = 1,
    ODD_PARITY_BYTE_ALL = 2
  } check_type_enum;

  /**
   * Enumerated type that defines the modifiable and non modifiable cache types
   */
  typedef enum {
    SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_NONMODIFIABLE_CHECK = 0,
    SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_MODIFIABLE_NONMODIFIABLE_CACHE_TYPE_CHECK = 1,
    SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_DISABLE_CHECK = 2
  } master_slave_xact_association_cache_prot_check_enum;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************
`ifndef __SVDOC__
  /** Port interface */
  AXI_MASTER_IF master_if;
  AXI_SLAVE_IF slave_if;
  AXI_PORT_STREAM_IF port_stream_if;
`endif

  /** 
    * @groupname axi_generic_config
    * A unique ID assigned to the master/slave port corresponding
    * to this port configuration. This ID must be unique across
    * all masters/slaves of the AXI system configuration to which
    * this port belongs. A master and a slave may share the same
    * port_id, but two masters or two slaves cannot share the 
    * same port_id. If not assigned by the user, it is auto
    * assigned by the VIP. 
    */ 
  int port_id;

  /** @cond PRIVATE */
  /**
    * @groupname axi_generic_config
    * Name of this port. This is used in transaction short display
    * to identify the instance. This is copied over from 'inst'
    * attribute.  
    */
 local string port_name;
  /** @endcond */
  /** 
    * @groupname axi_generic_config
    * A unique ID assigned to master/slave port corresponding to this port
    * configuration. This ID must be unique across all AMBA components
    * instantiated in the testbench.  This is currently applicable only when the AMBA
    * system monitor is used and is configured using a configuration plain text
    * file (as opposed to a SystemVerilog code that sets the configuration). 
    */
  int amba_system_port_id = -1;

  /** 
    * @groupname axi_generic_config 
    * Specifies whether output signals from master/slave IFs should be
    * initialized to 0 asynchronously at 0 simulation time. 
    * - 1: Intializes output signals from master/slave IFs to 0 
    *      asynchronously at 0 simulation time.
    * - 0: Initializes output signals from master/slave IFs to Z
    *      synchronously at 0 simulation time.
    * .
    * Configuration type: Static <br>
    * Default value: 0 <br>
    */ 
  bit initialize_output_signals_at_start = 1'b0;

  /** 
    * @groupname axi_generic_config 
    * Specifies whether clock should be disconnected to this agent. 
    * - 1: clock will be connected to this agent from the testbench, 
    *      based on the svt_axi_system_configuration::common_clock_mode.
    * - 0: clock will not be connected to this agent from the testbench.
    *      Used to disable the agent as per the test requirement.
    * .
    * Configuration type: Static <br>
    * Default value: 0 <br>
    */ 
  bit clock_enable = 1'b1;

  /**
    * @groupname axi_generic_config
    * Handle to the system configuration object
    */
  svt_axi_system_configuration sys_cfg;

  /**
    * @groupname axi_addr_map
    * Applicable only to slave VIP
    * Address map for this slave 
    * Must be used only if the svt_axi_system_env and svt_axi_system_configuration is not used.
    * Typically used in an environment where only one slave VIP is instantiated.
    */
  svt_axi_slave_addr_range slave_addr_ranges[];

  /**
    * @groupname axi_addr_map
    * Address map that maps global address to a local address at destination
    * Typically applicable to slave components
    * Applicable only if svt_axi_system_configuration::enable_complex_memory_map is set
    */
  svt_amba_addr_mapper dest_addr_mappers[];

  /**
    * @groupname axi_addr_map
    * Address map that maps a local address to a global address at a source
    * Typically applicable to master components. However, it can be applicable to
    * a slave component if that is connected downstream through another interconnect/bridge to
    * components which are further downstream. Applicable only if
    * svt_axi_system_configuration::enable_complex_memory_map is set
    */
  svt_amba_addr_mapper source_addr_mappers[];

  /**
    * @groupname axi_generic_config
    * Indicates if WID must be driven for AXI4, AXI_ACE,ACE_LITE,AXI4_LITE interfaces 
    * Configuration type: Static
    * Applicable only to MASTER 
    */

    bit  wid_for_non_axi3_enable = 0;

  /** 
    * @groupname axi_generic_config
    * Field for updating slave memory in request order
    * When set to 1, updates slave memory in request order that is  even though response
    * is received out of order, memory will still be updated in request order at the last
    * data phase. 
    * Default value is 0.
    * Configuration type: Static
    * Applicable only to SLAVE
    */ 
    int update_memory_in_request_order = 0;

    /**
    * @groupname axi_generic_config
    * Indicates that the monitor will check that recommended number of transactions are used      in the locked sequence 
    * Configuration type: Static
    * Applicable only to MASTER 
    */

    bit check_recommended_xact_length_for_locked_sequence = 0;
   
    /**
      * @groupname axi_generic_config
      * Indicates if X/Z checks and signal stability checks must be enabled
      * These are low level checks performed every clock and have a performance overhead
      * Often, these checks are useful only during integration phase. These can be
      * switched off after integration to get better performance.
      * These checks are automatically disabled if SVT_AXI3_4_PERF_MODE is set
      */
    bit per_clock_cycle_signal_checks_enable = 1;
 

  /**
    * @groupname axi_generic_config
    * If set to svt_axi_port_configuration::RESET_ALL_XACT,all transactions which have
    * already started along with the ones which have not yet started but are
    * present in the internal queue are ABORTED.
    * If set to svt_axi_port_configuration::EXCLUDE_UNSTARTED_XACT,only those transactions
    * which have gone out on the interface will be ABORTED.
    * Configuration type: Static
    *
    * This is applicable to only the Master in active mode because in passive mode
    * or for the slave all transactions which are in the queue are already started
    */
    reset_type_enum reset_type = `SVT_AXI_RESET_TYPE;


  /**
   * @groupname axi3_4_config
   * Indicates the way VIP reports error on receiving SLVERR or DECERR read or write response.
   * If set to svt_axi_port_configuration::NO_ERROR,vip doesn't report any error on receiving decerr
   * or slverr response.
   * If set to svt_axi_port_configuration::ERROR_ON_SLVERR,vip reports error only on receiving 
   * slverr response.
   * If set to svt_axi_port_configuration::ERROR_ON_DECERR,vip reports error only on receiving 
   * decerr response.
   * If set to svt_axi_port_configuration::ERROR_ON_BOTH,vip reports error on receiving 
   * decerr or slverr response.
   * Configuration type: Static
   *
   * This is applicable to Master in both active and passive mode and to slave only in Passive mode.
   * The default enum type of error_response_policy is NO_ERROR and is user configurable.
   */
   error_response_policy_enum error_response_policy = NO_ERROR;


  /**
    * @groupname axi_generic_config
    * Indicates if VIP would use separate address spaces for each tagged attribute. This simply means that,
    * if a coherent master or interconnect or a slave attached to such system, recieves both secure and non-secure
    * transactions then both transactions will operate on completely separate address spaces and result of one transaction
    * will not be visible to the other.
    *
    * Slave for which separate secure & non-secure address space is enabled i.e. bit [0] is set to '1', it will accept both secure
    * and non-secure transactions targeted for the same address. However, while updating memory it will use tagged address i.e. 
    * address attribute, in this case security bit, will be appended to the original address as the MSB bits.
    *
    * Slave for which separate secure & non-secure address space is disabled i.e. bit [0] is set to '0' but, configured with secured
    * regions i.e. addr_attribute[0] is set to '1' in svt_axi_slave_addr_range class via task /#set_addr_range() in system configuration
    * then it will accept only secure transactions for secure regions and all transactions for non-secure regions. 
    * With this configuration slave will use orginal address while updating memory and will not use tagged address. Hence, secure and
    * non-secure transactions to the same address will affect each other, if targeted to non-secure regions. However, if it is targeted
    * to secure regions then only secure transations will be able to update memory and access for non-secure transactions will be declined as if address doesn't exist.
    *
    * Slaves can be configured with secure region by calling /#set_addr_range(<start_addr>,<end_addr>,<addres_attribute, ex: 1 [secured]>)
    *
    * [0] => represents separate address spaces for secure and non-secure attribute if set to '1'
    * [\`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:1] => RESERVED and should be set to 0
    *
    * Configuration type: Static
    * Applicable only to MASTER 
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE    
    bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0]  tagged_address_space_attributes_enable = 0;
`else    
    bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0]  tagged_address_space_attributes_enable = 1;
`endif    
    
  /**
    * @groupname axi_generic_config
    * If set to '0' then Master VIP will not drive overlapped coherent transactions on Read and Write
    * channel at the same time. WRITE transactions received by the sequencer will be blocked from being
    * sent on the interface if there is another READ transaction to an overlapping address which is 
    * already in progress. The same is true if a READ transaction is received from sequencer and a WRITE
    * transaction is in progress
    * Example: ReadShared started at 1000 ns and WriteBack received from sequencer at 1200 ns when 
    *          ReadShared is still active. At this point Master VIP will block WriteBack until ReadShared
    * is finished on the Read channel.
    *
    * If set to '1' then Master VIP will drive coherent transactions on Read and Write
    * channel as it receives from the sequencer as per other coherent rules. It will not
    * block as mentioned above. 
    * Certain scenarios that involve a store on the read channel sent out
    * speculatively while a WRITEBACK/WRITECLEAN to the same cacheline is in
    * progress require that this parameter is set to 0 so that cache states
    * reflect correctly. 
    * If snoop_response_data_transfer_mode is set to
    * SNOOP_RESP_DATA_TRANSFER_USING_WB_WC, this parameter must be set to 1 to
    * facilitate the transfer of snoop data on the write channel without
    * getting blocked.
    *
    * Configuration type: Static
    *
    * This is applicable to only the Master in active mode 
    */
    bit allow_overlapped_read_and_write_channel_coherent_transactions = 0;    
   
   /**
    * @groupname axi_generic_config
    * If set to '1' then Master VIP can drive random snoop response for
    * WasUnique (BRRESP[4]) even if the snoop_initial_cache_line_state is in 
    * UNIQUE state.
    * If set to '0' the Master VIP must set WasUnique (BRRESP[4]) to 1 if
    * the snoop_initial_cache_line_state is UNIQUE.
    */ 
    bit allow_was_unique_zero_in_unique_state = 1; 
   
   /** @cond PRIVATE */
  /**
    * @groupname axi_generic_config
    * If set to '1' then Master VIP will allow burst_size to be less than
    * data_width for Atomic transaction.
    * If set to '0' then Master VIP will throw an is_valid error when burst_size 
    * is less than data_width for Atomic transaction.
    * This is only applicable for multibeat atomic transactions. 
    */
    bit allow_multibeat_atomic_transactions_to_be_less_than_data_width = 0;   
    /** @endcond */

   /**
    * @groupname axi_generic_config
    * This is applicable only when interconnect VIP is used, this is
    * applicable for all transactions. 
    * So if set to 1, then the interconnect VIP will always update dirty data into main memory 
    * if it receives dirty data from snoops corresponding to a transaction from this port
    */
    bit memory_update_for_pass_dirty_enable = 0;
 
   /**
    * @groupname axi_generic_config
    * This is applicable only when interface_type is AXI3 or AXI4
    * If set to 1 and axi_interface_type is AXI3/AXI4, system monitor will update
    * the port_configuration member axi_interface_type as ACE_LITE .
    * In addition to that system monitor will update svt_axi_transaction::xact_type as COHERENT.
    */

    bit is_downstream_coherent = 1'b0;

  /** @cond PRIVATE */
  /** Helper attribute for specifying solve order */
  local rand bit primary_props;

  /** holds total number of enabled tagged address space attributes */
  local int      num_enabled_tagged_addr_attributes = 0;

  /** Supports four state memory
   *  Default value is set as 0
   *  If set as 1 supports 4 state memory.
   */

  bit is_4state = 1'b0;
  /** @endcond */


`ifdef SVT_VMM_TECHNOLOGY
  /** 
   * @groupname axi3_4_generator
   * The source for the stimulus that is connected to the transactor.
   *
   * Configuration type: Static
   */
  generator_type_enum generator_type = SCENARIO_GEN;

  /**
   * @groupname ace_generator
   * The source type for snoop response generation.
   *
   * Configuration type: Static
   */
  snoop_response_generator_type_enum snoop_response_generator_type = CACHE_SNOOP_RESPONSE_GEN;

  /**
   * @groupname ace_config
   * Defines how a transaction is associated with a barrier transaction pair.
   *
   * Configuration type: Static
   */
  barrier_association_type_enum barrier_association_type = RANDOM_ASSOCIATION;

  /** 
    * @groupname ace_generator
    * Defines how DVM complete transactions need to be generated.
    *
    * Configuration type: Static
    */
  dvm_complete_generator_type_enum dvm_complete_generator_type = AUTO_DVM_COMPLETE_GEN;

  /** 
    * @groupname axi_generic_config
    * The number of scenarios that the generators should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int stop_after_n_scenarios = -1;

  /**
    * @groupname axi_generic_config
    * The number of instances that the generators should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int stop_after_n_insts = -1;

  // ACE
  /** 
    * @groupname axi_generic_config
    * The number of scenarios that the snoop_generator should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int snoop_stop_after_n_scenarios = -1;

  /** 
    * @groupname axi_generic_config
    * The number of instances that the snoop generator should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int snoop_stop_after_n_insts = -1;

`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname axi_generic_config
    * When silent_mode is set to 1, the "Transaction started" and 
    * "Transaction ended" messages are printed in UVM_HIGH verbosity.
    * When silent_mode is set to 0, the "Transaction started" and 
    * "Transaction ended" messages are printed in UVM_LOW verbosity.
    */
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname axi_generic_config
    * When silent_mode is set to 1, the "Transaction started" and 
    * "Transaction ended" messages are printed in OVM_HIGH verbosity.
    * When silent_mode is set to 0, the "Transaction started" and 
    * "Transaction ended" messages are printed in OVM_LOW verbosity.
    */
`else
  /**
    * @groupname axi_generic_config
    * When silent_mode is set to 1, the "Transaction started" and 
    * "Transaction ended" messages are printed in DEBUG_SEV.
    * When silent_mode is set to 0, the "Transaction started" and 
    * "Transaction ended" messages are printed in NORMAL_SEV.
    */
`endif
  bit silent_mode  = 0;

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname axi_generic_config
    * Specifies if the agent is an active or passive component. Allowed values are:
    * - 1: Configures component in active mode. Enables sequencer, driver and
    * monitor in the the agent. 
    * - 0: Configures component in passive mode. Enables only the monitor in the agent.
    * - Configuration type: Static
    * .
    */
`elsif SVT_OVM_TECHNOLOGY
  /** 
    * @groupname axi_generic_config
    * Specifies if the agent is an active or passive component. Allowed values are:
    * - 1: Configures component in active mode. Enables sequencer, driver and 
    * monitor in the the agent. 
    * - 0: Configures component in passive mode. Enables only the monitor in the agent.
    * - Configuration type: Static
    * .
    */
`else
  /**
    * @groupname axi_generic_config
    * Specifies if the group is an active or passive component. Allowed values are:
    * - 1: Configures component in active mode. Enables driver, generator and
    * monitor in the group component. 
    * - 0: Configures component in passive mode. Enables only the monitor in the group component.
    * - Configuration type: Static
    * .
    */
`endif
  bit is_active = 1;
  
  /** @cond PRIVATE */
  /** xml_writer handle of the agent */
  svt_xml_writer xml_writer = null;
  /** @endcond */


  /** 
    * @groupname axi_generic_config
    * The AXI interface type that is being modelled. Please note that interface
    * type AXI_STREAM is not yet supported.
    * Configuration type: Static
    */
  rand axi_interface_type_enum axi_interface_type = AXI3;

  /** 
    * @groupname axi3_4_config
    * The AXI4 interface category (read-only, write-only, read-write) of this interface. 
    * Configuration type: Static
    */ 
  rand axi_interface_category_enum axi_interface_category = AXI_READ_WRITE;

  /**
    * @groupname axi_generic_config
    * Indicates whether this port is a master or a slave. User does not need to
    * configure this parameter. It is set by the VIP to reflect whether the port
    * represented by this configuration is of kind master or slave.
    */ 
  axi_port_kind_enum axi_port_kind = AXI_MASTER;

  /**
    * Specifies the impact of svt_axi_transaction::force_xact_to_cache_line_size 
    * based on the axi_interface_type. 
    * 
    * Applicable only for ACTIVE master.
    */
  force_xact_to_cache_line_size_interface_type_enum force_xact_to_cache_line_size_interface_type = ALL_INTERFACE_TYPES;

 /** 
   * @groupname ace5_config
   * Indicates supported version  of ACE specefication by AMBA AXI_ACE VIP
   * Default value of this parameter is ace_version_1_0.User need to set this parameter if they wish to
   * to use new ACE spec which is ACE spec version 2.0
   * Configuration type:static
   */
   ace_version_enum ace_version = ACE_VERSION_1_0;

/** 
   * @groupname ace5_config
   * Indicates cache stashing feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit cache_stashing_enable = 0;

/** 
   * @groupname ace5_config
   * Indicates if trace signal feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit trace_tag_enable = 0;

/** 
   * @groupname ace5_config
   * Indicates whether the trace tag value will be directly reflected in the response packet or spawned packets generated in response to the received packet.
   * when set to 1: The trace_tag value will be directly mapped to the associated response and spawned packets, irrespective of trace_tag value being 0 or 1 in the request.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0 and svt_axi_port_configuration::trace_tag_enable is set to 1.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit loopback_trace_tag_enable = 0;

`ifdef SVT_ACE5_ENABLE 
/** 
   * @groupname ace5_config
   * Indicates if atomic transactions feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit atomic_transactions_enable = 0;


 /** 
   * @groupname ace5_config
   * Indicates if write_with_cmo feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit write_plus_cmo_enable = 0;
 
 /** 
   * @groupname ace5_config
   * Indicates if cmo transactions can be sent on the write channel.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit cmo_on_write_enable = 0;

 /**@groupname ace5_config
   * Specifies the number of outstanding Atomic transactions a port can support.<br>
   * This is applicable only for ACE5 ports with atomic_transactions_enable set to 1.<br>
   * The Atomic transactions include:
   * - AtomicStore
   * - AtomicLoad
   * - AtomicSwap
   * - AtomicCompare
   * .
   * MASTER:
   * If the number of outstanding atomic transactions is equal to this
   * number, the slave will refrain from initiating any new 
   * transactions until the number of outstanding write transactions
   * is less than this parameter.<br>
   * SLAVE:
   * If the number of outstanding transactions is equal to 
   * this number, the slave will not assert ARREADY/AWREADY
   * until the number of outstanding transactions becomes less
   * than this parameter. 
   * <br>
   * This parameter must be set if #num_outstanding_xact = -1.
   * This parameter must not be set if #num_outstanding_xact is not set to -1.
   * - <b>Default val:</b> -1
   * - <b>min val:</b> 1
   * - <b>max val:</b> Value defined by macro \`SVT_AXI_MAX_NUM_OUTSTANDING_XACT.
   * - <b>type:</b> Static
   * .
   */
  rand int num_outstanding_atomic_xact = 1;

 /** 
   * @groupname ace5_config
   * Indicates if Memory Partitioning and Monitoring (MPAM) feature is supported.
   * It can be set to either of two values below:
   *    enable_mpam = svt_axi_port_configuration:FALSE
   *  When set to FALSE, MPAM is not supported on the interface.
   *    enable_mpam = svt_axi_port_configuration:MPAM_9_1
   *  When set to MPAM_9_1, MPAM is supported on the interface with mpam_partid_width=9 and mpam_perfmongroup_width=1. 
   *  Only applicable when SVT_ACE5_ENABLE macro is defined and svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
   * - Default value:FALSE, is controlled through user re-definable macro `SVT_AXI_PORT_CFG_DEFAULT_ENABLE_MPAM.
   * .
   */
   mpam_support_type_enum enable_mpam = `SVT_AXI_PORT_CFG_DEFAULT_ENABLE_MPAM;

 /** 
   * @groupname ace5_config
   * Indicates the width of MPAM Partition identifier.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   rand int mpam_partid_width = 9;

 /** 
   * @groupname ace5_config
   * Indicates the width of MPAM Performance monitor group.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   rand int mpam_perfmongroup_width = 1;

`endif
  /**
   * @groupname ace5_config
   * If set to 1, it will enable the master component to support deallocating transactions.
   * By default, the value of this parameter is 0. This means it can not support deallocating
   * transactions and any READONCEMAKEINVALID or READONCECLEANINVALID transaction initiated
   * from this master component will be converted to READONCE transaction.
   *
   * Applicable only when svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
   * and svt_axi_port_configuration::axi_interface_type is set to ACE_LITE
   * Configuration type:static
   */
   bit deallocating_xacts_enable = 0;



  /** 
   * @groupname ace5_config
   * Indicates address translation feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit addr_translation_enable = 0; 

  /**
    * @groupname axi_generic_config
    * Indicates whether this port is a interconnect VIP port or not. User does not need to
    * configure this parameter. It is set by the VIP to reflect whether the port
    * represented by this configuration is a port of interconnect VIP or not.
    * .
    */  
  bit is_ic_port = 0;
  
 /**
   * @groupname axi_generic_config
   * Indicates if the port_monitor protocol check max_num_outstanding_xacts_check 
   * is enabled or not .The max_num_outstanding_xacts_check checks that AXI master and AXI slave 
   * are not exceeding the user configured maximum number of outstanding transactions (#num_outstanding_xact).   
   * If #num_outstanding_xact = -1 then #num_outstanding_xact will not be considered , 
   * instead #num_read_outstanding_xact and #num_write_outstanding_xact will be considered for read and write transactions respectively.
   */
  bit max_num_outstanding_xacts_check_enable =0; 
 
  /** @groupname axi_generic_config
    * Disable the association between slave read transaction and master partial write transaction.
    * This covers the specefic scenario when master partial write transaction is split into
    * slave read transaction followed by a slave write transaction by the ICN.
    * If set to 1 association between master write transaction and slave read transaction is done by the system monitor.
    * If set to 0 association between master write transaction and slave read transaction is not done by the system monitor.
    */
  bit partial_write_to_slave_read_and_write_association_enable = 0;
 
 /**
   * @groupname axi_generic_config
   * Indicates if this port is interleaved based on address to be accessed by this port
   */
  bit port_interleaving_enable =0;  
 
/** Indicates the port interleaving boundary. The value must be in form of bytes.
  * For example if interleaving szie is 64 . It means interleaving boundary os 64 bytes.
  * This port will access address locations based on interleaving size.
  * Default value is set as 64.
  * Applicable if the port_interleaving_enable is set to 1 for this port.
  */
  int port_interleaving_size = 64;

/** Indicates the group id of all the ports participating in one interleaving scheme
  * All the ports which are in the same interleave group must be configured to have same 
  * port_interleave_group_id
  * Default is set to -1 . 
  * Applicable if the port_interleaving_enable is set to 1.
  * Its value must be unique across master and slaves .All the port_ids having same port_interleaving_group_id
  * must be contigous.
  */
  int port_interleaving_group_id = -1;

/** Indcates that DVM transactions will be sent form this port of corresponding port interleaving group
  * This port will not take part in port interleaving for DVM transactions 
  * Applicable if port_interleaving_enable is set to 1.
  */
  bit dvm_sent_from_interleaved_port = 0;

/**Indicates that non coherent device traffic will be sent from this port
  * of corresponding port interleaving group.
  * This port will not take part in port interleaving for device traffic
  * as Device transaction addresses are not interleaved.
  * Applicable only when the port_interleaving_enable is set to 1.
  */ 
  bit device_xact_sent_from_interleaved_port =0;

/**  Indicates the order of this port in a port interleaving scheme.
  *  For example : If the port is 3rd in a group of 4 ports .If port_interleaving_size of the group is 512 bytes
  *  This port will have access to addresses with addr[10:9] == 3.
  *  This parameter determines which address bits to look for an interleaved port.
  *  Default value of this is set to 0 
  */
   int port_interleaving_index = 0;

  /**
   * @groupname axi_generic_config
   * Enables port inteleaving for this port for the device type xact.
   * The port configuration parameter device_xact_sent_from_interleaved_port
   * is not applicable if this bit is set to 1.
   * If this bit is set to 1, the device type transaction is interleaved like 
   * any non-dvm transaction.
   */
  bit port_interleaving_for_device_xact_enable = 0;

  /**
    * Indicates if this port  supports the setting of Poison field. <br>
    * - Default value: 0.
    * .
    */
  bit poison_enable = 1'b0;

   /** 
    * @groupname axi_generic_config
    * Indicates if the transactions on this port must be processed by the axi
    * system monitor. This configuration is applicable only to the
    * 'system_monitor' of the instance of svt_axi_system_env within which the
    * component corresponding to this port configuration is instantiated.
    * It is not used in the AMBA system monitor instantiated in an instance of
    * svt_amba_system_env (system env used when multiple AMBA protocols are
    * used)
    */ 
  bit connect_to_axi_system_monitor = 1;

  /** @cond PRIVATE */
  /**
    * @groupname axi_generic_config
    * Indicates that, if this bit is set to '1' then user needs to externally push
    * coherent and snoop master transactions and slave transactions into the port monitors. 
    * port monitor will not automatically sample it's related interface and hence will not
    * create corresponding transactions and instead will use the user provided transaction handle
    * externally pushed into the monitor.
    */ 
  bit use_external_port_monitor = 0;
  /** @endcond */

  /** 
    * @groupname axi_tlm_generic_payload
    * In active mode, creates a tlm_generic_payload_sequencer sequencer capable
    * of generating UVM TLM Generic Payload transactions and connects the
    * master sequencer to it.  The master sequencer starts a layering sequence that gets
    * transactions from the tlm_generic_payload_sequencer, converts them to (one or more) AXI
    * transaction(s) and sends them to the driver.
    * Snoop requests are still fulfilled by the svt_axi_master_snoop_sequencer.
    * 
    * AXI transactions observed by the agent
    * are also made available as TLM GP transactions through the
    * tlm_generic_payload_observed_port in the monitor. Note that the TLM GP
    * transactions issued through the analysis port may not match one to one with GP
    * sequence items created by the tlm_generic_payload_sequencer because the
    * GP sequence items may have to be mapped
    * to multiple AXI transactions according to protocol requirements. The
    * TLM GP that is available through the tlm_generic_payload_observed_port of
    * the monitor is a direct mapping of the observed AXI transactions converted to a TLM GP.
    * No attempt is made to re-assemble a set of AXI transaction into a larger TLM GP.
    * 
    * The layering sequence that converts the TLM GP to AXI transactions is the
    * svt_axi_tlm_gp_to_axi_sequence and is available at
    * $DESIGNWAREHOME/vip/svt/amba_svt/<ver>/axi_master_agent_svt/sverilog/src/vcs/svt_axi_tlm_gp_sequence_collection.svp 
    * Transactions created by the layering sequence are of type
    * cust_svt_tlm_gp_to_axi_master_transaction. Any user constraints specific
    * to AXI must be provided in a class extended from this class.
    * 
    * In passive mode, observed AXI transactions are made available as TLM GP
    * transactions through the tlm_generic_payload_observed_port in the
    * monitor.
    */
  bit use_tlm_generic_payload = 0;

  /** 
    * @groupname axi_tlm_generic_payload
    * In active mode, creates an AMBA-PV-compatible socket that can be used to
    * connect AXI Master VIP component to an AMBA-PV master model. 
    * 
    * Enabling this functionality causes the instantiation of socket b_fwd of
    * type uvm_tlm_b_target_socket, and socket b_snoop of type
    * uvm_tlm_b_initiator_socket, in class svt_axi_master_agent.

    * Generic payload transactions received through the forward b_fwd interface
    * are executed on the tlm_generic_payload_sequencer in the agent.

    * When this option is set, the svt_axi_ace_snoop_request_to_tlm_gp_sequence
    * reactive sequence is started on the AXI VIP master snoop sequencer. Snoop
    * transaction requests received by the AXI VIP master snoop sequencer are translated to
    * equivalent tlm_generic_payload transactions with the
    * #svt_amba_pv_extension attached. The extended Generic Payload transactions
    * are then sent to the AMBA-PV master model via the backward b_snoop interface.
    * The receive response from AMBA-PV master model is then interpreted to
    * complete the snoop transaction request and executed on the AXI VIP master snoop
    * sequencer.
    * 
    * Should the AXI VIP master fulfill the snoop requests natively (i.e. the
    * default behavior when this option is not set), the snoop response sequence
    * should be restored to the default using:
    * 
    * <code>
    * uvm_config_db#(uvm_object_wrapper)::set(this, "master[0].snoop_sequencer.run_phase", "default_sequence",
    *                                         /#svt_axi_ace_master_snoop_response_sequence::type_id::/#get());
    * </code>
    * 
    * When this option is set, it implies that #use_tlm_generic_payload is also set, whether
    * it actually is or not.
    */
  bit use_pv_socket = 0;

 /** Enables the UVM REG feature of the AXI agent.  
   * Applicable only when svt_axi_port_configuration::axi_interface_type is AXI3.
   * <b>type:</b> Static 
   */
  bit uvm_reg_enable = 0;

 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables checking of wdata/tdata only on valid byte lanes based on wstrb/tstrb. 
    * In a disabled state, whole wdata/tdata as seen on the bus will be considered.
    * <b>type:</b> Dynamic 
    */
  bit check_valid_data_bytes_only_enable = 1;

  /**
    * @groupname axi3_4_timeout_config
    * A timer which is started when a transaction starts. If the transaction
    * does not complete by the set time, an error is repoted. The timer is
    * incremented by 1 every clock and is reset when the transaction ends. 
    * If set to 0, the timer is not started
    */
  int xact_inactivity_timeout = 0;

 /**
   * @groupname ace_config 
   * If this attribute is enabled it will allow snoop response data_transfer bit for
   * MAKEINVALID  transaction to be set as 1. This behaviour is permitted by protocol
   * but it is not expected snoop response for MAKEINVALID 
 */
  bit  data_transfer_for_makeinvalid_snoop_enable =0;

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /** 
   * log_base_2 of \`SVT_AXI_MAX_DATA_WIDTH. 
   * Used only as a helper attribute to randomize data_width.
   *
   * This parameter is not required to be set by the user.
   */
  int log_base_2_max_data_width;
 
  /** 
   * log_base_2 of \`SVT_AXI_ACE_SNOOP_DATA_WIDTH. 
   * Used only as a helper attribute to randomize snoop_data_width.
   *
   * This parameter is not required to be set by the user.
   */
  int log_base_2_max_snoop_data_width; 

  /** 
   * log_base_2 of \`SVT_AXI_MAX_CACHE_LINE_SIZE. 
   * Used only as a helper attribute to randomize cache_line_size.
   *
   * This parameter is not required to be set by the user.
   */
  int log_base_2_max_cache_line_size;

  /**
    * Indicates if the address range of the slave component
    * has been set
    */
  bit is_slave_addr_range_set = 0;

  /**
    * Stores the log_base_2 of the desired data_width.
    * Used only as a helper attribute to randomize data_width.
    * This parameter is first randomized and the data_width
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_data_width;

  /**
    * Stores the log_base_2 of the desired snoop_data_width.
    * Used only as a helper attribute to randomize snoop_data_width.
    * This parameter is first randomized and the snoop_data_width
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_snoop_data_width;

  /**
    * Stores the log_base_2 of the desired cache_line_size.
    * Used only as a helper attribute to randomize cache_line_size.
    * This parameter is first randomized and the cache_line_size
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_cache_line_size;

  /**
    * Stores the log_base_2 of the desired atomicity_size.
    * Used only as a helper attribute to randomize atomicity_size.
    * This parameter is first randomized and the atomicity_size
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_atomicity_size;

  /** @endcond */

  /** 
    * @groupname axi3_signal_width
    * Address width of this port in bits.
    * When svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE,
    * this parameter also sets the width of signal caddr.
    *
    * NOTE: currently same address width is considered for both coherent read or write address
    *       channels and snoop address channels. So, there is no separate snoop address width
    *       parameter supported at the moment.
    * Configuration type: Static
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE 
  rand int addr_width = `SVT_AXI_MAX_ADDR_WIDTH;
`else    
  rand int addr_width = `SVT_AXI_MAX_ADDR_WIDTH - `SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH;
`endif   

  /** 
    * @groupname axi4_signal_width
    * Address user width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int addr_user_width = `SVT_AXI_MAX_ADDR_USER_WIDTH;

  /** 
    * @groupname axi3_signal_width
    * Data width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int data_width = `SVT_AXI_MAX_DATA_WIDTH;

  /** 
    * @groupname axi4_signal_width
    * Data user width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int data_user_width = `SVT_AXI_MAX_DATA_USER_WIDTH;
 
  /** 
    * @groupname axi4_signal_width
    * Response user width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int resp_user_width = `SVT_AXI_MAX_BRESP_USER_WIDTH;

  /** 
    * @groupname ace_config
    * Cache line size in bytes for this master.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int cache_line_size = `SVT_AXI_MAX_CACHE_LINE_SIZE;

  /** 
    * @groupname ace_config
    * Aligned size in bytes for the snoop corresponding to starting address.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates the size to which the snoop corresponding to the starting address
    * of a multi-cacheline access is aligned. For example, if the cacheline size
    * is 64 bytes and the coherent address of a READONCE transaction is 0x70,
    * the corresponding snoop address may be 0x40 or 0x70. If the snoop address
    * sent is 0x40, this value must be set to the same as the cacheline size which is
    * 64 bytes. If the snoop address sent is 0x70, this value can be set to 16 bytes.
    * This will help in more accurate correlation of coherent and snoop transactions.
    * The default is 0. If unchanged, the system monitor will use the cacheline size
    * for this value, assuming that all snoops are aligned to cacheline size. 
    * Configuration type: Static
    */
  rand int start_addr_snoop_aligned_size = 0;

  /** 
    * @groupname ace_config
    * Number of cache lines in the master.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int num_cache_lines = `SVT_AXI_MAX_NUM_CACHE_LINES;

  /** 
    * @groupname ace_config
    * Enables AWAKEUP sideband signal in the VIP when this bit is set to '1'.
    * by default AWAKEUP signal will be '0' when this bit is enabled.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand bit awakeup_enable = 0;

  /** 
    * @groupname ace_config
    * Enabling this feature will allow transactions to wait to send address phase
    * until the previous transaction's datahandshake is done. This will result
    * in unexpected delays. Hence this parameters is disabled by default.
    * 
    * This parameter is applicable when 
    * svt_axi_port_configuration::axi_interface_type is set to AXI3 or AXI4.
    *
    * Configuration type: Static
    */
  rand bit prev_xact_data_handshake_ref_event_enable = 0;

  /** 
    * @groupname ace_config
    * Toggles AWAKEUP sideband signal in the VIP during idle period of read or
    * write channel.
    * Asserts and then de-assert AWAKEUP with the range of programed number of 
    * 'awakeup_toggle_min_delay_during_idle' to 'awakeup_toggle_max_delay_during_idle'.
    * If there is no transaction observed in read or write channel, then AWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int awakeup_toggle_min_delay_during_idle = 1;

  /** 
    * @groupname ace_config
    * Toggles AWAKEUP sideband signal in the VIP during idle period of read or
    * write channel.
    * Asserts and then de-assert AWAKEUP with the range of programed number of 
    * 'awakeup_toggle_min_delay_during_idle' to 'awakeup_toggle_max_delay_during_idle'.
    * If there is no transaction observed in read or write channel, then AWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int awakeup_toggle_max_delay_during_idle = 5;


  /** 
    * @groupname ace_config
    * Enables ACWAKEUP sideband signal in the VIP when this bit is set to '1'.
    * by default ACWAKEUP signal will be '0' when this bit is enabled.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand bit acwakeup_enable = 0;

  /** 
    * @groupname ace_config
    * Toggles ACWAKEUP sideband signal in the VIP during idle period of snoop channel.
    * Asserts and then de-assert ACWAKEUP with the range of programed number of 
    * 'acwakeup_toggle_min_delay_during_idle' to 'acwakeup_toggle_max_delay_during_idle'.
    * If there is no snoop transaction observed in snoop channel, then ACWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int acwakeup_toggle_min_delay_during_idle = 1;

  /** 
    * @groupname ace_config
    * Toggles ACWAKEUP sideband signal in the VIP during idle period of snoop channel.
    * Asserts and then de-assert ACWAKEUP with the range of programed number of 
    * 'acwakeup_toggle_min_delay_during_idle' to 'acwakeup_toggle_max_delay_during_idle'.
    * If there is no snoop transaction observed in snoop channel, then ACWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int acwakeup_toggle_max_delay_during_idle = 5;
  
  /** 
    * @groupname ace_signal_width
    * Snoop Data width of the cddata port in bits.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    *
    * Configuration type: Static
    */
  rand int snoop_data_width = `SVT_AXI_ACE_SNOOP_DATA_WIDTH;

  /**
    * @groupname axi3_4_config
    * Acronym for "What You See is What You Get". Applicable to the
    * svt_axi_transaction::data and svt_axi_transaction::wstrb fields of a
    * transaction. If this bit is set to 1, whatever is configured in the
    * svt_axi_transaction::data and  svt_axi_transaction::wstrb fields is
    * transmitted "as is" by the master. Also, in the transaction object
    * generated by monitor, the monitor populates the svt_axi_transaction::data
    * and  svt_axi_transaction::wstrb fields "as is", as seen on the bus. If
    * this bit is set to 0 (default), the data must be stored right-justified by
    * the user. The model will drive the data on the correct lanes.
    *
    * Refer to the documentation of svt_axi_transaction::data and 
    * svt_axi_transaction::wstrb for more details
    */
  rand bit wysiwyg_enable = 0;

  /**
    * @groupname axi3_4_config
    * Applicable when #wysiwyg_enable is set.
    * Indicates if the VIP should consider validity of wstrb in transactions
    * when #wysiwyg_enable is set. When wysiwyg_enable is set, the driver
    * checks that #wstrb is set only for valid byte lanes of each beat.  In
    * certain applications, wstrb may have to be asserted for other byte lanes
    * as well. In such applications, this bit should be set. This results in
    * the following: 
    * <br>
    * Constraints in transaction are relaxed for wstrb. wstrb
    * values will be random and may be asserted for invalid byte lanes. 
    * <br>
    * driver does not check for validity of wstrb in transaction based on valid
    * byte lanes.
    * <br>
    * Note that this will result in a non-AXI compliant behaviour, in that
    * wstrb may be asserted for invalid byte lanes based on what the user
    * programs. If this bit is set for the slave, and if the user wants memory
    * to be updated based on the transactions, the memory sequence shipped with
    * the VIP should not be used. For VMM based testbenches, the generator_type
    * should not be set to MEMORY_RESPONSE_GEN. This is because the APIs that
    * access memory are based on valid assertion of byte strobes.  The user
    * must use user-defined APIs and sequences to access memory if this bit is
    * set in the slave.
    */ 
  bit ignore_wstrb_check_for_wysiwyg_format = 0;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the WSTRB signal on byte count calculation in the VIP 
    * By default this configuration parameter is set to 0 to calculate the byte count using burst_size and burst_length,
    * if this parameter is set 1 then wstrb is used to calculate the byte count
    * <b>type:</b> Static
    */
  rand bit get_byte_count_from_wstrb_enable      = 0;

   /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWREGION signal in the VIP 
    * <b>type:</b> Static
    */

  rand bit awregion_enable   = 0;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARREGION signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arregion_enable   = 0;
 
  /** @cond PRIVATE */
  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awid_enable       = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWLEN signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awlen_enable   = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWSIZE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awsize_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWBURST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awburst_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWLOCK signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awlock_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWCACHE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awcache_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWPROT signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awprot_enable     = 1;
  /** @endcond */

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWQOS signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awqos_enable      = 0;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the WLAST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit wlast_enable      = 1;

  /** @cond PRIVATE */
  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the WSTRB signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit wstrb_enable      = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the BID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit bid_enable        = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the BRESP signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit bresp_enable      = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arid_enable       = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARLEN signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arlen_enable   = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARSIZE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arsize_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARBURST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arburst_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARLOCK signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arlock_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARCACHE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arcache_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARPROT signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arprot_enable     = 1;
  /** @endcond */

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARQOS signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arqos_enable      = 0;

  /** @cond PRIVATE */
  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the RID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit rid_enable        = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the RRESP signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit rresp_enable      = 1;
  /** @endcond */

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the RLAST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit rlast_enable      = 1;

  /** 
    * @groupname axi3_4_config
    * Enables AWUSER sideband signal in the VIP. AWUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit awuser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables WUSER sideband signal in the VIP. WUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit wuser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables BUSER sideband signal in the VIP. BUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit buser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables ARUSER sideband signal in the VIP. ARUSER signal can be used when
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit aruser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables RUSER sideband signal in the VIP. RUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit ruser_enable      = 0;

  `ifdef SVT_AXI_QVN_ENABLE
  /** 
    * @groupname axi_qvn_config
    * Enables QVN support in the VIP. QVN signals can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * All QVN configuration parameters comes into effect only when qvn_enable bit is set.
    * Any parameter which is declared as a bit-vector to support all Virtual Network in the
    * system, is sized by `define macro "SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK".
    *
    * If a system should support a maximum number of 5 Virtual Networks then user should
    * define SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK as 5
    * <b>type:</b> Static
    */
  rand bit qvn_enable      = 0;

  /** 
    * @groupname axi_qvn_config
    * Specifies how many Virtual Network a particular master supports for Read Address channel
    * <b>type:</b> Static
    */
  rand int qvn_num_virtual_network_supported_ar_chnl = 1;

  /** 
    * @groupname axi_qvn_config
    * Specifies how many Virtual Network a particular master supports for Write Address channel.
    * Write Data channel must support Virtual Networks same as Write Address channel so there is
    * no need of having seperate configuration for Write Data channel.
    * <b>type:</b> Static
    */
  rand int qvn_num_virtual_network_supported_aw_chnl = 1;

  /** 
    * @groupname axi_qvn_config
    * Lists Virtual Networks which are supported by a master/slave port for Read-Address Channel.
    * It provides an array of bits each representing a Virtual Network in the system. Index of 
    * each bit denotes ID of the Virtual Network, represented by that bit.
    * If any bit of this array is set to '1' then that means Virtual Network with ID equal to
    * index of that bit, is supported by this port. If a bit in this array is set to '0' then
    * that means Virtual Network with ID equal to its index is not supported by this port.
    * Initial Value:  all bits are set to '0' i.e. no Virtual Network is supported by default.
    * Example:  If a port must be configured to use Virtual Network 1 and 3 to be used for its
    *           Read-Address channel then user should configure as follows:
    *   (manual configuration without randomization)  - reset all bits to '0'
    *   foreach(qvn_supported_virtual_network_queue_ar_chnl[index]) qvn_supported_virtual_network_queue_ar_chnl[index] = 0; 
    *   set '1' for Virtual Network 1 =>  qvn_supported_virtual_network_queue_ar_chnl[1] = 1;
    *   set '1' for Virtual Network 3 =>  qvn_supported_virtual_network_queue_ar_chnl[3] = 1;
    */
  rand bit qvn_supported_virtual_network_queue_ar_chnl[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] ;

  /** 
    * @groupname axi_qvn_config
    * Lists Virtual Networks which are supported by a master/slave port for Write Address Channel.
    * This array of bits also indicate which Virtual Networks are supported by this port similar
    * to the array qvn_supported_virtual_network_queue_ar_chnl described above.
    * Initial Value:  all bits are set to '0' i.e. no Virtual Network is supported by default.
    * Example:  If a port must be configured to use Virtual Network 0 and 2 to be used for its
    *           Write-Address channel then user should configure as follows:
    *   (manual configuration without randomization)  - reset all bits to '0'
    *   foreach(qvn_supported_virtual_network_queue_aw_chnl[index]) qvn_supported_virtual_network_queue_aw_chnl[index] = 0; 
    *   set '0' for Virtual Network 1 =>  qvn_supported_virtual_network_queue_aw_chnl[1] = 1;
    *   set '1' for Virtual Network 2 =>  qvn_supported_virtual_network_queue_aw_chnl[2] = 1;
    */
  rand bit qvn_supported_virtual_network_queue_aw_chnl[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] ;

  /**
    * @groupname axi_qvn_config
    * Specifies maximum number of clock cycles (interface clock) within which a Master must use
    * all the tokens it has been granted on read address channel.
    * Port Monitor uses this parameter to assert warning if Master didn't use its granted token 
    * within this bounded time period.
    */

   /* If a Master is not able to use a token, then after this timelimit that token will be reclaimed
    * by the slave which, granted it and Master will remove this token from its reserved token pool.
    *
    * - So, it is important to set suitable value for this parameter. If it is set too low, then
    * most tokens may expire before it could be used and hance leading to increased token request.
    *
    * - If it is set below minimum no. of cycles a master needs to use a token then all tokens will
    * expire and none could be used to issue a transaction to AXI channels.
    *
    * - On the other hand if it uses too high value, then due to under usage of token or over-request
    * of tokens by a Master, there is a possibility of accumulating large number of tokens in the
    * token-pool of that master and hence causing possible blockage to other masters.
    *
    * - If it is set to Zero then that indicates there is no timelimit for token usage i.e. once a 
    * token is acquired it will remain in the token-pool of that master until used for sending a
    * transaction.
    * .
    */
  rand int qvn_read_addr_token_usage_timelimit[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies maximum number of clock cycles (interface clock) within which a Master must use
    * all the tokens it has been granted on write address channel.
    * Port Monitor uses this parameter to assert warning if Master didn't use its granted token 
    * within this bounded time period.
    */
  rand int qvn_write_addr_token_usage_timelimit[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies maximum number of clock cycles (interface clock) within which a Master must use
    * all the tokens it has been granted on write data channel.
    * Port Monitor uses this parameter to assert warning if Master didn't use its granted token 
    * within this bounded time period.
    */
  rand int qvn_write_data_token_usage_timelimit[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Pre-Allocated Token for Read Address Channel
    * An integer array is provided to hold pre_allocated token number for AR channel of
    * each corresponding Virtual Network. Index of an array element indicates for which
    * virtual network it holds pre_allocated token number.
    * Initial Value : all elements of this array is initiallized to \`SVT_AXI_QVN_MIN_NUM_AR_PRE_ALLOCATED_TOKEN
    * Example: if AR channel of Virtual Network 2 should be set to 1 then configure as
    *   qvn_num_ar_pre_allocated_token_vn[2] = 1;
    */
  rand int qvn_num_ar_pre_allocated_token_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Pre-Allocated Token for Write Address Channel
    * An integer array is provided to hold pre_allocated token number for AR channel of
    * each corresponding Virtual Network. Index of an array element indicates for which
    * virtual network it holds pre_allocated token number.
    * Initial Value : all elements of this array is initiallized to \`SVT_AXI_QVN_MIN_NUM_AW_PRE_ALLOCATED_TOKEN
    * Example: if AW channel of Virtual Network 2 should be set to 1 then configure as
    *   qvn_num_aw_pre_allocated_token_vn[2] = 1;
    */
  rand int qvn_num_aw_pre_allocated_token_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Indicates if same AXI ID can be used between two different Virtual Network or not.
    * - If set to "0" then at any given point of time no two different Virtual Networks will
    * use same ID for transactions sent to AXI channels associated with those VNs.
    * - if set to "1" then same AXI ID can be used by two different VN without any restriction.
    * .
    *
    * NOTE: if same ID is used for AXI transactions issued to two different VN may get
    * blocked by interconnect in order to observe AXI ID ordering rule. Because of this, a
    * transaction received first will block another transaction with same ID received later,
    * even if transaction that was received first, can't make any progress.
    */
  rand int qvn_allow_id_used_in_other_vn = 0;

  /**
    * @groupname axi_qvn_config
    * Specifies number of granted token a master can keep unused for each virtual network
    * it supports on read address channel. It helps in defining how system resources will be used
    * otherwise, a master can issue large number of token requests and once granted those tokens 
    * may remain unused reserving system resources and in turn blocking other masters, if it shares 
    * same Virtual Network or if slave uses shared token for different masters.
    * 
    * NOTE: by default it is randomized within range [\`SVT_AXI_QVN_NUM_MIN_ALLOWED_UNUSED_TOKEN:\`SVT_AXI_QVN_NUM_MAX_ALLOWED_UNUSED_TOKEN]
    * 
    */
  rand int qvn_max_num_read_addr_unused_token[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of granted token a master can keep unused for each virtual network
    * it supports on write address channel. 
    * NOTE: by default it is randomized within range [\`SVT_AXI_QVN_NUM_MIN_ALLOWED_UNUSED_TOKEN:\`SVT_AXI_QVN_NUM_MAX_ALLOWED_UNUSED_TOKEN]
    * 
    */
  rand int qvn_max_num_write_addr_unused_token[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of granted token a master can keep unused for each virtual network
    * it supports on write data channel. 
    * NOTE: by default it is randomized within range [\`SVT_AXI_QVN_NUM_MIN_ALLOWED_UNUSED_TOKEN:\`SVT_AXI_QVN_NUM_MAX_ALLOWED_UNUSED_TOKEN]
    * 
    */
  rand int qvn_max_num_write_data_unused_token[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of clock cycles (interface clock) within which slave must assert ready
    * to the master requesting token for read address channel. If slave doesn't assert ready i.e.
    * grant token to the master within this specified clock cycles then timeout will occur and
    * error will be asserted. Master driver waiting for the ready will also come out and abort
    * the transaction.
    *
    * NOTE: if this timeout value is set to '0' then timeout will be disabled and master will
    * wait forever until token request ready is asserted by slave for read address channel.
    */
  rand int unsigned qvn_ar_token_request_ready_timeout_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of clock cycles (interface clock) within which slave must assert ready
    * to the master requesting token for write address channel. If slave doesn't assert ready i.e.
    * grant token to the master within this specified clock cycles then timeout will occur and
    * error will be asserted. Master driver waiting for the ready will also come out and abort
    * the transaction.
    *
    * NOTE: if this timeout value is set to '0' then timeout will be disabled and master will
    * wait forever until token request ready is asserted by slave for write address channel.
    */
  rand int unsigned qvn_aw_token_request_ready_timeout_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of clock cycles (interface clock) within which slave must assert ready
    * to the master requesting token for write data channel. If slave doesn't assert ready i.e.
    * grant token to the master within this specified clock cycles then timeout will occur and
    * error will be asserted. Master driver waiting for the ready will also come out and abort
    * the transaction.
    *
    * NOTE: if this timeout value is set to '0' then timeout will be disabled and master will
    * wait forever until token request ready is asserted by slave for write data channel.
    */
  rand int unsigned qvn_w_token_request_ready_timeout_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];


  /**
    * @groupname axi_qvn_config
    * Specifies number of Token Slave can have for AR channel for a particular Virtual Network
    * This means Slave has these many token resources to allocate to Master and can't give token
    * more than the value specified here.
    * Note: Since Master is pre-allocated with certain number of token Slave will begin with 
    *       number of Tokens as specified here minus master pre_allocated_token for AR channel
    */
  rand int qvn_slave_ar_token_size_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Token Slave can have for AW channel for a particular Virtual Network
    * This means Slave has these many token resources to allocate to Master and can't give token
    * more than the value specified here.
    * Note: Since Master is pre-allocated with certain number of token Slave will begin with 
    *       number of Tokens as specified here minus master pre_allocated_token for AW channel
    */
  rand int qvn_slave_aw_token_size_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Token Slave can have for W channel for a particular Virtual Network
    * This means Slave has this many token resource to allocate to Master and can't give token
    * more than the value specified here.
    * Note: Master doesn't have any pre-allocated token for Write Data channel so, Slave will 
    *       begin with same number of Tokens as specified by this parameter.
    */
  rand int qvn_slave_w_token_size_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies max number of outstanding token request slave can grant for read address channal for a VN, 
    * in accordance with slaves acceptance capability.
    * Note: This is exclusive of pre allocated token for the VN  
    */
   rand int unsigned qvn_slave_max_outstading_token_for_rd_addr_chan_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies max number of outstanding token request slave can grant for write address channal for a VN, 
    * in accordance with slaves acceptance capability.
    * Note: This is exclusive of pre allocated token for the VN  
    */
   rand int unsigned qvn_slave_max_outstading_token_for_wr_addr_chan_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies max number of outstanding token request slave can grant for write data channal for a VN, 
    * in accordance with slaves acceptance capability.
    */
   rand int unsigned qvn_slave_max_outstading_token_for_wr_data_chan_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

   /**
    * @groupname axi_qvn_config
    * Mode to control the assertion of V*READYVNx signal. This allows QVN enabled Slaves to assert
    * token request grant ready signal for any Virtual Network of each channel AR, AW, W
    *
    * 0 - Assert V*READY in responce to assertion of V*VALID for token request 
    * 1 - Assert V*READY before assertion of V*VALID for token request, subjected to token availability
    */  
   rand bit qvn_slave_aw_ready_assertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_w_ready_assertion_mode  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_ar_ready_assertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
  
   /*
    * @groupname axi_qvn_config
    * Mode to control the de-assertion of V*READYVNx signal. This flage is only 
    * applicable if v*ready_assertion_mode is set to ONE.
    * 0 - Keep V*READY till assertion of V*VALID.  
    * 1 - Deassert V*READY after some time if V*VALID is not asserted. 
    */  
   rand bit qvn_slave_aw_ready_deassertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_w_ready_deassertion_mode  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_ar_ready_deassertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};


  `endif

  /** 
    * @groupname axi3_4_config
    * Enables optimistic flow control for Write Data channel in the VIP.  
    * The flow control of the write data channel is determined by the settings 
    * in num_outstanding_xact and num_outstanding_write_xact. Based on these 
    * settings wready is deasserted when the number of outstanding transactions
    * reach the threshold set by these parameters. This parameter controls the 
    * deassertion of wready when the threshold is reached. Since AXI allows data 
    * before address, a new transaction can start with data. When this parameter 
    * is disabled, both awready and wready are deasserted when threshold of maximum
    * outstanding transactions are reached. Note however that this will prevent data
    * of any already outstanding transactions from being continuously accepted
    * (that is with wready continuously high) and therefore can reduce throughput
    * If this parameter is set, only awready is deasserted when the threshold is reached.
    * This allows data of outstanding write transactions to be continously accepted
    * with wready maintained high continuosly. wready is deasserted only on observing
    * a new transaction which will cross the threshold. Thus, setting this configuration
    * assumes that write data before address doesn't come once the threshold for maximum
    * outstanding transactions is reached and thus keeps wready asserted. 
    * Whereas disabling this configuration assumes that write data before address might 
    * come and thus deasserts wready when number of outstanding transactions
    * reach the threshold.
    * <b>type:</b> Dynamic
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand bit wdata_optimistic_flow_control_enable = 0;
`else
  rand bit wdata_optimistic_flow_control_enable = 1;
`endif

   /** 
    * @groupname axi3_4_config
    * Passive slave memory needs to be aware of the backdoor writes to memory.
    * Setting this configuration allows passive slave memory to be updated according to
    * RDATA seen in the transaction coming from the slave. Note that the passive slave 
    * memory is updated when all read data beats have been transmitted and accepted.
    * For an EXCLUSIVE transaction memory is updated only if all beats have an EXOKAY response.
    * For a normal transaction, memory is updated only if all beats have an OKAY response.
    * <b>type:</b> Static
    */
  rand bit memory_update_for_read_xact_enable = 0;

  /**
    * @groupname axi3_signal_width
    * Indicates if separate widths are required for ID  of write channel 
    * (AWID,WID and BID) and for ID of read channel(ARID and RID).
    * If set to 1, read_chan_id_width and write_chan_id_width are used
    * for setting the widths of the ID signals of corresponding channels.
    * If set to 0, id_width is used for setting the widths of all
    * ID signals.
    * This value must be consistent across all the ports in the system.
    *
    * Configuration type: Static
    */
  rand bit use_separate_rd_wr_chan_id_width = 0;

  /**
    * @groupname axi3_signal_width
    * If port is of kind MASTER:
    * This parameter defines the ID width of the master.
    * <br>
    * If port is of kind SLAVE:
    * This parameter defines the ID width of the slave. If an
    * interconnect is present, the ID width of the slave should
    * consider the maximum ID width of the masters in the system
    * and also consider additional bits required to represent
    * each master in the system.
    * <br>
    * Valid only when use_separate_rd_wr_chan_id_width is set to 0.
    *
    * Configuration type: Static
    */
  rand int id_width  = `SVT_AXI_MAX_ID_WIDTH;

  /**
    * @groupname axi3_signal_width
    * Represents the width of ARID and RID.  
    * Valid only when use_separate_rd_wr_chan_id_width is set to 1.
    * For slaves, the same considerations given for id_width are applicable.
    *
    * Configuration type: Static
    */
  rand int read_chan_id_width = `SVT_AXI_MAX_ID_WIDTH;

  /**
    * @groupname axi3_signal_width
    * Represents the width of AWID, WID and BID.  
    * Valid only when use_separate_rd_wr_chan_id_width is set to 1.
    * For slaves, the same considerations given for id_width are applicable.
    *
    * Configuration type: Static
    */
  rand int write_chan_id_width = `SVT_AXI_MAX_ID_WIDTH;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines whether Normal transactions IDs can overlap with barrier transactions IDs.
    *
    * Configuration type: Static
    */
  rand bit barrier_id_overlap  = 1;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the min ID value of the master for barrier transactions.
    *
    * Configuration type: Static
    */
  rand int barrier_id_min  = 0;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the min ID value of the master for barrier transactions.
    *
    * Configuration type: Static
    */
  rand int barrier_id_max  = ((1<<(`SVT_AXI_MAX_ID_WIDTH))-1);

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines whether Normal transactions IDs can overlap with DVM transactions IDs.
    *
    * Configuration type: Static
    */
  rand bit dvm_id_overlap  = 1;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the min ID value of the master for dvm transactions.
    *
    * Configuration type: Static
    */
  rand int dvm_id_min  = ((1<<(`SVT_AXI_MAX_ID_WIDTH/2))-1);

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the max ID value of the master for dvm transactions.
    *
    * Configuration type: Static
    */
  rand int dvm_id_max  = ((1<<(`SVT_AXI_MAX_ID_WIDTH))-1);

  /**
   * Indicates how the information regarding the source master is 
   * transmitted to the slave
   * If set to STATIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES, the source master information
   * is static and is defined by #source_master_id_xmit_to_slaves
   * If set to DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES, the source master information
   * is based on the value defined in svt_axi_transaction::dynamic_source_master_id_xmit_to_slaves
   * The value in dynamic_source_master_id_xmit_to_slaves must be populated by the user
   * in a system monitor callback issued at the start of the transaction.
   * If set to CUSTOM_SOURCE_MASTER_ID_XMIT_TO_SLAVES, the user must define 
   * svt_axi_system_configuration::is_master_id_and_slave_id_correlated to indicate
   * whether ID requirements for master and slave transactions are met 
   */
  source_master_id_xmit_to_slaves_type_enum source_master_id_xmit_to_slaves_type = STATIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES;
  
 /**
   * @groupname ace5_config 
   * Indicates whether data check parity feature is enable or not.
   * If set to ODD_PARITY_BYTE_DATA, then only on data check signals odd parity algorthim is used,
   * every 8bit of data is calculated and generated singles bit of datachk parity bit.
   * If set to ODD_PARITY_BYTE_ALL, then on both data check signals and control check signals odd parity algorthim is used.  
   * By default this enum is set to FALSE, which means data check fetaure is disabled.
   */ 
  check_type_enum check_type = FALSE;



  /**
    * @groupname axi_generic_config 
    * Applicable only when
    * svt_axi_system_configuration::id_based_xact_correlation_enable is set
    * If port is of kind MASTER:
    * This parameter defines the value that the interconnect assigns when
    * routing transactions to slave for all transactions originating from this
    * master. This value is specified in some bits of AxID of the transaction
    * that is routed to slave. This value must be based on the max value that
    * can be supported based on
    * svt_axi_system_configuration::source_master_info_id_width. For example, if the
    * interconnect uses 3 bits of AxID of the outgoing slave transaction to
    * specify the source master of the transaction,
    * svt_axi_system_configuration::source_master_info_id_width must be set to 3 and
    * this value must be less than 7. For more details, please refer
    * svt_axi_system_configuration::id_based_xact_correlation_enable
    */
  bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id_xmit_to_slaves;

  /**
    * @groupname axi_generic_config
    * Applicable only when
    * svt_axi_system_configuration::id_based_xact_correlation_enable is set
    * and axi_port_kind is MASTER
    * Indicates that the ID from this master is passed through without any
    * change when the interconnect routes it to the slaves. If this is set,
    * all transactions from this master are not appended with source master
    * information when routing to slaves
   */ 
  rand bit is_source_master_id_and_dest_slave_id_same = 0;

  /**
    * @groupname axi_generic_config 
    * Applicable only when svt_axi_system_configuration::id_based_xact_correlation_enable is set
    * If this parameter is set to zero, system monitor will not do id based correlation
    * for any transactions initiated/received at this specific port, this provides the option
    * for the user to avoid or select id based correlation for specific ports 
    * default value is 1.
    */
  bit id_based_xact_correlation_enable =1'b1;

  /** 
    * @groupname axi_generic_config
    * The byte boundary at which a master transaction is split to be
    * transmitted to two different slaves. This must be defined in cases where
    * pre_add_to_input_xact_queue callback in svt_axi_system_monitor_callback
    * is used to indicate that a master transaction is split and transmitted to
    * two different slaves. This parameter defines the boundary at which a
    * transaction is split
    *
    * Configuration type: Static
    */
  rand int byte_boundary_for_master_xact_split = `SVT_AXI_MAX_BYTE_BOUNDARY_FOR_MASTER_XACT_SPLIT;

  /**
   * @groupname ace_config
   * Enables support for WriteEvict transaction
   * Configuration type: Static
   */
  rand bit writeevict_enable = 0;

  /**
   * @groupname ace_config
   * Enables AWUNIQUE signal 
   * Configuration type: Static
   */
  rand bit awunique_enable = 0;

  /** 
    * @groupname axi3_4_config
    * Specifies the number of outstanding transactions a master/slave
    * can support.
    * num_outstanding_xact = -1 is not supported for AXI4_STREAM
    * <br>
    * MASTER:
    * If the number of outstanding transactions is equal to this
    * number, the master will refrain from initiating any new 
    * transactions until the number of outstanding transactions
    * is less than this parameter.
    * <br>
    * SLAVE:
    * If the number of outstanding transactions is equal to 
    * this number, the slave will not assert ARREADY/AWREADY
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * <br>
    * If #num_outstanding_xact = -1 then #num_outstanding_xact will not 
    * be considered , instead #num_read_outstanding_xact and 
    * #num_write_outstanding_xact have an effect.
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
  rand int num_outstanding_xact = 4;

  /**
    * @groupname axi3_4_config
    * Specifies the number of READ outstanding transactions a master/slave
    * can support.
    * <br>
    * MASTER:
    * If the number of outstanding transactions is equal to this
    * number, the master will refrain from initiating any new 
    * transactions until the number of outstanding transactions
    * is less than this parameter.
    * <br>
    * SLAVE:
    * If the number of outstanding transactions is equal to 
    * this number, the slave will not assert ARREADY
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * <br>
    * This parameter will have an effect only if #num_outstanding_xact = -1.
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
  rand int num_read_outstanding_xact = 4;

  /** 
    * @groupname axi3_4_config
    * Specifies the number of WRITE outstanding transactions a master/slave
    * can support.
    * <br>
    * MASTER:
    * If the number of outstanding transactions is equal to this
    * number, the master will refrain from initiating any new 
    * transactions until the number of outstanding transactions
    * is less than this parameter.
    * <br>
    * SLAVE:
    * If the number of outstanding transactions is equal to 
    * this number, the slave will not assert AWREADY
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * <br>
    * This parameter will have an effect only if #num_outstanding_xact = -1.
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
  rand int num_write_outstanding_xact = 4;

  /** 
    * @groupname ace_config
    * Specifies the number of outstanding snoop transactions a master
    * can support. Applicable when axi_interface_type == AXI_ACE.
    * If the number of outstanding snoop transactions is equal to 
    * this number, the master will not assert ACREADY 
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_SNOOP_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand int num_outstanding_snoop_xact = 4;
`else
  rand int num_outstanding_snoop_xact = 16;
`endif  

  /** 
    * @groupname axi_generic_config
    * 
    * Enables a separate port/export in the slave driver
    * (delayed_response_request_export) and sequencer
    * (delayed_response_request_port) through which the user can input response
    * data in a delayed manner.  When disabled all data and response
    * information related to a transaction must be given back to the driver
    * from the sequencer in the same timestamp as it receives a transaction
    * from the monitor.  When enabled, the user has flexibility to provide
    * response and data information at a later point in time through the
    * response port in the slave driver, although parameters related to the
    * delays to be applied for driving ARREADY, AWREADY and WREADY signals need
    * to be provided in the same timestamp. 
    * Refer to the user guide for a detailed description of the usage of this
    * parameter.
    */ 
  bit enable_delayed_response_port = 0;

  /** 
    * @groupname axi3_4_config
    * MASTER:
    * Enables generation of exclusive access transactions.
    * <br>
    * SLAVE:
    * Indicates whether the slave supports exclusive access or not.
    * <b>type:</b> Static
    *
    */
  rand bit exclusive_access_enable = 0;
  
  /** 
    * @groupname ace_config
    * MASTER:
    * This is applicable only when svt_axi_port_configuration::exclusive_access_enable is set to 1.
    * This bit controls enabling  Exclusive Monitor for AXI and ACE Masters.
    * If it is set to '1' then exclusive monitor is enabled in ace masters cache is updated on successful exclusive transactions based on coherent response and exclusive monitor state.
    * If this is set to '0' then exclusive monitor is disabled in ace master and for exclusive transaction cache
    * is updated only based on coherent response i.e. if it is received as EXOKAY.
    * <b>type:</b> Dynamic
    */
  rand bit exclusive_monitor_enable = 1;

  /** 
    * @groupname axi3_4_config
    * MASTER:
    * Enables generation of locked access transactions.
    * <b>type:</b> Static
    *
    */
  rand bit locked_access_enable = 0;

  /** 
    * @groupname ace_config
    * MASTER:
    * Enables generation of barrier transactions.
    * <b>type:</b> Static
    */
  rand bit barrier_enable = 0;

  /** 
    * @groupname ace_config
    * MASTER:
    * Enables generation of DVM transactions.
    * <b>type:</b> Static
    */
  rand bit dvm_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only for active master 
    * Enables automated generation of DVMCOMPLETE transactions
    * in response to DVM Sync Snoop transactions. 
    * When this bit is unset, it is the user's responsibility to
    * send DVMCOMPLETE transactions from the sequence in response
    * to DVM Sync snoop transactions.
    * When this bit is set, the VIP master driver will auto generate 
    * DVMCOMPLETE transaction in response to DVM Sync snoop transactions.
    * When this bit is set, any DVMCOMPLETE transaction received from the sequencer will be ignored.
    */
  rand bit auto_gen_dvm_complete_enable = 0;

  /**
    * The minimum delay that needs to be applied to an auto-generated
    * DVM Complete transaction before it is processed by the driver
    * The delay is applied from the point that the DVM Sync snoop
    * transaction corresponding to the DVM COMPLETE ends. 
    */
  rand int min_auto_gen_dvm_complete_delay = 0;

  /**
    * The maximum delay that needs to be applied to an auto-generated
    * DVM Complete transaction before it is processed by the driver.
    * The delay is applied from the point that the DVM Sync snoop
    * transaction corresponding to the DVM COMPLETE ends. 
    */
  rand int max_auto_gen_dvm_complete_delay = `SVT_AXI_MAX_DVM_COMPLETE_DELAY;

  /**
    * If this parameter is set, when a DVM snoop sync is received, the driver
    * takes a snapshot of active transactions whose address or data have been
    * sent on the interface.  The DVMCOMPLETE on the read address channel is
    * then launched when these outstanding transactions are complete. The
    * parameter #dvm_complete_delay is not applicable if this parameter is set. 
    */
  bit launch_auto_gen_dvm_complete_on_outstanding_xact_completion = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE or ACE_LITE.
    *
    * MASTER:
    * Enables speculative read.
    * A speculative read is defined as a read of a cache line that a master may
    * already be holding in its cache. Consider a case when user generates a
    * coherent transaction for read of a cache line that a master already holds
    * in its cache.
    *
    * When speculative read is enabled, the master will transmit this coherent
    * transaction. Also, the master will support cache state transitions as
    * defined in second set of tables in sections 5.5.1 to 5.5.11 in ACE
    * proposal 0.27.
    *
    * When speculative read is disabled, the master will not transmit this
    * coherent transaction. In this case, the master will only support cache
    * state transitions as defined in first set of tables in sections 5.5.1 to
    * 5.5.11 in ACE proposal 0.27.
    *
    * Whether a transaction is a speculative read is indicated by read-only
    * transaction class member svt_axi_transaction::is_speculative_read.
    *
    * <b>type:</b> Dynamic
    */
  rand bit speculative_read_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE or ACE_LITE.
    *
    * MASTER:
    * Enables restrictions in the master for support of an external
    * snoop filter.
    * <b>type:</b> Dynamic
    */
  rand bit snoop_filter_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE_LITE.
    *
    * SLAVE:
    * Checks that cache maintenance transactions received by an interconnect
    * from a master are forwarded to corresponding slaves. This check will
    * be performed only if the system monitor is enabled and correlation of
    * master and slave transactions are enabled by setting 
    * id_based_correlation_enable in svt_axi_system_configuration and the associated
    * configuration properties. 
    * <b>type:</b> Dynamic
    */
  rand bit forward_cmos_to_slaves_check_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE or ACE_LITE.
    * MASTER:
    * Determines the permissible cache line state transitions in the master.
    * For each transaction type, the section 5 of the specification provides 
    * cache line state transitions for "expected (or recommended) end state", 
    * "legal end state with snoop filter" and "legal end state without snoop filter".  
    * This parameter determines which of the above state changes are to be
    * used.
    *
    * Below are the supported values:
    * - RECOMMENDED_CACHE_LINE_STATE_CHANGE: The cache line state
    * changes as given in the "expected end state" of each table is used.
    * - LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE: The cache 
    * line state changes as given in the "legal end state with snoop filter" 
    * of each table is used. To be able to use this cache line state transition,
    * the configuration member svt_axi_port_configuration::snoop_filter_enable
    * must be set to 1. The actual cache line state change can be done using
    * member svt_axi_transaction::force_to_shared_state.
    * - LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE: The cache 
    * line state changes as given in the "legal end state without snoop filter" 
    * of each table is used. To be able to use this cache line state transition,
    * the configuration member svt_axi_port_configuration::snoop_filter_enable
    * must be set to 0. The actual cache line state change can be done using
    * members svt_axi_transaction::force_to_invalid_state and
    * svt_axi_transaction::force_to_shared_state.
    * .
    *
    * <b>type:</b> Dynamic
    */
  rand axi_cache_line_state_change_type_enum cache_line_state_change_type = RECOMMENDED_CACHE_LINE_STATE_CHANGE;

  /**
   * @groupname ace_config
   * Applicable only when svt_axi_port_configuration::axi_interface_type is set to ACE and it is Master component.
   *
   * Specifies how master will process incoming snoop request when memory update transaction is in progress.
   * if it is set to SUSPEND_SNOOP_DURING_MEM_UPDATE then master will suspend incoming snoop request and will respond
   * after current memory update transaction is complete. This is the default response mode.
   * If it is set to RESPOND_SNOOP_DURING_MEM_UPDATE then master will not suspend incoming snoop request. Instead it will
   * respond to the incoming snoop request as allowed by ACE specification.
   * If it is set to EITHER_RESPOND_OR_SUSPEND_SNOOP_DURING_MEM_UPDATE then master will randomly decide to choose between
   * either of the above two behaviour i.e. either suspend incoming snoop or respond to it.
   * 
   * Configuration type: Dynamic
   */
  rand snoop_response_mode_during_mem_update_type_enum snoop_response_mode_during_mem_update = SUSPEND_SNOOP_DURING_MEM_UPDATE;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is set to ACE and it is Master component
    *
    * Indicates how dirty data in cache should be transferred on receiving a snoop.
    * As per section C5.2.2 of the AXI specification, a cached master can ensure that data in a dirty cacheline
    * is available to a snoop other than MAKEINVALID in one of two ways:
    * 1. returning data when the master completes the snoop
    * 2. carrying out a memory update, using a WRITEBACK or WRITECLEAN before responding to the snoop
    * This configuration indicates which of the above two methods will be used for returning data
    * Note that if there is an outstanding WRITEUNIQUE or WRITELINEUNIQUE transaction in the
    * queue of the master, then data will be returned with the snoop transaction. This is to comply with
    * restrictions on WRITEUNIQUE and WRITELINEUNIQUE while a snoop is in progress as per section
    * C4.8.7 of the spec
    */
  rand snoop_response_data_transfer_mode_enum snoop_response_data_transfer_mode = SNOOP_RESP_DATA_TRANSFER_USING_CDDATA;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE and it is Master component
    *
    * Describes various address randomization mode for nonshareable transaction with domain type SYSTEMSHAREABLE. It indicates what
    * address range should or shouldn't be used while randomizing axi master transaction based on the different enum values listed below.
    *
    * NONSHAREABLE_XACT_FULL_ADDRESS_SPACE :: allows full address sapce to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE :: allows only address sapce outside inner, outer or nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * NONSHAREABLE_XACT_ADDR_WITHIN_NON_SHAREABLE_ADDR_RANGE :: allows only nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_ADDR_RANGE :: allows only address sapce outside inner or outer address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * default value :: NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE
    */
  rand nonshareable_xact_address_range_in_systemshareable_mode_enum nonshareable_xact_address_range_in_systemshareable_mode = NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE;

  /**
    * @groupname axi3_4_config
    * MASTER:
    * The maximum number of active exclusive transactions that will be initiated by the master.
    * SLAVE:
    * The maximum number of active exclusive access monitors supported by the slave. Attempts to
    * exceed this max number results in a failed exclusive access read response of OKAY instead of EXOKAY.
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_NUM_EXCLUSIVE_ACCESS
    * NOTE: if it is set to '0' value then there are no restrictions on maximum number of active exclusive
    * transactions. VIP will not mark any exclusive sequence as failed because of this parameter.
    * <b>type:</b> Static
    */ 
  rand int max_num_exclusive_access   = `SVT_AXI_MAX_NUM_EXCLUSIVE_ACCESS;
      
  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE
    * INTERCONNECT:
    * Number of ADDRESS bits that need to be monitored by the exclusive monitors for 
    * current port in order to support one or more independent exclusive access
    * thread.
    *
    * It can also be configured with ( -1 ) to indicate that address ranges for 
    * each exclusive monitor is defined through user specified start and end address ranges.
    * For this, user should configure start_address_ranges_for_exclusive_monitor[] and
    * end_address_ranges_for_exclusive_monitor[] arrays in system configuration.
    * A svt_axi_system_configuration::set_exclusive_monitor_addr_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr,
    *     bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr) utility method can be used for this purpose.
    *
    * NOTE: configuring with value 0 means, no address is being monitored by the 
    * corresponding exclusive monitor and hence exclusive access to different address
    * may also affect current thread.
    *
    * <b>specail value:</b> -1 indicates that num_addr_bits_used_in_exclusive_monitor and
    * num_initial_addr_bits_ignored_by_exclusive_monitor are not used. Instead address
    * ranges for exclusive monitors are defined by address_ranges_for_exclusive_monitor[] array.
    *
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_ADDR_WIDTH-1
    * <b>type:</b> Static
    */ 
  rand int num_addr_bits_used_in_exclusive_monitor   = `SVT_AXI_MAX_ADDR_WIDTH;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE
    * ACE Exclusive monitor will ignore number of initial address bits as
    * indicated by this configuration member.
    * Example: A coherent interconnect can divide its whole address space into
    *          multiple ranges such that each PoS Exclusive monitor checks only
    * its corresponding address range. So, if it allocates 1/2 GB address space to each
    * of the 4 PoS exclusive monitors then num_initial_addr_bits_ignored_by_exclusive_monitor
    * needs to be configured as 29 (1.5GB - 2GB ~ 31 bits).
    */
  rand int num_initial_addr_bits_ignored_by_exclusive_monitor   = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE
    * INTERCONNECT:
    * Number of ID bits that need to be monitored by the exclusive monitors for 
    * current port in order to support one or more independent exclusive access
    * thread.
    * NOTE: configuring with value 0 means, no id is being monitored by the 
    * corresponding exclusive monitor and hence only single exclusive access thread
    * is supported for current port.
    *  <b> This feature is not supported yet </b>
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_ID_WIDTH-1
    * <b>type:</b> Static
    */ 
  rand int num_id_bits_used_in_exclusive_monitor     = `SVT_AXI_MAX_ID_WIDTH;

   /*
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE
    * INTERCONNECT:
    * Indicates whether Interconnect uses seperate PoS Exclusive Monitor for 
    * secured or non-secured exclusive access.
    * NOTE: configuring with value 0 means, interconnect doesn't monitor seperately
    * for secured or unsecured exclusive access.
    * <b> This feature is supported by enabling secure address space by configuring tagged_address_space_attributes_enable = 1 </b>
    * <b> User shouldn't use this configuration parameter, it is going to be deprecated </b> 0
    * <b>min val:</b> 0
    * <b>max val:</b> 1
    * <b>type:</b> Static
    */ 
  rand bit use_secured_exclusive_monitor             = 1;

  /**
    * @groupname ace_config
    * If set to '1' then VIP will not assert error if Master sends Exclusive Store without sending Exlusive Load.
    * However, if Exclusive Store is sent from the Invalid cacheline state then VIP will still assert error since,
    * that is not a valid state to start Exclusive Store.
    * <b>type:</b> Static
    */ 
  rand bit allow_exclusive_store_without_exclusive_load = 0;

  /**
    * @groupname ace_config
    * If set to '1' then VIP will respond to very first Exclusive Store with EXOKAY response. This means that if
    * no master has performed any exclusive transaction after reset is de-asserted then the master that issues
    * exclusive store will be responded with EXOKAY or VIP will expect EXOKAY response from the coherent interconnect.
    * Note: reference point of first exclusive store is reset.
    * <b>type:</b> Static
    */ 
  rand bit allow_first_exclusive_store_to_succeed = 0;

  /**
    * @groupname ace_config
    * If set to '1' then Exclusive Monitor will get reset once Exclusive Store is successful.
    * If set to '0' then Exclusive Monitor will remain set even if Exclusive Store is successful.
    * Please Note that, VIP will still reset Exclusive Monitor for failed Exclusive Store attempt
    * regardless of the value set for this parameter.
    * <b>type:</b> Static
    */ 
  rand bit reset_exclusive_monitor_on_successful_exclusive_store = 1;

  /**
    * @groupname ace_config
    * This control register indicates different modes of error conditions uded in exclusive monitor.
    * [0] => If set to '1' implies that Snoop Error will cause an exclusive sequence to fail only if
    *        either data_transfer bit or pass_dirty bit is set to '1'. Otherwise, if snoop response
    *        indicates error bit as asserted then regardless of data_transfer bit or pass_dirty bit
    *        values exclusive sequence will fail. 
    * [31:1] => Reserved bits.
    * Default Value :: 0x00000000
    */
  rand bit[31:0] exclusive_monitor_error_control_reg = 0;

  /** 
    * @groupname ace_config
    * If shareable exclusive access needs to be supported from ace-lite port then this parameter
    * should be set to '1'. If it is set to '1' then VIP will allow READONCE or WRITEUNIQUE
    * transactions to be of exclusive type.
    * Default Value: '0' i.e. shareable exclusive access from ace-lite port is not allowed. Only
    *                non-shareable exclusive transactions as READNOSNOOP or WRITENOSNOOP are allowed.
    */
  rand bit shareable_exclusive_access_from_acelite_ports_enable = 1;

  /**
    * @groupname axi3_4_config
    * Specifies the number of write transactions that can be interleaved
    * This parameter should not be greater than #num_outstanding_xact.
    * When set to 1, interleaving is not allowed.
    * MASTER: 
    * Does not interleave transmitted write data beyond this value.
    * SLAVE: 
    * Checks that received write data is not interleaved beyond this value. 
    * An error is issued if write data is interleaved 
    * beyond this value.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_WR_INTERLEAVE_DEPTH
    * <b>type:</b> Static
    */ 
  rand int write_data_interleave_depth       = `SVT_AXI_MAX_WR_INTERLEAVE_DEPTH;

  /** 
    * @groupname axi3_4_config
    * This parameter specifies the atomicity size required to check the address
    * alignment for a given transcation as per the atomicity of component.<br>
    * This parameter will not have effect if set to -1. The values specified
    * to this parameter should be power of 2, in terms of Bytes <br>
    * Default value: -1.<br>
    * Allowed values: should be power of 2, in terms of Bytes. <br>
    * For example: 8, 16, 32, 64 etc <br>
    * <b>type:</b> Static
    *
    */
  rand int atomicity_size = -1;


  /** @cond PRIVATE */
  /**
    * When set to 1, enables id reflection in AXI4_LITE mode.
    * This enables the awid, bid and rid signals. This allows
    * an AXI4-Lite slave to be used on a full AXI interface,
    * without a bridge function, in a system that guarantees that
    * the slave can only be accessed by transactions that fall
    * within the AXI4-Lite subset.
    * <b>type:</b> Static
    *
    * This parameter is not yet supported.
    */
  rand bit id_reflection_enable = 0;
  /** @endcond */

  /**
    * @groupname axi3_4_config
    * Applicable only to MASTER when axi_interface_type is 
    * AXI3/AXI4/AXI4_LITE.
    * When set to 1, accesses to the read address channel and 
    * write address channel are serialized. Thus, awvalid and
    * arvalid will never be asserted at the same time. The
    * address information driven on the write address channel
    * will have to be accepted before any address information
    * on the read address channel is driven and viceversa. 
    * When set to 0, activity on the read address channel and
    * write address channel occur in parallel.
    */
  rand bit serial_read_write_access = 0;

`ifndef SVT_EXCLUDE_VCAP
  /**
    * @groupname axi_traffic_profile 
    * Enables use of traffic profiles. This enables the use of transaction
    * generation at a higher level of abstraction.  This feature
    * is only available as part of the NOC product. Please refer to the NOC
    * user guide for details
    */
  bit use_traffic_profile = 0;

  /** 
    * @groupname axi_generic_config
    * Enables FIFO based rate control. 
    * A FIFO is modelled in the driver for read and write
    * transactions separately. A WRITE transaction can be sent
    * out if there is sufficient data in the FIFO to send out that
    * transaction. A READ transaction can be sent out if there is
    * space in the FIFO to receive the data of the READ transaction.
    * The current level of a WRITE FIFO is incremented every clock
    * based on write_fifo_fill_rate.With every data beat, the currentl level
    * is decremented based on burst_size of the transaction. The current level of a READ FIFO
    * is decremented every clock based on read_fifo_drain_rate. With every data
    * beat, the current level is incremented based on burst_size of the transaction.
    * A WRITE transaction will be sent out if the current level is greater than
    * the total number of bytes of all outstanding write transactions + the total
    * number of bytes of the current transaction. A READ transaction will be sent out
    * if the current level is less than the difference of the read_fifo_full_level and
    * the total number of bytes of all outstanding read transactions + the total number
    * of bytes of the current transaction.
    */
  rand bit use_fifo_based_rate_control = 0;

  /**
    * @groupname axi_generic_config
    * Clock period in ns. This is used to calculate the drain/fill rate in
    * bytes/cycle
    */
  real clock_period = 1;

  /** 
    * @groupname axi_generic_config
    * The drain rate in MBPS of the FIFO into which data from READ
    * transactions is dumped. Used by the check_current_fill_level_read_fifo 
    * method of the corresponding driver to determine if there is space
    * in the FIFO to receive data of a READ transaction
    */
  rand int read_fifo_drain_rate = `SVT_AXI_MAX_READ_FIFO_DRAIN_RATE;

  /** 
    * @groupname axi_generic_config
    * The full level in bytes of the READ FIFO into which data from READ transactions
    * is dumped. Used by the check_current_fill_level_read_fifo 
    * method of the corresponding driver to determine if there is space
    * in the FIFO to receive data of a READ transaction.
    */
  rand int read_fifo_full_level = `SVT_AXI_MAX_READ_FIFO_FULL_LEVEL;

  /** 
    * @groupname axi_generic_config
    * The fill rate in MBPS of the FIFO from which data for WRITE 
    * transactions is taken. Used by the check_current_fill_level_write_fifo 
    * method of the corresponding driver to determine if there is enough 
    * data in the FIFO to send a WRITE transaction
    */
  rand int write_fifo_fill_rate = `SVT_AXI_MAX_WRITE_FIFO_FILL_RATE;

  /** 
    * @groupname axi_generic_config
    * The full level in bytes of the WRITE FIFO from which data for WRITE transactions
    * is taken. Used by the check_current_fill_level_write_fifo 
    * method of the corresponding driver to determine if there is enough 
    * data in the FIFO to transmit data of a WRITE transaction
    */
  rand int write_fifo_full_level = `SVT_AXI_MAX_WRITE_FIFO_FULL_LEVEL;

  /**
    * @groupname axi_generic_config
    * Determines if the READ FIFO is empty on start up
    */
  rand bit is_read_fifo_empty_on_start = 1;

  /**
    * @groupname axi_generic_config
    * Determines if the WRITE FIFO is empty on start up
    */
  rand bit is_write_fifo_empty_on_start = 1;
`endif //SVT_EXCLUDE_VCAP

  /** 
    * @groupname axi_generic_config
    * If this parameter is set, AXI transaction phase level information is
    * printed in note verbosity.  Messages related to start & end of address,
    * data and response phases are printed.  If unset, AXI transaction phase
    * level information is printed only in debug verbosity.
    */ 
  bit display_xact_phase_messages = 0;

  /** 
    * @groupname axi_generic_config
    * If this parameter is set, maximum number of outstanding transactions
    * per AxID is limited to 1 for Non-Device and Non-DVM transactions.
    * This can be further controlled by configuration
    * svt_axi_port_configuration::single_outstanding_per_id_kind. 
    */ 
  bit single_outstanding_per_id_enable = 0; 

  /** 
    * @groupname axi_generic_config
    * If this parameter is set, maximum number of outstanding AXI4_STREAM transactions
    * per TDEST is limited to 1.
    */ 
  bit single_outstanding_per_tdest_enable = 0; 

  /** 
    * @groupname axi_generic_config
    * If this parameter is set to 1, all delay related parameters will be set
    * to 0. Note however, that actual delay on interface will vary based on
    * outstanding transactions.
    */ 
  rand bit zero_delay_enable = 0; 
  
  /**
    * This enumerated type controls the AxID when
    * svt_axi_port_configuration::single_outstanding_per_id_enable is set to 1.
    *
    * If svt_axi_port_configuration::single_outstanding_per_id_kind is set to
    * 'MODIFY_SAME_ID': If AxID of a new Non Device or Non DVM transaction matches
    * AxID of an active transaction, the VIP modifies the AxID such that the AxID 
    * is not overlapping with AxID of any active Non Device or Non DVM transactions.
    *
    * For example, a new Non Device or Non DVM transaction with AxID = 6 is initiated
    * by the user sequence. At this time, another Non Device or Non DVM with AxID = 6
    * is already in progress. In this case, VIP will check the active queue, and modify
    * the AxID of the new transaction to an un-used AxID. For example, VIP will modify 
    * the AxID of new transaction to 4, if this is not used by any active transactions.
    * 
    * If svt_axi_port_configuration::single_outstanding_per_id_kind is set to
    * ‘WAIT_FOR_COMPLETION_OF_SAME_ID': If AxID of a new Non Device or Non DVM transaction
    * matches AxID of an active Non Device or Non DVM transaction, the VIP waits till the
    * corresponding active Non Device or Non DVM transaction is complete. Only when the
    * active Non Device or Non DVM transaction is complete, VIP adds the new Non Device
    * or Non DVM transaction to the active queue. This ensures that only 1 active Non Device
    * or Non DVM transaction exists for a given AxID.
    *
    * For example, a new Non Device or Non DVM transaction with AxID = 6 is initiated by
    * the user sequence. At this time, another Non Device or Non DVM with AxID = 6 is already
    * in progress. In this case, VIP will wait for the active transaction to complete. After
    * active transaction is complete, VIP will add the new transaction with AxID = 6 to the
    * active queue.
    */
  typedef enum {
    MODIFY_SAME_ID = 0,
    WAIT_FOR_COMPLETION_OF_SAME_ID = 1
  } single_outstanding_per_id_kind_enum;

  single_outstanding_per_id_kind_enum single_outstanding_per_id_kind = WAIT_FOR_COMPLETION_OF_SAME_ID;

  /**
    * If this parameter is set, debug information is driven on the debug ports.
    * The transaction id as well as the transfer id corresponding to 
    * each beat is driven on the debug ports.
    *
    * 
    *
    * <b>type:</b> Static
    */
  bit use_debug_interface = 0; 



  /**
    * @groupname axi_coverage_protocol_checks
    * Enables protocol checking. In a disabled state, no protocol
    * violation messages (error or warning) are issued.
    * <b>type:</b> Dynamic 
    */
  bit protocol_checks_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables protocol check statistics collection. In a disabled state, statistics 
    * on checks executed are not collected. Enabling this has a run-time performance impact
    * <b>type:</b> Dynamic 
    */
  bit protocol_check_stats_enable = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables toggle coverage.
    * Toggle Coverage gives us information on whether a bit
    * toggled from 0 to 1 and back from 1 to 0. This does not
    * indicate that every value of a multi-bit vector was seen, but
    * measures if individual bits of a multi-bit vector toggled.
    * This coverage gives information on whether a system is connected
    * properly or not.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit toggle_coverage_enable = 1;
  `else
  bit toggle_coverage_enable = 0;
  `endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables state coverage of signals.
    * State Coverage covers all possible states of a signal.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit state_coverage_enable = 1;
  `else
  bit state_coverage_enable = 0;
  `endif


  /** @cond PRIVATE */
  /**
    * Enables meta coverage of signals.
    * This covers second-order coverage data such as valid-ready
    * delays.
    * <br>
    * This parameter is not supported currently. The meta coverage is enabled
    * using port configuration parameter #transaction_coverage_enable.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit meta_coverage_enable = 1;
  `else
  bit meta_coverage_enable = 0;
  `endif

  /** @endcond */

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables transaction level coverage. This parameter also enables delay
    * coverage. Delay coverage is coverage on various delays between valid & ready signals.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit transaction_coverage_enable = 1;
  `else
  bit transaction_coverage_enable = 0;
  `endif
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables protocol checks coverage. 
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit protocol_checks_coverage_enable = 1;
  `else
  bit protocol_checks_coverage_enable = 0;
  `endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables positive or negative protocol checks coverage. 
    * When set to '1', enables positive protocol checks coverage.
    * When set to '0', enables negative protocol checks coverage.
    * <b>type:</b> Static 
    */
  bit pass_check_cov = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables signal valid check during reset when protocol_checks_enable=1. 
    * When set to '1', enables signal valid check during reset.
    * When set to '0', disables signal valid check during reset. In a disabled
    * state, no signal valid check during reset violation messages (error or warning) are issued.
    * <b>type:</b> Static 
    */
  bit signal_valid_during_reset_checks_enable = 1;
 
  /**
    * @groupname axi_coverage_protocol_checks
    * ID value used for matching outstanding read/write transactions for
    * covergroups trans_axi_num_outstanding_xacts_with_same_awid and 
    * trans_axi_num_outstanding_xacts_with_same_arid. 
    * <b>type:</b> Static 
    */
  int cov_same_id_in_outstanding_xacts = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Set of multiple ID values used for matching outstanding read/write transactions for
    * covergroups trans_axi_num_outstanding_xacts_with_multiple_same_arid and 
    * trans_axi_num_outstanding_xacts_with_multiple_same_awid. 
    * <b>type:</b> Static 
    */
  int cov_multi_same_ids[];

  /**
    * @groupname axi_coverage_protocol_checks
    * ID value used for matching back to back write transactions for
    * covergroups trans_master_ace_lite_coherent_and_ace_snoop_response_association_with_specific_id. 
    * <b>type:</b> Static 
    */
  int cov_specific_id_in_back_to_back_xacts = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables valid_ready_dependency_coverage 
    * <b>type:</b> Static 
    */
  // When valid_ready_dependency_coverage_enable is set to '1' for IUS simulator
  // the function cov_sample_``dependency () of svt_axi_port_monitor_def_cov_util.svi
  // consumes around 10x more time. So because of this, the default value is kept 0 for the IUS simulator.
  // valid_ready_dependency covergroups as performance intensive and hence diabling them by default.
`ifndef INCA
  bit valid_ready_dependency_coverage_enable= 0;
`else 
  bit valid_ready_dependency_coverage_enable= 0;
`endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * wvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * rready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_rready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * bready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_bready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * awvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_awvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * rready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_rready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * bready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_bready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * awvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_awvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * wvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * bready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_bready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * awvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_awvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * wvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * rready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_rready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * arready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_arready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_rvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which arready need to be deasserted after
    * wready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_arready_wready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which arready need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_arready_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which arready need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_arready_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * arready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_arready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * wready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * arready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_arready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid  need to be deasserted after
    * wready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_wready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_bvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_wready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_rvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_bvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * awvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awready_and_awvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * wvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */ 
  int cov_num_clks_awready_and_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awready_and_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awready_and_bvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * awvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_awvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * wvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_wvalid_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * rready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_rready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * bready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_bready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * awready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_awready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * wready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_wready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * rready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_rready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * bready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_bready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * awready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_awready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * wready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_wready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * rready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_rready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * bready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_bready_dependency  = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates the number of bins which will be created for covergroups
    * trans_axi_num_outstanding_xacts_with_same_awid and 
    * trans_axi_num_outstanding_xacts_with_same_arid.
    * It should be programmed to a value less than or equal to configured value of 
    * svt_axi_port_configuration::num_outstanding_xact or 
    * svt_axi_port_configuration::num_write_outstanding_xact if 
    * svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    * indicates the number of outstanding transactions VIP can support.
    * If user does not program this variable it will create 64 bins each for 
    * covergroups trans_axi_num_outstanding_xacts_with_same_awid and 
    * trans_axi_num_outstanding_xacts_with_same_awid
    * <b>type:</b> Static 
    */
  int cov_bins_num_outstanding_xacts = 64;

  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates the number of bins which will be created for covergroup
    * trans_ace_num_outstanding_snoop_xacts.It should be programmed to 
    * a value less than or equal to configured value of 
    * svt_axi_port_configuration::num_outstanding_snoop_xact which
    * indicates the number of outstanding snoop transactions VIP can support.
    *
    * If user does not program this variable it will create 64 bins for 
    * covergroup trans_ace_num_outstanding_snoop_xact
    * <b>type:</b> Static 
    */
  int cov_bins_num_outstanding_snoop_xacts = 64;

  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates the number of bins which will be created for covergroup
    * trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid.
    * It should be programmed to a value less than or equal to configured value of 
    * svt_axi_port_configuration::num_outstanding_xact or 
    * svt_axi_port_configuration::num_read_outstanding_xact if 
    * svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    * indicates the number of outstanding transactions VIP can support.
    * If user does not program this variable it will create 64 bins for 
    * covergroup trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid 
    * <b>type:</b> Static 
    */
  int cov_bins_dvm_tlbi_num_outstanding_xacts = 64;  

  /**
    * @groupname axi_coverage_protocol_checks
    * ID value used for matching outstanding DVM TLBI transactions for
    * covergroup trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid. 
    * <b>type:</b> Static    
    */
  int cov_same_id_in_dvm_tlbi_outstanding_xacts = 0;  
  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates if user wants to cover all the id_ranges of the outstanding
    * transactions. BY default , Only fixed number of outstanding transactions will be covered 
    * <b>type:</b> Static 
    */
  bit cov_num_outstanding_xacts_range_enable = 0;  

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awaddr signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and bresp signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_bresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awprot signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and araddr signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_araddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and rresp signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_rresp_enable = 1;
    /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic_type,rresp signal.
    * <b>type:</b> Dynamic 
    */
  bit trans_cross_axi_atomictype_rresp_enable = 1;

 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic_type,bresp signal.
    * <b>type:</b> Dynamic 
    */
  bit trans_cross_axi_atomictype_bresp_enable = 1;



  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arprot signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst,
    * awlen, awaddr and awsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awaddr_awsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst,
    * awlen and awsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst and
    * awlen signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awlock signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awlock_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awcache signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst,
    * arlen, araddr and arsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_araddr_arsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arlock signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arlock_enable = 1;

`ifdef SVT_ACE5_ENABLE
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type,atomic_xact_op_type,awsize
    * and awburst signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_atomic_comp_awburst_awsize_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type , atomic xact op type , awburst
    * and awsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_atomic_noncomp_awburst_awsize_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type , bresp and
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_comp_bresp_burst_length_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type ,bresp
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_noncomp_bresp_burst_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type , rresp 
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_comp_rresp_burst_length_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type , rresp 
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_noncomp_rresp_burst_length_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type
    * and endianness.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_comp_endianness_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type 
    * and endianness.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_noncomp_endianness_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between write transaction type , awmmussid and
    * and awmmusecsid signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_write_xact_type_awmmusecsid_awmmussid_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between write_xact_type , awmmussidv and awmmussid signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_write_xact_type_awmmussidv_awmmussid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between read_xact_type,armmusecsid and armmusid signal.
    * <b>type:</b> Static 
    */
bit trans_cross_read_xact_type_armmusecsid_armmusid_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between read_xact_type , armmussidv
    * and armmussid signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_read_xact_type_armmussidv_armmussid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between coherent stash transaction type , stash_nid
    * and stash_nid_valid.
    * <b>type:</b> Static 
    */
bit trans_cross_stash_xact_type_stash_nid_stashnid_valid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between coherent stash transaction type , stash_lpid
    * and stash_lpid_valid.
    * <b>type:</b> Static 
    */
bit trans_cross_stash_xact_type_stash_lpid_stashlpid_valid_enable = 1;

`endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst and
    * arlen signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arcache signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst and
    * awqos signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awqos_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst and 
    * arqos signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arqos_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awburst signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awburst_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awlen signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awlen_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awsize signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awaddr signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * bresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_bresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop, awdomain 
    * and bresp signal.
    * The EXOKAY response is permitted for WriteNoSnoop for NONSHAREABLE and SYSTEMSHAREABLE domains. 
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_awsnoop_awdomain_bresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks    
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awdomain signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awdomain_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks    
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awdomain and awcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awdomain_awcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awbar signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awbar_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awbarrier (MEMORY_BARRIER and SYNC_BARRIER) and 
    * awdomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_awdomain_awbarrier_memory_sync_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awbarrier (NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER) and 
    * awdomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_awdomain_awbarrier_respect_ignore_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arbarrier (MEMORY_BARRIER and SYNC_BARRIER) and 
    * ardomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_ardomain_arbarrier_memory_sync_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arbarrier (NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER) and 
    * ardomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_ardomain_arbarrier_respect_ignore_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks    
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arburst signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arburst_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arlen signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arlen_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arsize signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * araddr signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_araddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * rresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_coh_rresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * ardomain signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_ardomain_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * ardomain and arcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_ardomain_arcache_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arbar signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arbar_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between ardvmmessage and 
    * ardvmresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_ardvmmessage_ardvmresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop and 
    * acaddr signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_acaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop and 
    * acprot signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_acprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop and 
    * ace rresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_crresp_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acdvmmessages
    * and acdvmresp.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acdvmmessage_acdvmresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop
    * initial cache line status and final cache line status.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop
    * initial cache line status and final cache line status.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_cacheinitialstate_cachefinalstate_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop
    * initial cache line status and final cache line status.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_cacheinitialstate_cachefinalstate_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level meta coverage group for read transfer
    * <b>type:</b> Static 
    */
  bit trans_meta_axi_read_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level meta coverage group for write transfer
    * <b>type:</b> Static 
    */
  bit trans_meta_axi_write_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI4 STREAM transaction level meta coverage group for axi4 stream transfer
    * <b>type:</b> Static 
    */
  bit trans_meta_axi4_stream_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI4 STREAM transaction level delay coverage group for axi4 stream transfer
    * <b>type:</b> Static 
    */
  bit trans_axi4_stream_delay_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level out-of-order response coverage group for read transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_ooo_read_response_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level out-of-order response coverage group for write transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_ooo_write_response_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI STREAM transaction level coverage group for cross coverage
    * between stream transaction type, tid and tdest.
    * <b>type:</b> Static 
    */
  bit trans_cross_stream_xact_type_tid_tdest_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for axi outstanding transaction
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_outstanding_xact_enable = 1;
  
  /**
    * @groupname ace_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_barrier_outstanding_xact coverage group for
    * axi barrier outstanding transaction
    * <b>type:</b> Static 
    */
  bit trans_ace_barrier_outstanding_xact_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_barrier_pair_sequence coverage group for
    * read and write barrier pair transaction
    * <b>type:</b> Static 
    */
  bit trans_ace_barrier_pair_sequence_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables AXI transaction level trans_non_barrier_xact_after_256_outstanding_barrier_xact coverage group
    * <b>type:</b> Static 
    */
  bit trans_non_barrier_xact_after_256_outstanding_barrier_xact_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_back_to_back_read_burst_sequence coverage group for
    * back to back read pair transaction
    * <b>type:</b> Static 
    */
  bit trans_axi_back_to_back_read_burst_sequence_enable = 1;

 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_back_to_back_write_burst_sequence coverage group for
    * back to back write pair transaction
    * <b>type:</b> Static 
    */
  bit trans_axi_back_to_back_write_burst_sequence_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_write_read_same_id_completed_out_of_order coverage group for
    * WRITE/READ transactions with same ID completed OOO
    * <b>type:</b> Static 
    */
  bit trans_axi_write_read_same_id_completed_out_of_order_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_write_read_diff_id_completed_out_of_order coverage group for
    * WRITE/READ transactions with diff ID completed OOO
    * <b>type:</b> Static 
    */
  bit trans_axi_write_read_diff_id_completed_out_of_order_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width48 ,
    * trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width40,trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width32,
    * trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_tlbinvl_modes_virtaddr_cov_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width48  ,
    * trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width40,trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width32,
    * trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_branch_predictor_invl_modes_cov_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for  trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width48,
    * trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width40,trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width32,
    * trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_phy_inst_cache_invl_modes_modes_cov_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width48,
    * trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width40,trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width32
    * trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_virt_inst_cache_invl_modes_cov_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_firstpart_addr_range_width48,
    * trans_cross_ace_dvm_firstpart_addr_range_width40,trans_cross_ace_dvm_firstpart_addr_range_width32,
    * trans_cross_ace_dvm_firstpart_addr_range_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_firstpart_addr_range_cov_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_firstpart_secondpart_addr_range_width65,
    * trans_cross_ace_dvm_firstpart_secondpart_addr_range56,trans_cross_ace_dvm_firstpart_secondpart_addr_range32
    * trans_cross_ace_dvm_firstpart_secondpart_addr_range24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_firstpart_secondpart_addr_range_cov_enable = 1;
  
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_four_state_RD_WR_burst_sequence coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_four_state_rd_wr_burst_sequence_cov_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_four_excl_normal_sequence coverage group
    * This cover group covers specific combinations of exclusive and normal transactions
    * <b>type:</b> Static 
    */

  bit trans_axi_four_excl_normal_sequence_cov_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_lock_followed_by_excl_sequence coverage group
    * <b>type:</b> Static 
    */
  bit trans_lock_followed_by_excl_sequence_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_fixed_burst_wstrb coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_fixed_burst_wstrb_cov_enable = 1; 
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer coverage group 
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_cov_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_cov_enable coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_cov_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_wstrb_to_signal_unaligned_start_address coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_wstrb_to_signal_unaligned_start_address_cov_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_read_outstanding_xact_same_arid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_read_outstanding_xact_same_arid_cache_modifiable_bit_enable = 1;
   
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_read_outstanding_xact_diff_arid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_read_outstanding_xact_diff_arid_cache_modifiable_bit_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_read_outstanding_xact_diff_arid_device_cacheable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_read_outstanding_xact_diff_arid_device_cacheable_bit_enable = 1;
   
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_write_outstanding_xact_same_awid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_write_outstanding_xact_same_awid_cache_modifiable_bit_enable = 1;
   
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_write_outstanding_xact_diff_awid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_write_outstanding_xact_diff_awid_cache_modifiable_bit_enable = 1;
 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_write_outstanding_xact_diff_awid_device_cacheable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_write_outstanding_xact_diff_awid_device_cacheable_bit_enable = 1;
 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_same_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_same_arid_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_multiple_same_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_multiple_same_arid_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level
    * trans_axi_num_outstanding_xacts_with_multiple_same_awid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_multiple_same_awid_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_arid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_arid_range coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_arid_range_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_same_awid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_same_awid_enable = 1;

 
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_awid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_awid_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_awid_range coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_awid_range_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_snoop_xacts coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_snoop_xacts_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_enable = 1;  
/**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_enable = 1;  

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_atomictype_exclusive_arcache coverage group
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_atomictype_exclusive_arcache_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_atomictype_exclusive_awcache  coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_atomictype_exclusive_awcache_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_awsnoop_awdomain_awprot coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_writeunique_awdomain_awprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables cross coverage of  transaction parameters with slave port_id for
    * the following covergroups.
    * - trans_cross_ace_awsnoop_awsize
    * - trans_cross_ace_arsnoop_arsize
    * - trans_cross_ace_awsnoop_awlen
    * - trans_cross_ace_arsnoop_arlen
    * - trans_cross_ace_awsnoop_awdomain
    * - trans_cross_ace_arsnoop_ardomain
    * - trans_cross_ace_awsnoop_awcache
    * - trans_cross_ace_arsnoop_arcache
    * - trans_cross_ace_awsnoop_awburst
    * - trans_cross_ace_arsnoop_arburst
    * - trans_cross_ace_awsnoop_bresp
    * - trans_cross_ace_arsnoop_coh_rresp
    * Basically, it covers if the transaction properties have been covered from the master to all the different slaves
    * .
    * <b>type:</b> Static 
    */
  bit cov_trans_cross_slave_port_id_enable = 0;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_arsnoop_ardomain_arprot coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_readonce_ardomain_arprot_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_awprot_awbarrier_memory_sync coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_awprot_awbarrier_memory_sync_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_arprot_arbarrier_memory_sync coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_arprot_arbarrier_memory_sync_enable = 1;
      
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for write strobes 
    * <b>type:</b> Static 
    */  
  bit trans_cross_axi_write_strobes_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for write interleaving depth
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_write_interleaving_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for read interleaving depth
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_read_interleaving_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for write narror transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_write_narrow_transfer_awlen_awaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for read narror transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_read_narrow_transfer_arlen_araddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for unaligned write transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_write_unaligned_transfer_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for unaligned read transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_read_unaligned_transfer_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction coverage group for master_to_slave_path_access
    * <b>type:</b> Static 
    */
  bit trans_cross_master_to_slave_path_access_cov_enable = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_lite_coherent_and_ace_snoop_response_association
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_lite_coherent_and_ace_snoop_response_association_enable = 1;  

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_coherent_and_ace_snoop_response_association
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_coherent_and_ace_snoop_response_association_enable = 1;  
 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_lite_coherent_and_ace_snoop_response_association_specific_id
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_lite_coherent_and_ace_snoop_response_association_specific_id_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id_enable = 1;

  /** @cond PRIVATE */
   /**
    * @groupname master_slave_xact_association
    * In Master Slave transaction association flow, for non monifiable transaction cache_type 
    * and prot_type fields are compared.
    * By default this configuration parameter is set to 1 to enable cache_type and prot_type comparation,
    * if this parameter is set 0 then cache_type and prot_type comparations are dissabled
    * in master slave transaction association.
    * Note that to enable or dissable this feature, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit master_slave_xact_association_cache_prot_check_enable = 1;
  /** @endcond */

   /**
    * @groupname master_slave_xact_association
    * In Master Slave transaction association flow, cache_type[3:1] and prot_type fields are compared.
    * By default this configuration parameter is set to SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_NONMODIFIABLE_CHECK
    * to enable cache_type and prot_type comparation for non modifiable transaction,
    * if this parameter is set SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_MODIFIABLE_NONMODIFIABLE_CACHE_TYPE_CHECK
    * it enables cache_type and prot_type comparation for modifiable and non modifiable transactions,
    * in master slave transaction association.
    * Note that to enable or dissable this feature, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  master_slave_xact_association_cache_prot_check_enum master_slave_xact_association_cache_prot_check = SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_NONMODIFIABLE_CHECK;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for snoop transfer
    * <b>type:</b> Static 
    */
  bit trans_axi_snoop_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_outstanding_read_with_same_id_to_different_slaves
    * <b>type:</b> Static 
    */
  bit trans_outstanding_read_with_same_id_to_different_slaves_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_overlapping_arsnoop_acsnoop 
    * <b>type:</b> Static 
    */
  bit trans_ace_concurrent_overlapping_arsnoop_acsnoop_enable =1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_enabled 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_disabled
    * <b>type:</b> Static 
    */
  bit trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_enable =1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp 
    * <b>type:</b> Static 
    */
  bit trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_enable =1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_outstanding_read_with_same_id_to_different_slaves
    * <b>type:</b> Static 
    */
  bit trans_outstanding_write_with_same_id_to_different_slaves_enable = 1;
  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transactions on
    * AR, AW channel waiting for snoop response
    * <b>type:</b> Static 
    */
  bit trans_ar_aw_stalled_for_ac_channel_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after nonshareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_nonshareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after innershareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_innershareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after outershareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_outershareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after systemshareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_systemshareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction ordering
    * after barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_ordering_after_barrier_enable = 1;

  /**
    * Determines if the transaction trace file generation is enabled.
    * 
    * - 1'b1 : Enable trace file generation. 
    * - 1'b0 : Disable trace file generation.
    * .
    * 
    * <b>type:</b> Static
    */
   bit enable_tracing = 1'b0;

   /**
    * Determines if transaction reporting is enabled.
    * 
    * - 1'b1 : Enable transaction reporting.
    * - 1'b0 : Disable transaction reporting. 
    * .
    * 
    * <b>type:</b> Static
    */
   bit enable_reporting = 1'b0;

  /**
    * Applicable only when enable_tracing or enable_reporting is set.
    * Determines if transaction data should be included as part of trace file
    * generation/reporting. Takes effect only if the product of 'data width in
    * bytes' and 'max burst length in AXI3 (16)' is less than or equal to 1024.
    * This restriction is imposed to avoid an overlow of characters
    * 
    * - 1'b1 : Enable data in trace file generation. 
    * - 1'b0 : Disable data in trace file generation.
    * .
    * 
    * <b>type:</b> Static
    */
   bit data_trace_enable = 1'b0;
  
  /**
    * Applicable only when enable_tracing or enable_reporting and data_trace_enable is set.
    * Determines if transaction data_beat should be included as part of trace file
    * generation/reporting. Takes effect only if the product of 'data width in
    * bytes' and 'max burst length in AXI3 (16)' is less than or equal to 1024.
    * This restriction is imposed to avoid an overlow of characters
    * 
    * - 1'b1 : Enable data_beat in trace file generation. 
    * - 1'b0 : Disable data_beat in trace file generation.
    * .
    * 
    * <b>type:</b> Static
    */
   bit data_beat_trace_enable = 1'b0;

  /** 
    * @groupname protocol_analyzer
    * Determines if XML generation is enabled.
    * <b>type:</b> Static
    */
  bit enable_xml_gen = 0;

  /**
   * @groupname protocol_analyzer
   * Indicates whether XML generation is included for memcore operations. The resulting
   * file can be loaded in Protocol Analyzer to obtain a graphical presenation of the
   * memcore activity. Set the value to 1 to enable the memcore XML generation.
   * Set the value to 0 to disable the memcore XML generation.
   * 
   * <b>type:</b> Static
   */
  bit enable_memcore_xml_gen = 0;
 
  /**
   * Determines in which format the file should write the transaction data.
   * The enum value svt_xml_writer::XML indicates XML format, 
   * svt_xml_writer::FSDB indicates FSDB format and 
   * svt_xml_writer::BOTH indicates both XML and FSDB formats.
   */
  svt_xml_writer::format_type_enum pa_format_type ;
  
  
  // **********************************************
  // Configuration parameters for STREAM interface
  // **********************************************
  /** @cond PRIVATE */
  /** 
    * Signifies the presense of the TREADY signal in the VIP. 
    * <b>type:</b> Static
    * Not yet supported.
    */
  rand bit tready_enable               = 1;

  /** 
    * Signifies the presense of the TKEEP signal in the VIP. 
    * <b>type:</b> Static
    * Not yet supported.
    */
  rand bit tkeep_enable                = 1;

  /** @endcond */

  /** 
    * Signifies the presense of the TSTRB signal in the VIP. 
    * <b>type:</b> Static
    * Value of tstrb is consider as 0 when tstrb_enable = 0.
    */
  rand bit tstrb_enable                = 1;

  /** 
    * Signifies the presense of the TID signal in the VIP. 
    * <b>type:</b> Static
    * Value of tid is consider as 0 when tid_enable = 0.
    */
  rand bit tid_enable                  = 1;

  /** 
    * Signifies the presense of the TDEST signal in the VIP. 
    * <b>type:</b> Static
    * Value of tdest is consider as 0 when tdest_enable = 0.
    */
  rand bit tdest_enable                = 1;

  /** 
    * Signifies the presense of the TUSER signal in the VIP. 
    * <b>type:</b> Static
    * Value of tuser is consider as 0 when tuser_enable = 0.
    */
  rand bit tuser_enable                = 1;

  /** 
    * Signifies the presense of the TDATA signal in the VIP. 
    * <b>type:</b> Static
    * Value of data is consider as 0 when tdata_enable = 0. If TDATA is not present it is required that TSTRB is not present
    */
  rand bit tdata_enable                = 1;

  /** 
    * Signifies the presense of the TLAST signal in the VIP. 
    * <b>type:</b> Static
    * All transfers are considered as individual packets when tlast_enable = 0.
    */
  rand bit tlast_enable                = 1;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TDATA signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    * <b>type:</b> Static
    */
  rand int tdata_width                 = `SVT_AXI_MAX_TDATA_WIDTH;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TID signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    * <b>type:</b> Static
    */
  rand int tid_width                   = `SVT_AXI_MAX_TID_WIDTH;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TDEST signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM. 
    * <b>type:</b> Static
    */
  rand int tdest_width                 = `SVT_AXI_MAX_TDEST_WIDTH;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TUSER signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM. 
    * <b>type:</b> Static
    */
  rand int tuser_width                 = `SVT_AXI_MAX_TUSER_WIDTH;

  /** @cond PRIVATE */
  /** Setting this parameter to 1, enables the generation of a
    * byte stream type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit byte_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of a
    * continuous aligned type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit continuous_aligned_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of a
    * continuous un-aligned type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit continuous_unaligned_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of a
    * a sparse type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit sparse_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of user defined 
    * streams.
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit user_stream_enable = 1;
  /** @endcond */

  /**
    * Specifies the number of stream transactions that can be interleaved.
    * When set to 1, interleaving is not allowed.
    * MASTER: 
    * Does not interleave transmitted streams beyond this value.
    * SLAVE: 
    * Checks that received streams are not interleaved beyond this value. 
    * An error is issued if streams are interleaved beyond this value.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_WR_INTERLEAVE_DEPTH
    * <b>type:</b> Static
    */ 
  rand int stream_interleave_depth       = `SVT_AXI_MAX_STREAM_INTERLEAVE_DEPTH;

  // **********************************************
  // End of Configuration parameters for STREAM interface
  // **********************************************

  /** 
    * @groupname default_ready
    * Default value of AWREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_awready = 1;

  /** 
    * @groupname default_ready
    * Default value of WREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_wready = 1; 

  /** 
    * @groupname default_ready
    * Default value of ARREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_arready = 1;

   /** 
    * @groupname default_ready
    * Default value of RREADY signal. 
    * <b>type:</b> Dynamic 
    */
  rand bit default_rready = 1;

  /** 
    * @groupname default_ready
    * Default value of BREADY signal. 
    * <b>type:</b> Dynamic 
    */
  rand bit default_bready = 1;

  /**
    * @groupname default_ready
    * Default value of ACREADY signal.
    * Applicable when axi_interface_type is ACE.
    * <b>type:</b> Dynamic 
    */
  rand bit default_acready = 1;

  /**
    * @groupname default_ready
    * Default value of CRREADY signal.
    * Applicable when axi_interface_type is ACE.
    * Applicable only to SLAVE 
    * <b>type:</b> Dynamic 
    */
  rand bit default_crready = 1;  
 
  /**
    * @groupname default_ready
    * Default value of CDREADY signal.
    * Applicable when axi_interface_type is ACE.
    * Applicable only to SLAVE 
    * <b>type:</b> Dynamic 
    */
  rand bit default_cdready = 1;

  /**
    * @groupname default_ready
    * Default value of TREADY signal.
    * Applicable when axi_interface_type is AXI4_STREAM.
    * <b>type:</b> Dynamic 
    */
  rand bit default_tready = 0;

  /** 
    * @groupname default_ready
    * Default value of QVN VxREADY signal. 
    * <b>type:</b> Dynamic
    */
  `ifdef SVT_AXI_QVN_ENABLE
  rand bit default_qvn_ready = 1;
  `endif

  /** 
    * @groupname axi_signal_inactive_wdata_byte_value
    * When the VALID signal of the write data channel is high and wstrb is low, all
    * inactive wdata byte lane will take this value and valid wdata remains in the 
    * active byte lane.
    * <b>type:</b> Dynamic 
    */
  rand wdata_val_enum inactive_wdata_bytes_val = INACTIVE_WDATA_BYTE_UNCHANGED_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the write address channel is low, all other
    * signals (except the READY signal) in that channel will take this value.
    * <b>type:</b> Dynamic 
    */
  rand idle_val_enum write_addr_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the write data channel is low, all other signals 
    * (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic 
    */
  rand idle_val_enum write_data_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the read address channel is low, all other
    * signals (except the READY signal) in that channel will take this value.
    * <b>type:</b> Dynamic 
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand idle_val_enum read_addr_chan_idle_val =INACTIVE_CHAN_PREV_VAL;
`else
  rand idle_val_enum read_addr_chan_idle_val =INACTIVE_CHAN_X_VAL ;
`endif
  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the read data channel is low, all other signals 
    * (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic
    */
  rand idle_val_enum read_data_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the write response channel is low, all other 
    * signals (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic
    */
  rand idle_val_enum write_resp_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * Enables toggling of ready signals when corresponding valid is low
    * The exact manner in which the ready signals are toggled depends on
    * the values set in svt_axi_transaction::idle_addr_ready_delay,
    * svt_axi_transaction::idle_wready_delay, svt_axi_transaction::idle_rready_delay
    * and svt_axi_transaction::idle_bready_delay
    * <b>type:</b> Static 
    */
  rand bit toggle_ready_signals_during_idle_period = 0;
 
  /** @cond PRIVATE */
  /** If this parameter is set, the master checks for any outstanding 
    * transaction with an overlapping address before sending a transaction.
    * If there is any such outstanding transaction, the master will wait
    * for it to complete before sending a transaction.
    * <b>type:</b> Static 
    *
    * This parameter is not yet supported.
    */
  rand bit addr_overlap_check_enable = 0;
  /** @endcond */

  /** 
    * @groupname axi3_4_config
    * The number of addresses pending in the slave that can be 
    * reordered. A slave that processes all transactions in  
    * order has a read ordering depth of one.
    * This parameter’s max value is defined by macro SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH. 
    * The default value of this macro is 8, and is user configurable. 
    * Refer section 3.3.7 of AXI user manual for more info on System Constants.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH (Value defined by macro SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH. Default value is 8.)
    * <b>type:</b> Static 
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand int read_data_reordering_depth = 1;
`else
  rand int read_data_reordering_depth = 16;
`endif

   /** 
    * @groupname axi3_4_config
    * The number of responses pending in the slave that can be 
    * reordered. A slave that processes all transactions in  
    * order has a write resp ordering depth of one.
    * This parameter’s max value is defined by macro SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH. 
    * The default value of this macro is 8, and is user configurable. 
    * Refer section 3.3.7 of AXI user manual for more info on System Constants.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH (Value defined by macro SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH. Default value is 8.)
    * <b>type:</b> Static 
    */
  rand int write_resp_reordering_depth = 1;

  /**
    * @groupname axi3_4_config
    * Specifies the number of beats of read data that must stay 
    * together before it can be interleaved with read data from a
    * different transaction.
    * When set to 0, interleaving is not allowed.
    * When set to 1, there is no restriction on interleaving.
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_READ_DATA_INTERLEAVE_SIZE 
    * <b>type:</b> Static 
    */
  rand int read_data_interleave_size = 0;

  /**
   * @groupname axi3_4_config
   * Specifies how the reordering depth of transactions moves.
   * 
   * Applicable only to the READ data and WRITE resp transactions processed by ACTIVE Slave.
   */
  rand reordering_window_enum reordering_window = MOVING;
      
  /**
   * @groupname axi3_4_config
   * Specifies the reordering algorithm used for reordering the 
   * transactions or responses.
   * 
   * Applicable only to the READ data and WRITE resp transactions processed by ACTIVE Slave.
   */
  rand reordering_algorithm_enum reordering_algorithm = ROUND_ROBIN;
  
  /** 
    * @groupname axi3_4_config
    * This parameter is added to control the reordering priority, in which svt_axi_transaction::reordering_priority 
    * value Vs reordering priority scheme.
    *
    * This member is applicable only when svt_axi_port_configuration::reordering_algorithm
    * is svt_axi_port_configuration::PRIORITIZED.
    *
    * If this bit is set to ‘1’ then transactions with svt_axi_transaction::reordering_priority highest value 
    * for this attribute will get higher priority.
    *
    * If this bit is set to ‘0’ then transactions with svt_axi_transaction::reordering_priority least value 
    * for this attribute will get higher priority.
    *
    * Default value of this bit is set to ‘0’.
    *
    * Applicable for ACTIVE SLAVE only.
    *
    * Configuration type: Static
    */
  rand bit reordering_priority_high_value = 0;

  /** 
    * @groupname axi3_4_config
    * The AXI3 protocol requires that the write response for write 
    * transactions must not be given until the clock cycle 
    * after the acceptance of the last data transfer.
    * In addition, the AXI4 protocol requires that the write response for
    * write transactions must not be given until the clock
    * cycle after address acceptance. Setting this
    * parameter to 1, enforces this second condition in AXI3
    * based systems as well. It is illegal to set this parameter to 0
    * in an AXI4 based system.
    * <b>type:</b> Static 
    */
  rand bit write_resp_wait_for_addr_accept = 1;

  /**
    * @groupname axi3_4_config
    * Applicable only to active slave vip.
    * Waits for address to be received before driving wready.
    * Applicable to a transaction where data arrives before address.  In such a
    * scenario, if this parameter is set, wready is asserted only after the
    * corresponding AWVALID is received.
    * Applicable only when svt_axi_port_configuration::default_wready=0.
    */
  rand bit wready_wait_for_awaddr = 0;

  /**
    * @groupname axi3_4_config
    * Applicable only to active slave vip.
    * Waits for address handshake to be completed before driving wready.
    * Applicable to a transaction where data arrives before address.  In such a
    * scenario, if this parameter is set, wready is asserted only after the
    * corresponding AWVALID-AWREADY handshake is completed.
    * Applicable only when svt_axi_port_configuration::default_wready=0.
    */
  rand bit wready_wait_for_awaddr_handshake = 0;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This parameter is added to enable the structural dependency feature.
    * User has to set this bit to 1'b1 to enable the structural dependency feature.
    */
  
  rand bit axi_slv_channel_buffers_enable  = 0;
 
  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Write address buffer.
    * The default value is set to 16.
    */
  
  rand integer axi_wr_addr_buffer = 16;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Write data buffer.
    * The default value is set to 4096.
    * This default value considers that the AMBA AXI supports maximum burst_length of 256. Since the default value of axi_wr_addr_buffer is 16, a value of 256*16 is reasonable 
   */
  
  rand integer axi_wr_data_buffer = 4096;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Write response buffer.
    * The default value is set to 16.
    */
  
  rand integer axi_wr_resp_buffer = 16;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Read address buffer.
    * The default value is set to 16.
    */
  
  rand integer axi_rd_addr_buffer = 16;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Read response buffer.
    * The default value is set to 4096.
    */
  
  rand integer axi_rd_resp_buffer = 4096;

  /** 
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * Number of FIFO memories to be configured for this port.
    * Each FIFO memory has a specifc address and is given in
    * #fifo_mem_addresses. Needs to be used in conjunction with
    * svt_axi_slave_memory_sequence for UVM/OVM. For VMM, #generator_type must
    * be set to MEMORY_RESPONSE_GEN. If there is a FIXED type burst access
    * to one of these addresses, then data is written/read in the corresponding
    * FIFO. If there is a FIXED type burst access to an address that is not
    * configured in fifo_mem_addresses, a SLVERR response is issued.  If there
    * is a FIFO underrun when a READ is issued, a SLVERR is given as response
    * <b>type:</b> Static 
    */
  int num_fifo_mem = 0;

  /**
    * @groupname axi3_4_config
    * Addresses corresponding to each FIFO
    * The size of this array should be equal to #num_fifo_mem
    * <b>type:</b> Static 
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] fifo_mem_addresses[];
  
  /** @cond PRIVATE */
  /**
    * The AXI slave currently supports two types of memory:
    * 1. A legacy SV based memory. This is the solution by default. For more information refer to the class reference documentation of svt_mem.
    * 2. A C based memory which has more features compared to the SV based memory. For more information refer to the class reference documentation of svt_mem_core. 
    * If the memory type is set to this, the following needs to be done:
    * a. Pass/include (as elaboration options to vcs/mti/nc) “${DESIGNWARE_HOME}/vip/svt/common/latest/C/lib/${platform}/libmemserver.so"
    * b. Set LD_LIBRARY_PATH as $DESIGNWARE_HOME/vip/svt/common/latest/C/lib/$platform (or prescript file if using dw_home build)
    */
  mem_type_enum mem_type = SV_BASED_SVT_MEM;
  /** @endcond */

  /** @cond PRIVATE */
  /** 
    * Enables the internal memory of the slave.
    * Write data is written into the internal memory and read
    * data is driven based on the contents of the memory.
    *
    * <b>type:</b> Static
    *
    * This parameter is not yet supported. The slave supports built-in memory,
    * but this parameter is not currently required to enable the memory.
    */
  bit enable_mem = 1;
  /** @endcond */

  /**
    * Enables address generation based on the values configured
    * in {nonshareable_start_addr,nonshareable_end_addr},
    * {innershareable_start_addr,innershareable_start_addr} and
    * {outershareable_start_addr,outershareable_end_addr} which are set
    * through svt_axi_system_configuration::create_new_domain() and
    * svt_axi_system_configuration::set_addr_for_domain().
    * This establishes a relationship between the addresses (svt_axi_transaction::addr)
    * and domain_types(svt_axi_transaction::domain_type) generated in a transaction.
    */
  bit enable_domain_based_addr_gen = 0;

  /**
    * An array of start addresses corresponding to the nonshareable
    * region of memory. Each member pairs with a corresponding
    * member of nonshareable_end_addr to form an address range applicable
    * to a nonshareable region. 
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] nonshareable_start_addr[];

  /**
    * An array of end addresses corresponding to the nonshareable
    * region of memory. Each member pairs with a corresponding
    * member of nonshareable_start_addr to form an address range applicable
    * to a nonshareable region.
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] nonshareable_end_addr[];

  /**
    * An array of start addresses corresponding to the innershareable
    * region of memory. Each member pairs with a corresponding
    * member of innershareable_end_addr to form an address range applicable
    * to a innershareable region. 
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] innershareable_start_addr[];

  /**
    * An array of end addresses corresponding to the innershareable
    * region of memory. Each member pairs with a corresponding
    * member of innershareable_start_addr to form an address range applicable
    * to a innershareable region.
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] innershareable_end_addr[];

  /**
    * An array of start addresses corresponding to the outershareable
    * region of memory. Each member pairs with a corresponding
    * member of outershareable_end_addr to form an address range applicable
    * to a outershareable region. 
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] outershareable_start_addr[];

  /**
    * An array of end addresses corresponding to the outershareable
    * region of memory. Each member pairs with a corresponding
    * member of outershareable_start_addr to form an address range applicable
    * to a outershareable region.
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] outershareable_end_addr[];

  /** Applicable only when axi_interface_type is set to AXI_ACE.  Indicates if
   * the cache must be updated with the protection type (as indicated by
   * svt_axi_transaction::prot_type) of the transaction that makes an entry in
   * the cache. If the VIP auto-generates a transaction for evicting an entry
   * from cache or for cleaning a cacheline before sending a cache maintenance
   * transaction, the protection type properties recorded in the cache are set
   * for the auto-generated transaction
    */
  bit update_cache_for_prot_type = 0;

  /** Applicable only when axi_interface_type is set to AXI_ACE.  Indicates if
   * the cache must be updated with the memory attributes(as indicated by
   * svt_axi_transaction::cache_type) of the transaction that makes an entry in
   * the cache. If the VIP auto-generates a transaction for evicting an entry
   * from cache or for cleaning a cacheline before sending a cache maintenance
   * transaction, the memory attributes recorded in the cache are set for the
   * auto-generated transaction
    */
  bit update_cache_for_memory_attributes = 0;

  /**
    * Applicable only when axi_interface_type is set to AXI_ACE. Indicates if
    * the cache must be updated for WRITENOSNOOP and READNOSNOOP transactions.
    * Currently supported only if  cache_line_state_change_type is set to
    * RECOMMENDED_CACHE_LINE_STATE_CHANGE. Cache is updated only if
    * transactions are a full cacheline access. Transactions with sparse write
    * strobes are also allowed. If transactions with partial or multiple
    * cacheline accesses are received by the master driver, existing entries in
    * the cache for the corresponding address(s) will be deleted. If this bit
    * is set and svt_axi_transaction::force_xact_to_cache_line_size is set, a
    * constraint in the master transaction forces all WRITENOSNOOP and
    * READNOSNOOP to be of a full cacheline access and FIXED types bursts are
    * not allowed. The specification allows a cacheline to move from the
    * invalid state to a valid state only for a full cacheline access.
    * Therefore any backdoor access to the cache to write into non-shareable
    * region must write into all bytes of the cacheline. For a WRITENOSNOOP
    * transaction, if the cacheline is dirty and a transaction with partial
    * write strobes is received, the VIP merges dirty data from the cache and
    * the data in the transaction and transmits it. If the cacheline is clean,
    * no merging of data is performed. If the cacheline does not exist,
    * allocations are not made for a WRITENOSNOOP transaction based on section
    * C4.8.1 and Table C4-20 of the specification, since there are no cacheline
    * state transitions from an invalid state to a valid state. Hence, a
    * WRITENOSNOOP will modify cache contents only if the cache is already
    * allocated either through a READNOSNOOP or through backdoor access of
    * cache. For a READNOSNOOP transaction, if there is no entry in the cache,
    * a new cacheline is allocated only if
    * svt_axi_transaction::allocate_in_cache is set. If there is already an
    * entry in the cache, the status of the cache is updated, but the data is
    * not because this indicates a speculative read and the data in cache may
    * be the latest copy.  Cacheline state transitions for READNOSNOOP
    * transactions correspond to section C4.5.1 of the specification. 
    */
  bit update_cache_for_non_coherent_xacts = 0;

  /**
    * Applicable only when axi_interface_type is set to AXI_ACE. Indicates if
    * data must always be supplied for READONCE, READCLEAN, READSHARED,
    * READNOTSHAREDDIRTY and READUNIQUE snoop transactions on the snoop data
    * channel if the cacheline is in a valid state. If this value is set to 0, data may or may not be transferred based on randomization
    */
  bit transfer_snoop_data_always_if_valid_cacheline = 1;

    /** 
    * @groupname axi3_4_config
    * If this bit is set to ‘1’ then transactions are only eligible for "write_resp_chan_lock" only after 
    * both address phase and data phase are completed.
    *
    * If this bit is set to ‘0’ then transactions  are eligible for “write_resp_chan_lock” after
    * Address phase is completed.In here "data phase" is not considered. 
    * 
    * Default value is ‘0’.
    * This attribute is applicable only to the READ data and WRITE resp transactions processed by ACTIVE Slave.
    *
    * ** Note, Eligible transaction are given the “write_resp_chan_lock” according to the “reordering algorithm”.
    */
  bit write_resp_wait_for_data_accept = 0;

  /** @cond PRIVATE */
`ifdef SVT_VMM_TECHNOLOGY
  /**
    * @groupname axi_performance_analysis 
    * The interval based on which performance parameters are monitored and
    * reported. The simulation time is divided into time intervals spcified by this
    * parameter and performance parameters are monitored and reported based on
    * these. Typically, this interval affects measurement of performance
    * parameters that require aggregation of values across several transactions
    * such as the average latency for a transaction to complete. The unit for
    * this parameter is the same as the simulation time unit.
    * When set to 0, the total simulation time is not divided into time intervals.
    * For example, consider that this parameter is set to 1000 and that the
    * simulation time unit is 1ns. Then, all performance metrics that require
    * aggregation will be measured separately for each 1000 ns. Also min and max
    * performance parameters will be reported separately for each time interval.
    * If this parameter is changed dynamically, the new value will take effect
    * only after the current time interval elapses.
    * <br>
    * <b>type:</b> Dynamic
    */
`else
  /**
    * @groupname axi_performance_analysis 
    * The interval based on which performance parameters are monitored and
    * reported. The simulation time is divided into time intervals specified by this
    * parameter and performance parameters are monitored and reported based on
    * these. Typically, this interval affects measurement of performance
    * parameters that require aggregation of values across several transactions
    * such as the average latency for a transaction to complete. The unit for
    * this parameter is the same as the simulation time unit.
    * When set to 0, the total simulation time is not divided into time intervals.
    * For example, consider that this parameter is set to 1000 and that the
    * simulation time unit is 1ns. Then, all performance metrics that require
    * aggregation will be measured separately for each 1000 ns. Also, min and max
    * performance parameters will be reported separately for each time interval.
    * If this parameter is changed dynamically, the new value will take effect
    * only after the current time interval elapses.
    * <br>
    * When set to -1, svt_axi_port_perf_status::start_performance_monitoring() and
    * svt_axi_port_perf_status::stop_performance_monitoring() needs to be used to
    * indicate the start and stop events for the performance monitoring. If the
    * start and stop events are not indicated, the performance monitoring will not 
    * be enabled. If the stop event is not indicated after issuing a start event,
    * the port monitor stops the performance monitoring in the extract phase.
    * Note that any constraint checks will be performed only during the monitoring period.
    * <b>type:</b> Dynamic
    */
`endif  
  real perf_recording_interval = 0;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed duration for a write
    * transaction to complete. The duration is measured as the time when the
    * the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    */
  real perf_max_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum duration for a write transaction to
    * complete. The duration is measured as the time when the the transaction
    * is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum expected average duration for a write
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is more than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_max_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected average duration for a write
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is less than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_min_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed duration for a read
    * transaction to complete. The duration is measured as the time when the the
    * transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum duration for a read transaction to
    * complete. The duration is measured as the time when the the transaction is
    * started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum expected average duration for a read
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is more than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_max_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected average duration for a read
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is less than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_min_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed throughput for read
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_read_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected throughput for read
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_read_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed throughput for write
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_write_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected throughput for write
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_write_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed bandwidth for read
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_read_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected bandwidth for read
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_read_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed bandwidth for write
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_write_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected bandwidth for write
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_write_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis
    * Indicates if periods of transaction inactivity (ie, periods when no
    * transaction is active) must be excluded from the calculation of
    * throughput.  The throughput is measured as (number of bytes transferred
    * in an interval)/(duration of interval). If this bit is set, inactive
    * periods will be deducted from the duration of the interval
    */
  bit perf_exclude_inactive_periods_for_throughput = 0;
  
  /**
    * @groupname axi_performance_analysis
    * Indicates how the transaction inactivity (ie, periods when no
    * transaction is active) must be estimated for the calculation of
    * throughput.  
    * Applicable only when svt_axi_port_configuration::
    * perf_exclude_inactive_periods_for_throughput is set to 1. 
    * EXCLUDE_ALL: Excludes all the inactivity. This is the default value. 
    * EXCLUDE_BEGIN_END: Excludes the inactivity only from time 0 to start of first 
    * transaction, and from end of last transaction to end of simulation. 
    */
  perf_inactivity_algorithm_type_enum perf_inactivity_algorithm_type = EXCLUDE_ALL;
  /** @endcond */

`ifdef SVT_ACE5_ENABLE
   /**
     * @groupname ace5_config
     *  It can be set to either of three values below:
     *  mte_support_type =svt_axi_port_configuration:STANDARD.
     *  When set to the above value memory tagging is supported on the interface, all tag operation types are supported
     *	mte_support_type = svt_axi_port_configuration:BASIC.
     *  When set to the above value memory tagging is supported on the interface at a basic level, a limited range of tag operations are supported. 
     *	mte_support_type = svt_axi_port_configuration:FALSE.
     *  When set to NOT_SUPPORTED , memory tagging is not supported on the interface
     *  Only applicable when SVT_ACE5_ENABLE macro is defined and svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
     */
  mte_support_type_enum mte_support_type = NOT_SUPPORTED;

 /**
   * @groupname ace5_config
   * Bcomp signal
   * Only applicable when SVT_ACE5_ENABLE macro is defined and svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
   */
  bit bcomp_signal_enable; 
`endif

`ifdef SVT_ACE5_ENABLE
 /**
    * @groupname ace5_config
    * Enables unique id identifier feature for write and read address and response channels
    * <b>type:</b> Static
    * Only applicable when SVT_ACE5_ENABLE macro is defined and 
    * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0 or higher
    *
    * This functionality is not supported yet.
    */
   bit unique_id_enable  = 0; 

 /**
   * @groupname ace5_config
   * Enables Read Data Chunking feature support in master and slave. 
   * <b>type:</b> Static
   * Only applicable when SVT_ACE5_ENABLE macro is defined. 
   * Not yet implemented.
   */
  bit rdata_chunking_enable = 0;

   /** 
    * @groupname ace5_config 
    * It is used to set width of the rchunknum signal. Applicable when
    * <b>type:</b> Static
    * Not yet implemented.
    */
  rand int rchunknum_width                   = `SVT_AXI_MAX_CHUNK_NUM_WIDTH;

  /** 
    * @groupname ace5_config 
    * It is used to set width of the rchunkstrb signal. Applicable when
    * <b>type:</b> Static
    * Not yet implemented.
    */
  rand int rchunkstrb_width                   = `SVT_AXI_MAX_CHUNK_STROBE_WIDTH;
`endif

  //----------------------------------------------------------------------------
  /**
   *   post_randomize does the following
   *   1) Aligns the address to no of Bytes for Exclusive Accesses
   */
  extern function void post_randomize ();

  /*   pre_randomize does the following
   *   1) Calculates number of tagged address attributes set to '1'
   */
  extern function void pre_randomize ();

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Vj5GCxQaanPTR4pdHIaHVb1D35mZ9+SU6srKFKwE4bQ3xMyyxaRN60y4Aq2ad1Su
lsLs8U/cz3fCXPPBSqacbsDtb3d0y5lDvMSNx+egWI2BdWHeCJ8703CS7AWne3pT
szs1XIR6Q3n7lNDjWgZtYDBYoXNOOkb3KQUOsvtWj9A=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1368      )
3rT4zYMcmTWvs87TGecF4AF7/6dB1agJM1dQHxFyVLWqiY6njTbq7ZPGkmQMQYIO
aCKwvx2HiYHAHV+TKa4OnGWIRNlToemlD3MwZijFj2dJUzk346gfxjOpNITxmGJa
pDlIyltFwQuODE7TnQESXtQwhqe1cPx9w50vRl0FCdeyKOa/8pWy4zFJuhVvdwxo
45jvFJASQnNOB2sNSeNLsNNTHRT4QNtN4NOv8DGHXvRhNLxDluyTO+Agm1UuLVD9
JJnNTQtJBfYiYS6QuhO3QCzhE2CCraq56v4aXMhvqoBUCWR3+6KwnguOFPndG4EC
tny5Ayr0sV4/RmQ7/jnWu4T1faLPmmdR0GZyJEnchpk+mAGezL4kT60DGJt+UBBE
s+Q88e7LsVjNPODiagFKmnuUR8kXeT2/UYy9GLc4KK2Qf+Rnt4p4ftd9xKj8+BML
uJn5UQvLs667yaM4x1SwHGqNYJsh+1lsoFTb8xHYK9M=
`pragma protect end_protected

`ifdef SVT_ACE5_ENABLE
/** 
 * Returns 1 if bcomp response is applicable on this port else returns 0
 */
 extern function bit is_bcomp_response_valid();   
`endif

`ifdef SVT_VMM_TECHNOLOGY
/** @cond PRIVATE */
  /** 
    * @groupname axi_generic_config
    * The source for the stimulus that is connected to the transactor.
    * This member is not used.
    * Configuration type: Static
    */
  generator_type_enum snoop_generator_type = SCENARIO_GEN;
/** @endcond */
`endif

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
FIxNcfXZes0Gu/UQdrB2U7S5CXywLpLwpUJx5XX17T/Rr0j9TEXGhrOL66k5mce2
pa0MCMvR8liL83+7O/ZBpjFRuemZlnTkxyz+RmLABizbaFM0uMyonVVjBD2rqn/h
26NeseKt+w03aJaxWXqTMRFuXoAjVC+YaixmrHOL/Jw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 14642     )
UZguXGwBbT0+RoI44/gh6qnRWTU53IlM1Kj2EGNK2txwED5RXi+n4XykQrkZCVcE
hWk+3W9+ZPPdoaRxfxNP/e3TjXxTnv66WYa0mj8h68+g5DSZlxGbl5hlmwOMk1SC
SnmmtLJbx0Tth9OkMcCipnL0GJLcgGmy/O7GomMMTiyAksXqDc7W9S6pQPEx0rbh
qDxlTXb9YWYk9bhqiqAp7ygM3i9ge+sUiIurI6kFTOczpkriyAnUWc38kazOnE4c
iCF34j/ByxlTPkK/Lg7hUNPOGqbxh6k2I95V+uie0931IrdVsDTy0+McFL/cjpl3
kmFhM6DASDMmBWleZt2iSqq5q0KiV7J/TXMA3LcRCHfiY5CuUFldmTPGVlhC/n1x
KpweY20Q+Je1UcYSd9QjyUo55kbd+otq6IscQO0jiYs9JDohyZ/JGt6TerjDGfWB
An6QfUHwRZoq4nJQMfMY07v0vLHehAGBtGTZLraIYlrtuhjnN1uQ9hDqZbo79Cqa
fY1x7Vzv8/zvGxC2dpCMLPat8vUsNXFdqnn9pFvzilcwYdFqDxYOXEvMCUTCvtf9
goVjkgyckag3D/1LKzNJwjxZ+fik/Bd9lycC8T8i0rfiAdWgd7fMRU5NArEQGUFT
WpXfCttohz3unuKWWabVgWxHXieeMn3/Es59aaLx/Vn8HA7iAISmNigpjwwa5+Ze
hKRSNCIHu4p0g6obJ7E6RuqPYAIbP5/7WrKpG5iKPl8nWlR8Lci+C5jTjFwU/mHl
0hp5Cfu9drxIqosSxs0y1CLaHH74N9c8oj3vkEdG5TFGfW/kXNJoOjWLGa/nw1hg
WFVcPLPAZqihQwP1n/XOjqv9AsAa1iybJGBxG3x+VOkVuVnuOjMXhMkQjBfhOhvk
SFVvQuwgX9ADz1IoKKVmmCLXymP7tuBHFRfMpasXNQu9Mv8sUfEiYCBOfDMRVXMf
aLQKR0duG0Usu6a05DTyuW5d1yxV+UnsDC6Kz7mgXxoseK6yE2fA+Q5mSW7IrN40
dB4DRdtJKvIQLDRedOMeGKnnMoa6kvWak7im47EYhvbOZHR8p7LA094q53hxVxu7
F4YBJ+5dAFJEM/TaqvkdqpflmCYB5KSLvgSN7Av+Rs6ORkU+4YY0QUuDHh4Pn2Pz
zzZ94vH5yHGThM1iI1uGW3Yta7olDKfGGuf5uOmRQuJKRLThJ2G6WoRNN4f5+Frp
r0bRNejLsduWLQVve+R26f1vKBhNMcM29gwAthTdzv7V8K1Y7KTZ99T5gGIWGQxY
y1nl+zpchPO74qX8vRRAFTIMivrgAj/kjpCGZ/POXLd02nrnSAfERnjLNe4cPv1S
ZOCP9N5snKOBb0JMNozgUOPN6bnlTRFM3q1LAj+5FGf1jpjCjeV2pmq2kVr/3vHR
T9yvSlWSUsDfQsWETQL8yWK6I6TmduGsWQ50sgAmjEvnv4rAKITp56YVg8YlG9nH
yvpnNFweEvXKismeKihiAGhisjmhNNP1YbgBTIONeBeUpL69H5oE5mirjRtEV47l
nqiEQ4sAHxh6UzsxxUm6zD1SebiGqM8+MvVSlgCv+/Apx0vE+FRmvkfYv8kH379m
u1obNBL0GUIdD0sN/XVgXGc1HRzOz6LBHri7T6VZ7LAqbZEFlSwomXIduPTuCjPn
Px0vigF0lG7PC63SxoDJfqy5tklYBXQqJTqazxSRCzU4OKbivCEnLu4bKk4k6c8e
5rcA55DlZ7pe29WQHsGt4ud8vPBwlB6viKmOn5ZsydSXfvaB9JDrxRgjl7C7qHh7
ksWxMf/P8KCTLcAA4xE1cqsvfRDNyXSxDvfQXC9A6Aqu3roE7ZSk2V3wVttM3mjV
chzkcU8Ji0iVDSmTN9LViD9KMgdc4xOoUOyjxieO+EKFgaGyU6Q5UzmaQFsTuXC2
oZxsxc6FKslQZeQ42C4sHP7+l5L31JR8f81R6vRXlgkJ6LBp1ZMPcO2me5Al6Hat
FfXTq64mtICzg+8Ulc9rfwlhwzYzZR4XNYL3bLkglnjnUTmjiLTyscMabJmc+jkR
a5o8zNNZlGW+N3tHnfahA9LiysdF6nQTLwZyWJtbuN+1LM/jjK5IItaLPsMt4Bjr
7YW3bixpsSZdP/B9WozkuK6NyCCT01a1GRo6Qd/sL5UJg0A6Y7C2d9l3Of+HZOhx
14abVNaMd3/tI+FF6CE3Ye7buJ22YWgyhm84gGA5rYlSWUjysQrhnN/s+eb2nrnx
4ifqm4tUzaoA5dHP7N3iwIFYn1cA6DmF1YE7+0/h+N5gBc3VHMXOAyz3qA5mFuiC
k/ViKS3KCWiJ0D5e4jcmg4Hr7Dzn6/YRRyuus8QKEY/RkYmC2Cdt0q808JkyzwKS
VLhq4XcDwi6bygezXnM4SfHeFh0xZFAkl1E8lyrVfA29Bng2g1feHKbjODAn/4rQ
FDX36lYZDGfhCw4WeB6H8FJwjRHQZTbkldaIwcmQ456W92R77trgN/bHrxJdUb7I
b98/7SLWHwBS928l4ooLwO6P1quKHDLYyecIOjy87GlZNUxL3eOVL2CMwIKK+gSU
lkurm0T6K/6N7XaxlhxTBY5WcjYvR3ovxedldTfcjQveDz5IzU0uZDcoK/vgyF/W
hDrfqUXGzinUbe6yVVDf+yHCdE7IA1+nBHegMUUS5mR5gEc5knIDIVcRAGO0DzVp
Yqr+lRq6Yc0d2luHOIqM79tWYV0bU2nxrg0oG9d1qBI+rlzvWmb0jHYpacftL3F4
9UyFSi/QjKlpMw7YJmCllPUcH3jpUzqB8mQzm1mIuhE/0yhKcrbTOH7kreiasMlq
aDguLHuAOtVQJSFB+058P35/bsReIdHs57VwbRWdG6qwmB+2GjwolhbJzccuOADh
/y1Zw06vyXUCwtaTjJizcsjnUk0Dcgs6Ci3idOs2HIOwLOZTooI5FAwLoCFYpwHb
cGaAcUdS2tQKphBcoSAqepz4JYrE8N/3iWSDWzvbIXDF6MY3oPRT74ph2QhZV9Oc
Yn1TXG7B44m/m7M9E1nIEgCvfaR3nr931XrN1fK0Swr+bJOCdBPYTxQibZXIlUdN
wm880XdVomCs1cYEuBoT9QNM3dzxjvOuAHA6NjpfhyLiUxpo5EHNZAAQaLRB+HkN
r7S6PHY22wZHOYtXZcfVEKiE6kqvpy8op45EsNN2hyffU2bO4pkex0s9wjrEeeQS
4jkpsbtwXjbQA/RqH4537NnXOv4SSQsiEy9H5EUAstChP4sLrzmsSse8gmYHwr9x
ueQ1zFiUkEG+ZZfm4DlWllZvFxPNouEqkN4PTwlI2UQp3rwSEOCJkBcdYawMRQT0
rF5PVzVpxswlcX0MMMo7KV9ABiqJiARXHvDrn3Ah2D1HakIaKXiOPiqFXYwN0S20
agw63vnP17BfXJ3Vs86zrNgETcZbmBLWy0OpCmS7AZbBlJbyG7rXFEurpGuT4Ij7
wirPbcDJb7AkfC+ajVGr2yr6J2N64Wco83r+v17QbFakj4Vi6J7p3oNZezeb6Omf
e9kj8QA7hkCe6kXSa6/GDkKLM/6JYsd77nBa+LzR/Trse3UfvYw3pxeBkmi7HXuX
RBQAZyUv9wx9zUqgFB7nlzFVYiuXWI0cO2f8daRP3L9TRRFl1BzNIxL6xqr3Z81p
SuFw6ZmAjizDHCtb2POu6lLJJqF+TZlKw7ZZXbtYhOHM86MhO3YbghG+Mfb6MZmR
42LlFea3sJ2MHUNmC76PiFt+JHoAFtUwivc6KIvmK1gdnSIj9jxZswEOX7af1jxi
Na9zgFkAs4IMyn8k1IntEK7hcH7yhBi810LgTy/D4f6TzqsX/FlhrKKLcv+avtn+
smf0NG9CohQle2Zpc/UL5IhM4gRkjL2GrNb6hS5fd5M4g+PaqTE6lcJOMLphICuC
JKIZJX59OYsczdP3loHdUXbqo3gmJwXbHv+H4dLW4/ItRxAhqSm13wO6aF1V4+aV
vFlWn69/1ZQvxN0mVW8FhcApI57UWCwNFb6zrdmFKHO8FryIGmGfinsokd9eobMA
DeIn8o5iXUcCv09n9aoNxg7eeco1wge4x1x5vu7Wyqv5M4UAzSldCVgUGlI6NDXE
2fTkiFSOCpHMNDq0cuGAdfNtQrL2FQrTyRzbhGbNjm8ZC3piZ1cVZHIxkefRpv1T
m4lhZSWBhq8awQmVX2Gott30GnKy4lyEyosGiesbRvasfz1eID0B8nkKL3E4cf6b
yDIx3WQGMEXdkRuna+wt/Kux9kkdBiW9qAI4aGOWBRTWnlfCDXyCjZDzUM54rTk8
BSYUo3BgfLxKOHo5Kx2OqXjOLEbKBqnG9UE9cZjqMcfhn5ZELFaKHFQLoW4k6vf7
FlEjlKuZAtBi00+eHa3Uu9F5THd3s2uUyMwgUJpW7SCaiKq7K0YVGeYHzGyt6zW3
rXRNK/s5sZaJGbvWnpjy5DnfUxt7c/SdPz2rtdKx/4EgQ+5BRNuWQTc4uKublSLp
tBGcPi1bwxE50Zk+T9/sp8dVmGPMjQXBDGbk0UHOfWEcRkP1nM5LmZQMNBlM6ZdS
7bQwpYpjXnisUMQ6JxocRtyE/Vfj6ODGSyAKTsO62Dq7OFBXT/rUY08jfWMNgVTw
heTLRj9/n/AhDysRc3FrBk99HBy/w/VALWiqvDJTELYhDXTnPS04mr+IKNNBOIUG
ohB1JCAds6MeKEbBDQSmeAR04Hw1/2xkgq2M/U+6jXTx2BT8QqkDG/8C4j4Qbx4V
icRPn/2RekZYiAlKLkk0MVTwDDdVc+10ew0qM69ISWbSZGtS7+t2I6eEU1wbfJvN
+AuevowfZ1siKrGNvuC8mbw5p0xVbCdyudvGKzFCr36+7fTls0QSpB/4NyzhyBFO
zRVLULYZqo5JBtH5l8M3LARVQmYKGz43Z+R4IAAjEBrgc6FKIcCSu88S5VYzDX/J
5Hl4qD9iMNz6it4ZEGDILfSIfbWxQz+1UAh90+ApnsRmjj97/BjryWeorJx+JVTq
8GmY2Coinep0AmL3/j1oSLGytRyS2aEBJXhQG0JAbmBPRXpH0JoCilhYi0x7baat
pItI/XVc+SrFH2kiBBBora3qPWCv5JC+08WY40fttEb48sR1OXkTkvVl8HT+ZKpd
jsyiFQRHVfTMv7DimLxK8QbjuMyK2fOZ1mQYP4dQgkj+a/4r7415BEoGLYicrNUt
UxzGKvm/lfJVn6MIuxfjD7uSHjYHcCfqNoTWowHAJ9v0fN0nuFxSWfA4EQwW+cCw
j61ombhsecdXiU5q2th3aSSfw9CEPA8jPvY8syOqtMNlxJanarJpTo3jgUeQmI4H
PrPDkklvYFs8fp/xhhuw8dz+OplYktJIdWuRquUTxFYuFnog6EkHIo0fq62NcT0H
l5nGYgMk+HlB6QS3i6oelwI5fHjEK7QGKRd/fybDbe4kVDdfwOYnA+c81NAnzzEn
HJRcvmLDOBBdJP6Chz4/aFCk8rr0Rhi/QGPagMG0L1bOd6tDeg4ugoaHQlS4uc7S
yhCMhrkVrc5rF4ME/LmVdIbmWBk12vaFcBEGxzJ3KYPp9vn1YTwCvEhWc551GM3Y
5S/b5PJRVRNGBtrUqNt74849t77WA1oKJRvqUdydNycq2TSYftnhPZHx9UdmfJLh
tl94kVzOEhtMqMT5DyEFNhgQBWCbZzrH+lSD5pYJiwX0seH2ycAmpGkULeYkr1ZD
g3fQ2yZL3gyLkPX+957VZ3/L+PL/XPEawxNwSqFAGxuEwoEoreiJHv8ynp0ck031
uSTZL83hGvXkgE/Ut0iXD+VIYpPvJ9+tzWmB/tFNQakkxQTSA/Hss+XiAw7qkM4p
qem5nEuTliqawFq15X+aSN1B30SI+nWJESolQ8Zq9kGuoddlCGjjxWAp00LM2Xj9
xrKVCYm/qKrCF0Sgy6KjRW6Ap3ItX4Nck4zRZDmFKDYXgjk6kosf2XR/Eyra8pOW
BTwimh9ZHK+Ee4fWpdkSvopt88rQojrODYShjQvNecVaqL0fb3FaSDBWvbIicUbW
f05VvwZ6LPCwFgJ9U2Bd/7Gd4o0JJS9EbBLj65Tfcen1q+OKYixec3vLg9cqf0tH
03jPva+nD80Q5YRRNSv4wDntdlDZ0g8Qxf8lL0PiACOIaVtJ5/BclVWyF7oj6xlF
Sbti9TArEjNB/eKUXr+w7dbhYTuz8PHdmqLKJenT9i39jHEi9sI3Q0zdSbt5bM5o
nYYUP9cY1dBevRiUMSjUwlG/24xK1UO+GGmku7PHqcPWvG6cRvVLGOnnWjWWTuqw
vL5JLvLcw5votv2kJ19DRuZAeypcj++Ka7R4cQrSllo8pF/qLv1NyG471CoMS4/H
CYeXuJTPAl4gPaReWcgwVY15ISm9q0LGUzL0GgYBqCQGjKEodVhm3nFGYCF74x3k
2LowalrG2o22NmiFBV9DShYpjwydE1dAmqdOAp+YrJXeU0WVrBrfW9keWliJcuKG
M6MxQXurnki1/znHSYqXnjXe0e449F2UDflmewbuxsqlDcW5VC62JCaLpmErm4Xx
ax/QrlfzJvTipUrPPXiDa5qnEa+AnQ3fXRUleCPSD0NFLoSLNekjB4B2y50PGPWh
8pxfezGhjumAtmEPzF23iI5L/HgirNJy2UFJk9/9F4tdPD3hH4Vnorwc5h+DXa+Y
oUdW26w0hF/ljFCI0VQv5bZd6G2tHvBp3E7XVJkIEc7qVSTlrCK0vtpb6h3LBLdc
lW3sw+4yEBGdQCZ2SBCtS+jf/wK6NaY2mdonyPuQQIrNVRBop0hfYruLe0GEy8NK
aCFdncrcu8ssfbZWQt1NbBCbGzHYO6dJ0faxp6acUG3OVsPl/WyWhLJFJrdNlkPM
fy6DFV5OJ/7ylYCTofd/y7F/vfHJ8O+wbxl0cYqRhMNGLdNj5sbwGf2WTOscU+RI
h5p/aPO8H6vBn4QZ/hAsp38vEvXt9paa7p1nNrYt8RpYU9QQRCq1Q2TAtTd+/XCr
iXR0+9ZKYNbsJSWu73/V2+/MELtO6prGWx8F1o7DQgde3y+SpRXwlDTS4VbcINIp
9HBWBmdPaoLuU6elV3CvnFD+HL/qCIZTl7Dv111yR/SM1x7dAx4fxUGJMBvmqrF1
itZvMP7vLbQV9Ofk7EoMLb1DwEhrOFgtqeqKD8P8/OOzmIK/X2HwxPK1hobtPnUs
Xaf+be7HeQ+qyU7xwcOaAFI6qTBXiANvXRxNx1ZdjCsLsCECbyxR5gT61rdicQQx
CInN0CDxKx+Yu4Fil18xkc4X4VylXFoNlJ3jjJtueeZls5d7wIrIK7Fz2PfPQ+P8
HUjbpMauDNJ8qd2FYY0z9F71awRRxaHWCAX8O0CcKzkYTHSz+5XWz+opSwBdjrZ3
Qo5AjDKh3kCJG2t8ZgULWJKi/UI9ebHFdQtosxAjmVypi489mBBX8E9Pnlc1uKDX
7Ox52ihMD9u1zo0IugzbXh6M06KmJUTo5K7Ez34rxSb1G4Ei1gZDIC9p0YkWyYg1
e1moL9+Wt4d4+pfG8TwfAo0efs3lzM7kf3tLq6yVWSn+fRPa6gUp4I6lNKCz/ed8
70v3Ule82hDIqW3namHhwbQOpCTV3/fh4ljojYbIRp9t7bX6zUxMHkbZ5GBMgiq8
37dpJh2K+0PkedA/yYwCrXEq+YTJL7xzfJy7s2nJAYJv33/yW8do82gquQAaTbpm
PKpdtiiGjhKeNaYnA8OT3MSoCvVRzWw0oZnSSBLWe5jbuGK0x9A+RzG0T9mjSkWW
V7DxsEePbOxkvExR4FCuYyeAK7NLtxlpvjtJmRnFDKRXyetN89EGJTKtqW8NvDdY
VWDvcXAHSYSCqJ4+97kLwMBGnOlSO6/IVBqSRCCquO+wSY7vUQU+rnPNfgm3V3sb
6O2dgmhi25PcsZWSTEYjS3Mwtljsr3FDDMY3Q0n+zz/HFdd5NmbF9CQn3YaQMVhR
37/fziPvVEFOzlbnEgu+UKkiIGojjYXbSBfdljb70hKD5Vdds1SfUyRG6Av4/YZR
IzM6MZpZsIOebBHMatEJLqex1e02aVeR2JYZe9OhsqduttGl4mhV8jUuV8P37CVN
J9Fqz3YSgJXFzZsNAo+efRm0f6LJwDwFbptFrtHHJnqnd3zev1Orvgpr8MTfcQY3
OtPE56t2bqwti7JZ+6DvwF0isvGEJ+JVstb5V89iA1eCa0+/qkx4ocP02TqgGTZC
mSpPD3cmGMuCw4wa8qoYxK7Tz1oFLkQiqMZa+cL/UiNp61Im/ZojeQdm7ZRBYhTG
ruLgB6Wh9kK/nDGwwbOJj89ktL/1G9i4hR4lWNOq6UPMXNySqDVGQEh117QZeego
3P0NZxD5q+TDIbHB+QOOvyAgDURk2uRN2HwiNXU4txQ0OunssE5EF6EPEh+1WLlI
ouEhMvsLca92Wh2x7t4HgzMAO9kb2C1xf7gal/bKMgdsvEv75NRGHlj7A+BcmWom
9nNho8QQ53l0oH85541sZ15CC5twF3KIiUCnvARiQFtXnJVzX1ygY9wa9rkHG+gd
uHAa68MeRAe52h1MCqquR/eQvPhduOfvfjEkIc1ivfsQdt2ST/rB1Qr6zTDSxBv6
JbvaNjY+WQfvqf+gvASvPmsIO7oRoIyOzKatPXOoT3edTaxg69+d3jUV+Uwy+mmy
hRjIdCWpCcZ0mjj7/Axq4GclMA3D3F2SRLRp2HoVPQn5Lq/m5pr+BIcrSkbYnuD/
FAebAok6FtGFkj/2zX98oB5HocveuGNjmJOQgpM6I0SEKtxGCfZMvQRyNEs6BmXh
xqQQ50/qKkMhwBc/QN7D5Es8Hvhqs6eEYwYFv9EH2R7DzkRO0UQuN/wOK+MphglO
IeQL4ms1s279s32zHBkK6KsY86YBE67XQo4kLC01/zu6IoXApCRdQR+fUkZkjBYd
A/eYHpJB6lh0wpPEgLrYdo2HFrD9RVRMLN0mfFMLC2c5MEHSZ/VwkpA4GCPv7zl7
MB0J/ONDrpKakK8llnhC1HZVs5rApWhKPF1vP9lveJDWZIajIaHO5HuEN2woQRp3
anD7102UV76qvVIXPvoFwCiPRh1xMUaAKRQ+AnAZJmSuy4DPO7OvnhZ1rFMltC4m
/wzFkG7DPsPCVkgmfL7QcXooWUJ/dAEZdlWRXOyyCY4FyOPsT+ak+ymwrT7Hsvvf
A0v6ziCYC5JWHiuwEYzF0HJbfbIxRmtSIJ9VqPRvHfKvGbCqPON0B4hwlhnIlPQ9
VLSyvG0M0dbPTnRE4KCL5NRcbRmugS0ECQK+SOGxp4X2NM4dzj1UFMz/AXGUobjh
RHqpzTi2GSMOqvLdFQ/G8r1Occhfo00G/VBzOWvZfhW8aRRVUfa2j0gmNenFrcrF
5nx1Dh1mOrVH9TQoo8VjcOD4NZFacH4bQ68SyB0oodL8Kqt/l75m2KOvgUhWS9Ta
C+fs2mvm3KbMozLhN/kK6I6LYzlUa2WKWvGfCSP96h/gTxw65YDn/eEAK5a80fiA
LbF5I+2hot0CmwINfViaLSA6mGp1K9I+z1dPJmouev46aSUMV8MmDFP6lpFyW8j2
9dd7s2G60R06RtyzNX8VR9Cr8wUtNFw8WfiN6IXiDlQZTZtWX30QNwyFg0WTEenl
IieqamNDDS2NUOGdXUBwnXgRKT1chu+4UvERAAm790rbHd2D7urj5FBQtPo+pZ2x
VxFYm7Sm/I+z75fQvVfGOE74hOcnDaHjpdePYkLvAFnZNaEka5q2BuR4gS00H5Ke
TfqM45l6AKOONy/p+k9vsbMt9dlBRTTIRTGkG3Tv8cppx1g2xmw3v8t0DAk6byU0
gj0ysv2oLUuw8t9c6YoH4NVqJ96BQ7AWnJkJbbnzX3WP1XSJw4/98HGQY0KdAGit
kq9Ls6WnGXDiQABmrR4PYpyirPimhQIJOVTv291B4RgNeHcGdKfr9YTC1pCY/Se4
U3Gi+Za/QB5Zk7W1jc+9HRtHk4xULSxf1UhGgWzrENk44plamZ9nTgjVxV5pyqls
IIXTZef5/mXBGpJdkO6Gm35IJ0jSselmMkvW1176ZH4iwdrbMS5zqk42v5edJ07k
NXlDDxwK93egW9VEtN+7BFZOncIINPeWwW3Tjx0h4nqEPRKC5xIRfbN0/LUOmnwd
eqAB79zWaootOoiSrCPg9k8IT4g60guI86OcENq0vG1TIDIUO8UZrUh3tVhsFbsk
H8PG/41NI+b+p78ScqIXhIYbC6kqvUYM03rctmr3nSAqZjeCYWhaANAV6AaLOA67
07qcc+fXeVwXth0ql0tWHFvp2wXqkgZjHZVRqGvJll1fJcqGNbzQTo3UmciEk07Z
4TYZ16Hb7CQjSrd1GwJLvSvS+xp69NxsKhXQPLtmpJOYDSTysm0/FZVQCZaJTyyS
VsSJn9VXVV03N/O3Y9S/p/dlcFLDjcbKxAl7rCPYG08UejWO9LObQ9CzGMYjVd9s
7b7Qej/Pmecmt3DfWFfsF9zE/LktrBRVoqvoNNcGpxhazMUeWaUqpOVxo/v9M0HV
wecmzqbVEriy5dfpxwPd1usZg2ljGd2KKOYCbUbiMGASr8OxC7Ua+zQeYYBxwRsO
2El41/AldQGb6rrioFRmVf5ibt76lFFTrh5ZIf2fupOuDXnXKm92IkSrKzY9ervf
R51VoYFXtRtHCniWXuYuoun49BPqBA6jLAFM/VUaAfNvX/007AJ9M//mQmTiduGM
0CczlhIcW/jfc4BCxkS1Jg9+R1rTD4vxGE80yHsoDrND+BHfoKg0/ikGRFZYgMgl
xMI9wg6LDGcMZ8rNICyjFYAMrjMevbKF1208LRfxJG0TEfcFlIggfd4fcaGAOhpJ
o6bBDjRFr27tXRaVIrRx2DgTD9wgAlP402a/qvTFu8VkgolX9cGLzsitC2PyGfbK
YPkofbRQemCORKn3XYVSgg+7kRyyH1EMxqJeXQUo2/ZQRhhHW9OSxaWD6I7p19nH
0CTQFnQZO5uefSK5o1UhrpjfwBAklfndGazL6489aDAgM8/IDxDbfdHAV+hTHfv0
Xwwj63lJkDIHTnhf9S0uVcqKkfAbqpaW1sx966vFUdbeNI4i9DdLJiqhtLjrAEgy
gaNAURmK/+5mVKi3gj1nRtcq9+oEeimCsTqa8M0AaGv/r1to7ZJpx6AtMZMb+Yob
8EwEpYUgen/RLk3xCxqconYx+zHi2ZpaWFme7QoVyrBx3vRAj6zMKQw/5IDHu5k9
Hdokfr70KA7CoN1WmIFsoYbOdRCoiJ7V9KaSOdKeSHktxXfPDIWeJ/wHrZiMB3bn
Id+ZdV3FtgsWO0hHF75MRDC4Kk6IzxUl2ucA1b8ImDNd4ZKtCVTpb2BBWsJ9IWQD
u1EuxZ4SRtqGWVweVtoLjgxgJaDNPUMi87zd53jsrWrfgXX3AzYN0Qked7B3oi0V
Curbbos0It58ZbUto9TvWse2tmvrVXRiVdD1O2rUe+wfGGykeINOeEZ8D2jpqqpc
2BsYIF+vnMrQx3YwYAGXzBmhK+0FN2hdIvmeUd6PC5v8nfo1XQCV1AOCtAdgosh4
bvmv1BoGMHK9rF2QCyWX+FgCzIlZu+OPrJpLDJjCnie2bZs4INdTiQUdG4thX9z/
TpwC3X3U7glIvb2RwxKJ2X5GvKwanDPSgrnuzAyBrop0iHe3ChNCOEwJM68OQjZ5
eDNVf1HaQjMKSdMpyhs2Jukc6l+LPrauDRLMg2WlwdhVbsMO9RxVEbdsPcoQBHsL
jUhswMRCTkgrSL7SwNOKMQ76tE9iF1AQ/zUlakbWe2xqve38nW7XULisPiUX6M7w
i2EIxnO99YBwKsfdys35u1X80gkmQXzgl5BaWMGcr/l7HSEpUQXEiw95OjrQ2NYO
ciSgiaplj4E2rNXIPUZ5RDsBiTU05R8vas+qySFoGH7g3GhVtWjTBOY28Ty2Ord3
4Bl8/ujREGHI65IgrihGcO9pJCem9bSrajlUi3YYHt09j+JRHbN2vcP08P06lzRV
5m8F/1C8YIcD8AxA4KQ41rpPKTv5r3yhtuPIxEo1zMWh+zLSyjiRAORE3d7LsWXd
loiMFGDXhquaJ++w90tZRz8/4t+y6xxs3CS9FzhjzukF+nhvf/3xR/kjYckKY7D3
7LmXgh3FHsw7ywB7zGkKE5XFYnLXSlKy3WNQbRLeP6G3b7kNo342OLprQoJlw710
0TrRLW3pmAJSnd1xJ8yf1JQGVK2fCyXnb0mJDcoAAgqb0wCvmfDj30zUO7QUrP7F
sbm1OLyDZPUoc5i2QaAuiQb4oYWC6DrOunABTQtVLlqbjhz9N6uEvvvXSSC1BpbE
6A/BVsewjJccUEBzH0UL8D8pwonzVzA5asH6WOXxj7VD4lD6hXMPVKf5sbl74Y7v
+NYFZqSoMcFJ7yKV8Ib0fChOR7bl3q5g963iIeUI56pgq9CRS8AJsmOhSR8Ln8e6
z2z9CTP47Yta41KPXbvcxXIF04MRiLxoGb20FWhjRQKMw2zDtArL43kWKWLhOPdZ
HM/q0LT5/csICaea2eMTqkXN74jA7MKiQafDmJxZJ4CenKhvNAqBVGrO/X0U9VeJ
FusqQXpUmXmFVBehVogWEITG3CG9+/L23uELsmo2nz0tAxo5kOM4Ky/jn7OWDV9l
jlqHE8SM1sRSxxkQbgI3f9Fdq9+0IQGgYR606dlBDrVY0QCbssUAqqLhrs/aWiQr
D/Zc5e/LjLrxW4lDtMKBt2xdDs2YK/OhvdZq3UGqp8OtE/AqbYmrGjDT8FwIAK/n
3BDfrTp8XiIIxXnecTncWnNTw+tR+uoEVWR1C9yyZossrRL2T3/nsJ2+xoxpRtJx
23/qQJ2wAlseQ//1lqnGaX+4i0bwxzowyw54azYRIdO/n6vnVWRD1ZOYNHExSAxH
np7/oJMTs4yDomqa33LFyQuvRwKh1ZzRpeKpnfCbvwcNBU/LUSnyEi8mUbYw1A3P
8IuSJhKmtRs0s6Zpyl1XaLd7UVvTpRFX33C2BDqTF7zYBYT+lPba82FvKByz/PH2
Y0JJUdtsugBp2S3wgoWpjey7ngCiBl1udJ+n8dTGR/lTekIVWbC64Po4IglA4V3I
DDu8g81MOMGQCE54YrgUBRzkNtg0KkuSfXTm0fr3HxjhVa8daD/2NGz+NOE3xUny
ea4I+u0Mp00LJL/zTKvCWhEl1z1kA+vsM449g7z3y4dxBpmud8O2coyQxp4jF2+N
uhv6DNuR9vbZjXxWmP/Y3d+ucV5BoRtcjyuMlfgkYL5vFpUXDXv395ktLhvfzZh6
KAZXvrMma2tIN/s9zdkOxvbYkEgNDQhUSfpJXatJcbzFs8SG+/SPfXdvmU3cOIT9
ICUaJu8PEJUnK5ky5o/xMC9helkPRDYFpjKEzr9UKPbOAD64/CVqlokIBv+XjzJQ
qZqVuVYIH68MEeAu6iNR6/W9nyMh3bkS5GUO+PqaYPD7HooZtW0hXHbgXcWc1sEI
Yeiv2ej5eBQ6uOiy+3P+iM5ohaZmUgHUcPNFwzqKyqXI/UZF73pyRKlUDU2WsdX1
ym3rGlqyaOwLF2fTZGKo18z+jTIMDJElUJFmJFWSZPcjOP2MZ7pQt22jM7TiyWka
OBLoSpZ0uisnRG3iiOeP1SC/ePflhET3Mrp/ZTgvc4lPdr2w+UWua+SfEz3CeS7P
IFth9WYVo81f7Wxfopkraan0OOQRvgyHj8S34rjWCCAZqyFKtWMjsmpr15Azsv0d
zzZpiVWjPJkkXtJNWxd+z71ZwdMEKiTeryJcVAMAAt4lFilY6LC1MwQmwZnolVFW
jbqcjmuzJEZgM9bm+bSvgDD2f/Owr8NNBmw6cukkiIsI/SL8nqGSuoGdI1WLL/WH
UgxoFNDVRYjai2+qhkDifRDERtocYOFtdR15pwuM3J47FqnesFKPaRCDfELw8PEn
tTt+dGiWVzWXmiQ8Cmgz0lorZODOqVt4SEA/fWUCEOMYLdmoBXJfGBMpwSHlw8ss
DO3yHKFM5+V+VOxJBfR5AvBuN2nJcCPMhLrBU0fLfbSgXomJOgX2TIqF59L6IfEB
GXbjUeGuMLtaLQkJZzmMUCWsY+rly2Qfz0DVc9m4JOYpSpTL3PhfLHr3JEs5nrle
VaanjqVXsTvwEnaBAEoQkpe/K8WlVnZXvZSPPb6bQsRuHPrbUQbHqBG+JF21RlhQ
ym9lv/uHLPy6l1J3vT1dgJyh4+v4kMihrnBDUvfaImM5thvxswaqu3IBJm17EFwa
COgm5rp4r/8hs+ZtcXBXrJA2z9t+TdtcpLVfl/UMaMc2+GfEJ1qBEAidFFa1SWgU
gzlbCJlwbNk3JBbIkP5jGVzNt0X7NGo5BqX8Kh8ldWq46ltL+vqIY9d60hzE8D6y
s400ODOcDjVn4VwVhzpmVIndzPmB/qoIw92iuwYPAtnec07lnx4y9dV/QtAShE/O
QhgxdPHaiyyFaAXxFmEost7aqWOXiPwPAOrZjAnzLf0KyteLLmuiw+I3jORzb2bG
NDOVLKKMa21PXZSorpwVDfoQj/8Q/fchmWhxzLega8mUzYZW8/mPTj7AiudYAszn
U+6SdPRvNk3qr2wYqg2r31mqWOtDH1eHbgrevP64aboxR6FyHrr+5iZKHcqY1oXD
h0rsJwM8dUVDORdAmbybWlZiHREoqZ/M+HAicltijHuKhf+GWhbtclhEdcps20Ow
pYbksaG37vQf7Nh4KVB02zUyDD9McyLhLWDziqZF1CfqW2WPGiMGbnfRyWEassTU
pAbX0fSeqPGOogtJAwqqahEdZxYcXE31NVsv7qiHjLgr4d9Rmr8Zd9DqTNOiiF7x
kdbL0eEDMBHxnMkuG4e/BnML5ahLXuklXourU0qhZ2melV3g/NVgvFnuNaCKzcWa
8c8g9GOxQMebHYIewjk3XYao6nkHZhkCwlqsLM1qkFETmI1x2ZMpWWTMBO56WV22
bIOodQ7y3jZGs3Zqh3bGkMWSVTwIGk07rvg2OYRerAcBJ0lBAbRvM3JZCAyg6nNp
9dNasv9n10uzaTnBcP+Nxeh1cf165CYE2ZAH5l9GN5FDhVaq9M5PUi9Is5mUQZzQ
VxBgRU0H3qr8EndeLqcZQcDHHOQ2/IcWUB1VsPYyoXLWWJrsNZKiBaNiARXIUTGe
OdE3feyyVKo2BAp2bioNbnTSrnAklJefNHkq78RMWqLhXoPPBujl0KuuLg+cNS+h
9clEKTxpPg0vZDCW1keD1wfpPebxHWcggzSSBi10Wd25PQesTqTgsoBtDWf2id82
kI/0QG765pxdhcTGekaFflhjYyITBc2Wv2dHLQZjcVetO+qqUVjIqTBJsMlcwX6q
XTcVQqbRPwKjZNRbmwUPRV17VJdthXSv2O/oqslnpaHiSbl3T1XPmcxGP0L8XmQb
TcCgKycib54cegJzTbyXAjMTMFiz2SSvo6ZBNPaNqad9iwB6cgjNDdkzF8gpGH8Y
YOyUuz2W2ggUTPpZkBcl6L0TcMhnAhsUsSVIbZaIUDo3VxRvyJCG64oxFo1Z9XLT
y0+sCrA8qjV73xFQYGPM7+pM5j5coVRX2Fx94z0ITI8TZ3xWJd+Bm2rsSechAKle
rV1e6Tq5DUgn9STg+M2qXxBGoPEhlPL+tMmGx86w2Z89ZwICY5ZJFIjE4AA7fb7V
DNV32zrxPtdlA7oLhz6HZujQI7JsghTwBlAssMevf3BM6UhyzBTZVE6T7tT7UgbG
4eThdFW2hkLabDUV+hbr3yVT+PYLJUcDBjy//1IfVTUjvakRX4TYcXH1scTYdCOZ
N8VFd8SleulcHckWvtQ/vM8lbNCaOJ+BPwwGg/L+N7D1re/f16yJQ856ilY4l7QG
PFb/4AaJxrGGjCWsjvrT0yAHMpGUIpOCGOJIqw6i7qwGEPYJXHu04nJLUfYNOOVK
9lYeBLUlKV0M8dx1CKIOdTcOvpiQhGMJmtVi5diMENqRMYzDoYBWZDqABXYZsbye
UcXZ1CuJhOm8GpUeIDvH5HvCTgDIevJOIKSY3aLfgmQClqnR8MnIGYx/Wwzd7q/x
xvxNt+uEuWEQmmo0gfY/nDrNbPuSgog8ckjtsqVMhxDBCte+79Mj+mc8nIBK/PDG
9/eqmAbS2Bq3vExHG/4VH89pwLZBNJJDWVd1zFXLUhIe2s5MX8nlSF/wGprrxcrr
fzojcsp2e5Y1lzwRKouwyz6DrnQyf1l+BDJySewKx3/iLP4FL7sV8VScBoTe7+qb
OkuTWU86mT8OPdWanjP5WEINnOBdwQcCpHCGfqhof7jhfBABfIBtE2e91tw/wG6K
NaMyylXGbH8iJw4YtH7b026gEVvoSeoDNFbtEdt/4PYrGcAJZaXold9cGJgeNOy4
XulglVuEWAJrDVmhqfq5CpoOElzf/DTD4SH/BIqbTBR1FbCSdPvdMMJBD0qp0YQd
AlE4LC9hwqRtmFXuOZcG/ZBJwSof4N9m39BQkTE3qqIK29MaZLpkCbMdkYFRKOKs
zUOtL+u1+lh4nFaxfBxAJLKrmVBPHEEjLkfEeIj3Dvs/YNTRPwxtyKP7qUc4lD6x
jlP/+dM41MCP2mT9WdkEvdGEOhy6fCQelUOH/8/Gv/mnBzpDGLvNUy3MocehK6Lk
AXOSYCWCr0be2IQE3OXsbjhSwxjXT9xwXzjF0GTYuakAdR0e3leWIJSovKKKRfS0
MTUvwHR0LERBP/tN5Gkwsh7D78pGJkdA/aY9ailDMohI1qvJ66duFsry6EeK5DFN
wW9yPA3HVn8S1bp44coRC63EaP5mUP5wvAL+K1NqvPwH9TUKJ+q28P4jKTmslRWe
BAVyJ7s8m4PxjxIcroyunJfyLL66ONnu8CcGcKQaqWiau2YQ+whZX0VeJXKbsNAc
KMjnYIMEOfFAFu1VgiB/HDh27vVRco8Rft5zU0FJBZrakLgM/6kwjL3k7hGm9I8U
ShgHvaStuln/ODpvVQC2Nr8jxkBSSi5yt165DosCGfrMT0yEueJLljYadkN9VETt
W5E5dp+auRa6AR8EjIsiiOCFw3H22hL1gxowaEDyX6uqvmfZXCnEx8mNbwUPJVqF
ZwkvQqocD0N/jdrCZ2LR4bpmuMSslgKmp0XThk7KEEjcDijVZ+VnWA3ZIXDF/kWR
N0gKlv2ioueaIRkfyq1nK6vvhPv+Y8Gqf+bixDIm9MMj0Bv2fVOUXtWrdxVvntEo
lxjH25DXCFCYmLpQ6Z55qbqvYDSwicI59WxbJuhg4pElqeSVVNQUNvfZjmRRL69v
/ju9H1Yw6cqobARcHYwqslv/s33fuWr3IO1b/U23yK4CD2VlFo3vQqMnG6WWxJxq
X0T4a7m0UmZhgKjw2xO95Ztbfd4vybq36NRn9zcdYgO2p9aP8lMotKYQa4phrkPz
J/5HVB2WxpcFUtLas9RJMvY9YYhW4A+7T3DFXUn+28Uf6y42WUaLdS39jSnFaj7C
z5kWuTFYVzjOhuvXsW6aMdRwyNOXC8v95l9CqjVdvhvN70Mf5mH9E1o4tToxk9BK
4IgaUL6hm6lBk5l+6RXsAEYadFqZgqRxLtrcjBw38YvCuBEe/XARA6Zeif8CtkFO
amfLjKSz2ZD6Gu6jOBd1EY+d5XEeqPWu7r4SVRNvT/WlF1ArM6rs7++7RgtIL3J8
EEvhY1sKqzSdT6vAaZ0zXVxbisQW5otT/ild21osV/JTgG9zyZgkQJBryq+KPt6f
rSuN2Z0WriAjbPZ9bX8EY4iWk6KrsXgkHNpWtC6ZONc=
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
AJBJcc6Cc9pg7pQkBHS1SGzzAcPgScCs1wYtZaTNqYUj1Lb2f+aqc3X9xLlQ9QeY
qdXUQ9AakNXWtEocKh7i+LyjETnt3QK/NG1hCtazH1dqwybmz9VNVnAzJLRPWzWd
ipDaqHWkb5FbA1vntsWoBi0h1UOZVf3pfuiwWUvAI8U=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 14751     )
d1r4J4BT07eG28Ebmpw3r++YdWRp0iimgjY8EZJP9E4jGiImHBSiOpvUxphXq+P4
WbWwuBePkU/j/Gif2W4Rp1LnTtgJpmkTSmYsWxgUK38ksbcBhIVuhD5OSt42QzhS
B0h5GJtnsUoxo6aKusW4jA==
`pragma protect end_protected
      //vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
HxiKssREcIGHixQWHHkCb/0zN0snojrmqCGTkr/PvVgkhC5+2LXV6npCI1LMMKtQ
aWwcKFGwNlyL4E18xgpuOopsfJr6O8cy0NlMAW2pB3GMwCRkIRZIiNsDW22/QAk2
p6wo6Pvn9xkJnuna5fchYHuv6NBb0nVGYq01WEHgPB8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 16397     )
V37Z+siw6LefPGErU/lppLUGMgAQsaoBTTQ2cVvJVd1ZDncWwEfYFySw4MW4kqYI
JpL8iFaoV3SGI11oX7K9OZ+6Np53a9z+v+alDgC567s79fmPwpi+o7ZQHcZiymtX
NjkuzdBlUcdvre0f1DWYOduvmBAGZ/bKsI2rq8L5C6MSN7Tlox190O9gbRMEJ2Sn
e4vTxW56T0xc5RMT/aX+q3HujwvP2148lx19i2FnYd4g/JC7ZWYFRrdwN9dRNmZS
QO20twBg19/Z+iMg2US3F2WoH9Q9WJoyVftI4fFqduTfZ9wd+T8IH3SjOGNjr3SG
brjU/6fWUFMN6rG8gkAAmDUChFWvI2xvjMyhjtnlDWBwRbqdgWLgq1++lCaq2y1Y
qPOsMi3tlLrHEGm6/9+oLRhQQ+Y71Yd1G54Vy/jkyPPPUR8aGig3CVElQGv5cpu6
985bIn4bc/ObbcBsgpBr6B5ZW2IFgZxDjT85MVkJRKoaYvOPI7LnmPX6LcpJhSKP
ITaS0cbw5rIsaGwmrnXkhE798VODc/tEJg2DNVruafEvrsXeUTCzGBO2AIF8MIzn
CLa/ZwQjMF1mWOxuT4holSXqy/nmg/CK69+eUEW0ZsR+Qw/METECPDeRwBSJ8I/H
ANj/OhbaxHFHPQ6GaOf9hDnFnzqLCYmAIFu87w+kdLj0WGLHPA3/3z4WmdPNO9l3
e7rqmMO6/ZP4F5xUBlovbLY+mbHZVJJ/QaJap5nVeocW+gqhaKgOTcFw6UaWcfOa
ndJ0F1/0dl1x+zLbydYrO0m/5nOBgYGNS9YV6CZrvL467pgFHCPKhQedb27Mi9xj
hygMy53Iuei2++vG3P1H2+j+esUdY3DqafxjUe5qB92DBpgktYwX/skisBXr+Ec9
jhD1Xsi25vz84peRV0vt8PyAbpPA93ICd+6h8oesPybpj5Uo+V1bs/l/HoF/3wWm
orugLjsgsmt0eM4aCo8evi4y7/ZwB6nAgl/MwLTwHDA89++aX2jKnbigUsTAbQeZ
ccQTUg44NlUOu1+uTag2y+A9k2vWSRLF1OgNhMu/YB8Jox9dkEVUb1SrDmTGBlWJ
EzVNgJXmbzBgw1MEhNKvwyQutpHYFQhC/VNYjf+trhj8l9K+jYj2QeqakQmJyyBG
vsPgosEsgj5BhY9B1/JaQw6HRfP4zcv9v8DF27vHZu59YTekxYADHXdBFEfviNOa
fdJE0ad2Cmj76jlKQE0izQ+2XipajBT0RQEC4/VPzxGcyEbpG6+pzxwlGBis1/bG
Y8zbpp/soAZH1W2fGQR0z9eYWlJmlFI6v3NHsiWafqCCxXZzi56zr4D6bHFz6EXa
BVRICqBpMFExu6qxLTJUsTM7bZq3PmdtL9s4/NqnfhvoO1so5jldr64r7rVMdKOa
Tbg2VNncDr8Jh1ajKxBCxF+NBTbjRqeJG5S1ni3qBx4gaKKuqyQR6TotUyCK2q3s
4F1j+oD6JiLhX5bJi4rFvGDm2evYfSfYTsGODw+1W5vVNxDMLW8g8ldoz/6KALQj
frMTE1/CX9GXnXyl/PtVE4wz3Sj7Zsn7ZZ0azG90K/XUyrgntk1xqcUBxUgYL18y
KpdS5jgUDlgUo/rQ9G5wO6iKWY4/nDcSF8ZVOVCUFjF22cGlCuWqxqv2yNhTkKwW
6/KjdQ7rwXI/0hDvQl+ZNE4LSDKkwzZVAwHN2Ej1Hj9urfz3ZHFOTYfAF2uJfhvU
qT7wH/wRTxFoEVR1ywbg6bDBVziXoDFIBpeODfCPcDQUiWmr/CclFWvTIhKLpgto
jEeOaS4v+6kTne3HCh88avANeSXQNDQ2AgKIAYa97oNO3hvqsjI23kn0Z8mHBxyj
B7a6mr0e8emHlaILVNcsJT0AgshnzOqhfkJWnRTXixMWnVOixl74HHiCstOcgM5O
YPfMtt2mhgrdILysmjf4iyEJ81WUEBNzwvOsrvBFqGQ+eIJeH84CjCvPjDzqTLzJ
jHZ1+OIqR6AsPsyg9ORcKxcM0K829+3LxT5SwIbFJGlGDX6mkL7YP7g7YEdRn0FI
3osD0PxiEdWbvpq8DraJh0epNfYNnZbTBbKI/mPMrSvkYpsrhUiipH0Xd2+OrVxU
qIYZ9s4fTyS8Ox9/mywcgL7lPZwgcn/5kZUuPnf3xfbifh152ik1L1ot0VtWJqSh
b1bLBwdastWq6Gbu1C9rfw==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
AngpZLGa9sZqv8Lr/QJenR7d5MgNkeREuocGHHhoovHZEPnhfBGkSosresgqnbT3
ZuPrQDW6OFQS+0dIe0zDBV9RE8ENTfT3V8NlDQStQOl6Xmr8loc1HbJZEVf5eKPz
LCM8vAb1GrJXher34zADQ4qdiZwBcd89qCLaQqeQ8S0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 16506     )
4NQnXU5QmRsSEr5oaOwvceC2QyYO1k5MKUpO/26gzAHKUTFUYx8Kc+swjjcFQG59
DcOpH662Qq+lRJRmaxgOgOLtUh/OsaJilUb/RF0MrlP0+bbxbkCDQXFm+Gi+MZ/J
+5Umm6w0HBG8zfmLzk4G8g==
`pragma protect end_protected
      //vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
fx7Mz6LOCwdaLePS7aP+l9h6Zxq64KqRpUlJU7MZGgmAJ1Whi/wPRtBrnXHG67+o
Tz3K/zR5cYBBKzzMXX3gA5NYQckogc8Y9KiUev8HlFQilsR+A2/EjiIQgXB0aStN
vflSyjFZLoEYyAvCEUahDoOTCns/AqyV1RLaYp5LgNE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 43529     )
p7PH7jFhztfDDt4osb7cHC4a61bSrQOeZ00G16VB0Ts3qRnS9yAkcqpWe2wxB8dN
UkS6k7QucjlDoz46IgdDh8TiexMNDdumUO2va3SWXSHPYqwRc2uYulF5wzOKg8fS
MUwMmDD+Dn3g2oUJmVGdjghPjBxhHKUy/RF86UqSdhaHfv7jxl5xrmyYBdkobPNI
IaHo8C93Jun+CqG4nJ/hrpVBI7ant4eL1gIF9kJ0dcNhKLFFYRDe1DgtSJMkiLqz
1xaNWGHtT6AejMEvSPLJ6qmRy3iHJJ0hjqLhN7RGrdDDWAj/OK8Jp0OkDsE2fJO4
8vHPEyCxiTLRae3OZgmw0NQUG4Yo9HXy4gkJxqR8TNIiBIwqN+LSKoS76wWxquWE
wT07X5DkseLjTK1ujfvCZNlcGLmQYRjg9jAzn4jkgbPxbRu5deZP8C2TfyD6JxS1
hFm1C5CrjjzMh3DpjLDIjxvBeT2/Zcq1VssqIYaBSl3+uc+Rg5WI1jUsfKc75CaQ
V7BB7CLlvS6xqLShRTmARiR6NquqNiFQsB+T+O0UXJhCoW5jkjbap+wpDaHplDcu
30uXooQ/WM4zWCjGEj5TFF0tNMrOcerWrwKZRqnalogYO8pmpGrUKsXnVr/NAdDH
e8R4rXEwCjzMe6PGk/khO0m3f9kM/ygS6WjS8gR77a0PWsk7pSpqOvJ2uxVUYi66
w2W1qG/Phspx+PjOaSGTb2RJL5nxWFqueSuKXfyT83UQbRTsMUndsXg++GQPnPpR
bJspdeFGUAmk5yagZb3STyynk2Apg4FSX9eXK8A4flt1Mo7FswAhRyQoECA2Pnsg
/TqGvEm0LKTUrl+DkdoSL67EbOwakA7YdktXdxkEXUurKhU7g35gbtajrlYHXdX8
ykNgN2KzNzdh08yJOoYu/NFGnhkS/D7xO/saxjv5KKCqT/1/aQimtN3fSZau5Ayx
9tXpBLDxL/5/f7QgOvKTzbt8NUZIxbZOhlCMOgsrpuLATCxNonf9Iv21QsJ4gfjE
YATXa1sWyBUeHOv8v2UzHxtAKmRSnyKJfUBLGqkPX88l4F6AauXQFOhnfD/PpzXN
vdhZsv5G9ABb5lQ+hfPmkYHgnh69s6QUjYfnpwzwNVrwMgdL6sQVEFSxOaIL/FKr
OIrfsRl0sdOjkUZ7Cp4wCO182Y8z300G4uHo/NO1+BZeSErAEM6JLJ65AoHUzKp+
i8GqJLFJTK7S/UPM2Qlak0Qs/Y3t+iXwhOttZk0+uF/w5A3k3w8LxdaJe3B0UiQx
K/QAIivVr6jmPHqVj/1XKsFBrURcOdJBeBgZRBZg6Hv6UvuO24xEinoFP/XgOrk/
RpVAqUlvu7zxccU0ihKYvmGDKqqe0XBVROB3NxHX6WGr8s/roCtxwEF2Clf2l9RZ
ljQ0kligp1UwCXZprnqVQLS19bmllZn+7uuLWOMKvJDBh4AfNmeu93xdtfp1vNMl
nFwXgBo/gJqsUIT8MQALKQ63V40jtEPwSM8vHZ89NYXftntVI+e6/odlJZ5aFnhl
cidqC98le/1H+0qztbwLpJx36OXxMVDeJtgSKFqvBTWwSg29O4XRLfAeS/OWa6YG
k9Ji4pzr0ct2yzEkPh8S/XRsxxTh9kTMZal59HT3WmdeX4rEb5aUfFgbyB1KSIl1
RiFsxHNbeaABBudK7ydrg5fAfxXOPDzyCZktzyc580D4pn9tkl5xadH7CltMlr0R
tW61eml4D0LaUdteY0BXYEWQHUm/ojQAeRsup8JXO7y2FX8iUvqftw6lZK3hW7s2
wczBypJfW6WnmVw/2Iq65qepRIATaZAb5b1Sl0Q70ikNC82PQeXJAiC2syBOzs10
q1V0NLIfxRWF/I8dc33Fm1FVnCq/ulQFOWq+XvxVMhfv/jaYiPsyEnFtQEs3D11B
F0PEEYXa2+RitUqWLZs/J0IsG1G0uDhJ4o6eOPuryukHsERAJmptaFcKe4VMil19
NTYTjI4pZXMMjoNdWGzuBabOFjxcz7N7hM41r3QUK1b0ksJgcNtYVG/mrHfTTgt6
U+bPbGGmKFA0FO2x8WZ3xh8gyv0jpoO282kHknjcJ+zlhZXX5wj+126Rv5p3jup8
p4jZn7vfTMzVX15zCCtJDjAk1Pd3+q/nmuKJ1zE4okC7B8QGTe0wtQZWoaM8AUA7
SU23Mv7TjcW141CdP3EHnbUP+ihhN35QW3NeAvCTiLw8aInjBjpwfbf97iy+N0/b
AEfr7LsHxJYYZf9XMaCu+tGzKRXv5RJD1kAXWWgH0raO0cpGXRaUee/bSjrnSep6
Y449QbwZP94KSWkZa+TSzJDb2lOKeMMTDZ6fcPM9AaXWJ8e2BEnUYySn8fWT5fdz
JKAbBIrryvtHDVH0brtUR6Swo8yNltqbEy74oy4hBhp3rVTNFgjCHh9l8YnrulAj
MqGgkzZVbiwv30PU0ZpfMllIpGAG2PnHIDgEPee0asX0XkAcmVX8PB87lC/upwsi
0yEuPDx0mUnCOTVRYDM9LhVZeCWt847d//XCM7KwAi05zvGAB9dbPUoHjkTuplbE
/T8cRDhUtBZm96lPJf+XMcVQ++QxVGxQcMzJi+TYpaSGgN6FSC3Fk6PdOkpRClF/
bkyv/1INvwB0WGGwiEw/6ZzJuz8jVxF3EcDd7puVzLUJLbgax/TA3QbIB78x/pgt
4Aca6ReRbaVdGEUruKCEpOKHwsm2EzhEu3ZlqTEJFdYSvgFypaxR3jxKq7GqI9CA
e4wkW2XIBCa44dVO/VHZYlFfTmlBrEwe8xNupRNGtMH3Xbf1ZYraOQGheVWvY5sp
ZyJdZi6twgyhw4Dn2zhRxQiCcHAMqU45cC1Ty5UOegdTEq3c8qHbJOLelFhVbC2o
+frwXS+MW2RDMRhyFutCVXIAV09i08+TjeTXYlJPHwfvvxB9bywQp8wsxShsEcMD
zFzgoQZZZM3kIrufgQBsdI+TbyGhQB5gr8eTUiJeanOd6yNpbD5QGHjXr90OLqyF
21pYBTDfosufGekWYeDkWqG2Utr7f6Vjcnl+8jYeAOj1MAz9CY0jKCYPex4U66pR
Zij51AvfaXY6HV0qJ/YARUhSEc2jxEM7PDsvULGeBDzfmFn3yVJvmHEucTiezyO7
l+jBQIT+IAvA2fwMCCIGzsYQ3dGTtYcT/X5jtjy27mzeobCj6iqCQXTM4cbBJBno
8zCuSOih2cOb3E2jKoTFcv6ttvE4UYmRcbNtypzBtVhABR3i1+KvTJr+OdiFpCjd
w1kZgTuYcOEQqXC7uPhWlCP5zpyaoUmbNE+5MrRFKTwpTIaRLEmzG7ftgYTEcAJR
ZLKxBiCDRWOzDE05f+nxVerW1UmuKo2f82wUqKvkJzwYDpx/byRQV2eMyYLtR5pH
llUI7/apRX2t+hpIXCduPT96NTRv65eqOR6Mc3IhuQtOzIiQkR1xx97EZuYQs/Ef
r0+ClAzTBLqzmr0CaHRtYVeD2M5SAo2RC5l6UBVjcTImTiujzZ4pb12/IU9CGa4L
gVznXZJk3PLCThNKDtfa0mWGFpEq5iOApAfsGAtyMuqE5hVCc6IRnK1GJUzPig3/
xcBKrqSQTkZxyhSNYSvGP0DO6cT/qCqzxk2pwW4mVF4m2jYfIuVv5457rayUVAcf
G0zaVPhECaJIKRKnOZ7/Fh/Prj8heVzFuuUmDrWv7II0k+hq22nqsDLgiJLaMVlx
QAl08M2uJ7OJ5B6do3xDnVXTcTa6znAAhGKRvmC5/58GD0dHE3eKPOFwwqz0xu99
mBGTc5FE6sndiH5TMzhXjZVfITG8+pQYdOvmYZ+WGHCNYSimpii/1Y9Q75iP4ntX
875dBLQDNutFdqT4HRl+VoVJm++2VdM0x6I1OAmSnN//eJuKgGkjUz3NARwaTNRW
cT/gXrv8JKhiaOT3h8po15JDnmtMPJPfdSN7ueOVxEiwZf6aJxVS/qtUSTt/Se5/
WxVy7znYaF9dtOoiytCEDzmDWD4Sl59cmW0uVNDNm3QHpfEdqym2urwFhj1vcp74
NQJOc3JBAexwN5R7H3aXXZoLl2/xA71HGUOZyJBVQd/JKCTzJrxWwjj1MYVzXmAV
v/Bevyk74EwFDQdeAk+9SSyb2Xv6Pkc3pK8ohlnNC3I4DqtHOBbcyPPetsRJdFuZ
kRQs/oExDmUVM4PjXy5H9/h6yx9f+icfFDciD0hePu4M6IS2/sw1P+0OE30BUjUn
GJM1LHUp+8PQEmKHSuggrDAoq3P61Eru0ycmWGVk/Z8YcYnVN9cfSJnvoKV47L9t
JlPyxLNecZGnaFy5Zq04G4BiwTYqObHkoNX00cHgL/2PUswB1MfDYjnn/3cA9e+j
uVQwTzCarcl2WzM+UqHD//Os/kfnB5zFuDXd9fC4KYEQtoILP0XEnxHDYHtQoY8/
Su/FH9GSLNV9noXzOrC3lynmNZr3yfvjUvINx+tv03iM9dGDTNvcdv4M6OsAOIo+
YIzG2wLznN3XJwlnwrmvpUP4IOYlgBwecIbOD1En2z2MXlzqETMSXyTyj1Cv/yZ3
dsMF5u3UmkbEHh4L0h+AtORA5aMB3L7dkJsmYOujI0CKlSyosczWffkbB6JD2HBE
ZhVI2vdqAi/21AJ69UdwrKwJzprYkx+3QxYTf6yFYanhqdagbSAWz1+CPYUR5OkG
kutcBkJeCejDn3K+d1cZOseidOYik85Pk93J8+IkZ/uauccNuxI+cduN5ZGwFPHP
qWWp3+YvKGvJxJdPts/WqzAfX+LG5eYmwzVuIS0MiZaahHOT8wd8oxtg+UgsHP7p
pcPinIcizt+GBYo/eDJQ0Kmq+jev90WoX2xlz+taYx3T0mXPDJ5E2yeBVEUb8IlV
WB78+qpI7zyl6xBBNKnAAbxBx1ymYOP8TY3WWC+XwQ8BXVd4vrdu6i0YcRlQjKPY
4LR2ufUtcb9ZFfgA1G8udS4b5nW03H67co8STj+9vIq7nAi1AvNLcIncp+5KkVZ4
douFJPlZa2iVa0n9N/QZca8UVRk1VkTOZmofizUXEwA0twihZ8+GDX+WePQxak1H
6TAloda1O8hZMExZLHUQamfm3ahS8NPRu1/MFWRyv9q3jhatSYs8A+WuU8Nvtgyj
iXHih7zRhFC1uPU+v7daie1sHu2pg916Vmy81Hm2bNGGmYwQLV0XkJiwQL/XJJY7
TQpD0tY1lzsUC7uVGk8MiQLu/0jxuHVziItfNcBeGz1Bsx3bKW8pVv2rIaq7I65i
R+7NJJ1q4wURDkA47L0IqNZDxsX6GjRXfW2LFxM1r0EvWwYlAO0NnJkCpxwgDS59
3ZDMEuq1+pEGc4ul4rEjB+Z7MUCQ1YBLTCaZ2XPhDgThddSEszoncplLMskH9Cuk
6VxxNzvgiPW4w1rLaxkfbHR4erM/M350M/r8WcbIf8yLeCAjf2WhqBOgJx6GwYF2
puJSQC69gWw+WoypRJBDdqJ2ol7iDaVLnq6M2BZjv+pT6935pofWgKZj+vFI1UE3
VR01giFnfKZsr4h0BQ3QrgaVni5NjRwD4VJaklNvF/qEIp6uS6ic7VrlA/oz1jLw
dUdZ1gpe6iMxuu5xVHABfvgOx8ONzWHtZvbFs6tC/iTT8E75pISTj9VQE7nGDjne
V/3fph5Z5QoupYOiFYvfAv8hr6KgIH33BldoDeHoc/15KsIRliODGkaUCVE6Dvf7
34q/57fgMBqzzKWUGN1DNjztLxHAUtBLIDZDWhuGC+XGeV0ZLKdisIFrpGa/0NP3
jzOWx+cbnz5zhXHQDdp1aeiLJeF+vq386JC3ydteR7BDm5j0dmSSGaYvPJWPd84M
zsoP3xkXVcy7U4UwUjI/nSLPazLbtX+pfBG8zLHR+3a2q+PcWVCXTfvV/6CP0ZgB
R00SBqP6r99NAsyUl8HZHa1gU2kkfQShfEBzTTW1s4w3phJVpfa0QG16aCHz5t6n
S/kuLSL4iPf27ZpcWIvfLdi36eRx22biOwZFl8Zom0p0c1EQib62pqkFkEYehq9/
A76YIe+xYv4Mb+0LHoFBGFIJ2j1FhpP9I3dtnJI/7T4f+bP6Y/KuEJONIOvw8mfD
9MkGhxlc1lzafX+JGqwVuFY7LuVK1RYzXd4dwaYeh47LYsPOXwASSSriImnWuu2a
7Jdnb9JjO7wg9ksX3N6BVpAvnUaWRAeUudhqjOf81eM+RpFHRKhXuq7TxXgDawKZ
Z2mYN2veh92BAtKb6t4Hq2zyCpzm4I6d06E9u29zj+p2uRv5OtGdUaCzznU7A1uU
R/p1omYVNMUQ8BofCAkKoKWR3qo8LNlyn5fT9soHvE7tknRQqaL5MGuPmkqHBd5Z
OmCoxYscQw1qwMVaO/S2OUo0Vsxz1XlJtmMW68jRcjU4jzJ9WX9K7NdJ1DhgyZlx
lgVkficb5Rb9H2nGz93dLlPbQUCInpgg7R2pzIBdoehQAO7VsNbxRvMpMo5fIzHi
sxIZ3Zxx0J+7k8whbojM8UI/1Q1g3wsnCed6hrxCwu0EifJB7m9WGTQEFFB51ReE
0aqLdCYVJs0w3O209GqefW8IRrjvBIZm8Zjuwcan+j1pPMAH9r3h9PEpTLVAxQ8/
qLrxncG3AiM77IQtppnMYVaBFuRCa2Em00/o7tdESstIfwpRh4MClQuMfFo2htVN
S8/4cYOy2omRDtFjVqbGLUBb9ie9DwRkO4DESDfJeXAvRGmup5Bd8PaSC98tF7IC
+ZxWIv9FfO6rOf/eWXSIEIyTAQSIcxeuF1o3I15ne3uyrsnlcZA+atjiev76EVun
sUT61pw4q7+cZga5276Kgv1t7NIb3DTE2XJg+eTNR6a/14Zh5PoYs22nSkvGfcJw
7E1ydvWsTFJH5L1qo2Z5+DvY8eV+chSM9P5CjeMdXK7aIpZ6uyioh3sXgawGBmSJ
hKh/1vx5KnWi14l63mthw2F50bX5f/L3qhBDKjPIUyYaSmkkAMQrYz3JFNBnrn5h
ZFpIiZBzywJEc0Wggj8y9Mf01lNKEGl1PouWzVLdpcr+mDFYO8eRl+1cMv2Pqfp3
/KmUvYC1E1J+EXeVSi3CDxwhyAn/l5tJ8x7CkKB+HgmFaVdWrXXlISVE4c43kO4h
TBx0I4Re+tbZfatamZjHKcTULWkPXLVb577dcQTVEATNUOPo2QdvAUVrxmbOQ//G
Txir7vYLxoobPdCXaUEaSU2udbwglX/F4fVac6hQJeYpJD/NcD9SDf8iz9Pdoo7z
V6LtmZ0XusVxdzBEkbYvSmA82Vi6TIQ4WyifTZJ4nFpDi0XZxgJwu0m2SRudbkWi
SpTA+OiEd7+HaKS+BwmX3+MmNqaMbr362g+OY5sHIlSeyK5SVyBUAT0n7qRbmz3n
mkyFdxF9MLIFsijti6s/W/XTBI3OLE+Wj7oUCrWuVsS3p9/BrBVzQN069ncaXMOo
7DKPxcf/Vj/7Le2gzRswbQ/rKjP28jjHnboO3xlsN/YjHT0j8RfBgTqFAK6nqJuT
u4qUsKLHGtcPeAwYTSImYdxPWidHa+eYzxsbxxGQTEem80gPgADOI/92QpUr4BlD
3NDQh5NbadagLTWpNqph5SyPl7WJyEpGP7doAxNhAURvb7Hird0KGkfJUb1aM2oj
PFwox3+yVpunv7HqvDRd4oLuN34kqGdYXcy7k32wC+87SYULQM2ZHvXBd7AubwC+
gzzvRjnLqCzOxO9NIO6+AixEiyI6fkDdUURFQ46noz7jwU6MBh+f/F2WTyP0Axfc
7AzkyVQcqBtSYmdsByPuEB3h461wulJydeEn/g7WcYW80NmnCRidesOGaKSC1CcS
3DaHhR37YIVLIyB0H0+yTSsymbgi4ZDX2Gw7AauiNzsWCzJApZILzzcoUVpZu+PN
trrWdkCOLBznU2F6X2x51Y69RtrrHy50q5wT7FxWNyReQMl4rcsccl1Yp5RrQKhb
oNsaJUZ8RVOy73zSuCDKjjmKVJ9LtSpMqvDEGtLq1kWE0pUovx8vSc5wy05tbMsw
YrfFwTZAZkKL8jK5IOXnBw+4PEMg5CAIzh6w5JVCNOziJshsD1PesAlkIyp1NEd9
DCp50YYQufWRyIqOMqzTKcrH57/0DJ/A0OgIF8AqkFn0/Cy5siG5p+LGatfopNYT
k6RV8m0w+KRp/sER3dwQFk2bP1IzjTHHCWfeCYxWguQJtDwIYVYzx/NATYbIkM9g
lBmyYzBri9rYlQbinlKIAARnat/1Szqey8T2L6vfpUZ9CsTIxTEu89vbuwjOJ6nG
xF77QGKItoRQBZ82fz7+gVk4Ws5xAsBKhzsf0ZEGxmrOMgScoJTdzq3jTE72Etfv
uwdZ/mKLv5hqzYUaOq1CzTAcFI+WuF87jdUkclAuwN5GXQnH7nui2YPgqSK+D7SK
K9qln39li+yANkTINaA94hamqxwzJt/8TwoJGBIZmZ8WZEVgsDF3CIM0Adj3fi3a
Xf3c0L4hGHM8e+RtFD++ByyvKI3UwySzC4rWBS74TfPvTJ6PXvFWXZjJd4yktYem
mnlDTpKaaTjQiTBiGmr3DprmlmL+pSVT+ti4flqmtEijtzpHcAaB1gIk2bhzbjkQ
DQcMByZLSzttVN5var4+zdogV+xUQ8A8VOIvbpf3v2lpHdgdQriOC7HIMyiyHFJh
BoCygknPEXtajBURxDVPb0Fap5hBufr9g66Rq2jcTo93D3Eh8CYhF6UJOllMCZIG
eoBAQmOW3VLRUlrBuYUdwnqsQCJo8i/ythh2Ym4MNhF/L25zfgS1SMfiNV8Kh3Yp
IZbfMq72piN1eNMYwyduB+JYTiqpqLfeoaTCcL1TEEGaLFo5ZxOlfenXjJ0soLgt
kDyhSTBUsdR2cXn/OvMJKKJLRVgfHDEMtP4c+Ae0upJBUxO2P0UUVIK+2Gy2nvKu
ui/sknvJLxBYz7LNJarAZk1dIqIpVeW9JNcJrk4Wno8pq+7jyjguQfDhSulbVxKG
pdvU26Nh4BISbOQ0yBOl4A2Se/B/7yPjlp1pakwUoORwQ4evvbXNdTpV66ho5Qi5
wa9/FAHFp6TkC4cMcwjBZ+XxYdiQox06HZ9vixkPTiK++tgv9PA/1fV5i2tUdCE7
UfaoWOGG/7plJGgDJbwp6jkipqpL3UVbsqS5WffYV92p769ISYvN3shx8aawvLdx
liCOW6TIv5luG6/YdUTxea8SbbqIPRZi3y1GgyUc0jFfd8oN2ng+y45s1aHg2ZT3
ZKp0QS3T53VaMvTUprjnWPJ/iRh8vNgygUJWKD8ydGdpRd9dzivnNOgrd15YKcxC
c84Ksaw7B/OTjujcoVGIIkwQuDxWvQx0TwZLuqkYqqnyVbFAgog4a7jKe30pxzds
yoe8Unk8rABrgxeurtc/S3iANtT75f0wmeizwNY1/Q1ZRXiM/D6ofDIAqSmDE9Ez
319gTg28BaHgv/6iqYsHWhJpCTPoiMmO7BrJTvUjnPY8h1+SwaGqU1fUF3XOrIUw
b6EGn6wIvuCzpRvnCqITZcDF0+bDbjvm3iUsEhu1sY4X9fWNj5xCMpBH+ysBA1S8
tjARGY2+JkrHDbuaOD4HE6UakR/w16toHCsHUA+ZwDy+GjWcZ8h9dz4RZfxhHIDu
3t0X6OBEbTdCepsomPpdxdvSzu57AD1XdTjoVwwmHinQGvDsv567FZfHbWjsL9z+
uTk4is+5V9KlLuEY65P6aZUTyvmWdc6nEKqUbJdpcRNDKM3GZPg7XDXJ5SpsKbAq
Q/1DTfRyRvRPmzj8lyfwI78RSpzOxx9epk7kO4pG5Xcn8H/uU9eGLZgnQcsVOe2V
4260kHwB9A2Th5jlRq5sC7sUTG14ywLLAvG4olWfdvpGqNh9GqzX2/QSjOVMhhlT
3QD0OJB6LdJXHuTfoLpQ7BzCpcMYCuYgCZKUpDlhZx0OjkbKoWT0/8zBRcYvoiew
NI82/qX4gWqqT1h/m70wkWLO3QJtV05g5sgUxTTGXK+Egn3yzWnim9YsxkxOEG4K
KmkG0/YRUTnc5aF8V6BswOS5XYQDptE2XQJaabBq9csmLQy1/g2ZmxzCEUGEDeb3
UhYFsnFmBzTREwQFMlWGZrhCwKHLaPA3xGaQDtLuNtr2NZB8V+mi4AOCkoctTWL4
CNfCTZyDBlgyXEQmAgtZIF68MviSIY5w6MPI9BFX5xSTtTYzhE8h4Cb/BVgeoHjt
ylJQx+nAxutyYP5lQXQamtouRQKOleFklXWxcUdkaCwYa+271xmhJNcfjasIIcnA
J8/CRNLb/U7RVMnJiGSWamxaLfLEK+sBrm3dK4KjwG6gh5PpZb8fm5QG4eYIR3Pt
CUUSI9VqRSqJTaa1R9QMUevUIv7yHL8pjDgEssz2W4E2P/t68WWyHZhPiD0DHThI
q28bjlcu2WTChOFawuyYk4WJ1x+xzEe1vwzVqk2GIARQcFfykqVbeBR8HJ52yIO0
USdse7wB1d5vOedTGzGDETD2SnxyoCt/HSq0Pj6L50eyUKi6MR28UIffGPlMJvLj
bmgePqDKPLWeuG2jab7MCOHJY3NHmMjMKyPItQhZfcTsdHlqVUFe0attK0VvEM2M
R57dGyOImgxVwSxOsZl7zS0uip8wNwONvdvnLyXS1USpthq3nObysOJnesqxfot8
ar7Omhvlz9f0mb0klz7FnU2Ghsz861rDAOeThk6OpyziabI/jc3ZPhJwhLjiuuQb
3rbeuXEutYFhqRpZRBAFc6dENxSVKxsAPo9E24vvhytRJQJwCWeGmQkJ1cp6y/kH
SURhQjvCUn8ptNWFly9BZTZgJpjNvCL2iIljjCuMxiKEI3FmbrRePKINZbUYeOYZ
UEBfbzR1onMSn0a5lwWHmKAegSFbptPOYXSKW+5BNpqC39x8ErWDaVDfV7vqUMnE
OgGqFd1YLGCve6zTXbm1Wxfx1lP43QjT8bzbVH0Vjp7U8n6BVd4oxH6O9aWfExLs
S4ykZOZA+TebGpjYW+w6zEomvsOptBnpS7rzqsIw/Ou87Ruy/J4YrWBhLiy3HA3A
0BuXxK92A35B2eXsuxQ4sg/AaGqRQejPiQmqYBLb9VzTZrt1/p2K84vWmj20n+qR
tzgo5clI+ZS4c6j2pEjSJXXnZeKBaWF717gABiX+QUV/TO6UQRk2TRqUxX14rzE+
82FHuahJvBF0Q1vU4uV0hbA+bpfbbEB145tmsMb7vy1257iO9g4pa0951HQXHlix
VE1XcjAzuhmR/V35e/dBSMX0PDkqbratKbETSiuRdgr9GfETc0aMmAck8aTryGBF
HLS9SEe5J8Uoyx2wmzxWHV4xUtitVeZ/+kQT8DQSjayKipqZCeXWmMTKIjIC1Y5S
06tEEusJIt1g0RZOlzJA4Fwvft95Q4ufwZXAZn0q1uho97XOSKf49wx69azPhqHJ
UT8bBoJnT6wKpyDINJiXXWhetGK4wE+O+p7MA8KxVuYmXE8bmphdtmmet344jOjw
tHV8dacO3WdATny+GuVTP8in0LCH/uTNQA2Z17/IhDU9fj3F9iVPc0wRp8q4/+D4
+GsTm5Xry0162wYHgmse5e6WsSGzXO2w5P+W0ijhRHFRJVQ+9Ibkccxy5cn3bPvR
Scu9b5pQqUbSvvlEE1iyE/6sy7zCvSQ+/bZzcrL4wTcBa25Kdn6oQYr/FS5oGVGr
bRaB883VXEV/H6Zt5O4JBg2/ak9vkK/oGdu5NHCXE/70+BZLoKSRdagx1ly4g/ii
jcoZsH2B9vOTuyEYm16mdaEWKsunWop4lDb/gCjiJ7Q0tNBdXISwUyOKTQE+CEzF
DIUenn8igCV/xVRaTpCK4blQHmoBqxpwZozv+V8Y6ld778ag2zpWMReTyHovhTny
s6+30WHuyrxNpwyEYl5s9HvX8R5C753mnsxXp6GxRo1xZ7NBiaRmyguoFKNXFJ4/
r01+iQIGG6czGxdv3YEtiQnedzRABtH7+T0fNPSpj6FM3XSxdP2BqIoDUS23szaw
PoB8Dk2bEV7ETe/jUeyF0MQUP/Uxdn/Ok8HDS0Zz7ZzjhHz5dq/uGMTicFh3t4bx
8qalRIusipjVc04+8KLSjz4vOu2C/GV8jvoKrQe5cKfPy0h9xScc1GHtITmzCdgu
OVk973GlL3QOsSokhMsIWGYREf8EMbYsOBZm+P/JDbaSajxtBj2xd8qDz7I9l1lD
ravERePpW1eltd/JKhH+2qQOJamzu7ESuOiW/Kel/TwbmD4NY9O83O1URPppBB19
ppFVLWVZ9MjNGzZMhzBK8ea9bfxdxipLI6CD/3QYitTCNwePcFCGcmngQ6g7BWRI
wb7v6Wgfzd/my8R+vS1SSI0++v298t8lWjzRh3hhR2dK1YcPsn8Hk3LT15QUNtRu
asXIdwKCDMqCDnAPK0lZ098e2B59h89IaL40eoDTWQdUq4tW708Kopcof64ZXl2i
2lsB6lkvfNXsl17MzDFym1ME891Xpk3q5QPqG7IpvxSbsvbsgWEclFqPVcP89gQa
2RF2cUrC50RpdIjS7VMbQw1mmVoO4sU46DLPPf0Rrr5/07+6lOIIxsTi2klxR0d5
dEdDd7Op7y6AKxH5yrX1rzzopwHEBlJo7MlzXVMVGrxwh0NcAwXv0Q4UqY7WZQd7
vdUSDd1ye6Y0nXkr08p1XVOel1U+lVLbsL05gQ7XNPu5ENVnQ+oqdKg5MweiWQJc
r6dCGGpEcGy2LzIaAmCx3LnQjLo/hbpqnglFU93MGw9Z5iaIcC738qdfFUy/jTsJ
Ei/iOsecCGcregm10O03jx36dBkO08OertAB+oSmjX7/RD3/lJtvbj22yVlX4gVT
SFNIPRrRvXqUtb5JpN5wM6nccFB3CMEWykZAzNbee/ntE0VbjhRJhlHZynfyyazZ
Byq7HVr6ms3Gfx64A25JiT1r6rHMiNnWmVtfzANZFcdEBM5XfpBR221x5/NVG///
Ya0pEHFEw8jb0NOukntmiwn2PSdxjOosgjcOkGtV98YnYXs2YAFU/E4St2H/NteC
SO1iIG1xxYb/bOAmzpf30LKaTXXwripePzb7mLuHXdr3lN/u1cLS2Xgnbxpg+elo
OtHxhAEP5LQzEpOdGwWBbiIJHz1Ficw66m5ZIK7f3vUYqcCCJwfu0kycZrIK3cqY
rGC8WdVl8GupP2n+M4vY4k4EE5MnebEBTCiSVZ7oIRCSpxuAV+/QdbEXFp4z2dET
sN6S/qRBvuVw1WNmIidw68JmruXAYO7kcYaubA31WNQQt9meg5KebOaqFwAuuKkx
ez2wUOTV7LbgNPow1uuscrlCd/ncUbstyTdXFXpnPssGUKAjB30NT9BWKd0+Fq4T
1W5NsEkfMSyPIwTQygD1p9X4PeprD4a9SyVHFFM3MyP4y6Kftn5DVbNlAIabaJO1
LNEGsRpnLHm0YsSDl7aCTjALSTDMots9r0SGa0uIkdzOcLm6E4gqPyoaM+aiZGYv
1+ahtD6Cy+v79cPLCk1hDoNB3Gf+BYpudrflY0xcnGg391xqM/zUOwtsdTiCkcTm
fxePvddYsb03GTPEUEwla1tQVss+1KMvUmTScaNCGolX/mWChQ8bmCKNTVzRZwhr
C7z3NNtpXfy02DCt7ih2V397txNOhutaPgi7IA/iFkAkZhKhzmEdGfoAs0tUn+ep
ZmJKRm4pIW61GLPlzixm+0iv/cwp2ANQWKnK6P2+mJWhB6/QWEP9uXZunYcpguTY
M4ipxwLi4fDSpFXxPcN2CXRHPwp99BdOgBKJ9LhZdDECj1gcFnFtqqU1JNO+vKhi
4v3dZcGLIZPh2399Kou9Bh/0gSV0pawhildR2DM5aOEuQLXxMBkCNWflGSVNv8zb
oPMG6uCz1oMoSO/u9QHbEFeJs2QHb+xcCCbB63ccCKVKLbecUsKWZTRjgmEIQORA
bjA8h120JSQJs9FrgNyDaswtm40I/fYBwRsd5XE01qUyrx6wFvmD0tcd81qgZhqF
vkClnzCwpi3lFGmtQZE8cUr6xNzN/V/JKLXjbtA3NfCsIlratputPq2N1+8ONzaN
GJUPnKTjUsTOCXY9qQ450u1oZ7Fu6HTyURC2fU2Q5E10V7XC3UWUd1zW89HLyqop
7wwMQ4679nYjSuZwEpnWZYGIS5gjnGk7vclTOje3Vuj3fl0fule99T6pllnIEoyf
7jtH4K96VouY/N56wHvwOafJUrFWAboaOY/z/hushkj3ISHTDEdsi2nU/NoSOC6z
gJ2dRvzl+G9H2xZfU/xFz6NoavFHq4QXTvaxt7HziEQsykt/1Ppdqf4r9u7MEqvr
egNDmoaOl0x8Lklkon9X7uUQwIY5fAdginfTPhMLUvt3l6htGODX8R32qwd8A8du
gDifnXrT+JwX+s/eAqWJJTnugxx0hxfhthKODlzSb3QsdV+bcyNIQgsyHlsxaex/
k1LcVckifqcHFcZEFVTKWwI+IsIbGzG4RDkVxqk0Xg0EpTdlc6o1vw+bi7m7KGFB
Lm025ez7BTDXONDW7V0qQMdCSAJeS2GMaEx7HzY53ZWoFJim0eI9qkHjcrW2mtTb
FmgrlSeOX5mUlrLHclgiknsjOnwKizCrwzEMpZUIs5+S3jkIv8i2BbdADTGY70nE
3l+9wI5TgYpj9cRN1FKYTaBEiNupxjToqXMEZJgIxo6ZSDIsegn0mDNYX+cbzGvG
Uj4MSDRDcAu88zKDjfnBP9CDtbFtIryHMznUvqYILUj4QrZs5f+Nku0pwNV9ptlb
TE2+1dYsgAa2Izlh7g7Ibr4ZdYBM5TT7xRpmU4cO/rEWF5uOHuG1x4i4qIdxopNu
TdwqVelBL68S/7oy99LV6cdVI4KQVEIz9YXziUf1GS4hoE/kDtlprilcQTCGIpWs
SbkghhjRo28w6UEoEN6nJscMgTw0Dm1Mg/d4TQ2QOQsYpuNdE53hQyeuhDvWP0mZ
IG7JQTwhwWOc+2DzzONEM9s+ZS/of6bO+hkf+jF8H6LcS1xZzsx7fv/iSZ4cJRi4
6gRYd4g+KI8QfDHdnBtttLp5UZMgibTp1B9p3plY1e07py5uM8d7OK4elqHOHbsf
5J/yL7h+kXL/cNYCM9WY3xlAROE5idfNR+cAsQr8EzkIxCpDe1sbFDsBmS/LxLTQ
YQSMRUZddjYSFed+t/GeI8R6CZgD4YGU7eNjNDgkM2R9Ed3Cdc7K6gbzvOxjd89k
aYS08bZJ3d2z0Q6JngU3T26UKBVqG5dBKldtFVZuugrfpbNiRiwu6TJgVq9POpbU
qN2mxWh3DSyo2ZgXMhbZSxpRAsJEYuvQFkajomnAYC/UapsmytywyzoVC3XzykhX
aymD7MmGd1zf+d3/yp3EDIaI6nCUgfGFXDIUuFm5ZPFVAzALXfiZ+my6i/Ght7Bn
ICJr5lLOsO9sNhnGvlRsUBDsbJOB5B2UXK9D6eBOsRC9NAYlL5SHytFTVpCVR8lB
WqNgZBRNLCjOU4niLfefSbq+0TvD7mf2LWCDKYVpdlM1oqkP25vfBzEws28R+SLo
bycXre/LO5ogGv4KuREM+Fac29M2p7P+8UbMbADd8D0qmC4C7S7eBM0hj0T/0RO0
3CAXTeSR1OfVwMWDU2590w+uGobdaUa5jxbABaGh0aj4kLBmbl73fN7w8SQiE3so
Qh6S8eEB/oICuA2LU9tjX1NlaQ4p9TrMX5fzItMtdQ159VE8D0cLe5jrTQDOvs86
NgPJqEWlQwcGzW8g2cabI0/4xURUIGrd1/rLP7TEDrfpAWKf2FOHLzpo7FLqo9AZ
g7EakKMOLQnD0iE5IDx8WH8hK8E06heM3p2YAU6M5C4xEdN5MG5TBipN6Ev09swU
rPx1VNinLgh32f72NWFKTTUoEqaA3U4Xx/2s3Ui9J7HvA/bVh3oj5jwqi2isVjTa
YnAqy/r6xLeuT3AgnRjs+uWE7bvIACd3lF7Tw6Du2LT3tjxRQQN3SwpeYybfjUsB
SHy1phSpxNVyO13r6RAgSAa1Y9KWcF5kGRVdgQXswCG1rwHyv8n9+DInirxhNcQK
j6rpAOWLUY05kmRgT800J7NGsJqlcXwHKiB46udI+KLQZRXBSo3UWU6VbqNmviJk
u587dNKlpOP3hDYTPV7Ub8OPEzY47pG6wOnQOuLdsxxgDW4TRgiQ+y/Zo+XPtQyG
baj4Bl7IB/izUVBbJyLmQMARhpGxrb2ZS9/DdI3MTOPWXQDKCaxuHD5WRIaZ5dH6
fWYAladJTd1AyQVPH8IhyqdViZXWL5BBMLgtu72FHVrfe16fr+MnvuRKmmHG9asw
jySRWHa1HUG69opsJYoFFB/B8nRAre0vm6rjQNYuVIA+YZknA1sB9ip7l8a/15rb
16s90AhqXc7OIjsnUQSzfYQXhSTSavDgYPj8MivNZVMQ2598yWYshS0SM3ziFN0s
V6jLJnVXwYIysS3m7tgJY5IJidsul58dFVBeDg0oXYhDRIXHj2vPvdoNqP7zeh+g
r1HE4KOuztc67nyTXQkuWhTB9qfXC9+q8RH/nCa3hUpVR6Fev0LtLntfaow36+QZ
bJiOBCHGdRFJ95/W7fmxWeMxoN7WLH9fKxvUDRSWk255qRbO6ePc1PtiuJ+zRxsI
FkuXxfJAS1Kxy6lZi9tPU9tGmj6mt3LYJS5So1w1jXsQ5PxeSYO3C5kCIexolT5I
VU4IKew802e2XHd+9Y6vYt8TlfLUMSb3WEtIYiNJ9rMan0T6bW7XV5Fck/PCLbyg
2FyopRR4iBN0nesRSxPx2UT2jdHDcfNQ5AFo99SCVecCbRPgKY6pAgxvnidYgw41
h8z577bbMebCjzpDU5mhJmQQMjlZv7KORObW3I+M9wUu6DNlc49B3TS1xZuh8NPC
5+ZbInVOwmMOR4pCxujWkP4H0SvViqQpSPHEy1QIbcwOAcDYP06GisfkkbivhVOS
9NoG4o2tQxFo+o9poJXmquNeroQ8da1qJlxbu2pLx4hg55kgtlEAZVXh3Z7TVHs6
GV1PqgUgXQc6qwBF1z1UCj8Hutet9Nda9oQzMcmBIaSKpMGWPX3O9O6WibZvm5uL
pPK65OO/anM677HALhOxuTdGH2Aa9tGz3jMBdynleq9HolpD0TI06tWkJpvwbP6X
ilGu1csKozag31aUTvz4NR9vtAIMp6ISYEaoZ9NwuElsmDEk9giNmfKIqlE7xqh6
PQZRCGvyL42xzEHplhi8jl6DVkwdsQO6nJVSqnKELrGf61MiXe9zujJRLlHfhu92
Hfs8rc6V5wqHzn1Erfch/Z+5XmKQI8MbZ2dilRTQFeCWbvlgnVSXhvGa9iTVncrB
V1LyAQyo5H4Ujh6t5AHq4Pp5cYywIyWDEfYKVYiDGXB/DI3tM7vxwfVAuHjlWxTr
lMmmtmf/PeMO3fpD7mWGeHX6tWOv6PdRHP5nkfzMH/zF10gdQV59FIoTxSN54hEV
5sObNdzOWabHCYFPtIP58OToRU9xp+ZAM5MTo9PZTRTG08ABzHeGGTCLQ0lSANz3
FwUv9Ec0o5qy9QWUvAs9+7WDWaal3WdEL7vInOHX3al0m+cQrdFSGeY6e6MzN5XK
sXDQ8ga6gfyazaRn5XDcF3B5VW75d2YPa63ZA62qWG5t1srLHA6cUiNeVD9b/z2m
MLokJfLEsCo7N+FK/kMMj+5aBhhhgcPtq8OgRQQJwbK6RqBwMfeOHIHfAj35QPGJ
WXAPE452LsgxnGAlGm0AaZgaL/bbvzNxk5s54pWrVSstFjjwTXZFcpIe705OnB+8
eP4cX2rE6At0jUU0rzMoIqfHEJccsDvZyZITf+BUi7eKv7acITO7ZCmJpZpa0Kmb
YXQtQv5FUOZzB5Yzk2V+nU/F2Cr2obhUif0DztaMVhXeL8EIugNklBzUo9AL6Zw7
1VbS+INT5mXybJYWixHD9kvorSohSTvttCtZgJxPYqfb7S0do3FEESKZg+ZljfoO
N0+rDfwjGSRuhBtLSBsEf9P/6sdIn48FBHBV1DRD4PdG2anA3kjgY21+06L/0oUo
CpUdxb29FFoWjmXuOP84SmNMYkbj/9HX5XSvsdPf+yQwXU7zb9wDKODSojNH6M1s
TXTZkSm7GW/khkPzgYsbpii8TZdlU3lLlkBTxNqB6H4IkAU0wvF0nKnEnaaDDawR
sVmVMtOSop+p8gKTWF2/3wOKD61miqGE6TEcYRKDejET0MALYpWE68Jgj2wTYcpw
a8SLKY+baZyH0gKXdf4o0ByHeDn2jOR+p/z7RHeHWdyfix1bJim3i00WC1ayzsRz
89WX53YJU8GU13P7xfLCh01+9VYX40ZwxS8p02tLBs2i0/SDzsSxP1/AyAvrr6FT
qMkEcBJtogXyAyCEo+YW8zGUTMC94b29n3UnIg4eOYmlu961y2zRukIx09n15+cL
xmZC1cSxDwim5NfBedv6rVHRM6XloUQzbfqVYuDUshiU5BIfjCW7uXOGRt7WEYLN
ukpWflKLVBZl1J5CzFZoMS4hd81sblDRDZGAmJi65+LvUpbieNe6Bk4ag+WNbDrD
/4taAeQ3bA+ybJXZ4R1ySaIi6r2RKhhhVf2WLduvzTUUFLTrnnUCNhZEo/gTNqvZ
s89Ke4DVozZt+1AfzeuAVOr/mPMKwUukxM98UbcS2lBIPgENIfqEM7EivNMj5a5B
qpSVCd5zUsfXDrHdONK9abyZ3o1ZY5OUy8oiq+kTYbB9s3tQvyqa8lDReFUnLJMI
h/sG6YuhO+B2ZsLh1ba1K6ngojjyPm0P/wrH1p4B+g5FhoVcS85hQK15ESU/TeGz
v4HYZIClMmGayKl7QRyPwN27QBv67vZNdQCZKWk8NlPM3gNdCB91gkHyiblsNd73
VuQ6r67zKexalkVqlak+R6lUQ/01Nyo9Tk+QDJY1jp3X0m+M2ceZHBpkmdhTMJDH
sRUlk3/to9+vR4jgaHDvmny2IDS8qtIbMWgmATKtgiZeNXMKULlOuf/kBdvnK91r
HnJm6CT9JQrkEBsT2mq1E6uOdyKH93mfP7oSZWs2bAgU47a8ZtZjSyRt0x29Si1A
PgIrT/MJPHWTazaDYMPP0XNAZvrVf50csFcLXi2wvXGG7oZSq6fYruBluaJgcrC5
aYll6Q8Ie3IHwF44NY/5Ishn7Ur1RP8yUs/6GYcWN0RF0BuyX6LJy/tUabIBLVAW
2CbSQ7DDxz6ZaNFexNpYhvBMmE2bKbw3Cr6I4M0waJSwxZEyBRtVZZSyspuCisjf
xgVwJ4Ql80+8iA3j/aAjly7QuK+1GaUzRWI5OYTovkEjnGv2Qppzg0KE7tu53d7L
WID1KhGafKOURG36PdW3k43H3EMnYQS24BIHLgXATQ126iDzF2r0ToD3BwrcI+oI
8/gcFTh+riJJcrVQzzBGI5RoPZGXDf0s6ena3cebUx4bd0y53Hek3W1LGRmxWzyb
lqXEI/T6mg7Azzpd3wLrfzRSvyylhcNmSTMmAUydjmQr30y0/4nYJMpKp/ims+lW
uHhYSBij4hHlEWmczlnhUDNtVP4AZ6+BNIejdXJmgseEKJkGwnc1NZcyHpmKLMxM
ucJ3UOKBhtEbqZPu87xxJWojdwpGPpRw5ibLrASOdz4t2RC5e+GQ+SW4udf1z1ln
HYWd1oNvC6rTlIQwoRtfMitQ8pz02A8AEYdRDHs4ykbgTgy9Y0vigd5xbhb4kjBQ
menJ68jM5x2SGWajLzMu+GM81qEUAb2RuDXMYlGuViuj566O49pl/Pw1fmDIhtSx
eVSaMkk8QTZ7iF/SI3gdn/QS337ga4wan3SgFPtFIMzCvoV1ctCYQwE47Q5uc9HZ
hLTo53uModvTPk/gOjcMCo/TG+ftWvTP5fIWeknhQdGL/YHqi2gmhCDIjQEIPkPU
TBDPp3DeoP7vIV1IuUGaIL6xTaxPSE1fVvNc8GXQ0e+NqqRWXFzYzvs3eye3SY4y
jYxs+7dYP6EKgb+ia16DJZYSkMAfjnAoz/p0YoIdQwNinFvovRZoX0JbBNAgs7yl
V9W7WObUkJJIF6lOr8NK8rq7bgkhJmUESfkH6ftkvI1NaUkXgNl8fXjEvfJwfrlv
EjiOegIXIgBTJIBHkftsOw0MeucqqOWBfbCGQE9DsY/sf7Ir/LHq7KpWMOvw2ynm
M8BrYweV2aYtQ0WhHVsAMNde8h2m8rPx6rN7iFaGn0DX8AB3mmt6uEzHJCjXiuJQ
PEhShtMFwRbI9IuCh3Knaao2Do/dXbgN455Lx1zw7cLRCzxDT6tw5FBQKe6Uvssu
0tpxoCdwOp0HJXaQta96owZ3OMMJUUfIwAnhACbu8Ho50IOHNmYkNPHcAOCCcoSc
1q/ZKhYXl/EDDL5NhoUcXhfesg2Tyh9zE+UhttPH7CgWEzzj3AOVONpiGLYKRXw2
MgGMeoRuEujQ6F+uiDf1Dd7Ye7Mp7HriETgBennozby2o1KGLcmTBhJ1ckIkfDN3
P9uogt0VVgQnxS0rdcWZCb/27Pae63e2wUBABuRfO4SqX9RY4XjkAm4RuTnL30Xh
6S/Hz6YsVfvPCdQATt+ne1DV2QUm+Azm2Tz09jZ9i1ELMyrUGBedLXxUSl7e3Qbn
GX1OP8rAj+lTyHYewQpaRQjuDkjd4oXwxPb77iNNR42EdwRrAdoUCr3FpCRLxYbc
MeZr5Sc+EcN/cfpFU9kxKPb5cX/ttYRKLdQfl5tkLm7up953u7ST6Olgzb7DiYJN
nmDMbzGIcbEH9sE0vOP2rDYQYh/oBhbQhPhkJ260157x0qBO7q0nRqe1b/BFMFnA
EpRzpXdtHFvu0u8PM0sJ8IcyzKNIcBcBhJrjnVlABDd+Cz8yBzAl/R0RXK0WJJKl
U5RT3lchVbx4emwB4+q7jqUXGgCD58PsbemmU2m7ctg3XmNBlJqvSf2yScLQUKjE
FQ3qyhBjbcLcXE406CfYXhVWq4T4uHEPiwpzIYUHCGm3ZMW1+gX5GNLew0j5jQNY
PRDHrR7k9KgQrJv0/HaXtaPWiMAqB8Y7kQ6b0cqHW/5ChJxbrg/hdxbYkS3hzKgA
GCZrRMxWTauy6pED1dLqXq8UU7bCbCQtVhiC53wtg2xJdWSxIPEQ0No+a92pXbJ9
K71skuVmE9jYr1xTVdLi6r+dDmkczjcqaC+tpYfAbphpkKXS3YRAjG801zvOtckI
GOVIwSYJfeauJ1qngoPPBuRJqjpGGJpNcLbssa/d5HpALsBcnhkKMCgzWl7Zln0L
N3EcUwQjuXynk8Y/uCG6NyWZtxIRrCce5PPj8qnNoBYl5OkFs662GdsMrXCHDlus
/Y4eQhWiFfMU82CIXBhSL6ldhE2nBZXriZxJ8UWHxcphzItMqsM2szIrdo+oCMau
8K9ZyhUKrsAwzJxQEOHiP1k6WH/liocRMdy6tkHtMir1kk/V4DjM9dMg7c9JIFKs
nnhSlTYAH/l/EGg/eYjYQjqtfNvmH+Uky/uKHjxVpNBQiIwRAnA1sJifKkOxU5kh
LO2iXzYe0n4PSKHrk7l5sfs0i9PqXcP2myiYq9z4jJlSdOTifWbckH638mIthssM
5q4P5ssvFBEKQZu90SfmWty2/0XeM34bFa5VfM2kpOlBLBPd5lBYHg//cGLv/GeZ
MlV1ZIU88usfzfxnnnB1ckluumzmZEebsaBCU3tzKQleXNCbNqRLVsvVR1w1tNa6
rAYP7YwmpW9Jsnoq2iYhLW3Eq/bosfIl808BhHhNeKF8MvZ8eSb2TyW8wWvEDE/9
XuAnfh5qO04SKvQccT2os4QEhQfccAswuwg+rC/YC+Bzs1XUaUlD1FTC2VvM7QfT
bvdc0lETRAnwm//4qk6c4gJZEHMdyIHWGDuq2eBaOxWQtd90pnrAgE7yr3Qdn8XW
wppWiwKHJ8/maqdkC5fpoul8//dEZ2zhq0wdx5kbXNOTu1IC93q32qs5ZENpLeZI
5Bdc3uVo61GNSsAhr8bse8RS2waEi8mMtaKOE9YdCs8ciQWCy76AloxKKzXae6NN
TMQqzTxzgCDIz/OF/7TbkTChujWFdDbZpxF3Moh8VNkiG8U4mzsq99cp9qrILmbV
1RXl9V72RpbDYsw8n7zB29A+yMNqPBYz1xNFuqB73W7klJjXs1MpXC2+0k5RcGty
LhfhlgCmFGYGbTIk+XgVoT5kC9/2y+4rxtBugQn8lMbj89bI4fFg54tffU5oKoHY
9+h/t08Cy0MLPmFrEvK0N4xxbXXhcsAy1jbx3L0jetkBKLKhcW8VzFZy00gmlcA/
PJiXnD630hz73LHoFrdtNnlcQAvEQmHrRulvCudUacuYC6viKa87Bfp77HWuSo/8
6CyqMqdanhbwzc69iEnGcg+PwbcvNZKjcbGQdwhIHVEkRcyR5OgI+QdnuEpocLqP
7lPMk4JC7RKuI/9L+B465Y8wPgmwQ6I9C6yJYO0UkFqh3HIzXxuY0kys3mdCy2f4
T0qaOhp/BjKtGNFCfpei4LrwLc4U9neaavsrj5quEEDMWCSMhaK/x1qfyxN/a85R
PGMJTY8eu2ZcKRJlWQv2pBnSASRn3hI1gdkDZ+M2xNiCaWjTk9kZKHD9txNVKjmU
UV2UD1vjL+rIj9vV3CFNg5GOuTpXQm8bH6lw5UJM8gn9GjuE5iRP6FM0PA3Nex0r
QDBqgDydgszczvEM+AyS6lkV9ZpIasUFvEXQmrwzIp/69RTfau/C0lwaqh8x3QC6
gvhqBZl220mYv+bFw1vk3Xd0PsR2Krg1IPbXc/oUxwVXPlSlTkHbDQT57ZNnvlyL
zuSM7zx5NI+Ci4wh5URVDns26QFhYv+y7YN01TvTD5xGHgF1WHdfw2vDAg2NspUx
KGGVWQcmU3LSQQqdAAE7jzN6qQEEGP8AFX9cLG38WUtnioEAoCMuhm4yZbO2D0/Z
TPH3QyqWOBJmj8MsDeF2lEJcmnbxeQj9bncZA10D2AwHml2sA2flAuFIrNuzf5CT
/msWlmn/OqQLuaThuZWMuCqHw/xzi7IOn2iNiA+SdFrwztzrpsdlj5qKdqIAtVGt
/SC2D8VikmGnsJYPlOhLhiyN6K34iMvAA9oTZOVEIZKDJFCmNqhHs/nWCvaY7hP8
vYDjerb1KRLbeTxyn/S3+odnYwWN5ptzqGL0yoPN+fj7+7pGvBDKvoEFwz1YOKBT
qK3kRTBXOwirdXt0uSoDIxDUSpLLeYRW0FdDcSd0y1kdqZBAgYLpQ1gSc6+oZ7l4
l6pesUC2S9ZCNJ5P5Cixx7JNd2jyrWoeE+yXgjYD70Pz/v8vxZZbSI0kmS9AqwFI
ToGQU4o8rZjQDrwaeEg6aptoCOVdOFRADAo+cbS9JMtg9/Nbke3OefOFS+sH58dZ
eoe+r+MeTXyy/FRfOp+odzebDqN9dyKlbjXYxcbJU2MZFvVObfotwzVL+L87kEQX
k90oHzRaGESKiBniH0uj1bTKGfc0U02Y30R7azsB189DQDdUSVC9PQx0UkS4b15F
lU7tTBtUS6uSQm/mjjcj2U2rV5aWH9ldsJ8z/PUJvR6dmpEftQhu90Kdbul1eUu7
D55lGrSUwUOi87loesTW5mV9jKtgrU3rPVp00gU0NUFqYsay68vV/lT9ctlR+k/s
i+eGp6XEfcMa7pU49uZfZpnidjcfJPj4bn4HKGnBYrnFSHzyVW0cCwrM7XX14D6p
dzzUb1IUz6AlM+NkOST3Gl2ECwsIyOGWmeJiETKn/OMnKyHtaLsF2ECGz9QLL+vW
nAkp4/9iNUy/oe2lkB5JADRRfFFrpXzgOpB+nPrT+jvHV9glt/w/R8vRyUNw+MBn
uTfqP/k4YExsDwiBAJ0Aa2lLdw+yaGcslejE7O28NgN27b+9adg81C+RZKlj4gC/
/HsbtOpcQZqRRAFm1CI6hSIRzK2gegShFPDVcTUmO6RfzCVT4UX7z/mw/GN7l7RQ
4Wo4KvyClWB2ZgYBpM6mpFKlPwRjcxaxxDlvtW3pkKGBAVgvN5+TRxIcK5vR1XqQ
LFqdlrAvJcSz2gqUXZHyC6u/2XL35KmZc/inbE8nPcUwHjaPV6QFeM8UDm/A+OUx
mGL0XMwg4VjW5jrblnbJDDLYCHoAdjIcpp5JuWBQoUi8M7DVljXhh3bQ7Lo+70aU
6i21DA2StGhh4Qi2J44UwR/8O1WKDsb6SEV18QL92X4ZP1XRZbLKW0dKFfje+/ZE
AVxsymcMFO0jEezR+GOo+DqPYyXB4xlnLMenTHuyZfaF33FJiRKnExbI+1y+Qqw+
pRgxTBA7vxODW5+WguK4oAey3U3L9D6mL5IiygC1Cp/MHXl4XD24TbNzZbfGyS5v
6qjJgcuEUEDhbQwprqFGg/B6DVemNrFbb47jcW8EN9uytfUfj1tIHaovD2PqyHpD
5mBiizrwqPCY66pa+uGrMnVkFWFCAx0KUHsHytZjJKbL0LRuSzik6zdumNIYvgIV
kFk4ihJuOKjIl6aY1c4POGtEpDiZ2Yv0c94dtGp3Bc8B+oVOrd1onF4vI1gsqTqD
1wRn4gpzmb+md3SQO22/AaGTP1aCPfJDqczn7hl42CL7ri2syoUfFx7XBlI4gKSV
Fs9QdMWMmXNA+OX4TOtq3kYj1l47qwkm+b2MjAX1JcgZomNq1o+1ORrwmgDvJoef
xlN2KOlAMXi5yFnGEwzS5/oRgMnkXaUKR9dskZ/uxzMJAREKev+d7JQ4Ej3L369w
1D7voLA5RtiP02+kWQastjnwWyUf34Zb6EfgGKl9XJJr1f1fQhLTGn6IY2KAFQM5
h0xFuzrTYHtK14Dk040ZZoE8Qr7uiBFi3zQx4SI0au/9hpXlx9Qo001dW5Tr+qz4
R41eGpeKk36yfTpswGc98U7Gwsmdsl93E311my6/UQlz5bzoR7my9mRoZOwe/sAt
zrTfgyGAKhhpWIurHzFRCq5FtqjSgWZi3iAu6X8b2txQHnwOMpXdKaEtf0Twajhd
xZDmeGVOOyXM7Te8dnmnvuF7u0K/W0Xpk9Q7MHfUjgDe5tTC5kq97Cr2ywI7tMUg
Jx713U7JoSn1Fi42fOhir/5MZ/5FHRFqoASD5N1VZoEk/wt8kyjEFrY2yo6wMl4s
Mo64eg+H7g2CBTO1BGssDZcZRmZhL3VGvh2qs2oTszRp5OQydCa/13/nIEw7KNOU
SnbCtbpJU2H3ZIS+QK5gxwVmZfdrLi8Gusiitgv2IfNmdldGjT6H0P8o26DGepju
aZEIJ07cL1L5ueKgw52b9WNuEY9ZEkClvk03601kT3GNwSPQmTKp+6QgWlMTz8y9
RqIPuUpjtrIHXqlkdbJ3apdHJoFWMCyuHWQT0+1vFFLiHMUgZKkJoUcmW4hp0XTY
NqW+aJ3cAHz/EzuG8uA8ugFcr4abuTDPh4USWgk5768eCthJGT39G4sZNhqtTumG
LqpvjDLQewCQWZSTx9ElJ6+9lKHpS1qzxt0ue5VOml92+MQUw9bL5ZnFBg69rRkr
7u1E0o20bZmmQpgk2lZRFUDxX/DIIDjjSLx8aCV/4hM4Wk7b60gF7qMXp1oStKRK
H54WmMMZrelbhFH6pFpG51yMhuUL6/yRb0PAHnIX1Atwp+IdeVT/hn74BNNUXsrS
tLF7CpDcWTjW1WV0jzFNWyv6T1G+xh4/f1CGVTSf/ti2YUoN1awwtLDL3FlU3rf5
EFDTBs2RxSSaf7IHHtKU+c6ex6t37okCTsGyhKweGzGsHD5T3eq+3Q+4ifdpqfGt
ScNt9+sS8vMJ32waoVfW0j4sVMvUUrhFF6RUgKOGW5KYa0HT3PM/+xBuuBlrvbgC
LqOc88+/y4oaPqkASKE5y33bVQ/3Vsf3oM4hnZDz3K/epKxgjV5fmyzZUd8pGcD0
bqOQKZ2vPf3/AVeGlgjq/3U+4mGYJDiXsof1naibQsImNfUnamyOe5Q/2C9Wd5qC
o7CyhVNwHNlY3Ir22DtxO8oOqyjrP76AuRcmUh9DoV5Uj9rUBhP63oRmKuONBsMG
m5XCvSI248vUcj71cpn5looLLfMiz33vIDOoePlh9UgqNOX6oY9JGoDIkRQRjTL5
yKNprIMMuiNwLNpq7SjxFTbwqh/CeZFFl60mJWKdk2nHgUfouZF+Rql9uUt0kJrS
HnjbuTMEN0drs0IY8I07rc2PJhJ1GwwrgqHPRn4gbiNoBgurOov2jvXUpGNDylQZ
toC6s8GE3r1V/qqjZva73ufpQLORv6Gwv3TVpHazbTfOkH2S0fher9nB03FElVP4
4egR9TY57EKZaBAahr7RhSg7fa5QoClge5HPWUzYmmUYWFa7oL4Q9p0VCgAnAdVL
LUN9ccG+mLx7qz1fZH/FgDovjwYkyDOpIc38dFL2Wnd0go87qibycv+4D0/aq5OP
rLJdjdAXOkN6geDuz19RxbQPAegF/x3z4ggbIFN51cwTRjUXSN+4wqBDAal7xbtf
JdJZV0NOrCz4tpi436Jn3sma1dY6JQbLsgU2uEmbDSw8GDjalRutp5jMhxdb6uLy
YzqFbPr3gl4kyQw/NXzL6LrQMTk8dB7LfCcUe52M55F5PKbcSqRqJy6iLh6UQihV
JaC++JSz7yB4llcp74hJDbqSqrNZBXn0vsG+MY0Vb5uu0767YsQAqkCcU1+qATXv
OQGvrtr10gjlAV6WYt2G8cex3zRnV54OQPWD2H2tiGZalrq2rnKS/OrYL6bo8U8r
D5lZOLgEwAx+/ONl8cmlIqmW7qiTwRkXEFS29ESEgeksjN/8j39+AoeuVAMn/uVD
0fiwogi8u9T2INmFn1xTfsNHd3aq/A1P1A+Nw96wE1NrtvyI6DK6u34sIb69TIex
mBAp0hmo7lwJzcM81fgQpoNv+f2dl1wRoyTKp7Anc5qFOwXrVQINPFkgz8AkFYQZ
/s1iF+VAbNYGm7vEbyYEhasEX2Hih1ovOFUyEEpNYrgo0oYmdi4/z7abPrOzaymD
nVRmTeO2fqg689NoskE1MgYgQRm72kw1kPfBOrFXUqhE/WkTjsHEXAeYyeuYxGo+
Ot/Uc2vgXjDpXGbSnkScXHQA6Y8YrN+LH0yStczDoxPt0llt+lwfX39+p8ziQKjr
ZXeOFcNUnx5Yb1qpxAf9V83hLdASA2un6SDLOG8pHSCFV57nONW2Szu4EFsTN+q1
OWQUyTClJdaes5DXrjNlxuu+MRdpLAzUm9NNwzczBtOtPNm+CbG7inzpWq1gPAhQ
ZIzh8RpWoP1z+jSwpMqVdfqi6Z9Vp9EwAekGLgSJfNEwZImgESgYy+cRwWVeQMHa
iW4IGNAnN9g0A1SvXWH4u6uYt8a62PjwqrndPPXZ8Ci+ge7D5ncipAEb47N1HqtR
9yit3fAJmwmBzW81zDqhpxXY9l4cvV0O58ayxgkbhkOwDcVg3tLzrxjqOdwPHXpg
BJJtvpoUc3mKTDpZPJWIlJhBNK00qA1wrKZ+Ntw6Tg736gim+XaIT/XossEuNS9a
JSpAot6+EX5/0yKMzMvOGySVhDhyCcPWfl0sugoawzrYiPbbofp8S/77cV/yvlvn
+ywHLO4uJDf2MEPYUwSgUix2tLrQx2oah7BiKXyR2xHeZDtWqhxNBSRnIgiupjAY
0PBEHT17c2URqhKi+lQIWMPaqq/WCasw6Dw4l3sPYgL4XwDx0VsABN9XlcG74eF5
ZoDLa/lYXt2DEWg5zaQQjtHd3vGbBYfqncZAlgurZsaY6hpWmewWr6NCO+XtOb0q
mJcaBv50ITirO/br/5sVeNmAguT+QnWAH0MjS5wbmzk3KRVjDkqqyb1NFf7TBUBY
ezfjJH4lv3eNExZP8l6EX3M7DpZ3358jexSq7V60WBqGmvSgO2o/h4glN9DzZjAW
rlM9n3HrgWP6m6MzZuBTc+xAkQpdLx7B9mb0GGmfw/495h7thq1FC4vifafAC0pO
BLSnV97x6QibnAYsEltLLr1Px0XtWdGas+RdYkGMj61UKzKKbdJSc/j2ag3xpQSh
ETjvocfoaB1yJH0O0R8vKoT8taxVj547dQRwOdU0dMQ3ihVhPeSE+g/jXvgG8GHZ
ECNvm+IbEnY+A6hSTWDhRoK9QjqIObII+OrvO66goj4BytAe1U3zVc2tW1fb8RTs
ZZxLZLK5H37pgH8bMoVkl5v4r4OzG8NP989lB7uMGFTHkudkAoUUyrlwG8cE7XcA
T8p1oyxzV/IBuUeWGx3D7ikiKhCH0CWxthwJREaVQgQYLAnEuXBLxYhpWuV7wiZ1
sn3j6DT1RimSopz7Gpi598D2PXPAczBQxkqu6bw28gtlPshcRjs7MCtleoqz829U
1RFdFfRWT5/Yihi1m9QF2y0t1WvI2GSyDqLuVlwDZ1jTP7KTCout5NnMpiH0mEtV
mzf0WbTXDlEsWB6/LAKGG7hcvY4/nPQJr/mD5tkLSwM/dpWC5377iBxrnR19wkza
1ZrAJmwTdWlk5EC9q4I5Zy8UQP7g5UE8RwQLj0elPDqg8O+LuUs1JD6Q7aXIgIvy
VuiJAZYazGoHiXnnQqV5iYaj4ORteFH8IjeEVEQqMIhHknPIXCNDrpuR4sya0Q9t
oGydgWzw3P4l2CaPMQt3aUrKYBak8g4xp3YGpNFvJhDvlqDQ0MS7dqe8D17f1GYX
oXsUjxrtuMN6eBHiU0h+Y5ZPgXGsXUSy03MlMEHhmdM17c4JFVgjTX5ieLJykGIi
3n61JKyl1Z9Efs7LisqPxzGvfYIv9e+374cgvhva9Z4QpRSe4PgWzWUv+bZ4MCT6
DzVK+8IVfVEP9LD4h9hkoxY3uMZeqwPmz6kI08i2UDRRrc2LxtA6RuvVaklW64Mq
duyPJ5iTIsllMBMiZxhxgvbmg7ds8uI37MVTAUJQ9s1VUjWNbPb+kYPzoVnOQXPq
gi4UJobmTCCrWJ8X1TL9zvBPTu8bSA372Bgj+ijEMgBtET83F3nbtoRZ/S+4NmI1
UFL6ECpNT92TIwZ5vwk+0+YRZkN9TbJythQhTob04CCZmzkiJUnttj5hQTmRWg6W
Px+r+f6n9tf9Y6ut1lFCrTp3saYmjVt/mllhBt5ZR3cDyHAz2o1mRspFGWUDXGJO
2ilds6CKf7ncmwO6dbMsn+RufcOKNA4ynkSELh2jYfMemvZi5sZ2i5SNMmu5er2C
ogvBdT6faSTBKLTOaWwFh5tjfGBRhsv3R2sIEAISJbiqkRIQqGs1GI5tAv/LnnE6
Qo/Vt/dS/LUat6Ten32xmu60s8b1i6OSHvtMITi3X2l8u/P0Y/5DNdlMjXM7OIU2
ZYPERRbIqZjwRDzgNTvvvCN23BFaIAY+htmko8TXimkVJtA7wO+OAgBBmZC2bDky
F8zf98AXN3DuXpQrldwjBnMKfXDo7d5CAnuF+k64/Ta+mXV9jsAiQP0fpQHvAvWd
ZJRjgamGS/OX3sxW/yVl19LSUip5QmXPeaVOtwmXovmKk5vS2W6Hh/GVXcnom277
7EUZGV9Y/DKlEZd+GP86pbxulB/zB0spgahqiEaHxhIUqmPie0RbFY82GA7AP8pP
Gy7ByqhJUL7L3ObWoHck+TrxIun+Ehxc/IE2WzEalhWUrhzHjs8622SqcKpiSlO6
8hMGe//bH3l0S3fsJ2I5esQ9J4HXZBJET2CxZm6grhVHHxWrOm03CZ4EMV7wB70K
88vs1jWS5KXG+if6AP+eCYcHbIwwROIT3iEbaBL+nihchkb8YDhWCj8y90rBVALI
titn4WEGy1EqpXTVVodlYjWumemnDzzfUtAZSXLQGLEHl0GIGmWMrdzaLHaoJNUz
tbKMCYwezAe9eGsXxqx2QsToiX1qoMYOEPSwxaoiN7mCIxD7t04RpnR2DLkjgjGj
fr+c8fLYc2xRfdqsoK6mUyIXnTuqJJ1pnWfTWkxAQeGjyJmG8N2eeqSIxsAHcnql
vSt3h3YzyCMl8CE3PTQ3HlA+R13gDqvLoLsPPfPltZfg30aW53Jf2nSre9jZ1lgt
yDttKAe4/SIt4GcKmArPkowxLG7DvIKODbjVI3YN5LB7d2X1AwtCxaCSLS8w88/B
/Fi+nGhy3Rhj/Q4736b7EalS5ef86yeElcIK68yQygcMIKyWd9ry47i9wF0NOhkO
Z6tOZ67YrgM+Uy/UnN9g1n/BqPt+b6K+t2enf0sc+CF/ANBX03Sx1eeyWnwgQmYz
RGX+43kqXZ6V1KeOqLpwOzJWydc3QxHClimCygElAS7H/CYrUaYnRdHuuIOSK7l6
fGV77YS7j4XHwZ46h09oiN2ocDoLrJ0cigBuFluuTXDultItqhO1Fr0nUOHhBQks
F5So3AemGUsS2/5Csk9KSJID+n2g+H/oyEaq9cFTHUjG03nFoc02+4kCEBiNd2I+
U64ursuzidDT5kWVnRvIp3BpH2lgVLdFZgHBXJuHTOEn6/I9DgiZo7OvYLRDBfn7
5y2+6x/gp1UeFA+YheQ0WyJgcDDHmsk7mHSJpX09pWc7PaQQO89/r+xLNduyRTTr
8UgdNtbPSQmDII3nzKL4XSOyji/fBUYWwAZ1m4lGyAYDmoCR8UQVbNfuazJx+gE1
EL4o+RaaWa/f0zl3EugIjsbdxLJe+h4No+3pnWNFSbSeI8+gkcjNILGcjdTcKzYr
W6HZWkFTsj9PWVF9xytrnP9HefhAGcKjApJEoJGU85a+Oo8TOMrhWWRMYrm5LEZQ
HRfFl1esDUGlGIH/OQmI8KViubOeMp66bvBC5UxvjexuZwIMTbC08xRyDbj174Ks
rzb/mVJTDYhVwI0DUXEIJ95XWS6kUEWeT3CLtdWb1fUF2agKtjf8taJ4EezVcQhK
wz88dd5ceWCsSfWWj3RcPTYNEkOfszRITJSoA77iPLFUK8Ayj5weNj6WRrftvJ6S
fcFREPjGpEY/ZvwYLleuTBHZBhqTQY+wD2Hq9GcI5a0inb5y4trrJHnjSkawMq/5
UD+KMERLyXr+ASmX9hFeTjyvp8JVLlcooOyJdTbkN+fwV7fogF5zl4MeyQq/KVi5
tGYG6tKnX/pu7NmD5HftsZQ6RK+friCsm8t9xFoR4wgvGUHCu1x3lATBRutQTvBP
MVJwx4s/TDBtW9deBDQN3f/FhxGDdu2b6ObhXcuyIM1Sp29nFRWH5mFrKkxStvVz
AnjV5aVJlhcPQU60FKYsvXzo4lIx3ypIQsL5yOoorUK3wLjZK+YtceBMrXTwnrpT
zfevr9LFDcG8Y9Cpt8NA2Km35JO2IyzCaHI5ThYvg/UaJHNZlLckUAjJ3b3yiwlj
M5ZdtWPQSDhvwOwTpVdZVj9R5S3e2jZwsVtRdE9spsddg4161jCdKnTudwcmYzkL
/m8tUaO2h0+mUEbiQN3Vg4+AEO2yQNO1v2G1tqzySXILMOQw5JTFuaDyPKUcZ3il
GDOWsEqSqxYL8bqg2h+V0UcYxDWAemquTMCXOrKrGmD5D+ZIqK5WfP9Uv59kVOTI
a2uTzadqnuqKA+aG/fHzjU0vu48wNL5WaDO/3WfokqqJcLqQKXXQIStdp/wae3mJ
dB8sGVCqPy/fxDpLR8S7cDpucqRDBOhSb5xHpX2doa+TPBNjxjL1zttcJv3a12QL
RPdTezvOnNyuIgaflbqoSd9OqWa71upsNjZkSX+1PLu86eR7vOiHceaw4tE0bMMc
C000V3TPA7syawujAsjk6vcebpLDMSkK2jfp/jvtp40N1XRKMjHk+sX4OXE0ssU9
pvVxqycRr+qKfFrkmFwLjkg4G7B/L2Wn4Q4F/H6bZUH7unTe0yCK8SpiDZv8e6DU
0U0iMOwuG0QCwQbfXwpA2dgF3/AgH/pWMyUjb85D1TCQl1UHFpyTiUFU/0bnTfwk
G4YdQVIdC/yQLa5lsq/T3P3vw++bZte7YL9XiiFyGUwtA5Dwm32klz80R0Z5kaY7
2ZpJQPJr/FS8/dILuj9QK0g7daEPv1kOrutGd4Dla/ZI+PGBTiBwZWP/uF4CDIf0
9ugiu2W3QXBU0gPZfzgrF1ZkJB55VP4WSpyHkwEcfoeDv05wTPLnP3lphH/s4/+l
xq7B58Dy1cJ+AAdn6ppWUepgw9QTAgJyppwJnSXGOY7IEPUFok4jRgv1Xa4m2gTk
j8tmEDCCFdibspxYp3oQATBL05Bv/FQrldonpM24HSjnJevXbzLJnrOBDsQSx0QS
68SEx/zjIeoP+AXAzXCsEe8TIkuivTiR5iWPJ/FaZ7swfyv5eedJkiRSzSSyyjUd
OMZoqngGowIGXimhpril4ks9SNiZhx8Cxk8JpsG9JdJXA3+uNH0Zkbhk9tcVPYty
XhCWewcojU3U7WWhwNFJVAATZaXC9IZ5EAiLa0E7/iXOI4OmbL75O9fpdghkqWl3
rDEzXxUfN6pmIVBqX0CtDS2JvroMBwF/aEdMTiiC/jn1YZp02/GICHXBF3Ya570F
EuGFDPb7SrF8Hy1RoBmR81+U/FRYJRLyDHLzeSMmv4PKQsCxXgyfeVXuRFdxplJk
fq0PNBt18wCEjScgzHhlAwXz8X4GoMzUOELsNisP33MH8xteK4vtCX/BxiTLr/qq
IgeUmUVoRzhfYjCSmp8L3WfLEPueYHnE3A4jDu5nwaIwUIOcVamAr046cZykR416
3Iwgtw/vk4zzKI/3za4UuL1ebW9uDfJf3Q0/oewKdLoamZ5IL010nftWNAlQnjoY
FjyYNDqBsHZJnbdT1a1I6bZ9IVA0Fc5Qm8UL1HvuM7w55KLFmXXXAxO6ss8OpuiQ
9nD2/w8J+lGTI4Fuwoll5uo+zoPgCiTfiasLOTAzenHBdOAoqzzmRw+TZx3Wtt6g
cO574PF8dLvTr9+oSqUGpUZFcUu71BmM9S6zR8YZCM6bC84YmZlTST/ppZccEFSi
TkBRaaNib+5QfgNx0tNDxlYv58wxGBPs8a1c2J+487TX6qx1ViSm62B+3sgEuwFK
w+Mlx1W3Errhnr3yBznF3QrO7cfOaiwzDfyQ0h0sjDU5hS00MEZJboEKjuhhvnva
uEVWY1HWL4uYwrzs3gwiVfnT3fxuPlzxqSJVvMVUaBcGuHgbmMQklC+zokuysOOP
xBNjbna4bR/I3ImtkyTvHW2eYJexP2xVLl976VKZ7DBtfYAOONniSoLOPUBkyvT6
k2ElmMA75dAuDUBbbz5n82MILbTXu7wOdHUn9M/kx13f4+F93qqDB7zA1YPPJDba
q5WAFvvh1oPa4l2DK/QrhCSosvLzCiVukSV+USShhg09hJXARsAhJdu7iHKT1LQo
3pm1RjKzNyXpyekmTVhr/8E9QxdewL3otozJmWc3Hmy4+/lCqb2gVuaRy1WuxmQD
yTp278LwAZ/sI7ScZlHreCokjaXccJhq80EGKNQbHMQwn7c5zVzkoN2zkmVwrxjh
TxWa6cBM8glJSK80osH0R/ectozDfGXvDrNWXqbg82FQDmtz02Phm3YDoa7nAaWJ
Xj+hD9wo9bGhPNh9RdoGSvp1rRele7KtxK5oBOSQPxEc6PGYF70tFYct3h+lwS+/
PtMf2wCojukgrApDTJCACE7gJF2ZiVikb/IhZ2cV3/qXZgqglBL6H5zpGmhLvyaI
/f5XnAaRggeH7SBQpYHX0s1IdAvk4YwqVWgbefUOmmbUS8sLlD5eOifCz8ca6zof
yJzwKC66Mn9eSFZh7wEZboDFy4cbS2YcIEheAqAuFnSjOIgZLCLvLUAaJjqwTCy/
au2gnKt5CmVYfcN2Ub9bddEtJMU9q9tOj2dYQbI9oSsR0QWtZuDvn8HDfFGpt7kO
Q3mMD7psxgn8K64JSxFki9f/xiN4Fq4QQygtyqtdcq0n9jrpgPUreY1RVn2ZoJ/D
HJSJsKUAfW5kinoTJEHMNqKN3hUFdH6EvD1Jsny/Yg7uOHgSGOdBTbO7R09xqNaz
UkgtkXyoyF8F6M1yT/t52x7/e+j/grB3qel6ajkgUEQ5XGFDvulFTdN2sdyu3e2S
CU60+V5+5Qk3BkF0X233ApKllMxrc8TdyGP3xuzH+z+jiYHeNGWwV/FhNTDw5o6i
V2LMqNH65y6n57XHrvXfM5ykv10jNEktg0uXM9V+s99XO0/NPlss+N3zWVecJHWv
bmBv0Ap3MFoUKDfS7his0lmTa75YTT0H8yMRMQ4I9S7H1VJv4g1Ma3fx1FkH+P0o
iGcxouI4VGRRBqAU3KL+O4ypptbA8SXIN9glD5XOmUqhmLOb7dSk1qjGoxcDmAbU
D/CpHDQ7kzUVANgMEVaecupZomGC1Uy/+ucYgOT7O4khG6mVgW++KnWfqmIyXyDL
VBMNxJhcw0U7lKc6tdXn2GS+0nJ/6JV74YRYoAtpaBj8rTnwyaBvE9oAsIbP5Qip
4drHqAc7Z8pEzmaxQBQqMNcVG9s3B6qiwpNv2wwUd3w1KW9o0gZy0XS/Pl5Lu8R4
SHQ4U6ZfvJiyOfTzQpzbS6+Xncyoqec+nVLfeXFUnP2qGw61jDpgt5v/L2IYVTiy
9bQODHmwBTQCwchONuvL9rNyq1/LSrzRoN43CjIptgCvRwM5zp72KbB8vREDxDPH
QJKp6pcafZBldN4AOuPj1MFsUd/Y4o35jhdq9iEDLfbKPRnUK9C57o03RIyRPwiG
Q6dzgFOIa9sNZLATWkkGl8SOtpVYJJ0yzDRr7XH8JnqMhloJuJsqnSc82SVw/fvO
4xNWcHifLHvaMnlIqRsX/zG9M06IhlpovDKKvAdMQHW0ZrWcDQxWJpRnbDy0urS2
ofk7FqUs9KIcHvI+579F1250qdkn1Jb7sJBM5XI3uF+wIc8BTTjUC8E/MhLanqqH
HSCqZm2NkDCTMFA6RzQSOYeKqYkRRrHQOaUY4CulLxlXRQaWL1h4/K7aSWVrZU2v
a7oy28JOr2TeSgw6z7NqhJnmsv7gzMgpgYdPU9AUitNlWQdRJFm4R9dEaz64Kc9f
+RcfVzaFvJ8OOSX8Ro4GHCgYkLI+y3PmYljabJDeCVHg1pJXxSiI0chL8lExTig/
bjNELdv9Z4x+BGx2h8srcdF+O027VP3JkzB4QlFBqpzv6bqKHWFfCC2JrsjeevD/
L2eDBwIOTa8bEMAOiAaumMLlzuabMwnNhfaTaW+Ac2PNZ7GI/l8hbLEtz8CqMEHq
MuQ68xeI+gcRy1x0oXiBD8jMlzjKQtWjfr4c9Lp0U/fJsSrgQ2NhsljUX/+IMu7Q
bmWJ9qnlakv46v9rCJpQiv1JfMoB3RmIwUKIC+46bptXV/FGW4uW7q3ofCrABdAv
U41CVKZRVZTIfLEPbNcle9LO2HysSb3wJE8SpW0NPepmJOHBnOiUrKi5dC6sUNmf
w4OwxNaUSQOV65kkM5Vrg9ojk/kLWWWoNAH92lQbEYavx7TfDbmgmwHjVeh9I3E8
f5hjsqeNvNLANYQcPz0JwfF5oKX65N+SIJOlMfoqOzOvDk1hV57uu5bDCicHrmMB
SNx4WnL8Uuv8L/f19SRKjTBcww64EFneiNsP0uNbTmjLv+aenTx+UxYnx3ucPiEZ
7Sso2yy/C3TK/jqXCAAEDCxtDuYnHzzMN/K+ZvDUVgesO7yqI4RDWDbatU9hVRCs
GrpZlIU3f6z5HJk7Jbn9UOr3vNdXNYzei/LEsqmxo3qx2+WObF97yPRql8ZeKWR3
8e8tF8NU7xN9ZBNzP5yaTAdkwXPLmr4bo+z3X0D2Gq+LB+nAuLvq/fkkdK3rmTyb
WfwoaRWzd3yuG1u6dSv6mDIkE0jDYlJVdZicpIdoyeXxz9Qohh9qT+NqxFpeNOp0
niD/Vp171/fbQxHe/sNqu+hSHe7dednhol22HR03E4diUVPRXl0AnSzx0IzzPxtA
nTrHHCvwaoiqfdWDWVmh2RV1ARPS8Kj5TC9gaWS8Fsrg2XlnYuZ2qmkdCSDCSmyp
UT/CZr6uw8jwl0pNPXvXt/lceIesDeb5vj1AK8YWeLMtix4o2lgIAbXTKoBWrs0e
HthAEvSV4hcrfTLsHLYagHMN+YMCaFJ1t1bwEx64mEJyU7sNfPdR3eA2k1BTplCY
QjsgupeJ7BKg3AzzCDytkspQL1jYNbM6gqnqh1NK/INRx+EW1zihmfGWMZloAwTQ
lfwQd8/0oaIL83v12NI60oDFCOX2xukcal78PycY6dE+jy5w5cjIptSrR+CEglow
`pragma protect end_protected

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new configuration instance, passing the appropriate
   * argument values to the parent class.
   *
   * @param name Instance name of the configuration
   */
  extern function new (string name = "svt_axi_port_configuration", AXI_MASTER_IF master_if=null, AXI_SLAVE_IF slave_if=null, AXI_PORT_STREAM_IF port_stream_if=null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new configuration instance, passing the appropriate
   * argument values to the parent class.
   *
   * @param name Instance name of the configuration
   */
  extern function new (string name = "svt_axi_port_configuration", AXI_MASTER_IF master_if=null, AXI_SLAVE_IF slave_if=null, AXI_PORT_STREAM_IF port_stream_if=null);
`else
`svt_vmm_data_new(svt_axi_port_configuration)
  extern function new (vmm_log log = null,AXI_MASTER_IF master_if=null, AXI_SLAVE_IF slave_if=null, AXI_PORT_STREAM_IF port_stream_if=null);
`endif

  // ***************************************************************************
  //   SVT shorthand macros
  // ***************************************************************************
 `svt_data_member_begin(svt_axi_port_configuration)
       `svt_field_object(                      sys_cfg                             ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
    `svt_field_array_object(slave_addr_ranges       ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(dest_addr_mappers,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(source_addr_mappers,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_string(source_requester_name, `SVT_ALL_ON|`SVT_NOCOPY)
    `svt_field_queue_enum(svt_amba_addr_mapper::path_cov_dest_names_enum,path_cov_slave_names,`SVT_ALL_ON)
 `svt_data_member_end(svt_axi_port_configuration)

 
                
  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

  /**
   * Assigns a master interface to this configuration.
   *
   * @param master_if Interface for the AXI Port
   */
  extern function void set_master_if(AXI_MASTER_IF master_if);

  /**
   * Assigns a slave interface to this configuration.
   *
   * @param slave_if Interface for the AXI Port
   */
  extern function void set_slave_if(AXI_SLAVE_IF slave_if);

  /**
   * Assigns a port stream interface to this configuration.
   *
   * @param port_stream_if Interface for the AXI Port stream
   */
  extern function void set_port_stream_if(AXI_PORT_STREAM_IF port_stream_if);

  /** @cond PRIVATE */
  /**
    * Updates domain related information for this port. Relates the address
    * range given by start_addr and end_addr to the domain_type in domain_item
    * This function is not expected to be used by the user. It is called
    * internally by the model when svt_axi_system_configuration::set_addr_for_domain
    * is used
    * @param domain_item The domain item corresponding to the addresses given 
    * @param start_addr  The start_addr of the address range corresponding to this domain item
    * @param end_addr    The end_addr of the address range corresponding to this domain item
    */
  extern function void update_domain(svt_axi_system_domain_item domain_item,bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr,bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr);
  /** @endcond */

  /**
    * Gets the shareability domain of the address specified.
    * Returns 1 if a shareability domain could be found, else returns 0
    * @param addr The address whose shareability domain is to be got.
    * @param domain_type The returned shareability domain type
    */
  extern function bit get_shareablity_domain_of_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,output int domain_type); 

  /**
    * Sets the address map of this slave component. This method can be called
    * multiple times to set multiple address ranges for a slave.
    * This method must be used only if svt_axi_system_env and svt_axi_system_configuration are not used
    * Typically used in an environment where only one slave VIP is instantiated.
    * @param start_addr The start address of this address range
    * @param end_addr The end address of this address range
    */
  extern function void set_addr_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0);
  //extern function void set_addr_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH:0] addr_attribute={1'b1,{`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH{1'b0}}} );

  /**
    * Returns 1 if the given address is in the address range(s) configured for this slave.
    * This method must be used only if svt_axi_system_env and svt_axi_system_configuration are not used
    * Typically used in an environment where only one slave VIP is instantiated.
    * Note that, "addr" provided through argument should be untagged address i.e. address which doesn't
    *      have any address tag attributes appended at MSB.
    * @param addr Address
    */
  extern function bit is_slave_addr_in_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0);

  //----------------------------------------------------------------------------
  /**
   * Method to turn static config param randomization on/off as a block.
   */
  extern virtual function int static_rand_mode(bit on_off);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(uvm_object rhs);

`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the OVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(ovm_object rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);
 // ---------------------------------------------------------------------------
  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif

  //----------------------------------------------------------------------------
  // Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to);
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to);
  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode ( bit on_off);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * Does basic validation of the object contents.
    */
  extern virtual function bit do_is_valid ( bit silent = 1,int kind = RELEVANT);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern do_allocate_pattern();
  // ---------------------------------------------------------------------------
  /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort. 
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);
  // ---------------------------------------------------------------------------
  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort. 
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the AXI SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the AXI SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the AXI SVT
   * suite. This is checked against OVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the AXI SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif

  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum value for range check done do_is_valid().
   * The max value will either be the MAX macro value or parameter value if 
   * paramterized interface is used.
   */
  extern virtual function int get_max_val(string width_name = "empty");

  // ---------------------------------------------------------------------------
  /** returns total number of address attribute tags which are enabled by setting to '1' */
  extern virtual function int get_num_enabled_tagged_addr_attributes ( );

  // ---------------------------------------------------------------------------
  /** returns address prefixed with attribute tags for corresponding address region as MSB address bits */
  extern virtual function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_tagged_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_tag);

  // ---------------------------------------------------------------------------
  /** if tagged address is passed then it returns only the address part corresponding to the configured addr_width
    * removing any address tag attributes appended at the MSB bits of the input address value 
    */
  extern virtual function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_untagged_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr);

  // ---------------------------------------------------------------------------
  /** If indipendent secured and non-secured address space support is enabled then it compares two address
    * attributes and returns '1' if both are identical. Otherwise, if indipendent secured/non-secure address
    * space support is not enabled then it always returns '1'.
    */
  extern virtual function bit is_same_addr_attribute(bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attrib1,bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attrib2);

  // ---------------------------------------------------------------------------
  /** Need to enable enable_tracing and data_trace_enable */
  extern virtual function svt_pattern allocate_debug_feature_pattern();

  // ---------------------------------------------------------------------------
  /** returns ID width based on port configuration and user requirement.
    * If read and write channel ID widths are same then it just returns common 'id_width'
    * Otherwise, it returns read channel or write channel id_width if rd_wr_type is
    * set to '0' or '1' respectively.
    * If rd_wr_type is set to "-1" then by default it returns minimum of read and write
    * channel id width. If use_min_width == 0 then it return maximum of read and write
    * channel id width.
    */
  extern virtual function int get_id_width(int rd_wr_type=-1, bit use_min_width=1);
  
  /** This method returns 1 when corresponding slave port is same as path_cove_dest_names_enum  name 
    * and is_register_addr_space for particular slave port is programmed as 1
    */
  extern virtual function bit is_register_addr_space(svt_axi_system_configuration sys_cfg, svt_amba_addr_mapper::path_cov_dest_names_enum name);

  extern virtual function void set_cfg_for_rd_or_wr_only(int mode = 0);
   
  extern virtual function void set_port_name(string port_name_);
  
  extern virtual function string get_port_name();

  /** Method to wait for next negative edge of internal common clock */
  extern virtual task wait_for_negedge_clock(int mode = 0);
  
  /** This method returns axi_interface_type as ACE_LITE if svt_axi_port_configuration::is_downstream_coherent is set 
    * If not set axi_interface_type will not be changed.
    */
  extern function axi_interface_type_enum get_axi_interface_type();

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_class_factory(svt_axi_port_configuration)
`endif   

endclass

// -----------------------------------------------------------------------------

/**
Utility method definition for the svt_axi_port_configuration class

*/
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
O5S9KbOuOKm+CGUaSBd+zGqN7UgDiQ6Nvw1c/Aze9XspYx6F/6SEPyvRmwFHxrPi
kWVyfNd7GNv9NE10L6qOezNyBLDeY4cgveB6MyUK93pzgmpJEnEXYmFYAs5oq5MC
rJgSBu2Y1tSOEbd9itAZkTgtn6gTdaIFAGOEnAbb3XQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 47175     )
bQ4YtK4vwY0T97oKvqekaeiBnrkUgwKSKMQotDEqYtvT8/ATJ7HwgjUBsW8IE+/r
btQdut5djkU5TLgoh0taUAv7SCWTb9LgS9MQy+/a8Wemh0Iv7sCt1v5Hbprr9uvM
NaNTHVDQm0100qEBTBCQhT/EsNf7YSjK6ETnWlxJu2QP7Wkhyg57yX1M20x/rUIS
MrfOq/HXzeQE+rYniSBxS5Tcbt+OGyJ3VDsbmqWX5SLJK8EGzCvuX3s1RX2a8Jnv
eK6Bni8QAd9f3hhme0PzFnHTrv6myvq+lFrJjCsVpi1V4g7l1SHHR8u1QkRBuX/6
bkhloe2Uo1TGmPGtmc52DWSiAfvWDofVHfhQZtcBkqriOMEYlEH/3/p2vfSEMeDB
8oeM3MRKx6iGhA2psYMV/StouxYzbHL3UnLnyGEy1s5O2tKyK4HJNR+J0vcLTNIS
0GFQLrsnrpaGZescRAT0tAhRQpFpCH7z0WwP6XGj7ioon9zV2W824D3axDfjJoJn
HdxlIx5gfhNbMOLY3dBYEwdnzdelOapmkRGapu94MgubpPty+VyXgsc6J3yOzJ2z
k2Z1xaaTlZXJGKNVdY8yyR5yEVW1DgVTzdkBdHRZ7DekpdMH+9aP/ZaLshgkXA9E
gINsRE7gihGTxwws7tQUetpQR+nhylrUifIItXmiT77c982aDQNWnmFrFcJquz1n
zcSQ4H63tkBG/kA2YO27VCK7epVYGO1+ubqKhyhqewWqIxlbpdh5RGw/Dv4fo3y3
wiF8U//EkDhDDVru4pkQPrqSHtQi81oDNRGWJO3Vuhgb5b2ed6At+zpMOYXYkoaE
ugWk3kObG2BpL8I1EJ0zH+0BmKabjW8k3vAUKGDg3prQ2ytM5sIzkOEy3wZskbip
VVz6MXja7uzDEOABB1lu1z/l2+GxhtJNqVxoNX6VqJIZgekx5EVL968jcIOCjDeu
qgXgDnbphknfLlji3Qoo+IWCQTTjdb6b3zzq1YIZwOAOtgRRTvTQjen3j6fAP2NC
IfM2zwry5baFDKm3At16NQj8wl//Id0l0kbMax+CVGQLTAhFptQwDT6fbtXdbwl1
54b8SnKYWUIFzetnbdGUmopGw2RaeibehuPS4RqY00b7VZtshM4p/W4D83Dh/huj
r3cCED9da5KcNS+6t3GW+7EsWhWStvEG1mogDG4Y69Aea0UCxVV+UAWV8U2Xa35s
uoj4l8aKOWiiQQpJ6gIpjF38GWzVWXEtw4MsUfC0qtz/qpV8li9QIEncLbhswvQ9
029Ze+KI4lfqFlcKiZV7elOoL3PJ/mra1zzGVkSDmfe+FVCT1QdXvt6Aewu6uxNu
/I1sY0mAITKrMH26SijnLGXmdpA6ye40ebdMvixG7IOjivJWgq/B65SZx0TzjJiT
nmp+zGLpLE3Gyi1wbUh9wekcCipLdGjxbt9rvgzzKbP2rIODVcT+B8SQQKw7QR50
aRcnt9G16Gi9BN4/lD6ToHALVqb8n9JBzPFEk4NxPh3RI2+JI5Car3cRRSUfePfz
Y2fUwfjNGjExqkMmyhQqHiWRVTAoDPAfNcqcfw8ExnQatO8ETMRVb9r14P7VBczg
P6fOSyRZIlA8A2IMm1m+hoUV4Rtg/EaZK7mjyNiIXge6NqOknGNfG9NplUqZQ4cV
FLb+GZKDg9FuhyXHY25ezUlsAdg6kBZLuwYmnNRSKBjwOItqfgMdekS9C6NvPKwy
21s7g1/mmPQs7hIo2mgSH9AN7V//kFCkRSa27erv6RH6xFUKAduz8jGWI8M8IfyZ
+HF8Fznta74KA+R3w/zN2t0Ei3owOcyw0VkDoMO0PLrfs2n0+6o/AciW2EWBXEu4
QjVvTEzJ9VBVWjGD2GMv/b3pM5QhT1GleoztzKC4l/kRcFW+nS0z9xJXpChIrlQf
X+SR+zjf9ndEi0xauWMzgpdsPL1F2H0Wuda+RqZbqLi4XzfA6xen+FeEP7syBZkE
AQJbND+27oqPsy/p6ykplcsh9O7U8hPiVVUlzdcm6CGSUZJma0o7fH5xfHKuDTSg
kz8Z05lK8G+8Q1dl7d5fEkcY3FisETNIp3njiP+9z4sBdocOtg1RQuCx+XfZg72e
j1DkGX22/o0opVTgqlvXYuJrxam9V9FErDYNEheSJO12lgSU7Jxfvo4VmGxr3SLP
1nmCiJhTMQOCOl0hhrAjwDcRH5lcQMUR2wPE9Uv/x19sgnWHTVQ4mFFt7ePZmlNY
a9cwiuJYgfRZi9Wknq/JgcF1iLKvz1JLA3OT8d/Z8K+eFHuiQMJsW7EUDgZZLFh/
3v63VJoJ1qhCyKmg6NGBljbfeVEA4tKAEkQiJNGoOm8q8ONUPUI8Uh1rJYDnjJbK
/bI3UMn1jQdLmDc6KkaW4y/uj4mpkyh4zHgcG1DYMNy38rHu12e+Y+YuJ8bcRT0F
4yd+nFh0ceSIBeR4Y1o0rW9+CqdFcreqlFqUSZSTElJCf2oo9WV7FEONxxPi5Ikt
Kopy9lGtT/D07U38JoFtVniTyqOpUyjXEkcw0gkXK7UuorinlCf/vKDdBQepnbgz
ME4WRZwsItE9wwuO7DLps78LZq+AN87ddYaOHZHzMNPPtd3AeotLUCPlA4PvLBoE
YuM/KYSMXcO2c2U/Q3NR9HbJiv+sJ1HzKZiWPzhM1Nbj8WJSaoEPXNuy+8qU3yNp
W542swd3en7IrJ9ZBSzGln8BJD8wU9qVlclAGO7FTsyos7JijlJ1GTyGXKhZ5rJm
3KjYmKPoZ0BQhXFrbtKEKhr8vKGI9RfOlyGIDX90vkiKbrcRJE87RwEiBYM89fmV
FE3I+bxM3BANX16q2Q+ExaHrtu0E5XXBca0Aazsp2D/nnOwT4HEzObvs0QDtTD8P
++45pTZ/08cDBanIwh1Yq8VdOV0rAEJU5FFPFbBmtUzVPdWTdDHXtQ6TCGxBw203
p2Wv0x+klomdknRfqgosczm3CtmuR+LxKtz1+G7SdvOhdE8sSJ41cbJjwCmINRnM
8HRqOwbVBwKQu9mNQmcoHqk4tbQCr7X2C3T2HijEAHrNiKW4tyEKU03ctt1Vw187
MFLn+oZtP1xlcda2AKYtBbsPJNHZChccY1onrHu5nNZzRinEbG/gALIgdxxWVxh6
iHOMJkmI3VFivmgGEQvADCRNWLUyrAV5M9zNSsH2eZ++LfyLSA+pfiQY1+kAZP+S
l3cfw01zMhE7lb+E24CZYN79uL47I8ed3LqwFWgBdVGVv0V0m/xWArdy+EevatM+
VWIedGEYGr51TKZtohK0Qps9sP9AFWUOUdO6ZzvdcKpY48ejTFp8VGnju819std2
9SPs4pvi/o/hOlOqZkmCDOXc6hW1snkfvLTCt8dsdGS92XSMT3jRdyBLpfuy3jrM
QN5GkxzeeDTyPG2iCQ+sF9Vwoxi5dee6Hw2pw6iPz6gBTxVPoCBA8Ww4REz741nl
YSJZCbjlap4rDse9GmT9LNauovzSEcTt+yfbc2E6xckf/eI636Fik7Vj8x9tC4jk
TbW7qDZ82pt6Z2N1SoF6PpdfHLZ/zYQcE/q5wwf3IjkTZ7wJ1XS2/uPS1n+HT2sK
AYv7HluW7ssraQDrtggUxJm70OJnFkqJiWTwyx7qLTspTxHNiAVLNpMjbGf24uzE
eMO7LbkRp3/mddxv703t33D0IQkY8zTafXEMrb5szLknMNzcdbzMom9IF/Der4sZ
a+y6ywuy4lRI+cbFV5UgmBn5Ordmls8guGMxAOu9ks72YfpV9kAeZNgkBXAuMkd3
ekVl1fE+hBUcyKSp747Qbj+nHV4ccROJrP+VF0iMSK4gwfwJkR88yzedc3ZW49eW
fc/XHFpaoYZxZ6Qy0cbist3wO/JeJkKJoA5OrQikNLEnj6y329AqIb8oesVgRv3C
rmwSUfXMmb1xPZyHRbLxN0sQcOCaW3yTxDzrtaKUc9Rn8q8PdkEWt3hB0GsNGVaN
QC6sREgMoMhQQ0uUnE6vTgL12sq+pQ2t1EJh7XBGO9b/cKOUIHBkwadFpPtarXwV
x1KjGQ0ROVQjC+eKCQHhcofDwYq4efCYMGaHpJnVHwrozrpGRBGVfQVq6KhqeKPe
Kcls6r6NfGFoRkJUiGj/eWy48ce98BbuDs8O6usqiw1Zh/q4NuFxAL3NxUZXKI9m
Pq17mLVuBp/mxjduSRJjQLvOdeMmgXsvFPpJzOy2D6xEo1BrEVeKZIThmi1c+v0I
Ilj7oeXpMkRkFCa/cVUz3pi4CtyxXEJM1ADTAJ0kA4amqG1CnXl2FeqKNCxw8Fdd
P28kM/fNI0SSH1NDF6LJgx4A8CffWIBeTX4RplQ3Ll88CLN7myAgMX78yRHnJ/nu
1Ca/UIms7Cq3I1QmWiHNumEji0al1tuHKH7rNiJbRXJAOI9xSO+m2TGOqFSRo63Q
lLXeNgcvup66EeJP2KDgnq/TctM2F9SuPCLY8g9UncNTias3fJ20TgDLeWXqQaJz
yfJOXvrvWUCdhY+mqGWxQlZMIAIv8nBTd2pDAyvGUmg5Zafc9U8yoT1a8/4tZwH0
q8cyGy0vyLL6smJkPrRSxP4w+MF1hFB/El4fZQMm1nwmDRGLmV8PkHHiRqKCwP+Y
RZnLPgdB9ClKCIEaqvY+nP0Gsl38wrlTq3a3FqWOD5XOgmcB8E2RvdPvbKGkLtmK
ziESNjLrGNH/bbpegk3hjTicsXNMCWCwakx20FLhG/91erpZZVrRYAQrbw5/ykKc
kOYUq2y3wATGO/ujU6+HpN97diu0aAn7H21R0nvQlQLETzx9H8FmNDRSdKzI8o9d
BohIaRtfV4Li49vyU4t4HjKBzBWR5gLjq5xHUCqWResxBI6IfqolPT+EHLhtiDpl
`pragma protect end_protected

// -----------------------------------------------------------------------------
`ifdef SVT_ACE5_ENABLE
function bit svt_axi_port_configuration::is_bcomp_response_valid();
   if(bcomp_signal_enable ==1)
     is_bcomp_response_valid =1;
   else
     is_bcomp_response_valid =0;  
endfunction
`endif
// ----------------------------------------------------------------------------

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
eIumUaiaMDaynAZ8JyBUlMNc8fkN4lr5JchFFCqDlkrGDZ7TfEXRcgYTwTjjE6f2
Z7JfNYOJIZq0FfRGEswEaqF/spZJVNJdx/zd+Bg2b3pQlGFMvbqNam+8TyuIX/Sq
iZPEI5MLmqYqebPDZVs4fC8TjgxzQ0ZSGo1BYiAD24I=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 394644    )
nVqrnCY4PSO6hKqViOkNvWhAGxW97B4pFDYp5NT/8YZCMIw8MulYQQh1BhhmJlVO
/bnwik8k7x2V2/mU1B1uFihdHYzMxbLC6I98pPvEDMni1/TZxakI0+JBtnpLWYEf
SgUxvK/fQAkAC8cjCN1+kxfr1XZiQWF9TtBwhYn9O/1O5DRE7h2e1YXIKdSeSQCp
S1PbAsSP5uxTGcFOYvH2uRr9ngQ5sQEUtX8u45JHXgLJlIch0y5vi8K/aD0Rafcy
SMT5T+07Tzg0lAdvqSJ99U/NH6FGrpROV9H84bGnq2y89jykTxlWrj0+mI+XpvFc
YL7EIfl56oKXD7dCvVtxkR0YyBDGxBWPqF4BKKI+543PVd8T2rXM1yTrk20eAz5V
eQA9ajxo/l2sMkREjWvH1Sg75XBTO0DzzEG7W/20N/v8jJt9EDmQOqBEzJ4WDG4a
fxSX7FnI1iCh03ksbCuVYM/b1W8ugqB9TVGJblsP6xF9YXATaXPlKoMpyGoi8S9N
8eZbWBTpL2upfqF2VZplG2XgbGD4AD3c1wVyB2ylbmETQflgeWZ/TQ0g1+0Be3LH
CSqdpGroayZkAZpUGSPoC2Xr/sNiHNe/pIQahlZmT0qo737/ZMDsQ97r13Lve++h
0SgJzQWv0RF75fEuhWbb01q8+Yx0l+ktbMjsu2P9O+AYcNRZUi8kAEgxOAkqxfmB
Ctz0eyYQaHWRpK0f6E26JnUHbMV4dmaPWVQo6VTLtIx+ap4RBgTZW8FHjfeZhyaa
gvyRP0e3dA8L3sGM/fUnWSXtKf1l+kYsc5/xJrZEFbRZYOoj5XRP9YtZnyHT8dgH
TR9Pkf0hEKBBfJVciC463CcxmDRiAYk1MqxgELE8RZEnP7qPHEDfzZpx3VOlMFib
nun+SZVI5a3a3Ee5bx0YBKH5vUM3P6a+O6LgZuZzsKCel9QhCG5HZizpVtu/SJCs
cPXK2OgPMjnmbWtIbeNXQxfC2/E/6UmkzHERT0xb596klTw5kWzMp2RZTvDEsTYw
3r2mBdnzqesYjk6c9tX7mt2pyM22ohUGchkFyBif+qr1WZTnJ/cxoei7aiAfaG3w
96erLz1PqwDuCBOdoIFYu+hLXLw6Lp8kanaJdh38CflJUfjHsowizCZKNRiqrbsw
Xmrfv6jjgpptS0WIhN+hJo/QP9kYJJagxidvdqR6eo73XLtUmqbL5kQ0JdZuLoie
gb4U7m94z9Az+In+sk3PJ0WrezmTIEVLqmRT8Ul5EDpb/V+gZiIYsM84x0rXpu/B
d/Q9R9oE4CdxcBWUYySoE53LBvlH31D0c1g7czMoBKCAej0dbubNnjLDzB3PTGep
b3chfcPx6yeVL8FPDCJ5JzDwgQAQyAws3p8yraQOgd/+qg+EXH+uHfaKgveh17Re
G0UY+G91UKOjPWLAxu3gyjGbNgWpyUppo3Ad1yDn/wvcEychFKfSz0sSkfNYQGoq
jCTJavlcOAIWJIOhkWi+HsHKo/c8I5++/+tSBMfRXf3Fx/5shERhJf6oTwIjhNVR
BqAhMjseGHGPwvHudQSk9fjPTg3DSpJH8wv288TPB71/VeaMsnkNfXX2K3flUX/C
0U5KC9S7pC6u7Oc+4eCNVqr6wh7B6TWV3dVSKt08gZmVJYJHVAS/cxjcTHPgcECZ
u9jze+iOvxN/30cSFvXVvf7RbBz6BlThgUOnOTMFlVTe12elAyrbphoBJy8WSR2J
w5iaZhspOPRK51joDLRLUM46ziq9VgEwoiD4Nyt4L2roDaBhX2KbZ9ErCKN7enki
auzx909J/+65214gYdRSlVmAT45ucgzEj0vvtgxkLYBoIjolAH1emwuPLH8e0j78
oa3MUCgE7vvpYCnRHJ9cXqwFo/PR9Qv90dHIsUm2kxzqQnWUzaShkMPG0gth0/tp
bpOd/Ga4GSqdWL1MRxiMeN7sh2kBmkcgAQcqcvn2hefIl9J8XWbUJMKmIZ9RF3SU
UnqqmGOmUZE2woDGncmWko0zrLxKHy0yTeBuz8Z5arMuPzmy0DfYKe3VvQIbvACZ
/IvLfuVvKMLt+xFdKyNj+ECrLh5u4iuzRMM5UrzWmHWMoP3yAPNhQ4eKNkZQEkvF
QvFUlNwdL6615L9wt+TMd0PCllhM9/rtfhcBayFvak4KRvmThDvc9MbH2hdOce5g
y2qEKQSLX7p5pijvSC7chvUMcFc+N/FKLOV8d+MVmvJfXASczVOPkrN8NfOHIC9W
5wzYb5mrPzO5BlG/kp4kdTYgBFWf7sWcIQhTT3KXrPnhTTuv50e9kpZNGmUBEQXZ
onT6XXzCl+u3SdO9ET3hIDdMBe9RavRnmepYfexYozhUkUqdjl9xdY4SQ2/vTIRY
q6DIWfCnsWnuB5BHxlnn7l8y26gsA3ps2rAFA8VjZfMBobGVd1bQvjteHwNFUpfV
aSd4i3/YZPdt5Jw32frW3jbRNIm2nC9Xb+M9E3PRGKmsrLpL8Umb48lmuDfATGo9
muISPYAoOWCIwAea1E8kpFL+aM0fX+osFnSsMMxVKh25FSjbGlDdFYXbxNibPNL/
1l3wtQ9g39sT/+9q4CLWjg+vtatJt2gi61A+MIBOgQwSQzWPDgHwbus3L5S+GtLN
sb6USaihNzBirstLAHgs7TvYmjl35oj2Sqdf++jafn/HBLvYr/BdWrLFF5GHZmSh
/6mhdxVNL5S0SGZCvmFC9g39wjVENBvHjOO75EC0puxrg0yB6RJOR+9EI7X3i71s
Ox03Rw6eJeBcuZ8QIuR67AmVi/InlccC2zZSTxSJyw+PSSnHdMU7RnKPjrnbwENH
PDrloe909DpSTPOi77BV1yW3EBMqULYya92YVzCj0oRzXsa25P4QVQavesA0T+H8
mHnkZmRsoHrp08BR1D+96PrXjvwYmM9op/CMhVZi90U6LET9pUfF/9Zm6qleLJyW
fVdujuGailjBonhvlx/WuFEDIXhAnxHcUMZTTHp/tAimxPizDD8lsJThhCZiaX+/
B9ptLelZA/+X1c9vZKlMXHgr2A11ny8YRqlsVAFmF+1lQzs4s4IwtbDEXyy22Ne9
tpIemg8aeH3pUyx2laqhSxZPWLHbopDG28O+AyJHAc5z5nbHYFr7nwRJ0mHZv3lw
sldy2o79eY35pnxYAkcIc8yJdVt2kxuw3tfFnespx6PCeFOCwcBhPfwwEa9SYvfd
mN4hl+du99/uBXJSuUI2SZ3OdVfvgfv0u7nat0KFId8ULnVnSmiqScoD0RuZ8HzC
LfWTPDYDtXI5npRD/rjIsjNpWAvCQ1MdMHPAFhm7AS1nCN+MH64ZUqoWimP81rpe
h58Q/kqvlN22WLJPQlpDt57fsg3RSri+D2Vv92jaSoL2MIiQrc1/QBGHDURH80Ha
I1dnJCdTNvlrvxEPfSAZTsqnU3/EMAkxbFm8uwLa3ZTbuQeSRDGG3kumLPB9LsM6
ov52kMS+tKzuV7q5zJTDFdCZrbyjuw09mlCK22qYrkdJfOqtms00/CJ72CDY3uP/
YS9uuPKRJSbL8chcJY1Mhy6ePgM178Mzk7l7pJbfWshZtXxmzOL8LM6YOdR6ZiVA
vtfxQzgTtiwVF00y8R9Q3/bAKXP6bYVzyYlwod7n+5xqJRCLrTZNHa7kgCgeTuJw
Zlcu3E5/LolScKZtUbQzvSKcQDdJKWRgzFQHC5XSgV/oO4ngXmb/YQKHAGJW5YKJ
WJBiftIYK636/zRr953qW6h8O3cqXyyv1l8Jluf1TmFR/qkgKAnx5aX0f0Xh8rO5
N3MJ/mSDnbDMjQZjZzO/YTtX9PuZz+YC05C/06ynCQfsnU1VbrUSbIWIMCQcHpDJ
krcJTOXzT5tlwseyy6NJYxBbPA73Pl3rdcHRNyLhrj2AntilGUi6mDD/82ji2GCL
FAFOxEhoRThKAer31YMOFpuZOFRHZSshSAri5asz/+8erboAmjGBmeZzQj7afSHp
OC42QWMYEOebzmaBYBvjyYi1I4brgkJrGTU4fUPlDSyTaCZDxE8rbr3CcezOkSNN
D6hzCXsWv+Qy1Wj/LL519OjCU0oUEWkjEvrsq6bTmTO/DUQDknH9++K+IUflA/zr
KfIN2hrhH7qpLSGh8/i0ngtZ+1lILDgC0CfUTRcoStxkD3c+snsaPv3FpedAnUgO
qO/ekvrXUWU3ZCW5LC2wXUzUXE7KA9rqZ4RyQ6yXWx9Dv8JlTlGf0+UjauE9JjNE
58BiMPO9v++u1ztt7nNjr7PNqHirWAqFwVw24396MNOP79SxPYHZ5KP/blvx9v5j
rcFEDqGN3RLO5RN6KuM9nqJESe/lPuFoTnCpKbm8QxNo3zMX2HzrFppauJN97c6n
8O8mkoikeV5CsJahNcgZvnA1gab/hI58rMxPIuQZSBT+CFzLa+/d/4gXIXmaMbgW
8cweAFxFdVviwyeGlD041RyD7iTrUNuLgB0BWiKCwnTyTw9jR1231X91VgULuyDb
/ENdGSHtopf9Zoau/wGVyuopMaALfyw/H1yzE9Xbim48vWwKLlZpXnvh3McXV2DK
gq/AfiWCkF+AiG4b4v/aeBH0qoqU89tlNSA/HcKNNqCbmxjOfLo6OMmwkTcmfjhq
0BXfgNwOPvzmyQfbFunBzEPM9DV35dHA+g/C+qouyAv3BP1wcruDB1qIgkrCkMsA
WyX7+RWei2Otlqoe8dFUSCXhtnatDObtm+h6RBqfXC3pA6KwGFHh9kcWHecV/NOy
yllFRpUwo3Act7RBQ1W9hcOB4P6c6AbhOPySfnXOmdHlOJ5qhEM6/VZcljGU+85R
tFcrGVvCtRIkSOqant+CUrs302uxlU6iTMBPi0R/iKpwJgKOUmX2XrIHubiBdATZ
Zk8otsyjnMXJ9pHZoMiLHrcfMMqHOu1EobjPbUAH1q5cqrTnOojPzcSWTMLh8NBQ
fpACKt1MKjARjik/FgaPjSkud7kBLGkDSgzWU1hFrZQj6nNc5ZvEi4plH4ktDuBa
um8nPxCWVlRZbW5j8ZW6RNAWU5UyfAkqEzNC7zE6Rj7cz38Sp5WYgEJQujYIuoie
eliRMIjCZxPXUcpN/xgT8tOjbYph2VseqrAG2fovDaR4AB9V2BlMP6OJeCJoeu7p
fFgSU2EBWyKjDfbAMR/1D2dKmWE4xYfQpcIUtm+PtX6Nd3TkwHbPUYaEy2ztYHa2
UfBz8dQFsNzmTxl8flzu2I4X6AkbYmUnYALTYRGEKDAmV2PluLeKqo6gDNCcSuk3
Mn2NetvW0YPC6wLZPyMWSdpa8mDr68KLAMVhnaVM/2YnNXSPpDyI1k+duOmRooZi
J6TwrYfng1kBk1Wqct9f5/e5qjhmhXJkHDlPgGxVDIYR16T9zKrf9iIel1ZN4X92
b6yqa/5Uhr4wq5abcFLNKlQrt2ELcdXp4eGfkVWIbnLqutie20qKMuS5jT+ooqrD
cp3rRECPTc/WkP/JOEIOCEtJVa83EuPMYb7SKC8QRS7xUxBN+0JUncdF+Oda7W8A
0qCarjNniAjEUrGXW8fbVWEWsJz2s+DxKBO3lA2+N3zwT233Cm2IWJW78+uFXm5x
TYFStQb9P5z0PjEVRIlAw4dnatyLyvUaDTVRMtkVVVE7OmmdupxQTLYjH9wSy9zZ
gEsOiPHzGUXAwfMB+ekGcdc6kh3rZLye0LuRMAae5nTUKUPPz3ianrGE1B0uyXRc
RmCfyxvalGveN1RxmQj0BtXClRN2jROb5i3LxztubevqO1AoM936tq+XqsnJhgP4
+CrjgWDVtcWTpWM5ABr3MnZiOxgaj1OLB/lWWqXhK9dC1cBlyo2Oj+PD75LPiO4G
pNzHz1aqLK0kWGOk02+KWcaTPB/i7dQwf26Ca+gdxH5UkJ1YhfF9oDGF8GD/4J3p
PrWuHJb8knz8rDn5HRlnj3hPMd5sNQl3OoSyV7HrbzlZ5Za3EzUNrkNqP4lATD2Q
RdzYiNsKQU52XaGWf+P66I3RQtO2z68LG1iKwP4fzBG6vQKN4C5w8lLlq7/SyDu7
2Gp+ON2O9es2NEVFQRq/w+LoFWTbXsYOMY6+zIepTLX59UnJ8RI9x6aWXfstOG40
bjvNds0x6nr5DibPS1xy0rVZMQKdfCUlsR+uBwxHvPfAVBYNLFgXv7HhZwDnLGRI
xLlnkFaXfTzizrZQiwz/Oe5DamShb/XOICIHIKEuX2aaBoocxzLizQbOQs44Eati
LFZhU3C1URCOyQKgVwpxItwighIw7MHuqTVtyQLAbFriZQpi+SuXj3/68zFuDtMb
nc3HjIvCHJsQG5IVu37p0uO2M9K0QknvxoFnflYf6n93U1vmDq3HjYTbvOIBFNe0
oti7m/tbvA29FfVvZdtgiIhkQQr58ymTRtjPirQNYLXl4pLVASxG26uldr/rUwIz
ieAdRAcodpZOMbU+s4qvc8Vd8Z/wWr5/GxxpGyU0liYSOghUWBtZCIjLH1myPEMi
zPYXi8zEiY8K0GyxwWTiuf/3t2v9tL2mJdA3u90CpxJeIrordvBUvyUw1KCKGvuL
uB3xSEEdv+1oHOk7NjxWjj6N5CLlBhnwwi32hSTu3br0GbZXpV5n+Yy9VYELCzms
bF0x09OCkXaJWcxLdIUDwRa0ZVDxC/10YECnI7eaesOv0VsUBmvd/SvPx0QjRedq
MTi75LTZktTmcNiM3xlQQjc7z/5ydlHgfuC+FpMpMJcs9Gl/eLffQtz1pAa08Hgo
k5ZFvJLfOJhsJ7hDCgda96j7A/YbhESt1bUHOEs9bgatfMvrmzi8YZf8ClXo84Ik
CchdREYZbMKwpeoo5eJXw0YsXse5ZdE2ki4vLgGc+esZDziHO5sfLVh38r34j+HW
lPMOUUg3r8KZYjJYOOoxjycgBlUNUjYq0MrZLnxs3NoOGmrBqAWAUpRkmC1BB8He
I+Yo9VvGoHfI3z6nV5HdsilVsPqmNBht6uCh8WsBg0r3DT2Z3S7/Kz/mh4Zf4/xm
9f223nrgGy+Hl4LnsICk5+JGwFXMZnMJQhRRyRuwBy8+HPRQ8LkPT8fOVUJX7FlA
QB6MvH1YJ3U7FZrUtmJy2X0x5W7IpxKnyDy601GkONMZc1pOp3I3wmyRkMdaVYzJ
6jSnJtsqOsVWYfyABNWHH8SItzgpIU8zlbbQ63s25zyg7rgNf0acPw6+kshLXeK/
1GEMWs5lFTnicrwa8HhcQ0Sn3hm0POEIkdWLtCLUvp/dGqoqRH+7xMT1KsF1/XM0
3X2UDEWULvMQ2H90qU9gjNOXAkZw5WEOxQbtwriNTfAzI3bbK9NbuDd10uyUjC+q
Yx4bv9lugDFYAv1GmmUzEqCPd+M6ky9klL+kwC5WJQAUaNQZNlRRYziJVInNAqKo
30GVU8k56fInm4j59YbPXqC1EJSIZqiazIp1wAiTyzYAUscItf2VtqHQ00vQe+FK
N9wOINHqzVz0fUJWf4u0uGKd2Cd1YxLDs3Olx89WRuEid7HmETMsH2sEjZsNjJpc
e6AjvYGDZzp+1zDIWM1zYo0HTa/r+zH02RTR2nWI1CFrwGj/11DP5GpWL73Z2Pb/
rt5V5RsWeR79+Zuzf17SVQwtW9fD+73NADQuJgv3oKzrCu49Y4lZO8GoigvORU1k
ESRVpRfhUlHfM98C+jgpHYksX9xUkG45PInF3o7rXIm6phNgy2ALoO+je3TznXeR
KemSNu+5BzqhPF8neuJyBqAUL39iJqFaNcnuO9e6sOeydzJLdjmA/cPcIc0xvw0+
OG7lpifMlSoHhoiakRfi9W9/vbK3q5O1nnOvbv4GuhC0FAX7p9fk4Tda60u3GIqe
UVPrLGHZgmyWu1PWm1py9jzIenYahfk+phkMBzIGx74VwO9YRPR+7ivk87rVLIN6
Xmp24dEP/wMRBxKyx4duchXh0i4goXgkXA7UVGmdwfdGTvDegu6VjB+D2VTRwH2n
LsRmV3f3NkQ/tlPtfjCdYuLRiumAVOG4s+lUWhoIMA4IOojJhMSs+7NTPNzLpztl
RVyvlC+D5S8yu4SewyxEKf8K61mB4glm9uhE/h/C/IqF+LpcyIG0a7MYDvwhS0Xh
q2mkUyQ1tk/ncjzjuaYZbeXz5Zbsp7W5XJeJNh975UalyJa4xi8hTzeSQ2KsnxBc
+vWBQN+Kcs/E8dQIlc3RnaYcif0dIz3Bexps3BaF3aaPAIG0HN8vhOEorEHfNf0g
H89OlQqrQRBPr2NaGirEFYmGPqmF4bwaWZF/Sq4mS/44/xSMXcU/42MXsTUqRk5R
WXG/6Fd0jLo+H4Mh3qhV/SMui8/L23dUpVGrSI4Nx1bY65Y8p4i3jKXmFlta5X5Q
8FR+9fxzSwKCtc3vinQF+c1lwIU+N//Q5Zm/MeOl7jQS0vn+DIMDeHgCittoPJ2J
0GxyWa75/gGHUo2tKZ97t6zsumdy2o66lFd1n2T2eB3eSQWc5ZuFl6XMMPlxyKul
fwQRizqmpqaCVjn3TNoqPD0ZuMWWqZf72bg001JnZRMc2ccqpDVSyLOLntfs+4w+
AbWMmBG/vbZ3PNe4VXXCbu336mruMSQXr7gNLKfJ5K+goAAIRMKHQHgCiVy7NLKK
jo5fNJmPFgjGpIc7TwyLoBYyYAOp7qFBiEZTxOUUQivbdph4g1yIZhTLkOjr5nO3
gHcoaJ5kFvx09ehSeeOEGnCLA0J8jArhiVIkNcIZqNV9PbUVdJcIP7EznWJFRf8D
3R8ymjQeqlldue2jc55rMnoP3i2uSXeuAXBDHajVQdi4xjPzEAsK54XMsB0HRfrr
rMLmBn9SOv6G5YeNXxdEbIA7Hxk9LKTDl7lRr9LzyZ0a9jZ0y3XnVyCeI265/L7H
cQ7Qf+d26pXsug10KIgr8nnUWaJZsY7S06PQ3u9Bmk+KP/ETC6bN3lgUVDCpw8u5
1SPu4ERyIDWqbs9xaMPy6d5rcZ2sQhQeZ4ENBm2Aoo3ieC+MdvpIKvWD2qDj2r3W
suhCaRA2kt7/fB8eGFZybg0g0ogDaq6lfg4h2a3JulsxwotPjBHN/QO8OJR1EQIk
n5+4CqWa+N3beR5mXMUs7MSvBkpcl4qexOQjEy31aynjp9cZOZhpXvETnxTXTfj2
aEiCwFj/hSzu7mXyLv4x7y+yWAtr5mE+a1dHnDt/tf/JUCDSUtFOUXy8XN6e0lIX
nnZBHC0ysgkm6VjDJh8Cvf5TENyI/TWlyHJYMbIzq8W//jUGmEHyfmgxJRlyozVI
bSOFel34d9B5pazHYdwDNjevrUfsXGnJRKflC86hmWiif+Tu/Rx67b3iJfVSGHws
mATuuCLJkxkRbPKRTN/SAswMYwXcM9NSJE0Hp5mg5Fck1yLEy8XvnKELYWIGne4h
hFeu1Y6Xjk1TzQZt+Ev/ddFoQ1M9bYh+D5F9mXvOUMRi/cOhv6EjoJ6AsmWplAVu
cItWNoI9MysfLEsDTuUYrZmG6M1Fo/+cyNItN/THHI0nlRV5g9ciJz7cuStWOKAA
pnYAYJYmsFDyZAiGIxHMPtAgvcpEDFQxg/G7edWVc0GKtYTYE+lr39Q3D9nLr5EV
sUwX22a42j2M6eU05GKwJwR8qreEN9IBB2lGvPfGXp3HCBTGJE4weeWybEbmllEY
7gTCW3tdBm4e2JCI9MLMYyG9yrI0mCSsZ9/gyj/xwmu2tgNSbPBgiYPu615OU16a
VvgM8dnIsacMB3bdh1IAC2DbAS+8ZxURG0UvzLz64Z7ykHc34rZY+O5O+UxOh8zi
Kd6kX6lq19vLjjmFPxpi8jf4yDDlsfxeH+8o/3dW2BiAE5d30gL14Ra9jenJazaf
UWlvLJ/cwJEkm8fviEZI6bf2dsgvIGLrkW84mayB42eWcM5vmmrq0jBV50TRIjkU
xifJkiasY2X9Gm4YTNCnR0tWo9+Bp9S8UlhAxPeEeEavcG/OABG7m0hiywWxG/ZV
rgXfbJBV46RW0049RXqMDzPD9dna88M07ZRfnSDG7adZd28iD+JGX1iVQ5OOWmSr
4dTeyFPyAhzHnxsIS74z2p7DozoggMAlAPd4HfeaRsFJR43vgMulIsrh/mnTbjW6
XPSIYAqTVw1G1d+N7f+GbyZNAaNP7jsJF7Tf2HL7TmKknJIvUEp5PXj9nVYurCKA
j++RDlAskt2+qUKktWM5IvTXiDcPfkIWl22LSUswRklQYuwxj5A8rSzXfRnud9jz
6welhbz69BN73d/dBRs/9GHnLom8QQaj+NUYl07Leu2j5zaMIOPrNQSoTPfv8bH4
SLdmiAJUd9Khe5dSrkPT4+CwTl8EtRam5jtMuFe0Do7vsW19aw2+Hw7VqO4UXCdf
MVOMlpP93jGEKkRQKYGZVv9BXpHDGlvojrGWKo65bDZX+p0deYsqD1ut04SvVtRq
Mz60/ZQf2WG9cRt3BuMcwNxmuRGfKXTEQ/RDRjeLq4ucfVWMBuLC5Qt6nnJogFqI
Tw9lp8rF0TFh7oFmdfC3XYwTHeBvJYOsIVWyzcbFnD4dDOyyGaCyeETiT35vW0P9
D19MX3U20ILggIOshSaMGckawmjd1SHxcN45oydbvnLAGmwsD7tNoKpZnl6FWYZS
GNvq3V577bjjgeafSVY8RK1lUlO8ZdeNNYXH7tiWaonCx8lkIQM/ONOajV1+pM0P
jaWZOsrbntRndbY/wejbzCBosl1B6EkKGghHDqpldwyNrNFAcfq064Y+z5iHVt8I
2AqRKRh4UAfJ8zy9DNo/3b422aOHHzeum/JbxBTLCQH+V194n2LwJadltxCPfwYC
RiQyEySOfnjK6Sr9XGJ/jJtHyjZ2NxDfnjBev69mGbAErtgbMrf3qYf0gqY+14bP
uPRLIXHXu+gHcrC3J6Rh1LgZGCIlrkV+ja1L7C67KuKzH0PKG+am4cjtB1YSg5kp
XSyGJYwIsEG4jIvEVJb8gy0/p8DOpQaWZQ9Mb9FC29ajCsxsaxQ6poOqUscCQ4Vb
yKYVxjcBUm6VBzbe0pzCTsMAiM/hTPfeWSAuzwfvbmaW23Sg0u9htW8/1OP7j4EB
9G8jqTqWDWYBojRjIgeHs1/CI7tpNqyLCDe1lFGe7qSVPflaYGuR6DLjVBcDEVq1
CsATJmNsZ1vaYdIDhf0WFAgvujx0qezwyhCcekDgN5lyLD+DTNt32K1WFjYnLy5F
EiHRSjRcAByNQG3ueRhxT/KkbvOqKOHi9ucKjCxGZYvotZjGTiyE2ofOvC4/lIxX
FkosxL25bg4B9USknNRcgBdLPx5JB+zSRG6nB1ohAlQ/f8Xr4DEkoCtJQP4KxHBi
ancEFO+fEVEr0OhACVf9Z0gJIwaANMgvXn3wo0g46v0nVMEBUAxYrrb0vRlCmNvT
g2uSkNO238EdHmwSoUt2vzr+NsDfcMBD3jYUcYGxuPL1IPryblB+nRKsmI9WOX/B
C5k76bYjmAi8/K91P1qRKFxJ7GKjHiASvEAQxDR1yBY/4G9jLs2nzWGobePKoIOE
w2VHeKENIzhsglGqJI/07oHpODCX6AzxIHmLXmQ54WAVIJBP0X6/jl2lQKVrbeWq
HY+JjgkIeOXgpyvLix0mriIT5wEKdZEfzl6BB0c2Akm4TfrbOCw4l8PhgS7il070
WGxnFQCMHgDoiv/+wSwG4XMfqdAu8NFag64bLptFaS+7CcOfsmTe51M40kb23R2E
c/ndG5QTVggXvLs59V0pqW44erSXV19PVdEsp8/Wp9GLts7Oi9djyEEjKMvrkPkL
5XZaNy/lFsNLJsC9cgVGbwwcxydIIKSNzAYAJJH78mzbMJeayuWht09Nc8rdsas6
hJF2dcE5g42SUhTQ7z+KL2E6i9QKiTWalEyyAmsCaMKJppcC5x3Uk3By2y3YsngO
y0RI6za1iQCKiVgGo7wlD1DZIaIQvuoEieUgwNNLKJglGO24X0lJhiR/rPvSBPN1
F+qq692Kwb9e1pIqs4TCBWVupWeio6Ja9rdErVQ9nzcYgaxQEM1J0utVec1GePxP
bOxQd9Kh42CDjeu3LL7+QA9W7mwV/AOMACMevuTj3PrvNETAXwO2FX27Fc1Aw0e8
zN02qj//LFP4yAvn+mgHh3WqdArLBmgb5QNCXjK5JpeOROrhaNCEnCaU1wJ7zkhB
0lyE/CzIQ0TYt/krKUZ7bk1+FPuGx0orJqb1FaJ+HjaaGrjKywcPNgWeZFkH/hjE
7YpcDzhowizY+N1ord4kY70H/JJMJVwWkEfZ1IX/waf/NFDfirXD1pLsP24qbHPn
qY3/o7mDXUO119yHgBMuMNb0nP+BhgBsNIWoL7DYC00FL0VAMNEgPnpGe2gmuRzp
iGaaVHYCQ0Hg7nI1nF/WP4DOpx6rc+QuFUZfPYYdlhkPcQBrY763RBS5zFpRrtEW
nnfh4goluQs1UfLLEoHTVXD+3f33MPx7xxtZW4Ocm7jZmw7aZZ6E+SGYJ1hTbjUf
7+8yOum1+zubLox+AiXbRsWsLiegyHHKaMISsWYtIwHTVOiNij7vDoIVqLe0TLmh
tBYObVl+c+cROurK5FY3QBtLrifMbfNzWLze5GRkrjvWacNjxBosPownTk9vun0A
rvfIPH+Z8CYT3iTuXhTQMtsu8fycIuzJjkOjmcStuUUCQd/8GavZr0rT3WYGibbk
5/yAT6762LP9khSJzsz5F10D2kJxxhIQI/YB24yuEOL6sf+3lfYG9NxDgPXHE7BX
QP/1Otj1gMAH8XsQhl5j9t+H46cVo89loWJ9BBNCEC+zHgXusDEtmG6Qo/FLOUXa
qcZ7Eji0CTuUIk6vGzT5wfQBtyuA5f4/b8RsUohUulf34yda4f1kMt4r0gVoCPr3
6KgnMqAgK2Th3dEatEDYkWRttcMl5ZzoDK5UDvJStRKFt/bDMHSd0DcVQHgCh7GZ
TD4OUkVO2JBv1mKQzYR/SYTMOR2W3YHe/WBUQS/hjIVaqG8FOrez6dyJqTRSExC4
fZZNeC+LLsg20XsVh/BGGzlZJ5/08XKA3VTO7+iDJP9zhogWsSkhkcBgTunwNmyV
pkxopeFF43JeL2kTGoCHPrfqdKxO6qk//FcUt/oAXFPzCAMf34I1iI8s2bgd3CBy
OIFHlYYP+EP6V1/7KKvxcnzfLLPH/Kwnm/3Cw12IEO5j4qu5G1CDl1xAsLUlVYoh
XwSaij/+nJywj6jeqyqy97KaZoP2cmsnKIkUoD1cRG+XdisOKzocWpmOfETlK0jn
bPBI6ZHFt8DEyi8NDUXTG31hwDrqTzu1ndN4BoBX1S0933hpKOfGP7MEEPwPp5kz
49NTDvDIwcYSx/69vA3tXlHAIpB5/hj/j3TjY9VC80456y8CMq+jD80p8wQ5yAtG
JOsxu0IevG7XMhKA2zeqlpGZB+6/koEAdAP9nErJMjnPwODUX+rbT31ZhgFrJgiS
nY7k3I7Oh6vF/FeMFuvmwoPK0bf59DUxpAwurEhw4qLuqzEdZBDfFMZPU3LQued9
YSAORfLixbdqW7pQH1nzsg8qcumK8WB4/SWeT609ASPUaPjIdsEq0XFuliUJqmWB
iwQZZa+gQeo3NnrJMoY5waZNJyov7z7k+8+lhdwx7iP7L80rw8UyHoK+rFf6jt8B
+9DHjzgvDZJILnd+ZHXdSqaSzFluYnPM6/yQEex1hGAG4itIK0Mg8Jc0A1ZVxqgA
VU31jPldIOPd3WepWmOmH1AnyJgChiqsMlDoik2zbF1brov02t482JoIsYe47JkM
yk9jGpyqtai1C0vKX51ZXPHPjSYlcnAPbQ4IBA01U4QWBrL0pq/TsAvf1olfeKAl
EUkfWBOpjWLqkyBd94LzkSE7mPoFJwupz3IEGt8q6fXUxSNyhQbl875HgucTzH3p
VqYr2CIphid4vw4U1NWhNoh29LwguivZH2xnyIL6KzF84XazQPwe8IkyBHNxByAf
l07cnZkRA38Du1FD/HwwmNi7utS7GntLEH2P1K0hj62vDV4flo9makjBIjbRY61H
G9yjqT9Oox8qk6/4TFVyAgdljDwUcaAr0C6ykIx3/DpCDGvcLkl9Cj4RFniBWUmy
w5Lh9UQBOwojl098OUhohTitLUPoqtwLuSJtTnaVwFN/b8NI+gVVihknI5HRhOY3
RBAt9UQ82dOVa9KPCRYpw1UGJFEfNfmPJ3SgaAv/gjldMVn/jKNgrVtoOONDRDVc
/7DZcz+KVaUemxQHaiLIdmuFP0bigy43jbDP0frKt/miSHhOelx1ykpYQ9coyQp5
wpQSE4L8unq+LM48k3h3QBKIT+UBZE54QZnaKTE+3KN0EkAlXkDrZcKZMgC1K5V6
C1FEXxSMHzSvMKol0SpcV3m2UoFue4BNChkJFJnCUAziUhy5EAxqq3imPO/VtjwG
xxAGzOgV34lXjAs6LZU5L220/bxlnJ4qhRW4l+8jihcXPPOTqfiPmK5C3/OSdEb9
QVM2nxDHPey64j8Qd4FjkGafl9Tk5Cio8H3/3TJaD+4qogNOtvTSYjbJChIidJ7g
qpD55SQgRyl8kBDY5LeGyGsT90NwLAzL6oGVj0zgqHUqh5HAFhSaokWSOkn9BIt7
WZhSUvblAi8CaflLJISvXWXq4I3OUlz2GBdp0F1wkCPTCIpRAzqfURfehq51xwwl
OPq0UnWK/RuuBoDzacik7lkZ3SJHiqwt4NF8R6sZsPBMBVRhWjFHG1uxIUKdrU1C
XK3+fW9MequmMeKWsJx8utQTQiq0ZE1oxdlozGOR4/4ewMzb69GMcm84lJlTGYTt
t2Z4TJ24tasxXt0F48ETYXLTYvaW4UI49g9J0g58op93/cosyG1KqHu+StQ2etkC
Iyny5d/Lt7sPX5IjHHvhLlZh8LWbP/kLeaT+PNtsm07gWO9hjheKA0ifFwGXrrwT
vcnbZnd/7TIX21emiLjg0gnI4uD9icDlE/BXHPuZQMmtyO2g83LjdrjX4a2CLd8k
eMwcs+mVa+/ACnB3YVHDc4KFC8UEw8Tplrxz2RjAkkBmwzmrZ1MVBpJuHQZ6UYoV
3fy/6jb28hbZlNc5FvUEMV8C7s7PiW7y8uWy5RDlSf51vtIQtREwdm5FfKnRM66n
ZJp3WK4mt96uTQlXhrTmzrmRhUa2G8ETIuFJu7hoc3HPXqyh5ZqQDwM/+mlikeO1
Xm2ujogs2GUuaNFG8YYlWqZi25gMkvNL6e3Y1YFU6dPtmM6z+gXHpbY7v7jc+c/Q
SykH6mnteUrcEhWo6InpBdYvdKrwAWR5V3HYiw5nAle9Ul229fEfrKBOaG35csAJ
E4QJKZwA6ohZ2u3UbM4E6E3znPs4yG+P3CLiNJOGB3pBKnK6cIJnFuQHkmRZElIz
Kog+lN4JZxtVHhWJ3knG/ks97rfT6sNryBE6s+Iupk0dvCNKX4gK4O1c3Yu1oM1s
hKJIQK2kd5uhU3RFeh946Adzn8SDbfy7q7STcVl5bCUipLutNDfbPnqJIsF53pG3
CYKccSRYJgWkRaJo0gEL6HTd79e8oUwvRK9xT9E4pEKC13aRkB5ifPFA4WSnSOju
z3r8KDnAzH9DvvhGLlFsGrBLTV2E0Fnbg2LDsyXJprDKQp6rJlhhzs286iw+qhvL
M1yCFNG2+4knCT+RQZoIaisGdIolJAyuc/MGxvyyvWXXJIVPc7Ix/VSxZRoOvnC/
SSl5f9MooS5lNAaofdFRRm1lLhUBNaDCJVxjnyts5hZY93MnIWIAjN6yYsmUJPCo
f6hCJnz4s6vVP63HS0WW6igVcD+yhxaFHzCBGGEnd7jItdWVwHRiwli5FdFGh91c
Jk7RshRGzqOuvkIEuy89k3s6ObINIaF4K3HzpG0O0U1NNkp3UbQuuF1qADNbNu6u
72lXObtqDWvojVjHE+gqcD9xnZKwLhlfJHdNs7QysQTfeF3riZM2fGxq6WcEcqeX
Txd4YrrpBFx2V++4t0Vr4EOgjETiwxP/0pS6wLIwJNZn2UOirXJOPF3Klrnymy3A
Ix8QG5H7URdoK/HTVlDoKSrockJV8cVrV1OrTcEmBpS5yyxY1HV9osdeIcNaEUGh
3BzssLM8/N2xroMy/qaUVBFnSw2/BHPkssddODROp6yeCTg37AdwZkHpL2C2X2ni
N9CfOH1iE4LyNmk+4UFN9Tqde6ADbPEcEu5oaNUEdyq9nhVwOLhqF2SKhAFxVgAM
mMIdilGlz3IO+JavAkD+ZV1WaSzyr0NMgGh0q6ky/UKsGihj8nMS0YhXyE4b5ggD
UBtthef42FPbEE+4TKWePt02VlxhYaFoDLkwiHnkrhwsZ3gQM/+k9KxZH9E6qF6x
F9x4ODI1LiKRdDq/zH60K05ulH9573ZiVVlQOVE8fqfjceXCQL2gxiiEiEcad3Bo
AR3gYT0GvK8M4opEeWBCBpLvWj7qcD97mM1klmD6/i1g96wvH8YqE7AlUsqBZQAu
9zWZdhM2vEy7mnsiU4nDXApqXwC1SbsEQcMwLpnMOA6Fdf5c8EuSPCtG8py3DBL3
U5LCaJj0qD2U6+ral/agx2uczeWTUAGq1PhhfWWCTgrqxT1lQ1FiWvpNv56L/xGY
TXLN0pZtfJtIOVS3HYhx2n58f1acTtamQcAnCvk2unRw2PHvGeolWnDm/QdiPwS3
TLjDnSB+XIcahUBjshaG8em823mMLCJ3D/SOT1P8pVTxfVZDq7gNFxKMQ+Zt9mwi
IZU2SW4BNrtRdv9XAtMSPEzX1QV+M66RRj1PVvWyCmooP7cWXbR4+iau7ABVqN6B
UZx6xaMBsUP5Ai9giqvicqqpazkLalh8fVLsbe4yVcGPr4m5KEHoWHjHieVmmBHr
zTkT9kmYBnQqGjXymKPzBzM7XphPNGZHRdhFEZJFkgXpoaamlen4G6O5Rv+Pj2zm
h4aRIMqjtsFw3d2PdQZFNj18fWSgURZmbRqHA3UNVKJtrTh/T0BaiehHNbukljLo
vaxOKSDelJ8mGUYJlznxB7Xfa5tQPMxN+GQDuxQXu7eI9LDns9LBJtvd9WkKYK+p
l6xVxOICHCb9yp59VKLOap/6LFVTT+q9y/C3pLUoXnT4tXquCx3fel7zHDd7a/b3
GC/Ik8NcEVpy+TaQFWc7i1FFXIm5kHtfWIEXPIOF9ZZZ01H52uMMJOQxaSyCTrw1
Ad6xQYMN5No+SKqwPCyL6kufRZYNPMExovbvxuOQJXuAlR4KmaY+LXELhJ7d1a8/
0mAbAVGYh38wDmn1kuWYRlVGRFiCJNTcveknfOVHicoYjr50J3fn9CGQr1AETbX5
fT1WGqFLqigF0OV/0tZd0HoPuoz8eyaZ4M9WONxgOfUaewRmNx2YgLxz+G+sRfbc
XJT5OG8a92l0ZH0tnE+GPaQQJYJAfQHLuUS+/qEjkevdSVXIPYpEsmNrLegY0l3U
nEOnTAvSf6dSmWkVRIr2qzDzaZszfqfjneHZsJmvNL2S1RwZOmfxe0aXI6EMbOBb
c2hGix4uFo5xFyYTHPMw7f+Ae5Qf7rAsO/ZeA7+zxDJiztp7D4IigAAoZ/TQ06eD
EMvWvq11zAPOGIX/FZKvFpZ6rOLx97CIILJEQbheUYF4rkFVHNPm6hwDSZcZ5sQO
+FBJGF4WlAwBcJGh+u1Qb8mx/3ayy5VUfQVFM5aXQzfOrizteNxdg6kKsJ3uhET0
XJSNnsKUp4kety+9wK2BUEhiwoTEb02Os+zbRqDUsaMQ0xH5t21l1ijuadIqcNCm
LMyNP1McTdhtsa0Xo5JJdMo8WxUhwA/cSfMIFlSNFQFbpeAXm2WSFpunq7iBnr6x
g49nUI2cZw+/8U7Vu6DpmCSqkTkZsA6Tk9Wea/lxrRNOF2DtMMcEkofe+Oq0wPCZ
f3kFXWVvJ5zh6ASc+wYnO27/PDBV2Cn1+Tow8bKq9i7TYOIWIHE6aipnCYPunD1C
ziyvU6f8+9Ia/r0zAmqVtL1uMaCFHW1bISxDwzD0YnEjHSp9zMvGk/JRBUKuqlJy
fE2UGqjyrrEYlRQaBf3CMdnzhTnWJoUrEH3iEWTZyQGzefzFjAPSYgnCi71agpFL
4tIXzcSO+hJm7/uAOdYSsFNu7d5hbIqkB19bKiU1o3q4IrHm+Tcy+on67+0j41W4
d0HI3lP0iEOtDAcbWVpsVeNbt+olR0dFdwyNZ89buVTnMiFFOW45YXARCX4Frk7N
YLIa8Y+R6CMobfIbNOoiRiY65vvTAxOhe+A6WIkkiUZK/vvGspYqPvhWnTMdwBE/
tWllSBRp+9j6uCJmgkp/lE7LG2M35yqHL2OSotvIOt5ogB1+A2i4HVBHgbm+LMoG
QUfbOFqv8wUnOln6V9GS7hb3RZZOzhjYvKDJvo6xuhkfVpUm/esuVm2Kp8ryNDHI
S5Ck6w1OoG+ZYLDqScxkB31t+9XEXar4308tjXweQnYBDcczrTQIB47MO7pOJmGQ
GJWqbBG09l6dPKNHaWhjJdJRvDxbVzRvb+uQYLCJS7vF9rm+migbBviCf87h+dRB
vviJLUKfS+J7mIQWLZlEQdduCekS5Yreh5GSiRqOPGJB1ck6jnHC5/dcYVXvPfob
3+p4UVFwvcww5UeZzdb1uBWkJnbKCRTVxpcmr//lWZY7+KGNaO0l+tG7BoWc4xUc
EjsEmov88T69OMlbtiPSS8vgEqmKYAqJokE6nDLVqRZyg6DouALttP3bkIHIKD0z
WGWWXjcqSjso2psyNsBOLlYkWjp/XyMZFELtSRYoRsBAcz/MGNo7ghtzV4w2zKs/
VjD/+L20QtD+BdrGRnGWRNfgEjHiCnRkangD9+xl49BpkmSOI0gDzObi/RvYCBd7
2NiQrokaKPLqmvTFbwmFuD7XON1OmcYkb+dE28J58STFGtWcfFa0vRO3ekkDU3aU
T/bDWE0OYyCnn1Xqckjc6mKzbGSrYD4cL41l1O1fCfyQ9dGu9k9IUsWRZQ4Ofm5I
dvh26BGM8/RK7T+32pdbi1Wvyq6xI96S6IFK0OVVOJnfRSX8pMH8BIsGNdnekX1v
77OjGzsLb49szESpE0rvqU4VuTMCXItoO2Ev4FzJZ1xV2t4cb/8F+ZwJ0vsk5/jM
Q7YuO4sXPEK+rMFlDxlRuartVCbtBeFJHrZCp7Vlal0IDAGACdiNqXblIv2ZbkRI
Ak2enek7kj++dAbVpjXRycIeWJ0qGXg0AZrYaOoYmZDsNKAARuM4e1NCXYPAYQyW
3N1waUwGp0gkfRD3CUkM/HbziBNV54R6xJZseTKFXafdu3mzrSmtBphX3CeJkrtI
YDullWKv48NaHcQ4opCeb/4wgAN0pl/HeTyNBHxsjJp7jyQZWGcH6UGtHhX68Zk/
wkf73LBaj8IhnZWmvX6oUwY+fevk/7bpCz3aNYa7Qv3rfi0Af0RfL0dPyilEWzSI
q4aQSr7vr+EWULilNti21jONCIklY+UlliFZcEH8w2gKSRnlyByIdYwbmn9H5nHC
GHgBkCV5WpuvdHLwmooCVg4XuYRToHaT7Reth2+c2Ypg/a0+E+KSzlKUD/PqTqm2
a21lulTuI10z+JOGeoYBhsRhTTngUafTFKhEb/9MJvIzIxnXR2YLIjYxtfbZXwDB
g0ulE3GfCy9bhpGA+NBnz2Njas3N+3VZoPDX2/blf33/eq61qsXnyrJYcIfZt/qB
luc3MK8x+Y85e8a5obgJBLkVxQ/+6WKtoimqQNy/VdymXXTsDOxE67SAiRwleyRG
o2z+ezBYMT3sZ7oI7oyqCjBMY73AKq6R8F78ThOA06p1PunSuUsgArqozHtTYMkf
TDrDp0atO5AOoktK/kJXgb/JnCiUU4DQNzO7RpAROevokoPyWn+XLVUQyhBPWNgm
GggOWu8r+NTLCbEMrq4B27OaHEF81JzSWgD6KrtaBHvP/x0GnsOlSg/nUXngZf2S
V+lrp/iN1WbWSjonKUBqdXnhKG6l/3RoSKDNcsyHcIEmyEWEAulCVXhSeVKrNVpx
qQkNOer/aWQeb2kD8LMhGEm9v+9RsXu9+CzzgaLDopmQP+AgHETEClQ+rVIYvjFy
08nYkhHjWeerpn1GfQjACSUsvj0a7LwgISoJx7/6lpy200ZHUjBHcSXoDCLjEevw
4GpDqZTjfWIlxblTgiIO1P0y+8JMnxLTRN7K/LdMMMEfyoE8kjAVNARstDPCO7js
AHNJFW7xDT+/xw0Sw5Tiypie0ySVwzT4PNNp0peaFZAmFvXLMoyR0B+dkPuCMdY7
HZ7W4bRNyg1cJQVXiFt2k33mRGbue0j9BKf80ryLLk00e5mM6IgWNKq+kVcwjtRg
UIzvbSwji9dHjbiWU/wiRu1rLQE2jZ1PHhfAqJFhWdGAEfP5m9M4WKZU+S0dhz5Q
bPqLhZz+ZK0sS80zx3CpVo3IF/4CRHPZkRHjAD/o8Cz5syGYut3oTDjykKgs2cTm
B3MueAhzeWTpv9hJ0tEUCjmF4TEuTEmCgI4+fvh9NZgjL4GGo48r6gcnBfvoO0BS
EMcB7Ezwtyb8eSmXjG59tq7ZefPXdSw7B9i50tLUKmCGqr2zesLOjQG1Ih+9cUO+
N7BQJiNYAh/Vw8OA60gY5T2JgQWc1u4Ljenz1gCuIo8QRgUoxwnEtP/2Qj6SMfUL
ovaF96Ynw4AqifhTs9O8c2vFVyITU8o6rzYQCRYFBD1TO/Qbg6OCFNa/jYmPf/tE
RY7Qyoq0AtJHPE0Kh8iZyzTEDjsF6GXnqLsSq9h5uWiysbmiX4ssA1Esme4zPfSf
DhXmXIzTzoBN2rugZDS/D0cowquSNXvlULgUjxL2xiLcYqr2STe28m9c7IlzQ3Mr
YWHsdfRoxP4BZ4jtxyJ319Jk5oOkKmCICcgfVhOvsNRtVq7cBGhDB96eR96GOyDs
dOIcbkmXOy6Qiy0X8lH8xLAHzpUdKs64ceX4oLZ1SWwlAM+aYhAlfSA/L5cjWRGk
D24U1zQ8AFqSyOlEiJmcqNflyZ6uuGi7IpWVALBj0LqFh8GFs6Ht+12Jdh2D/sxR
oia2wG5tnI3tFvG3rhZpEmWuV+51ZGp4AlzgQjRFlcGn1SbO/zpda6n2reSX5z/I
iKvCIPDcWpuqGwhc7iHnPAG9iOqJJ7kMJpww+iLAToKZbGnQNCoStwUWZpNzYdMs
Jty0FKM6mipqNlzMZD9pUD49Uh7uHyGa8G0yfrCfkfZGeJTN/oFzsF7Sr1CFNaOK
JipNNqe+n84xLNnxU1E+Ux0O06i62NSb8wTLWgjHzfQvCgWzZRtNnQCFfmdvdlhU
IE/gs5J08zRnD2hEIhkB82u+Egl4A2ny0jrceOBpTmyD9bRmTozg/O2lJbuacYoB
aFEyVijmwEzva9I9vIfqzio9/ktfgliHPDzDp7jr5O4jv0kPB0DI8h8snmpCXeIe
rkyutPYCMJhaLII8PunaAt7AydOHR/kULpuaUaimmkCoLH4R6rEYxdwoy6I1ESwC
to0W1A1gXqtgULT0cX9r22T3/K2adxNbE95Eg3dHqsJAWeSeC89yljlfHKXbaW89
m6kcY9lmiDqoHqTz/j2yak5UAtrradeEnpYsiEk3ZugQTaq/PD3mz5Ztc5b+dbQ+
MXX1NjNBbVgfKMDqPCjYdKh7x2Kpex/f2549tU0eisvumPfisy7mEN9EQk4p0nsT
kyXcdWDTnMtyWd8VPomfGb3ZuxvQSZJ0zsgLToHaJ1httwO1S22ImAfLpfNKpFQj
nrXLm/ctPvcWxbkFDSNEkS/Zvz7xO0PHWWLilOXw1oklKNPezbcAFmYY1cUFh/uN
7Yopvln6ZOBpiFNpSEesomCewfXfQx2eSEZzo9ialxC/7TEV0byny1NwAZQZABEZ
FyhLz5ZMCoU/sX3zZNX5udCXNOZtbAdZsMJY07piEmsyN1rD+zuBf2MGK6LMRF/E
EIxmsOnFwpnJPLqd/eEtU/8t+x0nyH78ed4Fxg/1Wt/eQJb0zrLYqFIAOCAmsicr
TUdbozJ05IFCVdM/8LL5nHYPlxNr8+oLZ+9S9FxrGll3ef4F2te/pE3DcRkXbnGP
U1EfpI8j/zKylYLcOBrANteGwLrDJlz6QUyE/5VLXGZqYjJkfH3PE0p9F/4xpsPM
mnwfM4p9yhwTWTRA83obkHBzoQHSMeKkuBMK8eBWrwYnRwISPfDnyXPs+f1igsXs
QyOUo1SOzJ6BTgvJb+XPyY1R6Q4IpzcKP04dRX3CLfgWwOMK1Ca5b3oy8YSMYXto
I44a1HgYvx4XLZap23I/+GieGjq9oHJAJMRp8TIWgEvtZQHO/Lm/Jnmz3XV/aosR
47Lm8cON8Rc2e8cRLrX/pmoJFD0McJH3KisoYjtJWkblZ9KcpL6To1vLRVTV4xhR
yBFAgC7iCowb6XmRWhCD2ho8FIk4XEuebWnTLyAJyIIeXy4urIx46wGS7D7rXuvE
6jrLmmpQQQJWi3vs9HZ3RDKZ+Hw+Pe1rSPVBoEvZKTeYDwx9GHPo9a6dDiC+w9Ay
ZpZT2Q6HdqDXhmir34XWwEaEz2x977c+eOxtkWTJGQobsfE3dMch4eLKqttE2Isr
OfnFeeTg6Qs6pX/bbaAoZ7K7SR4mx4Y8A5QgIQJu6pCXWfXNuu7sK9RH20N31Hxv
X2zk4IOuJVtSrMdTLZw3RGvPIR7ziAnFuCb4aZHzVAmyva+1t3uJ91GpZR04FHjl
Wg0azrG597Rr64xLjS08omKrZre0YUpf+lT/+4yxGuqNK94Jno1oHPJdneE3CXru
cyO5ZA6O0gFhVJ9BChOTjxhEOAVFeHr4b88KmA2rtIELnBgFOmXwdNDOHgxQowGc
ji3UfrGbJ7lYiAff3l/bv7X8CkEUKyVnRoGGIRF91sNWJ+zgeHP6LXCioARj6dhB
ESAetUGPZLuyhW4GfO3oWwrGYbbXwv9vqOc6aAnO4AVL0kcVDcOP5A1ly+GxD05I
naVl+TM/K+OWCMTtdl/AfX/n+ET8cYlEciI06QdlFrkRJ8oCRtItFQzxyqt5PY5W
Sxhw0de+cf2/1Vzynxzeww9s5SS874HQFhRbz1Pth775Fpw1I6aiZD6UEsH/J3X9
zhP5sWlExnjVcEBTA/64iMCWIwwx4dnWyNNN9VdqsN0y55KTd2/8qFZoFMe6Rn0W
dhmqOQj4MMKf1bZ0M6r+o7EGjXhg3Io5nxORS+Su2XtpimPkpkjFuEaPyj1bdltB
E5KCzssIV+DbK34aTLblFeLEKSnptjg8fc1LR29IvxIc7d1IqFRrIynWS5czXS59
pqk1MvWDXZWy52gmM7MrSqDXxDxBHBZq5Yye0b5ElE8wPGbLaCyQn0udcMTJxdkP
CCKI/mP+fFsR+k+UxnfliXQ8CrmDByDSEeyOUbem7xovZsEdqkvhXDI2DtHsRiP8
kEmgf8JMF0kg32HqBo31QCkg7TVF6wYp/Ys6vYe6dAkm+uHqHs3jDDIAkzvC6yjj
OKD/9mbodXsW0jnR/H3BJc43AjsAhtaLQlJ4GO+ZFY9wUmdwZ0suyguGpzS4zqHg
aJblTQdpeRoqsZDNnM2rnTT26Bk61lAV+G3UtI3dW6l2NXQQatr2eOAMu8x/b4W6
9uoLUtvJaLockB7gc8THW5+JeSEDOkObpWle44VcpzMjw+Aq1Q/WJHA46tvgE/bc
sI3yk84+RwomsLAej1jBo72JJqTJSiRZqK2MiPHRu85E/Iw1zcOTRPep9bGtph2Q
M2cc5rjnkVaKhasO/OUa+tfs5XI0rWbPEYkfs7mwbE/nXQd46MO5DFonALeSAPS+
XJqEgrZWv1NyAhf50yZM9Z//5MrZCIjpxHJn9SBlJRRv4xNVrbuM5ZBVg16SXfP8
atovmsE72/YoYqzmUH8757eXxJRwLHg+x+3cdXAPXBilu6yFR0qah0sgBnPBSCtD
yqSOKfs9DmlExrjPm6cKWQsApyNGeHTI0IwvhErOsVHIZ6LN7IpQzICKaV75mpG1
Q0Tv/eVXnqg2Ej6yCCQ2THTp84Y1HsdLH611iHfXUJvaBBGc/KlVI7dLN+qjyRSH
8QjkjGkPmOLO1eC1ajzTS5ov7FTjKFNHa1BD2wJQ9K8KvsZPSHDValX7c1MGpEgy
gZT4c1ysZlivCMce6CRbRiiz9iYohbB+y9HtZ4CVAMMP5PCc5nf1q9IqmNM61WiR
8NeEgAPcegoRg5SQCTPesSyvtSHBQkqN4L9Hn4XfsqWdFhhd9ptmcRYY/RT2Z+PP
ob4Lu+OY7JM1YOEAleRHrfdpfSHyYXEglSbW3lQcVGOaqATCd0Ex9vCL+xWHtATl
VvDsysFtLKE/MX/mZRN3PRyPK4JKy+eKBoevOaob2Cxtffdl1B+ZgmjKgLSUKkXD
RsQy0d7pZG00rQCY9YjZGeucm8UNJhrWYuSA79ueCM530MzHJTLOQph+Wr/lW/kC
eyi4ViqLUHatqeWmE4dVVjpBSSRHNg5y9nkNyX57BK9GT4m02mI9sU1GhvVPt9HZ
nu6H09S/dbMWZCEkS+oFFQrmQyDB3lcKEAeJMNh5+j9C1m4nwCOnbA/PwZUrmvwr
4IFIHICgGFL4Y2b8XIwyEnPzA7dTbWvSnNWeVsdVPdTAHxZNBsWpzPDSw+Hx7dy5
mesbhWpS1qn+8mJ0A7buj7/razt2x6ZCogvooNIr85LMqzgNzB+fKX90ZtnCpzQR
TAa96QtWgavAXmQhxVoIGArI7Q0im04ejED3jfrCOYYK+8WkR4KahoAccs64wcCq
DHElp7oAYaI9IZBDxXA2lGvmqNaYEmdGD2FvOtOOHT7MHRhQlGWnINRX0CQ9d8xh
jw7gZEv9F1PI4EDicKI7B9IcVji1y2kCa4Gevc3AWJgHxmKZ/BSh0ngG6cBNIqre
pJsBuNWu99g+n8mLBr33xSjBj90jWdQRugeCLKJ8GGPVojqGCGte5h3uts4wz2Vp
qoKtJ2eusxU9EkSzvyl/IYJIlS1LqXjKN+Cw/dauH+QOOeKkTvhZdobfWV05ew8o
mbH0h3zQdnMafR12yVnIsRLVxs4HwyLcD0xWcF5v5Gkww7lcka+Zqg5s3iLOee0r
kaEbQ5o1SCyxY85pzgKNamdCVDVCFK0ryTgnWoc7zkI8Vn7g9E6OFz87NuARAU6r
P9mi8Y4j9EI41RgsWqkaCbXgfUpwZUY0wv8TV0b5aLFv5PUDfVMJZ2Me6VxKakLD
CHe5HfL/iHC4gFMPrsd6oVLoe7blZocERJJYe/PMS3H7cPo4yLmNy6PR3tRmR1Y6
AEQfa4YTEjw5WqcYGy78J6jU3bb1y3MKI8GwPHfCUNguXgoJNfmVGAGysSa/kdiX
NsYmSp9xnYYHN+6rV+Q0M3Zt5UgJl60275eMSQVkKYOM6/JW5d9/NueRvSq4AYc4
R8/Whs3F7THkzJ1+jnD1XitdnBXOhXnW4VxCC8mh0ToTxJGlEvAnsmKUfENKkCoR
oi78IAHww1kBa0kBilCKeiAwo3gM3kFzlripYyY+azy2Ms5hqnAUNSEbP4BGMuik
QMTr+tsVfrCjgXOjbV5c/hY8MFyR98TeKHqq4giRdqMOH82Imjt6zO0ecWQ9ke5x
W+IB2Twx439lC29wCp5lreiwPE30TgvxgSrv1I/HWKk0vuHrIUBbs2Jvj+L+3tOy
EoBfuq2YNuV8JXN9iac43Isd+axtXr7RNojRfUrXAFnA/x023arB6vON1Kb5JmJf
bsdwm0Pwy9lyI67FYOjFZCKGNPsyMc7mLawXXm4BdOAzqlfmocThuezk3Mqb4bs3
eMgy1EgLFmFp6T48bPU8dY/Nq1csbeJunRzevcbQ6VKkw1yne5MGzUV3FHzsFxR8
I7NPlWCIWQAO0BpPOb7lTsiJiI5bKF7Rf1l/syJJwjtOBmx6bNZPzoXUnlplBvLn
D/ipvTS3PAA1QVprVY32372MdSHj34UVJ/qMCJTOg4v45YaRS30H4pk7Z8iwl7T5
zm9jasjFxOohYCtcMgF79DFN4fJpfA5Ud/aT7YriiRHXO6gV5qA16W03XpC5Ksjb
8PcTs9h1zX51djiDrcSwJggDhgDCmat/2r54e6NbuBUYU8beXb8K4JXmQdsDAK9P
Kxc4DhQmb1as4ojOdRxy7jLPHUiu282tbMvrcgEUmXdaiA0vGr3qqplRLAAl6sIE
Q9Vp8bFLrlLaxb0V2Vhvzylo4teekbcpw/1mp1F/1grOBknQYrm4/ivd6V3ZGL02
aSni6ijVbLSDj4/HLSSDRe3F2OGnF8VQy63O3pG3IWcVL5oc+70XdmzK27najce8
Ua7PIt95aF9kTE0jLGq1teDLCrdXIrQTw8AejIAE5A1E/QDcxTsnASXTh208YDV4
XA8+N3TUsN8oGqoLiYu0R2ZQptF7n30CiSDHkPugYp5rVPqVTAxh3yNH+NZj7DEJ
X/eQqdqEEzRnkjcaOw68GehlG3X+e6pxfUgHyvNTaupGCwihGSVC6PCUQ3zkVzSB
K4pVrmqWLz4jEyeBd8R25gjF1Rjf/4Mgdk1IxFnU0Ay/Z1ogfKNY6A6gy51xD27Y
+XJfmaFNaOir7QnXkO2oUkn6cAhymvk4tC4Wwy/iDSrWLjK1wGcDp9NAbB+Vn0QY
VQgiQHLRif/zuubWZ4XXGc1zkTSBWqAAKBsvp6QlRN2GHsq4Hrp6oblxKvAJnyCz
sb/s0eTBI3oRrgJr8wZLE9Qw01WaRUyXuSQBLuKVAKCe+39a5r2MfM7Zd9Lq1egn
9RiFtst7J9vQP2bZ1UgbNHshJmAWi/s+zlnlaue8ZAiBsgO3VzdI6lNLXGm59DE0
Ao6/nTjdHF/C8y4l7/Wx7c8tZipNEoF1zcZyC2d4A3R5EeO3PzEZjknZ3kcz3b/C
PPu4N37XDmxDGd2krxKwMxeD03Da72Rn4KpqpxcYQYHaDl+bt/3Ol30pE3QVwcKg
GExKDNrGBqoIsIbL/QrNc7Efu2dC3/mGf4rLFutUIvU8LNcbT7bZMw6I/F8JoVfs
O88aHluzvofjmYZedhBY+2Fx7hIrDh7jVxbdgj/uSSSadygnp92nsmvr8yHQkAKo
bw/qvstJccGT0Qd0gsHLv8RccZP04GLqi4HjpAfixqAVUStxNi4soVuYLGnotNB7
TuNAaJugtYjqX7OUcTtEpRUi/3XxS0DTRU2cd+w1MbNUkaBvaAINDRylIn0n6kzr
cXU5CQ8PKbOb9q2uj3pavxp4p/aYoaR7ZbQ3RixZuh+BNn1x+OxwdnsOJVA8G48G
AzFibQ0Ki2Z+Bp8pSZN+Ocnbg1KyNEDnHHuQUC7zqrZ3Bu3gv1z2M4bPnL6Oimaw
MueaIYMyA/kznLWJa6p8UJr6zyoiZ0d3qzA4oip6PQKLrtOK/NxD5OdlSCBnWHEl
M//AzYSi+QA0txAMPHr+kYdBWwSIQoZvS7xhirgEsamI5rsIoPBKCZ4VGPG7X81m
PfpS+P0apCLr1di12MzVPgBdbYIYfnrZ/4iNope2xtI8zBc0w/oc5v0JFzk1JLJf
UvOP44/ga/e5XuUyKSkCKw9sQXGN4vF4uXIRaKVR7hH1fqbbeBSDqJgbbSFGJ2DR
TxkqUSM6mHc7v8hyLwdqYJepb8kKyD4XqXNy0U/FzYBp67/TnJ8QY+VBaiYI7Rmi
4d3LiZfEnQhgnMO0C6BCiKioE6292Rz1Ox9n5mRgW1HDUb5EAeG16RNObleK+UMK
y8VI4+wWJvmJ0l2cXhq+v6XKmusops8URU4Etvam6ZIpl2joQqidxvTJD1SHXEt5
j84oUlKg2LgXDl6mK38MnoeL6EIVBDgq1mLWgrazrpESlgsgapcGRIMovCkQ7XgN
WFWk6+mFT9iVs7+L552v454KtLNOY8e5MYPBXYyXnzGvIjn9jZeOGXjKwddUIzX0
LmQtGtTScnNFTwiIwq1ar0LwJo+sy/F4PS8b+nM/J56r9mzHQGZZs3PsMXKYOndw
zjYNmbZTU+bd8fj7p96D36virX7yH2KYpCgTpKzvyaMLKaGj40Bp8M+0tet9bVrV
SDjq7GkCzjwx10RTa/41SapxexzhaIcks9FmDfMBPDjy541flQ37YRExtdyGjOyA
14zJN7ZJRbSCyfVcKMBxmcDxeFoe1G2Je32yG/fvVR3O5zo0c5+2lkrWopR00Bt8
oPl68hd8aLN8SMCJOH/RDkYFsUlC4XiXwQKtgJzZd2OINXdpMZP16kr0gMU+IQrs
CRBzXP8LPjZuuuyjpy7gO0pru0x31/VEsV2zfX6me6lA4Y2aW6eX8luPKE+Gj2QF
sgPvgoZnKiWYVjFe/rdUmjpaxpTe1V0RQWn/+RIQBX88MEX9eTJsunzp3ULGbDgO
GcMdCJb2zat2D8QkXliXMCvdhft10HPLzDL2gbKI0kpZZwd4At2QGGRT2yhQf4cs
zYB6AMuFuIm4ZIfqI3IQaThouHxwMCCgjIXiKALWwHpUFmRcaHXpXJQ3KJFBxekK
fGmLJNyG4q0dax7KMfSkcfqqlajc1cQsO7fS7YPhI5ernnczLCVNtwOBU2qk4W9G
ggkRQMyo4x4udNptizJYr2w1rUchYTImYmbmGGEj2WhQlW0gtnMXvQyMa1HJ1TUx
piBE3+InRRg3X/oeFFrcxACWIsh95M757wE7QKPko57Ay8OicrscBWDhOOswN9G9
ZP3lULBGkJC84Fw/en73kV4hviT175P7znp7OMfCCl1IDLS9/oStWvKR7g6wAXpe
GmlD/kTv3Rxnk+eLGCV1IcYl1Ud6AbiUKc/fM6U4kNKhZ8comd4w3qnWBCqmLE9O
qzRto8cFD8obGZem3S4Xn05equGU28nP5KYQxOCfYroJIsko+m4asMpWOYJC6tNW
tz7zW2jNI+FRjfgw+X+Qfa/yBmeFUnuvYnBn4R6H+8I0GRQSlVaFLlM/QwxwZCsn
hJW0kUSVs6+alhUHhLvuXe3GgggW3m6pRuB45faEaLX/CWo4Qz8F8JsKHRN3ywnh
PIomdPYpuNxi1hrTZxeXir7V6eO8TYIusjqrNWJK7KprZ3QTxrvScuyshWl5cKEu
kSNlbYbg9y3odyfCO42HaM+2tiaksrESP4LK6OtOj6vYDvWbYTyW+xkDFJLeZv+I
hGNkpm4l+4W1IkJCXhJo3WLtpNJExbqvqTBg3EKPHjmdZm+31IlxEGDTgx+BcFX3
dHDnzo6faonDyL4U3cn+AMRp7RC7R+aExujT8D5e9F5JZQ8lRx/ScY81GZoOLNdg
bWxXngU4N/2rgoMUnCCVHN6dZVNk5hsInHwwGQ9dH2hQMboVEgxvCeEjGOj6kvub
rnE8HVPAMla+0UIBzUkc7bTN8mYzNIDkUHptkB2Oxgk+stjA9fPbkRs8wRiNx/Al
CX+7+onGLkuOAAiBSILzGIf/+mmb4BXUOPzhL00FYBoAvMXLd+5ACOG4x3oqwm2X
3vE3IEYWpLqBwdrwNFZ1q0JpP1DHCK8coaxuEeqKIaFFB8aqIUxXznMpCt0Yh03e
a3bFNRj5GTgcOefTKMTz/BdoMKMmYuKCAeUSmZRxHPFElnc+4XIPoN6wm+ABeZ9M
t1xt//Bi2Eyd7MncgquSTQmjlUsqE2i8oaTTya6+n0kBAxiL6ld98UcoxO0NgScM
mnwEFE8+zLsu9AEp1YTN0dMoBSkQIfvj1FgcWy9PnsrpZaFv6+q1NNRfvFZMId4j
qu3D4Jc8TtWB1ZDPyueSdG5rnsIdiaZjsgc7R6abCjxRZ+q6lU+rhUJH/bkGPWA4
MQms9tu5kKUIxC3XeQCfu92R8YhvM6eYcB1kdVk9G/z6q61gNMBE/ns3HS/5zA7/
LrbWMxImX3S32waVrHT41OhU/PeTXyGqJpK3QIpT68fEWLgvYmHbzlOtrnsg071H
w64E3OYU2z0MzRFx++vf+ZGGIaRsYX1mD3ES71ceyQH6swHXLre9GzQQ7vMVkWWF
dXKoR9tmEfR2MLpCRLoBZUUnfO9ybg8J+IP991rkQt4q9u8J0zAhyuYv2p1bzjaq
+L0O+3Mp5hDL1wwh6zPQ2fG0XQF/NfR3q/SUxJjzo2eL1aLCEuwAKzi47sfsDMpD
dJrTTwoQQsiCKeiGX67dm1hKwcG7jL4r/A2SaVVsTFCtDHdbkeOznUZj+g9QjNvP
Z2PSAkQbk6xxr5QLD/DREUrw/08f2Q+3wuQu9PvGsb/6TW/BJIY7WZukf0o7W8YK
2LGveO7vMm4QNi8yL5Jh0FfM8RGE/7AeHB9GYnoyQD34/HbGTNekWV1kf7gmMwwV
esIyJ4mAeWpmN4+SCvfGckUsZv8uSG9azPdattk7xjXJd5J6NAg9/4PMzbS9G7eh
mRRZk4jMh3m1mgqwHdmWeYpM3tBUKOObO0ysYOfELX0lc11eQJghtgAHYERky6hS
Qvah0msFb8hGWHsv/0VbLyEpLm0JAViGxUvQyvLt6dn3eAMoyC4vxE+fepO8NHNK
0bX3gEBB7X7uGhhuBRO5y+QWrIuOCPwtS5xWbSUfn64y6b4eImSlf27Sij0GPISf
uSA9g4sbeCkExhX3BOBjANzFDIRsr/MXsUMyNu+bGbb7wwu+3IND2COj9zcUBsmV
Ihju/+OMNFnXGDQxyDBqLjzQFxn/EWRGX0exd0sqVvN60UdtenfC+AwCK7yo9Vgl
AoYrlqwnPKGEwkFAN8QFsCONuWs/FiL16UD9np6IWwfhz9ofcqZvqgHC1N2MsMnF
HJQY+7QX3+uXqrSvzeeZ0KLi0OhT4/97MzEQKsbyWUJ2CYOf0iB48c36+YgKuvV7
fme/m88X+/w9FRYdkWn7eOewmIXAh2oHaDjoPSefE8BmsQrk2kKtfF7cnhpHVsXh
6bxrMsxEJBcjrcU1aGUG2vJ1WbXJcTAWOeENvmCZ57ZhwFze3SGdo2gse7p0wP0I
v/knuGtaOWaUWn5ZyirDkL1KZHNVBRXKc53ZijEqNJSdvTPMos8wVhqyLWAEx2Cq
Zw7ciIgQF0ZDvj5iDIF75b4SweMU3j24DDaMuPrqDs35LxucdMMX8VYGQAIGRogp
fPvu/TwiUl+UAlZ6YbkLLt7q33bJkjxXTI/l1l4YDrJVj7u51dPSIF+mxi4i0/aT
+nbl+J7cVd//Qm7Ztpy6C8lJEB8IhZTaAopylsHKfnxGdK43KoxoK31aIWNd5jKk
OzXnWYl3pnuvR+grJ1J/xML1rUEDbNQPiu++5ffdekUiY6nt/5gq7adhs+K2/OjJ
aHcqmY2krP26/Op1KFtJvSsx8qs0tufqcnSwww1XBiFYhWoMh9oqidhZK4EXxmmU
aFA6+Ex9ChqhrdpJjwrEOYNSiUz51HTcVPhMV4vWI275BlUBWAA9umkRcqtjA37v
PVn3qQWuhFHPH5xLgLP7Bbvae/LveCP2o/0mRnLUw5wE2cF1sW4VS4EsHOGY188p
mSo7yoy4G6SVFX87AFT1CwUCeOl+8Rdv0F5sGw1hEmsjd/ZJc0gGz6/wujMD9ix5
IEtOThGqhUa01gEDDvcy4Zml8Nl9QR6XELqolWeKhSt1/qG8fs9kIUb+7lQc3lC0
CJWjIT52Ot+1Y+YzZnVOPKXzuoz15FYisEmyJmzE1NWlFOyd6qLJCrAFR5vB5g7h
VS0FoOofbkM17SALve5HXH6Ma680C0SvAKyi4z6Vrn9FsKpUdCUmcAk+i85oz8dp
xFaCVFTf//GAVGvyrpQRIjD6o82iwidvzcLllMitDCJJf2ypobf4VmRfmYhABBr2
PxKw/7gUFrCL52V7z2G6Gq9t3tttKdBtF59nCchnsMK2ypTllLpfxYUDNHWXKfDT
L7LHwt/pdxWzkAPyi1diwrS0wzt3CLGhL0uyiopidK2SMOGOG4PBBxptyrSiP6VN
pSI35iAlSdkSPubZt0b8PQqh3HqIlhpsTaWLhG6tQuRoYkCmQmbFZ7tcDzEFJ1kR
zYeFOROAa/fCrgJxK5ZqI5+TWvQm2/zd+lEDvnsrXDFpVIq/FoNRDMSww5g3XEjl
FegoVb8TzXjEmQfkHKSoykom9SUoCDgxzBfMy6e928+fUrpJUw9lgTGn0vrwBqjn
ypCg/yBrDzXbSftxzLrvpWsIWZr3q5xXQ/kxxY+9duX0TDeOs6xYm304jbi0QUJR
B8Z1zXU7ykIeUKysqnIdwMy4YZM2IOknTtXAqMTdYa6EXwEIpWtlxyF0mNaBfVwk
XyEHdPoekCxA2lgxAGkcHMUfLFAZHbiHrhWsSKbHd/8WeJ+pohKkdvWH8Lr8XRbu
fHfWaqCWRMEdfd0WsJzLgzw6ADYpkPH85k0nTaFgztk9ESv4VxeL7Kg3W4i5LUMG
P5ohyCwMVv5SP3Rzs6GCYtSlX1064RcoV+6YKEExCHaGKpWRBZwvAO1UbDdsgzUF
37t+tZjwEOE6BZ83fYGO5c1MszHVNKkGajsH0kkYllsb+Dq0Oi9wDDivw+Y8IMxK
3QhgJ99Rwq5Ag5bhZcUbazj6n4fezjoJ2o5ju9PLXAl4204liRyad326x9TFPh5G
xBlC9dOR5S0Zh2fCLFeUMbBpBsmVqFwL0rIqth79qBEFjogv4uO3DHulOhmnUXB/
qk5JyVQ1C68DglQtUKEeob16At3YQu/eaVEiOilPRH2w53LnoBith46dPmWUdctC
mws+WepM2ezPfhyBQFgcKqX6MGFvdgSwyFlFkr5ox0NGuE6nZjEq8Smi0WAhvYpV
8417WmH3VLlK2V+5rXbXVy3IF75YqEK985V7R/dv9B90nYyrqaqUUbugFFu8CCg2
HJAmfpix44k0MifeH63a/v/oMvc/QgYYyIJ+eaPBIPho/+7T/ICOt1k3xVYexI/3
EFCIPOYNP9xdkocjyIM0g4JIfKYfMJqbHk89OxbAFReRx+amja4wOHDPVYwJMDAD
u1fpSWWeM+bpzx//Y4MeheoX4Etu2TrG64vtJLFL06EmqrUbHfhi3j4B6UuwPFO6
WaUmgDknZQ8N9P9abei8TP+Gg8o19lQ6rWmgojLn9hzbVW+bBVrFGoHVAKpsZ9LZ
N5IcpoUQHjllZkQzvfs7NJETF5LqBqAiE4BOeecvNJWJi4va2557WavyRYXEuSyn
0YNEKG9DQa0recCOErAAW9VTirotY7buP89OR+WVsNm2twqbt7o5W3L7XBchReRd
rOsnDMiYfitS+IKQKqqdbcbYpE9ICgwDf2kenSeTNt4ZKK8b4xDFDQV2YRWZkDvm
Nmlv3Ui4CNrvWq+IT+/f+HVV4vKhngJBW7dEYTRZio1lKzbVGdDN0NU93iju25j0
kqpC6hzAciqYAZJ0Wxn6NAPiBhszc7KuIfTTzeisIbtqIsIBYC+zlmugYjZU9fDa
+hpaId7jZvpt9PzHkuh9x8P3hCrdTuMNGni8FlA96UiBmpEBwwI9l273TA+MoaCr
rPHQVNVGNoS4KBvYPvrHexiKyNBfWtsV5o6Gf1sqABG6yr3HsqDjwz0m8T72GHBY
//GK7O/y5OD9QsCDYX1IzVudr2v916Q0/us4anFugfsvSjRXSXxM3SyzyVIaiduZ
Vz/aDPZaJJ3/ruawOlytw4UDsXySFKjyGWCUhQP7oMhDcUEHTbSNj825gUByYJ3u
BPUcYGniaKBrEoUNrHWZuxLKDmPy/gzmNMrcPpzOe+ikUsWSqHczMzByfF/1MKH9
9e2fQMQCi8L2Orm7DN12CMvCnant2t7FuP9JimJpSUvfb2MR77TiElCSLAivPLG+
cHvWSIb5VPdkUBYaDeRvWzt7T4S3K38t1QoibPsREe3Ww/1zAoYbw4oEK1ZqR5nB
ATRkiNvNSlJmSmOQ9iWsSmCecd3DZuKTpgrAiXYzEowfUyJPiOQFojkyDUzb9LWO
797gmMtJ3f2dy+HeI70jtIiD4U5RRDN1qoZuhsTJH+HZaD2trITrqOZjZhJc0f2s
WBXKmomyrCOD3gpd22d/RAyUinGKXEL8IDgb9Otof1Cs5yiAtv0hOarlReOfv3+6
X0X5MKtAw+0Vt3Hgb5bqK3ocfE76tGBP+hmlPOTIPIkymVva+gOfCbfE1yCYibI1
YgQf7BFVmKYud5nUpaMXltcagADv1a6u+9IaJ03ULcMYWieN/PnbIoeeR5dxZSql
WnNEVv2lOVQj2Wts/Z0D7Nmm0agY0syRViQlXU98Yz7o2DlTZFqie9wtuLCgZuEE
037ALD7fpPF5zfRFx1BtkIschmTdT6pbfylBAdmqaZRxrxqKMFhfARPoNb/zA/Ia
ePMMwznp5wbogKKs0YOA8gJgpKdPW4E4fE22Qw0jUKohQHSpa0soAgz39XOLb7+3
7e/IKCERPb3McoQH2xeyDr/vYdQINoo5/AY7gfZEanHunAPb0wTe+YAEUPDv6mZX
JK4GhQI+JI8wM96hzoWqwatJ86yiq7oXDKmLrJfzQr10ss+nKRJKDFI3XBufNEdD
OjZNrbLWnYIpcEyWIXBvfO1JFbL/48gZVJYUQFDL+kWhb1tSrifL1kTWvtmp5m5+
sLD9DWsDBx+NeSIP/ijVEzKvmYpcz03n21W//542A9YZf+VcDDWJebsI/s0OK9Z+
bCnWfhg37awXAp29EDxGBaTGCq0WMV8eEDQ2sBUBAOg+TFsBmgERN/jwgUQyXacB
9ARvmQmcKR2wRwMaOJ5tz93zv+PvRZnxkGwhFSHTVwnwSITR24hpn0Wqxkn1oGoj
/j9jow9caS1M8IHacE5aqdMLWVu3HYt0hXS9+oMj8FgTQ329Gn5K22JkQwJYrgKu
038+9LJHOfSYoxegEmkjzXnfj0+MzccCxqmJopeK8xx/LDA0c82IvPWnn4FTwGz8
6QAsBc6Mi2R0uHiqSaqdUAyoGT78Wf7DMisH5dnF2NXI8syQ79msfTk4W2RC3UDZ
SkwhuysYvvfrTE6O5dT2u+BzqPvO+pfqsE04Qa8B66ok+CZ+7lrODqIehlX74fns
a0Hd+dh7C/8KcSTy56ZuF6jJdIUZehCfHTo6hJT6c2sYjgzPaiLU1YLrJN1L3kpP
NXNTRM/FVP70lqDx3i/8SNCkv9Asiq9CPfnR0wYF+6Vaadjuv0scMkje/VE8nagv
wRKNpJDnSKpJD+cOi4CXPh8qeW3FgIpltqm9tN4PYs5BB2FPYHzlJ8XLd9pkbjbr
sWjUW51D/9ErDkFpuSoJGaJO/UIVW+QtTNTjr3RyVek0pUsAMpHFrRHWm+1GVnwT
MQVmpwlBS9TAHZbtuF0JkS+89hSMfS5L7atoOfZBFeasgIC8hAkrLMi4Uux1L8N/
Roq82msb38GiZxwx7V2OH2s6ot/pELhP1s65aFhtPGpLsgCD+xiWIb96laA1+qIZ
NSQ45aogmqjCGlQiZRb+oFvgbFN6iBmu6j20FIOQUR7s7NuRChQAEOFkUPmz3fyC
73i5O9c4Op0oy4Ft5MobrvrkB+7FzfFckS4+bdHgwGuT2DLe6M9Vw+lqsmKf2dVt
4F/1ESqsZpC8h8bWM8qYScsp9aSzAjpEyO+ey7B6DUHeALKV/He1Q0x45ia69Y0e
5mnGQeOT5SL0866JIM4QCwjuhZFIuFD2jUO6YKrRXDJfahuhs9rNBsdpW1yPQ+XK
FNyU9b39dWPsSvtP1tHzrVp8C12v1UH7/Fwytjt50YT1AunNQrTCwuZf963CEIkw
+Vst/t7MsBkb1Xn49L5rvugpkfuM6WMah2dYJ1naFwTLw9jN8Z0Vwg1hwJ+kOvwc
o/q1FbBFjcaqiz9xutzg1VLVNMEIKB3J0mMBYzKuDplwLnxjhib58EfL8cQ2jktG
V+uNCObEZMsDKYyNFqVtLi74uslli9GjGXpJl8FCgHJXshDKp5BIjA7xBCn/BRYi
DrAS9+SMdfB9SjbJ/kindXKsjirDgLennOx6KDqzamRU0qFBk9Ju5yanSktnIQy5
ffj7HKJXxXKEVDZWsw8sZ6bSsCGah5XaEZUIOQmUgNTk6RuRz7cfx8rmxAY7Kv4l
hNJdz9Go2pCk6oQqO7v3ulPrSCeM3lyf8vgPSIsvjYoV62BXMqOhOY1+JuiuEHma
wC5iUb4GuwIORNeyYGNXiiH9Nk/x0uw2k5iZph6SrRXACuvZpmAQSeJYL4KPsIyr
YqCLcI+cB2fWozGYDDu7RWU9d5eLFwjcoYci5H8/nu8Z5x5pFou7JfidvpR7zwzZ
J9hpEwla9Mc+Eo9S7xacyFXc2SyuNmnXRnzA9IWZS82JcEC4AFH1VeIXE7uQCdjy
LoRsMY+iSdHOgH9EpzwaNfcYA1Ch4e4MpC1I8RhM/p+pGtMCaESEqX3nH+qJBzuf
Ul+1YXXnP3WZ/i822YCVgCeFidJRw4LDusEcjUHD745jaxSQeyZPnX58eQaLicw2
L3x1VoPzQYHU2XoY5Duy9A8JORdOWfhugvqYjkJdk1e6ZeOc2ufS/vB9qOONMkSr
Sb6IqffH2MfipHKGPEbx/7eS2MCPlGwdw3BJ3b2128uB+lXatG4/plOdQsOE7OyA
J85IYzaFs1a0nEXgh2iiJ6OB90WORlgceUpEtF/MXsyMvrCs6Pn+36od5vsp/On8
wV6U5z3WjcX3Z9/sRngsXymUVADl2PcxHmVMFzo3OxsolnTOklH9L+hGaBW118hM
NIHZZs1ZZ3Du6jBYcqe8Yv6HjkKE2hm74e6QiysgyWE0dbOvqkYyPBsMVdAnO6o1
a0t2rJ/qraWE3qHzUZiZwShyMFlWEfaFMYgMrQ99RItAQADgI7MtRYS4RNMzdgMl
lHaYeI/UXK6tLF7fd/4Tshdy/ha0SjbLOZnI+B3pja/Jq0Vbb14Gt5y9Dz7Cu614
wdDsr+DsffA7el370ng0zF/G4AiyknkFm824T94N1rZ78Hb2WNy6QTGwe6riKGfz
Zk2GH+V5LMYTrwBq97v5f+E1G6oh9YbjbAp7NImYaMg1wbl2gqsenV7d1gwMyuu/
Z+6HJm6IhTiix0BTrG4fDCnuf2x6LtMj2nq4qBRXK+7dxXwNrM0PInqGNShCp2GS
ibS9X5Nq/QZp1BsjxLqgiDLMFpHQkVi7l97FpiUFGJgPRvB7Hi2vpca9Pi+Gy5wU
hXIkW2gTZxRpCwISNUrHJIIZQOitcimfux+/RCMOHOr9K962K8FfoGISX2mEpELn
txyX+chC1X4b8js5XwyTjBblIluvL7s7f8Pja6CN1dy4xYpjRT4pFJH+D2YP1FdX
DtTowOOgJm7wxv5cHzNWy7lyMS7JnrIQwWJqKat6NaXRyLHx8Ogz6zwtC4OmgwhK
c4V8iKsExpydu8VXKLgS8MlGFqPmflsMKWKlzB0YDki4gfTgOnDxvWVIW4zi+nFG
33o6ZLWhSLtWxpt48IhloTtv7E9emswctGzv/h+Kv8WRs4ji9T37D2f3LDifJ9tq
BB2DVdar5IQhqcH1GHxoD5wTNKQ6E9nWujqTXAiS3PH0uJZreJsUELZcb3rnJSjh
0AeQny4cdY+FnrVTFvaBb6ATAQv9A7IxdvTrXJRUcM3CiICEi+4fkcXS7/6EoKwA
S2mFFrYPsARBso4HsmrjG8zAMcaKpRP0Q5OLBhcFMwC0r6G++rrtI4SPbmMf4Nt5
S/owq3n5XgYebgPZ2nkVuGFP9K4MGAPM18hwkA8bPstIVFelZD5bSMEolkl6stHV
l8CK7AkB/TJHk/9R2wrkceRHvDaexmBqbraX5d1DgvYs+Po2LQ8QLIinaGfyNDVV
IRlcKVxhQFz80rJhsM0q9zMWATylBH748N+ciPTx4U3g3QToQMdgDUjYotNZbzfB
GiLhTHTGT5RsGfUJEMXPTOEIAr/Sn4PIfM2ZbktJfI3hdSJD+Y7/6JncuPC6cpeK
s/CtMbTtpc5Aq7ci+dy/Lf3/PXimMFVuXrLsANEd9xH5h6D9guMT6dPV8fMQed3p
6Cy0OGoJerigEQpx8ymDX/tGGZh/JN2pWDaNTTRxcdr65M2ySMO2djTFLtrObflH
snCl9aomApqQXH88QuWZgXp/5NbEGCP1q8MqO0RUv36AnBgITE6inDnxd8XFHarD
ONC3HxRRolx/Gxe6tXZi8FcwyfeG5Ecot3WQvaN5nF0hqlI2T0Cw3gnp6n3dqNAi
QiD2YmT9sbL65FiTe54vSGOhqjX6JM9SpuEv83IayTNSWHGpmdULk1kPQmhzIqoj
ebEzhwioeUNgq5ptG2LU/N0YIducjhA8+aq3ijjGHsddq7oF4UDb2zwCHzyyebjX
ELzbRSZLNSsyRxBFJnSr+fB7udRMGjFZbit5ZO8EXzFYr3qxeZZ3XyFGTHFDW3Pf
5sNgFV/7fmjvOs9whU/xTTxGVLR9FJIPGFVGKJvtUgO2V3yS+dQ+k7vsGT5DeFk0
mgEtn4Dz7aJE43dagJWaXwjJ2Nb1A4IJgGXrBgJzeJGbJBNNKQts39qXKYvvjsNo
FlyLlJESWl7m255QggOjLumAEwaJuIHs6fr5O0XqXWWa7ZZAof81ENdJuKS+sWIZ
eVkMf/geh1ZiZqe2kfUwnu4tk+e8ndxTYZQqAUQirH6Gx7DHmZcSX90kBuIGM1fN
WsnaZQDQM4pAgkDffzsHBurQyBvjZiXQmu+0/Tz0kNtTAJP1XSI4Jq2mRcIlDt4a
tSEiVXhy3IncF5oG0OSR5gmXAQZv1PuccwRXhuDkjM7X9xMxBtHIfFci6um3t/YX
AGTOnoFYXMqwbioOwoN8Dwt3oR2SQvGBoiEu5z/xXchYiAkJo6Svtq9sbB2DpX8E
4THCPdyHwOp86TC+xHUmnvy0Nt3tzZ4pKqDML9qErS42pSJJ8lZJWgEP5L33fMH7
MJsfFjZoOVtHfCDpj7KvKk+US/FLjfQRSbRFYIXpcI/th2zJcPCiNbuOE5ONtJgt
OjC+g+ZkIdKnaNKPGK1z5b/hXE4oED0uLj+Twyf562nC4VN9RRD3pnYwd4+EmQdn
vjSwaRiZ20U1a9hX8Zj8ItyF2Sm3V8Ew/xh+HOq7GFyBSdcRhySHus1xDh6+sa2o
FDkvTW1Dr2tsGHLjWdfM7Mj8hpPggDKaJBY1C28dh4lZ9Julp/VFTjanXyhDrfsa
qeN52hl7L/9SzL8EJWvzy4hbkgxpqsgqQJN5oRukWOxYOXUwn37Kbp3Kpt2l1Imj
JrFYI8ZOCk/JrGNgn79eQwc1OcPwaciHBPKZjQor7+dK9Z64Pq1w/KRkcUHGs1/N
Wi6WamYfnM5+0h19oOjKtxElieEviIu+9WCqQ7z5O8npmyunGqIvWZKXILH7PM1R
9s4NKYe0+++3IxKlHNPcjppsgCqxTJmNXhkdSSzikzuM1QcR2x4xh9yQ1J0SsS5N
7js3IgELkZeIpCX7hdLO4qfSRQMaKJlhpPSctdPeJf9iQDmQw1952txbBG57hSig
F3pSz7GOJWLFYzJLlRxdVQgid48WVrno0mRPOTgKIzI4MjVkb+nP8cFQiHnA9eN4
uRglouVYXrsxuIwPKxQ5X/PegLW/STo5F4e9jgnLOqzgu5W7a1AsGY67KRQ45U1s
noGCnH9RJWYmri/CnscDU5FU5D4O9Ob5FjqbVPeCjdZrCw2oLyb98WDCeY09c5Ru
HPfXxeoSM8IBX6q1u+ScFDfvOZqIPEhFFGSNs8PM/ua2xRMVSm5NqeMqrUMSA4Vi
eR5/PkxKVdMIJCDP9gcQL+IkSScPf156v4UxigtEjNQ52tDoOMFRZO6pnOu2RRx/
Wet88bzgJAqB0c9zdevLB7QCa75bQune/TphBKHpvGi1nDX/rcOx8slq7UdoDG8u
Ilg8ynxz7vdx+8QL3IWoirjksM1oEWKxXhJg8pcVhMHnSw6EkC2NfpvOxvnhLJwq
/2JGqIV7XpL/glPkQJ+MM36F690BJKzg4jSGUGPDvGiZbshR/KS63IKoYLGk5VOY
OUzbc74wVyDdKvZ/taFVLs8MpcmBa1aRSw2k/uHv1ezVWxBCHhF4cC9G5o8VaEZC
QrL3TwRLoc+QKO9bPAcoeoDet2y3ExPs9/+Q+BAfneemnwZa7tL/Szl5Wr9+qnYu
63EIQBVyGhe9NZ07lclP40fxy0obB/1CpeNDyPyManZIMB0yESW7h0NBNWsl9uhR
ai+0ygq6zwUhqIuafRn/ywnub6BsmV7781mtTW84d6ccuAOe4uQoK8Q7kTA6X3JK
aoM/8ibnBLVpfEqphQTD8rwOVdc6fKhOmXZEOgiRn0F6N0r28PTEf+245gA7dw4T
z9Oaa63ws+CHb99NzrbfgFcCPm/FoXt8sCE4tZYdKchEBy7IvnKWFQW5Oe8JdwLL
a2eOspzBGkrekahOQmcoOXRikq+uzIVQYsVXf0GfJ1I+WsdNocgx+Jm5rlzStkv8
0rPWbMTjPslVzKysqa3Iziz6DqO7mW7UDNrPhjtJmUz6Ad0p2lXucAGMyxmgSxHr
4JKSFvyn0keUItYbEgCq7/mW6kpKnqugHZXDm9kctyIuH075k2rPOZYLp9+gCqt1
RXBEOyCO+QlaBm8D2NwaVXsNh0IHXGIfcnAPPZxBF6Pks+VQhr4duGPjWKYM6rxJ
g/LYRIG1NMVe0PUy8fywhE2QT0cHeRIjgboRllHibHziKhngZm7onxbDbIxKc29y
/E8FNnudyv+68yO5wgVm98vEIuJwwN3nNmsRsXBg9T3GI5YK86M568D8SbDHdQMZ
NiD3A2x1kM1TbRtrLOVzwYTzbx3bnhMev+TF1+VPEvWxmzzODfOMZWr8oIPz+E23
TuKbgBklMVK/M9hL9rmVQ51dQWEXaPyrJHWQA2p9r+96nGLfyii87bwWkFNDd/YP
5+sxcfZlHk1ZMuavOsMFSZyD6sJWfX9Pw9gbYsLYlxPp5iBTlHT0qPgv9uFQ+IIU
5nL0M7dbVtS45AaDHMbn0lZd/zEhUosGME4UgtxK+ie8KNEBzYpC6AFbWKSSzVnB
yOrC0s2158MRWaW1naSzPlKuPmT8rzYOmVWutrHp4+nrKzyl9prNgyiN04NEOfEc
SL4aJPUcmUEFwwiM2Ah/FwdfCZedm28mn53woDd8n0Pm3bVAWhBLaWkHY0crr5mx
tj8xOGB3o9/1WFDuycZtl/V4MyfrRXaqqI8LZnxDZlQd5Qvlv71xUbEBAiqTBfm1
KIcwd9RzkqjrTnwTZ3lXMdSu5YWc+deT54vSbRDx5hvMA+Ooqv5NzrOfDziDPWr2
KlrXdf94RCAjR7+/YBEWJ/Ja5DgYaMuH8qNXzuZDEO2Ca9ED8E6PXqKDSU+NgXBc
3H1xjC7Vs8OUUL3832VSR3+1enotRjoYQ188l6uWVlHDLc2h4e/oW/oUoxJweE9A
oqa8zEOhYKfJQiBrU+ioHIKk91Q/gYDOhgl9dv0pCbYNU1/Nezyp/gJ3zPx3NGx1
s20Xu13DiYQiUcTkbRw53u8SMSGoyFJ1mr/zMgjzvEN77ZCUdsYno3pMZ+DTmjHN
+Gp+2M/AxFZDCoLU93gyLTeSD1SUj6GdBeB8QoZz05iogUeMe9lMxYz+WxPTE9TT
u2H0OQ46JyWKFE+ztJLfKr5WJj1TSbPnhcBy5z9+OU3yzsagSrFiDqPgFulnI1lg
gD9vZnKyUYTrPpMupRmncNmyzaSfvJziea5e/9c5nyg85f83J5fEE4li1+OvWKDH
PFjBTTJQftQoeNLe0M4kewP5gBbqsc2PtYpkMSx9hUrwuyT9ILY7Ur+eW9gMu22y
7kx+qkU9p8aIRkLeHfTpfU6Fd+EoM4xluZpt4xKWcUYimtzH3HfO52fJxWvFbzRd
a0XVkh/k9Z0ayDrA51FJOt1yIQgbd14TsHMfOxrTgeJDsUHjYolYPQoe1VxCTnrm
MPBXwCC2RHFISDPGXeB+C9Dfz9uvkocnWgxCe0Ikbz0MKWqDMfLgsvWfThgVB3eJ
soaL03AePCxjkhD9LxGpjy4ghfYpM2FVY2G6GQUfSHMtS6lhvbUS32I/kn0XDQN0
sRWoAx5F5LefAfVH0L1vmwb5BWfIx7w5BjcrnRkONtk2ZCg8aDk6D5xSA4aAEmYp
rInmNJDsLU3vfhidZqy+lmYURCYgerx6GbsjPJIP7c/OeJ+X0UlyBYEG7ediJVaD
MrzWhm4nNjHpV8Ut6y8iCrqpXCbS2cbYXjmj/fn63dIAlNwOjfWiVrmipW0+Ht/F
daXJUWZGrt7cF+CbVhmcqnm+8JYCD9Qn8ByOWDa9QCiXXmD3czdzORe5+gCvmLhE
9331Xo3XtiTg1yxKVpjlOSckjl+JO0eHBiEC9QjxANJwIprb8f/6nuUjWntOkMQt
OwagLPZJTz+ce7HoWAQl9bdq5b0I2/Cc/AEsb2y4namuSxRJxA0krNuglsQtqhI2
fn7hOkqlDDwTU/U5y2xxx29k51NgAIkVjvsIvZ6IuBKtmPU1jmoOXqTmu9q70psm
mlqwUuVGSmaitGNDb1hX9Gzc3+xVU1ERYCjgsNvs075IwRCObVzKV8gBIvXZ+2uG
uHqRAgZnpRVK4d130of345u7zJI3N2qt2RMojiXKpLDgMy63b26hM42Hd9zr07MM
FjTPvNrndRMhy12pPJoaUZ305B2RFKkNAeBEM5RH3kSOm3BUEhKHqchrQ200reex
sxlhvmdswH5EFuP6enUriFTq6ZXdNU+x1l30NRKMF3I8XMJ4wdWJ6a+mHKHBRvtM
vClc8406UKt3llSqqtVd3Nb71tTUW08QZNjK0pZxycnYE6HiBw6BT4Y46jwe+/nX
i1lGB88SG+0RByHGfSlQSdVLFQGLPcwaxWUg3Sumtw31JGZw7PvL95c1X584OclN
0gr85CCsM/S2USvfy7VYckQdyy9cVrpfDVxKOyV792hA1CglEmRpyNllQAoavhgi
TnQH/CSh91IMdzFTb8SsAaeuzdckWv1Kl16jfHBJthsH/LxUM8+HSp0eyd9rvX8V
JHiti/45re4979zLkcbPTAmTmZgWH8gs3OUTVUFPowgalG4OEe5+XjzixNQqhsun
q91rs3I7on29o2659Ea2/GlpA2e+zPqVkNA8aNeHdmwE9Q1md+0nN/6qIjAt8iNY
oUVZ86tNKjKZ4VZGUMtWPkmbG9ZCkPTywhtF8hRKTfL3iZcTrPiX4yNLrZriwfLu
SyaDv+v3mxyM1P/wvxqG+OuK9kpSl20XRwwkKXzoPhG1hl7sDjheQhIv7U4Q+xJP
3F8G2YZU2ESKrAehZkjsULl9u1vBi6FR/E7kpg0pX7pGMH4HXZJ4Rt8f2RuQEVpD
K3IkpIgA6FhQf3LOCDsyXZzwUPQgxQMHigwyj2rDUM5Aceuf8kHziTz+woIt1BCz
NfGF6SXRnpsVEtdkVGZsxtK/9VMW2VRzENospssA+A+ac1qzq2QOaKIbPjFA/MPe
6aNIPWM2kPWl49htjY1n3NKMnB/yO53qULH97iJP/1P8prXldknB23U5B0tEWSFH
ZEbuci72Trqo49MB5n27sUQiuMM43tTvkMZ0vtxpkdX8WpYByLNHwFGJ++QoiBcF
0LYGwv+u1PwAlfT2D79DG33f6OqOWPeynKDLglPv2EWzn72fCuUZb6oIFoW6tIcr
tcx0ZKXoIxl08/5frRVblh+2BAEd0nuwkLIGHUG5rQPln7aVJE9UKfHqPqedOt0y
fx7qVSZ3NS8jH+GUEWfBhwamp8c9tebJq0c8gIfk0oXd8UwqTYeQaOrkzGzQYKQS
f0T11Vb7LLLx5Qn4/RDEj2HlgLvAus87n8a7hiu/SeXnpXEGZb+GUKFnQOWkub0h
ZrZJQoBNLbJhJtxS/BuCpWCufGLAwLEVFfoqeSHgDuG+aTyahJbZ6+4X6dU25+1r
P1Af9qQQVS+6BS4zOZRr2KCV472jlaBgTlXSn7XoRAJk9fqv/fWGsjeONsJCLEvs
ItgD3CEUce9m1FRBl9NrlsooVmXivm8QInaMLzHs18GcSj4ImExAU3fE4Yd8UJEL
1kw8xH6U2TIPqSo5PDntMIiJHHrXlCvKvn7TE1uVqhD3qYLoVoboia8u/P22wNPL
EY+0UdiFYV0yr05ddas+JjmnVpYiquHIL2La+BvcNi5ckeHsYrTRWxJUNcN593M0
FFhx57knBCigbeoQ4faaLU2+n4zsnuFz239MMSy65tiS2ZwUCdtUG1tIwWUfZMUC
aYz+aTa2aVi8v62X88XotYpoPVTTOQaGNCGhL5+RKM8XYGncfJHhBTEDyNugokFs
2ep9m5jwG7tl0tyfYRIySo3iS8aBwtSbev0iQKYttUKV4HSU2KySEk1v8Li4XP8G
E4syc2TEClUVGMJTqXi7Aj+Pw48nfyQ4pZ4HzVfTI2xUIbfCwRzkakWB6brzFHs6
Ow53rJu/FySp/R5DnCYlyPAQWOykq6WUE5WG8OFBDcrMYIAUZ0GL9VrbNV08upCz
OjQQrTMfavXPS+ITHeHwZ3K/wXFYZ4x+RjQgZcr7G08i/BOOph6BW682dcICsVQF
/TtPoTdobgD+1+XcIwUWVtyzYbjceAnPAIZ8X72YGquWkkr5fheRjOS0/NkY9GBX
bM87x1kIDVSEjnG/GsL6M/53BpaDPvaWR9Iyhk7v+r7NxEWBtT8DIrEzoQgm9mKn
6ISn+5AKa/9UajA3DqwPvBbrvC1E17e7m8pkeObm00Ib2eWuBAvjz7Wj9/frMa19
E073ydpGRDdE31YiVt+GJ76mwDIe9ABBXB03zLsBmlL4p2dAHSGIktuPytaN1i3q
29wjZeqVYSjwzZAoajTCA8SsgJ6Y+Pkij/Ubuc/AkBxDabOZwTXMOer9rL6AJR9c
rgbeLaNqr7x1j0PQ6+vOLeLswQTtOQ95L2aW9k27fTlSBG1SBA7c6Bm8GZGpzIoo
IXWmnRxIOPbNBipkEokYhDAIACXhAvHfwm/cErqQGfQ6TSVv9lj6RKNS1RLz33/y
oKmwsbxt1nan2J6IPWxk28Q8E4dsejGrCgDBJHJE8WAYAtWYTmzZaihMwyWgTsca
hbQQMn+6OxrLBO/x3T0n9JCAchE5GbyVk1Xo1RIy+jCOasxv6XOa0QWW4M4zoRyf
XmHbvjmNV/WCzRsm93nPcyuX/aCmLecALw1EtlDo+YuKcqnmzeitCdVrtaG3zvYi
DDL0+HASBDUOu+PHKtoMwWDsFF92DJQ4r+whdtnP7QylTSi3f61t6H3yd2ZpMrNL
HDkHtL75VPHg/yvl5xiPOiOyrOt32DLffU/AI3eYjwJM/KulChxjrmTCKbE2ppkx
EyBSyIEtPbBqMX3/R7lnzO0vUeKU1WD2Bz/dQG+LDGIaMt4jBP6j4VLo2yDjUT/3
V+fqU4F5emC1RVnv9kwSzvfryAxZJirgASusSilpX+ndB/WpX+lcyd1EHBYNqcxZ
2pKAp68aGIKtyDqRny3fZapxlEQx17HpCYqUOtQwmm0vU6A0o+ligqULfWQLjkP0
Y348aLmzCC7Qp1J6StrCC1RU4Y0bAZsWbsMUO09z/bWf6aC44UOJLcGdJmVmG7Vp
Q/CDVblbFyti0iP0D6rRIEUKXR+6BWTB7ZuKOXUSTqlFcUyl9zXgFZHK25iW7zFX
2abGjmyJ65u3m+JPPH2l3sUgNVrvfsvNlYBGsy7jfr6x9M7LCn0VA7iBuY5qASrE
ePsrRprAu+NMvOL1IuQ33qBLP0WW878lHjvgoyFs6QjVzbKbra0EITEKL7falws/
nbjV+0xYAcPFSQPBrY4ER1lks0vgTayvHRKBrHBFYQjsza2dpNwx8ZrPO8CAstX7
++3DuogAR9+1GF8I5lYNMtLdzI8c4CscneS4PbUXUuPdMIk8lBtSZ7ayHbv/w6wv
kJ7OaJqCxUqma7H866QCx98QBJXaBvUwraUIowdv+LSMUfDgcTlnjTWsMQU6hT+g
E/ttaP0FGzbvTtA81Y/UF4nTDPUTFQS+6PZLC8PLy2fhwFfMD9zCKIN1r42QUwJB
aPT0NLmTARizDPPf+YvH1c1fn6pk3UrqR8dTBWxqpLX65BSbN3b6WguktPglhYnM
JnS1jPn5GAv32R0micU9udE4Bs9CJTs6K8XecApUUNBepQn2eZNBsjsjge1foEiZ
SV5Ncfismzp8vCVBpgol4KWh1K/9un+JO1bqAZtseCX7oeN1toVN3AfbOr8yqi0C
ps6XUSXXDtTXzxyLppkGKVEQx6DwAhOcKRETp3/mr7zZXUEpEYQMv4ZHDSF+hMPL
hx2yZoytHAGqvCT5aFKCbjXgrioxX9THTC+OeX0J03MJ7IZrCbWNbCJSt8oBXNB7
vLG4WIZ8+gOa76IXcd1W1gcpTrgYZrL/z5y881Yn2p5BJevr0llutC9FmjzFrJZG
WxzD15fkg59i5pK79YOjQw2ds71MK77WNqvvSpstpQQMCboHD9AsUaAxcxR4UZBH
YTe5yvKZ5Mi+752agf1uKi3f0Wg6yqsFPVcMJSAvuuQaoaUcOfKzIrlUMF4d4Hav
+9Rijv3xlR8Xa/a+uhiQSroLqYefP/lzkI7yAqWT2KFmFy3Kl0a6pZlvCF5tOBOj
8XwvXhvJrv0YrAxMkCa3iI+A+dOGaI04MEreTwsI9y68xbXWxF7vAaZ5ffUUzfvZ
jlJdovwqaqIOAxFTzWiPg/RebV4/A42D+tjSJ0vFmcyRAbX13RbhOOO3N/cyUaya
qRfBBAZ6uPq12YmwU4xb4rcER2M+e+SYNHm4n1nBviiL0FX4F+4TRjrEFkAw+jyk
FS0+CltqhUJ8Kea/d6wwhpwNUzN24cSFnkzJZhY4d1wDukoMX4EkerwZ6zF2dfAh
R8fHiBY+AGhbsvrtRBMYERKZI/Ks9FM7Z0slUuTQCQdGbM1oGYz2zgiHzwt3eR7o
AlBj6QJpehtfPDlpSMK7nPvzVBCNdWyCKtLBxDCV8D11Buwdi5W1I7VnlZOj7hCi
cTY27GJVYi+a7mliRvSvdUYLFH03/t0m/edRpsrlAIQP19CzYxnQ26m8iDOTj6Pk
mjjJqrZ6Uy+pwPKCe3bV5CrXzuj0QaO9QF2c3VHnnQLZFiZRpTn1HTQMmnc47mme
z25f/XevDnsl4rZ5wu2ztw1QJxFgxSwij8Kj9P12tBsN9xCPQmlAlx5c+46XxQPC
Gl3e7pPbxDozxUNGiwS4oax6S84Zpp2cZ9q8i8f2A9BMw1ePKgIhq+V4ocCc5Wlm
6J5gtYFMO9OjqlLlS97ljsvzWg0xhA+sCmSw1M512uExzzqU7E8SHWsQduoDWtzL
40Y5D3QP6bm9aCWv9aXr2GgSkXiUnY53MRP3JD6M3JGAlht3McuK49DO08qGJy1D
KUVlwcBjZI2dYb4nmC/j2+6NPTKmkYjHtWpk1qWBoSfKsWHwrhFZnEMU5vG9vBxB
nH7ON5mSZCHPhnVmWFnW2aZz1aaXl5TFQuGpbHcO/mEGCIrDXoNXKOgISL3WM5O5
VOmcciA+i/gMo8RGg+zbRbko7OwCQJQEYkUCo8XH7GSi9UX2wdlj+mDjW/PNysri
83nIyDut0ulPohC4Azs5R2B2vHPAqdZZE3GMWh/nhlNqMAKwxkSRJwnesksgmhy/
GtC6+PkmDRXdpcvDE/XT/wdq9drBQ1EW2BjpRgEmGEkpHjNTfjdy7gb0/S5JGLmJ
BNNBUMTytGtAn54WQPb/QthDLubBTSF4D9lCvGGK3f2AdOdRKdhWKHV1RXlYaYnf
OTp0MyD40aLdaOpXFe6oiQL/GwHFnB92WKVnasxtJB6Bw5dJKJZLbjIVbiRSpvo+
8riVEXDXAupBz1mHnl0O9X2pMdjZ5wUFQp7hJPvjHhSlR0U4Xg3j6R6B1sIawAp4
QYmAnaoZPyuL5IkTUd5X+QX93WMoKF/nTFeeiDGeHiByTc72J5v4qGlXB3yy8R/N
VzMMdsEZNWA+PyAwpNfFlB2XqQ2+mDfRwWdD6sGeIPcmt1wpl39NPyFNs5K5cd2v
eCXeX1GHLNhFK9uNHI6intu0Um9SDfQEI9BMN/jf4JyQ+G6/fGkmsDcuwq6MlY+8
p+iI04l7HQ4Qnf82RF8dyIi2abXAKR7g0dG7uoUG2uVGGcA/Kg2TW9iMMUgBXauO
RfBEPRoXK8oA+/W9H5IhhDQcubspOpKXGcXZUvZMOSOxX+p8f0rn3VCnNNsOZRje
5eHDUDKe6Ztu1neXRoBJljoGpJKm7p+Jbw2hgqkHNCvhPxLuClVe1JWbSs1vOqsw
h8WcJlG9pyo9NSYbsMqxj1d65k7qZYRmfSGtH+SZVG2gmDYNhJkIR5xFW7TAbldx
7q//3UpmjN0GpBLKJXK6BVWk9L3CJQB4NKBoGhwoo6Jv6IuhYjUa+rGXGEo7qJcP
pC19qI7F9DrMu+tMYEDu4s/54QMIue16ciJQLc/AaIYwAFKqHuUV18MY12yMvoLw
i2SjYMM9Yax2t9r74hqzkPpal9xBlGLfx0Ve/QKO1c0+0g9IijPPoMhMTyyV+L7+
BXnQqFlISVuSmC8BN/yRAdhhbrkyvxtJG/+84o2oQ0aoG0hHCC91cEvnn0hziJhO
jgCEvBHFCM/I2/ybM4f+Af3brkAgw0A7RpyIXn+4KLBrIcnktDQ4T5qfUtUKTYc4
99SA5XjpJiLLoxyTRwuvuiGpYAB933KMqh2Etw+V04fGkcAvJT+vhy0VvkLvFdm1
GfJNs35DUYVyoOXISlg66yMya7R6z4zT/mzkXxKv22FA+FplhCGfkQsMmFUiBaJ7
8GHHy1i+Xg6hLJEkT9+lTUVZK/a/QuwgCJm5fPHC4vGmbAWetGM6pmvqcGIbIXVW
Zzm/MKR9wNEQtFZA/Lh31+i8wVG03xG3PqnvJ12L8UPXmIRpLn89rJOG8vEIOCIb
kiNKw3JpSUbA8bomiRuWIoQc1uCygDMxHRDCt/PVMq4cJ82dl63eYZuWHHfZ/Bcl
aCZrgtk6Ik/k0fdBmMYhjeJGhQW1T5p2xS9L7Tomhs+rGRShVqkwoB9rOQ9YWQrA
uPJug/QLzHlCBgeBYf7wxnqosUFMAcJrwUCSsrWIZeYh6+OhsSDQ6FtdIdhwa+TB
HhucY2goA+BIqF5kU2thwKzl8roRLNyJ0y3JcIKC+yoPL/XHAYQ5GTHQXIRwL6wU
isL4/1f+sRHUi7T/pCovPy64yYa+mlWZoRNP1qYCbCtt3bGjmI1n/g29iyA7Jnd9
txqO2fcOJKrkF8rS7ZCn0nc/z5X9bgOQ2fVgxKTFMUjQ+//BE7fk7s2a50XWnRvw
fNOfR3/boTQxb0aHXGVehcOfahZpJZOeAfyi0DvS6moa8iBrHuKHqlO5qflA59az
BzSvyEmRl+XZQxGOz/68vlj2Fbjil1j9lEUuI35+vvJ8iLP+TUcK4kgNtXyHaUAZ
ikFXZulBpA2Eu2VzmS6y1TijeJqYEFhw6x3L133ndQDK3Hm4O4uh5zLyy6PcGsT1
3II/yNn4MwM7n0k2ucaQdqG32TfCKQVsc6TCW11i7FPAMAWdVOwPR4HPY6b18ZYy
eBYjvPes8GI6MSHKRq4ctEROao5Zw6GwMIGjlKu+dmC+OsUvbAAj8yIadoMPN7Op
kowl7c5v6jjnIOZUU49Rn4xaPuT5+KMf6aCfwY/IqIGJdYdE6zsWh12B3OdSRakx
FbPRy2pOWReyWlQ2gM4x6LQKBzOtqgVcEboPrn8b18Fp9pAK2CUTdat5ij+N/HCX
6MW5+6Ra2MLUIRNTFopH80zKbo1V0akE9qUfOluHf8Da9TJHNGWeoalzOzHn9zEK
uiJSsUFyL1X6s4mSGdfAaEwJxuxI0mBcWDNXsJ/rrcww36S8L1NMiAH/Udn3xZdc
/r2KyKXJYnDv4laSwCwGQsSR8nLQ1vzVYo8/168yjdgKIinQYBWKjh+DXlBJ7GkO
5zdyg2wIKzrI5tX/lcfqa8+VYOCeaq6ctx1QgfstmuTXJUBGAlARi1YMzKQDpm4F
tl74ljwaSQwAyO1IQDGTYPL4mirX100N/H6UITvsPIQjfAVzoMj9jj8lx6txRIKq
i5QNX3bmlmOZgk+2eO90bfTMjV9muqFRnADFu+d7GewmQant59DIsd2v8qLiu+5c
SUNMKnN9wOXrjwsg5o/B6gX11Hjj8N1nO6b4I5juXUVgPd6d0jxT3ALDVVPZrCcM
26NmHvn2cFP5v8oB5NU0qUFOj8U2yYRo7NqLgg3mQcm225p8jV2nXS64G9dIuxn7
pXImtvCizV1bB4HukK5OeLyTWQ2YkEYYVKaPgjqf8nCA7BZr6JNgqJqFGz8940cy
dSA6BBduxXy0K3m7/9mZ+fZbEo5AhpkbOIg6U3nxlQQlXBwRIsCtY8w3+86CJ2FE
/fbm0E43G1vT2JouOuRY0/EVq95Az3Sd6yHXRASO1h+68qD1gb25tbPt0YzghCnI
URh+5GgtoKOj2AJyUzk4uBZ3sMnTLHx45lgqKtgThFSgM9gvZwCmjZdtRKBttImm
MJiD+mgvqwR2fiYXsVeYM+cBrHHBTYHeQ/M2ehNy/A6mQmGAqDGMQ8FNc4NHQ549
o+n1kI2U77ZRPP2uA9yDDYA/ZhjLf8YLGFaezxhnmL9jGcg+7rPQnFuX+r9oYMZ0
KgxmCbaSyVtfejAFxrHcBot8Daz83UqDiRHHtu+0JeQZwlfVxK2ttag86TXcR6rZ
0Jj/Ldt4YiD63sifj+ur8TlHBRN50BkjXHpHu8WKMFIpal72c9DjuJ6krVV8kFNG
zkzpixPqaCNnhMjNqpm2kh01Uy4rElhOijlTX7zMsuGp7s8dybUFshHHW6NkxeOT
8/HveubKdxHvvg+sU7aqpNTov8GkJeANJs3Cgb1FhvAbu78YEYtTsPaB+WbREiDa
ySqopcf09HddU5mkqIf+WcVcYwSY8WaclzcK7TqdTkmeBHi9daxuj16UsAcJ9Ktd
LwlcGuR6zAhZSbhuzvU5offNazHo0buAb5W9TQhofFm+7fGMKWwj/cujiBSNIUtf
xL0cFXamoIoquN5mTVj8y+JDKw0ZxAWIaJp/U7WkmPlrrgARCGcCPd9kll6deIgZ
+kW8OmKk/zZ8hdCoN5+Cdbea/dRYTkxxQRjPcIMiMrTCs9+yK8NF25t5ryUZSeRo
dN0L8XWHj1emkW539Ni5BSMIqkLE36vblZZ9YJ8CFheFo0nzsM/qAZzS3iqbjvo+
iE1LGZfRt23CUluOEXm8Cay2yf0OXUlbwMf4/XEquZcHvnUxvIjqnzoJsh19OlQ2
Qg6KRZbwwjZnFva2ZueQ6zsgvPqe7aZeDGoDmPD/bX1LKioKXN1ZNZ4Fvktjz9iF
qbCEBAZ5IHXR17TGuXZkZR+7vQ9VselfnmVXwaP5xeNk4ebtPPqhC8CYAe+9mWJe
598FO6hb64rFuOnrQm9ObzkkgBj4Chr6tCmFV2YXhScYgjsWPhTcCvbCy+5Lr/pb
TuR8Q0qrWH4UlUJBl1DpUD8/+uyaTNh0PbL29UKhtLyrqqNSHtFqoJiXBAGnREBN
CmwGCmkF9zYaZbdYnWWjumEcw5xX8ygROAPqGnLl284FX4501kfTRfoutLazMApG
rZd/RlA/fwxi6fU//W6BZDv94yw/h/o9GaZpAl4VayznuQzOAmTYsmZz0K64/RZF
oXcsVrhPZIEeCXKGu0UpWgn5d5ANrnFz/3OrgYktuTxHJf27KBZSDRc4xQNL15L+
gwacDmEHW1+tgQwSZ9nqZmbU88/IDN8rlEV8o9412BmEGIeRyWrHlrj5sELd6rhq
7nSCF5dlvtCMBzsrxc44Dpw5LSk/blSIK7J5KgepPWqN3rJFYgp8P8X/E9H7VmEW
qXMb/3h73fovky+HYt9e4Gk3yVQdz5O/jdkDN/885Ps6tc46SmD9oQGH2FAQiXnT
ZlS7IEmiwnYvV1mqkI5qtYtQzOM4D0jKU0VIJECa/UWKoYqSdlQBDcU96tqSt09v
emkcgFmdL2JmXqrf46tDTJr0wJhvGJ5CAscFzWnPOYswEAsKk94Obax6AmSLHlOO
Gjiz22RJtYs6KZpLhDgCx0trHFCQBaCPNGMRQ2e5bKbFFT93d0eLF3BT6uXRug3b
vAGZceKQPSpWY+s6DmULXl/+aOBXdH/tpLyWbCuwBV1S6WL9fM4NtApuBwbLhkjR
A9co8AyUpEKFUGNaCGcyVCvVWO2AMtKmR/xX50Qj1+PCRVFp2hPB52Cc6/LThpQR
nne3jjf0fIL9ySxZR1cCWUTwFCYDZrylSa85/diYhFMC0B9Flj8cSFYrQlQ8EIfW
IWctUZseF2xaXKCYfXINbEPL8NUr+yfoEVM2tb9K7axhm3vyldNTqcDVuav+Y0BZ
iTCRQT+kZWNJLVFb7f32O5REN+u/giJh5ahv7BliCP0fNPxLL43eKCgEspF7IFRQ
P3mifTAl3lpIPaUCqmaKZS3ILSgd/xHo7emgrXrZavGMo3iY7lAuyYMRGLS25ajv
JYe5V0iUuIVaWRX73uMVYOsDM4wpN0yt/qzq9D4GkbVUfTdJwR6iorPl9kUspr4w
BmG9eH4DbSdMlV8STyoVwGKlMxDPH70LT2viIybPf/nx4hEux7P0wWcEvacINoSb
5VXiGHkkNTpEco1gmpqoxvVQMPIUfT8jzVPCIRvC1s+VnyeN0qXXgk0gEZG+Xfc4
NNri6+lKqMS1HCTMwM420uzoxsYzvNzZoMLocJZI68jy+FN5i0n6gVrOHTYypllR
Q90KdFMVYvD4wG6wPPYWpVUPzApzJ9s8nEzTuROAlEqFTT35yk7InW7Cd/Gw5Mqm
r4hCUhYvS+MnollNLjEQ0AtP0l3Di5QHJNp075z1O8YZxDxWK+rqfnxSMWG5QqyB
dBQ6PWpvmx2YQcNLULGgCTzCN4MawVQuZ6jXbZNbu9qg/JOtWYhPW8F+w7etQEI0
JztLtZynmfBB6AQrGLQRff4v40l20uEMDMKW3oPP3mESOjVjdaZ64TKC4gwxCjJy
0n0ixXLJmfRR6QX9OX1Na2ULZfkHwPgce4EQ89mBS9eZXAfHpstV/U4BojUWma49
b0YsEX+gUjp0UESBAxGVi5OjpbQGAzw95I/MHOc7o4ufS2FmpKJP47ANr87cqneZ
cR4/8Zq8BTo2L5QwR65YOjZQ+FVTiXlGwf7Y91k65+jgrIu/TvQKWfrv1Lkw61mh
b7w5DpfpBFM1yRIgf1Q89NBiLxraB7WVVAHH/ULspnsWPlylbRPyh1e/UNMndf/4
GDkncu/wlT8o2je1u5iwCMPl8jtKNGNdlYRyTFJGJFy+dkw5DCaDtjW1oDdmEVTs
pD3JS7pbyfTO/KgleJ0bvEdFyy3BO/Ujsx8So2hBwbqbqmc95xjTkWKaRVcz23/A
INOGynPkrJMbMx2lLHOZl3KqZ4gU0gdQ1KemKnwdyXFJxqUYaIQPEIR1Pz5goS1f
JllGUkzkqsd41JrIK85pEFvL7JUMw92yel1C+7nmVSanChKHGEUe2GVBbMYaquyF
dX8EPbwe5HlLTXwYQ2e556CJkNiGLmMWqSN2Lg/BtLzbRF+vmsOTWnLC2ssngoXh
1rRgxAohbxMZtel0WqoJyU+2A04Vr7j6esIUcCbOSqhjuquLcNapslxXp/fcIsfO
E02ZsOuUX7GBb9w/kju74829lm2+3bFwaXttU2oAyX8rgDCdyhMV5GD9bc5+ncoj
9ImKAJt88AitVqjS011eANsj6a1GuHGdWvtzXn4tF/PmO8wioEvXPiycXdfQb10k
PPRkVweL6306zsKNv70B+JBDN3uGDxfGl8u5xWIjVMyFgbDmRMPIhkUMw29g0wR1
4JGObOKHXJrxjL4rFl37TqRSDDRV+QmEscx7UHdTWcJEFh1mgUloCB1XO9LEQs+n
XkySCj6cK3tFNrhnUrt7ynoQrH2p3qvGSHjpF3Q6NVDZckDNKE7L0ILMmFLjHdbo
0eolw2oS2lLDZfV8wp8Rnj7X3cYDbWMnV2UoBMcdPLCTvdhehbDFs2fBbj5wxZH0
1AZxksoWjjw002pcLAR6PEdIMQrqRgDue6McnU9W6uJMNrtE36Izy8hUlwAIJ0YG
rQob8AZZWVmQNyAnQcgTO7MJolB8aok14KYrHk0c+I//bTr4F83KPsleJU9GRJdr
qfgzsMKbHzX7VTY82BKLmUqBdbhxAmskmh85W4JpwitTZw5FXNwJ/bZwl0w/uCQ7
FS5K2aiIYYrxLU5+x6tCr+JuCW5Pim1A8NxYUhybG2Z1BuB524bEtFucqHuBUCgX
Ct9QlS5L+5q/mvF8u/TMye7WRNyaS1JShCJs3jUS301QdMstpJeP0k9CY6z5+yGl
/EWn/X75vN9PPAavPtn8TZrl0UtC4nt3pFTKeT+oaB3AqVDHOR8x34457pdQ8+Tt
xu9KSkawvg2a2hOJI0ieEv4i/fZ9U2/G39yzRcpFiek9oqgxQbcha+iBJ5OVf62o
Lfg2DoG9DGG+4Vj8hin5LE2T83TJdPw/B8qfQZ8G8EZ2nIvUBjvnHFJ9YBRCMqaq
sQaYitcO62phQl/bjfoA2/+XIdn5ys+XjM856mlpDWKUZASYD7MTaq9SqR8qIUyC
ZcD9Ul/Fps/R5WgarOVMpgWH5PSFVl1yjpAXVyyiKkSU5UZjMjUdkPpojJSqwK2m
cacpB55LyW8Cr7Rmc93eik25xeqJYF6FBBFrF2Fv+VlGa7o9fj97NcTL6ZUfQW2M
d09OF4DrAZ4BlLC1ZgJeR84o/0xT/4Gq8QeuWYEwdlf3Oq7b3SuWuc7fVAeHM7V9
lynTQGiufSPcl/vXedSmE2bFvgAZvnRJlYLdeTSbiuY9a8bQuZ8yrxub4NtmmxOm
OCmQ5CQNsB+k9a77LRvYyc9g3NcHYkxGU4QXMdeIm4hYI0Mrv3vI2TpLOxP0lLg5
9+1ejxP8Xx/NxdU3vQ/YLs4t8apXAqiucg+8bddzZCsCmT/7R2vzp96NZNh9QbL7
6xczvziy/CGWTsEOBuzjUZV/6lPEMdhd9lmRGeqFILPnCWbutVFcIeJVOENQSyxI
gmHM/UoB+B0PrYKoOQx5wlgW6KrIJRmEw2TxaBmFRg61VI51PY++QNOW9kIE04Op
e1PBO/8xuh2jTAeCAlT/uw2Sj1mqZAzufvXh3uqZxCydP5hW+i7n2QYgqKU9v1+9
zE5KZsu8EQTGTx3wxQLmATSgGHThj3PG70CTsLUmpAjxp4TLdsWN+F0DlTI+HoPU
VztiWHwvcg8K9tzqbKY6MFuKiw/yDXs8DsOKi23ajbKukoaKKAtfoHeq2jnYKUWy
UQJMJ4CabKAk1DYFQLzAUq+lI7ILtz1JLGxLAKBxrjBNRrnoEMCNwCaRdWnIRcMS
2dnJANFL6sp8xSTqDtT/H/N4cYbKQkAQtuigs+gj6Pk75Ske4N0eaPUiSy6+C6RW
U98FZPFKXYlbtF3X0d4MsKDw7clavzCNKBIdve2TzZ5yUTmOyRdWKByhtrzpIDPN
v7Y52kaAFn4n7BWrgDdsU2Jil8856jZaRyFhj/3in0fxH5Hextd6FiR/LMPsius9
BMo6WGY5yzxl5dy3WjuondRdqJZYsa9R5y4o2rPb6VVVYxpM2KIUZXqj79qYrxqy
uhn2WOMdal0418N6AdncY1BrfMsIBCL/stKZQEJ2SH4nUVqAGnbl7D9r3GK7E6XJ
ReZiWk4ByKbizKl5AHjlAAv8HP0Ias9WJtsS+yDAiAPG6mJaJUofSzILJI2iw5tG
5BlsVx5tuM788SxYqjJO8MDz9hLz3dqmwwPpS1l643sYp/sjMpaZyv/aI+5J6WXc
xhn3OIrQNYrJbzXgtXv7ujDk7837Z2NQwW1VoNok9k/jTvHJHrLmsDwP7sp1i4Dz
mnpOBNcslm68VBL3aSLYy5UaxrcZq6SJHeHeTVHHl0jENH7EZNDT/Q0t6k2b6sgH
2yuSdcX3fcGFQTmdbPaJyV+PAZrMeaxuCZjGqH32w4Bba1xk5J6uIfrCFqf11Du1
cbVnEnFtt/0rfC/BaMzRYmFW93ApxBMws8PWyCEI+85pbmds4Y7M5efUrw5rNZzr
4d7BWn0a9FnIBBtog7x4i01qpZFoye5x/7p8Z54YbEE3RjLq0mNKQjgygRGlzwk/
BbK7Xxt138TNom/IjytuMk5K/DDAnyOoHJRX+AMo1ZT/pImHcTSt7TDb+pkBIl7Y
gTFbOko5Su4suYLATN8MoKkz4bfZOoXbAn29FdsKSYcw5zBcbEGNwtKy1NYDS4YK
6KMf2ukAieIjALz7L9Q/zXTeD3y8m/veaOuwa8zxFMyV1vKK+8fdwRnQ2Fe2StMp
3HZCfx6DHr9f3l78hn1swsvA3tZI0H+/QC6oZ21Jstg8iGDQ4Hr2HZR/Hk4WbYlL
7/Cvvu7HwX+pPrI8LGNCUZFWSmKP77QZG/I9Uruf83pEnHY3OESZ47Ak0l8aA18S
YKPR31lLbjML/CabYdltadaWdz03tICM7M8Uvuxu+HFEIgC2GtsH71x9WFEN5kvE
BHaBQ+C9r3bMWQCkYFzBZ2+UXtoi9mcIvKda/ChTTPT8/GT6Jp045BbFqyvecA91
4TRbN9wb5sNzFuOwBdLlBxyiN5gc940Btvvf/KnjlMND5hmgqmgN/sLToQo9OATD
4tfIDJyz75D0qa/f10QDB9raTC0dqRpdYojWuE7vgB7tUCBwfEWRJj1nyfqcxgbs
ZD1CNdFCsAlDBz4fv2kBlPdApzcfhBL+nq0OPijLNm76jFpIML6tpijs+PNJUKCP
GaoXlR5xrirZs/uxEDazLc3BnPZr79x378fE9APtg8TqYWhWyVeQ47gybHYNMJQ0
NXe6IOnIJFlfL/wjZRotgU/kOymw69cHtqlJ+L4zzM3DbTb5qHHEokMWXe8PrWwg
glqLESJ4WnKdpcGAz4gVY/TvkgBxkCaNnQ53HqX68tmJMh/qzVsQNZWq5X04DRJj
B7PxaYPD98KrfyTvk/x5qNRJn2jfmg7FVyAiO0Gj5M8CDjq4pjmIBUTTlR+CpIKu
KRCwf32DhiLCVOGS/W4ayVI2y2TmgYTNrr79N5vXFPlSzdns2CO6bJ4hna5ZbL4Z
aw9j37x0c0Dlev07LhzXoqdUG4BzCqp2js55b4lXBrDBAgzs4mmwojHQys7bgbVv
p5H1XT+CJ17o6cKqZI8nK+ib4zSnOs+VXClaiCSMpMRhUGuqekEvKDtAXB/CM57A
Qf37yMw/wEpCfXLtftEQ/H/juJewfBtQIbBGz1qPbo/CKOjZidD3tG283+r0XowB
e2sbRuuzVGBZ5Jf+iUnNPnx9Q4n5OQ8x9urLq9sFtolB9wVYmjv4WiDczYcWvpni
wjV8uoU+uvgoZU412/I6X9+IhJLnVCD8eKaMqluSZmOq4say6UWhsWUA2V3fZySE
FdG01WTyFkIQ8MBdXW7Q/P5d0sAV64wjHKR7iDbBx+cxBml9Zvz2RjA+l7fFr8MX
4fGuRQkv674aIxAM1L3s2gYxcn8g5cvEXtaKwCsIPJlK9b+9Gl8AxsVtVm+lwU3s
JHn2lHNiEW513glcfIn1V26It7Pg9/+Budjnz1wEuY016b+JinbqUGmtQr3uds5J
2XWAKmba+/aNEMlE8R5682WBkp50MtH8/k61t+hrW0H64aVk+JUzEgWZ8H0Iaksd
Nrcwe3ExwJMPeebwVjfIz4mf+r04kaMztAglk1pFYzzYYKX/vbwz1ufmoMxPGKgj
7rDNwPT+p9XpvAhY1czVB6PvVUJgOiC966DfSyntPdy2Apg3ledv8Vin3tJP59no
RhE1oAOJTOqY9wfVK0IjULwOfSxiMW9GAhf92miXfiukI8MlADW1/eYiXwowtao/
mzrqYUZ17N3HMdWqGiqs7wvV7/jLPigJAxyBys/KMFcF/zZcd04wZbhJjrHt4xtu
snh2RON5DrfxhW1ugFDjmac3kSHxYqATZSjmp8nr7plrlfto9PDM7K9VO7qxFvPj
PeSnOUkPmM6ohtwguozFBP+cvToAj97oWvrdwlHWwzdUbeUT8THGHXUW2x5R38hu
JINcGumlrZGYT+Ijx/ymWgicPYmcc/Akh9d2b1vjqQhXXC9L5hyZqMRpALLx4Lvp
oPDQEGzW++UhACM36JsuzYUaCcT0t+8gRll+5yzRx317seFpOVUvUQP7ol+x+cOg
ovA0VbLLvekSanmhsd3DTfhavD4coYHxBFjHB/v0g7nDYIC93Nd28F9Wu7o0lYE6
hgvuzmBcz3GgxNOZ0lrXtW/CcKgTaUAxATtH+zUi7nm1hiJ1MQBjV9+dCEPDZOa4
cSEWIwShUGRfpqte4qq7TSN6efz+K+dZto5Iug6a4ZNE7/mUBpL7yESROfmglXCR
j+DjSvlnd7J/eMGGVDd0PW5Dpsp7L5SSLyMpXKURfxYaobJ6Z/mKnFmOVXHhgxAy
Fq79QUb/avS1vJFr70Xne3uV9B7nc2rdS7IgAZWmCbPMjcK3IGxHZ/xlXw1loOmr
1oPvmRILM5IiP9KWbpvshr0hraB0Qq2c+wJObS1qK3vKmEtxrZQoSi6tsR5eGxjm
/1TNwhiNk9HrI+3UdgA4x9GID+Ilka8qDOQmn/Zv6WgWNCZxavp/g3xbMkhQg0ky
WlGPUd/D5j2RwhyfLq1sB6JdicXanSxNRgwEe0VTbrsslZi4J/pIMzD4OtmHG0B6
091OX8xP8f/M0gaBzsP47aTsPxxLECvg8LII6dWzRu9wrCHsedAkdqvYFezPPx0E
dBj8DsXVi7kovMz7w725r1qvERpgXXQVqM9P/7vJxVhKTV7BUKoQSeY9sZHx4YXt
+BGsufzkxY7eJ+7d+WDEMXSmVtzHtcYRa6kj55GqKoyez0967OMDOujnxJUpXwr5
RB3UJvPklAj6cZfFMDo1XnGvtkH+XLOjztpI6sNsR+01r57Ec+mpvQ6Lh5IXwEry
nqpVGlN9RJKV7MdNSgc5dxVKv2zwMvB1bmMTQXrE1tFZg4eb3r/pwRdIxs0SUpNr
TR+JcQyjteIJOGFz7O+f+42N3FMoXWOXgpNswXRv7X3D2aXEQDyKiroqIrwfZg8n
1y7siriAagST9gaFw6Emt9m6SomqRi1RbLoLSsz8mxrk0RfMUTS4vuOoprePGxP6
lHaApFFCagHTo9eV5sBcR6MnyBP7HQu02l1c0wYBihVcHjQZXVOjLund95AUxlNB
pp4utqnINjw8JTgB1ScRIrqqQeq+8DfR1rFTimqLOz83K4v8mIUfipuKfs9nxlUl
VymgTu70bNpLuXY22LjgjadUnbM4oGeTnVVnGkLe+2tpa9WUBRV+BE0EetVPWQ5d
xFntpBzMaQfFWY1a9DQxckX2ZYAOUPnrk3OilQB8DPBWsgI9N0s6c4iqPo4S7n+C
hwQPEX5Azix5q5BsjtMR5p5NJj+7j1rCoCz2kckEbsFAg+i78O6F29xULbEruC2l
ihNIPa7ETIN2fQK28cf87gmP46+fssOQdbyUMgv4mxpKgTO0aXXdbMqIPKvfPm9l
sDnvuP1/GB0TrNNQH0+BIbDjiBtoCZMhlmP4Mwyf3IkbRK6f6KkojIDJMX/RDVTl
T9HZvhBAsVoF2D/psv3Olc9Mui9lwl3iLvQYfF+Nm6EDgyGAKzJTY8cnXqdWTp2I
9olKxkzO2SDfX6NWLP9xbtc8IDpzI+s7Ri2CGM/w3qVcfoD+pa0BwIzhTNOHLReJ
u+zcSf4JgqZFW8E7WL97+hSZTrDn3o0J74EMcQHqe0IUTvQKRQlo8wJTM99TPIei
yMU32C5/hGdaL9GvtWgBySyLgWLIBy/HzVJKRNNWGhfKEztvJRPy5LSwj0NERqhD
uyqvlE1Q3xqlTvdRu1NkjY+YGMAnNbmdbbSLEc+FNmIiCqNXN8ghsFkgzg8uKwtI
8frpJ6gEnp1DyjdF4tvuHU1/93wBb1IYRNFYI3Y2Ybst7U8buF1d86lybDXMfKdc
LsODWwaYPDSNWe1ob6er/e+KjhzhtisPRU7OYpzQ8cCwpVfWbwzVVxZgi3QEvuPW
k4QU8CHMwxsufkTH/ToMRCesGbmptDJcxxQymlJ5u1d/5cUv8D7fS7XV+xy44gP+
w7phrteUQCSAeazY543u2jb6+lVYRVVrFy7uYoop9UOkWumLWTLNCrTphJFBTFek
DDZkggCkUX6vnC+4t6CgHCbqxYY3uHFq9RPQ5wgoGvVQZBBYJhPFzNhG8gd+yBoj
VccNTYBKF5T8tXVelxDIiPcZsRGn1J9uZ8J1J2ShoshwztPdkvxMp0LN+AioOGY3
UuIqmQmc7oaLAJfauQXm3CzsO5CZb7YL2L+NA93gJfWNbaGWRFq/LzhpG+BT2bds
D5xdKTZwuXhJ20KAtZlnwvBgqLmc/luQ4i+/C3ln4FeZWDEdMhdZMj6PbwdgIC7j
RuaZkXjyrPCaIFBEndiKmRYGiHp40qNQqm+ye/3smU0bYzACjTybABSaDrf4b2QP
SqNA63FUjb0hXiVKajvkZBg1pjlR5w+eVIr8gfcRt8zxDiFh8QCU26HpbVQvBKPx
Pdugcb3+dl1yQTkFn8hndtds8871utx+mJsxhOlMbCNsjfLyviAwiS6Sk++73k9i
lJ9TudN2KnRQoPq41FeKg4D1ybI4CScBcqt0CPvp/RLFW2VZ4GBm2AyBm5hwjcaZ
XJqG08IFUCZTOUbzOtNZ2PLqq/TQ/7RiwGiP5MPbg6epXpv2qkN7YZKO2nLNck+t
8o/QVcSjUc1NtZrwyvUBO2empabfJa7JPVUZsFVVA6gi+md61DFte9a7l6SDlqZh
jFWanQ3ZogIZkDmDFmFD4weKfQa8YSe72FcfcXepN/il8qlsqRQHEymIcSl52r34
GfOI8ZQV8uIjldbXPxH2mGEbBgEFhrpHPqzgv/Z+LeWiH4JjtRNOkX78jHuClCrT
vJqecCshzeR7ruFu69mvLEbK70LWf8XYndgobbXyTSytI4QTvN/9Wp+/A1YlR/Bf
CEayrREIYCgTgFwpKWcLHTuKRDXZXSov8ykh611TyS/16P3qn0dZnTM2TajCJyiL
FBawSos+dN9uq+wZVchu2RneS9Nb586VCrHy0tfq39mgwF0oLniyde/qG+jQVW8/
E/PUIUhX/WJhpFq1s0sUHhg9GpL2ovJaD+SA7qd1TLUQWNOVcVSbObqk/EUWqOcG
iZ/onbjohSyn5RZXjSsZW7yDyQ4IPLj/aZuFGaxBTkKcZl9HATubz1WC+WBsLvTv
5MFR8zMIkuE8I9ucPo1LcRtsqBEPoJHyM9XPuIBR4FIeUUzRWN8Tj552eZwZEatg
P2lTnY9sLdB1OhrOkGTSZRaseK4EdzaWfWSUwYKzuGrxGnpBrMEQ4BWMREXfhQVb
UWJPoNy4eJz5fBKJpjCmD/71FaOF/X0ObuyM9G8vZWqocfcRx+UbL5JVm3T/K34R
I/OleokLUI7TJAy2x9UMfewcN2UuawbDChQsJRtjI/KWf0ZhVGpudca42MD34/VD
/Q4kwctq5ldDLDbSV9vgqflK/E9HpMDVBz5rqt2wBduaKOsvJPYBZs+5ygrHYCN/
YeF35QkfIniCPo5y7sNS7WI7LwACYLGxdLx+Hkdc7JDE1QM0Qra/jRrEYRhc65cW
bZcTYe9uru9MbfTkxakz0/5LiCeA0MHmzZi2ulwpVPne7CWzKxcFPYBA+9zLKg6v
NdJYiTnc6PtHAuvKxYoxGv4fbffvNCKA6rD094J08fIOhNlhPCnanBv8yUwFc/Qh
VsKXG8ilCIDE7Ek/wFtkbErMVMbrssg9SIp/RGp1H0jOkkWcf15sMuysseX2/Qjl
fxe2qBi2Tno1Yue0jbYv32oaWlIbS28N2+rbYLrPRcIhqkdTosAATJR6CeaoMtYC
b/9MdMgYg0faSO8WWt7hWl5N773akdYmGAPCCXnsXdnxkIXU4MRrEmsXWHngqrSO
KZtHr2vl3m8X1Xtctu/n6ODd+zuqtQC6iQUdcORI22UcBq82Pt1P2WHrP4x+cVsE
1ySmBtHf3nkqbusMao3WJK0kSdeetg7zjFZoP5mmAdCbAmiSPlGzwVMjdCTfLz95
9PFj6g+haGeGfEbB/XHrgTB8idAH9LAD1FtqrjBRr4zlFABbX9ISLle4+XhLMhBO
oSYEEf4kaqa3AZOBAECBxYSt4ycBXQU19Xe1smv0NY12+TjdddAE8lp+otDepzzD
9DvoljUCYsvDYLoR+wYUiA4S34MYGrKZNhe+IEKkmaWLDicKSl7Wh3wB4zFiyvUF
OmrQBd/YAjaJdAbauVr8VC6ZmmPUSvgb/n8RhSCybROyBscEt3UMiLK+njycl+m3
c5o7kHChUzMrR7CwbS+ywr1pmWC1Vg4XkjsbviNBpAkfsup78xlko12/n19Z+Kd0
SCedU0hEAXFTrhbuxJMBHKoBePylORfQR5tuLliVPY4Bb0dfOYzNh+I5Ruk+Fybt
YfHFdyZbN06xvGuSFj++eIi1Tq9ZI9u2kq3Je4oMKGlLySxoK/f/WRglvWVajgrv
4mAyaDArjfGgOH2Y1ofawGwojdSwaKoI3qkstebVyBim0SOcJxtq/ks5lri+1PGv
5Qym9Wa8ruD5cZIuqcDZXSKUxKDbBmg9Ld9o9PgQEqKmAF8LT0CbuWQVUJteo0uZ
Vr6Qka3GXdpNrciH3uEP/xLUm8WSFCY5TqwYQDPVL+POmokdJ/yRpc+pfJND3yvF
a0dipz861N3mrDuu5ft4dqMo1CAEf9z5bwjwvo9eMJNIWJ3jSFvZQuwzj1+Oo0iu
hUpSYMZLpKUoDKlj9QwcR9Mik3Na4XFWAKTo+m5rPxdPr1+d+OWW3PNKPPUsQky+
IQvE7bjYJZGCt7dxf03XHrX4IuvwcO2hAaXwbjHNtVoR/TlFZW22UwcElBxf9uIq
ucrYgpPNPDmCKoVPE9oSa5cPtlqp//29EkdNTsWH6AHZSlBS+0eWpK2HvPi8Uz+V
9UOX39TzgAr2EtB1y0BGRgFM9RfRkUfV6AR5TH10WZ/i7hBuwMvwxmD1B4i0qbm7
tHN/zyF+XH0XEI4oF4/4cE53jNNp/7QVedMa7HmacaI9AvhZ4paGwZMizcCEqZ21
PQreXbX5b2+n7yksBQLmOyIUngJPiigTXyJVVbiIBWlbjWngdGpltwHaW+EMbiRa
Fu4wdcnA4GW9XCJUqCmAtf6UdffxyN0MSp5CO0XpIkIGDzaiuHUvvCyHWx0RP9mT
zg7sirbWhOS5+g4sJ7Ss5sweVroqqCZw5Y9ziM/RT/8GsOLchnZHZIOnpwAu5IAm
Fx2WEzKHFVjbo+hw9qCGnjfcZu71Vgzcv+T6Btz7zszF/ba56rE5q+/v3sNi5dma
WPvQF/BqcjumqfPzEz/0xltD8Hr6uz8d2WoUwHZCQYHWWmzNytxZFKkNLoAuRzM7
3PDcq4RDnvxj2gaLBRKbaEd0o9ijwuPK96QvHIK1AyUSn88vs1QJpPRgsZI/MuPS
L+rYOCB+PUtvd3+Wc9abVq1OI089C9/GFiHpwVVthZknskwuEhlh20nvzPKQyW3O
uIVqzDT+Wrr5DlZN2Xz1excdcXsJ4s/AwZTaSiuWEonBfn17xaPARD59DxX7cT1G
BQbAqGxhK/w6LNxDoEJSqFCC9FRPXGVwXFyhWic6tRbElw3DmcYnYjbAzojMXQnk
ASVyN5c67AV1eFzn39ERrB5YacyWapYvuXGeCrdJWecjtthfAniO44KmVQoy8Vdk
MrF9R6UmccGKy1gK7ceBya2Xm/IvXC3szeQ/ydJIiZuxDvdpeWgo1aYavFvzDMjb
CgrkEWxnwIOTiH1sKqhZI8RPU5uXJQEWf/Tk/tx/y4j96Th9oEdgFboIwDA8jFtP
bjhP7wgFuYM2Qkiwt7fz0qS4nO0oE3RwmZAVzPKn5ENNx/eeM89jD9eKi2XAArbM
GvH3B0TJ4tNk5AXvxmYrT61A/Jmekf3Z/4q/qJxAsNiEYJBulCBQHuOOGdg1kbl9
rh0Fnhfskayhj9bDCCeaXkzWcAsRbA/FkZmACurnZMXFSz8cTn14LOG82b9wJ4C8
GRkXgOQ3tLDOs8IiZn/LRpKLfhpOkxn00VJ9He1saiECPFy+GotqYQj4ow3DBGq4
10XhC18lx+e1BBkAc4kLCllIMxrPiAWT3GBj+Jc1kKQSdvabUQ6hHNWYyJFe5dQv
yILl4DRz/4Cb0Fou2n1UYK7tO4OTPCFShBjSTyanjAE9RZPcZ6ZSqYOITHR5XEg4
+efy5atMzV80sfJn/i43KJYJJptKRvsh2ALyEhbZeXh2Kq4McSbQN6FrH+WMCz5E
c0mLkGd2fVa/PaOanT3FUCPo+YPx0ot96V21EgFfwHGN80rl4AmNFOL/rH9c0P6g
63eaTMDfDkTcYUwAVON3J2LVFiIdV6PPmYlf2I97N72ek6d6FagDekLeE9jxD2kg
CrIwXlE6iE+D3jLHcPf9Enl333MY9HxHot0L7M1iq0OtuDhbGtHtJEiIYC/dM5JG
Niy4YNrCwvaGelzfMOkCbaT3Anh1fxaVNlO+5EH9IKZzn1+U1IGIFUAyiO652IW1
MDmB6HzEMfUTDspZiTIYo+ndt2QIExZeSwN/eb/5m+js5xmuqIgW4LAovkuEhF7t
L/kcNEXyUuebBx9ugja/2gNysiDhzMgcLAsJYeVDbBuIueilVUGt1SvKWbU/q10Z
TfUG0E7PCEkAfO5RhIidFV5TxTKm3XhRtU+i3nIe21II8yjN4Qafz24WLDpk2ppR
1FkASX5ODkDr6Ifz+TfL0aQPGS6wf/7nDT95EPWNAzpzpBrI73YVPujv/OJZWcsr
29DDt56I/ZHoslH3CiwEehl1lhk3flFDxYeODr9Y9DUPU855nxFVcRIAEjJ4Wgoa
7fvAS0ldmhpXSgFhl84io95iSx7EJ2UEQcntejT7SHacEYrwTrZ8kdkSLTqZsHY6
330q53gWLZXSQKo+Iyyj25Gzxch+jltVsp9vpyZwDLKRvlCgPJLvjb/eshnkr+G3
jPmeTl7pTWzW/9CZrIRMkrursJUAKgooieoOG+wPzUrtnCQGlMFtkUVjOAsdv/GG
OI4RtwAPjA/yiZOI8pBbzjaLAzPoHL0vxzaTR32lyOvrsGXDPnoP8dgqEQmMRBt4
t3ktXHrSuDyLBpvuCILqnUojRIn+1DtvT0PUxEqhzmuaZ95vF7+d/A4Zcl/BO/F+
mGc98dfjo5/X6MLqJ7vQqqoLJDMYqu2Fjbo/ofgl/6mgAOuMxlXD18BRo/GDWOb5
PVXwnKA08pD32UKKAWrT6hZ9oubw3pURoiHzI9kp7D+EwsvHfUqcLwUYWOeiEKkw
WyGx6K7Zfdtx0HIDbCY65UNRIjRk3RSklgFxl09i7v811HlFIJfOfyhNAOxUvDRa
phdn2IkIQzsbODmSwkrM9i89jeTRlWP6wR2IvxX8nDh+39PI+dAGrrGUV0b3d2wV
9UHLtowUHIjh9gDUJIOqt65pZd6QwJo8/TDC7wFufELbyoGDHb8sv6nieU6BUnPY
IObQ+EOpV55W/4iEk/sBPV5knlWemz9ADX8kEvppIQ6mnBNgOWvrTOl/UzOWicDT
Dn9ZoasJLKR9jQJWNna9SUnXa023cxX9+BTg9Y6fkO9JkGUX2rPJBa09ZzA6EvkM
d8o7HHDFQLu7OEpkyqn85mTJ5mxtDaL4ci+bOm4xW0ycCRA4FsxqTXW4p5ujSMs3
IwsFiazDyqTkGxuX8wYkZL6El3/7iWvW6KlXKnqqke7XLcFJuZRziRZslOD2TKV5
i1iF3tgSJ4QKbRBdm3KIgsV2rw+rW9baKfxG1+sHWuGk38eoiynZeGF1mlvIiKg+
egMA+wizn0NmnS6/LFHiuSUrU5vvP9ltg6yDG+pB1rlFOp5+yJAEAyIPsXLLiusc
pCprSi6yqRCZMgkg0+In3Vz3KiiS0q0OIYmFvBR5hkx2vHZeUImQVqoZp1V6GlPF
1azKaI6CFr36ukMsRngT/5FAyQairlqfK98ZAGmYQ5P5oTU83HBQLgMA5rdNoWHp
Coyh+1J+BoO6leFS2xsjYZSn3fPg5aDlW1faSM2fr/q67iNsKT8q9XtrCBy2x+Fn
xEyDFYEg0Uv2h8KQD2fdFtJ6zc0QmZfYzXm4UYX9FP/bW+TaXYKFkOEo8TpWo/Xh
50FkE1pHfaPiMLPQ9usbXbPCvLL9RXWTCqU7gaW3BLZwpthYV+a18ubZz1HaK+70
jBWSSCuxEqa0wtzpaeIf801gx4yxYSwe6vWYr41k7O0iQ6We65H9KWZZSwg5YpF5
eL0eiVgb3MrT65yQ4r6JON34iIoZpiKCWhG8A8rEm0wFlFy+4uykgedFTYzEmEUT
idHWfUNU/x1GO1oftRRfCrNHLdB5u7vR/yhghFO5fP/f5sPiDDvxRjIfmBKbsr2M
e1Rc44kKV0XKhlbH0mdJjvCewqHwA9yUvnh6FvZcQP2EfyN7HDWXtSq74RDBawlA
FnAJhFzmlzQ20q1fNGbJo/VrCjDa9ZFF574tPFjZbQfJdiMZYcmqbRQFN2KnJD0v
bGtGcA8tsCYba+r3RTtYF7LDD8OKmIBfm+myYqroZ97ooUSFlnFhjZyB+y5z0ez8
xbsH+v+NnM1oDMbD4AgN1NvCOBFnPrOTTEwJfsVb21TMtutDhmIYaZRwGaLXw/Ex
V9myxfb4loEAz4tD+SxifSLmkQlA3DUGpgeuePN8ipv142k1BCFQEHPnvc+1D6MZ
AC5tMOTXpJJd4S64NRsccGBx/8JGseRnqNSFMBe8CgouTccHNfJvt64v8WZDWkrS
FgtlwakxA9DPZKWbLsaYKIx0IKMbCIqG2mfue2KLjDTNfaRv+jpwxzj3olW1tvQ7
ioq6P9avRnNdjBVURZdDvPLs/YoCbgYPNf4naq5MlySi+ucbXRq7O306pevFl9vQ
/8bSObJT7SjnkUFz46aSEDeZORoClx4wH0f1rQvlQ13ZdUVL9EVhA6pdGc++RpPE
WgM2m5l3fuz6La25jTLDaiOmVFx31XS4sSxfK1eZS2y8Le9Y7gRY+FpIH+OlB0s9
r6tdlEVSZl9VBhG3y6u2sBt228fINLc4iaVBfvZePtnjMJgPXadjMyxIoN6KdHdi
ijtpTbW5gnLBQHwdGVv1g2UKeovyIva0dRJiSM5P4yQsXrjaqSg1IHcB9qE8AGb+
JmDBaQ9K2/HF4CWuFvJtfeanlJv1ywAWpUj8ehXuGwJU2/4bpt1pwgGyMjLwZkZK
yDCblfpWLm16jx/BfIVZC45bIuPlhALqysCeshf0gicU5lpja28d7ZZ5EQSVOleB
MZFG3dEEfK5Wq6x4srF/lCJcS/D6+ApkMpgbUctiUclTvkdNHcMgGc0h7a2cctnT
hPgnGTNAJwtMmCxyEFnFfFZ+FW2UEV7c6FM7niWpUiqsBfgXkqs3yO08FvnVFY40
+LMq81xzB5R+qsAF1X5uF9KhScGdkDtZere0b13pma50WqbiaI+nJHAMd/OV1WUu
KT4gZqWi/5awM4lxywuL1XnH4myxHTpgv0IP+GfEuYcVoEykGpcSjpGg1iHgNJfu
19WLz35QBjM500WpPjhrm4UYIEd1rpMKkjISRBAZe9LhV57hbeT7bbCuJB/vDMBF
hgdYwhT25StZsbY+WH6VidgXRxtmxXRgZm+D/b9jWJp38DVN6GRNh9FSRpYkwqm4
zMDcEH1lkPDZIfH8YxosbVLxI1WnwTO+uGrxJHE4C1bIzKTOh7XO/oY5Y/7Pzebv
zkb/0fBDgTjYRQLU2eLEVbeWgQwmxVgQpCAogoVfRBHCn8lyltePqaeIYMwO3bpQ
Uw8TT7ppIc+qAE2XsKUZYGG+jsQPc7cb1+qV1mFZh5pH6Kov7FqTGZDP/qpN8HFI
98U7A3A3H/TIFGQzpWJY3zUlsdu2g6M6wJPHCiAqTrx+/f6f3QjDm2zTKVGV8ssW
s5LAfnSbSSjtGqSc4mYTYnP6OXpH6OWrUl9bMcrF67m7OEsC1ONoSPIeTDwertGn
+8GLI4nS8nhVNMdkZD5zB6cW/8dcGU1NysQM1qPQ7EB3uzOe9XUdURXonKn2FJnt
tm/t1FbS7WfJRwCeHwaEd5N18IE3JIku9MkjqADyim5FB9n2NzO5kFdjBUJlTCkK
l28quAPGuYHynlYqW4ylyG1dVXjVDi2m3IeDuDRhoxbjxB6I7HlvmFanfygKsJxh
7LZpTMOnh23bZrCr8oIZlvDD4Ia4gSdyR4QqnKTNJmzewKtZylpVXbt+/bt7UMCd
bMD5GUH5usHeO8Fg276AKEWf6Rh5JhpWhuGyYfEoxmedG6SsFTYgl1XZAEVGvb96
zTWJY7bbFgE789kb/ka5IsLbd0qXYIiIyi5YYEn9LnVLz/e3HP5h3vlx8oBxvkYC
dDmtBr7mYzZ59sj6WAoC62oJD7LCTt0tlKdakBGTWbtgMa8bmfRVN05wt/a6yepJ
jFr9NlEoKbQY/fjCJYNfRQdQdaFvPYr5EcSL+IgJAtpv63+ccy0wZc6Abtx2syBG
6tGRJ0dC1XCvXp8vV8G1mrIy2Hg+LVNCj2mJwiMFlz+DGdYb76JZ5cCflaHd2zsE
jlQiQFq6bIv2p1nYnRb0DgYgH5VJ0PKcoDPPQjyn5thaZ3zmL5WwcnEailvYUuJh
2y7BI1qewklOpJtfA93TiB/f+/cHQx8ObbDQIlDSWxYL+yZAzFoHG8q7WFBIA/2R
7g9TxL1QCLDDhqfJmMhGLDqGfeT+uDs9hRvsk4gctLYsu/bK8xPiyZ4A78sJINMf
OSLeFF9+CxbSvfJWhFK3LaS0SP8t8sBGrzW8Ea6Ikt1R9DMe4mobwj7586+rh4RM
oZgtxBdG9wJqUohQKc63DCsbnwK51eoB78Rl2qWz5RImwN2xWvo5/1HLan0dHFLp
n18KU1WiwIRqObkt4lGQOkX43mZPqYiM4eq/uNadlZ3ICTOkyYXr+4rcgV4/sOyg
8TrPrGTz3bzetKRUaLeQweXSiujpsIfZvZHC53zD0OZyZIqPHNsAzLofs1HSy9t5
hmd16xYsEJtj/1KxGCrBXuLs3gqpgZW41q+ZvNRl0ZrWZaC7JYCDjUr5vVQYuS9M
MtW9nvleaEKi4Vt4WsJq4omfRtBTipUDEmWxF0mPB6JovdJUopNKZUgdcuxr+od+
MikBN9Svv9z/yZZN5I1CHcyG5PMenU0IDoKA4jZymvYUONO2FUmYkd+2YXZm9NSy
e2yfyp5Ub3vr0CgxJ8qhWTIQSi2tGrt7KDdsi41YGp2fmFFGtzyGormJ2Wr0ri88
0xDlNn43TfZ63Sow8Xle3b6g6iBc1ek0P/uG5cPxmGUo4rRTpbk9uUNyB7eckb1J
ZMBw7pI8wGzvWeOcWPJFtSIgMIgxcx0ELGPJEi4ZUWAqETsyMI3FtOUV89tPvIJN
zlSGzbyXvZt84IEPWbz8y33EFWlqufIb1v4DwO87uwOeN8Nlvzg1VjKIHY+iRWnO
SPUpAr1P0vFVegq9Wf3DJi33Nh1jU5DdbjmR2rsiUsFkREvZM6+Y59s73XnTTA7z
g1TNOGf4fAJNS1hNYRuwsfowz7hImpxPu1d+dIeJ0Yyt9ZdZXUI2VHvIDLXjALAY
LHjARhTk46jq37k0kzrI9lrBOACA4/EWLWp8DO9JQcG0omBKTBFrOponHnEXhrBL
hT8wwlCY3Gs+mgnQt4C1N5ymKQnVCHjhoXF+FBFOxNJPw0CneAQqJiV280rhmKKx
i9d5X19GCDPKaU2bVlcTLcGazb37opLC5JcM5oGt2X7vZyzwZ5h0PpAEzYU/zCg7
iZDvU1foAblNQsO7eiOC2ZSDYaVCOLq1VmdyzVm0hZJMNS1Jcw+xc4AOaPY63C+X
EkHqZ7CR0ehMwDdWpkIDXmejalMyBrPA6TcZ6bea6b1v7uQ7sFtuoUsX7mL/1gAg
eeXvoAHQin5bCi3isTQ1bDUtjbUuVYJAV9GEutYkwQx3iHVN6no+3UhgwmOYkzW0
6b3iZ7PEVXbGjnxZS//uEI/QThLbJfORw8FN0liS0CacwmGHR1//bIDjfUWQS45o
lPckAbduKMUsAmEw5LI6IoIlpCQfkQuPgIMR0liAFb6yKdVuCRK3uGqj3IRI5bOJ
FMQBCNlKbpGG23nmLxfxqwk9UXcnHK4R91zeKXCFD+IvDYBRtAl04yEe9ClMfhWV
PcpwRgfHsJFndESoyelZJm6EJMhpPMDo9pSjO+EDXZpaHPR4gYPdJbqTHEE+U/Ks
4T4+2PwYkhJDvfF3uayP3wLdiFbxjvGeZhGdeB7EvZfPLJm/g+FBjsSFjq8KlFO2
R3id2+Q6PtP0WO6S5xCHXB97mG9nZhuzgLmt67lapC7Caq2o5t46i5pARsqqDsr7
tuNnxW+cferV+JHcsqGL3+fMUurMUcbLIcQq/gj4JUD6u3p9/021UKRycx/3qFfe
pvm5gAh2GCfNpLewzPAmF/gOK/VtwRtCMHUaDzsZkRX6+cR+t/BdljsVwVyy1P6q
WiWGdLQBXq28Ji/0PWgRK5s2nfxbuYgV0y9yFKvds3dCfqqcAqw0OMVxh0ffC3hG
o6E0sFOP73hVPwsBuYdQ/4aEPg9xCZWczQaw9VV12Ex6G24HZFmWZW/yz9FYn+hY
joYuZAW5j4kCgJTTvs3VO0TsyoD7V9j0/EmQDxs62scSA58RziTa7CseO9dkAB2I
q/m3H90p348XusYCXSxigGWCAJAMcIIKoMdcuXDji0mTp92HilayXqizV82i5ILM
WN2shFPrOANfx+Zgao7HjtyA7uRE2vGNojxnCKrQPOCG4pQb/FfC8Vn+iZ5ulqjc
I7u8/cd2+OUaKRU4tm3EIl8kTy4ibFIicTB33Q2Hq4RdVC+DwajgETveyixyCF9m
6dFcn8WK7nuWDVSItflvD3nB7VIfuU5hfqDlJG5pbfLe7oQIEiqywiKqqLqumVdq
NPiYQzNu9IH4o7FJvvUqC02aGjBQOscqvUMKlKdnaX0/seFT2sUf8BIbsZ83glhP
0zJMz0oM8z0zHmhCURx99mkdnYuRDj79s62zpoWxVsfTAFC2a92sAsM6VmtaakyP
/lP2dap/rsBfhMQikNK2ghOtnu18C7wBReRTUVvYpFE5lwRwBGvW4Ho+Zqbzxk/h
R2vn5S2cuDe1ZQpjwrHHVlDl9C/TfjAcPv9dr+16jnV3KL4Z3r6aZbsFLj3lHy3W
ctsVzcypNZwxbQoiImLCnL2REHnjBp8it5U/3s8VGUxHHhVc+FN8FcO22VUYqACB
1+PSIwbP8Qet5bJ715X7VvzV1eTNE1z2qOHpPIsUqGop2EbcTtO8Q9GllbfeRU4h
0dJWKN4Fv2CWvKMZ2fMIBzRXfKTt8szmG3z1x23ARToe80t7UlzarMCu1PKVqMfF
zKwDepX110FFfnacE0pFDK4PaF8ALCPIdMO32OAlWIS8BO3tngiDXs20v+9PzNld
U3fDvXJQughpdQE+TMjky0liLTFX2MHZ+vjcMwDuymYdzJBDuLu7YSCqMX89E2Oa
UZ/tT4/Q6yCvWJZEddIHorVHrPVGb1oFf8lt2I4ZM9LO5SqS1jIPrWQRcfrza8Ih
cQY8ZfAkcvKuJvbFGDpphfYXLgQ87ln4UvICNotpGENHbqhx8NqAoe4p45jH9CLM
OuITzeFWVcruvtdatHmwyqeHaiRp58gGMnU0QJP3Jmz4UUBP5b1IKVATBRVMfP+j
SOGX87veKLhBY60bPAeNNy335XA+qLMOT+FOYtWxKrUl86szaQKbTZsCSrQpok6y
33oFVsBlyBzwipAVd42lZi6RvnGNogM65a6QKHIho2Y9kCaDavvBk3Nf+BEuRKlE
vLj2JLSkD/THfG/csBA2/9z7+7lb1jlpCmUpH1Csftbbvp8y3jsiKGILbK7jbozV
79lAjRKK/tGafG2Kc6DxEWz1+rsmEHJF9d8g369sO6g1nRx26YFr+h5Oeectn/ed
fy53j0h97BUkLCPL9741y4mVJmQeYG7JA9MKfsT/xdIL9W5UmEOCeGTAXpnzdXyJ
IcaefNFxIr/QmbR8QGV0FkCVx6GYWWj49ttx74fmXfzE6bJcBD3gFUDYJCIp98zn
delYHljU5TwdiEy52J70VQKXe1PFemsYEcjkySXnZqaXIbrsxapyoMNp9b5NICW1
QbP11vhcu82bh+jKCtm5YbckCotG/6wAotnTU6Ytv/QbT8kWSYlYMUTXAZbYNWR+
Oa++bw3qVG5bzteptBP/3/J67W4j9mSSNsZMATwTQDkD3ipOTGrWd2o8J4ZYi5I7
epv6XBf0PJUwfdPmklQKnucypqP3rRAuuch9qBFI0tBQyzZSaLsVp5l1qjYrqJUo
0ErvnEbxd+NmWb37/NYIeocHmv3mUerTDeSCO3kSGx2NxQ0sPpKA8vTXsVPoALy0
V1ksiFNlJM/NAZFl+OqWwW1EbM/yBtpLVm7orxQvMYSBrWtdSltdtZNUMN6Z5vvB
Ue+XQZ1PhCWmnqOI93PsV/jVP7fVN1RgZr28kBxqEjSRriAewB+Am26P6Jmkuw0a
Dq+7XfT2JR8WcjHnOnOQ9K8KehduzwVBOZvnw8LlzZFh3HAC1k5oo6OnmNagHI0Z
H94gPgfW/sOgR9UY9M342GZvl+CpXXGLQaNBD+8YxZW66aS7LxVr/tg6Ips/E4kd
gHg0POHimqLS5s3j3B4JGGU8s9xIq05kcjAaQum9Objv2+Erxc/rl5WbRHF81EAr
q7LBf1RzIGKjjJVq0h7+6I+fxHrUrM6GbiZReaieDITnudNrcQIZi+6u00vOJofQ
sNBe2Idg+SwM9/aMJ7TBStXqZ0XfnnDkK49DYqirvibIQWtuUCT7ynweBuY+usaO
d/zk19qT9vdMWbZi56ec4qIvPIKxy2e/fKZbrn60Sp6Ogr259J7QhMNrnJqzKoED
yyC7gAC8C8lpf3YCWfy0VQDBtqW0K5ACjAkVbmm17kE3uR4tzV15aQPgWQbPnROE
jRZ+mWHYFSOwtd20cOiQ54tTknc2W9HSSL+ZBLKofn1Nquc0hJxCusDaToKXPczW
Yp6eCEnyHykM+tM9xgWwFZuqsYL/RFnu6GFwK/I0CPPaz/SqbuqSddyLuUYfDKyp
Qxi3P0eOsbs80qmQ425MawXqDDLTig88YQIfwhk3QY8NP/wSSMSlTGfRRVSRFzYE
u4C39F7Lw1s9CSs1VlQmMHqwA6noKg+Bwi7C8uitllMQHL2CFUO/HT3yjq9ZnSNB
i11WE1856CFs55qYT2cxWm7S7du6dVFV/XWOjAkw7e5mi2pwEJkHHJ/zr1X46dIW
05Rou55O7g65KMTuhTsv+H955bLKU64U3Roivg6kDqMoz5R7VVi+iNFGt7Sw78yL
b7fu3BQD2KfHgFDhFVw1ycuG5VlpTaqvKTuOKQffwVs7vpZbXr1BE1GT4nKJ/i69
yQSMofqOrq7EJjGoVAF3Bl629EOCuaRIjwXw6N+uGIZTzcKbXC8caPvJDXcSsd9o
z8whsT8crqjEedD3xje/TMfMCZ3cuog25msuf+ISXAXusP/NZtQ82H/d0eNUzUKL
VAkr1IjhIxVp+qEFY+j7ZxpvBAfTt4ngvXDWz+h0N+PsIdoVOCQm9tB5VrWVJkfX
HHxH3fcbfpQySi2wZYGwTFFPLeNTHSG6qZhwFrf2XaB38XkxX0s72hGF+GWKiuhX
t3WweY9W1JmuqIX3hmPL4txK8sv9DOPq+sM4jI0UTHpNean9CW/gIJk4rU1hGyey
oux8b6Nza/C7dVqhWUWY/IOhVBUcA/aiLPcvtxIMKnydg3bD2xXMHDm899CTeHdw
XKVaizWRhdewMduTppSN9IY3TqqbljV5aWN+SonYJXnGZ1PRL5A9vboWJVjdfDLu
t9xjlp0lMuw3CbnCog/ridkTDSzR/Xzt370LyflznjK2E+/uDUB4DDCkY1hRpwtk
zstqRsFak1jG3RTHeEn0FCpvzKJEsxx2x+ih/Dz8c1oeZIBYDOvxGDkPzR4PNEBQ
4W/9nEZRr8DwMm7KGEgnJziHhXeUomfYf60WOZlHLOiXntidlzMkDDHOemXykMuV
Kae28/yplqZj6lZOqASApb0mdl9mtgwKZg/rfe0XxrDf0tnMPV9KQ/AjCiU7vAHP
pdNiGMXeLZmve2In0nTpUDOUdnF90RBU9Wa4DGLm7b/uiJY7qq9AoyL4j/P78w5u
DouZEgsIyccFRai00VrGwLw8/iB8JKL7VSu1Aahw74Ukb6km1wpQjNRcI3XGRxB0
cZ1606GSG6cCmj1Z11c9L59K0xO0GwC+53V4awLLPNYNfUrUQbUdiTxylNnaO6W7
1BdDoVhQ7jCASZ1pw6315mPRpAgZK8BSRo3wxCXpTTNixWYYCrw7Av4v1FOuup1q
rUF6gCn38+ZRM8YLl2oAF9zYQps26muAuQOEulUehxumobS0xZebon1O1khMNtTC
DirwBkdNAAYVg9ovGITCCb0Yr6aMXL7UMfB+haPfl8LZeWpjbmQ5Dm4UPWxQSb+p
Nsfc5gRw5KtRhG2jKpqf0TiELS5qpVTjXBd8HQmpFy7nr3+HmYcsa4pIDCQKyPQb
rsfA1W/tb8KX7LiGgB8Q19ker1b9jpVMjaLJCguE8ar70jdvCD8wNk9/RaC22g27
A9MLxmIi8YIzCy1c5rv4NC10SCJBYX2qBDVWMd3C+Jl87IlTB4JS86vqP1knflxj
SLKLx4XTx1nijQGT3W99cvZN4568atPrmh7Gl7KkyANcw1zgQxymYxrP9BwsC0xR
e9DaOI37nu/PAIPShVjx//kW++jSPnmjykLwXRF/99iKddsn/eJd4qTZeqNulqyp
aBQQdcErrW/DeQ3WJNkVLEjVuNY4rfVG8znnQiui8BcMeSyEEZ2X7fIiww9qBTtV
2JJ4mWrRqCxHb/ELq1oYqTn3HpP8sMSO39LSA+bBOsdD9X+2koFn08dFb9/X+k2j
CCs9rAMImKfK4etM3TF8yuA8qlXeeancUWDcqPmpbZEpPR5Ej0EWDgOveFc7XHpn
zJZ6H9EsRbqdlFTspugeOPVg26ammHE3DYugrwglK0xU/go78vnKPG2qvBQn3aDB
wALG8U2KjCvrldq/3ekzUgQFDZymGC8sPSTji+y/51I9iq/mReC8reZEXtFG0sGm
axiIVfZzb+OHG0ncs55xUIGNO6lgDOqMeWeVYMOtn+Pa7fHRhyC/cZCsfRwlZbvl
6O9SaK+ljViZC/Of/QeHiKYP20zw6pUDgAt1Uyw4STKvb3Vf6T9NcOauP9AQY0Yh
avPt2XUwtsb0YQTI7Nc4TnkQ9qWuB0eXEjp6T/Ib9ROxO7S6zmF4kPNekznE7Wps
j0jQG5QwPwqR/TYK/XYYK+x66KuJr1vsP5PxBMK2YIu1bFVZ6p0mnS8ylcagOzOB
5MyQKyn9x7upU5j3g16HR4w1f93kqailuvXCf5ku9feMnO8fjcE4C+7MJeCjcze9
6SgJkcG8OFKUn8eXHphU8avHA22QZHB0Rnblm/WA0Rovz5GqiO+yN7wZdBhPwJ41
/0Sx2fTaAJsVCJ1QinISL/9U6GN5kieOxuSou0rSAH/oBZbAMPUFg/X8CGSqp067
jxbcAi5szlZ6NLs+FxjHL5TZHfcYIyUNhvJhp/Emh8aAVIfnFVOxIdPDB1voqY3O
iumtuC3DB1oZv++lyudjChgJ1E0xmN4u+tqu4h2QcOKREAU8afv7W+NmAgcxcUcq
cK+AmynS62wz85PzWQQu5Qu+s8p56kOfzeLUO/SaXGUA5bZVCh/ZJnPbM57avdNu
0IkK4Gh/w9tTDsBQnff9MLAp6+vmtojNoXhRrgx+rbnMPi7skYHBXdZ2nzA/94Ms
9Tx1g9UjCK6+f0OEdKyrsp194wFMfMZA8xb7EF5D6n9+x1EXuqsLclMAjGeTL2Dj
AzLiHcwCZcp/eestsikys/MmDqeI6Gy9CeVsi3UYqNZXjqF3WGzTWG0oOhbTqsqD
bOA6I+E0wQo3Lr6nM3gDvfm2t3Lb8Ud8t3mC+eW6nfpMdw937qs1Qq+vUTPkbP42
9en3IuNsbA6+eL6zHBQWceK39tt5ssyBdsSeTpqcd0S4hZ97e0EWgfV8dpcp0Lh0
u7S8RWJHN4+xCEGsH85DrKDarENor97/CTzMvtuxDPj/pl+6XWKEyGuIAov3Ihzj
T0mWovhq+wOZ85VeLJ5NUJ+VFlCIgmgTE2ebCeVvbqvpDyZXTiOflrGAdgHUOZDL
ckB0kBS9vYmnrztEuA43nCf/+tSpwYliCTc3nlJlxmGLLeL3BG+9/spU/Q81ibZr
Xy1a7Eyi+JnPLjDJyt8Zug3IJCTdxVnkyFJRUaW1rvULEPSJGeS+iLRzRqxfOaGH
m97GCmbUQAfdpUWhRHt1x2rnhsAWB9fLLn+x5BIAaWFaf+6wyBafgaZt0TeRqKdE
cmbY7Hau9B4sXlppWnGyP+NOefd63lAtVOdrJL7oFwuifI9BfeesO9O1AMYurV7z
LAOrW12ezmHqoIWznp6ACW5kevHmWHBYT/JwHcyuEy1/2Oi6bnmxQwCiF7h+NVRi
NlH5vRe5hBa4YIPvJmQwExbIsXa0TxAVPnve1MMlqSo77T2Tvc6GJmJhBwNt8d6s
apfJzjdVo1/PY2WIY54uMTiJ3ixGPLGTdP54QCxhnTlZ4gaMynEMTGpxusyNRi3R
1sUHk1e1IUWcyW3SIwQ1xB5EQcttld+OFsn5NAmwL9Yiq9bCSghaJ17Bbl9/vijY
KeCNT8UoxSLkkzwsLlaTCy2Fze/22nKAD76INkwzPb47jAI+eMVgZVKLpgEiFbf7
IKyfgLxVRVyG8IRGGgpfQ8SpjVHt7MCRMjEh6QQFObR/B7y0E8gNfubAuhlaFOCB
v76W/lG1D1nCwTq2DbW0aLOV+QBiGSLh7lJ3EQcouzSoE66NQMBuU39d4eKYLsRq
YWdMGBg6etqlrDePMRiebrnlhD+aSsM28trMdd/TxiDkNfjoh3Ski0s55W83lL8Y
BBwD9jfDMu4STO5hxpKFX53uEgdy+4tnRTMuBkb3190ao4ncfO4nlGkqDomgRP3b
TYp834XN625DhisMq2l1jwj5J77ojfklx9cFPyaBrvAnYzi67Vr1k0DHNmVBEIjB
Zc9kBNsqunRLKVy/aQhYnHGmIf+gb8SOIB2n5f76+o36Whr8tbDdyif09fFf8ZnR
D9tDLi65zM8Wqxo4EI/hwPUVNqGgxzrPd6cHpir3nuUnSab7uf5IpBdDh5c141pm
/epzksUOhoGeX8IUgcVYa/1x4jmHeB99mqRBQHQd65VCwBytjDHUS2yU6WJyTQ8V
YXJxCafQIAS8oxMXb8rs/zaXpvSE32fIp/4mVSsf6WKerT/QKEwMeKe1kDeZ+h37
qJbyGBsGi6Qjx/00xF268j90POZ/t7Em9zdKSg3CWw+E1Fh8G0NkRI+z2wq45SqO
nOw5IEAWatbCkSwv4qtIpmU5sLa36yGYIsPoYn1+2HEEODh4irPaukSfEvTsXzCg
Ah935VfA4GS40mMqu424404YqDGVkvoxVWLLBhvDf3lTMrc0bYEwE6cOWGRmDocS
yUb2FFegO+hU+7P6AXs97EZRnV5mgZ5Ag8p/HbhQQuKQ5KZqK4X2B+owsUsGpaxo
XrRl80VNa2eeWBcFFSrfGpe/KvxQI1aP4BHTR+prh7yEo4PjXNnjtY8yCl4cijsm
Ea7TDZArsiNPtgEwZ8odf5/PZZwOioRREJM+/e26AN3J5SrxX0jEbqFQYnBjQbHN
CJk4kl1r+iQscE4LBLiErMmBw2myPwFdfihrcFmTKtuTsb4G0WImzOAe1QWtud4T
gWFETedhkT19spz/DORl536jISVibgjCjsVatzp4DhXOs7kqnmpM3yIMcNaP+4T7
vgypRfKV5L2/tcsFO0R+RMXCCRCjxv3dS6zaNccZNafzWyeAaKO4kcjSfO4p6ZjA
Q+nBnfxnNggwtufCq0vyJXdc+ZiW9VtzA5krb4ZicbQqDN0pURaY3EpTUGPnRT8t
vR6xi6ilhp+Y1vRD7mxMdmVjXaX07cedSoIfacaKLycP3PgGkw6+PwBr2sK0dzaW
KHRn7DdB0PoHw7FFuICMpeo8mOkkc4JTrS0i2ubya+lF19rDgVs/e1eP+eypMje1
o+Yr+QWIyGomx1vvpqLIPs0j2hylq5S9yADn7QCcdL5fDrevErvocEcvc7J3h991
VOBJUkxinoO1kz5/wdHibzN/6loyMTliwOEWJOP4fq5iMRv68gKJjkbCRvhOuukA
XkHHoDXFkZG5VckPtqFshnqM3yZX7Qxyefg/OTxyAa6+0y/qYotZTt7gVUZfPWSH
4MxdwJmyBgURnjlQCkVme0FLVRdHsdulM5Ni0Bgon3tVfuf94I7+bTH5o6a50qc6
QGTkLTmlEKT1WZmWSCy4qvhOaQf3wNieQjC9L6zWbSOF9se5r4Rx6g0sauINHeLL
wgTkXpirw8GI724jnU23CBR/YZq3DzLapIf0eijyotniLVtXHEDnx74eCXNZuP7U
KhAEJZG6Dg+u3+wPqoyDcIu4EvvNqoRXI9WMMWzjHAoSm4aEFo54YL0ltEcGh8/1
VjSPy8BuHnREM14jKl//Ya0T6SeBSAQqrocs9F8Ksv8jrXn+eyhZ1Q1OT8YFOKdb
5hhCE3vKbw21MRDx5xnMJokAC6w83v9Q5KEz2+yFtVxlTqfYCzeQvwgReAEXHSuT
20hpqBOBF5pM9+yCtzq2+8LLyQ1JYSMuNVn+gRcZrReRX5JsMVAjuUz0q3eGI4Q+
CFM+gnwvgW55todBURkjJFElpsyZxNSoAMxfbAM2gMSP6Fffig09FtnuFih00FOj
poLYKi+yp3QQfs6h9gGMrSMsNQ2LW2dTF02POcLbRC3T+iZOk+FPTHr8gddmRZaJ
ooNilb480DRlx0Oy/dC51ii9gopsEDfGJeXf4hnbRWAEYhW+CpJUUeTBsZML2Cqj
BP/rXZtI+OGxvCf5jG0nhSQd0km2H5YTxcoEWK5KFqrWVG647OzgNO6BeBFWUHtZ
J04uve/KJyy2VgpHOTWEdDGnQI91Qy6nBb3JntFnLcyT8uvr8/qH/4o/juZ3xn3J
95pE/Gks3poN7BTCKYcuZRL/Mp8J+yjoTXVQ3lb/XB5Se4REHuuCNhDCQowOiF1c
um9cyJMzN2Qg/6o63bpTPse3lxg/axGQhMdcb7MHCv5NdNJeruI5eHo6mo3SQKfe
emJNUw5jCm87ekNffzTadVD+uhNEMDsKW/Ri7gdwxKHX0cXV4qXFJD19Wa/H65TO
I4+kkSg9TUkuPjWgvL3ns/kYc7Wtbw6poHYiy3W5+svsjAYbZarzf8/ltLOEKqkQ
GJ4HSV2YcNPVKdGn69MUPC6McJeYROxepJcMnPCSpVOYCT3R0NYS1dGEE6GN4JKe
pb1+Mfpdg2YBAYE+ScCQWbRiAv1qJQcnLWXWx7iHLOjmUsiJ8KYaYzv4TZJfLK76
p7QlIRbRMLnnFhWVBhIPnpmiLfgKRi1WqjIYKZnHrmqodjYDYLkbrGM1TUyQ+2FT
Dtwc97fg9toHTOlncZWJJwPIxRBpWzABB+r0G6Tbc90I29uipkHoy7L5DWR+NO49
i2Gi4nJDmuwm9+g8c8NwGEwIHZuFWvA/sIjOcmFTT28Ux2A4ex6qJbGugZu9VzBr
bWfLEAd+XWd43ZmMt9R2gaJlL4NgOhyC93b8AcYWXT31dsPXaiPNBNCW2C50Sm4y
qM5jd0FFztUdVqPtxrVncphd8FHWE09AQUYDkLsVYv56SmD22G4ZvAzld+O2QQzs
gfuwy+Vy5FDqBiJH+4o2JNxl1yc9IAGfuKTJLbMn3PwMOtXsL7LXtv1VV+Nut7Fp
gPv6q51jzfJy3CREMixnhx5XesGVrCYx5y+Y8SNS0efSgr7w80YzNhVmk8jNKxgd
ZF4VEWyqzp94anB7tTbM8u0ZGVrsW+HORLwvp11NEEw9aPqYDiychZfx1RvXsBr8
9N9aDEdJ6ab415cyGSg2d21BdxnTSqjUNqopzc5k1I5BuThN1ga3e+JnyDZGzNM+
7ECt2FyO7hfmjF++9uLvP4vAnvVE0j3Myx7Er02uEwP9pviM5rOL9HWPOGJPUBgX
gJMYnWKZiYyvBy5QCWMxh399XaNQMM62UTeH12Z6C+mAVY9Sg0CkkTkGLtemwYiK
yrHHkg1ZA3BSloxQ7Dp5kzMZJBhRR/LxUFGLrh49dtNWpeq+nTx8Y52JaeLU1M+t
0kFE/Aj5Gc9HEXCVvWV5ZTyIU3lgr671WDP2Tuo2WqZsNVPj4dUGXalprmjOTO0F
fleLK0wKoVHBuAtqR5nGKRAjR2xYohyl1sfOrmokKaXaHhu1xGEV+ZbTzojXOBm+
4lStABe4L+oVZ74792DHm22NWkbgpM0/vOLZPVUAPyU9zPFUdIZEcbBmRxSSQKzv
rYZvR3nGZyH7p4YUNsACTKlK5OuYsMeDFSQqsNPUxfq1QMHFlbR7vEs1zpFldHlW
6KmT63l3iv0ElcjBCbY5S7TLS4iUmQv1+MgreiVQmaQpzVrmurTzloW3qPjyfOlg
x8lwWnRmH2vM8qCl8Yr+Aq5Al9cXEpxMltaDAE4MEUuGx7PrzI3c7i+wuePBMWKl
q+8nwhZqUdKiviVPZ80WhBMbOpPmu9OBSHCiB21WBeKvBFm3cZNM3+1AiaYE1SB6
3emGd6lM4e2seIsFVC+lxyOhmmDHqHmPwds22HtGc/pPzycC5BzRYeDkDUsO46JC
NL8G+CNAWsWzSDTpzaFnSCIS+oQ6+3/NwXSNfvCxcGaFTvYTZy6UQGZVTIZjnKnm
jS7vqAqFqU9rRfjwiaS4cNcOZBxlyQD9cF17pamaSE0XdKs0pSPHuD5BdHv5pkQj
II54lY4Yi40+VZ/epgOnQPaRgbESYE9oaH2SICxo+qT4DHXKtGZmwPqI5dGqxfYh
51bsM09cRYSTYJ/kcXsc0Ob5tEiwySlpab59Oy0FgZKEKAxiGHhqjy/3RfQ3zTqR
nga5Je2kePYEu6KBieWapdbW38t6zSe85UNiSaggzUD2N7rdOZ/b/CvptZ0PxHnr
JY8gu4HVXOI/CvlstrkJkNehV10XFgWfSgwYjAGhppVCFnZjoNEOXth3I6dt7w5W
ug67CpDCyGUXkDldllnLU51fMSuU231o5DBE25d24RfDifvXNUfIIAGkqKbYjSWD
IB9e7prD2JANKhWNpwiTVfbp6hSWb/kZxjyaxzQpJUrxTPVR8i2CFJrknnbC2vpb
pvHi46ImXv3IuS+70TY+tyZvhoMyyfmD8OKlOz+AyqRxxXJzgTGw7fvAN4c+oBB0
0pWZHSgwrbg8RLtEU1UXqaC7v9HaKH5PbbeXya6wDTrVnRF2EA5Ju+LQzcIPmWOE
jDge+nN0lqyaBOUhfh2mtdvtosZF++bYvTgpLWwdE6Z3stbiER7OKz4qkp9EyrKq
XanbPdn3IbEhzMME6vDYnzE3t4z6LpLkA91Gwl+JggjGxHdtqRW5ytRyEvsYb28h
+TnKjajkE8zkm9+JufLlBRRhEjv44eYAhu1fYqe8DipGNctVVKZWEba1Oyl7zqJs
dryeSOEy+p7nk883mX2eM4wKT1Ytg6+BLTDJ47/a03rz/AO49e4WArNdD8aiKVDS
wPv/P2L2IP7VQE3NvnyTehpwLuLbJXndG3MHGVnjlu+IE/WPJOoTpgwQVxCKTa0w
H4OdKobQQ/fXuXnk63cJ4u9I+Uc2krPAp6VqsgDYTlivzYN4Jsdu9ObjBQR6mLKj
xfp5YoiMASHRXweGXFSoM6JynMbdjLOEoV9QMJNhrz09mI/DVRmE0aKM/flkCpLs
MpculwZvk02RZX6+t3jIwYQu7PvjqMayy3FkSrgcD+jps4ZhB5JE2SNjIglkWyJs
4BYWvMzK1a5nM2aurKrNDTI2OQ3o4GeUrLmDjOX9eH5ElA+3ikrrr9ovyMoiL7/t
QPR/E3LF3HZZZDXQlQEOkQOHDrRv2h+2/fySCDZrmocJ//GKnMsQv6bYHXvbyQCD
LTmAFdGrJx3vVAPEF9JqvgKSYo/yOkuZn6+5L1wOghTq4qlXvf9MzLexvQVKyzQ3
Y3EY4m8u+3aQUGEoUhiRv/dp2kzChiNHOImBy2L5ZbRIlnYZLOz1Qxqlm19ILMS8
itNBIWuCMXT8X7qCHBQLyHsmDso5DW8r3FusJRZod7xeryJWp0i6J2AYwQSShZbO
iRzlNxKrZ0kn2ht1rJ780SEaCY/IuTmQxqyEHqwv8RFmu2cguFwDPvNEevFnl3gK
TTeklyoRqoOarVRUZ18/8GScCHd3ek79yj+eeR+QW8pHOlAxNJ4Sw2YZ4pNuVudv
eVnn3NO6pOb84oQt+ucVnnXU15F2Phyd+s9yDvOSCezDdPbPOdwqpfpLle3clZnf
bSXGEMp2tCSkfedi17J4JIiGOZUva24OdB6izgngfunlPuZk+pnUAkVydQz5mr60
WPOxeq3SoC0f0xVLU3oT7yOgZmQA+ha25vPT61hzwy66vehow+EM8A2NFU2LrR3e
p5uTcRnoKQ6t7meLyuaUnfk7tpJq6ZLLk+J/rkKYkBxXPP/IGE9zcUDun8c98D6F
cYzN+EFg48kPfudXQpv6x2/d1fJBpWOQ16PeQ5cLhaR+K4WBHgPXkazZmw/ycmn6
PlDm4GlqUfvASVO4+l4DQcBZE65iXbgGHfejOeox75O5LL83+Y3WwC6YVETyHSno
+YmrvRfxvdgmXAqH0rvfOKKTyVRb+8nA27nft6eWaJMKfHugEWO5DNUxVzZOFjc9
DHqbSOf8tHdGX/4vbnfE31nNviAcNfMAOdvU7dUzvRB4gkscMqb/jSbJzkFdVMD9
/tlYS6Qzu6/qhQZ4Wy/jiSGFvGHLQozf4zNd7Ovuq79Es2opnE4kRNiDPi6c1pvv
TA7tFAW3tLUWNWYQkCPb3JAPrIg6G7AUSWaLIAzQclPLRDGzy94uXYX/Off6uAyv
1B5rlTX0HH/kY4JLhB0B5CxEGms8rEZW2y7Pj47k4G9P/IlacqfFBgcIXNaV4mN4
4+1ROenmojDNCXp+w4lA8sLCTNUYirv6MSW/YvNcJgjpRv2ocnQeqNBaJOrVPD9c
9P9fnDAXkaP0U+bb2546pzT54e5sjYEqvsH4IOTK2KCmuEWDqdIhvdshzK4hDatW
yYr2Q/AmRoHn6CmL3gzb9YIFU924mifDIUbLanVNRTTXhR3q1CMS3vXIQrEk3E1b
JhlcHWXcpyuaAcVcJqcs5zStcLdNTHECNxBiT4EPLpEvDrIBJUC5wmiT3T6gN1BW
NTHN81azJ2LDQ8wQ9EXNP/PPUeDucruYjFDj1gVsjBzmYxi+HJv6nC9Z/qWphZ5e
HHSI/j5W6NzUKBel0nt6BWG6ILnSzZArefpjeXRTNoZVH8vnLoDwtpp6P/QBlnKU
PNtrE9Fdw2bBdbGaCoKkIxB30KdrlSrOyj/OH/s4S6cuGqgbmqlqA5djQS2FPUYk
u1ad+H4sDY0SNJfxzthusQwoZgO93ORuLRvJmqAz1oYePzQoao6fTJ09ffVFJRy3
+KODADkFAg7qYqcOwuBuSiiarIYeoV6WdWqTTUojiJwoPojV1L2KbgDkjuVj7mas
j1GX9RkyzC2kdynxgsJUB9M26BVTE/K0AHemVuJxVGqbqMHXDkrvFRYEDEPXECSH
dsg9u5vCVV10NJDjPKEHQHXuKzu9E57fAGxVdzob55Iozi9KecjkJSRP6Gj7f63u
gaDeSq4ZOPD1oD5lmIP2ZEn/xNuR1Ja/K+zqq0SbAPHlsql2vP9LJBXu/fBwNooq
hULE7oSH/1qfeMqcAi6qIw1bKH07PhNLPDGqhm8EmcS6MlVtA3popGKpmhFp9arI
LUDWr3KbDOS5TBzcL/sZX+vd6aYtBgGbkBmx4DDMfqEAVV1kqArJFDdzgMnFpxnd
+/xU9mrp4A8/UVNPomCuphHjoEAj3FcFn3qNqWcqmXQCLiEELEMInhN+7TQ8MjyF
AzpjrnQOgmM69t/71F04GlY7sxq1BpVyLjKwQvAcx2stwd0Zh/Ecxkwi+66ayXXf
3dD8UYZhqf6Wjk/ucfqdxYN+qYawgCJqFsFPpx2xXhYxf9kbiveo063mAUskaKP3
jHUJGhVkVjTYJgNrGIltzwfoxS5yh8BuvM141U2Y064rt6/09sNw0TSQHDNq+w25
ff+6aLoeL2/rlTcWlwh1zgvyd1ryY+vnti/PuPhD+nh+14ojaK5y3iyUM6Ht/XuP
S8cC1Im3K1foCWHla6mqZC72Ti48B6ZnyQa+0lSHYQxsiNTv+ocP0bYrloArJCVH
mZYzfOp6gzGiMVU3mxv3dp9PvL61glj7QYVWqYMNWYFTqTnZqqtN5Y8vylOoui6l
h6uQlh0dDwh2yMxKtQG2amlgu0zCiCnOb+sro9zisa9IVIwJQZPggQyfxe9//e9I
TB4Y7FW8A1um7ARQAWhlYRcjunS+stBJOz79ujD+sHaaHZoYPRHgTZ++KK/8Lnti
Ilh4xsw3hjFajph3FcUugVw59Rb5+/UnFOINp/3CKrQAsdC0SUGFIFWBBUYUWy7i
J6K31i0Cg5apMugSvIFFl73znmToFnYexaQsEj0SvdRXGrpt3dkP4cusOq2mm6GS
a2JgGpBBauQgeVZnYd9TgCxrpym37MpQJX5Dum7n54KDBU261pOvZV4Zl+rH6G49
FA9K7I61devPO09nR1xfqlyICjbAICeUnEnH/GPdZmQNaIVp/pR2ffVmAl9V29yR
Y7sOBe8tIHJ1IXRm9hBRQBw5JfBZx/dXVw7wPzkXY4UMlovJmMzSpSZiJMJI+Zx0
QmIs+Zymh3zGTmA8lwHypD1Kx87qqw7BBPgszWUe2Hpmwx5AQ8Gf2Lh0WZJhL84T
AkUGEHziGRUgwNqMq+M5/drxMLp+QFmnGJzkbWkuAxXcEQzRtfGa8kESnHTRMqjt
6yd41UyT68+t/JStH+naeuU3f7Ed1WkoGMFLb+KDK7alN6gde9ul1/SM16nfDHKy
pG96P+9xJGERenRf3jufLrca339rbFwXOsWwzX6ll/KhiQ6/HEc2Zycxb/5dSoL2
+LiY+sJzwSpuDMBJ+skjzxTt0K24s3vubYxSR0fMZGObS/zStW7Cb5TYHrwsY4VR
M8AtC1J6UEUx/674bqqHARUbzgQdyhK9ajT1jQSxViQt84uCcS2tiNMhWb4RBK/T
uFPcAXz14ZGiKCFnyZFJ0ljVJ3++VQFY1BK23a2QMfRilZCTSN08Q33NC2u7EiAx
87qC4kvRdRx59p1Ngp0y3UsxhfwcLVjE65ctrvyTttj76eNh2QRgQBJzPyTM9hc0
XMsZ5obRzDLrNqLwkaHlMfZXSM4fZrvjHFBOw8eeABxig05iBNP0goWkAiQzmKtT
UoPkH1MJlwaA7IWGVDt0AUG0kNv5qP0AcKlINv1j8uNsQ/I8I/0vLuCDPH8xJJcn
tWXla91JhkW81UVzz93Q8Oqcg91DE3LBOZUjV6jHVkzYd8zteE+0q9kUIHcHPrvQ
/7dSNqNXnYQcWt7oLWCB8Yvkgae0pcgDsU2wv8rYY+YknGeigoFtWfPXRbNl8AyN
fr62Bq1/3OQqXGEjmNtQ4lyDJ0jsc5Hz4KcoM2vHnoCedoJKnX6RySZOls8xdxER
IlMvbVJN+/5bPVySb/jokhhrfAwy9O2UZ3N5Tr3UeAYldOxhuDMvPHMHwsuuHJZy
JVOuXUd2w6qFOzscv357cea5OMlRR9NRo6nVv+hZIKNXqi/y3PZWsyGbcwdmISA2
u8GsnKAjir360G/u6uCX1XuTBgc3+FLgTIMfAn8dDG8X97INeDPDdUotCf1VS3yU
5Kz5Ijk02JKjb4MLa0lVIF+Qqwn0esUvF/W85vjGWtod2TrD5IbacCW0AfQt9vSX
wbMVmoSQw1ScMQVFq6yLT0Mm9HpA2kvvASI/qQ71ZCgU756k7KgDwel3T4v7kudO
7LTCmBD27MA2yhoFHbvtwXcovK/UiE2/nM27fLFrqgIeLX8e9vgXyY4ynoJIO1pL
DxScBeKTzmnpO3FmIrhSiP2Kyzn8H193Q8zaA5EmAVY3VNiYv/R7oOC9EJ/jVd6N
qcVNPKqwn53jyvwBtyjAJARVqSPeNEx14m1D/tu4pUuyqbNXgCUgpBd05qyIBsop
XsOcfzLabEluTZKv++svwDanfX8zvQ0F0sNmdT9lc5Wp1+rFU6LbGoV2a0dn1xSA
L8XMugFb7cj/Q6Zl/c27iucYCmN0Qe/tBiSPOxYEfD3em5jWPUK5BNHXowwaURcC
eNWZYKeXt2vDhpXKuAHC7nDQc0bPxL7ET1l+x4UAm3GdqsShBaqif3JEa8yhcp1y
nCb78U0ECUxX5hLTzmH5/pPttfa1Z8m0MuF3Qp5S2I7Ua+1rbbYWtqkD7GvbNCD1
XlU3ow1XZVTPfc0wwdB+/LoSuGTz/3MeiJOkIvWatXy+y+DDsK5qKgrKCwismz3K
uz0Lu61uVk7HIaKBUk4CPkpjhlG+EQKENVWub/I3x930tAgKsFRPLfT+1QW/Vd7c
P07usjBFaAvduyTER2njhsZLix/O+uqldqr6CxT/m8cEELuoArDeY+R1XLXk32iJ
eNjxJkazEAhOmHmtC8X/4vrjWMR3iwDMbxvkP0iFrAhlFjTPHcLibZ0mMO9tRRS7
FtBOb+yNGBOSyW/ZJmH1iU6A4vl+wm3ATJXnwhiFUvsL42huEF85sxeUvENJSG/5
p+fzDGe9Sr2UHh1kC3oE255JIZsagfPXbDaNYDKWVCULImCfq8E1OL+RbV79asKA
GQfQPV/Phd9gN9ZCDUbxskhdu+Ig3VPZPxBvm8ZTLLQSzmbOj+LmFfW+RM+EJxAM
iuPSRF1wk3mdH2x+stl67Kya6jwVanuV1+2g+2S52feuqMdlHSJXeU9fi1GjNlfA
woWF6YydkEPMH+cUwcp6Tk3Sid9B8DvCz1noDsf/HW6PboC55sHfq2PcPJgpjFtM
/cpd5oXDtaxAZQTDAaN/JuRIL7WvdZSwo/XtIjWYsLoE/q4/rA9uJsi1K0tHceik
5b7McmFJTuqNBySAwB4GQmIdN0dWA7HU1oju/S7VmFyvipnaf206rVdHWBMZ+9B9
Lsoz2fhD7RulS1oqfZJUh8J/jf1eSCbMgCy6s9YhjK2nxKWAzqVKczI2ZfdGq/FJ
kmyi5DPlahp4NCMpcVyS/kOxLwp0dyPuOZll7lH0AvQIpondjuSI4NUjOxGbvPxp
2xoIxmX+WKPy76c8GE1WhnVwrnZHZdhVRD1RT8Bl5uxkDlroMtk5F99lkQO7m8bC
Z07ivm9mJkaSA7undJnTje6/XGiU9g5+mMiRLrVKjAtBmJyTW/mo2z9gG9Fg87v+
+KL/ZKoqA++X7L4VfcF2dzQ7AVfT4xeOaBGeROxatK/NfJFBGg4H83aZN2YK4pxG
1cga3zSEiydRWj7EQ3Js47RMeXXVEGD7Dvzk0fTaTnSTCdj8YRNZQUqvOkoY1lBS
6xzhcSoAxZvpAPhFBP/rDEPrwExuruIjR59fcJVDG1qazeanYjDFxAAQny9CrHap
nO+BJbQO4YWPmaUBDDO2ON8TDFT6hD+BoeASLw6IYb1Cp/Dal5LUYy8yYQHL7e1y
0Q7xPhYnWmQkn59WQDwax/WaKXtzKAWxR8uxsOO/uB7FjkIpcW8S2v/Eioj825Ne
LgokRCqHWaSuZGNxP8Wz4ePM53+BKqZUAGAVzfk58uJKeZQxpNRDkRU22iJFIsIR
XCcmP5uUQuj70KyrW37D4KKFLNLSKV5DDQXgwbVxiZjVVvJPBq7ecq2X2eiNWfna
rQZmhPb89aNqS1Kr22g0EcEOKxgla5gxrEwUx1//z492E4Gw1ohNkVH9dPiM3eTX
dFCH80W4cE4dc5U0tL93Vvxxf8aDl5LKqtTIzYoP+KY5JQuo/zTKJmBhZnBC9HnR
KqJPFDjSAWMenI9Y1UOUc3+5QpLZb94E+JmRSw+3VMuRBkcehBsJJWd5FSVc2iQY
h5aTNtZatjvTTCkB6uUa1IYNhgxmbgSrqMmQhHTtPfuGZfU/krvgdhXUo5o+xmGZ
wWQ0c/PMj1Jo4YbqN3zh1IJ45XEn/invSkjqEnFzc1TAuq2d+LLjnu/aPWr6b9rc
o0rxkFDEd3BZH/duH8M5UJN1mTw/NzKUIwM4LzSR8hoyrymS03orwgixotwKvsEl
nv1CX8ZT+bOV6kAt1TMYnVzztblpvjUa9wY4szm17a6ggZSmRE87ciz2ixNTLcQi
+6mUsyHE5e4vThBpQBe2tWl2f37Vjnv/JFGmpqQsC9bDiUjGMXHojGlRJGeTuT5M
SN+mhN+/FoURM8gb898L5FNR8effaKIGz8EMs5Rp1WC/gmCZStBcNGOS4OG3hrYh
CJinva4cE98TPuun9jBGa4Faz+VJ5LSii5Qad/bJ7g+RD2LCyC3KCI3bwRw6VI03
Tegzqcg8ShXNyNupG5H6SV58CQjbq20yWWGFyzIvnum58mgCf6JHrTdXchlojJEq
EPF6a6mRIr7CFNa2YSe+Do1oy5O8kHFXsUIWtWio9OsoOQZL3X3cykAvmeDFOf7N
OmilSfrddisXQUxocbbV1sI8dJES84AYPoAo6IQ+Z2cVwImso3+3Z7ct1iWzNcEV
H3dCR/UeT35C49ktAVEY7QldAFwSwQOLDgc21YZm6NmwhvgXaLtHMUfA1B92g1nD
Gg3VCuE8+bEHcg9HhGGTxun6bM7gVi3X5t8gIcyhY6yV4ykfwOgVvIllm2KtVWLh
FlhffG9GaCGor6n7risAzSYDF9oxnTVRXA0K9rDq9VHGdujZZ5h8S1ipDMCDvqDt
EINRlJFg2hBiIi1ShrTNwLDLcTfM1jOF4nJvAebBuN3D83hhHz5Rx2zwojBYTw/s
FUYWO2/3HKWUyswusVGjFf3wiL5O/UfmkcgzTLSnrZEasjP9lpDv/eTvJZZQYAKp
CyXSAEZrz9I1taRqKMODbZFmaubEJajVb6MZf3zPzLfVYqaaS3lHul1fXkMZzWC+
YNxNwI9LMGAxQnj2Ch1gJB8IG3JGhEmTuJuCwaLWlOeQnSQtCorJmB7+iblrnE4O
S1d3wK7RqwnAqEIK+liywGeTSpP56BF9VYV7s88/6X8+iiZoLxactteP1IFGHxuf
2YCGGZFWo4VW7f0DuSRjw7AbuBnWyDJTRM9Y80fts9I/xvYPlAeaPEZaHhAj/HBB
NuJp88zlUzmErQamTsrxvVEqVB61IrnSv08WYc1lc+CerVpHk/XU2tXj0GWQG+iG
Ft0gsxzluSSR37GRa9q7uKGAl56JlYMHukb2iU7R6O+1GqcbDTShh8VD2CeGvRG6
nZ/vjqoFcV4dJC6XUSEdJHGys/wkcmOwNIX2UNcJ5RC7oA71RDiq+dLfbcYnLAS6
iXcXvWG1iS9ogi1gMMMNU4Dx2fhoaelJlSQJxi7ka8Dby+YI4REp+U/dDrQ/I14q
u4VuiQjVb8PQ2VevQ77ibO64SJunYv8GYL2VZHyX9DkMpanO0ze6PUtOo7vfiWT6
wccZNu3pQkAfks75R1or0yFLH0cBZER2YAyDQ6RvG5Du8iK7SESNKxBRL9M1nTKB
J4IufuulT977rK5yCeV8s+TE/1E8YdJ1UqIkvEFxKZhnl0cnKqHzMxA32FDi24Ng
GvSEcz1jwlXRgNNJrF8Nq2WeV9eLPuJ+OM0qBy4v/9lY4h2CiLQPLn12wwmwVYgv
o6SYy4YtIH8AYVBBmz+35sS00laBFt3toUKjiCLLB0jvmwcUk+pV6E+GC4XnE0MW
Wo0ytlVsKgjZH600QBbG4rfXJqJOkGfZPgaQ2cYYLMrDIooOX5iHmCPhIbrqxmlC
3RXmCFypieA+4zZUYAeV/DebC5vIfsXG1UHknVZ+7QNRNKhKkJARaITkLDmfGuZu
5wFqMEgo7gh0+oTaPOxAGr/MGkaIxtzLd3lPufsaXV/RXDHU2a+N/prOVTC7sNKA
vRrGxKYP9lVuA8OsQel1Lz1xTaH7Gml7WQoXfK0U48sGJaCgz9XrJwgFs1pmOh3p
eUNECY4CMZREQGSOizmPR3cVorO1jPV6hAeL6+jbQZFFbbe805fETEQpHSQyHzV7
L7mI65sTyj8uKiVKom5ctR5IPiSjJ9iG9sxp0ftUB21+34gyeddyEhPoBFgaE7z0
HOMFKsakIdRwyFFqqgu2lREflnOG2KuIXtQ6l1W1GNPLtBTng8vk3HM+ZMapUj2G
gaADDBYgYniY3CgDdNiUk/bCkU2v4tbTSyMLrnNFZMQp4nnc75AroeU5J6DYN2Zx
O309XEU4PsekfGL8DbTdgQr5tAPBqhGRaAob/PxEZdf5Pzg54eh9tNLq6Q3Gbvwj
a5hgcA6b/39QCifocZaGhCdknJYvKUG3AqUEnCfA8gmZccmiUuID9BuVllnH71CP
UQMqi4TgQyzTYRv05HeksjREW51OeGSzH3PhRfSJ6yWqgBxwZYWcSrbz/TWu4xrS
I4xbg8Kiefkoqcgi4y6FAJawKvTRrRudHGf0mUMnNwfl1LFn3tDhHIZzeor/eKYv
IbePpMM6+ySHQMbwSFCEIguhkP3YNkQB8ET9YU7ZXT1nr12fhK0sHhy7MbqOUH8g
7Z8PEHfxxG5i1qucFFVU1Fd0lT0mPOzLEoQofueQuxobGC+H8hC/zxoLiiPIvB6W
5gcipfbfcChtHIAl1AhWUvfW9VGUC2QnKWABeL8pOcNOIbbOEycezq4FlJ8wnBh1
zwqujKtiJTTOYF5dTNNhzMPg/m+yh2HDpfbiVrgcWAUb9LlMYNdOqsMwWzb1HIAv
Rg2XM5MSw+kgq9zgb9YMYaEKObWr57T3VfNpkPtND9P63nz3lBOmmxLuGDF09tIw
LlERpEtumlIyxsCa8npTMz2ktc8Ks96/E3ykx6CvkbWFos/4QF8iC8PG2pfMa2/1
4netasU4lFL9Ts3gN9zOQ4sqZKH/PPRBAlhMqd/crdstQGm0+BxvTTvmxDGzP/ZX
w/LFAa99WBn4ej0j7ijyMGmWyHsaYUa4+Vp88d33v7DL7z092NbyOZtfIFRMwuLY
/8E7F3FtUre+gj6I+HkeUOqr41iP5V9761domNd5AuwOiMprVveUGesm8UGp/qGi
GVIA8v4x2EsU2YZ16oUW7TLED/rbhFMqoyMhbpjTyNSVX/gysFNnksM9GIZ3kFvM
mhRogQCoMhikSoMRaApRs/sg8XkKfJl9JY1cEH1BYjnfF9Gwwi400zxHQwclt45B
3Vr26fwl+cXX1UEqeiY4taA0Nr5/51zGc1WQJe6RjZLpLkb1XlkTo6Xc+UZrAPfw
qYCGXtJXQbfU+PTERoSSKlY3JydCU073lnx4U/xplTj9DhN1u0QSI8xfEo55Mbij
aeXKA+1RmRNhcEYv4X57uCbI8e4CrlqZ5sZAqRu4/lYoKl5gD1MLtmdFNegYBTX6
plaUdesw7rEO7pmDZU5i/B+Ixlbk8t8iLnWpZeveNgOuOl2m/NSZeoxK9+fm60B0
C3aGnHEc7DJTZCXK5+q5U+3TypHaP+AKrJy1k/t9OmbVAV7fJn4Mxb6Yl6tjhNzf
MrDUo5Z7IellG9kvJ4po9koqg4y80ZTQ7Uw/Quysd2rVXb2/zpRBT/weKWizFYpk
ML/VdQu5/8gxqPp8WlJmxRgUCUowUXREtOQfe0qL3nvs+onc6GUm3GVxLweg3GeZ
960aV65zo0BwhCm3o8sWyHZwpccWvKfzLDT2v9557I6g/3lodOihRx7TBmITIf1j
/vhjbPzAjqL1u5c/9xUYGNvEJIeojQAOPA+sJe8EFiOpjPSliBeUJ5ULvHQiMqKn
aJ0IBEuroBRM2Kb1QnBYnhRQguxQOx9Zn7pTu3FXKdhYUchNUMBHgqwClk3Q1Bam
1wcnD0LefPNOhbajii+/Lsbfbt+a72woPJdhHC4cmkzw3oRJjou/QQiKSn+Uktn5
LCRQUWuEynuLFhuwEtx3tQuWb8hIJbcNA3Fd8my2NpG5HXq+Mhg0faZ9KW7vHaS3
M9q+U67JBhisJ/ymFlS06uaiMRdCxbAOjqteJGs+n36mhhkMtQiZn/cYKLtqOjRb
b553XV21DHTB1Qcq4VvLVJmrzvef1qk/3B6vNXTA5yTTlPrjYNOxzbZFbBEThXLm
X9Y0DGpaskeiWBx+KCDBWQlsSDfDU5cpiK1VMQlotLhh+u4w5TuRgfdNXdCo2y6l
2UFDD318J44t4BMbsTr2dffLd4Zop5skXCbn4XecW54E7JMNdXFifSA1tf1kuoVT
0pNn3jmmYRsb2qdpxoez8CBm82ltgf0FuQy7rf+eo6G2GR5qykJ3BWTS0Mnt3lq3
nRA22ktAGLLKogkD+RaPHnVBoRMszmPcf2bCEXObwfmHknOJgXuB8H+Eg4TBg6gm
K0UDpLU5mgzXX6rzWLQ9D6G1x4G2EwzRrozM2s9JiYEtalTPInzuZlP9BVX4PhVZ
R/4BWlYgxd2TQuDKJ6F0+x8U+q7KINOGgHHn8zyYCMbgpBtHY6VHJclUoErLtP7w
vBiM5IDF1ZHkmGDlV0lkkiP+1jpJYcR+2xKVYHZvRKN1G3Lnklj+eWNV3QiEXxAT
+d6vggW0f6U7IixLXPY7LWdAhnghDXWrCNKSpkMV7BsUakdEvNc6s5lMB3sbEPD6
Yh7mHtyQBhLTD4r5/wLl0GxHqyqa7DiON0U3oSTTlgpdpjv/XucxWaKPVILm/pdf
yUWFCJRjuL4O7J4D29mer/nB36K2J6wXTxdcNKHFj7Qcil8suYgEvO9wRb8qr8dD
m/KLGnW36dPyTT1vLGKN9nImmPwJwtdvOxl+n3XoDVkRBVeO1Gihe90k39VB+QH4
M19W1Bog3mb4qIAPE9hAJnttou7UmQACxMzZTsJb4PrNOXqqR7CsA/S4uEmmFgOz
qwShmBdJw2OxHvSk8eTjX5UMORCOiG9iJKpiuqMo0CZvi3aX3OiwFQb1EjQ8I6gj
2pkYjP4r/svYg9C9tFasxKfX/5/eomtjOGuyHd/Yf0ktvk1oh/NgPTeigWaG34pR
jzgF+Ja/eMRwV8xsdk0flMTi2e7eC74oncBcmRH9jOUkDDmObU/pmC+zA1WLu3lq
vjL+bxcdwyBNND0/xleI2LPSJwywh5wEXUFXFiN4K9oia8f9gLB54do5pRoG/i7g
fyBnUWUpSAFK+/wrCLSjhDZjoPaL1DTZX+Ry5fb4pSSUuxCL+vgznpmFv0YeAmw5
J0IvfusGfDV/Iocf1mpbIp42c4ITmkhBz6NW+5apNSNoydvAiqUD+HplNqBTgFH9
xvu4CHjDPoCv376O+k75ltrqxiXKvMdtvX94dDqhEwd5KtJvAnaUfNyMkZB/5o2D
ShSGgVYQY9xhGMT3Qiebjvg8ptS1Nqo+gLQk0CgaVzn0iU3t4HHQY4KsNa/Rjgy4
rYUOpD4VK9PzMdoFAY8hCUYiYYc/9MeyWCKS8b+euOzpUEuCART0OkJ5Jts+jQRT
aHusHpYcfgylbRRYXLnlczpmlSnIKQ27oO+iwT39uI5kvf3nNkc3vf4totKJD9yw
5Wpep3nO/O1RKBc2CMzx1sCUu1mXbp8YBOaKdunTIDEjICfqkgG64hqbbHaTjJqR
5J/SQu6mz4PtE4/CGjEQg301tMDc1p6gmf0ylDe9dNYGUsjbmDssiqrvGzN1EMwN
87OZzvHPZW3Ig66twDz9QkDmeSOdxsgzi1lU+wrtk/Yxc7ZAoVvxHESiQdP7fjdv
uSQpRtM/ogWEIs/k59Y/Jqy8fzhuPC1Gt3c/7sYrp4b3a6HB9qnfqU1KlA52gL1I
b1P05hKFrz3CCSKK7KN8/TKSj/6i6G9Zez5bQOPE5bwtNOvRTGmARvXLIaReS07J
peRAJfcNx3eXLN8sRmfcleZFfyzqR50mHLZUiFqdCChLj85p/BCHDc5InQG4CI5R
9sf0NNbAEexMOWMAAyo1+48OTAdUejkGmd1zaZP1lvuMsB+g74lpVq9LIXChTCUQ
U4IFR9kksu0oaZPrv+Pc4GryAExamn3uZ46AbxqnyWIOSVj7+w+YBT44E/Bdo2rT
faWmBphIgQwbt+3g39BAU3fwWo3s75d64n3nQVb/hoO4u2kB1OMEyHd0zfazTwd3
xnm7Q8pbKaEAlQRmU79nVX4jTHyIOv0LymoCU7PJkNvv9U6jWoUxPVL8UFhQne7f
4WFRL5wsTJGM/uhtTi5xvZqwLzSGMmlk50W83mhtfrHSX69CqWL/EK4cq7XbEyYW
s2hlzGkMCEWMpOBGaGOi7j8BIEwsPLFKCoH0/5gm/KwJQAczY8uZPLpBPz+2aMKg
hJSLpe3egOagjHyc51hnC39YqjrtWurCVb+ZSVSVFvgtdPtMovgva+H6B3ix0TLR
pyM90pVPRoF2436vZKd128xyc254HwdyxYX1P6pTR8RcH5Dn3ZB0Si6wpGykaOtY
o/eLWum8IL3BFsodU5kd18VdVdRtUcPfnrG0ZHT3ND0uMXtLvvzjgAX7NoERGODZ
69KIhOuv4GL76khHQwQVJmpSBcuqMiDS7ZTLSuamtj7jHz2fcPx09U3RTRyOmjFU
iNLf5R21HjjA3UFkdMfafjp3iic3QBmjFwsoTz+776lh47NPuAwpJ5YMT++QWV6l
UhCX58KBZ9EibCFjiPXczebH/O+Ni7y8t8NTwhijSXp7lX6beqkPeVuull4CuRfv
YMvik+kv/cftAEooCNNvPXUqGayYQIEL87d6V9OSjx++2gJF50I24eou7oyT8Z7X
DPPmGQjUu/qJoqep2rMdMnmQbLRGPvUuQLCknnLJ9J2jb261BzSJZJ15h9bAHn+u
TVlpz48CfyOkHdb60ouFtBGPwVB9FSWB4YPUxoFqIC/Xnn/Hk03pT6NI4AGBwRM/
aHXDf9PqSZG6kprnf66h4jo1nLtqIo3wu/fTI07WQN2sRUNHiNk3dsCu2wFQrEe6
49Zk/hKTf1lNPWFaquvqkKTfPFypYqnlauLgDHeZ3MuP+zQL2RXRpHe2uNc6ETXv
NOUQYPZmB8lMJOhpRWDARWouCs4cPSukFy2eQD+G1gUVnGDR4qk4SjHK1LOWDRnO
nOHHdhKJT403Sp4lQhUc3L3g2Nu4FKCSeqPBj76L/rNrUY2YehUj3p72Ol50c5wk
O3hJWayogET6+N9Xe+Xr/zL0UrDslH9Cbzn+2zRh/n95PxlIRt0QjnZCPG7/bg7Q
k3uKB752d87Kp9W45h88B6N8GyEGsR2Dv4C8pBeRKqG4e3f+8bGaP7NeDAod+kcE
hRifyRIhDjYWyQ5cXO5/WrlJfxMw8zSf0tt9s5pGrv519v1nJhwRvATJa7YM5ZZ9
NRW6lpQ6cT6TbUIVwXaEf8ZYl5FUFCquf/ypVJ+PPhWbgR304Wxx88Z97QcPlZct
whzS6A3gNQaYkTi3FFwZ08GJ3B8uDIE6ZxG+/iOfgI+oabMedPnb33J+WmHiZi92
r95ClbG8Z3lYoqZOMf8FJ5acGohnIoQPGpyxIKwWIYE68jDp7Ovw8BnobyrUX9CH
Ad3iWfmukPMpawPfCsydrVodz0Ei/P7/w24/qLK8ineQ7y2vFVOrhGLBMpbI6s7w
oyAWH5QbaoyLf3c3gsh9zvBj5JYIDCzkGbpDhR0BaT2dAwhBkbuVvjE2jPOT1bmF
V5ReAta9xXuTte16dboRvFZKgIJ3XiFLGzOm2SVmBG8VrQ/qUJOncv5IRMN1H2Ia
sQzhE23j8BZkGc8PokTCKrKTB7hX4uEh03cUvsyJtlQ4NJZyvTZMn31fQKUh6OW7
G+pJhOwstujPdITTJbbdzreiqlEYBxOMiOWchVsIxxymGPTau9QlUvHtHbxEyuvt
9f4ipWhGOuU9MnFBK+3hsTcdfYRAF4kB1cye/c3fTPINgNQ3WslkbYSpnSDTXj52
N6CySjowmk2JEweTRdtZSHlZZ5CLNfNMIUlkWRzgUT/1jBA4lP/gTxAwZq/LclRE
tnPnjppy+Lo3X4jzImg2JfjIalyswIbJYhaaufov9prIYK+8Z/DN0Maaldv6ViRL
24wRy8lTeN9Z3dhJUROq3SrEaxX/kzJPKjH7Cf81ShzVdSo/Vu+Fr52CMWwJfxaa
jC2jovwaAZ8CVS2++KuADwS/Ge6hqnc0HUS8n8hsmqk/UeGiMEzjUQ4ZzLleVN7r
hrLaC2a5rVe6sFaiCFxVUmWTm2XZoPvf7cK2t0n5pBEG0rs0ANX/1F8kxG9jF5Zc
PntH+mg3ypPZMdFoPcrSZyrrNwusUx23hKcZdj/mn77U/JdXheWMVu4yiTwUmn2c
mUOfM2z6bmXQHxBeySRZQAAJ3FbG2IqgwTjF0UbNWIFUmYdyAeuIzFkFWjevWPJv
K1td+GayNUr+kiJiyHmDEX+f7dzAEdH3Afu+2xTgF8WxR1qHol0slyPBvZmbtkrd
DN+20PZqKyXCidldwrmfcZUmV+OwyRDi6z+mCAz1KH3raXg8wiavu6zOBmRQxMz2
dz7V7LkhNfmm0cxpXnzHLOS+xFfDBbmK/Moo+kbUmIHIsj4XWMfm44PprMB9sU+F
ZnFz5uI+5pjvCf0aXD0fM7EUeCC0KK7Y/7HCs1fnZKgCXkgVm3/NHzLT8mxgTWL3
HNhKNhS26yMGHQxZ0dKAaTxp4RbL/HbkZMhIkX7mPi+YGZIun9dEgQNv4RQTjXg1
5mUdRkFBxhUsU67sShOlmkz4RYLBGXlsThBXnKMiWupOUmZmBC0yYcrIV79JrAXR
G5KPRQIBorKXNZaoOF4zUDFm1QXNg34LfGadFYIOF7zOg3ZYmVyY4mQX6JQ84T0u
H641FLEilsHJj0QGSbV3a6RMpkXMjgsZAqXqPFq6TsUmiA6TlLqCI3inB31zpZxA
z5AfPBSyF/oditN0NCUJ+9vKwWkgf1ul/p00C2zoFhtBTTdI826T8B4SyC5RAtEd
Cvp5fHikM7CoWn+PpO1YeNIeBXvbnv+OPjBy/KBKUVGYxrZaXHGu9qIt++cIQVRR
qG4wFNauLbqVzXYJhTK0Fm9589EwpsfYDDthS8U+pyYxUTH4yqw9+AcIG9vOAFzP
QMtrBdQNcGdNIp82KXDKQic5ACo5ItSauLNatGCthmIxRaPqCtgOyFv/0BWNkoLb
jImA3SRPnIpCBQ4UNipXY6rjNjbDut5MEloQIpurdzORy0opTDHslmc2LYNflXsh
mVvOwSEd1r/cVrJ3ywY2G9oL4b2BFfUqZyZx5gX8TF9Uc/LtRuvQskQQEHvsw9+R
5SZmfmRscEphD/Sk1adiMuv0CLg8bv40FvA3zhgdp8kPlqrjnRgcempM9Vpskv5d
pHiEylxk5bGBFYRQdfgKM4hXBRYgY59jxIYAZAApkwdziI8PjZ7upZkG99rqj9r+
0U87U10o74ABWVRmAdlHqVEiTuh5z/SGcvgs/M+I3/mqVYlJheKmwsSoLG/L3iUd
txQxw9UPTRHG4Uo7qKcYObneTKTUM1fuoes5zicVw/JfKz7kouJOy+0ioMD3QUxS
/EkLU13xN74qgx48NnfcGMXUPrUVXZh7thYjTThtBrPnAFvT69rUXYMQ20zteO0y
qwdDK+M2dXFMh7vTr+LSKKNHk8NE41Dm7s9pe9pXVSCZ5eFyZJpxm8cxVTogzYPt
LD4n2GadIA+/EfAxtG3OE0ZqjTyU+jP7Sgv8B5riDMlAKS+if97r1/zughkHAKfO
D2stg9OfynMDMEU+H/4EroGpzcrU2P1UUtmh7cF8Upuf19P36QVJcm4rzC+lPScT
bNsRp0uwhdcZOzsMpfq5Bvl/7Gv2mJ/ZGvkLwpH1qas2VsPsTReST3A347iz67MD
ToIPm/J21jk5lRsjA4hikAjoX9NPNRkjq+1+BK4cy92pf0WFgBUa+EgBgHNdm/El
mgNYbj28WFNf3ThA4lj0EpiwH5mxX9kjVszglINHgHym/NBHPbxXFJfKxIqQKa8P
HWxSVr7adeBJdmwfn9D110MkSGowlQ31cs9k0j6iXDzU9+f3hpg/F4l8E+pyHrbl
QN3Ng6bb1oA3ypuwUFG/qXkgYwNtTGZnnZshFrMR7T8uyZ7GPwpFoNsEfy0AnyeZ
AexwhfH5bKGNWLfFbV3XkkIJAgmiSMCufqYlKoipQ6hQY5mlGOAHpYsJGrrdTasn
YK4By3JynrFDotLBVu1h9XEKZLq5Jvkk+vx/ZIjHeH68hBYDmpNCFZdEcuK6Y2qV
sO//OlWGMyEoALgEtMDnsI0dgGO7fpiThJDGGU90XiQp10Pba57z5SuP2MZxqegH
BHbhVe9WsH7EGHN/AhWb/fD71BEyBAn6NZDP2nmuWpjRgnl65WVprl4ShCQkW8sD
4ipAFX6slK+5cUhhdVk3McOMXMvin6QU0y22He5K+1Emmc8zvB4hr+CS7GxQzUi8
QlAYE1RrH05Tymv0FOV4LhPCjPqQErAHR5uf+FSnYJhUuSND6Cj4IZgzgdb+liqB
xifH7kxfCtiNThBSbO3Y+usx+8uU7HsXvorso8WWfzCxaeVsHxHeSsRE0Oct8D12
BVqXACQLhBar0dM42K3YIfxxojD4SiDijkQLNqSWIlv1AMXq7O54kQa1CK/TkG8d
Jc661H9e9nRCffaKRQu+6met4ZzssfP2NVt8Yj00F+exa9+CKGk0MZJ1OkgTG5uF
UOMRh2P8lGo9Ce1xdudeb9SoHMcfCnijkgsgK1WVoz4HhcrhyccCGJNKGs+xJFyi
th+6sXzfv5h3OaQ1rzeF28qYc+IPN1+pgbae49Br6KEIbfo0WQaCvaFiv3dWQITj
t9ReZeN0RU6pDC8wsIuQ9hbAnVjlqDXR4kuNO+wkbc7zWMs5C10QKjDL1+B9FlY5
BJRmzxWwCo6oSgIwk+ADjDeaYa1j0SXrAjWAw7ko5mR9ZMhX+Q92os2H3SVxmo7v
hpy39bPUXU7LeqdRg1FYAYpHx0HoTxUATMhCZoBGZl8C234PduYIAF7Tihlv5aZM
y2Pw0sLbTyoa9R8WFTwQUkpSgJhep2XrKfSR0nctqpGQykDqQOkms/8WUTcQSSRj
iNb1myX5kX4rFZWt9zdze/qWx+DL7fe1wfSSvgR/ehjo613qo2id9dNvpNEumsLP
zILWJ6EA9fWofvgna7ZR+BIetshhwVkxpVSIFL5CeGXvlnh2l6sjq7e367d9P6m8
ZjZvtxg9WC2rgkDomCONkxd0wjyihg7anooVQrebahKi6f6PBCJUU9DTt/eeODUF
f37SRlO6XBzVRaG0+b9Ly7ySFH26f0ZikTA260rZZ3DVmiLP/cEf1cGxz/yd8Cq2
dqOKDiaafD866aYhKSF2CaQOC+ZTIX918jrc3dPQptVXBIGa13EHJoFmY7PW9qof
LXHBrrkvt2Un6ppA4UZK06y4fOrVIIBXr4GHdrqPkNnGmITT69WFYdkTF8Xl/4+X
FlzmQ2ysb2vA8bGB8H3e0o5St0FenciyZ4JEIJeVp7kYFM9aCaJII1ybIu14Q2si
Lxge+loJsw4aES8zVFGxntuGY51NWTvIthpqA5vhxLTkAI5m44Y8uQqPbacha7Dc
onr4qAI/X/p1qTKAPyp+HnPLShzWB02Ga2KdA3+xS48aNAeP5vV+pAeYikV1Dg6c
Gxou8rSctDBkgzAiMd7bkCo1q4kORngtLnOj/pCdzAXw4lPCv34WArLAhaR3jG0q
4G0IzrtCufYUAsA1/Ssx1KJB3xPkPfjPb2fJuR1QocpmWXuCOhm7AD0SWVIpSmh1
qvZxGHA2aLcWRVq/PbYn4SrZaAvw7hQ663A2Zi7C19cbPSjWTfrHkEM/ZAbwqnmn
w/UWFl/z3D2ja7uEq3o7y4jvQUPOrN4VRmfL9aDL2S0mjwxP1/VRreUFlYHO0yal
lSChBuGBgmI5MrZm/W9UCI5EkU7jvtzWgyrbjM5/RJo6JW7QiGAixXF27RxrGncZ
Yo8kU3RCPX9v6UOTIiLEsXKM8ZQuHy8NyerSZiDiEAZGYFMKZ0sjm9+CXuG+biFq
HkPOumslTM+W/wKwH2GjS8eunrYWX6ya4uC7vKgBN4GAH0AGd5Ik0XwA41YDs8FK
1eCMYesQNF6Ry5Ai33e+aNM6EkEH9hel4TX++zaRo2STkb1wtL3/vROxNAxxug53
cehLeM5fDNyCnOvon3tLIzdwmHvQVsxiaSEVcBzdZ8audH7HUDldG1L87dEqXeMQ
Jj4fU58zzlRfr9DDBh60+NVcZFgugJskbHcHsF9GY/fwPA9XDxt4oX5jBVbrxWIP
hLiinvCJS4TqZcqPrL0G0MOtLNIncLZrJLIRj2wjb46k55afpOsdUq108PM4AdJG
zzW8QUYtxQWLr25NR30dBa5j3bPz8PzpKZ6Vh7utXbNTAG/k1rUmf+bDpIJ0x0BL
4L7D0GLwqmI96ddDoxDeikqwmDlDMChJhqrjxIiQM8fxpWpRVFmgJ1pmbrdyrWbV
cz6EBh9EdlPJX9wc90GrllNbN86TZ7b+x7inysppJn7Gok3y3gsh89JxJetfBvWf
fd+GVGh0qIOtciSzv3uPVW8abAINIaIiYfql5ra9xFxLhH7SO5R7R/lla5R9fDfZ
/btgHJVZTEATaYMxJbbKHnYJWi4fOwaHBwXXhFTEaIBReO9QQbVMNPxEEgGViOc8
oyZgTicQE/zemEbT6mS7NvELRSs4jYglnSZnQqnWqIdKNg8ICaxBjmWg8/TchPL+
E71VSfneBqMBQrzm/6YMzXlksoq8MLCqqiSY5Gev0Auw69Ma3sdp5O4CFCyT8bTG
52yRFGN14UKQXXSTEL3lWBuuIMG3+sUXvVVQG/qm9xYopnOdJCCjPZ6zxVfa5KNO
bKvewj1Me/8PMhwQo62mXsG/11fLdWN9Zu/WErOMaY8fZ6Yt7vStiZ3dU3MOroFl
my8bKbGjYxo1QuBxrOei2aj/NQwx07x7gd2O6ngfdvaww8jjoGN22b+3rVRrZt63
FE4hWwYivwqHy1ROIq4y1ROh3C0SsfBY9R/da7OuZJftSQCurNptRelJxCG4rPHn
1eSipRaSUrw2ZKR+lLVf6hzX2QaXid2U+N8EFyC1Tl7OliFXT7othz+nDGhev7H8
8B8O1QKATiq/b4N+uqbhpUyhOpAoWqoaJ5vxra4QQLyCfcq0Pv5zBciZ7KuJRXhw
Yr7KrDqWrq1jt3fMlFj6XS8gkuUfppGq71mz6Wuaeh2KJFgNPdIjoUTB+uwl27zr
HErE4b3cfwpFaLOW/g+EJGj5bLVQ3Li8/xtMGWOlHS6VFLPQBwYh5iwmpG6kgMzr
gQZExUifzaxUFceUb0jwV4+EfkIGFrMOdmsxOEgwer3GqoJOZY7QhAxYdyrYHzpe
5O/oTF0fF5k+WFhtBVZUQ74/v7Xi5fzVm5IwGFHPFl/z2zeiGjd9tpKSNWCJ4NYO
vtRLhiUcaVR8I8mxCCIzo4ivpdyXnaT1nOgi0iOd5YRYNNWP3rLobTqA1nUb4Cy6
V0DWIP54R2ZaqrExsmpRmMWpwVydE/Mln/YlJnYzO7Kgmzr+PwUNCXcYNNiZhv2E
tNiPUEdbfRFK1Z04kgtDQBXdXPMz/A61miVEkw429ZjvzHAP02FbomAN2Nh1yLYq
m1Xk/qvahC4eF5iaAPjmP4983crw+xHVWRE5rxaqDHoS5jG6tYb5JhQUKEEhKwu7
ZExYdr2g9SQMTMrh2l6NEWf8TAzhCvxQwHkshbF82XpLqQo2kJnF6eWW4nvaMEfi
VlRrq8QPvpDW4vu5/HRB0YHSjNdt7J2Zk9S9csU5mq8Co5e358+wuWqx58e9xgby
5y0i+L0hl4IPutkXdRedKFx88cqjtlpCTgjwUj5A0ucOVB88NfwrsdnaeGp7vHFl
nbF8stIsvlJCD9uIT7LYrQDuqdgppoDZmVLuzvExuhUE2GNaZ45GGqdZXya4rROb
2WK1KsiL15hzYleogNIJB6NMA4+xBK9Eo612hCOwDIqjWA4MxhTGNI781G8SI5+2
cHNvc1+ZVQU3GhHeHskNq7Jgf6b6IynmOuesJhDcabH0oZyYruGCDzZftsd22Sr5
bVWl4AdgXJomwoivKFGJP/VPfXR0xh0ENKvxZHpxx7yO0teRRKG34w1XbJ+uRa48
IpCK5hQMh+jLsadFkCQSb3yBhT9a9VmMYwVNtsDvOMIH0wzZgdWRlL25/jDRk8ZT
kbsckdYYpz06pbNhWQfEZKfgZcZ9SH2ssr5Wkg0FSU3cL9mvFMAPqm6b7SuXDLAT
M7rCugbhJFfn0GKi+yJAsCd/C5u+MSoUMpa40ffOs8SgPYnZSLzH6Z4HDo9a8QqT
zpu8YLBZf3g/9/p/NM7W3FkMJicHTs2ZymUJ+SF8y8mmk3wTHXW6WyWjXqmgq5LB
jDEs/1fStFxHlcJhn1fCkmjsMMf94azyZNwsqfupBFgE5zKF+TvD8VlqbrqF9PYq
4oIv4y6KGo4Xf9g00nBC4DP9I/6IZPE8f4s0ETqmlesUDD0MP8O3X/Wn7P9gCie4
mmPUo1jLWzISnjCj537bmKD73T7+5RyrLx6j7Z9vK98BYBAx38Fn+Q9iBvqVPCJP
WOTaIVfcuBTQCpommnPMt2z9ChYuMwpMvPAcJMD1sflWrbwHMWbeBRxHasVYZc4I
9bnPkeUTMLbCLEdBwdJskZ8AMqpU0BFPazqqbEYNfXsUodTCXAxE28NOeCSdEBJN
sUPfjcxikQ5mQ2+xjhR7niLkwuGxeMWNP+o7Vnj61Nt6IgBYIFjK+p2US6wUKJJZ
HDZQlcw/Mj8GBIlLGysIwJk+k1u3RWpTxx8nmKVnXfJs3IX7CzGtor15Fr93ZWgO
SRmABsMtTFR5sJI8CL/jEJg9V04eNxJvkVxkTULEgzc4XgtC/MDMvTD71EZZRriw
QMB1HW2puQ8980WJmVWdidwChy5iXoFhhsP+iwHTSSbOHye9nGnam1Fw5Jep9i4x
UgKebMk5K9JhZIP0tgzMYseazMLGjPzNOFfwGNtCqRpD5Knj9BeNIIMVNsLD66nI
V+EVZMQXEtSRPRsM3CJdwe0HstSDCLTxT9lYARtAz+ZummxgQQtVDNPOTXrg2N1x
0gLrcJEaVsxVCkuJY3ZUGQy9B9gifXguqG2r4aml5WE4j3OkEyhgxL6dO5WkEHAN
qbUrAf/6k/7Ea+oCQlrXitF898MlaLdCmuLaQD0rE+ucpuXc/ot0Oh/lAf7OaI4p
2B06gpgrzp53bx1VdQke5CHfdlE6eWIhRBZX8zFi4FN0EAaxygdOVN89R92e0Gn8
/3DCkI1wYkClQUK4ndMCBlk+kQLh8uKjNPZiE5FSiWq4q+3r/2VvS3M2jwMJUYwc
uu0XTPzNjQ7WwZ3ZcO9h3oQUMsOHlPExwnpE5ztZmDTe3Yel4KH5LDVxQGOp1cQR
CzX4lNpDBqc7ojF1Ps5k0faOL2Puwv7TaRA5vrkV2kySaCKe9mt5wUF/DFY8G6CS
MbYUPF97U4HaeU7EGdDuBkVtFT5ivZQ9t7rCoWVnEURBEm6d5lPw4pLVgY2Uuaz5
saSfjRsWc0SJ1eotSBwjpQJT5oPbLwrqW5E5wUKebQxqgRihfj9oA1SfRTxKNXSV
UuUBn5jf77IiRYEND0mKmXJMU0JZX8mKY5iH/UeRaDvzyYKuKaIJz9dp9Xiio8jG
3HSrDLWn1vRlFavQ4rjxM80ma66qyw9z9fTnplqltuiCkGlRglj9jDnMlR+dElD/
brpiE9IVYkdPFWChGYzBAsiAOn0IDw0KQFQfDwPVPYp1RzoOvgY3/4auvc2aQWHr
7xZLsEn5+Gdvnl3HGxcWRM+IdthTeaWEx6JzQDE1eBxlhN2hLwtbrHXx09fh2aVR
ZkKS9PZkRx66pEuFop6H9UgbzGxJ+XXW85Hw+CMCK7jzt1oYW0jAfQqjd+rvKt0a
uYuOxu8HU/69UyiSPaCuQG37bLu3CIIDILSbderqlszS38cYmKf8wKnIMO8bov0H
MX6/pkjQJWlbhZk7knAC+kQWlB0ujZmOLtz3tl3PZYTZ4vu4gbW+Y6DdB84ZtyPQ
4ulXp8A3YKdm1kz6Wshm4WryUqmYcYhbpNKC3I3Sjqq+rO9iQujMarY9kl0kxKbV
ZDrHkY+Oc4ClsOj0vpSL0Le5abRRSPf/Ts7qwaiIpkaMtd7ctOlF3bC3uxgrTOTj
jValB1ggBItfNoDYT+Q6WWsjESa8ZjYmsToBqXHih7+vXkLhIXJ3tAXrX0DoUQzr
RJaVqCBLgsXhnNaYW6gt0yGZ7lFyiKtBkukblJ+AYwRFVmi+njoKo9r8o7QEINZF
0Ab//yck2BKTWFiIaEcIwIh+Dy5hI1ecNVQmAEXVM6jOHcgQCMXrLO62CCzy2yQt
CuVZMaYMt72meQKSngkHNqIEwBeCK1zbPEk33PODv3KY3PfRUdTY9g/cMwCphP66
/2PiodWVWvfH+CHjYe3PxfcIA3OqEa3h2ADi62C2JJoDmFNAu8coiO5Qqla2smoA
AXcwyUqC8/A6aZ5NiP+VIOmoXiXjGMIyWlaNcG3182hggM+GiX4RK31LMd/GqhJT
TNOofmz3Hw7LvnDDY0q44DM8j2APUlhX440vaQFRSjOegGa/ti5ATzQX4ilpDUx+
/Ugtnuxl/hfeKqllsZ2hodrt7oRzVPDWLDg+IEXphipBAw2ydGZbza8yGUZe+e1x
j7mhogXP+hAG0hnAJ83Dbclz5/trFZF5z3HQi4pzuzac3emGZxoG8BTmAIERfZqn
TtlyskP4tfW4659CnCwRtJoI1mkyxE6Put0vXS9dK/rfoWAmI9B9DzSjAztBSH9x
MEZHJTwbsOHxxxvJz1PZj+1sS5uDFFSfzVNgaeANecHr8y6ADBcke5qqIyYPqo3p
stY7eSA0hbkqXBzOQLKVI6R1fJ/hDEFSRzXydRXwPaF4e7dtIBjO0QbZ8GA4ppQR
FlEET41YE07WWIXH3IwxycOQHL6qHZJSOC/cb3hg1wH8v9f6wjko/E8gZ2ZSqjBX
HOdshhsqgVYq4G2wxVnJsZRPP7wo1/tgUKmJObrGEy3YHz7qMYBILg2ImB55A43j
/mdKGfRhPerq9jUoXwnElRQ5+/256X2mZ+K/TbNqTmmHUm3/TLcR6eTbNoPBWaiW
5I63poQJaMyNRD6pTTINvERifloE6gbBHFoCZlhQ+9+8JFW2lXjnswMUOQ5qBX4D
qirVvn0rqfKQBBWlUOdg9QzfI3tJ9cNp/9mA5zs7FLstXlW0yTA/azJgLwXXs8uA
5fFJs5Hg20ziCu9rVVel8dg9V4EA4a9T51i25jixCKZykOBUZQjPq0bwYLsI4+Rf
6KQRCa9FhTYwdTQR5EUToebI0lJBjPGIvDDkoimx/uZJb1Z5kKnHM7433VfjArC5
6QUQQkD2aALqVa2N6iRNFiUNp7sd0gCt9nAKYNRaFv7IPhIkZvjhwH84O0dH3IFn
WqecU0rw3F536KenePk//OkpEniUO1vuHLGZ2WkqEZ9wl4Qe1TLzaW80w37JTUqs
OHVrMESlWpv3xWTIyiKJb17yRcAOp7qtWBe1zSo8GQIWiUSNPRjgnIjz91nsLNwU
90Q4bDzfNJDqKvAkhPe5VcBLYzydjbsEvJQ2bBd6t2XfTzD4PAL13nO2KYAxxATI
SFrDEBXTX+9ZiGMSz5klxxX8UqDxewfaVdVbxZNsUyEw0jY1H5axLGPDB9amAIgn
UGxw+fS5ddnCkPZymOHUR+c5HhDI/UfCJ6P+S9rbY4FEmLENDD6vrI8qo8HhKzCO
d5bwA3ZfedxJjgqz2hpyBRmeCyyIy/wIDoUqTa8yAOfMydh7JsI/QEvehmMihlXt
tTRjIgOtVK7GB9cMQDsFprUFw3gz8fNUysux+wFItC//bChMfC9VCngfoqwaNdK9
H7A+Wb3S6ChJ/AbGO22oiaE9qQMa4zqyN8xprnozdrRVVbtM45bc5Rpfx46gqQwo
xE6c1KyrZtdqX+53+R3RED8I3mH7uPrTDkzeiggqLPZ5Lq1zroIM9Lt3AzCd8Tif
ZI+QKALs9zmtAjoacmvxm92K3ycEQsifQUsG/TGhEDeXMsIuvKkmoirNf9gH262i
TwCropqR744C73Ei5OK4dOwo/t+9zQsSShfwUX/k5nEwMs5PHi5Qev78e4JSTya0
SMXCEWc53cR57ckUnE2C4T6ltrkVVGtuMUSRVr//RvIz6HcFV/n/Y8Mvt5uoTGtu
rfwDeDahanpzyA0nAJEMNJNE5oiOIWvlBvKQH+5paZakd9GMuyERMZ6cecf2hljg
fO6Dcd1FKA0KQ7tLKpiDTTs4UIq4wNf7BXxxafnC/qTasNmCHnAqWaxhsQN3+rIx
lopzFNmxXYSnwAdFHUT9t3E5koqmMhuX0ldRxqW+twjM9cXjH6/YdXiGnl/DTT0e
ZNQj9KfXjhR6tkPan2uu0aHO0irQCyApLQE3IVp5rIFl/sOBXqKrMuTwk7JAUoRA
tE7R4mPqrmqtc39m9m68hJ+C8m7cHrPVoECn6zInFYF7juKaNdfqyvKnCJ9lIOHY
55LYu72jwEark+PJmnfyLDwPEGb/qFpPK+vXy1z+L5hr1bX6+iGKq5mB7fpVrovB
qHDN8NMVZg7hph+C+//PwFryn68aG01aGy+HNIf+yqVVDK43HT4G6jSdUNGK5lVe
X+Gl70uDGkgYT0c92dLymGpEceHuSTkKWhe3JFn+8IqtNBRTOlaoPlCkSvLe6bnM
XKpwakrdEbhjmR0JS8Nz2lhhtb2NjDEnsCdC87AX1JPKr6cceHpiKBagvlEAUSgw
X5wf14S9AB63ZnU44AWvCWpj4HdjVZFDzVT3eJYH6eSOH5/5eSMaDLpKei69J6n1
2To1jG1De6tPkeJY4wVCc2/0uZ+I0G0mnLfUGAI/3AE5ipRyjbk/razIr4wZ+4Cb
gMyVlLDQw+P54SulqlMkErDzDMgigQ/HF/biiA6oquqLpPi4B3NWQKiWfgq9YO9w
EEZ9RG+R97YhipV4BqBIFXKgIX7VGa7T/KfdL2w8KfZU6LiE2pE/rW9NtiGoXYnS
YiA6y5f7JgR+ccHZsMnEev3t+uhpBCtsf2gDpa1JtNEetS1VJnThtIk2OE01lXff
XqiLuKqQITf67f0dSZIKxyGCQpxzAHkAV7B0VaFpDcwFz4aNWPTnGxnqJJRMj6ax
jPvCXtl9fX+jja+mzCQA+YC2pyoRbkJQUcO7X/TDzJQBOAp/yTmb1kH2NiYvBoQW
/0P/ExY7w82Ffej6XWBrowiINKpht8h6zAEMtg0YX5QluEzX+1wVL3YxOUqulPKV
E1YhczE6uossQHi1Ib1DOlaFbKpp4+qWWdCEJY3vHGBuPrTQoD4xLIbRDp61TAVB
MRzoDr0QOE56z+Wc6APMkCw9ODHEcIQzmQeFsrov45NaiB9TY/QU1tcXqf0/Q6Gz
uQWuivWdEdMI6B9b3+foLjosOv/mHY3tNMC7mtWgbD46puFpn8CoO5ZlPrmAs3Uu
AunngTkktJvKOXTmZrPVSZJoAIp543p0Fa6Knka7NLh591UM95Z2C3QdA/TsqDHt
crG162Y2BXbZLHX6XH3Q33stBFHhcI7wCxelOTlLsa+3kxrOkqxDBiFO4pRaoGy1
I6/pYTFGzkkhNtFXdqYHOu9ZJ/WXmHMv/Qxv/iyuPi/6YmRzduuspdHtNO7XZiij
JwBjC/ygDtg0aKYh0JAx8epUyJEi3+0c0PmU81bwAJpHT00sUUNLCRrSUAvJQ/tN
T43P9oeYooGiVRYsVrIlBKwwHKfYzf7ng+qYd8sAX79lsH8TQaxd5gCJ+EfnMgyF
EfXvDU9lZjGDVlfV0ZFguSXhkl2KcznCAaWnNby9ZHNhSO3oyuWAMVhwZzHosZg8
elc3jp629xLO61Uski4z1Zo2CxLuRygybu2fL3/8i4HjECAv0Rrlf0RrxdxkBfq6
fKeteXHFLKFv6awVBqnehwRsW111+Zmx53HEdKWgxaIqdv2awin2Eujw3iwdfJkW
7+7u2Z4RD90UV1nw9K3Rbxq96dqZW5fn/15Pf5NUGDm8l6mbBanbeUhJ7KSitPQ5
cq43723hoL2t7GduQeJHJMCXwiG9HCOskaTGLgHRNrDEjzykMP1ADyzKZGx9kJpL
1VwMTno3FsihA4d6QwU5UuQEeK9NII0GhC9POKKy7o4afZddRiob7Hdxb/DGJGIn
LTEgHhALYC1mocPRucUBMUGFco1SLWCGkHieasdYSsZ+HRZPYuKc4ktxdyuWzE5I
TsCZ7BESBMgvxRYlxeX12SexVpawQTOl6rBkSIg9LdsEeCjlafMaZLyGzARS6ktH
fhJmOgVhoDopxEZVxGiJw7GUhbC5C94YX3LpAJOCzICrfMKd/jPfyph1unSwgni+
Vv7iLPtaS1vNq0G9nSuWBFInzqR+iwEsNkFgUzRLjjZXpvvfcB8rMbZrJACQMgTJ
tdT3tUKm11YbKWes4QQvbCyVTtzwqKM0opSfX1+JixJQHCSedHnieqOtAMcv5a+7
kW3QSkp3iE4WucJ2nCwkdnKWKTz+YkdPI7eIyWzjSrvd5vciVSusuyMop0smrTZj
OVusnHdD6CMvyWUYE9r+jLLsOi4p4nkwajMoVb7Ke0S7nxewk2tO91s0k4xeJsBy
lpMBPS9KFkF6RiBfxks+2WKogxF5kJZJ1c/BKFC+9ER/WpEweVYw1sg7nwjeOXWe
goCN30fmOu8+OOpkBBGW8dAnC2yAv6/GjwrpWMswB892R7lHkLcBnIIYw76hH/0F
sDGTlCM1V9pveTw9e+SVViCieM1pZrnWGu/5x4Mz5Pbdjr0z9rHUx2qm2WYaMQyL
QPCoIhifFUKZQv69PjldT76EZyJxnnwx6b8pLblCIS0CY/1aqCYSY992tu2MJWW2
mxf9uA1mfWSf8mGJAPuafMVvgiD0LDsFgPDZVrMvbtNTE7VfYxnx+Hi0grtfwgYV
lwPgkTgol9hAWrbDIr3semJUdJUwCUqRspnR0H4iwMixBBACKssOas17jETLTsm2
f6C+kg7nBDvif1k0gJXH/sTebGh1H8adtScQlVVdnEJZJ1JL0yf8qi9pUP79OoYY
LA3CvHz8Co76KHxOAw6vbv01SxdW40tN/nPtth0RXcxT5A1WIlJrnpAo4D/DVQQB
taWmg1sW5YdRvfDbUMC5XA1uFUTbF2q/gwrd7dE6v7fAwFwVJYmGcWTpoPquR+yF
HmVNaA0P8/fmVuQ04AMrDaxhwwnvh1k/vKnpPr4fQi2Ep1B6cDu9B8EgbZk/WuhV
uoMhVXmYBr/UD+cmKX1r58ejGgK74Y/m2MsnPVHjpVWOIMXkg/UevFxEaajhRSZp
Il8gqEgKx9SfkWt1JNxCSvnpw6gfWO9ZIoljWnPKkKgMSBSVjCAoJ7+i8KGF18AN
leRBl51Y2dZ0XKlNYvFyUo3+idaxcXBVPBICh4WQ3TvzHo+FSXn494mZQAG46+wo
20OJ6bOHU1uuBMae2cNulkHlMedewwDKgoAKiCJaYZiVfDpsEMhesfPph00oPr6q
rhzTNjUr1NiK9XaCmtGGUv0FM9dh1kLKFhr9bTefr4rZazrR4ZF3aU+TNeZ1JTkO
yhrfRCWYOWBKhU3tCnIOEknnWhH7LdDWfOMkvu0wklnI7jLVltTyvkmhwofkXpMx
Si3CRX+/7D69qB3gjR0RheYRD5stX8eU4jKfcsFjMZXeRws+eU/e+Ujdf6SoQ8Eq
7xeLxXiLBRRjvmDZFnQJKaM7oa1cIs26YMDg42EOhxHawggT2DtEpPVtdATWJN7q
/cUUHIbiHwNAL1IAXoDOo4ppl2ZJ3jWJbaxgTmZpRiAdGFVZ8C1VVMxHMMZOxrlN
K/y+p9xVTSvWXGzvvsyrvXIoA9Ce5vfOLAVMDDZ+rV8mmHmT2DmF32y+3rNLotle
6FVWKGJw8YVaDQFAI7zPhyc+7TqHuR8MfK31bsIIsHZc8vGi70WL9X/JHFWdD+Ah
g2n9amD6Gv9IvdHhPtdFbQcmPESQNHrZatE+mBUl5Q+/wExnsdxbo4xzO1t91Sp5
G62K4/kiI1AVAs5drAEMrW+/43CRhQTPxKyTR2YNPV96xtZHO7NMpSPJgvRX2gN6
UOQBCOwkmPXvNSy9ywCZT53iMz4hF0E1MJG6t49NHCsnkZdDPvwBlgs0NBuqBd3l
wMqal4CabxgSzSYW6CDEgigYAjWAgzx+t0HZ6MjbATndgZQxi5UeAR9YWfd7/Sxv
591AaxH7sydcSo1JN2nKGaDGogx1FUnjgQjxMhIEzCrPpGYDEHuWVQrzTjoWivtG
3sOeje56BwOGnsx8SzZODrSoREAzB75Y2Il3N67deLGHYHFzK9VGUh+hPHE98VVI
FA5hrdSpdY8FnOk0FXoWIVrtytc9G4EmteDENfebsOqYtg7coqoMZjTSotq/kgRg
/HjDNz1WRAwL76sIJY7FTCbhLt+z4TqsCyTJLPxoUDYrHlfj3KLhR4aKLCTkgDJ7
yhMrJ2eXyw+h2ncq/iI0+5dDcDsrtyUyyYc53aNwOKLG8t7DvyM3hG6BaDYctCfI
rUMDGx6AhsMGFvK2RHi3oKgPSqJMLO1yFBpakWfK9ja54Z6aIvh/H9LMBJsPJPd1
zSGPbrDK2oC4+icclq2QRir7dDeKEn62aXVSmrq+AgTDxxVbVxULRUv+22GSMjmd
7tcH1MZe+wpr6NlbRGDAbkV5XnfMrArMHEJk2DImctd0EkZ8OOTA6IGyeRve5N51
n0gKpQCqMqVxGD+ROf7RMnPIzQhwQYPhGEriA/ME4XccewKoQVWbRj6atM1Sbrlk
sUghoMPRJD/1Sfxha6ra/kLF8u/2dudoO9EhIQ4oo8wU6gq7ghOmA8zczYB3aE1F
cQ2XQeoRlLcv8w0pRO/vVSKMgkO8aBvzv/mRrv1f6JV6ScFEKoLdAJga0S9RmADU
YHyIVxRu4v04k61mdNp5PnyDm/y3TOYA4psB7nElNVCndEoYWR4/fOq6r4GmIghE
BgaYeLNLeMgJFBQAgAuu0XRA4VYZlM6PoXMbA1AIST3eFhq/jGyCXQegxPp3s36k
ohHW+UJPkE0gKfbJzC8PxmUJ1PEa8KsMhYlWp/Ra1Zq3aZowJyvu+d4DeuKqL0h3
SEJYO926lFSUKUzA+Tb7WyEySfNtkBiW1brPRHFpmS+XsaxDkzOCkpHAy/NZ0HrS
CrpV3xMYFAdHh5ImLcWrZal9Hf9A/D1/p23oX46OxFlZeELMV49Kyww2rg9L0jSx
vfFODfvjIR2bbIsJvWvdQSs7PVrbWD51S6qFSCP/2WBGqF75uEc+YLp+NlpMXC7k
+t/vVJiUxJeb58T2l02JdmV/OwfPxe2pDzlllEEb9s14gHi1BabUdx3Rj2JM1jwL
/ccAWZPyJ29lpKHQ2kZLC7TE1mqAvNpo21EomlG5o5Rtao4EN9bzjyuy+1mIZywV
wqhaS2Z0qpbuyCo1hH+9tfNSyVHdycuCqXeAMd6dXM21YhKtpHG2ccxoX/5rw1UR
x4UU4NC7MvjO+nR6v3vovnt8kNFs0/3xU/NYIySWZY0sjxSQzKzrON38mbq9wE6T
OS9pnqZvpggUc9G/wYb47jT6Z43rzmCebExygkJ76Q+IRDBMMj2OxgXuDzZp8jPg
RhLrqSc4QE4/+Qlf56HeJXq5t2wi6a0ybyzoKbmiCPSFayZ2mUCeFHKuiJdzX9s4
KkJ9JTRHBKmihAJ5GP0mCDW8vbf5tQWYzn3K4wC/4LpI1iU5p4h5vbaHyFMVPogd
adEWuSxbRLiaq1BsllMUaHU/dbFxrp4Gq7B7c4GInqgAWs+Bvu8lnHMYgh0npzoo
SnaOpXiTKmPkoDGEEofqvkehdPbUAWHhfwhSzEaejz7ykoo7/kZwu3VHD5UvB+Zz
ABZA4KtZdGjGseuJivKVazoOziI6UhQovJQXbjsauvgt6kmbcPmpEFRVwBeOk6a0
Ho7lRm9VggwIYyjVhtVHPgFTP3zw8LhkmqYJGdCwbN0QAiMdb3c6vnQaxnkWHlEW
jA/zE0XEHQ921Qcb/XN/LWOcKIzYtdb/KxPcXH/gzBifGiAKE1nNznlvtVq5rqw+
Ow1tYvKkYzCeRAVPqxt85YB9EED3yiIB9GVBTJnden32cTw16S2sUjeqPCMlBont
d4u7Fdyj2fHQ+bVO6UCxJoS3b0RWyTnbhvqvJpyQfsuZav9cn3MvprD37xpuoupi
ZiizOyPiNUlXnoENDtUEKcu1OnhdZIlTynU+qvLsfKNEze2nmkSjsgGQ6bf3Cw7b
/1Np4RRQULtY55JfkXC7vrV5YIPQucTodgwQON6h6fA6v299lgyWgrMtqBe5mcp0
dYuRMQPAfCsy1gjDTMLlhPWuSX9I5CGhPizlvC35hcnExsKIPos46A8lMBSlY8j/
jBQoY2mbPfncNvQSnGHloddj41My6cnTKnEXuSzocfPRiR3pvVndB9q+cE0LmtzJ
4uE+j/xZ2Jg4956Q5GnLHc6BSU39wRx0N74qr8lygRSMacOkTPCJC5O2iY61TkKf
9KgNZNW2WgevEUuDSLPQ9K1G6troy3FBlPT5Xf2pAzmPT2edevUWtQdULIXG/BPK
u4xTbueUrKOXSea0ioxqZ81E6RsRXDARDn2GP1AWLWZUoRpbI3ofkjN4XFf2ytkF
0ZlVKibk6m3R6ZgtjE6quo+WrmzrFKXmd/EVrcxQNr+/MUUUamcxYMbeXs7jY8lF
xUBucaDTsKAxGycz3luK01OiLEf8Qb7pCCeB9V0V5YRpAZVNc95zDJ/fHqhZipJe
tT2Xa6VE0AJaFEDK6DdvrcWPsq3GcR0Jztqc/0wPNxy7YG4dLsSxwWd1hCVvv/sM
qNHLiBYeJpNCma/RawHlqngRPDWdeI1xh8mf3hAf3i4KwE2wWH988/C41lHu4E/O
yxTcz+KEFYQYe+PkCHaijSXydOxiuOLO23W2eUgyhZGgH4qH+1SQ8u0eD3G3ydFr
Yzwxc85icPuf1TdVl9s7dUQiXfaAeCojxA5Z6T3QYMx4S2SA9lEovfzKdD3oitXR
WSvM00q8xkrHiygm0U4+4eI2RdFMy7y12P6en5mhj+H2p2UmSbVneT+QCpILj5VO
PQxGKF1JgcWODF/zBRoGtsQIh/a1kvSur+6qt3gzeSHwn+X4LhZzIAR+mt7wYB2b
nGOpCFrnSgKX8Z9zNwC4R9zvd1zZm0FrkSLTk02hQr+U5aQ1pc2VBNu0PHtRGBVS
+FSGDPqzsoxrNwSokUktOpsv4XOQAn06cYrFPrXAViMvIffhDVE5a3Th3HUvoWd0
JC9BeEujw4gJp3cyMVrWvxoB55G97kV1nbBxQlCfiN7rBVilM+PiAXuAGXdoN0Kg
l4cIoYQ4KYyjvsKJqHSKcJftEbKhBUGQgAHHy7dFt57YnzjrQyYY9jxFOoytIrX2
JaRqa5A9iGrNwSMlm5Ug6tiXGD56qlyBjorR2idVoewoZdjV6UlYRy0Xo+hfNTzT
oL23nlJbwlzD+1qWmo/QkSBDfV11cXSYb6S7H97MW3oWW3nMAqk0h5v4/7le0hmR
GOpWqLPlUdoTlJ3cz6FGbJBV+PG+i1QZuga+tvS3sDTCdVF9VNRhXBUGNfGr5dTD
mAVQG9rbwkwD3ssCSjr2zIhB2X1vW+gJMrNmXzmy66XGI0PedBqWiwAD95qcDfGP
91tX5ySQr+ddogojWQDIf1BQ5JUsv14ZSXrT/n4IqOqAA30ELtxpoJ046KNJiE/0
lWuAo/uk2lcbh252mRF3W2Lu4dh7cQM90bCtMT4ffIP4i0fQ5ivgZkMXWNxc83QY
7gJodsMtUD30X1ocFDoLyozDyrBgivms+UbX6SGSEGvqIwWfO/n6i0iGFhOAbxKT
1bJrm0C6FZnmpsYok5bDavXu6zXUjpot82zCc+fSw+kMsmtnBlrTedjGiAOTAias
q2mtLKSPTItODOj9QHAv1cZUlTenCL5ltNMTpPz9+cqW/lFKTXHI4tRp1pco/U2+
jmMOpyhrIhFu/fDe+OYKZEea07GxErm1fz+NO1siZDyiIwOxXXOH/aFjylExCuA/
gCQfzX3Svm6aMiXy6mu1KOy515XkAnRYLRMzIS9Y0M+ePAQnDKYJYQztJdR0F3yF
dFAPUJk3ioH9g4HC1qT8xTt92FIw7WrVYYPc4Oi3PvohQkCcuKImnpeDFc13QwWk
pCtORia11E69RjJyJuvq+t4FLRe/TlFczPeqVAZ7Tzsk+dLD6DcDCcw80fPYUe59
Qvc+vaqzN5iG+WmoBIiRnOJiRGGUv/jzpWrkN0uuNxKlwRqierp2svgnC+17cVqM
6uyzLVGkIKgX2Tvz5F9nypRYiIJtOj/CkQitIefNrZakTUXDypfH8dNcT5XxtBpG
dqnSzRo5iizxYqd/WSCml4bEk+Gx5erhcUQKPNSHE97MOunD80Lx8D/PKTcxWyIs
6U2Me+nYQcKZe/edEyTwvYvhj/YCjQfVa+W1zqtJqa0y4iNmDA32KaP7hKRuNy+c
7nM3g5R1KmJ/AoyZA9iXDZUv2rscFw6qq1AJvmulLELB4tCUNXqFg10oixB6i14F
hPSxv0AIwL4D6/6F4FD+TgQcrYdgnzX7gJm9KAO4zE7Za5vjhwDzhcDqPxB2LPrr
xSteD7pUDTyBKWvgrMCh9s41H+17OYKATkpps3DNa+Q+a0yjLBWhQoYkgRZNy/JS
HrRE89v8/aBheQeOj+hfbinV9WSOs+yVgjyDe8OO1EoQjmkEsKg3+vvzN6XpG8y7
1QBGrI6rpAsoDbNtlxCOBEW7gaPhpBsvtQJmZ6amNkaXhSBeHXQbZjKCSEoLxo2x
92d44OSeGGIveo4dp1EQBvDWGx5VHVYucmuGYkfdy5UfuLA/ADIva5QGL6Y/s2j2
gCiy3WqFLovbShiiVeFA96JUwXA8Ks3E8Qmv2YUcu1j837+BYxV6Zi8LSmNdwrPK
qpsL6b3DQzDsfiLzehc/JejtxjmpU0PQjLZtACMZUd/P2biTkw1R5H9fiTYZ5U03
bgngoKoSX9WGxKitsNJ7Dxb0KAxWBeRkXv52+C1PW/lYn0CunvIlA6rrMy1AZ5AH
F5da3ViSfazmscsbiIKZ+G2kPvdErMXTySwhwpSLKSDCsxgI8Doh77yRv+E6lVHk
v6+XE4a4nwHZYSyw2vaVKzzzXzD2Bg1gZaZ6Csbj/i791TqRa0vboXaeAJ7DdeJh
p6DbDDSfTeAd53dE3D92xauzLA3ph+ckgG2AIpK3uLIdw4ZqWIWE8MpV2p9i8oG9
NsQEH5IvWAbfFScByKWUCZeC9wH5J7idTitZ5xKioVrcJzZRYHHWGPrz8ps7W/Yl
qnqiMMvCYn0bZBUfVcquQDVhcLhIGPfBuPxEl5MKnMdgQbwX9QZsDJOODPSKmXYx
3BZyJm6YaeYI+Swbj77V5FP6GugeB6S++a0OMOzZ6pJNNkylZ6VcfF51pw3J/Dqa
OLMrrp/sJmAmZc45/dgBpxrxtoIWoRzGEUdDRDWU9G8Ham1HNzkLZuhw6DYff2aJ
RzZf3YGKLiRvElfREkYZYEmT5XeN0Kz+QIZsaoIhYgxodhuxRM2N9224+t4xxLDs
D8XOJnxW33X8jp7WWXZxyfTWFgjDYYIdZcBbDj5qcB3AsMDiFi1ZxvsAXkWX8bVx
XZOe/H7vBPevA5gR9LqjZB5EDgEg7Qa2oMkDcdqd7sZi4+QV3EMn2XzeyOAjtGTJ
ZINcqJzHPyd7qfBR9kxTAGeAGkUW94gKK7sjFJlNjGLJ3FnFccWGD/VAxmK3NrcQ
zmt2sErfkLm0OGuDCqzVvAbYhxATeKKUXgYqc02LUpPfxWzC58KKT7gNixChdDna
vGu2np0nH/XGbsGr4wtT7Q94wGXa6grIRW0s2Btj2AhlsikN16RHERCHI+lJG/Qi
+idcElopYPg1WsNQwgt6xRqYdYfal6csLyHlyrTErHq0srt3QO8SgZHdwoHW7W22
W7cmYllY4oRRQhQincm6o53yAX4oAaffHmfmGvPVih1NZF/F3ZYEQhrBuZBSWdQ5
3LBXYU4FSHWBkGaFJoEk9JQ5rYxWAKWZVwC6Wv0L8XdD1SsSHFxQgJoUc+9R6FX0
7zySJKvcW1ue/qjFoXqop0cQxtUHWEnfadoKoLTnS4BVf7kvESiMdikW+lSO9bBj
ik/RJ904eLDSiiPelnJLJe3BV+3mRf3mHWZINVrhvrdtKFq/jgNdPd9G9tmU1Wrt
inoe+eaOS7xZz4AMvdv0hTwR24U4e/4Y6VB+n2IOU8tGqIYuX59QsC1KQ9FBcGxX
BtJhykEhKFWSlH2ZG5UFSMxMroXrBRYymyvp6DDfQ2dOCxsU1+5Va2+WXwlkabg9
ghrIQFTTX2vCoKShEhNR6ObqH/hAfaIZ+EhpurtBxDYntZ6vjfbzHUIkWhEA312j
h9yyumU8hM3NjKP2R2wqaPtsmOhGqt7HOnEEmSRNYH0opcBRffVfisZMqTQLeR2j
1wF2nkBG4/DzF1LFR9BCb7oSULaNLFGWmqG/HGYGhs3QJbZVA/AEc1GElNYjTZ7M
r8yL2Zz8xczt6PtwopT1gp6aayZFJTnwLf9RiwvcHLJgzBD7AIi/fFcyocuOBT5k
KcHUzUdkWLRBxLIAdY1yTMlBuMR0LPwEryakC27jVoVzyMjDuHN3gIW6zpG+UPGF
TkWxyO5UcSWdeSoIVk+Vqp6ddTCR2iWhURpXLy5ME9S7HQxKi21Qt0L7GwOtEutk
y3Kbas6wXR0VbEbpjsaGTarwUTHm69FxoRk9YUw9wwML2l1Kt8xVavu2I91gKWIa
X3CrEk/vW4yIMNg/Igv0BFT2UQfwLBWr1vtZYlk+eQRTK0NxWTrf1mcgs7NwrBch
NO+F2FeXdg20GsPxda/OwrljxEl+S+a9VKfn6DIMoviunZccXjJ/9D8iRphXN3qZ
U4XGW3tYunTRbjzH05xuzNltUyPBE+pCf1dMlNS9wOFtFH3FkUf8kofU+gpgQ4Tr
kxTCEkz3dXZwCz/1m/mJDbYrENHtYM5ALb10JS1dQcIPTstjHHrPIovW/1mmhSYN
q8btCOowopj8iUBkdc0WtlD1jDs5h62IseafjkCpd3QyjiVt4bGkyR9HDre8N4OK
CI6XAfi0kmgDk3jAc/I3C+rir+7vwi56ELBO4tHCzIpdV5AE2CsXKH06FqygEPXG
kMi0Yk0wfFIlu2tszrdSpYSWIjf0+fqP5IxOK2KPiihyDCeovX4tiuyu1aWg34c2
JCkl9kJRaAkzPSIM0qYJ+SP9CjeX5qUGqwb1QMTFX4JAhP0I2i9utdjUoZwfvE9f
zcmV/YHG8gUye6ARjcLgtSoycOG5xdxA6wb05ytVLnk7z57rxVfGUmJdruOdh/0L
Xk1S7H1ro9YJM/0mSiYIKenuXIM15Zs/hia6X3IMEqZEfDpraUl8YgSOn2sEMrxr
udEmfOhV8T8XdpHQx5pq0alxtw9nba7Q07qxsyLyMfP6CVktUnAGM17gsJtVd6bi
ax+dGYprlmn7cdPJgv4cNailQ284Kcgs9TIxy1JR6DiowlAhnaaiJb93tS8o2OCm
0mxr4dS5w9ufyRHbLD65OeK2ce94YmPuv6Pvs99qvQPP91x6wQmPX/4Rxkh3XTex
fQ7f0QJWuLOI0fGyIOIbhx8dse9K8suDKOBUz+GDoo5JQawKJlUZNRVumK4JfqBF
sS07KfDzc5zxQC50D1Za4ludwrN+rZs7NpI5XQclWTQGL0L8vT3GzpU5MZdbKuLk
TViI0MUyPMFPP8PSqNI3dgNEjLmg30GiNWLSAJhXRc2IJNSlPhS5KcZfjSD/z/nu
UOmd7SeCnhV0KVGVJ9bQIcFQI3V3K/jUaI29tmeVaajMscnKXw9Bq5g0swYq4/rL
6xeBt50aYoTgMfAjleVXOfDd8AfaJ8Fu8sFtXxo/XkY0Nf/RstPHd4LaeV/8chQF
2ONjwGrJTjMWUn0DzuHEUl54TtVacpIsjBJntamsMDS9P7f53QInQHzxHyw6wE9H
gtVxQASkp2MgjyCPa+66xsqrNubgCaLbXBQ2y0LI+wAA0VExNe15vrUsSf6WUa7g
v9M+grXLrZ6xfCDqLoQm/HqRIyINro55bfH8Aj5wMXHe+goY1NbxLwBmOcdJSdgY
E+CRjxeqDibGKaUso6vs2V2e5Zc3rfYm4skrG2kbTxE+clf8qiA1Ni1aBeWX2Qu8
rIEYXs5BCfjFEwHoFtO4uL4ZrUNf+XohFuxVhDwf9/QcKn4HtCaT1zOiz69UWDID
kbUAIJyzofAMlpaq83EP1R/vLLQdx1O0vSWAwV6Yi9N2vskF4xBAwzPqlOpI5WQy
9PvtfD6FJMHWAK+XUzZyElnfxOuabaoBBGPO4zBQdKyon0HMVubYRJzXC/IL60qO
LLk4A5KPi7qfCGDm4qh4OTK925pQVK8yAhkymDR9d/WHJk64vtvhsH/Rb6KXzwHB
0zUt+ZLFPMV7ccJIRWrTXxO/PCflS8FSpLFkFFGsIXrPp/PqGP1p/hmW0FI92B2a
JCqrdTHXBDtr8ZNKI4rSxHhOm9k39L4zJrfktriGYDyuDvwd2Uyw/Ifd3GmVZBk2
4m0GdaWC72kI1rDl2qraCd/YXmutwFRYkcF6/kxVQ38zDXzLsf+wPI6zVTSbJnD3
TBDSCSxqI+WgDSEH+Ll/SrabY9PmmnJgZJy1NVHEVbxaif4mNIpkdAs/A/f3InZt
CWOM5GmQSVbNKej60q9nzYznvGcsw8fm+R/jeS0TokFTha2YAaUUgVEiBHlg1qJr
iHwo5iRhjU/KTsDLcMfmipFsmTReCIANKatICcLlZRdti+26qqk5jHMrz77R3LY6
5+aJ8zNo14d7joNcYhX7dcWbKZ6F+zYQOFnJPeow6JP8ehbPFrnjsgTq++y9+YBQ
agVJqDawkknxL2LqSwHYfToN7xk1As6Mhej5gx2KnvGEBnGR+EX5Oj5CQKd7K0AR
RiXmnptVbD8f7f+rffUqdadnax7VdTAQSXZ5EnNH99QlAwTFFLRlzfG6HQBcs4YT
qhamdVtVlrNQQE6yeAUTzEYDwTbeoxtxNQ4CjqqKxTg6P6h8RWj2ktNnuzGmSbyD
It931ihNDqFki4+FF/410ifFrqQAptWMVYOpkvFEvT3gmDxapT3eaQ2kW6FcgMJe
5u5ZEs3YpyBn6kLVWawXP7Vxl3B1wKBKfbSihi3qbfiKecBA6AbUgUHMtPiGa82E
PrxHVH/dIALG+vsghKKejFelOcjQ8uSUOg0M+OvkANM7pxM5+Zpz9xR8LDPeTCvb
EdC6x3PD3Cn1eDns59yzIGMj6kwWCDu8tn/QuCb6ojB3l9wT1mrHU6wBm44VufO9
hEWXLzC682LyIxpk3onuLHeHq5wwAPubwI4/PNwWyldWvdOggEKTpHkXdves3Rfs
6qkVGRW65KNVW6g6je2njoQqC92qiSTmJr7IQP5BOCE5rp+ahbuEECp1gXF69was
e/IV8uZcZcT/xRkcmpilc//U083RglCE8dKUyxblDT2IXQ/REFf1C9patbTyUCfI
ESvBCxjs3bdW+kBCtkJmJyC9zb4Lg9dutewTKGU8NlMD/tNRxN04YZ150BTCkgKC
jYF7Ojovr/oMbEmR+o+Dvt2oVBxZP1rqrGIGYzbg4uq+fLjlmIRRjUIEBRnkJvGz
fPxhPrWiEdKTca9UIYr9anfMhF0u/vYcsAdqyUrFDV77d0w48z33Ma4Ozwmil6f3
7CdS8MeS+S72uMQEKTBlNrnH5AcUNpP2E6niMlsf4bvSiH/VmKJQv1lHHnoGyFCd
uiUQQdIK1XeNPhTm8Zk7eXCZrx26vtMwiM7Zh/YmqJxfe+t25Vj6ouaBhC9PfJ+4
G09xejVRYo5J8HpVVevC8gXT4aj1dgkgF7/eXJLTZyC/+YLdQDiZrct25jKPhgr5
wYCcNaa21vWviz/rA1BccISv76OxA3VO4avocuDZIyQo16S7DYyGscmJmsOIcNtC
4bEzD+VQsXS9zbFB2R6daaeiKNk6tEiJc7qiAH6y7KOoPKupVT2FmAbqNzD2mlbD
jje60Mzalg9iozOPxahy8Ea6UqottWDHbhL+W2I/js2/tcYebSXa3sUTVHEXW1XK
0VtRLV8hViBYQLlO00+U3qcYXzrAP0gLVMU2MmxfFYdf54qF+WaNxepn7D/3H8iI
kEXWFPuEfSF9k7cy8yiedN4VtaG4rHBepbiqgj8DAm5Qjjtk/9iEKHsACQbLTdt0
cc7kd6Eo+a56fvDcwJ4LH6pM2Tck0qwUiaAsEs7vxxPuT8viCkNeFJvDtkdgnp5M
N3Arj6kvum8/AMd+jPD8rdUOIHxZCMowZLH4u3+mXbrlbFRzYSFDwOvv2X1ZoVOJ
io3ekM/7JMiqjXBfVBJ2JKKSexHgMSi2Ga2JiQsGduWLCeNMiXNZR3DHoQHYptZJ
VChx2thGfyUvOILipBZGT+1vxCTNU9f0WJan5U/E03bB51WMF7qfOcp2SzDvCIlv
iO7489CmKneThZtEkVcK6MNgEJeMVyLnZ159cVrrz8ngAQSN/VM7LVk04bDZM3Yr
fRBXwjEJe5ed/++F3+2Khwzg7CInp81ewL+24QIpWYhh7WdoWA+Xc7hSdi8MFKjs
7JrD/0NkAhSaaYRWx4F4QrxoXXJ+M7auXKB36QBVVMBHYHT/XjylwYsSWE1jO4BB
kBZ1WRMyAylah0zsFL6eR5zQFF1BJpwom/1JSIW+Za1FRxLNG8/Nd4jF9/vUP5nY
2ZRinIL4aqyZvDifqOV+Z1vcAJtcxjnNVLi6W1qRNc7c9lUf0NElWz3VPZEmKbVD
rM8c+8f+xvZwDTgQ9PsFW+lE50YI82BHj4Qx3qI2gfDEOMItassLTp4fpJerVGlw
6Qjf4WeBSP1LlX6Ibqyljkzu+qk8j7RaqJF2qTxQ8kxAHz1pdvuMyEXnuN+rNdhQ
tS82tCQRUW6AQF9Cc+XVIsRGnz4BMjRv/LZc9xLUexrY1EzOnS7+HJhcdLCv0+Ed
CzzXnag08P7ZzBy0XzIY8UDhhsJN7+0GbjOkHi0W+xHHw9pRRUsQ88SR39muL723
WIsrh+FTM3P99EH1jdS67HwNVyRyZ/HY577X9mu+RzUuTXCy09LQ+bhHiuwuOucR
quhJFalByJT80Ay8gpWtkq8MK/9z/r6vrGQO7fs0FkBXuWMlO5Bgi5GdlgKtT//Y
Vly9l0XuwxbKWd3tMNcZ6twFdu7md0p412dzWy+A5Lckbq/sYBg8CFs2WbyaDmja
tMA6KmIJXXaRZiJsqKEsAa9fpBE4UqUo5rsuE5X4Z1wvTd483DM+W64owCY3Z4y6
bMBIx5zpWKFwkWDU+cRZ4nAW1q0wQ5Vr2BXMCxanBwSbRw2VE0cnOy8F84JNod/S
pG83vbEckg53YSa4EOIg3gFjkQ91vK71/aLDOj9vraYxpq+YE6PpmQ565soSmJVe
8JGabujN9PJDuy2m6x2B8KsouMu6BWaDmiGWe1ed1n/Uh6PsnYwuIL5u5v3M2ePb
xC+dWtnk6ekzn22gktBPZlZ7H6UBwDs+F2dRUf73DfiF10UkRBcYEcPLkn8/PKXH
NzKdY4EgMY7+1/qxjS7rpr8fIjhe6Xv1G4G5zcGVSibqMNh8OOlwDOhkfnZzYg1T
Wp+UMqs8ZLtqIw5beAg+PFYZFYNsrQFv/i21OwN8wmoezOIM4+u0ZWM3myjT7aJS
KCxcvEBFGJAOcVlr/V6+kOwAOMxdTvNIGHD7yAgnKT/C/uiTwIfxxaYGbl/WFn9f
F1LYgxorD1RnlB0VrQwwqZFDmWayKcvmfSKWzRa8SL9IqswjtYE6piGbF5TxDzEd
/79sArIJeIGTjDbHbBBaxD+UQjQ8hPPsrtQW2MzVX3QNGQPad+knTRIVwrZJ0Wxf
Ba6UTHNw4fZmJmhWXZLVxzxdZRsFI4LNwksRE9jLrnFKjuUzMoNdgCb1PI3Cc1n8
ZVuT8Dncjq6bbNrmeD3l+tUmFLYqVmxD+jDEEcC4kIsmvmsMGRsE1+VGl06W7haa
R3FsZxirawoic3b2RXJYsSfj9+eBMm1uAXlBifhnGLzKmnErS3gB/J1CAK93kz2L
7bvQnRvvRgoWcomlbEWJYZ85qPysGMHIB8+E2w7KWpQXomy3oUx3q7ynj5SFKRSb
ApjVL9RvI/SiqVZqTCPx/pwFTMaeyTMkfzsicmgSzye0Ehq2Po8Vdf+m1pmYUiTS
t3ZXudnF/6qz9R+kARSkbGWE05KjnM7zF9W0JCy42FaxNHl4SwvOyhoqyrXECxAl
t8MXqw5Br2X2KHRy0JIeFOjzK2k2nIOoKfbwR1rt0FQWOyB2K5Md5u6HAT8qU0Ow
1BwTneddhAQHwJmqnyYGqN786QgZwH8L62sYStmMgXZ9qHQnzn+1LfV3fZCaZo4I
FkYZpBntUiR+RRJIchfNe5FNcllMQC8Vg0YqU4Nhj778A3xDvoia7NMwJNdmRBIO
NNrp60QqUlWJplvuBE6e8Qbs3RZmq8h+dqZHRzflP4i81viJsChTAGavkTf1hAXK
1xgQMiHDjLT/zc32VsAHYzbVFBxCeKA1aEedZnV8CPo2ql0NtV798rjI89DJNKG+
ZZH5UXS+Xj9r3DE4fWQDJEpzhB5kaGBQvx60Az/JTfbMiImqT861nBssYSMewWex
dDyZu1zHyHDs5kCTL3+MN9/YPGAZ8w8bfOynmPRJ3/FO1Mq/ORkSy0tGBG2EjHUN
S5H2jeg+8fPaC26deYBTra/Jsv3KdabKnZECdouXfW3EKYBMlP8w+mkgNVQk4jh+
Q4Y/32nwHJYjyWEE7t05BvqrnZSSekl29RAyvGfmEoQOJFN2vbiYux/fY8Iryera
2N5Qwv8gdVToWTJM35TjY+9RHLeamAnpwUKS2dDMZxGt8YlNQs6HwoRSTxYDMZ+4
nFs26vGvk8bhQfnuIwG43KPNmcawaq0rUNmbQpwwMYY5Ijn8/9q0OnshaQZjvRnL
giJYvcqKIsjr2I/ZrQSMrpbe7w0kx+HFoHCnxXGH3u8pRn6sf0eZFaxuvBrdfZCI
1fRJ0MLFIPuN2LwoSrrwrK34/QhQ2nTTp9awpTCI0VMwfDlwaKp+HhauoShXDeBm
cAtRbitcV8vRuNx/53Hpdqq/QChFmzPEhfl3kh19F79Yeg0eeN/Pmg/gaVs6UFGR
CHSKo3GbUxNRzWofDbgGeB2hjGeDja240LBDnjgSFTIbaozypR5h9BRg6USsWUir
pLfEKQW3cJrebk0mduJMOt3OTdPJOKICxWEB/uynZccH3P++a0U0/9vp6O3Ln9Nv
UZ0LFCJ4wl+fU7vzmpElrhmca7gXJwy9Z3nqXr5M1bBbN2mIydA5BXws7y5fkDbP
2MHHviSILQudblV5fKuKbgxTwMXdwQfD1Mjq80gVromYUNfogm7e5K+z8Mbr1c4/
MUUqHa2ISjdahfdLsBEeOIHAOP3JLAmTo5i+cQZTPKj6WjDJrrkASpr0RJ8aKmNd
xmldA3X3SHQV0S8r/Dd5OeWAFfAJ2RhM4v4CPmtRvX5kBr99o32EW6Cy9FdVc1aB
w33A+hA4zOhXcDydddp2jbvc4tvZjTkNvsYNTxvfITsD9NuI8jx/AAntupsKdftq
iq426tM/BeNKTY7WXrlcBPt1qx43Y4Wah4vj3B6ah6qIFTqiEsmsatEs9oXKzDJd
dLG3trA5vOneSe2GWyAXF2FuYPmBDtgniDiutVoKto50MLfEa0PRzcjw7fxJbMXm
9cjXFA8/h5/Jxn8FAQCEK7JdhjRwvXo9r8IrSac1T4tfPr9zLAJiotMJZ/MfFEeB
E5JYpstlS/jds3tGsie+UKgAxYoxqyPpPAoBGCCIar7tirf+rRHwQJdrtOY8kZSn
tpvVdzW+dXjmiw4pjOdL4+gu6zDXvHdSlf3vtrVqt7G26ROpPkdEHJgUDh+9T+3L
reHI+7AJw+PM3uD2aeDqCLHeZEkK0nWnliBqVblndTDop0/NDfRmgDsti+CKrEcK
aQ0qsWtC80SNsuxK8tdWjmG1gm+otgq6Sx/cLRd3Sl7uP3IDNen2hf95vIbCnqIu
ccx8guajXSMCW+5BEuLAoCCjTBIUnJyDICJZV8uFCYu/EoXmVS41R/l6EZm4HH2V
Tt0F+hNXs40ZUIlfA6shV7KnPno8Xjj3AnG6CxhV0aqGsmOVehyLcns6RYqmmriw
sm8vPIxH4RajIYQKmwXSiDcSKMq7cJ8gIMHScrtoIiHpk6B15uylPQWTHyQH0v7x
2J95JSR+XKs3rKk3/DdPBwTA/yfphVCKRGKL2U8xGbm8SK+kloiqcXTb/+Fj2uKz
I0CX7+7n2ID5V031M75I/V1e5RQEtDj6VVp64ek0GeZMwNVz34MeqPaVyCr2nHrt
aGnfwpeNu9Q47POmieSjpveLXoXoYl5vrMA+62GmEl3dhhGfd34lknw33+A1EQlz
r+T0qQ1eCb6XIUjqnS7PCEAdauLHW+nSX0ivkj+VoCf/7vnwhOFI7aWqBuVmuqxT
Xh7pOVmyoM7UfiJ7KgUgSgu0LjuaEfxy5dUwZM6q4SknL5Q83NEh9+rHHiIQKgEO
AOvyxhY97y3AgYRWc7OgtuYMi1OgAB3VesN1yihiJWWVsslINWYZ0HsYLRSTa0iK
CE04Iw7JUK9QFtvCuRMXok26gJiYbTma3AehCWcD6dA8M8mKb4XnH1Bfm9WOhsM0
VYkKLq3jZHQJsHCc+wMElGjXpI5ww1xS8ciFmHw63YYBqE4uBvtIs5Gy0NXZiAbZ
2lmZcuJ4vmtq+XcCKV4zpqIxrJh5D1JP139Fyj6PYtGFRoSUAXVy6QSYtv6T3KdG
lyf25HR5EjgEIgseRCu8TxfafZjXVwGjcOD+Xsv4lCTaVDCZuuzgIkS7dns5/qBq
9x2WSeSiDE8KyquNmzFq8/XdipdAvn80JParbBqffVoQyD92p+uDnHzc6QUYYqQ4
tr+kZ4KNgKzETkmE9TFVhDz0Y+PrCG9ihgzXbcqn3d3sSZ2v3bgSRwGPHW/ZzXSV
htzDQnIMT9HEyVioQqnSidBRjlUaWDW8aYwv5WPr1SoPDlIrE7OV6Dndo8uw95A0
+XJ709AGurqK5ya6d/dB5m0XY8255uccFiF9aWMYUxHbdT7MJ+gDzomt3KBZ1uRQ
wIUW0IrSOCt3MwkKQ9Ww+JcW/Rw/P/6i1nM6hTuDcgMX9dpileWi3vhBErTX2Ody
arPRwsDF8EOf/F5rSOXOu5R64RdPBOcPhSzBPsWEeHV7SJ8YpkKW0eSyeXswwb8k
0FeTIqIzzNiz1Yzxc/hRBgatmbjUxgcGLd3XKKLIlC/Lt/mDlC0920t6aza9tHfs
hepWmhqUomX759srX3wQA1H5oOax8mmtSxutOc0XhgUmgeN9LfB6gVRW6fkUYc8z
Mjvv/w25bGu7ZTmsGnPmj5s2BSNQJFfSNM/uhM3T0yJmqWYUpOcKjX3SP6Nwp7ki
DUF++Hd1LGhKo6WXQ4X+fIsqnC5afU2xqZ9JhBx8CfW2bl90Nq7BSGbWWpI2Ngq7
3MZ33nhi9ObUXWE6NG4aOIBcwc042pp6BoBgi8Q7Ks90ZA6gN+3umQu3bNBBWnl8
Ipf7oItz8hz6HUuzecLvCd2BkYSd8u1kCLXsA5QYdqXI1gdlMyk2DDoQ1c7QP5AC
8wYyRGJFZ8iE8hxb86uwc1RnvAgd8M4jlSIOVhse+cRgil8Zda19lRl9U2IC3TxY
zDj07aom1sRg6DHHIgOh9vYhNFCKFCiMNvx21G+qgsiTpFFp1ptUczXwq6K+95yc
BfTxfjt3A678D/xaw50IRGUrtHYxIcbb1AoFHz0WCcHsMUep2JsmHBCt/EfjYafi
LEvzm9qg+6e/g2YtXwsp5ZYFWFQ0fNloPdIV7997jxfNqvNbJla7hbq4n8GpBSZO
v5X3g6Jy56QGlONjugObiJy4rG4x7Z5YWStw3OGnxm48sURSJmVOmbk5a+bpGuE4
T0xlykLylZtNkEwq/lU0BfjoycgTH/8f7i9rCsZGUAtMUeMQkAx/em+I+XOzBF3l
63WVSongxGyHBWEm51nLySzwRLtvmrwOj6veYYIGqWfpzP9/4FBKAQODEAThkM8g
Uzvy5avpdGyXJ4KDZ/2FQ92PHid6qW18AT55rLhkSjE6Rn2ivhCcjlgNPW1pREui
538/RpWfxQ9qVgiIJ7irUpPwlNuXPa5qAQrr9Jh6sAQs+J1ncuqJ+VFyn7FZxfOa
0dQPjpdZSVjkega+V0gOp+4bVPARkW8eKaYh9aT86YqdyBRXlzBP5TJDdkFc5tPZ
BNB5f0DhV5YH6RqGPH+t/O0do1IC0HvVENoqnRg5z1o8QDx4hcoCce4tAl3kBf5k
I/K/GN+YGrCfUY/WcJVwlJYGUvPBDjdlvTAoxRRfSnLiVIF7EQU0hQbG27Jnb3CO
/ri8zRaCeNMUVkD7akwS606eqhi963DCZwqeV+CT5xyHSyE1dKE6jtlPJubCNv1d
59HfrjKHKGOaeXwGegXFV6BEw6fTElWLWwym4nYo1txTI1Igglfw3/pPn4gQUSmx
jyR2kizAkHCSOFdrPQ5RalGpNZKKGoyh6dDGnmBbyDAVFDw7zIQonpYt/Dn0lh7D
MGPyVjmw70GGoqgkFBKuu0xv3ebmgN36HfOYJiXMJrCxqHMsavPClvupxwAezJJW
YOZiQ1Q+VbhhdlmHcdp/LUhYWS9qyxegUFTfM+TJVuIYh/+PaJyFgI6BX7lid9mh
feS1eUBhcY4XY5+2gBMPVqCbjc3I2LwToMg8JBhL4XosnTurErfD2taq6ah95t7B
tKywY2keqRiBEAzFrkhS/HzqQZxXP6nU2jRWBB7XKsMIiYOGEyUQhKvzzjl0KB6P
mjANGIHZ/WskK4yh9S3R2NQTKcUAvHiqyJWmeqR4QNsOb9IZDs9mTWcFFC15SdlK
8oMkHM9mG+wlXIt8URNe4BTiGosS88bcT1kECZYT7q05elQgLY8n67uN89URksDQ
AoSldV5MEvHrzwbw71tODVQtuvAVXiiWhn6IMS4MNJqzhLc/MjJN6UoLJetE4OGx
+2PaJ+biWcA+Jdlk9BSKpDsEnOtsf0J6LT5Qu3+LDHTpKVwcPpod/nqAPB2Vun+H
VcoZaqY7SCAIlQ/mpg9IdWOVW1tpJ5p/ipzJ8hN7/W5PZA6xhaWTRdQ5u6SNWluj
dZ8szFnGdg3p2QHxCH3cA0pgxOY6zg2jZN7tho+qSRgqHnbKutPD38s/bggYRLvr
tIAFRlIsdSw1qj9uHYVdOZ4iPRQv+mdooei+rX+Gc5zRs8MG9Psns461coyyNKUR
tRDqqkSYpEUeGEeDbZI8pjaUgzy8TapDe8iGvX+zsCZIUZG971OIC2RpumZWB/rK
0II4doLrsGulqXVWsUUj8AoDbZlOALiwb0v0X9CTvRgVwFk6HIibGMl20XpUW2Yn
eeEoQt8sds90kFUAjHbsLQMlLBglX5OoKkbANM9llVp18WPMharHGb88YS5HHuLq
A8H1n3IsrmJEc7LfmLuaQX05K/6LlS0zcdBtW/YqyjGRim26eXGMgvKWuqx8gQU1
e5cfEDEoBpQBuE4N0XZBF+ljmAedapzm4vjH1Z8Kky9gRTjY4yEC3wjQs5ZxO9xP
WYJu0xcWv6L70B66n4b4TxOp0eW6zRZbXduGZQCPURyVbA4oTgAmzJgy3dTcKaHz
sNRgXA8L1chyQUP3HkBL/rF7XPqmlOSc3SZmLAVDhGoep37mbOeMOLkyQQ8CFINg
fD8TYWDnJ1LKK5F31pA1B2O06h9sQWTBC2tf/w2YzDS64x/AX2L49AMLSia6DGhV
sUZIVTbxQAXvqiPeo/REyf0lJxyB1Ql3xFYh+TIe8my3AudAecUS82pyU77pQCnq
kgkuN9fxrTfeCzA6w5AgLxoGQv5j0V+DGtjTJuANzNg3tjI/gJkKm/GSInQKImAL
PgHQa4Cr6XGTDa/oVXdlo0BUKkCSfnDU19UAxc80yhVFWlhbACGl8VIigVfNa16A
TDUZQyilFE9KleYO8nY4jtOW+muPbmamU3c7jErh9Ex77i5rmj7OsvsRwAcAMM5E
7/j2+sYDxooyClgrqTxXe5JLt8G+dy/9Nvt8RpTEqRLqGEypsH8TZtwn1BDdvQs1
kElRo2+LqVi7bnwCQ71BzGSgabI9eK+w1vqCBvSW/pUqzOqPOaXSOSwLkWmCkbPQ
23yZ8kzqqDxQTamr68XxCEgDMMh91JbI+lYSIoL+nepyd1cyi+zCJjHJJQEszjgZ
O2rq99nVRnWamzGmxr9z2TQHmvktxz/mE2pxXbFqJOwrzjXqDd2pZvzvZVJkJ5NF
zXEUSmv8zZd3f157nyvauC+8EgTSAec4l+kvhyqJIL/MI6IajkPUcNNIpPlhrxag
7nYvj6kUcWC/Vw0rsULDoCjKKV5brT2qm23US0Iz1Gl/VyWSt48CQKjPNj0MW6jE
s1nwat5VjSj52rf0qoyEsjgTYlWKI1pVoRHHtDzzAg43L3j8h5XZoueVeok0GjZ8
UCISv8kz4EZf3NrWNAD32dzVOtYX24F4BjzAJDS6+qlfLLaA++c7EeeDHYzGycCP
lReA2FwLuB7b3lGTYbMpRHdAoxUVYB3Tzo6TIiZ7fSZJpNiZWzYXwp/bHd3XLNj2
5J2zquWlP49xdxS8dE8pKqHZ/og1YmjmmKCy46px6hoMSl3nepS8Qr84zfYYkQhx
RkjCIsR0/DWPsJl1sKhYKcVe3KxuqQx5XrL4rgCjRI4mHqzTAF90Y5nz0w+kvZ1H
0wQB7RUe5/flNZZgRv4FGfDt79DCGqJxYCQXIuFIunakJAcdm8Tsc+EQFQLIBfro
XvfilHMGFGZoyzEQZlmaD+TBZTCnpAmtAsD7XmIM3oGXwT8BRIyundDqp7bvo5gj
1HVcK6ggTtKjfEPGm2IJtWrcMHgPUxL7YaiowXiLjjD/+cENEumPyqcjK6pfgLWw
n+dltDMcrOlHXYwtErzTvxXtEHReoym0qCO4dTGOGffI0VUu1JhMlggGFuB/F3r8
3tUmNp/wML3rHwJbHoMMjE9feWH4wpL9/qWBFVsANg2cXuLRAXyEVhSZbQUSZlYh
FHEwJziOfvq9c0DyutYvslm/5SAIHT7cAXpac2lDsDZNBTRxNDL8mCFoTtt0SZUv
VUtkH+JBm8o6LriAeqc5Y+lvA3d6UEVlRBXQqHntzotSr+rtJwjeLsHt4eS1Wd2/
j+Gp5zsfZMUGtP6H/a3B4BFJ3YhQoMsFvVhMVIFWNex+DssCR/uRI9ZBUSkVl4iF
UiO9Rumx+QkDG9953VTC3jHtTYV/8veI+GRn3tpZNqUmpPK/9f946OpOWSPiSRqM
VEjra3G9VKJg0p6Yms2CJD9TQcbRC1T26tg1akVrpp2LGG9oq6+PwZCWhDLqdtTf
zy0GR5Rkmd8ObrMkJ+ZnLTyxhqYcVUSig48mBXKaYyQC7SLUZyXFvqgdkpL12/Jp
P/6DZBI/hmNnBUThhTYv7LUfVn3Kwjnh4PqniSy43lDEw2KqAlt/k09CAgVOSPEy
i3ulTf+FtppVPZhk6YIJaRq3F2TVXRQ9nuVvPa6nh+y8PkQlIBBitjbRntvmJ5ix
w2QIIaXjo7nFnWtHDvnHwundhTJCpozMext9Gd2HodnH/xK8LtYx6hKjj+w+/HQb
K55/ARK2EBD4yqJQGdTyHX75j22I7dqqC3KjzelaHTFF3NFPveAhf90zlLbDy2CY
J4c9fyi0/lT5F2EW9T21yLf2HC1QulTJvbnsun6JCbD0hEfp1XbKEg2sfD1CtJA4
Q3DxQXcHxCQozjLfrwv2G1DyYDgp/Y9epC+BmX12ai6q4ZKxg1e35AjTsecutuVG
la49w3v5zmbmEPjK2/+dmVVM3zdqKsL6+oHBdiiTor8o7uXj9GQygX1FMMfd28eR
qMkoi4lfmSTxOaXuihcX2wm14hp970C4Jdahy8QvMVmmtu4CWlLBss4C5UMg7kuC
jRfSVOiXN373dfK4XnsK44skq4JZg63dhzslkQagieVnQlUyCQ7mOvg68IueqvLu
TVQgF7+b+gC0iRPkxBkBl3/SpnvzHYkLB0J2pOJYZkPWPVTzGa6J6nHUrA8p85zW
61oIsqwC5lfuICSLEGcMA0aOhWX4DP1gZd+u7CIR8wn4CaYrohvA6v8Hozs3+WY5
puX4fBCaMlTc/wY6xebd2Axxlf/w9d0IorkFHW+d9cUlV6kVYERQ5t13yyKAAvwI
uaaQfkbGZVF1TFqudIZ2k9CkyrR+J92D6q2B1urjrrSSuvBDXHT1LJbPQta9/ZUC
febcTngE1z5/72BLs87ERBMr2ZdaP2+sCPpdpRDkPjNCBol1Gcibz1MX0rOMx1rQ
ufLP+GRX91qQ02LDrq/oh9Lgtm4AOhy6JboAsDhb2N/WmaeuIg+clbiK86WPu26L
GZSi6o6FAOj8gwm2KfBtkv97cGPc/MZdj5Ey4ax7LQY1WJFhJv2RjVFc9eEbOn9m
xiHx0jQ2yXLXu5IRzJ0MU/oc+0IiB2OzaqDn2oyCT0zDm57mY82HfzJkbBvUxA7N
iWoK1gqxiDfIAG0YTz/apj+4iE+Jrv4WodNBiJfH+Batb/o/akZsNvGeqKqLlovU
9WmwOTeU8sKzselKPnyoUCzOmJYa+PAdRxwG/B5OLLEq2q2bqXQqGU4d2wc+rFRb
RR/pbMune+FzdPe/UZIG1skjrsffelfwE4J19kagUN1XDuiEq7uTM+MkZ4htwckt
fLcTtmjmHLQetC1+Ui/j8xbaaiABoem2yZknatDAalYlLiHLaiI+tY9KPX7/DC9I
i10KFILtIWjn2S2PdLtMR8RRpS518RFKAn1KT7oPRBdGvzKFFwv6m8XUPMkY7jGe
9EWB7vFx+tY+rB1m8HHtlgr4I6K1fGYaReCvAQNmKQn1vzwtBQyC5QT4CWnz9UcU
26gJWbJhj9I/cNSCx0k80hlfx+JjzJCI2pmZZrMwThCYxOk/4hz9upY04+xvDXVS
CUiCY4f1sIhD+R2o9lp0usT/uLxaw/kxlyGz8NF67nTBFGlQsLomr7GFUub4qgl/
8NtiIy/IizycDptvTUeCUofGdlSdHXw9ntJ2JA2Wnui/L/5o2kphBFULNHdde6UV
XauTQlD5Krcks3zRUTN5zOJUHhZ13nGean5ERefldSiCcxObeZuXEJHr2VYUwMdC
/qppDeSgfjQ7Ds9NtYKDy1njq7QpU55reReds4WI4OzzV68zlYPHI4ZFT2nXczhA
8mnPcHHs8mah0XrhjGQBZ0sJp3J/PTonZy0kbni9nK+pZ2Plpin/6xJ1gGKTTMuh
ClMEP9tMk1BvOX/vU2k9aBK81vCC3sazs/z2eBQwjpN2jB7dQUui7jJpTQ/8sIaq
hRqd4n4w+PaHFDF9xC/clMtvCIIzaqCHLIl+//ppCSwMNXtpb6FOQcjCuo8foAap
IrrUQRRK0M4pmNaTQZN+F2mQCh50lOi93PYk8FHxAtIdzSfYmQqCUaFMkT3bvGoF
eGhwvKOGQjyKzSUdmmBxEHCeYY8mvCnzHS5rGdjH4uf/B6f4kuAKIiOQnjkKkiyJ
rkrSc68Whrxs+tzI0i92MgJLWGBLEcvbD3dYuSdtn1GrwQoWTp76X9cmXUSasK96
N3weIBuLhF4damMZ1Bg/gcnU81T484yOrJg8o/Z2d5xvtrD6Z6ky3jpTC/E/x5Hd
udhg4E+OJ2UHXm3ymOBftOqXo5IP86XAQl2//RCqotCmb78UuGsd8WerO479c3OZ
rMeRqLuVVQggRtoR/OdkR8iPBKgi+kqT19SARI38MdtnH9Te0eME3YC1l2svazyC
UMCD0k9zXK+nqErEyaQwXSb5ynDyw4IfqXvt6bN36fXGpNAXU66G+QlpHaB/DMrn
PmpqjqYkKAcz4JrNiykaej/meVi+2h4gxM2oBz1tFGa4y/lOBqADOPHLrFCRWLXz
jumZhPtCIlV3ZyCZd6qzj61BybhZbrXQUhHkgtpGmSp4vOFWozjK+htMLOZ5h7Fe
8vLNnBahjIwmu/0YLhplmLDIkMy/rt68MfPsEuinhzKUYFzhrOsEc/lS9dUREEz6
nL+55Oxai1psOaK2RAx2K6dzqo7Dw92N4M3g5X/f9xgNVGRVN3BX8WsPrENi2Uxm
5LyBpfm7LmZPZlbt3ySwyrnhqnGEQRGRBfCYa5Zx4UN9eo6MBgyP8F4qyuTSuj2K
nHt/m7p+6lDxqqzEfIB97V54xIjY4VXQBkFUQCpgEjXF+Z09ab7cKV1p3zG5LWtE
5dNY42qylAFY7bQ3N/oBLHrHpa3wW62KdMH2l0rVLRaHCaqaUrvXuMC6VqiNl5T9
9MXk8BWODP2/Beil2MgWca1xKVGDuDY11DEhi+HorESsyNHmEPI996S/oBfaBPJY
SJBOr16C8g6nQMCxFcHOGR3mymcPCHqwqiZgPWsp59o1IGgaFeyhogfJFOwhFl/F
XIgBvZLNpu5jwxaYPGBq3LDEpX0GllhSpRufFAZ1rFH1mLpBAhV9BnOzT5Qw1Pwp
Z6TfMVDTqdivqD1sgPyMHQLuXlpHxUj59s7/c3CpEUSVyDWQtARpiV7FgjKR5tM9
H5PIO744jXcE7yK4XYtxsBwo0z0WftNkrxTGFgWBe+Dn3B1HFSYy+C20qGmWhe6x
Kdr3Yr5wk1O//iLROb/Yhbr0rdg74TqpGJTBejkIlMVYzYkCgUROEtkLT6EwqhFW
CqU95c8loC1VojT6XOyw7+Nmrq/yNjaDV/F5oYBuBI1K5DgYfyrvR/X9n7blHHZ7
KN8OHnwQMQd0FRntpUBy8WkEyEUZGLK3urLG79RKopDblqumnv3ZC3p9ZaJRrhq3
GSlyERuPDiBz/+5Lh7kV/jRPSonVhlFEoOfMsu17uYVEg/fuJFm2WxhJH4rxGos0
4LCsIv58kKA9VEkD8a8kv8VgBzoTWJwblp1S+ethdcgWM7TY3OTaUcYp7VlueLfX
167CaNa0m9SvzNKTKQ1L5tr9lqeA2jsLXoMQOtuQTKxRBCTLEnmRw1ENO3fBxdG4
h+Qev5ipetIj6obxZ6OT//JdrGAyuUhu+tYj7Li5I1H9K2dxT9O3I+kS6QRIfRMk
xOyRj0hgQEObryEvvTTjId0SBAORTnmaeogwvGeQ6qBdbsulnO1mmGYBfP2e1k+t
bjwTSTRc7+EudQvVK0XJFUVxNiScPtp5BLZjneoENwNrebP5qiR1GnACvHjL4ie0
96N8EkxkbMyXhLDlvoR1todW/iPscazvGWLiolGvBUNcX4sYaTuF8qMag9cHMvz2
WUzAtUoTbXBTJp9ujvQVUZqK4CFkQHZnqNpDp62i/SNqk8YC+XXhqKJmsJY4I1es
wesAi3k6KSJ5kbKc1OzIIGIOw85B2DWEUwb8K5Oro2jTkcPw+sA+MTt593+gSZdR
SZxpJErtrKCu6d+3hjgk1AXxZgni6ROQtdxFaS4t2NxnCI3SVpfldnC0jC7wyapP
ssK++YQn/976yue6tp9pENJb24K2Q5W1lLJKp9LDU3jKNq3Gd3PLnP9CMmofDTcZ
GrQjPSA162fjhicUIJf9hKu6J10TiG5PCt7ZMfI+yS9039XmaWL9j+v0j6KFu1fs
DpxRrByWzYQla71lANXgCDfxZVDQYqfMw4nlgZm94MLS1nyRmf71qEWWFeSLZx2G
3Eg7pJV6RcFjQ++F4kE07AzPm+5dYSKBG6P/rVdjVYzc9AYwoAfZNE8ulf6EQZOl
AzZ6jWlpjV+GV4P7JqqxE4+wyKOAEs0Dnj3OykWt5NlAoPhnt4q+lfwtbDwSJFAl
HwpFbSjTVi1GpZYwSsjAE+jCioQJlkCSpXw+OS/yPi6eb5XaMVZj+C4TwABacYdm
Lk7lMuerGcK4Sc89pQ9/7bgCgKXRRkoa0Py07e/ZFigHctydii728NkRZG8qZk20
NZFyDHny1HUO6AajWcpuP0x5B2KprfMDAC3WO2rp08MdwhaNZR8k+XFPmX27vX+s
dkghWWtPhUVHae8uhvagaWgmYPeY+xn2E4gqHXLLXM5d3BrGGqdNHU+RZBk5TYnM
OUfeqVcffXM4YHqDxkGNoGMhtt3I7G9RN11d6xnAwxWpXZCRDJCH+trvyEC6jrsj
t28sT65fA+lVtPKbU2EgOYUpAkBVGeCmHRQcE8KzSBHKEKQmoL47PeT61+AxSMXJ
9b7wuZDmbiPaR/qX77rOyGVHtBFASZmOY7IRf76bpQL7u1Ap5e0p92tUlc/BwKQl
ZfUIdAAisSGeg2i6ncI8Ln53D/sZzGZFP/airNhh4VBG/vieps6isZnQtxU1ydxA
Y3B1d2rCyN/kYy/L+uEykCz9HVu0OVXSFDMqwW1EB9XiofxpvNB7rfYWujaWsxCF
0T11Tme6mx9ZDlanCeCLJ9CuIAip5SiUljN8LWTPMNGKOuY8cTRdBUJkIutUSsrf
us/wtB9PEtz7mpRDfgVENoqoXY+GATTE61NUCd/yEEmJXPaotVT8Pj0RvqP9+89x
G0+kTL8a69NFzYtkJ1nhwptEb/eaAdp9jgL22fc4UKiW0kc8GEWyzllKUYEQlbtC
oWG7DRXpuwqAYMaZS1bakHUTwfbmXQB6nocRIL1SBYbCxFeiR81Eni2NMv1MuiVX
86H3A3BkhjDgLa1snxKilOvlqpS33vUB+0pTIeBHF1DyRK8Z2/45NQMDZcCHwXbN
YNwfgudJjEDbIWIwwKbvvjDzaRpehhdy1wnrYPC4qE1eUABsSuA8EDkwlibkqTiL
df6ve8mUoOa7RVUTbC97zTSKINQQ4VEa3h3izDL3p1UNgknR7VGPE9Pl4tNIL2iZ
tpfKUTr/q4yo1SnUVv6miYjzwRJIgMNg187GqZe+meogve6lOQ1/XrABjpyBS9DB
+1A/0e/9pczFHl2lSnckVhQs3RN4cs4FXBV9t34++1yaY9CifbS+gmzhzc4wlWnm
hMrXTKuYU3WXJhtcWGzKOy5bw4TNwlEFLhSRx2eOd0kZXbbdgFsGJ1J/GtIezmU3
c8n8pf66mn5EFyTv7AivRFDga3claMpTH4l3thuJQIERi0OsKxG6UbXQYzmsoNXH
RYqtNSlN9OHGbjzWyBbEhG4gG4NsPOO7Mu/Wd1D/b2vVeszthIHaNOZH/+jW/Jcu
oZH/q7teUew5uAlLzykifJpdI5jgR0JckA+ExyXknmxcC63riRzDZyyU1fCuhmn2
b770eqxfBv57IzxnHxyVn7abjcNE8n9QPg/LqzIoSzCPweXDmbRG+DB1bwJvaT/b
1SHWgLn5fXRxMZ6XGo8+3Y9PSxUBIi7kb+z36llaSU5N+I0w/e/enX3aTTMKVT7N
aeRwhV/rvjhxir0yZfgmoC0edZr2PbYF+i3SbfiCRKTiWvbY+SgW0qm+435poT6v
6Zia5QD0c8+nRJ6nqdegelZoXflRaRgH+wg4P219vQDnxH6dzs5auWdzYuZx+jdJ
CCczzX5xfIWH0aEldr0P1rnIZ4IXdLxq5cG+EGUlptk+RS37LAx5qrz13Mwi+Jb7
9EUQklhA3yw/XOiBLIyF0aRtdKFJEqV4GGtQOJh39qQ2Vidz8Gpw9PXrXWAmCkQD
CFDgVk0+hGZvjjRJ10iZoDO5EPK5lggT1EuKGnnW2JIPf8jl+0aqXAdTNI99pIvL
BH49Du8bgynpZzbRmUrEQ5sL6IJ53aSlnmvBT0KZ98AZVjYVljV6UWX7AmH8ehZz
K3V/iFr8fhvY+ZdHc8Hoilsj2c+e09dyFsNyY0r1A6nxriSt44RhbaaxbNzH0rjt
/31iACdoNHnsap3XlDABkzs3rjvOASmbtwnfZsBCmP+Xm+b1z+VCkKKRr9ddqlNa
pCxyCer0w9QDsJJliMk9KUyO8YGJnmYnZJNuc3cvGNzMGqNtIbGx6p1V94pKRnKT
b37MWZ209jc0xBAwz+82Il9fF1jUOJ+/eC07TX9Iy0OSzVxPfqotJDV8eFPoaEL3
T91y8DUjloPOHz/9qkxJCzOKijZc5pzXreH2yg2e1EvqRlO4N2O9BPPSVW2DYwzF
CDLsNboE9sx7L6absDgoqoom1y5V3m5AGxj6vCIjgB931l7Mtat0QFDFlpC1xEUX
fVWyRoa1mRTbUgkXWCvi7RlNMI0VQ3YjQqQPW+wKdneaCaE/Ckv/mPU/WIGfhcz4
dEX0F9WlOlRQ6pqJfhw0BLKyUFNo0nHFmc/zZeBJMrAHpjmdpAgpyelCZJ+oHDhz
rT7/6+fxhYS3r4NtJZC/0Ymjz/TD2uh2WatILAyIHkASLdWrKBL2+wtMdSrYAe79
O84IV83HA2tVszw39HiadRUAhqnmdD/ifkrOfJGivu4l/jppBvQDiz92uPnZzKOD
XggIxm8Px8x+u84J9lhBVCUln4r6814QARDBtMAisa8Cz85ZWHef+iajGx5dkNVk
aWYJB/CxCf0Le6mpximud03kkJ4+PS+fvtCIOcNUFWhZhKjurPHCRdB8xT9/asdm
c3rIyz3T/kwByh/L7Ytl8yAKO1Hq5bJRith1LyZ31S9gcBOk+/cFM7JpcMwBuF8p
pSiS4lMmM9Eagbrrr/qxIFfeUbW0EAJiKyF/30P0rvXj2vHUjarjVWCBOadiuNCS
csiGlnrCKL1CxhDlWhYIlH7ZU+40TT8h1Mwb774iUf5YZqOvyIMRqbl9o+gxmSAd
f3roV8GnsLWiC1FeHifNL2HEXy23VFPFeFhB5Ryf8HSLqFGAt0SsjLk2dvxxFwaX
e85dx3uOKXDFNLD2iQ5CP/UoZg8skbswtXphhNL3fA7VaT0wJg5gkYSVPlKUdcPT
BgDuOduzTvpg4txdTVLqa3+qVfXhrCgi9f0fPDCcluwruAgdpfa8Yb8KlBjhRnkc
6THF9izGCcQKD41rj81/epMjdJrQ43u+pfjkKRr/M6EDWKbEAoxM+Xkz/lLTrE5x
fpRKs1+s4UclsBe/wEe7Qi4j5eXnDmLfXQzlyUAf5X+0myRnAVFwo5xXGK2ql80x
9I4mPafZuDHTISanUEtP7Ji396z176mSbnjr/iCJe6CMSD1c7+AopU0Dq2eDD7G7
UHDI+12fFW5XUs7sTqVnbDuvtqceTXBkILQWZ85dcjBFZs81OebDBapz0dVJPL4x
Gx/pfeylCK1t7vLNrER7WuIccVwCuYPCXDK1qhPz/fjTP+9eg5zrT7Zrhfsg3FxZ
rWcsHEmD8ENqWI2mdwptDLRT5GXtRvJecX/Uv6juuhu7ciQh4nisJoCRQkCTwe4R
bmEnpt4hZB4aRh7A1j7pZIIutQbyUlqMRvEnZcn3jz4QNwYP6vT1Got9wGCV84LW
y9eXmjDZsYK9FMRpGND+4jSS8Z3OKw9LouMYQ4cXmykgWsLKn5yWTQGhrCDoVhsR
+pt/2tHjNhsnasV25sJOjaP0zlcIHbhZkau01NzwUvT3pV/RVv/yPgGe5HGvbdno
CSJVgc+YS+9OuAVxhil4aypxIwBTO3tKJ50QXNle9YJpTwlgVnkbHDqlru5ptJY5
NkggEcwVdMq/0U5jPVmp9OJ4BLG+Z1Yz7rOfR/vBZlJwBnMP8swnqADtMPlj5RSd
9fKbPOf/9PWdoqKZqv07wHGION6Sp7FdhgWdjw5iWTP4ZdRVwTfxKoRp+kMwXzYI
6AIxT1NfxJAfuWVZRsZ/lKJFbq8C1hAcSJOKcNxl+0m8jp8PRzH6xzqUq7F27dsX
YdahmCxDPsL2FQeXF8JUQFEmMjTKMrg1QE7o9MG2pCxawgMQkjJvOAvmqrLOyPgG
jvaH4ycnE6HKPVOepaNSWhlU2F1r28UVoixltMauiIixEXfgz2SCyGueVAkzdMh8
6rhu7TE3oRahH+p3Ej/x0cDmxbSzm3PM2daZfeZyM/PU9QS983yTrM+2dGQlRbom
aaJ418AXCIKo1rgk9putR4BHrDWd1PGyS1598tq2bFMdHqfrQoraWeZch60WD4i5
cEfJopceVaJMSFsDYgaJRUWaWI4yEKE/rZhs98k8SpofsY7AezffuoOCQgHI6Mue
FG3TFUG/4onVgo7i4AtNxI/JjihPM+KQAsFktzAO06zFOSMWV2x4KQSvI/wNFC2Q
nwz8rsUFrGk87obm/BGgycJi1AUkXvLy05AVillzmYNCEAc/PsLpCD3SlKsUdL3r
kRy96TaSWlyGu4FuL/R4QbAuubC2E7pGb8VMLHcf0+CNiLNsQZcOW+pDsUxYOAsu
T4PEsUsNZ428mOjum7F+ForXkEXo2Cdc0bzKbsmhHCIxhNcyaHAdZe+0T3t+PIKK
iGmp7ZHH6xdjQyxgYlg/palPdKcpSyeRnLbfZ4dJb6iKv+bGYRyYMkUMRhqxwhVC
ZOzg61zLro+svaLq9K7LwWRPubOOFMuO+yLGNlTfbgKRS210QaDfvMYbMZF9qvYf
RDfRvjE/3q28pgc6san46X3QmP8SSywYHOw2onB0dANJkpcg6fGutQiH+2572bEi
rS+Dizn0yIvRtVFTWBjdqZLmgTqOQxxuM7DlWH7fD0NfofyqxkarwcdWp+/KHBUZ
hEWZlFg61tPpDgNEXbV6PJGqoq18MKrYHdPuDLxPyT1h/NPDuZ/EAOChPpXhynAC
o5RT77TZVzldA38UPUQxwpq69iJq02dSF+DrGw/sj711use12A834w/x/UuHKUeP
K7L141pUNnn4vxxQHMyd0fPyEz2srOxaWwwNe/NU5h/P/rkXBgdVC3L2f/0+wRjC
2q2rTQdH8aqQX192jnKYzlCrNlr95642IUBoMy4kxO2eBU7KuQpEzPCtZImzqCfn
vYP78HYwUsBL7aV1ES2+0AyICEqsTqBfjcLKMBtL65maTD1qMS2W6Um+es9NOyRR
jQe3lw1xEby3J1kRfLsbB30FY/btbNDw6OcTnJtbL8nEo0IyfxNFRkSG6bYJ6OsZ
35oLaPDV88XyfNq7EfYDkeaz2rICkSv0lvNhd8f5WyxM4+8LjlUCD3zwKdiAc4Ux
oon9mQbnxGIjznvxSpwuxINS+poyJySQBiw/BIhqldzdytwvVv8yjvH9MSmHYTuy
a1K82sb0IpLf5Buo6Wl/GbWbI2KF2wc+3RcDfwoiN2T5mdGVk8MdAVaSQpprLyNp
uB6StzzFrrbcJ1DslHkZaejsX8+hQOEyiNBnZTfqqiruf2MHzFlW8vLyneVbnOp2
rpbzyB9qawsfMa7fuWRRGulpEdNn2NMGOTgOMMD86OXYOokJdXeKHQlR2P1XCqhE
c1tPvuWp43VX83IZTx8aEKUdfTpTkla8yCivYNkNc1opiOuOjPMHyWU3yi/z0wq6
84T4ku008DQ5DmuDvg4UVF9Z7/2kyhE3bvCBHEo49G3FyoDuWMl04JVkCHy4ybha
q57StBlqCpXyZ00hw2sf5J1mfh35d0Aph9enT01svR0PqX2+9xtnGk5yRCneOH3q
JVNgYR8ZKMI/uSWCunV6ujcvCypQ9+DveY20omQw60k3nkgZTuHvyuYRA9OCP24x
OzvFFk+YeGINxB7e74WI8bFfi/oSa1A7tfpVQ6ZfavI16/QH3c3pRcX5K78BoUI2
vX8/Hs+mz974No4PcwIhA0akvvzquDkT5hRbZutfXFjzWw/EiTBwVQIriMBsjeL/
99pyK5C57PeOzghvVWpxzhEumGq1wPUZn8TGjepvJuycpSss7ScqOgr1ppMY0XPT
/hP6bW54ZK2MOX1VVziJSj0xCdUYvQ1ahaOVtb7/PNhXXhYZzhOeCkZmDdQCgUfB
xSm55KeJTfb/2xvEw22l4x8mhN3b6DY1zk/G/q82p3Cu7wB4LgsBYQAquPGfymJu
M2rEpmwNmKQgbEDxFep1Id2PKEp8eRnwskdIJMmfxJZ5nkHey8eUBWgYs11egvGY
R9PYCVsgy1WtEFLcuzgNxI0FdhUDRlizZhIg57QIwRCugms1Zhm5KZnXtL4WPDQu
VZ942Pw1xuA6q2EUE5GphgRxGfHOhlvaHcGwXTnAVxnpx0wKGbkcVzHlNZbHAhLV
piKtLnLvHgxBpjae0rjnslAsFNB41EfUF6qM/9mx9NADdLW6WUft2jUA9L6L5kIM
BxzIqAkl5uOwHUlsKKZP+82HZB5MsoqXT5hHJ//oSimVRXmZ4UdJqGpzyL6RxclR
7R0xg3/mMGfxJzqzagBBdardQMC9NZ0BNY2Bhe5OhJ7c6Xs7vFRPECjFtZ802YbD
O+7ky3XlImDAuhjtbPObQX2cuN//n9EZHnb5VtmYmWl0LTbtA3Gkl9kw+gWWWUT+
cULr8eWCgxSEKqXGhLuZvemFoYK+1GL0IO2G6E1FsTxsO2YOxZXZjrp59SYjo79h
q1x+v3oswbN5Q9XTcO3MNOqLq0Mtui/+ZJiyD6dvGHEpq7qFiY9NTzh/otKfGW0B
8QPOsi3XeWZYac+6DSCd0PqzQEAyeJlk4ZT5KUpQ0tKdNoGhxfSViZCY3ab3W9d9
0DW/rUzerCwIkDLPJJcZBhWjxa7mBxnoodwhVY1ZE4GBuNvPyFgCt+hW9Jez9t4/
dyDZw5AtMPiTco+IFGqz5nRF2hRNq2OoECRT+7CJSDFOuU4Cz+ecbEXHEEeYQMDM
8Y7YkwN4wVlDSUb5KypScXmD4OYJ7Wc508AwSoPV/mwPqxAWkwXbXNnvUSYT73lZ
sW2Sxihx9nfiifn/v49RSSQKFTvVlSlXpCtXYT3JN53M4Wj9/GJgVBqE0bS46ksm
Ze2e8tMj83n2QbovOK+bWVPP1r8nrgihWIvodjJ+8GRG3Euoz1cupEOvaLykjU8V
E0wSA6A0fylfEKoHsMOH4sCL9cr+r31Nd7LlPxyYlMltwxkpXmbQgDv+ZX9+3qtK
DMtCftTy4PpECiiw0QnUUGwpShe6wd6f3u8sw+e5WizgS//XFNbI9yR362YpI77W
9w57jxxos7eg8IejfGANu95aUyVlsTADLC1drUoENup9/g9VPTlGNfXcOttp1vIZ
aodR5eaN3En1XJMiEG0/lY2I2iCQVwZRbWH+C/C9Vhvx6PhTivF4gMqoBrCSSDgq
Iwf+ebOc0+NjnJqaX1YZk5a50Tyr1447WbFEyTScDg5wmaae7N6tBgvAhbksrvTK
HSvzT/p8B8/+VaE8TjN7SNzhx0iJYTqTg1pOc67/eMIg9qLIAjiDioV++zVP54Yc
cG7CEi4Os7LNAzXgEwSQZLcg/GU+KO7dXqFJPDQVZ3UI5WE0Hj385t7KvSUkl0Ix
cC5otMqc07istz9rrnpwgMpz1I1hvQTfTKknv6EgckmtdFJEBH3azcBprW6vz1Ju
prX77+aXp/sTMEcIYRi68mBR7zZy+IbXTA+X3+ER77JA/3pAC2vO7oy4FQiE4zPu
JkKApjqhagu6Kgvy+drVzd4MAPIdXgCuhM1w3tBkFylhZTxeLe/pmnPFN4/yejVU
7CkxcA7EL1/NL9jV6/5sf5i/Ucp8ZTgQZMW/IRJs+vyKF1XDobp3bBXkIXdHs37a
GpISx9kfCx0XrMZrQ4oSp+XGff0ODSxtRIRsIv8EGieXuz2HycMXLC9AOjVovvuh
2eu06aythpAxlsjDaXbYK1zO/WOUkc4qEG4XPQdTQkEmX2foJIdeRwYVa8TO6Nz3
AAs5D4DtnUKbioBfrgnsA9dATQrGHiS34+oiEY3LMxMN3E/ucmM1xWUTvPXcN9p7
O7B5CVhpMBw5Vp35Be5yMu9T6PbntvbljQtRhVI4GYvhD/z4ncgofkJPj6btdjMg
4fs52K+5aOVJHzCNky7TGVAbIUbyzDGSgUpJ9ZZahB2Q4nu3MHE1Xk5HxYNG6yjQ
xACNyUCUJV3mJ83mg5BmmB2AMKM1kax25bvVB1xnPBc9lKNxbvSYH3/hKhtzDSUb
DP1DfCvOzblF05E9d5bQblWDw1qd6iqXzhAGpq/X/zhf1B0EliwkJEcOGESAeXgc
iHyr9Hqe3rRKO9wZqTG14wNe6KF6QmD35Lij/RZcPHY06MBE4TvU4q60tBWJ7sRf
06JQxLPhsdm5oe7he+cSfqy+EGqXhT6sOcN3Cdu1PA7FG8souVWlaqbs6+QrS5Ek
0Jl37W/gtssfys7FGYcBT59bZnDQYf0sTkMKMNlHfytYUwc0CEG1YuDPbjOMbQxU
DLG9CHFd3WP4gBZ86HS8S9NTBOVS+sTjsUWEd6t/+bPzv5Dwfu9M2sKULL/YSLHT
R+EEXeZdzFkcgDobJcGu9UiOTe7UMvXLklpiRkqYfoAZjOAqpxg2o02QA1LTpgQ9
4+z8EK+2hTaAzYkSrCLFnOnbl6BvhCIHCcmh6WkR+//yA+JPztegWZbiQRtV2fe6
03tj4BkXc0nhzfvx28C3q7oLeBEd6CbJiuNmZ8aFDrS01XdyE09YCD6TD8pVF5Dc
tfiE22Zo9vQ2oH2oD3Ueef2NIPmmgHRnIV/RB2Q9cSkVeik6xhqHkQ/IEYQntxbZ
m+Z9GHIsWx7OQHDvOSy1EWwD55BS8MM8NpC2q4EwEoKyqtDQ91xbJi4Ydrkl2XEn
CjnQrO1Li3Q+y+07NbUANKWlIQJYx5Bqc2JUbMtJdAWEcJu35cE4CfIxRSRlXln0
f2xd5iYn1/q36aObErmOXcfmme0we9+PGbdJrFrlsaRxRtF5+qd7UIFw+vLCl5iw
C84W9tiJqaexwlwQAvdMEOcRPEhNvDC28MqqZxgyb43UqvYmACYyqNZQEuCxm2XE
ljjLGJnEgJbCv8pGDHaEWcLpde/Iyfl16PDbZYRvL1QskNpGxI+eLy6CWVa+nN/1
PxmLvb0D9D8otjhfBmCc/NhPxMmCLzDtTyP1n4ALqQo478l9gG+cKksxgWYjz6tg
FKeDaavsu9gjRqt6cKP422yJvlfVGxPUmbmh/E4Pi4h9kdygmjYwK1wFkMdPNESi
D2UP//T8KhLVhdIoNE14Lp4KnLhnFm65gAgS9psrawo38mVhHJ3LnP/NjBh3RvlB
01Botp3irz2wIzgD2wE3vSQ6tBWYNiExaIWceIR6sc/R225Uy2OcMk7Nzj6lpeJ4
gSy6r1qozdXbAqWR6TQfWvb64qrSHep6Bu3JY0ENYsVtiMkp7zOF9i1AOhSubcno
qt/QQcLiGbbOKQnvfG1ay6n/NrJTEK1I5VGdYCGWvx2uqDnFjgFGQyxE/lyRMxJB
VlFOUV6FPrBSnzmQhQ/pI/VPLETcPABrbE+GBjI1vuvNEM56M85EIgs1VcYxHeZu
Od3IXdsvC9hMQXgMfJ9uYnNCPeUH6pQFORMlr3cL7VYlxWkYioZbq4QwF/Bik56w
uTxmb3sDu9c6m6SCqjsuVIFrcdaHngQ7rhO3RsItqRiO3NXrZGnd8xYmexrAttMJ
8/POtj0hOcLY2PYT+P0+51icXqy7xtuzZVCL/dnSeDpTutKjz6rR4kiUj1YiACTw
Z4D1YGILo+eblnoDM4WiRsh8pnbCuQtFOrC98XH0+B0u4Lh3Vh4v9DzRNkpT1l3e
VCNvbspOkIYk6QY+Z7Mq9necfskOgNQtyE9vQBfB9SpdTo+W0YLmqVkqu7beWFbW
zY1CZDW07uksr/Hkacv3npoQPOs7dZu36IbunNH6RNhbjmv1Od2Zsje0Y7NCViVg
aBMkIPcJGtSClrsPeo9CoDXW+1/vD0PVRDg2C1kCIYHuvXwmS32xaVBKgeFtLnI0
HZrFo3llVe+sNRiqCk6ILNQ2vKKoh9PavPXpR4LOZhbhXVXwjJx10lr3e3S2bsqG
1iHr8pAkyWN5FUgVFCahQmEngNe+VkxO1aZ138TjlHE0oTM8c1Rle/xD4fbn1ODc
oqU6imXzu9/V1yH08swhe1MsxSC6FP87M5oFvzwrgcg0LmWLY7bwgltFo/EbZ5ur
Kit+7bxJ5/HJXhJqCLNoauySklI2TXT8SH3LGxULgjJulsb65+tALAfdxo8EHiHJ
jKcKP+n+g7P+Ontn1agq4S9kpWLg6zhputWXyHzBZmCfLo/U5HuCKih03EKmm/Ng
uO5Ne1GTccUrfp9mPjTQvKBpLp1PO+kQCXL9gBMbQPDMMX1Yf2FgxaiO/s2PaFPq
RQZvTwv9pkj9sdSG/tjOdPsdqiew28tebC/E1UrzrkHil5q7DDL5sgEdwh53H64b
QhRJ7asWESXfOYIRIPABpYsLQasS+9VHpjyHOiS3dZD+8W7fLWvhyR1Z2RzBB8XY
DEwGE++14gJk0KRsyK0OcLmtRAioTafuMTcc1yUvzXuy4+UHAbGQLcLFz0d67jBr
zirIeqIGA4pt3ZOLQ7TgvWcS3DosTApHWx/qxy5ss+HlvkbAiVY4QE7bkSBGB5em
JN1XskXERpr9t1s7cLbDyapCmKgAFSQu0vt02chij91tLEgjUjoulHzSUGKAGDkH
rIJReXbx3Z84jQznFWktjKd2GA0goOh9jQf6ApuAmGIE/eDovAFP48vthpTgoCkh
Of4er9xuYrsP58cEKUXv4PZaOuiZAZF13cwxS7sAhWEbSajXpv05q0rBpQAdFiLq
CXTzqfOtk4DqwaYQTOdjf+71Za345H85o/Z90Ksag4YjnbeYEJ8k/tJPHfmKCa7z
EAPr8SXwhuxwOhB6AaA+S+Y2CIMqaIVPiAnfhvbKMUVaimWj2JZhpH2+pMF/rWsL
43Y1YxffIcapNdDpXv67jcLRWYxkWBuPqjrsl0Bg7yuO1Q6UyLyT1bvHc7A+p8+l
QCXlpSDVZX2Axoy2yxXJkeu/HQU425b9tHerz/d/hL9vms0XppHkjehWPGx0UbD2
2DkuBH7U/M/73Bg2Ao2ooZZTDHmcMgDJ7AfD31o77LvPlc3vTBksTCCLxUWC+upi
oQwgUX23esdOBSp9jqW9Nqol0LpsCOIKPVz1f7Yhqg39ybqZiM/kcsnH8ZLDTvBb
jG3G1SLly21s60LhLfRMfyG/V+ypyWLktqFIulFDoi27npZdzrkRKBy/a4WibyX6
Cd7s+83JRLVr50AZkSULk1LD95aMS9nwMRHv6CzCenQKCf+idXZ5AACwasmPtuLe
7P+fFgprKkMQcePQLFU2M0Qtefyc56cgWk5Ipkc/HBS3CKbH2DHApHf/qeP9F2kE
EPzk5B0nxfpF03jLAqITyn/8EbPdxKKetcVuyPx66LIPAedYshvpYo0MchDqXXAR
1YrRfPXRXywb0uUF8YkSpWfVBy8DAAEUiUKvmRyoKzjP/dCqW74nTuwko+7pK9qV
5jH9jLIX96fhUpJ7tWDGFVJt+lU3rfu0mk8o2lei8I+0BhIFlUlNHA+pWGyr2IYQ
a4iYqK9SZWj1CjolY90WgRpNhnlpSoir5OzQZC8N2kTrW0vOpWhsrDMUGKBIZkhE
iMURwUf2Obf20XWiGfdx+Cf08JBDp7Z1BkBVKAggSr9HROX+Z3B4fzb1YxdxL0jf
jifciaICmA3jQrs432m/69sUy+Q9GrEdLs+ocQkPnhR5n4fNEcnVJUgdSJrKJCKf
nkT7FGEuWisdI/r75lu6Jq7/RDHMhCDOkB5a730WHW/y4Ax2ovmD2r/zBkzZ0/HA
HtEuApqixZmSBgdNcXC6E+kGa4SCP6lJLuzhnXTJf2KqRpYeO3AR1ZBoT7pJQqeW
GGXcHQ/j2QwKT27o4S2uFVQN3IEB/VIWXSWZeXj+2d47UBhOjmiEgwICJP/gLeo+
I3kEuSSdDpC39r9SH02dGuO0oUHeeAfNeJDuPzRXh15+BHuhR9avCRkh+hXb5dbm
kXxCg3K+75nbrsejNjLo9tFfI7MVkRIfb6IqZWNwS1NzsY/ME0hYh2PWrs4/Kzfu
kinUxLI1vPJtbleROercfNK7V4/9Xxz4FRwOyurvTm1RUt1GcecXwjDv3qmiUwUv
2cpeFhwQSI1tQIWZqISNDlvO3okj/udFQNxDzChVZqZWOSA9R5AFMDAL6WUeBHWu
/PVL1iGNRXyTkJyyTubkw/5mVhMsr7f9VAwMlqR88CULjAfdNgGPF7AaSmTQiGo/
FQ3N+l+IT+aO4DuFN8z5rJqNrNdVJQjgNS2EREPLbC/CKhxB+L0qPjeSs4JYkpbo
EVCsvCxQlQiYEtmmDKMI6eFj28ovtz6YplHWgwGEmH3uabacHImqFWt4ga7yC719
4SWQbdW6eOXwlS+70qcvKOBWp8smEthAOgMXBh8iNg6QduGcayU4rC81ZSPX4jbz
xY1Id6yuP1ynTmljDvnvqgDPeYllnt0rdNL3SuxAadT0qoyZNqtmtnoRjG2rMIkg
8LTkL4oRi4L9OVmAyDPYP+sLz9EhbxUi2XB/84cM8s0u+C8SgPSkraqcpcRy/lek
SaYcoP4C++8+Zy3pzE7ID8o2xYDBxselawuW3BTkD6kY3D1dtwXiTki39RxD8COS
ZDGoHZZgwFFqd56LjnFSypFJYFhkCOhMRvtcghfIbFvtKMtFta4VFlqC7EebxYE5
PlRQTaJ6ayyYQu6lwcqOX/Jx7NhX5G4Ruys7Ib7UBjXWA/S3OgK5EQANSM7X3uHB
mvqJMcBhZ2rjgBSiVcJCN9g6RP9BtYogXl1DcNUD/tarqqeKa8tGn8mcshs2QGpr
57dnLbUOeOGYyeemp7aFaj/nH9q2kmylB+XD4CnDC9YfvfR5Cd6qQOKwvJlVdV7D
DKZK0Ya3bAhDjlvEbYvOPUhtbYb1tnsolwyPSHfuk19+PA+7A4jiwlajqy2MMxO2
/cIDK+evZcSBSNNpelhoO1tuBdKB0CWJSPqRi1BT2aJ2eR/pkbbAfyhGKwsNrYDP
afBFSHa9JacMzGuv8QXzKm4k9/po8fP+kfGsvpLl87QCseVG+wRhHSUoa8NHdhw8
bMmOOGkMlCmEoFJ6kq3ONcgR5p+j+1vIvjOQ3Su40P5vZXV7F5guh3UyLPhfS5lE
gToOftcxTMjthqfF5oWPStCE0zMD8otQFRui3d6ZRNjWKqjTf7DN3M4PSIQb+mnx
RJoXoxuzqG6I078T8KPFyzqAqE5YiSMukK3LR3wjvlf7eFwDmheZqEpxmzGuG1M8
q0rT7K93wX5OlDmlZLGnQvHG2L/BEterD9vCLHcXZ64jLD6xBloFJExHTHtt5Rjl
VHNHjHYGPaqzPZ38L9Vvnv/xc3c8twXiOvXLJdBEJCTBoA46G89aMyrJEhymhyQ2
qrpH+j3pTs3EojdHqinEp28lxymY0gzp13ZgUxTYJfhsT8rrgvx74OH8M0ColHpT
cpukWJ55u9EwJ9c6R1VM6pLFmNFos15BygDO0jt3UaQoJSUmIgbeFyOItlIbjBhu
88ra1ePaS4/PmzI3uMCAdO1yZRFE8jAa1ywVriJUlcDUwLoKdSUymCEGlpv0ojI1
fLe4CP49x20EJXmZZI6Bbq2ztNJrsbbvzwxXVQlE+S/9ZwnEMcUpLYAF2ImvKbRl
BBec5MR4SbQqhD/uWEjeQlZnWWpG5UTVAoq7ycmIyrpN1xpjbeVcfhVbaPwT1BSw
2QdFwm+ryjZDYTPVtQ7EC0jj46EtXIpemlx1IaZJZQrfoqvdetPCcXHXfyEVYLYx
OYa4u1CD2j/VXss01x4zNxarFwSj6T/zZQ572P40jKcV0rLHPZHEDk66oEquHV2+
Q0MndU/YdIhDAp/pY4vFZvIjb2oTgZsXijhQZoh2ZWJ7R4kSPpejVS7OjgRgOomX
q6DfMase5qr9hI/r6rBdbY+tHdlCmoaWj2A7XYaqOy2xGzIC+ZEsz21cLi0sxuaf
LOf/j17pdBqfhCwHHHth4/TkCXCxcEMg/VfGCHGCEUXrlty1JnQrAqCGFCMok2YD
XCyHoWL8IuMlJewk87XmxR2lWLJjYVvvlSbDixOL4ZbWjmTJCoK2UTL3zop3NL5g
28GGHoyiip+xuQDImuHiicsymlQvBlc1neoCgcC3rhF5LLtwLoUfCZ23K63uCU/m
VpLZjdeiDqy+zS2YtcXvl0gKl92naNcpy4JE+ho+VJ/h3gFccIEZIptklcMe1QJ+
59WRhoWV07NS5KLMCnLXQfi0IRrr/UFqSeaWjLJZ4pJAoBRZDjWpD5JTasl0y7Ke
iOxplNUce8VkeIP/uY0wyeJVkkZk+i3nE06V71Rm4bt0hldSlV+RjWBptSKeVUjy
/6B5SyHLQyUlbhwhj70fSQj0W//WXRrEWqw2ePC3Y1gXsqbOC0lgXXCkJ3R3EtxM
7LCoRQVKu8VjmNYk3QK/VkydYWYEPSSPiV7ZhfXyo1XyYiW/4XQx3wxF0yKJy+Mu
Wk00T9iGyv52f5j4K8dNpEGnSFeuJc0mh3YtTGlkStoZi0Wq5ONGnAHBVF6ta4sV
B0u1s6UsoWAEdBo7m7Dx5YIjY2Z7NgTBBezBLA5SDqm+1Lh8Dbr5xXpxtckIK9nA
GvtP93Mcp5DkzsvG3ZnE91O4Tof3yDvUB+z6C6x9omaVuBfbwAQ5KQIlhzsWHnVr
rS0o92YZ6MlqHlF8Tw7rMK4VNmw+Vj4T9WbcQNOzDqTD+9Q1QPb/bdxOU9qorOpK
hl2i4u6t3kylaeSiV/ERL6mnhakJ0OrlPI1vgSJ4kwfEz0sbzybgK4Jog/FrOHOh
gr5VNaNnqLIpTglsC1TeSR9ddJu8eyJE0g+16k06c8ob3J+RzPo0NR5u7gGbEA3+
q8V9OD9jGSZ79zfZOoaz63nzAH7o/txbc+GrrVrqkgMjc+AWjEWcZP3oKBzk8Iir
Vw6pZrHc7aQt2vZCptwVmp3rCrjig27Vc5V8cKb3GWmJRiIZV4EBQEO2vDAZzPb6
buHSNqVHlBiErMrP+3HAymSpSJTbyZlIL6pIGDKzoaSZe6qXjuxceOfY0GwcTjZu
qGVfqYy7vYvMV83o3YPZxQawHpRvPyjRmSeVbrtX2+8+pAihcXF0zJTEX4Rp71xW
BXwhh+BmIop9qO5jvcRS4nog/nUXcbJFuea70dl5beI6JubAjte+4ZN7VmgvbINk
J9Xg+kMpv/oMYfMJEoPppi8Arc9WncKMtIFVSWsDVPnCKYBo3AsgEmQSnT5TcoNw
akL/kLn6MIHIP493Du/G0BPhpUtm56I2fhkE5cw4hcLyACOGIJxJgnDT+W6IYxRk
pGtrnCJgVsaHyYQoqeqQRCnN4V1v/jWI7YkaCPQpx0Bsz7bNYPppkA+TSJs1xh/6
cFDYcr2fJGY5wEe2IDnzYAU3zSwoOQzs+ONLDBjWknABISxH6Icls0kt6vqxEnIy
ayAm5jk7hu9VqN8u1pj0JnXXAMjX3or6v3WX4y4jVwJv1HlkvmRAvS7Bo8DseOrR
sp9/H4P3cL4PuGl/31efnxA3suyULbVOEp2m4MTU7DRTO7aYrx8c6woR3MD6slMu
E2bVvJpdcnR8XzShvye7qqhNbUa5X3DeFJknTmrX7517zDjqcNFJHpu9eeYSZWi9
STCm0iq29uC+C3sMM+F1iOKqzdqocsq7DFJcFydbUuRjnflbXOnbGS4nAIKp+H8h
kTOHB6YlPhXM3AFQT+7bb34poB62qYBNSNr+iaFZTGZZN1bMp1KVjx50ci+oytAe
/8MJ8PAL07I+TGl6pTxICdcKX6LRRgO/4Lm55mRHeyC72y9XpvRlJDaMEp2OUkLd
cfd9E78+u+QXQgP41nCIMQnk9rIiUeKcp0746OqBaxUsO7gpeEg315Z1vW5btaXx
bMcGZ8MeAW2JmjOiPoSbh+YFhJHMFvV9Hu8CVKj8U34KXAQTtAD5lDr65+Wf2hly
zzBb/iLvogULvOke8ymB960phzOjMtTex0k8AuWgWv8excfhlu+DbH5L04Zg6Mgp
G+NsyfeEwsnz13xxFEnrwK3lli5cejhLU8Yo+uNWRRk81UMg2/BTbTQRkPHML79G
009ihEExvjn1511q+qHaahWau3NLIciimvNwf8KioVLP5vaJ52tQvZ2WG7q9GByF
Arry6LL+KOWdQEtQztC7dIjqHTuXwXpkNTNKfrccIiy3qk3+SsaIWPy8P5UXDdbM
XWYLSsbTOpwv85IqsrotREAtca7pwYiQxZGAKWMUfXtrmm1xsURXVMzWIwZRbATO
C2NkS2eHku1LeExgyBWOMzZhGKXcvLQFZ8Eljk0Nj1MFpEgWb1j3NQOvg/y5+JhY
uRquUY+rq6a6QZdfB0pJwKZLUrj/w5ykFbrn713ZKi0KXi8mYxsQRwdnaiPZByIt
ayuE6kKzTe/WGYPdXhLuaiJCLnXRehakLwyt40UbuDMsrWdZCHp7HB3xolDOXsDN
Z0ilA/cPKX91HxYylvyLkkNl8FRm2zARBm3vsaK0c7ncV9zBhbv/wYdJqkbW9udv
sj1WT3NYWCFSrD1ftbFbCTX26OCTAI2Q3r3USHEuA42/H25MvgKE6wfHVOYjmkg7
OocaHi0hPL1SJCoEaB2qukx/Ivwu3jafLvBggQPFqQpeRbiyOs5cj2XGbp5Ud8gl
B0jaOmLX+QI2GROSNiSaV0m1s063YOj2oZuS9b/9oH1eZCZOJTH301oZn8KydDG6
R4K2W11YKYc6mdsQ2PYilQO92hzUTTFuap21iXeBXyvWFVMolgE/U9i8AmkG82U/
42yKwFpx4FMHQog+sscmuqmXN4Z7yggGh48RlSTTRoeTmL3BhTluPTGeeYq94580
SVMM+STKsOAVRkEdl8qa6YQzLqnN/WX/LTPUaID8DWUJB0qtnu4sOfbDqHMPmUbV
C5KGotIIDZysSlqQ4iaIKtYGbhCXtP2j9vVcbrzgs4+FyiGB99rM0oNay80kjUNd
LkY6mbpTvbUHL2keaoAZ4W2T6TfTSP4fZVyoR/7trowgcJZgAXN4MnpYWAB7tj4c
SRfjouoo15PNpMxjuzlpYMaJUQHNKVqY/rEsU3TYTnoFNe90tguHhOpAZ0TDROPz
qpdpi0Za7TZwTK1BDPxQdoF5JmmlbhgGPlYOE+icBGt++reNMqr2pjbYVkQSFF1r
DlB9qole6f/1FBsBPjEkn1EFPjZrWpIEg93EQC9UNr0SvS+TMlJQAg8ZmJoFrub9
NJ/rRk/Rd5akuJD14YbBqdBl1A2TcO2kz1HY++dIPQz99lwKimowY+Bq1StlxEie
xAsgCPXFVqux3CB6Xor8heJqBu/wLmghzreZklYbyfv7MqnZzVIn708brpUF+Rls
iSPzdBJE08hhCJ+W7L6f6NhgBFDBNlVcmiFcBcsHDS/MzDUmuiHQUE5FlnUs6GRX
VyEXWiFMCvo/JHzOv/NsZuEaYCkWYGZk4EgpCMJsNvIxzGRvUxan9PS1s/VfJ1OI
Sp5DQIkcNrfYD++za3Qm7Z7TYEDbePyShfNtftjlrvv9ieCTgQFRUY6bghQ0Uw33
HGJ3zSTbV1nZs05wq13+P7Et/JPstMYu9BtMnYGq6sDYLVlf1BmEOsnH+G/qbBt0
i36L+87GzEQu6k9D6hdlbORz+B0tbqKDjwcXqImL45dcUzEOqgtvXWfshJC73erh
tuhdU+fdPEX/AMsoQGVNR7030dfyBDtfpepBd4pFTtc7LV+S5YBEkz8gAe8sny8V
J59dw/641GSDZj8UlAuUCeKt64le7KqQ22QQKmQ0LAL6cH0pqzztohb7ch/YZzxQ
H28hF31Hj14itob3oI53GWmj6A5uvWiEEEFzUyFvncYjH1uCaz5hcFulv5PCzgPP
VDYJuGssbRHZijxKvoC/p2Zeze6inxleQy3z1A2DBJjuq9ngXSLC9yGQWKZyG5Bx
8aeJxCuM0Ro1liK82U0zP80U/v2ZD1JSrKM0fl6bnKZPbCIly/qlVexV7Z37GHDj
ygCVa7A7+K/89DsFFczDdwS2APoVj6pcAvTU3/IpNJoesFFiml/3YqNq3Y/fxHFt
E357RDpcaZMjooM5/FwsUGlnxgJcd3hrer7V/sQ8QeIYB2mzPo+6HtBbkmpR03dn
fPR9G5Eza7pjhAahQh54dhXXNUr8H6Cb+Fw9SREDa/PSK/aLd1dS5IWB1bQnkGu2
n8TjdgPgXS5PXEzw51VLA+7oI6n+vMUnh2kONQjouRCeDMk1EJWxqpHyB00wb5si
g0Q0PZifOZnT9vaM+b+cKVa87pDmowhD6Ld8PEi2mXlnxSQlsldNWuOq45gGlloS
UzcKByFYOEAyQxMRSKAQZOEQMq7dmtnYpbmHoVjY1qaX9A0ErXkynYnvDZRi5V6s
YXaKZdrWzDVMd2ehlIFCr5UmaSBkfcGyaFzxLCSQbHvdJwbjeNhL8ZkLTIwlnqIY
W0ms3bMxuGVD1Yu92KGJllKCPlQKDDRL6svBYLMRTQlKZIM/vIb6ToqB0tpYQoCC
KbzN6I9Z0yW0DhkYQQ4nscItcRQ6ftIlLt+Ct0tstva3P9D4Gkw9+hQQcHwnsy72
eEncxzA6CFxNgPv+9jqIErHZOr+l/QYFGson2zNq4mo44Bdh8B65WA06hcoXrtYw
KfCwLf3tlgSh5Klf89Q3yiBPhB9uEotLK3v3UArxof1mld03xuwBCA+XgNmBv2WR
ROGW6/jFOzHaaDnpwzHyXPBpHrOFPkk1LxgUBmJ6XnOHkLLK7+Kn++4LFJAy7Fvm
rSLqP+XuXvk/dpaqTnXNJEO6s8PK2Fk7QmW4Nh4Hg3lxR3wTtcMHcyF+lRv37ayz
22bom9HZKCx8uDazFXtnQN6AWuM7gUN1Qs0YpjArfTx5CbSh9OUiKQ49YM9+mAwI
JmHXMtXlHhd226pIg52wBx/dDu8E7pXEJClXOj8oIFMluPCiiCKqzCVEEBbYW+GS
P0bP/zgoQMGU049SOpXu25MCjGbMSeJdPhEPtV/qHSy+JV8sWaA4aAkDdk2KVHd6
tRgApzCGEL4wRTsUnPrTw88kufnJJWKK9sq3QTTrHlyE4ITcu75QqtAJvz+B/kv6
MS/kIMIOgJVOAGWpBNPR8uqmGnAkxK41lCnCvd+fCN7pVVOUnuOHZc/KELC0rvjQ
57sVtLa42WDs11Ps4Vqhhc01kaY2ft71ZnUID2uVZlE0cdyCxR28VufqiJBi9EQH
CpCsh9nZUjYFfCxd2gFIlTstmQqAZJ4CGVDbuLz3a0mv+6jwwPW7Q7fB43F5ucWw
od8x4lf1zqV0Z5P4iMFX0mRwaX8A32lP+dh7nr4gdwrQ1B6uBlzwJ/IwGmkdQHwk
sFbidOgxHUzltQH4ljLtJyLkx6TmwttmQ6uAmqDl2v2v0AiXIKU/JujP+kSXMG/S
6YUAihdxsZeRxCvnu0nfe7tAQchoVGfmmePsCc8f7fn5KRwmk8YZ2AmttavkozLL
czsKweC88BtRZQL4cm+j5fveSBgMdHUsBAhzeAgoz22P9JOAQYKgP4IhJuofxQuL
La++2v1Ai1mK5ipp8orkoE/8tO+GLMfqdrcZrjdC8nt62VC6jESGqvVNkj6adcSH
e17JZfLUjNaDtnMd9XZdxp6PWIwUNF0/+t8XtWAYj3n9DwzfFK4yUfBSkOegDH52
R0MvJzMtnQHPuCTjPVm345aczyxhAN/Gpe5qiby9cI5Q59gNaiTTmMlGiS7gxa3h
8roNrOBwYePHzve9vCW9JqFVeBCnfunwd3yi4E3R/qGymJuronGnl3TDNA945KHr
B0ZOoTFNaQ3URzZepxdeF5aKO2PBA4qOa58q1XFzYMuAZSOwxtYm4k7TjPtIBqyJ
5Ra7rhojA5wZtfdsanBH8aliVpcwnuTf+DAVMbuGYK59TlHAUX3hxoC9folgSpNV
xaVpX7knANtOLauUH4kEfJz9D3vUCXHsvC5i71c0Z3sNcBohMLSA3FEzBXpv3z1l
F+OSTlBTMAZ9IjH0cDPBn22ppdoCksQtzd4a62JWHNvsphCQVFh+M6hcnc5elZDi
f31tSyQqrTR7KARCfb1Hr1Xs+i9NswSuMG6h5AJ9ot/sH0jMWcGY0CMdDOAVEVg+
rfCM1S/daGRiMHmtpeCcBXIIDnrCi1i/CPxNLaMlqVdthapFzA0agrTk4SVz1MrN
iUoRe4BlD0A2V98q4BVGKM5EhtgMborXR6z+ntutoq+FsYOYtm9hd5nIf1W+Zcte
ZBn05P9PuBTpkKWyjSaG5KWb5PuRPlf76QY2lQagxaZ1H+Ystrg5z3Cp4Q8b91TE
Bax8Sufjkr7u3SrHVpDJJUv53VchaIh61l0GikHbKCDvNdK8WvAw0J4ZjxNBgg2+
VKBLycX053ZUjMJQHGgtFHhrfn/9ZrlpfTxVPHm45k/4tKMEyvepkUb4uUgHor1/
Q01IiKHCL/6rNhpQy5OYzsAahh1hjy5Bkql3i21xCIE0jn0YD1nGtO7GF+rQLKXP
pWKTS6xSZZ9s9KxgazXD1t2f/wXoKItupopREiCO9t7O3Rf+m1bRo+vyRcfKVpdp
UI49TK8MmCJXbyILKW+gYCYNikp1PW2lHKEPcgXfrDkzfb+CROp6iXQ19JB1GrJ6
T4yiE0P/1cwlCynQK9M1SPF6O+KB+S/dZZR+w2Bc6eB0cF7wngKHMjeSc+N7CRlh
osMoLdF0KWPil+VPhojpXtS5xPLK7aSUThAsWG8kcw3PkcHCwOWYEI3kDbaPX4sb
cW3iVEt8jBN2gqrPWYbvSngsHv4WK3AAaZRUKNXnOGvCSPwQN13Nie2MYcwM/fxf
5lWh5c+B+JeoFd9B01n6u4mEZZky9JlFqFQF/P7x+ks8ljkcDdMNpQRdlAcFFa1A
4WJyAOVt1QAtyVo1BHxq9EdoOLL6G1KMjH5lCuCZGlgbVrvw30t53rByCRCHE2c9
0lKD2VVLkl/gaReTUtEEGZcAoiOdgviswbFGxjqEc5PPLIL7CXZByINiOcibv7KC
mT25BePWBSZEmcqHSvZkFQj/c4b/+ai7Bm++SIJTCnOARa+8AxDgkfYDCxKVKvE4
wDC+MK2kVEQn+cO/M+EM0ZlEJaSVsXo9MD5PqtlZHe8wvpC3RdLtcV3BHyI73DYu
KoHShppA1FTEWAQhlMDzGPfNSWiqWQWMTEXou9kQ9uEPAApRm30DrvgA5g+TO8c9
i92myZORqam55QPYPF8loCTNDFJr3a1GlP5vXjcEyRO8sW3iM5hTfJB/KbhPQEG7
f60byCLdNZKeHHpHLeJrTNQUbOSAQyunpaixr4qsn095gtkyiSFOklur8OKKFMJy
yVqJ99AyJkP1/ceH+4N6KlwvS7b6aqCU/Orev3JgWiVk4ms7YcddEdZR+IXoODB0
vqrI9t5OvsV/I6NPT8N5psdO6yduc0IRAQ+dI1mxG4zhQxIYLEetgaw7O530Hbie
tD40FFgyHOswtK3Pc5+HSP0V/OXnSiesDP3P3Qre8OYZMjJDiErCMDL5YE+dwFqJ
kW4XSmxa6NenSJxsU3Z9FM3ds8w5MKAPSYxn3/lPG7Ys0yTpZuMcZYVgN+imQadT
CNTZU1ssEy2MYDiXc4cInH6JDpCc9iAZV6RctnQ146GfvwB9a6oeQ0d3lciitI73
nItrQAY9fjWLhV9lfBKvoeYXFs9aX7rMpeG0CwlDdvo+Bz77FQ6l4UuX9L6JiDB2
P4VUAD52ysp9/mPQwW7PF4OqrS9agAif/Zevo+Wgz/3IaW+HimB8SPAx1CCWj68N
r0lcRtKxpa7ewK6AwCV5ysOxQ2hg3Oi0Lum9OWz5vIiqvhfaMyjvYvjqrw69Iocf
gOUgq9mrqwMfT0Lyu1uiUwSsjduad8NNJIJxwE8P4H2CdO0DneA0FNqQVmIVtMjd
k9m/mCpb1XenmyG1G+hDl8jM+G9aO3XLrw5vVa07cprgaboMOzm0NgHVqjJHN3uS
u6Dpb1UzTPmylTeTMH4Mp1dRgOTDLfUDcxQCx/pCLxiCzY6MoMQgX3SZtFZ4kKFB
EY3y3nlRByGBHpKuk4rCHaawvmPg4dlIR16UzSBsMdom6VoAp3nbMhRaAb6AyhA+
5d0fYURYDKY6HYDm+a7DQavt8BqTzeXUda/HCS/Ru43y2w5yQeoCfoCeSdBTcGpv
h7JF4Fc9ZPKS7P31sIpF4qcexrjQRSfMKhIKxDIRwQ47q4h+eE7vUpcJWvyVTPiq
nrJj4MDT6brFimUTJ4v4XLqZB1UTtMZOiub56C/L1KTj9adez4ek35bHldEgKLHH
mZeZwtJ92vBzwfO/48os1ZEz6NPHOh5VYLqhWUIISgbdvvExR185ZrvuYWiDDhBO
MUTYcMc2iqWxDUMrc35yq56EOqCMXL4kjq/GAXlKArqB3dbNVmH8v1DAin5qv4Jl
ETUynsAKYCn6Q0jpBSUXXp0BhPFQobtTHSL1G8BB9rloYFre83Dz0GkSdiAPkrx3
kKbwKqAg3sjqVJdvlyufY/hMhGHuCwbQlXEHA18nE7rYSI8WkFZek2QnHsrhOKdq
G2b9HzbePH1wVbxo1JRD6TdZKc9mDSYPyV9dTc8T33M/+rYfp1gk5Vr/Z5bCi5Jl
x7j0t9kB3a/y4LaT5e0OSWaLS7wppOqOpihyBHvYf+1HRIvDBwbbCQhpq6A/VxAW
Csu1CjccMlGVynUoMY7gv7mUMeextRJVoHRxmd212oCvhIBHHUyie1v68zM4ZEit
1AESSMtcYfS4Q2MBty7NjsVK1n3RQI4RhoQJn42cHdcBfTcVz+1aAsQ8zOTdV0FS
KyMjz44YyeKr/S2yQnmq/2x7BxnSbBETW9vHvNSgkaxt75qs6RfLu3cmTSD/ajOh
UPqkjZhHy4zSWWtphp1UJEDpXqbeoncJglVa52Ucvq0J0M2U1kAflprjyneT1cFf
WiPg1t9NDVnwIWnMrL/vILVzXkzfMeJn+otLyn1/eegQ5xY35intg8bfoYxZO7MQ
eE7vKFF3stWTl6q2wkXi/DgkDmgJBc1HKyrVjKWvLzS/7rTkKztA+H3LgAr0gTn8
uZwOdGn6SK03AsR3hs6K6jUAngFnT8oBbtV7m2II/Vie8HZiMS8CUzYWRWn80lIv
fExYTQQ4jZDxmL/beXm2tyzuhJNYWUwL7TCtOyXJwo9UfqUcb21t/IAtBY3y2+Rt
l/t0dDLi8v2Olc1TnsAM7DV3g2rV9RwVhLqFDNGMhCBL3lYzVrABgcxoYXXT1XpR
CWp3Ka/Axj0j8E4/UtULA2M9+I3NRQ6Cm3fZj8EMVM7d0qmsfuka5ET7y6cBUKG9
y6mZl2Ub9h6oVKiWVkSBmcdVQPq2VnnhydA0YIx013N3B5BhuF75RMjxWisLytnI
JDQdLWIDBKdlswW5bsoh7gFIVziNAPVD6M+t3nZVQ6ousUslQNUGEgxffsX2AaIQ
ax0+UcPep+RLR72jKbCRyNwj5nPgbFU7JFe+QgHuwgUuIZQq2xbLVMACfRz9uvaj
q11sCoNHLM/1DuNPtW1F18nQiwOrNTHtBJhwxM1fwlf22/jEVr0+ZhJNzMbslmwO
824HYwv6gbuJsWqT8+7qwOBOzcK41xzwBHRWslxeqxuUJIHBVFcSZOB5v+t6NeFe
qIB23yOkgXB+C8xSZxnpj0kdABFYHOTD71U5OCmJqsz/Wve8U6mrH4fAQom6G6Vk
WtEuzU/nXLBYb8GrFmHuR4iiVB4NfokrMMFhXcZhoV2LfwbpPrx9Y9H3EBQ7S3Q3
3aEFT9UICZFI050Y3xqdBsO5crahOM6Ox6xBrmaDg5W5pAcrRtu2RxWd6i9YAPYa
exc5RfwIAVhrrPKbgZyWVs5YqfpizTPY164Twwd5lvbYjSLZzmxrC5bg3x8jnZKB
4KQy+2Ng2WU5rSIqI1YRkTsSXy6Mxr0UveWmCCitCqsPILDAEVv01KnjRcngTjUu
JS0CDuVFEsAbfgfWhNImDxSeahVrHqPy8stYM7aRsB20xMRzVZ83vXNjX+NMdpcC
Mmi5B2YsFgKmuXn95Fx22rhxU6z3O0pbGUng6tUIKxnxNZhXHfliICT0zJbzLpIC
Z/eIgAOC8d/kVHzc4f+7tJGW4JP/k1k4syCetd+qikCysCPHqgJAZsmb4WYYqk3Z
IffJRVTNV+iDtKwO72RB/OwYwTsjUIuBFr6s9fUPWDoRuO7sWXJIvwyKJHLj7qjx
5OlKlDv/5oYclHpNaOIwtI9PwMn5RnPgvtvsH0/Q8AKd5Sl1eAvnGR7cutuvHl8F
mBOQosE8Gzx+5MFC+u+3q59M3N/88xzUXBVIGqGK37Bn9IV8PKFwRhTBYRWwbBpd
/jQubCxPoB4WEN1MqZfhSUb+3Y16ieNXUcJgwzf+PZxfgKdT65r782CUlqPMt6yx
7xKbCRwF+jmsiRt+Qs7BfiI155I7CUJ+knCPQfEmogpizPw1BdxFaP8gKiV/5sZE
VdcoSjie6KWGvgwLbuKWcQR05MRWK8IlvAD41VSPWXTomNO4C2DS85cPoI//YFEh
7bZi2tLXKGfaWTRJ5G+CyMRLGKZ4IGs6a10s3KvCOW4tkq3OSmV/fFGeoE252zA4
8KiniqUPyCRYy0oQKo/cQ1YQ23w+8Njwiiqgo49V+gABe/5HQMbaqe+6KOVmLO71
hrud01DhTW+FRphmHqGqM8ecPgMgxX5CIIAz8MKgpiNXCxpESKtDTBW5kpyK6Szr
dAuclgh4RHI4Z6V3ZfcrL+XjpnLmjYCSOjQ4tpNpqlYjacpkHM+Ztm+vGr0Cfise
DekOPsLvuV6k2zbp6BSyTY0MqfeOAF9aaiHhfFt3msrM5Bz62b0hSQO4WPDmyYy0
OFGXsrqwv82CvXHnjn2lDMi0A93c6crImVhrVt0AA/wqdD+cwz9nMsifyiAD70w4
3aDIt/5mCbKSbs2ppQJQnb1rc2SaXzhmEAo3EFbOy3OvNoPr88bQPyKB3G0v2rMV
4GdjmAbgmcq85xp8TOyqf0JKemPI42uI4tLwaaUEu2akEcA2tVf3eR34BC6ySst9
PNfQzyU+oTH5/wq/fXyggE3cC9zKl62DKm2xE9aGcFD6PhTINyMVZaKEYBRwQymT
tMb4EzJOJGwCl11BL9Hbjns8n6UyAKa7KxnNFP8Zc+29n9idWtQ7zKHUU6wT8TK0
HaJzgJihsKxTNz6XhOdN64E0LvRCqkDAIypdlCi0rb9u3IghSgzheNMBt6/3dJj1
nuAgYfASLfC8S33BRPCgOvyWoIZ0NXMD7vv2nFYrYBtuK5KbZ4IgRFXRMEX9DeZJ
5yJKr6q2RX2FEDjud3pgTlwv4G986J3TWapGehknYamByL4dnN7/ywgIP2FjArBG
W3c+I0QqsHXNbOdM/2XZdJ63BlQuNd8znS3GG19WVEwiF+j27WXLcCnN3rCwz5Tb
jtqSV8DUsAeWh4ODu7hxszonE1VW0zuWh4K1paRp0e9aS16toqWvlkWHUz5hpgqt
4wyIY+OafcDSuwXx2ZUXQRBe+dZ9x3pU4Qz6/h2aVoBszl8GvjU1BivBAAhDr2If
FMGZKgGAHLfzxZCgSk3vBeiXsrxhQYgaPV8x8J1zQppf+data5kQ1q1q/argeiww
qXJuXYf4tZNk181+XM1eLGUnMbKBWP+v+js3KMIHnVzWJjUwyZ2ZRlfUJQWVzgT4
Gtzs458KNv6FN77A4bVSULc4aizQePrGm+vKkhN7A3goMzi5H5TYMzhHG2f9aJz+
FKt2fkTzqsIhy6HgCl86SCLlRJvT0ukO1TROqfIfupwQVKVDoHJNJOlzVYDYtWz6
a/K6I7dhTKIKEyhgddk4bByIJQd3hCEigtodYZybmYuPXzodv1BQelPfHws4LWAA
Iz0e8xdVO54gpFDGCPZRB4pOW0gCJbsbtsfNs3Rmc8jLngToNrN/DHDf0l3t8TbD
GRFkpYzuDYWLgSylQ31S3XE0penTYxqIz0ClqRBvk7OPMoQhwZZRp4WnE9nzw5uy
RcGeSDQKuCweo1ISEoH56ar1JsBXMNvaa7U1sC+fMhqYzm9ZH+oP3VXTMGVO97iN
vW5swSlNg4T9w8NrkMiKjsWgA0MOwIxdz/U/2oPvPqhn8UbMqRDCxF8FdRvn6Bj6
WXor+9/8Vl8xpGsHTtCouRIro4rmWJYL0Gaebg8JA6U2rU4Ki1kJP4KBsa8gIyZj
1Z4oKLsB3L4GcmKLe3flrJptrxTHmyEJ1dhp+VpM2vsinDAsEUAx9d+EH5TFtH1O
nu8qU51uQ+Z3v6elnarSU97ziX/cwLtyjntp+qCt6a7kMS4G2ykJ0pIRyVWcSTBd
Uo1coq/Ae8rUaMDDgQK2cpbxosd+090rZZC7KcdVy41qQRYB1oa0yLtLqWbKVGZY
nfNFr3UYY+eOHtjzIyK2sohQBbxQbXCQ6gd6nze1fBlKxSpk0cF+VxznRM+/8pxx
DKHJ8LTI6p/epT3xahFheUSnkIO8Fkg/X/DQD4tx+J9Ki7bKhCHOsw4llBq7DRrK
IG3x5aQtIM65rQ09zXXJMc/eL32KA4IeQl4YV07/ZquxBxw6RERzq275/JZoFwe8
qiV/CI0QstCzCK+z2Gku/De5k7mZK8St2lAxCX6qd4c9EboC/HMsAj9wmhhVKGFi
tdE6ncC4CuT8k0lIpF5paPKrHCU6aKqAJ60DKs2Fg9Uv2/mM68wM+bfT1/VJ67yo
TlJnwoJ/nqzqefaH88JtbXquXALgjFlxFuX0ZZ7Trk7fu1fmluoVKVlweIP3Nbwy
n/pXMNGJSTlu5I+3GGmJdzWIfz9Ry/P+xH65zNMwMofZ2U3+QXPhOhfe/Z+BAONm
okzCNFBwDZTxBK3SnZx5r7shKwn2nGDa5G4bA6zsx6LSufpl1ukugPJ9Tg02RK7o
2v31S61SKQ0AdqUT/rVMg4pOZ1IPsBMlpsrS2Qy7L8JwZOscDmOV2X3DyHTZhZPu
jK5aNCS3Mf6KpzCMp4rlA5kpguAmrop9FsSIvlZtAyriUQjpxdUyXv2nJY4Xjmk4
9w18Xlac48jYIAVAo1H3HztHgIqAYDc3yaKiu3fPraIctLcPbxkINXolhEu/Kijg
847S1UVhAJmavmjbi4UBFEd9zCkWouj/Zi/N+9cB1OfgIzqq3cusA6/aamZwO9vP
FYTYFUxR575bd+5au1DkOxpgzWtcw77ztj3d/Twk0KtMXzAHsRC4414lKqJW7I2D
pE8awlEAPXxrIJ/Qvn4ewpw7ziR2V+Zvk+Qp5aRLQ9ero8KbuxXWgj2eDQyTN7v/
yLyZLEI+se+0KjbQxQ7kKY6P73uU+kHKhXS5YBkhp+bLduVNcsoaIWjwlMZwInih
sLwL+vEfdWoOckSOv8ehmiylTF3lkBa9c2Nji0ShUsQt3+A24pARzpEUgeEU2mRm
elyxjeGHHIec3xXn6wG0skjn+y1sFzD7iSg7824e4uRvPJCDQ5mDcXtq9DEu+CaH
vxcBBWjalIrdNfcnWE4bYJ7u01PskM7z8vNkF+xbSTVhvMAN+H6Q1gMifMIUPFPo
6e/WNH0ErY3koFsYFJ3mDXkvGD5aNEC4THGY5YIEWSCkAUu6/KBg9SHOqCkCkwnl
7/tamPI8+cmmsWv3prEgtNHLldJWxeZ2hBbgAUfqiG23hpS326njSWzCyvCJY7ld
my7IMj3JGlD7kjn9LRYm5iw41de4REQJmKOgSZ7BqmKFhJOg487dtc/ybnq/9gek
J9vZ/rhVpVQOhiDRMMRnzQX+p/rhm2BQ/RBJwPfRVLB2tose/ZH2glSOzK74pg54
5CDL28shtjGep01lwc3Aw9+QZ7uAUOQeDwK/twfBtTogJrUbaasYoRQVcj32N27K
XN6nC3LskYtKWpyauMxcZGpDkDvSK/HYs8KDVK6VHKc57HRwYvB3uWZRVJF3Kpz4
IJRbx/Mph6pS5Ilu2IUYwhswLh3EkS87FDKTWKGBVtpGeDTVQp1IPk1I4xp4DXZk
0yhKS+mzcRxObbm+b61c+obYVDJDUvSTMxJxV1oNX4oCy34FHr4s47XCeDHOzfzc
HiN5ETkJ6SdidKaVsWQnHv7XVihtFBeaRt62wvXq/MNk462Uoz2Hhu2BSnl8HTzY
79+dbg3LqxbFNgXACh5BK+youFCAtWFbFYxwMJfavWP4LtOK5K4FKJvzyqON/6t6
PSsA/mt+2aDufAwjlUjCZemgcNk/I/l/8FwvM2koSHIlOayInJPedYKCjbmLGwF2
oinPJrT4wLXLdbu3zORoMEjgbJ6Hql8bqbDLYp+EC/UKgjrniOCfaHDigXCLAkj3
EZo7GzU/LVvsmlAmQpm2etjLoDltlI+Py3hvhut2Q5m1gK/JWledazWgc15hWWXV
QEdUbEg3Zz7o8llsTdzTqNrBkwEFhx70+lvkFGkM9ETEWkGjZ6Y61/VSI/JBRcxS
E4w3HMe2omVTe3LsPBou3Iqc8LldGXG3Q/qHgE9GtLsedhp4SLmuLtMu3Gofafsw
kU+IukbO0BagLgnWTBiPgUPkOPbWtAz4f5ZqTxzC5BIC6hPF3vMt+JW1R07MJvvV
phNrDJE8IE5cAA5I9OLkNr4P8ovV8OHNWRyLt9FDgytTDn5FKIeCB+3cmWo/e3a4
tXK4eXh6BtxmiO5tV2QzSdaI9L+/MXGO9emWZUxOImvoSv5Xf6TyaXZvdi19s9az
CGAmZOmUWhbhnqgDQK6GrdcZkvXT2uwWkej4JfmqqLoVnN+IR4E1GzC1+rUNVr4o
jLHrBYEV6pqXcU4i61GxUhq3/w/7w0dDaD3xvVgCxmujSEG+I5imFd3z1lHzdLEU
IKvMErCKp7292YnDHI6vcUYmyJ5g5Ovz80gb6+wgdrkO/H1oxPqDjIwEena3WHj4
htMmNscEq0Y7sMHbXW2quotQeYeAVRF1k5U0cNfl4XE052Qn8OlXuIFqHSJdlRUu
fTW4gw1mHRWEP0o1+ZVMxuPHz8x6Od0XmdSXJXYrwDtWgEhqrnjOHegQtYJN75/b
x1kQw5rosq1JvN0fHKN4O3zZVu8ie34JBkSmI//qecZKI1h9DimqqdSv/OL7xr9j
clyyDQ115ckgMD6RdNCPmvyQOCbpJI+YOj/FUZ3B1XcbMK80H2PbpDJzZz/xqX+f
ajT2maFRsF4CnFsxwj9ZQOIpZyfyLEviKvRGkRffNE3+f7JZBcdCIiyh3A0xmGTi
T5vBrQMhWueJ2N5jIwnx0ZqqFYp/T5Sdaq6Wjl9gYMgymPurHUCcFSumh4PlDRun
Bai1DIw6MbjYEWeHiCv/wZ1JfF/DoZvfHFQ1R9d06lRGtbWhytxZhpYLfPqdXn3U
KTbUnWW+Xme25VAZT0wlykQUwJW/QDQMbXNRV/6Ic8+GFqEXmc5n8xmGiMFSSBHh
eDinK0grb9zZjV+EgQt+eKciVo+16uJNPQ4mWY6IS0+EcSagaXygZ3kFCRxgLI/W
e1msL7+cXzxa5rx+vfRjS6C89fwcVzPe40b7puDVWMP/7f1XsP5OweQatFDX9dMZ
c/nS5kWEgL7Mo9Vi8FBXa8gTefgKVyWTIy2TAm0UHu79NtB8jqXRqaqUPCVcKzft
VgMkUax8RBC8P/WhgLxWoSy1AJLWjmP+C2p8T2zdXob5a59SXwAlwLs+BbvQ6LiE
2mPrfWhEaVfbFzOjgYfT3RmVGjOcUTG+vBG1ZR1j5ue773lr0qo00i1uoMPva1DO
Tyk7pZboWEtiRs3eGtT1T5nc6DLJZ79MrfcSMa3inm/KMJIlOqeOFOiIId+AOter
UuePrgCFYR7/Gn3IOCJ+g10qDEdqzPHv/JfGkCzHtTcpsolqGDcS4DpcLklu/YHp
kKU3p3qotyAGM5V9WqV+IY0OUGGSPYnqrySiDnxOoR544bgrc+v1g5Vq5IYr5UhJ
B6Jh+hdBjzt/dfkDdUFmEfcYvZpYMLOkZL8HKhLYpM8EsmPzKFP5nWel4PId58Ca
zSpuBY0z///ljlUhKDBEOpTLy5/ZEt4rifSB2uYX+R8pFPJGuWyzXfxUQTr+dQYF
pctZcSNUTV5CvqcyEdo0yvuqob2RwCnRngN82p2sJtrx7b3oXTS379TTcjuJGyvV
5Nqc8ASVI3ynp3c6Q72gmvVxxClWyG25P94Jd/u4U0qR2uF1NnC0Q0zVq1koIgwR
xslNM7HxkDxP/ZOOUITHg+GytujAAMWqM49CDTRo3P1OUTlJbA5xP36a4F3YOvW1
gMJOPBxm0IC4DIt7KwfIOv9njYZI/Hg8VNees2A4CJzlSATHF0/AT7ux6kXJT3ED
XGGkWcn7noxLOYBv/2LMXaDU2kkJnzIceAxkBncwx5sFrXgMnGu93HGAY2DiBh5k
OXSL9BB7TGE/zaw1OdXGcEa1H23KN5OMgHsnihZvI53Bp11EBUoKnTU5Yj1NGp5I
NUsdLSWNb/KYF+7PqxmtqRZ1MbAa++LPAPeCrtFuzmRYbmigLPMPg+tNpJMBxMfr
Nu81W6Cad4HpUUraP/SEq/TYWclDxbpqEK1QW0eFe2Q8SsCHmZR9AhJRgIw1Scdf
Vau8yXykH5XDqd2nuA1FG72Uh2Mq7uHyz2wlRvYCe8yh9KHkmobNn05yDE+GqsCY
K1bUhJ/erB8wOAfsZiCOAQbcJKxlao7DHcbXGp9oDBKkNvDXkugWR8lZeH48svF/
pjkYJFJI9Y7I4FekYtVQSEZTbx4FruVw3hXwJOf+9+2/rfK+rybmYQAo/8qMN4pF
RZYP6s+Cmh9MJryD20GiThMIyPaHlGKP3yEqmCi0XGEOPQnIEuFpPNL0NTBlyrcJ
qFnI44ou/oCZSprWmbBr3CAd4fSeF6ik9ixMGlm7SxqcxyXAIU9pbqadZeSueBVQ
Htsx3EJVbfXtfWGgpoUxMM+pZkueFY3Tvuh9vz68oBhVYAwZNv1ILKO+XFxslHWq
s9Hjg0cNViu4I1ttK1+zzNQ9aS2mLbK3+eXoDOOCc898b8aXTuvCSP98+mL6afQs
ryNULgUaH+eeY9Pd6SJN9EXI7NoZJKZTLufK8CAn9LhPi9waTAgcX30SZAj07cDY
VL6bfPF0dN+5WB8oE7oF7R9FQpsxMsy5hYrMknk2K87i+25UR504XXISILZjmG7T
AemJtsR7HszpsZU3lk+jG4C3f2KNIxdDN+q4Q0ZEqRB51Pxu66ZWwH7Uz9WoK5Gp
6JK3O7LbGvXKhwrT74m/CCnhyaqCBiUdFB04LMblPZ9hMC9FvlJbi7bnOpLdTP0F
teASc8x+wdXpkyZvXIVLn7+1LbcDzaVaxHZn+BohXHGGxM/xMuGrJs0OvGHV2fM3
wSi/hQss3X4OKDdabH10T8zvmgs0YZu+tL+9kZe35fadHE2VbhH81spTA7hcCDs2
jzOMEiUYXivfCc8Lh8VrFV9LWetA9ETayXf3+4tMdKLthT3gifFwOtvCaf2s2/6P
6kkT1G++LGD1v3g94lT2HUpcKhahRfpaw1k4oEQOxbdvP/QvRV0Elf3v7u+86AXR
LOL7IKAuSByI5nnbvUiDx4ZWqa8Z3hH6c1Hb5t94jgfEuqE/UZzhO8MTuPY8MJl5
5M+tbTiOZQDs36EFcSVP34OjaqbtdAbOjhruO21VjGw9uhCPaE+TAoG3g8be3Nn5
lEX4ftjnzxdfxQvnDvryiAI8hNVuowQ7RpMtViTBPF5ZFq3Cc+Nmt6o2qMG0khEp
J256Ft1RjFnp3367D2Vpfzc9PQCSlH3jGomeQHcTOm7Se05NQxAanx2HFj3Q9cZR
q5raKf15mNhWvUmO8oQPkMun4pbrc/W1sjET8+TWugNaHfNgSlsI1Cp1xV0XozSD
LMl9hmqKUToAOkL+/Xkv2uyj6pWNAvcHpIJkApTpav41xeakV7N3QKLraHhZFa9G
bYMaIGxiPHL1ck8ieXf4UpXbXy2YxcSK2OieOerStAHHTzhOLYYd1N4usSjFBXyM
e1WnHX/i1p2nc8kh5bQ3H+fdXz8ItG0tOUYugwU7Bl+U/lqdRDubVONqyvoRefvV
pPicO+eyuFF+dSnNhOLvi5/T70H5CY70I3Y33Q69EWbn3Ydn9uvEn8ekRjGd+32R
srs8ReuFNtnVbDb+Oo7bZNa5HL20zQ3AwQ4/PKcfoJ0/m2U5yu2PFUo/A8dc3ZNw
YubM7b2FZrafw2mQ16TOihG8Zervu5KpmSH2Jd2pkM8HXUuJqUV0DS0bKMZneT7H
Mn76USHxwOv27kJ7yYhTRVRB6eBsOWyOLqmgJAYnPh/R98V4e4mjez7niwPeP+Mu
TZcouQ7cstqGbMdNYt0JZxqkcrxF9layKp5AhuqIf65h6vuoEfembFS4Y5/AD8tE
VK+8Fu91YJETvWFq6n7TogoazVQQ4izdRNXD9ZFlx+oRbyyx84HWhg6G2I4S4WRd
AhY5HWhfwo6cag79/lSyJM9RT8EIAeY3AGiaY4wtWWCYg2PdmOaiNU8ntCnTPDwD
7EHjAjJLAbPgnUGxg8scBERVRxB962jFe/4BGv35f3eZOSHDEdCsoUdWbWLsxAcK
6CwHNK/P6oyc1U0K0OVNpVYVw8xxW8mYK/tURvFya81tKNIanbfjgkzUf2s0xbM6
wS7hwH/31+4Z/jdGb4Ms7/EAMylKn4Zn+86yOtBprtsOrfLj5lLBTjC4OO8ES4Wy
xV5tczpd/T+yOGqbFrm5aO+/5/4/twvcJX8rCOTdpTZ4sZkr5ZSc5rVtvskF1cx0
7bK4X1GgFiGGxH7I1yZxeoJi0i+Leknwrn0BxDi82nVJRH5ySutlH/3/mNk3mmOO
Hm8oEzwtr3NH3lHqn5YXAHecMGMlA3awrhn8anjr8YyaSfQzR/Zyktgp6RoH27Rp
Rg9Jf6GsjBCGOi+je5i9iYV9OqLv3FUhKBCBoKqZjk4Nh8vXJgAkp0ZNZBqljARX
tMilg/yDad5Hki2HxKIOLgs67bJWZq2t+ThviDkj4csF/Pm9XjpRzFS5BUIeuwQg
DNchkAMpHnjrD6rA4aheHqvBzRAR/jvtruraLGWuqWwd1iFnpowRd8pKG+BEx2HF
SFvcahGvd3k3XUQWyqwkfr5latPaj2XncKgBcHT2hTnbx7XTbpW6DuhF9pWWY8IC
g0zmCMdgZpJaaiy+raTIhqJr/LgdCOgJP/XTSZ5iDQkQfrddowmeVRXoGhq9yCSP
iGGXKHXl6HCou5WcygcKamt7Wzys25oy3wOCeDMlW88O/fWjamyyjVVEGsefXG3A
WEaC6DW/U0AKOTm5NYyulbcjapIiZ9dZkvsbA54P5a/MOhAQ17sy2hkFgH6e8DII
VXG7awFK88jihk6x8pnEP0kabwLDhLgbfsnBGEnJuc72+uJ0b2EXsxRChz9lJ9n7
CvHD7JugnSCsF5LJU0eMvm1DBmi1UeacLtOWmoLiIgHYS/uesdzECxx6c7Uvdk5k
HCBY2vv3r6Mq4PAWxCWm4n0M1eELUv9rW5LGWQlnvw1oPSAN9ue8q8OXq1lMGttL
JvgK6c7rVnEtmRIXeeBdHx95iATvGbfFfy3C1pBCPaGjb7Be5e9rDXNB1zUMTYL7
kfMsuJapaiiIVyWxGyRpMriwv5CL7MqUfQWYUUNoucEjO2b+/NsGKwSkNJYUDwiV
RAAlR6Q4GJ2L/XDnka4I1pSNu397F+nI8MdeebzEY9t6Aa8Xwj1VXPoWb+PMrA+o
eCMygw5naCi86MGgn7lSir0AuOi2UED+b+wU6oxJyxyUIvxwZiSuQGiG2WtqEwyH
nj6ysD/Var0dyAdBnpennGGUSNseLy9fKHhxn2LvKkKfP1QsbGYvjpWXqKjOHkDg
xcYmj5/rbjeiGEZ7wEdmQ/bQYc0cQBYVBTLSdhzllGpjvj1QTmWu7wZ7cOQYXwq/
7eHd8ILG9vyqtOxonoyDaevMK1ucqgWunOXnrn3orYy6Rpya7v6EpQG5EMn0bv9C
9nFi0L/5qIQ9/yiJIvkPdjw1dpWE9EIHt+vORuWdNq8Dpg+S2dFeJ5hFHUyQ6nRe
vPrUSkb8uwrpFWvLJh7LdtWTf+kT+X+yHHiiGmI5kBDsJFcOP9xfms46SYNbTnJa
P5mcWG7fG5pdoQ+ybE0AWiXo4AKkk1QMd8qOGhrjzswbjqNeSETtbXBfpQrMZ5Fy
t2EfSGcb6kNOae1jQQnuZyhnNE4XknM2j6JFcOgvo5YmsXiuN6AHzxO3RPrzr5tQ
JTB5BV+osnngzE8QwxIhqdlAegDBEYfmKxb/C+PMc6XcE78bzUdJ5eCYGcpHsaYT
LjoR7YvvKUBYf8LFH6LbcyZ5v5OM5oLuVpbc/8zLn2ZoO+c9JWWGwYWfHhpLQZhK
PRc12gPqX/3/krxfw8Huf0dj59aiy9Kw27eQduTt/JwCcK3covkyPqhgc2ou/+DO
7flq7cqo7zxg55LRtmGHUC0ClDfSmhzLWVCDh/9Zds6xsmpHLhnInxWrCabQeGOJ
PYBPxYotX8RC1UQnk2dAV/CYqLiaj9/XTu1mtotXvRciITsHMM6gEzU6uX3GsuWd
qS7t7Mtw08MgHS8nvyOBgT95aAsuFF/2pXvX2/fxjQa27hl72rIAV9uFIxxXhCHy
6Goz0Z67noaUoagYuQwhAgOkFYuox1It2tW88iN9/uS1WLAyNjElsTis2lOloOgp
LPXfWhAnJhP9tqpkH90ljrM9x1+Yh9pneGmET3iPlj+WHYADxeurRygmdlfKfCLU
yk4HcyvQfmqzAe8J+B0CJcz8nd7w0jEMWkrNjEd0HI4FZIuj9PXMkTr7Q+TpEuEU
kNW/jopA5TLGKP27u2ulaKjASBTxAzbydh4YiKusbuuF9w4wmSO1Hm6Ungn9/0c0
R7d3fUEuqFHWurpJjLrtQ14PBThVVyGPISdzopX8+xtxNtBYMKHA0r+du/AkZVfd
iCcQosokazmAoV4EXetwDZpz/CO3ID/D/V1nSKbDCd987J78Sz9SzE/UtMmXXABl
ERmrh/4BdX6rBcSGhbQ5HiUQNDPDBnuKO5VEpy2drnTJs7jQ05HVBpS9MSu01PP2
EXuWmgs7xntHei9vtu0xDZB0H7/6k7qCfiC6iXnTqXDgBRA1Trsn+mHMC0G0O0Eq
43w6IQiBOc7VCCPVh8eS2UouiVviGdodnNMkJDLKYu07zC2fArZQDjxOgK8RvJpX
aoDEAGIvsb/TzHhIBUUjajG3iN0DBNTrAtzffuz9ykYAo52GypNViJc9nDfPLJea
KoJZvD91MgBqxTyFbn0jdbNk/pTv7ajolvz9SeJOqKvm7/egbPHzy3HyvFmoNspA
XG/nNbib7CzLiOvmS6U1GIc/Lj+RMLGCic3Ek/8b/2uxICN7UCxg1cxXugNP0SJD
uVB2v936jZaCuKA1aZsE/GgZdKOQkAhlrMT/mO2UiRPNCJ+DOvqFDjjR149iv90B
NP+TzxBgmboqbKW3fjCWs7t28oPbvbwKG3GU7obeUIWVhEfpDapMyVxQEUlpU7Kz
um9NbCKTE06Vngm5Pdy5UKod5UWrl08hmVBUjkxPo0TyAZWQJI/qzkYpZBnKvRzG
F+bFW6qgESvWqq9KxMf1jsC+nJSfrMtdZyKyo14gbKEmBceB6KO5EqXj1HbBoFGJ
BKCatobgER+m/XQFsnhl2irryEyQLnzfY1ze1z5rzqRC8p3rqLDDaq33ofxD8bLB
PsjGLPZaJ7jPwitbr+SdTPR/shYnC7oKfEv8Ng7NSIv30fzbaHCBCy51nny6eBdR
ahIPXTXIwf1pV5QMu4nPd14m/4PHHh+fO2pOK3Cj0ImUakVA3PKfIOFpIc9iEupG
XQNB/B5losvo4c167xVJ10FY4LX/5Fexr5VjWrXtMKkXl10bmypYddzFnh4sZS5D
vO9/SL8EzZNKNGf1dq+Obaswgh2ekbIxvo+7mmxcxf72UPlxPQC4sK2BRtwIIRcF
khUB5f7WLDSnq2pLs6PrC0WB7v2HR40tVAi/vnl2avXzq8qQF33RUOJHFwMGWtls
FJw9mJbjXWfoiH8eHuUHqUxyS2kf5blVePIdPxOerUM0PJ/tst9LQIKK0Nod6Szr
uQ1Y47dzWU7+6g9zNFnW9Rz638ddmYs9QWHL9s0sTREbdsL6w0TMSY8b2uAD1CDN
pUajfMvKjTgSVBB8ote0rxG7Od+J4qUSIPgWbILVaxb2r9K6FWoB5yqW1ag5cwJA
cVl1+KJAxb6Jbvnd5FwA63hanqy8UxdeVEopHinmtmOsC4Ig8HjyJFDUTfHmcUbx
0I4E+6vPI+o62u3LuWu9ixt4hhygifOYXlUCb2N0gw/VX0JJ6SkN9P9S4OFmyIfm
DWal2ZBlUwH9YeTtATIAFHe9swEq0a+1SUJ9UsPNeIhmNzXkiy9Jx8lwPu+AzJ2C
DCa2guftRmUXbleQTZhqYkupQojVu+C9+40Sjl0HBPEoS4izkSk7TgpFXggMohGI
n7G+wQzogq0j1cXVHrlFG2uJNvzM1RxoozCFdNnPV4pC1CqCmDDqDMdmrDwRfaPK
wIiO17OYA7ZAtmFcf0Xow75Bp5UJMHiZpUEIrQ902XE7rCtmp0w5RR7JEyln2uwR
lMo/DKDvSil27FBCJ1ZKbotKnqI0koQjlqcWyjN8YXaW10KXULUXPh5k4cfTWTYA
0n2kDjp1+5++PscWGGSVqnrzGPjEEij7BLC3i9K6CwdwCw6y5E1dZKyTDnhbzhTz
RNiREBDb0sBtDpUn/jZnHMz0k/EwgVxpQ7Ua19lzpI5lOe6XpFKZJVjGoZNLGTdZ
T7lPlGJWd9a+8CKiFTa2FDyIaB9mZAvFzb82uYJ/9RJCN7O2rjxKSqBBbZZ3t0EH
Qs35AcXNDsuDKRYZNMhWyFC4Sq/V9GBZ9YodFxBOSxIHdv0p9EGSS/DJ+gJeEIg8
Au+QH8SN22z6nGAF51uIvTyvhPttTyQuumgQQzgg4fPzD+7Lwnx1EfNofHaGBvgj
lSBBVN3KWkCqvwOsBBiA7Fk6/Tw/kIwO+VtWHasYe4KcGFWmK/eaL4LaEbaw+bbc
l5N0aMequyma7YCohn4yVOokHJwG3Kucqzc3kliaFT/8pYsV1ScnGpnLWN/PbRVh
AOpa4wR6Gn4W3QgGO2AAXhV3Y2AMcXvTKxLYz/tenr0Jx7UQn5KRhjvLdBnckVY7
bwDLU5WyRvagiK9VWCwLGUESmevg+VV4uoNr+W5zpvaxbhPCgiAXpjmNvtxxTrbP
brEFNpD6lfa3ssE0VdprDthhoROyMFUB6IdGjA+/A+3ltxC0zhruKtSfUCe/AFx/
fnfm+tiYJ6JoP11MDTeREtHkHdCEaFT0rm6PNsLVuxrLM1nC0JXwSnOR70qa4AIa
Vf84zExZsYjKn6WTY0T/xHOY9DE3FPM+NLkcC2zu9gqNRzia9gnDZGTqpHflE5MO
Jnk3faODyQcfhpN8yJgCjqlHoHKr5D6WsfgvR3ZbCsXHNtM/y1Qq8DQTg11geZE2
F0NWnWEeR/eCsRcNyeVtH60IaaqVxEUERbjfa16jfCnsGReBJ+PvFpxAjmfhE3SF
2grWjTDrIqlmHLR3GAHUzn57gcPhN924xw8ugyijFM+MozJUqbn7F06mJUXKOMml
9ivdLt9tMIpeQSNUsbc7l8s/adu4tp6ZiUZ0Cei+eqCQR+zVIKYQ2PcHt9jx1HVO
Ks+FxkXxgZua4ehgqrxrEY7zl3NYncUTEGeKFbrZIrRIYv2USgg2acJnj5r1xeV4
9FniWnN3xEeEp3CbHRsS/BbcP96B0mYJzp88re+t0/QR32ahLKpTVTA+QNAjn1Eb
z24/CsNInL42twxH0WbtvagbOEB4j02Ig/FOrXUGyVZ+kepQYimKoPhRQkqSXFLB
z9PeiMc5M0cwxhuWp4UVqC/P4FHpV+TTvMWl2akcGjORSfbC3OcsgjimQn4KBDaK
MlazTXmrCX8rBLWTHE/W2xjZKLvjiM8uSheZsdV66MnGFxnmkj2f/aVsR4b25fLU
Erqw9trdON6IZejIzmpQK5VZMYhA3y2SYQLNuX3tNEf65Io86DQH06QUMbVc8rLn
LwPv4bWCa/8U79xrZg5nVQhxZIbvnARSy/CaTKN88Lqffy84ALyOgXmq1d0tSMn4
+OE9Wd7/DW1lyIDoHkc0mnAONbmvVNDuViEzsIQl3iCAENrGjsy9U38ePomhKTUx
bsWJSW+qI3t9jxwLJbV/0mOqovnSNASgBvJCev05LdJhUu/wE4plAfXK/Y7M2yRg
w9d3ym8V2iwQi7/N1ZLeiVdoEhyRvUfRTul++PLAOJeAwlQ/2lEPfdL6v85fkk9+
TRq0ui70ZUadqnDXOeM6+1VFsu2xwskj3UEDHEsIDwxlwtqXsTuaVks2Jc9U8qFX
tXxyq0IeVjH/qcFqyZx2s/TgSKvDgMf91cqluTZRNxvKarIRFLuqmkEHyb8Z81hd
Rjf7gLHSJNtUGcyG2Au3uiK/5+QI0sb+TRwhzpVDsTzOdCLzVXS52U7jzSX1/S9P
0zirHOlS78qvZh7C9LGbnwi5Ax8iwFV+xlfm+WXLQ0T5F/LJhWwVELEosJjRrIjR
FFjxiQuKx4AkvNybdyUJn7MfYnyFxEGRq6VV4yYwM5TUwK0K44j1aF2m7a1ZvViz
ZCUA0ai+H+HEYSCBxJJI2wDcgd4ReQ0ocgBWgCpLWgF9IO/kDP8whK/9++6udqkL
yYKX/QeHQf38O2oprcVGWm0sdUK2azLA77pMZ3hw3ySaTGAdMpaaLdrJF+gPt+m5
o9xx0yP5Ogu450YoOqu8RDO4Pb5i21Le71LAbxwIJtGeweGM+/qvAP3wavyJJ/ka
/R5zJo4CqjcwZIuJFCGxNLkFpIGD+DHIYJkfjW6vF4F/dpqxE+K1QpEPybpmOaoT
kqZiJlGcLT9N2OXzKRGGxHXU1TkcJWWNwIMKNF+1k8TM9LIQMXcBwSs/JPU0MYcb
0kh72R2yJ6T9RHUm3vxGWRZFWxW/MKka4mPj46oo86l/oo4eB1RHmiyJ2vGULlW+
JIBz+T2//WctRrSLCGTgHuqXKYWWLNIwwpqHZFZGLvAjxs2ScTsPwkha4ltkWm3t
EIX+F78mQSApvXiUQ+F66hQfvDYZdS0MuWQZZN/mx9w8/BvVNvh48cnlcxBbfrzv
YLJnZ5++7Jy20kYPljGCUVsGiG/6H/mCIiX3vr7Smvgi/IhLHUXc0CMaNmxDDivf
c83CQjjLI2aRbWOA45E1vfzv8mhdhnihW0rdVhg5sU7m5N7HjNdHrUluDlRjoDOt
VCPsmt42bGEKNfwCyKna85rV6CFc87uuMWxqdIkZG9v7DKH36D2hT26ZxRX7DdbP
VO4jdfuojoSD0LPyf3L6LELQwywqYzkHpUhtXMOCllFtlA2F5WMTD+9CJopk0+xH
X9FHSGLkIdWdu2UXndPr1My0j9TmQRPSznTJuk80GumXYKKIE0pdoylwDbqJbBBC
dTp52hS4ThzcgCwCFYlg4cUUH09FpL6MiBVV5rBkXu36WvFfsx2yKt8OnlXIzyL5
mgrupfW8/fCOHQLyQQnx1tteey4UpPVA+YSYVfDPc9g4S9Wm/PNkVeNprcmRPYlj
h830eKk2hRlfI1pajN3mIPiyO8G9YGXgjdj++xNYyJbhn9ECOuHQjEWng7VekbFj
Rfx8iOjdn54S2hne+tVQlfnUmWtUj59hU89FQBRjDkZBTtSfLE17sJ+ypurmeX85
G6XmIfi8ZJp/QAvyhZ7flLFQ1Z7whDdvYCYyZqTZDivL/UfrAUhA1prPvY2NNDWT
R9NyJp3gMbHLqMXnQLXE6chvJumCx4ltzcuSijbGzHFRHsQB5ysb4yh6yxHi8JfE
InSdbTXmfp5BmanKviCk5jpAHV5sinKz9VSbSZ2WdnCznD2yTP4wKoD6y/2bJ+c/
DE7f7AlBknrgg7mmpexS6O/6gwlCzVsuGEO33deSLcCSm+LATYJ38akJVXUsbDzO
PavHtXkSvBjl8OsWJHj1Hefzr7MB1yJhQWawiPtZIh29rDp6g4uH2Hk2BQqYl2Tw
Z8MV/wQhu8oGPfa5DGAOgGxsiblm7bt65MDfTkofOE0KwXGCCMsccG1boyTzZ/Tp
XMOIVogD+2/HIj2a0D9Co1Z49Bwzz8lqY6tIFtU+Oi02a59gPW41RKgRthP40iU9
8MN30i00Cz/fqHNTDql7peiw4nG6BXdD6wIlITehTUuxmBPFnWYYLuXew4Fm/0Q2
Dgjl7YuvhfGoz606sR56m5MizshSc4zZq0IKROhjgQmFdEtR5RLoYkt6AWNhO78n
H5fkox1B4pGq6EOCf2WbsQ+ddbzMy3fgp9f4TFhoMqrF4H5NLL+DmqiF3oW0zsjz
iedp+Ak0mg/yRp93LgXTNvRAdiGZoXo0k/vQYndLcQzFDWkqZuUDVYmSdDFnsjOR
sGCcQ2ym1BIhoHRUfb5LWrWHCOXeE+xwsJc/IiPmxAZmGe4q3/G8DJ1PhFglVkBz
hast+qHZkLPCGyCartferW4mHIWwDHPU6oApxb3qoVzHvjOe49VinAJRJBCKRoIr
845eB0KV/OvHxhaN4an1ueK+KIHCT3726TGPPJnWSu5Nb2pHsy61+3OgooQ6fsP+
AY6/QNaJ60Lsqqn5OFc09mMXOjFbi9sIBN4Zj+hOQPxzxXXBZ7xlL58vVfGcuwVZ
HpG1qkDuioCGab0hYVbqTPIIyiHSKwo9j7JBd2YeDwlW2OrTkTYT3GAK5gITmrje
62Wpv1itNkdyrFp43fvm6llQgmR1H+hHqSd7sDm7V7lx1/sttbOHubayy3Z/zdB7
lk4S9eTbuf3HwFs/90YRPNiY3mpJ2Tr+DpIcefOkVxF0LFh8TeG3nWy4i+qV2VFZ
xfvqrQLC4dOzTDcADvFYCPFXSBuGq6ToFzrgIYUJjyppuEFtD6+dDs3KqltSL4it
zE8x7ShUsUmHv5WehqqDfjy8Sc9estdh4xkKZyy4wu85k/9qScMYBcG0De2oOl44
yC8mOP+G/Sj7hnKRB5BwzVnwLEOm3uwckKZjr0UnWDInruSpJW6JYY9+ObjGFdv1
1imIpPkSDTztSRYElZhHJNnuWSw5cIgy99sbLM1Z8jjEEMDlSR+eToRzOMKOMX6b
Gxt297dhO+getw98b0WAfuDGFBjg0A6Ft8KngxvSqHr95czaR5rNHE7GiTGjYUof
FR6KpfErr2VUGeeIE/hy/abAgBzUgLbk0it/l5KW767Q0Oj5LzU23TMu90NWeZ+2
8lXCBQL7sjKNXyh3FMsA5SxmIRc7Fq4qfrNVsTwAbxIdGChIxN1t57D4FZFDe3wq
CLz5iH9yUvp5wEuchSo/gFegpfZwqNXi7Gp1R12FOpW431IHhArvd4xgxe3xVjDM
0t1JPrvH/rB6i2EEXeTddYpRqgsAlpvAeNuByfwELWMweQ0wEWcbH3vCcbN+0e3Y
IsZcjQxmPCC4XJdBRTzgKOGOer9ClJzAgiAdTqYMScSsJnDMwtIQxvIVhO26QwzU
IdgCmLvEDEgIbz5n/vV1O7SEE3beKZCRABBh87m0693hCy2ITMXY6TIedjdvUTEX
zPP3M2aczGqucKyUqutKi1zo5xyRfs1p0YhkAU5X/mZwiRFwVWm6qesZ3LPllrEH
7gbdzrnUgITEL4cJGL32M93Qes1HCo2mM+PNnsShW+rzAlGwO+DMGt9/50dbNsyP
IEdWBa5K2GFOE8MAGBXvNRpwfYXbN9e8rw62Fe5cqvz6Xxc/Qxi7PDB22OTf95PG
Xxu7UEnqTHa7hNuY5PE/02dEbM7p4WyZVz/lnjdVBE28FEi4wLsiAYYZbJDQyKzt
rsKl3JB0IJJDLLwsCVT+vLxqUod5IQsoahWdGdH8DuVoK9n1fQp7OHdx1CvOswQU
nXb2/2VbXOcRqDbBSX/ubxfKKF940pP9ucBprb+INNhWysphx35J9Y0aTs3oyj+G
lytbMVm1dZltjQgtxudhBjYohJcTMBuGaQ6BqDe6YKELGGtsfaNUEx13z15JQuPK
Ta0J+BqzZIOntYU/uQPHZskEbG+Yp7rkDO1oNF33AVdoQzX0wCkLWt1OPRN2IzAj
qgTSyQomT+nidi1+zwPKgyVdfWzo6wriO/NmKSYHHBR/zB9dRzspRAIOyyQnBX89
SxwrzcHVVWaScQVTnjK+4tNLLetzxuyom9+aN+46TbVZN6CIW+h1A935iOhZ4YUz
QD9i0RpFaTiKZfGTr9BsJC/9dvF5DcC7CYpZXEN9IsNbZPCCDXnznKO6DMdaT2o9
n+zoTl4ox8wqxUMvcuo0kcGb+5v8Ac16stDzjShecwWt+j4U7BAARDe1+ocqKvB/
goO/ZBynqY/QdvrwF+o4SX365jWEnVXf7sNLPPDOqDSxeKVx3aKY4rBVPQbRBhWq
qvX/T5dS5UOgHD+55a4aHnKlW5/4UAnO9bmkuQ3lvIC8gWRuWMeM6joaR8RPIoWT
Ty5IKpHwr7ywjc1ybNEt+m5Kdt/ksQ3caKW9AoKlrB3Ha7CRjnaRL1lpxcNNLn2H
LrOmlFsAKnxtJS11rDg+5aIzcrVQJ4ZPK15h8mto2VgKZ310AVvKv/aA48n4qbMP
K5bcsQbQ5DT8k5mV/ymVyOnmHMFYOwxAYUQAftieEpHH2XXuSoqYt4MeoVelIyXM
ar2M8IBysPTarCOfKLKuuekJLi9GFi7Txnef2lAX7Ku36MzBfr5A3WHP//G5rNJh
d7A4iJ7GODYFODrW5ZhCfk5Ru9Yy8T8flCUKyTFpK1cy6RXSDoc0pNpeW0Pj8I19
5orLrJf7jlk3OQtTiLnM8HdtcNqAGdKz8OzBk03aTxDi8fUKLoa3AQCWW1uYJ6SP
iMUB3fIAnl9rAUbk2ex4msJZfXAHON8PsNYcDoFiM6e9EqumzB4jIA0kBfj0SLMo
tSBdYbhT/EAKtFN+PD+CkRfBj0S8mcjsz5zNaFPk77a/h5wvYZEz3UsXX9TG6WuK
AEpdJshadj6GQA3ftFuSrAhgxBISXJd/U1xZWiBJZo5UhpmIprXPle5hmtSheRbs
Q8FKfiP7MYzPtfWvSsT4baxVo+Imo2ksUNFTpd3e2vdoez+RqaQzERDQty64ZbbW
CU7odhaxbG7cHWbcYj0q4QdAnxtJiPSAwXHFZzo6UXcoQogh/UaOjhP/6XW/P+vo
HDC3TVqZf8vYBoXL6tjNUR8YLDRmcAgFPY4PQR7q+7s/pQDd+TML8IStqoOmghWW
kYEJygOJnUsV4coVsWT9LYp9Ua2nkDyhtpR0BBbURwiMpWWADhlSdcMxfBQTtC2B
4Tt6Qbmsy8NBHRbKTWihsoe14tkIsg+m7grj/dt+EMI5yBxCxUDsv+EVngdhBxsv
TlVHiRLbWMnMe5TYIAd5X3UUSvz8kBmzysJTB7TovOf9f4fEF3S2Ve2hHpUVzB+B
xyE1tZBBesDDthArOD5mueBgSkwQn1TfNNAQIm0L5jyCFsfycDRMXWklRWaZ7BjL
8ZVJtRSOd5lUbzvnC4q0aaNwcUTg4pSJrVgAWmfUNoSccvnI4WgNl8mFT/aaEeaM
8Wp9VM2ftEPestZIg1rp5HKpk467ZwU8kUShex3Zm+nvxdkN0xBek2pizkUV4+1d
VF1XWm0LtlsPnzIXGFbe25IamzPK3ecQU8s03JXtDM7qbHadDBN3GLZ4SvAGo0h8
5tV5C/hhJ1jmNOEXUhZb9lntSmfPTNBnQocZRXmw/ubBYMTn7lti3Xi4CWWHnjmE
43AtIxqzkj1vRVH7XOue3IHKW4wgL4KCBQ9m9S7YhSSoxfSnb6YIX705ypPuUCnk
TiI/gn34Ma4RNLvmu/Ty2sYDuYwXM9otqvr/uKnJXCBz0LWtFiyS+fKzQXA2+VTB
LXso7LPqMJ8auMj2lDT5rmJvnfKPywMBETQu227aJ3iKbmQTeCx1u8/1B4EuxbcE
X+lMGYqUKbYxIzsBeXSLZWoJAA8/bUpn4EG5jSUiiTj3v3o7PPmj1yCftzGz/6zC
TjWWQxjXq9M20xY7kvsBs8hfKFFjxTvL2gmGVQjZvp6hDQp++LiJ4HoOiX6aw0th
g4WTN6JP8Jk6cAMdWbXQ6DpwzL1jzS5H6JDMUXR34uUdQCrPoo2q8XHnU+ULOWvE
8CX8wkep030mh1KE0WBShiIFNsHdCq5C4MoyfPd9eK8lih+WZitt9OVHAV6lq7Cn
RmvwxcvuXozQ81mX6YDPT7YsGYhCZbRZVfp8rFoER3n36NCFdF3wa//1BAaqA8cL
HL5ZH5n9VFrxxOmRdEmOA0LFiMVch1CaFfS5XumH6zOUc69/9JIwLWZ9WQU3B5A7
svSdV4elSxqeiMnIupbfuK3Cj9V6+DxVPpwQlm6aO7l60KZZSmaixAspWWZlgvtl
XdO6FE+vkXvX7i7rD1cjnpkRpS2DIlflnO0RF1t7tl46ZnTin+OBhyw4Lq4LWsZn
0EYTnb2/tEtuUHmRXYslurbjAfy2iTsGplhhav6dChYKEZvW5oJHK3GAoRZvhdlf
bA3FePxVzhK6N9Vl1D3glUSZ9nXpLB9DDaE9OyNQR6DfRV2QbXq4UikvDKqmF/Tr
n1450jKV0rlOQvZehD95+CV9UrxndcbmwKTAqzei08EP9fQGdbFnCzK+Pe9ZnrzK
Y5622H8OsTMkspR7Nh75uLl2X9/sB/yLGZ2BlopjD/m4DKr7H17+vhtH/zPvecjL
/bIhBVYm/nvTUgGmrUW504ljLaYmeNGM0XQ0PwpUiG+QGQ77GvgZfQmPaeIhIeIB
jwIax1EOL15tcetTl48O1PiYuCI7XJ30ClgM+11/9cRQ6c1CnDllGnqXzXcWVCL+
IVykLiGagzG801QGXpSrfE9eqj9Pl/RSbB8NAVHtmElnztBKs7O2Bcjb43SubhXG
ZiKtsuso9to0iTL/R+IK2Ug5RXzAkWbqQNGBJ5/B18rRxz+c2ZY8McJMF8UJvrzI
UWlokIEQWiXsVJh2VpjrytYjaj1vhNf7GHdCh3VotNBMDgVTW+8uXKC/zxaSD3ki
1wXz9OmN3CmEqLh502S7aG5UPEZzvePH/2G00gLwooiYfA3qHEaQszlxM0fYsJWW
6oCHYB+TLQEd2nKtswlqes5Ko75LQ1QUStWIjqokicMQMXAzHC6WxaSCdwltSr/E
dU9asgeLqUctlpmvRVPPXbLtceTzdVASry+Xbp192Cka9k42NnwoaNr6ONndOs8V
a2Qdgf9/XySNfLFwrgX+3oKm9SNh8POp02J2pEBhrPw1bBkntvspk9EqA77xF/Bx
XZ5WraDjbjG/V/YXYHDibPsmawF4KSGXW79YkFPW4MRJJCCqZX+Lplb1aGfvUuqB
HeWfiUm5CEHeHBmz5k3wasUK79rgvt+AO9aZyinqUKTcrdXyCN6Wf0vOlvmLoYBB
ZV+BJygoiWo/A+XOf0zjsDzrNkUIV2MYup1suFs5mxcGLuCQgbrIIqlhDMrqHFh1
6g4e6wVoJjwmfPmUwzrQixuf41bL/1pvOiEwT8Bt0iYjnZjIAu5FzMdySS4Wqms/
L9vrcERJeaqBFjK/CcNh/TC8BT0xZh3FdtRYDFZdBq0XfGxSk4tm5JhqLpb9Q737
fxYTSeiXCCHYbHcLuiw1iZ7FQae76PX3rJwNAHNAwwHR1JAdO6ESbuZVG/24w194
OLGTcwzHHQ2i9cPzmuEbu08+qWFyVwxdNcM2oDXgxhAnxHynFO4VlQI21K4Mx2Aw
5sspq3MJs/OZhc61WDGCK4HbDC6Ij+NkPnJ3K0VkHH0Cu56S6vA5d1rWFg9BfGUM
hrSUpfnf7162uk9cEu9kBukBJeOSBVjjyZ6/X2MVDAcJJ2S5efelRC7cbDLw9d0d
L4USBE7cyCkIsbSIxDqtu9/F3j5oLmY0A554mx8UGtEkYFIPf+cK9vSiT1mlwX8E
sAHrp5AyhUIECsxlmj8tAaF21UDA9jMeIWtd4SFM1wKZRZhm2W2VOfPJh5Ph11K6
S6fWWIQxLU9H+legQsxX3FR5AFANfxMppG3/x04vvN4DmeARcGewTGRQ7dAM1Oig
IEmPp66YMElDW45kQ64xvtAJt2kkBZBJFeNCm+zZ1Al0ct8+oKm84OAYAkbqulMh
VZHLSvLitIjTovt6jNhvBy0947MNX/VCC3OKNDLYQKj+AC7cWjv2PYOz3SpBZtHs
9MmEyo19qgLw3mT+71Mh0GWL7FBu2DlfXDjFfMJDbvlCeBDn5MLqcA43v5mfARIA
AtqX/BRtmIcNp90YoegEAp5WTdq12B6WHFsKF2vKeoVYMMPhekpZBQvQkmsozldn
uIxBJHR/ZepKX9YqpDSFstvl6DqXlByxbkhOUf/CrAi00Aub+guz0NQ0xYDW2oUS
lqdiC6kBcq20QkeUf9DVX0IxI8Nm5NHbKUka9oP2HDgcKmiQ0caimQ3FhhsRYxS0
izKOns3SNsWCgFTk4Xaox7EkDLchO1aPmGCZwLAP5i0rZrq8CkNatXXTgtURr0g7
z7PcG4KXBh3cckBFtj6yDMiHdVdR/TOeFmNse7rXagTpk4P9Lq0RAkZG6MX5skJc
ZqrIVry5/9Wn9gblCySr+WheCdh/7s5ojpoNdnW5mYgtSwE2qlcPdDoEQ3aGU7Z3
O3GgnBjzpvMLVaXy08t1OgyBkQqVl218y1M5iQLcMdZi6VODjIF56P+sXyGJtQt9
Jzja9IQqYSsP557Rd9/Wbutz/67EuVFBHdSLhyS5x0PeXyneCZQ2+IET924guBl2
/dq0gwoKNjqGh9qgy9tTgKCQXgGkmy1wAf1SQMUAQ2TGdFmKd/WPkEIMqFpTxR4T
lX3rdYPpcqOx5GncoYmpbzhmMlbra0J8eIxCQMDTBTvF/NW9kWPl3jgM4zFXB4Ut
3e+MhJ3PrWJlyauT55vSJR/mk3lx5svyv5KmS3CAd+uopS75ADdT43BJyL3KP2wO
T8tM7D4DSDDNeghZhhNJPfCJw1T1C+hXKjMDHisdRQCqjEYZKJeanay16kdBRy7g
NxcPzuGyyKQeRxgQOb3SclD2RAmNkNhdKQDIQEGUIMLTpBTXGftpbo0zUncmyvLn
8OhdJgoKnrC+2eFeWabw15Qci5NPDL8y0LvF6ftD0A7TeA7nJ/ihTgKApFU5YeHM
87jxyUmULwNXx0Yw7YI1fiz/+s3eMJfyHrA410lhcQGlS+jfSXlBB2zusHktfWWE
Y7zXDwWP4cv3IXQIkzVIuismiRxvbFouJtaAs+8zrJmtT7f53nQGgJM8t80FLCqq
RgiUUd8wM5d92GszUi7J2+OwbD17/i91oprBSMI3lVWFxH82UCeFGPedwQeJy50v
NlfuxNEEpDJsQDXbLrCn8p1Y7ypDoC0qTWpfv1kbrk3fBP8GvhRuUQT+rzpZ6g8Q
aPcT8xkIqtVfd8frGLzzVCfEQA0kNEMKJQq44OHWoO4Q3wcG/ghcqanOoxuxxADq
kWDXOxIOZQF9TtFQPtk+vCBH13t4ySMNKmCL+QCFb8ZPms5tRqr4wexrP2xhWfM+
OfNXsDiPt+dba41U3zouMy3gbgVpy7pLxS/mEjdiGbHn/3N8l32XqIdeP7ENZsQi
bzw/EkzdybqivQS990Gooj0AH4j3v2mBqhPdIrdjELSnY4QredVFurqFjz+bnmcQ
1Rtu+dilWhC5GtPqChmjbfPRRDJjVgEqkF1TZzYDPkdV+t0p/Z1GIdEWyUJUhcUe
FjzXZMsfNawH37GvIo28LnEL5+LTeVn9hk5R29BReldhbeCoGmQt6D35G6aaRxee
Q2Qwxpd1+yRGDXpDlPdj6ZaiqWEEnnwbTfTglHcW67JUvI8gAZca6OhBmrgJ4d3x
3eNIsLklYhqtnVxDP3rk8bLLpBZF0kCgtn2DgipYng3VMUYNdGoQ6RYLcMoSKbjx
T+ynV0NLKLKh5CUZNIN8j03VSsq9v5qslfSQs9Gt0R2ip7LZWezLZWeSz2a+2DJ6
6y4mp02AiN9LT56FuTuKISZGUX/Bp/EOblXg80yffFajdoGwZJtjjcE4BaZ0IqkK
ijH/b1CrwXYovgKAA5ezBXAzT1bFi85++Ga5fvtcEj6u3d03POmG40D/dO9l0mru
z9Lbh6mk7mUmcC7z+E6TH51Yq5SpCw3NH3Mvhh886APCz437fLR2zrtXdtUetqe7
6JjJObN3aMfRCgsUILe8kB7xVClVILCrYF632/W5O1aUThWUqjatXgfuQhwEYot6
SaBdxWo3pVy4/xXhVuJoHv69t3AGWxjCdSWTMhbqrgh16LkNGfK7DDIUSbPNcOWS
op5/gGuoxysG5ut0qEoYL30Mj2FY0s9+IULAXrFEAAf+L3tYEdCxYcdNF0tB2+y6
3Yz4fnPV4uoYoqRBmp/CVW1rfaZcmfO43y5FV8m3DlqMm2XTvuxNkunAz0cyL7Ao
UWcIA89OOOEzQ+VtpzOJgmyGOmgGS5162UfF3agYcvAJsWrJlcfUFqBegjiAS9Hp
VI6Gd+6nQk31T/z4Y7JSH01haBPoJ2F+6+LisvMo0yZbU1qoELxPv7GIMPEIixH+
5WCjHoH7qYOEYUFB831trtPZMyvC72Qw6DLROxE0ZAMVx7JezKWTGEvsFeAG9z6p
B/RzHmjrilRMNqo8dXungQ6giJWJQXjvrYC6ha/FSqePJCDpPvFOv2iYYoM6sqUt
yOcpQBAKDAZn10wsofo71UYnD7N+p2oq1CD603V8+ajWZyDtu3tgtrI5933oe+jB
6FXqx4yXO3LrcSiMXcwpKS86eBN0K9aEbYlwcitCaiUNqwLBGIv4WMh+mVk2TgVb
TW9UB+E+ogxX++BRxcGF18qJsasmp0/95zMoO0xVz184Brs3Hywea0de+og0z2NU
l36oNF/Y+ragY7HbSHnMHGPiSqXH1zrPl9vmnrwsvHyi/r4ee+N6Lu5Q86ojuVox
dLBiS4iBCiiYjdrnuSPO0ABXGA42gY8CntCjwoIVbqCLaHY/3PIrZBg9Zlwz/OXs
Re4SfpwDyWDNTGIk1Civ0HOq53MK2fz0YIsiwaVXGGvVih9j2USDueJ+u3AuA2EK
ASvgK/lC7LKs9hZriUF0pE/9Sd9sT6o9nMullLkPw2RPBYP5L9ATDITNf9WMo3uW
0S37InFITsl3uLPzji9f8mt63RVkJcyBM000HT2G5Ly3RZfPEI53Y+fZHfyHCFPh
QXnNtrbts/UfGdoemjFZJsIiPe+IuPM09FDGIE3U+m8rKGWFW9pzoIhslnKdPRWs
Beu5l7/WkLwALaB2bVorkK/n9ci7B2OzwyC2+S8tWMnIO/StzId0k3pMnKfNxuyG
kCUAniLCmenCnKRnrCwZDDLy9FvNYbOYpEXa3c1urpvENDnKYDyQ+fwW0LZizmCi
rB3jmsTnmUUeDgum9xtTtYoQREHq2D5EPA9yOS89aAAcybsWBuAYGagXToLZBoZW
hPa4ioxt2RPAWR9JqAza7l8Zav9gNsakhIAeD/E2WsZc0JKxvxlLt6wIvzmoHET8
fJm4o7qGfNDMvxQ7z8aONq/ubeq2UrzM3qpihtjLfpFQgz3xE1JWjDFW6cub0Xg5
GQeobTjxTaGJ8y5jBPuTeqWk1b6BqG9N/9DdR1d4adovQ8RjjWdeHTYV50xHe2J8
bcot12PhEAtz4IkcFrcXK5k9Z0aXbGfmH7RcuujlDRs+FNbxSAHVS0tEyny2Efnn
Ja84+f816XhLrkNbZ6486saxrGLaosV5eFkt6qF9WwZHp5lK7oPADYnvcSUyQx/X
Tr2A4IpC5tbztgxPPtxEW3d6GkuLlwvrtjo/JER8jnhfpbq6NTKeNJSPDwRLi3bk
0nSNjOIAyPJjSlTjvW2WDe7Rh+uFnAal0bX79EWQFo1WSlI2URtwiVQB5L1yy53j
YCu5575YWiWBbvSSaHCwehnerXifbW9auFMX210+orfdvZFbo5Ml0vaPP9vfqE2d
J+OHrt9acYBkBtJOdDoru5YbMC/KMlMNps16OqZrKqz6U40xylYyq2+d3dhdn5/a
G4Zt110GBGVaCdjQYfXgi00qnck5ZmE4+8gRy7nMJxOpQaCcByOHUyaPyKPLMXOR
8uulnEgahNGgPs+/BuEDWvZLFF8ZMwSVPRJO+TbJWFRhpHa+ZAp4qbFeUW2+o/LU
QV57E3llG/82B7y/XibwqlkmJS/u7P+HzwKlg6Zn2DXySlmgxm1N8DKtRDvncUOX
SaTcgu0U0wYx2+OK3unU8za2aAF6p4oKjGxKOyBdmpby3E2zwYK7MrSdGB7hwcpz
OgcLgraqecNRpG7hHa0UHpsg0xXziI3evnvO6mVlKBV7tiYK03kk2pv6QmUSvK9M
UBZjqdQIWKTLZmbj+c/RO7KlCb6eXsiJo/fdBBLnXwPtp3kpkm+Mrv5C5mlo4rE8
ncib4vDkBdbR2BVxmMyjYm24DwSgZqixKfBMW3mCUTMNnxRblgeS+NgDYTCLGobu
Q8kNCv3Fg9En4b1KF/S50NGSyU3issLHFZv+7PYrgK1BW4h5UxZUP4+Co+lRedA5
cZg3IfS33nKBPTlcwKLZrWOwuKqFEwzE0wJ0sUCxzuu3I1APB0AfdU9E8mSYgSHI
3OfDATqJEjMMlvVIafLvo+8G6zfqcr3trT9eMqeTib0rWzbdfYBMRrdpE2HzAF24
I0aP6pxz0WPJhZ6KKm64e1P9N7G8ox5yUa8yxVejFcIZB7X9xqearfiHv2LPyHBW
VREuHuJpp7z/2/1gUtjDxZ2q2RANH2CwyEllGx2cLV52vteRBTK1AQ31Aup5KIhk
BVcFA+7XMl+ZYHdKgbKjupg/JkV2afHoEjdk0r3kfBkFWG+iwO1WjuhxNLkW3PPf
IPjj2adPK6j+NcKuYeF7zhnwla1lMHrrNtjvWzmEfIMP5GS5UR3ucBURLKt7WFE2
E40gr2ERpvE3e3JvR2l5N+x/ICpIY1gkSK53gbXCWNDeelYp6hyymBC3+bp+R9GD
LimpvWVvWzZOrX5+lVioBGcZLOFhKi4eJBqZj2mg4O9C0hBSEmS2nKQqpzyS2MmB
T8heHLvmNfcVAgF1H5FvyqpjYQ16dwxLuvxrNm5ujcXz64OLRA5NuFpN7tYgHloL
zv227eP4f+zAir8wGLPIldaH8uRDPf/TsnoM25HnnxF0icrMJi3eubdkEsjjNye0
ds/YuVdanYlg1l18QT3CjqzslHdM2Kf8wWvy5D2K2aC6GsbqIwc/J3Hmd2J/Rmmf
2oPt4EvgZwCwjSEZe6YO4yCKtakW9uSwmnccMoEmKofH9KMI0EQJNO/3juYRwuHg
aIE/gNqskMvhdwwH/O1gUi1LvCUaVBL6KEvAYtx3SPEToM26zgMa7IVrax5gZFyr
FmFlTl6j7t03v5d+Yn67UnTlUPUE4HbOde3/of0PS6KgvXSleQn2myLDi5Himrua
00grJ0ITU+yyunDKOn5xAjm/++UhCgjexBes+aGW6cIXUp0mJ3WllDc1kLCIcWCF
8dBhqxT9LFn3WZTP0yKZK057+wW2RkQFH9WdjhN90NObC+lIgMIREhgvgaDdtRXv
ZcsDMJ0bxfg7v6zGvaUr09YSgkzPWQCrTqfjmPG3D6LjI7vf5SDuEjsSkJGPdri9
4tp2WGQUnQddFgS8UP/vXR/0/LsuuYhCAVrbPg4EPGHhdfAtyPegIllazFSBIwiL
LVWSsu6lMMO6kFvQSGBCJzu4v2G+KHu2TY+cZqGmSB6i4AiTmfha+p37zTqv/8Ro
B7xwqfzOWAcVnxD2rfEx5A7BZF1lhhVCogMqnPIGxZKMvqnk03Ime8SxrU+LS8qj
daD3nCICo8jCWXKy15PM2f+aDlBUQuSRLlKSK3e4IRj+azXEZSt8kG1U0hxp1n6K
bkw15SKd0fHkYPZNmflBW2HfcQaPPX+81+BgbCL0AlUPd6Fwwk1k0sM3cbU/Fs7x
4Pz/RuxLqgHxKchM8ULv2XJfKCqcz/vQn0g35H0Qi2PcD/YOrs8r0gmMfnYdsHDX
rqFYGmqDVf/t+lwPh/+K8Wjr04qTrdlt23nd63+6ZijAtcHWb0+NRMs6xxq73Ne3
o++qq0Hg0JAlxBDd0usKQ65lFQkvdK7WyYrcxM01Wsz+Ta0Em0YS9yWjUa3I+rCz
3hYRGi5eXVE1MaF1llWxZ1juN+b6Hh/7xGmqEpVe/A+q5HJ54Bh7zLMRGCylZgcZ
lD21HjWA9oEDKd5lGLUzHCIZOq/nhRX6ovfYh9fRKvQqF5cbuAIbalFxDY80gVmG
9izQLnAYXoDG9aMTdhzXs7OrvBqnbyqPV06Sti/uhHQa4QSqgd5JzncjV0Qd1+br
PHEurjuy8zLgnQ6qhIIioaJ0dHgWXMQkhg9s60kHJZuUNKO+3LIae0EWMquHJLEe
obT493k08rKlesN0SwRNZw2/FRbeEIqh8rBMr1RAL4t/C/Ca4iXgDGga6u1o9+hX
rc3yl6vFT7b0NyV+wJMlnVtrslM8eWHmK5DbIibMtnIZPOFQWOhJCnI2/cEPGYeE
Yw5PF/kLkf2i7J9jb1whJYTLUcJj6DrGcapl7sU1PHkcXdmMpHsiZnoeSg9+oe73
vCKLFsYLu4tUKcrgmnDLBkQGEfvdbqL7K77onp1qFuoVhakUn1ex8OoohilWrTI5
dmPyA9FMgnjIIm3YQm62mBhRWsCgTRWYaqwqiM9MJ4Chdu0AHtiXo9vXcWCjBsqF
xxNrtf3w5O6Jc7ML6/TDQyyuCL++kXRGk5DEoou4P1Egy513UQ5vj2hzZXlFAIdc
/dqBV4WLuqaPnuxgjypvx9CJcqz+2nvKiuwUgsuHB5ou9Gu+Zk0gPEhy23MAa7lJ
tUAQUR8GZEYbk4pR7sQKaFsZGAus4EUHs8DF6GvoSqonfsYvDA/mZpfEr7KRil61
OmYL/CvIz/cUxg0K+MmOUgw2JCgxXehPBAhhUnVQG9WOUIVj4Gaw5e7r7MlkytwE
iPiNcne7TLsC8kj5vp1k+Kduye1IGXjoLyzOyN3TJC6Tf8ZWBlwFtwNP3h86W/hC
Rfl5LstwPZPHUAf/AqAndyCIDRM5FFKG9hLBCmi+jlM5PafKALXkMvz3v6uPo5h0
kt/5AF8wl8WnDJcOfMHycveXDDaWny6wa+LmTMZeLRH4CVqKDiMzO9+cUvR5Hrer
pk97yN/kxq9fHMHWbxpSW/P3fvoJeEcW74zpuVovVcPA+Co17afeAeySkRNK4UbL
eD1BRMAuivwd44ZlG5XTLXm3lfFJgwra8pFCQysuoB9y/JvoNSjnr4A2kWIDimI5
7ZH85WRDhsqqD5anrdNnD4VSihCNKhS96/SxBAHWMQ0HtE5NdjtzKVMstwCNr5Nf
MVneL6s9DLMsq5Y/L5qqTxfeRX6qZ22JLHjwYNetXCc6Qf0sYAgFKsP7AV+RkSlw
Tl0aKEvZLmVFzNChf43cYMSth71F6xvAOO8CEJBAsLMNW2xwx7XgEFJpUdH5r3rM
iPWXXU74YipzcWoZQwwTAf+g9VxS/2tjfffT6Fbh5tA03W1v1g1WJhgQ2IfhX/U6
qN3AW8Zo9LEgyTKiKOQfbkYE9MJEUykWhqCvy/iQM2oCaM5oquylj18/uVT5uHL3
zP37th3Ahg3WfeIOPtyYNo/Fe9+F8Pt4928a03qlUqsrySjdPVPbGuWA3lWXWqDw
XLZwAogIm4eOgHAh2+4dH2EkC4q02/ze6BLsWVhimr7r9iULA8MIWgZJ8fY6BSUI
daWQtcOkhawgbXBJMSGhgdc6lenltEvu7vukXzk6ioYA+IIdjPOB4DZh3GK5LW0u
PqiMMQAboxq5y62I3bemCP4PfmRX4TCjdtaxql8ay+10uL2eHYyj8PyIqNz0Vjip
dnW/caE0Pe+izF0ywlNbqldLEte4OORdnG2aUfBoio9FoxcMz5fPa7vJOEII4sm1
Jzty8FCO4MyGkLn63w4CVDrNdFHH6bhG52kJANTV3mAR7rnZELqXY72rQVH1EV64
zCupvny/ARXOBiK6WvW1ooJ3rGPtZnPq7m2X+Gj5kQbOVDe64IFcmHYKLTtb69MS
raqLz4ikfedHfAQw0HW528P9c9Zrt8bRDuNS+srpmozQp6CVV8AGCWBbNi70Zh7N
f1uSIY4yGoFO0kzC4DKNXAZZBoTd/Ivs1gznHw3DYRaI4IC55mvAZrft7CPOPQJj
HjvgD79zpIVw8Vgynn25FhIMhTwidEwVSq1kJCb4k8tldtQpMB9U0cuIX5ykesfT
uzniStr3e6BzZor4dgPgA5VoUs9XSdv+amIPg0ScHmj8qP6z4O5IVV6xIscalcXM
7rq3mMjnouiAtrTIX6QQa3aylLsPCKAbCaIC+Cg7DLaC96vIgOrxRqWkQ9oyZr+a
8coOLcvKT0ngQTlZ1C3Ym/tCVMHiP66SeXXowgJOZWBfw+0ZVrSyL5JE6rIJ9wmg
H1JI4+fPIv7l/a9GNffIJUBkcJugJvk4wkZJUdiSor7vTg3BYLp8ts9M8bTh5Hkd
2fh26GmEjJap+Fj6GoTlk+uL+MLI/uacr7KBNEMpRKL0y0zKGijwD6nDqOSWcdfZ
wYYrWvLzPfdL3Ny7L2zRY1jMFZWnqzVZFKMPdUV/lXpxdAofdk9oJM1qTvyTids9
3tm/nhSGjwbDpkBpTO7Yf6+KGXKvTyCUtWsgmgC4fU3MVB/0m0HLW0omQrGzUGt6
xKit4khsWZSeOrG0CSMMwL9lTQaBjihWMmuLk7o7KVANJPD8kBHjRYyGyhkDkDer
upa9uGPpY75yPZCW9HWlkSNsUXepmnYSxbFR3yrtz9EWhqFnTDi87UswYCYWCuNb
qzMttqU68UATcUlmh3zsjD0Wsblo3hxiPQco94l8eWhJ9CAn2jj/rHH4VefTUcBg
WXgrvjScM24+6ryvGnw7Lqwhn1Ba0ZHFPePLP8SBu28u6mDBohFtv9LOLzEhBfMv
CTbJcNmpKF7q6xVq7y7bGhUe189WX+drlUXlTFtK+v8CKAybkNPdITceEtSP/Esy
ots758Zy/mzXMnCtSSuyKO4Ms/XSyjhJeCezGNTnbLJ/vC/YQOjDrgaE9TMXmcY/
ccAt1ZIpMb8GEoaz44OJcUaxjtLDMv6wmnL01sOV+tdRSCSscBFQdyIOX2F5EdB1
84WepZ+NeQr74ugFrOLgnwERsn0j84ZEwlBWO27aj1fPqxMFmhbAm5ElvlZDc1Ez
E5Y6wrSdt4vODn3VtThfzuyc2nFjJvND8NvU6ef2SAK2vlmRMDF9lOGsuF4SDw0K
tSN1+hSpqSpJyddJFCcMNfk5i3cjEhIuLqOJ3Mj+vhRaivYzVqkVm3issDtHTdEk
C16Z6i5NURqftQig9Oqt4PCTwziIec21afbQQVLowFMNccxu+p1PJptXf2C2VXk0
upxfRPmaCGpdb2BZSWN+ACXBCH93peQP2YaE+80Xhe8in8raomV5znTaw2hMKHV9
nHGMgq4txWqkP2vGjWTtZ16lyQ7taBxJEk7EVlxeyFLN5n0RxbBylsMmkz1spG+E
bIxh9Fq2UNUCxPv2tFWbB1sGCPEyuMlvKJXhavPHzX94dK+CQ4O+TwBhjnptXaBU
2OaV+rFTtfnUFsrSKKYC5+K0XLTIPJQFPw8zcVsIuDvsAh+8v0sud30UPTZs7xUE
kw8D8fBKq7QjV2wNncFQQcYNsI2NbpVU2Eu+YMu8rSYC+j2/l1BtHq1JeB7gexNW
aIQMkBfko8IXU5UyFk8vTDYRvhT1rP+f6rkY5qbY6a62UcV8GYqo8tVacdDT0jcj
2XQlOvM2i6ilYo1XVYn7L1L070BfFgzZ867U2sjwJBX87LTObdMsjwLSyumiQwCi
8GgPIXEwE9+Cs63lYZX+el8Thc5pXX+vVLQf7SAWbzteyx5jHpdmQarVa7j7St2J
jNCoE2MucFUhc4sGec8YOP2hPqCjYxyt2UPiBS0nFw+8Zp3czXPc8nxDf9Byg4mL
H+9IOt9yEK7KmUUmHvcCFkjJt+gDY7CCh0O1RGispXsoEVOHQENl9LzWumOpnuEH
F0uhScdzLOIjAvongxIOoW3TSu3ZM/8tqsv69PBSYysHHfGx2BLYinSCcSQZFPHw
3KfQhjEL8NmKWfJM/p8xWJGhRrZjHwuUHmg3R1UOgpqWp7HdM5YAaaMfLG6rHLrc
Vk7P6KJdXq/jKIRlrfmwoVqxcVeWzuex2nUegr321PzufDyGoUFKVUzpFxJL6KM2
jF4aMHHmkIGJx/42G+MX5HcHWz1jOurDVnlP1fr8cv2TFfg+qterU+EmkIwDkcmU
WquD5XrcGKhBN3FSh3qcbBW5r2oG+b0qLACYqanXvAyXRtHptzcvdnB2PD58ZOuv
6zEm48+ZMvw13mPpwZaKhTMjKQE3KlHKa7MhTRT/fcNklcx3WCE40Fw+yVFvKtmn
8Lmx6pYoUjo10XCUjTX9GlxHHtJFHtisaObPVft7WQwSBZ3VxYePFCW/kLSs0Lge
ym4z5bWiwUAAJxNxtvLsJYM7rTeQYAipHLRiBJj0O3ukiRi+8ZOfx24Ta44zU0gZ
cBzyLVG+rJGSCJ2+sOMtD8sXZPjuPwllqP6Yv8tFgkF/RVTkolI0Ek697PwGegBe
i9Gp/HZCei+pnaKLGFQQGcMEVf8G2v3LpM+eGG11VGhXR+1SzhnFBpue0YXmc03P
uXuVHB0VmPgho3TWRIJP/y5cElCuMqmj/1pMlgQxvFw3QRRKNHl9bWxGSSkoKdys
9gMDhffvHKDPqcs2N3VxWp24VGbz8Wvpoyiux6v3hr5p1ACFHc1I0DtuFzcDfhR0
9Bbch7sjDtLdmokZvt56Jn+CxX8HT1l1Qu5H7BgS6B3N517d7emNozJKeMoA0PvW
/5eszQJUoMjir2MeD61Ooy0iTVlts+Kr3sZKUe1NryA1n2gwIZufemm1miv1srir
5NZx841jVIV0l21SrEBlv17T97VKFqPenCZuMfB+xCpqMcbj8VzCiwzC7sw0C9GL
AaoZzWRpdaABM5YdPFEf0/2n3JpEpERUlqJ2F4ZLl/+Um/qmTtonEdbgRoHCl46/
AOqttoUESV0piWP6ZW1F6FqBkCgEm/vY8CY7+8hNDfk+D1siweeWKzSNZ7o7y60a
sMK19FmqizepzKlinrlOq6LQuKHvUgshDpukKBervr0NTxrCg4OXUyxoh4VgzwmN
OlqWtK+R7Vkf2FDRmhA8aLIbiVeGRi2D2B8TVH4GKM59Xi4VxQ0JdpdCfN958yER
siUZiPzYSBumN3LTHY84L4lKrl15XHgtBs8Ccbhq26QU8ZBY0eUMVDHvo1O6BETU
EjiVUBaxxbdY9ZR7z0Qfilis5sMlrllzhTooPQzNfVo0+xqhBLe1mXIb6jhTQDIw
YnIU9v3tU3B+lWvymcxJNZEIUv4O3TLRoZhpQNW49paWVHV/lG7vAfaS3M0SE1BJ
bFQdSvrPFo95tkh3HfK/XjF3+kJAAEmpvk/a4uIi9MJEdUXZvkcZtIdIFoerPqs9
iv0GPXlbZxpcgjfI3MNu1Vd6e2TRdUiGat6mNRo5eF1LZhh8u2jPWd6BO0sadn1j
qCz81tBb+gI84ve7hWBQKKRMVAZ4fj4uI+AUL7m5nGhq3RNLZphaeNCB1QhVyfr+
ApsfXTH/LXrq1DI5sbcA9bwGDrcvjnQhz1Rjsjxala32hw0VL7hg0wO3/ZvSvX9C
x99FrspocCNErYJEnQdvemxjF6jOOf0/A96TUsiuLOyLu2C+6u7bH16YzmQs6det
ddqjw7UF/iEEtber9URGJIW26KJa9IAw9IfJOO6/5Ic2MBOgicUk488U12vsG2QY
JWCPsGCbeHIkhfTi0F7s/XBV9ZN7TuZ59hdOt6cJljwjN2Bgh3baCDkqtQjQIMGY
hjCwqTc1R5N4aOt50m5qQEdO/dUACBsMCU3YaeLR+mLRHXGYLGapD47XMBHuz0vc
9Jm232VGhYCrYNi/UYZwuisKZ+LWsfYNWoDdvYGAFjozyXPodLJsNJcGm11QBDkv
HmJse0nrcUay9KG3aQPi3yLbfzjAmBOtIBoIU76RZVAwy0Cxe9eVZ3nCgWuRO1o3
sFz7rMvaA1GGuJ8lZz90td4F4aEXDv3AJBeJSmoFxZL0Xtesvsc2D/+V6HNNTGne
Y+6K3Luwbx91Z9ep0zYB81tjLTJ++fPI80A2SrWvlLp8Ic7GTWYaUqnePGoO/VHg
9RVDpIKpBLBWZLh6DZctOaRn0KZH9vFNbTRnhJXrPMoEnmWsPIwdpG7fJWBiPWre
Egek+CyoURIejf1/RPDszMj5CaefFyOeWJaGa+7kzpZNjJnh6jnb9tnw79ol4yX0
fTOjiHG2FGGgMcm6BkWCJMPXqqeCwh9kx9+wz+OtcE6ZvdK/Rjw5FUAag7Ut7oGR
2XPmWYv2t+0gJVs2UfpS1zKjpXuH+2S4pZP0cbcgqoYKJ+YWls4htld8nMStuEoK
hj19bRsIofB6lhDnEbwi81Y160BIG1eysRmcGvAYsq71EROvVutuiXa0iJEiTxvw
xdNffxjKGPoiVQVpNaZ9vUSTs4bAui7oGtHKrXrGNw9Y8fow28/ndBbw/ZevEvRm
Thy0jPfsTJSBd2VlCRE6naCkzR/Vz6fjT2kgRu9IVfTT79gugjigYnZyqzBRvKDM
9Atlq3E48i/5ZSJxeIeF6mBp0eMIwFEFjWnoADkkTl7Zf/weO9e6x9TJ5sqH/dws
CsxLNAKzW40msgvUQZ5x+3+KEInmtfaYxttwRwbQAq1t+zGl0fxv5KtVFrl9k4mJ
XuCYKk+LsgIOdpH54SNwT3hWOCro8V0ZnrXpih+JTTvlYXQddKUVzh2GjMEcSG5I
wl4mozWPIbawVGB/bDkT4PyX2sZMPBu/yRp69iaeGiQ5rzgs87cGY5MwFqn0oSLP
JTilO9qZtxongt38d2CvRre7fdcBR/SwuuAxCmek66kcd7T76j+afFGM5CQsw7oQ
JFELF7+40Itxyqmn5nS1YSGJC2qvgAk/rdKoS6rXDgQt78tuZN1fT11IWNbcuxI9
O6F+GIbd3+3kF7i4fOmSFaCHTMGfVPNOOUONNCTNGqhwASMvojazauXH1sj4EbCx
arotHW/p6ChYLtoTSPDxelMFsTv1Bcxc3+hKYT/FwR7OsaPZXhdKs8ybdumbI7kZ
sKcrCDWm7qeThM21N9hO1zWZHnzSGCcPRVW/ODJuIYi3UvXLghthRGlqGbOJFnt7
6ARqMnNib8eyso39C0/tTvM0VnF9+7yWb0xqYDSLBgSi4vWRCCI0k+96bgt2SGvc
AbjfV9C7wlY5JM0qXfMnSxPWsCLmhL0ABkU7xgTxzKRZfErLQjHGAW9QkdssuNWv
1Mty6jMnE/g2RmYJRYM4OkU9IxpuTKvLP+FTlTfJRJopSf728s0OdSSLQNHsxG7s
pm6LihNflA0MR7WYXXscqj21VqirQ17Z0PM7uuxW6yXk5LX8hAXkXIXxiHDSK3MM
l92XSArw+V6Lr5trqw6nhKTeTcy9tYCVTIwarrH02/uj27qn6EnJedfJjJY5vgpv
DDPfXfXVTEf/l4IeSNFA5G2RlOe2YIb9GYvR/0xdSGJv0KpVjqYQjHNE/f4f/Ti7
aZkNVmIufT0S32qbNKNNEGfFvU+eB/d8fvQSsERW3jZj5os7+EeTmvdnbjNkrgLE
iJ6Qe+OAMdtPmnsbNkWpqVJx85pNgiTWEkIVUQuPXjxNhUgcD5jBbtKLZTa0QtYn
CQ4Ea2TbHE9wTYtK2zoBTiYN684nlxNfyk8XacV2xdqBUnoFdRO+kk+OnSoTK+XY
b2RNedEtEqryWzPPJSOo/ZetVqXeSjQK3eBJC8yRykA4A6HgZEwTEoxkSg8n1l5j
xdn2Xugc3FZcwHa4TyNIstlHIlJc7lWxj2JMLEQabnXh25Bksv+CeresLC+IgJnS
kuS/JrL9wqY7UdU39g1QkTGUp4ykn7vUEubnlNR0O8ZLSjVX4si60qJLiiSoaY6N
lFv30AwNG/oMA3sqXU9oGNWUzLE/tg8FCXgxE4d3jJtO9RBLOrGw/LGWj8r0fd4g
LhNibJWgXdsUq1XTQIuCnUX3DQMypB8XGW49nhHOIHXf3scdWwVMg6eVsUr1xMMe
z+m6DjI1uW6LZzhdqSmZ5Xyv/6jJ0YbsRtRWjagrVe3OhPUdxy0yTYI8PXMEChyE
TGX7ruRUyfRqZVwi8EePg5ZWUXWMRZN2k8EJwISQZwACAqHKaaTnUQY6XSbV9caz
C+yAJaF9x0XGGOC0WspdeQCa7P02YWq82tJegQ3xgBSUqzUb1h6crQDRu2UDjYci
swejwfO8iJZ9nI+mD64poe4M7ZLDGq05lJGBmEL0Bkeb1xolaE2kYq47xCe3cNee
Sm/E6VwsA//8b0C6hioOD0Ne1L4PIp2x4TSx0UAvzcpwy/+B1R92DM7AvjEkYk6n
rP2GLyiyVnXmAkMkEPa6R+lsiLYHTlztyiRHi+SvEPQIF/3u+HBbGKJqyE8mLr6z
lSl0wXVl8UrtTGVIDloaewDUs1QxfI7FPD8QQvFCASx3Vj7ChByMXZjhtDZQeqqj
DtgZyKbO/DT7US5ZlXtxEhcupMF3Mb3IX4Iz0CRp+UgJ3dW+NZpF9837ApHyQkOm
NPcv48WLcWdYzh7mxd6Rz6NIjf2gRFStyZxqBSDocUsTozc1aJwHlepzoxOTzYwi
o1LmV8Pj7NnLa+y8ZPOCxqO7Yb73x0ugg7ltbauswDCQXyCSOMqhtWOiESUioNhy
ikY7/ANImvHIzKa9qUiq6h+yLyGrevZjvaqd+FfMxxDSJjW3LZdThWOVY9od4Ysk
ZrPH2dw14XH8dKg1iIjFC92eXZYps74Z7tH/bNk79OqEdrTeMsnYyNETxN2lgf9q
LLrFY80Z6NYCNxbsIY9dszPf4EfSPDQC/gTtGy90dTrBeXcgFEJ/Q3EZGu68T80v
dio5O5TsrQLGFIuh6FO/ty2gn0Rs6wevVcid09Sp19IfEBl7YjhEePhWmdS9+TVM
9Teobl7nJ0aUwmKC5MPc+CP33H4KiVL3MPyLWn5aCiciexsiBYQYbCLIZGLKjvn2
U9ByeadavaifixswLFA27e9wASAFt91qobkGlGmy6pWOPesfkZZG/zGg840NWmGz
uzHpUlPlUwgDLFejptWFOEXSiS+1i9HS0H8LbYLDJYKVoEbtrVkcyV/JyxIgbm8M
EiSDpApS0hkq/awnnOB7w2mnH/6sCyvyylNOlHwxAU4awf93nZYG843oF97B5erx
YohBrqtLLuycZs8+8QThIrbNsIfbixjCj9V65toeYxqGf4plAqaf9utKAGSNYj7+
+GzZXZwfUfOq7XjSmy+gL3crTms6AQ8okshSBUBRwTyDtx4kQACsrHD5NFR6AYZN
YHeUFGBW3thAYNziMYyUwKxI1yPfYt/TjqTmB/4EuZUR95OPPm6m/aiFZB/4/Kqs
LbbjkY7aXeXvG4d8lmzDGNHbwOqgdrMpFAwynN0AyVtv/FqXNQMA2pDlB7RzSCl9
wqL3nzgCj/ZyBiGdDZRkZRnGIBOhgr12jvyrM/dc4k6B8ZwOKKFOMBsLYGsAL+0K
9CCkSqt0qxveSr/RYBXlKyjrf/Ytosog44lVwFat2ag8yb09addMzfDdL8W5CJpI
6b5I+KlgVQUhyFjTVU8LLhlAyH30W+6NC0z3/b+1vx7gaRT3j7+2/crySWNIL6I5
KhTgkW0b9U0jd/HbdCsYcdZ2LYY8W65reSyXETksrnLLxoxXxF9g7M+8TtxOa1Tg
1TfoNZheDgmGDy1jyyOeZ7V6BQkeluP4hKztnlhgFFOzEcAg3jDpw/PFmkzqgz+A
f129nkuttqjSBmJWKziTeksCifOixm1HUS/9B/nDFeaAW1P3Ivzf7GYvu7TBbYB/
cEYczoA6M73yIt1Kj6qk34NJFbRpGn2pC5z0CmuWELEI0sJCXXVtrMOgQ5jf/vlN
y0JapUXpms0kBOftns4fnVTAibOueWVpMtjZoIZB9amuAjBGyQ0SO98IjWrI+/ka
WWQzUbAo0CjP31KLdIeCO+4/FDdCZqIztyhoTQaI7hqzVOGULy4YcIqpJqdDZy24
COW78zx2bHOjh9TnMeMfQxvPSQnj6jVLEhGCUppUbl40gLydSdbNgom2hk3zl5Nv
hKxcLBVIZGXK9uWXebKHLmkGtk4RS8bAYsiYJjsErJdrxsn5jaYQTb/g+mntwwOF
KOfGSb8fNPKx78NOcbYPjaPeMj2x1vUbmvwgXuEwWAuAvfFvTPqmsoFEpJs4yPbd
VPYnGEIKBXlzIKcHqhdHM0/tfC8wgLexY6rd7qBJJGscvQDFPRLZeNriBnu+wwkf
5UsyYgcskW5BjFMFwBPxiKeRdq/nmxU0q1RW2tC8RNWvDBYy+3JGde5xqikSC93P
yugYD7atQqmc8F+bWdC7MgO82RJUO6X+35Gw375rXt31/pGFL0qKRiSyoqT30Puo
Yix0fleQxKZptRsiSS5WqSIYxCtbHP/k70t7JoosUDbIHmBIH59ALdWr1sihSrES
fVa9z8oWvEAUeQUc8xH7W6nLGTzGF/vPN5rP9BNCeKQBAU5U5l7vnj8zt9YR45ax
k6E2pwNgnc+4RLD+oem44IY6FZ4UY/1SmN5dpAeZmUvGvayt9Qw/h1ykQla4wqoj
PA070QOcRkEeLvz/CHfKg4fT7HMSnY0u55WHqkSF7Wkd2U9AVvzn7A85lF0+xc7f
pdu9fEbhGgE9nrbZNljIOxM8+jXjcy+jkSJEd1saMf3w7qzNCL54KLyA9gUcn/fc
s8KVOSPc86hq61XHFvMvocX0AINPySs9ZSXRmGgFyo4mV58v/zq/9stVbL9Z5Fsh
IC3fsd1c+70IAxCAtDBruGZ8Zbqq/9qapSHXEjZnn2m0fLilv5533rGiZq86yVrb
Vpx2bV719kFZl4zIK1CgrUe1j6+xTbFIYKldYf29+NWnRRDAUO+sZE/6BMl5hCmf
sQtu5xM0EflzB1ElNHHqrKAgNbET79emE8wDD/odspxZ9GRHcYzgq3ZDRUMQ9K+T
xqQJ3CbRQRCC8kDKEzeqwbB5YGV7aVuTuP8msagpnj317UDVqEequjwqtFVxJ0eq
lrUQ1zhRZpaGtMXj7OrMdwyzIKyDEEhcOBXCQldEnKgwAwY/5hLh3TrlbIHsPMvB
uv5Dp5/wxm80g0jnJ8T1cX61apx1TnY0fUCIBZmkuC/6iiplsezpDsYuZhr8SRBU
K4kGOrp5HBLGBbck70DQIdLVm75OAiSEnU7zCo+4XoGmojd5YWt5a+vyf2Dg/d5N
qByP99qy000O6jRi1mnnvPYQW9oZ/2cr47qsekO6CD2kV6NV+pBWcdUB8+I/+jui
NdI8gbgxI3WRWbYj0k3EL828miUzhr5Hb4USi+0tdZ0OpOd5pdOXhK329/VsKSyo
gGXZtTiBAk1qB+nLPlvS6H4JTYIwj+omAtFij7iJFriStJmHWdXoLzm2bm8bLCfj
Qr+3FCEvdHlg2U3pFAW+4XSkbr5SrMkPCIR1PLn2O6bABNIvLIFlGyHwvUAdyEXf
oZn0cdyO006cRCpBtxEMenxIzrJNRru2mjJtAvtaRAqINelYR+7VprPNOHA/ldMy
OlUEZeFUSYa9F8pjIDmvKU65zPTJDZHMuvcBQa9woM8bPK7Xnjb4IKs6u5YVzInv
is8TEKTHqKilGYWGTkwNlw6wSVPVACXDfm/edJ7q1XhTAG/69IuYK6BdmIo4Otha
oxhOLWQ5rxnS/GpF0HVREvxl8tYWu9gViIdD/6zh0sjA5ITEdqXfrYeTjcrMlWKR
jozhQzhD+FhSoR/K13BthszTxmThkNTslpvgy16qQmRmyrgPqytMg0+vK5vvIySe
jnJRSrE66ST8pUUsM3rB60PtqmDQnXvSyshhvEamnB+aOYQ1Qj4tQ7rV5x7KtQE8
N7iLdYkiDv4a3JgdAKPZjgj6Ds+IpDMoEnjhY/WL2eaZojBvXKxrwzafqP+I6YTi
sUn568cn+di2c183QtehbEjxcLc0HkPlBxkgUdCEzquho8lKl/AI3QMmhuVqvbgI
zhn8+C5OUvVJG6O725v/JUVorL6kum61oh+VqF+kQPEmqREzvezByeFOjwShDjLX
VpYpg7uxvikxDFlQYlM4cSV+McuUYf55elm1acmsn//8tj96UzAJLqeOMKy3nPgc
XKPF63svl16q9YwpN4GzMS7NyWSh+15UuqDwkIhaq/Knt2NX+2W9smSGnreWEBOn
TM+ex8zk2lfK8VJm2tSkqmHKCWnUcZqGuJUsMkbXhdtGP8/qXkGObkwuHTSdboO+
c0JdSj/N5GBGjGYGS/dWVMI9GF4Iaflfyh0vLFN0BG0rCa2mvC0iKSXRwiAFllEE
Ag3YNFEtA+LEUmQ7DGAzwGwgfV0IJuYSAFL0OxE50E3i0vzERj2nlLoEyqZrXSfO
UyoiKdvkdz2jG3/HGsii5XbmOUctFZMRYp9LJXU8AMTv9dlvCD/bEvASiVezFKhW
qzciVLtKgfiJaesTbXZNA823aFidonZf9m9Wv2ZPGfeiAqNUTXBc/+6FrvkEj6PP
GZgT62n99bHp3R1RpRvNLcj6O3TRtY0XbVE5ZdDPbXXhrUnzux2JdFgWCv0C5uEz
hs03Md0bi57Zm3ZHNyhrkQlNs6RnrMYBdOnKyyBcghBN2QpPMO6vgHPgNmBddGwD
riVMk0AlsmJsIotdphwbTA+GEmJrBtzn3J7hdXG+kHCIN0wdy0DNOZXOhWCP2epO
nhga+Hdim6FdnEweuNmScz0mNggpaRulSYuzLyCEYkv09CP1ycrnSycLnzCVJTv4
vU3jNCP6hccNO6LCSpOQmXOR2cDQl5O6FM7cdeCWY3gxNDt2Y8MlfIyXgXC21KHD
RhgE/1LtRzryN3ppWZ67UUJx56Qx6GsRGDd4zgi1sDkJAuBwE7Q0MCJbTuiCJP6k
EjEYrBS/76guZ9q4UMiFkJL+EoxlMJeZ2tVGsPPD1kTMmgrgdPOn486H64xbZ81s
8bJ7+VHQmgWdU5xqSZ/jM2W3y5nCi3viJb74ZNvUSEzUmwWXZCf2aLjF7XercTM4
wHUtjA/b4iV9Bp22894H8fWnVz9fsFVZvbnyCWOaXrkmqKLha/ErdxhCszvI44OH
fMfhoPxnlIjZmXGU2OZwOQNX5FAvlokGplLLPeoFsDwFHSRwa7KaPBMcESxlQAsE
7XUyFwcyjK67ZIkgcVSI5X4ZDpreJVwe5PGUE4Wv8YyvEdkUzjMojhHpSUrdOmX4
WCVTy2A72Vb4MKPpAOnv2/i/xvwsVVBRZbYpZid6HKTfG4ex6q7PxfUgUHCskUmx
HWOtwTuY6tF/Bk9VGv5gNrAuUaHfVuqX0gnJolXWSMgGBkyjimPrcAScKtEjdaVN
8qXwuAM0qdAxH4AcVwfMTI0DZGrVvY3sZ91xYowAAV246fEt1bzW/216t2chmDFk
pK3qe9SuPPBHfz+mAe00FW4ZRsBwLMON9/pM4BJJhp6EmR6G8gpRg3KZmFLEiqN2
pJAz8vXWHqPVE9aRRA4UeAavNAA81zB2bgZccUINWxIrBKAvePmrdW1bnldaMGWZ
si9hEhBqxFRi93eV7gu/qDC4k6sstCVXbj1JZXJBTkclrh0MalzOPsM5BpDb9Hcv
IlpdsiGBu7DjT4gXyqpFGWimvzhJfshkYwZ/31VfeFCEpH1x2OcQ+zIP86jpJOHN
feU6mDeMIsdrhA5BGGCwdIB8q7sRHuWkSiFrd7Cxd8AHvb0MwUY8SWssgU5YEmwI
j36KlsyzofUTVpUbcmMm1uztd02PjMBA+4HVWS/IKVmq3ABKoZFCUTjHL4+vqXJy
6aCxwAobC23Yo5dfJ0TFUuFZuM/Xh+INg6ELcisJ9g/Dr94wG/ETMGs8k8bmJpR/
8pSaE4IPO09i12LDzjJ+U0dedUXe4ZHIFpaRBupTnNfhkD366GALZh/lUKpPRtPH
YOQFjeUcBtkD2aN32CSZRKNA913RLxOuV8td7c1PFJAUhHHd2FgMf1/lGrxPaD+q
Q45JqR2HQ4vqs/uXiNhKOMudkrJ53OZZDhj/DrEHvUTnF9mYY1z25UDAzD+1otls
cozbj0xTqpYL4kaCIMj9v0B45d4EHCEP7DwX//NjQso8kcpqdH/xZDqFG2jh3TEy
To7qNMjEwkPFpC3iKK6S55xUH3qm2TyzFJ6aQWb7ds8Eg7kGLVHOmiaIm8KTqx3r
NOZMkXC6JQmBQ8HJoZ8sY9J85Wuu0YVxLs7m8pcII7E9O4/QqZKFXyMVJqBj6kVv
i8L2LTYhl7XawjrDGHjzqn7fmBtqCObYJS6NJZGfKE8chqvADhrf6BRr7W0P5cWS
F97NP4Th2CxFHMtnCNxOin6GCzq9zUzkwiwOT+f2rV/ENV/OWuY3zHFbu7mhIO48
m1GcaEId42p3Du1wPnxR0ihbJFyAQ7jn0fQDCh+2Q3sYB4/HKFhQZA3FfsgCKSCD
oJQwsfm2ghDzhTtnEFdsRmb3+JwynC8YSC+hw5MlXphsK+aBkUMD0HJv3MwAwsH1
h4WzUQ4Aant2AOVr4g4sLL0jKpe5moPoSBSOjcx9jPTDXKQE/zbuVCMaKFYL9bLD
Zz+sb01z36aMbWVGBxx/dDHXhTl15/WD/xU50qvVlAYNSxM4hLEVX0SOk4p7pKFB
O+l7sAKtzAJ3k9YFeIBeD2J8pArRAc446yHGWke9U/nJI7IYs4HDUuLpp7YUYF+R
6eD/Uy9/RF0C3qcHNrgZYWdHqtu4jRcDTQZ49qaQFCYhbUax5G3AIk7QM5DzkkT2
OOSdL2CFGke1rqX3ZSV8fJG2lek2LGDATXC8cGsbh/RHWZK9eMo4W4PqjUEl59uL
pNLMXt9TPFV+EEcaxyJS+K0Kxeu9E4kbbQr9d4QvwvpyGeRuQyOVqQibkTB4BtMl
mswC2Wrf+Uq6ZZqvMPyS/JBa4YvPs1M1W6L7Qnc/xx0SRF4dKs0tHnNN0nBLN9W0
NSLHZPEKe7qljCfvj7nNienIjEuibgi9yHePcOhnryeDiH2upHR3SbhmXtsXDKjS
tjihe5yEj7SY2lsuWf0qxPX6ssy6bqHNjS94kHrDLGSbsZ1TClKaAYQtuI+QXrtt
48ujs+4WpQALhvyX3x5jCFrQhQkmKJUF7tYXHN2+73HKOCsaNhV0IQtfrRACCOmC
V4Ge3b7PftZwsc07YXzdCgfuns5LAL0+DCZvF3CO/UpJQQMVn8CeZIGwwBsV0PwM
h7VL31fsP5zuwbyNsq7z2Q6AFzOxlvcSsCMELZgTG1N6LYm9lZ1cpXi57TQGuxS/
lUwRy/X+nJ1iFVPkYe/o+zI3qARAyJjqc9ir/nw3BmaFP6m6qaIIkz+yVVRshwVE
wvHYtLb4pMsMsHpLwOz+cJp4AZ2VizVQHORqbfueAot7/rjNX2HYTeXVcLR+ymit
q9UqnBxB006uhjOGLQ8f6hhQL1BRfSa0CuEkirN1iZuE9kPPQpdlrPCz4EhqH2If
1SrR/VVE5Ihvll5Qe7jAg8MzvSzTnI+4/d5JuERh8Al+ytOXWYvXeoO0/HvzLSh3
b+daIk6uw5AfXS8TzF5fP8y2eeEkADBjXUfGnczF1HAybyVakMjHsWvAKU5gkWkD
xxjbqg6e0wvMjjMwj5Q4a2kcgenv02R/cIrW2psJ4PVZpWdJbSTq9dY9ePqePNeZ
LOd4OTG/MXXlXUc9tNRx2KTeRUh0MAjHtHCzBKi8nizbyxUNedsG9pnO1Gsbg7kk
/IdyqRv8E3bxghcw1QWSKBhBpe9QPsL+dSf9rhn+/RWTCZXLaLjYWJcds3Qsd285
mMRwcqxqWeSi8t3Tb2TeVj8QfSMV8yy+E5F6Yyx6bo3GYVGip9xlclKwGl9zBERi
yb8GowdesIxc1pCiwYQ345kJtaB53nHrsj2RWPVBMriQGn1E7pRJq/ZoQyyaEViS
VFK547NSmHxLrjKMTprfnXjWO+XXfZAFKySOyx/tTBkr33OKuIObXhCacgHWpIdS
rMi7mT4zezxXz98U5uhZt58IUXm23SC+nXUVdFrhP3oloHqymSDrllGm/84Vtw02
+QaRzSI6mVO8MKjEHYj9uYhZqFzuoK9rdCCfusRzutpyIhS2pott7IZDX0IYImMj
97p87F9h4zH2vWtxk2/aNSvWXKf3MD5U/LW14pIwx4/js7OBi3YNrOGnmyLgbvTE
N4lN2CgAdIBgHAsyc8YStCaEJ6ImzHZWKUS4S15GXqFBInrQFuNQ2deLxFNJv5bP
+5a/kPwvfvjr+DD4/LKjfqkhU3vg3kjxGzQRWUuEHYjSSRNGgGBTtX+6XNPhRAQ2
Q1WkNvb/65yzjmzD0uKftzj1cZgrAdH1s8aqwGLrlrABUOtjPlwq8PNEa8Llz0Nt
kyu4nxpqOKpU8wJ5ODzQEhAIhBi60YfuNS2oRsEUXk2NcvhR2ngNPITPxo7x0kU0
ZbBjtbOWvPqkn23gw4U0FbidNMzkl4ZarTTTISbJ7YtVeaeDPfRTflhbDiCv/CFP
4tYMAtkwHjxApxzXOtLMXfCTosZGGqKvg6SGrsr87+jXUhG2seyKPy5iSRNTMOml
+atpl11d5Tu2W3EJ+ii+Mh3toONkoiTmIq+1Q11ugunj+9zS0JAdJbwY3NUI8Egs
GpAv520XCACj2xQvFZ+KFpiuqm+c+sKSf2UlQrHM/IavZGoN5LYqkKTJ6vIe9KKT
g0N0ovCWdyM5SGvtggAJE4r/u79z8uUHpPRPfkIZjUJSOWP+w9UfCtLR+GeU5r8J
atab+F0gVRyMIvoBa0MC7XNIwhMZwo2vsFARFpPJQc+WfQwqlCFckPa2JxXGpTLX
tCQc8rgRFFkgIhEuqWLpN0ao98ZAscdfQLSb39R0rZQarwLCyp8d+8EiA99VbNTM
ebF2WThlyt+aZjy+mmoWrTfgnUO3T0FJn76JK4EyhcWCJcbxlUfcPzexqSrVqUO1
D4+Fs0BjgvrT7B8nP6Tke/DbiaUvhO+iGkiJDN083LTbXefPYHwMusJGDQe/1tPU
nbJiUoccClqkbPdI6b6L+YBJ/gbs5QznOzh6r7eyLrr3WUVVHfNiAGPP3wP+uyTN
TwwngL47kMkyhryKtxS9aFDfGSutPLzuFpPC+HFEOq5af6D4G2m90Zj81Ibbdjfr
JGHEGE95XgVOQkf7H+RpBDiIna0y6UhE6khQId470IGIRYpxOlXQCyi/ljU0dcN2
FJJgr+Dys3z9BfH1Bksw1ATNBpU+HaJ5qQFB2U3AOjnvc+N/1MpYboTnmjhBUYJX
bd1FWwebfSopnRR6xNqaZy3zjg75oTCDC0kT0gWBHPVlH488rNCcFh8kFBwGdf6m
gDEpWtshQpL4YLGMwACUGmJZwyBuvGZWJpwiwyRQj2d5vIAifCxqjirMoJ+eZrg8
K5VtW7P3JCE2Lk4LchM+0GFmG2w34TnUMjfNvFtnQewdfQwHfaNkhu0bcx8C0fYM
kJYbsHXgbYXL48GpAYXPlTelGJshSGLot5SIZwjmBPR9e3pNYwQLBRvIuVCjUELH
ZDZY9CPy7rBAgcGGGE4cDjDWkZR/5749i6U9WpxHyAx6lnI63I3qxGpc9Pg/vq0W
E+HFg2mqxwZQrS+tV3nXugvhSXr3euMpxgBTx0Nz8LS0pihdebuSCqjmrVJd2Ipa
1/n3sBvjAs3pzgjuvtme5nlRsH9lWbqCMkv3k+BlYvXrtqEc7CLxcYdHa6IuPw2l
afhwUc06tRPIOef1xFmwuUSH9FXe48Mmxa48srrQi15F9xuqFSLhZ39ILGhdOEVw
z3W5Y9MTpGLnI5R1janrHqBIYAxlVoj7nHc6+s6rNupUW/FFAdKtATbVHyCgWb9o
IZfrs1FMM9mTSpa6WQqENWlB3BJysu1B++MT9h2wkIQCqiwM/O/ilpz64f3HNY4m
+xJp4fgvui7t98/84ae9cL6ZNwhwYyZL1BcRyD7giolLWQFTDxkWGbyotnul7luq
4Im4xd6iR3usXtxBOzfx1Mbpsb4JjEgnF2cayFHdxgnhH7ZDgTu/svEIxv7E15q4
QtuoU0cdMX2tBlnHYo4DiFcfYcorqw+h7LFZmSNylDS/4x0JjyZyPtXQvR6tozM4
/ccTQf6thioPNsnt7lAmO8RSIg3e9fS5WWFwGBI2gGC+c5WNqbQso3+FyURCZOAA
EjLcxMU2QuQRFrg7LM90OvBNuEtfW84gtXz0kgDaEQH+vg+RjcjO60GhAH4OW2Ph
1rT1xisjgyCKaz1wP7dPy0pIzfnMcfj595FhpUBk8IXTLpMWAx1QB7uY0NKOsCL5
mDf7INk3a7f8qmv8E/Qk1ZoNTnk1+W9NvWS5mZmJVLiPjsUTzAAeSWVdayGo82Gm
rgAa2xP2GzSTWJTmoIJqP+Vhftq7uTGGBouJT4M05MEoGz6pU5d9Fqe64mVd3rCX
MNAg3IPLLRTXyWr95I9MGiNZbZT6qSsiHokw8CgB9E7dL0xJA+dIanKEul1B4QD9
VtyMM5o3NVcl8mXfyRUpssBBkdQqYbnAu5cWf5jP/GBup4EikrisuWwnwpL0NILO
90Y5XETpb4/1f6Br3p8EziA95tHYchzAn7ro4JN6u/8X5ux966pT15fNeCgFS36h
SI3IjZh2d9ClkhQwDYsRAgkvPKzfE66YKZjgc1Qu4nBSwMAH5zcCuoSBVzOaAVjQ
RBwIhdCQndgePL5VdX3OuMYx7sm3UUiqM6YIcdcFBNtCRfPor+S6wsueSwyGHBBl
p2lMliaUECCyYqJxcI2ENS//9+bfM5eePKuTN5yKoIi5nhnTGZHhFY64a/pX9/h+
lYXAs8wNBi93uY2IGMsJIQIufhTPUk6nUrXvFBUUrbLGbnenZd1oIAxGQjDQhvu4
2HDYADn1sl2xofAjwj1U0l8FIth/FH0frHv03y06i6CGZAiEssHslM2+LLWuhb+X
4VPS6f2LBHcPDcvJID4/kUYVCMViGARyVhf/zdZ2Yj8C+umeN6TVeJ1TAppBM260
EQEv+J5DzN2AQop/K/UkC2e/5jPX1x4gPkFc2q1Bp+2MZPBeLzdv67ZoOW8ASb+y
QwGPEbxnal/OEBsbo0hjcf7DUnbueQdwJBY9nvPgbXsS64+oyhRy1McYoOBxS4v1
hoME2Ts177ROhsIRqIwJKB6cWD/qQdKW3Ql45BfxK07Uy99HuIe9T7sRbmtcnc9T
2lnugYeR8iiWdXT7aM+xImSNYtenCwY3hTpceqyiw3HjZX8r8pUUGXE6jP1KTfb5
hE8zF5iJM/Cm/mge0oe3M8Tkn3MX1nnPfDfsBbidQnaI9aZ4bfZym8SSEoEe5bqo
w0HKOEw66bWRXudZJbF7fW3pD5P7dHOqDvzRiKYgryCelRaiFwN4BaBJlC6BQxst
OFPc6YG3flecynrSZLXB1DZkqCXyZ5q3xYOi+8ipiLoZRp7/1BO4LuSY4NJsMe0Z
3Xz1ynkkaGquwz6H2ccS1MeW9iWNGoDInNsxDbWe/oOtP+sKDzfuCvGd5i/nAaBN
I3CwJnSC1qBtTo40vziXD+cm3sNnOlinDdK0VZA7SN1cJEwv79gtUlc7/3xMjf1s
TEpkk6/N6kZScjAyfBefTYy4r067JoFdWBME+nMhl6LgpCPkCof4NQRmXVVDF8FC
per5YOhUd6NIm/PyOcEZJXDPNCI0m5KmSkLBRy3R8h1dDT4mxXla5TgTBrzg3XNs
CK6UhN9u3bfA2EI7f4qdzYuoMu6rVBq2rbHNHbPMcjSXbz+5OO59XWWv52v1d64Y
2DjjS0pn8BWlXAL3mnx2dDh1ISCIBwGF7sCdq83S6BUEt+bYR1/xYhJhm0FgDheV
6/iAcBdgLHfbu0y38cUJHWZ9xZgH+2JpFCs5DYxYrn8YwfkITOgMUJD3y7OL+f9t
O3RSXwHSgJ0vGv+BpP2byg7pxVxGqN7pIzD/uji06GzK0O99xMhThnxUyIQrmEBX
mI8H09UGYvjPZOJWl68dP8VWBNjD4DMk0k0P9zIQBX77IN21/xOT2mE8wPHTKYsA
WEqYPbAJwAlyqwbkGTdvHCzmEJCgjhIN8ormj+1lBrQrgpD2Ceo42EvnSjcEVTOL
vqZjmfOPynRgAoBLADDVfhrBB+JNQbXS0pJGG3NYqgcTZGzD+hjBFD8q1z3gCfFf
tmjA25krZBbm5OWIbj7zJxlVikLcbgMW8ABD0EsBVlUbxNdZwYRRNzl0v8AQnDHW
wBAxp7mzST3IEc/8uBiAaB3rSrEbFXGQ/fyYtO5Y7VZqQWgrPwf4u6BkL2nrHmxd
je5ySiQF0309T73/dLuuHgImHGcDBS8h2dWwnOh20GqA4uSbUJiXSujVY6Ww1J2U
88/EWL//Rwy1sqYUjP4HGg2DFc1qCDWI0kIWlukthX+8nDzYquWsjUEWOm5ueJVf
EIBqzRkA+wNMZY/Afz/BmfuRVMEY8i0oYnCzkhIHrq0qz47zBKvp44tz9Ilv0yVg
YGwvfunwkF5ZjH1yMg8Y+1xHUdEAsepNWPgZFlitgJSeA1doclEuJYv34TEJFF0c
C5oa1gpmdYUSMyNooi4Ezp0f6Ubnef8Mynq6+JaO5nCkLDSGnd1uWcwHbh1vWC/n
/692+cLoDVAx03Rg57akLKBFJP7VSf6hPmrehPSxFjjB+iWJ5phYpb5wVNWD7+f2
E90ULYq6vziemrvRyBck6ntB3I/s/KRtRP5X9wcL1jPYsZS+3jjEqULTXJuD2Ay3
UGqiyVnRpZS04RofYbeO94SFn8n1VjkfyPhiYdltpVqYAaN+rjarD06weca5no92
eC/09oiziQP5lH+xWQp4UpZ4szuDnAmI15Qc8+CCN4/1LHajUHH/S3Ip+YFU2S2o
GGfNzA/Hf17LeUOoPOnPTE+CjZHnUQf20OiihTL5LQ8YkqQzwlShfeQ+ygLCJDu5
jMzfFD1B0x39hy1/OnRJHivX7ViC6Nd0TA60Gzthb49IsZqJtSgwkITYCaP0t0T8
HrvOkL9Xrqx3y9HzMeldHuaTLLeAfeTh2o2QTX26sJ1kHD1qvZUEMW66r8vU/8XK
Or8AkV/7iAb7shZNqL2Hojk0LONwj9Ouv1tLWiS+I243wcPb6/5MGLy/f7AelRwm
u3/PVf3bjoMz3wxjKTif/WsmB/ftsmos7MokmDsB9yKS4zCEePeMQyX537T9WHT9
5lfPlhYWu2GXBBRfBO5MhTWt8roXit5SR9fj7votMNDRcbIa0ptcm3rBlZVZ/ifd
4AMshmnkWcn+YBBMU9c69LGOFhnQLxqAWrmsU1K776kgrqaPqNwB/dbnUlmel2Wn
7GomuuMNxS91i4PXBTclY139z3B7qguJc64GrrE6P99esdThJLfzT3Z9EdwUlzRd
QwLBsmGiP9bVGRXj8aLH4tC5Jld2tmQyaWVOylPXie73wf1JfHHPjz6x6yq3Q6MW
nc8ciwgSDxz3vytKqJ0osELUPozMjswJtWH/RsHFcnOvkKcp3xO7J5XQBgLtG+vJ
PCXgy4inf4o96KnrEpdaSxWD7yVhqNyqZVmkuXjjV60Tw4Yw6ue32LdIpyTFysxG
Qlp2dQwcghnDhJ82BH5JVGAI4ghDqnn2J3qzqOAPp/cEqX5oyQ/ONqrSLUG6JBSr
bRG/3DG0N4mq/1TXe92VbnO7BhIFQn4958w04kJgppE5VYDW76ktCfFzgNyGF72y
SfjYAXIIdpC9JDalLJGfTGZr6gpmpx8hdgb5B8vjBmHvdaftHz4J/KZxRRcOrXO0
zBSnjh2RpWMVBTIv/H4r8sLGIPZid82fE3yA2D3Ek+MS9uN+VZLT+D2eggdcrcDk
+e/iTWX+9S+xCZv0AOuGF0Svbvp1HaER6pMw+v1BWr/0Lq00AqEEmPHyazQeYHSJ
vXpse8A9q0lP6iUnXnZBD9CnOfK9ePtU7clvUJZCsGWdeEp6DGG+6kihYJFyByOs
/sqBUiGKSrPUgT04RKuoQgMHCjXY+xeS3lBeX2b4fVB0YLh1JTFdtZuMgHB36J94
NKwFirv5vYUlK+qoag4Ep6R7oQ6Ijs8Pmf5jwXV+ASmOCdKSZpGVEDar+zhKFdb9
et7JAPk5k+qeSfl6OsP5Qg4x30CoCZ0YhFHpLRKeeWN1WLSGQRD0t+AhAVlz1UR+
8Nwl5slboDARahuqmr7U1UnlqTVSRjRj+j8BBBl9AFfjoFFppdtVHyzGvJbGRhAv
I/KHczbKL1A1yoaxzbqr6lVjtsVJ1ujhtBsTORbu2ye68isp/RleRa1lwDNeZEbK
p0VFudMmDgSpsbhYRVV9uLaL7RKknflSr916DDb2GJlGgTxtu7a8IWKiVIEJfNde
xhXbz6IR3GjA1dZ716XLeacYlb8M3DNRUzcsfFrByPU16PCqq/SAOMnO+VN9pN5J
c1Y+Bh0sQX8rfeu4wuUTVBJLoEjwR4vE3F/m0wPwhadNcEnlILT0nX4MoBlMgTL0
4SDJkN1xJb8terS+xTnf0rHHJ6II11447pE9pnHyM0RdYWN1O2FK2ymTxYLFFBob
XXt/6rLi1mWSBIu3q0fhQ0CvBNIGadVuhpYQIW+QkvdAmRlBWemN7xuzu1CBfP7O
m0goKvBxHaGCleQUHxPoC0rE8i4pyymTPxzNcEOPQ936d1BsRstwzCfJ0V+ZkJ6K
3szbKOa8qxCUAu8umQpfm5GrDjTSfepWfjPq7qvsEbaUltzESXH1NV3xLR/fwEv9
PTXTXOLBaXA9PrDbKK5ZMLAdXYj3bAM0R5E3o78SaR5KnfjHBuTspO756rI783H/
HMvWg1vAMZSg84aND6o5DZSn0UD7xfsyALhBoit1zFR45ekS4uEpxrdwEuLf7Y/r
D5FmLKhWQx1iqAVtLIv8IX6vHaqWXShXA5sSLb7wNhOWs85zA6z2zq9lpef0L8h4
RJYHEBaZNvr1YwzXbLBnnzc//Epd4uqwjMFno2FE1qkLFOtAvK0PXfPZoFL/W8ly
+DFx3Naqay890d56E/UNwDiHQUBYMQ9ZCpd1WdzkRv1MohPfMfo4LoikZa7VZxWz
91rGvXmmWQc41eDQyBPDH5nMl0NHlLp3jsTFnqFmYvTkruVMocBJwZtINeSe9/9T
nQT3CZM/ohe+OtgVr4GQ8GpkgsObSDmk5VBdwBhE9PSnlfbB2JG52U/OV9VKJ/B/
KPxg9hDUzw4RMX5WXwX7dieojTcy5AcBazkmy/wLfMN11ISrxKGEwAYhyC8BIGdd
yqwUEYXNCIO6n4uimnKUGT17jayFSHj8MU7Ue+QfWzlFlXh+AdZFzKtu6F3fAtbI
eTvoMMw02UoxO7O33jnrq5bZ1g+mKl6QC7Sbl02U1T62KCT4c3K8HZ8V4deSsyAd
FzyE7lvzl3S84Nn9jNb6weHrmrqdKno7Qj/MYpTrPORM2Ws8r5xFBw2YHqEskv6E
mi4SPcnaWjhGT9DGrzn2pUktaegyW/FmiuOlKx+hvOSS6rd8veG7V7IgpPQgsGNZ
qFme8AiYr7WiDeJ1X+iacQ+yvbc/UN7MDdjuYVXYxCaopkUrZ8ugbkSLTLsi4yay
3AigV80mpBOyzYYj94JZuEOqInYWGzIsTWZpSZezluGekDSfyHBmkLgtg4wCFNkK
i0ffT1koWPRaoAMBYNbOjCmRF2NElG9OQjCQITyBdap3D7FfsnIDW1Zj2JocI45z
T5JA0ytUgffe8+5BaQiKmwxZXKv/U+qcXp0f0+UIB6bzgebPP3mSDdhesneFNZoP
wfxwD/Kf6OfXU3xjutBWX25Nel8k6372WByUfES55dJOTJfj523H3yswaUBVYihc
vNewVb10khBpRb+nzj1i66YnMyufToJ9ykJBM09SJCIpyn1PSwvh/UGAGvnvLcoo
iGWFJDXgtHFKpwHpSrjF9/RwZp8dvDiEbAjYFE7khdi99b+Uz5o4BVP8LUhOThBh
FCc+l2JwZE8GQ2eHF5kb8PR3yHMsJj23zcRs32Q1F0vpOwbNx2bsxSQEBlGds4HD
yzdPu6iqHcIAL98GyI5tcdBJstFT/33IqcdNccOrOHdOqqhJVffZolXEEUaXbcFr
txRo0eiM3vp9V8k+3Vj4dtbngCwdHq5byk32pudza0asM9tkYa1+4Nbs6amrZsBC
WfJFfEQf5ykRdzFioN4PD8aZO81K/h8+YBNFlgHtWdSHW2fv78w6CwkPkd5SE6O9
mCMOL4lJBF/Yb3EKzDaDpvJa8b6YRDXjbxQoJCOJCda+RISvp5wG8j1I9TtsXKg4
kl1yWd3CiADfmipDwg81uUfCN0wgGNTTxaL5JUGV7l8EkLZb3TSzDTp8c+2QtqAP
JXPnfdM81FPVCSyokD5LKnMcvX5fRrWfeGpnt4tvzjBt+1ypFYQ86s4uSUfG/Fsx
6J3H1TaQCzdN8oTy58+CZ+NmmHsLAl1UVe3xmG39Cn3WUZY8WX9BUaNwIwi4zW4i
4/K2JvWOlQxdamcrff9N12c2x6GvCzuPI20Q19Wa6Km58S1bhIEMMjjkSPsUMExa
4tnrEzkTgsyC08Nvre4zwRmp0TEKXW5fu33VrpttQqsuYLmSj+Wj6cVB3gwFArh1
Zd4IWBQANXxvYr6BnOLs7lqWKPh5GfzMyWLdrgjhPjymw+iLvVPnUr9pcyw5srXV
+yd/PllIWs0S9Mg/8o5xhKhNYH+ezqYyWZKWaPQ1frAwAbZwy6cP4YfuajIRwN+S
8AHBJdbLKW2S/ybYOwn/Gd+VJh2oZszIXE4U9g/mJ9ewlMPycn2n1lmPqyekfHHH
5D+3KX35Iizfe4T6dEraXik7rHqWU+8jkX8NCDl3ZB2h/4XPuCEhG+d+K5DM/EJK
++/nwjmgEK80xKZRXKCr3IwizSPso+bdRco8AcyzRXZ69qA1Ql0aaaxr0D0j7m3N
OXnOhZdcv6L9fOi/cu44fVSCmpKAeR3FaDr2cSWiqx9fpL0v5lokcmr7YpiKWZp1
p72+ul/5berE37Y+dBpFlDlHaQORMtiYQF7qLDb2WtPjmkVhok7xq1XCzjexgpZd
SS8O9iBN07fLPTAsl0RfQgmv4jv4ez8pe+SHRHyg9p5DUyrl+K/HNym7sjnEgtaY
GvmUIiBSEDn2E/Ow7OpVFUqye85k/9ONjKkkxY9XElyaJvqir/WcvrkI330YJXUh
QMFvGB+hq4W7xXpfzLNR0wV4m5nGzL4UqOqW0PBHytAp3F9Ncj4ngfwKl2O5cEQw
dxENq+ZIJ+u/0q2vWN7paCH7JwRag7G9lzHHmwqULRoZX0O7IZFPXjZGgrIO4lQt
T3FZih2+qqQdq0v/0QUVtGHf33M1fTY9gPmNxVsoDAfuYCXXwxx/lU2K/3ri5i7y
dAJ9cqEkpUo6ycyLwWCLqwcnUeASkvWox2r5r2AKbkFrnAA/pBPAHTkZkcRhm8P2
1vvlySvlHdquhUxX8T86ROg8Air/L8cwvmB1KiGcfhYfmTcMJFXB9PFaX2ebdQFc
HFUds7BV49iwk+0SzIBVk7pGrivQSB7pH3IABlJk7oFLuMVGvx3ym5XDHvaQ33sT
FeC5hEwfrQNWfY6rLc6kHo4Q6SfiiBLALRfvs52BBbeFbBNb2OVCa6SII8gbYZ+q
Q5VFMuNCtbbAMdMXB+1jhruJnjwb44sjExCZDnm6X3KnEwjZVL8HIslGvPJDRE1S
ZfPuqxi6FBsq1lmJpqY5Vlr5bLzjn+CnTIpQauK7qIFlktsyvRwIK/Qj5pIQbKq7
qp87kFRU3cGSoxHy+1eWtL+JtiiTTW/hDAxPZBTj8xpSjgvXPFBb9o8KcRnT7DBi
eMDTr02ftwgWryd2aA7pIkUHQingdkgIFT3yjTirDKLmgIPjhDYQFKGNjRKSets4
zQH1n/gRwfl/o8uTaiKy2hvC8DmELnHJ8p/lox0yedY1iclmLz5PwJxCKi28p9YP
AbF9v/lDjx05LQi2qNCetiUecXFKGC4blrM626DNLifO/W8HTBFnFOeTMCbqQItL
pw9iumA1fYJrsvxwi/Cu+QWRaNqfSG/vZeRKldBM7gajgKpbf62v/QRMb/O8/bM/
LOV3xd0XhN8XmEzGEwWAkrMrsp98eoll8BqFjDArPaYlXOGGWCqD9YcV7ApiN0r6
43PBij+UjQ/z36xH8v7MN1WOchKsywM9a+vVQvhIVBDG5wHF3MggXhW/NA019z2d
wUJx2EQESbBu538vjvfJNEWYiSTFhI3tEQRVDI5m0JM+pqwLq3vh4a/XYDTF1GIr
sX1DsJIA6WQ9CzRa6GwMUuoho9wgA+qIoXnxK7F++ughY5YatU8X8UU1EG6OPDbZ
OmQpFZaZBwIopWxJ4MDmMt14jmyMUChgyOe9gymbvcG2GUF7eYepgcOdPJJpq40l
8yiIpGMoJNcUwQk4x80vIXHacoTvGLur7n5i61gtn0qU6Xjku6/6CDSI8RBrlmte
9eskDJ9EEojxSAR8JxvU3vJNcVbi4dl87XYXh+Ec95JOXQBEFnkJ63tJdqfQmEm3
dg553tx5KEPfXKlFNTaFMYvHaUIc7KdKwVoB/u+bN5pWdWAxKH3NfSDb1G349YaT
X0qj2LhsSdnvmdGXbARFa91e5feHClWrudwHT2jGQv7zlH6dngM90UWs1cgoF141
YshYifUpEnokyNreGkK1cX8S30JTTPUj7qReLg+6Jq2I5+YCTtuzdRup5B/kL3vS
dw4mHkQlhIGZnw7K5v+9F+Kc2ArOvrh7x97FlnMEDv2Q9rf8S1FwDxR1aFdhk7oz
DgUra/ggqnMcjBdloPG/hRARve3AMnPloMWXFEUA4WhL5Xrn/CgJs2tygvUdDqDV
Q6UiMqi/y7VyCvyEg5EBd/hFF/h0WFAkLNGEhlTu8MLW3GnS9X/52j6WJdESYNFz
Kv6Uubr3c5AI9tZM4lvzQkNR8MXtRY8CMpDGWLwjBw1lhsj/kjFeB+hPHi4utNLM
pR+f2OjsErPUoI5SFFQE4TFmI5PPN86Zy29Kw1/kvt7cUIwtyCmHjaEqInleOEKB
8qVM9+yV4qVP2WksXbKqKmHtrfOte7YK7/Vchn5JKHoFQZXMF7IIdWlBSkeA00F4
oysqfaSo5MbWFclRr0dNE5hkzh2g2swTYBXTl0V0BJW0SeaaNz8SzPRcKneqOZe1
UtWmRk6zAOfpNWUAwMM1PtE79/4LqOEXQ5ieiFpv+Pv+bKpoUHeAMKDO4oMvb12z
6yWUGHGgLTmhqSWYW1YMuTH9Gu9QNzSb9QNFJBZ/8NT2FI8FzhCUKyzflv+Sveg/
LIsQo8ackxslAQh/Cyb27DL7MLdsm6rEZ4FzkXKKeb0I6BINiB71ZhmBVNwHpGeH
PIhepnwR3ynq13pRC/TMOhk/sT49JrksMtzHLZsh8Yyf7h7H1ZYBTL8sya4gewaF
66zxJ1IsZfh6dBFH7zHJ0Fr2MoxsGhZsBedKVWYOMsQbzyn+yDe5Elb141asOnqM
NBe5MK0r+V1Ti8RsOzVmxCIrZduXrTfm7EXR1JZXfo5U+PUq/l/OZ2miT64+2B08
ZPjAWynqaV+j7IcUN2yHPetH7kXXYNOBJzCkk38WuJ4Oxbw+a9OWj0h8XnBy79dn
qDt8xaOru9apEFCdRQt4EZGR0d2f4yIu/M5pKETcJ0vw4iMhRw275fviaBf2dPHV
QVDQimhyo8H7/XUMyJUbFZO6pmmvswxI6VRUkXErdumjzo7lBMOZpqxIMb4ig1eg
PL1fS4jj180iurIYylyEuTPDpeD8MKtrY6aHA5eOHG6RXRU1S3hTrrAjnLOLT1Ed
ceUAecuND53pIwhNGAsx7hKXKFgirVmtdCwG7oANa6RTQZo5YwdRj7wn26wbG+a4
M2rJNMdS5QWLg6JNmk1f6ZLZtXhvOS2Gkw9JGbtm3aabER7+ket2y6nz2xfuRWMc
RSBJ5eg9EeFudo2JgkGCxvbhVPi4NDrMcqYy9Aivxxjt5m1gWx7QpOb0afF7U1W+
rhNhE0htZvWS3CRmakHnSQ/SCSju9jfcn88G1+6y2TQsPwL5+gvH5l3Jo3kcr1rP
3Q3JDLp/v6rO0Ydck7X9DhMmmaAJN6jKm1s2fPRG0hGOJZoN4mmpQiyKuWAthdz+
jDpDYHx/6WFUdLWyDiSc6rq52U5KdtFfZL+epzn5LT1Ne1OgA5/aPiyHYF2x5Bxe
zjVVDK5aKtwq7uzLNyBEVQkyBzLUyWu0EIIA4aBujUaPZy32QHp1TbR3RNRtp7SD
hKX/ZJIYentHSTQ//34BTionoAwW+V/tHwQkuEjceMLzx0xLdoff8z9NJhicobai
eF+mlArH9/7GX5aTft0qCVC5wJd2fYw9es5D3KTYf8xh2wwxGGm4PdUTDYrWsHXN
AYAnYAn56IoVavkyjQLsbUwW7NmyBZAd4RLlDLT/sRp4iKHusI32oahgxnlU2omw
gfz+ThAg2BWX8pxouDEFhVhelAvNM3UzWsePh8waoADs5trAa9sE3ZvwW1qpNbR3
tl7JZJV5Ski/MQZBEMLOUPowGwltwnQUjq3/NuejSYCsqpP9yQOeOHQzw4+b8WOf
/xAUwXfwqG23bz4zp2nPWYhtMnPO+WnFIu1/Qu+rwC7hTWF/QaYlcjCa3y5jOeLG
GlZ/ukCXG3KuHhvmvZRLHo907tWJjY6be6975NRdrlZRO6wSvK7ug0NlE/MEfWM2
Vw0YwJizPTCofQnUBoaCNy/CT3VKcJUI6vAa640Z1rp7XppvsgVdM8BE5j72cvwP
LFfEEmW9ZdNC+5M2BHQ7BSnCyeha+CZZ8ht6E2pnXeVjBVbH3pry4pTdihwRzBS6
sEybJdxh9ltOWTuCZf+4X+jw50H9RqVpbCcMMwNr2R7BjaxvDxMGWavRzbdJdF3P
kH3DIPLlO2rAxMtaS+gMdAtcRVhYZO+q9+NiojCfytlK5NOLz8WUUPPiDPc9zIXV
y87g10OnOv53rkqQ8vHdoA1HzRAJHOMbZcrzjFAHpT+gBvrzyen/fLjF1QTI85VE
/mhxH7pFzckQ9pgMzmS8mRESUc9gjDeA1WUWwotIwZaAAM7FP06YSMx4Z73WBKT6
9alVdTgjOIalo+x5FxEnWw90jJVgi0HQ8z8vduj36PFuYyhIqN/Gy8BfAx3lOnlr
LYyGfvrK6qm8i7wddxAOOoAcYU6qQiWfS1Gb7+9oXDyGktG3+/5KQXqL8uGjxJmL
Av9Y9Q0WwWcYgns0mybR7r8oJ9nxKfrXW6a4L7ZkZ/P7UAPHRi67lVLDS7YROqgm
EOklURRj/EPLKgjuBIKX77QuiIatFHMENWM+GAlJZFW6Yc0CvZKneKPrXgN3qL95
gPt2TjefMueMf1YdohIqZj/BfCg91hs7uwqP4SpaskpfMqza/VTHzZ07OckoIyqX
tRQVkiQ9mrymj708Uy2gxlf0PHT1dWIevutdbnAdUWoGaz10BcYVJ6fZit3MBvkg
yqnFGbObVyVwNHRevYCufFcFf+MXfFDXgHVgqnSlnrqeOqxa7cD6yI7ZNwKDvDCa
aG9fsIbaY6AIso6mRS/42vh2wcWB8cBxi0twLJRahIgAWwC7UKTvm6+wTy4ucT6K
ilpVGGxZ5yjFt6sv1yAfZGwts9jkIa4VIF4dJHKpwugP96zJAkMm5U+6fcqSJ9wm
LaKs2zHFswYhZh8sLSPI9p5CQnyevyaBqTTsqvA9IGiBH3FuqyFVOvmhoOfiepmH
K7etj0zPcJIa4qtBNsbQX+jxv6WDpv+oPMPbECljVWkC55dihkQE0zQSfou461zP
QsF4NZHfUUGBXucDYln9hSrC7LTUNKs8MELYsS7HHTV3OMvg8N3A+i4YDntk7yz0
F4ADf7gbmbjnNGyhn9SoXkjdEsbbGAkJT3CGy+lDnIn2rU5xQUZFmqsnay6ZDd9B
lCG051GG98JfqfjhnpxPKNQ4SMIcAEQpPTFS5MsE8E6cI68wBsVITZP6LKIei5XH
A/nzxLI0y5fSg2SVLCmGtmbPqxmnkloyQh50OlXDGHI1gmV2gBAjaTRT3NSIM5vG
J8s0Pb+nUCamBH1rutCAr0bVzToZojmf3RaDJ62iq6P/ii2ACkglu66CVGV2++lB
hGyBFzEsMOwgaEd0r8+ziSu16L+fcD54Ualmk710s/WayiQT4OZgOcBZizn12ySi
kC+0dWtBRxmxg9+lB6yBrzRHL26r6aqnhrsKeUcbsx0vzQhU8CCoJuxCFoW+YtrG
YqpZqpu9um7rX4LG6eEiEeRiseTKBV0HvhAnfEGgZ2Yc45PStj8bL1Ufo6M/Jt9I
3VvADgQBuH/BVYlY319hnkV8WStmrpOPYe3FS1Kl4fxJha/ucf/r19/WDZeXt30H
mXcpIANtVuw5B9qqh3OrXXVz2nnch8nlH8zQljVLLRIdSBtOnipbxnnY4gEFcU0I
smzfP4HIrRIPlT3MV+Is7/1+yGk/fwpPbY+b2q4wrv8nYQInX7XfcugWzuQZu109
x97YzQ2Y6XSUD6ALXvv5BcgEKchgcOp1KmbCMDOl5+pj0tmuQeOpuo9Zb1MnRjhC
FDEIakZZwnkKBg2abNujBXTJ9uL8D4LPWn3l15dZ7UlnGWUKJuvE4+xnUqV07T2d
Ayi7mf4NuKiuwmnSbheEB2cUpG+QjE10hUiYGujAYx0VAGacrnOsNLm5J4aHecY6
fq5LSMtGUwYQSyz7WDQjYCPv7cJ3I+doRY4icUFahTAT1NPm66rmifStN0RbRMrM
7j/8QhoQ7zhH71e7IMcIxKQbihS1hdGedh0A/f6aACLIdMeV3SIPNBjR3TgibMm/
dKMSVUZWCVErxc66e+S1cVbZlHpKprrCA6hCU2jiW/FJcuOOfrMx72duv27/Zodw
LnE4wsPVZ8QO6aHXrM3qlSoU+DFCctd58Pg0InHb6C1P2uPMgr7Dh41ZH2XE56CS
dbt1qsox4XGtMoTNhmYMkk8F80tiu7iZvFLegzxqDBuH9UudWMkNHtn6YCqGEWxc
7+eiT+CtBiVqIrvHxpuoE6RSgWlKOvNdvyTS/nQreiwhwirHCEuMAEvzfJvzw96t
SCCGSOIuMDg802MzMcKSYmUzFI40g4trWdD2iJ8fgXRttRm+1Xx5oqmEGFECaHeG
uIfj+cDGbg5WoV0bgHpJQQOOTDHt3ntmp8ANgtihQdoUFul1cF7qLFEkrkzGrlZR
OByUS3BiqFQYV8kPY30sMjJAPVKyLaM2G7fpvrR0Pl/18bH/z+ODuGcnvLy702/T
ui4nkE+MezH6YMbeAZMp5IrhUQGdh1/U5m5ryghqTgoxqjB0MygSltoalm/+Gkoc
j/O8Mk4yStpkgpI/HFwunyE6ScSkWLyBC2rHWMkq9Zlf3ffNKPotRwg0hSOOQfev
ihpGiT1vq3wNbyvKmNoSIJ01iMxePE5hvqGOgmmqRtJqIIFNnT4NHkKUdWrn1AyF
qnQwgjtCXQZB91cChrrKIH/dpHEZlthXUmVuflDVHe92DSiIc7lzt7Z/YEfidn6d
rRlbH+1f4R87zZJnk7iSvsHLSo/xJt52WTvvp9kYVE8NI/bL3KnONnlC9bsyqzFg
Dw9uD5bGnAx3XpBaJqTXHNIMUM7/JumoyTzYmmkx9qP0XHczvmeymtBBMcST/pAV
DgSeohSRVPbY22Ofrq/0fxyiSwJbsELdzeJ0Lg8J0eypQRrUAbvxG7kx5psQUns4
AGmWNCCMdsyDb4qPEmVasOfgiUkC6ThRWXVHnvNu26n4DAFDLTt8qQaLiAyNYhwS
JdYmxxjZe6QnKXeFG5d2z765NzxBD87rih3ck1jx8ZUTb4WOWVvLY8xnmbWEJ5EL
FYZ9dUcAVl+voHSKBa41LfxKZ22Il2XdOX4+3kx5LjVob9cdOxiqZNqBo3qW7pPr
T9Pwb0J1tH4TluiWPDrQoXyYulbEc1AaKajD6/ddr4pdnNpEZwRVEbfnC1OAqR+j
f4Laqo72rNffAwM+LGAi5o+Znql8171gaEUsUQCXK7vlBA8xKUnsfiGOJ0QyvK8w
7slfTDL3bPn8aHUsGqfH76KTVX4gQ5F0brBlWcoJFqrorHFPerndbgUMhUXvKnMa
gd2zFHvI3Ou9xnvMoiHNz1q0NcjicQyaf71HYDTdDMHOubcWRzekCG2kNx0wgG/+
jmI601fZfF1m40whwvM2/iHnQmQDowAIsCyeNiJsvTSFoqaQTgwGhx/Y0fMflnkT
f3k5ZkoUJy1VP6owf//EFNHnU1sxUGoQj5z7lBuwLZwG5qHQW6rkzhJafOb6Xo/9
igoYhKMk4fXViZa6/CfqiN221Ld/cHM5cNf/QlFFj2mo2Fwos1KwLR0p8L/41l2C
jFjms/IL0JJFEuHQ2jNH3f2xJB1zjE35N44kvgVBO5pPkkK3j0ZIVyrOGd8Fb6Jx
IgmPMeAaY+CYMB/mjXU2npYZjtrrKQeZxMjSJ0einTDcW3lOvtp+IBZbKHguOpZb
6/SeiKS7D4/QFTZvy5wsEEpiU9gLNFPjAMDAVBjxp4WawUItO6t3nRGXbJy+0S+w
yIXAQIE/DFBNgUwJMevSSogVi0uU08TPmzO+jbEeTazgXQy0Nw3nJRrAljV3d3zR
K7n7tiNbLcgxfwLn0qkn/dSv6n7cxO7zORuNWR/2AFyE//KTfWGSFjpjPrEHFexB
nUEbu2B63mO3SFzG0Vqw295NzMd13HwwmzceqsQ9NjTbkQke/8b4IaRCsOfxi72y
T9irYMSmK7mxipbdsD2DgrqdO/hKXIoP2xzgOfk8A1hoYLWBPnJLa3EHCAwVSUjn
/X6MEQd31JWGPX1H4qoBmu68PATrzETFsyVXswVVGQJzpU1Z14xRCVvuJipy5hAL
0bFkKuhuKhlDfL0MF5T3gAs7jNdHIIpS6kiofmE5bqqvM4PY6N8jPNx39jThyHL1
cnBc1ZzvvAgtXHuMXX70EnWhMuCCDSFQRXZ3pSSZcSsNllbvelAt8T73dUcrwJcx
JcQYYoUX1mX3Vqofu17JtXCSQ4SN7RgtPHUWo7JjUVMU5rRqCkUW+TVjCNe0lxGy
Pmrbl2Zaw068vSqrWXvhwiw1dnnXXsfWHT4t/owKTqpPzJSBYlHLquuicsAvcWND
gA/9UBc3h+zrYp5I62HUgKyXtHUxJ9MoJHSiaN+Yr22InWPWWAiIMbUCRTiVG6oM
ueAQ3s+z/irA2RuvCbZzwD497ST8uIgvNUhmul9oEB6NbodpFsGTok9SKDnG7sgA
9v7UJV5afKNes7HYe1nykd5VCg4MDAoVvtXoPCENoBpdw6fUAnQNr0Y1hKZbRmMS
kgxq2AxEFc0iaqjYCZegHtj388uJ8/0aGrLxdurIr114ag604GN3IItYLMez2qkW
6N3DIm9g1BVU6KnTaIkaDxeS/4sxxF9HjIIUYeEHpCgu0QSO/XMl42g0QMqeSejw
nw9TDvxUaqE17v9pIojTl5x2MW4EUXGTmYkHxNDlKDG1l5Qj8mDWTqeGpBNH50+7
ktWTvCfzCxKxjJg+8tTqMgVwqr9t7kN9JB+Jbogyxo5x/t9bjlnGeseH4VR6Ypsp
fqIeMA4OtT/lzx3XkE0M0tfVVSa3oMYdbXUiQ9Q4L/HRiJfU56Og7v0Jjanu5RsN
nYrcLZ1qKq8S/gD+cngAvLiO2rHWe0YRTpQLAnCnCgkSrDVuSoyQVMlbRX8gb25T
3f5ZwGWE8aMWSw2mGvuXaTrBQeyWmyDvZhJz/t18cXJfhaXTqB30uN3csTwd+PCe
VL746CQJAueBx/eG2nS7WVzi5gD69G8JvHmOGfSgtTNl9vaoAnt9O0Jc4QPkUba9
0m9Xq1kBwMEXM0Sl2LmFauvICDUvcrD7VnaT4KmJlxW3c1VRp7lpgQEl4jbv+vTV
oRQfTHYQwXSh41Wu0f1tfFvlUsGivKv0EZfm/BtZku/CV+2rzD8JkucAOICm9a64
j+F437WFw9MW8zX6Mr7l3Tin7vSs3TNGHn26y5cJFjuux6PWz/pKNdUMScmAYfsq
EKLYXnz9qL1g6fNki7l5xilC2YFVI/wARU7cTUWgOEMDbWlxEJSxkNaZzV3igmW+
c4sL1TYYBeLOhbC/sO5q678PPvYQpDYS8/FEjVUwchujt81K/0PcwMFAPuBWPlpI
dLA1XGmk9/YaRTSl5Dms5XF0H4poCJ1Rg18K9wV/GfXljzrp1mbm7hIoE/jIJhoT
marTaPoJsN6BKkI1tu1V5AZyPuw7halnp+y0AFoAD20Vkd5nfP95RXRslW021g0Y
0Bx4CL7H/vxHXI3snxSIgugL3kVCREvq0VFMjjEdr20pBp1swypxEPr/ZAg6k/8O
k1gHOIMxRG27gb1NmjX7mDbVWNKZCUS6+iZBCXlSgsMKQChmJ0dA+uE7JfHz6heJ
b8W5zhWrv6889w5J+WEIl1fr9wdDe0fMb4uDmCB1ylf8bCx+6VPNry/ywtNgs8Pd
n3pwcXw9T7t54y1KUDsRLe0DhJeQP7pXvOY6s2hi7st6TBS4EiI10AjkYQL1WBVr
/xggk7LKtF6akGyCn6V7jwa8vzOQn3BUhsEj8CA4lRAntkffM6KfSkwQ5K4UoJXF
qBW+fV++CzXGVJHha2b0dpFoc6TG+g0z21AlyeDQUNxPSCZqaP4xqdKZHOpuDdZQ
qGquWNIVfXg2d/A1ihCCsw0vHQiwaw+17xuBSboYfyeHxmNJUbvQ40YiuXjWST/A
JovMp1EwDhCXtrr1mq6Fv3HN26oa87vOAi1mJeTJXsdPEBq1lsqTR1gxdXo4M4Af
mWQxARggwkZAy/XKOUIlv3p+RCwHpy1T/nCBe1jnYfOJV7qLBblQ/wuxOqtOlFHS
ZrjIi+VCn4fvSLYs7W7w4IjZaYH6Q+uQRVcHnS5Nblnchmf9DwOP2Wh26pYccnIF
dGTtn2PmWpiHjn3yi6AZRQkv+5K3Kd6N3UafFHqwoN0ttvq2/OcdSElZyATlKN0B
Cu3No5PLgzIJoqDGmXAAleHlqsCR6a8Ke/+d/+13NfiVhBtup4viXZ++ckFqwLuP
SHS4Jbj7Rs2AH7XwtuLuJyMQJnU2bsZKgwqGLK6YnoylBzMSvlkKh02BJv63erDk
qQ9tKKZAdmbAVSJZyQYDFWiwiwsxHQIk4uKGoHs2jS/0DlidiFjmyynElF90plUW
kTTGlbpdwNXAUWH18yRc2FpBzNpCKv5eWuWiAKKC6FYE3pacMkiXe9uv5CO9w+6B
y0qkJpdKWdNBR44Kwxe3T0ucfkL7sMgxG3wFx/8DNVX+YiU6R+uCZZI3e+WZElHr
De9xZfsrSupExCcBSLPzcfesvMRcVQvfpMxOjeTwIG9vdCHLLRy9jU/TyMz0OREi
cNeTOV6AOmfSt92qHaacNy6L48C2ALMIM0G3OARmLkakaPZGNf1qhpZhsn1E3RL9
x9bHIt6gh79UYGiiaJQzA+BP2n7JYJMrravBsl7ptQPVABPcRvTXiod+tlgdCqJk
dqENgbYkQP7V7oz9tLv6uH1e9NkeZBcGX0NWl9TDg8N3ro+ZJBlX+RzGCgFXZTg5
z87wCl3BV8V1br6s5oB3rspq/m5rNfAcxfIC7bzMwHvcpANrT/NhFt1T6qlahwQh
+NSvt2zqd/HGl65RUp0ZR3vXr7s+kp5vUDJe7rm++GcB53F3No9tWAjqmk5d06aM
vuRrFeBQGDY9TYuAx5423iF0rJo64PQcqcdrRNXLjxVXzye+Egnol74sPsDAW2X7
ls/JZJ60m81mvqrsWE+X5rQjdL/trgUCd32j1Z0wEHjisklEA8D2VtkiU63talOd
sc5+mdobq0zcz0+qHjE0w3UJnCmUCriJyHk0/AcKPL0Zc+eDjKZVPWEW6HaRl8E9
fEav2NkVoXzmINAVOcXR4+lW+waARDfd8HLiiYx9ikVRbPD0sD2ST6aQzILTfGMg
36G0KQTQEWa8ykyYU4+V/PcN+lPSNB1WjM0Ys5Q4p4KT9T7XnTNfLBBDXqoVYPvQ
TEtRbMVjVBVhnpkXkoZ3zh/M2aJkDCzwHrvm3aNanOEFvTLFWt/DgX9anIDaALwE
mTd1e2vooS0UgPzG2326NZvwgGe0uXynJzZ5N3fVECCvft+MoVSib7x3EzbiprQp
nYv5D+gbrZiypR5DRDk0RRh6DsrKYkj1moeFtTJW7SLTXcuYBTn29x5uS6xxYGp8
TJF8smtVN1Aboav0HpwW9OLaHFO/Uj2Pgv6GZt09Y8UAMUqhj17TiG0tyagUQRbm
EWUccJLZj0L39k9RX86DnBZzffLwa0+caFssK5luTwTH0EoScxUUhmwO3QcncsDT
wCH3AVNUUy+jKhQLzttFJ7LdnPIOHBThNaNtCjyT3II6WCDEEjCx82nR5mmmke/w
uRo+v8WTdm2GFoTeB0ShphzF3eRJIpAscqIunBQStAYUJclKsAxLZrkPtFYEf6nl
6hnUcVYV9ZHwNb797IzNQkVm1Z+zYdA+MN5zrFo2VYDMVUlREI9AT7hXIhba5N36
pZxeS4IQhsV3GrAiUeO4R6AfFsboRPyANA7qYv2tfI9hIqRNywpyyX3rFV+1cDkw
A0ImwQYooV4iAwr0HXkKGCuOiLQfgNVnzfgzLBIdM3gAR5FtpJKpyuVZ7iF8EtvV
QRdZVXdCcOEaDemZDgX2buTGqsOAWcH9xi3MmE5QWQoFX0wIfMBn9sxXcnNzLODq
ep8RddJ65zLSC/tpDRFf50NNkUVLNM2HmNUS6Z3tcaN0Q4VDh2mTmJNTB5g6loQT
fYRG8bsb1gKY8NB2ZqNft+2QN25wnBf0NTyREpgcHPWyscODXofX92dKsC17xU+I
DIrP3dEbO83K8n5ipP69sihm605G3pIfZ8DZzqEIRxDqP5V1o+uv8TqMn8MIsMlX
kpd5E7/EnfaEKXJ2hkY7T3glodTQX1+DaoQ4Bv+c4G0jNycBKYYd6PjsHQaAS3r4
oS3Xx1H724WC1BH8a0pvO4wwG9Vr8bBcoICOZe6K+bPHrZbBH+MJNhOe8Ka9/eN0
+oa12OXx2gqloWcvSPUW5eTI4QqFTiLkQZWV9rHEHBK5w8Lb3Sl+F91d3HUBZDk9
CNDIILQNCX7ljv8fRFjjvJOE6WyZyDn5+kfTJr/OZabnzOyOFFmuQi9hdejjPsvZ
irE0qHQ25VFPu08JAqz+3Sulue+HIpzRvBlGRc+WRgmuJ7CV1DiJ4S3Oxihh8Ai2
es8iC9PkF5vh7VCmiT8GdIR89Po1WavdtNnvhVSNTjWh1VTZ3VIWAsp8rseN6wfK
jE9jYqD6qA6Xtny4gGqH/N//9zDp1GMMS6QMgAd1eDC67E1wa2hlgiz7OaXV7Bcr
V3MkrrUUYX++OMThYSsIiplMiSHe+W6GyvB+Lkt+U6kbaAmhCvYm7o/LPYwu/Q6M
0eVFi86CbqaMkbdR0jEd2r3Zg0nhc7Dc8G9D/IMxwMr2asGVA/v73OhLFA/JksXy
mmab0RraoIP7FFH0o0zYCav2p3kE7jhUL09JASmCnbi4QpdLAiKh2G0tAV7caOLO
OhcJejIJIvhOPJbR39ocmIkI2P0s96qS3rLz+VcF5crpn0XrpDTXbNPyB2Lgw6v7
dgz3h3Q6G5/CaaDkMz1GuttyE6osKwGQkgsfK6wwgP78ufFdIDO+lyhWdSrtx8Xi
HsL1pMHF8ud5IlhHtBGwlrzjp5myWZk38kDfb/dnXAMD53h3ZNYNS8Dj484yk92T
MFW7NXOkQ9tRsfi2yDPa0uQJI6V+7P71h47hBFpm3+9tlIdxfAJfrZW58OWtP/Hp
tmeMBE/sjj9vwuruhEhDLoFs0zb7tg1rYyaMXHQodDOAqriMSbMS1G09qn4VccpV
fCh2RSS1SoIHacA/AZsoy302bBmpgruLJahUhCpqnCo2AtievacZ0pgdcWfB7N6f
/zBwx+YUFDKcW50DfYcKlLIRsylKp7affXDKrHAr4IcglL7TVH+p0gZQcGiIB+Js
O4DJo1KPBpzIcYUpFtjaF1u687yc/CosAMhlSQBfK3LKfiqx9y+eAu6a3UVyY4zW
D5Z/lWYooK5FjHEJpD7FmfsY8RygyqaOxhzgXr2k8Dl6yfeDonxGXKdjSh0PAncE
T7uS5EENp0kroYzVBrpqvNT0ZYH0e8UFyECBfvLZ0MMyxSPtyn8q4NRlytPApiwp
ieucsOi6j0cOdx12yisr5fb2BvXYRH0Qdjc1h/w1fHocC13jCTl+o0Aa70/rKv3e
MVYkgJtmwdQ1+SLKJfT+6b08oZNvtx0YlL26Yt1L+x1RnA9UYx8Lvmwa5PJ+NGXe
BAm0gykplI/3sM3tEjJ17zzR7HXTunm8/nH87Z/LzU8538XwEhUiMxVXMy7kLz+/
xd92Al0Q6AzwgdHysTpT+BIVHWvBXhmvxbouNSq2Yzev2N0sugvh9ksngQZkF9b0
bwt4BrD1K/piLoi7lgfYCkpVMoo4GmmSQx6jnVCU8wnDpyJl7Fc/MWLOeax9+11O
B70VATINZ5mEmarl222db3Rid61PAjQqX7FpWxebki7/sZ3irPokIN/tonTXLQCn
ddcf00kT1pUPSvJu0jNF2pQzMynVhXEKRxu2Przq7FFMCMg+QwPHm1vsXTJu95Sx
2wLT1KeJF3SxdUyWJnTYwcOFEhKWBrFRCGolxm1Wb2aWTbI3QNi5oBA7PIih53xG
q77f9GkJJ2Zw8aGnH9C1f2m9MqhytbX6iefpnWOsGHvRFj//GcATjLYBDPdh0kwC
e/SU4Qtmjh6QIukSQmeIG/Cz/gpyLBjsOPE1Cg98dNim80xaIZ2nCzFarV6f7zPr
q92spV0NnMKndvgeZ7YttTa1sYuX6zjF5Z3qj2WyG4+4qfybH3cB6IXFCgSCsZc+
+i8oVQYFkLqHaILhhbRbk4AKma02K7thGrRe/GAP45f0Yp7ZFr4MDrkeb6DZxwDx
Ha+pXR+vdazgsS93RGdRXhJAeGpEXwSH+LbDL0MA6kcPPwFv7RmyPnrfeX3tP2gd
frfaPB92Jhg5EW2rJvnXYeL6AXPvsT4PoXwKLbve96Xhd2ZuDkWmow0GCJbg/yAl
QIQ96SKmKEZaSsOiozJsSZBLdplG+ko1/vTIGbBiTzEFFN3Hms04Du6PXZdph10m
IaQmcTCmhfImGp4NYtL/DnejR1iVxH2WYlXH288UUNkeFp9wz7sgWuDHoyFfTjPY
bhc/ktRLYtLitoXBNbCJKPA8X7vBcypbyIdZkK09Cm+cRwc3mzFf9slSmAG8CBC/
fnzel/mKSyqGObFLAIpS04zQKXLxOdgFCGF4WPQ8pNlM/O6M3oXitCeu4wDF1xEZ
KJy5e451B3oteoG0BamlaftRN35WOLLK05UAwyPVJTQY4CAQv3AG8f0es3pruLK2
THrN9SB9zhUAmOBvIWgGH9e32R08i5h3MA2Mvdp9o5QMCP/9vFSrA5dLXc6hOK5N
fhGthpRPQH6/bJqPMUIajoJczb5VGEAAvYcS2F0PI0Rpo/n7PHnNn0fzb689FDw/
flWB8kIk/lyzQAVZO5eNNlYp+ICTNnkBASG4bFq1qALJPbYD0WLibzdzbWwhlX44
5PZO3qW6iMMahog6z7jivLgej7lKx/4oM39mo6//e0lZj/aoP4izSCzQYiJdQYnw
BLLZFC2X+QucpXk6CPQ2gw2v4A1JOfTG8/WLPWo6ANz8nWheTRlvn69OHvmUT6tf
ZAGlW9k7+WfH6YP8q2LV+4R34HGCnn9pjkWyIB9W+5UYG03DnQtMnZikzgJ48mIm
WhxcpgvzIQAhZUH/xRC6wCgV6ROR3nSPHpm86LA2D8ybYfmjXjxDDxjc4AhWq4oa
eBFsg6wPNg8GGTMv6jwtylsjqKEZdsPkp0KS4r32UcXDTxkezK9Z/IbVnD9iyCV2
lwGEuY9Vl7mtvIN97PZ8UyXiXPn5c2Lo7L+ho/QxkaPgBDxzj29Lh5pDhukqS8sf
Zz/Rfl5TNADzFizLRLlNDjz3Oxueyxnv1YUnmv1ftLAhQSJf2rqAoY5hrK4m/B9p
m567rfWJdMWSi7Z4XcFQgm/vzoPV42hGkRBLCOtfs0YIUXYB7ep0DLxqMe38p2rt
UKm+sBZBhUfpx6wpfe7zppGY+TFBybR7AgKAREbPQLy8fGat1P7WjexHFWDYhl2A
DKoCsvjeQhvdtQCj1+Ujr4xksfYRyLO7WNTyWPr23ipDY/1p2PptCOCuB+98A0J1
NsPf421ucfFd2T1IZfabuZV/7MyByT20i0voQsofV9dK21/EnZk1kNgyr6kYX4EK
w2CYATfwjHc84g983S3e01og2V+Qhd51whU7MXLCoLFPk7pR4Y3J42T2iq39Ljvg
5NTh0JWVEnth4ofV21e2OKEFQZTmSjdPbqSAUgwwB3wfcrpXNNZsBYpzYElkmb4q
2YIvjbmI4QP3eRbaiXun06c8XSDHqn+zymJXOF+UiJMeni6utzBf7KhZpyW+lfX+
83boSlSi26eXK27PO2/k05gv/2+VxN1Myigy780pfUMm+OTaP8/3yT7WpANSmDCM
zHYln+d7brNeAY8qfn/7Hia2OZE8WpUmHNQpbBCRcDo9HfJ8euYeZqCycdTsoWXf
WwYglKRlfKYyDVxLgngUiR5YtH5Qr1ixTdHAvFpZx3Fw/nFxHn5vQ87ye/QAmOzE
Cp2ovPxMRbikd1HEG4l3S5y8YVwd/PQXfGR3+sBAboWiWMmtZCy6JHbeC0mXqgSS
7qyMqWJSwM7la9IiHcuNrTG10ElpmDBhxOabkcPJBdUqp0aro7ED7uHOG57dx4t4
YbpufzeL031oaoEtPKj8lu4jUKcHW8tfQ2TiXxI9lAyk6u5H2RKVg9fvbzVddbB7
DXRDCYNng1naJpSMILztkl8SURhq/J6hsoWh8a7iCs2hiAZG07no2yMLKK1lOeQi
Ot7MAlXhw2crRxuLTMU3t0eaU1Cb973apbNKA6C9AgIHWUmrzVeZDEYGuh3YzylJ
kpTCogmc63La1xMyAOQ+AN6y+uOe6uD7VOKUjMjDF4YHq87KbyxwSfQHrBnJg0E7
2zmNXPLST0xMfS1yQUdGmXdIKFnF5MDXLkxwWNUvH3mwWBSCRdAs7sijgiGGpuyf
mJoFsGvQB+T0RPTGhdOi4fL9nWM3bzFcDKmwBtGBTmTBR7+JgYsAqaKu4lt6GmYV
z86fzDj8SzCS/nEWcTNViwvWSxrivwP8QIiiGFVWm54McN415yqB4wcR2xym3UrT
uvtYd7k7/Mh/skk3kGWp0qhF7b8djxoC3hE/Y/ozbm0J7DXIeNGgbup9CTwE49DN
/xp5jX3ymnvikerPH6vn9Y6W03eMCnpuAd78Aw9u6V9w5uBQmTVAsDREf9A6k4BO
ej7rwuoadvmMop3Fz5/Wirivo+I6sGWfdFKvXQr6i8HIN/sddeioD2Fmm0N4hI/n
qnsWNTkopMuD0IYKviikdnS0kz4wXieYmAC2145/VZr3YEOCJs+XicVAxXmjslp/
yoNJXS2TiP4QYmSNRS8RCy2FO3X6x1a2ETK7lyJgQ3QLMej+5+p3keRI7vN8rxbm
9vb38tJVGjYD+hJI8Of2sJVIQ8mVN7wirPWZw9C+etSD2e4x8NBI2t36XQR1nYbG
Txqe37n7pulOUlB5BKoBqcf6+sIyFyJMbqCDXQLwhpphZm54kheZ/k4aa7zJSQbD
b2yxISjCcKE6buOG74oGDEcMoIrK7zaOlCeEFV2NPeTk1+BW00ANJEPELTjSVrOb
4JRo7q18eOP+wdGyopfCi/CxNdteeRkBvQd3N38uwJBlvhwVuiI1DiWv542sLsq3
S8gCtnBHN2I1hONXla3vODiBF0P2onDNdIMWrci9U2K9DYcHVdwjDPOKUCPvfbTI
tJVhZTmnmqhyF2eMmS5eS5+5BEOTnLflrMdbbsiDjbXJBJzYMq/Q2OFycZgkORCs
lMKGwyllFLHVA5/7bBnJx6YNqGAIuf0Gd4gIwXWcwNcsqDYm+grjGPcPfin2C560
oTycAZO3pRK6KEdNoI1AXt0VjpE54sNaKaz3s3JmgZoXOo16ML+dBkgfsSFN0T8d
eYueK0Vx1ri4TABZPCzInhr6/+Itzs8ji+65387Q5oHWDK6Ee86TXU0RSfjsZntX
KtcAKnFGvqM2CCvAo5F0/+cVSFWJlEF2XEWg7GPaKj42sZM/q6JgQ/QoZAdqoH4N
aRVhUNbojfJZiYO4VE0HHdyrbFdzeACUa45q5wvWsvOJN0Kxep+HIitrqGR+NNM+
hiGYE8YyLf5OrO86xgCQaVU4/19xId7ohyYgANAT6La4tBZu7hpyiCUIXIlRx/WS
IwGCX8bkTv5L+esO5ihWj5bf6nFadK52Ep8dFnhg/0Lrx+79OAh+ZBDORihNrXXS
kvegTvGinV7Q7oegfGlm1GAIcZ8QKXZvgadqCQyIdREZNZ1c6lMSIj2jFykaX10C
9eZdedncY05qsVtuqERvng59GAtrD6Po+CFjIyzeLkUCuHTHlSLMGskZqeIjh+I3
zmuf+Az3nVa9B9vqiF9Z3CR3OVecVzVtAQbxtQy0NqEcU4KcUcWHDw+p1AjRCHx8
KoGjas7VXn9gA9gQenTZY4ifmKC55iKlNlUzThlxKroPh+fNMcVRjwnGhJslvay+
+ppiYVmDNbQsUydnCRYadMzHvLW0DDwOA0G/VBktAeTJg6JRVXdyRuw6vUCKd/PQ
rgiykUc8gly4BsSoBr+waBmpYLf/c846Z5MBcXB0H+AmqolHSUSLtq/8oXYMjkrZ
rlcLxzNmqHbTh1qJcy2wq11lN188OFjYpHedApdba1HA2AbmtEM89tZDqLx786fY
2EYJOpHW6Q/233HrgtIfrn1daHSB3I5wr+gAlwOfXlhi6DpuDCfb0m/BEe7auzxo
pXdod+iLd350JUPnHZ1xytN9s+HBdVO8I3a/q41vLRBsPs5glCyNfRQZ8vJx1Fp6
kLVl1rYKpSsDoDa8wq0XsKzYEBYJGASwGkUKIEBdd2cVfZflONuSAQQzs7IUtaXx
DtSxIgqnIJ+7FPXHJlnX9SqBY3SoXgbGdMB/5pnyggmOrE5v0isKQNSHJ2GrkDmO
djId3FKbz44YiHqjvggDukN6Z9kVL/xGanQwt6JyteEgo4MAletHti74o1mLnuqL
i+glaTAsJJHewET7zjxIOE9N9mmcZTwvUtaE9pLenOMe4zuzEiDrYvqZYyp9EkNd
O7L9fYhRKrn9HyD4h5m0tCsUGIFPK99X1bHLc6WQjJ1RBmkGmRT8+KcXJtRNiHk0
oZaVR9K3iHJA95CktN/0UMmk4EYGJcEA5AJbF+YBej4Ln3/kmOOvpRMmMeX7Y5FE
anS9rjl++NAmh34YJDuxec6TYur9GT/w1ZN/lu/qM0XDR/tfCcs9EljkLjwa6EGq
Ax1fYijya8zREdxSkTxrHny9bR7811ev2Zl9pupJfKf41lrkHcheS1NCv0zF46aN
TfOa46M72Ztsb7d8WvpVWVCtMOxh9K0v8NMziR2j0WouVnlVyTUDzuZxOpE+mHEH
pWR7KmRTxkw7O12f1TpTA94HDn71B84I3Lwde+JJZAK1FDqcY8GajlICBS1uH/is
1yw2YtHK6v5NFeiG0Lg9nkkVqUp9JBkScEfU6ZJBuAadaSk9ZQZ8DLi8vCQGhqUW
cveoAb6alHw4A5aF4I4bdFQjW5S9GjTeCSsps8Mt2bQp7IF1gM+/cg1C3Fd622ZR
y7efaEEWIHW6g9r/fvOzM/HA9Zn5NZkOy9A5NsIKJRq6ChzGOHW3mKhRk8r+d2oB
3LDSt7boTFFIXhQ1Bcas6nNa4366f4Ze5ZYcXCJCtyJWq+K3Ogec1NOXkNOMzP1j
5d4tSPK91G4BQMDpl8bP24KTTEklfVvvsV5zOR1Eyoi4DFqCUCrh501nMEjFNt11
Be0BAlZQr2SNwt0AKdr4Ae8thBoC9ku+igaJW8LYOdUxpe65NyzEYih+W7OEU9I3
Ft4CGNFVp9XB9IAa8S3FKbOzq/dWPErgCkP4od5UoU/JIiHFjZ7ZtMEVUA/aYR09
A+qo36xmpwXBWE821g5g0SM2ZISkSMNjj74OkYlw3yuoAFIebHGUs1vpuOMR0kNX
k3eF2FNWVy7IkPY5Go1kxtaZpdYJx3f9ats0VbjtlsWrX0vFBhE1bKu32nuhKmAR
2DkqR4pwmuuQas/mboMpAJbIBtYrXaumKJAHn5PkgiIpDTUyRWXp8rEI+ImCxmN1
aGEGi2yX/nhYHuWXBbaIkWv2NYCd7bcVyNxo1+7lAJf3zgrgmfYGg77nMqS6XqFt
9TjZYyNUzF9am2LwGD5G826qethbJawfxYJhm2WXAPb+avTdprYDjS/59czxDwkj
EtHDKJ2ruWfjEcYO+MrPstl7nGOv27jt5Bmkc+IoYJw6ciYgu9jQfc2h+7099t/k
hHUB4G3f6vHhq+lPGYOHXl418ML4p8S4NBgS4q6KJMkwYYStDKvqzICEa3po1c7D
jjw862ChTa2uWL6bCyJ7GJoJQcjEW2f8O8EZrEZ1jNKrzNbAe93KtvJyAFKrrSBe
aDHSKki4cOIVtIt2ORm+TQF6LUQXISWwsPVWZwmEgTScROXPh/jPvbs32BXjNKlT
H6MjAl7g1/rNDLtY/t6p4ReJ/TWZ85nK3tEE0pCIlgY3E9vQCgixcnAOqvoiSJhg
nt8ec+TM4vT1XqixNcivuUMDhX2AThZam0hkX0MUS2c2Xhdc2UNq33LjX3/gao9K
nUf+CS2t6ZtMwkdoNpalKzRkJ2c9QY7EhDre9bYpCpxxq5pyEzda5EgU8NruauxA
inmWOGAKCeCkANAd578YY8Xj2zSfxEtHIdpZCo9/E8kR0G6ILfXtzC9A1bagiVSY
lPuRyUgzMy6DAcRpAyg+BvG+bcUguaQ3GgqWmWdjLr7lGBvgpB9QLwLNKdPznSQE
b33XzNU9saYP6XOzfvURK6lVcdrmDsSYwthwbXNRmnU5+Bja5R/dLBQZPM8CRCVm
QLd4vmSj9aE9okD0AJYMPFz5OVi6f6rrGYncDSZ+4Lbfl91N/YGUeMmT/j4mqwdn
qwCPnoty+qdEKT6dOqvYs/lhoaOGOm0yKEmbVV6+INznvtDeXxbGZiwYJ+aE4KrE
ijj3bKSusnzDwlbyNJ2TPvmrlnJM0U89BDA/wenXh5jN1A/xGVVEiRfRsOzoBWXb
CtH1qwZJijRBDm/mc8pDJ60bdbMphbpbgOXfVTKj5cMpuqdndtomZObd/RDZ2dZp
sTHrFiv7uoB5kZXKb6gDVmz9OTQyqDemlOtBN+njRCseHiUQsnLfWRx5GIMnhHLf
2rPQS/9qlkrGi/4fboDZ10ciKWWhGUo4w15RxWcnYRCZ3qUq+08xK5MHQ3iurtAn
F8G/4veovOeK6pNESFaQp/Uu+0sVb/sj3a9vE/AykhLkGP+H5YEkk9ODKdKV/O+L
YPzryjiTgCLv9g5erwuvrfb8V/GO5/eX8KWp3EUoHaOlGfSQ/mzeBX26KKa5gkJb
r/tRRJ7bw2O9sJYj5/6gf+PWxuN32kVxCFZSPZGWMT1hjbIKXFzQyTlJXxu4xJ12
8LCy26s25t32inkwAndN7BWv0uC52Sb4TJ0O1qAkqiYREcp/l3/jYADCuHDlRZ6p
JfBdkw8mwpbdrz+jlBJrq07G6qyVr0mF74ih3VjxbFQVxnx1rF6KXAxe8TBIJn/l
ECRGj6kbNTkYk+Hb8gHxmknmhdc3Bq9huTXjxLAV3kY4eYDGewEcBuW36cduLq7O
bgEMX20lvC2R3BVS62U6GXVPqcjjYSmKwtKUXETXM+rdGLLsc9bDHPrOmlmeU+Xt
lbpqMYvJW9pcSZOAB0LxVB0pbpbh9ym++oisciGZvyQMTPjm3Ewsfasi29fBCzEM
htIu5f5SPmoK6Ti501wyR1TMIxG8GOjVzg67FSTEpm0y8RE3wQ7H1gBBrDIfgpm0
kJ0Xk5bxyDQFdNdi+456FG8nF6rLXJB6tsBWQhm+LsVj5P8he8c7vsRkL3vVy3Oi
JlM/6O8uQvUOty/Lhx4xGXwwGHDTFtHQF8OR8rFrflkCgiD3sUkIcgzowNdCmRUi
5aVcriSB5pxx7RGp8wImFDJwgviXN5TPLGyh1VPL9WR6QOwrplJz1D/b/88LFkto
oi9S2MWLcUG5jkSi88NoE2QbhvLXvuPmVlKe0hX/FpWnIMpmWoZ7j0UhpbQUZxv+
hb5aJUHC+J1+AKRLFJdkqbTk/3RmPRA7Qiefw3xlkRzeK5gGBQ0XKDvJGMZbmkV+
0qk7N9pxGxWOSQQQ16SD9HSHJjbGDf4+SctePS8C5lL8ZlBqPPzAMwSRMVDayPei
XJ+C/yuNutMxiVl9WxyxAMTQpPVC3O1PT31TL+Ptm2/otTYncCaxnPpDDEeTJ8pG
gowudSFkpgRFOyTtw1N+vKTdYzTXStRzNLiLyaVGyW5GwO7mHWEyxnWhW/t81OI8
JoXxxNArHhxZ6FlNdGkGWWWNwxigfFYrfJAy1ffK7Y76t6jnT7HTnfAGf3YcLOUx
Suqt3uEV436tnXm24Er5avN7q4uxJIxb7VlKuJMT3LAb6MdpkEdl0JxxZggkHtIA
zql5Mq77glZSmdUYcKXAATb2th/Jo6SD9zGDa1Vu90+Q324A13ns40OsRP+wSnSN
zBJHRvYQuchgH2eygaCff/ljOLD33iJACeRHD7qxto9rt8W530fwdETc1GJCl4yE
8JjxSJjDo0Dd3UGu8oh81iH3bJ5tv8PlrDilybCD2Qwkxv0YZ8nygbQbsrSSo84x
XPgkbxoMTjrX2AU3cHm8oBJvEBJAK3Z4HBLuuMtKUl0vS2J8zolKbw4nsqsXePrl
tcBeKgUqLzRJDCmcINypOajiNYxEMaJXNw1xkEvzycGNWg7/x0G6utqP+fygPVV3
7f33QOtLvi+/3nhaJ6JUv9LVdcHNWb9O6QAMurvmplvhq/BIssK4ihfIp+A5Uc04
vJ5kt6Iyhw4JpdsruesWzuimL2PI+63hfysPhNNg0Edo+q5s5CmcWlvNPakP5Ld4
1tfiov84j099xkmbMdTy6SSpoU3r5HU52/7Rb7YvK8P7LfLdWxxHPKxWm/+/dT30
9CZbmfOud8/9dOVztVbtvlgzddhCoTY1gprBgSYBMi+7Bb3/5iDL100YVXlVozBn
N0zbKq3zgRXj+tjaPOy4mf7qnaxGTVRKr4QCLOGGS8TwNqq7shQ//BUgVpiL1JQR
H9zmVPuUBCvRyBeGYdCQsYvVk9D6Fuz/0+CLR286t1urHIfg2RxaBpIiaJ0eUgif
l+W3azRKz468GY8CVMd7mwmvUHIvXn/piQ4YjqC/56HZkdvx7R8N5Rhrk77CKaVx
9zYXixD7o2e7GzIL6lHa4xXsdR210J0u4KCvKu7kkOVDnKyKdM4LZFXMc3qJ5QOh
xua5fhDZS2KK6vYbQTrKvnNcKhlKA6mSDXNWF7xoAjqF7AmBIFcQTmRJCgME1lCo
lgrPbie71jQgpXvnYaEP0A48kIDseFULfC8aydCO80IA6G50hAxhEdv1UJvHaPHh
GAi/Ok2vQVnrf5E6iKEUKHlLh8GMhTmFUiGoq2LEh5c4Yx6tUy67VtJzZfrfHzHO
eFjixwo5/kF7EvX+dsscP0p71Cas+3MVx+JrlEY57eJVVXctl52WPK+V9NKMdm6O
5osREwruXmgXiDywuWiuPHf96jY79L+m7a39RD0I+fzI2DXiwCTP6zsKbW0FgYf8
fUxIWdn5uEw4ERzgyd6mTPdELO5+hTaTgBbkJx8thpdM+WtpO28ovCHy8a/7iPkB
TPrfEBVL7qrtfeMXY+l0MRTpImZA2f2Dtk8s3csZK7QiEA/ue0vH3xdvwAXlN3Xb
pltxcI0GHm5RFlZsBdxpaG1RP/IM+9cE0VruZS8Vg61b+GrYUqG4r/Eyim0llnLu
91V1KKHQNSWmqStxlkU3+iwnAHsXOAg9NqL3oj+dddvybmr3nCO1ZYRG/gCh67NG
bN5DTzh5AfpgoR66NwEAmgQu8fnyD9NUTGz9WiUvBIyb+w4dqki/1KOB0ZpzXbIY
UdQsxu3/Egzevuv9sV+36GXQMA/rVwsTA+/fT2rC62K4ulV8c1euYgvFQ3DSttsv
0EKK2A7DFBz1TtBg1HvPrcVs45zFGtmPjyFus5q/cvuudcx1VpaR05XsTpCCCd5v
6Jdk7TB3DmcdgeoylddGkeVUSwP0uWhvfXYW3okX5Y/oOEQn/pn68R3wh/wLm9lH
4uU9IQ1zo5538EBIIavfBfoNRl/QdjYC4g+otU6kvnLbCW0IG8itnnYFnnAYqOwF
z/JyuqkuqatqxwFq4oKns13b6+0R1iEs6fuLedtXVgmgGOoDRu2hxtE1f3JkigpW
/AWbsPJFk7n2fPKhHYTF04pNQPL709hXHzHtkYSKxZemLRHVFia7NCHFyYWk4mxL
OcLh+ffk//FObTmv1pbA3Bmdy0Dc4kfE2zOYls7uGzV3MC9jZ+Gd4XthGZ6Nu7Qz
5uxvw4B4xsfZbzGHSWjAezoTGw1vRPOAKgriqEOTclun4ONUVO4UMQ+RYJ3VPMBz
VgMvP/4TxUD4wLZuhF18ZCxkFrRK2hfQexwvlgA1G5+qLeNouEO5wQwvQrzFUZlU
Dim5WnHKTbY9oE2GPPwNDLFe1k54Pw8hwJs7lGVuQrNWHaV9GH3OK3TsPa1ZL9+o
Ej6nwnBo1UHeJS0qVmtxFe3kUS9ttlPsUY2eDDQoRBm/jQixyL6cTkd7ZWzOelRJ
KxCx48iMPxj157rrPwsYHzmuIZd8MMiIWXSJNSty6Ua6UZvF43B8TEudhQlrpnOh
oiqEIvG5fiWyHDsIpVh9MK5ZeyhL2dbr/776YR4QiactyGTmjfSSZXVpLA5vanAK
/9x0jQbIvi7YZGNoc96Yz51y/FgC1clHzVcA+iTLp8ugbOWYfp3Tg+wpNaUeb4EV
QmIMMNwvkA8uOP68Bk7A9TQdaWVFsNF3BY6JfhcDz8TWGQhSlV7kmYPH55RDQt31
uHBjskZjWOiO5WV7qQv6IDnTk+ilBwCPLHLdscany+Ob94NSZnQUCTD6Fsm2Ufxe
3Kp/nNI2muGwsBcvMBiFpOpH3J1LhNJQqyGwrJOBhaHtSe+Zq+2kYNvqW8xTf4XB
++DZKhNxy6P5tVBLDEJ2amjpchCuAJxxFz6VO6JvfxobZybsymHshu2fHQT0JIGt
sfGS41RorPQ6/qDzF+BLbbOcx6iTsvG1Ho0puOaE2Tleu1sAoPKXZ+g6K39wA5oO
AP59PtVbm9KcNdnDpnffGcwjm5wCl5CagYWOuICTxCIuziFXGfgdtLsgRnbgupcv
P6CMlqs9iJgFYOX+WZ+Y9l4BSO8+AmRWQJ4U6lh+v2CPBFG1qp23P7xhPMHrhugV
iXKQu6lNZVifQqyDw/O0IC+zlAnz5zLtJ6Xh0fN/1biIB0tjwHDCb9+T73Eat4Y7
jt5Z7XS9F8hokwuwn31oHOmZzm9LJywSYVhXyzc8vgdJCGRVZnmeDRZtno/BkVFg
ctTJqLO7Ndzyg/JbDXloesS8pglDiW6IpwWGFKoJwsdX7MAjjOwkHPyH/w7/Oces
ZK63B3hGVjOIjnSwUqviueLCOSiTEfxAdahLW3g/NR2p7qE6HDBw3pO3XSb+VTM9
5H22tzlMwuEz9OPAoazkpBqrHbwfs+xZL4HeSXG6ZOovq04cKCbtK2shdC0f+kXB
0AntuFj/wYgpSix/TQA6LGBSVsoKcKErP11Vm89tmfIjuLLSCHJIe/KcqSv3NRXp
rdH/dEvx5hwPVWYG5R9AgmtI6HYaGa1ACCMkpbl03eE88SeV5nPDkKCSIRWvBs0W
wzAVi17A8B76gvJr6uCtghV3HEmYxswQyuV5gSmsrDJuI8qT8xHuaNkXEin4m7Aq
KicbASXvYsFX3C0hBbYJOEMJSPHHQi6y8Lgq7G/o64WDQtfS4xtHE6sDMQ+W004+
Oz0idulQAWAVqIPKjXGIP9V03v6RB4C/dSJ4U7dWFftKn3lqEfRSS7+Aa+JGI51a
UVx+iN01IBle7OcGfk1j9mGSZsLRR2q+A/tpBTqmJlBoWKBarp0H4EV8j2d3R55m
DDmNLrWXYPsEK/Owq8tjFnud3KlrouKFCMpkGqPOKjNKe1I4QUQHlXOqQHwpVkHR
N9U+vliX3G/LRA7j2xptWO90UBqTyZiuPfz5PczRj90070K1lCUuBo4qS+pQSmGf
3q5uSEKHDDV+CkMvWP+eSkh78/nqCISBdNHFWXtM1DEH+bPEawkwtfmiikq04TiF
ldbuME8dMqh39QlTjTb8qZAt3xeSuH9HvGwFQRU99KPN0LAGwiXDehtSLO7sro0u
XDY2bYvowDpvw0+IuG/eQVUSJMnjDkQZeDLQQj9z8rwnLm2QrvRY7Tl9iE8E+nSZ
MN8ffYSR7887Z+rvjDGiKaYALuEyfEm32/iyyGT5JpREqJnsjZeAoc+vnqj8tbj8
ZyTuBPAubMAWc3oaJqtaK1YKP3ARXIIr+HpmdldnXASeI5mzOcJ8qrp2X/ldQVzq
uupy/esk+SawmBeLJkAYqMN9Vq0vrXBPLvHgfDwQ3C2A2NDx8vsa7YbgO5gjUsU6
AyPkQ6os/8TEje7oG2NYsxrpeQJ4tg/Rlgbrb5Es1zJcGJZwPonTp9/PPK2sHKX5
ccVmy7G/0W+vwH7AIAbKNvXywR0NGVEWpSpp5ML4l2cPbtiND8R912gHlebxUSsF
ttw5i/G9Y/m5hwcX0N6tA0ElAto1MWLQqzKN8L5vn/81/iBV5yugMI8lPphOQnxT
7AlbvYJQZcf3HKgakPK8MRnNPbDlzAQR/xp5DqH1ONAo+m1HdgkT9fBBLVtR4CD5
CAviEC62nOGqIYk2LI7wNb5GRlHFg6LmLI3IocYvRr/xqrV3LCn7ggtS8HHJlcs7
YXkcLu+3HlYdu2QRknW/0wlY1/cMS6/WObq/MDtQsRjkPn+RL/ELvoUwBXYYv5XH
f0hYLf//H6aXdd701GMRcpk+lFvA24oNdavAdI9VC4leuw2Wus1b23k3QLFC9ICN
LCOGzziRsZjldfv2icvbaTHTqJTKaggNTWv7z7yCQ9jI2VMLNdLWmAVt6OoC4Voo
gGOjwC1v+kKXtCLoA1DkMiG0tw8WAhSfa2LOK05QzdC7J+/KiJuDor5ldCJZykOS
TMI9BSActC9HDsv7cQeTck8/XKVdF7L9eYCPI98QwxAENtO3LjtBINqen+Vrts9z
7rV0IMa2UT861OClgn7Lqw532i6/QVZtG/f2hqbXboiZvNP5Vo6UM4OH8AO/v5dH
PlDRuAkLS0ZpOI+nWZ18nklE8YL8MOTSYoIj7Tg9w63fsRbmq2shQ6eavDuKaZ9Z
gn3uW43r0gGgk1kWNSvZIpCJ69h9YOM9xqZ6Xp8MHOxpLunyC0N0LgO6s5SXAaUN
9xyeQPwuJmldC8bwDwmW6yztwLEye2FcVWlAak3zmDiMBrz3c4XwXH004Ret7dts
LLh3krgb8CoIH/Rd+d/jWIvq7FuBH6oZpUlT9pbLES8jZ4ZnSxvf2cmBPD6HLFhq
HvNlFx+g6aVUHWOFVbf/hc1HNE35Nxq0Q93+VZk+OQOP/spk8efTVcSr/1EzSq+M
hc1og0gsN9perhLCIHAdJ4hqRF/2jXPT2R0MmB8WYa2lW/xw75nCztOmYJokLZ5q
Q4TgwhPiFSc/e2W2FDsFWQu7ubPevXn/+UiKaggRTKzUflnQRplOTcP4UtB/6PVq
Yofu1ZJicFMtZHTUpZO6wHaaXY9x/f8luvuVV69GsPf4r+BPczEHcLJe+A6gveZU
ppEz00BFkiuBKQuiWJ9BnNJv5A80Si/cSC+capes6nEPViPNGS9Hf0wgQnQp39CA
IwbAl1H8+jEnNAiW9WroOt/4cUPntpAV2HwN+RKnVzqlWyBtJBgddDUntysmU/76
f8Spx2ojdmOW3YnNhy3ojdDqmYeRceztLcnyx/sV6YPvavv3bKIl8m8GWBNUXRXT
dpgVtE2LWKdY2tdc4sAt8hlyEiAfCD1AY59b82qUALd0KSAXJKwa5Zr+VnBTa/lw
lJUi2VdV+z2Nk780padXNFYQadPhARNhJVcdfw1QNqrj0UCC5GBt+VbXUp/ZjPhB
Hjye8xgGy1ptz8n6u3aVozfvITBeEY2lsMhbhyH5tNg4Z2YWHJObFaJfMuzVkRo+
sKQrMQXsr5h9S0M4wNw1CGd8g8W5Aomk8u3uuNqYC9seU5bkX0+vBx/5tPUkyVFy
sQvc0TCrB1urQyveLkyqzgs6EzJF29L0o6xM0RU74KIJtv7x/onPNVqx8gAe1W2E
vpI3gyGqSkp8kvWZph9ZlX76bBqwqHvkKQg+ugR/mVdfI4MfQ83b4yGaIUqU9/uT
9e3Au7PI4ZMc8d90cvDs0lgZnVKqUYNGynoovAgWi+88wJOuKWm/qXOjChf1UB6G
YdG3NJvHl1osepwMFUZYuAktcF3YTV/mYVgwNkdhdbaugS6JdZnK6Dteq/v1GqnH
/avF7mKTuiV0SyWWOxpmf4CrY161jVaW1KL38xEZ56uEAkkYmEU5f1Ve0G9kog/c
sQQuOqSG2GV2ZeIs9uYk+V0Ro0yeZ/TUZZUyKDWrvIqJUS9ttzeCNkWl3EHiTgEg
td8z7PojecMoJ0X35qZytUasOo7UvLwxo81zwsmFNjtB068UOHTaA5hYphip55I1
NHrK1EtGMJd83dYhKcVjbe21OydF7AaHk25dJ7UfbXi4Vf//YavJOoB4Gcp5cg5j
01KnZ0xXubt6NzG/hd7+ro+tbB5zK5lFFyZcXIaJR7NNbSXdv6F3CjNVy6WB4VIo
LjDDUXP6Xoi7Pekgz0eoanG9XwHa1Zf70BJMDNyZ2gxPB49FmQotC8YG3kJioghX
5Oo9G+TS1AkPyRVyd8AqOvNUoDJvswOTAobhbME1hLrms6+UHLQUdh+xNeJd91ak
ldXoDsx9Qz/QggQ6pA4pkjSDHVHT0Af43Fm6xmysvlHAUS3X+FQRGNVDboaGOGs7
hA7W+8PFKLMoSn88kcThjBwgNgruu9k2d/96qk+zN43tFdrIedXWE6cuAa7yGDNa
PGkk61YpRVrs6XAsCo/70HJE958+6cCT9fTCO4FA7Uuyziv0S72ronFSTYlcJKBe
sZ4gwKzcp4cj5jegvM8795BV2Y6Wy8ET9YA3pjiOetvW8R2yNK0CPT70zVWTM3qM
bwx9MSh087laofPbUSgv8+Tok3dlTI62PtlCGUow3alK1G9RURF3wbGTB614pww9
/GFBZe0b2U2BV8R7kZ+ogZ1UMyORj3l945vJJM4VzxbMinAVYVKxGDc42kxqaf3E
eUV25zazenayAgio5S5CD1zOyruLmsRehxFFm/Tbaot6SPkhNI+Q7jFJ9qnzqKCe
i3l3ApagtVddH3ITcZ7zkts2QHv/0Rxm6MS6ehVJE4tgUcCvgQDjCh3mbaAMigw+
Lg9Duz28cpIb6TuRTYXNxNj+vyDDbKitaZi1RFWypIi/l8pj5hhXA8ZnzAA/ZzN4
dNstxAVP0FWYIu0ysKVb6TX/gUQU9XBpDPo2ZxrbNPoPhWNv94+9feDLCQRq2vde
K7ExYIeHoyr84W0nlOgWvVxu1goyQaeVdVKA0u53JX9eRfLFve65qEN/8+fYZdai
UItN+Xk9fE3NazVytwhsJ726nj1orzYWSTiwIQfesCDqQyaTNN6bOywAoTwxV3SG
ut8omuzfpMJ1pav3fGEZO0PAZAnmYXixCUPdXk5W4N3Cp861kOoI8CUnvrVacBaw
wtYnJV3axRdbgHIYvXk/1a+y76c+Me98yvohZ2g8VK6n5EkoDY3pzFNhzl1Q7Dqp
9cKEierb/rHCOBbyyTnJBcwT1hj2DR0dJrYfXjJuiMxH8shFL3YzdLSYSF/CQPL6
ssEzjTozrKK3eyQQ/AqihTXOxesyY0lHXO82UBSR1U1oCl5tpFaUMVwf9R21DHiQ
3FPQDtDqlF1tlchpHGFPAhV0eHg1Ye5LaqhqWKzDl+iqAxMhB/fN4e+B5IJGFO3W
0ZSwns6o4tlxa4TXm5XOPgwzYo5AnFFRndAEeRuxh2xIJGRsfoMuDBQJjI8YUv0z
Qq8Ws5gmCHjujICFwcWmSB26sObDGCRTPm410kt16uLlbNEdqhYO/eDB/y1319K8
VGa/gNbI6xUzGK1Mwme9EuK03yJkgThFFnq8wKc3o81WLkKu78Ah+NWPmuP1RthC
wWo6dxOnotjs1JE51oQ3j04xdUHUSznPR50/hyn6SAOP8rWScGuOx8P7Z1mIhREh
P0x+c8GcnhtY1E4sB3xnL5+hrty19isjEbcWEKZu/1oto9sD9HPdZVp0BHMYY6fK
yoUBRh/IIE4GKTrC6IxsovlXR4PDvPppOnf4Uu3vvihOYAmYwbxUEe/mVCEsE/6e
s7/CCTAUNXzvsc3AyCl/0SNlPVdvOKIn3xM3djllVqEF6AHIHHR0deyYd5DE+81o
cF/PGXQce4PL37kTNyWEbtM0mUalnGr4gFntiIRJ6H7Yi5RCHfNLd79tPwbnyzuH
L4dKV2Eyi+MThAYdvv5npembIfBGNmITb3r61X5PpzLTqMi3rcIrBLmDetOMQpvD
opR7SOI9fzg/GcxeUQZIglv93d2rtFcUHhExrYlLlab6i93mOosPn8zLYVlDu8rA
gBmpB2qWWfxLSBI5SkHh9a3hzAb2AdQFY6xYFOp0KbF02TAlexzQEEnSqMSvZCTy
gqHnBjzWFqzcUmyi4KwdBVAQazM4QLo2xfX7RImO6997GgY5yQnPu3KwwRIYrMBx
N0Sk+S9PZ0GVsYw949Y+ZnZeZcdc02nUHde9eorAxGr0W7gJxObl7pUgUlWKnD65
n5Wd80BjP03OFm19U646afAqmbnlmrY1aOcTpyeiU03E2vuSsk1/4OsrlUCFZ4iM
GtqeEmbCeChxoZBJ3z26dQV9RW2fvR0Zsjy0wXBgmRd5VjmA3EubRmjoM2Gtl+1A
IOntU9ux2zG3iJH3hQHsqjFf2t5pUcp3prziVY3680+jMkSqNXnK4n5x907xe4BF
PHcbXGP4g6U3K+0+kH+37n1n5ZLckS9+zzAs1/hjINEi3JK7p7wZagq6r6Zcs2TV
HL1HbE0mqZebvS0EXudzLDpy2nfumHvTi/rAs1HqTYpH4hB6risEwT5KggWxYKkp
bEkM/dczWQ9370X8ORtTFsEEYyQuHa9sw7z2HaHZT1dvwaH9L503Lb6V2ZgOSSBH
eHXP5gmpJLqBGsMv8aQkWt3bPGv008XA1k2Jy6LlzkegoRLbP4fqI8Z5JNo1AHmz
yNuP7Nx/4SNaB9VcpLBTWtqbza5YPTticDaFKwYhTlQrilNATHsAWI0il+BvocbR
G3CmNTnGsVgBsD5Y95/v8nP9p6HjVrgkEoenUxW2yv2K+wPbatL1NshfZLyHD3uc
kFrQzGgeKFiYT+w2SLrKAbvqNRjHEECYx2SREgFEjzZuePJCWzd6RGewIU4mMchO
8AZQIbmrUo4zKiSeM29odZwdMBfwInTWcNez+szhuG+9P+/IU5YylTonYjsKUGJE
S5yvXz+VJsOi0kOcCB9lkN/D8rWAT76+IRYvZuO1CWyUhJ6i3BPyIGoVFrQeNyua
XoyVaQYjZLDhyDsNg9sTPkThaDVEeke20MNCoEkMdVlYR6KOFdKMgV6M52Kr+cUZ
RpxVlZseyWfZsP8mXkBk+uvf6/eZsKf4CKSb2dkJGozU6XOLs5k+Ez/ar1QI+akZ
QMPFIAUTjUxatv6+Z4enUU+50UrPylVYybY6lStoUTbtC2TAjQ80bUBgyvPA+QeU
PX5wxV2n2KQ+n+lOlacj/0GcI0bowdKleihA1dRNQ5/YuYlvEsjxCDOskHCiH3Ml
oDGZhq/BornfFdsrq52UbT3CZKUsKqm51yMK1OCxBJ1Fqz0BnhEiqXXCqZ8xCmin
KPd4rk1TD+1d+DfXvdVwILzwgouAzQwWV67qz8T08hOMo0OVsKAo385zbde2UWbh
i4Fz5dOUR0P32FgGvB7XnZh7TCH3wN2fcdb4btO7XRfz/gFkUaW4Oyrw7jgRAERM
4UzJbi84PTNZlM/exTgL28mKmd6xYoyhNNPakyK7ZS+PuIyhzSDiyUGevizCxCIo
cz/m6Yic9+cIz5z5bvBhAEXxM84Ykm32iJg+JnYHabKTTkbkolDQDryKdhmdKja0
ttBV8BunDthlrNL02JlJIBOJFBFSPDT2yu49FL5NEFoJ0uCG2M95lxB8/axarc4B
D58S7n7WeEwiJX/u2zrIUiETM0Dy32OHHB/e2tkAuDXYjJmMAtMmjf4+bZuO9+17
yxj00I/7+uxE2EWVsiwvBrEsBi/0SJUEP+UaWpGRBRqjM8dW/WDo4veuGRr9vw2f
pTlgLfaIEyZhL37sAp2toq/WagDhf1nu+pioQPm3Ex3QDDUzP2vgFM80ScSgTo2W
+TIJAuGtAk2NdTv0FkouXNs1tgi18g6fSVKoB8LUWv7grecDatl6drHEblqVz9ss
K+Z9XbyUjaUq1mtSqYFKG5hLfvQ+zBto+He+GR7DwM/P1DcRr8JfPClxVHwV8/Fx
vRLFVFUSKFWVtm1P6/AST4OAWD3vYNZV1XDVEHxDYiKv7DylYlRuZtIwgB8Qb0Be
D4KgHMLG0AZSX0BQCgtAkwjcZ/0NzutTjwLpQrli0HiO83V1yN/0Eyt6qAzYp+AW
86Ed2aot3YZYZwBF2bISg2n1WIK2Tt3d/6p84wCaEV/UzC2rBKbFpDOuPvvW++ys
Cl18yNJAt+Wgyj6fVakSYrnB19f3GOvFOEDwF9ybdDui1ptZDxDVXbAN1p7MOQ7J
dhOrOQkuDGX24vBCCPczg4Q4MyNjRMdyW/m/7yKOCKcShaq1Wgkulndn35YVKqGw
Bwq+Eo02byoskxmh/TefkQBZUY1xR2UbNi1glVkOOte4CdO9HS/kR7lONnijeNMU
CTg7SLziUn2uSluO7mk2o5PgF3CI4U/f89/d5vBP9FmLj8qRUxZkLVSyrNltg3YP
H2uf2qme/+bFytVtlIs2MZoMBBKOSopvE/tJLTKq3oyB2ojv040USahO8uy1XTbR
4w6loffa2p9lfzz/SF02rdigqfw5si0ExicSq05Yj/tiOnGezkS86LiHDZDVEDyF
U16vRQTWFwIBMxowMcPfbgy2O0TafAQjohma0NL2+VFq1e20nl9qgeisvrPqQtDw
UdDmD1lEmZ0STKAz0HL44I6JG4N6SBlRftMszRtilp6G7voyS/LG4MF7kkZz3pMs
CZbA2pMia+Hanmpma6vsu60qlpnL4gWz94xcPdA+1L3jjk6gUAnwBwdegk/M1zY9
cvl3XUimJ9p7MQTobew7iNsF1I59P/H5s+hVjEGTJcmYOcDrimOywgIEFUVvArAn
8I3JOCoi6UYauwd3Wj17aX3ymx5STHeulq65KN/dsjBCdwPN1Zf2tBew905PPcJG
4/pHOO0R5s0VDZKCGpXxUBj1IjL2Hu+1j5c3ll+fOQbDcaWHSlNxk0Gqn5Ys5SUb
NJwLllZmlw6qoo1MZeiKU8TzIRDLIxkONqj6YHeV4kgPUXBO7Gu1nd20nDH2pS4s
RKYxNIKSssScyWjYu+eY1BustHXfSgQZ1Fb8FfzN06oGWP38kqQ4G7G8IM5wk+ok
hWCF5C5a/qJfnbg496dRrgXC5bPiZYcg8eKDZQlvkHQvUxP8IEZkqN5afiu0kcbt
QXUL3pUYb0O9FsdZycyvQxaW5fugjfPqa5nbhk7vXM0N/ovf8G2YIFm+ZbHN3Q5X
wU7qUaRP51kT//bf/F1BKK16j/CvnGi02wiy8HneLxpn/X7pAC6OJfkllTbfROeG
n3Co/Nb1vmGrYNCGvXjnkpOJp/aG88hj/lENZO8CC1fq05VHhvgJ8ReNkg571IK+
PBvbb9IoFleqJOEH8WmOX/5ez8ZTGVRVkEaNX6+ECL4XGQoOrbPfMv136Z6gpPID
JRrPciUTYZv5+15rCkPfbG1/tQadGvDjv5NHHlG2/rUoNdTEpkoBBdumxwEzFp7S
dN2OeN7tBjzkvr5aD1BXF77MB42s2QzSq7Mgj8Zr2djQNpvD3J4Gfnpf/YaTtaJZ
vfUQitji32viplHBPx0Q5epHAt98PrrSvmGvjqyuTPx/vGV0QnCUbrKEywJmE5Re
jPe6ZDi+u4M47379zQDcidKFRA1JCN7LGqC8j6NyqAIeITdn8niyqD/KTUFGzvQ3
EcKStJGBG0vbXir3Ms0/r7KxRE6nXB50jkTfhv0VtFRyTw8B+kSaQCh7vBWyGD8Z
y9aodq7cryYUUyLd2eT6u/Yi//U94hrkZe9icPzlRAkZ4iY7sjmqNZuGJLDON9DA
h2yJ3ENUro6p6kgvwKZuSK2PscFVfMn1jCkFjgMSVGEPg43AL5YvasTsuzvt2Ak9
aaDkV1h+J5/Wa4YnW0pDvLT8W16PEagddpi4fMFOYHIxabV8REMq4t3U26r7CyND
/weQZ20ya8xvPMZEwn7C8rQYAgzDMyxY0srQI3go2nM2rIoWN9+SxqWMc7WoFlXx
S18LvLNDLuMXV8ZSwuANvZb8UFy3fkusObjUTPi8vwPcvK9CWbJAFyh21Kg5bR8r
xuyzkX/yR7tBwlpsyTcIT/QEqUVO+ecNCvoakv2iciL1xKEt9KCbSX08NlWPTM5W
TmvgyM4Pks2yqc0wD+GcfqGi9mp8nEBDuFFPcAtBjOPcHFuTOr3RfIQWKa2OtJrb
5XKmzJDuDQ5MYaOe6a/o4N213CS9osmROE6Qo6vbgp/+WfjHxxaCjo2S5mm5l9GW
VlaQ3a0ehKe+ywiVNf0s/6XzVWt/fuVMp9w+z0feX23ioi7+zE8jDYtCMejBNnY9
oUZW06HaK+oTroEWk8uGashiplxl67kSSTh16/Uo0UDWeD+XW+n38HfacgKnFdxJ
nCV9sfYKlN+irH5C6fUGzfxDGc6i8uKQ4cPMvGGkIRxAv6C7enpqVBgfE41r3RUs
DOhWnmGNMs62oqO2l75f3jWvoVrQCSjsoZ5X/gfWQzcKQZkP8oPYkWLr2eSOh6tL
CP1Q+xkHVWwBjV/XyJOWLRslh4NxFq6dsaAzPcceZJwmUHuNEl5s7mv+8y70+iBq
+4x16tx5/ZLknBTZCqjWhD8WzeALVVotRvAQtC1rkRF415YajFY7Alnc204ncCHn
XQA2zMg6w6CPRf7EhoBk5HE8ajxEQVtd/jC2KyhS73ZO96ZYGsGxL/jfG1VSn8yY
tqMqOEiOC66rl6vTs71iOth5/FB6s6Ne05mIKU2lqjXu3/JWqRTFz8+/74A9nVoP
SsAYk1X6rUeACEY8sdh9TrB83gqyIZ5trdCIpyEIlSc1pPJLfv/jx4QhEMTqY/Xg
aJ5EoY+QvzKeXS/RCfkFpyi38HsnLFPf/GGRUgnChZcraPPXNdzNqiFk2+H7fqKo
StBM8pSzCYEZf9FATKDehxx7Hv0Flfb9pTA4E4zkHVEwRgl62XW3rJKuPR8cNSIJ
oVweEYC1n+F9SZ8K5Itu2qV/iti2XovYffVzXDVRQSTGaz3tfehBchFyFbxpSO9V
/VFEiTOyiRTKl6/isKmEXvZ/HtwYWGtBajJiQ6aZxk91C3dsK72DjR9aHMtAHoGF
AylSEDxoGY+vIwwWBI4jy0WliQ0XRm0ETZB8E+/UOglneR0QpS8d4QOwpItnONg0
zwhCyv4125MFzWp0MUWG0/LWlrm7bKCE3xzqVll4UKMleGd+2eYcKfW36iCN1bgx
Bc4LHbxxVYxNZ11opZq3ZIvSeA7JwQqOwb8OV0caIsVIseCf2h0Hj76RUp/DI0cG
xZPBHigGfEJdCPZTmi1vaFCZhaoYyN4S2GJBXLx5zH9FycNd4ZyjPjinmOcTYPVT
Dz6YkzWmErspe03S9/iKYB1+5HDJzUsSKZRoChfcEbvCy9hkAI4js9H19/YJNejD
3Kxj7y7KdDUyI/T/xzibjEkNXGbSfqoFMO82tGB1C+wC0B3rrUlqa5Fi/DHqL+Eh
oUQIIhtvjM4kh5ixSDJGRtO1ZQJ+90JPJsGgS8kbFds9Mg1YVR9cNDBo18HgEoAx
9P9yg6gPVFRq9Q4fZMh3cslPDHCXuGxQxbbOu9szm/69KZyFWZZtoIkiEI8tKb6v
DWVR8xnoBziZ4a/NaRSS7aINsNpzqxeIaJ44X2+vVqnbApV8G23xIL4kU4R2zVL/
vBQ+Ee6xETuDTfyhKxrypyuf3zxZsLU7vuUMdHjlwxnSiWNm+MkQIz4UFsNIr2pa
8TOflExfKLknsuSU0APojlDoeqHUnMtOdUeZRazop/2tS3WsVxftMIyG+LrBsSYB
oojwzfxawLUYAfp1Wq7+vt0GOPKDpYq0VmGuh7bsSb4fPkwJYVi/NjD5+DafqXAt
vfe5znrrIHnkjG6INzgiW8pHDn7IJsikhUp/Aov1Mn1ETudzPYqxaoH7As4w+Yts
mrKJ8Majx6LU3TWM6oJQxnF5gMOw/DCuPuGl0S0xgA8Bam4psVZxN3l8Vz+sPYSP
XYxuAW9Myr2Osg/H4HaLE93xDK3+hJstI5XmHmX1Es63SvUu5wblJNsZCYRDkFaV
HN1jXbvWiNUhTCed07wK/3btoscXdD2nufnJyke+cPmFNE0nGbPH3w9VuApjmd2x
YxhXWVqinDzaLG2Rt9T8yn62+NH9Z7gWCefiQgj11kzPZI0f/YyWTzj+HZmBEdQv
V8KEx7AbK5QZceaVkSrS9gk888GU/q/hBKOIfoG0XjPSFrAl+FvQFGArS/H+Qa8J
9XlrA9zKC3jhTF/v76Zo6T4tE6ytFvt6b1Y/wVV+JRDSjdH7YcQQeTUDYgfjNOje
k+krx4QKEvtiSme4auHByasonTiXeE1Y1KB2zvnhJjCF39rA5czC1MowuiOBj5Fq
F5L11hw7H2muuaWwvWskspBgtouLJnRj41zO9uVRjEJnb4onTqHG8I6dsBwpgBUo
NtGYk633f5eF6BJb8gzQhJIBj2yMtRQVzPc7u91bfwDfH/lsdMoPqMTTF0A80dVx
/XOI0eL+jV2SJSryRSpHpXtwl/uO0zK0951Jx10Ge3/GVfR1czhU63mxTAoR2Ukz
tMVOz1e0DxEAOYDrsMMNoj6MANDOLwMqlOx1xK1pkZ7admX0X+88RVQhrWAWrT4L
zwCrOdhmrjcryNnt+Qoo0As4og1RFLOONZU8xg/Swm0mLj1fQw0pK1avqyQPkvxQ
HjG9Z2ll1pGjpWbz7Q/LziOc4O43y9WCn5rzFxRYZSl8BVgOa2pIirKNbIsFvrkD
xpFbi3QruHqu0T0zTqprcCPOQ9Q475ESiPEueiEgQYShL4jYGr/SYewC6oR9m1v2
X8lt95XJ/EkgANQLAuKsQemoy5amdrzVnVAdRA2E65SYrDeS8D5xULDZDwGTzzte
GfFIl0J/zlmu3nR6gIqA1Kpg9l9qQFzlX5w5gTK0QX+S1s+aPearFvC9mxQcJuSU
Hq2ZmU3jW+VCw9I/QC6lZDFxp3xT7vfuXQDLXf0OgQcgrcTjmkznkOuO4t8i67gh
kej3vjmOi6kjIhktvuVgiuaWe0EMwHHIldSBAIWClOnA8ZJN2YCV7+GRASPD3mrh
fw4TcM3w7cQ0s7tifOKyIzkltUAD9B0OM5lm+BPsTdiFyOIutVs5+Ots2kMzBtSQ
ObnI57hIBOE+zyajwcruPPNRI11/B8unUm+9JstmGCCGgnAuxUAXOk0tm77CBrxd
43HOrD3f1BT3U9OiXo8GMTem3Em0N0haGibVJP10Huin3mrDOp5wmoClvziJzQBp
+Q1VtzRsZuOsCCyW8yzQ5gFkx3ojW5rDtj8y0h7HUq8zdo1EaYgX38IVS2Wd7LG3
TikI8bqDLrQA5/33/Sbou7Gw90vzkjIfXzmDBPNuJQpXoG72zA6rKuhSA1oy1ZN/
/DC2+35LAIjaFKXCK3qH3fkxPWUBXggqvwEmhVKqKfD8vMO91EiiO6YXrlvPlsKw
NE+tkLp3PHG/WbaRL4cqF7RXDjzefu6MVxIZgSUx0dcU8Cr4iD8AezqR+9XlgUdd
oee8ZeGxM+388hEc2Z1x3pHxPlQKz52IVGW2fmHx4VOo/FiLTV3FkPNmrHuML4gI
ykt/ztwYEJEYX7PMN3DT6GiogcSbczsiVz+By3hi94qx+ZCdKty9Mu7hiBtoULDF
odJBsl2NbwjWe45IgO46EXvf9tKE6dKpJd3XVVFQ1ZTCrn31ZMD4csOhfJhjEI+m
N7vswG7Kbqj9NI0q6YJaT7Qk4BMxjSicESdA+XEUR4AjIzkZU0lUKHjXLkwKGlb1
SZgE+OTiYUreW0PfZl6IOVSQNpFMs7lpOkOW3KORT/CdhHuw8A4/1uMwdsiFxNFe
UeL0NsOKAAHXCK+fKmss1nI5R9R15mVJ8KAGMg9KwoTdwGGeKbbNQR14NkXcfRaH
mggm8NY9lVjRQ27kd7TVq77xLHMmV0n/HepvHN+0uqfEXEXfV6aExA3tKUpJMsCP
1ZTxcUkPzJTsEw1ZN8exGhuUKWezPG7rxpxDZiHh58I5Aq/Qj/IXBq+ub5VV3Cc/
huRPzIH+kejZEYYfB4by9kK+JGDswDHFD/8O9c/k0WF3eveGciD5AY6pSZu/hxsl
mEp0CWtgU4sboXVco1tbM993isFB8VXQKcPRyQjqx2/CqUqpKMXBpcyYmJrbui6H
piertHoXzjTSXsu+fiFyJybLIh/33NjoHTaqT9sFm1WDZ8qDjRnb1dIWKqRYYKv2
RxKSL/qi6UYKOXQtpFU7wnfBWErkoRkKJUNiYgCkJmBYNgluNCPvAm+UsPKo5Gsb
Ogac2UJ8u9x3/0CHYIMBLbFhRU1Jy7MVmArkZ+DnzXGtYZy45fHz86JXncd7j8na
x4d31Y5MyLdwzoLRxY48Izyyoh4baHAFHq2s1TkT3NDuPCDZqsAIoEjPDdnJhqtp
d6vXdMxxzZET9XPvLSekbzqFttdftuQXY4d/G7hUTBHzgUSXz4P0Ab6aKsI4XeVp
++sju2VkVE+hI0v8sY21jiqJY8sP9UJjh0vfndvLOvqsVC04f6ob2+pK7SjGTAsd
dbEMjJWnclg9kstTF0LuUka+aAMLJzClhxNoiI0cFBOlJswLYn/oGUbzw70gMyZs
E1/voI4J6z4BYZbxWCggT2iCU1puTpnXbE4dvowGWTqehGbzHNxjJmo/gMHCZxPH
pFiXq+wMum74zqP4C9p24vVUwjzRHXo7Gs7vaUiuCjGqbpx9f9Sd5wg1vpnTP3lo
HcqV9KpyhbnGnHVxlPBZIB0Gk83K3zhix7zKDvpP/PT4SHIEtVNUeH+LGPuef/ag
ahwSW+jon/A8Y76m+FjVfDnyjVl+LI1msIOciVmkiw7E41Rg5zNJyVHngEzUcNhw
KDcwskkZLNkIP+IYMbTuHt7/8m91TBhg/gQIbLwZKFQa7Ch2TL67emxLwnuTYtC/
dqs3FQztboQTM/mEemHSIt2PGIa7eMTV0eXKNX2kC5RHXSKFGuS0AS/N17H0rV4R
neRe3xIJQccAh0WzOmN+B1gbNcX17jYfP0QY9RBeCPDOQUgCi0+nl9Km0NooU6It
xOevSjU8uACZdPiHBPOd8FSob40RQ2pniHbCP+aME03JCoqW5H3Zx2Xtv136nwn9
bIgVqbloR3/Hnmy3ksY92+F3TiIKzcZRP0XE6cfP9WrgvvpAd+Umd32bHu+7/Kcf
QkGmrXikhj0sXsx1iQisPLwf8MZXAFHvvL7Bo5L7pSWxx6XB2C3KP63c2BRxc2Z8
7QgPMU52+Ks3pk/xjPCs5m+xjBxTasGrZJXgOr9fq3Brivu8PpadvbQKKV4by0fB
2wrOsh1u+3dXdZph3OT2Wg9482v5sUpSCUcLUe0PM7kSLFX5FvSLtBgw1IA4C9dk
wVNPGfyVQzJ3Z+2tV7StFeWpg+5Bp5FzhxvwaxHCVHM5iSWLQ1LPe1cdHpp2H+k/
7INsxEvvyOQUuJ/rl3D2EI87/JKI69ygTp/0H/rLIt6BbUCpxx4o0zlks+ZWihr8
YoD+PTEnyfGq7H2Ddi3MsiOeaOoJmSf6QepkIHt4VzbynHvzCHNaesVy98Wr9ozH
IWfBM8pzP5CrGNcyEn3RX7WJZiF1VpnkjpbCLUthgP2uIT5TrGJke6AnsK8XMHzU
I9P9/ZAqraYi0/STqAEievM3d1SDAKmwnIGTjQWVVFYdHb5sWNXvHsGgi3STOu9Y
ZwJ9/B0M1BhnUX3VEpi0P/02D3hJ8X6SPfoIyhGISBVyze7fAMrmj5Nuf8l2ovpF
fWqgKDH7IjQEqRFtcO5Vxr1Ew/iadB6Fu5to6Je/8BwXKZ+lAR4hvOzgQhldIN6o
WDirISkcmP4t/NXuZFw0g9FmtggmchZ7Uj+NxSrNjb6C8Iqrp7gK58wdLTrdsnVH
Qd+vZ3UecCsIBAVM0KZwN2ovojBIMwA7+6LQ44erMag8WaoXrOvljg68OLFc/DFd
XEjwD8g2JlSjR2gZTxgOTqiL6+toHaz6dlDicQ5+cyQ58+gFovpEuolMR1/z9/xt
b7Xd9YpltIbOLoKNijjE3tzdatyK6IP14WCXn2IR3CU2i7C0AZ0Cu3H/mDLkUrtR
S2T3DE/APqPYqWURoczNHljdrgWu8KZQJD7+nUBXudk3fH6hJmdBPTbnR36XhtEI
at1BOCnmR/LY/NTCPYblDxmsB0zhoNcuU25PYwFmm24bHpOh8C9kdgkFlVNKT7cW
LcKWtAFHLycD+6jPpJlGidTzHc4px3oL3rsYiNw3vZh5nw9a/lWEMm4v3IxZm9PG
myxVoZgYAPCbQtbskYa6SqdEksV3nBFXdgI7MuAYXD677R27yKP2EHFY8yeeCRCw
eZATwsiOb6aWgLCmxdsy8+z+d5kuaKKCG9mqXwffIGkEsxY0QkYpIZ76grOgmksQ
3Kgwbw1AHU7XujcXI/NmCSKLTUNlnzCtllyBUyDlRXnRM97O6NpJHDAMaMHP2Nnd
XbjpNuiYz77jn04nhnSRRdNi7wD7GlVOd1GyiAWiVqoiypH/toPSeN2qsh/uBMpe
Aunz7Kly3jZjqMoq55FBkL815qZXqCEbjfHEC2lV8swT47vef/5FPP2PCVHpDrix
F/i1jb4rtACmXozFt2rdU8mX37UiMmdAwWPnqU1NqYc/doCwuL4Rtvyc3cU9rUAn
VQGY4edHnLsSEmh2YZ2WiWmJSCQwfVVYU4Jcfx8Hy4n/PQMlnUseiXUUxNUaTlUU
3JzPbEpveiPMq1oCJOuqfJ/QdfdB6DmtSPJEPVv/EXIYYFjImn1AMTl4d9NAdJRW
mQEPvB6tfmbQHb/LYrLjBAq7LSIZPlyo8Mdp4ZQiqIFa+I4ydL4GCxfAaNtlvTlv
nfE0eQP1pxlwnSc9ASHtWuuhjqHOnCwX+5VrzbVwf7nznjz2faKUKwf8YcuOFFHq
YMETvYLy4DtIFbDER901uGB7y0IoBxUJBeQscEk+MU4WiNimO3kw9lrRkT9JO403
351rdCzu6yH9xD8JTXpMjLM6yYay+RYzQJ8QJZiRA9v4RhfjSKd8PfAzdFHfe7GO
svidJTs7wIAETul7wAiAO2ZiASiUUfIsMNvYlJPPsgerASu30rRoTodIWeWlh2QY
mYyoJ9NXrM1wdFWMlVB7dHNj1gRb2J6A24k+GaXC1CqsOb/pbymUW4z/66qTMMsr
9DzEtQ996GTJMBmYDkWBk4dfloPqU3Q3b4zWOSNyxFHDHgoBlmv+t7XZsltrfWk7
e4b3OKTNWSi29j1jthRqQ7vbpQe1212b0yO+WzrMAvR2mEJnjZTCIVQLecPF8Y4+
JHgVgA/l1AavQi4w4Vj+sXhYFP9pnnhA09wOUbgy7stFZPha0Fr+rJGCPSPDU14P
9B8/Gb3XkVw8A5p78hfYj1ZLatKLCoerV38A/DORQy87GjsFz44XUxteJ911DiZB
Xt7Ho1z1KONlkuiQaIJm3QqEB3Wc6Hi4qBliD1BcinZIIjq7AmnfRLQAlhcjMm1K
6Q3PBWhJ+YrCq8+umG799oFAuoP/KKwmrJ/lula36eGyh/UMZSAojNvAjNpMNlGy
mxyjMw0PGe1iWoVxyLGDGYYfyfj2SwmMNQLTxAaQVD5fvKdJB9DfLXHjb0NWRCBu
n/8XAeigjphW/07a53ayeJXCc4dekp7tojA6lHlSbjV7dygLkm7AIbuvppwerq7k
vAiMY7wCZGzdmikqipmbYZqGnzWeG7hbnjesHd+sKBZ64U2Qh2iNnE5fMj4MLlP3
J0K8S3aeB2/ugBSk+e9jvHI2st4cljdljzPMNdDUn9bs/X3aPJnJQGD+ZtdmmwOG
1wg19slT3+dHIs+rOztCCG+iw2MRO2osAqtWG/ettjk8NO9lnXuIZvQjubSkKEsg
W7HSM5yka+QzgOPQHCvqs+yrTTVC+1ayg5rIZ81nskjAaXa+o3WVjbs/YRrXx9+7
LY5YYHHn/fe6B1+a6hObKf9T+iOJsZfQHKrVORoMcoZ2TdnpFNJe3ziFqxcqezQI
WUwZHmPJQhcLc3gW/zXdDB38pvUVmnhUCM5Si2/mN4u9AYYzED5SYWJrU4p25Y6h
fFwpg9nDux0zkqGNU8QH0OQB0s1km8r5k6HN850/w3gQsRdRg+Jn861lDpnKL/b3
BgqrCv3ZykI+/JaWeChBj69Sqy4rzu1kFPshd8ML+5xtvDglWrJqUa9m88jDyOWM
tRrjsZaUcLz7miI2hMhCDPcfdefXkGR16wFX22ZJVusp650h8nxP7slhJcH/U+u7
ZAEPC6jLUM77w67upznUGnzZB3ZeHstv6qjg5ymP+uLpsz6gVZVuS2oWwIeRiZi5
FlSp6ZgRkvm0ywTlnGpZmpecX8wQZEx0OgVONLoq0tZPOfJAaDGf1QQ8VMeeRyNG
nghWZpSSGzmM9HR1tcncNMtyLg470G33imoSlG29oIwXeE1EpPFFe7f0/bCMKpFA
rR/kv5NDp5JC1FGjo0YaiXLkaqMeUXR78+v2g0g6vEYOzszHalYro+1NMZjrLuyE
T9Az1/KvYfWtaUdqhfs88+mOjtrGiWPHkWwaoQ21PAMDia5y3/Yp7KGIZFfDwBXg
yfxbY70ovEMcWmUWgLlFjNTpiWjBz8jRdX1NRUj3e39hzArMgvWOFnC/2ESOhrnR
hZWHILv2QO2t/j8eTLTPnZXz1v8IkyxdKqYTZ0rNtu0J8LQRxz0/7o/D/6Y/uBj6
mNbqEtgwVb3X4eajR5VCECDdpjG9dhUpi2lfBVv2ke+Pn/Vfp8V2+ZYgZTS89rDH
kgr6PZxvej2ZtYymkM/W76h6FbhRrQ2X9eG/XpIckByNvFp2RMtZk5wv58qwKuwp
qPyKVe+NMonc5pgQVsoyRykz2EUDaUbcaSFdBjMIbk4mmSIz0WLbYeCPzcweSI+C
cjSULx0aHYP/KdiJWFUwQCsrjQxv15FQWvMQhPLzSLN6vo+nc5kj11+3WlMGhwwH
eJJYuLq+GyjRgI/ZGCxU+hrwpIlgMGCpLjf20O5kEiGaAmBlkFLRlxUhYRlp4iWr
lPg8yTvJhqypmje2gHKjT9eqEUVc2ZBiOQWMQxp2Obko96S7Wwbd13sMkXS0hCpQ
25KKjYZ+Cfh9hAzVrl+1FBcc5XIS03JSzwoZiGZ6sapRMXbCUA6ZNUplp1YGzB2H
EFSz8zwUiEKdSo36DniUMVjptvXZiLtS4DLt+dqocZCzn606gHjnRg88kfSFevk/
Lmua/2aaIoPBqBL4oIm/9Vdx/3beeqff+JIWsdMne8Y49o2bNjoMtr7QPzs2Wykt
OX1Z3VjJgciXallBrFhUH4CuIToujy6vBXHMpPqKDTQs0RwHhceuV1NKeju5AvrS
jCFXr3Aq+M2sW6jf0r3TTPBboFRhGN1PLhIUUCyVBD/OvGO8qJTgZl5iiwt05mhl
6XDZoC9++CUdVQxIVwUhKZyENWeBuegCzX5pYque3OiC0UIqU+ChKcwFUZaDRkR/
TmZ2IqA2/d9EaXjkeBF25DXpEzv5taAzf+mKlyYHeMnYZq67QHZvXCDX9xh4mcWh
HQWm43EeuDfic8RqtivLgd43PjCzlkXe1mnXI8QiW1KbDstTByoOE1K6R+xQsj1M
7D03ZSyIe6SN8y+4Ts6TYLrPpKGVBsV3D14auAv+Hy86BTH9hIHWnPldlFAuC0PE
9FDBRbZBvfB4PybgFpGkcBx/ld3iZuKbO/hhoOAE/HUbJqvQfqjKhCJa4/zCViGz
8KT2d882IRb+hpeUdrTXvL8SWs81SJhT+0bVix5v2fRO12TdljXZM6bv+eKzvTES
WDO78Av/zvD2u5lbmV06OPaQWoE5iWIKZv5SeZ9wgrp8kAG9I3g6r/0jtsq6GAl6
dIkcSA41BXZ3q66ywYG4b9Q3vVHW0bRsZ52VsYIxgEmeJPNHhJS/Oetj6pjNKUpe
/Bfv7329Ro+5kyUBm8u9HaqCkHxPSRv+T3Ysuz6CAJiB4T1FKg7bNV8uMqpM+EXO
AHnspppPuibwuT44hUg3ssgKK7PyU1XVoHi6drcHRi2rENz8fqWsCyVoqSxKYhUN
4PoQ871VtOzlWwsAslYlYRh53MMLhdG3uQJW3upl0M5L4gWclmppvG3SEuwgqwm7
1f1MoFKAE+bmJ0yxq3Z470NNvQRrKidgF1Lopc2KYb2aV3aA2OlVHmHi2YmWiHbj
Z5Kjz0vQT3dmSFKivG/x9OM7bjyymjpv6HV/faI0FSorIIngyhyZ+gPqzEycFJFt
PjHAMQkYzFkedaFiDxNbgauAxDPUZYrQqSlG4SZmg3qZ5AS++H+dJQL4Ubs/vCKI
Jv/TauJpG1Z1KnbIXE/YbZgu3i0hlWd9nXIONYcVCI4Wegjy5Mjxe0DIRNfffzvr
3uibKnrHS8Q/HmpMHHiHrGf6hkgc3BkNQtFTnk0Bacml9m82SPmN/pJWuHrAUwX0
ENic2AhMH4SEepQ3EnUOSUiqQFFdJwyE39ya7e1xjcx/hUIiUp0JekrjERVU6l7E
B5IVPDXCfDxhVHQW9P6H3MwJSsS0Y/ycqdfcme89RrX1TFTRmBNGlyTS2MeoyaPf
0ec2IDM1uPqsGHRGLCSdORoVyZD4kbHWeog1sLMoMCpNoQKb7Ks3NwhZJJEVkQZN
IBmIzUArwjOP8aNpkthqe7Eh7xIIID9DsE5X/J+E1BCbTIRqSiREAJr541cP/6un
/zJDpJnCPklinxSBIweKk+RbfofVRc1F5nJnkPxCYlYdZqGJP1psiCWDgUo77OvF
ycNi9g1wddruWeQ2/0/QspJJr3JfDx27nKiXtFd6e8lmofo78TK0hUbwNPoFBR9z
Rg19dUFlkIr7eaxli4ALczAoP3cgsVc7tpBUr51koIJoJev5G+2gaPD1wgSRPi1E
1HcoA3Q/rvrhGpUQjtcC5uKUFKlWJLEZFYq5zWXB9urwEILupX1rBQh7BegXqft4
1RGagaonZJjYvro2q7ay3TeTokF3SbLh5iJCKY5Jlwbfo8evxxkvus7Q+DY8FVId
maxBrD2Pa52aBwfZ/8Y/lT+MWBgIBFDtM8s/b0XkcsQ42k7hSqKF5xPhDsfZMfgS
/I5oib9ZCOXwg0WpN8XEKgmdrQcAIGaPAe/Rm4jXi3qEDf3wXOcAwWbOtzQQa6Gc
2GmPW3lR+8NfL+Zrx7HFT1VZyRkZbjR8tLjuz8At+iBCmryK1rjKUjuzNdNeKrG6
be5d8nHOCw8c+UmYYMRJSIuhA8blzqfNDduDQ4UCrU/FcHBGklrY7bZnUgYveyum
To+gr0CibpnEwK7d99p6VB8QtDE02x6236WuapcyofLNmQtUEADQlc+ELn7/41os
DmRDCqbEwtvhukmzBdY64JRhGD4TutM8fikA9+3tz9Zoy9muX4l5HhkgRhFcMZ0t
yV0/hj+/XKJV+6KuaNVi3hJ8MHSCeSMUa/03wUQKShkUmC8ZtHWuksMsApfQhHpa
QgKuEe2aTGQUQsaaFJOW7wqHrTY2OabCqSGWE/YoxZl4QKyo2AEtVGPysbokTS2w
Ufg+QaC8AjGxEmkSbPLiiy0PEi2qLElbe6+T6jZXNMpUZaWtSnnuHl3itcDeyXNk
FKarLT/V1RmbAnkd9+Sx8FphNfIW8aL/G3uiRFR+ZuDbF7Of1pFDQ/88X93oX/u4
XeA9PlniHdkJ1150bKZJo1n5ghuDyaKj/tvDHFUmg9YsmUIxrzkHwNTRndOxF3h7
Hkc/uEZNVza3inEdgc/weiEwoh73RCS7zqBjfONlKE3Q3MVj0sN2Ikn68nvcXmiE
tgWI9JJ2rEvn+pAjZlNIiziUWoIbSpc+4RZFzcGfGlw1wJ6Qey8yTmG70C/4jDRT
Gq2OGtHhLqx9DugLDAd2zcuA/JMc3S9vcJIuT5rQRR23GY81ek0wsxbo9rDNaz+e
wUsJid/ovHlIwH/yEMVnY4PaS28VdFNNiIePr70ywK8o1YqBnElRyENgFTJ3VYk4
m5dxrGKPHbQ+kHURUa5wKW4tF1mrca0pDrPLxEZUEO0Q6XIo5Ajk2pKMeAv9XTLa
OT7qkwcX6RPRyN6S/crLmea/DPYuakOPxZNbqRIfpGSGewwBQBcqnRujxcVcbsXd
jBBbq4ByfSr9Jcs4G52Hb/FxTVbUE4UmO4hIF9RZJfrxnSux+1U3w/urz7iemduP
itNb/6lWzWF3tBWW3PV1C/RDNJoi7qUDQRNTkyHyTxGNKvM+eHvpMW9sw7QL0Aae
pcd1rbO9XmbucYCNReQfZtWLkpmmzrlbZuDCKKVdLHxp/srQ7dk9wbLOBZQVnxGF
ftJeIBWXqCeKxUpSYqk0qgvdSGQuRk5HNHR8a/JsMaLxTJVi61WYcw2958JHK+XC
xq2z74i2EqXIiNXMrcbjt/C2lXhaU4ivHrZKqJNh9b6wZcTN3TRdpSux/c0nLIDv
wW5hgjaO50iUhD/j5U/nEit6eYVK8QL8aVu9Q/8qQDPEQJpJ6LvEDN18Zu6PJfnl
ylUwRmH+CePVNe/vWH+0oDjmNMOGzy0lS8VMgHl1EwLw7EVlpG6ugGveZ2cqIOiM
EaGB9MSa2jxrqT97xdJyRnd18VlA35i5z/CM/hEcQh7ach3oC0+h6w1k0sAmzxff
/lZv3sl4tyhRogaxYbktOrqU73V6a3/peGkY0mv/Hn2WNKsKH3dEyOoYdkxAxsO4
4vmo0g0X+BsB9F5PrApEfzSXaQUp9QU5uQNLSWxpuSeM3o2ItfjfOfO6neuRFfeZ
1IHqOGnNNjbxXnc66oypJ/TP//nzIZ39OzHhC4/J7CDA1EquL2MPD9uTckzzaW+7
3oicGcauaeegyvrME02fp8OOeTAQAf4SaXy1sR25wyjK85xl1qDztLZFt4bdO3z8
asXewPu+DeBr4RgWAaev5+ZlnWRczXmVBegPfnDx8fQCgPaqoxRe2N7vS3RIZ3Hz
NvIY3EETBXHtzAXSGEhGzgvIokxICq7iyoK5XH2rVgQdZtkrvqkS6tQD1LyjUiyP
1QHgcoL69di+9fnQafSGmC4QzJY+I98HfqNGbgMr+13s7ioQmu8fYGC1U6mqGcC0
OKnWyJrQeC/GCIIzVa3BaPGK4+46bJt+g0GgkYIq6A6d7+2kquShxUFXwrTCgoJH
Mi14/tGw7XGfcVXEBswLwPdplX2KOj24wHcRk5dAZmT2qObKVD9yJOq4Mpcu7AbC
+5SZygddSj7WdDOaj08Wh8FK8S4T/FqeAzOcBX/46BO+u2cDKwaXfw31l1uW5m5h
4orzamu6t8y26+BEohvjcqKwAPzsBa8UkDzDaHteH9ko5XrcaxLXNPGNNi5sZnpz
DRMd4JltQlB7Aq7xAZoo73r3SGJQmSwGZ68WLd3cjXnNFGa86xw7ZU4dtU+zJuMW
xgYiPPG/MGe/aHRYfeUt1wwFWEQqttFlY2lAtFwfSyZC1GWrOY9kHDRAFmyogtK9
oCxMmBRYE9eiaSaHwIlx+E0FVOipzgQERoFkzF1Y1U+J3agFgLEVZC4LiY3F007v
symr4fiz8GuDJf9ZchVo+T4NaYK/hgaall5bx2h5oLAQY6Y6L6RLbTmcRF8h4PVR
a5mOa710118BqCTJv+O/0sC0fEgeL6cbCFPB02Q4RsY3XhIhTHloUROIa0Ai3ZZi
pms75/kiAMFO2DkaORtrbhFXxJK7+eUTNjnMh0zxsoXuUC2p8C2+U3pRtVitfxAp
sHmqmf/Wph9Eq/fcGJ25gKFjrqYf9wj9F6fQdu4RkkMNkdvQkKJNm+5GOPfNRdal
bPThjIa/LDX4t12j9T38KCqYFlBRjCHylRMY+x/VVyFHyYD4qM1BBH4RSqu031pz
9Va1whNf3MBfUcdyl/v2kkoikv2s6S1whGYZ2UIgh5ggvWVX9a8MOiEIzABQbM0o
PR3Z5NL9954FVUhh62cZp8iqSJUmYEttuV4KJngZmtknCWGhOJwFRxjewE+pqOOb
j06slx30SBdYnOZGk4x0Iq6E6aQ81jFF9+AubR9IN6djzGXyI0mwvqE9j6lrMIHC
T3i7K2PLeQtQUjaaMa2g0oSU8zYmpEWg2DMtqe0aWvLTJVTZCVg3R2ep+diBYtZm
bKQ/rbSN7S54zfRz3BzjWXjXs02Fecl8WpNPQLqfCiSmWDIAo8iAx1WLRG4Vcisb
00LyQqqSfAU360dgXzY0s5XEF45LOuVOU3+azAHEtApku6ZZsMTiN29nmnjBYgKe
oH1rybI9rsEGmuvLrrLOwrcoQmVPDO02y/otLnFsA0NT5ynsqWW2XWLS+RCNVx2+
sbtidTS+jnzlDtal1nLZk9Z0X/kJBwLSzv8N1M8Y1KV7ilgaXWuvFfAanYRzA+cF
4Ssns5dSnNpEoX1QP3/oS0MluRadzNB4UxVEFMrg8AjHAR76qg3azCr68bjFIDXv
1D27cvrmpf0r+1Sykdtgl8fXQpwSqd20JlmLNt1AcblshJC546RDyr/ilwIkw0gz
mwGOIhU5YbjwVzhtNGT3QWbpAx5fRE69u4Hju5dn4sZl4UXTkIq4pK7OOiaIwgC7
dP+KMR8ipyOVBWSd0uEDBtv5vxHYFGuYB50lXFaF19kFSG9K073ZkbzzilctKb+a
7VLfL62we72M337ysk1/staO6A5n9C9qnS+s1lToQ23s8m2K1nvHXu3sSvG73Inx
fB58q/WWmzukrHM9SZeC31+0l58rXRcaoX3yy4Td+mPhGDgVQvxBO8aKc3PJO+cV
cNMZ0DwXSeaHpHZJD1RtAtUAbqxvdSTFDDRje5CGcQanvnIFflp8auA3juHbSFzz
Av7k68Cgwcy1FmuKeEPZ6qOXoX7JDHsE/t189deSa30T8htnYrlBJMnD4cI02cCt
D4X1lSFex+Dr6f2O8EQyc2w2GoU5m9MxqmbKEnjCdgm1M55m8oIDeIwd7XcbH76D
5ehzmXjkj/BH7Rzi53STvWVBiJQGYp3xMYxH/Hza6ZL53X/dvcVziN57KBOa9ZQs
wbCmcSPUY6N65ybYUrU0X2UZXD0MBzUuQyqslZLUG2EVsju5j58wDUwSlE17+Rno
1z8cP5q+E3IDbV8uYPPLTVmj42FdiXHMdRujQD8VGoJfj8LI57kHIalZOzJsRTPr
LelIw6VBLWRf3C09U0ZAIYWmifaW/meqGLDIrJartJPBvpjpGMLlmG5URk5wTqCy
4KglhosvokrCAtvsmqNSm9BgmQV0nM3yAIzM6FdkJ8m4FobDYkS62RpHjeolyUTS
WqIcuZ6XlsFvSTjTtgh62mzlikIqxVIAgtAnKsSifC4B3MdUSRpFwFixIzBZNgr/
8U/OwYxQ4hMPT6c3BskZqvveVhsXn+PqOxUIBd8UBbPwn2DYm05wGLBfNb7e0mIO
niCCJ8VAidw+HxBiHdOfW1ux4i2rXALefHRSXwDPR62EUlof1QMeqc/wa/ULTEZm
Dh4F4R6m1vwKVchXx8L+OfnFxZ8FZVs2xpALw00bfRcdbiFgovauaiGLifPggPRX
fhelfL7wlb1UWgnYeS0qLUb0mvAGht1SAQ35kjxH4Z3Pwlr+qlxefX1/gDwVDKlq
BnSaDgb9vNrLVlDVAD1gqlZfAr78u5wPykvsN4BIcehV92V2pD6WMXcjG+80fJIb
Li3e3gGNXTiYoQ3a1q6sJ7opRmZIfj36cwuK7YD3NWEyo4dWyTyPIKj4LpyqSYoS
FrisCi/Hf8drbECi5ujKEp9eiNjKaGu+T7M8zPiPM25UKsDNbMXCpHDcRnG9ddzx
FlLQJpS2KcpRzk6tjr7tAxqBgJSKVUTnLQz/iudOBRwaZao4XyGyzm/WwZyxqhVS
0Hmz7o9s5YM3tLdwMpWE0uVLv0zXdNnWiS5653kZdhXMIYGaocQ5Z5CNUnr0uEIB
1se8jKZDVXqZ1NDo5UjD/c+Vh2u19ZpzIHnFgUcEKUVFpOes2W403gLHv/DyN6u5
nhWHp50GE4wNLBQjUUo7JOC564QuR8Ejyi8YuBEZ5XeY8lrKNgCzQpIl02jghyyc
XIMuRobLzoN+BOU7PnifzKBNxV9Hy3ipRVgz+GIxHncw8VYnBjdC2a1EtJms39ui
3GcfNC8D8nKEuRJQgIqfnLC0iYMWABwLvtSEERnLNI31jwoiuRXyM+rtPrx+2U01
nvonZQGMXObspPzGKLw63JUcG4Q+iG9GTqoiK6YpdNISL2fTcN17t11lS8fpOpao
L6JUHIs6NitOmKTHeZ+DTf2CYP+ryWZ7KzAbiDOQ2AQTnuftTuWJrA/NyEpanMQ2
qfwiZ5W/a/vD/2ZUpr5iCxny8nWaHpAJWy1GmUKoQ11lIqBiCzg9042mLTphQKsH
+jNdsfBDr2jB462WNBoQpMdRP9NnT0BKrkuprhgj3Hjk0UhQKihAP6icUZ6470QJ
RSUxjc9AVil8VEowNAUnJ4WDJFQWTpNcMmOt3ULRdOWXgkVMinLAWOCoAUYUIpDd
YkFNdGQD1YW8DjghTGmwk5EeoMl1QiQWPs05k4fWh67wKIqwb9yYyeO1NxjNTo0R
07T7lnOE6UV8epUebzwJ5mEzgSiCVSY/9QaLmCdZwlVIsaLbZSrYaSsGBzH6y9fM
b5nUQhuNl4zSBJovpAnhnj0SZyn78TFxjFjT7whav+C9izp5WGsJGpfLAoMZXyxm
6zvZVk7IJ+sL27xn/683r1209+myqwbD6/Ec7GbUSinu9S64hqXtsGehP/cPFOtS
uH7XVhmfu0RJKgEhXVwG/s0xjpAD7wPtabPs0swe7y0OoycCup6s4y4/3AxXrto2
hrjA/9oGUw9dEUJ+8U16vJZTp61JOj/kVsxo4yRk1HpUWbqs9pPSEfC8QoYeEC//
391GMBeK8q1SuvISiwmtxze1BknMtiY/bcW0W+2zPgL8Yf5tearPwHj8gPiQ+JjL
PTkENcLHJCg3Wem7gUiulNMO0N817U7+W2fTnKhgF/DdjKqQbE8dUGwDWmEWldkk
rt6T3HDbFkLWzBSlsrfMRR4X59t0nDCMm9K08xpwpwhvmV48uR1N9QvQLllFecCd
VYoZ1BRaVqjI0Li5t3oN16zlBwwQS+Pg/fDJekleQnrCYHMjRiCmYoRF7UT0WQOO
SaftylQnLoZWWB0dJ/Gou3u/x4bdYTxlehpKdtUdyVCZkZPNyb1LzmZcK0CfYh+M
P68e0DpfM/yICrlJnSx91UhIgjrqzmZabLhLBsPaA88xOAJ7lrVUZyADjYagf8eJ
4dOzzzibQoMfG2BjHHYiDL3MoQCuuoKcWLej+Z4DV+NGxEnqSEbqU3s5vWUUbQps
UT94uzDsp4h9loKUH91gGqS3wMPvISjXDiEVdd6cXt8JBnawEhoJljZf+u8i8Plw
hh2v4fuTrzUouIC57g0iW5ykTrJigxfMv5joP4ZQ99XbEnQB4BJjdYb+OG0barh7
GCDfR4cTyezqFt9EPQij9HRwU5uJyDPE3Ho9UPaTGqjHmpECvXHtNOLVxTXSfNga
AN7lohVEOhAvvyGcg0ZWe+BNDRnIOuSWFo6skmAaZ7FrXVPVWk960Km1QoBY/6zn
q6PaYIJAaG/1gXOTOPZXxA3h5HKjJiIznr2EXSGBjX3Lq4W1e6NvynK6N/s/8KlM
ruwRyce0qcV0HpggoNbsfHWHKDSa5ohYXKLfq/sSkqpUx+M7uNL/LNyONFU1QMVL
oejgO6KhVBBzupd841rwmgMHIEswm9WWu9KLuiYITdcFyKY3QYh7HmaI0dKvIDZg
G1o/9LVyd6lDl4cZNAwu2BP+bcgDsYho8WCVLpJUHgA3dUx/pkF1vePq6ZVenolM
EeaJEPHpsCUQ///Uqs+Jmnt7v+qes7QxN6rRbkrz6fw31tiEncOcunfXO96X+JGF
/PuwZZr57gUVHp/cgrUgWXs5zeFDh8DavCLic2z9dOoph/ZEXe5YvOmoh1xIlxtY
C/uqnIp6/1bw5SMq28pHLrjoytAf4CzEjDN3MZvpMNDhc3XyTi8CAJkuLzgmd+40
xep7It5pwHMYG9/81sNInINhSaXs6r/hS80Ov3YBUzs+Tq8kYCgRXccRmqiShg+w
ZEh53xfJ69iIczUGB3N/Wkp+l4jGJyfnR1HLh3s0j1niQ54p8P9DWRZC2vxjsSmu
XA1fJujJ4cXetSAxLAaksO4HSQUYM7gXg2ZAs1OVESbPuqWn5iiAdtwRiJCnstWN
qqeFBtHSw7vWVOBo9Nt8t5DC/rzzvbroBnIOy8yPYEjD2pIfQ5ksWs/9bJyrGH1c
KhuNOKNP2pQw6hejHC7HqaUPHoDhqupLttlG54x1d8q9HCSaW7vOMneeqVrnCef+
xt2mOJDf8u9dM0odJCcTQ76fR/h59A6r/zrLO7nPaUN/PI8OCfx7pNqhdJPNEVrV
EQbUxF4NDSsg/iLH7VSgGMUkR/Xxz6Lh9aouq7xQ6+O92sICHo1nvtpSo6VcKSTC
6MqbaAxWAIJ5jAVvyH2KvSb3hOo66oRBErI6Qm7Iq/JXcyfwqgfgLQ7aZV/C6Z1T
G4PowKQxdCxcsDoreoSp/JOla9/mFLff2MdAc+g6Py8lUmafm+aNKKM9o61y8lzF
ZhqOdzUge9Hfi10eO9U/6h4vR7KjQ/ec6XvTUFP9wPXcLL7UklKMpDHrNflcguZl
GQ5kFfwXE4pEV23FpkY85yKvE63M1JyXlOnpPj1hcX23oL99+veSguV4FvjtXG/v
69Q5kcSADQ8i9RHN+8WcVVo7Ae9hOF/VftgPeRB+WIXPbHLjW9799WxixBW2pyh4
gq5rsoGkh7uIiY82+Sztvw0XvlrbtFA8jLazUSACAgWWbGpg4SusaVvTb1xKHNlt
tEPbtf+41V7a5ypKDAvLudPoT/Ye3QdfkeSn/zM153HRdpgkKYpfFfWzG9g40CiM
8Zg83jumpuG9vlnnAYMCxvq6jx/xCONyx+OWtlizrXLhdrMSsPukt81QPrtdx09E
bMaBxb68sqeCEaPXMlijSqUh0cgUJm4WpWNpMF0xNqd7hjvSWC9qrZYj1m6VMFRL
JscTuB8USA3KhefDBbh9H5Km8i0+xi3bh83q4FXFKviRaRgPJ/Tr/6Pot7vCAK6z
NGl9vjZtSrzOGCAOHnBlY+0RIfjawvySLeLyScicRiHpShD3S2ExnVWZV5uwXf9m
qqpS7KX2nIawsXk4zbcvwv1EjE93dFGt4vKzMCw/oc3tU+tpYepVTinNgsFOtR6o
VmI+cc0YV2ex5naW1JIhQzqvKRpI78kc1KuM6dclLoT4ysORLdM/MvatO+nQUagK
ql+Exqc0civOa6mgHWDVzoFQR0OJpnDomipyWPtl9IzlMt4cjFXqFczJXLDjKWl7
HBRRekkRPFNN7zSi+xBQx2q7SQYm2iokWEIGAPghU+14//b6pYOfYUWzT0cUh5ba
plKGNZfk3OLkBEoXD0tVUugB4Le5MKvnF7aFlgy6I5dYU5To/8EThY6X5zj1awDT
yaPTosuFbGwYpQFGVbmKtdZTM/lfNMIl9VpCefKZShRhhhkzyu+VIldbCV4vGcfh
vfvc/C2fYnj5g9FXj9rJMXWT4ZJxBiCanTuHjlCAos9AyaL1Ewz3XPUUerYtDuJr
mIs4yQX78ZQ1Nlx5FXImA9bu0J6Q4lXIBnqzviEsG30zLopXXDnPXB6Zycvg0Aii
lt9I5O6wsPg6fQNP6TdnP+7y4zdt6yYVD3jNCKwtWJs/PPAsBDFsgclICjg75y1D
8ucje93JRnERNZ0MbQ6xgy/0iB0oaKhAnQwI4MmNwjtBqs0fGR/+cVT/B5l6meBT
v8jMDJKb7sXTLofCryCYvJamuwxFWrtwH+Mrj56lI1/kmiLzVDIVl3fSFG/dwxkv
hMkAHRAcOlPQ+T5/l48a1asw5K/YCloT0HnSDJXf+Dlvw1TAZp7VcMM44hGt43Qt
YmQmi9P/12gYan8uGeURqN1UBdKPXXkAaFjshsIt/XDAso/heZsJNwDiHyhEr2ki
PXUO2w+G2V6txcrXAiaUVdI9ybxURuheqr90GJcekHzpB2k1yLp2LE8R6tOiBK/l
N/tfTs7FlzEnglZ2Du4ozDGck0xcOrj4cjjzbwW5WTJaOYiABgW4COjac3waW3JF
G+5m8GtoPra4q5NRq6sAcZC7wrCcp3AAzQLMY0zxZ69Y1uuG7JPPTyv0rKYl0MAw
XNkMXAbQC3x4F4DxtYrEndUmO/4zwRQRZHSNpqNeyZ4P38LIk98D693bPjJ80ciW
pd0MygP9A2nWYHp3YKkZ1eQ8f2FsdTi/R/w7kpR/ZEAReSc77UE5GeSzZT4+adf0
oqRfJZU2YihW8zdHurjoIufQ0Kt6C0Q/1HDYFs6KahIaajNdZT2BprbI0aD3s///
I071BcbxMo9psx72XoIQo2rHTqM0Mjv+LHfkQpBo2/XsPTu4sJnu4qS/O/+g1ToH
8nHogJxLs49fWrPibovSGC6FJByCGkoET+sKCSssct5HVhehoJy74hn7EQ6of+LB
nF65Lrligjeh7Md8pNagMlc4FPjNmscBdVbSpCQWHRfjNdOH1MjI2amdHHppyKca
Qa7LS7o9ofpuz/VJUiRqd14w7C+6qxp+BzMXr12iPxQGPs78DEwPs8F309s4swRN
KJTDqFE5jIfhrzK486FEUPuyOmw5VW7wIrH56nAvKm06EzJl3CWDxYLOITSssGNk
GJxKrcChVXkERW/mkdwDiKwbkrFfvVpshnOnD/koRQE2B8BW4B6CBCHIj6KDYiJm
DI++f9inlZ6KcQb+Jm1D4KbuaAl49y3G3xC5635/51bDKCMNripAZAv35NUXHdt+
rdYK0AxvAp5XHyi2FXrr+YIgRKe4wJcO75nFiPM+ZJpN1jPAkGnUm5S52EK8p1e2
Kk/Kw/oip02CxJU3oPxhNzbVgndhQPM1CPtKJ7ERC0ZDx6qLnOx3NvwFi6pnB6ec
crX5g0CJboPI+YZzKuZPyE87ngYDoqse85BThzVrOED81uP9mvO8ZHAV/ys/BSSC
RQfQ/CyHcurNYElknozb7XnX31LPR6UEm128PsslKOhnXYaGFcKEsFKEVOJSKYa4
Lpv/ybbGMZUvDGaxAG/ss8ECaB+wic014cmt4G7xGhBsner7RmSdtWt6AG0AIgyx
L2EWg+UqUAAdcRaDzJQCjiBsLxgwENG/i2wRMNx82pg1+xNOZ+yZbfNEqGbrUsxd
VkJvRFRlbfE7mTRlFOnSuxHYiHaVNjzYLkclJjV4glXW9oM11OPeNiXSPvEp5Fsp
duh6JoOOhYaGbvPFhycQoNXmAgxCHfMAGT7j1nwJ+shY6S/OSGDjRp9EUOGep3xi
WmuWCF0Vpb0M6Wj+4b39nA30BvjGdSEPq5ksyNDs7iPpI08ehRfQmlOeQQAeQO0Q
/JzGX4E7+KtL3DzmG16quRHEIOesWbCkdtJua4gzZiOI0f3OGqwr8gqPh6CDM4/v
1xr8fqtIZguDOzhBZavTS3xRzzWa546TVv8cTyOiZtDIhWsnlKGErpDN8WFHT7Ca
CpHlh8PjWDREWN4Nr5uRqudlAPbOw2VRqdVX9fZj+aHNOT2TtokZl3lNABgSizRb
8LvgwWUXVfsEBEAvyGmYIhG0cqoH9pIf6DKTnJPDm+YIHT423UDMb6Au7fYg3cLi
rtQ5a/TYS6Qmcb2iBY2iLFoXfVwmIKbuhCSfaF9cV4YPK59cXgTkGU32AglPkogh
zLxievbejXJmC6hT/vCqhlVLnNj5bkyImDY7eKAIVb1PYmGjCsO2dxgTev7eBDZl
7tWrAqe90vP1Z4hggwGi3Z4VO8mqJFw5pDTtfX5n8XG5mVFWCBaIrHs8l5Cpbdg8
BIKfIckwgmhnTFk28xIu4u2y6QH/K7+M+RtZD6egQLolS9CqhvHiLN4FOY81JJAF
luzrWJwyYzKyB5yhTZGlI85EMq7NaAXmCU5MQUqcBMM7TCwT40rQib5kmn4INYLe
Pgys1Ar1CVeOtnawgd7erGxJ8yKmkgYAViWOeLX1Ba3IC4IF+wKHMQ18YPP/QkQK
aJCEaCSEN33e1OUBai5fscBS1omTSrmNoBm1j/Ir7zaxhwvzLNASrhGepSspja3g
BSsPrY2xshbWtYlmc93SkGQajv9UuHiXIBW8PZL1mXgDZWFVYZYflCZgAV7NageE
/1Hdk/ou00YJsSyec9sNa3wUh5TsmXNM3hOtPS4f+ruh6+RP/kqL1Gx2TT/o3KO+
0ruz05YUEEkVnps6mY2VjgCuNlN9RLLV6FAPdU7Q8ra4pPGm4dZ9N9j3ETL0lKqC
s/QQrOuF4dYXdRtmVHRgjzUlkBJuU9H4NKI6XVq5htFT+IUO+PRvg3p1VHO1fiBc
ARyjLD82l8eS4AJ4mCJ61x25o1wlQXQystFaC2C93tb7Fd2eDF8FjUrk+QL1nD67
d791rZyZ/U0qaynsybFoi281NxrqKV6/QyhUv45vOWIl3UvF6HZlPMOUhdz/u6ls
J2AmlOK8WHQxxmuMMgwyOMsDkHUwRxsv//sV1jSigvnEXr3vZYkqk0Kqbc9tJFV+
9husnq840rIaY3d1CyjEUzGMHYfbez4tKhYCuP5+8xoHyHmXda4Ge633RdDGyEzz
EpyT4R7Y/cYF/+B6pGnI7t3GmES/XNR07PBAicFNgZ2hx0EjpeSa1Ju3mG/Swljb
yCQRnacufbwbXe62y2FRc9Hb3pqIsjipkKQexQjthzBrUH0E00ISrxx5mr6nwaYi
u3002mRHE1W61uCO1NP6hivn9etXNT4fWQOyFJzS02lCSQ63OLPf1b0Y/K5mXXKI
ZVvY1M6sWSpvWLGTbUg4c4HE4htH3NjSR6NmXkiJLCuA5IdAKuMqmntF/DvtoZoV
hyo0Nx5APKYfkXx7tAbpI+Qqou1sdGfNwQPiGE4lfiT7LNhycyqTWnx6cZdH1Hry
s+FxE9oZHF4vMT2ABZNdNNWCJqNoY4elOLYcu2RmCOcODxGHJB67TahwJ0VLcvAb
x+BZfV8EJW9n19e4hkxeUhv81oGfVTVQQXAP1EKHUlTUZbOy/fK4wTliadJigJNj
qG3gYsAWWBNtjZgcS6jAFnS0t8giLRrJa8OoDhh5Y1HtyTYe/VALwofYUR0zGP69
FV1Q9GtycMm4R0JydBiM7jASpfFunuFIzDZlK/pYUIuA+zDMuKbvYbJdskOmQnuG
pAlwiN2dBTWbjrQOaHG3Z+ghFYM7qXjT9Nz4UuaSw73SJEhkFzQmKbUeYJdSTSSx
SSUykkQ5o7l3X/QA2KFD1DkBvIH21GlVhSKdqR/K/mjFLuEIuCVnLd9aw2AS800N
2oYkhlgy3kaSuG+nbWv980YyhNxfz4Q0mgEIQ7O08VxH2fwP0dkEb3UchfyMLeUr
7G4b71eXWDC5OSH0Fo2A0W6DNpBFTPJQcp801MI0cu5uPhgn5DjC9d16Yt2dV6W0
IX4EUaKxnWUzTsZcrw0bK3jhIMSmdkbjpD66yrqgAUS+HmWu6XAkJ3tSPHxXTeWW
F6YS6r9w+olDSXI6y5ZjU2GBD7NBpQ69BhPuRwVrJfW4UnKYBf6Ccha63mHBAD2P
lpKEd6Kt1BlB7FSmytxqLBelkfyXp1fiY4U4vPTwC2pAaVzdc5O61rh+6BWk8UK7
tYq0yq6wuZxeSumHPv0a1gvAbq7L0C+C7yeb/MbKer+UAYh48XBIesNxBPgCqs97
zAmYlIPuKMy2m44w/+b1teeHQRgnmltwv+B+RDMLmPI5RZ0l93HMDW754vQvvnSA
EHeCfo4KA37NqyJMvVMHtcJ9Qq3KtG1tMJZKi3eWlITn2I/NYzs1etyG89nCM50k
ReOZrYhpl0lgyahEezStVASRak+JUvRhK34yXPL2VofWMpPErQS09J6cBnl894cl
Ss5VQqm2jvPuZA6f4xXN+ZkQzEXU/IEEdMlB/J1rRck4lSJzKIhbjIgtQGHnjjFO
uWBiXs4x+XAyZ5qH3eGDjkedOrclZVlT7yVuCABpZdVVyfv/F+4hBG3uQ2htL4aD
3hWHeXM1jID4tJe5DMO8slsLTEZC6e8reCfri3Y+EJyKNILCLMlbd2wEwvHvF3DE
67bjsEmQd+/C9fuPoB+bbAAuF4GDVxjxeBuXH+COE2NKWrz3+YH8oe9n1pKVnoka
irNmQdFglFBt314ZuZpJO87C3yqTPBc69tXIBGJRpjBr2KZb9tqQqupD4vL4dMQh
q58eOuUxeyt8Pglv1Jac+kRbMWgwfGMebJ+upatqzbutC65OvycBfuPspPQ9fZML
bycMhi+C6y51aAk4AzxZHpWfINry/FjEG2pjP74lhhF6gM5LIEPFWHN3FK0qbuFZ
hlJwcGzCnurhM0HpYhDmdP3lTMwcBQ/eXpj21PQRmD0GjLqIuS81ALDX4x7NZ890
75Ah/9nk6jHhK5EwAqipFRrrX18JQOX9l5KGcljjSH7S/6bvo3nNg3U5Y4CZ5wlg
BIV6/NB0MaVUfNFZH695CV436u9pS/rNRjW+MEhjxXexAAT/U0qdbnn/ubiZvMV7
lSawxfroFUCe9ZeTIOStA85Wqf0JtjZrwo+be0jXgNVkbn7faRXLBOPucDPGerU0
q5iiE+MDIO0rAL8w7xe199UzmCwRKNoByUVs0JQS7cTPJGmALZ4AJ5LX3ZZZMm8Y
s5GyNa4XzYqOqHUii9T8j5ucmdrY9L1Hkzovt499QJtxSFTFfV+4Q14emXNNhFzf
maw07QpZK8tR97S1f/JWGcWvchSPaH2TIKu7dlHehXMaijX3Arx8kmJSBAr790z8
6ZJ0ePKAWiPVyC63PZq1e1FBIDHkf1Qx0YHz9/gsMuiJ4pyFYsVFXNsxQgfFy+s5
xAPUcmoFpwQnQPcv4qVoTVGTFz36dYFt4rE3+KU7zL93V8BKtEN68B+1KcHC8kjR
xuQQLwHpHtF2E+d50NqOLeFQoRlb4+3tgIMPZ0aIi3Vggx697kP0z1xHt3sevxd6
kDlEbJf0++z4EeiJMKKYVHh5TFp0HL2dfMcwSfsUKpblRzOlQl+q3jAnjnCR6KFV
6se8BtT6GhviP/tyu0Oe/mWdEJT6g61z9+qkU8minHOfZ/+uEsWdJjCWdQmwaeCq
/vZMwzbue4oX7KG7K3Nvc7WRul+tIl9LwYFJTHef04qzjvi4OPC14JcApMf8qWOj
XBxoCBbnyAlAmysEYCJgsP9j2YdILjCBNJlp4Wd9+L9Qs1xrxY9g+XzPly2W/Y2y
23C1PbijGw7k4vRO1CfYl+MmIq/I9UYVeFmGv1tBG6zp90Nv/IVsG2u5vSIf40e4
0ZegqrjDNX0tRMl2WNk6ikyIJ/Vm2m6gyJVW63usAjfmzR7cMIPLm6rp+fRMCHhX
h9qKZbxEHxnILxKyfKQvhpwy2YmVGqH4TVDq3qf4F+EQrk0WWbTtBzSdxecdL8V6
6AuO3Bia8XPo2q1mDv6vruGTC0r8Uk1mxW1u1t4Vrf7vpyhyEEetpZ1esU7F1ClA
aGyGhq0tLFOyK7U0S2Kt/E8oAWmjSo74ADEeKY3LW1Nhu1TJlC9aFoSicmR3uQKE
IrvJQXZ1UAu/fp7ejRppDKhbDGhoUa1g0D/aARXMgn6nEw9BReaJwgoh+C6NkkYt
7ZuvhnYEeduL0546XFMoyONIadMC72t8aKOTSP/0IYc3j4WoyUKoGYY18vq3fOo0
037jUp2GmV3qHLcIBfzd10V031beO0IIenI/LAdIYlAPL+3upKnQTdWZ5xt5fjQA
c2br2+2s3va9t4v8imrUurVBnUldpQYfYMYAkZCyj5qd6AVr7jus666h5+RRWDsr
hnUxrM6GXUAG2qJJvtgownJ70aTlMYdJI+giro5d6983P4xCVno/gy6x+yMF9n0j
PO1/3PxbW8T4CzvCvKshE30/kZAXOSRMSmvFwaJqaZ280qVofcUzi3mTd6L0KdXo
V/OBHD7hlbbtjNJqUv7PJfqW4tvuM/qeYiVppoY7F1MMp4wHSc8EPGHzOSQ4M7fc
Yx4HI2OeYq6dmq9vM1NlQneO3xKaynEM/OVMyJbMiS/6hGbDICag/in0uF8h5r/a
QW32rweK/bHliSnZGZoL4u1L4NplbEW4ID0K7Rld2XtqlmauXzNBml0KzdPU7WBl
hxbLs/H1fBHkc/oCybdvXy9t3cFWTnMY9Yf5aAOuWR9+F4SHzEVMvkXM6WyR743/
GEitGjQikKdSTXGDhVGkwakOMVDtUgjnfYojAQinuRn19ZtTZ/ARLhx1C5EYIQew
L7H3f7dItUQ+bjD5uEIIUUev6HRw7EjEhPFJGrevHehhs1rp1qjf8cf/gNIMSMaj
fCXS7OR1268+pOUPXQWyiQrapSc86oGIq8fzEg9EbYOXjZzW+c6WR7Eb5xegocbI
2avDoYccTVkqpLnO1IkhC8b1MIJEX4SZakX5KHdNMalEFkWhLPQraIqr5mhX0w6c
RoCdudcvGFUrPjhsZhN+NRoGIc1LYlgh5Lyrp+3UFFELCI6lnRT5uziTtzJsd+02
JDU2A88Ijrt+DrU/F9nK6PrHwIJnaH39aMa9dVWWnU98I7K28bSnCtFjuq7uQh42
/dnq0XYuYGjZ2zW/cCsbHwXEKhXSOIw4QalDGfF2hozDAWqz8rR6n20tsFKggodo
x5XrvvaY7PwPBjOfkjlWAsA8chGLcbTEqOulOIw2JMI9N0ExGySCZobG3n9I84Z1
shzy3hzwogJNM79zGnobCvBP2HtxX92ZUmoGwPf13sTsvohyztxRT53XDU7lNo2s
07rnSN0j8MxLFudev3alPjgoJn9sUQtIz2/g+Ro4QWJo93vc1ILcaELHC+yls2aL
0gwmm/lpB4225UXBEyZRbO8g3euATdGJRZWxNUIgILg2bg8ouF9t0S2XR5UVmoi6
rdLP9Up2CBR5O5+PBp01TWrlyu/nL1oAqlYgAtzGDx+EQOMlDb/eBV1fwRRuSPJH
nfuuvRKkOkGAY4huc3qZzcb5wP1cWMdntCyrgH7IuxtQ/6wxf4eJzH63hzndipFG
l7hUmzmIIM54IuwD504c9EpNwMPeJFWiaPBsZz9w5yEWsrqkT88YS0/d4Di/8Ji7
S/4poh9vuJ4jcJiUzj4dmUT2GpAah4JWM3r4OCUiQYa0JZh0MtgVbAT4qejfIQdW
yNrKV4xRWYd7T/NCUf7+p19P8hM5lLQMntNgJoHcQc4IFuFx4OT0UBG66EvDR+bX
qmKCwtTmxapfv1yRpPWu+b44Jx3/ogcM9iYVnydkZyveCKUegTQPjN8po+A5ufs7
nJm3iA36cWps5nnyDvVAV3qea7Wlw6yk/NdvbwojPLC8M/h90Jd2NkP3hLOvtasN
ebugRpoWprCLBItPFdVgg3kv0/Z8OGGcLdDRxBo9RncMVu6EDMlyQp0a0T2moNlc
GKjDyCqrrwL/gBhfi1bo23BWcNYv7fyYooFI3GK296cvb/ZFsQT4DNXlGytggTLk
c8/ySEsaFJyrp+JB/Wcu1QLkjZYpgDavPe/GyRRpKU7g0kC+4vyr6aT9PUtF9mRj
GxuAsZKXCc4kFBv3jIPATU9upQeFhnlfx6pisvGAiEb50bP4mwZU68aaGIKcO6U7
RvF9lxg0fLg3/v0owYdf3A53ne/eqBU/fR/BoHj5orI0OUKgDWkOjNMm/3TtKP7X
kM2no4IzXjDvi+mOt5RmNXMzfr/MlUs8NLLOYomb0iOgwR5y3S1WBcagSgXwDgf3
GstgsQlLT5CF3h92bfVDLV6S5cL77s5WDO50GwiOuyqRw8M4mtz6Xn1PekEGMSHZ
Z9WwP6Kr9tA8Tnns8omGKNY9aj+uzphsVfxbMT0aUjnHJUrzCG1xtuQULPb9lvN+
ujNGDENuTnVmdCE+CEhd1ljTJgdtYlweAFVF89aWP5Ho2okyvp1FiD2b01wqtVyz
AJhFHbfKFqi1SzMUWl2WOd7aooGrSpngnx65YyzJ2uyNIMMoJ11ys2CuO6W7hU2z
rsh1GoaZw8bJnmPaPzOjjkgHdORObmXbCE3GFnzKl/7pzOkYibAiprP8800bD8Nc
kkKObGMAGDUKOywlOP1AxkJ9Ah69Rxrn+ealq3gKXO3lPmtj23BCAK1frdqd6gqh
lBGx5ISvI3oC6EWOa3chjSM0IH+Z6ZRZRtSpMPLcAfD4RUicL112S9Jsdjbc/PyZ
+If16oTHXJQ7ukXdzr75B9JdMCPIj7CTu2KBza6ElEpQF1trJlV00lL4QW3ZLiTp
jP6SVwIdF5LLCEnnCWVvP+W+U+2cw2LFyHlpEA3i/eqkhagMqRnjlsUkku+xef2B
GvdG9NcGuRAV/xIWhurqWlU+cJTbkVJgCxSK0aFNeq2pHEpzu4MqJpDyxPk16ode
cQVEFrQt+9PNB0L59sgUOfwOXChG8xc2wGunPGnGnMisioe5V0IEuHoGYXKew68R
NkpNcxwgR2LBBuPU08QSlcnK12oTV+UMi8+mW5RHLv/l4WXQhozXzh9M5eRC/Ubr
7pD88ewyV4I9/CDvJVTtLMoTIHuwCjUA61oElrrJcFQPvT1XhNtkCNPrUekHc6Q6
qAtH4BFrGHilYOjly3BzBAGY0EQ2o8NvhcN6XULoxg+rq90Crt4gMRelNiaf/yrV
Ecj3w9i8utQzADSyqiL8Hg7hcRiYSxEQ+5n7jRfcNfD2BRndcAwWKvrb506nz23b
9WY4Xp4Ot6pfnKkZ8Qto+Kw2e3+sjkhORyT8jRVpBPr6BotBELYmT9IysPQAuNoJ
mmxRb9GD12mrBgp585YFctep751BYvYFMUMBs1rtEDmSf2JrHKvAu6tYD3st4S4i
ttG9SloltTJyPyARnMTxlZKfrT6diF8qrZp7ts89xUiisN00GVJeLkkbrcsV1zPW
X989U4aW/XByX0CHXSWYbO1PiTTEx0ZeMbK1fhKRyhIjR1k75Z9K+edotkXxZp8h
G7Zc7VYHd/Tpe7MA6o0pkb0yuFRBxbhU9d6e1CYdnYQBrVGfQUYwTFRiquXTmUUB
Rpw+Y/ujUHcZtvXLdzdtV/8TGWBbZ8SmpY0LEaHJQqet6zkfsrHaJ9Ism8z4pbLw
2xUl7A7OQld3KWkOV7+thMEnWwWoqMmXGhL9xRGUo01pDrL7E3H1OV0ZIzEqWg4Z
XPQfK9cG6XGE3JyimF3tgjyGQB77Ir/q2rfU9nQgPbpHvffuv7Wfkhx4fF9AW74n
GXaxEPQAU7RD4EPfkRM8DokvrEHNo7EsAuKts5jYfnKUxKSgLZTosymHcTMUF0MO
7NCk2wvseaUttLhXfQh9XKWsU1CcDAhoPEZY8TYUthA9FWYnW3S37XE5/9xrb1Dg
HOpGuCydIpBJMp0YI6od3WR7E5oxwB8lI5Jg9K0qCcSi4n+YanQyIBJU8nEOw33Z
TmiOMuYra6IY9zYOSgzdVZVi7ilcj7Ud6F5hm7d16SVt0v/+Nuh/tABl6TGuN2c0
BD+uJTfGPVTZyKlte9SjWBcjGNXIxn4NyR+1GH58SZvK1Ym4Kkdyl2rymqaqTwKu
f6pWqBKMjrcr/JjlEdDeiNLdZMS3FA6+ZI6K//J97InBi1TVc+v3iUEY5HqDvMIK
L495KcQPUoivmEeJRe14x3TMsVQMsPfVkZf7HoxZMYb5AGT03hEqOMSukyERlfpl
YDgYMVIezhvMA1u7iLt3oxeOvnHcPGWGk+8rB+xP+Ncv8s9KTU65vUHDnH5cMAWT
u4RGtgn2YmgKIiw189A2zxDEN3BuMbON6fARRHJMUF6eMbsIYfhh/swpdC9E0hNp
AehJRLcskgsK2K2FA2A4i6D+PMdGf3Yu0uRbN1vw2mTdKjlvNHUgyjpJh9eGHzdH
G1QWlWBrpTEkwQCGj786V9RsyguVMqYtBAGpwbCUND/40d8kI01Y/+ZIfE/uXvOg
UJb72V9brBmNAc9cmhbNTaG8B8LUAjOg/p89xGNR6S/9vIWDd4m/IfyLVccnsPYH
d/u9lBVDziQKNV7eOzFjEhDG9rsocmu3d+CYOhOyxAU77EQjKPRH4IS502BUJaWx
oDsmZZBOG8JUcr1bodnRXdWX7zwJql99gPYvOzWvuIdALDYb2EhvZ1uK9NKowRf1
gjS4VRR/Ot58PgLweAQjB/Xl0Ej4gYhbiUUjL7MqSvotOQLFWKxSb0+htWTEL/Z/
j4CPDoBvGph4a7ydRyshxs4NHg7IKlEIDX7LicWLZ+Z+vnYLEFPX5/o/It5ORMuF
XU2peXFknGXwUcqc9BNC3EJsZx9MCxQv4+t4LWyLkj6MsOuTQn88q5NsdnaguUjs
K5tTnux1vMG3+ymrMjjqHZuTyzx/rZ+7ExYplVYJmOMBm1bFVFxpWBPuRNK5Ljry
E4bjYhk23E5wfPYUmAqF6U3KKooLxSQTPOnQDHIVT35N2DglWtsm3devpid1w5I9
loTOUa9c8VtuEegsCh/GA0uO6/Gf6H2PdQj8HHJYXt1AEvRZjXUeHPDz5jGWjfD1
tb4pX/IjJzTw0+hmW3pzA9psJ2lnG7T73VbULTqD3PxT5Cw4F6gjulSt4XxW5VMS
2c2UlxdfgJc0U8e/AJlQ+qxE/yaNfWDV7XzO3zVcQiTG3BRYlSgzbzkmJN1gfBFi
RYVB9WVPCvZ8xty1mfAtDHrCRbXvyw/zpwpt9DDVWiJ6bJNk9SX0F/CYrhAhWlxG
tTsfi+9QBt24Igabi1hnSp04CXnwEtnLSchLq3PGrz7ErSr5Q8hqmMUzhs3kkkhQ
YtXnjQ3A/9cpvCfs1PN871ICqTZP+9smnPYw5RaVQsrpuahBZ0rQB5l+iWFz643c
lETppzKveBkrnX5wRan71L3IGtXkeBHJbSIQFCShfv2OCh1XFFmlbDp8IFnPvyUI
i/ckI4oyvO8gMqHH9lSz5jAdarTi4PUY4GEK0qZBIWxWiciUsa6xCej8aasUwmuV
pgEVU5NxObqv4cHWt9YJ/0qbpfzZY9VCY2kGMCIKLaMPwliHOrFNnxofpE6kFIkb
yfw1oiVWsUTmlRyW00VTow2SBHJMKCrVkxjS/7P59Ih4GEfcGLUHQaFnLVgNpAuG
MQavnS/UDMWvWjFXi22R6Wp6m01FkplOqPlIIYCBtwD+NSBc2dPPKAdHf/RoNJnm
ZmME4ipXhgTCVMjJiaIfCrgw5XipZmf5ADj+VX5EwS69htQpqYHUN5fNbWVDTE8R
u+fnyiB0hlrzrpQEQByMiiiUxbAe2ofvzXZOeYodL5yJclxC3iXMzJwIQDxMZyRv
KJDsYea/9xwh9MeC3ojOUepFUB6rYk8g/8Wd95wS0WaS6trhUirNO07btd3BhVTH
VU8OhqQ4r+lpEmwf1ITHY9MK4aCI0g6CBUzvGIMDjQRhc9R40RrBTVBCtBN3XGYb
z6xMjdR02A4leM+kwu6WKOidNyiAc4Pwi8/eqaxizJigKKEILO4Hcd3Glog2cYur
llgpVSr8XiGfvYuz54erwhcXTtyk3swh+G90St+5eeJkgIdpZL+VqWjKzSSySF6x
CwYGJ5AcIvEabzPk4Wf+DPwIP33rhf+Vi7kR+vy0NMCSBcHfwvlmdt9lAQt57Yn4
EKsOfBMObnD4tJQ5Gx+bTxVt0Z3P68s+5N1yHoJ+BPv5YoHRST7A/ZiW5WNCnpR+
U7tlzlvhn22+mBkKVjymnzTj2gsBAENRlCjyCAm0t8k0QcaCthTf5B0/gSIOnsxF
XXNUAjcMbM/E32xahqT/ZO3VUdRcO6ZgcaB+4u94sJtEpom+sv7IE58jf9ASxXYZ
1la7QDiNYQmjBkdpW3nQKhSMRrmQHOJ/ahoa/a6O5cYltiIaZ5neL4bMYhusWX1n
NwSQzuC2FYpUXRoA1bibu0XDG0SNtAqA/lq5i4XOolx2LxyI/V6N/UOTuiLitbr5
WmH+xa0KRjFoH8PMKLNdtq/O7Tz3fcZgG0qEuhDLZzVB3gbiVs8CoZmm5gH/xwsw
Jub7r/EYDKtnwKEgyk8fPL0c2aW0Bt0Hl6Lvq/ZrmB/ko8p9C0joYrtJ0QCBuKuZ
aABzHU78C9aFzQYIlBeXvoxip1T5frDEDNO9jCD/iY1Dnw9iqhd1dRshTwP5R9DC
UQ0D8+hKUJeetOPLPyUijw7AMBTTyraCUXVwm2Iv7nFBsMo05/cs2S+ppz+Pd9nC
VRtlK3zldTmPn+vAPrFzqCGuc+jtDwKwsnGICWOj6Ber5N4vQveww6PDAL908pSD
44OR3vIkbM2+fttkA1UXssOr5SAgA5VE9Ye2zyH5oZJ+8Caas4xX6tKsnd05cwR1
bF8e7gKpYSUnIlfkW3ksyhlRA1iu0UywLUR8snaRyZf7UMCd5KmfaGBSjYgUeYJ3
An4/L5mdMwr4BiB2vsCtSIYm4/8Aj74FOLE+2CQ5Ff/ooigD5asTu9QV6/H7Cc8p
iJ4BzXa/XuWXAEZuzhwCGuhbKYki/YhAg/ClRcIIr9Vx+LEdT1ci4c2o8RE9hy81
pE1PWpc6D4oPjD1C01id1yJsE1eDB57KpfzWsoRT7fnNTDmqvxuge5of5oO/cUOq
cJAiZTLP5BPsoLc6+OtoCBNg9HucrMnMV67kjbr/9lumQkeZiF4Z6LYtppFixJYj
O+wooO7SuS88mlQoHFIcZZIbQbQs0/HplHzhp+R4WXBaD3x1IrEZsumk6BhWRI3l
DZGppU7YU48OcU3z9kTmR32ESyaDJY0rnlAfLua6wDGl5EAq6JCflYoWvUxd6KZv
Rd4XuNtxla8Jpw3f919ahvDSqexxwjrZ3pnEXs4O6IuREsWXMVxFrCXjrkiZcNwr
h/YWCuMoknmLx0r2wzzd+UtT3Lc0uaHyYJObhN8gpRHoV3COdM7HhCBxM3qDTcOT
HOUlx08qHgHG2ZZ3qwmgh8u2d2JZgK+uY93zFiQImu3/98kunn1ph9HOkXkhMZA+
0oo9a3oh7ZO+7Q+yDOUyEEpInPAA4EPd5LMHvYMH6xA+4lryMdFQBkXY66f9mot7
xGxCeh1RV8EL9z1dAKzrO6N5BRnE04NBcQRvCOIDucW2z0JmIwjVCKDYXng3C/95
6gNxkTM1lhwtfPh27MaSVwQTGwfGshl3nCv5yCHDm/WtFcn55zH1kUMhR9qyfeAM
hLn6c3dr0vyssQII7LgOyq96kIH23enYnJLP21inxYCFk6VfG4zUrtFJXP88WD67
k7MIWD3mqtv8SdnkJAlbq/w7DdkduY02I1v4/BAYtB+aXfyc7dD62jJWJCtLcuKh
AfiSShZsvwt7zvIbF2cAKAOjS+25eXLILmrrLvLyUoPy53XbFod8FUBOXtNlJuu1
5N4/rVtYbZWW99bea7V6YhdyMx3TNd/B69xsJUI5fK6snt8FdfAr1YTZ3Cccln8j
SwqR/OPQ1KtSYlGSX2AVbCZmWPT+rL099beXy4fgEiop9Bm3NEpO19aM47ijhuy0
YwIbzVyZ0fIp2pf5aCTCHoiuuCY9sbS9P07Ux8ke2gug8F17LnPNptzbpL8yfDbL
2kyAm9QSGI9rsXUPOa7n2NNbp9LE4kU2KV5Z4C5d+cZlvyLVvVdWh63zPQNcbZHu
WrzRRs9uRNdpNFjwWB7dY+W61zp+pc6S4hi+C4FODgC3yJUDl09najQLQYAtJYP7
7i8AaouMYRXjJfuJvoRDWd3FsqUVLCCNMB8A7op2lD0grECNYbnSm1wX//6EwC9W
lED5pF68RF2lQ14HRENWCU7ud97CQvvTQS3Aus1LcGbWHjZwisapFr/8VXswmdnN
d5AcljEXOkGOwXFnQgr3hs0LYyeFkpv9dwnH4wViwKXBGIFAuyme4K0ZYu+0qXH9
4LXh/bV+qydvJ3TPhsBydSpjpZ04imWL5KMDMFYqhzFH6p2V1WXEcM/gB4Q1qYCq
bHB7Hd+5ycPAeD5p1qx8sQrDCSZOcg3CuD2+gPsPA5LU1oCGMqv4TCw8tiEui2uL
a1tPaT1uLT49/xeeP1xZY+qUBcZlJE4S24ZFmeVfI48bbXLXYIca0KYHQ4Prt2Q7
rmXivfT6rDGAJqGlwYXcOl+6ArFtU/DLk56JwO10aJ3c1qtoSkvB+9ZCJBfWaA1O
J/NBKmFdIdMkY75KvY7Zkb33lOtAx5SEM9nvQdJ9KmcRmoa3nWKq5xUBpj4pAqgt
YtTMdHaBUeP3tUp/1bRR/lC81ZEKSa5BqSBme+2b+osxaq9KmndAbdCkpJ3sd0CZ
IVcGPsFS7Smjig9o5E4+7aZufOPwKwx9rJMRaxCAX15gva/G8iMZTN1U/OrHCDzG
QcieeBXFntbgaeQ7Z00lBGsSntLKlIppttU4YhWdnARd3ainqx2BdbM4E96hn4P+
N/PUQE4yafXlbKUeLm5ERDRfbm7y+HbKphlRsSj9O+2rY9lOL9yKqLQ1/YCBam6V
cZEa70eGy86f2G8WI3rFJyAVu1eap0WiKDWRUU3XaB1FJTRBkAPVXwn5gr3H3uqk
zAVnINyH7XO57++nv+o1ftmvXeP4mdinw0dt0R2XgswBKhBDmzFmiz+YAgoUxslT
L/hZjgP8GieJdcp++/LmPY32jl5ROzyXhVECOebw8E/7VFN20uxxOGx/nXtXzAjX
3fR6SbCpHKNqkuRYn6M/a3ZMTmW4EPMR60uRAyPsY+V/urWcCNJmtFvgZNWGwBzf
fo0Ipe9eYWNXF5pDWaBnRbTDK15cT5J3tyKQ0M8TGu+7HsjagAejDOP1CgAeKWkT
z55XxG6thl+gKzEQLVKQp5utQ166xEWS2Y87xEcRaniIo1bAS+BY2fE93bl/RvWN
jTNnbVoOTP2TtdzkTtREeWbVmepHTLN/qb5wLeaFeznO3OlwSUtZjlvc6KATmJeW
uXuVX0k2RqcyXPZ9uCtZfQM8bdr5F9FnrP2u8AXr5TAHycHp3xWEUx1gG6zyJPOw
YRiH+onuuP+FjtdHPJ/t15+EKLD6au/afyEZRVEIJ+Ietg3hz0hXmJU9dRJ+/CAb
1NKr0wdKyhQi0WJVKgsdUwn/ukmUdlY/5YWAoOwdDlQOD/IcLYyrE+6JT+XU+fvh
Qqc4ZwsSM1d8OLyokINdwaNIAogkVcabytQg3U4JfLrkB29ssVkfW+x2qddTpkty
TV1IAniFk5IOVL20CbasQUQLWrdWfaYi/PD5HxGgNBtdzWZLIU84AEbz3NVcpSaJ
dj2bxg+jMe5dImvee5EjGtEF7TTfTxzB5upAxSMNx/CMlZd8598X8p15IVpSQ3kY
zF8tKEUz3msLO/ZcWbDpGJV7LfqBBNtD2uYFtT4kpuWuf0inp9pN8rNoyKIu7xR6
/WXIwsweZALZwoJubuOpSSWr9pw9oSFIZx/VjEK3qh4ECHx+yvMY05XJwJBRyx3z
9WdEo98N0TA99MMLDszre0R8dshDgPdPbLZmP6Lr6r00D+chJhP9zroSUg6gE1JB
H+zJjl3nc0efLe3HpOO0J1JGhqABdlfm3joXby3hnLjsFVNKxUeMTA9fzooCUJTC
uxwuZAcoG/ntda+qPVQFylFgsDgVCXmqC6yfsYkVfdOIm8MFs8tGjV5+WKD0fvP5
wVCPRqmT+Bo9uI+i9ZxYVQBnVpxZz1jMgwNy2yoktZU0YBqPoFvftrclrXwZ5pQI
CBabDBBBr9qb9+Bfoa7EXrrDieNipsoi884BRP3fp08Oldy5oqoHELHvdKHaFLAR
PzaleTI8ZBO08ZKt1eT4NU01An0U/7LP600AQWlJw0ToGgluVtCq+ZxqfNU0Ymop
Cw4tnl8F85i1jSGw/vjv6vvrN/++GUyqv93x7gosrGt34piXISlsQFbLbCCDnyiM
lLJRi2OhGq8I0Agko5XcCzOwMQ6AENMMYxb/MfXiI7sQAo4I73jpBoQSkmPt2Asl
8y87IIBFIrlc0KNhAiiTJYAlolgNB4f01uUnWZwnBxEXBIxnRzUixtQ1OcOnwvab
ErX3RICKPi6Xo6BUp0TAUEODULFswTay9w8a4mA8VjLw9zgCie5HwnHAv83TWWAS
T9fs6fHwqJDub4ZECyM3i9og80VjPqA0+Yf1FnyoPK0ShwpPmlG8MHK4Oe6at0RN
S4zIyyDAH58PiZtaYwQY/dlvQqlpOb0L3N4wgeuPIxWOui83ut7goCV9E+LLrX7f
SPWdmfOTAV+fHxuSK0hDi0OoOyvTx18Jb2K+mv5tUjyIvwI7pN0yETDauTFb8Qlh
Hu/M30ZIiaI9CInlvF6d9bYYgwCWMl58mnuArWGqRyvgm+wn+VenAtnRMv+AvSnQ
Vuy1EyKXzHM4Xp7I0UopCdTLnPpSPJDLjLb05vCUSIvOyeQbt67rnnLeledIHjJr
ichuhKsMMzyXr/0oolOX9W13tBvEEty1mTEEH6QRAVrBXrDZ/azDutjmNBlXySak
eBA12WYUK5uDSBtcQhnBVFajoeJ36rG5pyPrlMp8LhXfQ+a9rMOurvkq5wPGS0Hp
Drj/LrRFT0HXV52f3J+Wmz9y0B+8c4ie7ndjV8Le8wYeMWCAWMuvsXuhokyTXrdi
9KwWl7RTLiGw34Q/nNs34wMOdyxxuv/shT1EfDGIqevsbhhGGAEMB3AwE644QWJ8
SV91iE4YP/91TorrSt56J+INHQKxa7YuOYWcYubcRPZHNCVb+wUmhOhHJx/m8Iz6
Cma2XMvPg0atdi6UXjjLxaD2V9SOQebKP1WMOq3jo/BCa8pup08ctSJ/iEohcKEe
hQAzHfgFXdMdgOABTh1Suw5+x1EcqIFVz1KXbCPzFB58kRTHVzEn4ike0OjDEY/E
5TGFgp+468z/PHFkouQy7eMjJwC2Je8u2JCAMbFWFdRQMKDlNLRxhtKDT/KtypeW
sOzD1g9Y41TM5IXnFvn8P0lwVBpKEsR9+q+DgieWklYnUmdcND+KUDYLGqGS0B5h
8LBMD1pOU+p1xAju3I/laPwwJkY0rNNkYvbPB96PQrYlzFWj40oSNYgIzlBw8tva
22FSLDNEJhydqqzBn58xK4etJgALkvBmRPFmNSJSTaHVRencc24S7HC8LCIHv6FT
naz3NGqB5zyjbX6BgWj46rnucw8K0Bqz+2NVLUbbiNWbPTWQh3YcnN8VTZZD84Sy
VwCnBVMYTVdryOK+n4lsjzvjbwnJoT07kF1FfpsqLuY02ChCB3SxaAzfl3yPzOa4
e61Rsn3qrKqTGI0aupzIHtR4GyzctHr23kIdNnJ5Xi10UhqWfTKAVnAd2088p8AP
Ds7P4ysPesfJqwHVhurJNnjGd3jrjanSRDP6T8iLYmK95Clp7sR1CuKmcYC7Cy6f
rIKnuYHu3TkOOllkOcbYkBgt+xI7PdNXhR28iALLPPjQrTvtaktEsbu24M+N9pxm
wvHiMFsBeGnJQVwq/1gs6hYD5teJjwqtrZR4SP4tnizngk7+Q1zD8rHobppLHzTR
ybHN5WQ2vXcM/XKs35t9MXC4fgMfsvvCBFoRrURDT8xqibZN3cDXlHRqa/Fire6g
DGhV4rd2ZkNo2VOxFf2ruUV/6qclQpfCSHx0Lp1s4bw/2VcFPqHAP3nwl/0oVSGN
KkCk3b744L+Woi500ApiOlA/N4BSujoaCH1nxVcmNGyunlOKrV7OMOW0j1zMbBjD
GNuZJMXtYSNaOssMxOhje3kcaK7y4rgEYmU3hqzwCzPk3Q9tjtmc+/G0zyOA0AEZ
11rYLUZ5pAfGvyypuR4Lyvyi4h/OFMp1sv6dGGm4HwGHXCddwJJFOmM6RaXRhGfb
EQu8tvtqfe59uP1twfjotvPVthIM4dSXOuvSekWnrOtyq/F3KdX2O0gSCebeTgF0
gtCKC+UQiivFS8nJt3NFkkz+k5oWgdxYc9Fv10X/zrEe13MH3B2ckJFebmoHCsiA
QXjaCVb5f6UPDVbzsQYWZ0LMziXvPOW4gRRU282mRPIaz7gfAKSSKftTH6jELspP
ePw23KaoQGdjV9RjXSY+tm0F9bzsMMj6oFPiadjbcnHjGI2doRANnqARwg2KXq48
Ui/Qp1ZF1UuCJ81Nt6FHff1aPjlvUNHKptO38hMMNAUUBLQlRXKbBvKLM0e84+OO
25V1B8jaqTvT4gE9jgzoEmdNLKxTwQsRgKgh00Oi2QxEgIDfd6ZJPJFEVxDOMclf
G02Po1/7ozioVUliwrWwWenPScLhVg9wS4yxWXG/JY0yakso5pHsEMnRnx00aIV4
mjXoYVdsQjBGLrSchoQSmkZIbmc+tbDISq3BmTd2w/MGDCDPSooM7g4+Nk1ekCmD
th7jol5CdMQh9b3XGGF5PcegBejgJZB2m5elz43Z12E5j7fct9NlkIprhvbZN/6/
DSdvBVni3JMukr5q4YjdenzCplMgaYsKVVdh0f8rK+NRqYYqoRSmKxnGoz2mY/Ji
qQjzyWHQBqcKezqSYDu0GwWfhPm3NSm3lqdMN0EGhAhC83Z3JbF914F+xlniJhx7
IqU4Nw5LbSetjhmEZBPtQ8hs0LU7WpIgYgmB7mvKr6/1B+ZammNN1om9ZAptfRUq
CD6Iee9mt9UBsy0raoerNaHwoKZbIyfoN0ZkPouvz/SePS/PJ5RjWXQ0xNIP2VSD
55+RZQHeFlmkWQuYAJlG/FyYt4hhASGDHxT6OV5zEdw5DRZic1K67H4vDiednkrb
7dHRkzba4mH9m1WV8YNLGB0oYsehxSaDCPVp+5L444Af+iOjW1sruWeRAahngHtb
qDAG+i4/8kSl4S9pMKEg3F4y8M1lKNiAx2XF0WnXNep5EfRTb/tLEaCq/wsC1qHM
tzQvABWVai6UmK+qLBOJxahI0Vext0rNQM8OvXJ1EBU73iTedY0bSxw4Ib3TXmZh
NmQh+/8FuwpzfCQIfwj1smO0MUmM3ud1r7kEVZtih0vq1wxq8pP9jJ589vNxDbQ8
neEiXS9tJHO/xhOVOLRerEJjI2QL0NiwejmyygDZdtpME1b+vyXp1RU4BjofEexY
wAVEGvFOCU+pRVC+xKJRt4CV4Ve2LvUJJ4JTrjnT5QHDy+GZeMahfIWhw3sYjFX8
BRSvY+J/HwqUwFhQsIBVCOiLgZzL85K4p9CZ7Q9V578Rodk8TQAETc/C7cXYzF3b
oAsxjB/Iv7reAIb3pYy8IeLw0xpAws/HpW0VUDI46X7p7zyjCrm8Xh16X94BDzRi
i6LVjbnOfTV7UEAiw0ZB24GyKGNon7fGbSGlhzJ0s5QCqu56gmqOlgSxR3BBdXbR
SdplTH/8Ez5elaSxUMG720YxStkI5DDYt3c6rq3EGE9DC43ICepevKE1Y3j6tUs/
fmCVlI+FHvGgMSkLViK2AhpcixhoPSofyUtJx9Np34m4X/XVEUwoaK/IL5Rcco89
8mGvSnbfKPU7q36+zOMwW/UAANQfNwMN6YlSahHBKjWeVQXoPl8Uv8JXWwfA6cjn
3/9X77R47nXWdi5PuQWT+teTa7joBtmA38cOfYwPBZ7vyImKAOHVB36d1s/9jcPw
1Gzau8Z2ip7AogmX8cXAeee1+xjVxjRXHDSmIax8lYDdnmq8NDYvcnKq1VMDRJK9
sOcgbRFdT21brgbIxWVihfCpRKvYz+wTVzOiYMHSbmcCXbw919LjonirpWR8BClD
vK/WEmbFOvg2ZSM3wdouzBpuVhP3PP0QFNd3yNM7VtXsiJbukA2Z8T0t9uvAn86Y
T9ftSAXkPEumtAvg4wfa7zLkVFtr/Lyq9l1mUkIHbxMzuC2GRTyH3hGgH3wLtqkp
7LQ+jQOkDyQd8lg2RcO82caeAgOK2VdRw6Cp47erlPbTxrca92S1hYxbd5ogTXTV
uDr0wY8f53SfhsggBvYA+YE37Jywxq5VLYK+HKAsmxf9zMX7iDqB46vEMPvWMTcu
oCr6i/DJl/0XyI/M8NKx7qqXI+ZZnY0HO6BgbnpbUI/Fy5dvILR3os1xHw0sTmjp
N+Z9IoZj4C4tq4dFtLToPIIRT0rAea5L4cdOOOVmO5NSLku9rCo832urI8g4DiHu
jzKmORmDYZ1oUzgy3dL1HYnD7V7EHEN8wBsZd7hS4GfPc2W/5iWTFXuW1QHK0uHD
o1iChXKEMD9PWUq5AzEcL6FVUuf1BYxDCaQIVFEw79pc0hvGuATy5T9DXs1pCZsl
0h8KX5o4f9c2D0ZLIA2LQEdaJwfPEmjukhWJkvCMe3WRdaAau7isoxW4HepnVxl7
7EvFFtRx4uIO+JHlgjfzkfIfankdcn7hMmi7gT0rF7Alm3AAXClWqyF011GfBplj
BcnxXQIMuCYQABo2TJaGY/jRWX/ANULpnl2bcCJWOYiVRgBZeEVmHVvo7/yg0zsu
CSZEIOX7QYvHbebCT9I/aSiKBuwsPvJ9bMjE+l8VHIoH4OiFuud8Io4YyTE2n5qI
C+2gbVKLLlSQ1xyN/fY96Ts+OYj8CBN5y0meDLerhy9D4W6rx950Aa2rsGLt7gJ+
OCGY6YimO9UKO88m1C0hFVkfQipMte+COeziqvT5QbKmOooPrC9Ws89MVQK9+QrB
zKkhIZxKIE4igVvZWN0AzylXTlFco2/J0RlleOsEMghYNLurl56Lkv9/9GjOl7kR
CfR/fPSvJCmjz9ArtTVOpq5e2n7yOQGBJlmfWur7VHSyaldRctu6RdWYia2mIdjO
4qG/1UcVIKYim6n/kY2+nAGkd0/AXMooD2sPLAbyhlSCXFb2ro02Sm6HaV2IUG9+
ONej+mcnmp1wApJ4f/03oLiRweJsGbJ6VrDZMq9hPVtP2w2xi9MbzQ2Ue+vH4fZ+
n7d2kpHtcViKqQwdW8fy97he+FkuWO5PF2PUP9kpQvrlVf2M18MXSKomE02HyFfm
nipgPC7nztMbnMYl8QLQbhXABAS62Ape679SaG4ltawmjE0iX15064rJiZH5kTLB
EjjT3TCpflGftJD/Lh55NSCtgelU6G24FdBR1dSgfipkrMwsyVORMyy/Wr7qDfGE
9jdzOmovYfq5BGN7tBPjfldnATP3WJpWrkJ2PGUkscoKKrYYeA1Oj/PFXCfUH7jz
2jwotzZSK7d3deEJ9yXlFMNLi84Pdshjg56wdqofh9O03DjFL+tObp6wKaFbtY8T
XpLGGZ8JB6F7txt0ZFtjmbyPK/03HsIEh8RI8jkVdagHgWye685yREhqZqCY+iXC
hQGUFELFbyt9oPvClF2BKInyPlhrQ8uyWkeeQT1VY+L9e7OwbaMsW+1pwLE2rD5/
vkiIcY8VQWYxirK5xmsDNzE/fsXVssqipzlhAUjWgjer495Ib7bFXDcJsbCdejVS
QlYwzX8YJo4z1iyJ/t+Ojs2NBX3p/NDdFMcuT7knBkqf/tYmwXn+6O1z0loqwQPF
unGtWyA2QvSYR3H+zjJEdMYU2dnX8HXVyAxwO1f3Z+IFOwoGMl0ofsMxyVRUxxjd
LT+SnsF3P1diOLxHcPYWUdoJ38BouxtNmQz7NK4vS6g2ByRGKfaHDaQsmJlCnVtH
sbp5WPuiOD5aVgoHKoJGA72IfOPkL+vP48CsAHxzl6CgOFd7TX/Rk1agfcV4GAdF
z4y+TL//SOuGFhokRP8HSWiWcR5FE1V+xaGeGa6XjflND0CfeIqtfbhVXa7ADa3N
7hPblUgqWQDM0xmneLohdf/PB6kJNQ7BKhGEuKn21SUISTURc8aM3OQgZKVE4E9e
A0nqWXBdhPaZ+fVe5BQIvD11WFPHliIVtzr7TPsqbTFwdvgAzuWiYe9cudcqbS4K
ZM08t0b098zgaucCiN1w3tBUER9F8YZlU49dGX0Tso9oDQ1l8G69j4wi47R9id+T
XO4BcJdodyphLpwmGTvN7bOIfve3n7Hhz97BAA8Qug2tOebmQPZ5bPRo/kBnU9jO
KjJ8/TWodKwfr2MfwOMFfVxes/7d9ZsWUDVKBvCwHNCNcBQJvyUIp3rOMy4YC72j
Pnr6YoAk93ZhhULMnpmAd5uNbsSiPIai0HQEAX6w0cr6KrT7HCcfAl3u+QVk79he
JFOBIf4/vbwqRbnOLLAy+bMS+9DcG3b2qqe5kErp1fXXaae0MZXcHTwIZg49ZlpY
bAFRYV3XICJLHqDYHhv2Dcd8u7ZdUpIwQsEOSlaDQ7xfeODpiT+HxLWvCKVg9ump
GKsaQIWupbON6bp0yhBGvK3NAExHwJjYWd42AFnXF/v0lleRCDZqHHRTN+QG4GIm
CKe9LzGQTXCA8amYtLxhcTy3uSeuMedMHJDAjyHbRD+m3Wnlis5cdc2/wnegcOCB
Sn+lYnNmjIbgSblZZ3bddgOGXyPzBrXnY7/rju/tN+EioOIymnFh3lWUQEzmWfr9
qbZUBDozQ4e1wx4j6+M3tHsqJZrJyLeIGOw3yj2EveC6fyvlf0lsdB9q4iLYcwYw
VfCm85byMFiw/dk9gkHJdlBs/GGNNBPe7X/v7b6IJTT6cw2xTp7tT8xTtRNrGFms
RfaLxv47YiyHSUUGeuCKVMAv6qUM5gkScIfPx1S+kS4lYWvpSxuLAJ1xYfXFhu5q
pkvGfoQE7Ntr+AiAn2tT4NzMIzbDfvCWB5n0XS+U2ph7jflgnT46V/SrYrqInTLh
DqqFf2OipXnFWqpOS/hDKz+sn5PYWmYsQ3vLAgvkKv5DEKtGl6GWJ4WezXPRgq1O
1Nh/d94kCLjmpm+BYY7YbIBIfRgjnynivyk6JlSMKrZialYqiEiusL9cE7Jw4/lf
oynbJWstcSvzcT5tQuo8JCwsUjYJh+MsqSVzXysc4X9Ip45EvwYyyRYpkc6ZTVaE
EzUxyIGPLxpAVeASyX+bgVBKNG5PXLUL6SpYREeNWtgMtAGlNW51JSpdGZ8++MJv
3lBhMhmg1nN+GUJnI128aWbhWbpCmidM+AdnE9E2Q/UURRz+BEV6PkyM6iNltZMW
Y2XKgTpCXYHVbsu2s8ZzTjj79M8Jlw7Nk5RmbR1/2Ene08YMoDRE9HlN+mMBq6VA
vBb+CwkTcQSElSXXeA8N8meraRN5Ao/kRLgiZeZbrcNMzAUbaJ0/MsStKxAJ64zE
FkoD7ROZ1SBpsH/V95unnQJwhYoyRFMLJ/iTmroHHT2YdiU7kakB/kFtHfRnI/6Z
rY7OT47VpSzNUHZU34N6o+B8/szQItP+cdtqhkgiQvqx7CbPGozeTGwg7dL7mTPt
9tCEBGYOLST04WpmJVqbICFuLuG/8M43gFyiMb9Nmy4cqogyj72WMMULEODYmVEy
vfbohBdglXVJsL8DUl/SS8LaRplQ8W8rAykCpD3blpikezMJyUyV0km8iYHISz8J
8axyYfk8t4/7dLT1uZcX4SlYvcPiY+oeWB+QTmHXxDID/Ep4zn383MnZSR040+hm
g/50ytp/SS/0fHDKZXRYk6NzaArJoKzI1dwkvBNQXPAsBUuHdg8jDFWGyEsFfQXi
vdwA6qFm+d6F54RzjwAUOEYv2b1oKkOYPjCMIEeAHkm/7Uno8HX88vO4/rjLhy7r
G97uolNpTde7pi6gGhy2HdbqHGiENZ8Tpnk/UhFjS1hXQN7M66ls3cXc+yW7yQ7u
QqME+GGdDEg4BN+9TQhU6z/6Qv6OTcW9xXW0DgCSvEqbO7rByfL8fh1l9n3aQjjY
RO1RBTkgZMIFYbC07ZUnA1hP658uk7dQHxcUkHZDAmzRozWfy3D6pB2fNGsoai2z
IpT4e3VMrCtUxgwyufn9BVQSQvAVjCbERtT/LGNsZT74WLIqRnn31vlJGXx9EZX3
5gLJeJKJ5Pl7TuYjv4WIHDNcmioocLFfacNLxZLidKPD/+4BZDo+hM+UWzILxq3F
wSQlGYuoxtdWW/kpkjm5F3lVrxMIZVUxd+opq48Nra0mXb2weHdxEyqmajinU5sR
+FdhUFQnYTkrSmva9NW721ccc1n4+6UoH1MWBv9lU6H5otJIAA15s+vunQWPCT5J
Y7x9HdXB+U2w5X88OJWqmOOIrpMl/XbyI5M9Kl8IU31kERJqM8CohAh2LVZjRiBW
pv2ATTS2BWYBm5i6JkbE7O2wT46j3rYTx5Ui4+JqlBn1+RtxZ9/KFnUjkA6grxns
NTmCAng/GS4IJarwBMGANJJEh4YknoPS2qANWEz8WrK1+eTKcGLYlXWwWUfB8lz3
xdQIh0OwgG02Y7uIRIuMJwn/aXKtG0IWDixg4/AxdBpL22F6blg7h0ark+U0aoRw
mokpJsQNqlBJ8rLCETcpEUGvkuPRfzRs1mhHrKjdwfxSjPM/+lPP7GzbLYg0MNGm
koij5vyfDcJU8aCdamVTzvT7rw228UkwlZG2hIqtbhkMDMi1DGlYFxdIzpM+jhMo
EU8VApK44iW4+lpRDSNnYEccnFf2Cax56XyK/8xDuslDj/07xn7OfkvWpDB6cwHl
8h3Y6bQNYY0aeThNRIMw7XU7PrHAQ+lHRwdn9GoFGmhrOGDdxBjHVpwRQBO0aczj
yDkvV12P4WR6tA9qQiDpe7LNBdsJQAWND85MYx1lorGTLzm5mkOUIDFQVZpd9o1g
uqL+ec/qAIdoBkmM+vNhzO5NEajtK8QV3wIw1Og6j89UD5Xjs0UZMqYMQgUYpsNO
fPOWuU/E2yCXWOuPA1pzd4lzqnmqb6zmBQejNDkMfElPOgCsBAqnnDIAMHijvzYg
TfNBlnV4/xfEsj6JfWCFcGdFsseaq37i6EFp3ayTfWNZ6CYNpcoVDPScidgV5hvr
nST7adALmpsg4f+Gpu4+73+WMXevwhZatra9XMqBSpX4PbyoFE/0l67ePzhfeJRx
8E5zPhU7veiC8nYMsmiVinqzH0vSm3QCtq8FcQ6ulXGcuRWf6ZpfikQf4biv6bb7
3vUnixwHChiQIziK9TEPApLUJA4RnRqRWF1gosSNOhrKh89QluzGd8wbAi2AzmPF
bM2LlCWi2llLLkjWWAkwDA5qyioBZtZxmMs6ktoqIlTRt+0ASztSsILvLjcHTe8j
OPz6a+nOgTNwkavbpHTsoLpMxSARafKky0pD4cK+axNe4Q1+0oxuDz+Cj5axj9I5
v302G0rVvze4ByE/blJagQa/oprnkLAqhtlv5xG/6TurAcDOZxjTEgdgLYxI6wg8
9nWaJj4X4KjyJKuv3lPHzPt35i3PNmWmPBGyjMjZe0hBRGg2zaoJzPibb8dEeBYR
efLB+coAHGf3MBKIA4Mc87KefqK6uwo27SXra158UDI5In9JkKIMhcspn5c6QgNY
193+gp1KxC0HCvfih104bTnK2Muu6Nf3W2wFNhtfYaYuMZcQ7HCLZ40jar/bHHXI
KTyKut+a7kxBEkj2CJe5QXlcf0Mai1aDdePNbM0y5B0DyX8KecoMCajZT7mPmdTt
qL9AOcCq7ppurqu6r+hR0MXplZx9OVWCy7+oKtUvANRX3sBmx8YcD53GZ15yxibF
nRkspf/jjW9JOdH5iKcefThMGx7d1l//cncBa4/8HgwM/nuDTYoPWSYJxdJE8YyO
8toOfdeQVh+Xtl4RvE8y3kI1gLpk6a0QYOL+vSXpIXi/A97/7EMPC8hGnLzIuojN
0VxbckhtmYhqfEh+uhELcX+C9QFF5ICJ+MIuDTOwJVqFeKcY+OxW3Ma34d7o6TSJ
83gcqrnMJrSNAovVyE2KMXU0IBS7QJDoPc3GiMqobvyaAY4LzmmW+EiOankzsK/n
3MJCY0SKbKArrlfAczkQ6m89XfpWPT1R8ZO43tM2HWWGj+PuEs+Zh/sxwFad7Gzz
4zkDfDMvzWbRUNQ4nM/Y3eER9b50Td6S3P4jFNkVBppumKyHHszQlxi8PvLJBbMH
DMMyWFHlM6AhE4/34wZm2sBb88U2yDMMKno91ApD3F3KpCsEvGLIXx+za0pgnpgV
jCnBGQnH1ywyfqO5C5vgjvll86uY1PoDSyO59/S4dGrx+NRt4/ClBE81BBa7lzRy
zj1pnnn8E/fr+9HKLSmhAU6tpPxDwTQkTAhpFHct3U195dCfelLBD3v/EGyU2goH
7NDyTIY4jb/4C+BXLOif/9fdYPdVE/yK6z+kkUw2zeXPIeLl0k2iH35rwgVS2zfn
b50jQbl0WNm/4HYDEo1IV/ubdTwPxU81PU9jx+nmkVM38/0VhN1vG0AigeeDdzJ6
bdt+OgxJ1chqZ6IoUgetR95X1SxvBXMaUsrL0V6Pbo4rNOs6VyWsoDsrR4XRasVA
lO3hK9O6pS+Tvf+uLhhIDHSm0+25r0X08xxypHQU9HVANOyNA0Qdi6DGhWiS/2Fy
DxHQtE2gQjv2LcHb9zbajqsT2KagXDw7J6wSPnN4lk1tPeH7EO1p8vRgX/SEeIJD
H7TCL6Wy+YbDGO5jAwCMkCQoZP9YRC+rpPpLVj60xG2CAN5bt6rztoGJJPrsXgtC
Y+LXKUP/KaSiEXiUSPhxus3QPBvsb92kvtFf9jImaLuQasyAFIgT7s8l3HKpUKA+
6TQO3hdGeMJLx2RevCPk9MTOCawtTlB1FD4Nokd+d+3hNRtE+rHXN3irG/pniMc4
h+Xzz+yMwcHyugdo5McJQotfxrDGQ4wuT5F2Dnvk91b+smLDpU0fbtfczZ9U0+Xs
H1+FzLJC9m/JNjTXD+qZ4QggAN+KSUiS5CM1akW7/0ytr7AGBFrGvZRAad2mAWi+
on59qN8/eIh7zrl4zN/C14NUoVoYitBvbH5PtbixIDOnyu34dvKf8KuRELin3k+x
9Y6bKBNKv+ijH3ikMsPT/3k3rnMkTH4JpKSVUNw5E3XLPjzhfShljSnggODanUbA
V0n3azo97q4r6Ivhv7uAC9IRY4pGIE82nMboVXeE6A0CkqSMGQlot1TZEeIh84Qv
JToNIYRI2gUZo+gjm0fGuRFN5Dt9VZR+m360NpC9jddwEoT7WMyjMaEs0oGUq52b
jrftzqslX4P/K0NbORzC9JwRAocUkwpx47qE0OpmffBk689rTjB+I3fREv5AA321
EEv5Ytmnx/V/luexolXtkApJHZHtTX3NCOyBfi/Dsu1IbKfU3DBC3cmJmdCLKnFI
77PXI8NFq6d4+fUwqTsEc/kbLr0Sjd0L8M2j6xjkFbusrTD7HCBtHh9O/vB0TtGL
2xWraZj3qDGgiF088lB0WTDEHC9Tt19BCmdBuDGxdRIvoPSmyiCOrIHMrOtZmoRs
t0r1mSZof5SrSgYupBMSfU0zFLrAduqOHsWd+49pYEzU9O6Zw1u3rSjm9W/od1bp
UWvFdI6lemPRJhM4BrBui1ezIuysWGxAsGA4A5gsd9GbOMRWWFysYKa6Vpu8VoVF
//D6Qs/2pTgUaE894Fp4jIBn63m6ad4ZY8gteptTY4JfHzi0zVxDmbRpl0r8qVGd
YRjUcZKMkNKsAw9wCdxZ4AF6SddWeqmW2PW/rV5dPHLaYN/ktEod6Ke5ojb4fyXM
5xEq1VOK84o/mX2xg6pfmcneP17JW8soprQwfyHs2j8+j6ySesBovl8IIWxf9l2O
WwdjD/G8KTpfYQGTrKhBKXv0yDLfgKQZdXhz/w7beY5NpvWpMNBP0CJRHvgm+7HL
PoZlR1EQmC20dLES976tk2iqpq4MoC8jBy+SQ51oqg7cfh8dqxKBIF7r7Wml0fXB
yhZR5i9B9Fd7nZjtp9hGqWt52i6M3h1et0J1WqcB+p1FeA2XSnWBGQhAErcMGbDP
jGtpvzxVFBh2aceWiaTSb0+558cIDCdpAs6ygRrTF/fbIXkN33ptzC0F8eRpLBKT
+Jdluhr0BmOJrSKq/t8hOVaE3AvsWWD5znXu5Wq1ZovzlagI1aHDeqNvOGaORqTi
rOJryXN660NQM0bfSLAw78UUnJEgm3HehxFaHvEgs5tEDb3nAx2kV47TYbyjEM6X
WiAzAu4oSdrpHXbaSVWEx7Fd449RUQ07C30VbWRrzZljfPzsBjokdhAxI8uUH25J
ZQMi+vaNsZQD4CSSUnRcBJkZBp9FfFOlvedb/5vfVKAGJ/nm8y/BdT1b86CnGMem
mSLBq2hgKpeVjFbqVOFT8XDq/5a3KbTFkjr9VzlL9VTSSY3op2wO58mRP7VJgqNz
+/8rnXNABNak++LkzqzUz3Sveij/ZbifXIq/RAHAyJZTs0yJafqJp1waZQUDimJo
uIwU6cAaYOgL9pTg3wW1OjAf766o0Qq0bTggYZhoFbQccLrp883a5s3dMMv9B3zZ
F5oUG9QjqWUkhoQ1GEweewGCsB/HwF+EsnuZP5mZzEQALnqyNVwgsKPztkGZbUrf
9wEly/0QEvfJjjzzC8TSIEstCwGrO0u7SYwYWQzH7jazSwHWCI0IKBNL2P0JOXkd
XQzafvMRq8Wn2G70Nzm+AgpxnRj7JbnedYyIYc8Z4DV+bTPr7YXP+/QKy10j5afC
73KK5HQIg9UVurhvVNfoxT0d//DMKMGaZAEJWLGzGjdlmw7f/khOURkZi4GmCB/f
gOjSbv0vuVLX589Ww0aqPd1TxtqxyBX6C20aGwdYyJnueFwXJjQdb6Eny0FTI+tS
2Ove5snfsqZ0IWkScfsZbM9zX361GseBp+AUkbBuYSzAoHpFn913uPQY9SZkyN3g
IhZQVQm8rOPYIaR7K3GTszTP2Yn682K/I4s274OvAjf3bRIWURG7wZuT4nIBqdcU
Dque3/hw2Kroe7wMWyj2zCwvlZMlT4T0qcLFLmQ7xBJPFgaiS6U3vPA+DPlY2+Ju
c+YLum+PSh0EOdWxXCa9pW3XTwKVva9o6GfKkVjGIQhCvM7/SfySKqE6vEk8V8oE
geQlP86i9NDOXFyi/TrlgzDfHG6rBfMxfcb08qg462sPFdTewKEUBaBrd0ikK5u+
FLhAW2zQZ6Et6A43OhoMS6nwqBxQ5/I7kVvOGWbB246Zd4lborMPACdy9gj8hriF
ZH899n0Z9uVoZY2joHdA4dJk96ZIdcXX5P26l9abFhWgGYSc3rdPGrmlokHHU6LV
q4u2XFIVPAJ+NSsjS0LvtNjE42dDH6NJAb7i8PysnpKcv9Y39Jk+YncohZpxAb0A
4KAm1eNS4JKL/5KGjLn5QDN4o+Sx/iCTaTWifHf9J6pLQGlH7nZlgI6JDc6IRfbb
ZBDsxuPr4itIcPoeL3pKPytstw0+Z36j6Rf3DlsJ2DEuwtfDd9jfrKefFiqu+DNz
WvPJgyZqUZ1P7/Pd/2ucaDtGVGCZiPqCC/3gTlUO0Nv+MceNarK4AUpDO33hAblt
oek4AInuq0nVPCgLPiufBksgUAU5OvphV8k+YY8ZCtw+zm53GByqlrTAaI1muvao
IWu5dbyRF+kA5Y+0B4dgmedJ094NG/At5F5Wa7YdogfdqXs10EYlpsZgJnxhQuHy
LQ43Us5fDHMX4notd2YiPkB4VFmMcVspQHl0TN5LG782S8LHlj90RqfPDL7Xrt99
5m6pJp3k1QXVB2KWwMXI/0WrxeB0zQjGdEVYK4u9CcvGQsl5yYGFFaZJVputoplW
WzYnJha+OoFuehaq/382qD7D6onnRK33sq5eF7IEq2vlLWOoVpMZy15flAz9Gb32
IExeyBSWWRVx5Lo+R927zRFDk+8TRxJT10sX3g5C0qh5X4yiQGgCqrSb3nsNh+2s
OfWqqVPYGOZTsAsBlNz7Ox24jkERNWsf9sMo4iW9qx7NTkXMvaMffvk75De/E7fj
x8CDAJtPRjHWPkyIMSk1VkXd3zOYTNSzD2zB3dLzOAOvsL3Vg8ecE14FRcAoRIWG
XOeKrPbzN3LT8Gfntfu2Cc6igC0sXDKY7saAau5pWihhGnKGsoQdinDpG6g/YAyo
NrODAlI+oWWaIyH9lI3xljOvQXibyr72/8MCMghPMWVyofM3y0P5Myom+b6L1ZQ+
rmWcVAMvMXpoG10osALGkBbGyE0k9UQE5LeR88AzmzAU9ZGWsmT9Pr9rj3VGaEWf
2HbCigy+GYx33OxEgjVkdLoS3NJVNClWhP9r3B+EPG4dtBLrU7j4m3lBOcRZ1fvr
w99W9N+OSiU9SpGWH2YtQEbN4VSC6pz5GIqjcdd0gIhFhyUW1JqRZz/ZvVtB5b0g
XDMTDFYY47DnZnGSooQH9qLUrzQ07thuVA6MuesFXsVOKVVNo07hyFQG7/7sgkSj
t274U3TFNk4xFcv0vmWjsHC10OMtm0gQhqExI5cRPxxW6pVdUkh25ZzFeqpHhC5u
jT4CbabpQNlUL7aPRU2b7uF0RGlBK6gs5n2US/mq60oEHlLH9lhPx1RcSVr2sSfZ
b1o7zOOUY3X/dfUzltDK1wIhgRag95kNemciHEaUphvAJDAiTPFxMLleJdz4D6el
JvexTm/3HtDmHBG1OfDepY/PFX3zfffS09NZrFEgaXFVaoZApYvLbtjTdcrzCdJ8
IQqJUv1K5D2KTvzm8Y4HDV0RzLbqP4+yfaMqneXH/UoFlXenqQwWeRT3osGZ6Lxf
t1WrW00B3RexwUiNmJ+xEsvWRCI1OCbMc/qMFnGnsAQ2d+cI51wciwyvH1Sn31QR
m/CqelxoOn50iwHup/OPrncjDP8RRWTWhQxFRfrkWLeR8jkGd+z8JYQZOa7oind6
tm1gO9MR0wMqf+onKroP5p8XhFQxSxZlYQ1BCybbpwGgylAauQvbvNgPZcD9qADO
r0KDH8knMFPGOI42XqrvBiOn7DqpSr4B17zW7R64g/XgfKcl4zMO9uD4C+fOMMJb
EB+cj7y2x0dsfI96CT9FsMG6rjM6DSDIPDACoAPT5U9F18KGeFiE5WtyP0P0P/Zl
WcYXWgBtBm4CebLVUDlI2D2FP3gUO8X7io50VVqi9M0SK95woOW4Y6s/mddDXgy5
SNiLKjmu0C6v+NcqtO1GpBX1lPesAC/wt+cJ4wUHLvyTQtHuCXylo4fouA6KjCMp
z9lGLuW9lAE6ZGQTdz5a5bdPWUGB/C10kGflZAUWuZc3a9aQ82jRkTvCTsGcTa51
gs3z2ZweE83ij0fgQ8Z4+Ctmb9mOT3CDRSMpewS81PZOH85ri29wuvNHS+qk0f1b
2ia8BALYn8g5F48kLVLr5sfqhkqwtuOWbl9gY+1InnGtxHhavDzsTbTqXOqMM1WR
FVXxGh+3eEC+OJlQasRaMLavFWXiD7qM5culc9R3TToEsD+KXRMf52di42LPBkLs
mebnkYOUUyJzAAa+FuB7Yx1DiKxEScH+c03wKCeyHY4tMaVB1IT4Jpv88LQ3tqBk
EEXyEiR7EpyVGwTgMOJ+/1E/HV4t1vyQIR5ssMv2q6MmsuU1cw7yx5R0mTokkgMg
c0jLHZjBz+cA/ziRx6uPwRMkkuTksRa6gzzTeiFHi5yrcuFtiMkASDnKNLjnOGwL
MdB74efVZYYDwsnmUvEnw4S/gTmYz8QR/HGluAYbxQKBRI4OavyEoP6AfDNLpIAT
Q9ciFXGcsoe0xpLP8t91/pbZhY5vKv5VNS/15OH390FH5dTEs/KOPxx7JvPzM8Mn
Rj/+lIsqaqqGbWKlmNLBaStFZsf39wxScED8uT6c+MS2aVbH1rCMiyGty30Z4joe
X2RxNp8/9Vas39Vp071cTqZeTK1BxyOliqG21iSY43f9ONrtmPV0ercOYTPl96Or
a8bw8nUoVkkr43K7+XnJKKpfbuClZCbGMGB2mmDdu/4RB3ZqJYBpLUbilxf90wtQ
oCLbDUb3EXccfuZo5UdCAS6ZbbN+k2v3+48J97RY3/yWFkrcmNkhNm+X9f+OdaBV
UCEOQCdcY+iDbhr2DPmge3//T/MCI8B2TyCxDsXcKpBjWzaLkl+8Shkg6voleyl/
uBmVS3xJQPxwWjIOLzPfpkG59ALH2835tUA/c8hGq6haxZLbVKBdpBMDYFkn5XGm
fHyMJu75oC0Zg6XYUVZTu0v++4c9ByiSgARGq3kVH8sijScSSyb+9/S9fvt0ypBA
f+ZbGRzqUpmc/aT1HPMxHdrmnTQEubawOovkELRiC8hzba2OdBlcKlhJq3mQZGhr
3rxYeVF1ncSWWPD8Jjhif9S6cKKDPmS8mGLVgDaGBavCgu090dVsBQnsru8ajY51
WyP1vG6M7yySL/AWW8CoHyhY+n1Klf+ImgfDfgOCI7NUwpu4qErITVlYx7mO5Bgy
TRGOgv23sYDtn3ULurooYFnUBBZB2WCKDvWfCss4QvyFki5pNJ+TNulLlxmVkUHM
VNO1PjWNmyJClIVk9ilafee7gL/AxoJt5r1TVX7GeMwZuMCzhfEET+t9K+Nvxa5W
q2yxRK/X7l9jqcVoKpgnQaB7GMSpm8760/5WuiIdnMhU4t1gWKTZgrGfjr+1TI7z
QDfZ9OTQ9pqD9K9vlzlxs2sqso32se4eoRVefEdqEM9jrR+c/8OI0Mg8VVxMauCv
19n8MmS3NAjQY1bFySQasC60ZS4FABTQwWyt1lkt7HN+CAO7rVbfYCW19B1ulT8g
c0Khjrs6dgmqVZDw6dk7BLohaaHPc0MmQ+nzra9Rhqcf1LIh4d7+d+zY6udWPqs6
SpEb/FVznCQQiGHI0e09R6PhunbFWZfRAKwno17K/GnY9fxzHb2EbAHdFr/ixWk6
CJDLmrvWDpHFzDcUKuo10w1ydcZWsfHZ/R9WIBnBjKKdCXXTIKEq+LImvPBT8WEC
mYNMHxvQHl4YLO21WUCFMbD8CHN/FO2tVJmvsaBO8t9q0/J8JijwjC6U/oK8S7wX
mEs+02PuaHt8O4T3R9xom2UvZwQHDFWOMNsPzmobcyqbtIBJlkfPRkT1bFgxZBMy
Alz6JlyzFxhR/Z8cSdc6tq99bgcWWrhFuSiG8WkqNc6fuUXTWxtuBwomHURM/0ED
vtpDg3zPuQIBmUB2UrNz5VrmzSdS0VgOx4gHQ7bcS0+4CS7OvxBaq7WLIzXycOiD
npBgKzdFhDk1buJzWw8f24BhCBSgLtZzuYLCOczc+Ig6jIRJYGpyQxt8Hj7rPVOo
Nfs+vSjahJis2eD9Lal/gx2KvP2QyjQxtQIQzcWbP4j2pf9tlgwzwPMaiLE0uxxv
qpwcF+DNoYoLOWdKGdCQ1TcOgBkYMe8hGNBhS+kZpQ0kR1Hy4CytpFgS0NkcECl1
r6DgyIJhuuQxR4PMH2UbLmGZSikUNkQkSZ1uVWaxTjnn4BI1Fe66QfAqDswmPcZD
tTndPKZ7J8okpMqCBDEZ7xCwarLiEb3Rd3NCO11Qhcu5Z4Vd1k0dEznUtxOKSU4A
3tT3z/UNaD12Hjh9YvCMDHu2IndSBDcSoZpcZq6PxO7Kva86j+zbaJHBie35RECV
BexcVNt5MxbcFmZghJCt4AkPXOqhgsL2QDuwTQizwKW9oJEu3O3zxPHuBhI7v6zK
3uRh7uFB7hW5JUm4S45cCvExmLrSi0nTox1B3kOd67x1SyWdSL6Ifmovipmzv3fU
zJrfH8E5RPVTW37MoE8YU7mpbEOl4z035mch3VIvgCPhWDrNxrhcJvj2f5deAUYy
sfPJRHcOeb21Qo7U06g+tnrDQmxMxHnxVmU8oyjyfJKkEG1N2pq6xaep7gyCLWKF
rUeS+50JmzSmwm1bY6kiNcNcZoCtcfOuf0Av0oFB8ZDol+1MLyaBVxOl+eHy9kna
dY601axAVnLcG73Dp7TAYAnZEACiGnI2lHLivl9XIEFJUdzSHIF+Tknuj14RF/rh
g+0bNS6U9CgxQdR3Cxt/Dd2T3qwzNM+2mGujq/yaGNRbhoq/HQhN+pnss1icKDlr
MHo13zR31V3XZ9pKomMPOIkyZnj1QU2hGwUZic++NLlS5gtC8Q+uEGOlQ6FneCnz
r2dbb0bJJmoX1BndZ9DT2CgETGTnEaGR2LWUO6AEBLWVeMZOZg2x7jeimIVrYcSd
tFnY+jZChH1mRIXW6doTzerSUaa+nYpJfdlqwXVvZtmlYLa6BSc4CKeI3jeEg4G3
b0eLsDlU6kZTr8GU8Yp2k8klQsaU3h+APYSlsADzxZQ6J8ZYlgnSLDSC8RvFwv1d
eforNXQImOm7dgrdZLhJmr+kiKNgNW73Ene9VqZYoruzrfo/VJesYhlS3F6OUQP2
f9VxyPTkhQW1mzsPPBvNtqs+1+oHThxznONpoxE8bd5aibT0k29tCtlgaBj0OVrm
DJsF4rzhHw/Bkd/2YddSzc8xezsxSNvwhc/SKp+bKn0KaFiVv4eTzKi5NUiE1jxU
qvecyMv04KQt6xuVj6a0E4ycYb5e+WpwxRVKXEi1oxd3qbfKwGGw9tOALUT/WcFW
+uNiXlmsOKpabVh/zJKPKfjkFytkasQbG/fL08Cw47IN7hE4/aXpZNQcIsoXQ64R
IZdL0vyOYMuDmR9Ujwb09pStlc8z4uhekm9W0hcARHPTolwVZZIUXnQXSEu6PJNU
2huRMr3dc4IQK7iVVBsjGhMhC0x4rVBPjuprWFWICyANNaVf3XpDENVPx/iHRwPy
KXCqalmcvYS46Yqof8zpe1PEwq2ZMDnBBlgoUl9/4Xtf8FhU50wOGsdr5ay2M3JN
Qul8B8Z0MtsD1Q5/HNYOEyE4k4HO3QarekIGPapxLcecozz88YDSZIHjtG1+I3FP
VuTR41CWt1Ca/l7fiY2bKW99Mqz9b23voQuXPUnB6ufh27jsyytSebQ5N2Gx7Yz5
DTcU90jIC4kxDnB/vE56lMW04s6WcfAh7HhyiGB7dANp/sweYaNh4ZB5BUghB+cb
g5eHgGVSMTHHZxd2pIeiMrK6WmZyWVWMr4ArVeAlcGjeOMXNr6l4e+wihR+oHQGV
qT8MksfVCO85NNSRaxnaO6tQ2aDUVnvcUcDO/ux2GRWdjCbSp8ahvwTqNdFguhQc
QHVdNvqk6n0nj1Mgq3Gb3Fnsf7rOxPg+ySY4V7uGkI2azQLWJDzHEg3Oplx77Oa7
V1dOIfZL+V6u3uDxAka3Bsht8qo4++U055YnAnnTgXltKsnFfKRizPTNLw+iJsTM
LdCweZUZ3ITNxqLhpfzCLf7yCQHxd3F32Z4lwV3SS7dQZdJ1tO2pd0mIiOkYbMlt
DXPpLRvV1oS/nkvbBypUpQD7ogcgArTRTDdc2lvHFoOaafKyJJ67afuMNvQ4RLbV
3XVnMVTnB9enBlYmHwLlbfGCA5V1GUM4EMDPfNvKlK6gqgmplXpg4Qr4IxVJwEjG
NpSWHmfWcoxJA3gdw/crla4GaFaXmhHbnSGJsBcXeELqHWt7dT+yr4Fyj6nfD3p9
jbLFSHSWDOW+txgYewYVC5OUlCYWTlSA62tF8bGbz9FTH5m6IayPsx7nK6viMxBD
gdZXG5QzGGflDVs76d/ScZJAxujg4cgRuQJhmuZoN+Jzrg9sJq3wHODlu/2lalyd
PObD6Djrd4tHVQX/txepnnUBrFY763fdXxPoIuxLwzuHMCUdxw54rvgYfiGJ8biU
U44v5QW080pnyolr2F427JUtpQwmyKvXr/jN8uhnTA9tTvnnr3AobSxewwxg7FL1
DAu8fQnEPyjbF+Ynb2hgcvDCWccjEvvyUBdO2s7pl0xuavJav3ZVyoaaEAPaLcMj
wz/xtRzX3+RTZh4XskoOehjptpZm1z4vNBzR7JD7cuDE2BtNHIOmhtwTMen6xNgU
nMO0PyFVUOETwvuPLv3DiFcsAuqU9P3JWt63XxMOKv7G7DfGPPBVKXIYlt1O8HNz
UBNryvlnayZxdjK+vxVi7bcbQCzMVamCb1OjMl44VOMeJdUUg4IdZJX0V93TiD62
p/nSYJSOqgG6SxKzo7sXfLERjUpjmsk/h/17RHfmtnAYDRzEcntDlx2m7EhhJvEa
t6rFWsj9ObL5YzgxHsj//oA6/qhJYHhK6F5MSJr0pmV9/sdTwd6Mz4158sWgkQu/
HzpAPE4JN99o9ySJiUBbZk3BJ8Or0VyPRfBNJhm5TN0hYj8Ktuum7ERctSFF9Nbn
tSupaw4hztW3sNCaLFAZpZGGa4sHNavXXC0g28lEyVsY4c3BJBzMITTtSEf1TOCo
9Jiplcq6T8nXbvBDr7PXZU0xrH5D+AwqBFIPYLsPoFyoEj9zLG/YJabVeNpw9i62
emD1yqaYNeUR6bEwHSGvP90koxC5nLvDm8gVpbvfbHXg5GlmjPxVODEVd4w0OYFZ
S4P4osqt9qW+rV7UAYvJQtl9NBnI1kmSGoap2LkiMI/vlNa/p9s8J8IUvJ+zA3wB
XgMMLsgYgBOR5b4bAAvB6qM/4swdZwr8wWJnEb0Lq9Fj3EMiCmHQo/b8bNa1rJ8Y
WYD26j61td0JcXKX2pucUKTOHoLh5n9207GE/qdVBK+2ziJF4lfI9I3kFsyogEo3
y/3Y5gtTSWOcI16h4id3NcmUiRlbxyicb4cEHuWIF2Eny4dp1gIlPXc/NNY9hL/r
AIktBbvINNzJE/Vn0diUm+R0w8dBp0RBZeZIKvW5Hv7LryDwlIA4YToea++myF2p
0mpDUKt6Ljs2dTipig/iJFDxR4HUKsVlI4yDy1au7KCvMDda5PFJlVdve9ZvGrOe
a/Yth7UaKIbdqd6oUCDjO1FbcalTtigEr7AgCmS8z+Z+SEsPwywJZBwu34JcgELS
fV2Lt96a1sJdT7rF7V8VWyFbSGbhFjnd5jsSSqRcgbsfpxZhLJ9xBGNRuAqeYWOI
QMG8/I69Xf0kDRPrWCYWor9V0dgBk+d57wvQtV56SZTxN6XEaI6oWHPVLUwbFc0t
QGP5IP41gm4+drjfsafa9fK2UqWMAWcu7A+0umHl1JxpTTWNTEOhWi+IZdhAafrD
YVmWpAmS64iWr3v3g6/cq3Zvx2/7i4SQkrNsDeN+BRyEu69+PIjkRZ39fsIs02Nt
9ZHeDxdV9eI1Vjz1VtqF5ii0gzRhT7unVVMZ1rmXoLH7o7evK4emTkfQaCqxPNHB
FqoZ0AEBEX23ZW6982TqNDwbnVyEmipmUQoR9xPauSeh4hjghARd264yi+oAt6ut
y6TMGy/cQGRaX+bF2mtkpOo0joTaVbpowPJKzD0ewS6NQesz+Z9xWhU6Lt32LIkL
MwAUJ52TUwnsyPicMqDuwnHZJOh5iRvnisD2/4CujU0fy+vk02xYO2IxNsJ8qDFX
LuSWfKeSYAJdoedYS4qrZbCjtCQR2QvXmZ0I4bZ6XTu4EwhwYAdcUSiduBEmvSyo
FIoYluzksj67dgmJjq4p/diE/mTBZTtj9W6VulgrfPOJ/dZftJIgbAOWjB7nXj10
4nlwV+n07NneMxmpD11+OLc0edCVHlQ5G5t8FCdjsL5vj6nRssgPkI2u+WQrO3s0
YZib+3lQr0IUj63mkk/MuQbEmTgFrpeRuXuKT45czYjFAwX3aMSTDEgevr7JSX/h
AlIfgtCj4kGXQjtYYI3g9FhESLMAr2Cqe/R0waQ6mNHXFG0kBAeTfgaB6eezSijl
jDupcKwq1gPSMzdse9EL7yKKh/koVmZ2LoqmvQpJsIrVryWXJDg8W0fBKm8v5qz2
gzbS1tmjK43ET/aSs9idOoo0HjfxkaxU0RomL8v2SVK5n2SVgwnQ4t6KegE6y0B+
KSDwaY8tfgbTJBVUW5LqSCUhN7lGLVQ5eWmQq9ObRQ8YqEkIQov9AYps7kUL1Wzc
wGGyM2tbf3XwuO+mh1zdaYmvjnLaEXsfw/uQiRvPynJaRIUFyNIUh8SbFQizJ0EM
tnov1Ocwl8sBIKh9aBIsl2EXKkyiGjq59xGpO/Nyr7bNroCVCRzXlWGARYxLW9n9
iU7ShMzg6HU1T1KK4yh52TWIShC7t+xPL643AaubASTTZ0pjCOJbSADA74RszO/i
fWIdyXyQjJtybUghjLBuNwQM69eaFyfLErp3vKWJRZt99aIg3yFK66l1P3n9Fygu
u/zcjf/1Uj6VsKBLQaAC4ZHn7dy9LD23yqQmfYGuz5nUk2SgxFsyLKyBdHM4WD10
X8uQ3KqY7vwvSjCgWHKyrd8AIEApZ3nVTvFshVagjHz4vpmWySajA8Qm9bPHxe2k
WwA2/4K+poSS47z1dc/s1AGC8fbwWZdz2WfeG/51699tznevY586P9/M5N9MFpQb
bLHO0ScUg7O9OPlKH81dCRT4VyCaj1uiAtTDz8QxjEmq3Z5Anz0+TbODW0B68M+z
nBk+Xa73Wv1lNd8ro4e5cxj8ZaK1+bhH5Kn80PC/VzoRkbuFRGLOTI+n5VH3Ki3Q
IP+4c2sqYz+wlnO2IoRYo6X/LjCwshomeIOJ9IwPO4OOnyQqP5c8xsbhjkE/Udre
wuDHnWp7Byhl10jMxh6BZdWMDu2lbsw38pZKRtxyf+I+KTtXJ1dPBS2/QYLT6AIV
VzTvS1xbuDn3g1lp/N5tgHxPHbXkMuUiMafHBIVe+1DvzoX0LMxDqlWr32D8NJTb
5I2PQmv4KbBmLk3X71tHCX43eqbpy6J/to0duj/KllB25FsDX2AY88eosTnKIuqG
SsgyTTyBKsWRTgwerp0z2y75GyS9fkZBO7gih1zRCCrQBVUcg+Hn2+/iV+FnttBI
/ny042V0/OvMkbzCD3WgoIqd+BCia6alN5LnEp7QyJZJFeB3UeMMjf1JksJPzY0o
3rkucT03dnXJwVtL/2vCtfOLHWZWVziPXoMHzlpN1ht+aOyu9VGKGNvUmGOy2AHD
UOjzSrdiOL/tlv0X157pTQa8W54qyjkknTaNGhIIegcI6yzVydbvebE2FZLeXONl
oRn8a7j3PjwM3hsuM6S79vYrngR5KVSy3Vmzvazl0AwOJ/6ezCr/amcjpc9WRsin
NrXy7R08CUX3aG4FdMIsv6EpQ0lyaR/y9OTHtsSGyNsapRMPaa6B3jw0STN6DdmQ
lbvpLKofMBPDTVrAKMVm+KuN5NWr1Q7jWypA42e24gZXSjz1IxxykydQ2Qx/ji3t
HueJ+BfkjTB4nMHwSodwi1Iwyl02aOfrL5fAw9h9GU2myojRPmXPa7BKE4f0SmiG
+a1YqXDe6ewtKWKqI+9nNN9x6/oeYGJaBUMJj/1D3MKfmqcesnbL6Y1MBK0V87YJ
S0mrO71Ipo4y+CQ7XPxNWoN1tXJhlf1cC2DK39hLde0QP6TL8LzZUjOblj5cIeCE
hk/tWaRVkPy4vHJ7WmsKEAsb234In0Nrt57E55xSfg+jocp+5hPqtW3LXM1Stq7W
UdoJHUdNNOBb2wgp03tX6yrhBOVk49IKcDVpTHLgE83I+41gbq9TZ+Mm+GWd+Qs/
13HSatisF1S6WvlQSKz0+2cnMecS+WslVEaQCC+XIBSmRAZZpV+A+FUdsiqCmQkR
cR6cEL88n4cer7AVckGLmtuQjuZeWPMjaNreFtTl6CzAhmnsJl/M+0gCicGzN4P6
J11VrzN6hyCAG1UD6U1n/BWOlINbQD7Y7jfNKMGMBOAgcc4lQwTDSX6hWhrThrRn
Blpmw6JTs7+zgTTd6NStz3g3J92+INUsFkn/vuenTJ+wqiIzJOfh7MCL/CwUFeWQ
SKJGP9qjSpxlJzmOCAeSBw+XzIAvVUFhuvmiyUpM9SB/Vz48uCeppH8spegE5o9n
IYL7BiKdAhL1xHvaWHTgVLU3Bl91n4ik+X3AKIAzfodha5HoBeltHYffeC4NxsO2
1ng30Qwl5NphNLCwujOxFsrpfgWv0aktObBTrvtF1IQQblKinWA5TEMKb1apJ5PY
Eec8pcWvEE9jxwc0F0TmB8HEe4OSCtTQNgb1T/y9H1pyjZEG5bfk2/XF6cDT3F8q
CcVl8OJrK21w++ovhuG1UG2tlkrmi3ghgWUE+redTqiCUZErShNWU6vhHJnkKcSW
Q4MFbmqBrFoPazrtfSB9bw06ztDXMdk7pNnPMSMBmAk85yQyRnviuLhYR5sd4ppz
8b/Z+4pzHwwjWGCiCsrEUUX+8HXYa7qiV0Cz48krATagVA3obfWwIZwj2D+5IdWr
RsY6KVyZWiB1VaG9BTFC79U1ClugjEz4NDvTJZd534KDsk/6NwNzT8zuV+Yw7B6U
L6LSn50HWyR8L9+ejsUm+4tk1NMfMZwW7XOUaS9fANcUC2A+pgk3kW07V/5r15km
/pLKS2rwV6KPcesJvSSlpnon1b+zMqjwEAdov1l00VoXGbXsgo26qA0SW+LMaaYl
xwtoXK7wzxu37oAD+L7eS41NE+Ie4miekgLRrgLkygVT60E3TtslyoifoXP3hXoN
v7NonT3tT+YbUTORYlEkSs/h36jSvhGmJ/5xfGzsDW2GpVRDPT0ceGIHPtPc/JDG
iEUpibt2qgTh9Dv8loxZZuivYNljHOY5BYsnbXyb7k3KheDGM+p7YY+s+pOQcT9g
F+V0zmla6bM1t+/wS3ghMd3ex3uwzxaXnuRcu6qNpMZHSGBPM0mjhPcSQNnbIYIK
qiGEGzp3cWJOJY+qkNp+1yCtx9o+xsKFnyC2g4l7UHe/p1TI1ZTxupv55lh7slw4
fmqP41jBfzknZctb2RtSPxKXdbYfrbhAQ1TBAFhCIArHRbqMavohWsZr1TYz8wT2
N5Qp4D1nUZqhTG2o5VXPssGR4ljqRELuNFFYQtssM7KBo71b1Bczafvt5OuoFNXt
ierqcED9HNM9B+my4luS3/3V1IEuODHcY5vWCoeNfJ2AqHjcqoNgYA2hnmrcIGds
npwcEojZ+cgPkgB4RJscWfmLEJ7PDxHOQj+S9oigqg0FnxO5z/x3pV7AevJ53tCG
Vbzr218x9TowTflU1Gcn2v7JjAeI0giKC+H3daZotf2/4DYcfkYnyc9b+PtSVXTI
zG40yTJwThzw1OpHli/aEwRB9YNCWTYzpGKB7WzQOOAzE0hWoCUMnqLJbGjQEkT7
cf57kOmBa+M5gWOw42C441yLRHr6W9yAmv0LQVUTVcSVbXFCEbg/hIB5bthNMnnN
Ot2Gb+0+p7vNsVe481aK2KlOXsmf2jrqJ5U9KeIGOQS7L5Pg4hggLBhisgUmnELI
aoHEtEpfxAwUMAa4kBwkHAJmfiRFrAKJu05jqJDniy+BB9HmE8UDg1mW6BLlRxb9
GXY6W0VnXFY4flD5WAb/riaYUlyRq8DXdNgUKzlTewJ+UCM0XBNqttSiU53vfea/
l7roQ9aI429D23bU8c7ekFSVa8fPaS413xmC7BYCNIcUGT2VxIyRUoA9xdkuOBAK
dY9ew3meZDm2YwdNCXSH0vcboNAo9hn6EdRA0utwbzDopMpsIghUm9v9PweZtw2m
ZCND3DvbOuFZhrh8I44mVkgzb+1TnLtORzUGd75lvNlrdpmdO3W3sdXaOZ+W332b
iElghdwCF2HQyHz2OmyeMPqVLB7/WYHy12nGRO1894oCnCIEmd6NiFpZn+cMFsNH
pdwBXrOYdoNK3JSt6pj9sxinjk5jFU8Wemv05N9eB/YelCOPcpy38IT17kL3wWPy
8taPH8BAL5/SaK35W+EKVEeIXw+0YxSz8WSGrOEbck/8vJLpKWBEGCXiIsC2IPbF
PmtLICZ4T2IBhC9jwbEDAlQS7zbm4p4y77BsqOzXTRZ3ejoW1zM8SBj7yhnIOyyB
FCIKM6zozu3iIqvBnAJ8kyWEFVfbXkP0PgI51/CTY8Vc9M7GlIysSPihkzCyHdeX
35G9utzlHJ+HHMAUh5BXaVsnn/hbFNw30hTESKNKb9ZvoLS4Zeq1BKGN/8a1hX4p
vwRInFXN28Ekp/wIPoqc0DJJydNpFQFxS/uC6FIeOJTP+5fGE+BgQdd4nkvJet+E
pUNEPHFty20G7AFgNkUuazcj1Zv3JvE+ssg9L65B+zFhzwvwfopkMt3JMOHLwMcH
gcxwEyI+LpEVGFav01e+39Ab79x/tqWJSG1oQVHe3jOwpD6z3ftsxx1f29Z7DZl7
7vz9euVzT/ILp14g7ecXPP5SsTVx7QFm24SDfJqrxEJGwjUEgPO0hXY/3+TN+AQT
mGpiJmlKWFcFn+1gChe1Vs7Je9xTm4hocF8MySQdKURDPqZ83ReAbqomAl/qXOkB
qP5mE0+srLZIZMxKXNsMjAcMpoQzl5tAqE08jXceeWepKNlg603qw8j2KNoj+lc9
+smmBLPK7PDnxwky0DsHPIpzuocIDKXjpxMNcPs4mlxP378hfGqCbLzxYB3NNJeg
xqq5+VPKqT+lP94TOL4P5haslWdUAvAWwts1z1mRnZ4kr7fvO+Ze5yUW4xTv4xwG
gwFUV4GT+nwX834DqjO3RXPuXaHfBR7/r7lrjVdPQmz3QjuLI9XKCZZX6G0SbXB9
xKBfXSxbnp5zjJnRpebhRyWRnttScCgMcpmDgSYXJvGwi5ul8ejovnsnI5daT/xD
qq8Y3oA6u11SYfARK0cLSaI98p/TpiHNsnL7tTYb2qAzWClI5pjy+e+XMqWrN+GA
ChrZ9KDft8JvSfmsWV7WuzdS7C2QKdApOGviuO7rECQGyasJDRNUsqo/4bQ4B4dO
19WpFAJczuJvrnTAnA8dt/HEM+orOn9PyF2d66tg+ksPiPOVX89TmM4c3sH1RB1r
hk/RX48fhw75pYgoPdkmNUjY1NFS/X5qqp+4fp8jD2G91DsFPPaMsIymjEOST2dn
JUAp3uHWr2S/qMVmEH2jF722vIERmSZelQFX7GInHDg3cmrAteNncHsqUzUc5NLJ
5s0bGSLK5eJ8riYDyiR37aJ6RJwmoSlhr/ypKWK1+01a24inoSJCBstZ2IGMFad5
ZnmkX7qdMiO3hRY+Vw3tGpCGwDW1n51FHsYeQT4nUx+peV2iWU0fT3rAF+445VHU
2baR6jieZoPHZuaTnGXmmjYEtWxzaE8QY+0CtgTHIAGdUQtzU9i54TqF34tBLS3b
feFIn5pjxQJyIrcULPo4oEzEFdYKoteQqULgJ4PZdbTBEW6aSTsb9uQGSAESkDpW
q21rZ0Tfww8eAZIAW78D6YUKOlvilDjlm/fljkH/j6bKD7YIUy6vy6VaBCxHCW1T
pJmZw1yhZItdAYtXRS+f19iD8APLdChXOHIxEzh82X55s9+DDEMeYaFR6+6a2hKg
+UeicDUFYTaZkbFK5YuxUQLR6IydsBsJ/pBIs/W0NjR/BANz+R4E4vLoragGQD9J
yB3RGa5G7CNDv6IARcFJCyABVA7UO3hYnib3Nj5TP5kd1fIdfHGNzMQmghi6XobD
nhnAtBYAlZMuuEK9LciHr4RoBmCN1OfvFIqUK6zmb3BV4kVU+LDujLv2WEMCsOLv
BIAtFaA2RzvBTUCBPmvf8tJbwdZl9zruS7EXd/4Ax/2ZJkz87SFOF+N5CJuYIiYb
tHXYjLEd7IwYWFONYdJGZ3O7PghwqKuhsoPdIJK8soMgpDk8xvdnRoqxDWH3puRs
w93pWoMSyO8bEMoUxbNYAnEa6Yv3G4RNDN8WIPHZIW9saUVtKzCUSjfL4HTh1AOs
cc5gc8xqTcSRS7mk/5vot0qBbK1zGwkGvulP9G4XbV+B04Jprxr9+R7JQ56waU2+
LRmIH7SJGYbYKXJpNbHLnmgrCxKlJ+hhFSIKsVU9v271E8Fi2sfpETujqxm78j4T
Hz37X3tkDCXVxEMxt5T1qRsaIlZtxJwCRtK2wEBfg28qzkSm8SqUDAzwVQx6woi5
5vz73xwMIHn4H8yq6XQVTkdXoDHHSpoNlLl+X1Lbkw6LEVgtLs90Wd8VvYWAmoGA
wA6PM17a079dHC8ESuxHZdXo13Yidri/RqTftN3sJLzUSU8Z7poI3MM9wvuhm1vi
KcFkz3DpF9M5gSkIn0iIwqfE/njBX5Teq3dbBnsh2esmN07dFYm08y0Ni2aLV6sz
QA/SGJ+kyFyt/smtv3RYEwLIW/+jr/X2lE3KIh/J5AoC3AfZOLv86bHDkyvdfJ15
qAisfDhr4XPZpFkg/O/YJR+ZRacQ60Hxr8BxNdYdTDlVsZWPDMv4VglSjZLkopOx
mk9GdMjivneQ8500IAh3C3yS1h1dmvgcMwCcR8suNVuf1riXRZzPG/FsUiMlVY3V
i9cYm6KPMMKzIupCV+xhSuHrM90EUsrrj/UzNQxfUUolvYrBFM0LFGLkSwBnUa5C
qK5dm/6z4vzkLuGVmWX26pNAcCFmtvM8MQsHOKwbCRL/d7GvouDeRONcuRbG9LjS
j1JNJFpRwKoLUhbwMy7mCJI6FVw/wBXo2XanmV0t04r1GAbQhc05ZCy8L6mTGCYh
qtvbc8I+4o/VDsWn7WF+oQlSieHtS8la5hPc9WHLEIyFcAWJJDgauDT1gcGJX/6U
12xs4PyqLQYYPv8xjtRek5Dc5VmpL6wF8qhvgc8kzNDFz55m1O/YCN9oueyEfT+1
1ghaEAPLElTBVh1ovZ0n0bwPyZpySGuHxA15Vw6hi1L2Lf523d3pEhuyfPWso7bf
NZH/WBtyNVp+BJ+BSFbzCnn7VNIhsk3oZtEPCSMCOUuGfbSpTMZQ2+UaBwpa24fF
9hfbu+ZT3pDuxUvcbihzdmgLDmQr0jV4+aTUrp+sG9y98ry3K0cpE8S9SH81EqFi
nLy9I+5L5P+yGv/9WXHbCoPBBWV0TZWohpc2HACBEPLNvw90YaUt8HGRdZgEQ5rv
j1EtrsIEL6n2LId1aCs7nxMynwLw3e335i/wCLhY8aBEVKRkSbzVijrS7jeVB1c+
8o9676NqbZOj70uG/xAM27Kef7wXQhmwXeiUrWX8ate5GMF34Tslzh0/YNscIPGt
jvc1+dY4MrGEqQLw7atgjobnMvI+vvhVSnL6k9tva1b8pNg8CaWvMT/MPVJa+Wf+
r1zwCuEBDnJnOiLHpqvdU2NSl6FX5kByxuLEwwfWP7AfCm/mTp1RIkwokWym9fMJ
UN2sZUQx7gOptFD2pNizYSJ55K4tdKmDHrq7jN8Ceoybi0hJC2RTlYiIcq2kIyLE
kWHGdkiSIojc3XsnAup8zDPPKN5t1af42j5pPpYJioFM9GipcFRK1j0/SOzuNF9r
OVTchBUSQvqtENMhyyzBANuC+CZ6P1Nn3pQiONEtQQPM1uI64v0hGnpKBBdJAyis
A0wfo7Z8XE3xvbRmzxjBOmgd2yLS3au5gHtnaeSEgwZ3QiqLjhjyQ+r67NoE6Pbq
YxtaGuF1Ctku+SLBjPIsNFmrE90f1zeMMhKwlwQYbCwqWcUlFceofpzu5TM13HTZ
qm7yAr4LYTtoZrMbr499d61zJwCsNCTNhAhc3/ggC8exL64/DF7IGoF64Gh9RRIJ
E/x1e8nRScoDjirTGNeKxmci83mn0Cn78SOwA9EM9/mj3bb+d0o+F8NY+D8+l8aT
N7CFJUpg4bVYHJGxpDE5PN3OL/bNyEmLLwrqWhwOxqHHztUxUbky6lAZnrq3FX0G
VcUthM3vsIK4Fxez4uUi0HjBOYntOyqKdUJ3/EJblyBU2rUnZckbehtRnWasOakM
U1MqVmdAeP4Rixd0B/HffQ4CtBpUOLzcnfeDBdtE1I4EIeEG8NG3a90czCnMYhig
ux7QjKo9pamUTfqmEklzk3zCn1tm9xWPL2fQFf9XXKOxfqmImfuo4o173x6x9pux
ta6ELlJXDahW7vtqUkbIqhoE6z/X+UBOn44X2wG8EgdMP6g3XzP9tCTWEwZK05Eu
B+7DELa4f8oJW8dQdTarQEJMc+LRHrs+bKrAaRfZbRGvqgyLYjtGzpGB2sIcH3fg
dqoneWn0qRJ9L1zDpTr7FvOCKlUspnW7QpqBV1dF+1mjsAUjVzOer8X0aO24QF/f
MZJl6LrNiGno2mYQpipYPNxnQzd5YZcpZwpQUHIBw0KEOaZSHSm+2qbwQSEqz/Zc
h3X8gmSFBzFvvLw8Ef+GTMtkGlnfnm/0BVgqzj1xzNtnc9Y5jQ4SmcCUMQAzpYn1
ppAx/up8VqiMNADiKIk6+jpYP/KY0sWVh7ihy+dd32Ykk9zsq6B5RrhWuDLKPsCT
6z4AW5uNg37vDX69fAva0ETKqFIevyD4wB1/lNmfgBSF4FAtVEUhsop6hQfJVJaF
u5buocyfXFNcZTgzChB8LjUl2+abnD5cdWv4jOh7Epp70Wz/z6a8ptZ9wfVNsVZk
0ngXYSkQDIHcMqw/dG3xEs3caEJms4QaJvc/VMs3ynhFaQ09RuI0m/sS7GBBOoOA
gWqdZwSpv7yLKZjAmhyG8sJEqNHEaIrFweodFs65W++l1qSdLjwxr+zuySX7u8/v
ep3awIvwBCy079WBF5M7O9r4lIv4E17bkj+S1cGlmngd+/xp1Oy7qwkU99siR/CL
k8YkuCjRmjszRa4pqhdI3WJ9Rx9+5MskC7JcnPuY73fUQL2Ym+I6OtBe3NCxxY5P
qZyvPmQztrOfUCihDkcXPtheRkCQShT3zHYyW3TAiLb1JBjCbMaNAEk6T+YC/Cpi
PQAVPSPmIBk8vGkiO/H6NPor0TDOlhrU4G376kzHouRA8fxmNdxPvxPhRvCFxN5r
rjZcnOSUBfQOUOIIUIXO2wL1e/HBoj9NnPVTxMCpeviDFiotC5EkScwZN+RsZurY
lPeCHfSwHOaWx6ugpVfZC2X3C35DgOB4Euqr+HoZofRV4+wr7hXXDojRHzzbjesB
Faxp5WAJkUbBWzjiaeq35YN9GZwISzIUOG4uQ9n77G70xmra2/EW/+tY1iudM0Eu
PuTFxo6J4MaXgahEPgEQx+N0M/drDK2pNgvbxYPuVMDkZvAY0VGjCLf0irgg0unf
rC9nnF6TtiuhYxtn3AYToYfg87kD5sDMvv4R0HceQf4TlBY7MSWcOjOdCTOY/ZAr
Iwxw34K6T4cglT2n4GcjGTUhI/3hVZGpfK//KJRn2Ajycrxwo4NGOX0u5cNfrfWf
A0fh+XpQhonM5cjCeHDqdVct5W3IRwsogIfwUv19zRgEweWEUFrJGd79Tj0t2vRD
PiSTxyKOBWGOxXQ6JwYU6WZHK0H8yXBFPa1Nu9f8BiIBrS2LGMQqB76j9PjoHEX7
JkMr6BhELTUewpZCZPc0yUKQ+YNT6x0y9hO05dWoKoFCZnpCctsO1doXDyNvU0vE
8V1uANa8XeIV89TDc7edXgcXC3uaHQ5ef85HW3iV9a13XxqYLwyBNp5WcYQOu4Jr
QxeI3R9EYcEe5y18icyxT4q6nfy2/bID4xL961ucu6/5fw+2iH3yjVzyRTjEdz1F
gDLv5QpQ33bcWIq2sSJR1rqeeWgp86m/JD6Kdbs4tmb/mSttMelz+eLtfMOYxiUp
2vkVfhtec+VpsMJcKgeLHDzLpViUksF/B/b67+L3p1X02sFEBzbOOvHSS4HN5QLG
QtpYA/v2x1u69hfyjjiHAI20IL+D9A45sdaSUKbl7JDoQiybzZ1dI6AP0GiIN77z
KBgJodfrOwZP6BJCrS5+xoxF55vHFWFCRDA+BI0y1jqYmHkCvJEURXZsFF8feo3b
BGXCmjBNbkXbL7JvocjWSOa35YmWwdhNmXDUPb1/tINocrU8atT3Ot3EOtzfPtB1
qArUkLc+C4bh0UMfTI1+O+bo/6+kbApKapqBcsstEYfwhZN8QR2Nkts+7+GvspEm
inKdnJGBn9Zf6X3uq7cKe9kOHf0pTR0JA+HHHLatXNTHzWjzKnnz1tz4cDCzTCH5
QRIiYQiwIzM71JDqMZBu7Kd0JfSCqdkcQ7dnYnQJBB+vjQvgY5Z1GVQg+qz/m7M8
rpwYPxUWI+EMZBM6nk5adBkC1iFr5kHQqMOlnebOAntK9sgzJaWtKEEtQh7hvOj6
LI4G0HsmUd2Aa/EwhHfMOmh13mLrw8d9kygubaTrfrKJWltzwRm6TbK/7kHp1E6K
UDmNWyfq5D/JA1GVeXCuaGF/8BAiWRScCUlij2N/5MbdyPRTYdczd9Fsy4GhvXO8
M5RKNEQKokX+19RlCCP0cfpskzyWRFR9yAZ1dvPr8hDgdzqrJt2C6NQNWj55AbqR
iRNNbXg1fiyL7UfOgoHNWlLyJ0mQ8Bxs4FuSa17nleq8H6DjS106mcDjV4rPDs/U
Sc+TedBFP+ULohIwT81oM2FPGiDR9QVEi4TkmHhtcp02vvOHiO6Bhjddihw0gCj0
c2svNso4fubBEv60VmOMDADE16tgVdKEqyDxJcJSY+1jiw071CeZ60D5YKAjs5kA
DB5owhh/VmRWPiOunKf10FUWQcIdXIomQESyTgcLs/WaS81QdTAarMZmhkKDeD8T
O2jta3G0fwj/fNgCQ/xJ5/eAdk+5TvE2O8Aulg+6mi+It3xYl+A0B3hHscIj7hAG
5F4dXrtw/nV69IGYRvbxTdnwLJzb6OZgtMfOZmIIfufUSVpAuEc8csl0KtUMFNYl
ftuAOZhDs/JelcMdAQjWo/na9CJHRMNGTHHh/qLD526P8vJDovN5xI+fhwT0AnPu
40TiX3kq+kr77yBPnO1iuYOJ23r5MiB5zLmaYgs/9kEdyaLKSpqoetfNhqvC9HGV
sjc1FR7gfO6HlbG3IT1vJ+gM82okXB1Bs+ZrPzN7Gyin/yjZ7W/sRl+nY7Mbh1LB
UFbYtdUjYfz0vbx1ib1shd1KnaL3A+yswvyqSGWc++DYJRtxoumtx379p1eBURvl
pnEz+GbAI/Rxc3JFz6dTYu3kWxI8f9/+Non7Dd+8L9imbJoW2UK353ago30JMqyX
tRYPGgp2wWTiqdUBbI+seJpwGjeGy5LlF8Yp7mZ8H3AXh5KLSNiUYkKQ90eFIRA6
1HNk6r/nwB+2VPAcV7TMx4hTPTjFHX4R16Mc4imJHXH2VMB5dUN6Gektw0UwAW7c
MMONsuafPBh4S8RoJ8w610hOAmPKQtNEPc6inFdwrfcBkbYsshjs7XokU1+yK+NT
H5oTCabXIa7uTVctEGGwwL4nLKNGTUDoMrVU42Pg7TrODG2tIBbFMBYyUSfvwzVY
HFgJ7+KVQhH+ACFiFWj0AibegIJnhgjcLUnXnw9FHxjDcWMp7RhveXawe2LrEa81
9LnYUqOpOsvzU/52eCH3ldzIAmuqwfaB4RVfCR35pZjhewL7vxA+se+eUzS90W8y
VpBvJ8b0gb6Kt9BCGNi8JeK26dFotusw6a680dtY5jBD2UIBmzA2LS8gVIe6PxeV
V5hu4aeKck1IJRtT5jFsnHaHd6H4D72jau6nPFF3lZPBNRM0XXL8c4IoN/RPAUov
5VqCx4SrAVMzJTwKfH6mihTAuEAJnMGqsiC/B3uSnhnBnXEguX58N4+/C5HjHFZv
3afCUXYk+FX305wWYb2UU3REhUBx5g0VN7tElsHEE1vPkAKuv433XhZFNBW4tA/a
SWJ1xMxFJtIUBl6cvFT6tL8On2LXlSm7v4JUUUkKs5Vi7FF57SGWDpP8o1JDtKk8
1vhsXBJfyc15o9+IJqCgqUJd8eGbsqJD96GZNg5kBWpc6lx7j/Mb0uTju3Q4j8AJ
SkAHnyA8n/VK2ykO/bVzoZYhAdHGyARWvFb1kY+zZrS7CYTjNFjJm59iUDmhbJh/
CPiFfwWGUtBQS33EmQQqAOftRIGCddxHieAcA//nwicDwd3zwXau4JceeTXm7tBa
T2Flkg4yUtWHF0AIl1/QLZU5HFr10zlWhqUxFl/Htb0XwOc15MqC+TNB0Hcn+1da
9E6M/Tr88R9GfBDKdN02p3V9egm3n5oI2M0+ghEYVBh96AotwUSlhN6rspaTIjUy
TBaMvCCgBLRf4HLsHQdvj8vFZ1/2h1/T1hXoBk+Ujo8Ol2ab+toXxAPag6k1FvDx
YJX4ArhFVauPo9qtuy5qGeb/anLKZ3Mdz6Yk508eGWS4xHFQXkOImoDinW7Mb++4
Tp5vvTZcwzVkEb0upykwaPgD5P4xplgYeVX567+eBYnRP40OeWNoAo0kUmGvGYez
gYbCu64Rb1Xh4iaxgzFD8igX7v745yfaIIbkT9izFE1cc6WOhBf+gDNs6F8UlZec
JuUBsZb7ri7A+aJxXZncviq9srcX6p3jckwf54igVfX1LzqmPzMie5sdJMaBn1lJ
EBdzHZAZtKmf5YKJfsF2BDXRN4FDaK+9BJtV7vLfbfpSH7oajuMVLvniztFUzP5W
8dQ4Q6QucXFe3pUMimmmC6OR9WK24cTygcxiSRaZ0j4inREIyBoPUnv2a+VnZB/Y
gzRjg6Usk+f9dAWsdFStU5IuapvB3nXXp85Deb3WIAtpgiRHYhT4rsY+75xhXvIM
h5wR0S5s+cxRzaRTtXlPj5KzglT2r3jIzturEn18m2igZHHs+SUWuEnqFEmPto9+
5NY1SBVT0C+bP+J+PxdYL3RXvCKsDptR5lqu9XfXOCrkDC624plh/4/bDuGpVGyP
Y5CVY40zfj/sgvvnIbGY/iB9hs2coT1c+7KrdZV2s78Zr+pu7jvMhNtePbONGPoa
7HFnCJ0vqk6FYEfoGLmqgKcj+KMkQHoSV21IVuEetDSXOcTqd3Q3CR482t5cZrGi
uEXQL8JPJVidigqKNFAsc/Oh052KWn0FBsV3/8tHGL8U/YFGF4kxerbhj36h0Bfv
KE8bp3r81kYK1gkcdvhlJZKaME1vofWjKGPC6b859FxSs1dI6ZM02ANxRNKOjraX
WxHdVdqwNVkdKy+L7htCZaqTpFfmkQjie8Xzsm7o4fx4uI8wDpF+h6Gxh7OVj4eK
x5VsIMn0PuRv7st+cVlgXSNEPHlktqbNgrUcZSdOpNJYCHFC0Q2pZpKwOaW3B4iz
4qRec9LOlvElU7+AdWl4x/OdHhIT2IJyUhGGp7z5NGAivHQH60gIdiOQkljeuBwY
pptynivC/zWN27X8ibryKdCAqCN8TNxufKQx3S1L50RTMrbz20WwhGimbCOTUv9h
EJMc03NXGh5wSMvDaTPQfvIVVx/ZaLV5KDK/Px/6tYM1GbU3EU8M6SGZTFpLwk+T
I5xU3RGgF8aD6UEg6/Th3QX88L+1093vrAmVZEI47iKvntX4DsCY6PdgGA3/2Hxp
NATNwEo53lIit+cIoy6COY3RLd2PL2tVofLvCS0Ma4yNNVxJoQM4wDNpTVTtp3+y
zINFnHcd1CpESEYkzvMBIw3/WvkkF8gxQpmvopr/lssN474tCKX5NtwXVUlrPiBg
kN53iaH2gbhtoXpOdVnDvXhs2gfukspQNNl2kOgo73G4xnYyzai4KDqllnzEapj/
lZgbn/5Q5qKWFOhFiCALQ3czkPKsd2ovhyqLlOzvUOgDGImBM1SStEnE4tA+NdY6
2U+AqbrTDyidpvQvzpnLh/KVvU+Q9kfGZ/TRf5qs3xqSNtl2So/LlGyXon75qKEI
3BxGd+jS8nP1sdOsK4Q97VYUDlC++dX23J/kRkTlYlSpyPWvn8SHfJddPU75GC3s
UTTWKT5K0jX7hcT/+4+wn/4YveisHWaVUo6iUDzv/mX50/YvDaMA72bBPaDUieAO
6wPd+OmJ5l8QD0ewZcuYM5D5hM8A5LL213Bd9HC8ARyOAPYuz8HN8FFt1wMuGLdS
V24Z56FeyrZRNLygCdDg8GlYSRoviwUgOlJO4lgkhQN4b8McNH7jrVbnfODLJ67G
6pyNVQaXt3c6w4k96p443+7vt6nXzYWJBZyUUj6NgrC2Mp9lM4BvwfpVEaGL0Rp9
BIHcjDWQbkoTQqJfP1hd076RwFLMf33MQmohtjJXDjG2fqCbZ3vs62XPSvtk9Gnb
opoJoixMt8zUFin3BTiJsXuszjxefScaTJ116rfFrp/aTqDY5mBXuUpS9khlX8jZ
2YlvOE0m+9pwDzx7V9Eq+ahxCqLbqxrHJQs/EsmcaomL62It0Ek51Iv+r6v2ScRB
Eau9o+7DxCOlBmUgyjIQ+m3uV1K+JuGRlxVKCN/T5rvG0Y05tU5pk/2zmEHOhA+W
QL7/7EI8BjFLJWKyx+rQwdtJYfJlMm0nMi2HUNzHWton//tCN0l9ExxpSBag4QQq
wQVBKFAJuBPdNirARadLuUR8WIKWR7zvtZHmBEGGPmpGpuzusaBJ9h/DWdLz8ZaZ
osQUKNr4aHsLZuO5bqktU+JesRi0la0sGr32oM2aZJyuyf1yP9f1eLhVvB8yPB+V
zYjWRH15zebTot1uPndgLJ6dKskYxLtuj8doOZkDdUwCy3godP5bQYVpHv0HgO4i
pLW/isfZLmnUnAii99NyUJlO7n/BrFZMXjxOFcDHVN0y89exmwk1V7D9XROSBF2u
TVR+Ht2fbJKtF+iU1rvmTGJV/qOIhKmPvxgmK9rJMhh9dJJyLHLYsRd0++ZrNDbq
vOIQAd5PcC1UFYN7b9qP9hA1ZKHfuLH82Q9yE6xBPDecM1q2+ekRxx9sVCodH5bX
XxB2NA2lcxs+5Hyrgv36UW/bpiBEGdHBZad/e+QULc3KvXYX+/dPwln4cY7vz9Lz
bJmN9UCZYsdFBjFXX7baI2YNWMuxFAE4mUA8iLwfVkrYOYgbqXIZPtxuBGK4+QbL
diNTsV8qNq7H/GjF07k1sYS3yohpOPkvEMuiYVIPxGclmBMVAtxf3ewcdkJzP3C4
4cyrErMBG2BZjE4VRS+aXlJmn4SpwvVR45bruWKJlqpSwmMO978zkU8uQq0VE2ER
/d+TfwVN07Xx7WpSM+HpItPrcTJln9fuphB2wARQVjyrsBpNzCIp1bkHXSZznnJ8
ica1tG2Lhdf+IjDgr9QaJK8qAdZzwdndZ2u6is4zYtewv+Yflrr41Ox/nd57KZf7
jOHXWIkdBSmuzN0a9IrBT7Jds4waIRoL22u4A00GAdDyA7V8UzHDYYVovqoClkuA
Woi/JI6L+47jb/z0/tnjD3lACKHZkm94CCDWxWtz93fIVT/6SelxeXoKRvm6xF2+
2xWR9dG5c012KOtfdYJleW7IKaWyZ9JUBo3IgUWgrZ1gqszQKvXc4j6IVW8A9Rjx
KmZFQa128wJDCqkCG0qY2Tnl0oXW49ldxFY8qYpha15yQdemCg6lPPmizDRbcsrc
muof8tubG4PB16KzKgSjY+dfYJggiQSpZHS7pkQ0ZFwQ9lpnHXHqQciGmnLAQy6A
c1s/WKiDl5b+VhQWW5fBNa9w72HVYhtnb0XR9cg1gg0z5jm9T0mEpRZd0UMITpMY
WHXfDz/OlPxyVGNcGv10l2I5JDJwYt4uwYpGJYRAWqyx28S4jL1dww/5gYcHnzdZ
IuFfDtvB4FEyIkLm3LKp7grP/8pvuZ0px3c7/1zQamSzVAoLcu9W0qsEsR5jU7ZS
Jco17eD+WbsAPrMAfFc7QM0kfyOwtrXb35zItWr6Y5A6Pi2zj2NHETWWce5352ZU
ciyWSuvMCg+IUdbbdv0IUT1zfPVVD77pTYG6toluD6piZaSqqgcwvtLJ6Pj6S3PA
3XDWuRBn80YAySIeujX3daX71mTeFua1cpHs8Sqf0nCRtKXRXIwmfmZSxqHZmJPk
6kE8QTYhIJSTPyMT2vA4PpOQNzCetpdZUR7YkfIGmAG4y5oqChU4bUaq3/o+FDLV
gYsa/EmQMhtebADKXLR5Gl9xdbc/8o4YxUp6gSLaxo9HurG38YVIyF5+B3xqbqtP
NvdzkV2YL+/6mDOpYIFoLHRFiXGedIvBuhv2y58hp+LtxvlkvvyWeB20Jw9I/3Ez
0wjIeZju7xLniB4twgx8UvUoP/jny+FeY4Ulx9C/5X0wvIeOY2j++bZeZLChYc89
3l35/JCF6HSSVh5GkbNz4ICjikvWMdH8rLFSeVqlklWSd3N/IWOcWo9QUkLau7ny
HoUu3K/oNBGrk1Q5N4jfrohdKI/QMT5SjSPz1vA6461a88uMiw00i+wF4xrCQ78E
S4s0ok+/vqlvB8yx5Zfyg43tqsy3qFJwEOfm25dH/kqpwOdkhc/njBcrZt93md7N
KtmEtLZ8dnFuQQWj2dFv7AIaJUWn4QHJ2ZfRRIbbM1e41Tlsk23/3rkVlyP+LV7D
zJQBwwreLhr7M5KuM7a2WHc7DvGKsNwdAeHw5nhduRrrAu/s2IgrdPXHyNCd4ftq
vqEKHMzBlc4Ly1Z4cwuWxlpVJ6ddwO58+/LSOG8e9oIv+Qq4bD0iXNUfIzJ30x+i
oGCrTCyV7JhOYLilBPIXIcKNjS9k1YvGi4gv3MToELZRGbOXeBJAiMtN8KgTHUYn
5ZfUuZ/IMLkE6SYZjcWizqwTNLOcIGAYs/ToiC8RmKm7c5ETcyaQQLLDIkgfFBop
O/VDvK5AMG03eD+xD3ILltDbTUq/vRrU5VHDdb9firU0mNjq1YLTBCN9LpjcCJzP
LZldfeKWIZ0WW4FYyPZnhmhzKVsQXVLp8iRDA8a/DSFVb7C54HmGWBOBj1e3+2pY
ar0jgitW2c4aaDlzHIAq8Ukhk0xstBccpryeChHU87NyfKe1FwukE69D+xpcda1I
Oc01FSLQQ3k6b7BvQoKNUi2C4RcTv92JDum5MiYUt0lwdw8S3+zH9KqWofyZZeCs
deni4tLv8kqTwAoPAUa5+4soNV79d/e3Pk/Cvk5mb8VNi8F6adLP0G7suhDhjUiL
1QZXGOu+qfPqRlq9HTyw/W+LeDebvn0w3f71bZxoRUzouuZ2wLv2PPVlEBP8gIQJ
arY9EN1MmYbuP0o7m7iugGOfVDB+LEGa4FpAWr+o/g2sBfvYjeSvArvk42oJlG2i
lE1cUTxU8cZga9XazxYART6WVzywPIq3vlxuAhFOJYagyotjuNLy1XY2957uW16N
xtcEEJOpX43Xj2swywt00t4ZFvJJYNs7hBdPviubwN4H/QwPN/v1Y/Q22baztwKJ
+nSwIP3eFNw1OtUbplVOXqOvMBukmjYkehiYT5IMuloLOvtHv8FBg20mTwvZLl3+
YJD2/Ebu9ynxphKOXCsULBL35pGMKs5Y+VW93tY3wQzIF+holnOM5JuynXgeHikz
9crNieBWkZ/FbL2GhzeLlfSv+/wqp+4aGSmPLLhnzo4ZIxkqIbcee3XUFkDwr8GZ
G+kSKrItGKaOZJQ77VnWtDSN1jHmDai8Ty1QqrzjdpVNMRpD8sQ5aOUBysCb0C1N
PM5EHG7RSwbU4qvFUYbE274G0UirXngzvZY3cVOf8rZ53WZ3iyZB0XulYdEwmQ6l
Q/0A8qTslpSfnYZ1dFoQhlpjealGM0YBFRuP1jbb+3AohihkCRfFvjOY8b+kHeE6
vdqcZhW20pODC1OcbKxkkKJGqaQ0I+xUqWz/evHKJv8L5KqCvubtmezXKwXE9Sph
BBHcs8ORHaQ46Om2RgA//zf0pqHcTnO+7URa2+nS6NJHRiykNMazT3YkC8NhdgPd
I6LKhGh+FFFavTyicQyHv7cwyVzTiwfnT6dkKxA4RiGrpyJlH6glUXNySgyOV2ei
HdWijPCZQ7MKFcyB9iV8fLxaYHSmqgLU6edxWg3U+rDosG8M1l7hFEtTyL4EKIaM
Ligm5kT7OobrMxNVKmieuYXPAUcNC9MFloCOVcobrotjTLtXybHDn+Zv84KTwG4c
/Vl2GRM0fs42ymonhBsuLKKCoB7cf4bojnT0L+a1fn7GVPXhJs7DbS77fHrn8PoJ
ploK9JPtWdvjhCka/pGODoo1erq+70W+VogbW+JnOfZ3fRIyjU35hjJffRgshc1E
gIAES2b0pb0t2GErPlNfZVsLIRVXAX9rdWCJIL0i3CRc8RGzKUeLtABf6rWxUiPh
Cvq/5uYbXuPxrpoYeV+fx4f4fptoJCChdqKA3qIFN0wUOOugmgG7gPeghbQjb1W5
QzMJH7X6nF9BCiiPVAdSy69JLqOt7+MwY42ZIOETBd0PqpXLf6yr1nY0x5eUu4Es
LtQ/MxiPb+S/mO1/8tYBYarthx5qoLBKO4QHVGRiaev6tgN+wyGmemDpFOJvuESa
IsNoqBElvzsL1gMcLlro/9BCTyDntHGgmtA6ZFsmZPwytOcVzOX5bpl5VUhM7qXP
NGnoD5/hoqyg9irkebFaRrg/EnmnEV8n3TEKaPcHOmDJcd0XyBMWL+aBHuN1RYK/
QCF4gtqqTraowqH1iH4xD/CnyMu0Td+m/0o8hLXdN6Q6HHHx8MgSxRTRPh4A/S9O
o7unwVMn5rSurGSzD9+XckEqxXnw+DlbVAMpc/Bjenwn2yD1tLfxtCfmoSfD2ct2
ayf4OAIMBtkwZoaBGWGq8PKjQtKcbtoBIhO36/c/MbJak1ceSKXrcv1B4T00clbt
esSsC2ZwUGM1kSucKRVocloPsrRd7G7+XLVPHtgpNzztVc8VXlLXQ6wp2zplRrX7
l4/MjTSe1RuXPeVo6W9yedlwEnzhMqTCnYi0/wCcHlltLdZ3q3GLeO8KqHKuOVU5
+oTF+mJjgJZOTaSYLfouk8dlAI9iLud9x1d7wkrU3whKLgRP60fcubkc609lmsJO
NA9dpWtfkZ56SVW1LfHZUOhXlyjhv6NH4KhwTrNIoF+EekVbyaP1CXgLZ8kOuq9+
8KJFsBUyNVEcX9jjXdD0+nmqipsAJko+gHaYxpQkl15nwkNst9KiiUoIaTOtW98f
hPuu/ipLFp2UvIRZLdhltQnQ6C/A78n9sOZ6cR59E41pwI3oTB6+ov/lgAuAQwy3
NaEaBJHoQhmsyE7ezj7KSTfNJNpmTGZGhkxUTdWs17hhL653X0ZDJKopEVyeXeCJ
7Xsnu4xHteEO/1H2li8/XxbH/tiNZKHLjaWsdC8f1Adq8c7AzvTITcSA7szP6DE0
heQnwB/d150DhVVrFt/CnpVSlmtUP5dE6v9MPzC9lToc0V9tP0ksMNCwAAwEsV4D
WMh/uGxlI8KpDEZihDA/edNmwEBISwJNpZNfHOCOLkv65lL3eVpzwIvQNbpjULVz
x3yBkL3FchF9Zxknzlmg7Js1W3b1WOS372g+XXglCK+lLYQFIHu+ZHMHjVAJCB5A
D2cEINs47l6/U2LP5AWNBqUbejMFYOPZXh17gMi7ao0n8F27ZYFJwJlu2MpzEi95
O0Bh0nPHKUTxrrugU2ViiB6tIo0u2d4tHHSYE4ThHe8khzai3WIt3UNZ59xqHRuh
palAAF58t34oTRlq9niOzsTpkWPFsEnjUca6fRHsNuZqPxR3kh5Adw4Ue0DNGmtX
1ZKjIj6iI85Z0MrbRy8Bz6uI79Xmub/whoK13HCQHmJZ6yZhIXrXXBU41Y4yQrIp
t+EawBwMY72G47XVugPVBP1SznpnsuRzjGfPqpCirvxKKXvinJXoeh4Us3XQL6L9
rrovJ7NtaOsGdhy+8OLCn3xG8leglYBY2gHsymvAWqAzURKcn/OJbzyLvMnFjmhm
2VujP82i2FYfTM7GbEMseb6rCd9zDBJNAieKH0RSUUMnfWSiAxsgM6v4A0St6ge3
7XHEo6lvdJw9cXF9gP3SfWLmSyUlldeHSZeFrgObONYqt7gI9k0lAgFwgasqg/JF
kgE6D7Th6sZd809Zxfdc1F6MMsCcNjnY6+fX49SkXVam/9rErWaiXqEpgCMO86LU
aynWNbH9K7nnZ5ri8qCa3GvPLyOREPjEQo/85dV8UKQ74y1dZsEj3oBBHha1ZfVo
YxDdtYa91kFUJTNrERpZCtv/QVXNrszyqTQoaHkDOgZ35W2rEF6Gz4IceD5h44m1
rHy2pVbsTQlTaQw3DvrNsPIQDz5u2vC22SYz4MMlFWeeAYsdUfBC+cD39RXxr0eE
fZ6eMHbFNudGfctC0uf1pt7km1l9E/Jy6Z2WQsG2w0Xo8Oc/2HUoVk3J5hVJaQQ8
D77fIrzJUvUJK21HHBCrSwaRIm4zHTf7cVchndXwqMh0RW9UgQp18OHli+gBRGRX
BzCu4xLHOFCzmmAJR4Tw4LvaBNJcWL7uA9ny/I58HdlHqktcEjAt1FkRVESoe0Fo
xHFezzhS5kR3B0HcFHhXovbtOrKQLYkhJ6LgbRWigWF+VPA9fgPvQezWCRzb1+ed
dhV3UTUSX8aoHQ6FNw0kh52Cn3Uv1FYHO4ssH/se+HsflINPn5s22uoK3Kf7LRtP
hCnb5gE8x/HOAxkCBOIfHxBN58nTGsYmlCFqNogRkQfqOYzCqff63Ew/sN+VXIdO
9kQAXT//yvfYFl1S9BPNIQFrJ7fFYQZ278oWooXPk6KEou9X3mzM43D5O+++1kzw
7lvZ9lMs17lfsGZTU7G1yiCZdhAIFLTVoXoCRWgRZeEZa0rYc67ez4pL5D4Q5Bah
icDmnMLDOzTr0n10BNIj79CZNBYdp2JEJ4Qe7ltu+MO7rBFg6vXmKDIullOqSI++
XzfkWoBT26SNIAFp9fppVubhYokizva9C/3xqb7O9GCJjtnxiwx1wR8PRLeVVI3L
4WeOasQNu77xE4i4jM0mIazIIa1WAO60sgG2MZB9avz9/yhozUoNE4Ap3qt3p3bG
Nv7Qh9ZG64GRMVo0Jcm4K7ti95EuhLZOrWngkYQbyY4eQ1WFDucQKIRupw1yrEPC
to1pJn/dprUBp+FRjf/J8xmOzriYbcQasn8zF2LYudDes2eVtmsNw98+DSaQcDHW
Nv9qGcNUI+Sy6iaDruWgZyhvMJFmOezPTY6P7F1x9HWIJW4Szl3ETd46hEr2qutP
JcEjBVFxdYv+ST/JTE/VTgnt0zbieXLVxEPZVTbK0gVnteop1d0THUhBoRmwFz3e
fsCN1/b3QRjC6xOv+viTnutTeQwI6E/7XDjuJtdY0PZEw0QIgEX7juPWjt1nkHqD
RyWX9AAk0FV0z77JgbEwBmrgyNZh251frhJ2ldVS6rShaqvkRHp0U1jMjQmOGLQP
Lym13Z/mSWJ65TnyV1z1aVX1kErY0/vKVe3s5YOuocW9BmTuH/ZlzMprTrDRaNHv
XT7eAjZsd/tIOA+zr11Pb+hg19ZsgNFaMFELjl1LFZqfAdpdfNuNW88TWPAg0NPG
4Pbq3TknvKVCezSPTOP2k0omVYv3d7F1hG9PFycN+UWRp8UmIS3Kxiwj43vqogbr
SD96m9tXr9zGz5quCQP7pDAUyX2EAgK4Kpiq/9EjwccdcBoI7Nx77U2TIGxrqy/W
b7nqikls5UMLrMg7kpKwOQ5d8DtoECL20havrPE3KeJ6pMtxIcX8fA3cWW9UDiGF
doB9iLG+Sx6DZnvpva23eB5zLXW4WpEl5Lo40/aUik0b9BpUAWW6T57NYrP50mpK
V61LlOkzmcrWMZ+piRdUtuDAZJODwctvpcbPdz1gRA+R8ZnAkxVCOTfl4tq2kCfk
2zKov9shmI7QO4k5ZCJmf+kJ9Y/4vUaoWzXuz8zaCQm9UZN4b4G4FXUTXflsWzNH
d/gbBhmw88FXp07svYsSGTyx1dBaR94pjabbL49RkfIszgsR3o+jEH3z1OTxlaD0
du5YOEwSk51s9OWEP2nXKzCcU49gndESj0iFAb/5K58CYWqnsLMoyFf5BDpo6FGo
VBzTkm5FBydNtTg0py/QYJ52/e8jtpsjc05+D22xftn7xtR/mgbe9gOE3upd9avA
gYC1h3PA271r5xn+IA147Yw8GS1CclU8N+uCYBjHLsQebBUIYBbROaFcQ4konuwB
GUbF+HA9Z9YX4n0A5+xv2Nzkfehc0f+P2C5xR6sX4n04m6J1nYJ9HujrA25rvAMV
/Ep5ydRpeZNXhM+e8tMdf6OcOqhwJqPv4XH1GkqdznQOou1aOxpvAB6nn/EHw+sV
edQrBx6jZM/3hnMCcdzXnHGbsLxafLuA2WyQbBjRLLdUOwbx7n1uuKB6QYqC4frm
3KuKLfUrf4Fp+iWDt7YdwyJtMsu2phWRtzBSrGTmbPkPTjjXqbobEtSc4YIJpes9
R6zhoCOnnUkPliDnPatOu/1bOjJcbX+UFs3IyuivMNQVaRdOdSajNUphvFx8KBqa
da/XMxpwDWLXjwHZqqNSXYSwphzLRvjdKxhyg26lni6vyYNOGCpV7RllNfjZ8NNx
ooj8i3QQkUoQJv2HyFjEBDVJB7sNfU17FLmD+3mj7QWYEZRREL/mzcMyAXHjPh5a
hvjcRnjwPY2Q0L7c2BI6VpoPdnq3MDhK/xA7453AYMF66voq81cBVUN/u2Nh5iPj
Lq0p6Ohz+MnHEYrFEIHZrnQsFQlPxC58pu/nE69oisia5lxJjOd9sK/1aTpsefF9
VHWGgBztbCsdZhjqPCq0CQk9NGsuY/xFlT/JqoXyzjFzmkq+0LueYMjHkdTb4IgC
LXvdhnBBut0X2Lvqxj1Uxoztgge8VDSPTCqW9DRFUmbxyGwxni8azItAYajwikAk
FpAr5FezlaXUTyakyhh7xxhEZrEzA6gYcBtCIMHap6xlArB5HQkdONw5OvCxGy5q
8+wajtslClGBS2Xogc0xPrjHQyuXsUrcYsz6gSMEvY89jovky2fpei/Yq6BofNl2
s8NhBO3SYh1VmMQ722ShoJGmc392sNB97QFKN/m2IyqTAc9a6vnW8GOv+IONPXKi
qyR1wqbcXx2h+0OclYEiQQO3EidECJo+psPXMxqH/ouwTdzMAjS7TZ/1rHkjHuvP
jc0zLTVloFwfSM3Pw3fQxGI8t2DX4v6WXIP9R1/QK6AHwWyZA9e+ywiYdEm4FapU
pMt9vlNn8Ie7c/71ZMk7Ct8Tb5oO8SbKsSLq8clcdBuqAhpPd/XU/2zcZwd32sku
pQCHMNgi+GaAh6XjPleesyDb2bBDE1zBPwJY285Nc0csHlOwOpinb5+I33Yj48g8
ix0XiFeuTDNcYTkb8rhb1THwzE/lwYtgeYizRdhMms3b5qk5OL1txzF8KirTBfXh
IYjewvEH2uPPRlIFP6ZgijVVdxcSejvJ+aNV6xiIVfrY7F0b2wBN1Ubh0Ej64Tjc
CaRt2cIm8t9f3aIFKqj9cg9w+oe0Fm/PW/YvlT3MG12r1BZsV8+Oroa1zYO/1XVF
xqKxCN5af0FKoOg/y5X8NDIprjeTihHW9n7/VKqphpskPnsiQXG7jeQrFxFTrN0h
5EAdcsAgQhTqI60A/6YKrdIJZE3rBFOalTD7KMuki6c6UvFePM7ZRA59Uyykhrvd
K2IeD+Tf6Fo1hLLUJGzQtxHcJUo2zNmd6WI+xkPRZcOATd/ttSfPBAZ3rd1e+fbm
BGfioH34W1Nn0+oVzuiPal8GOz2xt7OPwymc8UBI/rAFBueGjoLVfH6D/MsndCef
meTVOHz8BnsZA07ODr0BPhPo/j6cIcfxvY8XowL8ZPAkpc9i5CO4cKjy0EAscgmu
W7CeaPtG2rdXzTUVZksTaBrrLFwdphnSmNTpdqyS+tuIbShrEq8g7wijM/VXrmuA
cBDgFbUh0B6/Qj/naSI/D0ZUNB3DtD7l9lksT67kdfD1hYzGQnKMwtcs3qULc++P
cXtXXjPOpveQCfCQzSStEpRZ8vA8cZGycMlesv4aON3oLFbe+uo1cv/wCfSclFC1
mPCTYmrR1skAOuhn/F3UbwLed2vZUVVtJ6m7RdhwAxPEUevS2JFONAha9YdvE1FK
wK2s1lV2kmGgC+R7BVeCAL+Qa1b0H3bf8fd/aHW9UiFtxzxQ9pw3Hns1KOLTo6dk
Hjtd3jxvkbJWAvkHnWSr4IgH8VS5CXDJw4vNReUr0bhMmFPR4/9RENejf9wWMHhW
4Jtnmr0Cw3P7LKW+StrzhhoIsXEd34gFXh4/E1DrqImrO/vtCi+xngb7i+G2smUN
a331KxUYYANhWmVxeBBSrfrGO0Lkml9k1BX7rYnA/ojy1IS1ktRaVS3zm7G3UcnP
usyTu+TYzn7j/pVrfivkgoA9wnjaHWBZVHazrTcuGoC8x9dHfNkuVSLBlyeUHFPH
X933quBprnbQ4w9iwyOxHbl6hclFl0kBuixkTXHTzUDf1EPScpaxv/9AxDu3h7Uz
YRb+o5+US4GHcfYTQzRtNzuq0zLsxzb4cHhhR5pr3k9intQKBmYOeLFHIsEiFMva
alg+amJ5JMzI4DMpMcTiGvsCn4A9NAdgUR/BxLbn+TfBYgxTCrv7IDkmmGDheyPd
JTIYgJDbOGYMtVCMRixfS4j4caQMrzHUCL79f6RxXzND/AMVmC85ZMx94+RFeSxp
cBLX/dF1abj3wIB/URky40srUXmXa6hTQbcEpKCG4YhmFgr1oz80VePKgJ+9cBku
3Si0E38P3Y1LmFP7ByF6saBJ4AXv9TGzTDEo9XRKcpX9kyUkjt2GeqTcvV4pxQ7I
NEq/TqOgxym1TtWnJh9R/6suMrFU+RjQAZNVg//+b5rfexQioRmQ72PS3DTMjK/j
8xN/Nexe4An2d0XP06jKqhBdHfVjQBBUxZIBxsMpzHScg+ba8jtTNf33tmJF1UQJ
pVonC2/F1lA88GHSPO/bLczlEeBzUm0xjkm26fllHFz5v4RrlxGaHgIKzL4YzcE5
d2MDmNiogvQFTDt3PW9lqMF4iZ+5lOp9AZLh5cRjqUzpWSFo3oNe+pzbHUE5zYxE
agwMi575PX+HqYrwfdsW2vZ+bo7KUNRsracIjkXXuUjeLNN0d7tHSWWjn9ntvQiZ
JtYR7D0XCJcxrsYO0bIXDYKCvR2nP625KP7Ne3dIWcbO6Uu3vqU2ayj21pCSx+hf
HeKCXMzHzZztAYms8t1ELPp31mDZTaTnNBFt6e2evK3YlhEuEWo4FLTeaPsb7J07
d9anShyB3dcxyz9HIGwjFDfV6s20AmZIre6juZ5yHiUd88Uj+YA41T0foTUBXbaB
HJH2vckDQzoL1LMiWngImKKcLGOZbdGVOmbqX0x5rtiC9EhGzpNhPc4mQP+2p3OF
9KZTkFzghlVuy8856J5Ird2d8yYLgm1fxEv4ooFdmRGexLkYPjKFGkNFHvecUsB6
hb15GvwdN/jYwH3lNl+pQ2YwnsnB3ZC1LTnoz9oL0k7B04weIPRx6G6uygMGumd/
3jaEcTA1e1s/GkVELJlYxMifGhYfNDee2oDPnvWZKGXadVgpi0YW4S8gTH+KhDzC
ar2DLkF6vF0abTsKdR/RLvyaqsLDXZaTpU9BzVim/3NTg+gZkhJJm1s6ofOzwKCZ
6UTR5Y4ativ9lCEUlqc5L2l9LeiAnXFQjE0/P9ebjt3LgQpfHic/I2aAzYNa+M0Q
bvftJQ7R+GGM1drgbNshLPdndSTQNspl1rRiwvj/v5VCzA32OkLYfxrIc3P2269/
wvXu2RU5mFpaY+bwQzf9bsmu5D7W1xDMvbKXoPnSl7Be0Wu6AI89OTuG1yURCV7U
4gm25wQgqQ5GYhZEXqbM+Aeg7uyOsChe3T6VkPmXJW2DzORfYHzFSpI5wyoNIJV5
RWH2AZDV48Ual8RO/2tXn0f/kpKcXC92YSX/J0HYQ6o6g5FUl0CgPb+C7X4loQTK
4Mhl2S62zCwr/yEq5SpaTfxUj5ENV0UfOJd3QGvqtzbxfMmjcbGK/zRGCzn2nmFs
OCr1XJ+yIDZbdZMP5NGzOKmI3SPiQ22xgjx6QYIZ9K2U65uMjjYHmTewI9zDBaOD
OlCsbI2X7CdFuTUvMpf3MR5p6Qi10NAeZNG5i1UvfjfMJmw4fdtew2QUIJ7EJ2h4
2Ik8pt+ivVF9ldlDdJqc/koCGocbbzOziQnL3qjSeM/Ju3QMAMaHjuflWZnZwK4U
Fb61nlXj9fHb4DS+WQcAzUJFkUOtUROK4U3oMsOUpSCUCfA0ZabYjhrB6uvCs6qW
Agnv89nigPYQsH/0r5H8b7gwSXcbYJXxpnvFLY//32NA2WGG+2lJ2HL97eJdmdFl
KYbFHg9/mqUoRAkwOWeRFAE1WPc1ZuJadcdl6uX2A9YISLcGmzH92/s+5zA4PUVQ
56kOmxd4mC3aDriOeZY25dNb0KrtalrPFki6KarhWqn7RIgWk5Y/x+LLok6yf0hE
43bqJuJH45bkG0qgHtthlPkYuB6RYYngxjgtTYWc5tKGZGl3zYGVOK0G8zRYoJdH
78QZq4UZNWHl+v67+U9B+1uKIf0W5lgIGvUdKaibW+wdW0UQrMA+OHLIa1cPlojq
ya448HxoW00qCdXYclXa/em/JIg4D0YOBGmaBdzBxa/nKxOqqjYgwtbwZzQV8DRU
yedKlHATMQiUBBqQxNP6GiJSShL4CNkbE9BmbdpG6lWB4lGI6JHmGOXg6Azm/yOq
7Cy4/GC8+bDpYtASJF04sdwDxxnPc1sqqhJOu6SdFgHT/gcMjRl0Afe+NOkPA/5f
SA0YN0byVPtAt3G/UE98FE0YLeX7d5Ir7xJwM9CEheytPbh/bVIINBPMqpCe8gUl
yasM244lSGNuc4dmcL5EBXTonzIlwIWKa/040cGUNGmI/8R4jtouYqBCLCxie2zq
zk5CrEDFspey/bvSHbRivsDFl+iP9Pt0FOhFC5jKMnIEn5B8NmUNyx4dFFS1AYoy
UNeiWg8CzrbIu2xqWtli7tMNS6wLXqs/RBY6AVQzLfpSGMYenlpTIeBAja4+t9SP
3LM5hwiAfgmaPMqH5ItRb1lqTJDmyzNEXMYtS77UnbxCAJndBOP8kI9DWvmCrtVu
tFdCNglqY+pafmH7dXkcpEldEgxjq/sxHbHhrWo2qzHzpSwkcWIgof4q8WyItpBY
8Xs8BdhWw8lo0GDbYOS+m9cs3hu1YyoQi1GCOj6oz4ADoaTNrRPAgL0hBt2eAwnk
QyHJV0vzFfnQtS++G2c8d29Fj3jpvbOZOw6zUGkB7ikmfE4ASn7cXrgoieTi4Zyl
DfaMcJ2hYoBPpTCsZyfmyWcfnocDpW0Dq3r1bU8LkFnEXFjMOU2JophXKJVH0ISn
ziGiquH3GSjMvF/Owup6IcrBDduOKFCdQsTPcEkJlXPqUHvVGmVixGEI/dmvcEcK
CqvTNrYkkLpMEshwNgWrDCY8rEIxrZVbuiEjIR0HcqtPjErvbyofyXFgGJe9nXBG
TRLEIz5M8G8FLfAwHn0hQSUcCQF/xkSeQ/mkRdrT5B0l2JupplT1G+XkA5W/xU1t
aaH7CFFqKLrtP+lIa0ZYWzSOMguo3IdQovrJuw4Iy08i7cilqp7RGRoOV06A+4WL
qhslWmoQzMfZwfvqnj11Xc5/zcnD9svnTNq2rYvdQaxXq5qB6Y8xz6fi12BPKK+s
ZZ0In+QWom7tl9QHH/VsoWQT8VNWo3LbtIw1uHcHPZxxJVcYlZ+WzRLjWXj4yisV
Bwy7bWAOer0FcW5HqoeziRCGmciH7KdVNKHTWcV+gHvgV3SRDsR9yqk6Rm0OA7Tt
oEo1jKaGVpZa86++fFLES7VBJV1rsYQHMY0gJVd5vT+93XSjx2iyyrKYBBj0+8dn
Z7020TNJDOblEJzsFKe9DBhJXa4bOxCNgL19MYs4HpsqOkvVAbtq3K4hMmblpzEu
zDtA/p4ytZXlL+kbB5at1Ws2P9p2Y+6QNcGytcB+ymyEendbz8pHfOtzfu0IoC0c
OlDpCnfwCeuwfLkfkG3G+3E0UBsYj59TTCnadNhFRxBRvUtKKu27F2VKCjPnqeQ9
Cj+8jCvTliXMA58gEZPVKWUryY+5weBJGWiQ3njyqJpYp5Zr/SGdSyEm1vyZZl0g
Y++BcXRIMU5zJmPJHaypJTTp9ciLbSwllHR9r81Is+Jq3qJL2hylLssAvqK4Q6Qg
L8b4jmxCCFah2B/k/+WOqFLv8pVyAYbZ6SxChDmKu3LM5GrLkONnN5q8Pcz0kt+F
y17M8V2teCNEqqGJGekrcLPo66NlwMOeDgdX2uGTaCUiRua2HYEh4R/rx7WfgaeD
8DD7+Fw7rDKaHdS2WA1XDqUaRIE2PxahhhjtuTi8CpzrmYMkKFW3/ox6Avduol8Z
k7N0513I05NbYqxeC29vnrXWYl7zPqggpehWh3M6tY+KFKHmriNkUbq7sLqH71iB
F9voQmFp6TGwuBKqNqYePQW5uiH9XKejqfTcEc/gvixkneuu+K2irHpypQQZPenM
RUsqLLbmx58Iu0mMKjIR+IYL8sLjhFMDADyNAKnLjWdgxhK3aJm3BgpAUdaxljZD
VBFwWEv27+aC7HJaZRmGL5kezMdP0YjYlhnMXC+SBdFC+LzhFkfUZ9VIh0HqMRAf
Yb4H03HwUGfnnbefCw/crPlAnigZlhra5Z4M/1y/ucf/thwwPKMXrr0OGtGBHaFw
2V+6cmSqjjwWBANc7Zj39o6O1my5oomeensN0jRwj39q0+JvVoEpsPkKiRjMlvGy
53ZrNKY+1POb+YsD0yPZMQ/NqI1RypWiS/FFdKaglg+SFuPnuQNK74O6wCjPPODi
sSF4+rOB0n8UUMRTzYC6jErGWzgT9CAQYRGxp1YqT1mz0PNaG5IySNLJRFDQdH6j
E8U5D923WOOFQH9T2rlOCjgjIEGTwFo1DOEubHrlVPa+Ws1s3ReC0QAsIQ0k0X2C
J4sRFhveWxpPnKyU+FMXUGC78rLWXWVQ2S0/P56cYSrw7r25dTb5dvtWfXIBF943
dV+9H1mimjZBNLTYrRrxUFZYA+nkSfKIiZ0L/2jv4uxM0iDf4mdox/hGcims/aYJ
Urf92blAUNl8Ox2S3ASEbFxw1EWq6UhM2r0h/fPXhOs4zgQ/TaUoWM/zvxSDOiVL
GkIvEEhLXco9jOD5p3WtK2qcUwCidwNQHnWH32cj3fhfCzAV/uK7OCS6/5a8EcO7
Xi3mTLwVQ6OgEhcdFxLSqXlqmQDLC6zLOQYtRD7TZ6Etug6LGhE0S+9ML0ro1eRi
HIf395rfB6E26/UVsFRJQBh6kbAOgHHzJbG2/C9lPCjwe+w22VsZwBlwCaK2QgdC
yPdUni3wnMSNB2brPMbpfBsoOdSkOjHQ1yCOIkcmx8ZwXKLVLjDCI/8dW4TvntRm
yBE2yG8ceiLs2tjVd1SHV85dqf2O0DDdTKLdDRZDv47t3fLHOII4RyTNQGKCwJZN
dtSVcIwNfV+tKUAkJ3FUyATro5O/IQL6/dw3FwPPt57VLSMAKI+KmTlTmIPyE8+3
Lv+IS+nXWEaH7NqiqmMALw+5TMIK80hWYh/cQRkACIt2uD9J2B4mcqxORAtXfDDF
ZozbZNolR49Ywl+jSbEf5WCh3TlwdD0JhSgkjVDbLEPWqPFCc/SYZHhUtZJnTS4M
wr6DoChibkYK8NGJPM5nhWk+wrW7OzEk5inwCm8ZUha9+f3ejpoINuOH7ivJT5mu
FpHIQycJJPOJyLNPE+iXfiVV9tB8uTy6+k9UzYnLufZd1xkmjvfVopudBwr60Wrb
3Y4PAGuDDS5qxXhMrC2iebVntgd6jBmnlRSi659MPYAdywfEV/CGM2QgPT2DAfB9
0NELmaUGBRMyeoKz018Dm53HKb/p7DcrVSidG4h8O9e+FiglRgEp8bhttlR+IE68
tzG7hxyQyUFDGXTYYFNbqMrhU8wRKMaGBGtXNIYhq9pPvlOnZ5DutKtO75dzFQYv
zsAzHAZQkMhYNWMQ9nFho+AU+dJrMOxLLq3dh8uqa5z8EfFFmvqucdfZJc9/yQgc
h7cnIgub9lZ5+G/ubG8s1ekow6Y1rTxBg3pG9itMYhTdURtajkF/XpICQYqFm7ww
QVd8Klu2goSRsyvEw43pLyb1upygv9LvwClKwtHTZAvF7UfF724GTaCbm3KgKHE/
BgMDywQAYP0hjtJhjKVrSzbrP0495tLEiRROrt87XdYmfARU72Hvf3IBIP91w/Cy
G0A6ZsSz6VwqeDjCpWo295QvLUpcHk8o0pli1HZywlG76H/j/5mKiI7qIMczYPi+
UmtXticB5uyQhhHzekfQl3FB4lhMkQhuP3CrVkcG5i4G5LDlq02LH+DonDQTECnb
VeBcMU1R8jiJFmR4kSrRnQbh+Yf6wqGzPmBCZhSdlCapTYwW79hMJKYzRpN0j1Cn
eaklBpd4aYfl05EMZDXzn0+XWuawnbq0Lxz3fH7xPWOQXnUKYZAxmYQvpZBQopLV
lAd6irw+xXM6cpMvV5zvkori21MgsZwCSxni+mGEO6fv7kM1AiOTIiXOSDG8PnLu
2lKM6qryV68jXOMc2WHg0fcqcdd3u5Hs0hzgHG2WiEu3INW2Th3E8m3w346s2rR0
ls58aiYBXZHGYTKSWvWFb+HAKZJphc1I3keLs2Ro6a6ackMwKHNjg3m+5Otlps8c
HYgC9HfCZ58sDfnMJ8o+CmBCcvM/tYp1MSKp3VfxLAXrQaRuYWhMxmBNPy+GvaQy
CHrTpzn2AAhUsa/+kc/UG5cUCGvNn42Fi/Uz3E0M029mnW//v5EOouIPh8vGVrvH
HonfeHFtk/CyhCHHZ1svVw7VWsjU4VPJjg1pEzzHZWynM2HXJX9x4PhPvFIBg4Oz
eT44O+O/iEDR7x4JjT56wxPEl2X5ViYLKmqjkAkLPiY0Fnv/nbQbvw5CRcJnJOFX
imw98528Mn2v+lSYq0gcUX4upx6qc3MSRXWSkvsrEkgvumr7xZ0IEhlrWlRR8rif
7+PTPNxMrfqYJJcEFch4N149jP5pnSk4t0PqbBc/mUCr0X8nQwCDvI428rGvJQh1
v5mWFtMQscwTxw12AYQRFLCAr/ul00nJZwar7BgpuW3CUs/F4yUQj/cSuuw2uPKX
xGYoX75qm68DMib8fhgz7G5T2In9J247vaRxNBK2tVsGjVTeMeT94P46g+kmaAr4
V4LPpCdXaY/Tk45VN/TcQVJ7TfseHOtb7Lc4La4MP752VpAcbNOwKANVV6adIDqs
N3nOkAuO3qMh+y+srekAMexlUATyKNTr+/LhKSWFLd6ydhy3oq5zmYlbu737UC6U
mznMOc7Yuac/wavL+4Cy++VV91v0tM3zpFfaLS0u320T+P784eXFlbVJo5yI5+Cs
Hf6FzwqMIr48ryQslYM4aCxi3lKbgqWYB4cA1iRFPTHz071ZpC1CXWeKU9vyawXZ
JOwb9k6wVZva9NFdFML2Rj2pBKUORCU196KRG/DFBQoEsKjO7Q7NV7froa4Ayu3E
rMzoWOJgJYhuveNexBmy0nfBSfe0oAEEufJEd2ZRfG2PuGTJ6r137gCkRW/eLBRl
Tb83HY0qK7vYJjPqxE1wTgOj+nS+Alu37vbBr4RvfhQPrUYM978OmkEjtFCdxR0N
a07ghkaFtG6IksEoEbUHJEsMcIYyeWvQRs2asqsdBej6yHFUHyxb+nhXFQZOmHoY
QNd/AuCw0Q1N9h+6Rwx4RJhXobkuYcEVoQPIrFe8MbofgiHNWZ567AKNls/uGoCH
LVF2c+xD4kTGv8yEgOSj6BmjYKHwX2bt/Fus9G40l0Ht84r0uwn/MkXjSVLbNtOp
aHLWGiVVTsNGpvJTYkg+iMRLN50/JtyfzNTQAtzxgJnK/rmhivC/4m6+3yMBvyME
LNUuq3n5toSnrIwxzsYWukcrDe/eDxangdp56dWY4aop8pyGGTNcQwtDqwPW9ufE
C/N+/0/5ZRdbJhv8TXsLO1ONJzxnd7RvIuLnSfVVeI2qlPDtcNErJMJlz2XPfeWH
XnLvIDlmIYU7BxVHj0V47xUJ7gPnot7aSb6dmdL2G/YCWXhIvM0lMYutQEkzDGWF
lYJV5gOAWp5c2V/tIDb/Dj4b3MrqbipYxJrtk2xDXQ0jJaBMEJ8x+pyDohnAxDjy
KuDu9tD5yHJLS1mX3PGEREH1nppKcs/xT0KyRnvs4+G6HwQH0Blxz4uOUF1AaG4e
s4b59Y84x3vMUZQcOzDENjsePFrjtOpybtMrS88YtbfjNif9GPwMM/NHqxAkdnXK
WAyhtvxBb3R5/WjdNGcJ9M0zMy7oJfLvv+W9G33GZslrXaioTd16J0bn/wIxvnLq
OrV+NVGnnqNbIDE+OEIZadpAqpahve93UtPyKrY+EuFWPUEm1x4WMSktXzv2EiFq
liIOKsOBmHzcNs/yPxGDSznNMM1bD5CZJXLd63KN74ZAsV8dLft9/sfuYKk/7UwU
RsymPftu7Ei1CPNUWWuz8Mhqy8CngHZryE6bX7WZctV8d3lkvnGUYUyDhuPTt0ff
/0xBDF8OiaHg5fYBr4LxSfQzezwYa5VjDXv9XN6JOuOW9LNRoYA9SmW6WrIuY09B
TQmUroU0gHK+9JbTaEB4r/uXJHvBYtmk6bBjD1XtwNJN/bGGCnskIJrjkRPB5gLE
C+d4K2w5aDVnfURZgIYyqox8CfEOUucsBklcmQmFQDs5ch4Yok15VPSeE1W41e30
LTeQIvlnWH4AcJmZlSslLpjssj7TYfIhxHXQ31vQRfohp0gj3CPmZ80o0d4SSxLN
TatQIisChPr1I+QXM+aOHVLj0OIO1u2KOHbbSIUc01syLcDFSOHLZ1WafnGGWkOZ
nfM22Ddgpwdqa/IfSGhQIFizhkmi0HP1aDxlpNpijO5PCaQzcCVgwOMqwz0CwjDj
5KOAwNnD+dzr6fZoo7M5oKTUVcqYncvRGGnO4KVlXuX4EcpobIJ80HGZS0hnzklG
kosCHP4t/rv7eRM52MdTgoOra0oIFVUjVoF1v3UfU1Flr5pLeq0U7mZcFQuQ85Uu
wq5KLX6EXaFgCNpBsKiw0JF3xgzhRpDMe8nSW4ZPsUOtx8InmzYo8/vZ9X/TSIA+
4X9bv2Bydgif16uDYPe154YqR5yOC2ngnOfD4QnX9FAnDq43tHO3F4lB/BZZ1dSq
pEOAnBxhTul03dQeqs96hNoDcZQ5hJGIhvBK+70vsbCL0BetQcDaRCIdyCOQpuhL
SiATLUT1ZDLgCOi+HfJvIzqj7NbmRRrFjxpcLUWDqGja30gCH94QZUP6cxsq3hvC
sPW05v40dHzPnP6oibZ8DsGCZr3Wu9aeXVigj57OMfSIKt9dUGfXDIsUso9OQ++I
Ov8dfo4/Ay2nYXvWzx0BN1IPPnk0i//Mv/g6xBMMC6qsnAqv9SM//GRhsU0Gehq3
UwBFy8w+Xf5O+K//3VwW3DRHRSEPVD4HNPYoMpJZPvmBOjgUHC90+cMPA4UyOrxo
gFoTckVU8OLnQbD8pIWMWCqKTuAwEt5y2wMMmdYnvicloWZbRlH5CHRdyHJDEm2h
928OcXyIwf6flMfa6Bn2d1HNY6FuhcCO0PkTCMlJCBujDyeSvueM1fgn3dTKuYhQ
p0GqQeEfA9bsqs+bLTGSF6cTG3QnkpLn4/Y4YLDjJSYRO7KZlATOPcOnvh7mhLiE
giXbzkjuBRK1LHj7URtMfryhE+bkHto978ECCBGzpE1DJ/bJw3C5hvbgl2zyZIv8
qlNkmvPOclR0jUMggct4up9/jLNxgcs1NFVWhEj1q5AFDEkFAMwIWEKiL2hJWu8T
6bu3pCOCqkzGlmKmctqTbCB+lfB+QeCw1jGeX424tWRsRCiczRkj7kvQSC3cGWjw
hR0mD9HqCusYmKTYS3o8ZpdrEHEWslTl9VLWgtfBZoRpVhuGlhb7qbV+47+/clMB
EUc3sY5JlqBtpxpHiwz3dmFgtVDKZusr3kXcI+sKzhK80yiChWaHmQe66m7cRhwj
NfPWa2+y7eil/yACgztfP3LQpy7YXjGNG+iOHNXidcxtCGOi3CrpucvARIFUCycs
mzGYBSEfDEhiJVd9JxN5UIk1m3skeAO83aEn5CyELzr4ZJ9K+AQ9lcAFwLP84OME
c4cPiAL1vuIN7flaY8pSDMonEKpGUAq4VoxZYmRc01SRY33djKRWiOWA4ySb9FYY
H3TIhXX8G4ApwBOTm5EXOtH8cd7MhiKxg38X6mzx/e0RBYMHXrnKwBLDlsyulahe
B+0x3FoXicvdUB6JMACYr8yw1HgHTm4v+bJYuy4dkIMws2DBu1OjABItBBLQOI+X
/jV4Qo57Mi/2mhO226p/pft+lgUe2Y9leSxOV28FJ/5FOL9WAlaVz0jz/meUauOj
asIYn4CKOKWutsuRusQTH8CzFPvsCJFqoTn5PxcZgNWIaB+DypV+JqPKOdplp8YT
D2+jb459YXnbFUI1DzdL9mPJL3D4qhSQrsOEqrlyrqlQQ+6HJlDSYohP1RC8Gm7D
6aMXfLIbgGhrKoKwn/ex+0RX9PR9DENkmthYg94EkbhkBvbUTBdIp3/n/B6KGuR/
pq2YzxM7QvWSDWCaUqzwBc7ZJwh6BevM+za/FczaDTSk+Beorac2/rmcGz+EnCLM
bNO9BluJKYNWYpZ3NRo1a57BCXp+blJeR5SWGqxpbcWmGRjUHwHlqM2/F7W6pON1
XKDRrNQhFplQfAx5NyClfw5kh+rASszh1q3jvIWFMahkQfszT3R4wA1BD2ulNHSV
nvgI8FbMfWQbVEpdwEGjUM4S0upfTpupv3rsYzONDreUIEhIUW2KUfUZTUlr1SKQ
uLnTZEX5awzS+uVKBo1FtwnUkpEvoalAfb/l9AyVdii28NxBl/ZaeCl+aE1DkOCa
nI+PaStlEsdy9YfhnkxCn1lCmc5ntwTJ8ufhyEya6T2L2O/pvyNA9Bvw8ogCJUVq
qTAv7dwSDnp1QEmR0P319waOLT8xyVxW6vIhuzipNiTX0u/wcZiLvpLV89v7DSOA
TivYkCOaeKRi3d0upnXugwiKkgvUlqDp0Ynp4RUiJyIxVo6r0/egBE3+tPPjH5Qv
cRygwtCH/cmt/EN8Ty0RSyCKPa5cPUH6j8NDgwfZHkCL+gGMqTgu/iA8K7UzU81e
6SURSnMAGKi9w/rFktkQRk6KYwb1XDIpVDQd2LiXCtF1icKCbzXtFtaYfLpE3yzm
/TAGEiekwm4cJUH8teAHvxWE+B8L7+vMz41l7oPoc91Xuh20jPum9+3lwzU7IM9B
Dm5MGhKjAQ0C4/Y93Q/86pkG1jF1pCTZzd+AGM6MQZF6SI9N72RPdyjN9kYNJMoy
Iuu00ZuVeXaA8gZpmCEOOviJVGKtGe1JfgVMF28wAQ9dJteNLXuF2BeQVS9Vzmvw
2sCQy1YVGkrL4VOazl+Jk2kjDWsx83kcIANAgCMXsoV7jTtPfaIBXxQeN7g86QSq
NFMAxoP44iuN9ZhRTZb1xxlbm4M4wlyhfAzyZEToy5J8hqeeZ39h2AaPJPs9T5yr
pODWJmUpGomUrsaOnmddegvp2I0tK6Klebg7hw3LVdRdtqGfffOajneLE6QXrArK
VoUzJia0g/0ez6TFgfbHV47YherbJ0c0SzVpv1DtFuRvZhJDrooUBW7zTAc8miJm
0U/KUogFtqAzdntrQMd7MFX2txLlYNykzFQYLmpXSbLO4IrabqgsKMDrlCKtD1Ew
BeJAQ/xz9WbRoaxThHhdTOXE/wfylKztYRco+qniDoQ7LUeW2ce1Ke3+vV4RzeWb
dix4OKMYFb+/CaiC0q5DR0ucu4q5lj6ZpyPkOcrLFj0OaSkFk1S2zJs6HUgiiK6y
Fv2OHyjqQTGRc8umqxjeifIWibyLKjftZs3W4ZoOZ+fG5Fq37VKq1CIoWgh9dqnh
gGp8TutWVY55U2CQJIF69wSkFDlSkAzEDfpUqUhIHMYPpWw1FFrt/STFfSwd/oTZ
JQNU7P2ODmktpVrn1Idx7nzMbtC5FGSeC5I7MfNWcHVEB3dRY9gX9DOp1Dxg9v+Z
Pwyzcpr8VQOEr67Vc3c5v7R5Nf+6tZizR+yr7xEQAfXrqWwLKMQleh4vyCR5Dnsb
0lxV9RKTP6iIfUC/j7f3hB9YZrooP4SPPj3KpMlNtWIZMzSU9Dp8ZDYzhXdQ3726
4Pg/FbA7sVsLXih1FUJRYjCSZ2dRs75i1Mwlbxvx6nOMD7Roniq3p/LPNAGTNSrp
BU24d/Goq1oV5UfacAu0zsqYSRAD8sZ4WnYUm1S5akilv9c10cvodlP/pQO5UYRR
QACYiA/qaGsjri0mypgqjlbQ7d/wMbie4brVYBj2XF1n/6dZN1dzEScHbfPAm5NN
prSNHJZuHN8IA4AQHdcdR5ctPZiJ4LVa2KgnCc3fbECNaHAbr8fpVMDn1vDACWic
tQwMLSeXrFM4d/COCtmIKfdZO+m5jzXGvQDINHXi5YJVQ2OtSlcUDa3cgBoJB3Qg
dAn+dqHJ2/6nXzFGuSe6nszVkGS6b6nrlkbWOGlFDo/y/qbfiDOC27Ag/GTvW93h
D3DDBSyELNsnTU5nVeo80mDt+f3ZZTiRZczbF2TMLZ8BW2it5m6BVO9K/tDQZGIy
5IpWTlnUdosHMbN1UJ81mnMG1M+3sRaaRNv6nB/tr2r+sAxbSzNv52QhIFvpx/E+
2QDEChrnY6ff8nJjyZoj1+c/z/RiqR+aNesKM+aMEHp94QkI+ebXuUFZImhQYdil
5fN0+S5HETQF1H7m4DFhu44E2XRSK8XRRsiLUojW1E50gyK9wCeG2TcCgKdqqSS6
jP2TckLksgk2pv1iypal9mM45UEfgXw/HpWHKMNeVvEPMIBMUbvSOsTbFAYVzJNH
YOQAtorPkhLyrRHiVrC0RksOnUpVa5h31aqCJKzwjqTPA1nVk0XqPqGXoMtnkS65
R/Ws2PUlCEL+yLAh0g4afZdL8phzg80h4Qu7ytOrBRuY4K4Z6SIsuWJ9OKOSkNt7
otyA6oES/73G+qgaPHBqZW/Xkm5oD5pI8Qc6BSmaheBUb51HsAl00byxDuLfc8Ig
Spfez6YCxSkyk88cy7uN8QBzNElrGjCsxgvrUVIq0EUUoSWo2l+Q9qf8lhOQZwR8
a3eE1q29bp+Wb+VnWq/kUxB0YYIvUfHz1rpxnyWz33eb7ftp+IhoQevw4IUS7fMO
H+9mnKq/3giuGpcwOkjczjjbHOFRryrMwa+lIFH2bdIKdmde/Bo1y079uNpu7uw8
3UkG9VO9UKV3AFAW9SQTNSQrj4G6bg379nkZT7ciHl9LYmo3Q7ZrYO+5S9X6EjlM
wSmUWdpFpVuv1nQlE4lfEQhzEHIu4F4xZLLi6jfuTpbpPg9yMIT37BFZ8eOw8HIU
1IsvXH7lcSsTrRpstRznaxXtbQrHni125EAlu1oQDxiOKcM2U3pESUXtDC8nP4Vh
3RpUqOWEx2FUTkkZM1y3dEmtCqPGvwiMw5DWfrbbz7wqp1r8bbBGLxwPpU6XsjDR
31QLLcXyT9meW96yISvOEoATEKN3/rTdM4R7OH0SwsGab1NPtZZzXY5EBxAP1h4X
8GP09j823hzCK0IAGR5ixQA9CbJWR9rqRmRCiupxA1D21R898zOBdJPpVYLzR0Cc
Ro7dHEtynvysZFFNfB6Y88RPTbhXRSThqSU70UgCngE0cEXfruBBkxqm8IaW3Hxh
TkUuQx1ZicR4YovfY/lq2pIflRsHKrp7IwViNhYhv1FFD1T1rwCxM3UWFxf4+aKP
wtz1QJjaCWSTqxkWK3artZjhvMXQKxMlmImO2ZbJPSxF8pibJT+EpE69Cz5bD/oE
8mkUW9gnE8l6nX5Ato4dvsWlAYGpkyokq4+TlYYQBLG8HOjGHACzXqnDdfEy5J4G
YwcOrE4YN8AfMeAJ8iHe7OMLAoTiWYTlKmtWP/QhjmUYK3lUZL3BUXvrAbtNK21x
g93SH5lU8fjS+17ST7a2QP/3d3QqU9V1j/tbbgeLPW/dj0U/vg70RrgqKQTO+t9F
F0RZl5mk2Uz/Rcbe/11zxxIZNW4Yri5cIXFkNnbAne48LK3v/CTgMAIJZDkj9jCA
kYsQ2WG2g7D+7NO9+TVVh8Y0CY5AXjbI9J/mb1lkUi7VVRI2o1NId/hPAJyo0DDP
eiCrVs1AqRNqifHCkrRtIfw2uS/irgYV0mT23SKtk1x4uGyILNezgWIDWpawjer4
2IEL2/zTjSApdfzwhvW6XmafBxuxej/ZnGfuBHk/U8s/nl9aMS95I37I7Eplrb2T
aY3m/6V89HfsOqRggf4EJYGS/ef7nQCnma9LQg/+UyO0Z7wE7HTyw2vhOsTcOEsk
IYWCZD6Q6VBXdbijQUJNKIQYCRy9tuk6jhBSKJ+CJy4Rh0K2Og6WvEXB41ph/r+v
9XGHKbhcoMa60tSSTNx4O2JBWm2V+WIiTGwWjZikeJXYB1CL0e0DJ/HlC4U6gloP
ADqqyKpsZT534ffmu71/CSLsadEIC0MDz+IK6HANfsaKtMEscyHEYNBHeRJ5/2OV
1ucyLnJBRm1CJpOtaxYo9l/CBCVLN1aVzFIkh5RP3worgBfa9G1qRITKpWaIDESW
4hUjNi05FiKSjwsFFM1WM5mDvIo5RxVKQs2R5DlJroZCjlywFIntPvMYm7r/6kNE
NWn5IojT7Hg8vzpuDy6C0YOjHPDo+4YpYAYT5wX2KXRu95SAF5LveicMTr+eSser
tobbvse9SxEi9fc2OZuVKCHL5ygRThVc8FfamFb+fSJcuh7DACkCCyjAkMVPao8u
r1iNaZOB10vswjK3NtnSiIGrmK7vYDRFISSEI36L7cnXmnwIFwIBxFu+JXyFXWxQ
gdQ3njPZ7mOI6f5II/ExCHXW1FK+OE82aqRFqd2932vve9jkts5k2GfZdNMpzE9j
oHNs5V3imh3ck/UDGJl1c97R3dfnBJRqeUrEqkZBgShDHv4mB490K0JQFajwrnHe
tzFhOsEOT/9jZe4klbX9A3PlKQLxzVbuFYyg8H7zvZyHTnfkim/YOttCW3VMrutc
k33tCjBa9pyzxG5jqMc3AkljkqxTvZdMzDEdJa247/jS4LnphEFH++S4/MUA95EY
b+gXlIXN5SJgXNbypnS0geb9lTZ1Xh+nN1g0p/rwZY0b/xhs9IbSGFOuy/OBHeTy
YOCUsjMOXk3yqujUC+WzkfjpN1zTq4ikMOkeavpq7BROOZC99PEQEX52KiE1tCRB
5mKvQYqtggsGYTpxPXCND78AKmnDw28knluvx+rw+u55Fjj8iBN2bkx0ca2wUZ2f
V3tx0+8owkpl+bSsc919Tlqxg0YMNg/VGg36Yw85ck9k8WDTtKr8XLJPBk7Qx0zk
dVPbL5WW2AbTEUGnndolqnt6VvXDuadyzMJxvncuxUSssVmhcMqECHQ3oH9U91Ol
mOtpOpy3FakeotoKm2tQSpaAdWpcO8QZqySisPnuN5Ll5JlHuhfD27NwysbeoYJl
Qyy6nHvugmb5IVx/DNXpreP/YIYCfEAsJ+kAcPIJ/E+DioJbmhQUO51JqnU0QdA6
Zqe3npTeJF00SUDsxJe5b0hEAeLqddlk+ZyCDImEaJ28RMHHdJoyLGXQ7nytzOtp
kZuzcjHR5hUL1oCxpgO5fnpsTEagTSK/jvLHjBEg6Fdbkc+XMMH4FsfuqRyBrErb
fbR8untDDCDmX418oYDa7jI1+4i5DBdXSwA9HYYANe9DUVm0wqkiGX/g7d/3G2va
V0/qoW9d9LsuPK6U/ESU82NXajhhNg41nBOz/OFSdAOp7Gy8gm04RFe89zn6CgrT
8ZcIpMENWsdEmwREOL9ozeGRsuDR8A+OTzUWrXTY6LTpBWRLsL2aj0slqv+0HX5N
tv913qkJ+y6H6/G1ZdogEghlBik7RSPnf74H+lhLYO81/81i3tCWcSAMtAe1qSnx
TASt6TvT+99MMtmi3TqZYD34vNYzjnqMiU4LRwi4CVFiQ+j8z1hYbNrCf9kovjMO
x34yc7fogIG5UVq0UtUyqxbZMC4B3IbeDqh2GoNCNNXzlGzZWcrQ9zH+Wahl7yec
Z030sGNHWWnltbnKd8eNDm8LQcLoA6TFyTZvPsWlu+GTXLQn6mzK1ioipJqHH4SL
btKGa4YlSYVlkq4rFKLCwlwI/fHte9AtNqZvkadX5QP1SkC5a8KO1nq9D4kEdve+
7hY5gESN81edzrtYnbF9h9fi4WMvtFbIIltMJnZ8cxKrUM5nSjE7Es5HV2+NXE7H
rwt7yTHhjyo9MZowBGP6G//mIWFaBxJcje44b8/jwg2zGv6iqqO7o+agGzAZSHjk
YmXfjLCI7O8qje2Rl7ShxDLcXWLTZAQ2Aelg/zoqagXLKP7bjAQ1wcsI/+9ii2Et
2QJAbB17OixGVYcNm1TLM7jtvXRI898e4vWIBDdBsXXptJTchSRsFCWy+DyfubY9
0HPGQdgg6FCJBuNnGRSRV7fYo0Wul8eY3CNP1KuJ0v57iz6GF58QT+4conqzsuTt
AdrDgkii7Xnl9/dW82XhbJIilZGEuNbX+gvcI5U2NW/fbgnrl6ZR5n7mOwfXJazp
VkcZ6+OzMRm0WVP+JjhRP6OdhWj/OtifHxhIYGzyvR969O5DXvFH7l97+hiK8gav
N4Kdd8uyss5ea66PYK7No5kbtD+1MiYANpXblr/r6lppY30taxqWhdWF/X7kM2RS
icoCDIe/JYbMWbObAbyTP5CV5NpwRIbm9jtpW9KLFAS/v3tPl/VCpUd15Dpt/yxA
89hmfYl7E1FmBt5wbXUwVVSB/yibsluL9ju3a8AEhKQOq8eVjI5qeQHZwbKf4u4Q
X1UbGgIF2npnpvRLM94NJ6Q5edg6hLe4hkqkN0chJ0tdL1JrLZJ9l8mrdci6W7cQ
TjFUCZXPYecEe80Lsk5N/xftYUzSM5NSF/xhxMzUoyCnLllIEe02nQy5ii0Sf4TU
bjTdmDX7LcDFYvC5cKxuZmtnzEl/879M6IQng4FSZ9QDp/YYD9Q5bgNnbEemkrUr
WJIvblT9FM/haTDxqURvrlWz7Zg5ckHFfB914y92dGOPyFYzE9ZlEXogZY9CdO77
z1wDbnFFl5k03HDkMfA2gniEN78gyjv2KfK09Cnm0D5RnwAIcSQSTKPecKldOrJ3
EptvrAJLi4nPDh7knjVFMWGA95V5+FI4qy9+0yTF3s4ZxJgxz1/kkstcMA33Q4yv
0ym4Fr2qEWtMIgwpPfEiWsJTZ8hm6Y30krZMbSn/YaZiKGi7MwinipzBJktYYYc9
cdhfXtD03S3NY4XetXqtmoXlJcuOV6cGyRrGEHe0WWeW0RdD+3gj/LkAsQIQQdnY
AiqkAu3RceHm6ZyLhUFfuXsVX2v7PDZni2tDPhI30MkRYknHiClZY7q8HA6/pk6L
CfGYn+0fAQyQjvZ2Y0ss8vhht+2zzxu9zoMHGOIZ7+XRv18BTq1LXvQaBDM3ml4z
+wi7i2oxSqY00fTtmYZynI0Pz2wVbyfQosRkU6G567zdwFvth9GH1+ggMg+uKAmh
+U05UyZL9MJDIB7nC5Ud8WRrAfaRuqIrxLM+IvCc93ePFGsY2e0mebkkYjCdj+iw
S6KxCJl3dhy4PA2WlBIqEyNi42YYAcqGV9oaiM807kb9KyiI8ogRpab1K2h4bof2
YFuEWoGEYFLUhslUTHTdiLd9RmgZLR9Tfx09ICRwOm1MDp3/IVbTYUFzbdI0ivPJ
GvfpaM6SUsnPgO42s3SQtf/QGkbyvV1IpD5/wwbMbV9mmBkp1VX8wuNPpP0an7fF
XEXP6XG16DJ5h+CVxnFilDs8Btr0LN+Nn0SQXb55GmnqyjDTINqKd0QSCpkiE/uT
3V6PS1mG5d7Lp/YQ0HH6yZzBjBltRlR2Xshw3o8Zo4V9Hl0Yjq+H1QQ6WoFKk6Aj
I86AP8Rla6ghzOhRrhen55EbxWIRmhQC1zDAGUKQiM4i9babtZvQtq2K4/57v0n1
Lh85obAa7BlFPmcEMCjvMnt05V85BTozJQjoEkLlUIahfrtucf3B5dcxS8ZObh+v
f1OhSC7J6r+8OQ6IgW04HSOLvnvZNcO5MtXednY0sudI9edrqdbhAVHzEufzia+A
irYW2A9H2c2/jBdMD8XKRKnQuqrufsgbCGwtoJTMKpI0SulEmDO19CB+rKTs0ySC
F7DiLf/AGEwEvDrkFpfe81sFN73Oyv46aw/sNuSQJjJI6/mny5uB63/X4VqDTMot
M2bjMV531BLAb78khRsM396k5JkTN28Bpo5vldx89kqBGzN8ahaoIx/FmypOSUFE
ghHqlXsXQa660OO62tyokl/WCRE2L2YtoyZ8CHrItNYYQC8nyx+NZnh+n3F0mNvp
VCIT8V17wbmVkoxBGcyJAX22m36oHJIE22BSixZIHTxAQy/jh6Bb18aVoZOYAq8v
jDeCK3+1LKbAnUgYmbuxQ+Ane+puxm/pDFj8o/lf6bganeVviWdviRYrNiJJlHiu
0lJ1Z8hojKbkQui2GlPvbTf1xNtfFoU4OveqGfAJwdbyF+xffoksgeAXCvCq/pKw
S4WG6FILiEoN62T2QJLHT6GYMHUyCtzA7hfQzsf8jhPbpupcI+tud7/LaPCsXUWO
K4zKGCazNfxsAg5Ek6AKWE+8rPFFu94ngN0+rPCes0Yw4me3F2FRWW5S0h5olLx1
liXFzoU8n9nLWWENJoTxsuYiHkrQAMgcl20GV69gKlly4DIOhCb6djsUUs4b9hUR
RDXdJ1jZdV4q92GV911o5LlkweOPn0xGSdaOSxxOEmwQu/e6FDo847F2dgwIuz3o
CculLk2QKVFUNOeP8iwsFQrJggoXf2ng4oqVDKYaZdkURNTk1judE+2HaVsv3ftq
wa0+LeP3aGGfo7FEH7xCmFVUC8eZNcSTQVPGSLmQShpi6sE0q2pTeSHrUN0OBz7d
vTR2wXuOq5m/FlWyunjf5QXcTmbEmGu3FdA6DoPBcWnUnYl5zaEtkGr8CIEp/5rS
+SzNd7Prirp/8WAkc+Dpwc9c8jte+gN6zv/NFR37X9NFg/IcNFC2no1ljYIU/UjQ
Tt3iGveMrvk2C+AUko+s9m3uVixDgiOA5YlNr1FEk6sbYswaxnOAqHrchXL/HQO0
au61GFq+8fjSVLEqoE7ION/Ektx+clkCy4jF3un519YE9aTvrWmgQfRZJ9wJMzWJ
BXTjxDyXKf9JiqRFKFhCTbRhzUo/KUDKLIQOcV2QwhQlnnu5Jm9o9FECGYh6unWm
kVlKahI6au7387AKDnDDdfa4EeDRLlwKTRiNfM+6VgdGSKY8NJewGDaoax4knfSa
8bbIP1iHX4YeRMr9XjWMTYWi6pelXNOGq8Z3+R9kdAtUqznu+NRR0IfdYTO+8Zuu
JT9P+yqSLe9UdwLMIgJLpjDVpeJ9lsRv4zJHk1mRRB3t7IfufOSFyg1FSlCL92+K
OKaY1VfqFcgLeBfyNsZFi/lyoDtKmRCpmRRd147iGUdHPcdksuTvwRPlXImfp+Oz
BlWBfs1EqenldU4vtm7ryJi4++UvvFxTb4YlxdF7h3XlqWESJ+zLwkZHPZT+GsRV
ECP/exbsyYPoSSOiuWM2nqAm5ed8RiqPIzS/EcWUUuJUgjACkyp9N2jO5CtUMd8D
7H/ELNX5jVZEbQrJRu0g7NbixyN2W3uCEWOwoUqlIGFCicNroIbp2eusD2doSxMe
JorJ7ryhjJwihBRpMmtdY3P6V6u0epQsbvSl18l/AdO4Evcs7lWBs/8cY1NZ9JvF
wqJki7YCIUFImsK64TyXCI5l2lZjMxTAiuBeEEN4qjXskpd3ImTpg/V2gLMgfPEp
A6rZdlg7zSNzps1sl3CJRoS3AWmerNNjb23EEtnz4IqIZQPTxfY/laEZjaPy1WTC
LnclhkvCdPGx4U5Gykvb35FZ/5foCu8jbxLZuP4E59jREP7YDe42i/039BMbDLus
o5EjKjdnJcQ+/nHywcFTLB4xC3S5XdBlgoNlc+rCF+xq14tbwJgBe3mYjIqnIJEU
CBm6vf0AzM8gtWLY/UWXNBqFWYvOSZhm+7b2TkDC6tkPy5WqD1Q9JBiC9hqZka/g
7jsmBWdHVF5guw7xszz6AA/5/eUJ+hzBpO+f9FzKu69kloWaRgKYXoCsoUOd1vPr
hTjVSdCRqPn2kvpcDCJG5kAkSRKpT8XkEKyJEDGYNAYbg+RVWYgck7NuXRX7cOG+
vdlFfWLtyk5lI19fAmhrtxVqUal6c9fLWHLZy3IL4yOS15Y5Va1i2rwLYYuEIUDX
ktDT6Y5i8NOaoDaodK9+XqfwauNS0CGUXShHHoNhW1p3R2nOqe06V+WFEcAuk1oW
xuwED9qXsEaKKAw2LJvH6HDYMNjzMfEK8DG8Sn05iTIvE1owo6Y5UtcLOlutbRch
4ST8O1nCrr8djEjgZoVPGBJFYCkD5sSw7655uO3AsAHKN/XV2SmlEBAVs6JDTboA
Kh+yWXH2TwrgPmhH7QPIHRkBPZIOf4+S9AlPRxIuuT5aBX5R5daquKTxpNYvC7X4
mI0EUSecBQAJYVV4s+iK8i2Bo8awaFVTYoUp396/QSBNJAfrhixIf1BRUQiaXJ1j
pVzyhth3zKXt+juqrXipd3a17aL5X1gmtdkKBZ8VGQHJrSQpv8aOQINGYGMJV0Wt
fO3gOiz3XGcORTy3kqd8WNyVikw9iR4cZt550jpLnhmdBLXmlb81rzqMRFm5+lQf
ZUhppJv9BUWbSJjy53UrVsnrZgTXBq+xlaLpiTDK6WLCatRGz8o908IU1Vxpk998
lqv0d2KjCGQALlnHb05Ft4HnDtpGVzu/N5ZiIjsLysaLM3yjJwaZwO6wy+uf/rVD
8ppUSNIrgD/PqeqX3BiDpc40BFFyngQn8MOQ/T/jiyU04HaREUfmw3apv5vgw/Py
R/4lk1DlcW8wFiINvnrP4F89xEuesgfpdbH6CgxummjNVdk1l1mDhqhloh3rmb2q
mKril+jTSlaxMoZ9BTxnmILHOoWRsssbKdTFB6Plgjzvrr9+EbAl38ESmqCHoVlD
QX1M5Xvj4UWb+f8iMS9TFBLQMCcQ3NxsyYpsRTD0I0S+XJaxuxk8wimC20lEH1Wj
1JvTl7wjtyl/5+081fY2Pb3fpupnY6A8Bjwuw2IRbI2Rnt6JP1o/1k2fcnzh5crb
q2i45os/Jq+djspXkuMamO29GHf24ZcmQAlpOMRJZqLNL0aaQUrRAKkPAlrF+SrS
62L+Q4opbOiAV6toeeeOsXSICB3h23GR381jLW6Rm0NN7Vavm9FNpK9SWynImFzh
1S6oo979umgDoOUzwQd3PinmgqLl+9TFVDc0ChOV0H7Ot0oKc9gER9Q+0mnNMcMt
btVgfXNtIEYP98anOxhM8ikQ+TCXByrDpyLWYYl/K3q6eGt8IFskaTweBQvPw6kF
JdIy1RGCQOHx7qd0GWyZwbq9j/dXcSRLJ0fEGwNZplIbuzgMpnMfXHxLBkXxUid5
Z3vFnoA8+LlU/nWROhZ8RkEnaDreC6tVDjCl8V5+pmycO1483+F3P5+FbNCrvgwj
53r5VuDyQzNaicHDEueegt0k026HuhDepVIHDrMaSudQZ+vzWuIT4l51LyjQL/2K
etgxDtB30gcU0K6eRgigODW5yJ2SbsnJH2Vc4glebWwJcUxA/B5hwhaDFHTrzbaj
gDXsH35Q0NUsINKAiEb8JVrcPyEbVRtku8PEhbEKSmT6vtksfv9ZSf4hyXxPTMFz
CtAzwH0FkvEhbT0AgY29TtfaoK7JvbXLxtB4L/r0mw+u/xB2i7E3O00Vqm3/6tGD
Tuj7MEjhd5hqAAnh2raeXYhcuRUAHjp8WnJVJbIy98xON2Hw4NebG2+WJsO/0e7y
dZ24wOhYWXtx8jHYkiTCrHcmzTBxVnb++2xfOldBjZQvGxgCpYN5Rw0Wuy0OGCpR
DjKFVuF+dIchh+uQvYKOAumKNyYrOw5jhELj3BEIejaUpwG5pnYPvN2bDaSK4Ahw
czH7ZtPybJY5AFVz6oeqFbW6AxM+zAeWhSQAy9nQwHLLgTPxDhShzqD1uectW7Wi
9nmJJ5WMZajgUnxciAw/1wg9e8IhtC8YQufeA+ldPwNIG1z26k6euTUvB+8rvEXK
jZRq++aWtd1fI6HsD93YKjObJBVX2dWbuGev7/2qN/t6wlB7jx42MiqKvIw4neG4
ONkRyh4F1Yd7J7qlPez9++LWjRp47psRE+WSIUrr0JdH5Jw+mLR4H9ETJ05k70YS
1yJGkx9VxAtoX/oMJT0DFvNYbOz3aPOLV82vM0jFpa+KXkUTWOnmk5dxdADm4q4z
HaJr/tSBtcVotHkpTd2yxWHcIwaOzJZJCWWZONHV1/KHyzkcALZwlkalYBiu1QIQ
fi3OnbiTGnbJbrJ5QupFrEt1Qr3oi54rOBVQ80UuLjXMxdSqYqdDz4X39BVYM52Q
j9Vcxa+EYBTTtpmx6mbzMugM+9XU25K//lnCQ6Vc4BNrGpnfgzXTP4q+09iw8ExZ
2b0pTmTcddxS9cKSPr8O7Hz1vrQE+nQxP8zgDoA7xIS+Q0y3My0u0pw5gTIwhjyj
VV07FNa1a4W1Z5aP96bQjz/V9WSdvpBAQM73DZd4nMrY4IyGOYj14AU8LmQLnBW4
AINutZ95Jw6o9nY8WUKGxmHS7lzCrk+iGuAG80l10yRZ7CEhoTYKvuLxaLXpJ5ST
la1fJH21ihPiS1YlpeaqsWnA4NNDdU3WqHhAPazIsmS7nejkJR+0VWgF/wazWSa2
DbMISu4CmS2XRv7US/jhgNmHvcOmjmLjbc/sO6GhN+CgP+DnOaY4v0END6qmLbQL
ch3Han7n23W8Tr4NrB4rJOKtS0rLrB/3kClwvg9pc8T+laaeKqBKJXMNSIJSda13
wNHz+BWrZs6eBa8PaFAz2SFChmJycXPeWvWopmb9EcB+jGjWFUq2hHybE9PelWsv
g1JQZA/+hdvre6BnGm9QiZfz+w2DeUH2ZyJfZc5qZl6nuJY/5+VBYAe9NLFL6OyZ
nR1E0vwmyKGMQllnioCUiwTUG7ij+OQJ/gBkBiy3c+fhBiDoxeMHk3nnhQ8FH9tj
st8DGystE2JiEuthUqG1vtilN66s106oXBTMWGf8CKdFUP0ziupTrjNP+m5Ablxv
ZBaB8cS/Ab1Fsw3zu6gucE6GP0PODKa5KNZqUQ7bFt5mI3IfzRbqpR5O14hBWMd0
lco4zoPmK8n7nfcR59ltz6KLmqjFl8PeZ4iltTC0riTxv+QisbIn9R1RnNWthB78
nqQSZ5rfSA19GOUy30iXmJ01VAD+yCVdMSiAY+TekqREodFTMMRbudud2zkn2wvK
fyHgxXqn2FMwVvfCR7pgpUqxd1vNZzu1HSL7U77sl/QSiVKWlNf92pwXXOg7Dfd7
JvRZNJMflNB2RATB4ym03AuFPv+EA0kORjrAiTb+W0xTS0TYFpEk0aqObiHV9pli
AaAynd+kkpmiYfbro/Krt+7gYsPAO12s3NlpeUL+XA5KE4k0A/0iikEbxfQA0Cgd
wHGmY3LwLMj6AYZeT6N3c76/pe0tnMntUG6VptO9CEqsUWd6xCCOCD5S4QGOa6zZ
dp83pM7F6XF5mau4HOtQfhZyGZsmPm2IaENFLdLQ3r62tJKlK8vVSwanDqqCkTCW
8puZTkDbgmX+xxZAONmPZK4e5Dw6X1im338bjJhGSyZ41XKpxE338fVu2muXjeY8
gobSLTkJ199ItEEJvd1ScSXWkNH78Lc+c3dCbe3eyYJ9o35SBOS8jEtywgW8E8eT
hHbLAc0/h3xZaHJrv5go5u4jW0cz1Q/4xJ0m2GtfEE+guWvORnB9aZ9C6QiouEo7
gqt/MtPfHuZl7+0lW1RQH9zpwQxefCYP2vvjUsAtXfDvJXu8Z38oFd48WFHZTLjw
wz+cCYo7AaZw22gsSEmnzpLWCF3lMWsm1Br7qD8hHt4wJS75TkLxAWa+jdIU/JQ4
ivaed2kqfG6HOwOW7P8HryshBIKh0AJ0AK9IHxGX8rSOqnuCGN8MWoMBqtsnIYh4
Z6cToV/z4PAg1xSgp65vBOxVEWpAl7F5oC+qyB8dTrUBAk1jmStdayNb5/GyAPL1
x3RsuLk6cpRmmbYxpC2Dn3aoAC/LP9VkEbiHHCdGF2gattCjqoBruS57n0Gcmnbs
36Dx6SSMSrIIuM6Ad2AEykNdbYJyHnp+pNvMqa6Ab1th3I0NpK0lqm/bBcO4zEgs
uocfrxAZ1RGgZ6rBGPdSsKwqJjxakPJcAxmOsripWGtZQCJrUdsgSCvKx1cZfSo2
so5P+Awk9vGMx26NLmNC1wlVzufYIe/YAjlRiSsui6nF6JhVHmO61AacSOGSvq0m
btTQZI+Xz7NlRaO4Qlo1RMdEvRPCLjmd44FhmYrec+lcTPpzfsq/V64cTjlfjbMP
cObSvtzB84mk/rrNBXHG0iTI7FMfo8E8WMQqy2pF+FxXF625gKDmn51C67qJoTRj
WpwiTqs3OVGG/Xzdy2/+OMMKZyu18zG7mJ0v8ne+9gd6hNprNkFp0rx+RdqcVUUX
GGHx8T+MwXDFAg30cGE4Bv7+IRdOAI3mvQubFXDtNtP2F7pb9CoCB6g0FU0T9mK0
qbf3hGr49Y/motnGm1/HsChJTDIbqGz8I1WyMs+1K7LQ94na0Pgc/XTRHyyId+xz
dVBqgmsSxB1Lla1zZud3pFnSnl2s6OoNoSg5sgHqtKAec+QwHQQfqYdWLqPl2XGS
FGNqAmaYv+Fj6eR67+ihrUqd6oF4GovDk1gLvZkSr50vsIfvFAuFC+N+F3F9qcvs
xSshJpZyGDgBufJXzyz1eGzalTmb11/oVX3KNcZYis5RceiWnNLf/g4rcE3Cvpql
G0fOcPQPq6bEQ8t4wd8wTHSxn95hub1R4zaCPTBmm0XAq0l/Mpf/1KPkrzqA3J7h
kdJ6yIupAX1s67kEpw3UIKXXZLOdjHJKusvQLyj/njLEqra1o29tQ5p6a2dYBuyH
v5ASGckkvcU8MUQ5Jn0tfsQ1BYhI0aEnDBshWS7C1XFhk0v2bLftOEX7Qw1vasV8
5rieJAfIEa5sCrrP22jPO1/IsypNeAqwkkMJhWODM/SjkDLD49b4kwUCfbhDu+3S
+tE0I7evPKDN4cR/vv/aX1xSpYDhq9jkqDMQpkuNntbESD1mVHAXXnT8yQsvdPnE
HQ1VOFnPEH2DUnxCYV/EYztE1ERnwpR56crEUfOu1XMaEVwfz9KtSvpZW08uU1vH
iYb1uGRCRCJTO9EhxkRsnr7gnp/SLghbfLsP7O3gdBeLpvFjMO8YtSKNfWNri8Ie
69+udIN9K5wdsvZGOXnNHOuxZwHbwQW1slEQxIYCB1MYyw+Xtet7vnjjTZHtDuHS
TsGzu3KFqy+N8JS/X6vOFsajrqGMiouNNN8XG+31yfqKq6KTsQsIYWnWpsYOtawJ
6yp0lrP4jj9lTJGtQTzThq3GdaotwJibcw5ELm/7JwTl3VnZVQr2rrucs78+RaED
htzidO9TPfm7rKPU0INFctBEfdXM81rEmB4EPP4AYRsZcvPW/9RZKQvxJoqfq4Y9
S6y9tiZnS07GYHBdXt/kgnGKFsT1AsKsgeEEXCsQT+AP9GkJ4l2JvGD3kmdAuGKe
uWvEhjTk/tn7sVqNeOUjKCc+tHnVEdVblkTavPEq5FTFB5pcclrTRWsy/okE9V90
FIQKvVPWZinwa3HC+1PsSb9pH3yxsHsn/FtkLxGo+p10B0qc/HFukmq9Nrv0N5vL
MOUJJnWknTG/FS09jxP6qex/x3KYlm6k1SuCjoUObpx7ig31Cu2i6iNpoh5Xx54W
DrdmbfG2lOe/vogW0/pWVnICzI5Ly+zL8ARx38EuB7/Cppki+IEUq+jywQ4tj9O9
qKrwMqcogRsbDZUWEmcVxPtoxxqyB78C5ZguKAQKmuv97bt1mDP0VjidokdhDPO3
C/15FQU62gna+S7BqSipltF1dmkQxiAW8Rnr6rI+XFzxctwuewgzZHmhaQsW+esh
yMMklHjvNCXId7+8y9fH3uGeq/GM5f6PgFJsS9w5S7teIQvXP3B5gHyb3Pc6nk78
/Qv4zu1FK9sKI3afzJH2Jy//8Sf/SgQ5EmyBd3ZSaRqy6hXBVqncgyYBsetsAle+
S3hLHCODHUgCHOJpDSnhgWzwOcL2qE7FCKqaol4h1KC/XDqQSzRcyxWRWjSHfL+A
0sgLBCZHmpbUPrhq0VsIA491phlBWXUJY8DeJXj+f2IzxYROGP9pBmNtHyZIv1Gm
1Kc36F9FZsEA1kq+J22UcgtItlzaaC6+yEeuvbaRdSaWHsp2GYpO2yr1515tm8dU
3VajIR/DE1dIlYC9IZs+4fwpgiTqB/1I8zY0FpaG385Dc+2uedL2z/lYfHiTDJOL
QZXZpJkLGwD1dB2gNYyxNoj8crZWHpzH2FCNRHhdzdHvieEAq+FwwuRe827r6wSR
02YQLZjBqc9ggVK/CJNbRTdrH07rSvaPHxkX5DDDeWqmNpvydfpS/58uYO4CQcI+
oXpsDnUJlOKaiV4y2jCnolmI/BhAKc8jIF9oQTaO3aLz3BqisU9K1jUKCui2Ab71
xPfkRV5QpzKyzSYOwoR+F2wNeaej3kozGdWtc+yBkq9IScSbUfXTZf2i7lU1BbVv
UteqI3ahs7FhyT/2UpVRrbaxgNzdD3dIyxIngs36joTpKvJY8caZkGgqRnzG9LDb
WPr64dJRnNGfeKfBxBO4ZYNAPzuzfAyhuEXSChHeuFMVidZ3jYMU8k90UtO1RbJN
xsERTIfpJRDaBUwxVaXzghjzmxgbst+ZMhAp9zTsT86gsV2HfO+1CxFoDMFk4pFe
1TtFE4AcNMoto195VFJ5K33t6cIli0A/AIWq0HJq4Ok94U0/S0DIOEI7B/URfRLE
57XLSYMG2W8MCWfejRdhPfP2/hUKGQr5NicNbR6foYYb8YEttadmuI0k2WhtpVUp
pjKNRBbtABJlQ/D9dPAyvCaNJqq1uGa2oOW4DGMzuMXx+CueFB76yx9AjdpqT8xU
9O8BD5u8cvLorAlE5Uo8ixQEsv2z/Nwrt7Y4+XmskDxRyZ88oFZOjoXPZuiXg1Y6
xla8ZqwnLKZ8nnBSYr8cGilNHAjRMzJzeDsBLbXqHC4zQWUIhEtHvubW+xKi97IO
3qGzcN/dFxbP0XGYXnjGGZPxhQH/clOHiKV1+3lVgK4RY5fzQ0RHFjP6YWBb2f5l
YguOdtVXhst1GN3FynWg3FIJHYRUSd7OKyEFloK0Nwiz1DVneKyX8u2gSu/br9AW
mxkxD+GVWfnsxH/PvlxMeBKHAK4Ut3SN84fReHK+nUL/EW7M8jb2Gow/yuAoyi5s
sDcTozkcbl7UV2rAFqQjmOSpLq8b+kJHc9bOY3Rc2GXGS6cMwiSWO5aBBwoC87qY
9pc6hlmSqq77L1uXhOjXP3a+pMncaBWm6B/x0yLbGk+AjLccjdMxVnaUzWGUHDJP
IMG8oUh+2qMDp/ouANSGAgPiXhSG/GBmLmAGqk94JYj5AEAmw1st50xVxikX0G1r
L+z0DVU54+dkn46qWck3ALAX6miSy87isah6KjJHKHE0Bh32i4gxb7XlaUNEnP9A
mQ3I2T6vEYrbpNJ2+7OI1sdZ/+yGBobFI+bgAuaQAVadB7tJQjHy4V7IOzKq35m2
W6e9pAABaW13FC1VMrJ3Ek5nuyKbeKcjiHsOMSZMdDV6qDCVb98EdaYqpW8vd0Cr
DYudSwBxfa46KOO/xHabFgylOJEs/qBL+DekN4bqp7GRXATGlutWdZCGG+Fjwrmb
DFW1uwEzMVzDeY+TLgR0NDf1oxWZtrPAzC2Vdd3dX3n2qfw0jA79Kpnj+Cvx7HD0
fG0VZnYJqHwM2Bfxqmp94Wr9blrIHsFRZ5ZpIbK/ClJEN1YBJbtmNagIMr4gdz86
YmymXYU2qFfph9XtDdNI+ZkZx2zUoiCMCi1RYdMDUfHfI5nmyLI195Va3bFDcEps
QU/Ra/3/Klvhxp6UMcQ+jNAlyyc6SoUz99nkYO87B2a8Jf8Ij8+nqy3udxN0acdu
dpW9bQENu6c/QxqjC/83TGZdNq5ONkRmEdTO/4x1ipm7At6eVQUL81RHBPH8VS03
cs6wsJ4Eo68Xry+Qor5p53NupgDivVi3BVKggcN60DjRbTw3au3cumn3YUNYyyk4
TSLUjIgSbWmgIyUVlPbf2iX9Jgq9CPUp2+d4jKj/TrgpGf747j+eHrsdmLqPsQw7
/gj5DJqNKYpD+ykGic+T2b+evaQckoWczHQe94OkjnFfp2Hz/fJqOG211Ui5/NyN
gRssZoleTfxXcx6/TmMBuwsRfVC3hAFWjtCE1wqL8hKyWFo69fV5Y+D34I/MoT0b
rU6XugnWlU9yPC/yruUz7Zxrp/kzCOhNIikA9OhtW/aIb1rZ/8/oCooBT0PvbI5M
YmOpLeLVMZSCRt/r5CKALMJDMgTdKDly9JxSuffy/qkXITEpa61Q9sUh4EdvmKy5
a0S1YEuKobqthSC+F6Y5XVcwShIVbjKc40bDOsLqJvhmf/Yr8o6gCq4b+9KiLg2R
I/id42ohhkJ9Epc/nDX6K6jhLdei/16NnCE24SNisHXCeyOYe7LfmO4WkpCdxccM
A58+rI4vnTN+vMxEedDNbP0rOgYIQPJFrWmkuQfYcEHSDZfaeO3sENfeLDNhq3te
ZdHlqSDMfj4yL1m38Jfo2Z6Q9PSYjBmgM2fjRg4vfXGHLtP+3uxFiayLqJ1U6/wY
wC2uvhZoB9XFlAgzQX6l4iH9jvi2/3ytlK70lP/KqQwGyX72cAo8ICPqCAhXfTfG
Jsm3wo1nCYBCA21GGKcgk/k9NvNA8/pcUjA4+efOOd73jwZT7iz7QJfyVy9pMU0K
y5w2TNjoxPsu/bGoguI8U/fIwCIRnCsGrGdxvoBpThvobsMD4WjAYF2wgsv6KUdO
shk6yzk1PDvzafsS56UcnOHrn3qGmHU/0kowAPQDoK8smVfYJmEAb1vl0aY/rrLe
L1jidiiGt5+zB8t8Ja60mwFdjM0e6C8fS30rYQQ4o4Q+5QhlJnWEohMEOhPtUcHs
pTaL5LCSK9FYJp3J2W9ZuCf0FwHuAa6YiVjshKEN+3+2kdAfyqSUZfzyqh3V0gur
sal46JPDQWrBYCKZRvy400CYtALld26Brc4WNTKptW3SRWN3Oac+V+/ZhlDvqhvu
2Lw2ngGybWr4P/8My/lwqCZFDC2LPOUwL7f7ykQmeDEQAvMnRv5MOK+dnxP2NkkH
vX1kA5RZBeVJJAdm+aJWVRph1D+oRY9LnRrvwxuHhbRxxiG+m6T2lJ1R+cfFf9Kc
oKQgUk89j2SG54mJPkxCU1gF2Ww2S+/zeKVVuHPSneJvQ7xs6lTxh9pco6iw4Bhn
IAA/HEE7PYwEtITQ6ms51ayN9vu2tU4HkU7QjLXeN7K7Tz4Kp8i67ete1IQciwZC
X9CaGvDBhLBfq09faPHBgMP0DV2tHu9ZBi6bMivSQbYm4TR3SS8W+jFscbfeuhIb
Yla1JnUn07YlC3o3m5eKEGi/PQ/CCdXJ4QX4x1Y3yRJFizDi7WF15iV8IOUXwS+8
eCH/8JwokrkpbExJH9x3LRzWUSiei9OcEVUPQZrRQkKmGUZAe6rqy1kfAeLeDnH5
xS+D89v6o0i2H7jdzYTnTqF2lsZb9qTM4xKIl68fySB8pKMM04yeBf4MbvBBFhhU
lT4+mNfOVrKen5dTMrywWngGng4E+rqSaqW5purhWUnEZf4YAmc+I7Q7F2XGKz58
1Nkva0qiuSGwKSGXMpnF3HQnmftD+7bK4pvBG+PasNB7bH2OsA/IDoYKGCOykrRC
lqtoZVeCjn0n5KeG8J0PAL8v07JHmMUK16C7kJffswQT5Eb7msqg97yZjtxpLihU
aFEC7uuCEzOPcXEkM7k8YKL30o90j0S0s/Xua1iYUljax3zyKPQMQWc/Psh8Su3Y
nFun5Tj2uz03JDy7p5VZ/b+8ZhFnvO+GOV/5a/kjafdJLCCAwWGkuwi386A5Zw52
KfNnDyr6hvvg4ZuwDDRiS/eBuE+QluS1GxmuwUaW3Zi6oEWVEKlA3iPtSOf2ZSVQ
dmYzDoaokaauoYNJfMajMf0yFdTuQaDgJB0ycI8cEVsw6m04bjYEzUXKeNiDPbVO
wG82wpfirOaZibdHxBG56w7ZG5DkiqFHuzT/AdD+Dt8JHosz8osHYS9BRBraC2C5
M2164yOUmkJUnz+aKzHOxfaEH0DfBHwpQtAnMzdLH0U7dLShb54lFQx3ocz3Nh9r
6Yo4viM4mT7W7Nhhrk1LyMZaGFDKLW1piywBj5Cpxrg+DLqQmgr1u2Kd54pH5RD8
+bI/LhLrCjOuiYRtzn7G0sQD2UxX/OCKJy9Z635eb/Cw3UT15FJwJcHqWISV+PTg
zR5B6ZlHp0Zy7yb7kUxK8F6O64mHm4ADdwhRkogqHOiaN0xDXtlfDxRhPJGSfHOO
IQZ8RRepRFi+rS5mP2KPi94mzTPAfem/Mx6l5Xsd5fsmRU08FlE3Gyu5ONsyTybK
tWKjBm4Z1NP5xLEJYV7GRiezwSzRMCK6naawYb0SMgWIohdk9u4LGJj5EkIhgX9u
5eItXa3eFApC+ThJtB/FNSJEw3PSEtCNilybNwwUSH05cjOrwoCe2dezchWUYZ81
PHnv+xf3Dqrm+ZVpEw4LiI2HSyxgTgw6XHwiK7ozkS9bx3Tl4D0joxPER3brXdRs
fbPLHDFFYaoZqmP8EusJPTc7GhugOQJNDwA6Dnn3vwIC8lHD/rrYp2MHMH0oN+GT
hmbEf/3W6VuCwJpa1yKH6m/3VU/lIOXscqgLiKZ66tkTJdlDNRHC38GCeTKg8eVL
VN3UHaJo+C3fsYMYOhOSbBH/9QNdo6jaw8/d96S9AmnOASrnN3mF8LEyPQ8mnQM1
cYSj5ri/nlaYNbjoPiBvZhca0pf+iZyEqda1hu++5t0Y51YBmHfiU4FrNMTBSfM7
wMPalOoSfV1GsfrAiWTlVe7NasAhLHd+PdtDfJOr7+KX1TvnLNRdzv2kkFujE08h
GmZZ/3M7HTtkMaYLUBgWaLMgC6KXkiinulTIVYDz+SaRzRTd/i9zC0CATA2n3cQE
wiJQ2b5vDZxC6oo4eEXzXS8bkAh7qFgdDe41fz8zfyWxxOsh+Q2LsvXcrwT3viCU
EP+ndoJtK+fUPpzvOiUBN6GVt1QPyFufOgLkwWmMJzRikTcfhmkBSR1vGIfKbY4t
CK+AWE26PxdjghGOt03yy8h13ff2eLZnCpPgGsLW9f7Mr2tNmbMNhOm0v3j1BIlj
6kNK4gpt4dhmOxVcJ+Vb2QmppNuK7s922gG8RV44cHrbeZNzW3SBDVl7ubnZo2Q9
gjMin2JOxXv75zaBdA2IWCLfviWIPqatmhO1oDJUAmcdgdw1YSioZhCMLfh/xUsk
6Oy495WHBSQjp1Y5/m6HRuQ6xYXWeJrFwIXgp1DqGBH02wz8gYLHdF5r0OptpASB
vgq18Bori3Y/PFxi8Rd93FIifoxRQ+tkaEVLuIb6cbFC+uvIKaP/q/vlCIDv1mIl
+i/fD+3DsSBLeQgwRqPKxLORRw4ltYycp6SOkkNMIGkC/bhkq0n2SItL5V1ijk8M
a7WakK84Hn2SHYwZEPSOcRxHCDtgoi/hRIy1oRLA2+ef5g4G1U0WzbatBt/svI0I
UbLXBZg4meQsn6x76WMUbpT6/taGChoEy9AvH4TlCpzYtW8Lq2LS6B6vPb7VIyRz
pbb9R9qjqLnSLUgUwUbwkduGL10hSCXCXt67+eC7JDtv0fLJwlQxOtSapOy83HKf
mSSrWKy/PrzjEAXrTAZ5hpCQqvRo6BG7xMeZeonGO3q8wOdyaCzQm06jec+MQNas
eRz+GmfFF0UK7TiidcSrdOXjdArBLB/wwRFUwt6Fdo2vuJ4B7aMH0FEZzPGRlfrP
EDxS4aCN9zHoewJM2D4PbleGs6Rmqu0KF4KsEPf73HLPFS5jre+tRFdG2tgZl0HY
gp5i4NTcLYw5Sv+fusjSeODlTRqXeMG5EQo1iwjIelO6b9nv4YUo5DP4QkyESuU9
M9PFvx6dvc/A51gSinlVNh5exLZW8S1rbbm6PLTkBO9UU/8Gp180BYcJpQQOjsVJ
BC1cS2WIlpfuutm7wf0zCCNXvMixBhqyezkwvEAiVQs+C1iBI/5ZOHbIIIWpPkGj
svubJHYZFZy+FFX3mt66njYgk4jfBTR+b8Iy3gocgH9ElnD2bMOmC+S6RTRIAvDX
LrLBLz6TfEon7hH56nvrnbq+nfvvbGnp/OKclSwBULXNidOzVW0yBL6ds/3lqQAM
w71J6UHjsTve5ztT36ml1LOk7DJhNcZKuc6oHUx7z7fXLmn3y2AHbpD1Itr0Wb4y
BgIH6m/IaTLN7j0aU9mBp9X4jKywM2Qdk4Zkxyh9dOmyVJ7Ub0awd+vO4RMvjaaU
hvCMGHQPcLGfFPexjUavAMzmNhNpTKf3dWEh5k0h+HCj0TFrW57VKBj02iJwtv5q
IP1coUQ0RmGiyHZehoNkJOH21HiWqbwpCGWxQ/ZLd1yPPBJiK0HlTWljeqaBCge9
DpFok49ohUHHCj02ObaEtwV04oFtaMfwhklwK+zcPPOeTbKQOH6FOJNiHDIXRpaG
pnAG7ufUPa2GYlfnDZnQV2g/YxChTdN3NX6899TiQDBdYMZgDydDY5RIx5dg5sJn
XmOU7xoYf3OFXG084bqZP+vx6nD9Z7fiPhunJnTehEcACUvlBFpHQgS3oK+lwpLP
8EMzDXe6/aW33cADSEJbsM14pfsSjz8PLB4oJ9gnj0Qyh7pLrCg1ZS3ULrRk6daR
3+Jd2WXfHzeJN+HedCIK0L2NoBi3NWksaSa1GXXBVfCgWVjdyWaBBSH8sLEtl6Pk
S0WhsjPbzLi1+nY9Of5dPJ9Yfsgtls2wAW9IoJm3peavSbdPZEyYTw//kPsOBDCa
vZOxH3sL1P7hwkJaUM79AIdS9nVNFGtVDKv+4mtrsviUMSH8M4hvngX52261jjlc
lpMITlmrRlmncCLNF5m065ggZ3sCROdiEHnfQehzfcF15KiUBvHOLpIhUwYV8/QV
n5ohCztYQoBwRM6IEqlmzhNOPHJsSmEvnB8vhAVPzLNyXzUuk3WcdgaCuGR24dQf
JEcFRDBFz09cChkHyR4HPZxGiWKB1s0Ff2OzZ4Re37jhlQoG6ECOn1V8XNtseFCa
Apc41Ahcco69PtQlGgOSi6gMen4giOMc00jRUlreuvwvGtGV7yTrEY6WroP+Mo2f
dtpz0FDABR6Q9rl7C6uQI11kPbnEg2DCqHd/7e75VRbGhkHeXShd+IP/O+RLswtL
YZ1ey8VM1Wx/eNfVPwrsym+SxxJbiy84fUT14nDEPT5362A6oeq6L2HFYwW2hiXy
527abbOefX+ZcZ1jQGc38WCY0JXJTC6L5pixlbEoy4HujveTumTH8uZgdWGrVUsB
6Y08kaIBlesanSNWvfMce6vvDWaJaLkxU0fXoZTMNXjG6fKkyZFv8bGmieKUU4IR
IqYu9LaA16JJVoVS+V1JCv5UcBolZunZqj03HenT8rwaywJtfjYVBrYjPUOnC+yA
WIx+ju7cbdsunfRzvMXYb8BeEf5uq5nd+6YeOj7DLy16B9a/M6m/EQlE9YTwUG5L
F6bHhT33mFhVwtfl3kBNyHRkYLOJz9MlO/PMlMMVxOjRXkFxdX04r0m+2SJYgZJI
NeeIa1KNT1g9C4byY1908YuBpb7yRF+4boqMqadQnB/VRQUmrtz3OryQcjYGfcaX
/V/UXnf2nxZE4MBKRH90DtCTXrW7miEU+NOq8OfDkaOmChgiP9n/r0k5xmwA8BFM
xlO1ZBjpcXQq9LWUtlOeuXh4yrfivCZtmAdCoAyZb82zO0jRPM2isluQOOiSLiAP
coW8m2T7IVJlmf7B92J2Ou1hgDDd3IMjRy7cK7Zqv4vCr+jZ+EVnMkvgPK6fPAV3
iLxmT3meSYm3zrdHMRxbk8C8Gml7vDBIbaM928XT7v5X0iNOXvqHt9j3WTkIt2Ap
My60uSrgsw6ETsgXAMTjXzbg8FN0DCpqSTA0wjZRsVTjxRYyYikqd4zkIWDLLb72
dV31YBrBcvcRh+bsObeTMRNRTEgY91FUvHDMGkJlGiHNZsUZzovMXf27eHZSGiZy
rXik4Oglu5fNI0MOjwbinwnFLJ3GL7D+SyMZdaY18w51JQMWp6MEZlO1i+Lkf0ER
zWhuOGK4EzIme1HkCZNB7d+vvtEBVlqtxH0YfdsMFhULQhVmnWxonKTCmqJKOFdB
jr7m0UjQthrl3JK/jcKj0V5+1V/hkLxL506mxhgvcBfBwqNkjg+AL/ol7I8RvMEi
9G7IRUatlNJJe9aVuIZ/CleW3VCaTmLbqcoZqeY2urJgVZpaaC0//DoCo0ZiUvOO
hELnWfgT8elrTyo09SaXeaLIldOT2OEfFg1qonNA71A3IJj9d0hIwkJTKpRiHHC2
NDH0nTREPZJ9T82d2wsSWx0hwvIvTrfOc0JEZq0AhNgSfuK0OyrUVCpMZPREpAVg
aq4IWWCWmHEouclQZx0Fpy5g7fmWFRozLEZapJZfCVrKYLBv6BV892dtMN68yCng
TxeYAxnhHmIjPnesJvV1Ns3qArcPBLCj5sQJz7wQaHlgVGhSlQit40341ygjdgrG
6AtAnKLwQpMe0zlZZb9p+7FeUTWkS+dM9xRkoYqD5r/GHiHLWZztqYlCyxSwin1v
flam9+uSZUWFRiBvBuxzue/KlcRNWbg950UQCh7E3rXSlc9uJof2b5iQ0nP2hzlv
ZBvoq7fyjqmeeftirTN4IbtXVKunIR9NfOiUN7wsriKk02/76Ud455Bc63Q+bsi5
gdCYOJ/6WZVycv+/LFcHev2uG6hVThBj/XG3+0LCOt3nicTK7nchjM2xB3nPmGev
+Mx05HqudATRgvlflb45LMPL/HkeWbUUDHqAftYsosThXidk0psa+F9Am7XTkXSx
02PdDXhTrpMXkuuATJvGz6TK59RbwOrdRlNrxln8z2kIUwnzLsD7Mb5HzlTuam2M
vofoYOkfWekZzeDRPbS7PU5DxC+fv/JdrI/7uQWpni7ZEI1jdMe43LurMcJyre/a
sfbBbQ1/w76+fMgBOCOTMgQreIbdJoVUglSbj1KSKQYyTzsAQOSS9o9R5XIF9q8c
8DKfEBz2MPIvFSzMAnUUdXl+AtZJx9j5oaJVIZxrw7mpK6F8qbt6Eq3uIAGXitPx
qzoCOQPwSLjzsAM9kPH7l5UfGU7yJ/tt1jtKEmhiYSd1CE5aqLTuTCAJpxyry2IL
UHQwc5RptqL21Yx0U6ThYsOPcArxP16xBaSV+/kTuqwWe2PhqUxwtUVBZSeaaEBU
UHL/C5F4TUlEZXjTujZlZEYpUlOwg9WS6kFFdPhRvdfyTPABQ09j2a775xXpE6QG
D7K01eW11Ay7k8gpAeH7imbTpcOV2ViPj8X6zongoNB8BSYSuMkkIwC7cxQ7qXVa
UTlpEG+1khageeQmRIC1oqKVikWGnOlSy4JXJaRj9IV14/M9q75uON//dufDBvHw
x9IH3zeQu87nJR9NXZWkyXPPQYuzLm2IJqAlFpSwcg6e5uH6Zmue0bOw+PSrKGuC
pLdeFDvyg8HtURPUIx8S8i70e7q2Hzg+Wq+zp2r8z4dCxPpdHdoUGJGhEjjXeHLr
NLTWKC5t0ijvMgRNybcWaPgzo4W2vsCjizwZq/EFZCFaNzcTGe65iLUQQuHe0LIZ
72LSTGCJmZVTMjhpPdfqvuRNMJNvmzMsPK1wnKGenrAu2r6fiZ5VGLa/svywjrLh
BW8qL6MYCYqfhYBUW1KuLKgnR5WhqgZyQvIc4wtkOIwpGL9mOcqcuZIpKByALr5Z
o2Hlf3y9dF28H2D4plUR7D29MLGYt905obLBDGYTrauH1PDJRafYYJc7sfSK6bAB
fnrAYYiZViSqI9e0pBfDDovi3Keqq7mpvZQ1ba5N6r90YWOv6D+HFfLiQd9SlUnE
5JRbWVevSsMbP7QW0+516YWkVDg63gl3f6LGylIQlRkI31Iajlj1A3Xu7OztRViv
alABXn4D8DegrgJzKmlg01GiE6fjnRQTFTDLRGgwVFr0kfmA5YHDPF2aSLdKiuhu
s4tnl0AjPyZXx5gaXIIsNyax/hQswea7nGVSQbgq9kLkM1OBSBqZyRDe4WXRJ10J
OJxJLQx9aY92BNC6fCM7zNnTuzo/dDxoOm8MxNAm+/87EQchIlZfqymgYyb73sTc
nOAWjOPe2VV326UcgJ7F0jD2bqy7z9sL2WMM5H4vECuPcYktOnjH2nZjejktW+qO
6GQzN8YVgiQ4xYYHzLdmUbk6jzDx6V6K4czyeiaYPIcITTIiJ6NaSav/Qwt9j6ul
mqPOTRgIrtNYhyjzN7nQUP/VE/Kd9e6IU2m+vWRUyNBWA2xuv3aZuO2rxaEu7wBm
wsZ5dtTyV80HK1ZzRQpzw1hgnDeoNm3PPCLK25BctLAap5R5fXEInb9DLTwN+TJo
SLkBgGItZ9VmSm01e0yWzrk7yy5c7DJ9BNBv485JhtXlDqHEMqV93/pcCQqCHtt0
MvTZLGJu1uBJbwcNGtftEMgy25plsznKnh+D3Z7y4DYZC/a1Fh9UlPKXIk6YeQe2
Lh6t87HdaNLCi2krKPAJJuyMrXko+Nqovs1aMtYXyHZOBhnQiaL0HYKYJHK9Yo1D
EAcnR85dWW9T/Pnn/hvRpLH4oEgGvA333tgK1+BKKW0VzWsuSVWZ/EAC3qk1lQny
opXy9tchYqNrk5YLhOE3Mtjh7zOHzwS4EoI6mIdr0TO+YAd6vQqrZzFSNqrq36pp
JeqcuRMIXWPIUpQ0goTzX77riW8uCEil/ujazVvYonOCVN7MrxproXNZI01bDl/L
/Fl5YCzBgaF2EuwzSLn97aqXA8lm0lb7e+h4VrH3u3vg5LneBap9fbK/8yP17sUh
qR9fD8CLT1awR3Acnwbea8dfdy+Q466vReldRAtOoRxtrZ3MYPeohwo5VA1FTjZL
VDmgAD9rAHnA0DqE1p4lpb1B1aoDZjEmTyIhrkhZTI3XvSS3R6MA3sQCp4g9MaCW
GNMMHbf7Z6j9Aad1zXOJxVXQltHvMXTfpLOov20xvazxAenWQRoP7P6jBvkeONW8
4EQAPKoz6BfhxMKsqVNoHDsy6qMI6EUhvUjFO3RZ9g3y1Sc3TSqrDoqGHoDG5E2E
6O0gCyx4nuiijfvDAb+WwhSwzgX+RbqW9G58bshyhiXi8nJN2/bMJByW5l7lRkxA
a5t5jyCayGCn/rhQZ/CZTxaOT/EQFczO/SuYUmhZhL09OMBFs/ViJbpJ1JZqEHzb
pr4WTFznQZsGnk58yqjse0bCIMJwiaehBFVeCoanPJ3lQzWIrmsEQr6AX+JzE+Ae
rdD+1NPL9zPKlGczrHBU0dHMiN/fFJ5fWySqjWuhE6RFdCTrR1DJUtCe0MT1zCA8
tCzURfWwF+efEMJ59nNaf8Jcu50DsWCLO0OFeQJbLghej2OAemekAVpWAWxGSEWh
rZbknBErcoZHN2smDpwR8a064wxCiqeavVF7pjxa/8VSF0b25Vfdq/Qt217huB+A
Pgifoeph+iN+RmFmoUhcCMxlOLYK012cSNPP8NJIsZCHwr2nizCEcjT+nWqP7CcE
BJWXYBmUZ84XOyJ2QUAhS02pssGT+ZL1GmSbawlu202Fe+np/l4nh7C1EDxzPVvK
VRhh2IDsohDpq9mQLEJhzWdKRwXwDBo4+yKSyjscXuz6WeCc8Og9psWpYl24sGGC
kGpoocViFc5WTLr0QrukevgsMgV3X3MvTfvcB/EpFIXLj755qI+ccyobL9ccR5ZS
7SnonAsgNkj/7EBUgReAVMr2/CqunNZkj9zlYXtYKBAQLvvT8fXuVuuXkz22klKb
yiF8UKPHCwZQ51FmDwrC/MUepXn+rhxfxmQa4U94EA6ckDVRY2RMbQNezawp67fM
W5wLMfD0rBd+iQiwM9+zedmdT8pYjdQiAIROZjxWoGyEN9Ekz96WNvypW4JWs00I
jQ1C81AGu87AOUANYDM9w/IboKosglvUJdRizZsoSFsMAp9M+RLVP6zaKI8qnHYa
lBiYJ5YTMBZ5R3CzclbAKUZmgiHiXqUAw74LyDvAUhwCmkrCt2FH32yZRrq6CCnD
dVGzLx9svy6TRHCMwyNt4XEtfA3vWQc915+EOL2gScoQHRQMHxRwaqCkaW98vqpO
XqEJBD3CDDuvF+Q1RPy78z3uWAyxuSksq5dtmgQS0tjUZFpd0yLtHxdXyCrUKSRf
Y2mgc97COdCuN7kjOm5O72asMSScuJQWYduoN5oZi6EZLw+ew/Wy3WnJQiwzCofw
wUJ/vUfZR8IZqP9ZUnGwNYAH3FAe6hRUjYjZuRBZKcwQsesZ61F03nCqU48N9HNX
FzxCU9Sl1mrKuTS6u1LMeTWhdrn2aseutNFYLh1qvxBPp2BXES88BensoJDgRJho
AvRtBmjOfAhIFOu7nAQAm3VvYhGM+Sd0vrsiVSUjVLlhUvzSgVv2JuF/1uMzyIA3
sIHXtuaSZgPFr00Gp/SSlnEp40IEvV4Edq1sIoTVcvBkP+Q6i3E8XUavsxW2CUMq
fBIVG9MxPARsiZidF3yJel7OCwaJaN7cSFa1/RSARfgdlb2wTzYpWIox+BCRhk54
GMSWG5uPlL0U2ok7LA1a99udrR1vv6kIpw4HPf+02gdgO9ym2v+h3dEg3UpHFMUg
xklyUMAogqkilFyqYPrmwPjBmpBBihEHHGC9pXF2gWzIh9mrEGYk+1BZQuW/x9BY
K1jXABthEfHGCk4UrTz6Gk4lxhiN8wY3xHdHwKtoaej8OG+FxmXu9UglEAwhxokP
/eP31Ja00eGe5yABcwCnB0YhG32iu3e45DIP4yV23Ic9cb8NBeu4iSYJsBg7D/hA
mBwFrWFQQcIhm1cvC61vIbJzPBxsElBUvHrVAKkT5sNtm11yHgOyJ3J05moQQcx9
lTgXCqW52EdQafYystZsFN5PO0M+C1yjUC2k9sWTgx+gaCdTNOnw6XA+NgNpmaJ+
rr6O4Ert6NtmRq7TWG+bRIWOL0OyTqodPfRiJOk8l+kRfHEJ1QfezJ+f9ZzL7+kf
GohcnjdZmODvCwGCsKBpJnRR/KzrYXtm1lviWUfJ4GdLuQaTHTgPMun4qjDJI30p
3k6QXR2opX0q+aoi4oSTr0Ow+oGheftSqGXjML0LRXDQlhBOOhd8spVQcIkUg+2R
cuV0snoPTLgErd6xVaexPJpCCJNfeJNj3mbnoFOWX90kV62JyC923NlU3QnYHHgI
BfkG2pZvcFsQXE3Uko84T0H9MrlH/HXbYEPgX60uXOxZcNoM6T4+cvxuLeiDQFVB
DgIUjIafQWnSTiofrAjP756khkh0oIG3sVIK0ztIrA7bRvOVO01WDzwCG7TMypwn
6rz41rNPhbel1zS85JRT7xMe+jxIUKtxuZS5KiZTU2AcNJWxseEO72KDof3rMIa/
0GL2j2CHtwgfyNsR7ugCEv1VFOtlbSUaREncNXXE9BTwgMEzZDlSsEvP5+OI7otc
az3MHUdB5BNVUL4txulstK2XOtA0zDPNlsJte0BBuCsR/6QOaZ36sTtgZSMA1Msg
KPeCPk24c7mcEK0TReS5XeJZKx98Bz7FK2FzikuzXW1qR+vfAPbbkycK2rST1I7V
1UsMdIi8xzB3o8CzNvPQNG0cCbAHM6R5S0SQ9AMRkwED9XzxLa5bjEJyHD4Dbn8c
9ALxE0N4AVZWTPHqktXQU0TUamBVeOdTp4XvbjHaURVGZ+3cSro+lEmoYTgVpCD5
lDYh+L+mdO8dzncEDrFK1JiupMkCyE/egG1rLjbqxe7odeAGfOcZmAWGJEjVX64Z
ztvfptlqArBWm6HExeopJA73RcKcd2bIsx7SSyUA1umalHspbJ8aZzeGZRTPQ23C
4HdAWMhi+rQyomelF6S80zFbfJBPRcztvhmfIMG1wRSjgmly2n1qE0BXVSReazMh
HxhZLd7XvJHSL9WvJwJDh7m66tG9Vc87SgIi6Il1w6rl8G3DU9yi+U20qxehjMgj
RXMQIA8XPAe7vTOS4qM7s7dC6ymxLCtL79UrqN15VSZoS7xvLxqYda0pi6g0X5Sp
hZt/0pscRm/2VQ9jJA2nqvshdX+Ia4vYpLGaEcmL7X8TStnQ19m79+ATkC/0QTzN
gWgb3XjcaUaUEoiAeJBqQp9qGEbm3v+Gayups278LPum3O56NgrVYzhX83vaduaF
mQs/ij6v570crLXYJBuiOT+UamzljzZADzN2shNgvzXAsBf0dyIzzO+UVZoyxvic
rcKZQgof+Ant9lMwYObGluN/bKJE+rdmox/NBG1y2Z1rKSC1h3xCLkQedxSZfcEt
+pm3yA0E6zbFDQu8N0vOQyoJvTQMdGadBLeoy56D3Pu67TE6fJVLrPEKWDe8Hn2X
NXEMWMwvplNgfkVUmFoAhBZf1+rrNUOgWUohEdb6DCjyjKVrraffnfShr+OIrxRm
tFTd7NMQi+ZxsedAgjH3UWaWVTpcGkgX8dsnY+RqXa+i/eAzRURGnF7KnGmP6uGz
z/G+CVOFlLhp6BNmUfsKwdl64dgvmZBbUQfUD8PY4JfbEcLFSbrDWHOUcJBX8hq5
nQycWzQ+dr8MbQElsTJR7NVncPqB1cOJzb0KLQ3XvlHhfhE8ul7vE8WT+skjzE7P
p6LAfvej72a7WyAiBc8PJ7sN39Ud5Ooi9IVu9z12pXRVpqFDEKneq00qBrpH4gNl
WP1ZPxtX3kx9W1Qsr9RBbjFtyATdUF33tlo0GIGuXQEoGcV4keVwastEeppfITrH
yIyBrGytId4oY+b3QiLK8vpKX+ffPeILa+wHmRyUbDRnDyEqbRQf2IzbbmiZFiKN
SH4yaem/KHjjQq4HwEiRqLGOO+iE5Jp0HcwEc6us/fHr05mecPKWdSGcTDJcYPoy
WVLtT9epBFQyXsvrzOE4A3DVlKY/I+1HpKByxL6htdUWO9baxJ86GnzbyDNkPKbt
pr8fSM3ZVn4ovWnT6n0QKIO2RItyPBPTU7c2aC2pa9l6+dLZfC4+K+U25+GSb7ce
gcBFkjqhopYn+YSVvjrToVlhSRUu43ZvWnM+E4xR6jDsQByGWUrPkDbmzm+mVkRy
Jz64y+/oA5vwbnn25nixgXqobuwQP9FBOHhsgWDaKp8PK5lWMCrQMbiTkVTezZGg
tM9y7KjE2WMrQJiwgfmYOm3GOeyt59tlqTqizP5dHDKXPlA5JBORUE5DONHq3gx2
l1eu4c38bt7HeL/dHIqSf7X3xy0mqTmogecmdHOV8lBPQNs6n8ZyLFsXhKT9YxSq
c37S35ZGdZJL1u8snSFpNIoTeYngeud1wQJ4eIabCfn9wvyny10pf6mpDfqlA+Vn
DK90i5qAEzXSYJp8yLbafDj209ee9E4uedAul32iX76/YuFEvK6+FFBBdsJW2wKJ
f26TzMm0fMtwcdQJuULkpgoCtHbXwD6QLilpXNuTQsmjAXQZxwcbqPq8PQCNHZoS
EbeGr7yLOiXQeRXCBvbuf7iIhUB3nUI+4toqRwOOLdE8s/6TkpU5AGDMTT8B9kIC
iCKV1SrTXmPmPKZgA/deVu95SMOHDpqGhj9VAuXWZUhdFt9sqthQSLL2PgVXMDeN
gQtolNHdv1Ou5bGRdF9gGz4xi7Is0y0G6sj+QKoznizPxZ0HQ+NES9+tKXo4AvLb
YPHEOh6KDuDgeU/lcpf7NSMPvRxuPOz4d7BKrI+n7WaTSx/TlJfzzGwmAK3JyKR9
VLaPW8Ulv5+jPH2W8l3sQrWrFMQyRgUFJFzQWsqLCoBoHOvOEtSxZP2MeowGzeXp
4I11n0S4G0GGacyayTgjSgGdy++/DIRLDVJzudTDiruDNs+8mVirl1IvwrYfBz3p
NewUj1a2cC+aN6ceY8LVNhQjLUixwo3OULc0i8nG8TSG6+WBqarZd0qfvMId9WT2
IcRePY9wuyQePipNTPee5eXW/sqg+yopswhqIu/XaxGwnc247p4xV3gxDAzQ1t+j
E19cRecDcgOTWRVTxx1nptd51mUDUwyGYXyyG1x9ARCPC/+lT2G9r2/JUs8gtwu2
Km6MKbePDHlL/gn/DVR6YHmwZqZqhmS9dAcj6vdYcV1Ugp4GDKBYTy//4t2/FiTO
wB6IRfVcQolqarc7IePxJKIO8F0/8PlQOaax2ZxSwiN41RRk1MdarDDYWEI2yhz9
/zAillyaVku8yjxWn2yjvdtyedhsqBNQ9NaEa8RH9bh5EbFtPX6DV8e1OAvgnbc8
Vu2nV9WFX6s7DkOPdFmebO55sOsJ0F9sTFm5RW351gLhwm2RaBLpOz8nMWYfSdlJ
fh/kTyKLMbeQhp6UGxqxejmpDa+5z5WwdEfCvDPD6QJ21YZ7n7cdaT4NbHzNUMY0
I6phTBZVJT/trnAtzrbMyKtZEqAfoXA6v7uhlGOqLnvFOvvnw/b2Asqqk6/6gJXS
pRcxdbx1eRCcR3q3c1TnPmumN5cVKHEfN5NAxhsUZQZBLb7c/9qk4c3kQ6f6qxTs
+RID1QnPoXoO8gmSfTiC5/6gzVYbFu4R+1kOiBGL7AgNDz7FsWW4eAW6hVcjdFkl
J8ivDUmQVQ+l8FDebrIGFS7VUVs1ZstmjuDr5tJxxa0YYSBJwmgQ0GcxLSrPwVcb
/XzeZddWdZarVN9uvKXIQDD3RpJtnALRgyS60Dy5c2Gk/0xlDOGKFe3nLvRY0iEf
kpsT0QQ4bsAIl+jOyyeu6Hrx18DNsa5i0wYHwW9SF+QCDDlw+97LWGw1a7P9m2hX
ef1FlFkSx6Ic3I58pBnRt8OswwZJaqinjYleCRzPzAsFMxkvbsvIPAUZCOFOc5tz
syd2b13coE56Tuql+gBybzVPDd/rc+Z6mESfFk6QCX7Gv1Rixs/qxdSEkOaMr2Qz
+Jl05jjjXM06yVW1rkztk1TKd/urRm9aTtJb8RqFdMbrzR1Xtvb0E6UqdIqrVb/j
BN38RWmSvInBKsWUwb0ruowMFf2mYf5pqveqlJnxm3PnGRodnnIEKjLFge7naiS0
jHFzteVSbF1IMGqzIWytgpnfEPiP6LPzIEI1wFvcw2ly/HpXxx5PgRY1bjqM1/xU
pyPSQXbDtvJUtjILlmb2BAFcwlE4INHsQGm7uh2EYSEoQF87saJhULZn7/Vrrc4x
+2pMElhuXCk4tjHIreWeiWkBHlFoNRi/sdEqjIBzJiJhROGVm6n8dkfj3LKcsWmA
zdRDw8+/As4NOFtBS5eXyOyRucNH1cMDb59LcXI3sJ4Fyf6KXkpBWgeMgsSox0BK
KBKra1dq8IffF1/EODgQy9C3rgwMh0HQAQOK9CyWwvl5ACR0ezE2//LZAHTzD8Hx
M1xX+9oW42CiDRklHWkzLl1WNQPLHV8OZJ774/rJpAFCYazXAvC/WxRw219ZtJHL
8Xr9DYbHACm6prBYL6S+FnhEJK2EJQuCyKdDaamhxYeWapiVa7vLAHBWNo2KCqKv
1TYg8KO8SphlWcBbE6GY2a6xMw7QTPsYtKAzH1dknoSH23+LnUsJz/qVzy8ZoPcq
KvMat9F75a43Sk6fwxCQsnr8nsoKdhNQeTjDRLl92pjQ9XGlLkv7O2xhApz8ZkC2
jbT7EjFSDj5BVuXCFaQcMXJKPvxtTL4ArAZbiQTNMMb0Gste4qWsR/PrQqeAPv+5
oKUVUfdU5Za6WmhsuoQhviJ+fSNcdXl3IBPAneeYMnMyh0/hDU0gL2j6UJw34dnB
lvHDq9rAtIIva/0P+yjef0lqwXqUx4HdOAKXGBA326ezzsftMRtAYLIMzgp+E9NI
vyRgZ1YmGD7DZ1MX9uzAsh5uwCK9QcVOCKWcbmDmGkr1OI1d1lx06nxp/4HlU3ec
OYHDiJHnmjyf7fd7sFgVrdEp23fLdxHNVnlTq9734HsskdxDf0pfDvKTeiSWxKDc
WoRa1NXQ0K1qWgmodvXfDfESdWOXT0DefJ/34r9jeP1ony1KTh0zGukeN23aTano
rybSf8ZC+jTOXkJzvsP6Ywx1U/V6W3UkrKNavt6MQZNLVPAsXdAiw7BNGzx3vdLR
g5VcxKvpy5pnXhDaQoaVVsH3u+O3zMnXu9NEkTUcgs/gSg0dtlBN+upwltZqVPb4
eMiWPV6z02Kh5cMtX3D7Hu1yeLiup+ALBYUM2CE6hzSCt1lG92wSDcPVuA5mwmFH
7XBakGVZnRsRh7rLGBPP+VmB8xn3xC6fB/A2ksAZwoV2WqAoBi0zWrt9D5pTS0Yv
X0q3YvmDij9kEUoimA1nxj7IMQPC7b6rmNX80eVZGC4cV0JrwbqApb8ijLbwz413
uT6O9lBEqgOLBfdeEgm2XrFd4c3NckSGs/QGcw3ZntAYpRLmIi//AEcSJv3MUiP4
JH2nYeqwW+7x/iOtUOYnDkF00EVfO2vKNFCbWVI1BU7fY9UqLwNQ/TdN004CDtPo
zTqIIR2OpVdOMpQiAIGiplNAVve/kmOMi4KDO8jyrt1qDLepIOHpmcFa+kjoZbpv
n1ewRoVxyghnAZi5ylplMKjgITMnv4I0ZCVCtADNt4C45O1pek8M7LMOPW5qzQhK
+66V+vSfdRtU2hkcmCVIHXlOsUiizs68H9BeyCMTUEunCCFA6iaGvnXohAcAV1oo
2r4Y4+ucaK0h35ZKHKlER56cfpLvO+mt3wqTBqrtr+F4c9G/VbKhdfsVZEPaJE7C
0nsPXySZCS+SQhc6biBw2h21KzMF6l3XiwLQHBfAFzU1Bt5ItdUFD39E9NMPRBUD
htMBimbkkFQ1EuqBtDu/902wDDFd9MY49nSo/Cyg29HjO47/w9qgFgix9jQ4U3lf
mxTcSkIIaPpP1h/+RySU6BhhZXhKI12xJo5O4/gatkw/VTC9WaSZkSrFSz/+QZSN
MH285X6pn/7FDw4QK33nPbf5u/XKvE9cdNPBueq/fEQAuCnSFyy5j57pz13koVnq
qWrQPVpZ/PV2nmbWMj9NSlkqbqmrNcISgICdGyaq1v6bbOScRz07FCnwPWuhF7qW
B/6TNysgWFUpgbQPu5E1I4ZIkImOVffBCvEyUBgkvCY9dGRPnSp+qANeY3UteRoi
m5QfbbDVPjp04oeW1RBxlwZjlPfFIZxQxy4V4W3rRRYbcQUNbpkJ1+RTGKFzlEPl
39Z1cdnkp1kP1FzVlTw76paP4LiBCrNH1rk3qgkBjl/OOLOtcRBKyT9CqJCoOBXm
QT0vQ+h+FpCD79fTH7pMN+TKOivGlwOG5T6I6kFQSDFoXahvz6Q0iLUFsVc8pnHS
/fX9DBWnGbSrqsgAaFOeQwV6w+n8rmij0ebHlGI5ucvtm65pIMai2jXDi1UiPiHm
r5PO2HTQLkSjivQuKiXIkSfCslYO0J7KG6mY/SFVXcin6J9JOiKd2fan2xSONk6Z
N0oNA2hJckE3kKVcp4A+oYoBigWV9UE5KW9ABZyglCn3Bq0NrM3LcCm4JhvRKM4B
g16Tdm/nh+7FB491lbrf7lyK/gfIU81aR4zFitGePPIdUX4x7om0QIl+RsGw75wd
53C9t4K65IG/J1dOqH+vhfcWYklsuD24TaQXQVgXibda83HjOw5KWXmQkyoYXsK9
5pnEhABUCVgbwk7BOICI3AsCfTweAtid7f2t45XbvoEtp8Vi4ZY9M2hU3oPkbgpT
WEu9F0ALBZAUIymW8XQ0PSwyJwUcET0gntbE402Z26CDOu8c1/7wkaxagqzlXPC9
cne2dlT49RSY8TJxQbeJcgaGzXPRMfLvDvPT+ZOikldFnHu25TGV/dD6JfUJ2ivI
gI4amaGk2M1dazVkNxYRiauIQNrpVaLVxM3JbpyWikHu4sKGnUrD9fdYD6iWXZSU
7KdfmQJHp6P7LMjqwrTlJiAqIyK/OkgI+zGy9DDC1uBn7mhC4rTQiNZWk4SccEzM
92f+3ln/fSoDtepvoBVB6UPe4eipyndJ/CfuxQ5RHLKLUVq7QT4cswqHZpssfe57
0LLXr8ft4tOVYgy90azoaVLNmTSBnTBrAQthMWlph8aQkHuQbUc5F67JeGBOPqYT
dqWoLKa4x5P9pyY2yFMAF9FjgwAQFJcwhZfbth82tMExjESBIYQf+FVJafOizTMv
MhmC5cdcnW3eei+AYN93ex0nuyB6Io6u4h+5nmMlDpFej9ooak40mqGoHGrYh6h8
W0QPngLdExalD9Qd9zPAfJ2+GLbVlIryeopf7zZtbNQqQU6gXCYViTjdqPAYBtoG
RrgRDlxQmbcKrcexsDycdpn2vjFgyAEXsukDxX+VmG6q+MuKY1S8Pmirf2gqHs42
etWajuhWq3Ih/BwcwKh60FsJzYZYN2Ky6Det8GSyBLmGo5a8NYiYmJAW0RpQ2IBq
JWPvFNYSEoEaNNvtvbBD2N26eTVHpSiiQQ3w0Ssx01BCEGxhSS0PJiNAZnH60lWl
GXR3g+bnN2hBlDPzMwlHrWKiPIICD4SCzMeQLrXOW8mkg0Zt8rK2NdYMLUrgtOf0
bkZzm2w7GAECsuL8BTKH4OEy+JSmWM7KRHoL1SGkkDnkvENv1OR8K+AantR/pzkc
5W3oJZHW59FqFhgYBogbbsjdjbRbRDPZ8dKu5LL66VBgJTQ+ptJ+a6/l7YDdJUsB
aT8ssNUuZen8p2S+te7p9oPDXt4R4dNNqSbwPRRuhPuQtjFJOSMuKgGvP55EnB46
EY798e1LoPHjjBx5lO0uTlNl8S/5b3O74OoUTdRrArxntwdh2M0Y2kMf7d8SKnRF
tp56VZlzjyO/x5N1WdwDkAk/V3KEk79a+l5mc2egojyUH6nXhTS0Sapa4nK9nR67
dTUTXhuOfWW4X0wEUmbyWndCByujfPdp3PSu02DxPlhrJpIw1tlnhgCDqyufRi08
ACblsJ98+ZDOLPgEuHIE35yZllj9XLEPLMTpHv3kl9uuaCPcLLJkv11qCjR0vRN3
UQrTbdb0eZ6M9YCebF756+Xz9EcEtp52O4ciBSB7/xqY2Lc4XLhGWo2UGEK6NLBt
P/T20+i5ZIuRC/XXtkR8Av5O9KXhg+yq1j2MgsOE+dG7UH1mZ7vOKBOXTLPH8Wst
H4qvpenZ1jthrkuVAsxkfFFrqCUWJ8wQZQOpphbsQERWHWXZcffD0MRywYJjHlF9
La3PmwdyhdPvm8VV2LaCW9TCjY+sO8EFWdEXqZyQ/w5gKgFZrIuY1PNxjuuTSph9
zDQKvOzPua84L3DDvUMG/Y1mirwry3eACN4y3ap1+SPGl8CrQpNczbgVzLc/8WSQ
lCMU581XqksPi1v2J5K41RUIvsxMnoHEGdopInJy9eXEQHDCVpdckpLdjb2A+8BC
CP2SX79bC/S0n80VZRHy+wUbRDB4ZhtwrjrxHkawpJpRP+PgMrn1TIoU7n/lhMZZ
VdPS9fE2POhe4ONLBynjCA7efaqFOQG2uJlkHWT4sW6oVV0X+dDS+g+TtBno3+/d
oS94s1VgudpF5SI1kUl8fRa+mtjWKdSErfTGUCNCAJ08ft31E0vBSRTkcMYjeXaY
2deC8YqFo55ioa64obwEBoejHTQnCqjGLYm+lGq4SnCFpgK7+w5gN5qWFQD+FDFE
QvULwbtO0FG9pmCHF+QsGIqt1Nl0hTAn8Llm7oxyESND/QBlcPMVKDSHGCLwbktE
f03PMAx1k6ZiqAQYWn94GvE5sh2FjqWvDP7viC2EK0m3gE+302Giyo9LA/EtI9w0
bt0Fsbkjn5pAQcpsaJ7/QbmcNRSodY+M71ci1m/3Fv3VGKGwSP5RAqjEDsigliFT
pKRUSNV4U0RrKRxmN00ixnWevatm1ysdyxXXVRxVkk9bmhL4KmkzrpIcjVJkquoC
H1udmpPuVvovBAih+AYF/3r6bUu/ZDPlL/BVmykX1GOewbC0ilo4iyzL7FtKgvDD
6khxAxY58YS3B17IXgJaqGWyysXJA5Z1UbAtL+C9Ak+QYzX4ofDRLFsU7lj8rm5f
yd0e8n+wB1ZLB4QCyCdqNDZKg31YLXMSoWeo9OeK1Oa++AScdTioA9xN9I/2OAjn
yoOxRIHHxIhtVodhRdn/u/4g+8Hh9rDAYFjAT7oJWLdkToMyI6/7dzd5vT2w5A6t
mk4YBfkdB0uTVReWVV5hFONfG6v8r4ctQwGTXJZEk2zM1Zoda1eppitAXsJXiA7s
iVSBo56BpRrLY7XhyzRz5lIjuL7pHJoEVYQYW1Uv5cJPUVhmfA8/OyWMoqDGub1v
g8+Tj7aJS1zrzsiawYi27wYqZvUy4lE0yzuw6c3+U9oLmzwk5OcgqnTjmZthBajd
8MGR/VKPwvXAPN6KOBPt+zqn6Z0m/5ywXALpdBx/XFA9mqcyt8Psm6XFXccbcm7F
RrYXAbxqTp1N0WqP3MJlrEqXdMioGILrW7teYm4MQ3fEuw9vip82Yo8ZLyJmG4Uc
a6/WneppqWrLdIj9ImaCTdx0fQfCU799Z8LrE/82cPdDhmLG16qPLWro4oz7lJGO
PAOLor5Sx1i8CqYPSq6W3+Zx6DJ8gWaqDnOPhDKX34DS2qOaqd4amja8MOMW60fW
KxW8/hZznoLRfcpVYu3mjHeHAQZJCjG8SKn/w+sbaBk3t10aFJZR2jNbewoLGaQQ
57e7EbFrfcCZIZAcsjesX0GTP31IeEkC6QFeBYvVeCwHRHzPz6iVR/XjjmwV/2BZ
qy//urlxHE4nV23tFKtUdXYwQmRwE1qds+ATdX7qVQYR7DtWWSuK3O3SbBBfab77
1hE2Cg1J2cCDHn0FvJe+8Ud+0kWDcfC6ZrSNNCLxvyhLX/LWhgxLmTL5CpZfWCaw
moocltRDO8WkX5xC1M+g6jDWZVXtY76OyeZNG5wLu5em7Gx5ADthDIX4XJIKf1hv
Mj82Qx84sR6LPFFik/6Cjh3WmWSsLwGwpAlbpb2Q2AVLFBmUL4Wx5DaXtE5rLMkI
GiU16jD+ocCf6lHWCIMOmzFbA+sSzsxiC+2iTpXp+Y3bqhCYl8sPqEqXSj9P9SjT
K+kKidlxugeBles1/NZEO4atC7PykIcmPgXAT0cmJc3LNjHmznl+rASMs3sjdFgL
/44hacsCRdqeEbKOgr6CcCV3L/gD13ricRmRAlNWeJsnd1AKdRXQSLKpozfykhFt
Z778bp95rLJdhrsb+32TaROfGcqLNlvrdx34uYWt0W0j7jKrLTAt44Otah3GEh2B
Goir8prgCcGCLO125E0sbLZqPeq6Stzz2rCcUC912zH7c4g6jsL8AVnE7gYjShC6
Gp743G814MTshSOWnbs/FLgPhR36XCAzgsW8UxWYybUS4+7GFZKbrUcSUenfhb3q
Kzx3AzNetLchjk8qCajFRoa7EFq2Fykfm1Me7zFxcl5MqrZfQpOj9P+Af0AlwDqX
V+/YSI52HWYLeJGWswa1RVNcNaMtXsUdBTZs4b84KDIovophzwVESKsFP7PPsUVW
pDnIH4tVxeonFrYy4qaCrBLSbibdBnU6WleKClDZNjv02YuVfw31yiialUIT27cp
XCYXq+f1IB4iFGKS7veWBcSkmPLDFUIm6e1i5wT/tl6LjH0L0fvkFZJvtpbC8INk
5cgtf9l7OxmkAmkkYuvRZu53o1KBGgAclbjFleWtS/cw2QEjvdmwqA0dcHhQkd+h
NXkqbHoz07F9hBirpYaWaYOUDO4qt8iAoFqRa7fVvEU/KEX0g21E098XhTCGu9hm
E2GUHr1UnoCIK1j4fyeNI5Xn0yeOtiXLmyx0lzvkOOrlyOwKT5tZ6XfwICg6RR0U
3qatapj9EA6Q6vXu5DfX7c9H/NFiOUhyYTc+NuAlsiWig/FVw2LDcSYkqlOF3zqw
eVYBb7/MCWUbAhUqw7EdQ5ncEbzqCQaLLlSc6Ni78093EOowbarm9+pLShrwsW9g
yDdqHhb90IUftKRQaZMGzlhcDRSC20GHcpTiXLbjLqZuNlKzfEGs0mrdef2ZNViW
DkbZ09gTV4vYIynLZkrVYQg6uMqSNqB2Se2KcFh1lg++uLX/o/E6j90ft10+UoIG
KyGpvGxmi4tk0tkg8sU+fbXbix70VoD6guCToeKpgjasYbpqp1eXlfN/gyEvwSj/
Ai8uE57FmxTx9I5h9BzZ2WwN3qsDWI2+rJQqGh2kpqfe7UlOUBrBPFG1/4Dr+vSY
zQdvJpolwZ1PRxilqPP2/cBGyA6/L8J/zh7aQ4ATc0ve7taMUv/5dPh0NxtIx4yz
LWU+IWBgZ3mMhVN1R2vqfi8x8U7DXFDEhKR9j/PLFABeMCPu+SCYtkH53/2ze/4N
jUx9wN14xFkbHwwB5E3M27cibOTcZ8zB0kXAh0vvAQKMMpeWYlSP0VcJZ5BklruT
62qLhKryO7NtwEPWIZ3zUdYChJ9jTe4LpFgXIKvPXMFll+1KOBSpHx4hH1x1bnGt
WBPrJBcO3y6rVdfUhWYJ+JdrgZn8tOslzT3qc2eCywZqFAGurN53JYCONyXspf8i
cqbpYr+LJ4wc2tzvgqiaectYWNTfZwlf6IXgmudy0rToT6s89aRS3QYiMTiTB6iU
RtjlDVOa3JJumj1M6fhmdVXBHtoDPmE03C5eiZrHOEzUCVScpqEn/cKYPB9S4b4Q
JTVe/SUB0K84Pf62nlzL8O0u2kKdXbRxysVy/8aS932kJeSOdQ/xJCFcV5C9HaaC
ntiD6eqv4kggf1czPl2ijDMemVYLmCy6dSYVESyW132zlI3LiCkcujS2VJUWC3qB
4yaTsQDPPSS2oKs4OSpeHo3dF8UA3dHEtxIjRJ/gDWAOmroUi+H2cvWh4jO4QWnt
ybQPGlIsisB32uOB6E/a9LwgOBCyMLIfrKFGAOsANFhtsm0UerxhHDamjl1rTkyd
7pMrgzgmjlIIJ8MESk639/KfRWwVNof+uYBQLdBBMosd//ostfESztco586D9O4Y
y/RjxgYpxUSstblm7exbC/EroI+RtIxYxY5Q6AfEsUnOiD/Vaw5UmHd7HizlTuyJ
fr52h60xsFSLGFEEQpBJlmmrPjZUGRCfd6qeyu1MN+mynBNzTjXocKe+sZ6kYXSC
WavrEPwEknwBlcmxCCJrRgoqls7AnqEXc340Vl0H+4hg43fEyKyz8ZN9f18yDoBM
uCCJpurIh6Z0ea7vukDlXIrBwEuX3ZX0GrHmXoHEymDJg4N8crG738DKZuPK92e5
6KNK2dAdPWC1spisLQeSYyYrwQYacjx3kWOeEVC+1uBpf9tINaCt09jSiqdq1FiD
mHjPXY+GbneIDZUSyJpHCQgpFL12hQMS5OgAtN9FUEV+KIrXdZMTeAd87wSegpQ4
aTs7OpSGPxnImpkpJH+Ub1OWdK2/wGzvbVGRYUh07Tn7/L2Pt7TTa3Q46uhZbTNS
smFIQABLj1C2aUtiCb+34eVyIpY6uk2+TTpW3kO1rsSDv3GkQmaUW9EYb9jwV4ZJ
u6AyoXDTrELeDqKVZx9Gc84ZuSENmWHgLxTPY84AX6oYaZig+7frFjqtUXLdqqfk
elBpij4rQXtNrx2XBEEVEKqJN7fxb9miwWyDNA2UTcv4Njb/YzT4nTKEHGrxGfrO
FTvS65fK/uYeeAJ4orWGvgVUvl3zywVFRqXAdQVej2WefN8PYX+p3+KY9WwI/lDx
yf7YQsdFWAfoZrtCANhdBnddNzlWZpbzUumN3TZum1jiDKAKH9UoYu+6d100epaU
c0ymo5PSAZ0XpH4zrVjCQGa2tGi1C0EtW43s5mViduw7Rz/nqPN/e6DRh/Dgb95W
yX5bJ1WkUiZHoysv+8rpeRVDQrzjDHK+ftvvgxWjBq1ELC7ZFngR9d/fHhFd1A2h
q91HGZGt+T9YFJQP+P2rqpFfNEgFfqkqPYga8uYEtFbNZ7UlRTj8dDh0jbw7wA7C
4WQLYY1Q75CKrSM4ghVeBj638FeE7775L3dNQ9Dk6NiT+8X5hw7D4Ut2/a2UWBs2
aFFI5OPHNlft3R7TCMcADc7neqi+3LbDxsW76neduFbVQidgLf0ikMpXjaSclpFH
OJ97oLt1++1l5Ql1HjyiXEI8CxqQFN0ivbFitstb0TW8HQZn8s5spLPnDf+ZotNB
0mX69m/gcTGjGmEVXv1hlvSx8G3z0jpNX5+9379aHxWXya13vAwdUkUPpehKd6uw
8vifEdsF06ZNCGcQKAcW/AYU3Lr8jwVkHtVS66rkvNdyyYBeRULZ85ZgOby4J1t3
FOZTN6Ud+zrhmtRoHBNrcJmHHBpCS18TT2VBOmyfxjSoQy+S/cMhVEOiTyH16bea
Lk3iNMlnRvl7CczuIxCOn4VApGjKpPVWgPMfcibubS7wKPvXo4k9O9+btgEG4zBb
nFmBLapNj8lZRijiqlb7D53th5FSP/PRszyfxVyLpUfejJuuyUzro+dBweZatpiu
MQuGPRPVdJ42/AurSizfjvFLlhg9qVlvxbmnq3Q31RfsQFMoB3l1DM/whpd9OYHD
EQpeoHJQlgO6dTEQCwzFJpklAp4q5bHMa5U3VbchAaa4xyLgiAXq8T0uVAMaNSjj
TPh9bFZfV7OTHbkmJezjFjNGfgEIlXloWCuomOH+IWHwaJ5kWZi79Q1BLTUUQKXW
k/6hBDZM0XHiyFyLyWOljJyJsaDsMijVHNltscrNsU3ydTh2NFEmKQbKHu31YY+Y
sRIYri2wsYTX2w0QgAQbof+M6f6emtog+66JHLqSAEetM8yeOZfJfo38dfpa6PQ3
GZRwNowm2p3QNsF8L+svpuEf3z1tNmYofjgP0izfkiwPAGHvIKPIzRgxi5agL/T6
EOOClYV2hfj/s2ZWRUeJPDejncpI4HYQNelKnTd9d7+MPIfitryFDQaHS95eMuW1
D9KrIeth0b0uC9wV/1rjUdSiBLpb4zXEw7f7luS8rNt6JtPo2BVbhIfBpNR3fvLy
bOm5d/HwvtgpMQOj6Bp3h8PcwPILgdZCJvrjeK+qgFEs60ieKnxSzlu1I21gr9oP
KOj6tfFqkmwQPAIOeri/OMOnFl+S6sMwsdDKAjTf/Jr2Qrz+GCTS2jI2kqEOIUfd
yMOeXc8rQWWqQNxvsVgsgmwl7ApyGRzzBYFcyMeUF57285CwhUxY+oq9aXuygDcl
qOI+AusmNGJy8UlFxiWrQFmvBy+HehofcfpOvaFm0huQd7gF6p6dDnSJk7jZjY1E
kKuT9pfXelRyVEzfApd6bac/2bwojI9RVFANejwuxlTcvEx4TEwS3Bc2ttIyvbaK
UoKSKu0lwdfx3WyJboIxhNYTHOXglyUahAdmles6KIaZfhhQKua6NLm/cXk2HC07
5kKFDL/xshnbkFcl3SaHfQzh2CRznqraDUw3Xb9P8iEGbIa3Ky+Yx80GVUvuKzmk
c9/pyG2FGs9SERStz2CIowTyUNopOgGaNdAOLE5BgPCFhBx/YuOLGHDcj2fGzv2u
HuM+0SfEq13JYsV2HbVKUunwSFIFx/ldA5pYLTZQfhoFiwIScrSdSIi5Hui/IyYt
MHBiGRAmSo0WvbVZOR4IhN00KCapkbc4TsuwR1yss/cjCKWMYCsKfWg8DjH+apIV
mgyu1RfDkncAkvoUFa7/hMicIIvEclB5HzQqnMXUFglhizfnVJsb7ff4Ma2j9yeX
ucovhrPw5pDwGPur+VMMeKGveEbrE7QmsSXsBWak/wwic8r/d/Q+o8DTZLwqRA+f
iuqdCuvpYs2JabvL+lA7PPxjOa9FOLNuV0yj6CaEuCp8hIQEcE4ny2lR7IbftDlc
DIKvCfkZ0Tr6w3pBYForznij0Mg0L6beWyxKicXA3oyK0qneuEYd/yXDvCaJtqMi
m6jYSZD5wqLKQPDuopY0SDeXH3roxrawqHlER5DldNcaM/ithlyZnf+paBy2gdGw
jyXxsyIhG1Yt657rP2SdqllnSRsKvqH9NVfwbLitf11AQoQKsT//cql/DIK1jO39
yj74Dj6ZM3kHwQV9Y9Y9aR2Oj/kUcTUfE73WgAvsj44Ry6ht+MSO02zB+4AdkLhe
1+sm937ZMzX62IwDm2WkOh+9AQVK2XUp5zDpTfLuzVHE4ozbHoqzW44LT472zR+O
UxHGLlNbPrkEvi3sjrIKBpjGqUmpsST0T9oUtDnRUtq+50iGSYZutvUfRVVZLCYs
oCbtqoH0dcCerQ8tgZTVrXlGpx7FG6iUpnH84bDE38EM+/Xr5KU9lU7tapQmiL60
V5r+nJtzwkXckr3LHvYFfaIhPKj7zNEQsmJGtNIRLEv3nKdaFWZBBeCptCxPKn1I
iEgi6rEMQ2UgcqGJ8NDVRjMvtgF4RFCJlXBLQQsauUwwSVYdmUj4QhRsDQAylMep
o5kYURLtc1nSFM9Iy+AFNJSycj2QFgrhDTlfBKCP4BsH4LMS+UU0MJ890MvGRbNV
B24gTSoUy8c/drrk9sxfWxsDfbwtoAGHxiRKJO6adqh5jP1f16NPZ9RN5qODLDKx
qWQ8d9LTnQ/u4E1lYBt4yhhgfLOIWI0q/YtV5fe8qKSNdppLLUhgueAmELm1iIh/
xxIXeD+tuQkFdb1+0TXADrwKqnu4zJqgzkSgSrKEJDWbZsZrcWG0TdL7e/TQxs44
cFhdW+ROo21bUaLDWZR1O/Ds19riFSVZkTFJ8KgJa8j3sIZuJQyXJkFVEODJL8i8
Ta/lCL0gg2gJm1AhaQ0E9gY6R1F6Lv8RDZcjqtq8MbOefuO8YIz3kIv6kys8/r9s
8iJR+R9vDTBd9LlghQ3TuW76sA9DHyDG6dtuLysz3g/pz8HPiImRV4+6Y1XXsuhE
d7MeYsNbgvCZF8rLyWbiyvN3xtf+2wiIsOBlJUHe7zYp25k+FDKVRrAMMu0apsGK
F7uNeRqOpYzh6/C2XcGi/VyxxStTdf4m3OAJqo7/dIUKjlt+JuiM8GZvlGR6gdRH
xnoc3VqwI0xwfb8c58JguIQUkwD/IIVOk0FvxY+52w/9fC7d0fZnSSklKajZTGdI
hdlAdot8h0F0o+5SH1z0qjBnqkQcnBw57caM3nHyBsF40XL8BTKydCvoyD/BM9z1
gkIY+9tgPrrgTc30pblUgEgRBoY86XIC2rlBPvPl4P1mvv0dQD15jkGTfWeKJI4/
C1V89y1bVlkG/H9c4iALZlfT7vT8Bbrz7JTjm5TJzaMVbxL9mHuE6AZxBPZkgjnK
A0kb0snG3mMesn9dqHjDmSs6mbceUxSEJnP4GrhgHmwv5RszEYhTHfjHop6F+/i5
Uqc73G2KPMd4eNBmmohhLcEGDYMCzZg/5zDQwdf6MwjvIJqJGhcRKuMBl5dspvLO
V5A5G/Rdr4CRoSpBbkWCLl4sy2pdq0UCc2NPETY0N9hEH8MpVDXigIAEZ6EMEcpc
ukgo/D+RLeEgRHLfgN61AT9LD0ADUhLrpfvfgIklNtpfSQHSM8skS03IIWcRq+hv
qORC6gjxv2+ehZG92FIvO9RCDe5eyItIiKXVZZVpysdA9vHKu30sdnd/wD/u6nfq
PkAO9Xn6pSwVui4Mb7rwcWo2b0KFvzrWhDW40LCbKMYcj6oRNAbzqSBY/yL7SRZ1
aD8BnJFEERNIb3u5H6WQ5kT3mOYgRfSlXs0Z58E8ey5/hIAdPJvPktChlqgjhVzx
7D2JeukPqKy2prmeJx50giUx4P6Wkoa2TWF6+cu+JodsNercwxtySkam+DsJv129
lhWsjGDPl+nbvpLB3ilwQA7UxM2aAuctbZ+rwLrnwpxyplEUuA7kW3fMZ3QeVg3S
9FWwRjIebYEd1fBQIXFNJglT5w63mphGXFfM1nQqS/6sA/vXGHzildESioIh+8Nv
q6gHhUhCT2sPj0Kk8YTd36BR/T+pgfUDWyatnZlK34fuJJgD8BADXoxxPc6bkWyI
NWk2hrw6Nak6JChj8cJqe1LfgQRzn4ofGECszy6jA8Viq4gOoX04myQeLP+p827Z
PU9zZhUtQwnFGXYWRaWcxxrJjHUV4DM+vPqOQeehsWUl3VTBLuo1u7sSuepGAH/u
2aHvyzKLLdttdvWg8woEyUeN43e0Omr+dvEFA92DfKPQQiXGEivhmfcod6tD6EE+
dVx/s4NZMekb0IN8M/UfrnKa75PFTR33f2Zf+LF79dgn3qJHfBwfudfFeaU1U6R+
wIUDNP6HJOUwW2e1ljwp2EQVIu+G5juPZssI+0lNpd2yX7p8/B+BQeTdtZOdZTT4
a2Q1KeKNU7ILsVcNiykdHu4Ikr9zi3cVtrucHXoaaWoZMyzENWeDfVqBf7plH2Ey
EtrhBPUPuzZQ8DUxbOotL8Bo05uTJTNzFAVnU7ja6F8sqCsnjAPB9CYgs4D6d8Fa
30TKQCV1aPMLTkTg1VXSbNOsADuDYa+bTmPSPNHT44hJZaSbMiVM8UUHLaE7zh5W
Z/qSdlzgcNbMeGHDknM4T0yP9u7Sj2o/3fe50GXnfvqIzL3Sd8lr9FG6WrDQoDpg
MtiVnXiy5jAHD0rbfBxcdGpcPdgeAR2H0ZNWJsifdP3cxlMcRaFLUFczcSB1Xs6u
iBOr7wkVPQqz4kcfvURBvsZzzCEcYF8MgW5rb7m1/Fw7wt7Okt2PeKwpVaTd97v7
DR9//wsXmSn9uqA0DHS3kWHAifgLwq4wXACjRW0G7Sbyf4lA6oRz6fvNUtW/XwBb
Gx8xVbA4vP/PCfcZHa3OydsQXFyXf2EVgP4fQKRtvFU4nWe2Wxm3An5XjPe4pxwi
/8tgRPg7xQnlOaX4EKsOvO+5DloSaawRvXlFA+nA76XHRbsohLz7yfaoDj0sN5Y6
tOkBXeIaItZcOP7i5eLLddaORfM9WbQ2HswDpjRmbZ+70+xGe+91uV2MEPT6Fqpt
yTGqHQImzei+vhPVs+sCEjasL+74osRrwGCe9Nmt1Ebv+xfMcMYqSOcmp2OuRZXO
hUcL+aZuVmkfh6MyhrTWPX2vQSZx1HWnvJKgQ91CAfsfywniKTyZgX+08LhEu/Nv
JibmzOjdYrSylcj2jOy/aYtSumHTvhIdSvCv3OD4hO8oRd8q90eH5P+ywZkrKZWa
jqzRGfIfw5mDXqX71E6v1I61MM1e6FJvzI/fR8RG4u1lQR+xeOCayVlOjEyDETnF
vE9VIkx3ti0qAYXbLJ82DhbTvClBAMpL+m65Ri3YNQOZMbS35F/yy2+FuPBExDEO
qX/RjyDEyepznO8HITbLUi5Ra2wuszvF5TsnGw+kYoTZvTAhJAh88nbQ32Saqk1n
GjASNaiAGjNxwEDxdqvPT1VyvvVQgjkcHG9j7ztrxm0ko8DZrdJ1oseZ1bkUGNOL
i2t8TsDJpkrFGZp13+Hr14zNSxjZ/IYQ0AfZc8WwHy0fQMs9FNPWbdz5NqhlXySs
Mubbpxs3PUqcEzZGo8QtUD49npvr9vnMHPdHyYSds1He5O0gdhC+jzLoGI1gbFD+
c7FmfK+wc3m4jikshyMFCSa2D/ttpo7+z+i0W4xLtA7wH60Tur3IA/pEC8xUOJkN
04OHLeR0mpTdh/HbvujQJSlSJWVUb882MndZyq/XdQORPDr7ybkIkBwYPYAbz8+o
BtDvlRnOY2EbEr60p960S+whh63NEW3X18twN/aDL688yBGvAMyBXOR65F3NfATj
1bG/UA7pxU8YpOjFIk6113eYdMuj60mQdLfXkjGJe7vjDCn7NOJcnqgVd67S0qU3
bkAcoYnRb4OFc0NySsUni6PIgB6XdEhdQ0SpETg/KjScIOu6plag6XPScTMXOfiQ
1mHEpnDjxQpWMOGMbcv1lSbKpzFPZofBNGfHW0scjsXqg1kVOWQs8nPDOkP87GrO
J8I94ByzAJcd4+VpCzP18Rfn6TNwQSmue0aUFWYgDoiluo35VPT1hxMVbnAyIZQz
2qbNHRE9i54T5BY2daqVzKSxir0Hb2QGRjC9+WXWxmUIxcgqwQQYT5RHTEKaIWXx
IZXDD0cnYZWBVqbMQ9bsA/C62pP6Gri4Myas9kYf3slNSPEVwzK2SS9XTih+pxLS
N77FLFo9aOmqvkEt/bcd0ZSbd333BcyuYk7PEoqbeRgNJZeAsjbvkXCNHHomIpLU
EMjwbCTldGRSm9aGKzb4QmWzZD2jCVqt1Hv0dY7LTeY1r3FAUllGoCwuFXIdRano
ylzaS3zsC2M7jDqe742Nusu2UubwBDtA2z/14nUKrT1Qyc8qkiyMisdusJfWbEU4
rM2CgneUkRWHkyBzVND/gnFgDa8IS9SCWTpalCg7Be9rHj9LHzEcxchxqhOXrQ+q
x2FecdqrXlzTEsvToihbhq4bBioHBTRKeJ0V3MfgT7bmyFlcCr128Z5ku/2cimFG
AleqRdSUIDHRNu7CFhOJeKZJ7r6gLS6oRiEQ/XXSOlVZaULY/KKArmo2IoDBvOOk
l2OpuQjq+Ct4wvhAyhFPtuirxQVw95DgXfEje55KGwn6KSLWE5zXnlrlcOrKke48
nDg5C+UonbXghuzJDIZomJNiiX99jh5dpO1vVD4uFom+01c0Hd8KDd6+77RwHm67
DJ8xI1+ife8mpjsNwHHimA76Z9K2czrDR30PfDKvWnfOIgQzEgkjPV5gmkgaI/WU
ZSvYDTWeawvOUDcZwg+LuBzTd2OViLi1ftO0UJcKsYIHwYTrN0fycv+9AfErp9Xn
nCxcni0YytN4pFhx982YPBEmobm2yt2kowlxmCQuwKOZ2MPt9RKN19+91+w9mlr/
bytrelE2PauS9iIzpXEFK4C9UnGRygZfvwJPUAxUfZss/ZkBlYH/QT8pMOE75w8X
ahUBfLmWso5b1WH4+HsnilfN7xlvLzhjEt6ZNC9UXU/EIi1AGlP6iZ2i3kkAYUDu
j2TSNZ1c+1CHnQVy8VFnWOt60hh/Z3nAIHK8V+acyLlUOm8t35Wwx/hkcSxnEP2V
jqcsd1NSo3TSNm5+ZIcttUl5H+HUJfzMBXgJtcOPrXRXI0p0+0ByibSgPheEodBB
0yz18Mr0Cfhv5nFzuR2KWqGWcY377vMpL5nIDcQmqa9fRgXYyYHARBDKSnEXlGFr
tJ/UmTpJsHq97LHHCK7BSMX5Q+S+tB/pTNmaYew/G4WDdp1q74g8bvo/Mw0evVOi
A3ej1cPWM3i6i8P40HFIHb16ZvNR6gZCRQ28MHxuzHFbBqU7DSqtCRbKwF8Fo8qd
DCsdsguUEFHSCaMkM7joClMGIdtcvEfF+rVRPqrT3oa4/FQOsJDZQImH5aZpnLDa
El+zlQ2RAThso8Cv1SUqZeFMqeapx0xwHnH+qG3PPBdpzotlvAUTUnmVIz/1d0Da
gFXk4yCrIS49BL1MJKiAlw4yTdcurkKzL5lUQOGuD9ZtWL6NLuydsbPZHJv88Ow8
/FnaFXKuQ4mLgKRjQhTgWrCRPaT8/rS364/Bq5QmlezFAwHjwAWEMPZ0NCneNgtF
2pmAYnKL++I65KXljYNvdLLQvMlGIAU2JTvBSj/BEzr9MjkRK1xpz9NPdUMJSyxf
J35o57fxL9OtJkiXHUVQSu9+uKnCEceFkWerKut+bGD2uEESPwTyUKuvWe+mKLpW
QCqSIcDTqROC9UkTRUuHGwwYnIj4LaQFJufedpc6w+ZuGJDxeWjLSX7pszbDvu5m
2SiQ0TKQQer+H4v8jr8FB8XQty+RKO79Lw0yWmtQ/EHKYNwJf8sUhdqXZCjTwSL8
J+rBEm/nCIZpKCcGYxdrRk3D0xFrqHiB2nA0exov0nQXrylOBD9M+EIqNRIisOhZ
oZpACxsB49Wz9ysvBnLkUIq1h2E4+swtJBlyO32mQ1GhPOrhvoc8wqBtk8D24Cx/
BHKmp8/IM71xN5iSHR9IOAQvYMPg4Evwjv/yw1CN0zlWt17Qr24+vHaXq+hEQ80F
0s4vk1NUcGWb0u+EA3Ah/A3AXR6Dywu21B9gBHr6BTcscqVqajon/46bEvTUTxed
0PoX0b5veEhsr8IRNSSgcEVn60IgUaf+P09V6gA96j2CJLrd7t325AAZNiLqGYPk
ybOp2UXb2E7ireKviN4iWdjpp5lyH7HFUEJ6VAA/nwRjdM5CpMGmIpKTDzRhPZYN
f+Kg4g0wDiM5biwVq/anKMG6nYXJgLfzJ8achstWVJND+vcr+L+0YYn/e+Nq4FW1
R2+Hl+ES1DB/EJ2ptVu0Jf7NVKKPVA+NXd1XPPAD72hmVtXWujoGO02LKRFaYAMS
wGo7jtxZq8pdlH7DtI2suZdRfAFUMMz8dqtN2VeZNe4OIBBJ8tezAxnZAlfAE0av
w6oEzurbDaHV1+VZ/oGHDYoURP1zMy9yLqHeGtERU8x1/b08lJV3KWIScbtsnG2b
5oVDbCMOJGUHS/YTgHP6yVxWON9x4jmp5MN4NsQIYAfqwCEswcfaXTYq5BpygAdL
03Zum3v6oTcSfcUKSZ6YhEcsOLTFHaR37Oq9qH7qTRxuJvamZSdRbyE7BLdzVCUH
BwQH98JjK/4oQvCFnER3DktGEAv/DTVz8YLBHzsXxRe9g86Pw5N7x2yCKdLTa1qm
g1yvNUK++4/+JnCT8Us7rpYR1y17PSndf9tLHpLRMbyDz11FdpK6ZmGJjZbmzb+e
VvG4axmtTtVq6abg26LmbFNdAeN03iMn5PrTu/Rs/gr7llw+Huv8uwn/6iSWqI1w
xUQYYLFiCdWrS2SgX7bT8usqRpJdxeDmLwydirDvyCduB3kDsipmnsiGTfFqHOmX
4u4CnBist2xVU/WVdAfJdGIHHQgJ0I7pVXneR+DV0joWQC4ZkrczLfpJOgh7Lr6u
ZySyRDR1nWWCh5Kb5h4KoYf4Kkj708ciO4Y/8hjHolf8r1G3kxsheF1V4OcdFGUX
mz++4FhZVgW6LXF71qHONxaApfzdFwKFhX6UXFRKXM1N0kxhtzZTPjkh/eawfDwG
vO/h8ljY/fs64XRvatUOtFNY014Sh8lDU7+zUoYbW+SYqs0jlu4hIuo6SSVpyx0A
dnD3xdPt28HGpOh9qijcYCTqqfQfXR79GALyeO2iGJx/tGk8mkBWjlO7SjiiYxwP
P4MWtJnP0aez9BNX6II0h6pDIK0jswRo28+kfW6V8wdghYQ+tYTSYDcwmpalU6Hy
M1f66EwpVG3Igth1zdSb8pJR2A+Yxi/PN1QppUQUlNJBT6SbvMUAXyf7FtTXUk0R
elwwVWIsRd3AqNzNkLDL8UgQ7ncfKKRP6bEx7cDBoQ7dtCbeYKuNMMj3anH3kKvo
rJdCPa7KoLOdRqsYaXD96VjiWS0Y/AghiDbkCZmDB6H829qEkVFon1WtANEuX5kl
0BuCni9h8K9dL1qjST5tlt27/Kk2z6hLF+l+AuFpJ/rkphLgZg0Hd7geq9uS29a5
qPRYMu1kT6cIWwF+oK20cdLpx2tvzaAfvSZawvdEKRtYhuTedIBS1J4Jk483p8oC
zEhLM3Ml089m/kiPKgAEuCdMIlmyQHQrQH6Kipd6L4uk2yiTEfH1nmRthjx/PnzM
5KgDWInvU7PtQfIXgtRQomAnCWEJA1gyR4/e74IYvJSSbThBH5ivEw3kXPIH55+L
ipcqlIso1lbEE0+whMHhHG17JmdMNPTyNo0/6UzvNgBCFdWnm4tqFBXeqWRn9QTd
4PFWIA09Y67ZMrj/RoG+bNftMLpg5jtNu1FCGKdmuBHxi7/rUGIPslnGepSUfp6r
KcabeY7JKQ5RJLq0+0K2AyqI8R3f3Lo4wZsP2+90DxTKHmEcmlQkPD9TYZMyH5BP
d1vLTzAJO6TwqRU5GFgw4yKoweWeQ5K0Ye5E0KRCzPs7XgEZwD/fpS8KhOJh1+mN
88nmnhmOQLzC1E3a4r+rA8f05CZ0Xwz6mb4r0WdmGzHBD8jSsdmRAMnY13vj708u
+a8qOhs4u/rVfM4wZQdYsgpvPdKMzoSFE2HJ0JWUYsACQcwUYfr3qIVgcY0pklI5
TOgNcIOtyvCYBhKrnlJj1yDwg+6x7X2eH2PC18PszufJTqTX2Z+sWNo6iA3E2pLB
Rv5pYUqjMd4e6zSwrmLukz1JhZgu4CKdLQEuyekPlNrSmQnuiPKtP7M8CrbSXDnA
bpJHTbrpxXf/yuZdZa0ZgxOvFeUV3ONGUzDz52i9lw5XYvDsmR+G8JUNjP8E4KSW
sgzKaMA3hdty5+evQ8B96TwSop8ob65d5CFciVli0OhqVnuQv6aAygXtDnX4fjSn
LLkJyuFoMJcwAdWg2DPw9GT+RQKjQmd5eRYeUk+r82N59MqoKEHJsLf8iHER9y05
m+HlXl+PNe6aBTgt0Xm/bZuulnk2ob5rJyVMTp1oSvFNU/MTX0efaAY0dfw+RDtg
IAyynczTLmC3yx2Al0/jwlcRd/HlJ7uMV4zwtrUNXVAKQrpAW5wOSWIoAuN5IUym
oRJ3qHmLvUyl0N9LAGBfuhNVg/6TuiBoix/26ANxfEz2y1f5BnoPeASBfmnLlckD
tCt2tzSMnuUd5IwUm7RhSJEoGMP5l9p094ws3gaFsbIy0HQM4DAG/E+MvkZ9+gzR
0hZSwR2XHAQ87WXKw9b10uwOUNSnEt/k5npGhgYXWbgJWJEHxLKiAXiD3euNbS5F
Kw6YIQG/Sr3Ud/6GSbN0uyN0ctpG4lu9ZBAEyynJzlXi/TYVzzenNEC/PFLLhTPE
IukFp7BUIEgItLGDSBH5dCpSuXjQcayE9MsEKPHxt41nnOafz1+JXA+N/8kDBsh0
2S7/3gwn92nipo2k5DpwTagw8UaBzm4oz/1vMvh8Adrb2e7bxZ5O9YXO0EpGt3xV
T09xzfJuUi1pCf4j8eRFy7fKVRn/a5TOGuX0jtI8YH6WYw2iSA06za2alz9cR2kS
qMaTHnd9G7sV4pc6w3qbOPu/ZtxTVzF14QrQhwpGqhr++vzbAZSaPMEx4B6A7Sss
l5O88ZRIxUXrMevRx/u6AI262c5cYu8RdUYGeTfG+xwEJBGy3tuGU3UphX5z5NzX
0qHLIzEEFIcvKLjbzMcWG1XkP3B7cxygyjjzkAY+X5rNlCyPl2mTnRUMivHkFCA9
kChSKbcNecvmz5zz8wb8rzJ6OmDZ5pISiagYIhHc/lKAZwOjCOgvQQLrhy1aoG+P
qjGpoavwkRHkwxwAxcQPKyhwlq7N9kBOJHHJMPbbmfSHn38bJyrPRGHryfu51Qah
hgqPGvNO6mA2u7sZws+BarJJ7OKKOduGxd3YLsxrg3vNn6iHqYOR+XjfzX2/iBBJ
JQT5iUmTul3hywvn9AukiiLhjHGal4Qdyc/xL54Aa/qBA/BtTK19mLye3nKx2OgX
11BfKLjFVVAmoWcbfub4ffooFswX+T6ydLftqTU/cEqd24xmNJVF2qXI2qi8+hG3
AKNmTfoMpaYgkfLdRqQq3sGz6ZzNn3K+WJ9hrVliD0yWBmoHkuMU/9HcRzq4c8zv
r+BET/NyGAG4AnG5kAUtPzwwSgspmGbUEE3pctI2OgXvnyU+CUfeBa0SYaj77CBn
aYX+cHw1ilKjM6PZeSBVpAjRVcYdvHuoj0RDMArkUqAd+c1OBymivr1oNTIe6wRk
hKWM0FFbkCV3xPd/RLWHioSQ7M6h1fYa3z8z3ueGODDQ69PnwNeN+9QhlyCpHF2f
TYT2dBZJVw8/a698Jb9gAmWpiGLhis7D6fVqBBlZdT5FXGzH5dZBSl3cMkASmn5F
m5ORTWIBAdGGftS25GwP9XxpWUiTHQASjDWlPqaqEDbvi4RZjXy1TJyaHmvMKlf8
LBI4/rwzisbJez4rBqCt8jmXCWh2N6cQhVqYKBK+FB8zMoy6UovPVFSwcLcNvJPU
w6YKYkfUbwcNvu3yhWIrmdtbBCMe8nENe03bWDjqHPNWRYHGIW+7PkzjUqxLrqxY
cUgJ6GbfEkE0FKlsbKSKTuYqqJUCkRxuJreAqI1CJ96N9qH/gj4/A+uxVNS2bBBi
TqMX59YwRASHUTB9b2z7yretbqwzsSieg4TUvQaXA0RY1oBxhUiohIsYJmEvYspv
M1eqT8Gsi5tn+tBdE9rJ3j0TK9szXHIFx+mN8c4hyZ9w87VnGMvhXeDsxXFEKphC
gePsJubMY8Y4xoSxvvIXx4xI+TASm97gJFjBx9vmy3MIryueWFoC3SJFeR2tfZNl
Rxi+iSg06qHvBqTAAKNc03RGTUXgXDwc0pCMa+1fhzzxQXWVEx7D04xavK18oPkZ
KsbYZhNPYxtPaI6N3tbsxXeRrHo+qTU+6w4eXLhmKCTIW9VrYGpH3G/y0DXaxqPK
CRR+AqH9+TRMMrp37QLwVnTlXwaU8U6pRoLldMXcltnqxeBPxDclgI0RzPSOBOXK
RRgVPKwK5V2lLB9nEwD+UAjymo8JlWuP5vVz4oNeRYyMMoWmpJmnLylp+s7BVR23
dyE1LI5hx/kOnU0YTwzK4TylqCDHJy7jaHpw7J2cCc/fboOQ/H+JrgjRvtMUimsA
bNNFkhQasL1pstxu9VbAnMEbcjEf52cZuyZwapMsnwV8PoyF0DubOR9gkWtmfH7a
toK23f1lb/0uUW5fXZbFuf1BwCO0I/sa2+XN8MbeKullOQMS2i1S9zPXLMv6ApvA
ppKderKSb+HeK8P+4pWRmtqbZ1sTnSqpGGisrAuMOnVGJu6zbWs6Dhrm6x8rxKYP
2zukqCnc2POlcmoivF1X3iA7fdLMbo4dfAwMty6DTugV+6VLJeIRsSSGBDBLrC9H
sdgUt7T5SqDEQi3BIAtaLwjb6JTwOzItN4m/YdaewLBt5COcgwVwKzLfL9VyVv7b
bLVZw2TLM4jsLFjx55E++ZjJmiep4qYs+y8ZbOkSDRDOKq3zP1iQv4ktSc4ot74q
+ZMoTBYP3745TJGsG2MJ4zzooNenLbkaM0xSrRu/zInwYijnSXq+5IVbzpQ4cn/R
Nr4xhqWMns1yj6FXMYT80eb7hqKmH4WGzVSSRMIyCsNit8GuX1gKphnhH+7Q4qvL
tx4xp89AuKo5dCe5lHErfF2rgd+NW58zN9UFfWfN9H5rcdfBGOs7Al5/NrgaInF6
RVhy4ubnw/MDJMye/Q/lFN/VzdhSDhfEy6H4wv7ssV5ifw+oK344dX/+7FSRoxBN
lOntdIF+V8Q9DVWQMYSZUG/xgEgP8T4aXtuW+j2WcPmVsS5F/VSMPoQV1RRpOupZ
1fGWESrm6KDrE1QhesqhdSIB5aKK9yf7yL3cJ9h9MatxzV1cxhZGmUtxfrrTSTRX
L/RsiTM9bZJeyFH4vTBIavV1q7rYk/IlA0ey8uUtu9baTqS6OLitCQDsCjsrZjrC
5Jeq+ribjxt7TtX2ikekeiyxPd/YzGrmvYpNdOilb7qkUbvFPsoPnQaQropDkqOp
u3+PlVsEs28rxA7AVwaCTIqkxXgmplWjNJ9LwqFTlnT8RZGVMiw0X3cwsNRPQqnM
iC1nQvZJNcHHFhSmvgII1+sZ2a2OGJIoA31aQ1mWqCjIBiuU79FZkPKMIiYOP1GE
e1xyU3LCOe498/Wy2TVDBqBhdOpvtEDRBlSFGj4NwchAmaXgVwi4AsR6kP6S6kOl
EWRotqVtUYMM5mT8PrX5594h9aOyzMNgkSB7KxohL/Tu2sa0S/72C4yoRmCJ6SnI
iH0wUQ7OT1G6/0BXTD9Xdw196vS/rDwcFAFZ8WGn714ipo5S/tP9Ujub4WJG45w1
a5guAnW/0FZCCI4ylBxmp7nzUtETydHLcNX+8x/C7nTWBDKPME6Pm9XMb0JLqunu
3GcZn6Klh8YWiIhNpkDSRId/UC0LzCmVKxY2lC3puJqgbMjtLhX4iM0J0SLXv3hF
QKKad5VJ6GAKyRGlUkUT7Wc4vzgymzgkzsPBrlU5aWtvdkUE2fgXpc/quY62/Ji5
fCpZ7u46P+7xDzlubGjI3bBpCyxbElI0TEdFcFLNePG3yITRTsCj80vEq2MFbTir
BHDvI9Azno6/z0CxtVm5b096fDIm7LEDAz+68CNph6G2LfboWOtgOjIV1ASDvHMf
ZBQXrQUpNwteJpb7JD32XdqhkcBsqwxI6DpjyCMr8IaNvuyDKUa3QHZjybCgMus4
NRVvcb0fcxdthvvSeHnrAqIckQAxrYmRzYIfPpQTZn/ddwF4lc6+i7EnfhgsfnIH
MCeC9HoVW59ooRQMsdAD5cfAuXp5I5wqZyi/M1aW5/6mVayjkcdQXdLWHVXD9bv1
xqu2Z3o4NL0UTQfh4ST1hQU4MzsB1ze1cQdDpJsIiR7wKqAVoojOeg1GQvw5eYNE
Y6p1IubpEde8dFnHjWx8dqgJHqvNaTnH/x815uQ9+PPBdmulzUrJWjg7WXtu9hGm
xw3t1mc0OL7abGC/3ipZv4Gvch+z3JmYR9re0CUQ65zOH+MleWXeh+TAXAgDMbZ6
omOoFVTMMTNUwnJ4mlkqUehMH2cVcfPq/T4qj7IQHVDUTDNrkG0i2jF+nyhhIShC
5ZwlMCB89ScVm5/wg1W1Cqy73TzZ1G80eGStZTZNXMQbQiI8Lbh1LJ/bszWOa4L9
s+kqPWB5h0zsjmk/8CChRkp5nBWVYc7VNH2wPZsqsCZMqKVYLAdss1oQ+yVy6Vds
0XTtIAFXdcLuUmw2EouwjzIkL7tvMhDqMuMzl/7gSCK7vnK264ZLwikNODqQN1SR
sYe5yInqCqgPjnlU5My9LaxlaNUw24MiSKWp7JraXFaBv6o1ppo3IqNl7oT8BSwA
/4IDAZPKgNpt+uPOhS6ps1COB+FJS/h86T7A7uKt5XMq3wgzg9pkZ9y2/PdioZ8b
T84NY59hIlxF78uMmD58Ofyakn/uscm4QZmI2bre5Yd2xEPWLTxmAuR21VJ4aX0/
Cl5u4w5mG2tkJD85bPzUfnUvhBAiOEDyXBhpu4AkgKlLEWvhKLwz7CrwJl0gcuKO
XOl1+Ood0DL5Bnj83ayqGaP3WQwwvWhtHOoOYHqnhkTaWiPOzDO1NkM7p99JW4Zx
x6CA/3bmCki7PqA3X+w13pgOgQwpzAupqTld/0nliil93SHWi8B4CEc5wB34ttT0
aiX/Oc2SE99xVFV/z/DR6BWlKRz2Fk5ypGHG+8l4XNYAtzNsq5mpdUcMu4BDwTV+
vVZzf9uj4adfQZwMaS1gNHH257M9ORh9clMWsXrWcJdDIYPAIskht81vc20+uBHm
d2Q6x7UTgKr/W+Y3EuGC036CzNhgdP62sx5cgIOBKLc/RRsAo/NDrjaYGaC2n8/D
ejEYCYWVSmwmtU/n2ISPq2W5kJLKyTm0OKgKDL4gjCSx50vsl5Y3ZdLfwW5T5TDF
aJIFCzFXpp0LpqsjjgCZOEF2HSiWmjiwCLfdxI7zw2FFcW5gtnD5LDiIV/EtAmRh
YQfaJ9QWOhG3sQXf6BgVMl8rrfo7oLy+U3wWjARcu5ygG5Y5HLrR5ZuEBYqG7mmk
efWvn6i2qlKTELHXiOZKVSUDgxccisjYytNBYLQhjnDZhtNm98sZQ4IAy/Yd1qjO
ZJLEzMEoQ9AlR+omQn839RMoSf1JMarOWtcLGU+XDiib5q4kBsorrlDG6fwwYTkW
PEs4mY60SlJsZpRzhpBayuQ2VoLPFsXuVRNn4CTkBtyChCRG5uboAzKsqT1DMvm7
0JemKyimpWfk9TaO2QD9zJ6YE6AOfvE8ilEXMlEE4mMq/0kF6tKOJUDPGxXUOFoV
3zSAzilmq7Vio0kljFw9RUkcc1p3gW9Y4cRqUMEEw2sbR/AMbhrL4BvXKLStN2jT
yzuQl/iyeIJh02a9uSZJA+5xNJIA3k4Fm3jV4hQhNickhe9bwE/cr7jxkLSj624u
kV8jyJLpF/tmf+WFfzMALNFUB9vDMeXBgQfTHA6KxlJaD6B+SMPxS8ozIM/r7Ps5
lLAtniu5butCEAOah2pZ1UZo3BqbbPg8fdvjMMQesz+IpZAdooXgfldkyHGJzCEV
ExjXicW0swYVrs0G/C7dlUOwUozWj4GwBMibsRUoY2mjo5QnEPqpluN72uOYo0df
df2b0eFan7B+uljdgUW9W3/puJlFW+CZB+9jPNwWl2RSZX3ODb76HZgrD49aR1EC
iY3VYG/ZyRlGEEg6d920h9i5Da1vyy+ILy9eU5RtGBZjCdW1xzTL1BMqCkoL1S6w
FAj8VEkDiZbCGGR9Dw+9DBxarT+IpzPYEep+cAoalN5f1KPTAJlRhaMjh/moZEOU
1zy69g0maW0WXlfrJeK1xWZM8jl2FOx/hq/ZHXGYuEkS2AqipOvwZh1XaWde8cjK
BGi6TlsjEWPMj8zjsHMkAZUd6uHS9OcszcLhex5XRjdzkxnUgSEuUFtUvhTXd5Sj
J9bjKuSkpdWyrSgX/K81UrrGLzsRis7CgVVci0bfP1wwPNYxrSotDtDpDF2zORJe
ir9BCVqAXwUI4P5/m/GCmQ6RZdWxWLTqmzU9FNSs/vGhDMWHNoslizwdTo3Ihcta
LtCKZT7U/5f5poD4X/KEndyk2UAui1RmeSnjDOfGlqaTT/HW+XBcS2JhXg89ULe+
9Yl7sglJCF+HEPa04r+KAxQ6e+3kewr1NtGxEukn16NCaHutngzYGSE4XhcTS8rW
Fio9v+JvBC9p69PnbOvllAflk0Yw4LKXZLfGKRrq++eMfNnJHlKStk+HNp0WAK/j
cqdvnB//P4DW4OtvjObzBdBpOJ7xkdLL1SNnQPfB0sgZIOZhLR1c+r/XBdzQz6ot
hUeg66oq1DMVyr6RjWT7UIrnnuCY0vu49FG3QZwoEY4RmymYT3vKV59OK7/kYOJk
v6w2EmbqwAnOGS4VJwcjS/mzx+U/CeTeBwKszJcG+PL5npLwQZnsqLI5dR4TtKvr
FOg0kVIWiYvWroNz4jpX4nmQt6vT6XxMo7ypt9WMNPV6LNXC7su9rJH3qR+kTjB0
4gB0k632myDKELxS9YHr+WPWy0cPY2dhatpfIYFirFaOP/zkaJMx+OiTcj1x7qQS
C7sCxtLyPzEiIAP+idsKoWI0IaTCe/W9k5nrkRYRyl2qWcaVx+uYJ/T8poAJo4F9
cJRC/jI4sdWILO206M5xyB91UCT9F/xKGmi9dnrGOED+MDr+ZH723ZQs+oz+8PV9
5umcawOnY0rAs02fcdavIWxdOWaP8NdASj82VqJK2/vPMdeX5Rg1aUdMATtynvdW
JTTyyLKtEwUfE9PmpK+VC4/nNy9MzVw6sZxSo7kMpKQsE7naZQzI7t8N0xoQXAHB
K/YU180FdOeNLe3y/cy2rh+kBZtQiK/5rT8+ElbY3yrOBmdwZttoKMz3f64ZEW50
wt61TrgAnSfauOcU+BjP3OKZw3b73QC8dTR+sOGTSRzT9h2NBU9CAepsPLOdpGjA
WhpxR7kAD7545tZGYhv73kgnx/U2SHmC/YBxJ9Sm2nl+SjDsVbUrxm5PvjTvDjUD
tyfnXfxtcFIR5ri7X/WPDVFr2dvaQ2aJBbpIu37X9US2gMLrUin+lIrLO+xIbEOV
fCwB2nzQj5aR1CcyLODBOjZcHnRB4jiMtRR1++VQ4wni2xNhLRfO3Xzk5s+Zbhny
OrQESFnlkAFeTUhNTBZbfFkIJT+Cg9xpT8mmXn4n8gZrey0I3jfcsgXvYKKeLx//
vTnNIBIjaP9eZIk+rxm1eLeGEa2wNI5FThijTsEW+sHrM1B3V6irTiS+u4GWOdJG
alM9PNVnLpcUdEmsb2uDVrdriR3qcIzdjF4TqUPWOTxj3DgI0Vn2LSzrKpHmJdxV
+HC8hdjYIPzgkLr+SYZKLX+r+XFHvn9OozkYUbB0H3sFa85+GGlKYfTdA3V2xi0s
pfcI0Omhy6T3jbUu0YyzylA9+CARV5w0RWU5RBD4Rv9OfH3PXL1LT6E0coui9BBf
4M4F86WPhxvDrcuLnnGr1XvOjzdBpDh52bQX4Os50FOb15FBOaEaAujkzuxcfmGA
H8dS7rReQh+LjnWS52C3xL35oEGqQPJ0dAmPRPQVEQpgQalVGRE05kzxBkQ1f6Qp
4pix4QhCMGV7Aoto2H8GM7xyialRxzz5iR9gTH98uVLYz7GGCb5/Z+wAHEyLX7ZX
6q6mo7NM+U4dXD4PCWjBzHoyfT/LP/hxYszZgZvKHJMVnxHAvWfdPt0gKDUVn7E0
O5LdNDCGWD1L1WFT+UV0oAkG/MgPTdfcG1Pbx+/YL7wEDrbYElq66ylMKJ7B1gOw
/lOhB0TeSPpT5Hqjs0g5zIhpaV/JkBZJsUpcgHw1/H76ifrhyLvR41uPyGiiHbT4
uEYF7iO+1zwGxgkck1RrAUnqg5Bvu9mDg1qUrLpIToRm5XVK2XTUYH7NpJxj55xZ
YBrhmq57BOdwN1bFVCqxNqZu9Gf26FQiaoQzFM2nuwU9TYqpxrRR7lnVGHafa5/T
PoJl4a4OPcHPayohItxtLd1JZxmUlYrTTI2nS4mS4BRPa8ztaxr0ylpcUfyZ8zDU
WxKsg8qIu+KK9fYsV0V2gte4oa+UGf4wx/NlHk0pHvsEmKCV3IWU+kmS7JOOO0yS
daf5PJyXn68pCiYJvEbWxjurD08nJnuSsHRdSckO27/RQPPMzKHt9BkP8/YxdAz+
tenCS0ZQ5bhtU/u62NxjH3oFlVtFOxF5BHKqvWbzbLC3jeH1O7e3EQ9NCqaKmIzO
C3Xh7miGMPqTz9T4e2XBZzP0LBRnPcrV0jcIZHSsELlQDco3FaJyper/QYKzSqDP
hziMDmk31Ea1CUDMxpdDxWzRVHYI4Hg+HTnVymN/BjvtpO7GnLn3Zn/br/kJQWy9
Ae9LuUFYrHgpUXDsgEojfLzZGG9yvMW6X2prIQwCSTdTbM/h95CRSGOterbN/e46
KqCdjvGObI14E3T9JHQkI0PSLA6ZKY4xhSNG1Hu3MxdpmXGtH3RGq6lKeWfDrYpG
N17w/F0gorMqKSNpFXhtrfYxW8swMbYWeTge+bmCdmOExLGd7tLipe+Tk9mrgaar
M73eYLOG8Xb/yqSFpls+RLapxSNs/HphJKDsmr/G8lkS8VYlgA7XA7mu/ms0hD1O
9RqfpPox7Q0I/U5RY3i00bW4/bd2hS3krhxjd30hzSNZcDOQdSR1sEpWL4QbVflM
8TrwJE6RroTz1FsXxmCxv3tZOXlbmadTnAZE0VqkWd/imB2m/dL8wbp6QOhAC+40
W3Zo0Jc5sWobcKeb0k7gSZM8mIj02vDhmnOu7c/saoSQHjS9MNWR9233TVjS/IYn
lE5ZMh/rrDESc2VaJ92yVxuVuUTSyC0ol30XJmwDuKr4D4LaKaoFixAoTbb47Ca4
WRcwPEupknJMGiY/3xKCSsVr28xAmJmFK4ZE1QDbhgfVHfRjkJ0IW0QLoKXnwlKC
yYcYNUG/EbMLnRwkgZGBpJzAzCsmiW5lTzPbD4APfNp3DlxeDhtHtvDfG8vzvDhi
BF34Pcs2W/6tywgeHeeYHcpjDRzZfugUblnEQxVRUant2Fr2xeeaCcF+qDJ27Qi8
jiOX06EvzWyd0Cy4IKqegv6r40gHUtEJsu+8vQ7kOOUPlioVYxaPIH7afdqA5ZC0
78ZhQ0mof1agggY3Cs1lSEyHcjBQZnSuh/p+dSw/xrBcEjkOOzFjpthq9pC9kacJ
8KmmWt5WHkEHdCYgkhxlRKfptPlnJO/H1gjsven8gJRaJhlQLVfUkGKob/+DAoha
PxyGMLUnOTeN0VhOpnO7AX4Oe9yiQvHF7n9lTUxM2++/R3uwgEe0LzQr66lOu2Ob
pWtDP2by6zaIX67u5QN/wFXajHLHQWyksg7bHHqTS0r8y7ukoyE0s0+Y8AKw9qHJ
I3SXH09abpDJwR7F2JtJPKVIollbOgmOwWLkIBonJwL8PQr9W0LmzUvyBeYyoOgs
mCMmYPajFmZMHfOBRc9eHSz0psBhQQ0IDtKf58aqeLQx+90Emx2Ev0iXtWGHjWRU
bf4DSPQfdaeoE/xEhO3ZAMIyMKEtTbXkgqu8m2x1vmbqzo8zMHY/18X76B8v748m
CdKom7o3U91eWqR9mWTRP/W5tZwVJ0TNZOUkq/sGG2Os9cbdZZsZ7bFEqngGWHeQ
oDDJl4d2SpUTei1qSdl3JXP2s6FILl6B8mCKjnV038CHx7ZR83M0emdB/DbU9l9W
SsrQ6LovfAQpB8rrU2Gtksu0AlrqHWBAhJt06XE5JAky/kTmKpHpYPvEKi/EH/ew
cOdsKKv5nA+Q++KK2WIG0wdkMqm4w1dup+pnQYShVwJnKvpW6vVHG9xtbjQJfGeS
btJy/zeJFlq7s6cVTDsN+zyFa8FjIbY0+aFDB5/fdL+OqntuCLCvTlQyLZE7AvR8
X/mPCFluJcglrPeqO5KCpgy9+4MX3/2wfTLWd80iUhJX6+/Xzld3CT/ZnC8VbTj5
hz9D4lEP6G/wd3n7RuDHspfuhxo84Is6mmGkKnwh0/nkeZVl1SiygEjrJ4NYkgL3
ikP7xi3reiotJkq+nvyJoe9D++LxleHfEIpnTON7wX2DCsiyCPFLAqbA1V3DdRvz
C09G7gWS5Qy7gU3t8E0hpNSFmhwaWWzJDrluVTz2v/KbEFHVbck34ilPuQzU0HLR
ZGFMj+vmWwMcBHQ07jd+wRFqWayIgWjfrcPR4m3SBCxDtBeniA6xeQmwoflgKSBQ
0daRR2aBnLjhFkvF8tloK+YeciZZ2382X/9A1wVNl67jpcUnWCFSN6C5VMZD/tEZ
KzDMUZPgnWFY3ETn1zM1Y5Wda6qj3zo0UgtGt9mj/M7t6renghXBnx3tQyEuQqPw
cpmqPiWF+xcdEIg2EtLeiFkjlh63RU6OFeFJoinOuWIb2fV/ltOxh8v0G7r1eX+C
6ax8SY66Ear+2sfAIVbge+7tqz03eaXBzOykbMCgrcQqQpUj+3eXpsOuxxyRxVMb
kYMyal/1gl9U1y3P05qCf627sHCK8IIrwzgS9Gd1tJnmpYLZX8qV+puvuCpuEAVs
GneI4qVB8dcccLvjtbTdovGO2HGKhvPZkDAwssbIC16nxfA6Ga1wIBSUzdOcJGG5
XAp4Mi1nAbiu5IS6dotG/3A35q7iKNWN/sHslxkboMijESp9j+nXQ76WxUSk7to2
V39YyYjtrSyQkziPKEi57MooQhY6ry78Z3NDjn4EfvDJ6nHQUt3bGvSHb52pcV0r
5jTIdnyAf0ZZqVUMgyHGTAc8m9rjW/EJZV94BBT7j264Q2EKaT+PNSt1/Aukyx7V
MavFEnizWbq11WV/uQCioIn1Ibi4l1c5JtbR4bww9rWRnUI3Sf+PsAy4IKtoJVqJ
1EZ+05h6PfquDyjRIQpmHInMKeXCwJO9+YHWdYVuiPsGlQmpWLzsDQgUzP0TRagJ
zR3+JKXcTdr19Ly/ErzO/nM8Re/15c+NvNgXynaIs/rLBxvRw08sgt3N9Iw7Y9Eb
h+RD6yqURnZ8x3W5JuNx6kjkWnQ6wY9ubU58s4qy7mNSDWTuEHyo4VV/gPKOo4Oq
uia+8wI3koWZGiHId3EF7WlUHId189FotACdGeFaOy6QihG3AbyB/vxEOpruw8rR
hmg0mR3jiAgXNHE/bg6jWOMUyKTE5pNwQvdT1WCZoc0YIikFtNDwLIPH8DzoIr46
g7fTtx0paN9kfGJAmEnsgp99Mlhg36tHH+AvTXfSCru+LzUIQRctKIP1EKnjgWWW
RV9DGSsWDVElIAduix4VA/b3FNCk67yalrFqmCGwuKtQDJam2lDewFKXnmXC4aA6
x5XAMBFb/hYvoXTIjE9XUaOShlXGD5CKENGyam/a2aZglb3GoZvc9WYxgrubMd0g
ylotsgwHGEdGH7mDOv26589L/lZ26vn+2MD1Cj3RFpdqkFMvGcgma4559Osfj+Ee
uXr8HZfyIp/rTRo8Ue7P+pSw+/+k1T6KjaYYF6jjGyRGXr9t6lOKIUOeCZXkGI1h
UL50rKxkhsnhBxVa/DRTve2eSIXvJIR5tOy5C34m2m8xHSLyrKvMhnSsm1emWDdg
JU6DtfAG8c1PmkN6UoBwCIbAusHstpC7gC8lHc5/EjcnRkkKo+kia/ZUcNDS07U/
4cL9mfv0bAJHqZJnwJPquHPBtGaFSRu0VCaSd5S9mH+sjxPIAydpo6tI6w3MYT1M
GbYCknp0/q/nsVhr+TcVU44YKQIb+eoomaeccKv+e4E+kUq+Ol1l8qEYBHCo9RCc
Vq9osEB3OPfIt6sXlNK/1ol4XhBA3MyUMtjgfjVPDlVWlwPjJGJs0hb5EeFaQkde
a6K8OIReJSeSz1T+KnDS1j4tmV/Mz/Yl0BQIe3pO/yrqaiGAJJ7ad0sj/DvT57My
iCinpY8gap3MJSycXiHWyT1WlQtSyGNu7FUB6llYU6dHZsFPhp/Q+SHDu60LNcZ5
rI2R8eDdkmn/owhmoYdxyhmEriKTDDk8jOeUaYB0RoKxqdh3WtT3CIKRk9r5RVGd
Pz5VhaBpwIsU+aDvC+snGuXfsAtTmxnd+DTb6qnDCyqkDV5+m/lXOU6t0kbAcbCf
gJepYaSC/f0YstilajJoL12oH32VN44N71yNvYi1wrVXihgZ3bAuUOq3oAmHwpsq
ppl2B+q+3XTXD+y+nElQLlkedVettE408cLUQGQNxZZWnQ36TcZrmi3VbAQa/VBl
PxmKAPg8ka+V7jC2bKePTk9+FK9U3nLyI6mvAV8ZqsgIfDeM7k4GtIukcZuh60n9
mJuWhmM1Z9GQCOoJAjX0/6wMoUVgjt5ID8lFwEEkBwKStRn+A+l6HcfdQutTZZaj
2TmKVYm/do/Bost9CCfVmcN2qLsGXMJEiub2+p6j3lgAqP/c+FOA14TGPBrsjaU/
bMbpm60010h2CIYmiqM1O8APC0GMdCQgIdqugjhDK1JzSIewyCZwax38qrHQWpv1
94gOshKtPLkRISCJVpaqw5fNexJBoGV+pnFhttxOM2byvc3h+kRQpA1ZdrHYwEAU
52L1XLkIevfmbseaQhrvsrmv7ewdj0fWHmOxs/l4raKRjVw3P1jLmslGmeKwDf2l
b5CajbDORNd0YGFwNFT69EFop6MZPgXCL+yCzqcC0F9OzeFpkQTw2+H3/V7DlJCy
2znSQt9fpZoypAOQoKh3vL6fhjwLqfUfnybNirhMO7pVJbm+OHNlgo/ZxvBKFuld
vhdD/XmhY92igbB6gShlaA12H24tPtHBHgADmpH2DyAY2FVWBG5TDDsdvwBK7VnY
tlc2A4O6m5yJEb7y4zIfcjopASsywxlY9idnDaSeUhw6VY+onMOJApvuJkmNh/UI
QxP5a60joIUzP0X0siTFJDph1nnffbLZP8sdX5xDwMoi/059ri/4mdRkowHM+HWI
ftIZB8fggQzzSmbClsa5UEpPfTzaxgWRle4AIc4zrbJDqME6bWWHd5RQCJPzSW8T
jrERh0+7tQj1EefQ5YGfK7re1mUZow7rJd20otKQLjhqNtrC6MIPyyJM8aLQWw6A
rSzmtrrw5Bf/9Y+s2Q2JU5p2NaSSduGFYQtJg+TensOQGNhomWv8GuO4OQmsXL+K
Hioz7lCtADRofm8DSi1i/76cgYqAgogF1dOhQOspSr7rhquA8h9Ff932Xmn87YVC
cH6HTU67IiUxAZNplU27qXdYSWbYGlknUOyw4VoKojcmiOvLm/kYIdzYzCmWeA5C
oB693XBpYF2RGkgMg6UY7TkTLUKT/Sgdhf83dqhQ7o7LXOwg9U7X30Y5Fa5dXyiu
e2qyZImdwCDuGKAEo7Slr8G51/iE5DBmm8QCrFMB6ObOn/Mr3rdZUOYu0DNJE4lT
no2K4eGp4J4Cq9JrOGzR9iyo8TV9Kcrc3m4EYKGmUWdBu/c/ezhhwTPeXva32elf
o2zgUn35jR1G++No4M20Wq+PhORYFYWhvK5njggchzaaQh2jtnvMbMAwct1f7WAc
wtnWNDUPvv1k3VUWyHsNEExdJAG/q+sP8F5sgXVAsQgmLX0HyqVimktKnbSLdKAN
sFA0WNkcco2wzdFYAzp8DXoj2jKS7IsxtlPrYZ5DvW0EULJbVTnr+PnVuGeDKg2H
v+Cx+lcIQbMi/biBlzbH3Ms3mw6bPz0zxW37lYnmCFY8wTOYDnalSEUfUM8K7c0p
XUlzu4BglNaJkHgOwci/4dErjmtYkhZUpODjYx5sCHSnbRSjtroCjoKJ3y1E+mON
6OpYmQtEUzWKwRcHVdRvK0xvINOHdgGENRdHTW6eG0v+INUy8uhFvK0LF2iJAtyV
dQ9a3UpHJZ322AOZ/r2PLFra6u5juad7H1UCT8Pwd1jOPdeW6qzu/pv95pxECEL8
DOOTh/Qp4I6p19YoPLIFKI8krzX0h0wXWpzHJP5i7N2u+ArBmq5HFqujIgfsgE5v
PUwEWFJz+q0ntronNoB35PQ3VulQd38ePvVClDSw+F/CzAO8kDUppEFB8tSDTwlV
XEDHU9+CZ64RhTVgQSXRwJUD9zxXuC/egEXqD2GBYSiP6KBaOASVGFsx5eXjzmrZ
kJuQ98G4JCWiCAGUimQSXqrpHRcuAce2OcLlr5uhD4pBY9ip56cK/c5JJhxYMp2v
zi9wnCGg4Ermd+jEVk1nZrCcrAtGlF36y029+zFrleQtprdaDniy+1t0xlaRoMzF
Kc/Gahb2W4EvQGMnTxIZBxS16YKY4NGf3bxrL0Kxr+9iUS8FXd6kUcb654ZFi/Qk
evZRl9t5OGmSirNtTd//b4T8rRIzTn8mA81BX8yacxgYpKGPhFloUAgwyE+MguaX
foBlnRFoeFgk2yHGrf2BxcQkKqi8fIJKgGoEJLORSoZYyc1qhI3zKn/aCdFCOSCJ
xIqLnsd4NAFxQ7przsiLrpjVlIXE55klHMw0T4uX6hbCx+lD71KTt1zKY8RQlIZt
QHeeY+6snJM7Ct/ZJGp7ux2Xw2zox7LMGXtTFNbLJw74f9NKHWi+Ef0TKPx0Alw8
UuUJnZfguTlDpQoZ6++jkFHR88o1e/WSbSsIpr2kmNRjzA3IyY6j90HBJpdToF20
XyBkre/zBce4nXQ/sZfAPS2v/++4OCVn/+Rp8SemPK7ssGDCeVasMAZSIW70nsxl
S7y1xL+2snegHHKz2JHtzHXhQq7m7k2o5RbTnojCm8WZMZaNCq0QAIAPckTBL9OM
dD8rrMCP3ugIkPsXLJK7Ie/6sJj+5Qu3MubxjNZ5AQZdUTaQeyBniqs+gQfHHZIr
fiM8G6eNRpsobaVOJ5wZ9ex+cSodwjKGOQbSzsR6vt/m2LM0iAdGB4B2/NCem+Mq
Cnv4UnrcqcO5IUNvkQoCkmy2+mEYXUPOEFBmg2xfUZuEs6APfidQ0FT3ak9JTvK3
Wr2BrnDD9lj3bhmJaBbkLcyG/ME4seFMB9kXaDiA34PvQC3QXvYthWpxuar/X17E
68siVcLZcTgtJh1WIbLGam3fT9jx9O1IyxujZcS+fG5zdVITqPbZzB/4f+DASrFh
nIpKNuSp8rvPRzflbqeYEdL4k3HCrNW4WQzI/MT3pGFmPlnR3nhNSvfl0NsRPml1
c6fOuHy4xovdf2ZqxPq1coK0aRy79toYf6vhUVXbObH9qOvE5ABlhSB44Ovsml7/
qk4bkf+uDFtQNgC2xXU23At8eqJmaNiWebYGBWWj8KKQSMPJQUbN9GVRqg/i+YmX
65lfC2kws4YwvvTE79RODecTiZYploniBTGsxtHpb3HDO/wpI/zqdPYEruAKoM0f
NHddxGp++eDmzMw4TCgwZPqd4wJba/vrg8qDXcEHSIhNVsIkPrdxvNoCsp3GJaqs
D8wL8T33ubraqWR4ozmcEeka+60xV67UjCzLSCfBx7ZkEJYQGa6xLLWJzoLXtXKv
XUTMiNRiRnQ5DCSdewqjTRe3GGWioMJQWyd9zbXpRO/vHg8Hdz79WzxCmxeGMcGl
gK80hMVWCyBazz8HO1mvJokkWdnaHj9mMLQ1fRtj+Ec7O5aFzvXCZk+Ik4EepnfZ
W6cPuGcxq3EiO+JDyIijz57k0RGIVacF5VkUqQq/3mJZV6jcyw6i8Q9y3h2yKHvU
58xYPCOsGg3i1+C7e1hU/xYjksxff9y7JVKo2XgfTCne3Jqc+zhh4NZEhUX3hBya
mIEX2AqU8nYErCQU7AX123B6lt1B8KoEDW6IAxyBBkwLSpnQ3WAfqF7YpLBCOqZb
H1Nb+Ekx5BlwluKUVTg4qyzfpOfXQLj0u/4NJfK4fT9hTX1HqXqnnXLgvwavavCl
qVM8j+vDZ6frC+0hcrU1sjkhR46fuh0BWWjA44s9M2XaabMDPjae9UEfOFyZVM/H
bYNx3V48zRGKV8b9gsyQXVUWURMp5oiFnsg2fI8wv+Zu+eZO9eJiYGcyG1S7jXh4
f5NI24oP6u29dxszdqaMHsLo27O0KPI2MdAX9RTIE+iyQbk9omh6DChb5Q7bG077
hEQvctM5WiSNy2o8imGUU+krEKPN8Cav6+JrwXHxvNNGE6d5fFdQNVsjhFg4EC3I
6ONWFzSl7IFpVwCGgGX/U7UhHqmJueCrtyKDrAWag8ThbM2vRxRtFmemzp4AxzJZ
IKLQkC8H7TLe8jSA8sekgjFXZem9QzMzQ2eMOjOs2woOiKnbKqSABdxrqZ30FwW2
bpArmJI53o9A9r/aV96NtbHKBy0kkbvXCBnVepgwELb5vJwcy48DHCwn9ypXoW2A
Tn5QpqdVolCGwPBSmniUzQOO9fD+li3fpnOnaNDxCjh0SCrumWkqyY8+n9n1tx5w
1BTOEH+y44GwiHFuIvnoM5hCSiwTk1zxr6EEzBnyYsH+fCt7oW58xv4+8W53ErRo
1pf88NfzgKpzBmI6ZlC/GJb+7orkf3FKTmWd7hoObB/HVkv85PKlq2hj3N1e4kja
b4yBfC7AfGU3e4cm0HOuNwy0UEMl5lsRpMW0dvPOhP2brj+R+Mn+pc6qOU1WFR7O
NZyBhhjrsb7Ijso2zJPCCxf8ocTPqK3HayV/+qDds9qaFMAUwN7dPWbum0Kt61DO
c4EKzMf3gtfuanlNIK43Gae1J2R9Uj1xRnTVg1M7S7YGFYSrJG5/CQw2ajr4Fl2a
g8nBd7ixWTP7sMPcG+Lw4p5IHv936Ua+P39Z9fuRxInMbbRezYEsVxhgnshHzo/G
YVME1eohHVqh03mCv766wRD8zjUWD+iOjwtNmeD90mgV+l9rwMh9vvEamd7scRiG
jBuTZrlJm//4zdVYnb7snTuy/FSUQGfjWswiTUe4aJ+u96W0mKcD61ejOkDPr+EO
WXXQahhxvissSaUOZnHKX50qjtyzwsDOBVf9Di1aou2K0qLUVuWfVfQIfPsb2WYh
F9QFQfyVlxCURR8h00/+y2FoTQsU0hyhKH35mjh4HUAUFaGSP2KCeu+9265dBoAG
tkc9A0dlKxk5qvP1ODCBjn/r+yv2WGJkl4jcpI5Uk/4GV74v6MWLdbrLYs5g1ecK
Byzy/gvuhYFf5jNffn//f4K/OzyEROagZ+1qskgV8fOSH3Ox7SP9BPJNDbrcAG9f
FKgoArzirQ/ylPg4jvn9nMZR6udyfgeREtfKeWA9Pf7jOrY8F1pWg8LN8QFThHfn
2vnM1uFlRO4MhfAh5mgrqClNVMOMqRgIpH7MXVjk15WHKxb8nejmkbvT3IPkVL0Y
4/e8zS1jQewGbgZtRRqec85C9uYhoILUC4vZyNwDeZ7KsHsW2TGSmFwM9QCuQQ3t
Koxinc/kY8+3uHxYzaHak2djH6q1rUfaKS8OBUtk//p6B5UZ0V4IHp6bd2+wt2Og
TlPFhFkDqcVDgr/p0J4+/gEbfptlbT7hGmeuwlr79WAY/ElCqmJ6YMxe1B9kxjDw
0XFv7MIbJZH9Yn80+jIA947cItZB35KsZ7+GZ3JGY+AjgZpGKw0PIcg6T5GNK/fw
DozxlH/IEAXfOC/XvVq3d7hQgCnqX8onSeooQIGwpgdYh/r+MrInqmFS5SGnW5Zn
Uffz3Aad+IUmqbLS2w54vtUs2mDITE3hEQCDXWGZ7ehVpi+Rhi7fWO+M7UipldMM
ZQn7rIy0iQSoaaAWsRQMQAmvR0GqIW3+PPh3R4PSVuEy/s08yxmhHY+cXpfY024V
oaGmFtwqmW67QddNyL7TTHjxw7FvYInDIIeZcw325ib/zLN6uTZ2Csl6GlLkEp4P
L88aXXavFVpKZxwXGk9bqfelcNgIpRHWLIjLNhUJUbj9anBLvHgYXglugQ/fw5G8
ds8CH8R0u9C7mLH6xV9TjNBDAP0zhmIQOh5XZBa4omRk+coLvmG9eT+8MEcFrUYo
4zQr3fsoKBWyTWdGitRRz5JVs7tyxRtiQVkXSXUWM3E0L1zAv6OlSrAbRpR2ouLr
ZMSR7br/XW1d7sh2gBRYcj0EUy7bIa3Ak6zdmYUwv3LxiakxlNHUoK2lyUA/iI0n
VnlTpmtOqy0xgFG6g+pHAq0Y+6lEMnRtFfxB+DtRxAOANO8Ef6Y0OSYszDjj1vVV
U8+gAWgX6x8rLEdoTRQJaq2W9eY+RVKDizIXDmxWJjMLU2rJyVpOjxH1D6ykl9DK
SkwRJw2tKeyEFxewLmai2xRJLFSubFIAY3NFzx7dZewnA+HtoLeNxvf1486h+HSi
KYpSAssn8poty7+axER2lorREds2ZqwTHiTlK7u+DFn7BGs0Qe6wzXoBscK5tD+e
LzqdIhL4St/l3MT9DZTTwFaI5Ol1TXIOSUsf1Mg9/AOkI+EsLE+3GdJp4ZpLN2Tr
S67SBtd9zSX1JP8qLIcmL4GSbuvCW2ni9flCAW4DZd9k6GdX8zf99mVqQ/ULj6+G
A+pAURrgPy5bVtuj7ZmwdNsTsRYQU9E+i59kaF1ASP1YBROIv/VjHNKSB9nwy903
HHQRkFwoHbxT9DC/RqFrQzzOe/0Y6e1DARSWs5D4IVYVY5TN0iutBaxf4GdgF77Z
EB/KGhtZDm/ZFlQ/AGMOuqW+Il8FpZS85NLXCT8Uysip61/6vgyQ41ckKAek+4K/
C8ubz84sdtNWauevnu2S+uTGzJ6k8oeiNVtmz9wSIhC7ofe45nsf+5i7SxIZD/+a
6rHx83XBjwwR0s/xnR+IMWAQhtpYxaJkYcUb9Y1qCXcga7u53vO27xyFTAUNz+hZ
ku1NTPqm/NKTrXJlWPE/T5AFpg6o8g9N0gip56TqvuTR6vvidFRH3R7wSl6RW3dU
tfVDeu0WVbI5RL9S0XYPasUIEA4s4PMCDbK03PeFk/uk8WKlHKF8ijIcqLvCwqeQ
G4sBgokJPixy1peNvDAhrG5HuUeiuvggnZC2o8e2RdQLvMw7IhnI6Na3D+iBgvN1
UpARHz8+qmymfSamQUnEvD/iPkhLwS0VEmjqK7gE8X72F13Rz1Vw5ZfkR2TPTuR+
njN/5QbvoT8gRvev5lnPUt1jTBxtitW9bpWqvij4YEUn0AsFcxv6HtN7JDrDpx/s
O0+9K4K23iTyTXg+81/M37LwHVMTpGOh5vZTcmrbS4HDLIrN6/Mi+j/ysNjC1mAT
RommjdSpG+2YIrMSSZUVEZwn3XmlwYN/oppnCEich/r/lMnsRiivaHguR6DpaSpH
1j4ppf7qSs9wDU1JOrRncF9ZbRA87AEmbwbqs6IRjFPfIWCAO/vytrcEFGH5XHXS
rv7m2G2Yqz98WYHkHly0BWNKixJJCkkVFCdq6JG40JgkNpKPjIk8EsyUbrYyvFN0
afBLyrXCd0LtXsmzkksHoFhtkBiqlO/LZTZ8ySDC+HB99QsvRCszmLFqZHX2YRLE
TICv2lMYoU8syvij8hUNQfp0BwSPChmxyCz1jtqMEMhcPhRdyTDfK5hYPbaPUsH0
0AX/MmTWcbFsAp+ESBsWeuSBZebdds7sYvogCY/9ABMxcyQXzjy8KxB8C+EnI2de
qUCbLXlzuLNMY2VDmWs5kGDgDssDVFJlncvWKRJfAiuDvd+6+ZJIxOQgYjPjoBvZ
nWw98rklKlJ8tYsMj1pip7tOdxDpy/iYo3u8eanP7mWmVdZIh1eoaZlauhQg18v6
Y+LbDnbNxpU/+p4l8wZl7pAWgQpW3VzA94Bn3NW7ZQHWeujPP1kRPUE29xqw8upS
e5MJ8/Qq0lcapTNQDrllSlniIvZyeU+HImKXOs1ysbSX3LRxmeZR3pVTpGpDeeNb
Hh7spAL4UcPA0IWWyFX96U6kfZA0QB13spjuIDRe4gogPpSNKHdMVWrZVLS97ctb
5lT5ERNOu/JIe3meIEUvTT1hNJhr7S+9u8lKhKGn0SyRQHqPhAZFjkQUgTjq/a3n
9E0AE7ToDHrgH/AnXdiu+sy796eEJ5rVLuS0tPR33CIPt3lMr1ZHOv54q8w4lAIo
L2bE8ApKa9MzKtoyFvcdj3JEt5G5kIk601HSoUzXg2ZevsmHxNg1OGoGdxBBEFoF
g+ZAs6gzyPFURtkgpcGynPyECnyNFzE1u4rCz5qgiVsc+ulEUZTFN2AjItEhsbjc
QR/8SB3uECBuxvfKYUIMOPB0GQ42YcPUbIvLbZM6p6jeEy9A5sO9lmWL8D0rAvHR
SMbi/dwNQ/TeB1oCEivUEi2qpJ0jcf0m1BNXL8EZ8l9LDsH4DM2XYHJW6vuQUR5k
LeJHKIZhEB7lSGZBJZqugLixE2QBH74QWAxtug4+k9c7Tjf3gEr//zk8xRw0HX1T
QI8RIeklJDA3WVIfkZ5LUxiZ2LyLeENkXJRfarjMIVp1vqQF/fwXk07Gf8RAxVHg
AgmtL5s9YlLPGnAEuksfF8zTTdiKYAS7uqzAJNnrw0A8smhxC63CwWkrZQ3ahF32
DbjmCoLSrbPnAkQo/iSuxgzRUcavfw+2E6xV3Eyfa7f8h2pqLMkbrZxN2e9x3y4e
YFVru9GJjz28me3YtTLizszJ5wLHYb+A/a0wm5vmIEquWoBgJoDbax8dgg8XW76r
sJMxVC41IlGeIrM4v81222Z9rqz7oJVsNZdMLlt9x1V7GRSC1vtdXCYFvq39Wx57
kZxR9z3/MjgijpPuk0HR9aE6t1Ino4PPSrqj1hmvUYtsy+yaBgcMkyJzE6yh7u+a
zZB5nAPudLqoA4GQVmnRNqwwO7VzDnUk7whR+6zagZn4NO1jHaOeS7zfgoT773DE
UgoHVxGzKi/IIeYaU/aJiJRznwGnJ7cPiX1VgFOevM9G9/vy1wwRT6iQTQC9Brpv
VPpY3rkXgAipzRSS5vsxjOyBWfK6FrLdXnUjz08Ed4ay8X/qRD+JSqTkrY97vM+z
v5A8k3EydYf7ik3h/bjT06G85JD82PkcjGja0afAs/+IOREy0vqCTT7CphWn+0mc
qYa1zqA7VV8c5OIrQvc0mG3dYOx0VxWjDuRwazPdmfQwf2bmXUnm64wvYmh3FAN8
pAFgHIibCZ6O1j3jzcDpCG0FQLGYqgx9aCC9LnYEb3c78Z/iwhci9JnRk+qoqI3y
oBVY21vE4932jAFzya+RjL1yomOVt4CAroVaQ3DdNYskBHqflI9HWk+8u0QrIBki
QXJRf+MjuzDYmAVnT2b/DhG7384/F6/yk3AzDnoSIh+avWaY9YLCbr20w+wAU+2m
+210P0MceLcOKF+KSe9piaN620QnQUt576Sw4V1SZ8IQq35BUdauuNzAg+L1WFfQ
LpVJGeHYMBuzNdsF+lz/vJpOHi07dOaLHO47XCbs9sLhPI0y0PCCqeLqqBXuBio5
32A/e/35jpFludp48Wwu+rAt6ZI+zlo4fFCNRrtDqFLuXbi8y9f1mFMWUhYiB8xf
lFIyfIjhdfvgggLbonUyxk1TcIc3aqyP1caRYeXYOjvDT8qyD2Hzhb7MLGWVcQJV
8CpdMMgHYSjXjJvWrvkqBOONXmMaeVnDX3Cgn8Yag2DjQHh7ggV0jxEAPILj2cwz
bNQ/WdWQkcj9eSTNUP3T1eWNUxwEyQstR1xuAKWeBHFb0NIl1nNQ2hK2fCOWPgIy
rS9Jpq3Epg1l/Nq67kUnH5wziiO6dQL52a7g0gd6c0WXkh4Xq7JkL6nFv+t5hg5r
rGnbESs0otcT7Lf7oTALmml0mzceo0k/ABAXkZsj6oLTPe7a4Zi/MsEgqWNmCM/H
Kb5mmYSIGhY7JlDEeEsECNldPWkT3OdWvMM/SX1UFj2sJeXI95Nx77G9OWDTrQma
ahPEuLCvnZ+N7Jz2xSeTpUk9/AgwJA7/WUe/SGIaPpn8L9oK4fNt+LyCGKU1SEpS
P3z598wm5UPdiQMG5pN9nX1finyxsC8HerbThbzHiO0svp3l3Kzr9sretdu4ShyY
SgBxOxrucRozY/Qzj39aQA6VmFOJ8C8X24j6zEVkrkg2u+YtfQCh25cB9gkepyc7
0KibKo3dRsEJxy3mGRfudH5BJUm2gm4qe8XIUfISPhStklw2VeYkFKPibb4eITWw
pMdL07UfWWsN7jjKnnxUL5UmV+tfrPkIY1PTC/ZZJ9xTwqSXWCQOvb3/4YQueX0F
5DZAbpq4ZrWe8SKoAiQ6KMFVibfsAAxBc+Y8029ok1Jer/QYtKvnOo/vaZXiQtIR
dFQ9gse5+Jr5LdmZ7t6NRZ2VkdnDeQfA5+xNhgQPc4Q2hRXhjt++ZTvrt5kPglP1
cXl4XGvT+8O0Dp5CCMHxJ1Cna3Rk+yxIBt0RK/MrdUY/n/WOD0aqrLNA6vxJG22X
2Y6qr86c1FPG72XOzyvWFAY57dmqn+p3jfQ1o1Eo6EIFPoRpEIPyEG2XGwsGrshl
Q07JdD3LOx4ET2d4kkD6kYaqLb3cLRhEQ8B0yDo87NrRxRs0PZIxI4uWrHt4Ph1E
1DLfMYhJeziXqP+L9jotT2SToQrBBHSRCWbBvZWgj4kR8o2lbkfKdYrnfMpE3F4W
1RvYibwiffrtNZSCx/zs/9QDgzASyu+eog7aOZjnXu7sWrqlQKpjs6wXZ9jClH2A
aEZtxVVKf2JWraSjGG70WBTHrtXmIZshxyQncyVYb73aXtmYALF1ASLR9cbpL+xM
WewHsiTCyVkDL1ptMmPvfnOYZw63Q4fJnoCpFsPZugx6QXpIxjyYDlb6DRUmIsYU
9S2B92RlIwHdb452caKgqSXZFvpmCL043AhaDPFaQpSdIsJVQvYBalYJhiUEzSkR
Uhr0YeJOAJGE76hvcgo5mSOcGOr/Stn+RTsqk+MfssW2NvU1hUW7CkcwNY+iT+3P
NlIsHYESacjGAdhVe/cWJHrSVwFWRcy/yM8F3FuJ1RLpRuZDbhgs1Zj+hYuEnaS8
cOQwVSbp01kc/rmhSXegWXEMXkFYB15T+sliZz8HPXcZ9KM6YN8LGOQISmPVi8yc
u7d1/nnEqAzK/PokZpzpHpWD6tNe1S8izdXQWDVcOAbnuJBGx/hUtB8b/mreEoTv
ADUICh3rWYyhuUZLUT90cz3DaxNAMnZVLZBj7HQoD35BYQg/dyY1x/K7Fh6nWSgD
+dSXOEVT2n7E0Tfgcg5z+wMGa/pus8yWwSJeytCFRb1+L9x0LSxbJmEVm4WlDApz
cjN4eFOiuuzpxtypvxFLKgrgIPskHE8Vn9x5NefYDoFguInkkGskyx+m81YxNi+F
S7aPVo7pd/ceX2kHPc5DFr2CNMbV8ZxNDgHhDizu4/oLmS0zDvZb4Yc1y93N4Ljf
YTekcMOL8Bg8J839ZP/5V9PffyKkt/nhoTvmGEndMe8Z4eqO+1I+q4bCLX7GXq0u
KoSID/POasr/95+RyrwpDdjIPMWZDvXVQEK7F1oxdEXLHD0KHLvKB1Suudo4nxO/
JoR6Rgaffjg13f9XxIoyozPP8tpc58BAc4WStiHlANNKDNwbyssWKtYh9PaxEbk1
NTQcLzj9cH7gJ0GQGu834/vZbsgoym1PQc4/L0eHxZQUViI9P7fJyKe26jjO7u3d
WS5xVlr3jUR9/DY6HjbIa7clUwgVDZc1vWUyvMcMSqqUPNorXp8RZw/sLyICUZ4u
+up8JxOMLLApTZE8olN5YEfYHl2xix8Tg3Eig49yatOQcgmt5dp6YZHlPkhCbou5
sWU4DN+JCHYk9xT0XPbM+c/m/qblRVjfpZN2xl7Cnj8LfKi1ZxwWp04aZkx6N6Iu
VgDx/mrXhimap0lZAT5yE3hbwTz0vBAcsAM2sQ4mzCVdxRwLaLncAtLk1N3nToR7
g/G5XB4MwRxwlCwZMS1ZHfUCWsjFI9MJnZ7G5mkt+L3yt+cy+2BPvqoBt/64ungB
2iuTqMVBfragDVHXWRagWGgyBtrH1MI6biJOPz2XUJsui1Kz3F6ceDih6fvLWLhl
Kwq0NOzmyO/W3dcUqT6xMPZstmzltiLOXiPSgLS4SFouMsbRyHMiH4fKYWC/trb0
0GUBAQRusWxOXUwMK5gYu9+Mt7VkXp11P58GPZTVQoOdTCG+lo897zt2UxdfsFD0
pX1awjf4UE1ejPL3nzR62Ty684ySxXfdzW3Gc8c6W+9p19g7uJ+UXljhseX4g7+y
BlWwm8WR7E86lVrbIJaeY1MT+Ry6ZhntF+bo5PJsEGubfbD75eke0D8BYMsG9psq
vhuNhtqPs3/uTi/CNz4py1MfA0qllSzqXvTx31oIb96hlT9rx1doEKbEPTBDPNKK
dX+UChtA39oiBqqMVL8osnqNTR7Tf+MDUnaoxIMMD8WpLdgk8p/cw9lwlTl0zRlY
c4QaLBeZ5skdZhFZB8WoeVrM4BvyGJPcRK0Qu2s8TmgAKMvucIdwXtIjncnQRmEa
/srsoYyMRxM7O1cbptSPFJ/Tzx7iogJbFYQsdWTPFYfCnavSy3p6Z+GgSTAQ8Tuq
SSiJbBCCwmMR0i9bQWxA3GSOlxBj3U30i/myapPto2I6Fes0rgTQIez0CmwO+8O3
FN7z7A1wZGN9ijHfuHL3XVLzkbTfHfPTVRZTaXHjwxhZ8U4++bUQrLcdXMZX16Yp
nb0uKHkG8+1caA6BM3WPKINkGSjqV/AfzQ9ZT82ezxIVpcHH1gdZjkaO5kfjPHd+
e0II6kIUgrycQiw1yDUc0b2x8QDZno8mecXakp8xrjW4+N0BSz1VNHUzjhmcTW7b
sQtU0bLLLqdWLju07Sy6JU5nPsBH6dfGo7fnPYu18sFxZqX1r5R3lXyk8SEh8N0O
bw3ZxQxr+S0joQ51Q1A+j+BKw/1lM75EHn6fiSW9PAknSKkIbmry1Y5fFw9+jop9
/S8o33V+JRNMFJ/WkWz8FchR9I6/sDcDJZTP58v78TomIsMUvButOKks6zNDkwWH
aKMVEKXpK+knid9+DMQW0g5JmjtzY0nW4PUsVXVHToGU3gaY0sBDcl4sm+wCPFql
EqSgpi4rBhai9dT9u/6I9adzIhSBAIRDmiwswQvN0BTtK/rTskkWQk2UON2TAdsX
yZPQ8xtT2nF+Y4CszypY7kDC08Ux96G37GKzyL25EyS7LKq0GzrpljoDT+6481J8
gjnkVDQHjhK74+paJvMboawLVPhllS0zy/WOmYkT6qtUGYaUGQPbOezU3DxerrQM
/MBlVarXvhhUHr711ndoG4tkcnkFqF1cnyCnmDwlAl3l2MAaCLNZ4tvhpud+EsHq
60xV0f0xZLa0CJmp4GQh0aDvzpX6ZPQmlFCJKY2IjKcyD0axxV3qYIO0pkYWUoUa
lxAbKIqDmV993k/Xp+0ssAscuVKgvBKtVRzdys1/co6SNCmcutwEw3E+0/em37nU
uIFFf9SJ+Q4zwxvHU6voe+BcKSCzQWkcmqbF+Ek2UjlOpu19Og4lkRD7q/J7BYUh
ghD8G55BJsbr1xrfn0ZPZSh9VHBs++eqdPWP3LqMU++vV+6hBcJC1FYhf18J8/Ff
qgxy9l2zVDZgQdUmwS7BeFg/JzS2T5JEGYwTw0TVgsMmM9rKIK5jZJDErRdFhcD/
Z0NWKCDJubeWdZMuxGDhEECAwgz8emHbq0ylRmemhr9HcavjmBwZX7B/TRCPttcp
770DL5X5YRLOrxtitzYV0gm+rZ+ybxh9SzineWrQQFjSU4wyr2Fw9qBSqfXVsAaP
rmGDb3pyF8YbcLcLBWTd0c5LseMBl71fjlTduQRUOJealj8nunFmDqMSTt/7x9t2
nlQSR6Oa8PUTt8s6IYWi4/fnjkfl1KrYr8epfrvTJ9MFx+mxZRqn/yozf77YGbPa
3ltOJEn3hxIKvYTLW9VRyfHL5Ktu2zlAUpeeDI2LdvgXpTo44C4t/ZML0JbYb1Tq
hASwXJxAxU52m0cHzByIirQpZfsUQWfaFz0soiIHK0p2gLh+HMPSyrV65MNLpiUF
pZZPgUftQZcPn7TP+NgKHr09QpSZ0/JuJArMI5OFgWVL/t15MZihpbbEwl5II7ng
BPNANmf4e5a5abIPpOQF5nfaV9FOMSu3oDUw4KarZYXD8LC+Q6jS9jtunSzOHazZ
/t94Nls//xqG05d6XTDG5eqM/GQMiFSwPjzGgJHfqN/P7udBCkfq+xAhOGjwle0B
fhJaOOyBYBA0/zbG60e6VVNTldF+raYbtqT23Xz4IwDAgbSchvj12AeL1gHjjW8B
CeddKN/xbVHQQU7YawZI1SdcGpSVwzBcMPp/RrVySt7BEDvkeIrRKflt5+pS+Nwm
fp8cnSHUE3BnR6ddkdXMbIRbhGBg8T/ziqvV95BDlor88Rn1bkcyEasn4/b5xlZc
sXE/DuxhOTovyxP5pZ0iGLtfEdI57DtFaKxKEQdo0+10/Hvn2Q5UEGvYCjiWA0av
ct5d/tgptkIkbka2wQbY08bA67nbVkAa5QYTn9iozGUykJpkuI29mNspwxFjLMBJ
UsqzxyWAZ3Bx/a4CWwKa99IFta2mjxlorNioBtTU4QtJPyv34rMU/aKS00SZgOfD
CEmfdknFDWDdLUQf6RTIG1yme1BeFUQ21VYWXhUeMzL7jcjO/51ChPs7D8rLWBKF
GdiByanOLeoAdYtad6MP9qjuOvotHkAdZKCVPS+iSJrMi52hMXw28psWt4hiiOE0
X8mkCUYeBz8g5pLHQ/Jh9stK0hI+PygH4WTe+dh7BtxGpUd2yAN4GyBlUJez9r6L
Hs2FM9BOGtPhP/31+5ArfjAGoFlKjZCcrP+KHhmO41qSeU4djTOwFx0nJuJXK7Ua
XY/UU0OPx5qbZZ5sy/pBGBPV9I49G63xlvASgj+BWBBPAhIkU+SKWpRcWG9UEQLT
7pbTBSdiudEQxC21xLI6DrPVydQxvY0qd4IGEMk1GVS5mgap5foY3vYXndG24yT3
oNsVzuXJF0ajoF5Tic3imICXTsCLABDF79cWr6ZM9vFX0VFeE+v9kM4k3ZhztGT/
08nHAb/IrfpUXzkPttIQVPj7M4SbJgbTWw2dNkwXJ4qHAcZvuIkKYUgeCrwvGM0R
1ZSHG3HxlOaCWj8TW/3aQZMXp0DIU38EA7mj/eI3NuKZDJwOu5HEnh+rw8mzz5DN
XPWSQ+weoJNukY1ha/eE0Pxdk/SIGDwMEFAToH++zMQz4J0X3sgVu/jx6ckAbFlt
qvnvpZEEnOu9cw8ceE/DwLY8FUWqorlJVt7V7MVeJ9sbpR6JxRVlRALCAjmfbxbh
Ob13p8KwSTQvzOEjEbq2Nl7wqzq76Relg08tI02OY26y8MSgkdQ9feOK3SgBS5x3
2Jj38mp3/cbBaAU2b0CDSbm3x1x3EVFM8uxFG152AQap/wZMsFP6st6kCpQgdcEL
+sSzAOSAPwwIG034/HygYTemRVxrKh/Z2O3OyKT+kAnrMUjvk1zNy36+M1l0KuRk
S/3Sft5LyrI+IIXLIKYSk/Oj+ByTinPVZMMak0qS6ZaNrfJ2VT0YphNKFNSgm8gQ
gdu5LIxH36LmV0eKXOj3UMx6fxoB2+qezUANT3IjzqAE3Iai8ox6wOIfKO0/9I79
/2BuHszOuOnNwB50wZ1czrPRfoqmifkaL5sfpQ5IgOLr558NMxTO7cCSTApwsWAb
IcOx4IVQDRjreB+R67UNZEiRsUSqMs116IOgnW5CQSWZIfo5F6oJmQhLtcAaBkHg
FB65tnyZShEsOH+967k9mXfDszMTy9FgbH9yhTd31BiS4fbXHVhzji9+S8Lm92l6
qQG0yuCVHC+m07TcBjFCNCVMC1KPGuZsj8hl2uCQ/k/ALgPsGGX/GeohXxrMphnt
iVcBH9/QQcMLFB8uQiGTFZrXKYs1tC3BObyv+HUzaB0x1AJI1B2s2yY6xjtvjVZC
kSeNJFbCxFYJUg+3lwbSBmcsPwcktsnFs4kvT45JBnf9rd7afwGIgz43A/7JZB20
g4Pj8iSCWIlQRjJtOWtFihqPTXC9ZEUA2k7BLHxXVP/Lsrt+0jL0d/rlUo6sw/mc
fGtKKf0PQuXCOUUvdjK0fCqRdHf4sxmvvXQ7NxkUquCYIDtqqP4lvcVfdeZE1HSf
urgJdlpmr819fvuxqdeanNAVhNZ3yWEtAjHnam3+iK8JmpNfN1pY9TUiNai6i8GT
7VONkk85HOt05YbmabyAHuGXFp9IEy3wYoQoI9yXcRxMSdn5qoIZu860MlSZz++Y
7vK4YuQXYqYZ2iJP0ZWicuLA219rzJmJy0OyIzpHaY+cdgpzAHXaOsGXY6lSFScl
hv6hjZRGttCNDjqSajZUNyqDsCZmoaZBrJO+DrV/k5ulckEsPjoLC16PXDOzDkvD
dvwXM18xfawSSLBf/fw4Q9tSQcTFBZl2guQaFHE8wI1CQsaYu8Qv3h4YDkEsOtUc
HL37PLl6d6bsOG6M2YSFiqM2f2yCQNVFUGUU98ffQ2MP2ZsCdlT7r1z8veWQMH8x
eW5jIP7FRrz8tCWDdOZ+JdbhfmjwcW0aaGI6c0NcKV3jeQkKxMvZ2x5ccZ6OiGIr
+iZ3yNkvph4AD2NWOuUk6iAwIxMiD47LNg9pFo2hb9AiOz6n9Ic5IO3O2T37KBq9
WUc4ZaZEAfW5+DXaqY+ObJyjv49Zx2xKREqcA26kDbV8VXdLcGnBGVtXMhJ47VnN
wtpYMYLX1ulbuSaVypTGof98YOAsyUb8RcsEU+UThXNR0eubqASPErj1ikA4xn4Z
/GoTA2zKHRSktjB/l4npJaXQqAB4e/V7sED1EhuUiS7i9/BPnQZZY1CqmycNFP62
X63DnvvTpVtfzVy//IQCckXmEKhnACTSmsiFkN3pH+DqWynTb72hX51t7r3LYlBR
ROi30uBM/KyA7EUtksOqimZ2FVd/2/I5vRr0p5W4hv/HsVLUuKE+NP1GU2E5DaC1
Rl94oRdRvq9PRDkClV6eEbuoU40x8Wk0Ks3tlMQdgBsmsSXJvAWaLzwuOsAr9w/C
i6IGPh6RyH369NiVpi5LUkL7HYf7VsGXlcNdKpJ9mC/G/6XtOR+G84PnBO1d9LTW
5hCRVxlKWt6lwZ/sjqBNdAMq9dOdfWckUNRsgcIofWAERG/T+NSPgn7nJfB33qI4
RSPhl5ZkKU/YsKTYdJ9zt+I95Pt36MXvXhWr4cRDQxWREOkrQ8Afb9RmNwq49G7M
BLJ9w7wjmt1HQTl1sV1J7SUqG+cqELWLr8I05Roesuo3fmq5daHmQ/jjIR4Gggz2
MtVYVVPAD7fIfnQrUL4cBJPaxX024VL5h02jHLx/bwZdjcrM8owRNiAYyYsA1HL2
I1cqkZmUFNEZnzHPl+Q4sFP8Feu1fTaUPNhnweQOtK+0iYxA0AWugQLX110CcCoG
mMiUYt146QKO3HoRtfD9x16aY77nO5dfEZyUz3BD4T1gtujBNZmOKBepN/cjsWe8
Hg1JmDaLxPrNwTHH6h2frt5VIYh9N0FPOU9pSsnb1MQ0y/5uNz3lfs1kwhj3kcN9
RtEqUY9fy3R8zbNLn83QUPMnt2J2YZP0ZMxfHOW9HbPfcxRY5cQkjzN1xFpL6NHQ
8/lwV1z0XKJfG/D0wiag1LqjuHa/gbfYTaUwouU/ajEoRAcsoEqX1W9cnLlK7KjP
nmhs9uu9WR0E2AGPgen3vzFXc8Rkp7ZUHpD8VRV1MLnoNGMvs2YEDqfcERFg3q0P
83kWMlbSriRNB/SHJ83rWamHGxhekXoArZCIGow5KD4no1p0obcygsMFBYuIrK2K
udaJHXEzOhtdc0cQIc4Rd3cXJkOiVS1cCCSortkkGUuHdWINAhNfugWLTaoUdo1X
qOw+91pqYKUQF1xFpqvIYwfOabx7GYzvZ2UTnP/ge3HN9emrd42iAsl2D7fRVelk
rJob8RxGDfoWZimzc8NsH0bJGft7SnPynszFpQErWu/Ugm6d1SWtg3Q0rgKaF+2S
6iif5umSFJ9uNkKI8l2+rjKsd8BgBOS9MsBUEKek4123gSPqUeLduxj6Qd7ahMP3
fd+Gr7D+BO+rg9QfisyENoGBVAEC+xEsCm5zCuGmyMc5NFG75Ni/RCGLt81knpd/
hoJ+b36dhVbg5ZlrguxGAFzNdOKurV/D/Ku/WwpxEyJX1NfF3ncd5uVHL8ZVnQWm
zUsQeFvqvnygu0bNCZZniL0dGAbjz47FvuudSptnmDBmMQmpu75on1SQwsE4SB3E
nHvCw6YPb3sreEEYqVxcaVzV7N/48N5jTgjE09f3r5Tk+pAjCtWEC9fGTZXqOpR0
K+N5dPtt+S6p5mDWSMZxdfLIF7nYES4UN8H2LCIII9ZvitSSNgHKRyge2ltmTEa9
zZ2ScWfPkIysLO5mw4Nn549ho4vEIVtJqhhw9KSTuczefLXPkHAfaTuQx4i93jhb
WmyKypB0TJ0SAkMERhfgGPQ37KL0kg+fa8BW7Pje09AxS1h7y0RdLmr63SEYiLBU
3346BYcwRREZx+/qqCqOT0IlMvBHzo+tYteIDh66PjNHnaWzwZ2gmkkNZgn/abEV
Vh0kOqQsFFfbB5u/+LsJbDZqq+HRGr5HNgczLUWDLFo4DJibCpdg50dAeb9zoI8N
BbvM+mN2diWMC4sdbpvBeEa5HNR9gGv8MskysQdU1xBxEaXlX70Al2EMYZFd1eyw
e/3tAbYfjukW0/qhz3SztjXOvr97ENdRu/gw0MimunoQRYd5dONmwo6iigsuoMVm
EkQU0uFbIGZf+5QrW/NBCCwGnR8I1zrAvDiYVWWfWAk66Gu7tfsMXBug3pMuQWIM
uxdytfyRvEjUbabJkCf3W5zpPG0Bb4LUzx0GRzt7VRYgoa81oXwcMF2S8k6aOCHo
AtM4SFDQDlXlnAwZlCMrzt2tzjSmqXnV9bfuSEYgwoq7bBcLNZ0aMCUoBsNZmqvR
e0UT/Ir2Lpjx95nnZruZzYo9aAomC/Bo65nD03Vw1P1VwNhoqOhDBALUQcwglSeG
M+ZKjGIlHRdbSbadFJi/wsqa5V40QWlmjcfhw5qXXCzCOwDetJ1rF1k1PwwjhmDf
PB+UojsT694ng+eFZN1HYx7psiF3ItAw43jzG/JUzSWdRBGwgDj0NEd14CFJiPr/
swSPQ92Jn3GS8LnAGzvOyq050CWvRbXivLEjXaFz6naE8ovXt6O8Cykryl79GZ1a
LxJ5XyVOChhUltxfQwrL8Yqq7Rcx52Wkyp64JT//PATnQslWwD8Bh6R3anLyx1L2
8vOV1vIw+5geJ7X1exifUWi0ppEO8BVqJpT7+dhwHrWfyN6Rl9ib5jICMyS6Ea3H
4L1Nrx3tlakDgq9XGGDOEdr+N+CkZWHby9vmg5xRumBoUYaScT8OQeFlflNYQHOn
92pmlBM8xl/BX8OF0ruuG+SSZqjsDlSKmU0GSjVCt6569aaEiBA6hrf4RwiI3mdB
Ry0ahkXBQ2CoU7Yf5XSHEGRUtoXO8IzPX+pQ1RsISeBq5QRP2fZAGAfTjjSFq8rO
ZYqe3RAlomE6i+bUzfigrH4MHEQvlvOLhcN1El3EXXbqRUpP4e17Mo7NXgLlQpEo
5mzQO6RsGG1e8e25JK7LRRiloXGB1ThCm0Z7V1b8LFZ33mMU9L+l5Fh7x3Ixfu+0
xf1LyrIPHaMhkBvUOgAm5OhPde/K7NPCxxvja8HI3KQg1keyo9sbgV6A/V/z7woZ
wAD10i11R8qhhQrDom8HTtmHQarztm1fihsvZGHtqtzc5m7eTcz2A20sskx9PkRW
x3kb9tUPMJjZQusRdpHD1XLQF3ckpVuJjQRImwotxsSgChdmqNRs2lgKLJh/badp
MWe5CmcZSk6X6rigqWwy7qpB1/d7i3jYCOTFPLOWUCcwMOX5FJCO10c+S1T4v+/E
bqD2FGwvOLjJzo4aoJ63EClUEVT8poR6O2+kr74cuAzXVBjou40qgDj4eGYYoSU+
FIQYeMxM6zm0ZOVGr3CvK8Msp89Xq8SZxrI2MfLsBXw7Rs57KimTRjJ6X5R33kWa
jKO7nAwc0r9bVppBX3Q7i9ro+zifqRXnZtHsc6aGr36ZU6toMr5B8XmLiplDZI5E
r6JYrCjqY/Hdsbd1DpzJ3hdYhudEl6xjngLln+xDU3UXHz8c5MVPOgsM2NJkBhwf
SFeB4GMemd++uOtkhu0q4RpbhqDv/6lG6fxm7n71lWFGSLwALzRo5OaIHDX3UNv1
n0N2E8LFfjzYc/tbLrnp/70r2PbBdIIDOYBcJmG9zRqOHF3a0pXSdmWGPXbi6Blw
FklH25XYbpePNVGQLu40VGFYOWsqggijWxEUOaOEVweE29aXcnAxiAA3VFHXNPag
RQX6RogKoKisEDwKphSG39tVU6Xg99RwgVuJom/azSHh0n25GKil8KRWGz60lsSW
iKxSxsSBjh4ZIe0ztVFXb9rdAFXO7+eYcfh4FFuJGSARjrOEsFo211GH5SHkWQWX
HaiXDvWv6H8wGR6mGWO4nRe/xdfari/adE2DMfb3hohvGOcDTKf15Zl4Zb04qwdj
5q5Flz7dAQgMSeTLUbtrmUlj2KzhhNnpnmBrMUQ7i+LGJ59wp/eY18o18SQePMdG
jAlEY/Pk79Tld19cXRRO/cVD6gGOC3gRlUm7mC0iuyVlhEdVjc197ZRmH5Kp1k75
QjvlXi1JofZUZq3AGA5w/UrZq9a61Q+X/6XY1C5enXY0DsiSFO3fv4QWxESlEq8/
Us6iwYwALD6M7DRCvZZw5FtT2i8goJcjpLLRzUsEF9v3rq9fE97lKRaaWYnczczr
J17jHtc0ROZeSs6wIUb5E77U9LPnpIBSrNQlfZAMKC2J3jA4NbV5+OkRS57Y02JX
sFzArBINLhHiM8N4+RkAz+orxsWlGlXhNMc5Ks0gUZ7fl8b+AnvRz/1UmsAReBGU
BCSopp/QSbfZLDcoamcEEP+LxO4PL/U/JIR1Ez/nH24SIyuzN0+cDoQukFhC8aIL
r49lNxf6Bvx8e17ZOaL7iLRTIgzaKt0O7rmj+y3JnhcpoNfmTF1hoqlzuWecIl1M
WkpH8BHfiAKJYZbBn2JoLUJRHtpkSXlT2Ko/+bMUaSw6tMopMSurWSwcpxyyt0rz
n8Ok6HNBQq6KT8n3DX/XtOBTyPrZ4YYHXTS4bYXsCvJSZv8lmMQHaJ5djyaF5I4H
MnDSAMDj2nZpydyCPHMPIQV8XygQIw4jq2MS8AQu/goyE2R5UJnGbOSrI70kyq7w
C2ZWXInXQ8Xt9VR0zFOFP6QbebdUT1Y9re4MiSt8xHqtIY+XBkyBn2ytv+9hODtb
pb2p002tpsppJ7FVDAcZgPUXtUr3gxGrIz4cGfyy/jgJ/1VHCTi42leULiUwvZPA
W6+HWX2luQlcO98A8D+0dua/5cm/YvrI7U77XECZo+AzKAEuuwR5mlaX68gpgC9F
q/dD0ebhgdB0/5j12Dmqnqy8gmR5WKZIZAPUWtnRdAvBmeTcELSvhwkcLTJvahfx
JVTCx8idPk5VnqmZer5kqb4sjiOMlwQDP2Uj+BVnmxYIFenE89O5cgdlPhzrRjDI
H4vcD2x1sonRnTuFig4xdJdRnmg0c3sI+f1qY9FtSmdTUurRWT57TXaagYbeuN4u
kiMCXHb68pUbSijE5YlFGczCdkIFfwNXuHgp01bdEsMwdNKf4kq3LcF4APO6k7pH
I0ljZMcuRSPlstt2etVzumA++4z5cEZkq6RkcjF2sVNVGh2WMtzYEwBlkEqYutY3
g6dAwaltgg3trGqAuZUudppiI2bEDUSxn/irH3OYTloHxPm0mNDehcVdQspa41Ho
Tjl+TGAY9Csb0yV8lgqkxQhYG0ngEefGfWAIZ6i7/SCrYE8/XKHFwttameftmU12
x50BF9sxPFOtIzT59HBrambQSrNp1g3fVP7ndjunyX4X/hVELED6ruEUjQuF9X7H
I5UuJTWoCPbV1juE9QtA099bNogmQLRxM3Gk5rex48ELeQOcUpkjRHwTEmp7bl5e
g/FFK1LrSFcP3P+M+SW51t7g6DkEYQ+4yeXz0Oo3V1C3RFTsB248fX6cJVERPhWP
wprCYhGoncn2UFywMWZpC0EygGZG69rPaq4CgCvhKZmZHGjQVxbVnWLEr13HPstn
WBUGuK8v+aXWq5VwG48vjsc6LCKj5cAD3KZ7MeedmepBFFZpO9beUYhk0XyxQAVU
/EUFEBA7xk1MWZGgHHPwXRs7EcS9MufE5A6NMkx4ih/HYZdGHrMEHF5H2QZCe9kQ
tnlIg4iZtppUryx4vdAHBl/upy/9TsM6HxZYVv+thIdOeB/3n6lORkSL2AxT6mhr
N8SlcZU5ktjMcbGoxN+ZTtE2qsekVkohLqIOjNr9LXrA0brhJJm0qTSXQqEpuN/x
dmuE8Rg0lMNRUQxfmADpSMIKp6xq3dNHuFZvEvqVYGjKSQfInJsbC8qTTVSXhOUb
GxNWJhRecAWcKbnEIM1jLOnwuwrf2HRCiknV1R7RkIFmYUCrz31j0Y9YDa+53jMo
YGO9AcMuw6iEb527peGzoN9d1MjHykjIQXDdPG7KGQfXhkYeuAogXlrfaXWsT6uj
QV8oZ6PFoUvRxe9DKyf1axz4ThEaoc3BMQfqLurQ6JBQmpkzobsFwVeXFen7NFFW
ZgxGhiGoXjfXkazc151QewNjkKoHhKpoEJxQM/eEaNSVRTM+OKpT6YPQqfXSgPFH
VonG9agABaL00Zb3i82J2/UDT9wNt6C3IAe118bvfmzJKoIWt3I4zlKgnJ1JZRGp
DTZkXcWspb8PUC6hnsdbFg6IxZl9SCKuJkC/ypAGicVQcgxv1OIeMlYsPBYq9Tvr
/c/kYAsyQ9ecNCXbyvIB8e7KUMGu/xD2zeNro+80ZoT+9BSpnjAin+ENLt+t6yni
0xWctaBaNq2xZClyFyXj9NPWZzYqc8hFVrxLf9pmWr1k5JXtBEQ3Z83tCq0FkOlk
P7uzXPwEXUzZFLCWnk2rtcIIf0C9rwXERYv/O8kzMOVMTBMCXhaaOQg9ae/Bz0Cy
ClODsBSYSaCyHjoMj+exqpleirOiQnvCy1CjfCMxsu+rpCcs9sFwI19oehEfFmV1
vqMeyeqSGVwcEG+UbtvlbyPpa0q3wkRQACP02g30/zZcmGppZ0Zxt9houj31og1W
xZjCjuPHQGv2OJ/kQTl9ad785FUqt3QrQNsPPiwoVbJD4RVyO8MZKrWm5ELbAS3u
jNdTApHCDxcdCh8DtU9VTEg+jQAdPezQSH+m4R1upH3irODsKQ/IPgq37ZjDTgwP
txuRU55VozFl44HovElXsCautIcF95NqtfMcfocBs+yx72NZ8ksEMLWRNgi9H+dU
EHacJgfF1oeY0rY4QV7sM2moC1RgCjhH+7rQUfyLd25PSXwu/QPbJ6d13u2hM/Xr
xiPO5Uy19LB2eqnUQCDAGDuedrDLf8JoabPcwMakm6YucxLw0juyGrrh0ENwkXIv
AZ5C3+8/75Be9tXLMwaPUB8is0tq74GDWP9BDAQ3mI2eueoD2qKC0Mw38dpfMaLx
l95KNNBXnl9x6yfA1rbLujGlWZSJKVzHxsPPxvpMbQ+wHWLgcGiqHtj7VPKbIMD7
ofo9cEM4IAtQa/0qCpECPqM7mkGf/TUboALLYA2bbqfZWrKeqoqgRDeaF8TvW7l3
ECYzOQA/WfHdqQPDCGnTLV5lhpwfekji103QsfSEb2NdMp8MdfT8K49zufpsKlfJ
yBt85k//SsjsgnfQyNRh7D/PWYpQ4nY/pl42v+w4Z8wJgTwjkL2m52pouIi807xs
/USqnVSqT41KD7DyUBK+YrO8hzr0RNfi2Wog+tK0cO6EiJVRjBcSHMTuJz2RZuZz
diDlWkMIbeV5UE1f5Gj6V7O7z2Jt839AzQPhqQnNbIf4Lq7E0gkufzefMiTMo1Rs
Y7H6vizIItjmms/3Qga1uoa3DxCHdMnegF/UaH1uKrE5a734Y5H7GPldyGm8hh6J
ZVyfQHmhu2jeDpmN4Qkh0w6pPGm/4Yz7kfNsmptd5sCy5RupHKw7aehEegAEGCAW
HslbxuyBab4tpqjN+i1Aat+rmMTo5vuPBxDbxo82oedxTtHEKzw2HtB38KJQLYD1
MYh8a5AZlqg2bO4UZ4NmXyYZU9KnLJTSkYwTo1ltZ3VRdl9E2Wat+J1wsbno6C4Q
9opCAmgPV/qDCOIATwlOfrj/atYIhJuYPxkepHE+M19U3H0B7bOf6Ge5fsKFC1dS
H0tc5NTuAXvcD8GKaO8JQoucL8/XmjXYf4QSNNZg15mhPd0wz1PDAoftvDAylK9q
l159/g6xVJg6afKdK1lv0SalXcczXWILtpljUIaThD/rvMe2ancfyPvGfzmFZRtH
xYc8N4Qg3KdkZlybaYoR9ukxMYbH+vwSQK9vKxRGk1405gqu0SSQ4vxqQjGkKtw3
AzG6f6ATwj8e7enX0iz91tshemxDsGqsEbqStWxk0QSMg5NiUngQbd01qyPYCWs/
QkeKS2MKtkO4RVVSSorvo/fEEOiaKapJxWcd8f5qWWQRYo29fkkwaJM205/YQHU3
dU+WW16stgkWuE5QDpbgRhUHmRbtTTkyygQOKRntmvZqMVhActVZ1P9Fw76GqIth
LY0oVCTtPaMcSWlppfV4AKXVN2k/BXol+vyyDC/zObfCqWMY1XPJdcehJBIka9j6
v4D5+HqBrdS2T/l5KLT/FxN+yCJB119LFFazt+xRrhhsAZ9Fx4VWD72p1BLSNNRP
379d8B+4V00kELZN/RWbHKo1GheR9lfkXwIGHhSIrlgMWOrNa1n1wVBxkjcA2Oqv
Gpo8SByQN2HyuEa8n8dxCDR9tauGCAb32bYccZNLoRhj7LLDWuoLIp7L40aOzIde
dbZbRed0R5gTzhtJo2ANUop1Cs3aX3jHnGdoG3R3HDuWo8eZ1hevpyhDF7ywKbil
TH/vqskshas5cIyRjqmCuBTO1GMkhvjwwTajME1wuPouqrh2aqJ5aANj7UYWO1f2
4b5AJ/AAJX4IhCceiktsMWBLWLA9s+G5mYGxY7ezOrAKe4QVwXvva4Wqr7MiM36o
bhhMqrsEdS1TA5UfxrsxW0VU5fATnI3IlYEPUuf2qD33/ep2vBeX6etTRvuexTQo
03yfz/DBDnYZOPJndHILBdeasjFUxD82l12FHBvtYT638NTSJmsxngivmBvl4ASE
zKOMmuinvDblyfXxxKyrWz3CyvbW9g8qB+ulog/D36bWZ/utmw+0RIRa7pdOOlt5
DXWUXCSwnjjVuYP3zyX1+WNfAYDs6Q1N2XdhpTVlklq0uxNh5kAaxv0RO/bDFKP6
Ss34md9UGZRyW4/+WXFPCpU6bP9eWB98WD9s0tbggsR/ouYlXU+IE2Z3P6Vf0Nl3
8ccMDaHT4kxR1vGNrEWWhB7MVbY8i1BqkH3Ms1fB86tqh5I8aRZ/sdDR32BWe5JH
Azat63iYlZk6ZmLfk3z6YNr3NERuAx3u6xvcxAdkNJynXr9lNG7JdzoP8eOOUX2N
me2ijpiCSt4mqTB+EoE5X+dK/X/fG48nmZ3TxlggW72IngrL0yUUrDzYSjB/adyZ
G6tH5T9WMFdcrzz9LDEFFHnstlGOMp9pEdKHHcvPwgeTH497rm/mmcxvX1Iw3Scg
dVGHRng+9ucg2C1GAvKIikoJE5uohvtTqx7l1LZki2KkwdhD3es7DXR7R9VkAGVQ
Dfi1tH+jx1p4Bk92MiaXz6H2nV6Q5l1splb4JrZCk/SlV6UvzeLIyxTz1HbI7O7+
4STpxngATmr+KQ9QMswsCtCeJNNR7ijO+AeXPEz6lxcE/2NAt7k07PWJU8L2kQ0S
8SZy7ipDfpDxS6WjUZHWtoL/YlVYoYhul3HjVeP0pyLc1bMM6liVpIEuOigIu6kM
kRzQ/Czd5lfzznbyXKPnEG98A9VkmKwvtwlF09TT4T+TYMWrTC1QH+Y1iP2q3uKa
mGf3i+9vmfnqtQaQUT+9VYjhbjYuU+AAnybLanrw436w5jndWOhgoFu07XzNQvBe
xYwiNtHHnDLSKIp6ukwi66fyqPm+fIxdHRjmr6EUtDTOGW2okIlIDn3+62DPAuUk
PBB5XdOB3ITI9AFwOjp2HufgU6P/NwbPbMLqAw7huTyVlw03MOk1eJ6HuMfnuPaW
aZ5ek2QN16Kq4T9InpjxeZ6jAqesQi+j2IyhZp/swsF6IMsxaedXhXIEDDmF19am
SDLOZBfqMH947cWpHW21gBPlkkVPnusrh+5HOnSKnR3BF4IkLlgcD+Az8VH0Nak/
m7gjNWk+gEuTkiV5SP533So5I/1l8yt5NIRB/cJpyoFJnmjPtmsF0d5q5bka0QzU
jNjIsvNq/M7KM1fhB0tmMQQEdfZAiL21uUq0aGjfoImsUcvk+0tZDLb8fIoWFGGo
sJdiUkO88C/RX1ZPjpBgc2apBsxfqM5Ypa0a2es8yiM9geoBjrSnXKrDYqOmofbN
gqvGVBPLLkIaUlL//HPdZwYZoSdiMgDWJv0u+QUrmY78EEwIfplKSbUEp3j35k6Y
ml0fZdl98kudsXuIm2ZRoFrioGg0Zg46yDfhwPdVG9tH8eMdsCAcBhqC1H96HKNY
SK0qfbePZ2+AC2YJVESGAks2Y2apxwPb9Qa7fhtCD1LWcJ38xTed5+WbnkK7k6m6
GHXt4XCHa/4x4FNdIOTXoQXC3W6xaur6uHYSVDLVcXKm2yXP0gtefhNsFOeWEIEU
qGMF7TJkFJMe6f8cgkIL3IPvhG8UYTXBycfrKQfXG63915hw2uRVRXFyNHq5Af1c
Cy562PtGKI5dofb2P2iGPQTfn+WlI8cP91LkyNuiz/zXDthSZGL2TbymH4gT8ESb
X0MdYTHl/1e3UzXhp1x/TphDlAWsk40Fk5kdyz3LEtnpuwj8SRVS1hsQzgp9DSMW
yjHnZI+s50BofmGQEPefN3Cw7nhELB80fkXoEE9UHOC6AuB7+qAs4UyvRAgYkrc8
m842Aqw2RU1ROt93hFTxc7lixTCMvSFyWQeopIHpKEGJ03pc86lR189oKYYeM+wa
E+NA64p1sqUXrft1yMHPKjfFQjFJiJ8p627CJGWxkLgmQMmnaP76jEYYlZppapPM
2UhLI6oeN5Zekv+e9yu/dwKdQUCnuoRmTt1VKSiT3uT7nIvG3U6o3OSYxT6/JFCJ
Q3t8w+olo7v2n/kV38QvkBjFgjn2GB+BbGr0h/KEYQnN26wwxX7hKnqQx425pmUf
V3dklGstMiow+nOIbUD2fRVjpqpVdGUwmclO3lKCmyZA0ar+E9TcHNkT2Wayh7cP
pfuMa5JzaILORVyp5hWGmxlEe/8RI5Ce0JYx25BH+y34mLxZtQxgwLOiWuZa9itM
rDNAU5XAQ+q2YGufTCCzXo9VepcTLkE0oUjU2LzsJaSWN0hKaxFnHqkCV3C/+KOE
c9hmQGFHwkOPr/7049U/jV1IR91Mx25aAgOYERrSgoxFfl/7l8D0BaMkzGu0MJUx
nPCELHdIVDGyiOVYHUj643pPoB0BjyFb05rxaFt+gbKrAysi6OZWBKbQzqSltLq8
HlE3shDG79nIETL5PMA5IilwLw/dDvtYXr8tfVPHL5SLBQ1XSGba8KsaehNTTyrB
geGEQoB12YlVoiTECtOZ9wJvamnd087NPElmI5pBhjdxxhUT1rExmSLodWPq2rrU
ssRMDI5mzXMPiKgq8u5C+SwwpNzPLNg8bF4hGGsJOeg3ukFZIW2AZwP0iSU4+R2X
f3Xv+RqIHanvlpPEkeAcZQuOsD6lQxUQUJhiau4q/f4yW2aBXJKqTUgUEliCFWuG
FfJ/WKI9Dk25Ygv+0E3eA8klbuXeh8QTvIOaQQXGp4fPOXKgTluiwRPBkaTSDoVX
1D/tjbE1USHy2/lDbS8E7KgGkBCBZ4rGdWuESIraxkEjzDiUHZRJzBURnSaEKtc3
vK/aC7LKaxp3imcSxMlcEnO0V1mn3oj4piWgUEtSb8khjCfi11PjW2azIchY105r
6ZdwcRbNNC7QBgWTJA7Cx2YNuc2qPfQPi7qfMI9L9QeQ+LuK7n4SLzEcj9gBOAGa
hHXOqNbiyxSHdkrWUXgrqonDw2knyU0eyyM8JBtBS6xJFR7M7WdCMlqC6BiXIpRG
btvyUac3WsDP3/7JpgpDsesswXPCAwuzo7VSmpi5vrqdAI/CZWey4wOteEL7CFw4
0HFDkbUHKAPJoC+Ud/YM8hy3yUgE2CPCCEDS7CiMhPVeEpiQ/K7kVQ2US5WrSTjC
MPKtEqvMkj02Re8jzuhHQR+ohjO7p0g+NDClutOaUOifOO017Ir80ZpLNHJ3lgf5
+cTVoY3bBMD2smK21JeFaJa2rLrVl4bbk9owTXHj25jne0OJOonv8yxulQORo2Em
vfyGRKWBbZCK2zkwIaoI3vGWvkuN9UeFN+kD/gWD6gB/XxuGOCBbcWHQLvw2j/DL
YYQyITqvUPrrUk9W20YhqtYk2GsziFdSqOMPGPv5RWEWlyyS7MsnnprUkScpSFhC
ok81Z58ELPTRyi85AGBrM6yVvKXRQ45jIVPiCn76Rv4N6qk2u49YZGExPHmpBfVh
X3/HSR4GUoVTIRARk0Eptvb2jdQ37XK2y0zKRKmyTz3tbznlhnJM4g0+a98ci9oO
bMxQrPz4m5LQQNjEnFGLdby/EF4NqXmKlLYwNCg3hxwfswmg19e+w7bSZWBfPnMD
p74p38pVGVSj0rg7jTlVUglS/OlxOCYepYnyqKHBFs/YPbmTtG7wC71b8IO+9gE5
25I0yXnH5Q0RQOblKXihTe/H439dJDafMcKDnf6S9hmRRnznhr7f3ZbaY3GFNjDR
5uWGeSPJUxLtHh1ATe82hMU4/1EToIlyqWfSo91bhdcMKZaIiEo84i+W9Qyu5dsZ
YcGh+BHChXAVImj02vZ+/te4L++yKDN3qwH+4GhHNbDTqyTIOBiXt4yJBZ+6O29z
f7dUvfKl+MABrlmZq9iGdsUDQB6cD885B63mRZzJ0/vg8xV0xOZbyu4uEuDM3wCT
G/Ts/kXf584MPGpqMIRpLiNoMeIaQENr5MVcrq0B0LntfKUNVEOvNpztZNAGZkJ0
Xdvkce9Q8ZNe1Bvm/MyBQMzf1hyTTdYj7UCO7CaeJ+8opMEddV5jskEgDv5UvwLu
Z7J2dmbGUuDNzrm9w4Mho1IUFSDQ1Mff4CHN0GoY/Q3b7VN62UidhjLBOOInTYfC
3sW6Qpyh4d79iWut7rT1iLq+xvFxkhYSl/zH59l4ou1Oeporo6moEd1TLZ8yQyFI
5AyjrHeYxhMdNPKXyxOwWzu9beUVfmHhXqYFBvlLOnsG8kkIRim486xDlE4x4X1T
6Pw6qWcLGhaORe+v0leDMcNaVlk/xKvk2agrMrgGTy+aur5PTVAgY+uAsu4P5YBc
bDXoTtjagbXeh4IPShIWQfE5fYI0q3VlVOIOSL2+HcWV4KOFNHaUT1w+3lYjDRHN
mNAIu1Iy4dRc7DfJ6UdcTnfdstiZaIADuxuMRYCol2GBGHewmL0QM3s2XN9SOXqP
mup0JYafVhs3uJ1mlAuaNGs+6WFr/hD6+IKcaCJJ+Cwhctg277XBPDoi/vWd08WY
lZlRJDrZpfrzZlKYmQuLovRt1lTjEJy419JEBSai+aGjE5cpIFoKIW0gL1Pin9Ws
AEny4WlGrJIeg8mXhQE5kF0GpM0Q0NM5nE9Y1fezGl0gyD5EBzY5HYIIvn9wp9GA
zL3J99X38/yk3/4EzU5D28EZPIWJu8P6SCBA5t+2YUqOXtevhIG5a2qVM6RtqsTX
vad0aMH1gBuGMJ17qFSHsn8iq3wWLQi+mm14VqKcxqpEP27tqerFy5EjbtVlq2LQ
4o+AvII2SKwbPIS7nqY20hcZYw9Epc10Fgy3lBbgOXrjvVyWps/jEuasOFGTsJCt
Dq7vgf7RT42vdh5b9llSp4mSe7te1nOVDnTlinjTmkFih7RKmGAm+BKlqiLZpQiS
MqqEmn8lAiTnkU56LRMc4249hafYtnlo4FFyFNJRtLS5zW7DjiloNnJKLS3sJchk
O9iGYmoEBSSMY+O6ZXukQMK0/PFCQzdcaoo86Pl3nX/8lNwtLZ6wXNFYHnTxI8le
ZU7vkr/8JwbL1er1keE/5ng7fmPsGOwMrelMUZKFkYM8tuuFun7VjbyChP15i5c7
DPR/a4WSfW8Ze65NFUQHREF1GpwvlgZRj9jdy7in5IVGHmSEiyLgfhmEgctpqocl
Ku2cqS5aRKW5rZfMxF9MegLpiMP3j++bu2cBuskzAMA7o4NH8eXUuzbvY3acNI8X
yQEdx0WFfQSFti2F3+bkqNSN/LH8PJbFR44q4jK2+ufeHza60iri+qerJatXGaCV
I91En4FH4x90bSGvur9FOy/HwdPg1zmLGsOpEaObiP2dUrMhHqS3b0NFgme/WiFi
5dl5jaxBjzR+dzpUDkx1oRBHrpLu3rxanxcmf4MAl9AjEmari+47ZLMJ+NV8Q11S
qVMPjc59hvvR2iaxxDa2LPgf8ItCAoRykL2fQe7rbAhdPKG0o9V8pCHghkpSVpB6
XjUPQfGVwm6MplhH+A+oRHRB82lWdfV/d+zilhchP7rpNC3nvywOlZHD9dlbrWhG
vYb33+qfBy/l0NR9oLzY0/5qJC7fS4FwgjX4WqJgdVl6qEu/6d0pbRcl+Yjt6xia
gZGwqlpErHjjeNZnASG1yvapTUUdZuB4tDa0/6OcrXjHATNZ/wks0W10gMQiQOHN
F31Jfk8qlQXcVdt1hyoyhi/SKSlAEh4j2bvRU7AND5DqY2mkiBvdN90B2hwiTNUs
3Ib6Xb3wqt+jBMlRNdlhAxFVjfWaWr2gCLQkrImLpgWBpsIxB3705sYICWNkIoRY
Rp2n3ktBzm7qlzzZXM+TTei9a7Vd8O/9B8Y138L1mD/8tco0tZp2c56wU+iCqoCq
0G+BSl4qyyi6tA5MLX05Cp1eKsa0qADnSMThrkeTraRDj+31U+jeGP3f4Fms84BD
zNJC6sTI+6xgYU6i8MqAlHIut1kj0R7bY5Pvm+CkqD07M7sITNTrKQs+lPhnFz5j
ahuP9T/NSus4QiEWcIk9P9NhFY3KpXIVNVwedTkvetVG0IrSInnj2OtWC2LXVdka
jGIvMCQGJ5egp4ABF6WYxBszWNpP38Q7gLsV/vVI1fERtbFOPElMeNhfJYIk68Ud
8HaBiIuAgpKQcMPQdMLiqZLLlQEtaW3txsAI+swypLgmf1MxbhJREUXL9PpcuAP5
kii+tkt0EiPjqzHXzYkTQ6gE6OuHM8NhYr6nVMw91D90iL7+3rba/zDlktQR55Pp
fEnF6gGKOFQqK4z3x6sWUEfvaIV/6umgDaz0u/66gZoVAm81EUCUUrgfT8Tsmba7
m072g2IbDh3qlGcBCvo3Opri7P+UAERJ/jz21+RXuHt7fBbpSFHCCDMZiIFBTLJK
ZtBM1oY2m6BiBseobBEYkHsQnHwzTUp96RBGVB5y7yYEJEzmqcWTPmzjq/N8Tnxp
inzMfvN8DFq1227dgyMpUXJa9Qo4G+usUTG7he7fCx73BKbtgkYVoRY2WBnzEoiM
zMmeZRtCCNOeW1I1TS56J9UW5ha/a8ftpc7EDsiiQlyqGTQWdo7U6NJgR0Xr/rgu
juxruRApsVsCfdMQogYIhe3dmvRngzq7SS9szqkGkUrS993YQuxlYB0rpgAlobHC
uEKW/gII3NonkZQdmod8ZtGa4TkjSo2pzpcEv8WD8hP/ozo4Qz4hcaAtS1Ie8Wlj
SniFyl3b5eMzhMY7HqpgiQC3y/PnTaHEG4zt0Vn+i/edsd5LfJzGHz3reZ2pnCHc
XNM7+nHlqaX9a9DlS5JsJQDGRBkfw08NtO9dc6xsbJ521GUFoSbzwpqyeiTB/OG4
Hvo8QTnTPxkRfFP/C48ZNyUqZssPnqt+pBX7hqiFHH5cVBRQdbSspIrF1tS15xdK
ACBnnbyiZyz27UgqU+Et5Pp2pcWaNnD1EdRAj+zj2Bt7Scbp21K9T83TYSdrDrBf
tP+Bw2Y85i8YEyDtUEY4sa1NuW72sZe02ViTpVPRLTIoUfUCHEK+uTqps3aOYXej
tZGIncox9LJn5uUA1eL1W3fFByJix7ArvApPjnAsGNqWekfCtAIe8o2aVoL6P9AD
+dD9Zem2Ks5gPUlx+C7iYHSQiebu8EW45yblN+sfRejMAG5lqRkZKWWmwH5wUUse
WZCZrWPomlH+cLye9gjubN/m0FsdAOa4oMA0cwxYkpT/E6xounHDr4GvBEpNtDwA
UcBMyQjDPEXgWQiFTfXDV5pwmQsIYZl9kjboNPmHloHFEatkQyJ2JLNdKRCzs1cs
7MkI5LeiPTM4MHgQoMzrTuntLuBKQndHszZj4Ue7nsAo5Xmpmae1qyy2xTBtzoA2
1VUKlpbB+4l61nuZxnGT6Tl19aCMeWGjAZZHbZ5UFClQ14K9q1IW+uziJmOc3o0l
Si16+5/gxvzv0lPpOufFkQ5M+stzTvbYzc0QSbggdg0+ZpneXwEDGym5gnsPfjEQ
nRw9km5WdNfIwyqdfZ5BbLfaruwVzMPXApZovZes4PZPU2ZlXZiu0Q+Ls18qcTf5
zN+EhZ7iYHxwbKKCxiaOg2Xvd2Nrn7t5cSXr9B+AbFjL82QlklDHRIH6MksiklpW
pPBvpFK/y5DxvzVjIu9Q6bA+ieRcqhrBHQUS4txtRAG1ws5gzVsxSmqp0GhfHOv3
a4CEO4Yd/99q9yax87lDb4XoJ7F79q9BIs3hG4ty8pyawnto5WltSBR9fQPQkgnv
YmXGlSV9/waE+S7OCLlzgjY6uAwgsCLmpFvUQ6utXj6RQh0qVj8jjG9X0XJGimip
H9pPVfgFOUiLSq5A9QuJtjMiuHO9Lc/riqrU+m/Qm/BaEHaZPxabyJU4whvhynwV
OoccaOwdfcm6AgVWMbVhLpToJnddA6izNF0cvZWWaA7QE1vr/T0KhgytRG/fVfRL
pEXeim91f+CMnA0vsrrdtlPfT2RUqDkFS4d8CPix3YC9yzFMhpd8y0iFmMHY5TsJ
FRpBdqjPI+cNZ6xjWpb4lqkr3DCMQK2Ht4nx0PNhGSn8JV0bEDWQ3teHM2baBMlX
1vYLMhVJRKeu8rcbpI1rZYWqUvv86+mjhy786Ni7f4bly4SmykGpfr/gtQvv4CB/
hRaHinM2z7Qk1OIgPFeOzinpCqx2nDcdjlu5Ouo2ttaZNoMZn+MxxelB4sCG6kW6
eHC0LLLbmdaNhzdljSQUjpUrYxtDqul/IB2++QEZuh1pe6AxEG4rUdIUx5zL3DdM
Kp3CaGYxanUcFsEICxlB9uIcYiETBC4uEqeXqerE6UFj8uihpg49hVrXFMtNplMS
s0chh7DdFA7JdB+N08E9PPH9bWnV2Qa3cAWTWdLYS7c1d6+W9VbNKRlHxT4Exehe
VefM0TVgAsLbLoleX2uVpqm83AvE/mJ5tMY2Ih5ai/PzaAhnGioZrK30ezme3SGb
kyjxomQL4nJXGGWcOuK/0A1FmkYewKxVmsFQbk+oZYoT1Zw1DsHfH1LXMBehm+MJ
oHgUKdusFjflk1tZQkR6OOfDr2MsRT5JY9/wTSEMLZd7IHPRn+0z0Bn68YyM2jBL
rJx0pkJQH4di11RoeSmhwYoz4yeTgRO8gU5cS494TIdxRm+l1mcAxk+Qsk2JsK6u
P4LNGWqW8WoXutn7yo9RPSPGZcCO2gGAUHjJiVxFnakfT560uphmoEuOYpYDl7lz
KjCcu+F1tfkRtJz/BqYUEJzLY1T1yslrzKyw1tR+DW5vzydwGLuZB0fz3a6UlSV6
bvfWmvErW40tQkehoRy1EFWscXSgTkB4wYnsyKK7MYeASJX0GHdZT+vXQshk3zCT
pgB4EuzYgC5RBzF10sAw/kaQFTTLnTFj7YztukkyQt9duzSjH3B/YV0qzYxeYpvN
bdbjBckmOSz42DplggjCzr5YZSb5gsd4p6+KbPc83f6PclA+xNDoOihn28Orh2nY
tUg+MCJPEMPGBQIDtwCKxq6M/Npm4FbaOw2kYzEZiMNlzceHJ8umQ/nE058V43y6
uHSBkMsvAokszQqOVYUGs2lsA7Ej+zhdSTRV0CB3NB6r7uYvai9zT2PsZdLBr1L2
qHUfMOoS07zMOriFeXwD/f43Kykr/t31qEnv5iraKoBwFrs20TrmNTJGXI18wrlQ
Nq8kE1f9kNf9Fn/HHwJzlfbrgLyCAm+PHGLs2Q4J1Y8jk0N5y0uBlPzJReaTIPk0
BDBKEk/ZIkSoWTtfd00rXAT+LtLdt0AdU6UIqfCqbJdgIDQ/VNf+eNHQMN/UoU1s
6k+LMmPx8r1BC2IZJiE2jEemWlz2g3IOQTC+UTS/qd5v/yjP7xZP2tU86ShBamI1
jmG55aeubf1Bn38gpMeEqQQkaLFRrtDI7qrNcbv5HA/FBbwVU0FlRKs1bVosFLPj
Fz6ygkPOPTVqHDmxJ6MmjAXzhJLups+byoi3X1rFWt7Ir41P/V4ChFV7S37B3+GG
hNP5Lh9qJlv8VhljlKZQx8LL7bX+zHP5zjW9XEVqOIh9CdryLqNkesB8Oo8YtCGS
kQ8Kn40ATopQJs+YQSuJ+meRrBkDl0OwzBqakLRa47bOi6OKOI5G2QgEW0lJUGsi
+ZY+3orP1ZZ8Z90r4F7NfBs8gOhLRaEfKJ6sSt6Gq2DAhoITtwuy1P0bR6mOPQn/
T1gsghXh4/mpugUkB+Cqfv/isVQoF8/5xACvaBrXI7yWrbJxa0yK0YLN0n1yjaPb
ooX/3XAz39zg2we8CsbMw4k4z3Y74i2B9BW2PNxCi2rxiaMrrDU0HDbJj/JHPgyS
ZNAqDRLsUPrG6lilfNRRdwfJXd4Rh6eDAZzgjO0b9Fd30od/Xx0U3IO0WYRZwosT
JdFfRxDry4CatMhMoog0dQpav6K1+Pxey0w68yhxXSSrJW0OufZ+w7JX2f0M+ZWy
58n0R9z39GULOWOOKbptJ+1uhiSWlBTOTZ0CU4Q9a/x/Sottb0sgkf+IQGsloOhl
Ww8WvZPlsuO8kir0mRapKen7WKLRwv+bZPwjH38+1gP6m2RQ97SAbJ0f5nVZ5jNF
UxaDCOCjCAidNU6syfnDtIf3p0FiY2RXz6FlbIwUsqVh1IS1af5kCcEgg1Wt3Baw
nmC1y0uoNQcr4nTv7/MarqX3v5gINtcM3PgJGsAesbfSm37gAEw0jb8SYOwQ6k6A
YWVcTUyygNi2m0BdP7bLB7mmB3nJacqUAkMcOj9xcgRLnHJDLnImkX+lsYfejPxc
qSQxgKU3nA3ozIKuLTh89joJQN9ofUUkzBbYCWjUR3mvJ5IhLkWrUjAije8Pkfnk
BN+gtkw1JtzQHVdjek4wUZZzHP3RZJLd1VCgrxXHSZPZzGTEaDQQnd11qQaJYcgd
L4peorUIlHkd/eV8JMgLPwJ/IiIr6726nx+i6nEd5c1UGqDZt+tFo7SBrJRfWrvD
ftlCv0EFweZf6iYHdzgiGxPB2BHrbSvJregnM4qdUalYeJH0q2ZPuC0j+QyuRiU7
kzBe1qnbk3bWHkPyOPKsw2R+dH2iEh9aK/KCJmMYUlE1GzMEgSmExlFYjTANsxIM
un6t2qj41/OMMAiMgowZ7Nv/IYFCwYz4GWDNjQd+UPwZ8AUfIzLoEB9/utlYngQD
/6Bb8WJd5tDhGaYC1PEhakrO9piKmqLHFU4ceAOTSsbEWqTn0NYVjETt1DlY72+m
HisGOD5NPxmCMz/W34DKUD9k5g1r0uux+OHbEBsQSrZbzBayp4aq3mEE+Ow1087A
XdVaW8Ify9zh7lCeDgQFqwM0++He9Yq6auo5pC7O6p93DkmaajZdZ1Cpoou4R1cT
48lLAUMneiY5Oig2BSVWC0dd166gjwJkZV1M+fX3CmBamgtFWWtMK1GhdJM869R8
wJg/5eVR05TZ8jhUVPfo3cBvAIQljQXOQOlDCvCBPdwzDoulZlLcamHYwRGkvQ7R
+HGv7Mnzy54jsaOthboOxpnkZHSVOGJNo0NrF/ZMXrd4U+M5tQEF7eepDGZdvS5C
SupUNf3LlCnfA8kYXGUqdZ+IuPyUIlO6oeVsdYz9bRXV8YFdBdaowPYRU735f2fM
8Xa0KF2XyFI3DKRD06guFM8aLkI0NkEgAH1aXCWNh+z9yPCOy+HlcLbTVqZYvLZt
wKM1DdWhZpz66dt0dtk4dO1F5xDc197oORXzfTxN/fPOrGK9r+4IDHSwZLVQKJSG
Jzo7UGSwL88lXrlCto52pOjPO5enWPq0oChLbah5wZAbCNCvLI0FeyPGTXBnADu6
735g2Lm+KWPzMPBlKCQbYv1B7HcB029pqZrhGQATtbaMcuWXyM80oBKPelMf58iv
h56KT98uQ8I0Qyh+3s9n8U/pW44/FGW/kfwja7e1AOBH6YCHOilQJf12HJ3OHKmn
KdbcRKWqNpSKJmBeqsx8du53Mi+nFGNwYy2CMG/NoOPUjyhdfN/dnT6oQw89PE0h
SThKCihalK1Noe/I14iurN+0x/VMMVvKSUPFpsHmmy8VKstS2siOzkaZFymv2pJ1
N00xcL3runJYqv1r3l/hu5cNSS6d5Nc6pD0B6d7D+MgK0inOIWKJ0PlCnmqgiT6n
xiOXjSxHY/ZGnbwjOtm0IpxYjc9BWjyFZIarj2+mke05jmTLDydmdYTeny1PKXXm
Kh5nVBsmK/Nu979hXu4fNqkFX43AulZnaOclO8S2cR5V49RKpjZXklBoZP6UAmlf
/wrecT00KJ7gNsOiZqOeIbeVhZOrJ6oIV9YpXVi5kbcv2nmO60rTdgEPEk87t/xD
RejEzFTLanc87z3CnGzJlE/WLmwBbh5a7c9VPQhjP2JG/KbvVRnHJ+DlJiX26/VV
9YjAAowQdyd2nWkpnP6Wb7IiyscQzNUPAnmOQ2naSbGIjTmXi6tkw+dgqlpueeRD
Qsky90Jkcz/vygcIvHR1w40mGAsBkXGoHhfNaNI5onviS2QeuGPJOSZD4bxKaN/R
YrEtLolGMIfIYzgAq1giVt22rhmL3OM5o0DLv41Rxq7RPRVF66eCoUbDHJzOfXKF
2iggea9+qt6Cwmvzngx9MjVYiQ4UzYitgJTgInzraboR+K0KtfP25N/ZynIebMto
Xw4UfZthYDzNPEliW9UkS+YspWvcy7SNCmuZyYleLPBuKOj+9eGE2BsFCP2A2ZTk
Fe4xRy7RuyRDJljMesMkzPPbnVX79JdtF7tDZ8yn3omCc33KCcFdAC+2IzT/JZFm
Hho6drLd1tSUg5BVbMdNDYwU1YEqorVaUM+kWYNNdfjmBpouE3PDCbRUWKx/+huD
mlsiTMRI4+MKiO1B2b6KpzmXefpu/iGTZqVV9NwxAaSO6dCx90UNoi2mRYCXB1Km
FYlUqyvT08Cqg7tOfmYMsBQCmNGf2lq18OwMqhBG1JldnDmRQIt3i+fWcT4FheHN
jKA5k1MEc9wgoTKkBxLE8iuTDxZB2VGu5f+wLNXyRcn2IDZvW3U/QTALPTaeoi95
SV8TPvV1CGpKjy6RxEqNoT0+NwKQwvA7d49z01qXsFqjlzXzmV31le8JzCr+rfKV
DaUttkrzX9tc20uJMsR6AQAv+VxQ4CNVOzvxkljNBvTt4VS6GjpNS+TpkX52YClk
rlhtYL0uCfgaUj9KnvnwgK9ovxxACq5GjpLuqb3BP5Tlnb3Zel5UzFT2bDVL4QjW
gkj4aMLgjzNA3odyEkOrODaBzTSOJDMuMiYd1stz6yUdqfc1p50Z0GMmX+I/CQ/V
xBUmcxZsuwnRzPecKQnnwYLyjRnNtkVmabSJ07hoPhLj1Fg4imja1MhTr/ZuyEgy
A+LZJ5SSz3JrCMQ5PO4VgLvvR57kLsPYbh6VJeTPQooBjTYd6sXVEWVJEWphTcnO
P4yfQN2eRJEqAOQW01XPUsboKV0Ut1EmHQFRCwgEDYiH38ZAtOJTs1jK6WJ9qolz
3/BORF/fwNwb23JpOt3v4AsoP1+aTt6+mkSPFGPUAGnU1WF0uIEO+84B3oc7A/1c
bT/P0Qv6WVlUzpt/UkZvslFH3WQX+CYaCAgWSdEnnxrr4sEx+YipN5FRO3PeNyUb
MBcUldtlnNEThJNvcXLQFfSBXTTcyfdxil2Z089eGefhOsKgP1CHEENqW6KmCPiE
cERz8ly+PWcg8ir0qHOVzOPgwY4UM9971WF5wWUoljpikRAalypb0GpPS9AAmoBu
/VGqOgGaR4kqAsZmOenwnbiiazvtIDaT6SOamTgY/R1foCtn2NbsLO+r5HchfpHg
J3KLFCd8NNiysEEKSpDCvd2+8LVfWkXfaJywqEDmqdIlcVpVW6R5teJzD+4Kg1Gh
Xk/xvs5zU1ueABjgTZtQFFklWk/aEY3/lWKO2Wc2MVV1FbJF1+0A9Ye8ouGyZDXn
pg03XDfc6a37aVxKkBxDM2D9TCbKnXgzJUZ5h1kjzqMrWbUUPa7uWngCEencxi1M
0VTDQuZxvo4pkrNEJm7ZoVFT5pkHcNuCJoy8XHoZWz8Qd4238vVh0SxeI5wN0v6V
Oh4Tk541LPHJ0D9E5P0abJxeopkp/AsUiEQaMxIlFEYD7wDnHxm95AxttwigxH6q
J8h6Mo1P5JnzI/pB9/tnDeNzyukc3jMnO5LuNW4JhXCkU4Ql6Pgm3hfLRwrhgNPh
HRhy85vDhobxrO4LA3CcBzwU5xtdlAZm8M81XbRArF17k7j1D317YuhDrhTJPoh/
9E83Tvi2Z1J8VdYwirCuNZWQbWEkOrmuHbPGlgXmuMERB2YLdJfsAr9VaN1tguzI
jLUHQMqQuNJcFdEai5nBRVIw4ksrmOwAYxTtCVgoubLXtaYjPIlzhuw3NeLyO9z7
g6RQaQYiYkI1T1N4chONbw2IDDLhPsNfKoeL/qw3dMX1528ZVvOlnm7HmT+JIA/g
s6UNKny87hacgGvt044zmf5N33rdrHXfR5h7l4q1WnplXmPq+nqkY1/k51E5//EM
U0lcBM1dAyR8hpm5jbiLYkZXyU20MMeODyZQF1f18D8Ua8NBvuCPKEJxHqn5VDkf
l1wkJI1B8/9EhWe+1SeJPP9nugpT8UhCcjaBrXotcI2sw5Ve8DXXNTitDh13Btzc
iSw862p4lIRnB2TGsYWEpIXdpL6FLDMsiyB/W4q4A9yvgr0cjHy9h9vjAp13AKQL
xHoVSovVzIy4rewDv9VO4O7d5BSxjSMVVAr77vLoQdnvNM6rSgz1jiYJeKcclLJ8
u07q9wsmK/BowPOnuBuvwMxP7qpayN8LDLKge3qT4M8rtLQCx0YpyvyXC1ErrulW
Y+5YWPN7q2F2Mfo8wWD8H6hvuzOYNQtUSTNSviAe7bkM/eXdKH+vywHeur1hcFL1
TVUH0fSQ79+U0lG5eH37CCyKtccL/MotQvnpqVlHieeHilB1Ayi4ui0aHfNE+VbX
cO/Mkw/gitc1lfqoCI3Yl2uvtLEqxgRKuncS4jAPEvkH1XNelhVeqfQ162p4pYMk
iAqZM2RtXUMho523hv5nxoA6JEk/JPLySsZPa2FN2zeuqqzTF+n+yNhSuAz0agGn
+dR8SNR5cEbMQtP+mOtE5sJ2LGsiJp1nmd7NPIKmXtV/LTEZuapcZOoLjm96r6pP
NdQk/nvsZDe+6lLKG6TuqAnkVrH66pfFr5zFiLLoE+eusdrdgdZoPp+LSP3gCidJ
VdNdlQwb252w+VowBAlSkd8o2hjCNM6UKR0Sv/1P/koJFM+NN4aYlObIRZuYg5n5
jTqIeYDbjMCFS/DshwVj+h4QHRdwZ7nAFsfOTEOg8KD9l0/daehoQZD9x2gY+tCT
q/HazV73pJSz+fQklAC3SUmYh1j7YglJ4ekwv5s6D9xbqqry+LTCRbtggg7ZsjGA
yDyTGTEigAULVGT0E+xN35XlKOdfQY0dLSUfeU/2KhAiEK3KGoO21z/QUefMhIBK
6FFfffsR+5nBJ2BuLVEc48n443ED2xRc0bDQ2Mgr6oULwqrKFAsw7HWJLQVoQ+K5
Fjmj1my49jY6s0OJfV8/JcyGhkZIwvUv6Wx2rTZ0JZpQjXSaDuJ4QbzV4V5WaOBG
o2bX0bvedNR02qVlz/eqB75i5m5HX7fLzTK60eLuKxQgvuxIiTcYvonxYFE2+O/w
xRdxFBygfvkMsNj3cyMlaJnrz00nEQ61f9FUXQxJY+tlbqGNarw6wGP/OmyuX1rJ
f44KZnELmZAS/q3wqkT9ufTt+YFwMA0T9mV29txL0dxIj9raLOGTM2oDVrl2t9UM
TGO5glQo20kbCwRpR8blgUYujV6l/ekE6mmpNuVjr2uIJNAhO8fDoj9pgq3mP+WT
n2Hotv9mB7IfgSg2Gtz/l/gjvMtV2oJYmjCbdhWQJn04xcX248PBbvRFcaQ2ugal
JO6Y81DsQtSKR1DpEJJzUnH+Cem7WCcJrQ9D5u6WcKEkyINRUOYLgLWK7ShjKDb5
REw9CMNcb2r/XMo3NLtry9oyt0HHnTvP3CFKCoKCkdXaSJP+EpLc66Lx6/rsBg09
1qdtNH59RIxB5uzTmuD1hoJ9youzOqwRBeChJ9Tu0SsAad24wBXUjmCB0Qb3ZCfn
M5M9EfTwkTTXWQDktnUt5rspUWcI1xVGeFr6LM3bCmmieKGUuDBxEj2FirxD64p2
STgLJ6/jA4J15oTYJrWVbf4vvmXA2oidiv7F11/5kEH4815BmXshGeBqFV8dHAUw
ZczWqHj8t6xa71FyBGGfKpGtD5b4pL/PFojWh863sb+aT6WTVFq7yq7jcXRqRr/A
IxrAj8NLpjNm/ibAMS3q1Mdgkl1ZvnDi+Jen9ne6wWObtQwPq70PdvgxnJLG8mcW
omWveWLC3OEk1NmB1irOUbsS9C914Uda8SNGvOjGR8wN9lxsiYZbu5HtX7cfoxLx
A0uwaLtOXsOyGRZ+KQzrUCKU0SCYLfEAcGSZcLquhkRm6LgCGFFRy3zV+0dg58j5
+8YPlO3hOyuGATcvChS7kGifC8G9hx4Jz3eHMxc/J8r6Cn9WFUjrlZK1Y3lClkyn
fLyh8Yw/bpGhyiKY57t+xfJJFLM4OqVHq5ozsAW/i9dJWCYeKEsCkQl18+S9UjNd
sT4hG/Rl3jxXYehNHGTicoEGJENUWVjgmvZM9R8ZMEaYhBldeXFcRnqJjFroCgzc
U68FLlFBeJw7GynpG2gmjHBWtf0VnLHWkV9AELSlFlouYU/CBQS876qux08nB7Mm
gsaEbYn6ewCdXvFOtRpv8oSciFNNnMdku00aJaIBIjcdCbHvDYsmksfpzgZsqt0O
xVpgjWFh3Y+7sy3MWrixPbq6yH2AtrdhnAmiAd0bbPtuZJCmx/BHKioCdP2RvJR5
dRsQb/6xtTRcPqk0Z223PJRZ4FBtaDfRBXGnGzGKm3lAi/C4d8fN8DG5kj9+IeEM
Um+YfUm33SaEZmPoRhyrHT5d3FijPmcfIxCGUSnXbO5IKxIIoh+/Lr0+uZFn3Sbv
c0wRAIOxNMYm3Y0jhOd9IQ0SM1uMxJ3sPHovfGXl4Rf3IqY1AHBFr38F+DFbN1jY
yJVXrMT9crxvwgh52cEAgLFigeIncdiPW/eN8xZiYKJeIg+WsVqC+OQQ7n79vlsT
TWKYjHGbZV7zVQJgV85FgGVxJaGKGMCNyt5dsICA1565ZMm5dF+UUS67PZBfsKCb
W6XG9t/RikHpN2uO4RfQr2jWzW+Rc9mo1R0n43EUQwq00xTwEMvAf0/5ZVd1TyEr
c2Xm/TW3SfblO4K/h1upJWuY3vEgPMYhDM+6+d/CuEJcVavIZgW4EEe0kCQU21Zd
ho5CFCv8ILRbN4X0te2qbcO7Qkpa9q00JTS2otnz6FlJh3D0ZRk0cgqs+PRSBBmz
qTmD8yKnDau+ezN/U6w9mz77/88l7TnSkqmXHiE6oSGrebO7HD4cHA1yVCDyiRiA
o9fcSRWoAALoxoQInaf1GsUIP5SaCENtOLgplrcuxQrI7z1HNVi89QOHDG3NZHJZ
U/A8xOcnSMAIDT+srypmSw1yFzOD6c5gK1t1UbF+SvoOGXuHQsWDigwXl1M1MrPF
EGomg3k+RTodrPvaYW/F9YNa+JbxAwfEsaqtcFq+2357QIvz/7N8oVzctwZqci/9
71Yc+cJUiwD3OhahreauAQuhD0FauT3AiK4/3b43Xd/pI+ssYt4LgTGtnzCHH3Gg
ahClFLJYWUEBOHFc/dKa1YjGvU0Iv8FUh/qOZHZyKWU3kljyEv0soPK1T4mOjBWb
j8VG+XHP5YJVIlzrcyvBOijOkEhL5DOYbERdJXh0maLgYEOBUxn3sAgOfs+pgSdN
ZUhnBryP9RAVuzwgF2fEyARjHD9wV9hl/J4TotGM233ciiPLgAHD4u1/7FAyTFxD
kbWy5z2KOfkM3r4Hj8VuhJEC5MZb4up1JOkREQPCzbISRqpXyIzqyxsrnqaMxV0f
KpXfYrLm5DxL+EjOT13XFnXqY4eYpPlv7rXAPXqB7uGZjtPy7KY/HxyBT743UHNM
SMMq9uyhIKsJ1RdRvWM4d2PyAenagHDwH2Tb/DohVeDBHsWgaITYZAB79yr0tTL7
NK0v7NHxXLjdPzo2CtO/4jemLkkwf3syCpLiMaksDOOPrTsTTVJ/JCwSNS7IIGMn
Gt4afxkU9snOBKRBNwvLCQAolYxZY0IsvhExCKnF181hObIF3Ilmwzv1BKPaGvmj
EtgFaQ2aBIPBdiwgQuEyQOAYY6fOlPw8kAqyzYkBknD0bzZGBcQ9v/sTouaBCkjO
mKYD+ZOIX+chPltYaJn9CL6XcYtS4Ug3YQBnhaiMy33/E9VL5c1laNUVpU8AQSw1
ku0n8B+RJmhphXBn3ju2niLM3K5XIWtcBicDwWAIynIHDIlAWrPPF18yMvEuQOgM
M0lHjvRiOzSd+bX9tunE7ibADJEgOKvabz+ukEswu61Q89qqad2ZXgBFfE5L3nYZ
GE6/xsyk4W0W33i/SeGczGT3sJHprvMRiCXlAb1cvtBKOyRTqC6ZyBvROYMjpVzY
viAh35me+gcFgwhlTrhe7n3dM0ZXQF+CpVBFmcP22bbDiJjatHfEfK7kKcYUo+Ay
+nMlV+fyrMdgpY4whG0gaia4qLnf2VHcbsSR4FBH5v5SYMV/y9FsKg0XFfZMG+xK
nZRufG2uM4LDUMzw4R9+xc4vBPMBNqPaI/TZp0OzheJeSZHA4i3NVXXVnSRa5w9U
xrVByzRAQ9HzDrkSxlnapMmRGjAMSUklcHigmrGb3b9MshVan3TYT0oO86GBQpOc
dD/ErCHutffSstBAijbhJo1xBtVLYMiPIWVd5j3RSSOTiBRQQP9m44Mm1X9/mn0n
pSwI6X/iVOG5xPYRQjfz1erTv1yny8YWF8g1XyY1sKvEbOAEqSGTDMefBrjKKBrh
J/6I5a4Hx9tO8JD0na8wgIVt99jlVaLQZSTMYplgaSW5fTkrzcaw7Zy/YISnezfQ
xafl6tgnafgNS5ZqCZuCroCdxjkbFAxkL3Lg2AOmDdqibRJnfXrxWURVLl4rvttQ
2iMiBirIQhwpN6cnuomIdqrpSG9AFjpoZKYFntzWXpd68qSjNJcyIX89t0j/bC7b
ZzDQhpXAsWF3nch6GjGTLoIK0PnCNAUvMuTUC5HoK1vCSH9gzLcHgXDv1Aja6FnO
At5zWQ0J1ahE/kZ+3tP9Se81nCldzxPKo0vQQb0cXGIsYCveysMoW1FnS4HNmzn+
YK5jxymtXoVcv/Vs9r5VasrrFWPUBdC3X2kgxHzGamYXMhTmdczQlHTfcq5KW2qP
eeI63TspuDx9Qr124eKSLpYWsh6Jxui5FuL2ZoF/bpjiLkMRfC4CuYsqlUU+3dBg
OpZ2ZTT7SCRD9p0QmC5nzz1pBakds4/gQIuOb7aOB7/dLKTOEDStEcB1guJuwT9b
N/NN3Y3zoiJlhKEvEW8vqRqkfBMEUmZmnvKPhlgkMBcwhX96KiSVkluIiNRZ43a8
u5gMvsl5Oy9RGK8yMWduFnFuZdJkIiIDhgvxjQXyEmo+D6xpMs94L4bF5/GweP7I
RtcipZutbDGaUFqU99zgPJ4c3rX0Ka7GdOA5vZ0c39YiWTGrAVwuFI+pviCCMk7f
2NDV2LpdNH30JnzUuCPUqPQzilBQanCHhiFfQflCAtJVJL+R1QVkwEbXqziitabP
M+L7kkWQRWPMjXNb7jzsBdtwNdCxKWTYe2q+n5LtdN72MadjhNwDG1YgV2p3XjEz
4N1K4ktfs33uFUVqZRRXh92qmQ4/37W1mtpDkvymUWlpo0D5EiE7MiZSu1F8r7U9
sl5whPhVer3VNaP/1DkPe36nI3TQhKs1JO37uPdwmOBOb3+ygLHzvUKE7ecXq0OS
kdNxAq1HpwL64INWfOOiVEyaxBt3bGONn/N9osZdngM8x/e1o2vJzqHpBVcW+yaz
4VOWzrZ7bhprqnTRjSSrKsHoBfoGJVR09xlrr1c2HzVg8gEfGZ87AUSceHukb4Vp
nR6xXpNhZGnwIG2yajKvn5mFyVYagzy4F+lJGGsCZIglig5XfJov/WtXVUIuXe7d
YdqT78PcC5QdcvyWyVZx5v8rfqo9/MuvFr+ZQ1rbFexUQKKCf411F8R3M6bSWMEG
tJ1PWdAJ6DZ/PZWn6Frt3IovV8yTyE6K5AQ98pgvhz2yNZHH12m+1BKFHiGTfffB
p3sUmej5McZ0dHbvyWNwnnFiDH1hGVdahSan5VqB3GI3VPOYrOp4ltA8H0+89DU/
EkDju30unZZItosWRWnsnkjr6E6zJG+IDKGb2dEfPWgondNilg9qZ+HVzqTbRRd4
QwWE1tZOZkJVAcLIN7PZiDDBK/y42iRuSeTdXBTS3HhxgKx+1VSMVQCoPz0BQsR0
gFcIxWdl2L+9iyq7bit5MXa7V7TsqmJIkvGUtXohRF9yeh3r/aaNWbsQEx/v4DEC
+/t9463bzAkj7H/x+KthRP9obbFTYXMh2csQjnDB1Zw9/C41xNnf57YU+/WObev/
0ryR8VL+aDZX2do48jA3jSOsNpNsLhV87mmKUhpGVv6d+jnUjar2s2kvBbUp5fjx
V9UIGq+yS+4oh5u9zJXZ3BJPn6G5ehrmyj9sW1UjAkwLnJd2tM4mquVeFW50xh0o
5tvcaLZSDkMYKOabAm1Pq56p16GL37LQi2zF9iX6vbCSGas+vl2o0ggapDm1S2Yy
CTbaTGoRgwin7PJTx+HfrmORvxdpbuOJamVFKBTLAEjZp4vHrNuWqYxFmv859RLp
zPXVJ3giuHrVfcnOwhjo849+u5ycTPu4/T+wgOlRyg8NL6Njim2zUTJV7eS5nd3t
stH7tHHZcWi4UxzYkGuiNrp65NBhaS+lDBKd3q5aWlaYQ90a5Tm3AAc9Twt68gzz
OtxvM1c3/OMfUVYjMBZKHV97UT0SViZm70ATT6GBcI9qiDcbLN3m3+/n/HfUAXga
mMDkiW+5INTcN/goJZRcaSBYF5pSh+mwZFKrTepOc3HJxc3B9SiMYtyPyJhbXqLT
A9BJBiKbRNb6/UQfgM/uV0y+03D5usoGUFdaKFUhhqbGGeMHLxYCVJQRw9sM4YNr
/FBtb+dK5zL3i8vyVXXW4J+E2hzXyuevzZXefL2BKKCPDwzAY/Af20zORmYdDMCp
Lk8f5bXwlw9MDrJ2GGti7EQ7aVDy7EEKIIXBkX0UMmc/DitM6ixjxEGB7mUsNtLB
lg6F3vL32nO8QrK+guxNx3bQWgem4CdH1BJb/UsNOLBj8WcatG6NyfhC8469spuv
ud6iiTcSkMUGX9HOU6chz6A0yZ0eCUQAvMHkkiMRNE8gg42/PZ8xBaKFam/Xmeev
N1Emcc/DCKp7lSDbiF04F/haEgbPrQVkMZR+VvjTckkkfV2IZ6DiLsxZTBJgZbtd
kHeRPUaA6fu7/GDw+BGjWRhooD3gaRtk7YmSa6u2RvuEif7xH7F7MzXQg3rurVW8
Q3wmuoa7Rghxqsfph4kKaFpFhlynF28XmTIAjc1YzNR99bg7hZyGvruRAw+wRmro
N1CmQh+pSptg5sKqQSz63TQd2rs5hzfK3b+HnN9bB6DHRDxqJouTn5eC84McUw2W
TRjvlbxz7LBIuIqTAftCo506gJKO+Yl9PMTq5m5tDjbsVp4Hk3/tPk03GfAOJuuD
YPQung6PObtd9pZx0krwlPaCJCo+g+9oJ8Qi9VJVimisEfyiwxeHkR5m136TlmhR
fyU7xZJTKNVCL6gkiAmSFvbmNgiPW9YpUngbayb6cl6nVuCfkEBaN/TAx5yiJ6SA
qXOohakFDu2S6TpyBkDAZah1sPasjylq+sJheRUNtU9JnvDQdTzkHa/MKDSQME7v
wBGB4KlQiRfUZ8kEEBtWiBxRGHdT3XE6qstO83Nxl2Ec41tWmH/0tDc1FpH5i8TK
q2FQGs5gZf5Rz5y65lMYuSL/QsHPL/8vqtXRYurjBJYhW+SswLfhDIaU07Ql4E46
1iNtWUvsyZhLWkeyxojDLKI9H/2KOYxSIQeo9uL0MoaSF0kY/Ikl4FAIaHTUG3RR
HhV+sf0AbJ4IP3Wzp7zpYg11b/SKQtFkvxbX/JoLkNMAuS9P6Xpl1KPk4UZB3P2f
P3TWS3KDczkjV6sNriMJMR6nfpk2VMjsYquLGURslSzCjE/q1qzrESjui+QFqWRK
olt47sr5b+6pGgy0dc3fmMXYMfONyXBQUUxZC+t4Hmxlx52bYMroH+MFXlWrHPCS
Xnr6OBezoGRVi6flkNBTlecG/1sODeD1TnEw08WWOsDHHMEeVL4N9XahHbrtu3Sw
uKe/b6HsXQMLaBlwk+0mn0gORrajyQy3VoBtbq4zS0O5iWwAvHIs9wntOZBD6t+G
xdZQnZ86pU7ELSwnxzDdMCS3QNcb1zDgqDn50CoB8rS9ZERRKAqVAp9ZnxzGt0Ov
CZN3x5h0I8iXdDW34fKVpK+s3XTJs2XxJWG0lXPVcNgFHmBxl/mGJmmx81cNWcLw
CEBaC3iIftbaurnhmzJPXBfw0sOsrmF3hYKDfEv2DUWAApTrjTC+IXiQnHzAx25s
8N2R6TEC9U3ZsqfhapvDjJgYfLS7b/bDUG0AwL8sc5PqoyaHbxVn2+6AZzcLEzmP
0B5+3TXynsBSSvLhopeXbdJKt2rcidhUet1b3DkV24Sx0qkO2OIsKjxId4152wnO
OQaYp7U7PVJoMnRG/QKgAZFRHd7oTFJTxmxx6LkPIzw7YnAO/00N4pmvy3jzGyjq
jfMj36mzjbX1L+D7BrtNruVfdwRlkXOlyQ92DOGbylsBmIj4CBv7qK9ZZK/W+yl1
fQ3xkdzeIkna2uIGz5LwED6Xr1In8MqDNAPG+cNHFOc3XYd2Bc0doZh4YAXwu2yu
CSGJJ0dG9GwbAcvKeSMWtQsYR6wUsDy310vBKMVfDlTv7D1kqugOJe429MJ88OCZ
MrBOrsxkHt0W6BhjfLeNhjiaK5l6/B284xFzhsiAWT9hmikodgmd4e2c+BVERtnH
k7Y6ssC8XUarE1yEL4Hh3+02VcVlGi4NjY4MFHA6IR/76EwRXMnx/J1yto09Wmqs
CK/FiXx/tvr+jlhlBrtFENvFVd/qy0YMowThQgpJYyl4JhI1izmJLVP3XGHUfDTo
g3JVLcrN8TCTsM3zsf9RfwmvrtarvsHth5PrMSFm/V1Xp3DkLL9ZoVPHgIBWhhaE
BN27fOdy+XgtY8ftr8ZweZ6ROBh/zqivzu/PM98uKVs313wToQVMWmItcTgVT5wI
dWBIznVVbqJ/hbBhFmBZmLM69yt4zLsYsYL+6FmcAWM8aYBATai4FxIakSraLuUC
bnOH4WqVLagw2wJZycNJ2MplncRu88e72B3DMgrUdWG1zJNObeF7FJFjx6WKZ8nb
GEBaPzzLtfQzXodwq5LApKe7EyDhrL6ovgsqaDCPIqCO4mjJkwg1jvjTks2JojdX
5DF+bPgIkSFdG9TR8zGbfltHxlAECczph5Iyx0TV71oBPI1KvyxhHm0Ojc0kG0/J
Rzj+FfCV+vcuHitDIf4/qVHevX6mODyG5++EPCpXIwKf8BYjYWa6XlCiXY4nztby
+ax924Z56X6ZO5YdaSh7Pbvl6Gw09blmxbj5M0nM0iyJeStmz33HRuHPnTdqMTS8
oEciAZiZdjZpaw8+f/XPD6moMLIebu2GVL8wKquxY95NhqPFOaKb9v4Occs/Xd+F
M2coNRgYfHzDKLo/ry91Gt/vuxEkxX8IDg8NJve8CE6HqU7SxDS27QVOYjpfKcsf
8z+YKrMzUhUb9ULxOMqvueyT78K9Xt/YIYtM1eHPxDoJlGG8GgI0rqmIMtso0GKv
Wjg2JdlFIT1vST9GTGtpTKdtuJCQ0/qqMTINF5lHGGhudJ3siQHd+Vi+Yi1FhLeI
OEhpq3087eqEpYAMbqLnWqof8ojeTXvQi4slKKAz3Td8M0P+MM7z9zhPXiC6R9wX
ok9FgMlARrJgIKmUdJECNlurKtI7mgjGapIi0Nv3zdyCcpeiWtjlaThb5NqEh6vy
3JQI4Ufn3enxA/v3iunX3GmZa3fGVbIcr2skjYv60qV8ps5som6L0y/jr7s1gY9O
nLJj1Q6MgMZ8AMwy93nz9nd8rQ/uXXsmYtAQnq9CffSTlnooFjAui5NFZ3TnnpzX
XyduLi3c92NEGUfS46YGIR171AWqNkTJ0ht3J+q/FHgoLmbrGSgCuWIjY2bPrYgM
q9llPAS9thlFBM8Pp/nBT38+M4BDNI/kvb1Ihj8INHOxO70c6ZcFh9PJf6UJ0v1i
XprgqlR5mkeK5Drym3UBvOO1/c6iwhU+EPQvn50/SD7isOgHGebb2V3umCRmX/fe
3bvCaDb2zP0ewx0+LzDntEnnp6lDAtoWusfnV4gwF+gynXd5K/2Sq9cUf2vzKb2U
TFBcgkQ5RS/Sn07VWM6Ee+m86EO4r3dwB11Ifqusi4Wg348MW09KpgzW0lEUt/4v
mI8r7kRjO46Fp+RDwHI1kFZNDQ0GFPEHncDXE7lBROvn/zAAFf9pksNb2VNTkvk4
pcAuJgDJCWVPt2xFLWDu4/0816k7sWLZCBaSHXk8W2S8F+ZlZXTbpyNuVquMH+sA
nHz7CZ7n3bpDysS1i4fivV+rS4ZYg/JshFhzm9vra+9LPQiBoaK4wjfOeD8t2WZ7
NTxUkYU4ioCUY8j2ErWv9bdihN4+J1tRR3MsLZO/HFft/1E8YwFDDtrI3nYUS2A6
+Carkvq45DUQ3KQEWQBqvRHvwZF0o1Cd9uH24qmSFA48coFVPmRxBBkR2JSAz3gz
O+R9qNS5+bXxx/WzHKlwMaqO7fvrbECVSIB2rI7ZbX9HlbJRFVSHR/ulX4nslnTo
kSx1c3JzTmkTjTKXJqHx+r5BwB5b0PLjTQ721r66WClMy6WUiplC4Stm2hWBC5/D
RBBnybHs6hZ7d6SDc5+bHey9IilUGfnRgLhvXp9p7UBBZ/GS2CZeOTLCyVUM6FMk
gUiQ7UCrTujQFzdX8Rp+VHuepoeNxRs2UHqA+8sy1gYdiqYIHWhtqZnBgKHNdEcu
OaQlDolQxqUmZ6xfKv4pCyEPL1cEPTQKgKRqnpYStAhmc/96qB5YtYclyteqJPd8
22xW6XcOMrJPiZTykz4jCiT9gwwk3F31k39HHcRNuOgETFJN/U6omIGAshcXC0ZP
+VkSc21hCvq40TxP1kypkHLG+m14eL9Utx/arATOBo/y/EIrg4cYcFtcS+mGjKD+
GRL9oAbhr/h7ml+yTgK76vq4Nd+7edb/1OX97G29dXdm1j/QuQi0W4UBjsTKkXQc
UbWPR/KFRXNnZE4oYTZZPejdI4EJpLAKxyIwlq2vKcGe4/GHnD5RVAnTytKc5iXN
MZQ1vSMb0+Qyx0CxWOe0oELrpiNjZmI37XNJkv53k48mUWAnRgKDzrIJuyLQRshK
FvaPZuD6sgJBSI9lxO1NDeR2dNXEBQYmSR09cmkQM1fxwyrArhwD0z9cuUBzvI5y
dCgAlL3dWvizJmiyiJqKjCqaSLGC3cSbzjj73e5o97YJZHpLrGmy6apQY7qb60/8
BPce69GabNeu7rfGgQsVsPGjItEY6PmQe88nBoZ3lMbLDHRjvWCY3XOWY3mzUQPn
2JwR14fodJurllkkJWqPKxXt0N7Oa8twIUax9Syrh6giv3v8crEEGb7kOHW/V71C
pxYeQbPVumAc7Pxq9QcNGNCdreDMCk8PwZfVgy7f8TUTliQ3ygvOcZYPa0zlTZo3
3/WeUjP/2ufsrgkoA+hkfKXGN/vjI4mdKzASz7m23T6E/5bcBzlpll8gZ4aP3zWw
/kAwhSTL7Co6hms8J+OBuwHEe55+X4KjHGPC+rtWglXrMQfpUghKiVDxy4k4yX0h
BDGjxD5oRiP955JCUgYHsO130QaKxgXBZpFoMQo7sduM6JaPKns+l9Kk0oa3kzbA
iMTctr+og7ftm+OttyuffUGTl95NnzQOpgHi47kMGsGmSWf/CLgzoig0OqCBI/0N
g0KdnQJOxecB6/hRF8ALwQUK9aIeK5WmBmnvvyARrLKwgROvMDdX5XWhNhn6e6mu
bsXbF1MwxAvAU9irptEEZxdbTHMQDo65K9FO7zummEdrXOEpaejwgIHphucSVksA
HgIfROWm+G7u8Htb3XmcVktV+2sAzqCfT/iOwJu5TZvWN1YkY7g/UOo5JiiZs9Rz
P4dRXcsbwCreYaCVhKGp2gNIEwDqRTV2but4jRz2XiVX4KssirpmCjQ1X1PyebJQ
MztM2zlzZM5Xbr04I15jdHFyAAe58vbFPycjGxS0cBCJIiqQ4zibCftlPSZOz0M1
f+4y//Sw0DuPNW4YxBlQ8M/M43eu44FVDbwxepS7PPCMVa8kN6LemBxbt9U0QCmW
EmdLmnTXFfd0jBEz0NMOaTb428nJaGYX7If1pO0TaDfuSFOcAXzXFeRVfNF62HKe
MZHrVMmzESB8Wrh4OJTzWrvyySgwNcL3Ia5L9gKLodiAZ9xXyZpqz46NuaAphrJb
svF+brpkK+ZXxzDIMVmcp0IAaPnwH2o2rAPKApGR8k6P1eYImKlUub4/kVziXk6p
Vm9giLGGQKff5ZrQNamtQ3kjukdoD5RlMpin1AUZr+mxmSrVXCv9Kk/ri8ce1vyO
11cQIanTd+gcOiVVNUta/V6EPgsV9JKibhBgJ9tozw8cwx05Q0NPTIHh0BhJ2+N7
dVnVMBq5Bjhk8/C1a1v4INp3s4EM1/1UmaAiGKemFmzWXnx84qB4aRTSYKYmER4Y
FOwDuirQFskMd284sw2XNiMKF+wz0rS8iLjQMD+5bi/PbRhZN914zL1cZOcouWwt
NqcXVSJi+ZAAQvJzhiaceyRZ3IXrMIFitQsNwJXJ7tTvas/TnLtLqKenVIHPGSVs
4h3gNn1Iu9FOw4LLudvHIA2E85P3BkSrVWpR+/t6uM5NcFBN01ZLZkdXDp1yi6Z7
lyQGm2sj/yE3CUYzqHbRDXwuGscvnsOfS2XpNZ0yi8C5Jj+1313E0eTXE09MogGN
ubDZEahmX0qQxta9NCDnl4plCRD81JicKmGaE0PmkTpoBnmBDboHbUXjNA/Qf5ff
YxSHwOqjJdljXUsrcJJx5z/cGw3fKzIPQcKKDXvZT17I96qoOjaCuVKi4wzxn8v+
8fIHyelS0pmXAWFddpOEIDFMTqieA7Wy2V+E+PAHa64i7cjf6aSEMnTknlZeB5ii
sCEO/chQpUg56HuASMH6ryequ8ZYWnX0yi8fqS+twqFsMg6Dgorl6prJVJQJlov0
NbAeNrdgdcKoSrzmvgg4IcrbQ2m0oiNsNu6xv+OMeFegnKI1DIMp53AFjlRl+41v
K53RcAW1/bbpCHkIeO2d+quS9/IO73enCN82UsUhywoG2e7fK+bI5qy1Q/r5HNd5
4GFqcxndWE+SPMo+YzX3Zce5b2ua6gogv72Wj5rtS7dWpZdaGKcDYgVEnb2ybGIV
hJf2Lvg6XvcnSKEFp5n6jffsD1aLnI3dVKVEwcvPeexur1BUxgmeLatwJSF8rTLP
muJ05nyFPnaI90UNyGF+kc5/a553sjY1PkWy5KxI2BbRcV90C8wVeyVm4vLIYBbu
dkvBa6fSHjdMqHvjbBTqx/Ett81VJgpIm10Bb/wqQD8ajC225l/T+WpVCEv9OISl
L4TZ9sAyFsC7HWWacl9d7ydzD3A36d9r2d7CtXRo450BoSBrG3gfcpCaI3fDWIky
+SAp8XU/en/gB1F/2jdf0RZscwtOzfiIs6cd8w+kORbb61aNiA0clec30Ku19F7g
5A9azHePVWs7H5spFXWwodLODHUL6pFT/jSAqariSVPNwhT4OzdiNbF/CMbPh+h5
fXFG3MDqXatLIYfxr+T0GKEqRlPiNvwU67jOBIHXLZOU/g+NSWnPsuBXJq3HfugJ
xxCUaJcfP2GoHfrJx9xioZ01SPJCj+unJCrI7Fh8gyPvODuMqW/1EXpOusD/zjme
3d0qi1hyEL5ioAzrtkhykFYXO38sWIIYoGbBwSHodpdE99MesJpa56u+v3DdMh1A
kIsp+1T/hOVFqRL+ocJlviwaQc6b/oL9E2xvb8QbGlAXn9/kx3ftqyW9nAMQ4eXs
NSMZcrLlO2XQfPlIj3oam9sjr7rfoAHh2jMpfRAZSDtyQxeqprxaVFvDS5tBi0dY
jsvNHHEw4Ij1n8/OKxYZ7LJYfHppnFlB7PoR7jBtx29zilfx4PC2zzwJG3k09rvu
XxaEOScajNpdJIg029V7Cg8cwvL8f9n9+PnRCorf626exAmhjzZvXUy55ij6Pj6p
nPV/Dkk7EwsWyywc86yC7NV68bAV2B0yQr6CHDqhTTek7cujDPhyZGm5FJnQx8Nl
0nThV17xhigzMClSBBUZmno/a7WsYHb85AFKDnnLA+a2W7QTSfI4s+1J42VH1zMD
EKGIU+NWSKiU7f5ugjNjTz9sh9pP8tNdg2clMG2jW9BHo0TGeD9RaTNxek6hKY1U
KIYZflqspTnxWkT8hHjjBCSnksP05jcdBJIRqelypAnm3ek9rONSvIVxcRzfmtYc
KGwz9CTEsHHJfylubjxyGTwRrjASY/pUedn8ucDeJ6jFYfYP+vQbw3bEgUP+XKxy
6xbeuaYHCvOqr7skEYFnGjxmau7BGSHRuzCTlmxLfqnl3I7MnqDh4SMvGhtHbggp
IMHjdnK95GLfamstV7Ysos/gZaQhpbJwa4e6vbU+yYivZLFb6FZi+tNLCQyk7P+k
Q4qYjBkL6tN2ZNjnvErWt6u5HAMpcWAH7blaRitaZHMgRG1Kr1eql41hMU7MrTvO
3JVPD/armzfPXDVpVIRX5MsDhrVoDheWtzWVeILP7uSjYIXOVGK2/GCTGftk1yMh
Q0aCmBpa6jx14hU26XTcrb21tK4jfPe6fxjD0jQONQ4NFIf3brLx6CmDbj2TOQkx
scHOhhXo0C7IoztlxD6appO+Mr/ZMPg80bbAqaCYk1WiaYxysWpMLKITtoQzWejN
dDwt2ydvw8PZmJ4kEmrYGkIPQVLowkYJZjzyhLU6byJ7J1Urvgw0xD2d41AO5YxD
Hg39Oth7L19TDSbyCiGEK6/3EgS/ciwN9IBVP0BmBKYQd6+xJRVRiNnrgWKepyJl
F3oOKfd5Y0897SKoyuR7HTRKpapZn7sADFzcRKpVKweDQC53DlUCeyehVVfPbFnP
eR0WSznRUMeyg+Owq9iKHK8rwV28wjw0f0LNMAkEHpQmPp4sB1QjC4VQiRlM7XJI
vTbi5UnvqbM3Y8Cz1zL/UrJCWY/Pllx/l7GE080FJkjymJH09Kuxh0oBoImhl21L
hYV07vH9SrTosdQu49bO7UGOa1EAldwnbtkhYQeLGa5leYXaT0OTaUcatSdhuKfv
XSsVGVlQsFC6z5ycImf254ETS1mtoCEMiQnSMqoANjF8t9hkfPAXYRxHEdeALCYK
ZmjZqD7/rPcxSqLy7LmxmgNkhXZ+nwvU9GP/BOND49rcZQPoz6VLNwKO4MouvcDv
W5cSjDk6Mj4jC0iTDnvTTl12j8+42T3uD6lH/CDmwQYX1xHNi9HYaSDtcKggWTjZ
QBY58QEa7mTKRg1XaygQiwWpWf/zErSI2OQ66cS7/hMk4evjVwlqATbt+0HGNdte
BpBT/G4WpL8pm6/U3VjmuZAvSiw6+jbSO8Sg69Fy16G60WjkNo8HMlJcbsNX3UKs
ICLkBgNtoshA+GoXZcx5GP3CyQpx7Erm6bhaWuGiLa8Qm28O7FMi6LRnclU8N1EL
RQ9j7kuMpInVQoCHg5OGtWQerLJtF9NyvT3podGhW6ciO18vTZqHy2iHk9Yyn3Yx
ssWXzz28KL8RXF1EI8La18boQFVTnqM1HUHbu8hUmtSkav3eigOGdGmFxuF2XBw5
vWefaIVNrpBLj/q18EE0S/XcAiDRSEVqTXR+8QYuul8tWyQP890EJPfGi0Y2X1x4
oBLjSWmQbfa/Bqi2nGa1IRNio953sxXVpWdSm96qex3olyz3Sq+IXQuO85qUDg+5
4d3LY4WPfXkyEqmnl/Ir4DSm4f3a8ZzdFslRGZTXTD59PCaBTZcTEwvQQ0ieh8om
Hi4kG9xYZX6tDwS4ILc58CxjjGX66kk1qTaGKmDODEaZRlQUgB/axpnZgclxrpYI
fEdP1MqKMNfpu0+WQCqmhJXIr3+rgsvdVwVDq+su/7MhMKt2w6ZMSq4gwt3tL4LH
J7dgJqCljNLxW488sIPkg7ZSjrtSmMjzx2CxAWdNNhzchsOx++k/oMXVHsNLQ27t
pzclXh38OphAAPLym2uegY7c0FsjFUoWro9R7cwd2G+qMAitbbsqr30ARyshINp5
GVatCBrUCRXvblTeIVmlcme/FxYN5afFSXaYLnaTbqkCMb8ajGsNFjPz7Ib3kF+3
4b55+bGq/IVlzIXFyYfSuGnHvAaAiFw898m3+3DKvMlPEOC7WxKESLBL5fkqtHy6
eo7SwHRgoyF5WKXz8Qt+BYCQ//lOrQ6mopahYX1NNkzO5X2NRxmxaXhiE8ZWPgrB
iaYwClFExLL9oEtJz4US7Ga1gUZOnr4GqJzfQB3nGCcqAvGxIBr2jvAEKNMfmDVq
6Z9UZPLMqfKUK1uRJHbp17wmLQst6dMWbOkqKs0ffxDrw3sSKh5CXn4K3eH1FceR
8ifnFrYUwCMA8+Gu+zjfRH21Bq/pAydjIc3/e+moKVzkHK8alSsrLERmrZH0ovVV
CPfuM8mmejHXQ/x5hX1gLyFUZZCR7nNdYmwkESkkr6FnHxuxY5CJ/QbHzvBPzIdX
pJ5BPTVICbgDBFKDF/nKgeYtlve665aEs+CX9rJcHhEzQrHv43mh2TIBAJ7ga1Rf
phgcvmir44V1/V0uc9WIbj5Az8uDgd1Qf/CTgsiCNg3ERzuag3XUGyI0aJ8Tz/LX
CIv/5hi3+qFZ1Dx1BEo8fhnkA+jpuqN7mB9WSxLGqCk6Ds9xBgOnZb8ytRtWIMfz
8CEDXUj6JY7Bn38vKMqxfKauql/UdDtS52kq3U6SGVb7dzmhhNRCw/ZuZCTikYY0
VDFke3Koq1f21ik3UZOaOLmBAmJEKvJ1j4tIP+XlFeOtYWJcKkqbmcmZHEercB6W
keIkY0NzT7OEHeyBB8UwL78wH6vHByoKIuEOiPvvtfhdT+VYWJiS9U92TfFxXxyb
UYzHFP+UMNV3DHrjoPhbq+UEUrUdnd+uQLzL262ZtqS2/PRo2bpULTFmOd7FD1TG
bHruzg6aECCH9vQlOLuDWYwUZ/4dEqA5gnsJgrLr+CvHproPZJBD7mNQXFM78g3W
ZC301mrfu54Wq3/7h6pnN1gqw0WaeHvJG9ib8prG1DtwuY266mZy+HLm7v+kMH2o
bBpz95BLCfR/scYqI7ttqWqAbtauyIkwqOl4sn7aK2kH/O+t4kqJ6gozjDAny5RC
hq4rKsY7iUnc8tE6z/Ri2GezBrKCkaMdhamh9j2BHjLmtJVqwPu0xvrC1nkYOFe4
jCEj92K7iJRI9HXObxkSIYVReh4HoMILUokNJ0g17MDkqG+kUSPEf79Oe9bqe9Pg
ZxQXFxWog402m2Dp16htZRU7dyOvwHtSOJ2Skg7x1Eam9y7GDcE1dvUUj3VB1Kpi
BZrIHUz6EMxMNWS1rZpT5q9q+JeD9LfzbgXfrLnlLYBFuTnEq3sFeXxS8Q0yApAf
9Y2onNR/4jYtfm9JI0wI9WC38p7oCx8LLn9mwza5k77HY8ulkOasD6WSYDLMsgrg
n5Q4mhsbECqourGhdIMoK2pFbbwGLE25z6PGYchpR8/WpqNb6e/IvXxirD51pP0d
d03lJ9K5PtR/qDh2I7bRvY3JhWQUboQ3zGgZYwL4HDcNC9y3JpXPc8zzhPjXyZaj
TywXFqlidF/qSUYq+25KjQA44HCZCxbCCAFeWsS/hvCQuJX6uJ9L+O9WbNyOpChr
9CyKEf11SFWJ+0KIGOOjPfmfallhjPXEscfeC+YF7eEyDpwLx2LrmepJbyKwQgc6
k38VkYx2OhjaCSph7QNyOHJYQ03dl5YBpSQG4TNOqHtiRPmf5N7Z7UZC8TE6hiF7
asSxDBMN0Ie2UC51qF5ztWJX0VKKi2SevjoolvUBSxd7RYKBamBKtQgrhtdoqLpg
1YaRlcv+Aj/8TZboIUiFN3Pu9hC3i3TZYfM93D1C2QICkkEF0l9Xue9ss0Qv0usG
NgU+cLNKyJPsuoBkAPSlzT6G0DybYfDv0dZqWj8b8VqtV1iytZPahrhFs/lOZ/p/
3Yq3qLSov00l5ChgcvyoRJrGb1lNWmIxZWUHN/7W3cgv3sWF71vwv0kG6LxFrCyX
I8Zdf50EPYzKS8nFghuScZN0sZhkZwpTwxy413euev3ZCW5tjcSWIU0WmvqKfxfL
6pXlKMWy+nIjdMzSfn8eIJnyr2rRhLzQbI6QuvWaQkTqZO6Kef3RZTq5yn/oh4vQ
vAtHSJp+R+jIJKbP4t7QiTf8j9nBV3GRIK4UkTwoghrjoOPIHQxqyCLb5KO96Wzq
0KX9NY/mxoMvjxUDUwETyXn5Z+uThdR+OiFNWh3Ra/21vinQlrGzial4tNp8G7Ws
mwHSjYZhgp5HnYVGkfjKBqdTKoTLfk3VWKB5RK4Dv7BO3Ik/oJFvoLJDFX8VnxdW
+nPKgFmqWcU4NKtP9GKvpdePCcW4pNMJMea3I8KvQwtuifEVAyxErvrXLzACBcHU
50eBAZ6GryfIHEBJQoBtZ3DfIWdGGPAmAkOcQs8Z7Cm+ke2rHUhVrb0Hvl7y2yYB
E+m/t+yleeUFQdqDTQW/AJd5MQH6y2dGh2w6cUP/ZuaYQSyoBvix6erpqahNF682
TyCb2XKDAgdNIPrHwq4FVSpOeopzsYv0NZJsn8bwyW4pjdBlk0Px5/7953jQFNfS
KHERMrJqJdX0bESEXsETqneNpCt+f/p6NMUTvHR/uM3RXi1d4kDH7IJVjjwyjfMq
oRO5e/+305xDTppREPmqG/G9RjXDXVMwrUhiGd4cqyjsr0wmCM1qTqtNMUn/GKiz
zaC/JrXz2CJmQ+D7HABOkEGfyVr+HbkI7+2nAsn1AwIbJ4fkum84aDEJMqlpG76e
O6qJOGFuedhtZH7lCDO3y30rVclJtANn1z4uR48fRWTt/e60x2xt1rNwywDUwc4i
P1U2Tt5XQyoQ0fp/0yt18vJeUJwgEydw2pvo1b32aRfQB/1BazPTI6Lz1M2n/LCZ
Atl5g0184s/kZi4oRCo4CQ13z/ha4yWe0mzSlE/vHmxZHtB1Kg0lbWoI4A77sBUA
VpL0ua+HDLNP/K/11wc1MZt1fU5puhL3x7J5gLFFdUgpU39xU05HkpSvGb5MQTOG
sAcHOIFvuDYCdY14c7wNOYpkTK8p618APIh3xbsFNT3dJerYLIE9nFpl4Lk8Hdue
mvflsWxkbJ8Jk1gOVo0qtB0ZVZ0ZIvuKrtQD2E/XIIrdXLVBSNuPZ3Xvl1SjK+V5
prfyg1YiMCBtZQbkvhPTiQIVAXZzDVQyjDFiXoBYJjFGQ9Gb8qLfQbguP7uwLLxO
dsDEs5MG/VS/QfxkDUahBO4RtxnU2wipCSJHAemyK1zt9fYg0Fit0lYJMht3kVBu
w4bxkm2i084NtDKUt2dcdW+CJ8uql54vIPc7PPLwDwMgNITak2CzUIHI0DiHN6WI
heYsQiXW5bJzsnnx7ZT03anwJzHq2k6g8T3OWLck/vZr9gh+HnmpSkpRQjsnFn+I
YpQFPTAqVjNqNkeWzX7TFXqoxUusjoUVDyuo1i/6+pIQa4FSHIxTOwBJ4ZNy9/iO
up8P0JbepWR7iiEfqwFqRdQkDWKw8psmRHCPVWQtRpJEO25H/7t/6fM59j6aldad
+KS9vSngroqCpaHDXqygEMJj/kuHK0/KPUixLTZgLjaSn6rXZ6U1CfVFEKAdf4+o
8xt4v/uqv1qQuSG1w9F83wFmKaL9lpAH4VvuHxtPwsGyOUl350vpAN1FhEjLeaY+
lIV2S6jlB5YE8FwVtCwr4IK18ph4RJY8LucXU2tBlRLz7jtwZunUBUN8+7KLPF0L
nbWJmF6LXmaTYCZ3vuwsmsboPv6xIY0IKs5wPUphZi2zdrYt4hhWgkXIRnBogEgl
T9AIMsjDnBMSF18yocxyzmgEDJwm6E/WRveo5a7ceOvpJW0b3XrCqqBN4HBdTtp9
ash7YNP/ANbiprWfTBpo8suuNrLFD8W2KmN2mEGG4ZP5c3nh8F/Nzv01rvTIltl5
+6DrNIR+jskAiY04TPLO7wAcjZsvHEMQ4g5JDr8PflZLOcJH6rgt1w+5EQND8MB2
JTj0Vu76hyBLAVfLxR/ywLpbxBgeR+GOCIMNSsIBLdysP4BZXSGeWPLhG6uOQmeU
tHRh8qChMwkXk+wWYFw0QXaSpeRfbWu44Avi8SkoLIFXcxpWA5OuKq1t22XPyjuC
LkTa8CTiTj+DjUJxI4lY38Uu9K3k72UKdv11n5AIDfwGwwz8+2QYZYMkon4JJY+V
l0weXRjECt3I+IelL3gJXowVN14P20JJRuuErfHRezvj5HVcyd8rN7qOymk0pwTx
hgJ+XtsD95+ZLntYQXev24/bncB7P1fD7t97Ijox62yEzx0Zsegj2w5p5Tv+WqPG
SQUgywC0Vu4wJYH4RRXPsBTxEMKFso4w+FuSkbKJk2WtSyjPe1aLeVtB97ImWSJC
3t4k4RfFOWcNj+fbKsCzHBPO99V0GKDM6CfVdemVw6CFUKmDgHWVInaDVitz8g5Z
OZOqgifEFLmDUpRG0Y39A+IqI7kJe5fiOu+ko5L5/l3a51BqAxGiy2zNeQyfGyoF
50n3cMgiosqjV6IxowGuVoWDvEsUIIqQsA/QKd7rSTIsGRRu7Yk6pOieceDph6Fp
+oKxjnUL74lsVUA+mXqHw3XgqptzlOeSOu3JwX1Y5rn9QSuFlxiwkhPwGw8oRyJe
HgleJc7etsX483bgbGe+AIdkaMDWlcGsfO+aDfkCZd0XMULyEarB/Z2PPHFpFAf2
7SGMCcShKWhjlHfTbUib92neiN3fw1y+7dsOe5ibV1NuX0rj23lWVP04lmFtYl8L
3aM0jgbm+OPnpfzEpznzlsp0lM+BFrE/bmLwkUmla5VzYzqiAGOSVmpTDhr4fTV0
Khe3nM04wiXd4lxvQGHihCVEFp9CCoR0ZmyNc/rRtIxf1th9hc2VhzaRXz4xc4a1
bGrZfrJp1o17RCNNlqT2DwRHvyknZ4h5KgRQajuRCmeOeSE6NcB5Nmo1O2CVzCuj
WFKRMzUuuMb7gLX5TdVlTK99lxnIj6Z8ya2wIxxcLl8rWPoshQTmhocHIfnL7WUM
yWMzqWzt8NxqeTi2FEkYltwSMmOv7HGgDuuu/vjXSKRtGo69dvQk+2nxLBEmdKCu
0qvk8g3KqtHREPqr4C1s9htyj59XroSTfrJtsqfrVVxOuvtaMwdbOmQtHpQWbdzM
Q3Vla9VbnffpW5cB8qyB4EkgdXxXBhJw4hsFBt0bHELjNyFRpiON0nu/MDi1NlrZ
LD/BjUcxFhLpGHX1kFDBAMr5Qd99eu7HyxK1XZzX2DBWuYZ9UqzK66TCr3hGB+iG
GBPwgPQ9SfMRoiM4Syy7h3Ig12y4SgZgUeCAZnLbiKle3zZhlMphL+ajMM8l8s1W
2QXqERNsEjPTzVtGhORDi3Dyl5UMw0dos+PggTRC7/unItVV7jZUqmaiX1cfjUjH
xduqsevTUo23eU+gCpLawyGnFnpCWeIcg+WEkmLeNqvjr22iXA9hyYmIuimtrpon
fq3QuIzg2rdIsEcpPpIdYz5PckOg219WuWUajCoEfMkfWUyHlCTO4PpHDeu6n9te
jp6Um311+/+5gF13NpnyiEiZ93WXPy9KoaucbJjhoA7Hw4Si5JvliW9o4KLWPbN3
cgFaz8egcOfPhafOXmFgEAYhB6k0sNUVVkFEcZVGW65LTVBMUjImbl2cs8u0RbXJ
M8/UAqlso89LGIKfPneQcsli3bGUgLNZMZ+NubPCjsjuZbTrRo5T+8z704i06Jjk
mD8DE9PabuRxeveUrzoiNgD4qp/KOpvH+VRQik0D+s3jAk2JCYF0TKj1eADNlDcJ
UxneaTuj4Dq8Nm6PiB08ZOGkmmnGc+fQ+gfGzi7MbgrgQidM5TnaERXtqmC3Ltw3
jZGDWEw9ptXNoI+C9wQg4LSgaG66oEw/HVhM9q5kdjWTkbeIsjL5h9n2lAUmRv0P
NNewemjpHHTAOEsJYlrAp3w0mUyQ5PpaWYq3+Ab0bqR6UOkN0qtdgcffPEY/MtFN
rGuDXXY/i1f6kYM9/88EpsD2PW9jMXuz5V84gyB1bjQZssuVhZDCaeytHbyDEZbQ
G/8hL3p5TxfW6u9mb0rVeiJ9mExJLR7Dpsel5S2iLuE1UKOgpI60lfEJO1PsJChs
TqgSxENh8vChD2ZlJ9YEnHXFMj01eG1anNXdbdn0ArS8AZBsI3XNdJQgbYDOeyJA
Tjj8/B3L6StnufbXJZa82fMEM4ncA6UChJAjlNjN76Wm/JpEPeOG/LSV0JEAhV8Q
E3Nvb9zBILZZTXA/waIoLsqsIL7/JbKrNkBaKrWGoukP68btbnxxd4oYGq7eZkCl
sCZePYaFP8v/yChhAAR4xvvmHQ8SN37dZ9WxCZkBT1QN24LV5nW+jzEoVa7KZuQM
utdHEKuoJFoXPjc+KNvZ6qd+Zapr+1cRFIXm5ofNsrwYYJ10zGN48enb0BiuqeJR
fjsZKziJk/zFXzl5hyzVEV9x2EQ8ii5Xy++vh5MjYs47hOEwCbWimYJLAJEt7knl
EMfamE/uSSWGEujfWrhQ08k6u7oYyNXr2sr+bQND5/uUG7XkUlvEy/QOj0geSn2E
aFz9jAXIF7KtPDAbRXcrQg6dCy0P98ZVgmeNYkOpKX+NQxVlT9h31cmdmsxVO7RE
7UNdgRJpGjO6O7iRfVmdlrgk0t3ezYJPI/8FriW4UUkfLuaady9zZeAlUAme92Hi
SJ28CJa6MWXyz09HWQVo3T8v0JSpLR6n63bEcdWdBVHc8wsCuYToj2Yyx0D7A+xa
kYxu27na2IIMOmkK5tBV35e5KduVRin0t7cERc3NlhtYtLh745uLx4s8+uo/wDbk
b5GFSsUBnEHDzVgHJJCd8Dp4gcHk5ZKbYo1xm1JjAqUO3FfSP827uWhZrCgSLTBC
4/YTfprpp2ikTo0Qkv0Hn7xVf+dNEhCt/d301wOMmvpH/W+KP13f+H/ku7YPImSN
J5Q810uL8+S1ZXBInefLWlFexK9TnyIGapZDSfGj1zHfghh/0VZI9PZ1BlZGp0ho
jPKCgB9imCFSrAmJPK7SaAxYG4PXGQjXYmmK2P0mC4NLwAU74EOLGzqS3fx5GfiT
vT/aiTAibm/BxZxesPneUP+Y1iyowjqsuLduDmFtaDF8vTyU+zCmFmki6DPT0VMH
WRNBwt8mp8GbLBl+wH741MZg0LVyCPycFAlWLCT08kUIN99SlPTyogODh5M5tWX1
dSz1nIGL/RlcUKhEYkc/mlGvtRS4N0OpuHY6cIdpiaRZUUP3FonbOeSIhnQLEkWC
FmOB4WpM/U7C92WrHExVGV1CcjR+TajZw5tlTNzNBDvwiicTb8RPer9Cl2Dtb3bB
JXV1Rk0cuOfIcpjtMMAzpnMmB1OpXBdvtJGRpXP6iJDzoKLn7hZwDc3ZjqeTLTRu
Ta1SkD+IKnTBEd7gr3VdJF7zpJ63BP0lobLUUALlqARoBbt2bAu9kixLDS5/MXSB
JU33dqu499TTmylpkCaKcJGo59W1jA6sZp+RONbj3fQwM6ou9XClUJq+NX/HdeVo
03t+HKE0HxidQFEmWoRa2znDspRdi68A7xeaKREP6jsQ69ML/BcwwUSkWYWSzyXM
tExowpmGJhOBzmenKlnVOTCuFV0Ad+dcMba+OK9YKJ+0CdYz8hEaRSST9kgWDDxQ
8KhTfZbIb/t5F09sst78/GONzBLveBMks/99g8jS585/MA+EXBHNNmYsWnwXGfvX
OZZSn9ayhiX7WxL/8QvyStsaC0Mr0FB/I98vyE4EH2CioEoqwqKGuHW7szShzDUh
lfR19V949OJkFDBqNcSlXZHRDHOLt9qkyxGPgW7ocEiz2tycxCLWeO7HMS9DSpZI
sD5oeCwqDiZ2Q75Ax9dH60fkHAFa2wWCnyPCuNwAOZuYOlTLNFJw5YJk5tOKHnJS
lO1JvgKVQjAwER6OnD7nvlUepNuc4Oah46p/TyzUUqvX8oSB9D2SZFf9FpekNS0n
Qg87ktfWQyaVH5NZP3IxnHxoIV9STBmYvz51moGio1udFVB0HnScAzFvLkbvWTon
BAehKNCyD1mk+qT8N4NfWJFgophDoPMI5ShNg7qGbz1CFegmkbob6y0X8FruzuCZ
RgMlQxLziy/8TggVN3jujxHOuqFmJWtSSi+IgicBHCnpZ3d/nKXhlqawT6KrNVeH
EPja5BnYyYOaTMdotrnrNww0fvjxCDCS7zC0qT3w0Rxk5AhzwLPJ+qCoQIDTHXUj
QIFrgypN5Fqu9H12hEDo9tbxEzNduD9zietD1OHdZ07kQnQAtRgV8Q2w5koIj6uy
m88nf+jFYsiEP5GtcLhuKL/gs7Fv65SJW2rHGCpPshdid4C5bMgoPNCxbl9zn94I
TwLpRwig/yNja+zsO7qBKbpc8SORDK11XzuEMOGY5wIHnEGPru2ERpkyAoynYcot
0BwGQEoJ8Wnzv22jz6mIWPGWveG1aLLSeNLoRqbp2D/y7iJc7WUOSVVVAmxFbSGJ
drikWxtmmMAa9XUh6H85ehzCWiYzGe5RollNcDL06/eDCePxWuaBBme3b2nJc2K3
qqKS8FUHScPCnwnjxHs08+rzQMGlfFcm/hHUIaBBJdtByyN1q5jQHSeV/0TAf++g
BkLCXidqSMVSpvgIpm5N0Pbh7RHLgzfPy9LDnhOBD/jiFnlOuLp1gvTdU9iWMo5r
wRPicRyKoPkzqXdoEFOCR3Ez3v8hAtZ4S2rLNA4e0TqhMy0rp+oMJVY6tnLB/DJJ
MSJty8h5dAGYZAribqjKZEHoNlF1AP9E1rHNnQzXSBHwJp8AaOWVt6BdK3f0NCMY
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OeI2ebRAIpHLxMYD8NByQNmEU+dzfKpwTrFss/0VtUXHvX2jT9AnAksv1kxFBeNP
vLhP10iIISceqxoj9RCFdQyFB3Iy9ifnLKPrxwyfNpRHbG7NEsc1Mrx71aW1mz29
7q7j3lH+85Zyh63fFRySUfyYAGu03VCja4Xaoqtdccw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 394925    )
D3F0FrCxDmpm9+m8br1cV+dtWqn6YWGwwrBCLS+nFGknhffH+LQeCWINCgXxNhzF
l40t/SIJU5PQupMLQZpD9IPlRWxhoQpg6f25WD6qHnhg5TtYgVkF5kRf6bU92Ref
7zi2LlTtZjaUqbMzp0f+pKhpfsjdzIMRMZh6j3Q77UU5F4WtgBemfsDqervSEzu7
mSqsKdMzq6Tj24s4MJ3gBuWH19xwH7oPOw2sBGV5SiNUz7sBizgeutLmvfkJvHc4
weR60YLqnKHx7wdFO5mjOa7spDpbkhAd7ho6BUvPHfiDRypXOIe+/POstMKnvCFa
ht5i/3gXBCtJ1VFN/oFXu76uaoIoONEICO26QvskjI9PdcTcTuc4E/QiOYAFwBPx
`pragma protect end_protected
             //vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
hX9+KlJJO+G0Uc9h9u/slLEHnzXBs7yQIeZCJ0hUfS46SoZVLySVZIppZpyk82f5
MzqJS7r/InrZBbuRmzRNZVzuXVSXcJUsbKpC6MrkQCIGiO81k4Vk+DXELJcJboJ7
VD1INzsmhygSXajuq/5EN4eSuLc1jdkcy2OfGNwmrC4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 408306    )
AjMsT4XhEjsM/Sk0z5ysXaNlAZYA6AYsbaB05PYjtbNLiYd2a/H23DjOWqOL4oWp
q+BZuphnGwuvjgDvd44M5V9d3ISTQ/Ifv+ig8PitW60kOW9XsULTNAZx3lENDssq
jZiucgrJt9GiSsLCGwvUvuMlG9qE3N+B62cRd3fitIMnsF4Nl5TOUzViTdkV6LG3
jV7I+KCYpN3kU3ytnBKSllcVPalnkSdNkUqgx9Ciju7cWXca1hW+pRxglaUkPCPv
ILZcnmq2aqABwVjSSN3qTa5I82tjElZTfsuj/TqkC/XwFz8Ziw8TSEqYCWkMjHju
Y2rO9jb2lqHZYpwEEhO6rQEe/cTpqA1P1Rt7J3w8YbMztoJwoIA6tR/LKJQaypwd
0fqRFN4jyjGl0HeYOHWnSXY10GqtBxO5ArQJ4POCYX6G2j129kAbSzUjZ9yXYWNW
/K9We2S1w/gcfbkQxxB9khFa2NvHYSMpGnpm+9Zy3QpzO7NH3mD2xh1ntzXXkMsA
G0gMkF9lb/yViD0SOCjlmbWMtdwb5JYL4aaazzXgxA+eStmuYE/7s1n5QqokLYy0
SiU4OPBbX3emr4CpffZlUAnYg7Yn3WO7pauM+UBKUNRM85heKI7/EYkxrEIimbE7
h3Cl2c2Ghi7Km0sL3X2OVcYHU+TCyNqdTCpIGtW8ppVao5f717WiLsrnMs1SpjPr
ifsJ/BhDhcj3TNOB6C7ezXxgJI1bMlymbfwXV4CdwM4DsqTqbzrMlCAIm9Zu13V4
PdTTNkTQptw/OQ6UH2VV7bobvTUP/LNE1//y28RGy0POpVxPQHNSuzt8a7mwnWtr
PagFB7GZnKIjRRbtFPBCyH00x5vxS4y8gEoRrAdVxBqICANyEpnbsVeHxUFSyOmC
1Y16Ct7oXKlwe9IitudJgAIXSFdfrSQlTjFZ3hFrzSV/+203eWv5Z53rSYzl7K9Y
PlSlJk24/AbCG1BqHa7q9XwvmAT0Wamg2QSGuKN3CWc60gwJT7EACgkf6MoJ4jQW
v7Db9rMvfudrgHU16NC3QILdmDkMQTlnn9wWoqwm9LcvotkFt/6hAztS7d5vdalU
ZbFyVePEFT1rVu7+QITjI4zNdncU0NjAl6Xtctm5p0P13/P1rTATAVqB3cUxbxuM
X+IqL1Rve95fbl0J8Glni1rhSU3UWlA/O19ROUHPw1tj6Ygw6Bduid5DqASQSL8u
xBChbk3kZhlwJkeQlhQ6n+qXeUzyYsiWJycbQtiR4N3IGbYTQeAcZKITo63HsTY5
28JANDx+A9eBin5g2rsvWa4Lf1kxJckKroGjFQdEmUSs4WT0Gzf6c6BIyMMOCBBr
zEM/UUnrCdxY25NwFtNKMu/g6wfF5tqfraSjHMUx8YCnC6GmSGX6OJ4yQ09VJ6x5
veKIl3FtQFfQZR+Fzmetpdii6r7KPF8e4SmojkasIfYL7coKCKmaPgWvNqa0ecpc
2yFlyaofMGkKK93+cvm34B3zlcef2yZ6/ukvHOlH7stoiLF/Q/554Yb5aM2ZqIOG
Hz6T7kq1KvaCYULshs9sKD2j5Gnr79bZBN9YjEzVPPiUPK2Ljo9jIBNFVbdbCJ6p
S36IqcSuX0dEEWI+bPOQqkX6ild3s1ozy4cqdsf9gawlSg9GQdFSTQPB7xlXWI44
9oCRkpBiLclU/xx3sreeAGNvVPKTJli87LdytbdGRCIKMJzb5bPhvANWGxrYr3Lj
5zgfz8zYJp6L28sMPFqo3uu3XlB3D2l8G/aSqpVEYcukYTlnThX/dw603x2QXQM8
2wiVkaRoOFUcIgnu+o0/t/0i1cwmGZyavvcUEzLw+9goscEiHlywCsDD4u6dTM+T
9LVVYNFG3I2vr3Lc3RrvcGwqWDZuHULostAhc+1WcYP0cyzoELvWZILpHpHl4aAD
ZZ0MycMeLZXC8tyvt5iNyfZyhOb9TR91/jOgAuda2eLRn4lbAjOEyq0/gV7k4V5h
bg6LrV3RdnyjAIOWhxPK7IbNgMp+iO1uO85cJmqCjxW8qCTQw/bWFhWmjoo5Awt0
UgGL/8kTuwqEWMHvj07n7qleAd6yI0ehlMpG6gYqzNSPKHM+HAdG8ZXVOQ9c/mTL
06tNl75Hm4BCj73ZgQq2ke6tXxCq8Y2SsieBGW96JA+6V9RJ+Ni0YwtphMtixvuU
su3Nk67QGUVA+48bJuQOkrnNRXSh8dO3v9BhFYJIMqHlDvR5y9wVBBPe54PlSElK
Qpr04xcZlr+dCXa78JgHQvvu0ItjvXC7wdpqr6JFt6Z0HzpgppYwWSJT6mgqBkbC
IRpeSGNjwkcZSRdxiKQ6I+7DbV4GqVfjKsLHdGXhAkZiVh1wx8GBB3w1rfpll5Kl
h9329LcqQajq+ejBIWXBJL3TqojzUDL4bGxrMn5MNILPE426bLk/zUuuYt7Nt+np
LtXcTMTd2HQ+2zqiXU5pxcgGgbFySiMCOt/rzZLFscJq1NxdUJ3ECuZgUc+L9Ujx
J3roaw/zH5dh9YWnfllSkR2CRXNCSMPSlxJDUMREO01+jTflP83C23mkFyG0D7o2
m5DOg1NdGgcXwp3Vb6mdl/nfsHpBYrepKEkGrbwdBbtvCWOhVML7eiqEPqZzhw4q
aq0cVKDUvf+lu6pi/CPVl8S93t98fYPupJOazQySNM3k/GbFE7sonUx2Ry/dw6RY
Z4x1+5YFR5EPKODzfw3YXkcuVcncD9XY9xuJsFokWAyecQshzRcwcSMqtq41gcFw
5pgyA89ZGhLQDwhL9Ao5JS/TH+9gBpXd0b/meP438z2aK3GlyWwQaRA2QFnnZEIF
LZo02AVhoAkHJlJUs5BkQv2RWlmplZ3IOJCAQgYUfbwiebiveohQphDf78MLluyC
dos432teCrDJZ1qu7Z4HOtoiAIMlXpsDGSlwwif5gwQ7+RGO9/MH4iHfOfZw4GM7
p32u/20HhgwAYwAgjl3GLRjLUnIr60EdzeZOH82y4xDiARN0BREO4qRVCEP5klbC
4J8WMJjArLX62z6EuNHqiEQ6e3PufZ3HTYBihzEKt6lKDej4zJlAW7EbhEQvGV8k
R8buQimifywWLu8//iByq/43MX55HMvveUnlHZQfQh1ShXvr7R33vhonW84g8BX7
ReatflsAW8izT5cLzkZc2PZXeEQ1705m66qkFLB9vO1K3rXGP9scKsUatDVgdrAs
spLg3OAk3QoHt5wr5YBb+amnN7geGulXKoZZTBGwq4uFxcr94xAnTXUCk1lKHYvd
ZxPe0R1bbV/+allrFImhMVi4RmX9dBMwzyPc8aemVo4vqWLoi5LbyHqYBPpqZ0ox
Qo8I4YKNoTtP+FyXu1bEHY7faSP0qh4nBFa2GT1PIiNnprjkCT9iT6eeRyHwXyVs
OirSZsBk2/jJQXVgpfZdFidvwjy5zk+7Pzzn8RdqdWxqJcgNSqNTBE2sUZcSesUE
0WiavyQdzRJ21ysk6aP2NyJNXzPZZaMiNBgbHWtD24G3TvX8CH5rImnqax7m/ddt
Wa2rHD+o5QaayuczXvT7WytRWPjmwwHugfQ7Z0LSto8wZT4Ubmgf08r+774H17kU
Ap+sMu1ckOLSGmmsSUOyQuZaZdMztWMHp8PaUmXcYe+8TmmwAILBv/HJ+ipg6OEa
7zpZ8Q+xtrAwnmvqwLc4i0LnZfDBwmspQgHicdkChEPbBY+qPbH7EDRive7VB+UV
oPRWfUu7PoVeeXVFtb/E+rLU5IPtZ4QLubdqi7tYg8/lQSfBiA/B5JkvNgdJnGY2
QAXCtKhlNhfRqYQ2zyiO+1zRZrYepx/VDMqMNmHvOts3ccUUx6dLeYIZJaNVoECt
ifDzPeR3nrkJWZml6p+uxTJTpqjc/P9VBojpvWLuy56nwp8CAovphyIGqcdcMNjw
qBTYvAumHJr3GDlAVyNaPHcyeY09bGhVKrjEKLfJDsxiMoZxgUp5GltZ+T3AAPsI
SbBCGs8RPc4c9WT4ApVRp0WTbuVm/3fYj2fZLLGF8OGvUD5E3iLmewG9c2MmYQDH
JqrTQj0Sf3lE1ObR0hE2zp4dfZrfF7KVMnE+x2EfMfFDXYgZriK3x/RiWRBEdi9V
2n1qS9eScaQHq87pPZ1mqZd16FWiifQcm18f+azHZgTfVXYPty1BA5RyrrVUk3Vt
IieLrdar/FQjVS/ePfCyHyxjXKlJ+KeC2roCk7F0X+gRuX5qWNF6drHO8fJANa2g
6xV7iLwEuPcUfW3bbZ5V8HksBxU6DGOfhH20mJplVLCWbb2NaU/cJlLvik0d4bxV
W/NNl4W9pBXqhaf1K0r0Qhi5VRClkdh7q3veoW3IkCc4fgkWNAvFPu2yxx4FPKL3
fHZRoQ/olWxuaB6ig+rL22ofGejvAJUrlNWnZUZkMXVoyEIdLaVCvUawDznhawOj
2VKxOqQq9WaLpsga3fagPf3KKxMsDYSMEWdQrx8b/MwKcDFwVU09uv6JPo4O7MH9
5srp1PVDxvv93bsFSwlLQ4P6uZBo3W7Mmo37d1RF7+4XiFPv0/9PrMBWaT3xlHig
PxCsjoq0S+d4y2V/qZQsSQn+GOexquqdi9r6bdM5xY7epv0bRZSOqhvY+9bX4tqV
B1OSwyRmwl29NggT2ipIHYzwwyok9dQ/weV3gVNjAqFRWS0hDDlmMiO5KXZHSj+F
l8qQ6cyq9xGqmpy5FeZF/tKFr99a51e6sJrRuagTXyw0WUtD4jCQ2stoKgJPDkOn
y3v+eTjk0u+Zq+NcjSbdkRso5a2sGAU5LjusVITm/OXDso/RiAGhrEJBioCAabPZ
XqW80sUJ01soibVgYgTfN+SVpW72fXb25MHxg36CqbErFjGfD9otOzRFBaJB7KB/
6WZy5bBXgexUsudW4yZynvoyY0Ehc9b38MgOpPsKAxAvZdrKkhFwS/zds1zJUZXu
oxRhYW9Yi070K6qzpJndr6CW/385Y2ruiCeWYNk3KjFnwPwbDVZSi8kJ1wPn9V2N
Fq0oJ+P+QmzkFAYdHlvCs7gpltBhAn3GIjMyjPVQHMuYYc2qS/mo5NfkXy5bWH9G
hW2EvOfAv3vsGdKMkxEfKDqTWOu+L+yKvWALNA40CGyIQShA4YLe5o9RmbdFUgaF
BBmlUvf+gTZ+efn5LZdw2KJxWeDauwxQCj5gAagzR2c3NkRZelwkXim+me5Xbcuw
GXb21OiCYi0btGhvRLsG0dGzc0IjRTYu9CyWZwB6ZpUmw0ATkvd9qyJvlwOqeOcX
VkdcJNDYTNPO3DMkzb1VY6hLzbbLF1HqLDeUCjkaDG8cBphp1Omi9h9o3HZex9Ai
nUKsS1WjKzxkNcSaxhODke97w4M5fAG4eWivnCt7jNRo6JGcjrrnQ/pIizfVWuAN
KRGLV/iUvtZBYXQiXWzn2lusNA6WgurK0opFpRkqTIKeJC2Zl+fChcExtl3VmMG9
Y3w+D1eS7mZ6X2LPD40zl3AsHZM3KWPFTzWhSR1M8Q5bjahXVhrvpqbOTKpKe6s3
LglyIQUXIYVYvxPq1henPefzI+6fyHrKJR9ltSctktjPlKusydAUwwPkvATod8ll
sU9Zc+GN11L3iiuyZZK4UxJrSbBPmDR/Kw8CEVmm7IHLT7Y1QWqkU1z+tyaMRU6i
IT5veAAmuom38jxGgmFtlsKMbc6SWXl71gxJRXjnB5oE+0Y3dxgEFs0EAAu9UP7K
BOXIG9j0ol+tkSICqmM3mVkXur4SlBAD4XILra3NJj7wVRw2MRH7QE2FdM3v1B+Z
jjEJcBrQtaIr9h/F8SZiZ99o+iPDleKybTEa0nzAS5+iWeX/RKuabKfFglJcfEJk
FDSQmlvbFH4Nmo7vkEjdhOJxoav6Z2p8kiOMzWiCEQ6Wn/xi2zgEo9JIR5Ne4Sme
lIDyM0GjtBzmQ76qtNBgo4Zc8hTjbpqBYkNRCdIYuOQjB+FJfYUWu1Tm/aXUao9g
Lzboy76v7NHRahzAHEKzDSq2KMWBwNn66S2+2EDIWdk5oQxUan6A/wCOn3NqY2i+
R0vTCR7lntITU1TYO/um6m3iKMQq2NT4W3FSVnB5h6CwbT/u+HdDh7hN38UwQfZB
E9kqVH4+hmVU310C81G/FgRj07Xi+1V+cp0CVWOGTuYDIZnAUcId/Yku0w3aDUPG
IOoSUxjrG+XFChDw5y8JiCKM2VkV81HGUsyMKgCkKdv75TMdvS7deetv435CS5Wo
f1h8PXUZtq4iuz20K863A91vqi6/aEhp2guyyOcfXEA4Bv+0G/OILft3MawwIlrA
KnMLuMPzivy4ElHtMHF/fg86aLhjCgM3H2yttEhp7ZkXfpIVsFOOavmKjCCyeLUX
uoyr4RP+/Res4yIQDOBgcBu4Qdt9LCJGXmivOvOhFDWRs8ejhIEgKnUDHpzQ5kQr
IwFqkmkCgeV6XdhhxbPwkzeuVVOjijabQLldN6Q+0lje2wrNsBdN+GePROq6gL9D
IJZ2xQXuD4R6FdSA3utsO6tWnop7Zxt7jKeWAJ9vMlQhLIArEZoAX++qwTNuI5XG
xtXKPZlFFmWXBy4jXj9uDmbXQABLAmpdPsxP6rNk2LFKm9WGNHU7EpMHNYLvtDTR
prjKr7YzEq/uDCNvzRy/w4Vc1Rr2olYNLDsXEvlUpU7UAG/JUnFz0betFAOEDmmB
2p65udnXgT7ysIeCIRM7xWMJSFi4jnFSCR48NOadVLtUWTEyM78eloYlTrlb0UHl
TWYo9DPov/B5gkjfIHrvbDGFn/mmkLuUjstYuW9Mhv5buDhXnJXBcS2sZy73Sj6V
jsMSN3ZuAx3I7NEsnbk85r7sgRXAEVRKJpJKWQwd8Qo9s9gzxl37yW1CGhs74G9h
Yvrv9kOd0QvIPrthrAfQJDQXG+S0QgKJVPTcGCTwWHQ+p4458veD5vVWTTzyxHzp
Fv9gOuRM3ctuY8oE3rmMdxSGXCx33WaO26KZP5LvsYIUTIcPGyswgGTmgNgOyQ8a
mBX5iG4dxDt5Gu0Bfar4e/kzFF6apbVQVMOiMA56v9RR0AvOUuduTBiTv9NjuZc4
U7zKlZoQfUGc19ce0CrBu4UN6o9PEh6nPav9ezKJJi797eEed+Y2G6bRTbYsV4AX
cFxmW2Jij3YIOFD1RPSrx5Wh+821VmqqjKipCGskqNNDuxWTHeeHtHgWndX0xSCX
ciyBG+ohJcqAhywtetALFuPHXVRltYmyPwgDuQVbFwSDvmlt+VleTsJRoqA4eioM
KM+Xwd4mIdKWepGoSgi6GKp1zfUKR1CFnoTUTpyUx0SSolC9ZCUoQRf8kZvuqODt
eUIjkopW4XxbH5m5C3MACACJstdHjGVsyf17k8lyOEYhIVn1A4Ip01CXg5lIuicQ
tpLEY1hxirA+ApY2QSY9xw8GuGMYQmco2PHIkoypl1sfEjgNF8W7mx/P6MAnrNgv
HMpl6QAtSrbKPpqxF8c4+9oXYGFVlUa5Ru2nCr4CgDxHk4Kqwy+THPOdpnnjWL/D
8Twrc3P3U9s1r3cMLcrMIUm0U3HUs+TYXzJi9VlgnDZFpDwjUUL6j6k9sX4uQvHy
E3cwwuXvGvrxBlDAWyle5Kcs46OlVzEPyrOflLZtMNurIidQgGjq8g2ZJYkkxoIi
dSU4Sp/mBZJs1UiuHlpgVLoe/V5+q03NDc+IwcaTEbuu1hH+F3MijoXXtVmh8uyr
R1+CQeT0nXQAWpS4T/Ncg53Xrz7/flp+UUd+ma87/EotmUxHC+Np246LWPlDI7Qd
7vqdBJgRPNzINhgP/JZXh0z6upCTq0eatNt7VtSrx/zmxoU53PQ0nEMMT6b/D6cu
a4JBjGJfkYkA7BH5RNnIYdWs07j7jfUvtEIGaNqlUP0NqZT/yqVZFQWy96Y/1XMw
GLAkgld9Pc2VA+lF2yNf1ftqZAPNb3+NAAYWDHmuhbk3WHCsIAvqDPt2oujdd1/5
pdT5+gHQlAa8Q8ikwgnZ8XA2IhvlR21/scDGb0oVvE+C5lgU7aZWd5UrZg5arnKQ
rwlWkM/UFxKzyNX5PtbaKxNfuQh9EfTmsWF2UFVfLHlrRUW49i/w2N+vC+F6hzNE
e3PfYcBBWEr/B9REBjiWUDASYacI3OgLixOPbuyoa1JWHd/JSrJNS5j6mXJd6soZ
We0f83LP/WJaOdP1jP7drMxYiNLIcmD3fxX6g0WP4LFYVytI7mOBMXa81Idbm/Sm
Dy56GDXxKgZRpeJJW0xyBpPqG9D2Gn5qttzgIEDgkgjV94D0IkdvLnYd5e46AFhf
K91u1rw5PzV4GOvQrNjwwRriZwPMFe1ae5IkhZ5Ixs/3Lr73TPXoWy2APTq/qag0
Esr/XLmQ7Pv2WGbMno7Bom0wt8JyQmHZV5I0P7ctZfaZ8smSHQRU6g6Dbn8UOl9R
FkoHDx4dnQ1yhq/hem5tuWN2uXXiZ1KDGIGl3M+wgHGHCK/knmgQjtaflvjoRma5
tXM4nt2dGamIFgw4dLz7WEW67iMWhPzvam3408RQBL/t4Vw+a/NNg1PPEcjooRQ7
aE8aDHnC763p787wb0vPU0XoxV5Q0dGpFHHghni80XaSjjs+ACb/YhYgGVUFedxZ
M9e7hU7G/tNLlZFdFP9TGkSsWXb6HmP/UTBJkvWBEO7EVpACNKLgiq3mUylstswN
6QmaxGRmNvwxJlynl9UT5F4/RC4Bko2+/ZCAQXBnL0VrgJRRLpsADvPz33Nmrw4B
tZr4UbzWK8D/zIPZ6wVTiwrzFNN8zOr2KprtOYSWByZ8tDNFbRc01ssMBpAO7hqK
n4WRpc7kudEczI6pi/yoOhIV7ZTcJapHDZWffibm2t4RJp5ZrrbgPv92Yt57bBlO
riWcfE1f3gAUE16s52drLFlvGovBbxfVpa+ZkHWVuFBWDAQaXU9Iz1oG5VbFz16Q
1/UlR9KMQpMX8+oPeSnIAatMkud2pCgRaxGKW1CitnHO6CxnyZHus4LunbdiWJty
V5YVKGklyVIumfEkGNIvrEzTrcl2nkRS9wvfhqQB0wtH9Tc7Yk19WR6aPNpz3RCZ
8cF5OX9lLWpp1urahs/YcPnWdlDSn00X5mdrBdg+udU3F+dqFL93lm9svLDOPXnX
wDrAlBYdlkVI05NrXi8/lShessBDZyXlgbryDgdkO4X4gPWUGJe/QSLj/tyzJKVu
9vikyaVglXQEMJ6WCOYqW0EpiBFFeMu1Qhc4QIe4FC1dPfEpbtfCSuZcaEiL6zkf
DoWVVXBY/BoBzHNHizuBo+jAkB4WeNXVb/heKcPvcWBA/k0BT0CbZHten9fCQcX2
feoM6LPGAjdFhEIiF6axIcbhj72Km2ot/0KKluG0fOu6SpMXnI0eA9aPwyEtYqSN
p2m5OV3AuG5VX65V8CQyYpYxfCRaLr9f13PKMMiKbh1nziIhxE3c6lIp657zFtVu
QveooBIWUBh2wsxPuxT/JpoeQJRsmMsXFNKJQZOg8gQ3whV/quMlCjuODx1Xh34o
9U79CxymrpkBJvCfsdp7zB5gvSPQv7c4xNN2W7XLcSeL7KiFDltKgJhv1IPNOQn1
AV754drqzvZbSKZd7HUzc4L6/oNejIbuJKZMNG4KpflIqpC42eZGytHDzksnTHPw
g13MUoI7EYdg44WnsxFyxGPu65gLbqxvI8hj/marO09G06ubB+FsFX0XkGRqlkt5
6hYCUZTjxXA7XYkDhdnjJRZRd8qE9HuS2lbTdO6WWHY8P6xioiOBmMQlVvdE8lJa
MwviEirahpxDpWdEbJY7sQY55eAJqnXhdxAapbYSRRqnGPAJyIts11mpHsZd+Mae
MhYZQUq8sBC00p4bFCVKCI7my9f1t2Bm7ZtrLT07fl5IL2iPvplwVxgcCbiZ/VQ9
PYIj9DkpbGHZ08J+c8JGdTIdVzBXFNKB9Al5Ok1Jwdtot/0A8BMI5irUqK1ufW1s
tjF3e/WBJDCtf1b5zqGSr5KG1vFqpbe+4/BtBvP/zISsgsE0ctFLJVBRmdu05l4Z
oeo3bCXXcsamA18TvvzugPc3y+FpU1BmRYOAJv4++MB/qh+ywh7DG4DgoLAvU5/T
Lu/zpeeng5FEzDTtQCBve0MdMCiJKJRGZCXoNZklsdIAWuiHMUSxvEv1Jwb89Kpr
wWN5rlWt1LfuhVnX1Dozqt63+4qMWnmvqtZqfHka51RNA0Q+e/7YbsHA5xV4WGjs
g52FlgwNzxhLpASUL9wcrtpRFQ++hYxRv+GKAF8AAuqx3jup1dgtb2nNVQyhAmj8
aACzISF4ktGstz8JGA8gNesSCbc+qGcT5pAU1lyl4TubbvOh4Ud8a8Ei5aSmUZr4
coCFR0k8ZPCfJtZ1hKGIsd5isHsrMeIgJEkMugIXuEVUz/M5ywemslu/CEi3izmh
AUjqTd0Q2tO8SRdvPnOje+JZctQWapcb0E1yxSutGuPXA5QFw9SRcNP8Fbus2OJQ
3qmdEpQM+MgMs22Dotj5bQR+lB5YaOQZqocbBZPPHjVgNDcG6vJ+cmaSE5JttyEC
kDSvNCJ7Oy5GfRO7ohtR6UWcnRBLZywaQ43EFlzAkM76KhvaYgacOFp9QThyLlcG
vAd9r/7P6LhuIHXGF0QWOUZvDIhIHrfHT0H8ky0/OclT7oCG8QxH0xw/jiCejReS
hFC0FHBgVD65xuttlbYuH0NFrZm91pjDGeZOSugsEfiTlAIm30FL/x0LBXJD0EAf
aBkTMID6gHFTny+PEzJ4Sw4+PTqV0U8abenp9Nxyd3oQr8zxEP8tvRps/DziIdLK
zNEl9yf7wvCBjsbOkd/e9WCwjmoDYh6cmqpCQlfORFC7TnqFWSFLn3osQ3mLRPbm
LG+9DcmXh1YWfpVtr8sBXctHz3ZpKurhXVfwGKPyn97/xT+0Q3dg6BrTT9V0GT4S
z5fMY7Ryqz4fOc845qi0zVp5uaq5abttCoG7atU94osb2bY84PsNYwvgFiHy1W0P
XPHi5FIdPbwPhIpmnVpoNvoMiy1hwTKQ696APQ4vdHwDDKUffzW74yJBpBa06wFy
cUM+UutVdfT+A+XnkKnCN6bMfZom6zbjN5bZae2vVUJb95Ea0dcYlecw85j0Qv92
8ibmEQQkKXkJZEdpLuj3w82opBWVf7hN+T41wUIGEAOvl0GPtwxBf4z2hP7EDdYG
XA4sNwzuc3TB7bz/TXLswcWKpVEoIckqEfpJojwuAIpn1lzv+GkMsZOrCy+xjoT6
tzA8sb38sD+7OKz5XkpYoOXxosYgjTC0aHbVcaBen/YUDRD2/QylMMJFzYYGAcbF
ktbzPtPh07MC7qZVNwSyTdKDIcN7sIJZnC6n1haVI/YI92IlncnbyzWBcahlbZgk
P4nDf+F36FpfRwVGC2Eu3KgTLARFdTxhO62W+fUZxOzLK/U32kjouhrxH6JOYtvI
AKsraGQwFTnx0F9qlmX2tFkDHgtMHRKgQB4lZn9LgQXlHnGHOcXvil+/ovlfhxIM
oUC9S25UzA8E6DfxuB1FK9l4sNpLHRmGoc1dSPI4vVSxvGi8mvFh7OAJ9KnSzGvJ
o0XUGzoaaDoNps82HwJ0SrXmE1Z5jphTZ7+Zyqn81vQ761XSqfjtFQ0+OBtOUKuE
EkN1r1wjkj9jjuJ8VSPXvxLmH7RB4jW9vWOPxe2m3KcrxAWrWMNEhiZ41SVKTT24
ocVZmTcNezuKGK03b8cpLjMAl/ywl0f9PnqAMOlC84d8L99a6IEHMGoATfLPSX/4
zDx5lw+ve53DDH/fXz5C/sYqX808/72P5lMijYr8ypyR30HhBRaw/5010kCle8i0
qfNxVDjehLNNblQ8+W7zY8miXL/Y9eNGCjTXggDA5NnKRK1BtRFWUOmnw4pPNowH
ttkcaNTupupyLmzMJS96bqCu5YbPQVx6bXsKV0nPvtuT/woLUTMpQUi9CBs4bm0S
7a7hYTR9VuOytbIKQkWDyg+u5i79Bv28bMgcaBMykeInFRszVIR9zn7jJ8QuHLlE
ONS4/8e1P6HTbnfK/MqvsHXfZ/yDSBlFjx5v1nM0oq/jrDZck7Lu372Pe8HKWkOu
x77ugDT+8DK1J5u/VfGYcFRBY1D8ppX11b+S2oZ+8SsoeRQ5lUQ3E+iqz2qPWh7v
XRu0ZOKeeGQUbTu1soq6x9ZvKyuBFOF/ZbkBOECp4H3xnto9Y6QiHgA17t9os/nr
aPUR7iic/mUYlWS8Xhwx7qgWvB8fb9DkbwMmKndXpMyh5zN5YSRCk8DE/aLxoo9G
doUkMvH5E4CwQJF+IONfX0cM2CYhLBLVdt9kBzV81HFbgsaMtXQZfloqL9YAV3QC
Xs2Q8En2pKp2js2InYIT5W1+jdo0hBZmvn2vKwWJ50Jk5naSb0+NutzUsyifK3ds
QHjlDwlFkhca3GF8xy/kT/HSNVEGJLk2jMI462r3mMVM9LPejft1iBh1rMA6ER8Z
SxDoURNWLOQTnbyhIpqvNzsbrvgB4ezdyWe05eEDAOTKZYc4uyd/UWzIhSb6d8Gu
W1MXEq49870e54E93Noi6BceH7KziFQfaDzaEa1pLAEyzTjPRbLjbWTTYVB/E8hk
oeHczQkbvANsbhP0StpyPye7rMC7cQTNYNozOTragGGA81ujlJgTKegVkvUrc7d4
aZnyXlLiGmz96+xFut3USS59lmpXEB1rPRpfRLhktNbn2viS97prXERFhScfkk9r
XSpUoNzxQBFTINa6rZd1XAcsah2mkCG83e96hJWH+aMvZjcPBKHK28FuNABDIgrY
QQhJ8P8TckETKRbkcXf1sChYrumeAJj7JszcYD3BJrcAKYHAKTsvt8Pb5yuPULiN
rNSgevIHCmq+pmLkGAXL7K7l5GngES6PH7Z+ATl8pBhhDDZpdyaClTLhG7tUEt3N
Wan04sNtNWOfOU54+7yIFoZdNUTxW6jcanjyi8Jdb44tjdwtWKB81CooAHvQJtDB
r2yq9UjG0dDB+jCv7PEIYpSP+RMmLNWyam3KzWBiwoLNzMI/rz9Aljn0ixe9e7yY
lBgDoJ3d54mL36rkVwe/jgiyypyDOMwli6cyFkf5yYGLXf+ivTw83fkcIENQ9sxD
6qWQyHMb+2HgpaD5Vh2849s1p7BeTq41NnrRt0NzuA45nf7Fq46mFAdTr2uLRAvQ
ifGHTT2qWKufxW5wt8UCl+4csdWWmUkITx56V5YxfmSRf9ucE6jYVPFnHhzqGY+O
RP+ixTxqBBRJZmTlxX9zRNg0lh7DgRJ8LzJvsF6vaFxBQWSZsvUceKojNe/MamgI
yV6PTzZqMor1pQ4h5gdNUFmZ1LDK/s28wQptt9c0vxH5Huqh443aK4JcXLMVhQ0g
pvEIJZzDZCtvPv/BdqOGzxLZB425UY2rTdTRkF2jtefp2Qx5JiDyAu2nlqf6aW0G
cG1tAV/1DiC3q4mbStvz5xFlbzD7YA/hoPALTRPqvwFrt8Vf8olE+x+QLOhGj35F
Ffk/DMd7G656hJ9XTpBy65QssS9u3iAVgq4WnVcps/UC/lg40cV9SwNXLmTjsfo/
og5byI47zGG/+Vijn/MZU3jew2WPhuD4vP+z94mv89xO1RWERX11TFGH3tTgw6iI
BGSZOzKvy2A6SviYGhlj2ikB//gjoFAmbyVLf18WdeyoSF8UA7peWuHDmQTvhpXE
jg0DOlg5ZI57PckStOKCfxX2qZCgOllIs7PIEyJaAkN+rfYM1N0tAKB5b93wTVQn
THYAKrgtiSEsTTMngq/oB6SK+iWMK5CXODw4TYUUOvzh1QrYFU1X3lELcFjJOG3J
YtqCZfR7efhsT5SndVTj3bPcROAKVMfFK1vqZ401yxqmVOlJnchPCmc0o2hoPPXg
EWbs5WllpHXmTk2kZ26EY11Cn/M1Okm5z5QiaLflqNZwoJfPn8O0oTUkacAPqgRL
O/nwMmwI+X3iOzp7Em1IKQyW3VbguzpbTA4Mb89D6zFIrKhDfWN/IeFeladE6qKW
bqnhkE6KSxnW8fMgN+WVssqwlGmvshBXIDLC+ZUdkF27O3xLgtYvg0IvyvMb9EhC
zE3lKK8/QAIFvD6PelK+j+YMMMXNt3f4NdoFWgF6LqOf+ob+49ob0YnZOZNBM1JE
6f63nY3NMG6G5eQZUmIJk93H51ypKoHpxeVI72ppUY9kwdwoXwOiIe3zm6j3XtHu
UpciL/ob4xT81m9F5vpsjtvDOSCGDWaTH02Z09B5NRFCx3DBIIFBtsb8ABJ8zhDD
9GsBTtE83erfm70s0MBFNdQDdaA6Wkd7Zdx+inaBwaUzmaXoCQ/Zr3tus9NrpH2F
mP6d1jF5wlGUDyzHAPcU8sF0azpETQSrhnMhl1i/WKSgO3VdfNdFgjokpc+iQdaF
6PUEbdapYAoXIj8GTC6XLppCAbvIiopUaJ377TlZIlGeF+8Mh4ezYj4Gp12SOVlD
jMt18VW27ebA7EhYxdcQOTFxGz+QUm99oNV1tD3vFAmcyAqyb8lD7Do5mMCvb7uI
LXtDgKBHPjl5PRMIUp6RSJSVPI8ZJhzj7Tox2IDlj3c7L0BfBxP2Qa/LlVUJOyN6
vbmZgSVl6szuY9oj/I24OVEDJOjteX3PbE24MsNO7hnn2qT/W+UiYaYhbis14QYZ
WUBaqYP02mf3HKZ9SMnulexrcjktyKx8DYP6/hpKfqyf6rbl3j9Mv6ayNyQDW41O
1C3Zabo2p/KHsxOZRf9BGY4qRhQgF1uuNx0aBKM72IetxCVonbPdtvv8ScBmjggQ
N10zp1eMbWGVrLWEE096gKHTQfKC4wlyeih2xiZaFexNs/XOu/8sVVf4FTE2Tjk+
Rp1dLMEo1f47Ai2lk/G/36Dy7n9oIFW/ken4UvJumk19Ax2BhaHyoMcvjpepeFX6
6NZ6gD3ETI9EX151VNsnTPjazofnsyqoOXA0Hcs2qGFB6zQa9BRXPLRhoSmdR0uM
P0bF/6bZgQH+tVVgiaYFUXe9+RgDCpIiSA4uTpUxhSk4HnQ/4BimSpaitM7z0s7V
kAKKQscheSakAxLO/zBcn2watU/zcM6QrCHaDDR0qdK9sDOT/Uv9k4Pyy8VVbbx/
MJOoYzlPR/Fhep+8+cWhyz99RZ8K3K0/lPiysJNeHBaQliwe9IHnCgQmYloWpM4L
x2wEwS8WJPCeP6ngj07yt5K3NdRJTDMtEsKhTQhsVJxUEOQpYx8jh3a6POsKxV5Y
iotIGOfhJCWyFgmpmI3UZTLODeEuCd3T9f0AtS5rZ96LOxbQPP+qZ+fQ8ixgJJxS
kDcUqR/UNq9UmMcsPSiHzC8hlojZomhe3jt/VmL/KZMdQUuY5yQZ1AyqHOldF8Lg
ACfgdYqrKe9vCZJ57Bp10h/WB1sR0poEk6/bkb9mLHkkGMuSFtaVS1K6JG9TDo5u
mSFfDqvZ5cPlWFmjyTyeOPk47583x7tFDp/shrSCuv6LgXRxL1OPVn9IsQO0ndqh
95t5GBEYQegNYUbqdGWPs9naS3HvY2FayAWtvAJUvpJU44paVF8qytoc9KZtCR5O
unPd7TYqepcBmxo9jA8IELLJPHqyGa9zf6zlu7qAngeftg5DPrSnmHaxd7EeZVFB
ljS5hIo+riRYKxMUU4rx1C88M1130vwwfXcCPhv9wxYmgpSIWdk9hubvOZX9XCgV
YeRjHAlqLNidHXLNqd6cn+JUBuEtz/C4KvFH6iHqxQmckB7d/7DfAGTMnh4NduNS
lzurDOoi5tzC2Tow0lsdPM8tmRN3yKBTawOfFztJoiI2oesNcuRTOkDKppM0gVyp
VgZXG11etX8ONOpmlfNs1ivtSD1wuGKLBb0+/eDFbNIyQ34g7Yo7L9cS+KYcm2Yo
O5mvzlV0aYOsANvGpI9Yuez0C3t5moEXVhmW0dWrUzOuyasTLHD0xjxItutqTGlB
yJojVPlOKsOaUM5YaVojq7B7jvuESeETagaDNNzoz0eVOgJwkplZaxVjB6AC/ovS
cfb9b4IWWUwRFH4sEElSoS6RGVjia2TapTADdqoPVKwbtaWD3R/y8jZ9uH6nIagr
v50fdgBO8kMoXWhgX3IZrt3B+yW7fxg9d4rBzMLlxc7DQwQJo0Pxoz6hkJXJ+I3r
WBV/fcYOC44PZD8o5Uu59bDy4iticDgmK5meSf+2edmP+wuAl+0mtQY7dXh3eeui
3PB99I00gbPzc5lNSIFKtAe6zjaMFQkmRh0DYWNwp5Mz1JlrpxsL948l7PcvKstq
Kty+LcroIXwuWfXAliP/udKga3ldArQ1V6xlmn4/C97JqUFVdPguSeFvAovenOVS
TR/R9Yi5MDwqYdv/FGaPgNK87EjaZN4RouW6x9F0Pc4EtIvmX65nDRP/epF8VUzL
9WM8qbzTY6+mqD+2Y6PNbV9hRDRxoBKe/rogo9g5oke0QG6O13t5qDFeotI05v1S
WXA1QXeH6mwn2ME7NOwVVBLk6IvGmoo9jlVtQh1crXbk3K904x4aTg4aBHa/DCFY
j5Sr+PsbZXSgMhI9+Jv7KMkX7FHaqGsH2NbaS9gOgjTwN8lZcobqWulX5QRJDNYm
AnruEMbAPuQ/aHyKSdqW8WraWe/pyA4kBddkALqE+/joxunzB2xdjnnsuLV42Ei2
oioLQBZHY2GhC/2ZlALKlN9Z0YkxP3k1bMZ1N9Sf3ryXmayZZplaXhegfn0D2eql
MDHqhq20foa06xNPMpXk868hyiA8n8GU9yEhPl5AMtgJTOu2fdiLZ3y02EuG4xAR
n361Y9uWXRHBnRLAGdclvgREjRG6MBg9j+uwZRNfd3DeMUkk4mi6oZd88LDvSm5R
wDY6D59S+DxbXGpElSVyadFmRyUYV8ZqpZUrdrtj5GdRK8Bd1ZHoYQ4SiD9kTtnE
VoygXaVwYrxd8oJdOKeT20Z5zFH1DLOTk3myp7eVE3n4OsE6kU79h5Bh9KH+nTPQ
sdvSHZ9Uz8n3VTGj+PYXyDNl1arf8M/sHq1SEQlIH1hd3tVMnXnaFRWXQWWGJjpV
dPNhxT5JPBmCUINkZruT9+tyceeTLV0f11uHy1aBYTIvzEMwGXUfNHCKdfA5W5GO
WWmtsoA8kLmZz9NXDVbdXQNnJWHN0MCQJ2dIGh3RYIvExISH39UgGjFNzBB2l63Y
sdEOE6OkTB12k5/6IreQUYYk6lKOm9R7YptPiYbyI8EwAN9E2y2IOq08lwbwXUwK
rRzQ/v5mBto99mvvoxhNFqBdMQXb6aF8zpLveBIwpFtWdw1EAy7Z9FiudZt77GLr
uLwIA10myyTBgY3MHvRZVdIGyrNa3HwVwiCRuAM58IbPiD5L1V35S4RKNxNdHEst
6W/n4l/wdj7klQIB6AXagvWPChcHdtz3x3nJQPr5f0+OXTN+iy1dmqsUE+63UleQ
dCIn8KEdBw5bR1C0Xx33mrXRS+6sn+9Zbpujt6HB8flbP85lImu2nAULu+y79b41
hY1Dp2J3tqIi7fQzwQZoInR3KFkilTiGfZ/UiAA+sBdDmEqR43uTaJI/J1YNShgl
vCrjU6ebGoasTO9wzBHLDjiqb/9nECuf6ZACxLcOe0iBJK4kSqPAyBKvR5bTvMm+
i5L38SrHZ/oi8c66TUNCu0mOF8VnxiYFrvOlJzk7iiz+g6QAvEuYMNeq4YhPzpVD
zH7PcFk8MKy5js1sVqBLyuVBm69Z5/Jdwx91P4R01xhQ5CkaQ02GFUlNS5km6Wki
6HR41ot3jGbnHy4mntIveQHtm15W3lP1dG0GKhV/hpqab+TDXKIgydKL3lyq8wHU
Zrrd9LNWgPwi08klSLXQ5ZaWrjEG8Ux/5s/FTXuZxJs5vw0X8eOZfNaRo4hQmZ+u
pW0kB7Bax2SQlw/jiMpotCfK6uAodKIWYGZWh2KXt0jJ8hzCO0BXVv7iBdkcJlxu
`pragma protect end_protected

`endif
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
DJSW3zEWMBzGu2lpcFvpTHRYUwTHw7LPyAM9s+4rKsHeU115MKAu6WdFHHIRzTdo
zQzqBENgbOiDUNdVqriNHXeZhPDj4sL5+g13L9CCs85PXx9Zbg5V3b1Sm9v7MjHe
cJI5UBZBgJdpAcbhQ/+1ll/DaPv8kswcvHnydkDpirA=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 408389    )
L4n3Jl0jI6w40oM1r50QJwcKfucLsRmTkOc9Ba9c5UPVRLDEXdk21lGbxN5dMEAj
KaYsOq0DCZzONswluhinCpVgIKFa4TjIsm1O1h1d50EFCjKLTd4K0sktmsXnHDX6
`pragma protect end_protected
