`ifndef GUARD_SVT_AXI_SLAVE_MONITOR_CMD_OVM_SV
`define GUARD_SVT_AXI_SLAVE_MONITOR_CMD_OVM_SV

/** @cond PRIVATE */
typedef class svt_axi_port_monitor_cmd_assistant;

`protected
UVSUO6R3bCR98T6d3#ZN3291(E17@\8QI@O:K[1SQBC;fT1QR7ba3)J1]dAcFJJ4
eHCA2_C&M(9^8WX8bJ)fKWMAM8-F8XOH)-M<C/@TQH<c47BYX209YL+P?1CD9d)#
Of<.J=JfO)IAM,gMMS8@eXIcEF9B^65.)<IK5IY1YO;,-Z_gQ>6d]T6]/60OSSUG
:[?1EdU7OgFTWHM)?2a/3dD_K92&?9=?#f#M/Ta5+I^=dFeJgN=3/IJD^Yf_=Q#;
UVgV?V^4)]\&DYd(^K0fdH@CN@P\7,G9fH2R?Rf&2/;I^&8@3KT([+RL&/aT;@V&
dB8/SU6+KMQ,T05&/57YWNbW6?93SbXJN-^T?U\eIY=A7ZJC^e86_2V;+WM;gJ,7
L=9U\H9748eZB\>Ae?GRAb96:LDNKPaQ]Rc3E4_)&6:).TeZT8V4GGOQg?cZOC@)
RWMH-QBUUMZ#Cd/]-KCHU-bOGLSO90SH<:O5JcFA)ebP)SSP0([HR#-5WM>YWP\;
#Ka5T:1(_c\XW5T2-=@)a[,d-QQH4F5M67\3JTD@#[e]DA36>fb4aQN>@EUZN60Z
OOQ&DQ;)HHO[Y\L2QCbF.&;\<__K?,XZQD2GB]S22;fK,&X@J#H4_b[?b<aB+JVZ
-)geJA^:bK?N]5W1+a73[[-\EH?PP<a1SI]B)9N=1GdL?4Re8N;D4J^WfQ54^Y4Q
YK>>4Z&P&O8B4=>#@0Z>VO(E]P+P]Kc,MWH;G9&0M(9AU;4D.]b8--f5:8CL0>6O
07Z[@<JFD##OA[LN^a/K@D,dZAZ::?aI4W>;/Zg,Q7OAa#I>NE(^#HDRaC8X[YA(
L<,6QAN#UKRcYS>EgA\#>O#IdGGYM8H^fIRaJ@S)]O/955SVCHfZ0/-.,_3OM@_a
a.46T&CF&W&d-b)LcC<<O:d_@\SD2G6E9,Z&-c?U#PM>C+<XN>aP:EK=a)&Pd5(c
M72B\4eD[ddC)MUUS&?+@4@-;JFEDM.JK2eN#U3@]?/g4Y>/?G5=E<TPAfC&1;M(
7MS^,7VV.6)[><46<T<CPf-/cKE-+=,:E)/GK7S.[EL48BI+;)bDBT38R?c\AE3B
dY(bg>6PX4V,WDT];JFN-PgDP:Z?Xf#_T\2b2fBPe<J[Z=L+ZENWeB95&-5F-NO>
#C/UIU=OTaL6-+=P,/Z=).3QA]=EVb(f5K8-&M#=AbL\QUfQ[Q&F01aWDD+/X7[0
&WgCAB[TGK]0fI7JOdV:8UUFM)XTag4QCCDJ63A<..JT)6Y&cKb5Y@<0MBV9)[<(
1Q>>_8O;S4&@&JG,:PH]f2L;c.D(;IKM?K68)9;-XfRcQc211WRJdN>@M.O<:Z;=
5Hd/2)f^@ZJ1N>D48a20(b]&DKJa,0-TeU@NJ_PKHT:E:2_6A@/Aa;-2g?e=OMM4
bV?C_B[TT3[K)&N(G&I/bBSA7Yc0BLI7OZ(NN6H2OMBb1;VM?W6.]XDP>b03GPd/
6^&9;SMO(=5b?dY5^A<&ZC_/f6C7YT.@IV<f&?MI2M?MfHO84<eFMOHO>@=)Z91.
:+IL0?c\H<R?&K?-6ML0N6eQ^?HeaaDXH(T7)>2Kf1M:bD=9(;Y92MbYDG85D).4
4F<CEUaG56^2DdBd-\J95TIe)7?VY\Z&)IN+L,A)O4,46U<A,0&6c?9D8-8RJF-d
SL5\U,Q2E7]2c#7Hcf>gc\P7BI7/bN.@aBXJeP)J(5eOC4Ve-W-@Z,],Z;S-dYRE
egIe25=H&T)fd821]0_CIV5NF6](bL[Zb5)^S[\^7W_d>9&M)4]EF.O(Q(E_MJ4G
CRePCNEf^ZUEU<eY7AB1&4OX9b@14G9,/a-3&>4faHD.BS31&Y>@R8EdDOMOY1T-
Wf=R<]0cdc?0ENGL\XFR5-FL=J,>SZ@f>1.1fb\b6c6=IM:XbIb8E?>=O\PG595,
#S4KZF6;J]HA6NED?@^OGDJcMe(B\)&RJ=-D(9U9&c9dJRf.M.Y+JRQbN9deea;a
O@O2;O]g8Cb2a?a1K517]TJX.;<^3_]KYg4W,^5A;)f,>1.<Q?P?/H:4.5JDFP(]
.bOIC@a[[7>Z:L<V5VHA&NbdN(gb(JEN2,Y)S(dXWA/V@=:&;.E1SX?1GZ5Z_I=?
6^@RD\J=/&8.g?;bMbHEEd@0Dba3F-U)W8]AD_1@M8HQ1KK(<4c:P89)H+:]JCV.
MT@bYa283eE+?@TZAR[eL,4#K<JT]F>:?8)P83bR(cC1A,5NDT?-_7a<>?8_^e&E
BE>,H5AfUE+WI11#<_J1UgT(W&^0-\WQC)+(/,WQW:B^C616+5P=aTG68&c2HS)X
S&M?=GJRZ=;Rg+IQa5(?\MQDPOgGDYP+5S3JQC8Z7J95?=_6QK0?B,MNVFTRU=_J
6;R4&g]N,d1&agO3,gOe762JE34LdX=F9.PdFQB#A^[Y]#TR):8]PY5ND[YbG=OP
4L+5<#?TF>3Q3\LeVV92+I(-2XbQdN&S((A(5/ZR93fQ))5d@K9V@B:E(-FNYCI=
I,.Qc&GFU6ZA)AO[ad;>H?R&+[2AO)IUa\@X0b)cLbV#>8F0^Xd&GNb<7-^+T)?O
@8G)c]53-L)F<AA_LPQLTUVHPb3_AeR_2E?W<=^?&Meb@J)b;MWb^eA&a&_Q6&G9
HUQ>O3AKKJ=b],>aZGFKBf,<TXbLNY;8ZRJJ2U@<d=:3K&5[;8M_YM=#XYYGeWFC
MY/2HZ8)-3U#f=V<G(78TIP4+BE9,6OeO:0/[MUD2d@@;-I)8_K9M1W(;NaTSHc9
Y3T4Se;V]:A-a(KF8.YEKa3,4,L;-ZQKD5Lg_BIL7.dV5:[?1XN?\5<0@d9^P?eS
-C\>0&XSg\CJ?X#LW3>^SKgP_8B;HT_7G^=)?g:PT-b?^bK(L.&5595@]9R-O2QY
6KcV&L)H5C7O>OC@[=W4e554AP0/FOVQC^P7:+85\M_\GHLILHc8XORAADDI+K>H
cbQ19fI><K=>@QFI1PK_H@d#Y2KQRZ:NP3+HK4?f19#<@[9DE-/08^9Xa->TJRBX
H2[.N.2P)Ma#3QJMC0M>UL9FV\aQ3+>=-:[8T0,.JP++[YbHbK0[_S5cDF&Me4eN
C+7]S?SGbK[1VMF/JOSS(5BZOO-,Y_f/6JL&Wb6C<RJO3fUS/VfFW1V&[J<ALULf
A_-#:TgWQ69^<S&e2f1\d/BP]R&49<Q6QMDL)a5:\3dGZE0Reg-L\BM/YR+_a[AI
/W<\IXHg885G\YG)CQbX4eSaM.Q]>Q;c_ORKC<T4TV85B>CbJK:I5Y_)GgPKUJ.I
@VbEF8g?R,Sc>J/cc+&DFC=?c70,LFe7:?;R@Q9999UMK\9T\N/@4>Q46N-X8+6W
d9(GPQCc00_&ON/<bOH?E)[J#@+&aDTXd4B[3=CKY\(+a#BX:O5e:Af1gDWg]=O7
@1>/RKaR<<@I\==M/U_dQ79OWO]fT(CO,fd=+6)QZP,X@H;ag/LF2e6LJ4\FEO5(
M+CI&4Y,[1&#\44R]4EdCXOOR/.b3WGFa5J,<.UVbBKYEKT]CZAS[;BVd#\IBW63
F#E4)VG9Ue107E^XdM,S7#NagYV76bM9aBNa1MOgg]K9:Y49X##DXRJ2a)EW5D9E
8Q?+WQT082=I2f@W19b0F/U-cQ[73P);#F:eXGfd8bURKUR,a_M/VL&Q9,cNBYSV
4,Pec>ZQIEK63g&NaTZ]@Z2OG44TAXGYGE9_3Zg75.L^9@^,.GGc-3U4E/bQK4eT
V?b+IJb\^]NS5D;7Z<98B7ADgGRSE@2]L=5g),6gJ\5C#b#Ha<=fP.#OcbLO@1^C
7aN-c+LDYN--aP&8]ZfgcV4gc-F1U:[&9BT>TG2Sfe.;J/QE^JR#RA^8LX2+SW9H
M<=\;(@X@a1IE)]5cM67C&GP6D.\M#K>&Z(OaCE@b[TM+_Gd^=MR(YdXX:ZgYB7]
0f3#_dG9,?WG.<]BZ.KeeV>+-BV0-[.,).+H^XYfDY<W6R9TS;9.WSUN1Y,^=R?b
dHO@RHLYRP/]5&>&K[A/GLPK3Ee--Z?8#HU.WG&L:BH:=O5>g(8;05a5?<5>c4Sa
J\U808Z&Q]fDJ-g7MP?UHGTG5GXS[88B.fZ+:PSWKbXQ(QF12K:I>GQ4,NW8H28@
7Z9E8XV<Q&RNS+Y\FW/+?U=AcF[;&^g7F].;S.D@=Ab[=#QdJ1<5&1)K;&G@5D)J
>f^H(X.GASC^4HF^MGE_\@gU-a4Q.OQL>OH9?&G.B>CS(@V7UeG.=Eb[<=\]>AE@
(ACaKWA)0g.^Va9GN9D55#,7Ja_:MCa\+aNK@Y?)D?E(HaNA_5WJ-2>)VN1A<UJG
D.T?692YC)-5Be=4&4<Y,\McW([Ea-481,aa=eHEY1cZ61e.3JB\TTL/^\=7fE4.
5WE6E_,@YA8_LS5T]-V=\Q+5V6Id3JX1U&PW->B_[@:ZELf5Me@V24\X.AHf_KS6
2LK397?D0J.IF[ZVS^44OAZ[V,NGCPMKJ[<(^K(I4:fG?4:eKJV&^=1J8>:[O?R,
#EQ)0[H@-K7@bY](>]9;N9dfdd-6<U9B5,OE/>M2,N6Cfcd@B^X&@#_a8IDZW.])
VK#\2fZ8>-Q[]9<Jf:6U;Y2Ma;>?a>T<^F=C_BGY6L-/=9/R1_1DbH.\fLBX@c,B
QT?>9A;)3?;e@>M2/8=[\;;;4/>HcB;@>Y/N>?dY7+A1OMYW,Jg&BcU2W2-3N_5c
J&+.6b,T0Ig)U-FMgIaK^8,cYA8Vdg=PAg-GI),Z-D7@&c)1+.?B&;#gNb18R)_e
K2&[GPe1STbb_&.Y?2fZ96G:12^gV9b1-]6QeXBPNg1&.#Q#YP&UbeL4(H<L^dL]
,f)1/EODGW@/I>2bHWIf=3Qa^A0K#C_OUOT>_IDL+M2+X_@4adc#]3Qd,\_:<V[T
TJA+?EDU;PW?48N65RbQ;Y+#e-\R]UN2K,F?Lcaa=S2e=16IJ7[,U;/C24>LW10^
#^25.6d-Q:+\DMO3Y+5+_)<2PHW/LFfK(<<4F(6b8TS,VW@[)Y4SG@)<\W^2GQXN
4-CE,8&_XC/_Zc0L;IA22#VeNDP=KFb\@K/RGX?1>LZ;_2@3^Td06[S.c.d4V8Y2
a_e\Q#K#/9CL+&;>02;BG#,XC5OOcX1gV?DOI4F>OO;Wb),T_G]^gQWb(IJBU-I\
e<4]^XP;<AUF7Sg+\42+DY,KG6YLSdZ);P..&Dd[O[YR]X;2@[WXbgKg&9b?\IH2
0\dGG[6YT+7da.NN8d,ULGFeb65&/aa5,]<T-U&FBg,4FOFHf501H/Z2O:Id/25K
7f?IEWOdB-T@8^4W>Q+a?.RZBF9<aXNJTZY+Q/8/DZf(M]#D_R8Ve#g:=@71W/:a
^)b_cX[88a+0TB?)&NW3-Q<13a[LKFgVULE/a,LcaFH6,>L0(+3S6WTc#0LfX=#>
d>?b):J+2[V>gML.d?SR?A^_R4?]]Ka+S,_?9NK(9b&MNd@[3(3[MT4M/USf#Z3c
<9D6<;85H-Y8^)MENY)>E#RTH/[6SK]@_0)X4I7bQ_V#B/BGPDRU#bJY@X6S>2a[
I[cPR=..\(2B&.bU?4;/H6J88YNOH8QOQ49;#b7^#HG8.VT\]A>RKS0F;=O]EX6<
L#;O[@3T#<RS)-4?KSZ5I6SL&SU[:gP4K#&U>SI)DWNURg:F,S2H;J#IAM4K=[6(
\FgPC9<4b-JAAOOgQ;>4FcF(Af^bJUZ0G4KKR_.+a92@3Oe^.AI06WV&aMGFIKF3
&Z2&H1WCSDYOcHR_^CdZ;BA.2Mdb_7FN@[HW:,].@+V/RD0.]dX;bMg;(D^U&_/,
fY7E&/BI<6IK9#/fYNUe_T;1XWRFLU>(>a=OO&\TA4@da;Q7Z=eH6HS=6FMfaggA
&8g(HP6R&F;=#MJRfDd3V/(3V@I>eVXD4<AD33-[DX]BQMHJK_[P.e:QZ6X,#3-4
66>2S/WHfc-b28,M>5LO-e7UWEXW+P4C?]Q_]HE0f\fdWT0ODH\T>eWQ>^3g@^df
0bCZT.MY6\(/D1(TWT?W[G<f=)MOO=bad;_97a8fZ426UU)d@JM/.^-<+T(Qe:eb
gV#039-cfRdE;0<cIcL+I^2cAI8[7?WdP5F^2HB:9e[#?T2GA+.]ZJ3529QZ&33@
1Q#OQ1-O#&c<fD.bW+Y^31B_1Ba\XJH[24.?86O&:R[-).=RS9TOH^00(7UfDZ3)
-LGL52A.?FJ(4(^T?OSc/NeW5>JP@&ML7#NcW,]c?KQ6eVL2A6C>A&4Z()T7[WAI
La)5-2g=?-H6,KgRZ8G,S&,L\JC30,R3X\6KUM9bQOPT27D]<1b+@:MWbQ^^DQLX
B-LFVIJ@:b2,WFC]>=eQQ&]_D]K3ETGF1V5FWb[D^CCL7Z9X-[-&gB-8&5-f-ZES
U)599fR.RH3SRO-N/R0XY9C.1W,GU<I/b4b^S0H.[UF>>/E32C#&c?Q?.GaGadO3
caEAG3Sg5Vb&(QIW_23gVaJ67eW<gbfgS:/@b4TR,6\fD4GcSKQ>E:R4fdXDE_)\
/Q4T.E]=)E5f>7Fa=UGKBTF#feYHBa0V8TEd?ZX4\\<;@Q6S088Q+\6WBdc=f_GK
G-+1<eML(.b96YQ.=8G2--[33F)f,:23C5;:Y?bA0&#4^PD8&>bOMUHVS;]]QNV-
D0ALZ/V2LCNJR7U,>:Z,>Y]-R]4^5:^AfWY,5O54JA]I;b\<Y:J/YV1P8Z+CIILg
HTU49c9B.EU<HXMX3D7U5,UAcMBUBPZ:=N]gZ0CLPFC#Tg-H3:S2a;@dL3f313LX
P>RTdD16cU#44c-dB=C.DQ8]&_.b=@;NH5^dBU_\@ddMH319]g8_TRMAJH+5@bGa
,PX)40f^FP.<+^56bfV0KA8.G,]OB7]dU&g]DYN@6U3:eCcbg7XMe[gYY2Lg^8.A
_#&M_I6BMDIMGgd0ZVO<<2Bd[,GR.\YY</K;aM5(=:.1PFFH6@WRf.Ce]08IH>+U
[&F?)EV.5c/A,Rc6/#:VWB>S1(#YN/FBMN+9FTY?(gf\DZ^Q7=@>^YGS,<-]ecVY
[>T@(&E#XN=_-)N_9N)>CZ#1)NBSbG<]]@\X[,3]b212+N<G5NW<H_+b.)O^eZ#N
+7Y][Q;)VDJKV&-4cd4IfR^VT8aGIfc+HS8JGP-R2e>d-;/GB+4+AUMbT9a^RZ1)
#;Q18C3bSM-4TJD>_MCF5;Y^V1R0DJ)ZM[R\#gC#-Sc1[6P8V##6^WRE??5N[C19
XQ4[V+C8_NE07ePcFLF;GYTbL-.e)B3YQH?1^NaS.bQO9WR;^\TZ_+/FC-C>fb=2
F>\d7RJ4B3Hd@.;HXAaa1MOVA^/A5]UKKIaB,V6H(<^dSQfDQf+CH(A<WG^0fJb&
,T-de_-Q0BYdJg..Q>a\&A(FPW5-3-6aeT#\>EAaB2PH2.][FZ?XFg#27(LLZLgH
f-Z8eR4Dd+dSf;a--OKfBQ+3:?\?03<Y(=H69-RA2+I+\1<Y95(=S)C1V<.&WUFC
_f>5@I+U&C)95O?/:/c:<PK52T+ZFGT4YPGYP7&aaN1c5@C7Y/Wg\]M>(]b([,6b
#EW@_C[9F67XLdW+=ZI=\bJg0=.VE#gA6NDJ^W7-V\GNe?Y:Pb0T>Q-/2GIPZ\3<
[gR]<5ScZeePF_ECEKHL8+2[CNKDO>WTCHC^7ff9;f@a.+=ScT=0fNZFF4MOKG-5
Pc8,)T\EeO]4LX&3)37FP&\Ic.d3ULe7#,<;EE60>R2>(SZS4#d<T6-;[,1PPKYS
/&G@f>&NHZ=UbBG52VO,Cd&CdQD70eIJ#E\+eC0XN_Bc0EdM>Z<8cd_X+NK)b>UT
J>f;@<d8f@.272@^)2)bgc;Oe1<#]BU=.IU#G;,J+f.[dPF#+=,;3YL^[\<Y#T0\
37#6B4SQ+GIL]3#U_BgSM^_CSY0RODW2IBb?KU4,5N\E13ZM:N\:0]J-JUC8I=WA
Ya+KHTA]K&ceSE2Y<NP6WG=Z4>CF/@&8MM3SLTB?_W^9(M<HRd?@-G8=FE1TQ]15
/aR5C>b:WCd/M2ISVOCJ;^c8NAF5g5DBCZcOEB2Z(d=0=):U^bFD;d#,a><18>5C
3,7YO^2ZQNMZZ;.N0NJ>Q.U_9=K>>N46T#b=3?BAJI7\#TA9N_S_dgYcV\CUORM?
^7W_/G@M7+7.>F5X)6cQ:/0@NbK3,^,bNLCM7e(DOLUF>ON,D+&Ac_e_fR)J0AF3
\^EfI4QYGG>eG[4?gYR6/:(Xc8a^D<H-?eg1W3C)CLJf9&=6cK;S=FO<Tg#FcK79
9SC^[DC<\6_@S^=#>/B@5Jc>FGD)Y>OWP-e1HNG&.9M[HC<,aIR^-FL4QA)7c@;;
F@PV:O_f^Qba_R#=^/\8FgPBIVT#N)WLGb?6)R+2)@,Hg</PHS4BJ@FA[d9B?TB1
YBC>50AbIf8USE>fB>CYL=Z<O0.fWDCaP11QTd/^T>S,BD5HDaPU14Ge0Vf@fP+a
Y/@6b#Na?bW1f^dD(9<,[=R@O,PW?^M.G8CRS_@/&XZ[[-TV?2XJ+&M][^[WbB>O
T.P\=2VK[GSgDR[5+HO;9,8AZQ>4UF_1g12aRbNO/\P):]>fC[D3NM]NG/0_?=MD
CGB(T5LB/e&S=acPV4?e2X;a\<C])g0\QN^4CTTD3Ff,Xe&<?bXK,bBFF0>?2EE<
feH_L.fX^].A[033>041DLJC)+80HNG0LL,TMDHS1AVRNA91g89@Fc0BUTAY](5?
gZ7X+^,C@ZDb0b9GDO[9a)=VF@8c1f&M@:<DB177R)WObA&X<5&UAGPP4]4e?V_D
NI6B/[^STL,9L&TaNW:[ZZYU=\QH&XaODf?JBKIX^[H?eC\E3)@CcTUO<e&[W+H\
O[ILD4?eYa.EaVaSN0=S/U.G7V00aX7:(cQ:;9AG@M#=K@a#87RJgBN,_)ZFOP>6
/K8^WZa=1P]dQT#,VU)Q_f3Id;N3N<[.c->aF9EA?-&YYeI6=._V&,PV]SB(A3^7
SCPE-V&SMDKgdGc/R.V:Lea(7LfHO&bK>)&][D)T1NA>\14CC&&1AO>WO^:Rd;>#
U6b#.Ff8X?GZEK?J2d[ab<1B,VUWI8+TRNfa-;IHI<aNSI5W>LgI[NJV\86B&eb6
cD6Ib5Oa^OT2Af3+;II:0cV-2)FJMWM>ca(1RP.@]1OX,f^?T_We_\K[&c+bV:D+
F<5L(>)fK;]1a(/Mf4:Sc[.T8)c#XJ:6KQAKQ#e(_J[I5;@/O?][I4N4LJ9+7\Qb
,/2<bBf6\Y,>OVA+RZ\F2A\K:0@I.<e2Zc7PQPD7?3SL(KbU@SRFR4,GD3R2^DG/
H07MJ?4PAFP<FJ8F5f6A#U=+J&0,=PAUGKM(-#BH89>J6XO\OCfI-AXHfL@PU1Ze
L\FP):H?d:.#(@UB:@CRGR,2DASKU<FP)05XgMYFLC4J-?Y;XL9PPCR1QNJ6R?<4
)dN\UH3=3G4EC+4e[/^#@5KbF5+.E[NfNB;9\T^/[A.&N6WfP8T=addHLWWC3TbO
cX@;>F3IT-N;GbEVJ^IVMLG#0c&L+X:+3d.RR+W]Af1F)9?b6Ef1=-Y6Y1Gd)XC/
],^WK4>f+LU^-:--9PA\d[D(T6.@#g7-5g.OgP>ZPU#]Z3[MA06YbDcK1K3S6#a9
BI8_<fC@\2Ugae[E5^UP)#f7R-GR6RfI1_[-;/c_;c[g]ZJO7I]A1=7OX>Y]YR9.
329U\_JIP[IeWf;44d.<?>Rb+WL:D^K.b7_A)\_eN(]A\L_P8X-9H2R>;BWOFSZB
f8UQMaVQ2FbQ#UMLUNI25B:T7Ye&/2bJ,[^Ja,TX(b3\dV5Y<JfE1WbQ8e>W\c\A
7^f7Q9=d[DB1<_U5WM8E[Z,9M-KBHRBJSc43F^,FPF_D^PQMWd/[CED,T4bKE9Da
f>.DKRaP(9aBSIP,^)_G[4IQQV]ObJ^>L[[9[+<0e-8-0AZJ?Z(\>]f,M>Z8g^JG
JY?<PSP[=(J,2KMV^EbUc.247#DN?\,8,\2[)OE(FW95I59PcEX.fHY&NBV#_-6:
MaeY[J+(O[Od_c<b_#I]PU@)=?2/U+I@-5dA?6EQedIf+-66Uc+I3X/+bg,/U+1\
B[LRA#\Z>f(RWOV)gD@/HLFD15(LP2gKU[eY4JRA[]f0U8O<@+#I#gFg4f@1FDSA
JL6A+TN@WJSYccfI^&<41YQbTb3cg/>]-[@g,U6,#1HW(fW(QR[d#Yd7EG2C<7_A
A=Nb)79.Sa-8BgH(R]]_67HDF\4:F9@T09bfcZL5J./RE/8aTP>Z]@(N,A:82CA3
Vb@YB@@BQcB7:#dL@L,4;_cV5LCEEQ>F3IL5bDc4VdRF<10Z.+X3_=36^01R07=U
Mf>>NceaG3=_IQ177c8M21+0J=I/O>S#Yd.?:^21;^E)BeNB7=(3)\6O230\[b.)
c81bZ>fDL.FbA6\F00=/a:RW4#ZHTX6JT8_)77I,QaB)T&[Fa0N.EbV_\EW8C8<G
-egQ6G5ed&SCRIH4D^_?Q\KJ]J56V:1VfR-X9A?Wc4LY@W?VWK_U\P,Pa?1f2@4S
(R7@[=^D^Ld9XJJ-O(XDH?e@+IBWRb5UPgeRfMeN;\D679cUMM-89H(1d7IR,0KP
\G_R26_YJ5I;]R+<_>C2f/4+JJ7<+[I[.4MNDZ>?^?C@5g#C;QPBH@9T\7\QN\<F
@QYUgEJ.0?0SP_K;g:OH0(RA1:eRd2,<5e3dGHGE-M?L,EM:LI/eTdS^:a9cD3_K
#Eee>;gT&;R/LZ)76cJW\];#DGb-P=,N7)P/[LOH3(#3#42@82R[5]VS;Z)9R=E)
N9aK0+AGdTFRLS>8YANcM/:&cW0>ca+V&N_6C)K684c89DQ1]1;?_TSIKO4#707T
RTJI\P2:[X&(CK3(ZFg2DH1>2A,05LB=(J^662@:O1XG</FMO^.9D4J_3-3DC_LC
8BX1#B1LW+(0b3LU7>#BE/X:31f_?-VW_FFP2MN35H6bD;d#TI])/ECON]aU-3Q)
I]0YIROa1B3&7MeWLY8,]GP5E;G&KLJ9A9dbc05-,9f)E<JU85/2bWR#)+Lf++Wa
/)LWW62X#[UB?Q+&6+=bY6Fb9IbD8NWbdW1MZ+f\A5eW#Z>ad9Be=?P#LRBH4(]E
8AgY2DN2A2>2<KU#;JR+2S,Eb]YF+J)6bECfBGYQ43^WG]?^g)gb7<b94?0f[>\Y
-56Ec:J8(H0;R<K8]N<+@\VfKOf,>3MZc?3-NFK840Kge-fMaQ>E<9SHQLIKEZN=
#8E_WX/,Z2eB^@@\>Q,M4XDd<EGX7MVV(8H<d8bPSDeZdd3@?JCb(dNNHXK=DXKW
H8&c1?[+&(I-eC9ZCZ0CbFCb^;#HRe^f54J4BC6?[d(BYaAc:(V(C6)aUKfOF3?b
,LYHOX;,3/H9[_++K@]LO4bT1F5U.>Y[##T4,LW]#\7_?PZV:1=H4VP599._-:.^
UOT[<-gBTdD-H&TDHQCfRU]a,Q@=bL8EGA1W,O617T9;5@,fE_0P@P?)@.47IR<D
IJSG[FDSSGD/75e75L-\OM\5+b_CY3ID:U,L>23Q.=8JHX,)P>=B6S[D5YKRLWC0
)fY((&YAQ)63eX]H>Z8Nb1EST=IcN4(Q>#b,VQ.>]II0BJcfU6V)geQ+45[;I5K4
M);=.<3DBb[NHC0@+^0KKbNE5EI7M@d6763X<DRPP9eJ7IXe\a)G:JZf#\)b[/[;
5J0(YNA/c1fB>4BOe)]WEM+3fC0\O_](P?(&XA/f:\[ccHE&_DBDOd-4Za2Q;=JT
NAH0_25\#CJ:&7XDXSG38SJH+H7+<B>@-RTM7Dc61bFZT31fS(4MO@N(3X)3Q0G(
9;5GF]QcLK7eX?:,ZDTX)_00bM@FKdYS.;a1WI\[R4=U[9N)C1@WA7-OJa.K/Q(Q
_=UCb54LU1<K[Z)U3DaFLAMHRNM#?Z-gU?G#6Mb&c/\8,TX&2NN5DF-P0^7F--F@
#]@N[C6?GS/a@3ZRI<dQ-^Z9#KK#d21/>O^c9,.5cS#LFEXJdW97#UUC#2OL&V?&
eS=U[SC]Pd#W92K80ST6S25&8f0\#Q,S-1E0G\&J&A:Z+>;W?CAXSf&YVgJ-N:-D
e3g86bZQac,gfDM0cW.LPMK>Z4SU<&=\GM:#1ODP?\:F>d9Te=R2>ZDd8)2-7G<D
.G:FS9WG0FTN[-:K/57<W?(,?<2+#N[]\[8aYN^)0DB7GI=@=+>8Rg9GL0GBbe7O
NDZRbWDbJ=,VA6CJ@?BHIUU,=,7Hb;>FZ>B3]ZT)PTc95^(L]e\T-NQ:8H3a:QV\
>:U?Od[)P4DMFVb6:S38VRHX[PNbNe_DKd^MT9:#VVffET0Nd&TORdJ5MVMFG+M2
&UaFa_I^OD+)W(ALX:9VV=X2)R/(\IDb<K/1G.8C<&C/>81HRE:HYGO\T:<@4eMV
cTfd@Fe4MW,?-2_0\_N_H<1_,@N(-dK6OD0T<,VPcIC:A>],)YM[A,BH4IOX.^f/
(P5NPV\,Y,c5aLSEN;3b-aK05_,8J;-,AcaaP2QMTfMBd>C(YJ637.BEDV(BD)PM
Rcca-?,4?(2YT56SAN<a;+IKg,<aOZ0X+RPb;V].G2X@6MbaEXKVEU+O^6MXPC>R
A.Q&B35K9T3W#g^5a=S/aX=G:.>Z&>7Sb)GgH.(>AF/:;X#LE3&a@IHJCZ.)J;M]
:H=9FV9^\2#VJGXWb1[_V;JZF3WUOWX4]MFR9=LB7#/XbVNHa(SA1>aeEWGPR6]G
,7YO5a[.32UO^5f?X+F:4]eG^M38HRKdLMd(56:KGCH/N10O>Ieef>9QNY>fOf[-
\DT31Q=/]D7+.<2XB[Tc>\@1ab,7<eS-59].RCc.[/>MA[&ZX6<JgU-6dXM6[a^\
+5-=P#NAR8U<T)X&5P.B+9Ge13Hc?R2J)M(@N/6<^(B3Q\3C:d3X7f0A/3/>UY8[
F7+^=0<_2dcEGgH64RBLIQ)Z2)-.:;=dDL:B,J\/N#cB<>YHDP9QR^<,@-=8.3QA
EGQf)^cXABRCXKLA_Z-edSf=EgW=;AHEBP=PJQ4=6C#a=a2>3WaB#aVBHI0H=LU+
/:a,7c6)]8S6]T/af@C\1I3[0_,1]TN0eI+)8W0-1?8+V9eOA8.Gd-5=G0ZXA(./
2?@J]DZT\]&_(V].A?IZ3H99Y#FWU<-69f=W=NTc2Tb)6d7E,QgC]V2K>UWPYC8[
DQ^GR1>caAcCW)7_G/9+I)C:aI@H.4KI-Z]2AXdAdZ>.I7QaJg>Q9538&:041J8I
GX@Q&_e8&K.)8aM:D0<BED]gAVK5O7(714DN#M_Q)2#D@cX(4ASg(:bDcMR;(cWH
;M?;&d6dCE_&L=e4TK)=\_P_@O;76b4T^_eb,B^;TD-<MZ1_L:::\d0,7e8(7_TZ
-/X^2]LXAO/KN-\cUe)?,#6\Bf\EKCL87_\P]B(WMMBFYdV@fEZW7cR4XR6YDT2T
V4Eb<_6a9I)^/BW0X=2C/=CA1@0X0I6X#fGSWaQIVTQ=78ORE8U4<NX7Z8N:MW)-
_X.^[_1SaOBTHM/0a?>ROI)eGWXZO:IPS&C&K[X^?G\DIFac,GQcL]Z0GT>e+2KD
,+e[=S-U4/Kg-Mg4F/-E4fd+IJA(DL@KQTCT@Fc^D)DfVYEBc;Z6&/)X,-_5c]C/
H9Hb7&^2LPc\1Gf9[/R^MNHZF1Pc5U5B&SQgRG9=<0\5d\Z-XEZE#d&2^6Z[LAW[
&[B,,B/XY_K:\8(2Mb^B5^4edg6(cC>U#04IT=fa95J@0]\/P8AdY.9+BYea@+EC
MM/5A8A?0252J4Q73ZW>BBfdEA;@L>0#<?\P1AL(YC4Bf\?=&J/2LXTZ@fQT&9:6
A[3cWS)WDERK8?9V=^/gd?KT2ZTEL5\-^IfAL/@5CS_?9/VHU^^76G)&V3R[WdZd
]=3R/U42Q]UO]a81Z8\716PJcc:<TBN//QFV;aRH;_LJOD4IPfYGK;;,QCeXC^6.
,RX7M;)RKfIbY))#@TZ=f@A/-@Q@?D\a[HYbc4:fFMa#cSXP&Cg\N-WeP0ZY#Rga
B:ZG)?=CaX)T\Q@<0^6C_CHcYSaZ]A37C6Bd)Ma&&AG6e5H?<-gO14_]-]Z(VKfb
/,KY624aT_cQOYE22SC9fDA]@/,B@c1;,f^=,]?>;I>+#c</R,NM=0J37BRE7:\K
aM+:3=CCeCF3^Bb19.<O4gGg]f[+EFPZ,a(0Q\B/1dP@HJ;4a6(F?369IS&OR5_2
Q71?HW=e2&b/U+>.@c(U;#<6ZZ09)398JOR<L0G@F#5Qb]g5=0P4<#&+WA[YNfdE
2J=F^@dY,7FbA_d2CBA[^RI=:0f_db&\W-P8Y=CHSG4/URaXEeFd1)+Xf(;O7=7[
=BdNK?+D/+F]gN=F##8/H1gT40>)dg2aW/#@g[ZJJJ,XgC+,MSEGfO^N@/e-)>cc
0;&gK,2V4P4T0HF07Y)+E<O&RG68F]9BBSMUCZA<QU9Z.=Q\^YE)T@e<D:[b76T.
.:RSCYdHJ18F;WOdF(+/1H&5\>5#A7&5X&TGZKZ&TeF[GEF?Z\)PKU_&aeW3M)6b
g;Ic-_PV31J[FbNG)a\Y[00EO?D>Q@,YZ,cU^>@HMYAf]V7O);P,--YIa23GZC>I
A:=BBE]3/PU)^^Ccc-PH0RDN]P1WC,EcY.&+.db6EV-B5IJG;]bCN;C.8GTJ;,#[
=]3IR5,TW(9KGCLQMaFA3KJ1U\@6aE[A\+FB(0,9WGU(+WAV<M^gI[6]FQJQ+\QO
CVW[-;[S,_..eD9c0AR<P8AYCO7<6^JWWVSEd/1;K:-2R2BD-_M_CXXMe7RNC)61
C+;T0Z[dOGJ4X&\&_f.1JE<#f)X2XGUbQ7VR_.(Aa<=[;A\YN.+<56_IL_gf7,<0
/S_WNRIO#KET.]NQQVbB#O_G6ET34Y6H5+_&DCDF&/7\=HgT],X6L7&B\Q>gA=(P
WO>OCA;HgRHO1>aMMY@)X6/R=D0,e)J&ZEO26@)E?;dKNJ;I[H#U9WWW[WT&N-d)
V;1We3.aW.<f@HCF8ZMVbEQ+.AD651@eaeG.GSJdUfT(A6^3?GYAUBCU=9-V&WN>
=ZADU6BX\+3c-I;Y#W@SI>Jb7O2U\4,_)f2fJ0>OX1^_54U)FfEMATX&MLcNA-Ib
R[agGPN9_F?H,S:SH3bB7JKWO4\JPMR6dGS#UQ@:,Y]>[BZ9J;Ybc8@R?FYB/R89
a]9U,850I=gXfZ[3.J-FIaU=U^@,OY1JP-<6,;P^)IHCL.FaLA41NJTbP9K^MD2d
>V0gKRK,8\(1,OY3?;XWGCM.cV&R0;I@<OC<b.9MV__[Xc85>1b7C8?;Q-I9,6G+
[[NOOX(ZFK<cG5)RIWO++9:e-8XKgNG<1<a@J)@#7:+N)Jc1-T\&HZL>ZfI/;&GY
_X^KX4;.6_.?.b55+JC(5J8f+CeD+ddI?e=[eTUdB?#9-Y9bVd^8P>6C3DOK&2R+
,SW=@=PL350ScBVg^WAa8G(3G?fGIGRR6YcU/WCTRO9_&5f#(.f<?ITJ;_g?6#6#
>)VGQ?eb3ff<,V+OX5bRRff).N)Ze[S6U0MG-EB+SNaf&L.LSY8QFW1gge?2>YBG
CS@PF7Y<99b&W^W.dXZ48\7X&\I;gd)9EAK-Rf3X7CZ[]^b-<[=X#8F=5;?FdWSW
=VKD_QJ/^fZb07f<)>DODPLadD5;3GIYH_J6-DCK]2+/S9;5aBeHR#7EfcLJ:#:a
5AC91I/9W?.Ud>4cR9^.BMH?E)M87-O;[,b&c+:gFI=0A]_^C@(4?\?OUYT.?TFC
MbIg7&(=A64ZXTU90SY-?D+GbIa^bQTC@9XW4cG3Ee=QXS1I#9F-I[<:>06PA=Mb
9e<H>eX.Y\Q,#.87;Q6^0eP@^P-378\BK:PG05^g=Xe7eL[B0L;#PT_5R\e-;S3g
]/+7[F9H@?TDOAS4eDb>5T1[g<+S&6d\YL(SHRICCA_Q@F_APfKSX?GB>>(TS1W1
4b?49[D[NfQXfDY(Z/_.cF/_)KIRP+/;14__f@<CVgY><D-bIAN;&/L?dDceaZ7;
1-GM/93C[>4+g@09K-;4RBVcFGS<=XITeB7_)Z)-fd/bJ:Za?04c7e3XBB0YM8C8
<SRd9#LAb6L,O:[>NS#eCWgFNB+97A@E3BS-(d&US^]AR1.;GG(#?&J-(IL_;K+G
-Kd]A.+PASRJ]8K31?=FgaOSHaYE/HK[K+,aKKP.[?DI+MUad@)1dZT5(L^4U]^Y
X8e,[O=(O2Q.?,H?+aP)MB]>AB<XCD_Qb2>g=aQcg?V#P)d@=f4g;H7OC4aSF#Rg
U^K/8=caPcO\A<PBXO0\MXFOE[&-@L+CZN\.d2LSB4):M0-g5HG=?B?].1FHS:87
ZOS35T&dV[Q:aZ[FP9S/+,MQ8HEK?C[I,@ES+EFEeb.>.0P5O[6[ZH>E6cWQRXWJ
7W>F\M@N])g)LPAJb;/AM9bKF8_6?ZdHKHL\#B_>7Dd:4C6HG[_gb[ga98(c=McT
X-N4B[TE<\XMb_02c@SQ.#Cg#gbDK-YC81M.FZ@Ic1@,e.H3];1_>E2DfP:D0J&C
>5B].N#9OgDLBGZGVe)N)V4Q@<Q.#4,?)Cc6d.ZLZcTN6K=,CcVCJC8XO235/Z=Y
I:T\56SdPLfgW=X45M29W.c?.];MU:g;_-L<GL,Q^4R\@DVbYZD\V^0GdKWD61Pd
.8b^^AV)=^]=X7E7T?eeK@JJd7d^R&7\(8R?C<fU,4N<IQY@eXa+JOg<:EedW8@]
K.AP@9C8D(>_J)ET/NMN(_BA.]0<)XGX.)GJZGMFXYd<C$
`endprotected


`endif // GUARD_SVT_AXI_SLAVE_MONITOR_CMD_OVM_SV
