
`ifndef GUARD_SVT_AHB_MASTER_MONITOR_CALLBACK_UVM_SV
`define GUARD_SVT_AHB_MASTER_MONITOR_CALLBACK_UVM_SV

/**
 *  Master monitor callback class contains the callback methods called by the
 *  master monitor component.
 */
`ifdef SVT_VMM_TECHNOLOGY
class svt_ahb_master_monitor_callback extends svt_xactor_callbacks;
`else
class svt_ahb_master_monitor_callback extends svt_callback;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_ahb_master_monitor_callback");
`endif

//vcs_vip_protect
`protected
CAb9WU=,U2EZ?3T2>(gA8D1FJ49(ZLU4bORD#5a2>1Q/CS[G7E/Y((7QV)5O(CRW
.&2=Hc=J-X2?ZbH:^OEc\K.1U-JK<-PMeHIK4&O),#MMFOV7VLH)]/JK;,02)a.#
:Z1:8S7BVI&X(UBeM)77SAIc=:>IfG70FN1B=</+1H##1ZS[L>GELHOb_^-a6e++
M5B]7D>IR/R./1/S.ES;6Ogc135b#XWIJ=W4E1aUFL\dND-gJCNEG279cAE(Y40D
?X-13;0TB8[cg#+D-5DIaLGdEIZfeZ?.)0BMe\(.Vaa]?(bXS)30d\@65L9OT:5P
H9Y\R-/?C-L>KVg<CW6>:&P]7_dT1CcW0]LM[ME?]699Z7MHd.D4A592\,Xb)6]Z
Ud=e_7QA>4?O\U_AbDO[<cKG,SU8&H@4fA<O\KeE9TWDd#.be3U=dO[XB35ffc8M
-9WI1b<)(1>LEB@G61/IGTMETU2JZED3;W1cZa^86O4T;(QII6KTK0W)897O3A/Z
KML:?7LT=TAJdU?HTA2N79f>MUIK9VH-ZQB#)3KK)SE2B4?91PVHY[(b^?)C[+)7
VQ<PF9e-TDbBIO(9:9A+&;BXSF?U0AF+B2UW16ffSY0D]#KQH)1[J6KAEZ-MaN+F
.0OLU.:I/>,\fbAZJ(Mf,/ZC]<>ENN.B)?2M9IS&L6>2FD(NP@-P:U4U_adTH/AQ
FOfRfL/7g7,-L\IQ6Ob\UG4[b4?JfbVX,.1.R(LQS12JG4,gfZ8:GG][[0aYgZIb
U8PQCD=.GN@T0ObXWX33&83]EF4-I.-N8ZI#C^MBbXPH94EB?@9;VD_@adN^O23g
<^]428dQ2:PC,=SS7&<#9/4)6fb2CQ<JDb.ga1aL[0b_PTZ1YJ::SPS/gC]c9L):
667#[ZCPEJN7_E+41Z3>cR=.eDS,QNIRaJ373.O\g]e)>?4d^#<ca#3DINMHUCSK
f[^^C<]O8/a41H52]QeMId:.S#T(_FP\\+b>.L-6&\IZR,)IaS9L>--&JJ;R)C;F
:@P<A)\d,7Q\1;]T8G:Ab#W5OH&V?\+N(+3311X@U<UA9F\EZgDV?J^agZY#XQPg
e>-W;8#QQJTg9GM3,\A#2g?]KG/<1=_b@aMWWAa2bLTc/2HRG]GM)]D#MKYH,JO?
]5N95]5Ob:d8M.F27]bZ5415+3K,OXP[.H\2E8eXOR&NNH,+,+6HDNZR=TQWbPBc
_OI6#68deF\@6C,H88f[H/N/@)XgWZ7=1KCLGLPBB/LJNMAY(HPT#(X>2J\9e(QL
_TEQEcF1Gd-<T:7<X1U#Q7fd_d]WXHGN9)(YUf:D&4)&#Z3S?MEa_KLJ/6)D/TLZ
IL>OeR@Z\g45Vc,KL6+bX9bcB&^.;U-VZ2&aS?GD-XU,<_FH&G,bHF=VXDICCC[^
>61#Qg4YYN/:SMJ:BSO+R@PI3;110E(aDXCLEU-b+VS.cJAP5X8BPSa746A9cT=g
-P;EC69Y>MMfS:3DFZBbLXN^25/F8F51M)8?+E]HUOL)K8dQTIGA_dC/SEZXfQDA
9LPS2OJ#6D2DR,])@Tc;e[0IZ>HNTX+G1EDV^@M<McAOD=ag,)5PGN.=dUO0,A.:
MLW8VI>F>0@7fU[A](U69?U@\,bV]c3L?GWWI8O(80OHXCS8=QH>dIeQ-883/e[+
[]W@D0CA1URa1?,A6c.eOCS[O3Y5,MHA)(,>^bfJ:fOM#EB]?+N8R7S?F_YBR0]2
MYI/=;Zc@GfSQ,8)D&=^KY-Z6:Ga2^^LFcW[G6Z_(=V?B;A/?7HGP<[TS[19;YQU
^[/0?RV(5cCd;599:.B5NcAVJRVeHRXZMCOVL[7?NU:)+CZAQ=;^;9_WH6_138e4
G&4.=:DN]7dRdg?YWIX5.G;V;eb&5GDR9W+=DMQKc+a_^cVY]c\7=\88e;:HU;O\
B_cCGcQ,fN9KLSD3,,^d1X.0(eGTG3C5[9RHQb-OaKg^.+d?d2#Ycd^WICa48,E8
^6LP8bWH#T\OG[1_0M[F..K+@N495(G8HL]8:SSI1M(Y;G46HOX1I?E.W2O8#E#\
;[F+G/8MfC\KOEI_\efV:G-ED^YD38-4O+N4R1?Q;0fPJU)((8(6G1:2Q=&b1PAR
dad,FC6=4JEAEHa@M;@&=DP&XHQ#?=04TIUddPdcE\;5&PJb.A&O.(gZQ<IfGX0c
M8<.ATDBfFVb4eWebJ&^(0D6@Nb^d1K=(65QM5FZ7)Z/Q,HF_N<]d6bK94.8[P5C
-=Vg9N1E#(LU/]Ba.)c_P^TR43PG]FRDCb]7O^SXV=<S^adDHJE:GI;<B0\<-gc4
<+6J:^;4C0c2[Q,UIR#C5;SU/A/#@28X>K>]Kcg;]H.1WZdZ4-f=XRWS;M_PLK[<
f0A0.@):X[f,D,F-2&9U2@0FTYRUg,.(dK:;.f+TT=A+M,WeB61a,\,d.8&HG+YD
gJ[VI+0<82aTW4+g+X]XWC8J#ff]4G^HffW9E6R1Y8=;OHC[=9@/BA>9&(aMRUeU
f<HQE&N_fVV[-PB=5\/SQ-K;?52/&6V()TEI=S0SC=VT--+-@Cc,^)J;>(D3AC4R
Sd>JPcW^4V/9<]DR38bEg+U_RT.#+]))XO;INNQ:Oe.+R^TOAJ,\;FgIfG1g?6Lc
-Z:2]HLQfTAHLKO=?PCPI+@6[\Z,1ZCOA/A./?)=974C1G5RPZJ0.dAQ+.#,X/UZ
N/)0W/PYM^PNNXXU5@),[MJfFK,d_JM[&=ca25U8=8O5.4W\I6++70^FOWXD5XJg
D4VRCPaCJ]Q]BLG?;Z=dQ(+HV0DfKM[&T?c-_8E82K>,Q>ZCaKUb8J;Y3/+e(Q0;
=@5A)</HJ[XdHI6:@baQKDdL-139bT>>7a+2?Q0)#2B706(V(,gI1,]IY6Ke__9,
f(;IDV]C3aO7RGLP20_e4;aYVc?2^eU--7PF+NbQ=Q=O/,&5G&>7:MHOcK3@UA6g
CA2\dN294](_>2_YPY)>8#UP1:,KHX<@?^KVcP@_K>7<L^JO/C]_[U.=[A>,B0HH
f[Wc_15E1MLW1cP@.>P?bFUZ-PJ;&<00_ZR#.L]AS4aQ??JK-DeFBIARU;[2/ZXJ
)I1F.AN;R,?+<5E4UX/H]VU/9T2VXU=\Pb:HPA9daNd\K=7O^MACWG@=R17f(/R)
UbMd.Lc_FYMC^FS^)?TfT\:GC>QY5Y^32U8V,3FUEY-T#2KD3EH6OV+_b]:IZQP1
(gR5/XT_F3]>C=C?_\FE^0cSC\WgE@LRB)G.<>XZWI2H57ObW2HFQVT-?d8a<6F;
2_CT5374&-4X\&2:.H[)eg3I0VBPgPe/?4e:::KA#_=E;=bf&F-Bg7eN=K0R(adO
[8_(g/K]3Ne\a3C^@7T-VS]8@M:Wg#YQGI>B8@[K+(B]FK__;5O]dgJ<_fGAAUEK
,\Oc[A8W62?7O[)XLO<J;5J763K:TdDX7g<<&]OC2>eMA81\a=Y_6a09-g)AfU/Y
Md[[3e@78_5eZX,@3D3E2f<9XXYd1FF)INP+1,=TK^R7,T^>D1--C3GT(P4>K2eT
6#/IP@-C@H297HNC?:03NH#ZWTZH;(96Y<=+eYVHN/V(;(V\QZXQF-aAf8c]YR>:
N(7A)C:g(E&9.KB7H8Q&:+N\37]/B@ERVe[YHOS51+5D/:<Hg;2Y/C;E9Ab7I/+#
dP836R84S.S#D_,eJF&J3-a/.Q[C5WbE+aePe>E+D39^#\g4P)IM9/91+;KFdfV,
cf;^Gb7F\H>/DF4[-[6;O5a]TG+.)O>EeQMV,P0F,;EKM8PV7(6=,&E3&Ceb?fIZ
RBS+Gc[41(/B[f;@ILV-M3OVRSXR;=:7.^;,>XBNROg-@c9g:bC+93]5TP+8GY@e
7U2,:_ETF9R5bX1&FI?<F]1S6-[V[\)U8[=)\X49&Va=D1HRXTLJ+bSYKYK/)d7e
\F,LdBd^]JFPOb(C&(afbMRf,cF/GVHgJM4#IUfM3C>CI@Z0D.RJca+PN7H^LQ8[
F/476C#S:=[-J]cZI:0SV48:f44E0<@BG\3R/@e]70X1_]1&E<75C3b1<+Q0E=V=
V?)B/BDS<=OCE?:,?QCaf):e2O;KG\&/#^=J?+6.4A[&Z=P0PZ0B6([YgB^^9;-#
?_c&;e1VR^_:I8YQU.^<GO(_L6aSO+(N3ceaUKfJ:5O[2T6:8+);Z44:3RS&[E+<
dBJaYF[I5F=DMF:1M]N)-0>>\=I/6R&:RMADb8JB<4#5+(Y<K-fcT71fL9<]1F)K
3GFXefZ1TCE,9Z-H:#KeC4/R:Sbb7OFf3(L879P2c;MT#G5eOLFcV-5ARBFU3SfO
Z^H8e[LQ(<]T):/bb2PD.H9dGY.Dd?B1OQ5KED#6S,fB>OY2-^MZC;JP8aE<TC0T
a_.MeYV]Se[N-5V0:3-@dbE_NJdKTLKPUM.adfIB+WKf_=QRcL&PWGO.BaZ@TbM5
#TeWJDL,+G?.[?HEJ<cdW8,^G.+N@3.[D,YMbeQW_#+&I5AOM^A0.90WEA29\>ZF
8N>B4;JF_,@EdbWS.c3WP,QG5dVJ6OCEB3S/_Wc]Y=:B-RA0B2bG=Z#L2]@-E[RK
E_Ae.)c2AKeP?VQ9UGN@76P:KVB[0)?QfQ9,58]3gWARSV2@KPbg>0d<9f^d;]F(
fYCcV7<4+H92I=]N-,^I=Z6_03Lbe?VA/S3:72aXe#0P&_\<)EA8:SXL3@UKZ6]4
:fI.GA[\+D74)&BR9B73KgECF=(g^0PMVSa?D8L&GS22;/FW0=_6fTSaCN-VW?]1
)E8I/R&)b+T1/6@2@F3fLX_7QK741Z]H:GF]I0T3a>aMLI&[HJF.UcYf8DLbWDe^
e0E^TFB0>>Q6IH<FKRVgNAa^G,0MF;:Q6R=9:=O6(5/1^G&[Le=_VK?0-A<EGdE(
TW/F=LGA/PN6XE4_T?4^]=4@Lb[2fP0/[],4UMPH43MPU&<7CKJ^YQYf0/4.R_32
GLd_K7K4;JeTI08-S+==+,@8abSZSWP?TgUfQMD)&?adJE+HY/fVB3dIK\;DbHU]
D8::=,b#TWV9(M-8(Ze+AABTN&>_,D[<KRUT1c2YHO60gZ=]IR+O?(&)._^,?E&\
:49)DXM)[B]g=<N2Y0H,?;M/BK)[6F[NP1e7U]V&53b7PZ1fOPZ+Q-LB=D4QCad/
V->#DV++PUC0+.VR)JgZfOQ@NY9?)/7/W>@PH(H3X2N?1#5OV(?\P&692R[+4R=K
F7GP52>J0=S@Q91@VK3H8=):QUeQ0RA,T2Rc,IZ(Kf8^UFM@7A/]0fXVdZ=50e/>
M,A(O,_TMV;/.D7aWg]T9aV01&-I++D+HJ(S;Y:Xf@eQ\(YRNT>0f#aBL\OR3QI_
Y<3g+WZP-4J3XZP9MIBJY:X<TMZ/_E9Q7_ENT>9#EY/[Af^g0ZSV,1X5d9(#L41Y
SN84L2EBfccIVR(QA7ELNE?(N;7,H_>?]YfCS9Y7<5?7QCZJfC<VM=fU/=84Ce.P
[\RH?AN/A>>7g:JOf0DO4d22,Ka>b.3dC]L9-PWXaVK\JDQce_[&10DAS00&,#2C
:Wf4^ACSC._[7G+79OAZG+Q>Oa[AZI[/TH-\.<XdCe1,:0ZE?E&g)(61.bY-JW3I
N&R=)OYcg[9UD@MGb&Z,[+3O5C_^2#\Wa@NdM20&7V<C>,XQ9T<:?#E.D1bUW-LV
0RW>R:DJ@.Z+_B66ZTAbMN0Q9I/Q6^)K2.C9G?f<8MBA21Z:)Se.,&RB9Mc)ZeAD
@g7[X3>7N6+F3g;R00+?.ENa,V[+3a+?72DgfTHC^8-<aSeOUIF:KWc:f#c[VZaZ
6V,I3\.^5@(W[ee\K>JE^-FcPQ@^UW^Weee[5FONQNRE-H(TT7QY.@O#(7EXH7&c
-8-P?e_OV_eXQa,9DQUEGB.2V7F5&@_SCMUHDR#K86=Pee0c9O:LS65299W(@bTN
0+b/:-HgK3(00>RNXGD1N^[@1d8?2YMKDWYG#b.QSB?6&X?SH)IOOX(A&E(#?Y#^
PYA#WFc6O6SCAFW]#X2>RY1FXLc.;ROJEWXS>d>)<cg)AMZ:N)gJ[;4-UD3fS^_S
(8Kd2E6+dWWE/R5P\50b7V72\94\H&QM1;^,aWE.WHVc_&H+JLaRPE.?1ML^TQ<=
1?,56f5<+_J(DdLM1bKPDPS3)M=T@<X5A1.4VPdcLQ>Y5HC)CJRP)BXXG?@_^c2J
4X+D+4Oa704ASR:Y:V=S-d&RP-RV9#20UB/5)<.F+#R:Kf#BEaL_P)Y:Ddb-UNEZ
8/-@IQ)dH],ET30PX2Y^QNeX;W)RN4502EOc(_8+3:C2+FOR.d[[8IZ8B;TKLU19
#fQHPU\(>L3DN2\DdLe8]>I/,KVL3G;,:,62K41GE/NYL^bX^DQ7SXL9\aQX^_^O
6/-BG8)GDPII+DUM(4B>)-Ia@LEg?L/b@AcK;I/8f8TGEd7+\@6;,-5fBfRT,KeH
)?UOD154A?.K]Q:8O##<\_5.H=YXU9B/Re/0MT_5@=DVX1.NFDU<=D?cP?&eaSEO
3#[>N9(YOeDKCO(4OVSG_Kf0+Z;Y:K12CR3V32Q5>M6Y_g:6f)b_L4=_e4PV0GcV
EP=E/)U:\=HI:fg+X54M>VSdXd>c>>Y/,P4Ee0]#BW5Q>5+Hb#&(>d3GU;]NN492
gL:TcAfccGZL1Sf8^5FL^2]BNIJ9Wcc]5/[YO(\=FJE6_Ub]T2#C.X5KJ;cI&K9G
Z3TD(QIfYaS]c5a,D=^5-]I21NaPC((44Z1R,,?Vc@[H[>QJ<]:(7Z17>4_Md-TX
VBLYDU6M:GI0L=-GY8.U(_S(G5.0@3;RM-.4>d8J5b?bXf,@E:W?+^/OE:9a/PUO
/:KL#54^a:FW#KGZ^-a=AJ]\e\2Q1#8dC\aAUD)g3P5#gUaH+=5L8/:c)?0I9Wg\
8MeA9?NTG)6MYG<-<ENT[3g6=6P=De;Q0T#YE\Kc\3G@B^ND85(AdOU;+8NY2a=3
2\UaXU3^I[PZ]:.L3+=3<.YN:MAOAeV>0RIZOF^L]M(C+,WKH(+)>GA_;+SL.MA?
8/[RV0]3Ta(Wd\Z=0PZ79b(TT;^9XIR=9>>^.UT^/9^Y>IZ[G\E^=)<Y:cbQMd4]
5/;?]e(:ZWAXIUVO9NL;OaT1&V:(c;MJ7H7N3NL#]FS7PE)RX3K.U3C#2W+S94;Z
&JaHeWR0)I:NI\d/]cS_.bU1#?G@<++)->,6F4BR]=O;@(7I.,L_#^\SbJVO,[8@
/\97#U>bYC0:4&04N.d]3BB6aSNDW3>:N2G;F0SWgPICc\AbADCVf1=g;F0?I6I<
+SOQ@Z^,D:V^8AKded1.O)f_<UIeSc<c9B+GH,^3OJIZ#P?OGLa;PZXFgC7EWFI9
U[4IB[CWTVYb,M&7M(abg@9bR\4dJ?WO])f+YdLAQ0TU.AU-dDb:9/:(TW#UHW=g
G-B.F0WJ1a_EJ.&)VK5b,JMcUYSRgOC(g;b:/:^LE2O:7Q=FC8-Jb0c[NVX]A.?5
X<J[cUH#[NVXN:Kb_KQc9ZWU8VI9CI=eL;&dZQBGf@O+UPd/DYP4L1Z/:C5BcN]9
4-R+1)YZU8@d0A69J#^d0D\;Y+3+GgMB1RO@9Y=#16dH25VZ^-G91^P>/5B9H^.C
5Tb?3/.YWE)I1YI_AA?\gK4L\1bD4+\/?.5UQHGI]W+Q.;Cgf8d@BQOD-cbb47XC
SBC88:N;Ug@M;T7/G=Ugbg;Y.UTC_+W(_C14D-;X7[EN)ec^,7/ePK>;aSO0L]4-
Y<M8RZOM41U>K+DG(HREg5fLAYJaDH-+cE>/]G?>T.CF=5T9-#0fb,U#8<DK=fLB
UeX]D[YB>1JKZf;CJ]X993_RGaWB2^#4cD(cF,d\H.600c\5C^??g?4U5]6PN&EL
8fe<V[G+<KSI0Z[C+/PIaI5aWNd8.6TMeRP(^K>L/1R</<F[WU9#b_b?SgL/AO3I
Td&)9gf<U&\1F.S<IA98G5Q&WN=](g#KJ87MQ3d^SX>a360VIf[+4Z@9Obe24D8:
-F+HZBB89cL/0Y<X6XXGcQ/ZVdSGAVMVAb3)#WT/VWeCIaHPT9_II4a]\NY;7bZG
c8c)[NDaC[X9V)#+gIC^IYPH)d#@M=-];IL5>EObV=(;:;=<(L0_,gZ#PNVAX4O5
C#12/;g?VO>=KW(PKEY@CE-1d9.Y+6babcZAN?#R.,KJI@9#:@(AVfF2@:\=N67N
UA^RAK9cH#-ZH5fQB^X_,\/&[a1+OP+gMX:S[LI0BF9OcG.fCH[eU95R4eYSfAe]
b9#OPgdMZMFECEM?CS/(H#c+MVG(9/HJL@cWed)9a)Ya&f\ZTKL[,G=:D01cNGcG
QO[?d4Q)XU<?82=fe[7?:J]cL2_^-GW;R9C3@TU?P([HAE5X:aVVW<5R/:Rc0>MH
WXFdKYO+e2.KAY8XBG2.@?d)P5XWW]6+Z<\&Z/d5RH)6?.65Qc>+f6/(KKL9)D&+
15\S)5#=FCP2#5#@XL<Z4W+.STVU,\FPC2HXe>a(c@AgcY8&+?8X?7Z^QP:b[1X:
:#,B9B/D4M@OebEQD;<^VQag@U-U\0/-T,NA^U,c>4/F&V?OLIBacV96eLE)aA)b
J@]X3;WG)M/EYQM(]OD_:&-1faDO=X^9:K?C9N.I-,P9#b)4=b,+Q4b9@U];PH7N
>4F.D1Z[TXPW<@T,_;<-[RO^XWd+)0PEBRPf38bZ&If\-:f@df=;g5d>bb?#8Ff:
7U-c:)+ER^:J:]4aRV?2f&;,NS4BN3BL\POH[:D.>3P<E]4S&GBC;)^CMUN:F;bd
KL&Y67Q+<8f)gb+3_FN]<)=I.V0:&@;?AD,:7Z_4WM?MM0Y5d9>3VLZJVF.7\CY(
Y-0+]3cED5M<1&<1=#cWf4ed-OL-J--dW[YR:JZ.A&A/3.JbCLFGG^JCaN;D=D2L
D5:^7eCa2.e-]2[U/XAB>eL;Z6>(?TEL(Xa4[1(UZI]P7+]UQ<3MGNG-)gceH)<V
,8df)eM+eTb?((CR^[H^+SI6^I]&QM=U_>fV]N&/_4A]T/2_1R,4#G&2+2gON?0K
CZ;7-^587O^LYX0XY5,fEF#[^O(VQZ;-VVN2I(Ue]9G7=Q9RCUaZ&B;QdFTI9L9C
0bC2BPO\fPBa/RD29F\fB7JB)G317geXJ.cJfNcd[]O0-B?NZ\U/+4+1&AOIF43C
,3gB);c:4XIX;0<62DO[,4[]N+@S,D?WN+eBK.LC&R&#]Z4T20A)\f6a7fD2G[<U
>BT?O<g0-FIZE@[,+DO/13K&gb6PRT?9c5[,9bV:7,DM.,3_U2X.\Og)^0-B[Y.#
+8>X70;?Y(+71(ZA<V\E[#5.&)/8T)U>ZPES:&N@>O4,;4EJePVI4,a7IK@NbHB2
bdWRN)/=]6HO5gT26IVT,\&-02B3UGF(S-J3MdP26-)K,3KbJ\\;S>fA_bWR_Q42
J9\SE9_ZL[:Y-1Q]2FX\P][\KPU#+66[;#@VH9=Y-,+-QTfM@^aQ=@US\f#c;Q<e
AL,Y3P)/98d>\Q9\:VBC&Yb?4D/SF.=3,T(A_M85-_4<X9,/O,LI\MFI3>IX5La\
DP6(-5I]W(Ze1g5e^Y+XB;KdN+R]/LB_SR>5KeV<fI666I5UNWf,032V>99EC;^5
DgQ;M>QRSY@W\H0Fb(a3Q/OB+^YGR#>^SRAb;]R7dJ\0/09&VBU[N7<TJYZO&(ET
3eZ>K2OeQ57742BQ4YQAbE>+=L79ZD):(@K6>5&)BNeCgWZQ64\@:dMC?aeE8<):
R,1L.R9JP>4+Q.LQXe@(78&+IdQFX1].O#@[XCEXfYJV02AAKPUK^.a;4JeLJZOJ
7ZSM9;8=\0+CK53-gW2J4?,.gCe@=\Y;D@cLA?)b<J7B_R7Y311FB<dOTC_b(fA?
GQAM:aNT+?=?BDM(LUS+?,6E)&X;A?IW9<&M3HeIBBU&Wf&;&SVN</67Y7)W8gNH
D#]>K=A_a.I>]HDYD;_@?LX?82]VINK<=GN>eGO)80.QC,W4/#Y&;W1UR<G#.G<T
ZMe0IOa]MW3gEE7D&Z-W6dL_?+^5&5.\UZN_HB5W94cW0FZ2=>c#-bLOKKf]<S98
,b4Z:T50fIeUQ4OaMUfPAJ;>N#W\\L,g:/<DSF:aUBBPH5:EHPgJ+M3L@M@\1&gK
GK1LV0]M5]&7/9T1DNT#H=-_K.;+U=,V?\1=.NUHATXX0/D14^&)Z;9#OO;Q5gXB
9TbHFLD+NV/a63[H>GL,gcW7HL2GfIFIAIH]VdXT0KGXZ4M:fMPb:.R[@UY?&](D
&/7<(RT7K83CBCTLGY;1Q[]^LIeZGPOfcKM-@MA(/LZ5-0Q51=9>+4>X)UK)VaeQ
a2WLYW[ULW8S4Q;g(2[#C[_^Tg2O]FeJ_Rf98_+U6g\PS\\ME+ad>041G#X.X_@M
Ue-;3]Z/8Zd:=6_NX2#Q?gB+AQE3XR.E(d,[b#U/eDPB_\@F9+46(MO<9)>^cR?I
d-aZ,N_&-J1KUK=JT3B=UV@ZR=)Q3@#IY0CO2MX>=1V@DU<DMS1CAY\5^2T3J(1[
3FZ::5M-TDAUJ60JBQ?fWR[90R8&=;c>NBU/X13.;]eeD;L@Z=;Z4C8Z8d3-01;5
:(#X>XVMBX&QE9&P?2d0)2aCeO)-4IR=_8GbE4N>CT@:cg#4EBLg/ONQ5MURO0\R
&^dRVSR(N/LA=Pg&RI#9e)GL&MCO\&V7X3g@ZP,-L@?+fLFA[7(,QXOU;;]QBeG4
7_]FV,PH]_M]@7c<e[IO9MW<\=Kd[W8PfLX2[1E-&.=0:<:OV#Z/BQTfe4T6Z.4e
3B9=3@__e]aRS<(HO;5+?fOWGN8&)[U,?_EXBTfS@<V]e:b+(R[R9]Sd/G4K;2\?
;aQLJ2,P@.:DFZgM@72421@9aa/gNK/+BQ>QZI#OU^f3E5>TBNNHE8:K&[_@GeJ=
7PAS8-+<9f+B_J_[=V#/_+Y_VW)Yg6aG=,>8.0Xg4((?\F)KdMeMEI/HJ<4[3BFE
Q:bX)SD3#6+FV4\1N_FLFaXM=44R3bH;3Q#gRM\<:HcG8>XAMW-E0MYYb2E5&dQg
P-bO4;(M/O_KS/BET@YDN]M\G7R4+(V]?E1d5<9)IKU-AFGA+@\4X7aXR>@2T_-8
7f&:VfN<2G#O:8R07;0/4JI1cb=/8gFFI604G^dJWH<AJI@gc\[g>If>GYD?]8^B
I-[AKQcFPLYYR;:<3G.3<1+WN_<WIG5D.TU+^bRD-1&00VCV/M,NU\O1f+Gf==Y\
A=Q=+2/4Tg4R-4D15d0?O034CUaQSf6EDFXB<Y=;B;VGCZCeT2VaUSV52:K4.C..
N\<f()F3(\[V,S?R;V;2R0gCEB5KYaWLFaXLAG5(#IOZ1C,U29/aYVf0K#<0f+:_
0&]G8,5[a>=-SOSL=O\_V4]-8&@T<7Y:Pe6>6LW3B6S<Ra8@)JDIYF>I:NI5<bEG
N3,[7c>&^\1cDZV.Z?5OQ?FB((WD_H>?I92?]@CJ+Od1;WGf-0N^@C-DHc1F[?+V
Ca8Q=Eb/JU[8CVef2_O?\&E:UV_S[&7T]CD)J[L0^_3-#LPNZNE1g0EeXd-@,B4R
I1gEgg]gf@?,7SY0D,fKa+_e0L-L[c_T\-)BCJ@9J5E]c^BKH8I+<>)7?+;b(,d>
?cTcb;c&D-]ZfT67Nc3g[\N>?8A\OC(K+WbWL9.dSCW(\)B:5a=FF1^5OR:4,K;0
d[PF)ZfR7RMV871bda1bRQ^XAagbC;CTEE/)].K.H/>Ze14&-b@IgDULAKU9K1O9
bY24^6_YfFO)_;AK;<-<W0(e7e+\]0F\54_Z=[)b;VBH_,S+CDbGEG;QO];K;SMD
=4B0SR2BeFd(:VN@8eCb+(e8<4H\a3JW1NAZ;X>32=OZ_-B&HND5<=bMOfT,1C#2
1..^JaT.-EW(0$
`endprotected

endclass

`protected
Ud?Jg2IJ^O2=gF569P>b51;)XJB-4H8;]/:G>WT1REN9M_g?[4,T6)dM4SKc6MT5
>IR-S;TE[FK)D=(-Sb\GX17ER#SbaKZbL6BVXdZW7)eEAa7(e)]Y^D7-Z5Kg@ALI
.^L#LJMU[8]ON[KGW\-[^,&J<>XUN-I)>>9K?;432@?&_+?SLK5/H0&@D8cHDS^Y
X<F6d^@N@4[cO)??SR0Z9f&3MKA][.dfMbdM9WAS?LeVBbIM6))1F[]AeD7,c;fS
5=.d:N>#eI#Ue+<FZ2WH>PRNT0KW2bVW:Pc/,8Xb]Le<a3^?-FZH64FY2JT_40.R
LEK>g\Yf#SA<fW<?<=B7<&?1AC-bJN8C2J@K-8Q49c]Mg(gWd)2c;3U9AXRGdG9T
($
`endprotected


`endif // GUARD_SVT_AHB_MASTER_MONITOR_CALLBACK_UVM_SV
