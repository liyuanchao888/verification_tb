
`ifndef GUARD_SVT_APB_CHECKER_SV
`define GUARD_SVT_APB_CHECKER_SV

/**
 * Class declaration of each of the error check stats instances using the
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 *
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */
//vcs_lic_vip_protect
  `protected
L8N>9Kb;<#J40YWAU#(,0>]3LBZ<#\TD=5fBbPP77Xe4;U55<c3L5(RRZCKQ1G#G
@=:ABcc0](I]C7(>.gZ.UA?Qa1>5)K:J52SdO52FDGUR[FV\+EY1KOSX02[8aB^)
V@dXEce@d_)U#Bc@KXa&_Q>S]&,-59ZZEV7I3YZgf.R+R&e\ZF/e(Z9:,SFUZ6_M
6c4WQFc6IK]48RQ,RUY\&<CE]a];dDeN4^W(\2WF98+&W+CJDeD0=[NINYGe@Q<;
-QISLKKG88a-88\E4\dA#0\=9?UD1PFc>DSF+Sf=Z7\T)d&;A^:&;ZPdeeRGQ,\Q
V7;TB/.]U14R4[2Ucc>,K6RX/DDEE/0(P6aYD[9CFX_IL,#Y#f^c+gdgZMAP<[g\
A^OGcOJ1\=0P9AV#+4[@#-@T./IK^^-AgFa6=LdP.:<fR8&Cdf#.e_7_3@9WKD)f
;_88Y4YbRBb2YW_K6F2:f>XQ3^d75d#(?D_8DfG3gc@F/PJda;Ad9+QdEA4MRO->
3Z;H./E>&HU#&2SQQdG2dT9?EIJ3[RB(C^6=B:C-+T4O4-S/F4UM]]FMX=(&;C>,
g81X8PU616_,O&&D2f/KPcR/_^fAP7FS)c7G9,ME:c6;2gc^NPC6-Y(b644L@=99
C,Q9KF7\TNTMV70(_,TH7OY1+2:(E(WDJ.P2FVF4<P2b9.b5@ga9TXGDV),BUdMS
YfgFZ&<4O.cZ3UK?L9Xe5H=N?\X0\RO2>]PLF>04Rd]3(]Jb6-P1H5U-bLdW0Z3=
JU9eXI_)IN@@AbG73TLYM>GWO]AbXPS-NWIO<VWORW0@OK<O#K#0@\dSA2;HY1bf
\]#@51,[K)5RA(Z85__9#K8ZW5S0)O44>]N1\C/?I?[P1PCL=]C9fN<+<2JO0X-I
0(=PLO4I6OUL?XB3@:]NfHR.BdB58NEYf?\9;+F5/T@_(TZY/O-<4GaP<TGKTQfI
DaR]SZVRW7?<M^G?6a][c<4]V18fOI^K6F=F=OA1U9g6=_MSa?&X_2HTR7,I;RUU
A7QM94:Kd<MPGCI0e.I;^-5c^I7&IfJ\Y2eBV;)5^/&f1M(YPYZW3I34dC@&E#4A
gLDUW]K\O-JR+:V]F?TMJ]QG25X9HbdaE])0HfObI955b4+5T^(R^./VW8a]W\eA
g9X/bYA31=I,^S+EO[54N5NA>YEZM]X<OQZ^?+E-(fX\/><U0e9[T;8.6RQ?64X-
4AQB6gS4&8fgCK1Q6]7(=]_[.b^^<_La.c:EV4TBZENKFA_A^2Ud2)00B8>SEeHd
E2[VZg9?@U[&g];ZcDTWZL+c=UD+?K[O2#+V/,Yg4)7PQ+cEMLU3/>@96F1<=#<4
K^1cL<ZMHD.Zf:_EN,9S&[:^)B<>V<EX1:\J=.3_A(&ULQSY52Ac41&E>:+9XBPM
=@c<S(&<egBaOSQg=PP;Fd;JH0c1TVRDNG.b^)9[D<7M]>9Q/>?UWfX&MJH[[>g_
=;bO\ZQUJHa;S=HM+4E\)fV0E:794)4KB,3V=b5[(QI9dYJ;AI+^.U.G#2H:PTc&
AI>Q3D75Q&A9878D[.,.QJHHY-dbf+16UBS+.a1O0Q58&]GgCK9B:?LcQUJ=U+:F
/YVK-gdK>):c8e;X-A5,]PV-H)M,R_9P^)^HBaeW1.Y^H:4[&8Tf0IYZN3[F/6C/
M[7]),ZLEM8R1.S/>-7AAO?(gYfVML(N_gMDS:N3-U+\FE&,H&-GH=gD0GMb)ga=
1K7TQ>Q+?2HB(K]BfG[_WH>LXK=KC98cJ(YJ/#W<L4ZQEGV\K3e&79LgD_g18MIC
FS]3--6C<=e?Y(6PL_)SU;:EMN82T=2&V>HWMaZSa-e5HP51ZbK#A=B3C@[L.[GJ
2(,7YHB+&eY#(6XMA-7TgR4cYOPNSQ<PMW+81.Mc:6[/4T1<>],HDO22D9)N:HHE
,1#eF-Ke0egFAN<11S_WGSQRMP.,CdW&a^.[PK/]Ba=IY&;=C/U/S?-bH_24;O<.
/YS/e>NHA&+W+7;^WZ@6=TF?[0+WA>eHZgO#<)W45aOTM_N\aA?1YM/+X=f4N,A)
/EFPeY41V[Q])O6NE815<I^BY.-3IS_\5D9cM;SJWHg63[Ce5<dCT6PbE)\0?A>W
=.OHE-[.C;@QE@f@CC:X^64TZ1[JSaa#[<W95CcGEcLUDa\#U;V)=EfV3dP[01=H
<eE782F]OU234DJ:BK_9V,B,IDRaDKE9BGV-6/Y-g3_DLEF<^3V#>^,c>/AbePZX
dYcM\QKU@Z,cOJSIJ&#.D&?FaW]1P?>8E?>^2KJ2#,3A66Ac/JK^@-?EGJ1[1TED
JK1+8OY#A#XX154LRaWec2)L,8^XPE63fbN>IKa>Ta@M68ZSb:@SLR^+X8.79Nea
)JR)7fBR,F3KAW(0_@+UBA_CC=8d.74&&0UK+ZGaB.&/08aV7/U=2E2PUC-2eQ?f
Kd7<<?D^45KB]QFMffF#V3f2X(g_+\F#NCgedF)[0IL78b,G&T=:9.[)>QOS)RDP
4a4gNZ#NC1cJPeSPT=W45E_INbICde2AM=RJ]49.=I4(-EOb/Fc8&C[5cM=(6V)9
\AfNVWCFS:BUVJL:\C:b2[K5]AUIIS?396DUOBE\RJ99fc.,b[24L8D^OA_;HWTV
<.7V4YIT&e4L/b@fCEHRdH131H0](],?^?EB_WKM/RF7X8J3IeAXe++EN?W2+503
8Q/:K(ORMOH0UQLY)4YG5+(B:bU9T>a09U78T-a_LJ]HC_.)1XN<_0C>O;9+U^&,
.+C#79]@.R,(CRS3=,egVM9@?d6BU,d+#EL+BMgd0>7B\O(L9Y0+LE>bK-d(gD,2
+R(gWZUfO4KAUZ.TR,L+FF9@1$
`endprotected


class svt_apb_checker extends svt_err_check;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************
 
   
  /** Checks that PREADY signal is asserted by slave within timeout period
   * slave_pready_timeout 
   * Group: APB3
   * Default severity: ERROR
   */
  svt_err_check_stats pready_timeout_check;
 
  /** Checks that penable is asserted one cycle after psel
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats penable_after_psel;

//--------------------------------------------------------------
 /** Checks that pstrb is low for READ transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */ 
  svt_err_check_stats pstrb_low_for_read;
  
//--------------------------------------------------------------
 /** Checks that after reset deaasertion, APB Bus is in either IDLE or SETUP State.
   * This check will fire if APB BUS is in ACCESS State after reset deassertion
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats initial_bus_state_after_reset;

//--------------------------------------------------------------
  /** Checks that following APB control signals do not change during IDLE state:
    * - PADDR
    * - PWRITE
    * - PSTRB (when svt_apb_system_configuration::apb4_enable is set to 1)
    * - PPROT (when svt_apb_system_configuration::apb4_enable is set to 1)
    * - PWDATA
    * .
    * Group: APB3
    * Default severity: WARNING
    * Note that this check is performed by passive Master when 
    * PSEL[svt_apb_system_configuration::num_slaves-1:0] is 0.
   */
  svt_err_check_stats control_signals_changed_during_idle_check;

 //--------------------------------------------------------------
 /** Checks if psel changed value during transfer
   * 
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats psel_changed_during_transfer;

  /** Checks if paddr changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats paddr_changed_during_transfer;

  /** Checks if pwrite changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats pwrite_changed_during_transfer;

  /** Checks if pwdata changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats pwdata_changed_during_transfer;

  /** Checks if pstrb changed value during transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */
  svt_err_check_stats pstrb_changed_during_transfer;

  /** Checks if pprot changed value during transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */
  svt_err_check_stats pprot_changed_during_transfer;

  /** Checks if multiple select signals asserted during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats multiple_select_signals_active_during_transfer;

  /** Checks that bus remains in ENABLE state for one clock cycle in APB2
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats bus_in_enable_state_for_one_clock;
//--------------------------------------------------------------
  /** Checks that if illegal state transition occured from idle to access
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats idle_to_access;

  /** Checks that if illegal state transition occured from setup to idle
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats setup_to_idle;

  /** Checks that if illegal state transition occured from access to access in APB2. In APB3 state
   * transition from access to access is valid transition.
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats access_to_access;

  /** Checks that if illegal state transition occured from setup to setup
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats setup_to_setup;

  /** Checks that PSEL is not X or Z   */
  svt_err_check_stats signal_valid_psel_check;

  /** Checks that PADDR is not X or Z   */
  svt_err_check_stats signal_valid_paddr_check;

  /** Checks that PWRITE is not X or Z   */
  svt_err_check_stats signal_valid_pwrite_check;

  /** Checks that PENABLE is not X or Z   */
  svt_err_check_stats signal_valid_penable_check;

 /** Checks that PWDATA is not X or Z   */
  svt_err_check_stats signal_valid_pwdata_check;

  /** Checks that PRDATA is not X or Z   */
  svt_err_check_stats signal_valid_prdata_check;

  /** Checks that PREADY is not X or Z   */
  svt_err_check_stats signal_valid_pready_check;

  /** Checks that PSLVERR is not X or Z   */
  svt_err_check_stats signal_valid_pslverr_check;

  /** Checks that PSTRB is not X or Z   */
  svt_err_check_stats signal_valid_pstrb_check;

  /** Checks that PPROT is not X or Z   */
  svt_err_check_stats signal_valid_pprot_check;

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
/** @cond PRIVATE */
  local svt_apb_system_configuration cfg;

  /** Instance name */
  local string inst_name;

  /** String used in macros */
  local string macro_str = "";
/** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   *
   * @param name Checker name
   *
   * @param cfg Required argument used to set (copy data into) cfg.
   */
    extern function new (string name, svt_apb_system_configuration cfg);
`else
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   *
   * @param name Checker name
   *
   * @param cfg Required argument used to set (copy data into) cfg.
   */
  extern function new (string name, svt_apb_system_configuration cfg);
 `endif

  extern function void perform_read_signal_level_checks(
                                                         ref logic[`SVT_APB_MAX_DATA_WIDTH-1:0]  observed_prdata,
                                                         ref logic                             observed_pready,
                                                         ref logic                             observed_pslverr,
                                                         ref logic[`SVT_APB_MAX_NUM_SLAVES-1:0]       observed_psel,
                                                         ref logic[`SVT_APB_MAX_ADDR_WIDTH-1:0]          observed_paddr,
                                                         ref logic                                    observed_pwrite,
                                                         ref logic                                    observed_penable,
                                                         ref logic [((`SVT_APB_MAX_DATA_WIDTH/8)-1):0]  observed_pstrb,
                                                         ref logic [2:0]                              observed_pprot,
                                                         output bit is_prdata_valid,
                                                         output bit is_pready_valid,
                                                         output bit is_pslverr_valid,
                                                         output bit is_psel_valid,
                                                         output bit is_paddr_valid,
                                                         output bit is_pwrite_valid,
                                                         output bit is_penable_valid,
                                                         output bit is_pstrb_valid,
                                                         output bit is_pprot_valid
                                                       );

  extern function void perform_write_signal_level_checks(
                                                          ref logic[`SVT_APB_MAX_NUM_SLAVES-1:0]       observed_psel,
                                                          ref logic[`SVT_APB_MAX_ADDR_WIDTH-1:0]          observed_paddr,
                                                          ref logic                                    observed_pwrite,
                                                          ref logic                                    observed_penable,
                                                          ref logic                                    observed_pready,
                                                          ref logic                                    observed_pslverr,
                                                          ref logic[`SVT_APB_MAX_DATA_WIDTH-1:0]         observed_pwdata,
                                                          ref logic [((`SVT_APB_MAX_DATA_WIDTH/8)-1):0]  observed_pstrb,
                                                          ref logic [2:0]                              observed_pprot,
                                                          output bit is_psel_valid,
                                                          output bit is_paddr_valid,
                                                          output bit is_pwrite_valid,
                                                          output bit is_penable_valid,
                                                          output bit is_pready_valid,
                                                          output bit is_pslverr_valid,
                                                          output bit is_pwdata_valid,
                                                          output bit is_pstrb_valid,
                                                          output bit is_pprot_valid
                                                        );
endclass

//----------------------------------------------------------------

`protected
aSNQabD]QgVaLZbJZ(R/bZONMcGH;^J2EGdT(0DLZMS9e?]];f=]+)3-g23VZ9e>
Y-C:D>U@#b1)^9IDZ;^6Z2@47\dK5gf,dV.Ng2_UY-a\fY/+0_a5N(-bAd,:O\BA
D6>POD].8Q<U??N0OVWC<)(_f3RUB?>I_)eY(Y+,5:d:c#aaG@H0DV-6S?O4>deZ
/:.69dM@])A<FOe3&XMd30KFPg46&;D4/1-:Vb?0gGA/42DC[@@:eQAU\XA4[7A+
2T+O3KL4MQDCMAe>1JdNJNS,L#2NgXUFNJ7]b<4M_aV2D8K2#K@AV^7#g2::8J&c
]f&&F&/SWB,GI))dQ(-(/Eg106dCTTEY[e0B2X3ZWFKL7:.V[1;WYA\d/.JSSGSQ
1&)NcBE@@>7SNH)(@:[NXg[^5JWS)U9c4^68/U6G3[+?;#gM)ODb;WfQ,bV@dgZ&
LUN\H+,g@6./H_<M\1aUXR;Q^&M/eNV+BV[P8eML-XGg3ETYR2X@_/><TD+VR^1M
_4+O#NKfe/G^=6F,(9D4c9;JC(=TU]8NLWa(G<S#7?-\&[f_,[UH?+E6cW?Hd;K:
=WaDXe<#I,;U,P4H46Pc9/=UBDNZ#(>?/>+ILR=V])V>-SBU/0#&-P;0>#g;2XE-
R-f3J]3F9F+Z3J^gWOGB6;6KRLF,N+?^TTOVL:bSg-P?9)Ndc(;;F\TX]2Ef,=2H
MaR35]F&K\b5S-C/D@;ZXLFKYJS=80)=]>>f43_G0,(7=G\gb/26OWJZJW5=(N7S
8UZ@W_(KGL<3H84ZW=3VLe,TCB;<,-7[=PgX?]P:g?VN<<^JfX#c3@TY-ee7QSVN
U(^ff#39XOVO[^1:CY:#J3K[[0@VgLOB?<(&G@0-#A;,0L(Pb0QTA>EeFG>F9WbC
5AS](eL+Fa#0VMWBO]3O&bCedP6Pg]:H6+0QMXK7E[6SERbFA@B/\T4S3).60/(W
<B<^QG-eQeL=S;M6Z6.Rd#+dD@8:Y_I_A\E9C67KH7fR[>YU,F33;ZSH2E\T,HDP
bWMKG.?\FdeNBOHW@#_=Z1>)C;5+0U47AV5b0@e?;Ycc):N_#J[a]O_fYP^^F]c_
;>J2=;KC.I(O&<:T]OgES6L1c6c?J7\_6^K=BFRIHIfWT3DCFOJ\K#)f\)b0R<EJ
dUI=O4L>Le-)\6+AH41=dPV-9U.40S54.)P0;G:H#D1ePbB[JHG]1d\/P3H:1<(E
U-^eVD57P[^<5@TRC75G0QZ6,1GOQ/(MFf^@X(CVIS)dd/3NM_:W[S/P0)YRERT\
\IT88+DT]G2SP:-7BH+=R.dZ(U/,,9B3KT<RZ]1/GB0SEf>^IffXWGcVdJC5KTID
5-2e6AK\P6_bW-)?Q:-.CB9@;K:G.HJ<,K8GN#:X3&BAKVe=d,+JGbYXeWTJ&IYW
]V\8DL#(EXN6a\+b7;LRZKc7adRcP?PW^-=W<P_+U3,d+4Zb?-&BL#fcffc)##N6
4>DGZ1K-CAd@cRN>?d_Y\J+N(D(GWQHSZ#S8RT?L7F/GWQOI6a5PN14f9;]XH8(W
+OTY@0<,fZB^EK2CH^5?bMK8fS)+\;-66ST_[283c>RDF2da6,)]Ya,57II(>>3e
#GM_;fEcA8,F4#(PYUUXL=^1R\4.R3c3aQUdWA2aBPB810@),Zb[U^;;EV34DfZe
[-0KDVU>5^-dFVgAeS&+#>bW,R^JZAH\Q<6U,9:-B.L0g47#8cQd(<,C\@c1[EI^
^OLI4]L;N]ba.--McPg?56\IcAH)9_HS0&>(M@3M)7L_N?,/cTHVEBCNQ8?1DW8A
.aIA+(9Lbg+F&D?g<b#d)<ROgIdNX7BJfZ/97IF^N;R,\_SJ]/J7?L^26TV)T6^)
Kc-@3=,Z@2J&&WDM^GB=DK=6aC:?Q/&1Z>O;GN<2&5PfNU68@9Lc^Qb(\8360cXC
9bIZLY+(6Ye:KPT4H)JZ8K](;HOUY](8.U-\<+IC<I>Daf-deN;E5a0e6UCZY)GH
2c0T@.G9LJ)2+82C2U3@BOZKJ9P=R[T:71ZVP>3HR/8+IFaN/,3XG,Ba12AOR5\?
M.FD)5^,Wf[W6TSZ@F;@#XHR-.;&(GKZVF&ed@YG[2(6_#X3^M141-Y5VR.e.TAf
0>FA3T?G^NG.aNRN10J?JY6;#H/U+:4A9SW>GXW[NWFc([)b1;Ne781N>,X<P8&b
abDV<b@-a?_+>A/1.@W6^?&&cX_0-c&BF9I:N>Ee+b/(4IS5&[13<ZI.2F7Be2(M
c#&8KT/(e[_EPO2\c;gVR,H>A1+>A-X4d)7Va0#Y5ANK:SQ-N@_#A;:@EH5ScKC)
[;)\R)+/7R<PF<F+V3bX(EG]H9/PV46I<)15gQf&R/+ES:A6NEGYVe180&2UGDP&
#Mb(\JK#_&=2B:Q(CZSD6<5KFcG:P]B8c#^=VTe0J>N68]FC[PF+7b4>Y5I-;TM]
ITfbEVV2dLf2gV>ZB8T@#(S.eI2^K2f+YGI9WP[221>GWaS/Va7e6I@IT^],2:+@
&,)e\=G6=]+9Ma/Ha40AE:6dS(#0Wa2==GQ]NV:WTY6D43L614Id>YF>TH:OYW9,
Ffb0Yg69W7>-594b=AG^eF[-X?_g[7W3..I19OHL-67_6QU(8^,?=Y-EbG[Z?3L:
CPA];+1@E\dW,GVR+=:d)Y+VORg?/@W#VUG;D?QIg6d;:G;_/;A1dg0dg#VR)C41
NEN-a3Pb7EP941E&IA8>VU6:UGSO&Y3O.MG@RRVMN/[ZMF2?b^-?E3Q9Wg[QU:>4
:#R>6#@#,_<IgLU:H0WIO23bWH)BG(MB>P46HIbC]4BX:\N?7d,1S:Y&]/+&d^J4
>Sa7D5f&^Qf<,HOEdY/K#?R9-c&cSbL;dJKgeW1F1/\NJE6+5[RRAB3L6a;Q#54^
AfEKRJ+?=87&\YR3Z2G)3SPX,6\&H0;P5>f^BT()f?QedH4,OGL)2Q.:WA:>8AIO
5>Q7?\c[+W<YAEL#N0e(=?Fdg.G&_D04BBLe\;\.;,HAfC23[BF-V[b=#Ae:bF>^
G-d^fL:F?FC)KGdFaUbX^TD&^==IZ1D/CGLH<LD]B-3I1.=DJB0=U+@)K^aBM0=B
[eU(#4_L1RgF;J;]:385#Y9[B_V0BeSgAP?e\_+,(F[M)bVZJcJ5fb\@R,=f#EUE
-K[[Uf=EV7WcXSXK5Eae@-0aKRcHXfZQ807H5L]XIS((.B+1)6&8PUeEUZ?X_N+4
)51NL1K-[-69,>JFc@YZSV/_F&Rab@6<O;-588Z-ZL;BbXc[I4K.?\1Le22b&Y>6
-bQA7Y=RCXLQC+bC](<b5?IAV?P-gIE1F_4XW=B62V^HJ2D2SBf5W#9_Z)7E#4)2
;17D/[D@^SI<&]V4fR.a?XMdA8FEV,>VP72_GXY7:gB\/EdHMcITQKCSVY5Y6=@W
_d7E1OV#&8?T5JD.YD&=3(F0g/Qg)?XG[fL96#A;U2F;HJ3SR]aea)_^V=@VO;C4
2Qf##K_g^:F91Xf?F?54NCJ)E9d7>\;ZFUA?Q@P=)_[DW6H+I0cUX3M85WL880KC
)/N?d>.:QCb4VVV:Ba#RP]6P5BX=9Tfg@YNT37JcDU&0H=\BZ9^Cf?#@HKgb.&e3
<H.DZ3^73>)MG7a>HH.^e7UPEBOQ>f)U^-J?T-O?\78Mf+O\H,4GM;;60B(Y4&>Z
02D##E1^^YN-&+ZA(0eM,-dgO.Y]c_782^7bdc[2X[fPdDVd<24P]]V\X?Dc4,.;
_Mc:W?1FP6SQV;Y=^^L:^\.<IA=SC6#5/XNe.aWQDDM7OQD=I?U5R&d6I0)F[+AN
WcRXf9.4-VF#<f#UF7@WT&W_9D^&@096^Kd\T.(]?DLfF>/QM)>f]UNdGS[K9-NS
9G:93Ib3<A<14,IU)1V:1(BcYU:S+E(JFX62\]:dYT=,-2=RZR9#);8&AcT9)dTO
<gNX7?8PQV?9D^/IP4GG]T7O;3(9>J4B-(D06U^^WYQ86gF^?=#Fd8gG.fKLQ]#b
ZWf8UIRDFV,dS]_\C/@e^TFT^.ddI;gNOL:9NKD<_Ng>SbL3EGXd0>DC#UT?JYFb
WQX4UG+\?b?D#2\>X<HH&OX.e/8Qc@XQ4._=^9fLf6E/?Xb0FYB>&f<\59Yc7<>G
?eg\.FdRSCBMNO-?0e1<^=FTA2KLQ1HVL.HH_C4c>ROce?bH]<P@Z#I?^7Zg?I[L
P9H57@T=>4S>K15eR7.]=NfT3IG;EMRR/gZ>&ANXcZ5aM9=RSOCgMBc;U_dH:c1L
2Ud&&3F3X8G7Q[7UNLgZ=Wa2Hc+Q?@,.-^IN@Le[R(@G;[S?\3N67@MB+D[1Qa=A
dIZJ/V;?f\Y3JY+dC5>Md=Y-f]MDFY[6O389Q2Q\)K;087HH]T;G3)/E]7B?T#5.
O&?e[M8+TWF=GYGRQf&EcGKHM#[7CGf=CY+VR:KVU?_K-aA0E5/I8LCdY2+(P+Na
gfgTN7gXN::<FXcM_;6=1:2;_AM_7.EZZK&S(e1d6?5cb(U&e#=)L6@C>QW..6Ea
1=]e<;Jf(<5VP9BUG\VH0c><9bC5O]gHBGS5T;-\]@2V?d/_NI:f.JT28U9S;&44
-e)>2(=#R/BaK[KRJ+0TS)fM?8WWSa<BE6QA]68;_c(X]PZ_V5,3.XfEM81(XZN8
K&;[XD6_b.Q<8RF.=<7MDMV88VJMa3P]9eBWHg;O+FSJ>;7#[Wc8GLcb-O+?54;<
84eF;cAU]&QA1Z)dPV53Te2c?9@8ZA-6OA+ND.QIHRdBF(c=49S?>S#?]@:#H2N3
.)^[fgU\/@\6WX/?,+OOX08dKUe<_INXY0R=]0F(-^U\D(ZfM.&FQ9g5gNcQ;L7J
8]PK>G&C,]MW,8P?4SCH?&?+Ng8)/.>FcGO=_(WVe-7FF]NNYWNLaa9+MCT5+;MJ
3Te,DFC:B.X/<+B&f:d\1R5UPFc@T3L:QFB[RRG(&C6WdD6YH3bGYK-/O-eR/0NJ
4(>RVgT_?D(TIVGNEBRLEMcV0;V]Wd=PJa-Y+^G4G,X]OAP,GMK34D9;RX;c,TH(
3AA-FSW(7^A]aYT/8YQ)a9I3C,PYQT;655O#&]Mf4TW)7DJ+5a8/88OJJRQf8+dN
9-J32.OcZ&B58]WIX)PS:18/VJ.Mf+U5KaC45CA=KJEZ<E]WA2TJ;&WA+F2R?^6K
d1d=@#d<&@f7+9gG7V<82N=AYZO2,W4SZ:?WcMgSLb\8NTX#+,A1=)HHY.bZ-0)3
TOJ;0H[b\X[2&^=-/\=#<_RS>a/)F]2Q(3VKG4WSY#(JH8Y0UW\\UZ]g-/aWS/O5
C[Nc846AUXd3+2bCYA?&gYU(Q,SRdU(XI+]a_B)-N\=1_M:C@XQGbK\T=R_#G+(O
.6cCeK+T)EK_dJB.YXAX-#[-[IU^eL0F_S_EAGPO>FPI3A6eZ]#\&9^6HR[.ZCK>
7V645b\(HbEW@,HIM+=VJD\DVE@5GV70<eM=MIS.,=]O0C#&HePPZCN^6g+7Q[R=
GDf91OB/>@+[g^IdK].N75Aa?ag-7UZ74X?c]KFg&<+8Y6CgFRUW-++BG-0)U#R#
a7c)<K[<e^3.8I)MGBUTQS>cFaI)?:TYOR58L9J;FE/U#K3+00#&N8MNZ+>Ue7:<
dCVgQ]+d^>KX5E\-YfW[^>H+B[&0cD.gWg6S<LC-E^Uf_BA:MBfN#5,<DeCD#KgQ
<<T9[7VEL+)>BKZNOe9,NR&UY<,&,+0KD+IIL#_HA10V<=Y(c-C:Q9ZdJCcS^91I
^d<R0TT4g4ag21EQ5AN]TK-]a+<EV#;&FH5K_<APD;;M4_<\U-,BWJRQg,Tg,/GO
ceSKMe/-YE_<)J=cM[g9@?:7f7a:F#[0IaY@@D5[L7=IDT4#\/VT57]d+TNIc(?@
VITMOeB2a.;KMA>=.1JENFO34)Ec8?4b(YfWTf=W.g?77;HZJ^3KUK7L@&2J]c_(
BGDbW)_&W<e8@&ZCO_;UMffWVDMO-aCNK?HN_GEP<<MJWRGH#bG1)(R=Ba)L\,LW
1?\[9V6XI4-UA3gH53&X/1=eU.M;g_-3OZ5T]-)<FQJIU)Y12b&5Yf5F)PU3@]&S
4ZM8?8)feY<RDe+?>_U/=,UBBX\30S1O1;Ge+;ZH&e[8:eW:<SVV7W_Qf)T3U^7c
HG+CTB7STB@1bKdO>=/d\F@H)YZNHY#&I>cB(gcf]f=QGI#fA3)HcRY.b3N8J<B@
OU,0[OZWS[3Xd/)&K-7ZW:#T?MX9?Q[-L;=W1;EbS.U-D@ZU-KUYV687YP=L_DI^
XMb^Ec0fgRHDOGa2[5Tg-K2Ng&DBJ=O86DZJB?Vb#BL&G^UfE.R^c<N7XT)N&@G\
FU(@C1e/2Sd)aB-[&Wd0]_D:MSB@TfT=G59S1@[80>Y@\dN9RJBbKf<JO>62_J/C
QXJC3Q=e;(\_K3=d_/(<eYgUHW+1cW+36eNb?1(5FfM[/0Y&U0H1SK#JG#_cL;:\
@/(^1QH:b2G(db#PS)(ACI<8B)IKA_.XAXA2\FHRKH^&EXGaC9SW_c0;a+F)AK=Z
1b[33([KNcO1cH#gAI8QN=d:M<)UTNc9AQN8gZ-WcEPeEMA/#3BcW(fAA=Q[8#3?
(.b?1W,5O/P2SE^MRZ;cYO/B8J><L[^1JS6T3+AZ,???EEc2[PDMV&]O73Y:fJ61
#0E6b7fE?c_1:B^Bf()BDE#Wa4ZJ7JYS65f3PAJSbZDN:&g\/XcT3Z#b_-YId3?K
EbIa/,D<c^E?9M:U/GNebD>V+,S4>^gSa:dWFZ7<DXCab(E^O;T/IFH/>XAR=0?O
]S-Z,(ZNP0B\+F8-/(3RCOGO59O\-.Q=@e@K,^W^aeL;@24+>HLfPOO&?]OG0[+-
P)?P+<S<:ILX)IEDD9d/SfU#=8/7^L3gA[D_@2N;VB.HE/MZ=/fNH/4=1V[+2CE6
XMMf9.476O/+QC(QabXW=aZ[H,\\HTT<AMO]_F/U)FQ\HF55NS_[_1fX6NN.Re:)
?K::?a]D,&#&I5<Nc[)_a@=KL\^5BaK7IQ-(EH\LgD-AX8d5L/Q1UD^E3;.e7f;K
]9\^TdW[43^TDf_T-2WZ]HY0_P9M7</0da_1GJ5]Z<XGRH+BV_JS&YBcVZ0.<HJT
fNL3H@Y+]12X^)<?\1-BeJT[CL<Y1?Q,5,5d\9GGC:X4WMEFA)3&<dWcCD9[MU9e
R4JIZB:98;C:99[+DGPQ+/)5[IeJHgA6SHTLX,bJ^.U>FbZMI<GDd>IG[B4[006A
JUXODb.3[+f1.62EaQHN7&6+H[1.]IE;S=51fMcK[:Gd&PKW?K,C&+J\BKZMYFL<
QXTA=dVOc&9<M&Lf;;g_VL3CIL>==6+]FN9Xe113^TMRR;./\>L(FBUfQ9cg<BNE
3TP8W(W28;31\5LCXN,W_F^]/D5VG[V-QBO@<aCd9TP?KXe7^-+H2:.7A?g7@WTW
KfL.W&,@>;<.S[U?G\H7D-)\;3BU5.#MTL;<2(M=US0LTV6Vb&W#[g9?FJAa]9_1
+2@J]]65,,HP#=0E=MUFAYc60;>5UK,U1d25S_/XM&X6XVVZM=R:a&D;WI44-/_M
6g[U6d?1Q7a=5XY;:KPD<FAg5/H\WRM2::M[6^/A&R4<LJ9+e]QK+S.Jc6K)FNBU
g=</=#R-+D0-U67G\_W2&WVF=#WTQL85MU^D+d+eI-SLa4W^6:O@^/P),P3.&5JY
@AV:Wd\R:V)Gc:28BA7@&D)-:BH>X=CgYC)45@EHNR#aOFV.,1VVf(+_3b),<MM9
>@[Q->FG>]8R(F_(3W1cF5dAPY)+O859-V_<^=<[TURfEDg3CZ+H;ZD,4WI#.C2_
.\\N+51V(Y9D7R-6LB.&=G\H,3T<S<_:bO<c2EZY=0#]]BIY/0TL.b-&PbQeN.MO
8:&2g._YD(3bFVSW=c(\?;X[\A,<UL:38NS\<N=N#OQ>..X=#1ga[bS:H=#84>#Y
,I&F;@e70VKe:XT=K_eTA6-13WKS3bY&dYO1Ze4F1IG?=g+:;e@M0dFSA_R.gP_J
gWV]3e4XEc2C#S6O-WN=54Ga8?I>L8<3/,DedXV>77[+,@0:3BgK#G&>QK15&-PO
&JS,c&DOa31)9+DCX(U+/J5GbBaZ5CX:IcUL5],KE0g3>9-\<U7C-9TSgc3?Z=L-
H-\Ge3e(g24K1[;OH>S<CWaVHa28Q2X/YGJ;d2Y.Rd\)RK&YbZ^If_O[<8(3+Hc\
-G+QMEgJaDDgQE9-GIe+EY7+TN75:&;APLFUBJ0)\9QIJF6BR06WaE7\B-Kd8EY<
eC=9MLT+MTFE83TQ/PfAB35<3PY[<XZCRI-9B[N2&8U-P9@X=):Z(58-EY,;eZJS
Te</d1521N]27L_.(FZU]L.LBJINR:NW#QX-+fZ)L/S4-LLB&fcI[LRf9[D,P3Q<
5DJ.X((]g7&9P,,C7AU1XEAaW9G.JE[.SV:g7,9-?R/?.U-&J>^5O/-/TYIKZ)1P
[db<RYQaH0d]-4GS]L05>KT=:8;;[\-B1\N-1-)O/E09U00B0Z[6eC(XJVD6FY7>
Gd(V=X6CBfPP523b4-R=REbXEEJ2@ZP3>F;_6(X\7#;K/Bg9OEM7aE^Q.#eL4#g6
J.>9XFIcFMa+XBHc(YH2:40T6+U3(_e6;$
`endprotected


//vcs_lic_vip_protect
  `protected
M90?C+7TZY(;,5:WKX#[UMT\cGE4US/>:Y:IgFJF:]1e2?J@V@16/(EG:&5?(]Z+
J8>EAZL\aaT:(afC4TeHTMD_5(A2#FMeSg7.0]\X3b;H<<VA>CV:FRT_3(INZd?Q
3>U2IM:KOY2H8T]IA36-Wa3B?ed8:d/fKIF#9PG/7\O254N4>E\ZZD8dBI)K&1;9
8^8\WGN77NB@)FWN5I;VeYT-QFIN8:U3bg[46CPd[U]<M\JUg_Te7OUX-NZWPT?g
cGJc9b=IR<^7WW54EaTUg0@6]eOADZ>P\8<g,]B-81feXR0PJ;]d\VCYYd&<G?J>
#UUQC,+2Q_[57>e91,5g.<@3DMgdL79eJ/<,FJX,Q)\W]f#NCg:Af/]:6(b;_Y8I
YX,7A\U/aDV6bO.Z4#<WE1NEg9B&^]0]Z[SO\(T12H8FQ1NT.#/AdUC/,d2\5P6(
-XZ^:Z.,9?F\1cDAf2eCdHA[6AX<=LL&AU&V_GY,eW.HB\F^M[b>NQ[+-3FU9+-P
]2A7\a0I0QK&Q#15Y=e:S4ZW42Q&X+1?02STWTa7LNFHOG0C(L,U8Y_=Ic9Zd86<
.?_P/06EUX(3afTEDG+b-4eU)3UZK/5ASB@@f@Bf-,J9X^f@XMcOO?KY;/48Wg\V
.KH/daWXMI_NeXb;&aM1Ie5_Z=//KI><T-A<6LReLa:HG]@Y7Y7Gf\g+UCMM4b^U
:T9Ec0+\4J/4V)@III3>3U)H8fCSHU((>TJdaC50F-dOTbW.-VgD7)[X>]OPa&Va
^YY]5@87NVFZOYI&:\+CAP39Ne1W6>HS@/6.)EY#1#[VX66ZRLf/R61WLPDV79]5
_56c#2;BC&Y:fgFdPG184MCS5Q/]/-RO?H5a#9MOHPHUWW_IIRReSg-<J96U.3WP
_UJad_NOf>+XU,#FR7eA[=NP]BZ>FUVE?C88SAfA@\TNEC@<=?-@]+@^e.PebSTf
1P4:Od#:V8Q^C:<R>B)1a66>[S7VE[BfeF:\<LOB58DS5^,>O#aO7;/\#R#7Q&I(
D\<3N5+b]PX;bH]R.g[^\.-FW_e:@=,#_?8,0NMMR&QS3VE1L\@31;:?UO@:R<1B
+\Z#M-N2EOU>?GfPN=>#3dWACa29O3FM3bXT9Xe@9)WH_K;=E[YXL?\,OFOLDIO@
/4=2FWZ-dYR>48B>#c;B_<#:)04S;g@#[VPZ)E[MI#Zdg879^[RHLd\([a+9POA8
=^)X+.IJECF0H@(^[S]-G/V&d?P^)G:52OPFKDO_fYe-c6_#@A^6J6M=XcS347+_
MW/3GPDJ>U6,A5)#d(Hdb@3[ZE,KPSQ\IB:]##Z:.S3[,KS_GS,/&C3I\:=d(A+a
Ia?KA2c^2GHW-DOW=W6c1J/4>HgR\&a76Y6eI+&dMJUR6GU.8)DQ-=g0T]b4Ie+1
;F+0+KV\<bAMAT;Q=LVC@f;.ZWWHB[4/3@6JD]fCKG>gg;(_P8Z@JT7&=F51f_@-
F:,d)fg5aK==\c9J4Y#YCLf9G,6R[(O69QT\]g#g0#1,bc-+9-d(+4[41R):GI;A
,99g#LGd\:.S<:7SUdF@8LSe5J]9TM91c7F(7,-;KC>d?@2?75;72aFP_.4:#(8A
Z+X^3JCW\)VT.C:-=14WX5[gW0S?_56CJ^H7eV12[?K=__V(4//S=F+\^WE;N3&d
7C0FW:(2_K:F1EeXKP36DDEI_>&@Sdd[N&Xg:I@[(J;U4.T=8+SO6A^NUG]CP1/X
.]B7FA8=:]7+J.4W;VUHTd[<cR0b_E,)gMaH9MM<\BV]TTf.51GZ.bQKfc:9[/LQ
gF7T=VdMNaS^LG7BLfS;f6RZ.ZH0[>GR_;RP7@(9-.5H4b:gZ[^<2UPd)QXR4.G[
=X564]@CQa&2WY/>-5A8X__^9A_[?N>WJX#?-C8<>U?eEG:HbHPfHb,cf?PQMc&8
8UCLQK71f1Pb4PC,,c2,5><a:FKJ+4Qf\@eGCE5J#af-G@Y&/U6GR]UC&AH+TNI/
WaTPYDdTa;BI-><eZLc\@b/<I7OTBaL#2Le-eN-;[4baSMc[>dVS8JgD,]8[AHI3
D)HGE]631Qfbb6GfeV2:@b<VC:2=\Y>A@EEJ<aa_41WN&fIJZe@0OabGcE&LV;bf
JEDgL0]YIQSC]JC&0?[FD(B8/4H.\-Z3DK,G2Ka[O:#6/@3X:PI1M[S_ZP)+1UYA
0:I==Y>-M\K2H8bBK=K7g;0Q2<\ebU^9ZMY;O8K<g]Z8LPOfVW&]MR(S[4E+@_JX
(IAGF44,8dZ_b-#C52R;f88HC+VCbKV_WU#&fFH;1VN;U<K);CGL?Qf2KQIS.NOK
;Qc8G/g/-;^Sb66dK4;R4AA;]<X8P;+Le@^D:=[YR<.#JEXFXU?;)+J0_P.GC7=R
EU0JO^9VQF+B,GWZLg<b)6.Z\H)2e:Lg_BbT7bcddHTG?\#,eEc(89fPT&:U,;JB
.b/SHX<0T]U@>3?O];KP6,H=W,OC=VJ5DZ3e43U+f0D68IQ&+)TWc]8WGf2(#MSQ
WUFC\Z9dbI3e,P(EaM]<9<P?CB#VQVH]7<H]\3)IP/<b^ID?)f,+8.[DAG=3P7XQ
F?J3b8)8a@IN6R<YS@5R?+KRYQ-[.4DF@?49X?AcGC[4:_)-144+,ZL&&&FRB?3@
S50>J>9[/\-NZM3+;#^,N_I1Qa@;94?F9Pa>WA7gIONO:egH<5\bOM9bR2YdcDe.
X7@+5JgK\e7g1^Wc;g+[]W:G@)QX#fHMMaYWVb&]O@/V6b4bK?7e9(8GZ4T]dPUK
()P-a_Y.5AF3eRE3KaDB3WC?g__UEVLg1Z;V?8YBL:XTdMc;+9])ffSKRQJ(WMP3
;Q,W_8>aU7WQa1(PE.9XLE^)Yf&7A>O:;SO1IJF97c5V+<<6(\B1^(b/gZ8&5]?O
WCI4ZQ];X;A;=LUJG755@X8:-K+c^F\Q6MR?Z-_gZN0e)aFO+Td.Hc]@+]/=80?e
ALc+QH=6WI0.fTCaM=AJgUf.IASc_JbB[_8^QZK4#\TYF)aO>BUH<,_Ag8+O+NFE
S[9aQOL@>G:ZXXf=5>,;QK2#AKO5^X8P,2L,W&F7Q#/LE3MRHbR^Z(^?--_,TcR<
&A3X8DWX(PQ>3;(Q;gV+P\FL]\4\EM5B])3&B0e&c:;A_6[J\fXI/2(S\T=CD=#3
CG&DJ4d]EP3DF>N)^e)6:bK#]d.Ed^,J+6gBQ<H9f7+HKV&bQXDLS1Y^P^&UVX_A
@4I,2\/6W#@NAWYQ.?:FfcS#]COL9DR-SY2I)0DQ^bT.JV74fNP)=3^1cT90T)_,
1493X/bV(_S0B#[dD-?-bH\.0Mb,K2O&#R4ZN0;:6_8RI[E-+J8RM[YJQJ+[KRe:
8NMO#;c[\IS0<a20UFdAe?c:S=F/eKcGZ)23(:)SbQ(@RgN7&IR.L411bJD6HRDZ
)\0I<HHX2McBXR/X3.baAY#Q2Z80L[/^]EVVWBSY(b37+6)IV):@>T7Zf.7b?F6@
McNJTI-Xa+9>\;\R[=dGEKWR/cP_>.b.=W8:Z&4[ddMJ<,HJLc?L2_50>R+PfRV1
>]\LD(dd,?D=H7fa?,+9E4YXN;[[eJ2)^fTH/B:\>ZU<G,L;5[aZ@2Z>H9#U?QC?
RWYeR.L_?EQM^62e6C8bXX+U<1cOZg4aF.ETb5b[N(.WR<Y4\8R_cV:JL&)BFW0Q
BR:TcSIQ#TfO&bS4MCC?/Pc1M59M8^b>3gBQ.YO.[N]4512-2bc=I1--4Rc2M(R)
C7XB][/1e(&,PQf>f;@b7BG9-<DZd)3<:PVI</c&:6,=HR7RP(HET0GLDH&M_3J#
_[A<,Zc0M\.-]#8c3XEgFPOVb=N><g.>?d5#EVadR/T4T6Id@()Af4Y)Fb1b]A-S
=ecU/7bG)e)0.&V&ZH\SM/G^)eLLAE^/4@gRA2;;/9X^R78ZIaU=K><>fX2X@8-Y
-XO\c;4:,XKJfg@/Gf9H0WAJK,204FYEf;-9DB1ZAJAce?R>R&C>ARDZR+>EU(g)
UT7Ne-Og>9>LL]]T<4f-P4CUffO?E.9<)#SUHHG9YV1ZD443F;b,VD9[3.\T7P;T
OC3&,8fQO9a3US-,28YYU6f=2:F1;<,QL[TG^[Oa9-+L7;d^<(NJNA9Y6_c#\+bG
KaMJ-^:<->cU3]TL[^A##YdM8&->IIb:2XM:)0&<C]dfc1MGbHHSeG&6]<NPdOGL
?<-\2;EL@+Q[dCCgGFCZY/AObN+H?eZPJK;Eag^(>&&2]<WRT[P0,@G5fNa0NHOJ
e[A-?NVOAQ?2[e=0OZc-\)0X2:\aW-6E^1F(f=fY,HLRf-c/=^2>,26N#5^Z@/Ob
cHd;f=V6:=-Ec/KM/;V\OQ>A\2B;J\5IRZ>Q87\HP-D@XD-QL262:;N9V5G5d92+
#Q__[.?SYMY(;)UV=#=GMG:PRKTe;L^RUD;WgHU1Y_D0;>45KcCZ7&J)[[1\aM#V
)c59IeVH92(TB10c(;/C&>bE>g#5?g\?gUPTOTF[N=\F2ACa\=4U]YOG51([b\S6
^YHHT<HC)#e7LR^,_TB.)EFRL0436[WK9RA[QS?VI&2BX0KCc;LU))5I;gXgM_gc
ZX>GJ#(>W/PQ@A_aKS,,CN^Sd=b/XPB[#.8([(aY,\WO_O[6+?<];W4:=fSSPA3P
L8#-T96TS4eY0>83O>9F#V@>0IC#VLQPCEg@e=);Gf&LKEEBgS+?a8--MOJ9aJQB
G?16CMRNK<>_3ObTQV028a=/a9F-LTFeN-L_;[.M,eRaGC[?2e]f7O8><JT(EdU8
#6;&_6A,AQOM;NJedbWdfX#2=B:LBMAA0-Q6b;g[U;B]LG^Q=735f<90#X]:Oa^W
1C0[(KU.VgBFT&D[LeS.^L/[;1OgZU13a<7/HZU;Dc(d:OV6I[_>635:&N.SI;,Y
ELbV5FH4>F-e3Ra1QGY-ebN1JHA^_T;V#[O.>0&:1.0E)c[RVc+#/@I(22G[]T;\
&O4=](48N&/\W=T-(J^6&f<VF\0gA8Q#JZM=-_JIL>G.?CJ;,\<3]=F_T53G9d8<
#1)_\5PQ^^=AF:WHIF+RIY1FLLJG/LZfC^E/+Of[.ZB68&eL6SVE;C2&I1RdOCVL
c7gS1cQ3_#:abUIgH4X8ARd(^SIDP^)W<LZ-)16d;UD\S_@@/LeN&g9f[I=4E0BU
GLD>K7dc;(S4K\3B:dQ((V&.#<XM>8[_EE;72E4Kb58J2C;>5D2GA><TZR)_H817
9NQdg]2&M8Z7M9H&.H4E[VI?O5Y6ZE(&dZ,HZ,9R]eF^:U[Y/8>&Jg4P&<2RA3;=
&e)7M(_O3EeTJg0F@A_-SA,fNXab/_YEDE>;@]YGeD00@[Va7L;He^\I=X(P6=-:
GOSSV617JKKSML6.e@Ld4VCRD,GXFJfUX47?O,fN31D\I_OdIWPcQYd^@6H6/g(R
RG]7LXB(3/>:1EOM4)/f>LINYF(W\?/0@^T.Tb]d,I1b=\:Gg-[RU1eSDB4N4YMW
2KUB_2>B<eA8U6b6<5.3g0UVJR/KeR_;gJ@)F>5-Y0)U=Y_+;0U^M^6QD-,R-Y8I
[^PW>W.Hd7HH3c<LGVC@@dd>BbI0_N@O5)L=NRFVfWTc&^(YPTA5&VDI_9)#S]H,
<aVE#0Cc:1b_OS6#S6S/^\E)=JMOXQ4,VgR<f+dSX9e2A&0,)CM+=M2VT1Rf_(RI
e#@X62a_EF^g&6\=CK(AJEf03K_@:&>)cR[bd/XT-&;VPFb;Y9,K<(^.F0De[S65
8#R?1WY]f65721&X>5+8Y1PR):_W0)LHWca4(5I9(X-[A=P(C(H>21S1;=DK&/fG
]L]<9Jb,(Ud-PS)QP,4bH&K]cGI::@@7D6L-c]C\WM7;=9;.@XUg87V^6[c-I.5A
SEB=5NPGY)VffQ?Eb949Z^78=KKRQ>OFF05.(AY:JJFJZ6,VgP>^-\>NUa29_)>d
D(DIJG^1VdO[?&-F(_&]GALY2Y/<WQ8-cRZ)^Q,K>D&(+N6LJe.I0V1)?]I2RN>;
g_B]f9eQK44#Rf^H=7Lgb3I\,G90Y(a+d+-GG[\Wb?5+,L&_P#.UZ&b/bSCZ1b,.
Udf8@#U^,4HSW3597>;#d:]EG9g3S=I7UZ#\VQFbO\.\X4gdgX0_2H<LM=JGP)?>
;=VA#_0\#Q0]:JT&G2S:,3F3B7F&I/0C>@7;W_R?13]&<e/4L[(Ud6#=.MEN&,;1
gcNT0d5GUG6MN22G.1S+)D3I/D<6D95cY0TR00TLGDV>85KP#HT5I+A9a&S_Qc8Z
W8Y_UJ@bD.eT+>^J+U)R+0e>@+PdcF+UZ&_/_:[7Q=\JIWE\K69A;6HPI^PYJ8dS
L6MKL:K6I2dM^YO#KO6Jf5YR;g4B/_86S=a.:X<e?W<7Mc7=V/V-N@C4JA/&RST0
V2.(L;5C50@\LK,H+9ZX3(29DG0I[:KHN0KW7X(4^<e>c6W4d7:c88IX<-:a3O-C
-gDcGaIP0)T8N5ZJRCTU^M>TM?XS7+_RK+F&1T7LK(T&<B+CWRd8<1\L7(YR\81Q
-O\W.e3B>bfKfAIVe7&CBH7BQ+SOKV0[Ka[A^OJ4d]2S@g6O@aDYI(G=&>5/#MPf
b,I/9ce4f[?]W2:5K.X]eDQXLd\5TWC1XX>S8WCMfH/=,PgS(<8e&#b4,DN,-LA-
#^dKA@1C.WWY(/X&8;gV8]Q2XBE@<FGL?]QDggFJ.bSJ7HTLJP3/GXR2;8/=713:
>3U;bfILK/2ECR<fYZ?]IXXc#:IC&C?Q.SMMbfB^A+fHR6N/G@M3=,M9(Kf](7?H
UdF_T6cFN65)>?J(1[3U5;:)>.#2Ha(+:WKFO#DU<SIL=7^:WfYX4X<Z<:5(W?[P
I0fcZ1BGVeb:g]Z]MP^:.FTANO>G.ZR#0^P5E]YcNJXC]KDS;VeGLY.5fBLS+\cH
U_[fKgZe_7QF)Y.c\_S=@-N_ZE.c]KRe+&Q);_ID_&(_76\F?__7PU]H-gF<XVGB
YdFb7]-9)aJ-BH7B]C>ZFFKK>,CK\.B&g@gK@X9&]&D,)CUMbGcS/1g=FcK;G0]2
=YF_TG/N^Y>F8H?[_P4=^40b(9QG<+Gg7-9[(e-51af(HbDC^QR.C(1H@9Vd#8U]
2Q2UM@??(;-9-E]?e@HR.RX0aDGgAGZRS+8?e?H+?H?#(B(0Lc2f,_(#2GggS1XV
[f8WUH>>=faQ-1CR:C&I.cKEF(OE>C.G.5X0NIcE7>I2>D:-dZ8RP3bAK:#M_E18
/g#=3T<,]O2WDT]6;4g7-Q4D:3),a>d3(:T#)fdNXfPc5Q]a=80J>P9X13e,;1U@
-b9GBFcW7]Zg=/6]/P\G_F1IUU@5RS0H3T=,NSQ)[d:]P9=D,6YDA]EW3QJ@,0D_
.S\8+\S<IIQ8:gA)#J#TCZPNg6\-9QaJ^6Y(<MNX&@\>a@\/2FeJ=1F2dL\(+/Mc
TWDZeNO-X72G<U#O6UH.gY_2AGF89=);^;?(2Y[=>,R\#?>=N5ZFVC,6K?SZ>^I:
W6S-CDX]IdZc;agR9454X0+5<e)S:DV=W:c(_dB6V)D-Q;=_Hge;aY5Wf;T;:J6/
Lb/-63)S5.&AbR7J3LA-I.,K0aIR0):7FW#^FD#gFRE9D3#DPY#L5Z7]7]D#G\3)
T5LdOW[T9ISX+/++-;2U.+,(UZZ&DKe9:O&,Q\>T6#cPB]NRBa=-@BN/;cJ2Wf9.
f([;+4Z?(UEF.O,...Y_@FD.H7-J/.HFYJH[EGUR.fceG[4-dXJ4O?7.DBIY0ZV>
D(=G,H]fJ^7+#Y1^\LT@bgO7+HV\aLCYW-4WNAHG?BVT&CUgP96E+-;F?MY:[,bb
?17D(8V>N9K9Ff/,<(f&]4]WZf]-[4J)(b5cWB?R)Ma7[g#gC(DUJP4KaQd\Z;-V
@WE;G#7BX_9W&Q]TL/2b9/c]eK6DF610]A51+FAL>\g\A_ZLLYE(1bBgS4:b)H^e
_FMSPD1XJ+-BT)L?4S.X<9(2b3fe[VN5R@aeL-AMf-IBe2N2\[JJ/RW??Bb4gA(P
MbU;WM4b^)9P04LRK<EM-[&/ZNJf&I6aX1dKE?.aZUKK>[</(@I;e7,O^YBCZ0^R
AXW(2fI.-Q6]8UUe9>80B9.\I@A4:OF(bE5()TH(RbG>QI9,D+28XD:H[TN\XTf&
5JUAO6LOTgQfVP4@DDY)N(Yc<I>\@TI.<SPY#4-]/d0c<f4(VT44b>#(;bMHV4HJ
4#JNF[&?94/=->f=ab7a_1+=3d&39IV/L8^bIK+2FPB0f.<d)\BFLDIC^X1:Oa(R
b#;Hb43D<W@ZVK:,@,Ha>\Z50^V2O>]W.O;7OQ8ZbZ=K&XHC-HAU[g#HU^SegAA2
D]W(3F=>N]CLMO&e]Z8]e]&VCOW_S9fbdga.S@#[(&f<RHRbJe&d#I1TS4,#7@FZ
X+OcJ:6?/YefBFL7_Ra<).d7IdN/VJRGRHGZ2&[K4WY89ZGJ@X9PC-/b;=@R4)-R
W(S._&2fG<R?#/4L\PC1P1H&;4,?f0CTYP7.CeYP>Y9(Be3V3B0@I345S[U^M8D6
Q_N9c[[7BbAPQaO(([=@C.?)_@&#X<&RR]:CPgg9[bSfPfI6BbOD1TBAB#>c;)Z&
6@W&&GEaDFe(448eH+W1H=;<,LZ#:KeFA^?A@RSUX:Db7K_]SMDHM-D:2Jb7,g?V
1.4D@#GS(c\LJXJ@#dV/eO)3MdTJ:D-<+I)1SWDd_MdGKA+1N_B]gI0RFZ8X#M?H
cOM_S_YH#.>NeO-<=]c6)@_ZI?8Gf0N)P91<@&I)SdOJaS15@Y9CEK>?g^ZBCV3P
<WR=f-@fGRUE,\eg7dG-YEVF4>98RUZFQU.1=,Q?[VT:#XV-^G=H55IE=gc.BG@2
aVFgK5EGI^8TYQ6E.AP9C\Db4+CYNL#;5?f+/0[dU4M4SLM?JH2R]Cd-WXd8>^U<
J8@-MK5-E&:^7NG-bEHOLCfCd9_\#QJCYTP2e^H@e?dRc#0/\?&\U/PSN(N0[K]@
A#0ACSf5G@K0bfWa@,B]-8EX#6+fKU&Kc74R)bHbBUJESdYBR0VN6_=5dBJ0:XAD
6Pb-<3-=\X^A:&-c(8HgEWdB-/KR^X2_f?RDD=G6=?1H-_b-4_.HU6?R0+=Kd01b
+ZFT<YH+W>c&;3;1)XV@a#OS>YLHW\#3=5#,,2D=IIMggALEXLXZA0gS3HcYcT5;
R[.G;3>O/Pcf?1dO\<TT8GgH1]7CfAg0F=I)JabE=&><^UX^HI9;d9JL1bQ3.[CH
7R<HBL:(+=TH<PbNS@5T#)faJE0eG^VbB=,EJ<.WbY;EGX5(K1a4:=GZ];L=PR=3
O<L/=KdM>R?KB3bM1=g\G3N)GBQb<A2\A9b8N<KWbe4d3dbZK>aY1B&]._ZW(MQU
eI-E=0W.KUg:WD(+TbOE/GT7]3c5a)IPTLKFJ(Yfb7FKaDg?EYWBa>g1[W=W+&fb
3<XS:O4^\:HC&.VK;H8X245gIU4b0A2Q>K\@=6bJ.2&S04;.Sd@U)RZa6f8K:=Pa
(0\Y->4&652ARFc]2<fS=fWPYYX9\SSV^><ac7FOM6^b,FD7.Xg;):0=8W2_CI3@
&=M?^B3;AT;8V@)Q<bMN@NMFdINRM8MJd7d6VM@\fC;0F5ZK(8OggSa;HQ,:7[V&
18^O@fXg<TM9G5;b:^eLVcE@4[+K4&16_DXa&cfc>0482]=C_;)gVIFYH(Q@:RVJ
[_.b65==,K^DN=0XDI=NYD.S,.+C0JW[.7Z<C4CY.LZbQ\46B=Q[ISPb.bT/P89^
+:]UOfX8V^DPSHMCOI[9D?DR>#W9S,A>dHWTQ7,g8G>?bV;1+91QbOYS-+I<S+/_
g?_OJQKOQ?gXU+4ePc;2JW[Vf?I;-Y9J>1,d:f8_??-ZTBKc#-5#KD@dD&GYT4^<
UQLbA)??X(f+^[g0&Q+3R?94Z7PK_U34]3\ITE]?9YXd/IY<8E]4AO,/TPAM+_Z)
M2)7fWS&;2N>^>P2)6^F\B&=(gJ<P;;6:;aR3/,#VLeEWHb^#gL_GT(^K^YDA7^9
I&Qf(;KA0=K4+Ab8<#FCL&[+ZEJCSAfKDeBJM[SI_g:31SXX?]e[W7Ld:7M+RWKE
;Y)RHXT(-NW@I^XVd?61NeY<QaP#]YE5TI_E_O=6GaCPX?L/1&[7)V,ZS]O.c/=B
(IM>P7Z1aS;Sb2WY:24c?3J8;)3759e8^97R&G.GK>);=?UZ7:\?W6_?@C]_[=-2
JK;TV+LVe<3DU:PgFLPDSIBL-YX2PC=Y(J&<,a,:RI/G<J[&#TG]?/=/b?f)[^4W
M,Q.VdAa:J5MWfLC#]8\35/1_ASUY)IBQS\P-7-L<G,A?FNR:MQg^2)1VFF9_(b&
gUK@TQ:GA3UK0+>DGfG&D##a9#0TRH#FZ@9W54O#X49HQO5??AXTK4)4WBcGeeXP
#aUP(&6W2EF1M6a1Gd:3/(A#T^d9.ENW;B-WP#/^d2Q?3-#@GD.[_Tg,T1-<QfLYS$
`endprotected


`endif // GUARD_SVT_APB_CHECKER_SV
