

`ifndef GUARD_SVT_AXI_BASE_SLAVE_COMMON_SV
`define GUARD_SVT_AXI_BASE_SLAVE_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_axi_defines.svi"
//`include "svt_axi_qvn_transaction.sv"

// Note:
// Throughout this file, the term 'driver' is used to refer to the active
// component on this port.  For UVM this object is extended from uvm_driver.
// For VMM this object is extended from vmm_xactor.

`define SVT_AXI_SLAVE_IS_SIGNAL_ENABLED(axi_signal) \
(cfg.axi_interface_type != svt_axi_port_configuration::AXI4_LITE) && \
( \
  (cfg.axi_interface_type != svt_axi_port_configuration::AXI4) || \
  (cfg.axi_signal == 1) \
)

`define SVT_AXI_READ_DATA_CHAN_IDLE_VAL(val) \
driver_mp.axi_slave_cb.rid    <= {`SVT_AXI_MAX_ID_WIDTH{1'b``val}}; \
driver_mp.axi_slave_cb.ridunq <= {1'b``val}; \
driver_mp.axi_slave_cb.rresp  <= {`SVT_AXI_RESP_WIDTH{1'b``val}}; \
driver_mp.axi_slave_cb.rdata  <= {`SVT_AXI_MAX_DATA_WIDTH{1'b``val}}; \
driver_mp.axi_slave_cb.rlast  <= 1'b``val; \
`ifdef SVT_ACE5_ENABLE \
if(cfg.rdata_chunking_enable)begin \
  driver_mp.axi_slave_cb.rchunkstrb  <= {`SVT_AXI_MAX_CHUNK_STROBE_WIDTH{1'b``val}}; \
  driver_mp.axi_slave_cb.rchunknum   <= {`SVT_AXI_MAX_CHUNK_NUM_WIDTH{1'b``val}}; \
end \
`endif \
if(cfg.check_type == svt_axi_port_configuration::ODD_PARITY_BYTE_ALL || cfg.check_type == svt_axi_port_configuration::ODD_PARITY_BYTE_DATA) \
  driver_mp.axi_slave_cb.rdatachk  <= {`CEIL(`SVT_AXI_MAX_DATA_WIDTH,8){1'b``val}}; \
if(cfg.ruser_enable) begin \
  driver_mp.axi_slave_cb.ruser  <= {`SVT_AXI_MAX_DATA_USER_WIDTH{1'b``val}}; \
  if(cfg.check_type == svt_axi_port_configuration::ODD_PARITY_BYTE_ALL) \
    driver_mp.axi_slave_cb.ruserchk  <= ~{`CEIL(`SVT_AXI_MAX_DATA_USER_WIDTH,8){1'b``val}}; \
end else begin \
  driver_mp.axi_slave_cb.ruser  <= {`SVT_AXI_MAX_DATA_USER_WIDTH{1'bz}}; \
  if(cfg.check_type == svt_axi_port_configuration::ODD_PARITY_BYTE_ALL) \
    driver_mp.axi_slave_cb.ruserchk  <= {`CEIL(`SVT_AXI_MAX_DATA_USER_WIDTH,8){1'bz}}; \
end  

`define SVT_AXI_WRITE_RESP_DATA_CHAN_IDLE_VAL(val) \
driver_mp.axi_slave_cb.bid    <= {`SVT_AXI_MAX_ID_WIDTH{1'b``val}}; \
driver_mp.axi_slave_cb.bidunq <= {1'b``val}; \
driver_mp.axi_slave_cb.bresp  <= {`SVT_AXI_RESP_WIDTH{1'b``val}};  \
if(cfg.check_type == svt_axi_port_configuration::ODD_PARITY_BYTE_ALL) \
  driver_mp.axi_slave_cb.brespchk  <= ~{`CEIL(`SVT_AXI_MAX_BRESP_USER_WIDTH,8){1'b``val}}; \
if(cfg.buser_enable) begin \
  driver_mp.axi_slave_cb.buser  <= {`SVT_AXI_MAX_BRESP_USER_WIDTH{1'b``val}}; \
  if(cfg.check_type == svt_axi_port_configuration::ODD_PARITY_BYTE_ALL) \
    driver_mp.axi_slave_cb.buserchk  <= ~{`CEIL(`SVT_AXI_MAX_BRESP_USER_WIDTH,8){1'b``val}}; \
end else begin \
  driver_mp.axi_slave_cb.buser  <= {`SVT_AXI_MAX_BRESP_USER_WIDTH{1'bz}}; \
  if(cfg.check_type == svt_axi_port_configuration::ODD_PARITY_BYTE_ALL) \
    driver_mp.axi_slave_cb.buserchk  <= {`CEIL(`SVT_AXI_MAX_BRESP_USER_WIDTH,8){1'bz}}; \
end     

  // signal drive format - method name ,signal width,signal name ,signal value , AXI4 Lite disabled?,AXI3 disabled ?,category disable?,cfg_enable ?
`define SVT_AXI_SLAVE_SIGNAL_DRIVE(name,width,sg_name,val,lite_disable,axi3_disable,interface_category_disable,cfg_enable) \
  if ((cfg.axi_interface_type == svt_axi_port_configuration::AXI4) && \
    ((cfg.axi_interface_category == svt_axi_port_configuration::``interface_category_disable) || \
    (!(cfg_enable)))) begin \
    driver_mp.axi_slave_cb.``sg_name <= width'bZ; \
  end \
  else if((cfg.axi_interface_type == svt_axi_port_configuration::AXI4_LITE) && lite_disable) begin \
    driver_mp.axi_slave_cb.``sg_name <= width'bZ; \
  end \
  else if((cfg.axi_interface_type == svt_axi_port_configuration::AXI3) && axi3_disable) begin \
    driver_mp.axi_slave_cb.``sg_name <= width'bZ; \
  end \
  else begin \
    driver_mp.axi_slave_cb.``sg_name <= val; \
  end

  // Signal sample format - method name ,signal name ,default signal value , AXI4 Lite disabled?,AXI3 disabled ?,cfg disabled
`define SVT_AXI_SLAVE_SIGNAL_SAMPLE(name,sg_name,val,lite_disable,axi3_disable,interface_category_disable,cfg_enable) \
  if ((cfg.axi_interface_type == svt_axi_port_configuration::AXI4) && \
    ((cfg.axi_interface_category == svt_axi_port_configuration::``interface_category_disable) || \
    (!(cfg_enable)))) begin \
    observed_``sg_name = val; \
  end \
  else if((cfg.axi_interface_type == svt_axi_port_configuration::AXI4_LITE) && lite_disable) begin \
    observed_``sg_name = val; \
  end \
  else if((cfg.axi_interface_type == svt_axi_port_configuration::AXI3) && axi3_disable) begin \
    observed_``sg_name = val; \
  end \
  else begin \
    observed_``sg_name = monitor_mp.axi_monitor_cb.``sg_name; \
  end

`define SVT_AXI_SLAVE_VALID_SIGNAL_SAMPLE(sg_name,interface_category_disable) \
   if ((cfg.axi_interface_type == svt_axi_port_configuration::AXI4) && \
       (cfg.axi_interface_category == svt_axi_port_configuration::``interface_category_disable)) \
   begin \
     observed_``sg_name = 1'b0; \
   end \
   else begin \
     observed_``sg_name = monitor_mp.axi_monitor_cb.``sg_name; \
   end

`define SVT_AXI_SLAVE_CHAN_DISABLE_CONDITION(interface_category) \
  ((cfg.axi_interface_type != svt_axi_port_configuration::AXI4) || \
      ((cfg.axi_interface_category != svt_axi_port_configuration::``interface_category) && \
      (cfg.axi_interface_type == svt_axi_port_configuration::AXI4))) 

`define SVT_AXI_SLAVE_IS_ACTIVE_QUEUE_FULL_RD_CHANNEL \
  (((active_xact_queue.size() >= cfg.num_outstanding_xact) && (cfg.num_outstanding_xact != -1)) || \
   ((active_read_xact_count >= cfg.num_read_outstanding_xact) && (cfg.num_outstanding_xact == -1)))

`define SVT_AXI_SLAVE_IS_ACTIVE_QUEUE_FULL_WR_CHANNEL \
  (((active_xact_queue.size() >= cfg.num_outstanding_xact) && (cfg.num_outstanding_xact != -1)) || \
   ((active_write_xact_count >= cfg.num_write_outstanding_xact) && (cfg.num_outstanding_xact == -1)))

`define SVT_AXI_SLAVE_IS_ACTIVE_QUEUE_FULL_WR_CHANNEL_OPTIMISTIC \
  (((active_xact_queue.size() > cfg.num_outstanding_xact) && (cfg.num_outstanding_xact != -1)) || \
   ((active_write_xact_count > cfg.num_write_outstanding_xact) && (cfg.num_outstanding_xact == -1)))

`define SVT_AXI_SLAVE_WRITE_XACT(xact) \
      ((xact.xact_type == svt_axi_transaction::WRITE) || \
        ((( xact.xact_type == svt_axi_transaction::COHERENT) && \
          ((xact.coherent_xact_type == svt_axi_transaction::WRITENOSNOOP)|| \
           (xact.coherent_xact_type == svt_axi_transaction::WRITEUNIQUE)|| \
`ifdef SVT_ACE5_ENABLE \
           (xact.coherent_xact_type == svt_axi_transaction::WRITEUNIQUEPTLSTASH) || \
           (xact.coherent_xact_type == svt_axi_transaction::WRITEUNIQUEFULLSTASH) || \
           (xact.coherent_xact_type == svt_axi_transaction::STASHONCEUNIQUE) || \
           (xact.coherent_xact_type == svt_axi_transaction::STASHONCESHARED) || \
           (xact.coherent_xact_type == svt_axi_transaction::STASHTRANSLATION) || \
`endif \
           (xact.coherent_xact_type == svt_axi_transaction::WRITELINEUNIQUE)|| \
           (xact.coherent_xact_type == svt_axi_transaction::WRITECLEAN)|| \
           (xact.coherent_xact_type == svt_axi_transaction::WRITEBACK)|| \
           (xact.coherent_xact_type == svt_axi_transaction::EVICT)|| \
           (xact.coherent_xact_type == svt_axi_transaction::WRITEBARRIER)))))

`define SVT_AXI_SLAVE_READ_XACT(xact) \
     ((xact.xact_type == svt_axi_transaction::READ) ||  \
      (( xact.xact_type == svt_axi_transaction::COHERENT) &&  \
       ((xact.coherent_xact_type == svt_axi_transaction::READNOSNOOP) || \
        (xact.coherent_xact_type == svt_axi_transaction::READONCE) || \
        (xact.coherent_xact_type == svt_axi_transaction::READONCECLEANINVALID) || \
        (xact.coherent_xact_type == svt_axi_transaction::READONCEMAKEINVALID) || \
        (xact.coherent_xact_type == svt_axi_transaction::READSHARED) || \
        (xact.coherent_xact_type == svt_axi_transaction::READCLEAN) || \
        (xact.coherent_xact_type == svt_axi_transaction::READNOTSHAREDDIRTY) || \
        (xact.coherent_xact_type == svt_axi_transaction::READUNIQUE) || \
        (xact.coherent_xact_type == svt_axi_transaction::CLEANUNIQUE) || \
        (xact.coherent_xact_type == svt_axi_transaction::MAKEUNIQUE) || \
        (xact.coherent_xact_type == svt_axi_transaction::CLEANSHARED) || \
        (xact.coherent_xact_type == svt_axi_transaction::CLEANSHAREDPERSIST) || \
        (xact.coherent_xact_type == svt_axi_transaction::CLEANINVALID) || \
        (xact.coherent_xact_type == svt_axi_transaction::MAKEINVALID) || \
        (xact.coherent_xact_type == svt_axi_transaction::DVMCOMPLETE) || \
        (xact.coherent_xact_type == svt_axi_transaction::DVMMESSAGE) || \
        (xact.coherent_xact_type == svt_axi_transaction::READBARRIER))))

/** @cond PRIVATE */
typedef class svt_axi_checker;
typedef class svt_axi_slave;
typedef class svt_axi_port_monitor;

`ifndef SVT_VMM_TECHNOLOGY
typedef class svt_axi_slave_agent;
`else 
typedef class svt_axi_slave_group;
`endif

`ifndef SVT_AXI_DISABLE_DEBUG_PORTS
class svt_axi_base_slave_common#(type DRIVER_MP = virtual `SVT_AXI_SLAVE_IF.svt_axi_slave_modport,
                            type MONITOR_MP = virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport,
                            type DEBUG_MP = virtual `SVT_AXI_SLAVE_IF.svt_axi_debug_modport
                            ) extends svt_axi_common;
`else
class svt_axi_base_slave_common#(type DRIVER_MP = virtual `SVT_AXI_SLAVE_IF.svt_axi_slave_modport,
                            type MONITOR_MP = virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport
                            ) extends svt_axi_common;
`endif

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  /** Custom type definition for virtual AXI interface */
  typedef virtual svt_axi_stream_if.svt_axi_stream_slave_modport STREAM_DRIVER_MP;
  /** Custom type definition for virtual AXI interface */
  typedef virtual svt_axi_stream_if.svt_axi_stream_monitor_modport STREAM_MONITOR_MP;
  typedef virtual svt_axi_slave_if.svt_axi_slave_async_modport AXI_SLAVE_IF_ASYNC_MP;

  // For a snoop capable slave, this will be set. Initialization should be
  // based on this interface
  typedef virtual svt_axi_master_if.svt_axi_slave_modport AXI_IC_SLAVE_IF_ASYNC_MP;

   
  // ****************************************************************************


  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ** AXI Port monitor for callbacks */
  svt_axi_port_monitor axi_port_monitor;
  
`ifndef SVT_VMM_TECHNOLOGY
  svt_axi_slave_agent slave_agent;
`else 
  svt_axi_slave_group slave_agent;
`endif

  //vcs_lic_vip_protect
    `protected
BP(&@^.c<H-<E=Z_+e9=EMWVCM<+;;^STD4R.bRQ]#dZQSG(4G6-4(/_;+-.6@P^
CfeaQ?fO#5N5Ma;R(@@PPQf/[P6@9cMG?36Gd81W@PL2\^+A1#2C7#UKT=:b8]X&
AXb&=_=DPc5_g#WA]V\TQ0^,T\KY_@QT.I=eYd^7/9f\;TC[G^O>/O_#?H\HDMIK
)U.XBRTQS^_D9=?f5Bc.c.4&B.G?^/5-1=T0>W[@()1_e?C+@UQU+gQ0HTBFM(6B
P9A4L=b=C:;S@6A:=:_b\WZ2RY]aD[Y<U2F?Fc,c0LY32DAEbg06G^]gMQcJXS\2
ABAf4a@QD>COZ<2+;(:AY)#K(:I+F4U[DOSG?>AD/;MLX:@CRg&&aW;FFIDA(^b\
L(.6aI;YV66QL]>,ebO4,Y&^d1N6^1)B:ES(dZ0UKR9)c8+Z-@gQGEFF^Bd_WJ5>
>ONd;H(7ffg[KMU,)68AcZ,CNDEJA:f=VLDJEY5FXDD^G=ZW]JFaDP[++SD6C@,B
&9AX6+RfX98;(\:5@]g\.>ZX83W;-A3I&PD^\8gaa,^Q1U)ZV..=UM3I9H.[Jd&P
35:ZTZbVaVD+_;>?>e9<-NT+T::3g1?0afX^>K4Z]=bH&gU?7E:Y[GW0WG[A+M#B
C)M#R4<L+fO\g8&ILSF?YbY&M<>##HE8A^g]^Ye?YUY>QI&5g(7^_M:H;aVAKY1c
a?C(^KX,>GB7VWJ,]INf;dgRbB3OO.HJ:]3V)dEI9=b\[/:3B7Ne@?YT]ZY64B&<
^I#FObg8V?TQ:8,W8U=L>:dD5=Q4d_c6NGe\37U<>;TgH+8A2[/\UHYDO9RT4<I7
#52VIQN(TU,]-Vf5/b+XTI<T@bI\<Ca[B]W^N2^cP.JQfOM22<-/CdPMQfd@^YK5
T=E^,e8R:-+b0UP4GG@7E-UK#a[.0P-7YVBUgZIL1W2c8=?WZZUO<_)(XYQ1H>7a
@=W6L2>OE/=JV-<H:F4deTX1T?]&P8;_2AQ5dfWYG4fI3J1^&M7I/.7S6WMU7X7\
Zb0U)Q]-^8eGd07M7OA<)SF2YBVb-:;+aB(KQa.+Gb>/:6YJbM2_I]gOF5,B(0#P
OH;H5fPXZ0FBDL4#N5a#]@.;9e4,(H\B-1S#[^<dX<S,eJO[S+a.?-A43:P+dW^S
HD#I[[3V_cc7;EU5Z<]:?^M1TQ,KJ]A,1?KIfNeKWgd(NbK[XaZ[4ZaPDN6;RgeY
b-b:.,BfR(X+G0>H6TAc2VXIg=>67ZAS(]53R/4e6]2K:OTEV5I2DL<2a&EWf7<E
(f(e?BOP[2&54(O8YNXU4;B6KP3BO/WD.JJS&2^>eJ4:bWJ;5;,Ge[QI<RZ<G^.Y
HQG0fL9YN7D[XSCa-/ZDM@dea>18UU[+HFHZ[g0C_N/aO5b8B)M8,EH2@EJO&90[
-)ZQFc,@PAHHB;>[&D36,A980^;O<OJ&;&:KGQQJP_5JL3DU63.YZZ7;X3_6bZa\
/4Vb)fF&DZAedUcC#A[N9X4YaXPZ#EVWMaE6LHTf;LIN28T5JQ<SaH-&IB^&3/Q@
8G,LX6=[:3-.RbU>NB]/IV(I;:e>RGb5Y]V6NJ9LMR-P9BAg4?\?F/\#<K0gZGIV
>Nc+G\+gUG[_Z3>AZ.<F:71,G3EaV(NT02O5-g5]B7B=XdSM]FSA](5-5;fS0-D>
)Y:HI#f</X07G)aZ/gb1HS1,SD:R0LH&9:8f40]]Tg[BALbW3=.Q2LP6S]N&BC(R
66<6Ua[W5]O8=[f&<fPa4D6cXdU<E7V^X0S:\\T0&;.?;AW@CZAc)\E4g/CeU>A]
(9;-9b5135LV1LEF=O/@I-JJXJ384L@;JcOS6JM:9da)BU,e7NZF=E]B+XgJ#+?YT$
`endprotected

  /** This variable indicates the size of write response buffer*/
    int write_response_buffer_size = 0;
  /** This variable indicates the size of write address buffer*/
    int write_addr_buffer_size = 0;
   /** This variable indicates the size of write data buffer*/
    int write_data_buffer_size = 0;
   /** This variable indicates the size of read address buffer*/
    int read_addr_buffer_size = 0;
   /** This variable indicates the size of read response buffer*/
    int read_response_buffer_size  = 0;

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Slave VIP modport */
  protected DRIVER_MP driver_mp;
  protected MONITOR_MP monitor_mp;
`ifndef SVT_AXI_DISABLE_DEBUG_PORTS
  protected DEBUG_MP debug_mp;
`endif
  protected STREAM_DRIVER_MP stream_driver_mp;
  protected STREAM_MONITOR_MP stream_monitor_mp;
  protected AXI_SLAVE_IF_ASYNC_MP axi_slave_async_mp;
  protected AXI_IC_SLAVE_IF_ASYNC_MP axi_ic_slave_async_mp;

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
 /** @cond PRIVATE */

  /** Slave configuration */
  protected svt_axi_port_configuration cfg;

`ifdef SVT_UVM_TECHNOLOGY
 /** Handle to the UVM Slave driver */
`elsif SVT_OVM_TECHNOLOGY
 /** Handle to the OVM Slave driver */
`else
 /** Handle to the VMM Slave transactor */
`endif
  protected svt_axi_slave driver;

  /** Variable that stores the read transaction count */
  protected int read_xact_count = 0;

  /** Variable that stores the write transaction count */
  protected int write_xact_count = `SVT_AXI_WRITE_XACT_COUNT_BASE;

  /** 
    * Variable that stores the stream transaction count 
   */
  protected int stream_xact_count = 0;

  /** Variable stores the number of active read xact count */
  protected integer active_read_xact_count ;

  /** Variable stores the number of active write xact count */
  protected integer active_write_xact_count ;

  /** 
   * Internal flag to indicate that wvalid is received. 
   * resets the flag when it gets added to queue 
   */
  protected bit received_wvalid = 0;

  /**
   * Internal flag to indicate that awvalid is received.
   * resets the flag when it gets added to queue
   */
  protected bit received_awvalid = 0;
  
  /** log_base_2 of data width in bytes */
  protected int log_base_2_data_width_in_bytes;

  /** data width in bytes */
  protected int data_width_in_bytes;

  /** Internal clock count from arvalid to arready.*/
  protected int arvalid_to_arready_delay ;

  /** Internal clock count from awvalid to awready.*/
  protected int awvalid_to_awready_delay;

  /** Internal clock count from wvalid to wready.*/
  protected int wvalid_to_wready_delay;

  /** Internal clock count from tvalid to tready */
  protected int tvalid_to_tready_delay;

  /** Internal variable to indicate  arvalid. */
  protected logic observed_arvalid;

  /** Internal variable to indicate  awvalid. */
  protected logic observed_awvalid;

  /** Internal variable to indicate  wvalid. */
  protected logic observed_wvalid;

  /** Internal variable to indicate  awready. */
  protected logic observed_awready;

  /** Internal variable to indicate  wready. */
  protected logic observed_wready;

  /** Internal variable to indicate  arready. */
  protected logic observed_arready;

  /** Internal variable to indicate tready */
  protected logic observed_tready;

  /** Internal variable to indicate  wlast. */
  protected logic observed_wlast;

  /** Internal variable to indicate  tlast. */
  protected logic observed_tlast;

  /** mask used for sampling tdata based on tdata_width*/
  protected bit[`SVT_AXI_MAX_TDATA_WIDTH-1:0] sample_tdata_mask;

  /** mask used for sampling tuser based on tuser_width*/
  protected bit[`SVT_AXI_MAX_TUSER_WIDTH-1 :0] sample_tuser_mask;

  /** mask used for sampling TID based on tid_width*/
  protected bit[`SVT_AXI_MAX_TID_WIDTH-1:0] sample_tid_mask;

  /** mask used for sampling tdest based on tdest_width*/
  protected bit[`SVT_AXI_MAX_TDEST_WIDTH-1:0] sample_tdest_mask;

  /** Internal queue of transactions */
  protected `SVT_AXI_SLAVE_TRANSACTION_TYPE active_xact_queue[$];

   /** Internal queue of transactions */
  protected `SVT_AXI_SLAVE_TRANSACTION_TYPE active_memory_update_queue[$];

 /** Internal queue of transactions */
  protected `SVT_AXI_SLAVE_TRANSACTION_TYPE locked_xact_queue[$];

  /** Internal queue to buffer the incomming read transactions */
  protected `SVT_AXI_SLAVE_TRANSACTION_TYPE read_xact_buffer[$];

  /** Internal queue of buffer the incomming write transactions */
  protected `SVT_AXI_SLAVE_TRANSACTION_TYPE write_xact_buffer[$];

  /** Current owner of the read data channel */
  protected `SVT_AXI_SLAVE_TRANSACTION_TYPE read_data_chan_owner; 

  /** Current owner of the write response channel */
  protected `SVT_AXI_SLAVE_TRANSACTION_TYPE write_resp_chan_owner;

  /** Object used for randomizing a transaction to drive random values during idle*/ 
  protected svt_axi_master_transaction idle_val_rand_factory;
  
  /** Internal queue to store write transactions in the order in which address is recieved*/
  protected `SVT_AXI_SLAVE_TRANSACTION_TYPE    write_addr_order_xacts[$];

 /** Internal queue to store write transactions in the order in which data is received*/
  protected `SVT_AXI_SLAVE_TRANSACTION_TYPE    write_data_order_xacts[$];

  /** Stores the last sample time. Used for calculating clock period */
  protected time last_sample_time = -1;

  /** The cycle in which last arvalid was driven high*/
  protected int last_arvalid_cycle = 0;

  /** The cycle in which last arready was sampled high*/
  protected int last_arready_cycle = 0;

  /** The cycle in which last awvalid was driven high*/
  protected int last_awvalid_cycle = 0;

  /** The cycle in which last awready was sampled high*/
  protected int last_awready_cycle = 0;

  /** The cycle in which last wvalid was driven high*/
  protected int last_wvalid_cycle = 0;

  /** The cycle in which last wready was sampled high*/
  protected int last_wready_cycle = 0;

  /** The cycle in which last rvalid was sampled high*/
  protected int last_rvalid_cycle = 0;

  /** The cycle in which last rready was sampled high*/
  protected int last_rready_cycle = 0;

  /** The cycle in which last bvalid was sampled high*/
  protected int last_bvalid_cycle = 0;

  /** The cycle in which last bready was driven high*/
  protected int last_bready_cycle = 0;

  /** The cycle in which last tvalid was sampled high */
  protected int last_tvalid_cycle = 0;

  /** The cycle in which last tready was driven high */
  protected int last_tready_cycle = 0;
  
  /** this flag is set when reset is asserted synchronous or asynchronous*/
  protected bit dynamic_reset_flag = 0;
  
  /** this flag is used to print message when the stream signal enables are deasserted */
  bit stream_enable_info = 1;

  /** Slave Transaction */
  `SVT_AXI_SLAVE_TRANSACTION_TYPE global_parity_xact;


  // ****************************************************************************
  // SEMAPHORES
  // ****************************************************************************
  /** semaphore that controls access to active_xact_queue. */
  protected semaphore active_xact_queue_sema;

  /** semaphore that controls access to active_xact_queue. */
  protected semaphore active_memory_update_queue_sema;

 /** Semaphore that controls deassertion of AWREADY. */
  protected semaphore deassert_awready_sema;

  /** Semaphore that controls deassertion of ARREADY. */
  protected semaphore deassert_arready_sema;

  /** Semaphore that controls deassertion of WREADY. */
  protected semaphore deassert_wready_sema;
  
  /** Semaphore that controls deassertion of TREADY */
  protected semaphore deassert_tready_sema;

  /** Semaphore for the delayed response port */
  protected semaphore delayed_response_sema;

  /** Stores the sampled value of tvalid signal */
  protected logic observed_tvalid;



  // ****************************************************************************
  // Local Events 
  // ****************************************************************************

  /** Event indicating that all signals sampled */ 
  protected event is_sampled;

  /** Triggered after any transaction ends */
  protected event transaction_ended;

  /**
    * An event that is triggered every time a valid is asserted or a handshake
    * takes place.
    */
  protected event bus_activity;

  /**
    * An event that is triggered every time when address for data before address got
    * received and aligned data and wstrb.
    */
  protected event align_data_and_wstrbs_ev;

  /** An event that is triggered when a wait_for_awvalid is called */
  protected event ev_wait_for_awvalid;

  /** An event that is triggered when a wait_for_wvalid is called */
  protected event ev_wait_for_wvalid;

  /** An event that is triggered when receive_read_addr is called */
  protected event ev_receive_read_addr;

  /** @endcond */

  // ****************************************************************************
  // TIMERS
  // ****************************************************************************
  /** Timer used to track rready assertion */
  svt_timer rvalid_rready_timer;

  /** Timer used to track bready assertion */
  svt_timer bvalid_bready_timer;

  // ****************************************************************************
  //                        SNOOP PROCESSING RELATED MEMBERS 
  // ****************************************************************************
  /** log_base_2 of cache_line_size of master to which this port
    * is connected
    */
  protected int log_base_2_cache_line_size = 0;

  /** Variable that stores the snoop transaction count */
  protected int snoop_xact_count = 0;

  /** Internal queue of active snoop transactions */
  protected svt_axi_ic_snoop_transaction active_snoop_xact_queue[$];

  /** 
    * Semaphore that controls access to the active xact queue. 
    * Any access to the active_xact_queue should be via this
    * semaphore. This is because there are multiple processes
    * accessing the queue and it is neccessary to have this kind
    * of access control to ensure consistent behaviour
    */
  protected semaphore active_snoop_xact_queue_sema;

  /**
    * Semaphore that controls access to the code that decides
    * whether there is a snoop/resp to the same cache line.
    * This semaphore is returned in 0 time. 
    */
  protected semaphore same_cache_line_sema;

  //vcs_lic_vip_protect
    `protected
d#FC:^,<)MO4<E^]N-VBG#=8IB6+dFA2J=D59D\^R9WCGDU4dP7_((7<XB;&[\3>
[N=fUG@S\:/GH-->GQb_TA<JO-<#Y)a64Wc)e@HF\390L5G0eZ04-#CY]TU5GV\&
:AI-2JICXS9;VfI9OIM4(O^M.6efa69K_Q8JP0A?5D-VZP/Od2NVeJ4HQ]&W@RaF
&=91Qa)=7>_Rb[-/R+4AFg<WKIJTOL>f>dSN@c5T?4I[6=[^<7e#^9H,b:^gNU]J
THXPdG^L@\g[a)aaAeaD.:.CUR6Yd5?M[0^Y+@WCDI+_3PMG^b>FBU:Y+#G0(UCU
O_^M6-9+dADcFeaCW;IBS/BMX@AbZ)K7Wb]af(LaP.79<H6#NRQ7RCVH)RcOG:Da
<+=)AHP#Je](&fOZ;#M/(ebE=WEe>Lg](&OZ;c.35+5FU3:#>4]/)^44g2W^0)@4
DcV4d&HEa_;^RDI6f]JCBa[=KAO<C38EOGW4]8Ze@GF<F\fU.W#=+S(AYNT9OR\KR$
`endprotected


  /** Transaction that holds ownership of snoop addr channel */
  protected svt_axi_ic_snoop_transaction snoop_addr_chan_owner;

  /** Timer that monitors rack assertion */
  svt_timer rack_timer;

  /** Timer that monitors wack assertion */
  svt_timer wack_timer;
  
  /** Variable that stores the ACWAKEUP accertion transaction count */
  int acwakeup_deassert_count=0;
  
  /** this flag is set when ACWAKEUP is asserted */
  bit active_snoop_addr_chan_drive=0;

  /** Associative array of the send_snoop_addr process indexed by
    * the transaction handle */ 
  // NC gives this error for these declarations (not currently supported)
  // Associative array uses an element data type that is not currently supported [SystemVerilog]
`ifndef INCA
  protected process send_snoop_addr_proc_q [svt_axi_ic_snoop_transaction];

  /** Associative array of the receive_snoop_data process indexed by
    * the transaction handle */ 
  protected process receive_snoop_data_proc_q [svt_axi_ic_snoop_transaction];

  /** Associative array of the receive_snoop_resp process indexed by
    * the transaction handle */ 
  protected process receive_snoop_resp_proc_q[svt_axi_ic_snoop_transaction];
`endif

// ****************************************************************************
  // Local MEMBERS
  // ****************************************************************************
  protected bit suspend_arready = 0;
  protected bit suspend_awready = 0;
  protected bit suspend_wready  = 0;
  protected bit suspend_bvalid  = 0;
  protected bit suspend_rvalid  = 0;
  protected bit suspend_rchunkv = 0;

`ifdef SVT_AXI_QVN_SLV_ENABLE
  /**
    * Token pool to keep tab on number of token issued and available for each VN. 
    *
    * Following QVN Token object queue (one for each Virtual Network) is used for Read Address Channel
    */
  protected qvn_token_pool qvn_read_addr_granted_token_pool_of_vn[int];

  /**
    * Following QVN Token object queue (one for each Virtual Network) is used for Write Address Channel
    */
  protected qvn_token_pool qvn_write_addr_granted_token_pool_of_vn[int];

  /**
    * Following QVN Token object queue (one for each Virtual Network) is used for Write Data Channel
    */
  protected qvn_token_pool qvn_write_data_granted_token_pool_of_vn[int];

  /** Internal queue of active write addr qvn transactions */
  protected svt_axi_qvn_transaction active_qvn_aw_xact_queue[int];

  /** 
    * Semaphore that controls access to the active qvn xact queue. 
    * Any access to the active_qvn_aw_xact_queue should be via this
    * semaphore. This is because there are multiple processes
    * accessing the queue and it is neccessary to have this kind
    * of access control to ensure consistent behaviour
    */
  protected semaphore active_qvn_aw_xact_queue_sema;

  /** Internal queue of active write data qvn transactions */
  protected svt_axi_qvn_transaction active_qvn_w_xact_queue[int];

  /** 
    * Semaphore that controls access to the active qvn xact queue. 
    * Any access to the active_qvn_w_xact_queue should be via this
    * semaphore. This is because there are multiple processes
    * accessing the queue and it is neccessary to have this kind
    * of access control to ensure consistent behaviour
    */
  protected semaphore active_qvn_w_xact_queue_sema;

  /** Internal queue of active read addr qvn transactions */
  protected svt_axi_qvn_transaction active_qvn_ar_xact_queue[int];

  /** 
    * Semaphore that controls access to the active qvn xact queue. 
    * Any access to the active_qvn_ar_xact_queue should be via this
    * semaphore. This is because there are multiple processes
    * accessing the queue and it is neccessary to have this kind
    * of access control to ensure consistent behaviour
    */
  protected semaphore active_qvn_ar_xact_queue_sema;
  
  /**
    * Delay after which the QVN token request is to be granted
    */
  protected int unsigned vawvalidvnx_to_vawready_delay [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  protected int unsigned vwvalidvnx_to_vwready_delay   [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  protected int unsigned varvalidvnx_to_varready_delay [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  /**
    * Counter used to for introducing delay between QVN token request  and grant.
    */
  protected int unsigned vawvalidvnx_to_vawready_delay_counter [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  protected int unsigned vwvalidvnx_to_vwready_delay_counter   [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  protected int unsigned varvalidvnx_to_varready_delay_counter [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  /**
    * Mode to control the assertion of V*READYVNx signal. The mode can be change
    * for every token grant. 
    * 0 - Assert V*READY in responce to assertion of V*VALID for token request 
    * 1 - Assert V*READY before assertion of V*VALID for token request, subjected to token availability
    */  
  protected bit vawready_assertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  protected bit vwready_assertion_mode  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  protected bit varready_assertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
 
  /**
    * Mode to control the de-assertion of V*READYVNx signal. This flage is only 
    * applicable if v*ready_assertion_mode is set to ONE.
    * 0 - Keep V*READY till assertion of V*VALID.  
    * 1 - Deassert V*READY after some time if V*VALID is not asserted. 
    */  
  protected bit vawready_deassertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  protected bit vwready_deassertion_mode  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  protected bit varready_deassertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
   
  protected logic previous_arvalid;
  protected logic previous_arready;
  
  protected logic previous_awvalid;
  protected logic previous_awready;

  protected logic previous_wvalid;
  protected logic previous_wready;

  /**
    * Flage to prevent call to process_qvn_reset() for every clock of reset 
    */  
  protected bit  process_qvn_reset_called;
 
   
`endif
  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new svt_axi_base_slave_common class instance, passing the appropriate argument
   * values to the <b>svt_axi_common</b> parent class.
   *
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter UVM report object used for messaging
   *
   * @param driver Handle to the slave driver
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter, svt_axi_slave driver);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new svt_axi_base_slave_common class instance, passing the appropriate argument
   * values to the <b>svt_axi_common</b> parent class.
   *
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter OVM report object used for messaging
   *
   * @param driver Handle to the slave driver
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter, svt_axi_slave driver);
`else
  /**
   * CONSTRUCTOR: Create a new slave common class instance, passing the appropriate argument
   * values to the <b>svt_axi_common</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_axi_slave xactor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Initializes slave I/F output signals to 0 at 0 simulation time */
  extern virtual task async_init_signals();

  /** Drive default values for slave signals during asynchronous reset **/
  extern virtual task default_signal_values_async_reset(); 
  
  /** Initialize the signals to known values */
  extern virtual task initialize_signals();

  /** Samples the physical pins looking for key events */
  extern virtual task sample();

  /** Samples the reset pin */
  extern virtual task sample_reset();
  /**samples initial reset async*/
   extern virtual task sample_reset_async();
   extern virtual function void detect_initial_reset();

  /** Processes reset  */
  extern virtual task process_initial_reset();

  /** processes reset */
  extern virtual task process_reset();

  /** Performs Reset checks*/
  extern virtual task perform_reset_checks();

  /** Samples the read address channel transaction from the physical pins */
  extern virtual task sample_read_addr_chan_signals(output `SVT_AXI_SLAVE_TRANSACTION_TYPE curr_read_addr_xact);

  /** Samples the write address channel signals */
  extern virtual task sample_write_addr_chan_signals(output `SVT_AXI_SLAVE_TRANSACTION_TYPE curr_write_addr_xact);

  /** Samples the write data channel signals */
  extern virtual task sample_write_data_chan_signals(output `SVT_AXI_SLAVE_TRANSACTION_TYPE curr_write_data_xact,
                                                     input `SVT_AXI_SLAVE_TRANSACTION_TYPE curr_write_addr_xact);

  /** Adds a transaction to the internal queue */
  extern virtual task add_to_slave_active(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Removes transaction xact from the internal queue. */
  extern virtual task remove_from_active(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Removes transaction xact from the internal queue. */
  extern virtual task remove_from_memory_update_queue(svt_axi_transaction xact);
  
  /** Receives write address information */
  extern virtual task receive_write_addr(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Receives write data information */
  extern virtual task receive_write_data(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Sends the BRESP signals on the physical pins */
  extern virtual task send_write_resp(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns the consolidated response for the specified address and control attributes  */
  extern virtual task get_slave_response(ref `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_arvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_awvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_own_awvalid(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_own_wvalid(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_first_data_before_addr_wvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Sends read data */
  extern virtual task send_read_data(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);
`ifdef SVT_ACE5_ENABLE
  /** Sends read chunk data */
  extern virtual task send_read_chunk_data(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Drives the read data channel signals */
  extern virtual task drive_read_data_chunk_signals(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);
`endif
  /** Receive read address information */
  extern virtual task receive_read_addr(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Drives the AWREADY on the physical pins */
  extern virtual task drive_awready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact, output bit was_suspended);

  /** Drives the ARREADY on the physical pins */
  extern virtual task drive_arready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Drives the WREADY on the physical pins */
  extern virtual task drive_wready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Wait for suspended READY on the physical pins */
  extern virtual task wait_for_suspend_ready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact, bit wait_suspend_wready=0, bit wait_suspend_arready=0);

  /** Waits until the transaction is ready to drive ready 
    * signals based on number of outstanding transations */
  extern virtual task get_ready_lock(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact, int calling_task );

  /** Deassert's the ARREADY on the physical pins */
  extern virtual task deassert_arready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact = null);

  /** Toggles ARREADY when read address channel is IDLE */
  extern virtual task toggle_arready_during_idle(svt_axi_transaction xact, output bit is_valid_accepted);

  /** Deassert's the AWREADY on the physical pins */
  extern virtual task deassert_awready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact = null, bit was_suspended=0);

  /** Toggles AWREADY when write address channel is IDLE */
  extern virtual task toggle_awready_during_idle(svt_axi_transaction xact, output bit is_valid_accepted);

  /** Deassert's the WREADY on the physical pins */
  extern virtual task deassert_wready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact = null,int curr_beat = 0);

  /** Toggles WREADY when write data channel is IDLE */
  extern task toggle_wready_during_idle(svt_axi_transaction xact, int curr_beat, output bit is_valid_accepted);

  /** Drives the BRESP on the physical pins */
  extern virtual task drive_write_resp_chan_signals(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Deassert's the BRESP on the physical pins */
  extern virtual task deassert_write_resp_chan_signals();

  /** Waits for bready */
  extern virtual task wait_for_bready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Waits for rready */
  extern virtual task wait_for_rready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Waits for wdata */
  extern virtual task wait_for_wdata(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

/** Waits for awaddr */
  extern virtual task wait_for_awaddr(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Resets the wvalid flag */
  extern virtual function void reset_wvalid_flag();

  /** Resets the awvalid flag */
  extern virtual function void reset_awvalid_flag();

  /** Drives the read data channel signals */
  extern virtual task drive_read_data_chan_signals(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** 
    * Wait for suspended signal from being driven. 
    * Before the driver attempts to drive these signals, it will check if it has been suspended. 
    * If so, it will wait until the suspended signal has been resumed with a call to resume_signal. 
    * This is supported only for valid and ready signals. 
    * It is supported for ready signals only when the corresponding default is low
    * .
    */
  extern virtual task wait_for_suspend_signal_resume(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact, string signal_name="");

  /** Deasserts the read data channel signals */
  extern virtual task deassert_read_data_chan_signals();

  /**
   * If reset happens before the transaction is added to the add_to_active queue
   * the transaction is aborted and written to the analysis port.
   */
  extern virtual task  process_reset_for_new_transaction(svt_axi_transaction xact);

  /** Performs the data and wstrb alignment for data before address  */
  extern virtual function void align_data_and_wstrbs(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Gets access to the read data channel for this transactions*/
  extern virtual task get_read_data_chan_lock(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** 
    * Releases lock of read data channel. Decides which transaction should
    * be the next owner of the read data channel.
    */
  extern virtual task release_read_data_chan_lock(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact = null);
 
  /**
    * Returns the number of beats based on the current
    * interleave and the random_interleave_array
    */
  extern virtual function int get_number_of_slave_transfers(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact, int curr_intrlv);

  /** Gets access to the write response channel */
  extern virtual task get_write_resp_chan_lock(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Releases lock for the write response channel */
  extern virtual task release_write_resp_chan_lock(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact = null);

  /** Advances clock by #num_clocks */
  extern virtual task advance_clock(int num_clocks);

  /** Steps one clock*/
  extern virtual task step_monitor_clock();

  /** Drives the write address channel debug ports on the physical pins */
  extern virtual task drive_write_addr_chan_debug_port(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Drives the write data channel debug ports on the physical pins */
  extern virtual task drive_write_data_chan_debug_port(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Drives the write resp channel debug ports on the physical pins */
  extern virtual task drive_write_resp_chan_debug_port(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Drives the read addr channel debug ports on the physical pins */
  extern virtual task drive_read_addr_chan_debug_port(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Drives the read data channel debug ports on the physical pins */
  extern virtual task drive_read_data_chan_debug_port(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns the number of outstanding transactions. */
  extern virtual function int get_number_of_outstanding_slave_transactions(bit silent = 1, output `SVT_AXI_SLAVE_TRANSACTION_TYPE actvQ[$]);

  /** Waits until any transaction ends */
  extern virtual task wait_for_any_transaction_ended();

  /** Waits until a valid or handshake takes place on any channel*/
  extern virtual task wait_for_bus_activity();

  /*
   * Returns the delay to be executed by the address channel 
   */
  extern virtual function int get_addr_delay(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /*
   * Returns the delay to be executed by the write data channel 
   */
  extern virtual function int get_write_data_delay(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /*
   * Returns the delay to be executed by the write data channel 
   */
  extern virtual function int get_write_resp_delay(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /*
   * Returns the delay to be executed by the read data channel 
   */
  extern virtual function int get_read_data_delay(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Deasserts the ready signals after transaction removal from queue */
  extern virtual task deassert_ready_signals();

  /** 
    * Deasserts the ready signals if another process is not already driving these signals
    * This task is non-blocking. It is called when the queue is full
    */
  extern virtual task try_deassert_ready_signals();

  /** Utility function to construct timers */
  extern virtual function void create_timers();

  /**
    * Creates the transaction inactivity timer
    */
  extern virtual function svt_timer create_xact_inactivity_timer();

  /**
    * Notifies threads running on each transaction that a transaction is obtained from
    * input port.
    */
  extern virtual task notify_slave_new_xact_received_from_input_port(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  // ---------------------------------------------------------------------------
  // SNOOP PROCESSING RELATED METHODS 
  // ---------------------------------------------------------------------------
  /** Adds a new snoop transaction to the queue */
  extern virtual task add_to_ic_snoop_active(svt_axi_ic_snoop_transaction xact);

  /** Drives the snoop addr channel signals */
  extern virtual task toggle_acwakeup_signals_during_idle_snoop_channel();

  /** Removes a snoop transaction from the queue */
  extern virtual task remove_snoop_xact_from_active(svt_axi_ic_snoop_transaction xact);

  /** Sends snoop address */
  extern virtual task send_snoop_addr(svt_axi_ic_snoop_transaction xact);

  /** Receives snoop data */
  extern virtual task receive_snoop_data(svt_axi_ic_snoop_transaction xact);

  /** Receives snoop response */
  extern virtual task receive_snoop_resp(svt_axi_ic_snoop_transaction xact);

  /** Gets the delay associated with snoop addr transfer */
  extern virtual function integer get_snoop_addr_delay(svt_axi_ic_snoop_transaction xact);

  /** Drives the snoop addr channel signals */
  extern virtual task drive_snoop_addr_chan_signals(svt_axi_ic_snoop_transaction xact);

  /** Drives the snoop addr channel signals without AWAKEUP */
  extern virtual task drive_snoop_addr_chan_signals_without_acwakeup(svt_axi_ic_snoop_transaction xact);

  /** Assign the snoop addr acwakeupc assertion cycle to transaction*/
  extern virtual task snoop_addr_wakeup_assertion(svt_axi_ic_snoop_transaction xact);

  /** Waits for the ACREADY signal */
  extern virtual task wait_for_acready(svt_axi_ic_snoop_transaction xact);

  /** Deasserts the snoop addr channel signals */
  extern virtual task deassert_snoop_addr_chan_signals(svt_axi_ic_snoop_transaction xact);

  /** Gets access to the snoop addr channel for a transaction */
  extern virtual task get_snoop_addr_chan_lock(svt_axi_ic_snoop_transaction xact);

  /** Assigns ownership of snoop addr channel to a transaction */
  extern virtual task release_snoop_addr_chan_lock(svt_axi_ic_snoop_transaction xact = null);

  /** Waits for the data phase of a snoop transaction */ 
  extern virtual task wait_for_cdvalid(svt_axi_ic_snoop_transaction xact);

  /** Waits for the response phase of a snoop transaction */ 
  extern virtual task wait_for_crvalid(svt_axi_ic_snoop_transaction xact);

  /** Drives CDREADY */
  extern virtual task drive_cdready(svt_axi_ic_snoop_transaction xact);

  /** Drives CRREADY */
  extern virtual task drive_crready(svt_axi_ic_snoop_transaction xact);

  /** Waits for rack assertion. Times out based on the rack timeout */
  extern virtual task wait_for_rack(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);
  
  /** Waits for wack assertion. Times out based on the wack timeout */
  extern virtual task wait_for_wack(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  extern virtual task process_snoop_resp_channel(ref integer crvalid_to_crready_delay,
                                         ref svt_axi_ic_snoop_transaction curr_snoop_resp_xact);

  extern virtual task process_snoop_data_channel(input svt_axi_ic_snoop_transaction curr_snoop_resp_xact,
                                         ref integer cdvalid_to_cdready_delay,
                                         ref svt_axi_ic_snoop_transaction curr_snoop_data_xact);
`ifdef SVT_AXI_QVN_SLV_ENABLE
  extern virtual task process_qvn_reset();
  extern virtual task pre_allocated_token();
  extern virtual task qvn_drive_token_grant_sig(logic [3:0] vnid, string channel_str, bit val = 0);
 
  extern virtual task assert_qvn_token_grant(logic [3:0] vnid, string channel_str);
  extern virtual task deassert_qvn_token_grant(logic [3:0] vnid, string channel_str);
  extern virtual task reload_qvn_token_config (string channel_str,logic [3:0] vnid);   
   
  extern virtual task process_qvn_token_handshake_signals();
  extern virtual task process_qvn_handshake_for_write_addr_token(logic       observed_vawvalidvnx,
                                                                                                 logic           observed_vawreadyvnx,
                                                                                                 logic [3:0] observed_vawqosvnx,
                                                                                                 logic [3:0] vnid);
  extern virtual task process_qvn_handshake_for_write_data_token(logic       observed_vwvalidvnx,
                                                                                                 logic           observed_vwreadyvnx,
                                                                                                 logic [3:0] vnid);
  extern virtual task process_qvn_handshake_for_read_addr_token(logic       observed_varvalidvnx,
                                                                                                logic           observed_varreadyvnx,
                                                                                                logic [3:0] observed_varqosvnx,
                                                                                                logic [3:0] vnid);

  extern virtual task process_qvn_read_addr_channel (logic [3:0] arvnet_val, bit arbar_bit0, logic [3:0] arqos, logic [`SVT_AXI_MAX_ID_WIDTH - 1:0] arid_val);
  extern virtual task process_qvn_write_addr_channel(logic [3:0] awvnet_val, bit awbar_bit0, logic [3:0] awqos, logic [`SVT_AXI_MAX_ID_WIDTH - 1:0] awid_val);
  extern virtual task process_qvn_write_data_channel(logic [3:0] wvnet_val);

  extern virtual function bit check_token_availability(string channel_str, logic [3:0] vnid);

`endif
  /** Samles the RACK/WACK signals and associateds with transactions */
  extern virtual task sample_ack_signals();

  /** Drives snoop address channel debug port */
  extern virtual task drive_snoop_addr_chan_debug_port(svt_axi_ic_snoop_transaction xact);

  /** Drives snoop data channel debug port */
  extern virtual task drive_snoop_data_chan_debug_port(svt_axi_ic_snoop_transaction xact);

  /** Drives snoop response channel debug port */
  extern virtual task drive_snoop_resp_chan_debug_port(svt_axi_ic_snoop_transaction xact);

  extern virtual function bit is_write_barrier_or_evict(logic [`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] awsnoop, logic [`SVT_AXI_ACE_BARRIER_WIDTH-1:0]  awbar);

`ifdef SVT_ACE5_ENABLE
  extern virtual function bit is_stashonceshared_or_stashonceunique(logic [`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] awsnoop, logic [`SVT_AXI_ACE_BARRIER_WIDTH-1:0]  awbar);
`endif

  /** Checks if there is a snoop to the same cache line addressed by xact */
  extern virtual function void check_snoop_to_same_cache_line(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact, output bit is_snoop_to_same_cache_line);

  /** Perform ACE related checks on read addr channel */
  extern virtual function void perform_read_addr_chan_ace_xact_checks(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Checks if there is a resp to the same cache line addressed by xact */
  extern virtual function void check_resp_to_same_cache_line(svt_axi_ic_snoop_transaction xact, output bit is_resp_to_same_cache_line);

  extern virtual task initialize_ace_signals();
  `ifdef SVT_AXI_QVN_SLV_ENABLE
  extern virtual task initialize_qvn_signals();
  `endif

  /** Processes ACE reset*/
  extern virtual task process_ace_reset();

  /** Samples ACE signals in the read address channel */
  extern virtual task sample_ace_read_addr_chan_signals(
                                ref logic [`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                ref logic [`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
                                ref logic [`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain
                      );

  /** Samples ACE signals in the read address channel */
  extern virtual task sample_ace_write_addr_chan_signals(
                                ref logic [`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop,
                                ref logic [`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar,
                                ref logic [`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_awdomain,
`ifdef SVT_ACE5_ENABLE
                                ref logic[`SVT_AXI_STASH_NID_WIDTH-1:0]observed_stash_nid,
                                ref logic[`SVT_AXI_STASH_LPID_WIDTH-1:0]observed_stash_lpid,
                                ref logic observed_stash_nid_valid,
                                ref logic observed_stash_lpid_valid,
`endif
                                ref logic observed_awunique
                      );

  /** Performs reset checks on ACE signals */
  extern virtual function void perform_master_reset_ace_checks();
  
  /** task to sample parity check signals and calculate respective signal parity values for parity check comparision */
  extern virtual task sample_and_check_parity_check_signal();

  // ---------------------------------------------------------------------------
  // EXCLUSIVE ACCESS RELATED METHODS 
  // ---------------------------------------------------------------------------
  
   /** It configures response for exclusive read transaction */
  extern virtual function void configure_exclusive_read_response(ref `SVT_AXI_SLAVE_TRANSACTION_TYPE excl_resp_xact, 
                                                                 input bit excl_read_error, bit is_overlapped_write=0);
  
  /** It configures response for exclusive write transaction */
  extern virtual function void configure_exclusive_write_response(`SVT_AXI_SLAVE_TRANSACTION_TYPE excl_resp_xact, input bit excl_write_error, string kind="");

  /** Waits for exclusive write transaction after exclusive read*/
  extern virtual task wait_for_exclusive_write(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);


  //*****************************************************
  //            STREAM RELATED METHODS
  //*****************************************************
  /** Main task that controls reception of a data stream */
  extern virtual task receive_data_stream(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);
  /** Samples data stream signals */
  extern virtual task sample_data_stream_signals(output `SVT_AXI_SLAVE_TRANSACTION_TYPE monitored_xact);

  /** Deasserts TREADY */
  extern task deassert_tready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact = null);

  /** Drives TREADY */
  extern task drive_tready(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Waits for tvalid of given transaction */
  extern task wait_for_own_tvalid(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Waits for tvalid a new transaction and returns the corresponding handle */
  extern task wait_for_slave_tvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Performs checks related to locked access */
  extern task check_locked_xact_sequence(`SVT_AXI_SLAVE_TRANSACTION_TYPE curr_locked_xacts[$]);

  /** Updates response parameters when supplied through delayed response port */
  extern virtual task update_delayed_response_parameters(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Copies response parameters from source_xact to dest_xact */
  extern function void copy_delayed_response_parameters(
                                         `SVT_AXI_SLAVE_TRANSACTION_TYPE source_xact,
                                         `SVT_AXI_SLAVE_TRANSACTION_TYPE dest_xact
            );

 /**
   * Checks if the number of outstanding transactions send by the master are not more than the configured max value
   */
  extern virtual function void get_num_outstanding_xacts(output int total_outstanding_xacts, output int num_rd_outstanding_xacts, output int num_wr_outstanding_xacts);

  /** 
    * Returns the number of READ transactions that have started and
    * in active queue 
    */
  extern virtual function int get_num_started_read_xacts();

`ifdef SVT_ACE5_ENABLE
  /** 
    * Returns the number of READ transactions that have started and
    * in active queue 
    */
  extern virtual function int get_num_started_atomic_xacts();
`endif
  
  /** 
    * Returns the number of WRITE transactions that have started and
    * in active queue 
    */
  extern virtual function int get_num_started_write_xacts();
  extern virtual function bit is_in_reset();
  extern virtual task         wait_for_sampled();

  /** 
    * Suspends signal from being driven based on signal_name value. 
    * That is, the signal will be driven low and will wait for a call to resume_signal 
    * before it is driven high.
    * Following are supported values for signal_name
    *   awready     - suspend the signal awready. 
    *   wready      - suspend the signal wready. 
    *   bvalid      - suspend the signal bvalid. 
    *   rvalid      - suspend the signal rvalid.  
    *   arready     - suspend the signal arready. 
    *   all_signals - suspend awready, wready, bvalid, rvalid, arready signals.
    */
  extern virtual task suspend_signal(string signal_name = "");

 /**
   * Gets the handle of the active transaction queue to be used by other components.
   */
 extern virtual function void get_active_transaction_queue_handle(output `SVT_AXI_SLAVE_TRANSACTION_TYPE active_trans_queue[]);
  /**
    * Resumes signal after being suspended based on signal_name value. 
    * That is, the suspended signal will be resumed back and respective valid,ready signals  
    * will be driven high.
    * Following are supported values for signal_name
    *   awready     - resume the signal awready 
    *   wready      - resume the signal wready 
    *   bvalid      - resume the signal bvalid 
    *   rvalid     - resume the signal rvalid  
    *   arready      - resume the signal arready 
    *   all_signals - resume awready, wready, bvalid, rvalid, arready signals. 
    */
  extern virtual task resume_signal(string signal_name = "");

endclass
/** @endcond */

`protected
8GP;JC5IU:3A4F[43<,+G>F+I#a\D>E+XQ#=XRTG;)22)\0.e^OD+)L8a.^=P24\
,g)2UUCX?S\IC#CX&M/2Qb.U_@;_H#@;6#-.6&f.d3UTC<(Ec?V?=Y>[GQZf<G,f
ZRY95K,7KcQEDf2J3<c9X.1FS/#a&(7,&)X-TPRXa?56(ATcHS0RY[>X/,7](3D=
Ua(dJ4OD-Ob_NWeK(1&[FV02G[#B1?Z-#SK,2\8RU13<1B54,Rf\I2;6VL2P>HZ;
;B@J87b=PP-@J6-#DV^3GY:EUM\Wg;a7ZZHc0/O)bL1G4&#B-\04<ZBU.(J@/8A#
9_26F^^>/+=NA6<))9LU84_<PEIX6MDCC@59<LGR8R4:YO\];ZVF8JESe]5_H3KV
[)S]DWKA8Eg(MO1G/.Ngg8CUV_eF6R07R9L+.(aLEXLJ9]cKV)>U#f<UXc>f7[;J
RH#H-eFaJB47I]&\KV)NDX57PMDSHPLSM[IRJ.1#LDfbP,c0A+QM-d&\3SMO=OJZ
.5IGR[d\QcN[NU4Gg[2d<A5Z++1c\D@Y;4]?1=\,>F^9BBV7U3+13V(T#4EF@9(6
\aI>)ZOFGY.E8:,3UAF2WgGF>@;eb57>)g^0@c&GRY7ZER6-(#QK.bVc.LF]+dga
<@e64H]Xd:QD=H+TA+II7,OR^8@]MY9NBLL2=-U&fW3OcRHX5DY<PW_;LYcX2EP=
7;=)=eEVXF\f@BKF-4U^/]QY/e=W]8#U;Cd)[-3(4S<ZQD5=[?P\8ebBedS9)@L@
e#^>Q86&@I^@8)YPWZ7<VHC0[a_.HVNGBV)M?U8ER\Xd0W8)@;1I(JAd&/^^@5=9
+\VJU_PT(2G(Y8aDO)EDORIXdNZLV;;:c)_]d?c=S&V9JXYJY<M9=/dR,dN:],]/
AgQaU;G8_(6BP:<VfM^3VLXW[bce4:Rb?T#N5g3+cc)@.FQO@6#=?PaYM+VHJWOR
:&7;IFT-G^P+OOa)L2]]0&O+B,62a-7^]EB.FV6IUeV0.[E>:Jf5TY>/^<MI^&DS
VWd56]\:UE>DVd+?\1+,:>O_WKR=0Z>JDBS5fY6VW8E)7f8,AYaFeCdF8]EJ@_T6
I6704OcE0F)TPH[LWH&GOBgCgRLWJ6HBZd:gY^a(,#.75@+8<Q((,f)25J);F8-I
#\@c6MKS2eWQ8)cQXGWQY9:QHOOBc5D6_<=TBL>/O3,JR,/:L#O=KOG>fM1_ZE2E
<X@ddCB^C&:#+(7#]A(K_SU23Q>>2OGN+d\bT)L;6=._VQHM?CB6Ib,Q1L;@,2Hb
]J8>0)T.AV8YUTMW:RFE<OTGQ?HTS&?8G.MW_6/7V9cL5]/:T?EP+g29C[/E7\31
XU+T?cafZTDI32WF+&0_8:fcDEa&<ME5,H-\_@+fWe+-)f)PS,e]@abW2U\2>fd8
3gE08)&9fN456>G_XF,867aRZWHK,7Y;A#CG4V&5WJ@?<Q;E)U1dO/]5G1<9V,C,
3KfJ_9/PfEI;PC23DB5-<YU<g.-dCPUKUC/Vc=/D:V0Qc-fV70JWa9g9aZH-V+A2
c_QN@7CAA#G1.53#V/JD[WdNZb<Ig.9^b4@g<f_.Q:[VZ5E]g]#CKI+][gT.9]?J
F/5\-Qcf=-B:VH4Oa/Xf60.>P]6TTBZ=_C0582b2Qb+@JPPWD9CE^fbS7RQ2[UGG
F:FWP4VT4O2:aBH70H)2=5_&[SAcLbd,4;T]I7J-A#D\-EW#LTQAbaN0=/868C)O
XIC3-NXFE:W2(ebd-QR1Xf;<F+Hc>J#[90BbJF6fF.C[ZL9=A3-3M/?g7=T1N<6Q
1J[B>.GS=;3Hb#E4O?6UYI&P.7P5a<:30YZVPX807&^/YY&;GcD+Bd<aHK<UM,g?
_@:<G0BYH)c\P8HFBFP_<cFSVVO^_X<>b9(7\4R^123]K=MO&bVT]:e^8R9<>71b
::X]0&NM.g3T\C0LJPAe(e=KN]+)7#(C_^OaO33cf#=He^T1B9W2GaIZ:-HT3,JJ
9Y_9O7U8RgC@8<MEgCANOO)&I?&Ygfb7R#D4^,U3GeaZgY;f?0Y5+[7239>C,W)d
Z@[8Q.R\E70CF1R62#H5EYA85UEf7II/Rg>O>8:3F<6.fS@0V64Oeg/8fI<)GP87
WS@L)(dH,E:O3=YU)]?2[7^W,KbR@\VMG,H78IRf)OE?T)A-gCebc<CJdNAfVX:P
,X:6CI@Fc3=UX^B\>:ScH\Z:\H?9SY6?ZgA9,P-c;AO-EAIfb(1ZN<+EBCg3b\Z@
1Tc4UB7;C,PKN1Gf8<_f&F@eZ:fb/a\VUE;WGH,b2LM>)654J<Jb5bA0T-O?cIP9
?1N5Y-&.4I&G7MK_&g[UbV<=^_VTE^Ra@KV]UBKNfHHQ8fWC;82EN1SB5@I[(<:Y
(F-#7W]T627#M9K45@Y9f-:-#6BCZWP7LgKG7U_Eg^&#&?_@-H0)(;)GAC5Z14K/
</@801IQ/)SfPP2@1U\ED1?_S(I79NW\_[\9#c2N#LK3.+IV]2Fd,_KL3^=eH;Ib
B(J.5)][(XLNgY)(T-R[a#VJ2ADg/Q<MFV5+LI^(U@FS.dF[,g63,B3#N/R\<8C9
->T;BE24&aMQcUbcG(YA&<f)b_7OQ@-@3cU=T&[X@Gb<>B4Q[cge/6@;MQUWfJ\(
5&)Ce[;g(;)b>FGIWFX(.98A6cFK6TYA1ICGC0)0HbR+;<1W?I<?11+eg_Y_U=Y2
O[fP#>LdJUNS>:>;ES]b25>Y=#:.6\1V,A3/_:gK(Z92@\Ag9]4-H9C?^7HR1QJC
2Y<\1<MA1\-AW;PP@2PA^FVP(S299O>e65Q#<KI@#Z_CNbZTH:Q9BcQgF.OE]X2&
LcG3gcE6WEJ:@QQ6/-?X&@4F/[IVM<-X[2e+9f?8d#[3_Jb@;HcW=@Qc]]9>ORWZ
Af/5=2<J&b>[Oe5EYDT:U4d:fb+@-Pgg(BJVN#E0):-FB7PRdg0/aOM)]HdU&&VF
JAXdKg.KNAD;/M[IZ/[;X.E(0[^D4Y0BI9VS@d@g)K-gOdQ.5F]UKHB(8HX0E#aY
Z?g9&cgcE\/MY9f4=GPA;:<+TA?FUa\SHG#Y78O^9]g.C79d+3<1C6;#dEX0CY7G
aUN;_b</._cd.]1O4;ad:OT?<A5^,:3UK3;LBcAX>76gTUAYW<W(UJ^PQ;,]LOFZ
_2RWeNLF\H4F\-&+b#U8@M:PQHWFY77J->Ja-4U\B8d1<II0a;g]cQ?I3H=3IS<A
FJL;Y_@SH0KbF=3?EPXd9Tb-;>N813B/6O#?=^5,:&1ZY59.Y@@#CU5O[+:YE+[3
4SUC:b6?T3L:(94G&Z\DH+N9QFB@:VVE2^@8>;1e\f(RG?JSK?faA/-N,JFF^V<C
f6#O5L;RC)_c\:MFR@c5Xg7+:VMD&7M-ZK(M[@I=V/IE0A-P1-VB#Z(FQDc_Z)aY
\bFLd=gIAI&X_LBRfc78/_CYZ/PL/6afSbOQQS2+VLMY/_@Jed]C;Z(C-b<GRK<d
:4e3AOd8ETD:1UKEbSa5(/6b]N:/GJ/R::(GJc0Kdaf@BfXGZ+\^Y/_91MRI,eC4
ffaedX&D\B?GI)?V75PK,;U/P7<]4&VPW(NNdTe1dOfMMIWP1(D;AObg+c+1b(IW
1UQ>)L^aQ(L)1-T1WfH?GBNC4&;-RN?L9I1dID48?,U<Zg0aDXf1<3^.J8&0078I
dE1(IK2R<\/LX\6e_+V=2PeOS<Q6Gf2CK+BSaL:K<TNC]Lg#FU_Y_O#fG/<[Z[(?
OIJ@aMaX)@4_VLecG-99[QC+T^1+AS>ATLf^-Q4b3L4]aNEJ6<-SB:4/M\]T^?2&
7IO\U_F0JB9\+C/8e^61>F>8N87/PHK8f6D6CB1AT:g5)]NCHa^>.M[e(XAQ#Iag
GDGgR3&6H.=@TA+^^YW_R<>d:/Y.?YM[89?OHT8bJFXKRGVN)O50.I(+E6TDV4GZ
YQU2&Y\C94Rb0@G-38X&XS,D9c>aSCOgCSGU<_^FO.gFgZcA38M25PgXK/NWD;Oa
UOJ&a8+UOBG#Q<5ddTRZ>J9)(?0QD4QCT-^\V98:AJB01eZcIM^f5B,:GPT;P+UK
MZ+^(X+1gP?FUa=75-WW?];[;UE2H+QDK=789HKZ))dJ#3a<(^D/]8E/+f8g.+W7
\87UgM-066Z06gBZaeGMIS7AD4&aK<\8R[1T7^KU67)I(.1IKU[^10@<\cfLY3W@
:^[KEg.b;_Q^M]IL2?)d6cHVb<)eUF+Z7XN<MRB0[R4CC6AQ(UX9J9\H\P@ZARfM
5^H/acK82YNX8#,bYg],f;YE_K?0RRAIb5/b4\N>eS^C?0@41#]OgZQg,O3R7<]&
EZ&S0VB\26\RaFD._,W=FaWFLa2_R86BgSbVON[UcWcP&6>)612ZZ&TR1M-4-#CR
QJB+]V7\8TCEZ92U79SY-e+GNNeG)4e)RcRdB<+975DD\#e>b.J0If39Vf#g5Qc/
@gZB#_8/GG@86g,_LNM3P8(0+3[fHe<a&7cdCT-.V3Jc][MHF)fCfWN#BO5NQSe-
D7]eE--5-3/G6U20ZRgRN58,NEAOD5&=696RL8LbW9E34R\+#T7f&FR1UEBGJ)6g
RBR<-QN?9;M,3eL>d,QKa^5Z9)8Qf6,E6-d;D(_?d9FOUZUG,Q1.;0D<FGM_]A?[
;BFCJE:.eD#ae-_5[QU.0OFeVYW<2E1ZY-gD./E>Y3BYPOGTM[Ca8[<>d>+G\ER2
OCP/(9FVd(7#;FV1Ff5IcI=..:8B@))MPB>O[b<6=Pa-WN<PL2cN/aWSM01W3=:=
>+aMNBO/KGW,ZL8)U<\eE1(@Q-7]K(+Y(PPRH=R\gGV<B60-[72_F@_OY;/2AQ/e
?L/1K>3(:gW83XKKHJ3SOa(A&Q^E<5IbL-cY0028)\58[X(VF]?ga8\d)/0DPJ0[
<&/BHMGY;MGLYG2:[VHNSV&BN6ff1LU_4^9?1:CQd?)&;_J-dBC6<4J6\NNK\;?)
@<G2Y]H4Wef3EI(YSZ#7bAIRS_&_J5+B#+O?9TV>cBa.4-:P15EYUb.\d&Y37E<S
:R:>VT-CG;.^<X3fYg5WOI9GC/?H/XQeWeCJ#,6PF[7<RK=C=@e@3_7[81(Y\:AM
5.9,/4[.BH_GU8Pc,-\1Cd6^V+NgPDcX+<DM0?&PgM#V+fFUZ0>W^4#L_5WCF:QR
7/&]8(NW5H,Id#&d7>12[VTUR:]g-RMW,JJDIE;P+I6bI\.5\O.\JWZHVbLLd)Ea
T,=BCDMA54HC]>bSL1^HYeT4gP,^/&4NZg6S0L.)1(;\4_/0\6M)XZXa_(C>g^PT
I00-A_7B)I>I22^YFA&7]X+H8;,U/-3X\#CKJOf+5,KG9(I#6g++CbWb,Ff02/^B
M;#OI=YUK)VGc_+_HTfC=8?C1.>g4S5Y?EY2F+^]##BJ^:HeVbK:]J7-Q9C?Z#Y)
4QEUE<Q]EAZ-PR^B7B-:8L:bG)G=^(N&3H]&-c3ST0E=Q,:HWDX1d[QNV91(Y/.b
?VZ.a946eD@8eJ<U^\8DJ>697W#(QMLMN--?C/E/(Vb&XbWC/ND3L<N=YTXL53eH
c4e@XH\R>BI6?TM/<VXD+2)f@gI:]aWM(\K#V,JBY]6g_eN2CD-18R\2Z)=E6_3]
SSRQKL31<b=,OA+<df>H3<8.#5G:3/L&6/Y&P2fF.AaDfQS#0?cX8S4^FQaVeY>_
QeZLbf3f(c@@3f\_NHDbbAN(W^eHcK_cLUe_+D508LPX(+68./D/gRcPIKJ[<LE4
/B0(&E+NOF38(:TF/TJ=2F3[9RJ-DcO?8KDRVB9<0_>^)PW]JbYCgV^@5(HOD]X[
DKEBF^OOL_SB00<eB.8H^N6@A2N^/QXU298+f0M+W-D&HB]15.)V7[GN@I5:cDf5
E0,8dYT1_CfAX,]._.]CSR--#/Z=Q@b._e13Bga7TQ(Ec(bE3CFLD^.=&[VJ;CD2
GaJb0^VB)DY5/PQIGYB7\X>H?KXJCT5ab/F=,e_)7:\b3F+R_YWGDS.=N$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
@55WE/G#b1X(>?US:^UBT#:8Xf\>FDV#1U\V3&fbU\,Q7-]<[b95-(K-O;@YIU9+
[]O-?WUVN3<9aN<^Q(XLC^QAIc#L#P8<?9G4H.J6Y1=-HHDbXS2:1P),2c,4TW]T
)d;.#Y&2DRL)&F93CW3AI&_&#ED(.EF5PXNGgbO7A.b,9WO)TQEKNB8D9XT<WZS#
[D9P525\O>e3Q-@;MJQ=[PK?Z/J4YI@(6WI&df1Q,X3DTf=5>SCH[F^L4dg0\AT@
GA\fGQcea)@]W</#8fVP+IcH9SgaUI8Q/e51eVSF>Z.N;(>5.0+/4e?=gU>DEH,b
Na;b[&2;;/b,aCX0e5G7TPbMH(5+J>f]21_&@?e?OR9+CG,=8);-Cde6(be:(HfP
.+W[<A-@He_7_D8@[;._J8dP:N;Y059H_)F,52gaURN=B<2CVRRMM):M]5W=<#Q3
AF(NcAR?2BQVg?HbFVeaN>JFT+8S6b#SR5<6?.0Y8^S;JE,Y)#&TE;?GGc?e>U)O
[2^e,H_X6UdI4HZR_.CMQ,6>]=516P,dcfa.NNG:.W53cWRKS.[U^A-#S5IFeCbe
/3V55T+d^SZMa9V[(S99^C6(4@DcEe,Y8BGEUNQ,V6MDUN9^6Y[()]I]/XL4LaUI
1,.RT5C7Cf2e:,WE63UE0?-\#&-4eK&,<K#EHT-BL_+MA6\FWK:>&E>O^0gbY1+8
7^eP@gf<G8]eG:9[e2<Yd/A]P=;L)(_R/AB[8O,,DZJ/c-77K(;\SdeSC](M-,CF
dA<XdZXNgb1=fO2:<DF@aY^VF\+U59d<W_<DCY#DWPB,YKX<_H7N+BCF:DA,Of3F
H<[FAOa)ALY<W6QgL^PMfIT=506Yc,M^5e4/BN7N0c7.R)MRg#8SeaANHY.4>-/@
?6bJR1[3911XP8B/)KSfX9f5(W3-M&QP,\:NI[R6(AYa>\JN:b]^YBb<8aR0N7SQ
WgL_+Y8?3ODW37fN9I0eKOGg8:/TKgYSPL60Ja/6)PZ3T#5N=N#J>1gS^_]41-?X
VW_&?K;+M-a_7VWEDM;P\AX8Rc+GIVK/H\A9U=5ge[ggWM60TC/[-BcT559Od05R
[)]A7F@PCO7<BR87U)K/=Sg=P#]VaLT:0&e/&=WRZ?FNd^fCgR7Y(=/d-)^7MW[P
#e,&C\M-f540P/:+8F67#R3FR1e35O>UAa?X\fTA?)TC7CG0X1e8[K)5bG@L&c7:
:=9?8,K2BcLPZD,]NB=g^EdPJV5cWf.O;+(]D4<gT4O;XgWN:MI4J^HZ(^AZH)H+
UZ-RJ&HF,,PHg=>EBZ)TP[g#(<U6YRf:3IF3IfGVd&&2CZ2Z29KM;ZF:2LXT7H.,
/L:Z14d[YD(Z?XC-6BPA;]A?bZ^OXcg+?<OMZTCG5f>-+DS;A&LWFFedZG1)9XU,
gEZG3>DDG5Z:/Se0J)B#VIZ2B9B6@7IV-_Y6EUJ.2N.R,aa1Za&X(S^:NXF.=7:]
/VC+339PUdK5;1XF7&d9cKT\D+J5+(C?CLZISH;E_C2DX91L-d0T>f0-?bSEZX?/
JWK,TK,cZ#5MX.A#VUDO\[5?-I#+Z<:#4#(33(a7ge?0.^NL5a-ab2c@Y^^Gc5/.
\@8a-e9cF8_2N,)bQO<&Ag&fDBSg<^/ZNcKLHaAF\aa2U@dd?^Z0D+IZNa676ACR
ZYL+:CT/3Bd#&->785>39K\4e6.ZG2[gAZ6J()eb)XWTQ&e7CF6B?<8.:AI?CC>d
4&Ba-#UF0fOSUA(dA6:V-f^@ZcWA=@6&[d4G^^F(MSP[J9&<K\-WRfGME0I&R_4C
+b]2\9HC9+0,Z@(V66WZ[:J@Jd88^46=bR@g/:_LWR:(bX[;+(QQ<aFW?f5(N82.
:BNec+=Na4UH98-ZZ#-c[U)-7,/c?;KEBXB/UPbM\5JgB#40<Q,XP(&+Ea_<=/eC
HH06YC6ab0YF^[M\IZ&)#Xd#G7Y1QE=FgEK&A,YfDEIM/7STa^[6>Y15aT,#C_;[
/Y]g).Ue@1W]XNXDF<A&O88cC+X[?1O;dg,:GY2L<UG0Q_8eePH]V?H@3I=GR5>_
X-&HJCZa;YDH2+\E[D(2/R4bA6/a2)QLO>L#HE&1[U9fPTI<B:Ff/63E1M/b:LZF
gO>\aXI-(Ve<Y7,eE;_ALLL[Z[T>R.aS+W8/=bA0^NHN(4DPF9JQ#DLXJaEK6RO(
]A\Z-R<0,=GFG9.Q,P,4d10GK,a=X&;BD(+4)F0C=3VESAc2cHGe[H\XHA\Xbb<4
YBV>a@U\d#G+FTB,fGUBB)<V@Z]bN2J_d6U(>2)\J_R,.N&#VUF4g:S(YDf67?D:
TH+;/-?bU0\Z>INNY1YO:-2/8D6/;LHY#,ENUV,T.&\J?4U_#cKS+7_^>.1]_aa]
RfI&#.@bfV^U;SO3<9DCV<)\3(Q4+6,JY9@^M?bHP/<(LOaLG#HDe9:#@c_139H]
=_])cEO@&#,PD]@[ZcWSbA.[1JOf4MA6=ZIM2^MH[5MPWWWaW+ZBU/KYc349GaWK
VALJTbW[Z=]TP#.e<H]\.@\c0&.\?#CLYV6K?@>U:Ec=E?Z5S#8VGcTKSZLYEO,E
5Ac_7;9;g9]XYcXDE,LGY3_?dD1VdJgfBMDcT/8,AUK49:[YXW;e)U)-OUCa9a)Y
+VQN>DX/G259HW_]6c=)BT#c67I(Qd;9D@SQb.4SYL]_?\_Z:-TIGbPCD8;+MI_U
>N4<Qb11JQZ;FD?7./&]SB8#DSDI=#N2O63Wb=M1T\94EB(.#[H5ee.TI/dT4cCY
IaL7\=/Y)\7,S^Y7]Ld&cVZ4D#&E#S^U+g7_FK8WGPYU]POc6)0-4=MQLU(DB\C:
?.PXHL@gfN?.<GKASKO<9g8d9dY]/BABV4)&@ZD.FKK34CH>H\-\+WW\Ug>?cUYJ
/V/4Mf1Hc81?PK>)&/6O>d1Y[\PQ_fT3T;NJE4DaP,9dDTf&d>bZf(I35^]NKILK
<Wf+@(7.\^20.PYEb34R4[Q5c^?>M:TMAE:PVRMC3@3,YSfX.@04QVBd=YZBe36O
1F:1M1b^0,](41Nd1<HKI5=FE&(ML,KeT1,W;S44gFD-f7c[]9KN74MgRFF+g@F(
1?)\L]F82NSSc/+/#8I=0FKDJb)Qee?a-.OD7D,fO4?UO:SA/6T3fC[,0RE<GaF<
]8a+\4KddNG<P.N>1T=ZV_:OPX0^-GX5?-FLDD+_U[@BY94MERUA_151X)P-4b;b
ZGC_eU@H+/(=4B#Fc5<PY3?[:a82=HJ\eWC,fXSFbcI7[KA;_P&bIDO_3JBQPbGG
UJ:;aQfW^;V5@:LdbG5c((-K88,=0AQ[,6Fc[:(>8f/7WZfg;d6&-45Fa]8>J^\<
5+XM;67#F3&T(BgL5))dA:-..7YGdCNXNf>LQB>GUKdc\E8K\9<1.,5MO\GGPDgW
F7#:<Be#T9AeRU&2N6Xce0(==fLQI<T:eLLUUG/.Q-=K(c1.48LKYAZN40^QffVR
FDS4/(1:,)KQc^JBg+eXd5gCG]D<UB-UXZb79b.UMCM4]fR>BKTBT0bag#))SMY;
KG7e\7<302EN9/^(Q41e5(V)^Y3S)>Qb4dcCJ\6g)5<3?]OB=PCT#(\f&-=f70B&
ea6RgXPRKSN;E5P[J,&V968QJ;FCg3Ua&(77Tc94cZ;F]:DJ8BBO1WSOSF0;AD<T
A;RY(Q2XY6V-E,CXH/6C9De@N7=5T_6J+3<B3Z>Q^]SMcC0H:2[[=C+0PG@aFVDa
G(4adFAf1[#/=;0-2ZDHCFR/GBfBG>;G.ZC5dM59.R^\Y3BIYPb934_G/W(4O^BX
=>2?K>PX?;gfa8cCfPDW1:?b@ALQW99&=0A@g0dDMZN/T\e;X)/eG_7O<SQ>5P9R
4@M8&Z?KMRW7NLI#5ET>6BSaUd-Zb03XXPU6IMP>CFANT9AO_07@U5IIV:-e]DF6
4+I=L-PAU6R^G/1A_7F\U5>O,3<^g+_\JfE.O@+.CZPdfc3CMZ/Q4>A&#X-TDZVD
>(H-8\7Hea^gWJ0,a14,Z-0Ke0DWR+1^42]fJ;)FC7[3Y[DR]:0GAYIEg40Je.L.
d(/,]XXF&?7X?TUgXE^A7?=2[<7#6We0LD2aVE.Z(+\CeJc(7cb09-E.7GB@]a<b
K[3T9UJ6a-LTfP7M5\eDTU&]Ibc/6aEV;_g5VJBgSBdSH=VT:&SOW44:))4U/AC[
9?DVPH<;bc,B;bKaSGS/7L/LWTJG1<:fK#:=W\Sd]CFM<X,aM(<W\&FJ&38Sb>TD
G>>9c5L#@.KSM4[-c9GN(cSb1ST.S?@01=cT^?3&QNHeN_;?2&V(56=^Y^T)7PY1
Kf3d3QMa804D#c>E6U>T86S-:-/AEdX&,.&Yf4/(<#T+88abcg:_bTKHYbH/GWY=
;f3D.),8f(ecOEc7Z364WV4==#\7H_+K#fR[#X3UK-C;,.TGgM1SUK1AP#c-BSHT
A<e8VP-aDEWb.DR8D^1Q_W-6>EcFRIaOSWT3X7)IPYJC-#U+WA5BR[\dB(O>1g8Q
:Ae[5;PH;c+8Y^L1LBdDcDT@E_HBV[R9KQ3E8_.-8>B+CZ(]^_+5.V,O>_de?gX?
f<(EZ9M_L@=SAG2(5(OB<?#KV9.ZJXC#F86WaB0@_4J,T/N(IbYH/<T2TP(,5_7I
O352Q].<9[TF8b[;KBED)<972G)CAPN0SE8Z<G78BC:G<]=f(5;PYCI50]^a-Oae
g#IWfD4CL<<S-/JXBF(G\-\D?U:N7C#L9d\V-Y18fI4KWJ8Y.Y)D\[,53.AQZ@83
&\4c;c.Ke6T6IIT))50CB<W3EXg-&S2R]MNNfgP9B-5+Uc._IF:;6Q/P(fW=-DGP
8b/DYT[OCQPXD(dQ-:NgE./H4T2KBAXC.Qf=e/T#XRSeHeE\b9M;]&P3/D/SO8[#
>QcGN:\K\.8SRARXFd_VA51RgEZ=4BPQQ-RO-+Rc@7<K8gW_K^YEP&V9-B-f/=]g
V&8Z9EHf[224#^)FV3DB9-ARD#B8^7S0cAIe7Z^#<QM.+;^NCcVW[[4IAYVDcZFT
KD&KBdNKY;_&eg:a:fcJZKF;7N?5L(XY;&)T?&ARA<2I6baRW_)c9@KC38..4;-/
5]=LJ-RBHf]+:N>K77;HO.eR(3LZ&3Ze\X:bC2-170](Bd09FM1?\0d<bP.gf4eg
209(3+RTe9G/94_LI5,cU5IfTAYDeMYAH5OHKfAZ7HgN<-,X0(c^PNcf;ALDNQPg
48M]f@&7I91BECY8gG081,Z)0DU\dM]d&/.;Y2L,D+DU#[e/7:O(T4.E^Pbb\;=<
9+G[GUF<A3TQ.FEZNI[\]MAX5&],e^HKBe&fM3Y-\=<WKUR)3L0V<P;J6,/R.<58
<c\Og(c3eJW]00E,WXO.JM?B,F]K7/G0I9e@g)S7P_.ZG4b)HZHUb7d)K2GA#^+.
f6ZQbW;46_3;L:>Q7QHJ7(SRHaX--\@3E^>f][?Oc;HG?Ae+^A_@Fg):MNgDeP+d
3[F,<]VPe^H3D0H]2[Jb18eeS.LO-<X5>:]B5CV(G8A2e,RUBe)8GV]SM5OQK4A?
6=L)QXcVGR](:a[R?Cfa^aeL:K=Z.de3>3\b+bc#ecG3+0OS[^5;8#L9I3[\OLPA
-81LEM@31D0I9/\9>_&(eLK7]NBd5ZVLJFR(-A#,0@b(c3dHW9<JA\?0WXZf<OdW
FL?La:/::;IH6+C.,[C[P1<5\H#JAABN4AD9/9@OJ)R.8J#>:H[,\bgV;<9=_X4\
X+O]5XE3041K7(BZM)MNbBbcVN(&c&Taa:0+6Yg9BEPLXIN8@Q)XN3:LOeIYP)S2
WT[=cWX?Y#TLc97QRaL#QfUT#Y:.U-Q@S1bY<Q1aH>b-OeD:3D94Y;]\c.CTEE;U
TfYP^]49W==,bLc0KK5Eg8?V/BfKf72AR8PWKRKIS-g#),.La\@95/gM-UGI2YQE
d&;0J_@cFZZ(&QV[9Y)HF;&X#B,)g0Z,8U3C:35.F-SA(0GgRb/#V,JH+P4WXU^L
TT1WJDN4?c^&&aN00[?H@CW,F]<]g4IRe:BPKQ(DQ0NM::77cH8d=f\-XQ;5aAZ7
NC&_&WK_P\MTE#g>7N75WBc1,^0bW0.Z,.CU@[.d>S/N.YY/-HTg9B(Od5G_2<Nd
4Q.CB]\O^;#OJBCRY\K=KIIG]#S0989[@,HZ#?d\72=6b>e_^0,d=Ig^J-7GN;fd
))TY:QAKaQXB&AD33OMZQSO2P=]B\DM8P=BH<;28]J-8;6([VSP8Y6e,85c<6#\;
VL-O8>)a<OPfDdF_<6CS2AJ:H9&JX#ZJM2)^U[Ha(bQ,:b_NZC;ZV6O__N_#CQ4d
b++J8c,AVbXfe@D:BQ;D>PU)O+.2]-><-QEEc<(D-QAEZJI@]-:(Y(JPVE?+Pf0B
R36e4FWT_^82gObS4I/<a?I16IV][L0e)EG81ST]WI@7fFGAgQ(;VX6[?8NFJ@U.
E](YZPJF^Sf=,+G6UK5:@,P>>?5cM<[V@,dLH,IY;8;Q^f8??YTcS>#5^fbMU?)1
S49;2S&^#]>=Rf1>2/)0b-cK2:K+e<.,@GdA[VPGJB#S<O/dCfU<C-B38##BYOUg
>a)O\:JSBc6Nb^GP_WXT/R2DDIZI/9bRLD@@a)JfSW#]AU10aZ[NG5Ie(P\4bN]4
8HPPRUacfBMOe-d6&9NbJT(4Q30gFJF5;55\Dc)YUELHf[<0KJA8YTFS/e44+1DE
D1&4JMfF)f+97>//c1N0.L^PF(8aAB];,/cBbEeU@VH>LJHXcfg@^^BM@4.HJEK_
1+X^#aUF=RC7QUBbOYP6IdcfTgV;eB(bI(;,E^JSI(ISaS<L=6(4eQ,UUFP>dQTR
WQ8&g>JN.eb4.8YW/:\NBaJ[)^EB.--SO758W@;OBQK&>WCe17.56->S?gS-OJFM
Q8U5WW+BeL8QcXgTXaIXSAN]-DQ&F\ccD7BM.;G[,VOPM[V=HdL<W-3^<a/D5YM&
K1G9@6N@D>T@#T8#>>1?^NDZ&=7NNZcJ7?LVZ@DKHDY:=XV@&3c4.c?Z9fN2<edO
7OIf(gKNNZ^Wd:Tc\9&1//=T[[ZT6_B8@_0J98KXJG42MW,6?69D+HLKT8GXJ^Q?
#7&B0)W1,Ef\M.9+U>^@Hb/5RZG]0=aPD[WV_d=3J_;^)NLT;O23KV-8g,SBS+eH
_?Bf5-@N+4_Dd@cX+@3-_a4]93A_=M_b>=BAB_(-0#6]7^(Kd\7^:V:XS[?]Z:81
Z_84-X+;Y&A>eU2+fZa-Q<)0f4U[EQgc2Q4BOAP]XgMU77_/)^RI//?ea#OfAaZg
HQ,DE:gbTL50NXWGN8b_+NAE,#L;0QB7,FQ>O0C-B>)2UA?BI=Yb./bH[(P14\\9
&,=f>E)^AIF^RH)Q2QKGfFI4S)dSRgeR:3<5NA[A>.1dB,JWMDY#TdUIf@,\UGH0
_PF9?H86D17JYeHGLD22F3T4C2GO+d]6E;gMIXQJ@>Eg()#BVM=;Y+Td[VQCB+YY
.7f5HdZ]&CK<\#a(I\Nb>0ceB)bH<KDV1JM(Ydbc)=)08R[0cKf1)C92bUQ))U.0
4#Y?f[\6U\_^LMA+]KI>7L2O6D^.-8KK+<@3OeZH(=WVQ6\Gg(JW6Zb]D\>)T/O3
,c=85QKeXMWQ@/@#E82(X(UM,S0B8N2NENgV,+DD,7>6@a]@ZL9F?f:cf#d.WCg[
2M_If,7I[0ZfJK-_IH4(JGE^FaZZS;c5gH4?d;8#&R7U?Tb0<GMa7AW.0M_)H\/4
\R?b(W)6VEG07#D:ER<\\HdNNT[?16d+(04b;[Z0S-Ra80Id538UU&OHLGVNR^_.
P\=0ZL+BF2f\5gJO6PLJ:&@A(@1S;_UfaOZ2FO<@P.FEX@b\b3W#W/<.D,O1[HYO
eBZ,]0?_g0_80YV-DdUI?@f3:V?(VE_XK.>QQ53.#GIFA\NT,RIAI(L4aED.4-5A
0;GO0Q7]/GB=,J)=_IC1MNIZOP@O#W:TSZ5]fLM(<FF\V#Z,+:\MVIY4BB:c2@A-
O0-;##,9U9:;^AU-7+WFR20W9<&HI.]W&&^aG3XOO7INJE1e3AH7@;]U,b;b2eVD
F/DTffT&]&Y97,aCfQ[?L[=g/A),50@0M_f+=O7(&d1gAMeZMTREUMC--e4b_)f6
>LIUS(N?\&BY\#UPVM1/;@D=@,@1SPAO#B3WLF4SKF]+NSX@f:[\)LGg^&S<-X\F
@-6;4<VPFLUbc?.Rdc9YO7PA,L?BSe6V_AR40=<I)>:B+.8<2=U^_d#O&:aUDd(B
EPf\>6JTR^0ISIN(^Fd?Q1Re.ca_HBK-^f#abM\0^-VN^>c=4SfKO14E])TBO7QD
=+5TK4BA8f<L^NKCabcWf0DYQR#E-UcFW94803N?V;JaK3U6>_DY/EJ1R[;:c4=@
#@@=-PWYCC7.C32>f3/V(bJ3ZIK0MFEKEWPeK-YJTNZSc&c-=2+T2@bMa&;+J#QA
=#dI8;&/7Sd8]g)Y8X0bGc0G4KDWYA;<35\cSTJ?3_2AR,,NR9T^0V1XOD@AEC&O
^^8Y+-<NU>IA?9;&J7gXB=Bbb2E>2)-F9#UBK;d)^Q=CGQ;b2?H-0W?04DK:[CJ2
FJ6N@I,F2&S#:eT&-OS8Z(85W-^?[_G<0J;g@G_R4:2A[):TVfE++(#VK23-\(LS
F]C-f[)4IW09CW11K8d@,4JcSZCY56I]FRFXWZ<,=ESAQ-d@H7OgKZ2U]d#=T;LF
GTGSY4FG]+ZA4.659]Zd>HA9_R4b9+,RSH/4US6f2?:XL-U&XR,#NFed<e\e[W9-
0_E?FUZM,5[88<6fc3H2TMb1>FJ)f7EJ2bA5B8:?40dBUVbC-+_-I/#+_2VB3N1G
IAc(:XadQC2FC7[2]2eZ3,IQTG?(]/?KDK.Mg(c9TC6APbARJP9J]3M@]XdLE[]g
3BX?#/=_<713Q?0_R[V0I#;,OHb^g/1[BAVP4I\bX_,K7:0.C@:c;WIf/6FU)WXL
^#:eTC[Z31\+6SF8XC,G+PJ<9dK8L[dF8K^Y759?,[OF[7)3A5dDU4;Z^FK\X7#B
WJ9+G2:Z9MHe0<]ge>93L)B),&,d4\PSBJ<[3a(CUN5MWTA?H&O0],#^C2D,L^:Z
)g?&(K-Q.e0I?ODd/X;]I7ZDFC=S@0M)#-#3FY)Za_(UKXH?LY=<U7P:APcKVFWH
fQ1:W6d]D4J[VDB:b&U=_4&PfM)Rg24N:;<?34]2c7FZII<FYg]5Q]a(>/,G,O>5
g56U2&6J;\GPO+1L]9)Hb#7&Vg&0dNU)QNSH/Fd8FOED\PWD;/[V(5Z3U;_LIMAd
L1^c)/WM9LLU\Y5(UH?==RG,V<JY(&4H0M2)ZXV9UcNL>6B-D?g<5RC4ROI^c99C
7[5LOL(=eMV\X^SE&bc/KM]7]C&#b&OaJ2+cSBPIdXG?XBXWD4Z/5aV_e68c1)ZF
E82<O^d7BM^dN=]5)[F9/4+IaCV:NeLI49071JR<D)gTA9Dd:CM,2_[T&>)P-T=&
2S^2_WcZ67&YNa@Oc1/@YV9#=d8DWW0/TcM4B]RA)D,b7-Aa,Q2GTaA3C#^5T(cc
?\VC@)/>#&KR3:<38[-42O5W?A#AZUB(;BT9,N,@A>V,M5A2Q78^&8KVI78QJE3Q
DA_S/PFWfW@c;\/-=#EUbB-NTBUc&CYXZ3=Va4079JF9f+3d5=1b,Bd>e6\YUHL@
F,3_,Y^/7F_(cg_bZ4.&e,Sf-H=UWI>@(/Tg-#,7)4U_QYaWS42;70ZIUPW&]Y;?
9,&S1Q4XEKL]CRC-KgWWdMN)AUAT-g;N<d0KS4g##c[dK2U1.)5+B\PH3>O:a,W4
/:g81bR+I,PC\\2KBd)5GC@a5<1?EC\Vf(N\_G>Yb)?=AF>.\SIbQL<-]f2I]#<D
8P96FaT#O2N9aFIBUK\\;KMJ.HP5S9PK+EG+3\FQ]+V<FdKHP2X?\[K[>7=7O\B0
G4EI(C[E)QB;Qc-:D86P?I=+(CD#E[6M/UY@O]D]J.P&[d-TRK(F62XMW-X)2TGQ
eZ?/[f/8b5P/3-QR,B^-M/GVC]0N\3@fd49F4P0gM3XNWB49;[+ZWN:((Y@X6OG?
-E2,0gTTQQOfC=:]Q5VeS5bCc_B6;Hef7FId]E^F5#M3Dg)@_>R5V.>9-QA\\7]2
RP#S5-]1GcB7C7W,&T3>2aK=LR@a4<eA^3g>SdOI4QfQPG2=a9,3-3Q]]D;:_HY7
-^].DZ2^a=K3T2&5&-2]>\^/8R_E+L4_gA4CV0#\5Q-MGJVA2/TB]G^FT^C+G6_X
UAZE4-T?9>^ND?--RdCJdf5_&S0b-PS2cGRX7cOUG:.8U_O9DSPE3ZVReQYW^+;B
,5VF;&CTH@<(Jg<^]+B(UaT]OB1+VD?C+GC9dd8ddQ=b0X?GcU1cLf&SU:75XagW
8A2XWI;TNgAG[[)&FSCb8C1>YG-OMZ5OY18bY/J<.eEU&Y<:JGJ+22IEHIHQb^eW
,(3N0=CN2N0][15_VH(GL)^O>+I+GE:YT1,)LaW(Za,?H1)X.-S,.M=\GHCRQ(JR
WU,0BMZ5b]H3NCN,@2g]/L.LL^Gc<.M=AFa1@9C8R<+B/&KF_1#+PAN;LSQ)W=E8
30PXJO_<AJYJP^gH0HZ_5(=F]?-97SG)[,CD]d345NEcF)Z/X^&_(MG/WA&1@1[.
4?4HdGKg0HgUUVU2JVaAbb;1WgXdTZ7fRV6NGQVQJ&]/Z;Z;MZ>.BB[&4O8g#gH6
OE(C]2?cY5.+.gDfC,V1fAc[J1C)ZTO#TDL(W3E#/,0c^;OI6YC47dBUbUYFO\(=
VRH&QR4ZUT^W)7g25)51.g\ff)SQ/-+-9V3N8<)KbAH)N?.6?5))]#5\^\RK8RK;
X5P4\386@K9F.(5TMA)8C]SM57RbTAK6=Z-(VFN:EaB,.TJD)IdNaf9Q/[Y#T\,V
F92J@T&,eAA9W&[e>7SB;B=8A.MGM##M/+,P:eTcbVAZ;eVA2T&J]#cGdH;?FB+W
;aY<)PNRX<6CZ2C(X/c15MF6D(A8/8(cWdHe=[)AC0K=_(:bUC5=PV7>AdDNb#;]
^HBZW0(.U3I0b,66S_@),Pf392>FOXNce-=:bP06[G<Y\>T-9Df2ML,;Q:A5.6).
&TR/L6?@c-Sf7MFL@VgFgI]0[ZdN14KBag>GcPI3KI)/3B?BZ2a0):gU>\fM.#OP
Y0<(@ACYcd>?WL<J&\6;g+ab^/5@:@S)G)RROL-O_EV0./#@P9S_LUd=23BY7K8Z
MIBb]_(J[6b-1?O61YX_DR^b@,9_\dEWUK#_J).2Yfc1;?Z<G\f9Xg:_Me,9UgGa
A/UBVJ&J[W2C(F<F@KDRU5L8H;AJeU9O,Ag6Q@VMV6)-OdR6_^eGJEFS9.C[_#4U
TL5UdFB4L902&dUM(Z381=^#>JE^/D;BEaKJg-a8I[B+T\H1]5Gb8>^LU:FWG&WD
T(^@A>]-Sg(KMG+YF&HJ@HaF=O/Id_D6+M@KA1cE]BTDTKQWML)9^>GgLIg(Zcd#
RZCAEVD8,8cY(:4K;VO6VTW79Y&V3Xe?JNALI>-aGZ:\S&G.J[[J?_B(-T;_E0)U
M#\V5.41AScc@W#&LNRgdf#b:+@_<0Of&R:MB-H5CYKc+62aF\()]^:73U_DR7,8
F8c4[_B<8TP8KB?G,UI\T?SJNH+K5?#e_GLdLM([?/+K&74>^LJZ#R0^1B(/<UT]
Y0_9Z5<-c5V?&UeVYM34EBTKdFaIO&?PHc53#1K7X_\VRJfIDC&R;,=I44[b0^,Y
#F5M_ZM\[Z>1bYA:0XXc13F81?WaJV#M@_]),VQVK/.GATX#-UPZc_IUM_)a;-WB
W]?]Zf5YCbJYa=QL0[UJ&e:ZY?Cc0aOQXJ9f>#QWV1eGK\6]5Tg(:K+\Q1UV;cU-
eN=DJ(OL^bBc0g8X9JQ+NLR6;=70W_DLO9JM\(;b98fY,^EZ;bT36c\TBB6>MRD2
.We@-++>B?[HEaff.8=T+FE21YPQ:N@.bTLFMT>2gI48H/2<2_N]E]LRAFF&314Y
/::?D;7-]M<eF_g_P-4_e,_<=I:OGRe9ESc0Vc7L?AJ[(/f]:IW]>GMCYG9C2QXd
F[@A;7-@+U9Y3QcUF@ffXXM.IAg,,&Q-7NU17WSCEdLK@eQ:XBS26/C65E:,)WVY
Td[GDZ>QF)C+51KZ[967e+>c5\^F9J@d&YPGVC625P^1&_/Af..Z/D_PG12#4+5a
SUbED864VMee4/_Df9g457XIMIX9,Y)c8O^8#W.MA,gagV)0-2C+2gJ1S7[Z\9gG
c#E6_FR5>O?)7\<]S)=1+\_2_4XJ-.f&4M9PPLUdQ/_VDUeZI0/g5Gc7/6H^11(Y
->\E\4D_QQ+<V#\=E97bbN\9^<Uc(:/XN=I8H<N+.==2\g0]@C0RCC7<L:76)U0U
:N#+]#2&9R:d)c#SNNIPXb[bYeN/>DVUU9Y;]3E6^7eVDK+YLG@GE0I<EB.QFZ^\
4]0bQRK&MCQ)?>]&+NU+WQ@^:R6?)T_eQ6LLGB-XaVg;V#52=E]H,<0D;[e1b:YM
FQYFHKe^dXOS[:<VV(,+K6->)<ae8^egAF\1_)+Gg65<H8#0:VK#@d2a_\APF--3
QJgZ6f6C6g1CLS(W1O\gO<&\QK=?AJ(DcQ\<[]UT46Q5Q-)(P:>AfJ[UFT(#T><F
T,fPVRS(GT,9H7H68?S^bR_Y>JULY5ZZ1a_:aa:](Q#5AM+9].Z/F2^F0AWTGA4N
XOV38AM4Vg=LO5LKO?-/;Ie93^]_R6O0K.><^DX14YF(J-&F,FJg3F\57Cb7PAE(
2&(+R/3TM:gV:(?BgBbX+eJES#:U649-;@D85<N.0<S9+.2O,:W]1P7M;EN3O2#<
0/_4WFG6Z.@^f)Fg2/?O]TMe3+0XcGef4UV\beed?;FN-4U8cY8=GR2RJHRaJ_KX
0Jg#b)VD@21_80Z_QK>=<X)bJC6gdW4Da1@UAf@CWU_JZOEXC[CNb9WI]-<PI_Ha
../VG^c>)\N-R7NPXV_XH<W@2T]W783g&<9A:>Vf[F\_gB&FR:cPQG,7E(U@Ma?Z
f[7^.I\I^18YbeH9#+BB5_=<fSL&N\Q.[]A)XJ<.708d49Z.?H_SAD7>F:,Y>;IE
4.&MYYFK#M]=[_g299_(C(=dd6Q9\X6E\P>69+JC?[HX-W69U.K;O<Y5YT]D\?,D
F^TSXJDLQ,++FW^4H9F+EC^SUQGI9C33R6V<R])L3&1JK.IBbgG:dTXIgNCOO54d
VK,(Q5MVFT>K9L\E62#Xf3If=Ce/]<L(8VXMU^:BJUX]-)f4^Oa5_aQ7USg;.-J9
LQB137<ZDbM080,IXV:L-4RMBNQDJ+\87TR\eHc.4C],@_YT4O?@F0LG56cPR<AV
9DHB=K@Ed([Nf;+IOc62RAO^dQ>f)d:f47#dSMD_#H2B=LZJ:2WZ[J-X0^88(2Hf
8?B^A_AC0,TFU^3H+<E<;?1R\=54OE>;JRXM;V=a_/1bRI\bP8eZ0]a6ee5L]?F)
\VQWGH=XX15ddRBEc\Z+8>SeO.@]b1>72LWeM#&HbTMJdL>g6\M:C@A:>UQF[bN1
B_Z,P-@KJ)P:[X<P0&Z#3L0TgU9RaO7[Q[,4aGcYXD1Y==4-Gc>]O+\0V/+V^f+\
^&SU+:/ME\]<[VOE^YQ&4]J[?PST3D9)\)_1b/9,^T;T.@KT9JRTC^;?[ea<Z&\_
[D=A3H_#=gc)XRTCZBOdR+TJGE@fC28X&UF_W.bbJ7EI]3B1D@0d.B/L[e2];&>)
0Y4@EI5@-XQ])1X[)]CR\D\M@=)RN8LB9c<gRJPV2_P-.gUbL&cIb0LXAK8F1ODL
;ACB>:3IQFT0eeN,b?aBEC[HXGa=6e>P^\Z_]<f(D)]bYN3@79VK[Xd>c1EW-56G
B5#B].B#3+G-54TSVS((P.I3QT]P?0RG<^N(;?6Q;<FXC20&Te\=Z4_(SG__X0U?
RE?2D\IcUE>AZ#Ag7#(N>OfF@L=DE&?4Vb^8M#PZNQ5gH^,E:+-6X=/,Y&@/YTV&
^BX,.dZZT5,^;KSBQ;.<0.f2),S@CB,19;GWGLUfG(J/Y>0;-a/>gF/B\Ze(a)Gb
1[<\c]eQJ(MOEUDKCM&fP9N]9fE^NRVRVCHGNdQ\.IbBIg@,NgBMMM2e2YEQ9.^c
WJXV8:6[]/02IFVV#36c=U,.]\K6:X.W69QaX^]WNe8AIe&RU7J^]+(0<L\ZP>M6
c;OQYf[f_U6gWL#c,.-X)7/NP>^4<<IOcIf^cFb6QQO7&cE7A-:WR@&ITaA:eb>6
L.<>BbHUI5)NCLL132QN]=J4Q</Z(fA>7bTEPNT9U(fNXV=<b+1\H[X.=e:2+cMA
KOWR8W3,&-=XE:+dGe(4OV:7[d6-Vd.ebOX5SS&^-?R3ZF2HP+ZAdJV/f0DA,+LA
P&>[^G9A&CUD(9_RI.cLV\5ZATEM9ca>MTE0NM\(]g\#aW^aQOa5:^DGJ-0I?O]f
-1X5fIYaIY);B&;(:I&H;-eK:TcOO\Q3e9@<E&JU)G.97eKA.CCDf8@=c.P;8LU_
B-581)Vd8Qc;f1E[f3T60/?bfC43,dCB)bJB.ZN=)TZNa:a#@)]G<cNVZ>_V-MXA
F8PV+H;-@SU0Y+dg)>4b6R<IT/&bM-N)g2#e_4cJSg_W-9HYdRP.@1?:=+)UD,3A
8)#fMT\.8+?P.PNDfB&M@L7XZ_BHC,D8K4.OETRV@bUb5eY&7LN.,+]C6PD9STB&
Q1NcA;?W(8D[[Je#P^\T0VPX./^d\0YaNYR+=d1MX^H_ES;ATMF(9^AGV<MZYQUF
fJ?(_]Vc,W5E7K-)34&ZGc=e\;C3V-&W3.NF-T,>]S/KAdQ@eJA5=-0=TgRC#BBE
&)^4N@UHK[W>Z>\X]WGd7Z@KXOg)Q3>[<G8I:0DMQdcZc_9:XHa]>G/E.&S)UR?K
JD=0E;_<4;eI=KNePg;L(;&XYV^1W6QbIPNaEcU/\^BDF>6BfAd[G2R.+g:^P<<(
]>>H.L9;F[[U?#G(L>H)MG,D&6gNL:CHf<DFNMB8.2NG^8(L5?2d6A,I93HS19BD
<T,2;(5-bRE+\DLJ(L-,6UQ^fDHB0(WRaJC3&@.+3N].HYcGd+O=W-ZfC,&<_Z_/
:(feW/-NH:/]]K1-=);O,f(GCMD.H+-P\FRG^(f5/@E,3>a2]JdF-LK3&]87H)gf
P,/),>Xa51U6??&)/(G(d2)<b]532N_bBWMb,:_LL21Q>_e3eMO>8CMR#<EKD-gG
9H(R5/Z8=)=SFN/4N.?/-d4SQ#dS;:JL2+4DV)TT0X7#(a<EA6K=219B)<H;RQ:g
AJKg-LC>VHSb1;QW6E7?e@Z21[TSSV-YY[\g1)<Q20f4:]YL2KHA+JI[FeMW>1HL
aSYOfc1\bcP=eR@8e=Q-M9G4e9\&]@aC)>OUG6RFRa[867\E4^O(+.O)/(TZ^G&Y
eJ@-1E89a/.9&S?.FTg\T-S,:A^UHX+)?)M]c-<;GO#]IBUP7<1NU@3QWbS5[P83
+.Z^6UdbQHU=3ELP6fK0@Q;fHdI)+77+6/XCLN2cdW_UTP[5>=V:5WG9(:Q5LG,W
XOY&b8#5)c@N]Da<TTH2?dAINVE\4:?dC#PWEL6\0JXf0:CYBK?\[Oc5+^+Y?V_T
.\FD,NP7:T4H2+CII162RYW?Uf@_1UTXdA4PTbFdKFIJ7WYfgDM&6TO_9AXb4ZY<
aI\8MHaX?8EKfKUKXJGA0-daK,PDe-\bA)P9TeN+E#c:\YP#FHd.gHb#NE#6J)]:
^8ZQS\..BVO)M1Z9WV[VIbGAN>gTCVEFVTYVSFSZ^aXEb;&J\-gcLP+4/#9TLB[.
a#-?[[AT1)gXTZEV=1W9cfa5Z9U9:R)R/JCeQ+=,-3M<QR^[b\&-?I1^I_.4^7T.
CbCRUZDX(#K0EUf=JQEf@)\M+b<MMbTX5O+e]G<CZE/+_OSAN,&F)SE<AZ&:Q,J;
):;)baJAB<L(+S^eg:GD4BK&96^O&0b-AXN7D4ON0&)2^ZKR^7/T3=4fC)_7&?+9
<]8BbKY62XI[\[E#8_:;C<EKaBRI,V^4bT3GY+G1Y1aXaPPP),>4=H]ZVcV>>Ac+
+SCUPcV]+gc_=]YMCAQ<fOX@Z/AL&OQ5]d7a@5d=1UGD4/T3[MUU1-(gPI1FdFH4
?V=9-Ce0<7Z[^e>(NRPKTR)K@e]FP0<)]_gZ-Tg?e1Y,0/UL4XB;?]ba^NXeF7L+
90J_[.].AML=SI^?0T/SOS<3WB?Cd7<U74R@>G8d.D9I>#d4IP=EOSN1acGT/_K7
.9[PD3X#f]gS-BY1Y?_SfEC<NRG_,+)WYX4.-(7#U(JEXBSRLMFX9&WRfRJ6DX:C
G];f-PE]\..\@;;D:f=d,UQP=1;a(3:V)<AA>+1J]U39Z_SQ7Gb.FMbBZ-4<W0Q#
KPY(HYf0VU;X>SHBG(_DLbC+gIVR,0b+\DI^&\L?a-4P&\B#;#LCaG=e&26HYS/M
d=[VdF0KP>QZLLIJP)B_>V&BfC-9M]R[-GN+#\5Rd@3,1@F9-b;N2+\/[L;@SM.>
\,900W?6I18KN@/8(+QYC_B9?-:8IaHB0U0G\0b6_>e[,OB@,H<A2Zd:JD#V/IH3
V@<ZWC>cae/5:_3)f9W?N\OK]7DQUa^33ZPd&2#L1LOXOBLQ6X2&CCX\aUcY-<>Y
3WO/CW?6gYU2:W/FM62X+5@N-VH>,^Z+0NfS7aP6.UNK>b-T.62f@)d[36PF(#Y^
@KWC#Y:P+))_=HKR8<2QX1fV<3R(SL\g9.>a(ffH+.91XMMT\Z/:fH=W:dCBHJ8I
YP.MYJ(b;1c/gJU=,ZfW4;:Ac3[9VN=Y9DgMNB<C>V46^.MZ--@IICFQb;dfEUc=
GP4cA-(0A@Ne?5JSePR(M14:@&B&M>.fBX<L-[)>RGgE>XN6?<UYZO,d#RGc4ZK.
=:&1.1/P;XSI7@Sb@0:BOJT^9<2+XJaYNR-C5717a6]P;.9@+-,a<T#dP3CJfc-g
7(C#HP4(?ad9bH_\5PJPIOW<bc]=0^ZTe;>YPCd#9J&-O[\_642e26JA-7#)?gA4
:GE]2]9=5RD#JQGJb:=Z2J8S?B_:I>a9/,C.1dIHe121FT@9b@-0c:b6JWUN4F+J
C5bd54?-/FR+.2H:X\.LeO2Z<3cd00ID6M;(FLf2/45G,4TKNd<FE,+NFeS#0P8(
YFY^0D#OWH<((2TSB/4]BAKQS@KZ55LH^(HIX^fI06YULH7b?0(UPZ,e^VT9c(d=
L)FNL:a==.7)GHQA+e@2f\7W1]3]R&Y\7Hba-.DHQO\cNED5942S\V8].dMLA6=^
MD@BD<^MQ^=e_@=O\&RD(LV2dIEa(=O#E/[WV:EMBL5)6&2IC.BT;^@6c&ZXO8:Q
1/:]:C@EAK=\>()ZD)ad7J+ScOA:.M(TeO?f2[N)9dEF,Hd,7&Z+CgWA8ZZ_77_^
O);e=5c1gOcILIKWf<\LUO+88U@cdg1VJg#N+IZD;Z1Xgd[9VKWa_M0Y/;K78d,Z
I04;H]3LMa+O1IR)IYF@[Q0EHJTOf7@5TD,EOFEJ:f+c?22_Lb/:K7)O^)+.bRA1
5ISB&F.+M:-70@eD,5;7QI.fQ?FO]P-?SFD,C24,TL\6Q3@faGacS?B_@Ae#ZOBI
.PYf@WHM&HUA&ZM9JRgZ-I#d71cX,MDD4FXaLCGRHMX0UG)KZg+FF3C7=bcO6WTO
NMKa,^)&42@E2KVGZ&-0D=RadK=R+d>WIePM1#D(E7,4PI=+bX5U5d4MCfLT)GGR
S)T/]c_0gFT1[Rf2PW#66Xbg6Q((,ALEb/ddW3aJY=^LS5:e^?LYe5?VP+_;\WZN
_5.ac^W5PUf2#gH>c-=6Y4f?:2WU)/c87W#3?1N,Z6P/11C7&?FYZ3G7\=>HQ8^)
U@[BCT6@A3Ab3e+Z:=(#89S5NVaAJ^R:/caH:,TVYU,[\EeA>U1CdBg1L(V=OF4-
N&+)RZXeBB;TaWK#Bf[2Z+D5b.&\>&5;CI]]cDCJML^14Yb4I3)>=e.PA07R5F,(
1,(//YY[QId.O#JJB-Bd>]C1=g=Z<c5:c:Q.Y1d)9XgW,=F-98.B_J;&>:2?E4IV
f;<dE[CX:+(),),[\fcM+dU1=<NfCCa_^dH1V=G8;_\/VdN>,RM,D9H6VY^CJPXK
Uc6LGRFJNQ;:?^gI3b>b<^DR/WY>?NRMD.Y&N+#YQKO>N><YO=Ec9&XMF=N&S(WD
,#FPedbAN.0G]RCOD+#+KDFMaCY1ZeXf2]YSG,Q:BB1VL<BI)B\,WR[9Z.SgYegZ
GV0NME?0Z7fM7>@-KA.GE#/_6&4>6R@CgVL/PfKMeR0+&<[.-U4<>QS]N3ILA?4M
A+<H=GZ/I5/I]_3d>T]\PDbD[QVRMF:V9@</X,#38c]e]B><TV6F6_dAfU\<R#MO
JAdDO<CZ[)LTIa/dX?1a_S<Ea6N2-BYEEW#BM7<+JeKU:ZZO?DM?3S>0HL(cY<TT
G^LGd,CYLXS)<K>=]UIX>b/,PfAOR6Y@O5d?3Q[@6Ub.NWJ0EHPdM8g+1WPH&B@C
5B6)c#&AU6)?a7\OS@_XRC,K9?19b@HAI-d0Z8Z^NJY^YK0-_V\MUaK[5T9g#A]f
,0-Z=&Q96OE6g=0RQ(./7A4I-A\T>Q-HQ/;5S9BOQ1d12aKNBO)a=OcOc<-P:3RC
6F:De+0GC_7=4S@]_TX:Y@5=J5,FfC[<eE6gWM(c<=F/^_]3.I-[I,ZG0QH;550c
53O<>JM_Y-9@&FfM3FaOf81Ha=gN;OXPP6OXZK/d<Ef>OLD\L#1e<RNZC[03+YYE
.CI)5HW24E?G0dKb@Qd+@[]]?KHbH<e9cde.6+M[_(@#gJa2O1d6IU56D,f=F,5D
I:PV7PS(&+0TO+RM_\IX.C7,5(JR/7I34MC&9:bVdQ>]JJJMM(aTCbE\V9_aH8VT
G-Y=I-8#-\eeY#.ZV&A3dT;.TW(AY/TRP9,W>0^K8>,F1ML8JT[I(GV4>g81R]cG
.FWX<8ZLPWTE8,=G@+[VIf1^/4\KKJ9&LNOgg(Q?\=#.e55;CZZ]V0&8Z:^+>,5f
WONLO(RA5.6UR-UEdY+TCdUX27ZH&>B@+c?9J:UCb1B<(Q8dCd;-T_14c&:8I?c1
]W?e53\Gf,c<W)-ZDO(W-CE8A\f&?[;P;>[()E;GfB]4H(VZdN#U-Q=5Oc)D:VW(
PeSg4EaWP1F;DCT#Ca1,U]1=21bMVRaa(#<AOb#_e:>RD1NW@UJ.#N^fddR3Z[@P
;&N>XgJ0XITbW3V4+95eU-EQ3EIO/UUaf4(><8f)>,.2LZ4G9+J=aE,LQI>BRc7#
e6[/8d]&JJ?6]7J4775<;TO)^[?4Zg[_K^TgH/Ef=3#eT0aH\DTXJI)HU+3&cA]]
Ge[TG^fFP6@^2WU6NY7ZDa=e:.\0.?#N2:U5cb:)I=e6Mg0XI1/P=1+G8VbC?g0D
37N293bf&3@bg&Q[@,Ue@>bAfTaJf:[OREC?MJD.bWFG7?Gf)+SCVgA]DdYaRI-H
\c]^3^WXL-71,7IH=c:P<0K7O9]_(8XU^CX=+Yfbe2a)6XZ686Kc>#SIAe_;O?-T
KF6<1f9fQHU1M@e;)WVW/>Je9)2c682D85-OGba=:M@]Df9&b5@?_FQC5=S:^(gf
CWbU+G8S/#-e[1O,L?DGG#5GF>CYaL#A.HET=<(R7C;^R+e6E/d1KEgbR5&&^&(K
P[>CB3X8V<+U5e(L?XO8:Fd\:EINKZ>\/XDJ094V[0Rg\@Y)1\[K9V<?CHN-YIb^
#2P?UK<E7<EH5eU+^/OT9=RF<+b7ga\_;.<LN:Z14L90]-3&SbeXC,NTT,T[SJCU
I<_D_d(;\)fH4dBcZ[ZOIV0WR9\SH]-@(R2BL.4c97#[G#BLTR3]A=Od-CW_#da@
95b0,ccPIBFCU\3HeES@1Pg==K2KN-VKI;VJPdV5\FZ.^JEM[TE#gA?8,^d.ed_M
PSB/[@C_@#=J_E4-#DRAf?MQ8g#281NFdL^5Y#XX\U0HDeYeHdNCTH2)9OcPf2eC
D+QPe9_@<H;Z&3+Y>E/9+MSB+110;4\ffeZA,ME\D3V5&<8TAIYV5TM4T=A.54+e
X=dTbKHHG;;C4+,,O,&1]:T:(FU+2#4g@:K4(J0P?CZX.SK^g@He/:.4b3YX,RU1
;:+C+WDXcTP;^=GF);GK6&E&IT48b8<KAY(b<F29Yd8EHeF@B_FL<@e?OZ[VgE+I
6?0N>.=aF3aFZRFd6+L;(eUcd-,#9>6#-D8OdHEb;A^U(aWddB.fHWND63d?\a2B
<^U3IdWT(R/I\d>,.=RLQ=[HE]&5C,gXF4dTACP8dAg_@SQdX<RKB/Q4\=PME\2:
dDg;B6NK79Z?,,Nf(_/2\+G)D4#(>YL_REZ7TGCA3#U>9H:^E#.J?]I7g.I?,A:J
ZX6L5c]6PN84T60FZ^]#\Mdc828535R_X+bV1HJUVV\D7O?W@cWA(O?_HA4:KQ..
7_AX^fJ;K]#K8)Z;INe[W[W;.#C:L1V\R87S-_Ve2A_:_2=a[7B_0/G:A9NUM?4B
W+-K@TR(;Mf=<PQFJ7=J\Q,N]-5c/6<gb&4;YZ/NBd@IN2+IL2/_59eIX3gd]gHU
M[Z9ga4g03MgdED/(M&F2dD9W))/.[fS5D(7^e(MMb^M/<1b#^M:8bD/[?_#&SJW
BI:beC;.LR>5&3K8cDTa;/7,OOPAe]I>Cg179UL55Q/:T6=CRdS21E)V2SMQF0=f
&XY(ea5?dP)KT#EI&Z3N1IZ]AgYO86OcRF/?bZgP+=5=ND41-ROR8HEaKCQX.2>Y
X2AX#[e+:Z]MLPY)A1^W[C_>3/H(@.0LVI1PEfHWLQM^5(egWcf8UMfL14C,&:DJ
>?3&)O^?=B;B,#fTOMX]M<A2Tee<+G.)C8Q0(7P76P#(ZL=@UdC8:^D#E>\[eQ-W
-Cge(gY\E]T2(d.VY@A]e,,eC73.g,aB26-[<:b_#D(R/0J:84Y6/1FXX8Lf2R[X
?fc:CO<)1Qd_LCN[Z7cLKgZEOI]NMNbSWYT^:4V?Ea)b_];V6#X=LYMWDfd52K6T
9,=b9d,e\(>,(@U=AC.BKVXB.g.f0?fb8Yg#:cQ.Z+,4+)9,B848^IYCX,<]M;V>
FW3+WF7L4E=We?c2UV[6L]Sbd>_IVO2OU+,VeP(2fTa]7Ta?[CJJ4<IMG8<]9F40
9cW,EM.8@3^J2#Cf^1](NN7REgTH?&6D];DMIB1UM7Z5,[Q5[<TdAc\(DZ)^58P1
>P9&Yb0<b08:Y2PF^BZIDWW?_:_Cd=I(^1gL]QG&b..RXeT[Z[C:MKH6@?<3+;(=
]ba&W-e27K;6]=B=WRPAE>C\CLd_.3Wb9E)GJ39#REdHZRLYN\:1SJ/Q)aaM^#:,
eBQ.1b5-D+B0MPdN_W@C/<OS6KaP^V^.<2Z@^P]f8IR9:X59BL[AH&;1;)XI3.c]
1YVb6-RN?-B8NY7.A&40[];,ZIb&GF:bGI==B>.ScaZ&Z;1FF7#5?]+f2<;V&eQA
(.()RFK79;:?R6APR1_4&gc?]IfWJBV5P<MQF0?/L>9gg_O?SQ@Afb,JZ=K&4G2-
1@8UOa7M6(C.d.f4fILR/]9gAREP,IO17c8L0R5gLR.dEU#VH[Z[8;3<20c87A[(
@QIVCf37#LQ66?,0/./AD8Lb)CTZCP5H+bOeE1M\XMAR@WBP>VE?f^&b4?O7)1GA
XAQA=@XMQ&@\USDS3Uf)bX_Ec#;SLAVMDgROIHVFZ:-.X]@>eWA60(^#TEe^bKC(
OH)Z,Q7N>XO?X]=MI8:1SYf=6[/QYN.N);S+Z7O>;FGeP(M:ZY60#7K0UdD(;@7J
H^5;L2M6N02[=5Y=fA@S-U7.EJW&d)IE5?=^RGK@Ag@2&WFY3W7H&C4W(g>,(?F>
+EDT+c.DA-6bd_#VI\>#2aD7,F</T0):GCZ6L<UD4^QHX:eP;B.C;EXY6aUbBIeJ
DWUfY(67^^=H#e?HGGKA9@J,4GES7XQEYE/2?bY7GfN5NR9\7>,+FQUJcD-Ac:4c
5F&]T_/IU.5?QY1<DGT+?Q?(H8?-T4#f[LSDF+=#42N+4;N#ODKG]3d?ddb:<-Ad
N1ODS?)Ed5IU]WD=YC+X/M2]S;LW82)a)b;H[HB9\1daPeBfOFH;F;Qe(1\2TBU/
PFBCCGS/_f\3[>)a95>BggCa4&T/B5==.FE2DLG3QQ+N(ec4S?15K=cK:.c][e/:
.&<6+Z[.03:SE];1ZC>+4GGJe2Q:.O.7\A,Z[EU1L#>cIGW?E#Q1B7N6G4&bc4Bd
(aBW/5_a#1KMHR>;A6cI0SZTgXAZ=-Ke^,HaKG64G5,#Z<eH5=WUPF7#9Xcg<L?K
e+.N;@,_56A5egSC-.O<J6+;KJ)MM^\;M>/[BE0];aI9)1[-M9X1GA@fZ+PJ?>,O
OWT.YA5-XHZT3XU^?AAbOA[g16.&f=d8079I(8a7,OSDY82gCAg1SH;5U5L&W46#
5DOD=+_2^e8[P-[UR5\28;18S[W0I^>/7[?D=Y&BS.S49UXK#JF#Z=6fN4Z52+YD
^MM;#)?PXV7V@FR/0CWd3dH&G&bL@(f=]S<cg:Nc;4FDdf,-,BAD31,d1.G]E;B5
A^7IH?#.1X8O?eULJa=N?:(WL+_YedMA]\2AVWeEP11=Q(L\JU]U(F<:IW4aPSKa
G5;T597+gID9?L.8EBT&8f:1D-:9N90<HL\5,MXM3FSGWDJXY^c?7\Ed]7f?TdR+
1/,T[d:K;;&&GH<fa06MB9-^@^TeZ>b7#49J8-d7;S<1L61X5V@O3SaECWaD2^-a
7;ZS;S9>Ub/M:-+IMH@:=01R(&-?-PJf=4Y_[>VaO[BD=V#Y2ZJ:N\T-7Fdb?O\(
EW?If_3,c17ALUHS3P,N5]ULET7#<>@CT&FX-HO&_PE;(H7HSKQf:N-O.c@(?8H-
#JfJ.c:ID0J0(Sg8>/gW[Ecg87LM1TF0:T<NLW8)R=@CX?EYd/T[V2=<?9GfUY?V
.eBNJ+ICM+:,(UE66@(Q=0;Q#0EW9V8N))6>.G4eMg)b,X+YG#L?c.X+G082-#<M
F=QR33:LV+CY@U+<Q584O<BY:ZBCEf4:NF[^V9L7\__3_fU/]JSB63Ug^VA:fFXO
-7/eERV8H^O?_>6HKQ-?MQgc8XN,UKJ0;DN@fJb7R=;C53>9&\dL>:Qdg3][9<aY
:HE+fTf[<\4=3;?gC=-X;c8GT:(0CI>A1^EIE;1_Gb6-0&P5a3#GK797e/\T[]O5
(HR].Je&3+;eM53c5KU#JVfZ;0f,aTTYd?]7=47[(06TG2c:+E5MIX#)HBCL96A)
Q-_[[NGGV/[+V1DLTBAeCF5LJWEeX7SJR3V[H/5Mb,R&1gS<WcfEKJX8<EH]]>10
E,4?-N)I3R+:;CV&?4[^E[cQ@g^\/1C2N_a4g5^85VbdKVMV@?@NH2NLY6TY7B_/
R^)0=?B?\32M9:1VPY?NX?Aa6,-_TF2AZN71QE1B&@8/Ke/f+60+g_7+NUSN)_?;
>:Z[AN7^C;5P]f_/S[K)GS[Q@5MW6=@Z?-:IAUIG=Q=?;TCI)O)Db<@F3L7K?ZdT
3eILeW\\]F,T2:V1V[1=+0F(ZcC#LK,eNGY8&ZcHA>LaR;6+5?A>RV12PQY:T2B6
+16;1CO#XS4Bg0E^ZO9G_X=JCc:?9\U]1V[9\+#dL1-2]@=\B7F-M95=8#(1F119
8aRE1K4JE2Y,\ID2UZCB9/P.5VEEB:PN7L;NeCU@QaVe8B?4E[2E_P)SZ&C-=C0N
S2V@H,6bP3YW0.C75Y5B./9<&+[:WK,[C85K,]8K/OO<ND2&AdWaU#KS<MS:E6(d
1Hg)?#0/U.I^<>?S6/RDf3d,d&AO@Z;5[]^(7@/34Zff0e<=b8H?D^f9Z1>OP,7Z
N4gB@E:U:GKK_+=Q4Xga<UE&X?DLME&7b^Q:H(1d88.[,P;f0^8D_[]A=VQ:;KHF
9U,01VP<]/H/X>LL.+1A463&@e_2?cU[9N-QLFV4ST5NC1YI>DBI=EDO.J.:LQEX
7e?=R-AD0c4&C])9DF+DU[(R-A#LAJSZV4QY-KG&Y<Z6#8H;MYcSG]XG(g3<;H5U
T]3ZI\e3@\cF@bd+A^aE><9IW8ZL7<)c\(cNM:TLdcJ0K9:O;3^L=RRg4\f^2LOR
DGF_=VCdRD:IFMKgVUAc[Ta[NE1<7LISO34:38IA4>b\E]RM5.aZdZ3H9T4Lf=dL
@ce?&cN=g/NCJ(+>R3eVJf2.:OXCZZHE.=+KIGE.<C?>(aG0(51V\,MgP6b3K]3A
J5FMeUCTgN9U>>T#EOfCSfbd1B;X,?9cL:P6aS@:157UdB(:0#YM>/JY,TceA)>D
^YUGMX-[646]B94-/>7Q2#OT[C50?G:IIb(Wc\US-?F:MPV(QD<6aYDcegV#H,T7
=UGD/[#Z(-aWPXf3a,Dd/LEVNY>)OC,#R^OBS4)W>P(SW)>^T,Peg0C(5X_P6/(;
H+P_bTP6M1GE+Y-UZJ6HDgf8^2TN+><A/0)2\[a7?a;;=NA/ce_/gAE0P+)\..AO
;8NPN#43b(d4XT1GC_YE(XLdIU[8.M)cHB:8/C@A3L7ecN>5Y^4#7?CJ]GbS5f[M
9La>Q^\D,E4)9[F7J3VNA]P>/5=,I;HFGJN6HT]BaL>P><eg.WTJ-a-L\>YJ&f?/
d&5e:<N8?9TQ&(@=^gQJ[DbC6[:H=RcWVBf:d+<2gNdCgKc5^T\2C78U6?8-SCcc
&^M=OgP4-]QR</C-gOQBdG9e>[B_,0dL.[:TfAP>1RJb+-/#;CYc2bdBO(KagB)g
DHB</:UC+>9_88I,Y:BA3.Z;:IE99e-8\Ha41e2D]UY@/2HR3Y(P3PbM1S&LY?g1
YD_5\B]=J(1We=?L-]K\>_G]=&IGE>Y@2/#[#W/,EXgB.X.#A.,4Ib57F#91Q7Yf
]6Z,=d:6&@>UG-fDV8eV3_\/ca1]_TL8X..8BTg;aJgUNEg-.>TfAf:[2TA3,2;;
RDY[C=A.dU]4/DH#GfY?A_^QS_41M=E=AFH.TYW#^X3N/?ST6E7ZgVZE(H4F/J//
G7NW,DQ@ZaYc(A6PGPaB&PCOK8aJ30B140\MFd_>9=4K;#I6(H&c,C.31O=O74#?
_O3?H^O]PWYPH1/Eg5NEV?70UQ?QGP;EQeV=VD>J,Y-4M]9S>G.#:Y()<bR,CH<1
E..K]Ye?8S7DAAf=a_FC749UIC#7PSG?.KH/#>>Y41aB?d0HDX?OXIg+44bD@QD]
6>9\6TYJ3>cCUc,R)KTS@U88daUdH;EWd;M]BOIS<J\)+1Ae#)_[UM:Y8;,^3+4#
<MB<T:e\H6WF-\T]+(3Vb2Tc(JOb34DM/S:8J<V8MLWMZJZJ82#6MN9&3V[fK4Tg
[@5,T&NB?P6]Q2_egB?HXGb[6EB)R2?[6?#):eY;DQbURY):&[)W7c2S3;@@9<&#
^,.Ee/A5Q\VAXfKZE3?55M6W5P/&d^D(@Z030NST0cF20#_I2906VZ4gR<7I_F_Y
N=POcM0^ERV7Vc:3N=R+/ORgA[AgJOJMHJ=+5f(HeP0PJ6Y>dVQQ1U/eM(5JTT,f
7&)]:VQFJg\120)ATY8NS^H+\6\e?>-9S&.CG&#?QO#bP2T=b\ASTIZ0PfZe)2CS
_7R,WHSM;+30XHD\KN#P,;:N[SdG1Ja_+-<@)db:Nd^^a)G=RX6855.K]AUV?C@9
#e3T0RB?I;beb^RV\X7DeIG5CU1?]eXO^(TYTTNE3.EQ+;2Efaf10644WZb05c;=
=?-PGX4(E-Jf:.V9W0<OH_>M,MG[5g6.NC/+5/NZOe>VJS7)>D8U#6GW_Q3.&-Vf
32g6PFRKU9)/fed=D[5,PNKTG76cDJX1X,cP>]<bJJWG^W;O]@#[F1M>8U<2]b7W
edS)EP_N>PM#97f9)CAJYF4@GIb3Z#M\e-HY]JcgP:L;:IJ?&d-C^,g2M#3IU#S1
Q,#838/;.L<H&SKY).OIU\-bM?70]@/,L,C<ATR[AdG^OWY2@fdJ:4A50M+9>.aB
=^-O?7g\d[50P,,BX+AFQ#J2@10)FfVGW=.R\JA8-W9JT+1FFJ(\=9cI3OVJC)GQ
#]\(AZY<-7+cQ8B]Ag9&#A-4D,^:WYfabB8:cSDLTCa#-,NL_?d3[6Hd+Y\e/e7K
GOZbUBf:CX3PF=ND?C^_cR2JOd/E4B#9eJ+6\6Gd68C\Y#e=^fS<f_.,Q:ag_B8e
[4Rg;B>+(-DA1X5-,:MSQC&1IAe^;=de[Ua.QV[#,-f@.4_D3ST.H&&?SX&E15d<
5OE>KSYgbHYLE&>-,Z1?ZVJ&B=+)E;X)JU9C+=f.4+2V8,O6gV[5g5M[_VP+X383
#B@[_7ebCa)cQI,]1NJ2AaXT]+&);G@GBb+,?I6QLU>59=RK=?MA?FG3@]<?PUFb
XRR5+fY3:2B_0N_D1DI4Y7>fUK;?>Hb4(Xb3)dV[Y<SYXHR=7N3JUTN8[31J.1KJ
#GJE>,bH[;BS0Z@S-&bIf/>FPZ^_/6a@2OBY?>-gYV^OT0J;LFJ@VAON,4XFU]Z&
FMGUQfUed?Ec75D4c,Z(fHfWBZ(R<c@gb\9Ee:8UebBDH3EY7:/aBD5,H3AfWSb,
\;=:SZ62KXa5],=/R(a2?eV9VX(4:0acQ1+I@-R5O?>.V+[+C^.R1@g:b<ZPA)KM
a,.ZOg.N)IK,<9>R4Oc^8=gbdGNZN#(QP3MFCS64&>2BeUL87c^@-&g(OO0Y?I-T
>c6Z6ESV0X.[62D@(1^-L7g0/MJ\4,_8L8\:S0O)7bBR=34/#4_7-(]GX]_8>a3M
DF()]Z5,>,<VIZ.:\.KE[U\XY=F<)(3F?1ZM<KN5EL4^5NQH^Nfe4QDMOW&f\#JW
a5.b0F186XJX#MIfQNBEd/9E[<7>2SG6T#b<U]__1Z/7RZWK?]MgcT60(HWJT)J^
fR:G5H4K]BT)KdO7O70Hg?Z7ZP#+Q)P-]Y6bFTG=6c;e?]]U,<\YPTP5e-8MEJ?e
OJ0IHVTSHHB3@D[QRB-E#g&ddGJLB[Ua=WVD3f21A1XVf]aL,8+HP?aZa]cL]#[a
gLfeaaD&YN8+86PB8?-]0B,PfJW)K:MN-G<&bA1Lf)O&(.<D6)e]_V5T(HbDG4^+
=+7XZJ14VeLV_G@M&Y\bX-PM,WZL6<gC.2YRGT@[]fB?PgP@L-69#<E<\A/9CATe
E8R/M5FPT\D5a<25V0[M4bVAfTbYHb\[CQ3#eR9HC=_/2I;M0?/W=[U:E6f^D=PY
IQTFVC+D/J1J<dAdQH:+:_@J_KRY5?;;-aB\?8LEc@:BDWe-;,9WE(bW.)c5FZ5A
WcXBU7PC;:;>C?6#L+B:1a(UO9<5@=3J@S50,5ZU3RX()+ZOfg,1.?46C-LfUcVZ
^HXaLb/cNUDU/_3VUS,43;^Z#&S;I9F,/8^bSJfg#B)1dW)]@c2dbF^e(,(9Q2(N
>UF)[3bdgH/g@+Ha@^TK^&N7:Kfd:7Z?aZ[?5KB:Xa(RN>D@0<5MH^-I3OK<::,a
0a7_KT6RMXN8EEW(Nb)&3fC4]PRIH<358@I6/g[-<@NR&@bPb;L>RRFMd45d[TWH
0a/78O#dZ<C>;F2EIP85gfA(PVc>CC=/FbNNIDa6C6RcXX;;5U<1bCJ?[@,>AH6<
7VP(S3<)L,SN1e^K=K6OI#[1=S:<-^12G[<]<Y>f_;RaKZR<?dcN76YTU#,bS0WW
3=bX4HR9]>Kd.HL[bA.:?QS/f)GZ(>Q0eIGTZ+7)D8N=IKMOIJD:a5Y<0<&Y6.8T
X^UZUR6]L@5K-gV[#ME8L^:GPegE6>O<MV2M9_H<cAT<>/8ZCJL0;9TYQJ+#E0b?
(X]DFOe?ZJB495..1&]#AO8W(R5D9da=U\eB>]gG);g-,A38SMI5,SJC4O9>>=2d
bX,ZK][;]-\BU7bY#egTCWJ8\=E\_.3H3N7?dNW\Y\[NG;>^PaEaBX[T(fE-2OM:
\I2/;NaM#Vg:YL7N7:.5&)GI4I:/5IJ/=YVdFX160#5L[^O2g=Y(R_c[EGG0)51Q
1bR,G^.AL)V)ZLPEB>94Z-WES[A_M3GF3=d:/REVK?e8+>PQIAgA38OeK30^)Tg/
CBD(-1a5TOYP),T9\0RHb9#EKdNE/0I#UA).cF=f_,Q1GQW.@#.FKWH#.,/)<3BR
D7;#LMc94fYSB)<5-f\6\[TK0?U]2[G^bd>@=\EE=Ge?GU:7PADT,OAdaB=X8If7
B]QL&#6S0<e>IXWFJM>b1)877+HcJQ=Kg9UN.HOV^7b0^CG]VP2:\A2QI-0\bH8F
<(&c2+\?[U(,JURgO/8<eN[:XUfO,+((39,+a@eb2D]&e<OFX^&[<Y#.GV4bg=dX
;P6?\9D]Z0g5Ca<PBF0[BW]Ae91N54f)C^L/222LY2(H5K4WBCaK^0#>EV#0+W6I
WENX0XRL738<KD]N@C0@=HF,:bJ#X(Cc>LMYWN?J()=B=<bENC@.(1<cJ#VgXF88
g-cUPAeePYQLcSd_4=C0F]^2Wa4JBWJO9EXV>N1YB/?NM86T3JB;b,BWGg]2P:BT
a=N>F@]-a<+L1-O4b5SIcKN?cdfKC]9-RS/ELWL>\QLVJ93+UGTYBJM+(3)JH-=H
F>_,2b3bNQf^BNH&16T>OH>Q4G.7Z#I^f<T:TUZOEb/2S1(S_e4K-LbVBJeG@d9.
P1#@/4gd+\-]1JMTS/@8cPW:+C4/^;&cg3@6gZGO_8e3gg3Y]]/b.dE;,/K)c+DQ
.T6.,Q>IV8?RAH+[@)+^g@[c,E)95&7HeOT-QeDW.eYW]M5a]BMNHX(S0-Sba[eQ
IU+O1(e5gUbdK5;FY5(4:PEH#\g&761N]YJ[G/U7.EJ__J4X8+.-SfM7P+A/-OE]
NVXQd]=b=-@=(FeKHGcd.O(^]RLA0T(8b2c?(B+E;<@H_g\)35?fLFLAZPc8,GDI
W?6T2^3Od6R1fI1eR8faCUPXGERdS,C]MJ:DRG78^6XG?<>e3&Z+GG_[Z>Ya(Y;K
J.)WSYDb1)R6NF8\4,K6\,9QRN&NXNS)S;\3F(=)EGb;3T>H-Q_WfYVKZ\D:X,a;
:SYgD8\Bg&&&)Z5,g.Q07?SWN(;)\?#QA+GN@Ja:SG7+A9)=NSKJgFcXR0f?FTW\
65Q2KL8dI:2LGGb32F<N1@18P32FZGg.[61>cNM&8,\8+2P5:Z[\WUJ_1KX1.Eb1
Ic0E?JO?7(EW#UO7LAB,I.Y=<.ObC?5]G+6,@?O2P[ZX:XR:M&:V72PIg#(e(<0#
_1XfS];ULRI>R=Q)Nb((1T1Vb9->38+W+G,=XO8Y;HKJYV2@P\2FBS0KE^<87^dF
A=bQ+eR3\c.64gAD\\&b(-0HMQ8.:dWQc^S.ZV8bVS^EIZIQOfgXMYZdEGGdOTF&
2We<E.YJgOEM7=[:<&EdE0#g:CC45XJ0DHPOfNc1^e#PeEO6?a#aMT>>&4A\Re^R
C]/U@/4EF;:X5J.POJ@2.=aH,_=?E@H@PTWc]d<PQggWFOe.+U]ZZT&;=dbc>^Z=
?M42<WN>WI9DCW]M.(Uag7g:;GLJI]X-3>#b=N+2A_8.dLY0C&GF,BSZFF4I3SAS
ZJKU=\)V1g2J5>1#G0<^I)P(/+ETKGUa;>79e2I[>^-Kef;D,M+eO(&D.[KXEF>a
_f;/,Z:]N-C33<Wg5H5/DGTG>>4,_Hg-DJ/C&ZY/^C>_TKbQ)WT#FU@=>T.aX2(E
S2&P]da78ffJL[@]66E4&?8P8b@Rf8V>KL7b1fCJUF>_6J_Q.EM;2HE,bd\IL_SX
WX4#d)+D0EV?S#:,WA#=3+E(NWSbYES4fP9>[VHK>;V8X\P_GO]C&.#FA;:f_V>1
a4?>M2,&GL<cf5&T-S;3:T.51?FL)f;]NZNa9-&D,IA_)IM50,+Y:@2Y&5V2_.e,
8WCA3Q6CFQ,B=^^[d);^JTaJD][D7=+5M4DLS0.W@<U[WAP>C\]?QOT6)R7I&EQ5
ZBEQC0OC;#AG<ecDH2)1UPAKL-,MH82&;Ye505e@X_-SZ47&(P1;TAY?eA#Jd/J4
\GGJ/,U=G_+FHba^#.f+RKbYW(LSTYC.8V.O;-PFd.2O/c>YX,^9O;(:JUYbP/J-
,F]EZM-#B[bM<3;B0]Pb/gRgJB#(GE2/1cfY_5Y))37^#+8c_,6]+2>aOA,DF]1<
(7H9c8JD=f<g/I=.QC5^1,+,,(=F_HW&>^EGaI@6>@+KZ0LO3g5>VI<(Qd\,?f#a
]0&FJTc,FRJ7.]\4XCO/P.IQRSO^gOU(9cUPH7;G4/gcT+\DK>NB(JF/>QHB0.\5
)1c=#HSf0a1M5>@\NbW+L,Q/ALGUa1SG0TT/J0E7E^Q,[=R9U@JQDW=)b5RM23/:
F2A)@;\2PDOc^Z2FHA&/BXW;_9H7b2Y=V_HK:<RQ#fFcK/(W&U&W+?UW4?b8<UF<
[5N=\C:eOL3)HJ<9GH45>7\X4V9/45QASNOW&4SOSB&XgW+\UC[J85]82aTT8<):
<;,&X-AX^YB#Rc_T-ECI0cE()P]dVO1abadb>UO[YSK2-dJ8d;2U@7=WLaL-)Uc/
7)=f-4H0?AfI?DM)e=e)dS,LZ&\Z1-#]CIGg7IFdf6F=_VC\LMK[44VQY82>#,\G
+2/7A@E(\#:-,5I5Qcd^T>[SBS2(PK@#JfT?;,WZ9^)#8ECR=e15]Z2FRP2AA.Y^
E1WdU([\:0529GPQeT7)_<@SA@QFT@6NQ^eAV@\L]UAX+-Q_,UcF1J=-P0EE&L\]
Q)7:]@ZCa1T4Wf>RZX.?W<M[QIIfcIOE(E4dS>7\MV#->:(bB;eVeb>4(g-WUVQ5
dK_7])#EF/[:18ZXTcBN2#OP4f.JE,LC&4C31R#CEGW_V/60)7VZeSUMeC:edD.9
::3_:5;b)>W41@)5-UQ-@\[^f72H@3;CbMIH&RG[^e-WHAE_\b9HQUg3EfYJ^5e\
DU\:3H616DN<>Db2UWWg8KR3F?I_Y^.7&35GbNU8EMgGU8IAYGLN_Z4a[27KR8:]
MXK(9-P3IVa-AY=>A6Y:<1e/D\-&5:IYaY>]D<_:\^DZ?BAcBc_?6HdRIFRUMTQL
<0NQYc-K-2PN.Z_e+19?;CW9_UMSccgPL1/3Y-(X_S^K1XV3+=VM3.EA:D]BIFaK
-K[1eG>E[@CB[bXV[gV-fBR]OHUXd&G.P2I&/f(_JQG_V/RGbT#Mc831(G1Z9Q^R
;8I^GgeAbC7EFQ94E)&4RI[KV(YPV9CXNJ&-bd=86KE9a/UQ>O2P.4;9?DdZGS&/
.,E<TGcafEV>((aI@:DQGG9=[Y>gF4DVXJ@+&U[Y6N#E2./C][6<7A+5C3L3Jd)H
X</1^77;<f3#d&RC#C<#=^F>P.DdMK\a+d52fd4@bL;GW?[?;(d7\QeZ^,2dG.gf
((g.CUG.L/1bS4_=/]2TV-GRMJWNGLaSAaGY)6Z;J=;@+[_I?ZeGVY^8fD7]a?/B
&;#@/b1_#])_(Jb1ATFaae_2Y^+gK)H1T^PV@D[^RJ+HI^5PZ8,TaJ+6eD2/(a0?
^DFd(7=WFJaZ&/5dS^?MaKW.O:bXUc(d&_Q=b9KJRNJf9+7[6/QBZ:,QVIY<\KZQ
b2P/<H<PbUJ4@_=_C5#.W^.dKF]HK-I,UR)UN(LN8/1e_C_.;W(PaX)@5,bgOWVN
XGJACNG239=938HaUgCE3D8aNQ94=<fb(a4&4-]\:Q9B_,\<Q&O2X+&_e^B-_1g8
ZBaaDeBL6N^9?T5b(;T0Z_17XO_&WY?9G^NK1@f:>P+220YYdD:8Y),d57V0bKgF
a8[S38K1ZRe_]aSN=g2YJ[;>dQ5bC1B7;_[&_5B+g@?85]3[bE(P/.TP67F:[31.
?I-A_M&G[(:T.CZ)L\.>@UgXJc5If+&J7&8(17V<Q[9#fG#,LRB?c.U6@I<T[KA@
T7E0C12+6e,LUZC=FSP:aQS)WUI]^[_3<A:4>\IYMgKD#].c>&2<43N5DYD(TT4(
eP_TcV5B+3Z8\NF?d7K1>aF6fXL7SA=4J/g<GeMI?CQ06>dJEW&=&9W\0P#gGY4,
gF?_J,[ZPH)-9O]B7Y#7R)@;LU<8.1A[=VGQAIf(<Q0RZbPOR/3BM5_aaN\1\eN\
=.4P@RT-\-QWNA[QTKBVMcDgMcE(Y9+QD-/JDKH3f19(#VZ3^-5&/38[dBR>T[7>
+M^EB1FMYFM(<(H23ZR97<J3aCAS/Z[bFXX/=DV=P>^.N<Y)<^KGI]S2[g3)EYB;
3e0_)]7Tc@=84NC77.5W,;3c0H6#B\<T3]Gg?d2=McSXP++8@<Q6Q:f;9^a6<><K
1#;R_8U,eeWXb/f#)[\SgH5H@#]f/<d/P.L_(8.N=I3ba8&[Pf=6e5]B@aAg1ZIE
&:@416H.#^6TXM[c\K+914K+)YYcC.C7W#]I8YKa78MMbO,d<NRb&TO.4dbf#(gb
@?:<WUC>.AQfP5?8Oa=Y?7Yd[cAN9V4(/^N6+b0)_BGeYDbWR#NbIRSEZE/GDf51
VPOf^HLBacL;d[g9d5<f??UCaP&IV+TYDTKOX-=_@QFME^YC.)[dX1dO02b-CCg#
.^>37PM5GMJFN:&3+3UeG^WOI(O8A;>B.Z3Pb@TJ_e0bEU(d<)-OLdIFQE<,3f7R
)4e_>XdFP@&8Q,_T5Y(1H2,#VMENL?bVFM+[O95gcG]U-#RX>TA5>UG,Y+_BB\[I
cU1UN^#_c3Q:cIL7<3QK)[KOARG>I3<aPe^.T)CdF+Y@.70A+(W@U>0;-&)KIEYF
+XcWPX.L[LfG&[GNW1E#<AcU8:XeH\99R<a;K20RU>AGS?&NOfFL;M<]6A_9BLAE
HAG:COARdKOdGI]f@]EHY7T=3\N)#U]-T3<^M_M2-5S5c7ZP-KO1&BGUOeT\L?2Y
ffB<E<Ue<NC8(Z3\GG\&@gAR<^^DH,<NZ>0P_\+QZ6a6[SZIaVIN1=3WKZ>6YO>V
F]PCD?Z(T:Fc.OP5280+;AE3NL_=IP9).c<YE\K#?f_5KE8C,H9_D+?N=@4c:c[N
:T[2N(LZU3QW^\fPd7.a^9f1>IE#E2ZIK2K4&B,T=<M4XX/SBB/bg/ABd8@P6;_#
.ST2.CAZSde-W^(.]/C3O9Ig3BB5,@;>fR=d+DCEUD(beVUgRFOI-)]7H;RWf#S&
R]EG@25^7=V8#9e@X+ATNCQ=K\gK.P)MWNgX4(dGa+0.1PaFaJ>[)QIL=_5]aPX2
+[Ub892VK&.=7&,Bg4.-<WLI>(EFAWH6+_+A?Y9Z8V3U<5_\Y8J8VNF,K\]O,;M_
dATGI4P+VCf+N-I9JT;5KP3R;KR&Odb6b,.X6@1ZPU&dTRM]9ZJ3-MWI9UN_GY(H
\]SSTY?g[6cYJ(S1U:g5S&f\g^)2GY(@[]>J]:bH6F?Q89T]FbRDP@<DSe+NAR\9
>;2N9bWDJFB<6YFS5QfZS\T^A?Gg:/bZ4F@_0^<\Vf&#/_A..=-a0?0aOa]E^^;+
N4>#A2XRBde34>^R@fSR@BdH4.=NSI0Ne?8,&_V?\)MN#I<Tea&c@Na+HJ\9PEa_
>9\HI,bf,:PW>>5KJY(HZJ?>J)>I9_3Z++--/)e_.K,)Fcd2,_9Cd//TZ9W,D8O?
\c=V5\+)fHf7aV.]J+QbL/c;[A^GT_I?@XM_3IQ?9=c&gS<<g-[E935c=W@=[g9b
3EE/8?_.@W#d_e.?::CYC=8_fH&5O/7<7JHW2@Y,C-X<ADA7N)5]2<];FP</eXT6
OQ:WB?9e[5&(MCO(_X_S(/\GI3,f>^_O:45WMd,CgI\b;BaTGa5V7JN#;-O?bf;f
e2&6Va1d6aQD-0G@7TZaX[?dcWVOBJf]PIPE?D?5fcPdI=R?a;7@6X#M>:J7SN>K
LEg3IUA.EF1Q=]V-^KVP\8-C[\72EfeIWGYBT6M9[T;OYV&\0b]T19&CC<Z[:/HQ
3Q.B.XV_@+aP;7CWE3AJ&ebR]R?[8cQA-V5B_:&W.^MB^DM-CPA[eOQ&>AMH/VK/
?G;b#M5_E\==RG_bgX@6ZM,0E-eBQ8+E9JLX;U7_WbIM0Y-2-LO9R;TUd<N1aS?Y
5>a0SU=J;ZLMT-WBR:^S9E;^[XXNXLLD+E?0-/afF@9M[e;OOEf=SP6XGOX)]6eA
/I,O6#5QL/R.)4cO:,aE#SXKZ3<8Pf472SFb_=,f1T1Z_#PfE-21<Qa1@PbIT#DJ
Y7RDV8LTQ>Y@ZcNQ8cWa>BDVNf5HT&,93.)@#9g9C-afcH:3f/TJ8;eDf-OL82&S
V91Kg<.0N1Y]OZ(#.MXL_W8G9gEGW[d9M3cTORM0I(LB[ATa5/4XA,#X[5PLN\\X
WV\N5O8CD+.)<<?X3Yg3TFOcI(3f_gM?bc=7eRIRddEHe1V8)7BB]97KF)_P9AJP
V\[1=0O,,[7AYcbJ=3JD/WVeFU,+EC\>EH3KW@G.GN_UCb:cMba6AAF@H8SJ7LLf
-V8^I7LdEAAK-85cL;bM,N6(:XHV2DUCI)c[(+]BN-[T=d80S&U.d,aEZI[E4F)f
-4U]<7>2A\_0YFcJ<.N#LA/VMI7QRQ+X?JZ89H5I(60(AWA/)IfOCUXdCX+<dI<A
DS>YCHg3.+M3:]T)[d\a=dZ?#H+]3@PPP1G\fgM;ee_ca_4:V&NXTNFNHP+3D2_N
agSS.5_D8d\=Z&+KeZ.IHN;Aa,7&:XN&V4<TF^T8ANL]_-Kb:[I6&Z6F<(\AD8aC
NGSe=#]@:IaURZ>CU\B9UN&[-d5@G=A1/a^2gO;X4C\E(fK-CL@B428c\Zg(c_AD
7Qe+Ed>O>_?:[87#G[K]07#9fa0a-.,8J1;CbI]&K+eO8IYL2PKcMS=8?L\(S[+/
7#^gd\??[bA9ZYWSR08YgJb[IUaJ9\fQc2YP?-\0BE;@NP-O5FfV)V\4C58?(..U
@UC.NASa4Oe,RWNb.RAM@NFDHe/DR=P_aeNIND<6-M<0Z7[I)fg36VRDR70DI[C#
F/R>0&cKWI^;gBS(?.^,6VM5dKd/MdMY>3RUd-KF@g7(AY=)4LXCZd)27SA<RSe\
2b-=AS(HeO/Z+_aRIW:bS31(14e?bbD[[BCP6U2:6^eD\ZH6PFLAbe9SWg@9A_JF
FGNQ).OHGD<9?3^d4#P>]eP-aHX0RM73AA8g)/W?O#4@=+]5MKIR_XXf32Z)D:K-
g&SRR\,.N9RU((<+;</_#4C16OaeD.1=1/3C4(Q^;QLa#<H8B+2Q<.<6Z<b9d:6G
+,=#,QO@Vf3=9LAg5+G2)8C=3a)NX^LB+>;A@@_C[199ZaJ8;:ZH_:-aH)YZ?b\:
]?a-J,CSJW0=4ASB:D4bW[[&R[E2H/c=,e3aVgJ0:[U:XQ,[f\;)-_?7R;R4_V:2
O3ZW)\gcPQ0Ud0SN+5V6VW5_Z/15KU1KK,+(<FfX&51??J.NPT)dXO=2G,WL_4:_
dc67c)c3.a&E>VV76)7Td\[1>VffPL^L95f916YBQPCNB=fdBSR:8faGLFHJ>^WV
OdHe)L6X_+[;cf)Y;(W9&SVdX,C1@1Z?IYAO]G)(^OeIW]GQ2-U/M?^B&=X>7YQ1
2ZG]7ZZF<H3CF@B0aMHOQ.U_5&4IKfS>E8+(ZYO899NY\Va_WfD4=TED[_\V)gHW
0bV<@=aUX?Q<\^e1I-)+30G[\2O5Sa?X#CeJ8b>-.EQEI+WA6e3OQc<.WZ9+^TCX
JCJI15g=X]?3[PGYD(MbBF0J-56O_&YO+N,)VBD;fVA^3gZ\BOGJY?:fSdQ:26M?
\c.6R-AbF>L/9:3=I:NJ2ECQEPVd)dP6.c-#D5FDI)<6Q]/#c^GTPF#OA.X&>N)f
f6@Za)e1R4?1_9c<INQ<GJJ:YT;YPD:-O/GVfTfHc(/ZUL8\-BSMP_Y##/C8>fB4
J=1g\4;)-_-9?X9918&\CXP0IVHbeC:4L0K1L<#Pg;MC^ZUCI)e#5+2a@+6]XIWU
WHCPK^R1:+8\_I)K:&&S3cF+U):3H[-=1(][F2MF,c<61[=P^?[I_F1^:)]4V-J]
Ld[)+5?JAP.#UB,TJBQ@Y\cEWE9,6T,M+a8<O(Pd9R)9dHWQU^88_JLYTD3Gb\OL
T<LZ(^,#B=N#I+@-CY]R/5NF35ZMZZ#&G+)U(0:8-#6Bb)[ee2:/2+L[\A<D\BQG
3=RS^:#^-.YTT5<e/\O0+QLfeC)Qa]gX<+TW1e#+V,1ZQMK?,fVX&4:A:N4[&RKB
,FeM<8A>EDYbTTM-\O_##^EZQ]G,c<)[dC7(c5ZY]UYfI:fBCOW_g?Y_C(4e:3Y0
3cg^EUD2>?(R4aD]g2U&6OX2MV1#.#ZR621SNY3Ca/L.#MU(NR(UGVK0V+OOMO_V
4\,[ef-P7#-DQG@ND#T@[fCd;5KdTUYCda]HY<-,4PX4XMLDDXP?T=8^2D34f399
:0F;_\.=fRB)B[ReC\aIPcEd]=c#<FA,CDZ2D>^BO7b0c.^S=4(]S;<J(J0C@>,a
/0b9/D/8D:))g8#K0V5b3#@<WV->gDTB\@V>7]W=OaK2c7PIff&]OH^3S26=DeMb
g];ANB^<\T,2eN23&.XFEM4^+d;9=W=D#CL<],=[^)AS];FP@2gS&^5)@c#6GF8.
Hb;.B030R>H2=,9:>IO3SR53^^=XDed>TdA&5WWUg;fGHP<VD6NF)12AK.W\M?cT
FK2;))E.@a<],H,OJYHA6#a;b>@W\242U\N_3?eX.=eJ0RLeV_/D56:M+BX;IG&J
_<#1Y_0O>AH:D[Ee62FeHCZ//G9O(GZZQ&?5;+JMOd<KG<EgCXD>.,JOKN2PLZA6
Gc6B7K\2S[NaNYgU[&D^/@ZbD34;X&SddAaZg&M+SOO(5?RTM_bFVT8Z:53K/bf2
1>-Mf>;f-P_VJ:6TTEB/MI8RS]O)H,+Xb,U)bc[^T)&J:d1CTBFS0G1<1.d_?:^D
4ZJSb(fL7N<d+=bFZ/U(#G613X.CS;<->S?e>CH3a0LC6L4M-8^+bd/\K7dVORU]
>?[aLW_Z2I>+Z+GdeHJQ.]^+A.<QPGDQ)=]I,e,ed2#e5Lc-5S?6af=G95@T5ce/
A2U&JO8L5\HP,FWJ.Ng_=a<b/)#)RTV/.7N)V--Sf<L5,QFFFVD=C,9PV7LA0=0E
T14@&S2RC\:&;,E.8e9Y8XW6A;^eGfKZ/IH]7Z,e@+1cVfVDEF;C_]K,DCD4;)5@
8>JVB(I1\Q@f0,)LQ<2WHZ9]eO2.Y,&RANYFKPCJ2\R-R<(<\<9O[,6P0K^&ae\Q
B@9fbR]QC8EfS#7?V1_(>F[c5\/6UeaT7;(e0F&PdHd/>917HdUa(.\+4G2,+7(X
)Z@:d1W2>93^>5HND1,ZYCd0S_XK[Yd#NPECc+_:aaUc1MUg0;ad7a>B++APM0&U
YBEXBd6UXVY>6e:,;D4@^)N2U0f,C@?[gW?155Z\1<gI2/C?5]:WW;/,<,/e)c)-
D&O9/@NfS@5WXfFfNS&JbcB0N8L)10B4?S^?g?U@FDHZb&Y/(FH)M50AI];P>[A#
K_b>&2MGLc<>YB@XH9#&S.R]99fA-D+?6LL,@+CD6,.\LELQ,F_#GO&])cFE:30Y
CEdTF4D5)^<H+_R:^F^<OBAB@TLBeF<DX0BM@VcQ,+,,d#.][ZCbLg_6,&]GKYE+
@-V(cS;J=[TSV@Y\<W8-JTe(H8Z(7C)96#]0G>C+@a)PVZH-P._2b,;YKQ[)\gMW
_<V?1G5V?+^^KHQ:eg28AdGKeIe)BRP,c8C(TCWf.7MUgbEf8NWJD@cOY8.fQdOI
&g/TQ^;K_3M8N:d0CB:.9PaDG]eb-65O).XQC=3f7>15JONA/C>X\HWe[YOBa/bK
b2eVTX@aV\Fa]a4Vfa0U=d<P?W<;AR_M-TN7T&&gM7U05<)/M+3G_91G4(1TPS1F
M^H<GS2##\C&JK7:L\:_H_--Qg-^XC/:;A+<SV9TNg./\31ZJIT@L^/>Bde.;dB+
M&\H975aT=_SDY[CXf+Pg48P9D4?Y=OGC(ZdL+8MBRb?VXT97a?0FCS6SdegE?DT
UOVeJc\-P^(2ZBMJ[EBC(G5e:\3]PT.+Pa65#d;g@;2G1Z^aS6Gca(OabgOXA1UJ
71c=[HD?FM5GeJ2\XI]4D9L7F@BV6,P7aSa\:UU&c[df9TIWDJ^?]R\HOSVE-3U&
-BTcJ,(JSU_VAJ^4G5_&O+,\T_C[73d(2TM6:ZGSMWS4/#T9f:,--6:1;Y+e3QB0
N]9+,XI>+J.BD&G#:W,>\16.K#LS^OTWPR>@WH2,c50N2J;3f?7@WPc=T&@dG.X7
E.c#PR,:S,G?8+-f5(@eW-Ee,W)aA8J-+D9N;V=dQ,AYS5.3-+O4X?+Yg8(6N<;)
,_WGV67:3R?EVR.8,GW.AaVf;f>B3OUB100UFZOd1b+D<_.14N+gY-^7OH=d1XQ(
]5;3a?C?-VD:RBF=0U>_J/Pca0+_BA3I8,Te+g(:IfE7gZ9=G+X[1TQ9HWOaO.K[
:XF/78E[1IN4#X:I6NT52]a3\a2a>d@+AF#9DC0dD2?G):+8O[&;K4X#1a;M94E.
Z>H@RgaD:c3O#>4bM?X&/MAP&LAbP=]STR/JC5SJ+HDOb/b\+NT\48V/7R9\J1[:
H-_bLU_K15^C>ZTKD:gJK75@[GbG^X:TgB>fe&#D&I83:6ga0N&DR(/HQ&)M1FU(
+1\5_,V[cZ-T&,FT1/ReKC&\\TUW-M0=YM;>G>a))QaW3ga.PMWDC3Xd#8:Na(g5
=V(?.6?T_AGD83[Z8F)1]cb9Ig#SgW/V2N9Z]-MWXEGF^AH,f5fc@3&2\V9(+R<[
g_8[cg6-HDD-#BEMLXOGDUYC&7UGB6a@82\bUB04PQb?MDcNR<]+Q(A.@-B_N)V;
^2+]8-X.CS2>LA.Y]#<-XZ:XZ2=d&[8cHLG5<gS3-XHe^7.QWEgRX[WEa1/SXCO?
eJT=#c4_]aRM8O1C-9Wf.@)IFU;9E1XU5.)3de?=LRRRS,OR2#9<M.[@30fCC-ER
M]W,&16COUA<]=8&K^d(]51)/VOZD/d?SLe4SB#gIMcY6ReTJDg9JX&0.CEI.QbV
XBcc6)YAP,F)JR=TNSW9)5gYNS9dA6PEE>eD/+F>MaZTAZD-Q3?F1U)LCHY<G5=e
>Xb=V:=-\JBK[-bQI1.&HNFfeH9d99[Q_3_3M/aDBH9NFXA;:U/E:F:HI&I1F8N[
>GY@NE7TcGB;E3<:<(\S0@:O>T4dXU^Y#S5KcaTa<eB:c(K8F_b@0JFZbK)GbI=[
]7^U&d)4[.Z8LP0:4G@.QfQ/ND^<A72gR^/S&c8/>Y=H)<?VMbIC/G5I#.?O/JBH
I6M[NOO]:4aY[aT1&-;FK&^W9E@8VCQ\=-IMMU[[,-BP&E\SK+;M0#8SMW.gZ46K
f838G-C&R6846#2J^KKDVN:9)3V?2I52e,bO8./bE/:gZ:E,9Q8IEdB\H_f9cH12
NG_6(+@8G1RR(#7])2_GQRNZH2/^\@&G1>d.W&d+SHEeCTQ;M_IZ1I\CG>IY]d-b
4]-VM/I^1)+P,DFcG6)DF8aY9:@G.9gPD;:[T#d6CIB@NIHM80\RG/I^Pe0SNPf\
?)&WUR<K]g]aALf;XAR@e4La&&4C9C33RIV9AC\,0>O#K3SLW)F(^9@7F9-I3>ZU
f]c;eNB\=ODDcfUW3W^LS[@:^9:^(;__Ma7CX#GNBN\J?1,/M@2TQX14N24SZf1>
7H.7&]EPC=&#ZP\;EbRGWb0cJ_dV/7DM-_KAV9Rce.6F#^B<W=851D<7GG^@-H)+
<;BG</#_H,0c30I5#dPDB,BPRT:]Z/c:(gCc9bc779-FN=)-Q_X#:I#N<6?95=,c
BWAY+COB@D<a[WZePHR&cS&9A&\GY0/.4\^WL&KIcA4C9^-GB?KKZVc/<^(R\\7#
XCONR]_M0)=gdeKCF<#GYJ+2V4@Q+-F<@11R63&2N1b25f;03.c5S@c/BSRA#KGM
3,RbM2.aF0N<D:f2F(J>5D0^3C^fEOJ^Bd12JBB855cP:J\KS(N]5J@9><^\b)aT
^9Z03],_dd,2[>Qaf1J1ac,[\bY^:7_WMN,)dNaLR/S#^-9^Jg=d1gQ7]-3LeSFO
GQ<4e+1,,Q_/#175Z?X,f:-gP/_L@<#9Td.3=2J&4:.47Qd5T=c6KJ;^2@f[Wb8/
4d[;2C)TG=.95>6ZAMWC8)G>RQ(O0S,RYDWX0CL.];@W5YA&3_LPEOM6T&[JG/Ra
DW7B/Q)[B<31d<ef;9/?)RBSR25_2G;c4?L35NUDF.4e2QJEeP0CP-K;fH-E6B)W
+5K9F)[Y]U6,4;#PV?H9UQH_+?AFa<[VPg\<+>JJ7U:DfE+WEY=2^#-X6a#R:M50
8NJR@[C3aZ,AVQ.4O].;b@>0a14N:#OLB(&/?gfb-K@VM.^42SXb0UA3QHPB;I@4
TA)2[J?=1183fCZe#Cc2WV1\HD#:f[3-I\1,@Q#XVP?G@/+Z[#<WC0,1e31bBgJR
6?SR]DZ:/_;?8@2bb<49,RdGLGXWc2UGeC0KQG^@c6VGLf)OT)G7Hb+dA+gW6_EQ
9F01J+f;L>8?(00[XM@7^#>&N6158;<K3Ya-;^]DeYP#^.[O;5&HNS/I1MA<U:Qc
6V^X#VaO(c&(fU=H_XU9+::Y/),ag8Z^-LG487V@3?4)5YaG)Y\Z])#8J?ce?:_+
G62[0OV[53CYd,>M0+Ob2<P8<+TZ]3CPWZN9c@F4\T9?RJSM8a\7N8]0&ad]9)4@
O+\?c)O@,\W47KLNY?\aUJ,<8>6WJ;BZ17Ra460C8UFa))VYd&PQ+^ea^KT-R[c)
FWDMa>05U0C-88;9I)[d_@Q^>GRX#Y#B)NDg:I+2fZB)?DS?Qa(44;2JceR)P<SQ
MAX((a-U,WTJQA58HFMUe-c;7b3c>BA-<M6BGI,C[FMP=7Pc]]1b7_#(B4N=LQ1M
Rf0IQJ&U5R[+P7/X\,HF9G9Pa^5/NS^BCC>0gM.#/I(a4W/X;Z[0E(Zfg\QHLa&X
>0P@FG\TS1+YRR@?2145cA1B[Ifec38VQI37>M176A^AV9<DV0-f2WB=)]_F#4+]
^5G15>b@9@RHc0.&b=[=X>3@<N57J@EYX8cfI>FaRQ\0CSUWe]RZ+fL[cB;6]45@
_ICG6.XV8G9,>E#J3A-@\-(0[B<EUe_0Hec?)AVO0gE@f+UXMSa6g6HUTHS0<f?)
Qg?&8Ig25:N@@:^+fG-W3e[GbR>X^(eDY:ZB)7#d+:O2AU,If9:FIJ-GH5.bY4a@
F?(?)C9J/VY=^P3c0g?Sc;.3+G43G;N1&-;86VM/8gdHAc9T5C[Q9Jb_dR[.O:b7
L]R-1GLAD<M9,9JH5E9FQ:c_=5^@.4g4Jb#Ka1N4e:^)>WIK9NaZ@PfMggVF^QKA
P^CJ4P\M8\:2CedT<1CLaG>0-2M:(.dQ0.,VK.FZ#1,+@5c>3<OSaB]f1QRY>Qc<
X56(X\bVd5&5._>N?,P_ACWF98U[GMg=4EgMNHC20#0[3TPC8.0+E9ACXD_<B+W@
?;_/7Y3XJaf(+E8H5e[&>0C\Mf[[UJ_EYIg[cZPR#JLVW=UaG,L9\Kc;6C[RVUA.
\=f2:60ZCP4(>CQcfX6g3Mc,\(ES72+3T3GL9):4_<=F0R[-;7PO8AL,2PXg4DAS
@SF@b1@9[SY\]4ge0]_?NV>d/a1QKA_Df-N;EH)/IM\U=?Z=a(#af0NJa_-EVLPf
I-G^HHaT/)YQSCd\3-7GY2,3R+fYMH5B248;;-@.bb,[VM(cH92O:Na8,H<C3H_C
2g\Y?S7JUS1/@OCWA_#0b8OW=:C=0;I(1L,11R=W])a:Q&#2;a]DTQF0?>/f\U2W
M9PNE6GD3;/ETgF2\aRS&<6W6CL(EHg/N5X6-7^AeS[T9L_LDLN\2-W_LAQ,CS&@
.=1]470.F8/a&EO2/&(QGT4<:M:cg:,B_+6c=g8<RZQV_4HG[SM^;Z6[I0ZL[U)3
[DGI=\994ZTW58<Qa6A2XbS)NGEMZCd<2VYL3AVR;K/P8G80cUSPW-aF7D6[:#V7
KM1?&_4VTG)N22d2/8#OF=P@,.SJ;e[LcP@/cWL1ZWZH-=:(9958;U:(6WdUWebB
-PcSbR8K9&^f,L/O5<:9865URbT/V[\ARF5KgY;Ca#C0EYNU63Z2A<a\9-[LeK0R
(A8X<ND72OQ\^,&>OLTMP0RJDP<d\_gQgag:;;4eF7H[CKV8EUVXT<2<?GW(Z/7a
#V;8K6+N&D&VE8J]YX@IP5<\4.F8QEI\?\1T:B)Q&5;.g-__(T<:<X\77(0\3EX5
51[I&fOP(,(2@9UDDa&Q49&O,dgG,9eX5b.^R]_?d>ZagD9RF+M@eB]Q,c;HG9dL
-];SLZI4X1M9U^M=/+-L2A2A26RE\6R^:,6HHV9^IDZH)^9HSA??V]:FF.d7LcF[
/9aR6#=6(3Q51N63GLG/.Z-1+><B@=Vd_1KDTUU_]-9b0&IDO+D5:I,KdL8[T?@6
L+5_A__Ob<[2L(;;X>[e.&E6^Pc<L?O07=C1Q63aCKV(=&Re&?6.5,[>>+<b7IDa
6,/WF&=Q&.;76L:fG.C&MTD&?N,5A?6;PV,c.1b[ZA8<?b9C]X9>1V[bbM>YDRFB
IUQ3P6DXQYI4GQf4V>SN8OWg^cRY-;Z;?^f&>g2<e^ZMd0&/W5VK)[41>A6H?O6D
].66P<]Qg2Y?(/_:1S<NHF=(8N-8?9Z\&A;KLA3W>PZ/ZA@(SWU]gWD,[[0=Za\(
3ISKC1.d,g>N3OT8T,+e,G-&MAZQ27@;-6)M1,8g#a+PI?SUS2^4>_cZTe^F1,C]
9c0B[_ZRNLM_f+e-JRcD1eJdFY9Zg(8-4T5><FJ)FF=NYd?bX3/4)6Bg:c/C[H(2
)SPY1.0];IY/LA)YgUU=PY94NAA:Vd8NM:):@Z4fReC7LASaQ6ZbOb=Yfb9_\A&O
U_(QMK3YW_>6[8Af3.=Dd2L-&RaaQY1MJb94:G=N(g(/5GR(+5T9-+&G\?BZ\P<2
XZ+7Y=B,)gUFC]6^9&LQ5bW#N\62[B(,VDSZKJEMO+dRE=?D[(K8RBA^77RVQ/Z_
AA6Db8]X2OEJ];J+Z>.HI/eL]GCb1Q(;K4:dFc]#6]QP1&Z4gAM4#+OG0gbBN=(d
=0QgI_A:D-#)@X6W4NCgQ1+28MgFdCT>I)?S3H9VZR7E9X-g/1?(6WZWg<<4#A^-
Y7XSfNcYAUD3<e14)+HgPHMTdW/7>J-d?8=YcN=fL7J;(dfSA)207^,P3N4GPFa5
c#SEa2aM&)7V9YbV1]);JQ)/H26Ff5:N@eCVH\3.SPR><,B8BUe<[?10T&b,VDO:
J0SLU0G#2f4H2DTg;BaE>c;LAV^5d)077VD4__/XVS.);AfNQL=)INO[;Y.E2?[\
Ja_3KCA,+_7EBC:JI=K7A_W;5HL0TJW6W;#96__DN;&A/bS/@Dg=[?MY7IXEC23E
P28WbF\OIHLK/@-3<TY)XLV4G<Ka9E#a5?9+\9.:1=(Y25^5O6SM>JLGRZN;;HL[
NNFE4+2=Y/a^H91/e<b;&c45,QE/Q[M+5^7C6/c7P9RgQ5YgA3YY,_>_7)P+0G0d
O_83T0LL<P+A).aHJ[QWM)8QK(WI?=11a)W+P9RVDU8X<XPJSYE;dVbB.W@fA;=D
LDTJ&Q^Ge)O=:C?HHCK:dgbF<RU5L#/c[(:]f\g^b\&,FR;gb>EF70POIc4+aFPH
DV&)\JQYIEa>1P>Q;4OPC2:D^#J8^+KdU6XGN:UL@_CJ6MG)XU_QR]J7(FVM7L##
a6=PURd@_^]Idd3E#:KI@?S/+b.?,T<c23BYM[bE+c012.gML/C=,W^?JME#gKdR
b2ML-(UA:(AV)<+F]PEJ7ZTY/(dQ17CREI>KfEVd76gOJIB^TQHHfO38g?.F^?59
W(Q(IUJ99VC]/cb/a6.AP(gZJL>9dc9XDY)GWKQOHL[7eG]7=G84DB+&B:B?f:PL
I.dVZM^G0=&@?FbgF/E[[CeeA=W,(c9N4:@PKS=0P;CY2V\M01+&ZG>@P>CY2d&+
>\PXa=BbeV8PZ8a34g&9-\eAOGTV6O38eX1BS@2(0\?6]C]^bTEa2\)ILW70S9f<
b>GfV/P.,SZGM/^cG6Y&CU]Ua]Xc4\2)WD9/4JV>+CE8W>,M&dU[#BM,ZAd8/D35
A]PcH26O=d4Ce-40Rc#eE,^Y5&(JNG/RV?>d6bXgfV59O5L\8<6f/SL^)M(/X\4\
LB]LQ1GS,SR#1.,&;R(N41f^Sg9L13A&E:fB6?\FQ<GfU+-@QK).T(7KH6BTd[A\
@g;WAHd=\/#6;7&7N_3KX0eeB]HU2DJM9\[97BV#SFE;c_IXS@1?Qc91A(SM+BCQ
e:\J2JUI.YZ6USVHg7<PYSd4(gRGHGb8eF#C82b-BNT0/+LZ.B/bS/EAMUCK)AQC
Q<a+F^fM^NNbZa.:2<g?#+f0eg<[E+O/bcM&YL6=LVO&7X,1(eD;:F5b9HD7<\NW
;fZDQ^O)M>DgW04C[dXDJca?R8Sg+SBUOD^b_?G7&,8,QJ/:Q\bND[K:#^,LF6J_
2g0Z3PQdg-[8BaFg,PT3B@gV-[64cdV<(&=Qe^-.@288GN[:TS?0;3HWJ]J6YC<<
V.)7aa)V6JT;gTG^P:VW(W&QL(eJVIC:7Bc6&8Y9Ff;<VM#F#:ZgdSc6ETb<&/dY
0[.BU?(U+]SLFOH)7c7X1CDQO?PCWc4LCN2UPH/Z_;Gd#_.F+)IaRC8L.<;^a=e2
FG2:P(OCJLcdMTbg&(c=2Q7YAVVAEVQ;IH2XUQg\>,eJc)I/>1b(KO9MaJ^-b>C,
NJN0#U2JW#/X?I2#I6HQF#I432JM?O3(6F-MVY(66TCeYId_F813DO(2@JYD>KP[
d0^_T]?C5JV/I()6\)AgFR)OL/@cW^1d_RV^9bS7LB5H^V]cA+<?P@;6C<S3Ff[6
eVIeG3CeBE579;5RL[[N3,Hc0=G#W.IIPYRY1Y4BWXfP[D_PZU#BK7H-<-I4f[)J
>#P5aM;D<R_-Ga?2b3GD,3>=P-]L:7AVPeec^4QUS9FZ[&d2BNWI+8YAY(A-QC_A
S:)bPO2\7VZ2]FRBO?(;>UUdAQWM@T1+)[#g??XEIO7G&&:6?0L/K5WX?ce+gPJC
g4/ff>POc6UYPUfH[f-D=.gV]M/GaaH>dcG#E4SL#QN^<\+2I5,.B[=8MV2gWYRd
I.[]d6g,;.O2&cAOcIQ9??J(b.B&ER;=69O1T]7(IeH.+K?::dgY#\RICS;G5)\&
1@UE]UDMY(b3G;g.;I.N)FIHcZ?ZQf+,L1G/b8AT_5)\/X.;]0PBE\IXAVOW)ZBG
.CFX:8\:gf5deB_>+aNEL:3N@K#TG).#4^?KD_80.M5?/^KQ+9>^)S2cUfJ,/-;9
Ab;Y?#@Y[PgFD:=D#&&?DWdc6R<>>@KM^)2W:gf61?U#b7d^^fGUYO;?1aY)7/\C
^7H;a^,45f6(KD\.QRSZFfPZ?4@c7ZVD1P_+0-&]SIA9;QS=2KFWO_1Fa;D_(&a4
gK.]T4[<G_#R1dQS/QK^BcEHUOI(PbT/?d7>,6:U=]@T]@b.Dg6NJO#L-)Y)XG2S
e-9/(bE,?.6L9HW@33E>8QcN#8=ZMP#S:&d#a7,5gcIcRBOYQCMB2#>f.PLM&R(\
fa.URf6(Y[:#9f>P)c129L1[OF2,3B6KMgNGbGc#KDP;@K<.AW>OB?WR1\38(eBb
?1[7LS^<TfGMA&YOMF#d0XCDc\@9GY@&BP_Y#X6Q7CQ582/RLPG]^G+W)=[I&PMW
R+Q=1)8-c03CVEbPaZ9TB^b8/K:F.R04(AIMD9P8d#;(dK8RC_7[NOGP3g,b@EFU
:8[;fgE9)bSVFdDH0XYg9RNWUQUHOZ#N+\,g53TPS^U4e0SZNLRG(-7M&9BL4&Id
1T<T^CD96Z1:9H;g&5gJKK+O[RdcXF3?(_@[EX?RD4J.=(AC(eU3aQ:G4]\NMQRg
?F/J7W09gg+,QV0N7&Y6)FM=V6M0X;VNaS/SIgN,Y4G[^B/(;J8(X20OYHF1b?YM
Y19AG9TfKK_ZFL,&#5,#60a9_C&#K^dQ::8PF=bB50=\f^G0f<0CBKc4RMZEcT-e
I<ETBZC3H:?aFgXKT>2eMBMG^NJ91A9(CP/Q>BS26#Z)N&HMZKO:)=);e,+(@9R#
?3JCW/C08.5U4F+(1,:4_I#>-C@Kf1##H^g>?26bOVG6I?MGQ7OO&1<I2:e-EM+N
<cee8Xd1?gP(C-XLCBbM;E;EgVDLEfN)9,KE>1/P(LEDLS(HaI<5)S[.5PS;7bdJ
)/(,<F[4-6R\Q#XSJ_WeB7,=]LS?K-A0=242N_XEdPYU=Y._6[R3TdG4/H_ICc&;
^9YEX?_18N9G+W(M,+E3U82caC7ZX<SLPCSU,K?f2+/&H1OBUB:ce\f:L9I7Sf>&
PCc@d=aA^2b;?Me#90X<U=\-7@-JP.63DdeQM3^:aQe0X0MU4<b\92<0E=M&I;-Z
92f_HLNO?O\P@cG)GEK&K316NAUL>U(KcX;EPY^>Ga?97K88g2NE,]T[6GP2077&
18EN=e8?_Jc]A6)I:&6^(WDQM(;[4/Q0>-d<fDW6J_\6(c073UWGZ;TUIF<H^V/8
fEK2FB(Ted1LGf_eJU5F>Y59)ca5-PB,5X?=[Y/J1bTWF-X#SW+9>(NDLe2)7[\[
ELfbb&L2ISXWAT)K)a2.BGLMU.3:&)4M#FV/\KGPIK\0c3H>BN2TRL\+KMODC8FY
78C5#JeRYX>WX>1N.UK9]U^gX/Tg;(Y)EAS/b_If(Q)VE\U-e0^TQ?Xa#8:d>((f
_fVY):K4Xb9#9;(8a,9cK\T\@\EIW9:,6V(&_d4;:INc7QV+)0e<DaXdQg.;;@.G
.HAd/Y.VA4bC9VTNHOIG&BOY]6]bN2aP(2:+,/e13D<:P[G0AVaMgYFRD3K/_LQe
<#E4U<:K2dOdR9^R-IY86_1:c_IZFXTKPV8D3,W9UUPa5P8A6g3EZ/J9H;47[)7G
H@Vd;<.QC8Z?[-<J&<)IbbF,[+[FMbVPgfVZ@[b\GD:\^M<F=&Og@D.eRb8AAVg_
MJWDU/#^D9aV\KO]&UQCdAK-6Z7fU/=XdLI<P^URU>LS=UT=5b4^a<,S\KYW+-Ef
)VNg060e,.(Xgd^T8SV1D4X==_R2H5+E,.:Y11#G1^8>;>4<+QZ6/U68dGUWV]GL
TK/;2/&eC&Ra(=/QGL6+8;##GAGebUBeV)Dd&>7bM(>B0+G)c9?GJO-?Of@/\V?d
<=(&CZ/Y-U^a4C]De-(=7CRaUK\abeD-Xa/=?>.R&Ic4Q7114@;cQ^9f3QM@^bS8
LXd@BEO6NI=bcGgA:dX>N7?b=?b+VG)fEaYCM^.QOdUJ2+.M#&3NZT9>G,Re9#fJ
=N,^+)Y_YRX[M2)>L@WER>Zgg:)HIB2Y=>/RO1F<a7\=]JR/f6K+)@g?cc9S+L5-
2e_EBedPT(E+62DP<U7NRN,.;@)LKE2S@@F6?>D_N&gcVc7R3T_P;V#+aK9AVA6@
(,d;V_bEP^7=E3U1^a[^:,>)^2W44#7cb7#3:bfg@acf1:WMeJ/M8d;HR72Fc/5S
TLL)eT?9W+H=@]8bU[2BfZ^B4WfJ5V;#,/B^))R:..^F^8S7V^S07d&8#F19bVJ1
<(S]#RLY:9<MZeb<g?Y=@IfSgFA(?dXfe;a9O37(G+HDUEJ/I9G1[aE-HP-[bJ2I
SDN,9/f5?ZDTA]2OX/L?C_AE9:JVJ(g?+#YGF4D[JDH8IHd>Y253fV:OBNdfCaW1
&<QU,eaMYM>(]R4\&W)G:=G7/:D^_Wd]cUO2XQ:XS:U>&3M2&e0L,^R7;S?EeU/>
+\@LSVVAL4N,4IGc^cHXB:FZ(cZ0@6QT411e.deA\-PeB(d(fLC1d+D\S+@=8H=&
T&C(QbM6Aa^6QL(Z4+3U;8AF17)B)E]\K3X/)(4H.BM1c4MI1\]O;]5:>-OD4Od.
-\UKSW.TBIM;,ACfGT\[\0YfWa.@(@CXPMf0BPF),WLP5;WZU^dSfC,,aC4f3WWA
9gDPT007&V+WF.Og]AaAH@]WgF[2[>4]ebXU72IWEMTJ]4aDU;ADbTNe=b^b2?6>
C[TS+R2e@^#R#9)5E_HQ\2.HR43]RA9Y@>2UD;]5HNfMK2f9-:YLQ+8NL41F-O&5
2@@,/@FAXL6X,D0.SfZ76M=]8.R\)6gO<NM//RG&)7=@W@;A=EO]@b83.[\/.ab<
BQJ?^CI80N+JZ1HEZVf#[JF?Hf:G0Ke[&2&-gS0O9)gL>)(K6G?=XPaGQWEbNB-0
9cI<L.2>g6JP@.^4-2O>R9\e:-.)3CeL3=TBXPc,CcLUJESc8g;@Tg+ZXE(<72OP
QeTB&-/<)\;AHB(C(d:+0KOK/,@16ND#F0NYJF=YM6?^P,_a;deJA:KXO+1MNXJa
J;#Z5)4I4N_#P-85L>gPbf6I.f[YZ#\W:2H+87II/.<XNcFKP=b8&3<[Y.FPg?B:
S_=N8]+g18F[QJWBfJP(:PLWTDbY2VFdV/L[PS&N7,O#NI+Y\]\KW3e&)W&@aB@B
H/W<dF3-GO0PZd\ORXG;aC-D8=3016-&M7=Oa&F/7-YJ=GW,C__19K12.eOa=c:0
S<WRE/M?XYMR6,WPb\P?fLOC3NRS-#U(^+c6^VLULAgTX:-Z35^MV3F?CME,P^bA
Ob4D#.cg0b6FLX[HB9I:[ILY+d0b[<\Z</3HHKTgT2U/@[H;^Y2D.SUP[NC^33IO
KXLg8TfeZ&0WG61B=d/MR4XfcaH>;3:TMM4NeD0POa@9(dUCGNcP>[@geLd]e)5B
4[HcfNU>MW)Y91=^UdV+)D]G]^S,&FX/:4&&//_@)]geaJOBS4<K2:,I?^<?a]0J
>+(?=T]gf</0_=IH8a3_4I?D/Z8;6C_&eDIK9/6IH?A+aI9Wf)dU(IV;1XXN<H;#
26<60gMBBUdPC&ggK.G)IA-M9R[=,9:MPBcWHV7^92O@HS3-+[?O/(SY]0DRQ(H?
>2cA:F2(CEW/]-6P:V#+/,#V[?=GJ4G-3&f2[g:(5E.J&8@FU>dX83FaX91IHX_0
_Sba4H5P5P-YfG)O-ITYD:R,8ZNSK[9UME62)PESfg3,-P.(.M?U(a]CX[S;/^\E
^X]C\b(TU;BEV\QEXZ>(,+CgZXLNY)g4MM(]0aP\APfcPHbG87\SD5;,:&7APOXJ
Ed8/cHEZ];,<O\:,[g^\VS/]MfHfgL,7.&Cc&@(]J]5ebA1E1S_I.(A/S=9X)2.\
YWX.g,db?85PZDTSMeeX<@IJ.V7#R@L21Gg21^&A]7g]B=<:S(.ab_eD/K@.3TPV
bUD>0V<[8UU,HMS6FX(1I06?b]PWIf9XU]LeD21-cP59MId3B&/7bS5Z]2UW<aNB
Jd0K<9(;P5ZH;GL)MJ1g.beRX+.0S]F6GN3]BdRH,@bN8]fM+^I9)6:f-@Q[PU1+
,=TY2f^>[CeOKQeAYg<fR8<N:TCPbS,027#7E@+UY:;M)c@/KI;)[QEXN\DML-RS
\IcA45X#<]e4+SR5>&KEQ,P0dE6A0I>SW30HWY9WYCP,(c8ZMFY<,deG-],&KIf(
GfGegcE/]JEF_+O9)WRQXOVQP(F4@3HQIHQ:VN0fIX\PVY<AL(#;I2\J7-[38?J;
gIb&:R]B6AeB>YP,02K_U9XSXD[c9ZbeL_NW)JZ#8HKab<(ZN]]aaJR5@>DGM,:#
0fD+>[>RN>#EB7K?JE(/:&6afBJ3/AI49b##6J4@V)]aBAAM][9]g@>f_A^K;#36
B&QLQ)X?H;N/3@@0dZU1[8f1ED4#Cc=82BF\&N\D7;0\Z@@]8EY8[-=I?EYMbQE4
.5dMZ:/YQ^F#1Y\5HS7@>2Wb_=XfGZCQF@LXX,YA2_9D^=Q45D,WFQ@_YLQ[L,Cf
G-(3K\e/C)RX&5:Q.K+HG4d#DfQc\4K-0OGe<6JY6QgS4XdM]>T0/VWT;G6d@?)>
ENN3L+]U]4&Q(TaJOM]0=+\WCb_OKY7#Pf<O(IHWM8B,HN-dZMPZEQJIc=<-XQT(
;;4H8BOAXccDZcEEV:P().W/@2eTXP;&d>R80NMDUf#ec.a^&VL7C-Q,aYT52&,S
YKGDJN(I=4O--H3+O=8^QT9]8MD,ZO^9J^bNCcT\6Q/AE,5/)],4\L@-A9&^aS^<
&^=6.:D/7a4[V5Ag53[f7G@UVVEKdGX.-0)B:5F7f^FU3<0:/36)3<cVfH<7S\;M
KRKcD3GEV]&L3g#&+\JFTE3DD.2>gb\S#\OXeE?0Y6[=X4NXG:S[+LgE]e9SE.M0
8N9PW(CMP#X+UeSE@8=eQP&>9P=G@g:]1G^]7\,Q]\PX+3.^[EL4W()9_W4Ka.WF
A6GZCb1=1e6+;H];Z=2+BfFTQVA<.R9,)Y(^SAK>J)3M:ff#VOL>gUW)WG.#->e+
/:AZEK^@0B;A8&Y:-2Eg@]AIP_;AWURC4C4PD,#7;T=G:DKOKafEJ@+XM]DB7Reg
dd+_TX^,0U(ZN?K75,G1-e9O=bW#P-P8(a)J.&N4_G2:6Y30#HJ^4Ld=fd1&6?EJ
Pd(-<\X\(/:HM,]@SNW6EgG=^5]c5WF)dPd^1-MH8dWQKT1K7e[C:9S:&-J66a&a
N/6R=-8_&Cb=4,WAD:&9QIG:M<\\TaDHX4FNU(Xd8MFSfadZMV7cI_<?fZaDAJ]\
)Y[8fAgD2aC#;f(855<_ID\W=I/=b9K8MIX7L\07ECG2@[.-PB=27^E\_XBWAeP,
1NN9RGD^FPEV5E[<Ma8G<]J96+_H094Fa&J4AE@DJJVbcUFL#L\fgcP7\I<.=5cF
D?@P1JLCU&1dY-;J:eT+c\\AHd:3_,.bT#5Z>M&MX(CCJ^56BZMWb^,?#\dD^[RH
O/609#dA?#F];#OTcIIIF&T]M2TcIZPR=P<89)+GM#DM-VIJ2B[fdbGY@@QQ,7./
?8THR^>\g?WbVMCg0d4KP)aOFQNab?9;3T\5W/;R2K]WDA,CU,:7+e2=,,IMFF0M
7=\IgS.TY;EQH.bE]XGO>D@&b5TZ8C-_Sd=M1&,QG;;9(#dSdbAIFJ\?8]I<C=A[
USaY&D5U1dXN[@Y2IX3[&F6_cG</)DPN\JFV[L\HaD@Y3FC;1ZQAX[7L6TKe6&_f
3>=P4cE-+8;TZ]G6L33=f4]IfUE>R>^-1AL<A9(-RMXNUJ\Yf[O]]GDJAa&PV208
bNR;3b]L6N5X<H[LTQeW5:@BdNeUK\6VXZ>Nd4=7.AF#_)f4f6MK:@=6QCR?D]8C
YUGJ#@Gb[5KG,bJMg\9;F/1_be]<JVICX8cT-;=LL2_a5AO<;GbT0[ZW^HLAL)aJ
53@OJV6N523aBT;/JTD=\U8ZK06?JZcA66K@)K&,CMJ&?<da\26N?F6N6=GF-f==
@3D?LN@KJbA8UVg4EBJZfUI.S9Eb/SFHP(DOBSV9161T#fQ&KcFX,3_BeYeTgUWK
7J\aHA\./,-A\<-&T6@9AD5L=c#E-de/4BM39Y@+-DNe1B7?S)1HN5Q])-Z:LJQ.
B-V#HI@5)+D;LWg.Q#V\G2.)&BPZGGEb,g27eW/D,@bZ4cV)4#dB81Q8>ec4.GG8
D=c^X<dDfD,AK(>4+Z#VAa9Q@-UbJ#<)Xb]HXgO1N9Z6#SIaCLO7+\gZ7-/7DbgT
F5A7#?0EV>e;QM_Cg_U+A,R.-8f<J7SWPWK>IE3E&3>T4IK#-JG)Vc#E-?Bb1S?O
:c&USRfNRLH?9U_/=44G(,4P?NKD&5^g(#GGL.\bPRYEZWFE.CaH+P<>I#a?c;]G
WJW:-1-6(RGEA(C:1[.JH&C/7]EV=g892;/d/YN_^P+C:_6_Z]?=T43W0AULG+1S
N6UCVg.]JC[LfD)K^PY6&X]PfXc@CAZbgJA,4?c/;d[EV\JPDb@04?ZV;-]aK0(R
QF)7e_GSE\@[JC3;0CFKcdTTG&:UfN&18Q2?e,7LK72BcWN=(&IHKE\QO+E27\C;
E[2^KAU(f9-@HLf@/7T3&^=cB<CWK]F#a:ea2N,PBcMRE1&U\@59a_R;KO;bS]bE
e8RXY^7<^XQJHEEJ55E1FXKV:4d3^,^b(6MDb=(<A<L?C,HDZXg=/e]fRR)YJFE.
BN>@Nf\J.9d^/R\><.Q_=?IF./X:P^B5cgWca@(^cY4aAgT==Pd7F[+I8ff_MEaT
R)5/cIT+gJHc3-]a-W9adSePZS@BSfceab7=MG0_S2GK4O>XQB9P<XM&M;VF_0^+
4gE,_[cTQNK^>3R2?^:9)B\R.0#X;KV8OQ;4>G>A^QDM&H@bH&J78_5UKLM_\L[G
aJ0S5(Z?ET2f#1(?_)2acJ^4;\B3f1Z)<Xg.N#H_:&+a5<TLE\&f=[^Q50AR=:A+
N[BL8XG[TegM\B10eGPZ69)@7NM&ECM_M)U+[VK6CH:f&T/=/4CVQ,96WV\:W@#3
]gXB&,bW0B]@>YODP8ROS75UPW#7ZHTAS1T[]F):=TedF;_HOe?.Ce(R#2+ZRb^W
;?6UL8LI@^JH\ZESg9fG:@[(V40]^:MSSZ7[^7O4V]L^@@_QI\#K(]7-0^QA:4Y8
9:8cA;HDWcP5VB5c)dAF-H&E[SSR?;:V7QFg9O<]egKP67#\VMRI_Za7_gAQ+gX^
VD#UCBT>]C1&-=K_AOUK02bK2Q26gO0NJWN\EZGFF=dXF76LCG--V4O1(18:,M-P
>B6Nd;?;f1HDV]TEYVG+IAYd0R]\c?GQ#.T65;ZP98VcN)K2T8QG1fLb6ESd8\6.
T&=U9-E&D9F?(AVdaN[-b9aZ.6(FC)IIQYR]g+XD@B-#G63/LOG?ZT,/9N8(F(BG
_E:M+Fd5/HG1QT;\5>MOLYF6d]VTLfbO<-aS(]TIb.ce3E][:L+WX4]STP9Y;Q1.
A-8a+.5L&7:gRD8@9,O#,>=Tgf=\MLNbC?-M7L=ES:?K2SW?O[a^V0[\]YHdZdX5
eOb,K??ae7;1=Z91I@[1,?GGIe?)=c1a2(GQ?O_Z.(;f,g,=>;->W0HF^\S[FZ=@
I)XfXB@SRgBN<>J:)?I,M#B56:Ee_<9&2?(\03/AP^]2KdS>4QbMEIX,PY;M;E^g
01Nc4<Z@N]5cIJG)KCNP(W[7=;F>UB?1VREe7gNRF[dU;-HA3T8M#D\\O;W>bc?>
>+.e_USG@7R/@4+,O##,(+^Ya6g&Fd+FDYf0dGd1NBKTZf@31I7ND/_fbTE:T(&-
/,B>ATSEM,=R.X7b=\[]5-DT.T16cZLM19+^LPEF+R+:(0L]?A<8WTY91Od)JaZ9
WW8V@0R&DI#PBc8)Zca7_^]>/-QNO^#:8Ac)7ANH35R8XYDTO,XKF:O0UXKT3DPZ
9?G>Ma9FT#K6+_^O7.gd0SG94JV0D.gbBW:K;9JVN3]9<#I[/aTFaLYX2ACe[1^V
1fS7OI.^ISC+T[[<MX:8[<O()1^F3,K^DMH^X&30P]\]5;N1VS9+d-<SV8>AbgNJ
\&,=YFL<J<F4)\#WfEKTA/bg<gL9<=+KPd#@B6MLIU[MZN\6P?LMc2M]:?((3_?f
f//.5.aN1FC8;ZL=bOgJFSIP59SPDSQBFGUFe_NA\fFM\[FKa,+@0BR8H@L]E;6c
6TIB#.b99O#<U[eg]0.5P^f(;I7G>R\+?K2;P5I_C65=bbW)4,cTX2_10+1db86a
e_VS9d7R\&_B0b8R92BRU.-;RD3W/J->gT\[MY^;dE\-/M8a.^<]+J_T-W\[MCe/
7X)cWVGM^)WWF9\f@RZ/TTE8XbRe6V?8@-QLFX1[&2Eb07.DHD)B&WN2>eQAbSG]
0_fA[WI\M/>\)..KMTH,A6LJU81#bA?&SJ1.OQ)VgV.R)01S8/Yg=c+)X2[6KD8Z
0DP^;&J>+QB1(g384/U??OX#:X]adcX[G1N04]OX,<d#aDY)8@CA?MZW5]DH10=;
>IQ??Zd)+J1)f>GZ6/&A<BZVg17YV_&+]SdW):61d#3ISe&3F>_c:FVCA)X047A[
A\gO]F)E;_,R,PQ<@2)B,HO)A/3,\5L>(L@@3V)AHg5\9EUYY_7Sd_>WgL3_V3NT
KCFW6OOf_,edaWHJ\K727Tf.+<4WZVaOU:fd/]VO-UG/DL2H-TNJ&Jf>28<(WQ7c
NY^F&Q+&gSLZ(CROL/R5fW-0G=0gC4e^gb?1c;>W&HZ#4/M(JEZ99)a1@7F<B]&M
<[1U^=).B>\YYOd&G/O4@4a==XJ]5JIJ/a+K2VN\gJG#?,+MSZ7bb>)NH9&Y4-O[
a3=G0g+KLF1]0G2;:Qb]H;CT4@4@JdE-FY6W&^g9f](<aHfZ04U[3H7JF@J)7-O1
T0S,dCbWDMAKSE;P5H?]9M/4]R2BTeBcJNS)(Y)5fJ<>1R.)b1QYU@77&NZ57:SF
^K/(Q1:M+(9JF?+=-8a;S>CUfTB]29dX(S7W2&H:,LSR174R_cM;>Rg=EPObX2@A
[&BW4&7-0M#3:b02UK3ef>V[K=Y;5[F/XZF/:40cdcI#Sc\_S7MNb4R6+SDV]:9N
R2HdTE]UYcPR:_ZU1F5:I^#,H7GYgEF:/e:E^J),/#<I0N1J?ea\FLcXB<C@5G+N
-0Y>NX[+./5<CT-LbL0=8+&-Ff1?F14egd9+&5d;>_;BY22<fPe=?]5PF>?S&3ee
@+PQ/E3?W]41fgC&gG5cVG]:S)Y>#IT8TRQ\bMg7>V/J;b]F9ZJ1RM=&D7eeF,Jc
.2LA\^d@8:(SbS^4_KfJV95?TSIGc38Gc/0)+[RR,<M&JHId>+aUM(6>?>?10d.>
@L?_L2I_dVW5Gc;S3ZaHe__d41?:+Z<D8&NZF(2ZYdHM.\G0(S_c]\;8^G^8QAOf
baYe6e88dT1UAWNRf+2Z.T+;Rg__3+GPGW2b/N>egV://7T9^I=NcfIeO6(2@dNP
2N&YQEW)]KO/N@@^ZgZdWUTI>)YdBI@MIP4>^N83&4I5HW5.=LL[[_gS?Q>;E9U;
X\3WK0?++ET5A3_&ET+79/]5@O@6;d4RI1B#.e+>YJ-([KX.;HeQVZE/EbCb3)\Z
6_,K:ATXL]N^ZO]TK.98;,5B^@RbIVH@E>)C6Y=Y7a(\@.c>3ERbUUU.]E,@DYA_
/a?\DT(C&_eC&U;;fF6Hf6-bPUd8cND7(E<UI\H++(gOB,Y8aY6K/DX+>+C++\,b
#A<2RMb_,H#VT1V#PAf0^a9G=^=T6AF__NBFI;a+::fC287/E0VWVL+CF#3YN@6D
[U9K(WFMOPB0[=MK4A7J2:Ed#0SDF#Q<[baeK:R\d3ODM+_(@;^-F/3#9-Z79DIT
1E:Bb>4]8<R,BPRcE?Ra=#\+5EI#aO^Hd,cI(5Vf:K/([:BVQ)4Gfg\2bV/4.MD+
9.eTafP)VH5=B/a6Y+9LeG4DE6Dg<2;(]ca].?RbJP,(B8A7B3,&#O8/#^]I9,OG
UG^cU8dIa[+UA4d._/GXHfe,eU37c6K=SY5BQ?+@@cYOCJ(>>?H(a/Aa7]VM<UPd
ZR(g.d&/?F,R8Z[)QgUG4g98Gd>25D7H(cAQAcW^O<\S<f-,YW5K[9R@cAc#/Dg#
BPO1/E/g9N7?:1L95YaC9>HL>Q8Y>91&_N/6VTR6^-,42@Y=/J/(dD9@8ZAVE,CP
dWU\]J7S^cW-9R-YFU;^<#A1J1ZLfT+1G([X;U-bQYcA(:#e(79]RJ+@EE_OZC23
J7KW9MG?S1^deE2ZL[/&([TYX8DT2QF]T5Q^DUV\YB6=0IG+.-@\J2^;H<)g.],;
QdgX[+AS@eGC(6BNgK9cX1DO[?_KYW0;38:L8[NS(4Q7J=ed#&#JN:@6aL;9>C8V
.S-#0IgB:;>_3aMB0)O@63f5,CQ<UV;BVFF07/WZRIVC<=J4g^4bM:L^(^b75>B7
JSU^4LG:f/J9>2CB_fRb3/UQG^gQf0E.G>7+@T11.4U&>DfL_=O,80>0:,&,NgOV
KGe-FbZcB0_/f#)0(X9Vc[X-R-N<AE9FcA@\,44QRg0?_XWeL[8:SN_19X/7&W/4
4;A;2])OM-[8X/J;VAMf3=B[b<M_2#Y_KYc^Q(VV]FN<M=:]gfc729NU)+bD<V<M
6,G<2(#:aF+=NXEG0)?M.SMbMCI1&;B:a;2,]a=QDET.P&M.M9Z/aWVQ)ZL1/F49
2U8<GV(Gg=C4DN\8ePQY(7)RI<b0\[Z&Yc:gBZJVC[=BZDKLME8JOO7f7UJ@]_]A
7+-R@1>HLgY>]KRZU0,L./_2;IdA-J;#fSP:;E,@33cO886XLg02]XW@SK9OaI?a
\Qf;?K7UX;(/IPMLMRPR#I)HeD:\WK(DGF1<PYO902OT2R3.G<A_#7[9,gbUNcH7
@@UM=c<gY&Q5D5eTPIU],2-baadJ](AYL7:1:YCa/W5]?(?#T+cALK]2U-3E-YDY
LY43AK<#S]:@LC@70d_B((?EEg\U&,U0MgO/S=8GS;;?F#fX=(&#G-:OPf]e,WZ3
)V3>Yfa)^QQfg,g@&[8W&N8=0dGG)+:/A#a5IX9Q-gB1,a>gR>,+JB.JQ#9Y2KXG
96&\K,F^RNVB>RHdV#fBY:6F,/R1Q:g59R6&48-10)HZT>7N?[?a]U#M^9SOW4Tc
J-HJ?>N^,I(C_#ReXRIPM<AU3Y5#AWF.=]_E46GF2<f@IY7QTf+c276]@:O/WKe/
\66eaL7\];X33K:9FOSO2UI-J4PB2L\.aE94:Z1Y\_F,2:NK(>cY&-XE,&NI4UaP
UgQb=/Dcc_D.PG&8#2OZLWKQfU@KP_LGX4(+I^+0_XU(dGI>eNDcN//VWIbeH#37
<@TS=5LGMD>?D.=[6.JBL_QS8JE7P)Nc3>M[Kd5D@>[7OXR6[9I:TV>fSNDfLZ3O
RG;GfREMM#Tb@JfCMJLbRCdA-ETc;A/F;(eFMVZFV&)?0&]c:2bU,CMP&P01_?\I
A7JWIIN1Oc<1M\;JEO6g5c8LQR\:VYYI13=<S=2LBQKA.]MG:T9.&WWIB\>GYQ6S
UU+1(&fN]^+R.6[,,I)17G>e/8)bYeJ[::bBcS3R-Y6O)5-:M8c9,UB+2(GOJa4R
EC@>)X^&?S>11IBacJ:KY3M,K?P^4D>>\9:,B6#3aK0fL^P98J:?CU@XJ=VL#a[D
?5XZ,M.d()M0H71;0B#H&E.WR+SYa,;^QaOLNLJX8AR_ED@&ER^4=MZPId4H)EQK
,,\=/H#0aETXB,CU736WODCW:9Z-RY[[H]Y=A_WW?&#X2(:KO=,eIN3MF[XM^M-?
9O+aZ7K=4Y)5E\55_<I9#G.)&bd;J_WUAX0c_&d[_<\:HS3V@/EeVLLF=K&^RYAX
#ZcO;50(X48]2L4<bTZY(d/8.5E77ABXeBBEXQVcCY/B]0C>Q+/N?;YNFJ04dL0X
_RB/4a9#C[?E@a44Wfb^5J8ZOEKgCEPT@JO&_.?aW0(MD-fA7#7O.:C:EF\<9>>A
EL0B@;?0CFY9JXIN20A0W\K5W=)(-5SZ6T3AW+^[>71KJQM&=deRH]-^=1]+B5ea
\KSLJeLbJO,X;BK&gc^N^2.0G9eDZ[L/;JI/7e_&#I@0-E7,7bUa<#g._GZ96.[1
KCe(XP0dOMJ?YJFgF&0OJOD/aO:VWXf4PIN)(>3_-bc/^gX5W>M(.T0YQ9-6f4PX
QSJ8HT>FW:=\ATfeQ5L@f)S4&>],Q=B,d9YN5OgcQOHL9:]c^I:\<D#^?JJ-E(JJ
.+G/EDFPE\LN3AWYOdWHb<\=46CdC6M8,B.O@F4N4&6b6(KFPIO.+#T,2PR>.8g4
6OfY2.8:<SIN>\CUTZTS0)V(.[=.IUW@GX@=B3KJL1Nd(&QI3:886&T(Z\T=K@Ka
EG__5+FWIU^@UYd)U4+Ka&-]G@?Y43I&?K)&S)I_g\2;<Jd=V+a1[HTT>85WNbEV
CgUg,T@BD5Xe-EJG)RNJMIX@[5[PMX+ZGIe6gW]+YX&;P)AP)&DeS;8CE+(#I[4(
U4F>MK?VEAD1TMd@K#eCT@[+#5?cOYAPV3N]Vf;QM?:7KHEIbE+(4+3^C]<70R+-
<Y1[Y+3C[NN=f5XaR.g]gR>XR_f/fL/UZGg[.E8XDO#;MQdFH:5.b<g1PTQ+>-c2
gD;\eRLA0[C8Y=6<)J[QQ)XGSS5^J#T,&U(QgE5&(.YOY<;[Rf_1RSc4)ecLFa(A
_g7,=;9:HF5WP&W?;Pc]6\X0(<YTF)8Y2Q7FY\9N(I/aYGfWAGfZYC3:)bV51Q:-
J_@C5.;_.:1:Y=PLG2U-;Nd,[Hb(e]gOeH4d3&72;_LXdY9RL?C0I8^#O6VTZ-+R
RN(Wg05I=\3_Rd837_LC@=O#9Yb=IRaJ..9a)=b+,dcS)8>+MFdT79/C^U[8X3D?
\0,R9KOZ@=7XI,J7^AfDVLZCN/CX@MR>SP5L/_@,8&0WD;P-X-Wb#GVbG+W]KI97
G]PbL@?0a6EZ#GLGF,e,/52:@KXd-1]KZ4ES7,THaed1KA7#8^DNO]=eB8847IN+
5#HS72.^=-ZV[[)#EcGZQN2\OWA_bDCa\fKV-V&e5^GDK?16AVFQX4ZRJ,fbL+KG
c1;NV_]SN=[O44]VA0VT)\NTK9+Y1OCc,Xec<ZV,H;JY]]f/L5g7N\0O:>6337ZB
LT@UXBHYSKeH<:,&b.\<gT5W3K&G?P/eMTCc&ULEVN@gEb0Yc:RFT/<&2W++O#fK
@^1G/<G_C)C.WCUPf3.T)P+T(bN[^8_4W_AYW>GB?KC:dH<,,ZG/E(DM?;ZL0[^&
F?/CQ>=E_:2-@dDRc2T+JdBO5SDK_JbBBSU9HNc40@gBO@2GXPC7g)MQ\EIU^U@4
VOIQQ?N]^H\A<BL/@fS,[?^cNb2;XR-G:@NAbG[J&fH44UV:J,TV8dZAe3Jf+NfK
G)RSRZ)(G=eJ+R;,Xa7=]LKVd+W.4FEK87GR0Y,6CE;3-8:;-Q#E5Y#c+;IR2eQS
K]N>d_Hd2?,+;<XI-R#O0IgO#AIDe;YVA@bQeX:CU=70T_[F;45fIfN(b[dOb614
.79>,A;)Lc5K6ga=_dT\EIVDVc_+)0C._CJKbX<C<6CL<R=^9RDf9SI6@cc+JA-2
)2^5&:M=L[?Y[AR](1>AaRZ03;J/P^LJH&O,YQ0:;B[.G(:6SHQQg?.bU(aK0X6Y
LX;a@d^HI_^;+JW]b)D81&H<Yba86S\5a#^S8&+OR;6.@d_4[f:c4,b0<U#Ec1I?
fIT2O.9@[V2]Z;f=EJ4a3^B=G<d<;#f^G7NCC]N9B#^M40:GS:V28#>;Ia@eJNWN
EH(U_I8;BTCOed28JAE_F:@2&1c6e5aL<_#UfaZ54S>U[]bAHO\F;7N;2(5SQcZJ
(>=H]E+ReP3#H@GeC\1G9=D->;REU0E5D;V8U<)4D/[[,V=eU2)fRN?fX=+(\8P2
C:1O=C1+QDGEMUHWJLZ7?+\RbR>9f0GGJ.+Pf/c5a/#\UfE4]:3>N16J\>QX7[8.
4GAV&E7/W2/4IOLNgYbO8CS)65=87f]XO&,_99NOJNRAd2g])<[1_(X6O[.Z3bDd
A>C6HVWc>KRZ8H8X#:ITRT>1@W:2>Y\DMZ]VVb3KA#d2dEH#Aad=AC[Z40JF8GEg
N7WLg-DA?O\Z2f9ZNIEU9_F4_;;2#Igf595DPD^2dB7;FVPD0S+0/L0/VK\^KOb?
dc58a-REN#.N85#-DZ>8W\&:71J4]NReK\#A,-gRN\\Og)LU>>K_TN?))ERX.bJ1
]19>VdWN9@[D)8A[G[ZX#^/T#W>L0]:52WD#E)4cL-ZL/ZCQ)]W^MgH.W5_gR3-L
Z;Hd5MRKgX7b7:C+d/28;ICJb(Ca#4R/cWVXCW:8YXGD#2AI+-QdC7PT/]5H1e@J
Ie?,O5T-\IUTO76,3;W&CT0AAS^[HV4KdZbI^85COC)\ETEN:DD+@a1+G1X,RD[0
O&Va6O4^;DUR:O9#OMF3H>^a5f[+g(5VE(2]Z-6CfURK0V0E9/?B3WaM8eeI&H7Y
T_NNNWO^.Pe>/W_g4K2L(d[M@>FXJ=I,LCDUYM&<\0\0f(#E3bBM-;F:U^6;8C<&
f&9PJW(Q:5:>=-RY82eNLJ?>@CBWJZYI?N9<2@LB&KTD:cX(,9^<?=[&=cT#?>\&
a&WB./3-A3IQR2#S6O,_6UY:GI8WLPHX/M(T<#d5NML-RBa2^::->^TWXa>G0H\#
79B/AJ@L0,fR<N10DJFgKMB>dU0KKI3;(&O,a>OMT3B85NbWOe&S9A,Z79KEHA4(
=a@,aPGTCe[g2MEQg6/_)80cU/5K22>V/:=Q^;g;V>-.DE_\28d<J<TYWe3=5^MY
gE.JFAf\[#cR^YYeR6[-X003[B_.DIS&QY2\E&NfWI)R5<VdKD4M[R4V\[?fOd)c
-G;a0Y<@R=P[9L^(c.dQM3H1b46P(g_)ecd_19_CRB=1CXfVCXL3Dd2MLSQf0M_2
1XNI&N2fEGgM4P^CRW^0c1LXDK767X,)]?87/M2Y],N81QfXI]O0?G9@60)]6Red
O?,SPUPC&FX,5g/@/;?Og?UY-e^DV.d(/4X[L\X_=.1B0b@J8;>]W6E]>6^JKI<4
CWG4(V\U72b=SQ0=XgGN7]Z-3X0Q@4+e5\^=-6db&2D5N54SHfJC9MWZg3PCUa:R
,_HPf@E=@aOX4f50ffQ+,9KY0DK3O2S=?<HD.#OY8;5+R;>-Y7:6L1>A\TQS@YOM
eZF,0RQ,@<AagSa<.#I<];g+<)I1-Ia-@6dD8;A.Wad(5;;cBEeeRS3B);?[f1PB
gHbP-?Nd-OKaSXeGV(R-d_;V.;Xe+@^GIT(4Ia+63Qg]BROcUGe7DLL4gW62WZ)7
Q&Vb[gB1._H<2fC9>6.8bMf?V\[W.a:<@\HK=3c#M3&<38ALdNNfO^6S)37X,c.a
dYV6>gYGG8e-57/EKLBQECaGg:d_-7OCO9>NWeDbP(HRA;f(P7]TTfJWIC6)UZM1
L2XO+/E04.D.I5M;dZRbMQUD[R/VXVF7#_1aW23KO4\HT3G]<JeR31\Y:#IgcS[B
/^R@8,dcg=Q&:&He0AI5\C9<X1?fEF7(#)W6M<>.Lb<K(^PCV^9&9=7H<JJT[VA0
2XOb]CVVAIAO]a^D9_L][M99L>cI7cO+dRP1Y]P<:MPKH2IP@:f)@AbC#GWZ8PY6
W<NIFO^H>3K1<6ObVY5#I8:?,KC@H-@=dc/Ob(L_&[FEU+6W6dT:aA_Y,B(Yd_b^
V6IbTL667J5HX6]&/<V3Q[Q?9F2<c3>S,?]O_<3MQa@E5U0SNA]LaA#/T-WV\5&.
):@AcBBKE3/H-&^SU[S/U&>_cEa]>eR7Z\WF_<ae.7;\YB#OVXU0eX8f4^ZKX.E>
]2Z^JSU+OO2-WH]W0fe.)>IVHSOaaI[R>.7PWd9)U&b_S?^)NT2\-P8[4a@5W(N,
JP&cKH2R/E-\BE3>SBR+U&4A(CPXKE]UcX[5]++)dB\Q-5T5[6N)=@,GUQU]bOSX
@G0O&1f[L+U+?a,f,9/O?WAF<E+#fW>2.]cdgVU^Id>Y,=K89P+a@MB>R37N9O4:
>6\J>B=-+V\L)W.:_;OU#F(]#;><HRf)GMb9AHd_^#7/&5<d[F:-[&_#[UO\V?L7
RP?<bd>A;0.D.d5JCc6X1aR,6YbY,RQ6+1N2(]Yf5O23_#4<2\dVd:eLd2=A#=(T
<Z#_G<c=4#&[66+#K<WNWNBa<FNP55]cBN;/X0<0/I^a,[T#ae9KKcG+:=;dEEM0
L&/]J2aKUT<[ROH=F3Db69PI0WSM<<X],;2G&JK?]\@fN3#cR+cVQCf.aCM5_L:D
(1.4[I3_032(7;XHaAe7>;\;&f,;Y;f1.TF8-G&TXcUB5DPRHQ./JdA:^]IdI5[^
OZ^K-a@U]g)LIXf]KM<WO9:FO\PW7YRB+CTUdNUW>.FHD6=.[E&.\f&e6U@e8Y,?
ZZX4Z5T5JJ5#^:d_66S[(bFU)?]f^P+:1ad6e;=aZd/C]3a3\?^IUH(6[a^#XN]&
[H&Z9YK/G5V0dd/SLga<(=PTeNJMTK:.2FA@V5dF]cE6a9TFOW[^HZ;BNQ6\90]A
g&GR2-29;NV#gI0C&[?\^J_09<gZ.M]GTCQUd@KccdBfYN,AQ;4EKW;UETTNCc_]
P_[e_7Fe<#e6&1Z.X&/,cX;T,W6ZF2,3(c2TF8U[)#<C[LOJ0:dVND]/bcHG3B/,
2XA0S#=J]5BF@@=7>](:SAD4aXB&K<3c/J[6WFPbS[QbCC&;;@ddRSJ=\PeXVL__
MVN?>+@Z@8N23_+-8/7C&KBV?)0F.IceTa#(Y:],6\;@&564eQ&U0_]fMQ74H=B;
^.9>)JeRBE^Y&\;#Q(g@eA>aDR+=3H-770aTA?d-+^cbX28^/>Nd)LY,SJe_8OFa
K-->XZH)L]>,&X9JEGe-g^GYE#0ZQ/WVE_c]^bDU_,=1AgeRI4TL0W,&=#8<-WTC
DO8R.:9[7D&E0+J@356_>5_[<39OV2;]::RIEIIddd2<30-KF).=(gb(,1<3Z.Q-
\Qb&3+NO&?[XLT@(5CO&QG<Y_HS&WZVD^<KbP.V.-=H9@TEH3X./@=U]c[GI8MK2
9GN:5V=[E/6/5X#7V(U>GPB41L<E=GcG52c4KS6XM/<A>.,B6=89#\,dV-Qb+)8H
[;FT+4G@:3]L.HA.f.Z]GL&0c9_Nb>,=Jb/^UC+Ie^WN6(V+5H9;]S&5H7C/-5>M
Q(#=,2KJ=,XVg?2=BbbNIEJf4c=@]^:H2/b47:8=<6J:E0C-bdW_L4K_fOU?S-YW
9VBfG?F5cdM/<9^Q3QL#1G[XdRYZOH;@gcD_L)M]bR+8(eWc:RI^))BT9.&FXEI;
dDWQGcP;I;F[fMUHN0F(0F9S-g>=Le>cXPLVe;J#eJ&#)TY<APcTT.Y5P<dXH85?
??+_T-MVD)5,^F(/00QGgCU)DJ9cOBFBX5FK@M?d]#[SRe^]1O#W_/P?7bJ9dB^_
B2>,=V?LICDe>J@2ZG#@IcVL0\=R8fKM\F^UX5ZQLc7_+cK<cR3;F_E.SY8ZRY#Y
9f;HSA-&]VP+@H=_R[KPZ9BCaZ0b>OL1/[6MBDe:#Z7dPZ38W=;?:\3_PB^aUO+V
d&1N,/Fa_Y;TH-2MG1^eEFLaTL+9KKgUAKdN<:Z7ebc6<W]U+g,eV+>>8M2XCL^<
T2R\]04fZ?CPM-+4.:HPHN)RMHC0efg\6a8<8fU]\]+@<I.6^]+S^DA?ePa>_JfU
A?L=<fJN8/[<b4fW^BA.f2?H#V3M9C]:2P+U?b-/=JD\I6YC,+,@HB4]SXYQ8D:Z
VE\d7XI]RBD<#/X3c<_e&PaHPT)_e=9HUNc)T\AO.;PLOcT=K/ZCT[L391>[9dOF
@&cCbB0:3IGEP5T,3/H4\6UO?c3EHTI6GO[1/PAH6ZRVUFP.?;:>Y>+YL)5LOF-g
b3EbHJ2bAPQ1&8d7^-1;+L\N;e],Y&?<Z=/[<P3J9gd]/@3c_ORHH&NDg/ZMY)Y)
<=TbM9XEKUI^F-KX0X8I\EbBF(J>ac6Pb,1fF?WU#SMf49VP^8Ia5>f\cK)P52-N
)AVR/4;Q7N\L0Dgg9SD+KIB]G;.DEDL5?P-c-Wcb(IV<9b/;6O&a(<,/HT@]W2,a
&CYW\8fB0&FFQ45d=3)7QM9E:+_FG8KL&.R:/a.OR@V?51IcJQEF91?D-XgBd]cV
bbY^/4L)e(K75Ug)?G^D]YAdFPLAbCb1OR1:-J>SDSQ6I@MT1?NP:f@X3f3?5]_.
32WGYXPAFZRP5N/OK8eDgNOeRQT04aZTeYAB/-gT6^f1OEABBPGEN(8M:A)_IfWC
3V&SYC4CfJ+0fPN8+>UCa6)LP1d-()^4<bge])-QC;Q46T31#R2)?8XXT@0-B(+P
Qa]H21d#KY7f9)GcQY08,HAKZH\gS1C-4Cg-a\Z,@?02@fG>(P]/J36SWe,4?[,F
L1:P@[eHR_4R,[caXc2@FS=K=9\NR+5NM5MOF7YSRSgFJ\8f1d8b@?a2)FAad9VL
[3S-NWP-0I,[+1R;Ga>+)(2>57fI8/a,Pd(O+;fCY=A9G,V2SE^?IGSW)8)\Z,^d
V,e0?E_KfL?)2&GTIc(?^;VS.Q//(&R;(C(e<Q-T_8Q4Q/7Z1AC=/KJ?3@FdO]Ba
C7UK7D?W;RH_>F/HOJfX.Uf.fQdd<Q6VM\L8c4=Rbcc&:PcC/;dZ&M(b2fD6+dc>
c6O4cGTU^)]O06Jg^&A+D&T(^KO(:55/?MaN6QMFHK+6Q3YU7?#CQ:[ZaSf7PLCJ
R_@&GPa,8_g]SO.(\6?_(1YDVZCT5c<A7P&E^36J>,XF[F,#V:O>TR9:81?X:H#J
[.,X<.cJV2V2G[35Q;1:1?#SD:&MB:_J8))bcaQbZ><([?OJU_Y_I7bN-L&-K>]\
VWG+PT5S(&_3EENP6GK6#Ea:+eO;AQ;CX_\[MR.[SNe&H+6b9@bN>;:)eE4Se-cA
>#9@<-_T]#QXYf<YV#fJ&P7=65WA_f>O.6?@#?3+D41L^P_;+PVY&WfLFbML/?GZ
\WU3GQV#NfGa\?_#b5eW7Tbeg[f.9Z0.T+bW[g&AAAQ1N[6g\1dM9@QF[UQ14.\R
N]U\O^D[QIee>LF/T=fKTU]VJWVA8R_+Z>[;8:&RE#:S&B-T:N^HZ[U\cJ5QJM1L
+SM<Og7Lf6@IIS2f1bD,0,9^R-V2C>+IC:U_=TKM7OQ+39GK_g&:ZOIL8DWZHT2\
D6@K@f.?TC2V.E0NN??5Q45&97F_,76@RA>&@?V.CV/CZNCTS\CYL<>=-A2/)0(9
#3,NG:>^RWcQ)XW@O7I8X4[?+d)DP_\HE,E5=K6;F?7+V@&b^N:6]A/R\61;_[8P
BH7G(7V_)#OH,B;?dX_,LRHL-3/=V9fEAcL(dga6X2OY;UVLFO4YM3=0OBQ@Q;g1
3GQGYe#-AQb;cc?>eW@&+?c0?+=9e=_CSHI7^3_#NdSX\<K@+ZJBM;.]RN.<G=.g
XGNO<dC4O)S8BQ#8COc]>F1J6eMIW9Pa5NY_bEX,f9^DKGV=MR8KcPfP1.X7^,KP
eERS(J;]OAe\DTSRI;GUE>J]>+3YP7CQOVVPZ7KZ[9_C4F+S<WT=Z61BC=4ePOAM
c;?S[YL#LB&ANL-gLB)3Q?aca2#:L/2cfS)G]34#(>C0]:JG\OS>aM[_\1\IJ3]d
_(XXWE#BY6_LS&XCPH0E8X1,dWD6N_+F=1M-D+&?OaW_@SX)O3P@gAM0CN_4K1R5
\6ZA>6;MZ)XLQ\UdR7e.bAQT/]Y4=gC_LDeZO?282_AZcUI\JK3Fe#WaJ_TRM63P
TO_WF[gGc)^6@[_8#[_/+4Z0?AS1gE-5?MTaNQ-DY^@@H\^SP=8;DB(QXg;/6DU@
Y^73)3;gUeC,F>W;7cE-a]d_9PfSN+V:Gg7:AdRY3@AH[B)G40c+ZBQ10Xa_0M44
VCN^Q\4>b2#U=E++UX/bQMPU>,O^I?1\aA222TS(89;+>X]TcQ_=XB[S^H^60VC-
QB8EZUZHCV?=\RgU])?#OM8EQ+=H:0&a5.\Y:>2NCa0#ZV)]Gg>U>WEb<V7IA+K0
,17gS-Va\BDc2U_g\]Gc>=.TF&G\OUXb[S5X1O5P]E3JWB-E;.L]&2FZ,G9&#e>d
A^R<_O]d)K6,S)CH^F8Ie#B5_2L?,X\X6T#U;6Y+GeFFaFN9Z-8P=M0XD5_A;:DM
;=7g444<6VY.F2:b20dg+6333g/,#f,)NH_;BI&_ZMeDCCN,U0,:KAUBN^UE_K86
720M,8H1?FFU;C-&AFL9[K2_:&fR3SZfN?XWEgf^<Q?.SdDIe=Bb#?<.AV(\^+K3
Z2bU:>bQ&P5];&\3??Q1M_VdO?HI?;aNI0T)EYCPF]>:CN&E9D>A4A-&AgN@R7.2
bCJS;M>;PA;6I,(@Z&A02/[&OaLFa[8GWKF=<FS[cD=CTS/&Nb][CMSBZ3,[HR^X
1E>UFC6=021aN>Y[8\?O3S1?F2\MM7@)684(SM1JWfEQMcE)G-SSdPKHA-3LVU+J
[gP\H(T_)@FSA&L;-[(:\A[VBRJL>[g(3#COdL)QaXX6M.A\3=.W_R->4EM[gL#S
V-;IY:6a[81e;0<ILH4L///(15RMB3I_[d7_[IZ\gZKQJ@K5?.>fHgM4PZ0&\42F
>e56N-<I&IfK=6I2XN/2<K#@Z\cJ-4:?]8Z(Ma1-7bP:85Y-637\QUW=J>W,@V\;
=SYB:D2\I0G<+B6dc@)]UH;3N6.@JJL(L/,+A0R\NX-d5>4=(Uga_\&-35MP9K7B
O8:Rg7^7g8)eGVCXUgb,.85C.bXNH5UG5;XR+ZG/Rbc--&X04Kc7AR745?Qb[F+P
=7TUR/J]]C5_2KB4):c@[3B?Xa&G?&[P>T>CfO><Q@JT)J8,AOGcW[^1=L^M7(Y8
W-I.]f^Z#E5R:8S8;ZLe8@P#W.Mb/L4;,g12)+=B,LC=3=8SYdb54QSQ/g;M03TO
6dV(W95LFT+a#@.2T5Z4Hc.(V9=I#I09^9C-BQ9QD3HB0O?O1BXC:F4BQ_RD&Ic8
5,VU#J8_g-.C,BB.6JEV(GJ.f(H75__EXGHcc:@,_7#/YfY<fORJ?fXDUa9U7J47
)gI=_,_(7^JVAT[EZOAQ&//8F18;U,H@00c=1G#L4+5]CKJ>K[dF-;Kd1@.A-e(A
(b4B0B=PcNP[g)+:.IK8J_T7V(NLHg=UWQ5IJ.:Z2Z6NH5F75)WK__GX0&OUBZ1e
J]Z7Hgc/;YdRNS>^C&eV@g8YGOecBRR2L3-=b-VEGUH2:(^7LX#IG5=c,d?K6]M,
]5^0HOO?QR+K,@(9,KMMc7(+>9PEFYKb3.8:4RFV5WfKV\&H,YQGD76T+00BI7G\
d/7/5M0I:N+SPOBCgDaNA)(d--PJQ.,@?V8M[M@BWL?Q6LD7F[cD60;_],5CK2CL
cYHXQH46UKf+G;YSAH2LYfQ00&Wfe0#,VPVHN;,?Xd>G[Y20eKF1^UN#&X3MQ#d>
dUD.^?HVYB\/cB1,;^S2,BF]V-,85HK6:FPc[@fI9ONU>ZJHJ)50c#bMZJ,HA;g[
d,4YX358LLT]9.KT=UK5>](;Z9MMP]KWMC3][aXY0V\aF\02WHSZ1.U=eDa??\5C
)9ee2bN&Q=cHT)HXETN\MdK?\AVG(I#;8I.d.G3T^YK.KL[a18.S<6.70?\8aII_
-J;f^Q37.ecZd[4_YQF4T7=KM>b,_(SO\cL@bbR.dB+aKDdT4B0b=:[2_/f#)Bd3
XgBQ18I)/71&OQ#-^MJ.Ze<a(>?@42EZ/47^E^3S7@276CgTP?R6B9cL72-dKJ2@
e=R/)NW#eI_>YeZ)A::XfV+-0Y.SWQ,SB0OQb7ZNWK+88=75dJCZ)^8Q94?H)3^7
TCN9,.c6KGY2KNMWfL#3U@W+T=A?&+1V,48aB]?Z<7OW9QfPZS_gbU<Z=K[7=DWT
SR;?1A9,W=,HS#PZ75a+9OKBQNUM(]V5Z#Ka7;U+)Fc_O6gS3I-+0e-#9b-TQ9Gf
eN^_[6WQ&WcFI//#PCZ,DTKY2+H;I>+.BaMGH280D//7B^aU#cQX)a;X+@0Mc^DD
HN/WFI2(,87:ZV[8S=11fHX9M.25R.8RaS?__N57EYUdF:A8R<;J&(W0A7&KFd;Y
JJ#9dMPd_/O<2/1N0PadZ_TP.<Y7-L\A5cRO>fYEBP9]\:acTAV_90M/<\eN]=:W
TBA=8QQE[b+Z5<_GSB.R[I])K,X^K?9g0A4I0P?4:Nd/F?&.-TgU:a\\CKbg&[c;
dK1YfYQ-,e-Ge>80<KT^S46[#]:-EIgcNaf4DTPZ(]eVE8[EUALM:LM>f<T]MW0-
/#fc+GH-154EBFKA(NbC>?7B;4.ZXP&>E8/1<OAaLa)66+#?987Bc;&1U,C[I501
YP-T2e@b:IdZ=,3cb,Q+5KOGDS:a6:aYI82I/I<4cT/Q>])2+GJ(4-(4dMVIXZ#.
T.[/\BNf@G>UI09&_I6HX.a9cD>d6<#I>ff[D-De4dXYC(S=BROBdFcTIZ2B,Y5N
6J]?C_@IS&P3bEMLR8G)<T=@7)W/WS,(4,4/945MUPJM?-Z3XIPW/HgFT_#.BP4W
VH+:?KQGLg&/WC?S(Ea5G0d?6]GDe<CNSS#,f2d-.J-,Mac,Bgcb_C&[OZ>N5QBB
fQ_ZO/)?^YYNN^fdP>PTePdHQH#VBN)+/B]G8FL-\5gd#W))7LZ84K757:+;J5;<
f_LB5]0Sb5<G@5Jg?YG]@3@,G.&MMHJ007>aIR-cf,EM#HF>M6ESYNS<Q-=EH0ME
bZ+GI>dH/[[c(g.(&7(]6&gbd;f?LBPFId@TcW]0+ccfe8OHW9&B_;S.>SJFFBN?
LPD[52US-?Z/P@XW)K:8]4A+]&BM(QU>J3S]Q/UM\OB2aS->AN3WW)GD/LO:N/;g
_#f]=b(\YSM)>TF@5+0]=[+S5e9/a.2?1:7<Q7,.@(H<&\_1[0563BWE;+ER;MM<
SGUI>4N9>+B8bXKHJ#_<g>A^8WURb8gL296;/dQ.aCA=_S3_TMQcffUX:)Kg:c,Z
\/9]W76;,C^dGV?RN]JE_&/#6f[8X8?+:b2]:@@-EH3C9:e9=5e=AfR8N1M[,JP[
_>.L)+E&-[@A\1?=7G-#<GbX?90I-.L2@dL;^\/>PeBE7IF>X7GS8PP:9aU_L/a0
&Yc0c=5XRZ+<SfWP0\X9B4#dc\F+O>eQ63VCN5]^(0,&N?4&2)J77D>0?c4C[&>W
CQHbNO40cg-O?5D63_->8ZO-fF9;eW<]fg9/8),:1EQ4g<:<)4a<5OAL=4U1JZ6Y
ZW9JP2YG4<Q,P-AJ-aK=MCSI5Rd8MD3UF8[/eb?;]-2T.@,IGcc8=NY9PU])eRdO
cO5H^g1OUbOQX2,VKUA8CfNG3YUXLL62Wf/+\X5\a.=US3bCEDW(\RY)4(DV..+M
(?U0Ga:WOWT(=#E3(:g(a,E>[-UFP+3f4[?Q:RcS^OY3_F)DORf85GH\:NAC+_49
YIgJc<I(d6.0>NRe\#Ia.^S^UB:O>=7aeZQaISGHKYY7eO<]Y2Q^M0+Ef?JAda<g
R&.gSF4a:]>&2L(3H2I2)/Y8:FL+B\P-dO^T2&3<eXP6Z_DIY:4JI.BLAB=QAC)1
0g[)6,\M/WNN>DJKSI#[a(;dYD&5J7O]S-OV.?<BMbSHM-?:d;\9gR&XBYHZR;GV
J&5B/SNMJ9N&Q7TR(]T<YeQab4MM6RLVL;T0S9]3V<d@>KZZf#;a8M6a(CE.5J@6
9<]PgEI&ON0TA,TO\#g8Ac0UQ4D<JeJb_N73g3(_>W;;5aDXCOOY,?(/HXBF3P6+
:RDU/=#=E(9W1,(F<?5WM3:a>>791TM;B?2#POZF0#^-.;#^YWXHTXc@^ZI>e.+?
DB?F(1YK?,/HTN3;Ca.R/,JRLSDL>TSFZ:WQ2@gJ;KJW0EM:b)d&D.eV\VMOce0/
E7ZN&)f.QS^]=\g.cG^Cg1[U[HEMY8^@C&JaDB?)1?T\:^3-4OJ/A0f(M<a8d@^\
6ZgM??M]:#a\^-),5+9IU?65Lba^DEO1S0Sdb7).Z>Y_.:(&cFd^5fP4B/QA^@cF
@+]1D+DG,Y46E=7=U4N>0&E4D<C4@KFZT)S0L?_-3gR8D:;C7KB)NP1R6_<@)P#F
6J;1SN/=GAGLMZKB9EYB0XK?NB9MfG3;DTDKYEZ2@aH-NJ65^4#X&MCHMH)0M_H>
SgF,XS@E:1/7bI<MQ+WN)U.6;^H_&)F\Y[L(KWVVV,+>]&1GEfWDV[DNOJ8)2ae.
?bBa[O^AJ_H7f>d2BOX[fHJ)/\>-]cR3X(K].8:cZ.RTK.NQ+6C3[B2e/G@K\>_U
RO[98XHTE_-2.04ZN)E8bH.4<FB3.D#>dA.<gN-G>RfN]dTK7;HT[-cWH,KDO?Rf
W#YSNZ@^CFdHc=AHSLY8abb8#CT3/T&5<0A=.KSI,AY=d<R,fP>P_Z?U27JcHgO\
eVWCIZ5V(5cYHLF]ROSSJJOf27:X>R14,cP0[V41&L_cOWHI)Q\K,)&E0I@5JFa[
TCS7B/M<^fZIPQN-94(PJIb6ed>==c0D@3U.&\fQTCOY96P\P9a,D^B<.]T&H)];
S-#F_7e[BE---U-.R1:KEXBE-QW&NZ4\b7BAXDFb;BN;6EB-S\/?13b&NE<?1FY>
QG4-&&c96Z4M@4.UZ(PVcY9XRCGf^ZY#I[6:5J7N#9TGZJ,gbZ@NO2B3HKR.5#d3
EN2P,?>87gP+)+DMHB-Z^R(fe7DBE,3+fQ@QaaR3488ZWT@cf67G1)]TY9]af&)&
a3+V)7;7\O\IZ..>>+\)&I[6F)7KQKZA1>:b82#X/&a>TX;AV#[(=GfRX4ScT8(9
AD#Ha(8ELTVLX-IPLc;82LXELZEZQUb4U_XF+XBIaHM;;9])LJEQD=?\8Q0NRgV-
A+)D7EY,BV,??G5)Qd73bgeIa&g-6IbNCc\2:G8a>GaTK+O+CME1=O3cCB^SL6O.
QNTK+<6(f5M&7d#f>F)Mf=H0\@AEYcTCYC]GUKe^;&1JWI5NZ/842C;;_IP886N0
MS[cScfA]9T.?PX3gSJ5M3;-.b&:O5f.)4_&&@fVJ;7E:([62A;]6HeaH4A_&dMf
O^.]HEb?B)#VeWTE3>?cAN8;QaKO8,bZB+7E6.X[^M40E=[PY>^c^#L[JT3>MEL<
3Cb@Pb\>Q?T<PLXXE]:Va5XZ(R6:ELJ#f.J/]&fZ7BeUc79&8[EP=Y:6^O85+3\e
SD5&.&I3K)M_G>I,A&GDXDYMI=P+cC5#3PdI1e5C+VBAY^@N?\07EG7H@E:\fLYC
YZT?R/@WL:Zg?L\6FRG]&43d_HE;0[>(N8WATZfIB+5]4J=8CI3_-7dVgg)K&D@O
1CgSN<UU8U4CVR0ebU?9)G;1A7\?32f/8T86([\8a[?XE^W.4e[f7^_07^EA3VB+
S5)/XH/eWRS3#Hc36WZ5FZ;#1cL5<6cZ)G.,I6DBeae+EDU2;Kd>JT7L3BL4D]D5
C]fg7YUXAFX9c7P;+XU&]d?JG^(_:HdV01JM_1+^E#&Y4NJ/T5;P5:.ge#8MINAP
SUFI;6?S3HCH4K^LUM^OIYJAG\6>.XU/Ff8VH:\<#CJ3Z=0JEbf-=E\CZ5:9?.E=
@29W6fb6CS>@AO_^_.8UQe<9=bgC,Y<IN9XB<359WgHF#Z-8cWfK4C@,7KC_&><0
BV^bU,(J7&+4e/-@NF7]EYLB=[eDfA#K^>:S[+.[<T#@C_DL?=[CYcI6.3-fbT_a
F8MW9S_b4BN6\&R[(g/8A/;7<&(4&2])cQ58QE/e(LI3^ST5X9V=WFLWHPCEQ<J2
/3Z:&744^WT>@fJb9_9I+C_B)AYDGVT,YU&(aXMWC+Vf.N/=B1]]ND0DA;[:6L6M
C(3/KOdWQI^NdC38<cME:AECPA.RJSf\cKW2JPY&J[XRf7;S\,VE(//C^O6S2<L[
[KYMY2gg4<&>E[HcPPE/9I.R:SDXC\aX5]W6:](f9^:QA,F7NB2D4f8DFe)?JN<A
&/:19>8PS:P,G/[DA^P7RMRN;-af7@ZR4.2JU,^b7,>UZc1PF(0>><c6=R2C8O,]
V<?N]W9[O;MVfG(.b=E^1Y]CC0A,6H2:(QaS3;B,(b);AFKK9G-UReCL+1[.feOU
SS4\@RA<Vd4dd_=YK0K,VN&gI:Q+<f_JZe]Q-QX;TN/IR2ZLe#6\T=LN(B@bO)2g
c_bM7WA^4OT[_[E-8DJ:VLg3TZ./\/D@(ZaeJ7M_A,&fYPbgKV2/2\2F1[T4IaFb
00F-Z4+,.RGA>N9Qg<ebLC)+RLD_TLgOY<c,WgC2S863?1H87@XQ=eD;QDK,gFNN
1f0g4_efEd1_]Kd,?0I,^,8;XT;a(78=Y,aF_LK<Y_f:5M^&N.N.DN,WRd[<V1?)
\a0_+:0B)3Rge41#=)Q/6/DbI<,#.HIAGN@P)=WV^ce,Vb3U)KeZEbNaXM-(\2<P
/)cDVG<B\+0a.X3K-eVZB(Xe#A&O\bO=FDRGfAUEZK3RXZG5+7f]<H(+4>>TP10T
+]HCbG&IOPC_bQ.SDDVfBc5+g-dP[H292VZDL=L^^7-5P8.]U-;[RFW([7+aZ,]R
eM+JPF4S?:[NPbO>OU.OT;a0.XcPGYNI?8-cEGQN2#\QVb;(^V\JgT#V]FXQZW05
+-QJgeQSc_&OM6#+R/HP?&fc9Y.[;O18QTBS)K2^V54][D;(RN;Y2^,b;fOC>/Q(
,S7Qd),\E,1Y-]4=YGSPJ;:VU<5S]ZD:cW2W4U]1Cd<ADXFGXXRa:CGb8,)3US.)
1F&?5>-+GDP?158:MME>.O\)\7/&9U#,gO[cT@f90&J-d#A2DDeZ,<W^a\O.OTP>
=\Q1eD^2;458abd3&N-e^4]\QgT</]I17:S3)<<>AYAXB#Ab1NMN@-<<VUTWS4X-
eL792F/FP(^?Y785@C,Le-&<cJ;UFJ-8M94W^B3)g[#4gUe2LbXc;S2bE4KZS(87
16B_TSTX+A/AP;@c1_8U=ND,/PIN+K@6Dc8KJEK@1QdZ#N?\6/eU>LU#d-,F;>AM
5,P^4J19?O#Oeb&UZf5X6U;9fO_3C.OR2g&aY;0B@>c]JFQ-5@DD0^)C8)fD_<2R
C8<]PJ0NR?17A)a[]4DcMM](]N,dK/[S;>3V;4IJ,W)&NO,W)SLW<.^+JKXUaW/C
&_=52(<+O0?ZCA9=1bRF]ALY0HS55e)@<^Ca,SM,SPQB[b+D7<a^^7W8b,W-]2e)
<#Y8+DdQ8fdcP\7Me&?9THBUS?J-=+;9=LKCG&-2Q(?_,4T]OLFW/Q\M:cf@M_VA
3NBe4<C_[.J5f,DC^@QPBA.9D^)CH^=<(P/CbT.9(b;V].[QBD,]3_)=46<U11+L
U2[M^1;A8I1eeCfEd>8K.<#U]B)S-f+3TBeDLGD+>B3-I(/F)XV,BFcIDcO.MSR<
<)AO<#QNJ_U9QR(?UdMWNM(0L.SLGS4\ef5>A:SAZ_WBJ-WI2C-Gc143QLCcCVBW
]<8]e2U5E[-I7NHIaHE&Ec?bNG3?=L.(IdQSJ_d)+1\e1cNd#?N2+GQKKGbY@b?\
@/c]CLPX=E[]ZOF#D;)GGT?;^/8#+N,YY=(0\2O@75d]UYA<;VdbA(-NU,Z;E)0=
^bTH<@EQ9Z)eBF76-GERZ(M?B1X^=J09d@8dg:RFH^QI#\K)<DY?^S#OYH+<8ZNK
.S_Z\MC>3_4g)eOINF<F;XaY43/KVFE]+?Z&e9]O?ac&J)g#J:@=U[7[2I[TI.<>
(CUD>P\J-)0;:Q;LSbdJ+7ACL+ZXBeTK<@c,2E9]E7beZ;[LR7_@C7LL\M6DK-G?
E9V51^/VU9>J^O/N=9^P6189Pg[9Rf7#H_^0^\./-ZCADB\HD0O#DZ^J+_PIYWg0
Y#2<HFQ=CHbaO[OZ6EQSG<&bI(;6)<A57>3L2)\DgU-;.L\0.J-&GId@D5HWGdeQ
[JfO^N9+cE=W-[[HU4FE-9>V:SN57SQC&H.5R4OW-/06>),@;KcSG9X,1S?(7@Z/
:RNSfgN[QZfP)fL20A7X&(4/2X@KVN8eEd(6[?,)5LG6?4(P-=0,cF_@6+90dc;-
;7W+W&[IV))=TG?KNgUVB7=4fHba1&5@=+E7MVV-F)2MP2-K=4PU1AHD;94gXT,)
Qeg@:?O:,eFJ(&/,>Ef0bQ-G-D3[)P1]4-Q;JQS=.<W2,E\cLOQ;]YX[D_1+bS--
2Z,Ab9&)?YY3fDL62bCHGK\dg?)cX_+Vg[R0VS;@2R..0A(PZZ9+CULT^((\OeEd
O-eCRULW4/fA^-:G&NBLV-MZ:>U)UYE+[H[?6bA/<CU#CCDNd)J0F+H/I\5M9,_:
PP:UW9@XFO=M[0QBW+;QU&6+@J/U_eITM(f6eJTLO/VX0aPA;ZC-(2:T1W>EVRIB
.A:MY)CAW>>KVZd,BgZ\?Q58JPacFV)FEQ+,4/XbVJ>9W8GAD].+^;Z&5I-&Na7\
&bBP=SK\+3_U07N]FIf43d0d.c>VZ?2Z?_R&(fG]Z@_O5a^Y-0aX[bO_/#_ZQHR?
,[OLSBGeKaE3+-NJF442\=^\BK)W];F]_@(R&8^>G>-L^e,\V#9aS10cHWHT_e1[
FY6RJZ#&aD\?I>]<24,#?1-T>XB5e^a-D&VW?aT56FBOdQ/9A+11#;5Q;:(3SG/@
R^8.J8(TMQe_N14Y2fVB]QX/4MVT6\<(KP,8A3MWW2\6cK@X-C+Y1YZgI9SfZXO:
UAcO65H6#]cGIC3T9/,E)3d];2,D#@K6JX3)JP3M>93;0YBfecX90Ic)d2?aG.GD
3c@gfXIL?Re<NEXFYaQNY^Z9E#5=@4GB-E3BaacIVBJT4-g?XC/?GR=46<HGI8WV
PP2^g1SD]5;],DCeO&#/HfM=\gaf(4A06M;OI(Y(B<+@N.2N<YSV?VQV-dBSW>_:
4^D8ES;NJT2KdNI3=[I\)0>)R+M2@VcS.K4YDI_-DP1X1C<SI+)S?;dE19/B.Q#a
+a(TW?7Tf<TIEaY3(F#If^Q>0R)V-C0gO#TRF[CL)I_OeYg.9,]V&P=JEG.-/bWU
[c#\RZ+O(&:UbDU:aZ299B[f?[eS-\;AV#@[?2(U8V^HeHPfVREGb99J.@/A8Ld4
.76bT=S+/-(M/H:3?)c8JH:J0f<REQ6[N,.ZQFdC.FX@c(R=-,Z;V4\MSC,L;LNI
[4VLc?9a-Y^\_;RQX#F9/O[9E&<CcaR_e\a8d&3;8&EQ3&:?YEaMF.VW60(f)5\[
&BWMUF0^MA;:^G8eE701TH+,(BcS>B,ZdK(-U((VS\\1a:d8/ZPe0U@MHCQfEJBZ
A?3.WRG<_2[1_)/g@^D^#cA+UFf^K7DB.OE/&U,]MTd-9.8M9)Ma8WD=UQbQA;14
@:0M;M/OW7K,Y;#fd0QF-BQFK3/bXCaL<FB6HgTE/\OXXEOL>b29Y&Wb&/DC,+WT
BSZ9:M(\)Uc6MZSATPHE]98;&Z^XgbVGTW<fN-SH<<-,?([I1O]X?4/TTaEb_GAX
HgcX-eB<FYg]/:HfX1^-O.dZ#Pa@82Z,GM>&eBd;e_O3LU]Md44ecAdGN1@6?^6V
K/PAQ<^R.(FdL47NDJ7Z4-N;,/1Z\X_ZJREM+W)QU4(KTa+CD1>a(<c38[@3QA6L
c@)):.-/3GLTMBd@\[;9RYLg)\V4>f>//2NF6S/G][?Q2RaPFgX^B>&<ACF8].(e
I0/DNY<c+.6(R#QHBQP\RQV\GESDGLY-67/+\=gc/YI7Y#a\,VBAcNW^#)(NMXK,
F^JBQcc8FeG?71R:_L._E-QZ+&1>F1,I7T@\AMAV/e;JW:74?SRZPI.ZUJEWGER]
IJ@OZ,OE:M)QQ:\+==1IZ>SCbSJO^WH,_,10]P3K<TL-ZYAJ@_e5)eOROR@1&^PV
aY=cF@:NFF&/[cRWBJ?)Fcg=DDNHF+5XV6KgM/<&N@F__I9/WH\)d:J/T/KQScNF
5&4Af_;M&5@(A?M5(KXg+L.f(D-7AK(.]B0]gfaHJ:O\;a\WZgG2S54UKCY?b]\,
Da4KEK[9ET7:^0;)),U[#05KHXH@Z[)4Y+W;G;0A)JEbWc3O?YJ5<G@NE2Q/BYS_
(c+TV&L^;cRRP&C0=YPUAg//1H>5+K^fa.C_g)e,@(/A:DP8H0E;D/ga03T(dS;f
->)61J(#UBXN^MG])N18VfcP?&6XL(S>KYK<VNdc2VfK@7G9RPIObFGAL43X.O0G
7O>6da7>CB3aV;;C+C]]X);D5,5KR(((@ALN79\6@9X_M;PCbcH:[.@MWa#5GF,<
6=F1-T7LD^4G^I>-270(D=7>]?3g^L4)].JPZ\0eZ8cbG8P53\@Q-@9C@7b_CG\,
^KS:>f50Z(]-S:#GK>/>0_dcWTRf&H<&866N]0[M:6S_?\9(/D.]UH:KbF:a)f3U
54THLgQ?KC<+Z8_g)aA4_L<]X#>UXf]27Y=T2V2E[-I5J:K7\6.ODT2B(@KBV^4Q
SId]GPF6DUa#@Dd<[XN#(C#-#>LBdUVZPTW#aF##@:\X=VH4D4TET-A0+LX7eDQ+
(XR/V]UH[@XUJ;bU+<(T4CC+DR+2Z]#Q25,1Kd&Q-]?E?/JbEeRa:#9b3VHZ.KHG
&)#\UUWeW74EUADKQ]_,&A<EAP-4.MNd;ST1H9b-#35bJVP[9.X&M_ACFM),-ZW8
)^K/?[GWWL2d.9e+gZCM9RXNT<BK;V>+<a&+dV?UMD&fgT_F=.bJPJe&W+UJZZ)(
(DA,-;-.,-3]bFK[,IZ;,1R^&YC;RfHRDJZ\6.(X&N^&;Y.^KS&-&GPg3P(7QG4R
5]d[?eDLb.:TC;H@56;H\9EfS,-I(c7TaHf];3)(ef&#^U>^00X4+-B&0(/\1aQF
R-^e\g/<YVLP,1HF+(IMTEW1/b]V^4F:PIbXXI,e,A0RJ:;]#WMg,]@HT4VA0H:@
-6XL&KO/dW_Ye?/c..A,V5^;;BX](9(M0ZEIgR=a2&D)_+N,U-AFGXZT^A99bZf#
9f0V8b0SMNc@/>?MUZUXdZ/16[HB[@O^Y\E:W]LaK:BIcO\LNfY.2HUU9\Q\&R1M
/Ne7J]B]./9U<&c0ZZ>Tc\4QK,)P<AP?(3W-F&,PdH5HSLd=Y+gR.LJ]NJ(SJ]VH
PaJ;Va,)V@GQU2SQZ\A[cG:NaSM369TE@3\.#O^-41ULb?fLOTAE,EZ]bR0ZBLTU
9>/&FW2Q8A[]c1a112WY]_7>S+.3g;/6aaF@W=-VaMV_.]:3-?Y0Y;0QB4U2/]?c
]T.7);.EP)>5HIVI1QE+^\.OS.C2QA(KM3)YITa)^bB4B0Pa^c88<X6[K(Y]IH<D
PVAf(A?.1AM;Y-:R67)]MN)D7SZcN3W+VR@33FMKc5[:8K<e0a[2G^CZID.81Kb7
\OEgUTI.=cWZL4U1-BMaK7XJ>F-:ALK#O:aXfc86AL2MA6LGV8,Y@F\gMLABL+f@
?bfSfP;#]Ef<1\+8J<HI3;c\>M&\=S4?P>b<7,_NFb0\1AEP0#T7O0735,G?E/5b
9;f[_J>cb&&>_\f9604\P,&JP]_a;-eBdLL+YAS;]&M=6K_^<]#ca]S;MCE9RUE@
g;1L2O,S\D4G;:55B4)]U)/YQH+RBL9^BY5<4YC&9-V630T<@-6)@TY>K-B1#?@T
^EdWCFLV\dC=0MO]1=<.WQCOUV6E>O<g+OEZ@JTH(S<g28G,4SYFG^ES+d90K:)\
d0[eQ#II+8RAAbU62HT<YCL_0CG&JUB7Z?42OR&.@b\QS4O()224CJY9/+8/B+2S
)Q01[7<Dee&P1F8#eSEWQEJZ[5@6Y-])bBYeH^[-FY[Ld::<:I;)gINZg&#?3XS<
:UWeN;\&0caKNHgFB[I_L@0R5,SfeU9c:7a-ONN-P;B]W3MWI&g-2/#7>GdAMaI8
65d)ObW;3G4WRL?/F2/(6c]ICUJPg-LCQ#1301PT_0d]Ge=2f44IFe33:=ZRBf4b
E-BPY(BTT^f78c:R&\>\#P9J?SKO]c[NA_H+BCS-fK5,ESg.-(#9-6\?:0REKCKe
U2LGBcc0[G9;dfYE3b-E/-[aaY^8aOLBE3d1:fAZL5;:D?;#/L;<_U)Y61f#04IM
+(\K6+?U_EMLVS#]3(L&T^APgd7[)YC71d2cK9<RaR1U_QK>:ZP4R8egXWIgb=g6
^B#]YSE@E(2a/25:HLM;O5,N#[NU;_+A_1T8DYKOQ\3K(6H/IO]LH;_K\<WfNCG,
fd[MA7W+[<Z;<4Z]:SZ316>8DU1NZS@0<a(6S>7=TbW+VFZJHTZd&_Gf=<Sfa(/G
>]WBIb71-1L6fV<+OU#]L29CKefS5U1f@_;dPMTPA<X2YN>?&GYLbI(@[)dIF(Xg
ENP]Lf-2c]):IM58\2JHKG\Zd8:A]PQB1EJW;3_NU<R\f_,-JgCG=\?.QGC]9NR?
1;;@-W,OM^CF;/[^Me]CLW5ebF6\KEgMB.WAWB,.Ma9KE116Ke86L9M_E0IeI;67
D.7#Q@D;IeK2bOeU6SL7RfEI#;&.Va:&J-20LE?,&1b;]A<X#Q&@2P(UeN<3<G++
DV7LUB4(bFMRGMAM5bXFNW594cLFKf:+Ec,T:bR)-X@Q7L/L9-T=X-8W]Cd6P+4]
D7DR^.ZIRU3S/.DPR]JEDZRNMGG-H<OYfMGS;K&\RHB78)9+6ZQ(9F4U[V?&PH8L
Pb-IRc72^S.NFJcF0FNV7agfeI2T:g(.BEQQVIe2N+PQ;0J(M[IV_Y(@Yd<?S9Z>
ANaXJH@9)_4cVc216d-IfeW\=6fe3Q=)(WE+g<&@>QOf>M8DT3e9JKJT44<+_<P9
Re7=P>QBf5,<8BXHXgJL&)NSV\<+ZUB_97fCVIA\VR6=N=bZ7F[\8,S[W@B<B6(#
(7HOUA>E7ZG(>LCP4[=1g.I)E)^DA0DDLDWLBR1HLZ722.3Icc=)#.Wa0)?U<&dd
4SLe4IVV8SGYMbZ^OU2)9VS@ZDM32A0^eY4P]Bb+W;:@:&K)T>Y:AgP<UH/#238N
9\O1F[L2IR2+VAUefS:05a_9)?@/3+)gg3.)#HIQ7,7^^5W1?RWaK5F;VDf?U[OP
gD+EeM>H8,B=PN\_N1^9^2/e\4+acY_fOHJS[/aZ6d6FP2R3/S:dgYUX1S3>Q6XU
@V?R<W@DWL56#QQH.1?\A(eMcKT?&1C#dV@ZgTeJ@JJON=<8=g@Y6\644T&)Y)<(
De+.N6JJUWGQJ@CG]LR_X#9DfNJb1M6La\f7KV#WKLNBQU<Mf1E7(S4X(d93gBI@
0A\9f?AQRdTCQY<@OcCR2DF\8EZEc&/)6RBZ<6TH6I&>/5DXeY(]-X]?WC3I74I^
6:LX>6_KQFX(&N#efDa1ed+>+eRd133(RK&+6_5YP=I9_M3C:0M6BX1J=#Gf#Wf#
g-K<ON\R=6SQ8A&6\-M;+aN(+bMS+R,Y5,1G(?=#ZJ@C\G7N9?RXc>_<&@WX8Z,<
R9CSI[6CW-:_d+:[<+0Ogef:Z/E+a5-=0I]-3AKH?d21f^0dT-Me0;X[>#-]7:&]
.c&[,c@OcX0EdeUU8P3FG,f_XZbJ9NW5Z&O)ce#bO3=D>Lb7J)\X_FAcD[1@#bDY
^_<fXK_Q)_6E,SBOA0.WeLW?(+KC.AUg,&ISJ5XT.e5IL4XbePYb)<]E>5U;1Lg+
2>+V\Y.C8@&3TDG;((53Z)La?@GfPS/-PHR4NA(=U<7I6c42b5086?2C:Y\KLF2C
P65Q.UO;<77MWS.\X7A__9ULOeP1>#^T0\?OU2DIIZVR#A(RACJ7&[M9RV+8DNQ+
>b3QG9.@_^>/9RV8QZQ<B@?La_JOFC71;XY.E6gf-a8_Y[180KBKC^S7b3,I:6Ed
K^e/;bgT#SG6eCa5-:6O[-&VRA._LfOPXML9QJ9,_N>/8:M9e7+4Ma()4E4Z=]Ca
cZ@(_eaK^=OKNeGSMQ0?I&+fa;.P2I,K.7_NLc+WVF@93+#QID1E/<UY-f<M1\5\
_T4a]DOc<ZKW:0X8cUgNG=VOFW^e_3VIRdb5]aJdIR=?.QIG)7N/9&ML:E[8GN9g
d9@U9#J@41>.F6PA<?KQ2b(S?fCT/)-)5HRM,0(&K?F=@QP#7[V8]2&AHeddL<I;
0H)P7:6OP3HWK)X)6LE50DI@OVI)1#_4:)\U/M)PCW&fK?FaD1dB8CF)Td],9P^&
=T?3[,BQ<:;/>f#Rc@4?+bg\CK1?SG^)POA:-I4.2:HfF-b+;UcU2^93&1@e>,bD
^89IcaNAZENcL@JT8LOR_Ud)_.P)WZ^^PBSeDBS^]>./\+IC?FJ(S-MBZdD(^:/V
^4Ee/>\Bc=]STP3P52/^=8P3PX/a-DU2Ma/IBTFJG4(KF[gC/_&V28aT^eI(=Qg\
G0DSRW8T+TF/(Z6?=FQ-ZO3B_Rag5&&>^4]42/0(g7_-S^R:K=@]>F4DcE8)dLaO
fHSS(:,STc<f7WgEE-(L(EeDMVL#/c-XdI?BNK?:)QaWceE2^.:E?IK\9O\\>8[:
ccPR_dR#JMJa[UcU:>RB+.=9Y+9+2S_PQ&68]ca63+5T/()..Mbg;Q&)?UZ7HY(R
P4f1]>.HUU@g03SJFBP+8N0JON1WT70#9;<Bc3&QN)=6PRI=U6?LMeG+97CBR>Xc
LIN(\179D+MRg6dK-N((CB=#4aCVZX?UeOa?U)O<7=,bPgeF1[=+(e1M:MJ,&Od8
cCBGMYN^O0[CF]AIT7)1\P)c7F#:_;N.\&]9._OT&D&U;TH=bFgF>:7)X]Q[E:A+
?ZK8\Q4eB24I=YZTe3U-?M]_?2XUH8,4DX:fgY^d2XfSVHKQ1GfQKV@dQE3?cWM3
3U,LM]>;2389&DTZaHd51c<8YY/RNU.&R_S1];9TcX00ARUY<fddZfbFdI_<R,DR
I4K_7T]53_^;d;d?,.1.]J0GZ^/gII<QJK5@^&F>9[Kc7:FYI+5B8-^#:c1)Z4:I
EP&BZ^=N;QXK?]+U#[>LZB;PWJ1P[ZG&#e.;7eZ2QAIZRK@VeeKc4aLBG^?9gYN9
W[W802JJ009B?C[H]Ua03@ac8IG\1Ve3XNQ@2._&gYdRZ?6)bc<P?YL+3ECELC-9
K(_#A9UOG<<(P?&C.Hd5<_X7)C]+6+AD8#NQaQ=KfI1b<gf1F@2&?VK_MI&D#A1N
,4M^c:OIGWg2NUA)\25MU^3<FM]dP&[DBYLId-?a+S54#R\FD.955+/D:)OMDg;,
CC[E5OJg?O\&UXI,OUUKg<a[F>bZ?cT5]GXA5_E/?I+7/)XGH_9=>U[<C+3(Z3U8
<5gNY^9\0=dU4F:Wc#+-?3(DDTA\5\c]fGT)?\S3>8&0Nb6SZIB3JAPfWCDDEH.4
/HKCA&2b@Z=OF)J1&QE^/W-cgGSB=.\6^0LfZW9b^9-)\YfQM3QB1]5R?;4f=P]#
\-@C3/f[Q&CT\A]C1/L7=Q#Z):U[SY)[MT33Pa?K/#32^XA/VXT9bGD=4O9SWe3f
P8Z<XJT[I;7\XK<d;KFBea@Fb.IT<=eXV\8V+AYN&D<=9+Ic>Z,2&RFTJfFI[<B#
A<@O/2a3](4IFE.Ud?PEW8_>2?NO>=O8/E.gTCSOd@T<T2J)=4fZ4Z@^5UQFSG1P
4^G]<f]0&,UR[b1d8[fYGTQ2PY@+a89CdZGC<@#6>-V?_dM]^f9Nf[?G\e(L7C(c
5?1<6E6VL(AY(:>2<XD@7Q-,DAP6=C\d<0RE],17X[T=24&aWSE,;U[MH7G@4?)6
Y^\7eV_Xd^2.6;83B-AdDdUEDOK_3?S3M1#:T2?/XI\4d,0:P7fF+ePFNNT:2RY9
7AOUZ1+TQJAW:J/PWD+#HS=[9+K.>cIa8J-X6+fb70Mc@4bLQ#Sb6g8N4BZOYC5f
8X3W81;7URFgZNPO&+7C(&Ef/C>a8=-NV@9L_^Ig#-27^I?dCaP?PD5H9P1dS9/Z
G0339WDQ\fMK@;)JA,Z8b5?\\D/[IG<aU29Y:Z-G4/d:@:GT1aSM)c&H:?IL>WH&
KXb)G-UGOU:)(VA6)52E_;[5F8V]D/MCRS+e:?LU:@Q&1V][ZDF0+Jf\:E:(-JV0
R&gX)-Ec.EA59FD=Id,M?dQC>CB<X/-aD(aI,&<;e-aNXgUTTf=Z](YP70@,c_YV
,afIPBS>6/CM#eG&J,FNFI+Z.OWaU@->[HZ&F>\)EUSSeLK9.[ZY1F&+7d4#O#T<
C46EEae=U_Q/Q-)=C:I1_5:+dK)^7N:#B8g9DC+UKHHX(IP_8eOD@g?YRD@3N6J6
:YGHKM=D[D/<9T:J>;ONW3P1FN&c1d+UBeR+5X-,JQBMWAf)Sg&L5/PRK8]daN09
D)3U-dI1Ha[>fPF+Z(5K3@LJL8e,Bb8^004^=YC.I&.KWC;C=4<DJD9V7D/D]O+X
JcD8/PXfO:8OBB:?(.TZQ>XH+(PM+<AU,f9[<D&JFR7PTGQeV51ME-/Y]EN84H+f
JV:)^fG[0XW[#c6Z44U?LF]TMg8fR?f);-A7e15f/7PT-c1gCd)\AS\#<dQ^eX8B
]a=W0d(M>-N@>J4+Y)YeM>_\1]9SWEAGJJ]&</0::R8,WDE3X@?(TF\edS6[DM<W
P>6JC\(]<Hg\K,O:5f+#>:199DPQ>\d.O5_-,dg0THMDI_7QDY:.=,fN#1Z&@U<d
W9B-E?-LIU5P.Oag4\[K0ePP])R==B?N2eG.8+3_RRf529Z?&6419b_Nf#dXKfL3
2dP3H=1.W+JU5R.).c3SQ1-\Jb>95\cKKf,IZe;?0MfeILDH]1BKfTA^T>?P)^CR
4##5SD9f)-ZCE,0SB7_Be#?V1BZ20f0Qd?a[#=c0]@AN3YQ[7GY,WVO23</dKf0W
]4c@geBfJ)V@RT:JV^4OHSZe7XbM==33>M29<Tc134BJR23EC?ZR(<LH.:A.]A^0
&KWD^6\>\2Ua\4.JTN\2;c&8J&_9P&:VEgN,aGP04ZK754CA[XYgFc#-81E)Bc)0
];E)FU<MP#A1P+IOPaCL^\;B1O\ZZ7fR@]M6&5+Ye)?],Zf]9LQB\JG@>T>+U2(f
2?+\-UPM^J]5KTR#;5G2?TNb&FX#)XZ6,VB5IP3ae=AZ^;XJCXe80>[fK:\K=<=(
]6JU8fc5H<b=)BPLWHVOZFPM-O-+W5#Q^.GBYQfSV02BN9NAL3?A9SMfL?XA3:Ma
;Ke5\UAg@4(:6VRgKRQLO<HbCV5L-e;_NDf-gV)@P0]>f1\d#\=.MFD.AXD4@[HX
B_.3])O_M]eeL,&-:JH-WYLM^JY,WaVa7=30.LYNT=L;P(F9.0#).,9A7[e58NT/
Y@[eN[^:PP[6[@4^+-1]C>;\EVe5NH#W?0:JE#^2?T9Q;9Y37R.WcN&+7K.JEANG
d=_:GL+K7KQ6UL4CMY[UCIGMF^\RXNV=IG]7X9EeIWI+IV8VdLF=@g0WdH40NA[D
/87b.<.g-:HN^82]DJG=,<AdX/1/,LK<cKU9):g^Y5N7V/H3)UI0MLY@2),4&1f-
^a[OZ)I^MNOZ\IVNOdB1JcIY;8G4Y-;8/e<Pb+P_FLT:YR3C13K5,:\\\+Ua=;1Y
8:5PNN7fdb_>-1VV-J^5)?_43]RCV87-Ka6Y_6.-C[#O#R8N])K&-3+.Y8AC?W87
DMa()R[65QJOLA_]8P8IJA/A=T=4NGN(AI1afPO&)LP0eCK/[8aB>c5X_U=7C&XQ
[#_Y8DN4-IYZTC_SZ&T@=TQS([T4;YTac[#))D5_aBfQ@#c.KH4Y9<KWQE^P,@CB
aN]Hg1&[fEJW@<PRL1D+39LJ1=MDZ=?Ug/EV^>,.42KMNXNTKFT5=+A39cG.&V8)
,P-PUY2T3.E7UPX;:0/4-V^@YScaOY,?(@<EGI)HOI6U(O+a?BQaX(JX[@7\<@-a
gCRS#-47YDAS]&Nf21cI87+[0Dd&Qdf&Kf3ecNMX3f.ReO?^ZM<\&8M/5QOLG(=Q
)8OWI-JA>a2P&eT7A#P,fSW0A0A;]07(ALTG/>2b#HBbX#88e1+BIF,&J]N6aIR#
EQ,33^#GDE8#LEf;a8J#>8TLDWgDZfTKDDaSN=ff2ZD,a0X_N#Lab.U-[0^)0P6+
LX03gC]\]C^fU[N:D#>IO,8\(<KDM^J@bRf-57;P=:J-QP<M][O>F6+IC&YZX]bY
Tb7R42MTSbD5YaVPRfQ,?\R@+]/=44>bWc/,J)&/:OOF[ffb[:9RTeHERg0,aC]>
_1:W=fYDE@IcV,\>=?K=>bA8_-Q=UfH9##OG6KQHL.@95d\Q)G0&f,S5?E8.R]f>
9+A)4\@VM>]C][c=I3VP<1>=<_?aP7GRE&H2#F4H:MP7YDHA4_?G5aWY2aED7,3B
84fV3Q6MPR[Yg&<45Y;_2<&79U7=+UKP)U@ccf0RYKS:26&9PSO<9cW2S14,1UTZ
_;L,,42SEbB3UUQ0R]X;R(+0[3>g.&AM=[(-EN/VCRNM6,OXO<VJ[d-a=>/2\R8W
gC040aCH)/QY_g9^\,Rg)@-/LSG075R.4XP].?X;g](?QbZc8f-D_R4&W3+X+0JR
3KXZU\f;1&Q4G7d1#U7C_S.@U81H_GdY:@PVcdRU6g<6fc]L#,J@),-g4/L8cKG&
]2If;UYQ_[0EY^gR+[&\DBAT1O64#J.gV#g+T7MV-QG6^d2Sg\1S.AI\>^/JPR/X
Z,1#08&,4)Adb3d>@_M(aR4\MV<bY,LK.;7A/[6<Z7_Z9<OZNf).TKCa-VGT.+PO
GN(GG0b6YZQS7TX-gP2D[T]M5NR0e-+<]8J0e9\>9f-DB9D+C-eMV]gH8+e&X7EJ
Z0^(3@ZG.9(E&Z2cZI2>DC(D@4J:\gf^7f490+Ug[;gJV4:PH[:0aa]=dF9@T-3+
Qb81B8)K>S4g&XN;MZg2d8+CEXbS?64\\.(7F;RdVZ9fbfc372((1P#JB_2#\4/7
dNKY6_,bFEe6F-ec9AVaV<H:(M/Ze]L4gAACg]JWJ4\RSRW>#cT>U6O_?&_]=fNI
&-cH9@GR0V[#7eHe0VS#1UEQZJYRRd\_6Y:S06U#UQK\[UfX&a3b6TE-N_BE)G9M
Z4NLagdL.]^>A8NHZ]:P1]LeVE-G)#=BI<=C_Cb2SBZLEK1HZPA+Z,cU(2aYO^<1
f8.)P_.I-(8:F4)QB.J5T]I[K:U0[CRU8O/QTG(Qb[36SP0\N>d]c5e#W:UCg(Q<
)^28XISO\YJYb3S+[Sd;-WL#+=6SN5Ag+TO(QZ3O\710KIVddACdc)GI(dV3MDS[
J/c)F#)RZ14<OY4;,@KVJ^_Z]_3NZW#ZYH_U.5?G9ea&MXAcaQ(T9/<ZRH8Q&W>-
^b4dZ]KS0(5S6YX40538EPSb3FWHb-Z:MI6(dWHL+^ZU++:-?B=TCfIfGND5-U/@
]N^<T+M;1P2)2]TD.M?0:LL7IeT.;b][C,[ANGH<3Lg8(+:4/a3Q1;aQ^/CGO]G1
6-RECB2S(=K8RN8?FgB8cIGC?LF(fW/^_-^CK=>[RQYAF8a9c6Rdc&BcaJ<W5A&L
IWA+e/7ODg;#3)+FXg:L28+MOE+Q&Y_.bPUN^_BJ03.?#/4S+gDGE7FY<ME3;-J5
^QT-9P<D&-dba_7I2[+\@#UBY>1?00RbGB.R-I@,KDR38RNC),9YY:[4P6gg.[?:
(.DS@bM>#N^?6XHQNZI1ZG)?;#E_>_Og]HZ24[96IVR##JPO1RgH^T[(N;/2<Y:8
+]T3COJ72>Q[#0B[c^@192/-;MO1HfAUZ.PU:]WT3PHIN@^8^5IZE/>O:Z?_>g]6
H\#,a6XQX4O8HV3WXQ4VBN0XL-e[N9aNU,Y9_P->?(5YY4Q3(R9g?RZUQJUg&eTF
\5,Hb/SCdWA^d#(F]MPWU&.GS;WUV<EPB+cIMP>+5RZXW<d\M6Y\Cf)U#2.M_>V?
DH:f=+8(fg1-_&X96R@\eG77:+G8-2e#_P^?H-;[V_957g,/OFC7GTBQ.,VP/?-:
XQV4(d:4\R>ZT#F47RUYLdg4e_1/Zf/^5S0^UP=K#E)Zb^#4@bZ01L=T)+eV\2PY
Pg8J]8277PeX;)\?+\7@X[?=;/@UfdS79>cN41#OP_TLYgZ_WT9.Ka&3R>0(VD>>
K]/V>=H?4#S.E,JOR<PK,7@cMVF79\aE0E3_O@,\/QWOeXR4G-]/^J-A6bW\Z&/V
6[8G?&a[UDf?a]76B,X_N5.20JLbg]d@82P82X\\17Jd?fMW9-K2I.SL1aX4.^KA
2S-Y+#EG@85[?63R97AZG^9Le;U=P:A[9=\UE>1c4)U6_M8/5S0?8_18&^@Zf5f#
=PR=R3OfNZ4K+D)fS7&,=@D\B)G/U]d.1Y@L6G\O:fJ5R_X(F-?N>@UNPXKCC6C5
@DR)ccE0#,/R;Y3;2I2cKB86SEL/.-(GdN(BTR<^3VHNTU19ec=B>H]Mg2>J2^T8
]>8aCZK-_,JBAeF(IUR(;J^#U<@@#-P(4G21Keaf_AVbO?5cIFOeF[&.Ob@B<U,\
_bZR^4Ke(O_c^A[c_dB+(/WaRVY\b.5;J(RN1;D>VFTFda]J-F@^1,@GBG@HH,We
_0T/VVPfMI]70L-Bd]X(fX(0,Md(2ZB&KQP)G6VG\eH8ID;J:<DP9H-cO\&83_W@
cH8.O)@OW)D-=ZU@ZSLF?(G:KSe63_SaU>cHU:[+S#:?Kf4=3=5<;E4[[(P^,4O/
C22N@Q5S?8Q7cc&\><5:cYEGZML(?B]>X)>C__14JD0cgb-Kb8)8KS)]c^+V->RZ
ETA\B:CE74f_0d.;ffTV7D)\;=K1c4]X0X,gM[(04PbFaKJ83f#Q+8Zf/]dd>QeN
A0CVM(:_+bd_E&G3FN^F#/OUB>1K#B^V9#NZ>QO]D(_7gVT/c2832dLVI.D7,CfD
9>7N:SdH6QYBHG3LDCN^=EW#0UQQG>5S<3>F&T<cVV]aMR^e>U?_YZ058gQ1eCTN
TN+701OZf<9)5f_72<)9ATWDbA.OQ^2f@#P3#32+N9/\R9,cfORN+DY6V4fL?[)d
JbNd7[5cJUeFEW?]aXP\0@[(ga68C7M1O5:_3^3D#gY1N7W=8NI+H&Q4XIYY>1H5
caFCA.)\<VQ1eKR;c3a]gB#2KRLVI<-4I1F<<S06YY(JT0__CXDSHfNKdR;(^;:)
2ULZGg8bgOE>cF336<^3MaB7A@\QQ(,aU(3D:93:L9N\.K(S=?T8M-J7eAL:7b73
K?7,\)I=:W\43)(;3H-d@bb:d/OG]g]SV&fEbY[MWQFKHZ31<T)gIM58UD0X?RFJ
YY33)0d.4V#5U8a(,XTGG1-UYK&;:\b\^Sf&aVMZTeB2^@X5O7g@1V.6<YWL,3H@
8FX[TN_F.+QT0MRgJ)S+V^=CXRI[8?/aB9/F::5-J)BHP(SG-9/#747HOa3/)gXF
MG)XQSMZMISDg/#XJS18B3CP#ZIVD1QX)+;eJ#(K8c5V[dB+VPT1D0dB)=P:@&=B
UKQ7VOH@dW\)+O.HZ\ETMZc)3X[PX5NVYIV:O^84IdV7gBEJ&D-TD@TL25a+BG0U
d-E8K0V1SCgT>RA5&VXRPV41bV.BSD-dYPN<^b7BJPWKCKa)b-_b];Y.f8Yd+5.L
FdU5@PLeSWV]TU3\964_B13]QB3]e)D=FQ2LS(9,L:D/<.6+05(b=1C6?HSgM6Hb
T<9^cJEN_2@67^;RDea?OIc6f]CC/(+SD\.:,0OS_Pa6Q#,HUP)[T->F=V2^?Q=[
4bTS]BcQKe983N(,V3V9Sb^d26?e?8JY1J^a>3VOd=@M+[&;bF.&>KTTEK5)1geT
SWd+/52J0ENPDWGSX:8O>)&Vg?Qf7,:B;dabd+?#H;?_?c=0QEL6MO=@aS,&TV<Q
^1(^7(8>CF:LO4]H=bDRGP=\=0g>2Y]MZ?\0YScN3Y+9U?P^JOFdZ5VUeXc8I&=)
(\F.K:M_WZ[f<6;dM;eEM=I9QO(_Bg7N07MfNGA:1W\FBcF.]Y([aO[eGggXJUCf
0[S.0(Cf-TE.?UcRNZf/.F+6]YQ<-JGR-0g92647(6Xg-K&=aVU]?NdM&.X#b)7N
Q++O[I9Zc4O6]Oa,I:Uf,>S[/W861;?8=AJ4e>WV\0W.N;(e0;_KJ\TP5I2@&gI8
2F0M0d3=E@;#KI@9G0IS+IVaU^PSbYQOVEbX4ROBK9P;TN8V,AIgR68R#a0ccPUS
QgY+d4[Y5^cQ#0f.#J?-#T/8Z@-3.9I9DT=.g&<?7&E)Tc/)-6a88fG;EgEYW@^F
<YTTAc:QQg59eF&AdB91OG8VL&<I88/+ME>[I-1C:cX^UOa:J;6?4GQN+16K+/O6
1R7V/0-bL#Xc#>V\W7G:N//=TcEb<+^b-;OEJCD),__(5)^(UUD]I(_,_X]N5/O9
B,H2_@f/D,HSSX1=^Y4UG1L[;ZW#(6WNGF69\2+Q=AE_&,,-A(VWA6e/OU#:RNHF
D-I4)@LM&8.ce+F,>W[FDB,GGT5Y=KPBdAZZCOQ2M)IF8LY/9S@^6<F)W9&5G&.]
I8f+2QCXBP/ZM,3(X.Gd6E?#bHQW\ac(<Q??>&,]4]6L2B1;.=1:/R,aNcPWUL63
I9<R+][^,_Z@?FJB\GCNAMCE6J5DV;/H-&d:)<VFb?D(b4Y?1dIFZW:FYDP2Hf+G
-Nd]FIQ:cBM5DVKU]=McB6g@O96Q]]//e1^^^N4D]QF9>.CGcA^&Z1Z,DB831])L
X4,GS?G\@9X,PS-R@=IZ7[>O,S==J\3d(VCA7YL?@0[aT#d2]7QbQPR[S1dZ/>YL
1Y3WUBa2S)EE-TeS)_)CM.Qe&g2]a0<7U3XP:^c+G&W3;CEI<KGBGZPSHSYKUb92
EAYP14HK-+NcT3HK(@[#3A;).O6_K\&0Z7T_OC^dOJW51)IN\^1b??N+S\2R#LS2
U3?R6Y\[QA>=UJZ+^4Q,A=TeaCJG&3S.F(#^R(b,#dc;LfJ[KFT1gV<,0@LD;,:7
Z.fN/3V]E8T/ZWI6]9gb7=7dCK+#Q=./OaAS(@gRa\\4^1(@+F,a+.<I#C>EZ<-N
:1#cP-&6:Q=>O6RPBdF6aMKA8?CX]S+AHS?41:@XGd51,^QS?gYb(M<Xc/:d;HVN
]\U1NPH1+&1DHZG/WNYH1[ZEdOV4=6;L.Z6-dHZ(^gU[7;L&@ORQ?bU(MCWG6a&I
3]FT_8+:GAW\CZ=#W-Be4D^);=&)<;XUIYJP4C#^A&&>3ebOQC/+@3eS,6?CDMY9
,33Je<@2F7S;#DH?DG?09W-@PGf50.H4)A[[DYPT>\7<#IDf\:?.^bP-D\3L--@=
fY>ST5S/Q-[PNef-A__18XRSDYY<Gf-@Y7_8dcCTCRKK?M@MG\LE-;@C6^)AY<=@
M&NFKRK\M>>#&4Zee#e>RI^#Y?7,I8D#.-FPN\=>=LA<6QG.W-_<&W7d[K5,:73,
G0O3P:?g5SRFIb]W<:OA52QbZ9JNIZL:GQYHE1e)(TS6HO@<7HKR]<(CKbe_bKNG
?PDZNXZIW^755,#K4&VM1+J)c5&G_T4N46#?>;=ZA8fgQV)[?N#S-Z))R^=+NB-+
^1fNX#QVFf<dE#06,AB/aXTf?AFf)WfbJ87V:_RLL7ZQDRTE2>#S5ZTYPWg.c2:@
.?4I;eb:@K9Z.57N482C#CZTQ4>Web]b5-+<E6;OF-OS^1_DP\B^-<)aKG@:G6_^
DRNS)E9)2D<L([G[&OGV/>XH02QH]5@&(ZV64/cF1+^GcVS6g+UKP/M.F+JUV^3/
0V]OG3^U9d5VPA9S(9JHOY9=,CfY+872C\HbI#)S^LW_-dbgFS#IGOZ<3RFQ1ESP
bS,VWgLQcRRF_VU,8b<;#&:Y7;)cU&22>C+I;IH>6:UVJ2N+.US[[K?R(:?FE7G8
?5(\bQ6>8[7M1I.JJ9_5[(=N9HJW/Ca_(C44YB&3gYDH_;3AgJE,,c>@PA,_7055
Db[J#_Mg&?U]V6+A5/.gVSOI7--aY38AHZfaW6a?PKOK<J#1=E7+[OcQ6.9LRB^2
8fP13c?W6@0U[aS0^B\0B3[]8ZNMX7JMS;(eKc/579B3DYPB)TNR\KP]5cFF.8M&
D)?PQDXG\@)&Dcf#CKM>aN1gX@\;[,5b5/1J)[?G#YH=_3;LA;5<f;/b_-FLE?9a
ZR]c[Uef\5cRJ&:01A5U71Qa/>-P.cd[ae(BJ3\,T1=^^&eV?f\>gO.M^7QdD#V=
(Pg(gHe<5aB^UCeR^W-?6O#PO&QgCJH.[EF.JZOUeV:&0Hac:<SA4?8D5M>XE^N=
)DBe3c13OTVUIS@Cc_7&Z(Q>?L9JeA]a-=Y_</?OJPC[DDAW8IIb<;fHZP2]&@=C
+.N8607E9H:5WfOS<=X#d;PIF9,#6gMS.2=S?CE_<1=^e;S)X[4fS]K75G(d&@9K
e=>e<S_>;;\4OQYV(XW5YUV0_MN_V\g0(cX0J)(8:UOM/[,I#0ZD0cZV39d?JM;B
LR4E\7JMN//W7DO/UbfIO?4J&,D_d3UP6#-,<#=IM3QgW/.DP:Y[3<VPZ(d?<16#
d9SH;0L^#Z1BB4<gF](daF^,3,:R25OUFEEW^UebG/V\;-[B-cbC2+H0:BUfXMFJ
VP17S4FX[Fb44S[?2(O92eUFG+7)S.MSe\&^+-&d#W4.9<NFJG3;QXfHKN#+=bI+
/,D@OY.289V?G)6NSR<McI.XR&:.]C5?E]W;a(_,WcR/WTRO?\^KDeGCDW=&c2+B
H+_[7O<-e[cKBBZU_BZJ,JaFT[Nd2UdF<+M.>YM([6M3HG;2&]2-<YTE@GF_NQ5b
PFN;R/U,K\>6BbLD[?D;O(1:=1IQJd9.EL:0,^.ZYVG2K[^e;c>=bV[VN/caQ.EM
_aY;\?6C<H6[H-V?K\^=2?_28;O1Zb24&=E(AJ>e?X3LN#;U_OfJGTdg9[bZ83+T
GEMWSO>FK3AIK+ZRY32RKAcD[?0A>f:X2cYT+OXc72_,fT66@\<GRV/ge:Ob7afQ
/VZ\^#8^0X))N=)4_e(5.+D[KC_;a9TJM_?gS?OCVB1OYQ->4BK/d=Y1BVeKGB#-
NN\?&@+OV9HXLSB]d>J>J(M>Iaf]A9MFE:G&?F7FHN8Z+;R_1CJDc(+SD>J1eF1)
[gMSfVQb7<^9L?5KA8T011XdaPIMDa/PR(Qd6?TTK+B;D=^@@XPea(\+=C)F;I7O
(9+4a;PQ#d(S^U^2T:8(WIS8JdWfWf9,IfPS.1G1c(5^;E=BU#\/P\9dLb5):#RD
6JW?#J<UHaK?0ZEg?fH5&5\V,BAUP;EI]+VPW:[FIZ_QZ\<<HEO[A<AHJ,#DU3gf
J9/d@\42^DE&GH\HH\2f4OP/FDaB(^GP.<<L1JcZQXW9OY]d=U73.K4e-Ta+0TK:
@(A2SHd?J^<LD+J1g+Q3M_FF)&2QUFGC/84-O0a?I(ac]c6bEJHFKJYQ8CR3dg_N
f\gA-0,L9PbWO6Y0.:4.@,5#Z=:Jf^P-7&Ob7]fa28.[G\eZR6A0c=,b/S3f_<b]
_:HZc7>L9)7Z:(gL13WCVG(dScMUC<GPE)a]V69C?C7.cgR4U4e0JW=fWf6HcREU
7aZH&H65>5R\QZ(^T9ZMXB?RQIUD26G[50?RQ.JE08YcRTMb^T@A73RUE^8VO#eN
gb;-FA,58-?O4#T\1-J0&71>f[7A1Z4CObLK_CgSQf-Z8d7a43Td>(>@-Jb?]aY5
/XY@G_8cg:PS70Y+(2-.PgCO5JA2]D.Ga(+NQ2_D7SDE-C25N=/PQT[NTegR85E\
->)-:5a<;-;[0K;VM)Tf8B4VF-M]+-C1V?<OJOE2EcDg-^Ba[O.JHL[(7G1F^_<M
>MFXK/7=723d7aUH)C4L_6>GTd2beVPAaD;Ib,\6Y#+3.T7SIG<CB(8E9+P6R<Ba
gaac6U2G=2\[-+f5_.K@PP)P-H[<LKb3/.:cOWMR:RdXIcO9K)+1F/M@J-Q8&a9U
f?JCH6cTLER<@SSY953;LDe6,aeNG9O0RE^9?@+S:GOB)=QYF9c9X<0<OU[JE6I?
[cH5>_f_bc^c3.VM#3A.IN7[ga_Q9BW]5eL@1@aU4?.=Od]K3d)[b=FGGCPB=BI:
]g5JPRXC7I3QE@2^+9+B91,cRJ&0V^YC#O[KQG2Q4[d(TF0,+H\A=R8HY6;X366\
eQ;fQFaT/VS7+EWAN5X:/_f.>KZV<,J0_c]F06#16.7aGF-1]DZTd&0]ACOHYRcX
RDQ0?1a9gMT\+dK4I4TNP5K>Ba^2<a)N9I9/^?\/V?AG-aF(6>F3KPH7)g>XN5P3
<;KG;AGS?S+1d4ZP[PPXD4E=1A97(7:FWPX;7T4bA\d,=ZURI#U8eE_P#dB4C,^)
g_DJb?-Y^[Ce15@&TT9I:DSM#W]BcW#3A2<R0MI9M(L_DV@,Z3D2]Y2N-^dV2e>V
,1@#W6AMXdN8E35T^\90&Z[cF2daDS)f-@BP;&(4Ge=0^1):c(X;BV8G0XH1fC5>
O0:.^/22:R9a2=X3<d/&X2V\V]DY.e8HH&-c>9C3RY9,IYTb.B,N.IZc:6BdaVFS
1#eLK,P,<2:YIS(+ObaS>&K(<1N545/U0U0],_:HJ#5/eZY/6M7ZaZF=UN).PLZS
g@O(.A<R67PM:Z]:cJ^?[S:J#1cN@:dgIfXfS3XD.ZAe=MUW&FY>5>ZIM\I,K#E4
Xg1S:I.L?(9BCa1b682dQ2]HZ.W8O?-3D(4@TP+3UW.AT=b9RG(UZR^QbV\/LBBA
Wd2c^RI.O:CB+96J?A&+.COgd<>L2fJAeG\<9,7?d1@&dZC<U70?L>)E8AOM\C,Q
/[a08E<576TG;<BD0;UG5XKHEQSReIeSUIG4M,;e)4=GE=2VWM&H),JC6&b6JH0A
b0Y/WT9RMB@/>XbF)a9>SDcA#XJ_Jg(A,M:D^)5X5AE-eMdW-H1.V@Z#I@I,:^HW
fF#AOK1e)=>MFYXQD;;.0;eATc72^#A3_QKg&g4e9ec,37<HY-C/\99=_,3_,VCc
=I1:8Q&X3(SH\:[b.Q7J&=V+A.5C^g.1Egb[04(\H6RXaJXY,@d@7VVe/C?0:P1b
.D6JdNS4(D2PL.@4#]8c><_,2+<#5gVNEUT?aIY\F&5A?Oa4X;^2bM#d1]f2Q6:H
A]b[(=f9=D;d>T#?JN>8^1#F+9-PKF1NGV7d/[Ed@#DeKCU<#TR80P.GL-I,5D2d
8.7@?:dQ(GAML.O8AE@[cD=&][/&H#/A&;GA^;E,?89R+QPdfIZODVN-8Y+(:R;\
4_UKb3\,O)RABVXGJY?-O&;[OG/XP5SN(ZB,MA[9=QG[N[54TJK3=e)Z;TF&^4A&
X[fcT<@]3WQP(7+&/^#.NA61/-,;c/f[63T>\EA8ZLMHV6W8LW+OWKUDXa3Q06]>
^]@LBV4cUdf?QG_VV+1I;?L(e,X2TY^D.(.;4<#3&L5,N70[/NN2c.&B6\(29B?D
79b8W96aRUHd)[G^S(TJQV1?FP6HP0<.RAUMWWD/)\1Ng2L7c8V8#HDd<R(<CG;b
[Ra?SU^M7?C9IJUF:HS>1[/HK;eYDL;I?F7Ba:#c/H+2O.LUfCCA_?LZP)b;g[7=
ZW17JL],UgF:AF[FI\e\1a/WS6+#U-;FN&b88P@FN).L+J0QXTF3XW;^AX0?/]G7
C9)6MH^YW6bfTWLVSQJd-&AU(^P682^@<WHPB;S80YN;E0If1aR7CE2O-X(b-#@]
cFOAJBRGL=CC0+)W83(Q<S:#Y/J]P;Z5>UHU1?dJ/XB_IE::Fa7LH0Uab)H=E>[5
W8)@6:YH=#4/c9cIJ4=<KV,g/7Z8I[>c@QH:HS6OU,AH[@HQSaO><A=Qb0LL4/Dc
>3X#c<6c3>QSfXS2]Ye0AD;f603?0D2J0JE4Z)K@V1@C]-)Y6eA.JGIJN[1L+\4V
]bC//F8P19LK0gPZbBLTU<N8)JOQQ;Y?E<WI^Ue1_I\R,0H1-C:X/9dK:N=KBg8Z
5H-1aC\Gd=/YWdGLHG1OG5BGMXFWdL1Sa-Qf>L\-2b)M<.>V&1RG/F+]/]8BCNO9
B@\.D\gf7DLZ]T\;(X33P<ITe33\bPIJ649eOH2>TL@L:<M@@-T:bCN=)9b.2MWA
KH5IQ=_[/_MXCVUTJ,3eNRBR@,@]aACJ=Fa2CHM<UQG;[a@W#AD5f]@][>4#N)V<
RM(EI56MDEBM36T@41IST3WYX+1MO:=2@AXMb+5TfQ3\&^,1d_=JFS;88Nf67(;:
?<[73FP@bS7D+aT1ER,T+1Y=FC?OK.eg<f#7Xc+&;[EZMfGO+,9A]TX-_?)C0e,d
O5LaB7@RNZ]gHSH/(_N@K1L?cF/J2G65Z@DDVG^-@Rf8Xf-&,L<f./(V/#U)K8:[
2Dcc<Y[IW<EHS5.cK#;CJeGd>]MC/S1;bFaACcd[CF_67#J:?Z]?Q6cfcWWFbaC8
&c/<UH2VQbRH+1;1b)]BEHW@9(.)g[HS;T/,0:BP8-X)YOFL;#Yd_(HXecR7WaU_
;V\fTPH\@[LZEZS,Y3H44EG&0ABSD^KeI;86L.CBe/1GK/?W4Yg;.:aLIVA1Zf\^
PZWFQI?F;4?bRaB]Y/;E]YO6aPT;d]T#M#Hb+d:gfP4)e9b4L_JgFc,95fX(Za#P
?55-/MLE0>:-2>5CcNbB4QY<8F7^2L1=,a=G]5Ded,54ST7]:gZ[11D0J8f<Z)&B
.O:(-&Y1FgH-<OP9>^6XSaEL5-DaKP-DQ(?+912A,EfJb]6d2=W7=M^32FPd5\BX
N3I@T/L4V9#1]C+Z\KTZ0,Q/]ZJFG8Y0?/]&eGFG0J);Q9cdJQ_?J5],gNCG.D.a
QEDNB-f/=Y2X@UH2,aD2f<e,MXR=5DX@3=g?\Wc#VVEO=4AO:1CK\gWd9G[@?gg+
LK6(GA\I##K<R;gV[e6H\4.B553+3XE]ec+#2D3:(?8O=>?Y^9#-/H(Q,X#,&TXQ
Q#P)A^HD,G=39,D9QgTUD;&9OI36:HWgUQR.(&1?:;0eD/a)R4HMN=4T3).,#Se\
D/YgL0.CAe,/=LB(70=KTOCZF=BC@X(#HgT]@2Q#I#5I)@-QVC0>V&f59B&b\A&?
G^7fJ,K\B\ARFT(cYRB^V/^:#7U@:31M:Fa)H/KX1;[F8YX=Q.&VUZd?0I4QZ19S
Y<P5KOacg.#/N)YABNA&E6]dV>A^2,[BM=K:9N;NASHLIWZABa-D2I(;2#.H4f&F
?W9(+I5aIR8GR[(?^5[L1?BfDNA8K?P0<9=DB9\2.YcJEDIC^WEQaK/QG0UMgP>c
.2aJZ8F_]3CfUDYWE4ce0UQN0.#O??.5Oe,A659SHO?UZB<O6)H:@(F\B(:UU7J]
1N\@@7b]^QF>8EU2;\g_Kca>[?LX;:)]3QU;F6S5)+5XC:N?3^bFQ6HNeY(ac5O?
Xg863e2HR>KW8W22YWOH)cRL;g;QI7T&,VgDD1D?PNf_I:fe[T#5AV>U?2MU[&[[
VVA,#/Dg6U6X\K\>HeNB=GfA#(1/>aeD;)1>X,TaH<]gJHY.0.e;FOWQ&^c&\1CT
]NP7@NUXD=;Y1Mcf40)?[6JF0/WdcZcFJEfDB634@2Z\&)RY(UCR??6e:XXRWSF\
eP9c+N9DU<A9=-E:A)4888g(I6G,&c\VHPbOG;#J]W>a3^g+(J9[E:D#=E,H99b[
RD>B@KeY:1@VK]0AUO4Y-(25XC#;/]+JK=gLgg5U3J+(S357Wg?-d/W4HN7VaaE:
=,MWXZBT>&&O]RFV8a.#L?d;JS2a5\b\IGH.7TMK-?&0U.IORB&_:@21BWZIEA(.
6R[CN=.NHWLMffH(V5>IcI]BW7cKb4Uga.fFG,V_b2cUMbNQWZ/(^<(2Ib47\a^^
b;G;V?8NeDM-D:S7f4PF>,d/5:4T5&LCDb?A>/EUX3QKG/I@YXL86+H?FJPfN_<#
CT_K,^6VQZVQ,c>5eZ>e+=IBY<363J?I^eS(W^18<YdJM;D..U^RLBY5+;@_WYS2
ZZ\15J2&0.SK_?(gfeH?>G;g#[YDA0A-OME:gM;JPS>P8J8aJY>e,L]-67QQYe6K
]M&<gDa<S(L^7M\C8^>#>@?G82>1+fHXB&6cSdPX<FAX;9_I2XSUObVbg+:Af4U4
X:=B1E;Z^FP79,?\E(gHWR+6WWf0eT_Wb7K[_C9e6A7FVL.^,Q@,+3VfHHg4f&;_
T+,Qf2H59@@.@VI&b&1<N/P(?5XTAcTCDY9VeLYOAA\T0(eP7H^1-=T3Zc7D_0bB
I\/cJ+QQ+_&7H+H#PCdP\V7cI&I8&@b,.C:V&U#eZ6+C)2C8NaB=^;PRJf0SRW\8
[G(B7,7P2ZTRJb\]K,C6Gg7S<-1_g)3LD[6[/]:?^7AINGP\.XZ#4^&RdHSg8gcT
f(/]0(?X9Pd0aRO:UF?::[FdL&[?g27f3dZF#(fL7Z[@R?BZ5MMQc3=]7Gb+M?.V
,K#aNeQ]b7RB-7AeDZCYA?QB8dPdRPBb0f3][?XE6VZA<5UZO-<H.K^\>DXbORU&
.;>IZZg,[0cN;BGYN>1Xe>0E1bFYd&A-&MaUgE;K.g3+KWV:4.EWTHbF#VZ@fHa-
LdI>^04LNQbXdHGFBW.JfSd9efSeMc,FO\;(ISLOI0BFfL\6?FUL7KHc.#G+CTE5
+DADeaRDL#QC.g.)3\H6TPS>,0)-IgD/5\L)DYL4@UDeA+KeSA5&K]^HA34DGZ1W
^&cMKWJ_8E(QMb+Q29W17QDC-S3GAOPCeIP;C17FM/5T8Labg-cO(A39gGPPQ0Le
Og<X72,NWIQ^,+8XT8S\5^PgTg]XU@M5Ng0g+IA4db871R>cE_::V[NQ8<#Jf_-_
Wf1.DaI,2;Ta[\.RE>N;C.D4/\<K2^9I\=61&67\-8/>#[G3(>;.VZ->]?OeU^#T
S);F2IV(-Ze:5N<IKMIg1Ua[?fYU)T\Le\YKeYN.0,/FASV&&?eNM;W#;IS9U)5J
Gd[=Lb0Z),RAU/3]NAEUXBFF^6_.REXI-Abde[cbW[EZ[bQ>+eMOS<2+H>]1=&28
=4PDO/-;DN@F(7773QE7GP8?6JV[YB6CTC&),MON=B[MQ/1e01X&JRC+(_c8TLBL
FHKY6?4/X:Kc@\W^f^<aY,Y2YQGFKdOe]=G9I>1(V5L@dc8^8T-#YK(eVA5@;V19
9EUXW0R/]+M2(HV#[-5PMf[Gg6NY><2I]@ZW;TRIZ3ZI7M6:;UP>NeRdZ+cOb11A
3Q?0bSP@5+&B]J2f0V;#T580@f/7=00V^-4?\5/O&]G4(I6>.@52<XK)L_)PPNZL
P6Jg2VgC=1<&AN.XTa-(#USBG8-RIOZ]91.A1CbSI^9+c8+.9?2c97#=?agRZXgF
I2:F\X)-aFaJ76__N#:@Vd0[Ec8e3C+B05H\Oe.0.U@DH5,R4(4XNe5cQWVS+T9]
F86KLN-,E).2.E^a7;MfQO2J)CeU,#)MI,K4/[1;2e4bA&G;>&;YPf+LLX^II:;L
UC)MXFaC(b]<e8KNSODff,K0Z2.W9&R\NC/WCBBT,V+EGY8MdOd>ba9Ua.CYDE7Y
:73Q;F?M_Yd5\@K+Je3>PP=6[OFT/1WK:X8A=3@+TYB1N:7)J&5G(FRe=eAJ-.FO
Z]HUQ#XOHV:_I^WX:&-ZW6EOO[cW?-]e^N:Z@7P5b;Gbe14a:.Y[34?VXWT).34<
[;>9XLDf,\XEF<CN\8>Q>7MXdUH3P:<>EPXMPPc)CUUa?DY)7bSaGOW;_O_D=[,S
MbVb=([PI/a,#JOX]4fU:J+LQLI49TP04gGWBF&K19IJ7,)C?V/==;72.5811RAI
B/I^<[W;P/6YVDEgYINO^G^E6>OQe30:<_MGST8@+&\E/W<LZSdI1Q/b]eQ3?03V
^/_=]Dc_^<YI>O=aC(L2:^X)a9fB8P.YX9&KE8N>JJgTd5EW:U3[bb=2Df:8M:-&
eCD?2??S3M>3J6.M>JC]\=-_^bESg?d5\4JaDY<gO;f?eC+Q(8WLYBXe2U/I)=F3
&PD1RU)_b2/e/Ue3^BdA7af0=]VP^SA(BSKXAAV)57gKVF71#ER3::]=LXHG<PdP
FYX6V1ULB2,6H8S;DB3PA;:_A.=]g78WeGZRdK:b6XVP1DUJKKX?(T,\,]@)XF<5
6I?NR1H#)U)D3RJg0=@FO9HG-6Rd>bKb8BO,+HU0T?TTWdF&DESKJI55V=Xc&<4(
\C9>8N[<^^.>RY(@g=PWZUC[T)>YZS<(cb-3>=APAed+a1db;M/])WIdd1#2d0JH
2fO0_9Ac/=b#L#+)M[,9J@B]<.5KO-;K[Jd=<8b#\ES^HAWGe5PB\>::R_J>+14Y
U4V,M-3DaKM+TMg&CW2b+/+@@-Q=B-#[3Z(YeC)^;,Ae@f#9M(##9aB/AABY^SX)
@AWd5G#=Ec._[c&:[A<B[7QHTGY:T)<V@LS[#>\XHZQ5cDf9R)B<fR1GCb#c<PGI
948<B_HA7P_75M9aFJU&9cLZVfZaaa@AXSSYC+FVWV&PbMWOV_:ZJDK6+fgCG+X9
7b<OW=?J)+@@=O56A+/@K#d]YY6M7c-V9bcN#8RQ)T:>cB)_.=.7_E7@bJ(##?F-
gPQ_7bU4,@KgM]5UFg,3WFdN,T8N[2.4BL67)5&(-D#ad=S<WR3VJ(6FZR<-]Y/9
X:>91Y^GID;[@0HPfDPf7fVfIE#e6K]BV\d[F:J12d;3a3G<PYOg,Y7/]MERM^6Z
21R<DZTA23(]3JR//:X?02GOR3M&c7Jf/+U#M>?GbBXM/]0dSU9G.=T+-KX8HE1Z
TU2#C#f\&;L\Y#3G14_G>>/85;VfW@fGbAPIYE..1G.N2+d^Q978df6TeSP3PL+b
YHARLCAYcB\GbBIVQ:B]Y4RD/^K<aFW]Ag=&Q)1X&X0A,=fC1<Dg=PFTMV7->e\3
/N3R7\9H7b21V80-(I9LTG=ca7?3./G\8ZV7Y#^LT-]<M)-)Q<9UJQ9SDG^D8M\\
0EZ9;)O?S1I_H/T8-=W?]=@d@7WD:fV/T)<X1_2)e3&LN+Db]fD5f[eOGH--5@;[
0,QRIfV6T@]#Eg7H-K^B904cO-ec?9U4FcdCR7-c\;5MWG366(Wg\(170)0JbU1)
9H5:2IaN8F.;B2TW4Z_A]GZXV?gNg,0&:2J05:,b2Aa:HbXGVTM:0/_dY<VT@8;8
e>b8gE=5X-R?Z)T:2SR\A6P^aWAb59L)Rg_B-KO81>C378)TV]/@O,JM&)Z>RUD<
9T^)TgYg6C2L\]I2V+cD[>OG<@Z#L)2\-I94eE[dF+46/VQB3BAXPg[;f8IP;J<M
QIXINUYK5-QVPe9.^@@(0I4U#H03FI49RN\_c+6?>fce(a9=\J/KYCO1>VRbYGZ;
R105QcS2U.C+7aCdKO)X]^Q&dGRG(#H=2A?&PJ?b9\85&2J>=;,UXB>]/X-f83gf
5bQZ\GePa2T?Q]73c1@ag,;0W9.=.)g4)DR)[gg[56e9CT&VX<V@KA7\#+NJQ@B(
GSPSIJM\c=D8?aXLC#P0:-]VV<(c7I&_IH1\X1D#T=6ZQ3SQ1_+B4a:8cX00C/Fa
PbM)\XGea1]_Y_\T-(&9VIbQZaY.;K2<&K(B1Z=?\SPF0@APK?dVUO54Ub(T/.PH
CY/4=VKJ-E^Q#a_)+9OGeG#3dQ._NH-5ef?La](O4AZBKR8d6I.VH(RHEWfI_;AY
-Y<32?9V^,CB])MRP,X=CZ;/0VBFPe8S-&5aD:GZJ>I)e6L=43Y._C.YfZF\J_:R
5@2H;9V0W&ZQ68AaP/T<NbSB_VE61K;R97A#b_e;_WOLEd@KXEK;NQ0ceYBL@0d(
4B3<1KT?[?BK@2Y2+f]:W12[&4Q+J7GN_I6Lfa\GVE/V-Ob73124Oa2P6WK[dX1F
Y[4V#Y^@/K6\4H0e[4+3N<K,,P;A.:]dK)91A(+@CVKWF1d4-a-3/[GC3O>0[3#8
A-=-=#JJL^_0dgg(f[FY(B(cRQH>C>6cB=I>[\S1X2##ODI>2^P7H#8-fge[(bd7
_&_U-OVF_1aB8V=>Y8GUF4e3W#a5cTgPC49\O:E\e=aJZSJZ@bKK_8)PD9+-UTgN
^;\+2Pa?9446)((:06S6cL3e-ZXgZ6X=O<Ggd5gTR7UVUCU3c9LaAYNU/3NWY0.4
Ed+:Q<OD66Q9RB=;^bUGYNQM@(@:<WV>FG#,&EX:14B]^4BN,=D@&IdQf:C1G5GN
2Nb0V6W&dR9I#JUF93,_0gGT(NZ.4;LTO<1=OVAB,Z^R,_f>[^^PE0;02cbR:PAa
>XED12BMX_68&Z+gFYb2.5+XS,<W;Ib5@Q26V&&:.9cP6(.VKG8;M7f>FPRBM19b
.-f\W(QI17)gE#>@E>Oe:=Df>bA_;d:UHU_eU92fN?]JG1;>[(gPa)9>bD:^@=>G
Y7HMb9AIVA+?:J>aJLAXX[d2Qg#[VPZDSaIc<c8ZfQ\UR,B6FOgE<T3-.1(QQbO7
:]De5SX?8)D_FXa2IL0=(+&F#cSaUH9N6Z]Z7,-&G;UWXYfFFb/:b#0fd_GS4W,#
b],@d(#C/P5F^0B9,.IP,GbdWW6RL4\))E]K=5+.Ga-3=X#S[\NAPM(/HMW6HY=A
N,e<M6?YLa;H,0YBeX^_Q=-/._I@0\&\T?aE9&3U[&1c72LA4gNb@d0\J,+>IJbT
f3IK=0&#I[5&T#+Q&HR,,C^RM<9@55fFRYT]1dAZ[P)?df:SGd-76XAFH2M#7AEb
V57-1L?eEX2(6c6KG_bJNG7R]0I8>TPJ72MXW,eF9\QOeL)87VW7]?PEKX?Z5HUg
YgBKJ<dPJ26b4>d+69OW9>cA200^\_IS/J;G1RLGYTP+J.ZCgUd>TFCP-V@f6BVd
((GdGP7>G5a#(<e?RR#9>>G)](ZLIV(3=Z@S15c_;.;KQeCFD29Z,dMEEP+S)991
,R0bgOT-[Ydfdc4Q]IS[Z&E8\CLP^DAK@-]Qf,UYIZP<:_<Dg^TETK?;_:^_Rb-\
#IV5c^3gf[T0B28]=P98/fU6Z4K+b.>NCHG.]Y<E/)fd5gS;0]O.DN&]fV1@9BHR
QR2IQbD]QKQ2eMBGDTQYYNe&:B?Ig]gg4H)T\&RO=TT^EHDP(T#Se,UHaJ;[H\=,
4gJAMV&6A,N#I58R6YgdKQe^4Ha_,#WY>6DV1EVaD/T7f5FY6XSXK=I@\;5SFfe#
?_O[GFYC9J:Jg:&)392XJR>MLF<U/IaDM<dED9X1eW)[+fbG,g>Y-QdgT=YgYa;X
T/5U[BJ\X8ZeOHNU@SYc],M\J-WC^&_g9000eMCN&8N&<J,\ALgC706@^^8/D=F7
&1)I-T058Q6,<QYXMOGB3W/=-U-RU\=_1B0HcKYEYHW(8&UG\#.F+bN^Q4Y@M6?D
9()^;3:6CMc]3b2+>=[Q9YcFO3Geb[7<a.5&MSJO.WJA0Z\QgMX2HD7&OcO]JC:8
G1Da0g1>R;.J4Lg.VWK?.ATK(UcAO4#-J3[MDJFV<NEDVO(CUce?\40VCG0T??3R
SB^H;LcCSUBWYL9fP&7O[];8IaN)?-]gI]7bB2aA>(Y/S5H04TB[HOeM==CLR+?Q
H:PE9fMM4&?b4]b:HCI+YHB:UXFacS0fKY\XLL8O8b@;N)K9a/R_5R5Q@M,Q_A_-
dIb]eRFD?]1GeeWPV[g+FS\2D+Vd<AObU1e6Yac_MW-L]E6+C&:cU<E1@BRDe_35
TDVE-+(QaRVE7-0Jg7M23MF+5(_75>a,4?:KD&aU]C8724.CL]H5B-(/+Mae_C^1
9ReEWf;C.OEG\4MH5I2&@/eC-V_-\559+HX[5LaT=]2N?2R^(ZC?1PVBU](U?J;&
)ZRaMD1?-e>&07YcfK-9\JIfX==,-8_SP;5OD;UD]XX.KQN(,9L=-aRN9EKJ3J:_
NCb4.1PCEW4]Y#,^S:8D&H&Z4[G.]fD=\ST65+OS^>aJ5G,(6/Q<Q@K7;0IG;-&\
<]D0<Fcg+>:SRQ;gD<7X.9OS?,-I?L3>H4Ib<+,ZO#-#++T(QG(25a1HCWHV+F@R
W[A9.bKVL#e>(0L[>NZ)\Q/F=,ED9@(/->FLR_fc]2+454(.E3FU[fR-8C5/F&LJ
UDGC6G+E_D@]VTTU8A:X7^ZX6.0/3eNU^=&)^E,IFM2fF\.(IaUabc<?##RB[L5E
B-5Uf?SHIWT\C-AaL>\CST9CU25+f_K\=T-C&2C(7TWS/SI+d]DP:aIPfR7MU,DX
@::1ZNG^;F-)I<]1()AM@VaA>5H#<[6;+F,c^.EI(KcTZSZdX](H9cd1-c0=+6,J
6P;8?Q=&)ZP^A?.U+111)K.g5QCNWOEA2-Y#F]AG4<;L6VVd2&;&gFa[195]>6U>
^Jg[&eDI->@(1B;5g9WcKD?>?Y\GXPIO??T\P<#T=XG16(83M5.Hd6+W&K8X3d9=
0>=0#SS&DZ=;8AH#52-[X:68aLVORLEQ#VKMH3,:60YN?IVLRG0@fKaDV84RIOHb
)\TA/EbUG&8.OU:g9#,BaO8O<H[.]I+KED1<(F6RL8LK2RCaJ))1[VQP3T<2V\;a
5>5QbgCJNVHF<4A0W7>Q??6QFdH-@HW=BO<,@Va)-O@;E-[+G#LU7V?KaF,H=0)V
f/)GWOR,.E#)AJ)SI#DG\^f4V7R,SVG7f/.DAW@E)H3fN=M=gge,\TTH4LV2E(L,
=MMGLc1>L6G)\[.>eI70Pa;X/3?Fg4VY;KW,PHXfYAH&NUSVe8./cPXISfc8da&+
4eY)MK,)#/JD4TXI;UAJ_I-C>cCQMH+Y3M((e@2dDG7WB;J;b-87XdLS^d)<eDe9
ZDW6DP#aG5K5b8,EV[(G68WRT+g_]d2#gOZ05A\/24P4H5H1Y3S\?Q\N:CR/L+Bd
1X)OXa&:YZD7\cU)FAXDbRcPM>cN2:eZ0@T38?7NM771DWec,NRO<:]Q/9aUX&?\
(Y^b(XGR7E_F6-Kgf1V]1-cQURU;dB4_D)44R)Z4ac(X]0KLP6@b[gPNb>@eJ(D4
@a_6?X)-@5<;.D_PL?#2WaO:fNZeRG?,E?Pg0PT7MYRK#.<.E-F_9U1A,AGY(3/?
-0WaWJUgU#ABNT8V,_<e.GZV]IDdU_5eE^.e60+9>Z?52YGJD9/=R1f<f(=D8:#<
+^\7+^DQP>fLGOGJ6)Y2AH3_&W2[B\9OQg0:,<<\Cb4b1RbZTJ8P-De#OFA+AD<-
BX6:JM>4fV]#-K/YL4J:ZbV/O9.,#+ZUZF7_e#_<VTMBWAFOa<1a)2e<AO<IUe^)
(g(b.dXTSK5&8]fKL2-I542/(HG>#Rg2GZ=Cea/5<&54G=F@=E.]<\=9J+0D#-K\
MeC:H_E.\;0Y4J,<3Kg4&Ea5Z(Bg6-T4PVUgO,)0]&\^V=(L]TKL;QYK0TU>dK-2
EAMVQ:<E[>ROF_^0QKRJSKGJ__=cc;^9^RGF+]\?U)IBVAI,WcWf]I;I^2]6/b3_
G0M#@;1KQM6+TYGe->K/Qe8e6W@d>E/ID+NM+W9#(<\P_SM8FOG/PfO-cg39FY>c
beTQ+Z>30L&4Bf_TZYRZ9MJ:0.&,BDCS;X9B+FAT4E#DKEG/,BN^CDg_)<+I?YIZ
M/M9US0gP)4Z,O:C(YOXIbBUU0K@7=Rd-<M4JLFGb0RDR@L-X4.AL0:AREF//._8
RadTd.YTDcE\XM6dg[&>REN3d6JXBW[_,R7a].UG6UeC_(?X;YBJ@/Dd_6&:PC_L
@A492)9(b]PR/A37AM44EL3QeKP,R28g-[5S=U)N)G?#.0[fg#E@W+)JCSW-AE6/
f^IGULOWKeI\=M@FXPdWWV?G<,Me4H\=?XTY.GW^083S5)H_1L7f;JLO(UU<NRR0
a3?_,(EK4AcGC4@J8JZ)Ec/Q./HdVB6T74Cc;e-2U7,-N?R&0;]^\SPH6PRa/eg_
g6eed4>7C9>9fJb\/H#>[F(AJ8Lf./85b<SMD2+W/;?BWP<WJN@E9OL7f,H9SgeK
^NWIE[caU]XX&:8YRGd+IQ\MaFAAe6E<Vfb/?aQ&C103LM1TP<FV@T>P3SW93AdF
bdcfdX>\0S2TbS:YHYW2GeW2f-(CLfBC4]5>.OOHUE[aD-[N@H-2OBb2&U-(7+2N
&B:ZXV6[Z&#O&XX0_QWU\Q4M)VD^RPY[]5L>GE=;;#]R9HJSB&>^f:@[237S[9AH
3a:0SI1+:I72dTG;]<@/]Y?1SU5\=a;2F55@g1WO+O^CM06?\.2Y[b1^^Zb0+H@^
F=:2:YAOf.bKf@F\0+Sd(NOHN>G8X=OPTZTQe@1f/,\U@=3)8FL(VX))7ee,D\9[
=FFA<RL(T@;K\;@,gT=@3AB27XGf+W2L5^DcPU2-^2I1/VX4D&b]R[MI9fFXS(&]
-dRE.F#3797D1U]c]EK?YX9NPG_+:S2&NQ2]J8]f-RG8FC\+CPgQ&:R,N\0;>507
RQNR@GQTB>A9+./Q>.N3-HdJ0_2LPRf>f43?^9;TaV^-eHUJ&GOS:3KQS,_S/<?X
\F42)Ua/gQL#@LIJ>B^R.;cUXUdO9E=&PgDNU\_Ya)KAaLB)-\H4[>3DEM33XE-Z
[^.Dg4[d<<<,XOI9_d7a.:25;589^Pd&U_365LKY(P+)2-XQQ55adAHM?f.d>B/\
3\GZgZ5RI+XegeWSH:=AT>b1YQP<.PG.D914f6RH4CMEbT7D(T+HeG+\E2R=Y(:[
&d-cGC@;7^@BJ2bJ)<B#6R1D_>;HRT&L:+N05(B009F,RV/@a#XYdcYAGa=L-_Z6
d[6#[/DL([J:VT5OWGGa1PITZQ3d]F7&,S)WP5=;)&0TURIWS\BBSbe3:7GLNaJB
aH5(Y/6WdAgIV(Bd[>Zd=7\:Q7>fKVSb;CKR&&:<6>H\T=bX-2LdULXJZc#/dTO?
CD#3[[5Z]<O(6gc^Pa/[d,[[OaMZRZ+,C-dOKP#@I6e7V3K?YSCN))A&O&H=/5<d
/2JTe\I<+b5.-/Ue74I5g<@2VLDUJ1cV-Va,3N>K-CI7];RC\/5,YP);VJPd0#\#
4M5U_\2CWGGg,_Y@@6]QN(a\O1Q58ADT7@^+R6ZYfV\\&B4DJ5916P3(EdDK+6b8
7O]60MN;4Q__]B)GAGFA3]ZXZF(YcK;a:&_6:G_#W_LG1D2E,3;M_L2e-9?5Ng@[
ecB_?g#L?9=9T2QCR+ZSZUf/4CT/<#&8:;7&SAQ#-fUb/?aW:-.VH#IV0,(N#fcR
.9eWEXVF<bZ\&Ud<X#1f5-1=8gV>bQ[=dX3T7=LRVVV0)0NQIbOaIaTK5<JXS-82
d2T5\-AXd65/AVd4&Gd/1.KDc;_IG:-L#VPFSa3K3:1>SJUL8OJU48S8&#b]Be\?
6)QAcYWCEdR[IM[3JVWS<b4T4\.?5Hc@,?-/D:?6Q&FP79<?4fWe;d<[Db->aa+O
?VUZM3eVVY+_]ECSP_/W1(JCd5OA_+cOC-.f2eNY<ac&T)BB10Nc\g5L#YfGK&&C
,9FIXd32)g^&+efS1b)<I9CBZASDL_HL[J38RaaPGGSa>YbTLeE0,F+b3Ie,_I10
;1BSYMI_g8FQb[7O_/\MZdcC5d<ZRW,08BXaIA4a5ON8#7I),<A>W]3=J5=0(e(=
1g+UZZ[EK&ga075/]R1,^,>E;0-1H<E4];I25C=V_BUYM=_IeZg4LG[SbB+6PY33
d1HA<2QXUS5fZd&GVXaa\+0B]@8^]2=?M.E1Q,^V5D^JJW=YORfdC3#Ic<L(E47V
G+.72Ufc2eb2K\Vdd]]NRM=#]FL615@Wa&Ad9<I@Q)>OFIO.MdZeWG(bD^5Y\J7@
M:-VV.(8cLF)3:-TMF0KVXAN4c8Jf_4dXBfWg,CEDVUOEHbB?\4N,:[5e#0A=0Ra
G2Ce^+,Sa-/^1M0G,^HbGfcc/D;cG>.-BbRG@;V.96QTIE+8F3]G/(1YU(J:LJQB
:e2KfE;CXbOC]a#d+?Q&3&_Y9]?G.3aIJ?e9)c@2]QF&=_#-/O-JB(f)cAP+FH--
T:BZO0W,(N9=,@?<N_)D@gf57OQRDD>b;V([O;a,1&V40RJ7Gd67H?Sd/XN.>R57
=2EOE&TIB=C2?&>=ZD2^H.+?A9D+MH>AUESP]Cf?98XdO0?U>FcFaOK,L@IHH(4]
?7Yb8XX-?RYJPVF9bI;&a-G5LIPG7TY/=HPF#Lb4[JNXU_IX7bO;?E^1>H16,=@X
f?_Q63a^NBAK[G)H83)bKT\]d&)2<#]JL5SI;R#RXbP;Y55(=8<N_#<>C,[8.O<0
QO5,@;NRd@_QL3)?I6.e-5+TW[_5QP#)]Pa,d2OR/7[M#S_:?d;g\QQeK8F,.&cQ
;]/&BM@SWD&R.CL86&gcOWZ2EAg-QZAI0?XL0Y\NcQGE\ARLZQRf,.UNHaa&H4CM
B#,#g@7&@[ULGaDNTS5c^+M[,Ia)?J<W;7\B4e+G5BP15Y(#XED31F7]UQZL^8P4
38QLVc2+UKLH?N?(QdQ005><4a]43C53GW4.eUN9XJfRg^#534=RQScJ/9DK2gA\
V<aaJK+3Hg79<4.Y3.aaP0;C&:aSS.IKT#+&/B<#K_2+WHfPeJR6AF<c/aI;W&(K
9AJ]9)19<]M+cVD.7UeZOF(FTGcT,bW>f?1L@8#8BC_SF<86>TM=4UM<&<[,]7F#
5d9H;Y+O-SfWV89\U9]LT(I[6YQC6OESBA7<3E\]X>4+BMY16WM@(L0_MX;)[T77
/d>+T\5Z/T@H;FKHM=eHf5XXXf.Se^RWO?FIS^MgDR@a9;R:ANb0-#EP3-^KGX&5
+2\T3R.1RM;.@<L9cO7CbS&0YU6,d6(9A,9Y.@,#&1/0_0+dKR6S<MJ5C:];fT:(
^GQef<M^bbV9KO\PH4A,U:U8\B>/-XEM9gIO_0/_+YC5#L4RZ+K9E#R(([@VX?2J
BX&_17K/1S-^T_&:?a-0^ge94R-;<4K<I#_<Qda<29EMS.>Yb9MFETKCDA_Tb+<N
6e8YI7<ALf4@-^RaN28_&>MZK]JebBSSV8XM[4MaHB53=23#6W2@=BeCTI3=f&K]
aU,f+OP5J6I5Q7eW=5FSL96<AC3JPd;K^M]J\N2JE29-@aR6H27]1BIO=ReNfH7&
-#Z5FCXMC4Q/>bJa<>G3U.c=C?+TCV(>^XFgb)T9A13;DJ>e0bP:a=:I6=R=CN.a
7K9M:b=GPT1B7_5OQ4BCTgU:Ac9I5@#^I#cM=e7eY)8IZ2@P1cD9D(7MVZ2L2g1g
c;&+3E3>A+g70Q<>VdRF-Ua7Z2URZJ37T27N975a.SP:6f-S[FMP(\UK4NP1Z?f5
I9MT2ORe3(=f=BKa;c>Fd=).gc+fO<^(dbZJLR9>ZXX+D+DcQ738&9.FM5:8=HF&
W6>J;bK^29>e6;QY[40b\;:LEJaH9M^DHC/NERVZa(EN1T,g-AObf68;)KA>YTWX
5<L[4Q)g6AT&TQaaG4NL/JS&O-\MZD/WPIELEffIf#Bf8J+@BH,102M[VS+7+]K2
P3UId/J0c/]G\5bGD.DL[,;1eRO[>/X^)O#\)NaFR6K?VcP=<c1G@72Y)eT[4e6H
MT/+7(R:-C\)B;;^+>4-2Rf;9dW)R/U-d^W=_g)YJZV(G/8(>H=&e5#4,JX<]]b#
Dg=B;85DAF<JLE&C<Y:C-dTddLaNJ-,gST0F=PCM]EG9Q:KSJDQIe-&G?e\^g[Aa
K:)?3^A.7.e2XWdDHQ^ac[^bST;IBO0F9_S_?T-?<cTcT7F2_a]G;(-Ngd+@Z5/g
MR0ZDVXdTg4f,A,A2[FWG2AG;e;IAO@GO3M4BD//SG?C]Rgd[eFSE[Lb?(&D63=3
N;+4>A=;+8X9Z5HV1N2VDD9R\\.5+#-S4@6H\M&f\a+Y30Q=1]DF1]YXaC6UKQbX
Qge39^V-/@@R0TBVgO-<J1>G.=15)G/_M(cKP30>-e8Y>=Xf:(9D2<>;CFfMcB.A
:?4C=Y#O[LT)O_?0:06B9H-bM-0;TCZgIZ1@/\L:W3BZ0O7?e#Y\^95@2aXHC_Z2
]D<K\dIH5,e#W/Ia4@O6H(R^b54?.;B2dI1aC1DYH9<RE/bRO,3CRNO0]T.5gK:^
Nba4+I90\_I]CK1DL.0+RJ/_8;=7D034YMAZIA0//LbK)Ge@M&HAZS9=TSP2JIKc
)-5D^Y5eO;K:D89^Ycf:=+@:K4WaRW2T&dZQ?3V)e1APeJ#-X^)(.XPH].AaYZ34
>2::R9=HE?Ea168TI[+S^8fTVVbT(GfXB#b5dfbIeOY6WKdS[:2fB6:2T@09-ECG
C>AI#S@M8NS+DUU3fEUF=gEQeC#NT2W7Q#F@V+U8T6&TFGEX>K75HYI6EWRO\DCR
G=ME0R^g&M9YRYb:F7N8+5T@EZd&XIN2>?\M;CMUGY&E4:B7GUdccS(5+IW[])H/
Q?:-G&9_=2N-KB?YN.5VJC9DQ9W6Y]7-\f>=AG3_GVKcS\=D/+DE:7(0_WLZ0G&>
HO0^NCU\1^S6.:#2E6E9#7fS&.CXb2+[[PL#46/)a46><\]^N[Z[VW.+OBXE^2bK
;eZH[4GUeN.Jg/]NHI@:EJT=2D^4MA1W=V>K-R7MVHXST_Z5C/+:DZgGZ4<N^Z(B
agO0.D7K]Ka1.?a/TQC73G)K/<TG-IWO8VL8VKN+Ka@E9]^[]L@CbLP>)7]X&,@@
G.OTCfIGDF,R)(WLL^Q#3/2ZEFA)J0UZNWI&?HFP;PWMN5<(V:^+:@JOELA/>=9L
2(cD5&>:OXaJX@F&e0\Y?#--ESWP34213<32[f;/FbcW_Kc,a5_]<(Rf3DVT+;?d
+TeCF[-1G+&R+PFbVHaQ5JI/E?D5/f&>-+@P2[0K7)>SH0J4AY/e0&Ig9af;c\B^
BR=E.OY3@ICX?Lf1VX]eD1V7BW4ED.V[4K2Rg5b5W&a_G/4;GR2H6)O:4B7+OBWD
;-VE0ESD(?4AMIfHA1&+Q.T1b=Lg_;9,=.1U&MB#GNeKDW/;XOg]XDbaP6IBAS@.
?J^Y[e_(EPWQ8[JVFC,QT&EZ13#b04ZWT^e&BgM1P&]\BHc;g[R@:XEYKb?<#Le<
adF0V7F+4+9]4M[+-9J.D7aY#?;_TDW3=FYAQe5?\HO=BA1)MT\38V:(K]6U#M=(
&X22EDLBaK/#<\O#DMd.[Jd4GHefKPWOJ.9JgWK_:;9>_]&:L.dONU)>,DgR1Ze?
J&M/?BBG.8L[U;0Sf]W:9[<C@_FZ_#(B.L&L#W4,^FSYHTR7+\Y.JEadS_R9?(K(
@)GVH/)/)[(8Fd3\@NVXY;MB<76/B:e#dKdH=#_0J2SU][eSO@>],]I>Q\[,BU9X
]I-#Y]82O+Q4^??2J2@g\13LI8N4X&)F>>WD5]bf?B8N\JLOFG[6[(\0T9Y8[,Sd
SU64Z1/UJLHGfQ#QY&&T@FPEE-efFO54\NX4>MRG6b\dLTaKYQ1VFffHbZfD4^:6
0&db01g5.&]/X=.c3;(NW<.?S@I?^=U)PY>JK,Q-+:_^U)fa;;?0(ceCZBQX>;+#
ZNMEJ?2ZOJK>b:P7Q>ZKBV6EE4F/WL_@DGd5Gd\,A5WQM\YX[ZKHfVbcC85ff+PQ
cRD2E/C2@C;VW@N5;+Ic6a1d:;f]EP7c0f:J3G<CXJB1(Q/I/4EK))2?[\c9&&>c
UAW_dNK\W#D[\M/M=GK(@41_,J[]SK,TRf,7@YaNJfAb>4W-)<05eOcN.H)L4V:g
?ecRG5BL6UL@gFNV-[,WLX<F;1^-XfNVDe0WS)_WQ,^J3&+KQ4e41fO8(DF\&8G:
g3JWe?)1KPYc5;T2N&G/IOe3+^VPa=B+X1UQI@[+M.(U9_C)e-)S^:#:#NU]Y.FX
AM:T/WfA89QT6_fP]5D9HBCQ(:gK@,Ha^a4/;[<JO?)?+d./T7e:W9^@ZY=Hdf+M
K]SYH\-2gX]>Ygf#?/,LbXb;f0O)#@1=&NLD_-R#GYd3-]I=)[@]WYB0\[_&TL8]
PR2.:R]<?M.If&5d-4SfT8e#NA\N065>cN28/NbM8SWKR)aO_W60fe8S2Q]dT[<5
bBXJTZF-13Z.8C9U]A7&/4=UG\HeY#/eP6cN2)=YZIC5Q/g]K3g.AAW^E(c)4A_Q
TSG3a+G<ed1^.Y.c11YP_EHX:OCSVD16OMHF;@J(+PI@?G;PK+gT]IGFM[YZMWeU
a=f^,S4@Le_F+H-:a7#;FMbZR/QVKI)_8&)/5c)gC_XcPaIC)8+&Ybd8XK/Z.If;
2XMDg4VL#:HY@Xc[6/G73XH;VAC?5(f/.C^fMQb(_WYVR+&1K&GD;TP>54BJ&/.B
de#],-Rg=Q;(]/b)gZ<W1LTfHe^O&EATX)dK:I#c]6A9WK7@J,g>9ER4[1..Y6D?
#TXIB<a>9WT4b]MV20b36;c0C5DH5RU?fV;gS-2JCH1BVaJg?9ge>f.T]A.N@)T.
7:H_@KG>0=.7Y0dRB146A25?RR\-000F8:WQg7@#WKNKYDMRg)aS,LcdQ&]R#A6R
BG^H\JgIT2T?VbR(J<6QeJbL3&C]M0CReSPR.c1^]RHL7ZH4UKAI.9F>[/LL=@dP
/][Z[ODC+TRET+Ic3<g7LWB](O6?7[4GgTERag7^E1Y>4cX()32Z9&7^_6K<bTd5
+gU\XLV>MPCd@\CFb31caLQRH+C4_3^DG5-Ke,URG.CG_P,@B9M3g2PHCF(OFF96
K>]aTYAEeZ/EVB5XJeW?D<ADUP-)FD(\U,UbP[R&/S\L/2D<)J8NL@XL=BLJCJOe
MJ&B-?WP+9<JCHZL(/ZKM[W47AY7W63QcI7[/_#G1+W1WTB;a#d^]//UN#95ZM2:
51VM_8==Q.=e8Z^#(G(\<#NS>\E02-I-)41^^dF.2Qc_HL/\PS_bT(RGOG/f@,5:
Ce[P;C;T8:2M1FNI1BX2c.,;fDRd,YVXaTB?;Q6KF,1eE.<MONEDKb3ZOA:PfK2&
5.AXJH#K-#L#=+Ga.W(Q>gWcYW.EXQ&7QcN,4b?PS1.Z=^6YXQ_&Q^V&6L[(X2U@
?)MWU)?(]c?5)PKd)R^=A[F\^9+<ZF>6E(bZ^.36>GA@CQI.6:5?)<SZd)/EV.Z/
.+2ZeeC5/HPPgcE8ZaX70)fZ+c5WWOca&TOWO(_MSe:D_CbK=:^O]J<VdN3T8I_b
T=eaS;eeHCF7+A7UP)]X;H=X1_f1VI/,)b6ecf>C00.SB9D0F9^GO2+d-B;^S(06
6,25MA(Tc:=;;_NYT;[Z1S2;:QDHA-BKg31fR7M\J^+L@@..)=<2?^afe^+U)J/Z
=4,dQD,##+N@dDSfI#_bBG0bVH@3)eX0H+XELQ6N\Xd]H4<FPOCc>QG,TO+c,93>
RAPFfD(@6(JF7]3IHc[WX4W](X6+<0FZfP?_UN4b<.XC@1DPCJX+E6@<.a@9(@g8
S&X6;93MeM&6cB)O2&8=<D9dgR?>TG,UV1(T&6+I8N.\CdPCH5<Ce-gbT@KefZb9
11a,0(1((XLK:Z^RH+Q\8b9gA?)Vg4EG_:94C3I?Q6@_=D44)68-Xe:E;<fD])H0
[V:G^g#SI2>Dd62H(+JMV^7b-GPg<(QG\KR/@I-f&dE+57K)>#/D6)2.D_>dTd,D
TWZ[U#:>,E0cT=4>A+Y;K_/0,8.P439:=,QE?3#&1GLGTW#B:d+FSg:<JQO.=85>
?H3C4Obd&256bSXZd1M5Q&&<:F@D[fXH)UAA0202bK+EJEP.Xge.H8HS0W/2DD37
We?UaYUB&\\14MYFbT=[:YX-WRbOZ3[;O5P?\E9(bfaQV<Mc9UbbOY4?D,7S/:91
^7&QKM=FI9T/+,?J3f(@\SIb1aK3XGIU1KK_=ICR5-A4eP[3]KM>)&HQ3,,.GH.^
XIWV/UJeee=(30WX7Q7[E@08W;957;LbcFbM2,dE<,/fg;cIO7V\J+0gO25e[/N)
c1->U,UEZ(@=,4c8&4HSOGWX\0PCVVLZ8Fc@Zb:R-If=6Ea_c9YGXQ244-,^.;-(
XP<#\,)<AMb_=)CXP?,DM=K(<&aDgFMYS@@4X@?KTQWSe9fQQMXe]13C/0C4YS26
e7:&:.>I23;)E@MD?\N/>;9Hc_^,.f8G)4@]_?H3Q5Te?3_?PB.[P+(6Ca75,f;f
XK&U^[BC]b<Z1gXQ1fC]>T9M3PHK1[VUWV_0AUV6,(9+X5[0Z[#V@M;QG+P)/SJE
9.HS)[GVWSTe5HNDLUR.M8>F:+A\#=W02Q]<Y/J1L?/<_8BV.@NAIX-Z?1]DXRRC
QKSP??@O4;440gHWUg4G2ReCN[ZTbU?dG__=O0R?\I#O4I5YCI^_e9g-3MM>+^e+
;HMcI]8[/U;35VJfS.Y(M6P.:/E\]RW8:1L;Z1:)gZJe6]4]:d-G,U)_VQaZDUVM
VcZ3bNg-9B9+W\8c\6<?W]DQTb;_K8=QL2+.dI[MYE\EN:bgWDTaBR@(12)AcZJN
9KW\+N452\@\&_(Y@0^e@P/;5;O;e>7O)CUQUUd=ST2,2]&A;S],2cf&I@4RfdI)
AV3P_ccXZ(Z.?:C+AB.C2A/XA5?VEB>>?5f\V449^VTH:(YcSR+ZcdI76#8PT;P?
;_)=81\fS[f4/BB2cG^QI]fT38^P>9UBHCHUgYR>RWd[OX3K7cbd@87:AF7/Z.G]
59Z.)9T1W\e^7_b7S]Kf-P]]8/T2YMUEBbH,MX<C]#27B+7RMc#^6[BT)V4CUWPL
4)b\8AQHRJFR_XS?2QKMd+GeKPOL,]D)CVTWEH@G:5BRN)6N=eQDUeN_7f?B[W:-
FU,OdEb=e7G;b=S)c2C,N8XI5@L;_)V=ISef_[3SNR6,+Na6TeF:PBUX-1E\UJWM
>)eZ)&3M<YTE8Pg?=9353#UT9P<#>3Da7F_30QR9c_&Z]5@6)0d9a=ScQS0,^MR\
+N1C>KAR#_T:<,XR:HH(,b#d-g;:=H7OR&CbRNIYOZS+-K5\98+&\1AF&UJT=J(J
6@M+d&WG/NP-E0XX;L(Z]?-2a1+6,EQG=4Z6eN9\bW[EZ@c,b#+P>eD:209R]DFe
??91b0(KT&/H1fJWWO3R4-PML-#Z#e(JK-aAH/HFYS>d7J(bSa3=.99<I28J6>U8
0ZDK.HE^>O^N8N[SZ/O\<<8:&e6a#5RFbb]>>W06UA:Ie@ITR]Tcfae:.QSf=22&
GNTS,I3=#OUR6T6M#1KMYE=F<WVL2WDF,.-Becb].A2S__<WPYOdWJ_\AB115-fH
8X5#63(0ELE5bc1;&6FAQD,<L@OQBf5g0=aYYL^69Gc^.V4+I[dP.WE#P6FTd-+\
+Wf(X+PEX:/9?E@gSMVKD3B58>(@8=DKH&#a0D@d&b2J8Bg2=c3c4FV<1Z((7];0
UTdX73V1MB/7-F0A:NVTcEXD.[[A8b##NV_;Hfb=a@b_S?._(>,+7(FB@W@9Za2J
]BCN<:e)W4\Ab^33D=fR).?JIL/<S90GKA/6W,U(.9Xf@DF)9JC2.2^&<[Y;J?&^
,R1?O8#a(8PbS4dG?(PA&4=GHe7YaC^AC)<&cG8XF8CXO8?XA#EbK^-eU#3SA)5V
(A<GZ9R24)fL90+2TZb,?J-Hb&J9.bCY#@>7I@,.).<))4926bPGfBgR37^M5W7]
b?4JI^G=GDV-0;gRG58\RR(Z.3cM&[W[1E:XWJ)>&IEV]_RX3EcfK5=6<W)//:&7
5>bd<8YAcKUD9cGDf6E)?\AL(E.E7f7;gK.#Ede+F(SINE\U>8O=MYCGWQCE?A=P
Z5gSZ;G[IX)G7^b[0L3\2,&N#0Y7@(_QZ=U[U;fY57U4,dTS,V\O;gbVQZ\J:7aK
cS/FM@YZFQ3SUe)MCQS^ZQF\?Z7F@8,DBI^EB@19(=&Kg6#dO9a>M72M3;I[2)+g
ge)]>.[<.G_E,Qc@14L48Y1-Z,c-)77gZD^R381H\GE2D(&._V8D3(K8-1eGafSY
Ee.,KDZ^:KcXK\U/JX8\;^]TbQUC[A4HAXKgc=;)WY(YUI4:,-..#9UM16LaGAWd
0_88=4?_/13#AgVNI7cH5/6=?,CY5.L=>eN[R)=4QKXe16.G2V@+_>[LCF3_+0\&
\YW+:SMef6YEKGWEB?^GA0@>[1.:MDF2D2@1&],,>A5&6cQNZRg5J1a>D3f:?fXO
4N#eB??],60I(.64NHN4bR+e-1Y<P?#aRd(RdUPR7>4[+GR0W^KS1Q0\465P0aJ6
gLY]&(/f>X)S1A8T84P=5KTKNSL9\6+Q8I?edMgbR/5X=f-cDI:0a]9]#&NJe\5<
[Ed)K+GDHF7IP5,2=3;46U6-W&FLd5VA>CN91M;P7^,gC:GWJDfUV<EgB0d[c-AV
::#d:J7CQT^Q-7,Cg-M:2df8EX-G524:#BT:1?eW&?=g_PE<-ZE<,cGc^ABcTZXK
9XQYL>YH0\>1K^dQ-2P-4;)OB;N(:XgW?<&LJ98FfP3=U-_d@HM.0e]e??U@AXSH
#4fL4;f-f@LI?eWM0D]eN:)UXgaA72NQ)M)^(2NR_dTUa],GJMd,5c2fFRPZ7a9g
.NUEI]0e=0MgJEGe74U7Z+Y.[Y[g53BAO+PNLSI1IYCT]>D4-09)7N^X0A5[&;Z@
X[DMO7TgAf=W<QDK);/cZQUOL2<XUM4URZ/@@SaPHN;gJZHDJ:4aK#JfE1\;+W6c
CSM\Daf>5:>=5B8A](G>9^2cCHAV?dQDR05g&R[cAa;^E&>N0?K2EBJHG?..S9c8
(f=LP4\WM[e84BP-.^\d8M?9LWV64F/FPMTVN_H3^S=R(=gKE]?F?\^-F+87_[^A
(X)F6CW0ZfD/bAf6NC<POSEDR6T>-6f&VY[aFYB5<\WIF3[4W5HJM.6\#O[V0?9V
dWPW/d#>EH7a#[AARQeXYeB<NLHI>MJQfL?W4O4&ZU\80eS]ZB2^]+TY)0BVPf-3
MK>?NZ,@^e4IG@I\?BG27XH>NSUM:=-)FPY<<W7P&gJZ3bDM>MbT[3/0XD[.R^)K
>=_>)-b)&(]7?+L&Xd^J24@92(]PXMaE3/>2g&BRcG0aAIaPCZ<_D:66V_XaaY-K
6DG<M,3@)Q;:[EFIN?.8eIU493WN_>Q=-DE]2<C5ZEaN-JJ[1L@WfGIH3ZR1/LY<
>5G-fNY#WIgALXF)FP:)L8YM;WB\LM,8Ld>H[LS+e[Z5MT1aTgd>QTU-HT1Z&F2(
3HeH0?)20.^/#<9/&(_K5Pf^4W:4.8>d:#B3D?+H8.T.4Fab#((SF3fg^\(,?W38
UDV]5FO1?>0JAS)5ePQg\(].6e>2I>ORW,Cc?R1bKUgZKg29,FMF(\VEJc0bWQ@[
(=5UCK_^\-S\(:\K<A6MYa:gTLaFd=U4JQ9KPA9;@+;R_,N4@WCg^/;BZ^<&?[+^
e644M3Q^G)c\ba1N1Q/;@S/ZSXYKL+?ae_#M#M,CF8BE;LJ:\CS2J86_cUB8/&Oc
<]^H]ba\6fd6^EA;dKbP@21\3FKRGa#9GeAH0G>MZKX6]#.M+\7TbAWHBYc9]&b<
X\L4a;Y_DFF(WYQKGMQVbZc-QA_=caDg;@&KQ&>3aOS9YVQ<c:-FV26?EZ4=,H6N
P->NeFbf)^M<Ae2,J>K6EO_fG/Z0Z4\G_B5BID^>FbFK#^IS]25_79NOPJT)=#cJ
(DL83IL9F[52=U9f]+KZ\cDB1-7U.aZK;1T#UD?J1[H=OUB.;=]C94/.0O)d0)9]
.-\M/-VMFOL]J@,be\RcZ0;^V^).A.\UT1/9Z4g/TTaJ>]fI,1PMY?KMQdE][K//
ZDe:4>[aJ7b:;A[eX4AeQP@Y]9GTEcc]&23EA1dKg2VcKgbD7SY&Fd,R2[Z-4cW(
F>4dg#,\U3)OQEU?X+9Z&cV5fYMKQ&VQ/c8Z3-.[2SSY+SIUaEYOE9JUR?NC>\W>
)U,7WDL>_>D7-T9YQE-_ITIVV.d?A&Yf@0@N29HH_@YJN_^R)/PS;WE[5Z.Lfg?_
GU#d+H0A2&(R:V]GHM57V9SVCca@Q1VXOU2Z)SGAGbJB;E8;EJJ&KX9&M#X#H?X_
IO-ccDAQB;d,Ffa@O#[\4E[O7LS0[ZdEdG>H<FQdO9>#I<XDSE[I]H<\S&W=EAA[
P+TI?+Q<XYIJC0DYQ^[C9ME\_;G69C(@4RL])@],G?g(SYZ,[>a,PG986e.S5E:U
ZF2MfHK5YI(1IG&))SNL3JJ)a@ZX,V+)JA9<gN7TK-O>+CQ_E+^1/4Q#cW&Bag;f
6(Z47Ie0HYVH>93TDD<KFYO&0-#=P6)>1]#D,LBaNaN(6LV0I6E/aYH#L_CQe@Te
\aEJXe&aS_?AXO._F<\-fCW<+\@]D]>,)&VTOET2(A0J9e185f2]:X)W=Z3fQK2?
N1&)U[VIU&.7/1c@T9(HCgc^DKgUAWY#RFa&SW]0)?__ZJfb4R:&d[@>0dd0H0e:
0R.P2DB>9FEWcg)B7<2C+236b^_(QO?I=\Pa]U#3XD@GPL50SASKfZ1d.#2_-I]=
Aa_[&2KIKSQCK?Mf08(771?#Lef\[KX[N9d(#W_+EE;;K>JcQFZCRQ@&:]^e1PME
VT?8Y6\^KM7U_027#OP[0\d66+&7G7aXbMJI-BHC:3HX8DQ\1Je):4:,0Hc)Qf2+
?6UM+bS/3YGbXBS6))??)90PO[(GI?--(_.85G??3bGPD4/A?gB1d]Z#;)-e1L\\
]_LLgd7:ICPJ\=\66fg^>W31@IHHJ9D8e]-L?)=2T3:QV1b5W64O+#[3Q:E);.Vf
+O<cfM4L_\?gGD&DKJJ?U8/=:D]&(NH-IX]KJ])=dPfOMZ,#[GPR8==0Z?67(W)X
3COHNVNU[I=[:@J5<-B3?A4M_QaYG\fKdDYHW0-TB[Oc0_2BO-IeW82:D>&MKGa+
#TTCZ;<9A\&L0_XD:7NY?,MOQ#/=e,WR_H&6V#MYY-#60M=GMfVaXIL@P_^Mg\f_
9&4GQD@LFNZT1acV:44)/7fZ[0AeAWN^IW-?f[EBXeKA]).fUEUM=#\F6?Y#PT@?
cXE4O(5fa;IA:ILU,?-E)-]-APYd:VR\AW2CF4,HQLFeHPF_9+48@5P#^Q\g+eNK
-X>Z6FN8;QUg9[7/-T_N/>5.ZUZ&O9C>?K7GfAB9DNaNWPQ8&\19WdT]&E_c[BYA
+9^C]M9^2GJF5?1eRaU(>>:@CEX>.fDG6/UA@Ba9&d4@]>T9I@MZ:N4dKT4A1eJT
_4LEY=CQd./F3L;?H2GC,86Q#IAKR(XO<#/L&aTgQWRF;R2U)L8#RKILH,;-FafI
)MZ:;TM/g;bIPB+5;FCR>@e=ZBgM6BVK)X,7R.F>].dDf+5ceY2CZ=M?7CW2I?0;
_eUYaYCSL3Cddc7V9;/5+VEPDgX/+#/(8.(I7LX#TSH4-(,BPNL^VU840N>(1O;Y
d=JHLgfA<>T24c@3fRRU#MR_N(D_.-L?\IML62cK5MRASa31LcgM18.P(&-+8]1L
O,NLeY6cA,44gGRf[dS=06^T_f.+b4D=^g]E3G4ZCO2+&NKZV+L/#/&9[&RER_3(
)SOI;+YM?K8LR6F?O9;@6C]f_Rcbb)6ZR_X>1IP>&IS2HVJKY&A]Q5)[-8b]YJJ:
:]Jd63H?6M>A5]AAI5>9X-:?g&VTc456GQ(38fb_;R:,ePA-HFAdWIIYJC9K=6Y2
)DC-PfR_,gD+4cd8V(:c;NF<UI=P([1NT?B0FD3gVE\)N&RBHQ2^3+:&X./UYe_#
8>02;(F<SFC4UdYdfa2&_@4Ub7H,W<OWIK]_3JMc/ATU<M#.539g@5f6Ub#>aWL?
QC5.<\IWZOEPU,M+S.L-e-M2P)5gX7>(=e+T;?^KAZe+(O\OX-G@)6UaQg=>KZ<O
MLg-[U^OGaeVJYSU_9SHd0D+/)H.]:F:Q+BO+4OW4>&]]4eJ]DeRC)40=e5fNUG[
\.G@dZC(4VbET<PNcPB]W)G.S9M?/]-58cW4FQb&LWOXHc3VO7J#/C>(b8@MQJM3
J@>Oe@NM_>UQ@aGTS)/Z+S79LbV:C:BcV.BAD-0>U&-5@PK=ZcBeWR&/LDEI183:
N@)0XS(/LJ+36[P8P&A]BGGDIIg\FOB2+]MC31:/]<TL;V[g6IHN^EP+,PVGUO7T
KR_(JBgd4FL,b?-585eK0fLM37S9S,+3#=.<@\^+VHe5??Z2X2Z56dD__H[A\(LT
1949CL](CZ43O>V[@5b#9,XE-5GdMMbDB1@5a8a.#Q]CD/9CZ5?ALJMgL0D;bX=8
=f]TCJ?SP75>e(QDHS10;)bVVL)(He]ZL@fgM@^gf3ZCN,UA9<8\dM&M1FGMbZV^
NT0DWbBcI-9fPSTT9R-e.PMC=I66YFR8dM_5F.GVGVRVU\HKBY)R=BebY9d]7H)/
d1]/P1NbWYb8W=QMTBP3?):0Q[2;TR;OG.WQ[^YdI_YgR<1D/I@EcI[C6F6,=.K5
+Wg@\9^?aVF(3]#^g&cS9N=ZGHK(dX5WLD.6PRXB=WcUO-WN=)c,KT)AfM)J@a=6
Kg0<32J&T07\,<\X^MK+(=6DcEIb@4QOe07KJ)Y3^?bQUa(g/SW]eRROH+5?IH:X
^2GQ\gA/GCD3N+G9d/CMa\G/#d8T)@7H1M)<H1=c7_806DPCBD2[Cb?a.XVb\@=Y
83d9E\eUG3<K>@:04cM<T]7T[2KX<,MVN-S<H7CP-K0&,H@&03_N.]JbN(g:ZX;O
?;IT8ZQ6Hg;5D_aW+E&FRa^D8g\G)(0LQ75.>GYg<85,-?6@.>C@6X:IUVS;8),^
FH64FUX^3a)H.gPaA\21?>:A79?IeQJ.7WId+cYTJ:D&9S3XHED1J5+PY:4L-[3^
U6EDG[ZP0F:M?[@M;M&1a([)+:#aEa@[HI;e@0.+>4gbWa+DCRWUCdF7\Vf[@,E1
fc0K\Q8SKC4ZHJ>cJARTSRB@G1Y?H<8+T4TL#d=QP?NW/@=.?ULT6&1^?Jc[+DLT
_FQ<A#AQg_(JUA\#(4g8UDEEOC3Q436HOc(0CEHC;SL_/0CI95&I:Vf#_(I:a53b
b_;N6+;[A>:_E\X4DPK]J0^;_+>T17>-FX?[+K+/:D?aE4MH10eW;A?b7SfbG.OC
+_G-H039b=9=PeU@NB?X>66)30I^L.WR>TS5A@8d:EFK)GP\d;;K=:]5447X?a+^
X8-L.4?G#,a0?R+-Sf:db[\A9]<a5(8>B@LIXe46A5=[L9X]705efT>&HUETcb-?
f8^TR,[#edT9]eJDJ[K\4=,R&G:R[cRZO8O4IgQd]g6AOAZf4F,0[3>;]/X0ag<2
:PHH+^K6+S#I0PRC4,<OEDbLg-Fc&bgTY>A^M5ZZ]RM3AE)c>gDb04BBb3DQeC:Y
V[CgAE9[#6L&_Y;=O&DYSP+S4[#->RTdLG9@GO58X6PP1fN(FEF)1MSgA2CL:WW?
\05<:5:Hb(Qf<HP<6eDQ[8CgUCN8HSd]XaEWW@M@2f,FPE(e=,]cA;,^A_M8B&HT
IQca9A-e3fOb=5<VU[(#BXRGN.IP8\<M6)2H\2R6g,V1I/4cNG^GG#D:\&K(=UN=
YZ/]R7T?LMKcAQ=(XI;fb(N/(DR-._JXQJJ0UPLd-._YP>2>LAXU^2dIP</SB>EY
TP_b^MSGU[]3MQLe0,KIE\K5F:_GZe:596:Q=]>^@=MK[dVLa#^5P@JZSN[677:2
,Sa9#Reed29CY,).BF.-JXe]NLdJOc6//2KYWB0Q[A3>a59SK;__Q2b7e:,0=0H)
YLVg:8dcUd_HDG:9,O5:V[K_S.Q6<&8TDX0B+VZ]f4\,A7L;<ADXC=+6g=d/cOO<
:+(1b.ZRQ=Y#21)cd=b]V44S.UbQG];.fHROGXX2A^O@B6&BD[G1QIA00.,>\eYH
:8_)ZR+XVAZ+_3SK]BRW6O?d??aV1(2@(0=62.fIMBTZI:0C<_UP[[Y9:#[g60G:
5A1#GV/P5S@eE1)bC&^R.f&B=a>^5[,^2Z1,1e>^PNP3<gdX6K0G[(]C3L9-5H0(
P[LD0#ScB/.)g7?/d.KN.e(f+PU??gSH_Y/g)=NFdWP0GX:+;D>:#YE[:;^QKAO]
ALNI>c#ffC>g]G>DZ15KcE&+DF=Lc@W\2H(+E;:.V-Dc5J+d&@XgfKb1G\0baS(Q
O3,[/WWbM&5?5Rf)=PF@A,C(Z>OLFXH(37J:AF68(NIcX>OKBFQG(>(&N(^JR;^T
E/L>a?Y.66.a8-fJ\TLUJPDDQ1C9>FHe+H2gBMZS)EaUJR-,<T6-DRcIAT@8T<7P
?3KK^&^c+Je[)MG=+VG<V6V:DGS\)\0Q9NS3<3@::ASUQ@HBeC.UU:W<KN._a-+_
F1.R@_5,c:#WVN2SXXU@)1eK,SQf(:(E6#(7E]O1UF[,IHPD??6N4F<59\<Y14bf
73,TeP[>T&eOII(>FeI^F\\N.YZ\TNS.aUT#MT5(Tcd=dcU0?F8dSf7/&Xa8VBBV
:-N99F@\I33#XX]VNSgR#K]Og.LSM/_OX)>VbeV3WZ2EdUeT&8[?:fM?EW1)X1V@
c@_)WJ/1VYS<8#OdBK[W7#0<MI?EZXV>3;D,-/^YN+;J8bDPR>:\AUdON<VaX/2J
A?&3UG<H-RX(.H/8]?:@U?MV[664a\^\0=RFKT@Q)@>e<0bC\5Y#R9=8^M0N7=gd
W+Af4GXX7e0eJK)(&Y79N=J0TD.1E_=7/UP+5&c4[WV6?eU:SG^4#Re)[[?1fcF?
ZaTTW[.B3E>7;MFTE;Y#[LEbL>X4N-I9K<Z6JJ>PNQR\FHG-YA[UD]^8SP#c]U79
=7YZe<<6fHNK5YAI\B>EgG_+&Uf5F8IU<;_\&LN=ZIT^<U#^g]4e#,UAK-@8X5?W
10H\H+LF.JPEec=+G0^CY)>PbBV1b@\U/80FL]TC.:7R4JJT2XB)c1eYRZgZb_A6
^+WQfN^/74<?b4WY,fc3a8X2=ER5TS>NEQ/PP[aO^c/GeLPN3<(WQHAM:\>OP/NQ
5G(AR7g>d=K<NgW.#gTOF?]^2QND4?W0d.0._:4M:HK[+;9Cg8d(Z4#KbYK-DT?R
La9SKT:QCCd]:V>[E0P.AKF:#D#._4+7EXQJ<bH5<AbKTfSeK-T?c/NX_<15c3<8
C55+03NYKAR@665<T<^P9;dVS3f;2,8C_d3HKUXF8?RCVFGYD7WYb[cGVPSK(1:d
XG\^H^&WTN&:VS,U@8V/e<68UIHc>M8b\>-\5HRC#^GL.2<6[T\,.NLdcbBYQA4\
5:,^c5J;g?b(V[MX6+fI\9TK=2UDCLE>4#2#\/c8&,bRA1AA;9WA6FL\MI@<dV77
cJ(:_D>EXbUYRC<-@_G6V#&ZP7RIBWL.82<N#?VVKb1e_=)e:6a/R.R#\11NYc7N
AUBMVQNG[af,eK\#Zf971J#,K=fTCMMc_,CeK)0MQE,=5C4S[:;_WC+g,UEb5MXf
7-5O&;B<OXG6S<1HCR8]=96IG??BUcT8B_-LS[K.U<Ja5QK3Ff+8Z=NXT#/2B8&P
-8Z64__cSBc+@U#RfQA4g34]1aKBV?g@GZX-A03#\-dbRcFZ;HOU^HGSJ95:2=Hf
I,OcgRK;Fa0-K&N?-[IT196Gc.ZYWS]e0NCRP-QL84L^3?>_FD&^X?QJ@4THNT)?
Fe87g,P,C2#WC6:9ObEP>f9KaTYQR5)D8@\V25TAWK)&_?@]C,;-HJLf81FF9<dD
UY52a^Qf;IU]CJ&_L,_=C?O>,7c;4?77:+,^#-Q^fG3W1OT(?#6/&2N8J@W8@U[f
7cW9:J7.#PUCM^4LaV2A-7HJ&YTBYc=3=\0-(,51N.f4O+JMV;=f8BAR(PEfYKQB
PFBBS93)+Q^J90[G\;NQg&&[e[\S[8D4GTQ6.<41)3U(1bQS_,3CRU<RGFM#@/Q^
RV&9UK=^[H6)^JQF[e:KL9&_]8e7#cI07)CQX4b2&2B=?eY3LM6RR(1T(e5a:C/C
dT<\O;0TRF&>)^V)=K>5H;eI9OGJ/\_53bMS?;CS(???Z1,YeK>@+Rc_E7\OS0NB
4NZ)g>(Yg^ZDYgRVB)TDGU0__ZV/+Od&BXf4_BM[LF;O:DD;,>O&M2]9L^4RKdU3
4-F_&[_)WGEe.]>1cPg,Ee:f)a\MKZ/(+<]DCd#7E&^@,HB6]\Y0fW0=AOc)G\?@
,Id;:Z(b/)3DSa2NbA^TF.7fSXWeWI_XO3af0)5,E7_Tf[+1c@X:<0MaUA2YAD[Y
W0:cNOKJ_Y#7V[&)McF=[440ZCGEb-Yc70e0J5cgTf;6R(DVe24^Q1=Nb1ReBC(G
K5<\d@&GR)Y4<dYI86Z5:)/W\0ggacTW()5ceDY?IAg:T^3_AK=_]89XV:AM&75g
FF\6#aH9:(AT3E?X.=S]K:POfFS5TH_UC>K906SgC(1O>D65;_X&fDa#L=1D<C?U
P-1/_9YPB[^>W/3C->BH=N88VJG(I7\<D^9(JKe_W1e>D1,PB@gR,BAFJM[S1,gK
G6Cf#G30[P(FgHM\g:Z,.c+EO:74\(#(L^@-P1N)(FP,ffJE@\URX[J[8+7K>dcD
YBS2B&S#YM.TRW:<:-eND1YM9/3A\FBA@WUMDT2SC]g(D00AAa[K/L1&M7>DLPT-
<P6+g<J.K;6-?NA8>5M0XWCC2BV^X@0O=J;N9]3KW[.PYD5I4\-LE0O:YfI]EE3E
P1YZE=P(dOLVe\(QcR66fGK)LFO]QXF4MENbO\DRWN+JBT@gdIfKa=JF7(2JgRfX
7N:Y.>a8&B0dANeC7GaB[BSgffXQ?0N9Af&a/1(ZY31fK;^/R[)2#IQ><0@AB<)c
c[Z5Q4V:/a9R^Y)3KZ((F=85\()f)_C=U>V#JQ<YdaNZSN.S&:ggL,34#f8cf5+a
ZJ(&d+7&Q^8Sd0CC<S5Z.PCP3,?\6b#fR(QWMc(->J/F-(5)UTVN+R@?.@+5U?N7
Eb1@TWN#M3GTH+<1PBR;3.CBe9/VbFc1M2+(7_[:;,#bV/X)ZIBFX)SN<HT3;:@2
9PN#(d#PHZY2>GRT6-^9/YZTNVQG#R\EA8?B+ON5_]OHfN?gDB4g9.#[3_T2^\CH
JR\KY\/TGeZ&8c>N^E^S6G=+U4>?F9g&#<N]][&OJ=UG,7-XDX2RNWg;M9H9a13L
6?PXA.#3D6YdNdGA<.;Q),eK-#+ZL=A72E,7cWBM1Y;7,3Sgd+C/NE>KG)-;gEBD
RXeb3WAUJeF3db1bJ_@F^:E\d-=\,I(c,JMN#Wf;I5YU0WZH(G-UDYJb^[H?0>?Y
N?CD_34^AF4]@+.Z+dYFRIKaF@>N?8<SbIge;U(CAPYc-&[9U=EM-9a4R6U>YCKS
<aX(;R^OaXg#Dgg):aEeWS=)eQPIMN@EB^&@bHQ)KCWe?ZCU.+]W=cH;T9EQgJ&@
bQ_E[N_Vb<)T<TOSVTd_O\AKR#eP3TXQ(eL/NS27]4gIK3VG#KTA]836G:f8:-G;
VSd;(ZTDd3^VHL;C,d9_JC7X4OI_Ja(;.1D,N6c)3N#I/HY9U],fS&FPNY;VQ+@C
^<E4=7/S_690G3J=.3#/8ddP4LeOJO)/Ae7)>\SC5KO;gSGH&62gE>H9E9L<J&++
+dVYJEM#G0&MNV(8O.fBWJJAfV&YO+@cQZdYc-U(/_.7HI^>-AI29N<L_D5:+&SU
I<P34Zf[3YaN.GeR^5e=I3@g442R]Yb[B_/gd_Yf4U):W?4GTK<3&?\eJ0Q[5J,2
YeVFK?RfR9aU5a:H:ge5Pc_MdDL;KK[>DSaVDOJYUdQHGg4a#[Xd52?3:^[9HP-G
1148R=)I0,)E[SdZ]g36B8HDO>N=+e&IW?&;//X.ISEcSIP=NN;,6@3T9IY;7K#0
@87Mf<2WKMFUDVKD+@C:LKCAB^0+GWLFf0G8JT^YP>PgR.e<VUTRIG<K(;Oc3TYA
4,D(2HJb7SWOX0#[U.7[Y2f=--W95<Oe2JEA^5SH(_P+(N,#KJP^&EO:^8P-=>8-
;fC#<+6PEN2)6BL4+ICF1ANIBV+(L6_9V?g<)d^/(VPF-DVc6A?G]JT8S[<\RV1f
8Yg-Q--=2D]ZM5WVGSJS;eA@Oe8H&BZ^]-0O1KGN:cV4<^P=[c=\4f-W7:YS;DV^
;/IUM>;5NE\K:@NEUYKLRd(1g9_.0GZXI22TfN3\09(:>2T+)OL)ca\19GS4FY\^
O@HJ.96:+cIa+La3GCNC?4NCg;&<?5@&AB6c9(BO\c-9:6Ce:D,cfLb\\0dgN/RU
WWgQ;7.V.YLPGbRFc4)<D3HcCeJN//:L=)6J/\VD9WLAR6WXS4aZ7;F[17F>@:9/
(H1HX2BET.LBIF:/3JGC.T5gIYSb?A#+cZJ\8GL:0BL)&PP:.eBZ5T#4ALF)F)6D
.-]#;ICL3T6OcdIL1QZE^5+,AI^=MW=4]FM2:>;f]Q61>B(N:aXMPS^1K&2+.&P_
PF;,U2M8:OgZagC]CFg<SKe9YY/3A50_)_BPG]@&]@^TY3^8VX@<3,<QM)L.ZF2,
AQ@+MeM_\33&#HbCHQFAeS\\gI17,dL-CX09[?eTA;4fUCM7=FK6cK6fY3DUR))#
gXU2b4RN0,EEM(X^W,^X)dHbK2+R#U&Jd_I3@FLc#W\9H7SI+a;Z?OgVDd0JT&];
.B=6_&]f&ELa(=8(2@FI#7L>7>_0F566cE<PIW<(\+AIY4U=(H[[b]8[DD</#f7=
E<S[EO7#S7EQb>(</0JHX1OAZ41DLg6f5:/NCaJWI2(&S[YS#J9+3(cP@YIb7:8F
BcR6&Lc,dcS(XCQJ#Q+Z7BXB;W?W:ca)6>E6G1Za1>gW(Y4gK/O<gLR=@J#27(7N
HeXO(QH\f:V/N5XF.ZB)cTc:P]Wad_Fb5E68<:(,B18U=U]a9#ZXF5DZOHY-Af8T
^\^c1=;I2FgDZMG6V:Z:?N1=&J-IFe[GP[HD<L?K[]6Y29e>/8I2?+KHZ9]T.(MG
:N1Z6GM]6>MFV.5W#1+<66?M87UX@S65\T/aVEaN3@O-X6.d;^O09,K3?P#dgAB[
VO)]W4c&PFgI#J<&CKdg-c)1_ZV[\U.)(VC@1@>:;STV8;[,^PeFdeAXV(WdBgBB
-QC\6e29dc;GQWK]7GaX\_;26;:8X)5_ICO(O.F]RV8&,6Yb1NN2Z98V#DTC?DZI
];,::5f<AK5=E[C6[D)22,QXC#bZ+))@PFRX3#bKUYCX&26,0,Z.17U)K>DEbf)]
f3[fAFc;1d1.JB#_OS3I/S9N1YA<+9&DWPN#RD)]6R]1O/2.OKGV0=-DSB+LOb@Q
[T(g4R3\?__3R/]g&aSG@=gFLK+;<CC4I<FEg)ec#4Y)C,NW4#Mdg,OO^PUIOJ6g
c3K^<<@<7RIM8:E#/<&/LT\WZ&K33O;a>5.(\@E508W[J>^W<HVMG<)^ZY0Bf@R9
2(/9<W.IRNP+C)\IFL^CY=f,P0M7B1_,C+I-:?2NTf]GS=(PDgHM^SQ#eT&<ad[#
MFN;EY&Z57T?(<1>@A,Tb)WP(_#T8Rb5[QebPeJ]PX0]7g?QID[MU0E-4b/M=fTg
USKM)5VFVM15NdUZ;<6V]MefJ+.2RMbbWgL+TS-WCgcMc,26NY3N[?E,,LYQH3_.
_&LFBJ8LU(GeDW]=QG<B4>L96H:-YE+]NXg6+@I)J<=J.##,aOO0&Y-?9=[+MZQ,
b?UTd9LRL+5DYES1#4O#]1\&1(&M8OMF>?)M84[d>Z>Z[.+ZaD3dd(cA_5T^b1e<
NYW\CUb#H5KL(#5^WO0Q=&B?Fg4fGL^\eDRRQ((,>O/fQ).f38eE;CHDK]4;Z)LB
.eR4.Hb)aPG@T1V;X-LZI1/Ldg22C/Ab[GdHD2=EO-E30cB/VSS_FQW=3:c3O3-O
Sf=0<bV8J]&b[g5UD2FZ<ZHX;6^<dJHV7E5@[]QZ;4-ABYI_]VL)d@gELYTAUbL<
8Kf(>SX<.JaK-)Y?92AC9>+/W2X_DL6aO&4d(AL&SLT9HAPB=_N2(-5G]O+?4SAe
?Zd:Pe94;]@MGGNI-:6T:gaP,YD;-5b&V<T#R7?6+H2Uf24=I6@9WB&,LNRY/V>f
cgCa1^L(Z7<Y#@1U7BMF(GM]\EJ9V5;\]/GS+>G6C,(MF??LP?F@d)>d3.+DcbU)
BM[M96KB++KW45BSCT;/OfC7YJ1E-ZHGScV]#?T>R6OCVO-If>,@0(^C:d4Z\ADY
caGHdI1b<g+g>(2>5^W:TdK,G;\5O-bM@Q[2NLLDBPUG>5#,Bb>7bT]4Ha+1;H_f
:XY]<C2)U[AHU(;L_-]SNUXA.M4E<_5G@]acfOV7^B9L4WZ_IFISMGSG]\.\e-dI
PLC)0L]4A;MVc\JT^,fNb&dHG<J&]0Q-^)/>Kf&1J4^I7d_H9[V(W;V&(>WUS/fg
MV#_.CSB;[UU?6H,1a(M9R1e^adeL-2)c2VbL\0T5JRdf)[E[K9[DcX0WID>QgT[
/\D(fE9K[+I5.CYZW<=6EPbJ3X(3(-:#;4:dKb6T[0Bd&AW?-O@;^]IF]dUEO/8V
A&@D,b-d^OcN8,c/J4^/e4GQO=DW=(?Y(ReJg89,/8C53)gV^5+7>e0C/;UTe[MV
eA+YXCAd2_W&]fg5=P,dK-cJR79EZ7<B3[S+d)+HB3/2_b):IR#MG4]E+X,E.QNX
R)B.MZ_]7;762&J,7.?UF4g,0bWeDbb)7RJP.JXNOV6CQPG]..B?g.^/c(Ac\Y<@
:];[KU_=9GV9W\5HdO]J1R/<@\V\TP+fU[SM)+9GUgH#>ac&;[3eK=KZ&3fQA_-)
@#)QH25NKDTDHf=N^KCAHSOF977AD5aO-NdC<Q=?Kg+HaQFa.NW,b4GL0^_O,A(6
)Q0&IdR=W@A)XHI87O,c+J@TF.E&ND@eI-f8DJS?2(]1Pa4@LQfKF:=eZV>a,fdg
B\c&B=6c>AP[C+KA5A72TQP#E2N.?/]?8Z^]07B(56FTRLK?f(>;=+EXQ;]5gAHZ
70DR0FJ^)F)AY5CBGb.AMWeY>J6>1dAf;)_R:FQ3)1(OM\0dJJA\L(W_J215\(GK
IEYJY&]#ZSH1&NZ+VOXUR_1eQf_f\KaA2=M)N.D&E&TD@J^e0D>X?d6&44\5BgWQ
NM;MOSP3/FDC_CNK8M[DbQ?(Z&V/;;Mb=QC2M0XbV:;3@c-##SfC@N+[S+deaYZX
Q7^F?78/VHGK1b2W502^3F,^.;UF6+9-?]8Z4[S6-f=29L\+aH7Qc^HY@g(O0RAL
b>3G>5Qd+XD>R.])0,MOP0e+EO+1E,IJc1^ZZ@27Naf3COVB0JN_GQBO/&>((IRc
#2UYCH>YaIOKLb0PEHI]FW^WIP(WbRQ#a;3N8_X>d(_a+HgX2P@:71JZ8E@]LI7c
Q#X:^CFPIID@A87Hd.PMSW0cFffIXI<&8XVd3fZTb?)0LR3Hb,X6]18X/5NZYFN\
B08/MMU4&QQ/_R)K9J_2T_Jf7F(>QD.D,+_be];RU)(PZg:G4gH2<e+ACR@CAR\Q
5Y4G?HZbf)A@C6Y[I9#_B7C.S23+VBD43_L;+(F73dXNdgW9>M-(g.ZV399]-,LB
,(W^)^>SUN/AI@BeDH3[D+CCdC3&V(U\AL4:9&D@A[&b576FT.Y^5bK2ALB.XZe1
a[ZR2#KA\HN&92N+R#L4S8c/_6fKWE&&BT^UaC&)R5/VPc&):=_]C7PX;E>1IG^<
\>0[Y1g@9Mc)64F&NB/BA(:,Af>\B8a4W2TLXEHB8AY-(VaaZM,(6]W^MG?g12,a
<EAf4eaY;;PZS?FPRd9H:QK)XO.Z6,(/b;bQ>B-SV+X2f]=C319e]C8S8P<)=3@3
QO(X#TZN6Z9)4T4VaZ;B-,4b+b452WA0)>].c^\d\eV/7gJ5Q>?.db(PG[GL&<Pa
BDQJ;@dB@5-F^2JC([=@cYF64=/00M2\H>;7Af^>.,-a8F9^4:K0>PdfAbH_HEW6
dHI6R[,B1CDW,cV4@_QGD9F\b_UOR^?S<+RNFaVQ-Ld9</4D9Lb.>A3&fM+1Bf;?
[[^7/CA03/725>HT<3W/]aR4#c;GQdc,-Z-?g>Y;^fd7OI]SM3aAL[IRNd6((2M;
FXH2bUY[H1EV-)(4/#>c2Bc7)a^e#2bPcFGB+N8ZSKA>QL#N#6X56LD96RUb4>;,
4,R_FZI:L7YBT>Q<-eX:/6WGNPE.VaMWf[#E_TJ<)S1bQ,fcZZQ3U]13PRB&R^>&
KS&87ZZbOe#KBOD#H_F-f(IXU3B7)[c6F&(5/QF8G>SE_OE7/(MQ_V<4+f?W,^YQ
Z9a98+c:]@RU?@\MJMFb&384):S;G2)I2A+&46?75.W)6;=AV0)NHUTCZ_e=1,g-
UE<4T(SSO+_E_IK14,f6QON)eb.eRc>UePU,C.K05ESWSgB4RDEEC\THOc[Jd.]T
P-9Ld2TN]3J8O6WD?SW/SW^baT4U>S?9/GNR>D>.J)U^b1c\T0.[fS\R@d1#8#L]
P.B3g=PAW4WTI>,L;GK-61Z@P??6b;L^9Wd.GH6\VP/A3+&Ad_)KC0=NcQa<+;-H
bZU:M<#C<N>)A]b9a,D#::LM,(6[A0_,=L_XZNE)-X=a3Ug+7Z-bH)Ze#/8GR\CY
VeS5V.C,?\H3J8J[D,JTXX=.Z>E9LT)#VHA,2<FbN,>?^c32Eg,D-PLC:2H3>OfA
3DN+dC>=8LVbHD3DBRD/VHb_;.Da/1PW-6VR@)._UTTVe6\(g]Zc>-]g(/#g_6K\
T25QE\YCeCL27cG:bZW:,<N2Y,a))12O-<@6>A1RJ#)dU3MSTI]56OJB.PTKXc#3
3VZ1M@.4WK8U5UaH^:@7.LbF?b,Q?&:IP4_2J6Z<,O>[]-ZCcO=A4CL(3=1?2Yg9
]5>,9QT0aZWb.B(HEf70Uc#ICY22<V>9]BD4I=S8bdP<e&57Aa@]GCSU+A^AT6.<
D\D&@F/,>IJa>UQ>O+?]T6[ZXKT_.F/4)S=c)bAO2(1UZL+Z#cS&2F^G+(9_YgHM
BL;fG8@2C3P.N?g=/cB3-;9W)dJEeBeb)U^A@6+,TfC8])-<RPPN1GdNW#X>P0&e
\:_gbNR43L__Z8_3EeK&Hc6-1;;07PH&VTc8N?e+-,@fIc7(9b1cR[aaDOM596TM
cALOHc(I2;Y\BKedP#1]UZ_<2fNdb[;_X-_c>0&Q^@13JI+adWD8=#/ZK)c=cbF,
3];d0_?RSZ9IW_(G@Q+[QA_6K5=93T9D_DFI><Bd,_OM.(EH@+7GcEFM_LFCB<2a
Wa\I0;C8(,+A13,eZH[53+.THBV?c]_D/XIOK_bfJ>4IbF_,ZX15PO4aKROf;c[D
LX#B?8aPG;+N1X#8)@9UbZK36Oa.]T7c2HF#SD=L.>QRK+QPIDQWQeAc:fg@4OG.
W6DD:052TZ:S4UPOPZdN#2@G5Dg1\U/Z<MN4f(H()P^FP.GBY>T_C^\/GN@\BZV[
Y]Z6B<=bMR8aBOQQC>@.a-K1d8S)721WPAM+^aZF?SYS7(L@bK-M=?3=.M9d]W14
c&CSDC4TaTI_SYb_BEd@E7NG\A2Z_B>I)^J?JZ49KZgU8XdIY>KOI-9:(2;S4N:a
BGM5:aX(5<1CebJ44;0LCF);#LBX>U6e^(BC?CP4@@;]-QJN-L>9g13/ce,d-K<7
WJ+S.<@,8B6?V576GY#G<b)4a,Z3?N@Z+b07K2W6g.Z+@V3A_(T8XE.\EHM_]X&W
NSg^)<UYb,f?(JfT#&XM&,<Z;5OY[)EYXM0U;W6@ZaaZ+G86PVd8Zf.D(?,C0/_L
+TX-#&7^e&,82D/XAX]E><VcOQa)I_Q0=f)M&L]aN&>F8:\2bZ1.O:@+-c+4D[MY
dX5\OW=HD#2>I&aTT,&Ca>TefF)7F+:5)H/H4@[)0M2gX+]N5L+B/\b&H9M+-,.H
3-SYfN/d)<.]6&#E(5NT>DA52?9?Y/4OX-BD)A:)<&G-MadMZSZO^g#:D\=)dcdT
RP(6&VdKY-dOXLA.H#ZVd.X0LYeEgIW([65BMWgS+a8D?fOf)IJM:62^AX3&4KOG
PR6a(dP.F)J06@PL4fG4L>^^=U8eV.bDE)P&RDNT6BgO@(b2U4fS:YC0R34J8+R9
JbX8JM/?AZd>,C_X^830E-(IaeLSfRA[16<3LLdNE5?AIMLNGH)XH?.H>c9HCP/a
UQeUc(<.SUe(-(A&R^T7G94+L:U;fRQ5M/?e@06CXW?f_<9Pa^^88SPXT9;E^YK6
g.6:[@g?GJ//WY#dKXKF-MHdH&EASMSST@1ZS6FO(PKI3STF[OO]^\gEFc]&=B;/
&5WFV7L)VDgU[VFIeF3FS/08E[,PD1?&Xa3=CF((^aEAYET(@\U6M>bW]_c>#1Wg
BHZW0939/A2e/]DdIJ>M9V+UD83;JWD?Q@V_YaA]/bS+;#IA+bW;;S9&\KeFH&2@
4DJQ10K&J0f(5CEfR\G_<V>>EWAW.#@aZ)&<0#IB_[._X/S[G)3V&FT7+9/S86=I
N/)F5>>b;1^=#LDH/g+A\SFTXZQLb(;[#H.[,B0N\-C,X6ZA4?GFF-e4:aK_]c]<
(d/<.^B823N;f>3\Deg-g)F]L=SWS:(<5Uc_FBN-8&e^U&9&>7,DN;2Vc]@gP,;6
-:<PZ_6>G#?BJP25&7T(R<H3<-L5NQP2Z/8D;W&_d4CAX#3GUS7;X;#974:KZ(U#
L)1U=G?5cQEC&XaX[@2,/.ES;DJ(cF,5Gb#5K]6bUEB9]O@e0UDOEgHJFVL^_g<-
&85b4R##VRSE5C@\g5TM\>XC)KXA&C?TT.@gZf#BZU)^2GY86F<Z6EB@N0=Q^CR8
7ZX7e[=9L8+8L9G4U1-QP3=?>T9EGQCG3+_<,eWbS/fW>^T@PWUBOaeWJNbP^XGA
MIZ70g#BHb:5gJJIMb\/.<c9NL[5a6M3CWTBL=DcL66J>GeW/+@@YE;:bXeZc<d^
M,?5X0^S_#\ZgHGXV_?CHMBdV.J/FDHf[W5;0SLJ:\XO5Z;FHQbgO9788B)?gFfb
\ZcBS+BZcRNaEAFBff6KV?eCL+SUZL;cKN=K6I#NS=E)XXCY.g1Qd,QY@UXc,#Y@
;/^#B\.7bKYa@<@?cT&C<PaVeV[0661=Z(&&U&)@^:0(\D^VFc#UA1\2DEI)#EU^
:#39VM5]3J#b37cM6_BgJ\3bQDP-Te7691>CS;DM1I#[Y#.EW_a.@]\aQ^(DfI)F
YE).<Y6:WA;CN1Y]57I9N7WMA0g_IA<TN=>RN236cBJ=3U_>[)VKE)VS,d;26M^;
Y)dg)PeKQ>;>XLF6,>^:78#2d6df417VG5>d.O-adGBHNWg:C/6C7N.d=?W\c[HM
G-<<P/@Q-)5&b?,DLDV>>I5GVG1<.7-)4\WdU-Xa3<G1_cb\>ce@2H]a+NJ5>?=+
g#<MWP<XL3YY;dVSAUU&53H5e=G)Q&S\?<471A^\2f6FNJV\RMS/>b0.KZaA]]dW
f8MS[J?EODV5\Y-MPe6>B436-NI)4^VF2+42.EH;7WAHY[a?_FYWGF.LFdUC^f^D
T(9CbM2=O]A2EW<OMM8\1AMUP-Hg6QSR^#H(=bR6d^^&,Y&e)0Jd_L5/09OUeZ_V
c&(H\-]DPM?-OM:S/=6IFLY37QO\K0PgX7O6G6>?fO=fEf)-d;^b-)eA#/1FaIP?
SH0D)3(E7D]ag.Q#bDVc>A.T22/@TcZ,>ZATNW51BC,)6-W6MP])&:W0CD\Q3+W7
c+gQ/>VI^QdYH:GNTd^:O@FDX+D<8RN1a?#VK.1[OcTG5A.-^bI3;+G^ODI+\#B^
^OCC9#Saa\>6#Nc0XBWS)BIA8]cI0F+WdR(19HFd.;O:ZE.^::N:DI5C8T;L=C6R
E9N;G(gePEJGEW.)KaW9@BC[P=--V?R5/[2SH<2Xb/PeEb4NA3N5:JZ6?:SGgXG.
ZJI,H&];R+UWV7/cN_cLZ8BR.^AH,0N#Z8#NB,/ZO^M6T45+1=+68C8=IK--^LWE
&G>SDC/H(+e]I,Yaf#bO-XBM.<U@;Q(TEQ]EU.M1>49H^_Ig6_=]AAQQ:BD9D_e@
YV^Vc^c8c_6X.\NPBGALe=(Qfec#KN)4fZM;LX8g;3(2K,CZ^O7GEP+C/N6+(<bX
c?gQT8aDd>.;?&;eEO,eW1NId)Cd4=0&cFP-,]cJ_W\gGDKQIK])g&+FZ(BMJ\/+
S)[Ab:7f/_L_Yd<gEYR)Z)&W>D<AJA+RO/P<:>D_ZW8:#_(DF^TZ>992IL^7N(Y)
Kd\HB+GK.cJ-860W8O,_VSO+R23/#D_\X=S_;.L+<8DYdIG>V9O8ScUDN.^\;6M]
N7PC1\5BME[H58BX08;3:eg<4O:9gN&gN^eb)=<H^WS?cMR6)TZ>c1Ndc()AC2e&
.L],D,N.[ZRXaZfC&UPE,f+a.N=UPN,22bF@+OB92gU_bKFL3f:S&58agLE:Ng3&
77;XR6]T.K<B79=CPXM5>:A&d)&B<g8D[;CI+>YNb4G9(X=UWW(gRI=7YJ/[g)JN
-<P=^O]d.<A1fA(7IJ:QQ0NU0@SbRbW=M:DLRfG20TB#NXaAT=_SK:<\cgSd>M0(
]5Ebg9=SGJ@M1(EN;YVHP6JQUM-bFd\IF0+2MF1.)+WaTSW3.Ae@SE=[9>1GT[]-
&I5)eRS7?6E85#U(I?R0-de@a@d.O(7(dT^O(VNWZVL?J#]<G02N()CSAC(SWX6I
VW.PXcTE(3#_K88\X0Uf_P9+5RY6ZN@fLKV=,c+4+4[[VPHLda.1)cf3=__0H/(.
F3I.OSWgB8;d54IXQ&PA?>I)PU3X7[B)@]SZ[W._C6@RY<C09/#F+Q]<GU+]Z^CU
VEVE-c]&5C4>M57G<W:>A1;U4bW+e9+E8>DbIeD&[?Hd.[(M,0K8+Y@.ZXARA\Zf
69T_JNBDNC,?\<Ad2=V7Hf0QXI@&H\JH51CRbT,a=CdX5;A^?X?cZ1b6D>38\MbB
R.(ZeTL.OF:<NG6Z+7&;KOeET=P&9Ua2=KFG=]=57\#@d0b]B44Te:c^XF/=c_HS
EO_##LZJ7d80d5#0Y)YNUY9cR/2FW]T&\7.OR?WH9,D]P,<+fb]JL27;DY_8eP.N
C]S6J=),YLXKRMG(^5\OL6;J.5>U&EdP:bY3/TZT>4_8;RBF)JXGc7MYQ8X_Fa8X
YE4ZZZ5f1//-.5Sc/a99T+96:XacG<Q46N_5gg>IZeE802R-3,C,.W.B4Pf+1/Ya
/_4_=29ZD&QB<);?V.9&>0<S84,[C2+;IZLFTD\4>KU5N2\GZ3cT1<fR#]]Pg6L?
BU06E^]U6J2Q_,&QAL71MBXDXT(]KO0O3@H=Z3O0\FJ+@WS+G0L#(bF.MP2bC3L2
]A=KKg-S;=aNf1[f[8E].[[f#W0RK\+EAB5&B9/684MOHI<]F<-@-3^QC&)bV;G6
Sbe)UG9F@ff8QR)[+D-NGEVaJ4<TH]J,PU03#OOR9)&FX4_RB[.?d?U#;]>[.=dI
fN(]eeW)A\TS1e&;&_g/#9b3PQ]<(^7<.QGWcJR-A@&B#8PN3C_c><A1+UD:MBS.
O&=@1K.fBZ^#\FBGd?W(#4DdV0;A2a;X\#CT0?M&L-,&NY]O=F=PODAEDZ6eIJW#
CLHNg@<LScT0ZLT[b2+cL3Q[V4KZ?edWc((X0:LVFPWV##YOT7POg-<DN]Q0SOf4
SWG/,S#Y8&B3FC_Yb34@N+Aab\<B0-DU74BYf,H:L+fOOG3c/Vc+(+55J7a78ZRO
;MK+QHCUEP4A&C?36TTG8FV?<^7X[_fC4XS#=G4B?68\deZJO\4fMS4BS9QMW&e-
LF,+N[;G9PDYS<7AeEMg]D,,LTWfX^-@HWAJa>FP,8/46EPa54=:dW9?@9?Q.A4;
a[[D7_T/g+TR\:GBL@Saa=1FSLLc9SBR)8^V.40&LB-8B&04(HfD;g<:a#_ANMM[
gEV-?Ib+SG+N=3F)Df>d3;,=Vb\U2\4)N,(BGAXJ3+4=);7;.^2KKaS\cc#<P(K0
XZG22[^@dA,a=@eEND3U)-a&(&PEA3;TbPYc[F5.7Q<EARdN&\]<[0g1MaX\+PdO
7daPf6&ZX?B>Y-.RUQ/7)HOBbP7>X6#2Pe-g(&d+==A.>6_\]/B@G#3=OA[5]7Ye
T3)^^:4cYcW6R7f^WV^c[(E[ZbUPcZ]DFAe]A,&@&3DW1e.CJ.-2geTTT:_cR6e.
:W4X6O7&;S3B_XHN<XM@C:VX^<bICDJa->8U&6fXSH5F,UZgcLS-.:MA+bIK5?;a
MR=_@R9F,B[+(IBYc@._T4c1.3<U+cZc;X9.g<@TLAC&aNFQ/GIW?RIW19T(L&@<
F=c=PaG^3,W02+@fA>4ATBa@)(F]a+5:O44^J#cP3:^(bQ&3HX<ZTS2+2d+>JUDJ
/57,cC(g(_;efN/Y10TV9#.0Gg^KVS0>GbaMYZLPVe,2W)J-Z>A&dC?W?MTb?=J_
RM,fUGSLQ\E6^,S)GG3K?H/FRJ3Z?fV+;]GV;EK71PGUdR32C=-(F7NS,;<+5NW>
UH[deN&(:TT<H5GcLFK67)WD.>@f:cD?X40+?gFQ?eGQe&4XTP)aA>4)3f0[@V,]
K\NR.HN\L1d)Y-RQYXWD#/cQR^WYYV:QeO9SHAg),H9=+&RF56=4?XER7A]/UcQF
ffQ_=>_.[cFf.:@I_M7K@NU\4C/OB4RX=Ra_O-5&>_XO,TTMcI@H?=JZgdHM]\dW
=L41;21GHMa522L^<OEYIc.=T:_f\)),.aW,D7C4bN;#]gKS\A9dWeHQ/M=TZR@D
L+d2J9Dg\dI.^X[0MC6-1cg_;eFW??b)_[\U&695GfX8MZ/,DZ3@5Q^M/DgXMSI7
GNBd&I7A464E>6NDV0WL([EA1K2U5\+/G&>0#Y>K9#E(-49,-/+]+P>SYQ_?N=][
#]<Fea<SVJUARSVEdeOI\QS#R[W=gR,#]CD^FHIbabb75K].<EX0Ce+<-TFDBZ17
[./C6Q#]NXL&:XcAc6@^7U5&8G07)b/c+92=0d6U><_e2FVP/BcQ=RX/RN)0>R/F
,6,f9Xd]>dHXU0gWYK<aW,^=0Z<6FB3[G:[W,2F)Q?J?DBK1>37(W#61AFHG\6D+
=MV=;5;:T_+S_F.eeEY68#>HPAI.]]5P87B,C<c([PRG+R0:VVT>Y2d_WC@b1\[5
Q27GM0Q_A1T@/=]S4c0\AaC1(7gPeOB?ce[c?@>dSb31c)+c6f@.U]<^DA6@0I/1
GfU-UE:Tf+f<,H/Wg]?IC:G&\KGQA/?88D4T)cb6_d,)>N]7?0<OT4-EWH>6]3==
Zc>d(VJ6AU59f<fT<_5V-e5M<.^83e2-f4cW#_ZBD,_OBG/MgMWN]/E]18F(6@a\
FVafY=L2T0eP?U__,#N,SdX-e1@;;Q6a_H0@UBATVZU72(VGYdf:&C^/7aB)K&D[
SCLSRbFL^\JD,4RA_c&YNdCR81;CL>4D8<+g,AJ@W/_S(OKf:ggS\XZc>APcQ^;@
M,IAM=S8#QbM@S-6.APD[>D\IEc02bU93P8.4CKRTR<FF1(71#SB8J;>QP4M0>b[
CR7Y#G7T+2)X#;Ed0]]9[HJ9McLZA89O1G7R2\JRJN@1.Q,g[>:<FdHeU9LAbf[d
dHdUH;eQU@01^KLI0<;>.@&(BW)]<bV0]8RK1M5bRV8,S(G2P)#^P\A[P;Y661#J
6RNO&UgPFGVVDCB:c4T@I(CN.V4F@;H0P#KLHV#/^B33BHG>S\ZKbeGY>)F>T<3a
GKe#ISPg/]#Af]9RV)_4aSMRK[WD^4FWc3;R0BI;1U,2L:Fc3,)E2F,M6[LEb7Rc
3XP;YW+eHMD<Y/A>dC-)@EV#.L5X.ZGQ[#b:SV19A6.W2b&fR7V>N3#>0TL3O))W
HeD\\(IM3<:BY--RZd;KJ:/?W9HWc.2GVFQd.bVRGJKQJHYUC9+I=F@4IYg1^07e
#LO].&\@F1&YV(2I.Wg7PSA810M?e9[6.Q5C)USQJW/AGNAUKYfH77dAfC]O6B^M
T/VUFITL1,H-/>:5;_L0VG,@:2C6#7fX?X[VDb/7H89e-]3f&fUe9a#[;<GR6Ng1
R).WZJFYW,@=/O56fG.2X/Td+4eRLKI?[-5F3C_6P5@=[baGCJ=^P:^S;C6GB3D.
55Y3WT#F[]6-LKNR_JXHd@,H4dS_V;Rc>F)U)82?0d<3DU252bR:6NCf[&Za#9^+
e(&Z7b6O[Q?-,G];JXaf>Z;7>ZNbTLR34KV[U\T>IHd__:4TIe=gEW[1./J8CIdE
:SOA;6Y>F(57/L[TZ9B.Z1WLD9;<^aKITc[[O8a8W?ILL<Tce.MY-H1<;+,aM1Nc
B#6K?/EYB7-@+;<H:U+3LTU>3X\&<(0CW#7H6DEdX?B[[d?7[NRbGAC]A\3aeN9H
[4fcW,S\HR3U3JECA<gB)IEKIW>_8S.#3>B]9eD^(STYgF8FS/[1]8S9KN5C2=Ne
8KD,_U^K+8DGEJ^/,\#Uac^\c[0>g\36_Fe8(\>=DMM[4(L,=KGg(.U-De.G\UK1
/Kg.B6-F:;:d,P]W]/edCHIYQF0IS-@AG^]O-X4JB^5=/f8Z-#[??)Mfa4/])7ML
>aNMYG<V-gg84d>?8J_eLcS#LBaDR>\9\II;@S;#a=)@TLKNG);5Sg=VR+SPbEY<
:D53(9FG4g61F7(0S<2M.-9#,15c=PSV9#XZ4TN&V#LT)LB\R#(&.J]c.\5P\7FW
)3Q7]a3Tfg353>2YaBBO6N+G(>d9MY90B=Ka&H,8(VbJ\>0T[<.\T-ICY1UgYQ>d
O45b]0[UF6J4?70/eTgeK#P+;]#=V^]0S^:92DGLN6IMLCb6V4/\ZPO&L&(NY9A:
M?aV@:847+^/1_/c)[Z^&VU#E?4D>.>R4e63f<RLJ)90TZ[aJLL-&[gX.&UY?BH8
Qe\Ba2K85f@cTK/g]^EZ&XLY.0V)c91gb?-[B:K=D=;D#6Xdd]La--H4INP]^e+g
ULL;bDHM),Y=-J9Z/&JcOc+V.S)OS>@f>M>+fBI/Xa\(,QWQUZQH>QfgN7>F3/U-
D.:@eG/fBQTUgN./O\;WXEG41g#7NU0?KT86,,C:CKIASTP]UeJ41c\cG-G-I)7)
WF/H>&0W0c4cF12]4a[BV5#AK&X]X3;?faPce\db0##]=&5>WH[EUUTB(YXdZ0\+
&^2VJg,KTFE5NGHd^.KXU;c;^^C(4:IX=9H<C5(\+<]DedO]Kc;8)K.UD_1[SCL<
WFgR3H1U(<g,XbFc[2b1F=:2:?U[@.4g.,\cc([eTU6>O1.J;6(DTIBI#A@BN1X1
5BQV]/#b@T+>=(YF7AKPEI?MG)^^BE1@,<R,Q(X4^V:+f<86BV>1KW,E;4N\UF(f
K+J.0e3K#ORdO.C)I&9)S3/;KY.<(_PT=RZY_SbKd,b0^4(49RNY>+;:/UM#SRNI
?.FY1OF(-BKe<Qd\3XLJXDOa0;2Ob9VLJ-(f-[>_OLST_/E&&,\adM=8Ce+YZ7./
KW.8b,Q/7KWGCdVd2QB#]-13e2D=_\A1^NKCTJQ]WaDL[OWG0,5COXQIE+I<HO-;
D,.=(.gSE#G(bf_(7SOZWef9?TAQ0AV+E/NKfLO.;,+T@68(.W]P+eI47Eg5/c+H
5bBIdC&X+V/f]CG=Te,;KRXL6B52FMY(@6?732EZ;S2@]QTV]EIL[47N<&d+S7Vg
K:S/S.1VKggYGTX/_TMg<FM8BT_Id_UQ]&(>gY<ZQFGJa;C.VS1ZBg-GPLb2.6:)
=Ve4GJ9FZ=YSO73RCeVDM0JAfc0IMc5U1=bGB5Q?LT+?&+,@HM88T2I9\4?Y(,7]
)Ia8B3aeWGMN#:BPEObLB^g:<=a+A4Z2(\D-5[3)cI=;XE&<;4WMge92JQVdfL<b
EP^=FD)1BJ/dQYCaRH7DgSOBN(_/([<Kg=S>dZ^-GF5/a\D3gR=@2-ECO68JHA_Z
8/;2X]/8_>(RD.cAg>,]TBUYWcMU/Ue=27[K9>CEKI3+:[e4a>e,CJTBfMd0ZC+Q
1.D:#Kc;IKX=7309(.bQ>2+36X5V(O_X-Sc]4I;<0RNV@PQU4b5HOZ-MI.M#8IH]
L,OXBeBSfM6&9TL^^4E<1MDNXN[AQcTET)AS)XP?MfW?162Q-2;RSaUfAbM6L5d#
=-#@A)SBMANSK6ZKYZ,H;+)?=5VCM3?/BZRI[09PWN+(P5I\gP4c;UWT0E>aY@?_
W,b#3?ZV8:>EfbcEV6eWP/,V)G1H1C6S9aX#N)G(25_Z?KBCJP\<57\@?-gY-?=.
=A9GCO^BZgYXb?gJW\+O==?M0Z=0(P0U5WeHB>IGK@^S<)6/b7e.Y&dg5I9H]7:K
D(ZU@cMOcF#O:DY,FWe<C</eG2;,NX@L4FOda93=/071F(0TNM)3W\3/-,daPGF[
;VBC)]ZdggY&Xd73OaZZ>Z6CT1K\]ZJ2S7Va,I3AaK48N_WKdc))>dW?a0OPHd8d
4G5Y8\e5d+T)ef3WTJ52UeLBe/D,CY4W719_CL5eID\C[B@g7K>PG+XW:LUD6GdG
=\7RWPXQ^BG(63[&I;?M7,W4<.)8^IILQd?#]OaE2\5R,C.CCVL[;32D#YZaWLHU
(X(#gZdKU7;Lf.eI>-)bc>I7\Q\:<6M/c4gIa/US==MX;V0Y[ffO3G6U=S5e&[(Q
eTaQ&,;.Z7AXJ812\fS^<EPPD;E2H/A\.-/51S_]I=S1aZd7#g,+XA7T.#V,ZbgC
HMRIJEDH(EaHOFSSIC>FL<+RW8b)#_BP]/dXA^CBF>We=:-&^,@c<Bb[/@g:POPE
PW7R(YbN62dSBT+5C1C819\<&PJ()UV;6L2PN4?85T114FZcHS7f,_Q[YI,^GF?7
2+J@0CJP.3e\-HO,9fKOfZ]0gCdO27J_\?g:D(L1TYd@6U0^a@e:Ge/G>01,;P-B
S(C3RTZ_Pc1>&+84gK>P@cBP9@4GDD#<0=BNL68KBNX_T1><&31Vc2bW2Q2GbLOT
TOZd8MeKe)@JI(5N<T9HY98_bMeJ-6RK5:<O_BO2fZ2_8+;[=@^JAZeH5F^Y9,PD
>;(Y)2gK>/L]=4L4N9aF<><F5#L45agaD9;406Q[0e5,WdRQW6<@<A69WSI^8+P]
c>IU8EX13L;gbJUC-<,(.eM<eF.@K<Y8XIf)Y=GREPCOK]^2.4417YdG+ODg8@<3
)aeO(LMH>@SG6VZ6?F5<77g-I(]5F7V:ggC=^9VA4GX02:V+Q0AQUE-Z;^AV>:A#
Ab6,)AcR]2(/^7QC?)W_^W&7&^/58[/IOSY_#W/<1dVWR]a()Yc#@<H\a6FNAcAO
1bQSdbaLC];)[Y?6gS#U3cY^cf/RW+]_T8T&U8-4LYfA5U]5,:K2dIQP#4:#<<V5
_dKSD]LdFfVJH4L7a_>=+B>7T/VEd-5L+.fIaW/RXZg^:GU:#?5,;3,gU/H?EN>F
HA,/X/I4PGS+Wb4-<I5d(f5=N;L+[LO+O<65E<9Y.)b5YLSBcZ-S;9Re963(Q(3N
5Ve<SNO]SB@g@)N:Y7BYO,R6Qe6++R_FM0[9Y0XPA?6Qf45+.MRCXQ=7YAC/T28[
aAI8?+;A8E<VJ)&=3_#+-:U2)3WBD5HZUFA8CK[K./G[0Nf8#E+B:L0-1@9+d>DR
3d<\:SecUOcK?71LIS4]2^V,#QZ42\fM)7T78<ZSb=+OD#@)Y@46?(I.)LNUGe=,
):g&S-^c>e:EQ#EQ\LR+ND9g^)e#^_Eg5cM@66(+8JSdN_18bKA.MC6,C.PbN3[:
@;[&-3fLJ@BGS32eZ\CT&FIPF#NEe:ZL\J^1gT:F6J#2;^;VXC2\)#0a)SRON,.]
gU[LX:DZB^SZaXQcP5E0UEHCe#D^d<c-a^A,aI;??4Uf6]4(:ZQ=49SLc)HQFfM>
L4<S@FLSTc(F==.YDNac/eb&]Yg7(ND#\>F?#_A#GXAeY-2)5Be>-E7K-S7JA&9.
#?ILa]A/b92e0/-:=].F6bL5+V+.GIUed;X?RJZ&(XFQ3fV9@=-FL79K[2=L;&Pd
ACId-JTO;KYQXU+38&0(GI7K1QK8H4_OM5W::77S+[c2,IBbEB<fN=INY&MPcBHH
SR1_U_ZQ3J4Y6cS>X#R[0^A/A.^g)A^cU-7;O^cSN&UIW0^8@M3Fe?>;^>LaK(\E
(R_J)I#,ZKDaKH05XIceE&C<2&#:\ZZQeF13&L3Z86T)Y(S.6T_57aC^cR6?-.Qd
YH:PM<BHG7P>SJTMcba(Fg;:)M\OU:-cEVNHJa]>RP/GPRa\^UY;==3W44,V4&E,
,-c5gR?1H_,(<XF1(D?eeS/GCf].R/221LO:SZ<JEbC+@19KNWIUg;0;5cf\_?2?
PO95F6<:2Z;Q4S<FLHJ;);EV@&-EaB</#K8b7d?Tb)g0&&D5X9;;I&^a6@NX<fd9
B@DC])+C#^300A9#8P4/M]HS#Z(FBg23PX5:X9@0,B]I/a6Z&NLB&?I?2E]]H_&H
[1.Z/)[d2/I79R<Kc<0TA@TJ3f#-/BbDd5WC;;?V62\Sb#I].Gb@1QPf^Qb/DHD@
ASR8Xb^@SADSb,Ve#<K(5.JJb7^N6V[]1:T^DY\_g[</3D\(6H>(BFN[e&AS2+Xg
TW-W#C0+C1D\)F7;c/^US6,DW8>(A:dK8TMQb<e[.d3&d03Td;^)ETMc[U/TK_AP
PDT_WA/K+SaDdQ1;)R9Oa>-T5e]ZQ<X[0Z>9(bV(:M[#]OeG/bK1E3^b[Y)+BT#P
(IOH9D.OXN_320K/Q30@3^=e94JK,@@G.NHd.W1(-ZeB9_LTHE1dVY+@ID8gGF>N
&Z8b-?&dP&@O<FKO7=U740^8KA?L-I_LG(f1[0GOFPg-L=>21^&H0-61[c][M,aF
8OCL6K.,FR0)-PXL/ceJ&[(?Q3eK1W:2C85gCU8&BOLD3d,5[X/e-M?,K35]0d#c
W&<P@?05Q2<@I+F9\0&AE]S-IST0UQ:6,31D?=\_a9I37QA;\XH9)]7#:cLV\0Y[
BagMR&_?^B=CA4<&PG_ZF/6[.F^DLK67<.VL<=MSffK40:_Ca@FdLU##/W51YV_F
L=.aW/L>Q4KL]<C#Q#.0KH-Q-?]/8]4U.=AL?HT\,7X4b4.QIba0NaWK/?/Ka#5]
DJX.:@gd/>.)#^IdL\<JFDK1?+/?9^+)IXQMU>6@.eQVaUG59DaG]Z@]A>E-4FZF
]1>e-@?ScS(1>F[1H[]B\Z2TW6Q(,Rb3>MWK1I+,c7fP3F?gD@>,/^NR>7C\46L.
5ZSN:SSQMLME#Cf==N/UM>)VU9MX7H_][:6I,JT1SL,B5/SR))H8&TJ2MVLFe0SW
Y6V)M2Dc#YU&0N6__&O-TaA-T2F/@ccLgM?_0V?B-AX>SCd0aD&/S,[.9W)4RY(I
B\6XgAA=IH=@^FCH/]EVe9e^8C.[IAe_b&;Q@A<RYS3^8DI#^K-=K4@H;_RZRSDe
5Q7NH_\94G.E@=?]VMY&Y=0R?@&;3J&7G@X&5M8#A9M>;;)^>FIU#D]#7[(?S9MM
]P>(MA=bQ=3AO<<TZRC[Hd0<ZJ71+bL@KBYWJa6G0a6C4Gf,X7YeSKY4,7.F&Q9d
^#G2+Vdc/DH,YBJ5VR035X:C^X--G;&&6F#]aN#7N0V1VK.bF>P#?AfX]>9VUJg\
N4CY_I(>\Y_5ETC2IGG=QY5Cb=NY4OI^S/;HEXaf7L];?I9+EG::FWG6RB8[@eEY
KWfZ<OO&6767&S7<7?73U]gg3O5_Y^>=R4R8]U553ccaR[T@b=+Ga^H4H1cX4LPF
Fc(FI73[NAR21[J@dF+I=7[D5ZTbLWY)HcK_4V?SO34@a-W3<=4-J1cd450M#L9)
>5FCDHHO<f5MSQAIAB@9CVA/NeQX)UF];/4-_OY9:M=#K@R6H9_.E]2VYL@KNO_R
(979P<@BG;Be#RM=UY)-TF^PUQbZ5ZSM2-8A<F>b0]c]5,FagF0@N--MG:=Wfc5O
7E&=+fGTL+2&/dQOc^TZdB.93(Qg3WKKZ)aN?d07WfNVZd^J3Id,E3F;T1N9THdS
E]g/MG&.?GUWU8SFNO?dd52,^;Kbg?[bEZ6:)cPH(4J.ZWL=eTO]5ZG>CHWSa?3?
f]1V2-beJ0^#V&g>LK^^[gNM<\1V/H/\bD8f7LXT#J;+QH71+?OZ4;EN][J^B;@R
2VQ6@J[W.S:;J5CD+7TRe=?8#)2ZPRGB+QSe\[RLYE<ALX@><D3(]@)VagFY-Rc:
VY.gb8>1<,P&acY,YAYET[(ULX6N</013R^d8a>J/6dLOYdd7=Q@;D\c[H@5f3-9
15F^JY;Ae?WMeF=&;5C=;_H-G&U2MdKSFAd._4J>7gIZ?.]BI;U2+^)9V++Jb=EQ
(2Z#N?2YGQdQbS2YE>KCb(RH#aS7G]+7f_.M#W8)dV7TYe1(_+U3bZ)R?V8+Y)dP
d&5AC_)YL7I(fHET29,)R\b/7M=Sd=-SQO8>7OZ&b\9UD8I>JZg^Rf?5ROBW@7L.
Qeg1a.95>HUeN1-^K^>R/Q8OF=:BE2BU:JeQR][WAD;M<e3>-eLNP<fM.X77e47f
?=H-48_EaA&2f@d+),(U9Ie4CL=+U[=4Q6P2Ea:KN^\\B9<>A/G=HN_QLd\5;c6#
TX58M?01HM.6gc_PV.=4g1@_FKN)<Z\6AKJBT7?0Qe4;SR7JNeAD9NC=\SRJ;6GB
(L\J0cS8\Aa.VPX6Q437c4HW,<\AERUPK./BdE&5];GFHNc?dU9@WABg)bdT4\DP
V;-;L36#<ZF1-[S0<E_d@.ba=/I@Q9?5GH_5D-Rd#=Z^+6A\L@1N^/2HGAA.?J+G
#(,@Q;:9MKTPccN\+EX@cSFS+e9;J&4Ie6_?S&=>N8QNT@F\GN_fXN5A#)&9RJF^
=3GDI3D+J7,/<T-6AEL9N5G3XP08c^1BEKM1##1D=W;-SKKT.SdBZ=K-UEbY0]fQ
4M9>-6/2SU.52G/C[Q/F;7?Z:bC_V]Y806XI?]:J.KaM.A5UQ,0d#Q9-,LV;(DQR
8\F]P;aWF<XQIB)D435Q841Mf@;&bcSRY=91K#-,Y2M/2UWA,e2=/@fNeZL.D:1f
:;M^\STb3\[.H;L0_6IR9L+1eL<PX):^:A@2g_HP9a#PE/c-5R,(96C8OT)3ZQ3\
K2]Rb4UA)4HWB2a-@d5Z[UUb@J>1E7M6E47O.TMEMZD\(Qa/U=8G4F&+)F4&83>e
PE@POcKEb6(.gP<WUdLTW3J(D3KFW)+N2(9.[H=.L@WX;VN4;R7O4[\@W+ZB-3]P
g98A>]UCR:5DV#_e0M^>Q(d,;8_6[#e&&S+M=Ya6RaT(deXa60WKY91//^GT#W98
IC;A/J;D?6eDS1>7P)#11HWL:,-UP^W#OYP\#4eWb<b_:30<SRI5#N5e5(:a[K==
@O4;#[B.gB_V:72/CKKV8:]I?N]W)dI.8U=KR1QVY>6^PIE+>/8^G_GA#XH12DOZ
G-ZJe:DaNYJ,fZ41A(=2893M_A<FUO=J?]8TD(^c+Z0a16Z[_G#Ve;H:02C]33;J
bY1:cd\HdCL>YdY&LGI\>1MQT3b.]KVG@7c[8UKSEbM:GE]JWFD0ZO]ATG-GV/a+
Hf>)Cf/),aL(V>^WLdW(91((N#]4>O:e::-BH(.2C6Z2-V@.-:EN:SO8S8OG_5][
Jc7#(P6<G>J5fd^OOY4>J2[9L/@4;UH]+:+E#?1<&FD]3P(N\SM.[O>^8#SC<PEQ
cfbY,SVgB6U6\L^W>bB332)g_HC-c_3N5:6B7BH9dX>f:RE0<?eCNZ0C@VM\AeWE
LMRO=C:(B#&HA=-)G;(@dT]+-2P7::Gg,0REO[.;#5baQE?(HH)K-\OG].Q<FT,I
K8Od:gNQ87b>a=MF\OA6b6.geK]R=T]?,6Y0##(9I.1b6/0@.1?b48Z^a;CLWM0)
,f<Oa9^(g[C[g7^X>E4Q3G/<GHQMO9[,YJU?4\D.O)MacC.M?O]Q,CffE/DG/VU)
.dAY_1becaJ2aOXF(FC>5(ZFD0X72eIK6A/&ZFfB2JO:398U^/=&(0\[M_0\M-,g
_f9S1B4/&T8F]b=>JGg-6#=Y3#,b&FLCC7G,(AEd6.H+@DQVNSd[e6A[eDZS;eH+
;T5_1N]1PCEF:5GEb>6O]WA@1+:PITY89EGBe/,_R[5<9@(7P?>JQ>TLP1)>[?3)
f3Z;ZOLaT0G?OZ5R(73O6?/34W_CY:]g.-J2;<cc0OM@)C4N#;OYH?<>cQ5&E_ZL
\.GMg#2OST-\=e1CR+G<#=7JH&D,/dBP<Z-]IRe+=NB_8F+[IE9fW,7eEMgTF9?5
?]YF&201Y@dI8&=YI\:1:9J;^?K2K:690Bc7.^)aD5XaH(Y>[;7Pc71bW?T2@7AA
L[IRRCQ,D00J,Ha88SK5SS,,U;c6F5^\X>9efaWfRP8+46AAX:>M&O6VSHSYODd+
1).P?E@GZb#PE9a>T;++a_a9#]QW(ILN1d4L;[M^Zfa3d>K;JS/.^a<gf;QQb1K2
.F,2TI<67fZW7V,=JL4WdLc3a^5I4T7bU7ZRb2Lg6B&^[R+].VAG[QU9\+BUO#E<
L0<0[,2[UQ.-]W2#QScM#5IA575NgY?HIfFSQS2Y;V2=V6:5<fLJ^E,b+MHA^DUZ
f79A72O189WZZ_(7a3H-[@1,]LfFZ:+BBAN4U#L/,dA1Q#K[Mb,gG>(J,_Z73H<X
>Ie_1J-:3P/M.;/9<6XE18gO51:?SCgW#-Qb7Q8\e@aaG@cPPV]<@gNZJ0IQ<Q?a
H@]0G<;(cS_:JOM.1-J(_D>8/degH0L9+4:YM:(,_:_HLH#?cFR8D[cc:f8+W[OD
\W=^,?d#d[f4d]=YF8f)RNYO2a#YZ8<gY#4[W-^>Z]/Jf=L_&[8[:)Y3AM]@D;A^
1dYK2N:HT<PYV9@SdeFB.NaXR(Yf?3:PKREP4ZCUXSJ199758G(&g9A^4&.fY=;W
I;d2g3NI&EA7=EP@A&MY&OYbPC(JdCg7gaQ?:1g[19Q-TV>g:bA.IC8.bMSYG]eV
)#e13Ad<R+.,^N+a:49.gXMJ)bREOB<Bd.T,&.Xd9G;J(ZWBE9?-)L]L+_C3bf53
98Wb?^SO2@E)6b)f9CH5AU[TVH::<^aPRB+3BXHdV3@agP4TG)d@L#WK[>OUJ6N7
FH4GBP#I)eW07?=>:]e<0S.9PW]]QX^bKa@P,K0f&1N\d.TaG.;]aWX^;N3&b#C_
2D/S(-:H-373J9-7&H(AK^cQJ;?>E\R:Jb6X4OFKf127-RZb>1Z=GUUH9;MQSPbN
6B5E[9;#N>@&#Y@<..82.>EbK&1(&b9-@-,Ba4.fW[J-K^DP#0e/:_eE:.8#MO0=
a(T/KE_<\3RP)CLM(JC>X?Na0VLDEQ,D<CLfVF</\5/Eg?3X>5J?L7./AE^3Bg?^
C>V(RbJ)EcO&8INQSA7=0TE6>\4IH#IO4I/#\Kd,ZOC\_(L=c@6[8D>8D_E0.5+J
eg:K[VV335E<ceWOCWK#]X5M0Mb,AY/-JC&4,FLa3Q,,7/,.Gb2;2MZ\R>3?b8S=
89FJgg-X^#D_4.AQ@K[>LeWfOd4Q,Ac?#KK08Z/[?(g=\H<\@+F@,&K?H&8:QS\<
gXNM_f6cE+#Pd^J8BQ1C.-:bSKA1ZK-a<[Q@AaDP8cV<a+?a>Y4,T<N6#ILHg?F(
4ENgZCHK2YI^L3O>-/^;4Oc,0TXISe7,WE-Ua2ATg\>C7]GZG:3YUMLWOW9\W_7;
>/b.+:KT>a_QRF[>9eL>\V68^MgZMNPPZ^B__)X:c0W^IE/JA4:VQfK52d8FI6Db
;DKF/9A10X1I,E2/^fb)Bg+cS=U[W</.U5YW0@Z#T.b]-bG:g<6#477UE],>_=]Y
WEDH9?Z::1,_3^R04<QQ&=KTTRC>I:?e;)E<0d1U@[<N1A_G#fDOG[;BcWE9KOeV
8;^?g,E^I0#c[WPJ2+,\1Y.Qc3NH^@M#B0Q^#75J879X2UX8U+KF8H_D(LeF;ZL2
@5T@F^IKZd]g/;T]/9ObNMF-#88R[_:,5/_YcdRHP-)E3\UYOE.3&Mg;G(G3/FY<
Z<;)X^8UY]QPG9S[fY)L;WQg&e\gR?V]^2<I.8_Te?@1TPO[)YIOWAc_V42EY.+8
MLeN;G2b<]UP,IAUE4>DUHD]>WKJ;XDLUW;-bE#F4gRYZ^5DGgVYd\f)[WK+-+/a
;60/G;L22X/eM++I+N-HG:fc=B;H=)^b>:BMA9LgcM=MJ);)VU>(_#;[ZWI\(dRV
<VQ-_X:I5_BJ#XRSA)1Q[^^<N=eeW;]YOM,cJQfW=_F-@4:=;@HUHCBL6ggD&6<L
c@)U0<,fB+gb]Y#26;CI3#P+gS>KQ_]EQ0>DLZ1DP;WDH]cD8(=6DGaQ/(R9:LYK
V2FQ]:]NC;R==32]bJ9^=D<M@c0@_16:DV@.BTEYVG===HRVBaUF)9C]QN/f2&11
1\a2<MQbd3469:B(6H,d2W2X.@CJBH/M+-&#0JQ=QQ13-c1:B)g&fZ_AaYc+dQNS
>PaNACFaH+>ZR0W;CD73fYQ#d4fL&TP8]8.40QdG8>#1OTTK6)01L+3O^B5]g?J]
FAa6NAK]W+@^2cSD+XKJZNZ+>DZ_@&U-47E^QN3Bdf05^:ZOZQa<\dMFY;4;7Z,8
01-W)=CV:&\Y-T_\\C_QY.U[-dG@M[6@QHSP3X@2TB&KHbYDRaO0K9]b#a]>K#51
O<MXb<J87091+cT^F8Xc62W.fG9d@9L];=R5Rb#JJR]3cZA,CZ0KE.:-[9>:TR:+
5[bUA0]@HO2d&L=U&8a[[0VEBTT64fd^H=7>LMOdFXIJHK>[)3Wf@240)<Be@3b,
]e?QU=9X,(MIQ(dg#@/4ObVB9IXT,1E^(0ObO],)gP[(PQ286a=NcS3?USX]6N_M
KVf>]0AVe\L_M(:dWV&dV5G@Z]HQ83PB\@Y]2;<+NGAK_;A88XKBW6CZT(9XGdSd
d5;a/Ja2.M7DZ]BO0X[^;KdZJ27gf,C9]Yaf3P[8;DLX&C)PRBXUQO-()75<9-<Z
)@6HV9]a5S4IHMQf1/YGZZVE2<FYKYF7MEd7O?9Q6A-g9SM]FCC794^Oc?_f/7@X
=8249PeB3MD_6C)/>2+ZTd3Z7_VX>8^2+cWc/DZBK=IXF[8XB=XSU_:\R&^;1<GB
5>6V+Xa:aCg@;:@E-&+@K2(X1NKK.eVDH6TIB)(;2:2WR26f+/FQ]a[#=R<aNTUE
OO.QLcJbe)\B7e+K6Mg6QD?49aQA-,bB_J7e;,^<L:X&<YKND=9PdH,2O>127F;\
E1\AHa\KBg8;B=Y3gV&JY/YQgZdTVAFVOG#0@YUMB7&C2JO7I.Ae1d95<-814OL.
T3P&-:/cM(F]dBOAKg1PM+KNG=-f[2\=>XC=&JV3Z0YO#2B#G-,)ggO<c>2E8Zd;
]]#58_d<8a1RY1b)C^;+1^173BT^9+HYM?<]8;RS2>9;bIPJP19>c&<N(H)M#;LG
GP.C&)GF.IMbP92&Wf@Rf4K>N4Q[#Q:eHe,,d7<fVW1RY_T@3?,_K\=85PDM^W;5
&5(WRZd#/]?gK/dcRER/1DYI6JbZZ\8&?^ARLB&OCbeHY:>\H.8;/\T:6d7=3R3(
0.UDN7Z?a>-P03dU@72PG2#:+AYN7gKaf_6aBB)d.7CSH[FV7cG=MM:BXK?^,=^=
&2+Z,(;#,8/;PWS?U+4[c1,CD66N#,>D:bd&ML8#3-TbG4MRa)N5=_)S82HK@5\W
f6c/gS0VT^I>cX/9fYf:,DJWQZaVHD;E2f?N.MOe)]#ABJU>/5M2fROAE4^.&d.7
BUa#JGfEg;A;?VOP)cZT0ZX\<dTXb)2^CO#AQeYTF=6_M\e]#1+d\H(fJMT;X^RF
RI,]NOM3^+G>\ZPFgPPbYK>2H?gBOfBG@B<M#]9cC9Nd6U.#1,O+:V57Ge7)L4,d
OC&988S\gg;\X)?>+6@:TX9^6KB?>IebM>.0dK308P7[bg6?ca[IFW29BJN@Da^W
c1.<C8fYU[YLW+A4_eWU1IZD4ENB.6V1N^F,(5/7]8b1d07]HI9:HR5]2GL>f?0Y
ZZVXOO7eD+,A6US3B=8A:?I?=:?Ve+3EP:P-@K(P-#<eP\>D@bS4^g\1[4,W8_?@
7G5V8CUf:4#ARL\1_L(#bK6TEg3(W3KR,RObR5Y;<[JK5[,bQJ1<Oe.QTCU<=.1/
:X+]W.;U4&_?8VcRA2a?=G7ZQga\c<(^MLW^?dSX0LW(5:=0A@g5a>\SbB^#V.M&
Y2W[#NFCLeO\9H@L#9K09R/[c8EPS0OOL6^<U-H4a?#7_E.0[56;gg_V5bWY/Q6H
/U@Fac1XF]+dOd&^J3]HG-QBS/4Q8UMD@]H>JW4gK/?/YQO3I.GE#V#SNWVN)=I[
5:/Qfg,G;@A(]d>59/b3TGP]HJJ[IL/L57T)?bXgA_Y8f<;K<dc>#K[X8ZEXVW#N
d@7.1,S3deZ3eS8K\8EGc?SgOSOA/HP;<ePX&FKL=<;cA(S8PC2O-/DE5OdY2eJ=
]/G;@DH=--14V4>-1b2&@;>UJccgGb:<EB12-ZX7PLB[=^B?E>9&J3RCUbE.LaKH
Ra(WcG6#9ERWeNca0^?ZIG+U?V?C<0SNc;cREF5cdPI8E1aER5c>3OW-O6=P?+3H
ER6U4dYAeJ.XOVOB0V@8,/BAQ-X.cHAF/7[Z1X3C5OM0U,Q_._G5+?T:KVA/HKZS
fF@-J].=-8L:Z(=WI1aTb-F9_D7_.B,L7EbVX]E<K_0&[9\be&9VGAXX]__Y5IY6
7-d)d](aN]ce.5V1Ud>V^3M(=M2^#P.^7\7Sg&G+,?52N9N(b>W.N=_JE(L<a-4K
R7eAEXL,3Zd8B@QHO<cS3EZSGg,:#PG8=[AT>)c69L9O=BE:6TX71TNKf.SQWBP>
9(6JC3R2&cW9fee2LSc10FCH/KcIGZGe6fH+?eZUW91A&XLA@_P^GOUW[+UfGW_6
:\O7dNfZHad+[,B<QbB7,N)>@]M\>#:]]HW87e@WB81[1+;>Lfaee0Y,dTg^f@2L
@Ldag8&:#R:KNO8@L<9DJKKF>aF1D0J\Nb/YK&4.(GcF7&_-EBG?>6f<e=d7\I?:
SS5B.\O<]FGC3.2Nf9UdSc1)g[Z+P+XK.SU06.8TGX)==,eW#(Fa>A3I[4eAaL2-
5R_H=@_D06[DEcff5IN_M8]I?].NL.eSY3)CKHf+68J+N@\L+(DBLSYYI5]P^L.A
75K.cfDUJ,6gN8BL;TJg?O2;F#F\?&8H_1XVZMH?]8Q0I<PMbIY-DE0aXGf-/@9Z
&=1bc.WN;gG<R-F(_fD6FJO]2+=JP:<2DdP78PXa,4?@,6(?(C6<F8<JV\WQODBQ
V(TbIT;8Q3,=+>SGg3>\,&4Ya>05f>@;^&/c-;,9?a>0&Q5J#cc)IBXbQSW5ZAB0
=b)UTVVY<6XIALJY(62Xc@DQ6a;1)H+9;_-DBD7?cS^?+aT;X6D?KeNFPRUN;ARc
Y=DOgJX=6[4N5ef2dWcXD;I>N8.Lc@YTYFQX:_CDM-HNO^M>PXW/U+MZ+d2.P/YI
,D>JGH_L:f^)-R_S2H#L2>MH[Ic?T/5fea?A,J@)Sf-agfIQb6N1_;^O0S.#6AAd
0DRTTW.9))DF#=HQ_gTB#@(5#TJ&XJ;2d:0BPIcZ;)W<R)6[eHF_2E:R:T+[4/0M
\Q+K\b_?bDa>-#TfH\]d-Q[aD;&d&6WMA[2@^?_6cZJV\>QZR6O@GI9T-SV#e7MV
6.::71I+e:7KZ?9X#/SR7Ed[ND+Q&U?KN37e.I[M(@N^]5MdMT3.7]Ab,Ra5P(3c
F/6?&^GK@OO0KS<9ELMK2WN/JS,4/[LMU^PA3JG0R=2Df3PWCU8K?V6<0R9&eK.(
W;JVSa_A]],3S--7+O26&QM[81UcXK^)OTUU->#Gf@b_,85K:KgV<P:2FM[aW5-g
Vdg#:R:8aX0Q6V>1Xd0WFNX=\0[]H[7BM8FZSLXF9H2@#>f22([T=C#XI?<PXCG9
X@BN9\RZWZ.VPYW/fZ\:b6)&9Id?OC<Z_g@KK2?6cdI)6;V.5)[CMaGEZ-,fb^Gb
8L+\R6^UbA#LBJD1]MG2>9dY+_:JUOWCCQ.SEYMWL[-4>5D6Ae7LFO3VdHIgZ25#
G.2BB5e/;?RfFBJ[]\f>-6GE]NTHe@PCC4Nf7K>P6TE:?f&]T+1=SB@+<7b4[08V
>:H-N?NH@=YbHE?Y=Ab@&SBPg4X\Vd^JMfI7&Ge2:\OgZN7-,QCJFQ(4E#++dJCK
=KWf[dE,O>&>2/I)<(#Ce+B[FX2IU:(bO(=;_B(@F:JgW&g3(\f60PgZ5R29T(ZZ
;_=W_EF]A[./^EGPAcM+S4&I38#KB1-U8YbWY,I>F&>=B7)Jg_Z./TE5Z^T-[L,(
)aV+YMb>=<4UeD1L)G0KZU\J>SA@PC4E&4YR=3>I-\1DOEJA]_I.J8<d6^:c_3;7
+M(I[&=?C&Zd,aF#E=^O,&A>/4ZZ>/F>eHWXR>/?Q6\)7^aY0/EeNHI0Q(0;GP2/
+9f]AZK<L\&:<V,9NML6M)>QWB&5@1=T2659OB1V-T.\\[YJPLK]&K1EA<3N1c.6
Y>&3a^D(/>fe?.,66VLd/=b8NF\.EB4Y(4WNL1>?=PFBL]G&UET>CGcg.UAY0eU+
dDEc@KA&&H3b<[feQ\KASaaA:+Ze)S^YOV&UZagGOB9O:#Y#7C5^9.3;HJRO9R7_
:Le17TQ:O5b/].VWc/VG9U5b29UU58Z@4Y597R(b/4+?VEbdg&Bd7S2J/dWTKc+2
<6)9af#(G;2V,;Z#E;43+4RRdcLDA:)#/QE?2B0JfA/V/T(.TJDf#8.:4Db@PNH=
NLc>7<3.4#30dI>GS[B4Z9Ke0VfDDVU<,71?K_-8?5OHUC;N.2SV]5^bX@RIU52]
Y_;1,<::/.f(?3X+fgGI[=ZFgTcTfID97UMHaV_f=G32fBbWP<eS0(\J^GJPPJVI
37Wc\J@<92;Le@+D@565:#U>Y+UQZ0#=U1M[g/5c:BUQ]JXTgDcZCODFO2J_>NK>
3-Wd8[YT83[XBfT@1Vb_]XW9ZYZ+JfN#@#2=8aYY->^[Q[#0KIQM<XHeN?&<:+)1
:P(2=aYF7-P;X+Z)HG67&>DTf]IgPf73B@A,L?&WdKI9gDVa,cV4_fJR2ZLcJL#)
]J8_F_491+=5eY/(E=;9[e0d:C)7FB?I[UZ(1E63E\T;V][3Q9:UU?^&M1P<.bY3
#/QV):#g\[@d<TZ)Gb?7d,O^>MUX,;=<=@^d#D7J>7B:b1g(Ug;X5AcX2.LG(5Hg
UJ>(IS^U6X?OcaG/7cX8;f64NH]OX28>;^79_PT=(-\C.C:?1L82Q+:PH3G[#LFP
gU12YVCKT7D>QF3.V9LK<#(WMf,FaS1W8JL?@E:^UNFWeVZ=9eJb6MN8;_NebRI8
UB-6Q7d6OT1Z1=>;L_Q?&a#5[XODVf5/O+]@KL/.;L\P;8e?1F6,#(b:D-.97OW<
;eQbKG3f/RI7;4T.4U=YA6K/-6\)D+BH=.:,FM8(>F:=TF)ff97J=dac)-gB\[WS
WbP/,TC65_[XJY,-@WH8]C_@e)JU<?B[.,LI@TCF\J@107D]FRU=VX(GCZ5#RPU+
d&0Q)6>TJ<HM3E6@;\:QIS9eIY3+<R_Y>c:bT:XQ\WY0ELN#+A^WWJeePd)X>e_d
ENJN.e3U-[123OKCG(I3V2DMb.-9+6[&JYGe+NM__:R:>6WSF+4+[DFGe>&>>@?A
.2/31Fc?\KSZVSJAZS9I7I:a@@ZBB9cb/GgTT[B)63AIbXLT50Tg(I/GYbK?D[_&
>;_QdJF;MN.f5cXMdII?SZc33;f9bL#M#S9Y\5D>MRNXPB;=VJc1KOe1)ZLG\SPV
UK#gO+M(A,.13)fEW.UMf=5eA?3BFGI<9]#,F_>)e5QAc?&+g_P^+4]QA_H\6EML
DTAgW\ac\3^5E^6H.9CYZKF5=IR6&L-0+Y,Sff_\_@cJe5P9/,6&Y8E.48(F#9IF
XeJKa=I;eacf.(1HJ0c)#F+KLII@MDNCeb#e8V-_?5[T6ML67BSc4BReOa9_O8Mf
,HWB4^eWU8+H[dDS6JJBgU<1Z=cf4V8DL&@.U+LQ&INY2+2A\BQG\=^I6-J<YV>V
,TEDKe:F0TEKaIQ09_&#)P@&Q9K,M981aL;IbYW39)Z^#&eU+C;J9-OX9T9dJP5F
=?@4Q+ACY/&/#/8I,M/L2&RR(8Y_-ebFgZA(0SY;.:3^.LQ-c1P7=C.?;G>6Z]FI
Dc^9&QV[?f[OZ@8Ye=O8_dM-N^-E(6R8a,.6gDQ0&<N>-g>HEKVXUK><P?P&;6aO
W6NLHT-M85I2+5bWa3Y)L-Y(HaM3E,O1^G&V]g_;ON14H^g<OI(K0LfS&R#I_Ib(
H:T-^/-SMPIT9.O::7)LU0Wc_f<TMA6K<SY(Z7;If+2WbgaHg7JF]Q193QQ#cBNX
:b@M?;#f6SCRFfH-@c]G-)^+8GB-V<>M)=<;TK52WT=1M08XL@C0XQ(FC3bd-0<[
fd6^2dcF-eBZLL6N(VYA5gSbO)_12M?3/O=^UYdSe:[&-g[ZGY3WHF)NQYB1CBbT
UI4\M:7N_GNaN>S8ea^:9)A7RBSTc6\[b_Z<gQX20WV[U0K]aFXT,dZ(ITZFMF/4
Z_?T3;CABc6Sg;<A545#Q^QP;B#e]3\I4_8McW3_3IeQM?=(=aFM?8&8[5ff9B63
UZD;7)@@F2\GBBY-.IR7dOG^VL-H?<H[P.Rg-OXe-:eZ1]MCD>bFH,)[N2SH3N^]
_F.P4#XV,A8D-)K]U/R/De^U:TOP\F^DebYJHSJ[T(+UHNXP(cDRP/X8ZKF,YL;+
595FP60KRHP(8Z0P&[&<QW(CU3egF<CD-HW>9c5\f)SHa0;d^;09MLJd4>.f.(WO
:83GD;<)@<<WUJX4Oc7+?\KQO#UQC]7dW@=DVbVZJY3e8V_Bb5ACNFgQV5X]:)\;
@gaZA@HbIN)>0>6XNC5BLRGbJ5AQ.JHd2.;T8GQcQW.9X[/WW;/9119&]/?L#I9R
5++;KRH]QUSQ-W[G58[YU7=_6H7JHeY2(23[@B>F.<6gYIIc&eQM<&=/)>/1.WG0
[C(&P(7[R;#Xf>gcSY7CMH]]F^G[#bU-<-#d?Ff2EBc(]ZfRS/;?BY6c:Sc#f>[]
R28>O5A<KXXN:OUI+0S_1C2&?=MH<cE6H3E^\bbWN(c?K<S87\dLgH\d/ac\>V+1
QQB4(Of>;>K7bf:V(eY;,]URY(:T&cHHCe&E=ARSHCKU2#c@(,YOJf(5^MI0EZG-
QH#\9.634OS_A4degeY99:#Ye^S(3KK8Zf>FL860(#8.DC&8-LR,?@(^e_?,_Q8N
fe[7,>-LI4VS5NZG^G;P?;Zb\\I2JQ^LTU3PH;T:&f#bJYUB-LGICH(O+=M&aQXc
&GE#2#8=fd@2f&P3#21>WJ&S<A#G=VZARK]1GOPO6<fIIG)UQOg/YEc5S35PHe6R
FV2[WETU<YJZRRJJfOOE)Q?W<OPNB<R]0FK9J@=a@Y^Ca=7=AMLg?Ad;L@K##FL6
C;LZ33LJ.(a&I]1[QT1)&+7G>6dHfQcM\U#.@]NR\f8EE@8.J=^Ic6,EdEd]8BNM
:[5>NZab88&9N<5#_)Fg@N][aZ6(:/AZ\:cHF6</)4[O&ecMJF/7@Z1Rb1-W5&HW
YSTB_^_5e<L=g@:0eF:KQPdcRMQ,#7GI@EWA7HgU()D@,Pe0H0:.]S[,f#.;/C1&
OX@-C\?dH[+B3b;^XNOGJ]7+AU].#-f5UI2M[R1GKYA.0d,?Y>&@d5c-GR_7?(C:
O[V>c__[X57O)A.ROY?0<3d#FEeER)CPf[\=4A#eJ7E4BU.\\AI+d9a3F8,IR&A@
GSX,7-^&1/XF#cCW3fC?aVO)fHf]-dfVJ5M5O&.9.Z]#H\FXM\)U_VWY<Rab=LRK
1/=<_@Uf.+V>=?g>=U4JE<O.1D\?>]1:1.OaSFY5c^FF<K)87[+g/772FXKe8D7S
V[2\XKNO.,=JU7++a?4Hg\a#[_fYN)>3bTV<>fRX\fJ=C@FMdWK.;ZZDOQP)afQU
7(fY.E@e@NYd]JQ3MJ2eN@^67OJW_8+:O\^T+CI@ZfZ5DdeU0J4RN\97WW?B+RVg
(OgWZVX[FIX.H9W[;F]63>HcQ#Sg<.?8-CH,7Xe_Dd[6/PF0G=6-\IEK)S[SR&6Z
Ka1>^]5J=G?8)59IaXSCSd.O;NJ47+511Y\\OJdNbDIMQ=gJ[8Be:bc9O4Z93DE8
9U2CVg?>H31?7O/<CBfc,,E#-Y/9b3M4NF60dbXY2-D^OU[OMV,L:IB>]JN8[gI6
])a)?bR>IMMDGL^4J(LZK_JUfB03OM-cQ\\QUeZ[+CE5.QX&P;3LA73&VHDNKX_F
WgNRG>=WYc0)<cZ@^L>^YYY>34.(+NG=7#C\,J1.STc4_).B04L4P3E7KEB4^a5Q
IOPL7D71Ne9_.&\.7ZbR3KeXHC=c/B>ETM20,MKGYgf<PB)E+0C30f,(&U:CJ;)#
K0)=ccN4gC^CUa>?f95O^Z]f>4U;OMa24#;))Z3;8J2S8eL&[:?9;WEfQVD2N>Y<
4[1:3a3;6PBdJDK6C>P_]XAD?]8N.C9G).#(:2T2?#F-,_fda+CDc=&2)X]+XE&?
0FVg:aBcRd\8f-Og,OE2a_/[_Y:5eYc1/NALcPSD+=6&2YJdB^)7;dbK;daC:cB<
IfeSPgg_+FB4/K8?:6I7,[Df]-<,\^+e7WN]IVa08f:Y8J_&<MK.]HI8>;5:<X1Q
6?6TY>B6_[,==c2RWAcF-(L5-;C-aSC=/(K[E:d9459cYK5^H-MMS,1_&XXSX@B7
S\&C+c2/HR@:S;>_W9f<a1-T#_>Pa/]KBGY0/V(1XS/Ng.40QCPf#:c;FD7&aZ?b
.#cOdIeJ&CF[/?]&WeZVZ7JfbG:I>LI].OWQ+Y=YPGWNO/)2G^Sg8]CcTH.#&K[1
1D1BXQG,C_LJR(:\]c:<[C#1.D?Ve_.#(NYC3+V]#?V,3N1Q#aVVZIZ)e12+fb=4
,@eV^XGHW]XH6IgIaC&^BAH_S)K]PC?4TS1fJQ(H#I(\>T>>5GZ.ULO.@I^(S?D[
PJ\bK>>@4Lf1_+5gb\K&.RbD6)A2NAa2B]UagR8?bX7JafAb_GgOTcO_=DK(80a1
K+3MH2<K/-N@BI<:bH\d-e,+-#?B.F3D3ZFG<P8;584OgX,:0XZggFJ@W:_Q^1#]
1C86E1Q[Ig=P,SXf@G+aV)LNO#7-Q^g.g+QUS1@X+8E+##^A<;#g-#\#^e.BW1?f
eg]&#a=UC.S-&Rd([T/X5)5W_FBc.:?MP/MRAc\3N2-;D+88MTX0/)H0eS0RJA6@
_dUa0YS@O/Ga3cG8&[O5MR_ETENZRT6.HdDC(8FK.F/9-)#<Le/(3\^FKO+W/f8+
8\<b9\HS9?F^Eb/./L<E:OR^WW1PfdH\;(WQMR?NFd34E@0Q>75Of.^/aRG@<&+A
_MPT1E/E+6=WMK0)G7\;W3.[8(QP26AaWa&G(Lge9@,Mb:2F<3.QW<(6(UNg&Ud;
#.+;L6L6:5C>e#T]Z7g20c/D[eFfN4dBEE5H<;;W:I0ME>^<SQI-9J7;I72O=&EI
YQE#b#DXPTHS4<NZC.@f:U9LT5.f_-[DX3U?UI#22)S>aH/5.6S_aVJKS.d:P;#T
e+3\bGV>9]O@)aE;?CM0KY2gTf\Z3>:\2HPSN5Z,>4:eC<]a6eMb03Hb&N_efE3/
.5._DgU,V+M.?W-F9MA^BFYcG)Yge:BU9/+W0ZV4.c;3<S2U5g6DV^>I6>W6R#8(
^ACJH6Ff6VWc9M[4=C_8W[6701>=@?I-I/#Z8;N/&945_P5M3TE/F-5.E=efO]G_
bR&0HeSL0R@J0QZA=.f\&694X95C_CXW6QWC-f0Q+I02MT&7:G_^-RO&e\S^@,8U
]1AP>:EQUF@[[@SD3_PRHLIDB5^)c1UEg)\FAf_&3D(dT4b5;((+-AbQe@bQa^O8
OgDUOdA>A]3:6ECB2:R,+[53-@\&RL968N.M]1eV<J(4/a=?(64UaE0ceNI\,dG6
0AO@JNRF(1Qa<c>A@(c9/]0Q<<>YO(Db>AdR0FR;9VNZ+Qga05P<_5CP4(AS_=b^
@8.>>GWf9a&SZ95)-3aS/V+f^g<5SS.Y87[\B.E/H4-1J56#I/Z(A=4eNc)VZ/RE
]a[c5_,31OMT2Y<3FQ^.=7cLe0c]&(<^@Q/;VV:eYJFSA0PR\^+#>2_A@C:e_#0)
X:cGE7&aB[Y)gB<aga6/A[3^[CSI/8GUR5_LR&Cf<f)(c+R<J^A8NZ)g[VGe2.U=
<4TP.B)&fM&)/7=P=N3bX9aI&DU/ZDAIgXO@GXY(D=#P<@D9e.JDZ-)4]NPD;0dZ
Na<-9:#+^7c<[-VT&+>Z2M=acY146T\/g6.1G^OIYg?Q^W^A:bYcK?cf@EOIHFR#
)4R9Z<P9J:=g#^RF&BaKJZCb[8/C9dLBbGC-2,HTLLCDb0aKb3_G@E5\FZZBMX1#
5XMHORV2BSQ31SN(T]GA80=EWEHPF1=dJ2MB+\?0R@NVB[3VK)Oe-&UbETD6ag62
-:BG7aE^>CP1#?b?/TX0,P60Z?eB+@Tf+fT75cMB,Qe6,=?LA@Jf2\;[7&<SQIc-
^]C5=Ic]\<I^UBN4-V.FeB77R00Y<U#Ba:TVe?=W[H&HJRN:UeR(\^++&?J69&g7
a)<E?/K[S1XLW2(E2c=YF[#@@PS<UO]#C.[AgOH2#K5^-J?]UIf5fa;JRH0YJK7a
NLK2e(^F2#LcC(/R]bO;/S9VQ2=C4VF),7EbEg+R&GgPMZ,1>QZb@MZ.Xg_;?<HV
:fU75MHV:^E^1ZEHKO9L[2:8.CC-G5;83@KFaPGOW4T8VKX._F;Cg=eV85]C[-:b
DRD_U_gQT4<[\FTb>NML\RaFC,ED5>S:5fG\:Cfg^:B0Z?cJ#F1A=\2,e9CUYL+Y
,@+_UN>e3>cfO5U,4c;Y:AOMV:e<LEH]_-)AgN0O1D#WeV(@KBUOTB0.[NLT^b@c
5;+?gJ\a>NF229O[H0TdI;OdEG(J<BD=[d?S+Y^P4:QBO?^(,6L-QF7\[D7U=GOf
gRefA-,T\:8]1c9A7+V\.12<,dc\27BK)F5c<K]HfFPR,L:[QJVKaH964\)P3I9g
WFX0<UYdb\O]H^g8>SYO_MO+Z7H#7/2D@-^0=+MH4;gPF[#AS0USX8b&70Lea1CO
O,Vb)MSI[N)MG@[KN^Hc[(?b.U[O3+X>_GD#Y>N.-V?Tc//S_4DA#-+YCc]V38[G
VP77g\d.85P&A:S8:1)]O<ET;W<F1O,I@/_U5VQ5ga:I/^,Xe=;Vb[4BV:N\(U5K
7&g^>?UP&5eNGF1E@85P3)F5\6J8WY0,V;C#g(B&=0We+87Pc_;&)X.Rf:OGXGZ;
(bG:Vg7d2FQL&.FIUEMTaT9&4>6-0FJN-Y@C8eSSDGK#W)>QW99U<d]ZP_eCZMAC
<-JK=10CgXWbL2-b<7J@S1WQGSU<Z.CSN;H^-R?).J(::(bH)=6--T?8Z7XRT84e
Q,7dWDTFDFYONC6IB]cLeePIEG&7cYY>+4cE[HZAdL_fH6#I1K.^YD/Z52N6^5(Z
9?B#_-)5P[e;[:S;@T>MIKTWNOV1P(fSZ@f4M,0U^V5[)>XPRL1E=0^HKDgRMMFI
SL=-NR^)U&9(G<2,B45[U@+bRP8:\V<),e(47+II0/gc)(HVF7B8;YHLOKL[NHcO
baK\1@EC^Q0A^I\4B4YT0-(T<K@<,19^1eMW_W;?TZe^1I6C=#H:aV#&BQL)._-J
E:L&#I2;DSQc\)7)P^U8<dG6H\1;6N.ZG8AS1;0C<EP=DH/=W4@7)U?>J/-2N,Kc
:0?KFZcbVSC>VV<E8ZGAJaXQ\TeL_?JXGg)^ZaSF8NPXB2dP]ET0PYR-.H=;K;,F
f1YAC>A82c^EgS+Vg^_ObUa<@5=<(K,Z(T,DBFK>:J[5E=H8Q_)I^-E>DGc>FUO\
KKbA\^#\-F#(P7WJfQ4R66[e\3edW=dDV95DXFc4\O[cW>8S#E#MB_J[6PJ+)/g&
U.+=L3Deb)+2LFOW9Je\HRYeR@67YPDJe-/;g)OI__N=]Lg;e:0+ZC22bU]=[R)Z
/54YV7S/KMGE\J)S_?dU3KFQVLeC-Df=WY1[@,feLEGSGLeW(4LHeWW_5f4;?UEf
/Q<RVY&DFf5B9Kd@RGPFFX,8P2.ga.<O#(YG&^.]gA+4@NUgIJ>W71P0AT17GN8I
Y/:V20YR+SWcT-aTM:IX<Ve[SAY6#=[d:M_F22@#04^9YaNIB906:7KXK54)D0NZ
#IfAJ6XRT3PId@@<P^UA3^eKSC.I,?@MQG\^VC.a6cf(S?E0<2G]<_d,/SK8^gW&
E?=MPcOg=V]dC43<IEaW[6X_TV(0EJ)Z,aVdIbUC9):8AVLD2?MCU<N]I,0?XO,+
f5T&?f/CA<7>6_YM0U&TW;]5\0(U2L3_D]0[YU]Y7NB-:U9+C872>Y#1MaVLIR2]
3aT861>M23^^EfYBK7INM)1aFL(P<DDGDC:@LL<^<\d@A\><U=-6UV3LOeMT6bG6
R)1fZ_,,NOOCY\eN+81PbX\TXg,-bW/RC3U3(VI142P7<YS.S/g7f]LWaEgLf1bJ
+/eS&)4FVX;D/a56XFX&FNbF+COGMgeZY6@MeK4Q_Af@gQC]82aMH&[@V^_SI]^(
X<)@2W=-3bB8J4NffD>gAX)J53.TL_Y9a^5/gIIW/4S#6f,&HQRFRX,J]Tf?,gIF
.YPM]\-:,@;NdR:L7Tc(ERH&OM=DaWd9f_81V6N[C,G^ZBUNYOcQM&0M\3@F?0VE
=Bf]J5R,6@0Z_)VWaE+a33I5]-\#D-1/&]HT0MW12>/_IdK73FaPfRX>B[?N^15^
E2cb-J7fN><&+=M&;1P]08M:MfCa_1?aTQQYPKL6PQ38CEJe60Hb^:F70C5Q?B7f
LH><HO9-2Fb3218P9\@A93DK7;_]K3;b<@g.+HUL:Yg62DbA\eSMd^.03e)3#7(O
6)afSJ^YbUebQWD,f]<GI/P-Z,fBZGL_70#gN]O/,1IPM?..5IT+JA8]+)gYe/?b
H-)(4_2<[DRda@aAW3gHOa:.?R)25BOX0(53DgL+MfY]I>ANKV+)YJ4b6f,\gLTR
.XQ7ZBTMAc+dId+N#0G6O@14ef6K,7ff-\Z.Tg#?D@&7Pf-#-:0#7&N-=6I,MRU(
Z:?SN]/g65UO+(P5DP)Z3SaM=a\[V8?:eH2U^B_N-IKRPH0]2W5Z&JS;=VP&6-27
CY_QbF9)04S_JY74=Z_875I1H,2#PY4U4PPdc_J9abR/LKZRWMQ&eg+_cd()N6FH
;bg[61>JR?]NK9Z9CgDPY,J;5fIB4D8b#I4gb9+?[>1\-f>aY-1E9HA-/e@(:(N-
Q<_Wb0H^\UK9b1aSCU+d7\_T0<[T(0+4.f-/],L1=O]71ff\T^Da+gYCA]P?4^H3
KeY-?CM:R)JKW<32HD23BYX0CgAC>QY5C@W1a#ZRf1ZbI[H-4d[EHU0.N6d2V(XA
[gV3M-<Q,A1L3INb)2PM=?ZJCJO<2J=-F^0.8fT7O:YIRK[gD15BSH(QI)PI2A1J
WD\Z>dbO4[(QPeHX,\+8Ie)1#.2:B_DYW(J@QX^QK_ZM<4S:3G[VKYF/[6KfT7-&
(FL:G8bb23,ZfR1.X+e@[(<ZK-&>=?XEDfX_=>4f<Jc:10fHV-dWRN9HJV@+/H:L
JQ>4YT:5Y\AN24eb8VbREgD@EF>X1A=A(-04\+V+Z6<SL;dB1UV]J6YF@(NCAC2C
HSL:&&dI66aYCH]L0dMA;?dEGG8//AfHR+7e^(;fJ5HE-f,68/VXfJb.b_3/f3,,
<4K<Q7PY/ReVY+3.FfZ2aDPIaa.T,N4@7-OdR.L9[I^OCJ;7FIRE4R\7Rd6^b\Y[
&Z[?R4[R6gYV2SOISf29V?1;5CK[8WaE[+FZH.SI9Ab(+?W]4<=U4>;]0#[cZebD
.2^T>S]BdIdK1]MLQZQOb81@N+b,G/)X?P6ZeIG46T?SYY29@b?@UY4CU-\KUULE
7Va#;8>,3@;1=VFRG?Y\XB7P_X2gQ7([IDf@O6>E+EOWbRVYc[G5?>V,&,-W<5(e
U9gRUV3N[DI,ZE_@(OcWGd1If9DASK:>9DgHPC\-JfQa<]^/B1:W7VJ)e,75^S\I
J]@1C9T9Q7#JJ1RQg&WfC+V+&Y:JT#^=CX?F8,[W@\(:S:g34/.-<ce,Q^Z5Yc#-
gV,_F34&ReSFg:4aE?:-TaBSFAV:Z#ANQ.d6#6]NfVF,W;1cUDfeW?]6.-V)7G)Y
9FWUgdC9_BM>H&G;RU(L^aA.2^S1DfDHQ_]RMUcLR8<AFW(KVVUMLbC7BLaXIBO=
RF468L2/FTM\C\cQf0R+Cg9[g,]1dYS3HTA\_+#BBYK=Q2H?RNWaL;=1\7[FY9Ne
[KaR(P79Z,O/PSLXIH(Qa2Y@YA?M2WMR<H]+?YfGH96P0RYeH-FZ6O.1,3<V<Jd^
#e[WH=GWbM2gA)TR2H3S>ZD]MBKL68F>JNX4>D8a>O4?4RBOL>J\a4;-/-0gQJ-V
-fKHM,FSJPE-T0bNH]:+M&GCT+R9<ae274XHbTc.gP05D@=\V0[&,0Jd?0cMb^58
473HT4>-fcC\B<8])=.eI.)XcbI7BdG;,8[g#/D\^9[=YK\<_934@]^MSQ#W]LVa
?&g>P6:[-,#B7GVV/CgD\_1;W7CPO?:U.J[H<Z9A2b/:>^Rg<AWORRW9e7J3M_F]
;+6bI\+M^U(5G.ebX](ZGS,cgXaI:K+X=E_8gCHUZDI0L7RG=[[MS7ZbVd7]Q\P&
RU[2L:E&bgE^V]2VUP+2B#3&.6a)bfAO@<12X478R]4/WQ--W/3_K:_d4U<46GfT
b0bT^-Ob7cS6f@Cg<fHL>d1+H^Y926?1,(NBJ4:bM4<\X(38bBe?SV2ZLXQ9M:KM
EZ^?H0:OXV._0)T^FP.6U]@e+E\AF_6,?Z<a-If3&Cb5)C3D(FWGQJ[28J2G<ZUg
=\+6Dc/5#[7c/31.b;D&Z-d@Z3P9ab\?fdU9?E]FBc73d7B2G?>@,0<VeeW.,MI+
6^B&Jd1ab.(&?D,KBPb(>?QEBHUN9+Y;T.bIVJ4fZ6HAJ0<aIQZ[F(HL_L:7B81T
6C<Y]-NH9-CIgWKbHG2.&/D@R])g1U\gY)YaY[KScGETDH1>WcIdLT\6UR=T,Dc1
.ICY?:8HFd861Y#E?@MD[:S2G)8F&d@WF/(P>Wd>TZQL=73ZLD)+LR=@_P^LG_A>
1OBJ?,BGLUP<=KF]KHH:3-?=2UJF181<C(N)9PK\2?B]5S.cUK/HUP<5-_6.ROd]
T-e=>7]Y[-C0E<S7W]E6gHE[g@OQ?O#=B6Yce.H.eFb8]QO:Z#<@R3WUA9VVe7\1
V_+46cYAE+@gbcJELZ63-])1S<-@X/cV3N@K:(ENd\c[Q[[M0NOJ?0YARM7KG@e=
4MAC>7W==BP<-#D^Q++ZK##]cB?,;TC9^8Gcc[+NO.)e5L#KR[DZHO^_17Fb4\@.
V,)M#L^,<[3L(6J2\-CQ^O69#^-M2^J.\8MQVQ?[5bc8]6.(fUd\DNU2ABWAcI=B
b/XAB5[HRM#_.gN?09,K9E,G:34T/T=JD-A&La2H:R(ZEBW6V,N,KE[)_1J>MHd/
1LB8H,HPg?WLQAM[Z\).)-7=,NNT2.P1(B3[RB^\+)LDU>,+I#MJM=4O:Mf_A/,B
Ua2BV3T[X+0]T#U<U-8US.<@IJa.0e:U-aT,4Q\:2Xa8LLa55+(/_dU4C@_E(1/D
Sbc6Q7FGSF+aU+-M?G3525]=@7QOag=U?)@W^gD:BD+8D$
`endprotected
        

`protected
Y4R2Z-]_>+W@[#@=GZ3G4WRQV-:\BFa?/J4VM;afc=<HP17L1TK2()0K-EaV9dP@
SRg_eF-6[b+Te[[1BDA(dFRQ7$
`endprotected

//vcs_lic_vip_protect
  `protected
P41c0@/Bb2WW@FfPcC<D=OGK[D7Z=P>bM3Z[F#VB^7LKJ2aW)0.R2(#_+Z;247aR
3@^H19fC^b5VH0/C1MBU1X&-_1>ATA=X6\OO)/A]XOb3(/(J@>0RcVC._2^:9:N]
BY>,.EcI33KAU\6/ET?GW;87\_a@]3^(74YX:B2L+eQ.A8H+M7)MM_cM@UG-S#NC
9GJ8gY&1L5BMY8<G&W\:HVNM,BA.-gZ?3S.c1Oc@\;,D)WefW_g(D]9YI88T4AFW
Y5X+>.ROK(dJM<]HfUXJ/P]Ie[L,G71e;,cZ7+@YTaOGA3O-()Q8O]B_BJPLeWJ1
-,9M>IcJ)K[XT?XH-7Gb^6Jf7S?e&VDA4/.I<gM41A1fDK.ZC64L,O8D#RRFCg9Y
LKe1=a8)Yd1=E[HN^G=BU/6YL+WIQB3]RI\N[VK8J6F>VS55_N#O6&U+=73;ASaJ
^4QSJ2Mc@S^UQTg-8NAP2Z2S0fFf^6)IE&,=aSfRX2fB8&?WO2(C?B_.@)(^DVAN
.YK<S92I-[GNTb+ZV7SB8aGE(:CQdHG97E)NMCG:YCXFZE4dSW7YIg,RA3)I=5Y<
:7DO)4GE+MgU7Y4K;V6Id-\Ma\H09?Te>2eVSMXI&\DZG;9d2;28bV]?@5RZS#HO
79[25ZC1,6&XTA&T/(c:FY0RUD=V\QP>ddVCFd[1SIc0)(KD0HN,FXF#7K&Cd00@
Ff>=#dI,bNF3&K69f4B3J8gW(+M-6Z6M::Y3Y.[;UONd_]S(V8&XH-)04g2<+1>e
RG2Lc_U3?_aNMa(CUR-5dKY;AC=cNgT<S-ZE+_IF_5@H9.TO0^;N-SV/4\f.1RBD
Q(+4F&MaEL+(-e,;bCYWRfS=WR/_;_(727a=\H1.MT29>=N<M8EeQTX^N6b#Eaf)
+:>>W/bU/+-<a^Ld3Y[YK8(5U7,24@ecC_07If]72MgB#6>QeA]Y;V>9/CbIYT7c
/KDR^fJ4/3c]8Pga3Q<a]NP/?BX4-LXW&CKF]X=f\+YA9#;2>>]?[#D_&P_W@a7B
b1dc?7)1>8J^8=8\\\1[cC^4(MSA=Bd,Sb0+c9XXCO.VO;Ge1(RbL?@[X0AW9)R_
OR/C.OZZaNfbDA^<>HVQ?e[+RIbF@^4Q.4+QgGO-:^6f9_ND)44@f;_G_&HZ[XcH
d1G54[PWfU5/O6W\CNINYVX7QPb@F^c5,JW=CPKg?_UL=UCLTJ;@g3DT:39X6.?+
@R<R@#@SK?/FNRR<D?K920d:R;ZPQEMZ-V]IN.GCcBS]I75HERR:WMVP.;-eD25D
@MGZK-&YX3W/O7AVL[X&aWO:bV=_I2_7<L9=ddM(3&b0c-Sc@W&gWe^QNAHKPQH>
__bJNefE/\4XT=K_LW],GY:^cefJbP5YC-Z.J-_.PKT_AC#EZ>,9A+FL8@<G=a:<
V_H7&;XI7f2,(d-#J/Zda,J+6WF)TdfHE;g5],H[8.P\[?9+O30U^@1A69,8RL;M
I<&:2\.0_;:)N.1Dg@QJFZ#Y0Sa:e^WAHUX,#Z^#DE1VQ:AT\[ZR9?@O_)^6b5:Y
F9>.Q@c9PUO>[.M(H&4+Dgg#bPg36-0T4S^Je[RGc^U;N:K(U_:]3J.P^P<g)?_O
<7g6b=C+A=B0[WUJf:K])_Y5Fe[b>L(#9@DcTDgJEQeD3RIeX7X)+DL;e3X<E<AK
:a#aNY]H,RCR53dgV7G@NO(T.f+RTG116b1.Q=(<BUZ^0><#eSdW0Bg-e2eZ(E>B
VP>a=4UY+WS2LEaAUV/H=FId3K=<f_D.SB-eW;/?S@LEXH^f;ESaBPHfTCO:ND>8
ZUVZKG3H2;F@H[=T:]GQ?S[471(X)Z<<GHLbFDGA4VGV-EW:[Y?+@2b0L(DRD2QU
;+O:?:5N;RK+<[B;)PH[]348?C4P7&b#2f+&9H3-VL_RN=;0]W#^R/@W2a9B\,c/
_g[WB]GY6;/4N_1EELfF/C^T>G\Q/4bP/BHa;b_O/)g+&:K)W-U0;1)3Z-1W-+ab
&R7\,N>#.cAfN[a#@F/EO<DF5dE.e]/D.WQ5UE3=N^Zde#EN0dD&b:O0d_fD7PFD
M@YS.5X+f,TFZTEY4129-&O;(fN(P8XD[#.6C?Wg:P^4?S@93=?.<^4ZTd/2F?NM
<N^D]e;1,8Xe;0/\1JRL.6K_P\e7?d2gZV<T^_X7G6,OGQWEQDa>=0bYY7P,NY0\
&+eXL9,1<YHY>=W0,O34.R_B<NO2AIL]8;PWZ+//b-(3E04_<^W6RfdZ;B<I->CL
BS-^c.YA4ZM3aV8SXDb^K[AI7dVLS.QK<5IW]Q3IIWbg\B[5<>^&MKX@,#16H0ZX
2W.3R0JBaV7QbHGeZVOaO+^]-0)[4Y-#@1&]gR)O?\Z&cc;>U(+&a0E>ag8&2@b>
NY)Dg,Zd[Bb@<Z[EeR>\4-2\Sg=fCcKfJ,.6>4IJ[M-^UNQ\3(LV@7-[75Ved+Q]
F.+JZHF5=N_L7V8TROQ]7IHSJ1L=GA-X^X-AB8P\[<a0/MR#)b/e#W+T/X9fe=D,
:a(ccdf+]FRee4G^8/FPb-4_8XYaGUB,8)740B\3cEF)L)><?KBGXKO@/acbBHdI
\85;0N0b<\O>cU/4V):&,[]@IR#_JbIUN3&+a/BJP)TLe<=P8JYL(X8I<C,d0LdW
c9#fXR>fD\b\f@C/GHLMEd8d41X1:\@2\]g/e\O@=Q32F\1[?B:H7aP1-.IfWYaN
bX/09AC.<1M<1\FP8G2RcDaL))XS>)gTZ=Tf0Q5dR6aHSfa\J<[K>._2#DZfCa/R
9@g=IOKbG&F;7[2,G(4K-8_Ecg/Q_EcFL^cgISHB_E>7LOWdURG^UBU&TeYIgS1[
#fDa\fCT;bcH;+>SU#=E^J;ID8KUJYZ^IF\LW7H0(86D+WVWZAJ[.89>]&^)#K&6
2UZ2LYf(9WFR6;Gc/U][C@YfCaF2AP_0+,Y\>-C;c7aH1XV7b(80(\W;P];J_C:K
Z-&D047_M=#UC<8-ggGAJ;@OM\cPD-&1Q1>9W>I0bQ)#^P[DU+QJa7A7]:0=bM:?
7_.=NOf>I[F8X4P5R=c94VNH^O3b-]/8D#>eD/0Z@0+6OeWZ9_W20<D26W0A\-&W
XaTHH_@:1_1/71gefV(]Z)XD:^6<gc=IZCL8S>K#.UN^5MMB>0D1@X3.3Y\)7BRY
JROWRZ)Sf1Fg=8VUB=-26AYHBf1H,1V.-434gIc@841N,01,L[^d@X_YO[7H5PY#
)Q>LGdQ@Y]Ze?Q5(gV6L-;(b6bPUY3fa)Ad>VI<Bg,L]a92ZY+6GMdf?A<12gKUX
#6e0BLC9f,D9;PS7)>KI<0EYG9Ag@V,DYM?(7>;U@474T&dKMQIF^H#(BdT?[8M=
KVLYI?S7Y:LJcSWI-aB5^A.Y.;\9)Z:ccS4X_T7[\F>FKMQL1OX@_cZR)8fU9>]\
;K(\#JNAb2VQfY-@#<3FZS4cT,F>S?bBRf:dPDL@1Z],F@Gd&4G1b27(?Y<25.0-
5&6eR+2P95ZM/\Bd&3)EN(KG-C,fe#RH&Z.<X)SBORFf=)@V0+UeE1<O>NU;:2F@
a#K\;0?gR,=XUP#T2&fFJX@,4@&Rb.^OTF+YRQdE+R5HU#+eIO699(D1QHU1HS<-
TRT1/4ETKO3KWUea8K#:[ZM3\f/3F?3[2F]2PFd^,MIPN?P1AeKJ5M91NY]MSS;-
a;H8#4=2H05;@\GZ?Tg.2<-QF:c_F8R0>SJNLHF[RLfF[LN>e(L5M:_A?H65#a@3
ZG1?:\5]5@&B(IJ64BM3.(=NJIYZOg\(;X.?CB,@Xa23.[7CPH68_B(dVXJ:fQDB
HO1?&aKBM]a2+6>G324#N944]([NV41FZ;4[4\J.\A<&F620[(e\W[7g)5\M^dfc
eN:?af_FXM&\M74XR87^95>ab)W_YFYGBbG1N#HNe.c#_O[]PL@LV^\(RR[?3:,W
d58c^5[#H^aVd&UDKX;XeB)L,F(.ZMe4,1ZO2/[.U:ZVPCZ7G8DT5K5;D<e[3W.3
[MLb-a)CHXPF6_;G#^b70<6(eMMVJ=DC<)/VE&V6N2J&)KN7@Z629C.\]V5J;SV1
dD4;MAd833^5@0V2Je\F]X]6A(a\7Vf1P/S[E#E]/^_H4WLeBD8e=3^A;WRD)[D4
-@2YUgD<H\Ie-(,U]TX&KS5_/O?\KFAc()9cd0[1F:=K>&#2TNGDSURPfEA]@RH9
@\F_/I=<J6#/POeRc/AIBDa/REKPTgI[)^1V4fM^<V&U_Y/M&^R=Q5<^Aa@=T:Gd
IO::Z.X=8/:a17)#S,1&MUaNFZ7+\[E21B-/+aXE\RQ,BFQL:E18-4EMg),^]N0^
MP7LOF[_5@):(-.SO<1S2T.BF7(XK93F.AfJCX+LcYCH2VMeYC#AW:bP8dgCWcVN
>D)Ue3>[67WP]Ta^YS>(gI.XUB=_2XK(fbbL=MO0:(c06_SZVG-+U;HdEfI?Uf\c
c#\/>ReR:T=gQa2/U@CNT)_5HPKFV7F[?_?7-/R((PT+5\TW(bDY^b95H8G:PCM\
b]Zg:RL2,,58beT8E5;96aS@9C;[DUNW5Q@Z]0g)//>LUBefLUe0]\)UV^_O1_db
5L5dd1e2F[.^++56(/I1G0\B96e4]BV,BQPI)SRJ2MT][g\F^SBTD1,7-YFE[<P@
]d67bfMF/>PM5L.5cd]f)Af;Ud3K@():4P@)HQ))K/7b+66#e(a0Q5LUM3-VU_]6
#HU9gC/Q,ZZPKGQ?N+VdLH5MPFa;/GDK4&:VOSc\Qf\AgIML9WM>Le&WAN;)OeaV
VNf\M:-O#J]R<C+;P)X85HN?^c,V+]9OM=BR2c1N5@#Vg,eE6Q4;D9ZGeZc8Xc+-
>fe+4B(L\SP60;QFIQG0YS@,cV/f5A5DDD#<G_J8G)FS?[(gTEIf390YXLZ@MA(5
LP-]1LbQ<E,\He8EN<f2&g;B.R=dQP-P3HHWH-C-8fQ)&+Xf_,UV#6aR;>0O<K#?
1IbEW:ZXT6]._/B(A]Y)M6TA>MI:@.RSc-+LP3:-X@G+]W47K(/6ad[YO<G/L0X^
TOf9I>4467[;cERYa-f6eSe3ac)DKU0dXG;4>JWGeXc4CR(a5cKfa-DOaf1N8Z@A
XSWI73:WDS4DB7FF(;C=:W_dg:Fe0=SLP[D.7fKK&8;<2[6O#_[BRW-W[)V.Z//:
):GPbfdURC@Z;4.MEND,_[C]M4Ae_@FM9.6U93>U/SKB(GGNUS7M]N35>^3WcOA?
C[ZW0?3N4OPBV_U.NaTa9bW49(D^faf6KS8^4FdM#(+A+H_e;f:IcI.8RKBMZ0c3
&5O^eZ9R:JR/N9W[<_e(QWQ.:a]GD[FWF,W)#6D9B?&LB3J^/#[0TK2e630K2:7(
c@8=I7QN.5I<O\::,g\SZGE/,,F;W>PF9,D6^YaGXZ+_>E]d7bSAg)O_64(I1MYK
A@]F>eeXJ]C4/BF(Qda-GGf=RefMI-C]/N@85=NXAg??_CE/G?S72Y,g954_gYDe
/D_?ER4:MT&g4:dZE6QXK2E@a<O:=M)(,K\X@.[&aS^d];15WWR1ETCA^g<6ST;I
_SJ_BXXLY3S+aWUF/#KTFGG=b8T23dE;:N-\PU=SRaZaM5GCDD-7/S,U,[YD7E)V
\aHS62/5>SXIT#VDY;If+B.96G^#?7cYAB:aV8[2]=7EXD>0\5DXQ9?9WYVGf>^C
>1R#DP_^K(eM:/UO,cOZ3EEB0,3c828YE3TA\gFQI;3L,2I(T4M;_532=QXgG:MV
4NQ5)^IJR24[UT@0P@AR/Ze:^])])JHdHPDRWY9E^(X]UN/R4D035=0bIG<[4KLZ
2Qa-M.Hf/+dPbP8VK(Q>3W:S\RYOWM1Of+<QY;OP8<cWKB76:dgU[Td)O=SO.Jf,
S@NXF0@[[+:3+./Gcd4+[DY=6U0f\3]925+#>CaV2cIR]7WF:FZ\]/N>.E3L2F-2
I;JO^R^[?^TSK]?)c6V.?6DZ&/_P-U?b[0aPgML6N,DU>0\g]48a0S6P;XMNda?@
0+;)<3(Kf+,:eYD4JcH>(OK&HJ^#bV0Ma;UJ1G5+I0CZ=N)/A/\d@^N[VA<2/dD3
7SG99G3QO0)B1fZ0L^+6=eR&BBf+<(56-#?=H_D2EC+QbHKBZ>96B-JZIH:IfBIC
X^[e8#\[I1?63[cIgg2F&b>_+;M\@L7fC=@D85<1@GJMNE=V&-J\NF1?AGS)<)Ed
&::(M\=?[1I6)\7IT(U2.&+9UGOQV_(L&4,16]2f+Qb,PN.2KUQBCLWdD\M>-RY5
/O&gHZT^-W@15=TC-5HY.(Q30?>XKSb@_6_ZHB50C3,.WSR+[8Z]8aEaY6YU[<aF
bT+;_^?EZ7AUS;Cc:/;e.,[WQLEM<LHOZFVVHY[9DR[BII<705>8\GS<R5VW:AD=
))EDNV<c,4=AM_cR[DBJGe8C4[A7E30.D<YdS&b\C6SM0#b)?VH(^>b_C2&HAT^;
;-@/Wf;.,KHD0e8S<IE,4G;4&6][&4E.>?)@XTE#8;b^@]N9B_W:f)b8fA\CaZTb
B\H.#G)b,+ZHIS+V+1ef[+g<9?LV9MP2;Lbe>RE8\.]51S]WF^Z(dG_A3,6Y,_L_
bNV6A/6H6=Z&ZTNS?>A5AS17&,:A/=gOUQB507(__?7OF,d,dUPY=--gZN+#.e]Y
FUPLe#Af3f/N]L_D#g&^5]bLTa7(3M5B+)^K(H<5J-YNQHRQFKb_N\=Nf&L1Z<QL
BZEa(f)e]L?[8U6IJ7E(,<;S0_a5CLX>Z1cU)M>YN@B,JVQ;BdD,a&]RgMB)8SMB
EI@Z=027>GecM5\_7K2LG^75ISQDB,fXf9I<5,)&dH/G8PS]>b4?A55R#.0X@1.V
XVTBQg:;8]&]E:Eda(\7;aKP20^M#\TW[1fe]-B&(9O,K(LD5g]f/f&IO+P=I#gf
G3P>+>+MJZ#WV:R^dLg7G;SPLNDf[)V1a/-RIeC@697,KP4N8gWE#Y>L>>.?+V=O
OXQGYR<FRX)#=g?(UO,Oa:4.dOL>:_.H1g)G.]9I[1&D=d0UbIU)?/=4;NLgIJ3Z
MQFgCU5LYQ:PeF_,0SUJOC.-D4F6;W@\a^2N<.e2@ZM41ZM;0GX[aTTN#+ABUT#L
SB]:V<-bDd?MB8+?8Aa[F5GP6E-QPRNS#2T)COF=&<a7^J;(K(76B>^S^CO7K:D8
//+\87W#7)M?L:=RA@RI.9R.]d;93>P--4cJ_CBd,+CO1<Q)X72E@[3[OSIW@N-c
+IaQ9NVL,TS0LCR&b/JER8[Y:26CHRVBgb=2;]F_#^Pd[KRO]G]?YDEWWZEfQ:&-
?(3U2@_^1\S0[KVW6XHX<W7NQ<B]#=-OID/?R<Y&PVLe^71PT9ZX5@TM7Pe[S8Oc
Y@JV\XLGU+I24O2IbVcOg_0fAOBF\#O.TOTM,;9I]C]g;&6<X7S1b(<D+Le/2#0d
f6_EcdJUKUFIdEI/QCeT#87\6SHS,)&@ZDfdS_EONX5UUAeM:YVROH<YUG5c9MD\
Z^LA05:[UOME\&9JIES)J(9Bc>Z7Yf9G0TU^>2(FA#0Bcg3LVM7N0e2N-+PI((3)
gg:KO)BF?-#f6bd-GKNIN3.#4gODJ5a>SPFFJDZ5MZHIG4DB:d]()HILX6Q]A<^U
KD)<FRB@0g[O_45I[H+aUg4?S\D3(3bVHKO_c=).(bYS(<;PBDR?V.Q\JDcO9+])
O/6L(/_G>FF4e5+J=_dgg]XMeX<.#BSa29)caa<eJJD;+c;/\)G^6HJc4aC]=QUM
=,d:Z8+^F0?BH:g@f,6)6^\P6@QZF(]<-\C.c,:D>>>,4S0-A#dLS7cD-ZLIQfOY
7:Z>/cIG[D-Z?G\^]@K<85XC<J::+V26#OR+C5/V;90?0CEOO0K?=X,4#>JK>daJ
NJYGT7OTPC\RU(Od#\@XU_\A0IB8W_ag(BMM0ON/)3YabO/F(@-<LWR6P>5;\3SQ
<=.d2[WGIGHO8-2P,7gENM#>;2=d30KJOTd8F@&;28SL@NAU<bN3gfMR5:SS;8T@
HQ0F-,57fN7-Fa:KN6^fBJ^WXad2>W#_5?f;9Z3;A[X48;57J7)c\fg\e]cNLPeC
cD2A+8YNH/)1Z6-?b(CHa;dCE4^,9FaVED,M49YPa<+A4eEV@5B6B^bRLV0\Z&DU
[6AaQ^2CMQ<EC(N5URaea5Z3Y(=D(Y.3_cT5&:^aKPGb\Kbg,G]]=[MfR>Ne#<dU
ZZM69J5A&2QIN7RF[TVGG(YVQ3Q0VUFZM:JVF055J8,YfR7+c<=,,U85H6N^PWW3
(WV5K03fT?AbfEWP0KR5?(XE,O:2E52O/)f?T9fgY:BTRTAQM;Ud)-.:7A(Ff3;<
^V&S:O;C\CfSc,:^CD7@#I[5dS;CDO@@d2J3BEc;WUY20-(2P@ND.U5/;,TF;QET
b@>=f]UH@#PIb)H:XgD\5()SB0A=?_XYO_D_#L5;JNI7M9XW.NcC^QIS8,KQ2-\_
XWR1(;+U]PJ^#fN=D3@.SOAB.f;T@@?QM8AKdK&8E>&)/3:L7UBV@BNe9V[ASD<c
A)6Cf,97g/\WYOUge=GKG:gWHQf2,_^c?e7=G:#JO2<f&C5A+UT5M>L+N>V12A@X
?TF:,9^[T-<\bMFFP2Sb+Bb8e#G@59eRNOJ<4:>+[];@91HZ:&AN(FHV#M,c?^,_
Q#<.:MDG5Q9&W7QHE8XP,?O^?65QZdIO-Z:OB(S:dN91QN@;VDMDcd\^V:^:FI,S
^f8/FE8;>dH9)OOQe+#b<bFDb0W(d=HZaa:E,cP7^ETSL@UY<+H&:=9V[f6Za(NP
,Jc:d\E9,G7RZ8?]B/GaK56RfVR=K3CUff2@I0PNU#T[ERbAL3&(P&[BI&0b4D:+
@)FI@fFSYDW^V_T5//=AA2?C0.J-1RTAQ87;+;S\,a._4Cg_7?YfV0<aPS3_HM&O
V4eN7Xf?&&5-8@ZWg/f6OC4.c424BN^G[:Z.)dg-,K]0\A^U8d]JfKP:W&\/)ad=
;V8B(V&5?^b?;MCe1T:TdCX<K8@)Jg>Pg&@8GM@-cSN:>c&<Y=5XHb)-H/:PCf1+
7L^6O\2)3ZI0DI4P?2WZg[]f4J-(]KS;>^#Z2\c8RYJJ47)H_+B8aD=#&]M^U]SP
GbM2?5HR)5S=UaIg6HLMJ>]U+AK)^41@XFe0IgA:]/2,d9caeA,,c_,VJT+.]dR[
UFN5@4GX6-[J^/+eSV8.5+.6=^Q-E(.KL9[9A7X#^.I>>&:QVYOWfU7>3aUb\7D]
g5CM5J4PPQ<c@IJ@T1N+KJ@VMOEd>[^ed#(O6Naf@9?T\YcBMLZ)BTcSO,(OM5P(
LT&:Gc3dJ9bRgW,/+HgG4/HQ/_Y87f<+A]/P8Eb]QZ<E:&f)M&dG<;3:S@;1-V6Z
.2W<>f514?>89-H\:J0EOaHVAU(&IP-Fe,?(E&BC@MW\a:Z5)AYQ[[,0?UH7)7:P
L[S5=[0K0^\6;d7;66e@.LF;7M-/Z-BS<W.6OY@>7B9a+76a2,1XC3E#U0#JXYE&
1,G)_c0-gY.FW&#ZJVQ+E[8X+I)QCV2,&#QOW)N<E/KJ-_^:Ig/GRPUL98#ETW=3
BXZ/Mf_d?TR;/JBH?+eYD9S991]4Z,]9P=MLDLTZG&;-V/3,LaU3AXd>8,^H:2Mf
69N2Xc1P:(S0>T/)Q0-e6,DBD4G0L+1(dT#gQHT[9#]cf_LQgU8Sd>,YO;N2G6d(
_L:cLK-&^X_5R,.P(N[f:275Oa;[_J&B4SA/cL^JI(B#8X,OW&93Y;a#JRO;/7Aa
b<@ZLFV=L-5CTGN.4QGKFZ=NK-ed1e+aO3&-Pc;72cG=I4TD&^PDPW>@HbZ;C]<]
[-<D;CO?a[?HPAXQ.)E=:I46YR^^HCeQ2MY?LSA?@RU3gZG#),_:U[b?FL)1[&Ac
GG?[YT:DB70dWZWL#WNKWe9/JG>4\c^JK.ZP2]MHUQQ09R]ceTI6]IH5.UMFC^]D
\-/9Uec\2\YDeHbT6)>QOWP&)-aHX)-[=HOV_bV@O^OdG_JB.JeggR&8<RBc51U&
e<X^BE8=\(M<XQf9LE^:5PDa^C@PO#\a_)E#ePVD.<,?/GR)=VWb>#OggPEfK4/3
^>R8+PD9IC^TI#fZLd8W20]C[F@Y;9AUdY57gLD4L7(BS.X2gKHY?D0MYVg6[N=2
0Jf,MZ_We:LM42YTQ4b-.Q9TN<_,)UZeXH;HQ)UAK&H^?^0H3gPPCF32c_B?c;-?
RcG;2M1bN&JQFI(PZ>L&d,eKL4:0#[dUDX>T:IR?e+AD,Z\g7fW,cVZfeJHUYDV8
8,MRE,+NPT\BX4L[)KbPAHGF1:C8))(?S)UY:^K)=#bE],<Y=gZ3L/)Bf8)DNP0e
CH77A5ISP.FaB_e]5ME6K:HDGP1AXYK9Be85bR<(PS1DS5OcHaA;Q);2VIJS+Q.E
<Vc,NfbXE[)8#9OFD]MB]&+JSO=<,R+ZOS05V)^[e)VZ<bB7NS=^;&JcGL@GM.EP
_f8E^<+6+g+(<8F-W]eG1NK9ETJ5SW9cX@_MW\/A8S8S,5D75LFVV512Z5bEI.SU
BKG7)=<YY0I>2E<,>F&M#3#\W?3F#.]g(1ZH&-A<(8G-c>>4c_Z>\2,R^H2MR4.[
I-.0#[XGY]A?-FAEFHBUe)8&?,IfK-9#O^?)<8POSMQF>eSQTAU8]e6D,4ZIPF?J
X;Gg>bVeTK\:&3SCH(^b5BWU?15RUN::0]S0d^K:QC4>N:D]16/):2SG]#:\E/KJ
7-;1bL1Z::Aa++AFDJMb].a7Ugf]a?dT,(X#bG_></9T;UFNFMY1\#;W)5R8#BgS
BI+1_Z8=ZW1T+gW301-F-#E-,KPcP;<P0CW=\,+#-FMOBW/&Z._^=5GJQ/(#f)PU
NGE)XDHDgJ0,,;A[=3XLPN.NAV1II4#C:84I,T6b-,>0-38V:aN;1TT\M)e2/J.J
A]BHBZVb+(PeB74Q:Fd0TbT(6#5Fed5??Pf;^51fS7<ZCCR89Q[=L@Q&5>;KPV].
3=:>X(N>&HX;EF;W19Lg,RDQ2F8/<I7J,=6I>LL.:RT?)0c3^I:WgZZ/GCG_=1eH
/UU-[J2Q;aNaXZX>88PJM/U78a>dAUGEKA3[<5HR40c&Z\#9/+gDFHHeMO__678X
+10@<M+AaQ73bTM)g79]Y47(KC+E#??^J9SUU5+KU0HGC3PA<<gO-#4+9O_F]\H_
dF&D@eK3&K(;9G(OgT.L]=,?<RJH\<=(#1FZ=Hf&4EF74,T&B@+.RbTgO?79SORO
gB7e#D=F<5Ne>THaYA/];?1f-(9]_&,.:D-BRQ_QICGXKeN-=]W>I4H:NF_EX#<?
O+3#f>+G8L4G6).13/UFP0]VTJD^OZO3&CdKV<+9GPJ8++X<TG3=4^C=(C3AOM?A
-T;\1]]?g@5^+Ja4GP4eBXX16\UE<eM]J;#3><b;[.;6@UbVU_F5<4_:371(=098
+07-63e4>\U:4\Ffe(P/6&Y/MB;d=>)@Ma?]6d-T-aaIWSI(aZ0#JWFE#cKGS/84
J6#18C\K4OYNI#T0(EXP7V+4AA:bgPUYM&GD[A5(_C\-)ST3Z+>=@6GKK4aG^4_F
&M\@ZV#.[d]eDbGc)J6\4H,__/d<6.XFdb.0Oe#RU3NBW6[W[>-?0E7])#G4365R
FJCX/R1I@f.W6U/;1g.&KOe.A?YY[HQMJS.11g0(_g30e_V(BR,gPc=.A14(WOPL
^W>^:U(>9C/aV:adRTWNO@1JGYIGJHS[Z?DWY^5J(Y5Y^2]NR,3_MdLcD5H_UI##
FQ7?Q5]HRG[<9H7(Od]3L9eY#eHbGWD3WD3AC[5];:&ZLF2b2?3T80EX>7\LYcLZ
/0,6GE-HMMbeU7S]<;;NAK;1]9Y+,NZ<^&1?->=dB335V_;9Y4DPC+=YH:GH45d>
,a?/14#<+5FYJG>>WNF6gG9QQaM4(7OGAc;;\>WDQ(>X._>S8c4FXd&REaMI85<O
:MZ8#=-Wcb0RL8&9V?c9B-+7(HT?.HcO:K&6&5gX]d]8_72POM>NcE.8((>5M2a=
DfC9.S9b/E3&?9A,4QS,\Yb7.fg@#SHM;5Z3N4OKN.gfELc<T(24_PaYG?GCHBF8
I+4(B7b##Ld4dWL0DX.KI[d>XZaBY]IY&a7-_QT9HZcBPObg887e=LHD7VR6XG8<
PIM85]2_cU6[,V615D^5bPA2,baA&+@[RLG,1]B1HQ#.@W4fMaMSG+>OeIULB_<&
_=^YbCIe2;N3+eAfP]+ZH0Lg_g/O_Y;5A<ZE0&\W8:R9S^+fF^4265I-cI<Og_dL
]S#PfgQ^XRJ7165.;]Ff/>gP?.a<E(S@c4,W6M,^SY4W:?gM=2&[QABYU)99K8Z#
VcIWML0=)UI[JAK4G[5:V-&bd-J@V+I2g;\P1B8L7F0^E<+QUaG1]P<<&8NHSKVM
FXTHD^#R)gJI?R1U__f9@X.AS2HTIXJ)&>DI)a/d,XaMf4IYffVEBU]bD:<?@LY=
/2AD@XK/0dePR4VR7A<F88_ES.L<&LC756BW-I,@\TgH=/</TVEgAB2,]FV/:>g-
/A\V.EE]ZAS9+DI,X,Z+NAHT<[+[U.6O)F\TUA25H\37EcBAX79#-?.PAO=_cgH#
WKG?_e1D4Q>ST\8=?R0bXc37^d#RH;8HW>6E#,>N294@KR?ER;HW1O.G2R.BYO&N
T[AW+/eRK;3cLOGNUK/#.60gDN3<&fHYUC,K[VETHa#B_)E@a2-AWU]P^2B7-XG&
Q;Sd:Tb8=L0,D-M-U<84>8_c+.2R79J3KfG,_#5#fD_?dZZ0/_&93B0JgBICD8>E
QDI1]RLX#3I55#[P>4.;;Y:2Tg>d,Pf,ATK,=)<Sc>9I&^\R9I\&Q>_OgRe,,_ZE
:OYKBTF=._D7[<PP+H9;U=M>05Ua&6F?HeCc05S+7]DFc>fc#;VbKKOYVUSBL(g<
&&cbX<NP9&@J+KY=M-ET(U#O&:]fbLWd,+@3)HH2Z<g[TW6P\7<-7JEM4^^V216.
8Wc5a^d#7+PdaO8&GYTC#:cQ3Me&e7N\Xe@]dT,#GE1A3cYEWB@X<>4GE_9Y)f/L
O>#UZ3(#e2?PH<,/87;eVg[]b^Z@<4\AL?eEI\UcdXG]gRa[GSfb02V7Cf>C=(fX
J)\=PYA5XTMRYBT?(T4\\L3:/SXef=2DFF&LaAAA:F[cd^W?c@ZgOa_=BC@aM6XL
CT[f\FS9P,OL3;.>34LX/1af_^[-Y.ZTK98#5?L6I1VWceTTC@?OLJLR-PK+8IH/
YWc1f#AaV<T,/2XEZ#e]\<+7&YN+))TE_^U&F+LS=GR-I\GCb/]]BSVEdM-<#.DE
I@[1#&VC(=fTEF.TgQe1-XW6](I:57A2Q.(C1&G/LG^g;+9SGM-KEAKS-a9S\+Xd
4Jf]e3Ve@EJVUTA/P1:gDU^LRG)BAZFB[06edWH)BPgLO<Oa6\a</#D5?g6450]U
:@^+2XFc&NR[4.#GCXBZ_1JZI\NfSfe0A&?fHRINEE0YQfcGM.@bEc6D3DG5NM[(
Ta90??>:V=VdPBYc.I@PC0SQ^--GJO9gD:9EcNdN8NS-D,49eI-C,N+\I?AB+2X#
+G-7dUcE;7>\4&B-3.7;c46?1CGG/)d=SY([R2eQYJD8RA&C@?=?bX@E>CZKd:-K
gD:IW[VS<=1[W+BPES:58[\H-Pg4L?.51D?Kd?QQ:#g\[g@9.64U0P/62X1U3_Nd
<L1_.LeRES#GNS(L>.^T6/AUVS/WOb1dL^Ee&]e2;g2<,=?>,J@2Ug2U1U]V5KZ&
>0Q\JGVTQ62\;XIDFX[D:Ae@aS9#@AS6.47VXR@:R2[)[XFEVNJNgDFY8C4^E<?)
?Ae?H8>;0W0K7;/fS8?_X<WS)IJF9;X#=Y?O5g\>bN:O#@/6-JA1DG>>[bNb(79#
b7S]SMTEW;=:Bd#&)&R5(D48aU^U#BPG4.ZA7<=I9J8E\Z9Ig-P)dV;:O@&F6&JZ
WURc??=>LST28Z76\8@f-M=&0-,/[gN><MIMJ?_:J@\15=\CFD@IH=d7FVI?@_GZ
cM_M9QDLIU3J9fQP+Y^FG#1?R4Xf.R,_^(Q5@Ka\^WF/8L##=L#9;dfO5S8+0dC^
gXZ@2]b.Z,BH7@Lg]36<a,-[:#C\K(b&4DW-)=A:958-0BOD30</[5R(.3Cg9VO8
Fd.15W.7/#BOdC:9c24ULHWKQ8;T@3-N^YBJfIF@E2V/?VY0JV2T0CN7fF48eALQ
7O;SRTg#KSb3aZ_^#6GP8TVOe=D]-[\I^L^8M8QJ9;U;@S\/>^VB14HK10T&&<gD
E^Mg080D^#T(E</,YAIaR]8;>MWdU]4#21_G>9e.Zce_TI9O,e^fBGK[?>BAC]HY
^6#EI\BFMGJ/fO:_7(6>/>-abf4_I=J[BX_:c\IQY@UAdFCCc^RD[=Ke,9_P._:G
H61DXY4@PVZ7fB/TX]+;/+Q4MV4R/]#<YJI]PVS0.94>&e#(N-SOKdFQ&G2_#TTJ
3J5Fe6R-<:/[&_UA8Id0Bf;)WEY=EPH1GD[;3TN;QFRfPZb>JedcYD6#NYeMMEOD
U<e\:345390eOETZ&+\SKb9#S-:Gf74<@U(LR<f.2CR_YWN0Q&\L3e)LJgLFb<OK
^4]g2Z67>66UggT;K@>S5[(WF25X>fa);,WA;M,DaL=+(T;9Md-VT_5IM[eT\QEC
^1TU_a]REHAGOM[Y^J>2+?f)2Q04Y#a3O8EDBY4+>F4OAITYYd-I=\K5JN^DSHeW
S,0C<E[4bCKIHcdYDDTQ6eG_A&H_4\4G]6;P]_UQ_2<IBT&5[[HR#>gXOg)5RcQ^
^;RHZ&HN\MANRSR2DEdL=9L_J,:eeN3f9HCf):A-R?[O85\WD/W@+@#7U3:2G)-g
+a#DKFdK@<NM\cJB-G_>WP1RDH5S])eVN5I/XILNOC1aVIABgaS;a.0468d?T>eF
YbBJJcITICd02OI=NR-_bb]?]Cf72)?\NcLSPGEEJ@S]RVK&3U,@bYRF6dQ5M7MO
1QCW#^L66TfUP0=Ma/31)NWI-E9O[ONK4cR\D#-dI5EbDJNBUDZ<@@^@_:;dbd^@
f5&bB0US766C>K.T[&c9.Y@VKbO37.LIV5]a1P8\G0+^W(D;d@;7#<MJ?_T7b0NJ
8YA20>Z1W<Of(2JUY7RQ)#Ef@KW3?TGEPDX4(3EJ#S6DZ<2c9Q+[^&9ORA5,HH1C
3ZcQFRT-e94a:.2Q10C5][J[E4IZN3&T:6A+G7U#SSDf3CQ^>-M->YX9[0N/geVD
R21@O34V)W68+_+HSeedH(fYRgN,d^<\Y8?[WMQ+N;FO;W3#fU_L#gD<C24KWY6Z
cMW2Ga91IJX>.Hg0e<]]S8Md\P3(K/-P(]//&:/eM-+=c:eWa=:,_S_?g5+P(G8W
4;7B+QC&940=b<)1bN#7/+DQfJO#>NS5F.U4[K13WHg24,M,U5-[fL[])JgeLC@3
Z6S@IV;=45>44c>AV39Jc5SKBB>7XJW@PUM8T3-/LYYAQN49,>XH4M9Qa54C_7,@
Jb2B<VTB-ALU:fV09BF(-;GONMeKJ=^Z--a?:@HbE=G#<e^6S^=YMN&Cb3Xa\W;A
;_DEBR3Y7P6cWc)K;;a1M9-^@=]?OH:2UFLJO_)7;?,BLOD1\)^I/_&c2;U(3.BD
a?7@c^fFV(,OXPE0&MZ#H]aM5,K<)N&AF+\)E[-?B47KNd&=3H_Y@H#6V+6;bBK7
89[9G>P64>Gd0cEB&V\6/GS8MY+UDL(G0ISdIEU9g<298<\NJ2;]I??TDeS=9b)a
.8)4S<\VEJ>_#5-1#K]f9XI(#J5].fV67J]\P7))+EXIY3R#&e&D(JKc33LBMIA<
=V,9c2GbQLVYb.KHN<^7YYTGC<PI-.CCWS:X2;3K-]SRZcT@61Q0A,4XLb9_^K7-
CD.J]/ELXRT.Q^\O2.&Z5WM(,JS.U#c\EN84&4,LHX4L=L/#b,HM:gJ(c9S<Q/J]
P2Z3>C6fg:NLJ/5]]C+G8N2;Qd?<-N0ZO:U3T8TcGG_5M=<ccO\FU.,?O&Y#b=E0
>8g>:caVR?6QX8=S?7M\;4&UK7<^g<25Hb/93AZGPAFY#WVPHC-[[7Ac4CM38CAS
2Y:((KMa^]GTGA;080N-1fY/[FAe:2GQe9L<>d.ebe,WbEf;-V,dQ0c[S_:Of[^\
HdP#O/:S\[3bXQP1c&)ML&.#IIC3+:L]\AX6:M7IdK/@?X\aD-9de<17,6J:+(5R
1YL+3:(ZPR@ZZE5EAL+J?f_:GBHU/e.=7Ve#Wf0PWOa/H_K7\]EXb9]Z8UWNT6b2
USO5XRV+I<DUE+:P.GKb)Y(9;?e>KRd;a,6^:8?.ZHGe2Q3#NdfcSL+Zc1_0SN+1
BR8?AdTLI,<4;Nfc.3=TeDFE^K>Ze]NF;90\UO3e\RD>YB.LKE>^bJJIX,)QN7fX
.bd:64MQDI.E?dLVQ8c5^IYgH_)I,fE<#WIR#3Kg,DbILH>RVCLFXPK39(#KURR>
@:K3@4dJ)FV@Z1g;)g]L=\-+@83aR=a8VK2><b0S90P46D_V5+dF^bPb<SP\P7fR
Q>#I9=WV)&T9/<>cADBMN:1VNVW:eL<&_)YI=UO(_<Pg.+6TL4=C3d#6G)(fUNXY
EMTK==/ZBEX-BW8#ba.0a9J_1P5L05c4EL\3DeNgDB>1b#@)T/V+Y5?@+NU^bML>
bJ[9V8?8/S/F)::9M2;dU<JC36a(CP4IB(O-c#-Be1.BE^[)J&8Dc4KS.Lf,Q2;0
ecdM#bSZ3.<:B(cE7T;\E>DP-(=Z:&F^O+HG2Z-RE(/BI_Q<dP/)ggH03Gb5.M3g
BZD<[Hc.(d7]&66;YR3\f0+AR)A?CAg4?Z(/5-V?dO^R(R95W]N1SFM>X(f4a/3W
D(8=^ggV+E)/PM\1#+GD4/WT+acSS:YO^U3P>D#UX_UCBFU+..d^[:eP4XJ.#&_<
/.)TK\EQBd:g?fO3LC4Zg.;b&B+>_g0<)SB8GBK?L:BNXIK>W4K)N2U;FQB+:HZ3
GNN-7>550gHf;X?6T7J<:\-AF94I(Q8RUZIf/?N,\aH?c^dTR)HOd.HU9d[_f3AS
JD6XE;/)g<]N45K35IfG_c=b#ag&e>6OcI(feG,1?WWa:gZE6B8KeC+N:F.U4WPb
SHa/GOZT74@/P))@K;E_K#N:g3.+>^1>g=57ac5E_VOg^0IKDQ0B09KM6/)L):dX
[TWBf[,NOf[Y7IQ:#c^G4c+6INg,Y1QbD/81e9BM+#+e4KF\W5V72LFG3(M4(BFg
-3U-ZA/@c^Q(YUTTNSYJRN9dDMSa:?2cQFL)e4/.>O)85G:B0ZBSU8?2bZK>/IBb
c_X7c9ANd5^0I[Ya.5Y:)F8,VP99_Y74&9H0:,5J(LT38gL@bgTL?dK9B8DUS(]\
)H#@FX]\.O-TQEUIP(1gD[PQL<YI53gB4dPWg7aQ9^O_BID0COT0LIWC_U&V16K\
B^gWWC)ZT@42Se;](SP?7Z#T.b2/WJg=J0,8LS]cX;ZVAF-R9W1EV?F<eED-1/G=
WVAI>1<^E&e,Bg<M(;PZJ4YA93a>eUAeX;gI5#+L,A4F51NOA8XZ\QA?L3]eQVcd
;da0;;S#[-RB+]2ScVb_MLNF1G/?D=)eEGf^<@-@VTe:WcN(:G4\#ZEL8)_D):I1
R9RBQdef>8JGWH+-8I>Pb/UbgFNLOG:X\@\M9]DD#bZ9[LBN?PM=?+RM5SW@5&YY
,BH.JZPS2M:a#4+aGM2.1<D()?(=&KD<#?6JZ;^7,\:?)HLVOc6&Te..[<^]RK?=
9PU-I#\0c74<f85^\:TEdRgE7L_V5]RGD<YQ-cN,R9/=WO&4PJ67YX#BT6X3PDU+
K__S:b4Wc,c>Y2V+KKQ?DH.F1\f[fCKVcG#OM(c@G2YS=PTND;7H6bbZ;]R86&<(
&;W3QG=+4b,.F0?,;b8=:0XTKN88,L#HWa_AU^WSb:@O@2T:+IZa,X,VH;Q4OC5A
<dT)=3.Z&c+;8b+RB+.G\XT.E&E,IbJQgbd\>a7Ce5e[LZQI-M?+c2^1OPK9Cff.
+_O:VF^B^6;KZF8,_Y]0[-U\A2L-a2-;0L3D)UR>6&-J>WdP/KQ5fME7NR.d5T_.
T@<OI@,OOb3+6(&K[42:(P:)&\+([F+S#S.K9^E^6FecE8a;AH\=RPb(&>Z+Y_^(
YIOg/\KQ@RUYb;]\,K07FQ3AWL#PfP)N]d8@e0M6=Dd)T(VXO[1L5I3LGMF4ggJK
4Q-[_agTTNX4^KF)d?:^DK#7C7&-N6HL?8dbN]//]0.cGf>=;H(9f_&547&Tg:eR
0W[D_0:f#]c2N15330,DEJ@,)E]dIb4AG2b&VZ<,7<Jd\(Bf,5dA:9@U3G&F^8Kc
I/-KO6RB4e[?]2ME;E@1W<g>:^KgJ9QVQO0d37<.IHM^WESU\5G5+:ZF5PJPAVOR
dE9-?VS4.6NIb3b)-@SSLSQU:8@SSV3>.P?B-a\VZ4C<:4gDDZ?NAD<S-e?gJ-\D
P.-QFE7G0^6gS5XS(R24X7J^<\SVG6g/S;g>)&H^(.K;W,+N)g[EK:F\BPM6a]R?
BHL:1:DE_+.cD<N8,&<geU:bI(1ZQJb?<-aJ=--Na4;;fP=;3KL9,J96L/_L8MN-
,>=A3?@R1a4f/d56P@Y^EM-;ZeBW/21UT5.;Q^SDJ9S@2:W([,,P6]?e<fNe\YID
>)\]Q2f<;#+U_UB-bCZ96@=Oa7:(Ka7X_HBa.:f\FeJB:gRcY/X)RT,@FScEgA./
ZEW_,fca</aI@,ETLgEYCeR;IIP3&d^1@;<G1FXLOF(9b\9(#1OU6;8&V;4K+E?0
bR3J9+2S#5d-++&7.bK/9LJ2HP.0DNa-CMF>_)O-S5PR?3OZ&UB9B?dX:7.7(;Wf
ef)VVG@8&7QVcM.RMPaWJ=GT\S_J]A50X:LH;55_:Nfa);IAef4bDXR\2+eLcL/U
-ORZO(MWUV@_PbR[@J8_J18f<WaY6<dNL@LXX^cXG+)1f<9>I8(aac0KW4FVFS4^
+PTMQQ-Q0EdH)+)@&6..f,,TE^-gIH8=1W<31ed<9c(&A3U3W<?[7eaIASP.0(?-
\.aK6&XbQ7a.DH7fH/MI\NG?GG#I;9N(+A4Ee?392T;L9ER:VYHF;-FT9HI7CL8_
^6U)T#P6=0F9PVKc5c_(Y^DEN^QTgWCCbP/eU[7#W>M6?/;dP7J#2>MRCWYYP&;?
P?ea?#PJ3g:CaEREW8d5=d@:f9XEa3+Ze40P1DN+W^Db&a^fI;Pf&/:@D-CXBN<N
7+:JP4EM[D(#,@@Z75f=SXF4D49B>#]B:9O]7R6;3^AU#S#8B/XZ>]1U3HCB6DWX
,Ua\/Yc;(b4L^8c3_DQVSB@AKD?#U-O]PaXA[GV#O=]?P]9GFQ=-I\-TC<V+NE97
=K]7QSYJS9c^-2,fHBfgI1MH0AX#I-\P[G&H-(_O_WN_LG4g9<>a71&IF-HdH.V:
2O>FE^BW-@-@DZ208C_)Rc#,A22#V5MY(0IRQPRXZa3bW?DaGd4bCZI\#Ef18a^L
(cR.:9=8g5PG+0G[L]=W.IM>Na/[8BR]YRLeeO3O<]ga8FN4?[YCC#aceg=\,_N6
O@cBBX^LX0Ng]G;?\^:KZfT.EL4M,JWNe@D@]&B,@Y5Z,@&ZHG(^)TEG1;+-#LR3
/1W8O/11X7-eO&/NVMf2((-S9#U8.W,e9EVF<J\V)+,3(O.SND[N_D<#]5b)XPc?
7g63W]?KSE=BC@HYfL]??5)I]Ef;(@/X<61[]@cgV<1YdH..>J]MM:gdUF5;;TWB
ade]UaCJW24:a_G8WCTK8NE^TCTQ,;gDRTHF\;JK4,AW^O)KfQ@X+,g)TL6QgD9+
QW@:)0A^8e(W.;G/dHCBcP;FIO@.15>[&R1#0/Bc+;P)PW+VG.=3EcKF0LX>f,e)
^RCeMdEMe,=IfMeNZO>ZLNBR]/J77bSf\<W636Q>VJELI6a?#M</X.2276Pe2HEg
.(9;\<DN:=.<?M:;9(fK7>LCNA<T.7=+Tb(E(+8O/b[Q1\LO4?5TA)3<\>VG5aMD
g5KcU&H9e<;P^fF[-Q1<@_&;,#HC)R-6P5Ha7SH.R(H^e26@@(;O):g-5^A@1USF
,#5(YI.+Eg&B]Bc:8U1c@-Mc^[9/L54HH(a96&H>B#^?G1O&8a>Se0[1<M4ZE#5F
=;>U#GWd:Y2KCP#:H&KI5.QNWW6[>ef;[_DE?JefX_PNRAB,B@7=Q7c7TP:E]I\?
UCX]QBFS\]&<T>K?f3F_)D8CP(OHdI^1C8VD+0a98XE8]84c<0e=W:-3>QM7gKXY
/#TP/UE/Y=+#FSQEEEfDP3b3b5NK59?=,0:F+UL^<WX.K5ER7HQREaC&KBV1,<@]
8E(JBP@-M@9MIBK[VDLd75=ADID3BYL&H1LUT4#<TKT?>V-;L^f/4^]G?AHZ6O4T
;?a<NDXMFMT0C/[.M;&AZ&B)NY/PH>VR<[M:Ze./,E.93c07Ka-<+9F]\02@>cNg
V]gQAGc-9PA=BN2KTIN=R,G9<^1aR\GV5,2J-PNbTGB?H>\4Ng]U?B+D80d?eIK>
(.[2Q,c_a4G/bGTQT23JV).fP<8Abd(+@8fcbK_GXc^TaA2>UA9&X/Yd2BA1ORY8
G=b/g<]]@CfZbZQ8L1.Bf^HO32QZ4&D.GCR/W4.b(G-U36.Z:;/24(R5X&RL\DQ+
+]]\>U\<V:@:VPC5Q\@UTLL5<R)(a&^X#&#B+:\M?Z083L8@7#?)@\.3MWWb:D8\
V;..6=O;^NPN1:IL[VI_)9Q&MNQ\eAR07gRHMLVKBPKXN0HbYJLXbSR]+CV#>?5d
D]bXCH[8G=#1+YXLM]HFF;J,,?ZOK6N8>,A,3E=<gMDZ+C2,U^/N<eaA_,ZaafXK
(gdDRY>KY6&SQMaI]3XU,UR_.L#XYZ.FCZ8V:H<ZR=<;),502VE:g[B40WF+a1&N
11-3G.eK9;,WKgIU07JBIRX_V,.J8L-d:TM21c9d\V:@6fX;Re95]=PDF/=QIdQf
f<f+XBFW\C[_?,4<6K;:K&gU02X>P3Y:Re-^2bHAMDI,d4]O4,9C/;X6gY[M&dXX
:X>?L9Y(c#f1Ra-^[g,A_KR8+CBdb5]+6:(LOf-UTQB14H\.E)+&ae)_YK5W=dJT
;aYb&cWR\C\+VD2T\_Q=;c;=1gM_SFL=,c@9++X/CB(fGJ]8?N[_>TEgN.;GZ2?c
YBN(7aC1>Sd9a8EDg?0?OGE]I-AX;E5H,8&[aMT@G/?_KHBK(D@/<:J2f09d54+]
a,e5)I2DPSeK/aQ\40JdK:(@PZGgN>d[8OCH;2WVc.?f](ff(f(aK8.0=6NE)214
-FF;\<)d1=W0]HKE3K_EEJHM6AL#T#QPN?,Sa&-F)K.JK=+]TN[^(F_-4-#+:FE+
_/A1H;Wg/Ja2U=N5C>6^8IAXE(PIcAOY]P-MZ[ge<B7W_@MRKC\-M#7#+JL6I[VJ
A7\YA26@I1eaQNeAdaTf2]2b9fO<C4[RN#[<2;gKZ<@7J[=>TU3#1gd9TcV2Q,aI
AZOZ41XROB#3MG1W8b#0g1UV^CXISU>&CXF\YHB3^Y<MGZa),f:)U)<JDR),_P_W
:V(L(f.P;BT93?d.7@X_QIeJH?+F2<Xa7)WP4(P7d[U>N9@:;D#4cdV6VC6/CPGI
:2cD^=fAIFGJX.7K\2-6TAd67;aP=RHH31DBR8+bQQXK<28Ld2-2\4V&S6(VJL,X
b)QWD3X)L7DE2-VYY_M\+;J)Y3T?>f_Z.cVT>#Zga4>[[J;8>I,.UAML0Ke,b417
XUQL+R(<gf8Z@1DKI0C79QU^R0XIGO5eWTdBa&]@?>He#5/W&N?[[21[36C-86DI
G>Z]?4,=6U1O[U0Mb#C@F,g<G&?:e];\B;\-V7.1VA^)\F][6WMd\H6d2>FI4A=V
\O1^+N=7]QEH)Y9)Q:N>YC6@VNYL,27?]_)#9gSS^aDIHR([eD)3bc9Q:1)a+I)+
[Ve12^CU>X>VW256[-.WYCO-7Hc<_;Q.Z_&[@79a>CAJe7VHSHA?M#P3<(fL\9]b
bM@QIG;LHa58Z]@G;2^JUH#PGEbg_^d:BfIL]2WIQ&f#eWf9O_)]/f(dcK\#VdND
.O?>N0NH=P=O,84M;If]#S(>Uc-)(FTeCd6ARVAL0XLY]1DfH=SL9C/3BW(dgZJ&
b+\FMS:QOdYS1[S?D;/a?[_+eS^849GEHJSZ&_cgQ&_f3]NKK\IBC\[F@[Mc[-&7
MZ6]R1d6DCddC)SF33W.0MaCIL8SJfKa&>WV6G,:/9ccVN1E(I1.cG<)b_4==:S&
g=E5_IFC?aBgDL\S,Y5UT6R]2;-]a3D9(..F7FbLJLN===f@P<.d7Mff8>J^:\9H
V0adFaGO]G>G-c_c5cWT[&eA/]M&A2FZSZT::&MaM[FDOEKF:-^c>J72/G]-_Q(^
B\V,D#QRNP;Y>e]-A&A+N&#,f\b5,CO&Pa\RIUGWDgcD](;a_B=2I8)/KW/bZQX/
XX(VG^NC.eE).V6d)@@WQ1DV20=;c)K-d^O>]T/_-GE>fc^fXd(97R4+JRWD]#)&
RKT,=@[,TO8KS,9fVBMe[Og9f^ES5ZYa.EQ=(H2eX[3Z,Vf[&XYg&:/SLR#1?&>?
ff_7#4A_3CCMV(8I;&<F@C>A9eCDDT[IM^S_\?<9WgLE=,8K]a.e9)XdCM.3f:XS
dEecEL&3=6I9Ig;=D7-c15Bg8[CT]7</7b_KB+1O<eA[XBc79P=,1TNBK2d9?8SU
WE)QKEN7ZD:.J.CQLDE8T6N3<Y_B+6S-bM5UB2&U0B<a@WB>BEeRfa-,ZdXgI//>
T8_:AKGDNRS<5VU]N^g9)9ZJcf\3/NU^OSgG+Pf\)40C4I#[I9W4_\OX-3GT7+c:
dDCRK8AX?=JX<G)<B.1Q@I-aZ0dD-IY?5c<1cGKYD>b?(ZUJ7/b(OTG(YY<AdQT+
>MF(bcfeY[dfQGX3J=>D/>E&bc8c)aZCdI1Q[agRK=g[<S)&cJF3/d7AEG)(MS?0
e>FXB9^fcO2R->^>:FG_,4;=aANX3(.eOZ[FCU#[=,6e<@#?<JR0\@8Y>>#--W=-
a&/VWB4^_OO33BY2FfA\7/U6@8CV41\TD[X>-2?/^a+]f;+:4(>I;9f8WL2#b#P4
=@cY26;@dKVM(7=G6@^Vd)(F3K4P]^=K_JV,R.\@GR8P>A:-_5+59B>?gUbZ?eYB
+ZAHHABb:E[)7Xd8/G\MGU09gc#O_K)I,4.DJ<Jg.4]3Da/)3C\=5,;1(EdM.J2<
,AE&O-Y9GT#AMK5OK>58d_B=40\8Z,J^8SHB:dCUD_N6>cKD\C-L(UdY3506AcKM
X\WE0)Cfa:-4cQB.MI4(E[:Q36@g<K\28DOX91\IOX3<O/T0)TaLIL;9H8bEHCL<
]OI\J,LSS.9V_ZgK]/2[1fBO9YTWV;a3]6G:[G=e4DF[O9/&H=MF\+1[gXLVbJe+
VGX@./(VgG4=2UY(f1E-6EfV:[@2ARZg^.;>9cOWU/EgV?:RHQ()59<@Tf/)<4TY
00X&-;F<^2E,<B#af\VUb0<(\AcE/2-0?EQ)8#4QLEUS\]O=@aFA53.)-4QWd4:<
>PG7c6aI0UN_2_f;JbWW,1^)cXT^@###EW;WPW<F7MWL^[cWCSKX\5.GAf3>WDAI
5UCLXSa<TVJbB\Z=-61=^8e>P^;HaC+@dCNU4-FJ)5IEJN&T:aA4#Y^YH+Nd)/<>
C]N.W5ff8-7B3WWg@SZY\;4X/#0c8XXNQEO2::Q>Y^feGDOfgHZ+:UN:H&VY4^aT
[e@0\&gL<3V&UPB>P@TA;WZCB&d)3BaA(J.R\Y#AMW)<Z=;<G^FUS\1Z,?.aP/\3
<GO:BJ?IFg1g<8#LI8JD_\M?5=(:b65J;bGWSBF^WN0-79V=ZX;4_.X,7?b0eDZa
gP1TEbSXLRD2-ZD2(U9eGD#N#\+9WU]+5YdMfL01-EYM06dG0^FN2Z4e\a8[P_FZ
0W/7N4g5T.b-aC75b]+LA+bd@-/<JV#4aF,IfHM@Z=ZNBPg\We\RUCc:,?dFAX)P
f6b3#-HZfYAI:2Z.Y?F\D[LEP10JHF-fZ:VX+]YKJd9;-U5TOBdR)_2^-.V_dfL^
;\V9<TIR=+M;5^2D6/Zg2g?#L+BFdcJ:[T\:/<--]AG]@]ePa:0?]6V@0SR;6dU>
750B>.VSF)GTXJW)NH?;=H,06e,K5b&E_SE#O3EFf3>[<).f9@@2=ZZM0PC,LKI\
?><a/V9,HK3+Hc\YB0@fI<-d#g[(#[8R)V8SfV<-T:]72ZJI<HfbR_],e.7Ra<Y,
.O?,CII5(4d6-IEJ.-&&VZ@I/69^F,@(MT#2@<N-JFWOcCN@8GV0J)fZb-G&fWTY
?P;?,Z16+FNG35XJ>A(;WOUf+18W;c?51bO,YGWQF<<b1gKS&0ONd2E71e@@gfX^
8-b>V8aaZ^-,+Lf)GJCF;(.J4K=XB#FMETN.UP(N>PE9K.0=<I^f<gT@N30,^+1B
f5_VR=R_(3<7-LHAa7:>GTWdLUU6gO)54-O7?1.F_9G+)O+]J9__Zf,H4=N/JN2&
eg)9OMS[HaP64[5II\J6@((>V[NW\Y(D?0&Y1+\[7Q/(4;,[<A7BPS_c6gOG)dQ>
=#?-#^1XP]]VLYC/3=BQe\R3E&XZNe;C^80WFW3N9+FOQ@#Jb0ggFQN:D@<5<X6X
-@0>&F]U<:=)H:&;XUb2FQCTA8(+Oe4g?MTVXB0Gc9&d8FWbD&7LS3S>CHULbgE\
WA/_?NJ10&Q9=2P,M\8Pc:Y@+<F7IH7P1YNGP]B=3WO[MDZOK(=W4>]#<J2Z5L/<
@(W0e[Z^Y@Q>U9+;<_<GJRUAAJ;HcC.?RI#C.=CbKJ9W?=9>E-9^XK+9c&+b_#0S
7Y-8-gI?dOQ+0]BAd?:JR9gYf]7?#5B/E[a#c\3_\gKX\fEN,=/#/Z88bf4S5-E?
T02C)E10SZ]ecS6T-W^3IC\5U,P?<Raf:_H@=2(adf)QO.RJM99Y+Sg:X&V#025#
=TU_g\T5[IOXCL9gB^)#C.2:V<QUUFg(-?VK<([V/TI(\,+8E?bE;ea&+RH/5C1#
PY<\M/3Z=8,WX_IK&[&X<aEe,&FID?@Qb@5ZB>0PS-:\.&@F6H)]1UCR[0S+/GFH
e#)O5TTT?AF?:U_W1.c.,bU_aRAg_e&\;b3+_SQ9ANL5UBea7=6.7SIB;J,G-\.+
Hgc&(G#GfREAY=ZT=>7[c7Ne>:MT88T@0>.U_>S_O2UZ_66JgM&GX/Y>F19A6gd6
fd-,2B+Q^-Ib[G\E3R1#DH6,<6&.+N&cfZ@1OU0E^ddM9Ec22?..6a=QP;DO?6?N
R1-Z;f.ALIMZg=T/0Q+-\X;(.cHd&AX9GI<?AIO]HL1bCg]X6VMS]P6#A14)^b(:
bfFO[+7W523X^=VRb_1e>db4:dJg5R0_V+K>O_deW[<.g57,CY?g3f53c(DUCV=B
<]^CgI2I2\B-2N)P?P9G=DQW:?276Pc7VJ13f@WN0R_)f\J;:XZIGG#LOKN=RRbb
@I@HNK4<J@fNF[N<3J8DYIX/403X/cA,;MgZXGb421_gIUSG=22db9dcUL&@69GC
fEPAVdH1aLgdaX-8\:ege,(S-26P@,_f8PX]K#NKO/G\Z9@(5TZQCYK;4T,8KE<A
[-@;\HZ6dJIg_<<R7D7c49+1TD2QK&VEN-=S;XOWdRU.;FL+&cK?-()cE/a0D::U
__+eS#acZ_)=[[UIYEMac=PUMI>FU@d&d.AGVW5PdBe^V;#P1IH3@,)A#>0Ybbag
=ECB2R:BYB50>I\/HME3b-Dc7AFCTH5?R;VPHV#H3Fb(WZ#74R2T:/fY?W<_9:X4
]3afKcb\cYIGe4,Ie4:WCU>@KK[<1O[>\K+4/I5XYD8=:@[M[OO)MQVOQ1F]^eN)
Y+[KE0g-(X_<\2KUEXJ&a\Q\]UVZ8EZ&JQ9AKA(B7KIF+^B9#VGM#QG&?Y(06JHG
I8H<S3,Aa1<X5cPL2@a45PB9WZ8^O><5)@?U;I]_]:(ARKJO2cQ4^g:D(GVQ)aI(
XGN3JLR:Ve9&+/;+0@3/PVZcD>S6KF0F9A3d&G<)5<^Lb2,b\&MM;-_^3@;3>ZO^
-G392G:K:QXU:?;>H6[0GHDI4Z?dGZ&Q?8bGcg:5B&-C>>EQQQaNE#->>Af--S][
cH7D+[;EP\8,,f0/?5H0<@NKN?PP_49Vbb^2PPG4K9eL0:^ER8T,?<GAb\K9@863
^@;A-8-a_EaDB8.#Hbdg]I)_\/JTH2UEA2]fRRb/[R-1_;;_8@bBdN/HF>+6TZf2
3MGeV?,53d_KZ;Da:]EbHC@-/<#YL40>))d0+N@OXUPBSgASC&L[J#d&IMYZD,DH
Y@)4.a?E9-7&5Pa:]Z^T+#f2IWM/>[2(fT&._T29Z)J(X[7]\]e5R_4,&;US((8c
^>29DMTSSM2GJ_137d;#^dU]\dS>]6#T?Q5DICS(@P^c._-OUAd;YUQ7cAbCQ^-E
B2F_G?AEa]XW]YXBCUC3Q3?+\cWM7+=&ON)g#S5]NS17/Pd4Yd=2A@;AEg^EASV@
=3Y+;,T/8U..LgUL2[a2/&#YX]>6D<?<5XeD:3g<9]B&CIE9EUQ;[H&#(2=PNBY>
D.0:S,Y8]&,_a+V48]JQA>VScQ^,I,IUAVU2:&g_Y?X&F[YZFOV][?aaU+>:Q:8a
P;@cRAX[Ka(PP1>K3.J1\3SWdVW&UB]>U0E6(3bZU@740:Y]ec(R>?-8)?3(2:4&
E8W58a[-NZ0MZ]B5IN=N<GCLENbLf0&-a=0QCS\Ze)]@2[4+4aa+WO9f_a@WB[6V
UPNKJW&>VNA53bFR:T5GX,?N-Fc@eLGEcT^fH_=4-b#GL/>gfC.>-/gUS/H1b(7L
CK6ZUL4UUW>6f8XO-BV<\:W<F1->d8F<U>aZ3>3,HF9=DB+9WV63b0;T@^;#DR_(
6.6.927I3\(9IeEGLW=+;&VUV]eWaCY+V33Sb:+XHF#H6&Qf5A)G])+)588g9S4f
7#VL1)0)1bDg54\O9])MPWX9,>#WPQ_XO>E=-a7UPQ,a7]dc17HS:6OAb4&82/J.
b\Ib_F^IS[STE:b]=IabR44TW)JO@0>Kc@F+5aD>2?;7_C>?1._KPf+^>&:<B.Pb
CJg6QaCD?03/8W:RIW9(MB/714B5.4&2WG47BFQ7KD(FX>5=>]??3MRUURX8=57A
cT_db5?a)(eeE5#]dT[+2)XSV?4/@I9FJ.G]P[68H6V3a4@PZfBWdM<6,1Q\5]+Z
I40I9Q191G/b^3J_b</)PdW1FEKNK^RPOG_V<6G]2@Rb3];J;<O,F)87FXYBgfZR
6Z9FfKUR0Q/MceT]8])\2O,F[<.7KJ:@b7^Vac,6a0gD\+0.4\6)aT6[W8#bV?.@
U[c^CfZI;XUQ)JBZ/)(FBKOXLP/,CQV,-+9M?^&P0J;d&?g4VJ?540U>+;d/S(GH
;OKWdW-YE4?N#Z,4P,3\BbO4&cgTA,.cZA#):8f5b:09);gH=/A8G8JA81IHC>CG
Y\5^fSDWEf@&QCPgU+3\X3++,b=:f10Jf.SS2WC6gF-N1)8f31SK(2E+=+H=-5G5
4DEQB?3LO/(>HHbS&4^49NI:PYMG(YR=R]e=1_BX5dNIGZTKBIETb5EUaaU(AD<1
bHE0_KKC\2VTD4#L0F2)K6=B.P;4/(<G+\aN88AFC2cOJa-O(Xa7f\+DKBS/<c;B
UZ;55H,90MV;_gHEfC=S@W-L^)#T-UTRLW#^/PdHG)&)SLKg;R_>1-[RZKfQZ&/Q
81/,^1Se4C7bWBD3#Z4/d24e^-23GP0Pe48#@YHH8gY)^g6H^BS4b=aEJf)PKP+8
)Z8TZD:RW:@J@L>NeY>YS@aQO:+F>BcZYKC[7=QO9;M_,#T9aQPFZ,QVUV3[P2M_
W]HGf\b2WS\)e4,-P^:VQ1]BfI]D6H-?A]XSeX[]KQ6;VT8:H1;9VB3:P_TSH_PW
R7e\^/LM\\,AcY\a2M&A,eIX^0#IEDC2g(W78/^WY=#(a2-]Oe2WN6:\)5I;NNE4
9OdV-0NL?^)5NH-].?/?(A@LO.O4-066##^1F:3I1#aPZ7RB2>8EeOI2d.-?_8eX
H+L+.Z72JXE.Lc1Vc(bOTQML5&?d69H7Ka?J-\GOBLeIHXV\)]XKUc,C=JXAVbUg
YIP(FORAcKgOAV=WF7B[e#dF,dc0Kce-GG1ID0Og56=S+>V+;H]3UA[5BN:GI?gW
MNW7O_C+2BXb9G&DB&S?-U_X@EMaTN3><Mf./Cb3>];2a^Q5.8gf,cX@O4[S[A:&
M].a.4+FaAfIYL5,g/2g4-@AI87&CV^=BXSf&05.YF0+TYUDfZEA6e5GW3PfV-?)
f[X;#(&OYEN/;P:]/,#)((S8YAKN/Ibe.dM=6;4?gC:R,>OR.SG>b<A4,.KfCBX+
&f,:OEO_<)e6/LY)27>L>FJ7-4TWNE>a,/SA1/_FWb,@_XCFeSg5ZLaKXXMW\8SV
Kg:PK3::+eE6+QZ.HEJO>e/)bVaJ1eOE)g0aYNFL.+/fL:QQN=0#2@SZ7(S:DE?3
@e)V<FGJa/K&2]U>Y+3]VA,<e(278/-3.M0C((/-AGAd.+B&b1PD^T8WQ0I1F+,V
07MdW\g?=GV]P?Xb3SDAW1K4F1F#/ORGG#..=Gba1ZMBcbXL[eeJRY,#<L30G+3;
1gV@8AI(<7Y^e&:M;/[9FU,gR0_?_<^eJNX+AI4a;^9(Yc0K4S;<Ad#RT+TNXW@?
g8)aS)WEZRSg6c7/14BN?D[\ee7-UX8BQOS19GK4)JdgF\)BeKA2V6c6ER=B::7f
_K9CeIML.eE8-1W=P0IG2RION<K@I\Bf[NQ]=SVW>ZJW3cQ1>-<^@^bQE+K<R+2^
/W9Vc+D>FgX/#[[8)F\45)_]#Q3E<51,3OVcHD3(]U?C/a:TV]2Q>:@&T]&fbV;[
<]HKI^\8FP/IHR=&-c[<2H+c@=dMD:bLE.V50Y\(K86YIG<RM9E#YKZK5&RUA=]=
f07LLB>0NVQM1ReMRJFD+L_?OgQH0K[V]>D:M2c69-DgJ:@OMG:?Wa#>J)J8L249
U-^CJXX]N_GO#gg:9(a/DI5/1_)60C]1d:#d=Z<&3+aI#4F(QDf3H9)d24]63D27
712[>eN37W2FH;[D=O<bBEB=:EX6:K+_bdF-A>OS>Y&H1QQ\b\2_X)EJCf]14Re-
@@cFVJ,5cF#MD3LD\X&3gfP86FA.KAAHE6A[7QZM.+dBA(IW44&d383Yd#>&87A#
1=LZZb/E?M0/)A_;eb8f[)M93\YbQ5;B/-g:0<33V\D-+B&7;R7V#P?OPQIg)(,1
.\2Q#>R+G6KVMYT)1bc,/a+(A@Q-^:ID>_#>)=/:A2H</3e]>&4E>d)]dWVg/],]
570SN)/(:1ID(cK8egA-;,d(,b]a\D;OC:eJXW3Y4KTTa@>R3b26:IbCG5_^B;8I
)G?]/a>\YP0@c/>cM5>FgdN+9;LLg2WB7)aF#GZT13;#XJeT6;0LdX=/JK(99Z)A
I:<^FF<26YIP5F^IB<[S5TJabK.dQD9?50V7&:&&+S1;dGeZ:YJD/?gAH<K:&PI[
7K#f)XN+[aB::SWV.-;[:G1&A]cdR5c(ZZ_bHEOO7]9.9,cK+\F:2X-CN0fO]>Qg
JP(#Z1d+DD3fgb;BQPR<C._:X6IO()Jb1GR?=MK/SUP3e.4Y[,7(MS>^8gQG8TUB
JN+N^,ZY53W93NH#>Nd?9Sa584=[4YEZAI>+R^NN..^G3T?Nf:=@^Q&Q,X?76PZ9
\63IeL93-QSdHL?/2;_Uf_YR/B>I5Va/+6(dP0PM5L4>a3(JX4UH4UXZWNL,aN4G
4g#62Z3S2]@/7T?5DNAA/62_Ge:(5O#/9V;6())=\Z:SQK&__T#@RPT8cP<8g@+X
\S49LO&3_1+CRJ#6(eJ(Z^&F;SN^;8<B)ffPI_]IUDT,MfAPQUY;-d1VfXV;8N.[
Q\FYe)/^I\.ZUdg.FP3>:43^.T7Cc+>aX\BF=Z<2e\g0R[IeY8YSWSe-a8g.P53R
f]+(\UcAe#6g>X7R2M\5UVLCW?)1?4[MHT5B6GdA\c(gM_A14^,[,6e3eM4=?QEZ
)b0S<Oag0c=G\_^:-2_Zc:_G@^JLMWb/0@0?,bP>bD&:4f4=?N>WVQ<D,gBW/cHO
8QCOf9>CY[A;a,L0N9LS-7TX;5A0(fP9ZA0L(P+O+g:34KIP2e,2YQM_H.c,IWS3
J:GY.IaEW5\ZLH_7:8OJM8UHZ/OKdADJ6;aU3H4e?#+HUK)(e_)QdXMbX?DZ90FN
Q,Z+_&CeDNMY9BI8\TPTBN&XJP<ED/7P4ZO3e8&L(@9,62J)SIAcM,a-/))SW7?J
XKDg6T]JCJHKfd4f2Tg,@:AM;cNHX#7HKJFE(gOV\U<-<^22>D9HCLW^S^SdTD&G
R8cT8[P(BRFKNO_Z5@d#4JJ1A6CC#\gN71#QOV^D7XHT<,VF\>B[>V?9.cV5]^N1
.Ke2-U<L]c88gDVfSS-?_?6WSWd@=N8g8K/=5aK6^STWIb;(G6ac6S9Bf\6>,Rb;
K=63+cMc?3SZ5KJ(.7?/Z0c@DR#AUYgGY(=ID>L]9.GEUP+&36YbH>9Cf\BU5H;+
]XeD0C7VFBA&76)>BWRS7-\3[V<d^.;gIHF_9[?Beg;ceENBSWZVYfHP/ERGI</?
TR8CUP=-f1#R)XZY49^_7)0f+4eSBNYCR.UU0EHAdWEW]6eaFQ=J,9(-GE6T9V+U
Q\^M65S?7Z+c/f86&<P#6X:,L=+9093)+K(@50;P<])Y4:#5ZCN#V7I9bQ3)PV&5
T+Cc7ZMUP+66F=UL:]gZC_fN;)g,K36VZR(fbbJI<X8WM&OQ4F2L+;1P&5XQXRY<
,:\f2+DWB6J4:LY\P.^dN2_f([8cDT:3D=G2:1=:#WK0TFO,b4+DfEXX+16eI#GZ
;]?1W7B[AfI1C5Wa[deZbH4D]1/1;YR^])2GT>,-#A-],ZYL>[^_;Bd>@JR7E+,d
_P3bT3BFPJVAUJ39_P((F.U6S0^_4&PY8ZGB7=Ta681JQN=2Ad,TeAdDcNH[7IU=
_5_@f76,DdV)(A\Y(,bVg0EX@7^D\c(5JOK[6RBI-;g[QXO-=V>J4(Mg,]Wd1NBX
84dZEME.3JE,XF1XU#fK@CHVW:N>^HdQ+BM79B4EE7[N9M&@c9&8f#<R<Mf_fX;.
_LKba=?IMB4H7<C/d07M)L8O34?-^[XBX>9,gR2DLQ:AZK6Z)8DeQ=C@:UQH=0NA
2>Re,;@K(8BaKD>;ZePU<K22W12ZBU4c;_dG^,/A^Af-4,@Q,e/+0fQG8UYO]^YD
D4L+DU>V3.BR,TD5-=]XZG]bK=d4)+V:3SEfcaJH:XS-)JTM/D(3^#AeY#M8Y=G,
VSMKCRP(?DY#3aK?P0&D;G@VA45<b(FG?QK&)d\,A[#3VG(EdeU60J3L^44:g)-9
JMUEe?R#gRM_QZ92&[Q6&HDEYJ#+c=7JF>b6WA;[9a_RU^/aPN/:(^/bUg(,g0L8
]SaA1&?c,S4YPZA[/+J^8bR@?,b&PJ-;1[F?cEFX4cDCF;@)@)@J\A:FG.BN0:f@
.@#WIR(RcYKD]<M6R3V,cEJFI(V<REgF&g4X7Nc8_:L<IB^(a#&6K\XOb@[AUMP1
eb3YF-&EV_aUF\Q:>5FALLQ.&Y3#6WW3dNBA#8d_.LOceV;?RQ<3Z,=d?E(Y9Q1V
5\#,M?f[A8=<UAb18De)fRJL8F<C0&<?0960(BWU#Jc((dH](NULN);9@KB?>K/F
4JW[3@?CR>TAO+,S6fVRI+HX8K1gd5:M4?g,JJbF&b<gH6He4LA1XT.TKH(EWb5]
[Uc#T8dJZWgCaTR2EKTcfOf](9L-9BEJQ+1078N__:e6(\8G[+B_[fZE+.<1</B8
gISERc/?X9</1,.bCM4\DVAPS=(N4P,8=L^Q_.deUgbA:WIT4RM-Q--IZVB2&7;Y
GV4LJ6:,#@WFX.?ZYLGWWO6]H2\]dN.P0BPARVc1&E;T,VL7=#Q^#g#)[2R]S+YC
0#b6B(1DI-eRKM-6,RCN+L[[2P>]/?ac7c;A9XcS\:>#MT,XLaVOFQKdE03#)Rb<
C>E>IRXQ25L]FXB>P<A2FC^W-A8>VI>91/A>^/>LRATT:cWbAYa(>)L+MYL;+DGC
e@EV?;/R]+b:]-(B)AU.,b+,b6_XE7W[Gf--2:,33/Dg<STT8<D,U@EW[]C[)d,#
O5Z,a0bCefT=L6;-^a4##/#?)SK:S5-VL8?E^MCC&X1H9gK,2:f\c@fN?9G2;207
GD4R:V9T9DTJ(Zde5d;=4cE6PR0aWe<7RPIB4GT9_K;R?\W9KHV=V1HAS5SYDUfc
H>g7B1=815>WRPZ-@+c[A(\UN>PUWWI/R1gBa(df-5+8=UG29I7>NY@g\?7FX:5.
/QICBgd^C>\YaF_<L#^LW4TT#I>+CEG>#R;;?Z@f1MfXZW5b7W4fGUT?U80]V)>9
0@=d])0W><3X.CP(Y:cHLb<<=+]Y(OGMQeW9YSHT=W5:;@=7\XUO04f#fNK1TD3C
IgRSgIWYaYc=dVAELS/1AGI[\R#c0JA>6UgHM6V9Q[>;eSFI[U3)f)B?OSZPPW-M
g+0OR1Y+Ue[>;#IY:FEb:aCg\?4O;Cd()8MH?CCHZJMI;e2MK-4-dY8>TVL4Pd96
D]6G+:EC;Va2I1_(FYSfV<aO1_=4aK8<FD))^QOL3(1[X=Tb^/[^TR/a4K]?:T7&
AA2Q#Q0A)\1OFM+S>3?NB\[GF&Rb[U]])QGSG3NW:7a=e/&eQ=OO73HIIVaIY.KZ
aBV=@[/DU743-#G>P)P(3E)PbL1UAg&@:XLg9;O7d)L0;c5OUWZY@0dPULM-LM]#
M=Q>c@70aQGCbRfJWb_GT.Y-Q#G#UT^EPE=SG2+E[?ZBM0QIW^,Of)SU9X6+Y\P:
G/]bN]52c^\C51+;>PbgR)G-PaVZ\6_DM33G2:6;TbR#PII^M+(eXW^Z[DZDFULU
EKO_C72OO6&R[C_1)QWDJfd/_9:3#[H(H0;U]RbK+K:]GQ>=[gF@Qb&V.#:AECGP
Z/Z=Z)F[W<8[1)^&77LD_2P=4M@G?5cQ]TB_],Ta/Z?:QQROBC+0UeGZ0b;/,e,0
FXIa2Y.FSBU-@P7e/dVT<,.f<1K(?cC2ddMNU./^:5\eV)[f6=Y[5X^H(=eVOE7(
.Ef8+1]U0?1QK.JH##0M,=R2\g2dHBYT3Ud-#@1dS\#(S4SS[05>gBdfG+cZI?GX
J0OK4JRfe<NO3ASdT,g<_?_/60>PMK@H;60_-+d+X37Y+(:B.eceg1>J,^^g0aW+
9H@2I?N;C)2TP2MYKWR=6WF=[,YS5-F-U#3Zb&G:O-Hc_B2ORdCA098ZD.cC@.<6
CF>1I+cF-\Gb8H1b-9\2f9fXa3b/<]d,-T-B74=5.ZP&\<6b4/X@gaJW>XAgWPZ;
-]JG8OLQ#&X=GM7@4FD&&W]227c64@H:&2>R62_&]@;fBSSQ2H6M^7cf.3PXASf4
U23/[>#2#f[@2JUXQaJ6_Q_H/6X1OHVTL)aR])FIe0KXbHg7f06@=HUW:QfY)#a<
Z5_U(NCgE5EY+7PbNIA&Q]V^[?EAc0H3<\L+OgYd[>c5(LLcG0_LW--V[:[29O,V
8<NO,,>IYfdL9.YceV]+F]L1(H\aP)JKFNcV?dT:QD@c:PL>.^aTK#O6LG)4@WQ6
2f]LU+UC/C:.VS@0e0VYV5,UPWM?OIQ,;?AeY:Q3KSSN)b><7OV)_6V/-M38-#@U
.5.<cC8L<aWMI.+d(>TGO5C+U16?CDG_O6U5b0J(1Uc/L08KEQY+R<>5QV]Z4(&N
;(HV=\\5e)L^aW[Z9&M^e;ZA399;bUKc&(1&Rc,cDS.3S^99DW?L-(49^),OJ^O1
eX#CS;]ad>,[055:KMY5)&1\^E1F\6IED<-6VO?F@33P^U)US+?d5B07N3OELIeP
+=&^=?E&X_[:g6<f#:Ef)BPSH+#;KJ5DVJa5f]G75Md13^S7MP#d=.Q[:86PLBA-
BILYeO4YVNF;2=Y8H.OOcB.?VQG\6I#8(P^DQO)F?015abY>AA9=4?-)=F35e28Y
UD2M>@b#XH=]dgFQc/@#E[a[(Y5>>#OBB(7]@=YMF(ZbEOE^.aDf+3/67+^<6cbW
K=Q&G;3\HPgTad@G=)<V/.SOg\H<@G\(_:G_IE2cDL8L:TM_80?<@HS7I3?JSLV3
1S]R=T)??4\.9=86-aRXZ.;(UAgOM<1(M3f+&Y8=6aE&-K)ABM.TU&+ILEg<_J9_
;B3..>:8O-3e20I+1E1dFHF8F-MPO&^(0[NNQgcHQ].DU>7(3-F>/#L^bXY&I:K?
NIXST#VKMXcOfMX<FJI4&IAe=EbM9W9&JA&HE21g86N)Ia>>K8L^-5fDfI=)52X.
JZWX?#-S=BTF)-L.EF8W_M/d91?>AMb7)A&Qb>IYZ@;[PA;/QZ<G25UWR2-OF8-Q
R54E9LRJ>(=4a5(:Qe8FHB=JJRd<,]R;.MQTgQ27\(5e<g8W+LQUH9NH[+a7e6e?
ZSc>.]A?&.CaWN7f1J)?\5eD/D2b1g7PJUK;^N3L_LOV1&EY@OE3?-fHRPX6_VUX
&&eW8K)ZI6eZ&>Q7R0[XL6FS[HWg^O/<:@7cEPa:g1PASNgC#@dPXE>(1UR&/ZZ1
._1+=9K?>.T&FUA>K+Y_4/SN<8VR]GR_L2PU8PXNMN6=A[[.ZMI67:AB#5S52MBb
=T#BO12^87,d=#/0SJD8-C[.V:#KS[#R281SBD_BWeeOdX6#(5I18]?U:GPGXYJE
6;=Ub5#RE2UG?LAc.Hd5d[JL_:XVNY)3Db08)XM;ZFK4g88f./=@LKfJX4V<.]78
a8L1+A-+<Zcc(\Sa-_G^NK@@HC^PU4PPGW#36af(FM9[3g:DDPHKX9G_V;_EBEN]
+-4@B:2J;f-?KRRZQ#>f#@[1KC01LD346cXf<?/DR?-_V[bK&;NJOALeFbCSC4g[
S^.,#cQS_P5N:/NJ7_X(9NXY+f=YN,G<EXV-H[?-AS<^^(7O):TGJ]+2[8YdTZJ5
La/6TCR[IY48/#c,FFV_@e?54I749K-F^UQ]7gf0-<J3[T.3#fW1\[Pd\#&4B2;g
0;<3#JJXIU@>BHR?H(-Vb-1c1[<]d/X2e06-?-Xa)g;S0PJ5.83/OR?0ZX0>?UfY
5A2_(Y=DgdYAa\#T9gF.5>GR<0[KHAGA\a9Z]P4dQ[@CBI9CYXK&)cb[J^G2.A<.
;EA6W5&PIL@:&\@,SG#e7,A#Ua)G_+5G+#9Y05g?JSL2JS)\VgIQ5dGT]/T/XZaa
,QL&PT])J0VXHOe[[7,BVQJ])W;UO:TfO4)4&c_,5TJD4C0@#U>K\HY-V_)Q)&-;
#TO&1>65ND[+DHc)=&cWBH8LAfAR@=KEHfBK,QGW=7M3Ke=RXf^EPXaM6)bC\)d:
7:4]FT3N\L3^2f4B&U0[).&B(3D>UIc6cW>B3SJ)\Q@Y=[C4X]VUFV,SFPOM^4;\
FB&deFDf>3cIN>=Y7:DM>I9OHLOL209>5:<ER[Q?UBR8M#)b(JL,#0P67S[O73UG
EfXU?<GH=S0PO2FUf[[N4L)b[L7QY[G8ZI0eLC>GLFTdFL_a;+LOO4@1MTJB1WZ2
(C4+_K8<.cBMRJE-?LaDQf+;5P^J=F8PC?_PT6-PTISI[97E2e0A_8+c.BD7]J]3
5O<=X2cC.W#5NP7EE6E9I9PPZANa02]6Q+VGF/Q]2DFS8K:#CNHD+^)(.g94W<9e
=F&_eRXTZ/SV=ZV)DGEC.gJ[#=ZE8+(XKYM6=&CcPU<XO7aVTML@e<F=_3@_8R41
JQ6V&a\YFKK.TER;YC,dMXdBfdM33R[e2HLT731/EUfNCB>JS306bPETa\?OcC=&
KN9JK=S1fQC+_J^O_XcI:4GT4-Xcg+c,?R\R>]Xg@SXM^S7WTD61=>JCHT/OMYYa
ZVM:7]\WZ6]S@Ua\L=37WcC/:@YBJ_6SJDE^fXG4U=<\TEKH7,N6[_/eM]C</Y(f
W/feY\\#.Xa/.6Z?<M\750B=,9U.LMMc7f9JJZ&:JB+TX:?@D;b,CQ&O?=c;#.cA
e@R5a58\<@\5]>D4Z?B(0BR?6/FV(I37:d=d&gCEL@Q4_+FX^D]eaFN,U#3-F9X+
>dN?VXZ_[87Y5T_e9eT1geWAJGC0fT@9:gN8D630A,.b1:C29e=dJ_>3OPWIR]_I
g.V0YbA(>-T;)>NVAT^W75F]X/DMe/TRe7&4LT01RaYQ9gJO5RB<[OC<;cB/I^?@
KgD<3@.5]&6&GR=\TbA:H.Xdbfc7?KA@R#dT3,#4MX_.W(H=\H70NBSGV#ZdSdAV
e-;Q^;f9Ee?<_aS(e[TY3;U9I;=#,&ffCNBN_1TXNc6:7^1Z)fRZ2@6PFCcM2(fF
_/eL=9<gg+Ja01#-K<UC43\Gaccf>>W#/ALC1DEUPT)QRg[EO74OL[OJUY1U-GR9
5D97@N0J?,+a^cI97Pf\;)G9I;:6JAO/G2DG1e7N)1G^@4F/7Dg#+cK1._SFU5dL
:]]749&R;#PI2/6A8(ag5)7[8MPQ_.S@O&RQH<[0]SfZO?5B>.:GW5C[6c?Y[^3U
H;3=dHN49Q73&-KWbb6UgI2OIbc?Wb+9HOZYa^RgAT@RLD#F/P_HPO+E;FP:C-2\
c+1SI/5ZS<^\:,CXOFXZE\LSe02?T4,+796W)A@0NaP;N8T#(YbA013/HT5[-4Rc
VTP5K<I8TfI^G&+J;3,&81WCGQH^D(-1UTN22F[\PD=+-?3dJafdD]6B5@&RGHH7
GQ]G<<#;/EFMHWPfaeKI^Y7AWI[e#C0-ZQZ66]8MWEcOAL=U?S8C_LG@QBWM-gJ,
B3_<0EXA#AG.+bIdaRXbMde^20GH>,\<G)_^Gc:HCKX7>T\J[G)N6gP09Ie1T7RK
\,#7PDVPDCRON[T[Lg,>cDgNEGe>6D:dI)2W=AT[^,+d6-)WM[V(c]2B&W;)V3PS
?7f=4LEb.LTXcJ^KJMBMC2;Q)aU(.dUT#SICJW;bKGSCe6V1CBMB).?Fg-0fWZ6S
VEddC?c_-D_+\Pa<d,ZY-4=HB1;7[c\[6gg1]^U4C94-(=/7K:gEf,?Mb<L[AUV0
C,J)WH47,O@X/4d&C-RE6?W1OP^>EJZH4UJ2OB2U4V07U97=f6Q8&@R7NE3g8:&?
S&GBE#7X@=O^bRFS?b[5]10NY9+FHS_PcZ&5?eS.H3NLYa<LQ(Re=PY/#Jg^aU>(
F,ASSgA6;-/&:MdS6Q2J=LdgGFTW)3,^QTP)]P5M7MNV7Z60e+8H4OZOe&eSc0MI
0/D\^O_[)MVH4.eN;N,U+5X7\G41R_fObD#gGe^9bLHC\Ma.-Ke9g8(H\W>_G:;\
#4)J.bXg52W=J2AO0<I\_,NI1gSH-]Za=VF#S71X_3U-U:_=cQBXP?_62RaZ]P3Y
/d:,?<QD-E>,V^U1KFdMNJ&23#gD1#H;H;R3&+.PO-ZMg(B7?MV6:O-82>(T18(_
R)EM]HUO^<0f(Z7)1UGR+dd(S.g-;/>Z05?[8BD(7K+M&V=,SDFace[#?D6B19fR
DZX8IBF4eRU?A#O_XKgf#4+M>LMF3&(+XML&<d_=+JTD0X(=c_ee0@2TQ[V=MEb[
Vg]-AaZY:fRA<RY^d=;C,0K)<\;_GfB=K.L/KIe2b\_,)6+9[=X]\5.Xg2YD3VQJ
=9b#-,/P;YJ?2K51Ka9PcA?G)O3Q)6-_M<g+SS,f(Ufag2;HJ<7S,fbZIQY&6GE(
PX_d6=\2&QA#T9:QBcH=ILa]SW?H@-9/B>A)Q0SXBK)TeF;;PK,\&PFdP@=;-W&-
0d\^9<MI\e(]HDcC+@aDHE@\ZX^ABB\C4dCXg1_-#NKKXWdf8>H#>AE+FH0Lb#.L
CGaKOg.I4O#Bd^MI<e\>e)-8744DZ=1b?7\<Uf1;,WA)-IF)\NB/_X\b&>^KI#0Z
=9Xd;/2W9Y]QGR^5c&A54J@9.CZ]Z5@HJ=N(8FJ]+eCdR@5d@YUMWWJIP)WF)9W@
NaOOFNA;AbDAYeWR46TQ8#-&d8,N2+_\XRPWMG#O(O2-B8=K)>_>50<^YZ6L5O/Y
:d,^&T/KKWb;JRcB9Y^8:AZ5B,?3N?T38H@Z;L4N7Q-TWGF^>_0XgK[8=00ZBY>H
ASe[cT\K?YG\JA_KgcZUP=<BPNLVOOF0UE+(8=#V^,R93T,@eg^83/RbSGDG49W&
FH?;>W#9HXCD310FV>&VP(Ka@F;Bf>ZQ+K@BLVMR5Ve1=cWH@@[>(4(OF-[eWe3;
\(<:.LL[-/3D(#@@,#3U=&^N8?;.]C3]#TF)+]G0URfcZ#^<B83:;\2;XP+GA4F]
.8;(^Xf,V:2UO)9ZR;<O@3^R68[UFNDMV,/ad_[4N-T1B2XV>2aZ8fK]O<K]-QJ2
\?#;S7:Jaf)MC4BSFb2M,:JYX79R>84QWN7Q>?:O/X0>NKcADe,b]T2)N>]DfUE^
.7eR^PbL,9a4eB<84YdHV#Pg(62eUT;Vc9K?-aBEW>TA/7Z^45+JV\A(VgK?]1]d
N.0MVX/H-R+b22F>T@Bc@:[,)b<UCWZ7:4e1DOQ(J4gdUQA)(92LE2&>^\[XBaJJ
,I[9)6:7aNdM]+([0KF=06-@Q51H&1BB[bc&/]8O[)gHL=bcC2W31<fY;1054V#J
R&QRII/-e[+M)$
`endprotected


`protected
(S^AcUWO6&D(=8(VZR8(1Y1SO(M,eaWe(YJ7#bW1UL5M^BZYFA0K2)XK:>C[F=2c
d((7Nga(Z-6(,$
`endprotected

//vcs_lic_vip_protect
  `protected
)a9Y83VJ#6XY-7VHJ?;(<]V+U9>JZ\f:&@;Tg2O^3./^8V5?:>=Z1(#M?.7_g-+L
Y9/1W?/M@:O=d+(7g]CD=->+NaAFOR(.,<6[;3&eI8KRCfWHJ^GI\4g^(#RXW=cE
1aFQ[4c@9PPa5(R_Ife/;C7gNKA0c#eO<afEL8Q[P4d:Hb#2-&7^\BB@:R)L7>C5
;8G:\WbU(,?(S/7DGYa;15cgcce-ADEM#eL4.EDB9OE6,>9)[Vd^+\5fBW)N4PL-
X8],_,YS7ZAN#&F&R8\SPY+#V_7)7IIU>ZL-A.FOY.=&;94?F[D-9e_ZT.a?.;8&
E,CU.;2.L(>F-YKOGK4PIRNQDX<^8;>(GJIVRYJE_g78K+P5QaVXE4C.Y(3G2P^:
J,2,&P])T@71:RbRMd688K;_4;dg4TYN=?63-=P86;S@;<a4U.II13@0a_b#BDV/
]2#E9H#BW]3^9Y&X&),3e(IT0DOHc>MLMK>_:G)@G/=UeNS8>b-.K9cbRabZOH;f
(5SfEFZ@-DT7U4VL#6ZJF#:+8,c8J?0beN>L(H/EITNN]BV^_Q;a&f&CA>6@aeR2
74G0+K,T]M#3ZEcLZYg^7>Hd?317cEK;0gP,&ML6cHUTC]U[89E.]5[AUOP-0;f>
Q59VSN),1G/6W.Z_]8]-B3DN52[U@489Z9\U:5I6fQN9a<U)b?bN0XM=^_^:N<@5
<IJ9]8Q6-O72eEHbL:]?Td9+J>a_Zb5KX@+&;9e>(L0ZFdKJFZJ)O+7HMIb>M15g
:8/4<75DB[T5<ZMI-Ug+T)Bb84c/@:?;^\&M5WaY,8VR/CVL(R[QS:V94JI?\N1?
U,;_G)PMY<HaLQ_4bP:<48N5+4C8[G]_T3]=[J]F+b@-#2^T:]VG(dN(8dAQ<YF:
S=fEC\d+SFZY86-(8.BgZB;^R[KR/ETcI8G5\IDF5e-fJZ?D=c1]CTg[BVPI148<
D8J0<?AQ)S-B(?&([7JBNa&2_+bS53>c2(GJWJ43X>:B5F7b5@8C#VVB@XG4JcMe
JWSN34Kg^bKN7af2_X:3g4RNQX@M1)^]\7=RG#<7?X.T-3A82gQ>bLW-L(C2P4T1
@>P#9DHKG.b1GU,3NgJa7E85<a323?@ER[H?X6.P.]+eYE1WJBK+9P)_T=G@X:Z2
Tg\W\G:FFBBRMc:6B^:G2)d.Tf<HWGGV?Q@R8Z9f)U?:MM8OS#L1QW\HE0VU/\W2
Oe2bFF^?eFf0TJ;f]Qg3WFfYOB7=/PeF2R+S3Ec[6BIc>U?U[E9J+6a;Rb)C82c;
KfK:+&=.@)QM1/+QDHV=2g)fR.M^g@I(O8]TU8:<;PLN#]UPSJO(R[dQ6\:c\5Y7
N8QgQ[e=b_2;BM#3<b:]^V/=K?8_e\b(AQ+GPH+HIHMcXFgEU<8RWEFf?,#U:FEW
F+b-EQ5V&3=>e[EA/D\JP=_=b^Za&4MV>5J)JPA]@]7CFcK8RW^@FcWO;@QJ1=H_
\2-4K737+1WRDE.(:A3MN7T5PECcIc7/BHLdeNJ)]FQJA:d80QS_E(a3<a8ZE7GY
&0ZU7]R(Tf;a+SJ9&W?.)7^WR>&6W\VXNMT,cdfbd_8#[8JQb+FIgEI1.7^/[aP<
MV[-DcK@P,#>\aV5;aF(N^ZcB>)Z(Z23;M1@M6aRe,2Od93_B74IbPNP#9/?8BRg
c;9a[LfTR\,<dFJARDQY7BFQ4IU3&IeNV]&F)S1dLbKV.QD](/CaZY)C:I1P8VVJ
]-H/ZOJ?IX/J)7D&D3[7Q:aYOHD84C[;&_43\KID>-M-fef#9QQQ>c+KbeBT>&gE
Z+636:RbB-_/.?\G:IL>>7CTUBAO.(G3UI1UTP;1@G[<R]N?-XcL>:+L?#7c>ZgY
#@f,CD.?NPSe:J=#<5IJ.N<K59VA3GXffY&R?cXa361,Qg.L4Qfg,]cgb9Vc_9@3
F2>afTD>eV=gcF(,>]Q26O@N#B0d<bbZ/35Y3^&;fMf+T@eF+[9Be0dGg)4;gW-0
S1=M8WUbRE+O-0AS_,Ebg[,M;W:QA,84N=E4L#YPe)&[N[G88(P&G??.;J[GITM\
)HW#&[YC-C\D-+N2O.EY4UN#L:_\&I]7L)<CMf/U;3QYMdHAQ8<=dfT))4a.(=.\
,KA>9MU/G1G:IdW_7#-bD>a<BI.R:VH^NVgCH(\M3M&9DDX6a/3.#<H-BO?AP>D9
Za[ZbRXR@DS8#[EP,K)9-<b>62B@&YJ#5/6T5ABP8U]7J9_C:[.#=WaH#L+3bF@>
C1U_C8G,e;^00H46P#]OaJP2TZ(8<bF7_RRgV<A)2U3.<_\LN8ZY/:YUO#/Y/G)/
<SGGb^AQB3[ACUUGGHOY-F_b?=EL8gPTcQ8I@0;3@-9FGM8aSB/U]F&KFAF1LE.&
&AH(dQ0\_,8)=]Y0J^P<>M+JC(I\&2H0#3M)48#_&WH<8,T67c[B90:\CeT&&=8<
STT<.K?&9^1;f<\3#g@H?86\e:YB=^VH<N;FTE#;d;TEJX#+NOQ6Qdg?0Q<@OT_\
L,U,[W..E5bIZEXL1LG56b9>6)WYP:&4@5#R8,M>_e@b/TT(4++DDW[AJF-K-^]O
&LA8_SaR;K+de(45F).(F:#U&QHQ.WKD0eY=fa?O=G:1JK4MQ5Pb_2AEQ.TRdDNI
8b&&B]?Dg:Nd@g09eUgO<412[W02BLQU0ZZ1NN[9+0Q/6Wc9Cb2ANH6ULYVQ:.Z3
5R),XY(6<\\7+:\#G?PL\D3=d+TD1&^A_FREDV-GXg2OW,cU@]FDZ:OaLZ+[/OAD
>@+_#a]]MCOY9A6dBdO3@W(5HT>M;;WH0TGNS^#.C@FZ648HDNUE=MHCA@JWf>Xc
;+R#)W-[6IA<(G7cQUWLg6QDXb3/5/#g@,;aJW;fZ+S2T06[ZZ1<,I48&fG2IACU
.)^/&1F5g#,0+f45bWcMYe642MJAMCfYW&0Pbg)=WfDKI9QEK>]C##&L+g1U[(=a
aND&HPQ>T>0?O2a?eXY.b4J_X8,,N6fO,8]b/g4-V^[CT1/&/WGG-0_dL9>:+?bT
U4Q^+BVP[/XeWLS,-UI]\0DUI6=A)@9V:f^W4/L54(-W/T7#gWPJ?d;S&XA=[#4>
)#;19ZF\B5AeKU[^#e.V7g)DPB3f[00XaA-e2&^3TKL2=bYJ<3\c3IQ>>?V\##^4
d<cH7)CSH&22HS[a0;X=N6+O1KF032WR9Ye92[[X9Od_FcR9S509+9)H-SYeD;5N
38S;&XE5/B)aKQ[N8I,N14c-A6G)@R)aDLW0]-2BF:[aI@13WSR_Vb(Q)CE[(b=G
JLWE0U+N&M=eU8>JN-AbYKB_D/?L=0/e0=<)YNFKcfU-RNb(_<dS/;HLX#IPX4CA
QYH_>QF(V<\RXAOXa3#^N7Y6EWG^FIY)12\J))gd9\\[L-)gG&?H5WYbc_P+9?D@
X6E[TgVM1_g)9DB^)BO1]/?8CH,K-bK23:^0BL1Y=3D/d7ZX)ZS0C7cCTF.;3M\U
SX=_eK2<)>]2Ef_NUaEf0bZD,2a74@=a4.X.0>M:,aK;:Q5V4a+X(MBO,6SRd=N5
SbF,&aB=@(\+dBLWAVK@/XFO\O59SA3MO;:&X?1-8&N+-aaff?T5@8PaY+;CUEQY
RC#:,0ID=,TK_NUD6\]cVd:5#.F)P59g3>OLZSFYbC29./&]RE)@@9]-fbD7U>I&
1U-1F;I028[S+G+faV>_@2g,R;DQ8cZBX6;;A/B@Ngg[G&a&MRRe+,COH^H4U?G/
R(&[-&b()R3Y[#0_X,RB8=XC8dSL(#4GfHfbadVWT_aW<.b6@6)<8]Y66@L1&b/=
SAOc(;.Sef\&FT_3c]fbY]FGB3,VgeEgUZbV,MB0@2-b4>Xg8H(2M9Y?YKIeg:85
)[b[7NETUJ=7F417EPPC5E^XCd5WGG\NPBD8UeE&#^cbF$
`endprotected

`protected
#e=+UKB>&Pe2APQY:FW@7F<)1I2SL?XLcc^YFZc]D?5^<6MT&<,N3)7@4+T0QB2D
L@?Ae+f;6@Q2.$
`endprotected

//vcs_lic_vip_protect
  `protected
c>/TP1@5>Z^3BCV.Q8,02A;\9PCD3@SSAWV?e^/IC:bcg2-ID)[g((T]HDc#gK:3
SU^LKdA9TeH2gW861>Rf:=F>863\eLO2Bg>-fHeJ<GK(8=_685OU)eN8P9?>-L<W
b+VXUE[ZSWE#Aa:K5K<f(P>8^.&@RNa1?QR<&e^7=XffFTLZ8e],P87VJN]7Mb^6
G,#_<A;(FT:2AX9]bKK<LHbgPYd_dPa6LN9.D(K=(1CID[8S/e:KC6PKRP0XL)Md
R_GZ<A.7A8Q&ZW61<@/2/&-cG4)XROYd]_Z05^U+dcH)V/A>[bDW3:TMccXG51T6
=[-1([H^7]B-,U+N/1Q2M,\.TZYTfH+Y?Aa>SDVMMA#T2L].Q<ZUND:\1^;>L,ON
V.^K>BCD@a5+eRLTA;QK@_VGSAX4J<X&8dX8@O^4Za8D1KWHEcHS6Q_,R11,R2B_
Q?KTc0O/O;U)J5ScSE(4ZUXONdcLf\N:6.]&Ma:T(.D#PB3_V4ZaWV>>G>Hc?9MG
>J]ZQcF@3b:4_#9dRU-7H?RWeO(:g_=Z+05^DLKP;:>4&1>b;?G[cEXEN:c.=A>9
cLW:G\&TL[dAg2eONg0Wc/0KIb,d,\;[<,32gP#g889C[]IILI?YX@E+Y6Y]J;=[
F(bT64@4K&&QXbeUQ(FK+7\K5]HM[)OSO3^>DfI43@T3AF/\,Y\R7#@gG1BOP#O;
g&ccY[\S21Cab.^V/8Y6(M=S/HGAXQ.H-C@8I:OgBGD73</1R.J6NOSTXTL#>CA?
]XX3P3DRX+E-=-7=G/_ZJTf70Y2c\B1PF#[AJ3BQBRL9NPg#6b&?eGGQKE6>H]VR
4PT/C6N;M6]f6a<#9X_c4;^af[I@SZ0QeP#2:UD0)F3[ZTSbO@B_A-EXQ0dYbe:-
,6<D)O:K>Bd2b]9<N6E\aLL3EBW)U6S4\?:5I;-#S/VXcBNM6B#ePKROSM6/72>,
d6cLea&/E5J5MS\,G2;2Bf+b+g)^NJN^:-@XVe=8Y1PJOOD)_&Ae?M-JJ;?@-JH\
2748@KUYXdVYPLXU@\@GRPYa1IY6=9[dZ,P7.dZ9<\P5NG3<YaeGD0LD:_U7C.1R
gQ-DTH?+V9:B_J+D^/gbG:=:5FEO77CE^3;KS_^F-d1#Oa2fH</@<QKb\X53_e,J
[76FZC4:@@KVIPR7BLT/3-_DE1WRfNI72PU[+I>2XNcf=4DgF8847LS#fJ,e#gM0
;+EGZKPUDQ77LCE\>g+.39VeUPO-&Z1=O,YaP:\(]3XPIQ5TPSF>60>d)dZ;4\@C
LC^M4(8E4#QfDD##[(;,N&ad5]O>2G]/8DN<60U823KQU#M9>AATXA^>T4Y5#OcZ
+65U^J_&V6B(NV?,VY)206PTZFJ8L<9HO,Fc0gKbENP\P^_e5MFPP_SL3PA(P[-A
22F,gZ.<F=cN.F1ES?WI320?F-C=G3E,)/\_>6K7[3dUES=\I]daVGQ##->1QeP1
bLT6<133-5de8#X.+fE5]Z=0>2-ZU-(N1_>3:APCGc66WYC=bfLb2G_A2TKE+&N<
Z19]?\F-+J0S+SLeO;]4V()#1;O.X?P_YA.U.cQVD:C<E3e6YBYOKO&ZO1UORCAd
b:JUDR++WZQ#=A/ZLJUUMe2WA;W^VL#]7A_\YDGE]--\9bA3KR_QH,5PgR]c6&I1
b@//XRQFML<&PEKE.001/M(O?7Hb?ERYYdbfR9AQS)B@)7IRW@B(d]9DW9#af?c9
/UadCIBdG:[G,6HDIR>_RL/E77=RSf3Z9)V5&J8=9+U7,)KcF3<;a3Q^YK\Q_@QO
J8e;fg_]U>FCMA<S[ES\].DCfBU2QMN6EaNB8b.K3Q43I&dTHTa71=2B1F1U&+P_
UN@Z,\/953\a0eG[KZXS^aFR]@,S&K.@B:)fD<<OIPGe\^=b^LYLL;[TIR3a<d5[
g?:ANQG81Z,DUGE3Kc]OM>G1#QI2B#I9SOH?V[cJL>OQ3Mf0+7OUX<IR9La4I1#J
c3NSR)NJ7NA779JY(>H,.BC(Y_]W:8>9TIT^R\_gIBK_DbMD.T0GP-)TDM/-cA2D
Xa@VDeJN6/[c\M8N43,4IJ+-fNJdO>60e./K@WBdL]<XOK_2b-IBd-7.[E:YC&)W
?BP@ZO(2;IZGG)/eC@2>6^W@;?0cXHM?\X1D]e:P?2#ggO<+R-c=-Wb0/a5@FHW@
I,4F&?G#g_/B_EI8QV)11cE))E[_X;MYdRJ8O/S,d=ZCL0J,aQUT4\e\#-+A75)(
Q\[@b9H>Z(T;]6X>3BS,eL7X:(b0RH/&^,1Q0IJ]NXO>ZV&7)-^4cWL[CI3#1@IU
XdSEKME[+:=Z\c-O9ad4I8O^Z[:)EE@6G>N(g.A98P;BFDK2:0bMadSZUd;D.F>)
1:-65OKM^-,gbDcUT0DR;aY?3AUS@]Hd<0[W_,OIGF+W#DTF8g0:(,BT0[4=X&Ef
=ZY@1Kg:TX^IbC4d#KH+E@:g^M[D78EDV=A,TI-D.,U:ELA,#6HXE,9d=eDaPF&A
g+;A@)SUZNacP(IKIQCV[9:WQ4c\K5VZ[]?\<R)[/Fa.((c?c)8;<:^,V>AdW-&_
@3^0TOPUbR?9K?;XbaaU/L?(E#Wg4+\.22[CX6aD5WUf3>gB=@O(C3B]0<ZKA,4>
_]d[M48f\0YR3.b_/+Q5YBID[_8d0I<J#0]S9)K;aR622IdS[&ELX3P;GHG6IdZ6
f0JIa^;ZB0:&&ET)&05(XFa_@:C4MMCg.<O-6ZYG2Y:K<;F9Z2dXJfUg0U1.HF71
P9YX@@@e>(TZNX5;QL\YJ>[F<eV>D0W:&#GB9N\CYTZ<4-UcJ,VC7[G44WMZW340
)Z#Og[&S3e1+W\?\b@^FOQFG3#a[3B^-P(YH/;f#Y)1[3:;+4_^N@II^)X+0U8)b
dU8R#eK5.c]dG6@(JFRbZabNGa8(ceWB<6<cC=?J#TJ^&)BaF;f:g1b1L>O#AVUU
)UJW5JA5<A)2[V?J<+PcU]]<?)=R_HR[(WMUaDRaNT]=MS^4=RAQV\a4HHD[\SdC
PD@\.]+#&_SF&dD2KN.&\_,BZU<1OZ:==,W\XK>&JHb_:[IIVc]=&C(3CYTL8M3F
.83E><=PV75V_Cf2eZS:)..0e^F+?GJ#HYIcLQdZK,=2UNcFF><aN#Z()C3cW2X)
[+U6W#;QHfY4??->cE[8G.ZE7#]bKC>ZT:R]C(7E@\8Q30GKK=7N?d0U<e(g8A[8
8-NDENWb4&X-<N-#AV1&T(ZIUW0+P4R0CX?C3L2)H+JS_[R;CV_f=Vd1_K@e@LU6
YAF@T#UOM#RB\4S9,gXaLDeOf#gI6)XBKV/:U]RbDM@=_N#O#M-)/N1(<F[bSc[K
D-1#>>(A9R[+CKY@,AG]J/DW@UgMcFd)]@+a,89J^O4TS&X]UA3S=?6/==IfddYM
7&gZDe[W4&EWN-a?TCXe<(a7Q3L5<H,EG,dEcSA77^P/>^8-]>IX-fM)#XaN9U1P
aHfPPI3YGYX#-J(P^\2RK\f9F&Y],;#E/;9@OH8Cd:3JD-=-R>)0-3eF?fId,P_+
JPbeb?&LJTbIX_,Wb(3WN=?6-RF8GW9G<.Q^Bf^H]&P4^WJPA[3PRP>\(:.41ZFT
bb^J_^2fV-K\d967\YAHC+A+6_BN:0>W(I?)NS\U@e[XCZbZ1;aaa[Ca69H#U[^@
7UQ]e-B-06>:L69\X#^O&::X25P?:29&UCb=Q8Y/5f-@P:cTbT3#<4]VV4FTMI@@
)_C])b15#_LaOa;03J6>&6E&C__BQe2#^MSS?++1/L9a/E,&#Qd16^8,&+4JLI]@
e>NV,e^^bXd\O@D-b3H^Vgc#6:6S<EMEecB=I(^1V?#]cGf(3D<RIJHYF8g]0EKd
cD3],>dO(K/1c9-cc<1Jfff,B4H4XBSZO:(EJf6V92OWTB(^J.9N(W0K=c?B@1U_
dH.bIE:gAP4D>JDa&8W\>&,c/[W8/U)Ue,7L)YNIdgZX1//?N8J_?6CD@\3-.INP
UI;KZ>T[[(.g-#+MbDAOd7SSXT/XEE.9TEUQFSadA-4O=V=#d8Sgb_)aHTGAH_N,
,,6;fBSZUSRA\]GdQLTO#OK,F-V+AVRVL#9UGWDHcHL2J(-NBc4#JHRAd\dE0T1]
S&0@]gbdL]?A=6M:,\f].I7HK.a4987e=6c7#O#6D41)3?a>c58d>:8FBcQ4@dc-
aGGR^VFQDC(P8#gcU;2BQA3T9?QOPH]c:@#^UN_ff1<XVWB=:A0YA)5&HE0F^O0F
:T.8(Jf-TZ#bC_=Z1JS,3[4S)Wgg,:?RYOCG;&,1,HZ@ITWXfONFPK<0d2:2dG)K
DfH3_-P7(B(9NZ0P.WBUL55eQJZ,/eYa6X&;X+)I08>C+:.=B&0BZ=g=Q.G25g>V
/G2;bJC9Hbg@8dTg>FK]ILBge8F8FIQbcH)+BAZ]WKC;/>]:>6KeP5&UCEA.MfSK
Q_K:/GT@9X[gSZFCY^c7DDDRH.D)T2Q]R+dM)_(\Ab+bf6R],\=eYU-VeT::fG9d
1H#<RV7:Z1[Rd,QS1F,F&J3Hc8MAF:3<EE)TZBC&QGW2T^03MJLX83KUPK@C#GEb
.:.,62,(74TH@KQg.M6=+^?7/9QK:?[Lfc]\FMM4C#9g))-0K1[bEZ(HL1c8?K\-
a_PI^HE5@A59W]a&1[;(B<9.K12-W,:ZP:7-d6,G3^U1B&D<c4RSD6/=aR_1b8NR
GZ:A^0aN11+g[G@(RIbT&QM_L>2\/7]KU/LY#92b_S:OeMJK+cb+IYS-+Y952Zf7
T<4LTGfO)044<;+Z.ZS=DG/ED0f/+.;#,Ra2):4QS-ZgG9I=(HFL=<=VE16P?H.(
H?(8F\bG)/=gL34)d08Z>b\-M5E1\>];#==AUZY;_NCSYQDL<Y2MYE9_bEMJ015P
I&.3c=T:W7,\A3JNH@GQ1ORI&dJ^@:J&PA@O\66c>^fU#g&T\1.]8baX_23-L,9;
+WGaD-QLB&Y5XaRWO?c&c>E74\_db]F5DK8^9@]8eFD>e4/dE+D@Y.49<UXWaH@L
6TI#71AZLN/0e6XNWGS-80b)a>G_KQLG<QfXVH7)(26Sd8GWAPW/H>ea:J.7R_JP
)5.cd;USL(-G=g5\LHUD10M5U;#>]8>/,CBC^3e[#,7g,19XJM>J;[<=[QX9g(8&
a]HV[7@cF9@BC\CSV2\Og+S)FC@_f:DTHKO,6THbZU[WPgVZ=?-D[_>Z;@_VJ/_8
(_]SZ[>/L=G7_9S[-XNbAF<=Q@KSHWWY;FM6H,Gd<?V/K+;TgFf7K63_F[18B03F
I>6#SOA;N4[0\Gg(J^LN_XK^=D#@HQ&&L\,MQ,)K@NK/TZ;PUY8,WTd8GgG:.9JO
Q\V6BaM)>c/DA3AcM-XXSU^#L]gXWSF>M6BT/H9>H;^Z:NA:_W4M4Q[D8RYXERDP
B(=cE1=c1L/UM<]W4OaYLDK8/FR:e+a)8^8<P+/)/X36(0U17L(4>>6^VO>JBgDK
Tb&S&WLC3eH=D15NW,Z55:fI/,<NVOBfa7_)+AUIWE\_N1Y(D\QPVAZOU0bBagEV
d6[^SJUMPOH6[J1M\]P.9IEW\8,e>DD9&#KSY#7,&Ea4d_RQP.AeY\(VF/GBVc8B
9?ce)^E]dd:@61GMg,V<)<5HaU,?-:+f@>[YD)WLSA(^2IFM7VU\[C(DJ70]?\Yc
WO.Y+1>CZ[Y(KN9,b:S)BH;]I74(ZI#5)_HOI/+KE2FRR=@7GJBH(55=07&TEI5N
ZU6W_PA/7e.DHb^W[(4K562&DS0Z[.^&=9_#V3Z]J=g-B-)_gaI-&1L0@bc)EbBQ
/.UJZ&\VgKYU]6[R@/G_Y+0HH9NO9Q/f;.X<,KGE@5FHMa7RLD36R&gc<Aa2CY0P
GC9(/AI-3d]CZ<.))OR>c:-VUg/ed.aO/JCB9[IDVH(ONBa)/^:)5=ace28:O8da
L4PYOQQZGDDPQY.3)83(M.<Jf@A?0K7EKL/WA2N_<aHO2T@]:eVQ+.IK4AB8-1PU
U\G#)H7ZU?DB,?SQ<0?&TXJWMe)#?<3C\e_/6Zd.5RW#1\HDWIKU[S?)@;C>Me;f
CJ.G9YM#94d^MbS9g6[;fG\),S:K<U4&C;WK&AAff\T[\<7S;?9A#MJ4:02^bCXR
+\>MK<>).62gD,.-S&RDJW1YFeZb@F>#-<Z./YbE3.P5)M37402TW-I])RI+FE&\
\)>KKF<gQ.@gb,ZB::7>ED,THU)V@E4M+PVc6a&R+c3FBJ/J,\S=PKXZ[;&=\e&?
;a=@,O-;M7[OgY-A<=)Y_<5e0(-RD<Pd\a00CR6XJ[AM\DT;#M.?2MNTbL3RA/ff
0a<d#R@(Bb13MK>#QdQZBU>FRV-Y/ZM[^9HO</Pa>8>=O-9I.?N&OD,ICIb)/2W]
B#8[,M6@[XM,,XU>F=c1TN],IMY([f]RT4\M^b_A86cWgA6;^efddJ.@<.Pa5P+2
AQ;W+K+1d5VH;7M+ZS7MeSW8<U@HOD&g/SL1KdXQ8EL-g:;G\T48(e3X/E1^@LU)
\21^?9gTI-;P3,c^J_C6P?:gC[3F?[dN;b0BO<0O49QEcbK-25^dZKHTZf+VZT<4
g(;cHffN@d)&f_HBN9Q[]@Td_0QPEN\Y1/(fXQM1/1dK,f2gMRCAIY49f^DT=Q))
+M]@W-.W87&QH3;HfV6592K,ZaYRU_3J^(<QVHI40:_WW04Q^KP22eY)S+++;gNb
@(b]<C-G<NDDY<UTI3#:D>-93g&f#?DD-6bA@X^,Z3NG.@]/9+FW9SROSPaTP4GY
,e#1T+Y?QcT.L(V8R&/UE@QV,PQOH3_1V_0>SL;G8XbDUa^8PPM:Oe(BF,9HM3)0
-:0O]M^YV0Z@cUSc<D3#3I((f?1AQ\gJ-^OQF[b:e2;_+I30;_O_Y3OYT#2U_HR3
U8=2\RJ^B>>O1T5SJPJW_Pd@E2>;NYXR#OW)/fW4?J37<FQ7-=I#H0a9N9&=,YI9
2JXH09LG+SY@9aQRCN@0B@[6=EL=\/4N(:3_.R9-<c;T4(OcZ5AY?(/.&GC2R1M>
.Z.UK]J39@X---NV.0CLaKUN[OI)QaQ]7CI9AGF=?^3Bd3L/5X[f?19:J7aPdZ8H
JQLM0:M94\DG)PeF79BS((D])XU:YV4C^]cEO3a8&UXP>?9Q>AgeLfUGLE)I<;QA
RbFLdXV(S6)(ZHXE_D6X(X^-AL^IJdbeY<3SF02[0BMCFcA<D9-FF-ZeM2,dgFc&
cYe\QO?RRBD(aL]c>;MOUH?N+-3LHY2:EU#Na;3BK)TM6e@2:S5D\gcVNCJH1SGI
9/VWD76bVb(.R29KB#Q#+\E;eQ:H&FJS/)NQV]IOKQb2CRVbW3=R8FF,XS9B8d=J
W^]TP[e+,=[X)TM3V.\:72X[e&H+V6)b-Ac,/<?TYMB87Y).NA(@Yb0>a+MO6Hc:
Y.UCJ<S\?\:,DOeVQf^G</-Z;[V;37NG7?7-62]M-V.RADKMA8#_a=H8ZQd9[S7<
2R\E:I1FZeZ_P_8\O\+=V(##TaK>--<-0B^9&:)?&C+T2H:PW6))8:90I7[);&@M
TaF;:G9gK=F[a;[=a3-3PM>eM>Y1?aeR9KYQ[^-06]GdM/97M450MRY-<<]]H@P8
>9dP+D&^GaS&7RSK6bA3H,TY^UH7gcV4^EIDG@[@_\aa4Da]A=[SLM@BY5PX]+7_
UA9G<fK:=,[Bg[<[Q46PZ0R6H4S]Z[IHdY1Z6FM1(@ge1KQWdAVI-:#DGR#0OL)e
&Z-EG_QE<J;OQe&UB4e-#LTdfEEDB_VUSW^Ud6f(b\9O&,DM@_#,ORMf_c@32Y1N
9OVF=OOR<YgWCcd)WDGME@AQ)NSNfOC_+UdYR/5AN6fM1F&KCH#0X;4)Aa(4C/=W
?,9W961S)9UV)4@a(HOMHT28-G,HU0VGV0:f?Sg.@PDVH:)a9ca&1DC@d4a,f\9K
;6bAP<6Af(UO+e,ID.[5QY)7=&X161Q00Ef[:Y(BWaFR2,V;]WfVA-N&28gfM^(7
1/AI2R=_>eM3SB[fOe1[NUd#e3(B^L(V9BE1C@U/bT>QY=0HJQP<4_^1F7TCd^bV
XM2Q0V6Bg->5X&>7(4dfI#RdF++VB24ZW[BWX7E=AeY?.2aA(&R-[8NN>a+d35ad
MU?;FY;[7;72[f^aG,c8d:NAgc\UB\d=H4dWV5<FAAFd\R0B_R57P<[b54A&^)AJ
I[//,[Yc0_]P]C.G4,@&T&/7-Lfbf+aHUJD&RHZeK;8^LR@IJ=Jd;TR>NNbA4,94
2H,IVF)2:G:gHfN:WQ/gQ\:V\,Vc67ELAc0O=L:^,R-/9?MaY[05K:3SGK;CV9;M
b;@6FHT[Z53+&+MBFc0.>_LCKF2IMR74#3:HYa6UH>eD35;E_eRW?NB\1+6/_;Jb
6d6\XE8+AY&\e3aT6d4.WGQN)=VfN>M?BO:R#e?9^e_;<g0=BX=.>7&:KZ]4P:e-
RbTM[MeE92dA27#6WM?:Q&7C]=__(^c0?N6H?X7X3&T3S:45.dIB5\B/&?LF(Q&c
g@/(:YS2M<T#&-IR=T)a-1.WbWLDSJ]9a8T;9DeR)T]gYA)MBPP]D0(F\]+)SA.;
fH=MR&1J7EPNff&gHaYKZ?Q/eB&g)#]+?F(BQWIb_faWEJRUE.0EK9+\GP+36&D\
5bU4TT([N&T.5Q:Pc(@bH.9G\@4-G[E_8P?O2[8TSJJL_A#&5SYCV;bM/9K9Y4]_
ICXNbGXcXDP1^MQ=.^=P&b;A/cZI:<QZPF:^)9BFU+dG,:#?FG.Ta&@2V(^N\SG-
#3CY&DN@4.?1-$
`endprotected

`protected
P>a2&JAT^\@f2]^-J=0O0Hf8?S2GdXH3OLd,fDG?LOA3R+KDEeFO.)d@#H8HQ/XF
6&(^6Cf\^5Kf,$
`endprotected

//vcs_lic_vip_protect
  `protected
Bg\S9a.G:;6&Y+4I;C[?QSf)D5B00W^+Z/>;AOD+a,9KBY^VOH.7.(QL=>+>TUV<
Z;AQ0Z4NfEB7TQJcZ/>SPTO=adD@9b3X5KV0V9KV]UWaf;W_cE&#M:RVK507MC-T
;>C75&d[=aVNN6(<;PKXNIY]>69=HYdG+dR6dAX^?e3OD:dQ[-bDOaD1#ZQMXTCL
eY#D\&./&cQP1]KYBK7DSF3Bb419.[&BRBd_B0#SVGd;YF6V3d66;:N\[E+^54Wa
8cg2TaBJS4e-[_]cbe;Ye4U5dPJU.cdJ=8SF>fLgX/EPgdFLLM<B2e;WFX3g8BAF
6)GG\d/K5^32PLA])bF&@)DScX[[+dS>??C7cTP^G;ed8S=HD6HPWRe#T4U]M[D+
>YGb&G\_)9:VYdT2e/N-TU8^gQFf[aHHUBaSBD):GBZad9UD5R.W6>#][&7U[1PK
UH452dd<AB]=e9146Y,9B7S_#:1I7/f1G8^0T--@f/GHXQSeL)<OMf&;,#]-GA=g
e8?_11?R-XU:P;URW:)Oa2IDRWGD&3ISa_g2ZgS(KF.AFL@/_&d;+1MVN#W>&),@
HHN+3B0U@WY79T,LK^dDWXVe-T)bT2R4&[V[)F^VSH__X^:_8CN/5,/caHd<UDNX
C.55\2NaFg/79AgEJPK;T^O5UL)\1@75H=eT7N[JI<SVaRR0R<7XfCPO1E/I44CS
7dT+8ER,HDg5&3NWcW/6S_,)BZdQ&dTbPQHQ6MAd5LUH-3^#I_#0eVCeS4TM&SZK
Z1Y,7BL+HP578c[5/K=;&YJED4><G-a-6g_fQ3&b/&FK^^])AK58#JgR1bM#@,Xc
7/>2O:AAL:\,3e1P/BIYeO@TD^YB1c0./[3GffH=<COWN3:2RK+INfBJCHE0)B<B
K_b^f:O8TAN1VDN3fc2_:/?LaZ4H7G;-g&KHJL3fVG]](_;S9]KLUX9&M9#G2QfF
PPa@Oe(^eGJ+MJ?7eH.-WV;g&^/f=Y^Ab)dIYB1OQRNP;OZYgYV)IW4NH?LA>^(B
#QHgY.N.UbfP=eEFceQIX)eJ+]0_1R@_aODZf2d^/EdQ^L[(d[.E-0QN63RK6WM#
a&W(LgcPF<KX6CB.3-HLHb,?c-FJ5FG@X2EN@>6g(-H(fQ)_]J3D##OM8LYV4_.J
TI7M5P/-B#Q]=D2f2P)5K&(;XP^0D&MKTA6X<[\?cWGPeTQ?<B,3](bWXL@-BAN_
#JD82J4XK>V81,V3de2\\7)PJC&-J9WS,F&>TF/<\fT2g_3,<CXU(W)192VDcPK>
GG=K9G8=Wd6+MJ^bABAH>]F\RC3PD[<SO,28:E>J32^Wc#B&E(>&>@:Y84>G20LD
[H=7N(U6)gRPX+Mc.L;E#^Sd^3)e7T9)@JGO+.?:c[>8F=/S@#<D:gFD&;.@C[56
<NBRd-R@_1BE=.<)cc9bL[>9.FFW[5).&U0^[(5JTN2G5-P@b7gB+IJ[.VgX9^fE
HR\VEV)(\UYB9HZS_+2IE+M2HQ2T:BFRTBPXVW=V)+<^a/C05f,b417+9\9A_GQF
/GHCD2]f[KX@M8gg2F>g=R9+2P)K<XAc>8P#WN8NL=#Ke.H>=56b<DY&>A;\SVc^
]G^>]Lc@D>L@_6]Gf<5AQS^?e1N-GO982]TDM8>HQe;7H/P8V?A)=8XZ6=I9[])(
K2REP>(E(@_4UTH&=FCSO)IA<W).5/ecN(QeDMH<L;+XKg[gK)N[5E<V^-)1\4Ag
T#8T(eA0Ya;PO:8d<,KX&K487e2GgJ7-GDM_00b2XLI)5R:I/,f\\@a0:2BFJ2H8
PYQJA7-@-9;fP@1a\&0+;dA]agDYD2fLF1Q+C^:>S(3M:(L:CJIN?7.>c\#L28;O
N3O0W2#X9C,FaSE(VdH\(;F@P[3aeYbI-aUG^73L&^^H&-YU&GGX]7EK\);5ST]I
9VB&g^B8@Z,O=RNc.g@LX:HUCH[X]JF#510)8\G:<=9=)-e)J\0U3=,+RPeV&\K\
=E?W_g[ef8OU=J<?)E/+Q)SI)GTZ]3I<Y4X[U<2C6(dS-Z=#17FP\.+47Y/<6Z6:
TY^U7SN3Da]G)X7LK264f[QRY:c3EX4EDAAY2A.TEMOB9A?aA<RM@2@@CF85)=f0
<><G?+6F_(L(FC7I@+,PeW,T[K1H9dXS_.7<NFGEf;L[a,#7]?GVgQ+>;WUZD/cN
6HYQe18c[-&^MD<BaYMgHBBY&]a10(EM?7?EM9+.,e_0=f_+Z2Z:X491D0fJ@O6T
B::<FORU<Z[&0]:bVc9T<5@HMb)EbG36)4\QYJ0S,HUOgBM=L;g4@f&SS9JdEY4_
F8Z<d_43[4B7;?+EAF[RKTDD/YT27?Z+_GObOQW\-_)[d62/+YVUD]M+^5<JS]:O
@:U\Y[2UbNGA))cIFEYE2J=_b+IA/0U2POKD&@=eQSSS(=;[_;;\]&2SUU:I\b78
M2,ZOAQ?A.=CEPB+B<EK&QEEO]d=\bN=9HQ<DHZ>(0bVP.3.d([QgQe#SeG<&F#f
aLQ;/f:c5&a-3D0<7W>+IT.QM4P+W8T.Q=+KGY#;c1\bQ2dQX7);QGAV66<?91Q+
5Ra;=FEI(X)e;CE=B/;bTg)^)/-3&LgJcC7AE..4e=c.:MI,?3OU2EOZ=BCYDdbE
KG_<Y11_[U;3A]d&aI>>bcD)I?)0a3S#Md_D-Z?]CPJ4/VH8M1>[)0^(:a9cCa)&
X:5S;Qd>/EZ<41O0)LaS<OJB-QH3A#g@-MR5N:S4TMN5SNWBE]L_D8f(WHNA2T3Z
///+XA;;7WL(.eW&R1)eKZN7V=:-B?EOLfO#eb4R4CcaVO^cZMS)UT.;&H#O52;7
BP2ABf0S<AL?d;f/_G_L4(>JeN8\NQ:&/.fZFdcRYR_G./db^B2GD#Hd,PTJ;gO-
HKENBLVJ(FSOY5N6>Z@-B1a_?bG/,TAG^FI9ad#\OB]B(g#gc;f=#4&AAZ,MS-YY
B=]OW^WL<52&.+3;I:F68>Q3a#cK/@@K=<TNB?PF^EgJP33/,QeE+Z9a6>O8Q4#^
VaQbG6[K.?>E&-RW>;8GWGU#<@5;]6<LF2H,1.>:c#RD8JPIH)-X[9Ef1:7AIM)^
#efWM,Q^dRbOK#VKO8bMNE=U38O6/?FBXG:0TMA+[c3^U)ZK+:O:<\KF6QTCUK#0
4MJM=PV5-^8cJ&b8^HST09[2E(:>e,,N@W?O:[C.B(E]a0f6CPS+EQUNP89/1eQF
>f+)]=S:Q\6P)cYbE<KHSW1O2X8Z)P?aN/FD(4@IBH9e,+KU(,#E@/59O&;\8\LO
,:V7W)Y:9@HP4L^bVVgO^L\1^:@3KNR;[MD#Pa@&9J(gW^PJ4-Z/Ha[e:/8b1:0P
=8O,?TCe=:-&A9eY[>(&RB_(._Q]2+c48)8@D#JU3CU.Y/(QVOK<V+&;XPJW>aQ_
0Vg^?MR]W)^SeTRBUC#_^OE.IMY.;;aJ/B]KcSJTMP3K9CA+6^S&[AWECB@_dE4L
Q+EMX7FX,C,fY:QdR4JN_Rad;O=;93NSf5^94LVaU3:?AD\WR+BZ/[-\AJ8Q6?2V
](9.^C]PNb>;_VDYFJL3GB>C.;OW7H,9gQecXeU4a6-Jd0Ia55FdLgg\5PfeWTPd
@I6\?E1Ha>\BDVRM;<=Q5J\KBaJBbT(-Idd_XDg^#D4=3]#;7LI?1eV=@WVA;b63
LYS]ENWBURPW[9\.Z6>D]90[fZffOEJ1#MD;)A5X_7Q/g:ARW88X^,=^QSeO=+R^
TL[Ae,8642HF/Oa#LEB2b#RM:_R&03M.C>V\J;dfFV5N\W8J9[4DQUT<^0fUU=<,
XK<^6GBR_YVc4[FSX.W2cMH/__>A[KA+&BM[/BIb@7PQU1g+/3Y#eA#?=TQ+MW5,
0=7d;36..e7gS+acQT\[X/@_:06J3d#-[OAJCWL\HCf\LM1C@#EE/cT_CH]D4RBN
I_>[bW+8R18JUM)e0dP.OC/EH<D9+g)<E;91.?:?1EWV:I)eE(5[,=Z6^PSOSXT[
F:#;+c4SAb,0Q)=c:.5BcQRYXHN+bUeQfOc>GfE\N8^B:M2\D_/)]?Z,Xc2Z4;EL
/ZPU_^J1Tc60B7([+RfMSdXZP[>,B8+-Y/^R^7K]>&c</ILKHgT;]=b9O>;>QUf=
c:8)4FY5G^RTZV=@5IP<@Za6VVD\(XV8bb&58SNedO^6&egPbNJUO+b]3DS5f.2X
URRVZ1?=;5gf0]E:.>X]&#>G0Z,A0^N06WO74TDf[&4?0+BL0<9WBZfPSg(O?N;1
JXb=L=LB[X+X[=ODJGKP@7K^aK^VK.2E8>eR3DN/a4L:Dd/[3Z/1?)TU+&6V5^-I
PSEBJ4,I6HQK17<e3)a[T:a>E#-]4I4Qb.(@+ENOU&Ua5^PMc0<6EW1IJVN?WPV/
&RZ9W/8:7XOd6f;3,2^ee5OH5?28JY)5)Ge\HH,749cB<T-D[OM=;dDPKO;b\???
QOe+W<_/\.6Xd)2L]5R/9gWg^+NKd]DLDNRWO0&b_O7OU&I]8+2N)Y::Y[A2))]O
@-3ACM6R@TD]gL=J8_S-4.cPLAF8WR+4+9MP_9O>9.S<&e#4H_fgYQ([+^2EGL-c
,L#:T)=M/Pf0K(M86H8;Z7Ka@@U5R,fJU[Q[6-.J=IW<F$
`endprotected
          
`protected
IW\E#I]bV#CaQ1@>^4D/VQ/U):b;RRUc[5,f)LXTT_aV9f)>?AMX))8?>?C[CF,b
BIWTR5gY;EE+8DC;L(&aFH/U3$
`endprotected

//vcs_lic_vip_protect
  `protected
^;b]=B0E?/CK(>Y<,&PX2O5gU^=.?]><X4TXZg2[@a9>FU^>NVV#3(F/0,GWTZ.d
?JB7DOL?;^TTG&\\J4?Z/,>[&cJ#BM)[a9EbK-K:OD7D^AE2>]8bB\,A:OaafRE\
cW\-R6N5KIZE22E3Y5<(fF^a#+V=c0\F8eK+4^;\I^=W-,^WQY\f5O\F:W]-&NOZ
;:=BdHg=XNM8(V7G]4):/^<]aZ@\eV0Y[5,HJPEdO<FMEFfF&Z3NfXf:=\Q@aDS7
_B^JgYKZ_T2P8eLB#8TXG-8?HC((<@0A6EO.bJa1-IDH,=:^B+J7dZN-cd8J3E5R
L(IF[YeZI]-)RKb1Q12WMH^>F_4?XBCWU>@?]UBEE;J/\+T5G<5c(5J?/g)V:>9D
^>HV,N14KE?;]PMAA2&,3f;W_FYd)Z+d.d[9Q3[EIEN#^b12^.H2PAe7AE0;M][>
f6Z#.CCTY/O)9W#a,dafWPGM/ZgXFNZZa:1^4Fb5bQUCV_=[P+P:MD+5B=<6JBL8
_Y3:]Kd67H=2NK3Y5GE6LYf7M+J0IADV-6MdPDXgGB/LKbGQNM#U_K8SNgB87-75
d48EQ^NL:Hd:G-P/Jf<:+);5d(3NaQ&0;H\]=FE)@&KO#^>)fWJ:.aIAa]L,8EKF
e]USfQC8Bc@UP.9;-QQEESd57^G(4<=f#ce7aCC:aB?IMA;Y+8(fU+WCa1<[C3K6
3[LJ(AXLI4S9d^B6g=A?;JbXJKF#Pd0&3&ES.A(c:NE<FcU5G>M/]CUDR--D3WGA
0Z0FVcD;DHOA#+:93^?<K5_E3Y-4+V&O)f9Y5290Lf=,_^6+:)/J(N]:AcHZ[P#.
d]R=EHEf,+H)TaZ,MKNcMDT9C.8B\dIaUZ^^HT9JG\X-M@gC24JSM/gH-G7RY@H@
;&3a2B.WRTQ(R6OP371f=)8+eAE5I;<TN(fSGFdSZ8\9V65S@1@(DBX\\4[>ZQ&J
MWJ3L3W:@@V3VEVTc=HaEAC16e2ASE3[[U&MQ-M.e3.V]ZZ5,51b6A]QI3LN_]A=
EE<+U@<9YZEZ77HJ09LO0?@5]C(7\=X,LR8Be^V:I#=KRMNOS#Zf;dYLV,6;J&P:
HQ;<Z6URHf7LBNWQ4#[#QB)9._:A<87^J.)Q>dQ2;;-XfH/V=IK4QWBf?=\0E1_3
HI2eB(-PUc7aHTe(OC-dO-D\N=S<V5WcP@T/9\Ob-H-gQ-a^<E9.-?JPL.e^?dg)
^OZ+QNAb#7[e3Dg(##N>gO[5P<N99L1bF(NHGWBBSV+fG7RUH8ec)DP@A(?+[H:V
@EV84d.5T#5S5@6bbWXY;#_gZ.G7S3_/&M_=VD+IO4E2M1L\;Kd_H]]Z]4F+N36a
-RA?.[APZDG-G4IDX\))(J1\LDKQ+<8dP>>NQ21IO&?b&64</43I5F<a@45Ef(-#
5gc:g7?5B^,-K)gF(+fD^ef@=C+Y^F2g-+MD2NaGUNOF(@.+QF,SdXF?UXM^12IT
=I1EX.b+,,2J:/0_2](L-E(M-87Q:IQ-b\e)>EYBf(eHG+0,7&6c?/ON(Y-GRT;>
9P?gA8T[I]eFN)OMCB<dXgDM>+a)+J&R<_X<Ld([@G//C)2,+BMDC0+J@,BB<91J
W:\B:2[<9JUeK-2HCB1O2L)a.0&H/&7_:WKO-eL9:OaI::Y910.YL5EZOW)M@L[T
JCW@b#4L3UT3S/YU:_Z)J6.5eNLd]3^a@])^DfJEd].H8B@J8@F.Efaa0,&B(\T1
LWJcDT0H(^._I:,,IO5=5BGVDSPRaOO)CX;FZI_N8DB9OU^)aD+E-1;.M[92(b>F
4-<FgLVIYd>XSSLAS/A4TBF:0VdJ4^1;fE:eBQ)(\N\]d<P267R0\7ZZ,IC1Z;).
OSWRMX:7cDRK13_CMI5C]@9Eb8]Nd+0/L__bD72/\>TgbX.7D/NCIR7E0T[3-/?+
BVI?,5_LHLG;L=>0;09X<29EP/Z9_XRggWP@SH[^;RR^K0)b&VYR]/)?D##H(,C=
?^@F2L0FH8\^,SCcg:)16]D7SGF@@>#eJT/^\#_YO##.fYQ91#,F\?d?g-#][[ML
G3&1,-9779<[.JMfb8>6^>@UcBWXIa\9(ROW()VIUQ6c(Nce_]PTIB-<7C[:e<S,
9XO41g,P-ZJbC&6[fec#K6^5)@)V@>ZG/f__\51\H)a)4UWQWD[CJ@R6M/^)?QCL
4OAJ;2a=YDLJ^[:UB>X&(9#3,RUDbT\\J5ST=Z:I6I@cIGc)4:B7+Vc5).YA#_B-
H1^+]>Q#.dRG3M?We2#[c[\UM83NN?N+fQQDgUEOCSB4N&3W#=VJ.5cDZG4f=a;4
X>bO<+d(4R2=H6,>b:R;]dd@e&_.ND?PQAO/Tf7<bP=E]I0gfdG^9W0[IXdYSa\7
&89O<75Y.)HXgWZHI3WL1)2NCgX5I&C&<T^1V2<Yc2fUf7]f[5RXc70@XQ(.&Z8O
FdH4YJ^2(_]N\4F.<b?VSV8NRBQ?c_?_YN6EJ:0U(HN>C49NQCTJ]\O&g=J5\MH)
E#?J]Fg>6#9CC1,VYGZ/+Y>4+6+/U+(2>OMN@/;8PCc.f;\KgZagY0/cab+_73E#
#QDQ@d9J:dWb#XW4e93LH,MD5N=;P8W#JE;A+SM1WL4-CS4;&RARENd;+@TA9eN^
XfcD@@c?e:,QIAcF9]4.J27Mg+A?0a.4?/]O)2&FCg:@+EK,;Q;2(7A#RHCR@JE,
A4;\JNG;de5UZ.Q7J,:]KD-A9S:V_A=/0:N5[aW4CdM[dPMab\ZE=VfI^d[>X.If
YR7Q11N&>,8D7CE?KO60F^14WcIQU+SE7BSN?R6?)A6=HM<OH[JfAA?2(V_#C1LL
<O#KKAA?UM+PN[R4@Q^9?G4/J3>K=AL1(@G_=7ND2N>UCYCcK>6L8/TQ<#5RXVMS
+H@UPF#;,XRM\UXH6BE34TTEUNJbQbJNNB3_6^]8^f6g#/[G8T3<M(A))A+);FT0
B_,P>\._GIG1K&,L]8G:FQ<,g,KGE-J6>eC\Q4BM?7J3.RVSWJ&d&P]@a^K.79f)
KN><4Y9IXCWW<F2E&M12Eg,U93_--/dK)-+f;9&fKB:_FU;NTQ,Yf9OaW[F.TB#5
:.T1e/LU<5Bf4DW#d2#VH.KL,1(L^8Qb.1e_.GA_@<)NZVfU^A90MBMG0Ob1;<<H
\c-P2]CNX90Q,_(O)4N\&(d634K]<BIcHIH2Ee&B8<3_<\KVd+>/5Z-b31GYD.UP
._3d3O0]YS1fUNcIV=HNL?P(N_9?0<fSXUe3EE9G6-&,U<2->>YD;FF#E0<Lf:f(
>P8:O?EP30V8LJ5F#RN6WFIbLM@Q-H1A[0EQJ,@d@WOLV.)6IL5+3C^SW67_D>3W
Y3UVbR:I,ERc-/N2&EVcC4#.fCBJI8^)71DNB<(U21DB[FG.Bf0><Ba=4-S;e>-=
.9DfHCb,TL]B)46KKJJWLP;F5H92Mb?adL;0B]KgQBEe>d0QQ.DDFCFDc(+4?568
8I;d-^YVB4=g2SLP1@V+85-?/D2,@^)E&B)EJ3faW8PH5HOZ,gX^2(U/,W;HL]:<
EaN77@BXPGA[7&V#OK&d70;;#)S[LEEYO2c[NRY@K;-1a)D&ZC6G134(eV6#+8.8
Me3PaICF3.gW_GfX]e>NDS2F(C,Q-eO61T0.&5Ra>E//9A2K[DRaVf\+C2?Y^FJ-
4g&24g?3S(3T8@PO<-WMD\7#G=QKXa&6:O16c<bV[9LG+Z3;a#2L.>Z2H<Q;0)fC
FA_=#K:8:BLee+]47LWaR2Z:;&;=[aNFP8<Uf_ScF&6=f.@M?=dC4^:2WG6Q<>?a
c]/RYf[S=A1\[=:?OAc=RZg)O(aRe,AQG4+2IN1Q;42^B9KLO3QNP^76T&Q\c=GN
N5[8QJ:M7:5CA4g40C?3^)NJcRNTHONNS4:S4fC\\V0g0cN::6_.:3-ES6<-CX(T
(B+NK6YR1\d@BagP#fI&H>26Y8).0;aF/>Z0a@NJWA&-AB([#c::)IL=1@-#ZM&[
^7#-faGP5(1[d4SAgV2/bWMN52cKLOX:\_W)D3X[bJX:O+7LTbH/da]+B/eFC?14
9c>M@&-CO(YE9>:/UfMY)d,_9Y-+g#,U\Mb-+H;A_]\E<@.#[N3.G.7Z/2FJ&6cJ
@IZL4)UWJ;/NLANReTFFPJZ6c<14R:PZ#=156aP>79:00;F86^CcbU<,2_SFI5?b
P,a:U4IN)_=0NX.LOFVWBeBY611E@MZUH4/,1IV6P\NgGQ01=K20cPWT[EN+ZQ39
&Y,cafT-N@/QS7d4^#gF=U+?]).X)[:fCI?#e-7VB+5MFNC4;DcM4K3g;NNNNZX+
P-FK@@DSFdP;Pb\=Y3Q=-2S.fSU6Cd2YC^Wd4R]4@g4IA)J9;\g?U6X>VQF_CC6:
:[K,Ea#O\[f\EOSFC#5bY:eG7^.UfM3H@FaaU^?RLA+Xc-a-JA/7_c;>#@HOC->6
gX+&F,S0,e3d<&#?RI5_-N0Z&36D9;aPcFa7g:VIK\@eZ>g=XR\-eT[O[C5#BZC-
68dO9c5;O+:8P]X(X\U0f1LI-0+adR8P.TIcF^;/b#=Y/YB43fO^UN=dG9Q[1SJN
6OTO.02691bW41N):>Sc3(a]22?\F4/@5+8IaBRF08)VNTEYMT7Z#VB[6c(0eTeK
1K[88<]EW.KMeGeaJS+B-f_Id(@[)1V;03U]^4?4AD,d(eNJ;O9ST+Ja>L5Z#]3\
O?OFED&N,2cEbe.(#?[S(1e-(35PbNeMJX;b?+ZR,6?d@YbRI:JLfL@MSeYZ?\6(
[\W6A_-4^,&57/AULW;d2(7:fF<&7H<2e0gfKO-a-#d[XgRDBP9OPX<_a>JNMZ,Z
[UONV/<98PEI(5JSdJMH.#F2QY@T&-4VAdTXUK3agT+)Qe]?R2HZIa4#ILUZ?,:D
Q.[ERFY&MJN^68=\7#O1S[V>KV<P+aO#2\BVH,2;b3X44c78\D<#a\XJYF<>\G3O
94d+#@Qb@Wc;HAg<X0S2H6D]f6b+Q=d)L6D,8\372HD<;HX.DW8dFM()U@Af#IWP
PYDB_B)[E#<Jg?EG_cB:U5\5eF/C(W#/,f]WX_K+dO0I+#_QBg/Ea;?;MOYB=FQ3
-MD:EDX6fbQJ_5CGX;6O1(Z5I]-a@U\4e=8=6QL62g+=@GPf[X@A2_J(D:+.d;5;
V>b;aJ&Z.-1fXMMV##F@-_LA)R0/&;OA0Y,VMU?N.g>G-.^XBV,7>(22d)H\8QR.
F/WW.@ZF)OM\8aZW;G)=>bbQ+Wb1A-a=48a:C.[?d]_,C]@CM.g3&N2g+Z]I/7W3
@D9eWRWA(+g_AN?.8>Q-/8HBB(>bS@J>3]@C^,U7LX.fUU[\7-Nf,]^CE]9MU@9W
1=(VGGE[0[>)1e?:M33\IFKP/5(<7G,C4RdEF/f,&g<43<DDPO8UM&U.dQ^?1F@B
(dK#D@dcTNA>&OCV.?UEdO+..[CNSgLS/8d\&71+dgHLfUb.aF?W2?GR05V09;\X
K/eLTc=LEKRJ<WY0]P^KPYW3-Pf&GF>K[B#OY=:<^9LL1<8FeV<<YN,]KRQLFNI8
:W0[Y?2ZW5W^Q8[gX&]]dJ^DE]bE476N0]=45f539/dY0d]E)M<;+=D.N46U>G^;
a^3?&O+Q_dV8#S,<TbPWYTK:5cK(5E<WNS:\+UR+M(gcV.4(SJB<(NYPc#;\FL^T
:-Q=90L@8T9\1EN7g+/907NZ.=&]D\SZCGJD=H51,c<?YP=GdUCH_SZNF7X=BRd@
,2aA\G_(\fX)TD\3V\NG=Ecd=[48[JKaAO3Raa[H\JRH1cgD=EUagL\fI);J_<6V
R-T=A7CTFV:N:PNc(@OD_0:a@M8WKDaPZ\S67NAfZN?DIQ1Q9CZ7&(;;=IFA7Z0#
@3:+B_@e=IR8G+P#(V@3>C(OQF)(9K+18&TP5WU:&I9<P>U0cbMgSb-gRH&Zd^/X
K<3^_+T\TYeWO(F,[P/XWTI72JgRDQcFRJE9C&(NaLANL0ZQg9UYb[GKVe/c&f>/
[=1&EaSO0EKM]AU8/d(<^/UY,.E,Hf43CY;6Z8V7>8)(I.a&G7Pga/YTS.4c?d>.
>C]d_?3IT@AU#JN/B@80AGL76ZUMY,26dW<cV#=bOQA/KK8eOd-(_(];E0PB?6YU
L;21@5L\L5?R\;Y0FH<I9:9CR1-6ID#QQRO:>C-X4\TY8ffRFH:3Y74C,V-J^L\g
P>B)DBb8\9OD9+L6S==XEa:YDGIfJ6]_RQED@7>)JLfVAf-Mb+BR^/]CQ2--XR1.
Q(&>10-,TIU=2ZK_KdM2.68_TY.TDFPg>+P:X;Ua4QLUWQe:HN)eAW>ST:#46IS)
&AZR;Y9I8-HG8O7ZB9Wb42877(gY_RZ>;NUJX=bc4/V_VKgE7c>Z[=-35RGfRCL6
?XeM>&]f7)VBedD3,]Ye-O0@[PW)\4LM+LGGQ[O:W4--L]dC^C)a0VNEcYAd?:M<
/U?@\:5AE51VC3S_-LgYZa^GI[\NY[,U/G09F98/[eJQNEM=DgIXO]LG9_>UKe3C
BZ:e1+P(/X^VC&^Jf7#9[KU&0+:Ie=CO-MVaOM+[U.g?>Z\6_V?I;4.9EX2b0^\C
),WLURXW>FV5W-;--<Wd,F3R5b,HS=9C;=PF]fdU(^N9^QT#OP-U&fX::#WbY=)H
5^U@M.E[.c9>UF-<8&KTX)_(#JgZ?,_acOEHg/&5T6:&ITV;=#3W8aN#BL6S1OQ:
H@,FGF4+2]2KMJ@g1d#-fa=>)&UZdB0RD1^BB?\^NSWI8#-Z[AJQQ12J+D#CbGMc
B&SNNV=WPUV4;DV((:F<f.gBeX>+LUFH4d<J/7[KHAbcM2[=Be=A6M+JcCON55U(
:7a/:NF+2cK9f;;_A\OS[B5F?)Y[WL3@XY(^\JUQ,1#RIAb3+)PPD6\:dcH[L/U(
6]@;E#eQ-&T)\Ya:6;M3g^]V\>2aAG>eVB_-S-\T;5Fg41(1Z.E.KBS0/M&PT)2&
F(Z.RD1IG:6KJId=4[E:N=^(VP_O;X/BMI(/+::<:F.08R]6BYL@3R(411YP;T6-
9SL.X@EO52?L;9^D1^-ORR^gLN1SJU#U<@3/80\@XC\JgNa-FFdB7;(R]01bN,g\
WXgA-FV_/6DK=g^VCB]>+ZO_^,MH[[=DcNBEg6TW)fDH>G-21QSb;H&;OY:<@QPE
4JYFIb</3WbdI.feQE[==;0./?HN@S2FY]<P]FMf,XYNWZN\E2D.,QVF8XE(1[8F
F27#+KEK-08-9E7Y09=75>R;^b&K>^,\)>M:NZXbd/ML-YCB&aEQ3,>>4A^Y)UNT
]G=0_bJWTKAbBKS[M5GKEWe+^QS-&V/Lcc^])OHf?_gXSbB#3c(9cK0.__?Lfa2R
LcQ.eSK,:/2cb7;ZAEE/A96Nc9LFLcD&XGO[F.5U-bO?GF_.#F@@1H2BREHXYS71
DGAJHCH6\(c=QNdI[DaD-+5a_2fAg>#aP)g,>Y>4/)Q9G659XJT+?)]+KLA8cA6B
BRa.bFVF?SYEN-[X6BR6?<[/JYf15ACO2)0?1RL6=MR#JH#@eV_Gb(JNb&8#5LEf
/463NDb]-A]AYGK[f6L[9Y01P?2>eCZ<HUUcg[5f,],?4:P_T4VT+5+++6FR3H7+
V&>eB-J5(:(OD3SD7S5;+M)5K>14a0N?aZ2&DL=GFL<YQd)>Q>-[52MbL[8S<))1
GK@/TL9e9ac@GIY)1YH#M#2AY8O3#0-EZ=5(>4,S)(:MERVA_QQ[ZR6A/UDb>c+[
H0Jg#7.aYLV]WWda;9JGDLg6<]71d,CW=Y_OaY?d0B_DRK=/VXH?+e5(K]N3/O-d
e]bc1MQS772f/BL\<HZX64L#).H\<BZ\7[e.V\QAdGIFOX3KXf(L0A#XfOR6:ZKN
f;E6aP6Nf,He5MQF-I9EPN).I;.@eAg).\Wa(XTB[56<K=Y>XO\N#YM+HbC^DCCE
A+>V6+XY.b;OC4#I(aeXb-6QMce/68H@[BDY]IQH=W/S#3/#GVENa3<6HA9K-F[P
4]-)UXR=b@9/G)^L/FL@da+\YHc)P,a.D[cg_DO=,a9(H=U=g@LR5ASPA=1A65()
4M^GLN0.0EJ=R/a12J:AF583bW])S(BC/c;;0@A:)(-BdKFF&g>6L/^D3/JA[f3+
Y8,W__<@8JHaN/Sf^]2FYWF40dc99]/XV)XfDL>f\:OTVZTWG2,0f#UX##eaT-SH
/RRWG+PP+<EefJf^+[gC,_A.Y<]c(#\U>CBRW7FC]f1I)Sc?NA5-&X00&05QEf/Y
8gf[R(e^AF(60?LcT\;@;fcZ9/8bSP#?OG^)WGTFIVWYH6f0<\[(E^cXZSX<D775
XLRO?83If_7LG5g),R#,T^[JUQD9+@J3<)JBAD)F9@cJN>@CAN<9RG#a3\_2&26)
#R&[6eN\[WR5(BEWRW@#SZBKc=:c\XgQ&>a3E]R=D[J/UR^M-M13O+/OWIPQE2EL
6Z/-=\/+a,H8)<WKPe76(L75D9JTTL-Z?O+&RD6_(MTGM9GF#U^JbA2fXL7]e5:9
aY_VA1gAfO1-QW/#2B#?[aGKZe5aX=03M)/21\,HG8KA4__g=E,U:8?Ca5/E:IH+
gXYI4[9X]P]eE]6TO@J@126dX_P8b>TFTUbPT>V.IAZ;6G(LA0U3M#_=3SU1^YIc
>LH-VeeFBVR3\4KQ?VVb[0a+,XGRJMObS[/V?Z,W\X1.Pg#/[9T(RFaB<.S#;c\E
QdOF8&M7dZZ\_Uc:N180HN8[PY@=]?@EOa/_G/\SF^P2^CbGRc=0^HC37Q_3^485
J]=(Y5]Ig;^R<-_GAX_(+Tg8ZL)KFG?/LK[D+2ea=/CGP@ZG(?XH:9@IG>=+Z=Q?
>OX43-ZO9[6K12MQde=3]=FL\F5G+UE_>3.7DUN5]TK>FDX2Vc4ad72>/JY]e[03
AZ,I<3ePQ4/SKO]C+2.LBU/<P?:2U/]MCP3I<_X)/@.>C7ebB.O8\IT\G?PgPQL1
N7CFQ438<EG2;E\NN?,=Xg)fg2c91Rg,eMQfXC;C\;I9^76d9+UL_X/H)0g^<LUP
=@=1IZ?1:bfPY2;8?G)S.D#2Wf1N1_NQ1,E(;2&IOX5AD=+X\G,ae+&1Z5#262eb
P?BUe:&-A/6.MLZL4<a_,cd)>(M;b\:(4[:=\R733\/T?V-4&gAX=46G59^G#YDX
^4^LgV9?Y4AGT/14UZ,(3)NbHS3\,0:Fe5-I\K6^TRBFJ:GD^:N>5^HY=?Qb0\[^
YTI@E/gE8^B64deQ_;7^J(?U?Z3?e,BL48I7;K--I33U1[3#H>08]#R[MD;a?5PT
@SL;cGf?YF]ZF0:cGW]K^:9YM3\OHA4J4HOK>;8\Z>EbDIN<#O3[fAQ<5FbOWC5#
;We<#?EfEK4T>HN>#-[<?H<Z(N<_HLQD]:NFT)-7T46BCHOfPCI9b)Qa:;a)\7@b
0B[IgOd(+29[LAXLe2LGc3Mc7EGY2E5XD/,WKN[HfDR[VT,>4TA?2Of2HZ#[_XC+
9[KDZ#-aD\N(5c\KG?QAER?RX;<_@H3-?^WcN==1LgRg_8H45=97,]IT_<8M,8YX
#Ue>?QJLXKH:MGL77QE=/Xae&d[VQP2@-?ObDc)K7MEIWY@?HA.H_JOe0DB;DD/B
Q2>f<BWM@GSI=gN)UE(Y><+]eJHLQ=[FCY0/O?d/JaX)+B?:-HE398.:^68@4@/=
:M3edZ)U(.TO1a]f9LS@X3_S@41]:YFO[1O4>[05.C?FL#P9C&W1)G9/81WE,3;,
PF(^-:>-4_9,S\eV&Ic9[4^=5bI/1^fP60P;\XV]4eJeSJX(MN8=/H:P:A06WCV1
)<R2@]DWAX693)b^FeGX8O&Z+10IfGDB31EL-.M]2J5/d+QR@#:5C[).FK@)NP<S
ad6.X/MXH1e^[LAUWKFeDc;f/aG\=]B.;cfGP03\[,&(G[<;aPaFRc<.:)8fFO]-
]]e\A,@X6^6W4+&ATE6(:e>OMLJAV,gN]>F^_B67PJJ/aC&[F(X6N,A#A0S?<2-N
VYK:6\WE;KCa\\3N1AVg_T]SDaT-^3_Kb\2AL\)H67cD;Yba1Mf<:EVI0WcKX<#\
31<Q(fBg-;7HL-RCdGKcPL@&93<IA4#0M.eJVF2[#R#A=Q0cC&E@\=&(e^\(D2R\
_M,1OH9TFOCQ2#GXZ90IU@4)6C0U63MQeROT[]L;U(@Oe@cL?1AAJb<g7,LRWBSI
5^735[V/[>2GCZP(\ee68Fa-geUe:ca-8(\XL4Q8.3d;(PY)J-:8IU8662d8>Pc?
Be:)J&U<@I.N66?J+AHB4fZ57CESKZ7JESJ3X@03[)ZaK:C:T<c\7c1O#gAQ<FS3
EaKOcZO[;^>5UY?>#E:[XR35+.4/FA^+(>3N1:/EeM)e;>J8,0+X/)2.YH/A,7Db
+fI+=GN)5aK13(7<Z=8,gVHRTBX.8@D/)4E0;.ER7K?XH4N&-(/YD->_JU5KfD#O
R=0_S^1(4dRc[Ge@7aUV_7D/dPQ/8Mb.OB-=3;3&AL@\#aR/MI2VfZ1W\RX1:XNV
fH<TA:\9715A7?SXa]S.VTP4/EV2Rg)L4OEEI99AC7d[[KZ,<bB1WQYXS<+^-9PU
aJ/KHC.FX2C&ZJ4DZLceae40T5H5E;G,57bc40KOA133N>N,B4T85/&TQZb_[X8T
(X@/6fXa],c&P<H+=K)8,eRgR(/Ob7bFd<0JM3)0Q@7>EI=<#)-#IK8&5&OS(dCR
B\cf^7J1,E/F)+P<e/A5[/4VA5T#27-N;Z7X\)eN\\OY2482J]W#BgdG^QIXFfM<
;SU+,,9\8EICJ(__,L^E?-1dM]g]C\Y1FH]WQ9P8,5@2fB_8PH6gI&eV>8G]eQY9
(])+eM6,^1\eG,V3S35ZIdg@=:#BK9J);IQAM4E00d:M_7LIg5G;\0X-72SdLJ,Y
9OHCGS&e2^U217^6&R5.7R?>5X<YW:S)M<1UgcaP=D4PD@X47O7R:G3AQ-2O;99f
-RRfKQK_6(P=Q>:a1.19dA.)Wd0]]@+U+X_=O9eN[PeE5]?/BBOc7--GHOL8PJ)6
G[1>/(ga;2aVZ701P<CPPfd987?ZeKU;W_NU>D+Y(g>4P^@/B>S66,AJeJYL>G-V
/g=OC9,B6Sd5<B6I7=H\37cFAc^Q;H=_#P@g?-\V2-H&R><@POWb[P_d^^CeRc0G
UeUg]0W/(?baN>+<LAQU>)=A[)F_,=F5ER2;VG>MF4>HU3=IW\JNTf@bF>Ue6M9Q
gM2&g.QW1CC4^,\DU:)DORNBLf(4a0HGLM)#S9cEa=:a<H1^dbZGA-+RJe_/,(R-
O4/]YeVR1-3?\]Jb=Bb52VPBVT2Y\WJ?O6A89,CW14T^?fe^5d@(C1?,)40?a>4:
=gYB\;_f:NFGSe7f3[>PdGK+dBPL95I-@+YGDXFY&9bKd@V-P_F-+:ge]Od5_X9D
XH;KYWDSY8>L0]\(gX69AWKIM70C_]>06V[@KIHVeWY5gNHXA,.59>8L+W?2+OH/
^\Q@d&gd)Xc^5U)(Ra)]D1/HG\dQFGe)U(-XUC&U(+3)?2(9f/B)5LVMNg7M0V2L
-ZPNfJcbP7W?ZPR:ObY<M&DMe,K4_?.9Y&PKPPQBT7g,NNTaEEWEd41R.Z7eYHLL
XNF3(X,_#YP.7A;\U</P7)IX_a-#Y)9b,SV?fN.&34c<R<D3=BW(,4Q-I(eXF5.Z
8.T&1EeA3g7LG2G4OSIMIX12#JBASfVEW+6>S<V5P<:GcN2M+OD@BP\eT/BQc99.
.M4@M;=PO0O6fI]aH>b+^K?C/772_(:?@g3VZ1S0QKCM5@^84IDY3dQcLE/WAe-2
_A7T@..H\P[(_SbFAe=8aJ9[.9ge+_f;N0]OJ,X\W?@:]=,P?31&e./F3/.FR+Gc
GaJBH[4&IO(:b\:aT6T7.;1c8G[gG^cVTFHFZQ#PcRC<KLEagQN&FQU\3+(=W?41
JHDbCe)>D;D9D?J9RdLA0e,\X1R=K0V?#,Ba=0C_SN,c@d\3ZS;3N89ZO/G^MM2f
eff/\&ZIUP:V&S)\A@#=JW4)Va8&,U]ZWA,-4-LVT&\?<B8US4/)0;<>W6D;_ISP
6#\)bN5bD3_1<PXaRLYOFC,?QB828CU_9[JUW9g;_eT1^5?(B[\KZ-gFO2F;YIJe
L\1Z@9X)5ZGL4@MNJgBJNf=f?.H(^427@PRU9YM9KcNQd^V1F\G6.&>J9J?^+&9L
?QaOSEVFL726RdT1_3PK[W-f#cHc<3O408TALT^FJ&[AYK@FNZ-RY?ZOWUgc-GUa
?NW#E6[M.?cIA(A@Y83+:VO5:@GV^5&-CS7._=S++Q]I#MaC]>E\J]8FgG\.8:-G
W)GC@I#XYDVBB)D]_b<@6UGN^K;(8SS7>>e;7@;6SaMTDa@\P9fB7MR0P6D1=c1e
7@ZPadZSI3WU9YE\<G.->JH/F9;:?TQ5JFAf#]d&\&\W>(GN.UY6JF93BI/J]VQ=
aZ8Q]fR+df.bPW^(JP+BP#VJS+f@AKAcAg;YffIDfH:bfXSR.V6=//BA.:H,YS>-
b(Qb^BU;(#R5S#f6(JT&:ZSS4f@F,OR-1[>Qf&XOE.<6C)aQ#;7_T_D(40#>8^SB
C,KZF9M--;W4#Ye?cGUR;H1A,[/IQ2WN0F;MZ(S#:^Q&ZLE?Y8_.6^^0F]Y^F>8K
c+1)X9/D&gJ@BQJ3?U+:3Rgg1^J1Z3U&7Y6_c2ZHeS204#-1@@<,>S2=F/SGMG#c
OefYb/<:QcU;4C?DAULH3IKMUDObM<B3T@Ec2BL:_M3?(c3VN(e&)-\_XacCTC_M
13&7a6Ub[>+a#CJ.31L+4f^O:,0L9O@_L=dCLS]K/FHN],d.1=-Z:dW\;99]@U\^
#V:H-A4:0J&\L2f:U0]K#E,aMBE50-HaYaA,];E=1S8S9DL,dRdfa[#R>0:ZNP9D
7HeRU=L=LD+@([LZ95FX=7_DLZYW+E=UB6Z3(X\9(6fYJSJ..O2)WC/#YFXH8NBU
B2TXB-<@F490>,?H&#3e(9GCTfT.)c)1_>C+SFPVd(HKDCH;3;OD7A1#\D<5/YOP
Cf:IL+[Q=X;.UL0Ia)f,R5X\&X2)UQ[YF@,A68OEf++OSZfe;Q57bVOT.NO6Xb?7
M:fRX]36P_VA)F0T&N@VL+Gg6V7@2Xb8Z]1[)8?eRT=Lce@4PMCAe5.acBOB.-_N
LMUU3W)_C6SPHWHUS7Sf/@[<Y+a]HU#?L3+(7@]Ug,Yb@C1YD.EPV;YWGU[-V;M+
c>RSDN=KW(>O6U:@TfU2bVON;PMD)Lbg/0EdUT==)O@4DB6CJgbT(@6R46-FfK+#
MH?BFK/QbHe]-fV=04^PKMZQ2S98J&A\0Q8[KOKUS2J[b9SJd[DQK5e[8W,&39/4
Z4PV\D+[faQLfPKOBde[FCSV.EX5D<,BAHMTQ8)4E-g&1INQg2g]D;>4CUU2I&_L
C>MeO\DV<aY3@L[)5>O\\KE3DE7fB31BZT&(L>g#,WVK#8[S)c?eff[&FD.PIa:4
W/_MU+=I[43(MV-Jbe<bcUR#^3S,cg>G>&0,>AfC5f:M++<3(U/N+E9Z<-[X[M)2
)>R[dE@X[B)]YCJYRGQ=G65M&L:9aV7ZUJ[ZAQf5)#eV;g8WJ+a8]KGf:(5f/FI?
[_=,Y)gZ9[I2;d+[1QJ119#ONYfM@?9L]TE+Z;RF518?1)]#).C;B;0ga1[b+I;Z
^:^,OX0Y)WcT5_3^DG?BW_YMKQJ0cE8DIQ#C=^;AW(9T<=82c0E.X8WGFG15e[#[
))1S9c@H[,9^6^F#P;Q<Z6PMS3JBY8BN/.T;e.G0>EcDa5&6_2b\PC#P16J<.[IM
A@K9.>N-\EFWYC#P1[I.K=R&)<dJ<ZV=TW3XQc966\-7g5Q&(&\\T2,WMN;NYUd&
==eM8C5+TKU7?Oa-^VNWV]D_]QX(G=;IN@;/)C&7:?\GfaK:<X?=<BZ^UQ:V,^V[
bA1Q_-AB=,fYS@,HNY3U[Aa12dVIAE?(BcdeT7OK\:[1I#,JJ/Sa#c,gV:Y?-#S.
KA4;JE72c_Hf9M<cgQM8e[bd/>S,e^7C=@M[&JGL=c@GQM/gdO.UTV)]He#DZR\B
LBc:/E8C#26]N\/VUTF+VgcC2A1AbA^]F-G8-&YG+7=QW4L[8XYL32K&+D_NB(JL
3+7/C8ATDCI-I&4YQ,.-aB>P363DEAV#,R.S:)1&S6LCGWg(9S>a\9gY^A&2]aVO
??ed_WWV1E^.D46Da8(#aN^@F?6>_:TB#LU1fHF1-)7HJI\Je>C?a2<SQI=C-8G+
[fCWGS=7D-,).#bX02+Y[<)=e<K5WV;aU/C3,2g<g]DR4?E)CgVPNAUS<0Z=9/O@
=J]+6R0Me^IR4\2LPI[X-\^P_=+0b9\25:=fY7D_dH;3+[@d<M_U2(>+;G3FNb54
9:QcB];D5.gDYC-f\g>eVKJVE[fQg\(&6Wb4THR-7+?Ka9GGa]@DZbY\=9(9;C6c
c/Y]CfR0J&KI9O3L;,M^^C&1NO=Z4PEOG,UC\PF#cR4QCS,&Q3?JP>-XbbP.SLTX
bD<&@8HK?Ye]I4S2eg8JS]LFY#+_@]N2/I3:I]^Cg:2,L]<M12C16Z1VQ.GeHH=5
\\HO]X:g7]2\FeO[)=?]IdVJ/J7\,4&F@\7]6[>KQK5LRFW6<:(6b@;;d(XB1+,+
@MVTe@T.N3Na31C1YGN8Z_23C-43>UFSMH@)BQ1Y&D=VEC/OTGMTN6PV;)UI7bL3
^FSPSQX(/BW<7+?_KSN=d<Qea2J]MV?Ocd?DV\VI=8RDI(RH6:2(08/LG)6[MH/#
WNfc7,gdZ7]UgW&Fb]?S5+),H=#QaYXd2(7E1418d)]aN(6<F,b1H^&Be]-g/<3V
_C>ZFB-+f_cO:JdaI6aG2c43[;g+=2B-MT]G4N/H5?AHGQEff<IBaPH:/:Teaec<
4N5^;\:G:H^CI\JX0Rg0g:_8_CNHf:[O-0c6fcVWGP\S,BH.GKD/5TMN6fBJ[bTM
gE)YfQ1BJ,-=W\BJ=SQN,U6RFa8.c1\9HTU1WS9?MOW1CT_Bd]G):BKKV7\-/:[-
4KXZQ>.,Gc+cM+9fGd[>dCg0P,U5TN8E.UUP]5PfXb_[U+NDJ;SXHP][,KYHFL2@
F>d++Y6R^6ODG<IKTG0>;eM@E-ELR=b5ZQQQg5FA/M)b)ZU@ZXU34/>.KLe1(\HV
WJ^e6J8DEE+gbWHYa-?NS14-R-/BSRFQ#I>R)QfC.^N-_30KeV8RQO/I-FYf-T#.
EK9KLK2_T9I<0_:(>UB/?cbGNG8bY.W<:U\_a31U_DS>&@CCC,MaR^4-.,YN;F6Q
/]gGK.a[/\6c:_/g)JH7\]B-GI3gUg&]G,c/FeN]>N4L_CITcM=(1aJ8V1+6\+A\
+778QfgOEaTN;7?GD,FJHDJF#<OS:OQ\APY9\HN+HbKU5#a(2HB)<0/JFML7V#Ze
@Z98_\U@/OU+F5M5,JB9FO0V.?T&X#;.QYU8RWG:8cG5<W>/0A/IW6H6RX]OJWEH
MIGF\ASgI9I96CG,0+G2\GRUPb5?:>_.[=KWN4\T6[L@a:9;<GLXGYZfEeC@)fX1
S\=cgUa34K5,E1fU[AT@7XEY2R,O3NJ3N(K)7UW4F)N(e;-P.d(84986BUKHOa;U
f]G&F)6g?UND91QQ,:(G7WMHU[;a:FR=9#E>Cg.UO]ddIS4]?=OfKI?TNIGPA[):
X4F7Y<f_K9>9+D#B3fOcU@;g=;9QaQ6.(X\<T2=f3SaC<ARUFEf\f>)DV[A)QM/3
7JgS_/M04c#>VEQCL7-MT3&&QS0??Id+XA6/9fSE]Q;=fc6HbZ-QR9BKK[]N<g)I
5.^AE/6+T00/XPX3@Kc;_fWV4)]e1)?;EIS[A0W9bYG#]<XJ?S=OG=3a=C4@g;+e
9R:92eO-Lfb2MD;GE55eG-V_PV@ZP37c4U67]\V6@6-=O]LcWBJ9<O;;P>>KHYDW
6g;>-JWT+bd.SO+C&g)g^PZ?^.67N:CU>0Vc-HG3\g>KEC]Bf4/,CV@63.,P^d[Q
&Z]9.^05,]=>LZ/JXcR(=CD<EG\L@@/0a[f1=eG4-UT;cB0G1Y]IK<-3NDV]eUWV
@?_4O).V^bOAZ/f/DBZ:3;([[0YQ0+LIWD+KfBE=D#Z8.^-N+?4]9I[5<NAaRN,-
aP=:]&Ne[W5I#G[bY:f68;)58d>P+:3e4a:ZN)E&D=)f2b9_,@1KMQHKC97SF.4X
R8MRggE6e@ca:8(Dg8[SAWY#YaCDDF?NH:U?T\EJW#OF)Kg,6;UO<Ma;1\PZQCFd
/UEU2W.H6@.12<KLfH1\ee]CIXdY)LJ6XCNaJ=8AVgdFd>QMD3/O/B#EdgdF#<M4
FJZgE?L^U;NCf0HS,1KVM=?G:Ha@24HU2a:@=Z7EUO//4&0bK_6O][cT-OG.3Q4U
+eADB,Y_7@V._GAD/L@)<@Z&#E@^Xg\#<eQRK7WY:WXI-C+QEJ##(47P>R;Q-\@,
.e_^@>BV3YHe.O>[D=.e,d\<R[Z6]&UO^/-.=.:,8LaYX\?15AS4EWP4D[\I7+/L
R8\KHZD8(I\B@4Veee>;:M,<I@,SA)RJW^C^Eg;J5c.+cQT7<C]UIT-fMQY/G_;g
CW.L,KI)B12bIKX\XPa0faOA#A#@V/cWMPP:^GgODaP,Vb-DLX6:=J<?..5gKPB-
058XEAEM9M7Ge+[6c+[.6=&CDGY7K25.Bg3ZH)J#;RaXP8Rd]W#[dbFC)B/WTe&\
?]T4Ue,<McIC&]UBE^e4/bP(3PJ?R/U&-UVBTZeZ&4&78D&=a&E&MO:e88YPLZ1T
5#b^W;^3LY7TRPNY2M.2WgY::@#a)f-6B(9_[#R>XX:ZBY0#0A7P>;ZO8bRX4d;S
,.N\8U(XG93:#3b[WLO(3.e]Ug02>IcRC7WeB<DVUTfB/V]&/4bNJG76M-V4T[Z,
Z_I\^^]JX_7.eCH,/;@A?O#<?E^G+ELV@7<a+^L/H+4V5SXEX]f2H]+Pbb&Xf4X@
d8IRHOMEGE7ZC5[ea#c-/2;-^?VSG^Y;C:+GCgELFUce#(;H8S?WTg]GJ+I]DB&6
d#7BMU7>]U^6cYT&9ON8)CW-dV[,)QaY:=0AJQfK7.XXKaNL_57c,DU=M=\/(+N5
+?e)d&<EB&/2>DK;b\Zf(-FJb=^Q&K/<FMaf.2U=2SZ.NF__8?X]>EB9BHO#c<5a
FO\abPZ>fADN9_ESGE#T&W.18DF<.UZZZBTe#.ZdJOAM&.7JOgcNgK4-Z-JYAG^1
>5+9W?5?c)@LA>MKMD?P+VAI3,4DWd?#6WBZ+=fX:AHLT&UJ>=dBB\_#c@=<4FO\
QC_L-ES05NM+#P@&:18a+8<f_]C@_bL^I?1M9e.3?@DCF1gcD6gJT(#?57-1)]3F
RZ_X;TKXKTd)FWTAR1C/e9>8>>2L^+Ae<Y@0WdJ6QZ.\4;&Cb4.)58b,BcAB]fDC
C[Pe&:N-&\d=JW<S@DU(>[4C,(7-\>fP<gENPJCGJHH@6.6Y9Z[:X-(756d_IdOe
cGO9[)4\4XKU8UD<=YB3P;T,I?EZ/P>a;C>DL8ON.H,Z+N>:gP4BfFR9a-NE+B;?
eE2:_)bdSf^ZG1b>d()bEGR@RYC]G>7#RJ/UJcS<-LXJKCLg#W;7-NMY6/7FGDc4
_S/.6Cd>R6#_2I5A_C(Wg(XGF##MEO9[;,0)AO[#RHEdXPI6,U5EC^e9J7<EWPRH
ON@@+>CX]f-[dBg\?[g+JTADCHER1;MBHT&Mf,6(2E:+X.TA+P\?e\M9(RIgdF)7
&dN1?W0O6]7e4?W@/ff^2GgBc2Qa^=>K;JVRdE:VLDe]g/QdF-(@UYJ.2@L10VUQ
W7gg@/G;]+RY+S&Sgbc:\=1fc_@cK92c&8UVYTW_Gf9.B)g2;].S@^1BRWX@^\)X
D=_Z:6:4Q#7D7@.<adR_5SM)ecTfYR.(9=(A_Q\B@B+CaC&[5cdH+ZX-\]-98L((
:fa84&/,:@U61c&9H=&\FY506PFE4/E9d1D@R;b#c;gNQT>88g75Z(NF;=7e\P-9
eeJZROM_,FRORBW=VBYNZZWX&C:4UbEJ<NB-f/IO;S3BY&&PWA_=JC3V?U0BPeFK
HHL6VaOI1WHC18_,[HZ&]GI+73#&R[AfCLY6[1M4Yfb.H).DWA.=G\ACS@JKGQ.8
KR9;:N9S=3=04V#/P:W+Kg6H@YKN->VgD;69MC=Q^IE<\8[F3[bJKEX/Y]I-FN[H
dPQeWZ.59H[.eH4a24TM.J<@=7+e,@ZX4eCSOHJ4P^=a.c(NbTc<T:^b:L:FK<I>
aB_e-(BN/Eb(Q44EQOU5CU#2-^K4G[V^RXG;>=Xdf,dQKc-:Q<b>dYJ>XM00]L,E
RYFK-QgUZW[6Y98-Vb#&8K7gVGT1Hg:]&Hf&[Jg3:R7.=:3<>#3ffC5,.O)NR)ef
+LHT.LEY;ER]ZEZ0JSV?L<?(A(Ib8U1;EF_9]2-4+K<&<XUdH--[^aTa2[5WZP5O
46?HA\;I,K(A-W2/U;23T4ZP_D4ACI?Z2).:##GHAD18b:5=)bHYTP;)>W:8bG7a
e>=1T@^TCK2[>ca,\f+O&WIZOY4B/b9aLc&Ia:c7SK37IN4>I5MdI&@=,:OT(H;W
IMD;3C\,L;FSI1JO/)#SLP2_D^)8H?]S>U>e9cf2;g>C[=9.YA3Rb0ULW\<MKfB?
K&AT)(&fA?UZe_G>IYHU:#BZ]Z,N#b:?2a:^Vg<#XH-#e\-PES2<a9(UXTa:&UYA
8@X#A>4PM=<M(?^K@J)EW[+S5D#.038<TM?H74?JL],3bNMGVb-72.5F=URYLJ_G
=e_FT?a0eQFL2cJY=>&/@0&6W[W76Da28Bc-)NPDAPKZ03OabH9d/bH&=\7IS+)G
cH2O5/_.G.+dJLQ8+#5^.c1QgRQ8ecO8PU&.50OTX1/^-S6EA#>XL04eMC,XIcTG
KTg)46;1NG7DR2c>1#ONRF5S1Y)T]26Y>P>PE>JS)7G@A?5>;R5DH-,[[GYW>6;A
OC;\4e.UQR@K42;c+2]2e9WNda<a7MADX+W&]TbbXQ64D==;_77612bc+?2A:_&_
E(^g:bT11NO@BbK@FP=c[#Vc^F]&g:gf7ZD;3WF+-?2Y+DH]F/JAE<daM1HM>[M8
V)YdU4Wc[;8dRd<2WFQ0^;BFZf&N+N[fMSZCf)C^;ML70geUUN]X8#f:]H\Tfe#a
R^L5O4;Kf00]bdMDJ<<dWc:SLB3XE#3M8FEKNNE_H+(RE+]Bf;G)M\L<:X.g<cP^
AbAB4^V^DXAMXDYMOS=dJJH9@;O+g(8BE\+K4Q+YPeQQ<]:E-/.d=LI>W\2+CQ\,
?,/.(@1;U^@g4M2db/RR?YQTTD0_L,d=3d/H_&3VS;.B6?&[bM-I^bGVIZI#USZ=
]Bd.^6F\09/JFe@d46EBX7RK3]IY9dUM^:RbfdG[+NY6Df/IR\gM4Q_0d^.eIYH6
6)7CL1,?+f.,QVbA2]=30W96B[d^Q3cRL9+5cI6Uc?LLO-4I[EU^cY@,PYb=6fW)
g2Jce;V#T)SHeFMOLK<.:I@D4bZZ-[_<5=]K8U&9)KA=eO[-&NcUg=)]Q?P>V-UN
CbMc[Rc\eUB/J^;DTcDG1c^b&RA8/T1_89:M=KV;&>)-^+9)+(:]./RS95ZUGQ3P
DL,+KAR2:\J^BZ865M@14<gGW5Q34@c5.+g90@F<8O7Y[T(:4LQI=6HV95XLHJ4J
4>L+U:_-.HbK),g.[>Q_7bMKe9B8\BA2f[X,69f5;gBA&0-TBA^WJU6_ZCPO8L@,
8^5f^MT<FP0)8MA\JDK\JeO/dZAa#WPJH3@M>=d)Y8Q-X195FK5)3#RS_XDI;94H
#+?M?7.=a--Eg(&MIZ-^7f=f=Aa0-V&Pc16<[TN[V0Z8Ga]O)48,Z[PV?eC[#[+\
/Z9N-[I<>+YJ4J/&Y?5b:4Gc)_?SI/?SJFL3[=6Uf.]5[c@:b7;+9P\TZ]6H^aQY
?]4ZEBJXN@fRb<:>XL<L7WZAZNTUeCME8,#6G><WT)VBR)8_)XB@4XG5Y]fN\S:G
OC-A7QHbBG-fF#RBba<93+O7<I4T1WYd;RF3]#8MU,SR+cO+88=8WZXK[/aR53<;
eTIaT_0IIFK6Y<=L#/=0MY_QW-]UZH3f>=0,9Y@dH9##FU+LeR,G?W0AS](?FV2E
F#<@?)T(WW#15NG+B)_8L=fN^IQ8M.3JY)Y&:eXEAMWJZKa.e:9?T^X7H77:.<dI
E^^a_2dSO^,gg5ge+^@V,(A2<X\+)\HAJ3?06_H,1Y5+e1\<J[(dX,++T/<JBKS8
@M\Q_Q18Ud>[1I@Q2QML0++I28LH)f5==abIc@;@V=I/AcF.f6N8ELGH]JCM1SH#
d@/BZP0ePOPbfZ3S\@2Y,GA?]0Z)C1U;\A7@8C3B9CON4AH.(G^+Sb/C##O=QZf1
(Q118PM<f(V&g=GF+f(\1K@]Ub<KMQ@L1-D#-F^RE\G[@dDaN/b&gQ1+W<>ZIJ_C
eFO-=F/?aFJ96S&)cf89<6=BPWUUPU7BQ1^0O6]OMeD5J,E.4_J(FEb-fU)Q6->G
F>O@H96:9aO@8+,@_KM:VUg2Cg=8aTcQgc6Mf.eRbF@:RT<S^8-\+1FRE[UAf2X)
;IES5WW\)[CVJSc^&1V+dR0E+?VS6ME^4=Xf><c?;O/.c38/Ga5)&))dENVJIHDb
\;CIa60<(0J1=V2V/CX<QXJ@3^4-_=FM]>O?WaOMMUU>[X]f5Y[7cKe31S6.6]84
0WBT>R(cO7K<bZdC.#=gR/]>@b\[KJ[eRMG5N9QYLe:V]A)J9(,(+8;G-R)_6&=B
1N4EL+]A(^aJY+]@^588#SP;g>Wdb/L&N&F&1A[#,/bT9e#K(7;9_b@NNN<))cH>
BDQG,e.Ac@f0CU#[Ibdb\P=O4DOX0d2=<Jb]-Q-7]H+GNR#_\(+gIQ&?Cb8>TCV:
ZP?/-&&+_@G[<1>Y/?fWGZb][O5X<B_(df;b]_?0GGA6=BLdf[V]0FUZ9#__>fSN
/;\7[Eb,0>I[R3VQ5MP1/<SN-.;AV5#M)3Y.EE.>X6^Tae8Q[c,2a)@)KVWZYZfH
c9CbXf_TY=:aP9)&-b4]5U[_M:GY\#L&6,gfP^:SMaED=Md)_ZK+b.3C.BTK8e;K
12=&B<7M^-18^d2-E_;>076.]4W_O>I>5WSaC+9:?V3WA]=^[cF;K,YT/?f(J>24
dF:GL7OX]U@V@[ce]2HEIFb>.JAY]I]6.8B&S@e3L+S5,ITQA8#@ff@3AB73[/,D
BH3IU7;V<:GA]O&?YM3@+U\>UW8;^2\TTEd]:?9.BY9c7]W+feb2>2_WBI&Fc=Gb
V)<6_beGZUdMLUNeWOV/03_f,;#f.U7g#28F7cC0Y>dEH\gY612N7U(T:8:g4D)K
HA[NZb?D76)S>]B4M/gZ#cYY2(<A3_dEM.>6HC_=[MQRGdGX-]1BXFDCUK0QcY4M
]A>Yb,M.e+1SUTSD5\WRJN?R]cDOf9M6]c<MI\R&#HN4bab,1D\<d5/,XX,T/dKE
GYSWF\_VF-A[BbRU^OK,T;&?-[;WW.gR?3@-&_+XUPGT8Y0&7>+M22>J]+>[fF5b
KMJ+Xb:d&MeTH8P45#5a9-E>7,2E8,4(25S)-2VUOP6RN,FLZ=4)=#1NK:H3GI:Z
Tb4^S/cJd:AK3-)9,;,g0dZGH\d/2HfV3S(E_)[=#OQ.&f9E=dK)3d3BQ-c^SJ\.
Q)\:4Pg32N1.B,Q:65.P^cQ_#C>fRO=a?);I):SFD,H>;+f(T,O_9HI<X766UO/Z
K-]dD#ZFBU]fKORHOeLeN\2X>B6g5gf1MYA,34UC@MJE62P2F)TKP5,#OQWMeLBe
HKfU0NOK,[KI>N\:1IV82;SQ6&ZOBL+6<@HXR<<9H<Q9X@>3X#HMM5CAY(D2CXF#
+,OA93g76bZBK&Z31^@(db2S+\)b5D0.K(>3D?(I#B?+FOXM?\D]6[,H=9ObTRIW
+:;C.+c.4ZX6c@K1ZSYM-0&7&ObRcQ@+<eG7G+E:RRI#]X7#J5/L0C3M6(ZTV@>G
PY4L4=:Oe2M2W-?CU+@#X4Zc3_&#E3SSNgZF&AE&.U.W[5:H;IB#AZd?(e_Q9H=b
[cHZOG2d\D)\S8X\XOW3]#]KC&B:CGM5g.O?S[[dEF4e2^;W74R+7ReI,1H<U=E0
))PR\QMT;\T>9e#6bU368]#a0;<#5PWDQD5^ZT2gMQ)VO&aV[GDA+##P_/,HLc]g
LeQKSIWfFHHNH.;[#J=;VBS&a4I/f1G/S(?GK@BX-_BR[Xg?GLT<AZY+>/&Z[3UG
0(IWaDSM4AY-Wbc=:b4YgP:X=cef\aF/RU:I;Q,7,^A3<:;PKEMOe;b9RADdSe0I
EHNEH.?gO>@7Jd+B67X932\EZ?HKa1B&bY[^+T11c1#fNS]DJ\HU2<L]1c^DAA9@
1c:DI(6G46feN,(E3Z@04TDd]ET>G4YAN2J]2[a_?<b6[@8G;+RS;UO[AEbbSU:\
O<EPH?):?FI,f.^Q&CDE/94F+?Cb[#T_?W_:Qa40;e)RLS#-ICIbFB(Y[I+a.dc^
?=U4TTZd-3YBT+-_4O^:WSE,?66I,P23[F\;gdNg.Hb_NSJQ84B#(Q#@EZ9.WS\I
aHcE59YfF-Xag_<0#W1CV5+L;G\1@S#(f9bW2?a+;?5?KWPS]=ZZPXWK2D&&QCQP
f/G.dVVY4eNc_\]X79>TQ;67=K-^O2@^g1\ULO-<LJFZ6UIH)>R8fcb@ACCZLBUM
Z_4,?5Q07e?++QX,T3=+fPH&<X8G5;&R@-cD;K0QWPA\?AC,6([COE-,,Df44cG5
&C@RbKLUW@1)55T47PeC];J5f8\FH?9KQ91;4XBTTU])R:5<L9WDYYNABd:\&@LU
Q4]0)\FK6\/RMbUSW59)H0g4/E4=UM:=.U;-bU_4Ufg7Z_gGH\I2/8>2&6.937CK
U9F_LTXDY[c;L-O[NWUDPS2gB#X.IN/eC(B115EP8aE1T<cOg;YKT:X#[-+:61>G
5Va(R7GV7JZAb@gO#L^Y(G;0G>8WefTaJA6H#)@d#=VFQf]X>HP1#)7GLJTI[Z0Q
dLP?+5g>OG\6@;47I6&5903_W#b]D94I2S;f.9dT2b83RSa6(JH;YdeMJ#WXMO]=
VL,UDU9B6KLEURU@De>)WG<g@.,XE5BP3R<<G=+\>8b-./HVUT7W,VdYY<geU&#O
?\9dA1DM_J@/5C+NI\XdZO_(c1?C;WabK.UB.;f5[/U1WUR\K14fa2]WQ8D#UZa7
^R[OMOcc6,^aI8.7Ed.^^NDE:G&7@2NbH4e@5\B.Y:83=39c5I<U)5&O70QKeb4b
+aDbEXX7J+cNA#2d5)JefKAM+ggeW\QLL<?c;M&#<Tb:[c+R<7I#Q140NaBA3:Y9
<L6)(\(H-)RC3LPe9M+Y,,H+S=F:?87-D-:B#e#eaDb8GNP-HB^]e@E9eHK<dP8T
CeQ47JUFf;EDE/Q:;-.&T[cV-6#b6>/X,6,Y0I.@U8ZK4Xd7,G@&Ma^R-1d&:b6I
7L8QHN=:YN4=65XRO>//)-H8A_=PN3DCZ)MB=5_V(/7_UKF@,LF:2)JSIFIRZ7#:
4B1K\\>cDMKA7:9=U:e;W/>E]^\;aW-/<@VH4E7EZ15K_-Pb.S?U(Y=&6f?X;5ER
=0\8O/U:#DKbZQ+4J.ZeaC\9gZ-d3]CBM_S#9ULZK.I#g,KgP3MQ(T;6_FR&6>Qg
VA4eaA?MN&]R>c)3@g298O/>bJg>Y[KW4LfJ.2LE(94_/L<Q9g8)cMUHO4cfa?ga
<JA44_+M_(@0MTa:B)]3M@fTE^9BV)RV:;HN-^JC1S<a<+AXLdcQ>GJU@L7UZ.2-
HVM.M5ER@^,f1T&43+L7>2PQ/(4)S9Q5/.8Hbde6+Q7(R28YRf&<]NMZR.3)0a?6
GYQP>U7A3&DLRd[5L<\1:@F=Z&L:H93DOY\/>^35@I\Y4U1RNF/eYc8agM8L[HIY
KZ9,=d.1ZCJ[A)DH6A@KJO^X>71,+PPCG:?&Z]eNT-Q2I.RJY>1#LCf(.=_a=afE
K7=M-DG-aNEJf?9KBB7d;4Be70^Z<\^O6T;RY.V9J9Yb2MRe1HO41;?==FV>.E;L
/S++D(@G#>VaTT0Q4E:,f9.DNUE7[Zc2EadG#_9?=PFggRD(SP,[J8F=_ea)=5(G
JD/(5=UADg&gcI=+^^0=NI\0O9V]/W)c]g+]Y157a>CO)TT>6fOTBDbUXZOA)2fc
6f45#[&O^E5OeV523V()T[U[&QATLI06We:[9S#&YCXa7#WQS..\RH3bZ;F#82_Z
6;)5^&04[>8SYC9>]:>\.5K0cV[SAIG9Z]1E@M>IKTR<QSZ/(J61>J(Y6g@#&3J=
/?e:/YfXNT8XI>FGMX?d&CJ7C5BGDg/&Q3;7E3a&^,47]-e0OJ?<DD/+GR,[0b?d
T=B]OUCgY>WALV\eH>:>LeeeBK\-WV@[2HHQL_D/984R+FC^Q?@c0fNTR4,BfB/X
6:P21O,2f>&[]ZKGQAGN2EU(2VYP[WY^,L4C2WOa5X2Fe#)3^R(@C\VE5B:;aY-8
OF,J-N<&3O,KSa=V_7F.A-5MY5\W80UK..XQ?4dQ;LF^c91A,MV:(0F&P;gWI?-e
T&e2F^,.[SSV>[^HE92_(cMTc.<?M?;1@[bB+HRU;LPYJZ2UMGS0IAO+DgAF(.DW
8FgJOf.GUQUNWS:[Ad/U<CEY_5,(JVUZ)HRQEAPO46.:;Pc[27VJ#.:/^10)N6@M
E<,\5H0dML[R4B[/EGfT,)LYX7Mf(,B;H1U;/NgZ,MNcg4BTKPN6_+,8?&^_0G7b
?HL1dJZ#NNQe_YY[^??TTa92Ca3<[C8Y]^DFB[VRRRY[g?.-4>D^,F.S1Od6Y?cC
6P2&]E^O_@E:e;+PH^EWFW(9G7;HUTB2.VJAGc6G>@b\RY.(H^eSXO6bM<1_Zd;:
.#V/>P3?Z[EI<9T>NWU&G]+gOYbRBB&ERFPQ?-bZ5W1Q62.A.@CWI1D9;JM;OR5O
25[KeLW9A4S#JN>/)#40.#P5TR6M464M._=U9K[[S+BR&aM_1#WRag,2IRDIP#fD
07\fJ6X1KeJ0.fOOFK;(#KYUUH0T4a:UdKZ4D90X/?\cR#=SfDGA8+Y&Lf=K3Q(J
1,4U,0&@Y2fAGZ(<L<SM.O1be65c+/8?E[(R8K68FQJVUE5]>&&-(O#+a@g<-Va8
g:?=ZV.E@AV>Ie2Z<APX=VQYWS>[;bYR_A8_52eYeA@O8\8Be58CQVE@]IVA/D;7
b2MQJVJ49S[#JHKK=HWJCM#UT6H)Y^,g8J^O<9[C=Pc<B4bcNgV3Q28N)DI=K;H.
cO);L0TFO:WW<RG1&RgV&?)H+N>-LRga6(/fd^52+.]VYB_N8RdM^.MSKH0e\(AK
U;_gB8SM5--g_?46+Scc.TJKON8\Y(C/Jf6J9V\:1J2-K^Y\>UR(Z^da2.&]KPdP
I0<R4Hg4RTfQFLQCBCEc_W<3#3X_]_R6fWK)2(SB00YcVfAY@c1=2(]3c]#JEC6Q
N)1)JW&a^(9^[M@X+L0)O[Q\OYJGYA00[8RVK]&M0+AW0/2)-^W,(/OReEICKgb.
4M8R^3DALdR;-#/MORJ23/f?UWTC5g42ZJ[./[Za5d;V[FR@_A/@a0ZA9LIJ#_/M
FY6Ig:_>:JcE&QKPXM[@=]JS.+V(Q[a93H=[R#;W7G?1)^:\PWfS\#@Wc@92101Z
\674SYO+]F78+F)4A/c:g(b<P(9@88KDQ-GFc9HI^V)ef7a6e\VX-caOgBfJLNV1
dE]V#QLO/M5&a3V@H_W&[aF2).UQ@3MA0Zea^.7Td1;)WEP>/8RH#Z,0NfLQNR6:
&S<:5JP>dCNG=LUdg;:0)316^e-IfWe9T.cUf1Fd7NI9aa@0PH.61M(d:)025^6#
-\=_+4+)g66JbX17G8cM63DN-G+gO0f.g_YP0\#[A_(;[5-^X2=;SGD]<K,\G<JE
=a-^1Y.6R6>[CRZ)\5b\L=VdV^>Cd6O??Mg[XT&4&?7fT5@NIX?V24-B3;AGOHV=
ZD/fa7bG/2VKCWN(S<;EQUgFU/R-+;,+gZ7.<+0]&K]4-CV#b?MdIJHP>dOEP#[M
_@8_E69NaLc2E6<ATSg=[fI+)/0:X\<g[;34/QH)PQ0f=;=88e@QF;=8/EO/FYaQ
N3CeQU7[V2=I6G4P\=,d<RMX9a(dU2F=..CYH=>Dg)94dcDV,H:)B;W2)>D(K@13
A=-<;H)(O=OgZ](A54W<D9A&/-I.0R,,a8/TOX+/Y@PGD,#W=4d:Y04e3K&37?YE
^(\885cRb.[K4HE-Z2XC8AeVM,P.>8Bd@)=^HD^QW,76HfKSUNb8+,R&G,cF5)&H
4(\bI[5.gONB4/5<LP.1B;1d&IUIRfS8f=:A/c0Ub;2_5(@?LQ=Y8;gY\d);85/S
6<F]+ZGg^G7G]D.?//1Ia7.(W]GQY4+J[#X.V3O/4K]ZZ9W8.BR[b:f;?cRY(]7G
\JUcF2gJY,<=>Vb4cW<9T[5dV4g1ZAE891-<,PBJMeZUb81WLOHbd,QPHII2?+LZ
gfEd0\]C?BH1AGZ3EQF(+@0Z2+04DGfcT=Gce7#Je;e0_7agPI0;c5^^V2\f?E7]
GTCZ>?1RBKQHB@9T0a\SDJ_<dH[b?/[WGNYZ1)55I@3V,3]R-;P)I)fH;@4L)NVX
L)XVG4:^2U.G4)C2:HL&+:9M;>XY_g>#21bCOCT-7\RQZBBZ)R[>SF;DF6L4<d3K
PIAH8J,-fKO.[ZI2QQ..@2L)OZOJ8N/3B:81gX23J9S)ZAGUWgAQYOU>g[eN.=,K
=AKZNd<L@Hb&0PM7RVP0RB;2^9>V[,D^^GfM6_9K1G@L;;\.D4_]06WJSNT#/IF8
>5T>1G-TR3A066N5:XW8@X&DEeDX2R@e]]BCU4V]]@?CA42H92A/@B6GP,1e,THc
CY[QX2IEEdS;d5H\WR^K<ETUH+Z2GSRZ6.3-H3W?]J-.TO3T5V?/(L/^C:_F_UA[
-L<R#]BW_N5[a7AN+]YcB:V(W&AMWb#c9=O\c0#d(4cg^9>#GKOPH#=TL^gL0OQ8
=74QBab9e<aE,<LEJYC@g6+[ZN2Sf<;8R.3FNMFLae8(6Q6OX_:9>bIN-#R((OCe
,S2,7&-Z>O_=T.>FT6QPREH7ecEEMPLJJ]a?+3_5C?ZSWaK8c1:^FRY/2DK\3bb@
Y?.faY9WX396]K<3VPW(7Y2e3+>4C3Pg\YbN-PD..U2PGNbL10,]FA(Be8#3/(\^
K<:M9K(-4JJ[08N-_fKU:.gR=UJE+#c3Q6:bO=C<]c8^CGI^D<2IDELK.cg>:2fN
._BMJTA[=e4OM5>T7V2F;MK-YTRGK>\7@/+a=8&WW3,?9Q]E2H.RHI1I[T\D0Qg,
(&G1V-5J_:0(d&.\b,19AS-/?=>+^AKDL6A-LL#,(W+<=\9U;/\&FOQ(dWW>Y6Z)
.]C/)eRg(Q7)/Q^T#adDJDCDIINMaNVcPcN:D0U<c&[P_2ZIAGM]O+[:.H5R;A=6
9cGXH)93Z#;XeIMMGb1?\E+(<NR4;BGHZBLJ<,)[ZQD]^-,<4/#47-XI197_(d2Y
:<E&CT]Y9Q@XR>4B8AXM2/eG)A(/SfL<:@.W#.ffOFgQBU/0HD/C5\Zc,+78B9]c
E@JEX\8dg@[-QR,1<g.8I_XK^L2PJ7ED:dXBOXS/Y_-]SDG36EB8HGgH4eGJZc;b
<7O+4&W=P<>IM0-G_+cUCV\,(,E8J=;@L_:D2RDA&/_TA;:aX?#@efeKFR0P&][1
4]=UOE\RW.VGIPc-K^4^C_UE=e+5PYgMbc64NA-EW6D4<2,W)f]L1]XILeA2c_1D
BX:H;cIA4,Y/>C:X/_)DQb>5)Kb/R,C:=Y?9[53E+UdXB6;VR97;8#KUYC#\a12J
]I3Z?QAeVJNCbIUf5^(5g^MZGE/R2TQe#\E>a[C:QgW4L8Y@_aRH<(2RdWP4[dD7
C=CK70R&Y]C;.GcQD^H\5ZO=aE]?_RPD:7bH<FWW;A/@I0ScFE03HJ3HYGcH-#:R
[+M:.DVf[/D;V:M<,KZ?VN>0Y>PEFV1T3U>7W:_7:^;62a5N(9cf1;A@12&]&()9
:SEK^[g2]#4+STSBI35AcM>-PF/HG;6aAV>\.1]NI.BWX;WRd[UF=gaRg2dMObM:
#.PA6b<270G;8gASXVQ(\KbDD(?5]9>X+QdB59ZdW+M;GMX9@J[O-IWL,&KKfUb)
OMHg)I)AF>d?a#6+F6[D2)?S>8/bF:31Nc=@a^+5\+0]e-M;24N)0W=Q:V1N_3Y,
[R:D>RB>9/LI,@[GKb;#GgB;B[VD?D5d@Be/)K[_^U78#B,^EG3.SA9;]a,Z?3U?
&&9OfbLY9^VZQ=CZ9DA\A]#CF7=&&1VJLOcVD]aJ2M0-aI1Q14EcDF+RXLFGVZS\
DKR(=>eCMG#.gDfc1AKEUCgS3+>R.Y)1/Y(Z(RJY>M:JfZVXK/E0T3/GKIBPBTa2
<M47PT>e5gA1:b2.LAKb,eGIEe,8_>DQBIU@E?_>1[/YR0=/aE(>QJLM\g_PFb]D
,N-C9@;ScUe1V>GXbC9W;[(K?I4T#FU9RI1YW/gK1KbK2=\;.&I:=<5KOV]b5g1&
e,dY/X]APEJAV89D0d-8SOT\aFJ_g]/,b+_2RTUb#-#3P\GYZ:Fe?>A(+e?d\.>b
E&V]TPc83N]@FJW]GPfXaCCTa^VB^a<3B5Qg91f^e@GFR^E#;13(WLIMeA#5-UTQ
Q-@QP_4&<FfbPeW@T,Z\5@<P(]MT49M<:S?d\5:(UE:WG&-J;3eY,P4J@^FJ3U5V
NENUQD852<;G=W472Y;Ua4)T&HDM8D5LHOf;&J.P/C@[H-L+NETgDYL=L.TWKU=(
5a+G?V#KPW4;BBXKDMZ;0,.OL+@?>S;eWNH8JYI05R=7Z_90T&R,JY(<52C=IOTG
-\&9_G?V^;3.Y6QIS7,9E]@UC[WLJc?/4Dcd5A^[G(L>.15@I(NC8B7Pb@c-1fA-
1E_I,HJ,IL^);KTg=WgS4M(<_@<g;:TGa/7/+8D55Z8;U1>7O7P;b.?SS)6c_Bf1
1f&NX1)4g+\5)5M7-8;<16Hc8aA]&KPGER1<4deJ)3>gcf;B2VPT?[M]IA\-K\QS
d.9<36fSW+RF6SBY9[W4W)#/7D(7U4CU[@ICL1V/8C?]N&0g&NX8@Q(7;&+<ROPC
WZH:cES(Z>3YUaS#52fPA524N2+8c91dZN&M=eR^KHU8.CH1LbBPX#QVg_<+//>:
AdG9D@\ZB+F^#.&JPg)08ZcM5[JD1XeR?>I+>VY#]QQ,WO+X[;F#VGNcddUd(,3a
D(7[D8LVBP5N8S:H2Z0@&Z5G4(^QB/RU)&/fIMAg#;a8/W.eIC)+@G4HO>YYVTTJ
2ETEU<?>8Z.I)T:@[QX\LU/[RTNVCeXTSY[0<9J;#>Zd4cCddZ<Y3VC8d064>N:B
,FQ2J#--:;cX=H@N0LA-VEIXV&fXgaJ1@\#]RO.SWb/VK=L?Sd3U=02A9R:>bbP+
.F-6:D+OGN3RAG9A_<UWdGYEZUJ_[/ZdH3;:G<+S:4a)ZeDZ^M(.,_0J4SbS^4I@
Xa@:GX67EcE0?7B.G>8P==da_L9L-UOKE@3HS002+9J(CbC?6ORZ)&XKIVP[(\^g
=WQ]d]/PT+,\\(.5_J\7K/^V=LC#S[V-?L.8?XcQ3SD-]A3VZ:f)]6BDXTPH<&,6
CMVE6J1QcTQ8H:=M;+>QX0O0CD_C)D=Q-RFaK-SC[WQG[]<K2:C#FY)I1IXTWfE0
-a)6eW<bZW=3^#;RL8SVBR=S\T6L93C@XT2ET.-^efE[_6::M@WV6Ca=9FEe:G90
UHDZ:Y-+bGdQINE/M:0YO6DW:e&fVO4S/Tg2<YacCKRANa>#1]bM1(N&51W<_=16
ZJO+d9=4\,HVC5[PAbM@H\^TYLBHDGaTS(]I]/BLR#?>WA8_Aa0&\^>47L^L=c82
gQ@--^S/_bS19F^860GaLBXH>bdQ^8W<<4I-+&)2_V;KB)7V(95\;&Pcf;B-8DF4
INS7+,:9P\J_?RI,0D)Q?#-/TKa/ESODIQ,X#TMc.MR1S>BVDTA3^+&W9(B<A4XY
<e<X]F<dE+^Ed^:]\J2SZ#2Y_HQ&bRAF@27&522&DdJQY.]506.Tb6@+M4E#Q-PV
@8RQ.Dg?@JFdcE)/D-@2JN(.K144[8:8VfWJ<]MI(g;^8aB&-Y=1_A:+Ee5OV0b>
bYff[eB9;cD4?^1CKG@5=Ig5(5>VJJ__P^LA@XK3L2cB8.<CXa0(E86;&GRU;DJ?
\,1c7;2RL84=d(J/<5.Zfg8)HL3;K^[]8C&X<?^I@TR30(bFSLF._>#2=#>aQ9Y7
H>F<Maa/<#8;^VU9&OF,<If=W4d^S(@GL]G?fGO=U-MXZ(aPdUFf>eGZ.8,[PR=<
NA(3,4LUB880C.@EFG69IDV?(5:Y1_KfcG7JZE+JBb6PT(A4UNHdcd(0]F+?FbSN
:,U1b,B2E--c4Y12B?A?2ZeTbLYLG3C]8324MXDe^D)Y.N:ZUA&BB/dUK)/@MG?&
N^-ga=&^K<)<Z):2Q&PdY]EY-2B:S-EWV>C-8Id#XBTS4\,?=:H]b=T4B1R<e?T_
OdG<;,9Z(9+LNJb.@Hg2D#TGP@I^8V\X6d83I\g)bTX]TWN6&P+V)YC_gb<38X6e
6WgP[APGPMQ;N/HZM+KW0d6MV4.E^E8LgO,18a>ePSI4_<=f=M=JWF>gH-,H/H/B
O>;I#K9Z7bIPXSd3X.Q,0QR;=gI.SAPJ=cNdAZR6GY>NL=HTJg8@AYP9ONE&QJ>.
\QZJS9&:OaA-&;7^Mb608\6H02,F4^<Nd18?=3>E4THXYH,Fe:8e+W65+ZM34a0@
33]URE?\,_Z/Ff7ZNMEA>;>B51PY,^\fHG8R3W(Y(f73U;Gee3f2VOB>6Q4bM[?7
]-<R>C]a3ZKa(g_F@:e6D8M^1+H_(<S5UX]-&NRR70]e6=@cH#G)CA5f)I<ZS:eX
IeGL/71:-F4S[e)SMWSgK;.Z&W)YENA1XE[8\CZ)@:UQYG]S#+&NI:WJc5X/J0D2
X=0aN2c8_8geX[F_&[JVAXZT1A_OeV^XG/@=MA>a,.G38[XTYL@8T-1d-M]H7TGa
XIM&5;>#bE;f)_g#Q0Fd_N),WG+S^+aJVK-2J+F#)O[0+eD_gJ#P?A(^fLeSI?81
+76\X-H:,;7bXc)-2UD?&WQ&>KeCO[7,S=;faP]2<I,6=>_]:.&Te_W0a[fEdA)D
W[/[)MP39_3D6d#HRD\1c/;,.-^a+@<P8G7A[A[<1LCVg@(JH+fZJWF+V5=,.2;T
DC<FZ[QZfF0(9N?4BNeHE(ID.+S2Xb,,JK.gOB7[+2Fb3Q=g/FEMQPU)T59&@<8Z
UOH?:626K8\3R&H.H<=g@+gd-F+7fSMGHd.DD31G]F-_1eEC4FFKNaf.LA6#.<QG
_DOS@6f(f]\57<-DK5gaV4JTX,X,Oe^f(R,Y0GcE5WD#XZ(A1\-=.78N,9-;.)6/
D&.)WPMB69QFe(1J\;>6YL>A2.76YFGI0DSWa^Q(+,=ATZ90eDI@?P_^UP+,<6/=
;UfX70/L,S2N2CIF0EbgS0BdfTT07f]Xf,U.#=@#V)XO]#AV.]+O18K#cZ)J6YMP
X7O<8dHH9+>eM?N]ZPd(4(>1&bZGT0A;SQ9b2\A0^(J;_]aH(N+0/G[;KC2J<SGK
:A(aZE_1C7GYdUR>O6A/7bP@VT:ZU3f6(QS5#;]LGFc/I7Da/E+).\_HMKY@dFVd
ADf>.dYed+)IQ\G#759M&3Y)8SJARWBg_d0eYdcPf<LERb:[H7W^WbDVc8c^;K#c
.SD)gLN2S6b/MPEPU[-Q\0F/=B#bGX91JW1+VC[fc4ebb7,_ZaP40]bK<QMeYARA
:]+?P,YBdbD=;)I.6O##Y[I/,UX<\cG[c4;g.KZAXd>EIKe5;c;;Y>eJg-)Dd+7<
Pf3[U(7VOUISP\4gO8&=M[QL9b)a>^^a(XaX[e9/=\0P@]6X&(LTQHfT3AB>Z.6#
63Z>9(/63Zf.C5:AcB<\Xa^I@AA9AMPT9&,@52@N:FHd+.aI9e)_R>9,\DL1]XFX
6I0S<ZHR1[X#90G7QZ+16UZK3YNUWBY++G@g0<MHb\a68K^fd#33T+K#3K;]S>K6
ZPBW;YccJ&D-#]\Md,,H-R,ZB4-WF8L=c3GAZV:^_196I21UDGDFPSF2\>,SNDEY
((H=)bP3L@#JIY)0&)VT#,YINbU10F2/_KYKDMV2(:2EQS54?#]YZD6aGaMV.0R3
8eC7&GLMB8CR>R5VO/fE,]4bCSN5JKf\.Yb14Z@FR,,ScVC/DM.WaeO^&[D]U&2a
4<a?E+adWaQdA>0T4C1B8(b9^g+PE4:U(JLeMMK;NVJV8&C[6<S#f&-LZXD]C-,(
27E&.I;D\2f,+4<T-OR(?)/HA+\T0)PS/3(aI+e\Qe/AF-G\SR(N1[B/(9X=U-fN
97(+,a79W^+F4Y4()@f9U0X(b#,#T6X9Zd9/Y2Wgd\1)_:9VP204eYX&R(S\ZYL5
9J;1-=&J1BO9d]NV:;I8S&?1N=M]0@a1f#VVZ[M4,?A5K]FTIZeN5.^A55Q<LG6I
:>>4He7f<aY/0#ZY)cgPIG)#ZV=AWPW-CC6<-NWYX<eY3\37:S0gaT._Q(?LEb+U
^LcF(1U)d+eO.)33ZFYO@f5I@6aSL=2F:TI&89eDD4OD3IA5D,+.a?QTdA)MR>=I
1;<,OUd829]WEEb,Vd3a>JHM26M6L2\UDPV+5bETY167/Z:-4+]IO0]R_YRYMT,D
baT>[=B4=]dX4ITWECDC+(J._aL)22d?dVCFWOBBbK36VF]N3DH=/+VQE2>QU^6J
25?^eS8A5<XG^3XAH5+P,G^-1/DBJ-;_f)FN;,89G5L2A>\G]PZQ^cQV8XV\B7_V
8=35cPD>@aU0B^;5X:TM<4GLQXaY9Ff8+aU\Le_KTLVW97Q)=Z=gLddUL.Z\:VBQ
bf)O_BX(]&E37#[^ZL@EK\^FN[4/,-KBMP8V3/<NNZ5c\S?B(&<3N8gC<FC1+:-M
3&a4R52V0H90V#+X]?S^NcT_LSSbAK+XgIVVNJ.=+#F0A_?-eS,f@X/PcR4OG(-#
Hd>V#A@W28+LPCaL<2c9+,d>6U2Z__U]c@FC]YEGW>XFXH>J/0V0SB&-&\PU/Q]g
T+T49g51,cR5(2@YK5gNU?+d6dGF9N^fV.V+D=&Ga=9W47.YRKWTeD7D:g\fJ<^-
\>#Q&b.I;63EGFg^F&=CJ_b3bQ6Re<<U[3W58,;:SCe+)02Y=?07<.2,<^IJG?CO
a;]I&H6@+4@<)IaYP[?B<=RLe>CRLYH1^_RM&/R4.9#](fC3T3)]eO<])#43,fQL
S:L\@g;W?8<6-JZfXY20F^>D+6U&+W=EWB#D74gJ>1-7eZ@e+EF=8]fAH,U<2]B+
,Oa>L8W6.S2&Ya\4G:=)[@/K@T\+_/3ETFFVHL@4VN+7OY.V1R1-WA,&a5TdgSI7
0F@<f#g52^.2JU.0I01:g-[4cc(SWNWCAP59L9MJZfB=^M+@.I2FQA>Wb8J\\BEG
/e8F6HHL_R)#eA0]-[71/I3:1=g:NZ<EFVY<cB/1/5V;XLaM.S+7,[JAH7D__UHQ
H=PNL11.Ug,f=6_WNHQG5FB5(P+1QaE9De_H&R0(&^9?dg74g1.B)MVT,W/-TYOF
4-7O+-TbC:B0BVANd[@4RSe6:-H\:&b:gfJ.3a..+DRGe.OKA1\:L50V29\(dDOd
D-edK=)4Ac/8=bdJ,R>-^[[[3#T<,e-cR,FB4P3cd5UA8DeIO&>3FOCZU)==a?b>
8dGPbe.>WX30PbYPUe<0?ZW:)JUQBJ];g(f?:8bba.[8cB)\PM^1E8U,FE@/I+]E
-?HfHX@@+0dK0+:W.,?CeeLI-&1Y-+67MKSN>X&cGZ6&E;OYBNHVNfg)>NQ9<C#a
AK93WcPM2N?Y/0,[U#Y:GgA_Q8WVX:cNcd4<Z,X1dGEf0K6/22g3:J:cD+gXPZ#g
7I7bfE#Ac5fbJREM>KZ@<cAN:(.I3Ma=+Eb2MRH>O7<9?1)M/_&^A3-0._Y[AZYW
RRR;1X;TX[OHN-_C:.fBd@TTb2L]TQf<FaAD6R^E#1Q].KVb7Z9;0f@:e&_QNMa-
=K6Xd>1CNF=@6MKZ<:3;WA@Gdc7c>[<DWJT9EcU(cXU]<0f-(dLS+SOX)9KODN@2
0SP@S=)d-U+Q8;[Va-e.,P9QL2gagS4G.6+G<Nf2&Wf\T+?Yb],1N-2<eE+E6O;^
9QF#E5<X=4Td>\KUMYf=PMGJMI0)YY-NE(@U4J3WD7/YASWS5DV-D\g_DT<:(#GM
_@VANeP_D6\fYJ:W-@2(3::QMO;W)G2Mf7@Ze0Y#dg@CZLVLL]<2N;He2RL:9NdP
[aI:5I/^#@MK?L)Fb7afZK_E^#:?+/_G@^CYBC;d.IOeZ>J[EWXZ?GZ.Q[0a-_BI
_IDIBaZAPN1d4J]);\d#JK;<d]2P):-6&W/TBJ4/<[e[5(7I0DNH\K/RAW1UVC0a
55C_.3:.C_f^^C<1ZD04I6S:681F)V+D>;QP=E(b9c#Y_9O;^I,LEC-)U_B2,4,+
X9;I/@a8HRW<?=7A,E=b>VYW[.::d+<R1E;)>]9:]4C#(4+gHIYA/.S\_1f7?Md^
)7U6JQ7_,8@eU@?[N+J&)TH:O3a4&(bd4cS8BXMe0HQ<:P@0U])V(DSP,1)/WL0L
>W55FcH+MeBcbJV_M)Z[bNDP]_A;R,-6LSQ4gDTgYWFK_;6Zc4LW.:PU+aH_IQb5
>S\.W4,S^,S8]0Z.1g=4J+&YZSeO5feVJ2S(:AY?G>ZL\3PQGY=PX9M?N:3EF(V(
IA;+eKY(dA3_)365I0ZX8bH62faE6&&][UD@L703=@S_(:LR)<_]g?[SgW/FIfC<
HYgR<BeC4R<g3,gbS5W0_B+a20L#&3@MGD:OT]BTc>48JM[QGeI,\eCW2g@-MXZ@
I4JCgcF=0f+\Ma.9Dc7[-Ve#S(J/&Q@YFRa)-+N(f811H\1>CR#C0<SLeLOL\d31
LF.X^?>(:W6F0[@1b:Pf-f](Dc=C^=EL)LKSc/MBPaE,bJS2C2b:(a:I;\\(=]Y)
W8M1#D&bORLLf?C(F0A,,H(f-5#BQD&cVY6&fA1\<(06M:/R_F?FZb2CSE>:N8UH
J0YW.&OWX#^Y>QG(f0ZOeEDWF:I^TC:4b)^2=M3IPJVWZRG&;AVK\EC6#;(YOF82
U9T,9P)3?[R;TQ08HdIMB3;=CCN+;7<E\F)YT8e5eKf<][LVZU+F36X3)ROZ-f1P
>;J/eeZP>7>fA&/N>0W6T].SQ=TLZ+OLYJbcX0YYQ0O/^RJS8-Mea3(CcD)30(E,
Z15P726VH?\S;-#RZCF(d;@7b1VgXY7_7[2dTe/B^[&CV8UWF2c>9[+QRYD4f^1>
HIK/I8_[8Q\UI>5O7CPe97+?X04e@LGA>2BVDEDg5)K@GD\d@8@9;XP9XNZE/VdO
+0)N7-\87T&dWe>>eAV>.CDHgb.DL@]Q@8)Ce5?U:)97F]Z:(?-fWEeBQAKb7,M.
5E1-OD19:G+#Y@<JZT-:adE8,9OD8Y-&eMdC1Jf3>J>(Y2XMa]MQ4)Y+9^&LC+F[
/4I\IY5YY]&)Z?>DHS4L\f2b<eg>M>P7A_eINWKWFbD?S7?-7B_M7.XI4],+([EU
CI[_JU&J#\TP8I-)(S<L@aW9g((MRM?ZC+g0)G-X3\B#bd/^N^/.W2fO,,/UW:B3
cCf-&ZKE;I54UF=)Z.M/,94A_ALg)S-=TI:AKSVb^WV)^f04<T#P22B(9c0V9Z=W
>Z4D-EOV-=+fY]W;E/dOZHZ=dC^cK6B;c(VS\)a9AQHKe0^X)@G8D]eKH.8bJc)A
,Oc#baTKN8/QfN3]-Uc+:J0=3b1:gYK2WIf4Da6Jf^]>:G^8AP3VVaS2e]&@fF-E
9EX6P,b3RgC>c]g(A4:M85E2.C[XMB+[.3HA,HUE[&,A1CAQA3g2D)BKW;X&5][T
@4/QQgC_PU)Z9VF7fC-Q7Rf[d]JdX.PJAAS+7a]Z2G5YP3@02d4SWO6K5L>K?\_7
0=(MGgL#>W/8RJ1OV:83[dPKHLO)JfGA3#5b#&?NAbfU5PYRL]I>Z8cL&6-S.e-8
:BeFRBd?g2@@gM7?I4IgF2FOI/,1)+P5=IR1<+0>I@b7O7T=#&U^)O2IC=8<Uc8P
X+C=#,Ie63&\<.VU>R^<J+ePURRI.;b^@T,IUU+B-RR,-B7+,A@7_(U:Y1O<g7Y/
d0M+?<RH-4.PCfeOCNaJ-A/17MW\#;Y9Db#=2P1@Q>U>PWbIQ,ae\G54=Q7/YKeY
Qa/fQAUJC),17O.O\ccb[b.LZQLEJO2a[YS]=.TVXbH<5H)gUXSJMXg2567VgK0\
:B3[P6C9EV]T1dC;33F1OR8XR-_4^OI)PZO3K4TLW/36K^NU67b.4L41UdU+OK]#
OeQ(0QRF(L2U7Q^3R\9R73QIfE,],W)CRQD^8J_9H]af/I;KQGFA6BV\0+;eNK<.
d3+6TWF-248&VR7#1&bICU;[3AK<bYa\1gOQcUe\9aG+=V<7Cbb:QVQIWf5cQI@V
KML^PUU3\E71FWC>QfO9:PfB)8FA@54+@BF3P7H-E^TFKDFZ62;3F.K:<V,=CV+1
D#A.43+X^GZ[9TK53ZMZ3:OIg52gW=/_//U&90b)6S(,?/.EZ2aR9Nb:?T.d#cIR
fBd-4;@1.,(/B6a#0.[L9dFDX0Uf?YPO:c064<[JC@0,)]?f-B1QCge[Z_>EF>9J
0;#JWBZBY>DPaa_/Ue3Q.I^&AI1g=)KaJ=B#I>L/E#?^.8RP72>g96;&30FH.6Kc
<;Af\2<_GCe[CENP0.PL+Zf0,I-@gQ<ST7[Z/YT3D.SFUedWTbS7GZW-:@5FJ6]U
X^/.J<>429=c&0;#LC(G=XNTX)49U9E<6OA0USe)[GQY#?DE3+[N9<M5&8I<L4G=
EXd)bTN[_,c>dgF+e&9:fKQU08dQNOfBM/FaMbRR+#IQA:\M33P/V8M\QG,b-56H
c?X;/05V=&EcXFU.M?;6^7aS7_T4D<]F@-LE^=11Y[DOc4NTNRUW-[>&fR)P_I0J
e4,^HdM2C/OQ:1.93/XY?\>>1_-K<7fQTXO(:5\=3Y/Z]Y=TV<HcFeC8gLc)?),N
++9,?/@,A;9MT.=I:LX8FeS8aE9J_8OD5R\T,_L[7-bP/b]Va-PR[T^PMB591fJ(
\>E+.OM4@T2MX.C8944SD+YRC5+4=cD)g8D8K0R+RCGF)523B,8JUG@KVN;.\?eY
FbNRS3A1;d&54[MI0&6[3ER#^#N]@gSUB.T,6HbMW,>T<&3b1g+U)N\GIW302N2/
,6XPff1dL2+Q;LG9^KW]a#O1XIJAHGc@(U?a;TGZg+E-6c=RNL?XX4UJEQ#Q6eRb
5[MeFPe+>:C#&;VPM4?;WA&=](1QRM7FJ+BO>Y<Y\N-A;C#T6Wf0ZBY^Q?-PLNL3
U5;]@f98UT^,E\3=2#OU)=c.e2PRTB9/[RXZ.@^Z>A]/#@3@SLF3HL+3:733BDMP
Od9&\K<@81OOYf(6T9,GW8V_)7G(_7)NeL^(;gOF9THZ_YRD-L42Z03N;_dWPZ2L
1)W9^G-cPL._9A(DZ;<WXA,S_:.UVZcXL8eL\1#N,Vg3;YMWXe,;-#C5X3N1_g.I
aGc.<A>^L-=Q<7D^7S;Q.>U#8afTgKCQ(\DLfcJcGeLBd>&5N(85.3CZ@b8#43Se
VVOM-UR)&Y=eDX\=?gH?C:c)EBXK_,;#MT0-FWab^<[A/M@adbU4AIcSA?)fQdYg
07NFZ)1b(&ZG+&P-[2PMD:AKW^Fc=d;5,E_a]KUS^>YOBU;R]J:=#,HE^O5L6#H6
gUDCfcH[1f[P4+2=g5C7N6>X1YcR0J>Z1JSLA]\A<Jc_Dg3RdPG>:LG</&N&+7V?
W7Z.Xc\WZJP7Y+N7:@=]\AR,(3LW@FF]6c_<d_-S.F4XB2ABT#EfDUe0Y;.T(34=
Q6^O,+]I</0QC@#Je9Ad6NW#].C/IHT=20YHI,FISdIEeZ7-JcM[eL5Y+W)]7<?2
Q]ATQNX=0]U&2&E<(4Vc+QD42f[]LbV(QZeQ:a91@(,=e2;F^70MGNN+,Xd2=FTU
^Q,Z^I9;ga3^4YdKZ@:C4Jg7e7#R8O,&34ff1bLc0TaR&dBd,&]XTSE(U1KU^&^J
A;.VUaRTBdf?XU\TL,&;FVWZJDW:KJHdLf61(>JdC9\d4VM(L=8<)d<I)+d#PU_[
7KaNJ0IF)+\C5R.;0H#U_V97PF:([35),M9LE\LP3bT2e0PG&H\VV(KE4^>F,])7
^HP@C;L#4]7AYL_3d<)D)g7<Zb5(,_B(:Sf4NP4d8@RQO(gA3WPP>S+V?>,[07L0
@6I#K8W6c99K0+R=PIOWb:GA6eA2QSOTd6BVY81-9S.Q:?SI9>,NU#IIf830d+8f
6Pe@V#/NHVN7c#F-=ASUAW[,/FH:-[^V<Z[)A1.S5K55+:>b<[MDb:O-,?1G8HQN
f&@,CN[3F>7#V]OOD-SN+UTO=)c?(Sd6g^A-FCFYA-Z^G[T]0[CaN+]GC(_(gC@I
Q;@9Q]/K1#7(-,&;Q^>YPD0>3(=JP\>+?ff]bD^&RX3?(QI<Wg]U;93R\_Q9YOe[
JUd=WT]+YZI-2;4eSfBK]L-.O\#.0Q3#Z0[=gV(QJ8_O0BgA#^3cYM[^bOW^^-I.
:P\bM)LbKFfT+4G#KBOc>75>T,BHc/ZS^E[^OCDC/HXE=6SRY2bUB0adY)+4Ica8
f(QH_2<L6NGGgK+)eTM11NSS0MY=5cKTTaNgT:ZJ5P)VM_H?AOOO)0GB_#Q3MdF,
?4.fc.P_O.fYE=GgWO-<^PC:/K#2?F2FF7f;[0/_AB>+]XaX5g=C=E_(TYg48W_)
\2_B(I=-,&P,5Y[5(9QF&a;a\eRJ4\dRMDGb6H7JM4GSeI?)b7LRbXJ(N:C5RV/7
d8>Uf,G/]IRJ2L.B;<\[C^UU^1@&NG4XXM?4bV^SZWJHd\_OKa&(3cTIN5AIO3f/
d)@+1SCe51(37aa7-KK,69Oc-=Y=AAb1b[@HCN<aU0<aE/Lf2Ug^geW(XL(\=ZI#
O:B@W-6];3J@[SS>NW5L)6<HIKFC_H-PD-7.:1GSL>-I>7S3:[3ACC&(dP9KG#PZ
B+JeKLgEPHc05I3Hc,90T<BZf/>EV@-LK(#XW[_-).)EO?^^Kf<,Q-D7EB6@g#Sf
/0[C;^HTNab+AcJ;AIV<XE0[6F0e.N.+0H<)@.A)E90>b,3?<_+/:5-+15QOU@OT
STV7,+RZ&<K5\J8>Y=;W8<.FG0NES7W)4V1I;-X#Q+Fb?ZMN213EXa/\NK#V</,3
Y[?&D5>&&MF(YA@cPL/[Jg5J+d>L;EUGZWe/@J>-LZ,T6N8f9e5G3G^-NW(6?13^
I&#(J(]GX&_6^K[Y3=J:Cf\X;]DJCDb2T5?DM&V.I1D-=01_##4UIEeI46Q+?4()
NV9;O^K\]eN7N?UF.V62dG0@].5/_P=<aaL;E]B?Ig(V;:XL.<2#A2UBN[_W.,X/
Q\4\TDBdEMRGS]4Na.AF@Fd]&]BMNa?D]PAKKXF4]DMAJA_VFUS?M&]ebId_QK+C
=XIJMSZ,26[T-C^?.;3NU;9;]+6@>Y1?Gf-4(\DCXCHUC5WNc2TaB:P3@MRN::/d
^^cFDIa;.e(I2K#1V/O8gL]2_b\ER8I09d02ZIc/X,X;FKC;-9:0PZ;LHX&#G)C?
P.HEZ&;+X#3KgDV)4G?d,IKV?6Of1A3>Q8&ec^GF.&:QfDY@]Hf>cH0DC^N>C][&
X;OeL/QgZMe6fIL,<2BHW8aGVGHf2B)L@20+#][6b<?AG6=[IXBR=dZ)._2FdfHB
.D[,M+bg5b<R0G^LCT+IUg-;X55+TO4=D_>VbYP6AYRfR,c<(<eS&KPa)@P@,;LU
_EX[>e\(ZUK(gCKY?^>9)-W==ILF.2;B&8GV-MCAOXdG>beR\G6d9\;E1+4C]#9?
BUWBb/+c8B-C8(NZT<7UTDE3,682,GCB0/8HP]LgBDKfe>aRAc@3&S3T/bXZE]P^
[DF1eV&GJNcM5)2\b[-7Leg@Y#UPT1_LVO9NOCF5]LLMaUTI@DD?BHcVF4,5b]2H
+B?9b;EE9dSG/+dCYG#IX>;=-g.\Q(4FbSX<E&7NDCUAPfeO#,C\=I<==.;.4e[0
JIfaG6].1aR.@SdLU+[T_>&<;H6U&T-6PJT&C5bH]79Y\MfR_FHWP_e#Y[YcNZRU
LI[548(fIU<Y<2J/ZQ#[39AgNLdENYLU5WH#7?&/MJE2G2)NE<,aLfMS(>Ne@A?4
c\&Y_aYH+1b:+SSB349cZDD^SW\<U(dVT0&&5[Vc^G>_^3/=A:C[dd5<Z&YdJbVB
T@6cRe0fT]^3(GVY_W)=?VG3X+,LEWdJUO>1Ca27DQM>KS&Ia(^Y403LZQJg/7M<
[)#f#6a&]&^fBbTSHQT&;=S7+#OT4A+Hd.VgM2+5?K<=bUW4I_+&)GZB.?N2B0.(
72+OO4GPCX@UZeT\6@a#+1>Be^e@32>W@@:FDJ75/?A<c[WSEO66RG<M:)M#Q##;
,AE\74B0Jea9:4_#?VcLE+ZHW=E[VJPI772/+KY6,[f8:gZ;YR8g+a.A^I(-19V@
[D(^\K#[[/[YB[A(#1g)b\+f592+D4R(_d9gFNKW)4QSaP1gIIQ(LGb@XO].)a>.
W4DLCRZ5:,D&O_P9>fa51e]75_V31cN\d#IC\F:^gVYfC@<P2U@4f[?J4):.7IKX
US9\(M-[Pb8G:cCCdN74K9d1?]4Gcb]TO.+>^4bKU@U]LQJ>K\&T:RK#D29[CO(8
0d_QCc<fH]1[SZfWLZBUJD5J/NE;7/QT,3F)(SVL[4+.OGOS)aGWNU>Q9LE)<Vgf
N1GNZ\E35922<@;MIVY)=gPTO785-W:eXEUeLT(<5,40[f6Q+OJ;B00/WP2,_f)H
\Y-YC-80T5A;cT]A:e]I]P<a,G+FLP(A<#);/KHZ:D)A#F_4NWg<HJ6UA+&I<9;D
8Z]24X#G6YPIN;;PUe6#F2JJb_@J(T-L\)1I(dTTa8Hd2L+ZS&1_<,ZNcTL&M43C
1BaE<4EDQ4UQU^CR2>=7;)1b3MdUGefC&SEURGJW4VFZK2Z>)BM4:K/aeHWWb&3H
c,W?5@&Y_0Y10N^FA)_I7L9Y_;=f?FOc-W[D37f&96O3A[@7]0#R-_>g.:<?>N+_
O5HRUZS(IN;]WdDR<+@F=IGT,0d5_R(/D-6E0e[=Qd,,Q\Ba)I#a<WFN=TIKMZ^J
Qe(;SQWc<]H0QF/;5]^K,LO\OOg,V\fFO:=YK59a(/-ef7MT]&/G>7U]\Lc:Q])/
3T>+?ggAATT<-ZZ/TN)aG35PVA=Q/.c4UR?-W9Q/+/_0=4@XUd+?YOD;MXASSFK8
0LSX?ABK1]Of2/4938cEKO.TWIJR[ZWf-19^IDf;e-J>WcB\/@),^fP7-J#I3[Sa
TK_;c(]BRX<_7/7:5#\0XQ94;Sg0Lc0/[.1>5Q4DK#b&;,C[WFP+\)e8]6A?Gc[Q
9f7HTO5FJE=2.;(4E.3gA?Pe31eV;@WSE>a/E&cXD\Q3eZfK.>K\.5I>LL71_@\L
PZV4^eC:)H[J_,MTafTg.,.?@X@8QI^LN33CNeV(/4_NNN,^6[d+/I8,DY:^^Xd.
4J<YG6L+@H1d)UYM[=V5YLAKJ,9_0CPEKQ.RQ2P?_PQ7K[0KDQP2L&]6NA3f1?.D
&=#O-/dH1#Ud37XVYG:dP8aLLO]Tb1ULN.fBFcCA^CBf]H_:K^dS)ZDCX82&4/J5
AA)?2EO+\SDE/_aPa+fKE=?gcFS^LM#AS??A/\TD1Z^aCBY+\,AfR^W_e&aE8T/[
5H]Ef1?4f++A?d=g<B=-@;fcZZ+.d[)HFOAQO];)QJSKP2I+K[]Y4H@R3JbF1TZ2
ICbYS/TOQ,]#V)]_E@\;>M+Bc6;\A:]Pc>Q@:7,JKJf8AU7#aS1N/S,K7NDG,4L#
4G;Zg9<F1N9UK58-M(XM)/E0SH69?WLfIJdegK]4I5([I4.+VS1N.<[V4D2]0Q-M
&]BH3IS^<:?YU6#XcD6;T3(PfdO^fd4DKYf8AV@8SYCO<0BUR,g-+^MJ0GY@+(S;
VYKZa4<3P,/PS[dZcdFO8:c@?.YXAV:M3Td,+SQSSH6Y4#BCF.>_2+8,7]<]gVWU
KceE8Z@+JRg>Y0(HPF66f@+,DX7O-Lg5c&bH4C^cO<4/gI:^MaC5f5BJ3fD.4Ec[
S[/e)CV/gge->ZD&R\B^&f6#Q@OgN<d=;NOb0YDR&-LHacW7OGMMQ8P[C=JLb^CP
Z.@Vb32Wd#>e9;acO0H)97^=bDT0caAU5AN33>Te#+DEWX2J^@XH)W_e,FRY\)OD
O?R3PTO)a-CS5+4-5Z,92]-4/c)2-[+b_<ROa0>R4M,-J,&bf@-V[>MY&<bGSaA#
FRCE?24]d5QDb(]Ng)-QN2M<Lc)FT(^AbOMZ+SGRVI5(I75>Y=HWB+g#1U4MU?9O
Xg42]aIFW:I#[K>bNcAO9TVJTP[c2QNYbNBB<.ASb@TUgDOI<52,XNP=CG\c4/J@
2>N>LC<bJ)J]F#<UMF;8OU@BDLO.[d(L+,]fZ2F7ebT@A+1U)LEa0JIW&>If(U8S
,3L_:7BZ85e/MOg(FT]X&:(B^\MGgBV>fK^GN13?;V.&WU^<BE_M;fFa1N.:,0df
Z7geZ@,&B:NBHEYe:)9CWY@G)/.B9A\ZQ3<<2cW;+-_X/[NL>,,MI]<<-a<aAZ4<
G7Pc9D_W<9P=E>-NL]DL:@YH^GG#NO],g/>1=J\gabH1[45_KD1B\c?UZWE/,#>S
IM\LZQf9#b=7f_X:X:G((Z/&U0(N05&Id/7FM\ed=[aD0UM1[Ad:FD^C>)F+5W[T
)#UK>>U.dC4T<NE>\Sa3,-1ZZ04G[:b.MRPd)b@IG4PHUM-)O\453<O^OeX^(I[M
43KE.?aE;cMG^H2+S,\+/QGe]]]dK@&R2/N1#F1B.S6[7E]&6T8HC+\<106@QGB/
USSFC+E2ICQ1b>f8=#9aJ4,K#^NG?S3Cf8.T0eV/SN?.J.LI:.ZX&X8YTZ1V<4M7
(RWe[(:8Uac;dPAQ;03KA,\2(>L]=;FLS\H-DFX2eP+CecR-V]0F5]X2C9E@aE7R
?[6:Za[EK-PY\1Y:aC:9-1Z/4)-+M[3BS;JKFCZU_IC+</G:GZbLR-I\-3=P(\Y:
abK6U,KgE?1LK-HC4EO2]6^R3U)CE7O^BaYU,YN@VEaG.D_9C;1e66#>.@?C#7IE
_S0QeZ,S^dE9_M7_M4d@\N-X\>9,V->4Y=-_Ng1^QCQC[MafY,@+\WA7g=I(-QCU
bPN+ERMHD69>CYWYUFd-W5/01N=A(dL(K0H4YeEYd;^R5L&A-#+#-cIAg?QR@5(]
5BM]cDY56T8M@Z(DQ+X+OR_\XB-8A+2=SJ:X.D3M_8-U);]8@AT:b7c5,feDD-DO
bE4?eAHTP-1++ff&(C;S#f^X6TeY(cOAd>JYPZadVe2]deRAILbLF>6YFHL.4XGB
2#<9R\_YQ?_H+d&2A3&6(;[O?M(L29>dJ;A01]_T(VK_YacS:YKTUeQ9^g0]^c3D
C<;a6_N[@+HYCRHDH.U;&PPOW#JC]\+QVVS;X^<K,fP8&>YK+8LMKE:8aRa)3gBQ
HT;d^7?7c[98ZFPW&Jg,\=aUJPZ]JC;:R^C>#Q7U&WEGD961HC.AbI_,FT6,XY\d
6RHVeNb.3:&5>LWCbKM4>eID0)d,U9Ib.D.(YS-)JKD_0SNPI3Z3O</DfI;GGHV0
SL@>Oc7.FIb,J@\-GLbI-Xe1U8HV8<43c]L+K:1+e#_0T5Je<:HEZCXXG:bE-7^3
6UeNL616Af;@SA1\2:Pb5TBPX57F&Q/HFLUIL-S?&X7d#34I8+]Y:Z.GRDX.G)V;
=<1]&?M4158fZS\/PK4>/b:(K[Y(^f..A;T?^,b.GFLZK)J,BcLC)eR/d(c9+S1E
)eS6ZMZ1,1-eEZPS1<f/:(?O=7EeTWSSH<-(f>PX0L>Cg?NL?aCCg>b;<XK5VgQN
Gd&(.QEU5e9g80-FJZRRMR:;F43\.?#a5NC]8MN#=[&,[(>]+1^B-6ASGc]b4EA@
BF^g9+5\?FW8^MBQ@,O1D^G\CL,/W.IgY6W8M(2)R^d,6D#WaW3fA:a6=T+43c4D
T<b>99IP9FDS<e-0P\?0@\:(d_cLSXPC0c+@Ba;e-e?>d3N/:L)3,8Sf(ZH8@Z:R
^BDYR1P(7(af:_+HB;MTC2ZZK9?YNaRN59PXT,@=b1F7&U:)6D\Ffa,,\5AWC]::
eeQe4TUGa=)JaVTeDW@T=3Q7IUc@8;7LTZ0UQ;4A&:90F\02H)Peb(9a?O1QLM^+
H?KZgFF\)N5,E/AMV0/5EHEN77>0A2eV.gG6&A@]1#-a/5:V;/N1R=[C9P4dRbXd
8H<ODI#]16^?3]&G0/,RO;[Ic4\IgU]eVH5V(HaZgH]AWSG?AU-&?B:cA<3#43#T
=H-Q&?gRc+gL@SB^,SH/Fe,ZE[\6L1[bI,Ig4LY4).\<=IP/bCaRB98W/3fE?H@)
@^\a=;<@J-Z1<:.<1<-QK9b0_?WAFfN;/@)SVZ]_&0-H>T_PQg5;(C8?OP8J[.A&
__GB+2&?8-N0=Y(4(<ZV[cJc\+D8R59V(If6AN8e,28&bJTX[(7aWB3,,2-F/g1&
C2?ge&.d].Lg2<+IRI2c\FAa1;IK]bVXFf>##DO)6:7MCSC-:/+/J8<JT-857.AY
:3TfX9f16c86<5&]]9^fTOb5)-R2C76JYY7.</2]J()[d42I32G+<QYMT>:d8+a+
[[K&O)9a=?;G=IP3AP))M1:\Q#eMQ)&WaM]YMQ_C&#_ZN1<c8#(>A5W6O9+S1L)>
O^\4A0\(9A5^_>KWd:A&JKIB?J2a<9Q>670>)0cZKX9bWZ/_Z3F\FR:W/QK@Qb5#
a9GM[gCRa(GgO@G7JAAd5_-MCcGOeLJ7-;/M&][];+c<M@>-J0ZRRBQ7>Q9+LPf_
O##cQ?RP3PGfNVUV_[U4f4,07gLS9\ac(TS+.1_3_]J#=HLg5&CX<F#3KS\/P9KZ
1Sg@E5,]^4F.<66;6=;+7BYbJObIC@gENHH-6g8/-H&TSFZ:.0+IUB>OE?-13e94
5/ba>?gAAVQgdd1UbEELeC12J9Mf&b-&ZJSKQE&bH/\/MVe:@\?D53\Uf:#^29++
Y&JOZ(2)IH^AE921^5&cPDZA1KAg2CQ477YITCWOOYFb49[F66M1eAD0=TW[2K&H
IK:.1]6G9\3L1VQW1/6(,=<eZHG[L\f2EM7\U,]5)gU&M)7#)85bNfa]D?ZZ4cB?
AFX?L0Y\H)/]c:f@O@_L]X3D++gH5D4F86bN.0U:IK>7<V[QX]e&#JE+E@g/CA_R
C&72RY+CH_.2d@83<B,AK/6<I\B?VbDcg=U<e4-=+V8B^6f#/#Q2TSY8SOL@#LK2
5C</Z-R?[.<GI@22D6__W^FQffDKC/=QYA[./607MaJ2JX8UVF:FLW=-OH4:GBMI
YB6]@+_.bW-KJTEEHO12YOR]E3/@KITg>(3AEN]PVe?K5U=QW[,FFA4>F?R4RecN
Z_GIE9GU4I>/?-XAg=G[<M(>JXUd]YSOO(U3a?8Bd6cUFA\7e4TaP0[H)9#7T;WN
fI#[]cHYMBHQ<L1K+7?;Sc9B\EMS]D+S;^P(b.^YD^N:^Bc?Qe&75R;e^159+bKT
45V1:?H),YOI>KP<KeD=?ca?&31T&_(gUC[5QGeYW1?R;7c8W_f;ALe]JO.JbJag
#);@[^&L+XQg<JegH^G244S3,5>Ka0>fO(W.\)/]W:e&M@N:)^X.-)@JT7LK/QSZ
PT2DWeBB/,Y4_Zd:7/A:D=)PJH(?G[4B7J;+?YceKAF08U\J2L=[QeE(Tf_K>/.[
8..0Yf<72,.;@PZ/X&>;VCL39CV9,=]GY20N;/&dR))ANf5a-11N68ULEZD^SUU&
9K91a.2gRJY+7WN6=?P7A]N_Cb],_:V4Y)-BA1YLSeT\?FY;>bZMA(@,ED@T(QX=
YadO1N7gR4XI=S7@Y31)/NQ&aH&G_7_7KRLCVG39fR&BfM2>Y5W7;A)TJU\ME;R_
6Teg5#Ea-N#3G9N,\IJgd(;-_SLIOL@9fI(6RJM0,f7G<?Pf;#:^SeFVLf-Zf9?_
f2>I=Z\ge389O&H6bLNXb&]4J&>Y?)#(d^XRA,?J-X15Ag\8]SL800_KHYZ_JJ65
VTC@UPML?@EY/P:AY))UN]9U)?6#[:9JH.7cZO@fQ&;5(0c/C=JG<CJMWY@P4?90
O##aK5DT@>ZD7XZ#(c(Y5I]\eAR>[Q/cKZ@ON^4&dMJN[TcN365S(cM3.G1b?2UG
]1_>BTBgR6/d)I-.g3D(3D:<M(C4KZ[LMD7gH7/gK&7bFSWMW4@E&TU8Ie5PdG#Q
]BZ/^Z#dEW34/EdHJ&HUdX7A-eJK>7F;3A-MC)7aA:8E1(Y[&_6S>83AG<+SS7E>
8/M:0f3F=cVRa;<dVZb4):N@&[A77dO9V\=_+>MKF0ED@a<f:@WEfR_6I=+(g9b@
F3:YM[_5[7L3+g]<VRU?f#[P>78<E#]<CO/0=ZOB\F&6.dIN:QW[#eSWL/A/XPF(
cVT:F61:12cLFfQ>T\_7d,J<RaeAcL1C1Rc=W2C;0c9-J^f58CIPG7<XcK:8><Q8
ab#.+3aO]ded\AfDUC-O>2GaW=6UQ]70C_X3Y3_9UTQNL]/FZ(a3LG#<N\[[HL?I
7YU5UUX20H.VG9PXJ_TNLdW&J<I\8cPBXc[MXCKgZd5>8c4GEZ3)E1IJC2KCC]=(
C=&;c&H9b5/>a#f;g68aTcB:LO]Va,/,U+Z/M0#<R19LB&J(6@LYf2[--GC2PQaT
.I?d9SLaI4PT2;cZf,7_@:1TdW=2<[1,_S=GS+ed0G#OQ:P)<]RgY8\-SCUSce4L
U3]3dZ1#eMGQ2:3ebN/Ye&,J=]a,LD?6/Ob8>b3)a+g]^_G_U#]OS2;a9Z;>4#;[
WZ@6R)[D):KJAO51Z6YF>=P<,80>4G_,-Wf6Mb/<4TZ[SWASX^<?1NMO#Q8T@GBB
PCIEg<OJ#K<fYLO@(5T&6-V7[WLGFcH84G3DdZ?7g;5C/M]U=CQ^;H\6X3ZN;6C0
2SMgJ^5&f&Z5L,EY7\IGV8g_e:48@46?JaY>[HMAggN.4X-T?(JJ@I;K=Wc]M+HG
ES?X2>:7VZW]gB92;^65JYSM,)71H6+7GJMN3B\>+3@4H<f^-^TWLH-.f-Y_:RQ0
;c.N<MB\60/+@\7D>V_N;QHC84\5BRUWJE4g,=1]E.?Y-)LOcH]MT+#H0U+S@cg@
CQSJH2;)K^J(d,WaY9Pd,[Y@A?XC<V?SS<W@^80E^GIaJNFL?&)JBaO^98#J9Q>F
,bQDZ<8C2G4IfS=@5<Z\U6SCPc2)?J>XDG:SXe>1#K[b=BCN9+4PNM4dER)TH;1E
YN]\M[,2b@\BNA\)Ma#HRAcM9?Q[SVX]D@YD)>R,=>\31RK,M;Ug8?;P_#0&g:6B
K&^)[70-,OL;#&.b01(#)QLFc-L@0ON9R9JWUBCC-ORO@-E:/-c0/bU27YJMDd8Y
FeT>#T7KcFR\b.cRY1c]EU;;H=92+V&e,U4O:0e<()Y;gIS;)c^C^Zd3AeLX]9@\
;e;&Rc2Ee7Me,4[W@GJ2#e1ZE[QfJ:C2T/P=^fV@J=.f3IV7CLcT\FLX##@S_f#E
M\-1W^UPIBIV#S/C+55@,8;adU^DD,BC]#=&0EDY10eSO9?<]R\>O>R11e&8P@g+
_N@_W6W,LU^E(G=0(f@Y::bXNM6QZ8,/UdBaUA,C52LYO6&_6+9d_<@)<PE0?)<H
-4F)K1R4S^SaRgQV\\a]E7V0g2##=2,_08+H]YL[F[5fTE<K)IQ(0LPEI[CZX33]
410Y]Y>W,;Q3:d/6M/gee^[H)+JF52a5956,c/&[eA:\IBS8b(dc[Pd39fQB-DQS
WNKORCJ,OK+VF;g?P?U@G/G+E.dNdOI+LGS(gX-1]_-(BcV15^.+I9b_/.OX-:1)
=&LF.e3;O,6(APg86:[^a9cE]49\e\B3@bRGgB-:UG.16_^TW+X2P7f:W<0Q]D9^
7XJJe8R9LCGS2S8GS56IUea1[LGU^N&YRJ?MKJOfaN:5;2VXX^QeJ>AD[@fSgS71
0XCV/FP=L;THV)1L(E=XFY?T>),Pa,\?B:^?B3L3f_<99:=NOR1(&98eULMZ\g]f
[dP9de#11G]R[=C\S><0@=-eKAMIUM6.G@OD4QV-9g3S3AL-PO?JbE82]&(SPWVb
Ic?(gf<Ld;4]@C[(FMZ]b(WEb/geVK#G@&0g#;JLEA7Q5<a9]6--3?J[TbBU>1b(
E0ZKAY;OGgSBTKJcYHM[G)9CHRM4gcG@(N&#?CARb]NB7)UZBfD6.cK?@1_<:H@1
XbeZ(_e2GP^VUZ3L6S&L>W(+NS,S,E6(Jf-R5a#^5AMMV6g3.D_1F_4_b5a[Nfe0
Y=HdU8fC6W<[3]0,JQZR#g)J[WfWH2f_[77F08E@7[O&?[b:cFBOKcQ)L]B]+S5S
5c2EbVT8J@]0DSGF4d31F)GQ:.2JL>/X9b[9<#4S/;G2RbW6e;/X>&\#FY/405\Q
-/Y;.&KZO+H1WD6b/)JM1GTeI68gGNO<G.:[S2)]SM40eUJVWPC+ZMX(GT7:cK5a
,0:bI8.2g3]?KdW=;+Tgg.M.<TeJIZM95DPHYM+3/?4<5ZMGU+/fEeU;<PU?)H+6
UNE+8Ka3=7^;4-(_RK>W^gJ^VW0/A/=>=@c@b;V6U76N1HKeFb=1IP>F8LVU)X=W
Y_.#6V+^YfL(X7).CD/H:;(:f=V5K:e6K;1;D5c,)BB>54g2WH(B\M02=7WW5a7Y
6TQIKSK]8aA1AedZ)@^;5RX=PSK)&7+##;0_B7d:#0D.89@,VYf;>-5HBOE^);)L
0Yg\1Z6(QEK5^J,F0\2M]7NW^SKdR;Z=A4Q<0De<K.AJ;W\9@QJ1dD,7^>MY4&@E
7.ed+K;,_3^:>)BgFZ<UOZb0)J.DG0_4d9/D(<CLFON<N@&_Y]=bFGa:=W?7=JQS
c>fU@;181MdBeEE5-Z3MKd(;?B,,DJWS#b_E>QcbGI/T1R_L0dIVg2>G?0F&SPgX
6)U],QI:]2+;_S1,Q+eB8&KQ_>Z<8>]J?4X3aYSB&c_Sa]\DF/-3=&e9JXMDJODB
;DDUDCW?[4#G;LY;9DgN,^0d.3I.<9^;XLaC8)a5c)d7W>b<WLSE@OD2aEGBbQJ@
5D9Og)193SHd>;<4@<>HYg\/BFOQ^DKFX=V&dI<7I[8)2e>G59,.[TO+R\3/8/WP
[#IB?&M(]I]KMfVZ/LY9+-K0MENOW25PT]a7.NO&OdDN\4e-&Q0MXW#K^Gbc&:<+
+S7+a\G4^7bYJY;D4+g#4^-,LSgCf]S\Q4;\(aK)Kf#XJ-a)d]1(FBJIaRXJ#Z7C
;bFbPCa4D#RLW8:Y_WbdZ6[?+R+a2-.g[c]PaW]K1)\F\],9<,Je^=@_]2A9?7(F
,b;de+[NAWY\B/,LD@JNSF6fc_YO-0DGO3.LQ.&MY5aPH50XL8ZW6X?VH[+-8?e-
0,_V]E@D\G-1CO)^B1GC33,K[_MJgCEF\?W;AU@IN@&T=YR9?1.O+U+@:HVD0Q[H
eTN0N1SI2XB,fX[P2]5e-2THcS4I?Z)[Lb^T\PaE9?8YQ7(.AbV(+&gT>Q&fgST3
.dCXJV0F+.JMB?X&89P<OVcKaWeg\9]XbGUNRW#@#8Ug:.#-9L[,&N1bCdb/+THb
\),;R#XV6fX37IbeO[4]N-86Y>&3,X;0F)[fT&T4:+FAO31F/ccJRWAE7#S;?-/@
Bc:[GA/DLJH0X1D=&@6O@^IdM=<//@:\+LH4gg@\NdUT@2aL2F_Rg7V22ff7e#H@
;f)0d=YZ7HR:bV)+^F.^S2\\ZcZb+3\MB>K?L-UXaOd:C_g05XfX+#M:D1(1)\.3
P.RW?HD+VfDY.PcV1E=ODK6QF-VBS\-Pb,DJ-^6T8/Ea<A4^.>>-W^#C2AJ&W##V
b0=>-cLJQ6VWDBE)c3Vga6SZJ3)55\0<UgXVYa)G>+e>F89]7ZP\V)R-dPX^E0QI
NdHXXIZV-[\G4C/<;eX:[0I&9P0[+>?+XU:D:S1RUeaYKJ\J<f/a_HBedMMCVC2C
6I)1,fYV<(<ZF.2:6FD@76:/^^9=\5NMVH><8R^@;b(fIc3XQ\@WB^6UR=LAPcdb
fa3K69AQH5YFdWDL13W2aT3\7)dT#/E7fBXUO8>)d31YM0b8_-gaX^g&^@>T,3R^
7SBV]K(I7:9/e=-VX1#06e_GC>fJT)^42CZ5V:=P]1VGGLd-X68JS[.6X>X-J7GA
A5JXTXWZ1TVY[Y,dP5<+B9VZ<,^GVSXf_83BE#Y:F6#G12DcG=g&dT,0(BSMK:[D
f?[&/,=b(fC18AR6Z94KM>b>H0Cbc:&SV/:fSPA?1U(ECFY;BXcC>HK0[;)H4GN?
HR&gXHdDJ?HO\CU73,gGMd=8=;.;9bK-:_T:,Oa9b0O,T;DGScOa6[DAA^EA;WQS
B5Eb4@(1SNI64]<-B@BSIe2\=)^fXJ)aKZV-1_--?f>;.P;ad.Qb2^-W6>&=[;TT
L2LI/-NEe0<FJE;C\:c0^AEVf@@X_&e5OLP[^(e.OT^VN)KQPd7^d<?P2:gS)6EX
G97B\97OJUL[#W:FMM6;f:(U]WQRT_@fS5Z\&/MC,#.Tcg2@CEQ-SIdMJDgOJg]^
74)gD:&8(Y?AY;g@>cOMB-;cd1[a2PBUQ+bZ\(.ag]bE5fbCRY7O#_;1@1#6?#U<
PEXME6B]>1W0Le?fQ-gW-[LZFeDYGB7>FX7F51TF@E]UK.aC(MbTd5NEfOJa:?PO
_TU,PGQ]0Pc_M]&FUK:\Z97\7H@b+b#_\6KSA\a1bO>#G#&KcE1;D.SLZH:NH1GJ
>6DGeCJ@7d9&=\CP1^6DQ.gD0_\EMf^g:@f2;PZVW^.D,f9;;Tg_F8bAQ;-SHaBF
Y8_+FgI^20XA2S=5N,,@0LZ?O16Bcb<[fBJ&W+6.8]Q]_fdX8QHFe^BBOR<MIN00
LPP]1=D;+)XJa<,_S/.cS&(LCR+X1DaZJG:2bBc6dOf?<ZPgL,A7NKcA4Y5_00IA
bMeO3Hf,-5ag2aBb55E4RIEJP9._=2L\(XI/6Wa@@4C@a>TVQMe]TDDeNUCC73d4
0-SR,PJ1NCW3d],BD0=MI0W0[0B]PVd3gNNN(Y#1#W<4VP-B+K=OXZ,J9LDCR<?)
;4Z/2<:,BKd^d/a,b\^QA[^&X<PDN)bYSbD0JS=+19EKa=c3PN>R;+CC]5_D1c(\
3>JSKEMRY@(c8bfYR8LY/K^QZCA4[/34_;:E/6YO+>AGVf=[b93XOR-LV+>?E-_X
:/S9IDfF,_]+9ZU2DdF\aRESF9ZDY<F41?,MNI@Q=5(2S;9^Y+RHa&:R0eIf((_D
++)>RCJaA0-1T3,+c-T+;[E#IB8WYb7ZZ#&):2<2aK?]FR/[Wbcbf0.R2Q(aTdfX
d02[[;5GZYFO_31?OT3@K<bg:ARFU22O\C7]0BIB]=_ZOQ0cN:PE,<Wbe.?YJ?,1
C[fEE/WKb/]aK^KL09L:)e+Ke/3;B-I,]9MNf_8R)<X#BfP>VC=?Gd3cO9+5+Df>
WD/]G#@fEG9(K0g2X4,7.U:]bS<R>@&Kg11->S1NZWR2K3D0gT<(Fd5^/@VL1eIe
9X_+[LB:c&Ke=U4UHEB#K46EVf.e039gMgE]W;7b[/.,.&CL5)(UNc[W_f:GO8:.
Ic5c=#=bde2?EWTCW[<,?=GIKU6.,dD#2)U660XaN63ACT[d:I:Q\P9;bd?)gMWg
FXOTUb:B[J2cI?<TVQKcDTOA_=@Q0>egS8O=-IXX4A:7T\)#1S1acNF[6)?[KLf5
P@N7B\5Wc5CHfJ=+0D90dHV\0;XBZ3Ma+([QaL\Gd54cNFEgJ\.6fO@N:.a7B_#2
ae.954EU7M40S9BEG5B+4N-#YHg5bSB6MEe(TH77@0\FHG[Y(7B\SYJ5GdQbG/>0
IVEJ.>4Bc)gYZ4\b5IY9YWWQZB7O9HS]?E\T4f7HQG4,(8#+D=/UY1;K\))@P1.-
Q2^0=eERI?(ET72?]4Ob^K@?MHEMJCUWH)TMZLX29B7@?L1&J[+;X;/I,,08+P(V
)0)\MbGQ9]PBJV=]cL@[Y2N:B6DDD>Tf#VGe\^TW4R6f)#0]bM8\P&^W7dgZ:.]6
5D]#O&B3+OT[K7+\<S/T8bK]1V7cRg-OCdUSCD(8d=#OD50-QH.C?(83XEWV/P?+
J?5__]9;IPd;)@\+(>W\J.;;fd8A8g,0_9X&WA5K\Ze-bZZ?(4G(g[5Ze),,VHNb
G#C(W.?C)5cL8;D2/^VAFE1DG-Bg6b]_,dOaR,.RQ=YJ54e,5]2Z8U4f/;M3A9,[
f]=AOLI1--Q(N4<GfgYdX39.=UbW=5TTdIgZN&W2<9+Pd<P1=V5dA(NVKN)FZdJ,
=E[X:NZd-&P>NF)=5H0)_6GcZEC-F/-H/8X8DE2KM5>7Q.#Q\B),d\e&>->Ba-,/
64IGb>eK.9ONYOV=9[G^J>F:4aNbE^89+ND_GNY<9g&Jc&0CdISB]]:7=2[4RG+,
8H#RcIK2^1P.KG>R/b0O;+42NcdHd>dICF\#C(4^;N(.Bg7]-FAbW;\.bA2cbDaK
f_TD;E>>:Y>Ae-f)9GDP4.>QR2GKEgU;d.S4,A-CDLgK_R:)c[B,^.B)HaLC7gO.
fBK(U8EdD+K?;@W&2(PI#K:,YR[&IB5F?=BO>93UC/ATH->/+>E/FM1bFU[9=K:A
70#\BBK((C5KQYB6g5_2YJTceIKK=d]4R</c:8-/G6aZ_->Wb5edD4BAd;J:QR/F
>f5L8<=4c4S:)(P)U9:#[1fP.Y_:IM?]1T<@/d2POMDWgVcUS^PPH@(b&0&b]BaD
H_KE/PN_5eeM\bERIZANY4<4R]8]2ffaUAYIAZ3a^C0FXYU/\GJKAJL?&?eEK_Z^
UTS5c52)&NS7bX]A+^WNbPOA[Ya5J[55[?[T1[VfNTC/X+VUV1-T<c7N]bMF]UM,
QX\?Nb=#E3IAb.1D,6c-cV2]9[43.0F4E;=\/9#6-EcBf8,/0/NZW;W9fB>DTK51
O<1Z_(ICMQYH6fQ[G3ag<>C]VP@#AB&X+d_T0X,2\IePfM5@g[#--/H(Zd;aS&>^
dMHIXZKR#>L36>7+:g@/Jd<U9>K[AM]Q3>eZ+X?A7<e:Z+<N5P.e?#\[)PAX1AYZ
\IFFHWe;e+0>TdbBWKgYNZY7bJAU\#>>aFNFX\D()S[&K(31J=f0Kc8+;fSE?9RY
F_3LV;G>3)B:/EU@8E)&b5C\^Vf9PK(/[FXSDKg4A@X\?;aNB2T2#0@=O.SZO48b
,-Na/S-:7OVOY@K=,-9CQfHLfQ.?Tba(I_P<?4,,&8DC+;.]1U=:4BZSDDL8&UD8
S.F@Z73^_#B-R)DSFg4&e(/X1eJGfAXcJ=,0R]:Q9c^fV?6+HdB;0AaB0/c.==e)
EQ06T.W[0>P493->X\NDU9J_-^9\GR:2BbU[/Y#SNF4:<MI7a;:@NCCD.JO7Kf/9
-Y>@9_:[N4WXPFDN+J<eMM4H9W&6[fRXJ13W&?.F6+RV]/&aD@VD<;=XB(U2eV.S
:BPb;fE/Eec66RT@O\4X.;3\4V;DgMP3(e:L6W.(<>]W#Q=QbU:TIV\8CZH]BY4b
T-f87ba??YB+0+2Q<FSf[^91;&+KQEY]HS<1HE+B;8TN=528503XN4?5B+-f]?YV
LV7RB845<&DWI?_@Te27=_.KBKa9.O2a6I71&51@W5O[2W4ebTgLK7H@.E2S&.Q4
f7eNKOMUgY1)B5/IQ[BPE3#_6d@S30+2fCdOK&9fPb2A9<<NTO?_9O22O3Z^UM\U
>W(gVACCW52_[CT2X7@RUBaPY_-HMI)9L[#e(&J>V,]DWdQ@5Y@_Me1/D[GEA(A>
9WGOI@HA=N1(\3#0W?5/bZ.g2S<VN#7DO+,e6[(H+1\d@gd8QXPNQ]OF=)(:Q)M&
6D,P,NJSf>R(^d98&QB/0LL@KG6HOOH1H;39-#DN@;:&8^O4>LH,-BRYRE@3,MD]
7VK0BXaQF^+c<C\?;U\G0Pb_+3dZBgBYS4))Sc-BT6e@KNZNM0II0]JU^3L+_PZX
4PM;deN=f:bVWUAgQ]X)XC63#7N<&;+fReM[a/\:M9E/+7KCMG\e.T8W->,&G?/0
WE,,PQEa;O=U[gNFE7fI_HPM#PR-0T[9NGbaeXO#cgU<fS0#1DR1]UD^H5gR;N1Y
_Tae7,fAdL+VF<NXA4^d:b]OW@;McZLC&<),Z9U_P6(#(^b-,5TeW9<2D,fFR01G
M]HOg8480,@8:f4#3/30a<dW(HMAIX_2D_FbM#e1_bC0A+?-5aH1Ag0=>L-1eYNW
NO^ERNJSV#A[2XWaL<&Q^?R/5LLW261Z&O]UVAOf;63EC,ONSY)IJ#R:&)BWb3I\
D[1KSZ/aAL#,XOOM,I4DB;O+(5\)a+/QgF(-4^4Oa@/BMBF=.-Xd8L2F3G.0DbK,
KFcP6;W8\8fDV,R^&-<8_:4YYKZ:T<Y38CeYd5<DU-g[]?11)X;L+(C/90Y&K7Eg
5)]HT&&=26\L@D#PTGNd\eP/ZSL9bHR<FMaK.,[XM&D0f,57#2^KPD;H?NHdbUHe
-1>C80>f-4=8K(,?A2]HbC0cUXZO@B]178EGbQA4DG[ZUC@C7[g1G<^61:,R8.//
&3-^b2(gK=3W/NZRS4&81,22N]-VfDUDG@\-4b=FL@8)5D?(VYJUTPYG&J\#e2H)
bGLF_,,-I[^>eQ_gW8If7VAAUP_KRY3GF<=\Db0/>?AMBdG&g)0dMdYZ:_E,\>O0
G4e\e<<,]QX6ZW,PK+^,>1F-^\QKe#4fgcb9;5H=(LZ/E-LJR.,O;_TYb#?0LI;F
:[/gH.0#H93;aR=T2I8H_L5f@eV:Ebd0C9cX75Xb:SX,Kd0X/S_+,C2JA<1?5<aF
b.=9?0>NfRD_K7P7GOI;?6EE&#=;1<-FYHMcL=Fd+/a3053bICA6c8?O1L#->6V#
geZ:5WV3a0GFG[IY&@<;W2E\Z#8WQACF3&M>MZ,IJIF[HRY.-XF#R8^<:GM1N^0X
TBXg(G999<Qb5^a^0WVO(POKW5AC2(0T9):.P:>-0C5D;/_EM@g7TfK0GPIS2NB\
5_#]X>&=V,D8LRW@DKS2#H6WNbX2(VKa/:J_ZOBXVAW[,LVDUbRg&XT&I0TFEQKM
cHH#.MQ2B,,#\)&]M6YAVXGSdEL#I@^(;NRE:/=DZC/L5H^^FOTM:0B/()a[Lg<<
6#^03XgL:8Z(SSDM4D+c\gCTM:+H\\94_>,YB1]\#08f@@G7BQ>#[6U;A[23YOW[
>eZ@_L:BXE8M,@)5V]cNR);#[f1BW(A[34?=H6]9Y@Q#5>;N7E.4P3Y?ENdA2fVG
JL&I+\W>LT>OT1[^#P8aDJT?UQ6bdK-/ec5V[FDD&MWV#MQ&T#UY?)#(6SI:)e:g
#E#=2\01AG4R-]ZY>.#IcJaH8KfZM98EA(YEbcaeCfQ-4F1<)ae:H/UU:]d5F#UT
4A<d_EC:9IY(]FEU],&<XCa[/:KgZ+a3fGM93H>DR&:Z^)&-VgcR91P]@T7B9B@a
^AV:-^7N3(PZSdP[R;?cM9-]a:68;NMA(^YUQ?9\YQDVGY^3DV\[Ga14X0(geP\b
DO6K6g?=6+ARfJ&=#[(.aQ6AUY(@4LD2##(7gFH@LGR:2<b7KE_<ZU,bN?42EV\C
\H.Ld[O7C[:_.HI-PSJ\).E8Qf#<[(9^<&U0U/RSJUD#c(,c=c)M#=GbdLF20MH2
N8AAYXPT-EC_C_N,ITBK+<0^.EZ)(g/aQC2X07Db(JO-@OB#6O97V-&-Xb[9[Q@R
4(b>A5W&/I_H8@/;b:FQ(OQa1#J,M,5\-6=[8a324Vb?#NJRE:FRDAN1D3I0?)Q5
H/TE:e?UA_X(4Q;2.gRH][R#1ABHMC9c:aQHQ_(5/(;@6[7[:R<bZ+50VB)H,)Og
(>P\;,.Ied0Wf7)T)dA&B/EX=9[7g(_DM=cIc6U>LdJ;X9BW04,NFEQc8W;Rg28O
J+:;J(NY\a@^T[1OUUT1+]Z#3RJ@<8SbGHAX@)KeQeR#,,cWD9f[@_g48UC0VDWK
4O-e<V+FTcRF]Z\Q[Mc]MW7G-fMZE552<cR(;TGP7Ma_G5)QdbeBWVF75cM]9O)0
8XX\Ba\<1X]eb83?Q&.b.I3P1H/:W8J^0.KPPcHdJ=<[UHN^Y+:cd#TNdT?I3NA[
.a.:[5-=AJ\;6[eddZ\]8>2#-B)]3U2@N3Te9+D>G.f:#(.0=_50<dHP+H_G[,^E
/7?NYN1dfQFJ83>e&-=9[J&bB/_NdY(bGQ5&<^9I+&b\DXK?BUBX)4a]&OL(7cT]
U^WDWPWO[13&ONg)5<-O?X_L0/(BSXd/CG)W@<E<&)2/-ODIS]7M:EYDQ6SN2@Q1
d9@GZQd#+C8Y1W0IF4K+e6P-LHRd8e9+dN5Y_78=UI)cA,,_6ME(V5?eO>B0abM8
dcGDgC[JC4Obf8WX\U^EG[P6I4FEF7b@>g&Y^92C9:6DH.[I5,:fF9G)V];KCB;K
_I2ET[a8\X#@5ggL..5BV\Y.=Y[WTeg,2:T#M=M=9fB?\)I\R5I7@/6<GE,J<.E1
8LdBe45WV<35FgM@5Be\U,PPcf98/36=S3Ub]?A64&U+c0g/HZOJ<MQa25SB0,dR
8^dEQ4]1/D>FX](L,&YQK\/Y-0V?E=H?4G3Z:O)@T.WG=2]:dHPM=]fUe6a+<Vfc
SCYVH7Z53+E:RJW_SbI=OeH0b<O1U75AF4/aBZDNaOeP]@2Y_>6JbC6/C4-;d9B<
@Q+Na=M/REed3ED4Q?]QOI_eRCH4Eg]+JOCdP5d(SGO(P&W(N-G&bcZZWPBJI=2Q
SCW3LYfT;F5Z&EM2>A.8.WbJTB09[9N9\#3NH61?g<#:cRNDYMBbbSPW0=D[Z)OO
>7PLF3XPE46C[(WPK\(H2-@bC#4f&BEK6R)f-720]Xb_I^5=CVMB=AP-fG;[-Vd3
HcH?24E=6^dT3J\5U_Y(+3O2(3(CaObA78#3FA71Ve]Ke6GLE9(T(\N,6b1.B&))
f#\QUXMI>Sg>Gc350WPQY:=^@LTb^[dFKF:4Q_(#H([e--&,g+bV_0;BY9CdYD43
Y<0JDPg.P?^:1cHD&FbNT/T1b^]\43P/(Y=K)W>E[OaBf#\+bS+[D.E=&e+D<.1,
/OfN,7KH+<:<FSK)S.MV[2;6)QeXbQZW:A4Ia/L>QQ001ZIc<b[5R,;L#?@+N#.,
\@U@@WaC3S5\J?cT<//Y3HPc>OROeB)-5g88=9=2W1>YYM?+f75NE^bRe=?1;):(
K]XIDUK.gJeF3Lb#//5&WYb<.CY#_Vg^G::P28Nb106T)0c\8,CNJF-3QFEf#2Db
BdcYdN@6;PQ0YbZcJKBSA:O(WcPZR5CD=g4LE0L+b3Y^Q-_X<I<RKGe@Aa,O=aKf
^BADEgc<JU7S_O6.CL2TOFKUPQ6aX?0>Oa3Q3_aHAOXT5^DHRHAJ&?H18I-Of6KF
NQYWS<UYN9,U;fb[c_V7RQ^B92J4X1RV4HRVBPG5gg?M>?eK(_VUCBfKd.54U>+&
5E-&X^(+?#036HNREPOBOH_LS=-3M8DAG6.8Uc];)=e8#g.f/](4P2Q6&M(1:gCP
P#PI9G-aD+M>K6E,GRI0M^.H5fR;P_MC/T+\1b05b4KVYK-(2I1,IG4H/(E\I]g6
8JKc,T@37ebT+P]e3.PD><&2>-bTIE6K5IgP^d78=#3Cd8NeRQ-QRVM<^I1@IE]>
>.,Rg\NH&^Z/2+#E?SI?g:\;fM2a_+Q9.N:M8]ECb-1C(7&7d8eI[gX4_8/S10M;
B73D;;:OK&.H8T8e5G6.((G[K?L@Z13bTZ^@e5a0;HBM[DWaRVDf0+(4F6GTS?\[
Y#GNLHA,b2@bGWYU+P_aG=]4T<A@Y#8)-,aPX2E8CggXY2K1QCO&1J83-?LOU0K,
0+IG>-FMd<(F8^:[IWQ)25[,LDeF;1NIdM7Ue?218RcLJ#3gEG..6S;BJ[MBKXQY
Q\bUd9DcJP5WW0G1]Eeg)JD:<1X>/)-O-VAE;>/d5eW1O\SE^HS(.dc8AVb_UgPZ
&?gW2XXPGe8H&6S#VEP.3DKT_=</YaGZ6[L@Y.fN;aSWD\d\]-DL(8[;-8Za/)c+
],aCOR-beA>;,RX2cRP:Y)&FPd\WPFMCN/^f3<T])FL&2:D<4]ER6f-U;;#ZO=1U
LaB4a4M;aF)SH/0+(<1N#Oa#Tc+PR75+,MCXVTJ(NbXeVe(RW<ZJQ2BU<7GO,6T^
)0.S9@fIA/KGCeGTY_V,DL6V&FNUJ:H,VgY]XN533gC:[>\#\cR/ZSO?18bde_@e
/2ecQ[]@Y03F//<,8\Y0Z#E85()XQQR2_+g8@C<+1#f0EZ=]#,BT51Hf2)FK.R-8
E8\A];=M2-W.[NP)>,7UWQM;3ZFHOW9,gHEQK?I7Q8c5W#4[R&L<\a]A3<_UM#Y9
-1_4e)-a6Ce3g:2YFWBQ/H+QZe:FWM#.g1I+MUY5XV]6:UUIE]N?I>/2HY\RTHbe
deMRCVF1A),1KU=\UD\2cGLK#gF=_E>X+UN>V,e7TaO6KdR0F=^8QF]7A;8)Cf5f
5b+WRJC/RS1LH\aU:FVL)(8GMabM[][eWLWFOf4^7YS^V?B2EH=;HBXg08OE8[aQ
1UZZQg?0eMBeB=[f.gX);D)?+/S^UEI@Z5Z=ZBY_K8K[DASVZCH;SVL:8-fM=8dF
#PaIF?P?]QZ^OS4Fc6fOL&YV@U/4DS8gBc0Y/QEO=/cP@e\,g#+2-09?MO>PR8.^
I9:-VaL_O^c[4<6_D28YF_J/UFT>I@]\ZFQ:#9gf9PM&KU:KLV[RZJ=.//0SOK\C
5O23^)dASQC;KdDZTA,/=71TaPM83(=VZ>3>RU<D+?2DVfYB\BT6U;R5C7Y6QY-I
a-M0GELOY/)aY+g/N&Q:]6FX0PLVX[F(+C8>X4@[\>bEgI?@dQ9[eYcX_S0DQZ,W
EO);B<cWMQ_+;b@(b&De2H22E)&bC^N@7INY_,aTU^HC,/Qc0ES9P\>EF:K57FJB
dK\P5F<N2#^:6Z5.T_Q+(OA:gG^AQ8M+d57H0Y9(:Yc\c)\9A-a[&@+ZQ8[#8#dg
e91,@=AHGW[2U6AaIc+2V>dFc@-SHZcG4-EH/#54R?=)ILBd0DSd&B.f,0,^J6f0
e33Q(<fgCTd/KQc<<5#G6Tef.N=]+eaIV>YQ)XCfYYE#]GR,.\C=];N@]fJZRSRI
4GQ/K::e,=?B)PV]BD/\)@2BIa5CX(R4WeE+=eZU]+M&]>NXa5NCMQ2X:N:AKDAF
]^)JMMc)\_2DF\ZYf:FQ[D+_4FaW//FFc]dZK0b.9C5>ZO+PbHI[#B_@4A)Q3/fE
^G?f4POabX>TK5[?&4F75#(b1,g,b?#R>\7PbX<c5cbJX=a=Q2]481NgHQ(^+<-Q
L6H\/R[>gX5+LVY-2#3M&.F0T-(5.+W>NX;D:+).,XE&#g@1QYQ-E08P1@/D[Y[O
WU<#=+-BF/\L3JCW(23Ee5VPY2F)=;;_DZYRY/2RQ^BV,4>?fW+-e=)/(TccU_KX
0RgIe,D\37K<PIC-bH9-c:V&7^Q&Z[c^1DH-Z)O7)9Q(WOM[\NETV?A@03/7K4YL
XP8V,3I(H@:MEb9I574-3T)N>>_MSOKX[P/V>Yb]KBXPF1?:0LC(+=<<F-UEQAN9
Y56&_/&3a.?<C\g2KBS>+af?V7+H6>Y&5@6ZUb[,@W[I1B#>KI8Xb4APQT8H]B8]
22(M\XNRf)-7(Z)I6g@W:FR-a<#@A]G1gLKUA_e\<][5E&AcYeeRQU9W)(+\c^d/
\YZT(QE&(SJAb44dV0975<:Q;#+?N0)K8F#N=I,)g#NEFNJB?,dA5bS>->.=?Y0d
?CC5b(JDP+--QO;]ZX5RaCAgF-HP8U7>:gf4?aOT45E+[#Zgf(ZY2&AGCbgG(JWf
I8<,Y;R5L(TDN/47>:>6I8GYYCNVVVb,c84/X9T/#:/=W4;.K=8#&3WdOK_)E/&H
(?^-cRV;H&;1TR[GcFK__5fG][\R,E/W)Qdb/599>42LUK5U/#\[[,d,/^H+\OIQ
&\1YT70QK=/J:+UKRZ8],c0QcK^7S+\NP<#7/cY^:O/+CL?Zd@G)RG/Z=/TFId[C
K9=UC#(cAVR&62[Pc@(<d76/##CH&#&R8HS<[0d0GFW9c9ZSd.EW>KBSV/\8R\,\
A6#IN3fc]5eIU[6dF6VWMBW=^GGUN<@)AF_c-#-BH:a.IE155=V;?21LP7c^S.PK
Q-eGGe&O8@3=H#eCQ-R\LHS_>DOM4(8EH/3B:4MK&6&(#P9,7MB\1P]4[;,V(P7T
J=KWaP^DXNJVJW:N.UcDVLB^>3EU][RBBQXYZI4B6D9XLBR4=[3eR86BUb\X9e^6
R0H<YSEGZ7CE@TH)\>R&Ae\?2J3f^W]#(Fe9:@INJ[)6eG=04]IEaG,McdaYcP2F
:19Dg)YV[I/@1P@AUC_P8=@3;[6K=\X/R@-R79C9PeS?\g?^V0_UF^[9)a^?+4+I
f.f/46VMKeSZ9EK&JUaT6YB6&9KDH;1:R]>//d#IEg)XVE>AbN8F49&=g9VJFbL#
7T,dZ1Z(68-0;31/;24JH-7MVG90-eS:dQJ9Bd/g-JD@7ZHZPT?c_L31N?#M]63>
[g^c:,<P<d0?5\J>7FALe1-e?U[3>1K?8^)P=Fc+XRad<M6G-KQ0Qb25UdN(R4O6
E2d7L&eHfILVV<_5:cHD.>^;AfC^SPa>AfN&XUC=-RQ\9&P8I??,bGE3[\5g/X,L
eZ)>#O=527]-3BVd4_LF+c[HIVV>gTJ<SJf>dDb#M:]UFOW17#Y&U)B/b-K0;R6N
LQQ1<VEgeIE-Z=&=(XIS5209L#gLOP/LaEP@QE4CF@2G0Q)L=(63:WY3-IKeT2YZ
/-/=PNUGQ[WJ-FC^Y+@Mf>D;_K#O@=A>N-K+G]<aKI5012d0TV#<T1\g3];)f=NL
D;,dGaK#5T_b7Ec&?5D//ea1c@N6T)a/e/U1:S=+;/c_\V,WAcdVFLWB)N=[Xb3\
Af6J,2&.];^3_]KSB+5S5HD62a:<1A7;5RJMQ_OgJOY.+B<[#>TcN.<7QKV_@U&7
PH86&&U-T<[R:3;,;FIfd_6_QP.\?K2HQ5>702JW?KF,NEbNMK^X+WJH;92MB8S8
.#TA)?4/8Z22c<=BaW<QOWX4_6N.ES;PZG/GQ2SM0YHW_g<e3Ba_G=OHQE<]Ob@=
UIA@2#(QDY1c:[EQBcIgeFLfQ((c7D8&#4^#8De3U.\1>c54#EYbNFGA7a>/Z[-N
Sa,VfE^V/>^&UJ;)B9NY^4?b>4SQ1:4>ZX]HAgR<I[D1J?UG6@g-98^2UOgC@QVA
>,d]WD>8F?,1.cUZ539)LS,XLU6)&g-<eXU7M9?g(?G)T=C>7c#,8)M\][D##f0B
WYW>G3EQ:FNeD&BC=2/;d&X>;BS+>Ua@?Ja=VG_]V]b(AA25Qe&6YfX\eY[LD(>(
0MSB-[?4Y)P4LSMT0(E[)(KcD02^PYA8?4/19&I35JW2G>Md;PQ?e,,9._RZ+HXg
LPe^\^eUK@-A5N1bMAC\YaTGc52+Y_\IZDdb7-9)9PS^^V:F1@b]&Z&-^/VcF#fC
&a_8&UQ2f?CAd#)3@VJNK9+MD6:256[KE,GCG_J+FVGZX1ZEFE0?BC787NId0?ID
FPeEH]E<]A\CW#RQ@3/)1([1bO<-QTe[[4c>V.I;3e+&&J(geWESJ5];OZ3=WD,C
]eGKDS:_CH],e<BALd4SbV#M8<Rbf&aY6Ec,=)BFF&cJ#X&_YV8N@IIQG0+Ka0MH
.fV^KYUM1KKGW>S:#,-:2]c@]#[dJP?Je]A.Q.Ye1FYX8J3eI?/Y]=F)8[YJbEV&
M,;gC09W?.?7R<M&Zba\/6\&;R<@d+9I8_[X<a9)QR^EMFHQ1..d.KXTS#I_<,PA
?51cVN->(6<75=Q6]QJ;D\LZ2>c+,>-RN.-aT7]U3deR;UMW_>LUd?3A7X.DRLXO
>.VRG0.=SU&58_dWAaGYW4G3&Wg=.)Pf;H[(T+6dP_L)e&+.aQ;^[/>\ST0W7,C-
=8TKRLVNMGG0?S)NO7W3Z^[YdAJFL;Jd5)8U;?c^WECXK9C_dT+J05DTJ_La=gB@
cE_=ATPaX&91HR^LO&W.K74^T>0PCfMY@25HAWM>9K4bT]EKH\&IMDRa9-C(A0IN
K@A)S3<7WgDJ<&[0(=205WNg]<e/=,1\U=XETT^1<Z1.Gag6?3]F+1N5XH.AQ+7.
FH/0d_GA+/C=\bbW74N>+H3)ccRP.&R?(F&1.K\X]eT.[Z\93BGK_Bc1.OK7+UZa
eAgL3F&HRGX[1f-/7<_MS<K+^6dUNaBeM8dXSQ&@5TZREH@WBJ<@#]6<&5Ia4HE=
_)5B3[#.]4c+SLIR/ZZ/gN8&81MQ1?-UHV@T;+SXLgebKfP,X([^GP??ZfTK1&V3
?\NOGG.6&/Gbbe5e,)E>+8,6MVK.b/W\8U+3^NDNXH/UQR)Ze6F(\L6RceIFXCa6
I]de.V.),XJ0/]-;[dBYL?IS7NGMB1I(.ASd7VOe^H&gRU12_F<f3@IJL@TZ)gZ9
&DdA6S39gB+&=OM<4PG4d;U8O3^eb(E^+?)cH(C#K<XCE+HU_e]UgL/HA6.\0[[/
90QSEM4HA:E[<8,^[IJbW@Vf:K/b17e23IBOd,dDCbV_9bE<TT/;34#E7,[R@G0c
+B[:IH/R0<bbLSdI?_O,:-2Z^V9<7<JN?5.D6(GgdX]LP,8@QI:e\MX@6OL^;:JK
-f=(9@9@\0ae.PZZK^4N_#Mb&d:cBS9-2/]9X_g@5fUfO#_LF3G;&7O2=.)VX4XP
TMU,HSAgFM>eR^BdI,ZDQTV3WV7A\XHRZGdKF<LA5Ac.WQ]9L0d-Ac,QabUMc=4C
2f@V/DaeW^13,<U6(DA)<=]LH[=b8EN^7SJTAIWQ-WPLT#^KPM=[_YD+]1DYH;H:
M&>[FS3#8:(,Q<e--)O0A,#BT\0F<\L>T@<#:S-OJ/)Q,e[DM43_dX5)MfKLO2,L
eZDgJCDQN^R[ZecRc,I@H?X4Z3J7F/U)[,D<)GG7Oc=\-68&2N.UX+Z(6Q/>]0Q7
M65E9PIE:7KCIO#/7QP5^HH8?,VN&:QRd?.=I0U5C/V/KBSHcTX^R/9P08&NJP7L
X<PHTG,6=J+AT&M#+(-&/6557(9HV>7D6H]:D8W#1N9ge(Z/7)):N580>)2P+:BR
5/]-Y)N#][3F=7-ZL=c2CVPZW<.U7./:bW/0d&GL@;cF(KS46^H/<N#=2P0-]f01
M3<9V5<@)BbL5Q+MG[92B^Rc4><;/Y(2B+Ic[)_+K8J]&Z7gN<FWPNW4:TR1_IBd
O3MVG\=\;.,69T,,R.af1_S)b=dF-TN?PcEd_@(C\DE>E(aB]6U?cK^-J,\eE]aA
;>acT-=/HTT_]S[K#P:&G#LY>0D2dGZ\^)7eeZN4H=E/,^a;T4]G7FO;6YSd1:>T
K4;FPKRN>&<GI>Z@JP8,NOd[2^0GHbEVLLU9gOAA;#\Db>[TH>67(LV1J-GRe#:.
@g=6d(G=S2G#aK;,2Td=?C55N24dK]B\>3:X7aaH>baWIZSBIc^e4LXA4ff^QEWA
LDg9IGA\fABDc^#\6L.O5<#T(0TI1ZDb&PO4)L7@Ke;adS08\(.V8gX:(GA&9>Pd
M+G&0<=&=,&]YTM(C/4)RQY0QdI4UIEQF\9GP=>+7S+U/Ib;CGGIB^@WI:^K58]<
&TC+fY#UeI9eE=)86YcYB@&Peg_Z2;bSZ\#;8=H/:K,WBAfIJ=P:I=-Q/T)+I.Rf
DH_2AP72#eed+dfgE_GZc8>7TD&S,;X.>>T=?;N#H7Y-4EZB,Ma@9(>V[d>c=8XD
A0ST81\51TXa<IR9TB>#b[a\7(D7GD6LV@:fJ5O>c<JgeL3(7,a8,2T6Q)0=H&VU
WBN=UQS+I#S-65TI@1FH[^DF]d\:R;^Wg17T+<HQd3BJ_;EBebTCcB#1N/G]2_IX
[BIN]([XW.-7a&81[XU2f9_F2XFgBE_/^61Z==ScNF@+JD2P8@NV7CD<-Df5CN]F
/??0^#V#O)OX_<0W8Q.0+\CK\#dLgDE1eHGNXacXNL2UcGX:)91Z^1\I(/_T_YV\
.RDbX6TZ[2U:GXW.8X/DDPX&^5CQb/4Pf4UZJ6L>B[0K:+PN\-bQZHPB9B-^PJS=
f75YQ#OYL\e@E)_,#YS_FMPDNNMI8f8L]X1H12XS_;2@-2)<c9^?>@FEb?4[:JT9
TZ.b3Y[65Qe?T=34>ZCF4;?cOZ)dT4=&M+Jg)>_\aYT]Q/0Q:3.6@N^bMUN)GXGV
1:MMc4GF43Tgb3g\QO,(>eaSPT;O]O[?G(P]I\[.\L1fg2>bNfg7FI_[UZ2.CU4C
?Rf^eWF>AE+G,4dfK0Z4NbO^\@U?OO].4F]H>+>+G87:.8^9T[J:8@X5;CPY&\<f
70T)MccaE]b>\,?4_Zd5_1,Lg?RE[KRZD;d;)4/?B?,d.2(HQ)CIQ+\4f((Nf3I/
Y_H/HER9NS3fP5-ZO>::2UQZEFLG4dM5S8T9-&FNDMD+a=I:S<GR3_7B9T7Q1cT\
<a.>dW5b.=(@G<cPZcE]Q-#)MP>/4JHS8<BV2<eB6WYYW&eE\[;A&VS7R^TG-8@S
K/7;](;:_8XG(ZZ+5O6-:OM]/Z=\XF3.QSMOdKM3ef^bd.\?0..J&BB?-^^,[d9L
b3&C-]IWM?&TbSN(KKaG9,Fc,V)R<,K7e0=]P)[c^;MTeTM&7J+fEBe\5((P2f&F
36HI[O/8C:EEI:QbPGK4VQLMY?0V_9&C,L(0,UFO)BY<<e2/8KRe=e,EN59(4(IS
QN#N]VCgF^+Kcd..QI8@2-^?=[B81],X&HbI4Q=Q-D06XMR:]GPMY)V-6M.He=2D
eR27?g5&g);f:ZMYOe03gaHZHKR#eJ,V^/9g/Rfa/7T<WDbM6IAPDeXM?JL2UY+<
V#F+^G:)+R8<FU&?)?^B^_EP4^(JKfcJ-fP#4MDeBF@aRTS>8G/MRVeed0]_Q5MD
:5YcEB0dJYPK9:VSV])]I[>eY^?.#NV[U..B&M68\N/=VH=>3W7:RB[#7:V:S&=O
bOLb;f3X,5@bJ0?^b:#7,-+T41?/X&,.1#L9(8[0<7)4g+CX@S]M581>YYJIO3-8
S6#Z?#Q#5H73D,XZ?+T1f(f>d);gWL?>J&D)PPC5<c/BD,0cO)2,\Z8e19N?/=P]
f<..PeWMX[c\c:.9_C7:dCOE^HRTD[08P49FEVH]F@8.&M+C&D0&PcM(CReOIWR8
CF4;Z:a\fbY#0^:_=N[b-O19EZH2]R=WNNA;NRQG)7d/Y9eWCfEgd5d_7@PdJ?VC
/\8P]G_84RAMT(;;(YW&bJQ74M.8U[a8]8FcLZc6Y^;/E$
`endprotected

`protected
CWCbF,BI6J;9RbdBXU]V6_HFD(UNg>E+UEIKB4;P7/-(.]>d-6f=6)g4-PU(#=KI
NZ;d;+,QD?>,55,0V^^C)W-LWXYG+cO7g\3FLAMC,FQR,V0OQbQ(G&&2Y-.U5?+U
^?DILAAd#G4,0$
`endprotected

//vcs_lic_vip_protect
  `protected
Z4\:M(C&Ye451gIGANOLR1eG1EaMeT-M?#U9/#&\^?A)9C-dEbP<4(N.<d5UgG>R
/.Id(9]^D9e]Z2XX5<Te;_SE,?&d9a\=\(^F_5&2VZe0XZUNY3S:g:]=Y,;.ZXcP
6)U@GRI4]9g3Q=SdHC1W^XeM)TJ/QfWO:Nd,/5@]7Z,.U7aVTX:ef)_bR=T^Bb=U
[0IC3@R@,YZ?<MbAc^(.FD?N^6]DJRJcV7V1\eI#B1N=+Y<G-.]8a9BOXafIg8/-
.^??-\&J(ZC=eS9:Xd_X23RR>Abb7^EU5CECJg>SDR2,2]\E)9;:]2Qe_,G.W45^
?YXYOTODb6P(7L</OgE@VO]B<=[HVGXEXLRa,M;<HRTf-9SGQ@eXMc?O<R3[32gF
M8R,6//^_2XXC0R#\P94?5.0DYb[JS;[IQPZb)P;F@TgSe_c8NgATMN0_]Ba,I[P
?>OJ.T&V582EJJL2)P7EObO=/-8.#U-FadBO=e^fXd_Y;-1(^IDR]YF==@-=KF&c
TMXeGZ[H:SCe.HZ;ME(@N:;DXW>>V(\2<(83:[@(EM^C5O+/(-^^0U;(@?@D6Ya(
)MD=AaLf+7WG.\(W/&]<\.77:\=T(9)I#1+:3]0D&]dVPZLX;[0H\2JO5T8^(4VG
9/[WT+-]7;ac@F^1ZX?=:;KJFZ_^:-X5U3]WA&MU?]MNS9>IdQ&19ST5S07O=TcA
3\bKVO>S9+02d2<8M,)9PP1LHV]WCO=-9XdYNb:gXPGVJ41=?\I3?4DT@7WB5\1e
P(aT.8OU:Z+TUK.?&f<:<?56)]19:]XB#dbB0DcZ?F\a07PKPOST-D],WL,HWfRS
40WMRUKY-+VI/\fK.OA&\KSg_c+C^Cd4=B;@aK[<FX11_>,Qf&,TAb>?X8E,L/:>
W;B5YXc/V2,A-V<b\M.ab,WR>c;^_9&[&LG28I4?.M;B(ZP[\EZ+Y:3BaH<IJIaE
eXUT0T8gH-I3+@e:PM0^UT>?)>>dB+R1FHGD]+4N)ZRb-He]#O15gZY\dD0/E\JO
)?fXUW)f[\H>YD;P/+NKH:?&6=FOJAc>8<#?FJfH4;2NZdGN#AX60Y.>0DNJ.R7N
R?a/gY9](A4/e1#0,)2>R=^3U?H;IeUL(gS:d]BH?RTD2X<,==2,E2WQKE>\#0GW
H\Oe>Xf:B9_53K2SDKG9-HCRga@7Oa5JN[7@:?]H[?S.bU7PS^V+VO2&-d,.H@C5
0GC(7aL[B<K2F-V#?HfEK\#40E/QgKgZX<KKdS6LXc?T1#bQbS59\a;-5;;fU4f,
HZJM1&B\P>dgfg>.Q?TXWG3>MFP):DM/[@E,<G00;U^Q+@0e,]O@+9W.H1?T@5X6
WM:4B7<7?37(L&X-6aN;B(bdU&_DY@L-)A3.X9X0cF@cCWR(,g@a)O391)]N-T=1
gZ/V=-&R+B/AN>+#_[&>Pa[0LAU0556TR46XGdT2@D)A=LODZ5@=3)W#(]\4gO)I
SAP.P,7[HAMVDDeVfN?LN^Q+D/&]^9513]cO^_HQ@AU9b=VOLS,,b_IebGJ_[3XA
P1-?&J=([9@#93eYf_6DQ2@EWI+VFS1-DXJ,)_4?,Xbcf=Y8G:8.De3g3&d;(3>H
6Z^:;fZNE&S=R[;(@/N0/P/76F5NVc(G7U_9+[:_1Zg(.OgSLc>3_V9Z1J:,]S-O
DS#__;M1Lf]UY]=4KW.Geg8LVPacHa&RG&FR1WECecO@;=C20VfYeLd9:TfQ2FD5
+.N:6;HU/fVbA:#0IS\6cD+KNb8#SG5;f+L@.796&SL;H(?IIFgX-2(;N3V3d_E7
T2BH6Y1S?X0?91>aE9WYN,L_9Od>:PA]@_A^O+\V9;[M]NWA)HEQdAR?1B#\\(2F
IX2(=Rf<aQ#]-FWJ_CF.d8ZDETH.,[5J/].Y#^IYPLbScS?L4Ac/</c#Na3RT6cH
DfT-KM7K]@GNAT]-a>>]?-C(QGA1aRS:28_dRM0bGTJ34cN[,Q>4:I9^T9W/M8=T
P3+H&,Q<A)O:3_#;-gC3^d<#Q,EGORN7aY7UU(;]SJHI@)V,#+GB;P6(HB(XI;@d
&,#5<)Gf8aX@<(&S#0V#Hf?KQ#SPASQ+g0T<5^Ye()C(+)6060>[g.A;WV>4aQ&b
;e1;Y&-#X4L27,BE&Y<S?dJB8T-18e3?2BKR@&Cf2E;\1E][DTP58JB(V##=G@2d
\6.)NYeS#I=327+g[:93+64&VSN_>ecKEM7D&Dd?U6e[43_7&N=;CcgLXCe@QX_b
W43+Y[Z(g-L/V#G8<9XaP]CPf6eL8K8:=:Y2+)<N:#UN:FT-d#4J6_NROPc\P.;]
/.,:F#YX?1H9F?YgBPP6&#<+T7T<80adVH+K]7\8P?]Zd=5OBL_bdV>1LT^ZM,&6
/=^VPVJCe9B6Sc5M,3^=FY]gKWY:86IIELIG6(A+GSOS#bZ(AIKMNRW->?39PZL1
MZGUCTBT?AX3KOVEO).NeXZ;RZR))3R;)T24^<=,ZBXH^Ba:NI;(IXED4BEB(YR;
IN@^Wa+(b.4-7W6;=KS)AbM28-3VBVV\-A-R#?Y>,DX?7c8?XO=KY=N3BG]TN]<-
3]0[cAIO@SSAe>N\UR4gX^G2,3_TY3XGLd^g1I6G,&f((]3XRGfM=J,:@AEaOXWb
K+7&6F[ace/GcbH[91T:cX^bPYXT)@MC&&e07C+@(=S#.B,7#8[I>PV:XZDd0FM(
,SSXQV(FYE\L1\b(AN[G0MCBOXX)Td;EQO&<WV2[RCFPDfUc>8cO/+&Kc7UdPGOZ
9R:=)cM:&[@I2QPM570.M>YDU?a7)B:gRV1DDEHYSM03b,5b-EcW,==W\B_#QW=U
FTF#D5S;\GeUQIQ--6R;X-XZ:TT\L8VC^S([U([P&eH_?L+9)-a)-XY;7beE#^L.
L4]b(DHAIdX(PN>GdBcJU1F,g#E7..8cSK573N3C]S16^&1N0(DgRAKY<D@E_22,
g]R1A3TfH2OOYIa&E>C-._Zb_084F^>^Q03+7EQMI,&Vc=&W>,^15[YC(JQM<YH#
;W)C\ObS2D&e9Pb4RR/=N)e_6>>1T&C;_.A&K2YB6-W8[/Z:Qf?O<06;)FgdB-5K
V+#f:;^K3\eUU@ID=(A8OQYO6Ae24:DOg5N].b;K32\6(59>e+Y.5A;?M<_@2IIP
Q@8RVFH(1YeP-g<Q;N8EZ,J5MP7R6&&]LX-YJVC1X<>[1C+6K+VI1RGVbRU4?@H=
XU(5H,I_4DZP=J+;WJ&@T-U23/.a/D)8e^PUWHe6HN>U^VS#=)V2ZC-;Z)M,K<Q&
JZ1P,]R&KNKD31,TTABKB]dTU13FVJ=70ZE-9>89^M0MXB1L#eg]Z4L<Q6P;5A46
,>+eZU36#Jb\:6Q<_MLg#.?2@>TU_+bS@bYb>2E80PMFVPNC(##QGDV1K>0_e,KA
4DV1+7\g:LWCLZ5AZ3Q(5Q6a8cg]#D#X^RC^SW-8,:I[&C(E_KTIU95:H]gCS1YH
dOfE[];YQ0RB@MZ/?G]N/f[5M<8NZ]J;:S<Je6=?HOR0/g@Z9Y\TP0(aI<(P[SSZ
UcKf3=]+;VG4SeHX6S2)M63eDOMXW\b2DN44^[+1_[e^HT?W9MdOF)2XQda#9?aN
Pd(2MPSH8AT^R<))?L.e\&QV8,K[FME31e.-EGWTM@41EDHG,A)b;8d.3-:5,eSg
ZeQNO-_55>U#B]V^AMa/Q6@@DHFP1T;LB5B6RMLW>NR]M+G=,(aDW0YC+)0(=&/:
>YR=8X>JBc^/#=,^2&=@9eS0bNY2()LF/0Q;O=d/SfRf=cc=K+_LK,-;@Ff4&@NF
&@Q:PFP/A#(4F8H[CRX/Z>]B)I>d7K82C2MLBME/NW:Z+4:^N>Y3@3,QcHGdJS;?
,+8+E&:^Q;gG=YSY=X,\d6O;&+PHNaQ.]_,c+a8\g_EZG.295L,eD^/S#@cJ]\P5
RCCgIN?[KXK_,MGGJXeZ.gU1S,ARQR+MeNNL&/If^e/#M5V<8.e=cHe?Wc2^N+34
B1^XS/HGPX16)3GcP,\IK]AMF3-W\:2AQZUVB_2Re8KNS<EY]3fRSM#(;.eeYL)a
RdJ3YDb+,QO_e>2?gDebL\MaR9\]8HKGFa+Y1X_EZ&^(LBFM:BT8POa.SQEGMV(X
Je@X;/ZJNe2<f6UI9EUWa?b00gC(<RL;N&4UOe1TGRW._^)LKIVLBb#-)>[bO<0A
D=0c79N\;JAE=Y6\9^MP^G&D/VDX)5/-1LFc@;H&?[>-,AaWaF:c@E52TTH\GZ#G
6_f\[<LH5ISV\@1P7W(/1.J1>)(6@d>(,(\?F@8ga5e^++>5>/:_@#Gc@X1Wd939
8KR3_SN:0)EHZd;H,1J5.K:WB3Y,G7E7UJ)@BY3PL&J3A9]g<)<Q[ae@:ZSF+dR5
^6SXCS8U8d:,(/I=_JY2\V7CNFUaV;K/JggO/2FKHa@cZA8VS)T\2Z50D41bBMS:
7)TUZ@f4P]<e8eMN6CfIRY0E-cW;JNfdLM7(X^(7)VCWSI)Dbb05JD6G+BbZLR1U
JCP&Q0@)CZXd)+DN\g,>N2WEKQA[6RP@O&X>8WH)7:2Y)M++fHeVO,91I3KRD5#4
N?M:Ka+0H/^:JZD(T5>AYW=_L-^QT;;=VSO;bO\LWgV6fY3Q<cTL_[5RP[6dAWSc
A[;\QM<[FOUYJA2_E^EY/fBT^WL^]J9.=;^Y2b:-R&dX107eW>)g.#Q7N#+ZQ>\0
=RM2Z<_5dP_[)0BSeS#8AP]2aZSZ<28S@d<1MB&..2TB1IS3(SIYB,\D6(/@Y(<G
fV2R_,OQ^IdVD^Oc?0&(+2f-QdC=/dO]1E2MOPNI[P1PV@e?&=>6CQ<LOSGZBaF>
1/QCX.8bPKP3=KI1?YDSFb@=B<PL(2+@)EgVIb]F@0bZPa]3:dWX4cDIbgdLVF\R
S-9Y&&1(VXKDfK]KW]1Bb.,:#C^<)Jda?VX<CAJK]//d1W-bFZP.V==S-8bLA[Jf
QULES4bGG;a6f;^S.bX6E3N3CM[3DQJP:dK7d4:5eMEKX@H&9N#:,G4(@B6ag__4
>C4.E<:5QO?d,.6TQ]-#6>Jb_>9.2AZV92XI3X1<Ca+UF0E+I01DW5f)0KT/.(O6
b<B2AI[ggC\N[6&(NL7M&UW^G8^1<4HK>^[=0WXC.QMT5@L9#TW16^,c&\&-&5^d
/\d@RS.6YAL&P.8->[FQd^NTY:bONTa=,9AO8J]M<3JFB=NEdLG0X/:-cAONN7P^
[:^PA^Z50CAUX]5R5IG(/YD:&4T[RTR:(JQ5=?4))Ib[b6aeKWA\RWbbXXf6ZUd5
E]>(YTDUHN<7eTP#GL_9;>/&DK[3)MbRVY/1YT6BKc&a(;^1Y2g8G.c:RK]aKR:J
CAcK-RE?\HJag.DNdHdUD[PeKOVNY.gAa5O8\/K=:W3+BcA,f[Y2J+9IHA=)\I6I
ID[7@4_HT0:QO,W15XHTG3VO8Y-QM:NS>4E7dcJcOaL5HB\K83:]g1<QGT#^1-=9
7JcUT/Q3EZD1c1eN&\^S==MX)2cS+L^572RSWI)dTH56PNAbC429MN+O:cP+.P/Q
C(()=Y]C20EcdP^TY(_#BU4VCR+(GP:H.+21gM:Pa:LDPQ8D?K9Y7SG0J)50@6C#
L)7bKWNN\BMST3GRVf]6Q^f?U486@T078Ue6Sd[YgS>5dJHUb<_8A\RMN2)V:3Q[
\=(J<(1C18E/=daO5<bg@KB@TX&Z2Q6+URaBUA,V+#9CU8UNR#ceNc]4,<Z14@E2
2EOD3f:f)Q;J?67e2UOc;1+]4UYRR4\>Z#FX1WCeB^7cVX>JLWJcA&VJ>f(N],U>
1E2JLc(AM&fNW5<ZI:D3#fKN5D2GCO(.Q+7JQECPT(L]B,f?BG>S(aIE;Y/1;L5Z
W0^H4g/g)>:1#VFM5NcY;V9,a+B&OZ-)BF[?9ES]+\B/6#NQAgf.b&3]^4[[eM:U
UN>K]7&a;BVF2-OB#R__-_)I[g(3c6IVWY:]3[F&O,26bdJLS/]9JX+8Vc[J(H&X
+g<\XYaR#<UW;(@cFU)-SMc1-K<V^O;6896W92]F2<7@&Z<J97>S@7((]F=:W2L1
#LaZadYL6Q6:Ia+A)/^;#T1AXSgO<L78IC_)5e9ATY&6SCL^d58OMRVE,.cYD+#c
)K47,CD@O>;Qd+gCefYYQ6G5NFZ?.4:2a5^NC\_WDU/RS(CW8DG-E_(d@U.E]HU=
/,8#D7/YVM3KNPH&d;H0U8g#6S01<<-MWWBdeKM)RC/;)XQe?3WZMc@MVRLYSb>]
(8VM&JXW(T]H7VD=U9a\HFc6R]+-NVQS6FZ(OQ6A684,4/aYd9A_2@<Qdb7aAJb1
L78H\F;+;cVKR7M[]b]GN21L0&]=SM:0.=&1eI#W0]NNFQ5Q1:5YH+FB&?(fND3J
,Y[_:X#(ECKRPW>N^F8bVSb,O/H4dcYMFQfUgQg9FZ#(g8WEP@g^[2]g6((a+d#X
g07?2A.:LS^_TRGB@S#5#a_gEg<34]N,/:^#2:\]JXeSf\LOc&e;0C.6]\<R(OY6
TQ(KH0G\;V\&SaTfRe83P=WAGX++ITZY9_MQdUYFYF@Z=(,U-6LN2gQ4Z/CfQQdf
b91O)e[?VDQMV\/f4E(WC93DfBb:NMJ)W7:,7c?=:N#EIc:G+&gLHY0V+K>?CC5\
.B6#^:aSN1--0de>/.NgF1[;9BWE-^<F7_RBcgICDBc)g3cM@^&g55Me]beTQANZ
PWM=K1G[eCfAY\feE:/VfO5g6UVZB(7_ZPZ-(:U>&dI.^;PO.+cXRRL7NQO3BS7T
-Y?EHVNf,KCG:f^P0XY\(7-57IbB:9IJMbbOO+XD?X&8=L1&F^_;X>5R3HH5AT3>
KD\G:g>d=;+IYC@+Y0[58deKS8I8EaT-Qg&g=C4(0E,#930[9Kd_<_NM0bQY&WIS
WBb6<YCdR;\8ZD]K4d^OYCDT<Y;dcfa1/Y5M;(M-I>_Y]KPSa3FHUERPJ/6)VK9e
TN?0F@?<G7;6XR:/[)]3.dPR^9];CZ>HQ,\<+C^:>W&7<^5fGVF;d0TFM0&e43EX
@&GO(E(U,):S0E0[C58E/&5:X8KA7JU>U=O^9+QHdfbF8370S62@)U]@YP&bEKWf
?Y09(d[:+#R=IM>7(5Gg_JF;.Q3RM_.D0Qf2C>,@PG/>6>.^(bY5^:@P\dE(1)99
f<]N5f8?QWLeWE8=LLBcVUXR)ZWAf9PgI>UZHU.V>b\,<d7/##^J@[O9(#1\bMAe
]2J>1<N0H.Ub2c+Ofgg^#/O-9+c])LT=;af7AdYW-X7EReS)P-K@\2\(\;0YSBGL
U0:Q2DX:,\R<<Q+_GF2#c\2-Sd1_efA^R5/f;&ZJ1\::f99A2H1.LZf^VQ74>58:
eR=,DLZLQO;I]3I<1W8OUG>_>RFP+eVQB\gVV.f8ONJX0Hb1LHH)\7M([#=e>QDK
1JD8&_V[P&2NN(][RGJS]eB(6ET;Z@aV4>fA@3U(Bg[2f6KW,b[44XK#[G5/L6<P
/8YZOg#VYWcPPX;Y5.^dUe,MNYR?)[W3_GCEWK6cX_;VDZgDA[.;V/KOH8-9\KJN
ES5&K2>S\XLc1J##7^0#KS,UN<4_F^FdVX1GJCMTdV\9S:_L08gV]U:DI5]Ya&W4
VcEUe>.[UbSW&[Db/RZVFOUCgN8TZEbKbJ1)#bXOgM<P9&R54)MNT1F<)RG=HX7H
7E#C6-QH^[b-L>I:#JX)?f:EWJCgO+V.1H0[?4:E>,VV+3/?2[WN-[gSb,^L.XGY
^M0(g)IdTEe@CAADFR/=YN#O+F]+L0F.VN[]@f+OB@-V#]@Q;cE-[aEE9<46K9\-
ABE^M(#[?;E[4dHA0LRA]YRF5[,>2X,.NQ7T,DQ1G#<8#JW86J4(RL,L[6V^XJ;4
dI77f)MR)FaW-T&IYNA\7M>+b,48:+K-G]J(C@WNg0IDKf;eNDbL\Nd#E@=1J73<
BH#[BMda&+AQRRL#6Dc-cP4A8L5TEdaS904<64&\^Df7/-gMGT>\9-&PN[0\8(+1
->0R0FeF)A.KRJf&H0[<N:&=McH;WUQ8BK_&cfPZ^D<&)>&:=0I/.C32/_@eT.QX
44,0,[:7#MdVgK-D0aW(0_G8MFS;DEB-fNA^_J,[^MEW;)e^XgD.e(\e0&0(eZYV
7&KI#dN(Kf:[=7dQRT1+5H5/#USQ8_RW+\::N4GaGI35ANU&8#UCBN_GOGcO4G2a
P6[A[7aSb+@U)(QN>_5DV,/-ITU7;Y#K:H,<X<0gI@#HUC7J\ZR3PK5a,NW-g)C.
M[:L1@M;B1D5B#K85>F7fI=YO=C7<T80-50DKR\G3]P>UDJZbb=EPb>\MKC4]_FJ
X)LBQ;V,+#995IU1YZc]9W.d]PB]-MQ2MEga=9.Y01D/H5M0.W\YE&dOT0XW.DC5
?,OR;VFc[Ya)\,Eca3=FRZ2,aY,1SWB4/P\;C[0gWS9e8)C+f9E^D?T\e]#5&cdP
J?7:T?PRAdf5#JZO(S=@G&C.fcV/3V@WLE_BHWZ,W;cTPTZHM.SMcfC2NW-OdO3C
bB#5bJ^J3H6<,>;JO>V^RBG(^CRGS6\)Z]COS8F<<dI=7ecP3N<21@&[CO8&WaS0
QYQQGXaPZP&?Mce,P@PX-:.:&J/5fIC\F-GO\G0G^+]+dgEAJ_0X_#OAK_MULg-=
EK^^RX66ZTK5/Q:Y(=_7NTVSZ^0CX66+-C)Z_KR8@9[_24efK3Y2\=ZZ[b3>X[4B
_C1@G@41^XJB.=@7=Z]V)#>SGR42F<#dL(:##]XXdN.A(@He(I1U.Y>??<)g-Bd3
:e>@CATYEc+e(<:\<g&6[KE^)\;AG@7Bg9dRXX]A3SC5S/7PM5FbQ2R]JI6e=[bE
3H4d]QH?&5?cY(T&5+AQ..PL1EVX<fcN0(<RNR81\Q5S9;7Z>DKRE3]\J>MQ?/(B
N>]D)W<+gF77>bZ1D=5HR_BT^ON=/5U9@Oa04\1&QeOg,4ZcX16e<T2eL0D&[,d\
Tfg-eQ6B)IY_Z<4<O[c?MP/<,2GAgTW;dJdNG7MC/?5I+Q7(.<\18N7Pba/QbRT,
7[aQ_0M;L4\#+1Je@V5N1D6dL1]KKTf+#:&JA5&KM66?;Vfg>=@JQ>U9<G>F>WBS
#QM67MX<V&#2/T;#T>FT),\04IZ4@[=0U7W84]-[5JC+f^=4TT\:4R+;077#LF&O
0.(2gdRT[2B>&D_&4Q[_[<>36I:H.:_/f-RFYE31e\75Y1YFZ+e=?[Pe7Q1G8FXH
DCYQ.I-ZcHVKeF#WeKO1A/GN-X^J<S8C2+4:(_?-H<:@<QA:V#=HSE60R\(BX=[5
J42>^>9>^X..<F>GE-#VcaI+O&WWP2HC4\M7e0J#BN:e&6,\WcSKVYOB.__?9IC3
.a>2d?H+Q\.AI4(ILQOGN?M_cNcIMJRUeCAOEMMeR&Z0W?HD@)QIC-3LD6:N_<ZA
:e61E1[#2#7\5(AQNK=V8^P^d_1JGT0A6R(NQ>6JXXUgWGE10_^4TgDXVL/2J5TA
MD0a.M1ed1V2T_^J59e\J=?&)C3a\aC)L;/OVa?F3[cZU6d2==;QU8/T7PG=1T;R
a)&eXZH;9-UYB4Bd8BWOS?c&>8af&a>F@fAOO/+?R#??X&+7KPPB91K#PR:3K>?\
WC++NC-eS-M9C/NCF0/Rge<[4FW2Q.R>4dDE.@70(#;K.A6ICJ,H51P1-648Ye\+
X\[M?]SHX<^2WG+_0Y@U4YZD?f495<A/af-?c+?+J_RD>]3?CdEK=EM/.FL,&+UR
eYK]XH-^f0C0L7&9H^,6G9d-IO8(XFdg^=Y5?83UD@TS].\QITOIgJ)G-_&=HY&]
4@[GcbES#NX9e#KT>4M<[2HAbLb&A85AUU^K[@dD6[B95&IO7,WZZ5&<4BVFCO2A
4<.5T)Of<f]U+TM?E48R9\,XT=6[1a1ZMT=d[VYNMJ9VZRHM(HBZ7;E/X<DUD/=S
HW-A:2TP.-N/&b?]DW(_PdD&Q&PZR@X&/94dVaYWP=@D5D(&<W,^2-a6g1,IB>#-
=99455+9d<;HJIA=0/3J9cKdMIf9V[f.>N1,bVFIDV<7PE].aHG?3Wf=(cE6f57d
>OYH6(Y#,5U[c@_#]ZcQ#C0Q=5.X]6bMDPaP.15Ka.DBCaNBT8S?>).g-@7>(Z9I
5H8]54IQ^;@S#O:4RH4\#)LW2BOe#8#E.YAL1:LA=;gI(<LX#W9XL])52ZI^LOg#
=I?_39eMD-(4Y5;B6/H<.:[XH+7L&9C[dMC,73;gY/Q16^FW<F_+7=>6-HO:(d.E
@)RM;IU/fS4gIVD-8cJ5_[JN=772<g^HL=fU5]Q87;>U,RPJRC?),VTA-#,J&;NA
[^b@AX@dHZE6ROZF9#=>Yc_\U9g0O)B.4c[f5OC_61-6eQOS&H9cDWg?^Cgbc:=#
Ng/GVfN-O:6c3C^C=PXKPWHgW.H8^fL-f^6gLcCPLQ3HI7#0L;7bG:O(^c39FTJO
<\1.)S4+G[R):I>GV+IbQ<C&gZKaY9D@a#G?LSLNe^Zg93D@c4):5GT<8KF)_ISC
HX\7R^X/WN@?76O[?@&3SNQ6U<4Of?)C>]_GL(=,X@PFfNJ)#H)Ra]R)EJ;./?6f
FI37&)EgBc,d_ISdFEV637D2eY+9:))ES4NI+g5.g\=5C.cNeZ=13VJQF9Y8GI.T
#W@R=NC(/AZ67,R@9;U#3\,e,HRbPK>Fb/6YUe0]2bd-P=+3cB&@A1YRd07TNR/T
Yf^M>N/TGVB=XcDBfd3&)?X>,ZUAUeZ_?^[=ZF:EX542>.QPFSK.DX4N_&3L9.[)
U?2;L-OPKLdS&EAMQ34EH/b>]-,TH9d0;E>[L#b))2e6<)ZJ6=VG>AJRU<4>>3V1
9GKC+If8)7d\MZa_UdZ]O?UN2eHHSRH1,W\ALFN;-XWc1QZN>ebfN-.U:M40QPNU
DEe9H8N_DPBJFIP9UQCV6W4JbL:D9)DU<I)\DOTcb9P&SWWZf<D(NPcWJ2GK:C/@
cV#0=::SNX?Y1d>Y[7P<B1H912_.Q2M@LLbL)8.=19dOPFA=Q63<4.-Oe[P)W4c4
TA7#C+I3./.b-0XAf>G2DX,Af\:;B->/,CB2cW?BJ8)[G_>aB]b00C4B+X>[MXP>
WW5,dOYK^^aRH6SD<gQ<8aZ_#RcD(?0?SS[^a2/6_U>A8.(4d1I=T2,M@S@_8cDC
HF2SW^U1(\E5&8)0WD16>b-+2ND]Wg[?^K84^7TV-(LR[,?O_(7Q/G@[NV@+103Q
a:2eKc7R/;A:D:G\]40,(@Z;&Pe#S)(U9UB4#f#CgY\XI6:e=:WCE3O]a#9:gYVR
NN8S8cQ4#Q\M0PH9SNK3gG+P.S/D&..dQKK@@VSg^H_0YHECb7#XL,-&fTaA:04Y
GD-FFW,<XQb_;3=00-8(B:C&6UQE9H&?U[>5?ZX4E>=e<GTO#P4U806?(Q8-7a9]
QN4VJe8CZ<;aP73/K,==GXHWRO\G\.a(>3YGQRDOf.HEe=+aYWCaY2?=bLPXL#F:
<8>;OG,V5[.S]b;B]c&TMa[V+E,UYd,U^.NfTQHe=L:D2ff8>MS;1JQDcGe&2;UV
:7bTJI@/KPUIUaXEVf)=JA5bMANU?gJbL&>__DK6R0Z)P=Z3?]@eEeb)@Uf06=)-
6Gf[H9)IMEJ1f&/Q[OY^(eJL6fdW<Ve\\F2R]^fd=e.F4dRWV6\(ZV/+MS/41]S)
]4Y+MT\,E;[TS5AF)F;-8[\XZ\S?:D;-0PN#6LW?U,QGB,Kb7\/>=FN?GLV-Hg]d
(>FU#;A)^[R(e<TR)1R7O#G:,]K;^F,g)G^\L2]4KCCfDceeI/&//@8PBY0E^Z0D
A(9Y_6?a/JPI_H+&]cA-)\#(9Y745gR8L048EYfH#/+59(F)6W+=fI.Tg3R3BdJS
\>R6f8L/F44=9e58?bKJIOE[LHfa8#H.QEF3f74W->#c;VYa>6gXB/,Y1:4J\]A-
9-_DH>D4Ne/7cF2R[VZOVNBgDI1THE79SV^CfM_@-C;+T=H&+79(JE;TO>b[/V6J
DcUCG#QJHZN.C4b929^]<KfQ1+5JgJAX.(UM;]U/S9>4=Cg0LV_=N[Ca1NA4^A?\
,+WGP[8SXb+>F1A/g=0gH4/DOED_JTJ_DTQE&(cO(YC:VgC+8-<BR<N730=67Jb]
cC&^e[U8U48bG93/\HLIAHd,6f]=5^Z\.OL@^c+cJ+e^Y;-TVT<K[@@A;9T@86c-
QC6\@_<\>>/G#<KOJ7T3b.BZ,GD3d#X>D5QC(IOd=NQ^<U?GKaP+eeH8DH2eG_Ke
])a06J1)2)46QT7bDNTKB]FEWR)AabgNW6D5>U-d2BQ4XIGgeID+J+]ANKHQCbRX
BC6LN=[e.A9gZFBE:>Z.YbEJ=22RF?#PDc?)cEJG?/J+CQ\R&VPMGD<(C0Y@;bGF
3YD@R^QT_[0e,R6-P(887_Y#_b?7G7\J-FRZ/I@^#R/OE/A8(YKR6NGMBXS76EKH
-]_&L6\XDaEG)OD^YDW&0HDI8,,G(U][dNZac-(,NK,=KgSB\<&P)G>f\eBb@.M\
@\Z,EJ+F^P3f0DOIf2R[&b:4L)LG5U2BHE\ALV+d_H(-_]+9e0^DQN=4CZ:<,b<G
fGGY:60;3,O4)5bIOTJ&)d.dM=(HG>G9J<b1_fG8ba3Z#6=>&5</>dFQIN1eBH:Y
7M>T[J7#g8(HYUgTPE+>MC[7MBS1>A;+fVOg[&RcE;;L[\9bRI;HX6g8BI,#gEge
ZCNRU=-M]+<LgMIR#5:7,QL\X,DK+dP[eg&5dLV1,N1HEcU=86HMTg;T1e,bX^TV
0M@6GM^G/Jc3d(3[E4\-3PE(86RTV2S8E:&UfJQ.fQBA]P&:&VF<&RH0SHOGEbD:
6(C=<f3ZSNeV2_H-VTBMZJO-+Zg3W.VIaAg1#_(WfO)U^0A9OY#G-E3[6][@,7SM
82IgDF7Z_f6_;#E6(Z@b[449L=6fd6>[I>PMR.TaU9R=98bd)2X3JQV=F4R&^d?>
QT5dW>QB<+R/g5UgHDPMI3R(YAFGFO<_H.19f]eaKf&[2&/3bD2)Tcc=Ac06eRN/
@UAPOc=d8F\I(/4::.[D,)K_#G3#XJN+[,/dX7]9IA@3fTD_AKReVZOf@@PO+&SS
#X^(\=)P?F]B=\+c2Ec>53,ZO^82G>bb#06ZBPD[3=E5C8UG,85XC#aNeD]_?J&F
<J7OTYEX@(5Yb7>D4L(?e7_7/(]EM-0D1:K5HMG+1Q9&7_b5&M+<[2\I^=ZX_d(_
?<;/>I>>=\7@6_\6c\2&Q59]I49FGJ+<EJF<.R.PQ-D2&P_M4Z7YXX\E,fKFS=QU
beCd@Y5S2ZIFX,_d:1(4WABKPgLdNNDKZe8e/9P_L<#)dPU8UXMMK?60?U3WEGC#
^Z#(5-IP4;J\FAG:^DYXa[eH9UEC_E3(6B6H=_Z>>YT2@J7?@UD]KB2B3TVCMYZa
>O#HB?8);O^.Y.>(-J96LKZYcg.+f<]@HfC[[^SaA:e-+C7EgQS1WS_T8?b<&1UF
+\)1IJ61HCfLZ]/+T@BBMC1B0\]5eL]W27_V0VGF?(7Ta3e)\)+Ud,^Wd<DJB,R:
ZDR8@[2NSWQVB&RC,<5R.Z<^TTQ:IB9#A3J>Z>GK+<WYM7TN8Ief^1M:C06Q(8eT
;eA_A@Dd4;N>KAa:2T5J.0b(WQb4A63>eZGPA@&Y>BMMR]QX^=d9(N]OWZPa#:&Y
dRZX_P2gY3@RPEV7^9+6[J<H@gTe3#g_3/QNH\&g[]<d[&/]SMe]5Vd_<SU^g/Xg
HX(B:g+(G(0c4Je7&@I5>QD&V1]CE[<U1^S-)YJ-)W4IEV3N1bTJA<K-#2=f]R_3
#;W[gW&f(JH&2]EaWXT@+eeg3@DU_/@9K77PacPd7Yg4V&:1AXMT@;-8L+14AW02
aWF)YHR.cH=A=0E)16X#Rd;\f]E2K=GG;TCLUP=+FU<Q]0b_C7@KLJXP?9U[LS_&
GB4).6ZHI-(=TZDB-XFZ#E/B_OGgGH[V.-148+#<HeCUZL9(g+X&I@E8#cGK7_J5
ALe-5WI]H]>SQR40KC74P-4bLe-3G7KMR/<Z@+&M36]WMD+?H=A1GFe)1((GAR)S
E\9aP<)Y9RdBT\6R3#c;2Wb^3^eJ9e7C;0e8]B39O&0\ZJQTTG9aCZB\+12W[[&f
WIJaNZT2bFWL7B1&f?L6,7PNQPO+QAXOC?0I:e-AE;@_2,eDA=H_BNN.4]ScLSJZ
f=Z)f5[(/\-]0Yea=NfY:3>O\GH.0K>IJaB5XWU()T7J[CaTQa>VTG(a/)5:MEGM
]K1>Z_R<JE4VaLE-fDB770_^,)7+7Jg6RQ&-)4(_=GNG[JJIgUdK=QPF(<WBgOVK
_5\_,46[18N-,VISD_986KJNK4/ebBR<a[NK\EOIX#B<aCNMPN>aD.36a=3J07H(
<2]_23eEOS6T3E9LB@E3K1<H9L_@6E.0\dI):PF<N^)D-gM][=P454EJF+.@E-Wb
0\M#R+X&,JQE>Q3/CFNOeL<:[;54E-f<:CEe\\HX1If7;a])=RD6_&=e0fBXK7^L
6#3Q:FE+f80Z:@53-A/=e&:\0X[FV;3g&__#WQNF0;2XURC#Z5dcC<IWeKA/Fc\g
@UJTCD.(@39\KV;OABU#W_+>Qg.PWNG[E(Y;7c/-.aY6OT.^>bJ0)TH[]-T8?>f_
1:@<cNa[,SQ>N5KSd2MHd-f,gW>IQ-HN8]RTAL\Pf\2^0]&T+VX7#2M[X.\FP?;,
I^eJ#]@0C6(aS8SYA+)24X1/[V8?8/gGXbV/KM.?ZKbaP-R:NQca)1/5OGWUc\cW
bK<V-Y=9V\^bb/(1OS\&[Z+@M1H^+eG?[5bN+f4cGa60)+S_MKK;37@_(G>E,a8G
,=T(84Q4B(B4\ZY;FdF^1=5AY\+eP7+aQU76-,,3ab#+UeT_,XQPP[#BKB,ATeQR
VMYX69c:&\[Z6dUR\(ae5EaXD\(+3/(72JEJ,A.&ZW[/Q4HdC>M7=Xe4TM217J<-
[(^PA893Tf?19<Tb>:bHIf.6^G.4B_[TL:+#_gO^,4a6bH613dfL.cb;C)3Ye4>/
?<-\FF,(DXUU7&Ode8YYJ:RED+I&Vc]:24/>?2AQ6GNQ+Y/<KKe]B++Cc2GcY^>K
0f1(,^-[UNc=DZ]7]dXFZ<&5b;O@B1B2G):VK\KY\O>,3@+6B0IA[F>M)^K+N>+Y
dBA#U3RA/D_LBO-N+QK]EYJR-:-X(U-2TT5DG)8bL>?@V5CbJ;.-eB2A(LcXBV)C
RFO4.I.YISO&<2(F/B999==<^#,0)b81Z.#\e>_IHd,@B$
`endprotected
  


`protected
dL\#BM>VSg.<2@6>/5M2FL2?b[Cg#@_NcE[Z)3:0X\V+S2Ca6=<G/)8bGQDGNZ(Q
.16;<bf[b?cE,;;\>5F>6_2?2$
`endprotected

//vcs_lic_vip_protect
  `protected
#9R)RC6<F2LUVHZg_OO65Id)U_c#7L5/2G^K]ePK0OGYFZ\X,L>;)(/a?:UG1I5D
QaMKQQcSA(e16Fc9/HBDA(LRcRL_6/cFEP+Z+(B</cQe(97Z\@O@O5,dZ0ZHX8\<
f2[DcPfS55.&Ob,fGdT/d_:C==J.Z;e;Z>BESb8QYXH^eHg3.(89713G#YgK]6@c
RgZa:,Q_A+N7(:9#=&RV1KgNfLaAf8A^W7Q1&a:GA1NX5:(H,2:_I0&.)?P@F#2,
C0T[\K1++@8HaTHHQ87&4#KF9\e4d1WI3U)+gKgUQcKAebE6BXP>XAF]>CZd(/>g
CR9>>;&PMgFbB1(>Lb1:^[_.HFc=T+0fJX]16-W(>EfX?D9CO3(89cBN]NG][^@g
Z5A>b^QPbHU8[UfL-:T?aZOQ-4UR7[NKNA#G2]B?TXNe@aVGHP5CMIJc?1WJTDE?
HLJJYL2dXQ[DX)\K_QDKA^>&L(EP<YXd<@Y+R;Z>\f/BP<+-Z?]XGa^Z;^J0=a^e
L:T_VK133dM1(Tggg>=fP/N/_[Y)+X<WKQ&<P(fJE3T6]AF&QLRNDeNe5@aYaa5-
3#a+1bg6FATMI5-VO_/C25OLN=Z>@8)M/<?.J.S<XPJTd_,GV>5X\C33dJ=(T=C+
dA]>f8?cA@C8>MUe]HCIFEAdNcTS>Sg+TC8W6.[P)a4&MfI4<20bK<EE\6VG?c^H
c;<(GAZ;9/K,TT90(3)\Y7D(be^JBKK5CS@N38X_CC>9fOWfS,)F#E#FSTf(UY^G
2bW6,B>X@1;JPbLGA(7.+\Ha6^K@/](LT7P;JI6\#>[:R(?:Ke5X_>WK.ZDADNgS
-4/^O;4@A1EF,<E8O5<Kgc<MC;J]_(ZA3]<g\^C)aHL.d?V1Q4YQ?2N.-?@0,aZU
d7^62(G:#0PYS>(K-9:<BSdaP1OX>T7PC(B03#/N2_a0N2+A8,SX]\[Z.HRC/A=/
O-10&H0TYB582<4Z\+HR;4a3bI(K-4QE;e@S>C&K.B6OdL><HNLRY)C3=6U88ML7
RP(WGI.?P2@/-+C3;Dd/FM=E\78>G\bQ+E[&QNZ/K<[A=?GRfXMPQ551QB9&.^5:
<;FE3(?K.dPMEf6I;D[TM-D2Y_P>c5JN-.@08]aUJ[R2G^Ge@-RHDRS4Y(+EdaFf
[#;/T]PA@&>U115#;GbY/+S(Re;+>R()#LQ^@+VLFgU8]U^=C#f/Y.dD4A4HNRbP
d-[]]911L_NgF+7L\Pa3XSEA1U6]O/0B9+-\6,@+f6EQD69C#PWTF_g=&>EXaDF/
VWDR_[2@#Q>72_>-:GZg<.]\&Y&9Tf/76/T(>)RFJ&X6VH[S&1)V850[36FcTA,T
Q>4X]_M0<VS.A+FT@<XK(dW4DAdUWJ]OO+9&DUE.F>A#2a6\bMQ<A.D4>5g)V/-;
>^/XK7IdScG3#U6Q1H2XL(c7YE-)TZU9C?;L_VPJf@-4\&/5[<[+dQOWIgU?NQC(
9CKD^P3MUT1M)7HgS^1D34Xb)?(R3.,YGPJV:V=b;&B.=]UB-X^dYDEEID67FRB2
96[/A2Jg&5T9-e]PT8>fSF<&beTS6deKRgDS832U/Fe_Y+Q@3EDd7WH2^@,+)B7=
TV[8@.LE[YNS]L[OP,CH/O@Q@E;PbbKM3]TdRYI(:[XS4,52=[?#\MbQ+A&_C3X7
N0c7XI_/d6R>HJfGS)O.Ye=c(e6TdZ\IN>dU/[F^X;\eBb[&ZDECZ9HN_=#HCGQU
.<[3TQ]AI5bS1D_5d5)4c27+X#U]ZVOTF?V&K3]N.G)bWLU\+,M]b/HbLfZ4df/D
OP@UO#7LT0Gd\e;(?M,4AG5GB]H5:UX_44ac\5?b?I5b:.F,>?_5UNL0<2:\/bB?
BeC#Z/NC^:K+GH,DZc>=EV[-8aC=#SOBRdCKT(L8)W=QK8dMARF6R/V>XV@]K4Uf
)XB+CSF8+N@1#BMX3D&OX4HbBS?FDMTV5.J54?@C+^_;-e6P+?a4F8DIXDH&48.G
IG57D@g5&b<O+V2&]VEbO@2c1/F5PCN_I,9PN98^b0OMWM[J,PECC8K=1)B.D[(3
d1JHB^,]=L+UU5d/PBd;7.?/[92&L+9IAE>WSWX>1C\)E0?1==2Z=TI+E?8M);W;
&aP/AGA6g1cW1]dI5+V\_WbW)Pb1_Bb(5UEEU^[Rg:(;VG.QFVB-@1T4Q+G\F/H=
FEFFcER-cc6e/+27:G6U\A:7FON7+ZNS@a?GVF3:Q1RT[@fRIQ339gTZT]_6?A-,
_@58-UZ_HKGPYU0g2=[6Y7=UB-12V[3XZBe7)b7#A#EL28b;9G#.SR^0YIEIc.IE
Wa:d\,Z1@S?/Kg6FObP_-_a9O_gXf:^8T@]O<64=O&Z-N[?\LJbR.7[N,gP(1Lg+
T24.<Paa3HUF4;LA>GZ/ge[?KMM_YKT-/<L8dU2C2)d+aE6X)Z9RI-Q9=8F0QY)O
9S.fE-e,;2&-+\>CdZ(.F[I-@06O/6M8S=<FLe@;T<:fF/-.@JBO5C54e<LW4\fB
3?G@W]NMCeRY_0T46a=Y(U1334bTeS\OY[IBV@/KSQIfU-[6&YA\\]G]ZS1OCEg;
9V0A/:f91>OPLZd(fRV#PC5+dZ+=K92W^-ETD@TXg.#[>\]E=@;D6,&R1T4AU:OH
#<(/FJBLY\)RPADc9=OaY,=H>5Rg3KJA3&KBLF/eAXL)=4-/,IJXOKdXQH+?aJHg
>g1L1,_+YRIa,]0MZF99O.(U8H62HTH:S;]3?AD9IY8L<(CBNX/@^=CDLZ\(eZ.=
9>)T=2>)GCaf.C;AD[FJ\PQ97]>RGLb,LcgBC2Z4/BeeB\?@)]7Yc1AB3Y#G1;&S
@+Y(ZcM[JQc;dQ:;UcR)W?fEWg)4.GO/fL]7Y:C]O.Ya;L.#P1/QeC?XR?\/e0gE
E1[=<Q7b6Q^RSdY\1W8PXE@Nf/UGZ4=4e])AY7?;W/eL^?B[YeVBBI9aZ\Q5d8,@
0U\SONI_197U@_&];MYe@=Za.C?@,LUZ:b(JA12U=0Y24MR0NXO&#CM4O\FL<C6#
2[C^12(_/8;\5;J](3C<\>0#<PI8XZCSB_T)CV.HVN<KB<@6JHNA0S.QQ0RM+7P_
/@H(a91=MbV,eD9^OCcB\]=8VT7/9N5&3\C[1ZYER.-50J^VDAETU9)0G76DAF)N
SNDK;FH1@Lc^D/a#L9+dDQ#c(b7,;;d1^4g(Q;TG7T>G-TTB4eMdO;5O0Ze<<43C
5#<6D1Z?TN8SS3#CE>R3e_]OT;.A=ZUF:H=CUR1Ic@UQTg8U;I=Y_CC_09I5]2#5
I>6B]V/D0M?^XD-2[V1Ac=[I<IUNa^+62HX;CF>=R>O^OK,d.?Z7HG;;^Ub/\VV6
T)4ag/24X..@2B/d+e^g-/XO.>fH1@K\=Td[6]<N]A@[_bQP5=\]I=O]B,8;4(d1
8,9eYDVdfFb?/UZZC):U(5.c^B;0I9dT;YX[Z0[G^:.332IK&]JW#MXCIe3V7N0W
EbEK((+;c)O)Z76=PJQgV<=E2(=L+2C4PN&e@OaWBNR;QN8&a_f7LR;UG)bAG\&C
XW_,;&,L8XOeCHS4Fd)=,<7KU2F>NXeWcSLEB@<I03DL;e?V&2IBM@N6X5(e]=25
eJ/LN)6Pe<.G22c2&V\OaPJO0_<[P@ebLG-^@@EBNL8BJVCK;-067LgMeL259RZg
Vd+^]X@e6YS=W6F2f7&(eIT0)CG^_SeL2=Z/2VCdIb_Z7=Y2P3\;(<8T>980dNRC
:1.D;[:^g.]LB;#&;;LaQ/<)6R@/:1A]+\F8JU\,906L2d9-I#O#/]:d,S-MKZf.
#IHQ6WJLZP^[)V5ad>OK:g4a@^QQ;c()7a+fY8VF<BMI\ZeV6F)2ZZQ7E7c8\Jd,
g40,L)A3>@cAWab[;0+4RH8H=aRRS6.QU2dB^#?HG&OWRTTJ#.YXGbafb?Kd0Q+O
f;2Z&2\<D1BL0HGRNf99?M:bD)UT66()<BUR9fBUc0JT7SLAgd8V4I8+..\V^V+f
d0/cMXN)0gZNZK-TSI-C^WTJcNXU<G<D4.+UgP\[Wd@5:[H[W3<Cab=1bF=GcTBX
RN#XfIZWF>fE^/I(1@1)>\>J3b81__dP#b@,a.640V+:If=LR_M5L+II6c86+79c
?g=9-,dQSWL\C+^AaX(4Pg+Id^[ge#c(W(F_Q8UWT0X8\2R#3]9c-0>I]>8<O+I9
Z<6I;WgaI_XfKWa&TAO[B89&KSO&GEX@c<Ub-CZ:/ZU>U]0::3#>2G9#6.e+4I)L
SGC.NGC6a)<RE9Pf77T,+RD<3_7Pc?.FX_S&?bZTU(H\>g,N1LX\CSLcAE-.J:7<
Q99)B]^<71Z]BHJ::+NIN2^^RJPNfCf7A=<NTNURYd;/^Ub0)g7>P(O6-T^[_J_6
E8ZMAL8)R0<))E(0SQ[ICA\QF+8Kb(b.TMQ;Zg/Z)aLW^/[M25G,RFc:K^[A;L++
US46R7N0Jf,-414c:UJ\5.=40HeKGP5e1_H?C:]S3_Zf7,1BT)_^_ST\D/gg?1,]
NBf30FW2:&Z^/ZSV47#P(E=)(/b1Eg=_0NX5^:1LO0]+GfAaO_\6YdVeJ44WC4d-
1&#fa[dVOBbK.JEH1g=5)dT5Wc(dJaN>37ZNa(BGe;,5V+_>bg6WaZb56=<ce9[#
T=6e8T7d+F]\f?S1P(48BTc5\f,cK;7>Q?-A?EUJ;>8L=g7\abIc(<J(,WQ\)8WM
+I<B_5-1H/I/5K7e@+_.Y8[VTXK3dFeJ>P0M_BbKaM_)V--(S0U+.Lc[Pd:HBVW9
Z=&_[C1.)=P@4]PCVJDH\.3&(BeCXLf5<dW\&(FaQ4O]>WdY,QBb294D/87[DJSD
YLS]B]a2ZJ(]PO7L[\<9T6;#V\45=/<.Q,&IY9UNX7Uf:12GA]BCf_[4-e4@U-C=
4/8IYT(UgY,SF?7?U1YQYZ2U(?ab:XCWBD\C&M:C(0738R2?S(F.aAEQ4W5):7A7
MXW9DJXR5cUCVA&Y]TAS<&G1BO7#.QcPCDf2gF2@=7e,;]UQ_T(TMGVag3=61E8K
LXJD[7(;SEDCWX(2.@cYefQ?24H2Z(0?70.@d_:OcKa25cD>>L@1.+_J/_/IXN)g
OY;_fZU.Ye8P3^:C6)[A9F5^dDGFOP@)7?,=PWRKB[=EVKQTRabT]EAP4A\ZWVVR
H\(G<(E+AG1GEKg:aL_:M]DO_>ZZEc/I8eC)O,M<PX@?(FB>VO=480^dNZ?^K)R.
b>8L:OGQ&2b,0S4Q];,+IGgCF0=T<AEE]@9_K&#W#GWQ@Y;(0&+X\8dHV\B:)(80
8A6+)IH][)PCU1);&I?3ba(YBJ:43;3DHC-V]Q3/L-)WS(^]HeF6S6^=RA2<<#2K
VY\8/+)[AO9BM4aR86+,7][WQ4aP57@F3D]661aHFTdZ[M6RIC_?2ceDS_JZC\6#
NT2&<)AB)RQ5SceZ-TJD0LISP_;gU68Tg-0J.?+,8Y27D?N,?>LgZF,4(^d(@7Z2
2U:5CZ(H+\=(;N)&Yd6cL4-2F/#>A#fW-2V:.L3<N[6?=@??,<V.gC:[YX.-EA/;
G/HVLZIQU+FW08Zed>.6c@b#P-,S>-:Xf2/>3O;C,Oc[6>)6E7B@<D>IPN6S0]EN
F\S:YO1(<gB&HJ7Z.L0:3\52QR@^M\URM6Jf;,[&ba.=-6^WRgg,R><(X+Ye)cE7
KAF(#G4N>Y2D&1_&fAV-=G3P<<>7g=[\U@Cdg9gJU891-O&^4>Mf7.dS=L0bJNA@
><N@_:SR)X:1^2[B_[1M6QMWeeHN8_4K[E-JP#5Z5R74<H6&63+L42eFQMV0@-/Z
=FK5<\T6=>.UA0B1&&0Y8\@,:Yba;M]U0S>^Fb/O0d^RdDdIWY]8BeN0DC:O.#&\
L,<JQQA@ULZB(CV=WOBdL>LA2?A236RD-0F]Q[\Qf,?9APb:Q#M,\M6J?(9OVF0E
cM1?FVK>(8MUQO5PCC]?@M_XG1XFO,MSEQH5&OCbF)[/QR;BCC9G>(Xab\,AKdGY
g(+LgI7Md_YW+)\T&VB\dCe>FEJcG<K:0X)82Kd^YKb+/L)[#Jc9R#0U13B?P[b=
K.UCUg]69G]/6R/\4;?21LB<W67,-S6T3&8&:=0R:T/E&@Qb;H9_\GgJGIM]E8EG
S\M:.Db(X0dBdJ:9DQb[DZ<R9D/)f)]_W:CVV9^>Y0B(\[CM)9DR<Yd9\;a&<LYC
>1E#Md9bAL)F;FZCH)Lf,;EX+77JAR0d.&\0((].RBG+gKT8K@-dCaaJUPLPO#Df
LB>eQ0Z(]/\fSYc]J0.X\8=cLXQIGUIc-.g,\Gb]L1K+73c:6/M26cZ?eK;3J_46
<MJETIQX/2eS0W&:L6FW=6<^SCD61K3@]H=G(:JCXK<#;dZg1b?:VeXYR2GACAEg
@=+^(4@[_ScQT->>g\6]8JA.c\J3&B1@c36/H^OR4eDO.:4NfcPY0_Me2ae\[=VE
E(EdNa0G=UQW1Xc=>)YbWJ;_FScL\(K9.45X<c]L2<J,LJHf11/GTZf?+2DQ?+D)
gFKg2G?\HT)TF,;0/eZ\JNCLfJAZCHT+BLU\LDA<[T&?@.Y[/EG&dSd&N)#4S96T
L:V<P4HATf#@1L77D)6K9_cWD@QC[-1fUFC4&TQ#.Cfa_H3]+,S[6C]1U,NX0@TV
E8#cPV_4a+R&S;W5ZfO;DOdDK-GL+H<;?,?fVUc;R6O1eS5J8A=EGa<bR)XMQe#T
&_#f<9Y?)O+c6fb)I0N[WEN,cWB[F@+,Y\SFF7Xd7A=Sf@4)eKU77OX?FIcS@aEb
I(Q[3M2R2M3\5(Y3NM5_4KL:0?d(IDN+)ZS&@<P84[P(,7D31)NCEY0QZ<B.b>f8
[;[9S#_?H6ASVCQ:12+Ud(_W,#I<#SVS[,7W91]7DD_@#88,3bdH^A?8YVRR[bX_
>S3)8S05XI#ZJQ>771cDS0;V_Z.K9Sc.WbX/&.&8(OfeHG]g3GP,JB23BC(1@1b0
EC)CMN=/Q2DFcAEOOQ(Oe7#H:#,TURA]UB[E?PLCeJH<?fU.C14C-H,+c0VRRT#Y
B/d8B]b5]<(=Da<DG0G.H?0S&#4IFH,5DDB)@RC8b.DUCXe&67(bg]A[cG170T]W
,/P0G,;BacI))7Y/KI7J,E.X#GF2=P4TI(JDWR&W;:&IZN.A.FdH\b0#1+,\][\d
&5P6E\9M^K>9CIL3b#\d2IS](L)\/2\:5++0/-R/,_H>fCdTM;M#?XJI_c8XddC1
_eb6]D[[L(OSdZf1NR17B+2L23J4_7#W(O)&eMfEgXb<+\WaDdS[#MNQ+-;\.QGR
G:[BDGKYY5aBQF8P@P.Ub=-&OO7caO\)G#I-_#Uc(08VV1E#+A:b:0<g4;O,ES)1
G,BZ]B7Lb?>ZPe[+1.?_8YUIdS)#8f@/??([\IX9b5CH3E96:0B5@\IEYbI5BS(B
F/<I,A[G+NC>d63/HIX-McC_]DM5MC.G3GSF@Y7>YCE[\I\.=\AZKJAL_DF3YbRd
^TgOT6B<8OJO)A61f2_S82\EG&L&>T9CF>+=@R&3-JJaG]I&SJS>8HXcGXA6BOaL
78U:H//D]d]>DG^\H]2_/EEI3CO.H8BR-7C].A(R?A>5H#d,6/MGc\R,M2:T(-HI
f.a=2)Y,XU0_W.;NR.37JBgDQKVW,L/K-1YLga57ZP;ORE?fD_<c7J<Z@2/0]DQ[
]RN4_C2=ZSUc+2A+9R:GU<60=R^.O_]82Y@aF8DG^\PQ\E43SdG-\0M62Z:e..R[
]SH+bZ#DHPJgP49&2X=)IN1L3)8@gX-_QAX:DcdYA#@UUaeE04,(dSBaGL]\5#,M
2E7PGbI(=<bC]FgBK\I;dE+SJC>X5-;)]QVXWA8Mgf=LKW3)=3cJ#</a#gK1#UU7
ZY1,J1ZA_K.@;?D1JcbQ\F7R,.#>>D0XA=2GEL=#bb+aNA.ER(0IWD4X1fE5ZcG)
^P>U]58]FY/MAU0YPDd/RBUEZSaO@_O8@4]c.=S?cSGOI?D_5(V=15:W:)H]0L#?
C[C^\Zc?<=gYYbAH4Tc8XC&2F77/(<cfY><H:8LA+RA6&K(^:<A>L9G=F,bc9eCZ
TLFX>=BH6VE9&V1?,)C>GOA_56S._R.2FgfgJBZW4F798aIWSTf:VfUC,7)RN4YK
FB;3Da-aBTG:F=RLYeS,G+=42E[8.[e;XX?7\f\2[Q89T51Zc7];5bM#O,,W54#g
,>\1JeYT]If/bd;=YSgL_Q:T(7:YbcbEQK3^/)>,+1^TENN8\-79,5.>0=T=a-0S
OH1D2AQ6D-+DR1d\<>#55#RgZ2gRZDJFTf2EH)EMC_-S/,FAeb1cY90^B>?]>[KI
FZd9Q,K^K-I-U@K+f2PY<:/XdLZN6R27AAIY79B--D[C>G(.#a</1=WYN56,?cG3
864MBb&Z[73,.T#6V(NfR&U[63]AN+UJBCCKT;C,JD9OZgZ+,S8+YM#W=[9-^fZK
c-?V8@fJfV)M<.MD)64;O7U_MV&:1GY\MOM7DSGM_C:QZ<Mg&O#&^=a]Q<4VQ.V-
CVd,?)#:S9>O5.KYHO]H6fP,G7G7)K5-3<X5WTD1/e/N8B=cYG;CQY7-bX?3GXLc
.5;FB[9Z]K8U+AI>Tb/EL+d&6F\94Z0;TeRU]F,c]I^3eF=aW[+e4]d<SY][L?#L
FMZ<KS/4-&HfZ_00T/eb:Yf)\?:CVV6W2:-N4UF6&E&<83DP/(>KSGY[N;DZf\T@
0S.9-L:BdLLQeOKMF3&eL6N?NP@U&@YP>>-E81EI1,e.+[4H</--8,]db1a:P-d>
4ARZV:@]073^F]P@BB^:\Fc=)JG(.Tf-/KR5Pb(V9[)JLUBBL0NE#b<IXf]_NLc,
)K?@,0Nb24bC0IFBT^c[VJE(45T,-,2d53#BI]H7VOEd,g9F3ZU52JLNX?A1+VN(
])KE/eT_13.ZW/SbQ+@IOb&?)9PgVYCN:XI_7?(e(Z4??092DU@J2KLWHTT]5g5N
DP(D[fZ^R<@SO_)-<TT7X#Y=>Z;JZ2dR+2(URB(bJ9^b/.dIB_P?>:BL4^TgHf5N
=XKDP^6M_FKMI(2K;.//c;YCBL@35HIV9+;,KE45c1-;O>CVKJWaF;WDfa5V5E@X
F_M8Bg].b0]\[3)IA&7).LB9=,M0Ra@1W/+F(@^^Icc6U+LO+c3\95Z/JVX@_/FX
0.PM<:#7d<DV4/=6KZS9N(3H6\=f,]cX;>Za#.DXFd96UURTcBX[AZF\:[G??.V3
36Vg(C59XR?FO(1Y@cRbF<J#P.AA=1F7P[YI?]LR_3N:gW_9#ga^f^Q,e?2:RdTZ
4;9CU>g&;\Y5gIYCX6\F??O5/Zg]cRJ,??41^T:X\>BDR9(IG[D^W1NZcbYYe#.&
Z=+Cg(;/_LF\3&H07-MZID0bQFKXTg[E#]\HJCb&U_dg-I@3;dUFFaZU[GJ_)\2N
bBA6LBaEaL=(Yg-:I?dZO^5PgUO?LR\^NI]<9QZ0-PL:J&?-]IT59^f2;>QBU<VV
W/\0V7;OELL&/+R_QT8;)25O\.?RVZbBZM_]e/N;F_NLb5,:V6GJ;Tb0JT&-U051
Y0H&-<4U]^VJ)(3L;aDUCeN:&QC(7&Kd74/QYO/,-P?1<0F2-(^d.c@DIFCDJW,>
E)\5OM,XAJc6f7R)BJF@-Qb=G=4D<3Q_@<bC\e0O6?XgG^=G7-T-M<59E3UOaKNc
L@W8>:TOM#<M&K2T.^1.ZA^<OfQK-SSS4(RZW.=GSG6](f/>CVI0>61X0Z<7PPN<
DB=O]e;,7_\8&;1MK)66:B&#-H5USNeG3>T:SgK9HdZ(fW^AF#;1EL)-T4[SPbV<
3G>92\0H412B^5,IC8Sg3=^8]JaSNWCgNJ8Rf+]Y</_<T=RZ1]3Eg<GVO48N.-XY
7D)#[:Z^9QZ(1\gV##UI;=@Fe9&HZa\5BYY#8/Y>77KJKV)#,W>+UD</KEA=7P\&
ANJZU<WBc3K^=Y[FH_CUF-NG0LBOf<.4Xga99D5LE\-S-R#T48.49Me(>W4S6=RI
S0fI3Jc92?OHgbQR?bf9gV-DbV?-^<LO?d(1Q=D?;W32;4J#[e=Y@QV]Z\.24Z6.
\4A8aQV2Y,RH,D;AB3BH=ANg09^[>4[K<69T]WfIA>6ZJO306/&]W,HK#8XRSHdH
aFJ]G\IV+20@4X=DL+WCb^e1]g6R5G5\G2+R/ff/4)2dZK7Y9^Uf&c;EVd@NE6Z@
R8JdGbJCWFbFN08TI:M6&B3#<D8Ib<.Q6&ES=:FE)g-3S?/H6:UfQJM.:P?+LD^;
^Oe#ZL65G#=A.P]@_.F#6:bP/b=0(,WY/725UPP>I6a(Q<I8EV\Nf,+&R5eMW,W;
^&R#O?P)UKFa315/),QO2=,,Q>c2O.7Fd7<PG2YBQIKTHF7&?Y;dHK.H<QECX@)d
,JE7Q7,OCGWM2?E0Y8E?UNGedM0PF=(.2MK+N)-=+@?7eTP8-CK>L,D<g,fH@a5@
J;(X;2ZM4UT\O+_>,HU:3U,1BMSA6;;^8VBC:GLS^#QI6@)a3EJ+f]5;.VQcU+cS
/d\ER^c1&#Rc;(+/2Gf6V=-E(7Pcd=gZE3+J@:J6I\QUT433__X?BNg_:<]&5<3D
VfTb/->c;C=Y,d^HQcX[-)a\_gPVDSDRK?6DA^:6L6fM+CaX#:LI(7D^dY[9ZHT7
FZQ6MK6;cEZEe)1Q/<]1HPcLBePST;Z_ID(F#L9;NMMF(-0Vd)Gg\Z^)I8?RQ.2#
CDZ+]6H=gTNGg2U7,QYG?\U:K#-d&.SI^0[[AG]KXYA04>Y##4/WZGVc/g5B#9e;
^c>FD7LJEC0&1VcSd<TYHD,H++-+1Zf>.P105Z-?5[YfQM&db?_f/>5YaRD(>\XH
=AIg916ME21bCbY3&-M@gW8D223bG.<b(B1fYA17@O6bC9)XZMY#>I,/HEF1#[W-
IX+8f]ccWdO2(G2[bLVY.-2,;MAfY/&9dge,9cN7&PgU+]Xf.N:+2E[F=511b;KB
X)<Oc-8BH-=>1YbS,B6<W2YVC1RO@QB\)=<G]5=\PBW=0HF7[1_;EY/B\dG<M^1D
J+34BDZK1/bT?:.03\^5,&G2DZ2<5S&MbRUF94_51a24TJ&(OAA,>E,;T0HTd=TH
9[GQ9eSBVD[HT/+@B,7LH<Y&;6>:(?NBN>-5?9+cDLbQ,G4AP8LIT0T#E,G^9=\6
S#:@LQf8KUFOPC79KEFaQVTH;KH1AFQ&YeEVTgH^:>:-3_PV2AE)(gV&6W,)0dSG
\70_9>d6PacWRXW1@f^80R=4MKRKSN^ZHg9QII3RQ-dbXISYB/;.LY-JP[f&C^be
[T>>THF=F:]XL__.T3@S[@W;c67<EEI\]gY^MV)?5M#f0H;1>ZGMGQM^I\Ng3J<>
60O:^Ja)J5K&d>2M_8N8XYgZNF7OW>324=6NP7.J3>4]XE,/2N2YAQFY)VcHBMdF
R_<IYZcaG[PDgA\5NBE..aNVSL#H&I046;MM7HbBFOKG\U&@LHf=F=I^c:9X7)IJ
-G.)(Z3Wb,K4J#9,H&cEf[2NfYD1V0J^@K9BZK.-K_]XC=:+DN56ZEU6g]6)JIPW
^@1+QHLL51IKS12X;QVd:6NUBSdX,5F6:U9LMGcM,8Y]<2A>bU@+_c38]1NeAD/>
JIKQ.0U.C2aY4.BIA4:aJS-8LZ9gaX7[[\caDX\77>#)V^I2YBZ,-b+WYUXeVX/b
:B;EZ5?dG>b#I<g_-P1AJ5XPFH+:#?=^5?6-PWR<TFVT/FAM6D.YL0^P-?2T,67c
@?&0HGBEU/\BJW2d83R[B@&/>(SdWg,D,/(/6EC5+:be=X8c6@H]DX^=DU;COa;F
[80C0VcW)S,E^QB<DY8R#KZB[a?KY4.LF<Z7eS1^708c64#S>Y][DFOdO&;]OW.2
SaL<I3#1X\@IYfD:f#)b\PQG;YaZ+aETKV=T))0)6^,@A&S/cU,1E:H]_>(aM[LD
D9CGKN:dd;.H]:f9]<57F5O8#06Dd=1R7IRJ18MFZ<bJ^<31I2BD=UM4@Qc6b(+7
OI1<(Y-Fee&N>BYgR)Me[KE:Me=M3;+(e\7:(^BgLdf<3\UUL-7g:WK4OLI>D/U7
d#Rc5Kd58?R<G;S>&M9:]S\A3WIRFT_b>YP/7E2A;bP+I:-HbIf-V?@I&L_NG#4c
b\79<_8e)OLbY7UU4g+M]PbCLgEJ+4eO)G&T1]LZTKUUg,S^3US]gf7[>76OZ>?)
0B99K((acf9g66WcR3,9&@LC/Ya1eI8dM#&@&#1E(XF;EJ4UI?a)5g/82P9/JKL=
bCA^[>fcB(P&=g1A)(XKcY8E\C&eI>0P@E>D?6TA2E[4,^K]4bZ7>@ZOH7CLN#4[
.g/J/@W;-d1f^A5)Cb6.QILJ@AFE9@\G[.A^(JB]Y-+cB-FFd)Lg1:e;+dcU6OA0
&.]KYTK33b72UVZM6f[9B>G<2OZN=B)[JLP]3@8POXdagK3].c,fZdf33>gNH1QG
LL?KV,;WA..DL)aXBD(I\ZBE@\c/H_H\a+Q&61;R_BGaU,-H)B&Q[D;(>05+HT,2
e/H=.0@aHKM1Z955;)B+YY2d^S#0gLRfaR3)?(Q:AAOK>(eg5-6[ZG/_GZ75;9+E
5^M\-P+OT]PO#6P(&#K(OeW:gULAaSIXR0^4?]1>\PLg7LO+Q+Qd51gPZN<M1B5B
5YQ=C,1@0?H;Z2cY6K]0c^WB-MJMc+I.&H+0@+(Rc@d:Z)9b06GY=)>,\3IZZ57f
JW53a+J@fDPEVI9E]5bSPI8Vb,QZLM&R-@cIBb8KO#6U#;^#AUg;W3,>fg:>:+6Z
:Z0BX1?+FfB77,,R82SP+1;G(KN-]+Tb_>2c-61K18YKO2<aC&a.4]-PPWBcQMZD
NbAS_W.&LS-;aZQ5+X(?4](7.W<0]794AS&d9JS#>-FefL:/DW-N7:5f+9RG_^O7
[a6e596K>_]:cgQbBJ]1OeW8-f?@J33U;8LXGNGJ?JZfBSLVd[91IOG5U1g?>?VB
POTcS9e1UcICKJPH@C>daU<,JEOVQ<237R+dTQU@TJEQ16.MRN.N_KU><.WMZ/D2
#]OR5KASN\^MbOf>IV=?KcZg\<0?U1^D;GFUW[8Sg9XR)-[(gU]RFA1N#,S^Kd=B
1[S:GbL\[RM(PL.J3]Z<Gc&1-P;#F:cI&KfHfIQ@QF=4;<<.;4G(fV7Te.C;;a5f
FSgCQ3(G.L(^QY/d2Z;2Y#772UCEAYN0dBN0HG[4&)eO:HN+_,K;T_8/bEH@SX];
A)HSXQG,[7DG2g_Y5O3]QUgL.GQQWWS.JWNNHSPGQI_]QM,8=Ub6?TSN>dB3(1<^
_+Y[C0Heg+Sf=5e?E[K-BXEV).]FT3D,&016.\)LF[7PZ@aYe/WO2bcLeS?)_F.d
CWG6+]LU;\5b[)LS2U_YFGH-B9=aIJ[dHRcL]>fa#H,L9E-7,K<c\6b-.V;:1P.7
G]?g[G_SS>4=+g9;+0CSa(3d(f9A8d,08OabV@SV,:^J:E_/YP=DgW>,UK5G:7:P
6g<_0(aO;d0H7OZZ2;]24TeG=X#9P>dYQAO7/IfF9IB6S@LNKF1VL(9+N#??6QTI
34\GB_7>LM0B.)AQc\:e\eBY7c\=1QX@e4VIRXRBV\CQK]32MR?-A1Wb;f3B?(GK
K_<8LAP8;7(gSA,E.Nb&GfS@H78331I1KfBQ0EV9G[-P<D^INIT&?>\E+TZSB[RL
0(#:Xc;N;R7gBC\4HZb(E#M_4bHC_^]U6-FQ,Od?TMbU_@?G1d[@^-b53UFNI;Tg
QgGP>Q[[JK4QE/KdJd)T3\HUS)^=.JO.46<JJK>\?68WK)JD2#-I&R#\TfO27D6a
@L/M9>X8<RF;;bf/_YA0;:AZC<cL4f6=\^aZ8Q#V/._7Y;0>HeLDI4g-35+4NS.]
ce1LaEMH^294(4]6faU[b&SH4\=1<M[BMOR#d(K@J/G9U,P,KN3V8.VIU99;89f1
=L@LOLH[eLL5g(6PFM#HN[Q\H.N];1T5JA\)2aP58f-e_Q8C3],RNf[e+_A,Sd61
5Q/K<Z_#L]3(_A?H[Pe4DHG=Y+\fP[T1S:a.9ZJ&BbP2:^db-[L.:0eD+R?PKa/3
Ub,BBa0A6#=Ne6L#b<RAG\E[>&(MZDgF0bABgX=(2:g08bb1)14/4,V+7V2@<0,;
_I5U?^DXaNN(=,;c14^g/:O[@J9cF70D;71@FC5N&B_O,.8_g)\.]3bO;?Y,>V;H
/;ATP\LNG)@B/AD7#@B?I.ZM/O:&fYRT:U/=O,HH131L>6[7^GH^C8/U,:]2fe37
3Zg]dUJX0Td@/fO568[V@Ie(6TH3;_\T-gCJO.-^;D^)=SUX&S>fQ)+1:H/&FHR&
DI6U^S0Be+()JMDLgNN)\cK_U0QAS.fQUADK<2\64)[,B+/>/N#H[76\c2.YAGSc
2e/UIOYc=DI?[bAMFaGg/58ERUO1>c\MeUIE]>1U?I8B3f(-KA]7fbHP=B_c5ATC
be_ERH@3TG<K9D6&[aDWI&)([ae-BY(XEM_PU0;@b0AYS<8a6\K8EXVR+O^&Bc2X
I&(5fV^QQ9=&Sb)(\c]_4e9HBJ=A0=?c+b)N?c>Md@FE+)cPP;S7O?[JbT4Va83]
1-:cR?eE&WY2QOM;;I.Ua3)=W0>:.\+=GV:4BN<708(Ng]AIAHBa4VMVGZf-=#bG
/P)8YL8?BOABJ&^c[E>JQ?15J/5cQUF37POJ[..O?ZQ;LRaZGadO(1[36A@S:@Q+
f3NI]+b5_NT4X@0>O0VX7SbE4gH6TdGC2W(G4/]ZC?,fLO/P);V&/UFOK#V;2+I?
D5EB=FH2EECB/ee5M>cLK>>]J,=9PP6eUR5AGVUE2_U_G5)Q/FQ@>;L?<+BU-#):
([d+,4U.ZX<\H0X@/I(97Wb)BXZU\M\2CZI#ODLOC?DUec]WKF9b::;O3OU5B@2d
Q/D8McD2dYYEW3>U[JaA\c3bS@L?&LA=A-]]D<#1]-N1[08]/MZ2G6dV,:OX@Id#
O\BK2UU-cRNfR?eW1;b.GJ45WRH9N2E:5Le+/A]4(Y)c[/G>SX>cPfXIYS5Iab<[
4A#/<Kd_G=)AK:)&0SLFY/XSZ6d_Yf[I:CD#_dcgDK^/6N1.QUb]VX;JH49C^X27
7]a^EJ8F_[4\B_FJAe\]D44(FU2:A?292#=-c7.W#1d=/G&FXRa,=)=9<I&O#g68
5@//1d1]^/U2AM?/NYcfI_b(aXb13W?ZY60bbEA6\K9D@0/W5d5O&RZa\CY_BUV[
/R,?d#RgN(#]CMK[75LF++bL,AF^R=W@HCg_XAL#.\7fe,@@4_SeQAd6aFQ_a.b(
?5.^G@7TW<8KD24>CT>5C?G-O^cYI3dJ&XaB6816;<->L>2^.d74R+HHWN^1>9)-
cXLK(0MLN#a/N[e:G<Xbf^@;))e-_7/N2L&?d61/XB/?3I&SGgWQV<=XL1+P&/JI
eS)DS&?EQ,6I<P^A36KR?__([)ZZ7J,N;e106[FC>P-3&@&P#.W>6<6M6<7f;dLd
91:DGAUFTV(LZ@5@e+YNIG6W7=2Y4+<LgTJEbKO3>?)U<+EC4SWPW+L17-XXT_O/
+bWf_(?SQS_#f#>)]_E^[QR9.E^;@N7L)5)OGaFFPH6)c#EK7MJMEHF4K7J]?FFM
W_a^;V@c0TNdIO4L:D>R4(>>][9HU-SP;>]5LgY<NA[8@6QN6N-PHJ+/?(9e4(,B
B#X#=[MP04dAgEd?HJ;\-eGNLMN/<M[.^B.PHYT9^3FNSJ2dIF[L&&.3G>C?FbP^
0_17;2gaIR,(?+7C]WX8SCB3ZC?\E\4XOa:aG@W4c;;88+OVRKP&A;Rd+T#.MBTa
Cb73X9?AgNO#>AM:afDUYGe0@g7N=O0+<,_JfO(,SV=[1ZE>e(FH>&E(YDGR043]
M8_UP<Y_bE2^3&bPg3:U(I[UffFQ2dI/?FV9^c)8DKgc>E6G-f6#DfZUBHI]gFfK
OZ=ON;R--&AGWM>[6)/SV\7@_.LH?/9<DI7XXVM3\(5WV;)G^:9V_E)./]KTWFee
WXS()Z2I&a_2-9M0Y1?g->ZS83D/Ka2-N@6OUG3&O5gH/>X+aQ^f5KM3MO]SQY([
MV4aMQ=&2+@cU9LBf=2DG^-[Y#Pe)#)4\W3TIKU4ebEBB.A8YEAUB+[M0eL^(9U+
d&?c:_NNa2^)^-EN#eIK0)f,#9P@NHXcb?LF2\PcIcH=fMO?S<fX[f@aF@O?bgF+
P<AFW85g]VLKfGXTgHCD,G^HZU,S;b<eO&/O^I61=F>H<R/CLD54Sgac@VG5TIKQ
10-PgV.JeQ^Sb55)0:HKYff845>a=C/HS=>0?d^YX;W2d\DDW7T/f2).-.ReKNW:
AJ0JNXVd,#A772WWb,4_:#;CgF+<LFLRRK@6:AJ8d4JK\VA\W2Cbbg2<<:H+g+X^
+(G@5&G-eG<adOR_GQJSea-2GVa=UG+MQXO;/89ZgTAF?(BVfQ9U9>gWgDb@2SM\
?\X]96E=UMNN0SHZBR(QCKUPP3P6bE9-:NfdG0JC2\JE]>U0_N=V@\a->4UXV>Jd
2KB/D@N(I?)1Z/@.+[OA9JAF&@Q[Vd;527BQRC1:@,3I;0I@_fSN_ZGFRMXV&S1>
ST0TRU=<,PfF5Y(.R(>7&0(HP)2KF+3>g6e(d-.JW0J2V^>dd7TMGC5R\<@Wf-W6
.(6I<cXcN<D.NK7ZL8^#?6S?b1<2#N;F&IV4CK<S[>KS.<)@0[gA26H)QQA<AHP(
gSf72]T-]E(eKTDKOBVKdg9d1AAfBDV0_U&Y0NR[e&.@RO5S[[b^d::&S@\M?g4B
T4X54EdVPTQXOSEP6b\75&a,GVaGC>3:Je6DaKD>?47^>7HEDRE-YWf@fR]>G^bM
f0G\.=APSb>6YZ1#@:+C28J<8WMLFWe3N43a:W>,CY]ZRb:U_BVXT.HO?2Kc0=L\
SbaNJbZ5H[Q-T=&3S9Q&\K4ER[UZAeC7#&OE:LbV]:A2U5))A5&egO4IFFEO(1;]
75aY6MFWVgAG,T:U]acAQ1OMLZI_1dF-N;FM3T#2NPS?>cWJS7d15B].98b?OSR2
Y(Pg=TM]NHf,I@K179QU\TY^[Na5a[=[RJM-BG]Cc2B.Nc4:HU87?R/^?a_B&)UZ
O64?afOZ4PH#ER;<1DLg=.^Pg8/E&ReEOS,a+/W9((W.4=Jg.3f2GFEFLC1(\WC4
CJ.fIEW,O?,KBV>?PM4AGX1Wc;&U8D24b1-KM)b;5I7/fN^7_861OV.T26BPc>Z.
g/5S-d;D2G46)/S:T7NBK2@FLafF>U?#D/I9OA(,BcB.\2DgXL(bGM,IIQ9(/FLK
G+8MGf@<Y#Hbf3T&)@Z2JGB\\d7/)C[3QW.Q/(:TM=KQf/E2]0_L?0NP@aG-M;b,
B>>7@&Kf(+SX[_.B]1D]T0QYL7]cefVdeb(3DX:D1cZfYSK3BE,/U3]J3S-5=7XQ
>aE4K#EKJ#EV8Ng\(;3I5NWI?(b\g_?VH@3(Efg,.@9Z&8KfET(C>QXXQ;(87,D]
Yf(1#T/Eed^>PQZB_cUe@b2I[<g2B;/0b/7A?]O4CW,gJdYVHVaKGL4Caf]A17XS
9NWBeb7_cbO[LB);U@&^>a-=570:QQPDP124AOJb5HgI3C?&81QM?WY;N^:->&^Y
53AKdTJQ,309OVR1f@5KPA6P\0O<1.\g/3XO&Bd001g-Q+R;YA)1[LcT,<45eKL4
5<W-:BW=:U_MG9C@Y-+JG>C&Kc?6bYY^HP036c^VK11Y5>b\S?FgGK.H6[91^B=@
?g62L5bSU]ZX?QJ^\ScUGSU012>0=;Q\@--K@#U(CaQTZ+4;Z(P]5]VSNG([54<2
4?WW+6g=[JDV=&[a1376UcQAc_]ca.OZ_,>DEA.YS\XQSF(A2-Y1Oe9dJT.7fFXT
^2BK6165)N]^U4^ZK2@(Od-<_D&C-RROU.YID^RG6YA5:E>V(KSRSS-a<YZA31?5
YOL6Q[>;e93FP@/)I:&W#5\K\TL,M<IZ(fI;+EaG;;63-)C8M,V:4+^7O?U(CSeS
[B)WZ>^EfJF5_dDJ#FSL0F],4U#JZE1_bDRNZA-B0W55H=a#(E3&[Z.gUdU-9e(d
VB+BWZ^G8KM/&E[(/DGAe2,aI9CbA+9@;[PQ_95-OA81#-QDVPC_8BR-3742PH87
72FSB^6&cW/5.#,?Cc_B6?#JVJOMA>[G\fH?LBQN@-E,#<]AS2H(dZSR^K:X4D3Y
e#=47caQ=a>VbYHE=6^GMME</&/f3K4.d_P\f?0#SU1:KKI-9C+:b2TIeX)1(Y#F
5^A&Z-f49(W8ZLFLQaIUX0G#O]29=&6L4DO6LJe8\W8KHfKZ-6HZ&ID#1LMdf=JX
)@_E=,3QUV)K(V;cS.X_H(UdQb.,^?B.2I>_TEO9S\6feMaQd4V[,JISMd^)>.?a
M;Y474U\0cEYYTc<PT<G=J/La#,B&P&eC,#MNFHD;3MMAacRUVT,05J9V^>WOL4f
Q9T7QJQ7@\7)S3@_=\G+TdS_HHTKV_-W>6XacKK(Kf[F#c_WM+FI7LJa>P.Re<]1
Y^MdOcX]6FNCGa_<7-D+C?:b3AgCVafMSRQ@>aKDKP9[G0f@5A&-IMN8G]a)>3Yb
KJ1a(ba,OAI1/Se>BKT[7B]NT_?T?/,a5N-;19VZF<b+A:+gJE5CP8#2U+N0[7Z@
2S,T9TeQ4O28K4B:8K:E+8FKL7ACNbI7A<c;2U6U+G6&M1A,S>J/_G;BHBggHIBX
DcM<#aUD7C3,/\L_C;05G0H5RW#a[)-eZ)YD?H8@FD,Uf/):EV0YS-YT+.D3NM_G
?d7Z>HNS,28Y?:ZW0?;WIbY:62K5GfR7U7MD\L+]MT16dFLIb^72(;LQ<-LJU^[>
PAe3^GW,X4O9\Ha/[[XD7_Fc?532c:NSc_:(/D1X#S:1##GeBMY/QS/C;PGbQKJ^
YY3e\/e)dVfc^,N(5I.-fE^?PGZb95#B89>,edHcb/@a@QHBISG=DAZF\?72a;ZM
+]BGWb1</V>7b)Ac30@3)WEdV@9PMMU=B2+OEAP\B2>E=\(e00XY]ODKGd>.J9cg
)HNVYYX#+H.&C8:#;O&TSB3JUK:Ug91G8YJ?P:0Ja_]7AQA78SeSN(-8bb/cbZ)&
HQYM,DeBT1XVD1A=P=U:F5@4T>g-eFR@X672T9E=+ON3Sc8JUY3#(;Dd+\8W#;_K
^dWSW7KGQI?e/C=KcTN_:]M27+Y6RNNHQ4T(cNL9YG3(;[>V76Rd8H[^4I)egdX\
1aK@#DT&D?-(3C1AUPN@dJ59\RGb)=7d9&UK_Ub.79:Y@TTXUd1e2R&KeR1O2MId
</Pf3Bc8@OgU?9_8;8+95d;NZ&NU:-cC@(PHg+b5R;B?/(:1XggPBHaW3Z,].<X&
+/#/44GHLS;>J5HZ0)3.Ve\F;7FE-UASb3BSY+753\):KcR:YF#S1BMY#<;COJ_.
&+a]4UB6QA7==F,PGCU89JGBWY?82:M(>H]9;UNb[&J8eMV&c4(,7QQ^J^]B31V8
W>d_\c)aS/bWQE1b_]47]PHD@4L6,ZP9551a4UJX+G>U^?a0b16<gGRL+^M;&RW_
W9?/2R4(HDQbIdfdQJ&4gMPI/]A(9QE^)BD]AT(Xc6Q^]5<:_SdMfeKP:T>E:26O
JHad0DN;W>DVESW_:7YG(\=AJHE+dA1:CQJ7eJNU+4f>Lg=C3+4UDGabd@dGWD-a
C08-a5fL2&)(6U_0GF7D<=74;.>Se,Vd/-L15OX;^:)=+]U\=JC13UT:-<5N]4+d
+1F=@gWNTPeT]Q/AM[Y+?cUUOdO5\M9UGc^+?@1:I3YVW1_[BVe0bEB077K.NELK
:]ccXU<9&<LSEBS:(g)K[U316/a<&^[f2VH];7>3Ue_).VEFPc:/3>NF/1e&I6HT
K>0(X]01QDX#a8bVgfT&QNP4,-T7S,UVc?X(;N?e;X<&WC^(.U/7:#ESGR)H_4b7
8EaW<+>gf_\#@3=Qc30K:D5C#-WZ4@Y=L&d#M@e-,>Mb41#Y@_=IcHHeA.RF-Q_a
_U@;?1H&WI#B6UOTHN^,D+W.Y6\c54X^IMHPEGbVJ<.6KM-OX0C,5S37A_FA/f#K
)B/+Z(<Q6SUfFJ6\\DXJ##LZ;A-Y]e&O(10,#8f8HPE&:fYVPE(@K-Y;d/UU1QQ.
:(LfA[fVGM@gge5Vf>/bTL#WRLdXU^)dgJ-QeQP44BRNVL<.Q>SU&/;Y;[/eHaO.
3@8CX[D(ACA;6/&BU?eMM;2L\SCVR&5]A83[:-/#.J_1\NC,gaPP+J@S22^F&(7<
PG0[RGJ;ULN8+Jcgf)-OWRZ[]/.@X=Z2TS8&(GbH_D4-PgZ)VOIL1B>+B=44^=dT
WE7cHPMHa<bSa;_g7^@S7L(/8[.N:ggH51:=Jg6FP7SZY]Id(I]N_H.#1FO@T(K?
gSUI.3B9X#XT2gICHgW\JfE@M_?OB:\9Qd&;#LPZL_d:]USG?>UIG^.5]QPIXLJ7
\>>d3QZd[-K^R,<KP\@1Yb3</.DbIOFNGALG+>gA.V>H6;1/_)?./B<)TP7\7UW\
aC^B-<#ZOabK1Q3\74GZ<0&-AOA+W6?dCNW_:/A,LM&ZbUE\H7M;X\B^]#FNH_K0
]\)Y\1DK&:-d8gWNQA>OSFCSG6;bJ^&(d>K:&_^(=84#A-4YTB/_?Lb7b,-/@JG3
,5U+U?CYD<)=MLV9I?[e85BNb,^X;CP=.ge@#9@C&36_9:(ZD4SeC3b@,Wf3_/(L
6dNKTDNc^>T<?(Zb/DP.V>CZ8>N9EScE3X#<e7WJgHC^P.B)\c;Sa:/_U<J31MYP
Q?UOF6)fJKCK=>TP==Z;=Q[:5,CJK=I1-M-dOd)9+g3T)W]_QK^>8<V_:cM9A@MV
QMB,<I][^a<,A\TD216D(OJ5F06#5KdEH<>0M(OFX9,UPU#B.b=H8T^VFOU_.1g9
fHPY+48KH)2DN1N6a:\.#TH;,cYES^#,cd;Y(S]aF]6RI_#cRCa@BgX-<-O7CH70
SEH3A./Hg>6;#/CUK<I=OfF]D.g=/4eL3eCPa5;JLX_NU>OgaFZ#DEXMVUWJ,DTg
K,MeU@FEY#TA)L&YWaRMG^6[Z14f4LV#K;L5EZa;5;P;WU^ABJ^N=20aZ?-3.)cG
O4?bM5B6#KCAF8X<(g:.BK5MZZaO3FgXNR.8NDAJ;#O@7<-TFg6G1-;?DUJ5#+_=
,M4[]:=/Z@SF2BL[P]9=B)2RW^:L=_+0HD9\(NRV(XI;Nec/TNT<5U(]?dHLS8AX
cH.21d:1X6Ub+]RS)-#:0L#GL[0CP&KBOW(]^+PbcMB@BC:<#ARTD_]2X8FER.OS
KA_:/I;3NFE)\8>b+C<MS.-]I>?^O3]2HR/Ug2VW:K+8Y58faR<0P414ME)@>O#<
V,\G:\28+_D:Q(E4#P&b?K@JM##IF8D+L-^9.P.[ZF09M^@PRN7>CCD#69MKXE=0
I)7Hf,9X.LW-P;VPcC1-ASfUF0Ub)9\5O1T9X@FF&fd=Udf5+dWE=]-8.<d-f&94
J)HH(=>61UCQ_aPP?V(;[Z#@S3HBAE>,TG6Q1S,C><U:WV7GJXL[,G#JL6BE.KQD
.NPT])JN8W-2V93IQM+9(XHXG_?3-?Y[TW#P#d3BTRVJPYC^&B(;II?aFFC^W3H2
SA/T)]>+AB)fT:F@/-H_5dWb>CV+=4B_-,X&:1R:23YQV=K7T-@#c]FF58D@[VY@
0:IN_Q[D__3>-.>G(>)8G]f2\>=AR4XT:13;c<1K:35YJX\,L6/G2_KKYM6S<8C8
0d@dZ=\,B+JDY,]CIZccbJ\ET9Z26]43S1(7/,A/9.J]_L?@-><XFE?\].ad\\?E
9/,33546c.G9^K/fQf&_f454L0D-?[KIR?HA+6cI2VQGIY.N^M^J-]bN,&?S.LUR
2.U:,\E/>)c#6e_e,FZ_8:G\-PIH4M)J/XXOT\;;2)@65g&2UZO,bcM\<d;OP6Ba
FOc[HfAb/BA?,5\>LgP>ccd7)PVAL[/a^Z@bZg;X5c><;;:G8fcDBQ&X^:UH(Ag+
)=aJKTg8/NM1=S/3;Ddb)fbA&W^JL.)aCZ[3aFVU#@B.\2@1bbWPd:I0T8RG>B,H
=Y=e1S)2P,eD3XZ@^89@:=D_7I)PKLF-dV?L:D9S\&J0N#XR=4M&aB:B26aSQJ>a
(dSNB&a&f=fDGE]#?Bgf)<&D&K@>_5L<65[>.0F/V(A54gBF9Ab8_/edUL\SdZ)T
WW>TffNJ9(?J;BOD#P+Y3gU@KZ(]HZD+DOVK+g>-M5P1+TecR=Qc346-R>&Y)Tc\
e3@Y?->3KcfIY?IP82bQA09/=G:g,SWJ<ODOcXPEI611gBfW,#D3/GX6.V#RZ5,K
fIQe9NGRGI-AR83+6RXLD<PRX11?M3XS(ECbJ9Ff]5HSETY<9-&4&SW5C\H+GEcd
#b00F^FDH#\e-BE56;TWQ>+I]@3gR<O.:I^b+O_3NWFUP.QNgK8L@gf^^ef7OeDf
G56)9LM0E=Q11b4AIbe,P@L6g#GC1>b3AE@#4IC=O:5TWA9KfJccPdcEFDJ5F@M+
=c7cFf:P+0Mb]=:c/APB:6]+D6KgGUQ#)KFBeFFNFQRUVdLV#?V:e&J,TAQdZHO]
RQ&FV;-LHc)A3ZN[5edN;KYH1V#K#\-W]E:f9dTMMD:;Y#STfBW,?X,S7QBb._UH
IQNJ6S-3743g1JFFXb7:J^5,/9A6CYM(JgGX\<FI=[^Z#>^)gVTK@X](3[EfS&[_
bN/KCdGgM_](M5FWX7GcNYL6481?0V42<PeaZ)^8#-Z05GH:]T1AE<)+d&@BD1=-
]^41S5Kg]ZE9X^?G49J-4/eIb^1\F,5Z<U#BPf<g??2@,6TO.U(.:<53OFc=2^NR
b_5@#>WYQY:V-;2;C0XHW#0FbdBEC:D4dOY\^6:-AaFJ^f\b\CXa;g^)[&8MTW&f
W4]Y;G&FOEFL>?C4M5Og03[]VECN3FMd63bY^=>_8#=([JDfG.4df:V:?09g^bdd
C4(SI0H]8aOgYWg-:=KeADR;7eIKT<N@g^_eb[f3]@gVM5.H6=G=O@K[CL/4YeS+
5=\Fa2g&GE(-AVH]J=(3H1SeDSFYTOOc^2=1+@T.QO=#WKa>5Q&W<:A@S6OG54:L
[<,XUWd8g3VP<=^G<NRY3SBT64&]DYCAKTeZSZ&B^MD)#0JZ++968Y6>e8gRRb=T
U?X#>[YR]C,)XGQ0^BF23H^IM;B1PU;H^#2/XY>G2,1JI2M#.@g8;gO?LN?.eeRR
-6O7(60DMa#9&H&/;L1&?&3CJAEZD>?C1O0K(+N=NX3(#_@eDfQ5^NRd+EVb1(:c
4a1CJ2)G)VL/MXP.4ca47Ve8S@c1_KK3-E=3B2&:JHDOL^UJgNW^M.W8:PBKZ>:]
L,-69b+YU6eMHDC]dT#_5Ce#LM&_HQG\=-[-3#AQO+UIa(2,e5SYb+<QH_K:=WBQ
U2Td+O1UaPL.T_7BeF]QT8H/A0VY=XQ,5B>\6M#<CY(7ba2TY>KM^+(eUWQ\1cTS
.N5G];QEWIH_A&dZ;9WS[T0e4&a-8\8P-gI;+Q_9b>GWcJ+VR03YdV2PETB)XP1+
PN?B;dFaLG[B_EdC]6@1&5[&<e4Ee5Y+aHUP)H-,ZN-EC7D+^/9@6WePFZ;56g_>
fED7\c_MKbY6C>AXI8U8)d7:(3LH8];MOFOEDFEK\@ELOBefOL^;=D&LJ+9DQaC_
Ee7]=TARE1P)Q;8O[PHEKBUfA&#W+3E4KH-#R5/?7?/=fYReH8#]LOZ/(;FICPU1
;F=M\7BYC)=@0X8RL5R#fW7dSa6+:E8Y(F2KJ;aS6LQ2Rb.WS5X<#/P9E-),Xb4_
0g\d.50/K_ZC&dX&Na#>;b]>14S73Z\,05E1@63Z=?)]D,95.:TP=dJQ_#L=Hc0&
4UHX^85L0\\f&P]ZPf?HC)]d<<[,]V1S2E\dHVH)I@:NGf/O__IE.G<<U+U3M^&M
5_Zg&0,JgCg8=FI7\cV&OUb^LXI/,38(@IMTI0\e.\NeS.B@a8LB+)C/\3NHH-FO
/6=EC/:e+1>F)Vc[S&&W8W+4R>[G=NA)14]a5e6-c20]+c0]3aZ3M[aV<?<T#N3E
>.+>J#6)[5^aGUH]R8II/T,2YI.T5=67E4g]<,Je<Tf9Wa:(<,3=TDJ;9f:(cK:R
7:((P0XY7&#0O&X1+@Ibb9&4d:KI1QABQTXa<[K4/=K&VI2\b&ZfIObN>H>&15R5
7]PACd&98]S[,EUY_1dOD@F<bYb#OgdDWaP<]5\Q5.@EE]OQGKT4K;dPV8;3g8X^
E9b-+;a<Y40e>_NB(5UJULKeH:dW@.5]AG/@cZ\&.gL#[+5bEDBOfHHf#,(ID]&/
b>H5<F^FGdF),SXZF=FZWQ5@dYV,I=[&PSF4-T76N=7\EM=))USP^A<6YRF=^Z7/
XZPa4Z=WY@KgYX+I(^c;T<\1dTFKD.62>D0UaJ>[C]MX603\T+\?O^[4E3bC5e9P
a-E7#J3b#CC>7)a(Q)7ON6I7QIfcN:UeZ;Rd^#UD0XP\I00QOU)WMGI;1(3.g-D?
5N<XQY4gRR[8WT[]T-GcgdOZG=Z[2U9PMg-:;?]0RE\U,_^_+]U8/Zf?g.(YeYO\
HBIRT&T\1(S.gRE>bC0\_Qg/Q8+Hg:[7YOW&P+@=X2^=)(_Abd13\3eBY2#e:Q=N
:<66gM1;1\SVg929[\7>NdYR1^,TWRMW9\dR?PJ^S^JN31EJ7d@B;a>]C0+;HG#9
@75B5)_BWE<Jg=9:4W0WDZ2;^cNJLdQJ,VZ->,WS7R__&R&Be;Z=C=@cdY97a^F4
OHAeQc.HcQ_ONVE=R@;Qd,=@(Bf&FaZZOW5:87/_fPLGDE,EM:+McTCL09B/7NFD
Tag7;=1W\LW.U_e/P+_/^BC1I=]OL54[@XW(>E49[=T8PCYFXM>gZ.b?TPTDcN<&
VfCS33<W,H.b+YE\Q95IT#ST(N#fVHc\Q)H_K&?VM@a0_(b@)1(?<cK_PGHF6:-6
?UGZ378BSe5G)W.0+X66[3EGKP45I>BQGF#A.+SX3/HcO4_@#F7J>8T5bU-_RTJ8
U[bGWIb&QO6;(a>[:^(9GgOK8)X<dZH>EYWbf<4G(U6U3cU[ELKcbJTW2f&<P>#T
YL4,_>UP-A/Fg)O1@BD6;\&Z\Z5S]f0<46ReZ7?;JB##GPfO4WKJ/B73LKc:YAgg
-<8ZPb<7]UfC7&;116O.Q-Z?R/g4O@N.Z[G_dgM<E>FYY)S^O?Y]]LLY+1.UMJ0O
eP6FO2V=^P?>^?Q4c,CYe5-17Y1(_LRBK.(46A6,1BUC?AAN-eRKfDZ?N9\(@aDN
WCNa=E7[0\#@4Na<++Na4KXI/e0>-OS5VD/7Sb\)OH\M>6;D#O+^0O\A_1#b&>0:
gH7bTXI<5AY&]Y+&E(4/+@2dJA:<Y4GW#&f(<A+Z7WGEK9SK57eP<=fQ^@fWIf,V
:OL4SZIP1dIc.c+6++7+G3cER&-,>g>e@.WZE0&@bLH,IUC.VL4FL1Z_QFNH8a@6
F?O6?(cW&LgfN6&.^A-9IPHMLcRfXQV>=eACJ[5+M>:Ueg_Z5Z>KB+6H26[90K8\
=:5VaR4QI#2g77P?>:gJRYD1ZE81+0aAP4HF>NX]3^<UeNK#ZIK>^>8GY]NeFW]M
YBM0)5GSgbGLQ-dc?NP@gaL+]0_gY:eFc(PV(7E9eY0SSQJ]H&Ng.a_F66f)GKDP
:MCRKTbf+gDLOfR@_J5J]<Acf<C;L]aX>TJ(1E-/a5E+4d;E1BA7VMDY/A(3&?T4
,?\C>T&F:Z9cR56^;#c&]N[]A&5F=4?AUU5>f@\GTM1aX&[RSX44]G,]A/5DDacJ
6]0DbZUSZHC5V::XRdR7K-&gdKTKTLP;Y+TGGAG.OQ/P;?9+c=TDF7(@:b#Jde.^
-;EUFM3/29a_V>&HR7-=+HKI:&(@D?e;O[fT1+d#@]8R&\CS[P6ER+G,B6WJN@,)
\Xa>B0-gbMGH0RLX(E9bCdA;ZE_gH^9N;A:XVLGac&a[V0+_Ye8QM_/X,.5,#4I2
S^FA;P(g&GV6[\/]WH@JZNB1KV(,W^=O\Ne?cV&WM0B17-,+\ea.D]Ycd6da0[>7
SI<Ab^V\YH4?=IHY=aM>Q=0a0@e-F9CA[X@TH]#2e^N2?W,ZL[J]5Q5P_-(fG;BS
2FU0B.P3+1fX.YV85c=T>[Y)X(E[8)Qg;FC-8,#I)B>K-XQ0UH[e9183?9b-SV^2
cK4)_Pe]T,127Mb2VCMgc:M\C.7^()gV=<:LYFAMY9L7\(^CAB\2B/4DSO.R@.2Y
\fWC0I=\>>\LX3_A(VK:eFYa92SNE-g@>1^cP92/&I[)O+3RP>55XeTCIX=Gd]3+
CEB4UW=EA0cFUBMcTf(WI#9UQ\aV=[R+@(\Q-2XNN;5^AS?.[-NMN^+4O-e>(B[[
9_N@OfB,-_D@/7S@VY3Y6/^M+B9NZdND,-02g]IIRXdcS6DPIaZR5La<gZMS&aN#
G::VUGOA7?b944\Ya/2fUSBQ^&2a+O,g>OfU:M_WK:J@&MG+Y,B.D7I]2^Y\KE.0
gN(S(:+C?D\5W^1^[:Jd<6W_<W2GZ1bRXDC/,UOaaHIeI=JQBED(VGLU=^_aF-eJ
eC\3GUZ>PP[[CCA=GTM&eC9TN2^)SZ_4fcaZ1,fU.B,.#gc@5E_:efWH]E0FWZ0H
WS:)a<-\XXgQLe]=(SJ=&CZd6L:KV>F2#89JMR<P^@.@I+Pf<<TV^IcYN_?<DYd^
NgRH91PW1I0FXDA/Z6SFV<a,=c\N9<U,?_B/I5(?FBO2g&OPJ+47-f7abUYQ=<?f
@b5[?Q2@AM+<L4J+^,=>5M)aX]^3,e>_Q)LCFf(a[OfM]MKBM3XX(<,O](HP2D/E
DI\ZL.R4QSJBHB=J<;[OJ).GQGDD198Q/842fK>bK49NOa;(\UO](R4UH/eXZT(^
W[c:UdQBT@69gF1ME0Q/3eHb84gK#D_]68T:KJK@?-J=:XPCSA=N[4Y6:8=;a>#e
ZKF_25.Y@6g9V9Qe?\(:J[FKUdEQS>,G2-BaM,7-,?bXAAf)D2(GMT#f]<]f1P8A
+dN8QXNH7M0[RHE)Z.J/(KZOH&IP8R+(JM_A+TGBEFd4@,Q>59@G:VOe?dgSOT_V
5e,fgZ4SH,?b&]A4\,:,.e-[>,,UA=#gG?3eL2SU33L@A9X9cT,F+0,Nc5[??BEX
30a(,ZFg2_<IKVLJUEHT>GB9#KR\DV86/1:E2):8aLXeO97]GYE6?TIND0@eJ&B/
A5\TPa[:FLPY_K3b;=H:B_&-,6[MYb5E-Uf4,^BU7&Y\Y5fUBG,^ZYOWHOQS+9^X
)Qfd+-g5c,KUV9BW:66U9#1-dB_=P]K<_]8X__:T/-#c-N;b7/+f3A/X6dQRb@-_
BMB2Bd\\0X:KXgeAf+?EHLUd25-6E2#;J_OfRfW\\eRS>N(;DZeKN=>FL]EWT62_
#,9Q+\WN+DH&_<f\Mbd[H2VGg1^94)/[7#:geV7gdZ0HHLK/fWWI-R=X<@HB#6(<
A+]gSgMcO5IT_R,#N(\CA-LcK&.D9,IY7OfE(K^@_TR[gZbEEL7:>M(7He(;98XN
e@SQ4=PMVee>##?K(I1++_C2=3OdX9f.A41G9YAR\1OVad&NG-S_dN7[59_W1(M]
dF9IMSJK?+4W[/;bK]Sa&L6I[3^7PG6PHeIQKY_O[?8a&U(Jc]M5F4KZQ:/ZM&AQ
_a:>2Ka77_2,@\d+ef]T-0HdfT7]C/8](4>TNI_+LdgBUXM_e?PCPVXd#?^=0>Q=
ZOc.^.38JFWK9&/1>5ObbQL;Bf6C?@1fJbFEaV,C9]\:&+F-5]>)eC@#56>92HFH
b670</3gZcABbW?6+K[MV\&d;e2)_BY696I1Ad_3T==:g4<e-Md9Z=A.UO.CbTBZ
J=,eOP<K_0X#31JX3HWP-T<1g@:#)>-E4CA-WN(f_[#B:SKKUW<ASgYHRTX3c1Hb
,=:5MO[Pd+YR;CV)N4<=4@[/]I^C&4fK+Y/?C,X+AGX@-D/M9fR+IM_b\0&]g8b7
LZGg#3a\HR/E@HB0/fH+E/+?1]^;V6E;0CL[F;4daYgPY\AVR<\+_Y<bR.)YCYQ3
>=B229#Q./b/&b6L7]a>cQVY2fM/#1(U&VTGJe\\+d[b-TCXUA,,R]3AfMBI#c0&
e]+G@,\/;f<We1P=/F#E=S]^PTP9B.15Jd&KGKFG7@,&DR6#S+(c199.)WRP;ffD
9Z,^BGBcT^0K5N8gPB,babH+8Le;W[g7]Y,bK^5/H_bR1WT8OcA(LE,8B4I/Te7<
ZS+)H1AYN2M6U;X_-[Z#2<N01c0LQcJ_JQET8)CCUecT?N51O.[870N+<dLO?KB\
3)3/QR.O(,UE?3VKb:4)/KBbHQO3ST\WBE3/9;5&BR;-PGFT&27>F+CF(WUg]P+B
URVgN6Xa#f--;\+?2(_C?.d_DJNa_>4O:,#,JC9\d:F>NHcM6@/9,2b]fZH])M#6
BA)d9V5U#0@c1)T53W5f/U0DZaJ.;,b#X+[T7A:@fGT^T(JD.X^P+cBZR15[U9\P
G=4.O#7^REG_\@cAF3M<[+7e)H;]M\:V6+^[8^/H@8N(=fLAdQW816>?]>7;7#0Z
?TLF2/2c8]KEO+/NBFQ5NY[L/EET^)I,JH-U,NaWQ:/PFX)YH>X3T7cG=2bA67XD
2K29]Ic6cYCNdLDWb?D?FM:#,bHc&gYV4P21,1U#Z1fITT^d&^ELcd5:GWYd\JSU
,&=;f3K,TO\dEHECTb6Oe:f=7-/XMe]a6a4)X,IJgR<T]FO>=U,LV]/=EY3QaKH-
.Q^\/>Q2dJ9S&](V/@^>P[><03eR1FB-);+@L9PF02:JPP[N^81PPDPQeB7MA7+A
YN+7Mg:-J/-C]CTI=eE>U9MdZ+AAPA;9a<-gc]Oe.)>UBAMCM0I?E71Id_.(#R<:
]DLgB2TZL7[a9_C?2[HNU@4&B7_:>Q.aMIJW27WRZL6>:fYe[+ANc6>PCd/F,V)8
d&UZ7^P^5];/?fC,_B/;b6f]C@JOGE&65=5B3.Y8:WfBK.\f,_&;BP#5f_a>5fY#
45<3<geFQPD8:CJdCH+eTAeA9+I:f:T8+V857GdB5L.IbgA7Y>WQLeT/9f[D3cPK
LKDW/@)aGaV[1]+DOd0VH5DV8NWeX=)W9PV?6->#:Yc<I+MQHa.9&I/DfLH0Qd3g
fG:+^MfY]]A\:WL66[Lc#D1a<OF+JRM#FL^Y^&@S8#MS2CA7=.6E2e7;?0XdKD\H
G7-Eg<K+3W[MY)S.dINF4/@/g#XbRX0O&L2WY\3;=]HD2B+G]>Q(_L<<@,G.LXFN
4d5M)SNK;KB:9YZJb5I[\WW\bg\=B+01eNH1f))J[+bY)A\>YWd>dQ+T0XHea)L>
WM5W\N_4/J3:KJFHXTH(S7Q&\[?Fg\MI);f#cJRg,FGRQ?H0)0J_[3]V^YAa0+59
fQ2f237bebDYYOdc3dfGZQDKF()V(-Sf48[S1;);cX8c.X9M3X3b_=/LS@B[AM@^
P=\_VBRfC<bXLe[3[9&ZfQVe:KXPXa@0F2#>V]V;/-Yd>YYY7_TB\YVE^JeZW/R9
F]Y3LN817J9Z<IC.FNDSW]d,0@V/dL:E_W538[@P(R9,-=1cE1b;)7,>K(g9<[-\
-QPMfca0H)P#2bOHO5/OG]AY?YOH_431F#W_HA<&LR6;5N-OULMRUB]#Y7]Ne668
0abL399@cJ4;;aNf939-[5<(V@,MZSCM#\Dg?#4d]NPG[O_R?KK2S](R57Y,FKc?
fcL)9QE&bA4eYVg3Ie<T?#>PX6]Q16LF>If^UU5SKd/-^KEP8CGUGBSS2#U<PR4Y
W(EGS:GZH[&6[?]GK1a4Y6[DD3/L\,c0E]PBdSH:@d541JWb?,WP<Y7(WC3I.)&&
#UXB2K1AVOS7EET4DJ^#B1A(M+F7aD5I3Y,ZT[1(VQQ&F?227A7A7=GBd(:Z->0f
f)b-+4EIH63K<9))=NU0TP+?9@-;f7,b#9.OPIVQMN8I2U#0gLWTF0f,081B2HfQ
3NR+B5R[Mb,a&(??SO/e@X#UJ1-89069P2U)7-dO+YO44a]b(^0OVTLJZSPYf_+0
W5L-PX[5JW5[(WaO8R[6.P(/0N:CZccS/M<fA7M@:;Z:GcEZYH9AEf@O6+\UPBcc
f9Z6b0(F1,O<2+b<3fCQN6<bgN=5(6L4@)(HNZ9+WBPXf?cYRG6/+5.3:\UGLFC4
0P(71f67<V#R6D^dV4W5HT)1O3=B7,FTYc-,5_-T\G7(?X5PZJde0_?S)_UP4(b5
,\&KZd@f[IN<?TMCfPXYZI_P=b^-1ZccDe4SK-8#\QTGDW#VZB;R-GTDR=\+DRFN
X\B>ZfbcY#7Qd:]-TQGULU7CEf?La6FTZMgRPD4c422,>(M1a;6?UE[P#U8X52LH
-+>;9SJZ13)^agWZT5.?T]VWZV870.Qc;&&Te(PW,=2.T9U?FEFC5e=fX<()5)6I
87g?2=LHM\Wf4afa(V+=,XW0W,gU19T+Sg(YMQY+>.<NYgQHK5,2?@U=([0eU)-.
W2GP,C15Rb8LJd;2aS[<aX9^e67AdRXF8F2X6T+.FL=8V5:A1aJE5#]8A;ac,RII
gTIW>bF;OBIWAYXAO([YEBdUNZ,E(F-HNR:NeFQ)5g12>^Y:XYM#A7O5T>X]&Z0S
K#5JP^(UE3A=][BD+L,Ued<VFLX1QIKf_f6/6K:E<#S1NM@UWTPE<cN/.IbTI([8
X[92?e,IeT,5g&RONb[2HQO6Dac#.+)/=#K,R2,S:-2#C(]7<1Se_MBD-IXU>fPR
Z@DF48:.0e8FaP#bF31O8eSfV^]P11M24Kac8.S3aZ#>V6]Lc^;Ua-Lbd^]?;4DP
@_@FHLRZgEf]B/7F#+gTA-BK?gMM>6[XU#TYG(,>[LT2Z;49ba([70-Ea@e:c3Xd
7^HN9HIbW/M5V\?&GKAB(N-Lc9gI.?f6(eKD,W+(Ofd@dHa[R>b?6\]eR?UV@.b:
]XG6T6BK1E-7+<O:O>XKQITL4)XJL6]1\A)9f74gFgf+6dLJ1QKQEO;X6;M0+WX>
Xc[C(+[c2GZMB[YM].T@QMHX+3OBW3g+V,\[@g:<+HXb(U3#,^4R@=]E3W,JG#D<
H\f+(TA_9MB<.@cTE[Qac;CZgU737?//GZ]aLOJI=[a96AeO@-6FP6A=Ac2C>Pg;
Fbf88T:+,;_@.CV+CILgA<:)OMN3KSc^3U[(R.VFW90YW0#Lb&_0aO)/[a6,YI0b
?3=(SXKcfWM_=JQEACebT9S-QIWdQXU0^@;Dg^/^cPKbR;,FBP^YKYXR2a(B5FTb
gXGX>>\N.#@AeJa@b5b8K=0FTJdd@8^S[.._6;>87T@DI^^3;)?5?<59&_3YHH/d
Cc.I\+U9gfA3QEH-Vg@O\U=Z[?777/&;&4a.&EV6_38U0VFEf6E(VHIF/>T)BV@?
eF5PR3e^RH(7A@?)Wg_)7PJK&=dNN4OG_,&e8:?AABa],RXcE-(5g#3_^J[#V26<
A/bXTNb?Q^??_4&A=42\P9c:N8Xe,NLeA::X.Q4eaZJ>?<5<Qc[Q631RK?4(bTd^
1f6)-;b,ET?/6c-8c-,U9\^8f.J3cQ>bF:]?>O8=8cV\TEL2H=MN7=69UE]N:Ie/
a08YbbRV+P3]2\5aO6XA?Z7d>a[97N\8=K^#d<_Te,17P>;79?9WR&YDVO<7B0EI
AGJcKG:?9J3E]5C,C#/MO(bU08K6_bS5YA0.Y>UN-5\3)bF(16(<4;;A:^L6^1Z,
=VF]JcY=&d>AMR.2LQ;>]>X+K:;A&UWA9cK;Re1]/;;14DfaDfcV_<5,+:ZC2?5#
=1Ja0Z1=6,E1S&ID(+&OY6#Sc,TEE3,_,cWC5c4Xd3UEOcHV?L+e@O2K&+/(SceM
fV1_9KU9Y2RWITMO/#/=d(M?/525NFD6A<BM\LPO?75?31dc#\/J0\B&-5bZNDTZ
f/()/_U(#+HSUPIK;D@164):O[ZN;.1:dV7@feWZ0;3[ST:\\.R^Q]P9&BU<A\EC
bUYfB);CbJ+f;eG4NDBHCR,^a[D8W_e8ePW7/WWU8MM>LXN:BE_;)d_-J7g>,=f&
e,f;:H9MKD5^U5GX06Z2N#12/g)<1Bb&?)E[-@J_U+\LHNEQ(ca;gHFGK8Sa4;]f
HO/@J#/_>XfY2:\AU#IFScZWA76S(9(HEBYK8#;F9RPb6\QU:K1T]7N5N3cSE@Oa
N8A&8=Yd&KMc3?_@)/;LEB7E0=SB(eb??&/YCIW.4;)dH_a.YeDTS,)C+B#KO3:^
X7:&Q.D0\:FV</O^b/#gf>4XLP&CcPd0[Ka@EB2?dGCP_bc]>L9Y.>a6W)Wb_5LF
9B:c#J5/)A@OgOBfD_G80C>.)A?6@,a+7=(Z\9e\Y7eK6-fAg3)[(Z48)10N_PC3
.?DNP;b#7g,cO?=ZME),_-C-GT+f@11GZ)UQ,Ad5:HCN]X4SGgO+H#3HZCXYcIaF
NU:/GF;)EB.Fc+K\F>CQHQU([]V]gOM9Hfd]0GK?.N_D-Wc,@.EN,&-7).dO#E?K
1+B=Ve^eEEc\e4K>/gA3GY1Rfd)g2(>Wadb,Y1_aS=R^YV>2d=HR.)Q.>BGV1&39
JYeC_VZ3Va1Za\D&#FI:7D<WLgZ205?+dC=Vaa\9GeODV;<e.Q1+QK>1ZDVPHWSG
^N<+=WZ@6#Cf,O7YX[ASa<cCe/>5DS(.1L&9OOMIJS.6]>#((C4@+)0M[@TAaRJ8
.8>#_11aM[HN1eC3H/D9(@;eC>QNG;A3D+-/_a2:S@>9eDG[2IP:8JX9+?1614Eg
H7J1NL)BY218a(_dAJMXQYQE<GDI[EMWLY8Q5/)^)G-Ka^?MZa1:^.A/bDWgK1>d
Q4FZ<a#S9<)(f);B_GW[a[fYE9-OZVE^\K,3Rc^:C@H>TT7Q?XcP/d<8:+LfWL]#
fWGH9^G&a3IUDO\bNX3<LHQ\EcYL=78D^=.Q8K^ScP(Q:>@I/Z_8&#5&=CH(JUVc
fg;#U@@[CR-#K>f8#HC]RbFVMA@;MT?_4>KC=0ISdFH,YEFADd/<AZ<^S:bF.73V
;0@4&4//WdWd:+IcZ&4_HaA-,5-M)BM0S(.EH_dP((KId7/Va8[F-<>^RO9W2M75
@NFY0VT[2+3G?=Z)B)2TECBFD>U5A[UICDBe9S\V+Z,6B;2?O:E@Yf4-IMQgRABe
@eYd>YMbJeXH(_:EAM31WC<6I13g:CS8/.T<Z^LLZ2^(I2W8EWLfR8(L-Ra(2a8^
_eDK+97X+BSc-?aGAS72TO@)ASM92-5)P6I<<8=>\M,586,2+JOD#3N=,?NJF]&&
/cUF1=SLW86;N8:.=_[Pg:7&Ud]d@S?&MQ-6-MN_Y8OcS_E0]@S1C(fDJ/(C&I7U
\LAV5P=+ZDO-]CNL]7^<JNC;;9.KQ1F[=Z4PH^DX>47X[:0.?S2NX6ZVU/9Z)P+b
=JURRN9[YPDGS4dFM.&VL?0]Lb>P[314J-0/^QS)TU@+]Z0dN8ATa3g)_R;+6WYV
(,4]P,5A][b9<6HgM\FO;R^T=B3dR0;(?b=\8c7>Y5@DA2OOB5:Z[8aB]7WK<#Ja
O^?FbS_UK]G^RRQ;8:WRH@<g/(b9Of@(8T,D?(U4(2?4UH3W298R#XF:_-Q]4<1<
9GP@G;\ZFeB=H55f0KdPBfEKc8OZ;\_#(Z\)O:;M1=[U98I:BPBY2+MCUXdJ/QM1
[-W>>MY[b+\L#3E=0\KS2I)QbgBOKa+/9G4EGQ7^)5+ed?#Xb7/^<;>cOY)&882Q
0LWWf[I7/4)K(RR[?6;X3V15C_N^BCH/fg)9TeO@ccbaH@O(>^MANL7YdX>Q1bCV
1-RPFW26H-SUbdTXC_5;:IT?3FVZ[#FIJ;D_@7cg4fW_Lf.BJf1H/9_KE1[EG:d&
LbRB;R8:aaM5,B&^dI23cAfOB-^BNZ+2L=J9]>LN?0a4Ta/E>B#8ERB-E3#F8(WX
7XP8_;c=C<1Z#UK;+&@>C/:Ra2.3#FcU\1^Lf<0bMT6B7\6f82D&6)PAe,7().TW
a]9+].Y@f]<Q9RYWgR,Kd0-S5P9fP[77a+cPeY6)&Ne(Ib+;V08=#]=?bd8J#Z&>
\NPP14(T3UG+-Ic)U3B<C9B-?d_7-TYe#cPEQR_O4S@F-QTQC)[8bZe;@4@Ea.5+
1=7-R,1-GYVV_-/8(5BKGIYWYAMP:PD6=.Y[f(P)G_/<2-4+=EHB-V[d31XN-ATC
S.(&Q4OZX/9<;?0BY8-N8LN&OXI[H]?O2/?K=5VJ73=\,OE.3&fC+A[UI+f4+K/^
L90(D8aDMYS+M);>WKIO4<\A\WBWf3>[L)YF(7AY/SZ9aH-UR,E]9DJK2dgf<a-G
RB/&a;0eQA+#?>4&e^5?JbR[)T/<@fCOZJgU,XHZIf9WM.c]M20#LIQAR,?(BF9_
[-D3P&4/ff68YEJLcP<.\U9886-:Ob];V_HQAdXGP?KW^\FM\^J=(W^ab_P9NY.3
>M:Q#;/(E]J>b?NR[((&abcM\R8fU[6M1YBE:NN_R9&S<MbB@C=[gA>LOc#d]Xae
Q8-0c+X.H.UNd6V-&ASOQ@_FT0+Q[K@EP,_3_@ITSI.>c7=^&#MfCBUO<T<ZD[O]
8;D.62c^N\b\Y5.B(9aG+>RY7W.<Q58?G9?5_3d@.;a^+<&ZLEV7a3gKcSJ\P9#>
b((JFLKCW56[]T/Z@B/U]Ud5HQU-CXc2aDVOXN9FaX(G>SE)3SP,dMb42(+P\E]6
6-QKXK05NKB9<,PW&/eff/9=<=[>MS86(X,:4e_QeXBaVfQ44X2QI62?7^YHN(gC
TfK@dMaCRO@9Dd>>F?/33(J+8^9O+<W?JEU,2.^NZaZa#gU<?f2R.;8V3:]8/4WJ
[NP(#3AZba]YM<1,5\+FPdTe(W9:g&2H>?Q#c)PQc^R7G>37H.4CKKUI?CO6f(JV
_LDBKbFf^,>gc-3T/?VBX3G3N+/^41J.)VUd@50WPaND2dME0L>A)[9X-NdFD,U;
ZSKOdX9U94CZ-VIY).8[AM=+_9=.(ZJ<b<:RTYLU(9BK2<J7S6B(845O[?H?d0@J
d\7d,/VX)I]-AJDV]LA/8W..IKKcD;&X+(-5L663^I#d<U\#CR./aGK6QIP?@&G5
?gbRcN_28F#8C0AP2L/JIa_KL6bF,b\@LN@6Z;7<.A=eG##,^S;5]XYRA8HK-I^I
F<>ZH&A_]U&(YSCJ9Qg#UaW)BM3=6&VeK8K@M=HX/_P&UWGEIO/E&)24.D5&&F;[
-WP<O_L4U&eD<:FS_IE^_9#2(1(DAIA&_QA-Z/5^Xe+Y8CAQ3JCZW-LTKeP1]UHS
M3>U+]Y<?7M5Y/G06<#.E#3(>)\4FOP0@>;@@KE7REdM#@gO(X<OI/R<_4YgeO[+
F?ZZd\JW]5@7DEYd6C);C2A4D7_=[]a/)dZgJJa8OS;X=O>>KW-Q6=-NWd&QR=@c
L2Ee^=U9;g5Pe\(=d+/V.HQ.0^:<[CLW1W@c@6OZL5+6e/4BU(8SB:\+Y[6eE/D-
eINc.8&4,1\eYW]688+g1=4@=6b-Aa[TM9?Z?T++F&+AS&&U:I/8Ce-^?0A@-\H<
/dD&760((RN<:;cfV)9C4YR3C/J?=@^>Y=c#dNH7<VI^Y@M;ZVJDPS&GS_d7FA5L
6@=<>8)<PX2AdNH0;(UU)J6MV.XaPU\f24BF2<WO[b6[_D\=;34M\_Q,5[/@a=[g
Je8cD4b0bWFNTQ1YEcUC-@6B[QfXV<LAe)F19-Xg(Be3+9DF4GOSe^:\(K/@B<eU
fK4G+#):?/QG;Q;)D:H=Oa2&AC7caFF0E9/B5Z_2b/R;b.#^GG^b5)R3)[.L\AGR
7MS4Q21b?1Q:8L8&)8b^f,g94Z<dHVW(IEOAJ?cdF:P05LK(4O@XNV3]N,,NUZ^J
(1f7gV5M_Cca;;CZd(1d.[K3?:1WF[UE.S>df0I;Oa>ARFSI=A]3S0ZV982/eE@g
&5_7NFbO3\MBX9&XZFEg7R;OZL\O8c93+IMC>7^.D(f1P12H<HC#7>-(GD#>8Lf6
]_75(V2;.2^Va(\_>_8a9Ndb^-=V>1-BJ)CaRS2a&(,+;=UdGM?a;L[Mc2Mc61-I
SH@gEE9WE7)_#JUFYg-FLE(S4d+]6NC]C:\7V,L^>J+L?K5]K,0.3EBRRE&8?ZKV
YWW(;JX&#MOfF.3JD>[A.U+0BJ&4GcKddHg2HM8=)+Z\fZBDK1HN>7X_O/7UA]Q\
D.f;GO8D-/^W]NLQD@a-7GDUFL17&INIcLT#XfZN^:fdG[?>KaDV:C_&c26M53K_
ff]:c7^TQd4^F2J?YSWX#b0KR:0QBO:2S(BM-5LVIG\.&W3/1IWN^UY]9fGTe_9-
9?MR^1F<NPT8dO-L=fY33N_U]_O7BUOU-QfD&AR/);@T9.P3@<WY07>6>8\XH3JZ
V0H(VN\0U\d)1@)<GT>fL=#Y#ZS[9P[Ad=eQ,c2?R&+[(\D4BQ7.Ag]?dN8^cH^^
6G#DR/&RS@=[K#e5E;(S9&@ZBHaR,L/P?gP#Z@/0+WH8;A0P2-6JZUHX6IN0M5&1
ZGK=[33JM0<7D.NA5AH;XF(EW,S8bB@;M<82f&(QG&]^af@98d\G#X8g&W#?ZF[;
6Ze<e_<;[=Eaaa\5C:e:3]13IHT4@N,R7.+E[EZ0@8Fb?+KVF-)EHXbSVW/6IL^B
JXgf9O0LRa+UMEX6<>01Q-S&FT.+&J\7a:_FRbCK\)2X/d)1]U&))FfTdTS_)[W@
AH_3#>/LQ3d;f-[V;]FFY<V7X9Z??4KZK7f&egESKDIV:O_f;,]6KOKYe?X(#9_^
(@U@W/#-3A[ZD5M2A+d:Bc?YPS.UZ\A/BB(]\#?_OcYc@&D[c_X,:UPJ.+BgMbF8
a0C>Aa535E6HNJ(0C\#>G;#:2SB._UXdDD14D[[U,T)>Te&E?I-H:W,XN=#N17T4
-F);XAQ^<)&)0KD1LXc1S&.,H3YDD1GgA3;/&2TE(9@.QDPf^(HS5)8K+_RdN)<I
-d06d>-Y/IJaRL&](dND1=Q42FHOV1EKPI.Ob:DQW-b\a76MDWLO8JPb-990EbN/
W1ZK(OB&33>Qa+f[b2(FB^PcZM_TKa-H^T(\5Z64bTbc>4,173&T6&Y5D^),V7dc
YIf\Jc@U33bU(6f1aVC1d:2&Qc<)A^@JE^3<g86c&8g+,,FG>,QdJ\XVPgT9;.,X
3K^7;33/a<NA<53)\.=3R5#^C@8^L.T#^DEbT9LAa9<bKZGKEWFNUE9M?\6;@GDG
>bJ3@)5TCNQ&RJP]RXSV?-0C^S..ULd>:^_L1-ZYd:Pfg)IBSG5Kf9>R6X/eG3CC
;MW?)UOa\78-UXE&68>X(L]BVM.d3dK>BKT_9Q,.gEZD#Z2J],8MWCO^.de=B5A-
/@b=eC)ZLQE4@b\M.R>.:8P1>;@X7B^2LFV\T+b)@CR;JK>Re.IH1K-E)H),B023
DKWgd7.^e0MQ_50CXC=fa7(4[\>BCW)^FeZ;_?dPL+T>UZP?(A(G\LK5\&NEU\gP
?g79-N#J16D>F3df&X=O1-?^-efb_26=eYBECCbK2+<^G0d0@C95^;]^+8WR(gZ]
:AQJ:3E_>@b1U[8\&K,[6/TFf/aRVWeWQ?29Z_bQ8&VIcA1SKbN8ZTXZ_^f8A\EM
,c.fN:::)HLI;/W/;G9<1)KEUa19Vc]4e(&3WXEXOGFTOS<e^6fSeYM,CebL>1RX
8F>@:=KUFbAIIUAYgW<S?b3#/#;/0,I8U<,&_D)0.@A[XICW_G6;a60HL#EfW\Ce
c3L+H78JS9W#dF581BLYI<8TOKM33@?-cB5K=>391L?eUf;VP^@/UOIH0G;(KJ<d
7&P^O3E-V3(LP8f@;#]IYUT8?1O^\9HUN<#g9]7E3+#R9;XCLYae;54R8/D4VFF-
CF^fKO^+O>_7LRFJ\d(3-T&a\S,B@_TX>/&]PK-Ag;W&1f=OO-4^LI[Ha&E(C+KL
d&QT;d<+:Y[-7RNYfR3gDd:,[4V:N.f2U_]M0Ib&CP:-M&MZKf8.E:Z]b>McG?Zb
O?Dd\E[U^WX3aK)9C^AC6/1/ZM87:[F2U\Z/fg3W/PLcZ/][b46a2(9/<ZEV2TV\
aI2UdZ9;aP362AP_Y2D\K\g5IZ^Wc(TFW8<7KQ:S.Q?:gJPI8,C8.38E3Q/d?g&S
N?WFS9?CL:WPN-+OGRY0G:Q16CfW^@/:??>R<::_D]\Q]cYB3V=.P3CB&fbCdF9A
2Y/WW;^f_C\PXV+f8(<U(LQ\]F=;29Og2[CSYGbRUUEL@Bc^07CPKFXZEZ,X_Jga
[aA>:F#V?##0(I3O=2dI1S5?-CgbS.^@:<DPK\(,5HPbCTTPXV.+7I4g-@44JEN(
QaR[03@Jd7A/c/OV\R:_(#HRg#B:a4(cD9VA-#]AEHbSKd.T]a/OGdZ/W@Qd7PKD
2=(ED2.YDD[=FF&#&=]Oc,f>@J[EgI)D:O_F0-\N?22[:&BMgZ/1@H\[W\GcS<UZ
9b.b3ILBI-Y.LG>5KVQJOQO?V[/Ug]YG=_//egBJ0FV?2^Y8+EcN(:O-R@[VAHaO
)C+20U^[A+fZLT\c3d@+b?Wa)C[+Wf2b1)Y9b+M-V;8:,SUf;7Q0S7)[1/Q0I[S-
6eDUXNbb&>R+\AMRK)[:C(B12eF1W6#_Eb7+OW2Pf=)7cf:cbNY)IOA-g^WJS2<f
T=45SbP=T6V]Za<=8,0]9gHBSEII0,2J^/:1.gXAG?>KUXcK?dVeH>WV.FEI8?F\
FD2f&M\6ZE6(eKLeeU1a=H#>-/_K0gDH\/X8E31\7P?JJ\,FP0d#gJFK3#Q[=[S?
(PIE962_0B?JQ^>+XU@B?B_#-O[#T[]+,-eaH3eID6c?H<Z[g/]6U.\7\5#?Y9F^
PK?fTD1CBLW.@.&\JWP=[AT6>1M>1A..8CB)#5f7/I__e@MPDMV0P_54^]N6@Q6]
G5YUY#+G@.&[4^&JT^07D3?>XS3_E&=_(=d<>XfFJCRB>F1)/=V:Zg5M25=Q^MF3
7H@)GDGIJOR)X^+R#>V.Q&Q\F-b4\acTB.4^I3[W[@9F9Na[9X=8X\Le9+#Z<7EY
\#R,D4F_gB0d8Uf39c?dZQfPM>gT+AW(Lf7R)aQ_>/BeCG=JE7\^P6=G#4\;0ZU/
V/:dVM@/G9DDO,[0d.]1.1]bc.8V7S/ZN&BMga57H.dded[d:7]R<PBLZO&F^dV+
R;SR,ICV_-MfJN1;?Ka0V:e691MW[:G&?+X]F-Dd5Gf>DL/2WISeX+V.=ZDcA6UE
C/gO76DNC2RcB2-Xe6W^X(1^b_L(a8A).8,@HGZS]IQ2fWAV\L2);T.Y,b<aJVIN
>Q,=4g1f>P[.cM/RN?O>b^:0]1W/+(>MD#3=0Q\+W?TXAQ;F9?M-?-:/NJa&dM;1
Q0gCJF4Gg=1e9KG6Ae+X)Tg1+5^g=Nb0YNKTBZ;U(I42dGHI0ea02V2R=L\PdN/_
fX0gb6/B=EL.aY:Gf:U(S6]))TUA3V0<S[OJ7@g_G=6UK1&BLAFKOMVFR:_=E/.M
FP;8UGF&4E,:XMf1,+XYZdJ<NLGK](/<9+1bdC94dVUf;F-I\K3<)e:0b:+fOdNZ
5e1e7f^HWG=gXK#X;UT5Z@T(H-6.T]CKZ+>WM.V0eNbJ1<)522Gd#9W)SKX7[8#+
9G,de22;-dIfH+-,aW/[/KT9=0EJG7VB1-ga:9a79gc/gFSGJ@4^<eLRFZS;?ML4
W\?R;Gd>4aOW?e).Kc(Bg[9<9(+9@^Y#8?F[,>b2A&6/&3<&?.A+HBMdRf@.\-S3
,1O/Oe\S.]6D7UcdXK=+2N8CG;;YegB(NGG=XZ62aAEb(?e>a7^/A:?XJH6gA2#f
N;-X:8ZZ0Q)57)8,=CQIRUKEV)G5B7@IA?Yd\F7C3dG[JB]-QK[5RT[a&A0HaL>3
0[f;fS(UI\ISY\Zd0g.fE?:0Y:eIWMJ&BYg_BGLDW0d07GVM=3_DV>37X_(U#E8/
5[_&b?I15862G8_I.W>5-a&gKJQ0X>b^JcFG_24/2;>QGTU9\3R9I,,,9bLH17,Y
&ga<b-#><aAL\<:90P2/3_F?.ZIE[&1:4(6VIR83?DK&UQReJ&/[_GHY+1VS>;VA
,)TOKa@ERRb_O](3KV2a]C&;d+JFge@Z1S@7Z.c_<Ye2HW1P^1UfQ(1@]_#UW0ZG
G8T9=QA\4d:;=1(@W1TXdN,QQY9-I:P<gA4Qdce=?,XEb/(E54^\H:gO<b:GgaMY
>HAC0KY7]L#(YL2+9Nf=CO,,;EADGEDLaf9U^d]_]\3_a9a(OZ)3f\L::@df,aB+
&5g&2_/>9Od28a[=V0BB_3fZa:eVE7I8[Z9L&/-Wf^D[]dFN&(U.X9/9D[K;c./A
g);I@>8Eb\e1<(:aMWZbWP)<,:0AND]e+(G89OH?:W?>JCeeA_c;daP[I)EG,YL^
S4d-g7>^_]ZAPZFfP>3W&&E@43JT^N,3\9[ZLSW>Fg]JgbX(CIKd+(KU51gaEPc_
eU9AW2CIDXRaVVL^QEDC.8X.a1,7LHG&IF)a3RR=?VT3VR:X6+0/?PI3T.aOPNa/
KBd,J5.95R#EKO&R?:;4&9ID-Z#]CFW/c7b->?_a(dHQ[7ad=(,E0(S>+G?Eg(W7
8PKJ,_:BGNFOgBOW7HE&-1,V4b0,TN.1<OVB^5TD8#2bHH6X2b,Y5]VbU^e7O\aA
-F[/f8V>cJQa,dK1,QL:gb4L4gTL8@/H<PcZ9+U@/0b5&N6Z?gF/(T_7:P+SP([7
_f7Qe7LEX.:Z5ZQ-L7+,SU.-5KT_g9];/E8BD;g:]?V^<TOW2UcREQ,0GfG4FT;:
>60K8J>99GWSg?6c_4_/,>cRe#TW:a,1K6ddM;gQdV0)1@FgT4W&WaA?a501WTPZ
G?UL^/UVAD8T5C3WJf05F_;YW,Re;=MR&(YbQ:K7S=.G1RCAO,FAD15BS5eT6:5T
-;Wd3WQ/&d?L.,/#\G0,K[M+g^0NN&TG&aWLdW,aCW\HAga7J#&gb3F^J[WRa.f_
-2Obf??cHYJb?WO0gC/a13O+1/(0JH@g@ZA#N1<0CO=8L8W=\7:<(f?]Daf,?DgK
ZT+/E=\Da=7<CU+9OM0XM0bgfCXN&gbI83+^[Y1b7Z@,\1[K##gZ\Nb(HYAag08#
ETDffV<9305TF7B_@<A3/8TISSD+A.b(Z1bB7;^?:+[4R5C)]4[3NDRTVBHQDDIE
.3NJ60Hf+N&=[@eY91I0Y-^N3^(;Lg@1PIP[W&Q1>P]M(aEc\SEAfWE>E@-L9.?^
5A0@O[D+H/@2O^HM1Ze<1/_>M@#A[TQa.\a7cS1aga1;fV^7FUUPI@ICQCSZ];N#
D2Z=dCS@<EJLKK0@GN+T-5LV2WR:T/)B/<[FOIdQ6-,3XH8;PQO1ZPH?0\ATL[Zf
:W<?d\N>e#AU5,DaPXMaZgTPGJT+2C<Rg\agcNKKW39f[cQC;U&7&QH8#+RJ\#aO
U0If4ZL^X_^g[X1bbGPcBQ_K#>)gW01;Q2,+Je:<AgR15f9c_QWSM/XY&@L1VVVa
@>M_.KB>.3C2X49HZ#44K)V8?=g0UDB&^GEA2\[1?T@fPF1=g=JK#6+c7J^g#04=
M=E[(D9C-\cbgI&fU\OSS)\MT-AZFc#,@BE_ZbULdST2=(/SEZ1c4K(BS1UD,+JN
1;JCXbE\/VSHg^AE2OE&X.G)^+Jb3&UTS#?1V],SX+@a1&4b6PeXcY&>)&-8IHa)
Z8cF[;?8KcSbR8?JFBQb-X>.AZ]LS6L(a:OGT8[e_</JgH>Z;4;/0+JO6-T+M.95
V7I=bffP/-(\2E[D?(&K_#Aa[J9#:1R98#6gESJ3^5@)OIK#G]>MGae(6SVP):5&
e=LUYe##]#H@8[,#R?_W>)44V&DD)943]7Q^P,#P73@13]GY8T3ZF#+0^df:U(#S
X@J5JbE0VC6PX>><9HX3;;BCS7J5O:bKV_P[\X1b<K:DCd=GR.TD2U[4<(V8&\eN
3OAYNdMdE7H_DX-Y+P=/e87&M)_<&5W(?L28_#d=P:d[D,/RAbB)XeF#3#O^>/(F
FY&Ve9IA7FFXX1[YB@PXKNF0DE,YI=5U)TFefPSL_1^BZ9FGg--6(fY:cQ25Ia<U
&I4N^WFT01J:<R>V+G(X1MHKd>O;Fa/T;98N;Mb//0@G9/L7YU]G@8V-RSR[=3M0
GaPb2H0e;=OIST(g.^]F>5P&:,X6FA]E#7bSOD&gP:dRC-3V-aG7/<BXYH7G6HR8
#g,-E4P;4O)c.YXKH8Qg+,B9#YN/B&d)#VFNO)EbIT<I##\F/7d7[.BQPe_6S_S/
:TA1[,fI^>gd\/g>F^-YZ:V<NO8U?#PCG-V7/YX],PG.>I@XS]BeB\SXI2]032;)
=C;U5]Z=0_g4dV?B\-0?b-cgDYU.;#?R^4;KOB[Z04]=@-:>2b)L=9b>Q@cI2BBf
K7WNPU#24<G,]HRMOJP9c]g\>(52]e&-LP(dK:#Fd?@g(f1C=T;Nd3CSAS.J,B?f
BT0?CLGd?_@U4L(5]9LA3XOfV4Z-DJ0PcA^:()A>9193-1f3I15H0Q&7^40g:\[f
bQIG+=B-d:0Je]e8?+S,#(_LN0Za1.01&cdOg^K#BEB/#0?^^d#>a^.&IES^gg?I
KR]C<XT+0[GK4J3D38cCR/f^43OH:N2Q;c>+IE_T?bQ,NK);L\=W_,2aT6?YBSOW
JI.G#:ZHG0C\XgA(J\0,RAA)WV@c-:B2ZBcQdc79O9G8X[EO,KW8#I#ESS:S<LVH
L6.>Q]7C-MDfTFgaMN:/?:fFZ][bNG<\ee7?Kb9M9RL.=H<D?7]bOdE;.L5CL7Z:
S4YNZ=AP8X_Q2+P)fIfST<8CHQ3QU8Pe/8@3?PaTGV?>:Y;H:bQd-#g^1eAZSUg>
9g_a^I)4\8A.<)(.2?7+[3dZEMR<E?Xf7fOcYT,,;PF3#@\3T]e5ADU4[PW=X9J-
89AaY>gWEQgJ\;]/c6V(3]+),fFd_-#E@\,-)S^_Y#R@]]fJ&bBO)-Ed(:H=0:,+
.0QSdX?&;D.Bbb]N<,BL2+VAYYbZ=?T7_\P5)gS+C0Z-B<QNO+gJR,)DDS8cFJ/[
504.?#C95HE3))Wag0;2J0_9gdfPbULF=?3[N-TM^PfZ\f?68HJCU]3JK=.Y(N/O
B4&d1QR<4E8[a8b6[[>S/+V-Q)_Y:(7W_).F9ebY#[TVJaO1^F)9^H[&KDQ77Q55
gO1Z>LfR?W<+9<MW?NaaX7F9AS2]?7[MPIAZ&J?G.,A8D^OR4S(\Z4)QF1Z4.)(>
fCC\PT?CM4_K91T6[7>>@K/T+9#HKSB8;^ZZI5+M_aWD1GJB]S>_7QMgF,U7KPD]
9gTO;-C7gRK<dLRZ-C_29D6aD6R,fO<SXcN&cZ]H,H=A]bf-bC5_?1?[_TT&E]V4Q$
`endprotected

`protected
2V7@;(XWgATAc+,)SMRY&b=RDAa9bG5>DAF,L#g8U;G3J3.]73TD1)B-IOgWVA#+
Y^@Fg0I;>@I4]H=e.A_KZL=R2$
`endprotected

//vcs_lic_vip_protect
  `protected
F)/&8J8ZW^4O=U)Oed<.c8efU32>c5YXV:@W6)XO2,IX.L))fdV57(E[e=B0(DR-
7&?U[##6/<<UH#U7G^f?WcALB&a_68ML0TN?G^Y,FMc5\2g>D:L/OP@,3/a6Ha5F
E)9Q()Na2C572@>P)E[1L+N9KIHK-:C<-T;MPU.JT_#fP9YK5\+8De:L<.8QB.UI
DYFI)?2Jd+XB-I&SQR?+EZ(<<]d>ge)ZRaXM,)I3QaV>]>96F@.LU;I;XM?G(;-:
/\MR2AE(/EE/=+U_1?#SQ>aU@0fIRE:bbX;REc)L&M-<Id-E?NM2.F]E8H?:K>Q8
FHUWK7faQWE5/9fcET3g;J;e6E-09^(ZLV.QS(>5C;1^G4WT:Q6&VUCPC>B&:]B7
WJ13.&-JTR>@fOOUV)]PLI]DLGgb0W-?O(\B(M:\9a\FX@>+<M7D2#U;&\@5bG6g
.5fT>dObd.C&XE(?E+<b<SE-_f0HQJ))[>e-G+1,a>0VJ&K[Mc)OPaCX?P^\HV)c
E>1O3,NTYfdCX]@HUaJf2@8,Z3(T#WcXYaS<O:)6_Pa[.&9?45E/FPA]9S:LOO-C
<fM6#D><XT8#LIYGAGJVK)ec-Y2M5CR8R@K9SI.-JMZHJ8dDd.f6B#cL>+\f>W=I
,FLcZ3I#C,73Yg9[9/AX9_U=RSF;I16X=9Abf.WF9MBX4H[BS(6BB8D;:+TQfcSd
3[4(O]eB,CB&/G-_1V/c@)R..C8Z/5SNAR&C^,373,B>KM)AL6SHM;(_:V4OP+@P
\KLF/:K(Y<))(;X.eg:?FSMG]]A=-4R.9+,MFN:G8229(E9[C.c]35I^D:cfK>fB
CO44:G4W40Hb:@JOSRB+L;35]bN[>1G8^HeRaPA]QB:=4U=]-REL\;.KU.0ESH2L
4^=aV(0Nb&<65?7_]UK1KS7?I3H75FE#,GU=X_;8Ya#2&.)L5+We8Y6CaM-V@-P0
H::\<H^eLf/=[d2)H;X(?.4G[I](12e[1BS6SC,30\-L;:],P_VV]5:F089Gf2U3
?>>:CD=e]SV:P-N@#]OgZQ_EN[>MLf+=J_+O9[)UcNAdHP^J39&4O9d#18=b3AI6
CQ5LBfY9>,@bg/+-:T2MRNa[8R31<-QM[dBFL.&>ZU@aB=TDMSEcdS]AcS@^?6.=
_X>-GWC44f5cPK:A8)W=c#TZL;Ua1:=?B]a+LNQff^I@_V(SZ>25[Y^O(QQJ4J5(
.K3HLT23&]NU773Z_O_O>4ZLdJ28)(<8C9RU8Cf[Cd2?5B+?(9BS24bFQbfOTb4O
FB[E7D7)/Z_,J8<SaNTMAQUX3MY)1.=JU6_>:\I(,0L3<4JN0J:T85<IJN4-/[_O
SBf+(]DV11CY8NEJeJbLBaKE3+c5&LQKL-:IM:YF@+fWf>IXF<C:VfTDM7Zd,PPE
?(VDg;6+;S1>CY]K47C52JOfBO,IQMbY03OVG5N4fPO[62gR-]Y\Uc4:V9V4.+>)
X^gJ,&MQX2OIQ-EZEef)@Q]XcC9LEXce&?MdXZ+<+/(;cKGG#f4)G,[f?cUX/8Xg
)W8.WfAQSgcRUN]@W1&0YJdER?PE)4c6UT__.92dE<7^bYTU59ZKM8QY(5aP>:Da
ZA;_bg?b7dVSdCU1e&,g8?)K+(PH.YGYJ5C0N[HJ/KO/=]=3S+E+F#^;0GR/NUAQ
<F?4WCfX&I2YUg:>2@E&NNR^+WS\0T.K&N[X9LV&=?&/:15+WYeS5/>>?ZKY^H<)
2gOb.GPb29IP&CDZd^[@(4fSU@JEJU3(Y\-U_YKEK-4KLRPH8@,FMALU.Y\K19PY
\VC?,?WH0cO)>0)F\-\:MQ>VdQbDE#S:.,8X;(ZC[1V,+R<[7MedIQ>YCMX3W?1>
(:.=N;Ba39VCV/;>/eED8fZX+\781?T1dD39#HIddA.D(I-a)SZgTS8)8UESZ(2V
7&gKL^(QQ1S8>T7-[GI8&<,EX@^_3LWZ5F:/Zg5FfPA-CV-NHf7#gZ.0Pd@@J]&3
-1#CV.A^K;#Y25U9]3)__;CK+R0Sb)3+A@\KUYNW/CJXGgC\KTE&N58Y.1+cU=GE
=fBGE3LBO5F?90ON/6&NO=69EN2()LGgE_51K,UMM4)NMP/fDH>EeX+F/da1ge5#
QBW(e+J6__,G_0V9N<:aK\NKU?SV+UOG&.4c\_\V--K:E.fM:K<QE,aS^<8/4NW<
e#1YC]E;#;&E8OW?R]Kg>-9eDQ?dI\,MRWPL]^?(ZN8#33ZWZ:W1S&12cc&UMZ&Z
TMK^a&E4+?32X@GATTSMaF6:3EEb.Z>cHFU&O-2Lf:c=5>M.45\[8F>1A:@g&K=@
Vf]QC.>(B1_SA+U/<LRQWP[;#,.1?_Z;c8K:4FbgO\c&c+EF34LK>0K#HRMQ7)&)
62gKY?NZR0@cB#81@>Nb=e?CAICFSP_\KcGE(6G3B4-4D.T#N^^:0VD@KQa?]^H7
-Lc,[]N0eE+H>7e3g18gg)Z+VQVe^LTWS>6-WJVU,KN;G)L^QR<a:)<;^0_^2K]M
<P_5R?NVfX/WOWZ?4E0B/C/=c=MP#]<[SP<,&1<I7[QF^PWg/D#73YVT/dPECLPa
a:H[.NeeD?CD_d<a9(:12D)bb,bC]?FK#a-=DDY_>:T@bg<A/Z0T;=S]X)8XN#22
XV5@-QZSU/KdVY:JddScF:VXc2a-^GXGQcB<>?MN3AY[196YK=,<QUYgU+JPQ]LB
T6)C)@C\_D?+Rd/MV+OE8[;Z3<bTc7CZR1_K>5#L?Hb[86N)(#ZT&##2Z\T=\650
:E\d31+M9dQZ7?BHZZ71FY<2a.=6C1+3#M+=a<c=/-PUVB,)8H)e1;ZD;2\Sf3=A
1S8dc?38>]GOF=(N;NPMRQg562(b\4-Sg9T-+:Z,AZ5F-@EN7]CYeBII/G,9CRXM
fF8^++FR5C]RAR];f+]0QV.OV7)/\=C61.W)(WPMGF0@,IW(.a.FMY7(&c?7_AM^
(:UFV2\aTN153;dN1f4BUZFS[ZNWVd2&WG@FPba>6L?4I<a?<bOR[+QH?:Z^)L0^
gV]-e.QUYG[c7aA-Ra,_X^_@b;]KZd7Yf]^aCUIKL63gRSPNeA^WHU=\c3RT[8);
>d.WP+[B0[/Q=:LACdV22_>Y,IXD5g#0DG_/=P23?[b#@CT+)5./Ofc=8X+-HVaD
_D_@.2^^=(BAP?EN?[_31)[\6TA4:,aQ)J01^1E:cOdG^+c;c@cc8c+B:T7bT^28
2;+]9IU49>(?.\+\)4UTFF@5A1K./57OE#VHQ3QSG-[BN9IZ+L;;-g,>U2RS))=_
Pc\e]X?^3_A&4ZdS[P<>P+:@\2a(WU^9)ZLAKB@AL^3.gc_/2WgFbWSBKYgCeF;Q
ed(LF(EJ6G]Q.E[5P&CgQaHYKHHP<Z&.A(<.69_I+])DIW.T(<>3\?&MdB;3f_=2
+W9PDA23@FU,PRG;])(ZbSR:89X6PF/T:QO@AO__3]\(88&8FRPd+:D>f8IG=V=H
f,AS>_1_;<6G>EO+Q&CEb3G#Z8Be16)eAXQ1[dD<CO3U4)(?@d3Rd)J?C7GS,+@3
[]SF@-__M,^EEFEOBQ+(#LQg0KQ.e2X+EI5.>N7.O/f3\RI9.,9G786/545F76T.
3;YQ5++Y0-B7g1@M#8a?P9be^;,L3EN7A]eF);cEDUPLN(:d8VL]49R/g_V@4W23
I[:c)F#a.26>#C^?QESF104(Q<56CM(fAX.#EJ=?c<+C/.\J5=e(IP&/TXH[]W:?
C2.3^Z79gRXUF7>C]YD9&6bfcfVFg0\(.>RP3S5H^2dY\=3UEMQ/ULXH/Jg5SRPN
FZ,Q.aE>N@F&C\HTN+gB<X7d[aTE_#D;>79<P#4PZPGP_e:TH.>@:X[B3EZT4=^_
ZB]5.X3H_]EE91,0PGDVgG]\PKF^)&1_aUC@eM>e)A@3>MIW5c30\Y>NZN=<MDK(
>JC7H;HP=UdZ7#5GDQg>b9E/)N>GY^:K\)EIM?]1^@TTf#QF1,B]6f3RTHF(O?N,
1UV74=>#;.B.bIDO2MRL][5a_ZPX4Uf->FY:RdGC[a(\6;]N#TMbV:Y6?]IJ5F(F
P3-3A,QYL,<a(+/g0H.4#RK1)[#AV-:O1W]5Z?P3VL52.Re^W@MO[-6:F[24-OA-
(Nf3=D6;MSZa0aR<I1K.OCVSQ>T-9DSe=f<]AM/XL]Oe3:.K7P5GNbgg.;DPDO+g
\9EY^Z>U@B?aUVSL4-I2WG3X?fAcZa-Z1-d1G0fFUZ<MUR9dASY]E.,2O:QVc[NT
-dM>F[fJMAW/edQ-XC4>M.<J4A@/L9,-7BVV95QG#F8KHU1JE/@^L:bca<HIe#S&
MC1Z+C]MSFa98?X,_b]&NQ]#:?)2DMQ#HbU.9G[B)7F?(<VHGMAVQ+Z43c<+K>Z3
D_M4:RJ=P]3(2OTDZ=MBKJ62B81@aQE]VaN8X<^W7^a_I6-KQ>13J<@6LSF_/PUC
KN)-W]YQ=S;5eN:F)HP5U2e?#a@4TRRLGd8-.8aK9T.L1PW\JC?-0f;3[S/]7:0,
\2Ga9\UJ&?Gb5]Jb^F7/8APL)])9AJ(8RR>>R>2K#VD48fJ#-M5#+8.&E__#XI\B
B@]7DM2S0?XY5:BU&DX^LCJ.gc;1SSG.Z?ST+@+HBIPKN:7g;@-0-BV/=7@1S&YN
4/PPV>W+DBC3XZP)7RJJbM3d8(9&>0RaR6]BYe_ee<O9?Faf[?EfTV)SN)e?.JJA
0)EGAHO0)#2H:E&XPG4A_\-&0IKab&[CD(IRQ<L#GeL+8J<7,T-_?E(TcO9(C1;-
,I7bMOg9SO+:@bfb.f^a7WM6cU[Cb0FbYF3G1JFO)C&=O<f_7&Ue3g2RPI(c70?1
7-R:;X]7O,K1#?2Yd8&)A)3d/cYC;-KgO_^38:6&X_<5fEMaN2>QVTg2VWM-L;1M
dIgMMIc-9f-^YKG)CD2W:bLXK,e^,(9@Y>RRJC\>b1MPY)YA<,NFA.[I+=<8&]e(
O8]3g+bJAPU15&CWUZ_f.8/.,EMdM>,X3P?RX0/>NUf9XVXf61aTT<dB]fTDfBRD
=Q>>J2^PgK2D[=5R,XH&]^f<4ag&0OP70^(U.0f30[H[cWOgC3:e[c@M^NQJNTM1
S<a+K6a-@dUg5Od]Z#)M61QeG1K]7-)6baCYQNOT)_P)4:AOGC;,=W72OW2(a>:e
6,<2fgd,3(B;5NR##OP4L]G=4FO<S7P=[5T[&2^>C9XY;Q>CeD?a?(=gd_D+4\dK
O]Af,eg+^>c.S,YBO9SXPIJ;<WHCBIPY:2WUG@))7R_cgA3#OVX>R>WWa@?E5=Tg
>Qc)+#)]J1M0T=>+Z#8ZRXSBdZ7PT5+[fQ:bG((NW:/#0d4UTdK21]fbJ9@+S?_A
WNH/:NXX(-WR,BNA811<g&H4NP5N-9=4UE,:H?+g^4\G4T2ead98/SHHf4>LT(33
G^-L12YG5+HY@#H7#;?ZNC2C/5/A4/F97d+&0:)D0M5:+]<>;>Z6f6=I-V8SN6g<
,A+6f9-&:MU2R9X#A&Fe]?#?)2+14Ob1\14e4GV2Te],.^<NgRO&Ad[P)9[I_AfE
d&A2\H;XDEW)Q5[[\(W>3@JE9C2BOU(K6RWBCR>W=(Ic?b]gZE-.:AS>7J.6@1^[
4<d0)\6GF0?]PHQgZ#KV4;M3VY8>g@(fTD/VZQf9eRaJ+#V;e^Gfe]_I2ZDEB^2>
#g:c])7?b-Y]#S.B];<I5T]5cV\V<TTL;d\7_BZ^8\IGeDQd95U-aPG97=6E.gFX
(,K&FEMf\ed#RHJ7178,g3@FM6X@BG?+R\LC=#FY<,7U_,\Gd;CA&L/2;PPfR+^^
Z)[2S;;eG#B&82G#3>?LFVQOaWH3(9P\-T5+RcG&E<KcT/&I<&GM)Q;[[LdQb5;7
]3HC\aV[Q&4>;S<&-KJ2IQVdISH=,9;YcI7N3I8O&&Q@3DKe7/?/b8S<0L2OZ-,5
Pd/f(+K]V,FV?CYAT+I>HGC0][a;X#XGN7-VUUA^(NE9W?<[A0<L.CK@3cO/[./#
2;YJWA=X83V<R=XQ261_<SNf=2WW?L<OOZK-(ONT&0aQ\H;_/Q6.W2NS.CTWLL25
Bc2PLf67YVKSeDdUQg&>(]7b-dEcU?T:eTa?<HcKC\QXJ(T1F_eg8GE>8QH5;E7T
)Rg&DVI@MTJ2(8WeH\:+J+gL1&E0EMU9.^U2&:7:EF?.Fa/Gd[^CTG?[e[0(0Z=4
e^W>Z5+<YHD&<PD7S^d<5:9UeK=eW<0SJW?+YU,0+IWCE+M)U@]D0A8AZcR51_P-
&caS.H&KBE<X\[\c;A#a43#KP5/4H?J_V&[P0fB0[_4DJ#,WR(28a3P?&#8>-9U[
NSeb0A0C#9R/\fSP8#WNd0CS5J-/0Ha.2cG@A7.U1^OY(]1(PMPXI2_BVb-N@>.3
,O73L#QegJB_ZG?^B2K.gO5+=1(#G4a\AW]Q@M6,5(cC)\=E)P]GXR;=HCG9Q].G
IHW5.-/g.?AJf<eIFPNT_G&QLOM7C-X4-&+N5CaW?\R+W?&N[2gO&XP^H+c,LfZT
VU1#JSI&XKPW18I1RgSXeO:LKg;:<LHH4g/@,T49Z(#\GH61C1EHSRHB\?6JVYUP
QLHgcT8P]:=4CNH;eR,5WQQ/02a/Z>8[AaC&5<YX<ZC3@XGF24WD@EAG^e\R#F][
ASH;956>[9PCe+_#@/aTY1:aA]N_Z86TK.\CL,EdK[S:V-g,(5UKLU]UcSLP>J3P
EO^1CKZTU2@)fYR4g,Bb&6)#Kf^RAUHWT-]B@GYcWe.&@^Tg\0>EE=I9OJD4);5g
BbI\.:A8[5_?UL=/,D&I=^54KN1F+&5=VQIYU&D34Q&B\cTRIM@L1=87f\CSD)Z2
5/.#UN\0(1DaNB87McH@1@7fZ\7Ze8Q2KATDNXgK#UW:7He[V0b;4E-cFHg5UCT@
#FD]B.[3Ge(BQ---@C/7.10.?WNRB\RdM)H7YC;,.08:8A=ZWTYV=g)_==^=ZPf1
&>=SLZRd/E:0]VOS9<@:GOCME1,LBCKC.G<>OKC_BdFI&Z<FP?=ZbIb26S@>CHHS
F:eaHH<2eC(D=U#;+T2J&(?+aKb-:)CO]3>RONJY;+bb\LE2fMG1ed@WJDRegeJX
GD^c^WB.W\d,b7LG0BC2WSR78,4\IRdK_(?e&U3.GZd)_MBG8/DLeO7Z+]g>RHGR
df_F+-b8]\GYF.OQ3c/L,dCAQ(.@4b?5&YeAD5-2<56P9I:S1Z[KE_g(X@X_DVSJ
C:<IH6T5I-E,2CJO[^1G3P;E#(98A.//W]9MYQ(fKP[;335F,8B[EWa07Q7N6W=G
<&.<-YHZ,&4AV:JabeRbB0KKeY,5dB/a7eR&(T9P/]Z>B/?fLU#TGE/.\fBZV^Yb
8^4WQ@Y0M:4ba>U15YE_29g@Re[Z<V<^:C2OB55a+WTC\If=CX]1\:f?BeZ(gVFM
).<R]_dgI5aQMUaT8H/#&Xa[\THAf@65fX)f^0:Vdad?5E85L\d5ZMKU.5gQK@3/
:U1,Z?K.Y<\F.M@]RTg3P-UJM3NK9UI1A@Ed\5MK7aWQ]5_X32SI^G5LR?H\K(a=
9Q-BGYU0>RG^?JJ1JDe)(1#LL\E/3XNP@3XL<7J,4S#DA?QV-U)LR\0^BJBI61_C
KHAEI7H?F4)+?(Ia1K1V2c;a.c63b92GT\8](S5@gEcebH7=^IeI6EeHYYUBF])R
#(daKC.Vg#<Jg,b7F49e1A1H@W\\5=3-8Zg2g-A@HKZ==<YLbAU91T1N;9.#=C@D
fOUF90>4BKY=6_L7(=QWYg^Zf;/b5T3JgOFfK)6cGX].Q,d]=1f>/&0>D(T;B@FH
+H8UQLS_4FK5fP@aQIRVW=3KI4VM7S.6^P0f&VVc/-WO,G@H=#[/?W_K#VP8K@3T
Wg@;df13&(,bfO2G9?1MV\PP_PGP]J_f@5P.RC@C05\(AU[;+M(3(==<[@.(A1/<
d&1NRD99,@=:aOPD#XSa08]cSFDK.,FdCS--_+D[bc)9E,G[Jb819YFZNE832H9B
0Jc<Q?TXG68S,3C_+H:4X](;.9TZ.Gb6-V>,9LX4Fg^0XCHAGP\:CHE+BOW&,\>/
5IcN^P]gK@2f]>O.bUgR>;J\2;QG=G6&0-IY<aIgRSb59cQOBWOU[PIAJUJ5_Ua-
BK1O1b3AF,G+cKa=N(3+_KM(+R7BbA#-8\DTZV^4Y[]eH\)&Q6KL6fBUKRG5;f6c
g+U8fadKaLBS/RA_[TF=6Te5=ff><X.d:MdN]=_/&gUW28<Y02WX2P+1gU_>3a3P
KRK.;HFJIV#=R;f[1K[^X[O5]RUYOAF_=1M#&g<8\1MI9?<.Z;#?RSA:<9)(aH2Q
[KL9Y=-dQRDb:A>X[9R&SGG(<0+7O,>;F:cY63)@A(VZ/g?UeSeAT?->6R7SBC0K
0Y3Wg5;32LF3U@9__dEaHEcG1</_WT=X9QPbTP?ae5;^40CdbK7EO5N;30I?fIH1
ZU_Z_KHaY9JOZ+;-9#[F5_:ZF0;gQe53^D]8,K5DY+ZA0B94;DIO<gcPGc/WV<]0
R3[)=K?c:PeR65bG_RB@C(([TQaC>(d6:,AC3[VXN[A00QUUIc>5fDMf_a)6TEGD
9B5C5YZGdFW)8N4g&g5]7(AZ]V?S10eX480]9)RT_/L/2>YT1PcP1FeE?Z/K4]WY
=;adZcPNKK.MB-Bd-HD;I72[BE_78S&3R]F80L]#d,,OcLF_4F^,=RNcRPL]dL9]
UbVcN95:.4/TGAX1Xd:3:P(JVRc244HLDH9D2XOF,4g4D3-)6[B>P.MFK-Of-=g\
U]d#UTT7dPPHYPbg(f_L_@AF[&LLS\4Y?C,O\ACY)B:W;RPWS-(A8B#fF;0fKcbO
=B6H_+\BfBH<JNXgTA;VOY./0Q021^CN^5f=XX/,8IceQaD\0L^X?M6:#:L4V4Dc
KDT+5N0.HO9+UZI7S<DI,OUSW,Z@K:d9^A+;X/Z,]MDSM1d<E#27SXg^;3<R)XD&
&<]9M4X)L5aXT]+C5O?(-L7Y-AWSa_8JC92a@TUNY##?.eSKT-A(=e(dQ#\W<G#.
?RLaOY0HbU.aTJ#1-GeV9B7>H0bZU,._S\?d/J^U(.2NZ,.NKNTYXaP,C75Uc1CR
B(Wc5EHR4SKI.8b>[.3c(+.6F3GIMP_0&7.860OT:K4:\1&TCAID2]7)Bgd>1\B\
,.6Dg]2f,(FR41@4XZ\@)-BF/\YHV@6fFAH&X^OBG5]&fITOd>WR8OL\;^42)Yf=
aQ36PE2;(]?Pg>KG[3_F.A^KN4\N[5?c\ZAP4VMDc0NVE;b@+#FM-B?3491<S\3V
b)7[O:IE3K]CEJ.6^BZG]:6JfF)I=;S>HZa:Rege21=3U[MC(+F,gc1[(c=6VZH>
bB?NJ?bW1b5X0a[.[]COT)5Z3fDU0T#G4-Ua?&E//4?7-U96\?X^UCcB?^>3eN@J
(H98D2M4VPHRU]F^8e4AAT@C=+2L2VCg:DfTR3DbdS(0B:#T+Z&5&QF(A-)LPIWX
FHX^ED>^;9G^3913+JN-EB1;Jb411TWW^]f0ZV-BT)b>aCQJ0(I?d]FV5&6-J>1(
aAM;OS?P<8UY_=I]cR#-9N6d?(7K(#GNZ[_dfKK\2CC0T3_>@2eBP)W,=U67&5TS
-e\A-XCRB^I:SCdeVUAORA]X5HO]NDRVR2,&4M.fFVW,Z5]?Y0gOP7G\87V;(YNR
^3GDNe_9T;(a/.V(bKf7H:DVNL+L)?,g\]M9DLGHH7M1)[a+EH[S=Ha+&JE4WE,J
=->GcU_UUSE+H4[YF]T\f<LaSZH5aQG(Z[:Q69R8D=LfXQc..>8_#[U0O?,N,GI(
X4V0A-&Q&NM&/]5-/#=X^#=c>Z29;]-2Y[^@5Qa32.K2/dTXaTXDSBZb:)L8^)3g
@<A=AF)3.\/49,#ZXJ;7<)W58gFS-RDa\(eab.@7Xe;QQ))\a(7<6W@^BLXf0F@g
O\9J>4J4Z/A_7MOJFFU7-BcM\OF8C@S6?<Z4HS[;W68-6b59eg)dDH8V;??D6F_.
JM2/H?gVHQ5KWMb54J?J2Ya@?\/8.,cCELMM_N&OX9Y43;dV>^[=#N88)VfQXDHB
>>-RRdX>dQKJ7<C]=/TBa&KST5N5<fa<G;aJW3[3<88ZZ4H:G]L.>?CX14XP[cf6
(OJePN_]e?EUF#X/&)8R4YQ3I7;Z9S8.3D:IHcf9K18MD-G1,5(MY.5]LbOX<EA>
/NBSD64/Q:?C,X@C7#c4Y26:W+Xc4ZN:=[8FJ5-:/Q2PQ#X;fa+MJW8V5AO#H0X0
&e9F&:a3#.c4A+(V4,XI24ZT1,[Y8JI.JI3WTWeO#>N>IgOISI?J/^F-:T(BQ_Qb
fAa(Y.O10^\ADRg6#?I6^QVKFCG8;ZEOJQHCTZGL+#WE2FZ)g<d/[<KcQC/aXO45
XUYd-eXc)b3+TQQRBUE-5X+I(LB<1b#X6@N)I@5JKX2RY+Y2H:S\>(+IB+gaWP0\
L@2JK:2T6+R,e>AB5,>BD4OR<UE,[GH^g/2RNZM9YeJ&;/NODAM53[WYS2+O1F48
B-/7A3H(X(W,^@M,4?@e,dc#P-8Cb#FY-I4,]7[[WSgY;LMe#?OFNH\K?c2Z4U7W
gS>DD>1agg0A:QFEU5;\ED1RdHeATNdKBDd=e4cUUET4DJL7BJ2^X1c\dEL^\BZb
B2UfgDL04#QX,>c(.Of^T@Z&0@Hd>_,(RcgE&K@aG2f9d/#(/A[b):<9X;-9[W95
EQBB=GI,RBgTX=J=SbI+=&Q/WgV^G?#8,\2c,GA7]IWSgXDUCfWAf=;=4PL819GW
e;b(a#6:0_TebcSH<I2VFF7V8dVLEb>6-<C3;c6QHC/U>J^XS@MQXe4WRQSILC<=
QV]95R9+=73,Q<-FP\(U7^4=W\/6Q]4D?JC^\],9[U61WL37F:=A8;Y9gE2<2gLX
+\b2NX(SdK&E+aa<U-;3N3QKQc8H0<O01d2Mfd0J:IB.(ZJ60[]+TA=I]4a#]1?E
0]U<a^V9)#9(S/UWYd;I3>0_(-EL<82)e.ZURg93O&V?;E]51fN;>C<^/JaWS=D<
9R2FY)#]dAO;\f?2JST9ENcX)Gc1LZ.A@b1GPHaL7;]0V6,?T)8,@OW)QLZ.JI2Y
L594@?:g&d4H-CXacbZ9Ga/UbP=,[3E3<c,fQ)0PY>H6e[FXBK\82K=0d_R@D9+@
\FEWQ(UC#f](I<,R6TY&^.)92_MZMafUW@L]I4<&gUA)aLaeUDMAAgcG&<D9Ig[T
SDW_L^JP=C?:2OcN@>X<(cg?87WTCf9X52]?/_gC)f[1dT+KYWPL<1)T@5P3\ES]
(A5P:>0Y-_#IG<[;DRL;\?XKB&VZV-&4M4;P2e]>\65NW@F<&-0AaUJc+PU0M./-
)^\PGf>=MJc(eNB_c,M]L&&O4/fZT#SE<\-I]08?6FD.[b[KeI+O=<\7Y]+Be>_2
=A+ca.D:Q-gbd+aUTQ)B1^9.((;\Dc8TFY=,2+CW(:(2YED?b1]2c=<?d8#@<C]\
Z&8dLK1>]FU^5YV;)A9B4Z[<+]1P+_bAI>O[/RKP:,X/B3Y_b?;e<P[b(1J</gYJ
03MS/+[_gWP9<TMX;M[8;Ld>6K-MU7=KR8>9V^,0_[;YS=^9e11^--Q>OPF.SO^2
YJFRPeB(\@X]H#VGHFaB>WcNd5>5ONZY4?XT@dS]D?O;O=L,VD2[YY8V_:XMF/RM
G4L696Q?G7RdAagJP;DF8.G_HdFP82bcf4gCg#DP-^9daEOaeW;A5->V\K[UcJSE
RQ+62)Y4<]4^gE8bOD;JFE]J4GYeW._^.<RX+EM,e8Q01,.Q84,_@XR>=HeC4-d6
>#_XE?SNFRSJ#I:,U01P>?QTVWP/)fBH/R@?JBU1>5]YA?(_XMA.)1_cNOI,;^5D
T3[(\^^9OCJ9/5/;.;bL/=.7a@7)8Y1[6,<USg;.7RNGKU#]40B>DM<.HK]W:B&a
#Z[2;M+]>7L);dD[F+eEAc-eReW<+7f_OJ3G,,A9EdOe6N_QRZ+c+gWAcA+9=E>1
FMCW7>ZfF:[+FcWHf[eR3W_6KS7N]R0O2A#Fg+3J=c,PB?f&(J<(]g#C?<(8BNR+
_>Y@(D]O>,MKE?A;6P1.9B?MYT/M^#[e99XBCIeB0QY0c9DOKafPB7Hc-P_-Q+G;
<E?-4E:5b3aJ\21e]dM;(0Z.M)67HU[@.HOF^[[^)>^4IM3)3?G.--M-8A,+?3V6
_XDc]:.1Ie[Y?d1LW3^2;B4]_dEO]=bV,3+ZEPOY;T?.1DNW7[OYE\2fI_Q,(1QS
fc:P[]JbPfP,:T_bc\f8/AJU:;Y[?e.eGg(d.LB;6G5FNSG5>7a;<<VCRQ8,JLf7
Y&(A&)(Ped=&Ke?./:GX3>IVV7:(.MQ+dOL;RbP(2Q/L2]/6Y@dNWE)(?Jfc^N6D
bJR(YN8YOR@<Cd^DeB-X1&AIWW:MU91>\+d)J/(A;<9AQR]=fHY<X1eff]e^+9WP
>a@)(MScbO2>ILV14X\B]DRMEJ+-.83S\]4\1=]TcW.E>P7,17QX=.>DVLA\f9Rg
G\WU&6XRcR6=Vg5gAMK)Q><c3\[?I.LFVReM_2@6+&.5cN+9c#-.C)9,BTgX?GI&
H6\F42.a[6<eQ)aR&L&<G[:YFG9,H;=44U)G(efAFO:V.I]Dc(WI5\aV2e94(C@Z
[&TaWK_)/D\8F&>KG#KB@5c5ZSKONeWaU3fC7[@5ZRgeB[HR]c^B\e#dYHY56K0;
_D@51,90,CVLO7c.ALe3&O7_RP@^2.ccN=R&HcC-e&Y7R@?7^5-,^2XKeFK161I#
eR5fUT@?#+-P@=Xd)HOWXHXHM9^f+,HVUGUHgP/,48F+DXCeSH1DF@2cF82MU2V.
SaaMU2SPH97gc[)b:1ccVg3DdWa2)HPgI,#>U,4.\H[V2;5ZZGG^f.:A3;)K05-:
3(YQ6D^EF6Wg^[,5S5c&<CR5H48CZgI^&/Id0HEZA1FO^_L\3GI@<Z:M]Ja)3H&R
^-H:01;8P\MC,Wg>4gJbKF?CS&<+<4=aDPW,[9Y1S6,HF::cZO;1fA2?b2[8dQEa
\SJ\gScY_5HZ3S.B[707&EM2V9,C+5Bda>4gRVH77D&)V5[?NbH@NRa;?RPW__B)
>^FI9[QE-BQM)]3)/7ce354_/U,_5b6F\L-gSZLbZFROC+?9gaM>^I1-2YcSS,g&
GI^#+FVfQLK4.0(/SHfMO>^d8UQ<?>H6N2L>/UMWWe8VBAWI.0:U8(V<ZIN9bC-9
UG[f0cW4_M20@55E/Q)CGZ[SLK=INZWd?P?cb\X@EdCa_S-03]X<\/<VaP)H?-_8
H?>GJZO,0F_3a\WSPKXNSQbcdC.ZZ0IJddAJAEb;fF37;8:TJ(>OWI&^M.8Qe6=U
\0H8eGFU56)/ZA9=6V#R#XK]TaS;YJ,\YZd<a30+P&USa_NVT6?[a3e@d6QZ6;U)
^XMYL-;WXecXc=<\(@3@aHG[#:5/:4QQ>Pg9513O(?-6E-/eC8W2R5bKfV^0?]W;
/I/7Nc[_Ld8d<LVGOHZ#)S3>+Y,J]QW[P>=ZcRW\V\TK(B?;aM)(L0/44K9/P3_[
]#[H4,^:.GACVT;f]J1CIf,KC1TT3QLQII#e6-DV53-TY&04<<H5g:=d9O:=&+9?
DGPBVaGHf6/f@AT_S0TKS<&d0e5RAV])d<K6)IOG/&>e:J@(F(P7CXQ5K78&1B#Q
;\R=6<RODadGg(RA1))g74b?<#\C.eH7@D?K@faQUeXfX;R#;,[(IK@aRAA.0]+9
I/YHTdZ@F2;3&7)g>>BEE4&6),F\[D:H_Z9P9dR4W8WNX2:O#S+9)59)Y>BLAVXK
2F34(A+?6[XN@gc&d;)<YeP0?^;<6Jf7ga+MH(Lb)BG<^eP+)V+\1cWTGHa794A\
4_S79(V1,AGgON7L;+9F,YZf=D?RE0L.^)8UE\1AR7H>ZefO@e?P.\J^JS73O#5)
=-=gGdZdFTTOIW.KBS75+N=Y^8IF//XZ:O.eTYX)YY&KaS2CWFSMe+>TJ@Q<;Y#S
10Y:84@?A<6U,I73M3a2?0F^E>L;6]H?3YJ2HDY>-AA?+18N93LX1\8TDE.3X]MD
7H&^/SAAbDDf[:[V_Vf56aMBYaX2;8J2g34KFU-<Q&.Zd##E;[bV_W2>X8a[fS9^
]P55<Y4G)Ne^3N1GEdMLQD++GTU)g>TM^QFH@5]d7_d)6PKHZ46;-PW<]d]5ebaS
EaLI)W,a1ZTKOQ-\+TO1;V?PYVOT4aU[RS[EbA41A]eaQCKZ5;[GB.)BYdX>#93b
LL>1S0S\WCE1:5TF7?LO\BF6.AGA^0.^1^65C\LE[+/WcX)Y4a^BKVC/Zc+?,_4J
+Y3(M+eccYV;;B\-CH<YK7^d+QOHCP/9E[QK0BXZObEVR?UOHb=UH]93G#2WX^AA
U:)TUL[Y4b8O>@X(.^U4;V)A/LEU_U2d>:9c&=G3V@\.FZ@XcbdPUL<Z7C.@^H]&
N.N,Qb=a?_+S)d[\6gP8O::OD)LAH7N+4]<DCg]K4N#La;<(R98b<XGdfQGYY/7C
&#+ZJN[LWf/.0eR:a(?JN+6E\1LP(KVDfIQOK^3?:QMAa56>?EA6XH8#.1Q#(XL/
W@g-1MD@I;OCPSVgKUN?0;\e^aK&XDV=gK0PPN>&CX9fbO?I6Sg1aI@3^eCXQ&KX
N#PB^H2@N4<4^3B99?.-G6)0C#6+N1<CMY.g/K_IV>DgA1(^D95KLSB;:CC]VHeP
P,>8.:T9+c(?M_=4@SJ&/5G#&YUEGO)9OggHg-bX0f#R;(NLCXG9@?-XS8ZbWOKC
&Y,KA]\=gOMF]_5Z;S1I6L2PJO10)3=KJ5:GV4gKMB,X69.29a0/Ac^W1YHdKJ33
CdN<+;]L/;[FH&14I-D3UAe2&e#IT6\E[&P>DBFI+Qd&.^[1g+7CcYd&S?1D(d.X
9(1FL^af-cR^YB&@Ge3Oba6;g&SS#LdKPd/Uec=((U#:+X&93/Q;WFf,-c?_P\B-
e9^A+FN7YMd>?K&D-f_60EJMMbJ=84Y8W>;2CX9^d6CO?76M6cbb;35<>DaDCbd\
Pf1M@gALd3Q-,DP,B;gaf[^4IJX=Y>C/NK^S7FF?)[50J.dN9g)B@^]B:3P&K+(5
>EN?b1VQg\<F6B.LTZOG8c,5:#Q5A[bf=5Q-e58e3#.BSM95d_VY:;)#4CVSZ>5R
E+HMB@gc&faOe&ZY06LJSL&d_EV<,^46db#-/EV@_30D;6\B5V]Q<5<,ZSEU,H@V
f>W;@N,L<a)>,C=GWB7\a9d21g&3dZ;]6b/P^V0R8,;fOD-OZ6f#MD-A,[S:cKO?
If.Z=3N2?+6^bA+0<I.)L4_X0(g<W,&F3I@6?6^D_>SE45b3>G+(H<PA<9LT8\W:
B#@8USVI,-;_8=YW)=dV.[DI?B8S5C;J2Ed65VN]+W=[Wg2gTLgO6R7OK24]76bV
PXEfb(PSHRIO184(6IHX@LLI3#aIY(^E0<ON8@YY:\M26=O8V0/L-;;3)I6DG:HO
&)PaOY62[J5AGY@Qb?6]DPcdgX5[9_Y[J:7J9>..N:RA()ef+(\#5@:VM@(C81<7
1@:;XWV#O3B:XZ^>6bV(A_.=NXbDc0RO#_U8<U:5E.#YT8:>UC18PK8@^NR;RE?f
R@O2BSVU#S@I2SNV[7\2g<S\Mb<=Uf9;:1L94D:4268B]N6O]M4?<JY?Ve=EQFW9
9?e96R](QQ>L#M:NN-B,UcK:STd5;PNW7IN;+P1@C.WQO#1&[V7>#LPL6;fPIfDH
P@R]?gCX/Qb5HdP8L2g#JN\QF6O>NM2c:WM60FS39Rd?FD&TLeNLBB#Xf;VN7C]-
TJ\LS7g:efaDZO<3e<+J^></Y>:R@UE44a_-+D#e5b2IOG](KVa<;#6SVK=8H_B4
PQg_O]ZDM>:+-OWT6UKTMZJ\-X-]2I&\Y)P1I:.I5-#524gDI50,K@eI?-f&EKCI
N^e)OLI>UQ[/G--LeV.??CKe(3.5)adMZ&Z_AZ>2:]@K204)d1+Q&YD1AW);Y>UU
T<4S6LW,^Y;7A>3\FW8Gb=I)/62X/fD(N<@O:7H\6V\H:XWDHW,XMUMLL@Y5?AS0
De@W7:TLN-B)8(cY(J=RVc_36E/XB=+T=P8B,CA.J8X_75UMB4dH@;[(W3DWG=:b
4,d1OVAO>L8\=#\V?PO<0,/J>\QR#7FJ6^DO(F(VOTUcfPZO)5,L6(?T@>1Ya?2C
TE0JXZ<1]OEGF?:H,-SC?5_?b8AROVg5,aPKC.:dd=?L+ZA,DLG[K=FQB4&>g_5_
W:HIaWEE_QHcMe^K_Rc#Y+TO[R(LcgCS]KQ5IOGG5H-(#eRb\U0[;F[P@ZU,7aI/
Q#S_9E3A-WcS([..KOH+>WeVYJP0JX0)HgF0AN7@e1-ES\[1OSR:7XXTA+1,K?0a
Q9WTdFZ.4LS&,(Q<PV^Nb4(f708>M:GS_EG=::Hd4EI-1[U5W#P83;gIGE()>?SS
+R]KCTJbD<\f?(9&L5>X\0,bfG78IR8H\eM?HS-Tb0e+UO6U9fcZ35>b517C>U=F
T>,TP#RV:T>a?4J#Vg(cOELNGA0:B+-3&C]ea+.NW/1LSW_Z1Pg02_&C6@20S1;-
WBEe2O/)6L,B=B,]eN<?NagMN6U2gWBN6=gT,OGK?S?L9.73=:<@@/MAa/()?#=f
)We+Uc7I^.)6-4GS6#d.K+4_B9gSWH37=J6?;.FLPBA\B(]ML,[F]4I0,K>9ddH]
:Hf4\R8W4Jg3;WFI;0BYe4.Cb1caXS564\fSKSEF5RA;]>B(fd3IO99ZTg90C+>F
9]BbAYR+K(eg)8d5@4W]SU_DIRUHgd=OQU?:+OS:faBJBKI9aT)@3,/UgOIBO^b1
IH]V-;)^@ZbFLQV_FJfT9W36^1\@\#(2<cZ.GE=#Lc@0/;KAQBMU9Z<Y#:0A&dg]
DEb=EA_3fS7DBCc8N&LQBCP-+>GOVX;;1#d2\4?XU\)@I5-Ve=Pa-;^5)M(M2<V5
XE@WORW)RJ</ab6\2Z38^_][2Ma_<16L6]SK+Z6]-fc1.(8I?KN_M@])K/IS(ZP_
Yb_NHWQbZ[]DRZ)X8[?;RSg<,YGQf]6TCTPA4N6U5BaI(;7BF/6I&.,ODUI=8^,9
K7E)4Kd[V#J^:QN+8U2(d;dTC?PeegE81[\=2XP_K[g@);AS3I6RF/^^Ja5B-(L<
>M]#.G86D?>F+8g^@(QBSFZI0WEWV>Y#bZM6_CU?W;KVgN.OaGNcAF@gC,NJf,<)
K):\I95WDB=D2g,BJM<Hb983[,G:^TP]K_L&4>/dD\cO<ZL7V-S_.8;If4@8T4c-
_^eH\W8;GZ>[4N&eL^5-3+N4/4O^QUafTb-Z#IaA7DKcWX8<d;fISZ^H=.-7\+d_
^1QD_,=+^4aH^/:AO2NWF=bb\P3IXPQ3<7:DAN#d#&#?88.72=T9DVU^F0P4&D53
N<+&NATEWK@-DaR24gTCCA#:9Ta3d5-FK:Qb(eE6feY:[TX=>-V]\,HEOLW]d\Sg
U8gdag@ZW)#AGd&5V3KT[#5?.Te&&#C?^UG773.W?\NGS#P=&(2/MNWgVS&76D<@
,8(3=Lee3VgfD&]N.8Q98,S,g5RH?S+OM;IMb-Ud=fEUY3[WMR,++B(Q<6\Pb5G3
dHTc-4AXdb,TOP=8dI,&ab>_O15>F>BF8J>[HRX[8VRZ]40O^:=17X9Hg8f[,_GY
RED&\f;2-DXS5IWZQUX=[\VC&^2<3_Kf2df\Z_dc9Zd_-BAc8Na:TgbCFI(]C2JC
4=W?9aIO;5,Z2(EZ09<H?NI3__Pg\S#)_GF+/Bc7N>=1e/M8(1K,M@:agBA)HA+Z
_/Je0@0fF;2VCc>2?<6GM6Qb@L.eP&NLWfL@)M(Z?KB?/;PNc35)C29H=&gGg53R
##7dIDA>OeC+;bbTaeeT<@3Q.C;412^+:=)U@S-0gHAC5-9/f=?;[ZY107cM/@E>
O9R[][@3NF@ee@O>)#+0JK-FTV7G6X.OY#+>Z[XV->d^AC[E3Td\OO,IV+XZ+<Ke
dg&d8C<8fGQBBMDJ(,/JT_9<eR/P2T>.J=:B._:Pa5JJ8BEA46H/<#OWD64:,1[P
dMMQHFb?.ZGgFTK1Bf+_e[3;?(.6=+bO9;9afG-[I8/CKH4gXB@O4eOF1P&NeAI7
CDGg^(X=P>S(Y6E=[N;0Y6M7Mf+/CY06\,;Db70+OYOOXGU-_cPDHJ-SSAX>T\EG
IMK8fU3JEVb&N1F5e#4W?:[8TDI0FEcMAE[-,b(4[^P?IfG;3BgI/#?e2+SQ9\T\
YNL7V\L?8CAf/FXV(=8.SS4fg=TTdM]PFCIW[MO0b:2-,GD,01XJU5=9FREM&e:>
HLVU5-EXIU;^JC#8B8@7I)]DYO4I2b9]LM?>;J>9KY/]IR[O:EEZI82=+[ZI#Z?b
<CQS_KG-&LC7(QLD#>(2HKVO?EX_)@.=:M9G@=,4?[KQP#QEYB^MR5/3\6Z3&1^X
T-5.OP;7LX-5L.JIe7[N@^AM<LgU@_C_]2\_UL6?G&Lc[G^EY5DQ21^b&a,NL\J_
?#Q[\F)&X:Y2cUHWZFCN<EA1G-^>DT6_Y5,ffGcd3DI9:+@EYc7NICJa_,>=-Mb&
H15YFF/6c2gZOf&]1aU7JGQLGc<_R1C._82+YG1Q=g?:E4:@:L6Z#0]NX<JS#&7+
)f^7>^86EN;KVRUH4+6L;fWV\X(bH2WY[\RQ(N#][06GBVZg.(:0.UI[@N4WXH?S
9TRI@8\L.<DUT;S<I6Z:cHXX#<J4:agH+QDO9\JCOPX,SZI<GAF#)?Jd,,/OP>1O
W3D;GH4Ib[N^60a^:8I<G7P@.,_X:VX<(?cBb8ZeK=KZ4(<6ca\;D+LY?M\Ue3Y<
f??3)\M7KfV_ad-[F\[Od/K(66WU<X)^eVV&5,CIJ28fH@Z3U9LP4O-NK)?UU8[(
)6SREURa)>F>PP?2MRa>)?VY<P.bH5.;_83;7#OYPe<_.g=4?^6RGCEO=_;C5DgO
#P4[DNcT;Sg[WI:&Z.aVfe0S113aB>;AE;UQ53P;b,>XA]V_XC9]2:]#Y?(G<R+:
VC5G;XM[^W76S#3>JV>_ECIZQ8H]cROO&adM?N4P-VIFM#&(]D&03CTCdSDI_M.X
_GCYZORJVA\Z[4&&GQ.fEP;]MOb(7DF2V=ABJS_6JY:OGY)EcKENLZ4@?.Oc/.VC
UU:NT40<3HMNU,84?,O=.C6VRF0T6e5N1(aQ)\B7cDSBJYX?9<J(_72b)T>:\U2I
#M:?Q:K+]IQSH;7G6gWRV6VTF7EX-OZR7&&Q8]Z74H=;-U^3Q4_@g8AP.+BW.<N>
:1\2[fMK&aE7ABL;7/4/D^:2,<7)(@E:X_-YeSeZD9:8Na#F,1H?&F>K+JZWTA9R
X_8]bW9f(T==c>a(Qf/AE(7-G@OYGfWLd,+_Be?B1U0=F<]>Y,QK4gVC27K/)>bF
;68bc.Y,SGP@E7(/#g3US>,=,BX//3K9c:<:f;O.eC0+>=93TUW:fM]SGBf=#<1#
H(V<cf\B?PD3VXGb543UM<.>V)_fVdbO;1[7a5N=SE[AA7.OB=YaPPV[:@N0/8)@
)V>fPB+bRSDa?MB)GKCg=ULe@\DcOQL3)1P9PVKK67#WgDZ6T61K(AaIO7]18dGV
P?YZ;eM10:aD=ND@ZWBE42,f^_1Q+6:ac\/>X]cN0Gd<J:)L9>LFNI]1PPRHTBR5
H[NOcI/0V?#f1JW3:Ge,25]OMQUfQCP/W-C6FCeNAYG]=?G<QYWQ9&1X&KW[QV&,
aPSC?^QJ&/f+>-.QUJg@/EI#I]O@C3HU]9OD3/^bFCZ#D#)?N)<Q(G33FJ(Md=0Q
2aH<X9.05RYb-JdaS+_8eVC[Xg<OP<Ze>EIa&;X0+@R\1L8?C.S8K?a+<#IH]I,3
KFSH]DB^#1<,>XdW0ePZOf=,L9fUeITfHg8Qf692EfGaH+</YZBaKOVE3^Ig&_^O
V#HUA+;7a65YXg9WO26?=-L<:>C0LWa;;bP16/^>1BZX[Y7L(@e/9N-2ENPdCHdZ
R_\H]b92YA^B_2S10]JBK34dH+23e^.LM7?=@_5LQ6]TTF=V/b.I-N:a?;-+8eR1
^DW<6g7;0bN:PLWLf=PCUd@)TG[CQ?a/K(8W<fZNWg4>bO][TcH;SBfXO?F>O57P
@=SYB:WBD4I-R;8Z6_&>\/f-JN^ED]0(PZ0TI#_g-/.GH9/#B[YP4,(7DdcVG)8D
EIM0]8-#gGORd82F\fA@I9@H;<>>/?(b(@F>[VC0BI:_c4&1bA5^-8L/@;9:6;T)
#f##aT(GbY/+XAD_FN,XK-NK].XX3BV8G#VHX[II]A&2^RJE^98/b[7Sd=4]_?HO
2MUKcOfTA?6b]QKFKR^a9MTZW2R4]Y/@:ggNO=U--9V&SEZ<?1ZEQb2AE_@eEFKB
7&;=)Rc:0X\:3JGCL5gWaGT_(A5\D+\;^_6dA,^O5PZ4KEbYEbAW\KX8?W-O#F0_
LAL@ALBZD[.57Y(:8>Qf[OK&RSZ:0MD(@13&dS>OSICT=\CY(_;A+6,@#SO-e2K-
[/U]#LQ;:T[]e\KgS6b+63FL.[=J.+QV:_3L.Ce8N^O58OgV&0.UEB/27-]6]DL1
3\\,c:72ecICF#=6?g=X)NM2gLBI3JE-SJ:)P?FKaMZ)N6\aXG590/998P)9g\JR
@J0VHaXCRR[)2&XN(>X5?Hb@9(,CU/B&HUV\K6F4#&NS(PDR+_\B0e15/#6Z+UY7
J<McI.6MZ\baWH+cDCMeXWF8@8)egQB0??:XW6]HWPTJb<QY8^[9B]b4@Y(C@TB9
>DHNQNVZ_(SEQ@<-@>c@5I0\?V[P>U,X35&1?,&edKJE-aed6\BK,/>L5XdNQK73
/gf_FC7aYW2bcC1(&?gba;aXUT,P0+&:JMc(8=K;#_f9UJQ\/JL;T2Fa5)-^e1S.
7?Z(NcMgM@g3MHIP<=_<-aZ:BDfC4A::@5H>Gg40AOUT7@,E[e_)+NF?YdZIbgLY
KEQ<0I7.HVea64N)CUBH7)c>N-e)3-RO(P1Q]0_GCf/0<J<^^.Y)beEGHU9)BK;8
RWf6(WZL^JF(fC#\He8F>=.5LbIeI8P8Q7]9gbW2\(AEV4Xe[&_VUPARG5fQBFGG
TaD-JN^SZN0)d_[9]Y#5],8N+61J)J1T?3FEUUL29<R6;,FCOF>L)I3ZT;KJ)5#;
9L6:U&(KKZ)<\\d7K7)93dOMPXT;B;3S0L5fdAE+,4G5QEUaU;DG+P&[9\W2@@?[
<c804H?Z@-PGCIC[A-XERJUXM]VJDIUO&A?TFF2LL>KYR[BZ>B9SQ<2OMO6A0aM=
/.^YLY34X?La2/EK8UdF5J;^(EK0A>^VJ&N-H>9c2bI.:&JTL)?&)7eRMGH[&[6K
I)P#C<-4K>[fL^#>9=dOEAM\94R#,d[;F#LbfB5eZ<fV9HV(,.V_^\TF)>7fd2\(
<O,&-99@,KDO8ecdYC>+=X]WS2]V/N@OaQWc(QgO+1>5\<H6MFM=eYH/M&-)[O64
+T,G,L]:=IG@gH?O->AWK7]^Le.0Y9FU,O:#FNEV.5b4I\/&_>WSZ66e,3ZafM-.
c9(f:E63X2IX>Y1FaPQ3[-O[gQ<TgC<YK,dS6_X/5A\Wd7VcB21TO0fY&f6_^aAR
;]=aB^bAJIdA)eB\B6.K?A0dZ,CA,e_PdK,-&HMK(S95;/g+(=VI<A=<aN7+V=Gf
;^-J,/+S4X:ONHPI[ML3_D&F=MF37gNS]E4A:3;R\fAe7(G((>6@_,Z3^E1aeZ4b
BgaI[6<:=1>-;TZP?/_TYSU:I=>fbQY,R]UUPQgL?V[3L@PKC317af:[LX<^_^CJ
-+JcSAd\@=T&[g\^]94Lce4O7)K:PL6\E#4+b_K2\(42Xff;M[CA2Z]B7R@<,6.O
95.57eV=\2[gMX:+:\I>:aT#b(ZL07c9C<\+R7e\(@<JQ/BUW9[70KEF9(X[I5Qg
-MTd-(TgM)KM8&/c=b@5:U1aLF:7SYDJ+g]Y/T.PY3-VD3.U@M)DP-7/#aZUe3Ef
](JE9fA>P;7;AKQYDDadc;<MfK6S<e)?L&g4S3?@:d5ZE.W?[a/+C7B]32MccYQf
=#V??<c]3_P1;EDU\FZ&I_901H:9eFA=e=<d5E0/e-Yc^1]GK1MS2(CDd/f0RWXT
?K]S[UaB@QY,R2M8B-H4EH\(S_?1WO]5XTQOC,)d4-b#(,@&==2?\K]e@K[0S+D.
D-E5@#dM]QFGegA:8A@(&M&BY#CZR,E1(b7N>S0A-#JEX?5LD]P&W?U:<@6IW-^A
@T6,?BJgATc_P,dC.TWa&#d[^2WDP7[Z^gR/W8bYDVa/42J0&Ug/W^,#]ZFE[E+&
FFN8ge+NLKOYFC1LZ)eJcZ1cVDWd4U<?6R_#g&Z/]bRV;JIN]4CB>7B[_7&;.LUJ
BXbL<#^eQgH;.\PQ<T6^.C:[S>3&9gO^X=V5=K#:@_<bR(N2,D=ADUWNWOWd?C2&
/YR]\89]N3,d>LL/:QIL]\ZRD#Va]V;X?c)6_eH@=O728/1,1TO&X>>_=1E,(,=A
8e:Vbf7.K+,&BX@TD,3b,1D.3=XdRF@XQU[:<3WGJfS/F\<BN?:-._^MC)]CN+B#
YL07>B-RHGZAA.\?XFc[JD+?-gI;Pc,_O.82R(=1,K=?^B2OK+=FX[EM3\aCXDe=
2Y7L>FP@aPBARBJdJ3=f:]HHK:RUSW18#G\Y4:6P3XdVgcdJV&X_F:>RNHYgIMdU
D#E9I\<6_.,Y7(])Pg+/T87eT>LCgHg&TPFAYLYN.;I1HL08G<&bH)@1DA,:=O[e
I)aDM_2;3>)U;@UO79<aO(+DcUVFGAP)>5_,2#G_X]UU_=O[+//-OA3N]]/O)G.d
YPgg064AZ[1+-[.]S/9-RfX7bPZ_J9G71c>_]K:5LX.S)Va98e)HKP;RLX[OP6@K
X(.0Y4^55F]\74?GWbEUd[VFM\.6S),86FY==E)fLc9W1;F>YD_(fd,@<#_TL&@9
\375KGDEGF4<^aVYC/Le5>1F=bg.+ef.)T;NWA0(fVGVBQVO@N\:d9M[daY\@FUG
Qf_TG+7dd\D>-&U7N4RfEIDQdZ-M<E?,\[).A0b=X<TGKSKa9=g9.Y,#Uf-.adU?
>]V3,<&B2_@g8a6I#FLJXDNN(R,b_M,9P0eeO7)-9RY&L\\+f/(1C2AZ?)UF::EF
/9:Ja)?\FW4-E#0H)#M#[QM2F&+cY\I.Z68#g5Fb@cT4?e>UbXUG;/UfE,6eP^I)
-KbGL9Zb#;F47K@28S-,NVN]3FdaWK<\+PJbAOOeEAB\WZD/g+O(GL[TR,:.((NP
0@\\EV4A(QD\Pd),2B.g&X^U]JPUNOZ@Z9)^T#)DQY1LX5PG/Ug;S&8=:JAL_@O[
5[-GF\A_FcN4_d\5QHXg&-G02[E<JA.6#e[H.FP]2J=]_R,Od5C[K@?H/M.eJ&Zc
_b3^=/.Hcb0-eHd[)X5O<bAfTXcLZS;L?&_c)^M?5a.^66WXA()9/]fM5K49&4[#
LK@9N0C)JJJ,.^(N;D@;#GXc&41DgB_<[VJg4b3JXU0./9/,[MTAfB1\>=bMg8YZ
5=#.8Vd,RE#W;JE_d1fB1D-9)Gd<,Y?gV@eI@A)_]b>L5M\PJ(Nc/2N20d>9IE?I
XZC35T);PSg7AQVBEU@2K.[I.<4edTXRHa?D(L<ON1.5U#BVPNaZNL?6+)TbcV:c
YfBKc)L<aU5J;W;,U9fC=BC^c<AS#\53)O)#OQDN_Q646dI?]QfB2#6PGK)f<RWb
aK/Z7KR:9U0L8ZH;bHS45.:DgNMXa_cQI5ND\b7K0fJJ3L>AT#IZ5+f]3dPCA85.
_E<PN6C\=&]^--]+0V=K&J^>,>MOc@YNSXG-c8PK36a]9>9\[TcaABQ5@8)@E_Z1
T,((@e3;VFe&17]DD]:7Q(+F/8K2/&=\H6RLC;7:7NdYO&([KUB9.Xc7a(5USITP
8.>D&DaBe>16;f-Q#JEB<Q49NNb/[d<+,9gQCN=^<=Sf\O+_KB#[H^+:M&F\gGD-
2]]JF24^/EAOLR?5+]aP&YB7[:bDP<g>@6)RET@BH4cgGIZ^_7R\MKcAg[dU0LMf
b.DU85ZOeeCV]].+AcBcARU2YE,QHY+1OI1BA^C12EgD^R;0OJf;c3?b[aCYY]<d
0]Sg=7fHd1PPHd3?<bH-#W&9e8<YMD&8DF5&OKU;=92B@.GJ,-_M/_:--L^/C,T#
R<&H-U,R;.G&AMB#^DdS>?::87c+KS]ZeE>QdK]9T+SEVLJUNOH2Z+/RAd)C@E?M
-W])0Qb\UL:0/)/:&8<V:ZTU2ba>3,D#K1C=7<U<QV6Ub@Q>9EaM-IH<<g5T?G=H
[WEEUGQ(PQYKOfZ\;H^S.0M;@bE=TG/V@1WaZYfL,a-=P&KB3W.2<8c8_9KG/LQM
>TG.M/:K@79c/&L471-:\d;C^[VQZeO6dRCaXWcc;QEY/[BX92,R\#Ba3N)dcI15
_KfJ\>@=]/<aINR-Gb?)-I5YNdYc#.-P[ee[@7LKC],]TPD(;^Y?+>cf>\9?N?@O
D3IRHBVT5_(Wc\Y/KEfRWRS]3[QE#^D\af<X9&V+.&)Q\+(G4-3fdN^LU^?G1Ge6
/WBG6[.N9-WPT#S)Yg54B\POP+]:3O+BZSUG:27fHTNV(C_KbE2d9d#b(-D9[2gD
a;J<NIVHa:51M5#TBgILeX@Ib7f_CG89\&8@R-8)c9_cTLA7VR>(F2D<HQE,&\U^
e(a5<J9U.2UM:-]aHKN=/c1c8O3_(e84IZUWgG#A6/)H#.X/@[,MH+[?;Z\8N./R
HMD=/J&f6_F#NJ9U6P71I_-H9>YQVff^74aIWGbT.2dP6Q1TJCQYVVFLdJC3YgH?
=VJKab=UX>1J<_[WN=_^0-ML2BfNZ,AFJ:#D@P;e::-L1S.U[DDVX6=NF#URM-;F
R#U:@6(A5fU1b+Wffe(2L)<8#_LbFLcb_BDSd?GWdS@AP2D.SAbP52@CR3A5K)M]
bNfR1Je/^IMICR6YSNH0A_[LQ]LW:[PgE8_BTP4PJY.LOd8)a)>>dg@JG+UOG];7
OKb/Y[D,W:^?A^cN9W+B6;CU,]9R4)JXaFEfW5@\8T=YEWWgD64X(0;T2\ZXGM7N
,MD]1)C169D<7;da_(?+AcV/?#6MePgBbE7+B8C<F,34C_::)U:B/P/5e?GXRDF)
X#DS]#W-.I=P4=.2OU?A);Se)M^H]B)cZPRR^^#B+R/1@4-S>+R<cOK94Ag/.MH[
]fB0<NS5TT3f9Mb/.W9/4[8)c>DA]S;Q2bG;,e-R07S>I_^JH6gfUP+7PVXaHR;F
)+?3/H-/:E.&UIPgcf/Z[D9RD+^VUgT8;AZ+Y&>B?OU\gfSL=2T7-E&]<_YQJ/>8
Q+\EN6-^?\HC6WO,ZbG9+dg.7V?AJ>L14PM)(3f]#&<&BSUM,E0QH4^5\b>4C4_c
L>++fKc,::W9fKA2[+2]NN:Q2W@UfbN5,Q]gMGBbcPKcRW-5GICaXCGad@8GT38-
)I9HV_8>KM@MU&V&XXfRHFg</[<fVT,Q:67W1fc<\Q&8aN;>6X6GBKAWHUYXBc&b
QUFLBL7/>VD^aO00B>,L4<Z@NebQ[PGJ=?P-b7ddP>ONA/SW0Kd@b[dF5JO#8ce]
gVI<68+Pe?(KGGF3MW^c?9#;,EdZ:^eAI9dY&\#8KN=V^ER-H#:6MA0:PR+0P9e;
OI^&@<__54G+^Z&2N\O\^9fNM4f1C_HVPFF\QLB(J0QFcb>:Ud:d[#SS(:AY:.;O
/V[M5P>/^K]aOO6(SZDTEOHCZaD4R2dgR[<Q]>>YNZ)ae]NA:N4c4?ZZ<OU<I)&F
6dD:S,?0/DK,6LcdJB(cD8[JFbdc5UM.5(1Nc[=+-+0B]fb:/<;OOB\;Mf0+.WFO
@E#8Ue-B2.0,OcgY76T-O&6#,;>,:9:5-U_:,1YeN):-O6RJ8)^(YHK4>AEW(R-@
6-V^88;^Je8Z25)=J8]?:C,adV1V[aPe=W#I<Mbf13S:;H24_d>W@bN_gXWVASK+
_X#SCg+=6?gMH4AW>bV3eX>B1KC6,A[J+KCcVS>X-+MV<V/I8>QL_N7d5S72Z7J+
M>dcJRD?5FR8gYSS>RXD=(gQGI6PdM?\15B=[?&I8(U=_?]Y[C2IA(1SLB6>LPPA
BJ9)Mg435A-V[X4C[,GFDQDC+6B^^HV8e:5Q60_#^LSa,OJ1;;2HbVH58)c2H.Q.
fWL:1(1U+NI:/fBMQfdVR[)M+,J/DeAC\I\N.10TG14>_=R#00N@38F#MO.(g?AH
Bbfg6TP#2&+Q<D9TB+E0Kfde#GKG71@Jb7B_<9EM6W50?c@A6e;2?4/C]]7M474E
e\@^Ca3L,K3CKVeb^&,g)7BV7YHVY[,]-J4KaX(W7T9K]\ZH;D+b:Q2?.<D0DcQ1
=.,L]]C3TeaN<_YJ?W[R[DJ,b61K,6F&KNN=Y_3K-,F\?SWKQ3-Y9ZH0HUMLdf-b
F?D4+FOg:Pc]E1+f?EdZda\J[1T+d?5:+@FbcgO\3@c#<]S?R0VUZf_0aY14HH,g
d8-RGS<:b7#GL^D]43g@=OHE#@B)SH0/PQP1/9UbT&JQY[2UUf9N+L;8ZT>2Q;C^
E07^7116Z4B#IGI-F-82=WDPE4Eb)Y,\Pe1NNUIP&M,.LM<D#,N(18C#bFR8T8.?
eP&E]I2C,:C\_)f+@[Fb)=XS<Q,<4<_@HH/4&8+d6G04BPDL#-G(@LIID^^5LVF5
_RaGD)CF<aNbL8#<3(@74TF4Z@G2<DAFH,?8Cd^-Z)T^]JW+39&E[d[ESQ.^L/@T
<WV\L[6M4[La;RHX=?:H.Vf.GF7Se8f:_>PWYJfM8XKO-3J,]aVR;[?R:F+<g5+M
bY)<a((OG7S/X_P_RF8&/[P^P4V9bF(-Lb&H(.,40B8):F:E.B\Q:aSYM5DcP;&\
99/_?E_F)Obd;]WX.VXfGNNd&]d]egfd-.\3-^a+72NKU+LP2F^R@8Q5W=VR9MUY
g>,KBJ8b3f^AbM8,-\:@L&T;YP5:#/L;0(gT79U+_LP-L,T4Hd\V#F:W:G+@e:a0
OE]E=TTYP:b&YGa]D@R7PdQ?KX,;1eU/Ea#PVfVDdJ(?I&gWC7P5IKAda]+&_C<]
bAO@4^&g7G71XFK63+M]TbP@Z?ecU(f@SeDfg;,3@NKb()^-;AdYa2ZS4DHMEO,K
N,bNK3eED;:2MVABY;\&M3H1?/Mf/HXL;H5+C^IGZX_P1c<3@[A7(d;FZ5@Vg;V2
bMLUEbTbRgC:\T:I^a/\,B[2(C?H-bWeA?^DCH]LPJMK0cN&9QK\ET+G@,.f<81W
W,^3IPT-&BKJI=-4cH#NYCD-Z,B?Pa4,0YD@@VR>Mb,.7K)\+5=L[J@;]<+9VFfZ
(KaJ-NQ^]QJEMVA_bb_TQbM3Zd4_Wf\UQ;B\dZ:MeJ]Pa,ZAOOXOCI6)G(,:&ce5
Y158:Xb,Q+0H0\IL_P+(&dA65^JLdUZ6=1&50EgT6WO(JB0=+]ZWg0]@&6cPM8^D
+^Fa)43.SeWNGaR[LfPQaRX.+0(3:XHg[D8TWA(21D^b]R0aM;W.d8gC@_abfI>W
R>GCc3V>cg7)/#Q<Z;<8d]^&QX(,f)PGFT)@5g<,&^FCKMaTQKYeF?>DGb2?#<2)
>TSGZ2,e5L1H)4J?N>f#=[I#>gQDe&AMCE6BE8\6RfZ7d73aHcaKGd1NX1JeL=_6
CeRddVI;KA9?+;(-I=3AU5@I2I4c_LHI16&0ZD=YNag?>72]c[P12Zf&P5BB+G&Q
\7(2C&X)57PN#;Z?W41cJ&#&28<XgNfYTJ4AT5gSS1()JO#W2g(Y>\b63_9bPAVF
II[,<ST>)(_4+229(MP\\6HD@V74L;1R9H;O&)3_gR+2=f(+:83PTZ?-b=QK6S+V
N;e_4@S15-1.RY=9D?&L;P]A+=DePZg?\WH>fOdC[Ob2-M?dAK7)6@D?b4:d#>>Y
#M)SB2UE<VOf383@^V=J+0NQg]+83M]gSW,#5D)5Y^=O<#0cELXFVe5V/0^DNVS5
(KZ(^Bf97O>>U::9e),/T[^T3A[(8970X\.L_WG9V,TV:L5U;O,a;JA)8YZ[26_3
;,1e:#SR).W742YcX:Ig6T<H#gLN(<dCRD)^B9[TGAfD>f]5^6f(FDH=fS2^C.be
P92g/434EdHH]S+I#48e_g&P80Bc<]JS#@6Q&296P:f0?;S=8+1V]7K))9D=QH3H
<04N@#&;I@^Y<V<B@K7SESZI37_.1LE\g.\^?a.>@@[S_H?g_=\(dKIRZCI_?;:K
RXGW/E;QW7J2dE4T#g@R0L>?SGA99<Q4b?AP74?dP5M3Kf<CX@JSHP\YF>0_17@N
3I6>a[_/G.D#Ob8_:G8FF3_PIR-fY(6.<d/b<HI(gV07B6VDM;:\6G-?WW]>RX[5
<X)4e.V(bTbL8G(S3b2OPB)]N62bR;ZBUd/V[LbUbSfJKNSLUGD4a2=/_McdGD.g
?V)TY#bdWV;3GCQ./TDYKKI1F)&Y-\]?+-B]>VB0ggVQ(]eG2g=Ifc[,4?cF+N@C
;Qf<??b/--BMYbN<b.?>RU+b?2JV8-cXPP._X4\MF;>b^A<QB&;=]49ZC4I)D],0
A:ENXE1->@g;2OBgXANeE2#(WP2(9>fV+WZL^de3P]5A&PeSAC=\^GM,4,15S635
f,X:K7>fc.(K4&(P&_B+CJM#YU0T33P^W(6_fca0U=VBb&N=b@#c3.6]73E?KJ3d
:/FfEOZYacYSF3eF&)-Oa;.ZA[#@ZLJU/Xba3,5[Q:-:U7^PW_-SVD=+@Re55M)+
IVFY]g]GI#Y0S21e^OKa3T;NLWW0AJSM4a-6\\B;XD^3+bZR3?a&YcROJ#R0NcAB
739+F^GH=+dfU]M.Y55:)\YZLD#[e_?U;c1d?\Z&c-\f:LHQ0caYGd9:Db-cd9>e
cAG350E)T2T/T4S.7AY6[OZ[DKVFb&]R+=>0JZ@gIY2&6c)>,1f2?Ob0_OS+_8AL
V#2W5)#[U?g]1X;,R?-ENPN85PP&<gJYa?.7U=Y(Z\4b9Q,B6e/AUgY,=1PbWH)&
I;\#e[gPeOR:e-[P3C2A+5-N<PIM-)TZJSJ^;fL:?P#dW[I1FX@9ZANBf2XZJ?D;
5,A8E&B+;HZI/E[Lg4QH]OZ9EFFYDYA4I6C0XUWc:f4OLC+]B]K7e;)ZG(bS])U)
e@C:V[DfQ6137@#e:g_ALOPUOg&291X]C0SVS,N/F?W]C45Ga0bPbYAUV57(K.+>
M8WN3g&-Zd1:Q[SELgQX^8.FDQ]XgIP<EKRL4V@e2d<WQGA6<>?f(M+ET3;bNRBe
g^Q^;g^JBLRQ9LZE\4^1TNQ2X8fU]#8dZ;Cf.f+&LJB)2eQA;6RAL-L8fW4EK792
I0:MCSI+]1U;(:=f)d:e-KOR<KEP:,Vb@dNaI;LDB-a.MWVbIY?^ER70e_URc4Ie
b]]1([K?_4R,B-G4gbR[EFa\OaRGBD<a:EZ-0EaIC2&YTY[5?<9_WA^Z-](da,>)
^3GQ/CHOZ=dd]2KQJ1]2,c,=KOT/=1N-G<;MCP@+eObcACgHKa+9UE>OTf\gJ7Y[
6R)&,2F4I3Qb9O>6ZGR(c&<\FZDWLBBCBN<U8Z.V+-,=,&gPW.N>LcPFWWB-Qd#C
;XUC3F08L<9cW[A4cc02G3M>Q7G_FW3,U.#B2,/f+KX037M/g/d=[4J+IJ@???7?
5=L-E9K?1Nf0B>H)N\]&d.c-Z)_164>M\FQF_/(\0M&)bCP?RWb\/7\aQK7G@N/<
?7J,M\C0ETF51]G=4W:55M.5,6\-0N?0A02X(aJM\&(TdAQN(GN0HSeY<P\+<@D]
[L5ZAJ=HGP425DcNK)U2]:J#D/B+aBRKLcaII?W^3;F9S(Tc+F7JCLSF].2-\g80
#E?AfYI&^93:9Q#G<635-,e_K5E:gU4DcX_d[UB-QY?6#.;^<Q+\C4PND6(@R.95
FL-ReX6E@Q\cRA?.S;:TO4/X?C40bOUg4N;\Y(I)-/EbVAUWadcfT>7WR3LQ1Lad
/FaTO7-IKVa92>@Y[)FLWE_BCCCD5aJ)/LWb_X.]5b-gV9,?SO5@2NgENX,c.?/5
g)KTeI^/._IVWID_X,Ge;R?@FVPULX\1:JEb^aZf/^c0FW]ALA)\R.0W]6#A.R_W
\)#;Q0C?fVO.ZAb/3W6b#[KK_RRZUcT&RC@N&9Me7Jd=0;XeF[H+O8BE3O-/Z28O
LdM]197#.G=N8(1BTADeR:g-+OMSBUIZ(Nd60Da>/VcHVA8_8#R6W+aJ/RTY(+05
L2Vb;>0FUS>;)]GGG?<I6G+aaXYTc&-XI.Z)/gJf&P9M04)S+a8^:eSDc_<I8<5>
?0J]LP1A)U+Y4<C>RedHW]^X33J<;#C[b#G=5a-,8M7P,M_bQg,S,+\g-W>C?f+a
632Z5<>^,))N+I[PL=\L0aeaU/O,ML(5_dVO0=.).6-S.N-QFW[6?VK?Q8FU<fL/
O_<LTB>B<V82O+,cM>b)I[,N@JY<MT.#=GR,e^(]a[gHL:E=7(&0J(fN>ScB5DDW
&/.G^1;&P#Xg>1\8BIR(WMXE[bC;TWeDE65_EU6W#AAKNc<9#MeF]NAc6TA#9>;a
J6e@X?--g;WSOa^CSBS7NPg@GCIb,X+A9@V,0+S4[:a:H]P&KBR=)O+/.Y=^1Hf?
KgaeI7#4ef<Q4OFfG6#/XgA#KMa#F#O/c8<bGPI-2=28B5<KX<_4\S>+K:AIAV8-
L9a8T6T<?T8(6;6NM0]+?/]ZYQ_&8CRS>f(QFT(P5QCFD+?M^;G6<\_<W5^4D@]&
LHdLWFT.)AH(\/agbYVAO;C(Q^YAI/W4gCOBd6gP0=-N0aQ?TR=1=8ST\@2VU;1e
WK.LeZ])L-9QO5RCLU)=g=_Re4-/IdH<fCXc;.-/#9S]X#,5L0]7f<0GRR,LTP<X
gHR1NY1Q)AN5M_fX_H[<.=L=2WgH]I^C#+@243#\+A_c#>B_))B/+QR/1#b;EI>7
(F;YR(XULbM4c_=_F.0B@G9cZd6(1.W:6a]-Y#PVAQCQ,BdQ07KgJSa1W+ZYF(Y.
aV1aI/PO:&D7c>d)>K9ZHb\@M7V04K93AebeE)LHP<5(OXOAIT__+FNGOO(I@b&.
e?AUQ5<CD]L@#P4&d#(5):X/JXCCK/>.R1<XFeAJ88)1cI[P<7d-RJ,+4LCDfQ_/
AX>bcN370[??Kg:a3<<M&ZF6<_UU9QaG7_=B;&B@P\4?a\;\^7_<K..9ISB=LL-1
<6FJST2NXP+Ga,-OO4&^4_F:D^Wb<e26H4QRbX]9f,NSb])gSW@FM4Q7X5,XAV3W
PN-P1JHH7LLSfURQ>H3^J?f)(KEE#Zc_dH)XaB-GZ<fMD6\dLCEP<7I__@a+Xa\:
,FOBPKAGLD@]X<gOQY13^XJ#?)Kg=Y2EECL\T?dR7CB9DV&<eRc4ASSSH@9]T<D@
2G4^SPM\Vg6QX_^P0W)(?Ma]bHUW)GSHb[_eE[c)F>/c4Ce)VY7-,I6(H6eH.QEG
O?RTI9ge7O4PRRX94UPM6C4]1J&b^+[fZc5aQXf?gVY(:baPH>dd6WKXB\50=XVe
A)&S]-QX3#4,?#>?cIN:ZK&C7A2+H^Bc^(B6#CIHAUNI0IUIgK[aTW,[C1dC36Ie
K;HYYZQKaOY5f_c9Y312:2O<DZ/gOfURM,=#/cJ8X6.F>074C,89^W<958D+Dga<
Va[&YTcN1;2GGBac0UI/.SW?2\#\BJ>Q^R]IL=d;GR3U<_G:K-C:/7cB65HZK1:;
U<0L?[<ISMFG&\6\5=\-5OPE7PSN3W<\@Ub//FF<BWGNHEW<3]P]L=V;JW/0cGc/
#0Qeg_1C1K0MTa(W/\RBG;\_Pe7581.Vb4H:bF/J&F<c1:1]IKP]B(C]:61SLPH>
e6d?X:L=W8-+F;=6_G5.&C[If/G(&ePdH:ZF^K[bV3&[(P4._27>:[JM#1Ya@85e
Sf0bL@@0]4CVdXcR:?Da-?U:gX1EMG:RKM/b9-N&C\^4<Ub[6J5RPQW@XTD4dRAf
fC7PMNdKU472\B^3\G)a35_aS;YeL0V>#,@eAO0OH#;7b[RKG;T0R4G=aRTPM4J)
V).FGY1<&NCI/B;-dPZYYH-AUdS4HZ2_,/C+YE._C]A\<R9H1I#+U&<6^Z3dJR\=
.]S3g\gOKfTST092ZIA89TF,K.(#I]6U=T1a#I=,L1VaWa0SZ(09M]M5/11>7T9C
e1&8bd:YALCRZZ<T9I090dF_#/Ug]&[GN)R>F,eXNO1)7CM_,L0c[[850G6^:VY\
>L1AWTY-@9N=HJGS;?dFK8f,;[:9HfSZAO8ebgQgZ@XEWdCO-65Z4K;7I[.VSfMQ
K9.CCW7BRL<,6NKeIP9AUg3g8[W<QMfcG1dg3AXHa1FJW]INN67^6UU4R6^]J0VD
VNb+cUQ+Lc()>OPX^fE4#O-5RZ#b1904ZKeB4AS&7NS&GY;49\CbA-8&BU@];49T
N/9[LE@AQU]YWa3L)RYFNcCe[Dg7VgM&f:K(d>4KR.M0+f?K)Z2:g#bH[Z8FV2-b
>dWC1fGcFKP)OXBW8=MITC;VOEGWDb<^/G<W#C-+[=c^3,74H4B=D][.GO^[@YeS
1W;[Uf,eA?W]&cF)ECT4^Ng-NJUM_B<f,b/;U;1;3R.-DaES,_-W1GOb3fF<=H0U
:R^JP[:&V[G(&T38?KD[]UOZ;RR@f_O=T;XPH=#SP5M_@e&BPfIT#>KB9O&+Y-P5
:8:>C4[gN(&A)+a,JZ.NVeZ(YS6B.dQV6X#BBV^>(24+dL?><DF&dEE8fEH]VFU=
W9=O[5UXXKZ-U:ZW]ZCHaR7=5Ga@a]_<E5fWL3M,D,U2g6D(P3^A>2=:#,.LI+,f
]99\aC[Q&QA&HD[:;]5.ZVggAa3:NMRT>-AfHO2g9(>RQFN/X,:^I.;2QXE6\=7a
;aX4:F(_RV90aH9VS/PA3c+Z5Qbb7@MGI0YDI7I>L5UAA)IP]8&]1Z1,2_NdeV;;
D@<(9Ce;KbR/U,M5(9^Y&O0[^\4_RNR@)eAI8MHB8_&C6BZSY8BG&1S/U1&U2TS1
?AUY\I)]#,SMQfbI<#KV3ef9GL/LKfF3_6>]D.R8bV_dTf3P;S/&N=U<Mc+a6_P,
SATV3V==Q;YFWVfO(0JU2<BC^BLA3)56/dQe9GHO&4I&]gHb88,/K6K?ZT&e76#K
NY.V\0Ag(A#NXX7;f4BcJ,66+.NSG0-bS&N)?A#)34_dCg+2.QNYB[]5I/#g+eQc
L:T5_).#PJ6/g=DdT@T8Nc;K4UBO2P?=N7<.EL^-4-79>?[2T(YS8b\K\QcHY[O4
FP>^RR.<Kd,eG7C+V&SB\PIIY3Qa>Q<-8P44a6P(O;R)beD30e]4MJ\AJJZPY9+_
BTa4G^4718LGd2WRF7M>fQHLY/=WOBS<?f-A>,2M:#29ZBQ_1c;E::B;ZU6-2#DW
21Ad=>:V/GRd.G;aCf?2>.3I[geQ:W^799=G#^Da==ba0GXc/?+Q(O_PfJ.B9KMA
?CbeF_V4=VW+1OPG&)UcZ:^.6D8OE7,BX;9cT4[d[P(:CWHWO;:)Q>9>D>BNQ?TI
,;93.Rbg?H#<>U>Xe(<#VgJ,(g-=;XO0Ig3g-Id.c,;/1QSTD(>)bdVd#,S&?=WZ
Mg7V)Uf[222a&W/M-N=@I[:BaYNUMH/eF>dRRET]-R8-9[,fC?[RF1M41=D[1SQ;
4FI5@Q#9c)@O@RFQ_03DE;\BWIN2.9QUH[]&R.c\8E^c9?WAF[O#HY],:3\.Z1d0
R+#gNRUeUEa^34T9>9B9GZe4H0EZNRTBeW3UZRG-)(g3g)/66>):f]MXGU,8:d5A
b=ZX+&-6=Y]?;(LZa_.gPaJK;#DHC1SOaUd]eMX_Y^UQ8FF9_/WI&E1YA9B<>\TY
=#bLT-,+_TfN@I^)aQ2&JY=8SKR3BPg@>V#S<@8b(#L=;=SaT-&\V-+=1<]UP.N4
<9G(<84SOX/EWV)_WY-4>V7PPPc77F9K^Y24?Oe8C[723WO,BDR<::,19SC\Xd5.
#VG=54JJ\Ze6M^C<@WI7ffbe7U@?9.JgMHJeTN^/Ub_/cD&3EIILDaE@EJ,<1&HI
\8MKGc6\E8&W[Ad]6f4f)aC#X-OJgKRT2L:KcU6XX?J1_6,eP^.AU8BGVY5WVaaI
#1fH&a#.JIN.UHS55OVZM:^&JfU.?,/GaP.d0HfEN(-<CM[Y2aS3c1eE@]H-KNbb
RQ?CKGQ;,+:6YIDUG6,M.+ZSP]W)QYA\@.eO]/^I@SXK^5CCVMb@5W.LVf.HO\^c
\U_EI=Q_fW7WaQec=7SJCFM#<WWc#<b\_@\7_0;M_MZK8U6?6Cc9Mb8PYd6B55U^
K>0eTEE9SZ]&ZLRTVW;T5P:^]X?/H)=3\RDJ(>>2Ib.=U^^W3VLd26>)I_HZE\QE
R=RcS>UC>-FdPRNH[UM6A^D/KKIA/ANJ9/8deO?IL)D07GQ]L^b(P[4L;>.b9_bV
PG>JJcOe=DI_bacI;<K(TB?<1G^&XJE^#b1+OV5>dKd^48WFc.1GXbcETd+9BR=a
NKU_X7.,37O&2^]#F81,8:B2.6gAeJGZ@W8Ze-1_JcJ#.)^EE+eRT/QK,^Z/:A2R
JTRMUfP#UT.K+CP4(@eX,bc:HTOZ.EUL8^T3RCSP#:.>e)5W<\2YW/KT/VAGWE0>
E<CK5M;MD)\FB8A^S(ME1Hb3d8[gTT_2[B6DVD<99([aTRgd_cYT:6;ROAWd?Sec
b+@P[CMPOH5B;MN=7@:gDXH#UW4RBFLXPH8A#RSP]Y1:KN]c<?M+7NYP;RggR)a)
Qe8KaGD2e?S]6\SA4XW]6T]eZ?M_RURQC^gJdPafV7VM-O^eSfa?1U.GG0L_+SII
&50JKD4DYEHNE2#(0g_9^N.IE\CA@8W&:aE.:ASF.\\MF$
`endprotected

`protected
0,4,c1Q7QAB?17;0)^>cPV=+A?E[)259FeJR],f<B1TH9.O,>C.G,)\X1^R.7Y@B
C1E\A;UH]XY?+$
`endprotected

//vcs_lic_vip_protect
  `protected
2;NJX\=7-0HNOHbKE[+bdcB)W-YNUIHCb8>-5>.EYXbXMI^e>>F_)(\[R]O](XJ8
K=W,2cCS1XYJB#1=9cX]W,^I#]7ER\f8)_@?c?<g-AHT#JQKN1a[1G-]24\]ggNH
+fKYG[^:DQLgC^Y73184gZ]RS8Vbf?G><19VZS36Wed>c8>J71G(U7IZDKf/-@BJ
B0+/2#ga/]N+<)YOLM@LT8#&FBK1@]]?R#/C580:AS-6:>Pb>-<(e+MD\>T),9<R
F2Y]<H,Z,BWRV8F4=K-YdPJ@1R+3.Y@#a<4/:8L,eOe<2G^>GG)a=P3F_MWQY5?9
TCO<H^-O_CIS5GK+Q>1B,5SF<0Y=9FY&0e6gaP+9>bR5;>ON.5O&\]M#\ST65Xea
_RE6Xg[8d+V3?a6\\@G1:fW8g.DIUb^8VO^Z3,[>Y@dS4X7#R243e>[b<=)HY3A]
e>fYc<2c3/9cG4N19L<4X(.6=5]N((JCc>X\TLdS[dNdJc^S@^2)I8NQfB4VI8RO
Z&;1>8Z>>J25DS\]d=4O335f+Y]g:T&LWKE@-3)eX2GY?4AMVGTQ(VcK;[,HTT]/
&<c@YK^L4.?e^WX;=]^X)3YD/L)c0.0F<#JSIFZG8I_R8eSU(YZSO<R81-]SWIWG
-4.TD.fYQXW93837::+S8LCA7e2L2[2;[V>NH[722#U/I4V.bWfB)&V)#ZPV>3W0
gN&^a)J)cZ#CD6W0+]0Cb:NaG_D4]T44bP;,PGd;V-PM@5]1J2&7PJWFI(Rg:2&5
+53UQ)U&?+Kf8Q\b:J-C.UL4&gO1.[#bc?#-3@JNgYU#]Z(([#+BDOWBI-2ZP[gX
.G,c+Abad([,5<W0CeO0EC\T9W886NEE&Xc,A@#25);N(YW<E&Y.:5X?H2,[UE1D
Y(^N,._RX#HYa5L0<2Ne[(-d8=d_+.1::JO3##);(W?&EFLUO/?=LQ9U^P47XVbf
a<M0)UW-X9M.]ag@,SE:-PG6RLB;VJFS:@M-[33M6F\W1(g<aR2^Yg1Q\\fUKbb^
[,ZJ&IS:QVNS3MUgB\A;08^60/acXDdED8G=O(MO_UE:c7:V)16OU5B@I_dE8:)b
R:PNJf_&CI389aN-)KWQ/;0[/E4++(R1.W+DeTe=cEB_B0K/aKGU75NIbFeER_T/
_[LBQ=T)PB_dP)fVD5L<B=K,F]@7^d?@1F5#?cTYfGc6b=X9S=Zb;/=gGPGE7DAD
/>C]XJ?]H7(M:AX+04]M5?\VbR^c#ge8g#:ZCQ84)LeadUg6JcPLa0<T8#BG1=#R
S1(-W&PUd94Z&RKQf(bD;PX_#Mc976geR]<,QA2BUg6.JLE]7a=W=eObKUT2WH[P
XG#<+8:,b]G?+I4QK)@g#?I[(Y@b+]a=7?V98K#SFbSFVPDeBMdG+Q>F229[H[#M
L<90JFTIbSaW[N3[QXQIc:K-BZX=\_e+UJ(gQCEWZ8.7;=\T4d<0[.IX[Q]JPUg]
GRHcHX<A@-,:XK+W00]AQJTSTV-FX&+dD1LG\g=0]b/[(MPV1HFO1S-4R/80@VJ<
-B34]J(OMR?CO9?M2OO2R(WcVbSEY4-]_aM];F3NS+A<K(6/f9H#TPFS@]B9OF_Q
I<--HBSXYKA[\AZZ.64\3@[]R6S5fQe9RYMfQHT0]ZXF[-K2,Y;.;)Od>I11PR1:
^1VfdIEG.,-^GcEa&;6HU;TD1_&?fc)aP?@2&3@PI;bA;>g<:P71)GZ@Z<5N11a^
EP;V]CG(fS_eG#<Ga,Z6K,BW1S&,bJWCYUG9b0Pe(BHI9I)=<O&FYL44.O,;KS\G
:YZ;A_^R+J1#7KU4:1:&</@,0777aMOZJ^(3HTZ,\UAB^FKL@V.3<3cYIAd_<-RB
Kd([.Y.]+4@;P-=NS<<7D#DJC6HRg72#7R<3B\:6V7^eb.=)J:;@,ZNCIfP:59FD
C&80D519d:[g;bB.4S6IdST2HK]R54F(8,YNFT-,C=5BE6LC9O43;28HC0>U.>YU
SFb,@?5HIHV;c\)0H]>\]Q6,\KQ[Z.R7+5e(G?XX-Jg[M8b628@gYM>@@a7S]H(3
]aO,A>QZ0;CZH6HXKP]4T?F=.8DNJF/Xa@E8;Q0&Ia3@2\Cb.9ZYL).X)]LbZ3?S
6V?P459IPRYN;?P3eK;a+B7LE(5?/#,Te7eg.XCcNV8aY]<2JU0)U:#eT7[.6-fI
^L[VOAcP1)12C[<UA\c\bbU9=e7;[LMFU2&JFIGY4W54=YcD/b]?G1LNB5.PHZ]E
3Cg\YN0#L@A\MCg?\=E@eP;f8M;f3O[/#a2\NH?<N=9M-^<Ed/Qg_>-P;;CZXLH,
?I).6DeR&@9RIFfGDJO\R=7(,:UcBeeIQ#6bY9E@N-YQUg<>MEEcg8/?\:+fO/Ic
GE,UEd,+D2;M42^QXJYYRgU3:1)M=PcRgebM2=O=</TM,X#>&K-0QINb&_,53aL-
5DC:NPC1AX_,f?M)g:c1)F.\\T<[XP)2C273AMJa1V&+C#J)cW#^1JL_4U,bMI8^
cB#;#,^a\)O/Qb([YMS,J-BbG#Dg]7^WD6@U1E:3bUCJ4M-=,=&G9-UF6)XD&U9.
3ADD6A=U:46Fg4:NFB+Q_IB3&(9Dd&a).//P1+B2[XV]@+Ld87#WRM1K.]8ST)Dc
_HgUOCf\_Q8>C5-XU270)]\U2@&HK5\4IRC4IRa=OcN6F<N@0DH.RCO3Y3Ae1F_U
<OINU3D:(Ca_]74=<Y#PWWE4gGU9T#ZM2,0B+]PeN;KUSMa/NE4FRHC<UXbO@QX\
[XM;PHBDMb[]1CP.c_^Y#4;C1OVaL3P;CO-HdHEZ+556aFHB/SY?UWYG?>ba;_a[
>[dFf/P.ECDO:A&M.-Xc;-gFNT0UdY]S,S&;Nb.C=AB(gRA,KcI7IOFL>^^UT@_>
G5^>XNHK7:RRT]S#\U\Y;D2MK_bb0S4P2?ge2BOf5_-d6RQ-G5JISOJ(Z>b/=E_C
cMMF2O^CW.9[de1&M<4:;A,];Zd[1fUM2U57VO&5:KAF;WS9]GB1dYb[fdKDd@b,
H=R_\5L,b)c[3EJV[#;a?f(eU(>HG/HT&6B^?_7&+Gb2+/fLT@Z<eS@Ya<2O@S/g
=8-YGd6,OKY730/&BdXJQaVK]?cKVdZe=&,dH9<\^MLKYL<(,8Oe-YR=,aV,a7O-
;@T291.C3+R+WafS+,/OB)ObK-@#I9g9:[LgM+NbV?#B7bNeCV51OZP6)V7A0bC4
4M>.]NBd<b.;,TV.6Y0P,U^=6G&4Efg+cPDO67JF&1751edbD9RGG3e-Db+QUD(:
9H.S-ZaA3DX=cWc#e2X=3/f8=NO@?b/X]aIcEP:cF@L6?DIGQ<VVaQ],-ZB?,NTb
X[4HM];:DA^=7AcdWW^]5/2NAS@DZZV,&Ia4Da1dKbEI+^4R2+5KU^Z([c@Mb8g@
R.LX6aWE,V:+:];J)6;gTCZJcfbNKb2dBQVAH1&9fG81?d-T3M[]EdMO_a68Cfd_
.-N(aAS7].O@476Me_D-?UcIL)6=UaN-Q<&PR[eg_^P2Cf5DeP^.A<.G3YaL0B):
<WF.Z\_?O9IF1NM/FZN>6JAAWW,#a8Ng2D6f0<>C]OLg=GA+VBR@C;6NJMR3-:d=
cc(E31W=<NB08KCS]Dd:aRP8@Z&g/:VZd[&Q:U7H6<dWD9Gd\>=\S=U1K2>.>BMX
PM&9N,SgJ\(V8]d:MX4X2:PQ-fI>9(_E/W]XP6STSZT4-_DWU)cL4:FI,0)(NN+2
/XXVF2]3H3(\8W(94]b4:[g>7d=Q-N+[6gZ:3:>R<U]K77D,]a_HI>Y<38CYRH.d
0RV\G9I.)U>E=A[\H.^WO^I:MY]0EPY1@DFG?O<DPQ)g2^,\Geb5>R=)Vf)14#/c
AO-^83OfE2RafKA<fL]Ja2-V?8DVZU:Q9DZ9C9.eV:H@E=\4>E[YT8(<C\D2fbDI
?UfGCdfE93H@C(8^gfg7T]/[CJ2[fNJK-_dDYC1;LL?;/:Hb,/T5fNTXa8e,EgD@
MBT,E(fQ3,2#T=g)V9.X^MCF;MGD@B&Y]_/Zc:N;)G>1H+X-AZA/Z.?>=_=<9Gc/
YI2VKNY5eRTQWV>KK,#I4c()J^N+4aC_>ORZ,;2N6IdfK9G]48]H.8-/;c#A[H:W
[NYPK#J<+A4a,5)::\UNH5P2CWH3Nd-N4F8eNQ2g3MN9=FI@bJAXCF/U+:P&=UGB
^(/:=P:B^+DK0dU@]Y1XJ3c^+YN&E<P>F?5:WSM5;Z,e9dDG+/-VU57QDA_H[O0R
-^ACb:F9Hcd&gD/Z(@bO6@X.?:I;243&Y7TX)B<U96>RB<W/cU+,<@D0Qed,EZ<A
YI>?2GR3Bge,G<_e5&&#(C_?Q2,N-E#.X((#PK14XCH;KP:?N4?T-/e_MTb/=AM>
PB/.-NOF7[D8RMKd<Q_K[IZJ)PDgOMN9Bg93&87\AH]DbUXZBQ^M_?BMe33:,8<6
P<9SdL.-OXWFK0HMfePYR7U5d/UQB0UD>T7#Q8+K@^/(Nc4#.T;];JHeN&c:PXEN
&1&\[+O28;3V<ST5bF?+/Z+CZ73eeQb8AV@W3NXg^I7c1/#4],#_M\#ZYC00/^::
^\/P&#J&(dEU<;C?fGMOJAVeX#MbUWEbM,KdU/_dC9Q8T[IC3SH9/I+Ig;K+D\WG
_L]J&P-H+4RA+0+?2I4LWUgG7XUg=_ae:Q2O.;3NWL>AGWHZR0K41(c?CcSQLWN^
VRQ--3B4SLMBELGRa14Q<A(b=QNC8[-.-<d5BL+PQ3FX8Ka#>g/Fb5C]=1F&S.9I
<NGN_I>[0#<?[^J?&dDL^/]0Q^N#TTV2M.^Y5SK\,XDc0Z=>QaVX(7[TU;e8EXV2
-Vf56Fa4]5cR6aZQDe;W2S1FT[R^]#D,B/4g3PY:_KA085A1aA<ZUG/.NGCLTGN6
dHSA8)J:A<NP<E(F8QKE/C33MVc75QeX:/]=_>L=IY4RU&C(J^RLHPEM]7T1\MD\
FaNRIP([eBH6,+a?\^g?U,MfN-KS[A;TL[C[aD=_VX;,L3(,_XW\b+]_))JG(0PY
<V64#@4XPQ.K?WQdNQGb9UZ(EU4-]c]I-AI;FD<b8e>0Aa>U=VUV37JEK4:?=d@Q
7-FSfbC]C6W5M?2^c0SBAD#D4_2<_^9MR##?422(f(eQ55g[Z7eTBXT&Q5ZL9CGF
\:#[dZ-)ZE.+UMG9aK<def6<KGg8YBc=R&(Sg[#5Q<9FBXf)AO=XX=R>1NcFH:;a
VWRSP:G#_ZG)XVaGNfTaUY>4&ec_,:SVVX[PH8\F\;WH,ET_#U3D1N=TR-(Z6^>X
3KO-<&eW:aV]fD54I-_S;UT&a5Ie16,d)Q1R0D?CWgSSR4bON6KUa+e&CB7K2AEE
@8_T5eL,&,MI/O0HVMU^G1-I[<_.KCN0/4]JYO#KL:0B[3(Y(E_IgBX:eaM]:2KM
:T8>O9):J<FYH87AXaA1Q]H0<6S6PTF]R4Y8-9VO?3]GF/R?ec>2O3g8Ec?V+8[4
<XG7TPAZgXLbC6Qg3Facd(9/QFdQ6>SfL8.]J_+_H>+]-PPafABTRaeO.,2.5AJ.
\,S3[5D^V;;FF=g-#YI7bGQJaOfT\HbP^d-=\AVf;M6AQJPJ@+XeO<PB>T)UNg@G
aI<Y2]]M_R<GLMDPMRS6HO?Y391>ba@FR#WTUGKV_N;EPI).9a\5..M;ZI/PDYg-
fLS^)ZV_3H0FBPD]HfIBY.,\RR]gCN=2a&g+U;5\NU>]GWIg4#d0Z.#GN#@F]-./
FKUaGJ8:IT]0;/bec\MWG1BDb7#cNA?B+c-UbC^#f.<2T=>Ob\N+I>\,.QcX929f
UVO\VJNTU;+.3[KT>F\=TaX(Xb+]2WHZ8<ZOQ.fVM1TEIKX_AH9V3Za\AfRP(VAe
@.ZcKR#]TULK&H75IgHU_H2AA^PN//T0)Y>2d-H2N[FKD@-LJdKd\&CXX(c3<R0W
WRC3[C#aCPREJ(@F/fcN)3^-bQgOb_:3fA2[+<eWNeVF4)eK3)C(S??FQ-9[92SC
1@>BWAUYSH.@@G:AQd788A+.DCJIY7[+4./&A<7_GEK@DJJM>Z6H7[IR]/291=a)
:/4([>dJ(J=DO:-P1_VT<N#CJ.K>A.)GO_7Lec)Ff#0;-?2FSg=8,fV>[&[a/cE[
IW;:EUVV.K[IbY]_aL0aH.[U[d&bOQ375]VOGC#YSaS/Q[IX/77g,=-Zd1E;S\64
C>fU,g@E2/H@;5,gBYCV)(.L,,02b[11P_]<9JE>58NJC[d5SSQM,dAe.2a&TcXf
X;ebE+MIS&2]-SAg(K)&35A.R=J98.:cQ7T92e(]\TOeEgQQFVP]+e-@\WCE^Y>8
@VYCYA6_BJWU<=3[>Q;bXN^[))FZ/ANTWg:+O09#d#/)6c.F8CVCEYAc1IJ9H/]c
1I)?F_=I_E256KEC5D\</:2N:4ggARC];I]=PR&L);TX3H[<\B8]]DWaF.fB4(Kd
+;H>/&KWQa_XH+W4/AD7.EIf,Y(819b^cGJ?Oc)2FRR92+[C#5?KH:^DH7E>??A2
cc22&&G&F:]#<^2#d0T(g9WSg.U&-L(^@;4R</^.fb\UF];DP\<=<8V9-;D<32dF
?#3:;+(+gDE)5;ERAZBc^[XANN:7O]UT\GLF_Y#,dAYK[L(D9ID,BbHB<>-Ra7B#
5X>HF,S,5;T]GTHZQPd)MJTV&NcNQI[)MZC]^c/9c@EO>848g8f&Yg+3+](^=.:e
5dQ[9P^:?5+:.:S[V9EXV(DSb-;cZZV@OVM_7.g\+D(C(8aRP[VCON.(B3./<d4>
KA[6+E+E#c@^;X)42/GeD</S=(OCa]=3;YUJJAV(02[3:OF8&[8F,N0eS\:CK@TH
-^&DcHP-L^&[X&\ZA0JX#NUaa,baY0_6A3/^8AT@B=&dYK;[)b8\W)I=M#e_)>\K
ea@M#98?MfN^?RafRf&+)LFdL^a]WD7-#DYE5JB&B1bR1G<(T+-)Z+4[?\c?W8(b
OQRcMN];ERCQg>5=H5<9;M20;S/J#5VG]cC6G;bbeT9@U^B8.+eH5B6:]>9:FZN)
c1@M>5W:3=fRd]Ef]Te28K)eY&ILUR-W_;eHKY_>6SLD]D^E],Ye:5+>>2#DJ#AI
_DPJ85LX-MIb2E&;>,@g9<4b+>Ff7@>(Y[7@8V.91=I7Z#NK&eA=f&@bME,0-VB0
_LHD33TPZ[SU)B;RXQ1cJ2Ad-S+;N8I-P2b[>QF(]I50H2]9EcVAL1<a+\M3C2,L
(.K6b]bSNM]KF()f=71Ic.4=JfH?WI(TfC:&&O>6(;(K6^QOF4->9df,Cac1;ZIW
3.=0^8(EY7BELKK-5N+O@JEPT//fKOd#?.MU)bR>7RHg0S4dFQ-S,DQAY1/DE.B1
9^d]FI.8RJPc#QV)R>,>:gH4WTQV-C?3A280.RHZg6A07,2EgNZ1O05W4C,CSKW?
>+.(FX]2+&S1.Db#6_R2WY>1\aJ0+gZVbYaLC=PRGY?D3G=CL@4I&O2,fWX6ON.e
0f._P,ZZ?XQ\EV<SedS4^R4>^L9JX?:((07f>UA)gWb^UNOMQH?<\#>_F_WK7FX6
=TPXS=X2Rc7.:Z0HXf@EDa_JC+DN1b8S(<Q)9LD(+[G>84Z3_.FZC9ab=8fN4W:.
WVJbUe0]TcfLF(g5V#IaXb@<g\DAG(E6(2XK35a+O-1CBF/DN^McG0^VgaC?KXD4
e0O[[U]b@A:YMe2HZ^>S=ZC9/?<_XNeWNAL#:8W,]Q\01.V?g5e?+J7+1+DQ6]b4
N?Q^8CeN)fe\):0]6_GBJBB7L;LBCLY=O[B408B4&E=eSR:aDRLOG2A\QS<=I^Cf
,^;.cD42(.T8+7Q)Y8AcJ1MV#?]4aCTUB4?\9M,F;&<-Pd[PKT0cO3X=(T=d1@=8
L;Kf>7:[OT]?K&[0;CG2#-0>V6)^_d?YY8;?EER1HWQ,IGdS4AReMA8N6d.A;HcC
b_H/3YG3,ZAHM#5a[cD18RdCPX)[R_E<b+A7:RQHfL_4aeKX;XMfKNd+IB5XL\\d
4?g\AfT:c_AMZL_\;Gfd\#F3)e\HIFAXDO?.1N;9KE,\WQ]:U&3\?P(NK^74c49I
V]#\4]Cd9PIO2DcV^6TcHac;Ng,42afG5_3aV+XZY,\(d)OKLePC9-C:VF:[DG_g
KBMf,XZ[geL#0;^=5B1a:cX5N,_5&7Tc.Y?\<g6CFf&9B33OHc-WOTS2.[PeW=RS
O(?2cEWM-B5HA_/dBW(=A^Q]]T\PA;LJf38IHXIJA<OfZ(OF3<Y1P]03@CXg2)d=
D.5[8&d02\W(RZ50VK2X7.H#ZYFUGK<[^&618<5,<U^bHO,]Z;@XI=M35B5\WZ5E
+#<gPYd;:e):Ge>/+gMGOG@=KEX4E0N[J^UM9K,)DS6UBe:QZF.DT[=d3f;9SfLF
3,f9OADS[RO9IVS0])2#[BTS:0C+G/OA_^]TN[V\b.[RPS)=6X^KZb3XC8XL3QRa
F+N(Z7.24_,>7V7#0:[6>_#5/<;()?Y\<.YKN[bY@+&[E^)R6>5f<,g6a4VPW2IO
-OOR;eOT1+B1_SOESZScRY52.>e>@+PL=;//@#VPS&ebY0-NAP.T)F2N73GRXAW/
<R>f2@H4M5Q@U=9a-4.>]5=WOF&&g8e2ETSb(JSDR-NdTFO;0VdJ:b;A</S2TA;.
>R2B(;f?Oeb<0[IcWfe6GY_++<ZH-[E)MU4Sg&&dZGILI.-KeXdaL_Gd[RBHZUa(
Q1]EU-2QO9TATO@VZ+)R1<>V=e=g07KF/>fT/25N[a+Hg+N\bLMA34\f/Y_#@1/c
0?:Z323,<Egb^P#2YF(LRI-Ld\d2f]Z>E,&,G_c=/^4LaD0?<+9VCLIVZDV&HF2X
K?R8D?77dFPcYEa.R5]ff_NU8=YTGLP3#,Z<_HP.?AFSE)1;2dNY5+e;9>A+;9HG
P0N&S?(A.bGYW#^HC[&XW_PWL6bg+e,&ZPRb2-13VA>/b&5B:f<LP?BCgd(A@/YK
WX#L#2_f0D.VK@&>,fe/g@<.B_B6F5Hg:3LZ[+b2YW\J6De+Q2.0WPD7cG<16J/P
O1(aacFCAP)#H\;?^WTf#2g5>+HD/MDS>A2GR#<DH^Re[/H^I4;e&#@5B\8E8SLY
GcHdXU8.cA6ZDIdTfTWE+ZI94Z]:Yg[GW_GcNQ+S;Vb#a/BGaV(dYV7DRHdb\:P-
HMNKd6)OeKI)2gF]GE2I1_1c.>BVg5AS<NF4>=E6S:_S89ZW&,K/I:C]?f-&cOCC
_G-;L@/EY(Z=+PHT#B9HEZ^dST>E_0PGLg@E/XEM70Z#E5.K#PE+<^gLPb,Y[Na?
UZ9Q&CD4,]dXKeCfSJZ)MQ45[CSTAUPIMVbW3a;K:3YK>\UF?32T_(0-W4aK-e-K
ULgY\-;/4?#9IOJ([FZ@DD<^Y_)5PfL0QC_-1D2DPG/JHe:2G&Rd<EN#MX3:C9-;
NP6;>N&WZM_(T\JCV21&ga.AJP_;dC4H[SP2?B-4#V.U#C],]O/@(V<2AGVd36I9
P)DCfd@P#G^1gfdIL>c[f#?352.ReUB93;0QcfTe,L)Y9-a<7&7\PP]K_WQ[9LST
CJ;GA[UPaRbNQ;aG077C/E7MZJFL-_e&?D._SbdUK>B&(]K5Sc>d2eZ=RZ35GS_I
31e,FDUN_DI^#]_E6V>[;>XY<YT.XKaQ[N_47T_:G/@=Y[OP2-USLWGBDe54c<)S
04E?6NF@TAb5H8NJB[f,QIbPFAe1?.,O;4Ib=24/JS[.fH_-ISM=YH@41J:faZ1,
gF_&+2?Z@D\BD&dP#T?YJd,3Yb1@Y4L-=c[F#2(dK:??LG35#RKVJ43>A5;[D?PJ
I9/(C?/2/_\0,(;IT<DP+;3\a^a9V<=Z34L5\1E32_(ZFUgU#S3CagY&GP4T-Q87
Gb?Q@<&L-.>AH^&:MaGE>];C?f\-.-H+9+@<YTIZ^4?ZNVF;8L+-aT8Z_c_E&^;=
,H^J4&^)_5Oc^X3YdX(G.RVF#b)c+OP4Zb;f1K]DPYP8:cW5IMR_ad^Z=)<L<98M
<9XJ6)Zb1R?<K.I[SN:VJ_J3U)2MFT8T>?\QSb=5Ed@?>PL@d=0B3#g#O=DDPS_<
CIE+=0)^Z[cQ+G@O\_ffMPCZ1;cJDc.gZFV54O^\5-\]L6L7>/R8>Y[g2Q#Gf1Ve
Z-+[D91HFY;5c5G-L_D\D&O,LGT?+R8b6(H_9<P1KI6QB/UBeQfPAA_ZNg.4/f=#
>JCES(Kd)5J@VW0L@,#A0I@ESYJH](L1Laf69E9K.-4)+M4ZF?CVC40+59>JX8bg
&dGL>H;@aJ?be\\4g8NQMea19K+RE71_7@_[A9,F7L3SS[\/=&N[@&d^e.JVIJ_K
gA1DdT.2P.<.>#:C0-0,#^)W@NZ=XZeb4^;EKS6TI63I&,6&UQ8:/#cV\Y3(B^<9
Y?:.;@FEZfOEPNaJE#P9\YLYCS=dP.712Md/g5A5gTGXM:+ZLP?GOQ+JfQ8TXbA(
+))+7ZV.@Q5HXL^U;NKT,,I.M7WSPM/SE>6I34&L_M?^DV31:S6dVfB]D->@NAN:
6<BPY2V&X+.=;<9>._A[Z/g:cfL<+W-XZ?1W:6gZe4be<D;=fga#?G+WZEY2HLb^
)_09EY?ORe7O7GS:8(^2AM+6b,^MO^\K.ZKeNURP\1JIY,N8U>aE2S[PD:XaM/cN
)f]UD(F)&[A?<,.FCP]1FP8=9YD^#0F[PBC,3D8Wf^^X-b2-HGGfLB47W5e5]_B-
0Fb=fW3PC=<U82A/71?5J#9d&LRaK9N;GO6;0HG+\@-FY;G^d.=aF^+R4\15]<S/
<1eD]?=gS-X@HE7(F/:8-fZI_B8WaGOWI#\6RQg3)XH?T48:.UeW(YF(31L-A3Z2
gOFXH92.<R[@V<ZE5\bKW1&HC9IH>CV294[090YM:R4WL>K4JIXbO>/+(/FJY7<V
UcL-0CFBP;L7TWaFZ59AIE9fQ<^4:@1,KH&Q?A0;TN[J.VSb;)HE+0,@abV4^ZNO
;.2T/-7C;4]S[K#;daJLR(-W(F^Cf<V.>Z4Nf8ecb+=&?JWFMB:\)G7P&._FQ<?#
)2US_\W2M0Y2/5R7=.F22VRBE;8+8MB6/Y[=Q2)0J?Q-(0<;O=8C5B#2f:Wg,ZFe
eQJ_eC@29D^JP4XE0a:R40X@A?QELAbPM@cP],9ETNPQYb26]@M4#=a;62QI:\GY
?YLRfRWIYYN:;06Z2[F,@+8>91A[,6M8RIC2691>?U8GP.,LU,0cYZQYZb][^bQ<
ceJcQG5PfZ.&6=c90BATA)b,:&9&aM>fF7-Nc>0/XQ]0;9DV@]3f#Cf2c#bAR71G
SV.5C0UHZAMKe3-&(27[UOQf:I8ObcaW@de;I2[2/af\;(a11GKJ7Q:^I\;G3QZ/
&^-bB13J0&/b<REg^2+>AF3\U=3F1KE+ZbF>DIc+MD.M6:WTQ[CH-FT/.@c_Q@0Q
]O[<9HL#V.OM<I+9a.He/7+EN>2S]E?EJOHLd5J9VVNg+VHV3G<UAf-I44)#6@_U
S=O;5)D]SOC6YG=g3F:KO=P)CWCD@T<MW4KKfD.2GZ;W-87]:W=[.[63ZV6OeJ4A
,G=bFDDC?^TOGL=33+>O8_Rg#-PJAg/K39FF6>SI((U+0?(T^PgGbe3g1B(EZKJU
R_1ND5([PW=@VE4P;B&97,6\cg8JOH2H-?&g)Yeb3<L>BSA\ZaYY6S@:=7STOD1,
NECg)]@[PK29VONOJF&B:.[6;a_2X(;2I(6-df[;Jg,;T#HM]f#2aK346KAGRdX_
V:X+e(E<9&N-L5Mg@D?7Q&E8HFWOG?JQD48cHTXE1QQWH3Z(2K[QHAEg4^aeI?\S
0IPY<<==C3N2)#<bO:\9BSJ();.@9UV)YUCTJ\L0&+X:ETHB2[(HBOU&YO\ZeFAZ
U,)b:NF-ZIFRb=7067GP6FL&ADR04XX<DN]D7578TKWP>KFKA\?;]E@4@9MfgfdB
e=,]NI^=d\)UcU(:]=7CQe>g/N=f(Z&@A=9=]@?F34g::Z._7C7SPKC^\QNR.0XB
0L:AeDfH2bLW&gHM&)?PTHM#+94-0#.<-9/D;^X(4TXL5[(e,(@;]G)R=SJSUUdE
-Q-G+UC3.f)I0&-L<QU+]Kb#e/;>Q=<6UP+\^6<g&B^)RHFa2Y@QE/UE/VH46)MS
D2[G-X;]>&DSHSIN2#+]JPb=)@f].4CBA>[-+E\@Z?L(VG5NALC&NUWP_g44fOY6
3X8RF@+R;:I]6ef?/&9YF_6MKL+\]#;N+.7aI>GCITaJ3ED7[?S+:\Vg1.cH@HG=
H4JWVJRK@#],-BOb@-9+@)SCPL2fb2^Q:-9C+C0PXGO=IL[eM82B>==FVUHOe1PP
O^JDH<:0Nd0ZD\YJ(8GLd)FfVSdBNc./TDgP64gg_/70faRO=Y&7e?VYL]5W0/[]
=Y9dM^F5WF]Vf1KZP[TC[+0]eLUXV-UAZT@U-d./T3+L^?Z#ObL=5A]4:CdAI=]6
VBV#g1[[g4)Mb&6M?a[_-8)H74]I@BeW7GZ-[E2:aL/5]K)Vb],:RK)S=:@+TGDX
SD??&,be^fG.cWRObW9=THE<@c\UBS8Z7b:&cBL,H(fX&;/D?N[:2ST4:b[2E[A)
@S/c0;@R=0&2U<b:><U41c8XTdZFH-.4H?;f:P+8/U4]QWMPSU.FJ^ffAUYLL7X]
g7FcZJfP5XCS>7>Z..)4#5-3^>=3a?+\GW,Q9BgZK^^&Qa[f-B8=OXbdAVZ3@8:(
PgOd9Kc-FN67R):\LKL4b]OaXCD+)6(7J]b(7:.3EYTI(bL)4/X@<@=.M-NF62E5
<c.FP.3cM@45Fc-D.&O]HJR[c-aY6&4AdGUg#[-#U,JSE7#<W+U2/FQP50,?(XIQ
ZB3ag_(6Ba]FB\&M4\F_)ZO<AQ)V0PFJ]4.ODPGR;09(_B6Q,9X;G-?RfS?GFZH4
8UaJLc3MCAS#a8HZZWXQEG/SHHU.R407PY85F[(SVXN)Oe^3\CDB&JWd)K<,PV18
HOS.UV+YeJ.7].edPB@2aHK,.BP3)+8(AQ;<8>feZ?Re_7_S#9C[;GPS<Y-bV-XR
JP_-5GW;J73gH7=FdII#=-e=2N/Jb?P?B8U\ZXFGPba2WH>]3WXb)(\ZG<C2#=fY
/9EHNO^7+/b4P6:U_WeP1D#F\XH7FW721g:\XV8eG,9C:JA;A2O_,Q]9D\<6GA@8
9e6B0fDYK(5BL60O9eC#M4J^0Nd1e>U^KUD?cG>=DHCPH]ORRgGO]QSAG<.f/G]F
=\A[3cV0)HfNZ)PCA?K[/3T6Zb)V05b=A#dWV?[&UGX5-O&5LddeV^T_,2@<bI<e
,U)\2+Y=b^[(U2>R77720g.#:#7(&NOHEGg.gS[?0IF6._?+=bAa8XA9T<;LJ[5_
O1;#D@(KHOCD4,?#A8_&)M;8LfM:B^BD=[=1>&C:TcKeP:62FafD;[:&=EdO_df6
f=3PceU#\dE5,DG+RR6&.RQXSI/e:C#DAYO(Ne(HP/.CY(<=a(>eY&\E@B<a)WJ.
/AX\N;9CYKA&J.;(g^,/4cf/VKR)EH5PB)0A=W<3HHW9YcY8990H46SgIdf(JS==
12C=)TF@1QBTXcV9><[(S#8@7?.d+Hd@.[>Ag^Q,Y@Cf2AXC7aC,HI;/cPC]??gI
fDcDL9JAR#X3D[9(=X[HXW<<;eSQAV5W,G)Q\?V\J;A#E2a3SY1.;=<7)A#8C/,;
U8bgd-/g4U0^741a31+_d_]18KE1d9IEUU(F54HJ:V38/^VeN/_@/)>g.U7,>RL<
D#b\Mc5K(F;(Gb8D7/OgH3IQ01Y1RQ>TEK1:WADD\Y,CC^\e8#cTXCQVZ&+RVe5c
g,@b#<SS]KGUJa4KFW56A,X4c>P5=.9:T#&AG_RU4>.C4FL,X@+H>09K//dOGK,=
D#A-B73B@:K_/D.Qf\8KeKB(3fb(Z+RIbDRa\Rc+^.,Za4ec^IFO:<+ZHfeSf\?(
E;>S[DD6UId;<ZTQ-C+2FECSVFD/S:I@9:0X=?dPFbbcFGWUg[a5D)Xb<e?<NJ3H
,F25];]XORF//dRHZTceT7HJeR1&M?A)8?U(+T\=4)[9VI1AB3@[<K.V-:Z)^\aJ
9I.&C>R0G#A<U5H2I@fb[]/MS(0M0,H;XY\/2X;gWe>Y7a7Ug50O4C[]S:dY;O)K
C:+^e;P#Q/).3X@P6-I2J1I5)_5PO@A:&)-GJE5#_5JY\P0(+L1/3dMB9LE1HGDU
O2Qa/Fc1\)9T,A<Md;5]gg+Fda1MK@\?&+<TERIN<(Bc4#GaC[d)8J;^(_IcEbDH
UEgaG6\&URH?JRDa&OHB^(7=Mg[:L;;+-e[IMJ_S472S28#K&NVMMIO.PGQA;]\D
?(94?M(DF&Aa9A>DeXg06KZcEVK+H9f>H]dDBIZ6]JeN3SaD6d,NVZYZGSN-<WXd
?c5&d2Pa(9,CWM;(MS)WcX]55[WXQ>79e7eAe#Pb__<c,M+U781H8SDbR2IEE7^2
1LND>GUe^W_.b+#+cT[[]f-T3ZGa[#:X4F>EPf<119(WTKgO+I]T1.7::F)RM^+3
0B;1>WPLF<</Z^eZ9EZ.?N/>RSc.d@NN\@-)3]EZ.L+POS_U++N5.LLaa3cEDJVI
E3f)c^F3F[S^GT@f1-^dNQ6[,DgZ_-@1a:_TP<P/0a&J/b1XTK@69/7gEAO+a(DI
(a-c.f<9I+-EPDf[0),FLC&6&MWbcKB\g;?E[M]gO;PZUZUA<.a,bJNVBBUO:Oa:
Kaf92S4UeHY[&E\>:ESQ)?P)GXdT8>_(CJDB^IMd>EFJ<\.4FT]7:E1=646MZRPA
AZYXSWd->^W^Rc#AOGbZ&:Rd_K?c=?YJ3]P+Rd.e<EaU]b:Q9F3,aKaXZ_4+[HZU
\(V,?@ePe:--M@;0(95e8:E3^:M-,(2Z[=X9[SMQJ\B=0I[4E.CG5<c@92D\^?cG
FM:+RX6H/LbQ,=D[_c4:J/V3?HeOEIVEQ.):?>IU;[YXE,?1]M0.T[DYP2GF16#>
PdG3B.E<dI=CPQH6O7QWW>e85?VS^P_:;O7aO-JKF+C>B&XP3/6f(Z)bG[.VM40d
A&=88E<(Rgd2DaL[64?TBM4G+dG]./6DR[4>g2.IOd3L/.0cXW#-JBN5JO/=deV^
JC=#f/MD^94B:D+Rb[,GGJ;K@NJ(/f(bM57C\;I&U-cR?#XdBHMG\>.BP#(A83#V
:;Ed:C2^4EDGU&Z@NUCG27->38RS0A92<W@OfGHAPZHZTOG>6L^PbMa(<R]fb26Z
C^&GFLVY5@UR)?9CCLd-f7Nb8#B&L@I:4cEW5:><KAMdTW>8>&4KWBd\NW&dL)+O
7-U2f67.K5-G,+-5L9/+I<2)H4\1J=J[_g^)K2BK-1S<9_0O=D_@Td.O-DB^@f.0
.SGT)Y#V7R>ZI+9f_9@bGeA0I^]I8ZRUfXf2ABOIP(>SW0R>FH1/;ScPS-f]_<?A
@;8TfYA95W_H9[S^8cK&]=6ebX\/OILB-+Y#f0R<#c0<VcZ?@ED3-=M)_5<5;NI2
>-D_<TNXQO:(/a3]5-_IKH8M^I?YR4gaKSVA5d7b]WK4-B2)S7Z<9R6)C#35^;/0
95\NKZVW+?-8:0SY,\QC\6?J5T7bC8K2]a5+C#O]..3<P>BA?O^#U[D8aQ,#@61&
7Fc&7GB\f8_602G9ZEZWU,PPK&YaIPa;Hd74RcL28SURe(4.PR65T,DK0UW)+ab-
.Ne4@?G@/>U7QIA93?-g_-LTaW-XWbZ6]NYTR7IEA65Ea@PP1N]bC,A8WC=TDe;H
<)&GDDEXFBPUCMcM5S/Te.[(_\9LZV.=Q=(V54f[?a:<V+cfZ)@WTfQ^bP([egL9
cY8:H/K;;Z-0f_U?<89&<Wd7C^J^3AEL>0d?V]I1B7>Y^KQHA55Kd]G7WP:Y3Kg;
U>4&3X2<g=C[:^C&eOA.Y=[((YPc)I(SGJe:g9_6aA->1(KePTK;7dAP?&gd@H6U
.=1#:5c]ga[3TF<P][NKTC8ZYDcTZR-NBZVN5b=CF+&-@__1eU>._/.OT)@bdR7L
Z;-I+d;5N08XZ3F<=\KY>,QOZ?a=;7,E@b]J\HdfVW60[Nf#3O>OCCaLZHHC&56+
WEE4c9R:C^CA#QI6e/I.@R]V#4a4dc^c6^+/2LQ=A7c(SNBL7I\cAX,D7b=e#Q9V
-R6@U_)(-CJGdW\AGU=^2Ke&B009]B7GGQ^CX5V+;SBaQaPR&cAI>b.RC63Q2?\=
WA-AVcT[66g[C2b[GG<R;DSRg^6&fD:GI58?MRZ=?3>1d[>f>GN+205N@V-WJJIW
?F>Y\C[I<a,F;,fc=_&KX4P?/N[F=(cFWJ_Q)E/+I]:]8/.WMg\<VH=XB&(:J^aK
.?W]CQ)TEDC^e5==fKKN:D@&9>JCU,2,Q.EUY[]99^AIg\R3/O/=SH/19fH&47DO
^FTWgB_+WL3FJ;IJa40IB[T&T_fY=38SACW#fP.MDDUL:Q/g?6LV?ef>FAH6ED#?
F_RCY,;DEDIE+6#aY-K+Ab^#4fX:4T+1:cQP0[<e.CUI.[bN7<>W-.64F<dB0HdL
F2N7B]LPC1#+_]F]Xd@7PeK:H?U5A5ID:_.DW<&FR[B57:FJ+4g@<]77BHYQ\.M\
adC1.9]T#1X9<C\eKLDDMD_IMaP&a7+Z<M\VPEY(8Z+ES3bO)M\IU9UQ7ZJ2gOB]
<?](d\24fCRF^GaU.]@?aB)4P_ERTI[ZM=1;,Eg;L161TU/L/NG]/@?ZXKbVQA&d
@NV@W-S@_CC#]M+.E21:e?>MTGJVcR6S9(O^[M/#S9[WSdQf.@c.1aR(6.d4KfO(
FfX;e,/5H3?OSP;e1F/U_6F\OENL_=3TP\MT:B\8I;32N;/4-Lb>Ob^[\+G^K-)8
Jd6KCWTSJ1-YXP[ND\;)@e[-9PU+-J#600SM[91eb>7.=3E7?g&;F+Mga_>9-D+S
\PCG,366]6a1@X-g>-dSKgN]^\0DDaRQ-a_;TY<8Ff9NA:cFUf1H_O<WN.#84D&V
6a^NZOX6Z4QUY-0-:H\@gC<7G?13HK366b>DFL;+Q2PELa9dZK1F_[Zb]dU43OdD
7X5B3H<N5=QSIGN7]Md(22b[TGX^3VIRV(a+ZCMWeb/Se7e.DOYN:)d9?6cYANSA
]D:[)V1T,;W513MDUXE(95;>L](e&T^G;7IbdfZ,WfOQQEG.WYWRZ=DL6TFE=RVR
=GFM[<?#_bNDIP6<AS-D^1O?;X;Ibg8-LTQb)5HDKHT>F?\>8E.B_Ne?1+dM,&YB
A,[W;L1/VW;P9/:62Vc^;21\M^g-PQNR.L.8)KU32/&M70fbT:9SWW33CQM,PU?.
[FGZY=?H3UI+JRMED2fNG.E/AfJca@bPfaEcaZ-.GQ=e99ABR/eZ\DG_AMg::0>H
/R\cXA[SK3JBf===ee5CVNJ)?Y2e:[R<)A(^eQ6I4M#IEPWRaO-U5]4F&1dP:84^
(<)8V0=1PbaL(.C5?&g&O#LLZH2]L;2EQ^-JX9VO@ff:CI1<5XJO-WGEL2>[J755
F2.FMB+:AeaR:e&JaII^(LI60]EV.ZAU;:a\=+feR(1)792ERW;H:M>Qc>38K19.
)OLUgJgZ?6QfC2F8c?1,WW.XgZ?TC.G@85eA?NX_Ce#.N,<CaGRgS\\aLJc:H+PO
&\\Nc4?WR,L5d.5@Jd(QFBD/.^_Q#EY);L5F0H5QY-6VLde7EO.g-5[X5DI-5T@6
NLIVS/ee7QaB+B-2FLMIF3&<dR\;.026fFJ)]GX+RV-XE4c9dHWBM;_AK_MY2XDG
XW+,4J0J<)0+X@2(2-&<W6-<Pe0DAgT>G7@8BJ,bO87T@_=1gR]I2:VMeTHOUTc0
d,cAJW@,PXL&K;J(dbH7^\d?1Q2(Qd<9b_f1b8I/+[Q;_QD#7cB5bE<G6>6AaeV^
U/V)4=V.C8eI5^#525;^]P;aL5U;JbcB]3Xb&F/^f)HFVW1(-3MR,b7f(+6F[bYQ
[OYB=)&RdS7Sc9(7[Cb78Q@:+[6K-LJR]LdeTC<7>fWJ1d7?6TYAeXN(/,],H(K^
\+CFa(>^UWe9>&J0bLO[+UQ6M]g+;Q3:aW=JO[^W0[\TZKaBTT]#3[10X8b2SK:P
N\&MJ+F+UALF=6#&-c2<\-Q+ga;\A=QN>(D_TEY<-.=K=B.>O-VP3RU9]<0LIW-.
MHf/>A+8+IT35e^9R@6T+F>@S38B9+96?e2BT[Sb7+CS5[.KUf\W:(Kf(e.MIUcX
]&-+21caO7<&]O5N<2E//48&G8[6&)A(ZT0]FDe/(BQ5J2Wb0&WAF]#5#FEa4AK+
?H@-;N9I&PSCXGI9\0EcPZ\O/AZd86/Y19Y33TIP:V>&;:VR\RORDa<9TYLAQ?<V
SHgdPSJG@PSZ8a;b-e/-OP32#NG2f6+T?f/1/I..H7-;Oba2KE>H4XWUE0IF:d1_
U9Y]UX>Q8ZRV:d];WU0,A[/7b;ZX@2YYDS[M-3f>3MOCa8U\La&LJLI,F3V<I>6)
3J78XXTV5/=G39[#&-S=V9\fC.\:TCXA;bL=RBR23.PXcVV#9?_);=d7>ZI_Rc=[
>WMS@O+1@9eZW-9@;_-80E&.GE)f:E-KUZHf3Q>X3Rf-+>,b-aQEc5?I@GfH[R5:
Y&C7JADgRf+I8f:0T_9I&GZdYffFX#4Jc:Z0).+.8gfc?dTG_CAHaF6MbE^^dBb@
OZLLCNFSTE6+,g[1[0+-5GAfSdJ_P_7)5&-^8XHHWgX8Xa0UaVJ/J5/>=#d2QNe3
cAW3;:M8[d#CS9G0BFXeH=;NYN@GC0&g7f@?>;e+O4/#<LdEOK7=dPPV@+RO(BCQ
B\YK;7U[b;2_.R=FP<fG>b>@5NC-5../e9=BbP\4,B,PUb1:<_?>=5RIG?/9Q\OH
]XF&Lb3VW;^Y>>c#9Ed]IM9Tf)UDU215)bRNLRc,,K/Z88LKeU91=18]PWXQ(]TX
;N@<YBDbE:8\gB:OIe\DLQa7/cOVZOYQDSbC;)6F/PI1:Y7XW/5OPZBab29_XQ&0
gTf2>.A]X<-WdJP6PO/K&TcNLWP5aHIGZ#]EUL:2)CDDOO4[NgIJ,12WT1fIV+6F
_dW(?Z>,_Y\6;I590UYT)1K[C]^V<A6&8+#I9\6MeOL,c3Q<\J]:>f:LHDITb32)
/+@36eJFW51:ML_,)>E,36R)]S3c.-_@S(K+.IU/[dS&(IXVLIE4TEa.g,:,;G9+
()VZ;dB-=6Yc27[Ld\G]O6K\#,IC,-D:?-.BbHLOKBNC9+EcI\VXT/=AZBgJA9BE
C&b]HeMe]<>ZKFS4b/[^a9+CK+4f=J(@egYe9a>F@HV+#dGOL-5ZG,c8RdMZRe\1
/aeG\06)C(CW9DF7g\LF\L???[CY]7Gc-9a]9U8<70TWFLbWJ^H;,H9#aBC1HGY8
g+7A+#a\XPX>:-EKY:4.I,IQL;edV32J?S3VHUeGbc^(=eW;<U<;d+QD2S5>bGA2
@#f#+O:39<,H-PeM_2=4LSJ#DO:MZ;bWXPOVA:+EVf5.J01?)/13^:4e8&7V,P0Q
;a-NE,7e6Z)OYIIIIR>4&_+GE3:[2A_MFK]2Y(+2]\GOOZ8bW;.^/fULUEI/dPaS
F8W3[_.a.=3Re_03&?5RMS(TKUabMJ:F;c.RD3X,KI.beERRN4NKbaT5bD6=^f<(
NQd1K\:b1(T?[e1\CUKXg&G^DD<T16[WUI>56_VD_F15.J44S:g9&gCWDFF#81J8
110g:?S)3[QPH]Z_13)KgL5,Z6bOa@PN;.bdPG[NDfCEF4J,WF]4Q,;@c97a:^<_
<XOL:NS6GbLMd(NbU#ab_[7AGgN<+Q&V7I/gM[cQR]PYbAK^+\E@UQCM3?;/6Y^^
78#^4:g]+LX1\)4U[4DB_c3\G1J8BSS/D-+^PBfM5^TIf5dKP/JVUDMgC.IU;aRW
beTXd1a(/[<)+7^PMd@W2H,V(1Q+VADc@=&&:Yb1(_T@8IA+L(Ze]W>PIdA=^H&J
WgW(VFScA9ZTT_+G1HY;\N04MgAUU6\ZFaR;PB4YVLe+QA+(g9CJS#)VD(O3d5B.
RY1@5E6,#e?f6F<\^95)G(YLQ-_)HB3=-3-5[IQcC3@U,5P@ZQ:8++@/?),PC.0A
=]gaI>=1:g:X1&.6#=7-ZE8]1bWg)=&1[SB)M-CA6eg2]&LK2Y@0HaA[4)cW<5RF
L_&Cf@#]^.#K??cHCKADAN/#\?O\cID;27S?EODSf/[_a,9Tae#I;SdM#AWE,GZR
_D(:B4/-?+WfL6=#^d>g88g,9-D<PKNVe+QE_@cV2>.Ob<)?egd6/<-0bG;[b8MH
5J<7^DY7H]4?bT#I.L?3E1eFYG-0[<H@7(+;[U#KJ5D:f58W2D1K-+Q<)34#K<>g
/E[V1IbdWI/ED32:N9V=6Y;G??^SR1O_Qf=P=Z39eC)]^250\Qa=2OUYU9\AT2(^
,6KG+<DeNT],4173]^Y21T7,QHK#UG[&4eB9)1)ISb3YZ,+WY/bg4d+U5+]3?7gc
?C:dHH3@MbIa156JP_LT<O&_J>WMMK;9PUL;[L.U5DM6D5-OQ.^ZF=^NOFY1Q]JZ
=5F>P<4L27JSM7)_4#M\AKBU2I2(0\Qa-;\J<f8>5#gf5D@-6<\g7)<O>EX/aG#H
7@:eN53E9.S[/Lg?--70+Y#55c@TUN[Bd/2WH=I26X:6gEYeEFgIS7(<_^DY?HPW
KbG5M[QfDIdc]CQ=f1_2G<<8^XC8gTe>Q9,SK8]7gDPa,729R8QN6.3Lg-J@W3=K
I,EBR?@=O+ce.W=H(ZF4Zd#A8O99QK4[VEW\,N<GGH-GGb95I(+,FEga@K7R)WZJ
=6@LZC&PQQ82H:d)Y(&QeYXPWB8YU[2A):9gBX>N1(OR6&E-<OO?VEF)_PLZNS\9
S\]faYaZ:R.PE2\STKDZB_B.#ICa:OA<^10@T^XNfN#<::e,;40CL7I[BQL5?Sd,
Db<TKf.[T)XG,06JK-U;5cG=C&2e:.4[P)/KQ;9Eg<NYg[V._5eMG15d>H@O2?T?
,XHG]XWg,:M#M@#PC]]64H1DN8:B\aH/R2bN;;)NYKE<X[EHcaK>4^Z8AO<5V^+#
5SYE@8/>^IJ-F>2V#MO?(eH.YX=:?EU5@\ZYFD<CYC7-9MA755gHT8JcYb-d#&Ue
9Y@dC>cS#;&=L4NC@8D<8Q3EKaMANT+eL^)&LRBPg;ae;cH/a0Xe\a?HA[FR&=PZ
FOZ.fI9A.49(7fX.B[.AE1+<9.S[G54ONKZV];FYR(</_M0e&;Y#@-Ef)PCCVO(&
9]J28,^]-^N?)X#A,SXQ8+V#L>27Ea+<B&XUW)<<S>[B<90AC6<eQ)+K(bfAE3?T
O6IcLB_CeWW#-L/J\eNg,f+M-<>7+BaT+7=M@IG7@f\/VTB5M>aH#SEO@LH2Df;]
D&+aD3/S[XVHDS9JbJL1b?.7[7IE0-Qb+#W@KB#L3O6C@.4/=LPTX&E=Z_-_9B[]
2:f_@0XfTFP4[EP_5,?\C5JREJPTO<fW0],]NV6?SIf&a[DG.@c2:Yb&K,<N.faY
<HRa)LO/JZ.:QgZ_SSN2A56H^f;X1dYRYa9M//5eSeX^5MP1.P3e^cPCKSV?79S\
L\H89ZR#PXYX?IS(TWMbW.@b\0&c;Q6\G\.,+^172/cMA8:UY=S4[P)KZY/EfbU@
)-EFZ#X.042+T\75/.e/AVQd2,\PS(JCK7-T678f@A>gD#NF3(@?]aL5)=MU[9(b
30LN&XC(TZ4U2=[bU>>?.ESRCHYF^C4DW2PPWWDL\:f8?O>Q491=11BJ@T5RZ#fT
3:CQU+#:/@0]FP(cY@MPE8.YM4.57+2aKBc>Fa5V(FI<JEJ3dcQOQ#7UIC(0b2.8
]S/W@[\MQU?C=M[LV/a>P[Pc[Q]6:aKG8<PgW:=Y33c6>0F/8<4-(7+OV:2\)B.\
.cR/FKOd)c,L.)XF)QIJ5V_b<0I@abH1]+Q_-;4E8,GIU1f@b#c9^VCI9+MBg[eB
b1Bf#db^;5dgP@926^4/+:ATGWO_b9&.XVTDL8N\H7dU?c2W&]fd7EJHQ\>H,R,=
__/aAP9\BI=>?E<FN_2]GTZV,\9]c3eaWGUfPLY?OCe;NRK6T+^P7KSPMH,^d8MZ
NEGe0b1?<XR,d5e+??4M/5+7,\=K];g7H(6FIH+J7gMI+#2+,,/?DA\+Za:N&MVR
aZ@0QGe_L9,EK;[0gALDT5A[L?Q\bE=XO@bUed?.Q5H7L@P>T,gf>4[=>53BZLIc
OA<Jfe4.ORdP1==@&g75SIcQK=g?(W381)XHB0X^?W9ZK1H)AQ?:J@4X+Fa@U.>E
4dQYFX0JETDZY&5)JCK>-PKY6a.,9AI^c3gaZ)+TOX[>.<@:)4.,&::MN?36JJ7G
RT^#5BY+QZ75&L[:YV)JV@9D?4@Af:)X>O+6FK&+gK=S@<6Xa>+3?g2,RHI-QQP<
La5+52TX-MU9TVQ5=X?Zf+SbXUf>6Y?E0K[)eJ=eb8D4dYF4-Hd>R05;DB[GL?b(
KNO2aU95LaA-.#2Hd6FY;0PfVVF:&Yc&\:&JLI60,((G[2RY]><6Q+YM_R]2M1g:
2-TNK8cBM4GeZ\^H?V<S-.,GQ;>@[KgC#T8f)C\/g5a/B?9cB5<A296GUe?2N9XW
dNM8dZ&4?64?_BC]V0_2W=^T&@.ZE1H5&\UB#\/B\WX2OLFSfFIYJ?K;<#)R:X&-
D0H).:.NY-&\#0cbYe2#T;5FTK[D2]X_aa3;_@M2(6/KfGO)S.KVN&HJ?YdVK?Z3
;)KWG_fcJ4QdMDL9/0aTV4^AVa1[]K1FK\+#3Y4S8K++9.7CSV6J<)F=ZO<&Ne>@
W.4CSeUbZ;3B\f&50],U8]ZeWST_<<cG.9N0I+5^B>gI?+e(TZSVGbWL1_E+NN,?
:BbffBO6gTeS5O<D=X^X\91GDaUIdZ7<KgT(FR^>Y=8BbV@fEVAWA1\Nc-QB_@gD
3bdIQ+R]g<WB8(V2947\8&_:QffdA:()/3AZ(LeXg_8cHP3^P^ZK(XOWfM?\HY=1
LIKZ=IJ0dOcH;3\CH?WKJ;QSD#_FZ;LF]L?TD\SXfYDb_WZTTbTI.D+8DHgO/?3-
^R_Z7Z-IXd,[e1-9S.3E@CI1:L(EPbJ]c>T]:17I/?7STU1Jd0GOgW&eP4KBfDUD
;3H40ceCM<JI.#>a;XO,4ULe&8S+19f?-eU;g32T?B)?B2)&,Zc0OADOK]/I[F>K
^f(HAa7+_((FG^AZaZ+g5)geQ9[.W@JTK/U)XbdI7RdJBLF)Dc=):;I[,<,F6^4.
8L:RN/=^>V8=;bbZLBaHPd&QT@WfKVDg14J2TUA(^9X@0O7#G&MS+e_]7gRUN:7=
JeC+F8JGZX\:Y9L4JN:2LKR(SI]f/>>_1X:R><YM?=bQJ)Z0)//F[K_WI(/0IV)>
Bf;FO1=2YT2QC;P<Dd9Lf8B)9#5TY)BIa=3]J[cIYKPI[Gaf)74.\,Q3Z:M,7)?G
MKBDEUCJd7\Y39QKM(3X\5K(AF?>d5)Cg]:\UeQ7=VBX#/,=[2_cM]dJIUP55A\-
E9QRL?M,J_-7/RFgf.,,I9D<GF(BO_G,0f]?:)S3IRa-JHCf7-P(e##\[=,OOg[/
[J_X-Y-_TDOW1S(LNM8B#9XOc_dTS-]ffY^<+89]\IYOPWH@#;CGf>Qf=5T59C#R
Q25PO?I>N-9)Y:QNJ;:HFZU;T-f>K^g:>92^Aa.=.d56A5FG+&>@7Qg).e;ba]CU
IZ1YCY1[S-?YYda)fW]7cD[?GD(U_,bZcE&\SI?<9985>^5<<[1SMM6D?T6SAd=/
::;a&.ccg>LQZ/8AZ+>8)ec]&OQ37(VMA&P^91JC.&L/J0Q_]#,&R.T8_,/Fb@2W
<b_65)(]:\GcSA_)eXbCP7:95Ig\3cAA9HHYE+^Y/#A#[A)XHa3Lg<+fCKL0J@L<
1XAB?2f4JGV?A?a[VcfTOM&[[@EI5FOe9UO9/523B#X1BJIMLa^#GgX[N7M6\[Ta
g/Y4PfI>GE7J;DT+(FIeQF;-B,La0+Ue?#JKGRUP[#4+>;e0GUQ;R\BeD-=&4+QU
G4VH#NDH)T^HCeB]NL7cOMdX;e;PP&U(fYKLHUFfC@3R6NY7USY:b<X]1\1P[:b#
bL4UTN;S7G3WYJJ.G1NGH)IPgg(6g5OIIfJN^J4A+B<9XI1[QTVPKLO9E.:VVS1U
\\W1g8E0=2eVRHE\9<LSHdHa:Eb_);L#;G_12NIA=^>C<:XPD#LRg.&G-TU#]+GD
U<WTZF,D5]GcZ9SYcc/?OW?LBG6)Ve@&\c,US<Ae>7:IK/-L-EP]?,?_0aJ2J,PS
8.A,IL6#WDSB7K&2d6EMCKBOL&FeS?C>O[)Ja&<eF1a9W/3>G]a3,86Z:#,fL?Y8
IE7cf#7\c>+3^7IOAW<(C>Ve>6e9OMKCM(@?.T3Q<G?50eL[0ZZWYS+2]KO>4Z1f
O/cM1,GA_T/LGf8&OX^6ecZ&E=F8\</f,B/HZ:dg7aV9Rg<.8\V/FcK_QS:.7g-B
dTDg+F84@WQbTU[70(#fTOXXU\E3:W<,e4SN[3B6Z(?)1?GHb5ZJ//e]YW&VQLU@
H49G7:@&&UX;I??_f#&@J6T5M;U/R>Z<<#GO&IVVTS</)U.(cQIfRZCSNP8D@8J_
1?1/5+GV0K?b7DMFfW)(2WAFP5ebDFBD_8dVAHd8((-KWL:@AR##aT(8]0-_3,Z/
HJB1D]BKc/g,gTT:b&RD/\XE(U@O,A4C>0GeET5PX8D^N_1RcaJ@^_9WSC?TI1)H
002aFaA+9U0_&@AZ+gP?.7d..EdEVN+)^):)L@S-(WT=-P2M40]g9)f]IW91+N-0
-X?fdKH\Mgb0_4@@(?=N_6gcf_X(9EH[g?e>\6=cBYP0]a@TBFYG=L2W[ZR\f(DX
D#,MaUUU71RHE-HZW\_YPK?=1JcEB=4?U)Wc:-:^<g(>c+??2_Bd?+(Y+Y=])JP.
THgK.-VF.LJ0,Z1:3CR;8I(-@Ld4H9Tb\/dV:\T;N&1T:fMZUbOM,@X:MW?F,)^O
ccZIS8SI5f3]V\(:]DU&fa-PP)[WeMQ6O=aAIL4O#92GG40UR?7RZ(OCKDK^OX,d
7CM4G/_U]@@CM@b/D+S?2\+4_DF-Ub[1EfECL<Y.;KA378HS#&P;K^PKGd9a3O7V
DR_S([6[/C\dXXCMX&5=8QS/H^=P]ZHQJY1-RGAQ6gO0[^+X)VO#(#J-K5Z;7P:G
7BQQ[D<#KCQcDHI&_>/&^9;6YRC0<W38.;XTS7H11_C?D-H=OS3=JOA(KTH8<b5J
5)IgT1^88K2dQ#G)(U5g0P6GFSd3RF/LAGHE<Z\X@B+B2Te]#2[0Y,/WV]]f^AV<
GbbBY^DP@)dB.XMK&2eW</gc&F1S(^dCI#@<(#;]GV.=f?/I^+Jf)@/WK$
`endprotected

`protected
Y26^RFL65JG^@_Te@;E];G-;MJXO.C+CO6_)[&OKY:[R9JEKb)5(.)<<BMOXPB-]
CMFPF+[U?XP,)R._,#NOQUg42;;NQZQX9$
`endprotected

//vcs_lic_vip_protect
  `protected
C//7H;Df[P&FHX:-7;KBQD^/<UQMY<:afP^G(A8M@5Ed@egcP(OK-(VV7bg82<D.
IU4.VES)2I,:QMX&)9Z2[W,1[I\]D<PV;Jd\NaA#@4JeAF[._E/C[b2a7_>=aE_M
42>QZY&ab14Q]X.@ULNc5_Z,_[-TJ(QX;PbaZ.?W;dV7?4U_)^EEK_2-LUUW9\3B
&eA)S\R?:;O\<+,_D-cJZ.FLNFHQR96\VPK+7ZZV)\a^WV3A1:[8V8Va0[?VIf4^
Ge/B/B5-(Xb,YBCTQ&?6#S8=N@,H/^)87gfW4=;7M9Ob+7=e<B;EU45JVKV2eeKb
.>cf;gcYAIN1D)5Hf3ff;d/JVS9G2Bg2.^Q<]EbDRY1YdZH?HU<<dU#+FYd_94>Q
T)1=897dDT22Df]PV_LBC[U0d+Odc?@7,U>0UQ[ME+eMF^/3=+eRKNI2@JRE#\^f
.T-@L1g-\\7=1gDM932#,/Kf@B/c\a9gS-;gK[:]R4&W-48cD^-aWRfFGQ0fAQ]+
Dbb)3a[9.7eRN+J&g><.?0P^F1Q1&EGI48?F(N4Y-X;bZMA&,]fLZYPV6X3L7U\b
H_AE:FbC_+0_MA=_b_T\(,/TQ+4M_fI,JAc1J^[)=42];=^)^I6d+_2@=(,^KWGM
MdF^/N/G)9ER#@:de+b;/=gEaODNS_Q>GEfNY.CSVb;]MK2&U_4He-Y^,A58X?G2
&+4:a]7Yf?#[L]Y1><TU:H8HCf<O0?WZ(g[W#]Y.?PJB(_A(&a.7ZGW]E7LWVQE^
61+CQ:E.;5DaG@K>:[R/Uga\RO^OZ2-)6:?X+<TWS#ZA5.(FQ1D]ceXDOCOT3P>D
BbdEE]YY,GLR3D;WLREa@Qa,F0EMKIXb-7.T=fUV50ggJf;&/N,WLaF4OUR:XggZ
b3-I@M^BfAE83GK2].U^?fE&ReK5H/Y3U4>ZJE1fSX4RMRK9ZLIGMbDT.7_QEC/1
0P)626C?f(S(5S&=<.(W;YMMK;B0?Z9\:CJ?#+g7=PK5IN-e1>01gR0fL;XNUPgZ
4+&LA?&_[[Dc^\ZcG4(a+U3/-U<T?]/EF@Y027f0\8&;gNPc(4bLe(HFTNWD>91c
dc9DB=JV5L^-6>eEE2KC.NRUUN3X,&.Q+.Td8D7GL-2DO1O2d.12W.+YBC#G0;GZ
P;-5Na5N#S?^P8E[F\;)+],c7dSO8g[961-Q:bM)9)f0FUbZRIVPOX3PY0:63Kf[
R=K=Z[:aNg@a-]#e;57FMTT;W57STTg/5RXJ3fL6+50Z2[_>(8Id4@g6;?XKJYW;
&\W(f[eE](\>DZbR]6G_\4d3P(S;F,CA9:)+4C#>UGRc##/cbUW)&GEJVNB62#MQ
)dJ\-H]fcX6UEF/#1YF5>C-NfUEU0eTFb\.b.OW<K6\_H_.::E14cM))9K/I2fH9
0)-__^E4Pd?GY0FFMPbg-EU?eXFgW.g,/4e+6gE6Q?2>+Gef=B=_(8\\4^TEXXN#
(Hf^IH7f#-g;BNT=67c/EJV<Y7Nc44a8M+?QV[2Id3#.Z^X=aZFe3)6g:QB)736Q
g11PTHL[NC7;^Q=2/Cd8P(8I1^FDOgWTA(/++&]&e[C/E\6aLQ_XXaC-_fRH4-K2
=#HE?f)Q.#B57NLNU4>JJJSON8@aTIVY_-Tg>D3^>E1]AFbCRX]<c?#L=\YZ4))E
_,[,^ZeTS9#>73[T#fbM(<7@G#5+O^B+aYW_9PfY7/XYSCUC/8OF^^&4eP;Q&Ng6
J4L#4#=\Z<,NEY#\d>9f@3V#[>D.+4#;H+:?D:N1=OfJJ+8O8#21e5d?#=,F<_;:
faBPZ,T5cTQ,8_HA_#X@.(H9HfU<V\JE&@L0N8;\7@\c7)J2T\=GU@@(ETCe+O^b
-00OP\S8RD6,-:B/I)cW4]#V,(4U6STaCE</>I^abP,X:T0)L;:@/FS<@Cb?XVe5
CTZ[-dPQH0--:Yb4Q[P5\J,:[ITN/<XOH=a4[=a2U=BOCUd,cc:fa8FX/-,eY.L?
P,9d^+fW9F4CWaHVSX)Y)gRVI<7W^LK<G8UeG.?<=I,CVG#/W0(0ZB5?QJaA,?U+
E\IbW.URI[L07eV+ZA4FL6+gf/YC:R(TL1Q@=]CbBD8PC_Z1:+((HD-R@QB?a3?6
ebO+20E8IX(C/F@3.S5V:F7A1<GC.B&^=feS@91?A/5?<Y.=VLI(<9JA/B-KBQ#4
c62A5LG\CY_OFJKZ0JL<\<6ddBX\1TGS;4a\aeaWAGK:_TMKe3;47?:OI.350,S<
=#S4F+W#_JD:Y/E;J]1PC55c]-&:PD7(U?Hf1>NS5=N\J9+#E@A1VG.R.(QO)E@-
>aW5-JJ.0DZC-9b(CHJ9][46CQY#8:f3(6,)K#Jda:>9YJS/f=NM@]4S+I@-6IHc
#KXeUL6g^14&BYT[bUAQS;_-BI9;,>4[KDEe?(T/Ec3<K1RXBP#JCPI1baJ;\+M&
VD8Y)TPRBA^.?#K>-a>\36KEXAJ&>0\Bg[dVRc0I\_./+3792FZ9A6IJ-^N,U_;3
Q]Ac@>;:OUAdaf@d56O;aM<9e75UPDAMNgbfb6<P.Z-2]B.;99eN.aEN>U-FUKU&
)Gg(1<L0@)B^5\L]5Y;)PZ9B+J9HO8Z\X\#ceV41(SR50d\^_eJ>_Wd8(@7TaO>\
/TF\AaI7)8Z2D-2GGIQJc=6O=:SScFY]\;QfY-8A:98<,,D9JPeM0:N7HJ&c.Pf]
_bJA&^X@\HFNe?b2W),:H)1#=EfW9]U+-D3gRfHGg([-fOb87.60,<W:(41++a#]
.RL]<2I-2E;FBO97Y:UJ049NS^GS@>K;FN;5[JM/)6#Z@,GG)2]@AE4O].7^?=L.
)#=Oa;d7_[R<Jd=1F]RZ6M-bNX;N@c@;:<^)Q7?CF]F<S3,K:2KE,X?4ZbS3\E]3
=OaS#8BZ^H7e[2\A>GO\(]7#RbHR&4(O2PF+_7VHN?7F@WAB135C^5CVD\Z^dT0+
Xae5V\::TS\08#aOea&C=R;7M#V8UG7_fL-6L(AgRT]XERP0HY.H5dE/CL,G0.DM
SHVab-0MOf-^:EGeD@X^K]-=XS<F>Y\Z/6@V2P(]#78.eEd3deg1G5@)#055_Ib/
@T6TGJ#\5XDSO]^I)feQ-bH>+_UIc.UBIZ?BFR/B(]RIf>&Z^\9OQ/B&>6PKT.EU
TW5O_NC9.35X:@0/EA5A(F)a(aF,,Y_1g=#UOM6cb1Y=5+TgEeR\b1Efc/6J5DF<
H>WWEDF:Ude_<]6&QK[C9O-P/Cd;XH7)8+DZ?Q_(:[&ZJ8V-FGD1=<EJ.dDDH<]W
XZ#4Ag2;NAOc_;7;0LNd(#\Y2T,(1b/=)PIM^g/L+@M\VZd<Wc7R(aC24[gU\0G\
OcIA@1[3E,:#ddXRG4G/Nc>6B8G+C(F3.-g(\XRCFg-8>(d>D^B4@VYT.da]6^.3
bAA9DTgV>LD=a54eP?-J\aJeNc.],cBRM-KN+9<T:VX8TdS.U\E];L\,&X0bBN#:
]C&Wa&ED37K.bJJ\TL?Ue&WTKP<EP?NB&L:W28..SY9&)GX(?,U&_(0]7LP1;\g#
0LEe7:48LTR.eP<S][FE4(MUOT\gLX?E1BeMB7JB4<177,(D8H:b+^L.IM+F5YT1
dDODH-6G<)-K6.6+0d(GT]\K-3cO+d?IEFIY,[.</1P38;P92]H[\/(&R#D0_Kb[
DZZ=:F?T\W(4YggT\_OfRA.eD+SWFX35(^6&[=[N3a>NaKS]^C:gQV,:F^\cc2&S
dB#ICDCSS+M_UWcA+38MDRVFC#IMU@TN80A8DN2E/_6NGNHMcUUaOO?aBa2SU;/7
7/X&aOg7:5TJ+0@+4I]V=/9dc=(51ODFc6P;KZXG470]E>2U\4c58(?&2_]6c&MW
5bTV3/(YFI1D;UUfL79bO-1UF<[5NJ?,]4&fda-P/7LUBbZXDH9ZGK661cW<VAYL
0K8R1(0AWe]W8GTGWfS6(<BZa,g@P>6-gR7TH3G)K-?[6bQ+3Nf_>7-B[:NK3-Ib
4^dRDcD\S0:DD/@9Hb<Lf^?76-R]5a&RF7BeaU[O;Hd-[d47N);,+)Z4?SA/aC14
HSNBKC1I?M3Efc:6:,&6AQS]S/]AYLMB_N3aPVK(^_O)-2ZgRfe,Q]L?6B;+-H(]
TJ.H50:X2bN=Q4U@J\^R]>8TgA[CJ[;f68-:W3<fXg)85U:gd23;g5,WYPF>KcWL
5X-:S\E#S5:60.?A#.F;S;M1O+P6DGg.]a7GK9T)WTfN9HV>8e6N(@P171ZUa5+&
ff1,>(c21S:ZIc,3^eZ54#a8@c&T-CG/7X:(A;(EA,7gI^@6NJJca+-#=&MV.FfS
g/Y1HC)J&:],TW=WGQC8:1-2/bYcd_=Y7:()8YY5E0aaTgB&g92:N+fG>QCO+X5B
a</WQQ[U-W#O+dP.c@g[8bdYO;1@b4,g_;8cK8L,(FWL/<2R2P-FfQ8OaY:#S[fR
O0G03=bSCES.T0)Ie^)_M@KcAX4_/:;EWIQ&-Q=R7-+V.=:b0<?MAdX[F_/MXa]\
g^<GNOF,e#H3&P7F-BbH<?7)(#DY6^,79M3#N-3EGWIO#7LE)G&EI)K;g5=]5QSV
/PZB1F[c]L?TTEJ2,C^J\<48J;H6=41T[bZfJb]BU/BQEZ)?\ACVJ:OB/&J@<cI@
6<-FG@_/]/]\,TLI]:>>YJF/YC>4eXF+eB1IS(b&[)6&2TSWfFD@e@^3&[SfPFbW
DZb_eB+Z\E_Q2TS#D+S;F#;H3B([XL\Q+5b-?4#fAJU=aY)2<U<<IQRL_VA]WO(c
BEG,>bL&ZQB^a-6W_06?)J0X-MW0[HRH/&EeCAHZ#&&E1TMacJ=gT3J-Xc=9dI\B
GW7\PacDS5/GLP(:ADgLCeBHK=C1QUTHa[Od6b#;W+dEH.<JX@3<e;+L=FT<O-R8
/<,b(/gLTRLGC4LL\3gI,?0/+>):X]\C0953[J=-]J8K\QM>4T&A:f7:A5CO3DP5
_-&Ub#?SX=L[WK]2fDS.QTFU[b^G_)&&32U(g2CPN#^f>8JE\X</C3\?QU99YEb3
GY7_T_Y=QA4=fW9D^EC1aHBW)A(PH_=N?QL+P<ZT7\2=YE1R&C(a,[-FF+R@CKK4
XF22#H>9W]LegAU&:OJ<^[bgOJXNCI6]D4<E5B7P_gc\7K[7N@f301=-RHA[>&9D
c-U[,9/J>e<TF#]c^JB]^T@.6C2+,KOPF\C7DTYWOPENRf]YA,TU=33<+35_8dET
XF0T3b@gT)I.)VK16GGd#[2L+eM5[V4QKN,J4,9;CfIT4^\ZGUU7S>R5&HULT@5/
);eGXDa+/)Y-2OGg(0Ia&Fg:-^^b3cJeffE<P\1K27+O96CZV#,9<XdBOR8-)-dC
R8gC\AF:/.4,#YEFScE(OE3f#\;Fb8IJg+1-ef/I=<+VS,;HV.#42@&5>R:V1GTD
]==/V4&XITa/QdgL.HfV-GaWe=.2[_eS./VfWRRcJN]f>(9B&XW=R^]gXZ)K6\fS
TbBg.IaROKE2VK(-Og9a2c5141Q0BIA-7L40FW2]NKaTS=.)JHO^H-(5[]\0c/:-
>(W3K#7EW0J\?/IK>,:PF:?V54-_TC9g[b.>/Wb])>A_1;Xg/^B,PS&;,_/562W>
&&X@A61MJK2QcQ\9:9GB@BJFM-U61OHL>-_dJ=7/[3__;+DXPOB@2f1OBYa;EHB&
#X)V4UM>:gJ[)SAQWTB2Z>U1GQM#K\:M,R9)C&9^M.>,T9&:E<dP?3K5\4#d0bTb
-_YL_X3Gb(UY5S+HJcR(-T@U\D1?#[gOKRSZ4c##YF>)IY^BRW1P4_ELT-,W[a8Z
E3I=Q<KJA=GC>@6=@\.S74MXP.OR7c<W;Y&8_39=^;3)1TG;/fF)Y/ZW8^J;X&L]
B]c,/^;Q;I0VFbB:Rf:MXJ,IeMK7Y.B?QcddGRPTWe.3_^N1Z?DQ\;5+\XE94#-<
I=MfS\RI6BNUg(/-&9R:1R?,GTCV:MGB];;Fc?=<)f.#>3T]<1,QQ7_YFNY#NO2e
;763U(JK:=c1gYUK_Y&-OUbag.acJHG72[V-F/Y5PBb_;)BUb>c:_KS7(:/+/DFa
./>X3<V2<JB>QSN3@K.O;dcCMfE-<4&?+SMO,E@/<B)^dgf,f1^M:CJ??gS\QO.4
=0a3?X)_@EaKC]T??Bc-KHY0C/GG9O@8L[.&a&M?[-V)\[^J-#OYHbH[a(IM7U6a
U1<HIV>EFE<0]1.5(Za>@>(Wgd7HHS6QX[MeY\-,5P5BRDQ#g[LS^\PBdCH?d><e
/EM.DT5[b(<^b/#)O/5(XfN<f75UG&[/?]H]H?X)L.f/[FaJT(efd?8PTc&#8_@:
/<D[gd=_V3B-_SG7F)S(S+,6,aDM2)U\#PJgRX:21Fb>W3(1OSMZW?V6bWf^_@6&
G(8\1WDb(=X#D4#A,YDDcg7SIBJKLT_RQW:Z(/M8L>cG;]+UQ4\/2>^Y?fbLC>fC
HK#V/QV7<P2E.d8OcI?=8(fbYQ@]H8PfE0JMdJ<>29A-a(J^fX^HC_^a>(-1PG8.
JHTS2JJJ+e^].T6e&G/II&d)bA9f,W,\B61c2J5NbBCD#FaPDY8:B)9UM=Y0)RN>
_KD:MY3NPbKVQ1:e1M0J@+OS>[,6O7X2QT?0;4JU:,,MeP5PY9X&R,[V]E>^COYW
gD1&YN^V9Z/ML&S5W=3&2S1][eI@gd2CM@.V(\+g0]fB8C/XaJLR)W2LJLZT6<f+
:)\<@P,SB82Z-8X[2I]QM,+SR^?#d+/)X1&^<(BSeO-PE3,cNR9.JLeR/699M=ZW
1-5CV.LW>NC8UU3W]&##)7\0?V^1DL=W..VA76#=<I1>W15_N)fVIRHcNEb:[9K=
,5Q5M1[LK,c+LB@;D\/,cJAegO:]^P&&J21?@UOC9,dH2(98UDW&d#O=@ffcN2&)
0.6XFXbRW39eR[J9=5<8-K;X#=H+]N;LI&,>:S/(2._@YXSFVWB2b,-6W-fL6@SN
VVbbPF6b9B035T.8C@b(EK7O7dY)?+=aa.=DaZ^XO+_E0J)C3-V0P93R=7E-d);3
A-c>b86@eVHWM0(cM1C]B88Y49=f=PIVZ/3cd=#=IP.]g7]W^]/AJH[0N:M1F4BQ
0]=add#GS.;&+.],6BVWM3FS\A?2g8#.RRa/4E05,V3[&BgO4fO;7(;EJM:K,#&=
I2dS?=dI^e3][DHSBFJW)5/ZH4/g>b.KTIeC(+>>dM_MUdCFB?RF<?N9N6W6YP1O
V#/ENaHGGd]Kgc>2eF^Pa;a4b2-S7L&HEEX(1c:JZ>\LH>V,VN=?>[&Z46R[8D1]
W(&IZ-9EgGQSODee=Za/\2IX;4(MT9-4XDT\_]^L[CDNRR:=\2gLJ;ZQ?]9QCUDG
V6QNL62L,6IW_(Z=HI)DU:=HaAgPM8+K)R9\^YPD#=Q0CdAVNRJ+/T<(1Wd8e^Pd
-,S4Gd1=9f4WR&R&Q0g1HgCC1SgGFI<_gP/fN19ALJQ:PJS35Z&/6,H5R4TL(PJE
eI1&@)S;@C0b>+I:DFOM?4A\[a58^a_&^7YVY@J)Y5)a\J>-R+_(L_Y(O3TO7IYB
Z;@>U8>.Y3.HOIXe\_9de32(e&520<09FI.WGbA-?AR3d,974K3C4I5-E3e[U+CM
]=+E^c1<3KNFCeUdEZE:]3bf/=?#GXE:GNHF5b:LFf>U#+f]X1#.W=1-K-.SJ\c5
S@Y(MKA<@1=/.>cD4FB5_&Cb_PL.O24AdM/-C,WP8cAQ_<aS_9WSa9Mf>TO-749d
61FY7.c>3]fCTZRe[GIW9bdK<+gVQ5F)LHg2>=-_bW9,3V^baec&]3YD@_3)_M3N
>+OA-J2bPM:9aP]M_OML8.W?E@TB@TGF]VA,IJ9gSVCJ:a#0MH1?Z7<4KZ-HSSL@
f-b0DCBKNN82DUaQH@TWc\)S_6T,,aD(a<A[DZI39VcU/@QAQ_.1PA45Od-/c#HG
W-3Vb@bEJ\3BO.7c2B(<4^bf<8T0/?MMA+^_L6>#)OE,2]YT>NMMFKc9XS>Vf(DF
aEOQRXRR^.ZC:+g@:gAc0SBfa3(L43.(.e&G?N1R#b.Pa^bILPHI);5+S](1G3[O
A_Q6Dc+\9(eg&M_]G2L7/\1[P.1d8/CYH9g7FRD)6[dRC:R(GcP^@2K^4RF]E7S\
Y,(>Q<7X,?cV=-^9D^^=:+SV[E]1c3cX6Q@MQ7-7b\SV/>,94/.SFeO8]^K7.UKT
J#64)gP(\:<f4O,DCZ71VWJ@(.ECc(QHZ/B#WUL02\\UYX3;(F4N):7(IFa+8,K7
N<I-)Q<ZI?UG((7:M^f\OO2709<0GU]d(^R(<X/\eQXA89351cOUL-O#H(<_/XSd
YR_)<TBdNIaML1M\6B)T3G.^0O0#71Z_d+B4@dSV^6K7CE6F/W^\g9_IE-3ad2V6
?&9Je=#\/II]F7fN74RE@>YgA]QYH8GKYO:8+XZbLWa@fXJ^C.DOO3X=F33I2Af)
I?XOJ2V[_+NFQO4FDFUO@3,[E3)-W8RAO]GUAbDO6:/;H9WGI<LJHF63cV\B00F-
b?)V?Z,eV^#9=0;X<]Q>7+#G_2>1OS2QB.1[?&>d\2AQa<SAOJV)V=.=cc53KBE5
?_UgBF5gGXBWF?07LP[d0P,](Kg4T33YacI?YURLWeEc)7aR>NNN78&Pc:KI;&Lb
dB[+BV.N/,WI,Y^)VIGdgXO:d>cKWg1,?<M_Y:56L>c,^;8_S^Fgd?Bb:.DbYHfb
.AAR1dDUQ7=7c;bO.C_L=C<RC=e.=bZPIPb\eV<@@0.?.1-_7[IEdO0@bVO0TU3T
5ZWUaU8CU&;A8Y),TBa5,+2,#;[ZH(]@WYYW,8M06288:JS7)#;4>[ZK?5=4\ZM=
HaJVUQW4bY6#]=-.a4.@:=^,0(fNG=I4K:@Y=[d_4XKDM5\_?8gCD]SDd0+7BNAH
7]1?00DM5O01>B+9]LKCX<H\/IH,ATe2c.1][G+PMU[9GSd)4c:\Eeg-Z,F+8D7-
T([^B0<FDId_X^\b=6]S5(ES/N:8\V_ND(,^)aU25@/[N6]<#;7E#7(FQ4<c=;?\
:^&b=TRV,RfJ/gQ;WH,7NRKfZ\:-NJgHW+M<@\OIBX+QE5Q^K+[N_#@dKWB8A\2_
N4\6bBU0G[(ZC#]P,PM)JFWC1H[Z2?1>?G/e-bWeACUHXC7c7YcBDMZgNDC2.#,.
]\\\H9?#(2IDXT/J\V34:b7Kc.P&_)MC6dRL_JF(.P]SeNG>/-1ZU/H#&O/OA;7]
E-)?)X/a3Ad.<3ENe^Ecg5;4\[3_f;FP[SZW5@<L0/Ee]ZgAGCT[EUc+>bQLS^f7
CJ)g,[:J9>]1EZ@D98_(3NK-29R6gKVWLMPP-):H3/@@F(I=>)\f&c[Q913=8Q1d
ObD,>A^1N8(QZUSZgf@^:g0K36C,Scf@(LN<DVP+HPNEX)Z.5T]9;YT9^dI;54U1
g6SPPDc1MM0)3B3#VIEZC\-,GAe-eg3Z#O118?dF#)PXQ9E/+93YT^egDA#L67_+
8YQ9GRNNY27S^B>^\T^SEB[TU1_U3K2.)\^?4a#J.6Ha66O(ZaRc.RH>H4G8H(U]
Z<#RbH4e&05d\6VD8STC)V,QAU>UKQKLBe>cOg3:_1gSC+D9<QBH,&WU-Q0W/Q^g
B#;>+HKW()24aSRG(;D/K=?H-J/2N=7[7HZHGVVRASd0GK7Gf0C19e6#(1L<6BBU
HcLDYA]E6=ENQKOB_N2S(;eIdNAC?0bSQE1K,1H:==E^.J&HIWa3VZb5B4TO,6GZ
+QPE?O/_S]/Z>TLcDD+N:07b>;[(LA^G2D@a7))Pc3.3<@Za1K]WA@+=PRE?K)JU
:\H5W?c2P0V\gA7gO8-_W]SE5;JeEQ/D;9U6SV3fZ?3\]R/PZ4RYJ2&(/STK?VRL
5V=>_@#+=US)?DMR3NO(XO?UFMU^gZ_49T=-]91547KbF&#c(0c-=XM2L;SX0TM1
)bJM\dGcP)PH/Hf.8/A1Ic2WL(<0#f25Ue3)2+3#d?HOD5DJB6QVJ;NXZ9aG9,E&
^Qgf(6\^^VcEdUd093G>XQZ<3-.I#I@:=<SVR#e=^DWT(#8?U6=XH8<?g?0OR6;)
(V2E58f,X^g#/952cPAULS+FIHg8MTPSRO@)NE7d_.eJ+^aB&_?N#2#f2Uc<W=P3
LSS);_gKF(+.UQJVY.JJ/9MQdBGg\ISO56/\]0b6-cERE2fMT2#C-V#]]7Ma[E^/
]MHJY:PIHcc3L_JQJQbR,_9RN_,OTf+1.3-e=dX5RT)V-Jf>b/]9R@.UUOP8EBE1
_;eL1L+9BU/g;JQE/ETQa=80\WQDBSBVEOaF5Y_,PU)1YGEfO\N\a]FV8+X@@3D[
bD#e,MB(A8FXZa)NR<OFQR\<.Q/0[PM6]=LIG.T;(X9&NDHAVfG8FD+;JD>AV7=a
63>A&@dYECf3S-/)QZ6BL5PS9I&5P\@\2e-RSfX9Qb,a^&(M4bW24Ve5NB#S78I(
R7X,f;eD@\IDEIQ.))b=PT<DcE;QC>+WOQL\S-PZc#CX85KN#)9LTDMMd[W1O6S)
5#F@,I9@/_H;+dg+V>ZIPe(cR#@/B><CfK2(86/_+1:-X=6DZFNY&LMPARV\RO,d
GWgaEbSf8GH[FE?E_AW6e6Bg2K9ZDA?0:ELI^QWPPIa:[d^?9aEFC]dE5H6=N\fA
;d+=^\&gM>.WCFcP.+FU+a8LPS<df05aUB?]I-K30CQc.^8SAE^7bAK+?84T:07J
^MF(:)P3N)E<ZE/8REf<[b2GR->13TWIEdO.OP9Xe.BOLIgBEKJ)>]E;:,gI<d+F
V>0.1^L+YDD7?&)0Q@??BO^IJ1:BK&>CXL7QQGNC/<2?5.^>,?1?(KR5Hb[X&#(Q
faW-V+_L3e>:b+=eX0EdZ45WGQfEX3YM2H/JS&T@\e?N(M9>8K86Z5ADSXa1AOT0
XT^;TAY_GW,8K6KDKU.EW>XOEND214-Xd++Uc]E/[dK4g:U_JOTP_eO(TQRH2#-e
+b^BRQ@Z7Z,<1P^R]R?@Y)e<NUL)V#/7D70.TQB36_>Yf<;SD,bM\^JIIO6)CdLA
9<:GT/.@[P.&VAXOJ;)H/D/LQPMQWUCZR>.YA\JO0<bd.8[IK^N/<M96[_D:2&;)
0&EL_,fIZFANf@Ce33DGC#(ZT8ed4R0H48Y@@cXebPJVKEX5a<&BN2RW9U&:+\M6
cM.S/2&:X_3-AgN:&aZA;>b9#WF[#AF69P7A74F0NLK6L8\NOg/=#-(M2J9b=NYg
CN(_8D+H39/(I#?2@Ogb&I/:]-Of/N0RBb=D7B.4ZWODZ^,5#(_R.(V)D9@(bVJ_
=f^V(/GPFK2X8?F3/LN1SWY4:W<C?d39:Q^5]::\LPS:MCWd28LMa(;,MT6;E0L;
DP5>Ea6:[E;S__Kg/G#cYObgaQbEGf-OI\5_4M&Ug:AA?S2;X3=S_V-Y4PQCg^,X
;,O<UICdEL3)L.8@.(.A5YP65CLcCFd0^(6)3L9XIcBb[<)5SIGd@2LQH6Q;b9K0
f:7(GWVecZ;S?50ZXED))f75:Q^]M<L#ZEUc2?]<?g-T+=T153RD-88?(&.@;Lg:
E?#.c;&C@-JKH:TQEAI:_B?7TNZW&X/(a;_L>GL]@S=L1/QS3O/WXF9,PBZf)34M
]2[-P7V6ebN-;:4[.LTL(c\2[@?QPQ058&\H0Z2LeF+#fM-5KE01BI&W3DG3X8X/
]W22[()TCC^.^M+(IfEMQ&C(QJZOC<&_1A6P(H@g+42V+R8/=BLM\\.A7M/b1)D:
MR[ZX81a<>0OKPR+YX@-P(L<.<DOED1XD=7g_8;2fbQ5IbWPW\=f03?#aXb(H/;4
B8[3?LJ-OBYJ._99V/Mgf(-U?N0;fdBS\FHPQG+0=6XD\(.PUF4b_fQ7DcLY<?:[
]ffc?a>:6eY4_P8N&cMW-OJ_,=2-[4/+IQ&5?(_8cDJ3.J(73/8b_RBOG[L89#U4
:eV2QaA?B7[1f[A1O5F&\OSDIZN@ZM2CfEg?RPc91A@H65/PB&gN_S.AXF^aGGQW
?LUR.bF=4+gB^dKY(4C[CJeA4ZB;/:0@Zd237<1E-_]K4M0fb5a=8:<<C@6V&5A^
F<HE^@^RB]O=fUSK_=2\b#&:?62>eJY&MJ.J9ZOZ>YCg\-^+G;(1/;,:FVg/\74g
WEVYR-<[0Nf8.GSKL)USO3^]V<g];\3Ra]IY_O6ZZ]IRE4V3g)[=7KK#1MB+KFP,
BP8CGDTTOW5G+[d8O>GHGW@STfY73E+JEA=-f9Ef>ZR(APMG<VYHGW_.[>U^fc_M
@GHQdM#@<N-G_P<c4D^X7U21H4:a:7Q@FP&2GWY5)dRgC_^[&P]\\.Q)9B-_&-a)
+A^f9F;#3Va-bgbPX>_@J?#GI)d8OLXJ1]MZUW;FY(,&GNd1(^94D-b5Q7)QE/KG
)4b:OSN3G,1=]J1dO+QE;=)bT8U,MZ>PFd6TQFGc,WO^>P_N7=gQ?eIH)#60g>[,
Z^49^7M\5.YW-4U9TDJJfA#,b]Y9MD6X2=+ES.Tc@N_-D&/da/#90e)ZC;#Hgf);
#bI<YU_NY2V;d7cL082dXGHV,->adB?==]204PBXZ-Ac;[PA.dSC:GAB;[].^8K1
/_9+HXAB&6SMRZ^&PS.4&Ad>eLHN<FREP:=TF&eBT\]2[>?JLc?gQ[@WO?91ac.,
8-QeeUeTC;g>9^A,KH1WKBgWA5DO,N6c3,(]_0^(MM4.?26_e._acB+Jg[9W4C??
IS[OS]bKe5[egHN>R3b8+9gEE0PKFVD=;;I9&B(0MZRL[),KLCI6)/146.RJC3K_
UCa,6T#NT.8G3c4^WQbFCfCPagJA8Tc3CM=,^PU0B.4)Z(H3aN6F]:H.?KV);U2.
SWKY\C9bTHKeQ5))\&M,2>9)YE\X5F9ELIJPYU9WKLHS5O>RPF,RHB5P1#^148QO
>70RQVdF+f\<.L</Q?:J,YO&]9T2-0Y+QfU#X36g4011A06/SX7@NcHW9bZXJ7OY
.&GH-BNT@/5JBa2Z)eLWA:>CG/#5Te6;U@+fJ,>W17-0)4W9Xf3(2I#4.^.)PLg.
<+C+\9EGYHK\WE#CXF5)#KU,Z7CAOEPQ=(Ud4g2Z</ED>M=,J,:-GbEcIC[ZNC_8
g]e5XfDXg;EVI.[YS<8-6_B&.J\6+ZX(1>0VcH8dX20]Y.=F83=J1WEP?#0#IZbF
,12Y?H?X@/&?<</&==.Ee[/PLJQJ5OS#CW@;M;LAd-X708Ec<bPN?^J-69M&8eea
8RN02NCe5F8+0:?-K8V,VWJZa0d(M^d^HMdgO3M>.NJcP8AC.A>]8Z>K4=B3(VA6
T6]?B)^H-4>.CP6:NMaM>F:ER^.c>&28Xb6F=2HUW?PDOL@L0#\=bLd?\5ddIPaY
c=Bf+Tb&FS2e]1,.KIa>@);)AA_[119^WHARNdH1e2[F.fY1-&7-N.8WZ6_3##8U
.AHJ<-Q2D,IWJK&^8][&R@)=\H^@S<^<QGGF[;3G+GO#dcA>AbB,^MSG7Te42FLL
TM9<UY;RBPF&D+_Gf7L6BcTTPS^34RdKXZ\O)g7WX,+Q.(EBG76J&K^6;6F^\9WS
g-cZ:=eL=_6,#D8O+Dg/7&JMS?1:I.[+=A+4KaYD:03M6Ff-L?O[\eD.XBS<UL>Q
8=Z3?YR?<ODL95Fd\YdWV?<D-Ybc,@D:HU(.1Y?;.2-R,YF^,)E](F;.&#,H\4>L
KcJcR@?6<)VW2M^YQ4VM[8L\UX?DEa[L;?64bLc82(b#D@+dP\:aXD)Ub,=@.-=L
5W,gBJR^5LW1M;4BS@ec(7M856URJX(ZRBZJU\W@_^L=;L]7G<U7CC-/WYXgDNg&
W1-33cZ^c>JaY\F10+SPT\P&L-61(TMH52-;fEYE,Q1DMOQVF7L6NYF]MA\Zb_Q8
_ALIUNG:I.Mcf^^FLHO-O)MOF3CBEC-YB2=&RIM_,eDBIM83,(=;&U)d6DW&N0^R
eI?#0\c/R9B5>O=cG]Q7E?JbTZB;2cK0\+J6CfIA,MSg=g.9769XD+4DDXg=)M@9
9KX:AX0dBC<g,P#1f)/f&<M&0#&;6;cfO]f;Q)aLE6XN04-[Y6X(HV(^cZEH>=^1
=LV+OH^<3c]4;Q,d-+S<A(9#C=)eK#3S#dNL#]M/TS8^g01\TU?C3GH\]_[11J6Y
9Vg?21TTeQad&WVMU3gJc#4GKEc?BDWN.U-gB/ecXC=b@gfYc/PaHFLaLcdfU?/5
3J^M&OS::(Cc1E:bB#]E1:UH5bB-3]AT(:[P>)@@J+S/-:.EJ5M=@gN=Zc]ag+DE
;GSL?f&3+Ned8_b5HMWfIAfYaV&B8Y04dUA:S;Z0DA,a8P?YS20#B6c>6J^T58)/
V5JA5E[A@gQ5S^+YR9c=W1?b30Y#a+cE^VHV?=]?(JL;VE&K2?.6#T>.D6,I;\IR
aD7XggP[&.9c+A8ga^1&+ZefVJYV0MaQ7Z:f,@]2FDA#@4=ND;>_Y6=ED[0Gef6U
WIU]Ed@[b;QI5XVX9AOZ;9@0@VKAc.B:-F/,dOS^f)4P[NB#TGc5T=3@PeSd:GW<
8V#\d;YNV?AEbUe]P\AFUW6\U?EBFWFV(FL(N5NSbZf6(W@HIGPX^,E#GW60PS<;
8K5A937:Y)UZ3E<&17+X+TK/XeU4XT<_:=7XY(\Ba^MbEHLRU7A&fJ09+P<gM.O[
98RPAIA1fg/gF:>K_@H_\1a-6_[(T0OHB>&I^7?GFARB^?X<EV);XE7Q\FL(P9^2
24YD>W-;YAJ85D.?;6e&1KV^caZQDMT\NWX.[]DFOaD6N<:Ud+<+<9E,DNZY;Z91
<=UaPc5+dUF>;UD=9AF=E;&T#NU)0Y@e-)b3)E4g=7?QN2:,aFUD\7;1&;-7^=T4
1?K])=aI+Vg@UDVdYF#T[6Gc_@fG?^NQP<b^B)7T4HI,7E\(]WdRLZWJN>R#_8(,
7G3XYSU_L2[W4WXd_2,#WRf<L(2()@6a+Pf6/CN6c:QbPRTG#6>=#1LG\@2C\S\6
V4WG-:EICMPfIPT.57]a/+H[KB6YSAc7.RR7;V7J7U,NZc>\M&+RP1[W=WW?/BKJ
0CEWPBLdX)0I2RBL=W9P8V01@/E?-.AgE;(ggB#4JN=_M3?RJ7QHF[HYB/K3#_D@
XP6[QDNQ_EbWfFFIZQX<J/AVCP\d1W>QO:c)P00KC^bA-Y1bK7.6TOdH<gH<[6c4
KM,PM4d:C7HL1R;TMTMd:_Z+4EC-#Ic2@^/=A^DY6=4<9<L]4gVCG8F4c9a@&C.X
^b9)beY^_Q:S?0_;D<G;1H#,>ae;DWb:\6N>93L2TcQ+T2/R05dG=gIM@S]<DJ<W
N/d4@dY=+efe8d2RVQB4<-O9ZdBQI-4T(-bbUPH4FNS-3eH(,2[@VfPfL:HHZ^<c
R7(G4aNRS_6.7)+.WUb]8.B)IDc8f7eF_72AcI^8FeL(>8\V=RId;g63+Z5E9]^S
>XT-NB6=,H:I]+H@Y7:P0VDZe2JdbaJKe/Q9R9>AI8KeD.gU;BZ8[9Z6V2<?I2@-
TPY4e>D0<CQU(#P6Q:@YX=a6\3b,4MR[97LM7eX:gBETS_fG8,T7=D/B5,(&,R4=
)/#:Yd0c\?K3]&+c/;]?df49F6,MaP]:E3RND+9JW5Td(A4XeA/JRG0GRCGF7ND=
Kb-+;:)MQ?(63UEB8WR.M#c@Na=QE9YHCZc?IcM<dVQ>SY81:GH\?I#)dINFB;O+
U+Yd&UNK4]Zd1?QH[:-3>CV>MC>==/\(#G=AU07Le-\OD<F_63YD+gV<SK@0Fa)3
#ZLM+[aR:0/)#A_4cF/T89=ZH/dN#-TU75:9?4HI@-e1S7A@d&?BZ1EgQ+(cc;1g
-821bV)X^5TASY9@F4A,>^4N&I0d_@b;IE1=XT:)PQd5T@_CRRVI6#@b]O=-^LLT
52Dd2D_-<eH-O\G7F(-B.1MSN;CDf5)U>LBL[+)>&2]MTSLPH]ISXOecMR=+JN)7
#c>8G<W0PB9(VJBCQI+DcW]H4YHV7@])Y?Mc6_]F\E)#5E27dP^I0FVP\H6S/FEC
H<;@b(GgQ0JdH+<)B2W3QTEZ]3#7ReN8[4L\Y[3\9]PIea3bKCS2@+:YF209TIFc
5WCNOfDAZ]UYK?:)PRK\D^(FPNH25(ILcMGN>eLcM+R/4;Og24F5#L0I29F=Q.O[
0W09\@>)VM31DODR.H\c4V,5^/IUG8Y<W-#f57A+?KJ35YY^&M.,3KB,R[A9W-DO
D+]MDEXPQ(85<3>=F<^MV->XFHE#OI0g>(e0AZ4:H4TP.#eBW4PY1?/J5Lf&@H&R
^F14]8;/F)B:CO9eg01-/[5@D;O&+W.+P;dP0+81\H62WO[SR3[2J/3G,0S5aLT+
[FVJ\K&YWKBOSaPR(A:^4@)BJ\#B^?SM1fNTf;RK2RaeaK/96IKM1.1_/.]fV(FD
C>#T?/)@LW?-S_F;I[@(R;0DQ0W_JaCKS?@[<fAb7\9]XL&bO<5K;X-ZDYGgdW6O
aRVeLLVBMdKf)?O@d/^=+6g((Se62L1O1P546RUV_M=RO1fVQO[gQ/,.f]Lb)W<B
JXX=WMb5YPLJM)QBONda6(2MPVOP9RT>VK#AFY2/KTJ[=aES3I&RTQ@RceD7AOKf
U)NQ3=9_<R-c=LNCY.#FRFMdNY[(5NYO)bMMA[g:<YNRQ?3IB^>26b#:[06I9H/N
MDRL;-NOeSC[f86>^>VR+8+S-=U:E_8<eLPc\1[KY(;HL.R-RLR.&&Y>S8VP+^N9
Z>\;)4fXAZP?g=2VEXTMe,:QMKeN&GDB-@+J6+]37<>3;>EYO5gU2U:;OWRGTdFP
U;&]E0PTf>^53b9fYgZQXHd<DTYdG3b+ES;bG?1/b=DE;&J7/V76[Y6+(.\UFZ=N
YX(M:+),&O8_[g7>\QSOYQH]UK()fHD-dYIO,<G)^#SW)09U,R=]^d^7/GA=fC8K
ISLN1>L;>]?g=468V9B,5.?>?].GFW\IMBQcXb4RHOb&^>?^HQGYALNDXg4Ic0S=
_ZBC7)+ZgHH\IZ-_+R.0+Y4E)0+C06Pe3dL@IZ#R&;5CcI8aM9)Q;H59</3bU14O
H3P^HTIYJ,ZM@OM;/d+@C60+FCVL.(EdXEX8<Q^CWP_#39N0>KX5S3MN=(J,AHP?
W0PI-C(T8a0b-,BNd+WS.bGLW-@gBUHXM5+T[,a&5gEPG5YaV)b=?7Je#)f;c&RA
XT=MSHc:C\K95[:f^YW@N/+Z05<5^ad1;JDCJVdF<HFB1K,UKbM^7cMY\\+;gT\/
d3_K3VC#-3BeB2Ja8<eW/3LH)J[C+>ECES494Of1_JM&A_@Zd/?9]FE0bA0]RIaW
RD&@;LWEOXcM.c)4>51,SS1B)?f7UEUTRC+eKX,NLd>R-d9aV9K[a88M:gdGcC3[
T7<DRaBLV.K[eQVK4H9R,<B=;(0Z6M0)?V2=??Qc&P0>2eB(-\f_&7c2KK/D@V9S
-@=#+P5>0eU,92J9XcKMPH85Z=ZO18)ITBgL9^GP@#NTV657)<D&PS/6OSVf(fZY
=,&AY3QM?,bab6,,[O]]>Q>F@Q6Bc)FN\N0g-YTg^,1cN?EN:2NSa[.^&E&dNR7Q
KE-#M021N>FTff&)^?aO?-->aI8,c6N0J2f#@WScED2-cLZPLGLR>QeI3K)676=2
e54\I4[KXE,+C6@JT>^A7=E:J4^P)HA0=Y+\&-8;OJNO2LA0J<baR3.+(IA8#ecf
2]<aL.[0c<V&C_?Wc+YH)G^C5NCIbGNYA#2>g-+Y\\5d^A4-b[&)7NcOKEB?=cU9
1F>?FPPEbWd[X?U\KeZ_-HAWJ\;Wb5Rfd8A2B>c>?NL?YS0##_;R,f?2.QVHK]8fW$
`endprotected

`protected
<Y:9L@_I/=a]T>E.0cR&K.D:N;[7CWPe]DJeTU]AU[@3:BV0P/V86)BHIE>2SFCM
>R#[.(N6WfC]+$
`endprotected


//vcs_lic_vip_protect
  `protected
L_?f+B7.U&MIY_N>49@N-Yb[2VC_ZXZ:N86O=BT+-g[\K2:\]H_L.(5Rf4D&YY6d
7OEPC;^A&YLU.T^71]IXC&Q&9(cN#>C)AgN5ZQ:Cc9c)S\d7.91R.I;&)AdcOGTQ
W9?Z+5[bL[V6C3_/98?R<N3.N4M^AC@5(OAf7>9?.G-eMc3,_=0^4H)g&ZZcdQ(g
-]4O?#JZc1J=;K_>CKUN+<.[,6#NEY&^HFGd-^1LE90g[BI--V?)bYXfF2C(_.C+
ZW\Z[Z0,5T;IV([H\#F1WC]a18Q1\5)XgKYA@b2F^7,Y8G1aNM3,Rc[HU_S8?;5W
+@T5X9#ZD8>bWDCNJ\N8.b[.A,?\Ng?KO-YU8II[Z97.>U6B9E@4d^&;3cS#J3aD
=]56#aH@YZC^Q_f9^J=8=3IM+NL(5(D7CI5FX_(//)aS>::IR>Pb=aL+X7-SO07D
Y:;gagSgF/Lf^W?@L_;R4<)2Z#^a:IO\OAg4AFe4A1;1b.817c>DN^a:\W4^V_8X
cJLa@&8<#EHV5>+C?Y<B:@P,<,7X&gfYT/&dNQE(dR5)Mc/3]bA\X?UX,GgU&KT6
;2dY,\PQL1S=dJZF7d[QV[[0gA+?b@c-[#M:;HV]Q4B(R\fd6:LV0QK675U]SDKT
FdWWAX^&P]+.SdF[+K]^<X8&IVg;XIGUZ[]L6XX]b/7).>NB9dLT3DJFLfgFPc=6
?^1eIBG^22_2PZd;ZB/gQ3e)S,#?Z/KfS3/I2N@2TF;]5PHP6+T^J5e7DT;(W@cO
^&gCge&/3\0<e5D\cC0+^QM[LLPK.R\=5]>J5DRBAY=\YG87eB)LPbcNRBCM409[
VZ\BedNL(,c_+]B\fQH.UdJHO+WG]e:(<74KM/]OFO63;O=TCOS&B]53PB(LK)XB
:>BZ4fN\0E:g\PQ?;RV@>P52IGA;(5&I?O/71FW-OC>e:[1J/8-1X\QCa]K&#:g7
#Z;YV>#O[T_^9409^G#Q<@\VY>-XdO]4SX/[+?C1SQO2Jg+W@1+6fL<)CLIC5DaV
J-=Y\YcbF:Z9MaHNRBU;PP?6M94-JFbcWQaX,P5WB[N2EJc=-Vb);f1R5()#19V<
Z#YaGK[e36;b-a\.23XI=BJ@ddH7E)R#CW++X(2I1C>Y1bS>#YG;I<5_4,Q#8RLd
,cT8J>S[3DCRA,6,-H1>S;]4TR@-fGMC/cfB^VEaDMfVCSC8XP27W9N)5Y;:UQ/^
CC?IC,W9]JW-1[R,ZDNRW:5Za):ZXgAe<X(&;e-)U6.2CF_Y0TcL4#,T6&9^D]O0
?VJZ+/#+8[Jg7eVd4>2LHa)E.\U1_9P8X3\=K=]RZH,/]+ce;1a>NG3?/BEeeH5^
_93>YK[(3OA1)7[Vg?,IMaLA/[]g9)V_X[9?2bFg=\G9E9K7GbYg+:A@KB)+CMgP
/<_CB,R8(7(8Z=Q(2/A-A)9&[9M+JbR,FCdJ?]Oab]-;1H/f/0WbQG=UOD1_>]TK
DMYbb+[./@.?:d:=bYKF]TWK+=8S2554(T0D0AGNY>YcY^9HX@EM<c._:..8Z1^(
ZM@Z7@-627YYca(eT0<QA)g^M/f?3E+>EgBTT1ZcK6ANabFa0NA(U-]aDI+P:QT=
FNdg3)B5(XKbBgf[HHNa7//1QX6Sf/e75/cc47b;T81:T19AODR+Y:_0U.6[[Q@5
O5&(0G-fP@RO7bBLV+-8MeN1P^2HZ9S\KC6;A9^&7MXJ:/59E0FC+6P4Xa[/J7Pf
G&ECP+_IT4N:IVQeHd#KfdS-ANGRG2I5PRg4Taf#R#E]WTa[7Q=dPZ>2(CU[NAF7
H0-dS+2[QD._e,c;R>]L7cS=N>.]d=4@E<He7542=UYNN=T/2:_^Pe>Y]7ZdK^L/
+C7,X,]=LJ47]>[:-2@<.^_.a26O[E+BNM;D]B=--I/B65=-d82d/Xc3<SQ<:6LI
L0ReRGLN1\70cFSe/._O)T9TOgJcIgT(RJ9WN5U-/[Ne]f::H=AIYF+aJRTXD7OZ
WeD(Yc[^F<T3b=U][;A_ObE,7Df\-.ZaeV>>-B?4@U0Z/cRDGVd,BMKIB_UccY#O
J,gB+T>-1,S_]22S>]R?]J>Na\=9VS/^?3SKSBC:L?@\Q;)R2.a9\5V@D&#7.DJ:
_;K?QbL,ILXS9V/g#XD\+.d&\TQdEOMbTQB9P7cVS:SF6K^E@(SR6&2:\/3aV=F>
^.6e9J0H#AY[]HAaKa=eg3VNUF?3=YaJO]@7R3?&?E9U.<A7B2FLB#QPUJ;EVA9=
#8<XCO\/eN^K7^QIBXQe_=;KY\0-@OQ5N4>=J@+T?3^gI^[]@5/OSfSOb^VTI0;^
Re6M65fV1J?RT#1258Gb)?_bS6(E1[=f5_RMdcFJ^7^c9SOCVZ_PYC8P:UKaXd-4
DBZI6I3(7\5ggWOC]9ZOeW<Cc[I#6]62XS6B6d\+NcQ2KA@DMb9;2B-MIbC&XM;&
M0YWBSYZag^bJZ>R^NHL3b]O=CQMJd<F;=G3I00BBDE^Og@JIPbTeXS5E/X:QUbQ
aMfT-V/Tb_DE8.3DY5.<L4<-0;C^1.M0I/ZK#e,HA2;.J;NHS1<^X/CI[,X]ISCc
7_@JC]fW?^bd-MUEFdL&_))ODE\.NY4?DDE1RJ])ffZFXO=(=W,FFLIc8,UKROf;
@T)TR(ZB4?Z@WGSeVJL2C?dRWX0F1aA(&9>EdAK8gd2ILgXcF^JE6-(P#Fab7bX1
c&/\:2A(S\W=HBAF6>GdWF97XM3KW?JbK=D41Mf<A7>](A6)UU-_Z0V-9PJ+XUOd
25I.9Jd5).HZ(S[aE7]e42:\;C8Qf^H\5E)9?/WZG,(.JZ8,JE66VP6;BW))O4KO
HC.2.DVNXg7K.C2)J8V1@ObHO.G6[VP,HGgUN[=\AW/K/Aa8@&VS[H.c6]FPD&fK
c?C8SDJ2LW[0[)-=>HM398[;baVTc+A0f;S1N3&Of3Rg7NYV^e(?_b3/CK=D]-GY
;Y54g4#YCT0cFR?NQ:-B-1Q;7MR25)XOY3Q#1KVDSID+3^OH>L@4#@3A_.8,<][&
dLP&73EJT8d)?W#P:J6QZQUZ9]MGdbK/=2.\.^B5;=H+]gR593AH-efgWO@QTg#B
C.[PcX_OYcf<CY9UIMZROO\,R@XFf>92VWSI(U7IBa9_0B0J&NOXS\XAM+DGL+[a
UF@dFCd.,1R@HUgZGTHXLM5_E.&;1WR,[@2=.L[Pb)aG52AT:\MG2U<-+93W@NSV
2U<Cf_V\4^]=DY+>B86>F)[)+/[R&)g?_O]g#Y33>W:L><KbPB;DPgcC/AARBaXb
Y#I4^W-:^cFd0Xg8#JcW;/(OO/9-ZW/IB+A\[aQHc>&PffJ5L3]+,59KP<=7RIQR
2H(B#QFM+A?0G7d:_bT@I33UZfS?LS7NRf3AA[DO_Z@7WHG-;1+0OP/_ENMKU)+J
,AA_F.X>C5MI,G1@:&48NVe151#[<(,E3R:a@/bbDUS=W^>XEP=TF7[(-FL+&HM&
g;gTN2D68d?f_=a6DJ[da@.-6Z,D))9gbH3FdfL@.6e_=T67ZRYX(&DMV-Ie@D0S
&\6<HT4^,HJ2/CD^\c2cPE_I,+:BLb/JKI];.<dZTf.106PXGD\g,4T0aMB;3&NB
7G\SP50Be=MXH[)A-&\==46Q4351](6K08AbUF5VJD7.-gA)I>FH4ZI:QH&MP3gA
Ee,.ee\L<:YPdgQc5>9CM-#I^#PCa\VZ:@F-bfOa>CGEK1LZQfHP8c:\(J_U+V=^
455HVFd,6HNYU058,Nc,[FJCOFc#NFIX_3,;0IIJ_#A0@KU]HKB;JYfJD7g.PJ1N
7cD;JN>FH_+N@e-8H>)c;#6NQg9Z\[fIYMU.79DPUZUg_ITUZ;&)0;KN8Z#cVV+P
#&HPS?b[;TKQ_;8X.@F7dfM3]P[4L2-_\/^ZWcGYB-9K;_2[@KQT=O=B)MEQQ=A<
cPN#C)?SB4&C8M?KDYP&OP?.K::(T&IeZM(g,FH9;B]SEX])28=6AOR65.7b.UBF
(K4484B?<<c7.NW#?.3QTJVTd:8RU6Q)-66\_d3^c_UX4XYZB7CZ7&<S22+[deDO
_1=J3=bUEGO+4#XKJ]:]#aN]/SVG)Y]4QLf4F<Abee_2A\:JLd7IEWCBRA3OI#1K
JH<B)0@I/DH:7?UI/+AS36ACGeKeS6Y-@ZY/:I(6LP6W&HDDd9NFD5I@]>HDRbBF
5T>=326R(+:UJP?Kg>P-/--A28XG7fWfC5bbF^#MA+219Bc_6HL/O=2TQ;1Q,IfI
Mf)MdAE<-RQT8DQdbRfG+R&WXF]@QBY0Qa.&=X1=WA&S[,D:_6D_OU?<7-2CO_&&
7GWVOW)-,>KO=Hf#WcNI;dVL(MQHQ5H/)(40(1EAG2L#db#Z?e7-&7:G#I7)3:V0
VQ9@)OMdZ/DI9@<BIO8P(fVBR79<W+,\Kf:XEdITgZ;^EcE5Fg:0S5R.0f_cdRd<
b7[c(>HB@#D.G9=\4GFa/AK1/1</4E)Uf&Sf<GP@/+[Wg[/U->QBL?bG5@b[:GR\
aKd4Uc8#f1Q&(S:JLd?[0?A<]]/]8fH0.E-@&#M2dW^[EQBfM7JSK1,W8<BaSR1&
?S?G/MgPKYT450U>cK=e(,L?][.P9RD=P^UdC\-fe8<e)[#XT)?-_?F\5HFQG-@\
9=CbLgb(17O<P4N+]2_RMT427PgKQ+2[;PRA<FTb@Z7?I0P5f.XWT5TE+,?b<OM&
]bF643X((A[NW7feD4/ODJ^Z6?FGK(QKM(\H@#ggZDU#bAH4R[dWLQN-/[3[?aQ(
#KDf[Ee_DQ9XY1FXcJ?N\ZAJ1G1S2-:RV:LUcY[,IFXZd2W0<(,ZUFFC;GL]7f6J
^e80(-c,U<:Y26Jg=HQ^>RQd.&LQSdCDXBfCXK7D8N00;GJDG84<(U0XDQZd=:?.
(-PK2J8H0A;W)_SI^.[&7L@d5RGa:NI7ZC89+gIPW@(<FZ>.?#]M;+3Od&&<^8Zc
5ROFYAFWK(bO72@5]4AM>N>YU88&([gg;^P@XXg6WeX=[=,GN?V]G(=>e8.IbSb;
aXD2A5X>_HQE9G<Y0):/eMWITC\+H--SILXI[I08G:SdH,6d&1JH5HQ^^2bb<=F(
7?7@O.)YZ#[XdLMXf+R,>3L#EYCWI)<:8J-gMPVc^6;P\Z=3N&8a._OY5XID--&Y
R:V9+5BJB8>=9d0A882\<<RNP#K/#WXD:./gW)Fe^g4&0Z\8V6gK<],6\,-(Z@CU
+-7<>8UJNTONgOMFOXG<OLQZU3WIUJ,<9E?#)CVQZMdab>TRaFEJUF>1>JOQ&Ibc
>.<2eGV?(eO?1\O52dR+1@)@e:XWB5UcGN5.[<:4]N5QGD.QVW[2C=0-30:\CI8?
E#P2HbJN=N[E1^VPRFJ?JeM_MdR;/>M;XT.Z:f4-,.Z3C^W5&a<c7N:#FbJHMVVR
YRBP/H&UN56X\3A(,_dJ@5ZA9\c#M+C)-LT+I9832//?edZ4/Y=-LEA<88)TZ2(B
A37MX(PQ(,Ya[7/g92:D^GVI6#a7.O^+2HHJ)O.5]G;a[ea94\CG[?7cWOOTAAVP
d6^V1;ad^YGgc3A@NWY^23.MPeD86]7[aP29]6:P\^]M]>_g.\Mc:JQV]<NEfPFP
eY=b:a_?O2IZ6F5?:\SZF5OSD&FH<5MG:Kd+C\VVg0IfQT#c+0+?>=(J]2]AaOB,
Z&Q&Rg8IJ@Z8DUJN)A_<ZZK[b4W[9>eLYLT#CRJI=c4:^X.,U,U[E+P15Aa[GB36
2f1b90g45Q@?WKH@4ddYQ:QE<^DfZD\XGg8;X38VAfdT#7RS8]LAb5?2YA;+-2(O
DC#CL[UB?J^O=4MPfV@2(#RcWREG9QBSJFXf:<?^DGJ0_=#-]:1Dc0cWOMBMO;OY
A)F>+1S1XWa:bXBRc=d)g^8@95.d[4&\UY@Rcb58Z^<(+C+NG9>ACEAG<67NFJfH
DE_aJgN:,QD>:\@\N[1(RVR?>=c)/(-O:f][PMZF/B(Ef^]HCcGJ]eZc@J=?+CMS
>2;\57((Xa9SIfaW=.Z]#WfTV9RU2DJ>N2g>SM8=WT;?06G\cXg+MfLU.?-Ga71g
9^HZcO/4B4=O3=Wg)d026Y#bFX3I?5d2_C1Q^PdD\A8A<X<ME@NG97:Z0F1J_)KK
_<bc#3LAO\8QReJg,TOT>b1FcO[CD\9R_2Ib-f.2\-8;>:<_ZWRG+cT.]XSFa/LH
1;]9K^D;IU<B\BWab0bWQg:dN<adM/TI6P9IW?92?CaL(9E(DIH>)6;R,LR8:+US
KJ/VF^-J?TT==ZB]CE_D1gX2F2QVfg<F6WF88(M1)S7I3@=6_;gcdEOSARUa/9@9
^/M.\,_L:Q0#&]>8APXW1TLO-XgfHEd:B&1,LCTZVgF90dT0>JVFd)A(RCURGN_6
RNcD0YY1gId.X/R(^CG\I<W?MX1G/1)a]P\c4-I@4a4Y<6#f3BGDd0F>fP;@/Ofd
1ZCF/c<<P/A->cJQN/F9TO2N3MK@]I?G@_J+DV@>#=AC-?P+[a84G1.)1X__KPN4
:]./4,PRa:aHS^-Z/GDRU5O,HAA7Kg^d^MI9W35@XA/.8^7U?6>E\e>QfP:AGTE+
.\4,KNb:\;b=2N718W,.b@NU3N75,6>E:dVEJa>&_H2PFf214/Hc+6V-M7BI;)>I
8f<\gO@\[gfa6BQ-OT6/W#Q;SC/eeB6[/I[0eNM2;&d01\::dK(4F53^=U-V>YHL
R9/_II9E=A+D;5U,UgBQX]NC&M0-Sc?\&5(4\KBA_P@bMdTc:.BXe/6cB)Y\5f3,
aD;4P2e^FT^55PCMLO1>F]W:]g<@</V>UTEMUeWf[GJZFb>)+Ngg(MbZL[^+L9]#
8a+V0b@++W#X</99SMGEJB1<#Y[A.fV2CDNc8JWNLf-d1a.c7+47QBK.ZR2+gB\#
>NV&ZbNR?-1d,U[+930NM@ZPeX\@>;PEZAK1NAP#V\>32.^<-K253C3_.L\YGg,/
^WXTc(]E628)E2_<Q?&O/f/+B=(1/BNfG,VSMIE#)VK>=AR2<0Y<<-@:ELUdPdH5
)bEMQ=Y15A@M&;<We;F:NeAVPG>].@EUfAKD6EE#6ZeE:MWFC.&N:^I:\TcH2]KD
L_?_UR/;TNeaGba@A<DUL,P:Z:FL2,VBB6\:dX2@<P=78QUc1I>XdRf]H9=O+6&;
@FZ@RJ5YB-QDXD#QcI<^SaK_?_R?AN31V3gbaJ\D-1BNYS?6e#Y5S1SR4ULa\Pcc
+QPX\][89(b+Je[CGX\;Fg&>FNR,UILWe5<CCH0bUdTG3O\a=Kdf]<X^_R.D:7>S
][5^7J?-^R@&V+?0#D#Q(&Ce[eS:R5]f#U2D216G/CNP3SW==#TW)7/(\B_5#QX4
X(@>--?PW6ae<7634ISeLdMSTSG<c&?(fP6\0O1V=RIOCdSUe#e:\R_:C6).ZKRP
NBZ2g=>29\Xg-I3UeIU8LD5/E6N7?32GT.><RPTMfdNAgOF6:WUW_KZ8=7R]gGc8
M<SMY3_M.N6R](9B]gDaIRC_G?I2KWE[MPe70#X35WAQ5M[/6F^_9IM0a].=f_IX
Je+8OQ<CDCL1_Z@HfS),AU9.Q00aA);_Ke@3.8c(0HNG&Z0CP0;<\J\J&ZaY(B7;
f;O;&a1#dEg02JgSaZSP_M#HH8;64,&#YD_e^)D@dC_0O--J?b?C>9Ka;C<dU@eS
2&O06>+@I[A^QDE<HEF^6_JOCGc.C]AJL+QT563LD=dPRWM/](78Z_QP14a^Sf4<
Bg8DO6&0T:@;Ag9ba^-0CG(:)X66>FD:TF3Mafd2#adWVUCZ4J9[3UV:^D&X@cG=
3RS;fg/_>Q-K;>aM,HN-e[^K88Z-CNQH[(:A6^PH#04.\3PC:J/U,2W9eEG(&14/
:9F]C#BP>34J3=Tda2)_bS;96RWbY)_;UN98:Jd,)eWZ7@[)YKJc,>2BF][480aW
GgfL(dCF5aWQf^>T_.3JLa4+[-TS95&W8e@GNW4AacG^:_++M,?Y+/RXbZU&>?<7
d\F1;]a-L_MU.#.3egU;KT4W/)+dc[Q_[;K>E@\aQ(BUM?f&&bP.&5/AI0;(e-A[
W:@;fOV>2KQ6]b_PM[JG/UB-9NG9V9fOKFY7KJe4[S2eH_G74I7.[D8H@0UVZ,DI
;fK#JcZ^:9HB_;+d3aU\=JKUM:ba\I&g/DB_]@@U;PV:(gI+^]HAc64+9,U]7Hfe
3S,B+C;.^,dY0CU^I87U/_e7>P.CfC\XWdcQ_@g?U[gPFN&-\4T?1,0d:3=^CIT5
FEEUR:\,;G;=+&g&Qe2F([d6,f_>@8NXKDR:^[48:JdIX5=+=I6P.?BfSZ)ORPDg
#.bC=Gc?(bbX\2+R0gK[VLZMC(X2CHZ=,#&4,&(D49F086/.6YF4F,R-BT;9<Ad>
afBAZcC&d<7.1C=?KAM(J8=5-IDU)#P>?2)YdB^)d).gS4Y4OgU]b8HDNLHf)QQ2
OT.,6<:N/32I;CT\?C1\aZ&Z.BT.G5[eXIL@K9Y2V_X.d-V0)9(TEK39;cKa)6:N
(_]:J)\+Fe5)R7BQE\SW:S40^\:4HN5,E;39:ULL]H@d2>U&bBee78Q+:X-&A\VE
]=/dW.T>]fe6Ye\B3D(7MeeWL_-gELgE?O@X&c4Y[A91(H\GB2IdQSR<C_3.JD>[
<,^03/PO/3]YN-:I^fY[?fcL[4?<BTY#9#+JgTY\\RNdbX\E?]cS3TNF8P;SZ],E
gWY&0R\(8_3[?AO^:@gII04^PT[+3JdPgFVS-1CBLRRIMW\C+31:+]f_5aAI4^a6
Kg>C=b@X@EE)?>3<L0A8FNgT:HFX.+I=R?4LV3J7Ud_>I=W7=B3/G=8U^J;+d5a7
c?FLeX;>a(?ZD9YQP>&1^^>>.aN<YOY7&FR93#+NZT)GQ^&Ygg-HOK[4dDKV];ef
=Q2P6DFcUFP50^6O\VfI?^?0-_3B<]FK[XOP?ND9Y@08\I(#Re+WRB+I=eL,?a#J
?^[-d_Y2#3+7(EWY83:4.A]OR9&R?@F0OO=aKKE)<2B/1W+/MGUAYPTXEE5X1Dc,
8GIL;bM\\=;=MYQ4-3C/#2XLJC\60N:[Og\aKDT[LINSL2,W>]>0P>EBBCV&16Q?
7.\+a#AQOg^>2Y+7,bgTJOFB@W1[-e_E[_\DAT^C8/J6]D,<Gc-OHAK=;S)abbMZ
aa-5Gc]D24R1b+H5,L]b61=fX.22[CSb1,G@5@F<V-Ra^-+][/([bF1NSLB4]a/G
M]6@,XYEDfA?+1ML)R/+83V.KMUKDQ\dAP>=fadXFeb\?OCKM>/fU>@6g7[(_,(L
.d+K&eW91P5-\C4Xb?W7N3MZF3#BOJe^;aV1;(XN(X>N7XX]1/_eNXM/_;H@>Q)_
O^UAQ?<A\bd2,:.18)f@OV_\g<O2a>0+LI3GSceN\CS+CH/G74D&1U4?(M8T1=,0
BO6FL4W>?>G<24;D,/NW056P9&^^/^5?HG:QHL[A[aX?1_&fRP7F2W^0B6>A06;J
IW;8([?C3RYG)N+(,NOI=D;0.W2L:@3717(?P+D1]J)3[O9eFeZH,F<NRNf6c;^:
T70_/LGd70RCFf=AM#CVMP02L/d<&OLdHgbJdQB=^McM\I97Ebb<)f)<=ba6eQ96
:ca-0,;.eJQF#:aD^I_@(5+dT15=@94(G3HKYXIA52AEfET,d#:HU[];T\5R#bL;
&+01)5?=4cge>1;dc6;cXGZRTX6-9Y8T:8Fc?Y\D3DJ-La6\e@<?R1]+c.OHJ\4K
3ML?^WgDb0aL(_<L+dNM&g(PR^JLWf5Y49dKC[)>g:)9MNBf/fC6S\+OJB7.>SVK
H+YQ@-1,:HECCd+S.R#g=F4M:H(SUe2\9/0PF0=.]AHdZ8]2WXD?9bMR&ddYG>_3
G5C03>Jg3-NO[c;ZKcK)@1#/#;27aY8e)Z9d9cR>HOI?FWE[S/AWgOJ@[6>d-f-c
K(XUH]Q3V5Q3+VOE&>JD5_-I#[MB\g_JY0_WGba)Y0&@I?;=MD),#NY0c6KQ(]3\
>dFALMLEf/AP0)aQC\[/(faDcPT3>fUc8)SH;CaG?DJbBERU3V^\(8Hf_RX8cF1F
8,-HJ2U02aF5=M_43>MP+3.M(UceFLD9Ef6bLTe2;->-gYASEB2?C[N[O(a^ZL43
J\6MIK\7M+>KN7dgeA^T?g/[IGPPNaOdCa>CBYW9<X33g/1L0>,2++U#>3fffJ4@
L_]QKc:3)(TLW@)Q8c]]83)+>g-UUU1NU</8E36;6]BWO2&,OB&H04/>FA,]Y[.F
cR.CF(B)[C4M:]9/cXG@;I7_7&EO?&8UdAH=E&^LZ>?AJMV5GKY<8E>;c0e(TeJR
_;=K2ID7JCaC#:,bUTJTXO7de8)]9B?WIP?&&OC.I,PGNZ(0=]D7[E8(6E1@Y49W
;bdRe@,&f+D3)/U7NW[H>#C=QD97K,_W[PP,bGVBcV9>.^OVLP8fHJI3S,=>P7;B
+19>?_.:S,.=XdZbJ-+=D)@YCB^&bf1UQWK[)JLIJMcE0J9#d(9N0S24@G41V8f+
Zb>g1BHNY+:-,??2[:JaHL8d/1(V5DA9a#?<=cX=65=-J4?S0FP9_+D+\-1]9&e,
QRKSfT9X@0:IaO&0F6&5_MEDSP+/V<562R79?^WGUOK)?IBZJY/(24S^/g^eRWFW
QBY[B>W29VMBbd.QZ_&a4VBV[7:UJNVL5X>7_81Q-(^G46_G6DA>=)QJ3aN##8e-
)a0PN?Y94_HW=?4->97G\)D6c+RR:Q9XXMIIH+fY<OP7JG_&:,O.CDK[10YM8MbZ
>?Xa=_53<,PV^HF;B<I\<Y23(c6N+eTS]STRP<6>QgT&V<9[>VO-XK-JF9>).aEb
LcPLG.M7GF9<U;J9Z&:+^?,H-E;[<>?6e=+a:gac:cfQ9<YPO9Q(c,4Y;_;EAfRT
&==_.3Q<=CU<P3393F(]7HUKb7><FLM8eLA-cU5&WEX>,P18PGA>[=&^V7+,GBXP
]EXDcOPY5IG5WJL.]V6Q&R=R58@JC[)gG;S)(N+e7PJDU]S,ATN@CGV1FT2FD7cF
c)BIe[,0Q0;AF#\<#99YOc?0)?\1&^)Yff76[bZ]e.W<#76JXSC_/H;,ZP4faNFX
gZ&^?M1d##G5>CA,^2R:9\6HeH15CaDM+NY-DO4O)#.H6Y+aATE9SeXGEcf>PXG<
HF2(^_YTME;[QXR?IY:TU4L12&?c3NdRWMNGf-+11WN+.[bc.^fV1MB+:5Ng(cJO
P(7CV1/U9;/XX76O=&][8f@BEJZ+7X.V_a\J]G+2KOP,+<O6H\SdW@Pe+?7=(\S#
&A(2A)<?dWD\(PaV-GY/EE;194f5?cOPK<&@_)XXB[YPPdD?;,#Sa7:[#6Z:@NI,
_e;KL/dMQY.;+cgCNGDdULW4D0B7)#F?I^<d10Q2QD(IRIW=(1d\[eME.HZ.<LG7
G1._ZL:HH2HAeWID35R>E.-.VWbGFNBaO<H4XYcB?6/?#bZ=PEUD=T[ME\W^/C#:
=>&DH+42275<+TaJ(Z+O5-B]X:LXTKT=0Pg,PV)LY[b6CS@NS>SF)QU6Na?[_#<P
OF:&Z)N\6c0/6JeLH;OMFA71-_(Y_].1N#e8cTJ]7>V,70^Y7:W-JfQXO.7>A/cX
:Sa6.@EM[,+aH9_gbI:OK=G;)d=Ce/9#@V6Ng_W@f7Je7055-?ILbg(YNMg_Q<3O
>3d.ZA-?F(YOX27\W^><LUc9[>VM;H^G:A?&7,>F?c#TTQd>3(317,KCC5CO8g@E
M>B\B52M,(SWAP[DTa]/ZTSQ8@>+9L\(9138QZ+W7)aNdcZY=7dF]29dOTZgQFc-
A\8dg=<Y[>T<,.bB_)Y_CW=GKR=87?Q6e/#N-P).8EF2/V<M.ebHRN)H>8JgO44(
X.+<fE^4&9<,#J100I=:)Z(DKK1OKHg3(7:2B6ZSZUg4dfc\Na-4Md:0KHHX8JJ3
@@Xc^aY,:DSNV(\M3/IN6e#[\=Z6KD0TI:-=[RL2ZPeP:#3=-<J12^.BH]g3Q+61
CE?J]:dWME0g<8094R2N)HOE,72TQ]M.TgTSUPPeZZ&S2CF8;CHc7LPgc21L9ba9
IUI;LJ;WF6/F#W3A5CH<X;a;(XX73+^\YG4Y)-=FP(21aI<GD9604b/7NM]I_Ye)
BHAJIdPH@NPWf&d.3d#P0+?^Q5A?-aAA?)-=Y3A&+6E+cSe.IWSE]ZcYL^9#b6P>
cG53KQ:;aEM0b;^b1MBSOOT;L)UeMHIVT6+C^/HTS<4R>40T=6Wbd&B-6FTf6WIM
<-<N\8?_2ZV+DcZ>7_Da-^A>Q9]F>UfdD9]g/V(@I_UBIU]LO<1.ST^NZ0H/U5&[
dFF->;U[8\+fD\CK3NXH<G\(Ca[YO@N(U0:\;8Y>Z(Z0)4(cT6Q->886HH3#/JgG
9&:f.CQJ1Z]4]:NL=.KP/6=WX-Y?)X4[gMQ)@P9AX,Q0>8L9PX#GJ,L\JG@)9F7,
F/ABffBg_Z?-FaNZ#?/HC8J=34]T[SZ91+M+5@M8F7I&7(1;5]RGe5_DGLP;R@Af
f,)RW8dc)Z=EGMFF\;II?8^X77=#KV,W?0PA+L/gbRE?>8LS;)4Z>#L:]P76=TVT
0QO9[/IZ36SNOELD<UT52)\NQNLXPXVA9+-dD,(L0></D?L4HCeg21L)@,53f+]<
@&/-d-DI:([)]HU,@<dFMWF557DUF3OAc)T_X(baRY/2C-+_<c_NBS^3Jaa=T\])
J]WBAYQ:RFeM1Q.IXfSH3aV&aC16Y70)U)a3(IQ,Rb7=IbLCW]^[G\U-]?K@)egI
b1^b-#QQZ^NLcLO?\Ze7=CdVAWefR]B?>(G-@JNR0RWN.@Q3E#dNF#bG&?L^LcC-
?PD;Q/Mc]C_@B>O([6/b^FL\I]a==O<eD2G9LYVUU:AODf2ZVLf@:PFg>W0\ZAaZ
.20dCE#SK#29c1@(6OJDK3WTV,9>H7#KNb^e;_Yg-)BPPJa8MI2BB80N6O8GO_IO
T0cUKaPNgBS;\)?X0V0\L8;)a;R37@;MT(MW2@b;50@+VPT&0:DSCR\d&CeS@@DA
M0WH^S/LFMNEbcg@edT(O^#bP72D\aTa?L-fE1Q/:DY\P>.d^aF;gICT6KbTDA0-
9^I(XP1?)O&;6:,6Hd3+7]7/RE5@M&T&E_PN#]e(N/]@SV]^E)ffFT&gF/aa:MaC
RIHGafc<=:&LC\/=H+BW)gW+_HJR_>F:80MU]bd5U;9Sc4;<R#E2]MVAO@CJO.PR
LJE8d>:BQY:;7V:/89UXCF;Z;9O2ZeLD4L+F65U@@N=PY^FKb-=UHTV7e-63(d,1
@+XUaXCQ\R]]T,QGRBNI]/-G\dc]=O@RWDe>=/NOg@Q+K(C=DY3\G2+:_.=gIKR-
2(eRQPA(&)adHf<b=54D#L7;<;@1UKR[[ZeE#.A#A+OGe54MT(?>>21T>c_W/U]g
Z(_?]R4Y^U6G0BYPAGHdMTac^KZV97W#CMKCK_@5LV=V>-2c6aB/6<KYe^W[ZbH<
A19agI/M==ZC#:<3THXX/Lg_+I=OL8+4+0GRG2L]T45-JHBfQc<Jc8f@g>F00;?e
6X@O7HKXBc)fVPM6gMcfITRgZLAVHeg_J_?MQ#E.LDBB)+3Z#;]8O6)94-WPaA-U
.,>1-68._D8)3dZ>1fa5]eg].e+DKU-NaZO[]fJ3e,\\5g1LKg)]_U6_Q?IRQ]ed
,QE.>YD+8W_?=H@ePWU#PSRJA,@?=-a;Q5RK&70[LP@-=UPZP;HP,_SJb4;H/TN<
YV0)0X#;KDdX;UF42J.OZLB,RD0+@Y+D2DTNV;eGW9A,@;dY92C/D(IKDbN:/DF;
gG[XE8MgQ2Sd<>TfY+M<2@eES0[6dKK-;\7YW(<e)a+(6-8TTRJ<G?+.g[;JZ:MJ
E7)390_+9F#c3N^E-eW(V]7cJ-MEQSQg5J8g4>@B&5DPgEDM?5Y_Nc_FE]3,SJ(R
U1IIIUW8Ha0a?JSK=>4V.37cDM)9^(&99ceZJ06]_JJaHS(,[24<4GEg_Bc3acX-
BTRA(;5E[d?,YO(AJe-4_E8>,,<JP+:JM2S<Y:GLeGB;L0</X7MZ90VNQO.eG(K(
+U:\>B]FOA<NMJ36=L0#YdT222N2331.4de)f-@eC,7F#YRI559b2OJ8UPR5gH56
57P<FcX_-HB02cAU[W]/J&1Wc[7T:I0+f<G,e\CKKK&X/Q71/Ne&D;cIX,2g,44K
2<+OPY,b1TRI-VcAPeIL>1f>N7Z.JAH^7b=#<MR\A6dP4:+W3bK(&_9cJGT(J4)C
:9[RJfAc3,28QRfC4@]?([RTI9[:d/Tf0JW8AHFBP:,23<>56;2FebJ(2:SRc7QN
L@]c>+FX_P.YG.]J8UP10[_MC(R31ZFDNEaLV6@=G]K:\S71JX9)D.K-bI^X0)6O
g5G+PX5@\#X#<S9g7UG<9AK5=gE@=I=7+()1d:<M7M44a3_EB-,eE2]B/^KH@@U8
cFeDDC(G<JQ=L@f]3FW1P;LbMEeG].##,^VXWd[C5:eV]HfJcMGL4MXPF.JX@1-A
5KY#A(3)W32?8Z=g\QRUCfaa).399g0\SX#TVBA2FBK-09FdVM3.N<+#0JKL<C9;
+Wa6R5O1DY6)<Z)<WbV6;;4dW^R2HN]]3Vb@eEX(/GdO)F2=gd5\G4TW=W^Q0^Z]
X,a^/H\2I15eUf8-[N8^>TU-TSHXdQR;=e5/.,8=Q[F,Ead]7(E,Y4<[6ZG;8_RL
:KNDdEP9)bSXBaR?<g<I:DeXJ]DUK(8\3aNSS.B-S-5ONa-6EK\g(=CNE5FLAHV(
4)fKG15=24(B5I\AHCRI11PaO;^182?T#4bFW+XfV8PU(J=[Xf>dLI0gJF:?Wb1g
PMQfRQa4FS#C9F:Q&5:BGHTcf-Ud/EcA?QBc54geP9JD?2;3N<:E7_]<][83RBc)
dC-[>L>,>J0d=SO]_0:UJ(c(+G5-W7SdJ/P4#]Qc.XKIFGS06XR5=?#<@a/7#OC5
P)18DMWg,P\4=IX1d1FP8(H9IcHg3T/Gc/JBOb-J[JLbgR>d48BC/Z3Z+d3V=IQX
U9<S78JD.?27S?#PH5DP(S1#ZXc.(@ACKdL+IM3@3252VC+54YOQDFCS+I2/@YCE
&W:d2C(5.=Y=bK7+.N5],A5SdJ8.UK>?Y=ZSXZ\_52:GcS3^QE1E;^GAf&=cM,WX
6-;Ic=cNC,Y]W:99a_=g^F=S+g&A?WGAdJ[O7?2E5]Yd#=02@gKfe9MV.bf<.DW&
gda<L4_\)#]C,4JA9/HJ,?,G>.V)WGKAKANMX>S?,KJX8^JO8(1#0#-.I(SE-9T/
GZ)2g;:J]6a4<bY(KfGca3aZA_cN=4/0U>0M:F.C7GL2Sg597f&Be>JY9YX^]E8,
4dU8,16JCeEN#5Se\fe),d(QA;BQ4G_^(++;+2b)H7N8L(Ie>RTIU2S8Y-JEU,(:
e4LRAIcAT:MfeGWX&[&.M(gXJIZVHC^]cdEX:83.JURNT;AN1Qg/6>=NM4e9;c5Y
VSH;-2Gb)JZdM./A4Z214CTf.AJe(K4X3YZI_dGBZ3Q,2R5M:A?EE1#D#L0M@VG[
=TW#7a.H6KS:(/S\;C+RDZ4eWIP@PUK[gg2VMK4HLCBKR@0[d,B6KJDGS>>R]>-&
2XC+Y@OV6]Z2Ia]T>Ufafdg[9Laa3TZ_):0.)Z6F#+B/(+A:2&CCXDTFJ=[dQbA4
V]WPKVR]5;Rba;EQZ?HPM2(\\Ff0(8T]224R1J_H30Z\A)bP)L0/g=D,R]VXH1_b
+?V^60AJa97-Y03(ED&3FNE/?^(K1G(X]#eRGN2ME3TY;R@Z9^R#[^3CG;--ffgG
]<)RMX@SA=E6WggM67GZaBCUQ^+W#QJ4VNMbOb>Ea&GAZ=&;NEgI3>Z.])\48;-I
;If58bXT6SW?9DX=MP9JS?[8L(=,:e<&<&/b4)&LML^@^&&]1PGP;1NW=9PY\Zg7
,&]?MY;\RN_BeTQ0fN_a=+G;YJI5TR;N4GCEXQ=7]fG2IFPX_X1W9)E5XB)e+feP
;7J>?ZURYT4-RN(6I=<=gZ1=85L0)W^C&N[#EQ2_e=-^9>[bPYIe3;_#=Ya\aE3E
&_a<INS#Z306@--LWSRC-X8,>&WGN:,RYIW,Q.dcE3ET0YB\E:cU8Y@]O3#(2=_G
KO6_=1+],:;Y-ZZgF[8EZ[LaO>JII5[ECUG.BVT^FJ#,gR/K#ae4=.KUI]])WGA3
Z>W)WA;&WWgHY6/5.G4AUR4a+<3V0ePD60eSb+&\,5_I)401]B@ENd1bUF8IK]5]
3b<36R9;D<Y(V9c+J15^8Y<ME;GHBV&_-MPR93bEF0d2fWSH?FbQSSCT7&,Pg6ZQ
1Z(MQ5P6IcOTDW>Bc:>.NXb=:B8FZYFO>])P?Y)XSf=cSXSBX5A^?W0P]RD/_NbB
#@-Q<,eH>#-P0;I?32>;]X1N/HM9F5Q#[C671X<SLd)U+fL:WNU_?ecD(=I_<f8?
18\WE@d5eR9FBQBGff3;P6#JI:^[N2fD4PV^O_Y40CTVPFSddWY5e\CERH5\Z>Ub
QcI-_@Y:DMOZXG8a-\9c;-4V9KJ8=9a8,A3OE;dO+B4eb>)9e0D-)3)bQ=cYD99V
=ET)^XN-KCL5:,N]I.3L82[ABGS8>6/JR1Q+,4A,(.&2?S\d6Ngd3^)(9_<S\7;T
^;U35AVOV)K+BY+T(\bW_#7)PMY=3R#J\+WKe9XK<KAHO-A2A/_#VYJ&G)M+UKVD
P:c,]7R+0J<>]?<(-(_Id#,/B]ZfM3RbM\FBK9WX5(3^0fO]))3NFZSFAb_DKDYB
J_ZcTFH4GS+6G-W&H#dG^0+8e(IR?\bVN([8(QNS<DP4M;UB(C_1];CBEd&7>D#V
@J-#>8C7Y5>;H<<X4KZI.PQd]XXe75^XW2XH>B<NLPHBW5ZIaEEWaU(2,<QD#P\P
:<2_FL24WDSZAKa3132&XK:\-M2U-K[Y+d/EHg9/dcD&Pb<.4GC8=Z-A^PF_O?LO
M?&Vfd3Bf<X85;&20NU/TagNNWAN>&g4b8?3?@&MVB;B2g_[/EVg&@6:O6<X)dLO
4c.2G=Q=Y]YMNB:gFJ&ZW<7^_YL4<XcD_7=bNcK_GI;K=W]-^Y+VOJTI21JWN@@>
AV1MP[ZACQ1X.3d4/aH#_)=QNZ(Y,23DJc>DE920/K17fF,F5=fRROCG:7#@-4d&
@Z51<14B#76;I#_Y9H57E@\8NdGO5L;faO+(^Y:Yf9NQH4?eG-,\U<4H2,Ggf149
5Yg_TO?1P6H+f-VEAZ4f\R5S_5A7J4C?5Hc[HM7[(P1TeH-L^JR>S,ZD)^;ad4NK
BU+H(79\IU@aSb&cMZ/P0W441=3Y]PST)8cgM&1gYC9GLBXFDZcV(OLT]6CYY\.C
HT1Y6U6[g@KQ68[N8;H12B186Sb2BCO7d7.^^e:DICJZ[@4LO;PGd2LNZ\ZK7=E2
)gdF+IRd)X0/WdDZ6#^>8c=\cW@C^;[]g;OI(0:1ZJS+ZZB=W<^7Q+aKa2f52Q@V
-71P3]5RL#)7a^-9L^L?#^]\-FUPHW4R^ZX0O))#M232RQCY>f:eO5\:N<=0J<Hb
]EA(=&[UB@9d/gXK=4:N))-702dXID^29@DV:3Mc,EUHKWQJB?J3=>H)3)DQ0@d]
W36V-ac1]NB+Cb<BeXN^UE>1c8)F:O)7)POKZgB39UP+4C00_Q29?,1QU@(M+]7O
MJ/PW3+J6:#gF>Vf+.->WRUJ2#0=7#/ZCEN;VVFDg2=G5Z:\aQ_c,cg>?0f^RX[#
P=4:)<_&47#VSad@Zc2?9^9>-84K3&H>Fg4gc.]&](PO0B(eSHUT@^NeC[H1C]B<
G#RTR9?G?,Z-0XEfg].,Uc5Z1AJDJ@3N_WW4gVP_H4I#?Z:_a.gecN^?A^c=1Wd&
bK66@MES>dN0Y:#;dJ.83(E5(RLPMU(4=@B]dA)1W7&TMce@DXW+I22ZTNf6aPNf
CVD@1]@S(J9R8C\I.aSV0E1PP4[1/T]Z<AEM;02SOLOJ4BG-WJZ_dbVDO7_DbK:/
2F+)IUe3E;NCMWHdQ(]Ubb>D;B:=Ha/QY[O).-fT3?LG?+=SMHe-TdZ^WVV6W/#7
_cNH?\X#Ua_(+Y3IY6F-D<QObLRIg+<+E&HT29;ZQUNBEa#V^c9K7Mf04P;S,KTL
c[\,C8C;<bS;?KAJ5]@c/,IeES^X,;D2::<67X=a.H>)0C[,MQ\MX@/UZT6U]&R7
;[5a>gAX).RMfF)LW27TIT^TL14bC)90]G^:TKaYc4M>B48Ie4Y3FQeMP-6gaAaS
.OMMA.)-K&Q,NTJgVC6T\#H6=.:_Y1[?UVc;;8-8-d42e.G05>4QO.P?0#\Ic423
QVW119J.#[(T/-)KG2@V<>#XVRaLgN>M<PN/B@Z_+Z;c+ECgAPc7WWgHe@/;D3-2
2BR(/3=PT\eOI^F/+bB>V)@]]gLRW#1GeZ=d+C]<2JRTO6fG:#5T.G@\QJ^C>c2=
aBQJ4)Q,NBU@,K[G,6B^2;495(:;3-<P6_4]L4[[g(U-4:X)0E]-eIHNGcMLU+8]
J=-?WPJ+b52M,]AW__XV&fT3UM[CSB/0;XCLCfc-&8N6?VNKSQN^H[5X9?f(-+VQ
6.YL=V6GP.CVVdHD=+==<T2MTa>eD35.ONgV6gP+I/#RZI9^ce>;gX@XB.2?PD(@
8YW/ea>=eW=)Z1T^0+ZXP.V.E/bB-YeYEB)4[/IYE<=^U+F4]@I\93HWX<WLL:T#
[:9^8+K:bc](-9YYX;bVH76:>J?.V3OW@=U]H=f=6AHd7?A(gW;7cMNR4aMKd>g,
\M]/Ef9OA-&JTf<XS#2@P&Ug,C@?IFaX2C7)A)N#>Af8QOKM-=VPg.C1MVG,^7La
L<:T\BI85PWHX4fL0@.[_K><8c<83&D&DQIE+PJbf<]CY+=S+#O0/VXD&5F@QeYO
BNMNE9U:b;YN+=NV&)0YbL)_7J.A)E;N,NP,KN/dL,C0X3?93E90=\e:1]O<A;^c
/D#>@RAL\JV<;L&/4RA+YW<X_#IP^8=4aeK@#MS2HHD1MIP&XKU9B);\<>NE?2Ne
e;7b\PL1TBS9-^:HPO\6B===?X1AW.O6?+-eTS213MK,9fa;g:A+fLEY/gAdADB^
GI:7DD85Ng0#Z7#KPRMO4U9ZMR_57<7AQ(eH(HdHQ4(Q=>KDALgQ=7<4Tca@ON/@
B08)>c?S-S;85\AVU&.,ePb5XOK7IQ:ZIfdVe:9V74SeM8;(#/Q;;b5A+8^eM@:f
QVLZ858\YW&<OK,,5YE&Pd8@&V&+P>cRL_/4OH_##N&E^XUg3_.JYO+K??f6SdT9
8J[fII1-L<dgY[+;TZS0?)81;O,7XKb=c)9;6/dPN3b=3,V,e30d<F\(JZXPB&>U
I,e-b5W8H7L,:=<J1(ZG&II0O[/6PK?:?(eRLXege9.::dS+0>8P2Ic+&6[)L^^G
)IL1F3VgUKg:LM\\FL+#MeESXPJ\4RP]6N>e8>&+,A\NgWBNCN[E,5[e8_)B;XBC
C0IKb7aK>1DK@6=N1f_X9+]@I4W+ZT9]M4_c#C8FbX+=2\H__dDLQF&23.GB\=,:
J94P[C/.H\&,\DFRdfVQ=.\#I7QHQ^UM=A4gdD9MMFA<PGRGedd+UP>])A78-;[.
DRRZS1Y0ILbTW0W+[E8K2>=7cbG]HN+fXKTe6<bORVP=U\&4]YUL</-7[agE/F@Z
4O/W=@+LA1&]M?1E.3PEE0KFXccWfG5.Z-fFMeeC@IM3RUOcHD;_dO>BdNFM\f=F
>c?B6.>L22/Z^B750LS.,S#OJKZ/^?V?=eNQP_3V11X:IdRJbV+=.V\<AE@7GP^(
?O/1Z,6K6SJ@<ON&C=9d>SIQ,=f]JQFP+N@</C:=)<H9@0USM+,>LbObK<0NWg)B
O)>E9)b^,_b.@edV0T@J@R71d=[?@<cC_gbC7CK:ef^3&6/L]e?<UTg1P2K=NE8:
#S5f<#[410>WfZ1\)Q26++_M9e\FBccKeRYQLY4f>)3=YPHKLR.=38705?Z8^g.^
W(CPRP?PUKB2+U2)gFU-a<d#CM6ff832,67-a3KVRJS4C(eX9(TbOfDaa[^cOLfZ
9H8KFVRd/4gHV>.a6=K=R=N(_dF]6VKZ;cNFL.6;I&[.G;_WQC8;YJ#9J\AUT(^6
&[cCgD/,)&FC<PTf<aLT&WJ58eK+55:3V@)Q&d==(3+D+fJLU/f7?S2O].C8UV(0
f2]6c3c_c+^_Rc>SS0e5<2]K4:^M;&P2ZR(@.@#6dMK12)FX(YL_dDQ,HgBfR:QV
QW9;Hd7<GMB[KCX[]AB<73Q/\gM/B]=X4[(0]Y4K>.\NR..EPT:g75I^EG4L78BC
][97JM@Y&W(NCTD=dMMD)Kb[aaJ-#P>1EU@M,(b=Z+AM9KR/(5><#EdOLST]3>),
@S_779b6@g]cX54#aLP8EDE8]99HW(_./4OY<a>6-gBD(g&f/;Ke0abING[BR:Ba
3)]-gOY;HV@;a[FBc\1c@5APJ#W@fg@c&^VJ-aGP,ZCcge#fW51B#CO38Qa1_UU:
FbM;<Q4LUXg@X):?-M@Y_W_P2^C,]cR5JMI[.b2b+M8B<BH+<TJLVdMQ#06:2><I
6JT;-5G[V+a6dT,6S?3MeAa&[\C>>BBg[g]][b;-9J+B5^A,R&RGcaP@KDP&#SY-
7<OOC97VY9PNGW.f30LHKW1FQBb,:1?@ZI#\cA3HagR&L/AfMSM^gG87S1fSUJG2
38d;BcCHOWO<g;>R:A=_,5?P]JBXZVA[QM5ZX:XAS8H7TRXTSJ&@UF,d61W=DCW.
&PHE>GA72Q,2-O79c3;FEO<3ONW>]R1g1=5eS/fH/#;O=<_U0QH9](YU<<gW/8PG
MOg&cEW,,Ea>8eC7AaJ8L;b3VL.D[6MHa@N2R]^C3)5<&+A@9U7HSNQOC1J^(c5V
ZJ\3+&S)gAC,>[GN(D(b@EPBQ<IZDFB<_OHI]\2F6E5SF&L<GN;.De@DOb)/\583
\J?8beREMFbaX/WbM^6QJ7g9H69#IR8G0.U[I,-Y.URX/dcBCcHX^KHPKb[;U_2^
+c\JYP1B>B.KFSWS:?H4Kb)[R^EEI3Mf:>:^2SR)M=UGO.M]^6d-3C5I>J5gJ^F9
dT?cCM_30TS\>L/+\eBB]]ccYag@LHJ31UT-;1d+Ee-Y_.5F3gGI=D6TC>?O0:Nd
HQ7TX8C=If+>M6A-c?0Y6OaOb[1DGACY/;Sb=LObcIQFXOO>f6?LLK3:cKOUHV>b
6Sg.I@F04U>DKAOdeZ3VBdT108,OfU@#73X=XX]Y\Od64@YH8D0G[C1X\b)0KZRT
GgUH-=df[7)P-M[YaUJNR0WM6WP0S<TP\OWg7XM/dPXVWJWZF#P\>cT7APB0?-UF
ULaeIa>U5Y(=N1OLS#:GOW?U5AbY&[.e)8/XY:_5=/9<R#,+=4THB=@#&LIJP]B3
DcW9>9X?^R:_A56&c;.cK(NE9AK,TLV/<CNUeX_W.f4Tg,F>]D&S.2N20^,,ZNG#
cC;Hd^4G7fFIB()VOb>,#.6ZD((@JX#WeV0^J9.fL6TV[Yg;9^-Xg;>^>b]2:R,M
7-XKK#a2WR<0O?3CH8Vb3K_TNN&:[D+UePcV2A]dNB_^-BFSN1YYe22W9]J]06eD
3(.?e[fb_I7+3/f:1dM19ae[TBF4IaRR,cQO;W-,>GP9PTJTI.N9J-H;</XB^I+a
(<XNDNE9]dS^3?G?)A<=dc<;E,.MIT]K2Q+(2=T7Gg<3P+P1XCE7?WNc_d?5B+fB
AdZ@CLb7ZXAF9Kf<4W0U81<56J3TN)DdgFCb.#>/KbWDFBeeW#]6:[TFP>T_)A6D
WPG(O:0OCPS9eXM07M]ZCHA;-=PcRfZ99G]#+BH@AAVS7MSHSfUeWY_#P+R@&L5<
2)PV+1[e#67+\#HQd^e8>Q4A)AF968.3.f<P8Y;@V;Wc)+FTT:V1N;d?aU;a/)8V
LO,e;J=cS:OBCgP1]=58<UWZ7E(FcLYG1VTFDQ8eWb5K:0WBPC5/MZWEJHd)<><D
^2/R[&JM5f8LgcRY7SbX]Dba&)(b)MY):JUG#C1Df@6W5=1a:/9R^,Wg>(,+C4,@
])EZ@+7&b8X\a53a-\Ua0EU7A[&DSMLTPQ)OG67?:MZ@RIUE,0:aX?M-4a/@7IBM
c7fX.dcf)))T^&VER/;gD[HW\acT?Q)XBP2Ya)@-&K\BK)JbfPD(Z7e&:]9^A08-
@H/:9bY>\Z>K:&1f:S^L3d#>UDPFSV;4X)<^7I(^8W28CRC7Q^&]WbE&Z=@Z;gFY
aMY^7YUZKNWJDJdMeOQ:;SbBMQ4A]VdF(S0cW>cD,VYa#KI+2W_,ZJdPNd^RWFa)
961<L3JH.d+<deJJRSEb]-7b_O1?P2_T+#]7.X8817C^&EO##/=W8S=Wg^P)^]4/
XTggZ/Y.M/B@cZ1YK&UKKDNQ#70CeZW=NR;<Wf,Dd_RK+A>RC33\f\e[c4>V/Z?d
Mfd0,Ld/AN;P7E0f5C>W+S4[?V,Qb93G(S.2HK1(&#H<H+8H@\+D^)_cFY\BaA8[
<RA_CM8_<UD<.U9,36ARc#I\X/,^fC(EI14e#<O(/JOdO@33ZeX]=W>10\RVZ=4-
H?OT;LUCaN;<>T>)=eYC&ZWeIUC,J/g6g_:\gVR4,>MPVU^KYaV:?7Pf6##Z^]AQ
a&(>(P#S:f<ZePT/aC@:;J^;Z=eY-e-+FVI(BeHZ_&KAN;I883^TDb[fZI3aJK/Z
Pfcf8]/,:WNJZ?R@-\0EKW<C@^PbD&9W5<PK;^2:)S1K2<G1R?29_eWI3SdX@M6a
G9&a83=H:6,7HK0;R6R>^V&Dd2&6-G39YRX11a:5cK@;a\[K/O:6:D@\?5;19Ag&
K3aN.ME=g<VaG]4+1V2)GdT[.E^^fA:8<VOL#JFD&d1\906ReSdOE]Ndd@[3_f,b
LdSNe_Y>EEC105NLJb@41F4g?,O11O9B]aV^7/:IH/f\VA^&]2=HSS]4J5,eM1>:
]2&3^/c9TB\Y6,A?)b[-/HUe3CA,C[9S^Ha3_?HSUgOe&.(/[W/YD\Cg-/_]0B99
cY#_48Q5H>RCO#1fY=UP-^0=c:UX=G;4WW=K+/3BRZRgacb3AM+S@c[:^dN2I(d^
TZVVG6D[5#cZBXVVO512,N^XD8?\_PG[9+LQ>4X8926_3_^STED4NHHVdMGVINaI
.dY2>O6EPCF)2LHaeX)NMf&YM_C<0C?QOcB#f,cH1GSSB4aG?b)).-#(G3T1TEV;
UY(=;O8FEBa[?]AVTPA0(Y7C0QETW5DC.]:Y<V[9&MOPc<X,^#/60cb]B6&8PB[#
R8FgZfXZ:E>Z9PR5V)+(P&+WBROW0JA,-&RLaZEAUV[I6>+fd8OG<C_7N+I97RT^
-KL9=<P-6+^^X5:^74bY8F)5<+U;TR,;\dbc8XV8NHV\.:b<&=6SEe6d=ZX>)+\S
FF:8P#<0.5;RT6O60H]QY.]EbXE=,,#J4T?[A@5b_<a?]O]2(\&fL1]^R?RFGH&g
@Y/(R-0;O(Q1C_B7XE085CMK6[?f9H42f(JR29A>D\523Z28C@GJdU\Q^.S[G5b4
:F1.WYF:=MLD;8>7\S+)JUVG/9Be8b&&=6I;_GHfa)Y;5HP[cA<KZd;T(B7]>fg]
T3.Sc.1@7UF7^(69,(X_Z-3=(\)gb[bG)0I<MP>f7^&BCQ;F,N5;OET9F<abBW,7
ZC,5c.\Z:=@A#7<^,d7A_@4&L2Q,RJ.J)]\XR]cLMFI5_IP:/eNDRR3>R=C18f_1
\#W_/<YCFLa24P^c.aL5d=L>;aI_7>QT4,2Fe#)N?X_\W]>)^AM#B.PC@&O+;,MY
b\FPePfP#0X\?-2R3^K/R=>O7F=6/P^J5fd=c40E@(]d4a.ReO+2,]\HfL:fV9eL
:-V?S9#K\7V3\O@Y,2X&I6b5aB,Ba1=6^3caFDH1Ad]@01@@/#[XQRV_^;D7_\T.
RX=FGHW=-H?fGTa3V#?@P;G<c#<4K/@@(C@7(aZ_-aF5bJ;W/)D@.VDZ43=3fPPE
f+9UA[3Y)5d;W07b@Hb(KAe.:1R:a?(R,\;dC=V:T>B6,NA6&_U:1+5LNB/-:?BI
Z8R.b>bLB?O5D-ZN<1W_2WcA@ZFUD0SUQC\/e^G13/aS;K=K1IMU)SVE0Y2)P0\^
JB&Ab/+?[D]L9a745MP:Zf0\E1R]/\)3O?LF(2U7?0]bN1M0]2&_)7Sc(>FF]0&#
L4LXa,5W(L-N\I8I[gGd6<;@T6f]2ddQ1dQION?<D-.DFLY28>V\V?.=cV4X=BU@
O1;&:fG8C?])HZJ15:EZLKER@K^d;V>Xd/8d9B6-+[.2UDHO#/()],)X\+dGdb&_
6=OG7d9A6EW-V11,6\&J^TdbD+dM@L9#6:1bN.M;U@da77<_0/H#Q5gK==O,TNQ+
[:4GQHEe.+#Xg#E13TXZ+41fO6NWa@V8U45.E=c-1#g_O9^Fe\A6X^-KNLCO.ID2
NRVC&-R#)S&^.2.f7VF_.B:b\)JR+2gR0gObBBbTS?2)B4?e>K8-?b^/9S2)faG6
KZEUKV0f+)_07B<L=(aZE7AE;Q?A;@T@S@2GG8dTUZF5V<7+f4(S@-67=c47UGd+
gL]YG#4U,5L@E]])NZ?Pg3HH9:8/F1?K0?,5\B\=>03N(A7Oc9V<JHAcV^[R:(2+
b;e;RY#0IB0CQF])begW0[>abDT]f2@[99,ZE&cUUC_];20T3.R=We0,IXb(#:GB
M+6QL1cfH:d^M44J6]R(O6f[KXK.Q<b4\08?M8&7IHI-.E2BgW8&,IM-b+aZcYHU
9.#F2;_F##5e4JH@O_U2M_Rf;#@@_SgO,PXdO[02-5(E79_CP=f5PQ_.1C[CD=2\
1\8@9RF\Ef7Z9&VN#R<IIf<+MMd944VNg2HS#P42SK<YFeMRf@VELBT2/:4UV#.#
JfD+Q0b>a+99N5gCY;T9,G1IFfM7gR=\J4:HHTHOL<S#FJKT@^B[8TB0P.RRP0-H
4@EV_dK8ST()>d<cBT#(EK:30>.LbMKH5,LB\P19&E8;)D5SZTfF3)e^?WR/f(Z9
,3>;-/LRGc+FF[Pg[Xd9:Sb>H)UB]#,[TBE<HIEDA>g@L8>]Z,8>EWH=3dU+?><g
=e0+Q9,@eR5G>/VM1IfS7>MN=O9@.E(CU8H9JM/AAV9BX)b]XY5#.++.XEIH3AA?
K2f;\<aa,/b:L,OFXe:NYg.8R-.gOR,WgD_-5@&N[;:^Z.M)3KT>Y<1M0XV/W6&O
..cF7A(:g6/8R->A5\/\VPC#^Zf#UG)(;c>);DXFUb+M<a+fQO:2bQf(6-/ZPDUW
^MK_8VRU8T/#^TPL2C&BK&PdY7Ma3HEOSZCRfDY:85EQOD7\8@ON>_g<6;YeEC.L
,J_cRHg097DR:a\<L_57PPOKTVLD^aP\,IVT+c8;&==[0ZK4GRHZBFH-XT[B[DRH
NGD#2=Jd31.(Y4TWR4YK(6DfPI)[VH,cU0OO[9D^.ggJJa61N/T.OaX&D62+\T#\
ZbZ=FJC5+WC3c@-9d2+&SV.8+;9LW2Ef^R:&]f>[(5#2]UAYD1I:Rf)-80OBL.&&
GGG#HU+d0//aQ-?9=K\,>AGM<\>GEd(58bY,=[K>ecRDD<2F)C)4V+ZZd]V2<X-R
a-aDBV6/1:LOJ65<AQAE]LE>)+WIU)Y/cYQU@]STSO5J&aY]>T?0OI?ZSW4=@6M2
A/V<R]d1[;8+<.R60MEQR50/2&IN5AdO-PMG28&Q^TV?MR.+T6M0(?:6Y3YXP/EI
ULfTJ8(#\Mg+_8,[d@b&(8<_FU2#<,E?39[35Vf]@4(Y<U;S/CQ#9.=(7;\\Q;BI
?W&<J8GI8cTTJGUGC>HLV,ISIK&B;Z0T^-(S#3Z9YJW_LQ\9(G1FG&NeUC#T1.#<
3PGQeVf8&-H]UP01;XdT_F&_VFX^-.[:(^A@@Z7@V8aX+<Dg@e5Xf6QMYg9Wc,DT
CL-HA&-D?38)4OI1M=D3;VIa[cCcF8^C3]\(OWT1BUdgb4WQeDWUT<Y26[/2.BIT
&3\8:MSXJFX1-I>.#cHG3U<.PG9E5+f\<\7L>:5W36)7:D&8cF>e-f:QET2a9aL(
J(]_09SI4[KY#)5GOb>C2-QL?\gR#c)NY2<R?K2MX)6T-SG^#&(cf;7:0WQ&3P\=
.0]]L[cYE==R)3X/>dJI0FKg<<,Ec7<?S\=5LJF+Y?7KcAR),#YE,6==^I+L39W>
0#QJX=U+[VSM4.5LAGLWDVHM4L4I@VRd/9;Ve6AV7V).;4[AM+\&5<NC^BOSMQ:+
MN1+b+9&b-eHGGfaTKQc4R#),:]&?6K^T;bAHN7cZYb+AX?_[?(V>O/X@GQKYVG]
ccU>R@5dX0X:-MWL:M-U;&;[+]N5DXD_P>CUe1#__&]Cc?83Ed)@S&7e8KW_)0G,
O/;NOZRHW+a0dTE85KLBVN,2<WHA]c?]^f&Y<6A&(aBS.-MBSPYCCE2dPZ6G/X7=
d3;XM;7eReH?A&SV#4V_]MbaXU[IY4dN^]^g^@JCO2W+G^DgNFJ.JLT)4(-0^S(:
GEG(),O)N1,.A0YNT8OcU^_9HO<c\1e-1>A7TfQ)>,>.@-5EYb+K[/<#)D._\9.5
EAbe;7DNeKZ&,9,&^aN)E_A55EB-6<fX5:0-]E.3W.OM\5>42,]:2S#)2>@cf#&P
?.^D2HbYY8S2]XIRSTa38#VZIF[I)gRD:EeBL,;CSaBf:+e8Va738Tc7e6O-=/O[
6^2]/^f)?^<fgDa7[W#6L,99,3YM5)7?K2R5G:gT<LSdPCC0?eb-S3aNCbEL5FAD
e8K,=:ace?4,][-2G:]@-J3S#=BBV<H\FB)aF_1[>E&FP.bK.CDVL/W.d)L;YMa_
eQ?:1d75c5Wea76b#-&GTYN.1A^H)#&ZY3Q;+(Q.b,ZGPATUL]/eLL>g(34KcA<W
eWL31=NUZ-eVXgEL?;/5-\18D&7[(F)Q]O@7bR3HA@KLgU9#S2?U)P;bgM#L6cKB
UP3E)cQd6OFZ5FK4&:I)]JAgF5BGV<F^;&BJBBCA8(<LeW^5F/2F;;A[aQc#QY-C
Ba8@D7;G8_eK\GB8g#R[gG5=Q@](M?N,AacG,Zd7#1D8W@P?JRHJO]2&ZGPP4d&A
-U?_T&5C?^4#7&84KKIN-XL#e;N?:-CP^]?K6TbB#H(<-K<d\E:BMBKRS,];8LV1
&>G(_(U=d54g:B>)eA2cUHB1\Kg16;NL:9^H77F.S#a=BEg;XT,3TG9?/aC@FHa_
AR=>5)L.XMZ,M262gc@R^&ZBcF3>:KE:6+H^^7ZN8CX:<dd[UBF3Be2YdTLRO\;3
6gM>Y[P=//VB(eYd4AM7fELOX^Za&OASSU\aR-(\H66]9A)8O5&S)Uc<.#SL8IV+
F0>?C8R#C_W^XHG3U\F;&,Yf:S+(B0X+KGVd[<CMEG3Lc(?J/ZBOae2f^Z]bBEWK
>)c(V;HRLdA<<S4G^_@[F-QC]Bc6/Ig8ZIgc8O0a4^f5+X#^\;=WUBRIL0A\#ab-
(<9^efW45A0Mg?VJ):.N/32&eD,TD-Z4L+>.@D>R]cUXCdTHE5V3B+([?5CUZUD@
Eb60;]W?0\M[M]A5Ob;S><X2fW],W4gF6QGZ7>ILWA9J/Q<)U(J7NSZ]V965RH3-
]90J[3\^8ZFCY9V:44Sd.BIYd[(E_AHa;&)76M.7B?CN\D]HY+d)^44LV]YI7P]@
F>(;UG[NEY0Z.C)LK,;LZTZL&ASA?X>bY#e.HNeFL9GQCd#WgV0MFO38NbHGD>V(
Q(]Y\D;]<O\f8AM#/WQ7B<IEeIM/e#+6MdOXHYEg=R<BNRB&f)O2GGRfF+/=5UOH
M.;<ZW7II(#9R(@SG([PP+28()FOL9G@+^HIaOE4LOT9JQc7GY[NZ^e,X3[=cY<.
6MT^0RVH>]gLQM/0U]]KFP36,WZ7RI#@5=5_9^LOIBY]\/W?0R7TZ;g?:,9O-]d7
15YPP,JV1Y<F(4D6#@)//02&8M0E0PFBf=a@9]_Wb)eE6Qa+/\H_^A<N+B]5a634
fXK9IC#KbKTbC#H0C._b:SZ.-^bA2-+KVVTWFR)#9>R.8=P@)WR.W>,7[0_/>5A0
Yf-0)UfONZKF(+I6]K<_eK:V)_1AEZeHGVWK/FfH>?O+Ve(MZOR\Q))08T)B?O-,
]fVaFHg@EJ^-<K:\P3N8#YG+I0^>Y<(#W39)</P3/2G;#4bXaSM9(1O5eJ>,/9d#
PJ#Feg8B<cGcaYP-J1=4#L>IaNE?B5J@H/4WJ7651IKRa-24?7]BV3@/@O_<^;DA
A((<a>2.a69DVX:HNQ(1P6ZIUKFE1dI1TV]feLX@_4g7T,+^VT+Z3RU4)1<Z4U,L
YVGXSWD#EO]d;+AGCEcI]R^MFRF(CQ?UOVP@4159/0Cec:Vf-8bQO<;(dB.Y-g^,
-T(MO[11:+Rb@C;fDCS3W5-YLZF1=HQPYg<9[;fU_+V)H;B[Idb\;QMfc<D^Z4K&
:1<gIB\B,OU,fV[)>Z9T-/G6cgV+^6(L^.^P27@BGYLX:UTK&UA>B,bEIfK>[OIT
4NP1UB)H\&O74Q#8L_>2(LHc\L^[27].OHGQS?WXe?S?@V==SD^_7-0Z>]A7_^14
L4?9a3C6CO,agL#4B/dWC6&&H,O_QK9ZYA)^Q(QBU,IG:S45X6MUfKdQ:\76bcOW
YZAR\54?TUOIG,F72:bUUCV=OI)/>QDK[QRJK>:.Da/T4^U,ZTPA&\0YKL+6]C+F
WNB&;dP=CYg0,_EFAPRa3D&/:8F^gbdNLN[1eT3#:0)8-c#dX=,>e[\_QCZ+<2c_
]4>1d+K@(9N5((9gE>e=Dg:FQM+HYR(9Q]N<<BP:(^)IbOP&Ka8XJIC&;6\N5HA5
4JJ>e?&c+BbGeWcU9WUWA+I^NK\U[V-JIK0>BX=Sd9D6N,BIH7-)_VM#ZD7H?29>
J^OW=VgV+.Q,E-)WK5S,M)LJKP;EON1+R9>U,:JSKLd73]cUR9g#5<8X7COf]U6L
@fQFf.SF75ceH;F4W1YEOeCDTKEX5MY6Wb\I<EEP;?SAaEX@VbSX;eI3JAYI]X2I
AOCL?C:?A?[KH#gG:N[(;@KDa:EPD7Y+UPegI8A5RbcO[;[e3f+,2?f_5?RMF2ZZ
WN>SgUeP7@=)N&Q[,:R_+B4T2C<b42ZP/TeO]BKXG]ET8,YQF5L1NP9g1RGYUcCa
XAX>AB7#?@S__\_<M^_\cV_@SD.W#HG1C5[MC:B<L#TXB8fRF&L[30a;-7dg76GF
3O#K7GZ,[9?O#Ec>\;dFAaTQ?bA[PG+aTKT[X_&-078LW1SB6.3_>BK/-?<d(gGN
HR9E[P/7&_1fM8fOG8M@TZaJKL=7JE30]4-TE\?c+.RT&I=1C;TY8[Ea;_K-:/NT
+[R75]C8+>+b1Z,;?f&BCARJN65d=P/bFPZR+T-E?E[\.03N87IMJa;LN?70&FEH
[WbPPJ/WMN]^SeV5B27?;TJc/a]:/ZTGe<>OYeH[V)PbM.[BYV;eYFW[e8QDZ.b:
5T-b:/WSfO.eEC3b@\JJ?FX3:F/(OV;^a);,55GDM=Bg&3\)]If\5,);R7EQedE7
F;\84<L4#@FdMQ1)#WB#a0W]HNTBc+-.-BUL[T<PP>UNS@5SbK)=]?L5dM_MP9UZ
K),XKGEPAN55^OaOKO4.FIDNaA:KLd]g?QAEHaA6RD_3cD6a#bWV36S8dDg].N>.
CE1#/U7d/;HGN@50]D.B>(X+8eHf-><8T.7IR;P9UDH[M#64]KOQOdA>7>MFVW,d
5TG?S6,B-O]Z82JZQ&>W/SS6.<3#^Q<9WF?19#S?B8EB\#=IQ.YIJATJ]^fL\CME
?PRGY,;f+@71-2cTYbMaMdM1]dZ[cAP-^42Pga\&?D-eEEZZQ[^-^a:US9KW2+P)
EDYF0T46V2&-\_^e#2=D.O]GTUE2_ZN992[bQB;L^:Ic#2FaUZb9UM2eYXb@;W0&
&(BMHQMBG1gY/_6C9[TA;9g?4FCfEE?J-c4W2T?gU;acLXWS&FU4&.5IK7g,?_T:
D+WKS8](D+,(gL#41K_fXT.bFaBYL_2K)cT3;P8/VZ45Z.B:F#c7L&+[]9f:)[E_
K[CSE0)5):9(QQ0;3ZX;K<g1GN;;>4Sd().ZfI2\Q-P#N+&C]\\OG=UYX,A)Y:5S
8QG#8fa:UXZC7<OZ-1A@H1J=Y9V4:1MgD<9@YPA+R=BZP1(2+K-\QG+e65Yd5EC>
O@V;4TA7XW4>:H6:;X0)_G(V-;?e9^b5ODL5;M50f=_522NecDV+c:?.R\7]YKg,
9g@[GY<c:@cR9^L#,V]6W0A;IPaW/Z4Q7Yf\;NK>f@77(ab.6U\9@@4GK<^5Q?^a
^I12:KaG+PLA&-;G09MJRdKG+;^1@WC[7/0J9/Nb?,I#QU:Z&T3eU<c9cI1.IOLQ
O?J5/\]gR2][XdMC[:^=J<C=PRBe9QV/T6Z:3-1^I?+QUU;dc=;ROEQ<<CceUSL7
JQZCfBc3B^]d-[SbCcT9#F0W(Yc#M:e^::b28=D.V0R_aJ1<KU9MNOQ(90@ZfZL-
M7=S3:EfQJY^WL2V[_^:?KSDC#337FF1Wc7N=ANa],7.\gN:AB8R5d5R6M(e=2#U
Y6GZU]\-<-aHB\e:7TB&L,0+L9SVEd3RCJLe4:=?EPa>7#@J3U,DBB:10:<VI2;T
G1USfR<[I:AfY?WIC,@S;T(/Hf.H?@;EgYb7X_[[?A_WS]e]RQG9R>a@YNSKA@DP
+YNH@(+=R26[1B&=Z1<P_O5VF1;T+,?X,A.6<.-dK+g;a8)5ZQSC9#P].)@+8Z@)
J?+OB?:K6W74L>fg5]=?0GWO?<L;-+K&5U6^N2)e77@XCU(N&95P]1TE)]VC&FVL
==_K;2A17Y5de,V1Ad^)g@RZ^&P?TD0Od6<feFdY?eLX_:PWU.PQ6ZaT@7,8Mace
aQP1:0U+Te9F?DdQ.CEK#a=I)2MR3)2\/.N8#?UdVfMMYR+e2;[e0ZV@<?c3^b09
N=5SeLNNeK\ALBKYWgW7JgB5P5YLBO&Dd:Sf,=a(G+L(3If+eU.QH-M<4_bW(\A:
)(]D_gV/[DCf>RA,K-^[>/b>P]=S;PAMC+RKZLeF[-#_T2,EdcKeB^c>C3+@QJ#^
IJ&[ccA<A&Y:Za^3^(2.dZNVZWDPfbUTJ]M0N&a3W0F3I)7T/E7NK_3YP_9\+4,:
0>=D@/NL,GC6UR:VD/egFcc55P1_UggVIQBH&RWUCNI[5?,&a+>.XFN0dX+B:+&#
e,P9YYLKX(D]JY+HVQO0V0+;d#[B8Y^QUR=b:UO;/CDTUYGU0O0^A?FT(R71]8/.
,=Q:;Z9;R,^XL(d[TF6>B)3d\ZP>XM5+Lag&4KP>UP=3ZWJ7M<^XGD@8MF4AT;)d
@]b.7B,Nf]bU]L@6,0KHP+Ye16@WI94OZf;^fLS1\U]GABc+T#^NY-7Fd)&(-LV2
(d+YMTX>cJaBHAI.5?MaQ=-U-R:5<BFUY.b<^TJZ.FV<4)QKG(\0^++A<c_#^66O
KdJUA7Mg?4SKKJV5UZY_#g,e>1+KG8](D0c5<LfS[A;OH&J<(<a+G#7XZaX14EVc
DX;C<a;a;+WES@]R(A-J[gS5UM:Q)_Qb50Z>B857+RPNMg_^HW)65XV+.Q1bcG.T
0@E>@G1<a=>a/7]>BQ+=#R4Mb8g@9S_OEb370V-5TN=g.g1<bSX[1+e?8429:7IS
X7KK0OCT=)R_YB)g^BF.3&T9Q+1ZG[DQUWB2@6eQ7/56>N.E.4/aH^?89S[=SXL_
\JcD1Y+;N-=PARUFR21SS_[I6RNVVJ/AG(.5.,NXH]9#?75(aR6FeW41DVHO-3:Q
=H/PZG+a]2@MQ[C-e&ZR@eV\Rb?6K6AI_Q&)(FWU@gfG<J;62dJMeZK<503>0E\@
EAELBT5cLVK_45O.0A.)F]&#Rf&Z&/3N/M@-6?fR9^;34;]eG0+5S8;0(M/]C2?P
3?:_N@Q_BF7^CAV4)>db1M)3fV7;N#c5[LV;#ME]SYf,RFV[D:B>+AK/V9#Ycc0/
@Y,@=gK^5XY4I]7^?9.M:>6\>\OHPd1,9MT;46OO-c5_Ke5UA<09fT+Zg;b=9RYL
A<S/FIaMcQeVEG.A4g4REUO;:>bJ^5R.C1WY5M304&<&P8&J59+];R=e)N7Y6W<W
=Lf&67/Ya?dX-RKPM1>)168R1OYC/\@CFR5>B(6:8CMXeg<R\e:J-M8BR,L\D>=&
]ZGDFF_&MA&T#&8AP&Tf&/]d<.6d4JbgHJTK;gUTLO\GX[M>TH(OcDNY[/AJTKfM
g5MKF:FRQggY[<]:TSW&IO]LR-H;cOQA(bFeLM[V,5;eR]a3J@c0C3(4.g@X^]LO
(9cEX7@8<VK-DX<O&Uc=T8DMFBC^Z6.(L:CN83[JT:1&)CJ[9OITZEK4U&#/<ZBe
12\,U<B7>^<,/5MUIb=;IaN+W4YV[S.O<7ODD()MAF+F4H(\e3c_Z5Y1J.7aX0Yc
U.8_63#M(7E]9#-ZT\IMaDB:7?XOB&T(/YeaJaV,gTJ--JfNCBH5U^B+bL=SM2]c
AOe[WQKbPEE)[P.O/4AP/X8KM5fNY]5T[_0WFJN-FJB&T^+,9:1VL^)[@;0@aAV/
^N]4M1ZU6VFTYeOFC5H?C_>HWc_F]X,N9Qc[_M/dNBB-\8c28WbK,R_2Ee?@Z16=
bZEb7&9:D[/[)P&K[(>,.SdK#(g(=C4\IG97W@bV3.(1]E6b3)H.91-#/dYDdM5[
.9LR#e4ZNcGQFJ23V)Z+(?2LD&PTcCUTTbZJORgV1,>&Ce.L/YKLY[Qfdf\CRf19
b5KU&:def.cFd1.D=6GQbdA8#)13HUCL-^W^QASV&_B:d#BQaB/8g-+;\_7&<U:7
H)<QX=)\S+@cb^G(<QSaPeD4^<DAJgB;g;#KB(LO5,ReWG,;Q:>GWQ-(W;9HZ<22
MV_cX.(:FXTOfKK6V;?Ga;+PX>=WO=1JA/@]_/:fEcVAbD;FHAD-UYF6VWN.-XDI
6;].LL[WA2P,2dW5N==)Z,(&58N,D,<)@JFU6baa:,aX#aLO5C-P[=Pgd3)D?WG)
^6@=Q)O1Q\\c_2DP4N0P#LY:V/edP&519dG=fBfZ<dNJF2G=4d0WeTaWM/38UQP[
]4Z?fd6B-BcG(;=RSIB=[G,6JGNM<d0=N(Z)[__L\Sg-6ID?bdS<FO6E>T5::a.4
R)7J;(AA7X,#A9MT[6.^2Y2:^S4e=YD\cPGScGeU.=;>((8bf&D^Q,bPXRb.N6G9
_3Y3Q@>96G&5<f8C:6Td>&E>Z/O,H7N@?75[e.3=,7O8)_IBV&UL+ZT&_MWP+IH7
\-[C7JM,\Z8?,K[fY0>OcQ^Tg^fH<f)8_+W_ORfXM\1S9V;9CgeTP13KERA,W94T
<,.#ND3=08HG/YR/3_Z?ZKeCP4S40JXT@>.K[5PM#+2,@4cJ@()&08PS(9@E8+@a
CX@ZE;8g-,d1P]L_:;^K=JM;?06INHMEBe5=fGI&A/WI]aC[2LTC]@W]T(P.dHHd
GSM2>@XAIFLZ05Y+PO/IfT\@<.1]RGa.4fLc?=Ec?FIF\[Q/_L]3/@:MOd4LS(+b
J&,@(&NH.c^b9HU-M:E,?Yc<f4_3/acT\(Y5/g6@Q6Q\W,ZdcU@?g)4[0]bR-G2c
KXG42W1_D6]KE0NNfZT5=Z85#+WDPLP[X5+eUYVL@80ELEG9H40)36,TaE)J1agJ
.,dF_?(^>9P.S==fV]XY^;Ce7\V?fZ(LS7UX;_a<GD,[,bM@aCWV(T0F:7Me-4)3
H06c:,T=16#74+93[1XY_AUV1AgQSe-cAWWAZA#QbXE-4E<cA\T5\S,(\)#O8577
=+,P_^a;Id46BT_]L&ee4aWg.4fg7X3(:P4\bA8OVZP^=][^Eb-P,g)g0c8TUI3<
\G18_-D:a5&/V>0TIN-XNIV(8+_/ED2\[_ZMBKa&c/^E_.SS:1SCNd?Q[CO_G^L^
;IOIe0G3E_#5<cV4JB5.cB;#Ob#5>FKOZeAEBf=,_MWEffA=8Q.c]DUT8fP8M21#
N;I/VT7e>=2:6G[,AD+-@E,^K)NTP:0Ibc1.K&9RNMA6<-6e8V)6/^C(:BT(6=I=
9TRJ5;C:9dR6Xg>4e/+EF9NX_HRb0]06V+X,3Q]BLaLC-R^16QB=Ja@d9a^fUJaW
>dFCM&#,7);(?EbJN<T59P;-fb[05?9(FXWSONGE\T@YWfIWDAF;eF5KA=B]bN1/
da;D=L=b]PHTB_\=@H\BZO[?C;T_ObI/M,A,T;S&U)^6X,R>_7DRP=(<:0GeS]_;
DPNS&S5W-?OJ7(@XKg0UNg5A6d):@3\[M^(>]__HRG@#.9;J3?E_]c61fV/.f[.b
a:fH9g65JCceAZD;6M.fS:9<c#U6R89:VEN?4@Q/=WL?3[NXHA3U)Y@?b5XAEb:9
Oa]R/AP8#S/,]#RX?_<f;Q<gf:_LUPN,-_JKYW>Y#8?UPPcPDe@&=HN0RgV@^(G4
1dDQLAH3GLeF>[@)ZUPA_WB78_3,CZ6(P;XaeXKS-B_7EQ=Q()cFFg.a[-ZCe,BU
4<=LOOZNL=1RFF.1XCUIH,(]9aR0K@UGL9PcZ6072S&<>;Q)Xf-I_G+_4/#V>[M<
0QZX<5UKYa4\J<B28bf3EZ68VMXBNc5R:Id3.)Z/Ob>W&<>QIQSa0+<aU>,fM/M7
8&aFS/,7G8]71McCbN+Q(M,.@TJ_-?Fg+5>A4E9#A>11PW2JR(bRF?,+\H\1D:+g
BDeKB]74Df:3gJA_NM_3+<GTVbeHDg?BJ(4#gS)\&P=>XB6X;1[CX=#\3bg&D5=T
ON&(D[[P]+.e:3AdM4eEdV.gFE/dBP#^WO5(78^\;>Z^<+@N]B3OKBXP,^@\?X1]
@S5W0d2Y):-NO2\;e\bTR7\:e^+H2ERY0T5L4UZ&CN2-S#.0O@L3YDD3;cMgeWF@
L.F^P2=/Vf\YRC>ge\:@&+.25,DRbaf9VQbIdRL#,#FO,a@PP7SJ(L03gG+9D1^g
]X52]>L:c<e9M@&B;/NWYcB5A@/;Gd\_X>WPW;7<0Ce1e+0Za#3/g9#f)Fd:f:G2
ED1B77[W=ff[I[#SP?BD0g3+aeU&A<g/27UbP[H,X1BS;B5:7&.OHF>U.XX>G8UD
cd92BFYJ)-fD45Od6JWDVDL\)KdT?;&K<F;Ua1=TQ9PJL7Ycb/J29:9&VPe\4+<.
V=F,/(8d1=[2IV,052PJ<d)CAEAUWG9/a&-7:MK^YQ-c-7V9&K:g].+)19Q]48C5
RDOcbJC=KH#.-7C[E.cU7;aLg&\P21>D(<A?W(_H4X47U[)&9RCaAS=\f@S#94;O
4K.M_5d>GV97(RLONC1O^9CGL^)cLeYZ863Oc=d5.=a[L.1ED5^_A\/9#OeP7Yf4
Lfe;_H5\?RQBJ+f<b=Df(.\>6fJ\G<B+GG_.JR[3GIDGP.481<)-T,c,db-Z#GJD
;RFNJ5QG^=Q0D/\.^Z#&1#6B/N7a-2-KB^F9NW;E-Q?7Q>DIP6IR.\[5HB0:B:QF
/X>e>Y9cK?+?/;2(R()e5/N#=P]W7R;J)WG_POCA<>Bc?EUeK(V(-Qf6D/1L<?2-
^C^</fA>P_d1O&^JD+e-e4.<H;J#^<TT\ZdY[MAaXe)c74ZWBGV]TT8>>,NU=KG:
_acQ[<YDSYdd.U-Y>)I\63:faF:/I2X5L;B=>_4.^Z7<_bQT^_=+=V;5W2JL5LAX
TJEU^Mf9bMUdbf1R]]1,ME/54BB49&U6X8CYAAJ>Q/3ScTffdaJNS(,7CPKdegcO
8-eD4G[&SWf>UWN_8CL]3V0C2)W)eV3J+L@)J<ZJ,8RfV(4ZRgd<1F:\2T)-If_9
Ee^\].#g?G2cRFgb=HR\F,+9]TTB<b19W\cJ.-T^9+B@\TMI.dHJ4)PL2\(J_T+E
d\K(D?(3FNP1V,(gD6PWa6W>(;UFU5aa17/3]&=b-QZ^1bAC@VE^]3G]S5B+87V/
We9e6S/:7S]>VKF9:S&6&158TFFM@7E]2L==6/7W#^QETaa4b.FG.NBG-SZ<YSgL
dT&)YH6?Y2Q,3^Z<:?S>8bL/HS11J[T.d+fN9Bd[TCCH,W/;=R1<-XIP+V9QD6=:
6Dg/H-6/.A8A[5PfVZ#,Qg5dX15f9[[;92#1OGFB-/_R+FD)P>K9OgRK=,KH;7R/
>]M>LK-V0:<>Jg^/ST6;DRU.2+#;5bI;E6W4D5I^[PFYBX41aP5/DJ\ObB-F/2Na
2<E8RN;bcL?&_Y5\WB\?XMa,GMK?We7:Xc8:gLb9QME\dLK[1dVC&I.]><7Mc7N=
233HY86de@-36>bFQ<()WBfR.8V-I:?G7;81XA)/T=(_FH+MLQ&\2IFOM7?1MVJX
3&G3X7.]>99=:T7_dM/:3dY<J\C,9=HN60AJ,a@X;QR4ZUGMAJJ1b(ZST9P7F:#Y
SBc;G.E>^9O2L_##E.cD?IV5AD<M(NC+=+4c&6VRYgUcT\b-Cc=X4(U3E8bR0e.D
aE41B#-+HDJ)@X4[fd]HDLP+R@NHKN_?J;?2f,?eCXBM&#P)L4XIS7YP/,_JE3bJ
L=ZR0X+/9XWJUM8\]S7GDbWND056O_30A/6TAa?6XOA;T1>/62)L+=.<([e,#=NQ
PdFAYaWFb:K-cJ<.)(43[>8WaN#Z:,\DHcfQ/U.Fc1P5bQgPWcO=X@3gS:E;OBEg
&V#[PYe<?)X6V0H<QLTW,_Hd.[[P(-ebG&I]]I@4NXDF&<Ua)@Z@JgGBTQ)V96))
95g.Jd+94NN>9T3CCC16^#JYEg=4Yd9-LZY>Z^ZT?eL@N:L]X=FU]Q[<W3US9CbY
2d2(E3UFfcS6(Ub4X<CGH@T?^5\A7&0bDXI4LeW?(1<[AddeX@=-L:GS;Y9bf/,Q
S/1^EMRCWA;U8\Vf48S,?HGa3I[3M\b[ZBLKY=MN4I7cVP(0?L:B8EG]WB)?1XQg
f[Ya:?^S]P;e-G+\PWW0DDa1^McPgRc8OVI&c)6>G@DG\9e.HOVBJR[G49D<VK(/
8Te.=gMA<<I/6c/Y=&]I4ZCF.?VE>(BZBL2^dD-b64gO4RUO;+XSGUK>,1.,[VU0
I8MIMR@3\>a#,Y:VYI[70#6>T(Y\YD8#a4e]6GJIBN:\>3)#T6He1?-LE+-c-A]b
<D<=[(UPL2aN6:bS/C:EAKQH4VB&H;>O#^S<\0eeg[7NV[P#/#Hb+?aLZGfQUQP6
;aBBEV/gYK1=J^<X91S?-NHQ\EA(ce4?5&F,(a@f[6A8;R9?c8;X=gK35;,2BgN#
/XX:\(NH.d9W)(JJ.W=THJ15EHg/5?8;X0I7?MWdAA=E0,GQFK=bI1TD[;c[<.3Y
BXaSUN9S-G=<>H1?9cR\4-F@IZeY&#3]RL2^c^ATJ3Bd@Rb1RaY]XA21,H0]]/_)
2:/HC1(<KRPe>EX17_7&ZbWRF-VYX/Y9cSU;QUN2O>2_OYbH#2:W>/D3JJD4+30E
U?21KedeB=fUgK1)Q6_)0]D0gF6Md3JX>Z1VI787AN9Fe@&RaTA<MMTNf5M800]c
[+3)b(\a;539-fHOgRfTf+8#D/7<dB;L&=f^\b7AVALdIfIf6GTK7]>O&5_\K-VT
#M17Z)12P2WU85.gF?0R)@Eb^NJeFWPd\;Z7L_cM]0+4OJ-P19QK8fEHX[EJOB)X
6(/8\=5gS0eJV-##]2gd0:C4\J1YAC+WSWW2T1VS?S8:G4c:Bd2=Cd\3acdM)bA.
H;bg^dTOV74bQB@Ea0F51IPLV9H5KKFUgQHQD]C):X2NT@1=&=(APd#65V.3<)X0
NG_^2^?LO.M^__PHB7MT[].,FcgP;ZQA)QL]g@L[#7]1AL+KUJ5F&(N5eFKD<U>8
[_YZ<H,2dLd?B(@CGZ6a<fZdG<8P/U,EfM7P\be,d&4,#O6F5D=+?4(9H+dNde1f
#;4/7,SH^C6Ig\.X>NM&#@W\S]0:WS8[a[.-(8VV2NOP9UD@.0G7f_V8dA9L?KD-
Y?M0-P[G?dSYO?X[5ER@U7S=9O_1T3I/)EI^R-4;Y<I](E,3AGKYXS>aI>MRY84[
A^B7WdQP#@0MBK=^O-:gL6\:bQPgR)/YVM],C\MH6/GR/Bf:;Y17DKddC#?R>NP9
F;U=X=M[X.HcTEMO1J)NQ>5D=Gd]O6G6Z5><VW>S#,#fYTPYF7,D+6?Fd2YH]VA;
88U);LIJ)Y4LSUcTf\=>g3FR+X;,UV;gP.+1]cVU@/HMDc.1@g-G9+^+Xd(MCMG&
MeLcX];O2#aJ;48RUT9\f4<^8&N0.X5215[]Z15YERG4-BM8]2XQ<40f4\),LOUd
:()B1/IYL5?08Y0^]-B?11:[N_:+A.P#66-YHH)\LT,fK/QT6Q+@A/M-88N]^ADV
&3]6G<S3]D8:D?.,W6@RD^\3I\C-77F4ZQ>(0-8KP6:B#ZBHeb(1X@JQ:d^3c<R7
9:@YWEAJ1QH;.fLNcg8UeaJ<M_U-<RWTL[@4M6^TKVY]RE(Q,509E?EK=N]bc+aM
873SK2M]>VGLH_RBag0&fG;Y;Vc7C.[gH7Vf,9=OB9Y^(E/38f.U;8D2]=3WA;]e
3KP)=5gA0#=]DN6B3.BaDB#T&fBRg>cg--=OZC]Q.P(&f7H;&_:--YBEQ9fg2I/Q
N5IWK=Eb4=T2b/SdCM5PgAQW\Z?E2a=Z2gCPOb1;>:5@,Q?A60&3X+.V@O-C[^QJ
BH]WUU;4WTFP777U:CVTKQP3_:]f[,Y,R/^KC/CN<)f(Oea_@(B=Nb/Y6HWEWY36
,O,-NYKIdRXKTYC[F;-R6W.GcLI<<.<D5,9-,fG30TJb.V8]D,9.F]>,VW4?78ZK
;]0JD):U)[/SCUfBf1#/Y:YN#bG-(bg9+9eOZX6UEXIKJT5Y6VTX1=<NB.+FaN5>
QD:J?,+)>(R^#0YS#;Ae>K09?C0KK18CA)9P(85Sfc(MOP#D1B1@;ISKadO@D?@J
D.0cG8)BX9-[G-089S,JUIA9KUA[8OM8MCG9-I,RJ;KT_aMP.N:.39G#.BVN0Wa[
C\LW/_ZGIabdLK>X)M_U/8\GQ)8F)@eC?Yc2Gg2EZ=M(R7@9D<K:8cCE]GEKfN4S
/FT6\Q6a@]-VfNcJ_=2CIS2EgAX]f=S]WCX:Q71RU8&\b+L4(Z+3L;?+,SL=;49b
HH1Y&8<b36VYaU8eQKETF9S8M+9[R\bgHVS.g[S(JcYfPI1I-W;CNWGLcJW]M](]
fSJgPMB51;M^7Ta#?IB>/g^?f<OGL38?23DbJJNZfA>H^PTJ[>.2O2AWX=IT;_>F
_>LT]LVCc-/:3SW@\O_^PCEY5KBV8#Y?1cf;-5Z2&3bf=:/9MX+<9+V.1W#b;L,J
@OZgdaXPAWLKb(0?,eOb_WQ=\P@W\8CUB1AHK;AVWSWg_Zc;6V>TQED=^SDbBa]b
.+LW8VC.)WSSK(+AT\P?\QJe>D8e01J^&Q>J@9&,,P?Y,77VD\+&QVf=;=HL1E>?
)b@;SX.)&F8C(U59T]5EE&d,Y64;7c3Sa>dMM[@_bF(Z1KNEHe65Qe1af.ZKY_IE
),EB(R=,EaH):&^/UOAQeJ<H?#O#\3&:@K;>_5,EZO?.M1OZX+:HV<dOeeaG(;>B
#K3P<MOOIf?XI>988NfA_Fc@>.7:9(Z&XV_TZJ>&(99])g6:]\cY3HZg8F(Y;,QE
&+E8M9PdF)&F+6)0-YJg1PJ->?6AT70bAGJ3BebR@A:[_c\=C,-9CQgf)MF3VZNH
+5M,[bf=+0<<?e2CYC?IS@<+cMCfXB[0\6,K\DJDMYCg#JN4?P;>I#01/_<JV4QW
;7HC#0_U1a)+WA,XUNY-(TcZ3;TZX\gE<d)5VM1dQ=\K;_cK/8[E=R<-d]TR4YN=
5a\83Jc20)C6&6^EQ-K?/N3-)CQH:]ba7LE+D9#G[/P+WB41BLg)?7:OD;R+61QZ
20-4?eS<d/e6RNJd2#5.9Z2G)R<MUI4ac>^e3EaCUFPT;>9^L9^(c&#5DX1UIg&a
?a880:S9KC)/9L9W<YV4[F<IZVFHXYW\Q\J#8X2C6/K:Y1XQP\-F^_35e;/XbHQ[
.>.]]-,3U9MM>d4E/G=M;KRJXZM^1>83bM8CWb&_NbQ=W\.D(ZgCagW:26KC:X2Q
)Y30g(BF?BB]_CXS.HOH\H.Hd&?(.].=aG[LRWf4[6A4XDc6E\>?PO591&H<H^g+
\XX-Z?Bd<TB4IGdK3M:2@(-97=;(YfUYS7088RAK:UTJZ]g6DZ370Z\Ibb+)g1]C
,Z[CZ-)6\GD48D;]8&\EP]+6DKOLe=[MW6e38GAMB#)E)YK_PNO.TfX2:.AY5M56
Ua^;#P_LHW&7g8/B<g)9a:])RE-5R_B),f<N.ccJc<:?VPE.Z(/PX@85bYYHQ6ZD
>3Z\WM9;C:QLT1IN@\:V/FF9(,RXQ8JNgDK+A(d[6)<9KK3Sf9MI@7f@]:a,e^5B
MfP/^]A=ZD6(9S&^b&dHP@]K=[AIE7.:e(6A8Pc@(N_Y:YR?)9LA^Q<,1+=W0BU>
0,7QK](-K-&aE9:IR.B?#\4<&#U)LRS-\5<2]]^K_KM]I]D^BG9&aS+RWY0Q=9\F
CJ3a=NYZYRSV]ZH6KZ_3T9,>SNPO_3U(:+dNB(LQWb@YFB+V)38[OXG9Fd81M;XZ
V.WgUNDWH;D0(X6L+33cB\.(5<b&86d1^PWKPf\J2Q,4,g6A#XG<E2,Gg8JBXc;V
WeCZKaU?D3d^XN56:3@,NO^48bS5FER,,bZd-6.=&J\JFWYfDNT3M)ZVYQLdE3X?
O=a2GKP<IKd,F;./MUV,ORGcG+/JZ\>W&0Z[#7KJ:eD7L@a3]U&:R7W=CJ=XEE_@
[HH(&M55eXR):FYbF5:XSB0e2<-YFZ1N\B\?<^f<He,;N.PV9=,71@=I2,a_9O,K
N++/,KJ=?JD-;V3ODEO6YO[N+TG&a9.+>dcR.[\:LD&bLgHc^)N(BF[bPU/b;+G=
PXB5e87&bQa]31FP_S\Z8U:S&E1:?#fLK)IZ7Sd40>?AJXK=dOQMESE)3Z#UHP)G
I,U-14)?F\\0YP_(D7^.8AB[P3XM3I;4P^/2DdL2dNMeL]2()W1>_Z<7-E,_=XEO
1XAF?beYK5/]=UZ&@JX9gGKc4PMTRE_P.4TOD&(_AD6Y>&FeD802+/@S+M>5HcFG
eD]31NcKZMfD146QZK8d^c.QP#f3UQ.Ea(;,YUXO^1IW@T&X##8,#YT7a1Z=6>H5
WX3a5?#I&#LC9)F3/K>)[QSBZ\+3[-Y#dL-Fg=33NTT\+[g&3Ug9H==WQY(IK/,:
\9Te<92Fb0QZBG\)(?H61:V5^eDM1G-1MdU>NY=L=_,ad)>/1J[RNZf6EP/Re/\8
,5^N^_fQWe0RTEfJc[A5<dY\V8P&E(OcX?Q52,&?cMDI##_8d6fE^ZcYKH#.JcV<
=B2F7IQe@d01.)b=f\Q=C2^[Ab\_,_R.(F9&9XDd-2,UCU\ZV2HD31cKVT5:0W,a
d&9@Tg(;Z<X#/;ZEH53F+De::IBGQabVH)2VCd;FX=aA?K1/-72CW=?-=G8^Uadf
1[Y9>UM3g6,Lg,d;Ac:ZZS8[Wb^GddO9.B\H5[=+L/c+R&RM1H&NFCXIK[cNFDH&
8D7AZVPI0c_<+-T>_<4KbOI=:HgAMZT+aTdf(FUXVb-e\f#^0+XG=H_LD&K0>+<a
<)a:Q79P3&-K,&5WQA&,d([]5dbHa2WNRJ_<-\R##3.];/gO4f3ZdZAT,HXS\e,d
#M9DPE)f5NeBc>aF.A:_>He@0[:Y2_)0PXH7+ZN_7ERc^a=[&C/7a&B@Z_&P^PZ8
D(@aXINXBM=3>C2^@61(.\eIZQ1XZ=@VdENOG0V?Va?gPZ:Zd.(b5<S.80I8(?6W
b^e(PcL>U2<=9<T3(Q7.1;W&._>/6,,[bfF@IA-V-X>>a8X\P7:OMC>JY=NYecFf
gH)L@A86S09^N53UD@[d)++R2Mg1)H89b&#fW@J?V]=UH\@C_?O964[g)Y3bKR9?
e,+EG4c,b3V)-\JEBX]DRFGH#=f1JId3^@&ZDag@=(d[\;8F&ZZ#<Y>3;U#]+/:I
0MJT9U>a)2WCCL#\?8+UCJ.5XO@T85[bFN8EYL;BX7=J>IUF=X#\0CKEWU7)W4_>
^P@3Hb]?)?NIc_+cf3S?dK<T5F_(-BN4,C;AB^ODG-(^+S[S(Z[&AZNEa<13bB-Q
,?.R.B]T3P;d^^^3Xb8HJ=\dfP0/Y;LU6;TOX]KOR8;CRH=VV+c,CbOGLcf\ccV.
,,.MU:457_fQGLP#A-M=I+DUJ<dZZX.KOH(/,a=2_ZS5X1THDG>22&04P-aBFEI&
\WXS_b2KQWPaP<TGd/\8+/LGY4RfGcJ@<V4/VFUL&dO&>^92^A[fLV=SS0[#YEEC
M?c,a[T77=TGRfS-GG5?Y-7Kg9MND,dbNL==B-\+&CT)K9U:,;S,Y/VDU#\.0F7/
RSd-..S3c?AKAN(7Q:gWEC\A3GK#O^,8CYCbKa@E/V9LXcVTO)/B5c)P&.&,Yd\P
(Z^#9(4SV,Z?>KK;DTfOgce3?(]7?-?8g_71TT]^QLH#U?:31(:L3.<KQ@V,[g0Q
ZQW&OOQB?E:)#JQg_BY?@0FZW2W0gO3,+BCF-K0E@T&3H-VcK4-TXfC&5V_QX@@[
Bd^g^VK5QXKO/,H3D/9V&A6<]E\[G(;W[H\FG?BEV9-[Y0B&>QK@cf[UFK@>.>(=
4.9+fR4736UGg9V)+6_O8Y2QdK]DK@&0N(^@-&VO,Y0>-3YVgU-)\//9ICV47VLC
_R&/H-/OLPHQ/OaC3S[BE#9J-RXJ.e7eYR\EJF2&g32XZAG<PL\RZ&N+):KY0#AD
cSO=WZVE?=-PBE=EW51EV\RSZ6XbCM8#XM[Z.=@QSETORdNCf[8#cUYX?#Jcf>^O
JU;\&/Z-D[Y8>5;?U[H=C^>7G_c9Q](9J2BH:2[fL+U;NMdeU@]WcQ,U9ZV^d,^(
#V<UNe,3]VR@;]YL+;OR>GPaWc)(_/IdJB.UbSU&-cSAU/4PLLKK<43U6a]7a<PA
PUGKAW-^5D\O/_(H3eI#aHDU(O3XF/_X2P&IcdF_G)>+ag;(BbSPgYe@,4&V:O^-
:5^?[.,^+7Q.BaQ_C_=Y@,XR>a6=e8;@Z[>/GC8f-fD8[P@9^Z26Od04Uf2T8cX=
7a_[dEdgf,:FAAQIKM(DT3Mf4a^>835.J5_G4Vf+3_:[=JV&T&0,e)^MEd@(e2U6
,I1]O>8;1=FD3ERE/fP]XBVGVaDaR=9,0e)f^VAJ5/UA]N^5.;;\DHI5^M2Z?];.
WWKfL#-0[&SOFWRG1f1[M+H]XbEBfgN_YZMWE<[015eME:gSN-NBb2_AW+_-L8V4
_-HbR(Hc.]0#cTQCABP^3R36,F\[H1M-4VSU@MP:?QCOg^C]F.(K_6IFaaTJbNJe
6@>Ue=L8(bfJ)d+>KM-JT.&_YaEMZBT.N5_HW<Z1\/#fbffd.T]OAB]+L.b&@96@
-4,^(>YVC+6<D>a,7(3Sd[_L#)\(a=ZPP28eW\?EEgPD^]0P<8RZYW>@5N14P>\E
:QNV?C<CZ9b@CcARNG_d\.F(M)-_=,>B-(V>A,,Q7/,/8,gaY@5Af:f>J\1]FXXW
LfD0:)f(DBcSEN&^WFcTaAP(5acI7_]:(MH_]_gBNb..KOc29]9bSG(?d:&-_>_2
_+&Sd2O.Cg\YWXN4M>?Q,Wc,Ud\GW.dY8B[Z)CcS5W<S)0AR?=R\TH/5C-=?9-#4
@f9D+dFB@^5Z=Yc<W;AXdHd^7)=Y#O/6R9;f@fWLSWMg.35<X6]P:),\LXe=W,<5
>_0KTYLaC7(R\_bFCK)=]HbPe?CD)P]-V&\K@Od3#WCF5B-6&K6_2QJOe]HJAWB&
6ZEOP]:]F65,UCf&BD=TBI;X2XgA8\=;,&_A=>+;3KV,5MO_?@4VY+E[?,.GNU&a
:MIE;5FDL0E[D;UBCF0]MOWb:B[UaGVF&\N@eV@1\HcWU883&dfH=e6D^.).ZO50
=R:e/dXB^6AZGCX]TUGU4/)5)cA?,4VD4#dfOb+J>W0G_3BLQ:]^S5R[<:0dRLXY
H:)c=3Yd&>:0XDAee7@?X(@56B7I?fUC/f.(db(5bL0YBNAXUM_Q<)1Agdfe>JP+
?gA_JD5C&7+R))bMWTX3L><35LfQ_93Vd\#f+(=H5Y9D3Nc@b)[NP8e0cZ^[Uga,
(IJU3PCO\B=bAF^>GI6Oa7MMI[b0]gF7T2.3PeR7_SRePTSDUGI)NP9F/GZd^FVJ
#9BY#DM5:82gQ<0BQJK=<,4;@d/C-V&[&8;,@V(Se)A_c_4EI,VUI_H]O6^?dbf[
1e__2C>#7]A3KbCMEV16d-\aT?1eW]7LZUBT?3&G(.g:=Q_O#5g-O\=-O:U,5=@E
.B)T/bXGZWV098894RLUf&,EUb(&-=Y:XF.QD-?^Pd>&Q@=1(LBOXJW3X:GQDdEK
9;-J&S/R<2f>()@40RD6GM^FH;.&>TPcE(dN25-I/Sdf3QFd)^VT0<C5ePL1L7Jf
D0?F#WXQ^R(\VLgNeSaS-YD<,=&@71)0ER^7\GXB_e1<M3#@9VS])(CFE7f>NC(e
GN:?A>U\e>=[-KC0fCNfc>=,@OPGWSfc<F4QbB5N?G8U+^_METf)TW<-FZQg<Q;R
E#<;@dgLMB+:b2I8)(X4N+FM7fIc0@S0(Q+:.@34]gD<8>a?eF1I&NBHIJM9890,
CbOB8)BaG)=#Ab&b@Uf@K>&gg]TM=#=J<>X5Xe<8^KQMH3:>)7YL:M.3QU)8GNY(
3./5JDF3,EMA9L/\gU.cGI72N\XSLJb>+)BV7D)[NIA/3WZf13FBMB__@5X4H1HD
81XWOG7(L<).ENQ:OS5^6g9Z?XNIX_;GLK=MbK&,gD;Xa+4g0P]_[0K\5^NGQL;L
TXOdA<;F+HdDZfK3gK<#68TeH=JdU1J9eP^8Df(YEOg/E2V&b9.2<B=&#NRXZVA;
W)<@UGIZUWS;dJC_]QT&FXXGF=>d,=NQR;:f;^3+7-H#]IDI<7BY]3YEU>>D\Z5Q
(I1AIgE_)3,ee^@R,31:7S9TB(b2YC=(Z<3Z-@..#WL17Z?=T^J+]C.:\PBe+5[F
I;1,H)&O6CH3Q_V7aKW+AI4^P8&.^\L(L9]>:D_\f?Q@eLH^2A_#E6D^99EYABN>
9?OdD37Y3YG^6IIQ6>gN83U4VD0&U,506TdFHRZ>D,B0\,VO_MM/BLU/?GJZd&,:
[1&TUbU=9KBZ-8;#WM;0]+Y3L7bca_;gaV@(WT0PDbI4II#+f;f&aSLA)5P>ZY@D
_+a[=I3a=S8>GOMK\_YIE+Vc:-bRV6?)OX0,8P;-A6OcD<EA3BX(Ge=W5=U#KT>2
-V@cF6H@7S+N.=E=1\cA&XeZd1S3HHZ&4;c=^@1&ZL9^=:FI4CG4g6B6Q-<)6fO+
be/D.E5RO]E=N99D0U<T_4ge1UNVYg9>MV6=[SGR5(g(c=J::f-bTKA2dfLKWgX(
\@?4(E.LeaZ8]VSBOB0GQC]Y6dQ,V@#6H>PHAO@ZMSP7=b=e#eVZ@XKTJBPX)Q\9
_N^<<dTg5bZ>D7f8FUCN1TG1Q\@.5E.@XU6OEeg[J,R+9/2F;+)LD:@cN1IHgVae
ZD+=4KG?^2.-C7XCHeX_40gKXc:@b]_GN_b]/Z.d]6bJ&eWF5>FXV_^3bEgS@2#T
Q+<bZ7I5LX(,@8WN1QL_0Qb.,PQ[[N+cFCFU@g<G@BU8^)QRH(/+JDN+?EZ-_MG#
Bff_5(^4UASO1Kd@_+d+M(Ua83_8K)&2A?4.T-P,Xe(M&1&U)ObPE;&079cNZ5+H
NaH#dNLaFe-97IJ&ZAZ@IV066=&F]>2dHEGWVLP_5N.L(5bRJab?==H<)(DQ0eE-
=1G.5c7II#@[UNTI^\+X#?#)&OY-XW99aUX8)PYL)Z:^P=BQS0\IF9Y3aM-MSOG#
<U5e(KA(X:PVV[H[09;AA+D)NRV29X3DDLVI(CQ&V8A)_)#Q=JT;BRA]^&+U](,6
aP;U2c\]O]ad,U&cb_K3HMDP]_:d\C=V8WgLYZBQEe\T>+#5H(&^DfI4UF,:JO:T
VeZ=VELO6CX9:.f?If3N.UU@CaHf#4,e/DF1&b)H9;S=)5RLdg_cYS)3[#6+dRfb
FJ<.e]Y^ZT;F9TYT/[_6OW;8/e+Y<O&6Kc&,-W#DRHV6?ZF5B5U[1_:I[-;d.a#L
W&\UC[d53]-0K]I]VVP@d+,dc_J<N,BBBVYbVBfJ\V&?6R)&BC&e&Q;OAgL7OPXa
.;4ZU\6fOfUMP7aSX0-6SAIN[-7GQSW)DQR@/<eR9A]J/2V5I:_G1L^9<>C18,/^
f[=(C^005T)a=)6a<(QIUbU;18a\&:?<(&NP<fL:Q7H@dg_&[6ZHN:9)EZ9EIW^(
.P-SA<QK1C\F?)(#Kc0OZ8.dY+30:-/LdDOF^AO=.JU<X[W=[&=Y<>)H<B[U046O
(FT41QHS1=)OH&>=S[]>RF6;2^#S3(K9YLff(/c?3P=.W41Z-dBLK@Rc,T?fUQ\3
M7/284#SCPYFL,\Ed6QA.3Bg^7X8H+LLQX>-XOBQfKO6;_0d98+FdCY<UCdIJMKE
&eZ#L:ga40UBfOIU[9X&1AQgaRf1J>SJ&-Fcd_UU]LRM/=2+53d.LbR8;]2D(+BF
RcWc6a@fL-(O--P3Dd,_PL:e.__;B?MD8H10/2aR<FMB#9,3@A_B9HA]RI,>\BNB
2R4?+QDdK#NSP<4G&IXSGHF2N2JgRBA1fK?_2bReC=7e<6S;M=,]4NfFP(V+U<E+
TI);2,SQ?ME2^F.faWE0K]B]S[)7^1]P9UHSe/I>#Z4/7:CU3#FVT[B,6<;[\:VR
Nb@^,4f0F9QgJV2F^cJ<_9eYS/]ST9,0_=T_6^;Y&-^CaQP^K\G=^MK?LEJAC?9_
;7+VJQDB&GZ-S5M]KfQ.SU/,.U@&S>.C#bMgfJa^]SFDB>gHZS\7+cL-M5<#fO_9
VB:_d(c<2R)S1]9b:QD5##YO?:SMCVF&M:#VGY,=^<;_85H,W0&<S5K(d\1>g?NN
I8Y..K8?bE:YJ(C7;?6@Mg3^[8#]X<9TFKHQ=egU:Rd3X=-[.RSQ,d9]eCI(K/@.
/3-5?(Xa^T@(7.UOJ<Mc3W[_2N8,KEOC&Z#S<I7O//]JgV^)XJ-MJAZDXX-^-BaC
^7J9XSfK.EQe1G.R(S)<SRf-M)8?6B[],JQ?X6COTB8fbJJKKZC-6/;4c;9H(MVQ
2GaS[g)XLe_RVUF7KX7-NbGJT.5/.]c#<O6RE/#X4:?<B#JaM82NR7QPfBfB=6Y-
_,@c88Z0d&R?.KQ<<=dF&UR[XeaaaU&Z4OR)58F=L)7/S^Y.,[Hb7Y2._fG2VU3,
:VHZIaPB/^XH&#1_LbP>YJ.>RA&G6I5Z0eMZH@>(:U(C,?H->1J9]a7e/DB=McH#
H7>C8e\IA[O:b4Ucd,9NVD1BWZM60PME29e.)]9N\\&@LTE6;_\)Kge_eB@;fKAW
(6\K/ZW<c3_7(HH6&S/&#eA\M@cVdM2Q3Ca62N2(.3D49eN>Y,[(;V<;,\fQ@_,E
fbOXc48QKe6L9;;<QG/7PL@8=e4EBg-GCab+U_g0>V[Df>eFNR(He@S[/KPO=P+R
8a4g3(H8>V/LCZ<UNf(cO&<@=2Z+.U1&LV9A0Fg/[##=VXH]7V6K;a:&GccG+>9U
U7M4e,OT,+#Mg;2e1Jd3bZ+5F4/^M)@gC)Jb0CO5W21bO3gJIFN>/#VUM3.2L7,?
374N+LZ)(7.3\3Q9XL\)HgY+;WZ>_^4L9C<[AJfQ-0dEOUYDW:&OKWfF=SW2Q&[<
Y(+8dSTN<H/Pc80D_:R(??1^SfPEDIV>NZ>S)9G(#.[1Le.2P3SR>/14H<TgIa@+
g(<\?[IGP9XI1N>be)HWI9+D1VJYSf]4>Q8?@S,;239WMY^c<G8_[c95[g.+AL=e
7)B#CG>]FVg1F(bdd;FS(&0:;Rf1OG)S^S\YZcF.).c#<fYRY[F1D&5/?TLd:X(d
Rg;5.LRQ=e.bHHL;9O]-,H:e(R:;aEg=VC=\+50()/N2-\#GO\E#Z;^22+&N[P;a
9KW?2#S3H:VR?0O^1(OFFE=d4Q77Y063R1RcK&6X@3QIB+S+C939YXaa(UM?YL?c
WDKI,4)S0c-(Y&)?;V77g>ZCbW5/:[0_)&I>R3bfU/@\#<VVMOG8M^G_M<Zc5+MD
Za.3Bc^df5U7bE/V3E5QB]7WDb>aGNOO=LJ1H)(Ae.@Be<2c-[ZXeBW<<GYN0HJ#
IVR2IJ?WTYY7C;cGV7BM:]<aO=,0K)B9^KUeM^&A+&A=X&CIN3IU&I+bB^g9,cCB
[+/<6(P]O4,U_:JTE[T,8,K##K=7=0G:?W_Nd2[NU&bWV68JOATR&b:MX><KPA_N
QQR;;I:1\\Jc1,6);40gQDC#>_@ZOIUD:([P[IIcL#(HWfRQ;8]G+=P6fY.2W5U:
X&ZNa45agdH#aWTKGR@D#HQD)IM?5+U7HQQb^W.,^/a7Yd>c<CSTZ=b8GB>#LNLH
7QTcF=R.TSeY9[_L[Ob^(A-SbR2D&Z/b]KFU/&\LM\EgQMW+(J(/CJC9L=Geg4K<
8Z,W5A1bULPY\a,e1d6]a,G67gA,C62b)/gNR=QOS>?N>W:7PYJ4d((7Oc3db3eE
#IbX\IGeC&eSe4e+P9J\B<2E8G_eY+N?#O2M30>LcB>VeB+^1LSY2],8E,bcN/9R
8J:I6JP-KFcWTb.gGZ29?5<JL[F@3+&/VQ?^U59;G]&SLAB<==\FOIg^a=\+Kg1>
P3M][[B/dYf;SE\>^N;<75UUJ1L9_N=KU9]J&8,0&@PJHa?_VYXG\A4cK-T^W[TK
JNfEF(L6,/,cG]-gU&,:-VgSHBbF[>WY]6b7TYMP>#^/YD(HfONZZ;,d6\&75@WS
F0BU;L)KeJf;EOC_\6VX?=f[MgIcD\Q3b>#92X3.SJdZ5X@>H]^e2RW&I=e<HGS=
)dgf2Sd+0,gMd^NHJWIGSC&K1<CGH]=8(KGE[S#fL=8eRS^YH4JgP<J9ZY9J[I+:
[6M>84e3:J.C#Y[K5N9A-dNc72364-8\+/T4CRb7^/ZSc)A-#F^).T5&@:_b^4.S
Z@311ee[ZZ3QecT6=fXSV#G=LQLca(QcJ&KV5[D2811Ad?c)ZHM6AU?c_).:JF4@
<Y0G4:JIeWX4M#eG_[]:4H,[+U@^A)(ZY=H8C#=-S)TcN(3V^Ef)N?>MeP4AWKK,
,9C(^/fG=R3JCfE4MH/c:/,G&HLQa?8S]>B:8^P/#JKEZ)\U=a/+4d+T^+C1WM[N
)WI];ZAJS8@<6K#\A._G6B#)0E\/eBQLPDYH<].G^8,CRKC1)A:CH?,,\3]R@SE1
c=?:8J=J8L2A[A>02JXW8?D3)<e=D=NNTRe/R2>,@/+,4ERAH),D+(APV+Pc1cJE
.d@SL&8_</.OL0#:WX^J^;(gD^g76V:]Ec>2878A#1TbT.L/TAa28LC>c>?#O=Zc
Y<TRRD=I>1F-_ZD2NYPID^?G9/X_XM/L,fK/K.LX;L:JYFe/\b<ZKggf0R)WK4bT
Ng503fQ,Aa:ADJ])/TYRQN-AU[cBg08_^5\DLH&KH6T^U\=d@,2V9^YKWKZ@b9Y_
;4a8[D\D<<6TABXTI-GgHM0OMW)B]IW)^EKdP65cQ0SQJ)7M1_K-#VA:9;W4,)//
6=.DMRRD8>a-4KTc(2<SRU>L85Md7ZR;RC9C<dgK?H/TST&AZNY.1M[_R89B?ZHU
/g6cYKA+M)1.aRE)SgR\AfP--A&@GdZS[:H06I<#F,0gL_&g:e2.25NR5]\#P.[M
e)#L,,J8HdM//WGV#3CLFabXf9JI7H&W,O36=\_-Q]BF=8Od7V:-J_?3F(MVDIaf
O]X-Q+>\B6_BQSVDb&@>;;H)\394.YPA)+Oa,IM39fIJ\Yb<S<OAD6Q@BaCXXD0(
?8-QT??0=UC7G]PZ?E?a@,L)GBRA2S,3.C[)_b]?SA#b<)B,L?R)#[+X5Gc+I(A@
d;S>817.3<UZEgI=)5fe#1+R7-M6GKGPZAIA:^AAB5;gMV;JA8.KLA-X6eSBe9Y#
JOgT)ELd]?MBU](\UH6bU39NHU[_>N:;Q<BCV?J;<)a0Ad9EfL&>V0GU43NJ;:-9
HIeO(]5#1A?56b.H71_/#C&aX[:J@1NBX&QKEc;//=9JZFHbU>@:.]bf0?<907WA
/b5e0C.T<.)dXLL<9IR2PJJPMS#gcd8>d23MFCaD#N^.Zg60aA;]HAc<gAIS_aPD
_X3<cM4B2b5&fM65/6=F1/)[N4/RZ^..?C+F56F=V[/dS)1P;b?R6\S\>b]<0(>-
XS^(H(c;ZaXaKKGb4)Og;@IMB)77;J[^-MYSD?0:=GHV2OHO\4Re^D=U:Hf=T9>f
_ABB1)G>ZNAa7^G@@d&]Z@SXaD>cM[QWT<^&DbdRJeE9T,2gM3@D(YPPVf:==2eZ
SPO0F.-@(I0@,?U/5Q]/=8IWDXD3eG6RRf6.[c?[=AgZeI.@<;VEN4e]8<A/eFB&
T&[fe<(H\Lfb#^cbWN6(OgaB#<MK-+[fR\PK8F0Ic+b&3&\W]aeRX6;^bY2.(1^L
3<LH6NfP:#&/d5C+3AeN<G1a4?;4C&]J2dC=ZTIF8\++=+<W-0I+#f1e:3HgB1/&
WQafNB[<,TX^e.[Q1GA#dXIV&^-f8U=HM9gROa\g4g;aGXJ)(8JB2WIX^56R#\7<
DDe?^8J&SR/TABY_g_>gFA=d50e?M()250M/fQ5\Lb]5f=&)fD5)T=L1_)V;+Y46
^3U1OUeP<.E;e,8(,J#G?9<SG-e)C?FQ:8#1Y:Y[],4Tb=IeQ\]-X6TX:@+#QeN3
\gWVH5.<\?U&O.^RPFB[#_^ccL21PMS2YY=#R5T2?,?5Ae:-X.WK-LfOB),;147<
U5:aWDbeI.Fe0T;=(JH;Qd&N(=DKN-GO>YX<P<7&bLA,QO8?I.dLF^BG\-],)U7\
0;b=26RCGRQU\N.10XGLG#fe-C4W,/#H3_2>-4#UX2dbD<U6XH/C.fL^1S,.QTR;
B)(9b]:=VFDcG&ECa-P:-=^#c7_/&LgW,Z)[:2f9.dMHD=&H(B\L40JPa+gSH>YV
)C@>:C@<_HH5a>+@ZOXff8\e8(0<=RY>ST;7#:Z,\dLIY892HWL4&aXO(GN>-::B
HCGQQGg>)RG02+H)C,6=?6TP6KQ2N\K]LV;(THSdK@]\..+Va:<bag&JY+#+#.F/
39Q)aT8XREV7CdAG7[YdQT<eA<[aE0F7-=]I)[B=()&G^Y_Q_:<J]@(L&@35aQ7R
;NK(FB_PGT@Mg#cPO@=MMJ#Ia>X)P=2EFI]BW6H;7ZQA?G87\T+OFJ9-Q3BE5Udg
Zd._fB7gEO?A;ccg8J^M^GZ.DY6L+,TB>&gL_\FR=Ga8?d@&/BWBJ,G2G;?RTYZ/
J1;S37383f3OYIJa5W[U6C:0?@OQ#RM6F;<B6E>I)IN)UKJP(ef/5F3W>F:M[(5b
>=I6]B_7cT3@9gZJ-S@gES[H.J/LQd<]<HK=ZYffL9dXgd7\[g>=^[E4R-6ZA\Q7
]3H(3V0c_/\6IdVSP9M;b-=4<(b@.#@\9ER23L+&8PWA;?,@g\(G)-53]@=E\@D4
aZ#:.XZ.(QO5I5ab)c4]/f5:&SUW<?DA]LcfL&bFXDXd0UaG0AEN2P4IYf2^DU.T
K:PBEK=#dWJRUK+3bVJV.OG+HCK.NYAaAQ=EY2-/XS.(]Z>;IL411@^L(;@JJ7b]
0WFd[T^eGR9)Lae^g<1e10fFE0aG.H:#Aa\UZQ3;VMXg3fKL/NGS_,YO4XCP.Yg[
CJEJR1>4-0;Z6+]=B=?0L/>\g#@(C=:Z-KPcd(&=eK0c/F,FE2>\WEd853VV_7RE
90YEY.0<ge].a\:^Qf-YJGEQ_??92f\UV8,L7R6^ZD&L:14LJLZ;aQI_C._89;3L
7Md@QJ#(gY;1)AKZ]CJgBJb+&6/G58]7:1eRC2@W1/f6f^[;BC=ND]MNG#8Y+9RN
f_A6@1[]X+\b,/F+RIb]4Q.[7Q7bJgbcKPd762Y+O?P#,D;O7-aQDAWNO&U_)F[b
:(:NI)Y66(ge(=UNMG<)9ZW>5&A01eC#.H7be9KYL5^/=L5H?:SRc6f:eeXL:Ld<
KLXbIg6@YJ0YU1a8#^RY1>=8P>&2IS2,L/;N4WY?+JA(9T.)C)b-^OT5R\\N+6];
S9=?1ZSPHZO2]_)F3ecRN<_A9fD+EM#VCc5@,Yb9)DNQ)g+Sc10MSae#B^>cF2gH
7e,I&;(,<a@7L:HI6/9cA_c9Y#MA.K=N-8gVcIc#DT34g+d4V25?R/3bHZ9O<[1f
CTCT5cK;QAAQY5gU3K3B&YBOeVa5>7XLYI)R+YA1KX2B;VPBWVJD]FeO<P]?\a3@
5b(]USD/A4@AFUcN1,\?NMT&SHe::8N<d49LW6QTd25K>O&b8.?0Ig2,aS75;-ES
4(V6HDe78.E5S+XWcZKcQ1AD1g]edDE6]2g\12^EPWD&gJ8@DZSEJRQMAG2TN7D2
<)SIePXI]/\P+Ma+_bLbF[(ZeIYX[d>Yc6P1K=I-NDI-_\fa>[EG2:fUBaGP?(ee
2HgbPPK/>Q+BF@L>Z8Y;@^,[6&PKb;6[5LRV?FZd0EZ13Qa?IC(&.IcXK<PP<1HT
QZD2Y@Rfb@^gH:2])]>d<eUd-_M51VBcDagd,<G(ZO_UEBbJ=]Le55JA7D(a@L-#
-+CEOK>CW#@H?F77dW&c7eBU4gE02L#6cM[^,M02,QW4O;#54e8-C2Ec8E\5L1L;
9K.MgJP=;CKgMIK.@NUQQBSJ_V&SGbQf8d:.;=Vb/RB?_ZNHQ]FW#Z<.=?Y4NK]<
_+(0+U[K59=#.P\0NZSX;JfS<ZcLMKe@WacePP@AMAe.()TJF#b=^K_7SdgNDELf
)>:?d&aP:3F]KEQMEQY##T)\(RYZ/EX=_M5@Qd/:;;@?0\3Da_=?2U7[Qded@;R&
+b7F:(Hb#8+MVLD9V(_YG^dH8>VYb&XD2L=4.(/DY\G3b65GEd#82VEEQWV2YMMd
W-RWT=>]UE0S6>WCJAJ_E(b:Og]SS1a5GI)PA?./F^,6H.&13C_?\c>ZXV:>P:^I
^0GIHe0@>UY8eG]MU3UP/(R<LWgVXb6E+&YR&C=5@eC;9P9-d5_ZLd5CdZ49a6T_
c:^6T)30L71_cbbZ1>e0I3aU=4eDT94N;B?S6a>N2E91&47D5A4I@L_@Jc@BY&[^
S]5ad(G::=3&R5;QFL&BH7^>aDPfW,c51712<#E-#;PQTSbTg@a\6(0U/Zcd2Qd3
QQf11A\e]f_8f#U/7.@XDD#O1D76<1gHKNJQ>7+^IX\)T1UIT-[KMGF--bV(:]YG
6:+cf9J:dC\RO0<FB94Re_+/0_A.X<M4Y@)[\9A>+R=85<)aQ)F0,J9;=Hd^gS40
)Q<3QIfTMS&::22g-\(5g&NZ;;\4J)>NNL&=K2(9K=b.ZU3+(4)@#]70^@3KaAIR
(U&Ff,9U<C^6&4TdYO3b^H+c7A&2eT9[3]gL0N^b2R&b^)>?HeJL4g5C\4EGXKaE
3M=OcOe^B)+&P6(K+QPWV=H9>/7NOUOH@^/ZU41bXd5c_I<L0ERd#-&LH,0(D#@=
E=IZKc=65)TTa?&Ya;<LE+OD]B^,UI;,b03:ZdB4.]AFQ/)>Yb_-G@K(EDa;eMF5
]eKC,=W8D>]4fXAYPH>IbQL=0>g_-7M?Y=,@2UU2:1-]D012I3:gU,WN[YfBK63W
:@C-aL(8g(UPVQMV-NAT0-#(RY#aLS<T^ZR8g2>O[23PC;+)\Vc@d[2A-cAS+8&-
IK7PYA=Q1QBYaIBYS31J8=7Q-<_BXJF,^==O].&-HXHUe?1?U5.#O3ML==E@NMQ^
C4dP/fS?4@X6adCWD#:<NQWY:dCSG^,51G@5&?<dX;3S:eU[3];4@P1f@.GHg4YF
7<JN,@RRbfTP&ICN2a]2473d,COX^/6A680_)T49KD@(_U(;f9@9SNb/0gFC)X1:
EH7P]<bF,MFCG73,#f(3I>=EWW0.N_Z>A1a-R9743P?_UKN@g(AbH_1AQT06VE.R
Bg=93E_[;-#NW^R8UE59^S5-aeaH,dIY(DbFf1?#;5@gV4I_YAd=PU#J94=G6C@R
_4<&T:.+aYE)RN]^2d8<\NP5MS_ROF2#U)+\-OMU.<^2D;HBUd>VT\]E9+H2.8#c
6;DMU)Y-4)0@PH^OV.,B6WZdg)6MDd73+Y-24TTR^<:UM_M-.(:Q@.F/;KY[4@-Q
O_Gd0DBPKX)6VX2N1A1g-X<0[=>\)fPgdQOR0DJNU.)=5#/bc1\e<X;+SWNb?P?3
E7b4XKMEI[ZN74I:[4AJ6SFC:A_/ORAJL#U>O6bCRJ&LDAB&,J[D0DW\VNQP-FZQ
U#2ReJEF4XXR+OR,Q;a,9.KNA<?;HLL]C;4B?b_:e=Qg>3#d+9J6W2OEX\>FEBd7
P.0d4R2FK3AF\F+=RVLNR+&c[DN_d8@D4^TZ=.cU#9^Qc:E\54g:c&\@]Ef)<e>\
/>-YPT9)A/dM520Xe42HH4Y<9).2<H:AJWSKMD^AE\Md8OF];5YI+06QV-48^d-6
-[LZNMXVHWCCE6c=42RP68LG\B>e;;9XReGeG8Bc-aWgQc0P(G4-K.Ye_6]Ia=2[
/56Z>_=PC)&ScNaTN=;A.+4=Q/+-_Xc@2#Fg>(bMI^(K]9N:<G72DCMY.>ZY5_IK
/_,R;J1Q1e3-T??NLd\Nf3R6T6RB@TC_HI-d?K-)HT;<0/4^I7B>8/=5374JO25I
_fca06739]fS#.S#PG^VZO?=?-),C5CA73JD1.T+6-/QC4gEDe(d[TQ1GA+@a:L0
[.&+OYM&O^5aD_aa?3UEL&d\B#2FV6A?=R#91=90LGBZY@&MMbQ0<OdP.=5\c<gP
=Z+[5eOBU?ZE>2IC[QHIcLd)L_TM#CM=g)Q?VF_N8,\D(cY^H1DZ6HS2O<fgLI[(
eM0FdEM[B@L3\Y[3K2Lb=Rec),,_D^1?[F#N_HANEgK2Q2K=[U<E]Q.G_8Q>52=T
9d]#0d=\PS?V6L1(HD.?d=/]gL63@FRWccdPb.>6HJY3eF=@RZ>UT#=V6+#F[Q=+
XDV4ZA>D)_5U3)/]LeD1NbbfIT#P/J+W?RD,,OCec-3<-0+F5GC.7W=c8a:Q;(AR
=b^>W1b2)X]/DD;gU8.LC&dCS2;JLO5R-FJ=L4G8,G=V,<LK8C(9[Q?Q(@2+9N-b
8N.?Od;ZEPJ[(Z)4IMR#(L5>5;Gg3a>J09?GbZ[:E9e]):XZ35)]]GF?W:aDQ-.X
D?=)b-aF6U/K7.0FA_c,ZVb>[</IBG[Sd6N\7dNE3SV)Z]HRBOcHL3<,S#0A:b+=
4@AbFQVEcB<2=9V()X+6aCa54Ab&;R>W6(gL>23ZUVRC/S&bVG-2CZFM7cEOL5aR
8WZ;5cPHO:Zc)A8X5CXXY]B,1Z0C\PB;8)=eS5ZXPgYb#H?BF6KD=U]b6G3E4+5W
\N,APMUg^,We1;T,d&]2DSdC,UA^P&.RB(Y/cQ/J]g126RWLAf;716@4E/L-H]B2
39S[]5V5UMHJcG&g=-&/VfA5H9JJN:L@_,GSY4+0,8c32FN\I3HY)2^Ng#,,1&VC
Vg&C8L_,]GgRH41-N_bJXQg,f7eS.Qb079I77:>8Z2eS72WL+d\.[\2VENFKHU&e
FJ8d3^V_6-/B+1_C?7S]NLfCYf&C)YP,3HC8M2,&VOaSNQI8\WCSG6?GT_-233V.
dDYeC1/9.X-ARPVM,2MR(@T6<+fReG4_F^^fVV+_R@?SP6HZC>VCO4K:J&K)aT,I
0&Gf7<&2SL:7Ld4D&2\CEd+&^((])PU8Sa;8^^4TW0WJYaVHV,]3.S=-]X&dGgBg
=1,;fA14E=\c)Q?=_bSB[O4^(YaMWV49@G-9,0g<^<eB3M1dRK=T\WEPR&:g5?QT
LYaYHQ.aRMN-/UFAgPS@,5KO-U5-fA?PfX1&f&RfB^IPX.g0=ORURU<6[I>+dSMP
FL6#UQQ,(6fOdMXWH&N-(g-^DXNe]Q,[41N=YG;(0a&P9Lc9]D9c,C4OZ::9e/>V
J^4BMc6GGS)5>gF]g:EVePG_A3PVbFGg+)]MNM\#c;[ITg473Bg^+.fa=B>>5=KH
:PUN9\bV>0Hd+eV:LaLIff308bd#4=\+.;g>GHJ+W3]2&:0ZY>TQ4<W>+2]V@(dc
,0>520c\/\Q&R50ZFX^4G1Le54NgIdLOW=HDQ4L.\DFeBZ,WXgI13g;@EbQU6\aC
XB4C11eYP/6Y8f2?@<#N^N9cXC7XCAD7\J);cd]_,X(bcE@>]Q4=6<G5-f_-aEeU
Mcc9cOSO_RJ@FF)cd[?(EA2cOW_dHZOT?H:=]S9f6#e::gXA-g].M0JbA6R=C3Ac
\NZ]VcA^Y7Fc&:bRM.09g0@b<:Rc#Ng?D^a_dIB+(DfMK.7a3XbY@?U#78@W/Z^A
=,V#,cb3FL\Oa&&_9>9,d02S,B2?3\<I#@de_A/814V0\\5BOJ;XEA/H[&(2OUJ=
^B_-LI+ERd0=U71S,IL4>^#ba@HU_dM7=.>#\(QTPa9Z8cNKfJK=DCRBZGBd+8-)
AWH-JYK4R\T=G.0^fUPQDBB]&12cTee]W/^BT#[C-B)U-G#PA;/O18^HX((6I<,-
dG/0#3ed<c]J_N-^_L?9G((E75?4P:FZNPFQC)K1E9;OVFg00FSE9b?C6.PLY#g.
A6GfRX)\8MY&C&=MR(<\ZAJ/HF#eY616H1>EV9^C)13R>eEB(Z&,2E#5?M62DVVQ
/FEX0)U@OfeXU5ME?6b06[,B0.E4OII=#:A:=@.PIcd#._^J>#2;8YKE_,LYae7F
[XAD&(A5b(?C1CFAUEU0SKQeHV&F_<I@6?BFY6O+/;Y<H;K1^N8H>P:>-+D2ZV0G
&@_4#0=<RX_7U@A_>(adUI;Q4=\<.[8]bQORVPF9Z,]Sf=b=eEL5G+2A?B7ZT+d[
@>a/&a@a?()FR8c^Ra(.@TOIaBOf247;+0S.IM0-(=UKHPJM[S_2cQ>=M;2^?O)M
;IXIZ8g]WTW0U#BXTAJ;4I9E/MAU.3R6SKF66dS(eT7:1]3GB4dcET[;cOK0+g[,
9eH_c[WXL4V^69M:-:.E4M;9UJad190XC:g&6Z6SeT6b/3f[/\2]5Z)<W?=[a2Qd
-/MZ4BdB](SL9D8XA)/9GSI1W1YGH-Y_feH#BKL)83Y@U6#]Ib+_L8],G6@D^@e,
g+RdAg:#9>:gCP(.=8QO>P^)DKEf:.<3#^B]&bBd2e[S#@E\SDPdB1[]YNL4M4RC
I(IE;PE2eR=TEUT@eJ(&NA-QMCK^;Y]QGcaJDVMD=0DI5[LJ>dMBQf7H\M^e?8.#
4:f5RJ;F)3e,5H(4)AbS#ERaJO5IE:-Z+QZ4P13P+IYKW914VA<PA,/IEHD]^g/,
THA.dF1;Cd&4UW:ZW]&VYUd(]d_M\UaU?40:=e8C)&;5_g@,:4/Q;a[gKDc99:)N
;6#4<8X4_RT:DFA>Df4BbM:^YK/&FI[.L><.)](-@BO9_W)=U2E6(?J7dSdB.0.V
eP_-SXE+):Qc8N6[?E<O]4,OUc=@_dQ6<F8Uc?R)e.HBL@I^I>8284dJZ.P,U).+
:LNa^8Z<.&YH0/5(]M5>bU@+(C,/4Na08V-g3CWdCJ+:g,1B_eG.N\.Ob_^D;2.I
@54@eHX2.GOgS^732@V4/_U8]S^<>a,0g3VJ<Mfe=<d1]e=>?O<,./74.JE?_SW2
c]+7]f5bK71gX;XNL;X^RaM:M\I?O[JI<M<>OM:R,4RG_7I=8UbU[c?0=a+SJIfS
6V@gZ2IS0-9fLg#^BPKI<&W?<QG#3T=1QEVBDg#,/@XV^?3?UIa<MYF:@CWNfM\:
TYb;5432?S141C)?-Y=a_Sg@70PN,f@GMZ-A73g^d<US&0P,[2G)bH=LIQH^E=\=
WWQc/Z2aC_D\4YAK,LEcg;9f>+/aZO>]GbaJK=EUJX<=Q0>7bA+a;)AO^,]/^NK5
E?#(A>U&71+e3SbZQa7?&?;VN(LS@dbbA&Ge1g#T.^B9.=FaFg-\BfeaJ;J<U147
#5g<ZO#Z:bH@c2&91EEM_;J>)::@CQ<bVSG,U58I7eJOeBQH=VBSMO/<_fZ\-&_Q
V^\0TC<Q&GBU@JeTN/EJIBTK-P+6,J&86-^1VXD0(J<#&6=N#AOA3Y]5(=>6T37g
c6aCOL^P8XQR3bV?5F+@-3EbCM7I&760QN>9e=AfZX0W1RNaP,Q/[;2UG-,gHK6Y
cW3FK9/gX]TKZN)Yb^<9]<V3;gQ1H6U3VF^4D7_8g2RW+T@FFR-;af6>^S>W;/=Y
K>XHZ[;g.0RME?ZYLF3\QRR\HDbaIH-()#(ZZNL>E#V;BMX,)WJG9<)g^2/gGIcf
dGIc5EK5cMd+_.Wg;)gG9c\U/agOg-CPA9,;Z,]N^Rd8a[;7<(eS^EJ)Y/;.@g)U
_97f=6+9O>?EMZ7Y+OYKUVJ\H:MK-AAI-^]8425#U^bCPFO6/KGbb6O<g,(1\:DR
X3Y901[SI^gXKS2gE.-2W^UQ[]Ne5-dN\4UU=f?MJ/ZKX-[PUcNf/a>UA\XLAU\3
(c@,=A/L-9,UKg-MBCIW<@=Q>OX/VC9JT4#6&VO5R)d3ZabFfSF3V/VUM&UYQ&-3
=TFQ_\0)g4JBO^FZf3SG0R.(M0baIM@>/KNCJWKPcYTDU,/+QGC.<S6;LUUU/L3R
d5UAC?aZd5M&bT,@;_47F:VBGe7^1\/Qdd:BZAUUN6IfN.]^18^B#K)N3<R116/.
QR:OHK,Y-Y6G/eB[+>TbbQbfI&M18[Z09d/Td?&DL2VQ(5V##-W>bMR[\\SAZE5X
UJ;9IBG6KM#I\K(6eWZ>P7OOcdeB-DO?F?G[;.K24I.CUB04AKQ>Q-5B,Y8X1Y#^
53gTS.cd@Q;03(H^;T4:G8a,gUXPd;J78HP&d^BJE03>.6MeUQNM\VV)Kc_<Ae7:
Me<9AQ,&/;I_HT_,fQV,L<0H2FId41-XIa_Q;&;A5RHB=96VBI4_&5Z&=H28b66H
TJ38NcF50MY(g6IPJVbBMS#1KEE7YC7LKTR<_gN9_>_Y_U;bbL[,[/M74)?+63WM
?0M>f5B)3UK5@E]dJ-_.b_M[9AB@)ANAA)PHSdS):YZ:(U.c]B(2d@MV.DSg:+.X
5UYHTR=^^58cb,+CHT>K2g,T(:R5:J)a>\B:.(J0Pa1geYWGR]Z4;@8=380J(>R#
YXQ,\>P@PV.YOHRbT)KSK01R>4KMJG-=e(I/bc3W-b>X>2(c&3\\1/a&IS<LgM8G
VD?EP7EV8c63V\:&IJVO,+/\L#-BTP4<[TH65NKBO60024U_(DHdM3[Yd;F[VeQU
1&#HS])gcO[)b3M>3JfX^:EKV\aMRCW&B/;R:gb[THP#f-W@?##IZbaFLL3Ub)O,
1_I\D/T(1)_)X_6LLEAVW/J678CV=[Z579Eg0^AO>dcIM=CFD,>=fG8-1ZI,J<YD
K401X3?@c0L1)0OM3:=95ZSB)R\0]XT[8_2b=DQ)<+MD6f.V7<+H\cR1>I>CN\d7
Y-3;74;^J,(/RP]YU5#UM8V4,-@>4ND2554+R9=?OYL^7WL5Vfc&4Z4;81;3<6A3
DGa#d.fTV3D)QWaJ8SSReM?7M>[K++4XBV7O>:/N,FCcKTABCK+==P0dB?BKWFQ]
d^)7aC\d>#-gFQL<O33d>673/CV_J/1U2K90.BB:D_9LM24?,B3+R)Gb]WYGRUY+
;8^;#M+/_5J2?@1P]QVW(G;\@W>,e-.U)a/)ZeMNM5HM>,;_SSL8+\<=&:QII6<6
1EH#U;?Aa6-IS1)f;1?fGT/:=1O\<4@g.7Aa;.bF_F#3LR<;G<FU^[9/:3ZLfNP]
GLb7K++f9<NTZD>P/W>0F:^gCg]71^+7[c8:,>Y3XMd..I?UD6,4_FI8O0Hc/4HU
T)?a^<2.U#/fM;[aVa5@b^)77RaNL#<WW@c9YP,(Af+H6GBDabYH^J9@9K>d-=H_
>LX:#G+LRI_^Mdf([<Z,.KbU)T]g+P=DOEXBOf^Z_6<QMMJLP?MI7-3g3:/YD?Sf
0T3>-JAg5/VgK(?B,G+DBgVWK^RHBYI.Z<c,CR79X1\>_=P.\H4@eO?P&P^F8H,S
L2OgFJd-AS^f/c2;2<M5TI>J.1fT2F7dfV;AJCTeV[B<C^=Z;7Eg^S>VKMBPGMK6
N;2O#\,(AUaTXf7(ROa=)43]_()2F,N)_a>C6JDOS3gd3@/M)R?L5__PPW_(X4N=
Z.@H-4\Q9dAWG>U;@<1V=eZB:[5+PRT.3R>4\@7d]d8\.8bc1AZc0#7TbCL+SIE,
9.d&+Ta:8:HN_?Yc;c^1_LUKHCOZa977TW&<#A@YJdg\?d/#?EKgN>[PFDUPK+C_
;H]bUPf/C?=Te1N(LLW,6APNH<]KH:.XZTgeCK]D,9MP^+I@U)8&61,FKOH=,B(I
BP4G3[K]AYI\7I8#95#LU6gKLUXBH>8<,.D]?-4G+eA45M-:@Z\P;OTZ;F=O&TR4
<BAMC>=d,+],Y2+/^;LE=)^JL8P)WA,.HGZ(MVc6[AA>Y(1\^=?A?EE3^G/1TKL<
N8ZX)[g29]C(1.F#)bQ5:ULeJ?UD,CcCbS+HQ2TU=K;e1NK?ZAF:9H)EB[71[C1_
b/VE/6MR+(+QG/G=Ec17(L&W>6A-C.?6aA?\cT^CH6HQ]L)c/MW\7bXCRKPTdcS=
2Z<1fSAa.\(=EcC)8G=Da2\8C&9cULFe0Of:UOP?W=IQ5I1?3[E,bKW]THM@NP,5
NQI(=??HVE\PFBf[G03##]8IDfF7+0V1U-@K\JaZ)eD<GcGV(IXGSHNf_3,XW<e(
K^=U-+0/URDXX1;0ecPFB0:V?\=e0Y;.,HV>UU[LEVJafa#3SPQ.B+RY1J98R/B\
N7#BN@/RWO^M_?M,bNPQI^4D_XHC)@Kc,DcfFDX<5A(=F066+:XWHN]T[KEEVY:H
Yc(&4R6YN8JKRPPT?dMf1HOL&Va_gb?1Og2AEW<K<[K(;-+L<+FK+#&ccJ\RMfTW
P<,OXM6eV)89=[AIfVH72Xe_2?I^4aV\/[F-V_943^_XZJFcJ/Q2/a0+Q9U^gQe2
cd0M^YXAbNF3C:@GBd;>,YN8;^CQ[N9S(JC<d8+FZ:OUIMO]Q]3ZMN0YG;EIS7bQ
0d@PZ4YXbVM6,K+ZQ-fHKQPTXIHdQ@@>RLg8GK.I/V/0FJbVWK>P?VIJBa9bMI#7
=&<g-CRJ:O:8);_CI&9BW8g2c7;M)5VN?E1NL+C28f-U.)fVf/#&4S&49Z<3Z9De
Z72+SK7:&2e]4?0aCSPA)E#_ZLe6SX=W.UP1ZG-O5MH]/AQ]8()V^KEE>DHF-O\D
2731VS89/,TB]eVUDU8?Z9,(Z\P]Vdb.O)&LG#0f-#V8(f27D4ATA<bGXb)JC&[6
Q&YE?15JE+bEZJ8Z\YU,A6[UYH_KTc>OJU^0^U88J59=[LZfN@2/Y?PO:_<MI+d.
SP-@Y(:9[>>e=3QQf^L+)WOQ5D1HOeXEfNFG],F,&9HCB51;c,4ZJ..;F:CSZPLI
WE,,4N>24HZa2eEXbO_AU&N@6,F[WN:[DT^=Xf@Y#cU>7dA([V)/8/VbP;LOPWO:
,[[93@):PQ>eeP9][MFEB6G<HQG4dNHD(c:VU\L6@1#FSa0HATN=1MZ198\OUN38
RHW9W8DTPW\T#gE@QTL=_?S0G.TMCfL+F:@T_bec4IULHABfT?ed-?IgID#^E_1#
[U1<U?SPEWK,bA/M-SD8Z0HX>14EVNKUI)SY3BR9^=J_3(+a#2Q946>WE9)HLZ-V
6b0=R0(]FdE=X(-2eK[ZID?-Td]1A5e+JQ[CYZW77F,BC4dB=:?:e__+H6G#@I/@
./.R,E[b5:)/HRDF7;D7_B42M.+I+<=D6\gCBY,]]GaP>LcC=N,Z<)1B:/DTW<QL
(]T8Kd;/FO?a:gF^B[(2\^(GO[C#S+G(]9g8#8;/7fYOYU3\N#FTX3Y>??N8I=1]
X2GTYa3_65Q42(4aNW]=gE#S5(gL64?YK;bfQI\7(HE4(Eb]>VWW=eX?\@T)&:3X
5)6+EG::fU?,G)T=(HL&N\CG,[NXS7bT#&@(@9d40#DX=UW.4AgGA1daMO;JdZ7V
@.(9eP[42)P5O.Ee_4eC+7QH&d)Nf<D5VZf@#4#/YWa=F>A5F9R28B+/&=63/R;5
R3.BaEaGBTH(7J8+U-Y(2.CLFGIN=N--c6;d=I=&A<@3b3H&D?\cRQ8cB.5L\A[\
YXed9H]3;YKce@ZLSD]>)UKa+1b)1=&I;8AU-FRX-3<)5L(cfA;PG(WCEC3UQ[<_
E:RVe+\/P&WMT?9::R_7SdbYER4M+Y\Le6-PeSXf,>AS@T3B8_FP-Y1<d,JUI9E7
_;BNIB^NNRd:BfgB:ba^(F3fbb7VUJg&\J-J[MRFe:bYRd8BVRHSCNDZJ/MT(Z:A
@#GKe=#6<3bFG7W>N0-2XD>;G7?CNb6M&,E54XPgLZ1(cPWW39B&a[AL_-B4R0N-
-:e^]aKJY&=d@DQdM75Q&&EM-8W/#2&U8E>+Ad(,Z_O7b^>7V=G&d0S2X&SZ7Xb0
G4_()\=/BJ6C2d:HV748aB<\J4<83E9[R,KH]DXR4N:,CL<+@b2>/XcH3/GS/;V[
0N#21e_XO9:09^R:#d+4H<M-([,[XC[2>6D,))T4d=?SeT,0eKH>cNF+AJeE#6?;
bQcfL/>UX6?VT9.U_;I:VDbA__B3g[7#QZ&U3LVfG,E,=B1aW>7DERdNCF2f5)/U
+cYO(-R-T483fG]3U-2<.N^44YSe+YKM,U<;(\-K\;02AbY93Y?]Je)76Q&@^M@N
>&U5:DE==82a5ZTd4T3#dMC;G0B46/#:&QV\f_Q=G^<d+MXV:P.:LY&Y[b.(>NT0
+8XB)4T5F4-J^XUU(MELf,bCC##X>2FUKdX025-0X;?H-f9^KN@[b,P;@I&CFfaP
E2?OXCVGDeQ2I4gL:.O>J@9FaJgDba.WV[,Sd[AW1&1U5ITg;,,@eT9e-b>)EYN\
d+0+8(bLg9UHTUQUUJJ1^-)OE]U1gBQHUZN)JE:[PKHQ7QD6Z]4dF:Z/YI-4_Fb-
6TcV?5#J5,\>VY50c#58_cEb5]63eE21Mb5O9MPHJBaU6P>8C^=\OG4M>]:#:>M4
V.A9f-@O-AH-#<^KCJ_\5^>b&QV,Geb19M21aKM:V5^U&cfKRF9U0;VO8gJfE1-M
ZB,SDXbOV\92HN/_ZBZdSJO&K[a&S[YN0XU&g8K<:_5N&Z+:Ig#CAEVC&,8^D:-I
D@\.4A]5#]g\Y/RN739(G&=(DT86SdIcc])a;b-KV5;3XEIH)X>=41dHFM/ZRYF2
>W]Q#QW],RfG7ZE\#P7#3ATf28:SHK&[e)LZE<??<NJ1?;WHM;LOW7>0bVg)Z@VS
UY:#dH_+K@[f0H4H_:b:O;KJD-4^3<=X2S7&dB>QGC>\#FM_/\(D3SGJ3X]><V@F
W<&H70A#e>)P9#+c^f8_6C8W=:>a>3S#@J6];1OLM;IJb,_F3S?V^Y4+87IW56aF
<Z_#cZ1)\W@?&6HJZ1TbIT-.XVYA.(./M#[-(aQRdPJ.JH_Z33a5VQ-bQKe+;7>A
.WE21YXUXJ[Z42KAY\:Z5K8K_)GbJB(&3L:#a3R(Q.Na)9?Nfg[>JVBd@Vb6fDEJ
1Z[-dN^Q&JM2a57D.[KUQF.]d&f4,+P/S<4RK^&Y+57(]QT5V4aJ>?5#)VWcW-Yg
GCXX&8ROcYZg6=OOgC&X@-F)8Ge4\/)E9,JW=T>G^e=cB<fBA5-aTD&W7&ZaBR5L
J4MXKOFY24bdEgOMK7S7Z85RVJ.Y#-a.d^N.c@;]9\=+)<1;YKWg+DF+aK;cJP83
,F@UEK[A52A+S&f.1AI,]b>d-:KQD;X7b55g;[g;5Z5dgS?bF2@Eb;[P=;;,QFLT
e3b@QX72G6,5d/6;)8.(:43aGd3ca3VcXP?C[OP3(>NbP,[.Z0g:LQ;JK8GD9cCO
O]OaZ)fGLM<D^;&WR\K^6eUH5=6_?f15fWWRH_X:Lb.Z=c&eG9EWN@Z[KZTUDI8Y
5:-]U>?624CDOLI\AgTYO0e>f-gKc;G,_@c<U1_A9^-7f<dS_<#0#=SP_S2H@UWN
04#MbY0[@1TD6JgF:I3-.IBRFZ@DR1TdBP]8:VDG-fV057+DA5YFBP<1>G2(7T1]
gGQaa\a(@YJB]]?SUfFe\.\?CB-Y&4B4]f?>>?8Z;Jd+YRPDAVPD]CR[\DM/)DX_
d2O;N?0[Z;<+fQU5&W+Lf75Y^&S-),?8A0/FaPd:f>Qa_GLMZ4,a4.IcH6TP7IMV
DQTEV??ZP1S(cbRa)N>L3,eR/MT9;EN[>/DSTDI-@R6T9WE4KA2L1K/Q5[2:cAb&
cfbZ&)H=3F;YaE,7XRb(F);HX<4a;.FHO;=\G]EM(;LJM)Z]>W]c5Q<6?IVM7gNU
>G)-/5GV_(LR)TCN3gO6SRZJD5NVW6()_J1P+2WPI;-=[aH.gcO_Aa0<;-/(YS_#
P/Ed@_.XM+8[RM/_7+E:]P=74C)b^9^>ae,(,4FB#Z6;c]5AeBPZc9;KIM1a+.(2
6<BcT,4b=GfI5SZ<]ac[QW+(b#_&3=N^HKVR&]CX6b5O<4/V.P#L?E&KVD@P76V;
#<Wf1][bKB\+5f&9-<1KN5ZUL]ad5O5)6e^_7YR7HS?dL;^74ad8:eX\9FGZZ;fG
^)2,-AF/G]5#gXP8_b4TL&Gb/.M#OV9A:ZWV,ZgOOC472WbfC2cDS3_)24I]T_2)
HgZQ2WMC)#2,KTQ_J>),_Y9>Y;Df?;0=?VH=?fQJ,08ReT]JA[7RC48;aLe/VP6)
a#(BXbf(?VCDJ#IUF6H=<=4XaQRZ\3UNc-;&2<LgJ1fO\L?QVSTM.W(-&L0fc#_F
M+8Td?2.AL<GE[L5S4E7=2Aag/^AR6^FY2U&J]:1(b4K93;PD8[HN&K7<1<;WIeQ
]YcQ.OBL#-(cC)c8PbeMc,;>8PPZCA\cP_;]3X1OY5<6MSIK6S7M9J]\&=B_K:Wd
&55EZ.YC\G#+J@#\#MU+c8CNI/_ZGRW8J_-@?HP),EU[,+H<Ab?fg->S#gQ]@<T=
NB[F/DXU=,.<(B^70T[U;_3#5c_GE:Z;:JV][[UHfeFc(9G.?:f:QH_c(D&Mc9?f
039XS=?e98P^OD#a2DVH^bMeUg)b912<aXUa1b>^9CR^=7c5@\Zg.]<ZF9:L4Mf@
P#g1PE3H8LWWSKO.2+ZB=Ia[;^GP.QV<.16a(L0MF.V#N<&?-[R)7ULKZLW+,5KC
I=fE;H:Q9/SP:/2bgXc&6Y#6,+7-\f.D3O[09(B\R==XNc6fZG>17I\2HYI2O9W0
\f8U3-:\)3PVe+ZR@/H0IX&T.?TMcVccdaAZ8W8I9J/[LZf8DaA5+?>,<0[/@/9Y
,a7T6I/U.S1J+^[74N3//A<:VBW7A1838SAd46D+.d9I5SYG89U&bX8B/>&A#;cS
fIN?\8(6(JR5<<aQSZO81K2HP0:HEJbG^X:82]ABZ-V57.R+D=gg_HS&.S@Z7.TG
U)[5NXI0<BS8G3#,P5Gd11S>B&IFMc2T;,G,:Rg0V(ZS;/,C2:JX.LI>9^8P\-PZ
LM8F6EK],L9&BZ6d,?:GWc)?W/c9S49#4E7D666KOX<O6#C[U?CCbVVZF6?Q[,)B
+.&I@)0=(L(c6XdDfPfOOX+R?I3R.R;d,bYc1ZCI07O#E87KWJ/,Fa,EZQHXLWWW
9]7WRLcUDZBeQ/,f=5/8<.QB.DL@3Z=LYfH84+6.H&H8W(ddI<U>1L-SAQ,<0>WL
;1UZDTQN)bUP<4TTa^&GU)U(,NR=-7\-DSdGf<We;?>>T8[[22a6.d\HNB7Z7=;K
L<B\MN166EC;TVQ/PH[4--;C[76)K1/MgL8G-C=P0O?)Q6-Dc=^RfO2I,G8A,gHA
S;19R&?>9=g:/Z>KZfbVCZM3)=?O>M]2,a3\:4B=VaadY/HLCcAVUV7WOKc6Y<f+
KA0HfSTd=DX=;BI1EgeQL_RATEZW88F>J^ZMW;S4N+)2&FX^^;?&6>:SVMc-JM^E
BA682\a_.,RQ,[:[@,&2@S3-3\2>]\IE=aD/Nd8C\_?5+.AZ;45XBf2-).f3S+(+
5&e2fME]3Q>JP9QY/N\1XU-32Z-H1&G)P&69+Vc6-U=/I__2d,I/f?ac)K]W;a?-
GDbKV\/2YIJ6GeXaMZI>ZV5acBWI.:eHR]a;R4WY_5/G0bG;OUWJaG-_L18TU#Z@
.W#_Y1MGI&>7?49?4/Dd03DE@KE)W2a^VN##TZDCWOf5V?R43GeZIGCD?3bJYV/D
DS(SU5?&P^+SV^7K]1FU8O>:JS7+NERA?&IaORTIK#V.TaE/C=Dd<N[9B9H8EKGG
,ZdYEP=++5dYfK+A=N0ODK#R(7A[OgC6FR>XGL((T?d/K;e^HdF-H;SR8cY_5e_W
F^_^J#C3RM>SKf8KG0WddRbYGOK#FFETc@^SI;-T\64eE321?BO4T#N)3P-,_K5@
O=d4d)Oc+SUfY;)+\>K].>6VV#]g6XC?@Y9[4@DF^0aA08W2^PYLVV7D#(<N&V0P
C3?8AUN3(_(=G-ET2bC4@c@;f,7#0f^,P=,<fdPdd/5GCD87EHYL&DQMd_3HNYVc
+]M4W@S]/:MK+Ha=+/(+/KAH@O&D\?;.^ScPD2J<fBGScWS;Q.S/.U)8]RAM,dAa
0(KI)W-E<9\fGc9./]02IbI];B(eK=0BbD=,YUDPb@D)R8R^KaE5>PB+#TJbTE[B
Md44EDE9KW4.(+.dGbC?)(3#f^>c?NA:#MC9cA(?M9>;+>#dZN+C_JJ>fN(<A)-Q
AJZ:0&-.?;a1UcSa1]b=fbRDND?RObc5+dFgga2+];BN[c\=.8#<HI)W,2YAdXJQ
@;.P/B=S<Y7c.98SW>;?8GE20(G64DQL_>aSE4aYB#>L.fYY;\I_JW>33?O^)Q9B
aGgdX;90TV7)[=M1KaL_]<0UWgd37HI#5\PE55J1H6XbdK.1[N9.:UG47bP9?+;F
<,S)LSE2#EGYG8B:cA\-a+[@5T#H/S9gZdb?LY5SN,9U/72:R)-REdC4\#.YFI-:
W\a5@2U<#I\^DNHZ_0Z/(9-?RJ+JOQ4D[LTHL#f>:H8dNfT:]YOV)JD.gO4f(f@<
V3AFd6VE)SZXfg-E+)]3;dC<9-f4-70e&#Pg\)H,a;ebHPI/[+X<M5W]^,gb\DP<
c1=-XQc9]HS<XfM+,2K>RSP>afUT25:ST_+QM[F&WdKP,Wa+2cWG2RLRHNGad1KI
\OFDN];R_6BI>(Q5=1WY6NN/]g#HKgf6&A12G?DSU?JSS7cHK=A0I,K]7#SZ>\X7
C3fb=>T)[La;GZ<PPc,PYfUHQ;XH5<;I(8[MBS<4(YCg;ESI]+G=BT0<Lae<8X4E
H-?;=U3=N&TM=C4>d,+TB:K0XU7d-ga,;8FO;Q;W.\eHBcWC[=Adb.B3O\aT-\66
R/TL4WdX9+OF6),HE(45Ogg3VdLDb.W^(8<DNT3>eR/U+<\X^cC+bHP@AgbR]:R^
J=NaBR@W/bg727d8CW75PH#T2>T_#6;e5C/J++^-e-ZU.,&<I_O?PdI&MJU-7g0^
)6>.<N-b894dR-UV5[(,G2PCbPb@SQBSf3:PY[>48/5P\5#FgQUS-=R<eSV14=+K
3NFE[K[OK)7aB>4VA@;Hf6eEQ.B9N/D8;.#e+X);-5Z8?(LHPHO8FeP2Z#[g9MAc
1Y]IcQAa\&__B>[),aB/.,5FLg/7RP+O=,#9#Z1XXYVJ8.f@Z[HC;RG4MJ#91eb(
STP,^c8CM4R[<+^@&:MQ([>)S(W(54,_G?):?0H5-gTBHJAf<gO)5T8]WF@VW<6L
b[]R&+W-f[6A+DU3]CYIEJLP7.[[@K>K28-</Z[:aOHTc0eGeaB5&aJ?H+LBQFcQ
NRJ)X&a\>\;T6+FBQ#^7:=C2C-a:S<+6BXaRRa\YHRWBO3^0da;FKI6LAd@;9fIV
aZG&a/W_X=C9/#EAHI@9]0SJ/g7NM=R#;+T:WS&2SFc1YEf?W\_d]N<&BQ:/Kc>D
3SeNTYCXMdTW,Qe9C@/]aJ=c3SgWVLQZ;8[UO:YD,OIDAFAN6RAD=b)<>75C-E?R
:/LG+Bg>=#?H>eSUFF#[XS.EId.f4,V@<YUcJ#f5WTAfN&2(N8?>KO/2I4PB?_OL
6aOWYYUeIN4cZCKNG[^JYF+6^[Ya/SQXCNCI&eJ>ON_PAbfB<I\<Fa^=O=EB0(b&
1H-,DPaS-eM[61XGX\dc,[=V^e2XVe[TIM8..P77bF^8;7-X51I:HX2(>E+=-fM7
KRU\=a0^.X-T>Vc\W=;:HRKb/,FU[_?NMdDL.cBc-G0<&9/VK?.77TW]@8JIf^0B
L:04Q.c,,aJ)X7YXE[S_[IAeO9A1[R=Q&>](Cf_fCG+HgK<;U[ZAO/#B4>@@8Md/
c1BJ>3SRB=)I7Q<U?=2dN</U8@L/K^ZE>[]?QQL@Af&9;^C8:[L34#DT:,8L[+AD
64aZS-05FgN\\WF_c-&?NGO35&=1,)SdEUf&U5_1@F^B8BBLJP7W4U9Ha^LabT_R
GLf+8A0#5ALOY2TUH^LM#\gbVDI4.3)[_]aO7<9X1KZA.QDTc1^5::)-,Z;:U6T_
LLXYNF?>?4)WT=\<?A4.Q56fMJ+[GFY;6g+&_-=U1REZ))Fe;gNC7a)2_\;.2g0-
,?1&;P;Y-Ye6.HX<Tb8fI1.RXGC\B\@&284FM[)YHQFRa.#L)5XRU,L^,dTcW^0[
@4&MOYeQ0#Ee&VNQ7UNPH/E08+SVQ>LfIFIbb2&E,:dY1\:UKEP:#K[f>3A:0e1L
JKTMX[=BZg[O[C7?9+HQC+[F#:O)a]N3BO<V.Ig)Z#EQ<T9/eD=7_[\)E/L9HLS_
/Y68c&VQZ3]JN+R23)DV-^<Y^:Pa]2D^agF-D-#/RBU1P)^2L)GJ/\FcVCg,NTe.
GgY<WReWe?RF9Ba0?Z1X.@AfJGR>9XTI7^8I\9#LL^L1=94),:@-S@K3.IWE23NU
d<e)Y3eB<cVA]]eHFf4D:c,L_F3B;[\DV>/@KQ)0L-M[&@/G,PNIeK;FSW,JWK4W
O)8:6c_5QBAP>@Q7<+1KCK#-OH/R\gB;UP\@:MHJ(R3.=X+1c1&d.;BX>))V?:C8
W_[ZOR<CM,90a1RUN+.3TVH(IKK-9F5JK9C^^E\#)0#E_>G>7XS@6?7Y/f\?O6PZ
72f:=,2I];KcB?d.FOZ,G,I8XM;M/\UeQ2;L>A?A3:)0ZKSa5G6^4Jc4:3Z()Ga\
V<9MJY2T2457IM&FI=Q18f)C0:RefOWa7<K[cNVS)ON]LfS+;f.A&E54U=GS;C]F
ZNQB45\Zf#=E6RAbJN1NO1#>_=.QZNQQ)SH>>V_\eX1<JS5&;RCCW-Q?ZRX4./,^
?(_[P/KDDW<O\7LM7K(5I)P6IcO:=2F];9Q1<?]SD9/;\4U4NA+[TP_Ff1,2X9Y1
QF\eQc\b\E#<I]0dG[U5.Xdde2K(L9HBE;N)Ga:[g;,]T4gYJ1;XW.Y:dcS-V(c@
e7&1+0^Y#cW\1/-AAebB.PF72?^aBX+M7@ASZ8?Q]6G[D=>Y]24PEQ9OW3R,?7]]
7?>10MeKUT/R>fS.T,107.G14W5133.I8SGI/>\+:0[Yd[(O).=0I0<AO44J9gfG
/EO6F.NS6_Rd]]8L(.]Te6O)_3&7U74fD)aQ.aV]UJZDVVKB3,FT-[@^GBL,@H4g
6PNB7XGf6,&UC&(F::>E#_a,L[;HJU6g7<J_]=]D_I;F<^a4CIMcdKLB&N<bgM=C
3-U8-W7(\M+C+2<P?1X025_?05#gB@UI=d\[18MX-?V[5<(E^f-4@M2gMV,<9(Of
BgLeY<LfQSN\K>I)E^V+K\V9>?YDGO9J&+CLL=:-MgF-)_ZX14-Z:PAEG-;8XGf<
>RaK&P;=&S(EQ)03,-=U>(=^7STESANJ-O90DGb^.7Oa1Ya10c&g/\C1\d([5Sa3
1,?JW2dRVcN,NR1+P-II)QV^f#gV>SQ(CPOJW4,.I>Df6+NDYW+cc\[?_SY7-UK:
YeT/-N6@:JVaMGLg\7U9K)(0337HdP#,d]DSaXS2(F@Q462K-Nb[J(?HSaGVKG=+
>0MOAIgP]48:P7a-\,H@f;6(#87_c@(f6GK?dN.85e;V=B1(KWM\,6eT\?aZ@^)Z
NKQa9.\]Tf=PU(a).&f;c=R:8^:D@W\-QGRbGM^Kd<+9UaN5-JO(EI,:(=ICO;V?
=?G<cBY@,6BaQA\Icbe,_<CVZ5PQXdWT?.P2&-Z4P4@LD;EKV:9]DSEWR?.;TYfN
:DR<B^1<[N>[2Jb/77@;A;P1Gg9;59-N+0N=[bV-1aDTfIM<U]LTNDPa,<-gR7@?
CTF:aT6DP-P/SgFHC&bN/1dK#K(<a;(PBJE+WNZF8;aMG622SY6\a7cYJV>4+E2G
]NfO;d1.][VRbZBZ3S>LI@L)130g=YHCf4\-&7[c58(>]SF_X81EA&<eCQAUU_-:
R9\XS-Q].R^ZSK@@/8g^@4E:)HIG3Z+)L81<HeCc<P-S(dE1e6Y4,Cf_C,6=g<TZ
_UV0PX<V;W:]Ff;LYCbgMLcN5JK-EZXXZ8@dJV;<],K#K(N=KRd)51:]56/9C]X1
(&OZR06\(0#X-/-RN[[d]LTZQFV9EZ5HB.J1(4/?IWPI<UN4&MV?1=6YMTRc;=L3
Q\IVP;US/;M)4f[OWXP7add_:9bY-OUCQ5b(J\@#[N-dW49ZOe]AQIJFPSK:8)87
;^KgT)PYZG1ADS&@]?=]dQ1Ref5^CN\S-#@@WA]/N5S(GOJWb<W\SP\1R+M7aQP8
,aA[L,GGeV6)eKFEC=WU[+Q<_FP>T=c\CG:a4J>3d0C2Z+[\H?UQb<5f/=)GA:>7
I_E34N4P^aT9<:W#afVS0gN89>,(CggQg54-#AZa0=^8<7(fT4#D9M,a@@V+E3I9
MfA4&198d<@PYJUG6gT\4Y5KG/;_[d?<U1,]6D[K@F5.Kb;2WO+Sf-,],6J>IgUA
dVW14,DEXN5G#=;)U7F[ZJUWA?0I6/ITO^A#3U:I0[/NJ8Ac,B@eRYgRS5_3Qc-Z
/7##c/9cT/O2>,_V(YR&]U1AZC0e^6>IS^a-RSRAXcb5.AYC[MBA\TdZ_LYACP#Q
F+6_Tf]Y,1<U^6UU1D_^HbW\;0[(]3+#eWQbOJTM_<PTRbL1?Nf4_DLfKR5Q9&RT
GAJeV8.CS>.H\I0X1I/SL:g]QW&P2@F^N_HQfM4XIAPTSG(/JBSgHA_DO1V/>/IS
(Y1?QAGLPKDFW>5B=5CER?+27Z^<Qf-_&(R]>,fLLLJ-9L3?9CZbHR+=/fBaZ(]A
g^f_dT4-XS26/[+d4gb@00C:QAeJY/Z\D[d\-BDLTALbAFGBYC)4+ZF2Wf9VQd9C
>c&@F+RJ:G#fUeX2/DEdK3)+Y>/&ggQBL]:W<BS68K0BM=6@D-_^=\[<J(XJI<VP
(Tc3U?0B(;HK(g#9)&23A;0PS]PL6=T+EP7^e0NXGc)YZK?:Wg8YYY:H1f,Rg1@)
_F[gGOM]?a\ZaQ_B[CV=;6>)e>Og]9?#aSA2A8aA7^M1C?+QQdB=7I5ef@I-GPGY
(T_M9YG^IAgS(MK?9KN_MNY4-^O0aBc[FD^TbLO^O7^9[9W0P,W8H;K-J\dW+4A.
-)Of8VVB11e8cR@3H@6e1LCGDNK2)ZaQT&==;W2EN-(-0QbJ&U\S?(>MO<OK3C27
)EW]<(MbT+\CQ<=3ZB(2.^?Wf073Wa.(@fVK=eUJS;96D2(e\eJVd8TK8F(>(N#I
T=KPgKd8@X9[/f?#@<#]V>])8NM9SZN0e2:^=TB0KIQFNCU[+#]M6B9e^\1U=8S.
OSTWLd;Y@K2@,Sa&eUK1_K)+KUE4EEQ:0fe-?K42U58OT,N;NA_-#Ua?.U.H5)+=
f\Uf&09FQVZCegT-Lf(cLORC)5._]^d7]ORVN^/:3)JF>7H<P;8e/TUAbd;f1:81
&S>KT)]d(IaE1[1X?]gK+:e@&T??a4H]W#dK)Z1<e3cY(S<)EBU_JTC5N_TM<Nf?
&A\?63/@]UbUbI:eH1(__d)@JVW@Ue:/(C1WY8W0Q@[\7.c/K.C3HbMF+K[835>c
D9ET<O75cO6eF<S:Xf)DS2X43fCVH=.CfF9T)=S)IBHZ-FD/:6LWF@dIg/PE5??H
5[A\Z8L5-]L_RYaX2G#HGScM+K]?UKdW@)M<@5\KYc>M^SPF5eD7T>E;17(0&92F
KYVbfdUY249LV_^^T\]b@SKa.VI9D\94\abaSF?#2>9J+T/d6a.:(,#aA<Z(H<+?
]YHIR&2:;0L9&]VEAGGON=d31WWQG>:TRX<#O)NRDE;[>cTBZ4[LCZ_:ZNaS=E3f
VT14P8]+NMM5Z?BQUBMJL<6(QB.Q0_H#0g34-;7TVZ>U\W:+,af9A@7QcHcd?E\f
Y7:(/VT34,&.?LZ)M5D@GZM+9L)^[8@=b)J;_:L&Fa,/SXLD=>MAW&O;eZ71R#Eg
L_8PKQ1.c5eWYZ8OZRNLbNO/I,HCaFc7,^^B8LY/5MM<:CXL>]cK;G<^DfaR)ME5
<-c7[A4V]A(6&_EdJfAMZG:X487518N4>UDg.-4<Wb&LR)R_gC2WH\Z-=1\@0O56
Y;0-<fS/AY+71X;8VCf(2&#KdD2WcHCdUG)AEGKM&U?L;[V##)E\?=3ETKG2@b[0
NW_JR,/;HcZVMFaKMD6.T5)a_PGUJUA\e-(g?dML\Q/^,b+1FE.Ae,\cO;VN_I7,
IQJ.NZS=47I6#@d8UXS?(I;Bf5ULQS5@f1(XV<WMaVI)cFJNYUQ\)KXA[3+[0K5W
)(>eA(&73C3FLa3Y8@_BYD/<>#+a#bPgb)5;QB:XT<V?gCLQYU.V5_A@0#@&W=&D
35Q(3E?+=B#_^RAaYR+O33DBXYd>-Z,C/D[AUR7/;>T#<V6+Jb>2BB8:CX2d1bU4
ZV^^I-/GA14RA(RLST_aQDC0XU),F01EXV26J9(?#^N=(If?5AB=,BHZ.feD6+<L
+EfUL<?(a5<N+]HI@@g15O^(,2:&BU>f8gI,<99(1V69_1:6^XfR&0Qd.BH4_O47
E\=;b/&K&Hb&;8^\4dL@6X[Dd>NYTaJF_<(Dc9[?7+Ne1&KD0cNR)aa2aaTVHY(O
(^IW:(_1AHZ_<aC[ag>.Ra2:TY]]2[(3,(LRFE\X^18^&?aGWTW/VU3M5VIXbd,d
g,,5CV-A:\\/G[aC7_YMfO#_\-Y6/U11S)38<Zc-7#9cNDKET73\20e,O:FNHNM6
O1dSCT>(YNZ;;Lc=>XRB&b;^W1Q+=GFTX4>1W+D/^AcU,(2,>T#.@D(N;NS>\1^b
+DI8U@1[K/Q(ZXTf]f#?@BWON=;XVga5NH9#<.B2\_:H^,<[3M.IRag99L/Xf:\S
;/GdD5,R/c40,>9=>X>JT0OC</9AD\aWES.Ab@>;-afTH,3DJ+c\&PC==KJ4<SWO
LXc<(@9+cdQ-:NdT&F.NST4Q6eff.F2e.4S:E)4aR+4TJ=UQ-^PL;ba077b,,[D\
&If?JC,,Y+6FFE(+g&>5<@^>a2(E2K1K.E_Q,79_6L5Y>f7(3YKUWE\,X:U1;R]Y
<Y5:_)Q6FgV@C;@fJ?ZGV0aG.Q;3)KaZ#-5:6.TI/4A0N\F6QS^b?>TO6K0Q)[.X
f.YLHgIP7a[0=J[<V+YY<f8Z?CW#,G,5.=_6>G7:>L48H>.4PB8NRMC7f&=aD@fA
g+6(0SFE[V9P]#CS9[gNT^4+[Pc5Zb7ELM9G:RMO-RI=@R2ET7]5(,HR-O&3+[Ka
:^f#KQf)H)@/Sb1CdWI2X9?D7PgPW\YMef,Id8Y0&gK-T=f^SEGW6bK>:ET_+4M8
1UZFdRG[dF.d:--K>519(1db7IUM/JNU,8dSN);F-VMFW\59N3_d=0:e\]6bVLCb
AE?B71=LG:A)+7?>J8+Q(<6#9Mc.f[Q+dSZCSA?7L\L,/Y,6[:K<dH[ORb:N?P<@
#2I]ANG7D1[_fdU,Y)E6D_5\W;AP;34/B]5g?-\PB=F(f:1?.)>O2<K-=2aN.:Ud
1?XTTZ1Le9G>R=#6L\;,fJ.G7X?VB/C>BS2)AY@)1BUF=EC7XQJK=>-V:J>CGLGA
=S^P>e=2>gI\B-GX3d)c&U;PSR<X>&)a]^IRFW[_G_55-B@IBQ.?(Q^cQ_C)d4Rd
&W8)P6:+C)a>;#>W^@(]WHLTH6Q4.]S75@A84cVg(VcO^cL2b.Jf?d1J@Q@/LPd,
cDUNQI[G0<?ga4d/L_KV<M]e]+_XYfHdP?:^_gUE2O1+B0)dDXR:<:E/&XOWG/49
ZJd(Z60;>a&<A^a<.I[I8OZ)K-EA\[dbN:3=Q>:#LHA(;aNe/0MRUS)[T(T163#<
c\5aZPZ6ATP5L:=;P3_L]f>fH<._3OA2-H>gId>&G5U+T19\?>;LYM:L&J>_EHAK
/b,MS/If(:=H>DWb9M#0-OSKd40)VSMb0?I/>U/d))\F^#J+LD)XcMKZH2^\ML_\
LgWPU6TWeDgDF9TG8O\.8._KRMT@V6I,H=[;Fc[__cJKId4[#\,E8cLE_Yd/?^.]
X]2FO+4^LHO_W&IeG0eO(d\SGE@(@;BQ+],5ME#]_ZHMQL@fbSCD/(3]K02:>+,;
(e1gZ.@Y(L)13,79aTU9/?O.TY1N\(&)VScOKL[8N7eEa^7<Ea?2.^BBeQ(FQR//
^./O^(QI5,BS.cXcO^)>F?f;ALc,FOJ#[T4NBHZ0];QH=WFDGc]K]M6c/S0//N#c
O6aUCf?ZGD18d+@MeCNT(5]9@U:Nb+A7#G?)RJ#e@WQQ(D)Y_AYc9+.9H\-.::aH
=;T+7<.c)W5ZU\U5g(+?:@YBdf52b5KKG(1Xg7(@XP4bdKWe/dR_(8ZI>K^Dde[2
>6O_BKB_YEM3<E+MaDDDXAJL/-P@KbBU7N.45&6=FXH_^b_cH86;HGH\+Peb_<,Q
b^dKgTQG-B7:[]ZXW?V.L<B0TO&d7,UO_7d8\d>,M&_:4&T#>W+c3\ZQVVT)81>>
KTL)Xb95S/Q:W9<&X1Fgc_QOXN2&g9_82Q\Rg9GL,7g_)^Y+L=GL5/I\]N2.J4dZ
JXf7,_1V3HT@f;3.b[R_9)J+@(TDUX8QA77eD6_87g7)@d0,N[[_YBH,^[B2[U(7
;PA+]HaPcVe+X\K).<<9FITg+=ISX@]840\PC)c/c>Y_=:23?a2-]HLK)LGUb)J?
#5>8_DfNUeCf6?/VM2GV,);)RV/&KLN(J3GE>baPgKX)[7g1e@5+XIHNM-4P\(>Z
[03+ZFPPbgMZLcJ1^ZSW5JO@dUY@gIEF5\AF=I7U_F\O@R05<fg:7@F0ZFb)Q2H;
[6/HfT+@+fG;a1F.4DX&Z6Y=[NKYJOA31[E2H+TQ]4VOP#I#693JKCN7:dWdG>fe
-8dV1Xe#@e9LKP/Ve+f<@:9FG9NH[#YI3UX>UcL>T?X].EEI;[;XXU&cM.9AgV1a
N;]EYJdDe^gQC#0eK+Z=]3Z@\dEaR60NdYCF5eB_&b-I,V^aPBXBgaJF-ad5E>RM
eFH);7O..26(cF];4DW#?1C9#1a,LAJ(f(>>X+91WQWQMLSd^-IGd86;UN]IU<4=
S:ZM=Z&^[HCUUQb[L1eTJ@DCOAX-FeX8NRg8R9g]1ISb7O:P5_+2KEGGFH9+a>;g
W:X4W41UOcDdNZSVR@,=UX/Z6]0[4^&bGSJPaNSN;3(]XEJUN6JRce6Z(=g0=)NW
^/fg=FV#MG(dV=/<c+1\ERY/_WWV60U;P[cKHL^&I?dFeA.A:PZ#+(]dZE-=PcVW
H([c=ZJ+UG),16=CO<3=7(JKK-1ZT[Ng@H>O>S3,1Xg/RWPMX#L)V=ff5EM./g/K
KO+VB/?eMKXL\2E3VH]?B5cc95_T4:>L[QAF[/+JDa+e(RAZ)_G-[M^]>WXR2ZYF
D_DgEc2,0b[=Qg,J\]\^X6H.[^UDID7\1T)=]KG(?1<WX-PS@?[]Hc23Q(0K0Xe)
=ZHJ2;F:SQcNK2X3a/J)8Z?<]dHF+g?6Y8G\K<OAfdR;>;O^)P3-R6eM80J1B6[>
e^UUWU,F.;LN&<\GYB);_UJXF_3I99]CX;de>TI)A[UW4O^C=f,SPV?/LYKaW#bS
c/,Zd^:7E34QPYHP]2UBM@AD(.E<WN7M3EfY6[T\OIB?NFKKE,EJ3.O-GRec#1XC
Mf9VMO#OVYE9U.2&a5Hc2O?7&P_O>FZ(3,[I4eIf>]HO\W5Fa?NXM4C&2/HZZ.IM
872,<bSACY7W?6/&J[(+5bd2UX^aUT\P/F#SW1QgEYI4T3NPc(9-3+Df&3;MHF>7
<7JN3[4d==Z^>b4X<SeY,<9I+d1>K+TTT)NKX-VPFO01bPOOEG#f[E5DH-/U.;-f
?;Gd9_34+BHWHSZ;1C]^>I#f[?Pc;KX/+6-Z@QY-W6[FeK+45+b4c[DbcX6Y\.J#
R+Ace]e65&9#bW^HD[Q0=>TMa(N(MCfCe;0WUQ5ID@#Z?a#7_a_L)3R30+W&3cOI
WC_:e;N1CG]4O.(a#K[RT9fLPbTX-TM.?LdFA31@2_>)gZZ<Jd&<+TO#J)fce=ZT
cF+)f:8D5:F&.C1/XT(JS6Q>cH9TZ..B2FRN5)[VfXe+/7@^Tdb\/](+BMT^MS,^
1,IR([&MGf8^^CNE+Zg(60b&:Debc9=Wea;=O1V@-L,d.[4IDN;]&&6Q@QG/J\,O
47KMg-A@Pd7@@+#@U6dNACLAQbT1\J/Q9g/TM17S19ZJ7M0K7^0+WO5KX=J5AGCD
3Q86MTDQ,-Ma36)&L.e>+>N,5CF69Ba0>20&TYHZOGBX-5g)fcHI(6:7^R@=I&^C
_L5c?=/fY@cU4FAJfY/SfQ^6_@55C@9S</JS30\d;_4()I>Zd&/M;56eWX8/gO=Z
Q3e:a6)HL7/.ATHEf8)UF2?-bB8FQb2fc3_FF3W\^\6dAXWISUb=6\/(.FU3X(Z2
LYg=#&a\07/K;4HA^4K3;>f82#B]X^S/)8BJ+B1e?>#fZO#c/7GJ2?K&5\>F2S@J
f;1LOEeM>gCg08;&f<=,&[[0fd,\[7=aL&6KASTa4>,a)0()U6QdI7C.U=#PG=HT
4=f1<,<LCd:K:DV27_EM96Z6-&_eBBRe3cEV64_X>867N7^AG,Ug:YC2&2BV]#PG
0E7PBd3(2<JX-NS3NZ0Q4RC@=);/=<]WOKFU59N#8YR:8.cF;.^_Lg?T#Z9)LW57
S[\AQ_T#+4Q-:cX(:B/42/JVe0/ZM,1J<.RfZda9[A[FWE7X>@g7\^IY2KNb=Y8b
I(SSdZ;ddJ_L4N9DMG]+]:C77D5<WUCZ0KP(f>KT\WW=3[QV#E50F<Q^_X].?cQU
YJ?\F6X<f]fIG+fGM20<S&A7OU+?)FFRL:XRb),L7#P(<P0e;Y=X,,]R@Fg=P(QZ
ed^aY5<b^gaBP<ZZ=&g9TWBW]]K,R@K:fS1W0Sg<(,ELAcXJIOQ\31d,Z^HA(BHC
)>Ye0LK3S:Y,R@/DJCQNgLSN4J:=TC/0:bNVcVLZcO5MRa6(K/_E&4(+gQC9=3aF
]c^BC+#a:2SM[E0)KY=PP.O,F[)8d0T-WVKSN-B51/Db-BNH4&WgCP(@CP=_SdH,
[@VagJ+TF&Ad(2+]ESYK3B:8(Qf^D9Yb&Y@R0RQNJ_bGUP,bEELG6[bW6-#H0VG8
.>8O-;c-H&F&VB_Q?aXH[#DYDP6;,/C:99R6WZ4/OG<B&1_(2@YICJAAd/>5=-RE
:6+11KTQ@gN5HU&YZ-;@dYGQ_BLL<#?O+[FB](XTE:c&[.e\Da,A.1b;SR7;LL_W
(\@;VP7O3FRJ)#7>TQJ;g7f:.Yg2&Y49PTOc8F,TXcF3[R-I]ZX467fV9B-Ya5b7
IQ/;AIJ#L2fMI9PHC?[Lb[L<X54@X4ZfX32>gV.dJDT(1UM\[0@1[fb\LM49__bN
:7g\.(:6OUf@<a_DYeG7<EaH-=4/KF[8XfT=:P&J)MYOXQ_]8I;7JORZN0:XT1J8
O#KdaWQQSS6I.]cU@13_<+^OVX0EKT8L3^?R_>/&T#gTUVZ/&5H6Zb,-]4BSE-0=
&]>Ke?C42F8dB^_,VCaBDN:W4gG/IZ#.3S+.A37V]d?0SMF??(#A@7=D5/#XPUP)
e=DT<_F,S<>QH>?#175H-[Df>C/-NSB)5OJK)VKSCTOOLeP8NKTbK0JA,>cKJ]G.
H\[W-(GDIb#T\C.[;a9XA_GB)/?O?<A4B15RCbG#2:5W=/&I8PQGC:cU]5D>FP9f
1^MD]7/#>g:IfW-?]S+<1^e30d0VNJ[\PG1A=@VH>d>(D@>O;]:b?FK<>NPO6V.6
NBF/-BXSQ5)L_CVH,,5cbW-GeQIAQS5H9g8WgJ.b>NgM<6^3BZd,-6f8-LB\=K#L
?A(QeG.UWS\I67KJ5VI96JK>Qa#WN7W-&/=><[d)+\85ALN_&2Pg)PO?a6D-]_00
QKXGP//8dY-JfO.H=L;</,@5b.^K^LZB[O(CaA_P1=S_:2@3[:S:Ie>XQJUW1g;9
T.>;F9&E+eSeAdO^Z<[UTfDA)X7)#I1g>_3_C=g(cQ@5WP@F=Ha&QeRW3Vd<4[8Z
2MO_W:9DA24MMO\C.DG^D:@K@]1;6M[0W\)6KAgCTWR.RW9NCce6JVO.,eNI1eY]
7R,2_-80=U128-ENgHV0c#\ggKMTGUG@3HWP>6ZcfUg&5=4ZL_JK,:LURZ[BbDeQ
cgbSL96AX8,NEVe2.FU0@(PO@e&7[>a[U25I/2VL?d]gV09LI_1g/.D\FYF\_:7d
S8.9I>S,ZARb6,<cFMB.I>:2W_S,RRT8MCO4?^Y12BY9I+WX.O9PD,&0E@JT1/AL
[d;bSFHH#(U:)?31I2]S<.@OOJ5#I#1XWH.RYI9.L\gZ.76&:gV4].a)g_F6N#=9
&4dF0VT;/6c,[dY,0a5QJ>++Y:O=]5CgX09[,3a5-(b\_#a5CVLA&P>[PB&-#;Ja
ES2FgR=(0fPSDJWQM(CT8aDL,L:Z.VD1A-^3[U56YG8?PV<MLXX5=+_2^,g3U1U]
VN,cJA:U<]5c5+C>X[F;g4X:f+V:ADV.>e^;f:KYHVbLE1Fb8d^RCQ.W(Rc/0ZG@
H[2SL]U0M?5X@[bR]DcY]-FT;PL]405U[=42Y=TXO+@93#KLP5O.\;?KV<3&ZQ^D
TG9C8G/&/e<<aFJ(@6Ug6MBNGLBJ2d)T]_dMX9bfF6):9R,&B.M4?[#<#<9cPM+Q
ZB=N]dD3L+YFDN;?I6+IHUH1UE/>V0Y#N094MNK\_U5d6,5[g@BWTL1_1I3+JQ1f
2e6OPM]Z=]?XC8C]e9:>IE,e0//ZgPdINO7W8D?<[&<J2/I;RHb7TX:[/_PPM[)[
<13FQLf(718IaI5^]R]DI@fe1IH\^HTX^_a;G46#BUI/fcH+XJL>)IbMIYAd@BO9
IR4MR7:be#0:&MZG.-ed#.K&BLe^^A3a9I1_)c,9V]gRB=#5f]UTQGZPF=aP_dVY
gHQ@)bZQa47/5;DQK&9BG;+_4ec8g2@cY2ND[;&9S9K5L4R+4TV9A=3KUgC;Q\)f
K2AgeK&W1U4OJ>X2XH2,aA[6cZOZgP0FRFFL,4)1PH0EGKPHDD8H4L#Vf,H\4S6G
Sf?f?22A#P]:,a(J]K81dI-Y5_9OU:bKWAYEPO0f?BeWCAQ92LA<)_[PR>e=X2Yc
^If55&ALMb+X.U2MPJGeA2\^C;_Q:=)#Q@:+FA\,UURX6Q_<:^7\;;C;KK<\)UGV
V15XK(7EGN?NgYV+1S<]K+BT_W.-TQH@0[/)\;LAI@[8e,ZM@S/C@G=4G;(=<Za>
,]DDe8dg@SFC_+-,>N<.7Q<79[(2MdJI17WZOGIO8:(CR^Q0.6\[?TfW>@+6QZ.0
d-NXD4G#gL4bC<H434@G)69OLe8.,QKNLY]3.AF\6BY_LK7J:1VDOJPYN&X[(L]&
<O2?DdVDTJJ^Yb)?ZT1GUb(M.;SH<TQ)^4@M5dg,DFX?9=c7g2fUc:/LF<?X]C)\
FZ8_\^CM9Z7P:;47\;T;X.EMM<dBcU+#B_:@48PB\Gf[Wa8.ZS:aH[IM];NA7dBU
=2,K?fW/d=I7cK<B@N_1#\9:a&SX;2.#NC9Ed3BZgF9agaA5:-Aab2GIJ@S\5K@W
@)1e2aUPIK=b[Qf9>G;)<,1,CG]AMF02eDIP:8-@3f[F>L2=GYVL4GD^BMO&YU_]
dO;CKfT\U,FbK4:Q#-KT(3PD,.MQPE\Ic#,b+,Ud,@_Y^2ERQ_D@.WeA8^9MS42a
Y?aMG_51_7@H_/+3a@9FJA949@Qg(f-a\2=dM,BMJ_J^9^c62DG&1H3VTA.6]W1^
A=K#=6E01S:CS.2#T,9?M6fW^V?^6g<)W2gSYLQFg.IF-FQSKH_,O(+.U68^Z+#4
>C6/+6K^OYbf5P+W-\BCJ,P]:IHC#d>Ca?6f;J_HVE>,O=CQbV;)UL9??+&?O0UJ
/aWEB]I?b)ZIN:-:1gbH(Qf7;_]1?+5#/BL^FQLTD.R7(0V4/4Y1L.,6J<1S2+F.
T8OfgQfGT(e<&S3NcJ6D98X0IgLAI:OP7Qb09E25;0;DK#N@1>05CdcQCI^S#J)F
^(.P6B7VTU&T@Hf?35U5V&1BF.+SQ3C4)F\B/\U&-SJ]Q6-OOL=I<=]0OL>YM[C(
P>J2Y3K@3Kg6CA5,>EZQZd-TMIAc^C)5\N\+e8DA<d<Yf<N^E(\(f)BG.DWQ@A-2
gL-LZVBG6@EH0)F31N]5AT?EL2R3JN8Wf@UJ:G\+FX<&_dcf7&AY8@cO0O1Da5Hf
:S;2/0EOSGc485VSA=7MbS?_>&V\(SdMaNZ[59P,e&_4HR_:G+O3E4X9]\(F2e-#
6Q,D4RTOI.()&D2c\[/H-=Q-)<F+1T-LCGf[;\Sb&b&;2KSZc7:eQdPB@g-ZGYDI
(/6CWTVUc#c[7,JE0:HYY7KR\^IEa9VP<XdX3KD4:W80<SKd\/e>8e3a5N7D692a
ZBI2Yg6-JWF5[G[a+=)OPb3\S+QV^eET4IPZ4DN#fKIM;fDaZI8/#L=DVC8/EC90
=<1Y;+XTa/YZMIE@7/aS>#H^]Sd5cXL,d9;dCE@42F,?U)V5[A7B/FJfX;;7@_3L
M?c7C#2Xd.FKUDTKI#@K+LVNZ<B&]@cFTE2>WFK3[X^c)UIOYW9\AA<S]fFR_1EI
LG_7BK:3f4UW7AcFUMI+LNXSG]Pa259f]RU@,3)E32NeRI+2>4EKXc\L?15P66#?
O&Xb>@1P5W;<P<T\5,/BgR[c5_KYf6[@Q\+#5BJYZGI(7e0DOZ+](\fdPVM;Y0.(
2OS>[73W4DU&MM+]DLV.:>9^]JaTW6eB\\aUQ-8>YE3&1E\DP3CBA&J&XWEY1eC,
R-==UPFDdV&&T5Q?bZG.96OZ3G=[&2\8B;JXRbaO@;a_Zf_9abHd8c&g#72PW(DX
58C,T4)[WXcCSeTU_C#@)[K7,cY5#HD?F8LVAAP5?Kf]QO<XEU7_L2QS21U4@-DT
4>@X)FIZ.#Kda:[ZME)JdOK\4Y).MP^RfIaOcdH]Og&#:F:gc5LUEY3U)M7PBaUE
COf]7NI9a7WF>gZM0X)L95S@[1\/=PaC+IOY9_Rb3[^aS?TRJOVPKRb9CbHd1fJK
<+K6V_TE<B\>SA?2/0Je-(XC2_?gULaW8eB#(&13_UF&U5\R+f#8?V94g0(Ua9)_
g>:=Y^XF7Tcd;TN(&T)1/(PU)GLMbQ\5)IF)[.5>ZT0Va+QT]??Rg_RYZfg<Z0HS
.TZ>5,@<@X->](K6D-VOD)5g\J>\Ed?X2VR\4aPA=(dFZ<7IOb[)CZ2922UG<ZI_
\K]#@OS5B1S+<CdYd/2&RGIe\Q86WQ\K][]]c5:NPP8.0ZO<RJP?2^+^\Zg]&eWd
U\)/MZbR.M4KWA+_0@:Z7-^IR4.B0EZWIVZ/RNZ7#=6](\K\/dfbbdUX9>,e(M7;
T#<ABX^bXT_X=4</bL.YQRe>@\=AI+/05H6.XN^c5U@c.[9CSVAG^f^C=XO7e?.X
[Z7]_R4<B4^8aR+@B[eX(cBH0J=E51F0JZ4VfH3NFL/^?</,6>g\Od?4+Qc(K_:G
/D?>dRUG/5M=HO2cU,)?RQA.0R?dYQ02BE4g7gA<MgD_T),O+.YG()A>bT^aQR0N
aYf7;cEX#cb)C-8:Jb^9f3N86_^+J:CK=B.-XG@0?AS<NOgZ&IHK++LI^P784];1
:=g]^gVDdgBS8YSN[RbT0P@CXR(WeY=b4;Rg01c3GMO0Q1f)Xb;/-^QZL/&X,0aZ
f?2I^X-W0D?Y[0/J,OIOED1]U,=bSe<<f633:Ba=f6@8Q^eGSZ3Rb1^8PB&(A]S5
+B_<L<@[bg=d+LIB3#eIH=G3IKM^.K)HBAR>,9fBAOKB:VY(Ud\E8^^MRTYMc)8S
WYUNM+)VM1C(#@Tb_VF2B9&\7\9S2:>g?XYf)B,3COIIR@)EO\a41,Z,eO9SLbD\
V@-W[;6YJ&N;:e-9##Q.KP[)4Ef[a+I/8]V\QJ@.GH95R)C_#B5/Y?(@;[62ObD3
Z@F.U)E+:<KF?I;06(cb=I_dVYJKEAY].A.9W0DXf83N?PQTV&26^bE:^f@(&UaD
9LgMCU^1g:O.&-5O,JXPb-TS1^LWV+,#TNJ36D,;ZQOP+B.(Ve_(.;ZH80AKII_D
GA58aYFRIE8^[Zb)MYc2RW28Fc6O.X]O?8S)DDZS[PaE<dI(7LJU12+AY_9L@8)a
L=I;Ob#CO3-VRF&f-Q/17+ER-\]QXSUJNK[<N8#N-4MEN6T34S6#VYQ@&3gA4XYZ
GQ4&IfXg=/]QCYRI8\S\PdOSN(-R@&>.7LM&O#DG=cE\V46.(f>E98\KH_=5?Eb@
LICe[PCD20/9,)=H[+La7I.6Y8.dffSeBJe>,66e97BQf\b\.7^b3<9M@?L?L\F2
D5+Gbd?G/BaQPV>d5eQ9/F6e\IG]bB<>--BLT=SJ@=<59ZTbaKbF75L>0O4U799e
GR]33I\:3>1EbZeb6;90VIJHBF7a[#;a0LWQ_5FO9NPRVAfQ2LA#?0+<=SYHD_GD
b?5/>-O;E3^=1ZH+JZ8gP)O:P/KdZ_2QMYDLAY10I5bA#EBJbMVQS:6M.ZPdQC3Q
CNP2=[[H.4db2[SJAKFAH9/:Z<8##>ABY>^50LUZ;PDRRGT&@-^?f-<1\;G80)=U
0L:C&WJ=?==b1Z7>GZ.:QcgdSPBVOH>3,&(;IQ&0YZ9-S^0B,b-XWF>\WFedHg44
IZB<:,LWU[8Z4RdR^OEB:/>MVAYVKDA7:8dfgS+fJ=R,_XNE39:3^B9f4S#+K364
CI&4bR#X?5KI&QY;,],>C02&Ed(N^a,,Q8=CBc_+_MB@^R/Z^94RZR647J4?[TAY
AC]cM+,6>4YG9I)Q_[W46,;=ZK60d_gPGMCDTZJ>RT]4,aB;Y5VOM;5M]-[/G_;,
4X>#1=/cT(U4Yc3W<DUM>42W^gOHZ3W5\Q&+#N<46BBDVQ]W9WR5HJd?[-1A/C\U
-2A.Q;_TU^)-IM_fUS4dLEYSA[cZFGC0&L@C8R7f.c-@FaX(/g.&?Y5]8?;dTD_/
8#YeH&SO2TRDWQ#aDB^URPXFND[>&-NGVfB\GH7_[G)Hc@PVf(30c9+;LG8+CLDU
EC4TESST8?FN?E@DU_Rf)1e-K/PHA]V;I=>9&2(O>I9)EVQZN9+cSB3<9;;9K>G.
X11+@AbDMRH28^W#EV]@b@=RF>;/WLcT2_45T>/<]bU(dKb(MOTA3B4DZ[OcgbRI
GAS.1Wg\e^e2CZQ_/;cL#UMB;e)P]Ef>=9IDYKQ=B,<eE5W0c7<#fcIQ(WFYcfJ7
##Y=(O2>[?96B=+Y^+8dU)U_;C+2&SA]7>]4Q6;<a]);2eUa>@A\C5L1F4N(T[RU
E<=Q7B@gLJdCP&C7D,#1DSS@?3.9K_U]##AbL4K?TO6#PEc(L8B6RCJ6fD@M&_2)
A)(;c_F0GA>_^=d-9=+/aPC(_\22d)7/#O/ga@P6,cFc-:IE=6Q5#0#/J\d:a#)9
dee6R9]1&e5OaDZYaQO,AT)cE.&^Sg#Q1fA:OC]6E7##-=UV<=W/K=P.]D)&UP57
eI7-dPb>C)Q?OWgCU4Q[QN_3;a=d0MKACAc[,d(a-(90V9D9M]]C-_2Q(^(QTERS
XV1fK2Lg<MK0:7[J9=Q2]1Mf>U(LdFa0BdC+Y-L:U+e+68BK<R(.GN4WfP5S_Rb9
?T#ZXZP\X?X8K98I<3>3P2N;_=@))1/6(d5^bC7X;WSNR,Aa.@2TB:AP?TQGVD>:
D9]f>I57JVL<Fg//;D(K1=AAgO)R9(<#g\U5LgHZU@cVSZaY=0cL)7X.9Z9V<6-B
K]_;/c)>=Ia;XKRUEb:<;1ZAZdSJ:HF<\BPK=#?][3WJZ0Y2&^&&CTGQg2DU=A\/
)]CZ@YYAN0EH>EL:@]OG_K-1G00=UK14U6@YVF\TXU9A/Jg>_ZVa_7TS_[2D206L
>3([,>\Z_.U8ID,dVX;5g\-4@ZOe+dDXNC[YbY[.3R6<c=2?SX7bAJW=I4+N4^dM
U[KE;/DUXB30daDD,3L[99E[TG(S3TA5W^GJ7\IT(ZV8FK;MReUD7<X5Y:4^PX3e
4\H/Q1#e&;df@U3KK9bdV1EQ.)4O5X/N[LM0+XEPE<=HE,Zc\0J+ZSJA\5/>C1/#
2@D4L/_OdVb.;@ObPgZ=P=g5-/9B,UOgZ<8g276\R81P#@X<4&_VVDSdX4J;:0YD
S>.DaSdZA.LEF-\AIH1dUfS-;b_Z<[G1,4TM(EC02D&VJfN/5+E7O4Gd#PQa5#I9
(7:R1QfFU4/-5ZLDS2?=Y]3IM;K-;IGZ\M;9bX[H<2N4/LWZ&D3JKOfSOIC0RBMZ
2>YQDNJ9[=/\;/8)N[H-UH5@.Pb^75DSM_ZdbeBJNH=IeWI9NNT^1R).[DaH)F]B
_6(87fYEYfIFc8^LYPb->.VgZf;Y7PaIULY.g^D3685VaZXC=>1U-KGK9UedCT0I
U&(^HF<)HPJ7]7a0G.RV]XIL#aM>83g@J@WgOeS6c#1G-H\^GQ8\R1gaXcEQ&,)\
5#(Q3[IFL0>M#&9fS+9A@.C:?A7&g,9N-U62OVGgH8JUNNP=>ab+Q0@5W+AFY69+
W//:A=70?:?a,a2#YA5#ZWGT+RdCJePBI-(PF-D8X:(U^2A5VS.2\JM?I56,1)2;
17g>gd)a_4NcaM#c6AMBEZH:X<I5E#?A&K4XWDBNO2O(8VMU<,+J\-VC@&,&+E>U
9-ZQ_&RDfMZQG@:5E:V#I?=)fKcM]23\JM69&E\J+=<b9@.b/FBZTN5dY^\[185,
4[0;0AMWRKC//L1-HD9Z@EbMF0<WN?[BZDWI_O7H6I0X]c\V+\_&;9f==;+T5+g@
(VD1\VWO:XAX4SX.&-+7TPDV7:_Qb:\(CB2#S&@YC^>JMY\&=DONK.8GI/DK=TY>
JM.d#E&9N-_8R/CP^eGGXNab_F+0G?,2V(c@K4L?<?)e)cVJJ<UYfdcb/#GZ#(^1
5DKf[F:HDS=df9E_e,6aYJDJXTN3>S9^<1<)9>XIYMH,Q0/CJa6A=QNeXTWK+(\=
Z_2/@\PgH\=5?gQL[?G34PHZF&=(HAdJ)S,G2.HY@JPFF-IG&6Y0-6a(8KG1\_@O
0ZWN(9G9WZM.db<S[_R1Pc:ZTd.eNN9XB2>W)dg+CJC^LV.ZZBb1dC#ORLN\e]6X
B0(C&48=+>L\/+<C:40<3)HU1+M^D876+6RLJgJVT09;,0c#]LFTY>KC:6U[2Z3d
J0W)OIAX<2=@;Sc.a:Rd[S4[??80F2]&MdS4^01ZQD5/3<_:Z(3]SaQB\8[&EbPe
U21]9,ebQ>IMKgWI?YGb(\UO@,^W?9MAS&N/f1Be1VDU1fDP1W02e)H]]NVEZM1&
2b[-792M(:6O]S=HURSY,O@UGgA:X&aeA0G?9<7L<+T[D;CcT80ecbYR#91\aT#R
HagX[-G:g-e[KcbD93O,JSC]W&4F#g(L+JdM(&1O^Ye1P_MXB:IT7T?MW/H6gMYF
\FM)?H:-#0R8=HafY<6R>g.Fa\SR+VR)-bd1JUBC76SF9Z2AGWcW?4YFZ?0\[K7;
0O@9MYg^WTgeI;U=+[Y>&faaY#Y.L.H7202BKE28ZMR4F=W(L6@e#-U.C6SXGG2+
beQ[bKRYWQeaLN6G#@/Y+fA5@360,@&_fdZWc:<ICY\LVWGU9Fd]ObgHU#a,;&_H
=,D(eDZY93CK^IS1)DObB]daM?ESJ&Q&&??cD[SdR/._X2AL/>,8J5f5VG[]\16[
01Q(^-P(?e3&/HfZY^a128P:GZ0I<3CQ1K9&(K6eFDW@ZKPCZL:GBUNL[Q4eb]-G
F.1HRSN@W.?3JH.b?H4^7;0V/^c+E9bD7_?@a<OD)>2+@4dc-1^.Ef[,C<AS(H:]
g;);2,SOV]EGWY7bC9IHCQ?@L.&9#Q89JQ6>9Y31f@ZYa;69@6;AJP(gMA;.@U.Q
-DXD3_0V)\AZ8d-<#@4Vd8cQL,48079R0dE1[@RYKf&@P=Q,LY-a[GL<=2XJNKO[
Z3b5GO@9_Z/Jf)\7JHA<LV4Sbc8BN&>@ebYT(cVeDP^S(]1H,PcD[SS-6H5@__I;
[?#??D1S\<g4BTM0ReUaPVH5./2ZL_QA.X6#0IG[^@O5BWZC6P/ZU7C+LKQ[1J(R
D@4_VHgTFf)V1JT^Z,])S:W[@?(J5gQId##Kb->Z,=\XL,1DfG(JZ+1ee4E0./37
#DD&BP1cZ^O(/6F#B<LUSXf<3EBHWf4fQ\NA-5Hf8?PP[S4,@K50Z=HCLA=d/IQX
0,)L1/3?)a[1Rc(XXB/,2OS4aYAA1ND#LZJ\1<.=W(b)=c>[dGM_QT#5T@C?6b?.
dW5-,H^:cdY[MGIfgZA.Od(&ac)dcA;\CJD7:E[d98C@F[G1EaMPeBWAH;GKB<2E
b]X[^AG5)XD8.C>1LeWc=7]4B3K&V8e94gFV+VN9I_Z&IU#&AAZ9&4[WS,T=9@a#
FS?QPS,aW:P4T33NXgg_HJ+O+e1[f5Z9f/P;&D\/dU(<6F?<9([A/I6C)UD\XTeK
4AX3AZ(_I1K\]32cK3>f6[D]^F=7N#2X<;9>+\9R.IPK.B5g>5)5(a<^1]dNFbe?
b(-+\^a7;NHS>6f7]F4MaBNH-Kb.;GWDaK3J(OcV(:,0M^0WE3(Ob)S\PROR?#:-
@#T94R,Q/E\:8T4PP5J9A2N@4?B6fJ/C9=I4e#)==3C(T.FJ4d83STU78VdDO0Xe
:WN:]OBYQKQDW.N>[HE)F0^De<F2]aLcEeLVaV+J:1T[HA73.UAd=8SOKa1L+0)[
cLTbTY.15BLL750NJ<L7U)(e9f&aEU_+@-S5cFYbB.FDP:?8,9eWQ6W8/bPVVAK9
2c[RP5I4?+]5#OMaPG_55K0HP.,>)gW:8(U[]BI/BGRAA>)<[/FGOfRF6D[R3/D_
gCFI1c5fZ/28MGdMT7E]7gNKXI4c9<>/eNX^e-&H_]g_0N,MD(Hb1Q0W0\K&M6+M
1c-?TSPP:X-bAZG[1[:2T>:G7OF,JIP0F1SRNeY^If:&+;Q=]_:FFB-;L:C@7VDN
@dbUT&WgL6)CWKJ:c\^^?CX?5XI+Td2#\gf@JU.ML[<N,L^Jg3=]5XbHYMWG7^_a
6S92LXE<57d8\AWS>:3GK)8LQac5Hb-IeTN80Y6F/;9E1/YC8OAWENS;=#R?dgL3
SV9=g^KGI:1FXCTV3CS\dA29_M@1M)&R_f=0f8D47-B>U_6QIcCDE8D@B6:CT0RS
M:g0cK@2?<](QP=TN(QE#G)2.?^B^:Kd(YE.V^6[g/1<6[C8.3>gIg9M@ID5=^dQ
;T[O3C)SWgSe6(cXF?.>CfAH:(bB-0a1XEXK-f1ELL(aA4)H4W@RN\eRX1Q-DK@]
/7GXELWg,Id+G,,VJ#N?WR2AgTIX(Mc@ERgcG/gSFL]aI-+Q2Z8QO8JON9AUd^JD
L:NU8LC)Ve_,L<SeEQ:begXPEI].b<1G/=3e_[4/H4DC2HC_@142ZMI/,dWNDK=]
TK@?@.e-\3fDK&U(BK^>DGLZZ(]9+?(Q_]6CWcNCKe2#3e-5Xc#R7f+gc4][U_V0
c-&::Q8JQ:.\.)fV&9HdR=]X8Y)TA_XKIc2G5[YG6b\/ZJ^Xf<?:f=-F:#=AK.Eb
MW53FC&R^/+2672XBUCMfa:<R,&P0VL_S8gMZ?CTUG=d(gL?30]7H9-LA:H/3S5M
8ET=6+2Q21Y>]bV)X@gN,\@_S6H&)T;8:,UJIK=^VEQ5YbH#3UUHd/>=6d09]cF4
b2T1#:?/IM7,L>S]8=Cb8PEdEgAQPd^_<PO0G+\eO_5g+\0M<&f0:?LB-N8PSGQQ
aBAJ+PGAD([,47(,K=CZ_=L)S75-[YJA&_DHb)Ced4UVJU#(LXT&F0]G+HJZ@e+;
a)T>.<e-:cR7B4>.Qe-\^A?\df51:CTTDF^b6W=SfN^XFX14:LP:,7U#\WR1O>SP
c?2eYeZ.RZ[\4B[]cfLGgWgUMTXWVDWZ6D8G>D@G78F6+2,MFaWPZA13XBU8/T@W
W:;I)<C<E)N.Z(KcN7fdM3RUc(@\+U^T,(.3deK(deP5fJN\ePMUWd@I-,f1cT#X
[.[_)JTc=GZ)+UGeGIb//-9YFb;B9DXK7a+eTXNJT-9R#D47[^:6ZZ82?RZCC6>V
bOe5)2/dQ?5]#Mb5f0G,<f_S\b.P^RQbaDY7SVI2-bFQ<0S39\#K.][d&^DV/U,d
SW-OE?AU,-aB-6a^Z.RXKF84N#?.V7R+Z6_ggHBEa#dZ7+W\QE>W-e6X#)I:PT@g
[,0V/MC:^:S&PG1B=fKGIN.5gNR3]P[<d/d(b[dHQG#OE5(>YJc@^2PgC.<e^EY1
K&&I\<N[H)eTa/S.278b;9SKWM(e(BE&611J=[;6XXUJ9MB-^;1W8Z0dRaD./DZ^
X5N#V>,c(c^EGfD/[]CBdIIaEP]Bc=?f9C_+e2:CX4A&6[H8D:e#.#4PY\f5g3]b
O:[I]@VTb]9[_UT9A7VZ4&,KR,)&-<<5eCPN5R_@#QafBHY8T7MU>K7E.Z_JJ4;_
N>IR>EOUc5<-+N(GAe5O#C+&:,P]OOCKI6bFX#@L#KT,AeP9dS;XHDC2,#;6:X<c
L8^^Y;Baa.GNV0L5L#[?^MI;dSTUE72@+06,5+JDI@bDadCF5A]\LU:6N;D]/dHY
6+J:a(V\9.^Q?\ZL4^f;WI&LJ:P\5I6)77Z<,;e?[A)Ag/(;J7,G0-0UI1N0>eBa
S@@0ADe[A9&3V/@<ZE,,E[gDE+6d,J@&HN0AeUX<.UYdg40GGe2bZLFRf4aKc>)X
I/E[@/T<[A_]AKZW)W/\>LTQY?dCZ=/R728W^4^fD)9/QZa9^8dVO^-J[H9MCV9E
P+>(1BKg-LZYTb-5c@O5DNW-S<B4Z]8\PCE>aL,:)YQ)-=E0/81+BQB8MFC(FC]@
M0D)GWZRE#4JK4]5ZY25/\O)?ge#<YBK5M]).Z1?6@]1Y3+=c6QTF6GUA\-YB[2O
B4Ib<@L=\JBB,7Q@[d^<ZXO#R_,4a\Nf^K@AU.P-_aba04G5Q?J3NX@FNN-Ug(Q;
@ED\^/=LfIX/G-X8)g?OIU]Z=?G>,>6YD]5TCDdE?0^0Q>ZH_7JUXP(HIV<#7&\O
JBe_SO#IAWHfV_)LM]A>>,?I5#Q#FSL<\^LdXNP(E@6,9DPQ2bS#Qd75(C9FG3-S
dN&L6>b<TPR_FRIGW\+@P&Q9_?Y\^LVM<V-8C7gI+M.0#gc<[;(;0ZGP\:UF?#Y+
ef;A1ESU7(.Jg8d@8AAHF\D\IOZ[c9K#c,((_8SS4cE7c(cYX&1HGO8V[@e19Ra+
6@dafATU7P\30MC,[PRW1Qe#@?G7O4:JRDX:R?X[Z#0+BfSTe^_W@#=U@CN,0I4d
aJT#NOVQPHEF^]NUeLQP[EgV3D&9HcX)\N+@b:/PE5FS2Z(Y;8/c0DMdUF8IQ7HK
KNXc5)NE88d?=9QVO@J^&0[?P@[C@4^I?;Q=(FY6]Vf&Zf8.3;b7@WXf0Be6E]+a
Ub:Q6JbYGaV:M8W7Y6,X-Y5Q&3(a#V(5XK6=[AWWX8,e.b-XH@d6VT8MF6RLV8R,
5RQGVb?2GY+Uc&5NIEb/_>(^TEGK]S3M1VB6Rg4Zfbd,dR=?XO=U1[G7G5P9WTK;
VAZFXQ]_81ZKO@JHa9B=Q>f1D[,gL_S)G3g1Ggd_\0dL&V[MD<#cMG/:/EX_FB2^
GUO_D?PPZFB(&\+edZK<Y=MX;<SaQ+<\):\]OaT93P3\#UJ\fX?KX,+\C7QCM4H<
<LYFZCOO_T6BbF\[^;;E1.[\c<W9BVUQfDaKU6)R5\VHZA/3D6M3CW&GML>5b+/B
K>OA/b\Q;eAZT-8W9PZIZ,@\gFQVYC?L<Sg\2\PfJd_8F);N]cb9@,:W-g9&\_QF
,@Q6MJbD#7]4VX0AVOGD4:\)XNT#.#3W)A)+9M6aQPSE1Y_8Z/=X:>=WX(Cdc^(7
IR[gb5d(A88IH?L#6P.+.F06,aFM@c\2[O+N;T]G[+UG:7@U,.eL8cDH<NQ=-A)>
VYc,YFV7eZ[L@?CD?EgEK=#0GTd4(Dd.4O#)=#0D+cO8]Pc5QG9aRR^@=+DJbGI0
5^1#+&J(W<NedL2d;eOc>g)0T;X8C\<@87:_;NIgB@J2\IHDDZ2V>M.W96S7:?3B
eb=4TZNHEEO=?BNRF#5R_LAJ95d=b=],]MQY\1/&=8/-a;?ZfNbW7AY-ge^P+XQ]
=d+JJS\SH1#+ddL>L5.\Z6C?-F2F.0+;,b>7Q<B2L8<IA.PUAEZ;;B)C(9&c1J[0
M]Fae,G?.WP[W4PL2C2K2@4^a/<:.T;)25FK.I=YX?,7/?DVf=RYg1gUZ)8S=2fS
=VP[/^V95ecBUD6,QO2D@.E.LKe;Ve-&1P?09C-C>QSB0bVd^]D8)Zc(M@V7?NLc
Qg[6W2E-N9Wcb^WdVJLGdfJ+UU<DZ=NQUd-@f+9:^05c[[?)<H?6(Y?>GOeY<EA#
d;9<=bbKVX&bN).bIC_?PeE057d=AP_\B8UBU?:A(>.YO<K4V5Z=)NDQ_7;CT@Je
]#I5WaP/0bE?fYE^/[QMBIKQ9=:O5I>?UBLFR.LdNFfO_)267U4_G.XE1PY37cdK
?4XSHa4=NF:Q:>/FKMgc^ED[/YBSWYX.]LUf&<3Y=CV[YC9gJDS.KaVG6O3e)Q\Q
?HC3E4P@^B>PIOPF5C7I3CT44.;7GBHXM_,<=6/UJ3)R&P:1aP:?G#VEE-S/>I7]
F8dc)3_I#,#dI4P_;AWd\[LD]2=eSbeZYg8QTadGN>E&<1a:Hd=7AX<Vc<>e0P^]
JNFJUM;DgC8a1L3L:Oa\7#.XbJ?OfJHHYLW((2]U:GKV0BgG5fX0,[<XPBc9#7V0
,RYV;#4T?5;e]?4]c,<,:@dK/c48\PBd[/Qb8VI/PIB>XP?HRLLQ:,+[=;Lgb^;\
NA@Z?_Yf1=1#;[QBF,g(UE3?RKSd.X1]Z9e[^-R9g52bbb@dC^WXOG61+>?=;HRR
9=+=GXDQ8[.Z?;XbFcEER^:DA&9IL>aFe6&CDag;df.UZY@+[dbT?0+cdY=)4Qd]
]Yg2bK,7/D._Sa#^EH+(Q?]N+XH[BEFbc]dZHgbE,R=TIcPCRUgB_1b8IW6b1gJ&
\(HSMEa.XD(EU#de2BS?DEBfT5BQR#Pgd?P+#787SCdI^\-1>K</ZHF2GLW(2;50
ULKYNXO?b?LDc[@:>WdEHb_A#/@0bS.^5JT@B>bd9=L5YYKGg^#<090\#4d:5XNV
8g,:dUMd4Y=C9WCDDO];)@G/5\dbb].RZ75E?-7&Za;X?O=0d#,6^)P29_RcbafW
M0g,C3c:RBWE5@Jg]GYba,;gT00>f.3.DUgY2c>cb;BFMMYI]X^f]Q@cC#A_#/fX
.GIDPNJ0GZ_PB<,#W,Q<@NM[B(#f1.<VD]b#MJF?GXCa#4Q<)D=NbgF-Z@aT@DWL
(K6+&<G-b6,2ZQ6@V)KR+W@T1C#e:-YSRf9HQeD#I4^/Q;/-8c.ZO=dYKKTRcEP(
dXX)5faD56:SCB+DM3#\(8L]TbNgQD7<;g)4a=35QYK@7V;@:9\P+S1G3=<J#454
NK9&AURID-NG=+QR-a(b>[eRT.,4C]FPbf,O(L1<Wa.H,(5?KA4R3/7DDVPFOV;4
4.FVC@RD.[GgKWY@:=QT;^=d_7.G7?#>B,a2JD3Ce[RQSPM1:W)5=459YT2;&H@+
aaYS6<XUI;P3&eSI0LL04bKd.>I2f?\cc5&)LK\#DL=Pb0CdUKN>Y\^+.[aU#R81
F=ZA4GMCT3<\gfCf)E<:#1MVaD<JbTHN39^+>@a9=R4G(W-d&3-e_(/Vf-9Id(IO
CF+f\;]ZH)/6D2SW=G5HYKe:QbB&=/:BU05HAcB72fCFf;<#fddI9,FFd8VcVYPE
>OaJD2EOdFdG7>?G12AH7M4G?GdfW(1+&52B)D01bN-/95&G.@fTP;DQGN)6S[KJ
2OcI[J^2<J+NW7H7Kf4MM?GYg1I/>LfP\63Y2ZKdf?LWGIWF;EcZ7U&b#L7D+F/0
]/MN:M7gXJY/#ef\_SaLf=Veca79S-V,VVM:+Hf:ERce@IYX3)7SRP\WWOJVW8>g
NE8#c[<M52.IN/IR3L[8R7d,/^9C>U[]7Q41\C53,aAgRZ).>Q[9>X.M:DH^,8ec
)H[f2P3#-OA:a[H]8Fc0X2-@aJM:0dM4d,[,&Qf[KVFNBa../F3>QZ?UB5Ea&1ED
YP:S+-.aU;-UNU6D&B3W/#?P.LD1PF:PAD-.0>?Tea5?4_WJ)fcdb4Zd0^\2TE?W
7-I;BJBVKH&+HYO-\]gcS^0<X9M=FgY/>7Q0AW[OLa>?R8O(e/ZVKU7>+@T(UF)1
RUL2)]cCB&b,T7;L.J2)XeO+SL/VG]6(#:FaYH#.70<W77Ad;V\]XZH2Y/HJQ9bI
H/VPA/VfGDB9a]XC#H\#Og.L;<:LPJZ16?V&(4?<cZEFS5T>TLNf(+0YVaCBXWV-
7@;RQC,O2LB:^XMC-Kd@M9CPf_PT]eP<?\_M(2\)UB+._TaY^0M+@2CHTc[0JV32
;;&O]#P.-=b->fG-3:E\;>CKAg]/U)QYK1S2-ZW-+95WV0M=F7VZf;e;Q/fc-&V0
(0=/5U9:IeNdF=e>DfH.V(c]6X<G[2UOcZR9AA7aY_a6?Ka>_;>:e#G@K[fOJ7]Q
V30a2P9XOPc\1+K):^?M9<fMXGEZSDb?@)MN8^<8D):GX==,g?Sd6T\V:BE&&0,Q
RWSL?2>b+8.W8gR;#]@N4-]>=/8O<Pbf]a_W-&HVIe)SgE8(62Y.G:Yg<5cL.>RO
g-(JF-f@AGYd41;SAK6K,Y@=\Pg\<]V)&#B^0)]WFPXMa[SGG=(/C?HgHT^;N9;-
>2))Ye+KI,@:2@[U(caB-<WKRPLD09\^:]GZME@@&PD+R)OGbWgX>4_:c-+c_A,+
c\A;bVc:L64.Vg373-e2^V^S8TXOa9X;E7K]27^Y^PQV.S[ScKFUD/<P.ZQc\1EQ
BeE3K?YB.VVg@92Y9+D4(X<?38MTPRF41=U+II:>NSFXQ=1:S(A@Z3?&\D[7a(@H
JW&:;3DEc[B,V0#KK=aTE.28(,M4=1\gK24_QOJE^OA](S9a90MY):1^>-b,gPIU
Id&]aOeAbc]>YN61A];.<R^W\3M6@R3L(+e8?5SK(3N<c>MQU)g(&V-?);L;0WW-
F89QX.b&Z-GYIGC&Q-:dbGVeAC@,S><K6BH[a489eQ>48SQFZ6R0_V2gKb=<KJ_=
\3E\\F]NbgS>I_A=/OL2(<[L.aHY413RZH9)0\=64fF2)TW,SdT2f-e/GECJ:fW]
^[(_C0(eILTP0WZ^@c6MTUR7.8PKaMJ.A0dXT7A64S9V/;TAbQ,bGc]G\_@CN[:X
LW[;CYceP4MeY<E/ZJG(N_7g#KFP)6f_32L.@bPe#\:A+765-Q[=d?Z;H(ULRPJH
HQN9I/R#@0H1gg3cZ4M_&_)ME6H^W&UN@GOO8bA/?[VGU4fAf,^.2=M?e-\OPL][
FWc:)UN3Y:67/I23?8GcPH.VJ:-O.V@P.?EH/f8F/MQAE\]GRDE.1Bf^bU^PRP)^
V1\4T@1X@DR=N:(>CeHgGVX4[\)\C<ZBfOT;7b.O-W+\eEG;M)7NUL)P//5Z^T@e
]4U=a;MF,];)Beb-F=@(FeO2+K;HHPgQZU6;N.H#b^F;@1.\FK9D168.#LbYF,QG
<OUH(d4:[Kc;#P10P6c@9?@3TW40-9b9eNP47DAbBN?YJ[PL@TcNMI6,MBRJ],e-
GOgI4B89Y?T^2)cLdXC:^K1NQ1)MZMR73ZgL5J3^Md<2Aa&<DO-g@_9(EL8c&RAG
:=-<KVZ-3@1+YS+T_fB.88H<X[G)>_T6#)bLA^I7(88_\XQN[RPQ2;1[.F[6947B
=;O5<UQLTW]_,CD+5/J/9-dcU_HPGUb[-&9BgNgPcY\YA;9N^_@#N=/QgU845?=X
WQ06JC4YB,V8(5T4G5.OB:<:=<F?cM7X9eIID.TVDe8;T&K=]4.T>a>?g..5RG(B
[>[FCIHeA4ae^Q84&2SEe4AfQX1>/2K+8>TXG<>4C58;RbC.V1PL4\.OX^g<G,HW
<[:Ab\I7D^7IF-QGQ&)SCS,<4.GUS.4)17PML3><Yca++/NeE/?,FZ5(LQgQM?UE
S,=7L1]dE.V0bQT)IZYggLf+LdAK:;EXG,^gA1XM_I4b#@8.)^M>[g2=Hf+b#:)3
)\+21I_\B1a<5eU0Z@2a:F1T&J@.IF7QJ0/0MLSH:W=73(5>cK&.4KYYTB/6V>^?
FARZ&D+dO<+7)I;.-J+@9Y^V:0K>>-JB\6Y>&[?/[X[D.>_Pa590CdC__]Q7_LfQ
ZPN^C:fYgU)a1aN7Z??/0Z.-Od)HDRHHNDC-BW_U:?#8OC?(L.I6H\[?U@CcRUa7
>#[L):[Tc:;#WYd8>E,IZKD81:3(Ng,^F<E8d:E1,;K./g:;-)B6BC1[@:ag2D3\
:dde67@##ecDe.PK=([5&f6+PMK[)-dd61@.+AfJe>dA@I.?ZH;2d0c:VO<7HG.G
DB;a@b246E[-YUO12NNdTU8\PMfOeXSM1aCM2;[FPAV7V0/SYQBO0fB-/9#,YKT6
Ef;[K)g[[1J/5>[3;=H7&ZXO80+(UK=[6=9Z=SfB(3bE>BN#0IdP1@C2>?>7\CE:
SB3U4HRC?HVQM^5XHK^RQP4E)a-.RT(:b>^2&>8//HT[g\1268GG&6?M?=QcHBF(
-K7WHUX0.M3]5?&X^AFL[]8VJ26d^9.\^X(2.VQXVfSUN(Te&AZDJgM##8^)e1XC
:gAfC_X)BMMUFgD(F\]#=0AM.I(ZAP9cB.Mb>1AeQZ_A-Y;-TbHP>K8E>49QPcS0
3HF8NICf4:7?0),eJ;@LD)O&e<@C51N2/A>&,D>&T[CJ(3<O90gLA09E&\8WaE0#
b8TPa.;F4Rd8&GWD4I&bDGW&RV^CcQeT-;8.eR8HIDC307&(cf4&@>]?BJ2Q3^Hc
3b;bPLe49,e<F?f&&[C0=>>6/].]?T2QJZ3g--OM4K&V+SF-.D;0V3SAT>Y;J:=\
76D4,c;_]8eA=LN<J:_]VYJ<O8P4K/Z5.Og1d@C&M<6)gf.AW+QGaE^)4P^dAF^M
I8XNU1@.dcU+8gL8.GcJF;1_HSe38b+FJ^Y6^WQ:NRRD_>?ZPMD5A3aUD]HdA;WT
ed8A732B<7VO\BV40N\<OXMS?E/&/aCNaZ;,<R\GT=g;Te\-Z84-FL4\Z@?)O6<E
?c(7g1G;(O=J/>[WAP4KN>;R:Ke-X?1)b)X_.8YR;N_YY(1Y12Yfc;>&N#a-SX\(
4@)X@#W+<]?5RCG-3@Nc#0a4@WY#@I-OLVdJW+J:1@<C^[PH\Q.dO_#&S;^R6O#S
Q:[f13FBT2+Q#9-)cO[LC72UeBQd>Q@_E>X/&I7REOZI[ce7&UCD77Y<]0O^Q34W
d.>]L_4+T#bNA;@+;>TcT.TWM\e8EbGQH.\-12C_E4]M)CK8)NS#-317>7RX+cW,
3g1Z;b5GSH;WY02OOTJ4.L2_M\c+3^TdOa.cMG(QY[3EBEgHTHV1bBGI0Pg4W:T8
YcAV7-7JH2;[38eS70N]G1?JU/==R;RXAB5@VNHQ8]\FDPg.GH3/@Hcb].MQd^/U
IT&F^>&L//X<O[7f?<<Hd=<R3]E[?T,bKA&,cFP2Y?=WMRGYeQDA3>0>#ZV/UPAR
^d6=;8<WMV;?PZC#fR[QIY^80W<GT^]P?8Tf&E/7JeSUa)5fV^L3X-b2U2(1_d;N
NQ6;gf;_-I^(9-2V2&d=]A^M@8f=GF8R.>@X,;1,c9;9g#W.b,6bV7BO)ND6M3WY
c-H@2aU]XfKa2V#[.<Ff)QW3CbLH0#0NHCZ,IFfFBcT3_O][&Bc-;RJ[6PeT@e.T
XDc6f?fN-_(5]9+gJRg6?AddVK>@Tg0]Rd&E5XY1BNO7M>TJ1[RV&TYe?7GK\L0F
=?_gOX=2>0+1YI+,7A#W.dUPAQ?cSJ.G\a7XGBSS2KaTO6cNU9bT95\^)+;H&F=_
:\[TFV-0S^#@OIM>[:K:<g2VgeUYCZgY3RI7Y./?M92ID-ZSQZcO0+DK@5.2b>.D
)=^,=cff0[CA&=7?ER435EC<a10+Q<N2faXVQQ1ZcTV6S/TMb[#Ra:BGf3Z3G:.Q
P-).+QVBUPDL_90N9-4YON@V+XWCb7O_Y[I8X6O2Y6T=G@EgT-Q<0+ONe4;11D(<
b((gcOO2e#8-dNcQ&XKX7cPOPc8D-M-^47]K3I=I5M07=]05;U(S;LG9XdgC-6(0
K;Q?I(Z0B:DFLYYDMW^EG.8#TSX@.7;A6D1_7ZcZ0E^4:KDETb566\]2WP#<gC7+
RF:KcV+(d9,a@A#I@I=f7XR-JfFYYY_;K>O:X(6>HFNM>@5X3LEQ)g\=N@TPU7Cb
)-e,3C0B]UIF<\3NDBH0@3LGg1UeOXSf)(1fdS=E/33B;6(#?<7Cea6b3D.bG+]0
=]OCHJK8FAB=(]WIT70S<R4V5)EY6DK\b1\FYZL>U&ZXO\;f,/&PB4U5f:4);8;8
Q:g]\M/JZ^K?:>J[;LZFU#I0PJFGT_)W2;8@ZWU<Jad&W@M3WXF7OfHRTJScDWf<
:;D=&_=@9PW9>[UT9&LYCg\,/NXe2>_VcA3eM(-eR1f,&JCcS<0f2H;;ID2Ef0]Y
H)/P,W@WWaBXLI<dH,;,Q9DV?FRB^4=XI,VZO;;<)=XA8?QIRS)D?cbbW?e\6b;c
^aV65#c4RB@a-.Z87VAX1J7fbSGHKb.YQ,QcF9.4E2^-Sg&A_P4,^1DPDd0H-P6,
[P)cR317]72I2)E+Fc3cEH0XNZ5X)^a]0Gc&7=<K\85]R.D8AYVgW=XbVHP-F/)=
YaB6b?Nce_70@NHXU0:R<C5#2G#7@WJ_V9GQ18f2<[?I[fD_]J6A,H.[N4Y2ce&#
7[K+UASYO).C#]J8]845B>O/TI6e.CUA8VSHT:d<ID;<<]N#JLaUf-14YgVMA3ee
H4V<?@XFP^K)QJ^XOL#^8,IT?VgSgI#ZVeDZN=0>Pb9IS#OLgF^C^[##QR1FdD=M
C88+U?=&_G7B[c?BJRf[IRb^&TZZNG9FK]839RI-^0R^ODBWPLcGH]&\gSM:BcM4
Eg&DH.JG9DD7VNLb?6fCf;f>U&&^7HPE\E43b3&7L->NY^KHWMe_>U&aGJNHXFU:
MHG,V:2V?-a2)FIO]^G&eD_H(9#SHDL(>e@.&(TG)[PJeK6Q\\)dB:7PfQG_W@PW
FDP/f+Qe:cRSN?+=4f<HD?.>)WSJ\17ZGcfId&E1S;VRRX=]I]0GNI7GH4U>gYI/
[6:+>PX(@DD8PbXO7bg2@?ee4J)3;F<:T_0.35NEBT5O<VJ+D2ZQ>1&WGYT9]dK7
QaJaLM.J[#(c0>Pe[4&YF=PC.=7JWB<<-SXL6\:?_3I@S@Z@f7J2dT]fUYK_B_0P
gbd1#c^Z.Z+7baKa=fW]aR8IgMPK(@;9>96>#c9(W@^AH0]B_9PRCZ[\GaSV<+TW
/Z:M;4H74R@eZ34G/f5D=#9PN/fLd;ZIF?LH<Je1Q=ULWLaT._.7Qa<ZCID\=A0f
G29(d-Sb8)L,=36>V.LIEaOe_3,F9EOX-R5=I0Pd_M9&6U3=K334&6XAY+^b4D^E
dJ4f.L\Z:=6c);(AT+g?]SF:P=#B&T#a08)b5WCEfFWg8_EPJB>JN:33dd,_XZ2R
Z=55R[4_=bA)<>c7X]VJaK\KAbVVB3<,Je&a5.dAG)^PG>OOVZ97S;\F\H;B<gb,
0UW<>fL0RGKR.##4G&IcO3Mc+8\1aPO,BS,H/L&BDQcJ=d(OB[FON7Qbc2I\._Q&
+N7/+SWQ8bPUGCB[H_60]T:YT(-\G3,0<3ZZ[[>/E79fM[(@;7\>Ub(;Y,B7M9D6
ED_+V<.M)27Cdaa:\JUJ-f)XRb2:A_2:eX@-3^DJ45?cSCdA7-9-Cg.Y9<aDcV=E
QK(SOf0e4>6;@FG3=3A5-1e3OKd3@O,gPMOcA+@?GYa7)8=[cHD;V#^#5/JK7=B8
F,?^0PT?3Kc@c@@L:gR6bD<-V23\SW]1E)(]f@3e9S)(,1AX>^VUbQ?79A.gL66>
PbW6:+cK,F][:Z@:b<@FY<\Y[6bY[cX#XMQa6E67.Bf/CER_<6K)U+O<,gH9c[C3
31aJ5:9(bXRfA7-9E76]=T#G#\>15GOUfDXH]G\3fHg)40S8;T3+L[)+2B,Yd5T5
V4)UG<P+,K.K2B4bgUDdY#aPBP;I[2-^<7DIJPcc.87\5>Qd&,1^8(/bN:;(WUD+
UXN2K5T/;_2&V]cE<HNa?HYH@>cVeE;ALcg@Q_Z^(LWQX,/^d&^<VQ3-H7fQ82H5
2PYMbUPCI2983WUb)G:]aYK^+8bZFL:d7&QW5CbC6.G#@UA<O-91JVHD0M=?e,Qe
A,Z7#K\YV6MaDY/RD,a9<P)DUT:P:I+&-/Fg+36+Q-:O<S@0;]SaJ^Q4Y@bLT/H\
1</C+EZ@,b&YZ.M+<d1a0M>HI9fZ0dbc>BC6@@Eg=Ic&FLZ+=4-ZbVJZUJS.&6()
PB&=)69+<Z)feggRZd7KFc^OGJW4)&P-SfEW2KNIE]EfO70&)VC&CbbbGAJN679e
c>L(TY]JI6AI<c7eBdV&cJO+2N)YA:V2^>Ee,Q\Nd(,))R[M6UaL;^bTGTOK1aGS
MM9,DGSTId3\4-Z?Y^X)_Qc=>@--dQO60D>YI,QCO8S,^50R;QOW/(gBA4T=S.>^
d0NJ#EYK8VbT\5A_R0:IU;-/MT<M#3dc9eU-C96VYMR?B,Nc:GEPMMg=E/JX=dE3
CZ(@=H/Pf7Ua&=:5SF5FB-gQK/0-;9))Qa?F@:@+J:a;=YeU+5+2_.7<B#K#992\
903VUd@2Q=W?VS1A.,C1[d\P3NJ_CbE#:@:&G^,;JOU65=MBa^Ea;2(8[&-Q1>M0
W=F=5PdU^IV5>6b+Df3^OP[8IC,K.P+bML.EaH,SB<0c1A]WVJGVAFNX=T-:/V&\
Z48:)OU71\<AE:()Q]#Z7/,VHD>C4?3SN[0H&++FQ_^62HaV&.I.HXb1D]N_V<@C
8YaKQW)eQG;_D&:TWCFcSGgN__Q<gcc//.1M35T7[aMXF4eCJC9KE0L0#LL1E72^
A1ULN=&a(:8).a->.ID5^WXePWWEf4SJR._35=5,WGMZ,f2ZXQaTUA[\WL#W>5bX
/7cOW2XHX;8(<BaJQ1f#\?aWW1Q7\DYA+I<\g5P,26)dL@SAd0;E+RQe+0e^\Z.Y
Y4;O^aO=)4?H4B]8WI0I<&B\:TW.6N7QZ/g-D7Y.a.+eQKES<&\#1?V-a\&SIDP(
UQ;LIHQS]M=\#\P-,+JD,@3/&SVe2OF_H/Z:I/Bc/O@K7+=O-:E,U/JDME8gC.Sf
b)H]1TH?W,V^VEH]+O]&cSSMB9@A2^XQ#)B+4ULQD]<R)e0HIIJYKcE.J;Q3c]Z7
?OXLG8@DLT@3d2Y5TKd]J+1,02_3c1AF[BWAQUe&M_K#g]13S=8Q]SA[cI70AQ;S
7V2B>5<bT@P?Z68Yg<9\b7Q/9)>SWP2X=9U,\<[=R\-==-VTDd;R-<@f.^UD7^VA
K+Ne>N+4O6J8HL,c=IA?UW2)B4^;6R?L&#-c>C&5SIAdAI;A/U^)+=b8(WR>),6T
[.Ta>5[AJ[K2a+beE36IZJdV]Z.df?5_]]VIII1KI8Vg825^)ePHNLU=5Gd\WJS6
eB_ed)?R^@5+g60NIL_Zf[85aRLVD<YUAYI6]W//^cKLSL-AZ-:dc5aaKXAPJ[WU
\F02V_(:V@L-UAUZ,?NM#+;SJ[[;WB>;S^TSHTC?FE0\O5R=HU7YL5[H?b5gQ<&b
T:0+8A<(3@,25.1,[70ac=dN=3UA4=NF))4S]fE\e]-^D#]/:0MU>>E]JA_&f@f/
F8b(S4[#LKT<Y##(^5F]0B2XARdD\93aOPNIP-geZM>?FR#e4,=@gd.]:T+gRKIJ
Zb#.KN^VIH/RK(_1VAdH\.ae,PR\3Bd@K+-/=/[(,G6R.C31]\XgH8Z[)4FfMZ@E
,#>TAUeCg?0Z#0ZI?\<#DZ-\g;.b5AFF#8R^HWO\],&SX8INAQZC91,4NPL9B\S5
.#=OX#8PM^KB2.FRL:^07TSd9/2?9d?ZcI6b:&T&=R@1dUL-Z\,bY&_fM?8JXTTL
0E>@?#(2O,Z+206W1aL^@SgTMT3H2WP1ZD+[3>:>\9gVdWEB_E&LO^)G2V]8?JPf
G:)E]Nb;SG&64N=,gFA+gI[957C<R?;EbP^<2,SO;f=QLf.e.9AgLcBI4c@_;5EO
cB01-EB-E2S(VT@:PS?;7ddG&WWT;2>L#-OSSID.;TbWb\Y+N/.Q;Jf2?g^J63#P
cD93NPXfEVb:\+0U]2Q6d</ZGXb5C4aJBT2RGf(3F.7F]W#6LG=Z<<;5KC5GJY+I
G]83VF/.fe-_MCQE/bbEPN1Hee9Ne>P6.fZRRAZ7f0]a0<5cT&53RC^b+4/C2c@A
+_H3OFU6.J[7g,8^LW7T6L5RG1VA&0c2<6O,P4&CI6e:0;([#a5g(eb.Z4G<_8Ab
eJ_;I,]1K.T[L8/>fb]0F5NHD6K>:;ETb[A-N/2Y[+a#+0HQ33=OJa=dF#F_^OVV
<d7c8[7@GgL3HK/:Fg@6f714N0M@Z01JNRU;10BBeBZ.I?WQ9\K4<Aa5(AU&,4<=
NbV#1E+WZAb0+/ZXOXBB+.JWa-@Z\SadQIO5b&:NBAfB+BgdLc(/NICC;Af/L\6R
RF-;T9S3EQ\T4gbbOD)3fd12_dQc:DR.#N\P(&c-HKd-K>X<IaMGF0B/OOKP[.87
[Y@Oe_NcI+N7b_<UR=3@JbNNXQd5MB@f&4)1T@gVWFde?UagM/5f/CW06K1T4CG>
^9>8V4L)-VZ=N+cR=5\W1<_.EI4XBZ>VIW82MdNY3]ZGO#ZTDTUVFFXTgYD+SL^P
I\1>??=RQSTb^<PO]B@e-&,X_VI85Ad+FD=a\Pdb<[REW;5<QUIa(QdDJ,6O(ECU
6e[\@8<a+0df=1<^^,-V7B2Tf.1UU4d@^,FKW0:ZJ#>c4U#;CX0.1&9QOC\2,_@9
V:U]>GW3UEIY+OCVEXcIg-a[9Q^4@RVgZ&aTH8bCZ_\RFbT)?0R^Y9Y0g5FK;d>d
d.8g=EgZ4,OORR^POL94K^PF3e>0Lc1Kb<@feM?UPDJ..F8EBO?.J<UMaFVMAK1f
)<9UB5GF]#b:WJS@a40I>S?5P3;9UfRUP0XK<9H5:;?M@_K/)O3UAf\4QC[#R++.
NJ><ILa[5=>2E>(cFX++-0ET9=#N](QP>^Z_B]9Ne]f=]:de3J<TgD9/c?UK//a4
?FVYHVWYIRP\^J_>/<Z<2B2K@U<B-0gHLYZ^RG?)3_G:[]b>3b?VH6d7K;HHgggI
\8Oc2]cH&/4OVELCTDBG\C@;3M^@^[@(C5PfDZWB#/_9g7B@AWLb;?-<dBE7(]\Z
@]PbdF)f_1Aa5:2=N(.M019_&Y#IcWAVEI(:UG21AJMRPH<dU3PLT;(E/DG&Q,TV
G5LA.=PDCFfHO[6GG[f-Q8W7(DU^O4#4Fg\3XPT@cJ75NI-EfY_8e/dEFSb-;-_X
_ZKIX:6--)X9X4c7)+JL;2Y5;Y3XEWXb[R]0U.J5[EQPO3WB#FgQW@]]Oc6G19ca
Z?=\HJM9_OR-YN]\f_3662T(FO99;K2,O&^<IQ\=g]-J_YKIQL#U:5V3e?ZOYXNe
^,(S,>-g#@T<>YIKD+A\6KIB)YM0bO-H@CGeN?>)@6f):/Yc#@,&41K-ZY+9P<[7
CSS_-=][aR^==>(ZLHGc#3]6BV;&E,A19_&?RdDZ^;5?8-;c&&#RZa-\X</5Veb\
OO3X(00f\.fWZ8J5UW,<UKW8;:M.ZSELHOZT7#+W@6HT)WD_]A5W@b5cMeTU+7Ia
<3c]J5DZ^P8EGCOb@,5b]Y68=HIZP[e@PFg]agaWMGJ5]W.#-A<ZTFQb+J>6#D[L
_<1+e4c3+B85gB<Pb,cU84R(cL1W;2e@VQ=FNPKG6YV\FOR1WK5,a&DIV,+@+VRU
?^f,5RE18CY^U<J)Z:0Kg][.)L0^\RWDJ]=F:XCgF@I+N0EMGA9UP2;+;,3:d;.N
@@,3<FRc2#gg;]V6C0V5ZC)EUT03Q;a+VV=<H8<a_aOMaY7VTKB4UNM\L(4=NM[Q
GEU&UALBGYDQ8M--9C&P;c]9;KU5.bF=/?N4GJRF//Q#1_CB0DO9VU0X2a(0(6_C
74@4#]SZ2a?ZBP<4IPdMfBN0^d;)@&;Xa<YX<9#N?:S_89(J-a_6DU^SH\C8+[g:
d]EE+>H#+\(R)F<Q5-W_+JPY=P1(893P?PO7]>P>?Gfc)30+(OB4&Q,=d6C(Xd-0
f1[XN<\&e5R=&TbbRaC,A.6LDWJ^7Q@LX\MGNDK4M/cDa5M-=QAEYFSQ=5MYNN?>
c0Q<G,SV=F^_74SUfN3d,9ZLbTegU\F[(./FbB.A\WG:+-=cF5324#.QZK:HIL=d
H-/Rb9;;4KWcaEV5ORg,;K+8A4La,LK#6XS>#(G-]cE]UZMBG-YC1&8^\[CggMOR
8EG+VF(\:g8_829baKbD7QKBe\TR3<+WBX7HBI8_VgKS:W67J,::-ee_.ZIcT6:3
C@,.\1g^D437;W&F/AZ<@G3>CM@\/J=5YdJKVU__1]D0\=UVN;O^#a1KaY6&bFCI
W>0aLc+cEBMH)TJ>3=ff2^ZC]BeWCQMM[XW6/Z)cEU/((@0g9VfF9.POP_9L>S91
@)5d+5-/a.10FeG^/Ua]9\0+W-(<)ebW7E380&:5VY-HH-7dFJ[R3GNKdB6X#5LI
e[4TE24KHfIX])#CGc>/^dSa,<)QXT(9RK#N]J@N98gWf5XW5+1&=R(V):C<7cDC
?B)2\2##:9QY3eCL?-11Uc#OV[gMf0aE8+b13IX(C(\4QL[?1H[VD1-(DK<WREV#
gM4,(VA#0XRQ@<.FS@&\SgKF0(K2YD>D2cK^B;WaEY6S4\:]62UG+L>4+.HcD)RK
cP=>D24.dfM8I6^TcJ/P1#S\03O8aC-X<#Gb&X41R6JMA]36QEHD^1\,#)YQI8)+
&eE?K62T]U(@CDc2^^(Ib)(?WeU.#\77/0F[=R;55PE7Z0@4.CXK//X9OE3PAdZ.
.VU]92Sd)Wf&I4]YaD@edX,0=776F,EIf7=Q72F)GKPN&>Z9\#X<#NG1IC0@6Y-D
HYS>BC08&F89\g;CR&5@Yg&E4GO+#Q4TU4D/RH;Db_?VBfYa1XX<=G&?7c]+4d?Y
IW-Af:(NbW/>R4XM?:HKR^XUB.^0RY)e4)E]XdMERLU=M)=2,NNIBf&@E.O?;INf
g)L6I7bLebaF24Dc,=gg+b&[34VbV2b&;a^:=FT.D?C3E39.>C&aXS^C0PDCN5NA
F23bQ::-1_HbAZVW-@b-]2UV[:b7aZAK):F@XN4.((,14OdW)JPdSIEB7YV)\+-<
;S6>\I8SITUUaC(LHI,94)^AHB127fEa[d09a^[eX[=VLQ.e+@T1G=cOf6E42a55
P@FSQ,J&8=X<C&1gGgL61&+UD/3GABA?<JWX3G.?-5+gQ9R.bgU1_?PR2I4?F#TY
9(F7?IdD]87&f_Y,I.\O0c^LV2>^&#cK]:C0SeHe8_+[>R><GNUJKI(J+/FNS[g]
X/a^->FUAEZ7L#e[+D#Ma((f)SEF_O]dCO.[LYG\2L+VXR8E;EU(H)2(HAdM@U=9
7#.Z[]J<RHd:e]Lcd/g#TD\&R=c@Q=88/d76(OLef1;+&AZgV]#X+]HOVG=&GD7(
FCc^JNc1ZB=5UC(HC<UES#d4A&f(G#K7O[,DP;O)6ID=X9^O(4<6WHGL.<E]4NGF
-GP6L1N94O,&_D9L1WcZc;.]+Ie?]G>af>\L(+-YfbgW93TY7I3G@SI&QD1&K6_b
#\0[#S,8?SYMH/7YD-b]7X7Y(/64\9a\&eDE(G56BA=4V&0XGD1K&@ZUEYb:\C;)
P3d@3HD<KfY<T]PVDT\f=0a]1P.:gZ]A\()9L?^R8D&>GR?NV84O00bJSKC0c.:A
>L&\B5=FR?RWN+\ba18VDDZJZ3^T:a=.XMO@H003\4XV.L-Y>cI]9<4Z4.UE0WP>
#9.D3?=G60bPPVGEX]=0AFGceG+RET_eD\3K0dC9D#fKY^RW7()-&UJEP6BeMf_/
3b0FWBX67-\==];,]-:R5B/bc]^R]5,]#_#/YO)ZdJ+REC\@_c7MA3)T^@O)]O^G
f)AaAL9^cY?L>6=T[LRW@aA_J^[+dJY+GLDg2;c#HgGCAWKWbcc_aPM:I-V<RU6[
fc,P]#R]AB+H9ReFK]aKC[gVN):&\B,L)eZ.@RVMLSRc+a5L_B5@8V0?I1WGV^/f
&4\:IZ#RW<2CXG->97>WECJR^G.3XdX\Lb)6cBH)UfP6\:N7I[?+R0;@>B&X+^^a
+bO_e0:_AGG<=WLa8]70_ES?CSY:PZ4S.FB)&/G;7L_#/+:_Ubd1&7+@L/@fK^EZ
S#]F+2F^#OaC9R-aa>];AH0U92A7;+46fQ^6L&B6T@\:,E\KN[cE/2.R_<ZZ8]#?
@B6DM#A_b2BI]?8^UNVP,gMFaAWAa[M<cC(=Q;-e0gZ9:N#61Z8NG=74&;O+RdNd
N+3J;>_eE_Z+S5KZ/246Og[9F65-fD)ZgMK,VHO#+2+_)T@#(YOIgc9dG:,BADY3
8B;?@e0BEE5-7ba5.V+e?7?NcGGa,ZHV3;:=PJ8:GD,,8;/\M;a46R_^8d5V]C99
/dB2YUHP6SPbMK.;4KWTJ36RQZ14g@EFQTf(6.__C(7WcX:M\B&NQGP737I#+\<N
cfG5,e+A+#>CZd.J]VXR[?TJG8][U:HGFR8;aGP@80)V@^1\UST#PaCS]1=WE4NN
;E0:F^[bXJ]1:./9XaDH:F>_XA@VSN=-_\O.60U?LcMU-8dHf5K;S+>(N-V(CLe(
7;0PLdXV]EWRNRaH=.:fJ^1I:.Wc+R<0d1BKLg:XCC^/Y47VLd4SRJ[5TIFRAg5\
,:]:SEE=>ZRN/P>G,MBd_E^L=[^5P7f)9)..g+cVG+J8\,PKS@dUI[_H8>2f\Ca<
73^OBQ+>\RTgbXbM]X5L:T0WB6-S0F^YEX2d=[@PR,Z7S:Y>=:(,L]c82N^GT-;8
0d^[.1fYMf0@/<MNLXU_42G_f-.)P#H\N_UAb?(\C&V72=A+J(X4GN>YDMJTSF3f
cJT)[CLDO<Ng)5JV<^ZFN521P<?bO9TJ(:=Ma53@-@)A1aBRM&g^SX20N\7:WgRG
]I<#aB&#P700Z[(IT9U_;\QO<:3:2QW=/M_W-Tb]1NTKUd4g?>M?X2T=ZORPML<Y
8-F[g3@+2CX:&9?1T17cHO:Y8eA6B=X28-6feWZb:(cP+/1>I4Ma@-Z&_2OV8>ec
&bJY2W#g#HK\-]g:SXLGI(3eQ?4P7S\HZ^;>9PE2-#cQXO)QS=Pdg(PUYZGbJC,:
58;1<P5+eVB#IODINZ+E3^FYJ/cXP].)Ka=01-23IX.)TMgAE_;O]09+Meea/L;L
V+&E8=;Q_U\HdcO6g:^\56015]PI]Y&E6[G#&;S2-W1H#fC)+&ZFN/RC-K#c_-MO
e4d6F6B2V6M5;4A4Yc-,&>a<3V&fJ3#>Q>=_PBWf7\:bG/6.J=M-WdLCWXDJ9QA8
gM>7;+ge<9_A:SYHZ#&L)_5a2/)d?SNFCF1E7DG,V1CUB<QULA7U666+;dBD&<FA
]F55]<,&95I^:Q>3R1W3G]^R:?KE-4<#RdK^YV:dc<G](C:39bSM-WE7(R23]ccf
fFR\LC_]dE<L,<,8U+cG1@\WG5.=&F:E6+Z83.0T)<^B1eFTe&>[K)W(YLX[^VC[
&,g#_DU9,e\_[I3P,VZY&7)GP71]?3@N5A98E9beN>YUI]=SFW0V9#D^U33@NE56
RR@31)Y^ffgSG8OaY>_N4([DD)7Q?07WCZ8K-W&g<L06I9TdQc2+@L23_a^ZSTNC
#CaK<-8\.(fK,@PT7PNMDCW@#65UI8R[N-=Vf6dD/713#G9DDWf>X3OV;/bcW2J.
OD-6/=USWKH9b([[M#HT-(RZ(R5)e,8b\B^I,CTD+;4_/.P6)UELYWHKfSR4GYIN
V2<TF#]W2.O+Q#c-f.V[EDV^ca[[IPB5U@\Cf0.4XFKUXf8S:S#0-&a_T<)H45B]
PaX(5O\6,][JL2C?44W)0TV@O_\.G__+53^R+WNB^[?I3W<R:A1g&5^1V]BCgc95
F<)S#)BQYO8Pg,8=@SI<P8:UTSc0^-.gKTOP^4.O1)2CP.QACaS6DD4dLI_C_&NX
aWUV+73/-S.CV[I3Y2G1BPQV^^_eV-K@_E<e_I41UNXXf5[N4I@)+P<gD[Q@\7T^
CF.V4:,6YM.B]YcF&6Z>JBe:.\d40)QYI4SZ@V[EQ;bg3IA>E#aC/ODHN1<0,X?8
b#FP,MN=,G01.4g[=WE<A7X1\/O2?VDKBTK:dADMA9>&;2C\.((1<5FW:LC2Da(6
3.1^9/[BIKgNab0#[9YGQM.agS=dFL8SAFT0ReLY289XKbQ@;5PZHMcGK4J]T([(
c7?.,2bc]PWXJb;9aLUG5&:.0ee7;;JNU-)?F<f;1OG@7b1cYG7M0Ed/JeH,,^Zg
[,/W6<=2(cLN]Yb)=^@2)A5-VaO<=W@NdNP#@&(JI+JFZT4]0/[La,#>3E=TZ8d2
#:@)MWHZ7bU31W(eG[A94Yf8+^Y[CBBb8Z_S/W\)ZOAL@_,SHPLT_1_(Sa/V#Jg=
Y:ac02[;dOa;<H=I\5+2?gbaPIdRAOTAa4f^2MMe<-45[J54D7?TS0S-5]1edbA2
DP][J]G;-8E,4G[X,eT&\]3df:5,/\P,_Jc#B&(JX^aCFHV/ASg-^)/N-gHO<\>(
]TY;+A-N[R(bV;B.JC4@5Sg+ND2+4?<Vf3\Y-ND85D#ZSLcXbAW:/aeb9K3-X>J4
:YZ8]#O71>=F2B5PW&PU<.@I6Q1>M<3+X0IK9L?H\<Y41?RNN:LSg^<KB6,:aTZB
TAM\MZ.bA]D,J>PdQB7-Ff<9,CbX^EL)48VA/D,N5CUABKNF#A5WOXg(U7e#@82L
/gIJTaU==G>_4N&bG4PA/.7UY>A70cP(c5\a1B6XI_NBeEUV]DM#R.9Fc:GRP=YQ
gJR<=UQbXHGR#&Gd35b2_5_@aT5-:(?a>c;KbFa)&?SU1XUD:<Waa/fAJF7Q;FY#
SJ;C:]X-;aZ#4G&ffDF1c<A+C]_6Jcb.MEd#cV)GR<?9cg\[I,YN-^ZVK(L)EZVX
>I@aTC,)PE;Dd9eg1\^];-F)..ENJR]_AKQ9X&ZG^)eS-&]6g^AL[4B8W6fIHKLA
7Q;+HCg[(W(\F4e9+?7/d2>@IMV9KdSPQBb9g>d3K5:&0=;gU&U19P>)\??S/^.<
gaJ\ZL/.UJ7Sae9(+2Ac&/_X1fcJ+(X&:2YE1BDLF/C39e?_:K[8Fd/N(78c71ZY
1GDHc1\=2+Z+.LAU1Q5QLX;3<_=B@d[.5)DMTIgR?Q(Q9X5>bfQ;P077B/J1GJWd
a0P#2LZ#dDU(Y#SX6T&^G+2S?JdgZ5fLLD1N?ARPW[.FN6_A;;6HF6WW79,+KG<>
F=D<LCe.TYW/(6bHT6:e5^&6a2;0c]UOdRHbf^BVGE)K3b7<OLJC:;Q0#f=8HBH+
3+Z::#M^R<L+d;.;@>#8+dE[?c5Jf#<U#C97Dc5SYSS;GN:-L,AAHJRfSP5/+Y?#
Y=Sc2Ob46#8]V03GQO:Tc8Q,DeE,XR.NZf7Ec=(cN/_NM[Cb_4,:N<5>PQAYeHd7
bFI0AKHD:JDHVKE2VOHLHT0XH7D4ND[@9H.F6K&HbNK0SSC(bFgMVC]&4)MY:6c7
9\:GZC^U;70Z3NJ3:P[CFTCXaDD,+CMRFM8.C#F?4T14C_N]:_4T2F=V=@U),++E
94.&HY>ELP:>PHa4D[G8<];H<@@&baWB\K;d871-J+W/8OYVH03+WJAb_DTdEI#V
X[TNH1)G@87cCX+R](=0b_<6Gd,-DY98;2@f2?;?dOIZ;+WZ895X3>5cB?I<<9gQ
(.X^eB1fFI1-=Z?:YP(+X0:;\CT,9@&2MeC?_N)S/SIA1PL7EJWa7-a<.8C3]PGS
+:Meb4@9a^[-eMNDa5MYD>CV>I[D9,,8X+&aP\;aIC^&DSY:fGD+8EOM7TTF&09]
:)C9Z-V3cGe6&H7+cC9K@cE60e?6b[UU8Td@NY^5Lc&LX(8d,/.:SeFJbfE=1ZbY
GBWL,=?45K7@?]PXL;Q1+F571>FZ,-<#C:]2[58G0Z+=]<,+[?M>,P6.X.W=<Qf:
XXd)@eIE1:CQS18]38X@U#(/XaHG?UfLZ&g,L:0P7HVeg\;9(RTEcCe]_K4V-:C.
<#eN+XeE6OTF_2)/\4HZ,dG\]c?+g8R6WSGS0SI+>@;>c?;)-CggY1H@)^]J[d//
=V(bQJI]PFA8<CL,.\X/IDPdW/5AYJ5VA[g]]g02UbcU^_d@,LTfeA>f2T2+(]=.
TYOgEN,5IN6Y\YKYGW@+@;9XMAP).Ddd&TP7XR&Z,IY@<OHVALa.0bJIE03C94?Z
8.aa_(;1=d3GJAGV+g(;/cDPE4RNX_#3@U==.f0dI>4c&?6=P_d[QQ5g_/e[O3.;
d+gMC06[1Af+OC>U9LUZY\>@/:T_AdZ2>[_]SZ1cSB).>O&BXJ#NF1I[/EdSF4?c
_2@.gV6/+?;(U1Jd,VBWS>=,FLAO#0>2YHGD4FD6]D4[W=<VXcGR7V<^97HZdO/3
V?>Z0C0-QO4,,])e[FXOEI3<_(3cS+bD/#\4X=YAQXM(1-7X09bM?:\G5cE:Y._4
4:g[2.,0915cOB:+OM;#e)d=S7:bBeRK06W32b_8#OIVWcg.QR)-fG-L9VY;-[>L
E_99:19+5SBR>(G5B7(?/_E\AaP4,]F8&a82ebL#V)H;U55K\V:^ZFNLOB36>P+/
6aBX)N-cH9?]^,0S.N&>U#f<79L]CaSQ^K94TD1]L>)Z;.>.[\+Q0=A6TUOVY-C#
BNWI=M\K<(#46KHED4NFC(d.a<cIY7_2CPcS,W^g1P@8U1\=][:)L-PAI3UUf@]Y
2UbO7KOMSJbB#J_-NCK0;_[+2:_IO#5U\P3TU(gcYRc9YLV#]d,KZ-KLA,S(QH>>
GcL=McK;b8,4&cb#@O6H4)]#+COD1PSN0^eg8GeX.c2:CYafcZa_7Z3V-bGKLb_^
N&V&2X0&4OZa#JgU/S0H(3>I:RP7XDEHYX=>?@6\DLH>e1XB+.,a)E-J+S1)3R;]
X5POa#,.+dCQJ/<IHJbL0f1&((JfKg5&fG#KSA<4XSW5KLTQ=1d1IRSf\N,9574Z
7(KBOM1_/:#ZS\eG?L@-?bKFKW2VNL.f]O0WC[]D@LJCE6B#+C]<L6BUT[Fb3OD7
G5Q,>V?g-U?XC,cB8OZ?&e_.\NQ.?WSR]^DVZS=SQ@8(#HOO-&,L<>P929&dDe)0
HZ)T#M\(/&5B,>7.AVMA.9601c;6[(.P@eEA;cH_UVS]>Pc#gaa=RdOd89QK[=^+
D&\XQBfQ+N9\)HACY5TbOW\:H)MIN],Nb1De5\9:,>JYH]:3:55)WL_92;?bX=;a
JY&]2Rd.I2cO9G8Q6IP2GDf76_><FKc_+CZ]VK>9(W701&Q9AK1ERJ)S83a&WdH(
O;S<2/JaS6UK7_I^H20QfYM(4:A^148[T]KTKW;LB>+L[DfJZDT/6PY1)XN57PZ_
(-d5f]g;\4V/9LDPW2IDIY1N&AXEaFM:A^W.b48FBaD0]@:U3EVEKZ=SU3:)_f&Q
b0G0eYTg:B5G_c9ZG[KSRYg)OFT\Z=Ag)S=:^]UXZW4A]N[Q)LP\,:P8b2EIV@g8
VR;#_?1^H3b89gGd&]NL8KD)g2(C+T7M]#_UVE3775(Ud7)9QE)((-3,E8K74R4A
A1DXJ@.,LI_@PT:H&O&bO1N(839ZJd=-TRR,@cEF6WO:#-:>B(GDFe,-6V3O[7P:
A2DC)-4WP.9LS(6+d(#LCB+2)45TBd7U<ZA62ce0(4:X^/EeDXX)Q+M776+f#V#M
^OWdEVWQ^0L35X&dAI@@1YDeLg=B;H(X>gWDZCN?YP=cF4g(dcUNL08@DaC<+&/+
7^H8e:AOUeR71Te.XHUHRc2Ze)&eTW8+BBdX;_3)gcY8-MdSR=BZG3T^Ue&4AV)L
_@JcZXH]H^\VHAAWMB_SM#(M9/<Ac=7TQJgc)<.,[dEM\^9BEPAU#Y/ZW3PX7/NR
E\1QdCY,7-b;N#:E.65\X2PVHF3OJV.8\,OS#e/(G_GG#YEcUcD/2KGg8ZfdH.^8
<LQ6BOLb9^HbQ5OJ)<\F7<\(V+J,/M);cA\E@ffP2L[B:DH5Ia8<A5Y>KU-RUL)S
H]_cXU=L]CHf>JI7.F56ZH_HS1MQ<<3^1]Vb((Z\0LOP7gE\H@TM>X@cMXcZS>]2
585@?O2W(A-:E.AX(;CAa<\P]O:QZf,56eTa^>(G364Zb2_21F/^:9U,9N7GP+17
&K?G>?U^&HH9=IPZR09^2LD<eS[_,1L[17?@W;bXU6N>TTA4;</V\+OAAPI]6EF5
D6\1bP-_@3L<)JgbR+4V0<cU:N[(AQ70Ya5BX2ZBUS4:PSN2>A7Qf<#^WD(O9.e?
ePc+Q&&NTOI6PT\/-d.7L2,5X6YLSP[3I[#e]9[SLXO4VHeN=K+@++@:@_T\aN?K
BSI#]CMGOF\>H2#1/(+E0NT7dQ-EY:&.bSR@N6PQN=:gY[C=17^<1)eVVL6MYRgQ
RDP_d<)]-[]F4@ZVbb[TD_(XFUNGWYATQ#[(;A,c?K+?fG;0c7Ng\,>X;3)>;]2.
@WI:gN=J#7M])NDW/8T_E-TUHGB-(aHAR]@7#;P^QOR]#HWV+2YT0fJIR#1GRSQG
dH)[XgG_L[32&>Y+K0]1gZ3?(/6(a4fJ4HF95P4d3H::G=(H8^UD1F<fD]3b#4[.
N]BSO07]9QBO>g>8J^gC,d+afC4W(:Z7\Y=>Z].<0gC7[0#Q]]#_S\7&>P3GgE7Z
,@7JU&cMUG.T7HNJXLXg&\IXNO=&?BIZ2T;LRA/XFHO983XD:T(;@CK<ML0M35gA
(.:g803@Ga^gB9),?[3P0QBLNX3]0d4(:[4_?\1T]V,-D,OX;0=e)<(HXHba_Kf-
5_5M9(Hfb_3#0bU0,KfPRUB[JP)U4;-K0A&g&S97=[W,a]#T+_/\?-5HF)0R_WSO
1dP.X+4#?&:&83cJcY[T9NRcKJM9eX8L@QG1SJ2E1B,Fc,<XHQA)^M<#:^).5VSE
)HV(Q13BE.C,C_,PI[/N=_5^=GVST=+B^JSH/V1S0OTKad45@>VED])febMc=_L0
L3N#27A..4;[R;,OZb@aM=YT_3N,1bCX3J5(JWKU#SNG#cOCJOa@CP10LS/C@)8B
.7.@&4L+<g57L)-GTc^fIddg3JVV.MQ_WI--2F<OBbHJZCN]RYE:Me?Z16-NLR0\
_5X/7(g4f;63RBMaM[@e]59a,B.RO1LY;N/Z.O/Ma:F,Fa\Q:M:HE16d[g_RU)#W
CV8d\2JK&H+cM1eHdH]cJ?a8+#Zc,b@BE8c9L<]?^g_79a6&F+23X>XdWTT7FP8#
MJTTNfe[=e8?.[^[S9LS:+:e9WgN&,4F<T?C9_f<#.HNP)JBZ>ZfUWXb8+dEa_dE
-E+AB/[Jb1V?Y#+5?N,7#M#[;2U(9/K:DS<<&?59;_dCZ#+QRY==C>TBPWR?gVc^
V9Q-@0H,2HR+,B:.dY:3<X]SY,b+X<N]SY>7gKTG\?NUD-(1:TA3aWX)E-KaadX&
Y@/PTVL5QDaMR4;8S-NKW9.Mc-.C)8=3N7P@\IK<N0[.Rc5H0/FTM0:\2GeZ(),M
Ba,F/W>EA005^Ag36/(^T#.FfOc=27Q^JXf:F^OS]/I[1fd^@aH_5559RfTE]I.N
>E8adX<(Z^Va3:0DGBeCYLPX8\KTcT<R1JZS#f1RBGF7/fR(SeB7TTE(T)V2aP/P
@1K1QJfKA@-K:b8U[0KY51GS<YXZg=dYKZDW?2&+Q-51.)A[@JPW,4KAd;L+V/B9
GA(7I&6b@,385-T6bXcAPS>TCQ3OQf@F5eT6J]BObR?HO<K5g5B1cS4[,BRIQ#IR
B?9V8-6R1XOPaVA]Y>LCB+R;_-=+Q(/7fO)QKPc.]c/KBQdQBe,S9+N89f@VHPJ(
cb>+&4F8(W?59[fLDRAB+<>C:&^eXUT7JNXJ5P5ZV;V]_dg=IbHPgQ.D(f^[LW&=
4X8-dMP+dbc/7-#YD[O.,G[>367e;cG-EG[<2A1EA0]0A@A^P=.2?PV-Tc]C_35.
Q?][\M&4KYEN0f/bY0f92CD=,8;]>f-bgF;0PEf(WSD^Og1fbaeVTZM;?7<KAV0J
@09ed85FAd[+;1[+@@f0C&)WMKdW=VR6+H8&TBL)J/T]JdQ)UH(LRTdXJ082PD9X
EQQ2NgB@<V)C:-Wg1N=b?)([3V9.f,KKfZLJQ>WQ<IFXNW,d=V@gfG-?BeYQP#S+
MEL[IdGg(d_-2fUTdEK=CEIV3XB[.9OaECE^LfB=.;UHWg#QeO=HS\&/(R+4;O>>
;J/fI@L^O8T:#=SZ^8/Fb\YWD_(&_RQ?U6GV__[V+H,2Y1^WUeJ&:1g&,fe\3+.0
#:+2d27OLYY)KH;U/IgI+2>Lf_]a(K[C#^2LcSF.:H//Z,g6Lf39E1YSNT6.L&5+
885dWTS>8c^[\^<.GDDeDX2W1EX5_:,8K@acDeQ#IaR]HEdQ8SSfU+[?KLWe\Z.3
Ob/(Z7@J8KP4XZO#I<a3>E-0-SR_3AKTCU_AWC952:+[4bX<B[Rg.-e()WG&/.,g
I03_c@)+U@3X)(OOGQ7)IJ=B2_CL:EJBMNGG87UQL\Q-d4.FJTJfa-M@--P)PcFK
_a>\^)1</3c+M.1+Bg+?:G5.3U9G,-D)IL:X&EK+8ZBdWeQP3]+9LX<]ND^/&=0<
P^U><I[P__.W-eRKK1R/c..O87[N<C,ET/ee](,5D:#fHaK50eO60EKNP@a^1\R#
2MN+DDQ[ANF.Mg>M@\<0[d/ML36aT0O+_D+[Lg?\O\.@9U9d0+T-2\9JWbg(BaXK
+:,67OZ>ZOI;+,<LFC6&75Ve2?a=\0WC;[<-[)Q7CUaCZU]CTfL.K]JFObGKP)]O
a7O]NES7-3(9e;146G46:]D<A(T3/=[>_-65SS3f95<XQV7J0^^+(3Y5d.==XD-1
f=FZBL;X#Ud4[c@F#5Pf0Lf?B4FDBV(3UFgG_8FRY+5daZYe<LGH[U,V0W3T.Af\
#;L&Z]U1+/7LE)]^;fU-^+N9Eb=Y01,+A4)TVT2VMC#cCLRU9WFO5:]92UN)ZTSN
-,/(_0GXC9AFFb]R]7;1Ob?P>JK_-Q[?0=Be(ScH6I2R2?+QF724Z07_FXJ@N)3N
0<9=b+QT3B@gHQJg9e(#Kd+#dN/ONe9=[=^U]4DE0gY_XF.AN4;<CZ=EM#LQ4c;c
=3F7O^ON=dIARLg7(Z),+_T2\W-=c)+#I6[__I^TE[I759XRaB)U;?3SI<f<APGU
S3ZW8C7I+Q<+eABb)&=A&<g[6d#bCKc):<1e-7R-L6Tg@,8&/++PKW(LSZQ>7<]N
I5;1)Z]5f61DGaM:@-FC5S[Qd<EMB^A=94)f^UC5V?ZDW_:A]:I@.bHQ-@W=N.B,
R5d9Q4MFPDPP1)R\.&LX6YaUV-J-/RI?X/._a(JJTYe<.F,f\2(a\BUgG&0bWf5D
LA#UY_]NO&aOg<Q<O^,@+IN@\/6E[4\f=]HEeO^-#4;7@Z2]-,@c7<3J<NdP41C_
NK,H+b98HMG;T6>V9XE:Ag/d0Y-NR?[XG0,TUD=PK@V((Ycb;PR,/SgY;+)65f72
FGS,G57_g)3U1OY\/27)9:3E1fOa4,;5?&4:>TYSM53bYH97N1CZ+Na-T4W(FXE7
>OI@J:U5D#?JDKM/9YLIA8DBX^d=e^I:F4/FdA0NRbTYAC,Dd0.C);GLQ&\.&B_=
W^-4N@VB(F94_e4NT(U=_2L=M-dZ=Jegc==JgZ[)Yb9TS+b)PJf4Q^OEHRQSM(,0
V@+_cd.R\D8PggdTU4HW+RJ8RFUZa9CV]MP1a#V,NW#QCaMb[-bU2BEM)e0<]T5c
3bTR8\LW]dc3XL@1M9AOE),SVVS@99P0#)^Q>K;eG]_(\^;WeY4cG(Y.F2WGX;\T
^(agJ79W9(O>6_dGZV(3(<<,J;4=#NRHf<bM@[e>C-H6;T/LU[V4fSW?]I@2RPPF
HL60ZTEINLXKdT6dSe8Gdfg+@>)X/IVLDH9/K\6+K&_Ig+VQ0aBN=Hb[,&P(&;Kc
/3+=\dTQg,(@C4C)9BVA1JXMW4Z.0.dL<9;(-+JQ&,UZ-EJ=6[\DDX]Rb7G\49TD
N1e=,:2<;K&J)73A9Fd=732#.+SW/SRBPQO^,F688cdTF3bK/2bg/aUB=^8^W;F.
.H653+6T-ULBPE01URD8:=b10,L5S,I#HZO\H09_PD<STL9,YUe2QQdJcfg=/PQJ
KI\+]8-/Ke#IY4XY=+a@Q9,&O:OZOb<B.f4M&U_P^GMXKgGV+ZgUMY&3Wc-VBJX9
cOC+)Ke<Me0?g(^0EUB;\bD[CK<[cMW&a8BaLbGbe1YC4Y7=;.YZTX<R)(aYe(;8
DTRCdd4FeUUM1PGHgBD@<QWD8(I(=,2bYgF<UR<<#(>I)VYP?BMEW5SJJdJ^N8MT
7?80KWL7.g<\fO;&PMOQPU?bcT.F8#ZKL3,UgVUB\J;(C110^D;.=BEcPf88)1>7
GD?U^-^FVg(^@66H,C]:.O5W^AA#S\d<K&U>IKa=\bD5#;I..CH,&+T>,0-bdFNL
3/;I6QH/6:H)F9Z>QX-&27a[D1U=eB5dd[?6>YA9WRaSa8>)(X(T@?:56ge8Z\3_
X[.X2<E_)5N<=.T(CM29IM=^5VY,S7f]>a2#gSIE;gJDBa#1BW\B_N=Y4+F>Q@Rb
@[C=TB\?Z+>E42&FY/_P8+?M_+T&5VXcK.3XO(RLJc\B/NP>-R89=WH#^Z))gIFN
gC/cd0/[&),L#GCYO,5688ga<37;5WVEeR^YLKN2cWaSef<@P6]NY8R.9E>#:SQ4
LDM7XUN:2?=35:c93?Z2.(<]WKJW8W.L.Ofg)4<T:P^<GbC3T-a;+4@IOD@^Q/WJ
#9QM7+H8D9-UON1<USaDQIeW]TUcY@Q+EV3:/QU(3OS.;ce=<]:)-.AbD?cWgTgG
0>f0d3IVA0?#b-_@<#fUJ0=K\\3EcO@>,W0PI2fAJC#D+1fP+\D[_7-BC:SX>>Rf
9g6B7:3M[437NVZJZ)V2cUO4YAN&L8CEe,7g#=@4:3,ZRfVS(HQ+S=OC,)Q[D+4E
0FQ=C7GdO2AUV5\1dV2B(HDC-/D,B^BUTdKNGPI1Fd)ZSd/Z#(T]EO-9]M_;##WT
O+_eedc8UX#0Gc.D?PSg[3c]I6BKFW=)G]/_JLZ=1]J9Z5YRQABef_fcD[#,H38g
?_NDNFD+X/<-@P>AX::41F>,WDO,N]5;&2dX:TV>X?N\I4MV+TXPH9F03d<c)+\)
VPZFMN.#.JQ.N;Y=-P2@cGa9+Qb6Ld3TeK:OA,?_78b2B#VNO+MAI6(<-^YA>B7S
fOR49Z,RK.=21eL]#W4CTR?B9b99VT\J^LcC>&E6ITW6)f,JPXSLRTGQ=W.;QM/+
KIA1e7-g1W0dbO:]TF;6b(:SHfNX7fP;XI#Ld[\#+^;CV;>4EOf.[YgVGB.e.Y-8
)M@J=E/[FY9&c94>>^6_2\g.4+7;S\L,:EeU6CD(cC15+&Vb\06Q\cTO,]PO&:a>
6F+&Q<]JAN^=[))ZeO>,Q=/@41[NJ?8<F3-d+AI2g]2HZaUWg7OafK#MfSD1fEMg
7IF7DRD)&SBI;R#BWVXe9a)(WJ>;Z)T&>@f-TK8526:[U&?5@gWfa4NJY9OSeJ0g
>>&AKGDBA+:gK5cK.3>d(1fT<[G?ae[2cO\(BM<\)]DC0=WA0@#-0PY1_@F9:-R@
0a5&Y>DTV7QHAFEQ6X(_?-I1HX[C7/A=fS.9:N(]/\Tf]dTOAfcdC7YZ:O67G?VS
?gBb8(cf>cR7c((ESeEY[#=LBD3#3HWUPIHY1;5>0(+Y3M]1Xc.^C&Z8;L1HWb43
+:VXY[[V)1gNc6\5?Z>dbJ^4K2[TK,__\0bJK1.BI]<=FRS.L?;K,2H8B9I7Z?[F
Zf74N\^_]KKHX/Me>@TbY];b#aVMe^,J6OKM^8H6TNf3^CaBVVEg4dY;#bT<WbJB
^S2U#B[>db^17XRG5C-L(baSHEWe&MR-:g6M;>(.c2[?THO4C-S>:1YI6,3[.ad^
NVOP/Lge<g+F+7=92E)SZJXS6=@>9QAcSXGNO,GA4R2Z4(f0]VbBFe2:B_FBTWAH
PR@/@G/S)@7Ic=@BD0cC>35HS?RX1c6&Wa(1ZS:0B0A&P,Vf&]a/RB\-JY84cbG@
/-UbA7)MUBHA-2J0-VFZNO[U8CF[):Q)?>))_:]3XJ8H>.P=Y9SRQ0H5>_T_CZ+,
COf]H6bO2b[.,&\(/>)S?4ZX-b#+DbO8Z-bGWR/OSMB/]5US9AbG9+Ae?b.\g8Xc
8<3(c]A3S+Y,Eb^UY3C(2a-ddVS=;0[d02:1WADf.]6<K)AbB.Y[PU7:)GM&^X5-
^5^d7g&D:\4COg\(#R>Q+0/X<COO5+JF/HE>_;+8bD/LK?=)@gUfO.;]Wbc?,JZ7
Aa.9?=+/P8=@cZ=Q]:Id\@IeB.]CTR[(/UXcF1VcDGC@A\:KAAK\1C+N.@B(&7BI
76U08C<-X6M-RU@X<?V@ZM2,28,:G=4Mc^<5IaA6MCM:F5,L=:B]K,,4[^W<,N_@
Y;CLZNIS?&@64P&VF1A+SCI9ZJQ/RXTTgPIR(7AAL#gC&eG4Y8<3]@7&D0e2+(D0
?#S.3M)&7I_7(EbAe@8ZL2[Vc+;6NV+(d8;4Y-S30>=0QGL;_AL:GB.4=H@M.XW_
LYW8H&PM>IZ[<8Q]L>X4aT(FFQ7T7f)9P2U@HJ3FJ3:_+AINS5&LJOFGca2Y0&gd
H(B&V5A3YTHa4&?LWDNSKSgL_^8a:90ZB?VN(_#B>OQ]dO&[VcgOH^Z)QJ6\+_1Z
M[bJWWK6MRWc)&0M&9e+,Z?TK)#=fM/d=8>Tab\M@M;45?CNXPD.PE-#D_WIXc&K
KY1,6HIZ=8&9[bWf/NTfa7?.4LeGT3(e8BgE3gY^RH-9##d8H6b78+:eH&8HM/Q7
_IUQ3IS4D=UGG<PXHZ2</]^gDRT^MU14L>W#I#a#@:8g2GL3/5<&a42^Yg[YE\^V
H92EJc;-L3^c?dSPB-(V,_N&cFe,XUg7:DZ^VBcMb]C6bALXB+I>a?BV#/@=dZDG
GN=U)5)N&7bOP@SDgXRf;CL89WCPKUU3-^^&2E)Z-eOB:(ga)D<Kaf5;=9]=>KUe
,99WB&+?D@S#\H.4TTW/^=d2aD75MHg@:D:a7aQ5FcX==ggB(f<?UX[QI,(F<=RU
4b,P;M_]:L[g)Db@J_fM=X\?H5f8K7M16-2Q83HA;3/WDVE[K.@?e;]KT?)cDHe&
/O):.6;IZb&AbLUcX-_dU5[f/(QV6K7DPM75,5a@A5V@Q2EGN)\[XJ8UKHeaKb.>
RdRPP<gb75WW^cg&L)W)AP,2GMFCT.[PO-La2]Y-MQJA[VM>^^BgS8M1c^eH@=#V
8?>2O[a__W_-@[6#Z.G]\5E9@O)^B+NfO+WDZKa^(aS/Db#7KS8_5DGZ[Ka2V8(B
.e&f-#gDdVC>PQc]P7418aF25XFS6NSQ6BHZQL3.>5N@)Ic3gC7>6FB(=<HQ0<&6
T6B;_QXKH?LIfH.KO\-I;58f\VfI@#C?NbD7#Pg.g=39a5c-I2T8U),XKbeY0ST\
RdGOd:6.H6/<^IcQ,J-d8:d2M635VI.3g,_VUQR:[3EIef^BWIS<Gfd:H_:b(bK5
3D[&MYgOf/=+fNL)Ia2d3CM(c9?,E[\VGfI6MIREb9cU,RM]9D&@009fDNXgF+4g
IUT;6=;4IN]&.:-@^SgG[Ge-IYL2^F&/)R<bWQ>DKPDD)P:.aT6TC^1aA+O8N524
+I:F5IbC#I^JbaPQN-)WYZ+RLA#b,B283LeX>cI0.0;B^Zg,N+9Fb-&Pc2H2WGS/
T+Ke8+)\2:<_>.^eH]QX0F>b0\:JI:;?Qg5egbZPe>5T@>J;I(IGZZeNU+Mcbee5
YQX2CgROA[ee:TS_F&PBQX2T<ZgU3a-d3bg0MgRSVId9_T/EXC;(Hbe:ae1V?Z2G
JIAGIUH<^0aLKSZ#F3b9;.ga19a<N@9SXgH8;ABB1LFMc8[?9V^^;RD]>M4K^8.+
[N4#3/)FfB?37NaFOQSSU7-D1aD.[^82N9A\.^aAO(:MH1ETWFT^?3X2Jff,bD]#
Og?(WIP176dJ9K/e5.(6MDD+,]/B#D.f6>.Q0ccAIB50L95H3N>IW@bO.YY]:O5>
78-E5KAV=;1+eb_8H[dTgd)?g:4Mg;2L?#A#<2J^EYM<?aJ(3Jfb#b<e[c\eFPAg
-HR<^H\&&^g3^@aN4/d\ODZYbAbVa^/-U1S@cG2I?c/CU<>>;#]^AW7-fVA<=D7V
93(af9H8G-YK6P9/E:^-Q@1[-B#B5Dgg_3=&N8f26ENDf\N2_8e8Z&W<?CP:;++Y
c:T5a1+309A2L1\Y-[0#JKbO0KZ>5UTMN#BWB;+VP+&_b3,HNX7?bFP0CFd;-(,)
Q1.V;B>4VO5dMNX[F.&)7_P4K#H9^0f;THd,CC&.C#4]U@Pf8D[BB+QO0=ZEcIeg
NL)^R3=W1CYXS(6#K-?gX^2&?P,@:T/SZU3.@[PL8AaFUL0COb5@M3QC+5?KbgK&
(O6T>@=;[b@]g8O\bA:\^b=gS<5c/[_<_M5Kc2)SQ4gQ/Qa\d6GK2S5()UF5IKB,
Q(:)5M3;3^6^.BSQfC&93LN27\O.AJ01._DJUd<g>38RCHcMCA>3TJe<?<MN7Q6,
(<T_&IgCKNRSQWA:a4I1N;C,b6U6=U;3&^:_e0YLWd6[3DB]RPAGXSLYS^M];&^T
5\/OJ,[Z?Z;KQ2R:[]V3C?3DMd32D)40Z(e;/f:48UNEQP0g7<Z.=Cc-G&0+T2OY
]>D+VRS_=W+D7:eaZ#39IgEF[G;>I-2DgU5[(E8-A4Yb/&b6&OC<:1<2AQM(8g6+
5J1>&YB4-T?AAWQ/0DGR7(1HL0/0RUL/aa]]&]LEbW:0fe:01+6IcDf675]eU4OF
+P-[J-O?XT9F.P3(8MM\g-cH<7LOC1L=N[XXN>(aSa?#:b:\<]AT/&IW8=PE[3#I
?8W((UM8TDGX9LVafU[b;aJL<Nc1L;#/G8&gfW@Y)&WX@(GJ/F8(gGdN^F)56g1A
VBD<(A6<_e<A-]HM:QFa9cg4(I6eL7EZ1a[H0RC5FY<W[f4G5)RPD37XUcEFg\L@
aU=>=d7acd+)ce&M]]55>gW[?_SMM&6,3I08>7^/E1B(f+PP/3^L3A2Mb46(OLL6
&1QOS]-APHa(/f_HJ>HOf8f^)OGK^7R]79eDAT[_<,5X.5^L_-DK(&+L0b/38WP@
e.5IK7B^,ZY@]9<C[>c1A\-E.28b=PTUS],K7T\Bc#5_2MSS-ZPOT\5?R[HAD+-c
0[T.[6+Pd#04W,EYZO&M:=2K+f<NAXF;dbR.Q76R/G_]HIf):^<8O9<W)C?6EMOZ
R(Y]S>F6E)2b@3Q7U<BK.X_01&f175=-_]:.dd>JDM8b<+C@?b_AWR>F[]I:?=2f
33CFV[Yd(DT68_ea7P-L-\,fK@1K1;XL0CNaY6=?^__8fF5MHK<N[^DOWE<>6V3d
VU.E;Sf-+RVO8W<]]YD#g8LTO+Y/GGIc<TN20Ha8eO50D36(2OBHK@e.6&I[93_/
1--@57OeM.NS,5e:FeXHFePTfZ0>_QMf?7d)UKMIBN7#Q=,](/[TLLK]P@=9HP)>
VYQZ8R#HXJ)c^VeLZL7D:g0]WW76f>:);gMbI4&3V)RJ=3B,bTU:>DKgg,YWG[\^
6\8CgK@@)SaP<#]AeRN.#L+M5[RM[Zg0V)M<_#(a0a56&0AR&Q#[)?VH?)HIV;b#
<18,=(HB;6TVX:AaKN]QgE6A&G7Nd/g4[(K?bXLg+c5LK\a50gA&+.\Bf>X?V([V
AL_HY:fQ3PdV);6a&;RPbF6R\g0>H<:G[P)P;-eF:b;H@=H]gNg(S;T2Y]^]N149
SLRJ\RH\&:2[VC\NFFSc)&7F.Y5Ob.J45E)KeV@ZQ4\@,/2dd)X-#V198CHT/:SM
D1E5R&R-^e/+E[^&@H:Xb66a6?FY<G:dHe#EDV9),<T]T#^F&dMPSP\g0>@BSKb\
ZKF@ML3UEEc?#=d4]MJ/??Ca[_c#N[N1cT]D16UX@7/e9cR5]<E,bO&dB7dLW2=W
b;D8LUV,J#a#+K0DU>]93:Q)OHaU&/OI88f12D^\?6>F59WOKQ]b5^#a7<CJW+;N
ZRO]ZWW/36aO6BIb]N5a=-:6<7JFF)QVgbT=U1g[^36=\1gARQ6-fe:6MF^[U7b<
&AYEYE8g>93^K00Q(c;0c[2506GGW#b.GI]KfT4[7@LVVY1^1:D+B4IaEO=aFD4:
VBHZg,L>IVD,T:EM6Gd>C?2+>L#<^&RH]LFWKSbISTX8;98#HJ569RBcdRPKBGT9
#N=X@aI60I/+HFQ.[7ST&^JFSIQKD<K9P]=F[Z3bYd79&+TG?8GEDa&e_KNSg=XG
5-1=c+_/&GQ?4&GQSC,\ODLQ39GAK??^F?7-DHB.U<V1YYZ:TJ(aLNJ9/gU>QN(<
[5^B#LIOY(d5HK23D>I+]SX2K^E:\8;@+\SKKB&0@YJVe(;-H3Q(>PAc6J#5^.QZ
Of+?2IEJdZ.]T]W[&;^41a,;3A8C4VFI=d;MW27=/eAGLB\PRC7b+0aMXSeXBYDL
+-4@_&O((1&LL0]TRe/<PVDV&ZbCI)&H08R86QJ:4[CdXbF-&3dF]C,8e8+EA[3G
a:NSM,9Q1N4d\ONR1E^368TAXHICU5?2,Sc8TYOS4MVWE9<_=LDgTVAeGD;Af15/
;ISS2:]\XK^(H?.^Z<JDZV1bdSUQ/b\9C;(-YgZ054#@eP1cE_TLa_I^LWXL7e9f
Lf:f7)H3-V5Ya=,0E^87[A#aOLT,VY@)J7;M]R/K5_1^F_A&E0MILgT_F^PLgDd)
X6:IC>N@KN)6Wg.MY;E#Cc21X9+;-a=G^.X)\>E8[#/O+]YfB#66)L<Z;@WF7/#^
P</[KR&;#.:72[]2LQ0ObLA9A(P(OGa43Q1D,EA&WM82K,^9CdD3\.@]20e#D4R:
NLO?V;DRDfTLebTTNMN#-Q^T9gK2.#/1#&UFY[MRQ#HLZB,?>A]JP^X>&?a(Mc3=
#+aad9b[V,-U,TAR.2+f(IFIT8&RX+:HF<4;W2<GD,K9b9g:fL8eWa5++R5-1?+X
3B[PO#S[92c[LE<eMJC@_/V:+8[^K.[-C@+dK>HR1NS5-4+4.DcD56C;c5@J[,T,
#^;#^LS#HW:;Tdc,N7.T:4^\\g(;Qbd[P3<RI3,):WCFcXaff-e_^<N4aMM_1&,8
dDaN8T+TL_9C^A_VUH.[:./3,aV?B:e2bdKD;Z&_D#CO=>36:O,0X.aTbYY+dGSg
6YD6AZ/RcS89K.IQUKH0C)eNXQX=MbLJ:<7S\HY7L(.]O#)7a_ROF+H6NBF557<)
6A\BL+?AYR6YfFe^ANFI)2>Paa(7)fHI=?eM4MA>f/\B48?Y-&6[eR&EMggJJA5>
eN?Q7Va>RCF=I&<UAf^J_C[?>VTVdQ^-VKHI&1ZH,\/5D30PA(#3Q;92S?[3]6D6
U&?7EbI9:E-&1O80</C<^LZPMa[)fXGBR-T@)^cKaTZ]?W<B.6>ZgP1RHTa7JZXW
WN(#=+FZ?FIe6-a_\eY#O8LE5=7O<QDIYDc+5,&:e@F_3H5-Sgcg42=Mf6HLIZc?
b3JN8V_7_.[VZO1O7#YVA,#K+-.7UDL?S_^dZP5;8=5D+,->WA)IAOC/:S<+;I3Q
<^6^VX<C;)?,g]?,cL9</WB3-aF,KUZQ0H4@eIJXRJ<c&HQ83KfQ0P[cb<c@XH^Q
2[58J=7:IDY&U:=K@f?Z13A:PQ5@9D>f=5=&J+^62HPSX=R?AGM6K6Q^ZWMfNF]3
,T?4I=?2G;M^S,E1:bNeCQO2MdgCA)6;EN]@Q]:cE4Z_FN-cVaa+2eDH;@F=0#<1
(,dZY7/4:R?Z-HW5DYW@O[,6cQ/..Vge(-&a?B#e76,If0-a^&[UWaXcI@&)OXJG
/O(X^F0E&(b76<=&W)?,LL.GBge-0VTNCL>\TZJ@_1E>)]TW@+^?/NS]\TDEV@_Q
D<d8AZPa,gbZ7:9&Xg(W&G61M7MQ=20f4;&^T+JA-I)J+&eQ?Of6-])/YFJ,0(9+
bJ;)QR8MCOHRf>Ad0&D=K[8#(g\P3[A\0BAVP7cKU_7#fc]^]V0@#L0/6-GKRF\(
T[H1dc=(#3M;F8?>^Y\=KI,0Bc]Sga0+66Z^LfXJN?V^ef)YXM()V6)<a@/N^Ta/
OYH&,[BQY;SCC9?\H_>c\NK>_a@OF[44@CYGM;UV.?G.7\P.1,cf4#Be.eYP9R0&
2M2ON/UHSIf80ZVX8V[Z8LJSO=3X#ZDb=fN1?BDD87L.-,([#;Y+MC>X/2EJg\J;
_MGV9?adHd5BKMGSY57X&bDVPAUMUO#P93Oa1#W/X15b+J\Z+02M;L..?,F5@EfH
886>D>G=1-(4VM6C(EX9&=&aFD6E:TD<[=;aH^P\LV(9E0/?Bf/V]IG&YH(1f&NF
QFPSAP</c&[SS\G5AF@D^OS>>P)(L7@&/f0,&R#T:[W/CX:2d3QeO<B=J,6NFdB=
T<)eV;fUKKPcMR(4DO+ZDX2R#&gNQ#IDf1?8,+-1&6Z5]RB3]2aO1\]b+U/0@/eM
&,72)[8af<1X^cM/-M_3SUd/X_[N]+9]0M4-5_Q[:11#[F>6&NP,A)WDLR^-g[,V
Wfc2/5=N<L]MIfR+c2L9+ID57P<_T&\.-ae:&^,T>)[bGZc+<dVOX-+<5\S;=^8d
e)+-OL;ZcA7#-52,JCEX)T<TN4)M9B.-@S:KUS/?bNI].(R\bTf[QTA8cQU[E2J@
.U8I3]#W^G]T+d:-P>??/F#J>\aa5JW^K,-QG9]a4,2#6P?EQRbVGJJC5PcU>D7c
0aO6\2gQ>3QIcP-(XQd]^B6#C5[RMI(T9e1X+21:2]6EZ)e6D])YJ]6SeFfXg<2?
\@IdZfE5.E<SA.1^52+?-8A4;d_;(OXfX;1)TQTYFag^:_f<272fV(0;;8#a?J26
>8)0K>>WLLE#7Gb)I?M8Y>G;->(aW?HAN(H&3SJ5O/.T5eJDePd5Rc#7./]C)=/7
/PYM5J4RQR?E#Cd4JRe.357U)^+=CO:a^Ac6P-:PUMd^(X=G7\E9fL?0e/EJY#5.
#OHXCTKV&JTEKYLB8HP-6[50(;(I4Z5#^X/9=c:-V(,Wb[:CX<EYG@dcD#?SY7?.
9R?F-,#&E+B5e#]g/R:I#7VPC;]FP2EUeg>T4La^#=aE2V=HM?_G5CSYCU8J#,XB
1:1.5cSZGb,W4I0#P,RN<P@I3@7aAd5_R9)0J(aBQE9.3+<;Qe-UD_HZ7&0e;LL<
7e]ZUVW2SEX_KB=;08.1)d16c_H));KR[(VLWUT0Sgg@T<FE:6I)N9#/0_BdCF\Q
QDRGCegTP+A/:_Y#2\+OH5LT\Dge8ZJBKPYeb,_?-f#&[dR=,eeW?8YeCA7aPF-)
Z7/QJH2;8H2&2+K2G3AUdP08P-2bBC3=LTAO<7;YbUe[60eIH@Q_UPK.O]&B9>]d
2c]3>&aDcMHf<D@+?;)92W<H1]3+SNW@c=.I84Q4AG^AE\UR4[&:C/ERYTY:G,R-
O9=MO@L,=Q>JPRJCL8DOP9-:2Z2_#5d,fZOZWCW(#D]E<6]ZKRE3ZLA/16c3<:GO
EEdd@dXQaA9KQ6C=1DCKZfZ5TMH[Mg?KP)TR#)_;YEe@O?V8e=7eNRP-OQE:B0(3
&PX^NMAERAEKNANO18</H?dXPXg8_:98_^E.:I2\C)&D5/->-_L+8,I/\))b<HfE
<8HDJQZ6&A0C?RGS)_KLTCB,G/S9AB#gUJS)+gCgdDKaWVL7:XPJBHd-5A13eVD)
Rb)TO^VS5:@<&VPD@d:00bH(:IcfS\7/#<V[Vg8&d&LPJa0=XZZgYN05HaQgNfYH
([bJLFedMg-Q?LdU^7VNU:V5?L7AD=;0#QX76JBBMZFYF.61e-[.(1@G>OLcW)CG
>eB/J2U@XV[&Z@;)MY45Ec.KY:HW.cMPB6=If)abb5JZ)\ceSX1,4&1K<()#FIa5
6UKZ<DSET75cXO@Mb]K@92ZBRDT9CU./P\af=KA4>/T9)\2^BXN[:B=7I#a22Bge
FI<Q<-Z)@HG)Z+H4;/86d=.Y+/O:PLILPN9;=6Y&gIQ8W#gF4D)A7bTC315^\Re&
OcO3G]1237:SB3H>6:IZJ3/@[@ISQcMcYNQYdQ)B(N]3CZILdZcCI.6],R86K^[&
]bG#\f=@G3NNf_G<V<2NK?+.=E(dP](1NRg4c,9YF3-a5d1MW;#Q1;4)X(^R^PS-
=>gMT=-aX]I5V\Z5Zd+F<7\<-g:(Q7A._3Z:759;?&(@6KObb4-EMg]X#R5]YS=X
T;5N1D]R3QA,Q@OIg[@M+A5&T7^]b(@H&.OgM^:;DG8Y[3;<L3D7a<#Wc(b+3GCH
I-\f[>BQZcU>aX;Ce?Ja>4)cP/Q0g]3d=VM7gHbG8#M4=(KM)S@A@G&Bg@7A&c=@
1bM^PJ9_d4SS.4C-(Lf/QBAH8-DA9VGRHOc:Te&TY5+[ac:OK;#A.b(+6^I6A4-H
8;0Y?TSHHY:51f)5\aaQU7WLX5FRKG7B2_.=-D3b0E>+@5a[8ZcA(^PUL3)RJaXS
(,c#LR^EB5PFd=eH:S\=-@\CC2H_-)@I(#[#EAf\<@#5\/Y\LPGD&OYQTY?F94H\
H6TO_<>ff?88c?^Oe0P(C>P8:Z-;IEY@N<GM?(b3R_b=4P9\:O>TBH&ECgUR<D&6
,]S:cYJ11H#KSG>,5Dd(S(&][B:>=T9VZ4YU50gC-Se]9;aC>A<3D@P=QN3>U)63
:H?cLR0XaBa7S>[5O+VUVFcb<E&]Z1MIO6/YKL,8]C@HTLe3N:6PO&Bb0BXWeBLB
cR/6GRN^N(d[@5Q;<LH/K=_H<a;Z,J+c(A\U.g5>Bd7H1NK:N0&4A@T.8A5;\O==
e=_[KGA(4,bP>K4D-=O2^_/>&HGNYQY?R/#9.U5^+[H@<O&A(eRWC<(d,gcfLZQ[
.Q7NGY9K,./6J@IA)8LIZQ\aYDa_a+c_Gg[3AOF5L(3OIWd&R(YMcM._:K]P=-f4
STZJ((4a5/aAAG+P>c?SEA6Q/2Ma1@Z13,@D?@8aBH=R99XC[W-EgN?FWNc)BefK
Yc<^+8W]ONE8WN>4+.IJG,\[DB<e>(c6S_Ud)Z:A=9GHUS,(e;A7_=9B@[RM(Rb6
Ca2C:[Q7BTb3_bc90VZ3df#cR1MK6[N^/US=KaE5/Fc_S8dA#dEa,/MB,RPdJ5&-
;a_SS<DTabdB=?B8e[BN)9OI_W^V^be=>H17IQdB/DX:-]J[,>:#)?0c0T7#GA:Q
CcL_eG30PH:65P]#A01dMM[0DZg^+>RO0H5b34OMJ1N_Og_9;/SBP?DZXS+L&6bV
Qf4;FO/GV_>A-2&)DW7:26S?c\d#a,U-9FP:/@]Ha(LHMfAM\OI=\Z./(d49P_=]
A(fFdAgH=-I6(((5>-YS<L(:T4(b5PSb_#Y]CQeHWD8LO[?_@-T+G8+80]8;@-S\
feB9[SMeH;Z&EUJPX;>c7\a<M1_Bc4J;7O#@7_M3&1_;aTcAgB9.S,FNQNP9]1gR
_64#ITFbF,/.fQIS^NS1CC8L3ge+RHO_:J?2>bG3FZ=WSHHBM3b^WT;6.7(4<c46
7&C+;bKC23+L?M#.c^?5dE:-a[KK)JR=3Lc?X23ab]]VObA3[6[NO&J.^>c/>,G^
C>W,4=4Y,+]bPFWLJJdOEfSFKD&P5T7CL]Lc#I4016O;SX:IL.PGO0GSTb[T0\(L
E+(c7B#NaW_b#SMONKI(F7,=K/_7VI3Va-S>1LUf3WTPNQ(:=?CIBTII^?55&(0M
[S,)Y?g8:\D2P1@JNF)ZO2V+,M4MSb#?_]BE[^]TI3<PSR=W)(&OQYC(ec64aVf[
e)UW]MC]bSI\MYD_?V:3C4&KG^GIdcPJW7?gL>0f,ae)H5bH1+IgS&gS>6EAL>J9
4S&V17JL32@FbR.9XZW.E]]=H<MJ9TY&@N;:7K6O-U0.b[F7\0NN+\CZ&=8W#7Y@
.)Ic.#E[Ub#5eI9c^,+C_2#_+SPGcHag@BagAT\TF:MUI01#]0JJD/QF\9)<LGfH
5gX^&fD59\HZ?7>VObVV:WD@I[5,=SYVZ5gS&9,G,T[1?eCL1/(L>W17GaBg-W[\
C#,UXa7Lb7egK?(8Fb>^aS:35_+S^<<5]_JQVK+d_d6@2D-<S[XR]I:bZJ?)9P_R
/],5W1#GTH&6D:#CE=Kg/R8@4@,3]2c8Q\W3QYF9F3/H4]dXRRSOZf>cC>671)I3
,YXcd((-\UZg/]-KNR_K.:Adc;I[84D(U7:ZCHfEX2(WY;BBBR_SbCY9=/_W7MX:
d9UcK\55K7T7STGU+^b(=BPDJQcdb1Q#P3=XY<NKBMgJW?6&?_cXRSV6LVVZJ[QE
d)1\&I;b3(H2T.WgG[S@[MC@MEd->WXYdELX/+?R&B.1:SEFC=W^_/TW[C=G9\I1
(Q.Xc&F3[+RGANDU[JERMAcOdFRg^N7LRE3BgM;),(W6,c1ZK,L1>15E#g8aISR1
H]e^F3=NF@a_G60IPfRW>\>#)9^NKS-L[^K7Q=YM]WYLGf11P0\B,TT-0Vf^-V7\
WHSX]bC,J_(81DRE0-]?8,1(e+Cf>4SbR)^]c4MD18RcNP&g]BIUE::DS+Ze@8\X
8F=]EJ+-c4DAfedK(DEO>W<,g;Y0#)1aeC_/BD.=d#YD7):fJSB&Yg+OI5e75dPO
@MH7,(cT@(Z6Ka57P]T+[gFYg.,,9K/NQ3g&@W)37d;)W32B^&/VbEUf0)QV&@J1
-L=-P[-ZffJ=Z=9MeBSNQ0<7O)[Ia[LXE?K_=..QC6I4:2,;@VH<f(aFEB+&)\e?
,1VWbVg=gOf]Y,5D\D?]K&OcZ/9[A\^80#1,70^:O)NKdI@ITBfENT6BfNBcYCVf
X<Q2WWYYK)QI4B3D)=>N8KE53.Qc[YVV>05/XZC]5J5UWZ8[R,P\YFb)B1+g+f;>
]XI9Ye4BU]=JL&S=aW=>X)9HTES;H_faLF\F3Me=QC@^G8XMJ_9-,Ae9OG;JI#S2
VEL4FG#3/?<L08LHJ1@B5)8=BcA+gQKZ2(-cP?c2Z-S8H[\PUW#WL^3Q[cPWVN&K
0Ra2<_HD#,U&5.Ne&f[#SSL^Q=W0/,=BI4IgIeVXX.\5GbK+2PCcAbW\6SDF;G_f
U]-J@f0bD]7S#5Cdg@96.-L(VGY9^@BJ9Cc:(BJAWVS&3TWD[(P7.M1Z>5&KfD#X
b=4.4fT_7V8X+L@5,&a.)CLN__+TFK)OG#J0.SfP><Z2)KfT3d30D0F5-6^QaaNa
9YH=cJ2X.SSe)<04RSMS#U..Q,SMaE5K(H;)#<L_^7aUf(I)HGdVW8)D1IFAg:N4
.Wb>Q7GN5+SK-7[G,X/FWdC9e;VfS+dK_=8D-NG6gbJQ&cb[__(SDaC5@MF;#&8I
YH1g;TVY<P3#]3HW3OUgPNYU]>-NR]LadV=g<HcX^[?HS?YT^[LB\VEMA7&<ae1R
3YTG1OHfefV[W;a><U@:9I1dT<P#UecJ5X+/8<(_d.0VfEH^.E72U=)7NC2>MZK6
CVJ5W.Od,QL2QP)8HTef4I&>U-]=dNBJY#LVTG#&Y&D+PV9NWWIY(NNONHdG;7<F
eR//&X:TX]E,&>Z#7+<,06TV1_3\)+@OG6J0(HZB<c2.AJ-5eUg.W\5=e)?65IVZ
:VMUdV:/g25V-^b.eAPG>HF+/TY^&4dTR\b._]0Z,F4f1eGW<<#/-F/H(^S(S;:0
eV)P7945R;A5G1b&)#<UPDL\5L4.TeS=K?dG,a#gBD/fY(/_D/eP._5>RM0E)Fg[
3:54@[L27MB0Z<gOU^71/POaTNW\ME[3ZW+BQ=#?2/8_>YDFAK(R55=3FRJ3V;>C
)dUK:d[)#WgZACS;fQf>G(AL[)8F<W[]H_beZ^<dGV76X(dHdM1S\,7#6J:c)bD?
TM@XSE389#E8^aS9MP8OV-J-c.g2ge+f0>/X9IbgX8BXQC,?/c-\J6V2eO\EU3_E
IU>RVVI+T&(eGT<bWN#G?QPfe>>GSAB8(#]5CN_8.YgHFEdWcQJFK0dc/GP-C[]X
CIT83LVBf89a]7.&5-RYR9R^8\D7@.<dQ:2bFO^d+<:B<XeWIfOVE-bP5WU6^3<I
Rf8#cFOJ8^P;]A79Q4^)XII]A6M0<?^?BF[KEZc1NE/S7XTa]G(ZLgQ7KV_UF0E5
>b6(7bG+[\U^;T_R8ICd+6KeaE=PQ\g_bA88c#^CQ8-,7##JG8[Edd4:2:WRR7BS
G_WgS/O.-#)[X&bc[PC(37,EX^;]^/G)Nc5HOZX)7.>GY(cDQZXUT0b]YL+.JTV6
W_N=d:d]SP;R]=15UL7,^Vf_Q6^Sa7>@E-gf5fC=+ON>&V>d2(/AdO1)Df+V).:A
C5_/M5@D\&JfR+I-R3?8G]6>E-8S\<[a<Y)G=XV/G5EDPRKF]4[&B(25_7I<c\c(
/gZEW.@466OCL5^]eM@WWTg9B^M0DRU00HP6:eg&H:=G;M>-WIC=:,WKM9/CMLD5
W+QA-g9C/4aBPU>2(?KDMN<a&(&TRWTPSd<e]+]fH4X/O8DH[G@<?2BYMBT^#[4N
eN?&ZH=_5-HUHQc)8WOfSNQ1cLI/RE)?T91]D8f[<\@YKc079PaEA<A^_Z/gdZMS
Q]JcO6H4YeDc;NJge<JOB;,8=[NSO(YB5=0W(SeEaKW,0W)cF.f<6bc@,eU6=):(
QE;MV)7bWaS6F2H0P]BP2R>[a0#TUQ(+A4.3+AD(/S-.#[9?HIF)W+6Q+&&.:SBG
MCG.S>]<SSc7>P<7dCCS0)+3-X9>Z\I_19:DBC&VK[&I^T-RS?#.b)DE#K2@E>0N
/e)/a>eFC]bWTd[\ZHBJK61G5IE+M,@Fc4P(6dS,QW2J@2dE1+XZ/2#4.?HR>P65
Q3?R:g8V9^.V@0IT@J0(#-0;PeY,15VY,P2(RNT8^6W@C_a.1T-d/N0=M]3e>B>A
1ZA\N<Z54]S=0#I=MARHF^bJ#9R,TDO+gccS--&_0g8=AN8A3)]bKRBNL5MU=5=/
[BAV/I2=IC9F37;3bI6P35,MS@E;e8UaI=,B0+@_BGF5OZ\b\7fX.=TN)04]+0DR
ZWE;[b,6=_YBgWe21S.2G4L)UJN-EbF@3&O@(/?([Ba+/efg7:MQ:1<,.B@]Cbg+
)ga](eY;G5C8[3g1,_\WKZLe,:KNB3ZIe0T)7D>#^;.Zg=QV6W^<P5K#K+EYc[\8
=,Lg52/2/.VSfQHS\IATA1:0GEK&a3D(cRS:@6=Wg[b_F?P;Q18F7PESV<P8gMeP
K=.Qc9bKTD==+RK+bT18#eP]P>f2C?BT:6WFSYgCe6=3_Kd[=<Q:af7J3W.+AV7R
Bb(JGag9O.Rb^H\SJgfgLBU]A+_&-_/Y2PA8<Sf]:<I^JP>3+#>I\]6H(MUVMCf+
[Y(AVDC-NV/15;A>eJ34-4:XJO90Gg-5O(R;FE@#[[L\#+:=KJGTJ]>H:J]d4DOR
TU.^ON=g/S,I-WKgT3-N7/4A?=b^+8G-RFMV09CJ?H_UgP_<Sd(,G,_]P>)IGc15
)&Nc;+Lb=\)33JPG]<1-W=&5@M^80bS5N)@#JOaOEAg@cK::LaOKBP#/GZ/_CWe(
2aZ[+973MU^ADXRZT99_L\)&\\O/)K#WIBaWNAK:EJO6c.fd5fLP#6(#]+Xd/-Y?
ZEe<Q(4N5UVc7FD1X&&Vb74CW7NFTIcB^>@9[V-A,HLF0?]B8XHX1<B^D=LUQZ[0
M_X2/FbLf9a(O<)eWVDMRV54[5QVP-Z>eI::T)f6:_;BSD4M;6f\916H28<XU<S@
SZ5-V_/A1V#,aAJ&1@.-,DOFREZT4ETfH#\)_ZQQQ?\T^3G=F1&1Z/P^1ebK/)?:
=H33/@XR=XZ&g-)e.Sb6(6e,;gVX<V5_3#RXOJLG;=?Q,Z02V#7Z8^3=(7_9C_;U
G7+dM2YbXRH/;1J:)00#S73L9B0;9UX^1\LYCXIRN_)A&V8.>PJ.EHT+1]E70Aa?
J^?+Nb\,8H_3eEL1##T8g9EZ&#8Af4_A:.5?L4#^F+B3K#a;&R7V5>7[--IB_M;B
>Z(VCVf5Z@F]>d?\[2aTf^;7FH^]R/eRQ@\P=GZA2+GX<NM]>_bN8gR^V&f8>(+I
dAdO+b>.M<8W#@0O2#aOE@7gQcIS>IA8;8[f56_M][If-J3OdFadZVO\6NaXIEc8
8VR;B^,JX6OW4>2->3T;4;b\2OMEABEQdCY\DfT8b?&KcUO5QAS/e0KAP@)EF)5H
FN\XAGb):(X.,JXN>)^PNW4SJC^2\fI0OaJ9EXW]+4(,H+X5).g8RCO3E9#&//.B
638gXda9@R;bA#UB-88+Q;^9JFBg+?UZMPHDTf-90Z,3B&\^DW/8FaSM6?36A/6C
E:&e3Y3RfW3DGb])Y79<g3g)PMe.M#PN]/c:@HWbMC<IU]KNEOD2AXJUL81427(Z
-6Z22PC73J)4H)__;244Ag/2.@^/A0S<dY0([9f>TV[0;9DIPW=4EKEM.g;N38<(
W3)Xe?R^Af=<VUL14<LT]LKHFd&cPMR]10D2+>?(+4E5eYAQ<K\>KSHDN1O^@5dC
2\5]0VN0,:[@^2^502bgQ9+\Q7dE/3(@9U#Z)J=VAd0YSFK&B]\fU1#IReXQ][@6
Y@f=dLcR3GXDb6?ZRR-+RQ2FV(SVYdM[B,CQ4U?aa?C;#W_EX7e9+]\;:dCUY9Y;
bY)G34@aaU5L_99[Q/;5FN)/Zdcgc.V]0]:CKK^bG@fY@M0aeea-^3:.G[aF&DJO
I\3Xe@+1OUJFCGF#GW_5)R-=HX,K/CS+L/II3VQ_Q:b[3]ed^5eMgf60A9f0RN@^
0^NB9[6URFbYI.[B#agGe<N6KaTDESL#4a[T[XT_a0<SS.>ID9<g&bIM&;,FIN1>
W><YP<B05(,>?PKOV4X1X\Y_7N+-2Q].AHgU+PH)NbLN+.DUeP9eJIRU56(=V:4[
gc5eVRK(R(B>Q=HB\c;3MO?9fH^_S#;\,:#G8BKMZ)RKYHS;O84O0LK,(@]IX?Zd
O&DP>[Q,fMR<M4CXf5:6B7ME#(dP41\(ERd(UBT)aY)Jb&e[ad.<]:9e3-9QMU0Z
a[XG0:N.bS#&NH3c?L&E;>baS\&dCEO&ZXK-OUKgcPQ5[IM?9/L(+I:3?2&fL+75
BHG^g\,+^^M76OL@(MB3I2QQ^QJ2.BX8?U9,:5G-0#=g1#N+B1XZUR^C1E=]O_CQ
6.?g&@-SS6XOT.g2HG=G^J&A),UVVD1P[@5aZ9dP2cB?8QWcX9)dCGTX.I^:c^;e
5/QN+[IMRW^/+[M:e+cCgBFBT.@(-0d&fd>44##+[X?GU1IgKMg(S,g\gBGgGL1S
QVK,\<O/5+(UL6&R3E;M<0aK_]6A#IOg#VIU2G#:_I_K+aET@d[XE_dAJOF<D^Lb
0=<D:\_IA?ZBA1BEd[<Z4Y+cRb=OS_C4#XCI?e@UMC;7(MD46;@WR9UN#eF[G7?F
TITDUI)bL_[9cM;A4eDPf+TP@c-/8E-I@[4]LL-eJ:BT(VP>77:/1;+@Ma6#[AAI
M_2@)=V^I>He;c:65<YC1gA3JDDH#]_>OWV]eGR#X2\_BDCMB8^_PC/V)dR<4KL^
@gA@0SIK2H.W8I^VI<I)=NZP2=3RYcgN()#5^=cREG4,IIZ_A5CaAG(LP83I?R#L
cSI8Z)?Z]9(.NH_LN\VXX<d[SY;eTe16HD68bWLa-0)WP\[P;-M@(bUaJ1M9.:ZI
IM@+[0LfcVWP3>Gc=[-Yf=P;-CITXB:\(aSSML/PaT59S(CN3,J_@YXIPJb=V/1-
G:1a=@3:3I<HGW#OEWGQPdD>-\b:JA=UFC>[N9fca(We#b5]CdPFRT:d5APIWS^G
@dBc+DI.6QNKb/2U=<d@#J#+Yd6=)<:W;Hg/?32G5X2O131^+L,[^XH0Yag=)</3
-N-7FEg@C2B3_^-d+aX6N@L#>0:Y/+&3b^/GU:D+eVB?KV^-fZZ5:cL#MG4?/,\>
MAX,dPVf(EQTV&IcD><[M<<P.YaBLXfZ9.,H_LcL(L#_3W2EBWH>/>85d8bcG40K
_5Rc9CASITJRN?Z?.-]>ag.5>O\)M#E)U)5J0f#I3DGH[]&XQe=I?0HC>13=SO)C
I2dW)aS=55^CF1\cJF.S;/\\?/[OZQZ7/S)TSZJ__f_)02-3K#:T\=gc7D:9.#)C
+W+R;KA4JMX@AI.9_TBX]geWTDD]+4CO9QgfQC9J@F^]&629V<HfP01[9[R&f?Gb
g4-YHU[/DI-RP)=P/NeBCRX8RD1c5g,&[\4JO2Q3E+KTd(^#[-BFN.<+F<X>;LaL
W^d@5PX?=/=6.R<KOI77WA+C:=gf5D)KY)8,D/GF>UcV<a+L3JHWWO3UM><1e=Dg
O#)8TaXJT5D)GOM1Ug>05Rb#^G,0,?9;O1;L62=,W/=BF)gFd&U>(Cd;(.GD/\5Z
&8gVR6Y]9BD=MggLLMT+J^O8NE3#PdeIH>T5)aHa69D\+:6E.)e9-:FD#<+c2#7_
gU6=g84I8SCSZ#R_Z1e9@:d&GO]0=;L:/R)^AIAGC2]<N-X5&)2AT:<&3UD[#6C8
GBU93)ZO[<P8E#6dTLIg58W4MBC(<HeP?dC(QR#Pg-2R@E&(@AF/VO4E[M:,[0FV
Ye(3=-2XB+)C^24_KO_.K:_-^0A[5ABKY3]_>&>SA1;W@SY/^V)S>+_FcY.f&/X7
WQG?C7K5RKTP0)#6a34XNZ+&d_I61f&;??;E^c(TH[aZXK.K7_aI6D[_41d]EbH/
ZKC@-^I>=Tbd062OE;eMOa0G\[U95S0_:\Rg^GPJeQb-dTfa:)^4M+._;[.6J1Ug
9J7174]#6=g4JX==6?,23]J&HKZaN]O)R;M1Y^&4g+-&J_\fL__HD/9+;#fK7E_^
JWCd&-)\I^7.7K]6RDDDMAVTcQ-45AIC?SZ2&D?bdH\=6fVG/;6QZfR8^N=V\,AF
OX-5G.5TLa_@Z\bFHfK9-?(;a2BRXWCQRbLA4WLYZM@O@U[=Lg<<S_DcT536WGEd
DC_@8.bYZ[CKLBRYcN3Y=X7>+YSZS[R6=(#W8LLITS2fA?GRFZN-P0(7@?RD7MGV
0Q,-a5VB8\U1HaQ0e@O^)IIXbC=5[[)<(]SV^MeMQ]P\<LS<[aQ?M[Z7YHFH1,Y8
3TW,Lf\CT<BU<KT;[7/Ld=EK+QJbF\:78b&8;RG.:SQKQ@HX?g1Oc?_L-cbZEAHX
NRI&OPJAe[]\Z4^R61b=\?]4AZ(_^6f]ZacMHH3)+aG7L&+;6:C\6-&g<1U85Me6
;#XZFWQaWV[.Q>V0fgB^:>B]7G1HZ\]BX98M8Wg([-:e/M_RHG,F/7TDd]=57S2+
QS=VI-ZL6KE/cB=DfS]&YB_8+[.[F-\1BdOIfY+^3)^LJNTJDIfRO);c&NY3O4a.
8?S/?W#-8[2HMD308Ncg[PJ(;\I2\;^aDcWSfIGO[29HFIT7A<-]3)G>0e:EEHbC
J.e.;Zf#J90[3#PX&H>7/=2<U-S<=8.FOL=V2H,=[M>d50e?=_@DbD2B=3+O74=Z
U]MDB696U+G4#c^T8W@?,10IE7(5.^:DS)KXW)6A7KQT5)<&4C)b#3S4SbPQcXe0
E9PgLFTM-Z&^1^F191BXLO?<,QR(N&2)X4W\a(D@@D9IC#2[bYH/.+0E(JJ0)?^0
DG]2ScUeJ+cT&4TD;,\]N@>7AdK:JG0.2NKYaZ2b]=<:^<CX2/G)N<cc2M]=gA:8
X,E7&>&YcNGgg^:XWX_BeV@A13)P#/^39[SH<Y,3^117Y(G)RF6-#E[QG&aYI_Ae
E#HKZ+Ye;18-aFeP?Yc186,4c.dL<9[_^<&;=f5.N\KU55FG(B6d6.^>RW+?QU\F
[dTRH?FXA(+YeGf@4@W;@3J2Y7)=A)3UA^=[KfG3@:75,b2#Y)QD+?>+=ZU14?U.
BK6XAM)_K<1/,d1G<JKTQYG_EB:>Y+T>eHf\@0_Dc;#+3(e05Q&8=d7>.9^0ffMG
ceS<N6W8,S\@cK=4G1775EL:KCJBHQ&8NQU1=&(gD3@4<J?>@,#YKY>/#+P;M6-8
?OFBaSB&9)&YJA#M3FMPLSA#=cL\GcT>3@8M?,Kf2^P=DZIMU?KaESOe-CfG#IXZ
FBN7:1BEH;23ENQU@0^].c>&c5FMPE10^:U&VF)19J#(FHI;3^F42Gad7c.[\0a+
@dKQ7eM3J5c5UYU;),f15Ve48CJ-7/=CYEb9S,32a]6LU66S\\TZce+F9R>AN[.H
UGI@<)C)=E?DQREe#)e@LdV8D_X4JMW7/@HJGB[Hb3aQH7fB@-)Q,GO?XPb#RaPb
W+UIC[RJ=M&;8gO^W#&1)gZWL26NMP)b5Da+5))_USUO.]]V99H]73;XLc@2bTCg
,bFf88?A]YPY6TN_K.M3XHS\B3D=[QX^^LCG?4NX)2C(RYXB^4.:3TG2534.V#>-
gdW#=FO17=-\J^d&4a=@:?_c06[:HPZ\G-a4)LI;;OE8,)d=HMaHJWJ>6<=GMGeR
=C5_J&0_Ka:(+Q)44ZKa&WMK>\<R41bM^?XcF)g^e4FZ\FA.Tf12&^1+3([_L/g>
RR[L8A4/_UT+&<LC0CKR6De7;C8^/V)8SK67XS[Y+RROg9:DS=@DcdX171M3TPF[
^N^.]>L\R@-RPNKQ-Ma(;W::;Ja+EbI&:=Z]0=7IT&O1N/[(Wf>d^AY+U;O>NJ8O
dLJ]9-)&P]N@.>f-H[?E@f+<LMYP_gWYM;\(UI]>E3.>\U5TIN#.KfB#eCfY;(bJ
(87L:&.Nf=Qe)T)<Te->XdL4OQP:OUK-V#+MZ6?XP4Pc^-<7f6^]@\=aJa7#^cf[
Pa-:+84aF+R/e1GNLSUL:UW);?ET,Z5cJX1HE/;FM#7#N_4F,8b#))5.P[D<+EfX
FJ\^d<S)Y<>I2:IA6N1KKfbCY5)T-^C6[/d?5=_+RBZ_3@^9CC(4&7c<@.Y>2Qge
8DZDe7c&Y+ZWf#I969MQa/b=S5Y4EK8)3S^#@L\@ZQ6HVX84MKeW>02[adMJN>gO
/9RO@Z8dOWXgbLaeLT8>P&,eOF)V(27I-DS.3TbP,&WEbS^#IPWQgX0IE+#,[M5[
2?<7=>16-eZTc/aSU][/.A<d2-2/H]OJeMHKZS;1cC1GZ2N^M2Ua?eS8==cDTe8S
QGS_DA]&d=XBB>aHegYPc,/FCZ,>MWLUbEG@c/>MY<bSS_:P<N3))7>8TC3C3=,=
R8SRL6fH5d=g9(W:Ag+(1WaKCf?HPXJ.bD8LV/b/?=CI=7JC;N()APVTd2a]DRZ.
7DY79XEKe\GP@SI?b4KRDB74)>BO)3WO[#J:=,:.5PEea65f;WFNHEHGb_LHLRL:
.ODUEafK=N4HTf0RXK^N=Cd[_]]&67W^c.,#4g69.MYEXGe\0d_)4\eb6aNRBTXa
H#?H0_efIDcB]_a9&:S@LX<b4[=dH4P#aR-S1B:b\:13VQ95X;4?gRYJ^;X:/M-D
35T/),)&7N=09CGZ<6bWR4+105ESCdb>c/YJ&GeLaZA+VHU6;7N[LE[QTQH2SY5]
FL[)@g[_>P9[GX<NMVHFU&VZAbDAM1QO+Y^<PKZ)fR,g5VY5[1IG;M2Q43bMdcb@
(+(<_e7;G+B3:,HO3>^3JBeEC0H^+;U?:Pa<0g_L-ADK))_(3(>F1g6C:2ZBAfP<
+Q.X4GgSSIMgN]bb?<[/cUN(YAb:cY954g(F/>1/K1ZZ+@D#LbKI]]OXG_-BA7S@
[8DR)2b90Z4e:J\RS:&45(GK9/?T3F&bb@[41(2VZDO2]fa)^X/-@gJTV[#]KS)K
H4@B3M+UI/g307KOYL?C<+41R0A\S?-#(SOG&]/d#a/Gba2;93PHBZZbG6g_.@EJ
\76Z9&\@aB5SeD)LaU^\I697/33@4ff/d8ONd,@0=OEN^FSBQ,3dZ7O0,/&/U]<D
>YAd3L:.P_VH-g5EVf5J6>aQ]@R5fKFeb-]+EX07-\5dePe6\?)XgTS>E[CS:(K<
B>@.0e2aM[Q<XdL<=?2SYeMYINBSZg1g8<:R9FX_QM1X:Z.G]@-4a5L@):=)Lb82
/Ge\e<5Vb,?P\:5UG?Sfg<=K4VWR8]G>8AP)8:(V?8X.3NNf/?(G,D9IBS(g]3A2
0WZ<baa;9>9eN00eG&]<.3N/AaefgQ8[0A679XWEZ=2g7(+gMa]16G)?&dCSK[1[
782c]T/\f>P(7XB2a;P67A0ZHgcPO_)+H.I[X7HJF7/O?0)-2:BU>Y@[D:T]gUeN
b,KYHSKK^..GHGH[.gPP5Y0G:JJQ9V0E5d[]?c1/>)^a;IW3P1aU->D[,4T38>3K
>YPTaNb3OGP6=ZHF+2+g(RCA3SRN=L;BL_;F[W^[2QMUE[OABUM+MN<gM5f/MK#L
;UU1egb+Efd)R/SbH/d(LAT-A;R[R&#-ad865Y-15d?SD]Vf18.N#29/YPBE1GBM
H&V_M_Q6C:ZIGddUU#c70JEY2(CfdU;F[QbP2KK<a-N.2^PA40X,QFJ0.MgD7?#e
;5HKQY9DU.4I\K6\],(B^c2V4CO5NQL8YP,C^g&/?I[R4agZS_UCIg:W^E:B4H=2
_V[JT0@-2@(=FKEDgXTa9TdCV17T52N^dX83S29S5EcRb]HEL98VTQBU1gK]3#KT
>^R,6?B6a^A:Y<L@9R:U]RDBd\I+>8/2@16SIF@YbFJc6=EZg0Y3cWK>C,gd/1\I
.F0_.=E^3bbUa5=bTeWBcOK^8IJ=U9QM;<N6UgW\Mb7fPXWA0D@451]a6cA52-AC
J_A)UEQN?E0I/=ZRIO5S2KT+R95g^HCWF:(5EL3eSF<aJ1OK>C,]ac&aPH[(d<9D
e5ML\++U@8BL4S5=0aI;CN1,U=22F@#87@;&<>c8Fd-X#9HKTR&1Y^U4Q,:@&:(0
)9#X>Q13U43OO6P6VV.&@6Z7K^RV(FE5GbP53e0U0FdT.[8KcHE8=7\3WNN4\?LJ
L#\/:Bd9bEdd0>cN<VZUBJR6HdHXe/_:6@+?,FZ-6[8UF+.:9.2g\f^,CdSg:U2-
^EX]M=#VN3@KJ:.7@L[_.M4>bc:=-LBT2\X)9dF@WL:96487f,]5Y#-MUXVV\,C+
1-W^@2):I0@Vc8S8+WD?EZ(\SRZegV>&1dX9.4c>[f@G#4TXK+<a@1LMK2&CAUTe
);YV6)4I74E[NRJ0#cNFP\F5e+GLU5Y9KZ,M8FgPI+A^38I,YUP99e_;IX;T+)-Z
bEQV\aDVWWC,@]##D4RX8Q]bL6,E\7_Qg6.(U[JMXb&a17F69b5D0SBb.9XZAUH0
0E^\_9MPX/IX)5^CKGGSYagLV)P;aOcU0:Jg7P,N,dKG1QP\AL^>S+Ha6:W/1KIe
/)53)[Y&/,.T]^YTC96K)P^-4R4)=>75MDa)>0aIX1IH3GQL<NIdRP<Tf@ZIYT2V
[d8DE(a<MCT>;^\7_GF&V=@OI[>6_ZgbF)I39I:cJ9a)0IV_NP/L09.Q#/OMT.bM
>;aGKTH8)4)U<RbHQS7I;V9+UPAEeU[NT&cCOSd>=,&3CY@0M;/+-<:3IYgW?-Ea
B:Z]1TJc@a?e_K-XG^&EI>WSa,+)U.29TC,8:CM6PR7SgJ\ERE0,CK?c+Yb?59Ra
R>0EgZY?D.8:.VDE#5I?-1dPcK3-K7,5;KcNR-M3Z6edPE^9QLQO4bK&a8&8aeC>
c9YEYT0M?;YG3M0XKD0dW\1L-A+LG>(?ONea>0I^:b()eJb3?a#[&EaTO/[If-WB
BIV.GCJ2RSdENJ7Ya5V0Y9L[@ca,aAJKR=C6X;O/gZgRIW^bD3H5C2^[P[SQJd1:
begYS7HNNXffcU+GQ4DP6=g3#9D<A?@31./dAVd6_KUAD_AY@Z\//MHgM/V5J56U
O)-=X0aZ3-8R7^3J>L6:-T20TNEOC^FT_gfEcJ[,W8f,e.ac(e-A[cQLS/3CSQ[J
D<@aS.bdM@:Z>.GRCFI8d>G<W2<,e4Fd[.)-Y\GP\\O3aGR&6HR5Z&:88g_TP2N>
dEA+Q[P=H80Jfa[3X9dW[#X\\D5QQSDP3C)0TUOTYQf_H^KVESGEZ8_O=?&KBG7<
J5-@GH()NA[94K#,d6?d6f5\.=,2DY;(62.G/aSBR)]\]I_Y#IG:a^OHI>W6PO6L
8/.\?PRMO?6gP\dA^9NR<H#,/FOMZ,GZMN&#9gC>cNGMWIU=-MSD6eE6BBc>c5bU
^JPJ6<QbRG3LU=GTA0eLNP^CQ_6G=<PFXI^OfZN?B_PP[bfcO\#<+F]XSNWdFHLC
=gA1=LAg6Z-7W(C-1dJR&SD0b[UZ4@7BOKFE7W:d,FNXQ,1R-MdP=^Q=U5-DaJ+#
T4cFHVQN7[Z1)JI?NbKf>5Rc2TV2.4JH1XeegW4(U:WAHYX&D)QXYG:b9CQ\,gSR
d+1dJ)Vf))ROA1L&Z\NV^&KKFH&Y/Z)f1GcgXZIB&ZGR+XHa;;LAA\/4ZYZ010MJ
<[V8,ZXLQ:12O;Y(V[PQ>G_\CINT9\/Y(_:3COBI68:-a8^10NM0EVBH-^9RH_\K
VKZR]+@:/9?9Yd#?,/N^Hc.9(S(/Wb5M@@IZ<>6]DZC1NIQ=@;Y[4AE=<M4)=QE3
Og&6A[Y<CG9/4-9:#Y4B34PQ3fQ=Q[)/&Z:dI=2WVOO7cQ;5),0Z4TdaKd,g?e<#
c^R>?,HYA.fX6Y(bLG>f<G@QH_;DKG5HdS/^?)S>S6b]\4&3J&EP43G8]@&4^#9-
A\gWOA9S#_d]P@4f(Jb7+g<=b[_)gaN4-<51RfDdC)PULP/Pe5,G2AXa]3O8F^EU
2b8K\aaB65?/HV9#8Jg#<HdFdK3=:,#A3eT=JUc?S/<H]^SEM_QVJ>E]_(QOT\NM
CdLbJeL0OcPJ\)OS]&[1/e8K?@dd4,F];@VT?=U]gY6[^F/TCCQTDT#]:R,-:U@M
DS&/eT_Y,N0[ZO(V>6Q>NXO9R96C&gJ_a>NZg)>I(#1=>GBVI/+SZE#U][>LXO?]
4g:B@?&9(,3:7.TNPGNOH7_=)I;>H<]J>F,9U?PC+O(VK.DWZ9cS+IEN5e4Q8PcQ
5@[4<)XdA7TH3>gLAIO2:>4c7/?/R\E5g<>XIbW,Pg(J1.3L_DOFF#DI-V?5#].<
\\N(58BgQBeZS_B21_(b51dTE+e[F;-Ce(X^3gF;@5/g-R(X4JN&(G6XJKU=WOPY
)e@3PJ]FIb5V+1?gOAUMb3Sg[gXC95,NN8f/8fA<3KWJW.R>7BA-HDVA0YIc59.>
AU84Q)QOb>#SM(\UJc.G+P?W<IN4_44;.:)PET>B7WdWOBES]:R8L7)@[W1ccB79
.RT/cY43Z#Q3;7-J(5=d=CNR6M5e&(ZR8cT(D;&FM>_\5(11LZN=N0[#eYRD6ZK]
7Me_YLMb?W-G6J#QWf;dH)HEDCCV)[HEVTgCPSY.ceL]74dU7ZGRW=AW1^Q:I,IB
,[[K<_+cg>5e^.WbBQd+KeOTC,BDZ>AZ:TGM<J=6\ff.K#3[5_:F:&9:d/QAeOQ5
U<Cb8^E,\16.bR(?g,-QLEb</...[R#bR:7[RV376E:V6L<b?>OQ?@T94\>Ta@#W
P^:)T.^Pg72=1O63e.>R2<[L^g([XXd3R\eLL6X(OcLUF[69WY[..&Dc,;.QS1eQ
.[?P6NG-3/SOTFa3Y2:8K82RM<&P[MH[Z-fZD:S.,VU(TD5_M3-eGG#]>gCUAea7
R/83;)R8OGI.bB+B,<K1<c[](5Y7CVbcU4_>(Ne^Q?\S9<2.AG7Q9c[5VeGJ];>8
ZU2UY?LJ[Y2e]E4<>Lc</EF<-ND)a@Z_.\2U#[Y?RgaXI(97XQ_5Y?b#>B]U6AA+
,f_^PWGU/^:HA7AF.0XdSX:D:^G:L9dPg8-8^&0:LHe8P]-25E)7XDgeg_MKbD_G
H]Kf/K\:)+B1.GTW.J[4KcdJa0gYA)WREcJ[?-(:a#PC(MF^V3?1<HReC85WE6N.
\H&U1g[PNBACPgbXaIU09WQVIc/e]#QC&V)#?Q?G[AC@CXU1T@7YJ_0K8.ceLJe:
XA<89dN]/0d?:BKZg\>&Cb2+R9^LcQ:W_V>6>0eb=b_]5c&HT@B1g7:RLW5)FY:@
E-2]68BgJ=CNO:NT[JH-U0gag??Cc=2aBQ,:M<&52W+M1S<1-E/B;g.AU?3b/&?X
3@?0>1aWZ]&)19GF5,0-&KCdBaH9+RQ>XOPPU[^g0_LG.KG:d0KJ#g.KS.=.[FI;
IRVZTV?1-Ta^Z(#=GY>HSebd+M\8bGUL^b@II,/9-OEQA8<8=6c5D\FLQ8D>BD4?
Yg?M-]#GEZ=G\^7Q=T[^W;QNcYCB8MDW9P_-F)a2b>5E8_96eBCe=8U<8M2NEQSd
Z6aVIVQ6;9d//UdU\4MK^@>2gJS2f9U=E9XW:M;SA-gMXBU@)(&gE(Y)X4DS>ORF
H>E>8O-LNgJI0_>JP1;YA^Qa\_WMT4\BWC:F(c\b&1T/NH+S>&;@70cOFa)_WN-d
R5-Y+Y:.B[55OIHPY8,-:g)OBRLCC40/Q\F&cX>[?R>(EPHP//Q,N?:E5NCG<+2Z
3<7_S3D_/5bfCb-8E1&T-e0_#>MWVB]9L4.;)9ZM9dgJ&#D)KO(&gK#6_bcea^bI
<@V.F\-H=HGUN)MX;_#FZ&<FZW-bAQdS-f_PTK9ba:a;W6>&@DONRL3PFHbGQD/Y
\VY:?NTEaVD&PX?&1OXgYYOeFBEW@L]0ID(W3U_.VHI[<LbX8()36+(O@QgSE.GE
KFU#\MT\,IN6QdTI?8]gO]TBgO.I[cEU>KLHK_b^<M9VS8eM+.^?.QB_aG0fY-0O
:Z&G8eURDN32I)RfB3RM(NWWI?8cYUZ[F_Se#_#;+WI^2(#=@]d+;8eQPCRHV>WX
Pd\F\-Ne[GLbG8^82[RCFAI>PD7:BN\++a4SX@B1-gZMXLA.TEKbG2:N(I_fK-H,
YKU^ID4QA4IZ=KM&_<+,VA]e67[/&83BQX0DAb=>[L2P-T3A2,/IWJb87:U8d?9/
4J;)-=DN\.FY;F@Qb,=aW3C9/[<U&+.3WaS;F:#X,HEb#<SN/)aC0HKVN<aH68Y>
0<PMb9D2gXcEJYeATYO(+1Y)+Z@9DK.[;a=^g9NDd8_3W]/EU#IJN+:aS4U3a:HA
#-W7?S]SFUE08@&bWR.]K8\#c((L6cFb1J606Wd.0a/O6[7@KS&#Z56QZ7._>[J(
6MF4Z^7<2RZ@]f;<>P\?,T]5N4d^eUb8dEFD)#Ia95PY\J2A?d7>5=Z#7M,83GE#
VaNfI4G8_JE8(E3W.J630#TAY^1>OS)_dEWEX]GPFUZLXeIC-VLH__,a^TBHE\2,
YaZ8,0=70cJX@V64_;?V>Fcb-[P4KBV@C[Hg_[T]B6#(38AG#WISYY,bCGGeK,Q/
GOE_g1M5V,;F9GSOJRZ=KDVgCO3HH\4<-QS;>8a=[c4XN&+7Q3H+&Oa?13WQL/O;
+,aN#/B9^8AWfa_8&+G9)Ie>C84_S_LK9TMVY58NV_ZFL<aZ=M1.>WLW6f>;CMX/
14a[&(H=4:@)V(Q(C]TRRL2;Z&,\-/aO0-T.L8,^aJ5O1CEdV]H?2#X]KQK;@:HY
fM0^QUN?dY@cJ<P(?@QZ^>CUCIZ@/YT>[>.See:?&0:_SZXYb+?VFb8QGd>aPF16
B7.dC_OcE:+80X:3?-W?_QX:1><TE]OKE(YH8:MQCKX@b4f1N1@GCBBKcC2C9J]c
YX;KeLVbGJ)&=3<8CUZQFHQUQW:+)/Z_?I,J8@YP0YG>K[.X/Y3\Of]]U9LY@Ya-
5A6ggBG^ZJKR+QVHEG[dXGCFFC?H4WCeKHE0WHeS3c?KO40d9V>d+Z=D+7XWdbWR
\6QGU?FB]@Z\R9b4MFBEPe/_:Rc@M@_42<H78a8>HU2IgHXA@.G.Lf=&@39-3/?.
GGRREDaXfL<QfPN\aU=5aU(ER.d=8KD1E8#[D.+./M>OZCD6>Z#;;#N?e65a^/#(
f,_f.JD^\g?R^O79/[DE-MT^K4[71=O-7MJd:Q)O_02S>D3OJ5.bBYf^)(PE\HCG
7P.?F<gg4gP,QbcG7d0F)ZZ^cdd)&MN4f9)1MV9bbfaQ9M=:aC8+=TE5V3?O\+:4
8[\Ia]EEAGH;?SJM4PeOBU3XCSXbcF7dK;fSS_d2,75,3K67F(K.WVDgd.U:g[[N
g)4dL;O\a&=#?(718A.#.feW7)DRU4-b22=3OG7.#+[Z^0O2cLY,SOAUN[XL;dWK
;cYZP#^E\\O&KQCLggV_:YPH.<bV&_fL8,G[4K1NJEWZ9D;58XYET/81cNI4FJ5;
D3ROgRa1A,P/C.9X2.QY.6a_7FT9Q9.&):7=WWgY7IX>;cBRAEE?\Rg<:UBL@SFU
X\W1UL1?1OD(F\=OWWJ&0,+UT[+GB+ARL2W=^+0F-ONS@\a?b;@cL]1=f(;I,7=9
6L2A4R^H24I1)f+WJ&LW5N&.N#VcQ4+Pc13PT8+2^7OA=CVg..T9W)ZDG3#YcG],
DM:V&MA#71;+@&1#cC7W=K).2F8(XD@@?=c_bK.WLG^8bV?&MNEUX;1B]L5/K>Mb
&^0+#>BEeW#gL><fdd_0cANZA&)6Jg[eg3V),^]>XBL]6@dNEM>X(^5X;TG/1N]9
CR7]gTV(<3d;c-TRN/94IB]g77&8N3NG43Q(MV9a:M>,Ig4c-e51e]TAMGe0:X=,
ad6]Ec/53+K-K7TT]bdeF5L_eB&:+eS>#NHLMKS_>EQL73PK(T2)>(#df7BOfBdW
2OL\\OeO00RgXTQ2Y#JUB8Q[V>8P1&Y?G;:&9O6O#+K>;d9?V[^AWAWZ3.M=c<QS
#[8Z<eFAJeg&33^_e<DP00(,a)S]YQM38S4?g:I#SV0O<Nc@1GW:R7dV]4\PK8f[
e=C_,>c<3<6[+].C-X[^G6Q>2d\D<Z(P1K?/]X-=#]3XcNQV:GZ&9O8S20-=US<T
HG<21N]DNR:E.(1GF7J/b77ZIK;GLM_6=#H/JSQ@2/1&ZQLB[fCC1M0=<>42HP=P
1b_>b-GeX;H[\4Uf-#_&QK4F95Rc5&/:(QIg;g^a0[>P+_/PUSA]T3833/[g_b=+
U<Q?&GVaOI73eUO#5N1A_H3/gO8GYQ.ETe,G@@WE13XD(QXFaP/[^.:gB6EOG]25
ISYF_XQK_[BPT4--Q2=HF(=.e(UB0J@PaN(XV?S43c3XK_-O@C#e2[@DK]P_D>K=
EW+XV8TL^cR&>3S@(]XdFce-[;bZ0U2#4&P6:3SXM-IIJYRKB=\1\g;>fdeDVS4F
97N1agH44ZE)&]S6[=ceW@V156]8VPY]IXZ&?=^2dJFc=IA=9W]b22#WF\E^\:1b
(TUgYD-D]-]VVJJ,,,a9Je]433cL;,90F20f?=TL<3L,HPHCK=]KEKK+N10@.[7_
FEK9dc[c2DD?7<[(5<D_aTSBN1G#X8&3Dc,HXI6Fd>JAbJ>:_Jf:_73L>#ZUa]8?
c0=P2=XIbWX9IC;aR8?g20-Y+\F:@bP)A7OG4AP.MV9U_)g@<>VGN94WDT-&>9RR
7G\ZcE[39\5H(]64H-/[dV12ZB^>KX)4>UCa^<_VH2)UF316J_+4U@O+#:-;(I4#
-+<GRJ^faX;JR#ZbRZG<;@gXN;1R;^aB209IYbN43^R2P>[4;)<BO0B3].HV_@.9
QQY#59Rd)Q6DON.&LHU88L4EO.1]Lg)?b&QZ=X#,F^)Q@.@c]K@O##&Y+Q6^c+\8
M)b8M&M89ZO<42]da4/EFf;MVI=_6E]TQAG-W6@06FL:fOVCcFOPObW,He#GR,aL
IJZQTfM]&F/N/XI1.3-Zc.4MH:T7G8@(S6.c9Xb7-.,69PcVEI=DE2BAIW8[cfE[
P]f;@&,DY&VAS:e.eC7^6-_Y5-+DEK\@UaW6(Gc;BKAf.IW49C^1cMNR1>[[KH[Q
V(<7gU,bD><RUC=T+K<d9O3Y/_Z;0,Mab#A4SbX\5T-<63.Tc@+OJI/B3TPbXQR@
Q]4f1Ke#Q-2e\4g]RS?_=&CT/feB3?E04=W_]^PLK@O,X[UI,\Z^<B]D]:BO5dR,
Z?E.^fHITVNP5U2///(+#UP&dJDGT1WJ=VQ1NZ\&6SSK).?,>F58JZ-AD0N>62VO
bO6=M_(bE15Z=N&;Z5_#?Hd>G>RF.2M227XNZ??8M#(0C_ZWH)/XJ4X^NDMUf/0:
+HI68&9V&I16.5KMbe5-U5RCJe(e@-#NT=RdWbcTZN37FPLV_SZ3&75#[c#Q@/;U
29OM;VOX(;DG_\1f7KCb6dV>\Y(H5;O_g_(MA;G:JPDC@L8Q3ccQgKeE;#=(VcJ8
C74WL+^Ug6Z,MTDV9=/I,Ne[-P[KXQ6_d5Lb:DG;RA@7#cJ@NHIO@)))Z[,3.21^
,7Da_9Eg)#EQ[[4UU6]^63M/Y=5>2)36H4fggdF=2DV5SG@U_S1[L][RZ?E,a52Z
Q0A,MNX]e4[aGU+@8A@dKW>SQObAb@[[5;bDNP(V1BBVC6A0#eDdZTR-IXM]M@CX
aYdX<IR[P8L4>7>(eT3-&,J]<_I#@<UK/GV)E;+=1];&\7A9<KaP,/1:2&[6>_.I
Z)CLaD[g\ZWY4fW,gF2>77YX-;FT7&\d2\U7P&XW97#:dZ2EPG?VN3ed\2c#I[@G
Y=JS6HfD&g.^?:F97Q^&Z;_6Y^P03E\b09YXR18F,O<5S,G4@,e6QfMP_XR(]@Y:
eOa39;-YGQfB^.3X8(<U<-IYNK\>&N+/MEEN7fJfEf@/6EL0>b(fZ]+UD3M>.,+=
X1XH0>^gb>AV1,Ia+9>E]71K(fO<NSP,IBOQ9f-SBfANa8Y0JLe&eAPXdMg:E8KT
)g]?g&_D>beI(XOPH]aW)gbOSX)@9)FSN?OKXUd<Kb2@\Nc^>ECC]9,D[R>EOA/f
@32,O,5+BbKVGCN/7D\PU@TN8W.]e?>_^243U1Ze\X24PeRW;;O<LCTMIA=P110O
fGcCbA([;1=9F.3DbdQC.EU\VIHSR/@7=-4[?ME>=^M)85L+JM<6M;FRaPT[8@]0
);BWabC5K^=F(]MKfTPdY>Te#EVCEP&A5\f[,(MdgXb;KQBT&=b4VV3ff.WHcc)=
CBBWJ8U8X+O(g7f9JCY8Le02<VVRYC<B[M,&PYQ;Vf^fR-]+EacaQOX^?<Te-c#5
:WS?c9W59K;.KK[T[[?S<#2cU\]d#2.5Va?L?K#VR64&eVZO,M?a.4fB4S8Pag]R
F\1V230dEO:^gWN]PE)1IG_0HGOS(G)U-3+QSZA2I=_U8T0PI:_2(2VFc]D4(X^V
?a57)CT>G(Q:g=(<(T^_Db8Y(Y^fAH5Vg^IQ]GM+LK\RF9?UG^f1B>aB_5Y7TNF^
=dd\;1fUMGH&=&DH).N^0Y.)G[)=a\1HS_#f@IEW0Vf+14OafNG3<6L#TP2_E=+G
TH4.<K);/@b3]<B>8BANVMFe7DV9_+_Lf3YdfF0=-_W&X28:\C/P^OaG-4R5P=I@
\-=e@c<7bY0&JSg?-d8+Q63G]3\-:JD_?B9?DV,QP)>]6^__C&\4:.E8bPLZ(,?:
DNE0#<4bd<EE=CJ;gL[b(dVJ:Gg.Vc9NX?3+?\&Z96];9dK551?SMPZ11R3L#Ke6
I,4d:VX\9\&a<QJ/VJ(_PF7D/-ZM<WWT>AXVg&@U/@98BM:22&cCAT7dLBa?>:V4
)6^,TJc?c+&f,]_4L3RVOBI>(\A=PGS/X\?Wf_=0@599\?Pb=P4d7G@Rfe7+)f\<
2QT<J1/;SZI?<b/g#5HX[2LeY.g.Z1_@F0<;<R?]>_=F[^[A8[2dM+Vg6,+f9=WY
EM8G(a.THI9M^?B-:<d:=>/;RL:IAPP2C6]fU0gcD+2/g@;2M4>3E+RSgWd?+Q0:
;:?EPVbUaF6NV^D5<=B<UA@L\ZJ6=f=UV8Lc676db&C:911D.817G(J;?KGN,J27
RWeYX2D/J-d.:=EGTZNGDg=2QIE7Q(4RODeY@3KC0\fB6>.cPf[CQg?>.Z8FH_93
TNBf/J4FKH<cP=f7Ra)-R5b88CM2-73^Y^E&.?91PZA:<6)/S^Y=]0,MR68KEE]O
bD2B(<[C[bJX#BDE;MUU3/1F6)QM58EfHJ2Y8f?c@C&B;\bC/2@d;UW&B2><?P8Q
3,#2I[O3UR-@Xg>B5KC\;]0F1I&d-=+=<SDee^I.S;+]D>@DT@PYW.]73B=P3XM@
-b@-49c4^\.Z5(V-eKY7^48f4V6IOb6A?T-3e.9;0YL6-T?);8OcQN]L-aM-N>Wg
gA;9f6KI?Na4WU)K8eK]dfK=-X(KPagEWR^2cdT_^XELd2,JA;QTFNQWFO]O>-YA
XeO^\EP[]@:A?W6X.-3\&UHG&YCed_8NcGS>a\(U+AKO?CENNH\A#7EEbg&09bBC
;MKEPT@-BH9WDXK[70OX^_Z1)KGEV-T]&cSb&,0U=VV(3M16>4::O/,Q9\[7J1N6
/.3;Pc;O<:S9(cOe1@=+JBM7[\[I]I>A.NN2&e->,4BAdIMLX]&#dKED:A-@cUcX
>@[+7BS#FNUUO87HA\=>aZSC\Tc#G@Y(CX8-(?a77,b;#;f_Xa^Y\2=X]]KA2DC-
]C?(A_5=8NcDe=^@\fEUWSR7cQ4>V,XSUK17HN6TEW1,Kd63O?c5/_:Jae(SHB1e
QO,WM9?<\>:3IZ)C:1_DN:3==]LHa6(7Y2OHeb6,7GRQ=O<QR]5H?f&N/c+@H@+S
7Je<,]7(X_cXD-A<=M/#M6GSR>_2+_@/];F&X&Mc]>;K/A?&WNQ_e=C1Z\;Q4Jf2
>+N[CT)\R4]6_7ZUf&QA=/O-HC.[,.Qc^\H0N-VVL<E:@2:A]VfH[DO^=\RXZTCF
E\K<]gBM&aS.@A&7\68JYBUK1Q^^HeQJ,M\E8#+f.MKX/MbGe8;#6KD+,Z+e5B(F
d:EJ4UW@4J\K?BWg0POW()LL_VBG,g;Gc9GS3:Xbb+P?^Z-.NAQ1IE[YQ&<^LOfI
\,aIP9g5L1K5?;,3eI]PCcSK?3(H-E8]3^3PJ.>OO#IUP@AZH#SI:NQd5BI:3C-\
4&,IP[>+_5RH)a3+b?(XX+IIYRZQ2c:L1g@+VO/SW/#?fHfF<1)C/@.+K8bg,@bC
&fa\LU?Z\F5fYIeU9M_L?_C53UdD;TQVCeLZGC+CS?=f32=M8[&G[bJGT8A6=b=#
46D>1#PB=(-(8=YTW&A=\X)JL(AG9bbI8^>cE:SZ1b08WN+=C^W^#ZT=3#P>#BN/
9Fg3HX^W_\d6\9@f?FSc[R)76Ke+A(f1+aBZD7F\)JWR\17W-QG5;QPC]F#)@bUC
=d7I@M:[M(_CS5;OZ9I-,QAaLCJB9eEOX:<]fWca=c1)5^bd=T#LXXd4?Yca034B
FXd-<W^Me9eADK<?UOJW[<WQc#aFGNX7WaLfc(#Jf5));3<Q[gR4GF6N#NNfN5?B
CPI]16TdAf4dER>JQe\e45O9bfMMR8g-Y/^8R716.@D&EbKS.ZBA:8@G[&aEC9c@
Y.C1(3\-EC6S8DCPUfVfB?]2A]WOZ\)WK_dNgfD#.TRN/X)6L>GXMceC;4S(Ke:P
,DS9H9ALHF-S&A559UU_ZS0P^H]8<W1\@f?RW_&dOg@MF&5+?42ZED3U@g[Pf.Rd
-3YX-/ZHb,4NN/Q8&W<.2e;YRXG\23B3)6R=MOSPWRe:WMK1?X])/)#94ZW-16T6
6gG@e:6d6W-X(+[>E;KG9>6/4cDJcgA8b(b;=(UJ;[cLWK5Ie3XT7KEW<]\M5;<2
?H07XFZ>)GWeH=4)OYDPT[BE[.37&I;gc6LWKXNdK@f.;_;6/+Y4c1eIOVWU5VF?
8FcJ9COec(4646IU\+LCY;/JN,]7=b?6+5:Fa,+GA8ceYac5I1Gc:BTW_<-B(5fT
<24F>-&@C9d:e0ZU>9/KHDYf,^8Z/cBTW:8]T^N,51fH(6#T#c(D#ALJe7\f1LM)
IFHdPbT=)UfF_JRMRLeC3^/+SSOgc-H\I<P/2W2M7e>^8D;:EJYX:_BQHC^,3]bb
Ke:@[M;1aB\9ZV;:9M&[E@WY[LOU_,5F5ML//IDI#(TC99;DPNaOC4O0Kgc\R,0A
V\0K2Zg9C+)G@0X0XT1OYKOZ(-<>f9)XS(O;G:ZDB1g)67&fCbPV>XT^G8db>aX3
@,G?#:>AZG#[ECBS]?&_^RK^7G>RYL6@;FVRRD3==:21La(OP3>4O(6GIA14f;G=
g9ZMV.T.b?@02J[OPJg?Ef_6.W9MSID<e5&UI3T^_\;=MR0U2Q]DJ;+7MPgFIX:U
[5C7T1-5:L<N>-@)c1BJ#LBUfbRF/Lf=Le^UR[2f3T\c;-YTHWT^C2Q(>QNQI9ZL
c7EbSYB&PfG/L(..\9C@B(X<XbP(6M&YF,9.BF#d48,S>b-3M_c,9-4RAO,@[9]4
X+9-c?]Q9[=:.+UHFAf9RMb40/5NVWR&ROK.Ld.&F3CBY)B.)-Z[WaJdc]<]08^_
^G;X4Sb>Wd?8.D9^4=Pf^,M\WGB4fHc3dQPJYZ_&dA^<0EHKaCOS7)+I]WHK0\=K
-5d2F?Z&Q.I#da6#9?dIH+-(\aIFVRFab=Na5c[?-]GMTF-Rc9Hf[>Y/_\)DWbVR
Q-Ye+GIYaV5.KCV@CD,_1g:K4(Z/?/[63&U@)aJ2b4UV],@eG\Y5NB@QB<Z\9;AT
IQB]:g)4QB6cUg^?Pf].-ZE,MX#O:K]4aDa[H>JZa]&b1M61L]-+O]Iee(UMRO\E
.I7^MDNW(Ca,_,PM19GB+bZ6OVUN95IbEE#:8.+C5B2]::a&EY99X-2VMV:/FZN#
6gaTE&<We3#Bc7:QCQ7:FeOI7+ecYBe\DM7@1V^RfTcaA.,QI32/Ugb>WHd3fDBD
1?J0):BH6AQGOe/;_#7<.(V)?]M7OfRGB#<>1E)-5a-PXF6c:TFEBQg\T_=:,&9H
0QFH#^.c7HC(-dV;FF&8_??+gP.ZZ\)\WM?]-L4UZ(dRI\1K>B91W=PK:R5]SF/]
)YGR]&(?MBSRKMOL.X8YB3a8Z=6\/VHEE9I/A36HM<D\>W<#P(2>XI4eOG.0?_KW
Ud2WWV>bZ]>?\Jba.?LJZ^g51)=;)_HbUXaM#JafZK_QT.Q=WTe4O,F7(8c4GU)N
=^&VJa1R9.gHN@I@2GN?M1RHGZ0K?PeDdQ#08g\#@-OLE#_R_^^AaGaZ4e-\V8#6
0@EfU21\dDdKY=8A9@8MbF[O1/GC-C#D74Q)f6J,-5-<LC=P>6=H=^4S>?<bNNTb
VG^E,)\1e6>M71^V+[D?O]C,Tf,a3#.2O2G>NN3.BB-,<OBWSOVVGV+.\4]MEHA-
C#6W4WEJ,4^EW2AI@<0<XBKH>^C)U(2Kb./;KT:&:/]ONKS7cI_#M-T1@B]UUGD4
CP>ILEM-eXJ=f?:gGG)2BIW&6bG2.b@5<YUF9P,=8J:DgO3RO]UGML>K5CeGQb95
4J)Pbd4YCSKYK[R)&QI.5RQB1TT2-Z)[+,DCAF>[(-];I<7a-gL?<+,0J.5IPG[<
JG.WMaEM,AYH:6.GId?3B6/6,UF,7BGFWf77B>a0^AB.J0#P7-1/Y<NPZ\12F1O\
#B&,c6=D&T3O]7bP,g-a&U+C59F;,3e]]O/DWTD8HC=@d-NXR+9G4XB4HEE&X\Z;
XH0QK0ZaU>fB4Z2)YK#8I=f);N1H<X:.,Ic;=24UJ,.>SLJ8fS&_]>Gc&:gST-5:
[)MO##DMQb3Ec^TE4\\MCO[Z2)/(H:dgLT+4,)CM1UZ8aA.U:)71)ae&I<ea-Q,.
N8^f=,XZ9EXVYb,TL98KGNF(cOPVCYZ_[HA;.aX)+aW_0FS\eJB8DgNBNFbTEG7b
MZa/<1@5<88fJ/0&?JQ&JRU8FE5BPaR9T<FASeHO\.B<J@<a&0I(C<;d/GL2#T5J
=SaU5,>X4dCbSXYUdA-BW4Q[OO@C+Y[SV_dYd)-4G3N6X>?+(&;OTeJQY0<LSU_a
@e:+0WR,RI+O<>b&V[(M^&X7LJX<TEa4)^d8bDL<BPN=H)a>[__@ZNIUc7#IA&9G
EO^[_.B>00_+FP.8M)D_TZcO</K[?9abaPCW?(=L3OPAPg0+K^G4D(/2,c.+f@6:
:?QO^9dR^H>e_LC,FP-C_6,a@-,RMM8?#VEY:NJP5)HW79KZIGP&>&=5B==AgK1>
-S+fY/7W8T@0<7XM0Z.3IMLJIbb<b:P]T<8<)Z6NJ2TT?0,P4B(3VKU0X6[^W4KX
Jg7OG6I^FKb#N.(3B2S1;FTNGfc&,W,D8M[N4CZ.>518N^&/N?g0/A(.,O#S9-0(
OF:#+[dQTbYY[E/Y=]b):LC/-1\BIZ0ROS\bZBa)YZY]T5X,\8N\,?+\[8D<gc>3
-aC;K_VR_:ID\JX1.=W\#-K;3I&6+A#3(MI=S[Ge.978\Gf5TN<C9g4c>I6K-N,d
,bX6N<1D>,BXBVVaO(4MOZe0AVe/?2SU?8P/D^N)@R3b3>e:c.B@-aVF6P4</021
d7g+D2>f?JZ<SPWHTPC>8HVd+R34+5IJVaaDK;,[BbR<bEPaUB-.-FFf];=7c@88
N24&0S34WGSPCHTaI#.&[34GA\a>FK2GF9:M?>fR=/S1@A1dN;ZL,gVeS.)QDA8S
cKf>3W18_0ff[&0:3#I+e5+-&91,()Y2)DNaac>80VA.>cPV\0H6+MQ#8bE78F)A
#CZ_N5HgARN\b0-O+a+ZPW[/(bNCNIE)7D>=<cF\RCbD?cRQc74g>^Qf;^]B2^:,
dG)H)AMWTIL4J:>DA?-US)=44PJ/-aSXXB\ZC5-@9@dR?3KI71,R6A/<7GPO<UXF
:P5-G[Z/>ZU5g:@LG8fHDgXYH,^-799[CXgJR+&BG#Z,#f[3b#2TMU9L(&\H4IFR
KfDMJ6Yc:a28_.GAFgUF_bMP7Gf(B4g5U:VQQS[)CPZb=PYL]VQ@S2V?K/@3SDC1
+g4SI^fKc9]AfFU5LZA9XND@+_\,:W,c-@I5S:L4L@JRFY\:[)gK#9D<M4.UKVRU
X_Z9CO91DJ8-FMJVK8d\c;\@:&0e53+>/c@TB8eQBWH8AB\ZRbOeN\P6/U_C)Q3f
[);bIS2V+?H^B/M:eKP#FFb+_LI;(GZJOS[GJ-5<@>^S<QA2=LQV2)^5LA2?b>BF
f-X@=]UBECJ[aH/8VIO\dYW9A>&;.P13]/6c[(7V;Y7dUe<+e]fHg2B:/cTQ?>#L
ae.aO3X63;)5VG2F6P/:;GL&^aE3f[SHNIR?;^)I&N6@/1;30)?FZ+&aXSSKCR7>
@/a4<&L\(;g5PReJ3(e?]Cb[[GG7-MOM3d4_G=1=:ZadFU-FZ<-@3Y>1QI>?MV\c
(eSSCXLP/_4&?&J,3P>f.1X-IVEDB,(S^Q,W0RSSf;V]MKL:GM+3#(cbJS#>/TA_
b[24H@@N^KOc+g@XV8g/PBSS&6[C6VdG4aSN648/UJ130U8[\6Q9SV0.S9?64)W\
Q?N4GNEKd-]RV,<3Q_E55\,+Qe)0/7GS<C76+(ZZ,d0(Jb_4f;4Wc7BVK>Q:X[T/
>P60;A(+]/(b^1+;Fc=<4SaE53KA;MMeQfXVcT;F/EP([KMO9_Pb(Za8eLG&e)VQ
dY^;EW_QU?>X&1]G-<G#JL9WE(a.dN0XW:9;g34F_G:\&P2PX1C9RU=(RY<&6f^F
PKb^2He+#JLdML;Gc#W<(5J[VW?[=Sg-<cRRL_dV@#9d6NN.2?/052R?A2g@^Z-U
C-KY=G+86PZ,Ec#=g4B5cg]2WCK?K@/b3O^+0>-A[EWeP?E3+2K:D<g:</fFR5K^
1:1SUV;<QfT8cT[8/M]Kc@F-cW6fFe9-R4X8Vf.a1V&8U,+VWTJ\f2.XTagTAW9,
9[(T?KO+QRKFRd(_I<9W4:2Xge<PfVfe;a^=+f#.3TdZYA7Z41)2R/Z?&afNBe-&
>]D(gJP]Yg&;A>Qc=?#C;^>&EEgCc#FVI8DX_Q1JGL+dMF\8;BcN+IQHO[31;C:.
NR-N9I8>,6D[15VN:Ig[K3&QZ]E&V214_/c)eb5(1+Mea;EZ1c5CECb;(,7XM04J
F)VAI87_T7M;aeY:]61&W>F46E=1JL4Q32JW,QYe=?2__;d#J@Me=g;?@4[?]f(H
ePLI/;<NG6(:d5#P>&TYS?\BM7eMZYe&Qd#KHVL(H\RN=+CF3R8X;HY_<OgE\.K)
d[W&.RP+(1:WUL7T-V>9Zb]e@c@d/ALI-I>c8]+GY)cDcJFFPC<GdT77YL+;N5<U
d_+RGGX?VTLS)+bS?=JB1JYZf0M?f&]?c(Q5/9QV]<HbA;U9()._B<dRSR/,[G_2
[FSOTc>N\QP\5R@U5&CdM,PK.ZR.):\;[6@cX)dVEIRJ2eaGZ6b7=K+<=B(MOE?4
G&^>OJ_?b58/X@L1c>g,gA_<9V]=dT[UePgJb<UVMISRZFFCTZ=LE=[ZM8Y1B>U#
,Dc/_NNdg/c_ZCEDZ;9SL&I#@N]g6S\CSXNIH6c067Z-K:3<KFeR<ECY]<&MDU//
f?8\;D?[2V[af,#IXYg_V@4#E;]G7EB.AR2&FWWYGGcFd^Z#N7KL<RHLMa\ABPV1
#fL0QD4_dEa7YEK>b:K/J[b;=_#62JL=61f\&>ce7:1.BANXXE<6EF?Q2<e8XDH]
2<WbbIMd.bY/#<(M;Q8D-J]2c#XF)g3Q,D<UCg5\QcfMR.c&BESdO9e#21-<\_2D
MbgbLF5(@R#b4Ja(#3N/VA4,KD97NQ4Y]4T6T,BSc?&Ga])cCb)@F^2[P-6U6X83
?b9MLT4I6S8PRIdSEfe7L9NQeF@E2]Wd0&5=#(NgQNAA#&8COG+C^X.<H483[Bc8
X?/6A8F35Ic8;ScPB\[T>;UW?H^f@eP4e-H\L8?H;32?T&e5XPg>6[6C<>O<D2M(
Pb)&WJ6RP]X;M(J>5K2AQMOC-RN03I=Y)d/HGSMF#QdKQ:/&381LBb;J[[3W6?K&
fW)Hb]4A>4\Z504FH<A52<N2#4<MTL&.Jg3;\aNCU,,4&>2\Wg]8Hg[_c=[HA6?O
A5CLc[K?IN7.bP=3#&[+f;IYeC?HgJZP16@dHPB8RHgcBQ?H1^S)YC8]P5R^2HX?
B=,e<KbA-7#O8@44cEJ:GBMEG[g9fZYG>G9KEQDI6::F.L=LXPQfgL6VGcPgW8YF
D6&+X49X_OAc9^6Kc?D>Add93[a4[Z7a]?K+]Z,<Jcc7e71.)58M]D&IRFH?KCL:
[\OYX9Ma[fH&[Ag),Ac@>.&IaZ=2I6+C?&C22+EKg_VV:(_FJLTeU;^[O^Z:\e.7
F/>VDES<1S3-^268T,T?#1JPX^[-/[Z]d?b6?3QI_O5AER(QQ8>\19N:fQ=Tb4JK
D=USge&T^WN<d]3BUdeL9/\4_UbREG^/:eY]0E].N.cdD#4a;L\F]1Z1?@KM_]17
9H7IEZ>NBYCOAEAEfP=(W:@_?-DN)SS9OESdG;X+1N&XK-5V<dA3cC.OCcV\_ZLg
7:L;6e(8Y47T8O^UGMN2),#[)((,_[0Y=C()WU2JPb(APMVCfPf(V4JHF6+a5O3H
BVQN[QL:S4MTHc?,32M+,e?K@<]f0E(+1BQ353\CHXXZ>>PP;d9O,1XG;Zc_,8.G
+\UCEV&>UCAUYYH:<W6E)-EX=+K[OH5OfOK_DXR8C\Y;YY79aIeXEIX5QR#)#H83
NA0@V);O_K:5VQ/,GN.ePN4&8X=#K9?H@BGXc@S,D=UV44<0H>R4P4NSd_=,aNGH
aZ1J6@I<@=<RCAQEJ&e(N;URSO^aRd>RbF=(/;+4f7>,O@eU\RTCW,M^050M3#Y4
1,.XW])eKO5Sd/7)WadBXbc/L#IU?AJHN(4I8#)gfEg-9gbU-=8d6,C\X8Dg9IIB
V,WQM<3]JDNbMNGM0SaY(@RIB1bOU-NH7YI_@H:UgV2b[T0UJ/J,/9=/D>XCXaT6
/H6bgN33T[=FQXKH(O/:77Ac__;[NY>.G@A[#-;--A^G4_BOb(RN7MI7&J6Y&Yf?
7?2O7d,0N,(0GLM;Q#)2[Ag6+X<JFDN>]eAPNWT?eGAB99Q+23-c<8(SP,TQCUbJ
,BF-1^ZeKdgaNg93.IFF:_9ca-H=(QJF\<N(]_4g_G8?,W/9&HbaH&fXb]>X+cR(
9\)TKMPS9IYM\K:gSD.W1XT#AJ?YD>UADc.2L9,c.6U\_abQ]bcO=UJH3^1F0U[&
PK#S=).@^#a5Q-9HHBXK:=3YSbZG4HZTgJPXL^f4[E&D)&:,#,7KA7eI.\NC>BFR
J;K3ZTF#MI\;+Gf)6b9GecP?La6S+bT5ANJAf1R=JHS[]R?3=>SQ^9@=1(GZL[V;
2:_dYN1\ULf=0QKM1XL/A&:76.Z4K,NWcT;]F/]_3cG:)KAZ<F+IBF0:)X_UVFAZ
B;YNR].b5>D8aIaBBV&dO/?ACZE^0SZ&\M,^CdA/IaT,TeEdW5KME?f4UB-AV;F3
Ua6...b=TY<Y=5/A8?H#E-gRCKM[gDZ&C><]/QJ:WJd&WA5\d-/)4;L-AAcD[Jf?
Mc#KV#RNU@W8gL5H:VC3I;F-XN@5K1Bf#T?G)[7J;83XFUU=JZ3V1))Yb#U0RMb@
F/2/F4\YS3Q2\K#;:/=8E73/O9L>O[<2RDD3c3_\.F;>YXJ4XaM9;5L8,XA.f\_I
JB-cZc,I5e##E39:H.XX),X(?_Mde4GDS_3JH\7d;(eCIH.9<C-<9;a^&&3^WPAA
=0R53XBXK)EEHDXf7+b;gQQ=B)(G#bH:@>93&WP-bAdLMgcZTaRUH4DP^CQJbB37
W,Z_K;Y<>T+B.e42e&8=,]G7B_c?PK0[++[=T+)8=6J,2;[(?<KZ=;a?9K;B]M8g
)+fb\WU=H,]YfET9HN<^IB(_-FD46+K>VR_F8SAR0?W=0e2@P[5WCNFga+CB7:27
eWPbc,5-B#BIa0d4\)[TR3]L>JU>WM?RTIRB1-Z,ES3;:R.N&S>a)D5380JUE]eG
OUB+Hd7KDF:INPRF#@d_,A289@0KO:V7AY-4aJU)EK=CHb,<0/H:,^#)X>#\[C8#
=La:Y0d_fC;V,^@bOO,H0?0F]5^&B^#8#?E0@SYM?DHODb_aYZRMGB\YU)5UGDX^
:WG)4&\cPO)YTXV]F+2G5;b609B+7920=#^gK@CF1Ccg5]CEU>[^6A61,Q3/D@WK
[LH1TL+@DbNGC-^2_3BR#H2.A7E^RVO5A7UWc:Y<61_HTC_O>)]B<MR))_5b16WC
8fbEgf7TM=[,NQd=g8#a(0,)1]B\O#OX_b]_D+JVJY-:2=?gQe6)1O)_>N\GdLNU
]\?(Ig+J5Q:^4H/@ZY.@X[#U14MN#89[KDQW^e;&[D,A;B.TY.]:Rb?7dOdME6PS
<RHN.V)V_5IMc)A@R6DX9S&R38NC.dER1T\>ZV3Sg<_FC[cCMbF1P.#Q@?5[c01X
.c2\RG?(1C.AS_fG#AEa/03WY)T5\KW?;B[5_PH+84gGFC,)8Db+]-=-AgUgaW5J
;?8O;/Wc2..0NfO=\)Z^RVT^Lc9EbMD#6B#5V-P<e=ZA0/(b>VK0>7DbS=6&OI4T
UA07]Y;E4/I2JXgYGZB\W+9PRc=.^9;b<?CKaEa(:PMDggC5cTPRW,GGCT/@1;A9
6)Df4:)<^X(D<D#F1.Gb&+/]fT(]g=3H.\HZP[a]O4Q^cFTWSL^&e]3.Ed,b/E:?
\eRROf94A\W1;dcZR:B9XR)X<[+JMad21><9CH::&>(E5\Rd.T/1R6eb;b8Y46>I
e#;T47:+B9@VP/bZ1^1&CC9E^OSOPg5+8#OTL<@OGU8,7G-;=G+>1g4^BB8GIN=G
_7#SI5C)THX8@S(0gLd,-LNSeBKN7+=.W3G(??-TcfEOZ<L[b^?)4?/;J])L]gSZ
d\260()5UU2S,GM3A&ddXTb-&08J[RDB:[G95a^V8J#55W>7)P3=;0&O//c5XV>&
C_^..T:T,=A?U(.VO9)I,N+HSA@)&KMe\EQ-a[3\f6/@SM:c5_R&EPcXV&\e6Q39
9?3b;F^HKB0FMGBERe79+/GRB2NP)N&2#6dMN4K0.0BBc_>OID(+(=Ze7BB9B:X^
DWH3(d465/8\>N/_d&A\ZFEgQ0e-=fBf4S&)5eJ4ADFYP]3&67CGbD11@gT7^aGc
@baU@7;_XV.PdCVRYZB#-??f=B&fGSeC7_J.<)J<_#eVV3>JQGIe^fP9bRH3PaK9
(fIdac[DCMJ2AJ/PX6Q9UQ7@+\YVCN:W[/^^^)Vb^PG,74e@ee>+TCK@Qe</U5-A
T/2W4.#LV1FGcdL/OcCS+L:[d)HV6bCJBJV:)KcgJ.Ja&+\I5dVWWcaSE(2@IXVK
ILG]<>GJ?@Bd&KKdB1OR/,93DF]L44Y+2^Td;bd9<C3fg[1+?ELfEFBcT,6W>&W9
;QGRT,BTYU/&dLA#-.beHE_U[[c&J)1B&YB\38][X;g^P^,?<b3ZX1RX1C\_Nfg&
XZ>5W]:53H1cJI8^#4(Ia.QGg)CMI\(@0&VcNZ:SP2/gJUd:28N3<:K+^]f/P@BA
FZ#YWT.4:[9I+E)1W_bG[IZJ[dVX;f(6&fR2:;AKB0;KM#PN>Y1+@2C;U.Ff+Gd=
\eReV;T[)#Reg+[^?[/E@1dKSg==5[_)Yb@<:XU\8g5NcM.^Y#?ACZFYM.Ze[8Y;
+HICJ2@=Ae(9f)b]].+8g<R@U:c9WBL?IL/9Q_+;fd\NTZP@8FL3=)b\O^H0C)=U
RBDGe<&a@Cd:]O1T:.44U(51NNU,6[6]\GK_]B=OU7^>E.D.;=dMe?5(OB)4[M.8
fB2EJgB>^Y&?_<1E@I(<LN&Oe,SLV?=W5#//)C-HU)7YR8^P>_LId-+TXcA(e[,X
d-3Q4/6[)GcYPaWV7147YDBZ&JbbFD9N;Pg?2:)U<bV[DF_:bfT4[H.]a@U.;g-3
XE\M&S8B@OF4J#-a/.OZ6YQGEIPc99>IA1;&:R9C];09.aaD56Y:;P:I5c]+SJ7O
LSHZ^\IH0[/cI9+?B4MJ=K?Z)Z2M2e7#X[08b:V/@MTeW33LfW]IO84fV9-.71QW
07E]-=R8\&VO3[a-ZY@?9E6Z_+_JK-+[g#e<[7J1C()MJC;Ec>[D]QBE2eG^KCIE
U^\gDMR4KG:=VWTdO_T-KB&4eF_e^[DeZ2+a<C_PWU_Re:BI+_^:@STOD?3[LOFe
?,G8,N40-:(@8?8H)&3^NYFb4;@#IVE&7=KDHIfM>,S]8D&17E+/+]1J2]1eQ(&=
C\0UFRMgD92R580,@dUf:JQP>e/>?16FH]C_TI9TX:7\,13[;ceL+)+-9K(08)ea
0W9bPY([/LO=7M]cbQ5fIK]BcX+188HGW+#<bTAK=T)MC)7LebJ0QJMa4QV(a.\R
TL\HLUBfKcI6)E4:H9Y=\@KC^?O/R8c4T2EW#AF_\B&DB_g.UQ)c\1:Vb-B,c6X)
>=NNK>NJB/,=X-7_7^694)QK4;>]WS6Q58#/f64Y9#[VcIO])+#>H@/5F9E-d-OX
2gNWY.EE7/bGH2dafN8dCcL38/eH&Hg3J<NLfQ+9VGX:L&M<F>,Taf,e:?96B\PK
-Z68_:GL0UGN)7>#8/47c]-[^DYCN+b70#,&&?WK^?YMc;c,S\#D4R,YVg9<K-Z^
]8Ef.COS6//g+GC1:/S+AbQ>RZ0.#OUc42&-ON+Y6V3\Yb-9CHIGEP(;LQ>P,P&F
1,7K?LM[-BZ-XC.7=W/C0TS,6<\\(I;]MK;ZDdW3M7d,[F,8YCF-c7TT&Wc@LJI0
(573]bA73[&7[ZR0_/A908<edfLTA[):&1cZT_;7cgMK^Y7668:39V1Vc;&K\)4f
LV,G-afNAKP/G7S9^OZ#;Rd;b_36[-,BVcDR\cA:LV:#4dSHID0a3YfZfG@;1(cH
dX;cS#/=@N=//6#ESY(MZJcVJQa2>0S:dN,+cZ2(DAbX^E^LST6JA&M;/e6&DPQ)
Jc2_P)2I=DS=R?6HGR#7]-K5M>27S2;X7H9S)g+#^9R#0+(NLQQ,=N.S;R[:fgB4
DFSN:A(3W=9Z#f0R-TM&Fd0af>U)).N^JT_JQSga-TQe6C>dg>8+[?H)Qf\A\?/V
0YYaP(7KY=&gQ_D6QdI&O4XaBRIQ+JPc)1N[1/?<^X;>K@WGKEffYZAf/EYU8=UC
E=4b5W23+\-PL=#6]ILR][Eea1Y9Mb[JV<S:6Z-18,-)Qg88O0XPA_(SWNaKT]I^
U^c@81Dc:40?_S9G4[Mc9#XZ\C;#.PZ[NJ0IIgE2-6Xc5-<Z&Z2_17=>NC5Y,HWZ
:.W7dF5WM+\fJ]f?I3[e]2a5Q[0XFdLON6]Zfge(QNA2+DbgGg4=-L;f-B+TJ-aF
HRMDX_b1I+0/R_/WSVEEe[1^e:^.8.I0]CHQW5/O1B:6>J:XYA+I2P[U?C?]eVB&
)e3FX\MD&:CO-;_9GBW4&9)OY>71:c8?/I3NUVZ0ae8>M0SMKgM(eL)G_KOg&\B0
_aa)<VEcG-eX7;+933QMD;9H+49810]R=cG8K,N9e=;a+>F1fB18?VOcT#1NV+a=
+@Db3(VFJIb+0JLIU485P#P9)1bdF;2d4Z/A,NaW\;Z=-(<<Q9D^E0\4a/ZIE]G7
E]F]f9&_6T54EEf)VQ5-M6Zc?Kge&;3YG]_@;TNce0=]F1FMW-[_[85E#PPW1#OJ
+d/V#>2H83K,7GUP3[g37VN>/8)OBf@ASI,H&#[JRZ^F[Z&&&<Y^()#bKdSD^3QY
F3ZK03B2VL020](,P=Bg\Z>fJ50DFE0XUJF6e?[E+UKQSBYJS><a<\/_,O./f@,c
<M_W#D9?0@b=.S:0M.9<f^;<PU8Q#C+f>fI7D0+-7QgOR#V+aOQEVIaOSQMN&bP?
-bDQ2+VR>NZ]X,XbO3YU2d;3E[f:];HV7g0V@QO]+(3,Y((O7<MHB:\<HQH.>I+>
dRM5bK=0;)_O=(cA/CH^:UL:I7(F-LNa2LVe1<d.D:/2I=fMG1:F=JcZ5e:F4L4d
cDO\S31d<6GE>e\?3N+8;CJ#MSKL+]707ZBdE>L_8eIU2X\Tc7aUDV_@Bc1>\O>.
^JFF3MWLDVM,?RLHS1bD-8c)S2JHe<.15AgXPRfL+72R]K_376X4T,INfgEd>X-I
RFA5/\X_d.P].QR[Ba7:7::fMLf93TZ+\d^\0HS(=Dc_DG\&J/6VKTWg@b5M6S>8
K&MUP#AWg3;0<6VNPEFC4>dS\[&W9VZ^fgG2608FX9^+]-2R_CKRcg4U^=5/KWW&
5BT#RYD0aE^dTa?264W/&LG5[(D#>TH8R^/YNbV3=>-S8PdfMN,I18GH\@fea_;#
E.PU+>.+#POAcLJ<(#Y#G#\\XF8DYX0((5aHT0&FD6M&9\L3AE/Xc-Tb?;J^,7Hg
3T650326FcbI<.@aeT@ZVC9Q^IU6/b69GgQUQ9&Fc=W#^R6U^g7eO8T:dYN.+1FQ
AU7@K9#HX(Y4_Z=B6c=7Z;e(SVb\>=_b[CS>(D,6dEcX7R&6:&32[c->J<W;&4_U
Y2bF0;;DcF3E12FN8I>>9[fJOAcTPScOE&&D0;EKO#;Y&\4BOD:=V\&84Xb/P875
U)QTfX2BF7K;Af8M)K.dG0;2APW^ZdCE0XB42D@>V.XE5Dd>2O[W@^68:,9Ea1+6
/&9)5VIG0EF[598Z(JW58B(1X_R5a.g&>H?Nd2I2J8FTR[GI)3#HT1KL<c^e@=OQ
&UWaJWCJNN8bD5CQW>\I(W?a315](_C,R6[N+<bRTLE[2+\0,0D4.,R]HO59<YET
e1O:e9V@J&T3Zb?Y#A/L+T:6f;)X@8M)I]Y,T&gEJ(?9UVX;fOa2D8894J8LWA_g
D9f#f]4PHRQES80d]\##b#^[&V-PURP[^=&VeY86_:XdV)e._dY7DA7+A\dK.]V&
#c94O626gRSURH@T:0.I1+6+fW[4@MV@8@<4C6],42FR,A+PO\].^)C.1=9>ag1:
e3>J:A<+QCSU3EdCQRMX#3b6^B=R@N74JdJ66B.C;(<3bHN0W2O4=0\6,=;aZ/JY
,1a/c\_+(BPdZ142D,MOe]3(4-XZ^?a]Y-W/HOMQLP64c;Q/CW_aIg^Y#fd9b)PL
6H#Pac2R@5b4+,^d4;VeFFUA6DPf6Dd5[H+ZD[0\J)\,(7/3RO.XS2Q+)V17):#(
#UUR0)K(AaO=5dNJ??1<MU&;Y+\S(7&E_=@L#4NCFG=9>.<KO97N#ID9Q\0CfC^Z
F9_<Y^bgVX&3]dS3&:S@478B[0[#UY(RKG,fWZ1]ER(_DWcK1a_UVSGE<J:.Nb5K
L_Vd<IgSAJ77B\T#GV;EF1e-Q?(c@FT=#98#PRNdL]Ve/?YG7I\:A#N7>1TGUHR(
0XHa;X),V2/NA\6-g2,^6X5^S<f3#R&f_;5@4RHB4cdN/Fe/U\VOEELN+UUd>P:1
e<Kf>NJ^GYPECP#+DLN#cb02K)#FI.2W(5E]^g)5DZ_3^37ee&,3TJ&_gI1?HB&B
)e:FN=9gJP<eV+/ggM-RbPDM\YI6(7J9O_]@P]:3fQCLMcWR>?^1Ya.=W8-+g9[[
T;B0fZbAYO38MNHQDAWDQKW?/2F6DM;/EF&PE,b3R1@,7X8a2X@e/7P8?TXdII+@
)VRS;I3^fS2L/&EcD;f0@JK?.R;XR1e:SKE9053D]K6[3[]<OJS;71F\fY6E:#F<
)H>0(+/&47)6Y(@X<A:ZVONaK=]<0<]D=6JPMA5Y4G(-8ZRa]VL3/BgbM>1-g/2e
IIRUe+KH7BdVO)eaN7X]gI<&cXOMee:L.eS^C.@1fKG[F:;YX[NM/e9R;,;-JN0(
O]?#8T6]UZPEG_f;1-.FVIDHOb,H,SB6#:e9GT19ZD_HJT]LcYbQ\BSVHIAA&(aY
HWFEAY,\]?O>bOFa(d@-AU^c94_6HP7XFE9&U8c+RN4bK6](PMbgA@_#.<._3fWF
]VJ/8ge\I+([HOB?fW)]S[NOZd^EAQ#5@K8.Q;G;&AUg4,Kb+5P9&9Ee^JeOMGWe
.OC5YZU_E9MLRRYI)Y2VDMEdJ1SSEN=N:S<W:_OQG#/<V^ab3Ibb1gCfeY?@=b.:
6;b55[8[_;_4GG6F&AL3@KccJYS^g<DETR,R(g\@/02.a;UIX#^<9)c,ML,S^/X(
3J[N[M.U3)D\MCA<dA2RD./cGHS[GMLBTO2OF6cT@.5+X3Z?H#3fb\]5338N7_7V
L?->W=EKGeLF@TRZ:fa9RUAN;(Z<b?aU#3QGY1UFWA67L?c&:ST]8<AI_fD?,9-e
0#6/NbD2e@8W>[;YDX;OaXff]/#[RCM:13,X71e2555aJGG-<YIaNLSO4#[)+&G@
4WFD9S\fERAP[5T;>\5R_:C6CN#=+N\WNBdB7gbZ5R<()e9(^HT0M:\=f]cA71LM
Nc9.9>U1D@T4&--K2:RQ/MK0Y-e7UIG)K;.G?[McS:?5UQ<dGAbb[M6;Q8Pc0RG1
S_XHI+\F3=fC+;eBaN)=+)E-f?X]ATT<=_3:,J>>\2IZAGAQIJ/7#Aa9g?>^bNQA
(Z]A;=fTWR&af.?C,U<)B+;RLfB0IC4XPYL:0PB(/;)Pe2QQ=gD=L[#HNcE,KWZ@
A7BA\F.&b]eGO0gZISWJHH5E^)C4.(211P7+^G=4NdOX>+A[.EccIZXaN)^JG_5(
RN9-SEYVaGL4PIPSFbA7GW]e7#Da^aHG4T.RQPUa@<^>0>I5C[4\LDB5H;)6E/c)
@dC(7TTX^b9S@f-B\&X0H15Ic(Z6EBU.3/bb1MDLWSNXH?3X+V^15@e]B1.:HZC;
]Me5\-bS:EIDYH[[<1(,fR4eDJ9(3R_#D.&b+=(;M0gSK0(41Aa(OYUT1WW#S+?S
4C_J2SAgVED\c9LLG/,RdMTI1;)]QI_SZYDb<#EIM)&P-3I(b6V,9R-<b]_+/ML1
=5M[4X&IbF2P:77=#&:XVT/S<.^4;LAbTU9(Kg(_1]f5_Zg1=:J=L3ea;IXd&<1H
SPTBZ5g/Y=4WcfTQBYQ8>fL;VN]KbTfA2Vcg<acd,a[R;&.4X7AC>f8,-Y8^D?HZ
==?NWS\O@-?:?_&2(3dN@9:H;B+a/^10N2@fNgd^@F-CYT?Ie#dIHOTSFc9cKA)2
=<-/N1gIF^3BCO:ZW+R;M+-X[[:@[_C3PU0a=@ag]2YZ9UgSH/e&O55C[0g-f7;6
K>NQ^e>7-_H)9D?+2a@+(/R\?-I]<X9SZ0SQ#eNeP2[X<;?7E#2WT5_/]VbYE?D,
_Y4SKfF[Yg0SeZ\UC-;2+9KGG=+R9-e0\PaUZT;7YD-L#HFOI+I:?Id#UQL4cVB-
[(H@e4TS1<?)OV7)2XF0;L?C.Mg3T+B[eI/IU?=CJ@XWg;T)9[BLaLUeF?,F8R.\
L=FX&FOfT\F+5Bc>1]RFJO#9e3.\8?^NCG5Lf]6<37&CEQZb=/1aW@M,LAO_2A/X
V?=f+,W<)RP&]&#>YT,Q6,-1f3d=6SI^PLDQYOMdJ1ZbGD_>V#A=c\[_U\#@GPRK
]W.Xg=gDD;KLX7^\-&_d7QY9/F3g?W8&f.B/2@18IQ&MNH_8ZO)@\c8+U8?aWQG.
RU>>;:ZP>Z5W34-@XHR@1^1T_Yb7I^(FL.S(CX>gRC:QMPd,&OfYR]UB9f&_>e::
B8X#e[,;4VcbCVaBEEHVU>eeL#g)>,KKP6f:JgM2N&.1G65Hf(?Ea(I@N)R<B#dJ
F7R+S;&(FO#I_>M<67SDUY5&Se+O>RS_E9?J+?9UT0Q/[YT6eLIC&TA@RK<b-<3O
^0.fVg,^/VDY@9D3GaY[TL]07e@^R_Z_;VP3-#@DWJY@GL+c,N,c,>Q:#We[c\8I
K83>KBY6^;21ZT&[WI4.(Q6]8FRaL1eGROcK7F3.<-Q_P;;=bM-H5\dZ\e/-f>W;
7&c)\e7YV#bVH@+[PUff#g-OQDM+=3Wa7V>J-3:9JdeNHB.GZJ#:W?EPM+=<?g0g
6BQ4=H0(GAQM;2#E^XR;^(LI]5?H_1WgEWT_S6-;U^c33=MEIGW>.,[A21_G&=^H
eJZS&,F88OCVTZHP>GX&g3f;PdD:X[cAK[>F8VCQ@cUDQ.C[V)8<U1Z@M][aX7Q(
64)&3cF@:KfaN8)_]#-BL/?>_9#2-(ZTU9O^&[SKRMaR[87?g2[VU7HZZU#WWSH@
.C9K8GZb>Z7L23^JS,:#BA>Ie^TUXM7@)SDP^KV:2PJT\1_1EGe9QH5-]f<cQY>;
g,7+9MX=+NCKIfcK)eEA5KI]F4,5>:D^M=DO0<&K66e(4^J4AU9F..-_[GT#E\GM
0>3QKS>/TJ2RM3Y<fU^Q#7-#)+WfL4WE^D:.>KcOAAEf@AgQb?,.9[8HJ?13<Q6g
[51K>8M[9U\Q@B>V#7&^PNG=55[[XT2AbNUL.eP=UH3Ge<.&dE5e,I#X@VD:K<b>
fZc5:GHVZBX#b<(;S8dUFd=6<,#TDM/ATB@,-/.?E,+I1<c##de;Td<U[V/,TfXJ
?cD/QK^RVHQ-1ONb9WNVCZK]LL8-B)QUaUFV1?LcKOc10f+dYeHQ/OG/(T+EBaP>
&[R7EZM,@a(JaeF-06=a.#a:#JMLZ#A&GT/T.(ZO93AX)RYIH\#fPH-_GZV2_aM7
e<VUR\+L;X1CMX2>Q2T/\Y?0U=?85+;RY71@e8cOA274Qd+_CG&2d#&N<J#11g5e
3L(]3d/\L?J7O\#VJ3T7H4KggDgK4LRES=Gf9;FKQOJ+aIS2RV?@8-Zbdf,0fR1W
-[).;T:ZPB2gZ04?P07EE+cK?,:U09ae9PSI&-R14EFBIC8H\&aZf@ULCHe3KPS;
5d2EgH->ZW&.N>>c5G0AG:Ge9W#KC3J5<?Jec^COSS@2EKg)ZTDbB(CK3:da[FNX
2@SIc__,WJ+&J2RcFfR)dZ9,>X1Z&.eFRE]D)feg8ZM&TdFd<N=6aK1CIQ[Z_?>K
UPD3;:<NJH6-<9##?TO&IQ2=V+V)\g9(3\C;Fe]MLg&Bd<IZ3cG8(Q:4F(^gfC1#
-.65<&930:@@9D)16UMOa@V8e36H[0b&9R>P+,?SOdJ.Z2aX847IN.e;.^@FD_B@
&cW=^8<-JT0JH4X<.&?eCS\IZG^1\<5.5#=--d-IH;>gQR;QYU0(#JfHaIe]f&_\
?,@785TcHVHR^PYN+KHR?0dYAT80N,VJCD=^/</A^/66c<.L8\-ZC__>b=F=Y\SN
V0,J^+10g1bR/:#R2,+>a.D\0F/NYL+U7MZMDCeQ^JN(P(K@]?+_ZL[=)DcRSHD<
a1O]@#7E716@5=HR[,,2B]WgDc(K0V(0BXQQCZRAF.<D==.CTQ8?F5adF)V/A,Wc
>)H-ASR08BAAAB-7^2R6>8W:_1<abD;2Yg(#^<_;Dg_Q=]&fI0c#;@d#]4e8:d1f
H^<MP92=.PBDC4(.a5e.9?3^Y59^UG5W]eRBBN2OK9aVX)@ZA_fbd[,@+;9C(K<e
?aKF6:/03)f5RT^C>cB;E/#T0]^C#ORDR>R3:W6S3L[20_A-P@aNZ<<8[X;GM]7U
&DN/A0W1.-)f\^O)\2Y4/:4e:a9,4=TMB[R(K_32P8@eWBYAb4Z.Y8UMY;9VSeOL
b^GU.53ZKA.cWT).,H]\5/QVAggc(&Vg]eLH2gIF-,P-b@/Y\>2&=K9=3_d=@>@9
G8IcTeUVIZWU,;>\YT:7]3\AI_RDc=?L:d-S9>81>f0T2G;-T[;ZIb9\),F0Ha]0
+32QPVP?@6NFK\=3R)bK5N4aV+F-:8@<LKW2J^^><E=5A7Kfe\QY,]<;ScKdgOg8
>F,0CY)cM.Sbf:ER&D09@;eO)UT[A@c^.WOdGB,2#:-CJ2e]FdATHB]O(WG=PY;_
9(?);8BCdAWfX@F3)M)CL=XQ#3=BF6TG#8KaM4gdUVEP,XE^;0)P]?98))CFg?(S
UbUd1#;(8Ye\U;BR;SI2-8#NP4K.9<5GRGT:WW\@J=.d:5g8B?@AF5.Q7A1T;dL5
<Ygf1E15B0FJg>B=#Z;277]TJ82Rd+8130QQC/g.9=C[O3-W=,[Z:#+WZU,-VdF@
b_Cf6(V;U/V5JV1?YP2c,K:E.85\J^:V,6)6f4L0Y/>A,S_=RCTQ>TDb&CACKYSR
UafJ1TS8B;ff@:>&2^+(B8DRAHBc+Y<J)9H4-7WMfJ:-^PJDAV(@(N8TYMBW2K:c
>L?>BMgW<[.abSFe^JgA3E#;@N=J^4c5(>cbEBQF)F&4?4S[JB.;SVE^KW<CM<:@
e+#@_AgS(VVTB&V:^[b1Of.==gEUYBA4c(BXN1S<_-Q=[GO]S?5W_\;[M:UM]RV+
@6Q,10@(UZa4/O)(dYK#]C<_\Yb&GD:W:Bc#a]KT27S=Neb6@d0;Z?e_eJ4C:P>?
LV#_;;A0b+a\@&-M6g8TF;(YZ:,_eGK08[eTV47Q;(680YbMB4_>BHUUU_S[V&=9
OJY4+CCHKdMH,+DIb>JL,WT/;GUe-7CSafN(bT0[IIP5b>M]+(S.Eec\d-\bga8f
0>XZ>L&90UWDL0FBRBD4@S,:9AP,LV.e_?5dbRc6>2=2\I6T95b2XU<E6RTQa/aU
;KB3/I9b6^8YD&#2L:IR3TF1F)/Mf6Q63U]b5NA,C;.M&N&4O\6^87FU^-VD2(M(
e>5C]KO&Q1YbW5DVC^WC\#49a6P3Bc97>IR/.Q2CPH_;-8,@\2)()I1&>\^f@d-P
/HNM\2&7<Zaa7eg30A[OG[&XMPbQ&RS_=N-^&-WG.=;eDK=D#-7c2+#K7D:V[Y]Y
0c[HbOH9C:B?Q9#G6c#1DBEaX]_T9W(6VgA\Q3#U+_IJc0HR1=YKDJ5AfV\+a#]3
X,Y1?\\JfMLB:-KQ(5FP9f)EXS)L1>652T/a,S1A4QMRTF0e3TKKS1[S0K++aeA<
(R21);O#H\+D82W:Z4?1DY<b-8=1(&RZNEB^Zd@H28A)P&3cF-F\a:U\cGeN2ge-
V/O&dH_BVb=a/_9;[Z:)dE66@ObSa=<Y[]K@?1^U0A3Ue0SHa<:/HIY7)#=>G@c+
OH332)VU\\d)557a#UeI4&0A?b:Nb@0Sb/(dIJX/MR>B?E:3(5a@d.KG8ScK0WdL
)X/]@H?9_I,ABGA#<=U:=f;SM5MAfZ6-D-:XIU98<^?[06?8<10cV?G#M3L7-b+O
4Zab8V4EAAACWV\,-1B;f5I6/ONT#3[Qf,0+U3:g5ZA&98?[fW#de9LT37^aM;gL
+_MUY+[72Y>V&L:SR9?@V1;:3@eMfce(;-RQQQ;P\4RLQgUeg3@:&0BE8N5Y.KLK
a6YF1VI7/\U9T?_#F@=b#4[4XZ337\8=G.RBI,Q(Rac+CNP[3Md)G_PeaWU<YY-+
Z;2/=EGeZJU[A]KY9H]I.CWMI0-Y1Q_WG1Xg7ea_[(;.]B6QB1f1W_R::_c6RVD?
O/a&;_E3Uea4]V,A((Gde-6M)g.R.C8=bD@=,dLU8L_BRC>Z039QLJAU[O^S(Q3)
]-TYI>9\TQZTZ(aAUM4V[6>DD/:BPA-S[cD41B^AP>;b\eUDY45?SZR6OI3F8,YZ
<fC,EQdNKF]GH6d8Sa8^(\,6^R8TSfP+Jd.b>VA>RP5[G?MCX=XdDJYV1QKg&IgF
JKKc^bXT1VJHZIeEedDB^ZB:cN6N00IIZYYaBD-M^aI5V)KWAW01a2R@[1T5)1Z5
KYY\,<CY9=T])@T5KbfWBC6bJ_FV1I\0BOR?cOX4#JMdeWHLeYHW->H7GNbM&Pe/
O/<-4_c4:?MSW5?d->.Y95B@F=ED3YRC/)FWf1d6Y\WM/(O=G<MM1_H9)W@80UdV
.b-gYC^bELX&(_e8Ea7G9>^4XXWgT>9KB1]X1NZMY49cQDa\=7_YdPbeLdPA9VIR
,KLX(Q]>#<OE]M=_PU,B4W89&<<gCY>80_\D5C.1N<L04E[d#U=YIFPVY:bR:P5&
<+6R9^H?3DVTS_ea1IO]61KA22TJc[SF1X><C7.XGPId9OIU58^VZ,eDAW_L#F>>
3d8N]cW@?BW9IL]R-9G>W(J=-/AP=gbOA(WTb/_QT(Nc-4N(<bQTa+&7A4bL</E(
7=c-T4P;KB^G7>W:Z&#M6/^HdRU:=+>#=:TfdL]b:J7P^IO9]6HaV\]Ze\SNSdgd
P.0K2@-(6JKD;c^VYAg1g&4\=+\25CX\B3a\IR3O[Y3W@MMPU6,g+[J_,^SO1;gZ
9W+=4MGOKIFI039eD:T(d_-13C/Pd_ZH:eX@D3\,;.[g4I6+95e)b)/Be=Q^1]/c
HF_f._E8,RTM+7\K</GJL[(bO3NIH#5/Z&S-[V1:I]d+W--Pg<<AaFK^>OcY0017
KHMZ7,bZZ49D^g-?^3PRXN91+gg\Z36KeSaW2B.VS^?#Z7+#5]K9<C\_PF-12.^N
\H[[+#]fD8]SFB<7,7DZNag&1\TBNB//.,@&)5@(MA.\<]S2;8QFKZSN16S7#SX:
e;1J<BP)PY(eG#H>4N0;38OSH\44e>G)OSAAID@^^SN@aK7Fa3@+5M)V2fH.e7W;
?EbcQa>dAIVHP1V+/QQF]8[64><-[M/2E)Wd?)F?<=]TJ:Y&;E.?>3A>J0@#8&cT
fK1f[KQU5ce6HWLREMRL+G#fMPbaa16XZ@gQeE:6D,EW&+V(=&HR(a-ZEO32[ZEc
6@g?0L>9/Z=8=LaQBFX=6[BeEC)VKVZ.(P,0WVcM8b:UL@;b5@^B:>W&\Wf3Z,R9
Y[BPFGRNF5R2@;ffK^ReYDKa1JA0c&\F#W;0Q8XJ5T3a:-RCFX:A(:9ZZ7V]=Fca
__Z_Y,&9VFa7,_eSJJ6NgfV3Y]YbAN8\H?V62#Yg40>ZcLeUfYGE6aDb-=>>+Y[(
b7H&D[-1#?=cF>6\5G\7O5cSN=K]NS+E>?8]_):QP8#cGHJTUa96BB=[+&daH_J#
6N@=1Jc9J)U[[ZeC?QA:83H_,./\+^P-AB/=])4da:[dU_#OQ29)WIOCHU67/.S4
SS6Q#eBFDgS]UD]UeeZ4GA336cES@+BRbPHV6cWa(c^eNB6BNd,9(G9C];(PGgJP
:@LWT0B6L/I@Q:BW7d04]^XXJe\MRD7?SgS;f,.>(GP&1dTeZ13/45SSG.:6F)c_
Jb,.6@2P_2U[3Z,M+UZ+^FRQgRO(.&8OQ+G(S(NL-,ZZgR3MPWI.G()4IV@I<>0V
P]#_VSL<[8Mgd2R5>d@6U)?[WM#ac6@#Ne3-]7SFCG1I\1H)BQ]c?<EVQ&_dUO3d
aZ9O/gUb3JgJ5M0NY+VS@@C,/.WDNNU02P+&9Y4,?.CEZ@[<TD5Mg[7F7-[TY3bK
0D+IH1UATFQ?feABIQNDL=dJO8G2?\Q(C=8GT]EB^f&TeJ00O+3ZF#A39a/SL=-U
&^f2f;MaY#IB_#@S]4(3X:30=D+(SH[fI.c#bfC^DV<b2]cM^Gc^aF5<bf6MfBXW
Q0DN9^d<AbTe8QF-?/F=5)e[e6_TU;fS,;[LFeR&SVdDEYM2O&T-&Lc/+^]B]E]Y
AHFOe-1?J]6Xc5cD66)HaA..3?T\LWY-0W0GVG7IfgU27B;5#cAfF&JE,Z7/M7G8
X/F.^IPVA=dSCGVHZ>[f3YWRXFPgN^0VK1JX-DfcI26M8D]&a7:(2PMg)f^IMJPS
aUCg(5OMdACFYAUWU\+..LFJ;,e3a(\&+>E-7_fKZK(@\R)^W[VY94e&/2/3TOMO
Bd^Z(V3+@]KfZ]>C.VL?LKP1KY33W=PZKaD)1[HP)V.AOKa5Y\(U88Zb&@W&Kgg3
-KDL[E6CTBb/A2^PARFKP=.QS3=RBgQ^LFKNZS;@5[.NX#:gBKP?,^W,;ZJ1K/<K
TZ>O9b[29&0L(6c>aN0F/4Y#KRdW9@+5[=LWZ1/I)?.U[Qb(,O/B)DQP;U=I__\a
4PTLa^CP]>bcGbE7YMA0]U1.&FNRCI2INW5,38XT[^gf&QB&_B5d@0<<GNI(Td8+
]384)?^\I>8FdJTK99XG)D[O7;RNW.9#MJ0U+-c^ec:VW?L_C?Zg,M+ddNIA/O-4
AI@&\C75FTFc^#S:Y\&^JQN92=84QdYT9LO@(PeP8&fK^00efU;7F8410KJOUXRa
9@FY8e(Ya,/;-Z&6/b0B_65S1QJ/(c]M)SQ3DX]S-3YcELdPgYDb_56=#)]]S33,
D.#@#2G3.CCC\;A9dD7&B,)YO-&7P-O67A(O0T6aV.A=2PM(UF@0=62T>K).GS?J
G&LMN7N<SFI(#]@UCP=e;a<[;[SM7HZT1a\NJ0Ia&We49:3\d?H+H6[,E_)#d9FD
Xd45B9/Y7=/,U76:;IE?+_DWB:(9+MbBP]H&M3M&4(3<g,f4-YH4-2Kd=1+9:.U[
P<^RVNXOOH/+AKdL8UeT6I]?F^1XYcf[^PbWTBE8N]fKSO7,3RWA,d9;6JU])XBQ
FR@NZVHT16O8M@4H19C,?1+FLF.Qc1?H9\U-&5CS27G8bLZC4d,+X],:I\ZbcVA_
M4#IA<LQ[:?&FJ7a)CKVWdX8V;W(bG[67:R0=eXCSfbd0dPeKXUQ;O2a;IMATN24
Nd3,FIBJNY#Bf9&Z1B1P5H>>EGH_J9#H]5GXFZNN-_Z-\(ca4e#&VBYSZN;:3).e
UP_.9^V175<Q_H<1KS,6JVRNaX(Ef;?E]I#8H4L\L>W4W?:V[X3aPO&_1a=IQH(:
,<L<_GNGLL:9(89O19P2OVB5\V18:ZSG2B_7=;8-#HN\8N&KOgL\19ddgHODERa)
Y3cVA@,WTd:GO;ES<I&\X7#I6HNFSa#:7W\N?ePU#4:PaE[/NL2T(ALRBJ99V>3>
&]M:(X^Y)8d4f(&;AH-MB016EGM2FA2(:a;U]\aS=-5OL&-9;4@b=)6K,U,.MIOJ
1f8aVS>-QdMcYPV>O]U9gAIR-B25Z:Ba],bHE>5Y>BM?I<2>O?&4X8WTYbLGO1XQ
B0D5Z#V8/J>Y60_>A#C]@<0-^TW9f34O6KFDN&9g,eGE#-b+N/JV[#P9M]M]=cgO
LVUTcU4b0f[d.;LU_+X?W>0L=>b[6bdf9c_K+EXWB@dI\W-+\^:Z9XbT@6)<ZAdL
APaA_e\:f0PA(_g5CLF)e]BaHSQ>6-H-e]fa7c@P;L=UPTbVfbMfdX[CTADCJ7O_
W0FK\:MUU/J+B@;?P8OUQJ9DD/-[D(R6QGd_0RKZ0)ZNJ9g54#5S),A<OeYc<GPc
0c2&)<[OW<e>?S#9SKXV3Mg3_^S+(1fYXJ=4F5[C==a_.=-:,-LcTe=5>/V.QLG7
3]3:Pf\D,W.@7SV:QHP=PV;(\K0.gN,Ya<;aX_AJ6LWU)E/VRTC99H[AP+_eCebQ
[N0\0P.#X/FWA_XUO^1[L+T&XXK#<,1J[SWYI35\(I-=.,[]5L^G0/><=7I-Y>fL
#B^f2bMPZ7,S/#bIX_>Z:FS_/#YKM\SMQ<CU193c9GTa\7#4U1<gg&6UeS[b\dg:
+W(I/F;(aS46\ZJc5M4dU]9MeA1:IB:[+&b@=U-_0A<##0-T=VE(Ge68[^=K5JAL
e0\,aCELAC@f[85V2Tf=6H9L=)PNe_8X.,ODeDI#F.J?GK<]eY_?L,C+KM<\&:R/
?VTS)d.7RHW/F.4g8Df7B3#\S(.bPOW<;ecJ2R3GaY-,PeM/,dOY#@6>4cO44RFJ
XeSJX<P)-P7VT3fVC5N=..RB-Pb#<2I:F/2T-1d=A5\+-#d5?GaYN2)9A]?9S6U8
U,fQYFPMBI^UXd&8JGX^E/2,+:U)KYUT/N<ZGX>b,BDY5bc6SX1c_R&df,<^@RSC
A,^0T[GKTU]b2\@-&.09F6g@L4C39Z>Gd9BMQ?3PE=ET0E7,E^MK[AD/>/UD@TOJ
I@T.O8[CH(f_A1WXb)V.eDd)P&K4>3^F)^U(:/QWYUM22CgaLM(SPJE7f&,4P7cY
]K,6G:;FgM<BM@PE]f.1CRFO-4SU&4f_.6.eP5/a_0O+?)5LH@=aUQHR[(b\:]0a
MD:A2\6T>E[HeT.0Qd],#SY^99NPPd1aQP>A+X^?1_J9R4F<,3XN6\:.QbZ9Ka..
BL1YGUf9YZ4(]7I9b+&?JNeNFUP<+/fN?.];H76<JX\QCVI-BCG1C\.FSDF5Y/AV
d2]IC:O,8;_V)@)56H^)gD]-WbJ4ddV8bEGIUT=H9)1_@X+ZgZ]-8N7ObE6?T9?g
1Pa0[O@]Qa<G&:H^KAeEWF7X0fQ@X==C[HHS.&:]X(3G>?0,9<WTMNGaP(Q,g2.A
Wb1ZKCL(D[KRC,OM<Y5,3e#>DW2Q?I=R9_@5]=D)OS4;ScG/5P4OK??8&fR7V4/:
.6R-4aX+.#V1K=RHN_/bXJ7^.WMLT^5][B1f(T5<REFR54@efW8F<VY8:eRDWBKB
:ORg5I:]Tfb2_[b6F?/NOZ@M(W=,PP-.]:B6DaM0>)5.C.R]V[LaX>.9)^2,JI[U
BDB4SV[STNH=O)MS::)#+5T+@gSQ=K-Q2R\L07L+;7;?X[d7Q]243Ggg-1]Ia,W\
=TS-0=NcE[b?+W-LP2R?BS7)<R-A4&>^FDRV/8:dV6Q=JE2X\.?Z3GA(=JV_FR?_
4@35fSdJ_4ZbCCFI&<W1c:I6.Hc?.LY#Z[Q3U0_EeLMCRWR-C#->P]ZeGFJ(LNB1
b94CS5_7LV_1\XU>K:>M6G?)Y#NTc8VHAIO71?RgNVeF0^EE51REX?b7e20>,A>9
QN^[5:<g6]G<LZ;[C#G^a;AWdgbd,)9PUa&C_K?W0LLE-F97/ZS+408=\5R^>MP)
:cP5:_RRLF&]V_XcY>9)57f^@05U][3Pg.QbX.EHaHO+Qb?SG4AWRU?]Xf48.><Z
L4Gc>)(;O-E[.dY]A[^gL.fbWcR3U>b#[YbGK<2?N4b#OL0D^W/^H6MAEPM/?aa?
DW@_LFd?ED>QK@36L6CL#9L4@9c8LYPN^7YS)^T1)C2YXY/f)V=&QY+Ca:FW3;^Q
;-5OC[KAC@PF0_UbH-3]RO6SRbIU271cEJ.]L93A)N>Ob;KMHNVF0aI.[=UX<,=K
T=bCVS\4XW-FdIHI/;#LUMH6-)N6N)\Z+P&GXL#GM&9,Y]b#\LW3(/1d7Cc+9Wbc
A=aJ8?+[0H5A<=IIQd6,Ab@GMJUINgc.@^EN#LM?^@7U2@Z-Fb+.edED)e:G#;9d
8UF/VVLM:1[LT8Z8N@QAW;,,(P.Xaf.@59P5bU_=BU)b_>7&@gW=;(g#R5:DI&a_
-J7:,[2ZDec0=)DffGG18cOgINTb^Egf4H]&gMg]_B4Z@L(P@N2Z>0WMY-U.9HDH
S)7KJLQ;M5f[68EXa0=g]aOG&CXPXZ[5dPb+W=X+UZdc/NL8W8,/\A)VD/7<IR&a
0\;/a,RH(fT^Hc,\ZY?@\QS4K)Gc8&WG]C)HGSa\g+=ObA_57AR#O,Ng1d<.&\+7
??e;/4a^f42Z389B5cHc;E)52FIb15R)W5Ab0eFP>PcQ[V,K0=F?2//8HL=APHO#
\X\Q-]V>;95OI#eeP0TX2C+HBg\00,LCdYVKQbD=cU907=U=AI.XPQUMAK;Z4ZR.
_P\PY>d@WPL0D59_M;-XQDdRN7.F:@(CM?fFM.Q_K&0UbJdXdYUW(=\GO=G?2EE.
X9g^S[XPHVgTGMQ.c5)FIFHD1K-T&Fd43:C?5ITa[5SVYGSa_R,e],Ug((8YL96T
AaWR80OEHK^WQ\8NCC-1D:-_aCBHa(;a?EX(B#bMO;RgGbHQEY-O[a5^<RVBgGSI
1PbW(9BYQe4V(0](.<WQDA.K>;8>L\(_X5?ENS);bb+fGgSZ@(a9ZM]747Y0FJA1
f?U4e/_ZcZ:^)eY96;LGL262-R?+=SQLgYIbTC](N6?aFRb:(]-WPR6^AFY0gN4D
b&]b,A3]F=S465fR,@[=[63Z>BNTX^B<2=G71_<BdTTS00g>E,:(Kd^2(d?\611H
TD@+VP29;TP)c?M-VL@Q.2Ya-Bc2Pbg@-8MUOf>?5)>A747?+=-^7NH+LXA0?L-3
d\&\ZJ&^#H\1EP.MBE<31_fHJ^E<aH?O(b[,T7X9gB7E==Vb<GFBZK]-BeFDH)8)
[@PLB04#<I^U/-S-THGAL>XNJ^2-IXH8D6ddPBP_8\Y-^&6@JHUC/4?E&3<_9(9(
>5M&W8)gGBV8AH>7EOYQ\]3eDdA),a@7P9X&_LeOfCMbgWdVG70UBfWW^.TG^d^F
YLBDCgb75&)DK^&7M+M-?HVB4&XXSIZ0FV@<A^J6M\>dSP1C+/-5aQ?BRUZ,EW30
NGg&Y?+VQ&2W11EYc02fbFFLd,2>N;TG81)C@;B.4PPgdS:HK4P^9<eY/eB#/:.5
==B>4=<N+4M17BJ67<,KU\ef),CffLQQ>?<@0XL:E?-,@]:P(>cJS--aCG0;Od43
Z+G@91XA#:7Tc?^&7-\9Q7,,X<C9\A?dFV&LFeOMU)&HY,,CJ;^5A^>?c5,&82:E
Pf6@U1&WF)]H[-OM,)<Fa5/GIWcH\>#HO5;0gJY))X=PS]6R++253Z9OX<_I2A/(
G\7?HH:VL7&EPQE4fc1f8e7^1^.5]g^0>gOS]U6-6/#^@d57_EZA&[AV.:1b](]Z
H<Y<VXOD9:?O/LQdT7?VAfR)J0#V51=>O5).6EEEPIVJV#[..Xd37f3[:8V>^@.4
>]DD:V79OD<)-7QKY[H@P[JHI6U&HRgcTF\SEf6@g(<;L2F_Ya:9/>7c]]?+NYa.
ZG?5#MX6@V9gMDFFAbb3L#-7=]C+&@\#L,aI-YZ-K2E:(>ePP_CW+A])5&_F93TT
fQa?M&(bX0]aaBJLX,/+LAG^,^&S_);,E4,PR)TT45-92-WZbAe.J<<c)e^VTZ(N
B9aTfIMBZ1A^0+X0\3=^.U4Ke\Z&.)&YS\+D:BSIYKH@BM-6H9EQ?G;ZCe##Ra8-
?,LP;Ia(12OYf.ZIeM-DXR@UOV>@X9D/MD+Xg@-DfEN)Dd8L=QQIQDcT6\LbV>&0
@IVH=W?T=MVRU\FT[e3>9R^ZbB/-8WARLT8B#C1R9f#GWdJHAYO1<M\:KdUNFaDI
Sad:-\_Hf>G[KSQS>ea=ECUe0FKN;>a1)Hf?a^JIA,+_2Ua^-=N_ZUFS,gb=+K=I
F;bT/AL#gg1a?;cN@SCH8T-Cb&1]_=[b:9J9Pab5DML(EDA.3V/&::52YOH:)2Od
7Y1CZ.G\X[F9Z?X98VE[[]@):M@/d6)0fUWa]_B-1N&+5CX[2&c^W=D[#3Z45XBg
DCgMREN=FdYbUY54Xd>2<g^>1H<@1P@.^=dZ:(/=c9]-YEVeaAF@8U^[?6^7:17H
LU4+;TYP(?c#;P0G@T#R1,cBcd9[Q8^29f=T2gaXWA&E[-dG^,GI41.U0;\ZL3PS
b-T?0Q<VB9O&C)J5<@3f;FL(68da-2>#P].<[)+H&[>eEd>]ECc:QYbA/WZ11/a6
e46U.SI+f0R\G)P\<N91+W1]^[WS.cCaJ98.a23Nf.F<U[Jf;X,NRJX_(RbEH:1^
ZRdU@DP3+c//.I5g4O/dCE[W&V?15\;0.XFCSW,O^]W&_ZS,I7Pd6LDDR;7C0U@-
9DcF72bF@8@GEW?fd9=,0>U;,7NIDO:_063e:PKYY_8>:2;2+Sb\Fe/g-?FEL0,0
>[d+Z+8U6eR>)Cgb<XbZ.c(50b:ITYS;YU]U.QT3&Z].K0Of#29;_e5OJBa.:GM[
a6B[ZKBB^SF&]IYPO3CgcXX>I.:7a255#L/7_WW3P&RK?0TB)1YaI8\f2-9_D\OY
2NeAVRS]5Yf]PF8H5]SPAM=>e[CH35O^b>@WeAPDQ2c2X?1KaN;LVTcO^7(QSC0;
A/F0fOSL5&+[C]QX+<c@/QfEHJgSdZ>UVV<TG=.=@b^(/;22A5XM?cc296bI=A#0
SZ_3d(V<cbKcd.PD\LaP0(5AP13Q6Z6K6X,(c:XcEN1_C=Q)6W(XH-LT),@(_SSU
EVEBTE4EU39W0?[SMPG=^S>TF(TT()AG7c-)SFQM3,T032&[G>SC)JY3J.EKaY&3
HL;4c]NM6=(eT3Sd0B<dDZI/=D^OOLH;&7/7c6OQL=#WdQ,=&(P[B(91N\>ZS.a1
gR]3AdeTRMYXc+MXaCH]Z/4.-<S&e]:67?5F069c?=+_^U)cdRVC=dQN]KKGTACa
WGVeUO?GKTFg+5X]&>dcCVM48G[e<g/Qg,<Z]V)I6<2.#Xb@Tg-VKdU8>)NC:;=0
7&b=#Bg<RaVdR49O@Q+C(g1FMQ/@A;4A@BM8_R:e#f-+WaGD5)RYNB:VJ<UD#<R(
4bJ\=L,2a-Iac<W&_\7LG:H/S0[KX4BdV\,d]4bgeI9)^FLb6\MU:]>6C\5^6TVN
.ObKTYK92TWZY?>\UI@5T0=GA(KH/.Ng?4X8@/19S[AA.82)/)4=.R,Pe][N^V[<
5@cA4WP9(<AK=&Y9UCK7=0TH3F-FgD;3M4;A-cR^^#MF7c2(aIbVb_e1,,0MI3?<
<;Je/Z?<R7eI9RGD.:-DJZWDKO??KGd=6D#a56SUee@(^^\4?S>e,9Ra\;FIYfWN
_TA42J]AE/DdJF-?ZB]LC:?7;g4Z=UHTfEcACXVaDN)O<9?TL1&#[ZM(6gbgOU&J
_253=VY_MSa=+L=dHZaT4@Q1:S+[Z8]e[<&K>&L<S/g83;0<W)Q7I:#ZBf64L./b
bQF[;L_4WXHJY8\_(A?B<ZbdIOJ;dENa@Pb3ZR+BO2VC7=;3Y.OP7-7LVN@-(?OI
.;]<Z=26c99MD0^QK^E7.Y=^beLUZ?;+G-K\a.T\]](gPf0La3F2(;??9ZT)L/d=
a,P9#b52_7\B3+L&)e8e0GG@0IcZ4WaH<^H;M@8+5e\\,U9P8112AcVV#\_a65JU
7e;fC4Ya2<LADe:<?B6;Fa29;Z#\WbTUT5L)[JOAX\O91cTZ8d62ON7OgYRM:)7E
=X_d4?,S?TeI>ZY0[cE3D-AXUWOIaOQM<]]>2g06a:DWBMTK1VTX;)=9VaGAPTgZ
N6SIOI@dR^\Q>f,Dgb@P_<<-DJ<0gJ9Ac#ZS<1?1]C54?RdEGD40BRLHW80O7S[O
8P1WT8.43+_eQfQ_7?ZAf67c/ZdCL)\U060.;[DZcZ4fPR>A#4IT7B)BKEL04X>0
9?aR<EVbJ^C::fJ#a00>?Z5(XPQ<+[02/=_31BQ\TYFIWbe^1-F)CP^/8WP_b3Mc
e;_V5XH)fcIb8GTe]>,@UNf4MfPMOQ.]QWA1+DXE70XT2?L:-2G0Q+fSZ\WG,E.c
JFB1+(Y_Q0HF7FUV@0/\f0b.212\bC+8YNf,U&Y/HEc&+D>89(N&6gXK7]W1H]eI
9fJLL<(,b2(M[VKN#dN0E./&7/f)CK.Lf<?aSF4R^4ZKV)L8?9VA&NfW@F@=T,=g
3a:D[Hb=IB3@0I_59<7XE2F,b#7\S,,L&LY1/BH_;=):ZYP<W1=JJ+Y.f@_NSdA?
T)dTY6(?U^&?)NO@a&CWLZ)IWLW5SFPU<YEbPL;aCECI-)9)JS=,g5IM,]9K^WR9
K1(9WV\f/<Qb<87(0g>49_,ePdKEaWN@1e07c:abOSg[2c#=X?(Q@3Qa;@;)[^J(
&W&23B[LALKFB&D,U3I+:daGNBU^,Ec\RYGB5U4a7.GM=#&/)c8M<JC9/>L,CZN\
Yd5=_X#BACZ=>LGQ;fJG<8K=SI^R02Z^[9_<aRgCIVP\:/-R-ZEIc<OeIPVKN4V4
^0Kg1B/FIcNIIVR\Ve\TC)T@9H=\B7U7[SDN2:8[LV?IQAg;JDV?B18Q/.9ReL(5
DXP8@V[L4;MgS;-:JZ00?TDO]CC8ZGU_)Yb<Ie,_d0(ec@bP>\G@Y5Sa@Q+3F5U1
HH[EJWST7I^T+Y&K)8]ddd1PNFb:28;&.[KWg=bZdE-?d2g/,bI]=\_,.Ec-e-I9
X_fFM^,HEd5=2cX)[^K=cbE?+-L=[38GK^a0TUQ3/0/BcPaICUc<+NO<EgW[RQ38
R+JER97eN?,SS6A14^>bIUdPa3bZcGH>P,f\(079?.fL.dLb]/DV]1R;M>BL;H78
R&c=2-;UDLc&GO#-e2T9XgWE1c^#1cLYM?\:ZY[#9_9:<Z0YgL0\4TQd0H+5PE4+
X]:7R)EBK5^MbaG+7WVUL=(0^Q8b=\bAHOdA(1U3[\K>AU/.6<G0+VP=+URgVHCY
VAIOL6e8bbYHO4PIXF^BX>cN19S8gH/I)c[:_);=7N6gKZN7W:CLc+56Q835a[.D
XBKBR<5HEY)Le&=I@BK,^B:1M;W#3LYLP:fN\^gPQQ2=VAA)-Y\6O0Tb=J#MbWF)
OfeM5G7YTHHDG-b1f;W\(<T[W_JAUN:G9N@1aP.#[S93O;_0BN>1-@TXJYZW\<Hc
H626Gffd=V-UbfLY,0U9LC>U8L^e]a-a[++/AD-P9_9DQ>892>F<&SU]<63DA(+I
a2#5CMV#&@.)=.S^;J>EN<?Qe)=KfZ4YVLTc8c-S[&&W:Y4[PdD-FN4LS.fN5Kc_
YQYf1<HKHZW?QO,#X\e>I[PSObQRUG64L\KW@QFNeKB0QKS=<M[<&O_2?\N#dJ;=
H?\]YN.84dZN+)THWe6Ec]W4gYQ?eM<c3+EI(]VA9W;+ATM6)5KL^G<P9,-O:5)?
FW6c>SZ@Id2\RS14@ZC37;-Z,H;08\2/N0(O<3F<7164EKL-DUSDNe(RDCX3X&2D
5Q-LI/_&-9KSf;<VE+7[0gbMI(:RJZ\fIbBN(=8EMg/&?3RJ[0)(:7C+WE,#A=W5
a[cc_Obe&W?EL9/f6H.-+f5=565J7M6Y(eJ#7E#c<?6aP<BZ+?5H7\:G>4?<R:IS
KB/BWGAc_e.Y<;KP)ZR[KFYT--QMd;#6M6LM<dW];f&AX>3GH-3\(KER-@GYdV@T
<??H^Rd?&A)5-M/^789EeFCO=LGCH[b&K5[W]2:&79H=MT)6OE0>ZV_aM43J40IX
+fd;M_S^VY>E1g51T2BL+7a7+C_M.LH<[\<f.Z8?4W:WP:G>71:0)</@O+\W=S<A
\.3L]cK48JY3QA;3-I@;@]A+^e]Xd24TO7<W\]&UJFge1P2JHFDAP=?^\bODSR8(
a6?8FFG7.;>2Ob/GMa0;\/)&-f.<DOaYX=^1>I/\a08D1U].b>]:V-b8N<aaU1@I
-2d<HE3W0)B483I@B/b)K1NC3?[/8E@A,0F+acB.,7U1F#(IXHEb8<I\e.3-0@8W
TB;5K95cd9,XZ^:AE-LQC[(S/J4NT1Od]:U(@TVD5.M+_WM.8c<&PE7cM,VM[_8f
B@.C606CF.T,F[eN9f)-KU^_F@)b_aR#7LZ7E+P]&K.GALD5-WdVe;:OCgW>N7<<
^4;&A[^TUBW216D+[efZK;W7>M1,B)+;]UD\W.FPLZQ(04fEL-a:2P1Z[R7<Q3&f
1.B]I?^+V9:99^=PL<5/R<-SOWY6O1X\-)S,^&QEaZ;2JebD59MNCYH8APKH](aW
6P+R0dc,4[3D.eFD;YC/374HHLZRZaf@L&E[bgO9gO^+cXFJPd3A\.8>)DTX<?b_
E,=Ib&X52cN6/Q9AcOeSW+=4(\<M\dM^W(&ZYYa\I20ZdR/7efAWQ2dUbE:C7H9[
;\GZgOIIOKUe+4_N@e=K?VgYVa0eG:bO43KE>AJHTZeS?=e6ScX\W]1A]d)2G^JJ
V/K0C5@e75,a,.\.1cJd)+7>bSSgD-\^PD-F2SJ[774GL?,IaN?3^NO1&U4WSP_R
Q11/GJ[V,@G88c0fL(63O-:#@IL32Ga>2H(@e/0dUG04MA>9FV):6]#PZc3C6)2B
-E+6XQRD]5I2AK[/S&I6_RF>1>gQR;2IAU(,#^a/OJ,3\)6T<><8>U[5YIAK>d@9
9D14G_F0Ra\9B/-&bZ?KK>/8^SFXYPDGXA,9aK?Z);6MfdNbOI0XY+VJVdH10bYc
?9<SLA^GBOM[44MM@E=7/5JLGW:X[:,HZ9C0\D7ZD),B::2A[KYaD\;(^2fG?T,T
B0g4O1#,:4V70;IFf1W,BWL)&N))M39;+&e\G=6260(Q)JH6:]D?W15(ZR9EBPG@
JW6eYUG=TK859eF4Vf:Kg?Dd\LR_9eM?9CcL0([7D1ME?0E6;7XbTGULGQ/b7gHC
\H;Ha2@S0WP;QBA>c,cgO5J/c#cg[O1C]2E8F8XR\/T=+b)CZ.&/P&H:e5&AP/H0
Pb<@0-fKcUba9E-He^S5VX=&IB:F,\U-2LB+RG-<BDFX.D]A?0Ode)6CB)ZH&4S)
#UWOfOI2F@?.X&LfV1O)F&),Cc=-B?@&\H#\105U>]7NHK):+?SI2,K<faL2g+&/
_^V(C/DJ>U?U@51&0W#KDN9\<EN?c5AD1^6E.0293XJ^6XKa_#<#]6K\MA?e-[5L
9)^]KAUA<<O:ANG2XNdg5a@c3eN5V+E?^HL91YBeL?HZL\8:bRTbdA>DOB21dF3#
CL;a=(Ffe[+L9^+4L_R5XDB>2JXIg(GdObP7)C-_5?d+g(ZFZ#cgIBBS:A^E>=:U
:G-D(#N<:fQ/@.XLMB:?/d(F9<FR>)9;+\G(F@AS,NMIQ:CA-KSf.X_&(NC/2+NY
BL.A>80&FS6<PPO3HZ4K39AXfdIB5=,VSfQ_4&g-6P)7OPJ=-MCc34(GR34#_,-6
L9X<Xe;5@g5H5X<N4Ob/XIO7OLM#9I@d?Q^-=3,M\gC?,DV/X/7?>DJ#HLX5^Id7
F#T+(KHca>GeS=)dS55,E^<:<PN-:Wc>=N]f=(+R_)LY/b2WK8:TfQC.=1T[<aae
aU6+@;f8JQM=&R+N@<W>AHN0+G(9Ceb-_]8H8cX,[)b5JWT.=Q5-EQO,ZBe:TJWK
SM0-\TF@Q?_PP-U5#bVRcL2MRJ5a\DX3Gg^2#LJJ_>AcD>c8?e>];__;RM+FAT(>
Z7>FF\S-WK<Z<N#C)O\e9WHLa^(>6?W@S/c95_6^DM2gaV5]#8VJW5#S-BNWKIfS
H56#1YGXIORF(S7WUBaOL=abe]JLZ8FaT;/cRO&/Z_UQX&c6VF@[444MfcCF-=(M
5DNU4&&_19Hc-C8PNGCCc\3WK28BM)HF0=YY8^H7a]MIMB,O?7.aeTQE=28TS9K&
R-gecAafFcCY>R;.R8XX2PcWScHI1\CeJW1M<\,+IgD^-d;UK/\,>P61KFJg2G>S
F2)Kb800Rf\PP=)=\A[9g&RT?3,UVAU/B<3d7P9KH(/;AcXB=bJ+?=CEIW[YRd82
=a^3Q6)-dJ?K[=Jf#NQe\&cF\S.VJa\]=PbMYOE5<EOXF^EfC6Z5We,K77(-^?:@
b=TZ;ADKe\;Y?9+a@(6>QOGOA9OF9F:BY99XG&KCYE1+2VHT/R\ae.P)a<;c5@9^
,d99K.#0[8K<fOO-2[ZM8K,B[?KK#]C:\C/[VLOOEE.WgFX5g)UbF&&I40)UJA_F
Vc:=<,SOB,I#V0@#BG83a@COELE+64;,:cc99->W6.6#HB;M_[,=GQX5I^OM&=Je
JZLWQe9fN>?JI[>\DZH[X9X;P6,Y^-.76+@=9S#L;(=45OU@S&-P^:9C77;I)O&Z
UcVDOHGXbJPQ[VQ^KWf]f>a8Q5E?8b0@UALEI?_[J/3<AdLQ#LEIXT)C(7,MDW\B
#K?)@X9Mg66Q0E/b,OPAb+XN:A8H5.?/,X\>:dFBJMD,>NQ)NY[RcJQV]3e2=5g)
J1D)gOK<8X2D@6OT#[TV1f(>JD2/,QO&WFSfSR6C3\UVcK^MRK5HEEZK++;:8=\,
+4-K@5T6PU>cX9ICU_/1+^e;YHE1^>Ce52BW3B@[[,;XIPg/K&L,@+T&ZP(R&9ZM
CRcDIJeOaURL,KE^5,.:+PN-](J\MSKGG3>><\#2(1R31O71^0?JCQLaGe5G6T\6
)(K1:HH>2XHDb5^.N6MP,c&dPaP,8G9;4N90=C^POF,DgK>88ERJ314\W74DS=3+
+:d3f7D2M\N0N@^J)XW=@\WD4^Fc=,U]GJM-8,7[dS3UIHU2WAOJ@6UE1aNI:KVU
3O3IS8)CVD(<b&?/\M/XB:8,,WQKI?J<4E\_22(e\_-NOUF5?-0F7W>;Kd[bDW&K
>8_^NLIH+\egAe^d..-8VPbFbO&GG?FJI>OE6&g1RIR,<4]D(,c_e0?3V5U5Q-N_
NXe[.?C5K_S@X(WUZ=6fN89^.<KWIaGL9<<deP_4#(K:gM#O-8+TR/S<NJWXd0>\
36.U\&FcA6JG=Q^PD>8d,38Y_P;gA<4(GU)5@gIDW]P4gXbTF7#S<JRGFcH<d+,X
RS<-BDK55/Y1LNd4&5?8)C0.N_TZ&a>G9PU2?)UV[GB>T:6A8HZ1/0?aa>K/8.f&
52-]g+AOZXVdb8(:34X&_aYBTQ^>&1XeROR4W<f^]VaX]\SC\N9Q&5N:a>.H91M5
?JV10W=+Q5<CKNgLY7TW:+G=A5T5d1cT0RK,XWR)+ASaFZ\K8DS10\(-9)0C:ZK)
;GXW9&8E4Gg25B:^MHG[\]STCe._AENd[76H76ZLC=[MC(@Da70G]P]gGK8Q)Z@J
Pa5UMLXZY^e(T2O9YK^U0?>5bICQQ7KVfOVJbC4>)DVQ#7(/E(CgYaVRTMX&)+UK
D3)DMce9c)#;BKe9;9D0BbN=@8?LOI@364^\#Lb+Wd]LLYQCZ-;I5E]M.a^AZZ)@
YdOH>27C-3:6&9#FD5?.E]JLHKYc[ObeSe2D(#R79AHbOA,9B>Me=>caQ_[6:J?#
]_(b79U4gg)gDO]T4a(SgBU5W6IP:G&3c)]<a72C]/NH<1\^ZDeAZZTaB7Wb&WaB
R\VM:HZH))OLD[C8S_+G9b/H[FZ@\>AP,&=O(d-/ZBHNIg,0f-GdQH<V&6:S>+b;
6,Qa@SQ]3fNUO^/<g)4SA4O8RR@e4-82T@KR\MeBH0R^dM7B>,Ze_Y#S=>,3NAOY
^C]O@a+I+U:<ZDROUZg.WH<D6[36D?G\U\:.F@(6bB+D<ZQW=Q8MDS2Bb;A4V4D4
XI\W0I_ND=4XgC]<[=F7c(U(,CQF[>>5^F8HS97bPGZg<;WOHF>&/YFXSNL?:AJ/
HC8W#FQ0GEeKM&,+90_g;-7aTYF0]N/\7T>OE\G@8YVXW3VY@UO:R\D2Md<]gPd]
[K17/Pa(gYIT/39@P]E&-+Y14-[T3-@OC?1gBd1OOb1,ZHLb1V3.U@ZgK;8fJ3f0
?G^&BW<_IKA2LR.;5La:H4:DV.F8+Se,78UO^<JeHFKfMRORP0N\SE;E09[8+RG1
3(UTC]D=R9(-N(J6J&Aa.C8g)dZV6fg(WeD2Y@C4W^:e_;<A:eIJMTX4bd@Y>BP,
S8??+=P]Vg@C-#I-P._IcC6W.R#7_911^D>MNb=2g:b4bQ0&A=Q]0Qc0(CGU;4S>
N\PW6_.GJQGQGJA&\YY4342[L)Ja6+2^+U327>(OR5Ad<O=KX2GHB72^24e/8<5_
-S&MA#9V_0IMFebYJQDe9X.C7d79<_/WC_HZ\&H,a@C;O5Xb>1PKC9:MO]gD7EGL
Y5;49@g(]287a^2e:VYOO_OdNM7eISD1]X@3Lg?K.?-NVE:&a+M5;1NI(6@QAd(P
]C4NH)_4K&\QRASR[eO7:>7C0^WXbK0PF=R#Ob+ad+E7_N:N:QO-A;R-OD_g-MZ1
^_XVAXd3\aCNY>(dAS#,(SQ61@DK=31L[cNL(E:@EdT&A3=;HdHfd-.<HES?D)5I
e)7eKWJ057S)=/-CTQE]0NC#^;+19b7<R(/6\0]4WYH]4^8.^:&[,3MTUDV5A7,7
]Y:I>WCYf<[]1289/^UJBDR--VdZWU/KCJV6QRdH=I&6@eV?)C&W^?^OK@&CRG>4
#KZ@X8CU=H:49<0D+O7fe5+9K6-WA63cGOFFVF4XG4>d&dD7]UJdc0X#b2=-V(;H
ASA@VMI[\0(DC])g66)17XN^UO<=3E1c>EGI3S)g200VN)3Zf7@3fY?YI.Ef&L9Z
g4[<YI/a3TK.]4NCEBYS>7:Z9J;,Q?]>&;PA>->&8cPZU:(c;V.];)^3-cKg-[eT
XLY92218(FTV94JbbaN:3UR_YVP_Pe72)<HMR(>c)c)1QIe9I]\F1?O.XRBBb?,G
<EQ5@Je\1&:I[8D#AW5C50R?4B,?^45_dM6geT459V69e+6O-Z[,UIO#>]TKf<U(
-49SX(Gee.D_c:=IW7dR\,gS,H/F/JLb9Y4]3c\6-Cde6+YSXV7JYI81.bJ]<=;b
Cd],O:K2T&bBcb8L3D=8_NG1SX@?F7,MTXBYJ^&]CJ<[V+4YLCKKXZ3W4IXU7;bB
56=UW,Y=ZRL8g/DFM=?B<BFc<?_W)[5@+-(CHC#+ZTKIY54gbC#;?FO>@G9V>?3P
RZ3WAf7#^>W(JOZZNJ^QU/eg:^\P/FFE8,P=(:DLLUFeQ2F9P6ce9-]aHL6\K(I<
4bE(V,&33QT@\@6\:U/;59QE7H6K8]0M[KD\A/;;<H,-TRSP)#N\UA.fPL+b0]Tc
]U>OVA+7a36FV5\69<da,d0.6-Nf1,HUM0CfQMXcMdGZ\)P^/8,Ac(KJaVQe+(6[
b^V&+](MC#@^E1adWTB6PaRMC[(8eH2-eTT@E\<QP7+@>FLG[b,C/6Q66B_@8CZ?
2I4[Ua/La9-A#f&\@BYZECTB^dT_]a)^A7VgMG@b6:@C6R>]CF(-R3_\L)Gf2g/#
cVdU0L8W@YYU\WLKPMKga4DfMA2;\@FX^\](I)?\B;)=+0#[\e7Yf\3QKIaaJ7@H
IIa1Y1EHeGac0_f1J+K\>?DOVf][:058K3cP2.CC]a^=M&3\>PQf>0@OSVdP3fBB
]97SWVQOT[f)e\f^IH#D13/bV[_:d4&8[YaQUPK=C.GY-Vb)Z[MM?J_<573da4fg
4<)N2dDV[AB[071+)MaVB\3#_bW:]]+PFO?R)T=>b+_g8I+Y\(9,??2>Qf;bD5b<
W&O,[;UYV]N<KJ0+].TH>eK2LGWO@I8M3d#UHN;V8eV.&T0S3c&\QgXT4#MH+gDM
c#)C@SbY6?;EB9\YZEc/U5M#7]E5+IL\J@F8\0V6gZLY.#2&IYWUJK>GSMUVT^+d
[,REG\\DHE(T&<)]60GX=cB\F6gFc/16f;B-M:8S(LK?>.Vg.Ob5b+ARQ/4]dO8a
9NDS6D#b;Z?dUaaV]V(>J=NeJKY[eK#,/,3US-W2gCZC3D/Q.#>_&@9D(6/U/)6-
ZN^;\EIb4BDX^eI<Te&/M/cQ16]\e,98C#Y^AaI>]2]U^4_A9@GDXA:gS4_]+bec
+fM4(=dg,_U+AE43W4K#;CQGZ:Z?^EeAZ/#W[LeXI6ee:gd=)eLe0cMF32^MMLf)
><T8[:YRBLJOdQ>\J,^/+M_/R0(A4FTPSH=9P)dDgTNFTSb<g89dD39J8ePGI?50
><#O/H#67c7&<RbMbYQ>=;eCYJ.2K8[WZRGQ&1A^T^<,[f6[+T,,HXA/<//Nc4?V
O_KEZa9(@EPYe;U(XY-/SKH_U?S-VDd:NDH@4?b0NY5?IW<B2cDMW1fZ1T+E<D+5
7TR9/3SJ;\(K_GA7=K7_5><5c1KT<O&+gI_^@e1.MI&DGK80ABD#:8XaAfO4T<S\
W,Zb3<7VF.>Dd7f0AB79QBP9FH0PRgV6HG:B<)QW&L7M&)6CfWZMbDDYM/7M]FT:
g+F/&QZ@f[J)Tf+OE3.Q<.7ebV,8(cGB-4M)EXB&d@G(a_&X?-VO\L._aJ[52F7_
ZO/[b5T+KP)?;_21);+/#L+\?5Re,7X[a09-84e7RIAbbXGN2&EOU?5Z;HT39dG+
D751WVYB.DdT:L<Id1AU^<&3[37Q+N_-fY5=&?@?>Z_@a[;ZVga:W56&/PWK/5Z2
.bYMS2PE4Sc/K4OZSe)Q9,Q&;E#X>UP[3_faI86dY4MUa/V[+L:E@9aHbeMXP.^)
^c.-FFb9.>4BVQfG=[WDf35X_PcBf9I:E,<0+(V=P9\Vd\/b3L3MHa/+,\N7ITFZ
MfaBV(K4@SKDEc8STQ=SLZa4/5>:6+&XJE07]#>S^>dBe1T;S@K@2KL(W/,-8bUe
TWG@.=^23,_IKG;,a()5eBP/\;-f\cATW:S0OT6;OaE2eO2-Z2D]>.BPR8?>7JAV
I?-ZK1:21@PLK.Sae9&Q)A_H7WE7OO[U)a)CUA40RWL&#2WY91^AA[V::_baRJZ+
aHHC.g9;DNgbDCYVR+)72(YfeO@I?7OFKD2@KTR-_;^+VZRE-_[AQcc?U(fM7<4&
2:S-]4/g:<d-ET^G7@8FA#HR7eP9-Udb#:+?1@fTZ:-YBYG?07,Q\D=Yg.V0dNG:
,D9H7NCbVK=MZ2]^;ZUO>:AT,T#RZbNJ-,LVYEcJ/ZY+;3/bQHcJ-#A0[<)_7OSb
FL.T+[S.YIDW=S\PA9S&bSM5f3bZRH<:0U2V.6AF+GFWgI1TG0Xfa265T=]:]f\P
W<<a]Ib@#]SE>g(<BTU2_L0H33OW?_#477BRSd9)RdBgLJFc:=H[d+F\a7EA&&^Q
CgF649M:&=XO=PV=8RRSN3abf2H.e[AT^7CD#U>fXITbY0SQ^<-1<4-V/U1/,E2/
O+WSK<)..4/]V(Ya5J&^]gb1ULbb4Hg\)Ra72EFgA=V=06Ff#-V+W-1cCf+(KSAN
?UN.V&DNXK_\Xdg_SR(8KUCB7f2>YI0[[0>D-1#-Y[5Ug<.:<=S7[]N]\;_Y12&2
7ePTE<1:ggdWG,]2TaI[QG#OJ;1F2)G8Fea6fQ9<X9>H6RdL,b7R5YP82#7)FCIY
3+VbXf_1741SB+<0LT,Zb>HLOR:e/&Z;85<W0>@c)0=Y+;MSD:ER4-J#5SMDUbF_
FW72-WGObO/:Bd0ZUC@MMCE^;aQ_TZTd4R7Q>UKMcaO&R1]0^1Y&(/#MN(8HI:\S
7LRX1-YLKa6+1IJ9IAU6PPRQA-64WQZ>ZSe..bB5SV9HCa&2:Ag4eE[IcHMUS:C(
XY>M2;5BJ.6:.C/G3A9AZa67)4SP+#@A?&(8dS9L>^O,.aU\1H7S[,70P4;_:=V?
@5,BA/<Z7b>#cd&EIIMXfJ&IW6Q)43RS5X,7(dcFA[Qa)Reg.HL@YQ-7<?M0/N:X
E,ILDK#2UBA0TL)aF#DBS,SCZL80d79a+8>&2edP1AaS9.X-+.EbC)G4/e\CP-3E
]#=1P6TCNBcCMW_fN_+@C3H#\P.Dc63U]3H&4TTHSLf3;\K;<,>8U)BK;ZeMWIBR
8?33_fC=Z,0R?A+/SXHBIIW;+S>Z-GdDd&/b1U]GJc3eCZI.Kagbd3?D[F?[<\E)
ScE(Y,)0A@_EDCNf_T6dGZ)2MI]a0F&^7Ca=7=TZN34E3d@WP.E+.G>B?@a:O#a+
7(;2,E5D823dRW(\V-1+4M:P+&:6LY6<2KIAB53+GH]V9(3,WZ0cN37R)eZ]R.[5
g]E)6#0]gLbPM\V_@P\G:ZHNO,^[=A0Q1Dd.=YTdNRPbd5N4H8-2cWRV13Z6KUY/
/:K@98(:2EO#dK@g8X:7&>E:-6=\80YbR418A?feba#@XDd0-K;4/6VE,X(Rca>\
A_>#d/AR1@R6dDGHS:e8Ab+6=.c9Ib[FfUE)5<HS.ZNNBFAaO6H1?8dPW;)QSIR)
6ZAV[e]>4BG,<B.TJ2?_,)O:8;EdVL?]5>ECWHJcD,F7P(CbLfF]2L^QZW[@H[A]
MR:90(dR,8_U.WTC-#O<Y3gS)CYc07L7H\][X-8f=M^QNBR-_XZ57Ygdb0L&V(ca
=(_Og^US]1KCF?B[+0D::(LMRH66HYI2]VMR9(A5O<I?2Q6[JTL,34/4UaACI[PT
+9_EY<KMTU7S4[)_^A:]Sb0]D>)4&Hc<>]\C]VV#&2Z)J:70D,cCYgX-DD1+&L4J
/^.EHeNgR@QHE>;ZeQ^.5GW19C8(7M32fOVX2,E2TZ[]Y=6#<;VFcb;HRQd64c2&
H8KdP0PF?OcWc(Pddd3F(_\/9CX+dA7>;,G<bH6S;5gM1gCREF)Z,#BdE;d-M-:b
]JdH\:6GT/.HC<P?RP_I9\,28\8a;.E>.0.JOL0Je0^YWOK^#>2WNYBT&I]a9W>Z
K&Gd>:VaBd,Z47DLKR-W.4/75(^42_XgW?Wae;KW&4f05ID=9[&eXZDU.A?PSMb:
:X,U5S5/fN=+<X7U4&IUM;8#,)e\S\S7b-QS.Lf0,YFUcb@_b_J1O,ZFV._>XV-1
8e2J)2WU18f?QI,/XO#ED?=;C=MeUb3H#V?N<E4TN9e:PdI;LAV#=#EFe;g#WS;0
HO7G;PLaD+.#O_2(UZRPJ5c:M\6Y@O<#7PFIM/[4Q8&@.OUL(B(ObFAL612W?<HC
e4B.<c4@7K>5&,4HZH9S?9X:A4QVQ770=b<CYFb?PH9O?S7+7R3#T_Z):Je8)J]f
T;N4D3GZ1+08O@g&dLN=RH&@X+Q3#M<TN[,#dAV,MK+NI(N<\B)S#3J#G8ZYIc_+
^^OOa)VG?_aK2H<3]Y]P@.&ZUHN=(KIVS]UJL7AKa1@FFWGUd@YERUNK\:&&&73P
>);a9(OAR]fd-]g?_5/5+V]=\5DQ,=fcY<BH2QXLcaAd9Tc.(:f2@0QUN5IWaHMC
GIHW\B@/1=Y-]ee0@I)?d0EV#K1YM,e2:VCNL^?V&\cc(W]@Z(2D^U]eTLC=ODE3
6;+A9e^?LEW\WLXK#aHPPONQ4C/3:/Cg.-gX5SKOM]b6XRXWDOOAHIP/ZWQK>Bf+
W/ASM2014AN^dZ(=(/Z/f9NT+c_357b+JZ^+]HI8RD9>^2#=\NUZ[5T8NbM+L__5
QX6DU^YU7Lb>,d[0S[8]=.7SO3X874VEaG,e5DD?UdGe\Y9]a<U7]P]Gf7ecHGB<
=+ROeQaKMeV\T,<;<aW2CGLBR>NVWTag;J0#I8@=0BJb]ZP1b(HRD9/EP5I/6MUL
78@NZYbA]d/BTIQ]FS-SfO7K@a/U=H3C,\FAX7FYaEYa?,dL8L>:M>AdIc=W?RZ[
fb)B?KMY6YVaNf9HTX:DNQda92(4?5U2ND5gHFWQ&?N2;ICd+[EL9:^J:g)G&8+=
8P#3UM@U:Te(bdcL_/H=e_b?SLPS_^2\NE/#_#?#0<@GZ0e.\ZU60FUId#+4]TRd
W]DWAIdDBK7J+\(LUX<DZ.G\F1E@5SfA9_ITX7YH6QH-9ZObZG3JZ-Y-YI8Ced<,
<bK4J7J)1#T0P9gM4?U(KC+c.D77cgRW2?cN6>J&dg/J@-ac,>.0CcbHa.@D+FC6
63^Y79/<S93aNHQP&=V3N)I:Q=]HW9D2BELQ1aSPLR3dc@S:^H7[SWL__U<Ra#VN
(g;-_9H-\N]J1)I69;WIT4aG?@g1T28bdF6=Q0Z0#W.>-0]G.02AU+27FUe)F8.?
:Q_a35,6dQ_gfV3<Bd&RR#<_d[:N(_gMGIVPBFFD(d>P=eLIK][f9GY6CHG[5=5K
6\K2g6HFFfReb9WF9_:2aT1290[GGgI^?Qb,=/HS_Z-O=].C)_S&&1cFNC^ba(#W
/TD7:H+2W6VdA&YJY5cP,>MdF2d/c:/13,P9M029/V:M+aP17Ma\US\/Z,f200FI
);?.13L@BR6S&[V1?EcYf:ILKfY7BUH^7J8:H-NbB7dgO#XKT-7RC99.LW;=,b_\
Td_4e33]eG@?a[LTa9+M;QXI_#-Z&F^X2@O]G&#aPF;,eaN>#.eS9W7aPQ/:IE]W
JJA-<,Q62>Xg_(N^G73YUQeJF>a(dBDf+fG=C,BCS9,C7X)7DWcgEQB>RBBJ8V<S
38VW+]:4SE5ECL/R9590P]F1=Z01W<KR^0M,)ZaK3T-?8e9:XX#.D&<=eQ?+::6d
ZT^5IB-CZ+#8;5a.JUAHN+Oa&#_24[0BaJe^[;>2b0f)>-\O<GA-N].<PDR@R90f
7S)cF.2=59N-LL\OQ;ICQOJgR#E>P5JVL8;O.&S27B8V4G/MfS/e@RE8bA[H_?C0
31]U#>Idc4Fa,b0.M]EU(6SJ?DG6,-f+6CQQbbe=e,NF5IVMX=;^-OaOVQ63D/cI
6+H?Q^VSF.[F;ag_[HHX,>V<Z.[e)RI=4aYQ.2:ZNKFDO2X^2.12.;M.YFf+aDBV
Q-GH/(5^.NgCV43T)XEGHOfO3V__bB<8PGe2Z1HLFP@;4:1Y_]27GVC\UBbbH5H4
b]K@=W9Y,eZ4gXDN/g6.a,RT=L+b+IgTdITV.ba&^P:(5>ff0EF]P(OQR4J+QaXaR$
`endprotected

`protected
X85g2]/Kb.Q=#;=&M=<E4.R^R9(37?^?F)&\A&\)Qf^?4T;3](3Y+)Z_UY/4,64^
=?44OD;IB#)=.$
`endprotected

//vcs_lic_vip_protect
  `protected
P2d(#eR)W_#VD@^JH@\a+</SIbI17E9bQ;&)ZF75P<HF=a#)fQ^E0(B0H,[cWe.)
^I-bc-0#1<cTO:GE+9NX2+;GgGff\CMR42d2dfQVU^4&QR6c,HUf=@+KQ+:H?.Ib
?1+^;,B-/f4aPcK])XETdNA3TfbR18L=[D5g/cPd=e]f:J)=bC:Zf))ITeUFS4I7
X?C;Z:769D]M[&&4CZf+MGEUZY:bVF\4J;=R6HeS86S&[U=CcCffg4cI6=^\Ogg9
2A>6ebOY#@b^U:9-=:YGN4N+]9aFD<7-7c7BURJJXUC[AY\&\O#G&[dcObR5:=\D
D)8aH-7W?FU&_:3T?a+VKKfN8QIW@Y?6WLAL3.9aRf?VM#DVc<3NFfM-4d:2^\Yc
OST+&:Y5)F3I3[dT4/IX<W;9VDXG(b&gg:D868]2:BI_/fNA:XdLOVI9_1PQL_CN
Qf\/Q8E.9U(=HFaYS9dUaZGH)817E,=fLTgQ]]I2g1fE#W2f98<Z\^^57I#1:L>1
TLYg2QDZDU(aYY[NOAGb2E>N=EKa4@bNJId;/V/MSeR^J&JLOMP;BbY&Lb/T)E3&
PHZ+cb<07@8-5VFb,/<N?WE9V2dK&:45;a,:]-c>1SPU.+YB]G#feB6eM7E9S5ZM
UbQ)>[S+8(fG(GTL\&R]=C&]aP.1RNWTCU;,gCQN:2L:Cb02I=-@Jf0e&[.e(@Xb
Cf1PedCMV10;(S9JW;WTSQPa;I/&UKP+4)edD+dQ&AD/ZOQ,TIM1N87;cUA8_D.^
9L)LY,H-V:OM@<(EbMD3c392&+J^\O9f>M7#d;T#2B/Pf-I8?5KS8>d-SW=f_Ae3
#C(Lea(W4@:/0TFd2g,]3QF-SD);)gSVCKc_]POE.L^3LHefMXg)&Ne4=(=4XV2K
HPf(=\3gCFCU^MJUHI)])JKd:CcDF9A.H^6.3CZPG2aOgX&G6-6X9?/7?gE5Xg5Y
8?M0_bD@b[dII?:R#GQGMU;3aNRZJ3U/<Id@bQ8:bQ.#L;BGV)-0FP+:P^Y=8QSY
VW[<4[+d9[A76<FB:?)E(ZYOef;;;GfCN>cB\g<YS1U4.JK&Gd-;&/^2g)EGeRM[
gD=:(7#aD4(6JTK7T/;Z@eLQ8WIK5@7VEO(U[V;/\BSfZJ3&R&PIe1Ve<<@N(BA:
A[O8SYS?WYLI4\#@5F0,#g#RC><9_;<aY2##@@M-12dNUYOPfc\;R5=C_>D2UTE;
O(L(-<:ARVTF/Y1YH+_HVeZSAWd--WFOc;W(+OTUO8ge,TefPeJ]2NZc]30BEBFB
NY;77RDF_8^EE.c/.E)[0?\,A-&?1AGLEad.O,6H1N<1#<Z]:#JWNI,8(SLHe^A+
V.Nb>#1\K1^5aZB^&:N?NKRF+62:I.4<Ke57Kb:?];ffN/ZIW7#\-[F>(KDc;a,#
,Ua\17:?c@7Q)]\JR\-TX;Le:5#M:WD/R6;HJ3OCHDb7B]-^D]T/d<U@F/3\>fg_
,+#U1W-^,5cJ6dZY4@?e2Lea/Y>C?K7E#QD);@5^>,KO<LEcW+gg7,HM43?^93&A
c#eABV5\Z1R6<FF,VMO<^X2dNVCb,S>J>&)dP],ZXP71a=0P](3Ue+bM)fS5ZN^8
#=De-DK)d8[7+MEaSBIMX?B.OV9Ea<H7edK=5=##A^C)GH\W6-eDYf)2>7(Z,N:M
5[K,3/-#+I@_Y[LLa-#c\T1B:JYF\beZLc6dV2,3-B3][7AQ?NcL@#E0-U_4#OYN
2;]R+HEdDP(1\b&Y:Y1+?5#a^/_S[^Zd0ROJV/VUHL6]#ZIFfV12dY=E#TFgc=53
^cFgXSDCcBMO_DCBaWgMW]C\>gZ2ceFC[bS0VIK\[GLJbM@)Qf..EXA5C&E;E_Wd
:&H8f(>-Q@Y7]NeGD7&7^8ff1@bP:1QgF_Q14[\W&B9R/8M9SU):S3_U2e@/@,9/
NYaE=/ZK\[7UbT3I45UR/[gV[1)e6G825_(H<N>EX^RS??L+8_,9:EU35-G(^NA&
[dJ47I16P9\HI8HT_AB0P6d=PK_0[GU]P-M5E2KY1aGcZTGa8g3)dHZ:EZ;[cVFW
<.?fSA3f#U^:Ob.;5cI41KIb.>M(B1^IANI[e?-.BeIHH5-NY5ZX\B)[(=GV4ZV_
VgF4;W2DP;U];6[R4?D;O8eYE;XaSQB(@D,X=+K<@_W&.D=f:W4F[PaR28&H.0_7
)RC,L<gERC+gD37>H[Be0.P_e\AD)HI@-X7<JHG@OL6f\F8edM)=VXDJF15&,/\?
]>U8b_RR(JOKA&DB0K;U>_aT(-<&fC,.G5P>X;?[FVf6DBKd1CVQ)6O0FU-dWFZ7
:Z\?J\@\X4T8NCAURC#HW5;S9046ZaM>OTd;bP3&Oa>W)3&BC@C/_MI1f,5QIWMF
-KD39>Se:CX016G;5eQAeeGWBNHX<\0H8NE7IHAL;QQdH>@Z+NZEf=FVYBa_53J2
4-42@YPDBI,\g@YFe@e?8\ffA96g3F-7^4)PK<AT90cb-1YJ1bb<84WcaK;T0JJ]
LYGI4SOY.+/V08L=\ZXCN7XUG^5V9)bVg:Z,4f=UTEQKDK\d4/^XL<F4<2[SE>L\
7+3#83gOKB6G=cSZbF39-Q.0[_,JZ+c.24]c_]I-1P?L.65+LKXX/OTI+@.,BHd4
I,1_OCE&eB#+5AI4G_C+?[L+b:1JGeKf]GJ?a8]M/+24(e6K<[G3e3/G+6S?QBB/
4ZUe@9gZ&1OG\LV,ga-84[d+E5:K4=6#,1g44C/Sf1#L7F>9I[QM09E)CR[-4BC[
H&b2d^24&?Kg46XB@.df<DL#+#GM5]_:_dJVZAU2E1QeQ5@V()g#)]A_Tb3^=I;K
\/=X&V5XaPIOSFb?>=>bRaT0HN-VP@1ZNMN+G8^.5F6TEH:7J?:]XfR3+8MFYWN^
-0&;EFPI,XOFEW]^O)CIFGRUFc_J64JA7\,M]>8^<IO:gH_M4YCORV2^<NHD4)=Z
Y-TH2P-HecF;9Z_]5SDGWALZ@^\ZC6L\<ba307J4W/-d1P6?N>TUEAWF@37+2&fM
[gNT#Y31:VZg(DYIK\2N(&(0dGF5cILQ))Y+A<:)b^(cC2SX2PPJQ;7U9H/:MOG:
1^&9<0QN\Q4/QA[Y;Sf<G8dMb;8ZB22RU9H#Pd_<HXY>[2-^RV[TL_JH=-QRe<b^
\+BD_0.Vg)&H?=777FW6cSc;e^(,LR+HFLdXMWOVYCF.PD7gRCa[@?EY[X]ZWI>@
@Z?^1(V&0+2PK(ZK,Wfb[T<We_f,f17O#cE:+6=^T8.(DT6e?/^eALZRE3E2J\99
O[<Q=#M5Db61^);T<C,)Jc?f;C(?H0&]e.ZV.1&cR\9QPMC&B7D386L&B&QGE><7
AJDI6#5IU+-T>6A3bL2)EG^W1VZJV0V.I^]\,8#&Z,382,&@MB1,NJ7KH+Q\<d>g
M9SCQ[:/D_TBNIV5?,,_3^M.M+X^?9/KO1KIA,+MFI@U]#@4b&]3)[d3?\9QKIU\
UX-Y3P47(e/e,<#I-Q?H8P+IB)J;H9.V2/,CF;N+&9;_@McUO0)dZeV;X:UY]P)K
O+g>7#C:,7IcV=A]SWGGX/VKF?NKUYW99HM]63-D_G]>0gI>&N\EO046SBKF(WW3
I&0]DeK\:EaR14PY1KOde-FA0e46JZ\)C,)Z>eWIHU@:eQ8G]H68=K(57A6P1)OV
PT_:fD>2.N<KQ_4/VZ+\.dL@BAZ7W)KWW11B+6M#L:c8XQ78=Z/7I(Q)U-04IL5U
XbA\F/P1T,>T;M2^=#-9^A4RZ?^??[&\]1Xe6FDQQ;5faD5QH2C\U1/IN&<6Z73^
\\f<-H]0O.P9IHJgF=^I>d_g,7^J9BNEc6N_\0T;W(VB(3c9CL8Nc>+c=dL(M?SA
3MS[]aXCDd42^WP]F0eINe8EOJ3><Pac7V_cc5S8&D[g^7C[O9#I-KHD09,T6fg?
R0BN<MM>=-:K=9f\J;UW)(LB&2@K-U\H-:(Yd)fNL_6/bLO@YGZH+P-.UP^>=+\E
N?Qc/aFPbd9]3@aHMB:W..6^:8>-KE:Jb5GOgQ0<QH.UdgE-Q(3WM46:bVU)WeAE
21F#e2WCTQK@#.KbUM6KA[f./J#TOQR_XL3K.a(M+X4BV.+LY3P.dMD2f3d:FdQ(
K;JYb_X,.@-f<Q-,R@T<S47?>bBYIU?bES[2aQTQK5c&L<J:\._JTgJ.]?AfK9GT
8.0W6DV1S\8<M@dOA:<#aa^D]Y4c@(<d)=8Xa_Y(0K6Mc(UQA]_Z(FZK6:)C9WEV
ff8M2U;HcE\SH1S[O1Z#;LD=1dC<MFN]RIOeTYA9H.#Yd8V69/@>2V_(Fd[3TPFS
Ld0Y3F9BD^>LWX>]G82Y_B_Afcd_W]3Yc+-_Y>>UU^_GV,Ad.7D)]3VbK#/@FPDd
?L>R<0E&(V_ZS4REO.MSSP\KQ^JVe(f8A<1J-<W>&BQAC^OHT2GKMCeH4Q+9_VZ[
cQ?U[SI^ZYQ)#A93Pc2DKM-NT/.K-3GaB3/P;+cNS/Q6==WeSA;\-GF[a\=@XNRY
<+d.WC8QT74,/AG)dJI5/^.:;.INb)+BZ&4#3L=ENZca-O>G04L;G)d.C9^)NXP,
>[&=:#[F.<;3>96-#Ma-\g^\.LLJQA#D(eILe;G#ddEIgTWa-M5XXIKNRe,L.ZRB
][g,#U0A-D:>B>a4=D8.gWMQ:@_bRX8_4,AQ;f<A\ZMEB=dX2/DXX-2&/2?X8#cO
gN6P\)#)Z7<AScU_,/UR(eKARG@_OHd;/^9g&[<R>b5_.dN3=Q8aY,?:d0?FEcN4
T7d?d7//Wc-JE53g(F:]gP#BY9_#FG<WCdPW^NeUG61UBc//3@-fVI?)cE:@g)6U
6&V2&C.XB?AWe9(K7W-=J;)B->c8?5<4A_LERR=[#@1BA6.A<[_QY(YD7\06_52M
R\+,g^AI8e^3#<YC1[XS>\ff3d,<M^J0MQMA[/EB^1]HAH)#53M=(NX^/SRV^^?2
=S^NaYZFM;aD(T#_E3V&3=:&=aYV9S#4cPM8QD8S+_Fg>123f#GI-82^G5N9B;<c
D#?POWX4S+9dL._,W0CDJ_)1)M_-F4dA6E=Af@^:_5?:92\EeUI]40#7W8-.fDJT
,d[dMccKA/8<\?bQ\TVB-TB+dV8:XAP:1O^Zb-XgT2LgSOaJa9IHKGR9fd_X@#L)
YP3SGVQ#C[1FEZ5SU5CIOF^54EE#?4c&VI9[5\CR6.NZ:;_9UY3]Q[]e.N^W6LVE
OYIKS[+NUS/4138JT&dF8Wb<22ZWZY)?4[ce52[8,@cDa#N,?/NA&CNBR+9&GOFZ
@F8^T?<AG4/2KAgFF[80>VD6fY5MON6?.,Dgg-9dPAFO;L)<1cMNQQ[CV8SSYBG5
?]IS]58&4Q5?2.I.eET#=2AO3>#6cD,2N<6Y>R0)d(E.;OAZ0UDEA76ELH],N#Z<
,G(L+0I1O5=)#)JR(\T1O;cU;#2P]bK4cKg,KGLC-6\#fG(N<O&.NAN#KR,NJ?)P
MbZ7DV-I]L]_;Q_Yf+;eb>B+FP,672[\1:];X92C?WWHA_?JJ46ec1U^7dA34(=c
SX?\/)6L[)>MZKCT#\Fg_@/6;U]0<F?,=<2N>-Zg8[gf:F77((PPc.CQA:,UMgZ>
UVMBPf:]Q->VJ):#R^0_c>BJN5<J]+R=A-A)#ZaI,[K=T&YW@4A)FeBRCOL?QPB?
[U+DKK?9BQ<97gYIEI);bM5R(?X+L(L458Yb53aZ\BGaRRc];9O2?+B0T>\KU5;;
2=6;e/g(,EX;33f^_e@)7;Y&b=Le+Q1LQ:<_9eQ[>/-SB]@(F=<C0N#?#@A,MRJI
<6#^E2B)@NJYC-/8cGaPcEM&cMJ8FFJSM9fSW\U4#/De_YVeE2eD6X?HFa=:_5E5
a]LSJM#LV\XW.AId#/HOeZ#@2.3_V1/0[+X.Ve_0E41(TC94/_,IfdN#/ce9<bVb
5_4:;Oe?B7a4.g8>-(J+eD+e+T_X.ZM@IJ>&0HRdTbIb(^b+]J.5@ef:<,/C=V@F
&<#B4faQEgd9OfYcWf/45T\b/G6U[H(9aGN0,7BaV7(#9#EcN0\00.[d2ZYLgLL&
QD&9G&fJG9Q[SW.=Ag.JN<;Jb2+EQd#Z)4[C^0gP_PgBAJI)7#D2W3T\>.c5RNII
=a=AS&TO==_)([E&C@_LPTg^;5T6,(4A2<]JRT9[UA14H2LQP@]CR5A7A[M^M4^W
Q#-RL=II7c\NPL+=G&R&TDG_cNWO_\3#b\C-):=])A+D\N2C+]_=dDH15M6]>dM5
Q,>,^:/Uf\e:+4bPcB:bN;ZP.J)4]fD==Y?>e]_?^eV;/SA[=f9B&&Z^FS)3K>ad
?O)3(6H]XW&=XSGIFZ.g&?L#UE@R7c(f4LRFL&TE5X[6f(U+a#_S3H&aL8QGcQ>O
a48NWRU=WQP.<.X[8#LZ3YZAX/P/-B[e]_D=WWKaYDYJg>e;9]\\-@Sg#X:84d0W
^bNLL/M<KJZ\)WaC+)(\dG6ED:]cc[;,.L8^WZCaU28aM-OJ@)<LIgWULC]S5W.:
HE#f.fPGf[3)GJC?4aDd(?6,D)=e)=^Uf92Wc5OJYAd<H4bOHG08^5)+WM<#&1OC
M;N#W.8b<ZGaaB+F2@B)Le/N>a,>V8+\ReH52\W.=^9[+\^#[]=F5KWIMK(]f=[R
]3)J=aR(_(<I^9&=MZNAf#FaOd1]30&EWJLU.2N[8=P_W=(_UHI,WfY;S/&NJC<?
c3I8#)>.Xb3-ZJ)fV^^:F3S8/(]G4D7SP1\>^.-O?2J&HT3XMA_^5J69XD8HXD13
e-KE<.<G(NDO57/a67X7eM@T35\B7[R9cGAL;-FCK]>,E7b_7L,a^Y(.4/J-Gf_8
.^@#HW),>9L_9]IaIO,Oc+QeNZ7C<c83b\VM(eD>3c2X<RJ/JZ;#T3@9.^BPR4RX
(UB(PH8FHR3,&<&#:R8X-b4/YcBEDSZRH/J;.1]M>\bX#/B/>LBVMYFVe:<(8ZL9
8Kc^SB+8UQB.BC[O;XMI0T-<J-(E>D-K^FU=G,Y\R/aTP>TCFP6a,C1E9U1fZ14_
6NHbIQf[a=FT9@NR@V&a)+2&@[E+g7eEKdIg2XY.2,(<TgHcVeP.N_LOXTC2;cbc
3,F_b-@IfV-3FXM8NV8AU?Y7Q49gbLHA@cHEV7Tg8Z]-3TU638+L_Q6e:I0\b0Q.
B):PWF;3G@cDA_[aU0e=YdIH2f#57LG4N86:X&d=6eTJ?:\VVC=NUNO5HVaY6&M6
B76?f=8O59HY9.,,)R@a-?a78e/00A._6JM]SSKL?B:F:]<2S4HQ>E5bQCB6E(<(
D>GL6]:/7H=?:8A:SX+.659+02b&?:^?;/)c(4?4HWTU[\eOT)4M=Pecb&D>-X&G
FLS07AVVMS/W0eN.1X_KSNGd=ZN_OFea<E0KHH3fC=Q#B&c6D0+[5cgUX8e[?7+3
QA<8)[T8)4_W?XLa^&5d=LNb0A,^B[49MSR[dB&YH@Qa?MJ=cbVBQ8Yc-Qc_J5Vb
//+-_=WSVg3BF2.MMO-,dU\_ZRfe0O-:GZdN0):=I6E&,d\,TS:(39,NI&\1KP?T
RVMMc#=dT=5C/e^CHNe&,5:XMV<#dLESC:=ge^MF)FA1O)J0\e,UVSZec:1&.>AU
Sde_T@Q/5(b&B>6dYD>JMa/FcN^7;@-b4ZG_\Z2DESag&Ebc+]]V]==c(QC=[<B7
G,<&3Id,=J\&0/8I,.\OaAfKdWe)UTM?2d:gV3[^#AAf7[^XV^9E6DcU>@@:8/0G
<;-Dc/8XUdL(4g#17bc-HK(I]LLO1LTRR99b.P+C,?e1ZUU4L7Z5I0>,N_6^^P8E
ILC^QX(8MJ)/Y_4=\R/TS:7C+6EH=d8AD:V-G:aP5QU=]?O048a0GVAD48K[MF5:
(RAPXVgTALJY6>FKTTDZO^S:(P@ZSP9C:FMP2VLJCZQ0dOe[,gNMGLGQ721OaQO-
G>D,?YRHcDJLg7&ObRfU#YBK.d1Z=7_QNg-)-IaO48aXJf<g5VB4]eg6T]?g3,HY
KFc,,DPd7[aO_Zf)009SgeS/:Lb++YFD@>-RW?Of>aITKQ2@/1c[0fO5I0_55)N,
ffbH2<Q3\QS,>-AMMG:U,8UYC#?B>CIA5?MF7DK7;P?V6PZ>?-M-57C,TG=?=^(+
;CTBg?RYQ+]2:ffI3B+a?fFM)V@F7,0=b7#W_)e0)gLK4cK6#9NReX,=CK/MG\Rc
ID_gM5NM;R[9aEXXU2g,>;1gCQY\ReP/&XVTOE14ZLRV+HP;:ACIZIVeE]^ZJ-cF
05dgdX_.0Ke^M+M<;T]1)M:5K1J3V.]IB8H2O@1/4B8G-BC?HFd5^[W8(ccQG>P4
[g)UM^,;PLM,eC6-?),4O_.,DDdFDI5X7^.+aC<^?1J(.#=ET40CO,19@[^Y(1[3
LE5@_C4?+Ubf6A^&YW(c.QV]L94[=@2>5IN]g,Y=(-(65O.8MK-Y^KgSDPNgHOcD
_>_JXTO,OB0+P4b/RI53X.Bcdc5W>_M(&R5JG.PRb8J5MP43@\)W&e/c5/^I1B#O
=1fFZ6;X2\7@@PS?V&Ee4(0&gQ&+gY^K^DN,\2L;J9B8fGf631?X0)//MdLT7XaU
^c,7SgSM/Q,7=5QDG<RV6=R3EQI.##.d2P>?(O\I-,@ga1fZeaT4c]PH:fQN,Db1
cF-dBf@30[.<gX\UdGNIZM\U+R9B1EbPb3SB&XgD@0YD,.H1DJDFG6:+2^c@OP[L
O[)W0/7#SM3#H_0f53;.SAeb--MP/>Ma<JTQ^RR9;P1ZR6X,M5,?0=W0DH\TYKT[
8BebcGL-&?TYZ5@25^4&<?K]/44/[eFP4fb=a#\O.84.bfL^e#7X]BM[E25MB83B
(0_G/,082S5R&.\W_05.DJ\f0eW(fMSP#AHaVYLWAGRDPcEH<IE5MFOWTN(_=FS\
cW3SX<N>SDa^JNQaDM^3B)47(YBcgd7QbGOfQ@@2+_e?-)1OF6&Hd5WfNJ(TK26N
FT?(8557/fAA3af<GOJ_522D3;F;RWCQ9WA69e&#a&JCa@+A8d4)3S6+cbHRC-QW
eV3\5_C16<\OS,&#DM/]ZW-a.^W:1(AaN,[Q1<3[=g[1WX5A8e<15TVKB80L/gU=
&-X;8?5fE\(>:.WMbKNF<#JGN+RIZXGg8CMK>7F-K_5dDc-W&=QN<C6/=FUQUA42
;0/6I+EGX]B+=2K5R2\;S9PDBfHXTVgfU.e)g:_4557MdG:0_48T,P2WEP:FL9Nb
=K:S]61U>^2Da.RRd98WKMeb;X=2.EC.b>84EO&^3S\HFGD;\<:21SN8\V3NI[/0
QaAI>NV/@^L8W[XYaL,JD5KMU=H;;9ARKM.;+K71OZ#81:)X+R+NAdHbU5_1W+#=
HAL[=[Pb+.f,F6@B>7c<9#=-_^Ag7JB3YYc/d6^ad,\?[+Q>5Z,-.f7;J/AY)T#Z
N;3-=8MQ#.5:6N+gYL2L[1O2Nc&gNPZTB&#D;BY8;T]92L-G3<.&9Wd06aPW0]>&
3.a9AB,Vf&G];HOcKLXQ,abKS_Dc7<Rd>IG^M[GM,?I11O>=D,^X_JBFRSeT].aF
0Igf+==O\6>_8W22f.T^55Q,&,A[F,##[EE=J)g5),@9_7[6>3:baXdU4#4=Nd9F
\/SeBH2]eWXO3<.f1?]>Y&XU__KVJgJ(e\>T>S\WD0V^H;d(IVX\C(/39\KYA+ZR
RQU5B^4D[<A?a]E#BgURJ;HB=bQ(0^@3+U1TcG^\._4UH)NE^,_(>A5JAT\366_C
e:>B;Dff0&^^J^NE6>C\E5S-/25BAdCE0#76g>B4>(E/Q=FMOSAD[:B=C>1^=HYV
G53HH8gJ1]^a8W0>[[I]dIM@FUV)H\#B0<cFd(7DM(R9=&HdOgU-E9K4@M,?/^Kg
O(BU=76@<FR<DggT,9>;)W(JA3c&3#fY^R5]FT7R=ZLC<a_O5\L/Z:&)GXTd\9A+
(a&L1b4a[?)&S5);KP.;gNGGe[H16?VMDIGF3?L<Q)XD1N-Qb81CR(f.WF=C^0F<
[/bc@G(7((BNd8SHP2&]@g[M6;?&+U/,[SK0PF?fQIM]f968_.P=XO#?E48XRQ#>
?)0YCEE/7c,GNTQ(dL)-gQ;;:S4X:g,EVRCB&ZN1d:CD[V)NK^&XJ:K)+PJ>@HE6
P7<PC3\W5@f4F:MJ@1T&ZO0#>EIJH0\HEU(9+XacWQ>G+G:G9&c5C+N21VAP\eRa
U),=>d2)EV>SE,Ngf>YKAUBMDdZ^Ka^;+QTZZ&6W>F&4&G)&1f1.@V20?(\9+#;T
8EA6?DNV^S7?/HJBNE0/MGR+(U);f4#5df5XWH/,dSL0GU8C^4VYS&VE.DUGb]bA
VeFW=I.D<Q==>#2P?<7BA2a62V1T<CW?#DSM5RM^4LL(Y7ZLYadTGEB@6PZBRDJ/
Mf]RM86ff@O[F?AP>#<KWb0ZBGD+?<#_(72<gC=c,)2DVJfG2ZL-6V@PAV)B0DbD
TE(1O3,XHV,+;?,0^^9g@BCI:)?ePAJ>R)[E9G]RL>H_MWX)LNADRA8c:\.U4.>1
E1g215F8.I1g_KTDg\\SKHX-9GGd(R8802L3V#G-e)V@16T<Q\a@=5D9MgF\C7#R
FFG6.c:?Yg:+f:4?&ILSGET[C=MDPB/,C&R/cfe3&ZSFg4a\RU1]DI:(\<b#NY3Q
)Fa?DC9F20b3>\XSL-//WT@K2<cB:C3L7#Y4=G(PM1KTAZG_GFgEaQ#QKd5YCB:C
c)U[I,EBF8+3.Q0RQB_0L0G-[cWgY,O:0FA+>)gP,a:>BJ-CB\^Q6SK=ePK>]\dH
_WUB>8<Kc5d7AR_c_O6@=d_=.<^b<4HKLA@L?VD9G?AJ5I-?7-:H;DTb7FfG[?Nd
FJ,b[OBM(fW>YL,GK\T5fOG]U8^X1=6GMJg8SBM&+]7NDYUYR7W2g?fE@[H_cLcf
BMT1R0IHIa2OJT#Df_Qc8aS0>:,+(GHWU1Y?23&U[W2EQO6?YZI3]B[GZF0S<@fV
?E#eLVM+;3L8\X/g__W#(6;4ddaZ2YN0(F7,:45<J,N8?7=/LE2=9b;3>++ML9?V
/=O<O6X:-b(/b:CXJ-,g,.<>T0:[X.PB6L+[&TQJ,95)9R6FQXZ3f1G93BG7]7I0
@aa\Te4cU>N(_aNI1L(RWE_PRFW19eZ\2GHN7/a+]@[9UfH\5G.^1[PX<gaH@Y\T
4Z+6YQbL_9=@1.Q8=bY?b+U:\:#A(.MNf2LC&+6XD0]e-ZBdgWeN6b13ceVPgZR=
W^CR3)6/:d]I3X2f<HZS.4@P;W@fT1FXU/TH\MWX,Sb(4MI>9C(#7Qd16:Q,OfR-
:OB;Y4gQ37a[e5aF3.IffY(J41B@HVd2RYC+Y>U8(Q.PU?HEJAd_K\ZPB,VJ:T09
\Z]/.TIYT4La0735+f0\]UWWg=TZP0>b]J)(X-ZU5@J4^4>G)^?0V(fdgWFT?IPP
;X5G-2K&^aN2BT]TM=ac]0/[D17BQ]J1fVFV&>a&MHe?N=<fS_W3S+_JIE8Z75>=
IF5LXRR(UfeeNff[CMPF<91Y,V7@=:<KJ258?EQ@0/2/QG+M=;eV=/.D2,GTX^.4
9G7H(CSPfbBM?SQR2&E@J\Fd=a]Fc<d[ge02\:^-L):8E-N+?3)5\a[_(X)WJM=H
e5@Meab_-M&0faMJM9GML9(>:.f:[HP3I(Z,(_<\4.9DZaZO]f+57QMF9HCWDaH,
f/F+&=Za8C/O,1\/-?\aEK@DDEF09[Y6[(].Be&:S#-YC>4J?+@Z+Z^P4J[cK7DX
S8#N.&#0.-GL^CZeg6+XUW7\_Fc?&L.K.f<OR-1U,aQ)J,>f0F#L\:X(GZ+UM+:+
F>U8Q+O?)ceaUYde_T3Q_;RA2\YN>-+EE2CBM^]5XLO@G_8\Z/#>^cD_a0Jd+]0\
B6JEg/e>1HTP]4N0?_+X7A?.cY:f^BNV^:_H,?-C_]>LMQO@V-Z(^^@>_QV.X22>
O9aSZ98L^0N[R[Ef]RL=MPF,e-7B&f=Of#c/V:_@.NCB3(F+eFB&GO[O66L6G+I=
Pc;X@O^X+f+0IW0_c+4/0^UG?8I,N./&Dd/0^DLMaTc6N]eLCcZ:)5S=7Hg5IVH7
G5(YDVMYB^LJ^C@R>#,CC5JJ=;C)XdQgdH2d-:;K:>bR:KDKB7^>Kb;/6e((V)M1
&J&a(L=)OX5SSeMG0;T1W<,d=C#[Y):GC(9--c,G9CL_2a4f/&A;DU@A:<:4Af5^
1<EgRF^9N#O4)?K;g&TBJE#W&Y44?9AF=0BR6;]UYe?^.E#1?\))ND=a1D;E[4/T
<(9g_9Zd6IC(&.XV4SQ4V&G)8<X?Ydc0P/d,2[_/\YM_C[[@ed@JD6+>Q\>@J.O;
//24.G3X>ICRHZ&W4:#Z&=)KX]IPg62VD?__#R,(Y11,+?A/R8c4XA&:7OUHKaZ0
C=gFa5I&_SGfLP>]HQF=?/B@,eFP-L,g+Sf(H296[b6]>b]WeecBB0f+0@G#g=^:
,UbGWC:9]^WE;IK_TS;IC1d@#.,b?JLO+Y&P^0\\-/-07;5L/HQLUde7;,L5Q+\]
Vg/YR_I:73^2BN+5&#T:#-5K+)9+N:PM7.2+2K-Z=L5=Vfg0eNOW1I=d&-LcR+Ie
f)9Zg_[F?Ba/d[T29+U9LT@T1TTf>52GVL3&fc7#>G^++6?H-fg][Pe#aK8KQef<
NFPW>N--06S3g56.(?>QS+D9RI+)?8FN]TB5b_QbFL?),5RI7EffM(5+H:gG7=.C
C5B]fTQ)?,^NgC618<^O5O-O#>Ld@(S::9,S:&+2R_>IW^6SHb7K\<7SFeQC(BNL
,BEQI;Da9IfPWAgZGg>FJQ.HL]]3((O57S_BA&<R&\8?M)c,<cB?DJ^5>_)[ZA^#
:&,6>7cHINGTdfW/N6fE]ga[QRJM)6K?>BYP)cCLE.\S6-YB?NM@WIc0S&M^+VMN
d02=BV>FREEM@W,:NM5N&H7].<4#>ZXf:[LE[@JRKI3IW]HO)0<?f4PG+@/4Y2UU
>:#66A/WV3H;9D(+<e6+<W<PaYN^AM/YWWP_496#0-]?#BHF_>Q0CO06<?VH3FI]
0M5\SHUg7>+W5Pg.5KPa#S@AUSK.ZRG^1?3-RFWK[;Ab6bYa7V(G.,dG,Dc7;b)e
LD,DYKOMP@)]C9-YeND-6UK[Je8,NZSSX=)GQ\,^_?K4F2MIF/fcA)bOZ9]Z9-7^
]J]EUHUX^2,^<4-))4+:RA7O;0#eeM&=&K^=@.Q>196RESZF<#c[UXQ[.0^3-ZMO
&S8BVddP4409a<)-\-TE?V<#82ePIF.8c\-M?eDfM_bDVAeIcI#,fN_gL):<^;#\
_?3CYGB,E8R-B#L#6_2\MIgL/[0@C[3L(OHWY&6<-BVaD6A:?J?<8SE=<R8WGa^f
Va(SJ:]:4#4A9T,=ga&UL&]f\_KDBWTM?-9[(3AB0;:6a:XWU1-(WC1Z=6g23Q\>
2M2aTH(I]_I6<9P>B]VWa)\_A<17Y:HQXR=_eQb@Vf[\5DX)QW_a0.fgIESMA3e:
HW-cbgGXPCA]4=0WE3]Re.CG.J2J3PB?.BW9]C607F01OHJH_YC:7GYCa_X-;fb_
+T<WaYRULC=a)UG8.0<\Wd[T3OR&)@?D<T;_2@gb_]]K&ZDY3P:a;a<0LGG^H62Y
A:N+X4>W:B:_FY-fc3H7T7AE7d[5:f+35W\g2b]4c,0RaOgCHe\HPWIM^[SK=RZ>
0dLAaDfDE86P92_Eg:-R?P5Pc+XM/,e^]V]PW#J]<BEVIF3gB>.GP.fP#Ud.UO@&
\]TVII?d9Cc=7[1\&fF^B89A=82c=?Gd=6F\eY0RP9X/^T6O.E;fBBU(:K/dT:-?
=2AHKC-7ZUg>WJ+10.GR+Z5#.-W,2\eRQ,#V:3#/Z\8#@=)E[P1J-F7d3JGH<C[[
>Z;/XVF8@Ma-6\M?d[]</f];Z4H<H0dc(+^O\Fad-VH1e8+,7Y=SD=(e>-@D(2fJ
36GAa-8WgZ804;>3#;^+>Z=?YU;@D\5WN63+Kdc:R]6P@,D;KeIEQ&>L#998)[5?
841=>:8(5e2#EOPOMdU.9:gLT9KRbHR2\TZ1>\<[5->J:c7)OB1BU;1e/Md7@6VY
/9e2@=)g:+H;]S0^OU<19SQLBE^[-=IJQS,C:1Z]N\(\F\PdA:Q:\IOBWTH?K./-
a>PaSC][S,K_7<[@4:H6?7CAB#0VBV1^eUe+HCYD&:.>R-ZJ2:J0gcG\3^WMf0[Y
)ADdXL@:P4K3?;>dga8&6MY7]^3O+8S<YPXZB?;P-;,d=:?@G4GP>3YX75-4U4(;
&H25XN26^AX].O&fTD6LSW0BZFLdL^a8KI]dPAfR27K/c^.(5JO>,6Z:2P[C29?1
\UA--3WYcL7&e4JKW/U8Y^gA9#^-ZC-KTOA(NSG;fEDL8cH_R9T85,-X,41,cCUf
aZQcQ]B-F=gD-.R:#MOB-XaZ88V5B1a\AQaX)^N?0Y#S#Vf87XU\#T:6NaA7<,4,
gCDM26SS2c:P)LV#548a5[HbDE4HL-_SGDHQSV2HT)ee_/)&M3OUK]-2?1f9g.f&
Q2(+3:T_,CM(HA(-?K5.TQ6Da>9dCP3+/4[&aIQEQ<>WZ)4=&XX9JU0#)g&g\f:I
WFB38P^UL3=c2fGHHbH9F4(U6@L)4bV\-W>HUCVX;62O?bX16?Q(g]APCZ1@:721
4e6ASW#QWZN;LG?MSH#<.Y+:dIJ]/WT)-Qd4P1/-#M&gb,Id1GS0+TPIg[BGP1Pg
^)bb/6[;&+5;6]&NQgg=OH#ZfSA/b7#T-UXC^a&K:U#D=27WfSWNMgXVEHf8WR[9
IUf_Vc3G_a/<03&\-)aOc#)_0QYS9eQa18bG=6UJ\<N1]W4-bVb06<;Xf:X/1?bP
+b5W;6TU:^c;B,QV9,VXR@GD;Y7FMQJ<]0TX^/_/0NGa6N3MTD\OZcSWb<R]+e+N
^QB6LMR9>H2D<_C.D:e:#VHP2RaQ:TPD7c]D->Jc;Q^4QE^+ceUd+N:FTd#VISND
f7HaQ&M6>b@UL(VVSNN,GIJ>MU)K4dLG#_JeF,c#+;8S9]2G#86g\6\O&0=[0@[/
WM@McL?Y<^;I(U95+SXG&bY);WMB:Eg9gD#,271a=+E@2XW0.IGAC@@9VfbF<TI0
N\J?[WJdaVF#F9I7C[7V]G8<PO8&3Vf\3R@gW/cM)cK>DSU7MS&Ab0b8KZ,5NCQ)
AX:DK&RE>]T()86B^OSD.f_?03MLX3EZ@ELSUU>fF5@61UZ^+dQG6bf2KA#&].bf
1CE:fVEX(H/8Nf.ATFN5/+@^1.ggWPfSB3L1)TF4,8>Mg:@F>Ic@@L(Y>E7\\.^e
?fcRY?<OSA,PSIP:JaRA/RT[dKC\3cX=_C8E81aEe0Q?1O-2&0KbP#ddGX;F^b=[
9RW5+F=^1=S&P/^5fQ_@8F5R+R[-P;e\AbF_I,,^[dSY6=&@7Ve-c+b2CbVR.[d@
W4Z&Rf/A^G?baO3):If77C@#^T[Y\([:Y-ELF8#PEfZRRL+3;]1[N+>N1GC2D^WU
EXOa.CgGL@[8WC@b+=aTc(RG]>E>9eDFASW4BCRfe&1KQ-ZCFdTQC4.0V99XHO7O
7U.eF7\FdVV6d4T/[9Me4f&gW8Bb;I]_fdP8Cd^;C.g,A7GcZ9&Z\50HRT>(C+^0
(N@_Vg3W3MEF5F7R<&NEU);d_G]<I:-I(O:-UQTC1S6&<EGeC.AD-EL3d4UgFTV8
Ze-I)^\I=e\V\eYI8)#<.J/\H/>0-(]2Z-.J;JA7XO6@cZHD2(A)UG(@=PE@B=\;
PEa;:0gV]-,b_1.99K4^L.RM]XC/GOYRSE[HB;K;Uc+SR2Qd,02a@.[XIS?Cg2?F
CM>:2,/-3_-DOOY?VE5g9+dE:E\TKYRO77Z(O:D#255Gg8b:GGMK:OA36]CZ4fQ1
A0,WEcgWN#_/UZ=U+Wc]MG=ARDe,XZ2N9Z/gZFBY-9&M0>]037G)Ld<=@L?BH^&/
0bDF4;DZI:Bd3F-?8)&YV(WR<Q\8JP#LT(L,Sg\=1L4&5UgU/G@IU6B>e#:-f1<2
P?B:NG;caWS_8>\=6#ceO-YM4LEZW<-7c(VOIcO(\II@g\C@110)DN);+[[?>TET
6HR.L,C,I2VgT0#M<B<2LE(gVDJ>(:9M1ZC,V(,VR<[FM/Bg(Q&bUH^PTPdegd4f
T=\=_K#.ZL=M9HSC^7:7Q]d016fOBDW>(cc0b:D(/]125c_ENB96;U)e>ZM/MTbA
@BJR&)2=IgSZ]I75gOGSB.-@Z(8#5aJ8d=a5f;R@2;c,eT:I48B#@<2CA3@D(_WJ
3B\V-/8e8KFgUcA:7+J?9^L/CJeZ^7XO;D-[?eMB(e5ZL33WU_RAYA#(#OgZEDEb
6+OU(2C)0=M/4S-e6L6+@V.LD=:O9C3cg@31a+&0WHGR6EWZ:E6<K<M<adV7R;0^
5;GcU)F;15:fBd5>F.0>DV87c8L/:MV#&HLgOGU:cEHd?\c?8.42D@gP>-8+_^bY
=IZXGE[0^QSK\\[.Z:-9&D@Q/BX+@):@VZPJ/3N0e@6,1)CYd8fDD:V58-H/1>8[
WdJa\?@5@ADe=YM=;@I_LWWLa/]<6,/+?1+U2(8VC5J^@(B6-(P(I_J+;]OJYE9^
V<_QbLWS+.3Bf#ZD&bG(,_K^&cQU/8,Pa^U<E>RDCM0N:=;N]&34K8_bXP=YYe1.
>T[OP[<(LTBRT.)V+8,\=K7:fWcI-_C7d,gCL-9CKSZ^@:T2C?[a&ZRXRE=0^AdZ
OD74FOF0&c;KA[B6DR@.1\I&D>F6.E]dBA;#W[F:49+A/?:;8B/</?eR;EWQPfCL
,AC6A6OT,^J8I?9<S+/[KLU8LXZ]d=>WEe_[.NfBFFHBFX8TCOf.TVZ7X+dQ9Q04
^PHcG/</Ne&L=Z^>Jgc@)]g3IOY5K/?(VXG)b[-BeJ<TDME8HZPJE[=_,44)K8KI
0cA9[[U^&K47M44,Dg31,@RDP,2+8\U\Jd+C4OZ,J7.79_?dM=4fSSIE<Mf[PH7)
D_K_;H3\OTDdS(8\L;NTKFe^Rd8D9P&\<J=dB)W0QW>HObY6,E.BWC.X&]b[3X_-
O5SNfZY2RUXab#NC7T@[,IHL/dM33WXa8R?4NNO_0Z^:QJg>7;-,Q<]9TbSHM[+f
#:4c&I<KA0>Tf=6]NPNQ08YFg>Z61:.XgA\0A=g;:2DH,GO(T4KP6_;FKLgaQSIf
]&DKb4X7NU4P\H6F=<J32(.OV0844R:-3<7U:FKbB3ReY^H(M&N4GJP&)=?0^M+7
>..-^X18WdZL-H0V(dNPdS].-.9;3,//=JCHL^G#=P-RJSDX]W0\.2gWf5RW[:YV
Gb511935H&_]FXe>MF@1+?e:2H?U>b5?<86Mbd_DgTU.BNPO?@G1:ZAB^7&(/.\d
8c-LLPN#]8A,_S#@aBTAO_5?g52E(P3@LNEVN7:3UV8/HK;L()R(3>,:6g^P+7QY
S2Z/.)Qb+gY/?6\3.3+F6.1.^R>(\O7O[9d],(#X4YVMPS&.D9=c,I0=efV=g3>^
ZbFc+\:#EH@G^<19+TFA&>ZO/MWK;dBgM6abU<dQ6e\&R147Xee+41Q2+XBH_?D8
0VG[JV?D;gF-;1>1,KK1(8E.9OUSO4D3A]7ASGX7G?5]M1_BJ(+D<_QKV?<PDGTE
E(6J^_N6>3Y93YgU?d2g@B0+B/PV>9LZRY-A-?&KX7GIM\)3Y2Ec#YF0OXg29H2J
BWAEb6c)8L9TJN]O35QNPMN:1,E)(e\HI/&5@7N0F5U&/M]+&b#4Z\T)\#&dc-C6
.ERHSXeaX\g>87\+M+@8J&_RR@.^,.3bB]]MQ.;>E@He]Q<4aT54]WMLfTHX3S/1
Z9[dIB_3/GF8KDVTQ<E+.(@K\TXP(R_]:XW,65a>&b\O3PB.);<0GA:ANDU<7(W,
QZLK\@I<)D7b?@J@Tg.]c,+^]@U#M06FZO?@+=.VQHaY2A(YD;BEac,gAM6@)>KN
+caWI,P=YT&?D/94(H2[0IMF:A&+\8Y:C7aG;@>:7&RJb34,D@La@.DQ@&\U6G=c
B:N,fJYeP>M+&1N=e9R^d^F#eI>AO3JS2.#+a6Z0(N7f;N=F#Q1K^AE:Q^1ARJE,
UU,fO\?_SRX_?;L<M9JYQ9XYOZ;UEBfUCcBFVb#B:I9W5]2Ic>[SW?eN8XX24faF
_^VX/^#Bd2b#cGX,NKfWDd)D:M?0N,6OYVV]OEF,1(^=Q307BVgK8_TDbUGc.:8\
]H](FA1ZN0+KL2VI7&_(BQdDJK4/X4b,TKe=YAN4@P8;;5JdXa)8]d1]-JZ2QQ+M
MQDER62)aW#QQG+--(F>1ggeGMO.O&MRE=fZR#O1aD,1.0M_G^-d?8f_AE.9DQ.J
D1HD<F8>5#WTJ/gWa[KPCd1f._Od0M^+4<;+A&B4fTcUY)[g(dLQY(UPT_JT]^8B
.^=ac5/2RGGZ]/,#[-94HPZBP=;<K@):dSZ0EbFfYG+BYYG_+c)WT+OR#bfOD&FV
^Cb_DL3b?#KA,N6b57Q[]1&3<ZD[EU\P/^PW0e>ggX(_bI#-=HG@;Ub7:D:U7(c1
UZ6KQ859Ma_5MW6,-#6><f<304gHEG])XCFS1,.QKLSU1/YDL+U?gN+aKN#c5+?c
c/g;.+)=IN3<C>C:QUZ^#[)]aU9FP:OK3Ic,30.bcaSBEW3/5Y;e)OJDH\]&,7e1
fYAN=[gZeB0J_VNKSPEYRLSf\<C5)CA:7NVG&&\:,[b;.SFJfOY<Wa^RbAJT7TeZ
7#-&ZZ7E5O<E)4_\9X6C4X1\J,1gJ.(E4S260X1E0VOO.:JR;\#&J42^0@V)W/HA
5gZHVFVOQ=BJOa+;GM-Z__:e6[[/b^GT@30cf69_gERV)ZU28_02QH6_Y^8(b>fF
@00Lc4/2/Z0XeDZO]RX2<bZQM5e=aA>7E3)HW2PFO(^CDbYK#=\?Uc4ZX<W&80e=
LZbG1O@SU<6\W2cYYgP)P3-GE,.6TZ7;U69(XQ[fb[LfSeD\,&^]YM3aS3d4+X;Z
6<e])>6Q466LO.@J6N5<BcW19a\@C;bf6NQ23;C\7P5T:5(:?0c?dJ)66R&06f-+
^Q2&5K\aFD&G]LBB24YgUCW<If_bHIa9HG6?9OP+V+>S__bUCMIDE+cegA]+bL=)
+GAGc#H#.QKPdZJ1A[Q\b;L/7@<L.6=OB9-NRaSd-3YQ@,a=8,1R(1:84@8SO+Cd
7F?X-2X=\-&@d^/F#CDX:#7SI@RfWXWHVP1O411ZOg,8XgV9EPZM+Z7JP?XYB-&&
EV^JEVS/bHeR_OTa6RXHU_YBgYA@Sca:.X8227D^)L?3/[=L<cV3SF(FI=>_(=70
]K,L/XEDW1#MOe][TcTC5=g8,?d=a0dLaVA]0\Y3_4>)-APWJ,)^G8c?X2P,<M^Q
GT(5=P+N.XS<Y/_P,cG2+[^&RV<2+4,,3Z<&=S<U<-L#5I<\5L;=5Z>;;cU0,d_-
)V)M4RU?&ARL@A2f^LR?Q8=&fSX6Sa16F:Y85=fHc.0cKGgcd?TdJfG,/X;-7QXH
7LdPQ#gR&26U+a1MN-:9_[DQ&aEDcIEO&G:8TDUJ6&N])HS^;,OXbgFT+B1P],B;
)H-^a(GSR([f1Sa8UL5BRXI/PR,KI(6/(66AT3-9K?4751U[.7K/:JTKg-#4-fTT
H-f7N89,&J9/B.H>6?=D1:B8[7@PaD1,e?F-Z:#T:aTce^-OZJ8JB)FX]4P#7M7.
Gf;GVF&fL9G5e#e5,\;0:U[XJ@33S/F?Y)0]DF2>M<W-dGN(OcJ6BEE1BSZ;@(Y9
;8WDc^a_W77(=L@+GcAY\SPAb-XJE+QMJG-QT@:&@OZ7D77g(B>LR^ILeL_,+S?R
F2Y2Q0Je_2EaRB,5Y+f;I&-R1Y?1.T;<6&>U57RSC2^]6)?(IU5:=JQ(@F1TeJV<
W7E=C?MHg-3d,3@\6eaf8NTETab\Y:@N5\1\X5)ZbB6@;@cE3f4c_LA(ag9NE7]<
1+aO0D=L(5YB.[V:T6:c>2Z9HeZ4eV66J2K,=UB1N_:E?Q3ISKDe4@BRQA\B/cM\
f0)]OMDIB.0^&gYRW+BTaM]08AQRF,M&\S:Ifc>\&TBSdZZB9SaARd=@RP[<4aBd
JD:_c.a_f&7gZ:;(+?(NR\+a.a,bB_)Gg?/9e=QIVaUI;7P/cDWV<VCH[XR>HbN,
6Z#d84#0?2J&^+7cJ0U),D/CBW>Y3C\e@XO]]cR#E:1cE#8fFfbTY[&&5R=0]bAA
>M;.P]P1aFcM]XG9.Ud(;JfOdO9;&9.gb@dT+Z0<XC8JBcY=-\(20?QY^+bR-E[9
K23+7KZg[fLMICZ;EV2_V\;fT-UE\XO-6)9ZU0MA:04G/4P#?/&dR]D)aPQKT35H
C>B/?Tf-X3+#-1IU&-[Me.<=RSHQ4_ad9f0:GHL^//V+VFP<6AJNRG5H]X#(MKU]
LQ\4.L[KOF7)NY^)SC6U.?AJJLc73M61BHM2?Q4MKbdQ;@/)I7-TF2MXP3C&1O6/
M9+;+P0C^?@fZDcP[P?&UM82NM>.@VS,F+35\#_V+:8aB_0eXDVDc,RG-8RT87JK
g\);SDFHN#J,5M=dO75^_\dCK/aJMOJ_H;8Z&eJNGUGB#&5)0GPI[Z,TdT9,eR?.
LG[7MXWP#\fU#&&@U1Z?XVE.;eWC_fH]#3I2S(fN_+\LH1FQO:A4egB=Jc:db/V9
ab(CAf>0VR9dWCZ(ZM#4W.LJMD\&[Q0RDfON0WA-<KQC,\#;aXQJ&L:N5aOGCc1e
FF/NWePH+_C5VLgcFSY)4-FW_G]H_],>PafL@LVd-^=\[AU9#W]db8ZMW[T/AWGN
C])C6:&B<cF7/aKE);)W5UBO=IAZ^H;-0W7A<f]#\S7AQGLbH^-Q@Wc3(L@dJAb\
ecg0>+H(.P^0@_/JNaUPXI>6)AH1[ca6UKQW]BM;M[H#Fd@RWE.C>X=gBF=\CeG<
D(YQFGaGK,^AW:g+UbJ_VH581gX?(0>d0.@,A(PAFNFAfOD63)OV@bT.e;BC<,F<
7.:OSgR5/7E0OO<c:1AD94ILHG-LcWd5dDXH=>fb_4<DHDSJH)WJbeGF^XPL0/WD
LaGBDD1_c\6/)FI;EdYbS;((EMP_dZOb3XLS^;YLA1>QC5=[Y9a]dD7GE[^K3,QB
P]Q\E8QZM[#VG#:bELA\gUVHKe;Z7>WQGZCX_eHWTO)F2:&f&I27GJH^5NfEd/g>
B]AQ8\?Za6_&ReX7^D;GcdD&:3\=<&VGfP1904Y>FAL=Y(S=LQCb>UQBYc=Mg3Q]
UdM/Dd>OU<8@XN,OZ@2P]WIb,,>=^P7(/#GN-12g@)Qg2,+cS3dC+.G^04ZAQ+&-
E08aU:,YY4F\5\e@YXcf^6VPGfYY4D64#-b,&)Vd:9Y_L)TbY8ecHN^aQH0JM_^[
];EWg,F@5a)/;)WV/4HC:F>JFc&25+1[5Y2?(HO<=IcHNV+G@PRT8ffD5_NEB2OV
L72>=YCYbYD0M3CWOeM@MH,)M8NSE@fWDc/#XJSa;9M,b52&?E.@M?<Qa>9c6bPf
Sc@g=-^]@N-\_e@OG<?W27)b34cH46I/,W0,8+N^:B1e9CBXKX(#LTVcI4aY@6aI
EG_2(EF_@c/(X7&6fC<e-V)OCbH;PE5=?20[>WFL,K>9S^449S2-eWO/7e2#_:\a
=K70]+^Z+/_1R69<UT,\X0>0+f3SYc_bG[@<1.\4926WFNX>HQe/(KV^YI+CED2K
Hc+K-;S0E-Sc>+2Oe1CM3aM8UI\[c&]BHNR&?^1eXW=?P\_,S_G.Y[L:=Q#5DK;+
O(?,:1E-E,N18WIH7YPEG,GN+K>(2Q?=KF[?_ZDG9MYb_S]IHea+20A7F6UQB>@B
c\Q.1]BULJR(aEOPFb5bfbCOBVP:0R-YYS4@@1AcZRH\AHG-M.D1L_CQ]YA9cGHO
BE<6CGC9.RZ9P:JaN)4c<@9Q\>V::d[O,;OEF([Y]SGfG</aUbBR58+7;:]0L8]Q
A+,&#[fSU59YO\_/)+c[0fONdJ<aB8U0+9<df[R,/GQJ[2P2^_G&POGf1[aEAYRN
<@G?>Yg);agAQ_IDfWc&)F]C&Tg37QW<U?eacBU#f#Z[\F6^1B)H)),AIK_We<H=
eTP5]&HV(6]>Kd7>#P:4TP+Y[,L7VJY+\+0bTg&J9A;C,7C(S;MFL::5:1BIgbL0
PE&:56D.9R1W\/C@FYd+Eg6ZREU)H,#@1We&EgHFeAfTMNRa_.E2/:57&_+7^2W4
C-8-#K:>FV>Be&L0>1bgSV)2\=>WR0gb>XIR;C3:ZF(6NMKM0_@bb6DX2EV,dYX-
]75f^a<RY]E+eL]fg-9fSPQ0\@B;#?A;O;,\+JLWb@Q5K>C28ZP@WYV[=b[CU;d=
.57)DL-QcIY&N70_9M[aWH\FbaG(HcbP]]3..dI,fEK99)?5::6VP34A2,Md_H_F
2?FgSdWW.aI8:gaB/7g1VONNW](eDC0&Q<Q6FLLb28G;bc4:470X9GbWEF))13J(
_RSXG>fJ42OgRb=>2C1I1fK];DAc^+VN_TK@K4Pe;45J+N.+X_6E(>]H1HJ>64fE
^(:e5.3@F<D=I@W<+\&\GI^#=50VOY+eagFTeBUB&KXL=?M_XKK:GYSFOU4ZUeWN
e[KN>Z>TO.R/Ta]G2?GI[],V]-.dU?5A-Nc3-&KH/^d:UBUWbOHM<PRU7Q4d.N4U
&<[:86<6VgKAEdPH::0-A&#Z&QU>ebP,Q)BDE9T[+/80g,e>H@/810LBG>F78@dA
4&DGO9^g(eF#b1((dFMBLLf5e2U)4;J]E>8EY^F:d^QW.\IUKdFaa5=>XeM\W6cc
?=S0bg#eg,@Z0<#Z;e@D\]dP.P=LMPOQD;bW<Rb#,\geHTJ9&0ZL:.HAOWc:[gf3
?&3\O^[P@YCDMIO,cHd8PG>M;E5B>S#6MBNeS75fb\ANA+>@aIg.QWHba.DYMWDD
,c\SGM2(/9:;;F3RI0I.BRMZM+QQ]@bRR.Z/AT<G\4JORPQ/e@SBKUP\S+26GIM:
Ca&MO#1E=;CT<X]T<[7F?W9NPCTL3Z[/(GQEC5G\G?)\<L)Y#ILNM;A)O<XZN\.1
\/ZJHF^X;T[FP(Q8IeDL^UB)FZ_K9OF5C62O8G.+7M@&:Sa4fT:NV&a<R&10C;M[
+=WBGV(,W]6210\+Ff8?]\ALEA.;5-2K7^TS>Q8W0CN.c.)JTb9K,[fXF3ONC^RG
+N#ED=P+,7=)<0f3(H-94gHL;WC?4P(SeU&(?MRUI=U1@D8^ATITGYIVPaUAMfK^
Y\H,28CF:E@M74fW5G3]9TC>f^O8J)_;RPd)MCfRAZG.E-3JT=Q1_&I9:0f-2HIN
cNA1M/Cb8<#:>M:E?SW+#+-/JUc]DBIfa;dag<:GA17B78(RNE817)(cR915E:a1
Z/^6TENeU1+8A,)Gc<ZIRd:bV/>1WRCOG@&>F&XReP>G@=[DPXJ08HMMHad0MV.2
4T7KL2f_#@+a+;,c57<:5RXNYY3=&R?9W9^XCBfE.OZTA4XTQT9F9F_WTX@@LR2<
JT2MSVB23]CNAWW-MOH5N16>[/GQ_O#LGG(:[/A7@f4;IFg-CDJfAG;bX3NS5Kc1
GZ[G)YR7)&K0QOW<5ALgAC@DEbNERd0;=UT-9LR(6U:?f5.37],b##<05JW=RVf)
M:#43<P\Kf72E94VbCK@<SJX(]HF87<H]9G+NVN42ZLU>^76^OLCFbcW=AH=)+-Y
,5F<>95cCbX3d7[FPa13W@S3=@/B3KB27K=HWK]gebc-&I0=-MJNGU4[fYbKV9)8
;^HXHDP\PDgXRbC0/U^PB@TYgDEN#F=@C?Ed(D=84+YRDPYaH[3cX9f=<7/5E@7E
:]K49:gaER:Gd3CO:2eA3E_SEJ@/O&e8C8@fQB&G45D(J[CWa4XHAfQ;=X5P/SZ7
SeTIK&[d\;O@c\d8R+C,]6KMYTPf[J:OXT/MW]\A)dL,BR-T_Dfb97I4JCaTQe>D
(06C>=FR:U0(>fD3MSF6>Y_;WI[Ig3K_.g/bdU)bG<a[4[AgG^</_cF-9g6QeZ-.
OXB3J_HAPg17,V@7-XI7W^gI5H#Y.TK>8YQLGKMZL(:VS\H-0K=[F\5C.BW@8aX<
NL;@)_8d5@F>R/?]#Lf[F8b.4T.\X=[=#+67B3Z#EIQRa:-))gCL3Gb/<KCO_Vf8
H[4MIU<U<]H5QW:-:&gM)V<(We;cA6^8G1RJ8c--R;BXI>IaV-fdeUIZT(+7)e[7
760>fJ2OLcB/NVdb&C(\WfT_S,RT(fgAC=BcA(Tee-f@gIa,5L,R<.=dI3#(B^R=
-LB-KH(4L<KW&aY^9H&]WBDJ]]/7^f<R+JIT>>EP.O0Q@F1Db(F),=X8^T;g+Z>L
Q5\+a[S\JAc^BE>JE9O@O5ORc@Ug3&+<C(2S.HV]Y\S96;3KBPSLD#GB+bB,XQO7
<+6K#d^)-)@.,K.ET@C+#>LE4/gPU=8(G?9E2M68,-/(U?_I<e5J+f-EY05L@;F7
\Z#N;bdJ1C3)[Ya,.=eGVT,=Lc(V4^T;;FE2[U6c[]gUMSH-^1+G;;QVP?/W5X>E
>=<EH\+93?N=XP=8H,B9U,^81EVMU;.61=&4bD(9d_IJ@P?5;>-4RJ.dc8NM[R=O
9;LZ)V@@S<M.AK61X5AO:V7,cE-.(ZfUW3]5KJ^WfT@DB;a;6[(:eRFZ^_H5<<W&
/[[,b[\U>1+T_fJ8T_L^C=#JLHZ1b0(cDOWXO[4HO[>.6+=25Ng(8&=:AXf2TcFQ
dR-\A+R@&GaNMZT:He7AT>&F12/>=/X,2>faW>NT2Z2^_O&0\:c08R;[OB[5KM^B
RE)N5f0L60XLf)P]OZ>6Y5P#Uf05:MQda07OM/<-8UQQGX8,#LV25dRc7+P3O:I5
O=ZG(2W]AP.FAAL3IZ6fJ&_(C+>dHKR4Q>eHS<M0<\&WJ=S-T=\bP?/1GLH?85Pc
0(Y]dU/ZTZ;:K3<?BKT3J?TYBH0RHaecWgJEa4,9^#4>]\>eWe4IQaC=A(&a;MWN
/.<^c9]Q=TN7@(.5CDHLRKe#R_?J0XZP.8OM=X&@G.N4W)P/cU^#2W?VCO(<DWWF
/Qcde,<F)F;GGSLCV@WB1CSb3#K^=\I)#,gO\C@f2aYeHNb]=COg96-\:6WWXa=.
L?B&Af6@7^ab/+-G_^0.UAAB6^Y,_E\?8=8;<4D9;.F.IQ\#Ge_,4+KR9f+PGBI+
YH)+P(;EM50.HI?K]@:HD^G+58:8A.a9dNT^c2dL9&dgb8\BG.a8g#E,;4+M)\VJ
[3?O565U^8TC_)dB:gHV>Bb^]KbZF-RbJ;7Ig(bbf?Ob=_?#B4Z;M\&FgSY;/G?(
[(9V=[T:86P4f>KC^fKVfcD2[0RgKSM<N_AFR/?e=[H&e3QV3--7J/<WX]9cf=fH
b-;=WM;H,ee/L)geQM#Y4Ic:?.Z<OX[7gB^g^eTJB9@F:+89@^;b/(.XLO>@#b9f
^C0#,d(6<UL:_fFNaS5]7cS1@Be[Q(9TB]_FB[LQ0I._Y^1T;QOW&23)-(:/:CVO
FC4E[:e0L]N0c\TZKe<g@g7?_Afb#+/MQT-5<I2B@>g325>U>V5HH]H[6YK1g-2<
e;cX3JV9/=a9=:A+ZdNJ\Y#DcCW#LJ_+[R&cD/-@-cJV-ELaY=1ZEVR>X4aK(,U1
)QDUL#e_Q:-XY+099+-Ig;_F#L]b3G;WJ7._a5_4&Q,Nb14+X..Jf1CDTbN@[g,)
:gI:aVQ/UV/[[5H]Lc_U,DX+K630W5f5\_;@#a_&KC)JA;1>ARBbI3/d,)f7W?SG
BVK=9[4R(G]EV=e6K]XVCcK2XEND_CQL?,6dRY)_3F6S5E3MYMe3[M#X^F#Je-0C
9,0M()=A.C9eB#KQ?L\EJNg_A.bQU18e90BD,^@+N(=T8B_DM[?bKW4F3F@O.<.?
_#IH,4&c/@NdN0]HYA69Q0W>2==;RfP#55_N<SRGB3YS-@\R)<MJN]Ie6VUX7eB^
I^T0<[X75^XXYG9K>f7YKESW6B#;H1=eEB2Q+#)fE,:S?.G]]/,#_(7S?GSXA@LX
FV4@>-1JIR,GMEL>4_9MfWZ]0]QK7Dd())YO/23XR]J-U_:<MgD0Ed2_]3(V6VdU
;>2\;-N8@c00f4IQEM/b1O<>O3dGCEW(1#,D\8_Y:S181,OCGV(RI>8c8Q>S0<15
9e_SDYP[]6[)+UEdBE@ASO8cEY-KCe[<1]@4Y-fO(;SX2##M.,A/_D0F=_#?61N.
,ceQ9B204M0VA^b>ZT#\,_.OH>QM2UJ)]5fS:[L&&aH/8S_1P(+O,P((XU\6.WY;
#@(OE=UBgZUELO-c[0,9J/-8S]P_U(CI0AFJaYI)7-]F0_C8;F/GB_Ja8\>N,_3T
>\P-X.Z@cTL-,\a;XUW[YeG<W[Z]JHDUdV=JHBC.1@J.-Dg/F8@VgBZ=0AE+9aU4
3Z7@8&\2S(5F1L8[g4;7e?4903&?_ZdgNU@C-DT_^VgDLIR^2RZ-@/]MRS(K.B]2
83?]^7&5MUg,+FWNT&GGGc\3gT[&<2g)g:Hg@3EMQ_0aQ)FL0:8#:C)55O?b:_]N
dc7Z&.:TV6PG=#4J4B=?fdZ2EGQb)G+YKf1XQY8/HXRAYcaKC/&]N.g65afY4K9=
B+NP>=)\7;(BF,HT[PAe,Y4_Nd?P0b^TC5^0)A]EN=YQQH-@[RMbJL<-eLUZ>LG7
\.c<T\:73XK0=WVR(OQYR5B37OQL6.^VX2V(5SN,3=dDYf=S8<?L7QRGMbH(GdV)
=I7TeV]ga5Je\)<?Y^R-fB/4OOef2LSO5?&8^OTT/C:@J@/K0gH6>Rc_EHN(GZQd
6YC1_0YIJVEX/Z2NY-(P,D/5#YJHccB=X6W474DCH4Z7+B:8-ALO\:5SCDOQ#CQE
U)_#(f_7SJNdA]NLO;_ZCRLd/Y-F>D61CXC&/GWJLSSDfG\L?=:0B155e\Zb/2UC
<c#X@P_D&eCCSG.&_QJJGMcH@IS6D4-WUUcIH+<75aX&Oe-\0.6V;a.QC.7egb<&
D2e,Q7dZ7J)bHXe3;LaGM=0N,@+RC[TEFV)LI?=[^C?b4R3=C,\FNA(.THGEMOg0
,)Z[+Z/d-PD_Y#G<>U[+)Mb4D(W^;6)Id#.(g4_R@CD6HfL\_LLf[-&R;70\cScU
/+;Y=,0FW=CZQFNQX6[ZKSW4^91PEHW/8U&YQMW69L>:A=b+HXYfF:\8MbK(edLT
<ZM28ED^eN9D]APOTT#O,M<LeVU6;EX,CVDc3[TfT>GC=VM?Ob@eV^L\:O3>dDS>
dB<_&4-+SD]EMKHeYSP:MP;0X:DRH<bVJ(,I2P\R]DUO_cORM6aJTR@LN.B7AS^7
PQVA\(ON><JJ4SfR1YcZ95Y,+.-AYTM.(#&YR-S5NSK#Q7FM#_CfSP9baEF)A5L]
;OUbYbf5QfZID:;/bVS5.=LU3OCVVQW\d91A&/@-acVPc7L?CR5#&[K9T,K\Y.E8
eS21?Z5D<(UJg8J>J.5PR=FR6VVB=B1M72A9)8S:2cVSXd#R;3[1_LI7ZW>:8&2)
bL\@ePN4V?cS5_#M@Qc8[G5f0<U]6N51]CX^N,43ZDcLEPO58WN[#Q<6\DJ][D?\
/^@#(\)Ne?T9AM.;.\0>7SbFTUdg?JbI,]YSB6EELTTa>65KUdI#^_IVPf#-L\A2
(U2Q8N(e8DJRZ\EgG(gFH0=^SZE&b0F?VXR5D_XC6J[>-_Ug&Gc]C^B:<#.[\/7-
2,dA3(9V+d71+MEI[2C=LbS8d<g5C03Z(QTbSO)T4Y#71GOC]3aF]-K,EKX8S_cZ
<;^dY>^b>+SL3L/4XC6Y;VQdKfR:L-:7c/=^D^^:KIJC3:>+MAgTJEY@B.c(-YIF
>@;<5YIP^e>EWLS[@_<B6@Y1?Tee+70IY6DQ/K+Yb5]SBF=MdOCUNb(aV;MPb2/B
W_#a+;0bL7(O#EAUTb(0-D&7#)<LEZA1ZfKc3MCNBT<YLAa)g.&C1.Q?2U?Q6\>a
B_>8(_SFW5&N.5ec+FWE8UPLD>,OK42H>@5]?0(.AW#6/_>61.gfW^)aKD,W:dOT
Y8D/;RY6a9A:GE@]4_V@8>gLaW-EbPAIHN_>6\1f-H-B7@=UR&/;;P>.FB^,4:\1
Z;KUHD:9,U:BP6D1M.&Hf0]Ld=+;/,;MGa#[7[Qd:FDH.fS:JWZ)B/Z+1NO>LO)R
6WYO?N?/I=fSA2B[1PKU](&VNU1[6[XZTLAG(SZLUOL[H)Q];<6>MZ-Q8Z^<+R@(
/2FFPaWeLL,RD72c:=Y\R<_@@N@P12CR[#?PSJGL7SO>DP^UPgO_QP6.?#cWDC[g
3^/B1bY4(MYO-LVW=XT@70@YU>O;8;d]F_Z+4P>@Q?<P(6Y_5B,1FS-DgW6c(:M#
YO0AbL?SaKIKa9DO(P,]I8([89?^aY7>OJ7]8A>G:bNIME;<([]D<I]U3Ge.I>9I
9]I(6#W],P<>LA3N7_^-2/1fOVbU?@3/S-Hfa2:Y?-E7L\?KS9bTMR\MFE9-4LMG
^5H[<E><Z6M1.JCBIIHG_O4[+?_54]]JO#WAX6(<VF;_5R7Ge#PXH5Q2[dc@[<B,
,/,]Q,FLJfAODEEF3-KZgW]&fT0eQZP^^_-08Sag5DgBa.S;6U6J0RFYK@D1BFRc
9b.DF#=YKgS7NcLK7/&.0,<YMc+A[eK_dLM+D61X58P/A,Xf^dB^ZS7]bd6\,7LA
[gIUD3/,AG?a;]0@dW=e0I[5+>?3=/b?Q]])QBdGN4G)BOHUeW+Se#[C_MS&8G).
1EUBN]:34Yc#,LGMCM-Z0fGSSGc;FDHNT/4NY[,NR@0Me6A(eZEHS3&#=Bcf5eL.
T_>e:FOTQeCg,DaLTL^]70[T\@g1#Q[>OM1WB0G(1)cb9gI\78SSRT.g).\54#&7
.H^I23E&<gD(WX<@9<HRH=,.6=CdLX:P#_C/30CO;R7A9ENc1>W9fBDIf7&KX]OM
dH.HR(P=^5R1Q8R&#0c\C9I<^fc)]DgW^^JVSN6?MH--aB\Xe5/cg6A7Q:QB)H=O
:S0./JXRK?)0,JF\0X&Q?bL,CFH&&Y_/?H,dg,>)8SH&TY-b#F:HGBG#^]@LL8C_
R2)PZ:4\\+TeUaH(;F8JWWHZcbL\V>@=[PCDK]J\RP/Fe>d1L8\;e@3@GK)1[Mfe
9XbK/TA5e]e>ZP31CSK/Y^XX?fa6>->W78^;NJNV5?HNSb#2:HVH/Ob3JKVNC3\@
#VPgD1+(G3J_WDW^F:6b@R<NKXO,9[+N5b/BU3Sf\3e_?>8VJ8#N,H6,.C5b:.7(
QZQ[>7\RP1;_,1E1,DP0(.T[WN,H7Kf(B[6e^[50>e,AU/;#G)@Y77<XED]:K4\=
^gR(]8XcV77fH^,RV<,QbF5QSA;5HFD^+1Z2MO1a=Oc/GN7N/cF@7YBT)6b#d.+C
DR9JTUF0^#I>)KB:^MH&4>-)T2+(Y&[CZ.4O/H_H;,+cdM2NT3C/CX6?QV?<b]^F
FbNcgDaU\bf6@C6KOY5cN./@fHFH@C(f/f&eGZ#9V,FNA40_[LAZ7@W39D4c.e+:
eAP86_?-)R8>CMU-7^G95^1M)8CY#HB9XfS4CY&5NKFXF6L6gLE?ZL:bU-_#5:17
(H\D&#gLVZ,X3<b1>CT517P1J]a88RL6BWUNGA.cQ47^KS?GZ8DD:682?,Z2>[W4
60T53cH7PGL])KB8F241>#9]D_JIFDgNX(BQ/c^00@>1GVU26>R>@)c.M;(A4&#U
2>cOf(V(>aSPR@\c>5S+2I4HO]DI-WLH51OIf@Y.-&X_S4GRSH6ROS1M5R6\Ie)<
_?[T[^+)&R@c]H)U?W=U?O-Nb)BW=2?(5AU2WZ<@=dY7:,HH1&NU6^P?STXTNWXW
SCRWO.BU<e.1IKbF8D\^B2PEU/F;R=6>B#L;OCQLQ6XDZQ/9/U+RTN9,UK7#fJRE
eBcYIQ/ZI2Y-b8@ZNdDBA=QDGC[X6.bYD:N#&I3)LZ@f[EMQ2YL/\3@C.=#U\,+T
7C,27XF4GgKe^QB(V]V91KD4+5bG+>Bf4=O^_)f^Teg5F.dFKJaWE3RU_2fTWM5=
==1..P<5G)#8I&,c1fTJN^>0QKDA:?A@;2T-03(?52L0U(1)&YXZ]FZQJSV(T0J;
9Z5##>a5[?R(\I+Fa[[0-c2dAD@L>XCXP\3PZ</0_6\bQ-;.eA52]f<R:[;[NP0S
B/S_f.eG6BQ]IEBB79@3>_MW@F6B3bQ[(Ea__b_@-<:,U;5=;QgI<<7GEN7ZA2?(
U@abKJH4FYNMc7/\8XL4G/2PbRa.1^N=N[Q+--ZDWD0[LN13?ZE.R/KGYDf2PMB>
@\&d@8eb?+;-E#:3+]f;Ba1:N72]USg8e[]+f;<^;T7]_];2K8,5?SAId<=;<cO-
LA?4_c0#Q&=7+[#-J=[V?D<,M<4VYV_G]U9JeTf8U+N2gY\O6+II.5L:H569^/H(
,NZ#3RCRD>_,3/D2Xg/_C&;O_3Sb&89(aDXQ.[5QQKFK.-Z)&N_b4P\d=-.,G/S=
[@[H_W+1AT^BaOQPC\#0<R[@34F,3SPC\V_09++OcZ\C+0E928^OE.8>]ZaAU\b>
(:T.F;&<=.Cb@XUZ7NP-]>;C;MaFZ7Pe(;?fOC(),G=CYTcB;G)d5]VW+,D#QACR
a_^;<[)[9I7O)J4?J(URY/Y9=.RMCg/edL4HB3=WHHEHb7C8]GXG+(?2G:Q&7Wfd
N06eP;VN96]Z2[27^]fb(N.</4OBR@1,AS^)M^4F>TT[?;I-&Q\e__e9&UCg]DdH
6_eH=&;GcR,g6]eF_Ic+=5+0=O0&8K7L]]<,L6=Qd3S@W,MESLNOeG1&:f.#C/-<
I;a8Ed=0G4<-VB#L^f.)a2M-KF92/@Q(18Xe)M7U2[A<>O7]P>XL150,c0^eVM+C
Ve1P&M[E,>XaYX/D<#((0(MM9:=aH\2<;:=0;&MV-8))aCCZZa3?KEcPP_W0f:C\
5PB0#@>@O9BCVc^88^^@GP.Qa?a<419L@NFg/,+6c]6WgC]=0_FR\3);.bU/<V+\
g[[BWJAV.(7J<6e>.R&ZBaN]c3_G0#+MfAI]e0+FCHa_DE^(D,WZ]CE/P1&\Kc_N
;TZ1aJT-:9MK2V]cGCU@gXGIJ6?X:bWKfPCBCEB>?@.5JCaSL083YT:Ig+P=_ZL3
-IP9Y]\gT_:O0K\ALRb6If:=,beEZ<?5BcMT)Q4X63=TgD,ZVZARe?5O0F.1#^J/
0D)K:SU;K.3WJ7\)IW?B_@97=UN\>:F@c-/J8EAZQ:I@bdbD;-f02(J(A07K1SVJ
I#ISfSZ:1\NdV+X:RPb]RNRG&9VEM5=^)4ACN?Q]0_MLOH<142ZF3K=6YcX\GfdJ
Pc+=P?U^;\,8F4AP+C17F89P)E03Aa[M7,0;X];bT,48HQe]gfX,<)[[bYF=JH>2
#6]#,9(_bM04Q#AfgV,7P5D69DSaH8P.NE/Uc?H:X&_S8QM1VPPM\>G[URXH6C[.
4_aeVZc<_\4@^9L>UI0H+9L@b/IZR5Q]c3RdHG:)TILU6Y,7A9]/Z>4=?QDH.4X\
OXZ68F;#We+E6LTD4\&cY5e#D2=2Q2WR)T4Gc^^,MCR#+^;1\R</e8>cf4NDCZ>Y
_]=BZY&O?1.];=PCX:4CWNV.gA0c##NI/BWXQ\R9g=_c3?X^f_B?HgCE+fD.8V,,
J][PAR,S3<.D0>1C]38IQg0=&a-O4[[09_f,5UW7-U0FC:EFI6PPU#QWV>X[Z.7M
OV[XS/3BNHS:2YE@-C7RE.Ua+?5+O\YD+AE+NcY4gE^Ebb]9aNbF<bP],g84IT8J
@6^#b;&;dRX.+PI0JXT.H)+OB?KfaPR=YX?14Z4CM5&UAGI1XY)NaKXTRG+J8+K_
EfNJP4Qa6-eg+4IFQU4gGHU62]?c,Nc#DP5F^U7Y8<ZZ6I2AY,CK9],[YDR(T0W0
;J:a9-a:5V\J_F5:]f8=ELKfA/U<WUPb=8g8<eK-Y)3-P2PG=J9C>4R_45;7K[.L
B)RKM:._W1bDS3NF2==d)QS8GWUJ;P0O)71R:WCPE(7?J1aXeC8>^JQ>cU6]Nf-f
]ab\->e,^ZWC:VJG++)TC&18Z)=gW,FQ-M^NG93/OZCCFaa[A(2Q=AK^LcWCNHgU
FaHUXeV]6,S3V/N8=bT(OP,9]UYP7]fI[U@DggH1&c:9..g(?MVCM6[9(Af7)Q7=
3GM1b9;-Q5][=G[3H.TNR?6c/M<?d,>P.#D=RZgQV7[@eG)/DW:FfK7YXXDe7_Y\
CLHRdK[V..E.F?/QL_1[63IAa2SNBIBW][E,ZY/N#.EC],Ce,;>c50RJJFY++K</
S/g)H_NGDJ#a7I.fKVB19;d23#f0?B:^L[eE(6XO<)Dc&O:<MZV2;J)<UALWDZ@F
&\gfYc\T;^Y+WXJS4b8BE2DY\a/J>01]3\a0J+:]g/4GW;8JZ;(bIDVF@IVg1)3F
,J57e4(.c:.@JHTfEX-I.9eG240OB7F@g=FC[[GWg/BRRFIc@:2,&3IN?\cY[Z@Z
Mad=\^0(Y?10gG#G?XWMcY\AE(YeHV6D71M&&+4Zf[^5V4:e+dP6gHCX;EPaL08O
K[TC:P(UMJ20Z:)9L_Ucd_NV4,O.^=;HW;.;4R3[6fS[XL9FK]g8M4FY+90VTP(Z
E906bf;(SU<)TeF#9YBQ@a9/@FQdCZJ)G]878]G8+4X:Z8--8V25\dTH-[VZ,W+Y
N/8L1_B7?Q@^^?c(=6MCH0B?HX;153]9IPdZA8X,dLgXW&BSNJg^_P]fO:C7KD62
FMJVLUGHf31.>KbQCG1,5/;?VKJ-SK6-[_UZg>QdS97Z84]0R&WYWZ4KQ0N>2Da9
ce59I;ca)<d<d<;fO2)KX97a0HdRa;\53LW<H[5fd3N>c6YR,T-,Q[f:W4_Z[(V-
?WNLE<>N(-e8.Q>Ec4d)24;^)b2)^?g]71U^3&7DJEdI-NS1J<aU)5XCJ-A#R82@
c\&6a?T-XV1&M03/0US866cL.GD-cK-GeG2A1P-R.PP0M]>664.>2,<ccb,OG?Qf
U],D?@=V@cVf(RH/>Ef_GdJ.;RA)CW9e8W_6a&)4RCc=>\(cN:&HD7ZDT?EYcA6_
IdHRdN7-5/e2-#H+R+Kb;VN229H);OW5>KY20KGQO.0MVJ\:8(#,FLX:NUIRCe7E
cXON4g^8-gI>bZ[]1F72#4HXWT4&<=f^RM)#GNC6;E37.(T8>.DdK0S(26-=5&8[
e__Y8Rfg1XPCccDR57Z;IH4O1NK)/CURZH<+/HQdPAD-9H_0?WZMV(LI2E\O?1c8
AIR7\:J)&I4dK867e[3U__eSI8K>Le>5\#QW,?@YecF[5,+0DBOT6H;X^<bZ62(H
0-XA=5WT:/>T]FN6dcVO(;8URQ3FW^a]^R.\]f\DO+TVX;a_DCSWg2TEY#Ue/L.Z
f;6URSCI9QNXVf_78(G-3+<#YF^SfH2b,4Q9Me,XL)Ba<+T/GD/O[g1JPcSV,aX\
ZMe,36Q;^#2N(3<2VM@UUf4#e&&PUB+7VbcA?4P8:d5De>LTG9.b1Uab^--W:IeR
NMLJ4\D>8ZOCD3-ZaI,NMG+W1:YKWTZX5WD+T&WRM,VE8H4TSb5I8cZPZF#WMgS<
&#f(gMP^/gfD?>R<2\\.A6#c+JZde_U-,c:HJ0_ZJKHDYAA7@]AdVBMQfBME2a5/
AgZLT9LF<H>DZT>4[]f=A;?G5__QCAX/0-6f#AZ,R56A-Pd#dU.X?[BXfBE(7DC.
3-&HNDDBdN\9A.LD/SR.f^f7</ae:&D??.S(S2-6>2_A;/2-_aKXGM2TLDgO+-O9
_E^>^P+eD/M(<XE>8)?0;bgA;f;L<Z(8Y[5BY?)OAR4Sc42b._;)2N:FMU3#,6F@
[6N<I&WgZc\08eNSW02gQ./D);&aI3C5^SUAb(M=7AYY0VJ]_R&7EY.^FY0Q(IS3
S)>afV,=?V(eF)_Ge-acXE^[7O\HZ#L#NOD-7(Z?>+e-0R0dNN[UFc+Z/T)-QDO#
BE]NOcK>1;-IWbAgG9T\<+68WD_bQU\b8ZZ_?KQ/]^Z+DC:O^W?36K4>Y)>3[b#J
T9T3(/&01VP[RO6@\eDD##D0/C<ESF+F4Y@,O5X2.bZON3M5&&^D;_P_>0>0(_gP
;;EF2[:0QEB.?K\O+C1<F2.P,b/c\TWCU>(+L#HIUQgZ;18+<5>&UZa/e.&YFT[X
MF9gE5JU8]3?[OMF+\9/?:dcY1O1X(Q;>cE@(Y#(^(]/XYE/A<0<,4=Xb>eL^?.J
7W8AONGXbTD;DR-H-E\[AW=3aN432L?(+4LQ:=]J.<g>_R5SORf\E5N;P.GN(@:H
F8U==b,a1SSeaScM=03B8X1D7UV(VL15SKC(4gef9?=6JL7;)d_I]&R.]-6,J^;^
U=W]\<a,:>SeDH(_(E&AJdZKSZL8]\[/8aTe9,EHP^7HF:]8.@HI#dTE.ZYB7C(4
F[E@(A0<M7&MLF?/;eSJZSg+UW4N:8.&Igg#5#,,GJ+ZLMP+5B;^UG2;^DS<X/Y<
>HdMW[:YD77_D7>2+^C)1PcVf9G:>5Wa^<:<90f<D^Y^/,>;a(g:b#N]H@FH81gG
=&E]^):GQ^HCZQ&XQ+<\^NTG19\b>:TFgS[6N5L(U@[HVf1XZ@_/f&g_-^e9&W;W
6Y1:O0US+b.9Q,GE8U;6,A;9++/WZWUDD[f\XLG#3]D5d42@>ceD<eU&BeYY^W+.
E6f)4/GSYOWWFP88#e>,(30^>>Da&UHFCXW.b?dC,<?]9M[KQ:\2DQ9AG86b3)d>
]KC4#))PL[f.&2(N3b]VZQ>&6GY]9;@b;<CMbBeCYD&c_a6BQW&5#()32VcZ]:AY
bFNTcA)\Hfe<\b^A(3X#,/NU=CJNO>9b6HWB<-;C,9N]HLOGD(YJ1:Jb4OO5M4:.
.QgL<.QDOa.]T5W0?:#9.8-dURV,Nb6GL?gW]TE:@T)81^NN+8U=4&^gd+V3UI7^
5FAKL>P)g\+#W;5Mg;1bTK0DCWZ=6^4DW2>TDS(DJLI7a5B]cO3M(X)K2YZ)L,^f
J::VOQN.,Y1fH(3=+8P89L24US11S]CX8\CI/86TH(dF:T6<)>+WLdgb<>a_:WbK
JZW]>a5HDK=F49[0gc]<4R.G#1PY9V5J=?\f6P?:X;R2bNYLZ./12-Q4Z7MC^@Z<
S.[/cYY0TS)U;+HNCL)V=D>A]1V]OG+7Be?K?F/#;KQF9e^CGW=BIP71NH5bFCf=
//b<5YFJK&@DS\L8>X,)Ab.C)Q>[dPA)25TcgUR2ZTaQ-@[Jc+_A7Q[_.K?S5EN?
E+;OR8^S1K&ce@EV3cbC7QY8RNJfb+N@F2a]OfF1^)+6D9Oc?UBW@B2^R.<K@F\8
P((7-&:8[O-/C:FL;g;GA#=5XD/RCFD&#f3YFS+R4H7aAC-S>3M/I\gK=XcF(6XF
bXS.[-I>NU:;2OW:J,5P>Y6BfNY@@/PO#<7eKaOA:_L:-a1)X6,U#cbUASM;]@[L
ZN6;X-d.-af2BZb?_ZJa.3XE,N&)cX<2?_U<XGV040)X6>eWX0J)Z;&e#=^feTO^
cAHc4Ua+.C6RC/58P:#^DfAU\3=K_P,5J2If]LZS;d_KK1eb+&3<J^YG9Kd]>?Y.
5W>a.C5eK88]9)]?+6RKW+SIcNG1;A]+GgZaG32S^-&16EM]bEPcTBY5OZH+\Nb<
g?1SLe(<MFDe7&b2accMOdF5<Q,E^7X0N8)S131R)_/6C/=1NLU=c9e6W4W7bKgc
#]@W3WV,1MC?2>YR7=&#>D-.5<&M&>,MJ/BZIA:eF7UN@4P=Z)Lef[M)Y0&<eC55
W7=aE9]<->cJbE9BB_e,(e?QVL\#0)2-RH=1V&CgXV#7?&6b(IG+\[OD<J:(c7Cd
_F,A_GHG&fECNJ+>7\;Q2J48b?O.e.9;RR@DD.a:\3Q7B,G(VXd67FRg38_XE;X#
D8,4A-.6JVNaaFU.^GS.g-P.#E)\-P#&@H5S07##;237C+7G@5:P(g9fDR,=X(e-
UI:g-.F6abNeVCgS>^-,UP1=,+&-/7YQHQP8U)HG=YIINTI\L561+<0gZCM(<VcG
-S(cdTg>0EO,)aB#LV26;M,OI;6DY>11T[MGFD^>B[bH<BTaEI#[Z8@g4H/dXKID
=T?/N)T=e?:LfMNO<QaE(YP==)H9A+OW8OSE#LKH4&PJ]^EG.)F@La<\@T7I5.Y?
a4XYg(e13]RbG/I(#a_dKd<:D]7^?WAc&;/SN.W/<6Z]QAXSLUf4KK7O^.bUZO/;
2,1E-,5Z8J]X,&WY-#K<(:IAH4+4PTgQI_d[a:5T1fc[:;C;)Z0#_Q_FBaE(B11B
MAP4(34afT.D\6QP0(2PR&G&QI2;;SBdYVF6(_]a^30+74;>?,gR2@^:V.=I>WMU
1L,10O8K,CH#1:IN4S1H5+I]I02)aa+BHKAW&M3@@92.)gJ4DB&;&SOM#?@Q^-Dg
NQ_<H;dE>:K2E;K1HZ.79#Z.1g(_KCOGMDe0g4J#(O0<S4?0PMIWKc7>8SSV91^0
W+eU\3UYBOK\b-T.+JEeb?CGNMO\OdM?2Y8T&-VHM2H)+39YH?#V^B4[Q\QM.g?M
Fc<,,+0O,8B=M.3:TYYQ^3g^\=@CYHKCA8Y4Rf=\7RD\@#YbT8;_/)LX,1@e4]#B
@@;)GC^#&^87A85GO62F&JWG0X;[RF(1[/X;]Q9a3WI29,[SABbWM(J:<WD&<:()
Mec[BYN=PIX&GW3J<=/5.>FVbEQ,A[YP[)#(LMZ5:C[0>UG@V+8Y@6+1a^OYbT/e
_#+fLX>^_E1+Xg<E&[XM5OAI-@3;<5JY8UJd&e+X=C_fNeDD/a=#-BNT^a]L6E;U
c)1L3abb3XMa:^:R,b\]8:7VG_]>AW3\YJS&-86fJaJE0\]Ffe+dDS7J;=0>d=AI
<]D8A;bACcV+M&#TEBT(B)&C<@E?[\7eWd^51OTa[?=F#3_?<O7#>,X^G\,8I3He
7ZVdE3f7MJ@9[K_,+S0Nf9.\Kc]cOAb5AgEX:=J<P2@=Da[QAI5KIOCX30_E@gKA
(fBH[F.AF#S^6968_H&QH=F>)WR<C)O@.]c9W[f7Vf[O@DC[0L(2,P1@V@LCc?)=
FARN&#Y[AFOF]&b<g?1MNMM]:\G+]UZ<X4#85.51+IEf@a,AdUIg-0A)J-/,MT#D
=d#S/>Z6?e>9<=(e[009C@)aXMT2/Y0F?:;>Z_+-&B<3ad?R;Tg^UZ&9^e@1Ve7&
.&)>Sc<Dfg1&@bW<JC-65+2U,6TGTR^QB2OC,gP.>7\7U&VF_Aa&bSX^ZB_,^[FH
+^TVdT<KK@X305FD_e.+^&dZK)M;<)VJf_AZGV1,XTO\-<D3M1ZJ_,0\N2[I=2BX
fNBSWO-F]#WgC/]TMTI,-]cfECB^_P,2,5\N8gPV/5_@[Y22U-S=+->MR)^O7Z.)
I&(+e;VH?EVF][\:_G@&Z)<CZg,/Ja&4J4TXW\Z>K:>^R;.,0d:V2>8Z>bZ7H1C:
05>UXUIKM5LUcYGVTOcW^HT]e-80QY?F,.F)VB&8cD=YES7Uf5Z96HTe5C&O[CP(
CI#Q.Y@8CE[ZRIYbB.DC4IR[R=]GK?5JS8-AHAQd?)PF+D,#@-B?-&6(IH.^=:&1
X-Te=MQ7dSB@<Z[9Y>Z4AXEa5N+6M?]6LAJ@M]\\4;>NcBQN]K#^g>WFag8K338B
N.>LefdI93+0B;gK:?g-bCJ(W=(S-KcN1VQ62@S<N?@:=QZ1K]T^NV@)-F[NdR:a
X4N?_CT0GGOT+2[<I@KI]d7LZbT0Gf6WL&H@FG9SaKG3[7P>8fO,-;_?OB[URL+8
_c6^.KQcE@#9OG33]d36bTEF]N:CcMb9K^48IgFaAKD#e^BTP=[+OMYB2T:?TaaL
f0_cKM5ZCb<K&NA&;N<UI/O?:8?9]GM^XdBR@F.)?0(A?gfgRSe4;Y.HM7Dg>@_F
c^X)-[;c=0A,]Z]RS]KT8)LaD^@+=9P&8NV=\JF&f(f6_6W8:X,?8XC@,(&W+-;g
b1RV(:K,8>X<VMF@We;:71+dU;MD)3#C0AHNDDg<4;1QC0eA^<@46LeI06ad=BG7
a:b#N;7P]FD55JIU5<ZU>.KV,V].D?D8C;AO30AL-&<Jff/FgPFXfE-LDb;I;adG
CI>FG1=87S^C1L;<(d^EfLMRg/FGIKK<J6,6?)Acf&R[<.&8#)bL0;^__dW?JIA3
bW@A-N]K_U.VgUY&T=UR5\Wf9X<8[&1PF::9>OZ1/UHc:R#<@bAf51,]FdO\L>M:
f9[WH0cEC_#e&f55>N,Q]I&Q_5JHV/L,e.]IQ6afeIgE5R^7+=>4I=LGYWS3HR[(
NGY(d[aF<[:GWf>Z+]E]SLU?gOWW/]6]C7[;\W,[<(2T[6/(CGTAX_VZBe@JLM8e
Hg#=K0DQ+aU@D+aGIRGc>aXNR>?.<eF7L,8-6,;c1Teg;TQ#C4Q6\^Zd99+Z[2]1
EMN,agdJ\UAT]TO17?^Z(V?A9YPMQEcNI(XWRUQU+C7;N>PXLWI0)]UcY)U,eFL+
DM#U#Ae^_?JA\:UcSeH/FF8?HT#\.#5Y4K(/T2aS/X=7W_>8eN@JOYgG9a=)ZG,g
g2KEZ0?#^bWD1Z.c3-3bF;Qb;K#]I15O@LNbG&BT:@I-WSZQW2[8=OWKRN#MY[Z_
-:P8:Mb#J>R+W]&>W85e>.\)N+?1#P^e=,EGCfU//V1d@3U/ea629aO22U5J=EJV
b:a@\5R1<EROE+CUP:e\U3CQAFKMFWfGN2S<:&Q<J&O3:M57V_Eg=-b,&PE15ZQ8
fU\/@:MBPb9YA/DO/b:5.JF->f(O6=;^g=;6g#O)KU7MY-A/7=>Q8=Z#9I;H-<LM
e(9(M]V8Y<QWSHX[0;OUWe@dRZL/ZGO)3=E]/N\VFWDbLa6_?2;1g/DGBRD=,V>U
4a[744,^S]:f,ENFXC353IKMNcHaFgR6SULID0#db;.4O=CL88AKffCM+4_;O@[c
V.d,#4<[/(P3OZV2:50(LPAHE85TS65c1df;gT+//<+RL2>-egCL7&L+eBB4;>SO
X(KXW0,3afV1JB>5VZ,_+OO^8S8a[T4)+Z/03PUFT]],._[)\Q:+f:^PXYT>(YSX
K.]VU^],W2.9NgP[e_S,b3c7Mg75OQ=VI>X29Y?8#;J7USTETO,DZ>8WP:0g)a[:
KfW,JW#.g1;Q?)b6GTJRQ06T-)(DR1g\LTA&/-3<)GTcX5W<7Ib29(b#SLd.fFcU
=YdWDTYI,)3;4ac]-\f6M)R-CDa#B9=c-Sg751I>2@gB2Rb86+<2d)X-f#?(Z&H?
I1RV]3\==9[c[#GPN[ZSP<_5Z>:g^Kc@a+\F=U+/bRSMcE<]PaEZV2D,#g3X+?O6
+361R8ac_eY+?^>J)];YF5LC?eAKd03IVAGB3^4385:H;[<E+B@;3C:eKAdJU:Df
8KUTTC#5N1eE55/)IgD?CFGY4^LQ-[XO;[(]HMaDN.FR<.EM+)XOG=Y6>#b<J6dO
=ecFOgZ36[1/JSZ@<C)2]9[H@=g<E+B,/??>e#/L6_U?EaD78F&#Ja?&c.@152aD
Q/.f=QPGD]E36<89GG4,R,7KRVafGA^+7W]I[c8a/\,e9,M8Ob8&>)^@R.-GW#&d
G[#:HL\)f#+;Q1IgJ]TZTgd^]WIfL++1&;(]RF8<<e_+7O?:c7(M0e_F_C3a:ebZ
(0T&Y)&\:XPAHL8X^+DdC5Z[J3cNY[P)VC@#a^fd0g5f-)M?)gcND^NSKYEe&SJ<
S2=MC(,G/HK+)Nf//SL;H];0<J=A0;<7<,5+@/S[5Y&DT#[,P13RLX=ROLGM;WH7
DeOgMW[VQ/<<16,IWb<2aK/]Q;+3_RQ0X9UHMZ41BE_[K_5EFH/S<R>/2fP2>Kf@
<ZbQ&PWXg6WM[XWJ.Tf7BEQT[)G?8_Z(]DZ5>5Jb)O4OT8UObV4[GWcNZ#LP/#4F
>gC&-]39fabXf](H_I^#P0JQD,\3A=[bLXKX25LQDc>(&MLWG<R^(.faC<C+Qcb^
1^;UN0&fSTI91@S@G5VKW&gG-f\?X\9MD3f;5M?#1=eT@,3#2aA0_eMUI?Q94KP5
&+]N:FNP).#2J=M5.O5/X.ae/3_HXCL^aa8Cf_g;c^RP5bSbQ0SJ=0UV&:fX2NT/
5d3#12VG8d-KC+^(CXM@+O5D&?7)?b\b0=174C\(WKZ7g]-[TPAcA+(OO)ODgcM)
DEeC+T^]Zg\0+L7aJRUAW573ffeGcg2J&-E2SOHW59\CF&:<=+O1O95-=>^4PF:b
.S70]W)8[2.Z7;JD1ZcXd5K_QJTTGL+;T,ad+Q]97L3W)/;Hb-]7972G4NbG9g-Z
?;CeQV)#c_4cRL6K<PN\9;15+GAC)QNWgYMTX#9JcCac=:B_dF=Lb[gDMS_Q_/V7
><dB7EG@f2C6Z[b]]HB+fXg/4a6:=YC2]7#=>VH:+]5MHLM\1cW:])P#Tf^]DY3O
Y_V8F;U?X4+YB6JCSd8W.d<dVI=P-MGc#XJU@ZWbKUFd7C>:/LE._a]<QAg_Z)[+
(IBeTeC#EA:bW3#)Vb[/:[JQS<.=(_S-Ed[E0HCN-5AU,/F6(,0de/6W8V#A:BR]
Zf@R-#\VA#1H8f_&VPF8dg:6.@H(TPN4g[MJ8>>8M^Hf28A<3:5\Y=[+IU/E>=R\
@e?^6V2D.Nc&&3_DPH1DfL_aKMFR#8^G[cd^)=b)9<7c:]/@=1a[Jg7G:e=_RKG)
4N^aW)/a,JbYGQNDM[O8:(0_ROI,6.Q&_S+_MZ+D@\SQfAW01GZR?UOBFHHS.8<P
b^\-dCI-[->ZKGdS.\?&T\B>,0eDYE55^CZ@7GQKBBfEP,R^+;[K_Z/(SeAX[:G=
[Ne?_^K;&R/[1A=U=,O;Fg[S];HUEd5+Va-EL:;X_0E]Dg60JaNBO@E[.G:N:HMJ
NC(Gb8,8>cXC]=TN9f,(;F^FDF&V7B?R[/AZg_VX9CCb(_-+RSX]F5ZE^3,NR9VP
,1?PZRU97CbF1QT6QD@:.5/49)_MJBDSS4PMO:C?LIF1SI1XEY6E?>:D1<S#TQ@X
cPDL3Oc^Ic8VKGJR-YMGAdI+e@Xd@g.PVVT[Y>&3,R9EbeO58e9W&Z,9]U]AW<;R
&B)UV>b2MX@9X.QfEVF;-22O4g+HU7[77]f3#1(1Fe7^5eO5=6INcC2C8c24X]Fg
O[B9?GWWa9S+I_ZEN6M\,ZX2IVG,Va_D\<OV?[Z9G.4Y^c;\CKJ3FIbFR8Fd8d45
WPJWFdF0.EeJX[&;]7S?K(/Q3D)./LCd4T.\AU7>J_&>UTaA9?GFY;L0)H\RK);4
CTD,GaP[_Ie&(eLDS7CM/aAD57MB[)A(ULNSYY9)-SCd_QVLcU;f04ECPHCe2^-6
;AaV=25D@OQ(a-6@,ZT^:8I?KXZcN7N6)YV+TA5FJX\GC#\cBXJ349d22D[KAf(^
e+B</5PbQQO:?f3IMU_(32d[DDMcP6:_+_U-UfgEB94^PIG#KTM9-LL>(K4^:A?C
L/BF#J\e7O,,)6XYPSU@^)7N1fBA(#;29HMB>?fAMG/<,eA+49-?9=;,ELCe8VcF
LKc@ea-@[4_IL=TBBRQ7@<R1<I)O.W@:,KPQR0,8.V.)9DM=GM3&9._ED)3V4]Ag
9ZL.2d-76D/FVP0]ZR6>XSLW<R)a8fYJD_\OD8ARTKKJ9]V55B5S85./Ud:(PM7V
V9<RN)<,[b+HDAS5aHT^&a:A6&@cA,^&#^Baf-EZT[,ZWHDV_=H\+bQYg\:01/W[
Z>9Y#f;-E@efD);-8N#cM])T[?\O7]OJG3\DC:;4)(QM+LNJ65&:FVS]H&de#IcN
H3Q94PbEPcYD-KKO]A8[R1c,\9ea6aGM..J<ReA?S--04KNUe><A<JL-9bE+?0Wg
5ND>/[O);O1Se9XF:>2DO?&NDZ69adU(MP0e04CWYLAc7D>VSX-#/VGNKU]AP)YU
WGWBeHF97D1fHPMFAM)^.BI+6XF4(RIfXWeL,TWJgGMUb_D]T20fT-/6;=]A/(_2
P?,eLTR#5./Fa>6PdBZL]6NZ).^?H:X/&4Q]/9WF>a:375fD8f3.<4Q&J&#OJcT/
KP0HW0Z6.,DHF_LWS2;FLW<F9(FcIU.T(34NZW.)\.fJ[BV^:XRDC[]GW_ILM[6\
.2LRJ4XBJ^V3G317#Ha\Y6N5^S9@Kc06g(9RO;/[3;9S.fG[V>52DdcNaK#HB\TU
9+245RP>+,:/XS]H5+Q2.SWAR2#/c#TL1A?=9/NeH43,]aKUR.G?N(D\]F,?TMUU
[M0DWDK,Ac+/FLf8BY6U?<>89=9X_\2W)]&NU24(gE:RM]U7KSK_U9X-dJ3#Y+9Y
I/&/T(&MVVXH0D(MRDF7&\eW4#U7A&Y4b):@#?BAUG5<F\RQ-[?DS1PD2B<6_J#c
HS(;4U3JBL8/.V?0dXZ_a1MeP0DRcQQAK\KEUW;G:-ge\#6XF/ZcJ)SLV1?1(F2Z
].M?.LeeU:)LKH4@Y0J7cNS1)Q-UYX.Y[OA]C2T2;W2NJVf<g18H)KV-_@+7c9Na
@G>>Q1aLe/8fA.J>&/6P>TBf_K)K>WG#fNEPb5?K\DTdD=..cINJ3VN9TE=3K2E&
[5H:HZFc0>JeA&6<D2I<5ICcK42);K3/:+N+d\g;:5AADI?TE?d];^VYN3/U_;4@
79P))f3cL[e\<^\2)A-g]6(9e/-,3G,VPb]?37YZQ:3_C>M3L49+2XT)LeD1EWd.
I;]W(/024J;Z@MW-gJO2:f98^T_G]HVGI^H)3[5#&7OI<^9\<P:=9#e8[:fV_#/Q
eUc29FRB3B8J4/8ZA<FGDH+M>(8F6-P[>f5gb/_0f[O5](3V=<W#[b-QD@N4KK1#
<ZU;ICU=__4(#d&QCdR.Z@,D3B]Y\eNS>2C7@_&bW797C4Fe,Uea1?d#<D=G?8#]
/SU<F+SCJV9?:U[eEb&]9\S5#\E^[[M^M&C_g#7IeLHRGTeX/O4bE-8D]F:X\C:H
gRWF)?/[6P;,N]d]fA4R@@GVT>X:R)PU@6fO;VTd/dZW7/1:\FTQSIe#R^W3T^J5
=54TC?gYP<[-7KFGRd)CFC\Ef;d=5/+](^\NM5).C@_IE&JLgU6dS;M;<+6I1_(I
F#X;@eE+M9>DdR;Zc6S41^E,W,[7AbI_E15+W&-L\;;@[8D.>YcAe?/KFKE>K(Ef
0]H4_;5Z>^A\:Jd@>RWO^;PgC9&FPBML)H@:ADe@M,X/P>5-VQG3UY1g9B9bZ;?<
1fG6,(GAWTG#aO]]ORX[a+:X_U&B#VA,.]_?(FBd:4&fb[Q/fAeNbe,5,WV<V7Y,
SbMMf\L>AafcEIW@RdP_Ya;8BM1f(fTaB]EbO_)Z7[YTd2<ND;Y,LI:7LG1#^W7Y
]J]>cU&=7]-\LI0WAYMD8\6>e_X8cC881^=+/^\[VD8>)VI)Q^D\2d7FW(:E7F69
/fd)Jd(_@&0bRf/]2ZKd^\a\Z;0)V7L6R-./72/W<R82H&3^A[V@S.c[cX=V8EG5
/Y[O/a3?6f70cf;d<?+>P)M[:@KVB+0O&L\<EBCc2@SdR1SK,cA51ADH^8T2(E9P
R,[,W&0LWEIV&BETBL)^>[+/\O)I6.A3_WX+B7[Y.F5^42M+;PR1aX#AO7S4[geR
_JJ6&bI\_Gcd;/DA>0c8\QWX9@5,N-a:f:#3J3f^^BQE;[Z-dW<1WN7T2(,+.LFW
L#8X1X3F.aVY_L(;HG>7b(WK[GSCe2Q4N7_6I_a6@L><#9BgcQQZC0@-20-\fYI7
/,:<f4Z]6Jb2UfBVH6RdR@0T4gbQPMc#A\(Z\-O6Ldg?<KX?R\(9<fPb>_.8ZdJ^
L4;7/3@M&IHTRGWS;Pa>9CWf@2Y>HT&VE++7B.U&OdNZGeMW/1ZE7QM/F:fNUg/[
WA[5MJNVN@Q?\B.Y24BN;F>,aN8=N)9P[#B/F<[9c?_PL+aU?][X@a?^]1[W9g<2
(PY<V2I#Ea+)7RG2C\CDId5Y+,52+-U.YJ0_UD.NTIc(LN5V[;IR_@eU>.#P>;YZ
9f3^a[c#8-3XWXf:G:95Xe[S;7AY?]G,E4<^FIG6-S24R]=c8/ff98O#42C6DD)K
ONC1d,@T^EFC9>&<N^Tg\R@4>;NC@)Ge^B(5SK3.U[=(P^:-M4_4H:=a[GW-J49E
a:Q;+QDCL-6A9<\#(#,03J^A9@KX>;b7L_e^&@ZN[C[RO_\<(P_Y\FOYW3:8=5U2
//9:g.cV-G1.\Z)3\AXD5EOdgc3F-Uf1O1Aa<e4P>25^d[+DHF6F-OA]5I<2S(BH
AT>093c-#cR-Vaa_+7^DBT,[L@[EC0KgYP]G)5+K-e88PA,AENJA>-,XOXOEK26F
@&<HYVgg1VHb3/^(W_=4ZeC/d9a[0.E0\20Re:f?KME<T)f6d^g6:0LJXV#_<6NJ
EHG:e3^E.\CcLH2bDQeDR+(GO35@)(=I0I;[0^JU7c5L@CW]SU&95P387Y9K[U#c
17+N58U^71.c2EO2R>7Z6;)7L0\/]OgGU8NQ:VX:>T2V)c>Ab-UP=R>W[;J(cDEQ
GAF&[<aRQVTMRA59(-EPT;,O,3?VHKU8L[(.KGB,:T/@@@7A&K4);Y97:RD1eQH/
:.e6<fZ1O17+(0fb41L6KXN=7YV5)2QE>7+W5/c7H\KL&8^e5VKd?cZG9gZI-L=f
fLBJ019fSPbK92-e9>.ZG=LDGU#89U7YbWN)Ug90N-?fD1b(gUZLCX3]5ZMD)S[Q
H0G7R;E.0La8\DW2P\A:3,[@Oa[8/Nef/@\RL7e6MT-XJb)ad-@)cDYfY.#aZ\RT
:_+d25N?.QdTKR9HT2T_X6H/)EAWWJ4fV@BCZ/BV3<BCOQ1&_10&/#JR:2ID.PNM
+://F?F;@F60F17QX8-:##81R/2PE+)e5cb6P6=S7;daM-KP?K?EdTGE8dMLRFC[
,OVbJ^c(L^LKKONQ.\Pb&E4OBCS)?WZ2G,U0)eS^baTT;UBc2MZN:Ke39\f1WVRX
[+^)eNX+gYfHC6fd3[6B,XDGI[[HEVC)-D)b,^[\_gWMV+^0S@)bF1=E4]NOBMQ-
X#+7KFA]EMMQI,58G#(#R]I1P4>.OA78D99gV:[:#/F(^eL]YVZL[L+OYc:H9YWW
:g)1]9VDZUX2J>YFC]OfdFHY-U7)5f],&NaXBIO6+[_V+G?XWR8eH7+d/B9B[D8U
:2IgL[4E[H#dZ/#\?eX:b^IZ&2OeaEL^#6KKLV7A</gN3+L40FJ]RFLeC=JMQ2F3
=,C+Z6;U61]7R-(?QJGHH0DV2[a0Q<DIBYXOgLW@>UJX3AJ)/]ZX<NJd<;#D>>8T
+=SRB@#1,;&d)/S.[^4Sa-MS<5XIIXUc=<VCSK57UUg9RI68RO25WJ^\RMgO[d6,
ULT-ZKX@L10YZ?0MT?R\[de9S/J7c\NJ50H8,:M0-.L=N<a?Q[-Q[JCU.(Q#KP5d
D=<9FXXCWe/(ZX_JgULK-0B)8?:X+J44>/fVIA)R8c(b1;0=>3XCR+WMe-NZ0Q->
/+M@Z\PBUb/-U1U9Q:3_=\);QVM2DK&cLP,,MO@[?=NQaQcW1]U,^fJ55Z:-(Wf;
cfTRL]0J:Gb4F7C<4:BU5O8?b=2?/5>QOfYZ659;,TY+[)e.NT0ZZ\^+8d95^KQ5
LW/1geMADcWIZ63TIeASe1ObMK,+Q-7g?<STG4E9W#GMc)6[Rb+O+eNM(eUDf0C[
1&OVLe>?Xg5(X_)9PU3fDONQEXYA;:)JAcSKO(:dE/a)Fc<=8OU=@R0aRB:RS/9_
?BK9_O6IgaJI0T\B7V0/;1T(eFF//GVCad./PC^#Sa[RV-RB-XE<d=;VgK@I]#UH
2/X7^cVO:C=&?^XM#<(DVP)?GL(Db(HC+-(FG0A&1A4Ka)Y7?<_&:caY5&D:^F=J
7?()XL?/;#>:JYNW>gDYQDU26GcgW(<U)DeLZ1gJPf(\CLQR&_AECVJ7D4VJ^WV6
8_WVZ=E8HZCcb.)ILD8E94a13&=bH+68]I2KI7A,+Ha3gS,5U/]3-+aK<)5J[PL^
.X0:ONb7L#d-VI.UJA]XIOdD<H/fEb&QC3^[02+@g9I7c1AbX?IRK6S/+/7[:#bU
_8:g5cd.2F:OD^edI)Rf-eV7c#<8cOY<CPe2LgC[;<E[a44gN()E..A..@+/W2XW
>U0].V+=,]66U8PF(#13_Ce=d&A;=6]_WdNH6FK@M-2RWH\V)[2.#F2T+UVH]7J<
YMdG([OIaSPCY<O<C>>f2Z_CMBe1IF8/-7#],8&FdRA[SBcd\-1<2A:@\DJ40a&8
H(+e/b(;NROYN[>JP&A9>#A)._)AfTW]f;BafGcCRY+M>QSJM25?[e^U]0WFITR4
J#Gc2,GDe,8U:7CA=NN9);.R6/eGP6:Icf9,(;-:?5c[0J8BG)[-EUPR93(G.__b
M2W,JV[=fd:G/96\[=GS5;e1:Z)HfP2]+>XW)\.TXV4d(1Gg2Y-GUCf1=)GPVT/Q
\2E2IKRR-8g/EMH>WTA2@XA5Y4ZBS@J\7-TW/R0eF@2[#be-_H8Dd5X_5X6OT,/)
ES,BN4LO0#U#TbUI&(HGS[G3gX7>?,G3O.Q:G#5ZJ3TdL,aWF.DBeY3:[0@3AAN.
VBAA]MU,R.L;JN;P(;>U_ALgED;+&O5&1@R&IQaBRV^NSP,9PC&J=L(ZS@-c)JBA
fK)58<4+:87@B5CJT(d&cQ=&>K;ECKc:/??^c3ZN)8K>b-9Cc_#E5JCZXcP]^:<G
NB^VWJC6.Q2TM^JJfWDJ7J6^=:^0L.DFJEZ?d=<TQG4EaRN+5OQTY:PdDd&=^N>T
^YfIBdHb./)Pc3Y27H)/KV;,M-A247@dF0+gY?ccVT,Pd7@;,>S^FY\@)5]cXRFL
d]F<_M:UK)E2ddG+EA5;N43Z1^7S\V9g)e;,0._NCF0c-CV<5g_(fEC2,;+bgM;_
K30\Z;RaKbYA)WC2VTS8,[^Z4g5,URBCFN4?dd&YIfe3_8gEIN<A0F:D\:/^[H]H
ad]a9>H;B=UB#P9J0J++_bAcENI^U/(=O+dd\().5ZZ,X)2Cb_F,2#/:@6VH3FFK
0_d6UT6P^L)MDZ&BNK6D)A+GE=B[57I3EAd?XJD6\OY/fg9:g9(eOL#1=[FdN29F
Kf:L(@VbPZe;\(gO+5e6KO?eUYc:?=e4]/8A7]GXSga?]+M^OU/I8@OPKC69N^=+
Q:M9<>F58F0&\fY2RXP,8,4;4LY7cZ8&/&=Xe6AJ//ccOC:0WG08N.A6a94fFRdf
K<gG@F,GS\WLE;RADQM8J5\3K1R-V-H<+)HH<]VV.\Q8#-#MDN-SWLU53eU7N#)>
LFWL&aMJCg2Z[I-B_YX5IDZY?+12Dg4P09.QcAC?]WU6=J@WQA--ZS?]8&9>+6(K
a=N_36;BNRV#Mg=,,#[a/9J89Pf8@TCeU&R5YN?cB46M.O?KNTeHQ3+1AYX..AG,
Id9V7+,-ZD&5/bAHDV0:XBg53BT(J,0YD]YR_?7\,1>94Me09.(/8O_JRb\5XRKa
1F-DWTKLDPR>M5aVLRRF6,(56_DP]_1-O;b^I2SIGf4^^9C-K\aV,LI2N<W7Qa)8
Q.GW076QTAf.GY59<[gaVTJgJ#aBYe&)[0^#fVW:Dg,5@]3c-5K-C^-I?@]MaIY-
71^@23XI<1V-S/L_IDHWW_,P_9\O<MASc.6#TK\&g\N1>DX#@;^SbcUf(3P)MKV-
UOf)=GU.1AL<ME6U9g1(RTaDK=99.TD0eM1TZ<WV@92FE7F/\VP_a\Xf+dE15+:V
1d3>)?Gf=8CFF;ZNBQL.Of(;dGAag3J.LBO8F1T?Q>b\;GXQA8aP#Se)CC1I^0<J
-Mc?_=^9TB;L>M3f@7fH/&>YYM.P9<d;#EQW1>(Gf+B[cf4HBgVEFCT/6Lc@>B.;
Vd@3:9_VUAb2;5P?&<B4OPMKLW?M(D,cM75ZRF^DN9(MGQH3ZA&)AG3L_^;bARaL
TgaS3N:>6G6J>\f907FE9+F0eQKWOc->]ASb6gAPT,^GJL\=(Y6]55E&4PX.C@]W
N:?H7G^f5SB24\09TH;)=IEfdL:;c<U/+E=??.0).-__KES.TG6T[:J:]YT]^YVB
=Qb.8cQT<5Ig[9>([V3CQUWBVBf=KB/GQNFX/Xg5/K+FO97.@>X.AdIa.cUV0#Fd
4NFF9_2c@RE.#)1[Td_3(2+A[RYK17Y>,P:a3cgY60OB)_T>HB/Qb5+F.+X[5=_,
Ze?AC7I4aaDAMAY=-9A-;1]Q.,cHab631eR:TcTXI#J[1UZNR[/]d.MbG]J-X(;/
E6<5]Ea+D6XVRYaY\L^R@/\Z[DW363O7FG0M6_0;FI>7U4bb8+])0G=5<=UK5(GV
BaGKcA#^T/2]H7\/\4GGJVQB&?;8+9O2[WQ#B;f:U>YdD5,BY@=>N<4IX4IV19(b
6>X\c])1T..V(>5RRF]K:4_IVJbdUD<^K)cbHb/a6JHcb.]eD7c)fB1GTgQ>6Xb^
I80a[3D+Y8NX6fT@PR5EHMC-,fBVCC.B<1=/Wd\>K,=S_XgTIf/R-#.27GV550Y_
Y=)XZV+U+\X-[gW+,b/aJG5Ua(V\^;6V8@D.7&1M#gbCT]G6MPd;KJV=S8gAZ\2L
7KK:;8Wb&+e+EQ\e[EbY_K.<fg(F-@0V=0@]^,gUUagcWD@V-<GA^YQ]-CK?Tc&e
T7S-HbN0YI2DN?K:e:/A,_F.EV.TD0KHH@3YJL9)UT3<G=#-0BYZ>9.@TT?(DW=[
Wa<3Y>;S8^K/Y./AKNUUXKffTXI\+:I5[3N//a()1Ta+65KUM#9)/E.SP5aE^V1)
Yb)F_g5c;#RR3T?(d70>fHL+a9=e-U(6R8KgUd2<1I?0Q0&2X-TXN;RV[Ve2)#</
bK2Q,U/KT]Lea^EI_C0gXXe/7fW<DOI,ffDeb)O]R:JUK8.-Q@WFPT0O381@4H#7
H):KR5CO0M4c2O#=>)8Q?-F@E3I>;V[99ER/DXf><9^K_J]B?e09R(Hd<17U.Y?F
_MR#P,:0Ed7/]8edYc<B+H(Y(O/aD.,T(]E_^UWR8^B&gD=_Ada<;DeUBMcA+e3W
0NH>eY8Ke;.K;9,#XC=.BDU^Y6R=[?^?gN.A](2O)HPL;<#34Le?+([&@<ScD?/(
O>GTJCe\1=2M_a@DL30d)\3U)Q?Og&6dbDE53XL0Z:bR2OC8#4K+=[0751&cMV4X
1Y3WX?5NadUeHP),VBfS\,QfW(DUA5-OW3.;8L)Hdce6#2@YX((bUB/G4FK8P>05
M#VOg4cKXLNC#1VN>,[e3DBB31@G5a8;LbTR\-J>c24?HZM)^A>LQM4IT[I^_/\N
/9XM(>?Q@2?I^BfVDEUEd)^SeJS_g0B7N?\JKS&,9X>9USI;]&]K7b,BgQNV=[@_
c-H.O(9ScM,UP2O?CNfLSVfL6N0VRF)M\599L(dIX,N.X9C?I9K(X@N3LAR@6,;D
eJd:_@27?(KRH[eBBWX5YZ^c:22=a,?&92.:FA4;X(A)2ELgYYW;/EZ?]D:K-O4G
;GU2-&Z\^JCH@X+f<4f0^N\.I#)VJ0T/M8/.<&XdV]fcWXbZP14;e@18=OO@.gMf
-DW(a(Z=I:)X1Q3_[#9TUcca+DEBY,KZbS\P7)I^9XS<J<OJ85JOfJf#9EcQY9f;
AcbVeUaM9Vcd3W>c=MIZfC[gX?ND5WB<2#:D<@15TZDeb889O&3];=4bK,\Bf4EG
<&PS@B\Z+1+M-+8fJ];O-8Fe]L6,BG[b65LD?LZBG56)4EBEH4VR\IaWLTOB2#?>
W#0EC&Jf)2CHOG?f/F-XPFP.,A>7&OcgP6_60bE5D;A0V#R9c:cV;TJ8<=6CKT?+
X)HZ1)Ng1^DV[5I6,aJ6GL+b,>eg2DT&8YdIO>V@bI<#FQZ,<c1@][F@RK,DU_dL
?XSTY/&X.UZI[IJ0Q#BCI[009eT6?H#1?H5)\=-0V^6F09MW<dK?MJ]2=@KZ5d,5
BSZ_\P>OJ<R=.+(F@7UCE3G,TgNL\4)RXObHbQ\d[RL/&LB@E.(98RC\c.M(C#CU
VDO6SBLTKHPLCb+Uf@@HGUP:++aQ[EdV.0>C>W2@BH&&8X<f8>bXC?=Z5(NZJM#O
5LPHWG\.Ma=IZ\GQEG3#Q1Af89-?fK9,=M1-UY)EU^^5I4O9QL^:O)@C>eXK<eU/
^W.W=.]RT>gBa],W8Q)CR/-?:D[3SAZK8G.4=P4A9f^a@@EG2-?L7[F-\5U/DgQa
:aS7O0XE/<0OCDLR7U3-YSR661R.MZLcG1F.BSE^<7G?JLH-T_UdE/G>R9K(IQAE
f(9g,6ZKJPb/NJA&LI\KCIGd3d(R([I:G?#HJ??8WARB=_.=f;+S\-VGB4-3][D-
N8V[ZfA8,07FL/edIGR0B9#)EcLE\V@(FTVWd&.U4AJQ80.K,,&B47L<D/_1MW5C
&DFSSc@bWAX<DSbO+ec_f\Z>9QQRRPG1PH]DM7J]gDIDd>,#6JLc>S7U,&:[Q?S;
ZBc;K_W6TOF.6B,.J[UERRX8SP;Y;9Ge^g-H-@TZ-P/1b3GUN/3WA/VZQ5)51#\\
61[2Qg,3;>@=Ce2C3fWSHRMRA1Ra+SP?[^M3]S;\/@a0MK1Wgd^eZ08,_0T/&XOD
3;AbIe5Nb2.G:KN),H/M7,C9GPQ/^]faMC=4bG=1]\GVLC2G4SS-Ga[1E9R-C?#M
c>E4V5[X@XWKGV8\\f414,:Y[/4)b(:9eaeJb;b>5;c?3Z=-1]715+c[/?;>9?0?
dd=@,:N<L\G)F0@<Ib]G1#2QB-I93>;F[cLgF^S^NTU41MMc2Zd=@0E./#(fH-G,
+5+>YY6YO4D[IFQHUF,=,;SC?3ZI]>3Q#O;)=A-2]M]RYY5[d;KcG[ZB2PU:Eg9+
^SZOWRLA_BIOc]](HD)eJI+g;MY-.\0ed=J2EV9ed)VaEMP.4&8[F&)EZWX)cJ+@
<G0[A&+<e/XP\C5U_:;a?HG3DXa&CZP7U@,3V[CC((GFD&9+XEC1=KRP1AS,D:3A
_3RF3K>;;Q&?gY&/FSR-]2)^7;=RPd:;?(03O#g-2J?HKfKF5I8,R#(QOVF);A.Z
YN3BY@K-0+Vc+7:eY7ZADB7#J=V3Ge]D65G0e[aOFF.@;5?:a3<FZ9,W?IUTI10G
M9X:B?<:Y_F)b(BUQdfLFJfU-/MGSRW\V#K8^S>+6(+^9O=XSCW[d]/D/5-^ZgG8
NI]f#^cFTT1f-YTSD1D:^9aAcd6[V2@#A]];Dd,E5]Q-AL.#8UbW&-ELNCSKZ]_8
Z:<_+?d8&7OZ+(9WP6XfN,Z..M:E3KaHEH6\_&a#8&_WbG(O^KeMc+ZOeI8D6FC:
FES46Ad.5(?;cLAE8_@ddQ^60X&+4DfQe4X]V1YA:^[Q&f\>]HI^IUc;??IYF]S+
+^D6cM-6f+/HM-^g-=6A,EUC3eEa6S^F1&gZdI#]L@2A&-6SgO,52P0#.a(0NcGK
2a&I<J_<,4#3IO;^C/YU.8^WZCQa0Bf9O?]B:2B.L9XYXDP##(Vc6WNFH1UU=O19
D94NKX+I;I4J]FdIP6/.@(PbL>74dH7UgTVL,Z&_6OM;KId[WT2+KWD1/BMZH.;?
T6:J&S-4N>=8#\WQ[(:7KgX4aU_Xde.QEL,1d2E9C,3Bc@fNBK0PS@/4ZF8ZA^M1
M)\<VaV?ZZNI8?=,c)2f(3A2:4.-f9)I[A8ZBQ@22\\ES2d=6Z3&?D;X,>M_J+VY
(P)XU_1)19dN31gI;F\A8S5P2WS;G4,KD-ffPRAVa_QK0M#>=MeR6;-JHg9cE7eA
HbZ?_4M#<Wa(c/DG.Q6T<(Qg_b/&;DRJ?HSZ/L1QKL:RWW_+<X[@V?9A/)#BXC\A
?WR3[&8Q-C;eS4KR&+CeH45P<G>7I5X_f(;6)Hb7EP)2R()L_-8Y-efP,.<K7Db_
O\\)BgPO8S+RYKN:^M.\[EJB3Z]<2,@/,3RA]RBgKWU\\\[bHW]cBU_RNB]-[T@.
J7RI6DR87+H-RXeOdDc)/94=GSE(Q,SHO5W?]^69\)_Y;4O;BgJVa=IQF3JJ4LH4
b@5/_@a/PcX?\4G\B+&f>>X=FRLAJ_e97bT)Mg#\QIH5b6KGUbNU.QJ9a:c:[c_a
:5Fa:9f.A6g[O/;Y[7SAG_ONMb-QD4ef2?@Q/#O/[WHR?BRcXcPgTICCESMRQ&I[
OOC&@gbV:B],S][BTdJfK[[4W8?ZI,a88>#WJ;5_Md)+99Zb@faC(A@G((779D11
be&<^BY,2MF:/-YcFHc:G9P<->F4+MZFJ8OO#T\E4@+EQU=JA2L.^^McS-#T@U_a
>^]b/LcM^(EJ>UX)CSO/,UDWEGI=TfYH?.1:(CaA4L5WQN21d):V4DOQe&#+0VUJ
6IA+RegRTRg+X&W@FUXCPB-;)^_2>\&ZR7eTO.>f.-813F)QV61APS361ZON-[c]
>RQ8dW5L;2>;6JF5YWGZJ4E(0(PNaM7\+S9/&#R\STYXZQL?\_5Z8-7g8_3XDRDX
9B8BEdCEVWEGNdG0+<Q(f9bg,X90:HbO61&B\2GfR?D/\-eb7F3SYe3]RDQAbeIA
KLVZ->HSO-fZ_:Meg#GK&I]e+>7XE64DT8:dB_0-DNd/aWfFbLCF^L97bGg:f#3M
4#eP&=B]3RU:^59LSe4\93f[C/HcQ/3NZ/27K.DK<Qc#<VWBOSCV9RgP_R:c(S,;
>EbD=6JQgX0#YA=REI9ScZ/<^bJ591ALJCN;aQBAP_PE(U+S=\E4:[N9:I-]PcCA
)+.B1QIg0[#YIX(,e(#BFXGOF8NZFe]NT;])DUWC(+61b9d.#\aRB+a/,f66LN>:
EE5XTbfIB[P\?,[COILAZaKF>0dQ>e=Q1BZM0S29OV19cV#Peg8g3Re=[bQc,DG7
AA?DRdT_+CEU.6_NW8?)K3bed=O&6W@>D_d^3YTIE>ZV:/,3#Re]a3C2AY9I/G0b
P<@>Xc9Q_Kc9GDX@3@[MMX3Q<R5L&;Z><Xb=<YfM&g&X5\UMW2/HAI#AX[M:G,,f
W69+D:R@:I);2WJ?6]@;TU[4CM]M;LRN:<=g12@M&<P+3fI[b30J_:R6W>UW.XF]
c/PZ(8:T7PaTgM(5d2-fHE4DT#dDa,:RDIJ:2:U)gbNI+EQ96,:NHG58NSG?d[fc
OR]f3H23BOM0>b&d]Tc^86Ce05AIZ&93Q67Ea#?b<Ee:H3\b;5ATP&2\M^>(a@Qb
5C2?5\F7D46G6^>K#/A9F-cO,EHIG++>XB=[2=AWOB,1<ME0KD1(5gc?A[EG@A]^
A[/W&&f^GcTaMY:3K@S:U[?]g>X\M0W@7#ac)EC(/Kd@Ad]W=La/UFR]ZaZ,/1eT
I-PX9A=C/)5TN<K1T4HL(8VB2bg.&93X2,PQ3P4.>2<f\Afd-BbQLYB-:OWVV0(+
FCRc3Q@E2M>g3:^+/+(c(,U^eT429F(W^70MUf^@G^P\D/PXK8T739NfaF1=\FUA
cB0/-<3)6N_Y6\WFfBH@8_,1NY3CFTd>((58/Y7G<4+R@I#06D,g29+,HZOQP>T^
:U(ZENQC@0@beN_J@HKNY6T8S#CbM7^b-aa<5/ZIfbHR6TT0(,dNKNRNZ[(V?E#-
T88/HO]SA?R@\&&72,J@-/YQ0\=T;gc2TK0<D/-bT1#\EWa4:B81UFH18T:A:Z92
FW?Hd=fNM2&e8Hcd_@8C=,K3#ee0/U6WUYX.eB/?<PPX)DQ&W1&:L\>Ic+EG@+bb
>?B;d8Q,bADXA>6^X?2QcMI[NAD6R=J_.5/GcA5Y=D7aZPRXP<85.E04O<\[Y:[g
81,?1-IOS5:W)[a?QF4YCR)9.Bg-MT839A;D^XbGJ.cL2fIL\X1U[VM2Se=Ya\[R
MEJ)XFZMd9AA--/FE,^MR:K03W5\^aID5OEW@b70<Y670(G2)@8:2c(PKd/=7&c?
LL<Y4T(/c.&I+^?ageaO]2_).CFFRDQ;e)#43FC615K,I0d19L.dFO_<29-bC@W^
1,@gKJ[G.<Q\;&A2P.DASVK[OF_7U.FXO2@PF)2b[+?I;a?P=1A\E3+NR=A3R35\
e942S62T)eWR1W=SZ@dI17FF9:0K+;5/X8RL_[WBMZ?EV7L&(,9T\=eN\O=J0PKA
Bc12)C.JB:W0TV=O?453--I7<:;.6L[P.2X7@Y_EARM[O3)@37;K0;fb3Q25TWR+
4+<EF/E48Se8I+SbK])2gIg>&BF[W3[=DC3>7<@J#DI6,@D]&192Idc@R8.KT),_
Z/0e3F(\C^?]f<^eEeAAVe^49JaH0RYM+K<+C]d2?T&a-[\N;Uf5O16#4A2/&94,
2#IWW\6_/?d67.;+]CEW(PS1\QCLc]@K@b(&1,@.d?/ZaG#Fd?J6XGBId#^O?6ff
5V,^Xc0a(+JBWF/,R8X[M[5;]7J39YcD=VRBJSbJdUgO:Uf[8+AQ2C+&IX>9;_PJ
(A&M4T)R0:.DH>T3fT:b^L1UJBDASeOJ5gO\DOI1)g&gD_=Z0^67_1ef8G_D42H@
54f./,E2+Qb\_0E-]4U3]d=]aYYV)229(N2:M1M<^V(OWYWO?f^;(08NOVPAZ3EZ
M>Wb7:,]N8W_LfD=:84X08O)8BDYB25U+d[b_.Y7D?;Q](C7gA=AYT(Y;59J_Efa
S#b@?M[8G&:JdHSa8Nb(KLLC:OcJ#:::Z1FK1a)+88?(TY5R@68IP\.SL#c<=(:F
,6Be7Z9VOY:&Kg.RGVBUeO1^+Ng<6-Y9[<M2XP(K==HN:I^(.93F<UJV[^/TRV,=
U),A\E.Yb_YC3Y=]27XOA3<)b&?)_IQ&P.25)U,D+4E7SgS[;[X&DZC0&?:dc6Z&
&,4O-X1O#(NFOOLa,BRZ9JWe&?a+fUG#6S.);I.S=E@PB8XN)H?F9@<76Xf17DE1
YLc>2MF:+DbR&TgVK>e<(2EFeKEU;?F:^2a15Uc\,T=D0JFdD+fNSKBDc56#YE7Q
^C6DSPdBFd,,E^[e&6-?b+-d_GHg\\+HJ22gWQ824+=2N@^(SW4PfBcU9F;]2a,2
DgC:V[[)0AZX/6.XG@).O73),6HJOc]\6aHe,_8UAKB4E,-[#N>U\^DSI7Yc]J1T
DCZ=V-fb<Q>12L^(72EM+6(@\VaW4;@Q@9Jc<-E/W905GT3AKMPZO&3,M;O)R(gC
+35Q@=Eg1)P-C3@)6UU#M487/IB5&BXff)C0e9PDRIJgbY#>bI1aNF<g6.3BH18[
TX@J/QT\7]QR>ET=Z8Y7B#K-5-0cA-da.La(+WXO(IJV6Sf-f:Z-_X5T-.JTTf7L
]W5gYG#W+]?cT8/@_^^[3:97-_3_T4_C7FF;+Z@0K([;Z18T>dS<Z2AW&VK-g/PG
K_gKII]\+ZN9?86a/:<g396cTS?S>Z9b+DN3_/#VcBeb^V:H?0Ea:8)B_A#H&#8_
0RQCR>;^\aNWKb,&1F[.P-?0-NWZa.9-g)).c;d=d&ZR9MXVHX-2F94KP7fHJB(8
]fS6V\gF]BK6IeCT779(H;RHCBAegb/WX:#XZTM?]WO6NA@[Y.&YBKLFS3/QJQ&_
S]CeV,aPJBVTKLEcIJ([C[UYSHPdR2<WT<Cd>d4CGcfI@?2I81>9Ud<GL?0cPJUW
Ea;N@M;MT8A^<C;+0X;IGIaA&>S1-JO5WI>+<[>H2<5g(HCTZI39Vf&=@-^AT9/&
R4X&.DDSOJ39J#R-)ID5_AgKL3<7P[FODWCJ6Y3V?_PL@;2d.Zg&cB/;RU=+(E-C
A=N/9b8bBcR4GgD+X9W)]ATfL=dQg/FQF&&4I)1)_cDdM##aC4LO/#MB1(NY9FD8
EaDV/102)[aR4Z^dWe.S;T=+Z6X]<FgQA2T3(R.R(WEWHKIJ..-#gQ826-35;=SU
11fA#37SJ/&3[cEFQ#\QICI2OFQN9GeRd_QVS-:<K)>>X(5c-F.TK[b&Q=9LcJeW
CQ<M]3JfE#;(]NEVCS\NJ+Sb15WDcC=F)gPWL9I=4#A&PJ&Z6#Vda;g^),c.Ae=4
-;9OX3c/\ed3Q#A1=WW<?a+bYXFBTGbe/B=,T/?9<@H9+N5f?H9IR39.-/C6WP6B
,#&A(YKJ2^,dUg:]BfR.<>9]&9NQ4:@D+U[G97WA#0];-3IM9_\DL)TIY])DI8?]
[FXf2+I5,D0I:>gF0FR6OdDE;PgK)e#XGE_5]#&CXF?&eAd<P#X&cgMNDHA1>b)S
1\,cdZG./G#-N)KRQ3A,M<a95Vb75-S/3UGA;[<>RX65e#=a=33)#bQ0bb=Te:T?
cSNdLG2ZD0HI6LHJE?N@R0Xc_B<J.&3-2785/H]\JAOM+@V9=THY:POZN[Dd0&Y=
(QT-L@&.,aE80)cHS=N=[:F4X0]fX/^_Y.KP-N[2&3gbLaPaS?+HP1ab(-:<+4[U
aHLP3RSad=@:4),U+M,\N:LY:IN-M#OGg+a,&=gg1#OB#].V4IPADS/d,>^13a4.
]<3+#Kf89Z2ZB)H0.9?EbVQ36P7WD&8]2K9+HA8BGfJU?PU4&N3=7PR)5TffJX5S
/7X(>:O1\YOg=GV\?7\6-_=&17->b\JdMD9O7?DFI]P+)@_O;\YcV7dS,[:bB6J;
Lf4D4>b@94:@Oa[TY0[c>dKR?R>C=IP4LOU-7DLQe@6YRbK78-8S&/E46#NF3J<K
\-,P]7U=W#EeP^CHE.E\TID_e\,dT;XN&<EZ=T\>7.4cP4(6SV)NR@&^b)eC=FF[
T<18&8;>1W+dL)4CYOE>?P3>J5J(ZMO8A13SBQ]E6-O6\@_B,^X53:Y7-:T;Lb_5
f^bb=&L/14c3<CA[44EdAac<<@=TT,,WR5-<Q45Ag\BU(JMWd_ABZEN081)M(ddY
5:+(\QN)#e-R4/SFK&/0<-5;4Y,G8WaS:5O_;_LRH@YgQ(L-]N)VQTAH;OUdZTC8
6&))8fBd#(QR)(fH0YI#\KH?f&V-FXB;;eBd=J5SYN0&\ES&P_VNI5(TD<-B98cS
H8Y5XLKV-R]EL)_(KH1LDW?^1@:7_L2H;HIW#-J90fSbT6=Z[73AUf?A-Y@3X6QD
JT?;N=&eE;-O9=LL6\OZPXTcWd26cU/U=M5d>e@?CRYeV7AKWVRWZ)>5KB27SDHU
+TL[E?.]fHbO4G:?#>J=gI:BDFL/g4>^HD\TTHeDNF/B]aWHc2O&EYGRUHWSI<<S
R>FMYZDY?TEW:JC&\-I+Y^BI4(,5:.YbU6)TT0#SaFHTW[6&,b0;6D4O>#^94.4/
[=U4IegV_L@^2;D\e2/I5^:aI-4^eCK<Q9.HL]#W[J:#2b-XaXBZRCE=Z<J_@_I)
PYJ<<6X_NQHH-_K7<(:/]0-]JRF>QDJ)?)(5-Q[+=^cV6gG[1B57Jc^gb15)abOG
MC^=YcW<UUOcP;\ECZ<g7Vc6HC-,V;)Y4:OB460=e6=)\(HD<58_1Z7[\LXc/b;Y
e&a_MIXDOVZXBDA#>b<J.)KHT,MRGE2/.dc9:INQCF.Q^9c+]--QM_V@1NZ#_RGS
+ga_g_3X8A?BR>RVbA;5;NQ09:R1[[4ZZ@:/GCbS:UH?C#bK6BFJ=LA1<[&,&4#0
4U,/Ue0-A7\Fc^1W87W?aE^/gJJ6M]S&#PS8@137>ZXIK,.K)&OMWIRY,gF8FX,1
RARZZ]-e+bfXV3Q2EWcf_SK77AgA531V,CP6A57:AB#4F-1688E]0bKbfR<eM9Z+
=I.[eH^gHATC,1?<N:WR.86S[6g2fCETKEE?Y9-[LN58R[L3<09_B#SC6deAbC._
7Dd,/S0I-;R]J)K<63Qbd0R>T\&S-2RZafUQ3PCX/2X94VFaGP^]INUAKg)QS@B/
HY;[ReZ_.>_76K(9,AgN[4,TFQMbQQA@<LA@/55e5M>\(,a0dg3P8-JDT7;.@VY>
@XYGU<Z<Ee?Lc2-L>LV<C7Pa#KDTDA;C,0,9TR=_QDMcf64=a#G:dT?ZRP>Xe^(2
\5ILDYE3_.M2dBN/R1E8<J[E9J5A?:+_H4.407Se0W2K^Db9@g#B=EZPEQ?Y(.bZ
TM7=3/\(:]7BJO=\CSWJ.1c8GZWW^L,\R,_Lf4G1\8?f,//ZFJ-@::[PCSIHTF8Z
=dHBE;fG#FUAT,SeA@8BIeN.]<6O6LDV2A:D&H(bL=2RfQ@8LPJ;;/==+Bd0(e7d
J>6-5H[?b-SQaLX(eU70aZW5@&V7;,0+CX)F.gM4;P?D//b.eDY]Z,RW>I=3::P0
Cf)<T]=_cTV\)?DG=bC_f9;-AI+<7D2C4=#8N.7e5;]+D&b:Y9A_L9UJ8M7N&[7Q
OSK^3[?++N<+[.a8=+>D>MdeJPPB3\,HG+SO#g?_[0@e4>/+-ff^1/NO&:.MT53a
GcV9_6aU@S-;H:gNP/H5VRgS3W;/3>F8Rg_;OBR6+NV+g2N,@U+#XO:8Fc3/C#N-
bR#88[OQ_]_Y,:]12F8@+(dBHV0/>bGO/U7ePWBQBQ::5XNED]<A;UZRGOb>4EM3
^K=_S:@ULH)))N]HKff6;2a2GM@[IV_0Sg+S0N4UQJ,A3V<K+4g_&OY3L07dF\W?
P[a_I+HL&\(&9W7W75LX-FUeM=YI(-HTWHBPI]QV;OPZ_@Ea[^0PfVHX9S:d:ASE
N3\>HW4M5VgN3#AMISd:GY?P@G?O9dD@L)UK?0DOf[-cOC4U:>SX/\g5GIVD20SD
ZR2U][=O?=V0KE_(2J.b9Q9GV[-(R_AV6\L3Wf_&JLK&Z+YMG8VI]BS73,^=BVA2
Bc(:=)VM3Of\B8VaAKI&HE<N[94O,]ga&L)-V;_b:@G]N[<M5W&g4=]gd1Ia]HR=
&bc&#bFD[Q&Z_(UV-1K2bL<V(]0MEJ<?A60&bS?@IA;e_OeI)<1W4\5\fU@AUSB6
[aI]90:9LcD893JD@T:,TIGIcMHO\;@U&;LBKYQWU5I=QbJ1Z1_fQSWL\gbC0AbB
;@Y[Zb?+?CS12_^DM?51g\T9d@g;:&+IGH+3cI1aWW:fZ3XM5_EMBOd#:JUI2C#a
fX,Y<>@6^eOcT&g:NNZH3?_>dQ+eKTcGR)W-T@OPYT^C:5/>a+Nf:[CIO>;;<OAW
\b8eT9TW^8HFM9Id]7WF.T8b)\cgGWP7BM@ZSE\?HM5-)7Ud01HMB=]@<0IKURCc
_U6C9<]b3(a>A8F39VET&5RaS]+,1[>1gAI3&H,B8\\P4,#^[CHMF5[cHLQ6-,66
D\:L28))1>FJH:cVM8Fc>\fc&MeX0D\;GYa;N21e42M5=;Ngb_gc>)=Nc_4^.1>-
T_+TYc?<W19;/T9QL)RRJBB]e;U_gDSQKD2,(UKTO[70YV3K44HD1E\L0UH#HF6H
JYT)5+U6LJ2?J)EV;E1L8XG7+KHTa<_&@V@+=dYHRdFUF.BMg5-&;9XBPCF_.Rb(
cUcP;0T[U5S0EK.NaAP-e(7g&,7C^;:eV3d;MaeI5-9;cJ0]JbdgTZ9I0BB3-a_6
@6-_@ZLEBI(BFX_Oe61I=98dU1RQ=3];4YKN41C5=Y38&?N28faV:2C3Ga#8)1QW
J?RJ^1\#@:1e(?C@bK1USScF7c_/)[_bPJMO14c-U\Oa7Y]\V8b+?4?d:0F.#^YF
TgU;]OC(YG>[#<R&5-532)#U=/27geO6C+.B=W:\67N[>=:.83,TW?D4>V/U@QdO
+<_d3IAP#X4>P5MJ27A#9)L?9bGA3=Rg8-.3EY(2UJ[bT\T&CIPfb)+bUXECQR_.
+5C(-9RU3A1T8AdA-:0U(NXdRRN&8Z\1OCcY53,YGLf,DbOe\TO>R)2bSZ_KR6JX
L0RFGdR-^^K6>\JLM9+_gS/)I2Qb9?S=#6+OH+TK&-V7KTQE&[fO11:U2^Y\7:AS
A\JPI<W2/L0d(HWbM<:FN9eI?#D3SD2/\XAgU>#O7XW/0<;7BgMRM.GgCfZMS=&>
e3VJ:9Y8A8-Y-+8H.0/@;fY^@-TCMXS7@(U/EfZa2L7UV[.7[]/1+_<<_N7)<3dN
SZfNOCNa>VbMaH)7]TH_;\)<:6Id.TaW,2FZ=BM;[e?,H&aAT+B[AEe[J@0/=(DI
:0L=L?>6X<7LafNYC#<D#N?;TSVHZWbO_PaOYb.)Fg)(?aKAHA705d7Bc\>eRK&b
g):2a5-b.F7eY;6;ICAgP7EH[(>C-.T>GU)LA05+:[4Md>LXZI?\U9&KfcL2190&
aRMb)cH@@AZ^HJA:;/f.<fG#3@\V>cW<G5#Ha.c2I6bK/B:2B.MRA;4G#/-A3])B
:&.Z>SN0d?NIRKN)O.T3PBRe7&N6.B[LccI,/H1fE_)A[SaY\5cN3K79]L#I]J/P
)#HEe903:K>?S[=Y<PTL;?W9,gbbJIN,G;A@U/I:=.<BBOZL:9ZT9A_eJ4GJQYDF
VZ0adb<6]F]1d1:OX_PR;2_2M6:PJ-.e<=+W^XBc:)JJ^-^ZWb32V:gF8.7;8e4e
^-Pa:7D7ZI;4]/BA9IcDVH3-77#Wb/[UEJYOL;O87c5X#YV:Z<BGKDfVB50#?#4U
,=Za7;IAZb;V-f^Y8-UW?Q-A0;[->8E3@9W)XPfeGTYGAN>28CNOEI;Y;J[6,b@R
F29:J]XMR>QN<+:d<S,GBLC071TbEM#D.FLWG=C:&[;X(KXg:3<gL2H2>L#I7;4\
^T^c8eeH?CTHW<A?<@Zg\>R+;Hc5FD)+W]I87.PLQ[?/050=f+?[M7OU^NFf.?-N
\V:cW8N(PG.aNfM:OcACJUXQS5U4VSf,WT_2_W/6V\M?JN\V-07:A_XfM\?;\X^;
><_FU1bBZF:V>_YA-BLPZK-YNEN/QTCE:QK7H><V4Pcd2J17DZX.<_?IDA=Fb<-]
PDbD\Q5+,U(d@VRYQ/L8fJ7.#G:Q;O?K^bVM?f,f^Uf&:/UNF-MN5>=9:Z(O<]6[
]M73R7^-283=87EBcaWb?ZKT#Y11C5fc@Q-aT-]UM5P8R(Dc;VR/P^bee+>4RBHU
CX1g6=+VGHg7Wd_\-AVT&?^9-(\[X^Q_O04cge7HF.XO=I2;#QaaM&b:0768/&f?
6^;AVa[SVR]&N^F:A4beX>+[^6V^ZU2W@=C5IS#?2R8?O0#VFS^6aE221Z@.XATB
-YEU2OVCRKC-:0>#VUZJK)996CeP^,g<;W4SK>03^S-5+ga)I-e3K8\_>A,dUF,W
P8MYb^7JaZ_Xdg.G(bN<:9XSb,>XCdbSC.JK6XJ<b09McS\ZIC3\L^6+=:=W+:Y3
W62UI:14b7<&\APJ>3gBLU\A9]&U5,_a[2T>.7L&TR(W&OYG&/J\?^KV>b3FD9GC
]d5&H0g5G+&9_LX=_QJ:[F9I@U2aG:]cZJK.AR<S,Z^MD5H03;(J+E-ANR@F(VAf
VKI4-??E_aOS-@Y4#Q[/=2]SY:V,@(6bTY-X\PcYKac@P:HK/O7(5#0]RBNBUPHa
a&FZ,]aVeJ.18M(PRHf,4@c_N+VO46PONf7@CJBYdgBDU7DI6U\FA)8>&gP2\TOU
AT>##N81H)THGga7A21H_N]Va@T&<I>H4V-63g.@6Ua-RW>??@=ZQ2NdD1)eH>.D
SgXT7A24?=D7fXZcYL.d[+^H6)/9]UcYNS27PN4Z?05fG_Pf8FQZ63e[^:\X()=,
_&U97GF:/K@6QO2aPHJfZ5bTQFV/N/@P.?a?0G^=,WXe4LC2g+;a?S8-\bbLOSSK
V>(6;&4O9S7OJ^;FEG]WT.JF9aZ([E1ST9>AW;AV9&Q1DFXL]\QD#,J#\0,dcLfa
b#f&7OGfg\L>/[CbbG4N>#KLc-0R1<_N6:eVG&]KKVe0LP<eJAMc#K769FSK1UP,
@XCOH0T?Dg9,9(.4Y@N=fJ0D^b<TKAedWC-]Gb7Q3JJcQN.d]Zef(OM@LSUdK32Y
B&:-)3.HI>RBI)KQ[edJ,d9#=^-@]0Qc1#=gg4\7Pg<OD:d[5O6:^c:<1bcdN[@e
;:4c9YZF0CRb^?5T.#JYT<G.52I+_A+G\OHdA5J)@WMC(cEHHc]H86f_eE6&R3UV
BJbS@e8D&Ia(A.AS3Qb=15XM&;>GU/;+B6=9;,E)Kc26-OCcfD=f:2_NH+fBET/K
#F&C^L_Sd?[cWZ<\746a+L#?-T^AUBR^HGUf7<41,_^CTT@BUW7Jf]KF3;9((e/P
LN.\#f-&R)_F^cH-RE=,f0b5/d52?+QaT::<RScJ5PY0V-\>\]VQefE9]D#K9A)D
.IP>S>=NH3_W;5\S/H6H#8c#+DG@NLJ(Z\^e+Z-:B?U5gE+JJJAR<JETA_/W9d8&
N[._baVO:U6,<8<_ea_YGDgKNfZ>3g4:Z_^a-9T5cd6_COURFOH+2RY7:BB:PHT(
\]RM@BES+BXJO@73#\Z,V.52@-5P8(I&0Q,B&>Mc]<(>7:3^c+DeK?eIG66/YfZN
FHEK#PTM:W/ZR5V7TdcJ[S6>3SP9fYN15R<a]YIC3UWeJ@,c[L<UWK&dON:A<X6&
?.4RE.:]EZTg/ODV188ALWFCY-E4=:NZcV_QHS\[<X0N&N_YYf].PRM:_,>-e&K^
.Ld7]aDfAd>/5?4CPGOR?^HT3e.\MTNbMb[:bZG_Med24=^dB>3_4A;H&C,,58NR
5?C=M&ZHGbO4;BTQ6>-\^8=0Z28>EfZcY//V=Q:WdPRB\5:8RE:g,0)6e1fLD>M]
[YR2/)\YQR(=FXLRQb<QN:3K6.^:aD([>c-gEPgJG6>4RScEbUYK@L>YE.A+\.CX
NL,A5MK#B7T#ee1fa]/D7N6>g@aE/P^:.Z1XVQ<IRQKb-2.)[Q06\?.;5Y<1+/#d
6_YIG,963Q=6Sb(CIT_<@Cd2+7a+=bLeU5SG,RYNb6UU683]Z?K0\(^cfVeX]IH(
;2QJeF-AWfJL:.He:Q<KI&(a3&^OG/19V,/O#3E8YSN>PdT7A929EIT;Q#NbSb:,
ECPO.8I(9;?5J=&SK2Na4\\U9HeXg>VP?\4\]9a#;GLK:1OAfCO&M\06B//LeZab
;Ua)O^f<TQGfT7M#B^_?[GI#9.&=Z:J0\?;^#\S>T^K68&LN,dV4eVAcRg;RaJ[G
_#<>03/A:KFbC68-Bg,XZ2M<WAD8fa(\U@2c#e2M:#1HIQD>C/:5eW:dbOb3D)dZ
PI_HCdUb7.JH;1436^1A2:V6BSE[R:G+;L1McLG,@.,0FBDCaHBBEcOJU&#5.R_0
7E2&4[?[84Z/N\0/::[EWgW0a0f,W]RbIIF(\gAV:,5UB,3DcHMZCd[XNb>(?M\D
KY#DaTdg.QNVX14@WZG]gGAQQbG3(g&9@#@NRFa9E8N?gSXD,L-5c#/DeGa0dJ9>
QReI7bL]]PcDa_KQ/P&O&8.R/U)bE2_Y9Z>=.3^C#@B&RBN7N_HY1fe=bLa?DIZI
?#bY2+;#[_:FFA]0ecE(1^?C1bV[a3b6UGH?^LI.].DdUc,0?L=A>6QD4e8gFQ/Q
FTaF7JLX3C\HU6BI-d;Sc,?OG.&O=aGX)ERBSFOBZ-YfPDg?[YX_][WYHW,/H2/G
acB,_OLRNfPa&9g)XNaETW3]aXPeDCJV(=P>OeNDf=WN)YbK+/;MdL=5[:,_=fc@
+G#)R79(1X+8Tf:+GN]=?:R];;7G1O8XMV6E62?QM2?d+4g(E,L3SK[a+\T#4@-:
aPA[J<BPeYKcR7+H:-f4V1A+1ZXHcTSP8(6_@+L<Of[EVTgLPdbU6DPNET/E2#W@
@^L,G/UI-T3#K43LfA(?:\VM/>5:B#(_OB/T\7A0I:NgO:P7Q0<R<YIG[UKP1]3A
eHF<aB>C/+F3DdNB1M(@\@CWJc\>eD65g51K3_6VS&&b@>/.=YPB)H5HK\L5KK.Z
B^FLIN,D]@eF+fH@CX9#SL\?Lb/CY:7?Y9&.fH02\b0fB\F>ag4:#JAZ)BC:@OZW
I=.=<]c-6A25fVa3,)GAL+.FEU>KY0U0D+QL5T04QOA8aKAWa?;:MEK.QI@;LOTH
<K/VK[0GbAU(@-PYBBAMIWKAdUf,0d5@a(ZHUbHF1;97gRKd:GZT,#(,NaTCF9G]
RTd4dWS>1Y^LOf=J8?MLW@^PP#+>_K-25bFJc(Y?1P-8e(:OJ(-=ab+ABIc^2ZTD
?92KS@d\XD)f_g60M\GIa>__YS3.Y&JQgTJH4FAX(;L\A<)U(=<eV=0/-cNX-HBF
aROJa_V<.AbbC.3EY0QbR801,bO5Ma<HD/d^YYJFJ<e+G)MdJTLT:T>-ND^URNaF
>4YO(J15&7^]b=)UPa2)I5507a_f+GBM)HLf6^d8Z/)?3gE2(=,Ia6S;dA6@aP=X
f2X7;d1(VgCW^b,8)VY1ANP+#5R)/1/g9A2Eg6>98e+()421##-W3DC;M;_bP#@V
]FXCd)D#X\>7/U#>PU/YLN9C^?]X&GYWO\M/@0cQD8adQ9/>R[MT5O>V:/=Vd<ZE
ad&5[@+_Sd)H8b+M-&<,^T39XTU_TSSFeAW+=d3PA9MF2A7A)[_9,-A::\URS]C[
\8D=]7?IO&BA,b4eb@Q68W>Xea3RI,D#HY2]IHZ6D&(K;<;SR^Q7G([,_)]-<Yf_
I(R]BBXOB]A89Z4R(I?<4O@HF3Y-e9S5BG2+KaTA]:R>S3Za8C:,>EM46<Te1?>c
__875)?b[Q[Hf@U=4H[2J5V_]CR<d2,I[?;YM=85E)fU<;7KW\,KN@Q9fW,HMBdB
9^-Z=D1<L9F&Jb.-OH7:@&:De=BZP90g=^R/I=32=4(@4=.b105?4SgE46).^P.J
8#TGG61W[c9,cI>HR@_A:g+=\Re4J>[N03cG2CD?Z80XTT]>7eSSPQ[\e;e@f][7
?83V>,NYDb<ARf+ZO]e+a6D&.=Z=[HDUaK=3M]Y,09WK=E1>_SD/a7T1[?:04G-e
>B?:TA:[\+a8R/@0(7^J[^OTOY=6g1cDd.^KJAd[F,\/B[Q\H:>;C\/?.7)d+(:-
]L=-G1&^aQ<OWJSZ(+QF(W^PUO;KTB[FbYM6SCUMS/AS,<:>NH&0+29=))X3C1:O
_^T_-Afb<=]=6ZCdQ)/T>7gU\_LRJN[(L92S<cJe)\PRWL^7Y:K7P#7I5;c#+845
R9b0?<3=A<H-A38]_-XIC74Lg_5&cHS#eN+TV2@a)TYI/LS_0QgL68TgJ0[AQ@+W
8)Tcc;-=TW@6VAIO8<(,]\Ye9C^K&<gD4X::ADH6WAa(L]TLLEbOcRZdCf?f2cMH
f2H<)(?VAE\G+EcU_ZJ-a3YaKSUXR,2Y^39(W#UXC>A9.XH_ZH?TH2@ZB5f+bOE9
QOC+K&[S(9_?S70>;Jc&36O+78Fd2f?cG[GQ#LCeA-TAZ=D4ELd&:97gX\;,_McM
@@_<P+7)#35V7+b(d5aOd=&FYBR>U+BJIYSKCIN1A3e5UF+Z4?F<g-1c\S&1KIDP
<T]ZR^.PRA-49?Ff.65.Kb&A?S^(@_Ng3Oe)1E6WC(UTUOU[)dL)B3d8=6KFF7OC
c[85M)T#\3C4SV3W4DX:89#\6N)(;_[YFDd+b_7(X;SQMR.7<-L_Z(82DM0+K@(V
N<DdO9M0464O;HH0HL_<-d.@8WY:76L^GS]_]\T(.e-J<fYVd1#N4Dd<[4[g9V0#
Q(cWT5#c53f<DVB@I:f5)(C_9YW:H]a;##E1U2A?J>4,[bKcVf3@V+H(_b<E(&#^
cRV)>aW6,4CGDF_+NX5K1,DP+6_a/[_5R[-=K[5--/N,6?(cT)ZQ3,O?ZaaT;AGC
TE>QR47&YJ=#GOKG=TdK5QPg1c_/YX(LJ9gV,B<G/S^C#SYWE.>R)SaK96&_?C3.
RID14Uc-GKA1@<3[QC.5,B+P/=?BHg<YA,fa:gfgeJ)]-X^\>C)B+S)]DS3e0SE;
6FYPV#HNZ<SE.3^:VW6JBM@Z-4S/R3?^Z0_B7bM+b.B4/YR[dH#<bQVLePe=0^M>
)Z\90=0d9\WI7M30DG6L@JeYBIM##cMfO]@8D5E2?-9Q9Q)5#MX\/AA<OY2b2P,D
2HS3cKW2WO;@LSZH=Sa:a:]YC#>5O^5G.C]E/LLY8AI/KNK1,JEBCA(5&:\+CU<I
eYD4SEb6BfC7N=H3PT>X4:.:M8eALeD0Z=ZFR?)==B[UVD][a4C3J/IG6EPT6))<
=ZPRKD&C3Z=e1UV?+G_^8\gea-T5@-PJR_V)Q=#)RZ-A:5Rd3?C(/J=+VQONMG+N
?S@?&g8K[Fc:Ab(R2Q585I.)UMaNYM+Rb\IO)<M#]\#W\JR.=1D\.2@+0A3fIV-@
@Q3S)=&ag\,(@N7>N;gdCZ-B6bP)JR8gI8Ld<^Jg:9>UB,KKKd-;OJ,Hg::^O-(+
I[YD7+?+S1,>Oe,g+L1g1GK/?PT_-D_OM@2/TV+:Z#5QJ?_VNOAc79UC)W(0L:P+
H3g=f9YW-N0-#YOV+]OI2Rd@_KB[9YWf.NUV/e_6b[]a+L8Q<aFC2abg_:-GMW7G
#5;;M/CSY^Kf5U14&e2SHFKMR6L3/>M5J^fUF<A_L2WN@Le,76(8L)3RPEAHf[5D
BUbR1G2:>?5eLJ/NXDB)P_MM4VWa,5K_4+7XKASROELFB3&f<W=8dTf&K)1Ge?EF
)?b>@5H<&10e@_^[0.<>L^.:(TR;B5WQG2d\M9)VZ#eaWc#T-<(Q/2L6\F^cD(.Q
8gD]/9D[U<=A,,[W>IS>8-FbW@IQ37Ge&+=U,3A>H.Z3Y:2A_,<3agXZ_+C]TBT/
7P1RREP)(gEGOI\EF)d85;U))<Va_IA[K_2b@2E(c1MZ>aX)\)d)K_F-?02?@BML
J]0cU<;[1\gH?-;)<6c7BYW[e^3UO^6D40[W,&1UCG[?c92SB7F24-:=]9c&Ng-Z
[Qa9\:<4QJYG\=5_f53)_B&Qf[/;U&9]])>Je.PRM00B-[D(60cY3XLS?(R4aR9D
=M47>?>]4P)K4]f]T)Z0L3)-\EdVM,dKO@XQNXST?#H96)J\&9X5GTJ<G+5_\=VB
_OLZcFFQTN8]#8(4D[@SaNRU&#2RY\5[S(=DLJ@<<NLF=/5N4WD<1.#@JCOAHM&K
7^aMF#OG3fgCU_\a0?&\GRY4]B]@BJ;#<U09Pe0F>G0Pd\AbL;ZUd;8.]cGEI=cg
\N.&K&(WVSXJWCF7#eV^FXM:?Z6AeDa0B4GLC;CS\>1UW\Q.F-,0]HG3),8d.,gf
C]dZgce<&QDg<da^QgAI2CG\T:Jc.^,_Q42ccT#PE<:D];5S.UL=6WbVdR@0LDS8
74Pg,TPF8O)GBb>,>&OY\O,aZ(340?ffK@?ZR<;Bd?6BA?E8ca&/)W8XQg_]RN-4
@39OVN96:M[04W?V92=Z>OA(_g0U4;.<a)eTRc(fOAc(g&[U&BX)Bg)6TZK,((UX
RHIJNPH36@bHR>F7/>dJ?(UNg)QXfT5P?)[6KGWIQdP8Ugdd)/?8P.?20GbB#dZV
O63dJG>QQGH8;XR<9V/0J(L-S4UL^ae@\d/3C[-USGBg5.M15L>,C2;ABU9U)7A5
+E4^_>]@OUbY(0^Wg;]eMMR.QHH4e1\7KG\+-TC-NK0J4@U/<L&cNNd[,AFb;I00
1:NS=IS6B&=W4P9V^4:PKA6#;fP[XQ)5I5dG3P41eEPF6]-HVLF6ZD-X#O#UOL=D
B1OR=H3?^.4C/T;)5Q[Y8YF-<47#/b+6@]KK]N5C-ZQ2,Jc?[Ig5Y(bO2J#>J^=Z
>-^1\0A2K=P^1CR?VAY9I(/RJU61N;1&?g>Q8/5O67fA\RebS\[,F>QQfK=\6-]T
07-==40\\IRE2.\IYI9;ORALGcXJ=Wc=B4ETZcP:.cUdN4d<<TESKG2+]CZ[\Z?Y
Y6M=CRPFF)4W&<J6+<GGU1P:NRbB#K]RLRN8XSW/fQfOBWPKBU[C]7]IH_NKXLCQ
[,7/S:(?M>-gX.Fg[>O6WO?O+;8[Q#L)TVPT7\6/@B6<=+_JOI4J=eCVdSVYR-M)
VDd)AN8A5)3+](SL1T>&b2c?HMQc(b--@bNYe&X84b2gYg=b34^T_2MTS5a4BF:F
f<PSE/_H)-_a@;ZI(DM9WHa&_[DSaC>6VfUP=/;U]E>?P5DX(9aZ6>QM=BUIR2(a
&g82&KZA6TgFH<cN\6aMLK9(IHD87f[gMHT7PPJ_8.9X-WRDS)_C.]J#G^L91\)<
72Y:2N29AgRT0b7W4=K0UIDN:#[0SHZHO<S<fV<6OYFG_#MT#ZI#X([:dHI36NOQ
3(=a,aI,dd;g>HG#]7]56g8f^;\FfeAI3Y;9TPe#<dS\bY2X@#E(g((6\#(]=.?D
&dGQGDdT?XPbXW52U64=:da;HZ-T86^<aJ&^Q-6T/5Z0FW6a&[L#2ZKWea>[N@fU
e58)4OT:;<BJ8OMU?MM/#;0g?\AAIb0[CAcDB_CV[-M&;<EUUVS)LC9SdFHe.SfJ
66Bb.U8,_8&O<CKO20JGHB@EHb8-U<7W9Y@L)c]L@F1TdGZUAO/A2c1aP=TKb/f2
NE5g2=g[A)IW3.cbC+,>.VLRIdgR>X,_bXgB8DIFN?@X84C_:1VY38.W;;eA-^-B
2)YTLS,D\4Q3W27Ob2>.V;fT;LM7;KAVMZZg)aOgNE4UX5A2(:QG88#b=cXg@A.(
O@(U^=.B?\Y//GHA2>Q5DH[0R8H4=EJQ]RNB30(FQAR(NVBIa?W:LQ1Ee(7V]d3F
W<2bOFdU<HF8K.)J5af6;KS>X=^U#.H[g2;U;K0CJ:@@Cc;1_,C9]CAHH^+3GV9H
9WN2A#aP<Bd#^O8L7ESKW)(W[@(&bO8](#U[?aQ2aM\f[B\W>6:NX<7FfOTMG(_U
@e.V51HU@WIBR?\5,OV&F@?P-B3OM2QE6c@0;\3MQW1A&a&7cdPB4KYW7F^3[0(.
13PZ5EB&TP;D4>+:P@4698_;WQ8VE]EM]Vf#9RIXS>[]?I)3:Q)><VP15Vb5[G8S
2+123DV2ec]6\IIg91\DM;df5J#LRIE+9(7@18bS4e9/(A8^(>MPWeg2Y+5^&-/,
-1dQF,+\7\e:5FOV,Jf2PD=PC>A(@-#RVge,>^b]E<\N;7,7\&]-Y&DXNa6;F>I9
<)U<ZE9]:@FY#_(:5L@K9YS.-&DO-7]/HZ9U_-.)H^=N8[)=cQYP2F^=:Y>.1P&E
;XJ/U5@WaLRL-8UAD9;G@[d2(C0fG55.6A9E1V])R7e(11.]92;WRB;)FOHg1@TJ
0GK0\g=R)W(d<FC@/(5W6]#b?9B[T]1KL:V7^:\XcJ>(F&a_+(+/7g^:f+80W8V4
7VHb1O?]34,[0<L[[2?2;D_7Y&JZ8VI9bc_>F)UTG#Y.IW/:NEZ^@/DNQ/9\JK^[
J4,NGfa)3a@&F84/\,2?\5NTQfEC9?UbWMW;R?Vd/O&HO5G<@P.#/NK&#&DPOB^]
Q_(7+<?e=V-)&Y.(A3X9,/f,:,TZ+gX#&eYV<7bU5^-AK-PZD)FaP5gcZ?A4./[Z
-HVJDU75ff=]dPU@8,5I,@SQ5U01K?aJ?^7<KcN(\-KfeLb/;0BR7KQ9C>I7Z0Q.
M:;R<bLZdQcWYL351+IG1LF;f4,YID8^FHEa1C1gFA&baJ?0<-+,&6SX>_,cY63.
>-Ee:f,L05F_,_XGOgQbDV6Jg(/8:dE(5.;Ag-N)f)49;/Q2Hc\-(OYH/7(=@X=\
f5OB@LIV#8WF(^cXO0V,>6fA=^WSSTbOE#,S.13:c<d=5K[;4@/QfXO7=ad_YY,8
T(;_)(1\[^.2Q=d33M]?#LP.&=S,YJbR412SUI;=H3M].B\.[B0)V[_L]+[OH+Z+
X[///Z7cY]6+./HAdTHKaQX_<SJS4_ee&&<QL+bgNC=eW06>bVeEDXaYL&,Mb0E+
Q_adL/EY0E429\?N]\^aVN[84:9>=6-N=2V76K>\O@Sb>0U.Y;D-^93acX7]3I16
e:O0A+^.Eb,?)G\O_Zg2_#3^fUGI(0^]7U[O:L(f(DI-3ZQTQ?=e&QT2SMQMbRGd
A^Y\N=T?2LTdP_]A0D[.+Xb&)HSVGdQ\>FW/bQePVbC5Wc0(=H]3U?e.>^20d<4,
L#ZV9(0dE]cU<M/_2PEJ(B5&D01V+]C8.(H3LU2PX&9[=TR)OO[[,>(HUVQ-@WQX
A/>g3I0]e,T)@6R@A]LeE#Gg?U9M8<1;E[S(_L3c6,MKCbZ_5KZR>^8@d=FL@IQ;
_<-b+Jbf<Ya7U9gU?bbS7+b:c1+_GQ>;&U>63_V(Q>CAQ9;@f3DLZ_3<Ob8eBGRd
2F3g9FS\80,OLL3R>B8-KCJ\L-F;-IL<M;Q:?S=b]SQ6>O;@<ELX/_TI5Fc.VHLf
X9Z.V]_S:2QDN24DK8#-/9\1NbMC,F5M]30O>=[be[F?a[26CQ\^5;:DcR^5Xa\@
[8Ee=2W^dP:g]K\9L):2e--=TEf,LbRcG1\6^F0?@7X99M:HJSNANJ):fMRH)dD7
\#KBg1-8g9?VQN#MYg?Mb92EA2]]55dO&fbW_?3-M_3;W)B[5PGG;,gcVLE=fZ\O
K4Tgb=ZaTS-G#RE>^CY..OB(GVL<cbK=&G,Jf=5J;X/ZJBTUIc?Y0c+JIH&0_aE<
:AKE23=0@U2?HAO&EdI>D2S4X@b0VUDCOL_KbMM_dLJ14Q5:.OCW9]<CGV.[d[2H
;L?+4;59=P#Qc.TP-Tb2P1SB+/@7GESfbK^\cB]([+M>@@BMW+b+(F5WV[]R6LMK
WB?AACLQ2NgG10-EOI?N+baE^b8)5=1dU2M42N?2XM(5OaEe_I7\Y,1,Ed<RH:SI
L1_>]6:\gd&\X@,^>41J,N+_JL.1]B\TIDYQcZXE&>?:#5&[KP1<M^NK<X17JV+\
]/gYR9_C_3&EgJf)]<SGe;UVI;A0-O].I>_ZW))GWM<NRN,6YT4;X42?&dA:3R;1
Ja.^1#L1FLP7K/LW5Ze/R3c>H(TP^T6&DLg&2T@5(2=[7^9<>7+fNb#^>G)C/G8L
[@0:=6.&QUT<g\M/7_WbS<AZ2Q:#f51;)I+:J&c>L+>4=1KSc#[Rfg7&WKNX_gS_
bG.\aM?XRA:IEY>HeB3GH;eH?d6)gF#9YLC5BVI5PW>26BL#6]5\YGAY3FOf\V:^
g.<WP_1]eR>c_,:Xc:0O4ESZXL=4>&L9=fKS;#]Z/aGZ67GR^.Ygd5:g_B:TgfBN
>&8)J4;5f2A#>:I2/^CFdP6+F>G=SAAN#J<dI\b,2U=W75JP)NZ&J>\;<7KaacN=
T&FYHLN1O9=<WNJ6X)]=8;:GS34Y@@,/&I7N.KYNf^]2c0=Q#V;Z[fKbYHUZ@L<E
7<M;QcDd=(FTL?Cf-0d3bS4TV-L#BSP_-QV8X-Z(Y6AUXeJCU8]f0SL2K4PG6U-U
-5E0_4:?3gKU_3GQE;JKH@>)H&FTe4KaA[XYcaG)UJb,Y_H8-5G8OV5cTF_36eHU
T_JPXZ,&6VPeH6fY4#>QX_I++D-HK#a^B2^H_Ta4O&B;@\e(-NfM#CA_D/=)dARB
M=IMQ__7D1g<EC?/->c5F(&@?g2-]7<,LWI6L?Sd62eM(IET]gdF3^L+L&WWSMFS
MI^3378K>BKc:#)I5Gfc=OUQPY,cK04R[1WJFPa-7/bI)^2U>[E/_[9+1+GJ7g;Y
&K(M@QMH[8M\9.d(VJ#gKfYf7#VfV=)-XQCT26@T1Df#9gFCPI0P_9I?:>+RJFW^
TEJe],MU2TYCPF@0YS-VQ.:[K6V<E<R;MgJW]8A;=[:deHQGaWQb3+4LOPJ])=BK
YO@a)WF2JRDJ^_O-2K<FBIP.6abaZMVNgZIcWT-[@8VVP0g5A5e<>,=Z)ZL3B393
OL;X0JI0B)+2&K-.#K[26BKg:37BB2PObf1M/EZ:UQTc(D4&gTa+Z6YY7Wd2RCO1
LAdgH.9RI?d)AKCY]gAg)gXL2SV2>BQfeKU?6.7KFQUP(FZTaH@f/4W);d([2AL/
GFaI[>?,X,7KgLJdD9RbdM@I,eUY\d+b(a/(/d2B0\cLP+@\g8<,=A:^E6.]]EZ)
TI+,B14AReR@?3Eb0/B^b\AcW[16&=^]K4OL)LK7Z?394Z4J0:Y,5/^O=]J4YNg5
+CS@dd[.6dc_K3-#,]C>,V0]/Yc2+T]A_@@WEYF0_/ZX9D5,P>4<IYeHGdLWgMS;
HT[ORIM?g-O6B+NJG7-,A>+=;HTg?S64[/M,:5;QF7Ugf/-/Za,e4SANFaD&DV@L
RY\.WLE+@6,8.P3P<b8DM\HX4)RGIb=E&+]<(05Zd[LGXegW-Eg9WHa],>1R1O53
KM[\eR@RNQW>7W9\&XY9N5Z3=dERX+#(#+FIYY-Z1>G:U8DNEOPSCO)+<c#fdT4P
VG-b-P;#_&,_]B&gEIRDH3F/dOE3gcTYcde1.6P=/@Hf?OKZ?6S3UPT<#M9V703:
]=,-=-(3V]#?.BH3PE6JN8PI,S+I=G@eE=K7[W(SSK\5.Y;EEe0]63X_DLf-SQZC
MTT,(QXMU,GE@RFABdc7Z-7ca0HH+aRP@@=90E6SE9-DG_24N:>U[6d>eA9U]&FD
aK+F6Bc7A<0D;P1@\6=B2IC1DKV5H.e,P(3.4bEDE?dVFfZa5XUeLVE&]/888P_V
,4a[V<0X^Lg8@-_23U+c9YfaAg(PSX)3-1bCVV,U]@M0g70]2?Kf5)96?B>6e5Y,
RDFaEJWJ5DB244;^-+O1S2H]8EOQD<,-Z+Dc0O\RRRDURTWNDYb&#^+>Cdd43c,>
#<65B=)S[3)bUNP2\IRKX]8dX4]G=&R&Egb)8\fQgJS8U)d+IF=SEK=YK0)F>&X5
>4-7T0W>SY):;NE4S&&_.>0[[\;b],MM.VOH@ID,/8_SZ=KA4b9P1eb_]6RaN<PP
_4:<EGI<^7Wc/+M@KX(R-c;H\EQ=98P)YfW0>:3cB#eT=FUbNGOZ@V30SVGFBe=K
Fc5<Ia[WdLD8MVS)&2MBV6c^fV^MD,D[Q4:C=e1O-+H<2E,,gM\BJIC#B>G842G)
.9SEF=Xg<AgN;<I?&P<U+AfXd7SFg4@80MCLc,6c5QIQb0O-\\S<1#7H:ZO5SAKO
f3=MF<3fDb8MGG6P-;b2EP2_aX#,._9/7@bG=gQ#.cJZ93#CAA#@I]DCT?B#ZRc/
1EZ6g-ab8eC7RXgLVS/))#3(9D^d9BC=6D>#6\f8JgLP==O840=9:8Q&OA,IKEQ?
#Q)CMeYMZ+Aa;S\=9Uc-M[TP2<]7QB6]K@VgJ(,&HB1C6\9<\DJ]JWT?JVG2RB7c
4c1I9=HBdNOAVVE8Q4EXD-8[?/bKAWYLgg+L19f&Q/M</\fQ#C\L5Xc]&dURSNA[
&IUF(I[^c4^U11)HYT:V?SCT4#/IMPLMWe(MPUf/_Q9QRG]PQ6:FD>\0^CFRQHYZ
-]V7=dTWYNB__Q+8T<9dcaHQQP4g#7AgDXg_9@RKC]JB+_Zg+L\5T[LBREHfI[]+
<-(MVNGVM)4f=?+@3E0G+<D8=(=N:3N=bb5[@d?M+)L10b,dXSEX8G?H3.GE\5XR
]K;@2H66EDQ(,d<BU_RF><3>#e\IDXW/#^,H&/]N0/LE>01.Be,AVO]W1X>Rb7,^
\#a.MERaI2X2=_;4bOd.NT6E;9@GKLNE^G/=b9f7.KEd5G2O9bf^E.8+MA4\FdSe
/R10GH<LBUOcTQ(N?MX1M17#<HGXa8BOgJ75fJb&25K?_XcVcB6#EOWC5^#+MXM@
g12#AB4eHc(^gH/[2/90D&<E2DcfLH-?0#f_.A8A6,OW@<U4TQR__+)A#b-S(;:b
8QX/J+8JLD6>3<+[O61KXAB@TR99bg7^#1a:,7:Dg+E=]J[/d1JW<FE\\Tb7\]9I
Rb]2Kf9R=G._#\HMVUW/egZ-cE7b6V(cUO\0?dI@,I,.2<V^PIfa&-fB-AXR-7<S
AY3]XH-^1UJ[33cRYX]]8KY;NZV13a?\50Q;]S@,YLMQYf5:g>-9HKG/5Fe;^)N@
^Td]0aBZHV3BKXH,KRKKc7]PfTX_C&LP,ZZH5bg-6cUE(\1Td;PQ)]]:PbXf=(,_
-5TWXJZ4?;Y8Z(-4LO4HAIY(IbJU?^4eST8I._=#a/=b7M+>,)-P87H-H<BE=Z^M
;e&9>CHDQ.XIL/DXe3K\O6cBPU#f=,Y+-]ZAV.6Z]Nc@-d+L)e5J;,),@15gW#>>
87g0c;3aMI8.fQR=f0X4W5#eQU7VS6V4UF9<8/Y0_UFJXgZL]gdWW<>0O_/BA>^\
+Vd[3W81HDU_31/#&E;D92I92/(a]Q3<#?.OSA?db)-++T3^cdcL.XJ;P8885P5\
7<Lg02+;&F3^=IgOd^H/9M+g;&\F55Y7/bUd(I,^DDMM.c_U/0UJ^:0Q5JG5_V^U
&#LJT?U@.S5D;A)D^AcP1Y2/a9&6/Id&[\A?D><g-OECX_5/TR@-g&OGX_O9dXIa
:1LF:DZ?ce1T?DO:(QT5_-bH3cW,2;&Y?#bG,bGY.3KD#K^<eLef?+X#94Y@2aBc
(AK77cRdQEG,F9Y28H7Aa/XVOP?@9ZEcf?0,5P@2E;J\P9RNE.&I7)ae7.fd3K)c
B<GbJ=EHS)2:BbOX6<+L6<\Q>8]:EL,[;@.H;PXgB;A7B@+3?AIU(V\8V2X[_G=U
QU-gVD<U>7a]IB\YAF;UVd[)RA6?cQ(HVQU,G/0,0MJOO[D,+=/&V]9T#YfUHOJ<
\c2<_gg22A3F5P:QT:JR\YTF<1^7dHWY^4LV/KEZLX<MfLRXFN[Q/HPfZ>-g10:[
bC)7Z[4\5U3_/;I3@eJ9JMaQOPA-c]JZbg@c-RM,SD>7bZ(F;cc(g&,@d88HbIF^
C)WO^Wa^Xc+3D+;:V29=ee<eZ>cU2]>cBM78-d=?K;]1Z,H1Q9<8b^]O53Nc,D8C
dDe+SP_cd,/eD?\DKKMZT3NGD7b)TY[TdOI1YRb<b7Ia<<=gG+5JY;6e0N_M,Abd
]NBL^/D4D9<2e03VO3CSM4N4O8N&J;_b+^JC,/V4NFV2MSd.gW;T/J1cMB+dSCVQ
N3[EQ[#R=PfT_K^JL34<)b(2UBb^HRV1=YeeQe4YU+X/@Q0.FbgSW#C_a5?)aHL>
Qf(+11/4\.:fLbaJXX<GL@+I00A,KD@aHM;HX>;>ZX>XP?5Wec18.]\LK[Nac)49
3Y55IVD8/JSPA(B=<ZC#U0H^6VdZd1ge29\19#Zd:@6,^\MaA)4T3fK6SbSV2DWA
/EHYKO<#2<(.M8^?A/e&7V_Jgd;6gb)RTaN0AWFN1S>df>:cVMN-\-a+L\QT/R[b
D?=M(.9/25P.eJFg],(ML,c14aF8XP4VgY5;Q#GK[AE=@V/,UXGGVb-N,F8SR\\;
1gE?gAUHR6M##C?GTbT_]E&ZO>40H4AT4-@930&9(H/BXG@I_RU+4HAe5GF2g[/:
Y;?a)1EL-J9ZWd?M>&0]LKX>&cBC4]^WX\5Xc)43]8,BbF]@_)-gQ./J3^CUa5D;
e7FWJ:PX8?R]H-H?Ia4DI=g1f&7_YBW3S8)R.Z?)@acP0^Ba530A8Z77PYDRG61N
?UFU;F.649Se<UfGZNaQ9aJ&#+Y]DT[1@0a9P)8[UWL7^R:LR=.B^=g/Xb.Te/d^
&,4Q)<<OZMYN#^=5U.A=TPf?CgW0[_?2.SZ&^<O/R1?&V[9C?>(HHg,+6Mgg@8bH
L1.)CA2:>LT,2>:a8=T3g?2f_D-<gfX_K-,)F5@2L08&U(-X:Y?\4#+c5.e-5CS;
-Y:8M)@2C]S;&@8I5^,cX=Hg,X)[1:T06\0a6YDb-(O^>bIBUBa^VNWGATYUJRUF
bdNKQP1LW?(X:3U14+><GQI?(P^NM.f=V092:2L#T7OZD:eaC@2B:S49\eKTEf3d
^CcB<XWTX8L@F1c,1OT#I:b9S5&C1Oe&eN-7]B;#)NOD+GA_3dVO9JN,Gg]\IgR#
IcE^M:-,C])44)EA8:<-5FTV_]g\d@c245_eU@:d44K<gPgaEb/3NS4IBeKZ?U)=
INJDbCVLSU)XA-W@?f.ZS.1<>6,_5-T>b_:/cb-b2K9SSD]8b?@ORJ=LK0:K1Z5J
d\T1g(dbC=RLPa-NfJPY#T+KQXCXNTMR7,P]_VEf(&@4?U=UOg/L(Z6aT.AR/dII
5/#Vfc9A_UZ8E(OP><9_N1>TW;JdIF9:9&8<9Q5_3J1H+3K2_?:&S[?^58<;9TFU
YLN(D_D_fU>,f^9E=RF>0-U3?/6IF,e2_U2;9<^QP/VTC[fSYGI.HD_)^;MI65[R
.C>4c91da6@=6Seg+6<,,^a>A:&c+?WDX1#I_dDZ/:#9/@.(?8fNK3^BdTTHC:8J
408A,\5eRg0f1Q3,5:1VP=]MaVT)dS_PN^STYF&cGfAXP>?1(f+Q,CWaHBUMN]/B
R[@_;d1Vb[NGg39J#W9aK-23Pf]#dPP@38eXAUFD]XWG^B7_IIMI<.Q]-[^EId(f
01OXH.I2\1>Hge=b+>97LK2.C:GEDX/5TbF6/G:S:]aK\e\U&[\:b231HX<_6PT&
IG=LI^E/Y98PL1;X?_]FQ(1S#^0:HG5cc/._)b,K\9]1Z7X+[Z=ZbN).5f;#Nd#6
DS#U;+C2Y(:L902c0?NY6We0ZC]R,E&3FY2#]I1RddM_8AA(F8Gff--#VI>aeA]S
Z#8TAE:b[/Mc7+<OL14[^I#X3>GNc?]BE2MG=Y[OJLWCB1E;+4f@E>?<AH;+=;9;
J2S><0)XBM<g[CO^2/62)\eDQ=N#MMF9@WGEZ<V7.<^OY+Je>52<Q)FF=9dOfg(F
]&f1e:QVYJN<0WY^O9&<2fHJgb3[0LU=:G1P,e[<PT].RWNNVNdF#-N_ORIC&S;#
,1X<DO^/\)4??L;FYVBP@W:F4;0SdQIAbGBXa&?JFKWT.?^P7b+.K=>MHU6aFIG]
:+G4JBQ5]5ITW7Re8;\c6H,AWSYD<6T]@>YCI?-9ZP&_=UBc>LZd]FePJ)Dd=gYN
R.Oc^_OFTGR7Z[@/G[gaT,UI5cZaNc]XZbJR_PeP/.\NC=U(/(bMQW^BQE&C_L7(
2Af^BG7U@OXZ>+E)6J8HB5_^J=-QBJW5bA&1IE&dBW8(>.FF2C,.33_K2_I8D/UU
XSQ&EaTY5\,ZG3>e((4GD:T;M7)gTeF1VbU5F&R,Tc-IbXTA,;c<[2MN[3@K)=IT
Q^2PWL+OU>6QVa_&<Kg.U=S.(WGFP(H)4:V[^bcaJ53Y<A()>\VR.VV/=SPLBNY&
@VXNRH4R0>SKdW3&@.]4N/DAC4&DG]D>P#.O5Cb>Jce:#H08BM+FC81FeBLB3M@:
c9F80Z,+O,3/_@W^78Rb>IWAd)YFTfB#9Vf@STLH7+[?f8;VccUW1VKJ^DP<c(F6
@C&(V9P&FdDW?[dY2]B\8(9@26@=;GP4+P0b@-QY_7dgc59EGTHA3WXHULPKK\-O
Eg>^eK>:_A-HM]?8\DGW,FV;@c+_/5S_5/OIeDQW[gKHe>RW1Q(4M#71I?#/5EJO
0g6&O?ecSFN;?N7H^39:)Cdg262U0RYgRVH?82REH+935^-Lf]F-6Y,)E#VM#V+?
2aLFa6YY;JS=P.eQ47)Z@[g,BCHQMNJ:C[fGZ6&J:N<)R)A&?U#g2F8FFIGU>J/]
)eQBQYQW&JXR1N-1.P?,M=TWLXS=4085A0U:e.H/aVE@&bTSE>L]e8JNNE46E>UC
M-g,FL1X9Vg;RU)E/1M3.(TD_V_-RP<6-CDM>BFd[YS]Wg)G\PP1D;[VF6#W>eC2
@AJ0CHJe+6AD.SOT4(J<G&Pg]-46O+fC9L?OXE#=RbT[2g+Ac(A<d<L5Z[O#(3>#
?WT(H0)R-^VVc,]:@L-BRQ?@f1e54OWBa;F4<W/I24H@P:1B2]?SMYF0\1WW:acX
?6=:2MIT=WZ\OY,&)IA])9P=+AWKIOI7R;M.8\)1^?#bEE<FJTUUJ&SaL\da&g.A
_[63N=HS?M/6adZ-5)+XI0+_JMS\8P9Q.?-58M9X#/S56K]#?9&(P&X>A4M<.#Ze
9Oe8-2>A[:+AT@A^CWU6?5K/3K9>H:dgfT1?6f8NTX<O8:]/fca0XX327O#^5V,F
Lc=73[SHA2T^BgDd)ICVE@gPK]9aNH1&P7R6#R\=@_NTHQF<=3H6?IYPcAMQa<41
6-;1OV.@K469aC?:AH;1;W[E152Kg(:W8E_T7e\?I,7+e+<^aKT90QF-<g\H;PGa
4\DI+XYBV/O9Lb2A\+;0UF,)NAK-96826A21QX_f]cECM:85]6Y,d_>V)_O,GH_Z
LU6_XD+?KcLM_B7f-IJK_P)\;278V0&c;:)DTD@A#-dP&gX\ISO\L\DFe6GIALK?
cH1BW66OL4@CKAUa-g[aB0-;<_PeW_]U82RK]#YdYTcBH-^0E0-)dF,FSUZ6.QNW
_,WN@W^E0Yd7+fD;AL1><\OW7dE7)EEb&2Fa9eA;<W/KCTe-L_)9K,VRc(DJ.C(Y
8<\^ZPc.9T93&D(E8QF.G.^Y;\dO):JO32e[H(T6bGdAJ[9/f+3T+^ZUa>FV;)=I
NO@3[@TXY[FAM^8_YdSTd2.H+XcU715.INA?8\41gW1Pa_6Af3+SZX=@#C(KB9?g
5#0JB3\6M[f+ZaTPOTEWDLGI^4WE0-FS7YG]&-;0a3Hc7HZ:X6CB\..f^=LedE+G
ZZaJDO6_U2T&2+GJ4VXeI5S@4)6(C)1R.2HYJ#5fZ&Ee0Jf=Sd[e7McR3d55aaZO
/CD/1T^LTef7H]Q=.ZaB5;2M3<]VVY?[(f1)NbPCbLYFK<>GfSY.Y3TH=T1NBbC]
UCMOA>NZ)3>&LJd\02<(e@14=.-?_1C,#fO[Q,e0]JP_Af5T&XN1##.(6M+0;M.<
T?gF_CZ+;.632T/@-Y6AI^c2/HN)F7)V5YF;b]IE;aUeM>-fU/S.f0/1QccRE&cG
#0#H,_?;S_595TD1;W@FHJPEVF5;/gL-^^JH#&d9CefL#aE0&>JNT[Y.D-dK[U4(
(9EP-3g>Z)BUYZd0IY(V1I\MP#-],4DLQ#<_-]RC]bQ-E?=7EUAK0M87CX0b@PYG
D;5UC3/fbH7:3@4/6GL2f9L@^S^?]Add]TS4HVNVL?>XD]8V))f9&V;d\b8?0[RG
A(T\]QQbd&#A94aT;0?QA20-0==#ON-.>O;76T;NOdHM]1a?P#..B)>+L7Y421>8
#4NL1=&5GH/Q(IdT9SV,U<J(J^>E/C&eaaMegQKRQ)RNGRI0N[(-P0#:Y^JfKKC:
d206I-3d\dKMBWEVFD66#e^8=6\?89CM\\U:Q7-b[3C58g_+S=6U(JV_1LP2a5GK
?,?CZ48&\YL&+N8&)75_]gOGbaA+(4gKcb0Z=2QN0504(C4AF\J[K3J]L2X?&)P<
OH(]A.(_00;X)Q(Q?J)1PP.O_Pfe[Ib&>-b^F8cXYIKQZcfV4cP8A6V[PXQR>2PC
6D\?5N7SQ^]:I3EP<V->DJ60[TU;DK&UdD/3(5LbPN.[ZA]L4+9WCR0(_L>\(YKc
;S\0aHO/cWJ@++-c&\=PDHPWZeA5N[28(Xg-WAVgLR#5P8(S,7)[ZXBQ^Y+J.#_a
Gb?J&If,H<81Y2^P[BSC,:GaG]2JIeXdg03:Q1EaP\LA8Yf^AD[aX;O?9Vf0E;1E
]3,<E^4)6-WJNQ^d7-U+[_IM1@M4;&4?cW=D_;F(Q)f2&(/W]_>b:18OMJ<LVEUR
_eP<A7Z>)L_[cgbCd03<)/112aNI>WD;T]@:Z\[S[?9AP:d62@0LN45]C^(BHJ(K
fW=CC,)_?#Kd<FPG#f7PX2^]G27B#8_ZMMGVU<=5;HBA59\E4^ae3ZDTS(@[L5X]
,Z@Wa;@WbI6de<I&#9AJ#J;X;4_L^8ISTW_edf21>.@@F-HbdeS9Z8Y_A1BcX5g?
TUMReWQCZ:T(Of[#L\?eHQ:GF;8?IE[AW7X59RITgU-;/6GNf:8NP?RR^GC9_E#1
.1GB^IP8W+#(SZHHOd_LT2eU3g_XW-c^P:]U27(05-LTZ_0]/5Eg\0R_]D<P+\HZ
eDc#4?\C,WgLa;4U[gP-Q(1VBGCG,[_#LLX\K&G/I^-;Pd&>Bb7/KQ^+g3X#P-K]
QA)+A5>A;EIJDG2;ZgV<0W&96Z#D4NV(K\;,3RDFEO14ZC(\K^EG^aZ\XE31J-E\
]=@bESbWdI/d>I/.>></04\3Q7=-D)U#ac#&>-c\U1)FA,;P=/b_5<RJ3:^N56+6
d?,D>@MPaC;cfB1c?@04LX87FfI_CP_3<a_E<=[(F.NgK(CH3N<aZ35^E=W(BL>c
0OXb_:ZJNANY<^?GR\+4aD8((D_F@gR?\D(^:F6]aMcZa@PU5Fgd5eL0H66N8XR3
BU3P<>e9_2c-_\c+M9B=5aTO/:HbAM5D50UZ;S+W;EJ#fa,QfO_L(1DceT]A_NI(
(G0=;YA#R(aL#e;+aV@F<5V,UCJV=?YP2JIgCZ/V4Zd&_(bK;]F(M6+1<A+9-B)(
+.MKG&6L)(7C@fe4Le<cV_YeX83Dg5=VN_T6EOa_ABE2JF_72;Y^7ZQ^93=(I6JI
#N[.O>C&Z4^&WCQcE5Y5/OH9Ga.FSFcXaYC&3\6Qf;K8c23)?+(/aaC#+[.;@JUT
CXO=]5SFOUJC\gS#W>R68Y#<#2Ua/S/(##)B>ZeLTXGaT_](]@5L)?=?)bf3]J;X
&M2SK+?OA?;-=bA.E6eJbeTQY;=>/#_4H4(TJ50S8O2G#19F,La+0,NS;=LgXV#G
]AH/H@TE_B2\cV.FC9SLTd&ZfU@VU2M,KJS7PIZT/NgfZ@dcc4JR<&\Z+^7R[:N2
ZOW/eKN2,KXU9aB_a#J+B,8,=gW92-6=IdccfbZHgVP-8@(K:F^M)?]Y:JQ4-CJ7
dRBY^\-LKFEJX&3?4BKI@T?C]FB<e;FgDLPD,bF;46&>d72/8C15@BH,Y_4SRXB0
KK\.MLTR2QSafG9CK,6>9=Vc4U+306CD.Z7Ga[RJ2YV:>4+:;)#:UG02c[?cHd7;
\1X.b9<V8(E9JAD;_,@a?fa&U?R?\a^eR-62&?_ZA1\-IH()I:DC[@+\JB6=\H.>
&,@0@)>Yb),X6[X[^3<&E;aH?TD]M&ES>]ODE3;XfX>T>IBQPI;7fbZbFO?bP&b,
ROb+0A2I,]7<OL7>UVI01N)QV)^N]]M9QRNH-NZP&><VTG[NLJ>\I2=(D[Ob)^6a
G?0X[@)29]?R&.34MQV+=AU&=.fA0[-3\gJ,(d\H>;EQ,]bA)B^AG1AXK<74)LR;
..,^aPWD=P3(;-([OYC9bT5_GdR0eY98UORCbQI#6B5IBU\76CLTQDU0Tg;NO9_#
]FNI0=PX8J>SC/cNV11_I.+^;_2(5O^92c2A@e]>f>KNW;FcbR2@C^S^0O2N6T/:
98+YSJ1bEd-36L)N_ZAN:?K96B\>+3F5X6c=/KTAKG5eRDJX4c2<&C]RD)X2J&,+
_O;U<d9O;88e5G))b&Y3d39K-F]NgA:.BD/3OL)@W/.;a@.@EOJ31Q_JX,G>P[a7
@aM-cXA=)CgU#I+RE6b+,TT[2P2aTFeZY+V9AV?7gV_X0D/fMC;61dM>)@YGN;a\
5Ed/+f],YQ),):KSS?EX3YZQCI1W[;J,Ve7C5=::H#LgIJ6>Y>K<=;X[4e@Ke143
W0]]8MJ+1[J@BK31/((+BQQS>-=9._a4LB;SB)//<TBXDUWLHV6Y4;e?FS/6KR<@
F[b:[]@&7YC]MOPA83GK/8KU/:d#Ga)\(AI6_R;O[RPX7+Q[SEG@WQC9Hc+V]MVU
bYI>2QQKQU@N^#fG_R<M)g23RAHd),K^#Q1bOe[g0-WFa=gb;20_O<LQ/TO):eL\
g3Mc>B&0_^Z[9beZ/7<]\#f)13DL-,V]+O638M5EVcaa3H9>QI=E2?2<Nf=]&f&D
N/M6/OK-4CaD86gGg1_YbEWN92R/Y0;&C#PH<HA+@LV1X=WeB-N+R3<dgXaQ7HEF
HQ7:\]8:TJO3L(7_aC.3CRK#,-4\6+66DE7QcE_(31FWM79KWURagO@EW,[0]XX8
:-G<e6RENT/W-)>E^#J?2=T^?_?8<EX^TGb\0F[<RPZ[df0&;]Q_[XbSbQJV.X?3
7N9M(EETEIL([LO@L11\T#-H+>Q-.P8TA38;U_@CD>GS[ECVd<Q8NF8V=,b_c+_6
;DLW0SQO1#6>9\U/[OG_e(JLfX0-^I&S]-+N/MP6_UTfPb\6gC-6>2L0OGUX&VWd
3P>FV<-OG(K?C>[VUe6NIU4;ePXZ[A5^G5b]7DP+G8Y+YK(8ML\3)1KWWRR3H<eV
JTU\[7e[@PQVa97KGIA>.8IfJ.TN/I5?7]I1I.f)AFWN7^U(KV,31bZI93K?,9XA
P+Ka_)Ed=-L.PM0JX]K6gAHf@bX;e(BcMH:&@=]G=U9b5P_JbC:0M[.<:FDLb[(N
]32AOX)O6Y>f/ZXPbf>PIVX1fU,3BPJ+cXW89L9FeHU_g?+E/3N\X4WAFP=(-]?J
=KWC43g.cYTN_0f/]JfF1PGAc]NcC(:cT13_Z66L3Y3J5:c@X<TN[HO=0A-.><ga
1]fA8[._g&JB(W.#aSSgIN/ff\H3W3423QT))aB(SJ0M2XEKX:)QU)WbJa2S-.-=
WTA6C+C#/@#MJBGH1\>TOWJP[gWdC2AfCU27.@6T(+bZ\#VX3:]&PbgP373e=Q+(
,b4\C]b;#eGN>(5aRY=0_U4D8a.N/VK^g(S[cb7+<&^D;aJDR><J=W(7WG6^(7,:
5PA7HR\V4\466LN7>8ZK-(#,7?ddd0N&_eb.S_.]F[O)B;gBE:E+VYF#@bfe)Wd:
[6K,.SaR-XCIJLc3T26<VPdGcDZ=(G:O61GB5&\Yge&DRZaR(==[;6@9g/d[+[S@
=#If\b(K6YMUZWP1^([P+MFe;#KaT,2M1:#Z0XN,B,<^XBHIV+MfZ)TPQ>GEF623
;5R,e2?KdG6S9#I/><LN60#c.>;3[LI0T#Nfb-TM:O6_e3^]g;/DFR3b<>1T@SAR
4\1b+eSeUYaK[6QefaSLFR4]9YI-PG#7JC/>]_4+,2FY?=P>+>>WbIRJ7/1037eC
<VPR-+fAF7>:Q1edgX5f@O>FU>NTAD/T582#8)A+R&N<^^^c&JJdecUNfC?@\OAN
75SVAPgVW->cTAUAVZ;/9;W8V5TbXZYFOBT=Y70YB1G&F.OaFg7PZ@H8L]:Vc8-C
I4V&a^be<D/9bfSJT670gT1=baHBCA.A_Pg_=3f.fbf\9K8_)5[Mfd?SPa^B,;U;
.DCa63T6S3#g.]N8@2XBMG-ddAYY3A9OW>E>fE:LU;P^)VK;84MS@K31-O+;7_F4
1_N><,VeH@7LbYIBCFbG<^KR=/QL6Xg8D,CM6[a4GbSQ/M8cGD8I1M(be[6NS@A1
1[FM2MHcE+?[R.a)c5cRQ>.=ARO<bU[(X)CXK/ccc)LNQ\_&3.f[Y/;R+82fJ1@-
G2#bKBEH1NS:42IAGH.>dMOSceQ\Ye8d)YQJQ?U8_]YG3P#b#cKS6MBR1S;F@5aO
)B8?;:D^^5F+>g1bN4Ve?C=bMaMZUX3..^P?5/dPc\c^Q>H=X8?8KeK4>g]CHF_?
?<<X(b/Z.NNaNG@+4CHg:C;ET0:,9N,R6_aQR-,ZDc?&V=8(gAGd<5<^J3aSUYVd
V[#aAd_TWMI@L?HR)AScT,a#g9#^CYO=DX<-VI_@@7-OFIZLB]BMVF;G3+/53=P5
6YD2KOYVMTd?-#VFedU9VGAHR3YIb?72SKGC0A\T_eTHWE1R.T=ZEHd.<FSb\(>d
9H:eOY6Le.&C7MP1O#E^F)N0B1]]C#]D.8+H#P#gE(YZU62PdBQU&@Eb[dUB8/fT
=Ff+=242IWC+Z&TD3?c7QeHGf-C(D\Q/(0(dLWDcfcPbXZV:DI)99(G:dEB>eGM9
]FOCg-D2=3eD?P16O-F+ALR;_>IPO74S3>?U7A>_QPX7J\L1\>M@L(QERLbQP7O:
@d&,678#525HL?a-JPe,W3G:UH>+#g1UXZEc)X(^d-X&6_Y_c-BXUZ1f+QANLVUR
;/4VB[ZGF][R5/Z]G-a:=ZW<2^@.9<EM.Z,B@R#b/P>)7>e6G.1WQKM&DM.&f#:;
&,[aN3^fUJ.W^<#]DQeO>=06)HBf&^K#QU18)N/=<dg1bHO:ACU^fFR8=D8J_d[&
6.K0(^HCX9BMG7QFY(CI\;]ZBA0<NMYO+e-g7IV)Z(#]JR,=]C)PX\@/23N1b@;_
?A0?Re0Wb^GdFQG(9Q:+WT\\CB,:bU34YSg-#_&\>aIQaO#Vb\;_3;[+XH+c_Ld/
AGA&e49X7eaKNJ#X6.T:TeOX4b2#>/C(Y0W#0aQ-9,^5US(8Rc2cO]H55^QdB(=-
-B+gWIU#N.Kc=3L^(ZU-HSFU:MXHVg?UNOBbf,C#/Z?&Ke.NC7<L_JL9\<I&V;//
>gTR5S@YfQJ79;C_L,S&@0IJVC18&ILSZ7(=N^[]<bY#Vc3HT(BUgAAQKT#7.B:;
&64TT1J)@-fMYWD8G-g;PC2BQF\<4S(;D20OfX2#BQ.a@R<?.0#>(g@MJ55YT70W
V&FFZIG_017#T+ILacY+2K?]<Y1Xf1Qa2UK(H<\Q,aY_T7LJSNGKe0b\aGG/<K&I
XKE.1,F=dI,cJJ=VT5N;4=S[3CN&5X<<.OZ<58#RJE]eT^\Dd.)]6>M)CP53]<-E
G]EDb@gM)942U@RAbHM+GM\FE5B,Mb[RXf0U5Xe<3/,,C/_D<f\Y<fV-HF6gGKbJ
44-;9Y976<;:A/1;e7CU7SQRXWI)-B8YTD2[>RY)V02Q2VPW=WN[(+g3X&_69X&D
OJ;F-gL>8)ZBM<K7?\I9Rc@7Z008LgS_<#SgRJ:^9KN<U-CJ&I;?L6O8TOM)[U?^
@_b)_0[[a1?d]JEMW1G0@<ON+)-6KOAU?F3;4J^QP-7SC#gL)E,TLD_B/0&FSVWf
e)AE:,MNA(9LWbcWVe6B@>XYN;.U2>D?EQDHRN@#TED9X[g\ed-c;+]\LPPb21N;
]D;L6:]D+</?J8#.bN6\NNg)HL5^aI=L:#\UAC,/b-^(3.=G7Q\8?bF5dRRL24\6
I1Hg3c7ZM62).IMF^#2DPP:2?(^>OWY8FbY9XRg2C7>O?K;=7E8R=CO\]\CY>aa,
>(g-5CLe_&D;Z)/gBTJX;8IR^^Y3JWc6^D/9GHX??-43ZN,^1YZ9&:9gH<1.CJ2T
7_=>I1#E?C5>5>V2\[\FdL\AOAbY,]T@+bX,Wb@6_#KIZ6^\CG@UY>BT5O+?=5<A
cf?LGd8g/Bd:g-M2<g4_cMNT8(.+GNB?g4@2WL9&?YcM0H?&c_1c.Q(Y5T0P&?>#
HTVD@D5:5DGCRRJ#84K4W4JA3(9dd,d4[JNSf3g9gLAaZPU[E]+FLG>5?C)g?)>-
gGbU]>NZYMJG<1(;EGCa@--,-0/Yg-FPZ9J3\7A,UECJK_H[g)Cd4LIZ?7eLXAMA
WPLXAc<<-8AJfXUJQE30aI_R^EAaHcHZ[\VbSAKM+4g;^E]+=7T;SUIN\2U2b:78
eF]U#95GS7=<Md^C_&V1DC;N,&]>0@>7\c@,dM)[Ea.;0^1\Z3KB7C)bF[;:+)UV
V6-,,(C+DPP&F:SSE(_R^_S6F2I)=B\>RfIEgYCSW>fa)I)GXTbZQeBOPgM[gP:Z
KS#R49(Yg^2V<a,-DRNPb<DcS/9LVS^U@^Y\W@(C(_a;RWJ<&2&#^8KGYY4@E9R=
@DZU\1&Dc>-X5K(9\2<T/NaN^0UHYB]g/a6+JEa[<I,ELRSY:<GVNYeX]UB+.e8]
KL4_LMD@2ETIX?bN1:W?[H8a:@XC&2MK&_RfHF2L5)8NV;.7;A]JR[\Ee4,.D#LJ
N/<+DZc0Z5I8ZZ,S&?@-CR]0]96.<KU2VYUcN+U8+Y:BTJ@=B.,1_dcG.J1&>(2e
@^:=M9a+I4K0f<BAOX]1Q4RHM1dU7?T4RMGS9J46ZcG9b(Y>Cb2R)_;g@)UBC8BF
facF\19SL-(c-EP0F-TAU\VZ28dZL02G\=.2T@b45HB4f#A)H];5M&C#,b44a,BN
IR0E;gbMCKCU:\A^.D_<9CF7&#T)fWVZ/0H55EB\Jc/@0,bGZCZ\(=7P64U]e:e(
^\R[/P63&7D3dNAZ^,+AP=KM/d#;?K.[PEYfS7,CI1=N[e<74WL(K8@X/SH:ERKL
/30Xb(Ec<+P(bX1>:befMH.BNP;+6)_=>70WW@RDQVVJRYNF?;C]g6,]4dL2]][g
Q#g4LHGFSd6d35I/^a3/8J<PJ:0<>[\(<E\(c]</Z[-N-]QZ9D9fXH2^/85+EPHc
FTM<GXG/[A8#ZDU5E.8R7,O-/204Mf1b?-9f5N8(UXQAS;/2::Q[\427/CUXFD<?
&,764=+>?_G7UBM<IaA9LRVN0@\L?0Z4CU79U>MFL-UZZDe6R[G08;NFOg)HK5^g
WSb(WCd0D@0J)<98<CTD56[(CZg-M;/Z0/Ff^2-OA8V?eF/<DN)@_aBecX2dTg\c
YIc-&/gE4>45=cR?WLCEE_>\Q\HH=IKPGT&Qg>N<Q&H7RD59I+U1S#c39YRCJf5:
4012HMS/;f8SGfZ3BA4;VC,d>[SYbbB=V8&.\^EK]Ee7G$
`endprotected


`endif
