
`ifndef GUARD_SVT_AHB_SLAVE_MONITOR_CALLBACK_UVM_SV
`define GUARD_SVT_AHB_SLAVE_MONITOR_CALLBACK_UVM_SV

/**
 *  Slave monitor callback class contains the callback methods called by the
 *  slave monitor component.
 */
`ifdef SVT_VMM_TECHNOLOGY
class svt_ahb_slave_monitor_callback extends svt_xactor_callbacks;
`else
class svt_ahb_slave_monitor_callback extends svt_callback;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_ahb_slave_monitor_callback");
`endif

  //----------------------------------------------------------------------------
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+yv8qCWJP5yMR1qiQiVvYAP2fCK40qXzgKpui2Eqow7nAhPsFlxNSlrnRJvYoUV7
Cq7O/Vhb7/CelmlvwQ7l/ZUGXNgweGfn9PDyH6S2SbyZefJfxymiMYEsEhWMS9mt
Pj+Afup1taiBLFKZWB0l/S4HZKc4hZ/fzZNkSOjKmkDutNxKwclVRA==
//pragma protect end_key_block
//pragma protect digest_block
5iK9HjXtRZVlkK0wFQxVtfq+Wf8=
//pragma protect end_digest_block
//pragma protect data_block
S3Tav9kbApwADnxzNT6aOWu9b/+O8y7FN4N2fxXebm1NbWXKemNYXIz/8Omp2WTb
uJ/CKenddIgiUipcqeTUcsYL4BjqeaTmnfRUwAt/0I+J2OpOCoRTNUFqUDu4N1/z
9u138mlblX0rtpmXxog1+0Zk3FKkvEBpJ0ODqlaZI0ZOrKcst1cXxf1/fhoQIdBg
0PuAY2MkZ3RlFGMaFii4E/7SU/0fdYbVpXsFAkfXYUket5MaKoWqzxr40pTjEIhZ
4MkNH36mnLMuPZBNqFapvsRbePZO8BZUEyNIasqrrvotVCksqPG6PTXhw18qkrRM
A+178j2nW8pD0msmfawudTn1F36wA5jTF6C/yaPvJcF2zZSNogv97jSMWDTz8Iag
1GJdIms/HTIZkxHT0PZqYW49mklGc7ggK/ssECTfh5+EpJD3oPjvZZcFoqghsPFz
zO2iMqOuNPUQDZ7DJtbXHmLoWhfDuhp9SZIbHKtUHJaXNHm5j4/ERrjdNZckenOP
x91vJn2Kg41euUZeee86LCsvW7T9dDVl14jJmTHAB5jFNRVFkAV3mULxjIjpXowd
G2PwIn141BuuOUK0l887X8moZGK+jo1PjKiMu6bXw0nLvnlUavzFuVBNeqWSdxuV
lUE9xRt//polRUojY0vgeIY8bvfEQBp7sTnA4AN9UxRMEi30nBzKWkCHyKQYFDpo
MppauUkx80OBhCX3Fayd04IDfJI/6gcugZy+8f0kAj/HOYSX0sYG5kDxEwemDEan
der/s29SVUU8332KYVobk93fKB+pBg+TmoygQ9d7mAlLj3fufulRgOdTxesgjjWL
2ASZtzu+3gR/8eanzlszzN3cuihZZpoYnDTUpX4rIPPGYZSTcH5Fco5zBQJzgB0v
XMkw+rypp1ZGPjw9STzNHgIHd11xoZx/qeoUh0X6PBAggYGsQheB7zpGsjtXwM3+
PKXHBJP6WMoaPlMA7dBmKKEveQvtXtrzomyeUnO6CWEuBHR/FYeRry7Ouzos3Xrs
uQ84eTshP+87chOKnbAHq8DX5iBeYSON4y0nqUoO2Jc5+wblqKuPPS3jI+iKMKyz
7l+qhKEI1WDHvUMdGf3kp7HhDE+icrYgTCluf3t/pMqEGyfheTA3UMStludJ5XT1
5l7PCOxBga0bipDL0hZq7L/BXViWAG9K9W8ekm+OFeix987dVaZeCfPE+mdJ3cy+
CMEJdnYchJrCWStStutdC7NyXmMG4R1OQJJ4CXmqZBUK4dKGS0t12n1+tUk4ZF4w
AdlNtmHuLnQNw6wjFjqt60x+EXUObr7ra3M0baLdw3F9PlZXvVGnbGFnPDR6w/wD
SVBLwRlOPfbPPbqvoOv/fb7AxQmNJGg5ckB3nQ+7tpkykunOA+dbTIIVxKWPbrsB
gLeDTWBGJs6nXkplHZmgBbSIePMFRY9QJjO6ZzSqmZ/i9MzBm4pHUAE4AEsmkENI
xbWhD0jhCp9kmEOj2xsJkg0YcxZvTn0n/n6znyJqIut6c+6MTpeHheQV5a9PlXMd
gqhBYz0G9BfiUa4HFX/7DzcQ4xPNsxEBAnLHtTplZ257zw6qqCN8l2E+FFP2fzW6
u7VPX5fwPeoc6WtUedofiCD4+8N0jLYVsqcfITrhyL140EdQ/2gYFBbyCN01BXXX
y0aEOI7rNA0oWZEMvGPFjrujhNh9QAx1DRUBe46K1YWd77Hwf3kus6Q2iFyOdMmg
DfL8Vqt984InwIpDcLQINvH1VRYSYDedJXIpN5Fi9WCxilRiOdel2OKHFFnbNlob
PdlUL9MV+Eewxaa8o6kFq3SU9ATyl80RUv+wz/v49McZjo2NjSgQC58PF+49MVfD
p2YxtRwoBaM8LFGanO+jkgPio00ivAHLLmZgWWTrrFRMpO8rCwPLLkF2wilBfXWe
dh1yRq78VwOFJ2km6dDEjf0WcJ4Ai+vJlm6rmdQy8S7Sh7r1Ugz8/K5xC4/q6Auq
0LrKncmLmGuTA6Kl6cY1lf83Re18S9BTD8VsrzlINeJ1JFj7/q0qrGqG6p6G6meT
tWD9ijA7CLmaZQfPZy8zql09uRESx8Uw0YgKftCnMAJ0P0pcWRviSEFD9+BXXM9g
kiOM4y8nUw55WI8ACjJLJgt17Atrh1WXTN6aIfhzYB9KfaQYBSo45oPRlPUMsOqv
vYRDqW8Z8cLvKeEH4F+QVLs+iU27DRq+W1Anw2pXHjKet0tXyo0hcwdqMpD0Z5E5
ROaKc8XWUXudfuKN+R+yPjgsRGekTHJvpGHCCTVad1EgaPjMMKk+yldtHbrAQ0tu
iTQ9NpxTBz7P1+zvwaBQBBoVuKgWg2LtSmGI74TVNgT+xOozpDavArZisPJSNBV+
pG8gEgceQ+NsfsfPMjAGz0d4zTStK0CF60KmEiivxeN34LIe+jTTRGpwmS6fzzI1
NCwxzsWlJt0LD4IaAwYmpdSGoDrlHAnmgxd4F/8O2MNnK2su6r39ptS1ZtuPaI/w
eBJO49/AN/E7eLBq9Q8O+3Q/UmX7qtSIKBRzZQ/1usIo+gdS8XNm1qyv6Gi4oNx2
NdDQoeD3V7hQ9aI1A6Ou3Z2vlVoCTdLby2cNwOD8BH1EYTMiKG1KK3llDgBA8Yzs
8YBYkAnxdp/4w1HYEW27/Uct9X11yf1tfDE9vB7B5Oog5vSxh/bJJhC2ClDLTms5
y/lFCDJCshaaRcyURTycW9apxVaIFUHKgKLXfFRze71/6nJa6aBfmBLkbFdNaQBO
UKeGMmXXkC9KsGPDtqQSYB0Gltdvjm01BcI8BLBClRXAEAPHYD4/J0uri8g469zm
b2OCgINdYPuj/KqgPBgr0JqTXNhwJybXKNMTvhDYgwMN3+vnJP051jXLBJkX7RJm
HBWuv2foO8fSd5faEogAVqZOUALfPeBbkP/uKjLkuFm4KIM6EOmTN/vHGbPNVW9X
WZCX+abzsOPNSDQFDyLFKHJr+bEJk7YpbXorfWa7NDEg9n1UQ2bHJaqA+Df99d7i
xpqrCdyn5ldsSVvz3lIg6MeRXnU0fyq/7uvA11SngA9SYODFb0fXZrv1BL4FECFJ
z/xgyoRZKzGsoIOBHbdPu0htEJWY+lJXnlhFzSoDqU2rBdvxpttk9ZdZPtp7c9n2
aGvRO+eClQpYp8JbSkAAGAbFUt0S8fbCG9z5r7BpGQ4j7n8chkMc5ZGTZBQvO7dg
CmQRNCDVcZSlW9uNaTxL6zmbpbz/A3FxmP47XgToNYvUUoHjcVUZ85ueoHGSCgHl
dqNuWUTr+at+lzF9EWKMBjNtOEwWspa7UUy2QdJ2mbt8+bWvI+KEm5Y038fLHejU
B/5MAzZOUge5WowZCgYppZjpwk0WoJv8rFTqPU6N3p2mUj2aOuJ7uyMro54kQ37t
qwmPURMCWEpl9zRrDw83k1g1rkk8eE2eeVWwEa0+r8BDBpB4IyCdogby/4nTcK4a
ASMzYK6fFjVMRGXQ1zFkGMfJN3ok7IhAc5m/N1mT5jNPooL+VC1ngK7JB8y7Cwl8
ptofx80WD2fFFTnFGRe+ohBxiWGj4Rw/XMlsb+UabsFYQe8v7gBxOqarxBM/sVH7
NwG3rUhjOFmMyrC4cOffvee5PKOA3sgk7MTDtZ6ujJQgPgwiI/MkPm/K3HWrMtGH
A5dzzJZSDHy3rx1c4yYC3MDzmsSIXKfKi1f1PS3tpED/N5/vTCCR6AJEyDbPfHqj
s3TzvSQjdYjmU9VBKSjv5n7toAWfxxJnNIbTpv1Q+IRKgQ/P33GSmlIkl7cA8Wwm
L7hVxPpiIFtC7+iRwyGsO8udAqnm+4vEBACzNGJOTeSO1b0H2BPYmlI0nlQ9JVMK
762VsELDQMAKqZfHkgcqDMgtzHZBrmGhIgM1ic0LaucX2xympsiCYWwS+10NySOW
UPdPJ/VFxAJ1mUhL9rkKob94NlgstAJ111d7cgQySrJXbNAKecZRaA6Y3eQ5KFwY
ACG+qZtBCbl9dWj+R6mojfLj1kgGUeqUk6xkIVx0zBkYVF2dFGFc/OUyLUXdhwZr
dD6ZYY4QC2QvKT5TknZdQSYkspJSvxAXo2GCwM2o7eGyuVYV66AD3tvq1Vsrr1np
5hxSsBBbl3QmWE4Z78rHC1gQJ3Yi6/USBpVtHcCM0iP3NhFn3e6qg9dCIlKFnQ2j
HKbihaxN85inZ7JPsiv7rtyY2713Absxo02WJ6QtVopvtpYaRAYHAq46+Ol9L46p
09yUgMdA1s5BJbw6/NavZJBPr6KhE7fNZWNWFl3cb/frsBkjBWGorexQFmEny+7Z
jwWmiB/qSMX0OoYZT+19Uo8qIHZ+vuBRLeL+hYDDD+tAY/IMwT5nO+De6S4vimEK
UoMyhJYkfWMd0RobIkz2RZyFqC/Waj6ErjfDDqH+yOW72Mo7SMGOofjyDlu1ktlt
7mR/Hhcm1wO62K4EXKlT4HUGdeW+1lHk2iHPaM4wl4+XlxoT8Anxx5CKtmWRtU7g
/u1LA1463K26DlPW4r58JVpzB7WoH1uBvhPiK0Z0wlqZ5V8FF5oz/ndSgJx54e81
SzW4x9bZJYtDgSYuXJBjt1oEFXvatM1jDqByqPvX58AwcS/PNzGvtXWRr3SL0z1J
V4a1e+8MJS8LFCB0T3MHVUzGGMpZ1Ets4II8XQWyicIjxD4+Hdz8xbLjHG+KgZW4
ppfqOQxvS6szB+6sI9ZjMEnWqoG9CErm8VpKH4f7KB7B457NTjGMW7Hz2jYmrPFc
cWJRmh1FMPa5Tyh73qrezjSuADFKHUiEjCIF/6qjO9i9wl1sDENeSWEkfmwVh0yX
OJfc4mXM85tMdwTaIAJzI9fmaUk52JRsyiW9Mu0mAYHAnULd5zLBZZP/oYk9QxUt
jCyRtiJhj1ZYFLsbI3hE2MwYdVv4vqgrJwvC9sJz0RbZIAgPWMBa0mr6w1s0zXfb
J8E5EXIO9NkHiK0TQTPMx0wVs4NzRwXju0P4Grxv7I3WDCfPJQPd+cir4tvIg/6Y
p7PsZLzfCQatFak4a8xOs2EMNCk4XFVRoUJwLLSWSv/zpuQJktfy3E9xz2uPFGkK
hnGh+24tSE1mzb1gh4o8D7IF8r/lwvrUw7ck/XKTCXVjteQYHIZRT9aHh92CHI/3
TuJT3yGt6ANFTcZ08PL/qOjpmPWbvtHv9PDNxNkWy7+S8bqlzkIvKEksNs25fRH3
1VsLIrzihoc3qjjK7m/NPhMMzDdUVEpadtkNsGEcgDtTZOtkdGfVogmYuc3xXQTo
5X3ez+C3eK6Wwb7o/a519spFQlai13t8jBQoSgvkf5B0lxCMrePyVDGceKhcGT0E
Wtsf489k6bMiKZqfPdlDGdRRTvlO5v2JqalEwUByfYy9Xr6u+echbAsC3IAyeD5z
1eopTM0CbIjfhinHtI0Qf4eY1QPtfCSOwE2m8wT2Z890/jCRPoIz7yjFbgpOvSjM
pQS/jv1PYhDFOxfssvQ6mvushFqczYAmdiMHzKU6IQXoaXlhTXz33VP5z8fL0awg
xmAoRJ6TLnr9xFg5rXppa+xWLkWhoHCAZ8u9Am9yTuEXChA9I7f60oG0HwnLI5kX
T+DAN7j1EvzWt+8iQkDaLg/d4VjdieeS2cVcRYhA62CsPK1u+KZlFtCzg6HBKrSF
4k8089T9Va4DrpADNsLsqNtkGcZE/6pjLMLRF4U1hadRokhNuER2UI7LBBZKNDKQ
j0KpWKyAmRjPk/t1jbQ/sWRGilzrp4XcaRmsH6nDpwnUdng4CvCRnyA2r0wGyuGl
N8O6ueE5xf8CBSk/yk5HzUOwpFm2129qQkBsDp+xbsXL5reoVSX370RSRmfhwG8u
XOGNJby9zsgwrRRCqF9JojK2a1ND0igyjbxwt5WIYlolZOmyJitlgIHK57UonK+R
DsB0NWQOwkc/mksFdekJmEEOnG/M9xe5w+DOzVcsi0QkLPU23hVivRg2RTesgLdv
rugfrRtzeY8uGWs92mq+o6ONX+Kl/FYSyac1hqHEduFk8IosiNKc03nZS1fNfE7K
XYsmkbmfevI81ClSxfMkcrWT2hg3Mj/Qinz3+tX7Wq/L7D7Z1k0MfGc6X/Z9ITf8
6J0u+PgzzJEcAUCv2PndU7AjptYS4ZsdUUakHSsy5NNilkSpYjeBCtS9p7LhuV6X
fKRiYX/nbBTuwCrpCIRWtUxlnusQ8w0pfNYTH3qHkOJjVi3XiRtUok+2j3LHuVRf
oUtpuV/ju1i7tEgmgMYONrc0iVzjHZINkEnc9kxi5Dfww8OVcVf69foO4GmnylTu
w0F/NTjmI9I4FJ2s/Uj2oXVxTCRQTzZm9YeGTbOuOH1kJJAv6u8gE0snMSdjSV/H
1zFXvkn0jEHQ1HTZIoivkqclU5OCzzBkGFjR1K5gGxNRHIUdTWIiQAwM21lhX7+1
mOaWCD+Q/BZRJw43Gyot+IlWe072w1lU1wC5LCTkyQzofVckgAAkkGhlYcTiU0Ap
S2RzzhANHPSF9PryznGhzmbVPD9hKAQX/FtJW24aAe423p2wp6AnKuO/z5Y84WCm
HroqHDwo3/Uts2ioTVlmUlIl61iyW7KA288h2vXAwR7R9RZcaP3pVoeSRsGhFf5T
mW9cVxLpizri8N+8+g4KZeDmKxaAsj3mbWLywR5HtieH5+yPTxdb+hlFsMV9cqvP
VS5MH5oJIVxTY5VuFJr+b4V2H0ln5nbRCV2sRSK5kYYLbhVgC/1LidiiW/tV5sKI
dbCzIf++lSO0mEGBCI1MoeN3fzglSBWw/UHh4sORXSjIMveyN04SvH6a6GFi5lai
nhhFeT2D4WuNBpeDdk7M1l9bXDqolhMlzXykDp0gff9brs7p/r8SqvO0h57fQJeF
0+rS3vPWychQXr0a+N0Emw2GZ8rkLVOPUsGwHYdhsoU719gf/j+uQCulgRH102pF
5nKEo32cXRfFkeRyu6SSIf/1YnTVv4+Y0i/w9G+X4Afup/VUxUwBKK8CPzI54pRz
WK9JCF0oMO+Tyd6Tp3W0yNie8zY7H7V3D0mGS5hgrMjr7DaIOMkiF7MM+Z/tKvxi
NUJlGX0zkDDcvervur7HilCXCpQFqdu8ATR4AYpb3889jWLWDeaLrM4H5hJGqif/
vTntv8PlM6uWhdYr5g9pmp/aBn+UYyIR6rZSta7R4EVxmQgKDry/R807lYEXyTfz
OhEvGlx7k4BVYoviSyH4xk1SrgVrSqT6XcM+zJhrZIpYkk+RyL+i9hMd/CqISwxT
sxpXeQi/EMefkWgYW3J+G7CUdJIfmck0OP339y52mu1Y+2NKCKWg0npZpdJloLmk
OzIY1c1rXL7ekR+R1zrhn15QsCJTwwfEnV6Q7IQGEskY9n59abEBPrgNBtrUdHBs
g2Rpp9rzyCJgXIBG2r/+I+tWj75hBeKemvrQ3o3zJES3gObrzRvnSCA4mOOwYkIy
R/c9TdNqL0/VjQxu9FxFRB/1WDTg1bl7PF3y9hsODdb+J3/4IKYBuVLs5DZcWaGk
/5fJeHY/wbrFivwEjNl8OXz1pVmElUCpdZ13mebNADk3Og1kk0hwGW025kCQNd03
sfNTadbHgrL+5R6rI0QqQLaMmOiXS7F/M0vAS+Ku/ESDnIMn0oje1C/zMozIMiMY
eIADO6niYdx8pZYHaa1BVdVNXLOFGvB3ZecE2z8TbLrl0mRIqAG0J15em0ydqB/0
MX1UAi/jpp4SrzodHfhbK/5nZtyDA1XZIEQrjt0S4pYpH+I68uHTEhwLsO5MGjzx
5Z3ewtTHCJxGedd0OBhNVYq6vi6NR/83oEMGOkvHGmC4T/c0GsHvR+npaKGKqiVu
W7Cn6PySbQvMRcJZhtChJE5smXD2/uqH87b5MsloUnhn2n4VbPFDisGEscXNdhPD
Mmpat6GJwxtAwLX38y8L+PUsazgKp+Blwa/vvhWOlzaoiV3Y00BecmU697cAAioS
qJdwUVYtHyqE3qg+m/EgaKipI56IYgDUllT6YVFGqvOQhkhSfkH9qe5wnIpR9Cvq
PWy5wom3jux34/sXLKUabqht3mvPDg89Sz+SdsUIjEqbHfcJrH5JQSVaG2hWAgJI
kbtiG2ElBsq0ru6GYVLkjVB0uXeALSnXSJfMBBmobfrO/hcmY9/KaTl4rXE60iFC
abEeXUH84dTOwCKgaLetWVv0R4lQWZoHOLfGEv+E3nTT1BlL51j8rz5gzqREDRPg
LRx2Q8LwgNTFml0ixJ3LLy/ozgyNpEebhyGal5j1aohP+I6zEdkESuP5k6UlOvfb
6QvFxslmxmwOyuZn+QyNKAhAjUDbe2f6aW7y66TlrRT6GwTKpP22HZrrrvSpHUR7
1rnOjlCiSKmlACc1z5stED7kErnxJAjwM7jG3WkghATXOjEjfp7owOe/XM4OcGcE
XfOI0g205flk3Ok0CSqFydqQYCFsJ+zas1Uar71Lck+Q/AY+nVFGjIgPslZikTwG
QNgtAsYLsQQbFVqeI4pjItHf1pxe1cc4zZnbW90OJyUxty48gQ47qCIAn4enBOQI
sMv/Iz2GgSI+nfrzB4xmN361AVgtKX2S6D5fYH6Ip4zaD0VbDbLk9EkBgk/tfBmd
eLaKa650SInCFjqNI5Z7LAsG+GZGE2xgdwwadkzUUhAlz0IejALtcPidPUWMMmRd
Od+dmo2O5a+yKV4tlfbIh/A9GDkrniVK2OjdXM/cFe1rOYbu2N6sQ/9nLtzW3xqs
Gz9pwEli5fhA916J2wiY8PnAbJCaETgWBY484wCETrgG0PYlZ0ryhRu5/8LqoDJv
hy8Bd2b1xRwXS7Q1L1WTVJUN3IRq1vs4tVberIbOGUHkw0SohiFUOBkHx7TVaOrQ
4IDQG+HRNGrhm8W+hchueUEcQlkZO7z8BpmbP5hxhoB8prMTthBZjAI/MHZAWodj
y9nJYUtKXvRSU9mGL8scnSimsZD/BfJKg5FmkEb4pK+AMEDncJhK3NLAHkmP1paN
O+zOsNDxxnujXLE/egnccViiP/l+SmxJXpPDvIud2wZS2T/GSnnls1wuzkGZsGoS
AKQpXE5YZyjldHND8Xw9A2aNmEgopHqfDE0SF0XlEIYf9ztr0R7MWrotxomBmEGx
iGrd4f6/tPNWMXUPttpGu5VHSWx6q/2avUlv3m4bfev7Kus9SpsBUbpf0fH30eqf
NWv2t6X8igevZ/C96niGYX+yFekvzqUb3A0b0M3VoKnPdtwXOUUr4Xv3T23tG6+K
Snkg7HFm9UzCl3vQ5IYc77cXKnuwA26AJ9Yyp1kwxSre4cRzAi1YluklYkwyfQF7
j7lNjOUhXyWBoZOj54Qcn1U7si2q+g5yCDjgyFMSVS49zLCFAS3bT4/GXg2Vjn32
GgRIIUS6DcpIMXciasTTbj+r6UtRK4YnJJ9+lnYbhL0Nd0+I2FA6ZaCRRJhQgYem
vJFB4fuWulm8D/tJuIDRLwNKTRZJXoyYWHotQ/dVozHdwDVOnFtrQaO0DUk7oGVS
l9BOAQrnhS1777djB+nW2Kc9hVJDmVLO4sBsnoWt4jfS0P1FeUWrKOsvmlxmVhiH
Jn4S3tHututJnfp7PogWYgIoNOu6rGzjUW6bo1rmRDKIoL23d0cbEIaDLJo/o9ix
oaSi2Bq+m/EIAjYHCmwTu9AwtHyLZTNQ0xFRCR0W36wsUOrEI16aKXxZoEoKL50s
+5Gfj7XjtTqSTSTepQU7Ab1p2sUXN+Ko8kcDw8b8TbCDifXBPUNjUdBvo2Mx4QtL
ru8dVBHcafCBZ8LDy1XtPUGKuC3CI3ODJqcwLkruQS/33PzsLn+OHkQMdqorUWSu
VgUdxGzbgSOSUlqRvF9qeR9mclKtlCZHNjKuybBeyw4h5BIVn/jcB3W9MWwNaGOR
z9wtJl9EwEjLybLqp0IPcTKDQNHdgKvNPNbpWwaO9M5VFfGzY6/KPdlm1A/2FiYA
qSGdNlbFCas9sQ/7JyNv3zP7MQC8q7WwO4Vii+FUJAvgrX/yNLIax5aCHbGeZm98
TFJXGt9jIAlxT42cTkuOvXvAziadn0kK0YmiDWYxgo0LLTCbTBB+j0Mtz9SvBLHv
3Pk8NtKk3Zj1Xh/YQxhoXZf+1FlLBsTM/ajQANcuni5isgA3KQ886nrubGRgtbDp
f9PB4fVQSZSZLmOZqKTSX87W2DEd/Pw9iqDgQ3Exed/lqUSHhd1L2CdgZPMb3KkW
jVAuqLcDPLMfcStf9xNLusEAkKoCOcZKpvKxRXxkyBzLZ3jwB7NvoK9jOq2BTWoF
JzRGeddac0pdIR1qnpflqfw1eOMjOH2jCwG/X4sbsm52XAvGrIYX1REKjWQWlZTu
r3wjlqhQw3+9OInxGz/LjFHkAR45iA+Z+z9GbjKH2AN00iIjaO7QrkoOzZBpxhOX
7FttSq2aNKawiX5zjlZW+Vy9oyNhaKaS5Gs5QvGNpU8=
//pragma protect end_data_block
//pragma protect digest_block
tAxOrCC+ZrKzfKGO7dBecwMwxsY=
//pragma protect end_digest_block
//pragma protect end_protected
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
rdDXSKKRbiHgfTxRlWTqL2FuwHOd9P8EctubEuBoCmksfdGvJbCmwHCL9C7ZN/+h
KIruhBAOAOgH8ndbLYMmfU1QT8V+qttDZxqnX8bBKmK7pFy7fDtxcJvVaDQUPZXJ
tzVmAXVPVPyxmUrbyB9yKxp5KFIUSLshVFEHBCDUWwtVQ8gML03p0Q==
//pragma protect end_key_block
//pragma protect digest_block
THftKiKQUBIvtv434milqjFL4Fk=
//pragma protect end_digest_block
//pragma protect data_block
oWsAde8EFnwckN4qcjP0wEi3wtVG1vGCrZunenLPIDBlsgLr1qTb54aAAcUTSPn7
C6XzKIfzvJnZXNKMzy3pQDJzflY8v0PA0ROsZTHav2/GYDyZ4d68xhbLuldHflVc
h2H4S8MJkaYcboalrTwUMHW5nG+gpwcgXBuGjxyXcSzWsm9V7yf+mO9HZS5ssWFR
Y1vrZvq72ZQvfu+W56KB53h0E1qAftKDnO+u3DUOjuTU6c7seJqRih+qWJhDyvGu
4lyYw69/yOKV0W5VKCFc27u7ftiR5qk6eeMn+mLtD6S7ODydm/xiR4RN2psfUMrU
2fYQz0YO2AjsZB4FQYBX44Jy3sg3XBNluIUrV4xvo71LyFbvL2VvpSri11R4shn3
sa2UqMz+EbhXbFvUmypV+OuKPgZDPGjH6ak7vvG8TLCliZjD4DtXcjilS5Z1a9Jv
0rX/ngP5t2BxJMVEYYc+kyfHxdla5ZcZBHCDLamlTez15w6u2UJyg9/JDrI2Wrru
qOCddFpBw60skrtU/hC+QFprgWjSebZMUaS7aOseP+ewrkrAOSfDxqh3QUnCUzL2
Tb5ThdWYDbB1HtTgPv0AwmMUnhSo4FXuHc0JSndHJXlLeiE+OVWp2ergteT/yYeu
W1MGusXhthWtD9cA3BIcZi3WGbfGzRdyA8653LV6GWjrTl38u1wt+2c0fbxL5nw3
BjuuGWJYFvPRokiFWo3nT8ofUQW3Xj9XLCbHSqycXs1l59Jgmb+jtQc/5uEMVuxS

//pragma protect end_data_block
//pragma protect digest_block
h9eP5cXgDy5CGZtb0OUIt0FLRsE=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_SLAVE_MONITOR_CALLBACK_UVM_SV
