
`ifndef GUARD_SVT_AMBA_PERF_BASE_SV
`define GUARD_SVT_AMBA_PERF_BASE_SV
//`include "svt_amba_defines.svi"

/**
  * Class used internally by the VIP to calculate performance. Typically an
  * instance of this class is created by the VIP for each performance metric. At
  * the end of each interval the values of this class are used for
  * checking/reporting as well as updating an instance of svt_amba_perf_rec_base
  * class which stores the performance summary for an interval
  */ 
class svt_amba_perf_calc_base extends `SVT_TRANSACTION_TYPE;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ivl/dU7rzdlTohfxSWVdwdH6xwVi410ekFuybIkG+tNAQGjr7cceK1NCGNK9McF3
uOaoBPkPShE3GxDhwXLRUNj93a9Uv4JknIYX+gciJJJzNY2dD+p3wjYn71hABNeB
Wr63IddWZqrNaQFuISXI+G/08Dfop17lXXgFZacGoQFYaogd7GyWug==
//pragma protect end_key_block
//pragma protect digest_block
mxveVIeY0fYj0rQ8sta5YKtpc3o=
//pragma protect end_digest_block
//pragma protect data_block
vSYNlHTsu61/aphLKxWjuwKECY9LKuaPq6Vs4PRQHhatGAKXdYZyx85hJOp1aICi
7/SEZ5RyNSHxboLp3zkhEjeOiMpzgq/uhAQt9L6EPKhnQsq0JwYqlzh1+71LGMUJ
9XH8/ILHXL1f/+SzfLzO7MUJ67hRfeuDNSUSc+RURekEyr5IEQyYjhcQyScS5lom
XV+J2DHCYwVaRnN63UBmlp1/E6ERH6YtE4kFE9xOLVwFHZjr2KAlNEqekVDXsXvu
XbVPYwclUK6BSVzZg0Azl+yBiwB+Jccw24PozKc3UnLRVVdXJo1uhP7+afLNqcXR
BUBoacFG4/uXwnpHXX5wrWumXROY+9dQDBEcbQw3+gdqAQphQ1QqjVVyUHaL/KZK
Ef/eD9qi3v+O0454Zhpfg004pjEVWdTF88u0T/cglYaOlAxh8OoWIku/fO21m9Xc
HyOiDkm+mLcjYF7i/QNjSytOQAg3qhuL2EQt8PNdJtjhr/Y6P6CM4XSSLpZ/p5QN
uhdNh/bw0N9lT1KMJs/AGjWWDsyDpfgl+pAGqK8hjEdyBuZrfvAGoxpmm5EtkPjQ
WUQ/w2/eMKcNGqIB1WHZlTgsKtIcteKQugNUcyrwRrkktZsfTRZcgFoY+vL0X0+T
Tfw5DCECqj5mO3rD8K6Sg4FshfyyMS6DmPKzBmJfTqyMftLaXQcDGwL5WOMMDqT3
UjKs2bYsUxdXpKJUhZ4vxPjbFiIFOPrS9YET8d4NgeTnuf5jfpTtEzDzzPjDeVgt
q1oQ/0HnIfz+TbM814FbUed8rtqzy8l29cxsuXj4oL9UealGMp2VAmwalhGRth17
NBAqMN91Khjdm81o1W9YhckjUv1Qhe9Tz8hH/5zqv5clCj2yauuuDSbwu5dqgz51
pHOzeRjRDAMDVgz854dnKvBqLrFpEo6mtXl6t3rYuna25NctPGBYke1QtQzUyTci
wDQQPHNYy6XsaBYh+DZqG2TWBH6Cel/6hIc0bVX1j5UF+8bVAfVJCyEEgMF3O4X4
/egIJwP/8Q43Kpwc/0/Hp+9sqTuSSsIHJrQQim2H/TTm6JxG5J72BCe7bC3vVoST
s44LDASVfM0U/5zjRmu7pkBGEpo8qj3VleUKLbGD9pYRDeAuyxlqBx0H6Bqv9i8D
NKH+77FYzmYBInEvG9wSg5mKeH5k6K4Nckcjg6BSG6yRz/7sA8EkjBPrCK0D2I73
7z1MoJJoVBWWTX0hGrvawU9YRY+kcXyl3/m4MZX6208pJe05UZAe/2dFHnmVoPV2
kyz3eZNCB0wO4VImsIbz25UzuNYwp2aIUD6WauFt121dnUmKyNytDTwQVBezrfbr
RHjbS7Qyzf9WVfNGVG9DfKI5rpQye4NdrufFpGM47aaLcAun8DKAbchEOEV1lwlo
DqPn8zlEqPvCAAmyGByZRZZZ0NHZuxYNNo2TUPCayaMAwwalgbOg2HSDweWKGE/t
1cGPDmSSUsqpG6+Vpu1KOJCA6r6/KQ1cXFDxUFPUp1gp/WGBmBXETT0BLAiXytpt
EzqfA21GHszYZi1fYqDkjg7YIuV7joWsqwQgPRiLoR65nylc/ceTAYVAyfmNYXja
2sKcBrN3zkqvaz3pF1fwSuHT6RvbAwkY13YtjAp2O1rlnpBV5y/WNjuHpQ5rUdcj
AEHpO7UEIz16Z2ikVD3hGv6sDqinmokNZMHAUEu/nc1phbQuEUoOZY08VCyNYmsS
0Nc4GUqSx101uzGZXkynRQJC1QGXDBgRQeZjE8eLWubaENI3e530Htu2y/r16LYG
PsnYBrOVDgqbqV2awKNdjoUuTjc0l2v7zcnnR7zTcclZQqrj58sYGzEPw1xMGfhz
p9k4kXrkljEewroJCC2aH8ZdklsAlA3w8QXTV7X/yWe+mqyElQhwtfy3BSpFlf3B
kfGGLkN66vUsuCHzWUuX/45QXFTnnM/imJ+gc4YopS5cjDVuoHa+G7EVoaSaM9Ov
WbhW//gp8aWn+qyM5ceY/LTVUVCodoNfE0kjEyFcjFa/P4jmv01DQRuJ9z/0KwEJ
5P7KxTfk57vbfnsSWvh6kDEVt7PuVXLN6+jLwvEzCIEDrum58BXumxx8PdyE/Vw/
yrNiAWz3sIKYO0epcf3PAKPmGXuJy/UMTJd+xr8f82dMHppIh3vuVvn/BfUavVBs
V86yWSCPbKgYgtjdx1JXCcGbRO7qe2s9yGgRcQUQqiCD82xlUaMihvIXWZVdRfNR
oXm7XQyL/68sFeYQxNDYLWsIjNvE1Xj5/Q3TXvBEnyJgwQ4mCOeW1LM8cssXdbTM
2rXM+lxn3vZy1XbT4nAv07LyrPRN7nccSJcSOa1G2GhtD1NHFgeWYzWDkfcpQp8B
tJBd4S7Cl3zmQR+BFu5vnSvPCezWDJWQVUczq6gbZPBfgjmo/O3IuthSPJX6w2N+
8bVxfbHk3k6t/LGxpGNTBfQdIugGhqt/yaUK3QafpBJI88FuHH/om8Z7CHOmpmpr
EqKwD+otceM+3Rq3yK52jnFEohxI05SAX+YIWuioCIOxyz4hhMcPNs1JTWRmpj1W
kwEcRzt3MJZy8oZV4AT/4cGm+DV08lYOXZW8PJwAB3e07GQ3/jFb9cp+DeMRHq6o
i/OYvPNogU22RxULTaVkvabcbtft/XcfxbMiZxJU1vyZC8A0AvCNPrmTYdvfhWtB
4G9/28ykm1lw6tswtFHIWxJTw28MraMBTYQjorD+UwgeMvFzEGjsUMxbDtQbQBtA
FK+ntNeCxAv0sns9aG02i2W7NmIQ8k3PhWQ8D47bsnmNIFIqvledOTVDCsaACsIi
JEYs1nqNq1IOOGuaHrSXpGGNaW8CHBDm7WExkJg2Jw3uaOLgBW7OjoC95CXTcvkq
MIvEWhb0V+QwnjsfollKGHAE7WAVpfNnn/M5QtPFk3p57J3USAJIcKE/0+TymqhY
YPVX0RhO3D/hbfBhrOWUUtdSkH2Au+AgeXgUbkCkXeUgpYRe31G1Ty0rB+/cNucn
0jQ6QD1NeMuhcAzghtpdb4KGq0nQSsI/5QpQRt/rWopPjul0HX69BR52kRMdiQQh
hberwhDg0TPYrkEbiNTtu2VuFF9v+qsOXLhdqi945fQwB4YxOT0KsLqsh8/lBHyM
WnLsxRxd2zpGNj36aErTDBso8ue0s3jhFrRsKJIL5gpB11k13BiM/D6/tkiobfXO
b0mu1cV8NEaZAPcL9pqw2yoAyfOOfY59ExV/hzX0wr0ewJEV18BCtIDVtuGY8I3X
wSP5L/+1TmGzjSWfs2RdzCe1FFgUWKyuUKfpUuQWL0lAZJCt6biRvlWexn6pCxNk
qmXj+Z6vnlvl4CKW9m1hkuoZkWUQqQRle/AL6a3+hRTa6z8WQzk8436WEMLgyjx6
POMlqSgPNS1VAi3u778R7WyO2udOUZWTUyVNf5fJla70YZl6GKn+3O3875w+fDdI
j+Yoc86ovgHNrTAmWwFUuUF9k2qQv1c4TlQWRXLDNzyUrLK4srT9P8nmd8Z0IY0w
02dHKGz9WNJe8u6x8xbQPGkfNwFK4v3KcdNPqvf2/OYtdbdgSGRboFXgRZoGUhHU
z/0LoujP5EkoWktUeZqiO+bbO+2/pL/DCNO13YrGZa5Dj6xKhSkUnmuWCfrOe9Zn
jKvHzXrPKG26JmewwiviHVes3CzAw48lgDmxSldcnFld55kGmvj4tXnYUy7pzT24
LIJukco6FaNiJx+EY5QMZNm0TEynGUXOm78Iqu1gQnLzJOhhyzvEBUHVG2d12iHx
9JfIPnYuVDqdLWtxPqVEQUM2kiEzmfeW41aj6hWWJnohD4DtipwHw3RmfxiaUll6
DDSveY+AtITkaH4mOAiQdrw5jR4K9N/L3zayxHgjgTceL4suk5J/DYplwnAGioED
xX02j6PCZq0Mi43vRT3ZsB5CXKPfUlCWtUSP/uGMz5skXeq3Aqkn6uLAy/urQDWA
i5c0A3tvUC/OtLpsAekbpkazGKsrK7C7hl95RmlU+ym6QOzVz4Qo7JTdgjD9/yjh
Mgkq/Ef1Buq7T+dX2gKDT6coxb9L12tqCGXKfP0Lda+qI21Rtl5Nqh1AZmr++hV6
H5ofWUKI8DDi9gS2OhwMW1RoKoCH4uINJ5eKYdga9myoC13+pi8x+dZajU5Bbrlv
1Qu+XLVJkDFJlQhilV9bhUdCBpUHjAXlLNBax625cyjIQ2OJvYzXhU18HoDSUkj4
2cEniI5FlHMyoEAVETyQ6xv40m7vOLYv3BeohNuygJMn/2Ct+CE7V1fAoYvuI3iF
yrlAKr6mzFnv3oKaeLVIN+lrhdlbaCmD88HvzrfF/effmLgT31F2efOxIim3XuxV
6PnEEMwSj9ptRj2uNtxyrrr/iPCK+q4lkQ48SVSyo3RmKgUHtuZ2rupuflHrE4ln
2pS5dYU0rN1J7Th3ZzBy2y+Gt+h38KHaFez87ulPI6l8h2hecPa2/oreneY2R/0l
oeAscUaONSdviUM3QQN6NXZCgN/7WxMevLimTKRfvRL/LHnyTpBkY9qLI6KRC5zY
zNqalobsshSF5I88EO4pr1PZ7msZRqWbfeX3HC4y0Yuy91tqlzOSLxKBXQELtkHf
L+6iE4/9+TPUWq+jaWkqnvjSjaB/jqhNtMSC0jIWRPDepSe0VcDqvWGjpclUuAWv
x20LR/Af1Rbam8l3Yo5ZEDobBChbySeUpF+bMu32Ci7Nl0dBtyBxUBCmut2HFell
zCaQPrLfEmKIPbXHhn2VKbIiASDtubg5jH6eUR4n41h4jac0M4mBR7+l94kGAU6P
mX0EW6sb4638sIEIL/Z+mqXDS17BfryTTQ8OITrKsGX1BGa114K7HfF3m1VWvnuw
W+zdj5+GzdpFz5lJItZGzXzMSpBwlfyhuynlfAnIJY5jkHu6cxDzdbmeajqfaa4i
Is1qoJntw2DV3CJqzt8EAD8C6oaHh4KDQUaVpmVedI/Rwrtrk9d61tJyBd/Hw3Wf
0R+C6qRZn5QvZMNDgX6jwyfIi4EEtGesB+kyctW3eCnNF8rlI5VSOYJSqieVkCA/
YECyXM2qFMHl6eFZGa7b0LyvUr/VkJnt5aUWPPJTNdgMg5pDVMQpCBPG3o7Owho5
VW9xeTNqLKSPaj2dgJuu3EKing3MrTDBDbVqhoDBAJfWr/f4vpDSZtmoDDcv4az/
wwQuR5poVbMJTOap2eC84egmxa4+H/4SkzBtZM8P0x8P5RNZU9SJDIlkdlo5GENx
d+Q6TZce6QK2H+MFXqoro3hW4pU+lNaAN6aR8F2gHPg0dOk7cinh2uaP9U1kVCod
EDm6RzZhcNQr6lg0NxWH44yBv9cRYZGm6hyjixP4A6v9AeulN9M5e37h0buq2Pg3
ryw0L4QYjSU4IGhliLI8N/F7t4+Ni5ITLUxsfLO6TdW1omfEK9Iol4IW1C5LIvfd
gFDDCq4cI674Ex3k7UgEZhfypofM05NEOHTIpcmYV0Z3FEV+DvJWiFyioFOrKrqY
27QzY/jHVoYimM/HkEFgLtlLOCSQmOOKvIpjLxH1gjVrKwY++BBXCHiOlx3L/VFV
llWR+i6ox6+QmVfIlXb4rK9No58j4ySb4L6PYejynoSnFvvM22PkiOdcgWtU8t7c
Pbjo86jnA7/7FpaiCMpTjq/64oh+BKsYnKTr5Ldm0g+LBP3jcozp5fE+/1PHQ058
95hYY/1nh09ck5Hw+WeCmXm7oa0ZLb5GML78k9S8Z2eYAz8hu2GNDFdT8ptaQYHm
B/j/Z7kOu0kGtuIc674oyCzovefW7daB7+tbslbCxa+vDkCaIPJD7IfpN6JVYSg6
yr4qJbpn6tWNwW89xrjkNvtolNQyc4Ue/vblKuBmg6mJIPcslmgiOLRfdaTcqH8Q
rXhwUkg6yP+pKvhzTefP7G6d+pDRQcaG++zYe30B0ttHtjBjWRGexI1mGnGbC8uh
/VXR+XNNDzk+vXwpFALG3kvlUVpCOPdhps0O+W3L4s2CxM9hLsaYBNumhnTX9Mko
4b3mhDCHUG1Hy4NwAktzuqU0KSXGE1kLS1jj23a126TkYviYuOVOVu94vuNXj4FU
/ls5Y9hbT7kBU5JCRhRRK1c9H/KCySbFyW0Ed7mzVAo31NNEP1U44TM7xgypq7YB
hRZLh07Q52h6OpXkux6KvQ==
//pragma protect end_data_block
//pragma protect digest_block
AhXoQlFzAwnL4fe1VrMq2/C7SV4=
//pragma protect end_digest_block
//pragma protect end_protected
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
LL2EC8MpT+zQvJ/C2asYMg34rJTjX/Wx4MB+ZGOdgHTIpPahEzMOgXY1oruevXzA
pcgPLYFhUmX1Idj5ArGk74Vpaf8Api9DaoWlObqR8g17yD5n/esZJEpztdLRO4Uy
t/MUiXG4Uaktjf9wzqQMnW45YK5zFvjfo3si/QZ4n9FzfAdzikfH2w==
//pragma protect end_key_block
//pragma protect digest_block
BWZjBbHaOAMaVI5l5kpChvN7y90=
//pragma protect end_digest_block
//pragma protect data_block
fXIo7RH2Ljvnjw0gdNrQ9jx4ebum8q7aBOr/eU7D0XZKlb3qAP7KGTFCxinuB7Ij
Ssew2qxBpmwS/cblH+kPxACAjD6PKd7QzCnAducrz9aEosIqoUKw9fIAT43B08Fi
/m/cijFhxVnLFiuMv9sMcnPQYf/IyTJiTOfuWnWO8KDbvjWudbhNbskuFQA20OgU
S8i3XtoU/VhMY2y0eh5/jpo3CLEHQDKHBWqo+FX7WkQTtSJTAVdLIyPjbzltvb7q
PEgnYdvnoP+UFqarq/AfgbFtD3kpOFFmwoJVyOz3KQDKMZ9LM1fmJ7QDC4Sd4s0c
svRIT50v6j3npZBrbx4cSrq33pKTtAfonHQ2/LqEW1bQTPIlnVQmqS63OtTSugCb
RX7iF+3BkdLGoXHS6wfoOgzy8BZxp7VPEI5XvkMqdYYr3vKI5t5wbGtWt4/r1GFG
nbfy+iNDwoE77/4R54eETeLl9SvP1rQBjhnwB2w/HkUL3hgN6dWk5EtUCc5TRsLr
4tcprAUzuURzNidWEzUDEFIte2bHEycM9Tl5jv2zlBVOnalmkDU+muGD4idi/WJo
d02Z2BSy3neUyGoF/HULMLxFjwysCnnAv9E8NvmNYpwz1GJzovMzLRsNQDqRvS8G
S1aLViLAXIA5qt2Q839lPbC79us4iQg5a6ijB5ApvYbHryDUhqK1JKwWRGDPyFfY
Lb6OMoPtD1Qvhzdxx7R6MtG5gaqjGfoYtA1CjXF46lPuvhpcv12rgnGB37KMLHlU
gNf94xF2PghK6ezEm8ximy58ttOX3rbaK0TM6FgFUqENS9vm8KYpfB9hJ5HIiJIV
BmbPkDXXzefn8aAyiF1cmbIfvjMJJLCL4X4anhEfy+ZRsTFpnIOem6TMYypPnLPi
fOYyfw7Gw9lgbUADa+eNZJ910FP8nV1NO5uYKW+kf+9bnM1Dhg6hiwlIZ5OaS7ag
wplyz4EWbaDZ8a0hPKTC2dilABrkyXTwqWHbTCDYwNqhZZuGgNHJc6eRqRNFOhwo
4x8AhETYMsUCy6kjfxjfGzb6FBIMdLIC5T4edSMXTcH/uqbgCOPl3NcVkrtoscZy
NPYsNO+SJXodiiHmSIqv6+zaH/1FOa39WX/UEr4Dkisgs8pe5OwxsQZwQzdaVjAY
J3NkgcP9tY7uDEi8FUTIIwZdWMqYKQ2KbD9F0qXOG5RpWeo9T20brxtdcTTI79DQ
eZ8Y5KhaUFYb4Z48LDhH5hZFcKeLGM5+87Rk7+K9TCnY0acFoWzzLJMRUXYOAKCU
LOYK83NJbPW2d4aDXMTh7hfwkB8vxBvCKbYNXkhxlNaPYumxNzcUb0fPgjpp6qo0
GP/4NBvUcZurnrWYHwpvVC/CCKM3fd6MndetdK7gSYhzb93yIGYOExaUMj321PwG
K25jQIjZcgdvZDGFp+Nveg7zQESd+OfR97zP82b6s/ij2Hc/5CJrW1VnQY6vCKX6
LaohClXp/0Wyob12DgI/TsWo8huFCCK1/JCLNxskaGayxf9ThABe9Sk0AVlYVvhj
AebG+ZTL3FqTCWzMw28QBYKMZHWhv78zCQE5xvrA1KMxaryLlFwJqeOGIN+rSsAg
DL9l13cqF4RkzZxK431mWkfhh11EtuWZNGHbE3aGyYy8dbJJaDr3KuifEoobCW9s
rj/kqIcz+AcUr0K3qy6Pxh3SYWWCubUjmnN0i2ejP0EfhdGXmhTRcptWMDoQfV//
5GGtCKuKJBCTmP4qw2PnizTHKtGYNX8fbRB6YJF1Cc3g5h9l2sYm93SeDQXaaAOV
77mSChATBkhcy1MnZhSKZl3oH2XKnBjZJI98iHIY2DUcMtneObmmsKy+Wn4fuyeP
tFHX4njwFwTFyn/wZ57gwbYNkphydsni3ClPSWpn2KgcJ+90ieZDy7EZgO+L5lxe
0dF54OxAN0tq61QW+RoiAz8U4p6PKjFfIYzgIiLxKeLEeTCalD+RjgQ1woG8J1n/
yKLj8MXfqxuYEr/Bb63lYeDggVfazVhnchonGNDlbU6+jaIwkeWSxgug+FaYXqFw
y9p4qaotSAhlgqeqjKINVvJCAteP7GtEbKW7Of1rHIRMYUjdFiXg4tCRVMmQgVdz
EWvngK3gSh/RrRXJH4E+C1VWwjk7xrqnWL4MWPA6GwgBsDftbJEjsDC9vkAsM3w2
NxkZC4P9Jd5ORdXid/mYjbJltMtPaw0h8ax9FW1yxJy7S9gUlG0cBcUuIJANTY7Z
7yH8aFu2vGZBkLCJirl4zirJWeLRxtKUHDdrVmFQciCCN1sUs3SMoQ126s/1BU2b
uRt1yXbky1KEiBvwIykhlrujaCa6SQnMy2cHqjTM1/j0mwoZfVui0268BDsK5pMo
QbczeixKC2tAud7WqL4VstRHNlPEbi03ahoDAcChAoDoiBscwyGTi9p0tVsgoR8k
xZGnJdoG6Qw5aWPDTNFUWBJFVmwFPTBVvExjbG9iD7HEOM4lB+D8BdDuF7UDJgvt
NN3O6MuLPASuV0RrV9+aAP7f6l1IsrFDQBEylpPdpgYKT9kONsABaZYT86Jfhyox
TSQcD27H+6PDpkhXJ0z2jq7nBMWfjvsmp/RaTMkYPOEkVYsuRUerN6kgM3xSVP2p
zuq2HqyaFrIbn+UTmbkIAPyGrbjoSmAWg44acS7AEaFvVSaM81ishHuehCDnPvF4
/oPKO8GC7O53JLz/QB6ZJY4aSnAMjzylDXmyCTRaPVKGFvgqDaqwXM2KYdPWiR24
y1iyRhhp0Vxxp01diDi7ENIVK3BBSSZbDMQf4kvIOYNhLmMf4V5zCLqKZYNeOWxZ
fbGV2wHluERKWqtZQxL3bFbc1BPvTzbfF0OUAjruogGpOTfRN+v8Fauw2Eitwy9+
rULTmbifpqLTdouVxFrvkQylpfi7kAOQcVvEaUQf3Hc5hOmM63RbkzDx8lpZ4eQP
mj01R+PYe+mhjIZtOdXjm89kz1sLFOMkd1B7cBgFmvNev8LIHbpahhOa6Sic2qhZ
Pc9MMlmJNKgUkdb6SRlyQCaOwqpYmmpoWLtric9t/g1jkOmq117nwIaLcfbNETxa
U4pVnlXuIPDO4KPZ4OfMVATHBzyBoKGvcxQV0HN7aCLwVp3yImvA/MI5Qml8bZ3p
Rr1eJesvWeJ1WFnQIOgxPRN9z2T9LCVnZiPdjQtsfPVFrKWVZSjSokLFS0ZdwuQt
HrLtUfXVrhN3DVSSxib7jQetH/U95HrInK2ObSNLieuqCUto81M5frgS1oqVyqpi
pH7myJiV+A66A2YyhFWQiQK19q+6icgTuVsgR/tk6uFYAWewhYuZjWgudvShfuMp
TOjY/tHv8DFzFE6E18mlNqNnLdCA6zXn/U4ebDT2oifVdgbmxQYIWaMoiLR+gOgM

//pragma protect end_data_block
//pragma protect digest_block
vdHQ1bq3gdzc9rUuPLSTHVR2F4Q=
//pragma protect end_digest_block
//pragma protect end_protected
/**
  * This class records the performance activity in a given performance interval.
  * Typcially, an instance of this class is created at the end of each
  * performance interval configured by the user and is updated with the
  * performance results for that period. This is stored by the monitor for
  * reporting
  */
class svt_amba_perf_rec_base extends `SVT_TRANSACTION_TYPE;
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
B0bTyvm061rY+qQeZ+HSuBE7Gj8YzyRq1mZmjjqq3w8UfCG+35jkMWv3vADjcT2q
2EQMO1umgLY6VOzbXI2+DL4mnOfxOJSNAvKnOxweLKP5E5Ryu145nkXemZ6/IpV3
WHLzg5FhjMd34aMjateR97aE1lm6OpQdu1VedlkTxFJ0rF4/Fwg1mw==
//pragma protect end_key_block
//pragma protect digest_block
3FqUCeFKYQ14Ny97OBFl5h+r7aE=
//pragma protect end_digest_block
//pragma protect data_block
64u/+tFVRI0xFlyVJ/LG3QIUuzLU0UPIIFPpbIAr/9x4nOS1T+tFFseAyG0vXgFl
1lYIKTd4LsFf/gYkUtvqtd+sPh/bMUc3mnILUW36gQJhuK5LK2novysDnAHGlmfo
JJY4Ix61FR+eR98gdadLGEs3lq3ILTXatDRfUIiT+wyy9AbFxIsxBaIyKTCtcUw9
x6kj3LHLtSw5I6ZrWXrASUHHW+vAQGqPH1nWHGeyvIlDaq7iy5qrbIUXAkUeCcZw
N6Mc6Iy3mPdkcSsPTWihNTq0qu+xxP1uzW7K9TIdMVQewfuHUPRa5nzOahEPwdOm
oDmQLiOM9EcQiagg8COhlx5zIvKdoUi4Zh4ziZdzO6rlPx9J3x7P4pef/X+DAzZA
iDq/0sN9fGvEzPhhT1SfZf+UridiLqLU4iKlnfxdCroFGCJaZVD/iT9oUHIKL7L0
8xvkyLkGZN/EUL9EghZDM0zdRds9VxXMkODp95Vfjr44Y94kZjuEz0gy63wjStsX
jy3Yyt0cNGfUWBdbnfLKplt11zouQrfEiYlQzBUK8b3tPnCbuyklJBgICSTf40TW
xzouVoEpTqFzZEGJ/axgjIHFIU0GDSFX7OMAWA62h0I3r7idqZegJbOWf6M3Zdu0
ZsF7Bs0NNiigt9HSm6ZKqrTqjtxfl2RFjOO1uyrKW6+VMWWCROv8Pw1Xx3hCd0JX
5Ly5Z8TvQ+WyT6x6beJNqStZICE250KOvsV1vUHtl2KyDO+PyLmgs5e+BjvfWLb1
y2QoBQ6GusGZS88ERM62a/Jfy8Voc2YSI/AlwHEFPQd3zEnA0zs4x2GdX1OrWD2Y
XdFzxBLp0YyB+XBu6OYIJ57MlaXxyEtUPvSic4X2puCe9mfTMe+0/JTQR4alU9uh
A90sjNd9BzTypLHOyb4Mh5yGXIZhuqCXx7YaW0iyCKoAWYdlkDF8VI+wr7v509tV
qBmjDgaZUnSdy5phFuZO5Wyw+STFq5mq0cN1oY8vAhwbiysp/BG9X5BNNEQceT6g
rg3qIm+WwgQD7JVmijUEEwW50Uf7U/Ji7TkAqWUspE3wnfR3TJtEkjieb4e9iHT6
NNtGXW5tn64DMBQ/hgBQeSsgneSxVAFuL+iR8TL+77VBIgllxQ01SzTiZIym7ile
eX2mzYC0fRKLU2Nf9kGQoUEt2PtazUZkO8MS2uxugY/YCQ+D4iqMX7zeXhtwaqpz
Z+oi4dp44VnsmkbzLI8PkXEr1f0jx8I93i/uqgZu+zJZdhb6rlL9Rq1ikeJq9s2v
NgIwyRBKo9H+D9ClduFPUA7xrer8t0+Kc/1bpT6zZ7Fi7KT5K+ZeyEHDw5BC7HU6
e3sPSVIKeVPCxbkrAQgdlYkkNFO6M2ANy+WsuzqttHgX1pDYSLamuWMiKDbAhkcX
FRkyqjnmibe0Sx0+uITZu6OI8IiFwohK1ZutCVXG6LKWDv0Uqb63naCEDROqsdxr
pvMC1NqqKCQ5BBsKozDRv1tRCUQcY2gzNaeSamn8bq+XzunBWNo1arprdT1MjAcV
iVGo/UwBElCWNvptJXKAnZDCOR2Lpc57VONXLTVkWecdAG3VR9I7xUSWwAXUsBe1
aRFabuhCw6zAvJO0FLFc/o8HLMl1zWlCNHCPYsrWirqkNPaloF/7bI38qFcac56A
OoK9//pARzFGKx9bOUNN1Ti0cDaQC/fLLgTCPcDkbwgiIg378dttw6ljh3jZtvOk
aizYJfRbVzqyauNTUF6xBhU2y0Gt7OjaZ33cjBABJAoJSU/KTPTa3fDlaFVivdY1
iY+Is5vZCsKrybI6YeXUGZPgNMatLPwafkTPe3FIgDvJKQbk7JoqqTpqmwM4TwQX
wooEtexUHyJ9P8zNs62nOcHaNKpI3REdAKOqelWJN8+garcwcVgfAu8VSzKAxCap
hvevAtmrbtjHTOX+ObdpVhi4+hvGGwLU2oJKr0kyagP7rUZomT1WWtv3kTMnO86m
v/L78bvjRQ98Rffcr+av15HSiCZ0VqbfGEpA0FYlNDaB6sRngN0LYfSfp6rPBADQ
gPRcrMOgDtpbejA5+uGiWLmfUiEAk3WTHGoFnixYFdSUJRrLYdx5y1nXSD+9LGob
2rJ8g03/graj2Y5tvRAjtvJwW4rtHsV07uxv6GXcBSSU7HDtQfRoNT/xVmLZxHhr
sbipi3bQmjv/ujMq62RnuZ5UonuovL+8XQSz5LjWu8To1OYuZrAIclhBhPq//V4A
4jOJeZxdgBMp5CCPa9/rTHA9ktzklfqFQdUqUGcSGUoBTqo9wv2qrskghiatJYlw
95+bsn1Do61Fb8gzTd+9uk1WggXVL9usT/ILW4yBwpoZ6377WRJYAORBOvhNlMDh
BgQuRHItCLx4R35/fwAeXYamnViU12kog9QQ58QHh6aW64hIBJ4OBzXABhcBSXpS
kcDOXS+6C+tsDyTapIo9WaGK6aAYO3Y+ZB336vexffBxBv5QUyNM1/qb5Rv25kcG
FqE7CWNYI+pUE/T3GKlK6lxnryKSkcMRZz6ZZlJB/OkZpU2vW/CyhwxzCqAXFEpd
QuEfGFROsUveyncZ3UrdvGL9n6nUKcAAWGiRaYQfbL2Or7ywS29KbJm0mgMXR7+w
qwGeknV7s+UMfMl0mAGEPd7MyMOmeaTeIWO2G323MTZ+s47dgOs1zwNPpEtmYhDc
7TsElgQ48K/s+rWql5XFAl8SedN9L3iSTshKrvTNu3wrGtCEY8+Vf1PkOEpMahfY
R/3XgcR0M5QgHfH7WA+KYjQP13MbQJpQvYSvhe9fpAFfZb5PbJrj7lJ29qkKNjML
S0UJ8HXo1//AMmiTrkWSzQEw+jQ5Se0iVpdrRHm1lLc3XLfcJds0S6BR4OwZSCGy
gN1v2Fg7aKIKv6D+Csp4hQ7Hc8o5Tzaxr9SVzHTPyYTAGU1oYduaYMCfh9Ztnp7x
uvSX91eFW+AFVxt5rzzK8FwRouMxcCcm9TZP4P6STEevDyxClyNT44SkOr+lGJhD
PJdYBf6vwOLDh+tOKuoAtbAsSCmOIihrt+ukwd7xcjlmchpy3TY7vnCKm3AoCYsM
4yoa7/HhLFQ67KPKv868XulsMJ/nQbt8KokzO7ePEFArCoJmvSIklcn/1GMcSnm+
EacvtWTujgfjWxtyAjqjxEXxfIunxuy43Qx+rNyt4+Qqnn/80L6O5HqhCSQRUYSX
oC2/5Ln3WffXyDaas6xJh5TxMf6NlR8hcn4tr/PW6SsvbZn88mIrW/gVNA/ugIXW
VhRcNpX9Dbe1/PYk58qzM1fNacVOAqJ3h0cWBmQsImbJ+O26YOAibaMgaF9jmkHP
xouqd1dx/3h9pELeBDs4se3Qd1bFdMOa08a36AKk5Y8BcyTPHD1H/rE/FN64xXvH
NTurCUcBrO3rXsmBecoAB+/o0tcwWwF1jqFp3TCd2uIAH2F60HFnODHppmDKcoMi
r2x++U2vlXO25xEKGHZzH9XebeAcJFOxWDXcVPl3JDaFiPP34MTE7Cv3L9/1NcHg
gp4H9LtTP1aR/h0AqwvRw39pRDuoL2dE0Nd22BkPsczJxIHdIxpC3x8+25hir9B3
k+IN+32VIFkGRXkkExnIAWqkKYcykt3wGd0D3IENQ9G18vkWgxYt7Ffd20ItEWcn
92DjhlxwZBUo3keAdW+RtG1a2a4soSDSZlMw11fqheVigBbg4d96a6LfwRrAFlmY
CmIZCoPLA23prB8jrpMAMIhp5UqucAK2SlITbeur/qkz7bRwzeebYfDbEdiFtgCo
r9a5Q5sbWpQBaX/3FL4xd8W4+O02FaFXWvpl7C/MH77J6eaNHUiqDwrArW/cCplS
XBa/aGvkRIdpEr2NMH6XYaARdTZL3G/b5+x7WmNRTFamwNAW60W7VF63aOqBnJHQ
jzUm/mxKD231+dKrzm/thtW5IrVUkoiCPFmw9Qc7ZQEa+YXgJCDPDxXHRkzb6iah
3zpRu0xk21mpjfNmVeT1aEocoSRU9/RQgx5bTXVtp9mdvZpILswLBhGGlo4EwvYb
wBOekXyPdXMX7kPkYSI7EC5gjHlUyZgnDUXf5Oo5crUct81hAUfDAfvrlsKLlrkg
fkv/hZ8fgi6QehQEHMe4N4lsvgiT7rc1dHqmCk7BCkhYMySmfmW/yx/BnHBeybY2
E8Uya9YSDul6Ouyix7CQnhzodIrUwAOVgSb3v2Nleu7kea9e6riDg6TPRG+NVaP+
ZntuC0gTCPvskpFL+6FBSVypxv/Q7JX3v3YV4lwjgXkJRkUnwglbf1nPz/1MIQAG
U6ZUcvQrkIBgTyuoAyupoWGf3/RkyIJiszAA92empjjtVo7PSOFWep59sG1lvTPg
5+NwTGkkJgwhf7iF1I8UCxjrr38u3AmGpt0is1DwdFuxI/R+NcuQGCO+n48nCfxe
9JBPOtWGIbBn8X7YUBk4TyMj7LT7pPu3y6QGh8A1hYi8lEsMDYhUzFVhHmNQkE5h
q9d5ZOAmqWNG5O9ws90qupcCVacGF+M4hnUM1mTvhyG4kycBa9f0xXRpkiVaZM7X
6s6jVyYbXVcT8AbUmwGD4F/qKh6qKnAO+f7PMZEadtHBtw+gfgz5IalObrxIomUH
bhMjFTWYWlVYKQSKItw1aNtOL8/fSwVlFyCUBjD2QReIUSbKbZRw4TA8OEV+m5lm
fAaJmqoUY0RpdXYdjSB0i+rP//K0as5f6UfKeHOLgFjowi+Dgsnvy3ikt1ii858m
mxNqrZxegzvvTDPtFzbj0Z6r28hJgoX9hUF6oZvERq+oFhzwNnyqzW7iRFikwDhY
TTlatIlFNbbIpsvroEoR92HlXTAd9k788Ae5dnlBet1IpV1ftw8NRJq9C+3mmKJj
/EhnVV7AFSm4zOM+dYvimBymdYOIUUGYlSKWMH1ljouu/D8ca9Ha6ZgpOL1chySR
6Y5XmvI9rLJfa06YJB3goVz1cnMjJY8k0WuzQrO3X1mtZbgPt+0VTJY/loc7ptQx
I41NuJN4caWn4JhhsFOGFm506XQZUttZeIJ/nM/a0RBhbrZMC5IOgKxkU1Jw3VLG
13tjakGCsr6pUxAUgMpUOKrs791wKXw12VEhsWO/2xNKjMQLexHz06Pg/wHqHnpG
dZEaLuVz1tUojuj6uYnrjKBgu0xTjMS+0PXXJtJZTTWqqMp4x0uyNf2qpPJPAnJo
KdOxilDuJKgfrroPOtqvyGmk2Z5zLdIUY3UVigs9K8NC7bckvPeNf93KlTN8u4a4
dWFQXFjj7lVN+vT8wn6DPt/WoP7NpLvzWHfKgDUi4CL/NPhwFrGgXMuYFv9KIA74
OvMctaC26wkTEsOLK04Zku7BBrXkALDfx6om44UGHEsBmJHwDfKNQtAkSWUxtsq0
YFynR7yWGF+JRWcGLHr8oQCjEVQqSLeki0GPg5mvivRih7bEEjzrdJTQ/AHqNfx9
zSFmPogoEjNBtk4uvcgt/NeRCLF3J7HoX9XC0z+2NekH6k37CFUWQl1amf0t0stU
UjK4ypze6HGTUuH+fhY2G91G22HadXobRGzLm3RDCGC/Wcot/zQBJQGtkQJXR2L4
hjiBNuNJvkZz0x/n8keC+9yu+52TkJxD5mFh4llIflOI1wv2qyr6Mbbqmkgj8ARM
jmgeokktmv1vt4QuNGpYHe4PHomBe+Sb01a4F9FCRIOpO1K+2G88iGDzKzeIXyCr
5c6hP0Q7tFaCbugWNngKEQxafISVmpgfhPgKXC9EPgqhwPsZZ4eDwkCDiuf+u/le
857f0sihTEyvENw9GAXtVs/h+WjmlVD1dmc0HE5P5GnbtMJ9tBeW256JP7UBy74A
GpX5D3b3mcLAFVyJUtEf+6Ly3Dc+bM38WhPy8QCvhmTK/mGopYibcIAb0nSOciNM
kNm99dqN3vqhek+PNyxM2Tq7m1juc8I0A66wPhwtWN3OuqJDBXF5Sbkk2ZRP5jKa
tp7ies35BDQTM6Lq85qS+jPAbNZ5CFMGkTEWLqfAjlFawspUFZK3dFnXZkrZXj/q
TehDTAWUsQocAUz6aaHTFcp3FzJSNaluD4j//ui2D6tAGyjdGwPotRg5aRipSEsg
cDx4E6hyoyxDijTjTrwRBFokqdkF58eco5eHd2hJiPERO5Twel5/LM5FxhXrf26S
YEVQfqur4sLV8xFwojakC24ZoO+P6kzx9TOevODCbPR3dxh0vlCMOzDBbMSpt6PD
cMasrYsW26b9LyAvhzlXJC6tJ3oTf2urAtvKvu0mUahm0h6M0cvqmXJc2+RPiLEd
u13cb9lKrzuF9x9+fqyQpowfDhYXyWW+KSkYebSmxkgX+SoGvKFxivWDL4VhXZH4
lu2Tw3EL8kAAFHZxawtaLmwNX3AaKWMh5ZrtfENhBuQeQ7weu0yuAPF6YnB+vj2/
dXWV6khmHzW/c8D0brzG2wkPawrtu8DMTcHx1Wa6G5W/szSuwZMS7ApRIK6cAL3p
A0m+ii4mkapRjvisJUgMdKIYrbTOZqArRyXuOSFNAVeC40xlOrDVbrb0ZOubgsX2
VMAfwKbZ5snB/nxfqMwQ6Qe0qCR7PBhQDK+uHndSUMsrP5iMzzyYUYRJ6sJ4vBqB
11ARaJ0gIGowCsuZMfwTu0Efnh42BFBfztV5s4hhzFupSK+GLWPEnh24D730Mal8
Bn8FxZspELU40hLJpl7ct76tGh9gBjzHmbFgW4kKVaMCMVfi9GLnp/+zWvY5VXZi
Yyb66mH7YXOv3AFtfQzoqGRsC7stsZx5nVJtjkxhcOxEBITcmA40TGT/AU5Qr/bO
8W/6ItV5eJ1SHzwajc5alY+0IMQceQERKTtJxBqoPMaF0kqLOKYHBt1fYoqZlBbW
AdaP6UOItMf5tj7+kIXZy7WdWzrzPkJht1dLj9JkgkVgCSxNHq8wUJmDvy6gz4xb
Cx7bTDKt7xMXwB1XgBfiGmbL1fn210jzVuc9kh5xBp5yBQTgYFRy1kHxIRnBTpcF
3jTpw8LVhnB4Bv6HMBPYJLCEZ8g/KFh3xrK7ufKfVykgrKSg1uSIOn7MRvS5J8Dv
+lLW2i8TjDfQpD/IyYFuFjASeECNNoZkx/Vt3jKkgKnBxDxRnf9aTkfeSafTMZIL
QL8nkFcYEFgrXBcTJRvaxA53cUOyBzeXqRI4UF2XaIyD+L9N2ciskb0TIZS9K0jR
Ef4gl0tEVu0dCKAPk68FPhopY6vxVBT/GJARJeCrP3dA6gxWcS4v0/LOJuhsBPsI
3NVfwPLeq3Vw4G/xSSGMibsDlbVILdysUQdjcvGe7uFrt/TwaxktYVJrRL/T90Ao
URV8waJoK2jHJEWWzaiEHzAsrN8lYq06RB/5JZSUTRdq0RXDwcq4MDorabEK82aB
6yFiqr7uRWqtYw/zeLps5M8MEcC/Nf5yXfzHWfHkt6iQ8iH1HU79oix5NDvNOkNb
3Bs3KVEODrHuI6vmHlK0B1UVRsyp+I00qk7xEu3BdKarxjw4FVrZ15JpkPcNjDWk
KkpEEPG6g0sfS+IwVgFTXbk0/A3RK8+QrXHt1LincKMoCQFzEFINPo7ndrQcYhmg
6h51ObePxmInSl1BmgoEYAJ2KHmA7llzF+upTssMLZstVEs88rlo8rePdJpv7wWB
1p/nxr6/g750WXTGQ2aX9OGMomEnf+XviZYpxBfuoF4JTBwFvjTSEHb+8sAr1dbu
L4BuN42Fec5mq9etQuLzRo2fLAh7bG8NDfNMjmEBS6ANy1++ifikYDBU5rvO53Uu
GusA1XjPKQfbV2PaQvy5xPoEiMFbG+qBPeQKT6Nu4tQBRb/aaq1Mudp7cQWu8MrS
KS0eJl/zjz0CUuqOyaSd2L7ZQSbgXyaIjq7B0AuXJ1fUKWONxH1AsJPqO2motBrr
5FNAeoU6J0AMhxvOX3blK/ETQKqF7qjmGlRneLnKLFWeOKnaJufTkv4Ukoe4hWbi
iOlueeztQAFPytID3am3gkwU8tmYiI2Ob/khSJCZeK5sbwd5EQrCIfArzY+rx8DB
gNlCCkIL9y6isvHdfHdqiEd2WpkupzMAhiCpSvCF9NG4tbJJx+L3sSlFR8qSaYqB
Tf0PqIKQUmJWMJBk8zihINc4ZZVv30z5QhGW7X1y7odeR1IgE+XZFeSgBIpj6aM8
75y+arXbGstHqfeK7ifnegJwAyom3LDRT7XIWD+TGdBSM+rGUGWjNqO6e8tGT7Xw
LZRUbir3hZYKrQ69mjOYE/GgafMXfM7Ge8RObPy33iH9JfVqG6NyUwUQvcFinjc3
tnECqoxSVzNL9RwhGlOjFwL7wlR6vu8O6rmgrGEyXHbvnMSL8AEfTdXqN5YMq3Cj
vcOQZJ3yJ+K5SBsdMjGOZ8LJBusj5CFmFIwjoTNvFuz7iiHCchB8lACa7dta8E2o
vIXVyJk5GBdYqgdFn5TQP0CwvkPvMTLY76ML4Nqbilm0nLY/rN/abTh0eFL0cdfu
tZPQ/lcvhXYF4VVDvwQmRcxHUBRO2EuR4V2pk6+fiIl05ewtmn/pVnwZyvZBxWVR
fRwrQcMULnnrtbo9EgR+NO+flDZIVQTH8p+/Nn+zRo9uKY66kuPtq7hXJPW1SJV6
TO0aeyDx4u6rai5c0P4aHLfF1pKYJHUQxt4a0u0uSQ1vzer1u6NHYfGAvkGFArxE
sW3A9q5fiEjEz7puRGHgJhN0B12piUpkv5ZX1vhw61pQGLoTvmN4rkUIXiHQR2ab
GK8r02E575dCJcwf0kmRIsJTTfU7Pb3Rzo8Y9/j0wdiXwqBBOpg8qfIfmqyuUMWg
jzdfstYCrKCi6RWejKSY3AdtdxyG9wZ5V/GvmnI4skbevtzrUOzZjYSiaAJJ1zZk
Z2QnJ6cL+/OS//3/bEd1+oGGndxYHRQ7g8jODvoggZ60Iy1DoGfdnQrGXOQAyxva
VdKAnzC4bfqIav12AfJZNw9+K45jEXp/AWErMgQ9pIaNhF3YAaz0U+hsMeoJt2CF
v/xoQf/QL9c+iefqJXDWYkImfHKSwvVmvE9BaTDMnVJjHXubz35XN7g6CuD5J6Lx
//ehGe7CH/Pug1uVyL3pdabzK48iCgJpQiHPywjYAC2+GyAlxBnZvqBD7PPQH88A
GdoSVvfV8DPc8PYz5eBsaP13it6U2+9vWlXpV7NLC4GtXzaMRMGIOLfknS2uMe8V
8gtLTRQXit5K8wZdBNlCpHA9b3eNSYYNXhZErVPnXtl0SoFg2flmbLh/5843eOyy
t2Ad5MNmS/TgNYS40Ugz3ryK1caz91qRU/eVovC73QjX6GRmEu6IcbHNm+3UlraZ
TRhFGnhUHLm40lGy8Xb2gJL018f+rVAnkkUUn7GsxcTCz8FeWcdzFC4RD6y/xl9f
sXuOYHxbu5JqTHfjfVnFHcldsB6/+pjViNdOfIXsH3N/nxpzSeoFfWW547QAq1gB
s8AnXbkaPf8Z/Y3fsrMj8l7FTvHk86HiiaLZtKYVJM3ugA7hC7hJ29F4fluQ8V4z
0leWyKc1/Ib/tUkTjIEZTPbyDqPNXKrsHCZCcANkl6mSoQApvZrKLMgiMl1T0NOv
dy4xxPH8yAcwN0chQz77iOLGw4CjIGD9uor76k8Z6RsI26oMkppTKcYEytkKMRx+
t83rifhO10if9VLiNLq6lv9bqAk532nSo9F7fU5yh1s7NZNgabSRIDZH8yxeF2Fq
MflaBIlEyq3yUpRWZYf8rn6jYrgnicaeODODfN5ZD4Icw5U7o0RMBytMzIMq9D28
HxOetC+H1+PP1u81Yi4OYy7Vcquj3N15byrYCb0/0DxOb7AomZLhjMhVBVDR9jW6
evAfukunZmzP5SHGKzJ6MkNbHNqtxIpfm3HwuHsenu7spfb/ifOWO4UzLoYW+rVA
5eBQsCLuWesRXhm7jmiWAiJSrxVDAdd2zw8GlVRTLwyJrLplhRwYPi8bDDxdhSi1
I0ckrEUH53l68fdyBjjE1NDOV9MAmJuWPZm8iG6lMBP/SwfxwUKFdJhfTvSx5K2y
stM6ZCTb/ou7XnW6vFArsOeplK8Az4pgNK/lCvDl5oAZ7i04indrcALZsNqj8WBr
fPon7Vbkj171aXlq7PkxsdwF0dEWlQOJiKlhLGZHmrOfMV+RyUk4FRY6je0CF1Ui
XgFaqNlysT1BkhaG35V80P9ETTqG2NNYEZ7JKGLaZmZM66ropIL4v+VdVU/JQ4DL
A8l4/VH9yAB+PZ9mRvShFd6lBIMjVJDzL/xV7M/vyk24WthZ9Ozk5FyhkWZHSa+r
IlbtA5WyzEzKVmd0RXBP050OdLpXDenwpwCKqYYPjth4kvzU9a7PqK0CubbX8NwU
Adl69jPevjtnYsokRzzTDXJx2EyXvXnAHYSeq32+guMVswUOV80DY7XeYb+F2Mc8
icChgB0w/OB3JHp5xiidPOW8TuwcWoSMDQAG2xNvWQ8ehowohylZZ8jLSEKmA1Bb
aEsC10ptSq3Dx/5AegrAVTkpJzEy93Aienlm9Sg7xd3pAbMj2n+LKhhYJDMM4qY/
AgJajHzmWpI+yyS4Qi/xC1Dd16H/XHKeBEjkzmn5nNwAAuLmEBkXVUkl8u1LXego
uozX/nghCx280JqfjyGOBpzDGb8dvo43OL7xKopy20xvAAQSWu4tSlK5aPWl/2i/
IK21UcmBwBQesIIgvx5oKjVcEj8WxM8o2siA45kndlqNjep3qECp2o4J72T1ayim
aBUAgpH5VYOU+VFw65nN2+hyi0Zsazdqmn5fVCf6TMU=
//pragma protect end_data_block
//pragma protect digest_block
MsdYop3fQOkILIzJJqXl4IVcAps=
//pragma protect end_digest_block
//pragma protect end_protected
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
aZbLT9yrBiD7sHF0nmLZxatWaYbbvRMRavCTKfJNOTpLItgbS0++RuXD1LvzcUHW
Z8SkDkSXLHL2Uo2wvCRj93slUHpCmCjALoG+ApURtZEh/sx2yu/RnIfUEPBCVvdH
LHTRLcPjEMYwIUjf3s1luynAHyqDQZpIXyBR0PveMwJROjl28eKy1g==
//pragma protect end_key_block
//pragma protect digest_block
52R+hFbPEuhjswBn/Nq5gI7SWPA=
//pragma protect end_digest_block
//pragma protect data_block
AebPRxVWRcdFxsxc820/wuxlbi82NlygooI3lPPZXSWSJg3eLLuLbGLFI1EcsFVX
DY2smNc46r1z0YtklMnnX8o53DJ4Xf0l7dkRPlsQ2P0CeUj7w1mCsASfNOgLZcjt
NZifmjt/ep4IPVyiOsM7t8bq9rO7q3kE3BblMjgnK/M2gIH5c5R4e4kiQTgFij7F
iUoYJWatw2TFmltl8C0yUAm3buQ9Tn74XTpqbu6n62L8HQDQZW5ej0EJJ7ScqyN/
Q9NsHA7v53y3XRKTheaBF4s3Dnj1gyG8C6jCdI3tn68Q7qcUaZzDO2VLORhF8qhS
mP7rh1ghEAxtTPHp0A+zDoUrEg/xT33P8G9XCtNRZNDu8JUuOzYcxUy9cRJs1u2D
lQBUmGmaoqLlaj5Fe5n4m+j5p6mmOv9y84OyayYekrHah4NCEnqmzUKeaW2hSAwF
oNSJHdHntMoiYz2ssO/qKM+mxQuaEKchQKyOk7+H2MWvHxV6jPDBZNbTScSYlBMw
lg1Wfpk1bjaRDXScqw9l101nYDq2FEUkRqbmVEg1ZkgXKDryqnQlFSHxyEfPXXni
ankGjiaAh6ShX/rivDUHz//Eo//kuJytNxwgLfN50cX5dSoGLZLrvgOHOLioyKfj
5HzIZMiqQz098R+iC8MBUlTpG0Y9QKNoXUuUQpc895lSImtjlje0oT5Ua5Uq2yWw
gvkS8hGCFdMRQzL9bR6U4ZcgYAm1lMNT7J/cnQE30x/3rw+whOnRoxtoUz8JVZX/
qNykSy5NWMV+mPTGh1iHTdJoFaMYbWwkCCdhBrj07HdlnXbtJPlpkGW/7QuUjHLd
cMZCwmCMo/jex9vJtYqW47JecjF0vogdW3EAQap3QYbIqdcotaRehSc9BjVd6EMn
DPNJZYQN4owGAqWb+UhkhgdexX0IKiuBDpZJCUrkzFv5PowqDHe1BGXXqF7dV1EX
r1ajLI2rtxj61lX9Iu1aZ/C8h596gHin3ms5bmm+leyB/hQzT0rtO8+HiLhe3zJe
z2sQcXGjBCaH+CjFpn+/9qmU0dzj/mDHTS5zchEX8zhSa8glm8SOBitH4K8am/uJ
lxjrZKx6eCn8K9Nfov4QhHpv8LTY2CTFZGFptrTgliffNqvvrvo7NqpjgAAzNK4o
eQEm/wpgrU2EkGKr5mPNaBpGLhaZaaqGWAwwMxFfElQtMchjVmx30C0HbEWZhfGy
xtUAZzFddVCCiAZjURI0ThA+hapmyXE1peD2ffsBK1bSyxozHqZ4zTbaPa5nK7Nd
M6BixRDsxnWh1PFiZ0kYxUvZmMPpGJWrMpg2yIUc498+GNzKub333BTjdgFqLhKx
OwEAPpSQmNWpJ1ryLHuf3RA5Du+Y1+dUMSGeiUMgUY2VV1FohgX2ZbXkGuHlNPY3
pjeNgAGSqD8eQZVGoR0x4K58lVw197z7N/S0ALQy6FuouPd1ljUv98zXZCokTGRf
H1Q0S+LKI7CSwNN+vTxfS7YR84ULSbVX2rdyNRQ4SUm54id6geoLJ2jG1pODHtjU
yfltUkVp5dvdGYx9mPHfFkhNnJ0oF8f86vjTr4acibu4kDuGOu+vx2c48sCj/srg
MXJOYeewS/LJHxwZ5zPpL81xL7cLkq7sJcPzKu5NYweKGJQ+11c1+n0XpKy4cB/G
aNffgSqQtk+bPycIaMumpl5j49H3/WSSfrKJHpBxw+WDnT5q0woaNkLQYj+wSma+
G35YUPlKCp8pqzpV5LW9o+wlQ5RcpG53Nocgtwjr1TujvrtXoPpg3FH0+/Nx5bID
OojYdEWaiuENX1lGAUGq2FPAAtwRwAFaWI++cu988wgR8WhExVk+vz5pW95LHrMD
dyl4YFaiVH4h/PCreHW/rUVDbOxhRvWT8cJ0df2H3BnshtyOEGdt+KDc9gwcewak
hor4Yuy5HXNz0n777SkOuOa+gsiUNkUoFxeEVyvkNHodc9a9MHxYM817XauyftGH
j3Vd+xC7069IfOg1DsirHhkWww9KTolHsrWca3XWEN8Gs8wgoM7y2ZNDPIBSzuUo
mv5ftnr5soQBXzzDWa0Us+oRpcMWhJXLfXwgexliUFytjdU2x56bMZd+Jq0qTr7Y
2kSyMktjsgRcE6B3TyK3s2APJMEGizSQye07tj4vlH5XHmXLjk/zdO9yVS+J8oU3
lD/igRHwywLtaK32+fq9vzcSi3ocIYhNgtobuRx0NDdIwUT+7w9ko79KvVPZBvxT
sBz7/zo6kerHlJxmNNZk+VDNGFnf3Lle6pkNOwx0zrx2EjmNFpMkXkGrySLuilnE
GckvgsedrTzSUFNRuHRCGruu2w5k1N9YkOoyn1s/JWX0fUG/B/hVPJimPG0B2a1v
Qcz1yf+MOXT6LLTa2ei+1cGH+D9TRzeMU6kmqQolxh5+RI5mr280qkGJdMJ9ipWt
FiMyYdAJIlXYYQ4UwPNmUsXmNTD/FkOXbdGQ3GeC1ZnveDzmM+DADk2aNG33wdH/
8PqA+vFJOze2kZtNlf20jzaMW+OX5nkgKX5B0GZ/gMj0KseWz/UeNXrX6yjpkG+Y
BxVnmP9VMwjKpoygR3StfOocx0JqsPZpLhPJFpmf9xwQp4zFuBLTJNw6wdDdVM0J
HDCcyVCybD2fivxaEQVDo1QroW7Zk53XsMvqQvWmjx4gYSpyXBUl06ip7Hu4kwHq
E9Fcmd05nkc8TCmkjNu7Ifh5r+QSPsczOzI3+nLjL1HzcPSoF/HQu94z6pbS0tGf
RZNzUwHOVkfQpAbsXkpLvhOnCi07i3w8kX3ZJjHdLa1OtVGqXi6IYDfTfr/zppk6
2EgYFVOU8Ia+8QnDoLrKY9kwcmSvfBjgw2sacLfD8sDSi3LxDKvJ8E4cbXmHrlSL
/mqf8Ts9TxrPnVQhY0dGVvClXbH+oW1vG50jaGEGWN2183zSo10AsKfhUUP29ayO
rp4LqPnngexrVgSY8J1WUAsOxLmtiDqarolOHXLHXTK1CpyJPXEFL4ezPn/tkvNG
zCDWRkTRMXLGkbzQlxB3HysGkZbKcbv1uugUpx4Anh27bHC/MqD2xqeUh24W47o3
KBa0CYBaSgzDiuzDhwvKtNW7fnKXAh2OW2MuHY4Pvted2Ow91ANOmQhSg+2FqFpd
KMj3+xOaIiOw/PPpj0oJv/se9NPvOFY+8EhJNwuMz0ugsACvBbNTYtxFkLK+8ljS
H4N3BPS0sdTDvqqztVjuUuvhAeawe8JN2X4g5cyOVhh6+y5QlZFbozobMQqswqbO
kfnKxfiyoPBTRW98gRyik4VlDAHGLJj+s6VitvlgnaVCejD+UHPLqjR60F3HH8gc
+R1xoZ/51neINYtdzVGzWyeuPUmzUfbMD9TAsBUzwssebZL5Nx1RSQhtJiUJVRuY
McfJD4gW/p0xb30ERFuaFRYNzFEkrMIJ43YhniSm33D2xesBvxq+o3Hr7HjWbs41
+U1h3I2CWd1iwF9kz+AnmmK3822gEOv1RqjJ0vx6Ut5qqlONt9w2KM9Io0ltirMV
8dRrlXYxhGuabmHv3dXXLmiteQqijszer3WVs5ls2EwtXd+gYK2pHyF7zh2Q2ULM
1WBe+qjkx/NJyS6mFHOVCLZJF91tySVOrzH0qAM/Rhx/LNMvV/k/UuDODYSCf1Wu
k5Hnv0DkjOihdclTjFN9z+zCfKcQO+E64QbsucPkuP8kAOYEDFtZi06FuMlhLPOJ
wywQU69kYgwWwKod5MqU1KwlzyEWejPylPWB7u3PY3/khyvgP00OZmRzTbLJcc1X
h98UdYi7vYpmRt+6yUaSRw==
//pragma protect end_data_block
//pragma protect digest_block
39a69P7J/fgfejNJ965J1KRC0og=
//pragma protect end_digest_block
//pragma protect end_protected
`endif

