
`ifndef GUARD_SVT_AHB_SLAVE_AGENT_SV
  `define GUARD_SVT_AHB_SLAVE_AGENT_SV

// =============================================================================
/** The svt_ahb_slave_agent encapsulates sequencer, driver, and slave monitor.
 * The svt_ahb_slave_agent can be configured to operate in active mode and
 * passive mode. The user can provide AHB sequences to the sequencer. The
 * svt_ahb_slave_agent is configured using slave configuration
 * #svt_ahb_slave_configuration. The slave configuration should be provided to
 * the svt_ahb_slave_agent in the build phase of the test. In the slave agent,
 * the slave monitor samples the AHB port signals. When a new transaction is
 * detected, slave monitor provides a response request transaction to the slave
 * sequencer. The slave response sequence within the sequencer programs the
 * appropriate slave response. The updated response transaction is then
 * provided by the slave sequencer to the slave driver. The slave driver in
 * turn drives the response on the AHB bus.  The driver and slave monitor
 * components within svt_ahb_slave_agent call callback methods at various
 * phases of execution of the AHB transaction. After the AHB transaction on the
 * bus is complete, the completed sequence item is provided to the analysis
 * port of slave monitor in both active and passive mode, which can be used by
 * the testbench.
 */
class svt_ahb_slave_agent extends svt_agent;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual svt_ahb_slave_if svt_ahb_slave_vif;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AHB svt_ahb_slave virtual interface */
  svt_ahb_slave_vif vif;

  /** AHB Slave Driver */
  svt_ahb_slave driver;

  /** AHB Slave Monitor */
  svt_ahb_slave_monitor monitor; 

  /** AHB svt_ahb_slave Sequencer */
  svt_ahb_slave_sequencer sequencer;

  /** A reference to the slave memory set if the svt_ahb_slave_memory_sequence sequence is used */ 
  svt_mem ahb_slave_mem;

`ifdef SVT_UVM_TECHNOLOGY
 /** AMBA-PV blocking AHB response transaction socket interface */
  uvm_tlm_b_initiator_socket#(uvm_tlm_generic_payload) resp_socket;
`endif

  /** AXI External Slave Index */ 
  int ahb_external_port_id = -1;

  /** AXI External Slave Agent Configuration */ 
  svt_ahb_slave_configuration ahb_external_port_cfg; 

  /** Callback which implements transaction reporting and tracing */
  svt_ahb_slave_monitor_transaction_report_callback xact_report_cb;

  /** Reference to the system wide sequence item report. */
  svt_sequence_item_report sys_seq_item_report;

/** @cond PRIVATE */
  /** AHB slave transaction coverage callback handle*/
  svt_ahb_slave_monitor_def_cov_callback svt_ahb_slave_trans_cov_cb;
  
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_slave_configuration cfg_snapshot;

  /** AHB Slave Monitor Callback Instance for System Checker */
  svt_ahb_slave_monitor_system_checker_callback system_checker_cb;
  
  /** AHB master Signal coverage callbacks */
  svt_ahb_slave_monitor_def_toggle_cov_callback#(virtual svt_ahb_slave_if.svt_ahb_monitor_modport) svt_ahb_slave_toggle_cov_cb;
  svt_ahb_slave_monitor_def_state_cov_callback#(virtual svt_ahb_slave_if.svt_ahb_monitor_modport)  svt_ahb_slave_state_cov_cb;

  /** Callback which implements XML generation for ahb slave for Protocol Analyzer */
  svt_ahb_slave_monitor_pa_writer_callback slave_xml_writer_cb;
  
  /** Writer used in callbacks to generate XML/FSDB output for pa */
  protected svt_xml_writer xml_writer = null;

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Configuration object for this transactor. */
  local svt_ahb_slave_configuration cfg; 

  /** Address mapper for this slave component */
  local svt_ahb_mem_address_mapper mem_addr_mapper;
/** @endcond */

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `svt_xvm_component_utils_begin(svt_ahb_slave_agent)
  `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE);
  `svt_xvm_component_utils_end

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new agent instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the #driver and #sequencer components if configured as an
   * active component.
   * Costructs the #monitor component if configured as active or passive component.
   */
  `ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
  `elsif SVT_OVM_TECHNOLOGY
  extern function void build();
  `endif

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   * Connects the #driver and #sequencer TLM ports if configured as a UVM_ACTIVE
   * component.
   */
  `ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
  `elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
  `endif

  // ---------------------------------------------------------------------------
  /**
   * Run phase used here to set is_active parameter (ACTIVE or PASSIVE) for slave_if  
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Extract Phase
   * Close out the XML file if it is enabled
   */
  `ifdef SVT_UVM_TECHNOLOGY
  extern function void extract_phase(uvm_phase phase);
  `elsif SVT_OVM_TECHNOLOGY
  extern function void extract();
  `endif

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the agent configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);
  /** @endcond */

  /** Puts the write transaction data to memory, if response type is OKAY */
  extern virtual task put_write_transaction_data_to_mem(svt_ahb_slave_transaction xact);

  /** Gets the read transactions data from memory.*/
  extern virtual task get_read_data_from_mem_to_transaction(svt_ahb_slave_transaction xact);

  /** 
   * Retruns the report on performance metrics as a string
   * @return A string with the performance report
   */
  extern function string get_performance_report();

/** @cond PRIVATE */
  /**
   * Obtain the address mapper for this slave
   */
  extern function svt_ahb_mem_address_mapper get_mem_address_mapper();
/** @endcond */

  extern function svt_mem_backdoor_base get_mem_backdoor();
 
 /** 
   * Gets the name of this agent
   */
  extern function string get_requester_name();
 
  /**
   * Set the external port id and port configuration
   */
  extern function set_external_agents_props(input int port_idx= -1, input svt_ahb_slave_configuration port_cfg);

  //----------------------------------------------------------------------------
  /**
   * Function to get the configuration that should be stored for this component
   * when debug_opts have been enabled.
   *
   * @param cfg The configuration that has been supplied to reconfigure.
   * @return The configuration that is to be stored.
   */
  extern virtual function svt_configuration get_debug_opts_cfg(svt_configuration cfg);

endclass

  `protected
E:_U(^fP8ESa5=YT/)_Y6S[L-A/1L_+Q=\aDP.J1#NY4)0VgYPQ34)]dTe][2VHM
<0PVK<D._1P]Lb)Y@G5NR99#7EAP-#8_0LdL5=7e3bL1UD,DW\4@D\>5_6WMU(7;
bcUH\G&c/[/?VM;9,3D+P+F(f6CSFK7Q6RL/NC-0c?F:^3+9_E:&4?2:WUSA@8Y,
-90(RHMO)]C#6&KP/6Eb]_bM&VW]4+):KFH:_M>B#@Id+8V,^&^.&TcL#Q)9:YPF
(5NLWC7;F;?755ED8QEG?5H>NM3<O1)=I(5dGXS748#dB$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
.1eV?V7#>Q:OMEQ14N7TP=SM\Q,.3]=beX9X,Kg8<0PTTF:AK0Ud/(1gG9U6[d+a
A@/;\f_@.3^[WF>:<.KQP]D20;N.=S.OC:P)Gc&GcBK]-G;L57dVII+?0QS8AgJJ
f[YX/_MC,,YC@<TY0J@XEVE=D[0Q>U)OU];-@^f8BM@(fKP_>H==-7?#=3TY4C>6
)PQJ_5/Y12UcSbRH(_3_+QcK/./.gALb2VH;:e_,OKBVQDUWP&?Z@aM2FIF9)gfA
6;S5.T:21N4VG8R[<M-^^1Qe12CR2A^;IC<MHDP@/FQ:52(UDCaUX(b/O;dbUIdd
@SYT<=J53H5_F9D+;7:F\+J[NRM;.)TT97?BRgXA38S6@3?Eb[]V_da16,&)DQ;5
dB.TE[^gg_)RC)[MSJK>1OGc\_ZbY,Qd]+8&ce)-\P@H;DK8:?BIf5QFeK^I9+E2
Q\b_HY.XFKcWgA5c:B+YX,QF8EXf=^FfVR#)M61^V0,N)^3@3_?bDSbUd.2Q9BA?
2RQXI:[6<#NI[dR0T:(51aU\BKIA[KBOGR3E20/2#Z\(X?/cfD5&6.Z/3(FD?f?G
&#IKJM#4I[OMfQD>X;1eb#0,?LCLL_^#g71.1G0aQMSd<Gd[<NQB4F3/?-WMb#Mb
T[(JK?EefLe(d[AGOefVM0X[4/L;^P.&39E.,).&)3?KeT.+ASb3VSLf93Tf>:;c
,XM7JcLWP@.K\&?EY0H2HU-\2P\+bG#F#eOfef,^gYG2PI-/EN0_0,O,Z_?R+fd0
34JGWEY,KUMfc:V;G)/8NQX<LKY)>5+-Q5+XBKQ_17aNaT8cg;W7AD&U5)ZSB682
YKQE)OZV[KF&E=8:9B[,BU0ZKd[daI:ES.B.c4DQd1)-&C,E<O><+>/;W,21HMcW
,/Y(QM,?FYVXV=]MZ?8JW<@DU:@420=fHBM5e8,V6OQd][SOa1#WFM;ZE?153PVI
5LT363D=<DQ)bC8Kg5>N=0->NK_)Y?/cb@OD_@LUFZd/RGUQ1\H)F0L2I@ISbT/P
EA&)WMT.B)9deD(J2WJE>>8DGcF835Y><71G<X#_)d8^[-bVf:8S6QEZ:LfZg/0-
UE6fff8-_WSVSE?]N\fYUZ/1H0HDgP+?PATa7?G8-A@,UaBMRTE,\_DNfeE3JXWX
b;G3^,VE7_C7HXU@N]]MP\T,L)4@JGZYbKW?LCKG@>2;1cJQB>)4T&&[&5GS@bXK
1MXfaYUde3<VaP&1M=LCW5?0T019]b2(19PD9#Ag:OM<6X[99Of5VQ8?eY,0VXKV
BW7JB_FHFQ4D#0:@.GRT5Q)@bLDcWR(7F;#F7P,#^aa+3TcTDBY#EWDTMcVICC1.
D73gT<)3+V\U6GeZ56Z=:A4?L//HOc6+H.Xc9V4fAKV2QX^:-H4Kf:fJ.=MK_d/?
+FI1]/X-X02gNB2e@_9AGMXZe+/X0>?J/1(HF_,(L0U&UZ,LWFE>+W2^R9a0cTV^
ZJH^?)#aJe?b\dbN>IAW9I<@B><dgb/M59_3>b>5##\BWU&7YRB@b?+\:0SaZ?>]
BfM8_44dad&K09cggMP@#2_1\UC9JPXNB8/)@g9S+G>,D0a047Yg02RTR+7b+IB6
8IJa26YSa8_Rb#4f8ZAONQeO^^VT.E>M)IW]W\T1DPb0_K/Ng?/WY-Ub7Mf>.D>=
T(R2+/F1-?:21HRWe_fd_/2V2/)P@_LR/XV>6]FIP_c(E1^8/1<+J3A^;4(Q-&3[
ROHD2W:Z5=FS3R:N[[]_QMG93gY2SG#fG\JO=G6<[A(]e;#Y,f25B<U,Y,MEIZ1W
/HW2BVW\3]^2256)39<[6[;84TbTIe#YF)&B/V?9]W<\7T8-C)QUJIG6Y<7?VgdI
/2A1d,b::.g7?+-LS@&/:PFc_QcWF?X2WUKS2-:+<(/O1&_249]5^E7EF\L>BMDY
:6Yc:B/)EaAL)[@5KCYKKNU<OH@eT?&.d9S]]K&N.\AN4?(3)T>K[H_CV4cY#?1>
(C8^K,1e=3c8\.\^\=ZREL+LFP:7:GM^@.+VTUEKb\1\Y/^4KP)1[6X8Z/gO1HDK
,RT:RdQ-0b<(2TONI]-FQbAH#)_EW^[;SBVfGOPQJ5(/(Wf>1?LH2JS4+0?,T5Mg
+I_JYC2ff/a?Ic.:]N9Z#6&X2+Kg3AH_f2bP]2JCK78W3U[be2>+FR91AQc4:V\/
D:0dRGB1.ZR5662CHW4_dK=S8VLOT\M,6bI7Y@U.ROC[:,G)7].+?R(K\MJFZLSR
eA[D4/2EeWRDU[f->@_\^J1->XV(YH8-/Ta;f)=FE1]G,6DJ/Z8EC5)gI-YS&/c1
VDg2:&U[C&ZM:HSD/+>,EKX5d1SJ3UV.^fbMQ,E89R&H;Y5WR^Y5aT/,SP6Q0>g3
(R.-Z>RJ0,gdPFN.U#K?Q6^)LDTJEd62O11NfXF@2IJ]OJA?;&L6)[<]gVHQ6ZeW
QfA88(/A>9Y036FPDEI==(8UK]@EMY.DVC&^H/X2)U)fe,8C^.2&)=B^ZD92<PU-
#4]FG[C5BYGLZ^Cb)#=5U\-@cJe2U#8+H^@5,B)0[Vf;IKfE]G1F:;A<<d9/[D3g
+AJ=2+FE38fV9#c&b^a&QcD8ZDPA1EgO/cPc,;MF]E\P3GBWLQB2A<_^;.O-)<&P
&,.-f6<Q+LdG+T27+c0<2W6J7gD5+E0Y<bfQ?&O:A?L)cCMY/41EV_:eUTNG)LD<
07#9ZFQV8,F@4]R>G34YbdLY6e7KIbaO82V_&MGTR=,C/Y)(c#9]4Ac4Q]TS<YOL
U=HdXAbd,OU0;T;AUAHNO0);G3T@>\+J;_)V3@(4)QPPNARY>&6E-Lc(^6L.ZEI2
),/=?1GM[SV(e,eXOQH#VG7>H0N-=;PF[gVQE-DIK>T;U\_QQ1U)SQM.>e#@2[GC
FGeFXW2FaG/(B8<CE9D.a3P:H._&(H+]@(PO)3@.Q;RBX\\[<7_dA7S=ge\YF)J1
DXX^VTK.NZY4\:cTe6K-ePNK5[&SF\/+&,\X[e32HfF]@STU8OJa:/+Y=80gGO_E
PW;RD-2?3\.YgD-99\fgb)W@5_e\NX#G70;,GcHWTBUB[]SfX\33PbZH+[dKWIE(
[9;MOgBACK#UA&T&K5gc-R)5N1;L^J-3.FI^?&BX5>8c]O,ef=C??AQRM-e4G.Q#
V4AB?H+)Vc?bN#L\a\dUfR/d_&M1]S93Z5ZUX5fP4T?0fLMZ=g\2D>?g.MR+J-B<
TF;::H@ee1H-:&.>#<S^gA@BPYGSKG1F[S+9f=f_(R>Y2/fSFNM:[<1A&Q6E90G\
_R>=U>E]dc=:@0]7;Y]X:+XJ6CX+ff39,D,8c0N&/H\dUNH)6O8P37>DMf:]Q_LR
c?SF94<=d,@IALGNS+D5((9?,R=C2.H^JL,=@e.DX1N5@OAO;)AR\M1_Bb(0_De5
cU,-K;Z-Q73GTCD&L0(;a0g;SXgbK&5DIL0(Fag?Vf.S,_gG6\?b9P(;I-V#2HB.
,@dc0JB8=L(^1^78KRYRaGC]@V@bSA=e8UH(Ja_9]5&,3#K_Le1&IEa^6(?8<IAL
SH@bX([K[8cA1a9=Ze,NU[HL3c]+4YfU>S&T8fg5V46?^X<P38FH92J,94SC]YYK
Nd[(72=KD0LeY[9VC3I8AGR++M(d;/2)XJ/LH2V.?<Iga)DAgE5,=O[.34@X8e_,
F7e:8DE]O_.0=(MAed:_F0LW-HG7B2F_>dK]DICWT5Me4/e9g&L.>_L>fYL(PQFN
g\gdf/Udc/)G8FW)/gg^2g)T1><ZO4F4=.<c64=+/+0cA]0ZQ1d-4(B;-,c:+F_M
\C#)7I^;LU7bF.7KM9OXZ[g/->EOGH9[1-Q+(b4BRLLc7cYO_AZI0(T0a#<82CU+
aS#+ER1^\1>YV.#/2gg38da1,B,aUIc1.[VTH-b2]b<B902L=9_\=V\YJ4B09MX,
A[#gGg0TK[2H?CfbNc+Y<Fg-H:^4;Bc(=:/A[?Sf1>().2D.=&L)4b<^RG@^X78;
]f2^3I8:cc_a?d&XgDN_,c)L@<KgaX5SGN8TYM:-HEJcYMV7]a69?2K(OI)4EKd:
)b4&X=<e/fRY-.OZB_;#J[J-?OQTd1aGUNW))-Z&UI0b7>I<7:OO5YF,A+E+3K<Y
L?0gH)Xa[WUJN80E<>&^HH]B;d&0+eAe/4#.I>2571cYF)O6F_@MCP2LH]HL4Q24
7Ecf7TVYWgT7P1Y&XdZEdGGZCF(gK&f&aLTHXJRU?;J<T.S/>6BNJ/f=V/?(&__,
GM,QU5FcAQ3V@g;<,cW^-c5)/7?26We;[Q>C#fd-b=YDF[3K;/8H5OJ?5COc+=(-
ZXO&P6^I=H\-gH_<=82GUcUEX8c+?A^]LE90aV#C,P>(?L#J\7C1D#bZ?d8d;(<f
GRV4-bDP>3bI[Tf>UM.9\M8[OH[XCOJ)PL(bPd2e38P-b:#.\CMKC_Ce(X4X=55.
,g5K_d4SIG4]IEPZ62GW<WK2fETFD>5BX7A?T5DR7O<VUO->W2N0fIJS-_gGDW)V
d6:XK[>dSVSV(UO9D76YPfUM>=BKVPXXJ)3[@1@BLg8P-3><[CaM4KV:]F,4Adc3
)(W+^S&B62#f[4G(T_]4Y]C)97Gca.ID8,_g;Da#:/YAA_LTH^/A_f/#E&XI0G9/
04I];[@Wg8CDE0=N#e<f3PI9)HWT[/J[:];Y_QI(gNOUf_eN[KO-4/^Bd6LY6_&2
L+7Q8YdWc_;1#.XR/5Kd-Yc;+96;XI2)gMgRI][51RV:?U+b:f>(RHJfEKNVV7X;
T0ee7)F,(QKFAfO]3560O(HS?cM94<0TCP^f??5/<_/@&]PP_FZBJD4[KbfOJ+W@
PJe?UFbRN3]7BgXb5/#<R2H7c^\48:SNe06\-3SL;aW<@\QV:2UTWJT4TRFZ5W8B
gGc=c;UGYS.>,^O#6(Lc/H;5<F+O_3,U<.1f1KZ>:>=1,A^JG2eE.RL3M)GLb-^V
\<0M-0?dW8+@(gaA&I54LL?I7B8T4RbD0JENTAZ2^4B0^d:R,BE7<QdE,^,b7beg
TW]cDQ,8-<C4@@IRL7=Cf2aUYb#C1Y_abD>EA9a9Q7aNS-^gb.8#W:@6BTcUEcUW
b;]0;.:DaZ4WKWVO^;ZbN4J#CE35c]U@GHGe_R(H.aS;b5YM00PSNA2HG3YJ>(6a
A02J2YP9&L&F=P9JE&V6fU4agZ<X.UfRLFE//I6XL^W7O>/5_GZGUKDRV:RYXUg^
C0&a(][cgTB,P&)N4e.#@Kg3JL0A<S^e]3KTC^)f;PTGZV0ETZ/8JD)CD(B05=SF
[b7&4BS@9QF7NJL,3U^H=M7>B>;UK\Pb5342f.;e#SM&XTE+A5;Sg(gS^6Q#WTQJ
KR7KDZ=5]2&[G,d2[<DQ<GBSOM.gK)NfLTT-Yb^:LA:>??PR7BJ^Jea:5&N<#V&^
&T8N9N8NPWSc,F:VAM5QQdT@U<Ba6<N0NAHY.bcV&2>A)&&M;aL21U6,>V:FQXdF
P^LbOKQTH3aKJFf9PR5X/O713OB7C/<CGU<O/_]PY^_>YI5[e+[+8Ye?Q?N4W(F2
N/a/d0OUfeBT\ORCN3]Qc&WeZZR+^2QZPWSO<GcOP^9A^708E(>aLQ8^@N44-S\F
NAe:A&]#+);O]N=IQgF]bHLS)SV\_f+23;_c0+?TJE.d132J=PYA1?=]3YH8NYX+
@+;VU_QgVGH^LV(F))d=,]#3bdeUg4,-c[]8JdM[5Y5X]:GAC[#R@EbNfN_(,?eJ
>cAdS(JC:O/Y@JceS3R>J^24Y\O_\DM2feP&5bQ5bGRW/36a?\N[;:2B3H-,J69\
<:2QF(QcNLIDc69T,EL.U-7PE\+H1M2M)/66UN6=QF8-MA1#QU:>RHG5a93RY28[
Z.6Vc@_6cRO1&I),8ODBc#11#5gg3IHJCS,[;eZc)\RY8c0#eQ8IW<O:QFESP#7P
U?B#aQM=W2I?U;8>;.ZB:9f:&C]IG4#Jb_+/LeJ76aUER7<8,\N?@SFJH5fP\LH\
H](1K8-A/+_6&7]0/g2Z-KGW/H1ZfK5Z:B9Y&_ZI05:+QZf26gBa>36g?L=PKe3X
?-GJGWC6@JOR?F&dY-JH=\;B9V:^eQ40=<fFQ@\Y_-[db)]@SY9.@^^B\_[D_\4D
eS^]=B-6GNY:a.JK&_,6Lde.YbLID)F)PNZ\6FW0(F87-)d8Q7_UHG]P]CSE?e-I
YcG>QI#-d<^:.O)K@:__XFdV1E\49@YY#3,#9UYELa^cH@HS@2#&T7L65BVH<X.,
^UcD\)TSSMfF,3d([KC5.FQcP;/b15=+SLc<g45DG^_WA]9.V<U710VS7Uca0^ZO
1e12fAg]5@R6-;I/-]?8[#,S9L6]1a#M#-)_?I&(J^fBT)E+3.&86<W8a6Y0Uf+T
E@+.,eDX)gVL)RH1FAfP24=@3D?2[g)]V1]U?L4b(/Zbc7:G?U023&,[e1eG26T(
Rf#2>^Q?5Y4@BBIX5+DI2GXBU,bOW5N9>5B0FfGIbTC7=4L(W6#26@+O7H=gFdd/
:fB5<2&d.)TQ>-<LP,T7HbU>F:W<R+?RQY7fF4QbQDU9J)_+VP6+;N3[RPe)Gc=I
6KeaeH3@e=L0Xc,(64HG9G6_NP^+GG;4(,HcLD]:g[UXBHX-@aFBTLC41/=c>P;J
VU?\VB9<H-/PbYPKJI<]4>,gWC+7&0.GD1cdGNQ4)6-WY<4M&NLD/T(N[93bM<cJ
78d39U1e_8-7M?1P-\TOE=C2E^_]fWgNT5;e9^92A-&BgA::ecaTfF4Pc,?@DA,[
caRbV0B#,XdYENc:1)gbFQaPVK&:5Le#[SJ/VLNO4HD)6FUID4_;eR?gXA<ABAd4
#H:HST?GdcB5VIf[ADE\&W(bU4EbD2N=+6CA]:N]d5E<RKP0X:)c<OWN?;3)(9=H
;c,5eF.f[RE-JHa?]Y#(G&&;H^4SPCQGR=b\QYSMb)D3T6@TE:6ROEQB_a(?_g-K
+3W;BV6U]&U<YH,+=C)FYBWHNT=Hc=TSU0efc/2NFa[;[SRa<1DL,7(7OI+IB.Gb
Y2;6]J;:T)F?2:W@5eCBG#OHf1N+HANDC6AXD.NH,2H_Ea_K(4ePQAY(Pe1-UX1I
bR.+F1,RW@TMPZ70OZ-W?e(5@#L^2LgceB9c(T=^Yf\AfOWVT-T.RK8OEIPLO[a(
:#04fRMEIX7)I@fSA7V;:(@G]bZ,K8KafJNC=?Q4Pf30)Z<OF1E.#=3XYAe,74eC
cM/9a;R,A=L>cPU)W/cO/2JeP_@FKBEV(M,?56.0FRN7dSe,b/1fM>P\H+]U<+H6
<MJ8:XGO(#PN6N5)3VeSB)U>/7:CfA6O;3JC@D^SaHH>AR=8U@e?0O7PBGP7Td-R
7):+#-Ob&B?D>+1LMFZe40\OH1&WVZF^]W&N/3eFceVD_XD.EZDZ(.JLL7KP^81Q
KWHf\P_^^(8BA==W=AQ<8#(())TL6C&5(b;+OeUIFLWb[-4Q;,bRb-V1W4LOV[VF
5S)RTO7;=41ES&bR\cb2,-IG0_Jf[\D8#+0Ce1RE8agN2CVgfgL.9cYFFV=,c=A\
+;cHP=.,IT[9EBA?K8GcEb?<3E+QWdbRE(f@R?(HAER@6(W,?6ePAf\43UF=/c>)
S47@>+(g#1-NN=>33SXTM7H)2aL8R)>#LB&M\g<@(SWD?5-0<6BN(._VQf,EY4SX
Y#1(bF<CC)A]?>aT-Ta^RUGAK2;dfBY[g)]BB6.0Kg9W?P(R&4KD,_gH6O-MZH:4
@THKbJ^0.2U++K_U>7W@WPAIRRNCO,(UCR.g+UD_XNI;_?AY[_NBF;D:NW(OaG=.
MR84.^_e6&[K4>=g)Q&[(M4aAQPEC>,[#-R4_VB84,8XHDf.JVg7US45A61ZWY-D
\6B=&AggBAOEP.F@&0\eONf7VAEBZ<a)0&^?e-.PX.Tc].\7RSf1^(TZPaD<3-(N
JcJ3@eK;c9T<cWZW(C)I44K\VC)3>bL[);WZYZAI)&DDgF=#Na1\>&BE3K<B3WNg
M;H<fa5H):=DG:bd&J)K:Y>RN(,(1.:\FbS7DB1T-.)BgTf=3(C#BX#&XcfML48g
\7,V8/HYJ&geRa2O:2>ESDV?,1EVGb4GBG98G?QC\5F0)PDC&KKC,AVTcK](,J_E
Og#<<K30<)GU)R\4.E\WB0C=7Q.[+2OcA(HJLFgT5=V6HAJ0M4V](C#OT9F7.J[Z
/NF,\Kg==.AaO949(G@eaed4b@JMJD.a&Pa>&^D/NSE.7L_(U6@d9OcQf]#UNc^C
gdG7T0)1EgBcCDG5T?T2/C;SP:WbW;[gG4O[X1f/69JKT@IbF)OSU+;V71OC.]Y5
UFeJAW9eXcd3CIZ<Z]>#F^3UCT])F1K9^^.f[N?YRP:6O:/18<0D?VdfF/B]c-FR
B4OI=-;9g)29/@+EODR0ZZNP^=;:IcbIg6_HL64,:&FQ[H0E@3M?]d1Z&^7V82)&
8GFKEKcXXagSQG6dWVIJJK0;L9gU^\?fWQC9=V08V[6N/O\9>WJ-6QK2(dFNM6=a
IU+U\SHQJf0f8Q#4ZS\YdX^YYgN=Y&g,Ne7PEUQ>@AeAe8<DB_HT4?+V@03HC+C+
SVPHNbM39N#b=\54,^Z0OUDbUJ,6f@.>KcK7[)DBVJd<@_6Y+UN]+K5307)Ef\c(
@VOQ(3c^Ug\]H).TW2NY;9AMI1dIPA)HHRAcG5K#U9J4)BAT2OG9O2Q&#0Q8g,.9
LGUQ\LOW3a+^.2Eg5T0f(2PJ[]Q-Va,=LX/G/-=I9W.&__6/bOWLZTM9IT692LMA
+B9ge1XK/VXDWc8+5:DK.B]KLPA0^3\32F6VA.[1RO[(/TI;dVVWgO>Bd2;9O+0b
9;JP&J;cBU\5.I5YBaS>XG(=^E\,@c/=,OWD.c@b3)c4LG=9S-#1MK;KS[2.2RT9
VW_&+XFX75/HCN&fG)=>N+aaJXK]VT/@@(0J/?b:-d43HW63?D&d\T^L/cb&C]=9
SGeL(d+aad/DJP]^@>O.44X,H_I+Zf=ceMDb1S@L(O2LTUeB:.J/C6<7[^aeLK,?
8,^4JXDfXeY1=b=a@[/-2]C&75RCX\.3EEQMN4\<8Cc9=Ze3+=\(RGXJD)<_7c>4
8F=SZ(;;Q7&P<,[YSQ13JKaa6>U?NK#E;a)??PMQX[:Jgg9=RM>2FGSQ0#T^TGEK
7E.fKfGIDPF-g+g.ZeP8(ca55bb,W73]Zf^NAZ:ZZdd]0JcI@5^_,\7PbXY.-:1I
M]/]e:QIVdLUMNL-c-dD.N0U@(W&g4fT>CV=[/8QW1(\&-aU-7Tge&eZ(<6-5<fL
6Y0FZ=2gHdA[,Dg4JC^d6b;^FGYZ,FOO+(7=7C@AAB#5EaLQ2c?Ncd/H-6YCg2@.
?fZ-[8>^J^ZJ47XRVN6/:GaI^U(SK</DbKdfb:UYJV_MVZ2,?#MP:/I+RY[@,ScS
/25[cLD5=;(WPeJ3F\f#eX1P-9@63a;Vd>V)H/3FU\c5De0,eH,=1.DI)1:->SI5
=A@g>-9DFX&&H3-TY3?J3<.FN4[;E1OB+=+5TR49PdE.f=<fTI=dW#1=X93^(W/1
3a>EY6+b\E,Oe,=0JbP-P/R.M/0M0e8?CEJKY>S&O^T+(Kd.,(7IU.<^HE]A3\P6
P><=:LMK[..2c@dK10c^<Hf7TDQB5#g?D:HeZ7:FUHCWZQ.&27ZV.aQgDLU9c-=Z
@>2/?Z+Q1WHAVS..BF<[9aJOC3(+5EW1TIGTd7-cI7Rg(HAS>H(8Ka=M]\DUE7/S
cHDX&MW@d_KAXLCF+S:DU0cSKCIY(_bVFf#WN@?,]gcCK/]BX(YMeY3:RD[0F]1a
F7HNI(Z?KY[&=9,:V,cA:?>P+W-#Yf;T/VfMge246^XA&MNXTU_/9X]:>9M)Y942
#bbSd?=B-Y-G20[H-;ebg+bD=KBU@QQ[W;Jg^TSMUb#6U#RVDPWH,8.GAc5gQ&cR
JG-g.]P0ZbHZ.bZfO5O+/&7b2&0BJba_9EF2MK9VJ+\#KBD-/NL<:6G26[f_D+fY
=E?1QP[_d5R06]=:&+d,=b:f+;TbT\]I@c)#>-g477Nb=<8@>)&1X#f9aPde__;?
]TbK/+Z.E6(G/1D,^6c9<-[Te;T(+N;15f8-WBP&.K/+HO[4d(=#g8fJ=@\0R8N:
PPHaTL>6cZ#dW_2ZWLUJ<)]g]Y.BBaPa]GY1,/&1.:\(@]V7cbJ;Z&3;)[g>;BJf
=]e>M&7Z64BKBg/Z,L(G3>OZPgNC9>P=T6VON^X#6B,D];X9HGRU(PY]ad-AA3;O
Y\=;UeE_PDM]J/<:W8W;4B;a\Pf/X?(Bg149:W^eS5#4B8@3b-+T/U_/cJE6faf>
F5;M=L045#eP53e^gLcW2A0YdQ2BD#3]IaIN97A5CWW#G#6f8\A>7fMRCagT_TDW
bI;97I_&d9,/ZADHFC_C0]3#g<D@F6,\W>g3NDZ>d1[eeJ)?-J?)5EIQadRW[NOB
9><RA7UQda?YE^;Z_:#HT?.U/g#9dI^:H=E)^4>McVE;G4UB@]g1;S5/L<7d1U^:
gZ;5R./.ILPdQI9@PP=@U,6ED1d846c^L1O4:Y2CTCCJF/VQB[IU+Z>#&7<LOVa0
K5RT8HW4NR]Hd:LO-&H?.)IB/e\BNWLV[?2c^g,G_IH<K&bJO;c=2E(cVHAISgU&
^&KY<5?VOCE==R+/O>@0(RTG893&Qeg>GOE3dU3H=GAR-?g-U6ZWgXe^J[,W3NB>
JdgXJNI5ZUQ>Z\SQOMb,N14Q\]a1]YJCfS7=Rg)#)Z=Z.[ZETCe@FV96RN)0bLd<
ce=A5/a(D4Bb:(d4+CI<@8/TFKO[M@:2,W9/G>97)(e(U-Z4M@\KD1CV66c\T88&
2HJWJQ_?Z39?LJZ19:@P;]MCHN2FMY)^JE,VFGgZ,HHWH\&4.\BC&:[Q@1EIZ8bF
Z0e4Tf@3YBeM_^fU,ge^7U-_<7_8[65cB@RfHAM07e^)a4-O5=DV5>@.bTH2N>f6
5J7.,.#?;+#e:[<>MUB[8e<2:0LN<K(F8:DOUDUIQ;?8J4]=+.[?KE^K#gG;6c&A
)_9Z_4)0_4N]Xgfg[=<ZOc+D4a:T05&=(bCD)8;EVP?^W3]ZVe@7AD0^d4F/:^;\
M^^P^=1=E4K?C(Wf(0?9Y2+M<g>SN.@9Z6eD8+)Y#cYHC>&@>5G,#LObE)-7\aT(
3V(L^T4A[3G\@N2UU0([.78[^]VV?.c&d</b1Af4?DDZV\=9]-5RZFN&K-T0F5eM
2T7e]E_G3QV\JQd,G_SVYcd8E&P<&baGReOa4Q\]Oe3N,]aYDEV/Jc\LAYPPWV-4
b.;22LRQ>,dT^;#6NE&T5(B,8T\2EBe?=Z+X9/@d6b>BC+8#G/,fcI/-g?Yb4B2V
#2L2@[51>?0YR0@8Kb(A.Z9dU.E(]-;_f/+CKH8e&UH08ECbcA0W6N5SW60RC^5/
MT\D1+HX.S?f&.U@>:c,D<]96/7M(X4\JA)CbfUX:g:LSERaXLUB&c0:LA/(d2Q0
2=BPd5G_RS&6aB5R[\5UZMef7+07^c=R:TU,Y:TXLdX[(CBSQ=33#VEWNQNNFIe8
2KN7\]ISb2(H#9d7CMNAQ;;E7B7HbK:WBFGC4.F/T.V(2=4PbdM\#^RS1VBgEgPa
OHK3(Pf/6K#3L^L,MF4U?#]EBTYW;,3LRa?_cE^H^I/GeO>B.?^f7b6.P1IUQE#)
84\U[BOe_T@0Z?\K<Ye7KG=&]6YN+E#L4Kg+Z],<]?@8=7gPP)<QTPbYaRWa@a3a
fZffW52#<f]g(I9P,g=gONAC,;5b_GV.+A:/Vd\Q>DN1X)e+L8:QK5F9/)V@)UWf
/?K^YFMTHKVRZ?PCcDbZ#A:AbbP[QEP/DdPCfLLD\CX:1E1ZAf3a_4,4\M?+/gK>
S:cb1PY941?M0B_^9@,HZL^CEXA3.#?S>4:FBc=Pa+[2;^G(J&f2&&&/OVFe9_4U
(I-g8g)d9_^g5GBe1,?XYa:]L)?2P8,9\_]a.;8N\F#6HW31UEBTZ,bJdJb&F5P=
eJ&]eYH1[<c&<dVCd53OC=P[5-V=5=CL4H+<4;I@7(E?B-5+Q@4NDdZ7Bg6BOL4g
9KK+Q>88gI#KHaZBYg7R=RcC[>R:52A169[gIR_#/,15A4MG,/YK<Vc2IJIXJ[M_
=QFAgZfc<.:1-C.Hg(<cX^:&7P]NEE\UY;J.AW?L&9M^#+VZF5S^T:O#^;W<^=..
11?YUe=?T\\WM@W,aAXN&[V;TZX\9=)(CHEDE5U[AA/<,=56-Ua+0Z&3f^&42^S5
Qc<-UWXH>WDbOb0_SALXNG>C-2OI1^0b]O,c2Y6gX\-W5@P/YfR@FELeWIfL>TS3
.[UADBX][],[;fF#,^V:eXATU(5A8+EdH+HRH:E4\JF.(]LE+f668K8c+URK1\YF
c&I-;RVYDUQN?2W3WdU:^d89;)R]HQT4>HgIC@gUOQ[d+];U[@_/[71U6:(=PYF,
89AL\?4AfLQ=T-gZU9X<-0:H@AB_.]\H.H]\8Pe3I.8d46-#HY^a0&L&W+=Id4^P
>8JO[_5O:F9/KL1Me[9&&ET;SZ>TYQ2G?5OIZG6ff[9IXgDbKf_S;T(N.W,8P,81
]TDg8cE1<OURa49#LA.eS-SVf\2P@#R/3:0dWZ:cb;YeV.W^1=X089-E[,W2))FG
Q,;U+2(93VAf&R41Xabf3TOQ2R6fV?1DVPX)7THcNM/91S-fB44?.[4<[LL[+6=-
3GSE;?\UP7L7DR(K^:RJ^[=)ad9J6@,_+[>RGa2)Q(FIgWd#;U->EJ^^N<Y//T)D
?&O:/cUXZA2;)TGFJ>U@UGK+1YVND[fFH.aZY)^&=M32CaH;gJ4MOL@g&<UYXOL>
0aI,Y3R7Gg&dJdTY[f</53\<]3dOZMT_GD#J?3]ELO\_W36[=;c.KW[7#?.U(C9E
KTb?0E)E-=9A,Md(=a)H5+AeSH/18BdPI&BY8&TT^?DLadG[C2XV.9I&&^Y.43LQ
91I,_7OIeVJUD17,,g,>Q5Cf^OSCRRd6V0-1WHTE2<[V2<_2@M<HN20a<eFZK?+a
;06JN@DG,96gFa9_5^@-#AZ181&AE6XU<cJ>MeP/bH.01I:ZI-E^bIMQ9Y\Z;UR8
NW&-+D&H=7K-?3c8]-TH\FLVL=d9D3OT]SAC+G]S&K]#F8]URJOW\<L<_@YCH0.M
-1Hb\(>W@P1EB1@H5_^3R-QSL?W&8_a8(\LR=6ff8279W5UWWF@/e.+e]5e/D6&F
90B:<B]8-d0#bU&UAO.EMdVN33)fX5_3]5E<.6)>Y@WQde@L+ZU\&)8,QI\K@?dT
,>KKc:G?D\2:0a/(:eQ4H[MLO[AT>[WNB@,>b_VLeMPACE:e7G:9&a]GZ4LIKCWI
-8D]>[1LR-C@L=BdY=5)/KO1cCf=4;7HK?@aMS=a3A-W023WafN]^&GGE7Ra>?]0
=bR68.<4[3Y3UVEHGc:7UU/._.@gZg_K(P#e=97,.)?,XM/.)/0d\V_Z,_;S]<MJ
>/I2KC:1Sf)If.@b3&WYK\>b)+K3YT91?edeT5Y0JP[\BIFA+Ra&/Y/\WJWa;QP4
_+aY)Q]O:,^37gGgRFC,HE&(IG=3LC3+UR4PN9Ja\XE>>#K#\N==?eS)>J/DM74f
cAJF/#)15KFU)e&+G;^H1]]5I5>9N2,ULcLeCW+Y#K1+88Yf#Bc/<^c<+H?D;P8(
@I]\TGVZ&M:E7,e[R9&68UJ@,FMP,WD^1+W2b=fU5\L4RL?^ZU<-AHcV._Nd01XH
L_-R@0)SP@0OU=8G7gJ2FRS(HQ3N2A_I@?;J&VWOCAbS8#>]3WM7+Ig6S9Y:7RRO
NPb\T@VC;P059eHcbD^3BOQ/cKX+g2LE.9U58=_FWG?@,F3_2ULD9#(&5aPZ@fT7
R/H0@K,D/7C#7fQgQYKTD7JI/[:86-d/&Y.+gIFf)f,38MRH//9>/N]NFSBK?;],
&SL/fb2OgN/H12/^[1OP5&b&(^+M<YJ+8aQ>E?X&M]]\UY\QcL&KGX9]6CASWX9T
F)g&,4,.gY-K-XUb[VC-=-BUMG0T,Pb,,7=2B<UCW7(,\S=;H3\55T&Y7(..Q4E8
4-R/8bI0VFF_c@PXG]Y.VQQII&13FR68O9VD??^&O3Od5CUBecBZ?daK\QCQM#@E
(.QAE#SS;Z;GgSE7NK8(U8?R6/7T[5g-;RNWSg]6^E9:^59:95PKGP2&&FS+H_gO
K2N+S]SP@AGJKCd7,I^[AW<J>bb.]cOE,?Xe<\Df/&-c+7J05M&](fQ<cdJg,]8E
(/2EG@D.VAdG,<B:bX\QFZ6KfV8Y0cd8IW[7OHXU?A3G8YD6NKFf\e;P/90a6QV9
J?7]ZYTUTbHXb3NTN?IA2fa=S8XX.HN&;CVVb0;8-H2-6/c947XdX/?[ZF#ePP9D
TZDJ<D:AQIVW>M9HfFg+=7/C.K\J1)@^O@-?]=Xf^E7=3M;1RU2Ed]dJNKY3R@)X
44I3[AIf+e-c[>+:8(7Ze.db/TC;8^N3:P6J/K\d,BT3^Y0f@(.JcV([ea:I#6dG
=2adbH+@ggI+6XZ;)XE]MJ&@NL:Tf+D.f8J6#HMMKcV4dB2RP\5-B9VJBL9aYZ1S
9L00#Z(cX;gIaJ?4faCE)UF+Y#+AL)>K?g5.D)Be2-2\Y3&2b+QIE/?gAX@NZQTP
.)a+Qa1+QSO./U(M4_KUVRQT5TND[A:95Jg\aOeQO\(BOY=WM^D4S[/BK[RPQFII
YVL&]a\VaA]>JaH)\#U8QOaU7cNB]e+W\RKP7M(ZbFH<T&_LV0GADa1g4d#8TPN[
D0+3:1Gd=7Ia+2ag];HJ1&XFdf8Y\TU(]VAQ](VJgM&L)@7RQWd3L>UOIQ;YV]&I
;SHF-V/90EO.YPJd2B<AC?HBC.dfLSI3[Z7VW6@\VZT::_\K1[^#S@-67B;DIK#E
,-4e:H(G/QM5OD@CV=\2N?PaIF9Y5DD2O#D:PN[<]V1ON0cNT:aR,C\2\0K@X.2Z
TW17-AMOb;g+I0.TeR_NZG;QM7L5Nc;bg9E;cKGf[4d.9SCAQ6H:44f1(gR2cL&Y
K>Z]7CFYe5HVfV7YcaJQX]Q5T3S?(&Ha=CL.\C0fd9-^1QIW]8cQ],+bBLF,=e>6
U,cZB(0#6)BfbBF[G><C/K48=^W\4YS?F/,P.P)5Mc_[2FeG@;A+6X1>FCH04ZD8
K8LcHfMb6UE0J/?&(U/V4H\>bP[Yc#I:e,H9Qf.-4(<WXF0A,_M4GeBKC^W>ZF7C
Faab2OK53T54>=2,7.B9cK0O.Ue_ZYTe,M]Y9YJO1a>:2/KP1K]DN.C2XWDQYg,7
+7#ALM-RI99MRF\L1@Oe7RP8GaI\ge5.c;S8.&]gLP=N/e\^+JZ(f#06-=^)?CXI
;X)<MdI(dQG/6cP.R;c^0XNKEb.9@MUD(@SU<\H8ITcTP:<_E\^:Rc?Za0W8BgI9
,Rc7bB3+GBbf,P#O55Z#_BZLc2.ZdF&.&b:61^Sb--gbZZL?<@e_MGKEgJ;G;fV5
W9\db1ODLca4O_RF&Ba99B;WRg1KOCY(5^8g.NVE8a.];K-A,d542#KKFA.:]3g7
]8NUI4O/:Oe-&9;?J@QL,_]?F/gX>-_8^KfN/>-R(V1FM);Xc>,R^N;DQO@WdS#7
&R<D[(51_M_^H?RYN8\EJTBV-+_A<@aeeb-3IO;L)X;Y]c7:RYLVDX_g:LX;Z()C
L8c_.WY[=A_/)2dE0eNRRI]JT26@W5A;V#8>\1gF\0CHKD39AX2aR1d_b&GS8RQ(
WdP(B;S_gIKOH)?V7C1:>V=@H:JX3aPLKPF.-UV63bU20J&6f/JSfgF)]I5V0QWa
#6PP?<e\-YOaW\PS]]V5&&1bR_6aO/Z@97Qf09R/N63fYdHG\-20-IO#P4HZ=>CT
=9T:4;=Xd_?K->@O2c??[?HS651SN?UAXYA_=<CD)g)6;X#Q;#/FORSV\)4b(L2<
242]_)[88EbC91cPc3W4Pf^X13SMH[>I<+cUSa>OMZ&W7Ra>[(#F;CgPAP8GIff6
;X0J<1VXK\\TARTbZP6I5)SI+140[^M.WeLc+U0PM5S1X_ESAA>:&#;I>9YZQLZH
6P2F>-CBC-[.A-PF62.I&,DD0S#16\<7[R@#O;e7XP9HWA>GRX+8_d^b-RCYH&YK
BKVQM-T1,:##P,0e^[QX68dU?#Q.VbQ;g7_J>_=#5^C1)C/e9KAM@DXOUg#W\>EH
,NW:+PO,-Ec[_S9)_ADdI=gB,((>0f7b+@fL9NQ9&cdX]\WO.^:>J>SW/8Ng4Hg@
:/MR[2],e29P6b?)CTb]RH-,_@4<6NTP0PG\F,ed(f=>(1WNe)_L>Y[e+(9=RH49
=EY>53ZN2IGFa7Y;C2V>Y)7KT=O+2.)M<67/9TXYSYS\KEScKIa2;R9>DBQ46UP8
;[3G==QCP^[,,^5JgU47<bb[<MLP.5(;@SWNF50_TU+eeA6SD<;].K(H=LEg.F-_
Og)U#K9HFXDTEP8,C#Rf271#eRQF)HG1K3^BKDXC?PQJVe^]/_dEP9Q5OW8FFAFU
]b\:T6Rg4AW>]),?4SH[/0#W41)DTPMOdf1EV/f6aO@PB&YO<>[dL1PS9Hb+2\f8
3PBCPA\2OM,)Nb)7;/O>MA^Z1POUU9KR>aEZ)Ge28P76a(caaPR,fZ,JVg^&9SDU
A.\Y@]Q,]/Mb)Y\dPZ[P&ZU)@#1FE)[?9>bJHTI7;4.#f1K];PeR^V+(<E#aM&#N
\/&S&&XaB@_VVfUdc-@=24bT(cWb+)E[V,E4Q>c<<A,V[ZfR_4CL(CcQTRB[A,@&
6>RE+XZ:cR?(^^[CPAeO3[T<b0Ycc:S-^cOJW1_W(5D(J7@^caK1MD7>0WR)9H@^
X<R,M+Ud9XOO)e1,I:<Ta&g1f0P;&3XI6#QBK0gfQ12,DL<]F^\<A(eYgP3#5S;>
YU<W#KPD,:8Kc#WJ4RL+fQ>W?dfZLAZ=0HG[4IDI)IS^FCYDJ?2/3B3N^JK@\eD[
ZgJC?7L+P5(g3]D8NHBMFC:L9JGBY,bab3L+/PF:?_7#4&0H>g#FIZ?Had)NQePQ
)#8G@8KPg80&3O[PNWM^_c66MIVLEcO.(L6gf?BadER2N(A>P_W^9c>-,BZE_=ZY
380(>U:HU3&WAH6F^YI>Y&Ca-2\#Y2GdT^1:6e10V:HM2gaf-HMJSeC&6KBdZ9,M
0,Kf?^EUR46Vgc#E-Vf\&\;;:C]@bScJfHKDV;fgQc/M3SCbNL/+KU19S+CYWL^/
e+8[_^;P?d=B66-1#@@MYH8L&Z;bEe&7eCMVQ0[V.).d/0;9IfJGSY8NfSd1d_a5
>X0/5:5F1:=H9V(dV9?9g@G+aXY>+g=KBB2ZFA]UM:CW<D,)C8:]#,:?UfU)dgW)
:>=F)WTK&5^B>>,7HF65_>/PZ.&[LIRc7BLP)+4,XWG1)RC&W:,-&2)9UHTOX09T
C/56c6I_K2,J_:[/WUPZH,:Id97UdAPH#E_0O]\FaQVMH_?C2S+G2P<2#NK#+LM0
<7,fSUC3C>MC?Td>&7\75>R[ED?(FVSfB.\-ZU,:a)BQe)ef[A77O8R<>a/Y#0_.
Sf?f:QO4]G=IE_GXRQaJXR<QN@b0>370U+BL)=PePVV.>:M,NXSeU/AEYRH2WQTR
T&J^LQVEL#.N05@K8YRDB9@<4c])gB_bH?@4Y-6Bd/OZE0b1=8L@6VdW_bO,F1-_
&K0G-FIM-Qg-(_(\9#ZF&A;e+M^2A7W)7-=Q,;dV5I+/73Q+)5>-1P]#01U(#?f8
)\e25\YI;IP]R;:[L6FFQ:RX/XSTQV.TQZ3Jf(^.4^cXTMY\bW=<9HDI2M5NDN/.
9Ze[4HcfAOY)<<64WMD_)@JG=@O#MFbFGc70fZ=Lg:3A:BS-6Z2E^UeU0QOZc_T+
P/V#J2,/GWJ:()1V;/(I<QB[;6QDQO/1<Z45(AeWX^Y8YHf\A:BBPIZUCR7@_.CL
)31+FS5?UM4QL]]0PG@R&IN9c]#D1O:/G?1P\@P8XG<CZ,AN/F0K(@C&7#;91/G7
MeHY>GY2T?)TH__ZF\9P<@\d6H1b8(g#RC]M5e0#:6\L7_BS01L[0I:9/DG_9;Vb
(fW-QZL[O9IQ1/7CQ(ZC<)MCMDZQfe5<-+\Z-THd9/,.YU?(gSCQe^D:f:GI=L@2
(SEKAR]-&5Og(^420MP1C&gRSLD;A,SK4Ob7X+#K7,G9Ac&C,8(6Z;TaL6c2G>72
OC.SOKW7RP50NR6XdLK/fL9Ecb?b(.BbR)6>0+MLEdbbf(&PJ1\@XWXWYR>>(0E(
9X^)3IZT8^;D=AK=HFM5#MKEcaK,SEG2&G+)3MEBW1CJgYc\+4U1X50-ZI8MIJd@
&5[PB]4^OEX1][+5SVRdU/F4)_=(&8Y;4OSLe3VW#>3ZGaZGE]^RSAfUD]U4#N[=
gb(G.R?0BQVYPO,_<g8PCX2>.&Y0\OBNC9;W[4eBc6gMg<VW\&X5deCf0aWJ(E:H
=;(FRM=FP/3,8GIN974:ef#JW(eA\GF+1&@F.@?fZ<d6?F=(dK)-OBKUOC584>EC
9YVPXIFgTPNHS@(Lf\8aSSX2P=PG)a;eg0CW86?aWGDQ6,6aL:@fKA+gUJXDVQ?N
_A16IC2TOM\MCd-7/9:_JZE+/&+\gU(XDF0OB6BOb6?GQ+?TYAZ-a)?GO4XC#JLD
-;bX42DP>XRf8f<_O?SNS-L+QE4846#[c3Y-(aG&fX(,TISF2Q8//4ZA@7164TYZ
B]CF&OBB?NO8#VbSANLA#<Ja\YRD:2Ce5;#D4+8UYaW4C8#c?^HK5R[M2dA))+8c
J#704HQ[gcUe]a,Z>S2SP\7GAfRc(23-9OF)_,a3G2RDT=)/VTX_C_X]1^6dY6KJ
0P4OU&8_C<W[fA2cV5X]L9/L(BSN.#.Lg#K:T)3;AA(=aEMKV6^Wg@Z[7^+YZU\\
d:M6C\6Re]@Q-Z;3HA(b+d2,94YXNBdCSeeV0bOR30f9eNb0X9;W8;VdQG7.PW#K
)N[+I]7,B:[CO(WRM2I]6E:H/AfDcKQJQNXRN.;Q&RWJL/@Y]:M(/-G#+;\\)<\.
@EI<;Mc=/G;IKd[@(NYDN9&8eCNdEa/[4S]QH@47U0A)2R;EO?9d]f69#a7[ZgD-
f7J?d@/0e1<6ddZ):FW0.&05IMSP:Z2)dc9QA;IU==553cHWU8P=^fO,O75@b>]9
&6c>[^^JX:D4gWBe@-(1R&3dY_A-F<]S.8@Bbf#STgGO:QDg(f@A?f37U(?9HGIW
Ie6)bb0I)LUV,HSW7(VC]0/I4S)[Q<;PB2\Jd#+TAHW;TaYD/G<&dN7FX0QS.-(U
A<G99[dB(bM\<SYV-XIE\(GRdR:]0OO<;]Wd105b#T9Z>RfTRWf7g5:O>8,@8]YQ
S9GTD\->(YDJ/74d8K-TA3eWHH\_V1JNaOYVfUQCe8X)2()SKT&fEd(96NVaY?M7
0U99L@>=ILE_2_75\,Cb5V&V[Eb2g+(RU:fMI6W1@?d^Y\S/M;_GB(\46f&(D4eR
0V9]I+/S]c?P5X0,)Y;CRTHSQJR)FOU(Yg7G;=1dUB1Sb:VG0G/;KON&C]2A+=/K
N,TE/;>fY5QM#Q;4XfD-X?:(bA2F/6JL7[)9Y6<)da/>Z6=:[&We0_@]OE,1<@>\
Aa7bH,.0^#)#V.<H.F4JJ;2;;O_+Ig/TVDIM[63ORW;R_3Z;0W,)]7Z#RNE3?&Kc
DgKe(R5T9ag8&MUSf+H^N5[TH7c5b=7^4YO63(Z[D>K?GNKd[fX6VA3_fOCNcR90
PPMBE4S65[&0MW/GV_S;CA>:9/1#<5HO3\7I=UaJM8HD=I?#62QSg9SAMK_6L,60
JBA#()d=R2c\5-V##HF8?R])]35e(9fO9VI6:LVea3JB(3MT[IDCHG1@-^<0<ZLX
Jbd2T1>KO5GO_Mf\f=NQ),gB<OdR,ed;?MNVL+A?##L]^;_XbIcTb;)/HWM41X1+
f&T.H.]V=/UP(O]VeIRHSG[O=:gR12GE)?+3=QV]db9-XLN.;a2\HD.MFE0dKQ)d
6bLV9BLT-c#1._G-W>5UW(U#C^QU&O<KJU5G7gFDNLEN3CN#AA61PXZ\M--F5<0[
6^Ld95-I=3TP4>G4F8LWQ2bOfHYd6fPN?C0AYCGa=9I>>MGd#BefCa19(JXP7&?>
8,:=ag<e<[c,Q/&>ZMI0L):ed[O1a;1\[a&CT(KXJ9(b<1EI/#CPc8ZFEMA5R_I?
/T<:[D_]\KaI(egTJ(-[NU4Z75XD=3Y#8XJKP16C]PacRaW9YTM;]3,M+N;^9ZD_
RTfVeeODcDOIB_0HA0d=\)/V]@W:+RYR9#X_g1c3K5=K&10-=ePD]Sg#0Wc7TX/)
[+>QCHRg4>M2=J6#7(@6>_.G?KA1E\R]\W(Jd@U(c2WKBU8gP(2(&.<[XJXU(C>K
NO7PH\ZG[.KB/DO\.OZ+#7E1]-OWC\_\)aN:?7Yd[b^0FRJVW@[c\IJS4gb)RAW0
)K+FRd_ES-EH-S&<+XFa#-[f4S#X;XZUQ8(J.@&K#YVDG7bKHS/Re<,f.)N?67]A
L97P:Z[P((6bM&CN#)gX18:\>[#DH4/Y-3B2#?/eYI,EN0>6JTB;LTeU-6eeYE6g
C.QY);e]P88UP.+EI348-<?3>MJG\c\73UBU48K6S.EFI.B\NCBFU60CH;54(+R6
<BVUTL<596:6.=MVBBBdCCYcW3]C>GgVa8E>:YgTD->_\S7R]1AL0&J,RN/+]a+6
c8+I,IB8AfaY.&Z-;0GTX[CGB.;I3AR.=YI-JY3Qb5)ZaG>C1LVHG9V\>5g<H,a)
P<H\ND761bB-<&:IX0RDH3B-7+B+=2P<[3WOH)2KO]SGUWX&^L;E/GTG6X0ILRH<
6Z@fM53=.Z8aDIK_42f#<J_H[0XU=IY2g-;B65KX-\8OP@\CT;8P>.ZI4W6N0E^g
>@Xc+&8[Y4g;]SH(X3aNVSSa_g#M(5O^T8N\aa)5/W5JVT1O285F7D.>4BCAYI[=
UYWWYVYaH@+RP6QacJ5179>FEMS@LW1?&4D5=+)]SJDc212F&HPKaP[UDT:L285/
KbL?^fZLe8##ZP+OdSN9J#:M#L[<dDLdc=g0D0[HFK-)O=dC,gS(-OZ4ZGWDB2Kb
g28e:NTP:GR,R([Q6CR/]eCT:I\.[5Wb/D&),F8H=N6D3]:gKMRW.AUS-3X&H\;)
H&U\W#97dQ+=KV[0fVCec8DZ8d+c92HC0]C=0[31f.cZNJ+).Re.(6;B[2CS?B=[
&.^Y)TeQ#eUJI>MN&=,HX0Q_5a\H.VFdb5RQ(5427P,+.EgET:-,VIbJ(MZ<fS:@
KPS9gcS/6ZH&W2J5NeWP>]bDXN.D@,&F9M&F8<@0;1IQ8,#;2]7WC1-[#HSN:ZJa
J8-W>)=B9L+SO]NAD)NJ-(_ZFT^4;HY+Jba^C/560S0?U6^B?c>_B6-/1ScRG_T_
UfPFEA#,;+;5EVcbI0>f=V-=WfEb70[P_GBgMFaL^\-SQ0]<7AI,G;YF5DK.;\C2
U[e_76.FO9JaY&0I/T?W:/B17M+[.I9UIRI_1_X>ZCWWCeP&@S#3eQTf9494(5.@
eeA-&</-.UO.1M0W]L+5;3LK3GAZDIPKDS.Z]OW;H((@(ZW57Jb?gKNVA+1VY:#L
RGc0M>c11d9MWE5.SYT#I9c5I5NKIJGA)^@D?BAJU9B>6-)c26S,W-^H[=9-<H):
AR)(X@:MK_+,6X&_+D)FS;VIE]ORe_#/bZEH<@EYR1B#d7@SRJ#?,RT[]^61]:+W
(?E2G7+ZI)cQ;Bf/+]e-A=8@7\D\b#W5AM3)C0g3f?VO20M9d9QFP=Z-Q-c@X7U>
Z/^\+M#=D)BeH>X80&5I\_I#aDTfD-7YGIb:UW<;1_;fdN7ZNd+T)GPf9G)1,7VU
_e/(cV1CJ&YH9:D0<AQR(:V0P@A&FeB8QT\ae@<SVf0X0/-J\,#aX=1ZDBS_BR6T
P?>L07IBQ1C>7F#E6G8(7&0)Gg5X57S/8LROFP;C2g^F.cZ.?BO:gf65g,?faMJL
X&-E@^0J]>W0G7J7O+S:B]ZVGI2,]7=&eb2GYTA-L-+Q87H[I7@,[IDI7e^c,0H=
F=8OC#:O(c>#)FSIJGPQCIZEQQC3Q59:2P?V3=@4B-Abbge.^,Q#/EF78W=>MHaL
62H;J4b,]DQMLIf:G^^_>6JY,(<A-0.N^G)TG7<@@+HLP&+F:G^S^SK+QDVf4=0B
#&5=59F)18OfgYJ^X)=1S2,LN#JbFGLQ&D^ZGJ9b6ZT^NM6J>BUF/Q)Q]Ed4bO[Z
?-URW&LJ@JEGH3.C#6,T#(_3)5C3J7ee&_GF46IaUJ?(CZ(g=F=]^:>\1Y+\+)MS
L-J5b46L,+WBOUWYaW:3J<L/]\L\][@)Za:33,IP81YMfJSdga,gaCNKXKHSd+B8
TL#P2[eaE(+G,K\:O&/0dN>O-JHWPYgRQ<_dLgH3\\gE09T&b<_fb/#cAI9F7B)C
.(X6HOB2T_W/E]bS#]L(D=N36ZX-1NB[34=NZc,,4,NT@)ATU;8]DXKdO]NQD:OO
3&KXZ&,?OZB?#CGCJ>Zg&-^.X9BKQ56&/BZL:7AZ7QU/=eJY7LK?M/8.cec60S>P
4RCZ+9,8:Q,6)L0X[VK)<;FAC:CWfC@O:Df1S+bcKO6.FF8L\,8UE@S<:\-3-f&,
-R^;UB0J3FI[G=T<M[3HZUX@7:&+#C[/_=@=Y;]O[T>]?Z#6QY+Y#bHeM=EO5G;A
IV@-=PI2#@1,f6EFf7;bE--1e&US/F2EO6(P)Xe@gP^TR[KDNMfaL0e^7QJ?I,_6
/F]M#cZO9)a)B-EG9,ePT6F05\7+LX@B_S/&>_\U44daA_>c]186TE5EU,dQZ/GE
g.5\A.(Q@UO5a<G@M1.BK)Wcf+4+[He:2>N7c:PL4O5ZPF5&#Z,.B1dC:<LZRd>^
U.RL28IF136e5:M#Z0PSRd\G;:Ze:JaNaT3Y6.JeTNXNJL29BTUIIXXYT_=8;d5>
c.6?dIR^PKDIabH(Z+;<e539g@A/9)a?7C:W,I9V/70TP5+fS,2M.B_B?\/9@YaM
M3,O7<=WT90]^5-DGRJdF.:(\Z/:bTfD<(S+5@5RXSUBU1@#=d(B7@]GB:=KAEXZ
/CAU-9B;&7M?TPTC#,->[04T4Ce)(#dA>9.BcA93B441&X45g&NgZS,#W2Q&I&Pg
APe(eA?.Fd,XWd@#Bf<L,B&CfXP-530KX#<AC=8Zb[9eQ5>M1AgU<BO]a6W_]>[F
+SB5a#FJ@>?\=S>:R#[.(6T8+d7LZ0(6A_:+,MY_&gQA[O8VQ+(@D&I9d[DbKVY&
CFc0_=K6cH9QPAT)4fbTM]57+=CceKcg.<?&7>_^ZIf/=&^PbJ(\f394WM-2FRX,
K(2]CEacM-g4DWCW5g<bCKB>,A8LZVbMX6Z<_S=d(K-XUOa)OR9#_?:V\/<]L1=[
0JeDcIT=HfC_X@,BW=63K)KCZNDS7C7[E<(#,R[^)S2>aa^#fc91\;.:edC>LdD5
;+_,;cC]7,NNe98T]ABBac^b+B+9E\AQ4^Gf6Kc8?I,Xd-ce_FAGOMOZ9P]Cf)JQ
<Vg92HDLXT2JcU^M0b4gQS/YIU&LBgVC-^X>#LY5aM:@aEc-04]eMMR]LbW=6<0L
^-<CS0#L@U9e/A1AOUY.97bIYGYXIbP6C^L:.C<TQ@0NAQd=<[DJ:MMDDA[a&@_#
3E77,@R]:H,O3^1#d<9PLO)YaSd8ZQ?4c(7R/+BCMCS/SU2a?C;9=1LE^(&:IX1:
(WZ-U,V^HHJ)a0Y-5:C;HB_O[4][1ae20>7Z.TQVHBbDD3UYF&URDJcG:4_10A>6
:,1L02?9/&,G3AI/a,0WPBTLS6e\2dIL9ag5#dXVW+6d6+]e;Z6eU^--@T8RW46X
HJ.SP=KgdMR74K2AGD.aW?1ENL2B,HT42Ka:2XSCG0S)42Z2?A(P0OeH27EPfKYX
>=>TQ3MYMHJ[=X?X5[G=+-R+#b(J?EHI51DU7?^Kb2H#ZDeMWR4[-R/SbcY.f5?7
cAZ:T_[+V?6&Y&R.TNC64JPJ9KD0;gQOMU168BO]dcT^P:P1@8O0GS^RNSgW_Z:7
ZR6]0N]=7,8\:3=f;=SNGQ8c(X^=A(363U>UGJ_a?EI_E\0J<S2WIO87c6/4ZbV^
#.3&:VU<B(/4PUMa@0=>391E-E8+MVX/Zc7B6N/(>S?FW>?46MI@^L&+OU[2\-V)
/@W.QB&N.O[;>R1FMB(2:5QS>6-UBXSTP,<0f;RUTB\@g5R=Db/_8OYB79fXNT(7
K&(AS/FD1Dd4XY<e]U+V+C:;d:T4FL_,UD9-_C@/D^Xd8GHb1SLBWOLRCO;Udb6@
;S?AP^XUM>/<e0P7]RgXY5?H?C6K>.T,_#cK(U]@+K3R(<5GYbdDf@/0R[/7FK4c
PT(&QOJ:2K#PD3]FfCFdWV#-3Y3N1Q]@(W7W3C<B]7NFBAG+f+WbULc5dL0+_LY8
EIFS71f60MO@C(Q1NIc=/)&Oc06D95Q/ZV30NKcc_;6DIUcLL_)c_L&,)Mb/5bJ>
[GPGJ^GPGGLCR627#\Y2TV8ad_04>B/5P2CZVGJf9A6ZSV8aWVK/YH78gFDf2L0,
OO1S.RIdF2[M(b,<CW./I,b6H<R/?6TY19-Q(]VO7dZ)G:d6<3SF=84E73E9]@Y0
=,7N>QE73(H\O71[EZNRa9VR3M2<3,>G9/FE8M<3SJBcge1JDHD4Hd04a#HE:RU.
+]S?INKc1F0>?YeD4976KR-MS2>VNJMW@3GQ@U=8a<WB55IRUSY7/E[MMWO8LeX]
-,2&46]3&N^gQ48T#cZAa-&d16:Q;Q_^QOS5a-TE+.]86.cfS/QO;)M1,2=Sad/&
H(TE]\\<>A9RVZ5(CeMMJ]NL,);U\f9d?B+@U8MB;TF\_+YdR8M/5QPKX4e.+;H3
GXS#F)#0:Sf\+E7:J&GOd-/39BgP6C1TM5Ef9d]CS+.CAW]>#2=HBU^>g=F8P(;S
>b>Q[?0K6FW+E#)]E,R?DeRPPQa@P:98DY&b_G&\&?]&0)G&GR9f()GP[aT>d:PF
?FecMb>]bW)a]fUSI3_SQf8[e5^0[IO46.fNP,PAS9NI[A9Z:;b>,c(@6^5UAUR@
4B4HVIf1>>-R3Rb(5YD,3-Q6:(?>TRK-+QGD4[7cW.FP76F0aD.TR.b3>e)I/,Q1
3Ufd;/]WQc/_3dSH^FIDa;N+X9#NEA7RTV\QX9[41@LQaZ?+A@([f3>R0)aG8e<3
fD_b5f(BBJUb?LK;<0RKB91RAE42,=MGZ#^<HbOd&8/&DSY\5b@K41d-)9[,27gC
1IQ\\Y(U[ZR9D]#a5X6KI[:D8@-+N?Y58#I&/CfYE6bTRBQ@g^02a^CdAUO0BY?+
NG+/79>-?OV44f[Q[c?f#=TFST)g63?AbNRB-RV4c,,=^DVc.JQ+S7e]:Tf\6K==
IdFYN.JGIYH]\b><#^T#[V6RT)ABJ@<2J?6TZ+M/+SBVfDcS;8;Z79#3D4TM/L]d
gg^I:4S?G6PYaUad[ZTA^Cgc,@SbYT<T\Jfg4Eg]9@&GJDWE[5aQZM4O=3\AJ;9+
_9KY=^R6VXV9S31U/2J?EIJ>BW@__56#-b619]#Xc.DGY.DdXJ4G9TVE2LE=]aV=
,g=_DeQ(3:7ec[S,;JWZ@#W1\WQIEA/I(HN_VL6?TaZUU]\UE.92>3+e,-UER:7.
NJY)UOX5S2G+KY+^/b0-NddPF5_71?eSOO)FD^+R3@S5U=U<3I?+^VT^S^N0-Q3S
ef;T2-CUdKNNLZD8.(SSI#&]Y066G?RBU]dF]98NJQ)0Dd;9gRPdB0>04cY.YU\8
9YB4[;C>F>;5T>G+0BNTfR&,aG]\LWa+#IS5\61F824Q^L40F)c@:O3]7^M?SSFY
G?X<(F-VYU[7V35#XN#6b5JJYO3fAFUL3f]caQFIgXK]c1<GMNd<P6e]38+^1])9
U3>9Z&)A8U2CD,T?=7JHe[K:b(1/XbU^7DQJ6Hc4\=B.bNEL7(dMY3K7g:&_<AHA
^SAD24e(T(TXG-H,))+GIRED+3<TFT[,?Z^HMdUS33/&7CcHAMS1DII9cO[^8gC/
_18W0d;EIF]fQ]RIS?g]#&A2a^PQ9+H#OWKULUG>]8.VK_E59bbFH36T1g1SLaD/
1]:NW;7cZc4cG&><(9BaAO3&2CY0<)gGU?9-c4NI^JKR/O.#XE;,BC?)a?][1b7X
QZVXQXS+>O]5(P+&\+^Ug7FSN1YPd9JRe(?fWgSFNTVUg.+0a4=b,D5<AfLO1/fF
^S68_Yc<L,I4bf]+L,dP@-DV?gVab;L_)gC,=C?]3WFeK,>\.):P+ES^TVYZA_R,
fR=,Oae]MC7Q4Md7KLFJ+CIgf:OE+3\c3HcI\INe4@f+?7@:4/_&=T^-0fB.6fg\
VeGNKXU\.[3CE#-XH89c=CW)&FWJ(-GV51-56Bc>Y1aW@>E]X>(.GdgUMJcIO>8A
UMNcB1:5XaNY+FSD3T?IW/7^=d&@EW?NO,GIAgOL61.IJ#J+):M2)JPeQKYgBQcO
&C/RTYL,Q0-W3YA/g@[M6TSFDRSXaW@c>AcZ=+NB&.\AKFaCE5Y6I?d[\(T/R:1e
SBND7PL1T;E@LP@V)5]TUC6^290:7Y,I1?DaWAFFX<XE+L&gY+->ZF_U<[DOdFGI
&K_49<A)&;cL-2M^)5#/>LJ;H_[e@Mf)?TH;]Y?&58&,@6MfIW-D2f0KMdCEf2R;
)ZHI]7(SR:M1][cPZM_0W,WGQ2Oe#D2;f\S9@0R&d=\T2H8^4RVWSNYXZ:/NV&H#
@a]aR=26d7X_TTK9U<@</3RBY<8<b2/1XT6gN3a6BUP.aC2#O=]^Yc8;U(1FfMV.
L5T+=aB[13X=2F]65G=d[-]NW,AcPDHPO4d@)d4:H&:NeL[7c/T:JBZe2HQg2E]6
.3AD?]S>a2X,)N[IfV3X1U)G]+I+c@Ma(b)WY@#KQ@QKE-E42TPKLc)&H6>OGFX\
6,Zc+-Y5ca/;EQ4?,:1&=R2/H+X\PbA-1+3LaYOE_^@9cBPH#@gXF/.13JG-R=-a
:U@CIWI\6U(MF--b1^3?/JM@U^]Qgf5FLJ=Za:GY5</IaT5d_LYJ#-=UZTf)M#U6
e:\4Z]<6@b>c913H_P<<[[F/7,;50I7PUF)R@g_OTfZ>U4H7R]S0_?cT.:X()S\b
IX;\6QQ;Zc0<6=:f#Q\5Vf5I4L8]+0ee>X6(<TgBNb#+RV)+AD(JIOF-a^,?HccZ
1WQ_/?I#@OJ46A4-e6;._?fXgV#[D=d)<f<MUe6:&a7H/4<fbZcPVVY9^#UD5]+M
^[IC?a>QZGbNG<IbL,K>0^>++aN[Y/QddJ<2c(A>CE^4bQF@,?2ZS]?VSNJDJ.8L
?S2(;QZO/]9DT;d&WB;#7F<7cH@BEP,VP9KUI-^G\e/d7+CFDc>AOVME3LC@>#4U
O[L/WGB#gV+(4QHeeeAAE:3&6I4X<eH6UA#N5;b8))TZ9X>>QH2BIL]^SU^RQM@7
>?3]R5&]PFJ=KU.J/d+3HB/&bF)Zg2f+OQbb#Re<0#[4#JDU/aI-_?.\&8W33b,b
?:6SZ@Z+bOd?#)5gGXI@]P?^?3UREL1_UaTJQ#3c[(5MBHC=96Qa@/dFdbX7I4IN
KRT5a;T@4MJ9U75>;VG<4gVUWLE)&GD27gZ>&+X+<_H)^I0SeWV[\0J17UT6a)H9
U.-baMLIGGeA_Z,U/#2DH=gaa8O@UWO^0>P,)Z[)DPXWAW3fE^O_6(UIA@e6e/??
g(S6F:.<=FG?R9=dJR,0eNM(?gHR&&N7FNQ>;A2R5&.Z471^2O)-Q=B+,AbTb>W2
Q8SE,POZc&.QYF=QFUXZ;_3L)\7g17)@Pfa19G48bM[bcdgcfI<)bF>N,2WR_+WW
@?_3<QI1d>7-BGDLW64MfY)Sa2-3G5DCc0[XVX2.(<JBSP_NC6[8(Y?@M/P;&VQ&
B\C&3e4ONd7+XgaPHUP:D0aZIY-H=S/5)(<YV\Ace(&\^:=PAS5f&_ce[e9f8@\_
1XLG-V3H)Y+HI3/O1NC:KKfd+PN4<IQLRLOQDE=BG3V8_X?4^&4]cg@Ug;02Q#0d
8]D22F..OaE0#,&+b-4?G:8Yc7eL@B+,MD#OS#&/e83M.I.RTV,DK[M\,>#VJ?P&
]aP[)7af<WPQ:9\,&Nf.6J>F>[7X<<]cT<0]/_DUeI###Od82R_IBYC^gE?bD\,c
51f?IKVMR9daFD,-=aN#;8M=USH<?eKcJY?.+<8#-<5_aE\c\/ea6B=Q\IFO(_U-
aO?&P^G.])9Ub&QI&J<(NJK1VWePa<0L@ddAf-,O>6.[?f5Y&[K#)JZY8^H.9\KF
O@IPZF-ASVb<FF6Uf^O=20AJ+LX?>_BO7ZJ=DE9V1;7c[EWfC)1aEJ]TQ#Db;4?F
F:C:4_:]_E@9&AWR4Z^,)P)X.;;e>F@#E;A8TFSVf#8&Lb=I@,RZF^XO.FZ7cdKM
G^@-(ECTSc.c(M&eV<<3@MNcECJ+6fZBQ&/d0e:ZO)/6G.+A2B#G)CZU?J=bJ<@X
J2CY?PQ]Q+#?SOR&&1b9D>=^ZRAgdVZ/I5I1NfPEU2?M<-AZ(;8_Q9>.^R?@;CYK
4E?&&[cOP.3#1UF\MJ1M?#WH;Y;?9<OaTUQEQZa,J8+F,HS3YY^>5T@_P?UD:bI5
[M=UHH<F(<a3./]NE7O:3C-6+068Mdd+FWc_-H6V5SZ\MZ9JK3QU/+X5:(#Y;KPN
R0(gbFYe<8+L0)X4C4P.X)(REQMG.9\>>XBVQNBGf8\.1[5,cIF4;R7P^@U6NJ/B
>L7UOcK3Nd>?W_[cD8IFE8C9<(&.FQbW38&UYA#44?AXK5W9AWAPK4/@<_62bTDd
)IWMD-R@D6f:I:0]N_)87,TMf/5<EfKTfPM96/0KUUKKRGG?6[I.4/L)g.(>55M5
P]5f&/JK2[c-.A405]#0fZdAQE0AT8QB9g]M=NbRQAc9DP;[5#<3>:BG;C=C9.V_
Z?.+fa+I#-G[XLPRO^]AH)aT6d:X4;g^aW5^dSAAeZbX]I+\,T@_eX).C3bGfV?Q
@R-\7(0AfP31?A\L<[SP(WWBMd0@[V:U\H#0bcD&@-9LA==-/N3(fQ\bBAbc4T+#
I^VX#7B#JPR9D)>24=F[J]S<KIF.:RH+f61aDXBg<a]V2<CeU\1ERHBW7ZY7,.0<
B#IcXfUDN2[A.70Q^9DP)e@JK?1E=DKN6;+RUOaANV3=WCV(+WO-I/KY2(g9c0W5
<_N/CY2d5NXU[:J_^Hd>H<^]>b/.?W4-b1,U=+[d-UZVHP)\>c4D?<Xd64Fd\BRU
5Y;2ZU>,MQSIVR/X<5RafTL;6EACe)f7(4A,AB+D7SZ#9N?LS8/M/J7D<\SN9F4M
O0&8(H05WNS]ROgGB.,I:1_:dJ:1L8\\BbHaSbK0YbO&R+;BJ3>P:Pg9WV)717&>
E96,+ANGVO(-1U>I.3[W-Y=(QGJA1f@4C&AIB1_EI^-P#DRJIB,EH=G-Da>J,^[4
7bD-W]X(Z48,:0b1e:[P05K^=(H:<T+X7?,2cN?.>3e7/9^[:c@ddA10WeU5GI(S
8@D1&0VcD\LX(a^(CZb\F[A]N)]N(EgM6gJ8A@/L7T-3@T,?0,,NXC7H2aLUPRA,
2>0&6adIVUA7Q8a)3I@5D20&Z3URJ:D?Ld^>54/+HYO7JED2=Ibd+T=U1FUHYb,J
7?KG1@62>RSfYbMb4K0I,H-D/#W]B9dDHJT(YfM3aU#6_KH.&g\7VDfb7d#ba-9B
F&5M40ReA/MG@U.A;If]J9aWL=&?]Z-/4+3_FCbS)JU@=32]G1SCO0:H^^QB[SQV
5NeM-_.b?@]=LMP)(eEgO,L2A2,Z7XdKD?&&@+<TCT7L29B)ADUZLeN;bT707NUf
L?UbHN@<g)@LNA,JOFV_<92LLMUR[AS#2=,Q&AAR#Z21X)-I;@7N9BB1)ea=MWb\
NN?34e8_YD#f#)b/Z)[)a@Y:.1>W(9W6FYASBML#853/TPXQg9B4KMY;)dPM<VC]
X/L)._QA/NSQd._gJ4+E\_JD\Jg53YS:G-:PBI#0OD3MU?+6-1X]JeY_S=VaCBJ\
/EbSKS9-b42_&bSB7B<7=fM)@/68O8@]g/^6(:4Jg5?P1K/H5Y<dMXB5#8N-,#,W
9@PJ<D6E0a#&AFQFH6dEgSg9F1Y@Dc6V)2cWUI_)edOIEYY+NN(1U/6P82UQbeG4
N=W8&M&?Sd:@.>4V:U(@E+?.)FIBK<\GcLf.+,WB4<INc)7>>,dGW6_K,0.EB0(Y
4a_#Ba:\O8DI)0QSU><5bMN6:(eZ0=2.fQ^F#N2V)44(H.DC@ZLDF9SC,81)LeK/
^Cb<B]N39eN4N>\[W)L]eSaH65(N)C8\=9\-Cc4L2HF/GX?A<bB5[C-3_DI@P<:1
B@5OSPE<eM0[8#B<+[004&TIU0GFIg_.MJO^O8L<4=579U(;/3.@(Mb@BgAZEH3\
[)=7.V<O3/0>#?D7CV,:F43<ce=5LKSRV>_aAd69-\Me_C6)W=JQD&fS0J#dKNcM
@(0?Abe.RKW1<+d28B^M?\dbf[7Maa9Q[J#HG^<JIgFK.97f5RD(U/D5C5K>2:MW
BQg9JJF?e:>b2f4\IJ9&XD\,=Qa7Hg5HJ6\85),Ddac(B>bZMS8BdfVKRDS3UJ_b
+W9(_,:\fCCM+GXc?c27^#.HIS(NR6=#H>0S:1S_9@J7I,)4A]gGMP<?8@557Za)
_GOFf=e4@ZUJ-PQRKL7,42E=_42^_MVbE&M_TgBLY>NO<7.0U0X2^-DNCg&X2.NX
XLWLDL2O0O2QeWH\(_/1;OFQ2:fTaOCd2VJ)7@bU[;BYP[TK)_.^<I.).BXNAH,&
)V-&\b:B3de@.YAd1HL]/+4IZagaC:]R4aZ_)@=T.GgK9Da4<QXRX<7_a.-R;WI^
1/1@EgM0^@]Z8ADPJ_++g:5#BRIGXWUT60<.1_f8PD&3-[-]FIV#fM05HOX34#Xc
6#L2;1/]5VK]EVMa<>L\2-_SPU=<S#LE74P;]6dE\=&?OQ/cNG>P.-AAK=FH5BW,
MT8D)^b[HgH_gd5EaJ4PFI(S>TP7M.g#aI07P8S@FC2]&GG]WM//^UG)U).?:F&#
cbPTU/O)EE_AE28I.,BbfN4J67@5LN]gTG^@HX>AFS1gVU7@M6SJH&+RG38(<L4-
2DUNQCI^V(8S&aGdWJ&[/-Y:RCcCWIG?;B)=DY@W^W-I:e6M7J)\Z,T+d<.QA3/:
/aVX?;/N):,9[:M[Ye^7S@a](+FE:F^BAc_P0Zc?K@LUKeJg#&b_DG]GDa5FcUE4
PQD_WL^[+;SMGUV?Rf+[).[U\F(S-@_8S@f.N]>I9b4^5T87-@\UGe\<LfX0Y^b)
-2/Qb]MNeb=eNO:BT0dbUJ]K9SK^,8;NZG;&N[<gFT:I_MA.XEGg)0Y@=-)d:f@:
//bH;gbZGYSX2&f++Q,_(g.152K54-8RM/U&JaVNH8SC=X]b=9&.W<O1C)NPMRYO
\)-KZ?41>QY:OD5:JC]L5CKA3G@MD<>>,>W.#fCNc&L=&32I7D[5[,c^,Ia2/A]8
9C&BR#VF1S;d#/K9Z-Z]<8M(>9TU\Da/MB@Q\TY&c^=K9K7VQ?H2/dAL&3ZQR5M+
[?CF+6c4geQI&2gTM5<:Lf=JQTVY\Sa1V]UPHaBOBJJ1BH9A=+<L[+:HW-ZP?:F3
4@CJ4:^Pg);N2C;2;D8d:-5.X\f40cdH9T-Q/.&WeQO>ab@1cf71[Qd37[X,#&Q2
_WdL]dB84[/ITO/G.;._51]a@6ELR7>,>CSVd4^eU13;UW9^<4:W#6SATMS5Sf]b
.X>G#=J]-?6aF0=KN:^3D@<U5Ne8GT-@1CHUb^.YS.RScLe,B=^E?=DWC(+ZJ5bg
NQ,Te=Bd(U8UIG\fTQ.S^+E\@A@(RJ<(5L6H-V_&,0I1MZ/+F)U2^YDUd,R:f0Z4
TS4S7Gf<gRRaQCE+7R-T]A3S_A]Z;RN\Q3<=RQSg7L])[_F)L7O<H4-]V&c5&eWY
H(X<DXU>1)I0W,V?B5<4:[@:LbV/:[)99]5M13#A68[ZI/SMZ]\W)XG^O9OC+&(4
9ER,B&[5>XPO_(\S4M/KHg5?C=4gO=LW44D]-O)Y>eK16gU07&YWOGD^LUG&Z>gf
fQdZ=O^6=2]\WP)HH\(##e[Z1OQ#W/8AB:=7fFQH+2LDIEg6^e7fAM]O]LZ5STQC
7=Q_IRBRM8HIcb4>]0c3<1,OKF>+I[GZ(HVS^bFAXGM>&fX/V^;aG-=c9N#?>NO/
;R>4[0Q+BS.SA7D+Wd^JP:Fb)>3-@A962]]=V?BH^\Y0;:8/J,C[^&98,6O_Zc3I
RQbbGY&>=(]WRW<_ML?ZXLF_WX)&/YAd)JL/=K-=Y[XO-J)_Xd]GUTQICMb@2WBM
&QY9EcW;37]6M76IW\T))]ef6=9f61OAaQF.R1c9aY;&CVRGR#4@.=/ZI=/G/VW?
]B;af:0G#X]P&5Ue0=L?bM6FP+cUM3^]b\87<99I^]+)@GcRJb8AQ_5KX.<#b?>#
PFe81I6_(D<<W,&>]O3MJIg_D9O716,8-M;aA5W4/&/DcE6NARdMVWSX6&+_QFCP
;V0BH2P.O&?Q;>2:,9<#CWbQaN,4-/\c9GYHW7RAJM1;2]Qe=&@LVgc)P)V&ScN1
O2:[Vc&P&YYgAB].M:/20?[2N]J2#:?U[=Ge[[AQ=BcM>M1,RB[<R548PI_E.9cO
bVD)F7[;FdQQBX^Z-#JLd[ABCZP2M4&c8^gZQ+G7;N<D3\d,W<2_77<-JQ0[46^P
/&U9]Z3B8aa4/XQf&/d5>MOFM@\-Oced2(>H#SgW4?/02M1CXV^40eRK]HB.R7=Z
=[E:)2/#51:Z9I;UC&W&Q27,aHaE1LE-Ugaf05g+QbRI]?JHb+VH\G<:b_GZKGU&
5RNc.e7QeFUY]&J7R<bL1HA5PcOIeF)42L#4MG\,E-52WR2YHBG[2P3W0G7JS0#;
=(Kf@9QW#/_IO[DYRL/VE196gDKR]^beD)J.2MOc(FJW2Cf10eG=5]c6EWg#BLbK
K/8dQDaCb&N\>fR)#c0_0UZSTA^-1]@aPL-c3N4QT2eUgEc>,;?I4Tg(aLY.,@b8
HD^c9#:2Jf8IbU:R)72d;.]HA=?\.f=ALUC+U@gg0eNI9B;_)N18P;8S:O-S+#V3
eL7XMC#QVHaNTYJ^f#QA0(.2R-+dUFd]M<1B,F:E-Ba4YTHGE,YTg2KdMEAH<^BJ
;XAT.3H8&S3.3(4,Q,Ja&UF]/05Y^&VU2FLL=:29E=H<f\;PG.ML85W,>QeAO0(M
Z+)X:c,7C674.+&(ULS?VB6c[&38/0P\9Q:BLb]A[-1]f.H7:fe.UP?1^@,VdN[,
M=XUbF#RC:SOc7)O;WAT.H1;4K0Wb;#]0,;JZG5K5,EWUaf(7I1X#=]6;__]FVX-
?6DQ-JZAZOMC30A(FIWbD9P+eJTJ.=E.IS>^34#1J1g4>5DAPG=&-&DUL4APF?QF
[F;VeE9:.5),AT=BZ@-OM_+9;WCP<SN:dQae.N]RPOQ/7I,6PT1GDVHdKNG?[cdW
YbVPce_T:#0DW?eC:1T>40@X:Ie+dPI_>[/[PJGLK)>\MFGHJW/&BR+QKe@=4dd+
Q-3TfXfELMYB&0Q54GFa0W5KT]K6<@+eg<(#2Tadg1A@T<A>J)Z-M7P).(BHI+=8
N#]\S\\3VE4(D+(7C9.,?+BeBRVJDY>972/[UMg^bBa5-KL6ga6f^dU2K+54gA?:
(Ne+@CQ1M0a4.7H<^OION]MRc;cJ3\[+L7+A[TNMPdSATO-VXVL+ab.B&HeS(K37
AR^O)fb,V<8?/27dfE-#aD)OJ-SHR2<7AW]/6.F.HHTcaRX#D9VZ6L#APTW8+,BA
U6^N?\E9:=(E#?NE3\dTJQQJ^HVL4/8:/B(N]^A_+c<?>C>D3:Jb3RR_J7AA_E>?
N&>9JTK.)48ISD-Va;)VM4&W4-3.1JJ>eE&./Q1>HMD)]ce:7Q=KNH2G=5K_IF.)
1]@2>9<_;GO]&7+.gY_^[7aIH.T)QX4=e+09J7I&)JX(UFEUg.].+Q@7APF-9;aX
T[N0SVH,]@XAU+dRD#Z#HNI1H-&3(If_2TF,DXFaa9\E_2AO)&+G5G>MD/<<PNee
]>gc?\Kd]_F/d<2V^[ISPSB-9dI3EOAG]EKA=gD/89adS03NMAJLSMC&^,.R>5?N
JTbeY=Va=\G:,Q?b-43DRSKMHNN(;,HS+,2@4?R[:8(N^@)G\_F3V,&<:e^c?BP^
BE#R;QWC3,.,Ka,NZF]U5/ZX&[dX4LR7/=@X@+S<J@]_R6O:>6&Ib<T5PNHX\#5R
c\,1BZ\/LP:M&>g+_CX6)daL[ZO7QK7K]-(06S;.\+):Y,Mf&PG.?#KVF-&X<ZBG
N7b4\;R+MUa=-C2H1H7W:c)<LV+dL5eEa9DOD^4=bN^RY_g-F(6XEJ38+e:@(g;W
aYEFHU;8d7FYC:0dKDY4GVU(US.?e^6HVR>41P,a+TT?&;<:99TR7A?24I<+<aQ=
7+Y6FRFLA?AeOGS50dX;IQ[#5R3K@Ua_H,=..67Ug77,)R)#A+;W;_@a]GN:XR?K
e3fWbHQHM6^9g,eT&^/3IgWbFPIb>3EBCTX(W?Ma0F(@ZG^L9WZ2W5:aW<,D@=b^
)U;NU3>&>e);4NF:?3Y\A_[1L7Rd:0H@P1YVKT]J>,@U06f(dKUCBYd^>Mf=gKNG
S(Q]Za8[#X9#GF()+g6/6UEU-K6YL4:N5>3aDfMC68@c+SB?f^TE@56:WBNB,C&X
9/R.14?UCJL:X#QL>)PO<fQ0B?0?;G,#Z@0J_@BQG?C.(RgKREa_f/@R07@0Y.R=
Re+fJLVR()J-J7,c7:X77B/AHaE-,^YY_@afIH]_^KS8^Q<SR+JV+.],PO/=?];[
(_&6>X(YKE;CQC9S2]#5#1OaKC7ab/=G]LXUfUJZO,d)PQW-<-EMWGg5V/\R8FS=
X&fH5G#bb^FP5P).C-<59VFf_^9#H1QKYb1LDD^#fcEg>OH<];g/WNDg1-Z#T0YP
?9:R(BZ<g#_B0#aNJ].3GUeK:<=5e/A,PC4bIX:Xd2GQ_HFDO>T?AagLS6DMDK/@
D,C7Q8C=D2&;af&SFbZUX&=E\)9<@YS9KGW44W1E.M\=Z3K+fD8I0&_2KDM<WAWE
Fg92-)B2UFg5;+GUGZ]G)O7RU7;7D&J(g,2:OL\+BM^dN:]WQfEQ>E2J437+?bU2
\7@MC;L,2V,;JAEEY)III>SG^CJB-R0.WGB#Pe(JBAB:RKMA>0d-&0Tb7#JQZYYU
TgPYV0Pe[Y0f=9M(4PN[>D:>89>c5(15H44;X^e?7WWEM2Og3MZ_OWdXCDE7]Ndb
a52PFX1;XV<V;PYK\dH5I.Y<Q->].K[W.++@1Sf^9VF5.CV&X<:VL/P<.O4PYS\O
C=J16K)=-T(W1+3\\?US18M,39ILHHNS#705W.2\;<7Wg;H,(D>caNO^V5+XS4gK
07F.7C_ffG2I5+Le#g<[2R<VHJAF^I1Y/AF1O_]d5:MOUV>eZ)#]]98Ne,O(B.WJ
:1<;I2H=7g.D;+(MT[B/aWJO6VbCUU8ZKDOICH(5&9BZS;:@[]@@H/YA5;e3H+Hf
L5B+a\cYb7SQbDJ[=4]AK=fT993L?96GGLXSI&f5P:C=94ZYbD[gPc2a7IdX/U&/
:FfK3D6,.RU:d.7\W,A^]V5O&FA9I>7H_,5.c1TecMFTa(d@gRLKG[Nd^Sd\EaTD
g,4>WP3RLc>V^)a#H:f3^UP8M6PAO.d>X/LYERM)3EH7XUZ(.]:_Z8D#G+<GKA)[
19#,\;(U[)UV:<LLDL&W;UM;B,L(W&=^ZKa1/aY3d]g4-X_26]I7;D_W]:52V5dV
3PWBL)]5<#&=SK\[LdJ)G2UV@3)g=2N?WE?bSPbE&WHAX&;=2XE-I-E.JC_?7dHQ
\T-g10721TG(@D:(JYNb9?H.e#)G\IR.CO>4dVO#V./R5Y?LW7a@\^-<@GMIG(I3
21ce\PI9eDE+fBCB/4bPRbKH/-gVA7I5,Q7^5bE?=]ND)-F4gJL,@\<#KW]C0WM#
^&LGVMD(-&H&V@()a9I1/6MeF0F[7AZ(UZ/SH3I8[_TV.G.:V83&P4Y]4@GZ;7M)
cJ5W\_PJH0=6>Bd\-#93/4JEO[NGcXdXBH:RXFH-^C:\.&e9B(K8d)I;I]<cVcIe
I<2_+_FgT&9A[aaBTQ.)+OM]DBBfC@AKHe<Zef3E2O,L>UH&dBGR5EBf;ST1\Z1E
&1H/IdLf9Q;P?NJ)fHU5Y/ee34VfA\SX-G2RUYbVS;8ffcWD[US6T;)c89^,ZO?[
5bV<F]R0\PIDBM?^X?\bG7[QH8>F<D@[cf12DA9&(I-W(\DbO@Xc.=6,C5)f1M7\
E>&aXfN^/+ag7bR>I^5Y4YJ;9I7HHX+Z1.7#g^TWA=)26,Q</egBb.HN5CbcMOMF
+WFT-KV@aJA1ERgUQ8LSd[XPXD&X,3]L#_5CeWR#F=.d,R,P5Ve=eY/WPaQC[Yba
78BN+(gR/b(F7(^;AGg#/;XHY81IB;a^d.B)EZ<ATfaLU.U,[YCJ>,#:g))##&NG
gHC[J2LeL[SEAaF_VAHTdA)&BX>SaCK#@PIXbM=gJ7=38NcWKM^&8aIUgcYbMCDW
NY:Y@Z.@bZ79];L_K3K,SR(02RM^8EW8R.N71b;aP;MHEf9U=ggC<U@2IC=;R3Od
CH@L/E:#(2BZU^O-e=5&G0(D5eEA0H88&:f<1:4XLO&P=;.T[5.Ka;XBPKFC<[/[
EX.D8]cGKIQ?b5;d1Rg+d-e^3Z\T&FULGE[(7U-,M+Pb]4;WG?]Q_TK@YK\dHV7S
ADF?Y^8?4)=D^:TdeTA=0<(44H<P/7FFC/F@BY#Q1PW:)@L+<(>b),+CD6G?\F:X
IEM;^DgW,.Tgc,XQYM-.E/-9H>,WI5_+S=+G[;=7LI4>gJeJX+O8+]L&0\5=c9TU
.^U;#J#cebeA(ADX3;Bbc4BY3M9UN6UH)TFEd1_/#/=Bc;KVI][eMK)e?T:P)Ydd
5NAFM6G)\bf7FV?):TGIb[;J6;5a0MI[>2_c^VDH6\3fID-TYDFa/E>;0JX9,c^:
L<[=U:<RCA:490\>JS0Y]K>W/]=Uf/SOLFC7(0<S?MG58ef3dg[C/cG5)0U=f1C0
f+Q2,<7b,764XfO(6_+4ScgK#S=g7LfB:c)ZLB8)[5eMFYWF]2;Zf<^12,Va=P7-
bM[]U;G^3U8Jc6M^T1H#=<^Tfc,2fCS0]&CL+DN(]04W&<FbTVZ28g:DB+L].a)B
AQYS7&S8A@AFBMC0?Y@dS;(W^4Iea^-1-fF+XJbX]a+>d@\;C2:94^IH&2R]-EEV
XJQ02IaQ>S)?[)Fa)6f&Y.:N94--@3[]W2HTBf^_a?Fg.H<fE,;L_H-.<XN\KS?/
1)>@9S8T\9f>QcAMRY6V:b]FOU1-;NK4\EU9a^H:F7/7H5[^D:I?LF2c(19]cU;[
E7\EFOZI^APdJD3)&F0M53f3Lbf4CC/[2gV7GcYB=:UbCR(@PaL>8-0RFTU>5^&T
.,f&/cHN-)#&B@C0Q_)GP>OTONb([Z,P-:^M\K-.cSX:HEfPME]D#Oa<>PC+d/<U
9Qdd>2;V(dHY@ARPP[@/7^/V=B^4,-;XKSfG3/,>5JYT]E+D(Pe-R3C8ZQ@6/fB-
6a_[B5].#4]M,6d&7^WYeCZRHVV\GAQV;_N)2e\eT[@1B[OfOYJ@57f2R\;BPAUL
^dI:DXAE6)9L.QCLY&1M38\=>0/F3cATDED7ZQdZHL@aVL-H1K14H7WR4HeOD3J>
;4)[IDIA[>G)=.@2RQW=(:Mb^\NDSO/08QR:CFQ,5V/Na1-.J7-1_g)))cK(bME/
4.V-d(+:GI]GMZg[03H\VP9;#9MeWTN(3N+]=R6-1+C:RSX_](T5TQ2M@(R>E@7G
=73PYW?,;#[cW+M@IKcG(W_\/g(+^gA:>-G+372]O4,Cd&G>0#3FY=f]Q;\+96IU
VHf-Wfd25C?#\5@.c#;8+PA&3J4>e84Bf-GdNQ#)I2LFa4e#gP)/D)NMLG6X[9G<
[M[eX@MV1O\-3d7F;X@4FXK_D[R9>e;FgP[8E]VO^]54I-,.^7:/;/<6&bbR6S_2
CedZd(^F0XE;M?Of;4b:?=S)LZ75&gLfeS<TAH<?ELNQf:#KD4_.?W)K:45NAeFW
HC5QA^#9P>IZfd_:[@)&CKP0^LP,F3TR--YD1=:OH:WW<b<Y#S3g4(>_2<?<7#+K
(gR;B6KR-S@2&NXgR<T2<g47g8_7Z/GPEHG204G+[^=-:Ob^O&?cTEBR#R>aaS#=
,_.D1RbbZ4ae#<Y\M5H_/:dY>fALW\Y/WP02V;],&<E;f81Kd8dNg49U<.0_1X:#
PI+1I3Y<7;D5WUHWP;eTO8b+,+Oa-<@L>@E4.&PQTc<5)\0cQgL=b?3G2_aK8IK>
+RSE>_(,OA@L(_aS1J,d<=OdB9^RE.)8JK?g.:UFPJM6FH24Da<9/7&0;d00;^DT
(2Eb8X6YbYWN4_TKOb>+,7N?T<7Y2ZH<c?gQ&Q.TLYLNU.-d3.9Q9XJ/F0KbcM:7
/HL0(V_T]#-;7B#L4#)9:bYfK7BF:?b:Z,^,QR(gKUE:O)?d;A-(^NKIA0-O1fed
8A-88c=NaBC/SS,?S/=VL5O#bKUUeXdQ7PP582gS#=^(1_557GR]d-L[E6;.;Z_F
+MLT4,+Zc[G3G59Ya2)g5JMEVGDP5S]M)Fac7A.3XK<)a\F,E-F8F2_K]JEgR0VS
->7([NDE<[02:c--H>\6;4]-.=A=gQ3@PPdgYP\ZWZ&WXLO>6bIf^-d+I:_NC_4#
10-,XGY[0H[]3R=)CZ1<J\\SMb?(<)I?L7Y(1#RM-D4Y?<V8FE;Vb6(\,d))TO-?
9Q/G485/:QP#gXGSJW+GJ+:5__-eR>EXKZP3@-67)H4VBRN]TR&+Y<+?RI+<LJ,S
#2RU@ScW1cB_MIUD02W;Q)]cM,0I@^-7<c@0a]I.]U?8/T[B]bg4Ng;TR<8SZ\G>
MFA]eZ\<N3O#<KISd((2A^I9YSfDA^RZRJHZ)>1\(gD]cN-W@[K<_5P>A19^g)2W
cY4:Ud^C^@P;(9=fM^X+dTO3CFN/LP1/:$
`endprotected

`protected
QQFVR<.D4:dLJ8[JOGbZcLUD&B7/1Y>86YOd>gKfA#X)WE@OJe=]4)A6D5_0VgD\
1SVW6H2eTb\L/$
`endprotected

//vcs_lic_vip_protect
  `protected
.^6=@)2TE;M(4U=JdS5NK>+6@I1@Ic]XA1)PG8(,5-:cML=(gBaC&(A4Yf-AKKBC
NXB2:Zd?]IO<4O]-d.M@85G\=KNKO\BVeRD@)CI[G2@NS<YUV/g#25YS04eG6fCC
K&dTS1\M@RHR#S>RJHUR9;#3bRK=IOd45FM+U_K<>,aW7,:EFK=DE1SfOZC9<))g
_:3_R3\[62;I8IYZ13H@;ML,-<0e.AT)U__:=.f,8[02(D1df,BTD;Z<Yf35f4?e
?I,dfTG..12eN@?1^EEb^g#7C[faMW=Z[>(I&<K;@1,M:H:B/eLD_,O#?2NL84FU
5SK_SO?A16SD9IVd<QTTW<a124^0g.+1-1AgW[ef&<SHT.\Q9a@08X5b.egL_0@E
L]aOYH3K@WHJ8aI\?Y2J3cS46WLZG]JN6@@PPGX._&.^IWNSOb#PeS7X=@4.F)4K
acBKF9:PDCTQ>>AA&AC[/>/2?1\24KEYd(VHb#/gV]16?#DUP5?,VK1G7#-&:VB>
AW;EHHI,dDb.M?2&;WWVbK-2XcK7HOa(>[Z\^YaXgKBg&G,PfMeN+MP]&8cV2a&Z
PYc<W,CC37aMN\#5ZT>(M<,33\MG&XdQc7H7Ic\J#T1YGN4P.+;S(>IM.e8_;55g
G^;:&O]QdJb=P1+23IU+:WGU&ZVc-/d,&)>DWcKQ0:2.W8@A+@WGfK>b)3KCN;;]
1F_3[4cK)Y0.[VW2b,37N=VeTYHZFa:T1RJ\ZD(8XAgU4=2B+:G8=^O9+g\#?OND
T?)cZADb(+[PDC6.<JKAPY.Mf^#c>&Z6_[+C1:GJ[CF1?EY9c&fe?FB6?0g3/-6+
]92TK1J-TV5W1.#McI2L.deP.-f+R+NCTB)>=eg3S3=CMJN,g6PPWTPLXa.44JgI
IG>?U7dW6.33+L.IK<>50G4#7P@a-PaO,f#.4&d@3WVJ+P(&C,-QZ.HS@82QWZC(
I_(>WBaBM\@N?-30?^]6[[E7JWU885A@3PFfgdHCAHX)J21O7[RD@2>@+@gMEa@f
ff-.-A0?V&[L?EHR6d#FKf[>E7?X;T104_K6]9.DUECdAMG7[(4(cAXSQgA6Y/<_
/d?KG6\5D->e^(Q9XE_8S\#]OaZ[K@72S(YWZ(d[e=Q7+V63RJd];P>O2(&c\4MI
)8VP8NWF03R1<:M14&GI^VD5RQd).2,;P0E#cC(]dU_=:G_,@V\,Beg\&&D)V,/U
ee0-V5R]Rg3UGQNB3Y+gK;Q4T??:?X;BSN;TPMN/LQ,OG2M2[O&)@\:R/,B:PA3A
O.SbEe<Nb1.2TSN\;Z0L]/A-?#/U)ZM7_[_:ZGE<QLJU1DKTQ-Pf/cG8J9XK#\T/
4-GBMQ5M,=>Q^CL1WE?_3Q=I_6Of<_gFH-66ORaSZcHb#A6f)N<VSB.=U)N_8BaU
_,@3=\>BW-E_7R6,<I=W&Sd1J_G=UKD.;RI\]^AFEO@GA2RP^.;.QaDV3\2?W\Id
)b+UKKJ-gF2#P.a1,@5Y>D/@CQ@WJD3\DgRd70JC;[/Z?]Sb3MEN)eTG/eEC=0_I
DF>4BQPc(DYC@DP\CcKeAOK6)=SF++Oe;442&N^20\@_H+#3T[6=Z<S[f0]17W64
#V4#28>ET_TZRc9MZ)#OSGH\2JdR0Af@D(+3A]:ZI#WM<UPaNd=@;Z2?Q[ZU0T4d
B]X.1N>Qd,Jf3+^b]5Q]F]bbK>61JC:[.\D#U>+X,033bPI#+UCeH8SUN7&G42GM
Y#]cAC<)I.=c/I+9DP<-JT3eF13+L+F]:HRdEcE&?].ALLLVNQ^b^/PM1):GMRB0
H2\I]@2K45JeOgY.d@QUbJCdRagJM-R.#<QaAe>.D#.1P9-9C+^#D0,0Ea=PJ?&.
<>2-aA6.3^(MFEOYe;UY=VI#KXSPVJ?((9KI465HfX:JI1cYNe\&F1MNa\/R7,R&
C@f_IKcLC.;2EDRR_TSC+5P3AU[R,8Z7,d:\F5T7ZMY9-^e+PUc;K3/6[_7J(,Y.
#Y#OVP_JS3N[JF4dYKUW<G]YD;WN]X3a]8MZ_2Hfc8^Q4I2LX3_4[g@=(ZX^XQVH
EC8@=3^+8.R]S9LX(XN64CU536,=Z7/:,AFF4,Sd()8QR+^[>86L,fPVQ8c=7d=:
.R9H@Jf:[g-ICFRI#L\fHeV,e^W;O^(O\:<bDW@<=aSe8Z0Z1@a8g+5;a2XGQ?^+
3BN:+02(cR9I)$
`endprotected


`endif // GUARD_SVT_AHB_SLAVE_AGENT_SV

