`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
QErzkp5qLW5J3bTLdcdtf80YI63gOzKbbb0J8+gyr/+mGiYkXYkUdA2dktE0xQBX
SktCxcxWSv4h9kld1TbaQGWdBrpDuMwS3vVo+ZPtxfg+DUeuwMfc9d7wxVnUqD5a
8/mBwF1DG+0ulCCvqX6CJeoUgH+0iX2/lAAKo4nP+Fo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 83        )
tstdVYRyejBBoeZvb6BAoIatZ4vm4btIehzFY3Y83g4KUkKLPN7lI5SOAovMHmcS
Wyroy5LlmqBEnFWK/5DA80iwWIJFVKemgaOqYYxZPn7u8l7MFCUA08jt+vRYvT64
`pragma protect end_protected
