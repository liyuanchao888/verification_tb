
`ifndef GUARD_SVT_AXI_SLAVE_UVM_SV
`define GUARD_SVT_AXI_SLAVE_UVM_SV

typedef class svt_axi_slave_callback;
typedef class svt_axi_slave;
typedef uvm_callbacks#(svt_axi_slave,svt_axi_slave_callback) svt_axi_slave_callback_pool;

// =============================================================================
/**
 * This class is an SVT Driver extension that implements an AXI Slave component.
 */
class svt_axi_slave extends svt_driver #(`SVT_AXI_SLAVE_TRANSACTION_TYPE);

  /** @cond PRIVATE */
  `uvm_register_cb(svt_axi_slave, svt_axi_slave_callback)
  uvm_blocking_put_port #(`SVT_AXI_SLAVE_TRANSACTION_TYPE) vlog_cmd_put_port;
  bit                                                is_cmd_cfg_applied = 1;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  //vcs_lic_vip_protect
    `protected
>V)<7L=0IN\XTd8-&)XUgST4M&M\Aa-U(L>FV3M:WPeNaQ@YEGFY5(.^>).M#VY9
=R=NUKMZdY-<<@(1L3fI5#NP(./([K#_HQ,G8BbfB&K\7@XYK0Ia(G6W7R/2f4#Y
..Ba;[8+I?]fD+EC>0?W,JY[FdA2:O#+A&[N5\-TSK6,MM7-a1bIB@:d+P8#7[dV
cW7g#>:[X7>(6b=CR&5BgNE3gVRL1ZC&g&2;]I):B(G27a3/XKO)G#ZA>G?0XaA/
.^Q\B#g<#?T5E3NN_RV+W-^Y,a74P,(b+B9OOX^,BVG5c=&^?XGc\Y?WBf[]M8UA
aeQ\,/KC6<]CGI>Ge6)dd_\253O(Tg&>Z39^?Ya3C3S98A#2egJUFW+ENAdb#1IT
b?4WfP4[Z]BBXA-b#LR\XR[b]MO/8M_BWHAZ=\9e=<aE[9N)T_+4V[-5f2)5:>N>
P:fU]b2[6T6B&AF/:8DPQ9-d7N:[?D81/CAX]1M#IO.DS2]8FZWQ@fW)ScC,Ge]4
?2?LAD47KU?HMT#E&,]bA,-g2R<PGY2)D)7VBQ&L4d:aYc2eITQgV]]<_/Ec7G->
SJWC>6,=cW1JK79.Qa[E-IM;4/OV[96f)+F<<PdfGaHfK?]EV]T+L5@g)I/A+.a.
b+:/DL(SgY5?(cVMX&><BGaSd;9IM<4Ve_BK:a10-&>YE&YA2cda1:c,3A.T<+^]
ZFVR\[C?HA3bDTF1#4DW+..6,a,DB5+QO&+.C]KeA..D>+[eY501CSWU((ANZYS)
ON&V+fH>_BTKeEE<Se//Q(T:8=,)V?N5/K</(d6OCaW96Y&-F.8(^:W;f/[^RDJ4
:)9CE&W05RAW=M[JSPUI3cE[7N9>E8?^:,aFF2,>N,7GTLa/6>/8DQe0862G\-bc
&U,,>7_Uc[>f>.U2MB<Pbc/=\\#696ODaM0/SMGRG\72-O8HH4\:EL@R,DCV1)9f
S/82bT/H5JKbJK.1&9=@G/a\ASfL(9U5.LA&(f,g<CN;D]McWPbGX9.](bHWg(W8
Y)QFL3,8?UMS<#[a;IT),)9XYW[cT,2G(IIP-\c6=O:G]EX;Q)I8C.TMbLLQ9XB/
9aR&(AG(_98T]V\eC)+59EcPP6Q:84CeYec?Q-bdLSM97WAM8DH.CdXRO;JOSBF3
5@4T^_cRce,N[aOJOb9b)[cP6$
`endprotected


  /**
   * Response port provided to supply respone and data information in a delayed
   * manner. Refer user guide for a detailed description. 
   */
  uvm_blocking_put_imp #(`SVT_AXI_SLAVE_TRANSACTION_TYPE, svt_axi_slave)
    delayed_response_request_export;

  /**
   * Request port provided to supply snoop transactions to a slave port
   * that is instantiated in the interconnect.
   */
  uvm_blocking_get_port #(svt_axi_ic_snoop_transaction) snoop_req_port;

  /**
   * Snoop request port provided to allow snoop requests to be sent from the
   * slave, using Slave snoop sequencer
   */
  uvm_seq_item_pull_port #(svt_axi_ic_snoop_transaction, svt_axi_ic_snoop_transaction) snoop_seq_item_port;

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  /** Common features of AXI Slave components */
  protected svt_axi_common common;

  /** Configuration object copy to be used in set/get operations. */
  svt_axi_port_configuration cfg_snapshot;


  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_axi_port_configuration cfg;

  /** 
   * A semaphore to provide exclusive access to add the transaction from 
   * sequencer. 
   */
  local semaphore add_to_active_sema = new(1);

  /** The process that runs consume_from_seq_item_port */ 
  local process consume_from_seq_item_port_process;  

  /** Variable to indicate if the consume_from_seq_item_port is blocked waiting
   * for a transaction from sequencer */
  local bit is_waiting_on_seq_item_port = 0;

  /** The process that runs consume_from_snoop_req_port */ 
  local process consume_from_snoop_req_port_process;  

  /** 
   * A semaphore to provide exclusive access to add the transaction from 
   * snoop sequencer. 
   */
  local semaphore add_to_snoop_active_sema = new(1);

  /** The process that runs consume_from_snoop_seq_item_port */ 
  local process consume_from_snoop_seq_item_port_process;  

 /** @endcond */


  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************
  
  `uvm_component_utils(svt_axi_slave)

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new driver instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, uvm_component parent);

  // ---------------------------------------------------------------------------
   /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);
  // ---------------------------------------------------------------------------

  /**
   * Build Phase
   * Constructs the common class
   */
  extern virtual function void build_phase (uvm_phase phase);

  /**
   * End of Elaboration Phase
   * Disables automatic item recording if the feature is available
   */
  extern virtual function void end_of_elaboration_phase (uvm_phase phase);

  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads like consume_from_seq_item_port()
   */
  extern virtual task run_phase(uvm_phase phase);
  
  /** Report phase execution of the UVM component*/
  extern virtual function void report_phase (uvm_phase phase);

/** @cond PRIVATE */
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /**
   * Method which manages seq_item_port
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_from_seq_item_port(uvm_phase phase);

  /**
   * Method which manages snoop_req_port
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_from_snoop_req_port(uvm_phase phase);


  /** Method to set common */
  extern function void set_common(svt_axi_common common);

  /**
   * Method which manages snoop_seq_item_port
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_from_snoop_seq_item_port(uvm_phase phase);

  /**
   * Task to drop al objections if there is a bus inactivity timeout
   *
   * @param phase Phase reference from the phase that this method is started from
   */ 
  extern local task manage_objections(uvm_phase phase);

  /**
    * Implementation of delayed_response_request_port
    */
  extern task put(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------
  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void post_input_port_get(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the seq_item_port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void input_port_cov(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving the read data phase of a transaction.
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void pre_read_data_phase_started(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving write response phase of a write transaction.
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void pre_write_resp_phase_started(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_input_port_get</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task post_input_port_get_cb_exec(svt_axi_transaction xact, ref bit drop);


  //----------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the seq_item_port.
   *
   * This method issues the <i>input_port_cov</i> callback.
   *
   * Overriding implementations in extended classes must call the super version of
   * this method.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  extern virtual task input_port_cov_cb_exec(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving the read data phase of a transaction.
   * 
   * This method issues the <i>pre_read_data_phase_started</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_read_data_phase_started_cb_exec(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving write response phase of a write transaction.
   * 
   * This method issues the <i>pre_write_resp_phase_started</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_write_resp_phase_started_cb_exec(svt_axi_transaction xact);
/** @endcond */

  /** Returns the number of outstanding slave transactions. */
  extern virtual function int get_number_of_outstanding_slave_transactions(bit silent = 1, output `SVT_AXI_SLAVE_TRANSACTION_TYPE actvQ[$]);

//vcs_lic_vip_protect
  `protected
8:g6:Ng>(Ac8O_B\[0+-0d<V,\I#a@EfE6E,?[3]L,_#MSWG-H_>3(+ed]2)Pc.<
cZSJJQ8(AK1Ud6a/IY@<5K6.dKU1F9MY8Zf7[/_@SeZO8NKMO>(NC8(5f3RNOND.
d3YT3L5H+1OfSBFb\>:JIMIX=DA8NcRTU5::Y28^PP.cbEe+.CGRMR.\(Ca46UHc
LSG8&EE-IM[1<[)\Sc+ZQEZA8P:-KM;J@7J;S][.&#E4).EU+=U3P.D\UD053a7_
a?ZV(E5(\bOb#ZT15>;KQLZA4$
`endprotected


endclass

`protected
a]HNZ6cSY[)V>J<a<??f_g7Xf<)df_&fb]#1<^[701fX4JX4XK<#6)b7W]8MD[8]
QfPJYC+C3O3VTeED.^/3HT_@H<bAHASMY&##+eG4g2.0E]cZ(\D5fa]a>S[f_4U8
EZ=&M6fWQB)(6OOF.G)1.2[)>:>CU-ZHg2QS7.)IT,.bgefHD89J.4FI7#?W\^c1
3@S^6a0DGN6RO[RN@Y,+PJ^?INb?2,DT,;\IXX1J;\J(g@VOLC,P-fU-X)2EXLS&
M260;5>f^&SRf)<5L?(c&QSUKIKZe)4^1ELNTLT/G9RCb\/6M(,J@;Y,3K_dN9=M
J:(cB3:DJ)c0IZZ>4T4GAaPUC6DW;b\YecaY&IdCD;[?agGefR@.V_-#UdV?e_aD
L?:f>#Q.g_RfJ9WbL8HC?U4<2OSUb.G[7NQaf3bP+[Nb,WW>9D[ZZK0/@]EUAf4G
G&FXeE017+Hb]^^3.LU:Z/<P#e@QBI<FT3QYS3[H?-T.N]0CMA4LO#OYMJYNBfQP
\PF]c/YUPV>\V]W-::afYf7^>H@/:aaW@@A?ISA@Gg_GbQ7b2<\&?>OYL$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
5)T62MFF+K]W;M.I8\7dHd4_+?C7a;=1\I3Ba/eQCc_MLV=e/A4.(()gG^\5SZY@
RDbEI><K)#\17AOad>HZ((MWB&4^_<dL_/0ge?[gN?/+3I?[(4eb19T8eJR2Ba/3
[3EVYDZH?1],]0bfE1/3B1>/HJ,,8#Id75,>C3=-=?c8J=?^aH3O11cOXB4G/M[7
+d7#6L/A<=O4[IEVX.)Q<G-L77K:Egab+]C-G5[>#^^AGB#R.@OfUY\ZVbaGR+4^
K/),EG7;c2d5T\2a.(cC)1XR.^,RUgXS^UQ0Nd[E_8@B/@eQID6+3K8_AW^L+39e
_fYL^:L&J81ZddJfCZGWc3dUd/5BeF@G>+)^BC-gD6[_1X:^AF4Wb>\NU_WYU&@S
;&(f9EX1YL4;6Q>=9Ug\fP,/^5)#/,]C/G>ULPG(&?T#-0--VZaZSMa^\,J8_,E&
WQ#Q&ZS:CRM:LU6D0?Y=[(QBMae;==Og+2.<FR.&8Ye;<b3:6Nc<H8BC<.b9F]>D
e4@AH=XJ]cB)WK(6>/NV52+a&D[,[F^,>\:69DVOfZSQP5-]N244GSE8\^@+QS>9
b>4-]UM<I..,&;J\]A#]_N-QDOd=.9JQ3]HI<[c8XTO46b&;(c4@1fO(COcNfR_W
d)LAN51P;Y6GEI1<#U&OdL,H=G3f)Ab+bf=TO9_6W07A<O14(IIJdPL)(G2FOK\=
6T?6bCcULE6e=Ag#P1_]d)#5U^b<?7e2&GHYVX=+[1JYF_&6,M2FR]-LF/fIRE2E
^Y4[_CJ5cQ<2#e<JBP0>-3LBfBR/PNed&27.ASScd34>\.,[L#2L#RY#9>^)Y/(2
I@NLBd7^V(FLWM9?;QH2+;_>;TTbV5V=&0Y_GTWGa?9VU/eDCP8\7D)<84fYI\AB
#L</6O>BX93?RHQ9L:)Q(QgZ4?ZZUd=DCO+Yb:+@1BG#E\2^9G/0@MA3630FG_]W
FSS6+/bQQga97QJW:?AEdcBU7]@IS3YfI,@<&XF+SP>W:7g;c;&>];921:>(N6XM
b0I3?YT_Ua\9,,bY]R,0C@Kd1UGU80@ONUcfe^D.T>a+C[]P+)01EMOO=)WLYBNP
?#^M<S>1+_5XdgMT5)@XNZX:M,4Tg8V4e\?PC&cFG<F(2@[PEcMKWOVgd@UZ84E0
)N9U(-WHC>_#bJ/:H73Z^^>3\32bLO@(?MCXMG6?X^GP(ONf/YDQ+7KNJeP9fG-C
f^9[(1^F9\\1/QQObeVRKZ(4COR4Z765_Y?#e@(V&M^S=_;EI>-MY0(H)=V-EcY;
)@.U6DWgaCW0KaK=,>IM,JTZMAR-))eLC=I(AEWRDL2cUG;5CF9T:b0bc^7-4<OI
[+;&X(<WZHa61Z5,FNV(W+\YWEZ+H<M,bZ5<]_W03,ERG2-6;CI172MCI^4:YLC5
UG;5#42?E6\>c^1&>&.-MS7V2(+ZCB:?L0LHGUC@.;YNe??ba:/,dV,CeOB]NDTS
PH;eW-.F7C24ge>&PCNC_[Dg(=T##L[8&Uf^@d6\I_Q7VgTT]NbWV=\D:Se9IO#8
c[LSEO-,eB8HO@0GW444#XEg/(F;BWIICED7V/>9LCGPT6;+J,1BK=6+UUgFg_D-
15c]c>/#2<T1,dZ@+,&930[_c0N2R;82YX.CPDWe@aI<P6R>]&CRY8GDI77,eOD8
M)7-cXK4d@?JKKRIb2@K1>H\;O>b@Q^IbT31)H@OI+b]f,gY_.B[-W6RVbRaW5O5
HbG[&5dU3F?(A/VE&SZ6aPS#?\=/II09<X]d;S#Q)ef=[K[XJU)e2_EA:^@5A:2^
QAP,XP+XE6O2F(D3f6LK>ca<TcZH_<=_:_2aTDH#HXB22f8)_8._\-aOHQ=24@&9
&(B==e+^]JdSYJf.:-Na/2_#c<4G<))8^XZcE\Y]J\SR5R2J>b^FZ[DI]d\&ODVA
d,8IS_gUO1dV>g1461I>C.ZBG3/,FHV1P;0R]_R)9e(g8K6afN6(+SY]NBIO8Y=U
AZ9c7K_T8]<e;NJ,Sa#a,[70H^I<HCW:@aCGZ<X9d#[]@g?b5-e-[aC2Ff<4:T\R
:(O6:^ZUVW/OE=<3Q9O2_&-.0c3(WI:ZP,8K8]15bNUQ<ZOb@F?0?EdY;43I,Rf.
]3J.OeL\<T?/P#27<SQX?2bfKf19O)b+6E=dQG\I637?:]17:d7(?]/F[IETP-L?
W&XJ<,+(.\9V58^U\LF<IK&#][TJZ>?L5HD0X4^20NcdAO@_DE4)C4dT:Lf=)5<N
&OK(0W5?^8N;?eFI7?1/#</.GDEfZ@3Y4-?7117<9e&S?)]Y#LaW?1HM[?SUb_b-
^L2a#S/^[T1ddcSU)2P4I56V5KQ7MKX/<I:d<8/TJ[P9^_CCCU3cG6(W7Faf+@QS
03EWQX<ZBTga0-Q6;cH3NVY02\[I9X]:NY1dD/UM=Ib=DN+:4BCHe[)SH12F;3#G
TYg97:VL?IDZZ9JVTcVbOe(#VJUF\3\CJ0,&^@UC1cWO0XOgG8AS=XCFOQ\PMR8@
14YC3EFaAT5Y\Q43g29Z8E-\;c)/(IM>efQO3=YO>?=^A5@_F_O\)@Y[&eCH25c>
d_eOI2e7a=_2Q&@D>MNcI]Q^M4[d/d[DBJ8\RgYY@XSO0UD46OCEYZM0]V/4C81<
fFE(F<NPgd4/:<WYe9?1RF>NdPN6GQ4&:_=J1BEH1Q,KA=UL^4fMLM5FVTV@2MI-
IA_C:.P\N,=ZG,O5#IcDH\)1A@)Hbb[-GPCD(526>C;CB5BFUX6E9(:+b6SQ];LJ
,:SN2a&]8SL_[V(]<a0bRf^0&W#a([-E=GF,NRT#T;7Q;[.[Z[HF4]>KXM+eP#b2
[Z?H5O-)YN1)6ZAR8K7+[6^0XZ&RRc&HCKL3MU?02G;-c-a9e;LTb3=fN:^;U2E>
d;3CJP.eIbEZQBHILP&b8G_(VM.bEIT_,??F^H]G<D?cK<Q&&M7=<GfV<8;+,<Xe
7;W5a14)214Q2CL6S9a>L7(9,(gS2@8NaW:#3<8OYUeL61b(UeE5Be&+3HSP?)4Z
3fg1HOgHY;JIfMOPIeWSY_dfWQ9;?ZTU)/O5?S/Y3fM6Z5dEf00Wa-.MN\+_g<GI
+Q0_E\O#P2;U<7O.^W@2IdU8e2:Hga._]E,/Y2+Y-g+;?+-9GX4J;_eKFO1;HB=X
Ra1.],B7dP0W)f/QZWAIcU22X.FJae?LGGcXF>S+TS_0DC@9).Q1^[b7N3TOG(e6
I(=7)BR7Vc@#@]EZ(\(<+,U?Xf@eAT[B^O(8_]B^7g+9_,LXG=6IaH_\\LB62#dR
QA&31:#-F1@ZM7gO[CdT^IF,b\J6fI2aM6GL@>V7]9(SRC4HeA&BC_eB24MWebAR
2e-4QeMA+UM0e[R8KBO?M8UYfY=D_Rc4F_\BS.8g<8T\.^+aTLE,Pfd,#WKa>5KY
+6T(L50J1,=:J38NQ2>)AcAC;d/[C+0EFEG]@bFbF<F49^)aBbe&^B8bgf)c20ZH
LAPQ8@&S8<;:#LV,0YW^_bf9M-^&HO,]IOf=._2402bX:]BI2J_E51,f<8[64S,>
AefSGB3S5>a6;,AG;R;4C427^&_QLAP3KW^cg&DB0[7SG=_gD2beFc5e\7T=XgSP
,+]OSd]P_H,GQbJ4:AZcE-78=8Eg\U3EPQQTf]UXS)L<BDGEcEdU]F1+J3V?;fIa
Ea;T)6&4<BZKXL+TGeGNA7U\6+Kd0(]Z)Yad:K[EJ06J)^TA-OFP^6d:6X4I@?]F
L;L7Q4AWC/MKZfg:>e]T[/(OER(XceHHG[D>>cB:F^6:ILdW[8JAYR&7-CF^HKd5
H18)[dB:I>gEYKg]=9aNg?7GC5bD\;20G?ZIWX^/\X3c^fVf<:f2D,79_]S#_RUG
?Md>.ZS/-^T<-/Za,NBU=D<T<4b@3XMC;8:6PYOLAC]aD[Y-GCPS^a6&Y#?+;=P3
aX5<OPX-7VU6NK3bLZ^W/+HBF0+>DcH^CY]OGHc[G+HV[-fT7YHdZgZ#,Pa_O#-<
AQ>-_Ze3g.AI=-d<,Of)5D[OD@[H70I?5)c<#P>U4G0K)aX3+S(WI(3>f>0+R<IO
V:b(]V5OVAf5[P:5+N8^40K9?#8U\1P.ff+5c??fJeAe,d18=&G:,EbXMXe;?=bg
bKV]\e^CT[Y_XRI]Ca7\1=;&?-#P)e_B^&a3Q;1KBg(,c:WLJ7Z^_RW;Y@4GK8HE
J2TDG\2>\+>><+]8S][WfK8IdP.A[<:_RK)Ig.B.DNHS59K887460ZMbD==3T]OT
&<4W6:E\/;+#GLMKS[Yb1.];H=O]<-1FYV.P-X)WXK0<?4]<abBYb:N&6_Q]7:0G
0\P#1A-,+]GbED<U.0,NGR(\d^-LIK)IFHK?^.a\A[D\,D(<Z>L0Q.&Wf5ec^V^/
&Oe1(_PL/]&S[\RJc0F;SLbM71MJQ6cU1]fWEVbGRIT(fPd),dT4C:dP0[4(RO44
Y=(<Q<M(g-D0E<B0D;27d??a<0b^39/7(4e\89H?bPJ8#@DL[KaAUM8/,=J[;?=T
SY(5Q&PCUM9O6K07GcW1Qc36\Y]&G4_J.T9&1][-8\fea7Q<)(3XMFQQ^C,R-(C9
,JfTTa@dO)ZI#/[Ug;+VQ/A.,bf4N4/VFPF-W\P<6[4HX8J69\#0K5ID97V1Y(K&
:HeG3_M:49MZONBUb\f,[dL5b=+GH<(?XZAK3^_BgT_#b]3.;4(&(I_CBE16VA+_
IA4/fWG6OFUH8:UEMd&Y_Q^4QOB:\BcNH<QCJc]:+H4A1]AQI<?NW><@+SA##]Wd
_@(L66GHFc73VO<f^(ae-XHDQG<(?A/68[8c_Z&P@beH+=[17SC-CQ\7/+_-e0?Y
V&#gZMWb4GMWb2;f#(R1QK.3,e>2Y4SE1FXP^bK8?)<7^O<]H:/,d?]-cSF+^A::
2.)A@b?4YLT:+]QOLf;aO##,@EW#U<Y:;X4R:KdeeBN0<0d+I_eJ1:cGL+d5NGD;
W&).Y.-CUYFFGRX=4=#c7IBGR&+])5_RT811SS>V7B@#_TJCOOOXH6(a#d46_;=3
c^&J_[)Ue/BJAH9XZSDWTfA8@\BIZLP36[0aVM+G#0\>JYC>:FDVA_&gLc8[D3G9
U_6VV\?,N#38O]D57XQ@]]^S3ODceD0TO=C>[<Ec(bbN(V_2L;,eO[4)WG[^GHgX
:\MUM.b1AONN3ePg<f5Jgf@;B9.HC45+/\V58Q[gBI.(_d@C?USAa95/dWe(G71H
HA&5=Ed0XRYI[1O+KO(O&X->_g@(Zb?P;35#P#O:Z:?ES\BM@4FL8(AT-Q.(XDXd
],b:06L68FE7W2[0OcaXJ>>Z;eUMTQ4SVQ6=aEQB]8)_/@Pe@ZCIXDJ[DG(U,@Y@
OZQIa20XX>(RA#8Z79]8CU>-TO5F>L,FNM^RZ.W]c9fcTb(U^MCf0;M>,S29MQbO
>1:aV>,INPRU)?-;@SL@&VfEBX8P(a>,PMZD:Y9:UZUgENKG-,-KBT6dHLB;]^]^
4dPe_5<?(5QbIZ(M9>_A24&.Y_@ZVJbGT?@A<\K(Y&4JQAH2,gDWA7/cB@[Rf=-P
0NTbR=TbF2];P69U8,/(XQSADC]K46e/-f?DS[XRLfB9+e@)O9g=H70JG:eY39\;
1:JF7E_H/7f9,4@[c4X9YJ2#Q_XC0_3=dX7TGD_87b-]-e.+KQPdV;W]Ugg&6\0#
R]=]LYa^gY.K4-@@a](Sba+=[\+I(<FO1TLDO5MT8:Bg9T].CMY&8X<B?Y<#U?Q9
]^X(0KJAU&P9gM1.W0_P7Ig1[a\FAeg3L?^<6HA=@OXU@<d[>abSCYced;C_39LS
[+B0AX^@f73b2LfdFP4\&Z]<@=L-G,:aTbgLR3P\R85Y7B/\gb>?g)7K#T=TOSK9
P7S8#[e7]6)\)H,ZP2c_f4Z;7=c-C3\L-b;;7FX:O.=4L^RdG0g1&#=<F?6?,J@T
[@IQE)GY+OJD\(f?de8\cQT+HFJQULC+C\egMe93<?GWS_T.ZOX?;MSWFPe_OS(Y
?5f5JYdFIF(<a^4B8KBg4Pb3QJKc(K6&?NWA<=]<U/Td^U^)D/R[c_aPc&KdD+U,
N5LWA+P7EXgNdcD@^_&T.@VYD0+Z;F)4&GcJZ-d=62;O4JRIPWQ&W:G^>)</3DO+
I@W77D7RCaWg[/G;5R3@_]K\W>VcbY#a9JIFTFM>LM9(52-J1+?RQI-0(Q//YF@J
48Qg8S-TKVcLED[I_ga1)HM..B>@9Y06[;3_:],_=6Y\OE0IeDV83>WY(S<-#Pe:
0ccRJ3L-QC_N/8Y-NTRcAYZ/IO1?S<LPZ5CKFH-Y,gd2HU-.S[-US_M9#[MKL7.[
6.6\72H\?T1GB-:O<A)a[cOfOSD<M>GV;DEfBVegN3U_aCf-0K8>Y2S=d97JIWX1
R)e=^N3/FVRO1M@X/AN<TfQ?3)W@PB.I<F&:SVI9)U;8;O3Ke\;1e2(L4VH3CTKd
WGIb>0K@EHV79&HSK=+-#Dd^f\P\dJODc/.^TY5U4F]0H<eH^f5GcGW,5bOW)g6>
@c2)JIHHR[UGP6)W1VgNP4[<Td1K(,b&b,f)<50I8>3;c^f)BD4Y3C1T>BZ)eb,e
I39[MJ@N]J+61Oc_,.,1?A\0QVEBcg6d?QYI\:>H1<(c@1-@.+.<Q/@+1R/=2^M>
1//E=)&aHfI,D57CO28KNMTE+GMe7G=QW5c.&Lc\=S=[3Rd=M54,#K/VY#\GU[;1
YeTEKe/65TW(0_BEA[bXN@89XK@Y04]A>F>Y3aUQ#&^a.:RMYJA9DZPL+fXI#.XG
]>J-dV#@G,U^&-EM00H=8ZO<fMCG<95Q;HOd90TP?(GSA2^4\;<^HgWBdUf62R?<
(1(DcK([&b#\^@\Ld<TY3c7YN^gEZXI[:3V;c]POP[:,U8Q,5<^PIT?@F)O]T=YK
A>7eeAAG:(MSYHEdMAYHGKJI5@8-b.G->=B46(3=E,2?7Z@K07bC<[;TFTG(f\L:
5@M9:0QX#?89O9,fg=Wa#[cRYXOIc^eMTS5c.DCg6VKEC/JWI)44.;=T;S?_ZF2d
3(b.37HVMU]1N]AfB>GN.PY=[P)+5e5=_I(1],AObA#\\&?d:<DTB&-eeDddU:;/
8Y)1[1)b:7R[@[>?e=/cAP]&CU^C=7/SY(:1JV-+LJ4GE,X>WCW:1U+,\TI)[U,_
?YR&V?@\S\J<W&PPE6^-IW;<A(B_#N&_EeO\IJ#g9L,O:a2DPA;K2U^IP8,UUJ&3
;QTXKB1@.(U)e+?F7SU;bR)?I.RXfQFSLJ83#[]daO)Cd,V?W=5-b./,ec2fB,^g
8,+LAP\+W\c-O;b/N2;+=@8<Mb[)UJIL/f7(a;Y#7HL)C_JbD;d3U#0M52Z#>#?\
&b:K+Zf58G]8+WFec0REGDOHQB1,_eN3_KC)5,H,9Q:Z<52g0;)BJ1dB.3#=^TRR
1O@\NfGPYF7GD=1B,W87:(JB@^g+B;1L+C4<dO(N-)fYKL#4P?]b8MJ(K_/>?;W^
G=3=(5(d<NdNHgf]1D(3SG7\_8-2=7-DL?b0cL,WZ0AC6fC4fXPb=VLX6)X1=)/U
+4Y>/QfLK1XEe1&d+82f)43R^=339eE<e:4Q/<eWK\ZP=bLHa-MU\/dd,V0<DQ(B
V.fI7H#W?AJ>U6X5@X#O0e1TY;=,M>QSJ(PEQ5G97a+&WLK3M8T55=H6M#4eZB[;
&Y^d^?0d&a,2<J(4.D,;;G-=><<ZIbJ(,T#X>S2#9LeSa3E,E,,KZMc#JOZe\P_,
b4<Z?=g.XN]&M/Z/&M8Y53VAf55O:Da=,)Y0a_\eV]E#,TaF>K->YD/7-NE<#V3;
gMCZQ\>>+)\P./fQ)9Z4Td?(_&[-R9GfO9TUFW]#+N>C02(N3aA6&F_RJX9f[@Na
\:/&H3N;TBGcC.KHSM]_1gX_W:gX[[Y:&f;+eJ_Y<F&VRR?K?SNVeOeXU5bE?WAe
[gIf^ZOU^5ZKeF9]\4PPg\f[LC:QXdPD=49<H[CePU,#7OF=8OY9gM?(De;SRX#;
HK1FDZ6d:OTd=[QOYL/aE74+4EPc_21E]YYWG:QPN16,=<#(aC[>b:XXf#b0M?+)
d\&]F<&cgJTQdf<WFA32b<e>Q5f5T[aAO>LXgQ^bR:AJ:#YK@##PC</b.NNg=ZM6
AG6;N\P&>;C2(+-,&6OEAMMef@6W)9YbO\9Q24XZCI,G;PRXg.IJIf23Q3ZE^O8Y
BK?\c&O#fWP1Z?<\Y,9@^gedbg?WO\QT<)?\M,9KTC@Sed.4]Q7#eR3BN_U4J0?K
90dTBecaWefF.[8FdKT.@VVPFI;E6-cINMK7E;1;S,ea5,bCXc6VQTY/eDEgbbb[
-KQ-)?,_L-PFV<=2MfdXZNJ@[FZfL#_edOZ0O1]FR>2Y2NQ993Ng3.+:g#Z8BH3g
2ebHIcKZ&OW0@-a[OXXRQDf@:SMgH[:6^\M6,T4,6b9I=I:G1^E.5G3[eQd#c?b,
F8<QYCF(&^P?_RQ8Q=[N/#B8/N7_4P<g<;c]Sa;YC0\/=_C7EB#gW&\BY@9#@AgP
WdaO=\R4fO4c_S8gGSBH?H?F5&gL>MY2Gb9<T]:d6+K1Z:-R6QO<3:)B-&X;O)NP
dQ7[#[+QISO:&d9?)3BD&aOL0R<G40H4e<M-I8VHc?X&KURT/@bFEF##E<]J]3(M
5]4->8@H^[ePg.g)<Q?:)?\a0aU[4/O[;,UAcDE2)EM1BTH]KP.(/#0ILQPS+2Q=
/Zg^KdI=G,a)S0W(.4.]=]B?#2SZ_5K=]MUeP\(_3,XfOa9,ZDVI^TYD>DMD:G#D
&\=??1/+[e2X=bWEZU\dMdd-g8WYWC[:SLc^/3=IE_M9D?Z._,L\_E<dUEgf_.TO
?b3(=eKFb<[Zf=T_f^D+-OF5A+5D604JW]^OaDK;c,B#JFKLcXc4Uc07(ZF\1[?9
UQ6[_:EV;[[fV2Vb?MTBW53HJU4OUVU\+5-NY^@=ROb561R035>S/,#/;N+S:G^g
NP[[=fAS84dU9G;JFACA^ga^9OTAbM=WK:D7We:/_gZAe8_Q8Q9Tb-Y5BX&cLd>b
3\XOZ.49K]BPF<:XS&9+ZZXUT=+,b6UM)VAa:4+NZOf<;VEZ#&D/ab.bX,-JCFGd
ST2cS,aYf,RTS+7bG&&eDPfW=eM+U_C&YH?LY--XPQF7N\2Z=GU^(6-__\:6C),H
OW(=2]&+7PGBI_:G0>)G=3U5R+48EaF?&ZZ,S)BK;cC2J@P+G<_<44YUOC>bY[V\
cGcEID-:6K8,Qf.[].RW3+36)0L02CG7]ZUCY_Q=TEA^#7<4\TMK.CGHO8)adHSG
CI[DRcRV&&UQT(V@PLgNVLWW<2QbTP#W9.^3]-L>[0_Z/_>JMJ[NNX63+(<4,NM2
Z):5,V;ZD2D3+=&SHYD6M0YD<,)]Ua;T;\a3:Q,G[Dc@f9V](YSU+8.6U5f@>&:>
88_6YEJ)7c.G\(GVe38)#0ML=Y<=TB:RJ81FcMF^+B>IJ3J(LIG<F<QE@C3G^@&U
V6UOMF)7]#/gW],Xe,L^RXIR^PC82+HN9:V/CITU0M?-Ia.4#-?g1H_)U1bPM:IR
EXbA9NFH\T4>V6dLI_\LV+-eC4gZgD(ZDEZQ](Jd_9.W>5CZf<A_E;1=E/4SW-E@
LBT5d&,0(C,@cR+Jg@?d9):eE7LAcO(ed[geU2g0CK=TaY3@T?U^@N-JZ9NcW[cM
_K1BK4TQe.M:T/f;_P1F/4\6Ua4J2GUR2=)=BZ5=eK^>1,/2=cJKL^_+AZaQ0VZR
S#^[DW^&-f.a9HGMEd2EB\B@K-<IXL72&B2PE&Z<;+Oa,NHeg[CEbJN\E36VHg#>
@GC6a16Z9+c?_QBeSWYZBMa8ZRM:_d^Hf(L3M3Q+/0=N^Cd#Lf^#7^U@/J.gOB]4
V;L=E,5(P\GJ)\9BM<DJ83/930Y3YBX.2R[W6IYSB/1U7MTD=SZfdZ(1KGK08NQE
1S:80I^bI\CEaC4KTQQ4._]R1W]E(E7A>Ab+5/L+=W5?-#DS7Lc)1D(/C.3:7_aP
\cbb\B[:T<O2Z6WMfagJc_0V-VV.AD13+(1A0&[BH>P;-Z9_TEE/<)4U:7J_@)AF
0Y7C?+T6CZ?BP4DaH6:3JE[FfbBK^cg?S#5f+D\f+d@KX7KV)S1eEF75#)A;Td>/
W4aa-^;KC?4C?<\&YI5dgbfA<;g=7()DD54+XOD]&LT,_1N8I^55YGcZ+.-@@PeA
>P>_ZaR5P-2)543WKdRQ3cI2b7;1O->ON)0XcH1J\Mg/^#W.@:c7)^3C^J-\V4Kb
6?3HY1cGWG2SYQBSSI32+HI)]>D:Ac\S[6@7[QJ_fJW-?V&0c?+/3:Z+K\7/[]M/
ZE-D9A^8Z;.SD32XMK2)d&XA<FA1T#^Re>>-F&OR)2\U^&8S;QVCW-2QR/NgL^AR
3Pd\^-FF7#.@[RC0fOBR+3,)a^7ZQ).(g0FBE>?#-,2c/MgcR1SF5:(SE/<Kd9XH
2K(BDA;>BG.MeC6(GaD+BH-UAcR,D)NdE]BTD]5:WZKRBP_B34Y?M<&a[0;RPUYb
#5CBJ>BcI1/#;(Lg20Md>J_3,-E.OfC>PEd;D_YZ9N8D-SDJ7)<eFIF4O58B8@OL
4YS9KJ..RI@>B2G@Gg;<Qb(;=ZCV@QbBUL_T/PVIRU]K4:6gOeXbY6SL(NTVPUZQ
X.2\8FCcCM>CXa>/Z^V7+]U=-2QMa6IWZf:eO<>BBgZQN:Q>_L6[>-g_.gD?8NO:
R8QR5O8T@68[26L/8=Db1=?d/W&&e##SfUf?G<M@C^G;d^L3D+AQ=IWdO_cC0E8D
bJ[4c\]cLFY^8#0.-^.37)cA=NfVHe_4:.<C::+U6fL/,72/Z>BbG6WVR?GE-^./
8J.@T?b\[9Y;]M1f?SD>]#IH]aG>=M[N^0=MIVY]WABOe;/EZ,YW<^QH?9;gX^(_
]00-E)+OXRN7X#RX0?RNZeH?CJ=ULO0@51a.372S1.>R=fDf.>Zf>g-;Vb@D9O4/
4e]1Z?eFA&]P2P,0I[W<e)R[-GbSS<\.7:VH7-32#Sb++2R=9V9523C?JCLUdg-1
)Aef>NYV&#?.@T]YCg[YI,1+&8bM(=#AT6HGa=b\WSHLJ)dKMRZ3QU]eeU1SS#Te
X/Q,ZYJ/X]M\HfWb:WT<71)V>)MDFMReCR/)MbI[b+NT#cK+.24U4N9YK/I-5?X1
AV/IG(;NR_9a,;2Xea/C\[]Og4Za_IbC&8I74^EV(Q2c@GSOS1PME,IJ1.JD@MPJ
4JR,V+9;d0^\11V8+SQ^[4MBR^,<L<5<C=W4S+U2aL[?BW_.\X:7??+Ka88[gIW>
IEb]Q[,Xf5?F1B/JgA1FPNcBd):O?1(:@K4C[N3X,JQJWG3NT>IYRSQ:?&)KI:)B
6DGAB(74;:fXDKAR]FfD2Y;8>Rg4cd46GXYK9=\>/7#4,>KE9FCVDH.TG8U6;(P/
K],a3@d&c5&2BGK2(+HeGSJK2S-1\Y,eDcQ)bXK+2[+7M8D36da<-,4HCg-T\KV-
@eS_-+fM04:g(16_3TF_BI\C^fQOD?PP5-;bS,4K1Z&PRFaH^TNUHePR#6P1^[\L
Ff41VT:Z8?XJU?dZ[,^=\_S5]RL>=AC@(f.:P/VM33d1KO]9LgX]GD=1MQIDY&?7
gD>]\;?9_8f:B)?Y_#N@Z4?L1aBO->WNCUBFM+WN1(M,2b1O_89[-RUNFc#,HdCA
B\=fWFJ)?(N,<.E,2G5R5<;]Y8XU3R&?[WOd;)JUN/9K^Q1VM5>a&15T,LTC(<:f
[O##3H_:A,2P@YX^bD(F(V\H#d+[LSaQ-G:dH0U@+=@Z</87T&XB\Ba/(J571dQN
S19XAR-X5KJ>#NC?,5;6?264g[d<^fdaFacZ^[WO7-H(ME.O934/Z+ebF);@(;8V
TWTXC:K-O=#HJbVV=.NN^cQX,-,BOQeJ)#>@gDSYX,&eCP9T0E=^5X2@0#>A,d&]
H2A&8N?P3Bc4\5eb^S1)OZObMeN[LE\F>g;F?78e4Q&eD$
`endprotected

`protected
NNA]#4Z1e2S;.A+8R)eXQ5UWL];2DUP3/SGfX_9We8W^[Ga7K&Vg/)/6,U03FD=_
,/>6dFLS/8YbR=6a_<B8Q_UW3$
`endprotected

//vcs_lic_vip_protect
  `protected
7gG(-_(c/658YDAI/4QAP&T1,:_#IE<fGS(-8^EBQT[>f)HI84gC7(\:\@gd1Y)O
9O,g&@9<0FT/@+6ePJ(-U^T,EKMdTXfLEAMU-OMJ/+dL:FH9TI;UfQ+c)GKfBREP
;X;dY>FAM)HM0W<Q\)M8.aT#H.W4&8#Zd[/X?1]#ZDb8/S;AR#[>DdB82P^WCC5T
Q4K5QLYD9C4;d_#X9S40YUeO3eV11:ADDEW#D)/c1KD9/(1>WTT(dI._ac_=2g\W
&cd0]UB[0S>P5]Kf3FCYQ5X(g]_,.)R6(R(+@KEL8:f:fdZ?GG^W5=g/_[8ON^>Z
<6<CZAI)7b6HO:ABc/OC-NeLf_(;;1)E.,2Y4Z;(Y/XX96^>)5U[I1EQ>5[\^S#A
<5C:-VI:7AE3LHB:[+c>J6PfSU-@RUPbXH7)EA;TR?0?O_E2JF0AZT&-FYJ=)>QE
:BZ6;L>cfH?4#NQ8g@dXHbYDTS-</JK)XR/HP-4VCD^HQG4\[dXUF3)deJ9(0#HN
P(3H.,a[[KX2.;g,3A3^DMf#)Q=.DJ3=ec>F7ce3KNTe6\_@;bW[d3b(a(0R2bA]
NcCC8M;QV3U5cUXBHPHA?dd&I,[OdD&;U1L_#0OFBNgX6N7]c)QeI&c=Ma&FD/)4
14--6^>4+_.313g?5;e^-cQWP(/ML26(GLE+AOfIEOaC]Gg(<6ZJZe;BLCF+^B_?
ZTF<Y:=SP[&Q:2SEOd9>,4@ba#f1?D2NIS0fCD:MIVB4O/3LD@8D(Ygf)-Y(+8^;
=dH>3-C;\X+?9P1_LKPZPNVTV:-c6J0gM5+)E[7&B/gZ13dBPXRR.^PJ=K)XT;O(
cG@F9C\XQH6-V&^?JOXUBHd=2+XBX.&f<G=A-W=(JUMN=;+QYOAVQN\/Z3RffA:[
GAINdA^+Gc76.JeH1I=@F=5L:d(BU?V\b<4UU[VB?T=gINWP_#a<-9_W7A/-_:Fc
,F]dd_=O06R_+K\f+GGd8D3,-;1XB#-A1dFV#MNI6?T\+]DE4B_I5eR7SA3=Fed@
VQ7I[HeN<6+L_F;.X[]cD@YCW=3,-15L22G-\N&_dfJG&.^,:GBM#[#g6(^bRC]<
OOH^X/U6G;@\/U_c&M<FOa[1.E/51UO,/>2BNX5)B\b;?T>M8[Zd_XQ@0B^+T>FW
^/eg&KaO?C>^aZ)N_dE=<)ZN4-4(=e#>]X]OG,MVCO+?.AATY>-gD\(C>ASPOa3F
L0^f@cC,G8&>97F,\059G/OQ#YM/&/\]^>79W4?600_]9C?<eM_NJ1Z6B1IJ\B(.
?OZ[,cON=]09UV1LY#H<>J\3\@&/.M0g2;7PQ_RZCYBI+=XZ(eS0Nb(\1CbfCZKR
d(O28O.XPGZdd6Lg^-M=P7@DK\ee10=eE9XeL8b&D3YHTP)Me+0A^A;H(.>[YG(K
?;T[5C(3+R\1b4bY2WcW>7]bC;-VA^cg7H@g?=#6N3;6;f-<ML\2_bR:N.,1Y^]1
@T3H.,e[62ARV;c8S38#XE4VM8;XQKb)2gJXPNYQ]-W:?3-G].D,DY=NYI-^H0?A
(3a]Z4eg6+0<&?>A9\V)2BMS+f<&1Z[/HZ9dF^;=X7=.0=]O]NEDBG)Xb\g>afeO
:Ze-;S].=aSZaPf1UUY@&(7?Y=KK91<+-?7G)2A@)FAT?)#9a)I/<=aU89Y/AMSH
dOfJXY2<E74f9K2+=MXW3BJ@+WBG?N/5(R=g(,abc;-2?,&KBgRO5G?b;+DMW>/0
:H&8C99CC4SU:@a;ZZXC@\8c:_O:Y4ZFZ72a#4JfH_?TEBC>a]PTE>PH+gVGC<7V
&CJ^a2L2N6eI.(g6ad(3RXQIObf1MNZZNBJ9:E)L,_6=OI^c+^,1FX6bHL>F^04Q
5:W31_<5YQCG@D<a<I@?J,7X0#Z0@5FY&M<R)bR4XVAXBXKH8U,)F(:Z+3_97&_@
\QEJ#FTGKD4N,R\[2)VHU@E7^fg<D1#XXf+Q-\ZGbQQZ><XeFS00F#H):@;98T,V
0=;FITReT.PTYRb)\c0^?K+G=YJ+)a^#-:J#HfOIfXSOPUIMC6XR2d6CAE53M-c?
@^U<>bZ)Tb:T/8R:P:c#1b+BOE]g0?:[#@F^be;3\F2,X<\6ecJ9BAg7I=@:GaY&
4U6>P/\7V#G>=9?<(\ASG&#CS)2QFN:AL#P7UY]fDTQOH)E8(gKf^EWCC\0;35L+
feRQ-DU>Gf.R8>&;9\bMWg,d/-0KWS;ZN_I9HPUU)Ob=9FE4G>UX6W.D24_7P)1H
1e<I/,gS7KgAbcN&S[=(-aKS;.cgQeKW_/0);bI0AI3<F1B^#0(:\[d:^0@OYP:X
#5OQC2&/K/KN9SR9Id&b3aY8/[O(aC7^4,EBN>a7.=3?^4V:G8Kc)2)-65S\bSIB
-6Z08,W]@ac(F@HH90IR;TTA2f3OM3ZT.Rf&R8T+P8c\[Xd[@W+OPQSR>3U\D=fF
5Hb-HX:E)DZ1)aBS.e#LOYW]TP9)#D;ed<P.-G5:1Vbc0^2E#ZD^^7[0gJaY9fN0
CE2]3J2-LYOVOCE\@Zd-M<c?W8V6+9Jb+a.^_=[71:V(c&,M9)@c_RX8(8=g1I+2
Q8g]UE;\4_(8^cQ^I7]b+8;bH\U[<G0gPfICN99X/?N8_GASDae3cddYSPIGOZ;9
3E+<X013F-76.UP6HOcQGC0d(ITRgA+[F>I;_CBZ-I+YcV>WY6L)2+56G].HW<-4
Z./]\a[[A3S\KK&OHPCR)0D&61,(JEZ5@D.YYHWWc8^Ee_U&0T4#>85>]C7@g:B0
/f?O\G?=8bAYQR#[WG)c[EPeGF/a,:EB5:J4[P-L[ROHE1U;RZ=X)]b]/4ZY;4ED
_4C#M=-Dg&0Z^]+3-P?FTeY@Y&?2XLI?FNTC95\0<SP2(QY@I=X@[e]SM^.b-043
b9FI9b;].I<L8#+e40Z+S>=7+Eb1V&^C0.A/?+G4AMQH0I6R&AWfG+DW>aW5B28S
P5,T1SF,NK(<_0O/Z;8d9[JR&P6WC:CIeO]1S+?)g)5B\JQdA4Wg4A+E&-&PV8@K
1VI=GAQM2=(ad\_K5SfT[UHdKgN.QPI8WU5=SJA22e)&HPAY8c)FXc6\^[#bIaTJ
:,(gOT^GII5DY>J[D@Q\TTCJa>K\R4GLf3QL^9GK-R.Yb/.-QQA/L=UZTYL=MFfF
;MbNYJaF#\JAQJ]/NG+=QM&VJ)-Z5Hg-OH]5ddN5DF)dV15IRREU>3OE=/d4YMHI
SH2cPbLa)7+A9T05JXQ28[@]@NK+^&)5acA^[QI8OAKg,-FG;D0P(M4Wg9CEN1KC
bEJU3HPESD1ea5XL==KN935cA8<Y0g-1U^^HDSFQW<28>Ra9PH;18-abDU_]GTS;
<=0bg]#-P-UEINQdDg#Ue;J_DXQ3A)+6CD7TeaNHENdJD<]82H+D1P1/)2;,c(A>
Dg6:+^cc5OGB.W5Rg==8KIIH):H7;:RKaX_@>Q;D>--ddAg8,X&ccbO>d3g4eJPd
@39]#\Qeeb?XR+9UT_O)P.cW-V.V#O+A3OJTLf:_VNSBV<(J=DBEJ-5\,#G6J\A_
_\47.d18TX>G#N1]NGOFKaE?+#a<6QBN(Nf.e_)\;F]0HUPFPRVR-[3TIa_863Nd
TKT^3F\<g>+g2,+]g0;->.(Ge6R8P#aZb<aXIbc?V)K>,6Y9&Ng>bV-f.H:e#575
K1<//DT-PJ9KfOY655aCc2I,,Yd7HK/P@cZd>@1EB]D/Q+HK]@a8^+^V@/QE>4JT
J78^HafX+Vf=fAUNZLZO635cgYSgF86GAe_RQM+U12=-16WC9BS,F<#-NCgMJ[;&
;0M.7d^^U9d/?^e(]8YP)g3AJ1M]TSf\W.4,]c6I0N-Pg/@[,Yf>KL7+6RVRQ/J&
MF/;XGaa1#7Z58;])/7JY]Vc+-g,<Z[e\6?_g93SEHM4+X^C32&N@998fX>45NR6
#7+1&&2D)Z\@8]XV?^/g/)-W)K>ac\(6aCd]RPcD@&JMQG9>2,_V,_Xe#R0d=+N@
&<:F9IO7/;@g/\g:IO]KW7Q:d@;aP5NZA+1:8;)7e;_/JIb]4+Y?&_&^+-4(LI2=
7Z1L8\NEN1F3b,98P+P?eA^a6T:@DY7SRJAS#]^]MK1/W+XA#NaRAMJ]aZ4_[&)@
A;9JXASM>dT0=?/e4[(_Cb)=<,6/LNSbMcP/<eB9.Ebb,S\YO[GE77,4&1RWX\JR
R47R/f)N,cG?>RbI?:5=F2cA=E=Z[<0Pe96:A82e+.DUAcc^Zd.WD+#>HSN,db6=
2M+;dcDBUeHV:+CWPPdQ+K2]f@Y<d+HT9>T\\c@KaUe?)X:QT)DJQPRARUJ#UMMb
7M;O[LZZ)f-77<?2OWUg<aYM-@+J71,1H[5Za@S+^C+V]A;ET^.H_aSb7EVI:C:R
L&#f1C?04NX]>+Td_35bDC/cegJdHFH0Q:ad=Qda55\=]HGS:cP.447D)4Q^a9[G
30R&2I:BDO3/5=@#5G.BP3a1_9/_Y#WQX\PK1Q@=[LVREdGXEJ#O?VR+?C96a4HS
=bSX=00]K3.)24f16;-)-WK9),0[7,7R02K3ALAd#OccdFbJ(0Q6:D8@aD/\6\H(
QDYZE)7Y^1(fVW:ND3@,L_=/VSU>P4+11Z:gWPBO2P629@O,Y@DIIS+OB)@I:<1L
IMVPVBSKb29V2JQ022aJ_X#b#bZ(_911X+Y2WH(96ca=5<H47]C+SET>6MfeO4UZ
+eX+6fd=/M?CWBJGZ)4S_NXdY](FE^I-#,)Pe+ddd@GY/.UZYGcCE>0&H4GJg85U
+8gY-K1LBXV]^aZS5a9JeWf8PL?#A)BCgfWG9b?^E3F]R0=2cQSCBOX7C81]P:Wb
V6=Z7J&,d1J+\SCfK]S.AbELbVCUPS1<L#IgU./SOU<+Q<E/L)?;H,G(I_=JId.F
gVD\,Y2@>EV>B#1(3?\KZ:#dD)NA@@MJTM;K_Ra6Na_\RP.agI1X>eOE6VXC4.Ha
6PbBa+V,JEM?d^Q]+WJ+_M8X&NTLIZYgR7JZA\0#B8Q5_8ZK(5#@QMI_DW&_[<F,
(F/5QP?-+MgZXA(V&7N<1]1]EIQH5R^7JGO6CdY25GQ\6-@b6.XC,MAO.#D:GgbF
=_#0;?VP>DfEc/Y<FI=E8[\3Xa;VBe.8BBM6G0G8CNd<N5#RR)I/3+L6M/?<6M(c
[V2-\82A68RW+CU>+\_,(UfRYRcSR(=fdWW#Nf[&KZ,T<S3>[?84)c</&Zfc.XLa
Lf:FX-U]fNO0Q_6,fST.3RVMGUbI]MG708e6aBdB9RV8A6dOa1GY.\PM#O@3W/0:
3D)[:Yc<.^[8M,.&[K_HM>aC51.;S7SC5c<NB&XD.F@V)X.-(^5IE3Z-G66D(L1E
>4FF:C<:W,9f]^d:a8L4Q3_\#<GE#c-+A2.C9#CCV-[K8OR2)Y@H1a=VR)LTO48H
a3=8>H;:LgbZ;[S:3T4AEK;8IVZg/^-U_fNY[ER-0(?B6,#.7fe5H(@fGPMT_a)W
QXdX_b_/-;d3PKJ8OG\4#[FXASQV35,ZM>IAH7J8T846F[XR1I3edbET/JIfB)5&
;XOU]cFT?\S7Af(_FfdB5D7^:YcbYUd.a;ScULJ\/QY4:VJ=54[)>2UI/Z7J^=S_
#99Bc7UCbU+IGVgP+F=5C8M^:5d,XAeA+ZSUb/41BG3Q<^Z<]>0b4Pa5=>]:=QM;
[->=)IJ5Z(HW79B#PeLeK,a5aG8MV9+2VA>,aK(KVW79^b43]\B)U_CU^B__.@HD
:gddd6eE\X#V(B[X]T5EIfS3.O?_OO>L3TLQeBS0VE-B<eD2cUA_U@U&MRaG11<<
2ZT=.aE<JL,[XY8V+.0U-LUP^4a(8fL_I<,D]C7E@#AOb@1#,PE;8>FZA\CYL3#a
#9#e9&LT7VV/^^LEDdW+EMe^&fLF-Yc<0C68b7#>.@7W]b1E>ZM/:X#9<W5>\>(@
d]MB.Lac?UJWEaANCF>AQV^W[U3?g4P8G^cUZfY_A+f(C30G.DbcA=,\bB?gL4R[
E3d9&:b+X01g1;29I8?Q/:>-d4Xa&D7Q97(fSKRgQ6#3_,6..U>N892X#]W@1QX1
#eNHC,H8Y6=OPRPZZ<C6\DJ&f4#;?#4=?RdN1OWG<A(SbcW20P\U]?\#D[K<;)T^
I<O3U:#XIS:fEOb>V8Tc16XZ_DJI;3C&8K.S--T>K][?5Q/>&I7ICOZ(-BVRM5H/
9BG336E?1C)\>G+/L1aJYRDXS49U\,H34CH+F7Y/>\9NJ1bBF@&1V/;Q]PDQK6O=
.Y<:3Pf,V>>OC&8f:3>)NKf,Y_U-4VHfAY[f#48^Dd);d[L(D/)#+IM_ZHb:?EQL
a7f(6?Y:Le40HG7-6<1eYa;(#UM:-^;48+[S.^8QFggVCF-4d6MQ5CI-=d]+/5B&
EFVJg^N>34c\A6(V^<EY8;[O(B_N6Z)2=;4aL82.Yf._UIHdLQNbZa(;_035-RV.
b_Ma>2OQHCJ\WKfA404ZIJ8S:+/,QZ9ZVI.FSL>7#L)G@UC-.D5I^^A;97_@AO_2
(9Wa[:ZM@5@PEfO4Q09HZFdAIM(B(_-UWFcLJQN9<CS[2e,^]B7,ABK64FRWG^MV
5IZ1=(DeE.9#9A76@Lb2&1f+K(A??QWGf-:f;5L;g<EEW;DZ,8=>:HPW0F16(AYE
0G(,.2I6WHJb^A=[PBMDP=@bVW;.>NZG;JSD/e+cIH.-GN/6WNUa8NAJO38;RRfE
>XC4#>Z7X5N8=HOG>4Kc.bf3+XdJN;[8f0)Y^7b0(P3e5gZ1Rb2GC;@Y^ZJOHGUd
UZ_0Z049F(5C.e5NZN+f<JXMd09[BKC,a.4GH;TQZ9f_F9[#B;O?_a-R_?,>ab6+
W1JS>dNEY2PJVJ=,M;gQe#AdUbK.T+;=8,]g:&L#TH0ER^\\LPOR3K3cG+R@&)L/
V67:aACQ6&^<#KLZE(F?:T\f;Lb?TR-_dTZfb&DJK8E;Xb<[.;b\Y1/f+M/(g&e>
c+;ISQacVC,dYb47CJOOQC-I9@^+8MJ?BR@/;]6E(?O>.64Ma):-R>-EG2f(\X1=
g)W,1,K38[4<Y88gQ995Y?@&:2XHWNZb.a1KCgS<fV<P,YdN85VG^,BdEUQ16=-5
bNX(eXL5JC?.K=KS#@^=+#,<5bU>N0Le\eL7DFHD3ec\c]4_4<IR4)7=W<OPFc0(
LS.0K.ON#U:7>b8ZYM>FZ<=ATPMW8U(^d5gfR?g#gCg:IBQGcOD3&9J=HOID;dKI
g]]a9H1\16[QIT,;,=E.?9=#3:\bdY6eS/C0UNg2HeL+IdHJFMBWHNMFUeEJLI6W
fV^J]_8/Eedc1?X,GdN:IAYY-)/aMPS\FI^M^AMe,_[M:gH=Xa//L<B=]<NX=7O9
)EKa.;Gcc@^f0UD.TX:0I-a@HeVeb4S(,)XP</W<g.<>fSK3Z5Y,W/aG,5V8aE]D
f3)7;bK9D5e#SRQ8[b5OY_faC&]5&=&W,Q8UE+\[33/ZDF6eH.G28P28f9d1@JFB
PM5=T/_N/_;J@_Y?4<4EbX]EK^Tg95Zc)(Y4=DXA35,aU(2<9JY++.-/LX)GR.R^
SRS01L(;Z,Z/5/XE-D=L^\;9Zg\6T_SYUL\\7G7Geb_e>gK6eD:)E9IVM)4cZMGR
2ZLKg(Z6S6cf/(2<7(1SEVE@CO&MP]S?bXTM1gHNF,MT<a_H5/Y3d-?7[?/MHT@/
ZIgbT&K#-JQI^T#@=)^D)ZE9Fg:9/Og^&=.C?gAJ)#Z3gBC6+K/.D7fbG4PBYU:g
(</TE#KRWd2]V[O(6INQI<fA2-Sa@FHdIZO\cS;D+M)9L?<\X[:_Zfa)W4M&345U
XW(Ie.SE@C,YEHCG)c7f19C97(SDS^VZ4Wg0Q)V^3BI[6FS55KO&C^)HJ[\8F9=>
Zg6cPC2-@]:4?C=c-#H&K\Tge?XXC@fI)b?D/C<SY4e,fKZ&9KL+_?]<d\QCZKO[
&_&<+SO7(F@T4KNg,YO/;(C12K]_f@E=?8LRF_ICcfBS2]Jb?90<caKVOE,V6J^.
8e7^SUIL=0F(E^9/VfO[7d^E;Y]68a?;cG/;[Q)TA&=UdR,aDS56?7AA-aMgD=<Z
eIdY3<F61e&@Ne&#.e9@P)abPg3/[R4:0M-90Y3MDT+gcfYS8;UQH6>:C=3,f<fP
>4a#)WY_]LGEJ8B0fA>_@^D9<_O=3XTK9M:X2_()UbC99&@WJKW#gWL&[3(09SdU
fWD9^C8GZMBd2_C43O7a[2;^(REDZJLQfA?,L]FgJYdXbIM0MSF2T,9&6,@Y<\.R
\U#Q@^>;2Q2#,c=O[aQ1-,1&0NY]8,HB7O8fg[^B??bSe,>E=C2A^JAVe(8M<\5Z
=(OJQ&E6(2H4J0AIB+bS1NC_HG-dY0(?Za)U-=O:d:EUO2F0S_RCNDM,#R1^]/Ib
3I:UM8>[bQH.=7-90[C6:YZ&:BK@g?_a/F3D6HVO64f)P=/]-5a8061SZ17cHeM1
&L]P26_9]7]@(S8g=:@&X&NUC981HcOULcV?G:H1@,+#fZ+L9c5cOeSJ/C+M=0.&
(3HKBCeN@I6.&W\<4Z,bNSID3a6\\]./CScS9&gW<S4;J]^-@JZS,&a#@,\1=+^6
g^5JAJ@f=cW4:D<6&cAB=?O>3NN;L:gU4;TA?AN5feb)Pa2)NbBbd6-_>f7?P<6[
(Q;\<>&I\BR184b^M)5V4E3[eFKPDb4Y:DF?C)>V[d9L:A4X;EL:Hf67OMg<Me^\
J0eYPHJI7ZK9OII13K33S=Eec[)\[0\8WKZ.@::6Q8]g;DB:f156<I@XUC;(eHI-
=9RAR+@SG&\#6W(f#1XKH=2+<4c5C_N20gbbTFSE_d@W5@f=^S4B3I\_E>AF4fb[
Nfb.gV>#Ddf-A?S(#K)Yb2PW@#72@#1Ca+APAM3,BA])]543d1CMN078CY^F.dJa
\=]+L:Z>?V.0#GX<SbbST)=9P43@[.(7SCU-df/VYIZeT(\K.H<c&b.g<,Jf>NC7
f<aL<7I5-)AY>=(/+dbC)9Ngd9.,RV\aTW;KcU>48M39H2QD:EH_QDUgX#D_M&S)
(GT(U>VG=aFgg\?-E/?gG9HD:Z.A54bIV2=.I1V79>N9&ZV)=[1F12,YAQF>OPg7
XgPQ7#W?HD]O39@-@71#X4+_f#3/;5K&)XK#aD_-R8_L:eZC9&5Z63-4e\HW1],)
0\O,dDHRS60e.d8;.^K_d^\#UcZ@)QMg5HB<1AJGQVJR4QG5fY.RgMQ^f9a(L,R+
THAF:ES2fVO7R#..Q0<Y-C@a,Q,bHFHU:.UP\[CT7g(OO08VO;7++CJcdFR,^378
0@,Ed^\/O4VEAXLHAOU)Y^#SfV52Z:_,#O15dF+((]OXC:]WZ&(B78IBM_gH6I1(
O=ED[08[B?EU^M3aQDMITQ3I4MCHcL//[^P34Y0IMMLd^-)B_RLGMEGPPN@ONDfc
@4KX#cB)L47aG=DfV]WcO8XIX<D:9)MR.?K0e<9G-bd_ET?g1/gd7+bgYbXeMSbG
)UWQ=Y;dTYTIdZdD5?X46c,A3bIW3SD=K,/eN#ANGH:\?=,(R6Y/Y3MWf(:>;PWK
T3Q,.Z26OLDEIUfL#WRc50J)PIF=]=:MS,_<IQFgaB<@C=2CJ7G8<;<ZG)T1Yg]9
&D7#^I;3^)8+e-6A,]_>UVI,WALHM?Y2GBGZ:[Z&PEF36cdQ3da=fFY#O(NBW++_
He^B-?5V5M:LV9QeUCaU:,1eG@dINO0K1EX\eAfS.aI^NcHYT_N<2=#V&=\(>(+:
H[X0FK,20)Rc?^5gL;=)H(\8_S1Se^N\QZH#<WTO_:-_-BDGf=PeeT5U]O)+PJ4H
BN.gKJ?\8aN8EJfUW_0DWH_6X2IYOUU:[HdGK,#J,VKMgE\VHT>NGRAd[I-Vc1+2
c(b1C,:RadI,AN_UfW8K<4)J&?cYIU\,S,a[I6QA:eXF&(FG,YPIIN;E?<:2b&Q3
[3NNX,Xb=:[.FP4<7Q]KbN+<4PZ1\0<^EIA9<QdL(O#HN^=-PJ268b6Oa\(f:L7/
1?S_NXDJ?[-4:^-?\<81JT/9J12.W&&F^25V7,=NBWY=LE_H;J0]0aBFAT.9?9-1
7?7XQ7>gJ@_6DO[+-AHVWW3ggRD,.H\cRIE^;41OT_>]<F;-;1_DC:LGDX\6VN6+
4VV729GGHXA(#:>2aT7<3b5VF,]VM8\f/NBSU2IX-R.#G@Fb?cQ..C?U1UU/ZF5&
JXXS_cA)AKHBUA;RY-B&?2cf\cf<0dJKd4_\5=gg2CT6=P[B;@IbT]R)-5AQ)XU4
MCF)9SS1HRREBG>IT^4\]a>):H,@#1(V:SSV/>6/-)XBWQW+],I#2&X+Vg;_JT-#
QFNaT^1\9TcL/)\=#+H6Z@3V;fWEW6\>Pb+aSU@:9NLKOc0g@FQI6:4fY).=H6c+
78JIK?>OX<6L5_1KGX,TQN[3HHS7fgX[T^,6ac7-Dc8(83P[.\e+IdVeN0._8AU9
:<&BTf\9C3gHSC:gBVLKT=PDU\g?-Q00D^W)C]+F,Z6Y-R&]&LFC]eU@D,&3Af^;
a75YWNM]-XdJ<GD775\D1<A6]Xe@Q14b<]V.0=565_BPOR:6ILS?Q#U_,M>>.f)7
R)0:@WE(9US(d;LJJ_.f[3W-XVHDTL-4Z9b?B4=SSXd?AGQJPI;1;+6UP&JJ6OEX
93_6G>1\1/=.EZHXf;KC=-0(]_>8&#Ng^Nae(Hd.,e-M=60Z)C7,]fDU]+6af(D?
b4.-[49)YXY:V/\+WfXP)#O[ZYUXV7=-OJO@.MKJWRe=4[>QW_dFYWa/bZ?4<NbX
a-93N6<=N6f83;T@NA:_O:Qg:GN25bbT9T^U&3_^]C0.4+7-RK:MWWRTQd:Q9e;U
P.:8:&#[,B0>,c<TU4V+KT,aa:Q7HMdE7GF4N)_-1c0S,]QH<B;KXUS0#?,(fdaN
FB>CI(/:R#I7WSL])/\Td?3^W0;XIGa2CK,7cPR_,M14c@M[GPU?MR07;HNIC>E2
PYXGHAZ?8[-P2>+TA50LcX6>#,@.(cR7<<NNTTOBA4J0^;c[d(/M)ZCTcEXM1MU[
#N4;BbWHacXa=V6DB5L)L/H-7GMeH(Y5ZRV[IaNR&5C9>d\g6_b&L.+ZbgBC;(C)
88+&C83V&,cZ#<c^;FFT=]J5^GKR,^L_4>=7-&E#=[Y@aSE6..CaV66..](SI&SZ
^C0S]3XHbL;K<:0GL^MaU2IX;)Yg1[<[G^(MXd.1P#-&[Rg6NY9C:e;fDPWBcY8?
:_X/E=M28#CV7L02_fM3\WJ[+;0M<K1_d=[7?]N:XV5\RcP05E4.bf,>?MRZ.HL?
G.1GbVf2Y\3<9bdZG,bWK[MQ8OLPBLWB?KW^1)H?N]cdg4a3,\NOCbe_UMRRYN=]
,HJ>?aa<E0WP&@<=PU/?AZX4A,e.7<9ZV;JN>\V4B0#?GP.a,6GML+BER+g6G0HH
KgE/+4.S2B1Q?R9J^Q167U2@f.^dC7_e2ZB8:NBM<#]\77&eQ^TG8X993787XK_]
4E;)KXK7C:S=<@gCO3ccKWH?H?I[_BU2Yb69aK0WN[8&IE0dHb-P_5_087a@aS5f
f)OD;aX9S@P[0:.?K[EFd3c-G;bHdbN?bWV<?@d9@+Ad90c@eTdP?0+VML;>J4EN
TH@1SI+PN@5DcefYY[_EHH+AUIWd:Wea(<WX-F=P(2=M)QR?&&2TO&OB9YD8F^(B
3?54.,SPG3,?]GI:(DE(XGVPK\AOLDZ0RLf(Qg3R<I-<NR^/-#[ZC5V/cefBcJMY
c0-P35bB471:.)DMff6bI0:Xag-?8&c#aO=,8a0P]eQ&[]QF?#)0]]O@Z(:IFII?
JR9&Xb(ZE5@8fEfMG5S^AMM(Ya&-P+Fbf<aQ17=gR>cSC\\D;+Z\T3DQ^6M3(I#6
&9<1E)DR?A,QVDO@UU#J8fV&bOPT30,bFUY?FPT4NA]X)H(\(=00=HD\O+(G.;KK
+CG87feJ.IO\GR_e)\G[?g>dXCDBC;[V5T?NELK;dF?VA<9T,.VP?b98?0f&&aPb
O/(NO_KPN[:=9dP[L16H_b<LC@>;_<7g#eMA]E&A#?JPN?.T^8,P?T:OE8#f:\#,
E>9T=/D\#4>bg&F]=8-MC,(_KB3H/A>#8;4X3>cCVQRVTB9?GR@88FN5Z@=BLSOZ
Y(?#HG\e.gWCA-PSA5=BcfRaLMQ4V6f?Nc-S8EX.cF\4/A0Y@<c4JFB5_=40)<LX
[Me]0EcZ<N<>Yc0W=N29U&HJ]E;.#+]\NQPYN]YA?6_]CbG&^:T(/K2FVK?(0Vg<
6\=We=LSDYf+[LDJ0K/QC:K8YM<&/4E8#&L>MI+7C33aRIG?/.M0fPfOY<dHMbP@
DB\;WY;DK=Q2cS>US=/\eMSJ\5,gd5P=H0=0=O8K=UE57EB>83CQ49TLWS)K;PIS
9TE72;d-,QRI59TQ>[2Y;GUH#YV?(d7_+2X\H^N50VD^33,b6&CBQA/Qa5e(_f1(
eg_Mbc3H7U,I<@0(MNeHQ2U>^GH.(>O#SV(<<De+I]7<>=922O+eNJ>@b6XeE2=W
IO#f/HdJQ#He23._b\A3[LNYAN:2&YW_:EMP7g]>Md@6a2@?V29KUKB]4=-]RN/e
K[ebH&[_:3JX+>8P3S.M+J><8=ZKZWQ<GY1T(f9\RLZ)\IY=YVLO/Y#:,IR.6#ME
RbBRX2aP&;IRRGC2D.#R=^1<80:=LZJ^@fG;W2Y<?4;T#@.)>EGJC<I5@Xd2E7Of
NebWe=65)N+,Y46FOAG/IBKK#Z.UTBY_GaRE[1+E=c+,K/COPD^COd+5JE/13aJ3
38OBEQOeR0ESQ[;2=W=Gd2&\0dCZeDZbH_XZ\-A\\,OCLdcR.d@]b\U)?AIV(\_3
QGJZW@LDO-1bdRFPYV/)#387aFK7M1@VL#:(O&<R<c+/P?A)]TH#R[^VbUI2?R+3
9L0^WEO>F=I1T>.Bg,S1R=0FeS?2CLN[GeILR2WaMUAGEBAZ>I;fdQQG.H4g;Q0a
=DEdX:(fQGL)XS4:B.ERXa/a.7>=F;-bNQ4eN:ZTfQg/ONg6[?I[9;Z<c]fgg,C:
2[@QUW^1>Q^N69daJddY0;+e&^3Bg7b?eCN<?2-.WM\3<M64fE8@7d+T](F@KJ^O
T7aDf/)CD^#DVL>QVfI6b>f>B^cG<P\d83_Y4F6?gYN,BI-E9EEA8W69UE<\0:6B
)c3W\_Y\gIHG.P=HO6g/NX)#:<BBKH/IL6L3VBJ+4ICb3?a0YJ7,-.FS5WN9/P<f
]80CT3IJFL\-#B3_Q74VWLUHSO2;=UY]]D+Y0FT7c>7>DHM86Nd7;aAfX.;E^:dJ
Nb>J,9\+#AKC=8>+;03J5fH)gYVPF/)8A-T[6ML1b:1_;a<6#+cT,;&bV3W#7<:Q
1Z_7[ZU72)YB\4GUOXR7+f8b93;U^K]/e,WI8OZI]]DI+,@f9,eQ#2Z[(&d/(_9,
..C&=fKaG<[6NH^/.2M+6K[B<fd/>)/LIKD/6+Sb9DgUC&:aX2>_<LU[VVD/.>HO
ERf[Beg[&V&L>P137:-I;H6-bZ,5K?1LKLO8&e[fX<.1(<T+K[)1,Ya:ALY^W[YJ
(]<5PP62N8VL];]:X<C+=<[a;?]4H.F,7B24_=OfQ?3^<=-cLGF&a(>TPb]0XdcE
)TXX//SJ(S5I<e#LFGNCc[QSNEIM>[=NN=2UQVQ#geD;a&bYdCN60I[C-cP0_Jg\
7<\HSG:d/^_QF;f)2UbC7NP?DGTN=)G;U3S;5>0(SXa,N=<G,Q5[/Z_FEG64)_\8
8^W]4Q4TJ<>b/7OS785X#VA71VFI2D?HSR<L/L75F_;Z1VM)Fb(HfFU/CCL6-XHW
0L(YK;W3.86:,R[BAJTPg;@:UL:eeT4P#XPG523Kd,g@Oc(GeYZ],BP-;NYSNTZf
NR0GTJaX>=<EOSH?)I\W6SbXN7g5BH-gC\Nac+B7PN3368/RaUKbCDca]GUZ+4b0
)7HFWB2H5I[A>E3d3bB]cBGf5Y@#=C@I7)#-5DWP7?6_51W;4?570bX1BD,4+g7Q
7@c\]X/+=F=d)g#cU<=8g#\./OeAbL=:#?;/A0KPFUT=-B/gEe_fF#3d=;(<f5+V
^C>a-=eHR1/M+/PCDOP\F_f118IPVFJTGW62O9M7K0E,>8)//Gc^2JW3C-92WG)(
UH+7NT#).,ZL?SQ_V7,+D]OZ3?_1(?P[T\bUD^5L?:])JgLT<.GWVFWJ15-b)eR?
LUC4F8PegJRTBcDGM09N=dfXA-dFQ\_,<6]1a?KRaW>>XWX5D3]OfZWJL$
`endprotected


`endif // GUARD_SVT_AXI_SLAVE_UVM_SV

