
`ifdef CCI400_CHECKS_ENABLED

`ifndef GUARD_SVT_AXI_CCI400_VIP_CFG_SV
`define GUARD_SVT_AXI_CCI400_VIP_CFG_SV

//`include "svt_axi_defines.svi"
`include "svt_axi_cci400_vip_defines.svi"

/**
    System configuration class contains configuration information which is
    applicable across the entire AXI system. User can specify the system level
    configuration parameters through this class. User needs to provide the
    system configuration to the system subenv from the environment or the
    testcase. The system configuration mainly specifies: 
    - number of master & slave components in the system component
    - port configurations for master and slave components
    - virtual top level AXI interface 
    - address map 
    - timeout values
    .
 
  */
class svt_axi_cci400_vip_cfg extends svt_configuration;

`ifndef __SVDOC__
  typedef virtual svt_axi_cci400_config_if AXI_CCI400_CFG_IF;
`ifdef SVT_AXI_SVC_SINGLE_INTERFACE
  typedef virtual svt_axi_port_if        AXI_MASTER_IF;
  typedef virtual svt_axi_port_if        AXI_SLAVE_IF;
`else
  typedef virtual svt_axi_master_if        AXI_MASTER_IF;
  typedef virtual svt_axi_slave_if         AXI_SLAVE_IF;
`endif
`endif

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************


  // ****************************************************************************
  // Public Data
  // ****************************************************************************

   // Reset time Configuration Signals
   bit[4:0]   QOSOVERRIDE         ;// QOSOVERRIDE;
   bit[2:0]   BUFFERABLEOVERRIDE  ;// BUFFERABLEOVERRIDE;
   bit[2:0]   BARRIERTERMINATE    ;// BARRIERTERMINATE;
   bit[2:0]   BROADCASTCACHEMAINT ;// BROADCASTCACHEMAINT;
   bit[39:15] PERIPHBASE          ;// PERIPHBASE;
   bit[3:0]   ECOREVNUM           ;// ECOREVNUM;
   int        num_cycles_of_no_activity_after_reset = 3;

   // Common Control Registers
   bit[31:0] CCI400_REG_Control_Override	;
   bit[31:0] CCI400_REG_Speculation_Control	;
   bit[31:0] CCI400_REG_Secure_Access	        ;
   bit[31:0] CCI400_REG_Status       	        ;
   bit[31:0] CCI400_REG_Imprecise       	;
   bit[31:0] CCI400_REG_PerfMon_Control	        ;

   // Peripheral ID Registers;
   bit[31:0] CCI400_REG_Peripheral_ID0 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID1 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID2 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID3 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID4 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID5 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID6 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID7 	        ;

   // Component ID Registers;
   bit[31:0] CCI400_REG_Component_ID0 	        ;
   bit[31:0] CCI400_REG_Component_ID1 	        ;
   bit[31:0] CCI400_REG_Component_ID2 	        ;
   bit[31:0] CCI400_REG_Component_ID3 	        ;

   // Slave Interface 0 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s0	;
   bit[31:0] CCI400_REG_Shareable_Override_s0	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s0  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s0  ;
   bit[31:0] CCI400_REG_QoS_Control_s0          ;
   bit[31:0] CCI400_REG_Max_OT_s0               ;
   bit[31:0] CCI400_REG_Target_Latency_s0       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s0   ;
   bit[31:0] CCI400_REG_QoS_Range_s0            ;

   // Slave Interface 1 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s1	;
   bit[31:0] CCI400_REG_Shareable_Override_s1	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s1  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s1  ;
   bit[31:0] CCI400_REG_QoS_Control_s1          ;
   bit[31:0] CCI400_REG_Max_OT_s1               ;
   bit[31:0] CCI400_REG_Target_Latency_s1       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s1   ;
   bit[31:0] CCI400_REG_QoS_Range_s1            ;

   // Slave Interface 2 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s2	;
   bit[31:0] CCI400_REG_Shareable_Override_s2	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s2  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s2  ;
   bit[31:0] CCI400_REG_QoS_Control_s2          ;
   bit[31:0] CCI400_REG_Max_OT_s2               ;
   bit[31:0] CCI400_REG_Target_Latency_s2       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s2   ;
   bit[31:0] CCI400_REG_QoS_Range_s2            ;

   // Slave Interface 3 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s3	;
   bit[31:0] CCI400_REG_Shareable_Override_s3	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s3  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s3  ;
   bit[31:0] CCI400_REG_QoS_Control_s3          ;
   bit[31:0] CCI400_REG_Max_OT_s3               ;
   bit[31:0] CCI400_REG_Target_Latency_s3       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s3   ;
   bit[31:0] CCI400_REG_QoS_Range_s3            ;

   // Slave Interface 4 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s4	;
   bit[31:0] CCI400_REG_Shareable_Override_s4	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s4  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s4  ;
   bit[31:0] CCI400_REG_QoS_Control_s4          ;
   bit[31:0] CCI400_REG_Max_OT_s4               ;
   bit[31:0] CCI400_REG_Target_Latency_s4       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s4   ;
   bit[31:0] CCI400_REG_QoS_Range_s4            ;


   // Cycle Counters;
   bit[31:0] CCI400_REG_Cycle_Counter	        ;
   bit[31:0] CCI400_REG_Cycle_Control	        ;
   bit[31:0] CCI400_REG_Cycle_Overflow	        ;

   // Performance Counter Registers ;
   bit[31:0] CCI400_REG_Event_Sel_pc0	        ;
   bit[31:0] CCI400_REG_Event_Count_pc0	        ;
   bit[31:0] CCI400_REG_Event_Control_pc0	;
   bit[31:0] CCI400_REG_Event_Overflow_pc0	;
   bit[31:0] CCI400_REG_Event_Sel_pc1	        ;
   bit[31:0] CCI400_REG_Event_Count_pc1	        ;
   bit[31:0] CCI400_REG_Event_Control_pc1	;
   bit[31:0] CCI400_REG_Event_Overflow_pc1	;
   bit[31:0] CCI400_REG_Event_Sel_pc2	        ;
   bit[31:0] CCI400_REG_Event_Count_pc2	        ;
   bit[31:0] CCI400_REG_Event_Control_pc2	;
   bit[31:0] CCI400_REG_Event_Overflow_pc2	;
   bit[31:0] CCI400_REG_Event_Sel_pc3	        ;
   bit[31:0] CCI400_REG_Event_Count_pc3	        ;
   bit[31:0] CCI400_REG_Event_Control_pc3	;
   bit[31:0] CCI400_REG_Event_Overflow_pc3	;


  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

`protected
(dQcSb<^D\Ma4U2Q@HJMHM8V+<P]^PB9/c5Z/CB/4V8G7LBQ1;XH1)?X<E^:()DJ
=.SPd0cfPe<e]3^S3;&/ES-W4DJaac,FS\gAf\/5W77TIDP<;&MC=O=bfZe,6_8_
[94V,Wc4>22LSfYLIV?[2BF.N#B@&g,R7U^ZD<cB[=[9QVO\.>EVGF(MS?44F6P#
+&cRg-E&2T@?3;T(=^Z,?E)U48Gg)e?1J_KfQ8f>TAUBSNfE7(10#T[BaM1:g[M(
+1[LH\QaeJ,4^D7a?MGXS0)D9WGVSTId/RW2eOg,R.?;A0EeZ)f4>6[YQd0P8J0D
CKfYeH\6\AI1OFCUOJ[UTZ@1@E2.8R@ef2)cdEfHf7SU0NDMTX:4B9NPcR04YdX>
P.d5>X;[WH;_T?;^LeQM<?M.E08-8&L)0ZO?R-aS-c=&V0E]U0_aUGD0f8;SfcSY
d/=9fM1=S\W^.=<8Q?LIA<;W(;d?f]af_B&Ua4CJF787dN(4?Z8bMF-e5fHJH<)3
V[FIf;;d?JWJVQY]2ZJU\cJ@A));[.[g><>#&8M_c0TJK-fZ>2>7,POVW>XSHOI(
,GTKP;7cT)aU#L\<)]FO.20BXY_]:+5W0Z-FYHISYJQU6fg;-7K+RF:JPAddD@IK
gV:,Se)fAB^/(L45F1TT)3J&F>-MK,(/PL)).S+85^JSdPg<AabgOfDbBA)R/+Lg
9&_<X=PSR^MUb@KGE77,+H_()89gI.a\7fIQ#8Eb?&&eb555e6EF0<QM+EDDN+I2
Ab;HCB(aDMXMNLQ.8geERPd2dJT#CgP+.<0]P7_VLZFJ&]d29Q2\EJb+b^F4Q-.V
(CI6\e,()3THF:R?#W9VT3Lg1BFK?2YNSJR+d?(;6FQ:ff/[>4@bX>ETQMYSb()f
K@aC@=-0UfU.)<=5G7/;Rc=eK]_MEMJ3@;;f_&P^Y?6?24JC+_+],0\=0F<DfFGO
TOE\,>^)aQE5/>ScMMIM]WUUU;e3MLL4JLaF[+(N@PCDJ(D54ET2#0MX:8bQ-PP.
Z@4P4@@\GE.5Vb=,dDU5H[Q_-,aB3H_AW?d]Db^I,DcS#ESDP4PQgC#E:;KM,4Fe
L=VdNSD@FCbP[aaR48SVbd@-]RB1WA;ZB@RbV/7S9gLf.7YC#>eC_b)5=05_.SWL
Df:W=dNY4A;KRN35:CZ/HVaQf0J^S(5E<gW)^[D+NB44f>3cONAUSQ/NJeDD-b4F
S5WHY?()3(f\Q8=7VT<K>7VW?3QMS31&+9I@TBYQ=@?3\\+E<02E)-M3^f]:^RY8
+f#66P.e0TOIPJ3==0e6N/E;b</C43KK^IE]8BXY37S3,.OMQMYgbd4R.K15bJO,
V7D^1.G)gSSJH>e#?EJHFE2>CX5.^#N499,2T,L^]U_=#BcLONT>3_?g]TCS?&f>
BGV#E]0<GEHDQf/.PX,fI<E9&K453fPZ@J33T<@[,5\)f3)c9CDCG,f8A:ZPe>8a
4bPDJ.+F3CMfP?.TPd6VXBM4EBJ=)J>e#>+?L>VK(A;KfJD#5ePXAVVc?I>_4I.O
C-C5[8,)0\^R3+TU;]Q\UFZeC^TM_<5[f;2<KC8ecL-YED97?Y\H=GAUPL,bDC6J
9_8?R+(2-gJZ4LL^#/gT_NF3bB(4]O=RG^D>B(^EK=4A;MZaDgDX>dTS;Q_-<DJH
6AHfK@3gP.VNDPLWEM3VARHgZGP>_9BQ&R>S>ZNOQZ5:eGSD.Z7G@a-eVe^2]59a
+^ABd\)ATQgN5QC@N_M;Wg(\GXKOX7WC<PC./GUOD<Q<=JLG1(fd>\DReM/3KK.V
&@@5I-(7ZT>(^P&.4^bK-P0/EYXLZ/\26OW)U>V+\:)G&_],Qd\#@.LIdf_,(B;[
-LGAC]_,ERP7,7P[U^gQA+,?AQ^JA,-=F)Zf-9b_MLHPYI+G^BM6CLY+KOQP]D?_
8>_9Z+7H/CUb7g#UT[[AS94)S/8]RP^SM.FUXBd6Z]F^dcUEX[BQIM65HG#5HH9D
f_O2TNaQ[BP_aCYgZ8^XZZP73Sg:1/+5Z3,/0Y[60dI>\5f,Ga9:X=DHYQb5BD<@
4?)8_?1>7+T;HBHBVS4TFFZF[=;UgUOWA@6P<E9Fd#EG&d^S#?ZV#ANAU2BHKH:2
e>[=K4,0Ega=2P7@[>/0]&W4gV\KI_+#Z)N5AO7PS/,_7FI[VZfH&TPB/>1<8)V0
D3[P;_;6DX(4,2D]/64?B(=NP,8Oe@a;OT=)2(_&a[g6S[@S_c)2,]3V,GGXW)fP
G2>Y\^f6DQ/D3N-5_c:F6&Z4dT2.]0T:Ga?_BY=bI>87^YJYE2JJ(?C?ag?=f@9D
I,fUP=/3&6D0/=8ZTZ/U6f2IaL01(Q8\(W>,_1L4IEb<(>[[deCS),a^/OZT31X^
3Y2Mf&>LTUgYVD[@SV-dGF?4H/WO:-L^A&3eIL5NbZ#IJ:O\bcNJdg;We(]-S6U?
2Uf(?]LJd,c(8b+eeJ@bI;<-:O6Wc6Y)?Z+D^0.U0CEMb1KgQGFQ&^aHH-5]gAfL
DFQ9fH\/MGU1#5XYJE8#d)4Z)\6\MfK=O_<&g<2cH47a?.bW?,0<]&WWTE_\5U^d
c?^b_2;1N;J=7UV.&Z)V7^faa3(M,03W.KP1McM0-5C94XW[H2V]\&e_a^DZF9]U
R2X3:d]@1BUK6JWV419]4VAX=ES1^+&HTb#H)MR(PE?W^Q>]#[;)PYGDO:B[Pb?g
2^E-(EQR5<AM,/R[>C,V_J84WBQQ2ZW[OOET>#/7_O7+d&@STC)(94+_gMNO6;VY
\EeK00-H#_617.R(WQ/E]^gR7&2.N\[?<f.[Ag^N?<=Ja506Y^UF_@CL5VB(VW>H
RMg,)+1A)+>07B&a.8I#DAN2];]V<HEOJ-eC/YEZCDNE#I<DZ6Y:O_=48X_211d/
3JF4:O_PIDV>N0b=9_R7/70FNH4RDfDNaIJ8<SRDBXUQV.E\1;X6(QJ&Te;(<+XZ
MSA.bQ^3R<<<N/<>GN[?_7Z+BcHYb24MZZA9[^_5fF@)U@DeDS\G8L3)OgCI0e\)
L]I]?Y_2bd;?P^Fb^02F5[MTK1aWERBVd?9I.Z5b5Q,b2aDe]f())MA_;E(P_5MP
>[#V]I53O@Ta,XdVRd,E)3R2@&]ZWL/:JN=1SA^+Ob<8N0N9A,K,>Lb<E]]0_2,[
[3@<0Ve9J9ee=:fY[W(Jab5&Dc#,[QaG+c8U9LFFQ[gO^+Z9dVV<U>JH(dL--UYT
If@;P7ZK[Q_Y?RaHH[a(4A)JVL>QJ/YZ>Ie)(7C6,DdCK]U39.Yb0=SST4?.8G\b
UGENWRf(EICD\)^KU5/,2HX5Z<HN_OQAK=QL#1&B&063A3d8HOf2PF0.-P@F>&LW
#&2DedR[3B2LN&V?G;/b>)a2Y<<@)Bd;5QD#8C?5^:[f1^IW<QQ??)OKET7JSQS[
W8PT1HGE(Se8bGFWLIUV(P.9:83.d4)ED8[Y:7V1@c]9>&#<Z83>ZWQb5E<R4?W.
S05dQ-]UKBHIV&,I&7dd6G[@D</]<?\7S=_eX85.T+:4bHJYY8@Ha0[ZN91Z&GaL
-R52C8@X5)[0C\a:Wg93TA)L)UG@IJ>WG[01Bg+QL0)XA2Z8eVJGS#>@_FXgFJWZ
9)W2IJZ;.SL9fYJ_Y9-HZ9JV76\;Y7Y?9GZg7QH&#1;dSWS]>&06>9<-K:2T[T+&
YP\M+C&a2,OUP<CHE(K(WD-gW=\?I([W\<VHNa/7UWE;#ZbZUaF?cTZ),ZQEZ4@f
92+1)KHH80MBbZT@.Zd2\G4E5BE8)?VX@.bfCZCGVT.KMTDf(RB<=47?6F=_.4W]
@KOF;=;e4Ag.,\]JU9/OE-P?Xe]/U0_)#SK94R2W63.J,&_8d2_FADLK??F2Q\L;
RKTc+H5+<J:2-+92CDHHXZT1:Y>E-]S+g?GAUEUTc_dONa,d.=Y2-c??(eD&ACT_
feY3_,?a,UQLHCQ:Q\W^80?QdACFKF3=4dZU5+0D82JD6AdX+6O=:&I>)I(1O-gX
3@,:Lb5NM(H3fL/).R_)GHT==]UHf0b9R1[VKCIT=4F_K3^QG>Ne8IdgL>f4=?O-
@Y&U5=P;)gC)+Z_B-C;W8@>#NU&??TD:CcYYRZ(\&,V.J=ZT&.9M_NKM@JQ_\F7B
6@+X,OZ>9dG(AY^LNF)>.V)+g[VWZ]ZFM;#HfAN;0_\T8+a9<,@W<?bZD9.RJ(/N
-+J+AKE4PMXeHMU=332[E_L6@_V=DcQ:A1(UXHGGIXb)daD,OMJ<e0SePYWBEZA?
Y(HWgg..DT_5R<>>[+;^/b=5WTbFQc\[IR1TBJBbDKP47T)R&-LJbdTPfM[1D(UG
W?R(N4UD#U3>4K9I1Xf9YZA#=UEQF2e,-DK]K>L#8OC0CM0E0c]K,@dMNFEgP/Je
Y49ES5/B\?C\J9(.3+TPgO\M\P?->+V#T.)[Z8KNOTB.,B5_1OFc=27aQ:O?VdI:
.ac&,b([eR<3DSfWfX>a9Wc>U(Udg^P0)bOHQ+,^X\HUD6cSY7:6B\#J,:D0Ke?)
4F^RIGfB2N)N-Z;(eG4ESVK:NefN@U=4&OOT8V-N8][<aAI3g1bK6&C?<9J0Af&C
V22Y>&QF504<[.WE11_a&K<=ONPb#Q00Y:0=?3d[4gd7K-:M5Q]?&FSZIeOXF;d1
1SZQ=[51W(PES]4R/;Y>4EY/\Gb<4[NFB,1,UJ&/g8E>XY0f6ff9?F(;=#P#@C7X
O=eO6Y7Cad+2J2eB9^70[ZA3<^U5V-78R+H7E5[SQ,/:4:EMRC[eE>eT]?GO+RX>
BC2,KJVH^(PUT?+E)VX/C=T33^1_[ORXRS@X7G[5Da\/CNG#VRa,Kg+G16+GIgS_
_7PZfM.&72:\M#+#UXJe0C/JB=KR)H#cGIP23Xf?4>92+d2_VB<LfG1:R383Q6E)
T>\Cg>fd#XHW+OK2ZeG5\>WV&)S,YZ]e8>EI,A2=2P3:/f5eU_c.e1LD_[KGZ:QW
P3;ZEQaJ7g^,E6aNEQ[9[d)MeCgGJ-LV0U_B+61;J6;?[>L-2.R=2VL4SZ]<:2>d
TSNLaY><:EC>5gTGeTR&0;S8Be6AO.X0F#f@QYW@a36@#3JKdbf]>1(1W3ZQg46U
eVQSM4^SK?>7Xcd]>Q2Z&86Y#RVRDd#1Qff]RU;;_4^gEg,+=;M,XSFVf7C4SAVK
<\aCSfXKP,G=gXCX:2/?g?G;B/1MRMC0GX3>#0MY[U>,dMCSg7<^N<B)(,S5E)IG
P=gDL(?EdL_K5A+2+<YJE70GFIV>e5+(Z_\N,9>1d:?9(?IZd,/?VDFHd(#A8G-S
T^W=9)^])?^X#]SO618^#Qad#ZK[YTaV(;Fc82/F<aAU)LSV(&HPOb0[A@^g\_L;
XSfge=b.Y9-2dV3c:^QeM)VZVK6aQ@0H4D[\N(;NQS)O/D,A[YIB>A-(eI5YJZEI
MEWX_2ZR=;O6W.7W<R#_c:JT/O)7CBQ11Vfc9e7/<89P7YKF[^8bE@4MFNQ^d>g\
\c^cI\F\Ag#]aJ&_WP;)f?Jb)B=EEMd9;7cg9G48E,eA9-6?HE[N22Z?U?:B7GbU
46S&YVJS2IQ4I=HZ4#b0<&=1H;ERS-&R:V<EbbPbJC&&.R\)fX(#\S#V6-g_Ra7_
10VG=)A8U@N3X&.>.Y,5aE&.TDZ,/#(],#^fE-1]EF]-1KP\QQ9?8-2#JeZN5g+^
c8.)eQ,.<gMTc716JT<1QIS<7Kf&I>>f14SC)@6DVQ(_cM9fU#;LB\JZ6g,QT2R?
51IF8/Nf>,P.@P6Y?21ScD9cJ56BgMD#70?I)[I?=eIVR2Qf)1LJ6MEK3QITI0\&
JZ>UPZ=]YP&MMZ1+CB:Wd+bbSY&9@dfW&<c4-8Z^M>[[EaXE&Q.<B-HS>EDdO^9F
E/B\I&TPI3&P2;6Rd(75d,HLK/)?cZX:JA\\7:WK.M@L^QXg23DC.<FeQO=(G[Z6
GKV<Ae4^]Ya\/55]g:\XaXKb+&2DCCL3PM#af>eI(J;\@.__4ZHabLRB1Y21.P0-
1F@CS-[2US1Pb/6Bb0:NYE3MMTcfCR97T41Y4g6Q:_:P5]<;V451]W\?80+Y[[;H
T8=FBbOGJBd:6#3B):TaTLI<DQ.>#EA/;C^U1EQ2N0#CWWB70\K^^S_g/H93;ZU\
>GI98DR/A5W<_?EW?S6V^??HKHU2RIWeN.W4@PR5RgATUB8Nf02V^C?#4N#bI4:-
YME,&_K>/O@1eL_,R&N^81;P@LT^T@b^f7g94B_5RXJ9LeZJ[a1A;gCTYTXFK0dZ
R_^8RAg98^MEB_Z\10Ug4_H,Y<f,^JfQV@>&LJfCD1\&\2G3=Aa&Ef;N(LDa:,_+
6_Ybd]9g</,,<PCLNK(Yd@_EE)N#^e2./Of0C.O4aBO@96CY>@a0b7<\B1EE-Fa<
(1L]^+R\N.7b=b6VG:Sf3?KY\HC@+JRDG1d.PXGGK+HM,JfCA&S30aI.@BbC;f\0
RY<7\2U4V/+#F>a(UN@^UZQd5T+Q-SW\,bDfL&W_DE;U2fbISMDa?b7dQ]6:KQeC
[d+.>T?R8O\#;(.&(cbZEHQ,[fC8A;C(,LMG5W1.5JcIa8PBQ(<G\dTDH,fL@_6(
)DZBeH>Qc#E+F.\&FXX1-7I)PdUOE4NQ>(_ZbU^?=8RM[Sc8HO\=a873T98ALZBd
(0?8,E=C/IWVW,&36/:QMd<GG5Z9N-<B1=Z(b[cV?0IF80=(4)F.K(-,(?94>=/X
A._XDg@:]E=[O=P@2aIR,?8^2,c,2,:_;d3CC_;#/H3-bB1A1Zf8MYE]?A(3Jg(^
0^NW-Z56,&-(8+2[C<MP\WWF>-4b3-C\dA&[+51&-:)#d\IUXAYS8_X&C18::+BW
.6@-AWZGJ<0L8IW@Nb@dVeD6e/6ERH08&[&d0)(2R+fE6M<</N^V]+cFX>.+SZ9W
Y&@SV0cGE7YB)f.\-?[&@&LUXG-AZX33E6]@.?O>.IJ]Q2ZBWK-@Y48.]45;Xa9c
,VQTRe&,Z6cI2JR&1cPb;+Na^gMV7aY+M??G\OZ(>5QELYH:<RBbUdL/77EMb^#c
31)#=ePZ);NQNR(Q1SD<DHJdVgX^:GOP5E\FKP_013.(RMI\\Oc<Qf:-=C@4Pa7+
1e&ZK_&=O+#Sf-d6VI_ZgUDg6[J.)CPS6@)7]bN]E)-#&@0W5/f/,bV(WIcCNa=M
,d)R31c/f0?[\W-J,A@YFSa?D_.XC#@:Q:;IWaJfcd<E@Gf]<,dV]XI&^Z0,T@RO
9F@8[VZFU&e(^^PN=DE#c_XXT-H?;^g;H2ca:FNKV3\[Z:T;6FA^7E(#1)DOP7aX
a/:e1+8D8P<FI(87[L3^RF/6(PREG#QD&>b]-?E#g/;C44(eB06W&W,F/+XWR]AO
O3dZ+O\_R5-.DBE+:aDP&ZDb[EQGB1X.EK@g)a:QKNHFYEfSWf&VAMPGSQYYJ+&K
^2.^[(NQG&fL7(CKd6<8gAEW[<ACQXg9@9R][.M6AW&2/564^L0^f)=4?-bZ48K\
6:a-QNg6XMdM2O\e]^Wg06L_A-I3^\B5?c:/0\A=-f>;7W/<-f-M_3Z:F[)B5-9-
=YWMXR7B?.::<WQg__X-)BJ]G38[c6SI_F#<CL(:N;35Yd_Gd:B<..:UVEN8Z;d[
+-@e2>^d/WL]eadLa-8B_C_>&.^0:]M\[1P.3Q?RY)&?J7b2PN59(TA4T<M3?FVd
=0VdW@cG&a#&#BITH^C3Ua^U@_\IHX<92?T]>0Y2;654C2U/7<1UJEYDE@eJ15[3
c,)R2]/CH=XY=:JF-S)<bbUT[N^ebH6d75V<KH-D#[)[0)2]@0A(cT)1>f04/B;T
=;N>LVPMDBN0ET+BF)(P,=7<[W);eT3&\&YGP/4D4M7gI^=[cP^aJeF-;Ld(W6+9
HJ0B.1_acG0IN80JN7PE]G6D@/8/8JaaDQAZB0.e&eY1-<,;QVH#T9dMH0T@\NK)
?9g,.Y.M@HQ5OLF7,-a@9R0U(QZQ_C4bId.D6+KJO:UY=ARWX=a#3H>S\M+6A@4g
AW\O)fA]ed+.98T-1+96H<d2IX3=U808MMKS<#KJ1)R0UO0FC5Z^_0^-<2g7_e/F
+S<YNK#J@aTO.QgYW7?eO]eG2PYHXSDeU[TUc:JfL0I=UP@_GWRZf/Y+XaUU,Z]=
SO#3URC-;a?W15f7KLb8WLC;&K&;0]O4FSTWQ(aM>C&MP][@-0]JWRZFIQcA,D37
99AaT@]NGgFY<YT=<U>7E;?YX=4659SfaQ;_F];,(FZ1@UZ@;+?LW0M:b\:)f>cG
Q7&KMB=044g/),=Na=>C>4b9U]^@9@S9RY_TZDJ^VD2HbFR_6+GKbgCX2bOO7#4J
4-\dZC?Bc5GR=:C/C6#@f5W20MGPYC@<Z9WYfTW=-O.6F+-JN@7cQd_ca.6KaD0b
@\Jg<5SXfU/J&1VXB]d>_#Z\K]T^J.BS2BP<N#c#g6?TKgQS&^OD.>+]9WfHW(WU
XC@-O2UT&7I6129WA+A+<.Mc@_ET4?HA0,T2#\I/K&AN/):#6^]#9XgS(KV,Z&=F
6I7(3)P&(G]fUF->LYaE\3gHZ@A9:[MYWX]Sd>M#M\M(?B8</PXF@^LTVL]B#TEL
,7NZ8&V9P4B[W=J1RD+gG]]NH[3BT7LU6a-ENK/=#8DN<_M5dD,<V95X#F/K8=AJ
(),QL#64@_>.@W#94CZfU/[OU5Q1YHV^FH]M_3.f-g63I2.CP;MYb\4WVcRCBRFR
DL+-dX?3FTJ-/-1[Z)DZ66QB]76)d#-()QN9Cd==X5=7=]<ZRU.Q)Ra=W&L085-?
G+<27Y<#XOJX&24DXM:7\B>@.C@(G/(b.XCV<JB?G2]/QcY&<.(D?7Dd0P[Yb,PE
0WG,8_?=;[.XAQUUd#]C3(431bM_dH87_J;Dg<(T9aB+VX\S4@eR-6KE5W_\-1Dg
=883^1),5:=@^U&EY8Rf>2P[\=+RN5&+3g?/JR_+(>ROWS,[+1:W6,YXa_IK<Q&d
Z[7U6R:<^XWTg/XTbN-A,3Sg-#.1LI@[TN2FL1@<_-N(5[9X.YKO/N[(gD9aBNEd
2=4P7W/[N-;:2H;HVB)SZgJ]+C<V6a.f&/VB;OXR.L^g>V0PE(B,[WO,d^VK(c?7
,g,-.;4@U6T42D5O5S^1G/LUQ\f[L(b51/SJEafIdON6(I4B#QVPA<RO(<X2IGL]
;9<#FDST[L0\Wg/?6[2-6BA;cA#9?J^d\).dQ,\7<P#>O,9F(8PSMT1c7JLK[cMM
a/;Ag-CCgCb&1JI]7PHg^S@I^e68T?ae6JT4U>@C10B<b:0G^XNLK45Ed/]YdLSX
6QLZ=3[S#[Z+Mb69+6,GAJ341-;--SLPfU/,K40CcE#b]D?J84GZGgbIBA1YbA]^
MgLe@#I##R;MH8<LZ:MC#>EIWQGS&5,AH\T1UI4SSBDA_Q?>AP+WLA)<4O5JB@1a
I>0>4R/S3B9dPF>d30\b\#IC>3RF4=XC@K\P^C&:GH92;13?MUJQQ&N_I?PVNE[&
9_G-8+Y4&7J<Q;V3aJS+-NJ(?>3,eL3HX_Gb4ZD^H4[]5bcV>R@U9O9IeZP9J?a4
U3d@cA+)eFRW2#M2aOS:3=\P,>/X.,\JMGDT>,]R+.P?)=WLGV(6HAC)5V/AWN;7
60>IL+aS8aJ/ZI3-VafXEYXZIX>ZC<Kb1RdHMM[_<F4.]\eCf_4R<V73Z?.(S^^X
be>4MH<T6S^8He+-bBG<P/;XD/Fc9B29AW72P]bQWF?Je2/3IBE?TgY0U4a1XDL/
K_-8[^R&]5_G41HYKR4XCR4>;U(A2F]OERHY0Y8R-F9U+8K^)4MbGg06W<[gH_W&
g+YBgE#AX<H6c:/-e#aQcHA_;+U.C?OTC>I+RJ=7[I:208gbBY@7^FL@e:5I>.W<
GKR\\QWBb=6RgH8>4P#S9#(LPOXRA=BMa-@0W1<(aa5W5G6#=MeU:S8[8bI&3TGR
4QSBJY,?VN.O27OaT?N(b8.EQPX7c,/Zd00+cMHB&.:9f=[5W.]cB44,#S<NJK)+
C67=\T6QQ8-1J8X8f/^QXDI97+)7,T37DP_EV+-9I&HK>4SRK6(4]EWc&0K+TbCO
WePaWR]>(8)QDHbbLA682/S?CWVQb&#2HT=+NU,XZ[AQ/U3:7#dKQ6&C:;]g)ADF
;cX]N4+^U:U6-02dS]UD-Vd&P]KMK&?0D1^QfUJ\dY/-g^UL1:9]d_=6g[f=\6-Z
.>#ab_Q+fN@V&8P>T_3cd#(bC45f=J4H9X[.>NaVED2f[a7PK&^[7OeJ+VH\A,gS
c7R9;c?H^>MI5V\1PCR.Z->L=H2-Jfcg14@4#Y0bBd_McCS3A:;B5TMPQA1KZ&c;
Q7W((OfMMIX^V(e:9g^,I.;?XM8<Y^bD?_8+)?KUF:RYPeK:6V1(T@fW9)YM5f5+
W+^N3J5TZddH48_3N+//7cN,[+cN\b7cT8N:N2&RLI6MNW-WQ.7HPDVVT27fUD0L
O?XaF74.6&_L.)e#L]YO+3e<ZEF8cW[9gc,X79=083AMSUYd<2b6PUMUF0?91aYO
Y/RAGTDaKQeW#d&5WS8#/b3S-M=PP6eIE2R=fH.g=aD[K-8;Q(bfVF=7?#T4TM[O
@(.IEg7^+=I>7^/8XDS>=7,g^Zd?];H8S9EfXMAO/^(RaSV2BY&OQNbdg]W>&6\T
LE8:^FE2[5Q37:^GO(-5UOOZ:S_I(/3S8:/E7J+855/ad4&-7Xb:R4PLB=TU_PGg
ZCc5=;HG)b4#4U+QZQA]aW1J^1AIAMK&CCc\e#R3O#J,A=+1>\Kc&f1DCR7C)V9M
C_;c/4[\OIP_.d]).13^+L=7)1Y/(?a?&5:L?=)FM0UUgZ=K,U1c&gR2L[D@UT1@
&4N>S[+I1^@WV.Kg&/P\;=82(AYd\-VM=E^@7FbVOA])Q5[1Z.fUeC&?7NM]<a-7
:.,>\>-MJY0#U0g-d2L#g7PC-)]GPP@3[2?NQEAA+QW>ZE=,>b4:=-eAC+[0XMfW
d_319fSL/NK3?D7UGe2=HA5N&<eVRUEQ69N?__)e\5[#O4SY+4#@I,U;+D0?[<De
]<a4.gN&dD+PFT2-CW2gZE/]YD&?YE#/XU-#-17W_\Jf4e>H.#J^<MB/+B(4PPVW
XEgNcFgT)I9ALYb7E2-B<08S\GSJLGGbV@BJZ^g+LZOXTTcJL;?IX_)#E@=DgNd5
eKd>6E\D[/&3ZX]>(2T:&.AD+B).D\NNYD1LfYQON\bW1EL+L,7D,g-?fJ[.1>7P
Ff6?RD=#5,>@C4EW8d..+(8>0@Y3:#,W,EFcL8))+\d(GSIOXeSeOEJ<_c\48W:F
RLZZ^.H8.T+@e[eGO))Pg0IJ^@a-Z9/4T\dBVWPdOc_NQ)]bI?Z)),NHTB<H+FKN
H==AMTJAK:c,B4],(Qe3YYE#9M-1?-@=SIPYEB2+?X4a;.XK&N]UfLN1HPE1:Nd#
J[1d,VBM8ML[PN5(CdQX4OKT#CbFHTS+9IOO-9gXJ0IXW5]R?d9(T#=V5K7\K.1G
#e93VL01S.EDNb:-HJK8Mdb=BUX?_.ef8(@\(P2GA,IFgIdJAe/@,-#DAST@9]fN
>KZHcY:TKJb0LPM+UD&W?_dZb@ESc1S2gOU4DC_T9@L;[Ne=3<BV-#QQ38dZL(NF
eYB#-&5D#YGL>GVDN[P#^)1T\\Ia@WER#aB__>]N&3>bcM^+L,\R+d7G83DF5^5g
2U1.cVBR@8N^:BZ^\[?<XgP<QFQLF#HGBeeNWT\M]UcTH?\(>Tc;02;(WfJ@UPgP
QPCdY56V\1LZG]IL)]B[Q:B?GF4Q_E(58b+C:WB/LSVcAHPO9;/W8?8=\W(Zb=C:
+U#8;+Z8@[\THU;)XL>5=_a\8X)^)P4>IQ?>EU)1>.c-S.0/0HS?^\:KRA[@9D@Y
B_EYLaPC,4Nb231^ZK3:>T+?VPQ5Y@9+3C\2,:)J5Y.::@a:1YRLN2F\VT<[6d&_
R=U/4Be<R:d[3#<KKJ1cRM:NYe1bT_ZRJ)^eM,aP3;TT.R19YeV1&6/daT\f]O_D
T:]+:U:eP&F\>EIY=CE/6+&CJa,MdX#d.MbD=eOD#RQ/-6^+IO+LW70d/^S4+Of(
/:34G9I2.4J<&<4FF2^0gN:8S=CJX=eE4JfK6&IHK;DTU2\RM]E(8F-8CfQ_Aa0A
J@g=EI7U^&G0:IQJ+]UIb/N4WMfgHc]?9V#TYTLM5YGL_;)?Q&1A;37]RCYNH)&O
@7\9.b0R(S>@ZW5K<-/ENOU;0YPD;bV_P[<KUDK5C8HTL+Gf8=aHMHU8GLeH\0c(
#NVW.W8dZ=EZ\+6e(1,[_f\fQc#e\5>7,3N#V4J:#[b3LS,6E/FGF@^^R/Y2E&5-
]LA8:E5=NSWE([,ZfYXNIMDZ6K3Q-(&AE?Q3D.0#Pa(2>J@>Ka,K8Va[)I(b(T;.
P1LHHF=eMS[A/bUA2fY#SgNI,G9<Q^K#.EH?g&GK<^RLgN.JV?8[IEXc43M??I?F
)\D/,G0G\aS9fW0GR#Z[;V_QJMXBV4<QC3WEI_I@,e;;/g&6=KG?0MI_7-[;<EJ]W$
`endprotected


`protected
(LQM?\MdS3eWOOS1#U@Z-Z)BKXe,G=WBE,48G>5SY^dRB+[16\>g/)dR,BQ+Y2C+
@R3+eI(3==)J/g7@Sb2HAB1gZHgF@E2?QOWLc#L7[[+722Q-N^C5#\PUdGJ\Qb8>
D<N400Y9G&?T(/_a;]A(8;@MGV#I8)>RWb0A?O+HE&#d+-d1T&KK6cd5IKC0^M,F
SEFa9H#Q#L0Q:#7>240Pf,Uf?[/d;bDeg#c15fg4)6Q(M?P6aaHcS/:gaE]Y)_<?
/LGEL,P1:1B5YB0ZX4C9O2=0@39AGeOD7Q7LadTSND[?cQNHY+RP+gXL7&F;[^^]
T<9CDSL5\KF_KT)D((68+N1a15]0W0XX]:+W_K?\U?2LD9Z.(fXPg@3ENCVJ_](8
1\LBW@JaSMQOGQFF,gEZ?FXK56IK-3PDIB>39Nc(_&L@YeK2^-=\1fPYM?HcX;&]
Hc55ERfY2[C5Y-)#7YZa@;dZ7FHCF08bZ1:9]-g&G:THV)3((H]VK75d])86f:6Y
JE08XOFZU2cD[4]aN2b<Y_WA:WOB7aE158__83770EK_D2K:FK&>E60XC8F3X_gG
bR5[=+,3dF^OAV7Reae1PI6:BKPPQ?TT=]ZLPQLcX]._G$
`endprotected


//vcs_vip_protect
`protected
[5_2[P@\R3#c&;a0BeW+V=UK_+7_9+G[)U#C3W&]gY/BRMCP@g.Y-(Ka4IGPNK]=
aaW)#Pb\deaENe?;ZC\cBH:[T>,_BbWMA-WdZM8L\;3,,bQRK+==SD45UO>@K704
?_2S>2^]>\1+Ze\c8\>OF(IF5;a0gPN^U8-H/R3D#gfBOGS>c5gG)ab4H,X<FLT1
1:]de]Y#(INBRZ[\fGKT&IQ-W59_cg-O:SW3GB9E=bL(LbfdNJSC)[1WW3d@\D8O
5;(V89O&c\?@,+eW_/Ec@;[;^+2CcYdg6MfMX5d:LCOIbBJ0^58HH_)#MP#BKb5S
ZY9]SK7Pf86OT6DXSN:T<4XWDL\3J<?EPGBFeXM8I=CT<R4G^5=X(<5A+F[4@2JC
^_<gJV.J=)AM14-eP>(N<]cR]Q^I\K&RJ<I<^)J9H>6<.Z8+.H-IG7aWSE#e9b/e
AC17ZKN>PX475=X^P:9gf1=TR^-OZY9#U^QCKJM:DOCFbJTK@6,^^[J)89BI18gT
:K9>.<PNW;YMgBg@+?HPZ?g5U>[Y0HaYN/F8/4G]2XN?B+U.7VNaM&H4/ZBA)X]F
\D8VX@I;6@G>_Z9/>+-ZE;1N1;0XUE+>?8\AOGZHc_3L3U5O_db_LZ#V][ge=cPP
#CbK[YNA&@;LP<MU],V/4DB8[N7g30PTcYaM:Hg:Ja:2+f]KP5:OR>28?4_=G^5d
IDL.I+;Y3VET=,H-0/FV9ZG18HX?dd0Lg]9fLH)/#Z4cDGU@^4X05Z:a)Q&a)E:A
bX_dG&ad5PBbIZ&K>La;:WD)/1C3/,28L_Pe0G3B6)]V@gT)E@Kg)5W0&S7XRM&9
UA3<fP[d;+O\X+RfJf=#7Lb85:O_>dUM[WF4F:+VC?0B9INUFXca/\=_.U-E^;^7
8-T0KgR#E-[#/M=I\De7cC3K7?5:0SGR,?(U?KQH8F;CC&QNT,:VN@D.>OKS90I<
MPa#[39]8[)\T8d4N(/O?FdWe:d=7F09eG4/0+O[Y1DVFQ:Ge>-1(0K7_JY^_3SC
CMWAc\XdVT6QJX.C.\AM0OQSHF@390MN8CWV6G]?d.KTI>A>4MeA.N1gT+.C^aJT
0N:D[/a=GcKb9V=bWXLB/F98XcfIUdMWb3]U8eU#7\>+^2P+=>^^+XY2eASf<egU
IGQ+7JUCR::\A7.821V?C&dbg7#&YS4EO>3,#Te/^,21;A&8ER(?PJLb?/+eQNF\
5+G1_=T7?\PfOEY5&@CD3X&0U3I8gA=d#e)/I[b=EH(4<3NDMfQ+V5dUedId:GBW
M4S]I6R>,a3;NH(Q3IA^T-Y9NI#3;c_E>A243MaX0XLI#PCO;BDaBKY517N0d]9E
AV+LJ8@#1GKXJg2Bcf^T2M(4^=I(9_^\(&KQ8Y96.aL3@STSeFW-fR9FPX.Y99P)
H]1egEdKdSNVbMCYc;P3H4GYTfSW7Yc16f^QZd2F7CSOf7L:=+KD//Jed0b+b<,6
Z9RC<PGb-MeKT^J5DH.D^KVfLD+d\fZHY;9-:D#\TG:a=2KIa]8Y;+>KC]Q;D1b6
c@FZP3D+N=PT9a^31_C3_:[9>#;G1H&Q7)?[3^;=>HQ)GOTY_;_eX7Z6V)0L0a5Y
-3-:53G9B+CHH-LO_3B6YCa0&HKQ8UE=G-HaL#Z0LFG^<^/B2&OYGgUVH8(<KV0W
cW>[XYUT?,cE,PGTQ>.3AKSdSE4cXAXZ&TA\#ed.8E]KEE\P<SYOVLd)V<E=)8V5
+6Mca;2=#?-\78KJVJ<]HVGOM2I45T8E\EM12)-JE6b#?.6\VeBZ_D;W>2OWG_EM
VOL]\=^RM^82#&O4,1D?B]CDdXZ^01.3B=__;Ng\1Z>dIGP1D>YA1H,F@40K.7_1
\IO3_T#:]J3=7ZP5??fV.NTb-[.L552TQIbC[7aJ7+HK&3]c9fNeV3L\Z>=-(\7S
=b.c+UcAE07R7@4W&??\MR;)ED8A5Id:F]43B[c_DNQH,VB(cT?Y+DRPW..28#9V
,;PK+?4b@g[cgNa<g-09TDNJL@@d7BcE#dN6S2U2&.cERT.Z&\]^/91[(H+=aYT[
@X/17>WU;18\Qe(X1RQA7@3))/&+(7D&EPJ]cUWL]U@H#XOX+-4WMB[-(>7bPFCG
HT51E7X:0eT-@PKE^EMX+HLI[L.Ya/f5(217(I1H1e-b-1GLbRKGN^BINFVPMU#>
(BfQWC.,89<CF4(a>KdT3F(&\6b.Q+D96OG)b:Y_,bR1,Q<EfI@,#Z[1)c7R1;L,
3VW^fAZC2[^B>]I-[BdN6:NR#OE+3+EXcZ8S+PRQOJTX>7-3VB>.@aZ?f]-/A647
;K@\\eBGMaFe8BTA#XYZGROJEPW^J:c+]_QUNZaV\+bXWUfP7b&-7gJE];<0Ta^6
SBEJ>@^RE(5#c&K-,3FQS4.bQN6g9\1_]^<UafF,+7MS1Dd5?gG;R=0XC)S^X;\T
R2e4IK5Yc1eTX/:2g&6LD/2c573&6)e;_-:N1G_?ZI)A?cU3HRFK6W21c4EW?S==
#L=g]M]&^P6-+5DK4EcOMH>^JDa[2BcV?NYB]FSB@Na+>a[a3d92JH@8Sc4>8:(4
e#MIQC3HM+U30EWE/\g59Zd)9GXV+X4f1BX;RRGf>C<6@d^.FN7+DJbHZe-#R;B@
A8_AI6O#]42f[[ab]Sd<NUTS1GZc,#-FVKB952?D#S]G7NKcW6_#BIVBM^EU2IH/
/Q+GXH]XR(9gcBD7V\YM0S.=dUA@=7VEN#g>O=^+;7^?_Q[_/A/L#0BLe[eEB4Fc
+10SM3f1.?F+b(#IaFGE>NG68SQY&DPMSB75/(SVOg3TD/;J9PII2.b97SWbF(C_
>>52G^,V9cG5.IU+Eg81#IC19c-,//U=G#a<?<FP[.O0/8e,A5_\7CLa3>\)<4CL
7;E;Q&E(#CB2[A[4>?(&:]6//94I#?eG^C:>Rf7L.K#WCQ.]IYP2Lb=QBb6cN4<1
H]NYI,_eAME>cF(b5;.]RU8FeXP.DfT8YYgF9XaN8YK&b0XeQVZWED,34K((F@O@
E68^Q+e\2REf[HePR5]F+I@cRW5X=X<]c@V55Q5<#V)LF49\L=]-#Dcc@AR#JS##
J?WXP.3a/OEG)O?MMSX[3+6<M68^/2]V,>.S9:/HY[ANF7Q6d3S+E/T5+BVH,845
:J+^>8U.K5fSf]+TIgTM:CXKZX3YYE?C132B@O=2>d:UMU>7P0e4B17Sf(T#;GA^
BM_bN0V-+P<=38;=Y.LJMeZ-\KQ_.IbdIUTJZI,;M?L&ASgHP#g0=FTZ]Z;OIf0P
&R=[L=NP84aEBKX4IUZ:W8FAfUYCBEgf/fN,#67J#g7]+JQWJB#:(0T.P]2PSgRO
2C-3F:_e]dF_KM>-ddNKW?ENDP+BWZadDM9+_T@-?3IP+#X:U-QL<:cQRDMKVLI<
0N3C92Z3D5@E)CH(^XbL.edTIJK;39S.ZJ/OUV\W1L(Y0fK+Y@;FFOTZ8_5(2T20
82Z8>,DN624=(gKXC95/(O;>[.>KB,,>?EE)<76Y1T9_HTFP&fR:>g+A/;BBAEEC
>2b4Xb-X@dGN,AGB?-@a^[3B=O;eEVIJ8;(B>aL<S?a^\MeMWMCD6edEM8GYdZIM
BZR0(JCI[cPZe5>^-F9AZEe@_.PA\C2B7d;+LV[=FF3Z6C7F.ePJOR=F?TSaN&_R
S_cK90<E+Q,+TN)D8<:aV\HK[-MOX[]d;B,D+CGFe<UYf?BKeI.GFIIbI_0P+V8c
afF#Q9UX@L;CUH;fTLQL[()BC3KV;NaQJ7_Ef9NCL?0?\7Q;&4F(KLfc]ab:d3)^
9BR?0/5ND#O+5NDQF=gQ#\]Bf<e3.)fMgbPR8PWF^;TgZN,@;<dbg^/JGV8@ga#a
F.A7S8_ZK>@V()2JOS70V/_F-C[NXH0.b79S/8/J:<+1B<F_.#:-=U9ZA2#JXE@U
FY=I.LI&G^cXf-W[fZf,KZS@3]0>]]>fYS<7)&[5@:;[dg:.U<Q1^1IZ]3J?9a4[
6V;HEU8Ng)B8,RCO_59MXRTKRbIb_(b0KOU/-9\_b<3bWK/WI42I7cA/gQ,D4WE8
&=EREHV7Qc-,[_7Of([XUK^_ODY.EEYdQ<R3d<MD;KL,>(La/2CZ6^?JJN7XDSPc
D4IYOF3gY>26I2I(+.>[c:bN,ER5\dL)d@Y;PQ5#D/RQ9>,^J6N-#FW+:].?[fD3
e6Y?M+fA:,]2(BR3M]ZGO#2?DESe.L3TWb1TYX>dTBRDITDDgfE[M^\/AfQ6J^P1
<<_&P?e6ZE,WF0=U7?0SYHVR:&dNUZ[K(_82-;9gGWM];58_Y=?=;:V(Q1<Q1O=^
Q&/XA)WSVDT@6AN=d/W2IET=TMLe9gEK06PRXQ31JbcZL&4,RE3M&/ECNMPbV:A9
HV;B55+YZRTX;#T@5D9G5I\XJ\bY6LLT+[GH>f=CF)d5.U4&W(M\P>49?4A.I3)T
H#FQFIJ/&4?Z.<(2#bAJOC4._K079>T4YcWYJC[K4A#/UM.f&IG\,AKIRT\FL-/S
SP?\X8L9,=7..R[KG,[F=4(18T-FZF-.N)#5JHQ6E21PbY:3BO^QRbGVJKBL2e7C
T?S3)Q?(WP?#O<+>X72LcV/7(gGS1L?@:c,Q.SI4gAG&#eNf(L#E^JecSA:\?:-6
CLOB.&(=_1gcdZ(GTE.;DT4.3HM-BUA_YWV-TcfHIa?YgXaQc>(SNSFf7d84b6cI
J8AGb1M=dc=FcJ(QfV;e1D54F>8/KfW;5P:Z\^M#O^7^:Qg\\AXc2+LP?<J8OeJ3
O;;TD?R8+&^5E:RB[549@MgD3@d:6XH#c34G,/e-A,V@eNWP+R^RJ1.[>fYL1^[L
XX/fHSe6,^VA4P5)N17,5S27H,>47-I?H<V993Wa<Aa\RL:dZ+9f^g3R?)7;>6a.
Y&\E(R1L[OJ[gEW,#Z+S&B>WQ+bR;HK>PHfDMW@]b]9=[SJ]/&S4Bbb3AYT#Q239
:MSI5Q_OJ?+;<[1M:cWJgDJ&D4N_PP@>>UAI]aS\UJ@TVeI(VC+7/bXU7MH(^M9<
.Z)1ND:13SL?CK6C\LZW@W,B&(LD-f7bGE.RHV9(G2I;SN62+Xa?LIbBQLPF3V^D
fOD2+.f<><0JGN+fKVWGOg<Nc=fWX5ETFXKVGOXdELM-&)e[FI)1e^-2_[CJf^\V
7gQCN^?\TNO;I_NM>b7:#^,VfN9?XFAI[_SMPIY:86YJOWJUdEa33TNSZC_1FPS\
.I9;?KZC982SIf8=OEWK0b..Zd,a#E?fY.0AHD[FI3([_ee#7D5K]=a((I&D[VZQ
1:^:?JGd-:\=R&,ASU4ASX\#fSN57/UK]\T^GKbC_)Zb\V.K]]UO,7TP1KZY.@f,
.fD,IeH=^Q0U9VHX,/<;3TTBV_P@7gOG7,eU]V0cf^gW(+&Z#D(N.8Q_@^R=DED1
PgOgCYN5\#6ES&4@X[_,YJ\^b\=>;gCd,W(Y]9^f,__^,&gSTH,MKQ_dK[B5,2:C
B97?a,3BSCf=.0]c@g[[N^5TUVRd6d3UM;N9W)13VB<c\?-QgCLMF#=UBca.Od\1
-)H)NaTBc9Q.\HM824?aQ]47=<_T58SCE?+(GX,Da>2aeQZ1=YJ5)Y+OKW98UH/?
OAdBf3+_L&4:;2:)3ZNJA09H;e2I.2Q-D&U-G54>5?NLU/OML^Y0g,>9/d?N]T77
\V:W<+^0EA2_Z1b40)CIB=\5A+BR&UJTMQ)>eDS;AY7SD_[[&cAH?C50K@4/Z=L_
#3L<gUfZX#T:cRd=>aDdQS0VG_H=GE=+TLZ)]QffR_d05KTeJEN&bLU[S]_CcCGd
HbS=LBB6<CBFY:DBER1.4#Z@\>3bcgMg_^AIQW82aOHX#-T@>7gNcJZIW-RMT(].
aZA/1d^A+DQP[.O?@XM:^5<&R6>2\2#940;6F9CDSfOC,FHQQ[=.#W>Lc(f+_&0B
9V#f8XAL0Q3?PLKHZ[S@];e<T[8]c06-4WI7F>=1P1#gT]#\KeaM@5E,=??UQBWf
FE563I[f3,gFB:9QCfE1)9(@+MbTV)dP6RF0VHXfgf9[_>A[@?cMd47=OR;K5#NQ
A^aJ+fH8@4:6TUCf^(IaLC@H+3+\AJ2UE+6<P)T,eL^O&W)2+]45&ZUR9cSf7__<
:.&a6P&CdbX3e@OI4-^T<=:&.QWEWN,8f_[fa9-RQ95)GFLLB9WdD^&Q,A\F.A8A
)=/gQT,:G_#ZT2fG3ZE\;)MW\2L6gTK@N5@EDA_P@5H@<OI=>eC7.+FSA0<P<PFC
5P@0M1CM&:Pg3[<fZgdXBVU(&a86b+c<3=^XeX[XU1+8PQ\8K&VbXZg=gLS/A74E
@1UeN&RBU>4JC-N^R.T5?#fI[KQ//SE;EH[Y[aY4W1,Y>3-)(N=cgF+g]CSKENa7
\C7<97L0_f?.g-FT)1@EdP.T&-;F)YPN)ASe;O,GVc&=VDQMS;:fVNfT3e<?=N7D
eK3PUY_3Ob1:#<3K&1QL632D@.JL>@EE]]SC)YWbT-HY6T_.,I^G<M_b=M0M(WQ0
9.^2@b>CVBQa(LR^#R6#KHeRZ,e+1BXHRVPJYTGMVPfe6cEAA325b?590@?cO8A)
US,GGcDgE5CQeRT[58I33c9XK;W1AR2NM5[+7f2+1JA8D/F2=gOcW&B>\be3O]>K
YIbYOaAXA0J6Q/T\3SI_L17d>_-e.ff7).^=EC.badaYIa,b8&_CZ:+;;0ZBR.F[
K\G+93N@da.>Oe.(-Z\X(OQKR,G/B=.d;C+E+QdDW6^+_#fG[gDVf0OX<9dbICZP
0VG9]^DaN4GC9M.&2ZCB)@_\J96Ld5]10f:9UVbB<CA.&NQVfRK7TfD\8^PD-^6Y
E6=+^cFIY8CC_([IJM,@ONPPH3&SEV&HB3ac5Gc0H:EfbHdO8U3I].Y[0;=>[)e0
AAROZECcI8WaEPW,V]VD>=S;)VF.06G135g6Ma86?JD+Xg]2GII0C+Q[W#SK9#Z_
)M6GTTQOKe,b<(JcJ.Y>A:RL_?bA&06JD/36V89[>b/36-WUIKSZUeCF[<K,fPE/
T0eRaB_IHO3ZC/3dQY9O@fc7Rg2:cGF\f).F-XR&<D:M[a\OFV:aVU9^SI<YVGea
<g,b;@d;LPF:F)OMg@M:3\NJdQR],75f3\_MB@22[NDB.[B-^T6-/IWcJ(,1_K>O
61^(6EUT.UMAASSS=?C-8-B7J>9HbT5Sd[1+][3]R\Mb]5MK)?+OgQ\HF,66+(@&
#/^D]R](\P#NfH9MYVDIg<)dC))&33FgW.,+Gg78R2V@If^-;WN.E(\9#93[?g^e
2.[9@)))UHJ&0><Y;.0b@<c1Q12RJ16a[@GS8aOe^/UO5>@,FEaC)4_GdBY.^6]c
Q6I3Bcfg0M:?E7Te[N<Z?XT25gW/\Y\Da^e(3K3>W^3OMT89-Q,;fCY#b?OT:.cM
969>D8=?Aa<O@P(U+T0>:>[/.2VYb&d.?N5?L:WLG(H.OTfEBN8bRc;:,T&^-_22
X<c+]1S#Dc9R67?43?_F>L)Lf]33DC\&]\;PT?.,3Uc0]Q,_JTO^DL+=(X.&3bW8
Z>fYVZ1fPG-ER_cI;6B[8AcI6eWS7bO@.@5OJ+ECN8;(HXR+\1T]fgY@)23C)eJ7
MSPe_cJNaC6<@/KD^-6FD_&QS0>AdfII=XCWX2Rf>JgDbdGabR\I8e31QBYJ_3+6
\_CV4KcV,&MU>1EfIF>JadOUK;8SRJ(T?g6a&W&g&6G<g=;SQfeJI<S;^;&gKCW9
LQ&K[a=_9EFCfE7c[J@;fC6CY>B;\3F\Y^YC3AE.MJ58C1f?K-_R,_>dNFPU,FHG
MB==;eN=>XYAJ.KfVCOB)_6T_W^ZRT-&Y?d+)>4HTHIXK3J<60UC-N5;O4dRPfb9
26cE-0.8@KW;&.?M.>f]d7I&<F5K4>ZS=_09BdLI^(P<f)L)EALV41B^>&b&WG0K
^NOL#?R9Me[=BcZ<8FCV6fCP;:2-<g.?Z<UH&FS&/-C]gD_/>H5/L74f=/)Og;>2
Pfg5H^cQ#&U2gf-#P)J\cY[KYT3BD)cMZ]BG#5EJEN_e+#I]Q)JWQg:CV1^GBQ+&
V&:V83Y;[;U;Y=0VD;QKe1#@+ZIf-_edc,D/6HT<SBAfIUf#K/2Y?O0d.SQCNAeF
?Gd;DC_^(HcLYg_@+K(CI\e7<Z9:Q5.@gROfD>&[D6>KY0I2cURA/W9E^0FJ</00
VA<T1S+2Q[KTMMKE@ZeL<aG4B,K>7+O#2XNX7?1LC2#cR=/<NQ=9CReLV6Z#@VW3
((]TBaVEf8#UIRM.g]2,D)+;Ac6GF=D7VZ;LNeM3(=5YB-dV3=:#]bD<Q>DR2&>d
WNb9_RGEV]2cWQWT\=#3)7@JZE6FPIN:<IN^^;K5N3a<-+6BaP>9a+;@0[5e[R1e
EQNZgJ+@,\D/?.VZ,-Y]cBK=G;TXEJFAQ@1B>>8=JbMbgT1M#V9[fK+fZ[:a<6<]
ga/XUF9De65^V^HRDaV0[/FN6(MBa421fFBPB1[b:\\;0ZZeI8/b)FJ.;gN3AK+V
350cJ2)<L-RR[G:SCVJ:DQS)\JLDd@<,DG1/.Wg=d0@];-1C55]HMLE^Z;O;cAD/
@]8#BA3;+,H\/QI9&<,NM.E]J)EGB5/>Q<.+gFDH<<@FF7ZJ_;:LT^Y08]S@;#XK
-C2a-5I@FXU]K_JHU=S@LN=04<<B<aZGP8[Kd0>OdUY^Q;9P<3&?:T4<X53<S2:.
T_8->A,3W^D#fQL7c@/TJdM6A2^V>0LeSZT,e0IOS[MfI-BDY4G:+T:PRIO#9K]C
7d(^K)GdS2cJS4ReCF7f8BMcMRcfebWD@]?9C@Z.7#+65EK4f=,1ZR&YWWGE,@c,
9\/R7&@&g43M[T/-cM+L)/I@+A)@)T&WUN0/.aW\9eD>_I.AA#?@WD3ec5e\),@C
RE,OAaY8G;81-3:UX8Q=g?TU69PE/58KNa:))N;W:)A\?X^HGI-I.TUY.+?PZ16@
fV2D.F2/U#MOfPL:VW-^YC(L_QU3NNgKV.gP_C7WA=[ZY4(1IZKN6Ig4dO5X6T06
7Q9BBJHE=-4O;Z^f;<E=NfJ>CWZ\&F@N[@@a#_8<8_/>?/H(MK&VB@J=FYQ@2F>S
-[>.ZZ-dNSFOdU?A@T27EX8#&-A:Q?XW(,UPD(C4(;Ye<4LL_a9OTdPY^cJ?0<>U
-8,^;BeBV3UHPV>\4ML3ET??,MB,P;/^2FZWAG3ENCTf-CE@J>,g2G0,BF=TV+0\
0^9HI_HTRM@1JHB:ab=^TRUb:[-\5J,]#MWVXA)A.=<NH+?=)Dd3-1E8BEa2I/ff
/SLb[cUB<EB)M/HP3&FYR=27eM?WM<;^2b\#-4+X?U_EeN]>M5B2SNf+&70<C(7d
2,S,U^1AP65090JE/dB3?VK^5ZT.4B@7&:H#^_#@X>:a/2e0H+O8:IUMC6-D(gg^
M.(#YcBgJ19I(W3/1EK#fLQNMId2TR5.66G.Jd6\@P4cHU(I@YW\bV2,0,U-fCX5
d(Fc?5<Z4)^Z>ZGe\QQVS2abSF9c#J99dB]IKgLN@@aZALJ=.S)[3#3b#:SDD&45
gL=G9fN)eWIcHD8??98d?ER,CeN3]+^&:<<SU=[)70C3(CT8\dGKBJa,3gJ[^I:>
[(=JcBV-BF73^>[Sca/^#55-g&#Mgb5MFC-\J\bPa]\)CD0K,</5JC^/gY1F9U]g
M6C]?KcHXW]5JBZ]DaCM^_C8E[2=gQ9]?ET@4AOE+LTfOH&-9<b#A57H_WbSDND2
#fX^9F)L5SZV>b;VNFQc[2)J&F<OA)UYaX#:4&4XPO^[N,.0e8d[JBW_BYHaFg5A
W=Z^9H##dXIZMBe6-&X4V8?5)>MG0gN4<??14/&VFNKROOBf5eYC;4F5J-B#Z(aX
aXTS:.P/d=bbYDP25a3JbXbY#7)=U.HIb656_e6ZA:OGc<RBX#8J2Q7Mg^>9S2XH
X0M6WJA6D7U_(SZU>YXfbK;6]>^U=bE(dA\MO?6N,H9SZ9@:P?Ab^6WJ,F#+>)3;
3VF45JHFHY@OB>)A1Qf[)73>^.,G,O\85^JOf;g;>\8:)]1:S1DJ4G5>]514_Z:^
B.0&VPMEe1LWfC>UL.RVZCEPANfS]6)Z)J,5T(PC96=-+e4PGCYXO;&eYf69)69c
fZ?&=Z<2Gb&24Y:faf(5;2+UePONT0GHZFd1d#-b1/7dXV8=,.g.NL5?MKMT&fW8
d6A/]Y=Z>41T[35::@cCASZNBOXQ3MUSGfe[6[5JOEWJUNN3P<POgXKIKd/2J-9Q
;UNRQ;2.SF@4ECV==,c)BW>Df6N&7NL.<;SSdI0E/Se,<<XLR4[=aEG;STKSU]=:
=++XGK2T>95=^/\Of1(MP3ON1:VY#_PRa.(?gM\=#gBbZN?6ZGB&9Q;DQH-Ua@(9
2^Wf=M)e1LQ#2?Y6JZPAg)DGQHNbNOC<9M_L),BB2bNUV[C(2K0\KP[;Y1WXHGW[
c]-06RKg_R/X#RM,LU=b.5IeVd9T#K[4PH,5A2-g+V^3a[K^73(V[RU=BRIJDP63
=DCc5;:J()B;P43[b^>,/c/E45&NALGW<B]M>O5fc-1ZU]K1DIg3[URFM1^6P\5^
W2,deHK[#,b3-UP(J>IWH)YK/03NcV9C\9<7TK\Hg/gZR5\=fV>DTJLDOdA2BXF,
SagV5R_5+M+TgKL>2eQ:4L=<>(V>G[d\-cMCP[LM+R#8)U,a?W5Ge,9d;._/N>@G
6#NSgTe@D8V9##(AO)[SU@EH9R\-J=<VCYPE2(;\BUVI)D0Z7UV=#46:ePP6KOBe
0;A3DGVK7DQ.,?SN<.[_8J(0QE4CR7TP/RZdO/GbBA#<N2a&2/9:YNQ5V8YTQAdQ
MZf#K(bW+#dRbQ:eca2>G_bcX,=3[)N36?J_ZQL#2B9AL)0S?<YC[Q5,UI5FB)L@
f0FCG2]9_/;HTV#_EXcd6A@b@CE=+ZH&WdXJDe+-,&B2S0XgaX&=(4E3XgcNT,M5
99fU=E1HC.D+^MC+DeF\WS+9Q789LU-]8c3CCCG&fC-gJ2YWEE0WNZG5.T:2SDS5
,-g(dV)gRA=1SH[01?5@(1Q3G\gU]M1H-<BZX0N]5)^LYV(WT>ae[&/@VeL#XLN@
fD(1ZGQgDNI[_04][1)S[;1]cO;4HJWX&(SP^EY:9X]=)aS]I6:7C=]LP2/2@cX\
e<He_^&DBLB=3XUAWW7WWN-ANKM7EENJQ^Qa=Y\fLB^c7-aFL]RXe4]Ab4UA-XQT
cU2V:N,&G1W0TH>]AUXINPZ[ZVSA1OK4GbT-+5CE(W;D8>:H.\VMEKa_4f&)_fXd
<V0;>F>R)N_\EH[4F3MMK(A0LM7TN?\&+Uc.YZ/PP&DCVfb/474Dbg0,JL<]5a7F
c;5L_RaS-XX=e3Z)[g80EN/4RCE;C=7-c_6CY<-&96Q,KYU)M@A(e9?de4+)CY.1
R#d&aQ]6@X&OY8/B[;LBH4=;?fZ?bgbN:;U;URGWeOf_NI)W.+X,EJ/Y_/C2)3B)
X6ASO89Y9Y&:S6#@a>7M1U?e5aQ&XJ9V7#EC85d>1Z+f3HHdagL]88b9@LFe=CBd
=^)dN18Z;4@_LPBb5AR>f6-KU;SE/^7@TYQYF?^4YcG:W:TE.Ic&G082=9=R.;]&
?YJdK-2e_AB]4[S5]-^_UEJ0DYW6e6H,RDbe-\C14RG;[OL?@.,IELf3bcN1MRFa
Y8ZQ2/?DX/DNKPBNU?[##f6GIYZ#:I00]U8\8_KP4Z(V?UY@OA#F:.Z-QVDEA+0g
BY&@PMK)4[L5J(gdLJ\.304f([46,?FP5;34c(dWbf;3_^1H4I-37d^S)6U7@W-9
KS2OagT2Q6B1-deRVVM0;CD>[R--X7UP58=#X/<-+^,b#@9U2d3VE&//?IF0[_2.
\1\V?4(#PaGbC2&8Z/a_9g3IU-M8f8-87[f&=N6HT?;W1>]\G@4&(B6feL^IE/,f
]5B3/;TCFc1b:PL5W8JL>ZR2Z-\^JH+/Y?<fRc.Z?BVC5&VI9=/Va?]]4^/?I=bH
YJ[/]b7&Y_07.bTa-R_0S=UN4V3>=7W2W]/?MVDMKA[(>Kcf7T:U/<R5,b79>df-
KZf?ANF,7ORQ</a0YV@0\#X>?aQ[6])YDR&[)@b:d#0R1IO#LE\;>cYgXOG;Y(#5
g/MK?BgH[eK)PE#O&;(2N<4+aKXPHK1(Gd5IMFS:;S;MXE;\YN=gI?2SRVS3XgDL
B@A>A./D(&9Tag[HOU@?@+_VaF2gNMcUW72K8_784Ya9fHQS-F3L[3FU<98(Z_W]
MfQ2Y;f[Q_^Dcd^@8WbgH\,IM/V]eM(1JNCPg,FB9PbZ>&J1#W8BR<C1=)Y7_YDJ
:TQeZ9F0(QSXI/U.VOZ77Yb\3BDT8GPcSCLIT\/,9-(3GQ;2O:8H3#K@CM&Iba/c
:;cBa,_&W=\g,;\c^R9JB\)V8dLg7g2N+L?+[_&F?DSTV8d1<C8(9@[&-&L1OMCR
\R?\@^BLB,47\:[YfM?J+Z#BPb.V/[7/KGW,O<XYEOeJ04C&43:;TdV@\.=D.0<J
LZfJcFT[GDG]>W>KW_1=EM?/Je<W6BedU&9e7K;M9@X/>+5QS:P?RSaec.>a\Z95
EI.6EZ,5(]^-YTJ/M_\-F&#[/L#:=@W=7NM7HPYT2&TEe)Haa?T+46W+[R8WeCUA
W^c=2#gMY,UN98=#W<O>^aY(D(Q-bc7&NC,gJB-M7XIG+BV2>?&;@c/+f?HfEQ.1
2.#+LMDTHc49A?LW::cY>GC_]eg.S&Dg7NEe.9<PV?/C3ABd(;D];J&#D8<^26Y6
^GZ-\WOLDHWc.=d8>6./3T65\X,G\1:WFV7_/HTGYe\TG]OYCB^KDG^P=FRK;GO:
EEX>O63KFE&W0cCe#OLHR&&8YA9?\dQa?&W,N&;LHc3JN,KCXLT6Y(aBD3F^De#,
+^2IY4-]D>-Cb[GW6]V+1@6L;Z:daQ-c<@_JW-fGYb)\:U:NC483H>Q+6V9DRP@G
AF7+[L_^C^H?SVNJ9.K=\LPPT6.0P@:S9[UAL#JE+-JZY75<W=dMf-+NFS.1ZaA@
HVc)UcKPV>F<?I(ONV&-<?\183d)-WeX+^=ZFJ)Df2+CUMU<_6Z&\GDHD)]LLYY2
=^I(Y4V+5?\FNaTM;<8OH^^g_=9?G9S/>80NU]\=L8Fa#.+dL)WU(<<0J,M&2NT-
#NJ@?ZRD9f>3JV?c-HMb>BZ,NLA5-&KO.CNa&W@RNH9@RXKAL6c6NL0N21LZga^+
-DA@f2X()39-J^,V@)YE^\ZF\F(XLQIIXGg4(\IcP&T^S;I:A<2FF@-&><b0)LFa
+Ud>:Z09]IMfYV(:g[PO(MV7Q=?IMH9O-ZLa]cQ.(+E/UMfCC#<d@A0ebU1G;]NW
XZ\;K/Q;+Q2YDL-]a(](6Y2R\/SY2C8AEH+0g5MOVT:7,T>?BA,Mb?WfQ52NZLGG
:,LV/+FYEYGA2:PQE#VdQG2.\gB]1-3^_Rc6PgUcTR+aS^,\.I3^ea]Uf;>)#(d1
RZ-4;Z.+8gMd>XPD@FfD7@]TM54Ac2/Ig3N&gCJ\)\)GNcOaE&9:&<OY?FE[:3DY
0)W,GG/6(Wb8)UJDc8V&8=G58M>#:+]DDJAZRCUW>Wa?+(bg;RBY[gNN=:@ZIXYK
<QW:2aWP^V0dg9YgWV_==Od4M_;.DHUU.3&^8Q_Kg96g&BM<JF7S3MVZ>0V(H8UL
<HW1B4^+EP-\I<^^2[Dfbe,6#BG,b>ZY/M9(.,72#Cgfg8]ES9IRA_.NH3<dE>&B
e3#gdR19DDXU/?+L\&OY\?VfO7J\=?gM\CY:]G&[:2?RH5X&<2@Kec01#CI90>X=
M>;N5AC_1cD:(Z66J3,UXF5.H7e43^/bQIZ[Ye,AY^Yb<-M#3@Pd726SEa>YJ)(S
UBf\[V<aL.8b_7@]J0T5]HK-NAUDF5]F/Ab6-CgMcW5>;5.+7,+MHIKe1FNP.:&+
Q3P5@FdaAJ=5dOBaHB9d#:8)&Nd=@;&GS<D&\2)M-ce458KbN9/^@]QG6J5ScaOI
K69+6bb9:(CeNE#C]53V5E2?:]8^+/T73)CDS(-(d#]<EW,5I,&Hc-2+Z:342>@8
T-W==/Z,RgV[F-f1</\\g;J@7,P-\=<>9P?LM><2J;a_eAQ)C2FV]I#H^9-M4I\J
3;6>U1<D\<+&=#A:bD6IFF=0PeF-XP1Y.]SNCa&7K62B7]H7dJ:P5Z]U>O1[W&NW
,XSL@AGTYZL91d)[_#\^f2@U97c.[ASZ;Y@SC&168<N8NKHaC.J0O-[/-gEH4;:0
&2c/J7JNbe2KeN:AVC\+N0<e@T<_7b4568)?Q4-\be5QaU=F]&>H3)T.ID&Q8?,X
?.aU1;Waa5P/)KBKfK/fXb/;N[0@0+A4L3>U7FZKT^)H/W[8G_5MCCR#/bJUg91.
0.TPR>(e\_3NANbg_U?#NK&cG?D<0U5W)7?0=Ra4=a>@NSf=(B_@gb;L)ZbbTG@X
dSHW=EUX6D)TAWG9FU0^E>-5>6ZMR&[A,eCL[R<?0LeB38@gHG?OVAFCggCG-e\=
P&(,Z1\d<GZS(:^-9]IgeK1\9&dTX-HKF#..[7&3QP8dGe(9GNOC@C)R#>fKB28_
f>7D+\E=f]WSCRKH<J;4ASG_C^aKRH)2P-,#9HN84a?b__\fdK;0LM03QUVQW41\
HGPK+PVTYZ[UYdY:]CdU<N/>d^LQ24dd8V3@b6Dee)>U>X?YPIWB#S(@,RKE<f0d
J6=a]CfH./,DIOPL5dYVNV4Ng=]9bDWYFF#cf#IK(1^SP;9T+dA9AQG\5R/+5K5.
B[[LdKPH/0.6I@a-,R2<.]Ua@a<6[P66(N@(P#BB_S5V:Ne8DE=8FCg]>e,=IE\c
:,W^aQE3.:L[5(W-H5_7P=7M3O<9[9)\-^:+.3;.1^TDHR.2A1-G.]4/d)2C\)ab
;[,(&<),RXKUUZ/@FO8OC&e9?c&-5;#9@0b+Mc\SGX&M^L@\,MCVMQMJcb9O02;0
;654\]N]fR?f#/P[A>bS>^:K-M:0R^Ed<a;;Rd5\<X=XG>RT\H4c:Y0:;NPDI<,E
IVgTKeGKWPCNIZJ7F]+2VM?HB>9GPE)faLbZ48M58MWAZ>1O4CNP=M^5f:_/\b:G
>&6+cPLV?-d0fKQQ^ZAUO_,DW>,G[OMS6C7^R3NIK11N_Md\cCDVZS_,??)^6d1<
eTK\NV[4X-L,&>f/.CN(&<A2Q_NK#Q_a(ae2M(0/@?+Y^<g+F9L1OSL&\,F[/,RB
Nc?Ab>)?g8F6G.ZA4Uc8]VcBO@X&:X3E5#@L;RLbVM_L<G1_ZZ3\I/KU._:1,9]&
NN0Z&W)b:[A1D,W6c\(PCW?<DI<e.IF>>L4UWZC#b3_#f=0^>-Y=2^@(,Zf++0:U
;&S3-GbGB>,A-c8=;YZf&Ne(OK./\gBfV84D3[7#?7BA5DP8,_c2.<;Q;P7,3JX&
M^L566V5,(&QI#c/=L2;:#:R8&f(X/P:;EZNH8bPB]Cbd6cB7/OZ6(D-3BcggG&#
:=,L/?eCNM:aP^-AVJ1Fb[^G8Cg6:J:)DRIU2Bg&8(Sd7T4LAA5(3abR]DOCD#MN
M.eF(daTQFB5_<:?;fH=CcN/(B]?RKdg<:&^IE\LgCP;@^]7;EZBSadM/_RD?GF@
=MKZU\b09?\.=dGXbZMD:B&Efb<IAD\(Ge\N5e&G5?)Q&U(@YaR3[<9Z5W#UGa;T
CCR^C,T&,6W(Y@&=K0Y5:3.1@J7Q-aI+YEY0.5M2\J>7;-TAe35PHZ:,V0WfP(@U
].>A#=V@N5E?KP=05/[:03127F\\b0Hg5Xf?d&D=9_f<bg\4D:e)W<g?>#\dZFb(
?UF^D-=]VQaXL\(2#A58W#CINUKX0XESLJDR-2DeU\9N7d(f375;See(T)(QD)U_
?;WY_[/X^[,NcS1/(R>TZQ5C_1XRJ/^88F2N_8DCLBLaaQ>[,ZFW?INAf/d[NIH1
V0M4@(T7Z_XV=@<<35FcK60,]FNA\#E6Y]ceJU7@K7&D5daH=ZMc\@QcI\I]f),e
KCKI6=4eTMFe<--2_VWeG(EY(1?fV)2JN)E:TY,@]WNd,QUOW>DdAc59<aZ8,]2E
F988&LAe^L(fA][LJ4SA]B8T[XWZ7UE[M#E?^aILE@1ZKaebb=O@4E++F_SdB;+G
H2#V?GH@[3cICSQ6E/\Q0MT9)=?:B/ZVMS851DJ81Vb7)O]S>SY;\SXK3dW7H8-e
70K^FV6ZZ\e+U5H)>7dKTYY/0]ZO=c86+KKV;gH,TBb.44&?J4cYfY?3]eT8?P17
.^]&OOAF.b/]P/U2e?>3c84X#@U<aE.8MRV5L,29T_RED<<D>ZdC?fD[gW#I;WZY
YOFc09JD3SF[1_LR3D<b:\(A43cge-=Q]9XN[08U,aD#@0S+DWRYd?fT]7@c[-4;
?4Y@I+SUg,8UdTEO.a2]JND;G,O-Ke/T,IORJ,fCGXJZ@+W&d22330.NZ4GWXELQ
1I+>0&eWScbc^XA?BFEPVc<@W#.dNIA0_VDS\gYE.>;>S,5ca-bB>#5[Gbbd&3@R
]>],FdU3TF20B=B.@9]I/AEYY/#DGaD_T.Q\\^N2+I(D7aP=_&X/(RB1>(.>E_N)
,W:&N7/W5\-E[-f8F<R9;0;]A@_U&GDT<LM(=/21(>7CH2cX&S9#N:aL4FOJ8CL3
,-&V^8NW04>dKRK;:RBSXEIP\BGKC]e/E].#Zb#E?S==NEKL&+bIDX_([27QD)&1
bd-;6X1WOA[EEY1MLe4(VZWd@13]PHMeVW<e9J4Lb7P2bW-4FFM-1<Xb\ZY?=ZgE
b6AdA82-R+Y<AF3(Bb_0,>.2[-322]XY4<HD;_-;>YII6-@C09gf+/8RO>:?P&@c
efZVGA_?P9AL\P/SJT)_S#BTE/=+UX@600,I+@R+Rc8[I=?FRE<65^?.\gJ<@:N5
\D?f@+Ac2d&;09NfBd(@\IA[WW^.[+XL8A.ZYOfE/,9A7J=Gc^^?.EL1FWR,-FYG
,@=dE(0ZPd2^@NB)]LWF^,B[V#cB?\85OK5/(I6BDX?6[AVZT\eW7cA0#3+NXQDN
IHP)\?M#U42;.9=M^V///-CbDX((/a6ac1#2/@2;5QC)72^/J,6O_J0&g.4g@M?;
7Lc,4Q,F-0d#4DFM?U.<9C6JR9X<+VUfYT=]/QVIT7=adX+.+:<2?7/#-URObH60
->+V2E:@.G7NHO^_?IMc(;a=b9N[.8>=9#L#++]E;L-c0IRF<.P\OTA^H+LR[7ZT
(=]cBZLC?:+N23NXH_:@c)d,gB<DgQfH6d62R&)&\f++&YRYCF<XB-O#F>G@cdMe
YAd/KFT7#Vd;V(3T:[7S\?f&7aeL#,..;GN9/U1X;3E]a8ERH_+<&W[2VD6TCH8:
Q(<K-L?4P,0PZ^)?=)+ID/:ELIWNXSbDQKG&,Lfc,0<S#9W0SDJV3Zd\/(1^PH[N
NJ.53/I>)KZI<+.Z59S#(Nb+3aefQ,][T8K1TOS\c/PJ-P)0=06fBeRH[4Ya>M&e
@Q,)bT:([1OW)LE2Q]YE@:@J<Y9A5.QgfG#C&T:O5AJe2e+c=S(H,?gg2=a.5QdT
WB9@-T7<FGS\A>55L@ZT)&6O=fDW^eeYL[D^5=gL^^EC:_HWdB2MgOCV:H.X+[aC
/,KE-LX51C_);QT.3:;PAF&6b@G-4-,AZdaOc+(U95=NdRP89M,(6;F#bB#A>@^f
0ACA92;,>G<55HZ6V=cB2\::[@ZP2W@<a#PQFVZVK3e6O98SeECFU]J]_F=TM89C
b5)Y];.ZHR],XM<acGf7?fKRS#VF?Pa9W@8e7K.7AY91/UD44HK@;SRW9.8aG.&?
dQ(\59EL\?0.JB)&M>4.HA2Fd)R+Wf]UU;9#,G?]ba<X#CBc>>Bf>NX/C\BZ5NZ;
(1IF8A=fX^H],d40#05cD&XQ7LeBR+KV)#_BM)_6R:50]RYW^/a->g-0D49]AZD9
-G;-I-^QUT;11/d56/0,6?10/H;3:DX7]E18-(9Le0;EEGR(>;J;+&QSJT]&aK;P
Q7/X8L3154Ta5Y^\4LTc]]f59X++:.,\=VO4bA-^N+@c]6L(EBVeYYWA_[IbVL)b
A,BV:GNSg)DRZ6CD)g12Q:BNKCI@/KFC30/]-fELH,C)H46d^S3FB&=#?7_#L40K
LG_O?Ze3??QK+I0bM5eDPPGJ#T@\/7;_^72V[b<JRX6U,QBUFS7gZC&HfS,D]+Y0
Y=(KK>I5)1-)cC+2)3E)P;[\XL0W4G1C]IO8__(4,bXG>Ie)-.>VI6)?(+LPEUfZ
PS_=I)dB(:&ID@/L+4\4Za./UeAX9H_PH-(.@NCB?(L2)K,ZEDS7C;Sg>bcR9d_b
+7>+A4^#4@9LM,#N@ZY6O&>QfBSE-+R@;cO0W]5+>J-F3@-6YW@X.>H^W-]b<22a
WSNMAI/Q[3CQ_U?Sd4\PL;b6RSdEYAJ<(\6U>B+06eM?.]IO?T_;T[NR.Q<J3VDH
&0H/\dGCQ9c6-654\/[Ef9]UX93Y&?HKcZ3BTD<;(gG4/<^>NP<>NTZHd/-ELUVY
+Gg5U2P<PVaDO>#^=XcG\KIU0<31KS^WU7I3PXXe,[GRbUOb>1WFJ_BgUdfN&aO#
51d,H8Y7Oa5U(RecQ\K7\&O]-g[^E^&P7/2@KQ_I&50Z?SVReJBacWVIbG0#FC85
@F75=&e6f71[e;P.=LEfFXM4LcPcKgNPXcgEN>R#?#;?GF,JDTB+0T>]EE=6W2=X
X)^XKaX347#F[M_bLE4;5ES-D05@4=HY;]3TNe3(7\^@0[V/SSCWNQ5TE)^N1FZT
0473)\?KEaKHJDU@Dbfg/[?Y?)H_XY=ge(dXL^a7FN>E32cdNcKaK-L;1M+Q,)f3
S14aWVc9Bc#<[1Ca:66@3N,E)_#PK.;_;UJ0=#V(HHQJQ&PSaf[5FR<_,>G5CKN6
+NLE?G>HNKOFAM[TA-Ib:O+41:XO.8Ba+P1XPdFIYG1O1#\16-]\7@ffce0B-6+=
2.3+eK7FQ\[/XMB)ZEc]:NLU+-#\3e31F(5+K@8dTOPGBaT=<UVPTTCOa0-5GMBc
@?KHEgTX4[H=0LAR_/#TBNdA]5SL^Mb&?LLAVKV)I4U\Ye>1ICTb7WMM<b)]MB=H
Y+MGZc:[01?J2#fXf:FS/3#EZ>eK-IV_edaNO0L)E)V,=KT+/Z,WC=Q7/H?2<c)@
5+P7JMbLB,]E6PUE2?g<U>Z;dcbg^e#MWF9aZXY/<-aP2g/20?W.2Lc-PaIFQ<?;
Qd0_H_0K-XS6148d8g5WdA[1HDf1R^M9GA9E54B8^_[WcP2,P=fac9aO@UP&)#B3
,7\>Y6-[0eE_52Z]Z2U?<.D59?+MLC=88Q4X;HHESTS?^H]I)c[WIS&]U&5:&;YU
TD2\8\?5/F,Ac6N3[?(3BLc&+gI+b4TXd_5BHa+21ad0R/SRfD:9(MC-T)f>\ZJa
UF6eHAYZD<?)7):D]3XO@3RefLV\N-dUH7R^/??)B2f+>/g@42)U<Z6e[87WJ3VI
@H_XBc#5Q]-(WUa7>GVIT3IXB[@BZ\8M6HZeSFMd<PFV3<^3-7F_6[#-AKa]WYbI
c]c=W-GgJC3<9N<@P6I.O01<<be1Rf4Pc<AD.)eFHM81YZBO8,b2SKO?c8Y\N)6X
Y((41U+TR6DU=8OaEW[P+.PGZVf[#Q7?YO^?GEf^ZTKe8?)b5TIU@7X8WQHY_-NZ
D@,(TK9R>9;]d?3;&33F[(bZ/8Y;(V19fFBPI]YVI[=+0]XSTV/\d<_.CW&2?+(Q
2O]?R5#1B\=AZQ05WSO+fJQf?H3ffF6FM[P_,]L)Y-GXFUVW@\6GHTKHYd_<X>EJ
?(;C2\@G\1I>JJ/:/F;]W+.6Ea_:JE_6/g58C<:FWW1^1S)FA?7/)-<=)-/H,>[-
=EMW^@aBE)>DL3C=JX\9Wb9I#eCNfZ]E\f&/ZCV8c&;N_ML9KX;[2f5[g^GaAJFM
BP\8-P[\:O5IY8U?+).B[0C47::0WMaEBDKN31(:,Qa_]84TgO?ANMD>-R0SY;SP
<#cdLaFFF4X@J>+)NFFF#]IBD2@ZV316L4QOPRacH-C\cVN]gII+<&0R@C\6L&[?
_7O>9b4\PVF7C^EH+@MeIKZH^R8?]Hc3XW>(HH^:7MDFXe47LLPLV-N)3d?:]V7/
6\2?A:cC;CH8FKd4dI^#@XW\P1Q:,@ScgF,F4KgA(1R(@#,\-EF:>QO1R8XFF@L)
5IZ1b@>@,P<d/7LNe5+D(8CD]S=&C28TR=ecU3J7[edd8J>@)LK<d1Z,+9CdH5dA
5F7.c(5^DZG+?(6ZZc<]8AP1X23O0OcL@]@UW),R_cV8\M<?_6#HDe=E/OZ9?L0Z
EF.=MLI0b?Xc;1@fV\_fPOF^Y?-Ue<,N=fLN))(e>5?S-F+<B,ATL2F<-T;OO#S)
a9Aa\F9:d89[7T.FR_=3B4a?(g&#ZcbMaTI4eg[>#Mf6AdQP_V+^L\ZIU.09G^(O
^QUV<?FZ71S@-d4G_,Ga6N02.X-gNeL31S]6eY+3]JHHW05UVWAC02\g[KKc.:\7
)/;?gWA83bB+9@1Rd_b&I9f]b#&c(0CO^N\YZ0VJ-S:cZg#XCW7N\VeZKL2ePC:H
HA7E1NagS]?)J+7]K+?@F45LFfD4B>5=aXY<0;KcKW+Z[c-.gPLNHDI)#^3<ab-P
EOFLF(a2)fHGe&Oa^53<O]N^VH[b(RdL2EZP9TgH_Q#5VXcf?IBGfWUI-7NTO0G#
+Q&P.6F>R#+[=60+&]T7:1I#2)^e<B^R<OL7D>g<A?=XN-cb_#N84YOV=N>2/Z]#
2ANJ=<M4cO.&R9REb2KI7fY<;K,5YLO(/0Pc,-V6C._)-0bQI)4<IRD/>[?YW,OB
8&c2JODB4XBWD>0\TQ3OD-R.:+FMd0H,YK0CV3M?cXc2-GMK<gCd3fFcJK+d]36c
V+c7eLNFY6/+E;.9bA=JgS_:>cUVU105@W6^IUKX1RY:ZP(4Z62dSBa@,De=]5O.
JbH5bLRAW<OJ<IO7:[NL6/2T6R+1-D93S5b[1/:fa>:,<Wcb<>I\(6L)FBPbcA+P
3Le.,R<SXK6WMG3?_P]3M:9U+^3)M(GLU+(R[=g[HJ-ScX1g_MBbBDK6:g#EZ2N_
ObF3fNGacLT?/H<GU<>^cRN]RbY^E@8<27>55-d?Zff=2S<MXD2cS],b6)34L7./
(VGM&fOV7@-8FS[<#\5daU>.M1?SM1]EK12XVTD34]?\Z?,#:@L&g1_ETe^@UXZT
WI/a4S9bB^8MbI[BW_Q0^OSTa8BfX:eKTdOAS4E:@4]+<-OaIFHRI/[g3Mg8^I0@
S2?.@1M/PVJ7L5BDH\83f1D)Wd7?7a.<3OX@.X@XD4U);=D_DGJZ6aQ&fE8LOZL.
6](KNQ9B<R^Z]7]#bSV@R(^+OVZ96Zc6Y<S1O>X=YeGbG04HK8&UO_X3aHda\3H\
01>c/XfKR1=M(5^]_)?cPd,e^&Y+:JfUNS^2^JIae:K&\OWa+,T/.B_HO\ENHD.6
0@P6cUfaM9F2ICK>=aLKe7_dP,YY#:4aOGO^UfXM[RKV]OB(=D7c=6H3a<fgPF>1
RDRe(:bgf4TYbA@BeU-ZU0=W?_(b&d-<2,?\_TD&?(VIUB:VCY]dG_#R76YV=:R9
e,Ka7A@<@92V8+ZSCK4@O6[<8BS/:@F[;F?U>a?R/6e<0LeB?bQ@&aUCZP;4=2<Y
CV50^dG[(JDZYU(4Z0QLPN7DbL\0EG+U2^EHL0[&0e.Ud4]AY?0]ZaQ:W1=IRQFW
.c1VbeUDLGL7fZe2G4_L@MIF.--?\K:f>B9/7d/bfU(TAcN(\X@_):IAE65-@#f2
UF?b4Q_:cPG@0e8SeCWf.JfUL2G>0G/07=T&[_S^MJ?H\FE^Pf)M[P5VU;7YWYd2
9U.W?_P,&(F_:F[3UW9>CA-95cR@8gOS@J2a-Q]XFBVd-C_&Q,c2JHUd77C(PH;;
gI[\S:I9+;U/A&PR8(]VIB_-=f^-Z+ZRK&Z-N4DJ?>,=UfB3.V7XE75T/<Z<gKdF
Q-[1^@edO6f+A=BeAR5fN-bHKWN,^[;G9e0Sf?_4HM-_R7FY1QNU\OX-0I3:#D(2
e4+DS9M&VgQ=XQRQ-8LW4ZM<FWN(L2L/OKC9Rf.Y+)3KJBFQ6FcGb6g_J3&J\gYR
,Z.efUeY#RFAF/MTWbeeRSI^24LLS:c@2S:\1G0Z@-<J@E8=<Dc8]^Ae).L1?/YM
dV5BSXU5-<5A5Z7NB>X@^S_5+EP+a9/5H/\]H\b<IZGfUdMM<XGKVE3a2(?<V:OH
Oa-FbIBM9_FaKZG>;[<S:0g9JM9MRT).PG#6,\e>]2X;O6GceVBP):V;EHW?3:K6
:_.aeU(Z6^<c#HGQb;7@>3HTFK5>0g2GQ1\O8RR@;UXPcf,T:5g.7+KH0MDOX9?G
f7DMF(<5W=4K:.@JWLfAL_+LR]#/74N[5@agENC9DU#bG2]OBO(C_1f/cRb]^=ad
_S03ZM6;PDEUQ.O=b,-MRBTH@2dZAH7Pd-Y>Q[45g)0XeY\?Tb:GG^.AD;2C->aI
,BcF)?M5.G+2CdWf@8U[F;J@bK8+&9?]LLSG<O6IVCS1+CVQ]YJ6DKPeSRdE[=YZ
P/If1_Y_R\WgH)(>Te4L&Ae7&\B/4BT5N(#JALXb_QUbZ0@69[XF^X3[V@aCG,a>
dP6_9d[9W<O4+PbC0DdO)0U(cO<ROTW1QeCZW0-BYf-I]THdZ[FDT]VUU&83=e5.
TeS49<TZ>2<Vef+-7HCF9P>#N\_U5gLb@1fOU27S/50NeCX)9;Zf?\BW46JW5_L.
[f77NCKJJ57DG+]2JXFO>f3\5><[&^MKO#:bE\P7];.f:[5K8V4R=SDAScCN1f)(
0W-+H.3DPf,4Wa?3bPb37L(dc\U7KQ5);6.4VCQ9A6Q^2d_.f-Zd8:[4R(6JTG#L
:IEeS=>U1T]<=If,U^W&&L1K>UK^DbAPb.Je3>YX1;_=C<S]S+1Q4U>)4><\e7f:
<:geg7bB>/Q(C0T/#a?@e7&BI]f62.NA=-VDY:5LV,29,bQG#2844M44SO(BCHQI
=PXV,b2Ng0ZUYSI2?N.3J[F=fc:SKFL:XT^AK@9&9c.\f?XQPVQ1[ca.(G:Q#;H8
EgGU;VX;7e\8d@)=8&@faK[CJRS.DE(THL6UJIVCVb(BODT?9DEG4;Y1DUV0,KcW
H_\6C]UO,&)M9Vc(TQ.6^:.UY(51-bDJ1+R&e7<XJC,@Ta>8Z#I4X^3^AOa\YL]^
WO-@5,^\#I0eQRJE>6JF5eSL<KXQWCT:4UA;@E:5e&Q+U3-N-gJ),+]0.VE_a:&S
13F[b9YEcDZHY(T[A2_D_5>)AN:GRN-)1NGO);5Z-@9XNO1NO]5\+4>JK^Q?[],#
YSEM1R2+-5)L#O(R^f7HfU6?2]0),IK<4acT5Ta;8[cYW;]8a-\AGf2/g\/VO^4;
@100#[:6;IMd]GfZAI7,I81#T)R^?,W(=KYg(8^@V(-G5BFYgRCc1fac)N:]dY4-
O?^QcY28PIeX&T8X=YFTRNCeg/VVDB4-[4-&c.O<Sg8W0;0S:>#ec=c5K/ZNEd>I
@K/YL>GXSJ-Yd8Q(&KV:<H2aTc#K^DOK+479S2dZY)9;e4^Rc-D2Z6:SG^--06<E
3<Y,W+MHFg+/c/CLA+[_)VS:KM/^G&4Wc@7.2Z7RVQ&1#/[KT(TM5W,44).f_2W=
c[f3POMAcW[EdNHE\^-eH<aMeFf]MJEAYE_:&1NB7JVg:LW=MX,=#77Mg>fbPF=T
Y-9JW_JT^T=QT[Ac/5^g>UA@V7H6CbFJ/f[>G^/AQe=B?)MKWMaYVYKJ\f^_YXOL
dW+3([(]W3-FO0?-gbc=\,I45#N.L#9g7G0=:AeV_2G@Kc.UI0?M,/=T.3UTF4B-
><+CRX#?cKQ5X;XCDS-E6GEeJQ6U/1f-]@R,.GJS3a[,GHKZ>#N[WTYXCJRVadB@
BcPZKHR4fT^GANa[JbBR^K0c8J20C;eE^+QU:d/TSFEOcWc8VgK=PS4cS5?_F,d&
Q;&RfbSMcVb]NBK;G;[_\..f6F9N\fT1\(<4,XD0KM/e&4G7a=,SRJ;14&=C+SVd
.;:X9OX5OKJ??=c>B99\b^LWeR/RgbO292[G:QTJQ]5I0/;gUV-+))ZGcO;=].OE
C&J8.LQQH68;(g@CC-8((5-a.[C>_A9E7JE9?e/3AKCML9LdZ3F61eCGM1H3[1<R
OOWQ((83?RM<&CBGCd_Ha88.PME.@<2#a.;(aMd4DTTbg&02C2Ha&[:)\6[Sb(6B
4A_[WGfTT/RU;6,9X:Rd,F94cH=L;c9PQ.10e\.-b221,/ZKIK@Md_N[e)I19@Nc
P)72/RG1]a]O9>5=&-J?&VddUTX=]WLH&5^:TE.B.9+\1MIT4[^(9.KTDB7ZVF,D
K?#Q6G=:Ddc2L-e0+AdTff),7@;2cd,O371N+[4QT>97M,OQZ3fM(DY?=VCE6FXY
cT\,EV]K/HVO)TS>?[A@8S^4^I<2#62EVIMQ)KP#GGTGO1V/UdMC1U+LBAa+I(@c
+J>1f@\X/d-<M/:VH.H_a3HF.\B^M&H[5&D6YK(,P&-a&CDdP3P]/J@I6&,<6Fg\
e5=3+0G@H47A^\0>/NO.VSC\(M@RGcUg-84CK8Y,X_62^P-R[2;/T?gP:BP:0W?Z
[#gJA/fg<M8JLMK2/WCbQXc6JY[;,gJ^5#=E)F+ZLIGDdZdS\<76CbMOb_2A\0Dd
M^>1W-N)gL[<5(R^_-X9@A@a#cgI2Z]G:61@6C0Da4+,RBW1PO4_P.-]KCS-_7R[
^[O?.L68gG&4JdZHIIg&0:YOc.=NTL9#=GKa>MQcQA6QA/X0ANOR,T>UHFd_SD>H
.0f2FdS(F,QC@gM33eV1-=?IRaESC;PE]g-B1I<d)YGL9^37JJce>FXV9(J-[/=2
DRT2)L&gN,(^D^_@0#LZ##fd2FJN8?ALZ]?O>,=(M,bW^K[;4BLTg6Pc8ZDR2/d-
8Z\2Jc:H/52DB46Bb(Y_C;>6S^0=#P6B[&SY=&XW#OeC?45VMCeU3(W;3cW;_)F1
AM;FgP-C+ZHGacM?1-JC8(SbQ6ARaDO#9AIUD6cTUD^HIP@+7U^01LO5ZQ-+fC#?
/&6G)ZX&9F]O9=P0KI1a:Uf,aZQ:Xb?J[cTU5GAKfQ^IXV8.F^4=Iad+3T7S]fZB
NL&)-W]OCQD&=4?#+=LfL+2ONT2CHNI4_?J,R/1cP;[:L\7>g\F1TXXeS?I>]KV>
<f.1KH[MUH4FY=YBV5SgeU<S8(2=&;:.]d=f/Mf-/T;R@A/2f1S1=:5P+AT.W+W1
g0#66AB42-S](=J:fgJ@fYX^P>PFMZ/RD5fd^5@,@b2TLG1B-/I3TOW^Z,I7ZH:9
G&aEH3LN(/9VcRD8>Q/\=SD3MPe)U@I(]QZ1b<\BI5O[:48^J3\eU&^DNS8([?+.
K/;TdF:37c3B1=RTHX&+SNYH9;Y/TX1:36F#)B/.GBa+&@YA#4(ZHB069P;SH67V
cSV?=7Q4F;AK/J)2X&]BTg2XA,ED>]\.NH0.GH97)NWcOT_P@6)cE;SEP?ZC]UTH
M(8;6aVdBKWZ(7GFGRU?d]/JKXY<1LT,^\B@]\G+=URM>Y(09,,V^:]Z8?@60?NN
PM=J6c:YK(O,Z&6(fbY-<+(YTBW@OHLIAcgC#f1N2<=GH6gfQ>]VbM>M@_a(bB\<
4(YX6^X-0dK+V4H3>6F:&[D.2,:+7OZ/V^(YVQ)ON&Zc>1KBHG+YI@.(VEe>OE,7
I;X>(8@^BXQ0=gHGGI6&1+AgU?8(:eC#&Td3(L8;==YOA0&LO9NRNgc&^(<c06R6
70F#Q)a<YE&,>R,)c[5.-4WcEEd@#D,-=LWVP^?G(#-^5Ta<ZM++]9/0ZH6=]bPW
XVA)U<16KM30LA7=[+1g@S\4B+>JYQ[5;CA(g?Q]8<?K[TBg/EMBDTI#X7;TEB8U
5TJ61W<J>Mg6<E9\RHd<:0ZZJJ6-dB\5K7@_XA_dQT<F-_DER^^_E=.g?69A:cI5
aHJ>-fI&&/TD#WZ?VfZWS\TZ8,VdcLYM8a\)Of0UW]<J[c+XP\XXacQ.[c4-F,QV
?_4?.g^/C)R;&6#C6V<eT]6O(Z-NF3>deRH7>E#7Rg[8D#J6T#W6@C-:&eU)D+MI
Og>4HWC1V/&A)Y.=.,4HZ>7A4cT#MBUdV3FIB;C0H@DMRQ#IT#4[][#fMdb/^+cd
[XD+d=Q^>EQK=9EJDa-1U-I;K<^YISP_Q2VJMC9]ETAT\)?9_[AM;cTUV1U\AAT/
X+1Z#U6YS09/KRO;FY=QAf3aecZe/B.)B@]-WRUNVU+H.R0J0=;1QMdIc.K[#^e&
+<CKPbc[R\6C=;:aAN/P)ab8;Z>>#WN?#Tdb4+G@ES?,C+Q:N<5EWV6T=Q,)X8@&
_L=VV\-.5V:<VTg[RH0&>JQL,4\/IAR^8RWBZ?(gf@8d;V,D3R>861,M&#gYYK=4
cCHF3=7F+SBK8Q1JPJ<MYcT_\=:f+(6=bFU=;\1A7N;+EPT)LH<T1@+H57_+\YbI
)Lg4Q,IcU+5;HV\,I>g2^0<]]Y:0;gUZ0QI&UZCN><]8JJ^_CP99S[A4L13cWXQG
VJ0,a3S2,_HE/.);-GZZOgVbL/W;GLfQ\+2)#?e4>/:4X;BJTK+-&8R@N64IQ4CP
Uce;BJA\3[G/N)\M[Q)3VN19c-g<3Y>ANXZRc\OW6(WTE>IPd\0?QfE[SOO)1_TP
,[gHJ_)Gf670(<=^g4<#O6Hce>N,ZAVT#Yb6_JS)2;dQ0.>BdaGT:dF,)7:,TKg)
#9;20C4INM/-H4#?E;]ccJBV>f68CJdE0.SOZYJ1f57Z#<-dH4Gf0Cg?LXL>?VYG
L4YYB6+.@I^g)=/@CT4V+J[+X\9DcX0>e.LLV3[:3_QL7<P)d6<1XKN=#WW0KPd4
Q;g<S:SW.P:V^aVXBaJ)2dg]ZC<-1?#JUA)N/J1c/?[.#G[5H0R.cA]R^WV&-dPS
,Oc>LX9I>7d6\])]H1Gb0L5J1SAM1/F=K8<HILS>SA#ER;R0dTRbg?7#/gD<+@A:
<cfIGf]\-B4fVKQ3]KZ=O.V1WS0ZAAeKe@)KX\=R6EH>(WcKIEZ^S(-b@WSf:5Ng
DNGBNW&=1YV4_+VI2OPcO?A/0132[VJTf@?];U7RC__U9U4M5F4UU)f&/QM]EV^a
B;gg:3I4c;T^]aJ8:UQ:H?;9+G))5L6(0\L(]6&:WT5Eg\dZ<TMI>MRe:55;bM#\
]MV_55BF^I7&VVQDVbJS([@16=HG8e^@:#+B[_K4WBPW^b9]6QIWOM+P/M/\aR@9
M@6F5F4IFEGAaG2Yb319TEB,LLI\&VGUXMg87^-D>1c:gQ0b&f0&QB3c_70\-T>I
=VV@cF/O3S-6XORKMEQ)e?JX<OFTY^^M8+\],-PZBCSDVY,X26;8(Y/_5G5<ZVN)
H:Y>08e74?O,ZWF9gXUB@Hg9HM?.40[GM/<Z(H9A9Gd4Le8UJ-71BX230S#\&\#:
g?3:(9KB:KMI)C<c110PVa6;9II6(0&MQ/gA8[26OUN@ae>-bX&[gHS)TB([P]dB
?=D^db>P/eEA2A+4NRK]Ubfg;CWYB.8FVVO&I]Td[SF=[<UBZNTaT4FXTd8e^L3;
,G)T(UY@8^/b[I>GHPM20\=KeV#?983@d(W>dGWG-XHN5]77V)UJ(JCe/d&-e4;N
gXI/,c6a0Q,K>W5dRG(3T>FSfRd]+TY)E\C.SA;UR]c.R01RMdAAb4)7P5LKdK,U
,;VdS\IDE-&1/UON4ALaZTKW_,AD;>a9Ldc]F]Y0F-^3PYY,XU>TT]9DIDPbW+ZY
[3fTGSQ3]@979X_405T1H];WT+;[cNVEb(daVA>H6d&H^R2YbIWVFdE3CNRKKKGZ
b,dBU<FO=e7+4aZ1((?R#e+2TFN/QU-2E/53\.E?cS3:,ccFRW654P#;DAPO?#T(
QIM9:]1L2,^>+W^#[ZA7U&U6N&?[]LA#,XHC3O+ZT<5>dJ7O;VD+(ZOY6-,_.R_b
ZRK]6cLX0#OP?@PU0-O\74T0TLAJ=Ge/3a0#/&CeD#0QM69+7/Ob\7^c(C[1.&:2
641)B=]7@W6<)Y3-=\a]/39/.,VL01J^AFIYHV&EEBRM7A8+/+?MI_GRR#OA^73e
7dE_PK+S\:#8dcHX&H>\<]>]Y90K1YTH.(]O)[,>+-E(caWFc4#Zb?]/K8fTWLJB
Nc&OX5V^CH^T)>JFV7/:P&Y+(;b9)aaN)F_B?]@_-ALQK(S:9DGQd;NdR^YH+5#c
8C@&4Z(?-<];UfH#W)?O?=MSR)JYQS:P<=,7e?:edKC#(96S6Z6_bMHV7ALNF_1_
g\)Ia>JHODcT\g3N1V)^dc6-4?KSc6+QdAZMK9XUJC1(&T8AcV?NQ_TR3F\6GY2@
6SRO8BMCCc3I#AI),KWa+)4+H[JY3^>JZ3?U&R83a=+FWK.9.9d1+10#]f[O5K-.
CE=.9W:0.d/HHLX@\92)3.&)U8J=^2UIO:HB&-O7Ze+R5eYd@NUbeCUM-]dGS)QI
#8f1FF#>D)0_VAML:9Q6?-6>^4.(326PU_SM-H>ETMBEQ+?a<,PDfRLHKBf:d)@,
?QQaMT8gc#9aM8Y&7R396;U.,BcY,+H5DI#a,8?Y[):69\KJ7WR\g28;C4;XM-8L
(KMa11)b/f&b=\]7\;A\W[1LN+Je@WUCORVOP&&Dc=Ve5Y6Z,S7W1Ad3S]FF9;[V
3?GF^^]g:A-H86BO_RW6W1eFC8T5J8A<APTF#2-RCL+T)UV,GcZSAM2f?@Y/:/T4
EM&M&Z#>4]?e^GRb7_AQ;8L\6_=M\Q9cHL00\WK+8J\(<O8DYI,N;SUWbdYEb])O
0JYa==\YdRI<^83)NgGN7J/D&-b8G.@-cJWBDcd6P4UKd5:UG,U-dfXf[9c.Z-;Q
&.e-@@gS>7<AVe0E,0fff\D;.gBFd\GdC8TYC+PBR+,T0L3e5dd:?4GR>APS<#4H
>IE.&TE=3@9K+DNT==3?TSf?gZ;]A_Jf3T&W2^JI\]UeC(,-cXPG,UV;:1&7X.OS
\6G.R8Y8<83JKUZgX&35R)-EY)gUb&:_ZO/4ZC-PZf(R(X0-DMT(RDAHG1URA=VU
CM/Sfg=N;E_(I:3S_.)>Mg=Z<+@UaJb4G.TAC1I/(Of?A:3<6P.HcZK3E[9WTPWP
7<T&/\_6T:g>XU#BCJRbgH6^-\@&LJ]_0HQFeVQP)?SKD_,9,3f,c<3/ZZAc1T-=
E;3]We=g2aa-^^(cT2_PR^LXU::>>(0MX_Ja7T<?Y-^M;&H]Y.6Ug>@<YU.MO]-I
48RNeW:XXVOU=3PC@3T0BF[(M.23W=OD?2AMcJTP4:S(JOAB&QBY&D2PCY+PZ7NN
3AO4<)J:&5cR,SZ(&f#\D.46BEQ:\Kf=XL-2G1YMBEOS]e9KSNV7&+UWT9fC-X7W
Zd0LPNddV-+119#,PRH?-PFTgc)<D&701=:9[T&5&c@G?V^>3-HQNS6X1AMa7&1B
@9eRSaf)S6@KU@:,4WB8Z#01NQdNVfS_=;e>g?fLFbUGUcf>3658=LCR@<WF2Sb6
[CT[,0HGP(QCY@@M6V_9bH,QQM2Ld1)WUHHUW++_0+_6,Fg8]6WQD7-[Y@B_I\52
TRU7_63G).0dSB8J.RV4A5:?O8B8K98L,a[(AATKHDZPRfG:))XSQ8]T>-EZHJ7F
YGIbRP)HCgY^9I\C2QDB4S=+12X2_H?UT&YV=/-K<W1SU-L-?>K,8/23)G;&6b62
4Z,Kda/0QbE2\eJQLH)H#/+7DK+VRKX#dZVTSH\AB7,=@-bLO(bF7,ZH/#]C/+5b
,)P^2^K2.EB:#:P67Pg;S\78^HZ;9O-;[<&QWV20GF:7>bU3(b;5Q5:#aRGN7OI\
J0@5D>GHEbd+[W3UaSJD8C)<CO:6M2#R>Y=VX[2e1[Y</WaX>MK:V;H[NZ90]b3I
4]Wg()gafAEaW8V27B:IAa(3C4fe-E<F2>6Lf#EU.&^e.>fH<Y/:]#J15U#IfL/a
B]QeR+Z]KDaKB5C(=F^C_)&)^gZN0,1c86JaXbgT8H/d+UdEHgEG-+@\DdeZa-L&
M_K]?CQ5a23H4bCI:<KQE=UGfFYDf5,KCH0OXRM<8:6(>GVD-CL]RRGXV]&8E>@.
//?\<5@4&3aA)FO3cBP0#=BSJQXcZDCaVLIaV.?&Q7J9ACb5eBA\J&^2+B(?\gPf
83>S>;13704ZG+gYbM6ZaE+d,8PX\Q88EZXOGBOTNW93UD7_C]&OWFX0_FU/(-eW
Q3;NA?3EZD_Q^5BV#X@6-DST.?e)]9M+>L.J]O&,I+]OD;V]e<A];CL8@fQG0;CD
ZbJ7]L,(#6)d;4U0[/\).I\M,JA;B\6<ID@\+QLBX1Yb;(g.D-#CcK2\IHQTaHB7
+BIA^c2+OUA)+#JN<-VC.OgFPb+M\#QRe4>O\(]S]d@eZ23CO-0.f7F4eKR88#LV
Z=+J),>V46b2<b)JO)08e7P4)2QZQAK9W3EfO7C2M^Z6+J85TJW2Cb>UN<NZeS46
a)N.YGA1BJKKK==14HB@&J2I@77E(J#+\P@]_;&IW.;F.e2Z2S0ffVK28I^R^6I1
L<8-/B1HSKg,]5XI-O39,@I.eQ-c:+,O[3HfS,LLc@D-5V#\>_EU2[CXfN4C=2\7
1aK=5KVZL.<.Gg_LUA]K9;gd;,1MZ)MS;R\J<2V<0L:.PQ,;c,<7\g8GF?7MAOE#
_?451/?<:>ePGCX#C<X45UK+#MK=D0]UGHGd@4?W@3NJ&<>Db.Ha?]gD2d=@)-eJ
JPT9J3O#_:c,24I/&IF7+#GF8U_e_6AMfe@PA)))?GW97QJ)V@Hg&J,1(9887T4C
<YZI07(_HW2>E&(c-1[Q-7@edA[d;6YUL@7<SJ(gSPb:EX8bc84K^,AVP?;+J#\W
M,;0/1=E@,T4#aA1DY<b\8W8?=P6_0^]MYI<QVF]/5;bbf,=gVVP69eJY?=1YU?6
4g\>@T^TaTRg(g;DJKc&W^#J+]>\K=\B(B0T1fA2:(0H/IEg\/3e3>3O-VE7&J=2
47++g.P859S0(0U]ZYZG2+NY.1a;X9(<F-.>,&^BTRAO017Y]KN9a@;ZSL?N:6D(
GQ;/2Qe2?I:Vd,(AO437-&AE,JV^<fUBGOP:=3g:)ZA9.>OUO#B>UP0^_W]Y1/.5
OF7\))7S)AEDG;K\]4=Vac\;6E\T?58?6OHff48@^d@H4Uc0V23f4^cL;W8(.?UH
<>TY</DL46VR-aCPTK:DOc81YUfBFd,g,XcddZ^]+#,f:?4<e_DUcJ[YB6F5T4g;
I+f1KLV5,M3(<D\^@>1g).I)&F&<JB-Z,?SC[\8K9TALJ5W]W>W6MA9ZTbb(?Cc3
/0/5G&KY5>#FK#I-_WaN2:XY<(TPR-6^7.8d1(3cSOE5I#:6F;SK7Rg3?5U<e=JJ
-Z3I[Y4:<GGQ^@BBbb,gZ?Mbg,<0.]M/8Qb.X80L)\gV^LGF?&C/gd:Z2E=6400C
2W&&;Jbe(FGE74>-M_>/J99E]1TMcI-OUL(eHS:D_]d,&:.:SK\_9.+_W>NP=\U;
OEP8bTFUSN;7WN8AK[+K&N.Y]R^,Y/0D\F38H+8EW3SGPC@CUJ0U2OIa76I6K&(<
[A=eY])GEXe7Q4@FY.L(ZLLYUbE5\e>@^CbVBU+<7=6(ZLVV10-^JLd6.,;CP/@d
Oa5HR1TaH]M)FX-?-9?43:AYc/9a,?ddfLE1H0VbI/:B#YdQ?>(+:>5/^bYPCF+M
1ZG)eD7;HdUQWIdfGN2:a_D_SeM-H[_0.PGS/D9[ZC?(C<d8(]SI01^WXF2R?6P=
C<E0U/F=[PD4NdQ6(K3ZKac&&L4V+g8->,._XU\K6&O4TE4?NdcL0S)@cA>1Hb3]
VO?VcD&cQ_NWR[Z24D#AObBYJ6KFKHN>(Y4NL\-EC?6_XY38S,9W&>f,9Z&]<?_H
#If)#LBN<2>1G>6d+-;/+UQ8YUf;I3O-5&7Ka,;FK^S#FD1BP)^GI-5]Y6K9WUG.
Z54#f<Qd<g_/PeS>[@6@RVX#DZ)fLHaf;4F^Y+R0P@S2?B\NII?\UL7Fe@B#AO@2
92I;FKNPaR3d8f@9(B9ZK]1^1?G6F?d^6@VLKa//^A/9/&I=VP4M)aS0;VR8a56f
ffdK9E1\7YDZ5V.1\fV,8?2<\g=N&J[eQT5,I/5:^S047L,MZf7aXH:PWE10R^]_
<U-+?#43+cB0@K853;4@0W_K86=+SG1cO0V8?]ZD(K#^[UNX[B67G\Z&BMKB<)@J
^P?7ZaM&0DR_RBfS.Z6JWa)KI1IA@E?G(O#@;)UJ<F&INN62;4g;+\gV4:>:^/_T
Ag[c8\B996_S-JM^CO&XBXP(d#]4;:TcM80^.DOY)g8WI(]fCHV46,&LC2T62OdA
T6\)1fe5R3?CL^,Z:f4D2?;WaG]PAX)H)Y).,6(D-abG9\&DZ]HR0I480TJ2PZ]&
b:CABOSVT=BQ=^Ne4DJ-#EVR-c^QKd\#\Y7?\)bba:SH>Te7F0Q3?_,IeW_2L[G@
C9KL0QJB6\OdLT-KfdL895^OK.SXd>.6aO.5S]YH)N-:>Xf2K?X(ZGEY])3&(JL]
D=GPKaDF5A]4-OJ:9R7OUK]7K3aMQUN9&0=6IZdX>6B4S-d&/68LQCDgF<fQb?5U
P:EO4/;(.DJ)aTQb([_,G#/#d(,GDH2O-MU4XR3TN#b2O,+bU;_)CNgdS_PFQ)2W
aHN#c815EPTT;)(#9f-7)P:WOJgWJPAE-GffXeXeg_)a,.OZ5Z[3Pg[#]/94U<J>
^dE/C>G4.JL8,>7A_B>Ed&Ba?[)^P0WOU-\d?VEHe.-SPRQU].USF,8C)V./XA?>
8R2>ZLROf73TO:=7f.O?_bg3_Q4S<_AZ5HK>6Y96g:7SM)PXR4ZLB0,-YQ4?1K76
EY#aVC^C<[7)=OO5:,9-Mf.+a[IULOGZNd7VUC?A7&bS?]YVCL\]<9&eKMGW_.X5
1?=4>N=afaVg)+E@J]9155a>7;aVce^RWUKE0=6>gab7TCK@CUY22gK(2b9971Cb
;+>9UL\N;bSQ9.NB7M-1NcC-D[0e&L&c;CL82\OV?.1)e.b_=6(,B1b&3B7[#>4Q
USbe\6P8fIL)/27@CX8dK+I:c\AGI0,7E.cA+Q&?>Ed>HIe0BOVeX6FJNJ1cOW8d
/2Q>/&R3-\Dg0#:OaGJIVT6F#)JP>@g\0PUb=R^.7]^839H,@:RDUW9Ya=3RJTBE
Ze_:Z:EP=CLHB5B=M<PYc7OD_K(EO1R.?3[8LFX\,<T#_\VH_cTP:Y^e(7]H_TR@
M4S[>U4:]N.SQS]U6DP[>M]?O5Y\/fWS2>S-WHD-76G^E(T3L=Y&7:GRA);GE(5#
L^E9BY>WEZP5I-59)YO[Q)DA8NM2#E=g</c0]G)aER<NPEK)XG;7f\@D,eVJ@T7H
KeU&UA0BH>8G:>6P#RcV^0\UQUKbA/C+b()/L.IV:XA]Q+]=A82_V@\Qd]KALZ=d
VLA^WL.3/K27=.^>.E?;c7X-3C4J5RdGS)OAKEVW0D1K^aTBC^\7;+97E.9a@#66
;fL;T,,TJKJDfLD9GYNP-g><PCeHAB>K>5VPcR23Hf37X8-b;)OdRVL=[=G0T5[_
O#17CYJ&H/;#OU0QYG.f;S:>>VcUM5R<:X;UD=VG5+:X.(.S(eXSD2b9e+g>+cf7
_7KSg[@M7eVOUC\KZ(1DPG]W\+7>+DE_&=.F@PCOIF7M->@L[8ALAK0L7)I?aJ>T
)/MH&g/9E[AENYD^^NX7e3UYY3&#g6NJDPbP57-Z\g4JCD4,Fc2A9[MdKA)10BdV
F9HQV@ARG\D3<]?[_-1#CZ#bJ+2;J(1IPe]N&&CDb\&)A6BVN2)^8K95<5;2HS;C
JA@D@(58>+FRO3A_S]43#9IK_Hc6e.CKN1NHFa?N&V<VC.E.DM-WM>I6b2@2bfXL
e.(0VL08IZ:J:L/27Sf#=P89Jf)X(N&0He86OcPFT&0<EA.HQ8V/VJXJ_dcI-+.^
abQd]LG_F/W]+,aGRg<+Y\5LJUg:\fRfdWfJ;#MA68^6VM\TR7.I_5)CG#6>J:Ud
/;gd[Sc9KD,0/J+]EgSU@c-#5f#?)XfaP2<2&1>:/_(5f?Qf:d4KYW8TM[>:.:][
6fNb)6S-#46a:&IZC,c>dOYbBD26^.N/7RCG_7DP5FDY_:/@UQ\CcWHb(aO]e95+
S\V^dIGV)[LFO0gfg1].^1;d75N):>f.MP8V2X:S_1e0G@Z-KOY#.)7Pd;CUd714
A6<37?IBTR&&[+7d9KJWZ7:L:IK]Ag09d7bU[6PX5\O90<8,Z8a@3@K18;F6V[dM
9;D<X.P/_N2MFT6-Y_X6R=V_b[N^B/\6..E6P>)(0,bQa/@B;BZbXA2a9DAc5MRH
-A+IF/+IM&[DV^XVNO&?89<fd?>JDBG[=P6UAZ5&LH,?&I@=R>eW(IfUYY51(FCd
FTODHeBEZKTK:2=.4P-9+70<S&;2g^Q3];BdePaM-D?&KKO#SI[@fE-.a#L<TF?>
)IQGAF4M<e&08&-P6NYS.Y8S6JdI.^>V7YP<9,Y@VY@)&NL(+4K@AEc8=;L+Z7..
[0RN<3?<Q>+8]f_UY?gH@Uc#C@)gZHK8GY59?U78,dDO2/F_-:UBMQGc]M2gbT0-
/M0MQ7(g&O&N]Lf;;.(d=[]-CM@T2PWA7H4#/7-0UVIC[(,=2#BF8Q#;EIcP(4K&
/5>,LET^E9>)@\e4M[C_@2]LFSM9BX/>IQE>gT884JRgL&c(C>(--INS,e3#3:dN
M:<_QDCA]T_a-W=5?a>c.X<JgD64NJ[94[(^/;1a4_6@PQ_,B4ZfgRXIGB2a[Ua[
C&9,B95Ha9_-1CD-<_I]I8GKAVW:b0K05I1<GR[9F&[6BK8&F]WD^<[M=bURg_:<
a[_Y/23=4PQfXL=aKe;]Z,O^EfG[((@Y1aHf(16GO,#;C17AQJ@EZaT\.g-XbCf0
O4D78ecN965]6;IL1224dL][R6-^&7OGb3)./)LP][O1K3bYd[)?\]U)53B1^D\T
MY,HYA11]-+2)VF.AC7(R<I=#L&RX/CJ_D_VQ(J3RWdO@b:<6\5d?#R#J_([M003
Z[HTc)UH8)TGFfLb[@KZ/+A]CNE>&T]E=-+gI>M<L#?LR@RH#dbB/\1a#f=2P7()
N5fA\Z#7QBa;=Z&Gc]KH4dQ&+(34#U=WF5c:,AQ(=#(WNQIWa3O[g(E&H0X8P8TN
I],-ZQPK5^YcYdM/(;[Y5S05;Y&CN)ZIKXWHc\L6U2RF9I\3.^V+(Y0=SQEL\T7S
3adf?&JU>dVU::AO7_][1fG)af]AbPa--PEX&Y^O8LC.\]0FN_UVS>VdCOWC,;?3
/-(bCHHc=K#FG++,ZT51#-79S=AHCfSfK#ZVQfA,IV0a]?3SS_D]]\5JF@SV_Ja_
e54gQ03PWMPAOgYNfD(^f#@IJcEOI0MN)]DR6S/UbD[9[8WK,6/9)YSb0Y72)7;L
)#V/_J9P&Dd0[Q)JDX4>:#aAU(M;1Xb>S<E_-(R9>@Z592LIZ2@AC2UO@C8/3K5,
T\)KO,KQ5d5dVZHFZ)?>M^5G&L4b6Ec2-#9LWDB/AGZEU:WCF+TS3+]g9Ag#EWdX
YE16NDdg4La.-F.>d)[G1K)M056\C\gYc7\:#S<[aA>I-cfGN7T1_@9D7SGRHT86
]W^U?UD[DQ(W;,XZES/K)6a<J1[XX5V@\E,D+Z:[CPG7D@V<Za5D[&-FC3\-KUR4
C2^=W6+V,PZA^4_K,?T19[)<;/57Y)E.P]1F>Jb5AQO3>F#VI01FFTM5:fHGJQIN
dXTK7?@f]KPO]\^(N:K<T;T#]F8IM0#MOF(U95[Q\90/\?RYWIRNN)H/d#2]HbP;
6Vd(<QM3>d\PS/M?[]EA@JN>IJUSK)[E7.#[)Y[.N@F1ccOA]B3#YCdZ@EJB>]&-
[POEE+[@dI.5IF?1Qf8G.RHg)P</8Sc7b47=bND@LN/<Q_TT[d?.A^I+8b<H\aRS
@<&#.O;e0.=?H1W-X04N(M\+I/JPICa;0FC&41I2TLC@,=:RbXYVTF0a:G<Q#JI1
A4WMSI@GF+H7Aag.b,6c=6A)/(H8R&LA0FES3S@.f#X(2b;+>L<T9#eE7XROGI)e
g]f1GWE(Ob+GL@V&UB9K_c\.H2,C:61:JBZ)gB/-=c(R47>ZUa(W/0Id,J&]305,
Z@<YL:D6,2:0VbWe.1ML#B4Qd8X-Me>5_-0:T?XEZD6L&d+4#YL<S-HZMc(ECKKN
fTbJC2PU4f2=X<IAM.-6FaYVR.Ba.Ga>8WcN&2RQK@I/Qe#FTYV#6Zda-VY>4UO7
W&Hb(8S@::83e/16bd?&f)<\9YXg?a4CE@914d;UA]4CJ)^V0\M5_cbQWH[aeA.I
&:FV19eA.9)IY=^8;fcSB]R-Ba=L]V6?R>[I]RDI^7[+I2J7:1a11:f&#&9FVM4D
HG@0EeJG@?]7N0(J>5O<MR.RUcg7YDV:dV5fK,LX60W\-^g5=)^M>E@9L<[/4]FO
MXfN/7Iaga\WL:LX#?ZN.[C3A>CV-<dO(/?=J##H1L#RMTFdK78=WTD3#ABJCfHV
2S,dSe&;aG&1bI4;dfCMK(-eS;29@Q+ID.]Mb7b#MbF]+(72OC=.039\DOMYC8[/
^2DS;WX-=>?7OBPAB=+75W5]91C@LXfM2gE&4F\+_0[/S+LNI=eS#=\Kc#2fSMJC
EQc?6X#CNX318>[W[9c[eS][]OE?=ag](ge\4>.\(+Q_-C=S6YK:?g(>N7gF)\3J
1(f@_6W\>4K#-,>fXYC<9X/b&=VO.>MYKXH1\^T>b6390+D4Kb)2LRPaa66f5SaC
=CLIO=be,&D0Mb?U5)]KDN#g/[0W]K[(b#<XGRf?RZQ/<>T>\WPD;5eO234\(-1]
M[([+S(_[@JG,A,<4<[)X(RO+]_<59\dHMY:>G5;4PPCAH(X()64_^:Y:(SS_Pa>
eB);&F,]DLc.EcO489/2I-G\PNB,(J7N/D+?f1[LI9QGG[M@JH-cAOF<CeKd^MNc
0Z[\.&g]-25g0BRRNdEM[J@/@W5f69)[CHIfQ9Eg9]K5[_Hed]3L\4Y#7Te\H,WG
Z4&I>ZTA7>5(WE:>3^7;LJX>C(XK:KUX2,Q/],M7VM14[J=<R1W6,_])1[2R.VKC
,gN@S+N\cY,)9X1YU&TD\c\RV\A_F0+CB]6&?bONfN\JZ-WR.IR7ILV3L5[PaTfb
,/^c@0A&:d<=gG7e:/ELDK7bJd4/ROXa;7EW+Rc.VV8PZV]<Sb>JA+D[Z_?/JE1P
V3IQT]K5#VI1?HHaeFV&G,^?_]2+2Q4b+(8ED3[G=PFF2.T?TYE=Jf6Y(@5\RIgV
-QO@5.)Y6bXY6eV#I-a=Xe((@M^O<3dNS]VfZ[37692D8gF>+)T^63)O]b#PD<,5
9D8,+ad5(NI^[FC6cN@e2>PaL-]4+Y]eYMQ#]JUc(#Md707f,XUPA;0?XX<3WMZd
#cSOGC1d@O3CEZ?8SQE2+bc/L0W0+1ZX#QL^-H/6Q2I(&&f9M&LJ.JXd6)QL[06g
IeE+AA;<&,=,7.c0=Wc&&@N@T8#+ec8&BGGIE;afK]g8eKTL\9UTLG-KWMD.;_-A
R0[+)Z1(NQ3f3C05e45eHEg3E8FYHd-bG?N_b8P<R4U7Q80FZg[=O,T2Z]bC6W;^
M>=4<T-MQ_R<&dM-D-(Wd+?gfXMMdMJH_FO<ET?gYVc4g\GF;_I@]DUC=<=a-+e[
3W5ON4KTN\dL(2?@+Y5CJe,F53[1@8?).4B6;&O9g29]Ug&(6+gZeN\R#;<JLPPZ
4-Y@C:[\5<Ga:W=dOPb6M[?AS+CB4NTc7S#AWfH37&3;O&+(3d6EGW(]WKHY/\1Z
Z[VLL(:a.N0D;W&PP8&WdZX;([LZ+H7F2f,01E0g?Ac)3<C2eH^;>3M6M?(S6&;D
^.dL[Z+T0XfaG>>bT8)9.@K^E0RH&PP7@ca[M217G:=TFUT8PQc)g=-ZZ8(UeM9H
7&YVOV/;L>QAYb?WF<Ra+6JNE2])gPDX/X9cIE-]UQSb4T&B9eXGU9?(ad-72+RL
I/1,]:W4<KK,+VW;/@9e11C+]Wb)LF]LF9Q9B?,(\=Z;A5[EPdd7>f4;e]E(JfJ@
9+\W0BKR8@Z;K[0)g]OW&C-dbE12eCcSdNTeY8TdVUI4-f58W@Qf)bEY0K1cc=>H
^-V6<dB_E0,Kf.@.KZ#X+f@Y42^)8?SdM.gOY1:7&H-].6_NA&O<f(KX:];<(E8e
+]M:4M0c.VE?gCC&,P+f]+TJJ78EMV^7&-7,C[?-R:;UEH#N\\V1<LC\N&TS&XDN
L>\NSbX0GU7>V2a:@-a2KP5YM^d#/I0CaccB],bF(g1VZ/N]NI8Pd]5E#Ec]8GGS
)fS0^3aT.dV--XORX,6^UR4ddI,bYH&/eCf1M1.cM<f=8#=M&BPFD/VP,&;#O+dX
;>ScLW<c4gEeWFGW-bQ@fR(<B+:BV1Qc1GA77)g2>DOY.G#&_>?BDdf1Y@F:K0)X
c?4HZS9N7@E;ILFGJ+E1Y8Y;(=g,4O4]HeLP9e/E8VcA8)&QcIU&;_Cg@066Fa?7
M=6O-G._BXL.CR:8J[VIV(1Y>>[-AQ&]5?0_M__WOdW?Qg2c<O/>(JTF^0Sg=]b?
Mb1gdBMAS9R2#N(JgJ&RN8.&CU@T,dD5A+g_c7^>?&c8Z[aC,24Gf_+a5RWJ8/.[
N02L@-,@@B+PYU_\f#T;OKI:D8b(@D+KX(4f-bODMD/Q]/8cP3OB(9KbY&H?4=#^
0+GLf6A/d63fGFAA/5d2)A0>S.6-NWPB.UJb2>V#84eV??N[5T1FLT+a-C/K/0NH
ddEV0(87_K064UA]YY-a(,[GO]^gI(:7g476=a.6fE/6VH?X7U22@HG/c1_0)F>H
:;J4:R9^;SeB<.C4@=IZf5-MGf0>Vf\\ORggg5S^@3TKY_#feUD-LPP\F4\9].NF
\E7TPL[_#5JY5be7;OXd#76J]MH[S5Ub]d88Q6SM]:O5-964R(&Z8Ged,DU^)Kc5
2F7F^gUfa^c9Tb@.FKS@bfbKaZCb^5XM<4QI?Y-E-D.P3e)L27SE3VO(-6e[GRN:
,@-]N,J(g+]5K;N-JaAHY[MW4)H<cER_<,+?V2P9B2BDTTMT6:?Te>@fFZ7Q<^0R
;+a@5J58=XDB>)#2NVaG/NUY+NgTa^bY?(#,c-_+UJ3BgfaN]gg#0:/C,5e_(WCP
PPTO=9+]=FgW80KZJ<BbMg88)R;RCZ3N<-DREa2_a8J]8VZF/I9]C=ZH0COBU\</
6_IN6a)1gHa\&6#T^3UKLeUV\.)dWP#Y:):Ff1>8(_8]_ee>RJO&X\/7XHT8aDA7
.eWVLQOJ?;c]fe_7K;A6WeBJ[.7B?Y[_HAX?1JZSBQQP/_HHVgOA#0?FCQ)\0U3I
,]XP/IUF2NV7?N,[\:](R5^QG^gK<(-Y<+=:M_b#]1c9a0V6SPCR:_:KD.YDN2bH
+IR9R9WCFD)Fa__88FCY-YeHdO^(HdCOS/;CX;DbO4<A>>:;0aC+;&W)Y)I=V\Ra
VX3[&SUZV=V(CLfL0<[]P988X_<#7Sef-#JVKE:WJIY)(N2bK[0H@[JB>Me[,MN8
@c54aG(EbZ\\GD&3.fLM0eV-@Q/2AKBX(gcH(22VK?XUc4)VdVNe^DNd<L048B&c
9fO<b;bR/9c==RQD#=d8\FROM_Yg\8U#Z@gcd9dS_)&[5=-c10&[+^5[./SH8cP.
R.Z/N^0K8#Gc&1//J&We9_ULTT=TZ=-J?&D+Pg:9_\JMHUB)POWcP_XI.O[.P.90
2^X4+M@TN]aL.NMQ+I4TV-E4]JA\]_S)be\],_.G5KIA9P9E_S^bO:[QKNZ5c@_-
g:H4>I<:#[EGHS<=EYTb\_f5^JY-HD??S<>IWg<E.-Y3D\V6]Ge3e]gW5ANRC>f,
GIS8W]ONHaDB1]d(U<_A(F9N/TT9S<_40V.]<bH>OJ6R??6TQYU]PI\.ZB\G,6LO
AgGN>e9f#:R^2]7cLdfFg.QRL>;HHCTL6dN\-;?Ea7HE\:C?21;.<_0M;5YbOLR6
[QBJT_K_R&b_XSUd[6HZ)R<#&EfM)-GX9DY(CbfVIPF/3c1QF;JPMS:K(P/2Wbgf
eS_^^g2UFYPadJ99f&_47b1#e4P@6F^e+N,R6AOWI60.25QZG]a(8]RE[M(1[_)[
K;Q4aERVUB05@LBT;.g99U0d:5.)2)M#<K-,75Yb.Vf41TST&f;aV/MB^=90K:9b
U#U(b+1XN^JYUVeY;4;KbOR:78JKeSgD[;;#/-LI6]AN<]CfRD2MWaDXUE@3S]<6
&/EQV^G5Wb=1eaOU2fBW4G?N[FVGMR9Dc8:?EP[D/.g0I-6B2XUV2gHEfgVa5<F4
#12K][e+TJcPQTUUC<]]P<MY_MOEL;_[b>Rf/S[PIefc@c9_VbBR5DD.e&[4.+2X
F=/1FgJ::J4,X9M0J[,RM;d(JC]aZX4&9K+:K0/PMAE9e2S.6U+MHGAF9@Kb[fGN
[^f1H^W_d,L?1MbXgL\+)Z+V(WKJ2Be1(4I6<5beJdJ[];.GO/e\/4J/?[&#Dd@,
1/HS0L<5T]KRc]>)G&\T_M/E/C8/LWQ3X3HKN(M80;dG9T.1_c@#9f^&;.O8ZD^d
\&JXbCT<=_QS=H5F5SUfASd5g#QLHfU>MU;YYIfG9b:@NW,e<62Y=XA7\GW@f^QT
QSA?-ERTT?QG6&4\E2ZLg-dTc#P2PVO^:PcV+ae)f]K8&H;1&S9_LQI+9J]I=.O5
Me.U8g\Eg=(,gdO05gP>b@^TN6(ad/SeA+@[(aSg@PT[16f<W@3e3GMKfFDID_CG
_0,cd1DV/F+NaPS/B@BBNJU:=ZU3Pa7ZUg08EG+)ZA/_bIc@N&a]J,c<3eH==,P_
<TO4.-d[QO>146ZO-0=eU/-M_.XY@>^EK&S)4dE=<YK0-2eQ;_;ZJ&KF>)d],eVT
MAOSZW4E-&B9;0,C1-bP;I<PKa+QXPK.-gL55COA(>WP6,cS(B:>&_XORZ3N<.KK
f:WM]DTR[RDIOUZ@\b66.?@<,eK:I38bSdR,9-YD<:YaXOANR)0-W=eDJES7#9/0
#&FeO+G2W]9)?LecES5RP9g:f9[[9XdZA0d&#0I+.MPQ_M9H]8T(F=WLU1RR06++
;TZD(E2]:>bI:&?0TBZSM<]/W/;^FeP#fT2+@SKe#<?I[__c>O89>b9XN<<;FY95
IFO#7/g,:T<?[1+B)9VdDdDLS(=@Hfd)5E7X/Q[)3cGS2#<W7U]7f0_<NI+c]USd
7Q7bV+K\B=eR)Q79]LF_dd\QcV-5]0U-&GIOH6Mb_:-J&)WbLX^OKR=:61a\WA-f
IYK,^Q@#Ra+Q/\]LfJB/N=#^,1V8X3SH4.\1[O3&KgC+.P2f/[_^aTGQ<Q(,;OI[
(edV41F9MD93CN\[LBG/G#G0aLDcGLfH^V7_L,>9=QIf,T2G7TQ&9^g6LZbc]T@g
a15FB+,f6e#Pf,gYIX-]XL6<=\]ZO20BS95W,c6\UNE<f@8ALa0WNTDLc<5dU;+e
_[YHOYBI.80gKYYb1LT:a_:^L0:,^E/A>Q1Z_6;FWcHR78/)&.S]P,20YZ.<)Z-g
?-@#]?#;SVA#.ReCR_:&L>?f&BdB-06<GWaABfLU@GLHL-,dDL1@e&bb7e+-W;80
TCU7]^<1IEZGEQGTLU1H\#C?fA_ag;XV4?@]0_I#Vb)/6dZ.KH=fD^\DE[&3T,d7
01;65(Uga>-_/6/WbOD)4HTeEW(I_ZW9(\E#A?+VCUNYa=P<&\K<HN^)<JYFfQS5
LI/=5e.S5c&c>>O76_7:fbJA2=+_X=4MCX[.d=UP4.\&G5]+F^G/S@=;OeS__a6d
T7@]4&gV@&6ITRM8IcCcII_ZRY2?Q>:XY^Ad:RE1+g:PEH:dYQMZK+5,VO#&R2a(
IEZ9-E7-3U5g#3[&CIUe)+I,AI-@)(9,-T/gg^@/@CCZ]G&Za9NU\(T+(E5HMFgV
53DG_@g[BBSHC+gfFZ9P[Ie4QH[YFJU:_44L?DEX)^g/#EQ_H<+PI,G?=SC03VO0
6D>H,EU0VY8D):acDN#?W_SGIK==?dTDda;3PM6[&2[[[UUQQAVM0_;J^U:)SR2K
NV.SbNXQ++)eJCFKAY@Y.H6YK)(>c.4EFb[.gTdQU9#RY?09-O6PbE@@/0d2#&?Q
eF@P4&W192R+#3Cg.@CM?N0TF@T[&L00)@?L7A0E:AMKg3(&DAdL35VR&LO:+)\+
AZ+<B5354-A<V793NB0@0SCA=AUK;S47DU7AJ#5._?U-?N/e&_bdOM7ba<U5KSBQ
T,;R[</#5TgKS09L&E2d8+F54/7Ta6G&1bf=GeL:?Z0WR=6_[c_.;RU5g<VXKgeM
]QA#MT1\McX:G<<5c?:-f5/=)Pc5PJYP#X2O4WVRH@:aE5Y^,b6aXG59NO2CfJ(-
O@E-Z<U]MKXA@c/JCVT88>a5F0<-FF=^=Y]G95-Y_?_Nc@U6K+6X0C[EGYN0^(EC
cZ(aX5Ze_JS/RaS^;3O)[cB2R.LeO5Ne,M)MaFg39[g=972Cg9OE@:63aDT1JbD1
L68,4(V,;8ZI@16,\B5+I40Sc9?8SV\NHAUTf>6a\^fI&QVBc&E9#Q+9=HZ6fVEL
P+U0JR=3&/D6L1NDP20LD0?K6ebc:A_K4@IY3<]--C00P+@0B5KH8@SKc]=VP8,K
8f\GZddFY&C3C75K.F?dRAMMf5RV#>/6W@3A:L\9OVHE&.XU[4\LT^7>GL]a=[^J
,J)fAZcG>1H[Wb,8^M:g3QJ:5:G@_L;WT^BN)DcQ6e]&aZ:1-,6W-=85\L7^\X9W
SH6Agagd669aFEP<CH?XS0C/f\ZU?U<RJQX.[6E?6TBB4FC1Od/=PR1bCSGZ:;E_
>P?QV1S-)g:0P5TRZ]7UD/G#P>=Q>cf\=)NWP4XW\;Q^(,ES8.X\>^BeDdBM9ff6
,Wf;EeI-a,g\[f)gdFF>>1ZM_cU3)J6H7.P_5/;BMPY]19]]VBAY>^XCI>cCB+0F
P0.,8eUX>Z)SVcO=Yca@N8_WGWV=:FO+,KccJ/=]fTc>2XQ.@fU0UK1-+]@J>^dU
W_^)Le.=3+(&E-R/UL3/2<R_],7X=TaF>V3PL:TFX&W2>L6@UE688<X]Af]/RVHC
)<O=YCL1,QI_;]8KYcWRb\1W8FZG:3RN)6KX+T4^TMS/bdEXQOE@&47O<AFSP886
B#W:++K1X/+;\BM+=S63FNZD/@RM5MY[]G./eGbPP@1:OTULZ/a:e[TF#)@S/:Uc
KfFW-C:,JbOaW\MN#1g91KO>5/><K_FXO^^ZX/U=?;AaF9PNZMA+IPV@IAQa+YG]
VYM-#W0)&a0KaFUDV-G06[TVeM4@I,7U<WLN3G,JMD@#<>FR\49;<A<0^XQE=;8R
0DBVg=f^f:#B<Xc)UC.G\BM2XN=VT#&-P@Cd3[S#N,cfPHNGaK5WQ/>6eH4SW)__
F1^10QZgcNS]7P]EBG8@<A:B)SK]ID]?ZXS2.Pef]L0WN4ffXQWd1c3AH7D3P7R6
_We5MNCa,U(/2W7fI3\3Mb-P5]M]6MW=6dCcFZ43f?5S3:VT5.c?QWOKJB\?;-DT
P#0@TZX2=ZJ\H4:UC//?I7X#O<)W6>Y;eP\#3@,,?:ZH8fVC#KDY;Q8:HF+.Vd>N
U90MN3DO,?&YK=AcNZgF&O^bQ,E28)/O_7(bG^U:H>H8UOWaXe1gfG3)3B967&W:
MYS1.cQE9O&+BJ,3/.Z[ecTD97.1gP5XUA@W9f108QPB?.&VT,J3HfMfYa+>8.@5
LJO6)[T4?.cKNe(&-]^cQN(P7#,g1MV<2e?AU>G)>./HX_)TMe3F2Ac&\+Q]aI/\
d:Z_O1DFTN&J1bQMTZWLYd,ceWYN-:TZc999FN&GK24<9D6:Q2g,(4JCZWV=74\1
2)S0=H6;g+TLeCD7).??+PZW#eL0F&_U1#3GfG]_^W55+@F\1EU8VVOE&3GgQ/,@
B9U>9B?RB.MfN<R,,f0X?EMKBdE5N^&DP9QFR#1g\cO?ER1;,MJJ=-E?KScM\AZM
dL,d2;V:F#K>8(L&-0e.LTF93[GQ1SfK1&_7Z]IL5-<Dd(:@/O:cMLV>WC+1H;B1
df7PU\EZB__=BWcfM?&>[W&FZ/-H>RfaV?:Q7cR97R>+:1YS9UY_MPN4aH?XZ]dP
6GE[PW24MD-Jf]>R(bH\&M<6KP=K3?Hf88J9T45<N)+1<?HS.f5,>VWL)S7I\U@-
TOHN.2&/,W/]fNMYfWHbgUDH=Y7C-6a)_4/VP?0c-I2YeYa>O:KAS_F8@;fX[0@Z
D0dFX?@XBD^44g>_S3JLHHKDg^YaD<XYBLeOU:J->a,DE&W?CE>a^5\()4cAX+RH
BfJK2@Q[Vb>H;DD7bR0NY^?N6ROaW>(S\4^>0e@YYGWCRA:\gNTGY1:e3E^bg&76
CB6XFQ]IK\F^X@g(R:_Rg^11-[UP+W#>^1fL[e6\d<<XE>Q//G0P#gK)@2=Z,Igd
5,=Q4D2D4=(QIGO#>]8DLdAR&V#[YcIRcfU)F^,V3[8M75G>5=4=gdF66>[8QCO9
A\YUCA>T/<dLM0W/U;ZX6J[JB)L,g1+;/264f+M=X3&Jg3Q/UNfF=1M[Z:]V62@d
JC/9d7XJEHL@9b_c<P+I,e:L0#TS;1SLCdZ+T3/_8JZC)0bH@N3b1L5b\EJ;K0f,
[VS](4dI[<b6Ne?2PJe?#R=);T(Z#NT\Mf5FEGY?MMXCU7VRcJ@RG6-0J[3+20d#
+]))UaW#,811DGf+GW[T:Pf^\X>@;,BeReNULG<DRD:e1dA342U>dAYRE9S.AC>f
]A=_-/4Vdg^\DE_.(?ISSQ-JaZ77UK[>c+WJFFJC(a)W:G+6b:cU#<OL9]^,BfG^
M@PH.XN/#82c5B<b1dO94T:.FW37RN2HDA9?[e]P28R,-]-C[<Ja_>S2JDOYFB-T
#9=ge_/50B.B\08Y3ET^.C0:NR_@e2Wf@\(6\Kd(KcVH5/ZUf<3Yda-_>/.\f0T]
)PC+=I5@&Sd18Sc0)TIa]/fZ_E(4BTT4((DNJ#D0RfZU:H3#H4EBRJQ9C>?bQ_A+
Ac[W&[9)8-@?R(7>VJ#X:6U2;Q7^+K:bMb6g0XS+?HLGa9]g\])52VgF2Rd\e57A
H3K@T1O)4NTQ:_V22aL:R1[8+N&b\)1.2E>@DKA_d46:6ZF>O2MI<gA:[5>A:^.&
K5++&V@?:GV.4>(P;LgbHXKJ0dG1SBP/JXB&Ma&,52T.9^g76RH-_0>J3M\FD03]
BS,\SGe?847VW,IIfaXa9HLETe116Z:.C_Y-#DdUWNN)=EXCb3/Z(4-4F5S75P3V
?dS;#W+?M5#9SDFOPKN\cURg(G>J/f=S\g3@Q)UWVF6XF->?>@:620AGO[6Z#RCC
)X(JO^VRddDNOH7OCJ]gZ(Ebe3?g6VYXZ[Q/5a?R/LWJdg.YdOC)6R@;.H]c3d\.
Q3?(UJ5dO&e)dW:6@bH60^CR2e?_aRN>.ZV[(,g1;+.DF_NCdJ[R):)[[BK2]H(g
-]dA5Q^UXa;+V[7MA_+Ig.=]T>3_AL].JD,^=AW^KEb/@L)9@WB\<?9#E;e_^&6D
b@TUKP.c4,HR591;7:7SfLM[64/D:J&,,SN&[D2<eGL3H49e77>H,1(_^MG1N4RX
+JC05ggW[RXB+C(:L1+KS0EU@TS8O7GBV6V>GO]PeZQR@\PT<-f]gZ^(eDK-g)TO
CCb7HQUXMHAQVC@[<FXZIPcGBF4IK,Td-0N4A]]FQGIJ-_-eGYA:B@3#L.RTPUS;
Q)eCgg^f+aI#Q51<R9[HTU)?47fA&8eTLM41ACE:<MV\7U:-KV6/;(8c,:SHf;a+
e>#W+&E(#Y2.WM\5/0[&F2DbJ5eU</:1g[3Qf8RK/PgU&VQd/P<<MXMWbJCYWCD<
X?LPU/WUZXU[HC8;A5[6JSgI7QF[1>C/XQPKCC/H784BgXGK:IL_\OS8_.-B5?QQ
_3RM]3b>AH?>I](Q0SMPe,Y70.c=(SgDfO8;XT6bKg(H=4;^XR_Z1(R)BKcU[NG5
&ZJ9+<7A.:g7GfNG&)ZYG^0OS3&De+3?RWSBFV:7f[C26?Hb&8@;)&1GLD+bb.Jg
T?TYgbd]-T&/D4gU#GEe7XcN6]cR/;aKF(U+#H?VVBWNJ69d2.[e)(:]99,38MKG
_:0Y:Jf66g.T\XYWgJKc4<X[b/6eb;=E@;H<c]9:b0][V=CJfX[=?@GR&<].;-4[
cAKAKU]8Z7d23M1\KBSP)\)FR@,K633M&LJ0F^.2/@A;,4_./Y6T#T:1&LFXE/NR
c&=c-,2SOVN8A6G:NO<7BXMVaC3DZBfg+>A)JHJa7KYXVB2Y;_(,_[Z9B72.\PJ^
CWS#eMP=^WcBP+U9[g3RNXLe1eC\]CY[=9CBMKcJT\]11JB?&]3cZJ41GBQAf@J,
2Z)Vd56+/88<B.42a507ZE.[d.AB6ad/aU_+EFU:PG=^+^7?Tb_@g4]S:aOFR,-a
Z=aO=_dbR3?^MP,fV<Ff&9/fOR37;F;eb,Q<J9G+#B+)_FFG)HBe4@GE4JSY^FM4
=5X4Qa+De.dAfB3?SU>FVPgUXW.M/E9Q-@G_\7Z52K);f_7I0f0AY(#2&?Mga^eV
P7)LVP@Q@#&RbP=WfJ6-cHEPPP32@M^]bGbHg<-+2\.>QDL,/(9a(/XP2=>HT;dA
2<G<CPI/?94\g+2=eWg1DWYIRP(OX/5YgL,B\Qdc.SHg2V[O[ANI6&NK=M]YUaQ?
G93.@5Ae3@aCg]=Ld-CFX3?T+D17[,b.=A.>;gCONEQ)9D[1c]eSFOb(KPF@>O#-
GU:C82e39,#OE\.U?62RQbJa-9g[7I)3(TbcP^]7.7Tc)>#W)=NY>da/#-:Hb>AC
[F>:-Xdbf?J(4-Z:bTcFAVOQYZNa:0,<\4/VK1W?7EG3Y0ZReJe_@UE9cX@4e[8C
PL2:QL+DX6(V4.7GZ9=LZS.>>JHOeVVXY?a2b7U>X]0?5(3<,+P5=>N:2:;Y[Y0\
[Ec)I1DDEB7SeD;]_/W@VfIRXA=]#5ZK>B0>;Df@7]=Dab1\)Z]PHBfg9>,9;X/E
8I]Z(H^?TgEeK2?(g8[eWd@^FFQL?1QEMW.F^4+>.(AU@,:9;,Q&FRT:,P>5O3aX
9T.ZS\[e:]Re@=M-:64ee4&6.5>,LE/4RLd1XIS\bRJ+e:U84P(\@7Z:ef^I0)PT
Z&DB;HP(55dS5:ESNF>#LG/UCcI?HbQKMW/QJSf<X)#M1:I-P4WB.B/0@H2#B2S<
\>=dd>G)S<^L+[7E,eEC:3RKXCd2N1@R@?+\PYT_4(;gH2X^05^Icf45a=J[_.<O
\U_B(Ac@KWH+b]Se=3&L]aa__\#;MJ7VES^+ZD+QCSA^T,R<0dKb:^;He#=Ud/^)
(@Z_MdU+A&D;KZYV.fMD_<X2a>L[;&1+:X355[aQeM(dV;]aX3<)Z8:BN\QT7H&U
UFg0bLTDS>?Z&A[-F0-eCQLD4I9<^B(Lfa:-@PR;Y[,U9b3c3-^:,(:_J70BV)8\
/H&;@H^[8e:1-7C[cOI.IQ1WOO1PSC0#G.^&f\C-B?94W:T7a<H;:)]IU1((JQ6V
gHFgK5C,C\XS8cEW?_(d--HZ<\0:VRK1KeFIf=W^L6GG>)6?6NZ-A<V;6#GA?U_3
5J97&(29E30f)bSU=bc?Y/UdP7&Sf-EV/V^Qb.H6Tg][Vd[7E<E;@5#OI+D7EP\L
Xe^C#+M.<.7,aGSZJ@YBVW(6.c08M@LY/U^<\];Pc:fN3:0M+5fWHL++MeIN6;#2
8^Z#=2SZWeI#(:#F>&?cMJaTgB.(_98QU4MeD+c<36K)UOd2RDOAJ>672:TE@2;g
_2._N&/(EB&S)JEg9?bFg\K03LX3(1<>bI>V@+=;_=+21<gGeO:A&;^Da8[BT.EH
MX^(-=aR,PKV_COb_K[;S,cR(T)+E<a6AUFcDbQW6@9\R6JGQP^\Ge1^Y3ME\f9F
#:LP]Y]Y@bV^9C67[0[&Y\D&ALD[-;dED\Q-g4X9;KJ4-L1ZVSXC?T:?fX5]L\1(
G@DYX2DbCB38MRPASKc5:RM/?-[c[2b_]:)D602fg>T+.L:]25JPe.dCZUY1FbAO
K^<I#+H;E\\O[-34gEZBWTJ^d?NYU-=1CDZ:5cCfD:;6OINW=+L+6:0Kc0WE38IJ
HGOCI<D51RR-5UG?D)>:2d5\CSb(d5A@4JaZPbK93e_J2/(Td#bEBRcS.SXY+c<I
&Z2R(,;_H9WcW<Y66VNH@efD/B)LCXR@\SRb7]HJJ>WcR8cNbRcdQGf9Ub=+e(#2
R5CF63TH\7Q/WdKdBZ;0<)#8bA&/J]<K16b[<Ge8F^b4YB/Q^JWC<C^J.S\O4AQ9
^]AE.5&80XdHCTXa)XOf3X(9P77^20K[BF5;(-7aM214K&0=&8/^?8;^aG>g&I,#
/RQ;4g:f2V/<U<aM,.DAH@CGfg.\XVJE/4P6X)F@YSU=L,5=gD[0#+_=[7DG3T0)
\TLFBf62D[_0R&0/=0CX=B=U8LBHDS?FGLa/8@K&LUBF9OEH7YT,?Q6S>=d41/(E
Y2Pee^O:+2N72(?17a&@J2XCg?#=^cNU=,fcYTSHafa5,\0d(PLC;a;@gSAB8PWR
1I^)#.FTGIaZMQ&82QM7MaMVID),TGfQ&[EQH<?S9SA,J:@LcL9[:AL&LR,RI_GR
:.WdaY,QS)8L75J5XEM?0@b,+7^YTPI8AOWB^W8(Ye,C<HZSEO>1d1HQ8Z;(7Pd<
+<_1C\L7d)DaGNZLGR88K<WXPbCPSI1;47dY>ca6@Ja-EF;66[fGFF3;aC>YF?OL
#C<DNg3,@dBVg35gaL#&F:O^=V\DGN&;HW;7b:C<R&W):E)_UWO,]/PVOLO2Se,M
;D9De?c?ADS3]R4)VF<(e5bTF+52d-)RbCcXfTg(EN5W/]\/CKY6,\Tf]_9UbUdZ
S7f@#g8Me&bD-f6TQ.@R&NKBT=COL9H[<gC)aJDS:<[;(Sb8b]:K1C.;eS7NXY-N
Y\RM<9Y4/c)b^&C2A\d:(7CgJSV]43V5-4IR?I3;P>(e-aL^N1084Ca)FU[@=@:8
,IN_gA7OY[4UT>ZH/GJ-1S_I&aL6KU(9SV2LaH)d>H&-[,HCL=+J=B[K<.Q0HM3L
.UB0RVI1>X?Xa:;F=8WF&&f2:P]]ZOS:LM:M/M&M4(_5[YZ:E7-QH^a2XY<a?d^X
<K764WY]a.G[eK3#2VAGIe/[dB>A1/^gWR:IN18PI)K>5@W3KS?7.IX)g)6de2gX
QKa(J8HYKJPV^9Ba7(c(MA^O4QJ5?:G/>Y\D+IQXQ];OcECS4A<YO]U]X-,WJJI\
]0[K2H^0=Qb25^)eNM<#Z1a3:]G/e?ReebZ]Y^=eGM)4MMb]cO,a27@L,[a&RM&5
35#(8Cc5dI,S4TRV((BVFZVe#PW5N)/-E1)DaaaJ:A/0geCVb5LR<HG9b[G^[,X^
?B?2L=ec;LUf>b[ECJQZPXD8ZGXR5E(=RYe,/\F=-:C7JXG/IT,@+DgGO1fV]1c(
U=1/GB285W/<,)5GZ:d3Ac\]^<Y4MPZeDLXJR0/AKeC2L[P_Mdf(RS=WPFS3#AgT
2C4\cQZ\1/Y_SQ>UV<e]=@2GC])DE^HSX10MAM>?DDJ]d20:VU^_8UgIEb@8.^U7
@728AJZf=(+c;^VIe)3/V]@O_&OUWc)R9]]5TZT@f(@3S37Y.S-/gM:#VeI3P2;8
6P:b-VaXDOJLIBf@-9W5TH23?Z6?Q<Eff()K[G8bE[YEfYPH/7J,OCDII98;Z38B
d2CY1U1YDDJ@-=M;T9;08@Sg5@X]==0=.&Ne2[<QfeE2U,5)53;EALBBfS]bS1fb
4]B#eRN)E)5KfP3cg6M-[N>1@HE^(OV42354_<V[Jce_UHTa(O3fT0GNK#9M),>M
?dF3;Nfe=WOO;@JLG8@OZMA)&Sd5GAF3#EFS^F#U>U:=/N83_Hb<(4.=8M#M4EJc
,,AN)U?UH<Lc^6dCa[^(7\_1-\:+]Q35^OA80L0JV),H3eQP:Z29^;+Vf^_FM0IS
9^c_;()<_S_A[1F,IC08M(>c0IIC6\KUYe(I#A]PZg@J:gcF9@M5;F1WJ\+e8aTf
40bf?-ER.L79S>F8C/E38TEbH?40OS2b:Vf#D80+7I99>7J.H>WOdg>Oe4LMcT0W
AP_:\@JU_471B1S9H7BQ&U1HNPS1-Y65_+fa;BOW4OZU=-I2(?SD(E5fS:c&GVFa
#ABUHXfQN#8MVX,46,58NA+\7#S5.U6Z<B(IJ)QYM<T_K>R<3b)Z1c)U1Mc177:U
_bU3bdCe.dK0Z1W,g^)Pgd)?,XY7@F(a+],UPd9)Q-GHg<Xe@BfJb5&5Cd(\QDZC
I0S6Fc#f5Z5bM>[D+e5^LS<6NRbX[_T/)0HRMZ3@;4H\5>A,Q^HIWCA]JC/^V=?#
M8SH[=P7R^H?>45BL(,#/>c;\Ma?1f/;I4b-f6&^4eTH0T\P^\B;.IMB4:+XfV3H
H9H9STEX2&g.@8bJN-Y8E(^R4a8eD:M-8C8g?AdQMf2@NKA>_eVG9^fN9UAO,&E?
=N^=SWVBU_&-GW[VH.CJAW&1K(.-G=^H70:dA>^W(E;1Cg_VROc@).B5J6H,9-WR
^dQH.,P3dF7?A+9J&5Q@Kc9W(ETB1G1cMHLE^^TWE6+.gfF6BM1/\DX_3IF#\)fD
N7I\X-?M@AfR&=.cI-KIFUI.\A>bI/J>AL0Xg[1O=5G?,GA^W?V7c39.?EaDP(:\
301YO\,8J=:X/9\8HM#JcSP?:H=7N1&Gg[9WS&c=QL/Q#Qg-:C#OL+3LJ9=MI^B;
A^g]b:W)V0+AUN@G#=Z+[^6DR_BaAcBQ7__a-72M\\bCdB;8>N1e^TY_W=MB1CFQ
0Z8@>3;N:J?Zg5a;PD61&f/#(6MF#]LeQ#5,Maed&aYM^U9[)1#FMZT4)0H>04QB
Y@[JZE&5#,_D@ITTOD9+QLWW]UCD6QC>adD.8BTcDaS98gV4A5;Qd;:GdC_If:\4
_BAYY,O,D&)-76S]/;8#YH^HQa<YI,6g7N@<bDB++9c\LKJ7XF@TaZ0R8DR=#Y(6
)12JV5ZS9IC/+.1KGN(529U;IbaaYd4C#GdI54;Lg/H&Q89=af)X>Z#Xd[)He1[5
[(&^[JfUS;8,ACFS0gT]5]-CI9+b,C#\SIbO(SYYC6OWN^0;T3d(#<G0LFa>G-P6
5,S?38aFb6bU6=Q27<OJ,1X_?6L#&EA&GYWb>..SgP\L49cLd\CQXEE/O@A(?I^;
)JQU__NA_R<B<aR3DOCQ=N1=G6L&-]db7FUKQ[SOX^C\\[?Q[#U>bX>.^BM.&16B
R/QRLUEgabdM&1R<79>V(>6E4+;J^\UNeC[WEfC3fR^[L_0X0LD/\NSC,36gB2&2
,b<_B\K@&G2g#[BC:C/TS-Y9U5VMY5g);CBQ>Jc^H?[XU4QX@d0CHb)W;U(YC\Qf
[0565=-#WJ5@48>C5,UFVc/4..?fP)DY,;I^B?6[-@WQbd^f+IdGb_VAZ2&(BOU=
[B4)SX.+g0]P42A?YeFUd?+A&1B#Q/2.W<&&N3aK\8]&CL2?60e12eZ@_-(SccMf
NN11RJSSW#EP4PJ:9OH+TVJIYKGb)&fGP9eUW/Xd^6,8-PBBDU9Y.D]IEBdcdU5Y
e6eI_6\f0P.JT:<1bSdMG.T4@HD2@NZM>^J5TR77RF2bV?3GD(#.+AS.E3;9&_:&
+JT.3gU@4:RO9?]<.\#X/,g4&e47_2[.XeSOF3_VX4=/Y_UAJ>\[VP7KYf#/BM5&
M@H6OLKfcXR6R#16G[IXN,#MCY,=[,V;,.R;4@KB3^?YgHXSCE;aO7-\J:/M,^TY
E5(:W8E6f1XQN0=K(Q5Q[UQC>c1WWYH:^NWIfZ@@N-9eI(]>LW74MZMRS2RDP)1I
eX;+<._]]?R#;N:^9@-6cdU^gLfLZ8bFdZNTe9;WLAWR6dV2-/Z4^>aIB;CMN#N^
7;df1_9MB@DXYSHSV&X)XG9Q\2Uf.)^aO?Gg6X,DKNR6-?Z6#)GK)LEBgB8;P9(e
3B;SN.+(X0SCCIMdN098R8F]a^SQ(MLG1OPeCe[7+98Q2d6N_WU3I+F#O]RK<(EF
^/&8EQ<)eNKUUM[IR2/CF+4J79)-N7C[(@#&-NK)=Hb388W(cF^4]5;+XJ:\b-&?
Q\4C+AD3dVUYAWIVACAE3,M(^2\B7AC,(#4WE3&g@#?]5fZ2>.ZCS.-CZ[BI,_Zd
2?-7dNd^B?5XV)/:R)22)_E9K3&T.S5]fOAKE4K@N@.6B-L0P66^K-<.@8Q#]QBD
4S9dE<I51a:O/&N6Z[6)>\L8=_g-P?2@YC]4Ya4A.&DH5FF>@/&d+T/4\RM4@2O8
Ig)DO87B<gF:B\^QYC(\<V,(#6?A_6PM&U(SC&TZ_KTYcZ-ZbO[W,RHDRZ:S5O\e
1W1=#OfWcCWRHG20=afOT]GcH6fc0J)gTEK4gN).B#L17.FJ:E?I_Pda@ZeCO>-R
F>E3:Sb>Z[G<c8Pg)8DSQP#?V0^JJ,SB@R+5M_b@abH=bO/\\V^&PHER-DKV+GCO
(1\3;?61=AS#e22gK[3YZ?.aPH73Ue=2]2;eCT3YZ&4#CFW=GN2/8>FXR69MaCC+
N;>HIKb/]3:,GVHBWS7=c;D#,3-?BeST@f&81;P>W4e&E#DcBd7-.>+Q/HNaEga:
A+9?<YE4?&\W>W.+<A&X,GL=02/^H9O>5/>4GTTQ47L_U3_;;bKRR2cIE27GE_J7
bS_>7=GHaNK=Zc3,aOZ(V51<TbMb3W\eMLQ>^c2(98\+RU83_\^52/fb/Xb;IPbK
=d.6]L2G97)E_TD[/H<\],FcAPSHdVQc^Xg]@&EDe^cO+;;NfLO7Ug/VN&QRT:U/
dH(4+C@;cdVDL^(4/;K?dHS)+L,T9ME@.d0[eQ<L/)L=(]5^_B=]Z@2FPXO:]RC#
P3Z9F8P8&X1;--_J?(7eX4MdLNQELJB(\.IYDJdC\KI^E>GL,/d;Qg.K?BP/7.<^
F.:0-U[?=-KL9)2^71(:J6b3>[F_/LBJERLB:<N8;V<S@N@2V\-/<@A?G=e72ZE-
ac1C3GLgHZR/_3)W&Y\_)&V=CCgY7<=)#47+B=Z2YC@>:a\?f^^8^Q(#P9e;ATCb
LaP1-TL4N.0(e^N[JE9<C1aJ?dPSIUg)[>V8FD.Ya28U:S=a8??Hc9A6X@OWKZN<
>;W9dAB@fg4a;R9T9bCX^ME/V)IO;gN5O2f#b-\B;NE\B-0_]IFR,@&@?J[&]b0/
>D?GZ.73@4g/5Y,+AVU#S,]FWF.&Yf?0WTRMc&-KQL)6B=W.K@4SPYB2=X28;=F2
B=FfI@?70gJeE8+HU7<g;&R9L9OdI]e0S,J3ER/Yb?WH,CA7X?/?F+0P/9[X3BUN
I;THD[11JLg0^8_F1([TOMD#S,79B=PO^RYDYPX&9;A0K/g]G7XA9E/)?,MZ.;Gc
I#]g7KOMaPf&C?\.JHYa)VRD7#)cegPS/Ua#<ON[L6XEQE+R[e>E+)O]F7#A[0-F
/AZ=Y92gD4b@B(=;U07MG(I?.f.D>E;eKaNQSbXQ)7TU3-H&:MR)Y0YU:b@XB]OA
=B>X?)g[>d.G;fCR&NSG=M#8(4e;&&Lg0XOeWEb-6\I>.6a7A#83Wa[/-?)IZZJR
eFgFFN5BB1\G,b91HbQ]Gfe6O,>VH80-[9C9+E)ZHGS/#Q5X^^R:RI#K1#V_Ece?
b1SJ]]A^)3MEN\Y&59aB8B-9:<cZU#35(Ug;3aSI\.0?1,RP\NZ5)Y>9]7K^a+T]
SGUdQ&24PfcE2/CdIKNTNUYT2O_IIe7?:.,IJ60HW.DS)E.7&gFMU_fDc7#P>H50
?Q/_fK_B0-<bc9FA=Z^-O>^5eGbWJ4I)N;/3)_E,dTU,I,;+,3Q+U70fT<.WS\6_
VSV7IPU[)A8CL>c.;<7ES<9YBC/KJ2H#cARTL\J&@1f&AY4(#LG#=4LDaN5Y>Q[e
40+A^JEVQS:&?g;6J;PLY\)(AZT-P+U\\d)FDecNS6H>](.N/P3M@IL1?56a2+RF
+F+5[TF<.5>^42GD+XM/gZ:#22YG=3,OZT)7S?I;=ef)Q:1GFD5,BTeJ4:3Kcg_-
d0S#/;Q6.Aeb(f4#_ACb=+\FYVbQ(X&+A7^^\.7g+bMPRA3ZWFc(QeU>+U,f35UO
N]9BCO[EZEK7/B-X>F_W\dgUa/WW<\Vd(-_+5X?Ze<(UDW#cXE#M;b+-eK?^T4I0
(EV?aM_03EMK?S+&X8Y(;6e&E1)_g]8GSRJ8TOSO:\2UJ068\A\E974dBCP)d2)N
aRF@F)Qd=W?b>>TY/&d:C_Tfb?<KJ+HFKQQJYS532:KL6SVKHG:P;1)7X1>/.@@G
dA+&K-c?2MZ>]WG/;RKODU53:EeFNL)[[^F62X<SH?JE0FVI/\;F[NT51/[H:3.4
NQbTL26@)2F&e=U#]Ke/)cc)g\RTBFRA8R>_<7W,4_M>9^9PI0:&DB1;9:#&XVMT
bZOJDW>IFT3@:Y(220eB:PI8eM>(-YP\[:eJ4OCaAOJ3H;C(Q8/+))?]I=+DDD,I
Z41C6bJSZQ?S;_DV7PHJd:>GM)@Q@(#2B5MCR+WJE0&^ZYdKeICN<32F+Qc5(:TA
6>WC63gaCZ5)Uc[Q,gF3eY(^/Q<^5Bf3f>Ne-X:DJS./J51.L0[<=93d;NDbAPfJ
[cTgX6SefOIF8D#gYZW4+LQ\4[X\R)X@_f^7MC6M:;HJ[/#I&&+GP-HO#08aaH>]
S]H2G#05@[^:gH#-,;I.KYG-G4?>.P?1IM(PC(AL/BRMBEZ?dJ]L,B;c5Y5R&Pgd
g59VfJ5.#3I\CU.HFG:,8:85T,;QOgN0\C,(+<BW3^VB]DI7gFDHTZNAU?A;YgOf
QWPM]GS]MXeZVJGfeLR<f>K=gJQHV+M,PCU>Y(a/X;@^cIJPD#B,N/W.MJZ5O:60
eYRM&8\4GOgB_aVC5H,Pg#L+0(Z(-^J]L870T5Y5)a.A--3(X7Q_KKdJZ:X9AYW9
B.NCYVWE_@SOc5@[B8gRMb>A+N#2&?JR+K4#,?RY=L6F[.(e=,W4K.cMS-V2ZF2V
6ECXS=4\J)+T>J-1:.PFQa]Z_[]F+P5BI8\(S9>IBLg6M:]U6@Qe()1bf8-V/E+9
^N,\[ML.9S&V>8?&ZJFGI0=@A4;82B)VF4dc<XEN(\_c]H^4CA5T]gW3?JPE,+WO
1+;05Z=.EMacX]\d6:9V6BGU;W/,_ZMQEWGeUV7_QRD+&KHf<?HJQ<5_@RDK,W<+
V;UC@1Ob]TU.4<:E83O>0H,RR>(NPS4S:e8C;-:f)F7YD(KA7V48;D11U\C+dQ=U
&c53]fJ9_)UAEA-WP>C<Bb=bE+/J8>@bOV):#E#cSgbZbX=8BaAgB9);XO@W44WQ
](N@V1V#^Y)T^Q4^/Y^IB#)\L-CPRC]K1KP]eQ)FS3S>I<BPgc,K5JOI\Q;dR,/_
a81:NcIQ7O&-FL57+4EI<67<dTK)J,V3F;/XIA&:W3_==\L))>47WgQXc#&H8D4P
\3-gUH=E2.K0[U-:g;/4LP43&JQT8FQ3/1#X^GX<VVGL+Ng)]f&VL)>Z84g<[;.0
&-dQ37Q([0BF/<MH;K_LHE?:724G]>O?a3dK\]=e;N;Q^Wf@(;>:&@TV3TN#_IBB
bOXg,++YQS\XWc]^@Ea#dB<[#e=7cKYBfH^?:Y&;WUQ5JC2--DK4GO(4Z-V?>:#e
/8:VXW?=@7#XG[M2\a9,M4)?-4S3Tb_SPAKNQFfaYa/&JU3#PB\.34)C6_ge06L1
K;3gOUH&PY^/U@LaK4B3Tc\R1)Wa-M1g&@3JG=DT6P#fZA_)?K.OJbG2cY4_@/]9
P57Z/K-SXO#VH^bPA1([OMUY4Z31aOR@MST&/[?N-PS:WHM-X+0/ULT@C?<>bWL9
H19JH&UdWe0Z8C^D[LbJcc#Rd=(c_+5&AC3;Y7D_eCZB5-Bf7<43@JA<Na0?W52;
4.[Fg([6)1J#TY#ZKKGQUR@1V<WN?=[R+DIPP&[>]JVX?^e&XP7],.M@7fHKfCRc
NO9CP=K:SRE,&ILZQbL?BPc860YV>a.MXJX7ga7<KEJX7^e;bVC.;G(&T[0:dHfM
gH=X\)J7/P^1GT#]GE2K=4=d7,JgJ4U>FQM_e5P#V84V7Z>T)M?A5cP1b<Y:76UK
6CAP[J/VgXYOf1?3/G69.^IU&E,N[<2_-cX42BNQ[/dF@(+dLSRLcDJ(.N7[:9<Y
dU7^N5HCMQW+9d8ZQ2.\c-4VKN4=J.KQIXRBP^>R(NMF1\4+<#T7T<3D=fd2F6N^
9CGVV?M+D\aFYRGR0A(aCfDB=]E@cafYF)??N1ZIMaL3g:LcAJ)]]EP=d/aL:X=e
78FD]Yc2^VFSP@TRUCNCa>S;MC658eP&??7CL2)J-Z.)C[a.ID^d>fNUKB5(F>Uc
C&D0a38RH;9+H3fP?)c(95T4B(]Xfa^&<[FU5.(6H@W2&eRG3R9fK9-aCN0H2.T)
VLVH,(JYHA\c3YH+C.5[N_]PHFMb2eIK;2Y[U@A\bM@<<X[VX(YY4cDG4;JTE<[C
9V6;V23#QH=BG>Z;ET_gRb;V:<a&6@T/.c7U>>a[(8&@=fDV=\2+F0[=G)^Ee.PD
5;7;]XG\2&J\Y+;fO;5@Z:M5RLO:Vb^??IY)3GP=PYB<.UdNc>CUQ8RR3OR]WcU\
,0AXEP4&Y)KV..LgBCE_eHPdaL/U;IJ;_Hg[.M?#/..V4Da]Ve2DQW1T@2W1P&;Z
\<-+(2c+&K238ZRGd2+f3W8g5A8#R<UcWJ5dBV@\XG@A7#&]V&Na:=/VCGD-5?\&
?I\&H>9Z@R.?a+BaBHTKN\@K)YN,f_M<fR)XSgdZQ.(KX;_>Tg[.17aaMcK3Kcg\
dX_07#A=WBCM-.BVCMfeQHT2@-d5:2.)Z6(LdgLaO(QYf(?P2dLITTTdIK9(KD3P
^;;\NSaTD=>T/b1e]P(I8aNJ68N)&\gX8_[_QFS[8)2\ZWN33Z,_B8MaaT0/#4TT
#RT-><gD#IBS=US57:<^2-Z-3FHQU:T;_EU:OMPX3ae5SX_52HS^E&>9e67D?/9?
+:B7N9(X>MZ(UMI]9>N0RFgQL:SCcG?a=O6YCg/6Z)N-[1LY8+<K_N.(JI61K#)R
5+b<:16OW/J/fGJ&8?MNDN,O<0?)adWNDQMZ06?QFLQ(cB.>E\&;<;6-CI]26ZdA
PJ4[KKCMC,D78QT7>cAV.I9[O[I,LU&MRAL67AIZ-Q3+@f^=#L(TX[]c-)2H=dTZ
+<A,gI\eJg8e-[^.g@?6RT,]9<cMeC1[RaJ.A5V1K]Z?EK>_CPbP1S=aYU@X^(#Z
7<4(R9>/@E+==M9-_P3Eea-gb\L5XL1^6Z9.ZY:Z.#1X3<Q#W4<2KQd/^eXQUeNV
E_GBT+83>72]dP.Q;^PWOKd:aMGI]/fIFg\\:a9_<c&#)O^,C4?:<:).9VYZ4D3Z
32G2CUbTVZFgQ]S.bZ-JZ<R\DWP&9<FQb>0K@D6/791JV&<F[0D7DfX(;ZcEb_(-
0)7V)MUaR<ZY8\CcP4E?F\PE)8=f//1KdCK03?XYK#+VRdYBX@V8BK7Ud&ST.IRA
Q&Ug<L/3=/[C;,c2;eM4DF@OY]TOe6D8=e5G[Pg,QUNBc[Q7Q;d0<G,MANAc]_)6
:.K^U_a/Q>E?_7YLc0ZC.ZK^Y,A.4A=/)2O:B.M?:BICa.b@(GS><1KLRNdP,#PZ
9eU>Q01YJ[F7R/dOEKa)?H6JU=T52)E:K4b2^/3&7WRGY=,=b^GG#__Q#5\)GPbO
P^-]b+;]=BFg\XC-a(MX71EBPFZ32;d9g.Ne2U]eVU?GR+P;PF\V]MQ9MD&;B1/)
:E4#IHOW&OERaL2ZGL_U,-b//J_H;OEPe39IDI\;<P+)<8Rbf9YO#N-G0_@\I;@U
J99U;<SR@[;JQ3T02#RCU^XH.\]R,A65T0b[E6K8P)Z]2IHD&S>>QG4(UN&Ug74S
=4Y>2IHVI(/CbZ5THgLL?[YC^3(]=e<0:b]XY/gWVQ+JN)9Fe\AX#T(DENC.F>)V
[fcE5KUU2-+MOR0SHZ.63.TbFE&LedJDZE^b+<<WSf#CdDU:76fd3_cQK?2cd.@A
-GD5DD@DAa7b,>WW>L<+D[AW2?C/a#WEM\caCU#8B\Q<XFgUXa1/O>F(SR)FURRL
@BMQ05O]L9FWdK(\fXc3dZ9a7QD:1eW^07+]PYOH9aSO5V\G)=K_U9-K_;0Q,ge<
&X5\Kb&EZ^/:fG^5dIS:_LgY0#<6gT?8XXTTIS,KNb(PXJXR4??&aWf1,W8)T\Jb
KV6fW;cUXZ_/GbdHJ?3<0A9L7K.XDT11I>MP-VG,+g[LHDNHV-K4e]_DNF(E<c5M
GMP4Q__>Y(+5L?P6)2[5e2Y38SH<JaIbbJA<L+RF+NXCO(9\>S0RB5RFY21ENDN9
YLT>=^G;;MeRX3C[)P-]3/ZB.)_JKc#&Dce:X?-F.70X4;AfH#5QNbFHE<3?A+&8
f,.F&D&I)cT54eK17:(HH(INVY&1D>O(]Qe)dg,AKW,+\]\?>W3-51RT?fgbg6>^
4)3gVD:Id/1K;e[aUAb)IN]EX(V&;?30_GbFB2:SL19J/K@V=U]+=UbK>4_HK:.&
<#=0V=a_S;Ked8<CZgRN^g^O7#He7,^R&JHQ6-68\=d?/BC@G2F[HgE&M5NV728@
HXcX_SJcB@7ZXf&TTEXC^4[1b5_JTgIY-TLQLF(PP4&^T.?T)HRb3L.M&#E0=b>&
(gF.#[MZF)R;48\P:f)<O,KE5;2HF^ZK5HK^5QaJ9dR&IJ.1XgBaCaRAS8&1c2D_
H=>,2)(<;(2T2a(RGSJ1?_<gb/77;O06S5^,_?H#(cI?+CKE52eS4:]W:V0Ld@LY
fKVV<=/1S53&KX46Y7()I@9AQ6K.c<AGZ=?L^KXUDCDM3W3+VGD6W73&>T057;60
SNXK\&=M>b>>&O>#PCVJ/]I37>D5cAD5YYD4]-,>,9=]SEcZFEfUFaQZV/1T&4L.
aG=,>D#H^5IF:M_,bS+6?R6AYORFc?ZF9;f@)BE[C2,/T(ZUEY@OWZ>5[;Hg5B\,
74CY1^#KCW(OCS>;Vfa8@gPaPDDJ?T\J_S4Wg[c>)2?@R2>I9Xf@/eV7XMX@7_N+
0+9F@7Ygb&9Fe4H,:0,-#&OFR)BR30(#LMc3VA4H7ecWNI&/Sd&Rf8V7ZH#]TPb_
Z7cY/Q@ad-?O[4;,)6ON[QYF^96.83c)]d,IG0?)7d#4CUV,\86EP+W&./)Nef1J
6N_4)P3cb)3K&c/3ff\SQ2^:\F]L@-TBPI/H@#]>E]MBI.K#MD=@H5,M^PPf,-NT
=6GD]J.B=/f,,-SG6fgG844;3?FS1:6OJD\.[g)HEFK0b+?HMF=ZKJ,GNS^)eIP&
<eK[R=,N.GP7/;d&6UF/YDSS+=Y=GeC@]0<^AgB=&PU1Z8@S#c/J+[:_OA08[IfK
ag18&=4.8=<Z>[X+?@(Z2NR:?1HAE.V-UVF-\V,Jg]W+PM2QB44.AB(SJdB,6Vd8
8_]9:-A]bIZ6M+K;f5AScWST>fd43N<=CM?<HX;2L]bQPf/A3Z]_Z>-R23(,;>(R
P,E/=(Y^;U?6W/O+Ca6aP4N/B8e3E;+MB;#6,KP==1,_g,GBC2]e)B+>9YJH1O.J
Eb1EDU1gQMCb]Qd.?M4Y[T?-K/_c9JH:F.+<S\TN3PHGTL7<=X>\KTCe2YaHZ3^V
Cb8\c72f;U>CQe[XMO(4160&V[Z^27M_J48U0UYP7<^T?8fI8+(_<MMHdB:6GdaL
-RVXa]\@WCUP2)&FK8=Q#\H?+BTcS2IeN?1H(e1>OEFDS(:60&dTC7P0@JM-J^IT
^=DbS).YT9/UdWf6^HU>:Z6HY^9SM,/OP1C,GR^S4Q__g3cWJ4^bMCE#X;c)Sf:L
I(/=&NRHf-D4RcbT_QV,5_U_)[D&Oa^.K/J4^?8\B35aSF(YYCI&BGgKF4(A>0N^
OB5^fXg:EIgdTea39O&U:BE@RLbNRVM-dQ9&NN)Q5,H,?&S?5L\\HTG0[Q<e0K>O
g-SXR_\@+B@,2.3b1;6E/GY14#fB700#F]^FU+S+A_JET,I-48fMBc/&\VK&XPX5
QL_3&E[b&d?2c&X_BE#2MLS&+HUJ68g<eXG&6cJ5e?AFY<E1WSQL?b=]A70.HaS3
770^U&K([Y_bd78,:7e01QgOT>>1K=LT8IY@M^?QVaR^Y2Q<Mg6\>JJYTX8,Cb4R
a0)I?Q6\;[X_O#/Pf6\8E.QA=M?Zb4?g=15NJT>A65N;F\A@bH@Z;EBLYd;K[bRN
WUg_<7(N.La4a&@D?=YdeY[3cDS/d:eC3YB73g)WR1e<GBb?QD(WKC2MSM?+&765
^A)F,R;Kb?_gb=[L2S\\@&,9EUYd/6\^X.8[B@e951g5dTF]GV=_:gbCHZM/48Bc
;QM:F=PT0;>ETI13C1DC@-9)E=>eNd9&A/431HKO<,bL3Ec8b\&Ze2@B:3C#LLML
KB:ePVcUK#=&F6g)4LU2#X:]#gGL8;O[a#P>ER&VAT;FZ0A38S&/1cS&#\B[8-=F
XMJ=7QQHCILM5^edG:<(\5@adXNTbH.EYZS\1O>@+()SPQEKg&#3G/KJ,TPMBO_+
FGgH,J[#MHWe_=B:2+<7b\_NQ9gM[.eQ:&)<TD+@cJ,5T6M>^c]5ae>2@T2Q&]<a
KT^Gc7+ObK>G11e.[ObA73+#()YU&&]D9.LSgdZ^,A1,C:MXQHZWd9Y]U2<Dc-7g
7Q[B68ATLM2Jf50OHSF(MW86^:=]SJR&D@;=P<&F@W8<5)19)eV,FYR=_AgB0]D@
#>@75-Q_LAcU;G<5E22((HEC73GQ8Y,MTfB&BM.&0&Wb33gL31<g&.cPCcVe2)KC
,;BLP_/ab2UcBS=)D8H#W+V&8CgX;6L8H6B?HZZ0.af257,Of+Z@gND)RKZR/U>1
?NS0eDE.NPCN7L;A],ed>42R1IXX3B<QUJgN&)6fW-<=;I+<2:8/\?/X]eYY&P,G
D)>=KcIOTJ(=gE70^X<JdYB;?cb+&Q_FCfgCGJ4IPP#RSDJEXJJO-Y5-<W62dY=g
>K#WTa5S^.Z:WVE,2W:UW5V[a-aQ(NKT/&N\GdA#O<WRgE,I/5I<<(TO#_Sf0L@4
S4X-eBWdOEC#ZF)EC/C&Y]G2FWASBMVH[e0_-PS;]A<EabV7bYSG<da1;U>cLUfc
UUA\R9M[O6LXLc.IZ@];27R()N4PH=X&6OMT_-?GL9>:/IO(\KA-Hf[2SNaC)f;[
Q2eSL^W?W&+>c;YU8JI/Xd8g)AJV;JdcL+.V\O_T::=DW2[FOKd<E(dbR(I:e&M:
VOZ@13F>88[;IJ?[YI57IK9#K<c<SPfPNMK<#Eg--:@UA5-<)YI?30\.<KFO.B^Q
N>f<1@PO5KC.Nc#.VBZFbSS-&_VIeX]A>&&0C=;R#+]I7d_;LGFJdJg^<0C5ZX)+
-(CO]HZJT\SW,#.-c7+HECY+O7A19VJ+44BeK\aN7.=-4aUe_f1?\a+4=MQ&8=?U
TKaMcDB)6WU)aLASM>L8&-J,C7JIcb:V:]A++?L^WbT&T@I8Q:ebJJ?AW/8?B7G0
^SDXXWX]<8b_S,[2Ag00<=FE]>G(==Q=:Z(?B8fHM&dMCWF+4VcgGVfTJF0+/ceA
5_O4c.X/FRaO/@S,KF#=#A;.N;_a\@T<CND@1MI2T<HEBB<Oc30#MWG67Kg^Z&IF
fdMeIQ7UY^Qc(<(KR.8\[?5@>MNc5I+51X0V^=TOZHOa.,GZ:C#3S-adB3EcFgHg
B^\,^DIDBSEY:3SV8_5H8e1E[TUBW&MGUZf)NU,21\5LZG1_CLQ3TBbEP<Z?#DCY
b>WY>-IHa;c6:;I00;DMLN6Y;-Z26?O+?C=dP4N.<&NI2@BL&TBAa4E]ONPWO]e:
CI&=N-+.LTO-bM\QR3Q&J<X<Q4)\V:bdZ4P=\\2NBcQB3b]/JBYPXZ=A?Z;9A+fB
YO@+Q2QT<0[/>^fLbF_T>43359U_Sf\&1Ug3/DfW<<Y\J<e[-CaH0FN5Y/Z#G3;A
g>MK(38ZeeF&OA.AO(\3M><WHGZC+6G^.],UgA//9P9db,=QP0.OA-C71G&P2e^@
S7VT9)5FA/35GOcQY889ZMJ8BdD@eK5cT-2.M_Qbdb4Qd112A^#6DW6T&]4@PZA]
-M;GCTB\0A.K65GSLQ6O-CeI:/I@G_R2Q.OIcPMBQ)ZE<2:J=Z/d=\d1Q>6?Mf?1
fS6UH9TZD[=E,A)I+^ZA2>[4=^W\N20c-@0YJKKTH5c&.&7^V7)Z\P:KA^gg@?HH
f3.#A3YE88&a.5/B-6ZE^)05:QB?-DA[.B8.9.c)bY&3T+?+6EAH#g.#8XR+LV3^
<CA.\PO1Lf69>?;1)acF0M,C;O\6Z#^_&cBC@._^J1aYf+F:;ORT^Tba1_H&KS3f
?:KE@P;dCQ_X>CbcRXg0\g(26P9SLJX4[TF]6D2A6dGX?44=#S_G.U.-9X&)^XeG
0gMJ#/>_/Uc4<6Z?.,@91-C3GBSXZ^2(GLOL?3\=B98V>E1:OaQ4GLXEDI5);d8(
#<1(MS706N@[KbVSCG;E7N/L>^a#-=T[eFJgf(4e<+(cf?EJ,U)dU3W[H\T+MSCQ
\+JHI8^gUeD^?+[UPRW.[C89_F.K^4Wb?@KG)a_^4;/cPfCA\,d65=H+#(Y/A_Z#
]WZg=WRJPa8<GZ?06XfL4,gAJ\d0SU<1)dYa)c41LNg1[-@I8?;Y7-_A^WL;JW;=
.C@[7eP8;X0WBE@bQ,^f&8=]QRf14g.92I5O5?^1bMO\ZgBGa>G+4RZMZ;B81gGO
HQg8M=>R1VCe5]EaZ7_]aXc70FK.,/,T:U]2/T[X+MAX_L_JP1I#J32\4A8/>P8E
KVPE0c]V1XJ<U,FffBJ)H8Z(-O4c?W,Q0<dV&YJ-Ua\NH0<<PAPOQXHRc5^:HMNW
55U.5\Ff,,O=Kf-J^QK+EANc3;QVLGQfC\c/6bZWE,E[:.DD2\IHBUA?=X3^>;Z8
=?U.QZa192Hb)IQbIL02D,9YCB,Z6?IGdOM&a,QD)ZUG#8Q)@P<+4\[C@]FE=IN=
#e3+W<MK1=2,aHI2E4OPgN.C>@O1O)f-J),3<>_B,9VAAK^UUT6PB^fX9&N9HDM.
L.D^3,@SXUN<aBgFeJ^JU3DfSXO_ZUO@HZ83Q2?P22We_gNU(98X/8MGgS3Z,bN@
fJK0R;&bGGT@5VVa)]Ib/e_:#OMeKP6.7#Y_V@Wg7a62EHR7F11N:H4EV2c4?9+&
c6dWDR@8g8L8e\.Z[STEJc^d:@=DMQgD?b28:L]+;#XK<@gc(Pg1R\^\bCQ#.77]
Q3+>\a6;H(H;JE>L\TaD<RW#4AVE9Z>\A.L31dGQ#.b\@,LWcKbEY;Nc+bL&Q^eP
N9eVc]gZ@cSQ6(.&3eOH<Q>b8PL<HKXLI#7WV8K^:3D&G&X[Ec/4HN[-4Y6RCVI=
A],??]II:d6b)D\,#CK?D-LI5I<@Ic]T=c&^fTVYNR#d-\WKHEfY=O>Oa(ga[6CV
Rb/0K+Bfaf,J+fJCQbd.\O2&\:<_6e6Y.@947.G/eV>CcTgcCJ+RP7DD<I-9;GBM
W;P<@-BNYb@;WWJR9L,bbYKf#aLeaFR(J&R\7Nf5K##O;DHWB;=/M5PQYW2\^>(0
Xc8aDZgd+[K9]-CUSHP&TC=M^fT;6[CY&Y<R[:fGBbTP2Z)SZB:(;Z-^SOF=F6d[
UVD1682)_(X;49_TQL1C5JQ5;BNJG-5BJg6?-^(.E3cPONFa\D7J[/<#Z07SO,a.
5_C\aQAHb=a#P?cS3/:I^R_eTL/\abUW;<3\50+.&70Qd,2:Od:a?JS6ZW;TD^[G
+6B][Za\/CH[X<2ePNP4\?UG3B]ae.@FE(NL6>43@(S>--O&<.)@)7^/g72QN[<>
Y+8g@Z89MBJCd8a>D.P<I<LOA)ZY_,I9BB\Z2.CE[/P[gI1-V=f5D>I:&P6U)?ZW
+E\-IVaLD#Acc)9ece@=b@f6ZGJNP][>PD53@U;M[;V:,WJ5<]R)GecL4]LS1@ZE
_M2^_FRfVaAYDJ#N2WDVGHf_?EUO:J.<>.,L_?0e77&Q7Y)N4A?0?F#?KbL5+:BW
C&9&]7=<.M/7,UYBANV9(_L:_P?VdQEPBH0>-]g&(F68P7Rbg?6FYf<]c<I=,IPA
5/,Q54(A8E+(E[B>=\RYgUB(Y2\+XZa+dX@F<LR:4_^F5]-ESKg=cN.4:CXD]=.F
?-1\6.5DAcCK[.RC4;0a[]c.f,>N>&GC:dW6H:W>BBY_<Vg>A:MSG<AD=-,B0WH<
f??5K>&a7IadfAY(4[.M)M7X5#.NZ0:;a5>SORHcWgbDWZRZBdf@ed:RV8=2:bK.
aPgX?e-??dVVcK+]&^ADU)X/K3N8\47SH_L8#7??PL[3eFX6/W3-e(&Y-&JS@PDS
g=[5LaW.L7CB>_U^1E?FWPW6U_e6J[N]:CXLU9ag_Q9e5QVI],_d@7@C2@43UUgI
LCZPX@Y_<6Wf/S.^YM;S&M[b=3K5U2S(>,2;R#[O./gG\-KFCdR4/D[(+:[?d<?3
L[-Mae39+Gf#<<L1.O-PAJB(<.Yb93NBC]XZ&A&^BD\&4_N7Y0Ffc3(/@YK7QbNA
2Ke0M#YOU;?93<8Xc6f.VO./FSCg,/P5B3VQ@3BHAY>@3[Sb-#)fF449FQSPI96/
EdJZ6LdZ[5>J9g5/QKJVb1EFZII5:>a27#_d.?<M7SBM@;f-)@W/RJ^?4+a)Fe(H
5W.DAbZ6.6Y=PH;=7De=>(?7ELX^9bTX9P]b,T?AFFW3V:\>CNd?=9.@+G]X767d
?Q^5?>A&>.:B,d4f?dSYLD0,JN]bT6+1+TQ^9gA@B,bBJg@@[CCD/<8\@BKAJ,dd
H)^GI.:B<0SPC)Ee#CS2-,\I6^#\]X-10^JJb^fVL1Qc3.eC6&OMbU(@9D/P<I01
>f^+Ag0IMAE8E57YS+ASP]^7MPU+O>A;22:-SEYb0,W::Y4(PQ52[XRD6</PK2VX
<BQ;=#0V6TWK1&g\V[Efc+6O:,g]8dQH2Pgc3W5>gM6,B[c?a[:9gL12ZQDSOI2:
P&9J</5_(<cLR??LQ=2^TKT]4E&,7g:<,5\_e>cJ&0V1G&LeU/,:H)0TAY]?/eTX
ABgX\[=PSS>^Fb=@Q:FGJ)CA5I<)2PF2;&K4D\UZDG6.3eWg(B1UHI?\#aXN?7DU
K&97+/>N1=P&TU4NQDRIXcR>S5\7QAO2:7R@GW9R&eJBKBES;WS0b&X202K8T]+@
EW&VUN>+_46Y,McH9,2&;KQZ],#2\/14&V4X,+-3aEM/fC3R^<4@I4?5U.7;44-4
R]EcJ#=/[c?6WW(#QfAX#()XZ8#\JXaWeMXf:T^48G<,WIZ5WNP[V]gbN:_7,)T\
Gcb7c<#AdHNXF0G(ZCCE8YNF;5=dEN(R)C>+^&KcAa+bG1J8N9N[T@,S,,WSF7,0
&\G#+DR(7JD&]g<(8>Pb.0:ccfM99W89X:dgF12QF_(I7\37)CYbaZUQU8P@ZQRV
Qd#/CRZad?C)XO1&?BO\fG#YefM[L:?IGe)8&N;C0E6F4<<Y6\R7PFEfB[I,?^0=
U[15)O-KR>1aK)fV1XeZcA?ce/GGR1Q_C&L1:g.H7cL.9=>aE(H.@SY)LM1(5OA_
1fd;@0Rf#;c/P7KDXA4f:81S2AKC89V0bGDDKP/5O0eC;.2]8OY#Q#EFC/E/YT4<
cMLS<\a7W2<)=/)P(+<Gc&+RVd-:2.<PEVQ+a1eA&X+<@(W?@ff7T[PU&<D@5V.&
YYCV9Y_I^S&gI\VB)G,6GE4)JK)\^Q^1b^I;BU:Ub\^G=HLY0XGMJO[VM<QDS5_E
#V9DHWJYG:OW]e0>:.dC7P-:_Ea6LFRI\)Q@5Q=X:;d2@N6e?6Z/>_<5QC;,6JPa
(YJC\TFUT>.+Q(U6=c3>Za,@@YR)Od<2]P7HGQC\ZX7P(Og_W7&29,IRGEP481W7
34eM74D^)Y:B<PX27T0@-Y8?0.0e(>?e:4D)P->G,4WB#SKg)CW3a11+6(/5Y5NX
K/;d#BN,]D:af^D&3_2W)/X3VeRW7?E/P_2/b1.G)R5a#Z1Q:OE@3T7H_I8F1^=6
GX0U0N].,[d;QH;F9,68)8NID)<L0S+0:+PI97#GP7UHW<=Q44SOD46_a8W.fKRS
A[Q:?A]:/GUIH)DO?NeS_9C]F,^UQM(#:,.O)#7gb2YJJ(:TI^(8WTE>_#XXOb-Y
;fBS_FTaa#V5#,Kf]U_FZagW&(Xcb:P-DOCV_F3,EY9abefK[]1.<+Z&TRX3b1&E
11V0-;RdVSBdZ=@\.(g4bCZ4A]4QE4U(X=^I9LM+-TNXeWWIK_/WH^dO<[=P&5dQ
=P)I;G]e5QKK8EOR,M>-fJ@CQ-+DB6[\+X#0A]AO235W)N<8D0;<Z0>NV-46=C:4
&V.D[;?7),EUNR#LO2X]A8F6Cf^3PTBL<c2Q590]GSFP0bI:,DSI3M&N(OLOGF/_
&>,048bDJ]E;6fbDMYegB\3ga2RO5^f6JSG\Y8:GUb]cZNfX83c@eLO<L7XAFc/M
2A)ZLc.F/ec)C,)UKc^dR>b;f>,\+Ad)5b8]7/g3^D<L7:5.:F[2Cc^,-7K,FHOH
GA[JURKKdN?SEJ6OOUXL^J^U57eV=IfVcda4)WJA;\^WV/3N87MJ,6&B79VN-WD/
;-T-PJHW;X(40MdQL#D-_B(CJe<Q-Be-_):L#(gKVaE0Z]Vf1,^R;U/=O4c4UJY0
_T\N4P3Q<1:0,MAIO#F?QN;2NWW-N&[4;.7b_7YGV4YZWR6IT)b0P12-0f1#NU2M
LHc=\MPUN@g#G/<,_93eIF3@F-a[G4T_N(L;8DI:Z+EJXL8.(#UP#eRc#Pf16_H4
QT/Ice#Z?Y(9T=d&8#A6#.e.#>];<#Q(GIPQ3[&/gH=K1?SIR/H589SI?=IJ:O7Y
6OGEO-7[)a2?4c=HRg4Q6Mg?(JU(,B;_P/7KHe5I>IU\Kb;-MN3OI-?)+^E9/(]a
>0BY:S3)(9)??[)MdY@A+,OUfLHTR(e4J>0aS-_TLEWZQ39T=H@>FOSZ01\b0@-d
D\f,,IEM\49529J&R/EG.gFZ9G(KFB@-:L<T?1bPI=5:>cOO4\JNEPSQ;]#BRQRW
BB&d)X(]#>]M]=Q;[W?GXU8aQOB4?5f1IbNX-ca&a.f:8Q[__B_Lb?fKH4L1bKE?
5HZ\<=HD_P,(3AR\+:XLR3KBS2ZVRH\;_Z97MX)CZ6MUXPN)a=8.LM/O);#Zb]QO
d_^>e?ZTX=baM)WecKH/IJ:<LHE1TC&I9RU48^9Y0=a=PUC(1[+C;DC0^,5@c;YR
J\1HeM\=IBGAcK6FC;\.bA9]:7edDDUZe9E5>ZMA>2MM5NA31bf<WD2Z[Je(_A(S
^Y,?4VEMVOTfJ7-0GI+&JHfcVVF-U,?&EBT9TXPGYe)+^GUEG^CT@4Q[])W7(g1D
AbUd,e\H.WBKbPZ#F(F;d<&>PRc6gVDHIM(W2;R9\c84b0K)@:f+[8UR&SUIF7O5
JHXE(M2-:#=42B;4L7WFU;g0N2T];5a7[+.[g#e<BVS]_]Q.OJI(@VWLBB<LHcc8
Y4-P:,@I)9(;:Wg(UPb2,ROB83[5FP(0(ZbDfLTMM_(+7-D.F8fZ6a)PANb_DY0J
=gF):X\RV>:05Na_\B?069QG83@[11F)K+_+SO4>OD+\,JW1;_[2M1RJN;[&M3W8
eEeIKKH[<8cFT\RC62.3DI#1JEW:)(?=?2Q@6I+&[LLSg8HHO(b_4fX?^6^6e3KG
_3\]edP?gDNK;W&P0E^cMOL7^&.T8NT+d9/80f1UU:4cSN[7DdC)\=Z(f?:1g4&-
L1+=:=P\M2WOcS.Hc2<)]_G5S;^)9_7fU/C#d\gQ737\6H(K8N&<Eag0EE&LOM__
?I7;Oc@aQ_VTd3OA4LO:G5UG?7P2EZWe1+@cVO6^3UGbPF2UV+bHN4XFF.gE7&YI
V[7S18]K\.aB,@OX8[,8TU\W&LdLR15Z:^&eZ=>7G/(ZHc_.3a]YKM[S0>Gbe<>)
3@H>bg=+aA0;C/9W9[dVA<3>eK6/g/5J(?^V]/LJ)UQ,BNM1d-LE:,cJX:bJ+5<5
CW?5_=_gZ;_0B-D4+cZLR0^fF:P.)[8QFK>^_>NEUYe=ZgFGg[1O+F^gT):[@@G5
_<1+&dNc_3&L.:C^A2+#0BITDD&S),Kg-7VYUG4Xg40J@TEM=b>TOAXHZ]8AHB)\
VHEF]20J.+=6c\0<+\UJb+_=P68g#=/>990.T[:FOD6(8RGT>N^E3]f==<aVR17]
f36-=DKLM@?Q/YGB&7:f7H5-E6Y/aPPcV9a0Bf,+MI^S@[]LMC&EWS5;B.S.K\a0
C>@9^=2_QN.@JS0cZSVI])0REEOHBO<cDJI[+HF9&bI@Y1Z[2UgUO?d3::XY1@U9
QXAQYf8BXY(F@3J29=bWfd5[Z@B,&W,d/cQcAc;G[OR7M]<#H9-/91K]#63VOTfd
#KYReCgFU2#cQ?B9\ZR-1P;DN)_f7B^XAOb^C?SM^V_\0E\PKE5Sb</>()T+@9@-
UaA0df:4fI_Nbd7)3-6SAHCE>Y@eX93[Q_([D-Ya#DMZKDI:.;HD3g>^2V37=gGE
ZgR,.I:2N3M-Ad);Q2.eC4dYJ84610PIWcf+FbcE8DY9G2c]>/XdHR/;gCG>P;=8
J4N95[+/O@2#T5H5&aIW^-Db)b9gTL1YUCVOYa0,&(080FDOK/2BDI;J+<VO9EEM
<U#<@S+9XLCg?,GT::_,c8.U5_,TU2&7)11aOa>A,J&N6<9bG>:+ZP(5SA4J&_Pe
c6TRAIX9^@VPZQ9]d-NO0?DeEV1d8T#4VfF.=-Ng]@Vdg8^S7?&4K3OYbXKH?/Of
Ug?b1OGZg\eN50fW6/:XIEWM;M@&6;)]F9PJG]Fa>bfbK=;T2-c42,C5,T(EW/=U
)\G?.Q(V1#DOg]A_6FR,1XL/.NAbaO:W5c[C]<Uf0PS#BQDA,Q5T3DS2df:EQ#KN
N1A(?P3P1QagB)OA^;>2&c(_741f/QP_\e_a>NVD:fd4__>_a^7d\,1LFbC#=]26
6Y1^L[M\@KT6b&K[+ggacZ3Z9I^6f^Y<)?OJJ,P3S^MW/7@cNDRa_J7^Y(/Ca8R9
+&?[?;HVC(\BV@?>c^;_Se[=_?OA7N5N_+[]4DD3.DdL[/dBLNCRCS:_RcIdTH6V
fYgVS:R1BRN7>FFM?GA7.O+MEZC;E5HM1,?E^EGFO)79->^b:664UY1>DTbJ+J7Q
5Q@g/+O\KC/@G[AADL+4SVC#BD.T]7J2OZLVIHdMI?=7I/&C.Q7)a6&].ZZ=1?5-
<A_,RUF2/?3_cC4/^;\P-?_#]BJCAIfUV&LWF<)HY[+?Z(A2-)2C+fL<:ES(A/J]
?F.d3ZRY3gDSE9>2ZFfS=,3fKSa<YPXc9.5gHQ)2bJRU.cUK&]P_530#D:_=_4G[
K9+?,\X(Te(UEF1HV/-O7fOO,QCS73^B\_,O]>H0]#)R#+JM;X+A[8ZL=O=)3EDR
E=T^0+X71@;3(EAL:.WMIXIRW<:T5D/77J/.JH3_:83-4<IGX/[..F/e@^L3HK&W
;V>HAMP@,TQ#dAN=(&.Z?7gd6\_P2MJaW&@Ob^a=gM.#=U2.2#PY@95T]\[,>=_I
7B7;#g&(4+VXUV+<MD&.L@/=b+KD^245Oc-6-]a4d;N)H^fIBPeYZ8RB(4&W^1=5
B=[<U_<EUO_RQM(=GK/@@1NbUX9XAa68g+OCZ<78NO9EU/7_AUT62US];1COPG:4
F--dID?dbTDbY0-,1RRg?3>V;=M=g4L<#;[..^>@R;&KbL0eg1U3_g1:0L]@eGW:
Q-3aYF5D@[UB\7UB4CKYD41W[5XZZ?9R0^>A[L8W#d70_/L2eCT:7TC=GG(5:[C\
,cM4L517XL=0dL^+G0d#I6#E&)&.b?cI>\@1\-_^835Ee0aG<)39-\-:0?1?A/Ra
HfNd=97U&L0,1M9F2]G,YaPI[[AG1H2XF:BdeL>d;7^__,cD7:eWbHBJ[Q6Q76U5
\?)CK?#7/_@(:UGfE)A0I09dK]L#3<AB\.@/15+>d)Nbb1BN2@VfLf7):^,^@\L^
POW66U=DQFL@OU\AVU_E+S^(O9c^NJbcD=QL\K(ME)==&D]db).(b:4#7#AHJYV]
U_4IV\9^JQYH49-:,-DWfBbS?;.a=9c@VG>VM>f\EY^#B9f_L?BT3Nc^#aQYa4]E
)32GZG8-6AXa5AV#E4X\.N.d7,]eaF.CgV/&+CZLI.V?VT8]@>b.BAS4BM,6\9K]
><+XYD^IZ?:6+Xf\YFUG05O^VK]C^&VfL7YPZR/)\.IfW<4P[MFK.SK:>+AI^DP:
2O?JYC_JTZ-Z2Kb?HMK>5^D/-P.a07]H:/.HF1B&=gEV,a+@N)&+GcH4X>bG[<TV
[#/BW.XZ6Rgc]/9)GY<S:9gR0GV/\;WYAZ/;3)D:g\B1L0)D_dE[Bfd^bcT(SG-/
DK4)RG_0QWbV2>_,b/Te,MV?88bSM>RZ_EdIG&>,^aZTca_H;+6.V4HLD/JOD/IO
1\AW0e(f#,)01I;4-\0C[=URY7EHMg6CB6M#g3V5dRfH6c6[=)+0&a+cfRDMFT48
4]FbSWAQYe=;O)/9)9_C+VXUHa[M2_/1=?&7,Qe5G\DYJgW7N?6DOJ<4&5C,IBf+
21NZd&PcF_U<][:a#QAR97>C&O)49eL1@I:a/N-N]5Lb,c&I)=[IGH.(+/cW<](0
W:=+7Q2.d2dJH).&[=P5e+#Z>U^T4X6gc2HbX8P_J/)a?E<WH<CM<1?:@U8;cO^&
XeLdC=\8@(>_Xc8MB/KOIK1UOA)Ue1(E]\F?;EeS3.>eHfX6f[2V.,Y,?Z1;4A&G
K4<0\#FAJd(2)_XJFc-A0NXD;TZYUOHaI^@6c_&SU=cOPf5M5b80:K1&+38fd+^J
g42Hb#?Z.f9+?,+0g70R(Jbg7P.DUJ=.&+2RH_B\6KDNYCBf@aGWDce[+,FLOaaM
[>-6Ia&Q0/_&:(@E\bE/;M2:Fa8,48BOT]&IWc,g9H/9+ZaDN.:#?J,(:;2e&UL=
aAf/S2GGI[3]BJ,2:B@H)cTe/H?4;bgZQ6^5)aG(3b_,Z/PO<,6d=AeMT347Mbe)
W5@YR&SNWUG2)6;9SX7G;J8O2<QCH0KN^0:#Q#&;AJE4_]0)1&^K:NH;3:J8Q&62
c[\Z@=27OH7WY7>0[;L?cX,P<RJ^<G@<^=C?eT@9g^23.;\D6L>T1X=U1G0840AP
a/+FLV@[#)<2I2=EL+cS;I(Ke/(]G+_c2[/cQb;5J+Q>aZ</4K-+XMINJS:9N2fF
WWcQ.]P31V98XaBS.&g681)FRZQ?XB-TdH326T)bf]L325gVI23Z,T:X_TPC)IT=
bFC?Z5c_a@b\TfAe4Cc33T>8Td+-+QB+F)A3FF/B_e&YcHb0M^b\9:6PfRF>PcQ(
E>?,&]EUaR8KP))L4HgNRK0>...7BT]61,(O9EEF5G^-2IHZN+<8BLFUG?V>Z2SG
Q+^d1.?\?R)_fU)eNAPD]\S+eZFbT\QfX.MUGMZS/;[1492>Ad.LE#H98+C=O]H;
g<7N(<8#A^g&]SNdgNe=gU4;aRWI@.5_Q7Mf>OU)egH+\0C4O]EAPS4I=@LVX1IT
=eA8=E@83@92fe8/DUPW\d?HaZ)3^0D8T)/eVUA]dWQG#2[g;A@:&U]FVMM,E,<M
RK&9(ZSJTD<eK+^M(V71DX3NYG#b/#?C27ES7c:MD@V\?>?.+\=6\>:]aO-KLQN)
YI=eB/TQd/Q_X94A4[DVcH@]X&YEYDJ0FIfQb&DC^P]dUYgEcF4UZ2L>A);LeG5#
VT8D#LZGR5@_cHEN6-]dcE,bf)[VWI;2?IU14>(1+Y<Vd)1ZVP>e->aA;DATA8+U
.GH9LP_))2GKNCJb#;#ddg/XAf)I&63dJ+LFYKIcYW.C=e<)dF1SX;ba+0.=:OI<
G&XN;QP@HZIQ=L#<,DJBLLegec=O#9+G]fB)7>N:/a;[0#XDI3V@eE:@>^8.8(#=
)G(;FK>RX8A/ADK)F9LSIA7;#PO0e6ECS0ACY(W@UG;QSSBV(G4dOOd^SUQ8dLGd
Y].f=&7.(JO0NMF&.(W2=BHDQUCW&8fZc+,PA4.VWB>;B^PRbI[,BC@d5HQ&J9_]
RI&^#,E7-bSJ^55982d?8_;N-B9Z9SMV(G6WG?G.g;IeL\CL:2G+23d;7D4_(0d+
GGb21@F5&TW:68G76b+FfAa:-NDCH9\+TG<=YcK(XOUQ8bfQFOPMfS&Q_PcH_Wb>
P;E4(I0?=U43S<<gPNfb];6F]4B\51(OG9F(2-F?X)#(-E[2b3>B;[^A.L_VVI)Y
b?@I(C/;5FV4A:/=H/ZgWKP7gHcH+Pb::[X13#;AWKCCT/>3dJdfgQD-H?/5&2#N
+HD7C=G6JFEPP&CMRERM=.(V:b0=4(Re[E6_D&FWP7XD]@TERDFa&YIc[TJ_WZfV
T9@A-(FD17J7:aD&@]5gBCd?e67OWP^?1MRMJGg_W2]4RB9-W::-,CO2H^5dH,;;
L@RPa?M:1&Y75VR?OMd3OLSQ8;?FKL,d]_=.ZL+3e>E(K?=/:M1A/[e@^L7J1WOM
Y(d:B-+K[TBcV?=/\X((WF.M.[8J,e#SabK+g+M:]De5E4NZM/+[SMI?KT[4G_e:
[U^@Q28.OTBcb>:@[/;4-gAHV7.^YA0GFb^aJ9adK:9YFHN48??b>.cYL18/d9DA
Se;R5HGK5BUJQ#F+L:&F6V?20&c-&/-R\9Ea1^\SUZZ94UPO3:#SYefW&];fOS]N
=UVa#D)0GM-KC-WK&#6I&a[LWOI8ggIBa38&.>0aJI=(5/fV>6SMTdQN5V7PKF90
EH<^>-(3c<K:(>1dd6)abc#WK?NJ1[=BdLD3O)BMM4+YL0,@J6]M.^8C=G<6G;)=
AGf7;-EbC43=Fg,c;e0Q.GO.V;a;>/G3&<[AS8K8fLW\+I)TSI2050/V1[>g@/,b
[b=V;2)RUAR-HCf)G^^RIAaGG\=^5[YgbG,F@Q8gD)2D&9P2>]4/1D+WTO6><Z_H
VgNP:^A[.7dO\MS/Y?_@=9@A)-:f8>PX07WHT+ef(1.,0d1FL:f_dY@^=BCJ<&Q]
fd[SDYNS9?__0ZbR#@beE=)OPFHODKZ5G-P/8+1>Fd,fe?[C-O#SS[g;M&8^3TfW
=U(Ce_W&+K#8WOD]&QZTWf/>[(C4^KEH-(CU2gKOAULHV4TX80#7Q>[?O4<:<B[@
FLd:RL8Q&6UdFQUX&>He5c0a-OL4YJ^f4X54I=QY&8C_D(.HO9EK#AP&M5O>W[W=
QYSG4_L:dR.]I<M[;3,dBGFD<946UH)(8Q>Lb/8JVGL&EDc))Tc1>))8CS&U8V[F
eSY25RA7/bH2_&KFN-RT(48g71O@K)K[\JRD9=_>PY0g9JRB6,#9=\+gCL.d/Bd;
-BG=Ug.OGG[=W37Q=8@(EK5D.DHadT;G]Rd/a[4I,2?57&]dAV#(;VcAA?+;<0.W
:+)F[]CN(,B5?HZXDIg].ZPWRSU8bO0QfB/f263IV&1+5I=EJ4-@WB#?3(??]<D\
,(d@M=.88HCBG)/G/1&VQVF8H3D9OE8A0,bCeAN61[.T<L?GV1Q(/&G(B8DgBH=-
ZXc8?KdVXCHHg8@RER3OGg8e\IOMZ1?G84(-E1\Ac0bC4F5SRR+I80LC.7N7U7^<
_8ZN>I#bb8(SOXAY,..UOYXdZYW7]IM7+FUA#?G9[(Ac+<beZ0NQ;>d,E7Na0?P<
4Bd#Od(8dO^K@16H0b)dc-)HU#F\Se:eE;a-UVZ-.;EASJGU?\TL&X:9M0Q_<RHg
L;?4W<J0YS#2&NE1bSYK]bFX)@]d@I:b7^A-N6ZCX5=aCQS0HSWB#KCI/N@WKZZ:
HIY:&STLK:W:(QH(L&K]XeDYW:bO^96#c7LV/W2(<dV>5C4e[C^-K9)W:Qg1>8D8
8+Y0ee.]RV]:c,#7)E4eSMA@L)<S#O]+4<.Q^BG#1d#JMRUUPKgTfbVRJMSGSOg:
Wfb-Ac(g-7_VNCgX+.7RVA;4&ZF8IT@5(Q\Hc4KDD\(53=63Z<gZc^Y(a?OHAQOT
d^,a^<1J,Q\I;(JM/I4a]F&H=63^2+,?,1fdI]e./,C,-_65.N;Ie:\Jg_\X-ET2
gW):-<P]EFcPON\X8;b<QZ762\<FQK&(=abNbg?8LV[N7K?/_PTCIM];,.\>c-_+
&H@Y\/L;GP4=LA?F/OHa]L>(bHYBEIQ6+@TULP::Y(P9gOcFMOTfb\HICNN(4Sg.
#N0KHBE.>\Z44JM?HOb#U2eORPA]N;AP=KGV\UU69f&ASeSG80\2S(40R#I3b:2T
V:6>PX_[I(6Tg44-gaeK:.VNO<aU?@WQZ]+#;69BWE/LP=2S#BI3FCHdPHcdWXQ-
-3==d44].:;G7>=I_)9d\;Ie@Yb^T/ZHM=O38>WSbT+d-3?_]-EeB8F>cQ4+b5UX
UR_2Gb[eA<bK4->g10CXV&0/K)ZG3.R8.&X-+[]WH_#cH(c52?I9#HC)&LCDdD7[
c<-]X+Ua1A(V76:&gF_?O^/VUK(M\TA,IJ.\28(4,2PIA:8&6-?YXJ:-)Yc&-IB5
KPM1=0L\=;2UMe3W=NT^&.YY#3:CM#c0&-N,cY>#)bVJ+:5T-X#INcX5C,]XO498
1.<J\-+c9d_0c1(V:Le/6J=BQdH#c9,R.P5)JZZAAfA@\PZ6,Y4M4,N98B4Z2Na2
TRbSc3[08:b=M&f)O@ebFS7;BEa79OcYO1^V5f[G?\I<S;YD=J_72^(-<H,LI(UO
.+8HC=8\E5(&912PZg[]gP/A<LV>;CCQg]Z2+Qf2/^gDbLc+_Lc?f:S68QJDU5&Y
2E-5eF.F)-(1^eWN,/EB]M0TLcI\ad)R_GO)N1GQ6HbX;?\90Ud^1/[>:LOd[3JF
1/fe3_3X-C3f>WP(+:;3X&IGD@R;M[@b/&Od]?5_9+a/4C,#=cfGXFL]E/F>@Q<D
CX/Y^>QNQPc/7:I]Tc)A/M^?)@S0#=>b[[A8N?A0-/JW8fV^4\BGgca<H\G;Ue?O
&#(GdE/[)GY5JH@7_N9#4E3+:8>H\RE^5Q?ITH1=H47R+,))4#0H];1(),DI:]Hd
QW/X8A>VZLEX#+0Tc7d\HSe64+6L;-C18)O7&P6J&4VV1-CV:?ROLV1E7Qe/16GX
&3UNe\DfU.dB1e(L<1\#/G;3dC4Ff<IQH@3TLg3CaD,:5\;N->.FIHE#L=AO(?IJ
J:2BMB<[L-ce0]75F+86W]>,?R/VA0;GJ^b5_T9^XGZ\.#NSFHO+SJ\+U9)0S[03
Y)d/2;H#U=FQS5?(bgZHdE.?6;&O??0+UF];2-@;IF/KY>).Q9+)>97(IX2-fLJP
+b_;_gYf7[8a#6DXQ3L9^U;PC[,T4GA]RNN7FEaM/Z#g=JVDFWGKA=+\SQ0M162#
7HK#[\[ZOCAXT\eP_Q:LUT:N<Y\KOf:e[&Q^I=VNS+CV>Z?KE<c3]-7caRUSQ3RC
:E2BAdCHQ&LD1PD<Kb_bU3<V:dB=Ie-_;J\/dMFD63(Fg;4-CV/Q(E909XSV&-)/
43R5#.C^@&;d9#Ra^)0ZF2A#2d7/-)(9T.#aA\Df_@4?:2XH0+L)a(Tf#AP=QO^5
4>B<D2JE6g7+(aC-@J)dD^UJ3Zb?Dd4(46f>J]&7BfdXc&&1.-]JgDADGcYSb1gU
])Z=^c]EbI\F6ZR>-W<>Qb\;NC?^QL#Jf]@g-fN8CN<]JYgKR0M8B5&0GKg=D)#8
E(36SLZ8\.d^#A\6[)gH?UXeYc8f-;1fa<_1-TI?g]]U9YR7)UQIOd@/UNSQ?bA;
^9&FYeMdeX77?@W#-50R4-H3^PAS@S)#3WS8DTN<\Te&Gg?U;#/-#5PBQ9W153_-
1bJ4&#HB=Z\^=J8W4JS=\><BQ(+&=GH(XLDN;ETD^T^O>10OLOeX;5>6HBc\=b\8
CX(@X8I2L-LPWJC8)b?a[D?18Y5ccf]NA1@_GY0,U_C@b09\,SQ[@G:72bfJIdMO
^Y>M]:[1M9:cYZAO<VDgI5K-UTJO:/<g,8WHYQ9#R[,4(YAZ;8f,TBOV@[Z<_Z4A
\U&J#S609eI2R6[dSHJ_Z^?5VJK=+21\:1Z_Ta,QL>[^X^HVB4S<(HT]AeR.e4X9
7@XI1#7S<EGPZf<:2TX9]fYXYeBBSW-RPI?__CX,@Ua1ed<K(5a&7#OCJBeA3c+@
3\INd^-c/4<]IOe/[?9):,LZ<E8bE_fN35Q/LZd/6AWISM>2<\H/Z;8,X7=V65W;
=a#BWL?87PZD&38(dRP-d-Yg\:&DCbXY?ESfU0C#U2S3-A.RJf9[G9+S1C2DWd,V
5^HPN4C+SU=[KbO1^LD/<.W2eKd582F[RCS.MUXQLM/)f<<]8[PXcPM+M5M=XW\E
aafS<&dJ?..LBKLQKb+ZKd/^4O+[FbD9IcGZV>CTfI;_IEe1(CHIEFQD3RZ[]]8F
2PIH(JXC5OYSREQ#2IZNZDb.2)W#W/6IcX#:ST.X]F)X<1E/E;?]]I-W[[<Ie=\B
OfJU&#=C7A-^ge118V>HKF,?+6MWF86^KW:C2VQ6(.8/X3)#XJYM5O1K+e,4FER,
c,9DT2U@<aEQJO=RSV(MdfF;\X[AT#3)F@Ff??74S6(DC.FJ(/Q/<=MQc)K>VKYL
CJ073NXD4-F6fAW/9.Ge#3,2B@J^KDc&VH_Bf]gCFOIPMJ0S,AYgNJ)c(M&PMIBW
WYIA,+BS=,,RG1G\_)F_ZHY>IP&/M[3e(BUEX_JW0;#WOgK4d3HU27G_9R=O8QD-
bUWCYD+O6=;#G,&HRdM33a3.Z7\V0_(1@2&(e=fae6:OD0A(U\Z)>:\&A-N\&:FD
0cN/-O/J#^E@@RX7b,<QB)RVRIa\9+Z(NffO?X4-3=_GI)b-0XWAg,80W;SZE^KS
\gV^^>b=0(P/5A=fDL>1MYC)+8XRB]]f-\XUg_C:IF;W?P+HDgg+)T[KY_ef+)&3
;7]21BB7=V3](W\./Vg@f8U,>SV,\<W[V.8G8>d/E]g4)d@F\D)UL?:LLb6S^,@-
BM:F.FX(7(U?21edbeP_30EebE9]MY&_]8[0L7R>#\>Hdc,2SdMY2EgXF(Q8,Y^H
:U9(4;K^46.MHTQ63^.-4L@.>O<VbTcVAF007O##H/-)PL\CJIK.7(@^3G-4<U@K
aO[[Z+>d50^9&)VE;X)Q7E-VV]<^R=>W3UJ/G63#a.+YY45g@K]8VDOAO-DDXX[d
KLG+AGCELUZ69,>M)^9Ac_PW?)SdaDF&K#Bb^gF.5MVbXPQJPN\BSH>Qa1Y50e3G
EVa.(,0a8^/W[c9_/]595+2WM?aS@dZ9gQ55,Lg^W1E.1g5WV],.(8HK+B)J(T)6
d:BH7XV;?DT?3MZFAOQ\B_^R1,)(IeK]UKE46]#X;(+dIgR<9fZHg>bWJ_TT&<2\
\?Sc;ad>XJ9:?(;CV\cTLP?SOEZZA9,YP\JGIa]?3;\a@MJ0+/:4#,Qd<?2V[)fJ
=3J?Z954W2\GHXA[GVLQ_?.77O3+RP\.?D,IZZ6J]]=YdG>0dXG7O9B?]>R+)AV<
](6e[>(),;E]1IU9.S\<4(/F>4P/MFDH-IIUf;30A7A]NTbWG8\QZG<gB,@D+aFM
E8TA1a2H8Y,IdRZ;P85V0b960-:YNEWEIgD]9#6)HB2P8ffSGYdJ&We^=V>9S3\:
N^&.9BL-bA<6;8Kf]^K6W/5QV,A2(D5HMg]EQJ6_,0D9Q4IA.3fA]3?G/P<f50f0
L@bW8GESKG0OMVd\=6<#IE@_4Dg8W3JX;E-G(X#_:&PLM](=X9<@C>45P.1YLR48
EUeSR_KG9L4.:X9&Jd)7Y9KaaBE[QH4\4d9TF2N],#>#U-WW2D^gONH,Za(^<^@9
=2Oe/FG>0dG01bC@#Tc3Y.0NH3TPT+,J#??fNd?JDWfS7&TS/)S?JSL\VED>&_7I
_1OOeb=-4d4PZZ)3O_@fXFe+@#,V,XacT.?<@N9EOGD^Jd\E?d2&K7>]-__Yd9<Y
7gZW(&.6&POX,eH#=1K+MKJ^WR5\D8-YPXaM^:1e9FHZ]KKH)PU<]W>AAFE97>LE
YJBeHQ0&V9>+)L#Q]3:#X[9780=Mb[R_5<#Lb^dgR(g2JMG9/7DV1BIH;gU7_]bL
WV&J1>F+S[X<daY2b@0SNUc\+I>=5B=BM+<&YFF(_PCdUJ4.++80NP3E\^bK_@61
5#@[HL_K2cR-JfOVBJ4;+,/_UA=\GF6D4<\4aLB,,P^C5MeFM^>?e-=eMAZ/I=RY
<Pg[Q/gYUdQ(3K6f+5gQ+P_AU1/=OdWWdf4._E:I>MH-6R<_/_WC/E&fEV\?J?6;
#Bc8CJcPU7?EY7K_QB0288c@-8X=PGLOC5Q13@#K&4c@ZR1:F4FG)2GQHB1G740c
bDK@3MPRdQT&,Cb+_NMW1[MY148CD>d;9W[JEcR//97d#/GAPHdA[+e06@]X7VOS
Pa1B4KDCQPN^BgFY#AG(E1B9Ua+5-9Dg8H:8G7&(GfH0ANI^NAGc]>Yf3&fR(+(c
XFK]_2TWHB:.5]ILQVRd70K<RYc(Bc0X;?JO8WC,5^LOHV5)K^Cf,]KMIGW67(K?
[)I:DGIb^0+c9f7W:8SZ0Q#P@d7IB2;Q697W;7+.S:HN-;^<ZF@g<RVE)UKb?&cH
@e-b+3^DJDE9N8\]]H2.IccYg^^MA26(OAL)BE_9GZ,bDC/HX4H+WW<<?U^=_QR[
M6>+ZL0B2fEObH09VB11OK15,Z>E0Wc]^J?:cD:C[IaFOG\+WB6D8WK4TE4\VUJ9
CfOP.>(.EdIX<<6F:(-8bYLf2_eFR/g,SO=fIdZVc4c?Z^XR5A+aUD_UCTSHJLO[
S2@8C41c#HV(GS@E-<?#g[JN[47X0\_2Q^f.6GFODLO1@P?;_C/a?(#Ib<02I5ad
.LSBe7gK\81P_DGHM.M@MSf6H(gF?b:cN@[-Y,CF02?X(FB@=VTEJ+=+,HA0BR16
bU:gdcfBBbFR]VCeZ&6Ia7-bVB]-XPKI7D9,,FYN>GfHPf&X7NQZI2EXD#TMZC)2
0eC:VXI-G]Qdd:5dIL8?D4_S_N4U7^/)7H(e9e@S],]_g1a#6I]<86[H&CGCLP22
MDd,(c;/47=NeR,D;LX,N03dJD3+P.8cYGJXAJA2_(-,VQaV_50aP1&^P@2.<J13
Y@3^KB6d](=)TTL(e3L64ANg,P@<Sg;,27,\J.LT_R8YJK(8X<FUY0cJe@VgI5AE
4NPQ9K.M>&/()OR:X=[W84Jf2DcQe._)T(]TS:,/JT0C<&R0I3_II=1V4ELGDbPd
G5M;>[aY9/MQDd^+dbg#Z)(@cC<b3#@\^<JIMIQWHd5edg?\QDAb58EN0>YABX;1
\GMJGI7FBW?_KPF2+_7;fL7(\6C3UI008#&NL++[??VIYIFPRN@:Bf9TADD)M>]6
11UgADg7RDD8RAA/AHEA/PD^9:<?/D1,E8N9A://9IO>+Tb@X,\4\E50@2-X;fUK
)O=Q.9BeWY0efT=7GCR(#EYGPJ=50A<S/:N@;+bT5QQ,<d^6bQS):J-MfM[EGYc0
7-c=NNQ[);8+.4_>0B99__Mc_QMHL1@a;IgL.b/JLS@D@L4-Q5#BFSB.M,gR-e2,
eJ;8)62.S2._61&QgfL-8KT9Md)fSO.7(F17?4.?gCG6&eV:.U>VdVQ?bJ?c9.(R
M&Xg:cY3K\O<@WNZe-b)0QA]^7.IN=XZA>JF)g4FI9\C?DCWX#HMN8Ee9ff)OT(P
>+:UM=GOH<\[ZgMa1g5:O)=-PARQ6HD#P&TTeC^GNAE-,<4H1-5-?0=;e;]e(2M1
F5Bc/#2(,+WI?IV04?>dN>aUH2CO:DMXeE6c>B&M#;OVA4^J@U4c@?ZT].g1)C2(
Z)6[:f2\;-B0G8FY)W:5HOC?JKRaHYM4I<eWd9)N1;F7CCebF2Y@S2^,W=3QL833
a58a?UHc:M1JHCHNO<<A]7IA.fQB/EI>)aD\S\1YLRGS&<]0dQ2K[E9O1I/Bb,WP
\>\>E@\/b^&BN>5\Ud1W-;08>IB-K^Gac(449#2+/4^YCE6E-VM-SC>BL=F&@AA8
U(W=,[_g=140RRVLDNcN)@Y&3PB7F9F&)U]/MN6JPg.Gd^6^b+U;P#FLK&UG\ZLN
WN[C\.74ZfZOW[5//FCKRWJb;;J/Z]CKb9?B]7-N^c?Oa1G9S;:AeJ/K3e]WRR.L
>QZP>TC)5A?<KP^IM>9T5NdP<G6O-0\/(>2ZY4O]#KD75(b\.QD(N)R8R+a0H-(Y
4Dc6[0^4D7]>,9/?PX3H.B/(gc:g5cPV(5[.2R]N\#G1WLDNNSEMQ++??)bY/\:X
7g/Y;b7J+X>BCGV28K/EO<eX?0[KK[B.+b:2O2K,=,XU0;c8;fVH#E2#_eF<]/12
O)e=826Z^H&47YOK3NLSN&/;L7G,@;WZ#6\?-91TKSZa44;=_LEE8T_,\@aX+A-@
A(=R=bC:_g^@<]b.]<&c51YY<;0Qeb2P:PTUfW>4#4:OfSEgA1a@ec=8\W)4FWRR
,4S6\Z1E/WbBHN[c6ZBQEC6CCQZ6+6X:_DfJW-YJ33_1^DBT5_<3)c^LT][EG&A5
D62UBRd;J1WV;DV\/eH=(^]?X3NC9(]HQ:AZ?B94Q9PO5;IeA?00+]7J2\.^)6=L
(,&\bQ6Y3AL17df[5JXR&QIL,XI1J5bZ3KRX+\BG+YFZ5X^:&]->#BB#/fD(10GJ
g]F>SO^ZTB3)/B:O:,<><4?XK26-^T?J==,[[5R#b<EMaTg1MV[3\OBD,M4JU?)0
P;0>-KdAg\:QDG@bTQa?3d/^;aVO0>Q8OA;86=II6AJN0S5U+64V96DKE0J>dJc0
V#>PWGZWe[+&ZSf[H_U;dd?HcbGKB-_aYL3?]E#cL?Db)@3FfQ/2.BMPg#N-9F/c
U_@5^TR7OaX8^&I9>TEVDO_+2+P1edfSRB_e0@>-GaB)g;W@a\Z/):@4M=bW)^O2
#++RHAK<_&e;e-cd;73YGa<PG0Mc(&&^9\19_4a:./V<=&YKAZJ=O4Eg^W.ET9FR
(KN)A?5F+1XT#,Y#AegUHXd1<ZJ==bC&g50/;B5O@4YG#2NYS9Y&\<<>LbLAH61>
,2c5aUU=>]aV4<DSG(2V0;/ce8b[,MB=,;>O,^R.a(VD=\,7J#([@)Q,U>,KN<W_
g4ceVW_?D9FFOT9[MO;Bf=VYOBd7DTUf9eF_KRaWI<4;T?c;Cc(6>/eY9f40I9RB
PHeEd&c6GOO07bWMLO,g@&15cdNV9gAa+c<9_)/B];Q4c)YF._fLP/=Xf+S;P<RJ
c(ca4/M47V9Ee=U/S=KGQY&0?U;VBNb&+dQM;gE2V)T&CFNX<1e:c#4/2?^fH+N,
.LNPb+P&-OB88TU[J-EI:<TbB1f_0=TaL3](L23PO^)FA.98VL&972(9+6&eFJe=
gF#eYCJfXf<:T2TSRfL8DaB#CW;60MIA,aA>@//]S1?P4(^VG?AAce#;@ERQC5b[
W+4#H@+D_YFGA-ZQ+HR4Ta8JgfT_GBV/7-70Z9JOP^?D(<,.0]E.N_XV/4L+)8Z5
@C.[c;0QQKdC1ZY-dQd=+L,/N&Ld==D&,9BV\2X@;.S@7:BM&0:ZB=Q5ce,a3I(d
JI)@CP4R2J)6425&S,[QG[#&ZK(Gd(YW@Z#7A8MM+d.#&YX.Y@;T28g0FWb7=[8&
-DS0Dc1X[>T7]Z@J:Y7gaC,_5a8J:3cFeE@bWeMJ8]Wg+d.:2CfL(?:6)(,2d@+Y
+c-:9JH4>GPI8]X08>:4J9<2<F4I;5TMV>Ocace;ISHV@?K(C:1#HEWB@Q9Hf,+O
ZMT7PA.XGB81_-F@KF2\PMf.IPcDJW\>?gDWVK7cV?F2+_ER:34HV?V4#W^-gFUe
GL^&O3-.dS?+6XKa]WCO]HKGMV@AgYTHD1([8+OV;NZ4KF8-V#b3.R3#=17)I;@A
O-2RG4OgUB^MQ@&@O7KKF;EM#^#R4=I2LQaSB\1DOTY7:.6KP7075fJHPT:BfLK>
Oa_b-&<IY)H(KH^cU[gcFVR:^>/.[\2E5#ZK:Q\<1a&DgXL;O-,E/b=F,^cNe33b
HdAc/.KD@?gH_1P37R^X(],La4e(&([DKg]\G+P_WOHS1K5-99FGM/1;(9CH#A^:
&eQOg#L0Y.9.;E127WWNca2>_N)0:IUO=-_V?ecBRL-[8_1>QAU9=U18+^69CaMH
OgDOMB1&=],OVaLLNN4;EbLK-ZE]S3]bN4IOYKTLfMbbg^c#[[ZG-Z^Mg4E?:)?+
W]>#[1P]VF19,14S^e6QOM07\E_+YXRC2[/\b:N>c_WOU=XgLZ-MEVC@6(-G:I47
LUQTH-RYYdZGJ&M2CMAb)13#<[,572?1P=L_S;V=?=51[eJRA=Nd-5QB54_B:a[/
\^X2&5P7?CI)4/K,O[b\D)PU::fbd@PC<^g][][+UGIEZBUg8+D84aGaKC0f\J8V
&1B_RIR_Wa\\c09R9S(,7[(&<5cY&O(MH9^bW9LM5+@P,MQC&O&CbP7S\^QObR5;
8a])_a^-<V)>MV/TPOI>4QYP,)XbH005MZe@<g=F->F-?Z:Z\AOWS)1O4P^f5c(?
=F5,NbAd1<a22F6JNE)gPIA._E9TZ>W70E4/Eb_CeSOK)_8E?D[=e[+=1W)QLN5O
\gdW#[OR59cB3;2^]g3?eH<=TZ=V&@#EA347[ed1[Sbc>2<Pb/=04_?.<5>X>BgO
B3NR02.MPMTc&QG^;>]^3ZUCc@X.-77X-S9&88eF\dE:A8/9(Z&=\b(RPX1[ReYG
d0a^F)(/&?,7cM\X/cS0ZBJ_4Odf4TY#@^\K.H;N1>VQ9A)J[e6R/YZ1+aEH;@?-
aR(2>gH=aRE7[E7@(H63KLAdQZg#,TYd4c/=eNRZMQFcOcLB0TCD(=M>88695c[U
(Q6QR_HeQYGLDH2<@1aRY23)BOF3;&>fDH:B19W&X6^8+;RJ[QU7>YHT@-7gC7bW
44gd/8#7Rf^,OeDCZffEH0WB_MNQLc3P/7WabR<(FR;HKYVDLLY7.]A,VW&PXBfY
[^:JIfX)>CPXFW>R]/@Ve)b+DfUA_2f724(Y^HI-\@#dZQ<]C;45]]cN+,:C+D>9
)87=BN4W[C[)9_XK/V4K2)W=cXg^-c+6O6G&gEQRd/gK=7:T=H-<-LP;6&#<JFGF
=I\MD_eGB;&]5:7]]eVTPE+5+.d<VKM>-4KI[Y_/R@H.Ed?LC7>>;RG=U>214UK.
<1=N_L7<,R6&SYgVeaV3KeY8-H,\6L,FJ#)4N7\a88dOd@8G:d0QGHXc4C3VAP4U
W:UO)=GO;(@e;<:U+E<c_5bD;\BD?_+=2-.>@XeU<@S9Te:1[N>U5C(Y68TQ1gB7
+B_CN/P9I?O>bJ0BOLcW-3>,88,RZN9N,OH?LeaA6+MFR(1<5BZPAY;WFP_-KcZP
_JEE\E/c[-d,D3-K_C^&dC+0eS]aORZP5QdW,L/-:]&MHYZZ.AF+]S,N<)#H^,:[
#@2_Y_9P,JR-M,H<VfVF.P5,Z28d:>R8=HWd[](NH]-aU<HB4P^VD_d^YOVC<OBL
Vg],G8]BY-NW-CH.BST4C49eG6?T.(M]?5IX&[.5/-Q@@91.a#.fC2\(=Q.BdUg?
gY9ZCI])-feGY=+?[X27=E\TC794[a&:R\XbJ[0O3c[5=e?OF6V;F7Q23Gf[[8fG
9LVa&YS/_5YYYWOfX^:ZO5FL._6?JNT?gM]?Vea-(e.1VVa\L+N(T>^^L3PaO^I?
FG/,ZIWe9Y#55_]eeN;6[:CNLQ#McI.M&:OBHCBAcECP_^eQ6#&]T9(a]A_12SL4
OHSGJ([>D]F9F2FTg9>(_K=b8\Pf[2U8eb[)]TRaK&^P0&H30_7Te#-Wb9PV[;gE
Z8]b6D9UZK?S3A-NQ30JYM+Z+N#9Z@.a809=W/<HeeQ?HVZHX2((-_cSI7V3dL#6
>,dJ(5P(eaIWE9@PPZVCeTOE<5W-HG+Q>2V,N?1A/g4JEc_V1[VcE&g:W6MC<_gY
;>>P9:LZPC_<Md]:=;#g]&)F+,[DBI+P/J4+3g7?&01ZR7cVV.(,AR/I<76gZY<#
N\5@UfG45aS7eQ+D0)=&-@T7Z:WM9;_@U\e4YY-fOIYV+a+Q<J1Y<.(bPHX.Z@d<
=RX+(?>CZOcPb+U_@(,Q\gga<#>0f5O4bcNS):,\_#bK9+=F42G[9?I2O>^7/YS6
-+c1PK2[2<T=SP>aS:180LB?K:MR9F;7&Z6AMZe_KOYaZ;G]a?O]DM7YQXfDH2>9
ZA_00BbOf:_XX+6#H1AIV=UOYB&NY:K=?Z<MJd>1YFV[)/B;,--ddE4d=;);eGeQ
.Y#7/Za8U-a8)BgW>6D=-X;IM-cKC.\R:1\.,@1?MQYWU70M4WKI#c;:])&XQK3Q
,344JCd,Nd>>QWAR,d;6fRL&/W8/?G;(\Z5#,]B)Y7@GaX(e(SO,V6/UG@>f9c#F
XaQ#NL/<^d8WgEbFbZ0a&,O0IDVJ-L6RaQS=eX-b5T6S439V/8VDT+,&>L;8KTA?
2g2;;7PE:27#^&N>@W+&G;4FbbRY1&63,/bN[,#WQVH)AL5&.E_&,(&G6A9T46@N
:CUA6VQPZbZ2M.W;XGR&4caGXQB.K6E-N<cPE?+VW=2KK.&I=^#[LX?CeN]NX0\P
K-WSg5H#P]K\D;?2AJN\:Of9)_]\bS824]5+5U\[DEW+Z(<>TEJ]W-1NTDbP/0.O
MC)EEXK7VX<aIH?Yde/>#3-;WG#5.^[ZB+>7J:A/Q:28:>OcX8SX\>IXB?DP]=G,
^)c?g/+RJRbJY&JV)V5^2KH#PV1,>3cb?3SS,&-E0N.P<[LHK=:WSG2d_g6fP)e#
Re)=0Hf<]f(I_EA.P^N,WTYEL(,d3cZ=KZ67Wa051<,Y=A6[=RJOPPCe:0,3YPM&
I-3?QN3,_#GMOTaX>1&UOFAQUe6>PS?RH[=e_1:)FO;F1.TLKTg)E#9:TQ]aST3Z
fIAY\Q>Jbb:TPB#IZX_\8fJ>IBL4=TPB^F/40^@Wa[3[Eag5<bVXCH>e3M2AFCQQ
c>]JA-9gaR/4Yd(a?I_CC7YB\-=FV=S8IPH^P2Zf_+gfV;EO7X-,G8J]KR=I#AOL
b>O=(P;cdd7f,-=1VCMSGPWDBDHG;)ZaL&C[[a>Dg2.JX9/EP5Lf36Y5<K?&;27^
WC2,_TT+FHaTVH/LV<fN8IRWJ:HP(FT6C3JQQJ\[(c90DEfG/-:V&,7UOF-eV3]/
IQL\bDY^BFWTHELGZ+@Ag:48X8gV-7XG_6N?1-dI^&C2I0EAff-_,+eOQK8RcJL_
M>QIK\2A?M:VG;6FNN/SdJ6U1AR&M\F:#JADB6aE:O:U=V8I_?RS>e,0:g>Nd7^=
cVZ^226@O3EaV<(F/QVKOG2AE&2:AL(NbFFGUMW7;_edCY^ZM)NbTL)/@(Kb;@cD
[VJ:[&JKe-0?UeF-=P=aENa-^;-W1-<9KDd\&JAM(0J1;(B0.NYKe^2N)D\a6NL+
NJP#?3]2^7f.g(+5_(-TZaJDBeQT12:BF+[A[9dL+RGY15)L2:\\WPTCBOP,1?8+
#g53?N_8cUeDIFD-7?.#_/-9C\+0b7@de\L9^N0YAT@IC1XdBV-e8GL5[E<SE+:E
X0BdBI7MFY[VaA#R@L#?GYRgC5LD8VBbMRIJQ:)&\ILPY^9IR<G/WTUVJRfKLcgB
BNC(aNVQUP2^(Y[+YdGCY^+d:3()d0UX#(O\8GD4O+ecf6:4=<RBR?P55gK#MHM\
P-.AA^F:&B/_?DKd7K);:(]=U-_7P[VSS25YdOPL(R6;=ZFWFKWRS1d7Y/K(8IVN
PF(R<W6Q87JPAZbgQg?;<4EW#&_MM;;](dcK7WX)INeF\c0Ra=426cXDJ4))?#-:
WP:R@;=#GY5ePG+)Vd^9E[NFN9^,=OT];8M.@8c/#5(A-_CAc7E,_QMHQ3.V5dD#
@-OZO[f-W9)9.GA#(OKcI]HGJIf.S=C_K<;f^4;MB[[f;:I&5G/=[R2dL?eOc\&\
1WU??>W&GRJcf90GT^>.KMV2UH>0,WR<K4TVQe5_AQL8)M/\/XXN=1HSc7bG)5b7
2NZO/]SDg81;+@I-W)_UgU\7YR)#f_X>Q;SC3D,^J^eU>\gKPNYG-#G>Qg_0Og:6
OfOH_M#@2_5TF&Fe_1/a)HCDI]+5H<>S[UT+_C=)7J6GFLMD(2YX>A@]A\N<S6P#
Q33]b@,BO[e@+1/Ha7R?@O[=::IQc&N10&]L[6C50C1M=YaOFP,+QATYI7Q=<@GQ
5<TX<]V(1eE7]7>\5b#F.:QH>UXZ9c?B),MZAE#:?>cOCg7Mg)^W,B6SWDFX2GHB
&G:2V[9^1[<>V[#NK)B94J\:WAa+]I#14TN1;aDC^WTS<U:N?a5[&GYUTJ.d3YgE
Z]BTc:R/0F?SZ<-CK91aF_IKR78AfL:-4JNFgeG9/H=-WHT&GT1B):a5PAgC_HIC
/V9OPB=c7]Xd,a74cf<Cg.>Q4E?Kcb]M@:5eHNPPP3SUM1NJ\]<U.bAM@bZC2>JN
T,V^^II,fZ,P4+(=0XUXHS[@1V;O#JKgJAZ-&TTHDG57+,RERS+33G:?])3J;EDQ
B4KQ+[T8I[EK:<50Jd.-/T9:d:?[+d:E<a#MDW=3b+ASc(X>/^;RYEF-/&(-dd^2
32@A?CQWPGC;egWGc)Fa>8+HJK]F3S(>OAFQG_3)P-H//KJ^TN)4[N6H95F<;PEJ
P?<)TQCfI-)]:-]c+#[7XS&.T>_,]^R5W@0#cBPPXF^aXFAf\NEB<H=_@FLDdRT/
Eg_<NC(&@ZLER7g(<LO=>XI1Be\Y\CDX(C(.X3dWSe:&OXC+3d?T9#8[8IKb878\
RSKOd[4#a)b3H.F946/D7W+C#&#=)O/B0:eCY=@JI,dd]N+/1gP2INe#GN245R1g
8(SCCLLSR@G5gA;N51Qa]OCbFH3]c;FFHKQg_-HTe5])B_\WgMaXDL1=[CV3I9e.
(U&WQ/(1cN\,@II0O0HKgQF1fI@F,\RbDFW176?<YO4(B5Id.a,:+MI;1T#/I:7B
O@JAad)JdG;H0+URW7>?&b1H^:]AJD\PR\4e_MYUf0,8\3d:E@g<GZ4F<Vb5MHJ)
&/3:-0ZG+e3V+7cTSESZV:7d/QTFKV;,Y/aQV]__0FXEF+Z3<08EHKFM0J<[@Z4#
e87[WR+.N#JA/;>^Z919C3FX8PU+<,1/MVV>^?,^eOgSWQP@X]E4X0RS;6+VHJbN
:Hdg3CgQ6E7dTW,.6J>Z]dGQ4,E++^N=CI._cU,2E96K-@FK1M=R#YHUQ&Z:UL5I
e+)cV7W5PdP8+5WHE?^J9aKVE3+<ER?a>JWVZCW0Y5C4J>T1)GVK6SNJA2IE:c21
aP/<J[/((KF0+f;/1/7+P&d4D((\FU62ZYL^IQS[=PM+23DVS[S->-EZ4DNJ5FI4
^:c,I7PL8:4dcQ\S2>X0M[YYIHP;TUQO<#dQ9^JF3@8HUJYe>/^BW483UI:IZ/6f
X+T=EPPQSbFb_d,Y996NQB=VfO@eM-2=+/+TcN;/BD^8CTR/O[B>N,ELX28FJ02R
N2-9G\g0^/2>),aW,SL6;E;04XHV^^?;FJXZLMIQ;a#OGAg4NP??:B(.#\1GJ#],
/:VdL/-7]D_BTV[Yf3D1@UAT4BT-C1CBSdM]f-UcB0#KNN.138?>1SU/7MdN@a7V
1Z4<+c(/BP>3/e4XSJ&;T@:@)Q.e)>P@P2f+J/OI0^e,e#fN9?OI&e-5^\Gf5Cg#
T<A42_>bOFM;W=8gPf;O_@R-,7W)dQ5:BQ_7E6;GZ<?,Icc#>H0:8bF(HZ9T#PQd
Vd14DB^JO0A<0,C?[4],JUN7_-5VPO^(T+.^fV\=Ka9XP80C1REC/(9^MZH,O;JI
fd1JCP@I=U[A\0(WA10CaC@7KKKD4:KGV;MF1LGM7/aC:Qa:O8KOJRGO>)/c\J3Q
cA_^Z(aMGIgd?)Z[#-2a+XH9_@DCYZ9)4eUW-I&I]d9]O-M8X_MHE:>/JgaX,Z#B
J1:6fB\5I8H5>S[7Xc-(?eYR2<+EEcU3C:613;LYZLR-B4;O40)<]gfQ-KU8/aKE
=4&=G/G97_T=IY[eV(V;>V\Ea>_]DAYO1N=\d1O4Ia?.(44_=23V@7<<;&H6+9S&
dL/Y)AO#QKgfM^J=IZT4Fb.-P&2DD#R8FF5aC48>FaUHU;HX@;Nd;1C[2\bA7.@?
R:-+Me+JHb#G,M#EMGeAJ8bMIW3<S0X.4K7?+HN/:_U?LMPHKXS=HM@Ece:/PZfM
S#b-9R@@Cc(7&gI&Mb\I47WbA57g5TAZ#W7DRFeD765UQ+N0+HXPZ\>SQfgU;5ZV
^a[OWQI6VWF4>2<CSM8[e;4.5a#@^TRDQf17)2>D5YL=.Qg&H/7_(VS1^O^MYLf]
=)SOE<X<JZb2@,C53eQ=]D@OK+YH=_S#ZFI/WY-]E;MHO^\\^N\&Y<-\fL/O^#dd
\\;S;\244&_dad)Cb0_=5gaGM3fLG\22?O/7g7XAXNfVP[R2:ZW+4cU-)D@>LEe<
^4L.PBT.H>d3DZKJa)9UTBg:+=L<FZ+:/X=)L#DREBTB09K58a)<VTS.U22K)+a>
=.TY<QUa:MIGJ+2cL0;dNd==A<TWN5D_X([be#]M6>413ee.B^/6@9OM?af#_P?#
=D4E4UL+bFCfR0Ta<@#3,4Ae3Jb/2&81S#EZ]A:c5aRP:eNQ>2=NXM?MNb<a:fZQ
cDfN,=L^9)Rf,GVEK71]_\f[PMYY9a0@3#RcTAGY<g\F<,5P?W#DUfCILB?PM[A+
0e::0C=60.Y+5EF^+1QgF;@IYACP;d)e,NUL@a)<-8f]YFd^,ETT2e>dH@?:SAIM
?;D6LCF/O\?=M7b6R?E7MOb1<(WQc3E\28GNe4DTF@_b(POJ(A9UOX,VTQ0Y_fM@
6fbc#8=\;Of)Xcg-,4cQJCN8A&Qf3TZ79(^HNZ3S,aXTL.,XdD72JJg/:KG>LMD0
L10YE??6b2:MB9bb=0+1,N>VIE-SX>,#,#T#DK;:;511L<W<6>\QZe\f3C0@-\B6
EfUG8TP>.J+3Bd1dUf;O<R452UU1Y]7cZN3C&39]S3MU^S.@0[ST.5a_ERc5\>\S
_Nc:=^RI7KO-e=CP,AX,[=F6(UACcfSV,0>_NLKP<<B)FWSg/^59CV1818T89/)F
E<Kd6fE@38PWNcWQ.NFZ2?DF[.c5GA@;8WO/]<N[ESW1[d(0_HO)H/1[(5274XDP
YENIU.f;CO<LB#VHH[Ra(8g4L0:]&b((_A63^E3]T,#aaAFFD4]Q+R^:\e?C/W=&
-I\N;e3-\R,JLS^0Qe0<C5A\2Y00Y(GQeR+b9NHP3E<@UV&a0,TJ9LG-6D>/5WWJ
\-7VP?=:ZQ18=D^aa?EceY]eD@7,P:Nb&F7DUSB(^Ud4[(RBMQ#AcI#F855ORdI\
(0@9BY7]7P5;V6W#F,6X,1BXe-a5#e,RcH\BD.9ddHK&@cU6AeIHLS7AC)Xc-M;b
Y09dE/Y^I]1&FIC/5;B)^=Ib]07V26+,)28)&(^65a_9:0UB[N,(e\(/TT7.?_1/
9+W+(F]+9I@^/6I+f<QW\UHS2)N_d8FM_/[NR@eA<0g82Je:1,_Z)6]Z\Lf,:/[H
Cd&G-?5)RAe2Of4&G#PI^?=b4aH,OE1A7Ja^Id#2Sg@<4CZ+KG&<TXIC=fa#P\);
bZ&_4cX[::,XU?QQ+I70cedXQ)V=]&fc7eJ8,M3Le;DONWUDKb#3&I<gPZGP\TN-
XUNd@9^\.7Q:A54Rf9^A/UN3_@N.:@M0SC4<<?+_@CV[>8W@ND^)=&5NUG]c#&:M
#MJWbJ>eF&DggT4\\8<R72c2JU(]R6f\OZOac\E6+/_1FEMb)W3EBd40]V?<P0-5
GcMb;HU@e)fT6Sc@Og,HN>H()^daK^EEYJa/45KOS>^QRe-=#0:e,N,@V]&5&:3.
gDB;4A^-Rf-Tf@.;>XK<NH+/3N_e(eX<fNd(BXfcGc,=].I=IUZD_3<BR:R[TV/X
/\7P+GfA-fK+586,LW(&eRS7\K)cEO>4+84:;9fYLJbY>+.JCH\g<<c/96H.QX9D
E^2^_TDTJ+3.J2#<5]#DWI91V9BX3>aJIKDA(-:829<[<;TW[3b?7LJ>,5+6BG4<
P^^;[/PQd.>9I]3Ee>Yg;.GARB]<.5,+[M(.7SX,&L[MYD6=abXB.f)DWYL&Y1dD
:G+69=>P@_[?F-\/C8K(bJMfePSX7SB\K;6FGM__:XfJ6I,4=#@,?;\/eI\JeIf)
0DD1@8YMPU&O?gR9492T2GcKL?^_.TE=Aa^\_MCR>PP7,(JPbNa@&W2Aa1^^N963
4V#LBZH&IV<M]^JK5X9EG_HMUeS/A15[c5;WESL6X=[d>^Vg=g?>4BPIL;IB&d2H
W-O(=O]+CSc=Ud@FY.-T_\[\7Q@6GcEZF>@T3X]OK8O0YcG.H,10S&;X(6UC=K<8
W^<?T2,XAG.ZZVTg4NF4g9)YY6=,#MWXR:c,OH37VV.T@H/]/a_f&M<RCL^8TXO6
:^4eH4^^_KH.<S],YVJEd>5I(U)JG,5U_WJ+,6Q2^=/S/X,YS(Og9N(:=YLQ(/)E
92)OF8?@;^^eSIdWAYLRX:_\V1B?9Q=UE?61,WSN@C^:XJWfbLFOHfT.VJ,N2Y;.
EY=WOFf\S+RJG,7IE1->A4da7d\W,&.@&OY4@Z;Gd)F:BUO_Cfb(A;1>KNI;.M#K
(DY3_/50V/K.,[OP)L]B7T><9ABFSLTVYX)/:\Z9)Y=1#KZST>6gL[dY].9/aAKC
R]E?K:&VF]U),R#:K\2R>TcA7^PQTN/Y9WW084f.XE>/G[PIPeN?E3(=+(=>LE]O
08UgeQCGf3J-J>S>3X2aX^T7N1BFWM57R7],C47;[V5W,:P\M[4DX@4[/Y/MGR)]
I9ED9Ud8dGd\;[)PJ(0DU3dg(,-O#.bRVJZX(.gLScZUM,;@VFBU.NOXC6)#ETN1
+6F#c:@f,XBB+S,_JSDJS^><J=aga(=(D6=:@P+P)Ea\e0^O&=CK\&26?[c>be+<
7\D7S&9Wc?Pe(^7N/)5Zb<O7&-TDbA\f3FF=c3;<dE:#S???NYSG@0[Yb=0NbX=;
AL+P^Y;QPAQab1Pb8ON(gF:FfdRTM-XD3d[;FH5V4_-S:M4?GfYQ5\g:dORbGF/_
S29SID[9fgC13;>;/FfI6UMC@<OZF7fUX5>U/fB_:>(X7CD?bDCE/@CEZ8CGYP93
6/#Lf/bf+A:8F?e:X,I:e7QPd_PX)]ANRC)A/MR;Y7X#8=gUVOC>4E]YVH=F0DdF
WQc,O4,WSZ(E:?);edXc4Q&8-29/IOIK+QFN^+F;EQ86=FCKaO/.a[bM1HFf]g4(
1.RXR;b2fD?&9?BD?^QQ<GD,J+UC7(5>7/Fd[5PD(f\4,+N@A\IR@B5YBQC4=[dZ
cX)10293R-d_/(:J/3=P1d7^DC/]>[R5B:]7@+,CF@8N_10YgUbJce845S+cZT4:
Mc0(T\>UP/R;a\9SEaR/ZM8bdVZHS;9[)be6UMJc\D9LCcbf?5B52LMAD?a=dBWG
KMg&W(BV+IFAW^C)91/+R/T(+8PXM?_;FC7Q-de/,R<(4We<V40E?[OGK4[,],1H
Eb2@RBA+KJ5I&c=J[8+VZ<GBMHa3;0Bbb[N2,H]e>>LZ:(<UDLTTF@)-_2[O?Bc\
AC8[_9WUQWDQ6ebKW8g()2/a=2N1?^O6Y]dc2A=?VYUb^40fMK)JX=@R8H.R[Z\L
PM8)@3+]=+8]0BG9+?5IBPdICbC7B<bSgC^_eS2f1\#@\AGJ8Y2Z>VQ[U(Z)T/4[
V54P)CN<FE<XBBf023MZ]McbfA@V^O3+K#QXC&J\:S[7G;N-R+?=^@Q[N$
`endprotected


`endif

`endif   // GUARD CCI400_CHECKS_ENABLED
