
`ifndef GUARD_SVT_AHB_MASTER_COMMON_SV
`define GUARD_SVT_AHB_MASTER_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_ahb_defines.svi"

/** @cond PRIVATE */
typedef class svt_ahb_master_monitor;
typedef class svt_ahb_master;  

`define SVT_AHB_MASTER_COMMON_SETUP_REBUILD_XACT(curr_xact,resp_type) \
if ((rebuild_tracking_xact == null) && \
    (monitor_mp.ahb_monitor_cb.hresp == resp_type)) begin \
  svt_ahb_master_transaction new_xact = new(); \
  rebuild_tracking_xact = curr_xact; \
`ifdef SVT_VMM_TECHNOLOGY \
  curr_xact.copy(new_xact); \
`else \
  new_xact.copy(curr_xact); \
`endif \
  new_xact.cfg = curr_xact.cfg; \
  rebuild_tracking_xact.is_trace_enabled = 1; \
  curr_xact = new_xact; \
end

class svt_ahb_master_common#(type MONITOR_MP = virtual svt_ahb_master_if.svt_ahb_monitor_modport,
                             type DEBUG_MP = virtual svt_ahb_master_if.svt_ahb_debug_modport)
  extends svt_ahb_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  svt_ahb_master_monitor master_monitor;
  
  /** Analysis port makes observed tranactions available to the user */
  // Shifted this from base common to master common parameterized with master monitor, master transaction.
  // For UVM, it is available in the base class ahb_common.
`ifdef SVT_VMM_TECHNOLOGY
  vmm_tlm_analysis_port#(svt_ahb_master_monitor, svt_ahb_master_transaction) item_observed_port;
`endif

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Monitor VIP modport */
  protected MONITOR_MP monitor_mp;

  /** Debug VIP modport */
  protected DEBUG_MP debug_mp;

  /** Reference to the system configuration */
  protected svt_ahb_master_configuration cfg;

  /** Reference to the address phase active transaction */
  protected svt_ahb_master_transaction active_addr_phase_xact;

  /** Reference to the data phase active transaction */
  protected svt_ahb_master_transaction active_data_phase_xact;

  /** Reference to the current active split/retry/rebuild on error/ebt due to loss of grant transaction */
  protected svt_ahb_master_transaction rebuild_tracking_xact;

  /** Drive data process used for handshaking between phases  */
  protected process sample_common_proc;

  /**
   * Flag that is set during the first cycle of an error response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_error_resp;

   /**
   * Flag that is set during the first cycle of a RETRY response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_retry_resp;

  /**
   * Flag that is set during the first cycle of a SPLIT response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_split_resp;

  /**
   * Flag that is set during the first cycle of a XFAIL response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_xfail_resp;

  /**
   * Used as a flag to initiate the zero cycle OKAY response.  The value of the string
   * represents the cause for the zero cycle OKAY check to be initiated.
   */
  protected string check_zero_cycle_okay = "";
  
  /**
   * Flag indicating if a rebuild using SINGLE is pending.
   */
   bit has_rebuild_single = 0;

  /**
   * Flag indicating not to call the transaction ended callback.
   */
   bit drop_xact;
 
  /**
   * Enum which indicates the location of beat address with respect to WRAP
   * boundary.
   */
  protected svt_ahb_transaction::beat_addr_wrt_wrap_boundary_enum beat_addr_wrt_wrap_boundary = svt_ahb_transaction::ADDRESS_STATUS_INITIAL;

  /**
   * This flag is used to indicate that rebuild is required using wrap boundary
   * as the starting address.
   */
  protected bit rebuild_using_wrap_boundary_as_start_addr = 0;

  /**
   * Internal flag to know wait_state_timeout is in progress to avoid it be called for every clock 
   */
  protected bit wait_state_timeout_in_progress = 0;
  
  /** Indicates if beat_started_cb is called */
  protected bit beat_cb_flag;

  /** Indicates if the HREADY got determined HIGH during BUSY. Means that beat_ended
   *  callback corresponding to previous address beat has been called. So using this we
   *  can aviod the beat_ended callback getting called again for the same beat during 
   *  the BUSY or even during the SEQ trans type of next beat
   */
  protected bit first_busy_cycle; 

  /** This flag is used to control the delay insertion in reset phase and main
   *  method for VMM while processing the initial reset. The value will be 0 in 
   *  reset_ph to bypass a clock cycle delay and in main method it will be 1 allowing 
   *  the delay insertion.
   */
  bit reset_delay_flag =0;

  /** Event triggered when a transaction that needs to be rebuilt starts the last beat. */
  event rebuilt_last_beat;
  
  /** Event triggered when read data is successfully sampled. */
  event sampled_read_data;

  /** Event triggered when response is successfully sampled. */
  event sampled_response;

  /** This variable is used to store the beat data value once it is sampled */
  logic[`SVT_AHB_MAX_DATA_WIDTH-1:0]      sampled_beat_data;

  /** This variable is used to store beat number once it is sampled */
  int sampled_beat_num;

  /** This variable is used to store address value during write once it is
   * sampled */
   logic [(`SVT_AHB_MAX_ADDR_WIDTH - 1):0]    sampled_haddr;


  /** Event indicating that bus ownership flags are updated */
  //event updated_bus_ownership_flags;

  /** Indicates if I am the current hmaster */
  //bit   curr_hmaster_is_me = 0;
  
  /** Indicates if I am the previous hmaster */
  //bit   prev_hmaster_is_me = 0;
  //vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
BtAnE2qBF3QOlcJPbKXJB7JoW1ZOG93z9N6cwvq4qLNqGAeDiCFxyr0maqGFPkhD
9Lgp4tSBe3EoM1w8Fa/vwl0kXcwurqpjLsp1VmuUvkWU/Awn/n69VDMA9Wx87ryn
8mniS4Hpl9hjzd/COuigo1UuKtfP+vqcFz3z7VLT6mM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 470       )
1vr1dTpT8VI69FaWV5Ph9HlPk5eoMI219Zme5989i0JBA15M104uTlCSDL4z2zhx
1F0HU5FCoKq9AutrYuJ/utkofx/VvhabcdClSK2/ME5l1aMDDJPTHF//4tsoBlJy
y6/rsxMQvy7y+n9iJbOoBrqeJAvpy/uECpRvqFRsFt3Gi/40ovcADAFBIraCBc5G
IyyfjPBqVjDPeV3k8Zd12DLATU892nB7r0+uwTfhGqTsZbE/RNaT2dRUPORMkHm9
iVJWeCvi3w0FiRdtRUXrtU2NeklokXQskeJuhQG3susK2IOBkmN+Zu99MPbviPk4
KlpxJm74hv/QaPXVpFZB+/y8kyYHgOb3WgKixUlVgyzq/GG3eo9dj6+oLPNyC2pG
BoKZzG8VFZg1oRzTrgP0NVneZ54bGWZTlllsoBSVsy2wXoFqVBAJenfqBwx7Lmda
t2tniIrawi6PXI9z3YxB4eTF/fSEFzZD57DcOmqi+JS6nAYViCMCHB9NZALmWGJm
FldRGN0yuzuI7RLTk+Ka3k49rlKhhQIeBxAnTdM+4xUBuBpYJeUNXD6PZdZkKIb8
B6u0ReumXt+bVsT9RmfsRfJeGCkXcjV4MOo7Fi8/lnej0XHrqrcujVHvkoB0/UKP
`pragma protect end_protected
  // ****************************************************************************
  // TIMERS
  // ****************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_ahb_master_configuration cfg, svt_xactor xactor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   *
   * @param reporter UVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_ahb_master_configuration cfg, `SVT_XVM(report_object) reporter);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Issues beat ended callback for active and passive master */
  extern virtual task issue_beat_ended_callback(svt_ahb_master_transaction xact);  

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Update flags when reset is detected */
  extern virtual task update_on_reset();

  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();

  /** Monitor the data phase signals
   *
   * This method only monitors the data phase signals that are common between the driver
   * and the monitor (only the read data bus).  The driver (svt_ahb_master_active_common)
   * maintains the write data if the VIP is in active mode, and the monitor
   * (svt_ahb_master_passive_common) maintains the write data if in passive mode.
   */
  extern virtual task sample_common();

  /** Returns the expected address value for a particular beat based upon address,
   *  datawidth and endianess */
  extern virtual function logic[(`SVT_AHB_MAX_ADDR_WIDTH - 1):0] generate_beat_address(int beat_num, svt_ahb_transaction xact);

  /** Check if a rebuilt transaction is complete */
  extern virtual function bit check_rebuild_complete(svt_ahb_master_transaction xact, int completed_beats);

`ifndef SVT_VMM_TECHNOLOGY
  /**
   * Transmit response to transaction.
   */
  extern virtual task send_response(svt_ahb_master_transaction xact);
`endif

  /**
   * Executes the steps necessary to complete the transaction:
   *   - Triggers the TX_ENDED event
   *   - Updates the data phase status property
   *   - Calls method svt_end_tr to update the transaction events
   *   - Executes callbacks associated with a transaction ending
   *   - Places the transaction in the item_observed analysis port
   *   .
   * 
   * @param xact Transaction which is ended
   * @param xact_rebuild_in_progress Indicates if this method is called during rebuild process
   */
  extern virtual task complete_transaction(svt_ahb_master_transaction xact, bit xact_rebuild_in_progress = 0);

  /** Creates the transaction timer */
  extern virtual function svt_timer create_xact_timer();

  /** Tracks transaction end */
  extern virtual task track_transaction_timeout(svt_ahb_transaction xact);

  /** Creates the wait state timer */
  extern virtual function svt_timer create_wait_state_timer();

  /** Tracks wait state */
  extern virtual task track_wait_state_timeout();

  /**
   * Utility which can be used to determine if the common file is used in a passive
   * context.
   */
  extern virtual function bit is_passive_mode();

  /** Indicates if it is required to abort without rebuilding on retry response 
   *  @param curr_xact current transaction handle under context
   */
  extern virtual function bit is_rebuild_on_retry(svt_ahb_master_transaction curr_xact);

  /** 
   *  Returns number of retry responses received for the given transaction
   *  @param curr_xact current transaction handle under context
   */
  extern virtual function int num_retry_responses_received(svt_ahb_master_transaction curr_xact);
  
`ifdef SVT_UVM_TECHNOLOGY
  /**
   * Map a single AHB transaction to a corresponding PV-annotated TLM GP transaction
   */
  extern virtual function uvm_tlm_generic_payload map_ahb_to_tlm_gp(svt_ahb_master_transaction ahb);
`endif

//***************************************************************

endclass
/** @endcond */

// -----------------------------------------------------------------------------
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ddkrcBYq1y0/3MvLAeKF/Ti4eSxrlbxU3BHNSIwpmnqWVnoTLo7MsUKI32k9uJoi
RdVN8hU+QnejjSmSMdCiYwxUYa5WuxZasGvGgLpGM0L/8KBqUKNWtH0Ggqs98wSK
SVvGw4C+q6WKjkipBCLR4wAqpByQC+1wgecH4swFBWc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1933      )
DgGKtWS/gahj7SpNnhpogTgv7CVXNkUh8sn8V3VLzYd/fZcV6Cxk1OOKcBLfyuZg
rnV4aZTTO+T5T7PmEQqt0JXpqNpljdPdnT3h7bH1ZdEyCmsJr+F9D851g5ciNifC
zE26vLww9MZLSRNC+zFD6f9xIj4zPmeK83beFpVGvNt6QyuUJneCqyHvsWc9wkBw
6K6lEtn3NBsN6UhH0MaWebcXd9i4J7nVCtnWdtuaamRKxvH7rn6PJUGx9Wf0Volt
RL++JhMs+e1RyDpdkzOJcu5tSRE0+2v0qTRCwuGiBExzyNdwPiIXtyalvdgBo7xU
NxDj5z++eXhmunPW2EoVk+MXHgBwKaVcjnbhRV5gOlbmWBuvd6BsC/pJQdxERXu3
1fvo/lNxRvaitt+aFqkfKNrMuhigt/8nR6kDJ0f2UGLv2L4B3cQ9k1q2E5DM+srh
0V+C+BLHWPUq5YbaTVcCr/ev3fwqUxComKHyxjNKU381KPUeLjvykqChipTL1ewt
BynqcQXWuSCiVPYvvYQEkdMPynBGLmQQ3pjr7+EUxbWx+1ydZgRPIrv/6/1HNXYh
/xIbdzgocGfzXza4jQG8guaKqglgKJq4gfZpr0zJFxlkTYeIC2KUQ6oJzYfIGDvy
/E6xwkZBX4636X8EHKZqdqlJ7T3B23IECSqrQMdmJImbT7QemXNj0/Z8pk6SMyVP
AUXwo7vPDjPJ1DZ90AF5y1+H6akkmzv+E+i9LNcN9t9aTKpNyCURCW9M8x6owBFg
mvudUXKaevy61toWgfZaZU97OmxtSqbOCU11UJWg1WfdqgzLZNfKpiIPyrMRx2Ci
/rXjbN+7bd8DwC4jjsvfodZ4uH62GPCgA7JiUen2lbFxnBikv2C3T/bynIjgOYXG
Av80Jz1y+q0RSQy8w05vqzkofW1xSjjSBOv2f9OhF8UkqTeESQKESKYo+tFbLpIB
ATqsCMLIWg7mBHONgqzmpCRjGfYQlIi0rxxfxJv2VcC3zSx3x4M66GG8+wzYpOxV
ob9msR46rl6dryw2oSGuXFEq0Lh30g3LfnmrEcdSfpOCK7N7yigw/pLP5i/3u+Pr
Mot3KESSclYDfbKvAltNJrwGwtC9NpJHFoca3ZV4jitcO+5XvgXQk8rGLtdp/3Q5
KfqD38430iVYDKhKV68VJPGp1ERsKcAwsq9qR0vKD/T1JCn7Zy64047rsWIZW2tl
Ss3nnc3TveIcqR9qadPal8kvuZrClFau5VJksiWhHrXcPPeE40XmcZMd3xYf8OKL
Nyp50gejf1Q2JYAv1+VVwNWE/qTKSqzYIGeuxsWohxH61erWDFxXW2LmVewKCSvA
DXJjB+cXI8YWmGPQKb4qzhy60aFRUM52jkfLuQ0QLboJr1TWEN5cZT9e8ioJDc2N
bnHsJVicdU2OpEdKKDzbaS15JvwNaVLV5IP7Rp2B2Qqk+adlGeNTTdTRxMRyWP3n
8BRZpX9dAdD7Jf/2VT2kjyVXyJ5QeuzSuAUk3mtoClgKUlz21YbdWCx0CFsTIfmD
RwvrtTN8SU4wq5xu0AiTnb8Of3xtUj3fdfTKgFMRps7BG08pAnXarMeBTJ4KAcgu
wu3hmsKWW9DF4AvGZCzonCT+8IqvDo2AVKgy+t1lcIjM7ZtP3oFBteIgZ7dsmweZ
36PVM8kIs/f9iWM/ls/EC9wMas0K+siYIfDaq27tqlwQt68FuaLl7g8Q5lXzErFt
NgyaqHySmr22VX7knGVa0lFJvK17wklvkVZEQcW3PAKRMC/6ea/XQGjmcBIoS/6J
GZJArOrYGRsPlta1n5gNOdGHzyVFN+n/rzvT7j6Kd+jCQjb7NeMXWrR1BSKgROtH
ceyRKiGn8pC68lNh59qbb43QVeu9SXbJVk6hCf/E/ZrNdX0hTx4khbPCOM8qVS9n
4MZUb/9RpqMPEOsOasg5+0Uyz5/5ImhwkNevg3hpZBA=
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
QLuFGJpphmcw+fq26EcG6S/4ROoZH/3lIzGmBvOc3q5J35RlpyhcC+9jNvG0ATFv
r2tzbc4xiuQzIuNET/e5vUQdCm5A6v0mw4Vi3TPrqXn/7OTTDdJFvc+y6+C3ntif
1KIh63d+l/ac9YPSZtJFjOzPZZ4aM7+PMsHXUafs0Y4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 7796      )
R/cqz30Rq0eG2FnAL3hoV1igwNOnow37fxusXWrpDs3wFZNO/pyBO0Ia/AROmbW6
sz7mPrnQVaeiGRGQO8sj6Je0oaO44OZqv7xUVcvus8Swk0kAVhyXHG0a7Dnedefl
Gi87jKNK+8KN2oupDhnBSiBJj9o4HEtAu8E+XndSJxHoZFXe5lCp99UfP6TfcMIi
qTkCiwV7EgmzDm9Qdmzc50sUzUYSlyH+NCJm7QrT9uFppY9vwRR5BQTNo2YjwWhb
QA8lGjiCcAWHmbZDKbqsjQQmiNZv4rtAff8wwZkJ8IZkIlpyJCSej4mELL4Y/R9l
fQplgnS1MGX20b9xcFSwQe/ttHC0pPmm3vhRPXmVglK0DVNT2yj494GHErTYbaOr
zwNlhujrV0EIp59l1LiWVoDeiqQWGzHGCVmd3GrrcEdCm6zglpv2ejDO13Z1gEop
hapw9G6BBgL/K0FpRIob6FKnJNKoP9sDMmpXTQSQbRzt2XHV2zc2te26bDR5IFqE
EACv2LG/gfbNDscQSRL+t+4aBLlYM0l3562P2Y7uKZ3eLBeN+LnE3xVxFNmDUfyV
INgK/PaX9fclT/RGFsFRAyEh5KuUQqZoHE3WiwQz5mv03I3py2DGe7wgpXYP5MK4
QOK9ML9bZvsaB99zeZ7+Gx5Tdux8tinSBjyEuVa0CJds6SseoNEGzw0sTK8HEuNq
01N6fgABk3PvESIAk+7h+W83tiKkzidtePszFc34AeBoHjIcRqCpqiEwTPWj/N/v
5yt/Kgym/wyleHluHwXRIVcyMiWjxiKgJKkQMIaIBQi5m+/e70+fSCwSEi/NUNHo
DklW07ujBJnKQirxU2PS/r09/9yvp4I0ucQGLdzAO/38DiaBr3C2g8nEQM4ND7kb
MG4OpCY8ET4C1QwfnerXahJv56HwoGw6t/zCW6X47i9TCg5a4oviRqi9Mbka1kIE
1vbXfVgJYLs8XNne/YdNW/yLDfKVJ+szDQxWDEi+pwOqFsRNzvet7TZw7yB2fgFL
X+4wf71qCo8+Xfs7QDRfLfZnXC6Ug1A/z9Jg/lrHgY0etKBdfEvMb8kImRYeTBVr
N66d1KArr1l9Vi0jUpBMob1rqiPk6S8T7tu2PVmMmuOj3i6DI0Gl9xoFXY+mVxpM
oX4xRuDj4kVLWSdxu2NG3TaIlOr0fJv0wV/RSqf7Bh41asGb1qE3C85+sG5lFq0u
Jy0qDGvlSB8EvmFTVJrQC6BY/pkBzBqNkacZ90bccTldwAMdebnRdecntETg2I5T
t8D0Vpz1lHcTWkbr73o2LSpF4hD7GFKGYJpZjxVgzId47Hh6zuN6F6a1YtuE7+Ov
69pM8DaJSq0acN+Sld+sSc2O8ELG7j7cZAq9AbGkmO3h+OgxuaQvYuixXmZIa6Q+
ihfpsp02CrCNu7MvH9+p6CxkhDA8hfphEJRaeB7PEEyro+GSPtn2on5er6zHwC65
DYPxGFgSdvbV4wcSJfVuOhkck8MIJvPHXRqRIsmHUDR0M1zvhaLmtM/1DitCa2u9
KMst3HrGx+YHQj/P7CZ6BrQ3CIprJGXINMGgAQF4e34O7rx0tzJXNayuu8iCqgnV
wWko18gi/+CtZBzD389LfSqju6s15m3CX54LKaRjGsZo7EgHE2xx/793sURXDZ4j
ZR+E8BtGaahAq2Fyc/Yk9oolNenV0wsUPzfA+iLsQHzsEck+8OwcLBXP5eVn867T
wD9+NturY1SVsB6HxGxGEqMOiTC9vrq2vgyR8ZatL6W5t1V35+i0VIeIRwuJW7SY
bUNTuzDh4D9oPNuanCSWgaAyb2jfgDio+rHpNHUeCOva5tBJk4pwAHopqY/J3R+k
kzNNkn5krySj62vgrRLjOeq9oEcIGUWzwtfRcdwoCYAids4UsxmdQYZD55LGVcdS
U1SKcMDKUHWnOm6ZpXN+zc9eXicDJb0JzrhDEZtsWsaukcjelOLsQurUs9s1uVeX
7Sez4HL/NZtk2LY+UrywTDsN9/XJ/Sjib7Ck5TOlaK4yLoMdcb5xOwsKnibGvvvj
eNOyNnjvIN6RIz04aN/gOL5NkTPqs+V/42RsGYbVjT2N2tJzEd8ysGSwEA67krAE
Ar2UT1D2ZnIBTU/tjcnbGAvMG+61dyAgQ2r3fvXzHdPJ+snHP0wTRzmxbtpKRMJA
i7TH0AmlwHYn+gAdybH0ulaFFdoExstQyN1oPalfkqrNKwTVWbKsvFCXbQiduE1a
W3E0ALpImLtWP/7qPqUe2RwX2YZb55+R4575o0LVYvdtkgHI3XppvGwFIuHsQzoL
aHGxvkfUL4F/im8EWyzgWWYhj/bACScsZGakrWbB8OkFaClgbTBERScf7ZGoDJS7
v6Q6MBgmF3KCo91LP4vK8ljsJVjOwGIjo7GYlvnsIg7YQpjXnaVhJgkUUSVgycsC
ywdPxE0lqt1cTbEvA0ol+M8mGYmUhEryt8ZRQ0qGHRjyR2lZEDo1qRfmAOuczkSM
QERHIpPefJkXxLVFUgPm9z1v60SMOChiGIw6NHmf2nb45gvYNSpCYEhTfq+UP4qW
jLScIDNNgjA4otyE0tmPW+3zAUI8a/LPkTgh/iXKLy5d1XAGDcCMy73Cb8VLklEz
5aHyhrwIc+LsAFiZV0b29eU0scAWW7dCUIR6RDW8KJVEcvWXhg43rTt/ic0om1CM
bdEzr4nsKiC9WkQteZdaodCqcNSgkYP0vfGadP3xJxKszdaicRNHoy7TwmbwcPol
ESenA5UX3c5lI9zVwNbmYRvSKIYaL0V8TOYozQwbO/mCDQXHcNx2oAORxbCenxD4
NXdTGd4Ax3NUwZ8XxrkieVioyp7v1wAV1wdDpeZkXQWWnvUehDQ0XOXmxRXt9cP7
sheTKIHXUNicLsgYzYH5EkEHAoTQrGHRPXumNkRKCM2mcmPJAtSbdBpqoIYCZW1Y
pbmUCjiU/zIUSoY7hBedZ/bLNUpn+otKUW8lxaSNnOovqnMYFTD3BTs6v54E6uBg
vmsWwKlRBSS9UXXsqrRQWOkOYBama1YIFnbQWKF/gMyj9Vn08ljgVMEbn6CJFmCr
j8pWIgxWE4gbdcW+2aNzBi9A6NIUmtxXH2+LycgF2c9ulQ/vmCRUzr7dDZZnTIy9
Eo/IFJixk/xn979AJ2mh6imzMiH4U6c88mJGOUnZuzpYO0VsmI1ehYnLb0jHhP3c
yXs5JtE1I0BO0C0PlngDByNbyjxrot4Q0guToefUo7P8H7Wkij9w9g2PIAZqWEEv
CYU9ElmV9Q11vKiN4rGT0Vp3iNcnxlbGou8rEJdeZ37G5mzgi9mFl3gkLUfXnZcR
gkK4/uMl+3xV+5Ois2seEhDOgFuuTgcV1CRVY4IBE0VZUC//tFAmFbDT7g7yPwZu
DEmg0bvVW5wScynwP833B6+p3YBJQqYzb0WkwLaSvsISk+BinCC4TBNbIEsZSQIy
EE0TTt7GuuulgRF1rlhlgaQ2hq+5tpSrfx+T/P06E1Az3yOfnjRRB2xnjNorUwAL
2OdgVQ5qdVt5cq0Zz5hE3iEI4/Vk8ByYE1zWeyC3a6WO3dHqOmw5PYTOguLoUMLg
qdwFTZ4tAK160Y624XnTaIcgF0GfjGjLwkzPA6lSsmJKjC23Cfs982sxpgeaHWEO
6fb03Mr+nrFLD/bV9pyi0akN2GXA85UPLM25XUZw0vGdj25Wdj8/H6RHNOtQiOqO
NUCeER74Xw1Zhu1ed8IpsY1sa1YTZYTcFG5b+XFQ/Z/PRVHNwVG9dR4qZTzJ1PR5
z9hVPI7Q7wElh17xBt3Qfjpi4TKYFeNelLHEBJntZXqRFMR9+siTE5LVsXaUc/mZ
6967YsBDgh3Ri6K8tzkbr9BVOAdEg9q0ZJxPSzey5u7lrAgRJiRZgWNd2aY2pUA1
jfw19GjgoFW22zPQI1iSy0GU9nnMw4GagC9Ts9ajLZwN8c+HpV+zNRfyZEyC2xCJ
a3qKMgQveqVFeRVBOOQs1uRXZO03wQUPKEFT8mjdIWyCJofgZxhdl00q3KAv4JKT
G3J2CjGjBckM76BNlMMGe2f4HPVwyen+P2vU8NSFAsvSioGBOIncj4KzIDG89bSp
EY13Obp7oNpoIS2uykv0c2syknRPk/eLAE1EOr3LtS1+3omdM1ISAhrCwSXlHtud
8a6oUlYS/u5aX/aBv2uUextj+ad8vqL5Iop/01lhpfyQnvnVD6oEzvCV/XkLAc0t
fc377UOb/FlR2ovEHEUrzEfXmfOD1GfQEh/P8sj94/Y7kMHcn/7fBCRb+Rzffhe7
+3AMgeV66nVlMRWrI8jl9KusRzGOYNM0ADDWJD6d+X34llhf4lKT8XYE4OanZX+3
flAPyVHxU0IrQdFUOJXEXOFC7202jK62DtG5q1lLjuskwkMi5s6XKiOJ4KI0oSJm
2nNkcOCBOAxkYkuEJ5ii4SxfFBI0ymvxlqUoT0KoSErPX2TgUEMOp0pxJ05pjiYM
vvNuPE9KC0DCm9V4I2vxbW4uHjIPkNIdbUIgcWOcXFUqlJAqOmwEKMkU/Zs1gmBg
LUSbgQ5QqNul8cSDNdeDPtjLDAFxGs1C1D3kjlbd3fMtCu4192uOFTPgaQJrPSQZ
FUlWcH2V0eZ8ldHg+vur4Y1ipcruYCFzgKZBc9E3ozyRH/POpLOJ+seXSAJgZiPY
aMerhpZo2y5nm6CrNf9UOIK0fLx4cm8HNPLNZYOa6ek+Al6Jrx4C4o4VK+Q2IZQM
IJ+cyIxyQ6HhRaQhdM45ggIHc+sRH588pNFVZxMIlnn+/9J6zWVbngiYKX59BecF
EzObVklrewrmkJtU6R0K9na2aZMnV5z21tAV3VD9z6Bd9gPk9YTr1qoAk6eJIdPi
eiEhdjnca7Q63ut1aewPf55tWu2xC9u0FqX5rsl9uHkqKguDI22Epqw7mOr1YTCt
ycLRhjpnjZC8T/O4gnmn+sMt6wWmZKouSzyS3RPIxhjD2YIxeefySLsgN0Nm3jtr
fo9hW/308PhQdkOFoQ/G8x6IvHuD51N2y9WGJQr4f3vaYY7x44i/ot/y/ahJhJ3H
dIMWikm+wve91iHS2v3Y5FWzRJMPodTE/G+Sfva/ux5m0cOoMkuQLAD5Qp+5M+4x
K/T/d6CDZUvzUrGKshwqCkDBBLk60ihxvCUAtco1UUnSJKnJypnWb7VvPCJ1jZUC
YUVMrCifQdj9FvrYMCXmwfyrakErPblTJyFVIHb6VMOorYUBuVF455TnHJ4LiggF
FM9j4MdHgC97JOzgRth/N47lujGW9Sby8FBHybUHwMHupNOclllWXz3gcfFGbL0R
N9kEPS+r60u6WPhhYVVGXKfQZD3LFWy2M3CwjXoUJpGeVQGrDIxhY38FudiPR7Jy
UJ/p0mPt28kjVpWppKv5iFJqBChlP9zbUmD7UuKmj7mO0O5hASk0Ri9NQUX+lgLN
V8BmEk/MrBApIserThVOTyuLhomvy0KNSnXAbxshNB1P0alYwhQydsx12rVz0red
a4rXuNoF131CzX5DaSkKeASJrG5fzld5TbG9/shJIguOBZofhAMoF7Uj6XBLJeoJ
MN6JFonKd0iWx3QmkcTd8O7UOIkpKUa56iv6jWDVJiYLXFGoN9SI/sbf4ULLh2V4
LlLRw9sswEQBlNeDoCanJ4DI+j4ichtFjf9MyO2i4f3m4qyf9MovC+mrHgDomMem
+eXz3JBO0pq/ODn/lgcDeaxjw0QqhHtz87Vl1tfE1w/pJgRenJxrll2bKfphvtgi
FjL3gZUzsdznhCWqdCZhXDE3U18aj1bc5ttK8/7m6y96y+4zMFC1kk55juc+fRH0
sHqdXOuC3gHi8xIPAFQikQ/P7KJG1M6iiAF8kbbl/CePCzstBx+Ch2f4WqJVsf1G
H1if63amJsDedYVgmkMyyqc7+KXrMOxgEiIw4ncu86MTUs9cXnJO66nnh0sRVRZG
bGGDK8/Qt1GqJeMELCNLqbezCfhTd7F0k2mPq8HX8Y9rDgcAxk7puv2S2P9Hw3UV
4Cj2dQafZkLzdZjUggL6CxbRVtzOV/6oNq2JnVdAtGSs5ZsRTAQEQ6w00QpKbnoL
A9R/CDCmXsi7WODQdfHA7sifEsxzz7UbHyK4SLDzLnqxoigG97x3tu9PUlEQFrEu
qEjEgIDSwrqh3R6jSdD3MWdUPfl1g2S81rdIALe2CLNQwVZr1S3meUBt9uhoW9AD
eiX+OfbQHYYg9pBD+5dEQG1qHwdWTzwPzdwORX1yMxBfbcnT9hP6qhlH8zX0FC5X
yqedu06W0TidfOIiY2nL1+s6RzUZgX8skvYqsYZvlHWn0xUzPLQY4oW6NQTXX5E+
f03t/46mrlc11ShWZ1cUTD+9vyARfj801q7qhtMACd9Im3YhiXpsegQvvIJRwHgY
/ThoNhsIRIoCkAplYrjiMXNF+XFyNogbrLBTO4KZ1k76dka4xhHrbQxWgkoLTYkG
Eb4yXGKTvUrU7ZMklXhOLwgrny5Zub/7QzjG+MeAqxAKpV4lEIYItl9Fzj8+OzD+
H9SDfXEcBsJgSi/2KVVRpLcAFHKgxOQ4BSJyRv6ZEGcvzjiq743o6Mfw/phx+0Hf
P+gCQEulvOHXK+zArBquE1lupqb+EnGBexzLsw8erGgJaETGIsv6m+MzgL2puvmE
w9zeVLovJK8G0Mq6ZhOSLyrwnJKLEo6prTSIzx8mw9E4AGA6XUVFLFhhT4WW1ccF
c2JUxtAiUeMp9Y08VFm2uUzdZuN4tbpYtnkqPIINiT0Phz62qaXxpOaENp4iYJT/
cU7FDEmDWkdiFC9tmNkG4zKkhghLI9sTn01Th08XkE2nzpIcEgwiDNfRz0IjRm5k
irCoz0W8uowqAOsNmFbwxlbV/8qwiHynU9wlDURhglmU7R/GEVaTxUePpPh7BUYT
dS3qEZJZ6um+F1vYKTJOL1GJKYaQUFd+UxsJKrHcc5PtI3OsYE33dqyeItsFO+lS
NYpwpWk/Gf3hE37/p+Ul7ha61vHMQ9m2sftUxIokMHTJsqfUzJ8+Bs7cCrsBTkRu
e5AWbxHDV1rUv60x1mXr2hqupChaYRlS93XkSWrbNVQLob/QG/6Okt/XbHW5vxQT
Km13ZxNlaB52AmYrG8M4Bx4gsliHSpCTeOYA42QGK08bBxHVX6pAVPXhdEcxbAhK
nTL7AWK9GevQ6AfB5tyqCcONf15a5v0/N7DRVvMfmroxZndKkqE6aWCNQjQK6BkO
RvY55GcsQvesUBuTtCTKswr+Rfoi/MUYM7/rqeAOn5Pfn308mH0t6w0dsS5qyvPw
UlmRjA20HeguV/9ImPQ7AW06jQraeoQ4ReJTmwgPbnsXHfWJexBJJ9fxazODOK5y
IeOEPJ1U9+kXxgkPk9pPL4Tm5yMXOf1jrJYDl4NeABoG415KVaC7aKp+/EpKD1eZ
is+bJuICHR/pGdHGJrVvs3w0COe5XP90t5+ZDhJL3dK2OyfBRB1H1I7DaRzzMXMr
a2m4hWfxuYMzmVIDacTb44sHOoh0fZzAz3StR83RrucM8OHyVoEzCudYCER5rWpw
hcP0Cg9gJSUaF/J+qA7WjArUKdZzqarLt+v39oZKZLMBEiTGTOulaaCBpuyzmVin
nah1+ts1a75ldRYNLT2yYH1AXbKkKOhjY99YgTzbqErWpxGi6k1nyhs5scWdZJDh
axzTs1XGHdnJuj9Von9BxZQ8bS+9dP9Fe9KANTOIc9Ox1iusF1J5Jz9OQn9p2eZ8
9EHpjUaP4tJxcoX9Uu6fZ2V7mGWYNXEbTSzqIVXGVhCH9x7qxLVuX4DR1pey47e1
AF1G0Hdf/TUwabpUIog6yg==
`pragma protect end_protected    
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OX1XXSx54H2GrdYHlGozQtyF0VPN5rs5k1rmhT/fvVXsgPpUeRqucfaH9K5fW2Rp
/WbaFmfCznLUpkL9SCxmKoL3vgC7YM5ZF/abZBleWgRqWAgonSeM+CkDJqonb37u
Mk+rXkrXr0vhqbffng9RUPKlfnPUv2NCBK0pOdORWnU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 8532      )
7E49nM3WPku4TRad1Mrac3x40/q95+apYZYf5hhlnOZZNK4CvNmLFqGrfbX6Z47n
AMopPVNC6yzTYaICEH5dohedmRmSdDthGIq8PHZvzxHS0XBa4vfFk6A0XvUtz28x
MBJM4ECT78AYSlVIAjhINXpPjFOxKGgAYRGKOO7dDj9tiuBQb5QG9/xnokJiRUh7
j1Y50AW/cH0DW0tm5fzjCBEQURNL1f8J/BQ8tFgDewB/rfzPv1IBxVxB2ET6PrMp
IrEE18i+x2BzOZ83vREI1fpnkeYHH577zmD57DLWgiMzAIA5tqgX3bd1HblmL1jQ
JhoFGUUJQSclYQoci1U8cgMpOSn0AThJGuwca0Chbn3lyFb3UvQhtzOTwyC/YPuB
GfD7GlreCjLtjnZExE9H5FQCtm8mYsOXHf++BUB+FjKkypjSCgCef9J+uepQ8RXC
lpmgYXPxi5SkgXyaVONn8dQJqC+P+JCrO8KeXlKz7cyshAuiufIoh1kQJgrOC2sJ
+T1IE10z+CYvlHd73n9dR2F0wFdKnhh9L8uuU86Gm9Ki8b14UrpbREGDMquYahkn
TI/eDs0WGtIMSVRl93AB/RnHcJT04pK3Tx7J96fGIqbtJzVkvqQzGhE3X93cM7o7
cdyzeu3fvH7pjlfgT21LtNAWZWrfwnhemlmQpqdeV1mskUF2/lc0fGor6klLLb0K
7xxUgRkCYtn6opKymiSRZqWwVX2fCebk+kVfmatml95H2wtA5R3x5dbPE7VCelRz
LVVwosgfGE9B/C45h8cdJZOM/0rTOw/yAq7Olnserbmyjb18l9wMsD8Ql8udNQKC
ViXgu2CjWlg76N58zfUyAAguDLjD6E/EZflPwfViARonAjaqlJsvK1x+j9Dohttm
WrLHb2/6IGTtFP/2iHkjoLeKqKONp0gTeePVGOT9m8+DOAjedFJ30mifOZ1zpk/E
Nn+a/CVpx/HvbNX0/9hK3Xb2StGpdLUn1/0ms5CBHfQ=
`pragma protect end_protected    
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
mKn8m737hb23oCGdOJoM/i3rB+FIJUongkf9AHzB3nM+nT0l5Cfmd0fsaV7OccXU
hcJpQtYH6vZDL9TtCSgtUuZNz5ZOqny671M2e3zvXJ46r1VAIoXNqnp1AenRT+r+
zoLCbIvJjspINx6ukdZd0rY94EeyPHOwIaTU40DjNWc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 48327     )
dsO0HaxkecdKcQ717II48FfaSYHP6gULo9/5E6ynDOi/2ZPiqmgmyDghLt8VJ82O
gWwxE4lXWZ7NNpU2hqfoWgfyEGJ+72YLTKfbaBwZowRGJ73viH9KCwI4H+3b59tQ
IhJzxq57AzGP1p2CG3+XzDB9LDfYLrgpsrDFlRCzmYdc3h+cZY7Hoyogxtt6R9bn
nn3L9n3tK9FZYMR5FimrwU5fho9oBh5xBUcNnlgd45MN1FcNDwJ9ak9ju03nM98G
kELEo2aL/XLB3doD7mWfgERcFZitrlrkXyyCKmo+erdznSwevmh5+Cd+qO1JfLCd
IqwbF2xY7g/RJvruorUXP9fn5A533hREab8CEPheKQK9dXOXmqbFPE/PcpbG4Q2i
WtUYDI9r5Zhk3wEf6v+fZ01eNKGkMSF5ck1ZiZyN5H2QarXmF275htQJPNdK9ziF
dqEdzedZyIYUGMcIgDL35R2JC97PpCK7f61NwXPFahFZU6nRJFd80GmLbJWz7kdm
AtTr3HeFk3KgEta9tqf83Uc+5xY0In0Y4GMQlvp8dNtV6p+eYEbTIcOMh+fNfd5k
Y0Xj3kq9ATc/2UaYAvhQYPu+M75pj7pUJUFqKN7/No137FpU2fI/W3LO3At2FIpE
xfNaPJ1h1Z6Imz4QLookrCSb1UBCEQ+bV4+KkG0bYT6UcXs+PHogFQS3ok1Baaq3
QZlHogr/c6xqhoGJbSVHeIigfZ3ETwy4NAPH5/ef2oZy1GxuhtVFCd4XEPBTqA5H
7+XGnvhuP6fOrbnwnVEl+bFjaafKHx0gDXP1scPpo7fSoQNYxgM1ivAVf1KP1Hqa
ipGh5FDN1EgjNMcHrHckA4gdDN9Zv6qwvMKjGNHNqe8B2OgSms0u9FUSWYb4nclP
c/SPDKAXkWTwPrJSnlUs0XN4b4K84uXHBe/sL8YB0MgUKWaZyTjFIVTeSjH4ky5a
K5xkw219B2FOhGjB0mvoDwPAVCwBX03u8Zvoj1KSNUGmtP4WkM5dmuIMg9JA3iGg
rK4kXqj+yP58Ywui7xq4rF7hm67ymQtSl/dzAGl3RxDKcZ/QdRq1gdcOC+JFJGt4
0wq79Al+nPVvbyGc+4pF7nLql8dpzqqBrhrYMOiqW+KED3iRJctiETgnMNzP/ffa
qZvbzueC4biKiq7kcw0qYwHBnxDKwVT3+Y09JP9CUjpgRZvFPxaU83sID2Oa+9pN
jOSoz1fHGR+jzdBdAvY2Pc3a4v9Sl5UU8G1q6LNw03Cj3oC7ZH+cpOeOOs0BurQ0
2hqCF7/H+vTOeWNmYUCoYoDOO8+ES8KmdhVzGi2Eu+YW2z/1GMyDGXHbq3QGH4dU
OWFPxmzE5bxiDBH+u855vXoOg7AUtNIhUTfeWeaxnyUNVd8BK6tnshio7g8CqV5s
VniKh3FRJ+wMdLXlm3/71hug+AfdILwUCnV798Wf/EDPPBb7Lo2q/WrhomHnDE26
YoYf0nJcCZkijM+wMbgKuFZn6XeObKLf2NeYn9Fz5vC4z//o9haq2Ea5/t9XFMK0
ab+F0s5uEL/7cSABcGsfQoMsU9Uy7dbgHsYef1HnDN1jbNme1bbFeN2yFa4h8Lac
WHwJqNOkQKVwMO6TybtQJlTvFiLSxUDvPDyai3i2aJR+9WjpTPFjhrXvMn+nMP7m
C916Yi66hww5AdL4GbJuzr69kzGM1U0Xwfg0mU9w0Q8GT/2iqc4Rw5MRHdOwczuG
SUfBGD5BlcQohFVkbXp1tNfTFenkxtymPKOXNDB43eNFv4QYV2+4TRFYwFcQGGs0
IVaI60pgtKJAxjKuq5ZIk/nIC0w7u0ekFTlSvaDABkNI6+zCIwv1OuthAjE+8keC
Nnm1x7EAXQKHPfzGXPO2Mw8ws+mhiBQZm1Mfr5GJzuTC3fNjhGP+Mv97FS0b5K8b
dtZ+1GcUoltYbJVNStsBQRfzPNVeS8GL+JTVyFlBBCiJ7/bPnINstv55OuwmGyUw
BIBQlNQ5veSCvbN+KuA33a2Ki/CjmefSAAbhS4MTRZb0YiNmvDrufV3YgdeEBeqE
XIsE2Kq1rm0R68peVB9mOv0YmbUfSSDMrdyWHBcY1nwZYmCsmwu+zgIT1By5hfwk
dWyyG3dMAOrRxz909WFjc+7YeV/p4WoPlQYuhAhLR4lPf6hr0XhM+LBms5Zgc5zh
UaPCildcd83HXh3+53GhwBbdVLW2JWQe9Ur7sni8wGs9VWLH+O+n+5zNYIqUx72D
VcMLfERE034NDDEmIssRUIAYQy3r3Q2pXTc2sEC54HGbfAYfXL58BxH5cSLta8Qs
apxiDNKUALqq0PX7xy+xXcPgY9vCbH3rfVcr1TMTZkU5KXN+E10Xlfu61yUbaPOL
lBEREyFykcBeYohJO17ATs+pIcHVeEbwUeJ5vS6xOYubPt6bwyy1LERGHDmFi102
k3trKSE1gaqFGnzrPkfBgqhVXGCsSHCPP3FHhCbb2Gsa21KsQVA1/jdQnAMT3iQH
OKxCZLm3igDP33FkhQR/PjHot/hVO7K93Enf7q2845/qeX7cZmCS5Tarv6J7eVfX
WX1DNy2k+X90pVQjrZqBIB8CLvy5alA/rr0y8bdSZDQXV3ALwXhuZadhgpSV8d1Q
FzndZmPc9dWU+aVTyRsXoekuyEZrKCV7SBm39CmWb25JVr8KC9joJygBKh1RYwYR
8leN6RN8dw/Nmb6CwHsza4t79I60TnaHIqDpL3jNqzDTGKPWzNeOgGAryFTuX5qP
hdaBlHTLHrnl26BR0yS20VGyAexBtN9m4dFkvM211NrEKYHVsXbn667tYH4uUiSy
WroI6ont8GZBn0Q2vuDhJgn+asUg1GQdsLoaR/PeVJ04RXvlPRg+Ns00O/5aAjrN
/EMy1q4qrWUVc0MSdm4ac5ikfXVV0EcjFJFWQoEtUFJASvbLGHpZ1YaFQzpw8leM
AdUtAlVJ/03TlZpUxhlsdb62fYTV/VgNE/m7iD9CvzLZNgM1WIG7O+mu8eH9t0cx
HR97RH2ubK6VfDRFtOPbgSNagH1zO3MeiAy4s+0Mwo2WWMBRtRuKgFqAt1TJ3us/
jkr1S3sbjuas6sKWFY5/57VhYH+AVfVqvWVIYwzWBQGumaDBZLnjEp9FwjljBiDe
Zh3pXAsLhU85Ie7DzKSc2QCdHBfBpJFBeV3b+7nLJe9CN3qBCM3xPxZja/ENgGE4
24T2vQE2UALt+YerVYYCdEwB8OzmsjKz2v6a+EkZum+1HppLhAjo3A7Ro45nFCeu
mbQVvgEQqcUgAqY2wj9c/KPm/x1ReHNr9mk0d6gswgQzvS8W3/+LuJ/NLAi98+/k
KE86IGVn927VdSH6Er25svyruVAgK3cF6oDkokqdbXO1hrmDU5C1idgEfRM83fms
rOeswcL6OSViC2PfLU0D+B2MsCtfBFernViJ5MpMjFYPfy6sJ6XZ+8jsPakz4x+I
ZlTJC4hS6FFmJ6wdaTSEnqIl6OuIVgh7vtIl28/71zLcm/x3cmIRm3wjfDZ+Ka2I
O4wEThCGITaW2rgiDAVRvTHymcK7dmQ99HFo1smHKf0vGLtRCZ9EyOimEkL3p+6/
U1X20ccbH3xJF2VY9Pg90ITamXjc5IhQvnb2FspV/RkgAOHvcRe31KauRsddIUyL
yhQKpYqHqnxW3HWaOpi+YO8jk5Z1ezuUSSCaO8ZMC8iIxcq9RKC4E2BX1RQFApdp
i1x6fWsviLyCCxsnlL64Peqa2kxwgIAdYfuNQeHVeXsX4b7j+YOTFLPHD6VcEubV
gf1glDD4TuUthWcRLbtDJM1nFkKK4lH34fipWTUOEqfJUZzxF7YLndceF26b14cw
31bHTLj8DKK5LmYqHUS/2lV7XyAv3f81+mHfOu2t2JcFqTQpMPGjKRdVFRQJPj7L
9B34EbD4RbVlGuuwU3Kg384YSKo/Clb5rb+aO9rhWZn2gyU+YZ4Y+Jp/eORDYYvz
RnGyJk90AJxEHVj73cannzx7waHEgGszuwrRYjFrDakZvHsNRA3kOh6ZZt43ARNG
8KcJuH6edngaVclDGmbbnFZbZtOPJGg69cFyDnn7lQB7kZ7PZ4ylOhLp8T0u0wO1
QjIPH6vwvTPkkSoVAxC4aoTVKxcFNt0JI8y1zUsnNAGcoRFH5lWgQzuYyc3cnL6d
WYmQ8oiqbIjo1gs3S7d6nFlbcNTcHt28SEl1nOnAPhed+lB2RH/Z6jDI2qmWXgYx
lOGaPnfAKQW14KLpgBhC9M6jODDJ0+PPSMs1nEDyQYXbWUxhoiAifydQx2j9NNfq
Xg2T5/YjsWefnvJIrKSbcNdJN16vg2qNDFQf0cxRwSw/lhqW2JYaBnr/gZ99LDPp
+sWjUF7YIZP1k/sle4YWtwEvGslTbG0z6hV74yoUVNN6oskek8S9hcbsf2XX00py
4nQUEpZmG0kbHeeEXWnAZiTY6IIUtTSm8Gx9cUjeA+TPbFvqsNhdqKT3dnJ8bF27
4qG1NiL+rWJW0TF3CVmUa5t60QvIRcuTkVdI8tXnS2xLNg7dtJ/Gb3QPDp85g2P6
UZaOP53x98RhmtYmrZiH6SW7RwnC7yUNbizz4RJ9sKNZ4BGSH3hbd/EsVqIgAKXp
HNpn9Iq8LGiiFFz6EYWJ34AEUrKmO5I/m61IiYWlSZMOucjxm+bDpcJeJc19Z4nZ
SPcPqYFgKNoz/mCV6hDRsME3SE3IxBdNpK3v0dLz8MpV13HMLycofUBhgkpF6edh
2PkSIepM5bKyEeqnnGxXqlc2pgsQhvI3mw5Yve0CWJbVu8IK+kDQIHOzMnUZpHwF
gDOYaB9oKyc6DRMHGGFN5Mitu+cHlhe5kdcOInwuYpXdvW96oZ59HLPCBN3bqsxl
8w2bUyqybkPQobB8WV3aOrkZ7y96ewiC0qvExFKEINVwfZCHjY7AbMYneTuAiGQV
ROqh4Tozwjel+xpK+4xzej9yfkj5r3fqATzvyguPkph2FktR4HxQnvFyAUNQy6NT
OE73Z0CiLLoH9Se1MYYTvqXvEi0RgOm4Fh7sH558cOq/Cz8CgitqkHzSe2EefpkH
tuICgYdt5/aSNAmVpN6vEJTCMwIZ14df4KQW6AVux5H7hI+/XH0dqIeS0bhakUdu
SEoKwul66IKYd6Kxcj1aA0knp8KdTKdX+tj9rOmqNTl4HYKoyRVQ6V29e8MxaaQI
ytckhZvUa4c/7nkXWkzdCe/l1CI+hqYxt+FnznDEhJuFO6Yr0WooIBINLnKvkbI9
7nsfIDXF6UPoNP5zTeV0kFoazj2UYDBC+jV/0cNIUCAuT4zoy381JWip9haxT5JS
eBPWYLPCq9keEH4VYw3M+HrcNQZCIkRMBzvSDiejXcWw3Gdeeu4LZJPj9kVWSICa
ZHVc3/xjXI/phxUEj0+m0ilbTjMxg7cHyJB6dLEO1NtNTGIMIFZ0BU42AJhgG5u1
TrkGpLpiro+RYn1xgBbKkiTduFmPuEfRJtkq+sEWcFiLtbXI2KiB4DfrP94XRcFJ
f8o7BZ3XTbQLRhkNeSo8nXASjZE699LxAMPpPZ/RQMd7UCmt7+YsI9GrL0QY2cQV
TCM1iIUdMAtZNZjUC2nn7nfzM0YgyV1MLpmx2uXVRNTs6UCDQZ9JfPneI4G86xF+
ZHyaxYv+sfkqJjz0Gae0xgbDgVXP5WNtYIvYEbpE8EhACiREf8Ta440MIIOjCcvC
L/9k66gbloB9/ipyg2ZfG1g4Ub9kIvBwdgr7jFUAz3J7n746Ut7inzwo8P/ja2hv
w69bozOKyFjsLRd3bhOdlRrWR5AUeXvH8GFZHbDaByifA9cth7iKPRugGkKDc3I6
wpVtMtfWLcsDMJR9p/hXrTDaSLbU+Uh7l07ZOyH/FvOBzkv//KNgUZdcPj6KD1Qk
IfotzG1A5eDMdsxbN4+tsDQqv7cqgXueYKFwFXciojD0EdnXkH8Gr16/yRXHzakh
/nTQ7Wve29EEeW5s+R22EKwv29vUkG2RY5LtoMKjirG45gA2Kvtt/LUG0knIoz20
KC/eL1YvV+YbdKwVC6bQjK8ejCGEhJGKGwFc9ZyQQbCdjNFcdfxK0MG45wfcb1/p
9GnN0qzXv9nGJ7QddY+LEwiRUGQY9Z1/KdyDEl6wsMxAPwIFXMJydV87K9hz+LAy
1+f5NmOu9r+UKJNyrSMwryB3drcVZu71gEvVlVAQCbhTee79pCp3Pe3UK341goBv
+Lb1GMQzuhq87hlAQX2g4BZ8Q5mGo7uK4XyKpYhYxMadzWlrWM3VOs5RSPHLDgkm
DP/UkMWe9OlrW6OYBb83hmAqkyxmvLW4qNvlOIlZ8Ct6cnDwAgwi6MDYlqxgEKtI
0Skw3vDb6gxy7EGMKnX4exBAfcOibiTsmWYS3RWoDhDRbFNsAJ2KlseKWJnXLbzt
pLz/ny2xOubeGbwIc5hlNgV1ZiFGMLCVeEvULw6kRxWqRMsP78oMZFdv3Y4Fzpnz
eKeongtQnO1hJRwBsDSWGvtFJPAPr9rMzVOjLsRxfub2D8flv4KnPr2MfmHFeF2N
z6VxwbPfTGM+L+ZSygH1oVCaPVvLc2vrgFOt6mhItcn0sGwlfZQAhfe9A3XmxWvT
MaXl0VPGQe35dRsJpDeLjuqsl2NzM+e3eysX1MsI1qt86PzgfCKEvsWi5qXpN3FR
up0G2dJKPEL2zZ9O4/s0ykvTpf6uXCAQ4dAEMtAdOPrDOvKh2vIc6dbsoArxwnG0
7yQAMKiPs6vRzD4sfBN2jM/3wQC0lry8UE6tbKPq+DN4UIyrtF1cownZ1tuF5zpw
UT7iIe3UMI4w0WD1XpNMhkiUHnTUtLwfxHE/JWPxejeKa+LejoiK5OsDgijPKxqh
mbWx9JcE3hmDMtRo2Pd5dGYxxELqQRgNeO3s2cqyLnVytOwbn1CmuP74L82F3SpW
ZA7SMb150wyu2CEna54yvDHowDia6n+cTQRsWZD1ICDGvSVMf3s7T9sOcR7wpA+a
4xjf/6lXmVS8x8zir6Ih3BxhScIX013jR7Mn7CRe8xlLHlPf/J9hMKCpcSD9y0Ky
NYy6yDbvW1RxmW7rlEnTyJ4qCsVlEEZHOinFQVR59WgSE1r1P/nVnqQx5Ghobx0j
zWmR4Bmx8P7sgSn0TSSorYA5ywoRpTsOa5GMOpru2q4ORnDVe2EeYaWSrzKY+8DD
byQ8qEh97iuvAQiI8f8LV9WuyncdxW+AoFv1TJ3v53uV5dpFBNOpW+LzwFOllqC0
onSTxS31HS0AntQtn+LM+Pafp0gsOIsTgXWwJ2kdxQaJ7MK+5Zjtwkc+qr8jXNa4
KXUsCIPuMUwbfsMlCHeHtLqbkIcYmdxvTVUYNdqeUshA+2Ztn3zQFB8VwnRpQ56T
LW7VwANVZIxjXncvhN0nsm3dVrx+sHUvr5VdJcq5KloYfKSAJM1Vbt7JdPU8uUfl
NmWgwQAPEoM57gVCYyQykzRANqSad7IFxAMivtBLldIEOfWOfFr6DeY5KhgztEbI
/ngPBfzbrwMdyi/pLz5DBTtW2mBYV9umPd11pfuC+TmQOJqMczPsua76gTQKZiII
shRZ29DOwyiyvNyOGD147PTunFpEmFNpO5Et1yV1Mml0uy44jwpUzM+XNYMUL9c4
/PS3UVpocYjc3LfrfA4dtGKA9U6q68oNd+t3dXu8i0L2h/AxC4HfGtQ736ehhASG
LuU+XXteo4GTShrmdZdrHzhBLmzG1lJ4NAMJC83ain343SXh+PxZw8tmA7I+/yb1
UtC8FHktXS2odiLmke5pBZeM29FoOJ9r3u3euKUfZCdEUNZtK2VfIyhKyU5AykBE
gOqCusWBVM3yOrOjLXxKnpy7ExyRofcTCxBKMPxVWZjhAtyCl8X88Jk59M3pspIm
pwVEAd0BnV2bGsxOqMvuRJ/Qa2At87TehiO28xWHE3FC3bFtFRapiG0Tb4nuier+
YinKDcpDoDhh514aE7MxLE/6g7oS2Udz7QQDtUP4epF53Ieeo+beOlCYuPmeqqwb
+paxG0R+rCsiS+utS3LRw+2XZzroGeIs+M5Za558H2XVUwHWiVvtI3orDi+9T8EL
An8OIT77lt3z+hxnOS6mYy+ewc88zybrDNo+54zHsOLNnIgybtmETODHNbL1H+8f
B9MFrQJHHjtRwuXiCm8ceLJ2ASSDJaRi2RGl2Fk77RegrWNp80cblooXiHVY3v7C
j69EW9B+FDZL9rBaIVAC9Pue2kAN2707iDH9F2t9hnZp0I0O2+FX5m6Jr0AzGSQt
rmsOZQIJli7JvCEYLfYWOUAOc3n0kMhMyqu4X9mHX4iRrr+P8rrWaSajv+4pebiV
6dq/VWzbDXAO8PCSXbJduydICIV84qXhJF7VBzFSNX783GaPa3aENmWdV3Cxd5is
vhSyTaJjWk+NQ0GDaI/eCir81nKKbEs/Vf22kyjpIIG1csd8gk1nvPeJaiaYAML+
FL3Huz/HpaLe4+ETCeVc2ddBy5qEPRnLLmW9yZ3WqwqLJEVAu43frM5YHZKPaBLH
wQ7/w/8L7HZ6vktuli4vZIZEaTtIYY7fEA7jY/X+SHdtivq6hvSJZioP15N8PX0a
F2LAJKPsK6C48jVSjKJZosTw/2WDxBJhvC5Rc7MvxcUXU49CDNnlVLSWQ25mrkeY
qDHaieykdbBPXjwn6HLBBRSDjqxYyaQasAsp30pnksUCLz0Zvbmx91cgZJYPnChT
Bq49cz7L+w30wsyRet1UdlbsFTKlYZdT2FHWm2cXKbVJLweTAMQ/f+qd50PEIAY4
/oxPIvY82TbHQHd+RVjXCyhfsN8neo67ckdaRPY047YtDi9yNeYGyzhvatAB/YRJ
d2GcaLG7b1OQNLXPqhIK+LTNwCILzxsrvimgQNSQQhuAJxda1WY9H2i3tovl3H8h
G/lwQV+Tn5cYteOjVMkPaQcMlXjZfeSn+OJyV8d0140eIYivdLpPVnVRM1FRgUus
rgnLtpVUObW2Bwi6ZuWez2DQObgSRg/sxMYBmeHfb/9C/F82G6saTmyJDJAhu37q
CSkBUIcK1QVc3ot3CA/OKqH464bJCbLqDth3t9vDnL8zoVA8sdjxapMg/A00Lrz7
c4KH+ZdvohkgI4qKKx4B7Y/qcDCsNSKZ3zTxLTN1otTxZTPYd8PkoRZoRQqQ6oSb
v9osavj44Q5x3gCFjfv2YQr3aKFFPewHo5YEZExBS5U08i/tSJxYl9BJFTuJm0jo
bHc3TmjWDeV23Fko/IdiVAVPBV4V48+gtaHiCer6sMbEZf7dZvHBMfuURFi18N6+
ujjheWC5L2x6oD3lVW01qUuTfSPUB7tzOtcmNEso3A6zddSCJ3yxrYIASdO+iFtt
MdvmzkvxRzocElc9sKOnbQUrFggXl4vyT4PDD5JBSuKqlzMa72qcSYT6dGt04Dc2
67QPi+evIDR2AlsmE+txSveNHokZreNRwQmtgCnSxmu5mOJHxh3KbMKJgXcTe8fv
jyWxKP0F7qSZxlcv8tcCPYdy6/9zB2jR1u0MBUaWFhFlN34oLFRwsK0OnF6skHnF
Hzti9IH+UW65PmGt1+ytfgsRxl+/VRJGJmIdpdN9xD+g58Ni6B/0otQ+4Mht10KI
xbFYJcyR371fJYIYNfLBAzeYa3ZxjqWRSlKihuXDJV7mWCCbeJTrFnLoCBZ0ynuv
B1+2pT+9n1OTYuEoZfne/CN+MnqQdGYT5iGrVM12BmESDfr1sgE5Ts+dt+q6EXWg
eY5n3okU8EriFVwiSTekXsKb9eC4va1QOSrojmvVqqnDfFCqtfMSnP1WETZwa1P2
FmvB/6CjsX5NQiRJpKYqdAzJ5YD6LOY8N3ihBdYPmdjYunAjMW8Fph5JbOeKV6Fi
yiZKHnpwXpMD6pJLjX5rmfGdwonTKSaFe4a/t6nuCYnSUEnvILxHTWlNacR9QcF9
0eimFOgP8Ri6Q2bIQJwX+LLkWdwu5UhE6pesgy4x0RkmXByC9RYHEsn1ZpRdQxAg
2ptPfOspZnDfR+OaJ/rVwv/YtrfW6W+/ZUmitcoMdWv1gS3OIdnBD/GQty+2Y4lc
QUvW4cQVce8p8bbo3vbo+EEqP83JTlNBBs4CyFqepbyBlZG+XKwXZoci52jTFy0s
jeEkN2iWzgDKcvCQEnOfTmEQHOeuSFbtBNbX6xeMCqxbqK8QwFu3ktKI8MUY+Wlc
wPbdw//3vTHNdSLkUron2oynszbo3lpL4hc23PkQFbRDox8GdnwD3B6qGeLVlj55
xohB7vo3JBhEbDFMAe7rSX1wWQVuMZB0AL2kCzBG6av5pmxg10kANnilGSiJJ+rC
GX7cr90DNF8RVviViiRaNrpFiDG1cFk5QLdK9+PIymXbUMLUWWPF5n0NyXqg2Eer
bo/nbkswnAV9fh4uEHP0F5fQsVFf7Xb6NAF225qSGksr/xVGhHzCPXTE1ImKpwTd
LkPQd+suu2K3XsR1XwT33u0xo8KHwdtLPLO7m3bMjqCKBs/0fyJLvZTrFvQQUiQW
+thMtKHlcZzBigd+LhaRG1fU3C8ARgZp7JoUYCx2Q4nb/AkhDsSkBPi1aNUd1Q5y
sSKCBjgME+vg5VNagnGXQMe2mYwQPUyhkDac/iifUUxX0c6eW+oT9B2J/gpTEz16
nGlAu6UQc31lVy9J46hy2wB8WoqpVDLzRyvtyHxkk9ly9z+bKRae8GEHYUklvqf+
WK8s5YUDcqbXcb8eMRb+gWQlCUJvX/t5wn2KsSMcBahxotq317S9i0iet7a/84Ce
6of8Ucin3wZj1ECkLrYGwWrpyBLTK43cY5xVM9W7kT8L4etiIw1AXkLUwa/wkXOC
3pzV09/OEgNfcHo6p0vYntoFXRHYVi2QiWoPv3Y7AK9CmP4NstqQxcOY5WB1vZBj
MZp6eRMW44GaJSo242kQ7ZcSY8CGEbKA0sq6KQbSRx3hJ3K0wSweRMLJOH2N0KJI
v9naBdfD+rE8TZXwEl6qtlufOfcP+pbb8EfoTjMHX5sl37midq2tnLs8bgSK37eg
p9Z9fE0Sh9GFMvlU0gtjU4jY1bDF2dO1zl8Ke19XC1IVFoJ+vLQmNWB2e6xNGIhu
rpNx+uKnP7Lx4U65bCbYhkxx4cNNh6WvBGydkjBVwYgFjwUCb5VByh58mfWtxjHF
8u3hZEYyQgwDw9x7do4Fc5lcEK0OlGVQz+qrJXtX7UJ4lf1iBV77ZeQewdQ7z2T7
zA5Wm6WhBF7Xb24Cc+aiYLk0lt+/jUZQDSXYMTJQKCwlKqcXOBtkOCJeGcdZrkMH
8OrIRIkYOSPAc26q/mP03QJSlp+IMwIjupbE/Gm+kKL/7KqyaEZaS6FyWyCT9TCW
2VtbWtdYz1CgABkfSCYFpLEHvHPTp6AI3GADyhpnsY02v5tKCeoCuIP7mcALmUoj
5B7VHzFOC+4piu3BfKbTzZyE7u46QykSfAhun6QPZRRzfO7pmGbl5RwyYZfxYLXE
SRGzoPh4+DIClHwwjcuJiYpComLbhHNkHVXVCm10vZ98zahvsLx6FQwfUjhogBRD
Td1/VlNLwH2l5z2oCaHKDO5T4V3DkMWqGtmKGYitOymLl6cBIgBxYRss2fWGfpif
dOcZimlAi32DzLMf2Z0W2qVbpdfZSkTvyXTE8PlrGNcjrz9nHvFCE3IrXKMQLeg8
/xAkJaA8JHo0Ch8NOvSHvb3JSNfp+s9cEGSc4Nr8LIB5E5Yc9DZDWmqFE0OVHpuS
KlBpso4V24u+XUavc+L1wadFZl2QlbasKZfkvOtLPOA7J+azc3tKgXP9+BWLsDYU
rKQmAoBIfvOu+Ary12ZWkJbZvrIUwlzzQzYOkG71gMamyx/n4Xxz+3eZqwSVLqHW
0nJLn2bnIZ3zY3kEVrTym7NlSRXS/JM8HTjn48Wgarj2oyF+LPvgnYniDRK1DAKb
KDfgObvrm4fTvUdpOj5U2O85XS66MoM7nluZwkVLZeSYmMHMuJ8CwoXYTv8X9JaO
to4bnpTOKotemw8K0Ybkzw1bnMn1N3d8swFrV5k5s0nKK0dynN7FmjO7zKGCeqqR
Y7GoCPntH400SSRtuqlpxJOBi2nT+DVqVBCe0FNFkt6DcwpBB8+lUUmpUpB5OrqL
l7eNpaE+Kmv5d86iRu0dQUc5qSGYolXN6EkyrJ2Ja2ukkXUNhsMy7e/SYCW+L9DX
gU5smcAjTCHXsS0kAqXN5KLNNHBL2EE2+TGDAox99W+Rsy3+kznlcVPph1WzIkti
jI8UJNpVaTMu5p8isT7zyQwi49yM7/qwRT58cIFJkLELQtAL2vpTg7hHLP889MFw
lFk6q/KLNAys1ZMu2noENXQP8U6nErUjJG8kLg/syF8dUbftoaUdD8S+58taMEan
qHxhURjvdZQGj50sUyda1Kc/+3VWV37pTeFVpO/sGxbvYNnZHivAuubLbe48/Cnp
C6rIFbSwTQtEwsAEShDHQsNG/1JFGN6493BfES8TabkNkg6a/K56P+/JQSCl6NdO
aSuT01nQw8HZTIUS3mo9gyTJr8Xtlo1VNaErlKYxVBL9GIEv0g9cSM8oh6cbLHI5
S7jVXfskb16OZZq4UWkWFc08GbghmYTyXDg4wudwx8Cv5pey5XW+tE//yW0wpwlX
D1qWxpAtze3tIKppZRuZbFyTudY8vL2AZkUjK7SF0FxjdTxBaGGTSWZSozOv0tbo
vzoZBgo2eBd2VH5EJm3mYqQQwjO1elBHesb4kB7WI1A40xov0LV09c773AvNC6MU
cTZfOxdogiRCEbHP1qE/PGUlLTw2chYx0wIQLTsh4q3V8hDF75X+5I9qMa0q/pXN
wHnihOLpppRNTda8gOujS1xvUbW8SID1pcgXB9iZKJ54Su9Nxta27cyC3do+lWw4
IoRRihjFzHUG4AjVmTWmbu/BsJzn8mTmujnVNBXSmbP+UTGWr583RKSFjwGgq/JG
elsPwb0zMlMLSVxl6YfPx9TRENiSuVkIjxnhA/1hV09k4i5RKV8/n2wnuCZUzR8o
L6ep1qBlIVGB/3uIbJ6cMHtThoIid8LDiHEYhui9PcxxNNvxL3r/nE82ySVjnVQ4
ou5Ci/oLqhxd+7OfkoteYB/zLaueOdRn3BT2KZzRccvZrAraq3857OdAGyNx29/Y
JJ+myuvd1gC2hnGsKVabwveATpIHu4Mm1kkgaiDcgtjviABI31mG/HQnFNneHEmJ
cXYCl8IAxnA+kWU5eWJLS5SagGbZU1B2yXwhsdWx5DYNrpVcSvXjtdiLcmPavPGD
fINNDmojtDZTLpA3DsSXTSXtdo0NZO2pNCh4pvQDS6oHIDTE7VgqkQuQs8/A0aPZ
ugnq3earDaRCMlp4KL/XOdD3THkWjLJlb/nheEBMiYcfI07TiHvsCgUVgR2kT6eS
6Cwy+nU8TM/tbsk1c+ToF5EJ+MstJ3n8o0OYLgoS00TGWvg7fqKEUPZ7wUsG6dRn
eaaZCFrsE2/PlaqpaJPjMPiavrSvAsHEp1xnoFZRY/0soViQstBHWso97vWsMOSN
XjnI7Z8Vd/z4SquBIQmhYP0d1kf5cDNtxISv25CQ78sm3UTqpq8rocYJouJ1uzal
slvHoGkdrwQgvSLAzv5NEUk+4midYGiI++TL4NY0wCWqOjC1WUhWIDeUBADlNnEm
SX40Al5MXp6NcA/oKtz71UgzWIQeT2Ul4ksU9bnV9uvvFYC1Ub9TlYfCiomATJdr
48Wvpmyt2nJeaOIL6g97Lic9EcQ9LHkd0EopCFireM/ywmVK+IncFnvm5/Xk4ME3
KZ/q8y500oopgWqpKq4XCWqsK5Ixk+KT5KKmdtyE1RDdCdzinXn/0SDn0A3HvSQP
27sOECT7UXyuPRgvT/lhQJInZyP1wMWoiIk/mG2QdDwo/CIbcnRhfwgXmFlRjVVd
KA7Y6zJrkp4eso+T9NqZhug/Ozsttza1WMRShW3zSilyTf8vzIeg4uttR4KsWTVx
A4P2H3HEQquM4khvXWUphpjuI6yPnA9ZJQpfmKFcofMKD76Zpp6zvCBBY/u6WkZQ
09kFszg9ZOTSmRoEOz6gAPg1LPuCvs6ihXF/kARC3ibOV4/kChgBcJcvekgiIpMr
8sUVfDCcKZ3RN6t8jtK/7X8CyQnqDj7h2jfbkjAlZ5gcx0W2T6S1yEIwOvu3lIsn
aYMwI8uiN/wY8TPmUcfSIKKOohMVYtr21Fh7nZA4iZwv7KIZEOqVnbRRz0RNqsBv
u69uukenUNRyh5uLU54yzepV5+iIDKe+z0jK9eta7SEdp8+cM+WPM4QZ81OfUXf6
nOtSC48B2Mjyqy6QxFDnFrG85F9lNEQheaE72yGAhhhzaZ3Zwzk5Q30lqd08g0Bn
ChHEmQ3zY2jahzTfPCfOF/JqMmVu1Z4JAsrxjk+HndSbgjIXf3z2/VIMP42R6Get
jQBOOKEdnRx63VK0zZ61JY+ec0/uU5GIPY1kVJoPmjVbkaZqWtm/LNBXz/sx4n6J
H3JW+ish4lLadrC87Nf7C8kh0HZ7m+b9LnH9XjhLCUBCXupLssPAPU05HKUPP6nm
S+kxxe9lbYneCgQhoDsgTORUkopVcjCIWpCAdgnXd0I0gr0zmoQY2WPLLJpAyOMQ
Ttu3D5MqqjyE64B5XOSulxXMxDbaDv+U/HH5ugpF7rA6jGfCtrqVGSuRZWgo+eN9
ZGB0mg7J2BdqERHItHUNmGTtgdy4CqRhQJs/relehYQpYJ8R7Rv7xaLs2AkUrzPK
+TmQlbFk4toEHjnLniCVLiUjPN5WelXQPPlf7Qt76Evu4XX8lB6Yo/BCAeBscAI9
NRLtp7Jnmn9Oz7K+jY7dZR3dGVg4W9gy1OTw5w2iC+JMsS+Di60GOlk2lCdumkJ9
mLp2+qeVHf72wQexuuTNGHPcugawG/A8ykBBpB4yz8VOks3Rkgacs1KJNQ21VrOw
JD+OfjbbTU87e66N2YwpbugRWSVhx+or18ab1O00Y27gZKe4n5NWz1ChhOpoWc7a
rH6J5pw/qd/cTNRfAqXYRvOnc26hlMrvVmQ3SlYf1mCm/E2raDTa1wzQdUUI31RK
j4s9NpoH02PY9J305miVhBg8G//LPPnBnhrEtskdYqNDIlORSrnoIzRnZUPgWWl0
vhMxrU19av27Yd5rgCWD+wxOyM0ECkoeqABkhNkXXHBIIgqvuPHg0dGZP9ZxORa8
LGPNLbLWhFx2/562UfTKrOGNSQD8oSjzKNaB/2uZq4+Ze62pI9HceiKidSFStty3
Yxd5e0DPqccci1pmCfXFFhglq++z+/wGnlpnB5CRTClAVYui6TxncwrwpwE5fi0G
5DB5Izd0xsS/nWSarmQnjWXnLVJULW+oJzAT3h7K0u5IeD64I/2T/BF/a0YSsW2z
MAoWoqJfidqmJcN7ckcW2ZPwtE9q0TZXTiNSuUiv3E84erJeeyVkGxjjQRQTqKUh
8z43pjcv/JBcHkwH4MjQdkPQBmPYpBBz51QJ6u1QyJqfTzdDX7WGvYfV0aiGZCdy
6IJJJOz05MCQpUTERpqwtrfu2TiK0i0R9X44eaxLIIXqplJ6B9UFqFB+CurawtVk
5e+AGQ4RErlgIPCNlAs6rTvldX4QbIFScOYbZiF62me57l8sQ5LnccQrTuXQ58Qo
w1EtYzKlRh/wVjCChQykMOtSkF8UYFKdmYYTU1pjIowJBbFMFu6U0a505uO08hzi
yUGHYeWncDSZ1E2ak2/9C/1pS3WcTZMxewaXOYyEgG1Ou/R0cyxf+hbrXnC1ve8s
kuKNPcTujhaO2j0iCKY3md1+Cge1ZsTSCJHdUeFrLNx2HngliePFii2DjyJvuZRT
ba3SKzeOjnHpbmQ0GNMc8htEIrS60XC0KznuHpcNd0ZGP1J0UrHWyL2/TKDe+9IV
Jj2cVQgQfIMJkjscrCx6xZ6DNoyJKC2IHYgeLxPg1iwn2uEMWfuSeFkP25T/uvxl
7glT3YIE9UtFVPjXTnf/mYg5SE4WaxdbOmO9FcSvDWUiJPhyDz9wNWvuEbnO3q5h
biBIRblB/aP3c/NfA2+ACpRV0KMNxReU/iFHRf+OWnq1Cd3UcMp1inWsFUXyQll8
yL8YkEAPv7rYdG3MCYF0e1wEKhtIgVVCg4mEv/ewjtk/R2xsW/ICUWQRekBjl1kI
H45uqzrxNsrWbLylb3wsY29YssS7n/7sKMmLEZYg1ruTVjesjvUm6FZEsORUgPXP
+iuTofYlsjDnQ7NkIKIlKN4ERY4BRKiuK5X4BVy5//uZdyfVBnibhuHmBffodaQh
CvrmzFL+GqQmI5xeQxBcD47O6FH64+rtZzcIKSWHvqmPnngl6a1H4iii0QusloqT
Ztv/Ny8AfLI/IvHRL6H0qMJ3o/mBcWJuVtx9rKdYGIK6cdmuZw9PTTz5ulA6zrB0
XHAQ7zclnW7HTfd4ZJFp6PpbwDy681y3dGs8g+KFRaWTMMqtmvzprOVFuMiJrcEM
BJIJvnlOF4r2eAEo2bdXQdTqdzko6pWH9PaZ+dLVxjGebe9fBcMzRuetADepjHGp
5WktMTpTliBvnfc5V4mj8WJm9cmC3q/sCRp31k8SFIvaEYbkozmxMjDwT3CEVOge
J0v9tKlmuQwU4UfkV+CLJVCshoiJbPSk2K4vQlz0jRcxuUr942NVZGZ6X39i+l9U
NaD9Xt7uIXauJrP/wrMxGAmgbkhnU6xkP6StuVVXdHe57+wLeFUVmgf7Ke8fqi2o
qV0Al1PV+cIm5CMBqxUjYHKKQY7DWox1Q2hKF8byOHLdbPDl8wUFtEmnrHj7l8Br
mFwRsB4s65v3/lU58f6iAUcUOJqBR9f/smlWXhGaVaXbF4yiXKodonNWPittm+zD
eM+uF2oEwd6rTKGwGbnYeOoPToBhmtQfYzM7j+XBfmeJjT5H9FXLFW0SfQj0HsRX
k3Sv5pMDBb6xlOaQ0G7/f07wRzMI9yW/iLjTnD12wT1B+zOgcnz17BMCSvN9MtbS
fzQUUpZRC0a4jgXuanps5JkoD1FsNE3wgiPYr+Iq3GvtT5GxxiuY30L7Fzqc4uJU
gwONr0bU2revYBnQor2EbPLn9dy7C0QFVbcW/zL+tMB/2ezPK6hBtHP+iFI0uJOt
ZzhJd7a/q5roGuVW/82IB9vKiapDmkSRjV7c0551Skz2xGKWyrrlyzSGj+SkvXB+
qc4+dkFmHl8/ugXagFFFhS0+fFoUiJbkUJVFljS+BHvWXlo+rzBg5boxo2tQF3CY
xJKjR5rXGIBHo85TorN9cfIR9gdZSn2ilFLNmlgSdLWjj49A+/flALz6TlGLU8ow
rQs5uC1guKrUz7BXXTixcHtxsbFCkg5Fr1YV9+znVXJ7b1Iy/pAn7KkpX/2Ajejx
2Npujc7R1PwiM3sN/SbR5rzBjT7JqVvSujMjlFsG2ukiR9Ghc1UQPeU/bx3PZW2L
bI53GnzqrrRE5QE7eMEm9ZsKDL5AytngtOM+s0TIXVCeQ+t2TDtkLAV6e1i3RKQp
0lkZ8cTyXSbenywYMhcJnmTFFZpwyajxX2L7V+DNfTWRqtqXibACtGM8c/v54j/b
umFyjLuTeAhJkqkp6e+PlMMZihWU0+6E5mPL0OqEElyx38STWipPC/5OGW59ZBAP
KCxw9RUzWkZkTtXuaKEIrPZM8Nx8jj/X3Jn//aBaJbRdzwZQkm1AtZDKJgRa5Nv9
BLaJo8uVwHu2igN1NmpefHaemSZ2vh6nb4Fwz6PNFgeP3HtW0hHD7r1KDEf+Rm7y
0raZpQVPeG7AS3AwwxIAwewnl7jWFn8o1JTvfMqAj0IkTeIz0axevwBp3AYBjxEi
agkNWJKHC3V0YnCMkaeu3p0UlYrj6fyob7hujZozHZ6NtsRozPmJOOV3GsxWri/x
PWzSe4p3d3ZzCEs4743Dhet+UHMHH+lrSe5sr/dQYaD/SkUgV8aR6Qd56l26FKHX
MMAxG5a5G7WLNiLtNYX9J71NSbbIT1gzkSQfN6Wh20WJ3ig8EvG1kv1yx+fjA8mN
izC1ThX/DEanG9oPzMjm9a6ryq6GKvbh8VyuvcsPb4rAWdzwydiQxsuE5R7VcTHQ
emf2WJ7I5XgpzMYJE8EO4S7HwB7hA/Oab5pM9rocyIKdYtskZvaw3DeSfNvloCVy
TbyPvxTL/xOhIn923dKOcjkGN6EYstlYPKDxQw5V6nKd994b2BmSoYjLySl2cSxv
8u/9+2tMaNWMAyWX0dbObsHu3N8NJWl1G3+HLoDzTU3ZIpJ3PUQEsBBc8uvekmQY
kPAPyIlA0E+izbXleQbY6SmZa9LAU6ZkuXnlGR1anJj0VoPut/XUq1V2/42o9uso
VRUShRWzR+L485NVZuLIObvD6JfXKMWPZ/C1JMfhK0aHEOllaNpAkPa7HL7g0rqe
7wfORUGU336HhCVaAKjPCflgefbZNhQXc+aaenaULAGSlRy73ZNAoueNYbJ593YV
hNu7wUkkgFjDJg3bdMRZ3ykLy46cJ4nCIocDGUXk2Dz6/CtAXQAfaqqZYzF1Tbsv
XSaOABAXwYkPBb5cBFVClXUxxS56Pvu1GExZHqYLvc6F8DS6vHFDp6/IjnWViaYx
LKa72XhQx3HCERBbvf7P5VqN4wl9xkDenmeZSE69QHJHEUgk67WbRFRPQQt57MDW
Y94ox4mCpN/uQB7vANXTkq+dqoemJNeBvXe1D1nNa7/T6526XmAv47DaQGKTXjHW
v3ZXLb0HZCM8xnn+Up+SZ87JVoBXx8HQvEspPWPaZMsNtSNIC+mFr0ciFbPH0nOg
vITrSIAPJGIl0NYf4vPXbwfqp+FobfQhg7xW2QV2Z4bVrRP7yqVLJr8rEcJ0S3d3
db/vTD4p/fxW51jp/3RxwX7m+LyCLm13jRhwALg9vLh4PeyIyT70E7XPekirTneS
jhxXpjBUz59nUNlif77OSNPsaNyQ+XebbFKVvcphj23yy5WqyBd2fDVItVAZCjhZ
kZF53ivX5bYDEaL/pJuMXknZsIYeKpnkXfXPjqpkokPcQVNqkj6JZXsGYc8SiC9f
omhgCmpOBh8Y1d8cH+m18vw7WRThEW1g7I7P/pRcNHNg9dCDUrGr9dfHPBXlvP14
z5ieI21GhjXNGeVvY9hN60V5fCVJpOgoEHPox6+23+HpGOkqFwvYOZD/uspdVAbm
+zRvPnL7H2B996Xc7hxqn5fuUZ80NEAYCDAa3KsdkvV9wrkPbpGVHvJ7ItAbyacI
lVShtrKbafFpfDvl6N8n6g9JMFzTVhY0tPnK88EVIxUl7G81AvLhxLYFwbUWfvia
UGIc0GrEaaJXRNjVFM6tehSp3Z+0HAONr/1qiAD68JOdgd21YgCOW+XM/qn8YmId
w3VxNpfcj4R6X/GEC9gZYV6+HBb1wITptueuSzdaz0/M/IpXzoyAkVry48UVhtsd
lKiur8xI/mfRe5sEzZPkBrvnDcaZSzPLrmIVhyXiNJdEDGidvNv6a/GKaxL8nRkz
nnaoR5jfcZ7pZm8kGI37DFNmP3X8qhLl+5XA/GblyTNbnsFYOSDSJCBxkUAClj2B
L5p/xooqHTW3rmFd57a+dHneDcCJZCFRd3grFSMhKyV0CXtx5Z8Z+PnfkgOQshHJ
vuDUU/ZfW9y5CPQLdixdbvMo27ANwnzoAtJb1cLUVgW/wKT0ZWk+Ig2c8pIlNMCX
CilivYG0YFWbbZQg0C5TzCC6WXnkH1GTajDlyxO14DcEBLM8Zrn8wXfwIhI0HqD4
XFzLsiHp0jTXFNpG7+Z0SG8/P2gLyiUQTNTxEYkfS72w69+Soz7HqYGFdAwwNjGa
e4X2BQZ81ZMLVVIBFGTEraprlI/kTacc2NSVxq+I59cnkYQ2wXrCaZushY19b5Ni
t1TdwF/NvyT3F5+e5ym5J1fUnYwmn2Z8J0bydSQzgzdZ946IuFSUcZhjs7pCBkRm
FtRsYSi1+B5Yt5As8eG5ZwZkKL8tTcNXszSsvlr2ZXlXlbrJ4cT/zi7z1OPmp2oj
Af9H+WEOSFiQtrTLeT+fZ+mGZLSB4X4rqUgNu+xovZCTAgjs6VvqtYw3vTnfnVD7
34sUonzz+okLuaeZquAv0VtCfFQmXz9fJPuYQN6wWSS95zLe7pjuekTim6sPZYuh
Z1blTVrdhZ96BrZ4xr3obn9SBNrP33FUyGfdXDZ8yPwFXv+Qe8ef3D3i0Hrhrd0k
8b8vwG8PoVFrm/6XutC+ZknggATQwfyr3uHeo11u5If2zYzpI242zSlPGgZZhedt
bnyBkEi2eY4mjk65IYHwyqT/beNaUZFFf+nkNQ32sKrZIKFqOMmQiBqyc/JmO7Bm
QDZf2sy4vQgZeBSozT4yTA1oR0r+u7ECHhx5QHZ9ahQwTxkN7aDnn4VejxLvDieC
zjLGes1vLQ+3Qem2Zz3tQOH/sJ9b8xz8yiKa/IpMXm+w8Tp/4QFT3E6t7q0FWGZg
8PFalV5kfTBcV9h0mn3PCF15sW4eMYBLzFnwnUhZGbp3gPpzS5Z9WCMcOlevqCSU
rdZQA+KXSCVMU3/pjyZSF9aBLogJkiJKWkOJd2VsxPPkime8r1D+A2aKGTQMGzBZ
/yMeiYVcEWsCG3BYrreF8hrDXiNYDeQHdjPMjZ+UdY07ozx3CiMIrobWG8p4tNNI
gNEJ27ehD8+bl8s+ceK95kFzGG+TVlGCmD1whKEJWyuQvBX+eMIU2kdpZg3aOFiV
JMjg52m03uHsDYIV8CJ1pFdE9HTtYRE5pP7iWSZfKKlp0dYwFywqhcTcASqzwZqA
O4iZlWgyJTBa1Xu0yqPk0RP991PBj1/KMF2wR449fcJJ00LFkdkakZjBCezVk/4s
/xeFJ1dL4N/LDuM45P99yVGyf7rDXfnNTS2JtdsqKnyBDzfqynWuw+XspREndvVf
uEB5W12TCYJ/lsoBljo7wiIoplhr7LGsMYSICI5dp+HHbO5ADGBK1CcTbEKI2isy
3NPLY/LHr8ZKgOTfO0AGgBEulRWf2ceL5ocuGqmm8Pma9q/LxX9qMSPP6bT4rRDq
RLoFzul+lno3KblECiXTqrq0UWGr+fECMWLvwUs8WhY9eTSEGk6NpxLrXRs5JOsl
8ag/YkUzN5UbhlGsu3UXl/nv2WGxYIbtjfHEGgqa3PuYPoCGsGXKWko9gd8ac8Qg
fh/s62FCMSOZvCg0o9kLCjB5vUoYpKu13+EPd5H9Pi59eQMnfQm8jolS8bTa02GF
gi74W7szb+adGO2mxS2o+iXBdyOHD7o4jzTpgBQHSyeJzu7LVETm6heFdQ2QyqfA
tizupHRTlna5UCXAIF+HpR3pBL82wwmDX5CKYehPx+UbkP6wN5etlFTy2h+//RVK
KJAM3Lr2rCNxmbT7hVpu6zdiuvtehFVVuV+O0q0dtHuRjfr8/gq0gor34hYJ15Fp
pCkPmkVrrE8Q2tEhAR2bqc9zIpVk4RHuX8CLpGbOStMcHG3tSsGp8bKXWgrhYa4i
DQl2IiKC3tlycVFgSqIxcWNIpa/TM/zw1V7wDj+u/DtGAnT/RL7v3muNfyJ9RQmi
RUXBd9Rih6T6YUxYzUIL0DgcglBpucL8POe7FIQp2yaAHIiwbvIf3brCYC9dTcnK
xzfeRIdqMai/c9CxEtVs3rosI6VOqdBarDSLUfHlUKm7+2rSX+2TKUU1BVt3DZhh
/ubvbiHE8oXaeh6f+lllFKqPUEMqN5SIIkO/csiQerzauVrkAdygOYvtATkwichC
XRH2GxQ5Tm/cICSH4A4SvqpeMDnGeIaZKTeFDh4i34j2g2fVNXROer3+La/n9iho
Cdcn45iZ/F0aT3xMlocD2TX4+uFC834t9PUcaNkDchmfe/2w66BnBXUAnpkzBX8P
02Rpm5hDZ7IGnHuj/VfFjLpAJUCnYncPpbo6GbaF/NjNNxPVxq/U8eXE54B7gMSu
Mft8p4Q3/8WHCIyazChnbCtl461/gsVHG/DtVVhFJHjU3qyRuTDGqlQtTxFKRiMP
E89uD2/1rgL9aGI8dc36KSQozoppzLj8rqkPLVSUPZxowZubuVBfzxbvrAYv48sl
rhkHGLaPZs+TQX4X+HhKWJR2Ze9nYnENELFGdj+RsM+RIXwNny66HOe1+dL6BhVs
CI9SbDTWk3+oKe6ZBjzrpRkviQFx3jmA+BcCwi2w8AZaHl4zbSun22Dd+WNhOkPr
XxZVjDSX0Sua62CAbvoQUkoodn7Sn9GVel7possc4GoV302iQu1zsKwYBUROI5Ab
DD//IiUPWBmo3xCta7D4vKClyLajfQ5C/rFNu9hBRztCOxbPynMvcGGdpLdbJFPa
7mlUtYl3inS7o6w52G8RMJAB4mhAJThjnJhoA0WefcE3pj2MqdbTcfNyWTUgnWSg
fHRm2PpbLD/BpE93ICneOh8g3YUyGIQ/4V/9+A4Gqc4zWcgHDQV5QvY+UbPEG1sa
G8tr/vgem2Sr2u6dIwXYhCV9zGOcda9xCJcbGX1Y4KcyvVlIvyhRQxMyEq8upttz
cFjJmfZeoqMKU99m3zdpctUdpPPQI2SJswY9LviZ5iOhhAzuvLke1upmGb4fMzlP
GJsNoQyJC8dU81cqwSnP+Xcct3vl1bhJtye2K+3MXrnkMukMSW4TwOwwzjp4kMmA
y5Kbc+Zgbc6StSzxwCglaRIhff2E/8FhGAmS07KNyOMkT7dJ3JDTAvVLX0pgCRzP
J417If1GuwaBz9aAlvgaf8vYbypTq5nJsKc7yjyP2ZBvUU2WlNE20ty3PstUiDdZ
Hx10zY/q1Pu66cllA5F4tRqeYz8g6ACNHDdT5K3Tb3oZ9qAZWh61JOFRVPt/Usoz
tyce38evmmmmyikhF0VCTs8ebMLbhRdU/1GWWPNhb4/c7kS/WZxHtr48q4TwUQuD
R4Pq6SiawCrxt7lETUdl4QiFp2sSgFvs2t4k6bwfOx4tnP8MMmsbCVw8DaSEhzhV
FaZKCVkHHjOIlWSmlJtnggNdP3Pl6oyQePFYBAafJEIZpPyFpSaXNqrqRaUg9f05
OtKWkCWG2IOq3pYdlsnEAUeoRFhN8rKp84L97SyLBPrHYrXxmKcMi2ZIluPBmSSn
10P9n/kUjLtKyM6kzioNUSDuLIaUNiR1AI8sSmYU2rj8idnGLdp/AZ7jR5g1p+mO
lmVxl95fzu3TwcPXLOhLttkZw1sN1XeF9avaFn3hS9hoDKMmoM7BZLd/kpjE/hdm
YXKDfkwSRb4OtpwQy2h3D5YWn4pznAVcXzQN64pvn9tlMG60FW8gUgfwwsScgX4I
7j6S4oriaMmUw14dn9fHF9sYd8DILXrsGbY/v2dJ40hKMVpDRCGc9L9gfxU2PqQZ
7WtgxqjeD3P0GFgWUjQlD1E41p+dPNVI2o7Cg2Q4EnG2uEVpugGL4FfjYgyB460l
xNPwji+XzffOqm7hl7SRoTkcDBRj+cHk7LasFDEUUFl2jbK1K543jX23cBzigw7n
KbS119HnxuDzW6xrMMGOZrg4TFtUJyIvsh08DVsX7fIGHCSlQlUrmzfYITvoFgSX
gadlR6YTtnnpqmWZDNI2Tblh+DHzI8bs56ZB7UIrlde3AsHyFrSTSYlNP0ZgUF3S
EPn8GpTBWwNGFhQPU5FZ5Bvc15R0br4Apr3A9p+EW+o9UHbtbqILt0H4+yoe04ta
mFCzPxIbCvh+LnQ9T3X1VuA06myAyairJoz0RSe7kxB+V06xWGB9AHP4xrfTaDi+
bxU4ibZLkeN5fz7Lt4VKdKU12FwdzA5OkLTTsKDp4UcO93lwdmqb58ny7Kscy7+i
2MiKueB79nSDSEy56kBl9k1mOrpBxapSIVXlnmIYpcISpxr0wm8NSMpj/zBDu8fc
7H6tFbRmdNjL3/JSrx6r4fRJBeb2wO1rtsz7zKpWsA814wZMskd0GTcdvZ5Pnfp/
dpfUw9qbExu7IuitbCrmbBlhekeGH0pXd/14/lw0/c5UyTP7UamkqvSMyAJYb3kJ
c4c33DuivZ5MM4GENRPRi160UTkQ/fZpRoV5/P8Y8fHYXDF4iWp3dC80kbRAKfHB
+b2tiaDnO2zWynKNkuohpOKQT7cIKB7rPydXMt55Alxt/+XgreZKcXUzbkqXUQ0d
pJMJ1KtSh3bndZpl5PsZZC/RlmbMltP1WM68I9AMpnfGK5mkpylCx2nC5UIUhPn5
Xsm9UUvmVgdLCn4d/IgGsZPcUMhOm1tefQFuRs+iRKGPZo0H7Vnq/lIlXrcgw2U8
VLsILSSJ1Y015b8qYlAH7vUaOL1hC3vdgLyY1qxtAV+xO0eAnv04rY45qmsv+UL7
zaUl+0qZkp2mqck5wOiUCiyM/i5vwHH7tCHjw9eSJT3QHqIXdH8YpKeYr22D4ekM
D5MSMHKV+E6XQqjOhyCXC1KQk0Ro9u+lN8CBJt/WUCaUgLrfyF/bub9cWIuvbWV1
n+JSxUGpAcMa7Du/8x9vrE25a4wFRUDM9M81nmhhrfmSSfyS8DJXVvu2vLnlntuX
V1OxRFjl8rkfuULElJgbfGrWcGQU82mrWvXggPZ7XWVFAjyQMSFBUwibEGVna2C2
73Xi6FRoZTszfoLNJKUsowX9sXuwRE2+m0tW2ccmrKLmDYB9Dk1B1jidvEJNzUPA
uzRKxWDrZNf8Y+me8RjQUtVv+iory5LCGMfWKm3Wn+ToAXVpCbhgEsSzAJeIsxR0
/hNtpAIi7nziYY6T5SQIPhL2sWD+eYwxcamnjBBNw2ZN4ueRq24uexqlrwQaMJXB
Tmmf0Mv/W4iNO4r9DcyVBHYW9OlwbtN2oUVlAYbUVhauaizMxKYp+fMGXKYYmMk4
QCJpLpqxygiAp9ihZ5w4dPwHAFQ3jRCKOI0PRnsiLLDGMfXOPLEIQXyAi9fCxqZH
k1EYp33/BjNW9AGoHR8j/pg1wS6Ky0nGqM4AA0G2lTeHDx3OTsqXOQETYCZ4Cggr
zfKbgzh452sUyU/hpzv3B0A6BJSx42tN0FaINx7iT+On+8OeY36pINQzynPFvKRF
NzxClh3ymaHVxphzyiwvJYWtK9TaASjEBYW4HXToXBMKvJ/oBxDyYyAE4Vrxdfdw
7vk21GN0D2ecZRSaNuQkKTREjM92KXEf99v+wSQWAI7lp7nFLDyLZXbwdRAR8swS
2F6rt2CfjEjphxcYlBIe0zPc257Y6CsAy7O3ePZ3flQ7bbputzxsTynJLa6iUBwg
18TDLTMPQfwyJBQS/ElRg1AvFxA7eQPoeYpJfNRUV7MatKP3/0KXI0t/lC8nrPrA
r3GQwUNPC2F5JA1yC0fxTcjeg9ZwVlO+TNbo6rt6A+o4UFi9Wt7WQuRC9nRhnt1b
XrVvqnq+wKE/QsZwzqZf08hUncsFoGtgjIIQsRvNWS+TxfXiWgFD/1m3B2NnoAFG
RyiIPQVY8zb8LP9FmguZ5Mcct6g9QIIMEbKru0ytLD4SZsA/sNuDZm7Qc2SIkRvX
3ZvO0FlF+XbExaIFGj+n+nl9uT5U7MhnP0vkYVcpIFTbasLS/3izCAUWRRGhId6J
P1oesmCmOPMAisKp0T/nywv95QEmIbTX5Z/+R9FsUr3uqC/THBxAzGfEJW19sRBZ
afaHTjZ9rqNjExP0sHAn1dGrGM3mOJ8VKP0jdGIz/kUMAUcN8MZ3P4TVwuYvTXEo
FWGm0u05ZqtITDCO1aOPnDsSQ4jsKNdnkO3CRJFWMyP86rKJ27jC9hozPYcRqpWz
S+9WXnHrbxkvypT7KkxbCFslUTsUqTJQ+qEUcPEuEFozrNocyFtYU7iRA3IIkhw4
uzmpWZfq7wKEVAiyMS0/QlCSJFvKckAIKhjLLXdR0pOSbW5Chax3Bl+KenjYqYJu
5J/o/LtAJJn3NZ/AshIvNKRqC7Jq7J7+M3Vlk5r7ahfDQ8+s2i47GNRwlSNPWYrn
VF7L8P4a5c8lGlsk1m/+EcL3mEmQ5kccpROZCKh7NF3iyT6qY9rYKp/2rH+PX3dW
67eGC6nxOBekOH4MmtRf4xmqiWxPhv+bVqtJ+tb3wSRGf37RonrlypnkVc9heKcR
sX1WdDnX0wbiuPpwO1g86WLcKflHXaFKs673GJKrjg+sMd71/QqPjvRM/SwsLWte
3N+4bnd6v/ET0DyQ5xnnR8qZgztzoswFXOXzYglaF8i2XTyzch+mx1hOWO0Aw76f
NBoAm+EqVcvGgWNGM0bUf+p+ObzWQ7HotBt17JHFu/8mujMhyFYPZrVDBd8d1VJt
zZIFydnTuuSYtKIVIImnM/azd+e8UaYYgYO+FFmCnlJlq4ef69DlE0mp+phaeICz
JCn0t9Y8OxyPF8EDGaEMLFUsI2+4TxDrWx3t/zUz4KkMUmZO4+V6hq/h0+KYa6sU
soMGdjHbXRPcGmUknW0WYMRaZ98rtMPkvq7YX9Q1TLyl9eFGMoMzFLfeORiQu0op
VAnfrwGAbU7BpKP2PUqa4k/JQQXTOJUHs1GOGQzhP8medy4YBnyxdFsmGMX+fFzi
BQK48ZuQDlLprAgXX/VYyNfLKhLGBNQVmk2+s9TQt2Gpzzup76Pb5IPdEARClSc9
2tDFMalFBoCV5DTrkPe4hclJZDPMjIQW0Zr1PBsTav18lPBiUSTq/9GtTRirFYMB
shWkzjBl9I0x7bUiNaIatRfVR9JAjKlfSnP2XXtXNZOL3+OldYj463ZDjsetvXH4
nZu5+VCTWHQu7rAponsjtzCpL7OG+D3Q7iZMvv8GiuaBDK3uLkd5HPMnWvue4zGg
4z2WgX2rRrPnxZkLsk16FAAJNoLuigqIx+kiIQpLWnAXYxJbnHKYLsxviJ9sz1Lu
5B/FrlnVoWCgLWBDY3hTK0d2fDGMeVWvpwl7hcmjzyZ72optxdLximnI1Dmr6oSk
mFfTncdDb+yqAi56qMIVfCBFfJn/9bhGdRpSLUSXRsr9Krcf6IWXKPTjfn41CMEG
g32ZeJrjFLKzq/IYZY0EoecLlLUqEZc2bk771jFD7HHFWe6v019gNqVU+OQhpZBD
xJT5Lt/D04avlW/P0eIipx0ISLbihc565lHj3mcLfxW+KMeLsBLoEr7ZTE4HL1zj
SQryne7hl9gklo/Zim5Dk1ch5hlvUQsv4BAoxoybhhcsXbkKa7xykyawMEuobpct
BRFUdt8YZRioRwYXHopG3cCLIBersKJ63CxMrrV3/1Nc0K6paptuZiVsApKJFUCw
ZCQybCPrwQhuRgMmqlcJeXpcJLToO6HnJLs2pcBu9XKRHA00Dc26ULwhQ7r7tkEP
kyevK7McgTNDtgBKBPVLHk24ao2gysQAr4pmkUjHI44crpFs3gYIzqrpBhxXCaz2
jHsQjoTO0Gr/kkMDXMp7XLQVGBL/OYKs2SSKP1L+3vYuwlqCi93LlBIxJQWAE8Ve
BABC0KUZvyoc3rsprZsMc5GKexVLtTcE4m6/hRM7Y4a52Y2Kum4V9MxKg9qxEutr
55Hw6H06lKZA2KKKggY29lCdD0PJIbctI4MHh2kIy4XF6xrlSX1MVLAjF8J/UbLU
MeHY0d090ca3OdF+SeuSgzMSvMlrZlBXqhsntfuP3EW5oEiE7isl1hlk2LUxGh5Q
RLaN6Y1qTNFl6PsPLeII0wuDkMffyW+mphpG8+820b+2fQPf3kk6Uvjm6X9zitNt
wwnLBqs23B0CJSlJjZXMFxeWoVw6rvYRaApfheRib8mUJHtc7TwO8qQzAuJOqU6j
oxpFGDo1Z4EXKmx/3KiSN4RRJeJSc2PpLZqCD/JRjZY1A/oya4iV+A1GQXr1uMFl
nhlBIPXs+n4xZRkNYnpchscLhZ2LyYZGwYlR4tf5naNBFoGb+9lZzwKPsYXzQhoK
rT5I7nSs1M8ruosizn/lFYxUMOxwyELQbi5CKH/kuiRzITyGXYzJEkO1RiUcjiC6
0xSX7YDJC7Stgte3fK5n2PmR1HQFNsQpEJEm79CGuYcnopOlgHbYB6T7nyWXLd4O
E2CNEUZbpbFpkEgYG+X9Ma/qsnJTQXH5Ovf+JCRP/Syny5pYawjhXSbmC5XuB9JI
mABTkrnoGBivnsBJhVLwXL7xUhQr5c7E6ThncwT2RzYfpFqPMlsy4R6kNvBLK4gl
KlSe5+wK+d2igT8GJtmFRKppujBRyvCwgwb7h6kCmCxn4Cy98lTDsnNN7l8UkEan
/2Jsw2BDa9v67sX/JLqAs18PKIQyzTOtKydDQlb9PHx+iHocBOke1sFd8NNPdQq9
nQjY+StuI56x04/Zh+6tQb0UWzK7VsSjMoaNBMCBhjAxYkmt9S9BSsb3dWpmdz3n
bFbxACxq4uNYf5o9QY94Waa5mwdYy5MV6E1GtGxyzij+ZGmMlZNhbg84VfKuDedX
HP2Qp0fZE4nEXVqNHtjvpvH4liX0Dv3vpnRlgysLprfHvMcJbxBQkV3f9OY/DWfe
ulTBUGNjPm0gQaoCzkjVJHnYVSM1SYFGFx7DcPuhaXodh2e+FfLSffHRTNSW5Sa2
PHnTi8ir60wnAZL84N5lpxVJpqQPdoLWAzZij6sdXRAqiJjd4jdRw68+1fRRQYVt
wHD+fYb6yq1jltxklxb2adubUfvpL+cQgT2ZhvFuP92cJf35Ekd6NBkYz4/i+ark
+LQGVV6xMp4AhSKWN35nSlBugQxeL/ZD1M37NeXKgrrY4cdZiZ3/7U51owmX1VpL
UKTwWwl6lnSUwoV98AHdrhHH80BdYNrh8m2NNu8DKUDbUuFqoZ4vJ9sYqdDyxPld
N9YrNWzEW8l8KfndM3+C6UVZsiiG0BOCYZSFfESe/5gA7uqbDzdajtvuTr1BpAO1
QZ6SQm5gTR05qKmuAzvj93sjIshyLkBAIC4O4efu1L9LV2UiOxG5yL5ao/opefyZ
PvpcFSm4QPBdKeHXaMmxIPXJCX6bdSzHEkX5bcaTxUH09qMcYVaMtppmpt/k07cD
ivh2jpO+jmiLXzMD1PtYkTB0HIpSAU4BhF6jEZ57Unyry5cgKue+qzaMcMWqee68
SKAwm+auP9j5dd5uAbCKeZWt7MLGoBVnT6iXIEyOTo83lhUnM0el3nCazcNKuJiw
MxQgmYcbKNdM5PrYQIMTdeedReVQh0menRmJ7/3VIVOlGvy6J9X69crPly1GC5yd
bAO3qsbDPV16mB8nl0SINOSkjd+W6xaz1gaXcesquuJrIKMAwaDQ0dvHtL/6s+l6
HfZ5hmidHll2z5zMuN/cBXlvCKS17ANB1D0sprQyMHu/mfLh1KzVoOUiFY9woYhK
lAdok0+dzEGff3sAv5+nrHo03XAxr0jEwZwp0u1hv7JOF3nXDWJB1PP4eGABl0ZA
1YMV9817huDEC8Pr4xV2eON8IynqjK3IyOdCMXGnZImbdYmKk3iHJ1u3vaML2JMM
2nIBofV9b3m+UboifKLMnufBrL3NZZ+XdxWxFVduwOMOz3PsFQpgnoMkIWcrh5kq
sF5WTDq6sCxZ+EC/YftjxdUI3/ZPbzARjPL5Pj9py0AraObVFYiSyZZkQ8wWVIo5
IYWQmnqXnwbGjrAuztRyxOCPPjwUTmH7YtFaI2fkfFqdRk7YDAKlZsnNTS8XwNQw
az6aE2uV6G+0dU8/MJ25Oj1jVexScxo0aV3leSrrVL8jp+DHwVKP3PZ1L61Z/8lQ
ak9JTOiLmfuZBQMIg2Bm6lK1xrRg6sHNO8fXIchW0SCMM3v9zR7TwT2cXb/tOvXu
jPxR/ZK1tttxqcjYmx+29lGLLyyV686sv0bZF3j4qx1TcckZrFIsnPXwkT1mIzKh
by4D0VexOPowRV6hjsFG+3pxATRa9rIPRyqiwW9/qskzVnd2Es2ZGIOJNGfT5uSD
6D4ErBYcHLD54kWehXldX8VGXAN89tcJ16Sfqcm5MsUYvKwLp1VeufV0Yb1V2ck+
NrHedpRisNGFw3YyBXz1TmLNdjAmC+G9EhvDaxZOP2wqicCZaImeiNCQ4Tourtxf
ur19B4sM0rfLOcgaHsWAupqCUzdKepLOYqzGvjqoF0wOeulBZ3sTm1uFM+2nfj+g
jltVsMKczesZycvdx5UwX9Tj1vTy2lXmFjH2WXZzGG2kVr4V0GC+XKsLGtAKDM4k
TYn1aUEueBNYbO6FSUk0oFcB7goVTac7hFwXMjSITBZrTfJ9Q81XsQYezJN7vUP7
Bf3PRiuqhCF0Wcv273b01iwR0azSZgb3RtQm4B4tYWvHH+E6kzMxlI7WyxJNGCjE
iOAtdxIdS+Ct9t90e0pOQc6t6HEhQJAbrDFx/3ZNmhHftr5u6GjrsWDg228Jbr3B
cEWDCnOsN55avpNacrB1ANTCC6a2gGy8Pt6YXJ6t5hvIHzJ/SBIcsXzBhTmK6HGz
MjibYRPSYRMEDt21AYABsfyIeggGEd9RKffKAJuvY++wH9rD85XJmG6VhRL6rom/
Kjyo4EGbfoBfWGJlp1a85Lj13qGJXZGxUVGplZSWUeXQLVVqiJjJsceCaYEn0pL2
4mxlJcbzfMwJOnp5Mi5VmhmIg2brUJiCxanOPU9o9b48M3vWecS6SqyP+Pb2Y+wP
uhVJM6NC4eiFCRm3hGbWXPSU62lkjK/ca9UALSuxplcWp+LInEfdfoOorhpzNdNK
4znTISdOtryZWflX18DP8kpD0+5wR3wFlziNiuuoHglmqAcp5ZxTwhX/x3IO46HB
7kupf2noenz100sBiGURdHwiV/FWIpaXqypCZMRKLbek2icZV9wrUB2a7V8pACDs
QorbJWO0UZSWs7DrU3ZO/WHPM7dv412Xd8WgLfbq1BYa9oHy08+NM6kagOxz4iZV
icM1z6mKa5L2agaLY+lQA6Jbyw0sRGoISD/BliB+YUEhCKtgTZAPyeNytF5vI2EF
fkKXBAj3CRevxbsiyUha1cSIzuwmZthreQp6jYrkG3bL43WaNEQysafHlmh1Pw2/
WQS2of0Zj9KxCoQKgOpzE4LZzWWuIoD3WQh3UWM2wukemRQ+KHFlVZgWgaUa5bZM
eQnfzf/v8x7zDiVkZZSalmUxxCsyDcyGirTdEVh9HlQEdqFNWxuNvs1L9j7OOJWO
cpB+mLF9EZTYeUMqweqnW+htBpdhmeRa40SoXyVWldWf0XqhAGrCR0CUW2x/SDSc
6vx2wkFYUoCaL6fjoDurbg8qMz/IoVJdd2Sy0eWOaaNovx0ySxWwV8GsNn3vZsCq
25Ux3j+9bcw+UVR+pzmbU9lCDj7h+6MDmRhXWqM2QnEgYS/zIdxFVyP9VUH3KCy2
HAJZryx1CHBYFEji5YASUzfpJ2GlmjHQxvXmZJX+6f4PY7XkiThWinzDZr+JdgKr
ho2ev6xuqbC/7KzThnHz72L7aGJVFvYgz/SzUfaFpZrPwNQ3ZkI4WOYfpONXp5/C
Fc7U0LM7ubRyygYFXSbEkdOh2vZQulaABVbRlTWtWitNNySayp0IFxo5/A/8C1qi
ehynYIrJuTpdrlYEibSCTCBlxTuFIr/2B4Z/1Ar6TrD5wjHEqn8WDIkJhRRiK85y
BRIVTolDIa2XIcTTsO55yCyFParc+IFH4x0Y0Zwimnol588UC9CmGXf+vHGnfDMF
C/JGGJL9IF9nRnJbAnw1oVomx9Za2b84o+5hT3ukcQIWKRXPWtac3ag3TMkECJ9a
we3jcUi3aK3cLqkaPkLQaCsJHfPxWm3XMEMxjc/fE5ZG4dgiI9HoQVHS6UCu6XGF
GzrYtEkLk/OQtVt13XlWh0mqdA3eS3ffi8y5dL/vdFXZdSUO2P2qkjPXriG5vtHv
wczng9yb8pKEgDVBrRnZHWeuSSfdHYU3zI+PZtUMbBuHPgSw5UPU2zs+e9uDBK90
WYIdcuE341GzWWpwYg3zboJlLnorTS6LOtJxBOh4CxQ61oPonzzC2Olrgu25OxOJ
W7sGKQS141La6QUtHQdNT58yQCzzNBSDVsDHY5yRndTTULGKobWvUkfO0raOzJne
iYpGQjWZBb0fR0X3eQcuVm1EZXOFuaXcHm/HlUdrM2s4GEsi2WEr7PoDYP6w4SFs
WkpYidWPKhuRSE8fZuIMCEFSrNlcJEW2gfiRnnjA5YFJJ5Y6EOcHQYYsB3vGlpFR
qlehK34xVQsPCpYewz21D5UsYf8+hD/jEqn6/3ZRVb+xpWGLql/Slmjzv+/HBJwA
2e60jwywNai0tY+u1iHcJ0hmti/r9KiZlMS0d49o5D/I5y8Mu83vWcgBYMO93cYJ
C7/mcu51HMEzLCu7OLBKZGqpkmgHurGD9H6OGwEH2j9HEjGfA9HRJKj2/Yfq8xYL
6g5P/8waUhCK552+aCa0lMRMyT8dqzl4WxKwPsZGTUcCU3wqmLRCHLyYcbFSvFWD
6e0aXijO2T9hEhN/j7zS6KNpP6zsX+b9b2JlUfW+Bfmf5rMrQ33JttVXdNtXl5ut
cpdj7aw+EQrwyLiJZwGEsWIQDuSc9acEp5QEiaKN/OW7SRcZ3hoN1N50xE76T9IN
ahvx6L+BzaYksaqSsg/ejgrUuR8zxqVllNul8WJVtZnxCNKRU79fZk/ezZXo6ilw
pDLuUN3UITT4LnrNcCxF6c0I+tvCvgosFjOMrp3D1Gr7nl46ueuz+Zjw/kcdyFz0
HILVPcSByXvg04iSFftGxT9MgVIMySIoOM+pgfb7CeBgof2rS956NCVxjdFNjO4F
2mbRTT6mjePvdryoakniMJIHEyu0+0sEXnsMfrD8I/IxXxkJ9tikiU00EUojjd7Q
DpUpDUIj2TqzsFdjzT0Qb084bOyPxj4HH4rVUd7Q+DDAbUL09/TrJtzYIi0tK4yu
nOpGkwbICGJ90gfufjQEIgvzfK6z6kDSpGKNeE1dA6X4HTv/g1lECblBipimpvfn
WVbD0p84g8c3fuqhaTvjmeP9MzR9hgnMDM6yVoWaeb1hpo+DsWCl98swCsUcmO2/
dNSNnewYhYXt250ir8iljSGQA26IPrNBO79qigImrFaaJh0Wmw3XL3vVej8IaVbu
zOrrB7tFSr+qk/QZ9NPhqC8Jqc9ThOr2UfupKOITkzY5EL9D/xy+3BETD5sqVaLr
yDvbDLv5ryC+CfJ280NxqpGzJzMYHX+WbSwvoSVzQBbrmIES2NImRYj52QsVANxX
TzRK+bPkucDc/N43JcmjStYHoo4S9fIrV/5R+XCY1yzUtXRfELzKPu3phmCacYPh
i5b7GPbFvNXX1UdBCDhKi5305vha3cFJ8W5lKh+SPiXADxYu0gl2HE0hNQq8mOu2
43oytbrn1SKdVUsJwxIXoduXoNP0punTPAiVXb/xKEgTPV5cGGVy4sDnthebPm3B
1Tcb9qZQyLJYkelXjL0Uy0sxWdQUQjDbBWty4UPy+pmjxGansTc9fQTHI/EiJ8mq
BInN7IfiUhLlD2LkcIVMs5a5L52AzFBri7SRO5yWdjoLgZUnNd6alLWPilKXfWLe
LD5X8xJuBEaFg2C4FG0UL5KPPrRTBMR3Z8x+d4Nb7oB252K85SwEjSu/pBy3MAlp
+y609vCOR+CdXnm5H9yssh7zD+pLxKFyj5nEnRsNX+87rrjFbuMoUTOS511EyxPz
yyN0Bj4re8MM8CUKeqyp0enOrIWBn1tZpCNONI08jE2RY+JxzVmrJh+5AANwsav2
7aTQaaRRrK8A65ei6KpN+gN3FwM8tRtsAf9BgFwzelmC+0XqgCQjs3bsuEXPcYJ0
sAUcxviuEnaLf1TgU4R4spvbvYNs+ZZ9XUlfRiNSmxVZDvC2ZRAglv//P1A60m9E
S7csbgAaCmA8t/ab6auPe71bF/CREq2ayrYFbWJ8cU7kvI68QVA9Z6SIm+tKkqaH
LFddu57+yRTgjwm52WDQ94ciHp/WcVfOhmWzgsvMqt+vTIGMfbLVNLM1YCprQ1e5
nrGE8RaQVCjiuz5zi6PSSiiyG7n7GC+UpIRWQCZilDcdsb+W6vy9HwwbEkVLR5m+
z4DNByGD1w1KnKpB3OTdUBOi85AxrlhbvQlDtDiO9OR4iWb7+tXJJ5GubjBT8q9F
iy0dD83NyaOwbNB6d+IdnlA1LmPlWUucGplOmNbfySzjDKb+SmV2Y/5TYy4ObssA
2Pis6tqoXEfg87JBPcPlNghFQc00p+cTGwnhxmAx3CiJbrXgKDGobGa4ZRoU2Uhv
dKxTW/S7uydg4O+VRmqalggNMuRVzQAW3xXH4GoNPDr34azNQ8r/DbGfs9PZ28FS
DbYUEYVJ7rkmLpwktM4o6vnPhQA8vQwNPtTl84mcy0qlthexhpWzRAN0MXQICZ8A
FeTTuqe+8GNGziQ6u5Q9qg89tnt7EHMrF44C396BgSgeBdYC3rcNayoQABmVHPjR
6uXwdbKx5IDyoWUV0p1xgAc20F6utqlcgQfUERDfNwBZAk5gZhiMxr16I0KKT13+
iq52Z5wjzxwaXGRAShhLLUt4vkr2yD5JMHGL8itU6gH4ktpdcY5mDfnLBCLsiIC6
GSx2WSSwvPIw3dfnu3lPdEDMFXP0Z1MWsmBlVlM8YlHxGhEo/YnCp2vyLPLCeJPQ
5GGXn2LBADnEIVPMEtvrpRww9sRi0PooQgyXgHQLBQPBbRMduuddngNJWDGGtuqV
2O+aAguqz6dGoGGhs1ezJ87w3Otn/CuvwjgWSuyMZOWwITVcSH0ZbiG/n8CwNNKJ
loZiFRd706pcro8/EJBpl/pAIjoVr3DE4eoN5jcUnx1J6rqRLoMc47e9gOUW2Foj
AR/9NCtFE/0T2TdMFyAyFcIcJy2RpWQx78H5BwSUwMWmBeAnrm+yutU2+11BNvRI
xM51z+RuaEnZbwLDgJt1wWacTC6nACopVGXc187hCMnX3l3QzbUdOlquTY0uMYlc
L15iMlXKkqN/0gggDEfOYZG3qpsCAsxMis+TnGnSea/QsRMbh15+CiVcimYdz0eN
eWCadLesXQ68n7PMREh6PyZoE/x5Spz/IfjcAis0wX9tfw6kTgLOmJ9OnuYQtG4d
meXLG1r/00XU0gmsgI0O5c+GGdK51/Z1f9aD/QFoPDT3BZPdqb39chcqhJiMFa4v
0XCKHvtzCo7TQ2OXVs8s1xSihpVQSBzV0gac7Z3JizC31Y9PC1+Ikp6SuDQYyG0y
N89KMGvyaac89ZMf577KHZaFqcVYetNf+bf8ww1qc3qpbwUujkyK5dJWO2ZBhb/g
P26c/FR2zjcVZ9W8mN4g8A+5IMSb90PdT4541LE2nlZINFxPzCljATZ9h0u0+kDW
luheCAykRpM0T6S46FyJZL+svNmGV7Q1JXPCGvdoVbRwe5uWIzAWjXJ0ZlcF/Kr/
WoqAn3SNzc6IFoXd3N20vROwxzXL1ZqmA7DlCrqV4LQQuQ5jZyRqUcuj9G1nDhGN
2Ab5SWQVFoQKfS7sXT3OmtezzhZX4XbiZNsQ6zvDqgpqFHNR/DjXQX5qVIwEXpNs
8iou2DPHXUnuXbZ0OZDyeZdLb38rbnb87HirtmHphbMnG/EIzmVyW8pQwJHINTfS
/NSjuklH5eIzxddLUMJO+RVIuQRyAHNyZJeN43F84JJirv2fk2N8gaH2OnxGzVJ+
ebi4ZwHgu+5aBCPRndUNgMEgysd6k9bE393p34gF6rHTr2YyGMaR3EiXLxSwK+u7
ENHsPRTg8WkJmz47X6mSm9rILTglsOnaKLuHipUobWlMLAfK7p7orFdYpXt8+QVR
LdawOmiG1iN9csdUnLe/SsW5N107lo1ObPyE+YabZEECT80wNg4WSHZiKGr+SGGm
yrJYrd2bjEFAp/c+KEbzjW1rDvojhGwvYvUVNW/sgPOkHBFohh7yQfQY2+3jP2gg
svNUoNevunk4Ozuiubqmd2UQ9gLXVJen4I/LJvNwI3rQhjSzsuaU5fP0ANpaTSbl
DCMTxq6uqW9rLfgB6bNiVZE8l+9qEHPfMj5d5H7A0uDfLipqCv/lTucD26ly0NJ7
LkLQE+ei0NjG1h0e2toBO0BLyn8ZbsfuyAxzLd77kYrPAd79nDCU2tyJBHM8swL7
FECp4d6+uHULzdcLwr41omZl3rSP+Lxf+rGLDKzX9xv7H509oe8dWlTDAglfqfVB
1b4E8vLOdjQV3nxRc6svOrnhSitjHLPxqpXCwsR+yJc7s0N1K3UrYHXkcy2gHNUw
kc1ga1LT1tG/iBgGZWqa3K+pbkzcItOkOm7sdRUXZ5xhDBtQpRwHLABf1/ij27cK
kB2GH4/4Fu3o1rkypSk5ZvQ1a4/DlRE0yKUh4miXNmwcv5jJYnYw0tC6Yz95d39b
TyF1wTXvat6cyrqrpzewWQ/TCoec0YwM9w+r42w6r4zItYGKnosWxfjCBF6cec/9
A3ET7J3nmMtZyii/5C1y0/QE7kGj1RZuVVubz/vcTePgp4LJ62mBZdc4iqwRr7GG
3T8GPzbFIkMFpMqZMuMMDXiVqIzpvmkFoRE7fWOYBjdsb35aDeUNsI3hq54NPvA3
PtIQ4lgcWfCXbYFb5AowXaSFgtNlLrlCQg1DR7/wqBeYbo/Y/Do8cjtkkvUc+gGd
nOLemelg8w8cmoPLj/tP8MQLuilQb+pu0mRqhfFVF2jTUqTYrA/VlDYGpc8SzEF+
izJNFXJASwBv72Lsg4/Nx7z5U3ClOJfgpaqnaPt+jJIQVdHGUenT+DBtGLHGAs3N
V8LDSFeOO3UdLq27p88m8PxWay7zYtdrRD2TrUrs3JztkNlXwNyY44x+v2M+13/z
nS30/btmgKCpNXEIIwV+c3qQ7TCGfqOFh1bT99W+KpAkrIEqqil7xU+l3XpHl4E1
IOaN5sZWLC+6CEKmMkH/C3fZR6FdENIwF+63Gmol9/gDRGEmtONb73Fl7Bp6orjo
y9A8Ce8exHHkE9Eloc0b/p/4fmZ7dtq8FMvkA2CtkGdo+4NRkZHU1HDGvKUPUYzj
k0jJwqCv9Y49GKd/DOVVULu5VG0R1OcRTzXG90J+kI9tgHZI+Oh+dpQ5Ym1bQzXB
UhZ3C9gcWPHfVc+AoYrHa9M4gEMADnlKkvD6yGv0Zm6dnx+0WJvmDP2i2EmoagvK
EmvzdURtmpdS7QSmTJCSNIR99/S70Zaq2zoHB4FffaZaPpFNpKFroW4ayS974cFL
83lTJlxKafNnUK4omoNa+cTzGIiOhlaafLHSqQk5bAO4IL9W56lgJ5yWlo7Wg9fS
AITeblTaQkP5nY2d75Ghtzw1qY67/SE+rNGfDaJHSrd6rQ8nxlmGLJCurHCaP8SK
0WwnjWNLFj7NqrBA8cfisWOAOkNES4t1JGAMubeVQUML7kYwvlcxuNiv1eZRQdPJ
rJTzAEp7H816lfDzZQ1xGDlNLWMM7MEQU++iBlT1U9CzOLzVciPRiljuyQ1xgmeA
YYoOqmHaoo09MnWDr/11C3ZOTLuULbMSRWG7jZ3/US/RTISk7iLuBGOluJb5tSOG
jg8Tfs0p+osK/bDPj5pMGNDU/s5y+3gaRFVSZ9pNIPsrDwPLBpaYnpe0bMjplkVg
x0xdQGx8rsG3XZDSuWDyM5fCWVy6OhQ0GgkgS9WV54ArtW5bXLzRUtLEki8kirzr
hLktPpQordMQZAV4wLc+MzFOIpOX/fhLza2v8/WTtdp5AUox4nWuAUWH9F1tyKF2
fAoWEmbkoT68IFK+WQX0LQygAQnleJQzLB2yLTmxnaWikTfYaL6loXU+MbzHGaN+
P2Bkja3bw5ygEVdAr+ikPA+v0uBkcOLLR8JQzMzR7wIkzXYbbESI9UDnFbAXiJRL
DwCq3dGnclTUkiVnIHvglJIL9EmNGRZH2/sWdURRbAqxHl6mkzxyurKZJMluYrLT
+uBeYrcOfkGp6AXXIjqBI0TGcdUt9K4lCbFEhF5+F7wlLPazLtfT/GAwzGUHu4Ez
jq/aS/ncJXQQVl6I+Cv8Myjaz2QtAnkHtudQcjYmu8tnMF96e/YVKj0iL3yHZe7q
IxCnIFPMZNGiCUvXA1ap0LtznPSAyLqzL1SZTDDJUKkpGmlMfFMClFZHk7jLyDY/
L7lTJKkXGbNecicwqtgXfO6TLha9TGSsyQdxGldeq5G/6nn2DQY1JolgYlBaXDiQ
cqQxbCCKJrUnqm1R0HJVdjJeQAvmhAv+tV0a1IVJxZK+TZ3O9H9BNxkyN7IpnZWz
Zw3hCqBqkPM8667ficdoVhqhm/wXCeSELObm9z4h1xBbROfGvLwgvc4QyK4TrXpr
Fq1KoZhpx3EWO7WEG8l7ZUyyvG/sh0nwEkS4FobMUkDhAv3vPII0cWp75ho4GYCo
yqtLBmf0g1gy68Srqm4amHfNsu5g1qkCujMiff6NUUCL4dO09kr12r5tAMsdSEVp
0a3SKUb4kibxATS62tQ0+fkOmJ5d/0Kv1ljMWsy/vDWeNALXZqc/0VwJWAFz+0CG
BGzbhKqRH5S0f2+4JymywY8o2hf1OlcZUYv6rPP068yRT2QEnfXyQqbsGC2xUxAc
tm4h3z8NrfmWJ8OKu+FafplxDnE8Iz4j+bti3bJBv7MgA8BFTU5WyEZXnEtZvn9Z
zQ7SFlA7QtwVLuX/gSadjc9halvmI2wXYVv+Mo6goujoxlXJbHpsVi0ZU3iPtLOm
PCRepaYsoDdYJHUhxXr8V7zdWDcWfvMldFgM2NhM5yBRlWGiayiaMg1bfBzVhAhD
1sk3zqVPpKi+yJvtvgKryUrcUMU+JvkDCx38whSJRS55UpeDQvVl2PYZKj+BFQ4K
6cEpGhSsVtaewDBfuOuRufImHiHeJrl9d3EGxz7d3EsTA86/C0a34b2qdzWmMZWN
ElSXzHpS1A4zeIKppbVedWu4wKmN2NGXhWsqUaJaXHFn0MllLvYlfGgUIwV8pyC6
4OyyVAAi+IWoyi2d0Oa1UaPyaN6xNRqEnsC+V0ozY3ohX4Y+qtv1nZ3bxgwv+c22
fKCJ2m8A4YCwdMEUnplo7z1cxULYtkcIUvvhkIouvxHpngpOs/ZMQNtfnhWN7FN+
ubGCr8OUODLKvcXH7TZAt17/4LmU0v0/7Lp9ZK6uhNg16ASmig97AJuJvQ44HoC8
V+GiTj+/ePJvGOVjFOK93P6auEJt2WQ82z9NO7QnuL3nmqXAMf2LWd4UT6xt1BJY
Z1bLq237mnADQWU0qC1cRPEZ5RQcmV22IaWVg1kp0qN4Cmff58agN6gkoW9tdkNg
1VVUVjD4L9bCirOJF5I6giZan4NzaqZZvy+MP8/C5bHkAcil6EBF77oF2g3lvAIW
Ggx0ywc0zIyiZPVovzboRNE1uV3OTDap3NlX2fqXFpayVIqemuySTK1Yww8/MnML
MyF0jhFJQ8L5SwYZtbg+JCKXYPBJ0CIwohACf4M31O0MB6IeWauKj7ek5pTkwW1/
1IwEvdzVPOqxinP1xi3YVxxZSaVMuwwvypF8cWmI6VbOJ+5D3OdTqiqegaSDLuoJ
P2lhaosHmOtu55tBzV6Bo16Bnloo5Ba3I11wD+d9bDVVOSrx3TVdhB3DafQjqjwe
wUbYrNjrhFfSHTFfeieIRdnehpG2slb2PuWkgvxhsX7BKo1yZP8KK2pHhhHn4pIS
N1KH3ADX8w/LhjgfvfiYFL7kES4mtOMO1Z2fMg9PahNW8Sj35IpJuzyB+atggStT
gsJNJLXxrI1GhO+Ny3NT6qUgOog994fV+5J4FtwJa5yeDQnsrkQM42cJwqZgkXSw
aRupik2UwYkGSeLEex0pOWZqBe7dj59tfGPUsDq0ltsHqgCiUsJKloE3K+9JNtaj
9PEQrTY8H5nOZL4S6jhXR8YBeLMFoy6YsJANjutJaAV0wHw/qEz7UEGVje/iaUtN
caW7rF3apP+OglHRgTcoVRier+k2Me59AcYaFS5HAA4Pu8tLWj9xJFlJq/YwRuTw
jXWJBFS+/z/XDHJaf5dFUgp6KF6ZRXGhKLgz3D4Rt04iF60oY7MZ+QjceC8G3Q0T
gGY9H0gBS1EDy07iTK/v1zu9a3IWplHp7FGEfO0gq+zPLTyNVRVL0EUVyKHkajww
M1bimB4K7g3peJY1/eY5UF9U/0WrQiYlC0kxvq8e+8QVs7tS7oy1c91MnyZdYg7R
cXRTP9hQ9lSOG4iIAGSSdhJmAyI5fsA340suHzRWuMQDjofscfLD1CDSOkS6YuXk
WP/Ik+YjhsKrvXjH5/7qJLevmERWhpBHefgNQyfB/wR7OOUcaXyXH7rSbaV1ygwo
bNz5GA+4rDYENCzBEaJQsTZxLVtna0Ase0w7zqDgzaGlBxn1VXTPW0JVaqS2nbs2
GS6rELTMx3eqpRBbLw+22lU3e0WdiCmLGbAJX3MZJiv4y9I2RzcCeEivinLgoqch
1IA+pWjCOIyttwnIc2pmdzptmCZdZZqY+tBY0w9x9s8tqbi9xF/1cwseNOVkzRbN
n3+jJiK28QhqgfSWX5HiV6UJXba2nJLf8C74IDZGigG+gLUTveDQ0mhOdA007X5Q
TrammPcue0bNWAqaA70topMNUpsEQwg+tURrsDx50qBRcJnbUy1LT42/PKyfnJYV
NubAfoJ97rswU1WWc7ORomP/23CH2HvzCWT+OyaEjF00BZigBP6cif3pnexUg60H
M8awrLo1n/SCFIJFVQtpM+T9cE1jYihmAasz7diukdb95SClQ5DTzNidX94vx2DP
g22G9IG8gwgofPmROuI4UuV1eoH0W6mx13/M3BJmYaNuJKnGkWAgc+b8vAgOdEyS
CziReHPgf12K2DSSsYKm4pBe3YuKM3Vw5wsVNmMbiZvJtmg2jjPVA2xjcSiDz4vC
viR9Nsjv9nynMitg891bMdKNFk6XDh4j3jgHD6IKDF6JciSmSKsRJhMKkUntVqwE
d2qt8Ik37kUeBzuTEmyu/0zDfthj5MJBZktC+tP62d4kCj/nzeNAa5qRqA+7p5Lr
W7GMyqBEM04tmJ12Kid1ZIkeRG3yYgfuC8imdyrQC2PWqY2HqPS6oEOzpWtbAj5I
S0J00xZgReaYWNoAkpAzpQ9QK1syz26LL2KqmGNs0znBg1GS6/iHZj1eCOBFeCqo
ikiELV6FvTjISuI0zmozFQ225hADLzoeODGNh5+Yabcat2CaS3M4+AFVbxdz8IKu
qHiJEQmtW0MqF2XWwgOVeFLM+lhT2smzGD66J04IP4jNqMGKLDBc5CtB7HBDoOiO
1SQhjlya/cm6Ek7YCAPphEYsHl/X6SF87nYElP3vhQxqFvJj0ZxZPJKeEc7Zexum
UJJFqq3CxBVsnbLzi/LlNxZlygRkk8e3PaB2XHdG1Rwg67s/H3n+UTIg0mt18V2j
zXFIZO/e2hGfGufx07kmD8T0Lfegj88KwVTjUdzWRf1OBN+DEmkTJiDkUsO+wyCo
XZrtrwn0apfgyMSeVDsGLuuN6c+8+mCp2HrOr1CCBhPJUEriFRZK/lyt5ZLmE2XD
/c6mun3BHjHZkTWatGAUgxhsP2vWH7TY3rP3NIYEeU2Pxfz1y+UpRi6UrM3Ru4t7
r4eRxO11rT/K47ufTXtjm07Vn5OHEQreqTCd8yEa/gnufKYXwL1Nr7gZSfNJ13Rr
qffLNaPJXZdPjgRYazOFN1FksqW/JlYAgMoumOwaeRE8tr212yoGu4dnd5Voi7U5
R+kntrOEndhPFFluEUHBSPuPOHoK1aICKa6nSsZzne9JWqLP5ddZk+qAfDLtD8zi
6i1yoHUZE5irUUrBCzOKJ5Pg5ZJ1zqZZDRifEuMzj4sv/PWOh5jCWc2oAVKOuWl+
bUCpYjXNhY+lznOmtEe7Ac07gejG9FgqQtVFnHcf63nthJ+Gji6UlQOebg5hALOY
nlapmOo5WXQofcr4WhbP2379DHB83m+HlET7nOBBEyK0zC9nyNb2kXxbPnUnHWDD
YmwPCh3mHU4XACPeal9fVm4lrt9UsDpyxkzGD10u0SakU0Zs3fKWkYvhEzS6ATFM
RMGG472AuMeJf1UA23exLwfzxCAYg4ouWQlWq5KvMJbPekv16v/ZD3f/0eVIbnwg
fcf5mmXNsL5w0pGd/ozAlMtXYkJeVvisWgPJQ0RVJO5SCvyLoDA8txV2ImWtM6zO
u/hYgQpGpcAGYq0wwEfuUZy0z7R7z/3RPVqC1nIr+23btYB7jVx3StQx0IvT6fOu
2wZTAWhJS2b+Ef5EwQbKsI1SYkwk61Lq2zEl3xPr9Df45XU17aWDr+QStaHW5sXN
4IWWCnMnDMkfvCrgonDuXKV8LUTr4gaFmJ2AnWLDzXQ3uzcmOpmD1XfkmXN/nDRl
MfGFArUNWjxzQqTq1S99WIUnlAPCYerus5xXZe5n2WGXUv6I9NY29Sdu7xi4xnzv
Gtrd4J3VaJpyciyWBrbN6uZdVUCNSgPSeQx0cPEA83RaO9kUSHgBzIbPPnL8YdTs
MQgN8q0EecH7HDOL9v+uAaOnUCkssDihvOWXkW5wVPZSybyihH3glRvXLCTnZeZZ
aZSRw5BLENtO0pbvD1How4L5jc2lmrgYard/00lo09BqnAUlKijHDnctB1Q5b/Mh
/98P4adDKayITSWnR+eu/ufHcGap6d6CmNJE2QjNdSWGk4MtebvRRJy7XZRZm0ep
ikjuW8f63V4JySXMQJZt8uK5ps413ES3no/y3svZdHLIeTk+7Z/nU5L3aTOAa2Uf
TxeRCJwyc8wbW1/0yM7mir+200NLtROpOZov0u0aZXnICx4ckQBK0iU4Z/AJfCky
I577P9jAmMlZa7M3aTXj3eN6l0y0/uiCxPX7Xz1603xVcgFhRFAFnuT9RAJkvI2S
/6OTZ3rhJ5CYpxxd0WfaDedo31pyNJ494Jh4ewZQ2n2SJgnnoEqWtOiMs/wJhjMe
Kvymplu76EEh4opVCY1QzCuIip3PDJxpJjQxAr7E5zR5fLREHv/tq4D/9IGtFvRn
Cbbs3XGtioaqumQ57F93XAfSVndzDcSHZPyChFp0yVBRnazlWTtQtNtwI1kq9J+I
wUAUXDsFotgfKzJ6+lMogkY7lbbtVH/LwRU5zpOufj1z00wSn5szj9gzpApVSoVw
G2pnHx07bD8i6KnS9/e/xNYvLbDRCamwn6QvaMluFVq5TMFtZMIl3J6dueNl7wES
VTrHlmAC2GFzQZywgi103OFSGV0RBrPdWNCuD3nFIjWkUw9AeiFcrC/Dfl27ndKx
pID4KzIcnpv/D3f5KA+Dffa9pcvOqapAH8vk66w/Ek3EksVtsjTSpUf1VURy0GbV
yke3j+A4RTKVpIuhZNPVeK8FoPBzu2nBsbF/TnH9yZzHohpwTdGre0CapLAe38Jj
1mgqFGgWadXwOU3PurrOZPq3k+frXDv9GefOg4S7LWUcmwUGSjGg2wx7Fdv+o1Ld
fvwTtrp49al6VcVsJEu/CuvrJJXEJlhJ6gYyxHHQiLVVPuXyJhvn9Y1KvbPgwAh7
cLa4YhiyeZRzYgKiUSH5eCaVZAgDCbnf/RAiGlD3wfCWIsgOC9Et+cAkeukoPnSc
A/Ps2EkG4h4bkgo2pYeT+x8erP6BYajZT94YgbdQ9qTWJcV4/kr5/ma5xysC5Mt/
bUnWo0p5CqX+kGoSGi4+XBd8tfbOQuzN+t5y2LWkfH2C2hhdwQnMhWyami9MMjIB
aLQKBY8M0RuIkZiyPZ0UQ5pUVMNlyx2xBwXYi5MbBs4s7NSaT7ou5KWBQhCysTRR
qZfCqZrWEW2KYUj/cDH6NSr8otkyXOB5UKA42G/srgecpRB+rVRBVmvn30aOuZLv
4YTm1FT34djjzvT9sCbQPOv1k/VffpRwT8YtLTMxKXXgT+DrGcrRBmd3uJAeTjDn
TONJmkThttVUYt3BnUKvd3uh94R5SdqU0e42ASJGi/0WnaKrnxTxZvpBpy2wknlM
7TjcyFE01QCtNbm3nJOO87w+1t97qs1QqkeHwt2LCRlo55w9KD6otk4LxxUgpxo1
xXSakmXySVfSMqBh7Fpxmg7zcGKNYNhyYFSsrKannnYSph+n5odap9HNKrobFjbz
Ekegmmk2BqBe5VNa9uFoJ5d1s5K+0Cf2Rs4uqgzcdvdtdGDNswMIK0UYmn0FbPsV
mFGpRTHem4gzDz7XAPoVkz/GQGVjWUlZB7msbD48WgE7hmesknJmpDC/qL3KGPfj
bVipBjx7jIQvElnA6mwYBfsl8BC3ptj/3S6Q0oIBvBaZ4TgE/GmjnwBIl2nGsCTv
OlAzPFNSYMsr/8cCkALKsppMdercziSBOxQ0JmJxUJaiWdS/P5H8ttjSAogdwYfq
F5k8naq43egLcyJO0HFgFGyOOAGWhTI2OynaL3gvBavigksfGtOJbfXxPbTlLJfz
H72xXyc8Wkf5cE2eGLU+wu3Kt19fVN3t9Vu4l0obCTVsYFX+oddlQGWdD9hb07pv
fVCYcBEcyYGeet0/RADiEzQE5NA0ZepGp7iiSNQZ5/2yTUuDwM18Zzpq+12ntJwx
P5D/VCULx6GVW49IuNDJZkDFGTuB8G/Avs9Xr6jzIXHETtdMrJct1crbNNOh4yoN
n/uQGEqfod6RcAu2JKzQtFP2jxO45p83GZ43IjGKA0hbCNck3IBe3DDFjBSUEcjF
vgsXpCwxnRFbZXEmHAMWTR3VX2FneAnWJalLEthPz+UFl/WFJpsWHTt0AEMXoYFR
XK4z8z0luIv2kM6hwgqKY/PbERXpOzPJPF+ENvLp/G0WvJOezZZq1LV1nuGD5rIB
gMMK9XlFfvqGW8XuC6I+XSIBN6ggpEQo2XHKNZeqq/PSM1aKsnVEiqkJD1k71k8f
mQEinfrwVYwwyX8gDZGQezSB5MWwzA1pWzyXOQeSTtoQRtTxWFu7MNCYCNT5mFmP
8fi6tv2nvQh7hfTH8UquRm4qvogPnb6hzZSyFzXN/MZCdG+2RfjNszLblFPBDWt0
fcgTzR6sVCU0qfpiZs/ZiR0y1uyFtK3eSkiXGNT4C2i9CQ4nEjCdl+nBYyhpwI0W
NgEZGzN9og6xAhb0zcfuhjbZajL4tpoda/2ojTmCtnFEqem8Iy8K7rMrMchZBMl1
JRzTfA+Gkc3rC3iuFY9x14pYqU/g2lS5DgO0haF8lmDqNCfLeTuV+Pb9KP1EzAf3
RUZ1CKeWJInk2FSN0wpezSY3lf3/F5JTWU2p9zwGSdPTY+3xbNMLC7mSQU9Xn1a1
7NvaHPjapAbjUlfEuZgRMVZDbT1di6+NyvU7K3i+adFCqdB4mvwRLk89D1Ok2ZEr
sU73wGknGXvRZW/lGXoSAGCZnAJqJeVYaLpP7rNQQBBmv9XiJATtW3MNlEjnzgT5
QgIbTskflue45I9f3YBe3ZKlWwZ64+/WVCMyL16CVjdREiXUoSJd5hOTasTUohyo
d0bjbpy0EgAVm17iMIFIJEMnVvWGScobZC94umrHiG0o52eC8inkJvCLlmpGc2VL
/qU+CLdqCiNqPZ+zHisfEF+U3UDcyI/k1f0ZHSpDH6mQJZuPZdvjRm2lumeVD9Qd
EFd32Q1UKuVRHjwlYZSgjfXLcBCe7yqdM5yiHgDxtnKvYODE+SVfZ333RrEn59Lo
7CBIextHfLw9wR4Smodav5WIAOGk2ftyH6ITPKzhVEwL6TMPiC14B8k4juwmASn7
oghtwuWEBiuGD8Z2Ou4IFZ45eDG3Kvom9ZNnhgWDn8DgbzHP1D2mR8mIkblq5K5n
V3jPV6qSO7G8iA528qHRg9FtQMsEpVsXWmr5JVk/RCfWx/dZnT6n3BW2xTiHM8db
jl4sUgitOsiiMTpDt9pWI5HrIhUDafEJ0g/RBS/SatecI00ID4quWc+JomQx+8P3
CugeotpOCndaw1Xt9wGI2MGCitf/bhP+1m1EhJy/dZCL7opv0tPtd3HXc4Syrsr6
T1E66EyPhUfGUyuJiP1QEOso+Aih+fg/gUjYxMgPex+4uuJ/Wjaouo4gXAzeiz3x
N4lwNWFB/x4gXVkYZFEdxJDGkUyJCK032HEp4XHXMYGBz2bS4Q0GZb5O7RX/k4EW
1Wxfg5pxKE72e+Xr7w4PD4rZ2+SZKLvUyHomP5/u2qA+NqLRaXbZe7LMxpJI0YHu
m/hffCKbFoYnBO3K/CdsazY4MMlID2GTw6Vey+Hg5TmqtaN6bNw0I0Ko/0DsPDAj
9ez7UEVQHrHy0C4YZp+Swqy2TiUKctJ9rCleKz010vsnsFG2nYEaerdCnyJb3zl5
8lAD4fW2nEjv41rqDcE28UUds1OlN9rhWU4K+tFavoRplrRKG8k2wSM9YccJodMB
Yv0UAipyt2g36FJEMm6BsmCmaaTLjYTkrWV6dqgSGlGp9/zBrwHFJuiIeVeq84QB
eaTGLA8sPCObhNpBQcYNNPcUexTzOHGIK+QVVAMPN5dFnNym4iPtLqLfGlVzmbwU
Ln5VLZRTpzy9RsCyh1X2J1sUWrg6xyJ1nNk8zpQPorZVinHVyO5jNdO8ibp3YZq+
QuuLJQtvSXcZMJJJP/1JPVUp7aq/akzy9CUikSQLc3NqTemo71IjIMRrRCzIArop
FKHInTg2dCHHFJyfesUYSS9mtwFJ4b6bnFy2XGBWhjNsDZGgg60DcHC/KsHXfjUN
Kox2Wj0Umz8707C9RpvspNSFIcmcZyFnnf9p4UKK9Jo30s+uTjD7KSJhixhNRumV
uQTAnAyd6eGV883sIIl6YIk5BUQpsI16Nq4SYrYSfcW1dCF8VIQKQVKDemVAn124
LR5vspf5pRMx3aiuYJTIFeq59/ZfYqhWYIadUtqDyw+qSGR7ZMwKtrmDhr9lQips
OM9TVqZjq91saaAQVtf+HSSYwaLdz8t3QK/WE/euj0/tY6d3yNHn9yqUGgchDCVZ
pKxKkP/jFrEfLniU0ASbOR6OnzEAz/ERylmpY3uVsNYdY8EV9mcHtXf+3rbNpYrh
Us9/elE6/zhmT7fvBUOkB0JLcfD5cljnA2muEegfHJqXgkxjPTijl2Xy0t0kYff4
/ULL4auEjCJXpZpmnxTjk6ZMrY2fI6Q82CxP3Gjzz9nhrQ54MT2nGq2gHzY++vhx
4KX2U4s7/Ny/kSddISqvsLUdGVwXA8iHcRgRy+ie05lIV+R43cFDTpoUOihMxedr
mH5zC51trBlz/I79rmqIiDpWgi1Akf9zv/UECFvBA2SebfMOLNmlKT5dhfrbuxn1
f40GJ4RnJXWaG94JOp2VKhrweQ396YyevZysUFbUWOUNTnu9wUNNIwTW84bES5sH
0ruN1nRpWcET2ZiUcFS8WTL2Fx9T0Oj2kBv85MyPmkVw6BVj7mSZFFJ4jU2rDWBD
rESX+NqheEzBPB+3bw4ct7zTCPQvBocu0ffVxTq+8q7tkjfxMKFjqiFXQs0gyDHo
G7RZOVIf+22SBsb8KmJKnGYbxCh12hOkZxw4Pos9AIJ17vC8cUKxoG1AKs3TezTg
IBgcOU29R0onnj/3y7TSv27iH50goB8IY/DMaQP4famKyKbGhEYQ4whIKiBRgSMA
so7QYGu5forQQNxSYt88MTJRkFYL3kffBxmVdN2yUejwxB4iLNTwGTC2v2NeAy4F
V3PosGDObuXkGL8G+UTAWGQ/JYK9a588uE53ci5PVaRXSTmfXilERjsOOP1p/Sei
d5Z1M+1PyqBt4ADtr+QwD+N6vwTQ3HjTt9cBB1V41/w7/53h1YPLn3YsIx5bzH4/
9jMEria0+8/tu94kpdTlLvR7O66WE6KFbBtIxxTi8W281IiycffriOt3ir2++F/0
Za5DbJlwQIUZHThWs91oLSJ1hg2Q2Qw6pR/61p7EiGpUBewFFJ+OAZlXvB6EnK/p
8jimqjh4pSs1UgL4+VraDE0aul6K2okFA/FP7AmSm+J3YNZxeQazcgnrhWZi2xUR
1zD5pXLTnV3zbiyvNwur0iyk/u64cZ1X1CyOcXa+uPAhcgF6PDySWxgxP8ELGl+w
YztlYhVAGqiLy2mK2RfnxEcdHW6mlCSS6wB5GDYTp83WN5LdzWYGONzYd7TgffzE
2I2egGx6cOJVh5LpDL8wV3vdFCJz7OvjiFOtcRPge4zOi3GZLJI2o/TmjOKt2AG8
MYHUeN6ew1duo71DPRTG77vKX/kdhcMI4bFZCPFRrItzcShob2dD3p0UFN0+qD5l
rnWR3dlOEnzY45PeUl88SuReSc48s+eaMyLIZwX5WTrzP7HZEJoH5KbaaDyIXSri
/n6YUqnaIeBujLJp9il/hKLv2X0Cgse9mUgqF1BIuGP57fPS9VtZtMAwNfxed1Ji
NKHd6sHhiFWKqF5v3hWWpQ5pI60UNPUYLT2Oe2oidF2jMAWQDzDJQD/y3lrqQOo+
ajsj8/iicrY5GrdzvNdWcaRyhRfZmH4cClUOZXcXZaq5mmwZ8ZL5c8H2X1Nu0pBs
Yea3b6LFdmL1vikhrUFKNSXRrB/q/g80BjAWaLDWJWXRU4DW8+amp+MI2Rv7xaEb
ZY3SUvCAeMe9cli9SuhCSn8qj2exiHm5f7cQQX3JlTeEW/s31unvih5UWPcUnpsE
D3aGRrtw809Er8nf5thRAU2jUuTL20HafQ4nYquZ8heEJBjNdamsi5YWNLYC92Pe
5EN3xhFZb4fN2c9fwz7ZcQSOvnwwLR/N0jTdLk0OGuX9ItDgCLPnJ7lDFYcVvMSY
7w3+Ocv6TkaxkRGJXOtfYlBLSUNL11cfDGv+jHqZ7WyoLaYwdT3hSndzwLKIVWa8
fq92c26B+NM3Glao+LSNPDjWbd+e+JqVz6JyOjpiaPex6gBX+D3PgJUtMuaRfKfB
QqdO839borah7G/NchHWyo4R7FgZVZoGuUTTvUCJae1yeeyDB5FIwTp6nahkHEP6
mdGFlIw+hKV0LeH5cgJUiiPzxIwIxnwqKMrb5qjuMvvXNfb+DsIItcDwpuB3+pLd
Tzy59c3ZQZq4PzYe8dh0b0zz7knPdboFhRrJxiSPv/YCaupR5/JEKH0firaTiuch
hzfizuaJfBwbFQenJZMkL0vHOMXlBvzmwc2jgmEfvOGBrgM2BLnSyMc8YAfX00Ca
6u6E93om3WadoXj6tou3w5HO4Z1gF5tHotv7E5rBlAITTq8raQE6mJUYorRjuVBk
ibPdO01nD2XStrFcVIT8l6kP7juLjJbeQpypEVIsK9Z6FJWp/1oXuevuSc+ONhYY
1en0oaMgrxvRywHGf+cdZdupCAfEI/PSpP0vF3jNLTWpA4U5ODIy55OMEDChQDKz
FymznRnTHe0yIiAMhOxEhp34/M91xn1pwJBTFgoSl4u4PDnW6ZN4sSQ2J9vADPBq
78CChG/Pn1AK0Xb9HvO9agg64KfuhHLcp7ayD/mfHVftJpjNaw+JohHwA01YoK8j
nFN+6bn6LUhCY50IBt2O5KuvrOD0d+mslZNfDoajz3Pttx9+KVWeCNzbsrUE5DIT
ayhdmPSiUFe7Lt94NNV0tb4vsrWx3L/JMKrDeQOvWWTBQQLAMcljRoAaXnoFDj+/
huszsEtKS2rBEj82frz6YVheXhjTrcvKZ/thEL+TgLfD+8tpAUZH99adABU9NxQF
rZS5AzaJ7Rx7SRKZPCq2Wg5qzdyd3EXM1bTWiQOV5BdHTLHE5AhBciW4pwPvv6pe
VzIw+WXaFDEHRjpYyVOo714kUrk5k35A2bEaodNmFxROqJK1vsaBND3BibA9iJ22
ZBFx7HB1azuPnfRZC6suA7RISorxHyUwbnG5rxueBUq0SX8APkEehSsPvzsNrqFn
WJY1OzvEK8gwh48Jcu2cYnrbXKQXgAnjoKDG+yicIZOPdkGguJT1yvYIW6F2KZPy
+bx32t3P350ITqno9QAvmHcVkgLWWGqZChTq16y7SS5wMREkoKpXjHMJFY4YsRoT
vJXNSVmZRBKBhjauayvZ5cpHZsg6CNBtcbvcgmNnLuI5v2jZsTWmx59KUnvu3AoR
RjNvaZwj9JgwP6wKReYsBxpVvQOkBSr0FNpJbJOg8E7LiKH+pfC94mWFNxm2mTAd
6+Ah0Dx9E6EYLX/gM99waSICeiyb0Se1yv+Oz/BQCE/+b9j4f5P5sNBo0LFV/E+k
ZjKJt6y651amRzVr+bPu7vi6IRzEiEd2YbwlEpXYQ54JqSDCkof0ng0onaF+0v1G
1eTyO29DRmwhU/T4zzIF2kDj678EEuGPY9ZugBBrGu7vgjy6RkDGjn5WxyaF5KiK
hUrTQwKffv++PkPz8k7lxgK2/UOpoemzcVcYFFB36GsI2YEHvCNIvCFyzYbUCfO7
IyZ4CEu0Hm0Y4cf1htoNtHq3Vq5UfmXtet+k6/mn1zZ6SXm+AoMly6RnktNYD/kZ
OE3NO4oe0U2k+dJMtATK1fjd7rbMzCvhVwJE1C4uJx9XPHJXq4tQZrY4m6bz/Otu
HNB2+UHMVzPkB8NCXkGYoc396h+7vv4BkIOX0GWCZEepN60YbIs4m4PCu2AaQ1Rn
4P754Xr0pr42ch4++xnYN/KCaiMJIY6LizH4jq3c4NTTRnOc7q8k4NnnjuHLG3ea
FszUr+r9v6ZORLXqlKGsS3rvqXxRuPXdp721HCjUSLFDzPQy6NHGd1x8R43Q5CJe
+emVXMu2Dk/37XJJS5O8MhDL6p0rAVwnFqfIz55a7r2le2SVTXfteSqVrmpCznkK
V/d3kk4h1XJq2VA/Xvax52K9JkzNpV2I8L1ruZUVv9kDmI95g/wqSS4lKpA0OYII
hZhuMbwKh8jl3/Cc6zy0XsGdcS3necF/rSbzr+d7Ox/QqM7EwfOIEnHrBvJn5M94
4OCkphBILEib+UR/NsI73e9gWyToyhgwq11M57EhwNVAAVFLpf5JUWkJXUO55Mxv
LZPCnBKsMDyOu5LFXUtsju5NvNWg3wXdd987oAryFcM4axGXeibuMjEetSKGvX6Q
mgK3JjOoSeVkEyJiWtx7Ayd2OTzBD6V4mFf6FNK31mm39C72rJ6skia5I6F3diLt
TVhD3sXqCtHR119UTziu04/CSmEvuVKxmgIlpx/b0ke8ri/H5bRbDLQmRZTR4Vb9
wAMvH3zf5PY6WAglYq4K7wzYfaE/6rCTGV+csmRBjEytKyQlCnj6Xh7SuEFc0qRV
BDmbBOpcVtid5vQ5tlIaGHYgpBYl9nI1WgoAfAbqRwR7xEHvd2fQS+c4nb9Q7Gkt
vDlfkWFoz8nAYjvIn3tdOT4/2g75wfqcLOxqS7UxPP0Jk8mghkl+Yc144zjs8Sds
ObTi4/aMoPdFSbgEiWYVRsOc/SFl9mEqfGTEx45fGeuKTm4W4EBe6qBHzB4vTI/R
KVHfQXg6/1QReSpGylOLJohYDbgim32tR4f4TDQalhINnq3UNFTTZsPULm+niUhv
QfSzZ7pXQGNh1AyDoFH/FAEOoL0mGAJ+1i5Hz7ZAxGA8eaEv6LFNod1P4H03Zmnc
zjT5D/niP4bgQ2+bmIoSoGrIPnmlzCcQWhgecd4iFaBD4mSUIaf+goYM3xblLNCE
aCStCZgr1Z0L2FW57MJgNjnRafI3Zm0ylzsGe1MojnCriLYcB2LnGwNk5BvfrVdX
j+Pyf08xcYAAIbPd60pnLQ5/cUr9cEbTnUe3YzGL7FsKFV8wsB2Rdw1/JBP89Sqa
jp1CpzCF8S/x+m2yjNJOrD/CJEydSVv77ihRiiaww3DIh0j/f9DJLVe5AWYnNn15
lhh60AAcel4q9wiyRjJHRqsjDAMSnovuQJZLzYmY3eXC3eJZImq9YWrWp9oz/WUF
jSK7faixI8FC+WrogM27QpvqG2gH2avGrRKJc+iCcKUnJQHlcYZ00wycxovPF/uE
+GGHP4AMxgxYYbt2QlBVilYlU5FVi/UViPGGsz2bzYntf7d+hQbh69sHrC2Nigt1
TdKFNsGiZm4Y8T0eC9SJZre40M/9DiLWlU5zZTeU9gHmP/SzmU4Bu5K3wbPXJp/L
oo5vyCnR/xesKKVhjqVOdcrcfdQpnKpMturHDQTJ0szi4uDfcaZ6a/umuC67UrrS
ikzcr64LwrGsI2jYfenT4kBr9G7bwwqEwJF1XnqlR30p+9hJKkEj/ta84Le0LApv
aacSIHRLyX5iDVFbjaopC8GAKpjTX/wF5JhjybXYXzT8bcA4pZZkYTWhSmM9Amd3
p/KigE0/767op8JPr5T5nYsDweKrefc4qWFet8XATB7+xincvJggHC0yAD0nBhDs
FGVQJOg6qUYzuHXEqmklaskQp3vXjosMtQt9DfD8pY6laYfteonU4c5U+7jLkJFl
tzTUP2cWknjV8arHYNrwLv005CGNNDBKvsXlozmaWohBHqb3txIWsfRwHwqaqxtW
+98Rb/OS3aCN0DNNFw4ERfFpAH6aZG79qjsMms343kd3J3HNZZybajHxl1AcnnnO
O+132KvClcVEPrfn5N5KP03jJQchP/yXAFCXWJUB+MCkSDdt8c/PWUF5beti/wHs
VJ0WtolxDJszjqkSwQ9Uv6rHPB6T1uR1FWUVfSzbbvW01wK1qeuBYZpjhKrwqkUE
VV1m9lvIkZqqS/kbZOQE4gy1tODgMdj+dEa6KrFCXGxENA4kPyxK93mdZz8uL3TE
kuWhNaSl+pAg8RTSdaW1L+rubW2SioLEoUdYiqjUtreL7yfBs8Zae7b8tD3c5HPN
B12znykN2uZV3VdC4kyOOAj7Brs/Jfj0fhZ0g5nMqxAxea7sQqkqwFrKiHSUrMhs
eHwJkeD84qLTJi1mUOwdHhxoUmaaa5zktseyNT1AzISg80A9yTkrldX5HlcLAbzT
PMIliocJWyFxmsCA6s8hr2l+ruevdjsMl75yBAhWPBZSIuNoJ8/hZ8ZUtEXUODej
jRyCVQGoR5DEdMCcWCvq8HCstd2OD7exgAyNiohybkihfcNjXRnIfhhQf2tT6Fc0
V10wsPT6icEYyKK8X0lRIC0R/YGBTCcV94B7LFNpgqAnlRTPwK7HwxUqnHBL7UIb
len1TFVorWYI3ufCTRjfyaBOCRmxqS3FaEDhVCHYb3TC920LdZ8n/pbCGHn2PqFE
FGY1wZVTDpzQIbOb1ckegwCK+/B/MGnxbbf0ZvghMa+2g1MyDRDO/JoeQXG8JzsJ
xySBkPW6xofkSbWgFEJJr/p9ytLFkbWtdEPkt+VfcDflvn/259WiFu43FVZHh64g
K7uIhsxazMfQwFEAESkXMwvUtPhidfnTD7dZJedQas7YSD85iKVe5izTVmNIfBye
zZiNERRVIPhrhrffIpejWReUS12JQKSiwB1y8alc2v+eE+wuWrao8UwpneM2rzDy
OOnFCetGXyk54Digoj8KCA==
`pragma protect end_protected                    
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
iEkvoSTdMpBpgZ5AgBB7MjZqpzXUJjwRUG8zSSVbuKfnjWwYtSwelMts4RGhHUvJ
h/U0joWYnn55ShF0VKvdglgo0rCP2LfeUetlV/MJ9NQfTBM9mePNLtyqAY12AnC5
4+UKHCL1dLqaTFOl36Ww+JXMi1Auis5xH+t805cQGTE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 50248     )
GSgyS6lBX3JQJzab34ajMI8SL4XPot6+gxpquZipj6PQcgVMC4GIo5k66VB+oQtH
vZ4IHDnq3M7m0jX+C0xMyqEJ05W4wIXbVB2+GyiaP3r6WffJxt1DFcRVIAA6hHt8
mTMcl3mj8PEiaChElajqQpcbZfoBobLP8OcJaezPqpbPzHoCfOpYlalaliHr1lFq
jpBtH9C8mBZ2SDPYSi+gI3X/zDc9Ie2ZXOLuYSxQ9sKwvGc630+js0u1PBm/GQgG
KNc8YfpZrt+LzEqKQoaYsAv+FEOSxXAVI0Ewfj/fhcMiSZjMXyKjrcgtXSOaueAk
kIw/bW/Tz9iBwhnOlRCd2ZFx6NGA55STM7ioA9CC+9nPpLCyS9pRE9mIKnni+RSt
XXhfSAlUOVvxkUhcDh++SRleOFMsEy+prNjRuywHbjt4NAqQg9R/ETCFxh4fEP3N
QAdNPBL2QvKDcL+WuCXOxD6jZcuoOS9xuXfUJQIL6UcPBoCdtoPo1XZaCy9oyqAm
njOQL/7JN1APGGx0zYB4xtqu6UN0ENkcW+/dCw4n+t1JnarMWJNQqegISTf/yeuI
fEhcETvaly28+y/LWQH+3ZDHEDAmqFH4L1YTQ40MQ8QXo3BIQOh8Tp+40QHdPbXC
Pd+t9bH6xXMB9QBTOUZytw7W9mzcatYIbdmXU3OLzUxWBBgm6EAcwlzIp+DRyudk
mn7Psm6GQcEF66i763gfw2Sz4DVrfXCvH7ihLTdJbP3SAjfps0HH8flXNe2B/Udh
zKX+Bm6O3/RQpTEWIFkdBiaBbyTkCBgsMb4bDGIyMx8VLT4zFHlV2lvqEPg9yu3O
yTkSgUD95vgYAdmbjuoCcq/TytPvj72g9Hd3w+lEYWTzy1VCShZdEZa0biOJR8Np
kgpJBzwZXklPr3x7Xul13Izv0rBWpSqKwr05dhTe2MopVB1XhOnzkvy56ailW4GD
kcEWaXJPIy9j0XXY+ur/aZietP4QWNii9iYhCnfKtpfFt9irJ8tZmwAb7ESwmJ7K
TuP47Yc4AtClVs09UlPiJg2WflJ7viwon87YG9HfsrckqxfZ4VChasyoX0kGbdC/
YJKCOsUevdFPYeqc0FY/EnhAR9hxHK7RGaJxp9E1XKqlKQFOKCfnVfvzN01yFzCP
odT+KRFUcXfvqMdYkJio2ZzSXi/9wwXvnaO6SfQNY4u7nsuvBlY1b5KCeiyBNQqK
g7OFj1akbwOWROr6LD+dXMGp64QeC535e+00kQYYLe7F03U/YMxsGf5qD8qe1Xsx
KyEiCUtCiTl4LLhKpS0I2/VnKqny+JZ4tSwn5mFYRtGPJ0n+8fi/HhXl4FgEEqbI
gQ9qed4syXQur2gFvDgtxBRG8eErvl2EToEel7rzmRnNh5Sc719NDGsTuRTB3pv/
/ionD5bHIfHHE8TWNvCrNbo24jonzMrht0jBUZzCJP3SxDrk45QiVQDyxYBddDH/
nglUD00HUfcNxEWTdUbOYcitUD1evufJIYjwCFVtEVW+8lUYcwCNn1j0mtejKMCx
jAVBai7HolM09yvMNSGefrDs4N+G2YOiHA1aBObwZ60OSrc9OlvuLI2UTVMlL1UW
zOmDv+TStvNMMkjsjN6Bydh4CAWfM7sYs1l9QTZh6kMKaxYRrLHqR5NwCiqAIoPZ
cEg2YfUX+WwgLpuXyLzau+8vuTBZ6wA3f7eMCWsOusKfJQqNMjYp2pGKPFaKSGi7
oaqanTXoQMiGD13ILtSPFl54R+fuUsmRVhah4kbZG9JxEScRfIoBU6glBP6xz91i
1BY9c9EnZsow4cIgwMamrtxmDMK+YdTjzNqIUeLhpjkEkO6LXUCWoy819qT/ioar
hpq9cBDLLNH5byXPYTqi6vCq/rYOWLnit97uv4APBOcIvX9oZFVue55zPooBw2sb
3gkPFL/pSgshjAgOf1gFfitcLc47+uIencuUmI9mVh4YOr7W4D9QLaDvqsFjVdPu
nVEuZwK7O0n+HCSguC1fqmfj7W9GYKbHvqWzJe0x1IAiI9vWYwIryJHxput8Gev2
H4XOccQgV6t62tGMuRNEPOznLNy2TwqpQjm3JwtxsgZd9Cjnm5d3oTpXO0womCBJ
Kruub8GUHYvhp1NMPXkyG/pkjZb1jACFG3sKm5d7E9PoRFIXBQBXVbSyxPCCOlGG
FfyJrgiff3hXRT/sH/Dzriq1c6FGgF6cVmlniCJ9fp6KsUThDH5HyKx014vBg+Ck
7cc08JKsToSiT04xAk6v+Y6Q2U5WGQwDupxw9gMCCn19xdkPidXpxUF21RKUa79W
W4JiBcAwevSnT5K3HF+SwvzmgbKdinArcd4hhhQv7Ne+5IkA4rwa1droRs0KVfSd
n/9krZFGA9DaAtiLEtFXtlUKWQ1CUCunTpf2AZrbmj9lj91czyXPmDuym28BPQY4
OhmJWXu2hc4zqNV8RqhbJ0cjuyWQSmm29A4RZmZ7NaXLs5qa+G6ucICnaKLiFiyD
ecwcXWnusyJ7FVbK71KLIBxkEuYu0/DYn81QAld/ucRLz5CRZmEeONXx/V4DhZjF
tws31fFE/nL8qCbhdMC/Bg==
`pragma protect end_protected

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
cMzNslhWR3dNVGJQhmJRAVNpgO47Ova5BGHvvuSSZ0X7FZHX0eKPcDKyWydvP2si
paXQ642YWNXvgiWmCvspj21lRKV27rsPLuX75hnLUpihf3qnvV8a+h/EMKx+tNWw
D7tDut++122fchak6X25iWxrUtRMLf+cEFTatcrmnpE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 96624     )
KOt6Yb4n3N4+gAmZvq2XmzuGKw1Wv+3R4wd/3kXEzqwfwfV8K1M9Y7S10eAl3yiC
ZT87qx0LQjCPmOqWF3iKYAFBMqPowp3Mn7+2MNaIca/r6y0h4NJRzjthj0M0DlPq
JHsu6nW7fiIW2GJAlDUgCeV+CeFh2Iu2230+0ONBVCfe55KLYBULUQn5o76UvOGX
SRQDLdPBqGa01QZ8bDtQycjpUE2mbwdtwrHbkcLDneDuW1ciHYEM4Xv157T4z7+q
sYhZMsY3AFGtKpGni47pXynF2RXRd969mwUlPCOcJWdAtkQyvpH6X/znxqSIp9Qp
YA/opeBR9b9r31i7wOnZVhpTBSq5QPGuoJO4dvdZnlmj3cPDLCdTJj5fQ4cAsldr
f3DnP6VuMVkV8OiHY4b0FodyHnwOr92sblJEFHz4dyX5k4RvhpOpmTF5HjtIsfVZ
/ijfr7efgvTP/aELaYV9vKNvM0MBN/27c9LlFJCdKx18JwRMkwqVLWJqOcgg/Kwi
pbiQdqhBeBNdg9RQSWyUvu+Li+w4F6oxUZgxt0taTyGCPunrBFRYlCGnJV+z5CDt
PjeXFHIUDEw+WvpXL4wUgYNnXTtBgJEx5qAVWPi7YL9r90WI0Fa5VR+O15/TUtSL
D6txwU8rn8mambBrxSeoQ5SmG0Qwp/fj5Q95kqp7RDktUzY8x/9B5qSQjaMxI31N
YS3WtQQIVlXPNr14QXALAnV/44zodKJixD4z4/46O4fvvaw9G7t7ulfEaU4VEpij
sixGQsKNk0D4VMBa/V14Qh4/0/CMR7/7jcMISyN2A6edQig2l47g+qDTbbz+G5Wx
IuOekrTHd+jROYYQkxWpXwnP2OlO1isJh7pZFqzufmGopv/xR3uAO1zTjBafhZLH
ZYfmocRI3IIPffFALko9Be6yzeeEbjduC0096Gfh2n/JEXl1lXlaTy1hDREogQWB
tueTLWbtn7QE1yQl/mGbKn7+8k4uspfRpoLgeeReBM9bJPov3yIWD5uOd3bOoWQk
r6Uu38A1EHv9zGiBV7W9mqGXGmylZrABXM4TgaR9b9lHrMFMfq0kR4shM5wm660L
hTtxhPWMv6I1R0K+8CpedJ8IKhxWe9AbKT66WSN1yyCWC9IBYLjQhhxsbCM0ZruN
tOEEA9Q6d5LYrtdL1RtZNg/g1+kFAux8lu0vlM5V49q/0renhe+c5CTZq3S0QjPS
InYG31WoqKwVCWH8Fh2LBqyV1L3y4ZWMDvTq2PdxXAaNgSGs2TFdiHOdUEkgOi1X
vB117nv43jcqGhcjESZdZjn2E4H0cEO8uRB21rlHYE3criJJX4xCMWDl9GoVIhjp
O2bdxL03iz6QpcU7Xqx4iLI+I5v87QgV+gjsJszacsril4i4wOPhfbo3TxN/8J28
ApvcfzWe/biFupLhUxFbJkwysCrf5fhEcXtbWxGM+odHP6FQA0LGO0oiFjfaRHSV
JtSzG5rJQoukugkEuWLxQjZGKGAAZIqnB+c8sH00qYNgfVXtWB3EyxLTLvd6xyxL
bCKQuzrnYA1Kxy+BqhsW78jnKeftyi3xjPEUXp2ZW0DJXE5MkWEM3pYOYn4GMSRa
KPv+zxT0WJawahyAKwolqBnExK+3ljfCfD5FgLJq3eV2j4CXYb42b/O0vb75a4IV
HU4m9uCnAF6xpJ86Vz6Ni4H/KNA23Hj6kCtlG77eAyCs9IZ/cuaW4myarRYPdiAw
6w608/cJ6gqNCN8mopBe9mpfUa+0lWgT5ZJuPSnviYKx2nz5qdr06/nUy1TVjbeQ
QKDzvVOFG+rIQVJkJsVghUld9rSBTEmIkL6D7JrISwA9ru0NatB/XD+zXcWnJg5h
bgK+03mPB3/rzCuKm/whSYLlbSUQHZBOYj/h6OewaF1nvNe058jNQgfU2H/3RlLS
kUNv6JtshZWQ1HPYPUsLov36z9LvHY1MNRkWeUm7g+awedhG42kvtTv80a/ZfrQ3
T0wxkNA2lp2Gwgtkz/Fdm4iu78bkkq6ThsEyGKLDZ80IfCpzxVdCw8T9IKCecGUm
FHahsfpGaYhnVXxmQbcHNgopH0Cg0jTemQBIOlvw8J96TTrJb600jFSMalm2Cm5/
6A8fHl6W9NXEJsGcQCkPku6v+sPQP1pb/7pgKmnuAe2Dfl5Au7lcjEK3nAXdVsTt
0R0Z0nyLKrby6Z4Lh0Uu+zuQAzm2vbofgN6QJOj/97fX/O9ayItEi1tx764uWjjv
/ygSINxn//za6MmjJx/okBm8P8xWI92wczhjMjce0POBS0zqVl8SiDv0/51PDTjM
mxtKyRMIp9zhmMAqmcLFHhztmD00+7k29Iw0EYvsZ76ODAbjjaG6glWTy2+gx6KD
H0j/yn1Rq6kIyN5BmbPoVW6m4qRpL7zh3LLGK99iR7+LcsWoVFFYSNwqe3n5oBnK
vnrxIirIpfAaZCMzK0OhE+1DWtAWFkitWdxDJ6IJY9yV5OMpdXJmHTO8RiQQQbNB
8k/qZbVaVVTFmafdAWEkPVKTAXdqtObikLfftPtM504F0fM20VllEr/yk+Gwh+pb
OKIVDForCSvaCny9rqMH4C+byKopK2hoXTdLt5mgtb7ZMUf488IzDhvB1y9ij574
+2/jdvE6wFgWxhRQQaRMBadmN8PeqXn2idkOcy99/L2BH1iL1XJSMbQrrexa5cZE
gpd31YxE7/WkJSoHcdZ1Nb6rB6ziQstTzVP43eNvFGsDSu06vlwl0DGYmRKSVojO
xCLx+fthIXYDhvHJP4ppihccuttWf/nIcoF0W48bMyhYDyhrnc0fc+Ufnt7lKGHp
pVxLFEHJSxQUjZnQkZk2u/nDWteUMcr9neCZutLfPiBDoLCv7sWDTPPEQoZWqrEZ
u0fBTbQrh1E2PHyonRixPXpleLtkDeKwoPtYsc+8yv2JljUSrcT7l04FSBpKUmbH
ws4DlzyrOOW8HLt3dTyYMjyipfdddSan9F1dMVX38suDkBy3MeG5U6xmiROFgXm0
J5WqtNqvYsErY9Rbl2Sn1DPkZz1OjRBYGz8VFIWShsFdRL7uGN++Rnsz7TadXG6n
4UvEEjD4tJNWNGl/WumJoDeYOz0LCsg+BRThRbBPtMORRU4FE/flS0OnUAa1P5r/
fZWGN6HePefAF90j+7PZRQOFUWMFamz50hB7Uoftv62Ku+5ULcGKpjDXOKMdX29m
8lD57MMVaBbc9NZS069UNTPCxBPXCF4WXxYxYesODPGodBqSEfIYXSrKpRMnp5SW
VHjah1lMIwEiwihgjQMfnglk9TNCvS/pLyRNPqslG8pp/E/WwnioBeu8y8sITgkw
IwK2qiTG3rdYP8uJsFq9toDx9Ly1XHrx1F338mzv+qAVUxMLfGsZG1k9ssUY+Mtt
KSmwhi/j8+FU7C3RGYPwRly3gwE7UbWc9PbShqpdVM/5WRLXYhul4VdDEsk1YbS3
v39+szjyjL90v3re8nWua3X6Zni4KG+HTF+Qt+6f64/UdmOiOYW8Rh/Wf9qDnzJj
NhpTIMVQ1zrB540SjEYSLSQYkCPW9VExi+ldGtQOKJLX2bP42ovzOwSwNNdiETBv
I/CUb3E2UVuHCRfsDFffJ27RYaL3qtFza6qUrB2udbIlrlyzV7XSvizBKlOoSYUL
EIkmRLriDc64hz0hcF2XdE9AlEUa/Pz64/G1+Q52//awoqm5M7Fj9QCli2tWiX2Q
Ni6KluOJiuN6RBOk2cT8QpcyUe9fe1MGLXHYHwj4FxPMcTTE2OwcJJWPt36JpaXl
HyeKEumbAk6+xgeYBt+dOu9+F84XRcQ/I/EIZ5G9RXSgGFPC8HJJsh7n3c5vg4kv
l2wYPEi282qJpYHHAB8PvQT/AxLZodnT6ZgpLc/hpLyxrgPE5dESG2GG2zGhPqlV
BbZtfdJqa+tymIew5fb3yrNnqlke+aVUFK9WES+tvs9FM+3Xc6x2bREW/YTcVzSP
vnUevU438FZ6u9tjYUDREdwFun/TdUXl1IqfFeXVD67aNPyEnKTbfnomCtRXSL+4
KPZNcK/J+jRcX5/EnCszUgI/Ikx8+GCPEsH7InyAxMn2OqLT9PDU81vplaX8NVCS
FL6RihdZgACAuULAe1Ipr+sdzvenPV+nWQ8oIkajW8LJcKQnyXbSJhuafAuoQ8YM
yH8pXXkQ8zYHsG2FLFZG6yGLjEBlyc062TRJ2OwbTGkE84jfrcTEDQg+Fqq2Db1Z
XEn92XoHknEkaL6Wd1V+Ka7tlKs+VmfMjB1SXqjt5+J7DBYoQ/K3xhrWczSXJIt9
dGIUhiyD4EkDHbhd3Q8wqAIzTj0mz2PJKyMAv8NV1Bg7ikV8Rh4oNCcx39voaQje
ryi93p3UPnAwUMzg2KqJMrbiRIfAJ9o7QL8nKp+Kqny/HgeKl1nTFn1utHLDJaFI
O/G6Wli+sISAc4JDgw7kdOkwfO4D0srtggVzS7pIkm+UOiH/48OvYFOJOdRRMAOR
Dr1D8cPNrMN8/EYCfJmY9GWSrx+6o6fg8xiSTDYz64hfAc3vd/wO1bfKhGKiQcE5
qWAVAUuM1aMzXatR6kh4sgu2spLZJpiTrR27J8u8LF2eDvZVgsY/AA3Y5HjRF20H
rrSk/14Fn+hui4yPseGJLiqxktiH553gjSnr1w0yH9g93lp1GXXvW+RwbqiT+xXO
E/TxkRIjtF8RM/IPl3VSP6EXoDnfqT+k41NHE+Tpd81TrEyeG1inncDBr+XTiG/5
xu+33MVa/ViX7EoB4+6AkD4rnBdp9j9X0o4CraI3+j/Kf/loMNOnUdYlPdVsQGcL
J5pCFFGGihJAwL8V338/QZJLzdG5fKILtmPLuI7SUC8NMH/SEaW+eoSLXQKNu+HA
Grud8wJcvle8Uru5bZ4cOzJy2Yhe7tkeCVU/UKnxnpsD3fwLjVuEmUoclBrM0eXO
yGrpFoZFMxV2hAsAGoY0/fz5crQRKSJ4Ekp4LV4iLpFaUu+6F+gzJxaks3BHQpz+
R4cIM3bMr2DDLAVi0cRwfRyHoCoZNzGwBTOOHTXqMaWVGKG4xuXfGLDAzCelwl99
8i+qCpJnWULjtplV6SIId5zTf1pnHkfZo5m2aL58JwW1lrHPqJKLYsFEn3mlnOHM
Bareb22yW/xJ+X4+2iL+LSgHdoCssCe047vU6k24DK4U2DXPprKEC1nMSn9A/wEI
2SlE0Xv72W6cfUUHVMbIbnmOLWN8SCs8IzbSlYDEfKjCDIjx5tv9hyj/1aU4Oc7T
tRnPX09qJi7Eotg5rgOvaoQoE4SLb2Dt02DCOdaXBl3VmiGy722PxOGzqsD9bgKV
PbfcviqyAJR4Smzzla8a/PRlWBwyg7em54mmvYuSTm5iOIIl4R/bZibzqUx37oZf
p7BPskeR/VCwE+IwpPAOchJk980AyM0dX2TE2Yrl75ZwMu6LMzdBhjJVZU4I3p8V
Xvialq9CzAxOKdzQY/mMhX1TAezzeFQ2FEPpPEvcQSIk2Wb+8Gvc2ETxKf7kZsko
MS/jlVH/F3nEyccnv5ApsOcsOAwxhlGOee7mpEJ9qTKBcKbiUuK7X9dY+4bG6eQl
cSKqA23H8KDYcqh0uil8T/UOnOoclb+ViQJefqsE6E0kpEUeqTZbHh3fhTx7uR+V
BnBXACxaFcayObE5utU3VcO1uMTSv1UWJ32ydzd/3c8VI3+bv7dsjiALbTEiTjbk
iqXHaeo4RqnocQJwy5/tc1Y5JNRVWERQXPLciDy8Pd0xEuyaqnKNm4dBzo22Jaag
hhkV9ngmwjmwSl+jOg7UdpgTQvZYJjR0V3B5cFFoSi69eOQfnJLTOU5D0U7zNJxH
2i+oH9TNlKFEEZP4+5Z0YcHMu0dXqm2mfcoOJ/f/41Ae9HMW8xsPnRTgSLDydvvc
AehsVp0it5VdIC25YE6QtVC5q+GNsFXrAZZPEO0q7rczfkWUFmz3YXBLR7h28h61
9W67axdUyTIROxkPjiPuUb5LzF8UBpF3Zmq1Y/gVWAKJ35HmbRNlUN9XLpF9keBj
1edROEo6xlJ9M9PGfJ6/vGjG06YSV+O2KJJ0KbLIxjaFoRDUZvk0DDib3BJ6YrOT
cf7NYpK4jqAOMdb6itfd68jHK3uEtAtcyON4NC1LPrUIoVpC8WTRQC6VWLZmxHo1
eA4JF4e4axbQ5DsTWSbd3seJcfry7xTSPjh/KRsRq7OglYJ0cbxCrI2iV+wXPvvh
d8lN0UvqY/5KviDhn3iNA0UmtUvd8UsQs3Fw4ddis/8cIsyKsLAFiZOKeFQ5UoO+
ol6VGRaeJ3Io35K5jc1snzJoi7mtdafcsY+PnPq7xvb3dbXBcq6p/W+eToVZgq4F
/EEt0uQVNQDtSMIP7D2tTi2MdLhgxaGD/ioFuZkYo9SmUAgMRvKBFzCmbToSQOSz
oi4NkRx2uDaopAgUYGY6DOwfT+SaTlZiFLWXcaVRcsjOq08xkPsmTqm8pr87lVYM
Xd0zhnWXTgPwz6epAuid/Gwtdt+P4JdBcYf8sDZcelJ5UM8q/IHoHO/uoiZoMKzR
aPnhRKC+UCVqS/LGcFmo148t//L954YNGHD2c07V1mLj29mnylaH4BFUjOHzhye3
A/C3iCBHrAUmheK9rWaW31NiSbncBs7cQIQWdpR0VcNRX8FscLssMyFJtfIwxTf2
XyyHozK2bzgCEExYzSVCXroLzI+4alHcPuCUYTxEy1EI5lCX24aUrRXkSU7TD4bq
uPZD84rziRAXcvvKhlgFayjQqjU3I2iHSnL9rvEsLKcVrylsAI2xqmmtevVBLYFj
1TbVxHFgQ/83JbfhpJPh+gRg+JQarYE5Gr+tGyJjul6fq+i+4ZKokeQSdXLZSrZt
0eFsxcYqWv046NYB0r1CG+UE25ojeEa5a6tdpRaOGRO5NCf/1PElT7JzmB0UD47I
/q9IH/b4M9jlpiHIJ80NUQVXPpJ18TaRvR/4y9Ag3tKldst++VEEwWa1yNJ+Wjoc
E6BmT/+qkzb4OxDqGxi6XkJ3542vl83XarI13pOn4k4ivpx8t0OsLVnvjm1vc3AW
fMoPcLBS5X3HuFQC2+lwehGt8DYPYujACoe++nzB3LuD4AG/EYjqbbRgLpUE9svY
JJGsN8XknPnSgUtx2eS9I4egjfuI10tnlxCbkQZ9vqybheI1yy+jzkDXBxzxUwPr
nqRuw9x86UaamIJMqJx+f63fvouwznGV1+9FnvA8Pa0GkyhvJmNpECoAxk8Ik0CQ
9XRWydaIgLcHFwwhSY37EcBjreP/xtKJTAFuJVreFwlw3Rq0SKxQ2i8xOWOoPDzL
SqInEFA0DcnLpE8NOUvMYMqZbxb5Hi/MFXKKM7kCB6cu4icJNFsC8sNzFyqGIcvu
UCyJojDk8RGyp3cO+j1XdqqQNwfXwK50YNtEuyNWEKVINl1jLUFkQVNyF3CUy2Y3
GQdSYl79AuHjIRs+/GaiLlPlW1h5Z6sA9lNnzyrPc+I1fkJxsEWM/aVFj10co107
1CY7ZpEZ1rOz2CbI1FAh+4skrt2nAyaNu+7X4o6Ibz4D4k7k6/rhrrLQIxy+CvE+
iaxDPEWFdDMn0I1PYb5wH1FmLGfkGT2S4HNu0YW41husenb53bP6z6I3asPkVMA7
Wr1/6LiIBYnS2RwyOnz9qx+BIRRMIj4hzxwGbZSs+8AtodqJZL6JJHjgm4qgNsc6
OnhifTAd8JEt/wzDQUguEzMDunkXzaicXMKixCguPlWXqAunNBCMHAuYjxDlP2cH
XGaLU7lsLuGLt1elhs/nBOSrdTfK2WOzvlTiJyDkqdaBvH+v5igTHk86jsLB6H7U
spwKn3AmbUd7vYKLOPD+pgNrV4Y+tgsjuMz/Pxn8HoLEF1xnH56M0wgJBLM1s/do
wGHkAmYU+pJr4EMY5aCL8gXITE0xzn6xdZD4v7+CPMuD8c400m8wGU6CxUtb1OKS
3hxyFNya67UUCw44PdzpRuCjfqXqIPglaT7qb8fJp2JKj1/bU1gl+qRlw44cpWDW
0/ejH3Dl0Vt+cGjk7CGMGgCEIZ79Q+Hq6P7FR/KjToqCCzpXZ5JVJIpvmJiIQ9T1
ljVnpBoJpl7kDEtrP8PJfbBEE6CS0ULuUII/gY/y5vqbC0yBGWm9xm2KXZRHvBOO
oSWevhhNm6hl57uGrff7bNh4i45ixO5dm6w/wvWTlmYTHRyd8OjIQ323qDx7FdfR
E+htmsCJA4yl/LTeOShiBUS8nBivMGfcoPSO3xNalzjY93QLrVUmJaCkLkTxfe+w
Lboed6WkegaBsP8a/MCXMHGAxKFSvZAY3K2QMTaRgVJ7MIX76cLDA4UAC5aIr8C+
FMTLOlojIhc0eYXzsVkl1oJj0Hyca+XuCllNLFLS/9g/zS94uC13BJ18Wpd4RTBi
Thnjf3Nm3v2LSzleLACUX9V0PBnmdxc/DEtMliE5LtnesN83su6tlmQCmmsgcuB+
cBh4N5AR/UVNbIeGWLqFE/9PLUqBDJ5ZoRLdx8961xZ4qgnu1EGTlgsePIlBXTnl
gyiHPWJyjzt3zpFMt0LfSDPE1b+f/pLaCpOrGrL69g0Gq2r72EG2c/1fbwTe5eqT
Y9F0tfdYCr0X5MleTs0IT9d8YsqgQSGF52ayMmZig/Mgx7USNJIBgWw/zz/IctD3
Xow4i1wsh4C8WE2I2AMgLq+jnyMIkiwkZfEPQqPk+loFY6Uql1XxpVwgbFKrqPJO
p3pZgUZgfsKgFwmsdyEESj+TuFWvRo1Htehjhz/GWgS6chuEhbeVryJh0id3xVdU
zzPJpTrvb0O6xC2/FFeAFDALJRIv0DJHzdMTIgi9izSbBx5ZwYxzvw4ZD3lPBxN9
Ig2tKnqBrvV9rs+SX/iyv1f/gYbfWrgv1pUVJXpeOnKvSbbcSH7s5Q3MtOBBbsV+
xtBGMFl8NtGKBCTTlWBYtkVV0xRagOOhlQCaIL4Ew68eQb4BZar8P32FemKYIH67
7pPrcC3lLgxpFHXFMOCUWN7u02zHSHJiOSNud/j2MOYKbRWaVzCTYjlXrUJi9uSM
9fiJqYKF74m9joKp/26VZzY87SxqysrcFh1nNTUZqNfQsyuNLJvtqxrqXaqLQbop
7YvHXSQoFZ0QLVGrs8Df5YN9bIS2j0GuMjGuxc0SXPnLOQAvQ9+95xDNbIxtbmRn
vXj3DUx0Rc8OYwV6aRx8jgLyIqRBIW7uGdIqmXxdBba7c+5GtsAJPbFDHrQ+jHaS
YGpmnxg3uKgHPK4Go4KUEj+Jgt4r0sxz0aF4Hnj/lteMtBjdJ5jBiAjSKUx78iQy
4syV+afHsB14GeBtRmCuNEuKMQIUM8qXQBLWJVcfH8HxuIdwpu8J8J0Xz2z9FUbt
PGgL4zNP++oNCIaltPYe17viGJOLo58gWYLDv9akQJvpweXXySyZcSNWRLd9TKwD
Arh4n/dgyJS1nhv53ssDJ4ZuZkVPG5ps6mHHY6hbOT75AuLeXcVre6bab7bQn9Rk
RDc4d0wqEvaAqUNZzNxs6OiJWaf8zgiEU4GY32OSAna6WCDHEthejw61xuU1zm8V
DNnT9w3WSJ4yAvPqd4V9o2WETyy/eVRyjbUgZShPJSc+XFdL3a5gukXVxJn9ikG+
cZsmCDx9HB09dDGegFS30cNrD8zkK/vKwg8afoLgRh/RT25SNfZ5YahTx5AaHDdo
WsPwJ14C7JU6P/Wqgdt5I5f+mY0EgeFM6yV0Ural5kZRePzgi0zul8w2+RPkqy7o
3UmDYkGi2FQqcyK5fDHds2VvbeyOhiOIGvBPCTdH4OGAjzDQAKDkQjNkcahlM+Vr
VCJxsdN1uK3A8gNK7Q2x7dT7qkfjEE3EPHWAre7+5LXsBNsz5EWIvKFb0/9bkxZK
zX+RTsE3cFkibxo+AWMBkwLyLgdx79F5P6/Cmxa3OzMjjCDbSOnBMnN6vc8ooa6Y
NLrwGpD3o6e5ersZZOuGGL195ttVdcm6FzhL8FYHoKbOy+JkKTIwK17mkvE+ioQS
rZNzhe9SNMmD62Jydv+8h+/2qdU/AGbUyt2i4ouxUNSJHAa/ObWsLkEUsMXLWt6L
rACmv7mTouaPw9oKZwcFDUCFiFOv/M10m3JTTZGc2KvmAOFVe5XTvxapY+VQBPIC
ccnMsF4ovhzFgVd8Tmi88tSjm8R0Y/53P9RPR3IexwOSzEg+oZodfuX1JzR8za1D
qMtDcDkeRGYPFcOEkAQ/cRf3CvkG5v0KnT+WEygBX3SvA4ouySJJKKY3sc9uKTZF
9viJZxotsCgopXtW+0J9y7LsjrzxzljSpEZ3ZsygR4JwR1SbxE4KSFD37tPfNIb7
S80/CPtqCiRyBMM6oZq/Hq9ZQXpkTYYU2oXAbmG3upuP2KsifLvH+j9mwcC5zR+5
4zKtfn5deCWJhH3fTz4MXH8bdVP9qLJGlNP7u04nBM15AtuZ6sZ7naC91Ry96xro
mYZDJQ7gpJ7m6qPM95e37pnw3YpMEleh9QmnfsgRNKQX+iCL/7SvLmRYo24wdAI6
h0E/uFBzyHA7ja+4s1xTMYfxzZDeqsc7jOYQx8HvX9NtryDZu3iLnWDRXNu/vtxV
RhFRl1ZNzJZP7xKEM851m0Ddo6jAnpx9/OLCkcBZrP8LFhLcVkY6ktPmRJqCihHI
ifga4YRdah9onsEteayHzLHn1BF1/XndKjLg7Lm+GkCM6c165g/XKIYtC3jZIj7M
zTnOR16HAt9O8z7M5wGRaZV28IxPO6m0Fm0cab6/qJb3F91gpVHnydkSMpf8qqBo
0OIHlrNv9lneGIkFU+cuEGRMIRzTijJq84b1vmSOd2Yo0zhJ+VH1T1XrA/0eU6pf
XJxrD3D+OHrhnKcDOBn+tjrkdQQJUvrX2J4UqsH2ZnB8/rRuqBc5WfxwZz+FKDa2
Y7VOm9HexTEuBkCA86WAzs/BGZWr2SkdaKriWAojCK4bnZJVbPVKuwPVN3tHiXh4
qE2nSy7hqjHJlW/Kdy5OTFWC1hibmtOMPHk/r5gVl2iclFBK+jIhZ2cWDbLatf9g
XzQ8GIDBoGB38rNgucRzSuFTG/GKvAcm28mGge9NWDQ2RmXIFajW0KN3giO+e2Wr
NzSFvLUzHGHwez4IJm7UEyxMYB20F8ZR36ERjqshnTMVn/KVTsQ2EflTWOipwLMW
InSbBT2DUMDiZsUYXsBHOli4dGEuvTnKQ4xc7v4L79ey5amMnPgX09xmuANefqga
q885l0RiazegrqJ9l6gpLU3aYmdgNfjCJyk11NmAnvKZ9Yhl/In0uXfx+6JCnG2/
/Fd352pfNJwRBhmPbiTewuXMg30X5ypBVU1rAvCzppVRvOGtyq6PDfoZcBe9H0o6
/TNYUPoWIvTJad1+5XnTaRSWsBcjaGDgL6joVQQ/MGUsKvbLHUvdlIlqe+gi243/
/63+zGPD+JVHeuSmhxgqfyNjcIKFZ5zPgW4j5EryjoK/m3T1nsF3MC9yZeurRrie
NX8vRR0XmkrIh/eCYtwfuguvj1hSc6ht1O+dtWZGOQiPSlAvbZT4jfaOh/4EupVI
m0gjmFjAhU2by0WPMiUJfYk7B9fWqbJ4NpJrzhDvp4ElqWXd/NjiZRSXctj8gKrk
zWRdVhd3erWewWuP+y3wVtqBOlvn3cEBnSDW7u2Z3tQP/zL63xAmJB22YqENPI8z
rj1f11tAZbXl1uWnoEGRChV6ZeC6KMFkL9+X6KAwxVWkzByea04uGQhgDOr/a6lX
y3Mkdn5f8aYdRMIj8rmSHQjteCOQ4iM8y+YOMlphoV9O7btEYsDYjYjGKTIsfrGy
eRkkF0Y+wPXTOVea5EWVyE9Ia3Cb6mXEMOfrcBXWVZqtaHREwsMM2MVOKvjHxbiv
1fW66mxjX0IIWj1DWnSE5NTp3WtSyDzhxpbsdT0o8al/TGmcUwtgmT2J35O/P2Fq
zFKGIqFsoBrIm4oi8szqkllxqvY6jU6gYXj53esy1eNbviMz9EEx+ctG5qSdSaAU
YuhIUV6wjRZjPWl8i+3niotRict80fMfQl0bAvmYqFOeocFuR6qRMMRc5G4eUq17
8KgeBrrZdsVsBigQWlg0ia2hold5QQnbrU75e4aZnOVJ/IsOqT9ZJ18Hla5QPjUT
PtpDX1uRieXCzQosRl7exllUQp3bA9CsnRX8wJpCSrJp239vs2vjVFpthdkd62qu
q9RcrJYWnR81bVXz8ZNpgp1UKNUinD0W/lohoidbo6jJlspBHg2V3CqXUFOsnePl
TZ1+r1d7Szsd2HHyViu3SDBPGcwBOYBo8jFAO2FIGoJQ2BMmH2XtwLjLFQWqyF38
MQ3ICyTDsk4D6XAUu4j3tHOXSl7vkxFrpKW8+0v8SoxhoOBgXDucFDDkODkwpy8G
9UZDQIgNiGw/A2CsKuZvk4YA5PYtZ+ZzbAKEXu8C2F1ET1AZwT5rEclMN4dz7QA7
3B14DeWSso0q5QUDo3AtB2lOsAn5P/ryqW7HEgsP0zxxI5UcKz/7O/k/GP008d7l
hA61v1puCTs0S+w3jT/uTSN2p8R5d3f7QwGZACcR5049Tz8eF6YLWj9+UnXY4yFF
4TpG+OCAzDDNAnmKNmMobGVYRGYuWtxO4/jPdu6w+4BKcpz9GDgpbk03ursT8q/P
HjGIda7YjNqipdUYbg0VUu7b9o5mOBK8Q+2+oRj9FVQ6m1wFi1ACa8pStLE+w1gi
BNTVIiLVICflmhvFrJF/0/p7oJV8INKx0jDpOZ2rAWAHdClCxtMdxVOPSs3OQM8Y
AyvNiAy9u7/Bz/kb2jE86c8hs15FOa0UkV0QW823pvm5v83J1a3SrnA8/ity66QC
ouEtlhSi2Csps5IZvOiO/kdTQAmIV5U153LPk2AA0etsGlPtFWJVn+JoKajRnZR+
LZkIMlc1gx5UTxAGJ8w4yiYyRiLgPGhKDzc8s1d/9C2vakOE7rhbIlgFxKHAz1KA
MzrzNsuwzVDzc9xBduUKj6lO1YIYeY3ry4Us9Y/O6oae9x87YIlXTTQ0dsrUy8Mq
QtVpnfRybM07I8WxTWVNVHiPuZXwzQyDp1Y7BRWno6rXdOHTey7wSEEnnTU2V1iE
J3y5OCtWSEQBtANjW1epfWlv2iitumulU8U2uIooljjH4D4p/TqRbn9oQlim04VS
VfRh+Qr4DD2SyRLjuNJxG4S8ylcHapZslV3LNoPRJ+t97d5GguPBkHnDF5JxQ9QF
fYNzxTVzTt9KMLbchImloehTOkMwrN5xVeeHfIVFsgvbwX0YXi0WozfIitQ9JrX8
YNmOMuTyfglvApAxkutgeytmYEoD2HXj4pucEuqutO+aPWNzSowhY7StlVbC/yA4
ZVF5aJck7gpgwUqWs2qmSuP+En0uFbnNDfQxaBYYohING8xBnYz9wt2LlgxrnWCh
QtqFy+GfEc3DiM6Hfra+a4ZVrcx75YZmvwRLPTNpPgY0OXTIwHVAeo6MIquklQxI
2CEcZq3NiKOVjmEwoaHN7ByubboYEySQxFz4BHODwSs51RRf/mIQ/FvAvdYYm7CV
SmBDZSD/Pi/WOlCbrDgmsfeWHOc1KIPa1w9PJCEJE1DzwkP5KBkxg1oeUeHJk6yb
o078YoLucpKJ43ni7WJY+VBRi8TcZnVr7vUotpgyFlLtFmu0bOuI/XC1q1tVrRvT
LmYnl7YziZW38CkWUj7l4H7ukZakwtwLOkZIwnh+ZhooCgSnUqieXKhlhCwdkawx
3XIwjPv09lLjHwFFc/ailwBTkA/NvBGQZTklXXkHJhaMhPevREBbDrEdWoPEeFtu
ce5+9bvuhSM4kthxi7w07o8HtQoarby3Hq7+taV6a7lRPH8G5EBXfMaR7W2eQcJP
00J5ZqLfQMgH8zEpckLNLHvK2JesiwsozPDVk6Q0Pi+tqkYMpWaBaC01lGM0gHQ5
z3nkTRGWwgo6KlGagoxRZQidOZQtpNokERanLjLpnZ/G2zVtkchtEE1IF76Qv1BW
+bFsj8MkQTIOwfLLmUgLMeBYqJ0AN0ajvjY+XblWl6kQapNRD6xJYGzEFykMnOH2
yXQmD5TibsaWKjzCScddAZWTXA7OLAlwjn03bH8rHr4i6KO3jOOEagYXgFCfoQc+
n2aq6O/wascZcb1lUi1CJSUJHGKfRglthG503CbQjF5VMrNkFe1rGMGFMb+bPJ8E
cz1DrqBNugj+i94ryeE95JtNNyUyTcEJmaioXv+ToEqgMeCCALr+geME1vy1/Qkm
FbUgI/fvxr7KXicHzuaSp//anNMdFBhLFE5ZnF4mNsqF4aZ9EG5BWZqbifZuEPTd
2RPnEvup/z1A8jkNRpYB4ertP5G6QKprX2BtPK3B2L9m7goJ+FpwUNWqjn43BZXH
ISs1f/5TM+mJGtZEwoQ2WVoUR2gjdaVsCl7CEMl1u1A6yX7vLEyqmE0EpYtZoUzs
19OJk8g7DZpe8yyJ5TLpAjM9HEmZ+QDWamy3rCcwcAlsNbI+1rMoEYswbZm0Tf81
eeUtPBomr+dGhegjtUy3uvR5jkl1TwmkhjVnwZSkfOlcMJtC7Nknpzt6efEwbG/w
kGB2COtcqPWMlVOfOmwOUDYeetZGe13/iw2LlNvwAOKhbv/pqt3DIYzSIICIzveV
lInt9PY1/ygX0w5Pfjk6PEO4OyxBu1YJZmTX291RAB3xfUEc0onHcdzZcxtj0IS9
ddNX4ZB/TpEEBWUtGCqPojIa9xdnlFavojM8fXT2qXOI8XA4HvzizPKQwvn0u+7A
2TlHAD2YZU6FkzlZ7+yRE8PyviJ7KhT3RguMac6EpDsWk1Lm45QI9rH6w11jHJs+
Wo1zFDE7GQOEeF0+DZKbai6yp3xCdAjMrb/XxvUWP8MGnhzCO9VLdz6aUf7kZ3X7
yO1Omglr9NRcH/SrQ7lxX1HcokfJonnRBAAr7Nw6UhgPdbhghsFV3rhfabyVHHhk
k+0imnAQOzrnPxKs64I8asFSF2rzvmWuDLvulkYyV5VIdF/Ghe7J/MpwqXGrH4HN
dFqbITmFFsIfl56KLpZ/Fsv3CKxfvo9oepYMrB3Y99Fug4vbY6wVFrrPw8bDrUkN
jhA4iDy09AULsYAdLR6emdbCiu7HLrzyk+2Uxq4Nq8TpPrD1Aaokc2169yxK9zAu
1W2wSwdlQ6z1WYjPuZVMku+2iIr+HLyj8mKX+nR152eJHl5frXEUDx8cxbPZCmGz
kCJNn1VQlnI1cOf6ZsL1k3/AxBSdngaGGg5d0rg3ouM3ckyAVGHiNY3SMD57qTvr
/Azck+O/KqFohT6oqMvYmjnwP2Ut6vfcW3HtXHDB4fg8JXmsI70sg/iNjMXGySS+
4lzuIzrrEIcOuO/Wl4XZaWiYR9PbwfjU7ClUyrisf7O6nGLpYReXpXJo9DJ6lRjo
jxHmd836kWdwHLELx7QB8WLWepRnv9qZdzsn1R8pBQIEv0mM0RPJi7AW8r+B13xc
oBHP381z5tsMnrniomNUAWjYxes5Wsw45m+fSA6lNJ50wtsX4QRS9hefcrnxGDhD
KTCvLUNj1EzOti3VG1GPFB3eyGfheRfedkw07DzFBrku2K1KXuOBRAuhyl5eZZWm
DmQYVcIF2zLnGPNvRjfapXpoMLa4kUibxAwe5ar+Pl8Z/cLHtE/NgEOUqUP1lmHA
Fz/jz4imGOCUKr+zOsieiQmaSlntP0mCN4xLJ1z0vdTrD4EO49i0Mr3mgWxRyQGe
rWdkS4NFW5YseIR0km2eniTlOk6/gKeJFE0qIujOCcZj/Heut+2RghllI3Rja2u0
32cen60+QlCu+ImUpJ81BmMggtmAONGOfvXMJ9dyjwio+mtSv+UMIf+UEIHwCxUM
PK9zdAxuN65fkYTrPWAk2/u5s/+/jCuWwhTyijmAi2qDWcvz6/MFCK23sbk4s3Ip
Xw+zg/Mo86IKt7YXj01FC/z1I1KRKCT+rGBxnUvtCndxt4mzbK4fYSiiWZ1dtd51
0nxNC1kHafNWyzfdjkrSLuHxl5ab97jmZpQwk89eGAn6pP/GQD0LtGdENbBrqMJD
jGMkiMLlcMv46ELQGis3J0RvIOy1f6EjLOE0LMpX+/x+/1rgejmm9UPKbiQK7PJS
2FkxYkY4q5Dw/J2N1JSynlK7zCO0L3R95Upy7ozoNjapNDiM1z+1R0ctuDR65MUO
zHyDhsvyZW9MAg/brIdQx5kmHV+rz6tKuEJHso3gAT79XCMGTgt3kqlkwx0ju2Gs
E5vfuEgZeye05dRf1r5veifD/OgPhanamNNjC9itUTC8102JEp+CRQEtp7vi+pP2
e5uxo9dwBNgLoy5VVWPyHCvAHewDUQvMrs1er141kwk+oG+as5olyPvgKEHdHeIB
rYnJLAj7brCBlRospvpq0bGFKADcGg+ysJELveiXR7P9Odb/FJ3yLIFQ01LnAFgd
IQIlTPHusK2GBmExxT2QfOX9AnKH1g0RMEZqTjSE8UePdnXXWs5Yp97IK4UHl4hS
02ehPpEf/KYnFto/mKl1xKHSWxmQZlA7Szi4yWXB11cgERHaAXgu4T2IqdaUuoVo
YJ4f3yskj2dpc0BAvScHk12f0r9KLi4NvINKMZ9lpgdf9qHZStAKp+IE+/dl8Vhi
FzcHv2TRT7dXwr9UPfq7HSVlYbD/AQGiyI3U31/5H3cMbs2Sue2T37uxccbs8WpN
t4w+HlyYXJEEalNKwof7mSB0nZdfnjZMtYkL9mp0f7sqxNzLad98NPU3EsjiT0WZ
Dyoiuds/oTiC7wm350ea05z1K0EDNCx8jYbgN6I6hrjS7U0hoKDrIGTW0XjFOFXA
P8DiYmp6bSNd/UKJChBxYm9em8GJ6vt4n9J4oxrb2BAxToIsh4Je8ENuHrQBeL26
1F+QSl9bLS3lB5Eq77oQZ3rqnpyajmw/Q3WkuOrvNjoSz9S2y6LhkKv0pQR3iDSd
r2tAKPssbV12nKgQ5EleXvDEsMyO8G3JK6FfLmTmkNlg3t3M/JjV3b4K3rVB1IaM
Y/SVFn6RZ/MOB9sCOK0zTjumAH9C5WWc79wbMOc6dcCIgo60HkIJuGawHHCyh59U
7sloWH2us8sF55mDRQnKYgTDCtMfm46z7lhzUE3R9EEKCd3pDwnwGQAupjQH/8oA
IzDmV11AyDkHQT1qEVSVLAoYGzkeBtsN2sIokrxCXnHhgn4Dy6zPt1VLJR0Lqmd7
1N6qnmfifY8+pxV8vZ1zNUnl0wDJTGxguqpuz+o6Etpe3gzGoZT1Kb/Fb1kQfwFd
tLU9i/x1pUmXfx73pVV1qxSdNuss9fCIg/31Y24/V+NF4X+/LpQeJjupjjEb34me
J5xDWfkX4FcXwXbYs14+iBgv9uLVtGCE1vZlWgrJ7xIftK3BP4GVDlbnsTJcX8yp
JBQzdaJKvcWPRF0HgaXM+0f2ZApWA7WyCVMTWCHkSCOwIlv6+JXFyyFzkaTeX2kt
fx1WtEkt85Z2lSpur8DaX8nAZfe4OxhxnyLv0SacQW6SVwVveRdMqKGfTY+CHXri
aXJS4tuBmoLffqbIQv8gI6nMCPhT0EiwwJU5XsXV5j/pmTY6IhFLSDgR1gSb7jag
LXuqtXmQ67/ITCUT5fj8Kx73mhAXsT21GCLcHhyl9UrQvgtDAXfdxPVRbKPQ7l2S
zQXSF3yHF3FZuzLAYcSMD9FVrKWaHQu7gcoFle5zPYYeEZF05VH9+xnrhbrl17eV
ZtekxLBp79rxMIDTBALqkLh03DyKOAn/PE9Qv1g40uYu8ZIIAz5y4/5iNjeELWat
C6fSJ+vUM7cMBIpKmKJPg4ed0NgXPK+GHb2zMfPY7K4Fei5XBgqGtEnJSDc/ldZj
xuwivF6p2wvfGO2WFh9TpKEBW1f6u5kPdnxssXmE85bX0IXW0uv+Q3xZTf8RqFGl
m6PmjQjENSVrT0c+0kvgurXZOMGkDrtHcJWLUsdGzbrnM8Ni0HzI2rdS2mUbVdtL
nbgWoYAmKM57QRGlhlc5Zomz/z147xQQE/FpRzuA2qIEUk2qGicz7ViuS9j16Ji0
amPKQo4PejJdsLzP4irbnmdGAxp1WEtRJ2NsUOsgq6LraKbl/hs5Df67XgwGagm0
58GRabqYUd8OfYHp3BhadKRbI+ciorZmY2DzON00ZS6MUh6yDxd4tjarUqFxdZe3
R8F5/Q05RKC4JFPhJ+ie2F/ao6sJnMGid1ZkKqgSGpYnnzCupjM+FLxDJQh3w42z
t4j7yBMltfxURLFBxwFrc1A/uBcU9K3iWUCWdHpaBIwz49E5nYRIEQki5uAPfZAd
GBlniz3CmrcCJ6wzgyA+vRk8PcSRY8NS4y8vrmAuNcubgB1qkLb9EZb+mNNnEYuM
ZAZSBkPlWM8ArNFDoL1rb3qxfWffKehrgcp/26rc7s8p2hJZ9uC7Bx3eI3LsaKGr
Sn/GXRk2TJCOylLIb/EVQsNq7E65/4kIHpm7TMHNuFeT4ytllk+qLzXaMt/aggHn
xASjV/TPSFg9AYQHz0qIIEM1LC4YZS1mK6r+6+CyoUxVgwqXzGauWRfEPZFGB21c
iXYFts123jxOE+DLWCW73567tUSn1lZXafu576HH99ow6XlyAjDkUbEweO05FlUA
+sy9R8nnnWx/9DMsm6ZV+JD/dlsAL4XH+/ZKr5XRKLQ8cHIFNFusDxT5cJZ+UChE
jLax4V/uj/7ek6p7lNdFveS4vp1mbrkpukHxUqnKJLN7PXGWaJ7nj7uWwRHWPWEq
WRwehpmGw3HOta/6my4c0q9O3srX2UufQqN2KuGEGU7MyWHRPgNQhIVPZNSpPmBQ
eu7OwQKGL4n57sf2an0ABsAmhE30tKb8yqmjCsLDJIOKtlepkDnYHabXKwemMfIo
l18whrg/ornrzRyDQ+RPjcjNc4iGVVyzfFKRsuHW5CdqBULhm7X5bTspaQ2bG2aQ
0K3WVqjz1uRF6xP+dcTzouiZ1ma3ffkcY5wsXUVOyW0dGeBW+BLiIgeWg/k8nDzM
efN2grNHNMSMwqwUAOCJqkW1S2Q4KdFOP6LNfQIe7vAQAjihaJjHVts0Syk6uBfI
czBKbvGH6nbXg9Vqq1asXoYTLLvYK9SbVPjr5MzIXZQp3L5gjCpUia+XT3PK9zcs
bsK689cMQYrDdBHV02M3OPdh/bxkczJZgGjOhKDxHLpwwTzwpty7USjRF7lMxQTv
bZNe8uPwn1nkKSHQ7KS7MNWshM33Eh0+l1ifQ5hSyPeTfPjBmyusCj66kBK5HDEj
cGazsNJu3GWB0v09c8huQNXC3GYGUoNpTkzkmYvNkOMazoOUU/z625Fouea9yMkx
RSf8uEH63an98ABTvjKrZAvmFPH40Ec0azbChqFxpl9jyQlVrN8vbTzoYxGyMS43
JHUki1TOMsb8gsiuBeTq1wusuRqpGRIs9gjjtmI69kfvUQ1lNJcthiiPA5xyE+/7
wu0HZsGak1XIB03dgGcTrnxzaJnW1Tw/kq6YLkcgZnHAQc0bdNs602AOlAuKfg6N
DFFkowL+6hT1NiMxSE4k+TdBKiAKRVebTSfEBoFoLgQ7iVT/vN2lSl1Y2bF6Sm8U
Zx9m2TcEkoKKu9WpeQ711GjkluIKUzCSuu+ctrhV/Uy/eOkliwULnUfEwHqOjic9
Lu727Z9Vkm40AJhyovb/rK+543g9m3+d6JLTHcK1s/7h+jUGiEJtmHpVagH/5GZq
dIO6ktc3HyTzKDEu/W+qYUiRnByaxAGKQLvnNOzSm649MxdrlAGmfZlCQMDkPJ73
oAn621AztJ0YlO3zQCw28phM3TIpQHsPJ4OSq8cmMFbX+8Zb0i/XHwhsiC5WyW1U
yNQOVDnklUsiZXW9dC6V6uqCinRn8P+FYYCj4/zedSVKU2b0FHMiStE59M2i0rmF
1aev+mMQ2B0TFNFHePctZT+InYSVv5z18rAhhLDDZ7zzcBanpdwEy8b5cTPsAbCu
+oovRNbDu/68RMOe1uj7HuXvmKqtyPMc1t/i1YaOR0clvwkaCQT5ObEINENT6PSB
X5c5K672VrBGSxVnXlNSp9Q5JHU/+y2s3s+8uYsvyQO7bIZ7fQlLm4AhIE5XBfYZ
C2qseHVrag35sIBDArtffaKLeZPMoBQsTv6HaraJXcgliczzIMdBHOkjyuhbmPBA
TzFlbXVDDkKA5uYuBuxUAPK3dHyoXjSZfJ3kVkWlCIYKsiwdRv1u8ZVv05aI1br9
n1nPIQGl7qkOf9F7udBPHc+kUP57ugSEf5KNNUmupVj2QtTyxi6mZqOpBeoeGISX
DoSqCtQ9zcGxm6ixdbdgMPCXY1l2UJ9WLbQMXAMlKFXGe4ZyVjeRFMjdiMMVEiWp
Gkl5/Vim14y5VKBU8sYi+tTJTAFgj14uagSOgy39MvYOmCH1r7xbOaeAIs0wBIr9
9DC3FRNq1lbRgoMYbZbzgfQRJaUeEonwdqXbc/ryHRY8IMZpUv2k7GvOp+Sytdfi
TtFuZ0+b0hDK0QzEfRPrd8LH7TeB5qWvfgQRXcChpolKCiRhXZoGr+XebOffiLCF
rYV0btDu4wMTWBdtE/RuC6MR3trxhj0Z/MvhYBBECj+I1HHQosAKPEgboNlJjq+T
P5iv3kegKYItKYr0BchV8F0oY3SA5pgzkNiFYgjeacfBg1WHQWWZAYYUXF1p9+QU
akc9VktQYUk0YlL8SiF00SAa+VRcGKfBvDKLQY8DmtoKfP34g7rw5ndZT/OK5qNd
bkx+jTO64GvW9+NT7k19eSYOYqqVeRKlJlmkhOAP5l2oIfvOslncS0QditbsCpIU
LJQyzVKxOkpSqjk4Uq2XJ6ymXr2F+ay7oRFkBGgnLvXY71vQfj4oiL/6hB10ciVW
rvfwLc4SLXCu1JYMuBPMT8ANGLcVw00NzYBje1yHGre3IbcPhcit+A3A+CMaU6tl
t2eKMcpB+0jp1f4bqudqoVKqEDZUDTDXMkvx0tvaaKwP3qXNQByyR9go474zD4cp
fYDlqcv0vpOiNZGiEBNe1aU0vq6Guj6eoAu3nBx4qzhPFmDybFPZNN2V4buoieAF
GoRxNArlPYgcLBLN6CAlt1zsmuKEA9OqMbkwuMkEEaLlJWwlEX4cSy6QpnDDNpUg
8yBO3wBaim/JYTJ38d/jt4VN7avNbJcrX2RzyazSnvyWuYJ9m4dU46n0tKCf/TKg
SEcRDiLKrNfRBy4i0qzs7ATATflu0ppKf8J/03xQaW4cwkVG43RgDxiXg35thUMf
jICLi5h+sJbelgl4NVMjSQQszV8E9PAVIKeYtlY5XM2kQbRZIXYkxeKST8X7NhHP
e6Ay7zaVQ5MVpFv6/7qdqFHlx/T4ohM0xaKg+8OzA0d44wOEwkDgBbEqc7HaBPPV
G3IZPumIeokDhMX3Gu4vKF/SP+tIkVfXm0CoUIohW234pL7aYTuDPOUAC7d9iKbr
g74+rOH6JzlqWVAUiiJaJ+/niZ7BUW6IMt7oREBOhfpq7ldgD7KsmMOO+EBLFXX1
YzYWVRfN5q9sDgjBahgvpfja52eLMZoCC1Onh6mtmE0CPYIAgt0kzw6ja5Ylsz8i
Z0eyWBpPmWxNoIJ24kqFc75MYfhMW2IequZ6OBTUIB9IQPAUXR/L1wCGW2d0VaS+
QcpNkLeFCaDQ2A3GyRW36jALf5KHkrzZz5nHT3yYJn9W79js1NlNkhg2YtCmeXx6
mFhaBxpSAc7quSL/BqEQC7PaE8h7t0dRyN1TaGROnjvdUOMUDFZt7R7zw7ErJSAb
8D2kGtMfII626/ByABQ/e1rQxUz+Kaby+eL0LcDkXOaL74iEg8b9IpPc6Bvn3Oy2
7O4wQd9OGrRomfxlJnzWG5tTSPRtxXmS3J7PROUZMK/IZKIKzv7muCQ11yEJDU2f
4DBC2w2G0vxu2vvbbtmmwSPDdoY3Z3fj6JKObzbzDvQmXRFq0MQ//SFLIPMjuZDu
IZFcoUoiUDo80w29TrGl8YQW4KSnj4GhMciXwmGtJFoGm7l2eWx6PgKhQEKejVzk
5lMBjSDlM0v1YKXBIbSdTT9iVn2d+UbGN1c8XHexfYR4QKsWOFvDlxm0K0yQw1dH
d71vEtrd+W44t0Travd7tpWLpWKnnDkyg6dckOonLXPDXPE5o0Rq4J8sWP0slnd1
7aTiTzH61w7jOOIiR+k5R7D6oYlrwyIp9ASzBpDAY7UsrV48nDczo4QijmF3IS/6
P8avFWAE0GHoDpFH1J7ET598XjwyqelBjm20Afa8BI71Q4U+8Y82jxfSJLIayMUq
iI7RBhNesgtu0A6VBtk8E+Lhxk9sjYBzHEFr2+uEL0DtpTNc5MNxPfxIMfyCwYS8
PHjGqFt9V646I5oCtBGGzQuAB37k+9KuCs71+JCUICEIlFmm3rNas2nfE5IIwlSL
N3nmWrPTTL0YgUgVNThoizl+AUxiSB4nnDZl7GWhaME+P8/so71E4uPpgCqy7AV3
mI1UVcDMR7z8HQ095LaY8vqND/b/sOOE8R+GeVFUXAMXkjiPmHZUiJvmwEHUtOnt
pK67OZH1VoCFGb7kml+NvY/rzy5wq3gG3Yy56FelRqUtlxiNzK2gWh5FosQbyXOR
Jctv98jJTaEySNC8FzaDwq37NAig3TMiSNz4NFisW32WzTaAl64OaygYX4DcHCGI
v8qvkpGRuAbCOuCJl72+j9pk+xLnYO+iawoTSPXjrTYtwB5eCmTCCJnyUSXBu5Uo
rqudxgCd/fYfY3F+Hp+rISeJv6Zu8kb7B8lBiTtOQxofKGNgmE3/MKxvd9bINGte
N1QiV4iCAUxOgTCyRYDny9yyJqRbrjIu0k17uUoyjxf1rEHuBJar6YLuJVTwq/MA
QaqCGYR6Udj4SkNJfkWBEmKu3nMfgHOnFeOGjBGdVzt202iajrxaRNe04MSCdPsQ
acyfdNoXhO5Z/EQLhOW2FqDJI7gehM1yLIXsxjrJysKw2kPOMgdITD5RnJUoSyaM
ejvu9WQawiRxTxkIOniaVNTmYzhBThTEXhbAYwSLsCdcBUvViMs8EsDiAJeWomaf
y/Ua0bnht4hO5W4Uy5eFx+NNg+tAh3+BmAF+t9G3A6FT4FYV/BDPHeJn9NWIX/Ma
gBe/YTSSHXzLKkys/7+rWe2vE5ZSoYsNPOwhszXszpJ8Tu/TocVRdbSqTIYb8AbG
esqjpw9//LLKRzWDiaYYRb7EqZxMYL79hfqhQIgdYCSAZfQNV2xNVeQBNo7aHGac
c7cRYCgZ+NMUV+/K4iz9hokIv2Xix5r84XlDBj2lQITPdjaSjng3XYhPVtW0YuRy
jyUzllesBKMmVJgUCkk5Io5VTGjhIBT5YMz9OjOj0Upysq80+BRoWK52MOnMkQAc
5gxx+SzuZGxTW0Qc1kxISUVbQh/xaG5GklFzXsYr/kQhGJVu6XO/pJASZ2nQewRg
GeJTzAjkmHBgj3M+/kts2Ag8yh/ioNzwew+PPfK5o+f+oIhwMelPMvFdHtJAu51l
6IYgYkUmFRafC7KHgCMu3t4gFu23SxmqpRR0N1ZDu0ehQefpmnC74kWJQKODmng2
eRqoClaNQVvBT8s0NDUIJnbgTOvc2LXSS50Wf8V4mlO6V2tHs16VCCPsyhZn00Rw
ovdwUdzOa6E4PQD33jfZyG24JQmV5I9ClTjp48ms8qT/eSZMVRDFHMyjLUGbcRTg
vDpwPfdAN3di48A3PpRBmgSDNcjwM9SF+oI0Jhyi3XjY6Pcl5cu49NnYyxxAlE7E
JWKfUVvzt6cwhuqcncYcfWHCa7JJuSj426XuGPjM2Dc/Q+J+2RRDTRHYcAVQsC4D
M4xvJjDntrHC0bfLWbR25JY+CfdDbc2HanwTO4h8DIPhMS2O+akohe/SlKwTfwQm
5u7k/ge40Q9G9bzOIk6jVA1oI13GqSkpteFiA6dj3SlI/wq3JfeOGNxSUTG4oycX
yd/WVboMX4SwhZzoIIwQS29wAFq6z2vGutvvg5jRFIaEqQNjXGfjirBZIUjE8H6h
VER84z0st9T8/Q0t/AVtWPjtVIGGPCrlvaR1IpbTYpO8G8nREWZfhxll5BIYI+ld
+dCS15goJn8Kp6QSGo10PMKId/F7GnB5BVosn4PZ9+TyqbqPZTLLNij+niMc/a0T
pF8zIIFZEsJrUAmFV2tnrZK7TNDqO+99QBhG82VVRfqrx8Ha4OejWSGnPvRdzN6h
5S3HGoghbiiheIrmc0z5GedIXkDCvrzmbrUn/pkX6NhUINGBD7eZTnv2yKIEAAxz
8PVRzrMrp+D3oTxsEwlJZGH2HbVf4jQCpaXvACo+BEwCtDUhDNrpnbo+7d/JvRQ2
08rxn9KjLB8xPD2AAufTlsLxr9XaINb72qUapENskjVYT58WtXwHjFGhmjvLAYkL
/SE5x6bBLtE6s+I+wFVnlT0MGyOew0uR1/MZ1m/nJYxI3KRiz2QDY5gtyX19eu80
Su3kTILdADCFBexR4N+RpZSsS3QdO/cmifA2Ekz0eu+w+GASaiI+6Ronkj9W6dBP
BwYiY9E7JLV9PQl5HzWcTvIhcqTCo667U+WJnaKtO4sr/KUvrQVj6iCkovjJB86H
rzfqfpIrIy6ehIc4P8zarFrnVM0Kxos0/cRNBBHA9Sx37IKKM5q6z3MATVGIukYv
7dBKMYK7QQuIx81A+8ndt+7Bpz/8SToerx6bBcIdcBwL7wxayibF0mYaK5jltfxF
e5F+88aIIMf4lecuXHrg++69NhWv7CsGYswHYj33QKX49xPsIqQ8+al5AU0HfolN
K9qmqd6dTCwvSx/KIfFwZ2h/hd5oI2wo1gwWiXUlRVKv6wRwI/Nf7qpjE7aeR8DJ
uhp1TZMvF2qVV9B5gcF/pfqpdR2XW9q923uoI34mQOSUZAOQ6PUDp4pE689aUdTs
5vVCykGfU3MQhAegQRutZ850qS0QVI8Jg9kPBhwpgF3JUZEEKVBTrzhSUiyXhc3m
H7QiPQTr+tZiQqqH5Mt1tEZNrmoln3euhYX9AZ1Sz7ispnCYnwT6ZTeHmfmqsMUC
CrTAjj1W+Nf222C8GNIToEC3F2BEqXC8jK2v848TA3dv84YnRdxb+0m/XDvMH2T9
72GuClnIP3VhEm69kcID8uaIsRG+kp3ftPXfAmqM13OvJdheFuQoVsWBybBgwe5I
jieioWHnVnA+GXYcEfmI3aNW7IFTfxBSsIzFEUXE5rBmzB9jzm7fIiVqAmW91SZr
+KZAlYvkt80DBRhzq/vk4h6hQmodfLuPCrx2geRGHCzYvhRu6LZTXuoT4J0ltDUu
HjpAcPhIkjpZHpgbZU9lNDNQN6hOKY0YgAsx0CBSXkleTbdB1naeSbFi5nFmx2rJ
gQN00fECUwSapf61w/SosxovksIGYt+ND6ixvhlKsE7ZS94jcwv4UCbUwcSmLDZj
94/Ko6s0Iz061MrZ+yFgk8xQFEAeloNUDjFTZCFuNu6wp3nHKPvRY3UOspejaMW6
gFwM6frjzJm06mdq0Pt/ytK8PfufkozIN6rI2Png2QFcYBoaaicF93OMm7Hmgjwi
GwKwxEfcXBLYlbg3O+y/7HjjlC3khN/mUcTH1+/3NfPI7kB2QLFCbi0THXyMfU8j
wAt80LOhNPQDcmXzAtTCAixfWVTDb5ul33Zz5pTVs4pBUu4wICCG2MgZS/pJRrSD
8O+B7Ehsr7TprFT4tXOOfsZhksn0p6epyhQc6ZzB2O3Cmv6XYaCzxmA7RZ0SuizY
FssOOHiYtD/u8yHdAmqw7+nJ99YOmhxEl8mXHBerL3kuJz8Xi34d/Rz11fDC6Otx
1s6JVmOJ6I82a9ksSBOjidmLEhz9gfsqwWKH+MtKi2Mqo4rul19BxvMpj3dcaJei
j9rLxekY2NfiSPX+/jOmRM918avLxvgJGTjnd9KCcBr+ob/BNsPZNFrm56XmCisv
lDGa28qTN7rbf5k3B+wOlapYSgur7QJnpy2mgt+nHfxQUvPXVjSmkMsA7HHf4VbI
4AWiTGgIdwSKeWWg6pQPesbTfPDS/V942+HRerRBSeMyLK8nljC14L8ZDXOaqkv2
9A+sJPO0MxGu7TqXWvgBO4n0aRHfezJhh4AyvdiLUEcQge1s9LocuuuP0t3LQZVt
5X8pJFt7E6Ly6LDxj0V7rUHAix422MMM6GGYUB1Oy5dx3PmoHrEC0f+7lbcWvjz5
+8vZFNEIAISCcnuUFD8E5/v8IUwk4RzPe4k23QsxcLBj/BA8ll9Tv0B4M+hki2dC
GxNGx18xmCCZn1+DPTLuSSTkhl2Aya9ufdM9l4y/qq77Bsy3K11VywzC1osgXz7j
1wtLkAj+5WwdYhG0hvWG1Bu6sAvFdgcxbujWw52B09A5FLrymsq9Zxz84I4H/Dna
hK+TmqKAmwSpWMpDw8iphwdcUGuOLwZTGVsV+kgT29u2QR/zHfIK/MZcvRxDH4pF
A6uZFsN1sUICi7zb58a0kERflAgeJM7mgJDR2YmWbVqvsaMmHZ+KftP2KZ6Wmrn5
6lkCKMveuWN7YIeJBwKZ4YFRkSXVsQRornrb2WFXn0R5JJPrnkvvYfGjARi3kWbr
S5AxiyC4jk21JlggQdLA2rlU17RVAXyB23hGcSRpJc9LEnUofesb034qdplYc+K2
v46fu3p0MDJ15FmpVuhj6bPU7O2wFjFbZugsjhE73FDa/WSV0mSfyPvpxoDCYVrN
YCjVS6sa8qil02MfYcMXtANUkCRmN8ZR2m0pKCfPIpyvs0wUGLPuK6kfTeK8BKbI
pxOpYbOdr0q49E78Nvyt50j4EubyUE64pUeihFt10YYNC20PUeOHmSJRpbkHoOr7
gk13E0xjdnrbHewZNGyzE9woinkGaWJ6kvXGtJOQBE57xnfw0jOrjKjMxFfxsi8I
D4gNsLNoBzud25rdqO0k70HR4PXGXm53knHZLb1StyVzAXYaUdoczlEmw7Y0wkNM
ryaByM4an9ryeK86fPz/CgROhedAF7yBxm4RyShLGfCMXvx5h9Ts1T1QC5NFzWCS
c0stQzQf5lLhAPbuYSM4XeDHnWuo1unINbxruU9MI6HnNgVhlEXM4WTDjnJCQmw0
iessN0KxE5ommFfYTU8/BSZmhAhg2xS8f6Svig19Lsv8ztvddpe26namlIlNbFy3
CXofOLozTz1/0PTolQkGg9uBrp0gSERI+MBnm8hBYOsM/gEDKjXa67IXlwpkr2tE
YEnXzrDpC4IVGlq7sd3k2KbmzoJuHId6A9IqYT8Q+nSr8a9iwRe1CXvVZcCRhfY8
nb10juGCCOcQbeCZ+unEREUNnWdGGcLoGqqiDAZM+JPjXpIMIfwVO+cVnKD43IFb
Vvu7ANI8dAn0MRQMuqqUVtL2xHih5dE7cD6wrO2tmQWCtKrs7FcK5SchVOio/jv3
hlSwXBo6fpRz6+6/Q1yTduUbIGflWmtGFoefm8H5CuUqq0BlH3iiK7G6MiTLcOtv
RA1zg7P2HFtEERYk8TKOUyoUsbRAfdcjGRJxmWphVC/2Lxt2WuKm3FFLr4PhdjUa
cMddiGZvuLmNqKIclVIAcNFOLLtzaq6HpKFhYanrjr1HOU78EULpq2Wpukty2zVX
ljdhplvGz+Fz/NrKqGer8Yv+VAhZINHRbECV0kaJU31YKIN+G8lXlaUCk8S8kaKV
pJo82bJMIu1wSPt/Q2nV2f8dgC+dvvvCLPMLXSy3ptxo3IspW6MdDs7vH9TE3lgg
4NfDxbd+2vh5TpCimjuBmPwDQe36AYfEUKsxoPkoCqACwIAOcHRksJ84TwakQAbB
YlFJE8jYT+90tj+eynSdtqQPi+DYewe2qxMJwPT+Q3TemLdDT3gWffzwNkB7ioUZ
BHw6WZUY3kR4yeJGr/1phS2UZtjUkJFVvF/Uk7IGA5hQr2a0DfDJdzEs8PhM/2FM
mgKrDUIluyFjICujK5i/dtuljjGIP4H0Km5K235uW8C+VHZnM+na01hT1IlwCTXP
8rPuyw/gTA0qK4ZRKuGLDqOGHmMuQuvLj/4VyzaMGTJBNQC8W44p6HRlpNIIENga
eMV+GzgGEIehbnO0YcCh7h0FGeKue9Qy+etaCAZbfnjSxXny29SHaZdHP/i+j6ca
H6ZIQ3v+zuAY3ylfX2QiUTDEQ+wo+FtqjXpjZbdnIv4o+si0BhY8v7hif7n+/VhM
HIGx75q81q3t73wx05pIy2cKpT9vvkClY/ZfdljM8jtJGUH7Z1j4XSjptnKiVcJE
uxc96oJeqL+6UsnMpTwo0xtd06ysAODMpkKjuenHHpQsVjOCcBdduD1frUzE3Gtk
tOqjSptR/o6FElNCtG80uclqgZczAj5kb12PpC4djOp1iUxr7jWSDqCNbsjdKWYv
ZLBOuIqppwFMCpRQP2Q0hMAOCswyHyPafdpfDNRAZ8RBm/cv77maiDchQwohwCGN
affufYgB9Kc/Wz/A5zSvSlv0i7BC4kT6Ou8hL65xjEuRZ5qpAUomKM0l/lzooGZw
rO9ZkSvYf6/hfjtF+cNUK+H9oIXKVUS5gzwZeFhljmZH5shP55zU6ZpoVIKkKkEV
DY5Zi4R7ot96AAqP4m+9eS9SjR95db7lmeHk/pMi560KGIHtJTNog0c4mvXbbGkY
LCfDW8YQbiBz4swkM/1ZL/+pHIUT3dmycGch33Ed/PasAvrSM5W2kTcfDA0zGLFE
GCDFKIbY9+ubUw3BlZmYREuUgPxrK5LP3G65bYJxoq/baqsHslQAs9H5oImEPIzp
HsohNQ7Nei1ErSQOjf/RyE6UhlPf38uhtgJC0lJ9bxyCW3irIQ4NEEsVY3sVmdtz
yYVFMki88lnhDXAJ9bgOzXOdLowNPGiqiC36Ad49yWJ9ufyizUIw/3WvW4Dmpr9u
Y5qIo5B2H3+N/VmvvsnNMo5DCu5MSlSapqzEHjugngeXtiEp3foVenQBthbsFrB9
2h2mvRCNnkGtgrTfuu6A0xznXKkVOtEBqRLMjwqVjpaK6agp2/mtpaoinuL/gMUA
EQeDbcUkIR4HD1tZQoi5C8f/PsnRAvRsEZcB/JGAnl4qpO5o40q+xlcGWUir4ge+
hLem8Mxl75D1J4c0FomMC5yY9X0RG2DPxyUxTdEpN8ISvo5DYDAEefHHIeLf14CD
5ZqMiBSq1dh96feLf8QfPLYiFgUES8V660Ds1pxomIr3DklOmwltD/BO9FKz8AYS
/Ee3CXUkyTS5dMjDS4Bu9UoSdAFs1TWEchUqb0GtcnHKSjv5XR1R38zE7NijzMTc
zILXtVx/+nXO948l9gMxr1Vmsybnpk2e7Xjj/z6oI31ragjhCsxg5tBq2NbFu9kB
VbaGI1vavSafq0NUvON/9gvNHDoE4GqjgEYhB9k2p7Z+8wV9kcNwJ7YHd7IW2SOE
jQsMNxStqWY5BPfH9XF0OdLNAqSQV/JmAhT+5gBEHSrFcszPtdtKr2tkcvWv1zmV
GbNEN+fxM50CmTXwJuotIoYvq1TUbFQP9TNP5UqO2NWAgGyPtsxy7fmP6ZzBK8MH
3CLshza6C5QqHwL9GBkQZQ6HpaTsUu6CRR4Mx6lIigIA1DyolA2kDwZKtK0CToOB
wr6lvXU3oP7GU0+EtIBS+DurVIeXbnivzJzq9KcprDGEo8lfkgWi+HlOayL4Bi6S
IUWeq7sE+kRZqSTSkyoWxj3cSNozE6w/Ew5Z0j/UUZH15r4r/unQit9cXOcEEDKQ
sUN3eifc3hkL5wKIj791mXWnNOkE5sUd0pw2A0VJnFC4ZjwGnRIPysjQDj1ahxk0
xf7fs7nTBLjf2WS6hrLUhvstWvzZQ833V/sFFHRNP65q16UPSKPwvO7rf8mhMOOn
7FVKLusUpcsENOERtl6rSR8fjCcIK8OQZCqdheUP3ubAxeQuC/w5seyYcjCNOyJp
V2KixQKBafQODtFcOmfhV5E1CHY7GYw8zgxzxdpsDbaUn2rNGkhdiHGnczbyPf+y
UJ9y8KJbSMjA1PlqbycP9m6r1cPT2E0z2DL4lX7BlE566RsF+ceD1SiqyvCsKNqG
4nm/SRg2Ze58uL3SUDZNdEbIM6jHaTxq/82pCtgv2cuvBw1au086sMTL3LTv/sq8
W993xQZf/anoytG4KTHKUj1bOFHWjMNnRZkMSYseBPl5CWWYLfXGMeF73lDrVLYS
Y+Sh2d17E4LwE8/aed97MoNO8eOMwyPLBAlbAYTy2RZucbHZQ6b15RWYha1sdAlU
rRiaTTp+G59TfQCjcfjg5cfxvgCwwSEvtfVbh77+gC93ggX7jorQa0hC4bzmPnT3
nj1cVt60Jigg/3ZRlypQvQTTs4146V5Q8ZCKvUChdp8gjT2ierjZi1DS/PM4ppYM
795x7wp1r7KXPxAOzGjR0UpAGeZE7CsBmdkNI+Ml8l/dBDnfcabj7f5asf0WORcL
KtQx+8vBnpyLxPa0OBAzwq8loSFAIxysNjoWwMnRk29+i7S5ta6lgc8pKJ6swh6L
7OBLlZRTtppb3nAApVu7r/QyL0l5B/4aNYZ8idx/FAb/rnM8ttFLjJ0gEHUXFoXE
qnYtc3mJKymiUn6lx1tNQuZHTJ+LbN35QvJMFPLsxPN9dTwjAdH4LpO5d/NJiA6L
99b2nPPJgdFlhZVMzcf4meCMx05l5r3ULMr02ZuRTW6I7ed4U1mHrijy8v2e6sso
fOyzBQRQpG8WNjdatd1EyLvSR6D9bKgV1KHLHAhEWhtbZOnhE2XT+y3MTbgz5bpS
pAAC+QyYi3v1WSkv8SPvi/oIUSas78Qe6u4fqLS2vrmnIoAVDAI2IpWO76xSvlpv
jnviH8068EaN0FbdHJNXKFqAX6lBY0kpu9cYZWeKBOEcNnLbF7l97g0Nr90qIMXe
MLHpTbN+Mh6Lj8LBTByImk/AYJYxiuPMW/fFhawiyQgIynKodopNkACRDt4CfUpG
gEVqJhDtvnH6mCWtXoDpggdX9vJ+R5Kq1JFEEK6ygNZ/G2nSvCSu62YM7opY3W4V
Umjefsp1Nv/cz8p1HV4hAZ5WyWPABPdTdiSK1eSSBVW3FG5LVjwu8TYaoBqS2b4/
Uvo4Fuu7RYrVPO3NH7oM1QXlCTnzsN7RjifG3z2hvQczygBftcdRH34YaNUVXsVf
piMOQHyUUtGnCfs1+wQNoHQrADAdd0mlSbaxkmz0jRitkH3z9TBCOXMgjqnDYJl/
Zpjo+VARqLJTxMXR/9ffY14OY2SDvbUMHjsZemYSwhSaNNDYIKsjJQxylxTS2ROa
WZcs0GqzSA5zA9dVE7wXG/Sy0mhciZLz0J38PgLGzKav5Ab7opTF9CvHYHSpWlnD
Q8dLSLZpsongfjHD+sjQ6X9STJ8VxvKoqMjJzAv5lrH/d6dmKW9b7lnOM5/Zic0o
OJ0feudz21GHwzM6Sr8yEKNLWigNySxcNActN9GEpKSpTw9FvyzxAiSSwdK/6YBH
kWX+2eT8vHrGafIlENSgq2pZUMCa5Z5v9w3EV7rQA23cerXNaVvWClOahdfa38PM
zCg93hG6XC+HNxNZB0S1EbNB2hCWfqmw/1cthcU4S8gwaGp1H4TSlH7DnU2ATRt4
5wySUclZjQAX4M/L0rJ64fP9ER7k4q1Rysw5A/mR0eoDYaowD2hmWV03mYVhY03g
73UJR8Q6kI61oD7JCB46TnPV3BhAnsUv+lQgFKaR/n4B0IpQ/o4vkkx28JtTLFjs
vdwsTOg93JbBxNAieayKa3TvKc2pRIy+SuqUn8j2X8GeEoptbLpd1qdXOCBls6MT
McoMMHjz5zVQGL8tNSEvOzOtQHa3Z75QaH6SC1FZB/6Krfdv3BxVtUPs7x1F2THV
tp1PGBw+Gf2k0ulVGUCPtzSZOOR7Qpd3UTGKMc5pmdruEsrBJNwrrrw7S8//sBAS
zsxwQapmHFofiWFE23jx9gNe/7pYdmJCd6se2cGmCmq9eUV6qQgn7Bne2oVGxdkm
pEi+/DUC5/jzPhI5z/2Tv19++sMwSv4ik/L3+gL26LYFWXGpOz2Bagt9n1bPNn8g
txzCVPeEp4/t9G5LXkJUvN8ieocJjeQXE7JqIDuCboHQfFvXm5tRTvmqSxHHHyUA
YXhhagvjy2EI4tFnzpuuZgw0+cvx9it1v2wbJ6+buKNnPi5V++GdnrtNPouMmUfE
a/Zke924sMw65e2DHv/747QGoalpWZ9OM+B4ByTIOME0EZnudSi8zItjQ0icDYoE
abLxn6A7GV8IIFJ3klby6iosKIeViV9wQsIxlLf9qE/D9rjYX4PI31PQnTKJyUMG
fiLNmx4P3e95wDG8oGenwu9csm1+FzXbNOSNvi8ZSO7e3OElr1dsBYs9s6eAbLVs
Y0JS6dS+eX0Tcttb2Wf1mkGNClAry8+3ZdCAjaqqw8GuFSFoE5rpYlOMkPlsVlb2
kUxifv8Pw6X4riPLouwE5rawYb9i1Ek7UpfwlC40VmadtVmoSQ6AoLuDRYRfkK+o
/lTjyGFUF5VMxhKK6Ew3MxppmzRr3HD8Rdr3tpGZY4o9A3Wy6et6SaVpqRkZL0rW
mtczD7LplN+ryQuOxI7Hkd8wgWP8OEv4PoUW9Hf9s3gpE3iScE6ny8JciZnoW/wD
ztZYIHN26mtNbPuS9+pQfFFNNMSfZpuFrAHJTg2+gEIddkyzOdIQ8RZeIIXYno34
645OVdOKs+tb5te85og3Ymp2V5b2CNc0YeA6WjQ/OcK0PW7KCwI9tpzwGr1216XC
ZVUlwDAE7N296xpFes6plmH5asLxMbiESwTqEI7TwPmlEzmxzkSzo3OCNQDLAYJS
ZouSYRZNI1U8zA33dad6YAIdJ4KXkwkr2wSmhXJARio63Es345CfvJqVBtYf16Ra
KC3RDHN9flRAQQBjHM028jXp4M/C3jyj4DYMwT8FQlLLgOOGqeoBcaLNcIik9ta6
An/SCFb/zBoclS3ptAAtAIDZrLw52TKXTHx8Ai4i5MMvo46r8762UeBOTibDoUXe
kLvGn4BpgfTeUr0vVj/YL/97yFew9SBenSrbAxsreE2H7R66M9u7Xvh6e5SXFyeN
VWB9dIrjtU2tu/P9u1M6qWCKG4auV9E1p75DgzjBmk+FXgCVgA3GXVmq3dcaMeW3
vpTy/4vd702MpXB3LE41mMUQiHKWaDkJ8Tf0IYEdGJ7k8PfIMbpcVrXOC9UocLuW
jRXardsKx7OALIw7TwfJD7UCATDx+zxNOqIRyKySCvRQHVFaFcNN57UJqDgtnfYo
E5JLoPoLo1oI7xWoUEjgFmnNBKpWBX0sxdzg2QqLTxL5Po5UBE1tANTIK4raI6Rk
ZSVWyvwu6BaZdCjaybPaVoPKBgPS/kKqXjqAukIVBN9ZiG553ujQXknIjMg8FZvp
jFZDM8HVgwcmw7UbHz3gHh5djdmnruQegsoHy9HuXjdQDcKQn4893TWDVQ4sxNAz
lrmLceLWMX7VOSjzcvN4aPY7sy/5zAjpb+7qVTZBLl0hZ4yvXZengyFSEIDyHcUd
XFbJEFFXVU6C1P08+NWw0fT3AT5+afO8uZCqzFEhuEnVjV8HdW4rXG0JpEcA9n4M
5TNeTBjAgOTkOcxEeI1jDkrwFgo1lHy5r1mEtpDAzOtv6gpr6PclIPEbTcAFHv5m
pjZPxA6AlLCodjJqagMFaM84j3vdYNmn0a1prqYG/GA+j2khGHbUN32gWKAZ65OM
daGaXKCQQ6NNx33BGChF1lIoHMjk6KuKtWXzWfV8KbQVyYNeoUSD4F6XWtaWf4lX
lonPVsoMJCP+I5nuXlTcUf1Od3z+cm6D7lWQRh8kVKFdmL77HWRUqZxUXkngLr6g
LrXyaV6tvrpfcPuIvgfiOPTdykq+tweWNeOpvevlqPsEmif/1OWWZISH7TbrvNYb
J3n7hSGEURK6onKtGVgFgLs/QTlp6gdUbeBy6Olm2neTBqOBN5/jno5a630D/+Kd
x9t8OYOhOcXOeUpl67bks0dOgkzCb99yFqylkd7BnNGu5PZT7xYLuK5UI297DYhj
S2CjbhIHInNlCD9o4Mavl+R/nVvxa1gq93ZC9zFBqJVRIsSm7Z0oNw+fJyUZ1NaI
hQtKY1/As/g60wkhEXPTfb50rwjM6L4VxnNfkdAFlHRM2B/Wu3NoCOvRqZLVIBo7
pqEknURizbypVRhJO3ra0GcxKflWEm7FTA3MYr1Qb+8wMfV3PuFe3EJJSjQMwnga
wu8Jlu6OZhZ/0jkjugrwXKoJhi9G9Mxx70ofPUPeF4+AUaV1QHTGXQrLhi4V5iQv
+TSi0NX9UX/Xux0ZjvFF+md7BTyXgInyTxeyhVvIr1MARUIgwsjE9NP4OKn5xb/G
y7578Zn2iWVF93Mvzj05X2PkgkR77KLOHuRtp34xJCOYX0sgoIizoxJwOHuLfKQv
o1rtzL/MufKoPCauZqMCcw6tNgdFvMpHVYEw1lGwgVat2thqK6R22M7jIiutzg0x
tuPOlejRnpzeOS/0rOJM8HBHj4YQu0ThUMkcjcMJn8ab+mJMfEuM1AcklmkTId91
XEBm4sQYpzwxSkqOBuZZjJRrlH/9TA2koi+iyIDPLpXZ7Vade1IEjrUI6ynfHI4s
f9q0h/dpf+tQ0aTlMJaTW4bZZep6lrOc7bmfYqUcVybbv/ncjCvN8AQwjcRAHTh3
JyAQgIaAPC+Mt8G8jg+BSSDAg7hxn9Cu53VDKPgK0LcOVKWttLamcCt1Fst8ekz1
NDcYovmXEenseXeE9HGxLWiIZ/NJqhA+QIV6qLrVdsYgYFxR5c4hP61X3mkJf0rL
5/kw5swQfx8vqKWsy8eb7RE8HqiMPhrAQxWG4saLJgEXWkyZxgYRMgB7uz3GM0nA
/n2OQIRQmrd8ZhwIRflG8Z8d2oXojLA6ODkpjmVj1YzaBAWki5vx0n/crcchHgKn
DMPQPHRssd1D3P1sKjHtdCrIDnLBhOC0Qs8+1xkXvYGKa70Hh5ExNH9RPVmvg4Ol
NfEcvp7OnGUqks9N4XzhPsEv3IwbCE5e/uz06Ey5fWTw/T55yjy9tWGSlEZ90yYC
g9v1vyAMgeCSC1nvKI7BVLAWG4m5tDM3h207dnduaaDA+zNDMoxg8JTq2HImrLqn
9eDkONf4kD48Vk0/6qtq792L3QiAWTeNGwa15ps06C/KjLjV0vGnabcM1jkWGNhj
E0ypHwTS2jNZlYyADaVtK6D/Ntd1WgQ8MFdw93ymqYCa1qAKT65aPyXihjsYQvCR
K8b+pQB/8IPcXlH+fkFvH84eAu/BTl8EcgVyrmXu9Pjm6B+Z2j+r6hkJNe3c+NPD
lI0Z+hfjQdfPy5tJiwPF/4+e5qtBnX+jq27LGTsf7Ysggh78c8xaP5FXaALwNyf3
yACFhKJE9oYlCiLSj55yS8OSVRQX5dKQRGsMrW6gq1RQPSi04i+157HrcnNbpdG3
PfUDKSsABRL06Om151s4AiMKNCmeIVryV/kzAQivbL9ZPMwbFlGNX0V6chFXjvYE
xok2NLjxO9hT9mKLw3pnp0D4+9Hidu8FjosoMQTJcuWN6Mk0XC6jiIGLtvPPOzr5
1SL25zv9gK2/qcM8EsXQ+gTIp7sR6Q4FOpQKulPltR//1yV3cXe0lX5l/MkS4YQe
rXbyHeFndOjQkw2lmumGnOT+u6eq7G/5v0pYixPQUmYm1Dq1+EcBCEdZ2ulb554z
/ydNGuHETTOZnJhsPvQYtgb4qRmS4m76R7eFcXfpeVt+YyzMPa7iHx42XaOM0adg
9J5KhWA8UfMCEOYEM6sDzfVJIsneAXK0FWzEdDPVcTt6MYpFMeiDJ5K6xJLPSE9/
2TXrb2qLug5Z0Fu5vmaBmZHFZBOlKSbWEbHSOy2IhBfky519ucxM4vWTixJy+tqA
JVyTtV9DCEw22JBU70f8r86sz+G+uPKGm85nCf4Q7OCdA8CUtroJadw3mzE8o3QI
YcgQlaH7+g3U3RQaZ0V+bG5EloqYQ9qDT9xZn79PPnVhHxAhaZ9+pJwYdlqvtoQN
GeHL2+S5V5XV5QLP2hDQsxiyVetBbjpzd4bLZfIEQM9cFH01XMq/pVZUaijjg5F9
jN2Zb4+kp515p0gRtZMxnDYcrQx+iGVJsi4qi0QZYmQCckJq0l/fAdYDZMWDhYLA
iWwhcJqXvAu2d6smQCek2Ky54zrShINpXKANxYpV3O9pQoC1ZHDKccqQaO7cECek
/kuzU2ZtuBj8Y2LAhd65hTdlp/2LV+9ph023cMXjn3XtIYHyBMm9rH6bSBkhVgyP
3U68zNnkf1snjg+fRRD4I/acPNnXH+6xX0+w2XY0S+sTLA6s1a5y9tFXu0fFh1B2
4hRdJtcaHNZqx+ZWV0vADMEwicfidc5fVL1TQKpMkvnDGSGachbsvNUu/edPx8UK
KXjp3U01IQZuyq71qKIYWt1ChJn70ap6LcPjCFIhp47s6OJ8VAIQbD9ltNABRI/y
UXK8pK8RvwIG2uliTYcpPL2/4fH6urWmYPNCJ2ElbZ0fvqrHHUVP5FnhXz32xtMq
BwPrI47RnyeEzpoB3pQ3c2tHhJgNAK6vWdJMwJX9CvrvGGtn0qGCj1LML8W+XBs4
ReubdTYJfKI4lTlcPZA/hC7+yYMQmxMVnA0h7t/iHxYgKi/UZj7VTcVH/0c3hq3t
tjRvFeDPTkxSHpaCW8CIwcfpV+TBpa1V7I0HqSTx0HySLkzD0xJDpruHK8KyNrzd
DGKT9oAZ4mwPhOLJ8Vw4SjEt2h2f1HIYL+q4PHoXKymvOygbp45VybsIVs3Q88kM
GnlDJXzAJ/SbaKeI24sugC1U/rhNtxVatwccQE3Ys73+o7+HmzwTfRNm8OCC4XKk
Q4727p+QVT95tVoVzuj4Mn89iliXXb/iZ0aLJbkF5uDXeoAyYnkPc0DkdF1skY4F
0FChyqGTfGRcTPxaCSqz1gHPhJcFB4v4cejo18eKqyb5fDstX66wFBmumPlWo2Sj
oPXzVAVkgFTELyRvf5wqwbqoA4hHQ2gByASgID9XxJ+e3Vik0ATna3JOKHUkFI3w
Ztojh/g10ajRPUxC6NgfZRa14JDFUKd/+/L7x0OkXptLq2PhxL5pRuPijlDTzxhs
TSZu5qdxpTsgjnPX83dhRZ6ahQcTHYYWtegz5fDJHQ7aELnay+c2aR2MQyieujRU
RgGlGUrSO3Fn1qRWYnj0h8LbmWoFxDitvIeSdHmXvm9P0NBGNpUXLcn+2m778d52
REPRTk3nULrAgkqLqXrjpS/gNlThDfasIyRudhFLg/KLL4Oq/3Duywz73WLfrj4R
+GL4Y8/RAXPD4lyNt+Poctho3LgGqM69XVFWSUnSHgbwOeSBntIqE2/grDxcYcD6
hvyWeacU/jOVp+mHmBP5dqEqb4tc1txp4WfOHczBxmNq14cjXB3T4eFMx4dJCl9m
JmQWz8ZS4rRu/FTsg2SmyTBvTiLpwdNjodwdHEwLFigF+qcvpG767+D4Otfswrps
3/WkHA3HayGyHYPXrBKL3i2cm6FtfrU2lDNE8mh7E7jzARSUboYsaLJv+G8+tMkc
aq+hhTst1VxpohlHjlCpLR2ey5XWAy/BK7uIz8lPg7PDRnQmRoUFrUEs/8KAuISh
HTFEUMf8RfrsMt1U7fdBayiSX81d2PIPSDIj7vnLHiOSWyK+sOxhIrR6JG/DDI9s
/uugZmZNNIoPDUW39TXE5Con/0GDRV99/qriCGkmkxW53DqDAnU0J5niMEM+YcSV
K7vppUOYASm9v2rOxPDECyIaWfcK2+MY+xNmL888DHCa2UwB5HoR7CK99QTPZS87
KUwpDmCcVLIWdujLiV1d40p7c+lHRILdXCYjxvDYwuEoN/TNWFAM0PXem+7u7wEz
lUuV4XRDNxrD+lHaRFdc58pbq9Qf7ViJtYKzlDhQCgHRT/m6k/CbdyRdVItNzMNX
DWLTqBHLYEYeBLRKFHXlYrnbTn4OB7J07twgeZzvNCXAkc1MNfGpQ/kEtLrW2oON
4RCWhzV98CKSpsD+aRFZ35qyS2VDvvoBCYoPxK/EsVt5ERglTYAkZT8Xr87M2llE
z5/tA8UIXGHIMzLrkkgAmz88rld8uDGmVEuUo06MG1Sc+HDrxrrkVn6ErCEUs8dn
ZE9ckECixSVklVP5OD9mXJeJbafnpeu+N90BKswsJXl2WKJHRC8VW6JMde+b0fh+
ocxiuATD/UwiqSrXqEs9XjPwQnDDqdi9t6ABaXynPGcOofdQdlePzkPmYDtA/Lpe
cqb1t9tiT/MBnHuHIPqdk3i8Jmqum6V8JgzUs327+4rGNtP5a+RN/bMkiNM9WiCl
BW1NqQIg62PzTKcj52C0WeDQQbeSkS+n1oqqrYYdiVDsRncZTripr2LRfbZ/m45j
OpyjkboN6xd6TlQ7hAPp/Lk8UsY9dj3WP9STernKxlvbRZBMI1w2tYFr+d87Um8v
dJ+ruyVp1mtb+c7pzDOgRe2x/gKW1Puw4hsrnXKrDZhZItWKgDgMo5SouXyUO3mY
HXeGSgvvBSuaMTqYV1OEoyVOC6f0uY8FOzn837O/mnj8iVQzmQ0ZtEKK+ldH3MtH
ZP3iEMnHUJ/ufHEDb/y9GsRYHvgGWNQtvctwNwb2ZK+mZJgBXHoyu50nny3472h9
fM2prqzao5ajYwPRErox5ZtzjpwBTvYiMcAUDTN7ijko99HIAvEVCDtrIf8Kr8Zy
iYv4Ih7ZshJQLywzEiVHuTAHDnggwv/IWhZoSvrz6lOQl1SU9xWNA57m3Sty9nwS
tiKmbDl3Ho00sAN2CX+nIZTLewz2Dz3MoFwqSqOP2TKUJwgGcO9ayTh8u+EpNqOd
EEXB3ZEE3tkKDTGAZHsvbxdknZ6RzMcZXpSDQgKeDhWGvJnHoqDgF5WZUBMxrNKe
+XnoV7cCCecbECm9XqFc8nXJoAhmrrBoXZ6quxOnkb4LcGmxbkeqrhykeDpbVnma
Bs2WAckoIM7EhfYGcX7tktuVsercryOg7XrfxTIZHwf72+UE37giR7s1Q9zsfnAX
kziAxj3URS8XSGpEuPl/0fey5ROSWYf6TH4mbcqA8XMKSqT2kiT/kY9/MIeczDk3
FwDelRQON4Fo005jDFitgV80u1r4qvL2vPow7AifyT9A10Z3K/LfvfuIS/GzQJbV
UBMEZoFTA1UHp8wLPEQGyrcWZGMUJY4ypwB8+LuEr4Vo8y1MdO9fTb3swQfHM6Lx
l34ZjXa4xrrJj8nxNWFj269h/NhDhwUyd24bn6qHmvnBOFaF7HFXisGQ4/gCy636
e3nN2uN74wIJ8BvsH54q1Q6ff/MwE3ftoLOgo5/6nlWmEHYZBx5sBTPiQnol85nn
5vr96fi8ottbTdf3SYqw/M9/sB4StAdsa332xM8mld7xHet4oApBd657VXdISEX1
fm9U/Xmh9bKFaQNMznw3cYMfMwv45edKkfZ42sWkIllmGQ0ory4LxTCWVeD1k4Je
zpJ+YASJE5ysF0HRcAkMoY5aluLKy5x7HYIFT3mqOqy6/aazx16BgNbKlmPBBq8Q
JfNzF/mngVGdniNksc8Lhp7lRBEmRaEo8jWH8pCqcbmYmGzRo3s+xuzszLMP1vWG
wzW7re3yltI1MIRswCBSUiaVlmF2rTyN3chJ/00FBpdZUO6cFWFeDLLxpndNEJJ2
3RiNABZfj+lF5zRuB8dNfKc3ZzY0K9W4RCV4pSHl7EJnC89P+40ESXFndD2gPXQ/
QmyPbFndBOyplQFRllw2ML5AYjUPjwVicniUhDxwAuNwxlVyawmDbMEbrKgTJ7Jq
10ZqONnaGF2ZoqzcjVLCvhikYDia6xRy5sl1xyV7EUu4TA+wImz8DgPj8iqDxEkK
NlLmT2RakAjCvicC1ijWIkus481ZyQaM7DF+ug99v/QROv+EEWhzC/P6VGzC2X/o
Bsjv/RnryRZjoEn46aJXa+Pz/2A2Y+c2I8YnCaWZVG4APv/ysNqWYt0Sb+G7xihY
CVCjJHCK2oTNyuEGgvoKKFalEr7xOnl2ReEm+Y5vk9vUlYgM5Y+E/uxMXNbBMK3z
9aGkeNG4G2yps+kbbOQrKcaUxGrdLhTmtmcCn8RRV0C+m0NSlVAmZOKwwapUXUNL
RZf3Hmmw85D4r7IOWRfvEKzqGrTxJqSza25DErcwHsAelbJWZI0ULRrSl/H/9yI4
GMXJVU5mROfyjWaIjPyBhZp8QFc151gK2fh9+txU0iy4QCflEUQnAkje9iKZNrMk
QJgR9tZw1kWx1QNIDPtFA7k254ZQKw9lN1XnpBkdKGcfv7Dar8U7aI2Dr54b4cup
BWvPrgaUYANVbi9gEBI8HiPuFYKGcnEfNu7zWb25wqs1GXr7e8prpTzT6dP4KzsN
s3W1U3qhdERoKk7sYuVq1L+ilKKvy8bnIpi7C0iI9KpeYoPMazFffv0CsdLQh6YC
m54wIsrpbusQY0c0HbzoFl4Dca82bkmeyUndRhy+Mb0gBbOKukvKVeAUy/za8fVH
0I162YjaefWCfEkZ9G2g3880q1KuqQ0KHg/77yl2egJ87k//i85D9uA8hqYEfjD0
kjo+fqpJRmNrXlLd2VkwRg/DaFiJ42yNjDY6iq+5kSwlR1QQv/avyc1q9BYPdXsr
lvkyYGsj4C4QpofmwRcdMBo0DFWqUidL5MQyDIiVYKrLFBl35gnAez0yRUbny7HK
OXs/pK8fMgzsQnRAhmesyN8YYifO7XEz2EAX7//pdV3DWIRKqUm0G0Cswm9Tvw67
9II+mMiTuLqMv6Bk0KMWxMb4f49O4Yyuu3sHkYwE1mKDE5lBhP7h9MGbKW7+GNDW
uSbX1aGe03808mlH0mcQwL/KQ3dHN+V6+MmykqHjp5IyqP2skPKn9xK2P9Rontui
QqrYlsbG4XDvDr1BBmM+bI3qOz13FTs5X7gH02dEgmBCnzHGKsfx+7pzRs4WOg62
mRKwDIZco0RbbPlG3V3TgMXQAEFRbK7wtX3q2XiTUOCRXRPucN4KE4YYwSii2cLJ
hkB7Sco1aQigpzPc5oN741JK3l4UwtDz38zKdLyvNtFMYsflr41udVMFh3fgiedx
SCGeKxJb6SPELdBYDZkafjiTXqXsrYQHpbwYJvcCgPQIkyp8NsDhbBuppv0vePmT
QSN2HzD6BJ5+ziIuvHUXaGWJIYS+hMJ/Fs/xV+VZdQon7BvTGxhL7mASfAKN8ecb
pwRrm7+XRLWfLJ3U7O85fDAAAMJCxI5txKs4WB3bd2+uJ8OGC4jz42RsmUuXOayj
Ka5xP3HBlq0HXuDoVl1Au3NP0RORzX3wcIiz5rKo7Ywwb8vWfru1tn9FDrag8ggo
SixOndgvRo1e9/54a0HSEbRhayCdf5ZLyRjcJ6VYWAc6FHnn1r/o/Xto5Zm/dI8C
wyHU3aYCv5JGL0ei5rnhwvm+vmzjhnvedC6VqF2MFXkgaR7d2S1xAkGbvq6F8UKB
C09uYyZByuk3FAK4ffux6+FgRNT5OFCihOOq51+mS9d8KcCKW8sW/XMWqQf/FMMY
MLfHzFJ1uKm4+zjP24fnh9uUY9YNU1DyqRLQFzV5+gtfCZn/mZ2FXDu/sjTvyQdK
HyqdQCfmhfErKomZyBKm0PWzEe96+4aw8DjlYHrcdDp8++wESnBj8LbG94oNwWaT
Ym8m2GPQso1eFWSx/H1sJR4jAuYAEoxq5HMJTR/5g4BbVk55izzmrxBkK4U5KW0X
2qZD2MRkfji3Oft/RIChNe2mHwCD1no8wWal3+KYCK1DPTLt/2EhWjPLvOjzfDpk
EfM4hlPIBx1HIrbCOdMCtwLXM4/i9hkssO4IsRkGTnC+B7f9hbLRypP269BWQP8s
6jzc2P+OxL4F2J8ZsrSxf1hbfeeYUajyAtdhYjoN4jK4iL8wajI7W439DESklpYB
mwGWPIM1D/7thtaZMnKL0dfXnJX9P8ip0ZBpUdJtMfV1g0NC0xc6HvCN2iZv+Eea
T27fjiTT2CnBijaterheK8OJqhUbGswRz9gLwaYN+qSubLx99DaAgqolvJY3h1jd
c1DcoRPu4GkIRB6j/KK0toB6rN49JlxLZFwcC7KBnAF48NJQysRIrCxg6QOzp2tF
vpTM43F+qFYqIKHjEcIX6Kwdlbrm+IyP/nqLu6TkGghlqNm3RXsJB8/sr6htzI9R
CIFz9G/HUqFPAqXhX3kLAB0zcPPZ4MX6kYU2foA+TD5NKCRBluUByKWVo1iHb+EJ
r99nMewlsGkiw/ygMof8+1IKSMvjbLtBrWaI1ysdBW3kSvbUrL3HW5VGfan14StD
8Uq5jwp4mQNkhkZ9E0ZkVEMcbjTxmPKNUfM6ZwggQi1982OeYoCIu38XfGzMKzG3
moAYblxpjXrd/4pjG9uSslIUlOamYtG9upCeIvzhKZdY1i9sG1ceNAYKytpcXnVy
GK/r1XhA41IE1V27h/k7szNZ16tEdukOW+jHawClIqLEkpwy43YijJAdpHimWxww
5YrAW3HpmEx42favn2BsM84zYqzuDOdRuKQdTEbnmANfD9KWYg7ZGFEHaMeuxRFw
d1RAOAPxWakJSUOFTM3LVWn45++D6FavmRlJ7IooIMt4RS4U/mUncoj8Gj8ntSfc
BMYlQaTkaigQqdNjqhOVWfIRlCe9kGsUeMHM0ySwuKkP2cazig/CuVI1Urkvc0dq
aAbtnKXBHcxbixWGEg+3IJk+kREXDBleEzO77pzVN8LXjFWBkLL2oD/C75U2XANx
MmUx7NjBDUldLY5/NRUFcuQT3EGeBeyJHSXPUGwWgV+/zR01XPJExEbMVoITukkI
WbW0jOBtf6uWjo1N76h/Alv5dVzptoKAruQQDz1SM+2btJxO8bHNfiEzNZlSYQYQ
82LYnWoXPab9t1aBe2kncyT7HsFSk/Kvbu0Tx2q4sOiZgL6Af8ygCvi/T0YFFRL9
UErp2e0eBSqS562Rtvl/aqnpSBX4Kx7NrK9ATPEY/KvRAbU8Qs3gt7/mYv5Nv+IJ
Tfw6O18C8Fw1AYuRn2Ireee1vVTuKn50B/yB3IG9zmOf6IuEnBRVoW6qwj1vAnp7
YrprfrPTvEQAVahbTHLfWgml3Pwugonmuywg4JYh0fWEa0+Qzkdkm4TUxlXehWQW
Vw3J9+H9kRwnervPBhd+ZPFyU8d3hXXyg0aS2sccQ6EBEgUiHwQaDXxieekb4fEH
UMgBfgLnv8J1m+TM/93Txw2cUr+FaJMqfG+ysKieoQR6IDFGLKXJgURqk2XyutIH
mnFOnhqYVwodpQD0tzspHLvb8BwhiSOMD2Gfnqo7/awejKyJ4q/2i2J8QpFHVLzd
Mp3y8m6AHkHyHfbbKc3Ygc2UqbgopExT2PtrY0ytwDGTEZoraRQxEMBzEXiUBtbC
65GqK1nECpnP/38DgYYW/38PyLz+RXKE/C1p/OCAcuKpM8NpZ8ZtHFhhflV/0K6H
+aXsWXQXdlsf8yltE78afyhXbnM0cuvVY0nNuQ0+qW66dPfquXRGmYx9kolFWsyb
6rwDWwqBeHBYLUz7jgWTYES2OumM5xa3//jS41dGTK5+bLjzfEL+v9iYncC5XszM
Zw0Tu1n5QmhGNYzFWFjbXBK1ZPoBmvNv0WuyN4K1M0a4ZOO3mWfyNRQId7mJ72p7
543elDRBrA38I1G96yVw4j1JuYGGK9EszTjATUQUHMDwhm4mf9tDuL717IKcJ4o7
Zpwghbo/pJ7z/AuSiXqD9fI7N0jDMTjGU97zDrwliOpfGUkkY3m/0Bvp949QKQUK
JFKUkq1Wi0GxdpZ+i+mQ8fImM9K3iSuKydlJuO8l4hmGIhNtT5EP20HMn1cgIWWq
5o9Q7oMmaJW0korsKCVd9VD5nh2gR6jf+pR5h4hiVYOigxp/hZyVMm/MWmZfhnkl
RfVhW5q3snhMYt98Q4ADEXR3qMyW28PAzi/P22MAxDQ2ySUXrWdJRfxPDdGKUv7p
/zd3Iy8FANhrOg7nTkROcdiUCrtAh7EMmkeFljkdt2a+mR2ngTYa28XWWGmYTuHU
g50EjfkX+/yY2WK+Dc5Rem5u0RcpXM3L0BdWXzyedRGFr+yzwgI/tA57iqLdrdtP
PPR1lieS9sYps+4CbSnL4X3nHaya7msyAc7C+dTzfQwLcMF/u+S+QTg5yBfbpsik
sCoke4zRBM1a5I0R/7CdJTHuozznBO0gYWI7sym3bgDOnd7OgY3ZbC78Xncs7AGA
5oHckdHH1BsobOsGhkqBu3/bTBMGRZkbY2MHCnqT0Y50v//8/dTapacjPmFnb6Pk
h/Hm3CdrobRYab2BXqFTk7PmapDTFwOgchNtIewHvxvXq9yorXjPaR6CoksEWrPL
j2k81aPt4p+jIMbk5smQMejh36j+20BkEEhRddl6RWj//WpVz7jcLd2HdSTid0Uj
KcHNJIX39Yad3ypyeGkM5yiGtbFLCEekBovLsg6KAKsJA2vMRd8Fbas2So7ogG2e
Nze2c/a5ovAOBBHoQWYaeyLr4JAjfoLWKJToksV99dqUWIgzZyseHGE4HLdAGoHz
8e2hyhWHmh54dmghrhbUiM0Q4aC49GQjR+mgHu5Cc4c43ANxeSVVan6qTY5/sRl5
rMDqV7AdgwYEfmBMa+DNDRh5HjH/3oYo1ttnOIgERHScni0qV4A6XB/G4BhoHfHx
hUqjiBiX/4gwOXJFxfPfTnnxvkGJSg+wF6e+81pAFoSHOI4S6vLrdJvPDNFUWUN1
ULTIfjHBsZQqaJFOpkSgd6tqGPbHGf0I86mcCNkDe65DD6nNzRhXwDPm7RAoUxjC
gp0XXaIumsOYzaiwGkMl9ehKhEE79G6cGdLRxRZHsJoo47XGnHQiTXLcRXuXNNTK
c3sDv4/FMd3tTBR/wzYyKovdqMuACA+324Seskk1lnNnvcbWgOUA06f04UTJDd0v
Ef8DJNwZWwWsniXqWy/PkmTK6rbDIlnJrcm0+GkHmiE9yVm69MLtzlr+pa39tSN3
vYXfdojBJGNhVlgIhlLHre1lJ7+/hiU0f/JCgHcRsJPxoaQJdIaqJ/JW56NsdlB3
pPV7KilVGcFfdlWb5Z77y6ZXndW6r/39jrWphJyIAr/fMRsuaKD40XkdM5j8i8ny
WrqN2rVjK/MbrXMrzjHIkvXc/t9KgITlAbgkmUhwPkGVFQQFP4R6bkyw88xDoJBD
W2h9XG615Am7XeCZV3kZhgeuSWrh4xpyIyO4d04POe78z9Gey1RBGK69fK0st7eN
lWbEfD96MLBwl6YXvV3DUk//RW47bLVpruNrBPntZRDN73iXWJVIA+HXf/znCOSi
+c49dCUp/AH+UYDQyY11WrTTtv4/3dj46W+Rnibeg722lIN6fAmoq21o0zp1aE6C
3/mEvhaXzCHxF3Le+WNDunGhw4miqBkMxxKi9V9uNxUurb+s6EtZaSsp0IzTkgdd
g/7hWrDpXeODlXdp7dnMQu+W7cTlBDzQ19HgnSNi7hQvPh/mrIIeTymZRW9I2dMf
LHm8b8U2H6+B7MFlInyQkBf34QDzodFN7DR1g4ELT63b1Et8Z+7QkkbB4Wxsd5dm
iPFsJ1Pp2Fu2IOq6rb23OvBod8yymkyGWIge0VmQqhbv3mu3k0wVVBFnfWdwQlun
eswAwlCDHzwucA+ms5G03WW/porsK9a/7p33XmkXxdtm/ewDi286dtzro0I7netm
I313duMNZsJ2kN4yLiyfGDVwVtj56Lu35qLq+2h6VA4p0sK8KhxJSw3jsxSEQeVi
NQaJoHsKbQkPz/LOvXU0W555Hk4NQjTupnnS6ljqZv0W/1Q9UMRJljpmkAHu0Bml
wihN4p0WBce4s8C5RomurSi75JuufJCInraUoRyZWc5sjXdvYGETKt1KTiB0kaGv
58xcJx2ABKxO/N2qMSyZTUeTdg4QeeS/4wrDZ0nSUPUe8bVtugpOrFJH0UK6QFgD
2f4Khmjig0dQOJESmtTFGxQrYEGCd18NCqxDQpjae3HVPX3kEGnRj15E99zbbwet
MPUnYpiOltHVW36sV1c53XjVzq+M5PnzQp9fPJm+LDJ5BIAMiUCvY/RbsiVb4jvg
lQqHEO34GAjX/BzdqBRzxv1mPj+qsZxCpgJEpfEUV/NkfERk1HNRO30WEE5M7YFq
4tl6lme82yY7KURl9hmOizfhXx4trP4di5iCj7xahWOfnIHwi10xSbB2z6KaZQIU
89UmDSU2hvzHIb7CC+GjuLFvu7JSjlsnP59T+SzDKxQJuJsGQQh+SYV098iQabDe
VO2cIF96Rzt0/VobzIov5wUCz2m/wMLyPH4CbWoiUgVftXGyvbgBxURwnZcIhgUh
CZc0fxOx7QInB/UKZrS1yTl2rfOUqSwlTraguAuOoYiraZndSMcre4SUJTtM1qsE
I8oBG7sWQr63B3Cup7ltEf2JDJOD2Y+nK7vbKw8byj+vfHBqPGyoWdjzuK5T+Zqh
DhOtvJPGsBua48QKxJfgTGfQon9tbhkZ1+XysFGGtH7p7Q25poNCrETFiLX1DQVd
2EhTiyCDtJOLUkBRhrgza9KL1rAompTwhzcMn9/jRnp0wruXlXB5AGAgiP1u9uGi
rc8uBb3c7bjLzuq1wcc9l1s+R+G2LfPNnWGEzLEZ1wlf/Yv41daUJ1fFZb1uvw6C
fhnUQsA8t/jis7DZlp0/CA5bBPGfwOUi1R4MB9CTXNo0d40Y7Uq5uARq5BnD/RD/
0MuHx4KZYmD7ossX7qnTnPk5h+85RKFYwzKGL7JR1Y2R5krTiU73+WigaZF+oMYz
4dIMYIN8ly0lXDO5cI1uIqXhTiYwR706IBbeMWvUCwpLXwVsG8rm7hI+axBx2qmY
tOgajkgbBGqplWitgXIZpRWwpiuprQ4RK1l3vra4bA2nt30MsLFyQ/9UrTq5KVBg
bg/GtRXhfr13j3dOJ+6+mAID851rI/Sdc85lQYDnnB8HkFGN6FKMRptlnwEjHAfH
l3mlKQ7FZetLoAqbaOaRl2AGGJWx1ru6YEtWeGwdfKu+MfTHe2pD3z4y3vSroJT+
zlncUP71lyx0a+WtPn4T3NwktrVwkKwroudaJYGjthxBT/sXFUhMAVoWgzQ1zVP5
YCaOHZ16rd56oO10Jjcg2B+Q62KqsbJGYQd0Pp5iT1wj1iH6fqi70M82Ht77GPlY
oNFm2WnJhqCUfLhv25fXapEOB4wgE6HBDBv2T6/U1PLxo2i88ni9r7Z2BV/mca2v
s+VoSyMi62VvUeHb8/HVFkrYiMya2vkbhkcFnFxMdSeFNquujddoqHzzsfw33GUe
c9jcTxFTw/yYwaid+9PTo7jDj7sho/3FLoYUOejUtkB7FYHWPihAOXAyPY5bETaP
kFy2eccY/knfvBC41psiNYJojYfsV5qnHdkYM/jYHoWWUoUO2OCoPgrgsEAxwHPs
rL2p7LxFGKGU92zNPjxXZ5/LIvEPq9SPwH4f6Je10sXTdrMnEY0dlxBffIEHpHOj
j3hvh5KeK21E2xTjn/qBL1Wr764TUuQNXFORRlVGawC+bFXHOxbngMZYHPgVkrei
QUCCS7T1hT7REDsHdOYR+ma0NTuzdEyvZcup6E2ASCqySKqU4RhsxrhkxcUaaRJJ
tExhiuDaBNNOie5A5XsHw5+v+ztUpxALYCELhQxDfRXjNArVJfCu60TjYVjkX1lt
EgFfO9mJg1YE1B+LUFKNpPGPz5frDtfL842oOi8kfikOb8PQIWQg46SK5AmfDP9K
IiE+3eTvpluKwc4RcIWfemrl6BejvCMzMF8Ct38E5ZjqpS1qxW2J3GKjdhZZggKV
1KEoZ6HN5a9HA2J9srM8l/zrnsuo0rhSa3mOhlliG8CKWE8LLXLGHFKW9wL65nVp
NPcFQla8do5A+d4YQElwdIkKNRYBYTxjGEx5jl54p8roXL6mFb9jscRuq9JZprhi
QzfriugqvqJgfjtQHwUCyNfbwcbvHUCCfsDj/tN0aoiJERMLKMu0r4avnCdtwxId
NYhUnGZDpU+UC5bipBdJEB0Yz+nMTpOXZTTY3/mdu4nxFARmgxbSjORhcnx+Nk2y
fV90+3TYuvYNJf7UoVwRPVVrkSJajZmYliHm5sbDJ2Ecg+j7abchsfvcH9f4lyEf
Qt0UtfQz6RgAsAaq0yETLfe7e3KbECsyv7xRPrBWM/YknT7LqDvIBjJF4y0LzShI
tCPGv4Xu7tTc/zYE9hwQFTEpjUxUlsn5Yp+2j2TcZ5F62877wucci2Ip41u5fTU5
qlrZ9UDOSLG3WyIupwbBDqAtaF6/ObOFLYes44JYm4r7DwL2fqUw5W7OsFNsdVjJ
rI36kLktpmw7Py/SvFCs/DFgVNcqjyaUS+KO4KkSr5jjwSLyth9wjJpXnMcfYZKJ
B+UlulznNXl2Kmzhwk836tN6KFrJyW1IP+cd/J9lsLt8WdKONYPub79uAurI1HUT
Kn7Pq70Ej6v5QDcFuY8lBKrwB3gPIl0tYIFV2xXF4VHq/59S/nJOGV9f5U1qaSwN
I0HMt3sonuHRP+iDfPa1IQRy0aM3WEHmQGi4Of+nsgXHjxwed2kI8NKw8gGSuBdE
LjEQyNyKFue0xGOBXxB8PtuSFufprlg/iVPB0aFO8F7FsBC5QscJRODHJh9CdJPK
9XkcYjlNYR8PyMCo92jrhcSIKgEHOZlxKxs2zc24rjRHNYPTzbD8jzpTB+kmnltl
Vx7kgh5dWAjqXxfov3OS2mz5kut5DmPkp71PwL1B/3QkDPljwPFCdxsohIX9Jt1y
rw1YzanK4cCpc+FcVfI8YLlJJWEuE01UfcSdjIsRKZbORzcyQKwnD0a3s/Njez2V
SPBS6dAMxTBJ+pF+ZQAW3Qwee/GMD/8HQWxF3owmSKIQvMg3JSIBGiQRXpjo9QIG
xCIMX8wI9mEJ21EImDXRiV3TkRBhBlN/nvoKUc8Zi1uFxa3zgmKT33ZE9Yywn+oK
epYEKjSfzuBlIxgus1Fg2p+vnyJFciatLtGWg9mWQn8Hg0whhhwApdTKj2yqpLgZ
dNfiuNZV4AsXZ1bF0ZIfkn8CX25j0IvkluFGlknnudrGqQnrhlGK0Ia/fNxp71U/
CocSDbfo+ZGgAhvEMv1+s+h2AUaRM0mRlQ+UKRHCnGFss5OpQTzaVHXy1aQ5F8lG
ENaouMa20VueA8AoQYB+hRhP0KhQuLtDHiGDWnaI7xXik8uyjiQHHgzgDM8j4k8n
pXTbzvSrcCfe4BBJ3K8hp3GC+Qq4x7PunLSUU6Eg7dC1MhurI/eor0Qj5Y16bg/d
hpvYO0X1mRhr/QuTQIVckPRDlZk4YF/8GpdIs5sFqWk3WH2nDgpaQPqpOsKwwVIy
DdNVBpxsyu5u2TazL+hNlePbl7XYIQOeQ0j7b5H0aZGK1vI9srgl1UYO2Wdajq5x
cPwYp3Gpv+0nOQH+Kci6RdFyK5NHLgvQM4ZySHRnVnK69inuXlechVNVUm4+0Gxn
1pdWmd3rkQTOr46rvBc3b3fPzslTdmyzxXD+7YdhjHuFutYvj/FpWEe9RnUQekXH
VSCfFdX/lZEotILcKp6/eb8w6V4XRl+TH+VbqGM84Xlh8ras9sk5PSI2VcBHR0ey
hLli1qkp9f6CNaJ25B4mtzEYRxF52w4Oo3YQqj4i1drCdGYU0RS4dqMjykqE5vvb
sRFIuLMzXOIX2vUsNPDfG6BgYoBHmr/Ynt2Xu5NdMBojCvj9nIvde1CS0TKh9Wnf
Ol406DaRTS8MEKk4JzhPSlEETUgO1DG5fylgX3nVPaY1WeAwCtyGL8PpAxq5uzke
scN8e8sPn+OK2qD+sZO6c385MePYOSyjgFqDGAFotaoK1iGp96nhTtU+sLNT0mpQ
Opp7iKfxTPeMgjUsnLSVIxJezyNruirQjsZzsLnZYk5f7il+1/lG85Hv8vqpsbfh
4ESMbo8y943Hy4TtbjW4/4EYdHXl+ea/LE2qMMMxkrK9RlV4qoegyws+7b6iZkkW
xvVFCJY7zPs48Fid8cOyWPoMlaTg5KvvxPAWxSNggC+lAzPoBYNpsEmULUZsU4LA
piRClujyISOV/iXUxpS5uvOvwAX5aS4H6xoXW++K6s5ZJOwDHAZbwNmjj3IuZMcp
yZc3AVGY0uhJFaJDh9d5TRB1nC/D9yXJTFKhR8lMglfF7vSO+JLlxzszPsq/YO6w
IDtpbRz7la/rFof5ID/cn3O/EVaFaP2trwgHjexeZkWFdPN95XbOE+arekkz7i7G
PdcXsOpnBbK5lK76ip2i3e2N/75dbJC6GgXz55KlHotOegAs41CpKol67wyIE8Ln
8Qetbz+aPkfCXPK/fhxbE/wdNFd8ZMBrG8WH1OQy14kuHXTfu0vmXAQY11Regi+x
4m0TTgJ1UkKTg9X2A5N0EcubfP9rMp0V75Z84E4l5QJ+Fi6JmmMRWYWv3R4wHlHW
/43BQ7LWVuZ215PkElEt7kuHIypihKml23aYMTobg21S1Bpv13zYoB1tc2oh+GnP
NE6hub9aR+GHLA6BzBwIFzce3jiSs6dpR8wP1FC13W6yD9VLkjAM/4rXQ7GKvKeR
KXIikxwMQDISRL3Ue7IJp8dnn2OiKY3oVThvOWjvyF5tAJsZlk2xgFF5tIQoCxR5
LrbeKjIonTfnmapyWfjcXv3C5pjl5mvsE/eTlVDWcfHNBGojRsHr1uZ8UfrBWxzv
r2P2FNMg4pm5S8BUSZIDyplYk38uP0cOZ8UKZgWa/xwn9aosNln78P79JS4HFuyl
L2W8xm4W4kakxmJDIOAqQVGH3fTt7RnrtJ4UE2v5ului64lJFzrrNzw/8+hvBb9E
yzs4uB4/OQA0D6JVgz05+PCLklfho+iXst9hibpULSqeC02GggQhcZOR1RrB0DOF
kgJgjCvfKji4oqFpUYY02cuROJmlyFJTdFJhjSvFZ7deOrL0uryxGMFclZYiFtWm
cNYy32w1lUPFZLBToCwofsz3oacBKyZtL8g9oRJ60ohixFZS8o3Ez6MMe8r1UKB3
lhm8/IGouKOTLRWkb0Tc5tc4qeD+6qvU3f6bLf1Ou/4zxi5Ho5QPrc5voHkEU94G
wbSjh76Pv1qXgjd7n+7XPus4QuT3qTbTMUHCkyItcKx0l04SpQYWRzdegm7wrw3v
rLsr4fLmwPZSUdbaekXhMvcIArj4QBoVCZNM7nw/SUyRUm1EDJlcwBpq3VoTZhm2
mQgPobvz9eohRNM9kAYrBpkn73LBHfplvO+iUg3Y9OtctLNcOPUK0eNjnBEX9iH0
2e9GJGb7VQGGb0wbqMwspjP82zjfXMqtMcZa1ivKKCm+UvK+/y389HKcR7y7PPTE
e3mFeVHO0cSdLfUeeRL3D6m9JrKvFTyJXoK5hPcKyYmYSezMsRhksNdw+/1TNHOQ
ocM3LTu4x9VPF+JO4DMIn+F+6m+CRr1xWa/wSs0xGdCqLx++4SwqZRG3dy/QyPqC
Xfyql/heSmj1zoRpbHzM2d3KaQYTPVwBsEFw+vfKYEZk3JOwqQBE0PRBxeHavmGS
ynq9TY8JfsTjY5qwsupqoXTTR40m9vf3zfk13ZbTREPMgQ/w84DqAS1H+csNPUQD
JIqnspDLVBuzuXD6ck3yR42Usttjo0TT8DN9MdlTXqWvVV0NyDkQLu7BqR3S5CG/
xrwXc1TiBBy2LpTLGVEACJ5JpEpjvd27W9mUBrJC0RXBVufLEqW2VvyTSepalHPk
FdahMeHNmAFAnhwDXrTCN4uMRxD+pSq7nYjFgtjhzw/HQ0hAMOhk+Zz1rbHZ4FKN
VjcJm3iX0DprV5bDNdbqlzSI52Jqdhn6bqeutBF8E7LtmO49rnBPcSZztoWZ16am
eqd1j/XToQtNdMF3B/b9gLXaPBvdAmWG8cnnZuYDkPpNN2Sq2CWJDLklCFresZvl
8lCPBMzL5O1zrtHTBDI19W/V+zjaHt9YKAsemSvRyWcaStj0NPJECV+rLCYwYXP9
eK/qK831cLecfxnkWBClWXbeKOT5Ec2XPKDrMgZmX5IyrfNFhbLaQoFoOxNIgPxm
3trrRX3RjiTKltuD9q8E7UnZJHTV7NAj5jlk6DZVDKod5ChKM/PRRktq9nZX1g8e
aY6O+TEfW+bg/mtIGhMCgqU41cSSpaZDoo0uySuNbfmxe0ohbKctukacjeO22LcL
UDu6QKFQIeFw+McC9D/mEUdvSd0e7EoIMGUmHqbc2jUAvLMXBJ+pFgh5LP686By9
HDcIojKcY6T3GN5azAOpakU1znALCob6pMuHc/BINRHqfoD8uVE5mHpNhmUfpi6i
Am6Z4vn46HVMA5VyrfJEQlbf5bkIFPH49Cfgc3yFqn/CuOgQdDlBHsjLB6h87sOy
0tuK22k9G5kgKBRkiwMXX30AxnBjSFHJ/7eQOaKdbqMcTheAwFy9MArbs1NScJTt
ZZJFU1ynl5O7vS8ickgxcPRCbUi57DU4KXvkAoNEmH95Uy5o9BJYtGKD08ZLLocl
jQPtEf8KUm0VyCRQWfVCKu2h1h9kXlv+altZC3xGbpPe9/JE4gBCbwaxPQHRMhIe
78B8YrWwthKMt1IsLj/GPll2kN1OizM27sNx1n9FTFqTTvHqGlRglcQX1IVlkRdr
1KqAFM8ztzcrlBppckgGG7pXUiqOHz+Dy+bGyBsdNLJTK8pliU4ZzkjfgokEk3v8
zo5cb3iPP7buztEff1AoKA+2n1CZH/C93DRl2Qowddfd0f2YH8gSiv7h+BEGTIzw
5HHPIQvbT351JFDZv2RIGZHF4uQjZCL584MJPK2KWt6XenhaWPzQGpscj6/HhKYA
zOtXAUAMwNK4aV3W53sE6/I9EqqPoe425YpzI+Y8QruZw4i5pMesVowqwubKxXP4
ymtxQpVoUbi+aaLNkpiYiiXiZSlzZycm5GGcMEca8qr9FO1kHSLSZaPYVJ60TBPu
c0zJgMoNRAcI+LSeowq2tajXVR2fmki+9165Hjp9AnDl9C4sNht4aM5/FHIXOgm2
7Dix9Tj1alIHJmHdsyAAXKGaleoxqDo6s4MOLE0c8PyD+u7jp+g6+8qxAf1fpbbp
Jm1izXO5+782kggftCeNY6bjecD9kmwQpMEkhzdY8iOKJ5AWQs+M8A6HUXfAahC3
zMt0QL07mldNyhbb7JHRQiMA+hzGdMMFguYC36QTmMbpQkT5pR0XTgBFfNgwkrD7
Ks7BbIPnNOpiTxVlMId6ZXoWFrRm7TRLq2OB0wK1f2GwCXBouR+kGufc2Ksq6Rog
rkeR7w5tp1/egyPomhhZWRd034/HpmEJfHfD15goTqfo1iLr7fBOy6dOdDkxE/dB
KxQrPUdbP1vGbJp1hFdnE547Wy8xU4VMhiRCJfGt20/PJKTjNwfgQwyHgGmJJcjH
TYF/PbdClr9f8U03gq7hf42ZB1V01zpA0SapLXoh7gUYSzsdVZHaGU2M+OeZ/cmZ
AQNPsxBEqGMqZDgwn12QfgJ009S3eeluw8mHM6OyPnyB6VWOZCZMZ/Nv500vQMbf
BeLf3lUAVALGMamsdiibqeP/2rTD/Odr4GoBwTV4v4A2qRXuZLuBv6MMdtAnXRws
re1iccclYioFuJ1ej2vCSW97OaZReNS+6SFV0sdeE8B86DK4t24f2e9YI8c60OG3
PrfeEGF1RhUl7XGQ4A76fggx/aBLLxImFbYVYRjJ6NmY1kgaVnSAgbkx0vIWEQuo
h0J4A1V4EMGFZqK9jsmFJ0f3fmj2tcpBDR9iBtoOnJbldXe1Tn8F0V3VSoIVWQnf
eG87rSalfYlv1Lk6jMzNRCyOtQR8ZaQiYhw6XTEP0VruPe55ykVY2zngOJk9h94S
seFBQvp38/fI6x/azzigZCl4P5ZxoYAVA2q7gjkkZzQovqPBIySCaJiwU7U+pCRp
pqac8PXtEuSlVnO6c7ENEVqGV8CAazjJ72UvC7ctUHXqp2nT6lgUU5m9069ltLMK
pPuHSVLieeOwtPVw34TVljzZF39UJvECZ7spYve2UABArcKT0yWAW2UPDuLN4umC
GHmyOLIUcMWjPTgdNTA1N+CgdJal694bzy/TxUjCN3J4hVPACesBsD8cDcvVGmtG
eexO1V4FcyZSYPqAMUanl8/PUn4EJXjxvYxumFe6Km4nPAgcMytYaboGDdULnmoM
3B4dpS5nJXLMHtOw5Hs8FdHqlMwy9R9MzM+VevM7vLd8WC5gaiW0iCjZ3VdJs+JZ
qjTUHlXe4b5HHwC2asznh7GlWIO7bUMrMUbyvWaARc6QkCNcD2ISHQQ3uTleRhgE
5PBSk9SYy/K8cvulIhHEh/NRz24v1vyOnxUovTgjdTJaHxXgULf3Gzn8vlrjXS7b
5fgkN7rVfLIJtfIfNpJxJDQmv34yQWKocpgYHHSJ2VXa5GJuWDpQUDpfEB1j/E7s
dVDCWM3LxbPyZOwuiSXVfE9Xiejr944Hz3MNHABI2KJ5RQkO+lUbjwJH6PD7AJ6C
fgGPC962vBPunkg+xZeQGcrBIL0VfEYipf29x5AUzks3oC11LS7hd3YH+kwrxEWS
ay3r+l6IZkuHBl2B1g3fEQ27Hz+4+5TdE7SuWfmHNuiJvLo9zZ62rySGo0rbnU8g
34CJmRioYH1zpO6iwS9j4wrvV/jD5QzPpXyQp+Tse+NCBQK34RoJAXgTjIT7n+ev
y4Lp+2i3LuXW0YCFpagNa4ZKAkKoFgbUOYbTQcB6IlVrWnUwfWBwf8aNUcQnap9o
YIoFJQV2V6dBmVG91dgjV70VNXBbqXrZQ4esQfoe3a/XG7bL6ILhA04yHWMxQxoI
IN2tb6jYLhYTV9xVUCOL2Bz7DXrnpIM/3wABIxpldiIk+D/iyFMw4m5bNJgsTOc9
QuyAlM32yBzH2mxt2e4HKttxfSI3heKliphm9xx22nF7QwnWlpI4G92n2UW4LrjM
Cg2CAgCIGOm3fUUptSdCkmEs+blwY+8rp+mnMV4a5xZ/Y4e6u78EUOeZk57+ov+G
2dFfg6IRmeM8ug/netj8SjCwiKfCANrzGwR64Xp5ocGLeE7YMh4LbNf4Q4nyAP9z
UnolhnfUJ/HxwIEStuDws9cHmp+M5y4+waX00lmjATZf6zffw4S9I2nHsGRlJmcs
YYnuM68myYQ6VLUzeB4tOJyrm8EEXTEUTM29pkUdG8pS8kKQ7qYfYltjr8Uy7TYw
dn7dWmBK4komWFs/A6O+SBAqZV9CZja/ffo7TNwGS5u0ipW2yGS0tUygspjpA9QN
nrs5gMmYPNARoLjP8oW1pizG3qfY2H7nSPTEGjbqfQGXcZpf6NkwLAF1oVtNB/88
0KYXtTiE08kDUB4O67SEg+zhcaw0fBB4xUyeABUpNTvvH43rcUBa2y9rBtbWzAgp
5zcVRD1N9D9JrNLf0joC41AelRUm3W2G49xV15yoA8KkpQTiWkzXpJhAGg9xMR/P
QhJOOxAR5IhVKkrmjuPjm7xM8mnEXtWJnc/2pYhrm2jJ8sSrOexBJXi0UOY6EYRA
oTgnAf+2+4RUIbYYPVYnXgZzsQ2jdcvGojRgkLralSM8nksQnIsctcEqqr/iQD6A
iB/74WVywnRREPR2v4zVG9XOBd1uyBjbbdMTJjcYpbnd8iQAJBE8Ar1DTxpf+XMO
AaWs2yLpg32q45KcKVk1I9DAc5g8mOL2TiMM/rPoxiR21o9xoknR0p8jUpLN9kOr
Z3C+oHWTAmX74EEzRy7i7Zl9wiQvcMaGGxcmiEUozZZR7lE2UCe1lbnAV5WMBb1g
jJ9JnjjPNuZ5+XmGaE67xKjUtbmi0u58si9X6Cr3BqNm2qBeWpubH9gJ6+e2BR6A
lVR9faUcPe8oUmZZJ2n8A6Fr21FkP5FSGONs8GjcfK3KZz+s3wWHdL6Xm7pZh9hP
ZL8r6a/OenGz2Pwha8LCuLDlIkyNJhnRGnLXGuYfSvgOgfv3QtMgauxnC56bZOwV
QbdcQvsPrc6nknLZVaVVTfY85EThojgwrQWNWyxjqOTiB7bE14XUYmYAjqs7R4j9
pcsck0sciCIHOSy/7vu+0y5+EfoNMssmyJM9C0uRLV47Ifq+MQ30inFp/cDJSKP9
OnHz56daapeleJwcMP/GJ69oIui7ChalKUBt0lfjdoQW8WhRtxYECagxV9VDnJK+
c8Zm2DD1FGQEc632wOvPN/RZANGwKrtJZR9Pe5YgJaC46LcMP5hqccfGYxR8yQGL
aH4dDKCDHVMYcbY4vkdeOoYllqPX+NUDjjspxxZ8qxW0z4kPg5mTA8UJk0tLoB0B
W6UO/v+UNzvYsPF1bUfbytfMEgvi1XDMYz6BL4F1sQkTat3/VQfokVwzhh0B6UtM
aK9PQ4/2kY+UKgn8i74YBAQELChjr/F7bL+EBE26kAqKVwCyJ3E0NuPG9W7VEdE8
5kIFBR/MfAF9YDqff2xcpH3hHb1kXQmCbicxUNoPFV3Ybz8zzCJsIDPsUPQpEWBJ
jHJyb8FJISrkg3VQhLYaKaSBPMiL7/7SYfZ3uBoa6i0dXQb/WlC5cKKNxiDrhoIe
O5gSlOdEaOwLRJswvVi7XWXV7y0aCiG37b7BDI/K6q+rUAYokBtYcPj5tUsm6sxa
93hXLbS6jcy4pj79d+5nXM+K0WruCGIYPzeM1arOzPQbD96gj6CtOEm9TFQ1yz/F
YfYoCWApvRh7fHexzYa4yZjPf/xx4geBcbJDZcN3N9DGCJuiBOYhyzrK26aQCVA9
LnOIEPnMjtkbsf5/nX2idYcUS2PgmgqelMBnMTLjvcWhMeCM93hQ75cySNbtRPHH
8SytOnu0Ulazp/eAnPBikfRz/xCkgmSgN/RFpw/rSE+E/DoN3ApwoVzL4udbTUYl
a1gxchOvU54uNrwHYky33PjTppG6ZIfnXXDHDW/QvTHB8KFE0CIAa61DabN6yhpf
9IaohtNvIgJ5/juf4Nbw/BfErAPDIajxRxAupFt7ixobIBazThvluOMljKf9iGQM
Mdryr7lYlNuIrl2NQ/6qQfy8sfzL/NSzYg/LOFJiVDNy5eKZNu+E6miN4L+0QzpY
UkU9W7WOYgYK0gptBAB7fjLOG9Fw2GUiDjhxXcXI5fcjvrVkfrgAiCnpRxZlA6m7
Em8DelwMzb0GRfPPTgtrd60o2kwNADzjfzZc28CoADTsFEP4fH7wwUSI2h5pLFUM
/vy34NzdaHhIiSvRHWaeoLBsJRYERca6OlV60RCZ2XyxxEYUP47/FGm0evmDMNau
StPgbRDawdt5QxrJcmmOpuZzNXYbjSdqkGjGGLBK+F7iOjl4IFnrvTc304OrIDZZ
sVCjVXMRqJzuHT3rFQdyTu3t/n+yU7NFFQsrG1FE1P//E/U1yKyAZjr8lP3pzIyX
fFLJsxPKsO7uSYkXlyfRN8HVj9CH5aHde8J0+8EmhnzoJbWfycwj7JUMmzEkjxO4
CcjjPXAWOcMAzxLcuJ9Mfs4w+OHDkQ4x3G1Ss0PTlBuyT2/3iHtb2ERbdFl2biju
DBAMCS3Y/Gt9EaChYLIdtQFgXoYNb90mtfu8RlmsQLa2VHFSh8uD9202mBoe2+dC
0uln7Xxnw0dn1zcZsTgtH0J1FLoSOYD5JJdXnfHcnIaRWcBL9nNVkn1XfkjmFyK2
SaIKCxrUYosSCdb+pNt9WqkFa3T85gKPoh0h+cOw7Osr91nc8XC4sqdXLH+8qr8z
EFpZftzeOThEuo32xGOo4jvQ7hhrShxgEQNPvIv16V7jJx9Ew28qENIzcoWlQsZH
azaSPWEyFJejUNerzvBIxiU+mdkAT/7C6mQwLQ5l2l+/AOHYxwMRAyio5wY+GreM
M31SgZ5+6dtD5NsevyrZgUUQpK6E5YRvlrkty3jlY/i5xgHK/3VXkATxrWjSAtVF
pVo9DetcqGzsxzAKr/6FRBESQfMES/HZh5v+1RPWjFunBCK0XUeRUHFzk1axFVKA
HrDIwbWroQniI2WcvcQVHjSRmQMoH9+nk63yXc/3hgG0zxJ1yUz8dhPLTEABX2FG
kd/ltDbPvCTXj7hqDubJmetsHaQDfB9To2XKAUT7fHwuyhVC2zUhWUKXlsQdnDbc
lvo4ibMfiX7dawSnmalYFl42fjt0CtGZem1dpagYoBxe/7/6KmLt19Qof2dfl5+7
M3VtFzrRgfIOyZ2XbK4TmSyO0lqRobBUAfP/Q9EShjj83ONSZZR1CqR151mSq3hZ
ZonkbWoDgWqFRu4wd2zYNZ1KbgrGSpxRqJbSgMIGA5fggbZcp84M6TBdRU0tTLta
L4yS6HNB0ayNA/wTIEJpvRjTHXTxPsGoLLWsSzFH84IRjPBfNiMhNfZgzUkk70GB
RF/5w7E1pjLIpA0qUQ1t1OTRgL1wVnBU68JGEYTn11UnvXMqT/oDBqQu4C/eFntG
Mbq1odcbCw8Oll///Se/5QRDJQQBPklqhJrs0BY9+iTyGVvkkWQhRPJfpJkRUql1
NBBuzEaUTBsTcIaJWFjKLByQV9+AXGt3Clqy/iq1QkJH5fp9qFvHpAZUrqdJiNAa
Fbsy+wIYi6rlF1e6sRS6F9ZSb5vJK+WP4OCbVlY6aiWEg+D2m0+jYB7JWtv/l7yV
L6wgCiYoG382fp5C0pfC+rJcrYtBaPUMxpa9wdf199XUv6T/ELFTvrqPfQ2xpByG
io/Bf9x3q2rAzwumicduqDBENVeCJFp3rasvv7XGAwBKlV0T7xZpII3O/VOXFBhQ
p8t75DLUS6rrDmdofdXaZq9cze4u5CnyzHAE38bXPQMWwQDdQwHtq4gDnWasxoy6
5GQTPTW4iNSDlGf5BIggIRzV8BoBxZnCs6LDJ3mRCCzKRThVx+0tZvRfp+lOmW7t
aG6fZ3Lo8oWYjekdOywC/rBPWYUTMpKnFt8Mh6NzQg9CxOsFDaVmSwlKPO5Lfb36
GnOJ34NwSAyWZSe45xTzrOic7+wGTXF5k/gaVFWApl5+rE0V2k0jWa5LJN6nfHbD
3EEaqGFALMt0QmCstokw89/JU2uSeJ0DTKuNRMfafEegJ6in83ZMxMblUmmnX0q9
Wcwuor2hUuZvlfObcMBIyH7oIfqwXdQ8l7WV3Crs5/Gmb0v63BQOJWBfsxtznpMQ
NvnX2318dICvPVGEUH3eFsJ05ykFHlCgbKqgx6X0vNpbiVPFR5U5SUcY9m0d5Qtl
8KxH7Z8a+PL1+apRBEaQvYq/qzV6IVsk0YyHPNF0PH3DV5A5hJxFmV0wUe96Hz+s
HOPmDAwGWLwknNqwsPW8uBSQ9ur/vxCL4epm48B5vtSqGO7j4XTaHa1YalT69r1G
0IXKOfXA5YYtpfhkoPgLNyYihblOSxk/fa5cvbBlBgkb1RSDTenYxaoBg3lM2oyR
ieaNWx0k5qrFcQimT/RQgG3qzxLq5qmRfmnKJszzlMG6T1fznOMZmKyr9escKxZE
QJrbeSJw1qqpEl++xU5C5wRswYLlZwtLzv/xDzlc00ZFwu3K6+5uMuFxsvyxCjY4
E3ce1WWC3QB8Y1nEviqXynUBrTFDC6PH1GL7rPH6odu/07bS8mj17PKhrpmspR8i
k5Y2hFN3F9gz37p9fXKtl40qL38ag6aGz80TCg/01grZ2gWPolUSLcowmdcIpTbx
6h6Vjp/xj5DguwAzciW8hQoL3/5OKBQ+Eba1gIN8YPtfgJKbzSiPoVaUPJ19CmCQ
SPTm9Pq/3YtX0cyIosUIHRuKwbyFgNeQ4SyyJnL7jW7QahyGzmS001+t9zhJ79tH
A3GtGkiMsAQvP0x/TTFaveDXgkQp/tBtYVWylV0970T1XvxwT9qyjKWmdMKXHPJt
pB3PlijRa7YfUVMJIpp6IA3QQdeiTsL5ysH0wxsys4ECRVAIvl3KK62YWZdsyclX
o3TeytcY88RV9jvYSRcolm5wVtXmelcx8KvDyXxNEHrdkMG5FOn6aeVfw56OQCA2
a8TaWQ8wOCHaDCqIx473MtkkQIB2GrM33STnUcRlMxNr+4JDH6vWI5K40tGlto6w
fiReHnFOwMRG6vHVOX85o2GNSN5bQ9XF3fHLL2Nva/V78O1drbh5lR7nfTnh69fP
kuEZPVUi5scffmOahKZs8H+o5IOe1jW275W1zPYmgmpJCUcXphUQnc9f5vsTb6Vl
16bzoBRq10nYmMoJRr0kBWWWSCbSqR8f56ZDNjAq9yXr3SpidLEMU1JT1vtNB3W2
ljD0YsUACrQhIiSDRbCJ+t2g7Qy3u6hJPHB8WyGWA398TEsvpRXK8/TMIK85hgqG
eEps/ITFAsJXY7m43pjm48suD422o9DW/O5YnPpMYJ3SJYWX70yFW9J+cMntflEp
pftsC5c1zUAwCo5CYcqmAhhIQEc/szIdXtW3IU8wYGIXxY5kD9wmsZMHc2VoWys7
duRWIf/92v54HvFrrdmAp+2u8GzqEQRKs6MwMPLi9WUGezHgsjCqNlW6eN+JhOMp
/XoWeXabpfqPpt6Vz66qr0ZocMnVhhaVt6Gsg4LbO3qwa4fnLZSPj5pM6og5jzar
dOLRugL2e7dWAomvhAAFXdvjS1WudQRO1XQpvqh+thowIeXD8Kokyrq4r0RzYMY6
Xcn2jiUXRuD0WTiqEnDvKQ8nNWmplysHln4+EIteLs+vgFv2qK1/JKphla7Gx/Ei
reiQ5bHQj/g9GenHqHHW0FctwlWnnAoQfdF8G0FuYjOX/YVqrYrACZJO25yCcseG
qIbLIOwM8YV7Cpchog1bsLXfygrZS6Cz6umVhratbnIBJ4AxU5OJh0CszsyR6d5N
2/YL473T2J+6DYFU2aEUo2c2xSjJa0ELkvpKDrna00bxFjokjH1sDNzE3/E70O5x
arIxORon0ghVu6fd4Ukq7fwN2vltbUOyyA9MyRd4D0fItx2fe1YlglljpiE9e5ow
vo7JAok0i7uW2c5jUriN+EMBk3sZrBQGy4hCPtymKvRk8ZFPhJGLyWClKSgC4xKc
QT9OR8n7J1j/YYz+cssxNPVDj1lnSs8iW+A2hmmNmJOhGNd5uNe1qxiU8z3FmdUp
J56/Wro6Ty4cJZo20XiwN3VpV3O6noeIXVmXs+0RsLR1dJJhZhUzJZwm6jWuzJqP
57xNVdJpyon/tdHPX1aS0Hgp736QwJB9UQk3vB+WEWUGFTJ3MO4luEVgdnhMKF/H
NTezRPWZRtvO52DE9ulDE/RIdKu6ILYa+RcQ5v3GqsLBswYAcTLKzAZ6fRCvpWbG
mbhWZwcyZ92ux4uPB8qfYS3Kkvabx5QnsPik3rriwqsHsfo1sVpZ0YkVj6/IGnhL
H/xmYbH7YDLzt3VZDz8E5tutcN3pLa5NTC6w3Ismw/yKmWAIaE0NXCj/y0ISseb6
8S1p3gQ5uGBoPtNvMDfzF/4KsCYwxmlewwB2qu6TJ3o+ABqZGGyIH+AO2FSjcEOw
1duY8C9EyL7xoCD87TOJ5VCSz/WVA7wkB8wV4oXBlBaf/TzEYfxRIHBuHwXQ5yi+
SnI0U6VqcCQRQoiJ8CjDJy1zNkffSvm6f4eL+l03ppZLxAuxsvjscowY7vZUA0s8
Ai1KIcWSCSKgoS4Vl8wBWrt/O2RSQ7GABBLWCnq8d3+xk8/PsFZ3w78hawxRXpIM
B6JybW2ZAZMnRqM+pR1OZVouMFQaqxcMWaEOFSMPLmDFNOA28Jg8fmew5/lq03fG
PkHWiROtX+4cn4EMGM2x6dSkUhb/aJDbf6B4rbjhFQG5fwmNtBQtEadGW2zbCeJR
CaS3PUTbFiNKBlc5Svw5RVswA180go1l885VNJYdSV4shJW6ZToyGUT57uZz8Kj8
Ov/AGk7Viaqsev0VH7oJPtmx9nikOsZtwtfRFxOFRcFsooA2UhGjFI5xbo/gc1g7
92f+iFOf3ofilRRlCc5ZUPS633Zf03Ubvwn3+/NTTu/d6VBRvd6nlZi/1tsxw5j9
Ms2MLZyj3eSKH28Aeo1IOqK7xomv2BD7zbVOFTobtszFumyr+M6noVqlP1kfXIDM
WQZ77E1fHnslSKq9l4e7jg==
`pragma protect end_protected
  
`pragma protect begin_protected  
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
oDDCJbgwNhMeupcXD4W5IlvPWn/ww1bhIBCeSjom+ihwDzjKasWtACaAo48hzFSA
SZ+zojMx7rldp1oJaLN8/uj/pDionB5/+tlFRNScH7hfsLVudbcNptgaqLNVscDQ
a1gUrFDtgfD/IC4uonVuQEgIl6X79EtaljqgBjsHXks=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 96770     )
I11wjjmEC++ErzT1fPmA3p1JW8BN8e+PPdOaaX81FyV7QDQOnF3wJfdcMM7fSqcf
afLbWcRXuz04mHkB/CvvtpmNV0lKDvQvWpc+xoysQA4KcXdDNqySnwgFD51PtiSI
vgXQu4d4CJU+miVzsI6+LPdW1llOEadPs8+E10kr+dlib4RV4UDnN5T1AFiAYuXl
48kaGczOroDHBHD16CwJug==
`pragma protect end_protected
// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
TY2EMLzrnKSRk3UQwJ8dmglDyA90487UYPLER9ndnr7ZfLN5nlevlXJ8AeL4lv6y
UXUx90Dz22zVLorCOHn21dNJfUWTswJ6pgOQ1zlAI0i77OC9Moz0HNGiCXtUMtsr
FNl63Jf5WCnUjLwEtA0DLprKhfjkYHbPTTHSdyEttFY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 97016     )
jroSdR9HTqOcOmhfTVEZWKcBDevNgSrS23ceS29LgTxaBPaKmIaua5KXS0nRK1cJ
P5Xj1C4pOPPS11JJQICH73B/Sy7PUAyE3HTWDtYKJIah3ZW3HwtEbEwc4i6SViu5
WRpI+RqQHaPOJ+iqr+5KXsU27Ddk/+mVeDqGO54uYLxmt1RD7vT6Sg0+VzrtCbwo
RqSaK978mHEwd9gjUZd3uPtOIx+ZgjOKeY2dCSv76G3Ia2AsqW2/lIxRMo1N3WgE
5er2JLhUGDUmB2zKIKF8WvR/l03W2OODJqh18yqfEY5qHq8/pe2iwCl0XX38ZS5k
dJhwaPQLx7pyoE7pynIj4w==
`pragma protect end_protected  
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ec5y8blLk/7Sm9H83dlVC/jNlM93dZpf8+Wq4j++uerYa2qZSFZehep07FYZp87K
YfRc+6ALhi6MDVPwtjlZQ2g3w/mWQ4MhkDypuIKVIMtV8tbbB0zivCTbtTR+bDrH
QDVpODD4V6WZwnx0wL5feWqAicjAudV1vkzhhPedgRI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 97223     )
FYvpTTlo2n5EEmVLoOft80yII95Lu6r9dmi46PcPfyHkIJXPiKzEHhez+Hgzgd6R
TMMGd5Gh5aYcTCVawk1wOXwQZgabGOrmZilIGPuCcwDfMV5ZfBGOnYbR9Z2YqQ8G
DXSBUgfdJfPwcLuinuIHzHKfS50PYmJtCZW+5yOA2v2RP4rK88YDwaDZjC1B64/U
10zc1QoayAIGgv+1rDc9zXMTreBPzDEYArLx8WicFBasSk3l0Ce3pqMiSUoZvbiE
QVmupjSCXP4Xn9KHSquJfQ==
`pragma protect end_protected  
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
I83X94Em/tm+yVVbjDnnVz1pNgURPzs/Bs5n8D3T+nGJpj7/GVLC14YaDKI1gXkt
21pH6M4m+6FY2j+in2ptSzRYfA944qvA5PHjCG/4+oUyVFkoEwOxlkZNHdbrWIBm
EO0mze47c035bMcYobhPwex9F3xsc9Ge6P4UtEB+eVg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 101281    )
4wqJLFTuSiJzcSr7GcnkdHLmsG5mbm16NtlIOzoh/T76u3SvU5/lRI1IQsGvlIh0
CKVjmKgxHsQij8DATRVKh4e8bl8R0I4UWCcuKgN48Q0/i4naJP7+hp/t/XgL4g8r
xjGGw0cBgPKcjzMii5BbfT7PmFt4u/J7C61qWfI3Yrn+sB62tr9nTHgCyrLXBgwz
xMMi1GIZM+XIUFupcjbaejx4jCvQ2G3sDdLjupakJ7AvovaxkOJfb348eioF0hit
8+Eoox6Qpj8cUn9sYAHm2F2Yxrx9GrtbapxtVnGBZVAqJKNCxonuIOS7gdH3OjBz
j/EPuT4Xe/Rg25NaqjXTJGsAOzqQPX0ZkbIG1oCEPw+RYeS36oOaXeWSQ7IbjlW0
y3j5qwGtuG5YRozkDRsZVrYz/NRQ2jAsoFXBFP+88Kd09lxQSbc15SQvVVuW6+jl
fOYHNBhwEz7XyOF2LyNChNn99A3qfxGam12PjmTHsso2n0ht82c3OdI/gF1BwweB
mfzUuLWhA5WSgoK/ocmBnusGKyigFIEkWgE80elmNliZ4tu9ba0uKhezRHkg+8fG
2albWI9zrx3HyJZnFj1Rk4obcvjmdIH3rDu55ouJPr3lUQIuDJeIls5KpZ21262b
01zSNzgoNt0Ynq7Mg8hIb4iboe2iRbAF6NDXNJJwlMSOpSFI290USAsRL4tuxjKL
ZdgPmDDzSasvyz7XP20FjgxgN5+fwZ/pKOz3oETn6DP3neMcMJHXTWi+vZjz12Qt
2lmQtx5hyaj2xE2M086frQ2dzpjN28NOGBKFfGxtQyFoAUtyZWi5UVSEOdKZHrVU
QdlWXBpdapw2lypI2dsrPTjADoy99Dg39L2+uVYRX2jF6T5MwrD/To5A0pJdiclU
KO6PTp7Oh81641WeQBRK7rktviVxdHBYdl2H8Y27luLpN3GfxYbe7x/W/ib69Qku
3H+Nx2TnpSL96erzNsyOFXlagt/mIAe9IB+nsusz7Rd5eha8gm9uQV4dvXzIFq/X
fnCImGb6OwIlxL+L1A+9o5DOaVYLDdUaH6LwebXeylVb+nBln3O3UTqDrU0IuZl0
U13awo+H7s8frWbIGj2WZIH2WO1xZD9Hr4ZpazoL8JC2wwqREWo/FAJwA79pzBGo
Qi7h+RfsTXfu0Fp5Hh61uHNNrrnWjMOIkQMKE02dVzgN6ZSPAf5jfQ2INhkWcW0t
5Gjl+BovlQDLCaSdiZ8NuS2CwqKfQemBkedTujdXnXgbLUR4iXPTADdYBRFC8OLh
St8heTpggi70T89A3pCny1u6G67/N8O1b4hc0gnw84h3HLv9YmuInSzBKnxztSXL
n135sQl8T2qQPnjycD7SZbvB9wtYtVY4GybQiRjGSlLSymFkV8q20MSphyQUHgGn
cT8IQaznrZ5/YPsJeoTs0bErRODxqMTcTw8bIlXYMqWU9YN2lps2w47AeTNA8BDo
l5AH7XcDtn05oRe3lB96T9jz3VyzUQG0lJfGOwv0QTCAUyg8hh1vuKEqQqNmrzIZ
l/0g3R8vbVYi+R+ZW3yjDyitp3I8QDWph9gje+RxB5hMiwATGHZoCAY2aK9mgPsi
S12z7hcusbl+Uj/APdLYwDm+NvSoelC5MznefuS23vk0fuM46FSLCaHMynY+WnEk
U1/QmENbGs3rj3FJdmK30yMgXm1EdyZ1h7urGTwILavksGu3WESAL3lFzjIss4pZ
IobnTLyqxSfjn+7t32GAYriRpf/MuTkjv36CtPbWbYo45W5ryMHQ7+kRNn+/3+Hj
s3TCLcl1z4LfmNesx+gCkqsShNBIiBSB/pUo3AoMK3Wyyf5TPJ8epwhSlkjd2U6x
Gst5bbsNU/rY73RavZEuyCAw7x5gdLwO6v+B6c21P7HXMXHYHJP+uQdrhjDm/zpq
KJjfgUcB8bQd+N6UnOOtyMSdiI2FJRWgTMrM/zowmdyTP0VJ7bnqGzyM7tVjJXQM
qHiRQAP9/xPZN1TDXnhzFlNzQXMmUrRmKmqRDSr2z/YxRrX+mU/zRcyvkwR8eyGZ
sVXSaDmIPquEHDYT3J9+NoB0QsaYDXh2iklTsMyihYahXRml33TnX+vKoPNXmRPl
Ok6qZXnqbAh1YItSzncf3b+L+nEViJkBRM9QrtoYkhMLowCoPg1xGxoQO/zqZMMN
jrNGr36HG0vwgbTUerd7pbGV0ORFCxvaCgf8FcgNrzbCwe1GgEzWuOO5qjOS/e/8
A024VcfVcxslGpF9YcpT2tcI8ZkiTyEqbyiadlCEnnBrBjSrsrfHPr3eUHHYP8Q7
dQ4VjBDfimPc9lDMjrxspPkrm09n4FUQgKhL+HGEV/8t2MK6MutDkoWyugwVvKL2
WsHYaPCcbq+CrSOKEegRhS2UBpgpONAfDQBKETbKJc5jaxS2xQjcUK23GEqCUY90
lCB3YsA1mH5pG7n1VtC+maefNibQp4pNt43N2xW1UTfxQiETSUitTj/4MgWrFtZc
P/0MvhrOZXPDHS4sJ8MGf6UWCdhi/qe2r9i9OYsrWp8ShiAVI696ggH0/6ZsoNx2
xiqD3OHLbZytBuhe1eC3Pwy8l3NcJh0Yz/TA1eYcXL2LRD831hdadC+pnmEarUxU
DyHsI/VXZqVEk3+vPVeD1X5yxwz4s18tlVoIXoLIqC0aW89hS0lO8SlwY6PKYQOl
a5Gq1mx6pb5HcXa6XRshwCi/um5/zitmrJvthw9PwfT7DLC1s5kLXmUnCgy/I6lN
1J6inEhsDSFLhKhH5CLkHo3FeJwWYsxCExG2G9WlSmsfi9gqic5E3lZm1ZeVPCqv
Wjh9A+2F3FV4/qxvKhxonT9GyHg5kvJWU1B7RHwlp/KM41T8vLBcCc+Vxxoc0DNM
8+vY4LLV5ipCG4C1P6zrWyXGCq+ZdT33KSNRN49yZHZ0QVUJkbt+eQxfqTttms7P
1tk/Imw34b8tLZcHKzfCp0/Q3FUlq72esN+OMG2irLZ9FiymN4Mu67HhML0SSkMy
qAicGIjVP86Ybf6kI8GjoRL5YKKnlNPPKndQLpRvCDTQ2M0fRsEVvI3xkuu++ALr
zNul6xtxdLtFQgocavik8b79+qzRR7yr6pcdZ+FSnvFZCBJ3lVW8hdbf+AxfSq4I
NDYY9g2wKR5Pnm4fdxVZcz/UugtjidH6w4oVB/TaLff8f2xRkYDXX3rYnprQpk2G
SFTyHFwDoFwTCgL6fDvAhuCPjTpvAuhmcSt+gN3TKNwrSc2H0lhUtIc6fNvia286
kwKloyDRPiASMPQIcPNgyfH54L6QRWMxx3dZ0BHkWG5glLW3K8Wbc22ipdD8g9tO
JLIlIzAe2tole2MImEe7+6IeRw0vpeqmq6y6xbKHD4FMJLrvfxw6HAX8cwfGeZAQ
l5Z4KQXWiCe9DYS9N6DhxuGljJ3QpcdX/kmVFRk52Ay7i6cMH4F2gEl4+wN0hU3a
HrRBnDM5Xgm/2y7JWLtW0DtmAxONtcA+vRdJMXnzwfbxx4E/MX0BD4B5trRNP0c2
BmBjyajxxaoZ26gIxdXnecCM2TFXlqD/awO21nmR5GmS6Wf/d76ASrYNiMf4RALZ
S8U8OzvAiiSA4Ky8SL7A5B2s8gKZ+8DUBnBimUnmJonlvQc90X82VKESUzOSf6b8
alghudSOQ2dek1lO2fRahYBbVB5XwGArsN9mKKGS43Y9+gEKqjm3NFqr6CdknSnW
iNXzUaFo7k0QGyRvORrwe1aY5ocnylV1zmDqUWcm4VUueuwq+NnoKMIDRqg8u94F
81TIi0+1TOBaLjAhQvUoODzu/R9utbhfMR9VDmhmRvN25sSnSVjgGq/OyItBEYsK
pNqHF9w2ZrqdihqbaMIAMaXorOow09rzeBPQaFz8tWjBzDh2oYjGRdEF6tc7M8cB
wBMwz0m+O3Tm4SGmX2n+cd6SSQWqM9fUr5X3JY70BMeP/UithFxFaQUYPbtEOYyE
i2c4HMxPnOXaZYpKwoNSIZsR4HGJCo0MQi9+bJ7O0QZNw22oI/vQeHgC7U0jeFuj
O9iUk6OEG6GLK9TvliIg3el1dIff5Oew+/0MzT2aPYr6y6P6qZJZNf8hpUa6ufiH
VIouC9x/aWtYw0AYX79TfUcELQSmRvQfLFdHcAz8WCQcPsuC2znpqVsAU6h8UjmN
XfSiu3LQsjsG75jyUKqbAz+JKZp4LM0PCGvU1QmxuNG4Wbonk1EL4gl1SSyjjQOy
zBlYTDZRBcB1coqrKQCiEXd/l/kswMbuPzmR3fRH8hudsWbYS+bbdJnrPkEtXkTt
U4HJbC3rdlVJK5ssYDY9NtNtj7pyMYm8MI1+gvE1dDkp4e1HsRq8l0kWbs9f+St2
cqtEy9082pLejXj6wKxtoiF42AsAhGD+PK9GVHdUnoRH3OFbhtYR1PqYiWSzI2Hk
XOksrnUzmM0KzcYbqG8xlqY75jWcrE7+YlBxhk54LftuUpAqV2AWHHJNnFSZTxGA
VYIAKixeBxjNHJDslwEaxnGyKSenxys83kdaXo9g2Z2hA2d8e3c8Sqby4QtLGcf4
3Cf280svqyLjpGvNAnL9oC2EoqfpPgS8FtU3O7l5Pz5T5dGMJ9MBtFfbXNQxNkIl
RUT58hTxgDHYi9GW9v31tdJ+2WrOV1BFhm4nBx9o4n2isN6YqI6wW4OqovWCB37P
GwngAslZydNwGOIF6E3D4nl+tMYyUYc8/Ty3Kz7SRCLPKydq2R4MfERFhAJjXVWZ
L4Zt97h/uZ2yEza4AL5cKnp/8AS/JZavEmjsXXXAf0eJoHyK+vNLe715p1/9JKyS
m30oPLMEK+frfpzDwL2IYd0owfjwE7QaQ48fxNC+lzfHh0sd/foJ81S1BiyYOzHd
ELkVmRvHiDxV4Vy7g87GctS23lxbbKSZg7+8PxlAHYMoXMmTrBmti0HlgAF+liPj
wWMGm4O29GNJOhSZf1gvY2lPNnWS+5sIyGTI21aCAOdsfxpv2z9s6Fu4X1HIQPuw
6fIJ8fjmjSKGaOEMnVBFecT5VTh2ZWBekKlzh9i9+//WqcwOmEWz72ZMdOffSfZ9
XkLPBhjtMkTwHwLGX/dlB0lYMAGQzq6RpiU5Bz+8u61rQfMnpo+hZJkuzbGNfpvm
Z8jlWH6MSpQ73Tpj1Lz2P9xXDqo1/gFj1HnT1s2n1Hv+mv5jU2PhpwVBdb/5Cr5Z
W0y+Zm0430ZOxMrx/diA43rVo9xR21e32GlcgRJQYtKbSsjDWTelXRDHI+f65vYb
6qeKF+qoUuVMqKOfMqRgQZC6uIdyQDHXvGCLIXLMNkxoiUtPvhBB3rPF+A7gWLVh
ccOvJQeZkzwldQG9SM7FyaExVdtJkoJO8KkhBVq1d7+QjOJX4e6gslz+s8uwnRiE
VqLqD3I8F7XTGeDYCSHi68Uv8fhy6YcBbES3UB85x2A=
`pragma protect end_protected

`endif
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ItiJYNMEdGnrkAFmpZznFSBJ3pvKfTxaHVJR6TWfgtITtsZw7AiSQIdClqfF/xFk
vTs+8arQ7wle/3cfDhux5QapU8lsJGeD+KQg4fAUhpW7r6ZnuuypP+9RNwWA34MG
ZBtukiM4OguXM6/yhMjncPTCzNDnzuD6vkMg0XRRVTc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 101364    )
O2PWGcWO+fyaqaXQNQXlzGcyb/GpjGE0+I0RRemTPz/hNnSSuC4fumzF5+GqdDBH
/dZFILtgXvKz2/yEt1Wow1yu57VxEGLsVQnE1uQeKWHHCsb4hrJBTCApdhzAiiad
`pragma protect end_protected
