
`ifndef GUARD_SVT_ATB_SYSTEM_CONFIGURATION_SV
`define GUARD_SVT_ATB_SYSTEM_CONFIGURATION_SV

`include "svt_atb_defines.svi"

typedef class svt_atb_port_configuration;


/**
    System configuration class contains configuration information which is
    applicable across the entire ATB system. User can specify the system level
    configuration parameters through this class. User needs to provide the
    system configuration to the system subenv from the environment or the
    testcase. The system configuration mainly specifies: 
    - number of master & slave components in the system component
    - port configurations for master and slave components
    - virtual top level ATB interface 
    - address map 
    - timeout values
    .
  */
class svt_atb_system_configuration extends svt_configuration;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  /** Custom type definition for virtual ATB interface */
`ifndef __SVDOC__
  typedef virtual svt_atb_if ATB_IF;
`endif // __SVDOC__


  // ****************************************************************************
  // Public Data
  // ****************************************************************************

`ifndef __SVDOC__
  /** Modport providing the system view of the bus */
  ATB_IF atb_if;
`endif

  /**
    @grouphdr atb_generic_sys_config Generic configuration parameters
    This group contains generic attributes
    */

  /**
    @grouphdr atb_clock Clock
    This group contains attributes related to clock
    */

  /**
    @grouphdr atb_master_slave_config Master and slave port configuration
    This group contains attributes which are used to configure master and slave ports within the system
    */

  /**
    @grouphdr interconnect_config Interconnect model configuration
    This group contains attributes which are used to configure Interconnect model
    */

  /**
    @grouphdr atb_addr_map Address map
    This group contains attributes and methods which are used to configure address map
    */

  /**
    @grouphdr atb_timeout Timeout values for ATB
    This group contains attributes which are used to configure timeout values for ATB signals and transactions
    */

  /**
    @grouphdr ace_timeout Timeout values for ACE
    This group contains attributes which are used to configure timeout values for ACE signals. Please also refer to group @groupref atb_timeout for ATB timeout attributes.
    */

  /**
    @grouphdr atb_system_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable system level coverage and protocol checks
    */

  /**
    * @groupname atb_generic_sys_config
    * An id that is automatically assigned to this configuration based on the
    * instance number in the svt_atb_system_configuration array in
    * svt_amba_system_cofniguration class.  Applicable when a system is created
    * using svt_amba_system_configuration and there are multiple atb systems 
    * This property must not be assigned by the user
    */ 
  int system_id = 0;

  /** 
    * @groupname atb_clock
    * This parameter indicates whether a common clock should be used
    * for all the components in the system or not.
    * When set, a common clock supplied to the top level interface 
    * is used for all the masters, slaves and interconnect in 
    * the system. This mode is to be used if all components are
    * expected to run at the same frequency.
    * When not set, the user needs to supply a clock for each of the
    * port level interfaces. This mode is useful when some components
    * need to run at a different clock frequency from other
    * components in the system.
    */
  bit common_clock_mode = 1;

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * Enables the Multi-Stream Scenario Generator
   * Configuration type: Static
   */
  bit ms_scenario_gen_enable = 0;

  /** 
   * The number of scenarios that the multi-stream generator should create.
   * Configuration type: Static
   */
  int stop_after_n_scenarios = -1;

  /** 
   * The number of instances that the multi-stream generators should create
   * Configuration type: Static
   */
  int stop_after_n_insts = -1;
`endif

`ifndef SVT_VMM_TECHNOLOGY
  /** 
    * @groupname atb_generic_sys_config
    * Enables raising and dropping of objections in the driver based on the number
    * of outstanding transactions. The VIP will raise an objection when it
    * receives a transaction in the input port of the driver and will drop the
    * objection when the transaction completes. If unset, the driver will not
    * raise any objection and complete control of objections is with the user. By
    * default, the configuration member is set, which means by default, VIP will
    * raise and drop objections.
    */
  bit manage_objections_enable = 1;
`endif

  /** 
    * @groupname interconnect_config
    * Determines if a VIP interconnect should be instantiated
    */
  bit use_interconnect = 0;

  /**
    * @groupname atb_system_coverage_protocol_checks
    * Enables system monitor and system level protocol checks
    */
  bit system_monitor_enable = 0;


`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname atb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to UVM_HIGH or below.
    */
  bit display_summary_report = 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname atb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to OVM_HIGH or below.
    */
  bit display_summary_report = 0;
`else
  /**
    * @groupname atb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to NOTE or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to DEBUG or below. 
    */
  bit display_summary_report = 0;
`endif


  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** 
    * @groupname atb_master_slave_config
    * Number of masters in the system 
    * - Min value: 1
    * - Max value: \`SVT_ATB_MAX_NUM_MASTERS
    * - Configuration type: Static 
    * .
    */
  rand int num_masters;

  /** 
    * @groupname atb_master_slave_config
    * Number of slaves in the system 
    * - Min value: 1
    * - Max value: \`SVT_ATB_MAX_NUM_SLAVES
    * - Configuration type: Static
    * .
    */
  rand int num_slaves;

  /** 
    * @groupname atb_master_slave_config
    * Array holding the configuration of all the masters in the system.
    * Size of the array is equal to svt_atb_system_configuration::num_masters.
   */
  rand svt_atb_port_configuration master_cfg[];


  /** 
    * @groupname atb_master_slave_config
    * Array holding the configuration of all the slaves in the system.
    * Size of the array is equal to svt_atb_system_configuration::num_slaves.
    */
  rand svt_atb_port_configuration slave_cfg[];

  /**
    * @groupname interconnect_config
    * Interconnect configuration
    */
  //rand svt_atb_interconnect_configuration ic_cfg;


  /**
   * @groupname atb_timeout
   * Bus inactivity is defined as the time when ATB interface remains idle.
   * A timer is started if such a condition occurs. The timer is incremented
   * by 1 every clock and is reset when there is activity on the interface.
   * If the number of clock cycles exceeds this value, an error is reported.
   * If this value is set to 0, the timer is not started.
   *
   * Configuration type: Dynamic 
   */
  int bus_inactivity_timeout = `SVT_ATB_BUS_INACTIVITY_TIMEOUT;

  /** @cond PRIVATE */


  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
 
  /**
   *  Stores the Log base 2(\`SVT_ATB_MAX_NUM_MASTERS),Used in constraints
   */
  protected int log_base_2_max_num_masters = 0;
  /** @endcond */

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
BofdQCmibfZ6KhtIiP5Qb+/HLgi6c9y/NyoeW9nD2idGHav+DqIVvexfScv6HZCd
aBV99AvBKJOYKhlOm21Y3mq1jE7LwclHk2I+jnw8jhHu/QGCvWXl8VDcd918m/LR
5UyKqdrwvx3rryCuLzx6Ahl8jodmzCB2VLQwWHQXQVk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 2070      )
ilp3Juw9ORrUKE5al5o+IeT7avGDP6M3o4OIHY+9mBMI9V6JouHfF2vEgN3JgvUs
ep1wHvbCK9n2uH8GtOiQAPop1oAu0TD0tkDYqpqmQk3fRftjgohzeeZzIoeNFHzM
0r35Hhk7NRF38QYAgBodPyiRd8QwDj4lbpLRdrJBu1rUjajbDyTCYa48JP0nAxDX
6h7OOaIKQ1rNDTL6f65WioRGq2R0DtUzBuS4bqJ+zUQ8gl5ONtjvcbim+WUNJpFu
pKpFT28sdCTC++NAPrDTsJZufhR53Gh6D18y7E269nCQBpWlclW8my0sNBkEYZ5C
3Zi/SynVXVJvyIEpPTlwPhNUXwosArSvI6+MZOHw8kDcJY2h7u1KRItdA72pCTau
uoI80Ymf4e7j9CJjtf0tOuWr2bdBchyOHIbmTh3/ilSmzPoS9OCb0O2ETVHVtveb
W/sGEh3xb8wVQ3OVATc4aDzI/aiE4y+oXmFi5sRm6uasE/pIZLkwrQcNpqyA9qXm
WoO3AkT34Onj7zGnDimFsxH/+Vr4Mq7Q40xHpa8wQAU/TfzU7euhDRxepAMV/K0G
6adr92osz8HcOsS2KA0kVOtE04tM0EZMfCJVewr3rVQ/qio+IF6Vx/5zrwzbEMbs
NC2lJuSeFYwRDJuIzBtllZ5HtomjqMyXMR9/MzmenbhXNfP1qco4JaohkqfPxQV2
+cmxVwBE1hTibtttujW9QS/J8Ge5bIDhCNzZSQcduYek3gs9CFecNq/ckYe95ibs
K23Ed+5/6wmjIZM+38P5obNUjeSNoURBB9SlLwbkywK7ce9uSvCZhZu/tkQ6mfBU
Sxuk76YgKDbPdH6RD6GdEnygzyid4B2sQD6hBlcox+xDhj0vwsaJ+p12tv1RehQL
cjV3FbZT/1Fpb1AmMM6IY72jWbYGPsVo2ZbsXQSXO+EBFZwvuqPKatRineb665m/
mZTbjqEdz8UnmPpqt3/T4IDCovOviO9CYWe75Im3JFcR68xGDquHZ1zvVe1o2LR/
fGwyatpB3909vE+Hk44sTaLOOJdabKheUbKQomD+E0OqGqnA9oeSWlRSmZ08yYcd
YavgAdMAds5R3KN06eys/vSvdo6YUli24SS3H8XrarifmjMaAv7FDTkJ2a8WmohL
z9t0KZhnT99hlNCrN84/th72vyMDlKc9ZLttZaaoXQ/sT8DJVCJWSZJehldZXIHn
LhwCfAviGL3azrCEhO9uzReXNOBeZBFxRPTngCIwPNcAmEhJ4576fBXWCRsqfFwM
jsxYuxhkiTmFqxWw1/DqCIWuEDcdq4p+B6Dc98ETVhqb/+VeIQmCB1NQa3A/ANrV
tJkdixGGrc5pXQHgpzfz7QDV6SkzkyvEzAeX4wf445E2BvCFM0QWSb7iBKgXHCoQ
OpbyyqaQY2yjTEehffUweHO7DjQY9Obk16z31WAqyiOdl5kBuJLIvHmHsu6wi/sw
CsKEWGAVSeipQOGdIpQmB+/05cbYzMFtD4hI7ompoFywDiX2kzFITRsC4e/I9qmK
26OCMsq8cqyMHxSmFyNwt2IPV5vs4kZxIJyujaBdqC161tCnmPF6A9Iq5cFytU89
2cjncBJknlMP3ezqXHiDrX+ij0MJGauigQskTCjW3EtwkBxKsJ2RgE/jPqZgG3G5
wQRCVluZReKhv2Cs07xgkOjwMbuP/eSi6DffCD5dMSfzQj2QCMmW+thdmRCsRs6j
DQVOCIR7qzVjofpSl2nP+nDFz7obQcrTyUuSB8ljHArum2x3O6NEGmPEJj4i8Igv
rKQqIRasaOsNO/MpzzF5z7Zk/z9oziXVzQCb4WdUV1sjQ9k6Lec/p/r5qAHmMAs/
0GPImdTx0IqrrtHpPSCK31sHbofwbGIABsFqxmB4wV1AZ1tWv0EtdvQW9uM+2irK
Wnkjm1M5HjV5L67wNa421fmAf4xdjp4R7zC/E/YlG20gfB2D0mjXszTKXPGqveHF
tX2C/LYEikyAJ4pobzCgfpqAmgqkhL7pjeboHuRHd+a4lfYzst/8Xn3DNUgj6uaH
fNHp8jvXPWvCzMXcRcEHMosxVlErFz/rRZgDzBreE2JpwbK6hteQ/8eJCyZsTUof
cWsueqzP7VPLOb6mbrzSemJ5AGwUr5Tox4jAiTXuWryMj/JddDJzdjk4NwpPauSK
i9+GeJ7QYIbPsS650Vv3tC/EIRfBUb6Dr8Y2eLOS2shipb3HkA5LXHhFCKAG0Uf9
yQbKjk5f6B8yNxLH/mL20jJtHB8F91WiNOLX8z9owOF0SmS7LF6ExJkcRwy1o6BJ
OGRCfQtrPiTJRGOkE0Fvu5kexuQzdNK9b9Yo6MZ2X061lLKeWPKu5VxDMFL1v1QC
zS7KvXUiWjXJlqo1nhiju6ROK5Jbb+Tw1ATzROhR8ZttrmGP+gx1LGojAZfGQbLl
XhB6+TThgcuUlP2RGmS97g0TnRWhZZjc5IUUHzGkIxvBV/LkKn0BnRrdu3+ZvbZG
J8EqzNgtU02W5s0LJaL+8AuoGeXO+qgmRpKqzVH3O083Nu2ko1/T5Nr974tUENGZ
ySDnMDgmOP/nWr8oGPBJ1OdLE14zSQBjVEj7BISsTKh9RzCngzT1I2iWLvabn2g8
z8LxOkn8TeYHHQMTVYEEorzikRC5AHF7RTXj734xygjjcFSWQrOgBiLAiCrccLlo
kGFlBVhlYz154vPPzU0QKsOdQ63G4cnvYvkkY9j+49c/OH4Ulacpcj3cNWVHSZBc
GIDlJ6ntvA6walzvfS5nSA==
`pragma protect end_protected  

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_atb_system_configuration", ATB_IF atb_if=null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_atb_system_configuration", ATB_IF atb_if=null);
`else
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param log Instance name of the log. 
    */
`svt_vmm_data_new(svt_atb_system_configuration)
  extern function new (vmm_log log = null, ATB_IF atb_if=null);
`endif

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) calculate the log_2 of \`SVT_ATB_MAX_NUM_MASTERS
   */
  extern function void pre_randomize ();
  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_atb_system_configuration)
    `svt_field_int         (system_id,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (common_clock_mode       ,`SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
`ifdef SVT_VMM_TECHNOLOGY
    `svt_field_int         (ms_scenario_gen_enable  ,`SVT_ALL_ON|`SVT_NOCOPY|`SVT_BIN)
    `svt_field_int         (stop_after_n_scenarios  ,`SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
    `svt_field_int         (stop_after_n_insts      ,`SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
`endif
    `svt_field_int         (num_masters             ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (num_slaves              ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (use_interconnect       ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (system_monitor_enable  ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (display_summary_report,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_object(master_cfg              ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(slave_cfg               ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    //`svt_field_object      (ic_cfg                  ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int         (bus_inactivity_timeout  ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
`ifndef SVT_VMM_TECHNOLOGY
    `svt_field_int         (manage_objections_enable       ,`SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
`endif
  `svt_data_member_end(svt_atb_system_configuration)

  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

  /** Ensures that if id_width is 0, it is consistent across all ports */
  extern function void post_randomize();
  /**
   * Assigns a system interface to this configuration.
   *
   * @param atb_if Interface for the ATB system
   */
  extern function void set_if(ATB_IF atb_if);
  //----------------------------------------------------------------------------
  /**
    * Allocates the master and slave configurations before a user sets the
    * parameters.  This function is to be called if (and before) the user sets
    * the configuration parameters by setting each parameter individually and
    * not by randomizing the system configuration. 
    */
  extern function void create_sub_cfgs(int num_masters = 1, int num_slaves = 1, int num_ic_master_ports = 0, int num_ic_slave_ports = 0);
  //----------------------------------------------------------------------------

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(uvm_object rhs);

`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the OVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(ovm_object rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  `ifdef SVT_AMBA_INTERFACE_METHOD_DISABLE
  /**
   * Function set_master_common_clock_mode allows user to specify whether a master port
   * interface should use a common clock, or a port specific clock.
   *
   * @param mode If set to 1, common clock mode is selected. In this case, the
   * common clock signal passed as argument to the interface, is used as clock.
   * This mode is useful when all ATB VIP components need to work on a single
   * clock. This is the default mode of operation. If set to 0, signal atclk is
   * used as clock. This mode is useful when individual ATB VIP components work
   * on a different clock.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_master_common_clock_mode (bit mode, int idx);
  // ---------------------------------------------------------------------------
  /**
   * Function set_slave_common_clock_mode allows user to specify whether a slave port
   * interface should use a common clock, or a port specific clock.
   *
   * @param mode If set to 1, common clock mode is selected. In this case, the
   * common clock signal passed as argument to the interface, is used as clock.
   * This mode is useful when all ATB VIP components need to work on a single
   * clock. This is the default mode of operation. If set to 0, signal atclk is
   * used as clock. This mode is useful when individual ATB VIP components work
   * on a different clock.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_slave_common_clock_mode (bit mode, int idx);
  `endif
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();


`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the ATB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the ATB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the ATB SVT
   * suite. This is checked against OVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the ATB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif
  /** @endcond */


`ifdef SVT_VMM_TECHNOLOGY
  `vmm_class_factory(svt_atb_system_configuration)
`endif   
endclass

// -----------------------------------------------------------------------------

/** 
System Configuration Class Utility methods definition.
*/
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Lk9I6TcTXnN2bjhFOxfjVDO3yUUvRzTTjYxm2zY8J+doxmLM315lAdkw/XT/WeQR
Df+9XbvzT2yVoymcK4DkFvwowJPOxgMw5Q6s9bCDp9Iod9DOmQtrf5/NtII8k5jC
3TziCSIIRA/gQBTeiAwxcJNmKRgsxwpkd6uchbkJRl8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 2919      )
2UVuzCvqsM8DRJgpdhOUKOhcfstvLdU9lhuHFlVwI6gIhK1DlUntm/G4gkNWZVPc
RWDddH/jnAh/i5SPhHIA5TVmOiwkWFtNL08zBeR/nDCakPCrk9HbQ7Z0Y/8P+bSQ
OETlhCGx8iXYaT8558PxDZlqHSYuKRWMJERYRd13DJ0TclCO0dRjxHUqfqVxZvwd
uYSsNfsUTUsmiWjQdpaabpVdTQTCHO0rX5db/BPdLuyaXgn5UqjE9dd1FyofD2dk
ai6QeJuebvS3ey333iNZZt3pGqcA6VXK6xj8Tj9b1QDknD+TKZre71nDThw3sanw
b3iYc8LkqlPtElAe3QSq7J7Spwrwiru3qQx+dx2enEDUgUVx0kcBgHzk9u73whqn
rHeDh9SWTq0ORBTKkRUawH6pDgTD6ZleDlmVloRm8BnxF3anszeJhYlqo2vQpkN0
ntdgVF4HOFF6/sM/1Xsrn4oWbDe0YVHU7sM3MBtUn9DXxlaMvZCoLd29tRVpqAl8
4rklfqlFwYfoPiqgRDwx/JIv09nXz0i3HqXju8xiTgDtJTq5rIlDh3PZVTElCUhO
i69QW38mRXuwuXW6M77u7kIod3f8qNMD9Mnhl7mL+H+gLJxiQObsaEQMEK6IJ51k
2LPgQkFxETgCu00zWC8XInvMhyPHxv+0PvtwG+w099r6k9zjvtPl08YIbqTS7iIr
t56MXiiIbauO308e3PX/7y3ePkAsl5vZoiyNNC7FF3SyW5vfAHslj569T67Lhm0U
xGJ8c5vtx70rKBqC2FC2Xry3//Q+E9kKcfWgglKWVoQjVNHj+swuoKy1qFHW0eaU
wgVwvX4BJoQ8105nBLEEbgEEgkg7w1BDjYtSVMA4yY4AWQ2ZfvZOJZmy8/+XOWWx
ht/dFHeNLSBtBPU3mcA7UOvEfniokelCfbbKIvekcTI/Q6OhycT2xYCg3NeOJRT6
cgRjC8YbyvZXb2eSVczdFGOo5OgOaXaRhk1P7537A/j1eCmSMLFZVsIh3lsGUM3T
d8+sWO+W6kuqoMtmd6Nypqd+rcBgJ+Zr1n6A7AEDEf8B4GEWXLwedGdeCy3FZL4E
49QO8mEusGUqk/wiFUFCFeCxA6ubvXK2aye2h5Q5aQQOqi1tMzDHnpOBYc8UA/7t
`pragma protect end_protected

//vcs_vip_protect

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ggAnDGmj7WUfvrEqJ5+VoJFjLQtqcANtphWF+YRKAYTaEHN1oYy6180dJky+Z/Cx
1shlkG0hZ46XaQnVPBfR53raRaFsSdjXncY7l2d0Wc3aAUxk+ybR5ventUsgkhyf
K6Bv8tpzUB2WL4RkTH7vhmtaUQ8md0UVk3RlQwCvsCE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 64639     )
MGtxGGg/4eZuVMUii7FykNNC+mqPHpZRGI/pXXPWHbte5hr/eCDOST4T1tfhiDjB
xk2+ucB0obxuEmyYQ9WBueyRyCH/0XayW5hNrq11oKo3U+PFfm/FS7VXEhyVCFsd
CEJVPWcMaRu/OZ+Hik4XZpo2aG0skQhzLKbo02eLiEZEueo/pQZcJPsmu27vIsqR
BxmM72g9Zgu+cw/vlgCKgdG1TeGECK/d3CwxDWGFnMgNh/gXZ+otSHyhmaqApe+K
4ZqxWiu5jSLGb0lyx6w/1LpDXMnr91XTRO7JBHVnlU2ru1Zyb2iW6lQpMfjCx0yh
TPKdLPrdCqf3asRVa5e7tGY6zl+gkX+l9hEnMRZkcyuqInHmRpD+lMpTBYBQekGS
+Pj/9MjbV2ENFlEIc16hG8OLeCTL7W+iXpWuyQ++vAQCLaKk8e6J4QDdtWLx9J8v
2ulCB9Ob2ZLcEn1z6wO2qluybtVSKXZ4NH0Fagq+FXWXUS+lhJGxB8XebqUUaFMw
KYDlSwIPlneF0jv6EQ9LZZtAWuNHz00f8Jlgj+JrzYisG2YwkTTb0EFwrkSiVHGf
/I4fuGhyGCFRxehOFiiXVQLyzP7LVxtW1l4tZnAk9cq0DcKckfPoxnJIcKisgAcG
T2rpHaNJHgr51oIGMviaHwlWWamqBr4S7QBsm+9ykPZeVCcmzyjf6ODsGUTpmSqT
o4aP5qv25R+jlMihjpTFzNsU/HRpS2W/3CmRFto+B9/gQu1SkKwoafqRZ6SHoV76
f8v44pcDNtvDrqVvRnJwvANJCQUxxx+y6YMo/4ysYAwEpn9UPTFYkWLuVPCCWAe9
MBFbQowY/vZWURwORcYX2c8yyTSLnG8se8EP0G30TtFGiiltqWoWrb/wERtIQxkU
Tcx8uyd0+M0yP+WboZAHLtGggYrXw1YX3eZ42osIjzhsnhMVggGJysRnAfRUyBQ/
YCSVnfoGzEYQs9ixX/9MGa4beTMgRdh2twJmO0yFx8LpgVZ5uvjntCh13JM+xjiL
F/oxLonr0K9La7hK9heTXj6cdUQRLjn3smwi0rdtWHf9jOIiwOf399g9bce00rSD
ziGLT5n9ejeDO4Hxhh6GU7CnSU1oeI2mr7gsAzlD3kyIRyBIwpQuaPLA+lOouxQL
lnxdj4TJUisuT1q5vjJq1RQe7lOhLvJSXeOp2oXyuK11PLzWL9Lxrp5/Wk/t6JSE
muf24ox/sOyLTLOWR7hiH/Aef0GaLCGOjoU/BWiB4Su3fD+1Uh1lY323pT24i112
5HGf57C9spYBug/3mwjYoio9P8Ki57/Xwl0TSJ+fF7KmiYFXm5A4TuVhWb2naKX7
2PCy9gq1vfcQhvNjViylaiE8t/zvlWs+dq6kNsS1e3T1LbS3D8hssmKwwn8rRdo+
UKanLpad4O9tkfFiPuXl+nmZ+Ax59LFW/9Mobz78X7vAxyH6aSZj9P/LlPkleiOE
xWZZMcCO4NBwnGGF+IrKE3Kmov4NPxu149SRDWFOl5BOUwzRzADFYjEh3OOyCVfT
qrZynCj3oVwbK2Dauq0iYs0pOttOHwpWPpDq9UXW2QbmNg4Gf8fjkHExgtjEhemF
lB0UwFhNU7DpjJo2jLLNUxjFhUGhBoVjr2vD+j1z3zUJajfi4lwbhsNp8kC7gUGs
rdeZU59waAWp9W2DnO3PYxujTsHnrsA/PVLCdCWRM8KlX8gpo35Pg3FKgiwPb+4b
7RMa4NOjaSHnLjDP5OOIyHlaRgE7sv7kRU3K2d9RimbZt5+xJZNYNdmfolZMCOR5
U+K2LlThps6H+fad4ie7fEGjUfS+y7eGF43Fdz0NuqoOEtC2R5fPwIPFfDrQnkW9
7hNGyjbGRGUTBFttxbltZl/SUrg5wtDcKyzOA0nX3/r5HqKVGzRMIPuv688ep3cW
APAr2Ro+KZqIyI4S+yvr0cep2U3sdaW+NdXVtuTBZn52LPhFB5g/j13ZYu0dUVv6
hBgkFcZkn9JRM8/XBiFuDm0d4vhgHH/Kbr/eebb5+r/Z0z9ytQWaUxRIKjwJMT2e
wM5X1D+TBg94J6awR2oQQzceh+eQBGgHIt1jbzOegm071DRNeT3K8XpRI48RjmeU
LtWGNx3PBOnK5nFiyYhp3x7qglYoYqlxHY00yd9fPO5lMyzdvHjBIVm7xrn6Uj/w
TKjWBu3pmCWXGHMebe8+HIAvASr/R5TJYfwcJ+sReWQvKmcSX1xSLUgS/suSIAHE
LQlkmY5PNejrCXp/I6r57S1GO+d7njlVkVvi6neF/bve/DJjIMlcYxYpsP2ZifYA
TsOvyDTfK4YrpHdMqO3aZxOf8t1vooylBfHjIWmvRjz9qlk8aagHjKDZva3Jo6yn
3y6XFQ3RL2Oq2CyAV8psXKrVzitMzu/jysSVV3fV371ifd3o2v57I4nyJFeY4LmK
B5MASde+ASn2G/U0dU5x95ciHEGvRCFw8pS8X3Hj4sxwQ0FItZriFFkItIApulmp
S4mblXeXCpdUZjZQ48gClUc9Y0Cxhpv+j1sf3WvMvgMWLfrSXXz65oLHn28Dirts
NHX5nlgmtC/5CGZkamurHih8T7lBqAXZU7NKqvpkRiElVorbDCVm/szfJo6TbWUk
v6icZZ0g38TFMBV140zCOA2PoUICxVqJdELWw8u9oVW5kqhdHHkhAERx2h8X0xhG
6wpYuwFszSnZKIPo8tdbJdqDtz+Kp4m3NH5w9Vmi9RDxlOssVX9kNGRkkzivQeOc
EDz41Afc1XaEa0Tmu0PJyxj0qjTzRJtvMRZwf0LJA2Pn/G8aqGo6RsDh1FeN2mzy
65qskQNHYQqQmH8uFua6bUVO/EHznM2GjWcfVUeB8UhOBikuGacbdax9M5bY/cV/
W47NWK5AcnL9wfjR4SaIo0nGbkGX40iZ6M1VA6AZGcIhBTTr/85579A41kM0yl4r
PSxDif/5plo3hthiVADsGK4CYEsVux4HP5lG17whkizT5dEnZ+32L2cEpG3qjVhA
Z3dcJq/y+MNAeh7h/bCIUH81spffYZm065e9bvC4DLkK3KmHts+SGXLlYWJm7880
Qqya2KLaGuCDS2oCp5y46qnv9txeB0wCzsD5okNaHD0ho8+1ykZykL3mhk/3MJxn
wMYf4/23bd8tkQ4uc5zXbGVjvcDxPCfJ6T4CK/K2613Xy8C5KPo1CJVGo5r9EdUv
N53gm54azcs6JLTjq4p36Os/3UVElLeJ5A0STyBmV8Df+oCMojsTXg5sLgDfwLTF
Zps+003syPz6g3LxEQskTjg3dFJSV60p1GDRTIVp8mXaQtEjWOTnMoLeuZY1stad
k7Ojci/BWU9ISq5NSjNIso37+ITfxVvxQZk6vzHPNuXrHA/qQMLB1lomaZV30ben
v5m2HP8QcXc5kssc/rB8q5vAHYWXTE1BdmVhfhljUv0+Fdp3m3I3GdP1jj8n4lwy
B8H30GF/W1YhbSH7hPQfthNI91jgF7IIumO/cJRaxr6UNwEWQAdkQdeumVjDtjec
sXL1GNkiNK4Rtxqsj4Q/c+iOE95ChMoQL0SQgmiZ8P24TZb4mcX98bwxH1zB3NGG
KSNrI6pbEfShQi8NaSle6OT6OIa6o+7h+59MbtNTAb/ddxuFFqYy64Q2X68Jk1H8
v1lD4zR6yQTVKUfolpYTT4pmw5rOnmfqAQVYQBN2ceJuNf7TpG3R0Cu6ErlXly3t
iYQk7VHNqyPjWy97lGrgsoYk15Anosk+4tS8K1pJ/Vapp0wUpgFxoN8Eepx+c3QZ
tdS/VBcKWaN6OQV+yf9FKffAogxwBYLqsDpBeaxkrdDCbKxSLEiPGmwelNUKhGtI
Ct1HsLaWlRqs/ulI81Nogk5kAZWAMDMvhNPQfZmkoctAbaCndjeFotKaviJ9sOfV
FmGd5nB8IRzLdWcQ40oPORbMBkQ0zFq2RSF3Fekb4bYQ8su3U6WSgpTQEKk7BIti
ZWa7ycVrIdoYcItM9Tmv9mDtQYvDIyTv7yTKQ1DaiGjCjqVWGSqFKA4ztLFdsuvw
rBmxnUVRT1X5G6VgK22Da5L809y+Yd17K1Iu3C64EzECMUG5p3OWA9nnj5EMwjDe
dyLKI6/QvDH/Z6bq8gduUa2CMH8TYRsxh4vgjM6TPgPEsae/fwnyZDRlFyMItPKm
OMdedMcQAjlI/qPm0yEQmky8K1v9JkJlb28Z2rtXLHAMU7EFVvMeQQpnGv2gB+jv
mD9Dd5HdMdiAMRqij4z2m31gCDPQCedM8LXlgVnYKzAPHRxBrqpbvktECoV4VQ5m
7nFqcWzDEI5DHezDamBmeLo+a78wN5RCZgseqh//y4fKDUbS/g5ZrBfEZgm4Xu/u
pBRMfF1zBBZ8SAm5Dgbc6SaZZibHErFvWbO3pWLkBDNsou6EU7xlyJU2c+O8yvmw
hD86InlsFoxoRUa61/HKdHgsNuIvSckVPP4QxquaTRkEO8l6+HxKATOiXRHRvG8N
v4BQ/SwalXhT4HkXXvls5X31nXIwa0MYV9mILR0KxJL+XRQlvtFz6lFnVdAqCXBP
dFg8Tly93piWsHjn1BIbwc8MkRTTPiJRkPPcyLp4IGN2KeJLzPqccDrGHZAVudCt
47JwkuPc0JNJFThyOl9fy59gd0IPFAObHnwNxGRRpmcnI6RciL3FAIwdHzrwKfvw
UELjZQxPysLB2Skg8yubGHC6nXoOW8FDTHMzlS0TYZHgLw3/vys0/jYMhTRwwU97
DocCcflwk5CRNqhQOUnff2FEdbtGJehKG9SgedHldYPiZO5sjlWNNkS87l2+Vg9K
4m8BhDxtPlQhCj9jB8bNGO/ctZKytspZmxewGwx2Ny/GNRu5P8eO9W2uNf2y3xcI
wSUMaPs4iomk8mGaefdX/w1Aa98s5uKoYCzcn4fL53S6Jrd3G8NtNGqsopiHC/Te
TiDplLkHQE7HSU39oeQV5BAG1DMxZwLIbu8/fn1U5z5twfeQ3C0MslpkLiBS4XeB
q1gFnW4+LlpWKhP5+phb3WDddQ/0t047bHB/W8o7Rr2tMJ1ko8pGBIkQ93YoGT9w
tifVkLQEp6b2Lh3F3ibVGGpM3G1SnXdF/gyIeIVasCexrjH38GPPMp/znmUdOw6U
Ubw2hXSVpBgCueWB/Jj1LVF5Rx5ZdENtT/hwc6phGO4sc8gNV4qok295JgAWGgfv
dLFfMkSbN7ZoQMdmk69zppnVvHzw3GmRp45FpIExZ/0Xilc8AGV4LUsSIXM9yakV
nKGRhphdphYI9oRMFyRGJ3uxgeIVaemPxArt/Q2jzHkVzc/qCtiQ9aklSIvsX/Hf
fePGevnot10E8BW1rkSfmLWjnwKK5lgum1Lo5D/cwPlh/EcQ+i/6T7wjR+boahCz
Yooo7sV4OmCOcNdDCy4+C6wpl0gKcEs2Jdd7AL5JYImhzpbAN35H37yx44TvHNYs
eDHI5muEINnroTVvocDHoBzagEvGHS8w/dBJEOi0LNZxw3hQf91zc/oYG/Hb7kMa
uJn8yV4xpIsYE2D0U5ixLVqZCy6QfakfZx+hWyF/Tmf8IHrUHht+JOZN2TmVFDYp
WaBJ/BmV+c7tFSSnXza1h3RKnY+1Myp6rpfC7xqbyf6321Q/ChPdjhNkhyES0Lw9
Z7K4ovAkCpXmEopkwDjV+cmUKNcANES8kd1PdDgb7opecZjRl9R43XZtay5icnpX
/gDXtd+Q8HlKKymaKb2Yz8EA8ry8I/oSGiYtYAZ4c1FNQaoAVovK5BnuJAq3MbKW
my9GlUhQodHajqOOcor1nVKjMecGXd2dtm0Ftiy8nhvpep3RFe7x+dRGD3cEX/Vh
HNqC+Eh1uJ8pvlpAjiC1p88UCS6um/QY4Sn+xtuwfcoxo9o4ojsPk2AnGxbDaM2H
06t3ZoHcDqI9DPmRoyfhg0qrHbjaRYGEtXS+6SvU8iQ3EjuImS57JSnksrWBO3w9
TXX4GndH8GFiOlouzZlRiUNcUN13KRUB+ZSeO/++kGlr7qS8D93wNitcviYTIdX4
TkQBXc4UymdiTkyOYN2OwS08lNSohmK7dgcZ919DZEDQzTYJUEVhyBQHYPHvVhUp
6umgbCVsK4RIZIeR1xI1noU2WP99+WxwCbavXttK9GKv2KE9P3vzX2FogEvKMbDa
QsuLSanDPRnD8Zvj6UOLfvykTf8spSCx8sVngiGF8LOV7T36FX61muwhbaAF8mft
JtAx8FlV9q9TahPUr7d31l5kDNKirlW3aJ62aIzHAC38dn7y8zyOpbst/jttD8n5
ZWE0edFY7GBsAdz3Lk5BtSo1RRc0CaHRrReAw8pXL1BQONMJwLgVV9Mqy6y7JXyp
hvrkWj089ceEyuWYMbq3o9B22HZiRxQYJgZNAnsIHuEKrq2T/J6CZxqXpyyJbrhq
4fui/Ggod9Ez8i1IEpD4u50y2M7WMaO2dpQ6LgESywE13TvdK+wfWGUiRtnua8hB
UZ0nF35VDzSgG3l4OnYinN0asDyF33zoA5FXH3FVgBgzM97BiO1JlPNQkTs4m0Jd
gRR6LBasL6+DuTU48dx8x3WyX2r5k6dQK869gdxOxXwlx70bE+CmrMNjG5o5+vHk
pSKPP3wXDicNOMCpjd55haEQpKRmL/mixsjeIoTRl4pAwpw9lFBBEUYtdqf7CWYZ
YCYhiQQlmOcD564GFbyAxROX+bQQ2BMVrV0ABTba9ayAkshEqZsLWEarlhhPuK/0
z2nGCBPia5eN9kJ5YkpsC6guc9h3TFvy6UUAxjX1EHBs/WlpnikL9Jp46/NnD3gT
ykgyUmTSPiEKARpuGmQPrbeu83F7DRb8TuGx+NkgOVPvYodAIbG03W5L6jsIdS7F
l1rba5deUJxFxEyjhRT0arll3QkRUVoJJpn7bAdJ2rJKBRJ7Bw6O7oB5d7+No+Xu
Jz58aDr0ZPutT9BeF6vIpp5n8+Z0ms4T+wKKq2K1n2GuWUD1FRZOJ4ACXLO0yicK
Y8nPEZk7iYwwk5MvZQZ9TKUq8AjbUEr249E6TVzOsO0Z5RxWYYhb1tYcMu01ZgxU
P5MfCWd29ciNfz9hZkK+LPuvamE9mqqAAa7DS2CA579btVu1Npq9krbQ1CuK8EnD
+xmXMu/Vmw27fJRN0RmMpVaHx/cJ1xcodlG4ekdgvIXHEWdIXPgS7dDbYycNgl6z
Sj+dWk4ykagzH961MAeZaHGursma4aV9khb+PrtFp5N6spAeSG1qMi2ToXK3SQ4Y
QWDEu01gaXxYXdIRjfHy8AKjOnPJNRKMGnvp9kNRciz9NUFX1Jp6PJl/larMWZ88
kkNrrVHN30nzby5S3ycB4mnzp1ge9M8yebqTym1c2O/Y1F+mMd9s7qyvWMwx4Yuw
i8UCUs8fdGYP7iv9e6gyzxGRQhiBy9YB6Jkaq+JOBGhJ4He4s9dBpjSUMTfahmy3
jLTjpo/QscgMxieSMo0LELqlxfl/qW1gbrVGkdcnTv4K1QGcVZYxn0jfVmWVSnF4
lCyghIlfeOKrHsbUAthwMizV49vpjLw216fwe5t9rqK10EqSHvKIZHF/DBzqxNs6
0PS2w1foBLGTfApkvhYcd8aA+Zz183ccSzsSlcUQuZW/1PYCBgPuMgCYJl8DUsmr
6utgCSyRERT19aT1APNWOWo/pNSbOXUk5J644ICTxaRh3MmMIiAGyz9PlZCG0oqr
jSg4bmagPsTdpWyblv+DJqq7PSJB+YKJ3qdU0F1jqV0I6oJorKsHhDxrSra36Ats
XQK2a92XxPQQ2RyAMvk0tnFOODmByMX3pRpgSxEfI6YaxT9OEnlJ971+HBMuGF3W
7uReW+U7n3/mh6WlutbrFuBQzZ6IqTXNxJqMBQa2egDdvM+5FsFQIUk/nWpLWNCo
IfD3jdTuDFrhZ8wUtqMbbU5kcYgLnBy5WtbZud6ccl85+ztQrNxcws39BX9fhThE
J94Dw+MggZ5nP8jtFn3Mz+jFj7WvAXxwRW+M/FnJ3YviFHhwHq1JE1bgeDRd1I0p
Md2uz8Q5FEno3f/inKeVmbYadOrcMLj3BZAmKuoySLtsS2f0ayv9fLFSQP/TZwK+
V/TH4Keyy0rbALoR+Q4AXRw0imhX/i5d8dsSHqO3PpUq+1+0DXqiVbgrOFpdCxny
diVaxAtJFZ3OQoTwlPgSH9k9XyPdAiFwNlNARQ/d97ekPBzHsydOGGEFEElWgHi1
P6cZ4iioHokrxsA0zIrLZShA1dV09CjkcTiXoIgjK8iCLbWcO+MG5XaTcAcRx0bV
mgLii/1Xcu164G+tAXsmp2+dCa6rPbr3tnMni5GOC3895WaIqH4yGUinRfzkB2XU
WIHyALUuPcsLc3owoa437unzTsvURmD+UmCzv35o+rm2RnTHZ6SaEKDcCrKyrcGR
OR9s3fmOJMRAUkRF/x27nBnqYsJCIGYkWz/rYiXQle1aAn/ICX1YQaVztEtZyPGn
jddFtSK0rMBEKnre/5D3TgWJAxqXjWwxCxDWYABbkGRDqEojDtH98M/SQDZSJSMe
IMWbffHqtEIlhfShtjo4Q96BFmMIXfL7PuZRY5I6IQaJJ3omi5YXzOP/KFOlOe+L
IJvdmiFnSeC/5+1pyCmejljI7c7lTSSSXxFsHoDT9goXwoJo9CrqABA5OEgFAsAY
C7tIxDYc3FNq4YFH7xiuQYhxieZFZxSDQyBitn9jy2jebkQGAAQXabFYF8uOy/j0
P/dTVkbacYVhoyyLahzi6Yw5eOVedaDaySMuwbH+CnU/e9eKczXs5U4xZDs6xYum
SlCZGbdKQhB7tcyM4Ol20AD6SNuR3snLqtIdr6ldnA9ZvVzkFNJtWswA10pIqqvg
30IhXU00zdm8tpoF0IhyeWFZmynX4pgLnhe1hFn4WkBuiPihSZ88F7AjnERyrjzF
YtoIQ1Rbm5TkYUt8LnV8jPGiiZq9yq+KQFPXXXPmdi03/FBgRabS+IqbeKw9rzsd
ZNjb669YlFnEdEf8SXSi4bCwKhcmQdawGJuTldGnDNVc7PxdAWU+grPSEJ6+nQqY
nI19ZbccPkbvNzLUomkrSthx3cORwJsTDgZbgqVfhOLjuSnKEpaT7HPZ89E7WFlb
LpOm7SCXMsHWtlyxvqk5ilIhY5bbgHSWHih7JniWVJbm4MtkOpY/PvouEN43tf13
J+cdi9FFz7Z3T/1T7Za9nZAjGFaceQFiIaHF+vs5f9hvej6xPH8Wg4BwbkaiSDI6
7sGKdh7hx2QFvUt4MNoghH/zXLFl/MNurTm34B1pPh+eGlyj0vuDUr8enkxGBLHl
7h494RlMafA1c2Ni3SlL3gnO5bXeh2nqt0cW4vqLSNSiDqmhJj1Q2uakD8gDROGr
szUPxN5ifgJ3dl/4XWTtI9F/mp/WIE9cqovmdRJ8cGAEytYACU0nVnAI1dbQTp/h
6bC00jZmMsgaO0QOD+CIHghoMZLhGoJQi54ROVuN9YlGKZgw9DZLHZRF/x8kUxMG
ucWg7iCVTgEds+l+Tg/FojbnwNBQqBqG7PlbXnx1Pjt8q9/85LgRU7HfrKsOSEJl
wv/DO9mVn1IlEI1F2OAxBeLI73mCfY0DQZyH7zhoC25L6ss1WgQ9ePjtCA3/W7O4
Ri45QaSDm/rR6t+iwavK4r8i+X1hULYt+QJ9unV7l8G3Mxn7SDD9o+2dFlhC3SXu
8O8A/YP/DE66u8d2J4UnNRlMAPTwcUvMvm2hLu80tTQ9CzniToj0tbZkAMuztgZi
ProKksvs4sRMpChv9Y+8m/iF45JxD4jMLHlpnMTZ/F75G/QPdQbNO09u0PKe81Yg
ULvvPol6S0DTatXja2cBTQsFHRpfX9+/b4+RLrDO46/VGtK6B1c/vbzQiYpz43YW
XDX+5U/+PoZTDAyvoBRwo8mKA1goV5g/2uVAbbjGH5nCqRJDJQVvaRVPH2aXS6iZ
uz1Gyv1TRsCo1hNOsIpj83aHPdvHkH4D5n5j+yCBEZ/7JGwHX+nXua4NRpjlFmG0
wBGs9HDTJJcPugPVwoimwmOzOMkl6p5drL1rd53zn0EzkFOxKnvnIXxx3zwumJ7a
zIB+IhCjluVzcMbsh12iRm1cLKjliLJo7NT6MsKAVzWc4MqVn2NRhELwCbHmk3HQ
7nDNWi5n7uyi9iDuCZWPjmKFBjXVCJi4OmfWGbdJuHDRUoVIzv2wu7HW9b2hoB7Q
xZPFbrLtvJkZoezE1f9qLnaNcnrkN5a0eucCLcjbvrSSKMmCoKwRx7zs45W6DIjz
WeQJY0fbrQq/EzDv7AYDpUmrW4ubBdYcgD0eOTubp4Z8SNX3Sao4liWEevI5LB5k
x7/XUsklILeXhuxA4FH4BZS2YiPIoscjjfBC+udmjAELXwRJgsYQuUKripxitF4G
gVXE51+Fs97Rqe9ujaiNY8WP5iV8Gufs6bW9gRyBEDvGqAcn6yakOMuhR6xivHqq
b3YgLIVYLpLn6119f7ubn7+beuStkYtW2JUGOX/VTQWYcczRa7+7iU4AgmjeRKfa
zIimS5uheO0+PYSAIC2sW4J/tHX3tsrVRmJ/XsEIxd7kNJTJFvjBpqJh1pMkqjJ+
BDIyisfha5ASy2wDop7SHESrubVxzkb9GCE5KDGl4dIARjOwvZ7u3iDvW+FfMmzo
D2Gc8jknbXrpJZ39n/V9CbrPlO4Jb2CTGFCo0QoncnaT5ACq7VyPdfsT8Ah5eM9j
nsVxekZVpNRffsNyWVKcWsvkrMgN8pG9nXPgX2+wFK0AN92uVkpzG5i2KoUWz6xV
szC5Hmoc3e3NWPkRrn29gNO6aLZnLEg4+GMb6XSuQKVqjOozXhzN9o+OmaREccPR
ztGRBYNuUQmwuIOVi4edpAbq6DlGYh6H2yhanzHLGcEtTkCo9T9WBy7tcCE9af3b
lb+Dfd37dKF6SMnQqu9Eo0u+wj2xyoO/73uSSHpuk/5PC++ECxtol1eAX1u2Uy/A
1v2qJwrJS7KDulrPLP65MsNxVtbyYzEorarymNa79bl3zof7UPIEX+rCDkt2GGWB
pTQJzqN4GiYDtf6rIKsjVvTpmtDCY7WZHIE9GUDgmMxz7Vy/++YJUIvXSHBpbQg8
+iAIFchvc2BDLp5gC6hJ4xsnNK4tnWKYQAXrgJPZ1NQb1/uTvNhvr01BiPbGB/Ts
IRGtOcUEASl8p3AaOjStNoyWaDdnLXUfik9zPkNhj92ZJoexPq9NtfmQc6W9kXrE
9xOyoDUKlNrpJVFxUue+td0jGTR0y1Gp/x6hGiPq219WsjzIH5Sjq+Gbc+UP6y3a
/+FW9T+vqk0Rxfhy+B1/X80Lid0q0jBNza/a8x0LrpmC12UBtAFfac0rVmz9PSnx
Sk42qhpfCUX9RSs4L4nvedNbA1/4VAlcvsBPkbUnPpvsaCYtJOKi6RqgS97oziNy
iLPR/YScRldCr4rP11aP5UMDJ1kF9vnzXt8EeKbyiKMyBVQdCEEDIVhvjwm/jsEN
ZASwANDFlxFxvV6b9BsgcQcia1sC3fDgeM1ZXH8gS787qUsVt729SixtKDuG/oMq
Zn2dlxPqWJFICcE3s5IqA0QJrYBGDIMfM/8BaSe8daKqPMxSFbNDczMlzPOUikt3
GKdkTr8wfsQdE92ySadT+MXVLghmABStreggxtZKZqt9QOD9jxozMsjkuAHl/+RK
kmzy+V3EduQn/Pv8bRKFrqwU9eQXr1inJ1xqqUXjcz9wtjtUYEP62wpdBfeAfIAi
aHPAQW5Zn+L4PMuR54nzNjQuSRMQZg8HYr8kYbP3mJQ9QwzKMtLsnQIix0GsVyHf
k46gSV4PXbIygp0cC9BeN9WMSXtnYUOuVQGF8fDGKXUPiXJwB9NzG2cBvbJ+XxrE
CuLJH59tnWOgsXLlpvrYv+dnK+Ia2/0j0BUVFGstCuL23GzECtFmunSXY31WGk69
AnIMHuLjOPA8IC51eKa/AwBte9GmLAJfzI8TUKpoMy4JrBVxxM5Jy3d9jQh5lvsf
UDcIotlljs2AHWAb+dVEIeJKvoKW/HXQHk+zUHREC1L9Njf+KlCVKAo75dRNkbu8
osvB1pVDTFdf0k9jeVInfhc/v/BnP5+tOrWY8vgC441O9iqnWIfnREtMRNEjGTZs
O0FHIW1IILW5RQj2zeJeL1dl6P5cw9n6sRBbYjHLxaXKTXeWO+yvriRcNJXi6GqD
6UhXYsfypEjrf4nIrW9PXK9sTkZVmSM2dClo0tIfJjEn0yiR4wIiRXmMwaaNsWW4
bjSd6KKJPEOVED47hIvKh5UfzGaznqohRGQ3n3xRV0iBVL56Z3E9b4eon/gffYsf
STTWE4oIg9ggtzBczx1aKVriUt0F6WbVDxAvABsPFvP12CT1o9LADnaRi5tZqqxP
SDcSq3pulK1EnO92264cLctahEgCscJoqn6ZITB8TRSllXThibj/q7lB4lEpQanz
Fs9spNB0H/vnsbyHfHYHaqmHgrKzefxhoCPFMntKnd1Tei7HBAw4NhTOA6A3zaRL
iO5lDk7zNHq/RXMDiPuwxA1LsAxwjdviqs2tR6YmVKhAyM3v/JVtFE2FnZRIGPCF
t0K1hKFreuMocJ+5Xr9IPvAxRwwWqqAmjy7HW582y3jX4azifmdUdPzpzxX22l7O
fI8dd7Esf961sPfdRuMcrSF85tlaNyRCUdl5NiUsdySu9wOyFo5UurisR999RrI+
r3RwjlC9s1ECehmjOD/XfeySiKeuDJH6fNdcfypSQlwxkeX+ZQAv9nx7WCNGPkRg
5XJvGSpu2kN8EwRqLGrHJ1KgWRYEoH9IZcOnaq/Xf7wl0rRRQ/dnId7GLBT0SnVl
8VQB1vVMGXaIzVoOsb8LsIPkv7E9Qxy6gRvukLeFg4qMC8CxlR1MUunV8GQDaocK
zBhVHSpX9MnaKN9Y/3YtP+yoBlMLvbuocDiDbvPT4C8KZwVxiokjkA8/bBzFwH1e
7Me1dq+eyEEWyr11kMkv3oCk2PnLCGPLvSHDEqol/vFIar3iAmijjLLxjyCBj5zY
/NZ+uimIp5v/TT1rP6MPD8XXCMOHCVeYu2cWs6FOsPzBhTtQDWckFJGUWnGR6L2c
ovRaqS6voqjno7Ic4hrKf6/t05pqVtmwA5HzKiAYRgPR5y733HAkM7nrJupsfeD4
QJvSmkKmj0azJOoXhmeOQtTjfyLR8NrWYVK8+Tk6S9VJjQ0kYkls3rkqNCpx29K4
/Ef0O8YgQ29W8hrRWLcCvuhfyEovAiGnEfgf/qJdx0L5IDyh74hWVblZdQMdXYa1
JcVQmi6/PNLzMEzhOI0cIFu+Jx0tl1kYGrimooEBrNaAvE+7PeybGE9zD9NMQYDJ
iOuhq2jQgqzlK+0E3UG64+UsdIQ7kTaSUzTHu9vr4AYXeWfZq17ZyDPYk2lIjCa4
frAPALKQPZ3rl90ghaRSH61L8C/8DjgbQmNm6o4PJUvPz39v7WG6Q7AWPbMQ5B6o
epk65BT3vANUi1lGHPrLuPPrQtd7fG8gQOBtEpz2rHlbbss8Dw4P/+FdgkM/Eekf
84mty4nHAwLhyr/QMZFMsGxzdhyCxIR+BmY74S+PbWYRKnLl/JKmiynozkxit7PY
MlhGEJrpMyRrpPUKhnOVkJPurdTxLPdqquJpRGc2Mb6UP8vREf4TOrt00MxBDNBr
QfwWkR/KiV3J/WOD8psQbKq8eNi2FnsE+kOJRNa61Vkt4/Fib3KfNIJTi1kUheRA
onzsKMBV3lwsg6HoxjCdxmUx21UW51M8zdDWjmXM+0/PPoqIs9QPOqeBKZtZu0cC
t9Q0rs32JvBEazRXdGHgjp0NQC2QqNIFvtfgU88t/bA1YwwIsmuDvBRSZNQOEr8d
IzWD9D5Si/VNJUX71lATsL+NFzLAU0q5XmPMTOznpHlxs8rdkDSm8jacwDwlNrSU
asDfOAoqvbuVWoevwBP2SKj2TCwG2B22wRzDtVdDDeyHGXJtN/bnFW2FacBPLgyI
hqVrPFTpUJW8zZen3kUqdcafHwJecl3FBpQGoOydyX/QXszGEaNIR2fCgUAtXQ9z
lBXM/d9VXBL9Iw76bn7Z43iUVNwIWI9QTM5sQi8EMaaRoDaibgtJIHWK5z8eU4nh
DeChJYeaLR2Ni63p0ivIQpbnBzLCBG9TF+/6FAD6SiokCh/3Q6F0E16pZyYt++2f
MucK6E9OjeAYedPzt8kNtkb6EgEL6dKI61EHNApLpgQEoyK0ITl921PJ26ocOZhu
M8r7GiYO8+6k7ctDPTD0S0MZkZijixEx3QWfEjWFV6OpoYM0G3Nv/T+BGYhKAeUV
gf5e7Jc3mvPWysgFPaQHf/CsMQAIA9u/48/nZbPu0abQkizo+wPEIVq9pmAhyhH0
fp52qIOr/jjQq+3Xu+HoB/arR/nWHQ8x35KjESTPZvoYkrs5bcmFf+i4aPkfDUdv
Eam+DITI+izkI3kIoZPl6fMO7BUAIZIG9rX12dA9MiV8susddRNMXtsvftxNCuZc
MgwnU6px+akrlm2CGiLmJUW4CZQY5dntCY2A00F3B7gsC5Th8YeBx1XKH0MU8KXf
4Clqugn14621o65ndxSWgoLGMnwVCy70Tn7yCICFZMvNdSKm4ciwcZhydjmCcvGg
7MC+JEvKqtVoC5uzp+SwboSLIx+4mIJviOFaWaBHR6qJBNub19LnQ8mgsSxfH18E
2tA+DodiWq0jdIrabcG/lLY5kKnKXP5KocFte0rrknneou4cH/nYf7yO9TG1OKJ/
IQf4WB3I+uIcNxsPTtBfwZK/nfEQXDCOYjXQs1ZevJEpN8zF9+1EcMOHCBOT39to
d+6ax+kXf/E5QgxVXdFrIgqwXMQHwaarUYPQNagMxumjtx9WuWMq5D8tzXNW38R1
DKvJkLtyMVo5wobpypDbWdyx1OSB+hrjDwWV15WFW13p2ZukVgFNLhyEUmFH+fdY
FKQ2RdJRDv0qeX8HN9KqRwafjtlKqN6FhtUpbiL1qVJUniQpZbXxa6AikUBkOKb3
kMhCsQVuZvavLFsVfNLqOTiZt+7UYin1M7QfzLYpT7czzvDSceudvNP04jfLwz3F
294mihfodWFhBTpAzonjIxyzw2DsLLp9f5s59kvnYdRLs5sreXwoyJqU4f6uAzKo
D6UAFADGXnuk2Cjkn/3Iwk5Z5sMnYqlL/oJsHj4k7Bf2gBkZUD70qzZDH/X6i31R
qzv5R6ncMLfD7nqT0jxcNzKNwYBXPE9cgc2ZUwo3mmABuZDWor11IyT+0WEb2Xt5
zSwqzzmHHMEG9Xy2mVPPuVzp9dpdN9M4JSCuS9QGMXRKaRtSaJMqy8QRCb2SYX/y
Z3SkEFcGypjk/eRpj6tAT/36ZD3R3ZrxRQEqSLXVms9BlWHZGqz2J0O29eZocNW6
YlYOItrJy+2nv7IL6K5y1LZJH/GybJQOCrfIZq1uh0GLCuWO1CxXsji5UTAZy9f7
WowPSdhz1OeiDH7yUh2cWQ97stgoXQE/oF5JCqqkntF5bVx5PXfHgpLuJhnVKKBx
36/PbRhcmwM70VSCt+cvg6UxiFAkbMsqRsC6DsGXzhebCaswS6YZTElt9BlGTGiO
lxRc1hLlzSJhIX5XLSUnKPAWmanMSKLkB3dEsTmZwbOEYaFTQq1kiUz7E12LbNlt
XGqc5ZNhBYFjscsYVR/ZVgjg07x8R9cl0QdW8QMomJv6i29h5ugYM5VYA/dHpq4e
Zp93WzJfnxna9f9QFJDI4ReSdGl9W6t4fC0og94Qa4bTZVuCApwXNZiwXV2iTnHP
W7UE0tACaZoU9+YyZqHkHfk+iJEUy1GKA/2NT1XG2IIhpoEbzPJuiQe8sON179CU
9DXaPJ5xN3eUHuc+/NFkeh1dpwGZuJgmDYVs1KKstSF8UnlwiCJfXRuOLud1WLt9
Xgaw7g2RQPH3sb+TGMKfQQX8yf2BHiTjVmJzcLg5xBBHv44wv9rJLqZaiYSd6E/U
uvK2qsW4+KF7BpOJD7GSk5vpPyR5ipUn0RvqEYXY7bmCpPbHfNKUTz3ZRbitsl2F
g7rehRnAgnVvb37LvXaWkE7w0gd4I8tUlldPgkgrVTcLzDJaU3v5mfzxwhGG/+mm
8OV+HtiHXStKEydwwV1E0tM4aWuOTWKSCLWdEc1HH3vb1oKBHCx1kh9LS0H2516t
hZb2H5VzSRjAULwaVAjH/vyJYm/Z2ZYF/oVlXmpHKVF+Dw7HoKkU4GoS7wXbDrgl
ZDbcJu5+p5AZAidBXvflO4d1tArTp0fmxCQPFZyVrzek+hH8ehC6NgRAxlIu5rWW
SwshsNuDfxiFe066eHAOUWCSgZdaPlWBcetQR+GBO0ojVO00OyeR55+07pTM26LT
hMTiPBctb+gdyhyRmLhb9tUhVrzqyUkumaI1v5b7nV5yL1KiT6e1IeL3tQzogh3g
j9gT/3HViraDXiDZ2DC4TuIPXrToSSQ0vKcCkryYjQyIUNIbKO7RimqU/ag2gTfN
l3AAxyCdE29i3f0hAkdSDQXJnArawlhBvf6QY1rYJMNTT6ul6ZHxLHKjFe+3R8pF
1z2rw1r1G0DSU2lI3bPoIpTeL04ep8gWleObrPhsSiePaXFrYMlu44/ZJ4iEJnKH
bL6MBdpVpIwyfLNs+b2lKs345u++4jztZ7+NH6HfELSvwWhWtCYwrkiAiwKj+TVs
LEG0diwdUKEU3lS6P7GEzB2tOehKZ5HJ90VIh/zo0Lk8AJ9fn6cAARCu4ewF6EiH
B6nGU3gFQ4UTBmIdO1AGqI6T4lQwrzrD7q4fqKuQS++Mto5ttO6ujSAlMYHf3ja2
afCP4NxKq/4w3S3b2MwPHwchYQgBgl/+C+1D+bqUQzI2VOYAD8mCeDlpi63/l6ZC
Li2rMVZVUCs/6mnC4qh9MmjKvI0oLLHesNMe1EVJJvZmbDRVTpPybX6mVGlsyt+X
lCIxd/qfZpBO1UEKoCyTtbK2ARZTn6fuvghJD5zUboID3gnXSOlBSsAwZHBoCj9F
lft7rO757KBrhNk5FLw3Zknzc8lXTiSoNgqqOirrthyp/OCYAMhEq1J/6oN6n/D9
OyLkX5We0C8Ea0Ogo84fxSsfHxIdWuj3fXNvrm9dpSVxRQvW6lTQJ+1IyWPcUZ/K
Mii/7TKABS6B1ElER5vwQnPlhVwRRrEQXKglL5wlLtoOOSdt7/37/uxNKCgWgdKN
X9lCbHVSkvGzLJRPHQ+kmVYH1jUdG5BGOR7nbxJ07ztOpLPUjlMyebixds9bdeXU
kGeo/82EL2juqIHegJLg/mqHH7ZX5wafEQ3fMyHZB43kqJOx6SzHxuivFCLpB15t
/kpDJ468NYAz+FdqJHfedvkwNfgHCJIcN/5wdJxRezZ+2D5p9jQsE8VSAg2up7oz
BQTyI1gcny2XG4zwUOJ7l3Ril+UK/eEGZn39OmGrycMDd9vPxW68xIO/PiIhYieJ
lsVpDOK6QYtDqJs1egZS/Qx8R+WXfiPo4nNUKQXB7sOC+MjjNbGYvBLi525bteTM
DSHo0Ao3WJRbllCQmIAXR7nMaeXWeVSsshbOhJyO+NVBQ5Zjlr8OWbv1IUxEK73c
IXZJc3QJXRyEN3CMoNCCD4vk4tgZfGCC07MFVjEQs6vTbGQJflzySBrpzB1bkmd/
p0DFR4WAFuK4K5T7qewlhRQGz14nvgIaMZ0FrqvkEi5osvlY0N0QwB0e4SQ1WeGD
LoJU76C9LiGvf7UIsg2mxQB2yHtHkv2wMPocJl23sB6+FPxrtjt7Q38BppghMIim
E2yqrGLgh20o6cFjIMAtF0GP1h55az2Yw5g5p5zyZ6eRXKTeuZhX0DyzfPVxpQ2c
AKQ8zDzCOEHVKNBCfbEJysU1rVrOiJCxh3zlkF9Ux9enttx1Ob/uwL79IeirR87E
RZMjosqdCSkb+hZQnZBEsYeO3WekbVivo6zApNqA6TqP9Mq/kIb1WEJxzKlh2Z1C
k0HWdokAEtlLXABnbNSxswa8fR9tIvaFggzI1Qxs8XHDpg6JWWq5C9mWpB/VL3C+
mO1TQqXtCqN2rKuPNgIL0el13BwuaqTgARUKOoJqPvszj1n8rae8JnohFX5rqX0N
v0oxr5ybY7yIZb4TQc4yDm4E5nt72UiGfvo7TGWcLKwgwzzZeLUrgNo0vNkR2dJw
ybtquekJICRcsmw8yKpiHTXbFHQBRybae8yiS9E5Edb1Eun6piGLE1rGwswcgsUD
bXYbbSYCZEbHuAkWSYePA9TRmfE7ro0rxv7TxRlCP5zIizYBBqEGD5QYPpO/M/ik
xBnnkyDzwAs2EShzLq85lBjdQYtzwBxrMyvNUeeiYbUZhjwi/HnvyE59adWhbrMX
tDEhKX9/8s447/LeX+rUZF3h+gNPaO8k4W8C1yWJKwaFz1fffDJlGQcJO1vCfLu1
57dyvfPI+y57Jw+jO+BcRqSg1up7rPpns+fh/htav6X2gs/nxj3H+3/yPKepXD5V
ydO/rVBf6+qDywXCbEXnDyUPb1sSiRPwP/kcWNAoSRGMqiuvGIH7+jNMLPyMbcxk
IPGfzVzPkDpFkiMqSUzu1alKuGhXfjy1HnhgN2jfEwFmtXfW1X7EM6FkCoceTvbo
y+8C4FFFd7Q/F7SFG8AyKmGBBuz3N3fUd4G0rBVXTYO5x2zZJW3PZNPJssVuruFQ
qZ91TrbfanRmjj/8cQsbD+JCrWQJwEn+YUIdSfTMPaFKy3ifjqHAF3NwtrGPQ0I/
6r6IW7+vEkfFFNaGwDWv+1/Y9k/2EIcP7PohWi8CdOPbXuAtpiJCyJoPpco6Geai
YWMwyV1606moMfeJLZAPilW4eB4av0eY6dcCrzsxBNxvFlxJQOygP5lD38zIUwIi
dvt6hWAYTCf8TMz2zl0isJdYIX9Oar6DsF2goTkBT18QfctcHVB1R3bvkITHnM9b
UsYWb9RHJW5Rer0yO5ADV7UpfX9PeOH4a/0jmhQ12sxluJNbAVQ/2LS3OKKqKevq
bLSJIIQ6865xIryUf1oJCJ2NOyOgWlPLRFOAm5+IYHTTxvTC22q88yXiQ5M0x5oh
tmoNvDBP/1A1QUE8FWrJQQ7xrrgCk+B5C4RdIm2lR6PQGWZWYRJUf2ah9qYPjUsm
EYxhdZkcTVw1/nAlWe3XcLdVIezxHJhjI+3hh+0D1tS1ghIg3Ug/Yyg1V4FcQZjf
kQ7DRt3f0+8RGgFR5+DKqJT/qN/eDvzpfFp8W9Ka78xOVIOVpQWpOPaMq74/rr/N
+WoyvA41Mg1aUEXzJwA4SFpsrEy94WQmgLt9CXWzeJyAChxpu/T8fK5TN+EDrm3y
e0QQnKd67SIJgbpDpdymMCRT6kPLv59mvg0hv1HIVE15/G980QYvura2Fpgm5maj
rbF0JukpKhgcf/DHLlgalneJtq0mcT+tFi7v5xYdp8xhr6NWGlmTEfKaCU72SfbZ
n0Arj8NqQwL333FK+N5rE/DFSpsdfsxb8KG76XSKBDctp9YpCZd4HgLLfYZED79k
XBwtjpbzCotNx+ILuj9hBim5m1xEXaNlMn2m5MnmF12LXZdlmPJSSv8xFiV6pPfc
mK2XFaDmmw/3FrFs8IEPEuO5iFlhWszg8FyFbqUL/iY8kpdjuawNCIxVMY5jOxPq
nAzSoGGyrIV3I+0kgrd2LixdBpVTZHx0NHVOAiTtJ2GML0cDvCPw9KBmg1NGSmy3
Oa7K2gexFYY2mWzUnXki2hH5tZhUY+XeU5+r+VdGTpPFqlmCUlICgkMro7ZUx+eF
dONVstRNDY8sXbdjXptoG5FVzbPgnFL9z3OERXT4DYe+PiyC+obwm70M/4ZBakPd
/1l/bgbM6EmeXmYNynqwB5EAA29vs1UYPecQPNx8SKxGlWFuYIU6jpqp7SuRRztO
w7HLjRD1dG1X5Z5EbjJOZtc3BnzVnmyQQkDbOsHW9XY0dBgC9iDqlCgXYKstdWQ/
C2IO8LxL4Z+lXc50nWYzzrEP1P0zboPc4cDumwzaI+MxJ3GZY8K/JPkqDoDPsHo8
UVGl7PdcAIsQT1tdQOUyBnnDaMV9TvghcUBhxlapW+DET9qu5qKpIZc6kOnf1y3J
+lq7lh7HR9v4OaijARfQHVGKwmioawb2Ad4rJfYgqviMgeq2AB2aW1nWaTPkyruW
IzaOb6tpJ0G6xTSD29tE+lNDzMdy8DtABbekt/9/ghOV2hY4zE7fdW0ON/IRs20r
RZdru9HSMaYtp9tTRphIufB6kV4pB9ysr2JJ0Ngv7tgMveLnOGS4NKHeJqIVdnrm
UPfg9SwD1vCWEGhqsw6fGDB0cX5TtIM0Yssbg73CeW3Use5BD2NzZI7GfiJeX2xN
LgTcuttJQTn2K1CtxmRUkG4qOtqGrRnc19mnnoODuf1RxBvL2uMCIbZoGcMMEryd
X7+BRdj6PG89IIHXzKLVG0D8u6bWjC4cXhj3EFxfKvKqBHuKFyWxcJl8z9lYaHLi
7fYP4lhM+vejXdhv7/R0V0PV801B/MVDObJmyNyW3NjivVEscxpLiQfVxMLJrDQw
GP/qa153C5kkWUxwPefNHgzoO3XjC78Snuueq1y75wOWmzuSYrPJ4F0sNlhMQy1R
L7cu5srGpZ2Dwu7Q2n/0D8yd9JR17zOPyIlngizec0kjmy+719n8f7yBjQ3Bkii8
vf+TLQn4gwyyNz2/x5F4b8IUwIO0nKI9If/AxmXSw8cSzhgNn54CrikrHUtORNox
pCtNtDMvsRsoK0YeMlbotJ7g/Y02Kkoo1M6ebkRZlZUg0zTTkpB5EFovRAf5/9SG
5Hxbg4q+FPm32S7u0ruQPMUZw0Edf5oo8sjHp/rDHeH4mTG5wvIoDZ+1KIASAmoj
20W6l+vBNxrrJD1g5mw7OFkykZiLK8eVwkCXHV5+Q1+9V2Q6VbadE9yeZfSTVaXM
65yVM9v7Oqwwnd8FFbludq1lFmBRdtdTz3Y3dUOPSvNNVXrRD4+wd5ACOITbVOIu
R8PEi5YczjftV6L4DaMfbQsIrxt8XVEAZ9G7a23ieFHMgUJkOTA5VCW3bJXyGnbz
mVgo8sH8zY5eLzGB+CsH9uFPrlqHndzpzYlk+qLmOdunMXnomUoUssrFFvlqXr+/
tlHjq9/bBzgnXbW0NOTKxcXrLTXISE7CEN9h3GOazfUVw3eDy989ySZPUImRF40I
hydQCECcGA8zYe8uegB56Jhi62ekS/JEW0/8IOMavzTbNlANg0YIlGVxfY6m8eBY
UxNsEC8325D+aghJyV2T2QAFPHSnAo/Nla6KmnKXTdfY83W6ISyid0XgfZTgfweY
9Ftb2f1B2FpWCKwEFHt+oyXxIpjLbAJh9XF5Zu0ULaswAIiSpdoPa0OkL8ZICiPy
b/rpGK7qvHufH5D73i6f2TrpPKPLYvsNuZZv+bTuixkecgzrrg+r2UIJ9dvoX9lz
HcOOV4c/F0FTvRwWyCGwoZEV7VO3bQGd7/Pa3RzExMB8VUsVWqWpb3FAilDCTZbr
8yukJEKmSBeWPbBgoPq17UIES5o7oZyT4Gwa5FK1Q23mIh0GtCQm2vf9UFM7LWlW
8lqLY4Qm4HeIpH0VJdxOiGAEOYNvki2PMjCyt9uVLpjhCa5SzBIL/VM+StixcPJl
jko7kT45VvBZci4H64pWFqfN58eALhh++yfeyQxkHNhRVJiYjrBQiXj4IGtmK1gT
X1r2UnwEnALG5mqFq203SJupT3NQ6dE/R806w7cE96ELF7OcXkRfAt/sCX1W19w5
h4BsgMFVhFoKIiQ2uDLYcNHSVz7tFUXUhxM87gqXmdVFoVD9vLLe7baLX5lEdsys
NJptXFLIlMuI70Nhl+MbOA6JiBoThmhgFonFrw9+Cgs8FsZZUmvsNZu9s/yOzF3v
Bok9wcYEp9Ux2a430Y5jjl6xqtGX1XlYmhPWX3E17kbcJk0NLC4dGUJh61VOzbCC
cdJ7oR+3Jn7ys8AncM+sdH+CB6nb1ALjFtZlmXfcUJZ0ODyj6XpgJGUNLAaqVzL0
LUHuN/Ab3Sz0qQwTYsrjYAFtA0F8Z96iwdZ2MRPkWivFuix7r4pedfspOk8xe2fL
+WYlhf8hKOc+Wdm00DTk/REIOqL0X0Vug422F/Eo/eZ1UF1tpAyK4l+570vD0M+5
vjJ4dFRkINjDvf1v4ZClfv7T+6hfRxldwxcKUTKKeuEParqtsMqOxIBO5ZuoPFFS
ovDBxv2iCU+QUxtAyDXnuc5i2UUg46r7kc0O+t73VMqM6fEeOMcDFmNHGQ9hojAU
pRMowWEj1qZ81SpBs7ntxkOBCOwuJXOAmYZyZz+lT9W60A0N6pKZeEjmEhxXWG+j
75HjxrRvvP5mjOQAgHJydxWXRrXsswpqNepzXCKRzRQ2eqWOEExBYwUakNnM38qw
V1FLOoFpRXfvY7nntCL656aE7m0Rvl3fzrko44LEZj18eeWlHbejirglzKv/yMTl
03W1MegHM3K4ObhTPjXOfTxdhoiqCJjqzCLfdFFU/WyboAWHj1UvJzudfAwCKUwl
0bJMTRBDlJ1QdGS2uPufyX4abeQr0iPqjKWwdrVk49kgz5YUYp421PSKM3HNbdIq
sS2LmrbxAfKSuHbJjI4REDwol5MEAnt0MTcTQgtVAj4iJBSOIOw0ybF3ILvik05X
jSbANd2ec5fa9TwrzCS2+UC+4DkLzqzmCSIIhMh6N6dhvSp83AihDUMry0apOY7l
vL5SsgNhG7Mm36woYzgpYW9p6tEt8rxuyXyhmwb2t50+6fdM5GCkFA3+cgpkZeua
a7443dmmuKQYZczlTyyjNFJSc2vka0Tk7TwF25ngg5NGTp0fKFCAE0XDZuN0OOTY
RsXhrmOC0VuW2Tp3rE909RfR8kU2kJNTKHFxZgOCKFqzkEaulMAEBVBOGGkOmvAY
42ci20VmyoO7eZBHc7e4ZW00bbk1bO7wzCIYW9+jTQSVY51RfVYMeKjzPIN39gYZ
mH9UwpuBy73VTGpCkv+Pqq8mWN2vhNmZj47X3GkW3W1L8q59dt9eRCkzdgekohi3
oMDcMOChonVjbzVDakPvtmazlrT0/2jVwwFt2Eri3VE7i3IqVG0SkFVP3k1su0fC
wFVqKybLjyl+tImz5TTyWiAB4B2OJ2+r//Jq5Z+IPPGU4j9jnDPYWIJScomH8/cA
1p/cc4LOF1YpKP9YAJcBtLv775JGPMy1jpf6MGawzu7N7xgFcCTdlDEnVN3g9rwV
0rWU0yzjrjwpzkgpYvgOZIOsnc9s2xuzu3zK6erNDQUv/IWyHELNYSBEF6Qaqq5g
metAkILfy/B8TPzBpkjGIUGzAZPufiH9g4uNBUpSEKEf7oVI/sRQCSd90dnlaJQ1
a7X3nyA077saGwCnNjF3lDDRw3+rQbpi2MkvTqFWLnjVjOubxCrSdvmhR8y+6bfn
mPcTdTQjkormF1Nivxt5YzGqyOvPy88AYzlkmHyhZK3Fqo8CBELy37dlKC/e5yFM
kTvsi5axf/4DUYaDDE18TdXU2nZEBZ1hbb3jlE2Uco7UXOvAwJNw0FockhR6pxZP
FdTC7oJkg3/s/uuJOy+4FdwFyqBunUneusDO1eHq0S2jkRrcl0Yd1rM47NfqJBRX
kQ6a6+JTnfEevQvxzeTpz6JzHi/rCtlXMjio4WubHY4lJzUPqD6uBtt6BhD6P9qk
+dpaj1tt8hN+ZWlcZScR7YCg9aOg2GjzA5T9SJKPMtjp8t5SEZ5TLFFciThw772a
iEInWKcUhuasdOGnGepXcaBdOc5ynNgVdoogBsMlRxFppbiCfIRSEtq03007gxK4
Csl8WHhT6yrs63VJDxj8C1E/7YazH+XcXKH374q77jy2irAqsrGyzkXaimdsP/4p
iHQCc+JYaK4IGVrHkW9FhGploYG21/1BFp4xDgD2XfVZm03YQ+Py0VzriLZKtKl8
0QEjnelLazGYAhkkkv9qA4mI6DecOCEXrRV9D/PPhYFD70m1eFFmYryG9c8QhH38
M1vc3fCrSlg+flS+fWnCxmed7DXweCtmWBUIxLwG1b/0q0nOrgAyk3bkUC+VZw9h
tVkr81BQc3rRkzsU0s0EZurGiLZhapYErNcDMmgID4tQIsayRlfuztuVmqCXFuDF
KQ1TAzNbofhFmDid0H3/9Mti5p4NrhCwsXwn3bTn6ry0Cow8QrBg857ZbR9bM5Di
0e408CDi3ApPi7AE4QUCPws6MsIKQIm7SC7oQxOhsq+HeX77/8khh3lsJIBQ+y8T
dn1PvOPhmT2Yw1UoiPZOLHcVfg33P7qsTyNIgGqu4ZZ/0eE3zic85+gxLHLhjVzW
TFRcjqwJZKK8Wcq7JboDSMvaQRu0DFq9IHEW0O51hyK0fZXWdm4IAdGRFfy6paVx
pbjALZNaudsvvRzS/l5CFMF0eq7+L+eBw20P3i9idsJ1W8KGCoN/f1pVdR+ziUWV
q57enke1489uwjV5l7CQ51siZ+FlUzlN3FZE9w1A1E1g3X4WgvsgdOOpKEz+0GEC
/zghR64w1q/c1vESnmiM0FyTPJSzo7Y8M6csUSrL6JVXB5CY/lK1ROZ8tAaJGgkX
dqsbQ15GD2BC4PeTQuINmgYwIjDp0EkWjvrn5lQcbTT9G2vN+ZCY5ui4er0dA9v0
GWGHkEsFASSLkR+zPYrtGMOPeN3RBKVugUskFihlk6loIp9DAGS6J8dT5mMPFiVX
65yLdmD2wRcmAs0Ty/gGrlAj2KAXPKc1Xwf77roQDk9X/JRLKl2e2eMQYePy3Cnc
oRI8hvyyanxGlxA6mTJzEZoaMJaqZGJtdUI7iZlDqE1J0JQzPbiagaaxcmsh0+pp
TM3I1yx870nx/yxz3BB72O/M2yNaumlNZNc0ulyH1rBl4CYNNHdY9GXc1J0lob9a
AR5DuozLA4qT+5Zd4ZtFjCAFtU+kYbHk3+u8iyzqyFnxiJVVnyUl5eMKoqO4ESP2
0/Ipezag7eLhokaX7ceRo6AttE12IkmJNtQHeLpjXGzOJFZt8is9zjhoz5ALW+Pn
z1jC6dui8+cG5m+mIR5fkvgKaAmJVQhEYK1d6LxM/FFt5q+WuazWgTqBlVJoN7wt
sxBYBS/QqOpe+xfWh+LCYI5U8/nPa2FzT2zGxstBV6JzWOXZnIM+2in6yDMTvRwh
PRtog+znI2y3zNDcGRDmMjn8cqyMKD99vL8FS7dOCgnklugztNs0wPQUUMtXLRk7
Dxz2Gi9Whg1m8B037w9szvgsWXhpBUDjP5ac9QB/2q5LqnurEwlSE1uLle71wAR1
QTniaolKFFkFWWOL57jZMthAx8+E4072lErUrFkp+BK+fSgzOLqtSX2gdBz0j7Fa
EIxJf6sAmDE50UGpLNhVipe4iviBMW3wXsx78qRPqopOIFawcDxX4KeR+KjmPn1C
BUq3OF5PkHfhQV5XxvU5aMqQczgwVX4FAKx4db+94as69YOBwmLZ6Mynrd+Smoop
N4czFGxiLxJsHKo/J/cl6LyleksjDdJmf6EwU9NrrTrQqHCdbLu+1JaxwUU26JDQ
wGURGsUmPXgGrpciK7olGMs8Zq8M645y9FkwWJ/RgepYlEupL8XZ6jjBcuTUHgsc
n2xyQq/ZC2GaX4PAJrzKQX5QpAniGcCL6LtcnMRSG9x9AZCS62Se9MTTGiAU3jo3
naGyj+gQcwzpdqqXJ3Lyh7sxc2wryduY1Ovx5YVxz6e5ZF43ojepDgpDHi7BuPA8
ZS/t0oC9UAqpapWCJWJdMA6+tGgA24evwinYB48PNOFrw+SVI0yVpXFp7kCo5YwL
zhffrHzbn97g7W0E6cQC91uD1AJy7I8ILn1FmyB0EaWU13kQf1NzGJn/f4qP6Nnf
Jxs3lCfrUDnmaLHYxI+Arl6nQpo3G2ycYA2lpw7C6uXZlxZunUEhx5xvRslW8grB
nbPfwi2vgv3wbDbcHobmNevus9imRdy+QcuiyfqeLfOApN5aRuXdCPcI0OLfyvGx
Z4sno3Ev++MVmxpvAYI6us0Gs11izSZNu1Liv7u2YmB3eKbBpgo6qa9HDceXKnoq
+EPkY8BI5DnmQbubqC8DZJ0Uw4d8V67j9EMd/pqaQxRn4EuYldY2KQ7nKZR5kd0N
Obw+Mbfyfw1GiBxMr/YIEzRnrdrtaNBcAfcf+vbwRK/mGEPSA1y5OSWl/jkiHupm
O68rXDFsFRJDKUhl9atiULa3jpn0cyR0hjzRPM9cohkvS/tUiR5jZpk8hFCYBY7W
1BkNqgWB+JVNmZu5PP3FvGcKy6EAezDvPKyIKockodpef1AjA/PozzcA1AWVaLj0
vNgSYsFRH/r8Y2q9FoEkd3XDJ9tIMlRQK3d8H55Svg6jTvB0HGKqpFf04i9+WPT6
m5V3LTo+02yagcm5AwDXgYfCk42NfwB9qZbLdmyWwW7/0GjlXOjGGDKJE0vxCxsC
2DEvwIGDiaXa+UJEuaPu9LrXlLwUexCruPq88PURefZ/0ECwo0G1dwFpV7TUeWbP
qOHSxXAINVCqjGKf8T3uODuq9obzf/czC1B6jGxIibmZsOCV24ICjhilzlhgOIt2
ISCZRr/V8HGes/StGqGjUbmneICFH1AO5hau/nFiTWh0s9f6h6bCw+ieUKUNQisI
d8xAb+C9/Bd3VU7Me6fdToLc4wZPy/ksbwCs2hKwf55639rMpEPuZUz8HKBPnMLW
691GvyoIuMaSfAapNXOdR7QngOBrd8y/vH5Zc6q+yQYztCwWujtuIy1IC6TbAaF5
lq1AureCFKXNFMgb5/eb43OB3r8Hu1u3B987WNAiTCYOGXRVPlcq22ATCO8sxx1r
b2r9Kawz+jcGvJW0qTckY/Zq+L6/VSrPQNVc4hOQEEBpEhsYOmm6d+MTJLjCpc+N
Suwg15TMI4R6l0lYS6WItdKcCdU+g2ZS3gAMxXQC8jNTT7J6bidx0O6p8vRQ/VRB
Hzl0GRZsvQio/uU05PzaaVME5dr6cMt+ZyxGT3nC+9lYE2TAP5Gq2tOT7TBl4Pw5
9Em+bf0i8rU53HhA9pQlQ/KXudZ9WW+cxioB4gBgWhnqfVw4zqVLIYJa90l5bWZ5
KwToKAp9ejFrKMYLBcgtKDdWgMYV1ZNpkEsdn7h/9OOCm7dDtfr0EQc4SuHDDpqf
0nNrqrO13S7qtzt9oogvovvQKiPflmzXCEjClp4sbi3HzfG/z0vdYP32TkgZZVjb
3Cs/Sf8m8lE5q0/autBzW20lzupXMb9JKlhWFJcFQldjxR4Z3zxgOXfGBPdy4t+G
ohgPKd9hBfW8oJtBOItQYcBZojla/OOVWuwokFYgCG48vghqCBoEdm0WwFmVdxuc
/yzqJE1OgAExwV4dXClimPVnwsP5bjnEIlfHYrUIRJqxl3VIfYviobIBFmTx9Syp
fLvzfYEiLjxf5/rY4ScSRNoybkr8JZJlZJTpAhRow5ToJMCFGLLP1gUwMiNzzasa
TWnyqNuzWdICmXKvPdcjOm7PZEPR0irkt9ldCakrY1DT23jrXA7JNEAxNhUjRnYd
ZmqUAqtHRT/2lAiv3D6BP+1OjOMdaSMF4W2Kyx4dNteUhiA33CgzDtcH90BorMOK
kiVh44dnPeUI8FD4C9lNriuGkIQ+4wiaXl3M85cp9sz5JVcL+hkg4zH7tdYBv9KX
yYK66b0VgYhxesM//b47dotNYZ0e4LN2QeArBSlYHfrAXnOlFvcG3SHbsX482bP7
+ReUYW0n2VqEvdO60HvISfQnWColQXwj2oyAEDc5P36rj2BiljUNSEs2CxKqNiNQ
aXyrCvBuzFQtgczgVivHX/Z6vmOz7EDvrPwZHULstMiRHBbk1aH5N8dveGtH7e5T
vGZ9zbPm2EU5+PUZ3NA+lxtdVT6ZmMABzrQb4jqUrO8bmlB4rqbsu29O/Um1Fn04
k2W1ERd6pIq5GwdScwsDMYu1m0hDI6A04D7SFoNZCLiqB9SHkncnHH0T6G9odHxb
YIkwglrRoRDAoZLE9fvN8ChnNBgpPWHUstMjVc9pi0MA5jZhvimt/wfYkSZc1+05
Fk44ry8ccYXeAxxYeyQJSqD0JmvntFU/NmsfRJCDTlqS5arTQtxUwhEpc2g9QhmG
0CP6xJ9dnWCw3UB825LgtapA4kbk7MDjXXgSE7dF/fYn8DlMg+B54Rtmq5FameXM
qXkYMIvrvXcNvs5gk4qlT9uqnsAmson2osC8GyiKqwTnXV4wlushsh0elUdrgShp
bG+3drC2d/cCmfYl8CeK0Y1z+fiIE0zVOF+M7SwGrhgPien78y9Bw9AP95aO0YU8
8Zsh6npL7XFmPs7HoBzmxM5k5N5OXaHzV2+zvJIpexAoTWCBY4XiVt9rUZ/4rSx5
ZPisdluhrOojWU6TMsq19MeFa/VVhWTqzGX30fNbVWIKXq+5lYbD77kF5TW2mYbJ
zyDE0xHGa0xIBwy6HSgBBw2jrGMgNrwI0s1v3FzsVdEtILrFF6TRW/vGOHdEsWGC
UFOGo3HaB04m34TgNZBwBBauT19YohcrmGRCj5XRx/MvAE06cJyEMGGyC+wq8YWx
c1I0iSiomYEH6+H4LeEfpVacD2TBkbjoHtwbxeBGwLKjqaUTE+w83E2X/cbdDm4X
GuQYs7yFep0VUlEGs+Ht97/CWSR2VUNw9ToV9jhTWVpOjtMts4mle1b3GzyAohIG
u/IDcdiVyiGPa63GsUQtWfxOON9LN0q0g22eGzb/4JSKxtCldBU6n/MgO3iC+MWG
55xooUglECzDfgxrfxLAQJ+p0fMl8BO/yPPYKxWIiYprmDdA83Rj9z2NPp+PB2nI
RZ5P8+OA+lEfsGJWYhOxlf+4ZGA3mUbcfohC8Gq92mStgHeHJWUqUmlLYySlh57M
LszVXBwr1qipDCc0dQpZnPbPHrf02l7RLaP5aSFp9m5sEzF+PQL7FJfGZh5ylJK1
AzAMwRmsUDPKsVc2YGRI4PKz8rUknGUsfWDm4iFtGv0Zi8BYLan5gH5SVgPUEhXk
1qQMNL5N4+lcljIMmTGcSfrfUH1c4XFPlM6pg3h5f0cuCOU6HipaVeusUKuvNR5Y
zW/kDgVdh6mi1iP1Os6puP8Sbw1Nayc8JhViGftcki8R4R0zhk056ELCn2gspPj5
eBXFUuC7uYI6X8FzSouUFR0wOfgSeCi+69pwdxryLgB/oQrnTi89PaGY9bd0lqp5
rNvWqthe7bX1ZoAer0qbFmWdMBnVR1sgD6NVFWR1C0zpTypalXAFvObiEuTrHyHq
qz6SWLbdPNoBL41Jgg9WYYvV1hU5xe1KFPzlsyruoV3w6zR1Gr3wuK32OXtmdzex
vAnWjxnJV1ANS85RRNyAKO45cgp0+tqxdgT5O+bBVLYWt0BeWVZlx/tW6zU7Giqo
hg6guFZYQ9+7RqTdUocCKzQnc4bDeTGJOHXPkRItROuYF5WYPCGDIy3D/Z/ACD4d
xKcLdJ65rQfkUYxAAN/2E0XPgvEGWNPe0mTjfQfL7rgiYwUPfVLV0eLOAeJq3qNS
15IdXOjixuAZa3bIDVCAmyv++D+OFNdcEnj94dj8goGjZm3EJCZOpdvgDlWZJNhN
D6dW6LRPKLn781/G4P8q2HesdV1gKaG+1fQPC0ZlUJy/bYfz36KFu3sELsSXy8t2
Y+36S3aLkieJOmWK/sj79q58GQ6k3vN8L2qvE2BxcOqWKzz5vpEbAGseqltalcus
Z8ag/G34k7Ty7GYOa7aavb5AKBSz49kkmuSG7GZIUR2sjjUPuhhhysZIk8Hpv+D6
HtrQOirFQR8TU6Z4RDZ0lJGfHCX5Wxs9b83t1AidDq68fsxfD8IMX9Nfw2BxpK5O
+pdRGbZzsl+UuzcGHMoeaDiaAYNbFy17jzTdVHJXbUD0blieAmQqZE1XG+psoK62
krVtUi23YBiA3DGf1erzG+93mj5gYLQ+TD7ptPFSpOXj6ZFspTWwxWykM0XBgLa4
izDB6r0dUNGTu1tsh6XgyYLKTcD34gZIzvDMv6v1lx7xDmF2ud/KGo2nDESoP8et
geKw1LIBmOtAUMqQqB6OIsuBEehu2M80HNY9d+CfRxHmb9C0a2S+rCBJAYB3lTif
2QgUspAlMbP8NzYY7tHjGmItFE1OgwQ4KAjAsb7j1a6WxM9q9drhKGqqM2FmQcKh
qxKf80ryHtdA3cMZGdg7FTFDv/6UZrriCX29p4Ptvjxq9dEajAgeKlvqQa/4aE9j
Z6h16FfC+Fwv6P0vLJOC0sjp0X9AC7TaY84ywj2+CVbks4cf7ydDUdGQ4pfpAoSm
35coRP9VJeQ//uaJ4sxzhDDk5D+DEWB1eNTEr2Z4gOVAqI5IQFnjBw7zmjv/UnjU
SylslJHPkyAV3LeqyQH/scqmvEX315jt5WIzSznAqkcWbkXKBJl0URsVi07H4Ekv
IXbJSyE4QZIR7+HSG9epNL9g4sMrhGuUf7Buo7s4p/Qp+6xIV3L6oA2yrfaKKUsN
wtz8YUdHPPIeUI9yrC2qM96c8WyCw4VjhjpaeLox94GJCeyURo4tlTBQNdWGT+ji
DfDm9sr6HVgX5Vn1akq+QQDtjRdtAwNQliHW6TKRxFluG60mwOB6Sfg5+/kRsi8r
EZguQDgOo2jk2OO2csDvgWDRCs9Xmf9DbBIyyCI2eLsRu0VXQY5x8iSBd7onD39O
K0eOY3UpWvARKmKDMwpg8HS8SnrggCMcDXdseZxJcaI0SR4O0TkfOCKzfSs3i87k
AT3pdz9+26otJQZAipT/QAhaGFzdkV2mPTA0opE5XLxtA75+ajr8Fb4HywLfBIVv
mfGXszORMF3Ev3fZwUFyDAT0GH4FENtpxmIpqUTnkK8gEa9h47m+dWxPVZVi+3R+
LcWmsNERBL9xoWrvjDI0h1OQHYXDgBkbZNcfM0akyARHcfCDTMh5A11a4YNXLgjl
hlNAjrb61vQT2UHxqXO6obJKKayXJGZroLUcLVObfEpuHbrn6qwcXyEwvYsTf+vX
XCld6VNwEIXMd3XNRHZ56QWbumJj9f2SOhMEkVgVoJtrHpzrwoFS1Tv0semoxlxC
uBPeCocR6rPZ4DIUlbiJ8Bo21HGv3HC2bqTIchY+Zo5NbswI3rOW3+rGDXLnocoT
RNQapRqoKwgmMvfCLkaqCkWz/Ld+o7/xHgibqgWKJwy09KQ058rqJCRn8RSe4Kry
WxR0wel7x9Jgc4CUiyImwQKZw6He77xzbUa1P4BqeDq6koAoo8COBFoQC9ov2z0u
TU9MN0aawXDMU/VBhYUy9+YH0hYPH3Dz2c/2HGfgTtxzztuS40gs7YZxcVRCe4yi
5r+ZUGdlpuhXtWNXQAAJLLfX6/1jweUvH6iAgAfPBbLKekwZJhMvQVUBE7vH/zD6
HYog1RgL7kawHm4SosE30dDfxc2Y4mfCv57uQjRzlMFmGt7rTx7uUPmly2gP2Ohn
IF/n7R4xVnkLMtJbAtLr/J/2F6kyo15DO4bLBHcKPB+Qny6lh+UnoDQFn5Oir88p
2SWGgX685df+8oNBxrHuJi0bVmXiD0j6omkKzR1kpv9ergdyMG4DD8RTJnfpuUUY
4Raau9epf44XlTtAtYVicubCLiU3wvWF52flEzt03YPHW07n3CSLTKmAtgMVUk4j
PXN4jC4VACnfL0U9F/mAlG2n2ho1mNqrFLFGEUUlUKWKEE14IGfZFtoPWOnyroXT
zDdZKgxDo7MB5MreJQMJRu54KVkZeFi8AcndZdLvpTRQT/WbQGH6bzi/0K+MAJa2
yPNrwtWVf4rUihOa8kMBEu0QLGpGRpgBQ0hKDQLAHGGvbOea2HwgQPzxyzA0aWEc
6tsxc79Yw1pfLYyGbWXOAaTJYdlKywHAL9x1rgMHI8qqpAlMyDIiXuuA0NeB7FuM
2djhhs0uysjCjAn8hoBa/F1tAMrI2CN7PpHkMG05lBV8KaQ2YVin+Evm70ojHo9I
Dss7j29UrP3Nh5rb7wdUI3rYsfHI7H3KFk+4lOcdqeQ4ZQZpAOfqU4tGwb44+Kf+
2AoALAxN0/CCvnRx7aJaLNya92MzablVPLzxd4H9Z9a/KvysX12sxXlDGSxM3BBU
ayV6dKPJ1P3w9+ZTtu23kgr+gBtMCvsqXBTT66wUiQ/uX/KmqHwgrj+vNJ47PofT
uyKc3M1WEnDs3AQ9uM3Ago9f7x8zaiDfGFBW5m5m2tXQbZNwXgk963g3HeFrG+kN
8vtXRBg91jYBnOYTAkx3YJ5GSBcd4jTyRJYiNnpSrCKzaciRMVoIkyh2UMoNSo3u
gBonVvxIiE2LXWl1WLArLWwfkXcpmJ1aaJlwmIWkt0ehypwVc3ZlYZXJ1ItaoVjo
t934lyC5/p+bZ+YBALCFyBnb+7Xq0x3WmwSKxmWgjXv/Ham7W4fTpoI6CGQeZEu9
oewGUUVNfPRxi99OVRke5/0t32RQOa5sQqQsZjQrXQUwCo4M9rxcRSBuyKjkS3CA
bPIwJj4aQ/Y8mlGDbnupVB0zjzpSK9vsb29903E26Tt18apPtTzj2dyarr5ZC4Yz
FuInL6osB48gFZSDpFFoVwXmb6x+TQtqVT2n8pVFy+mZ5WDQs1ZnPaCkt6rCKkkM
2MwS48kU/9S3/5ap7a56ub03ekzwmc0tX8h7blHTWCfCxkpjjNYcE0qFSMoydZkW
/RSicOc8xK7ZlGmDohUY6a9sb1XdG2mbPjb/vS1S/BlR/+rfoSZjgZSePT7J4cjj
ZrK+MyYQfBCjcmWRRerWJ934zMzAuhwboEhIlSgbo3EphkgNJLogx86/rqnn1dYr
giDzVgKRyc67w/4QvDOA11Pxv5FMSXYLURbeUNiki9xBUv3ImuOJu6AyEWj4jjQQ
2BqiO5zXfAOvnbPgqwOxCIUOUzCzdx1NJwu1IYmMGyjQDp1dSb+PG8r/Ztyip+az
IJv40AlLU/SHpeciDG8kdlvoFp4Fry6XN8UUEfTEscgVdIvr6QSlxAXioFnXk6df
ytTRaqurYPkCbACEmQYyNdzitgqgsPpn1ODReaVoKhyGQEI3SJqTtZrkjQ6OvBYg
Dut0JvMdiowWZcRw3vH5qQInI1z2KTUKkvI4sflN7SdsF9SqKmKf53yAyyKwAaHt
lxaelllpcG5aeQ6k2prXsOZw+Pxt/lYQHEcoyGzQb0VoDPCt5BJH22HkqHO2R3U3
HEcFi/IsxynLWGo8MF5Xfhs6bJ3ucBKLWZrn7NwWY/JhFIpQs1jH/3mLccIoKZx1
3iQK1VDxpxkbWSkZRY/U9xVb0Fb8cHGuoUpm68EkuZ2j3sDhmDuhiA4SHhTLLM4z
0MKc57ruSbD751+MTWvWnLrbhcuAYN6deE4qUZH6a+kLYbzgcfxJozsHP2sudajs
nCYsAs14AcstqTReLSuxXnv6gTe1pnrXflqtX0so60887+IAzKahURC1+Fu7oicu
CvrpfyX+kchh4E61ogo2B2hkWV26Ef21tnpHy6IOR1bDm4Zi5GV95OaNbYeOKZfh
QN+dqQuJt8tWlLf8vMNApN6cMqe0WTjgUesMRvq4Pq/bXiisnpzGFWa7UrAhFXX1
5tWLMr+S2QfJXAJayhX3kej4AE0iQMzVWQBTCZqVew0q1rKwVCrk2cme6gjkrM72
xrIatNOkI2X3LEX5ypXq/uZu+jnD4+MiKv35/khqv2ml/gQyt9U+oVClpSY1GsW0
gtK5tBdjCgVQf5ltNdicEPiFAGCkyfmOolQKdh5EF7Zv4XonOmjJyaSnCrxB7Bct
5K/aJJmtEBIKwt9Dp4kJtB6Zi6T71F4dWAW1tWCj8e+pGRCvWSAOb3wLdxBx4P33
Bna4lc4H4nYoQ4Po2nS4lmlFHpHfAY3QsHSv7vv9pvvjVIU8GCRcAgZcso6fHQ+w
dL+K1wa8ZW8I4ir5aTk5Rfq+YOLA3ibC1+Au5aaAoBtAIEQhnNa4YN87qtiDvhKn
cae2Xh45i8sdtAC+XrSfO6yVDI7VHPlgysjtjLkSihyUFe9Ek4Pg+T4Rta6CUztr
w41oAstcU72VvTqFX9SBHcY9ORY7Dm1wIGNSKfkbSaVMr7eHilirZ+qvto2ujwmW
Cd3qeyq36JM3PnqNbyOa1IbavCP5g8ITvIW+idHdl+XoV9QG79mID07GWgKpPVWN
tKfrHL4G0cnSOQ0dDID2Ujeszz0181ovMTdUbPjPjvxncnytQ39AFB+Mu1TEaG87
UsLJ+s3izgpnY9AyLjUUxXLOmzFXGgg8RJJCB6T6cgHZ/rFBOJU1JrcFngZc39u9
3blqdYLrVaQuD3TsC2WGx2M52FOxnMbOk3iiZ/5QPyTnazCEtgwjOpi7IYJV5v2K
qMpAe1G3KE2kES9UWX77VJqys+PJwaDwNJpMWWNpVSaeiMXqUqWeOFB2e5pcNoUX
B2xkHvqB4K+RF9RZIvhxizrEWSCGcj/Yfj8ZOYd4llshX/dL6DTGfGpY0MPDLZkH
ZkYX8OH4gVoIDGzb6ZyVrbpWzTKBzpDvMoE6eYpXUtaOz291KpgGz8SbzD4wTItt
Yie/+IcgTkYilzJ0JCNhixDB/6jMm1CrMyePRqiaylyx0ThyBewRtnnh4TPNIqsV
8YkxKn/p1vt/1CUGaf+wwi7bYBpc4q6OBzX8DLXeRupt2GjItVjyTP3/daI+d52P
fZ0NXFfun/B1u+dCMMTOCK3mOkLvf1nxLCh8QAbDcOhLogZtJFRJNSmVEj9NvtXD
6au7KJoxvnVyTNLiPEmXuT+KjXqwWImgij3YRKUvh+xD8pCH57CEWQKAh9MLst7k
eo/p2KaLYEeaKhizv/6qC9At1G4IcCVn8sCJDa/saQidxYIpX2bidk4GP5U2wqOg
74gXy6L/T/as0qSBmBjG6hLBvF5SVBMySABHDYvDpSHOy27BeTPZ9usDws3nma3s
H6zVUADDcH7isfikfjYuv3BTgnhb9pg1AcqPvbQKVvglEy8Nohmj8B/ZpIpG4Y4V
4IFLrlXnGbnah5v0kIA0gEw39qpNmtJf85U1SiZuIkwjtnVYqji4abUzN2w0Ae4E
7xAQgOet4RvercEDMbM6j5dRVAlEtAKye1Vt+8gZpUjYavYmx1YnyFjtbnJ7fSpC
xhbDCjalt5QDH7OotVipubfvnrnuQh4VzoSoOBdRadhtoyqH+PlYPlcnxCT4tqBP
dc8ouPDSMOKohfbDaJgSxLSS5OExy8trkQh0OYKbCwi2kGFeOZ9z4B20OLFynPNG
ibfpJCpAjTEiTdoND99uf/HsFWP4clZKmY1y3T7VLAPuZRsf6tSo4QBZDXvOx0Ly
UIq4ZcAtWOgxLwmcJkQLqsUe1JoEYY4o+w+kA2MUg60HOZvIgWS/pVFKoc3b/bED
LtzvTRmryMcHjYitzkrMCbn3Sijgz8c6g9HNpymFyK2Wnc+olhHW0Cfd1t6RiIly
Hm6D3D4WUrOl2zw/KjNUjuQwG23UBbLgj6Yc1rkydGWqcaxC+SdsOE/8ORyZtau6
mXtj8JgVwWy8RhBMO48cDJz3/VNatxwAMcw5/4KXkn91c27eWF3KgzHhVBU/nuVh
K9PJ1YaZaPgp3osmLAqwxWZSHMy36LbCZSkeSS3M7L5zvAyt0pQg6BrVE08EtGvR
l52WaAqRw28nuphMsqY7GzZHwdYWLAmec/cjt9o3NGuWQfWXInWte8VA0S8OUauZ
/h4E4LblRTVCLBpmg9xh2pNKoy7Jc5F0xJVrU5pBZGgVzQmYBxTagv+7LSXNipJ7
9dBLJ1hBftXRs8ReAmGh3LQMub9FVu2jyUDXzeiBYz/OSsGWFd6lxkL7+6D6CYEz
7LEQYkpyOVLIge2DXZW7jK5rOwHTRxO9Fjh9Ew5iGh59Xg7UbJiU1AS+bkqVC5uw
12B/txJJDmqZLDNg9n/MJZClAPPLvfuIgf88F4kUQuybOiYpsZF/wTlIh21CjByw
Xtqp73rh+CxYpwqcg7U00Tur4AhODj4duDBWsqF21/FcxzcEsEH6p/CNJFOAHxMl
kqKrGpYo92q/ojtUWYQR6Y+tkUpI8SUI0nHGCwiSu437Uu4g69TtS3JOnak9DoFk
fBUGYMaXkMehvDuFYusGxHP1PKn2VxW4XBfAXZG/TMR0A2/caRibylZ0IYZBN/RT
UCAvaLqnIW+QsC60btruPhAHiEBvGuUIgc/cCu0wjdOJwPPrjLhg3QoCEbc8GrEb
KizYE2zAH0MC/DKojipDhPpEJ42IRWxatA0NkjFRMnn8cYUEviE91JwJqiGCPkrY
3gj4W/elSoEFmfWX4+q3uGohCreTFaffYyDcvlAuX/EQ5HY04UlrRT3XseoL3FOQ
exNVaMQzf2oiLPWriwh8Zt+jh0U7GqINHBz3uFi0G1VIMJS8HHAhTaPvOZm70O+K
3bDBuCIdclOR0Gqa80TgOylqzzZFPHIIfXCZu3SgIBxxOX5dlhzntr2xGxUd1b5k
2ifWDzzCuWIAo1iMn0QekzsjBlZvBPW4du+dDFu9oGQZJxIztoIL3eE1sYaGNvaY
oIw/cRlrb/houFNRFmuRZUW5wvtfux2hhVHsq9Ls9qTx/aptlFMppL6fXiFvw/kU
fn8OeUorevRKNYxmyIipWOmstO3OLCx0L0oGTYsvDaCf1bwSAp8S88Dvehle3rdL
ddScNqUBO+3YWWKJt/sBtn18jO0fMx51j4a3ykWyj5LrQrXvbVOAH2z9fPriLdYp
CKZzd7btpewlkUN31lm7J2m09vccj60hbDGJHAAHSym3/Kts9PCh+0o7tw5dJEth
rHjQuGqo9QEl6R8rpPGrm02aZ3rwK11dBYw1ny4EbzQYmJZ342hdleW6ZGdRgvVJ
wWqyMznqBYTxPkkq9lNCPH9Cre7ub57ZDOF8l6Pcj1YXA/FKdODDhx5yC/G7riTx
fbsAvHCHfnk5LUwD11A5ybZs+hSeG+OtD94lgqbQRIc268CvMeBmfV/g+tfnRSqN
H0uCfzLJzvj1iHHNac4ljHk54Z0dIaudTVJTAV1HaslFkBCrwli0hsUqYv6Ez8Vu
3py0ZtlMPR1CjggsloA87PLFImfuqM4GGIxjQtX/3XqO8P8QpCA6bhC6Z8G5FlMd
2W7p6cZv84o/uRsHJ+gutj6+f+E7upoBJTQsvhCnVKJkvlGRO6g4rUfVu0NnATZ9
6qYko7MSmn7e+Hr0dhyFZaBUUcJPmdY3PHepcLUM28j2c1Ct64u8hCvE04ElVUtt
YbX+w2qKJqmnVpDPfnEmPvXCpL3klHfZWvtFvSSv4y5nqrTUATz8+71UQ3aPQL4p
y+F8ZuISRN4f5aRuJXXYgEs1306OIMbWnqRtQDNJCGSLcozrB8y/CckxggCBCKsc
jQNXW8yuCJ+ZuOFd6dUo+ZT3O5PBCI0GzNlGA8blkzLCn8gLQx+oyf9W3mC6thcd
8Aa3C1xm1vt0voSzEL/bsf13sIM+A1fXNM3HUC71JyXbWp40MHTRIUPnte5phrH8
sbI6bbkjujxWT1x4iBH3DfXBW3rAmYHwh5kfxu9/UOoKOMddxoIpopOzHJN0M1OI
fmfl3q0swTDaQFVEHaBTEFd8jkY4EYt+AqdMBOWhYRe8ShqUmBwcjxUiLlZ93fw7
4zUBvDpd2Q+xCIfYEt0jjXeVyY/tUIbdLQmk8JvPssRYaAOAtd4U4CabMSalT6IL
tRyYUx5AcbPzhre3nb2WCLxjwfeCI0RncqS5DuMY1TnP/favxN4xVin8nRJM2Lt0
+aV41RdmSrhOE97MCKexyYMkyQ359amFbBqjAaoOoR4u5JJi/bykUPDvB/I3FtGz
gXljXYr+SMP78oYiihW3c6XixVb9tGEPnMYzE8azfij2yiC90lrygYNVBWPYyvbl
Q2nDbzUj2NpAbqVgm5839np9Zte4gwWnaEEAZEZmRnyeKrQK20DYdjUtd/zY7VY+
ljCPiijtiw9nRCHuXQve+xBtUr7+cGMBzVzBJoAWvw8ySytnZ1Iixvcz6xGVtRzC
NGFeNNcJaN1/j4CIH9LljDX7ug9HELhEPz+kleYelI5NNztxcGGnvwXO6v11fH51
XYq11VyDIHnfdPfKiwBz/ADC90DS9O3E6OqLcRgUcJSAo7sRB+T2flby85WmRXPf
UWMDDDGqO2naVks7CLipcKKf6ot0YBucI4W620H+cWwEQlGLhCjHMuRo7ju+tIz3
5GruqT8R8Yh3CrNCHay5J0GxIkD6iazzBIWjBABShPZPbSz6HHBVG9dijU9eOz1o
WWmMMAztQqFKWEnscFr+wv0QbEUlNDq4gIo0AbDeZTMSLV2QMs+IY9d9zRAz87BF
y7+al39uf/Web1W+sm7VzYh+O/v4Q0fAU1HbHwBYTg9v9oc33tgatmaUnxw8VTpD
dLZvTQpobuwXLp7otSejdtL/Mno6sF52P1ZMlB+eSw1sWs/s1IO7YnQCpBF8GJPG
x27Vg94PeKUOgvqNVP2fO67oZw1d9yG+AtRa4rdpj5LqrXfBS4wyMcPZWF+ZGhQd
FbnlxVpSbi11+XWac4vJZIyXSRnjVqzy2BVyJK7QQ71TG3L1sfPeqKgsLm4q0ijy
pnlJzGQztCHAE0GGGjH1Pl9JhhroF5Yv8Uxs79Pi88s0qKpDFBGGgbMdy2hfb/eJ
nIBhWmRQojJQ3m8QV/sg8OSRT7X3QMRPWSTlHv9NsbIJ6N7UbYtyazbW6V+SnjST
PKgvHsq8HEMlvyWczPaH9NiLKXPaJ+a/GXXEvs/OZGD0u6We7XYF/g1SMUU+rXLC
7k4/lyaWEjS9C+txM8zXnbjwpthfwYixhUeirXgIwWXEQTuPe7BLgAcxGQO/E++n
EZtf8d+Vvak6K0s81A9rro6KiLax3vRdWezO7FgA0pYQrqD8O6h48ebGnI/Ekj9z
2xrM644YqUzxsYpXRWpmE67dsmyqiK6ttfSaoFY4EI4bVt6suuI4f4gqKeBz7Si3
GNNdyiD9hwKdqyvuBeG7b59kqUnr12RfDsd8EL6zqEvce64g3NA25/7g6CQ95QXD
IjzG1nll9oIJy5KBQApnn8jOIfy1fbtbWrrgkCbvh5uHn4hgk7gbhVSsSKiHHOqF
AwjbVIZ1pvDg+HcMkXWI1SQYoIKfWCwG7L4roV9aogJT+u44GySqZOtcuEjjACSB
zaHHdVEKdx9Ye+PHMDU5g7PhzqNwiZk6xSrPdDX8/y6Cuo2+TxQSjjWZRpkGfWLq
DtQpcw6BC/I91fkR50ub6yYq6tqZGgUZgg4/ltdAQtTatLfk5zX+IQexFHhEUPZk
Hc2lkMN0fru4/xsYDPIpzCoL7DBT+q3sh7PTLDJd+fI910n+j/ZTdBNib2IDHiVY
IQzwOfTopfUgSKUh+Mx+MUaNMOiR7xRr3K9xvK7Czq4i6A9PjFW6+uid/SrQVZhV
QxKpSoFbYTYO2VJy09Upedo8Gujrs60iYjrxzH6qJc9e4eVopahcc1BjJFKlX093
O1THGkqFX+TlniWbaIF0WvLq5nAO3PY/xbv1WXIzAuHa8bFD/GYTpW/N/XKUOFQa
3DkMCHP3Jd/xtYV95apgVlKVy9O7RF6qAKjFHYIWLEp5KbONJDB0BwjjF1mYBghW
TG8sA2NzhnaTH0WehxX4CzzAflPSm2+u1YfGeUm2CxI8NUFtdm/JnSIUcyI/37fh
/L7LDcJjhik1LVZMoerg1ilV2FH8zL3yCeNPGyiN59S2Au2ftmp/xFJxk/vgdTvk
RZodk1pMKKImd+r1jOBmeqsATj+kUt4HgvnF0EilwqF5RcACqH2ptAL6WjPvzHBH
/z/1FXSb3cocv6hBJp2D8jnX5DCZRHC6tWSFfAz88Y/OgexG3b7f0w21Hrx2Qm76
djX/xobTbKu8PabAHJYzCAyp60dfgRrA7QbxYts16SUe4I4Lg7wspulV5WVVDSvU
qMAoyZuj1/UCU3+tXCtw+FPbEMFSwtoGNhs9bs0nloqkM9IyZZyheCjRHN2RKj7x
y+EDWozTXqfl+7p1ZIogSf2Sn/wpnxLWFp/T99tc+sKeADwzQPBFYYA0jVBJfYKF
2i4jsFjnfYG6k3Th80fZHA6zxQqcTa3c//7GyrXmmldEcBHtH29eWNJzWz/80ZyA
2UhmDAH4HIUdeqBV+eVPXAE6Z2rVJbWrK2vnf3Qx/cqbmtQMVFeyjuSsXipgju6B
+uPXYQJmvQtSjFlgg/X7yZ7zE2MN8qgg+hmghYgNx60cKJBbsmF04G6r1Yx1Xl7m
BIOhHd0SquGTAsoWZx8xUnw8CVm59++ID3T+Qd2naBJ9/+vI4RkMRb4NXLngKKUO
nO2ZASvwSoTit1vp2qyN1Dk48RWt3A3H/1qgHP3j3Co7QZEPtB06nTkHesiK9d/f
s2yeBfIo6S+8XC6V08zlsVd2qJZpDokVkLMopQ9kxtknU1CahSE0j+2MhCvtrGgL
eWj+oXbJwqOway8Uhh6dvpZPUvEinAf/VO2L4CJcqAawbU6jMTfKJWqQLZEvj/4t
AM+97HjtgTPTD/3JaUwJEC9uaHC9MOGYVyOboJFGTcZlcIkCNIAr20QsaA1+xfWl
ZpeR5He3QjvGpa4oW79aFYnalsW1lIk/bZ3VB8wJdACQ2vr3tA6UbTyhe5jLhsf4
GRFmHdgxaKUF2k6aEcevL+74O1QteVkJfUcMojybO5eqTKW/g0OUb1bKwEe294ac
0Wu8VdFd7xe2GJ2mbFapYgP1mrtA4DcFIob9bnFGLOP1PhP/skHpedCNKSrNKR/R
9vheaaMhEm8GthpLpRtQnvSWX41zyFkj6rEeAUSnDocmNtlAmT+U4/c2HPaBnC2z
RtgKtowdZnKoaWZQxBGH1UPIIV8T51bF1/ukQSNQgEk51T2cgzqPRaNSyE1Pe42K
RMfCqkpx5nHtHTmHO2xVZYlcBngqIpW6vvjx4j/leJRXvPPUt4UVTQWKrQiJelo5
zPLAEcknkQPjen09HnON4O1IPN7iMlIkeSWGI1s9EWV0ZNY03Pdvexqfyc87nEJR
YhPvu9eOAZItYyFA01usc7XyMYjNE4YJRZEd5Ey9GMbTo+AZD97X9kYKBdu0NbdD
+uTyWPc13/wVW2fQUIayBPBo0OFv8EK4G7VPWbEBexsrk9WJ9FtTS9ZJTT0s3/oC
5BKMtY7OV00PFBq0KdhD/xO37SsRCsBB8KAZqTXxtPJt4KasnWaTOv3A+kwSAHO9
fakWzhyEqgWEqnZQYFLrJLq1GFsPxW8sPTptCNwhNs22vACQGgzMBLZhqsh6jp8x
dM0PS47pD7XM3BRVyJC1Tv1e7klrStk8yoqsx8Wtq57hIRLspVQ45LomJAIpRQiS
KJAu70CkywOFLpAdD+XhtyZedCHV4uuqWQhvolDMA2Hiz6wfBIglIenk56LE9u03
3b6JJ9h3vqRK1fBcCwUdGFN/hGGKIikW/xXLrxlMDwWbwbUnNpS4ASoLvD6fkh2r
3gMh4qWTOmiJ1ErenJzwVx35uyD2uUBlSEJTJ5UAYYHo9cmgZNG20JejjkQAr8Sq
UP9tZLKqGI80sIFYHNb73joANw0l9+9pVpB1NKRPo1ziR/lRqqVGCmq1NHkZDiSI
UFbzJhRECvWHIhHbrmEw1uEv28uoarrh0ylh5aBg2yTRdOkxOg1GaHBr0WZF7Vby
uit2+GtiJzWAB+7Ft/dYZvEZz0tLe3iMEQlLkCj/zJpaMInY25mDaY33Hru7VViP
faQrLeEHJwo4X9n/wpn+VajUgk+QWnB86r/WFM1rHdY2teNs2b3P8n3pR7Oi/9er
8Qv+EWud7QXKCb21gDgn0L+xEvrprSOU7vpK8dVx/g0IfIuAFbzysGNWftoAs7Ue
NA+OQePIvIR1Ye1gWtLrTUEdQsITxabVct/ItUa2otpTQ0aUhSgoRlmM+2z1Ahq/
KfLO18K7+0wVFQvjG6Z96K0unGOzth3SFAyHX1LZ0yXMb89nnpORVuRW0UnZu2+5
QNYsRlZy6xsRHh1e05Q849kdbNJ5k4bc+plGU1TcDXfh1p3uNXPTZaU9X1vqHyBT
h4QUqauli5bh60porUpVsV/xJn/rcznNUhTsuKdpnhj8T5InqxiOHvLKVEHnyfj8
+nWgIt7EVYKAh81M4KzfeYhSPu7yjU7wTUa1r5dg6DJ3B7AUACnXSWMqcP45smUv
wO95XMGvI3+hir1xWMfQINxR0BgcOFFcgmgBUk+Z4/VKTqFdokRqrs5XL7kpuVaY
ffuWcGzraCEdV+UCFfM6YqIFin+xesDWurNV7zkVZgzSGt4V28odHMgsLGhv0Zcr
xhmxAuXuqSuJbeyIhDKg4Ui72hNAZ77kHUrWwGBYnOfs851lTclZiwb2pZTxgv6C
jDfSH4ejXrCFM7rEQEnFeR24EEc84HU/e09LMZvwXSr6e9yzlY3gndFK9bMWC0l0
x+ekIhUE2u0yuWXnE6M5x7vwq3cW+4vX+e4HbWgAgfp7vKn0eI13RI/Xd2vb4Dvq
J7obMsFFBiMCoJuZ0ID0slKSPRfSmR+ugPJjEUgNmYqteHLY1sdch0ey4Ahsv2+F
0OrGXM9za/0J3CKum+YGwFlzH0PCXNaCHUziCuGS+Tgcq6SlRkCO1jxVn9XV8YNj
vH9a6ZRbb2WHQE/r7LItDqHLNvdOTYAdRMDQDdJZRbPvlGtBlhtFxjrgfmcqlbV/
pDfJdvJk2sWRdOUzHxTdUckPLQz/Oc/hQ7X76NqlVQrNESKT+DBNtxzNI/lMxztO
AcGUNXD62OvcA2E8QtjRpforg0X3TusFDH2sCBDX4FKcwDTeMUDDaDm4fkE0rY2c
0FsIOolP4zmxo0W2vB2v8WemdxKHad0MdGYYLyJaMXuyImRFopESn9BvmWgrrXWm
LyYHUVAOBVDUgMNDz55UDmyFms3EaNNoly1yQRqfQsS2fu0Kn5D4PP2fmaeBoymV
hbW+GeIjU4xdKQkMI7so3KAD2mhVJ0Vv0+LZI2NVmqWoo5UbHbB7ytadUJOtyPLl
H44h8JDiMQ6aO7u/R6zS/Dpx9JQ6YOCaMD5SMmnHkFTpKq52IirQ2Vtk/yA1JtHZ
TeaMIdYKo2rRGhfTPbmTgUHEqgwo307HubZTXrc1zh/7LYECXivIlOXRxT/zJ9Kq
C+NaxrgTNgqwSUm7Ta6gbFZg9V71370qKLrUxJdNIydEoFNKxOSU5Y2ctSoJvGrS
SbFeJ7jYUO1uK4kUdpccoOEtfdFRlHKN557PvjphOCyJzu6SacRUAUPuv2A95361
/X6LXy0UEDv0xH6SQKUZHwZ+c0FMMNH3SekQPO0FQgMUDO1UffnVItGqlNSmMDH0
PPhkbqVjtZgUmPFerDTxm1WvoUC2lDh5ymFbXt3m/ZHeNtNnprZLIqMByRdI7eT9
ZAEX9HGQhDxmt03OOw/k2w0SCYlf6crJZ6rbkjg6xO/qL/9m0HAGzLKe/4fD7pYd
X715C1UD2KA8PE7e0R8laQJTzRj+Uf6B7F/aRk8BpXmMSjUnIiSEbH9HBioGgUWM
QP3OeQN9aebNHj4akfq0u06+uvSWggyClRn3w+hNJqU2lYx/tfnaGFZHB4E8sAHD
o/CiASMRfmOS8ILIBtLjHdvhQZ7HaLAKgkdLugF3V6RlUDF5DKMyJDB+74XeNwNW
jpXoGn9dLizzE+92AmSIB8pAZyAWke7LyuYopIOKsyykUAwJwPUpP2wWUSUFx49w
VDyVLfbIJ30nXcwpVtz7RBANmGrBlBHdlvWfOECzlqyTJLAR/1t3XS90S+m+T1zW
+0aertxEowwVtfNbjRZ2PM47UY2fD2+iprMT93nChjyUG8PQNMr8OAc7ktR+dq2O
mEyzTs9nxP36yF4XGOr02K4dbRNXmj4DMOgwEDX9MDeVUcftfwzuKEKf3AHgDScX
aYeL/bzL/kVxKHO2LDIyLvdZXGcS4ZQRSZg6rJFNzQ33z2sB8ArYAiZHq94bpgfm
pl8f6FFwpvlR5qfIwxmFFBpf1YwykViC62zh04UtYg8fo+GkIue5ETFRXl/tbXVl
+3Nt7/LxVQIeDvtlxqJP/3AAF98xj6Xpeec316f2G2uIk+Tfxv/C+iSyT6fpcIRa
oLBJlV6cZ4i+2UtzYksSyNtr8PRuVbtucdLJ/E3Z0yv5M+a8iJmgd4o5NDLGsTQy
MfC81Pj6rQXF+bFZTFzaSBh/MZdq9yrnoBtrHdkhRR5nzuKeAeBzDpA0MMUwKtRw
EbBbfj4muBtVxti82NYx+DCUvd104Rz/XQBDPGLSrXFRtvakQ8fWxWQJ7lu/Zo/J
Xd53X+rPsjGOWs17K4ll8KIdVfRUq2lYfmhme6+AhREFwLoYqM3cmFvxxGBUzwwO
KmWPrwjKQSmXdjhl7eLq7z9FZ9D6rizDYC6XgMyR+n7P1kUBC83S898yQEmJscFd
i/CAp/00I5kxVrWpnWClOVrsiCGcto4PIMl+L8AjHYyv1Hkr5i30DBzROUFUXKv7
qA7tqYhl3d7hXM5Jo2XaehSh2k75o4Bxd8OFw6EDwqKXoYmEH1OzBw5sg+fL6p37
v06P0ufTrRbqDVaCV9uIJ0yy2VpjulzfO3EobwSthC3fS8zX2ogNwCXGsXXHlUfn
aNpkCMx3KinOrvDs4eWDkbDgmKciyHdlI3DqZvGd7KWqRgHsO/75WhUTXsEShBL2
qUE3Z8AWHvs3AZatYOBuv5n4kC/gKzWKOPJvwJq0niCrzFO/vzXPmKcshEZWcAo8
fwOtJ69LlVwwTiUK54LEzvAeod86phUURxURbYP6Q5D4OF7j7l6lGcfBejtbk1nW
+8vs7xYtlJZ1A/Wy18Z5sHD9oC20PZJgAEEz7OfrrxTycRw0gypbKcao2QWSNepG
HOxxS5ZqOatcgaJ5a5cDYSycT4uJ0O6rG/rQ2vnBoIm310TkiWbdrYMSdxRHPUEq
cCQOA8aU8mEX5BGN3UfPc2HZtLA05HVDSigBSgWvbsXdfFjWNfYJbq/5n2qWvreq
G9vk7xy8KTZuY+gzLTTB0VqIVraNwzK1J5jhywstpHjBWrDopc7tJQcoZMUpPzyH
ryno7XwfXW7RrVgGXGX37UYal9ya463RcajogsDhddZ0Svo2hsJ7mrXYztBUuELV
84pm94dSCptBF//b47vqs5Fjm6BzQOEttmr0o4dyqiRyEvrWpOU09I4PZte8bERJ
944i4NVuA9cM/62q/LnkAwy32EAnuPMhdRYfxeAKGbGc4daKPwlOPO43iH1+PMGv
G9GCdl1aY1BoaEttSvPFwnXMcNBxluC8dCaYkt9QAQzQYgJKpTaI5cvcFBtH2C6b
FA3n366jVP8N/4b+WVCx7A7bwQfVgyNbWrhf3n13nykiOX6V7VAsTpYDvYtCa7FE
qQe6l1/DWcAVR01EPIo1dDvPj+Abd3nei9HBT+axnof8XC8G56h1PQoE/zREgQ8P
ouvYVigrHp1vwtXhh8Ba33mzUkzQfVcdQb3Tm0o4whzk84BCWw4lFIqFL172cwjb
3QMsEs5efGrNnEYMWoYVqvkvcxF1HkgaO8jqKOlrdVgs/GZLmkblWcmVv9754h0B
vZIvt44+aswm9bKc2m6KOM5Z/sAtJbvkxOj18plBLXqRZa1p/GW95IZ0btXtZkJi
UiSj8fmDmw/sBvzj7DvjaKg+Tn7EaMXfOtOmZiTYroZs0gFBQanaG3KZ5OuouoED
mK75orebCeHFK1ceNEGtqT0Aj52bCjQHAWyYu74MH/w4BRxpaHtZEK6FoWxJNvnK
41Rwu5lJZYFj+twRO8enLDvaaSqnNuPkOAw4lHrtB25WJgWCf+RUE0+0fH29ct2N
rlQwnUjrAMVN18dmtM6rkTnCxTByduySsotAMeXLL+7EziHoEM67iDJGVFW0hHxf
xU5UYQzzrdzVdaHzVgSrRSWHrSnQ0FNrsxVC1SJhJpXPknvbzv15sAg0Aak3alpB
8ANE8w9PIv81rJNqYYI34BjcbRVstCDnc/m5yJmKGB5sSPNsTmoOkp9bPsPBJ2Ns
ZGbdnGcqdC+zpXDatIL9N1wbr3UbfNVSb+D3WXuKpCj/T9dEBQ9U0WKBOvdDrceK
9fnt779DrcAqzZddZZF4T9eV3ZN/s7z1Wwm8YGUG1RnwNPZYy/WoNhTCU0CVQhaI
CGQt15A0AxYuivzM3glIlfaPEQZLsmfQjuW3y1FnbDxTigI2Je3GSOH4Rdcw+85l
f6563HBBzha4Q5Xwj7O/p2DsfsXpjLO5Bn0c0s8R7Vw2c49h43ogFhU6OTOLFa4b
QSQ3LIR28n7bHgfr98S0dAaBHLieEF1l1r51pXEQVASoaxJHXGTtez+0/aEEdTjK
KARs5f4+gyfZc7rqVTPYMeXhizuMdwj3byXudBG3WUdSSQm840S7NrVKPYuZok62
tyC0xFE7iPiS6HG/TtFBhQeNqhKzPLo1gMmjQlWLfJC6FMYfRuH77lEUFMBo+y3N
log9K15aMWAZtnrxYh6WBPMZJdW+5CmkNPJq7lhWyoYBiVUPY4kmvGz4mQmf8xUC
JZ51D18PNKEcSPD8ubzzFk9ni8hDgXhXRvSFQJUNCXabcSIBAr6Rom2niO/xg/Tv
cJHzTKWmbj7y/cryyj3s/P0SnphuwVe/iNI2YgGMUbSXFK+hpXG9kyXOTj9acVRu
quApJwPu8aFf8fyGVfqgvZUyctvnoC5hh9O2VfTUE6lcQ7bsPhc/JUx7WGSTtYX2
oAy7WDaJh+m+ufbrCVYsNDfLPxd1NU4JoC/aGRZoR/oMr1dQdjH4xIgyHm2Pj/de
lp+Yr7jCXM9VXhOeRDWtZ8nOPvcIytT5nXUPQJg0TT+UyoVYmIaFG/UUy8RezTuy
AnuBqQI4+S1XP76lLpwZX/u57Lw4yv30MOqgxJTagVPbE7gfG6+R6wxF4G1Rkagx
O28/u8U7DjNJS0PLZRKGmboj2fjnKRs6704IgY51p+/OX36a+lNQVQF9bu1ar5do
6G8BI+WhuQXnLG39O8LejPN1myrJUigL6sHcASBhBj9ykRGDUEIOBJf80Swk5+kx
ICZ8Qq2InThCMS+g4VJTEqg6ePNvwEPfrU1cfSbJA2WXrbcMojgWmfXjXCJ0Fkob
pr+Lnjq2VB1xjK7NmZyNTDymjhdtdxZS/WQycxe9r95O39ajrLl6MGKr5bE13XaE
gItfzT7F92p1TbXaao4p9V7+kTZwCwHIJuJQtmeO3m9XOHH5lcY35Qy+0bbrIzpD
TdtgdCdZSEE+qedaGOrJjtRsUlATuyv6JbjNbnQ/TGwGks4qWABHBCXmh5hbnN1d
nQsqiQ6e8Z1fKO5YzyfoUWBHscphA5pVxL8Ba2pqALIc7takdMLkZEFEKulld37G
jYYyYEd2VVFnCORQTZ6f4DpSpMc5MkUA4Uw9V3UE86bVODVKrNq5qyZBr/6Dsd5p
YlidpZgeuV5vENjlKv/RcK5QoehBbfHBS6e79d1WgGd2A38dn2sb4JUy305E6xuJ
H+T7Te9lik7SsXe4m1K1AUW6c94n+M5cvdaowYCRhjrJV9yJi04tR0PaX6USaQNl
Thy2CHrMG4XgXkuEkKF/wTMXpA8odXi8YY/eMuNE1hrgDTikPK4bwBvBh41h3SI1
xhYSX/IeD9C/gWIhim57C8gTWc3Cww9K5okD7BwSN4Lv2F90t9rMsKnAxp6qY8VT
ji3ExA6SnVG1jOpR7ePMA/9P1Wi12nn8mrkJ27TLr5zxK9m/5dq3tDYZeqnvlAuj
Ysd78Fr7b20iNfBB43PdezWnHwb5wewi4GcQw8WY7X0mR1BwOTUZ1OCRwBG8Z88/
9+1ce9I529dUusx/oyzg5oMiOoeVHuePP9hffnKFW8ZPhCLcdrPKjco72QUu6u6u
nChsAPKIWstrjy2rSlPaMQnuog0WGTjg9CImVKtBybGs8V+tSDOndzqxIyIVwE8O
vp0WaHClTnnhSD0cBFbYueIrZ/TX08pqCF5byB5rnaYNHTKOLSewCHSgovv1+fE9
3QlicA0dozV58Y+yd6+Ai7kfNJoW+pC4PmLypNSp32MQrk34dOxo+tM8pn4Pb+SO
C2tcW7fRwGyLVUP65vZq5bI5bBq04tmxm36zvQEh3Tc3sbvoM5HWEx4NBe7L35ms
0DrHNSwru3gkI1z2AQBojLeE2ci1gF/UDn8uFOSoW18LWy1ll5S74ULPYJVBRVSR
IYlI142qdWn+5LxwnpxocvUTiT2uz4r7CCrAm4XrJWGJYMCj4eUe51KgJd7TsWKJ
CtZj+wOsVLr7FjWICklpA7SseLDkpransqg7CXc5vuxn9/73Fibgsl1Q4Q0lCMjT
0EEqpxTUTT9VlVcMjG0DAq+GdZ1uzWwf7MBtOjwR8ZkN1avWnF7M4iG9xRGweZpx
Q7r2of3UCm7hqkq5+Pt/kxEvAqMF06nfzd4KMELgDlLyY+hisUJwDa96DMxyd3M4
B7RITL87AbIs7UDIid6w0tsrtAo1kbjqXnOIxt/HRu7jyw2L7itcZs3SV3hvOaGh
CM/RUEPyfqo6Ij2O5ySlVK2+A3CY03voGsi2/c4OXC5PFBZyPDDhEO+8Vvi3Lk5p
g3UH3MqURY1l4kBEt61iwWaPQUOBKiAakbPg1G0pQornZf8nnY7Gk5ehO2liMTD+
uhV/ZYHiG9wzusnuPMrdcXlygBUjCgVwlN5Wc7arww8OOJU9N4Sks6AC36PN1ACO
muNm7rdG8excHb4cAXwqOnNJV1V6FZFavCaVy+UVYiKuDsVMixdxXoMQrpYa8rkR
okMGXNRudp4cvlkd2HHoD5Lfkks/TD8vequ68VV86Zai+W6zyWQYQMpTHpQR9ZHK
3eSLAUwF+5RrVrOeSwLi8V36tDToPko+BckR8HbGDMvBGEZvPnb8iTqVlVS+XJqH
bEvet9VRForacYFwkVmmZJzNXMALmt249Fg+VMuoKiwBWft9wRqeXQrys3C3xn4M
Jt7/7ycGPQu7MDyiyVvyF1emD76iIWsnPnIuaFwEtI0TuQjAz2z2/jAoEDziiyq1
8iIckkHPigtoin1sRVJbV7vCDZWGpOpmS0C6XMEQp2B90gNMusmGJ/mLMgltJ76v
0FIkP3Og9JdiiGHJmGIO9lyL/myOcuBhpGtofpGmJs+2Qz6EcByKNMpK1IgM7+bE
QKvUdBb4Y1wbwkfjjKjm0IEqBGvIwTYKknunqE2hd59EFS2b7JEsgQXiE1oZ7YDk
TERKcjUl1WzXNIelMp4VGAni+Wh31kc0P+T4+IilAiwv8ozDoI+ZEroQkRK2RA2g
N8yUcpzagejv8ZX9nRV7rusanP8Xk2JkVXvdvQ1ZUP+ADbIV6qKjFLce6AdsyHrR
gqSEIefKTpaQgUSSCQyyD1XAwkm5VyRL3O3goZ22Fi8CUZcf0bDt/mGx8sEOG1yZ
OWuEsASRzX6w70LA26qoPkcATDZ9B7pFqfesHIXA0OIHbs+QWVr1bo3776sOCljp
Lca1dYVfj4/0Ns9Mna6ZKjFlrtNQGmOOuJUtoOidL6/Vk8mJ79oMOgtOnChyZJGt
Ncz9quITzmv3wxxqIKOdlQl3RATeAYzM7yLhrMe17m30YKnW8bHWBpo0G6yOs9ie
licQeISphBpOmKI0HSUDPVIZhfzrRTDs+G9J+XoOUkL+jev7199ArPXyoEBbtP4B
GYKKYNGi3lrUz5BTno4En2733KCFhXdHhr7oxQksAb3tEHKC/I/Ttwgcm/sgW3Sy
JQsiLtS3ev1vgYJGc+DKOuKs+6vIhwRWMKhQayWWbLJWZd5RVkEPjUte/Sudmm74
b4jI6T5M7ESFUIF8fPQxWH+sbudiKC/mUtukSz29BbGevdqdVhs7WUh9vSPW9cOa
5X0ExUS4J5Win9/EEYWEimQXPPYtjd+AgakIatDOwpvhC/3owrsuABeT1Tk6QGGs
/A9w7h7nKCVK8KXbNnM5kfZuLAWls77UatqX+Ef0EWQ0Cq0e5c5ksAAkrisBhAsu
VCHczlGDeOB7IEPq3P/vbPzNUfyRe7/uch51gK5cUeBRJenJb7vOq13LJ2ci91O8
h7f3yXbBi5q/RW6FIF5f43dSPtPCqg+QSaGzrm77iJHt/Lmk/YK/BoPzd2FdfkEp
SD3yFZVutoz3mAoqylKQ87OXCdLe2xm8aLLUtANMsY29CLFPPtLCYQnPXJq2gKF8
zXSZX+XXPzTAdE3HvGa3uW8iIuBDlxGg/109b+oK1VBLG2qDKQr0wRy+/EBmaATK
TiQdbWiaMTZPiT5sELGKgcYNfa/x6B77qgwxe+C7yKf2t1LbTmM58U38bf0/fF2n
i4jTF4DF7F6Vq2fLRbRORZqv7f51B/ED4uLVrpYdQu81JTOcSuX/kSf98Y69pyox
/bduVqn+AJod6TQ/EfYKG3zLaHey2ia4+bKAVdrQKYykJV4sy+0pzl2Mtj4eDsFt
3+7vZctMvralO2m8KXqqTosrWyicJy/dKCYJ9gI3ydFeQHCZQZjLvnsjOGUg72ck
HxHhTuXZO2LQbvBy4FT57k7pQU99rMnuYjxZBIyc9wc8sxgQVYKQeiMIdVzdDrdc
WjAvCIutJ3QTwHhw+katQxC1sYHVbYbIeuyj0Ltrl66sMvsiBYmToGIRgjGha077
BJ0ZYdxqIX16igqupMO/GTDE1pgi4ElVCPpc+UE3btKqslZUuH+pbSKbbC1G53WB
QmQJFWjMW9aJQKz/cw3H4Fsr9DwA9zsaYzRdMtu/U50w8MzxEjxbBRu7u4gxla5a
DvCQfw0SaP/P6xMId01/upKGIcPoHOlMZJTDc0FEpiyBfYPGwUWmMmFR7tUaTlDT
GYDAtgmyCi9wL97l2PdjEfzCrTVQjEi5BuWN2E0veWQuH5W23F1bW2OoOjzeR8Oc
0qAjyaJj//dzzVAF7RjWsgcH9EBPzw8kkmN/50nudtNWdjDPFWzuNNcxaTYICbGR
D6BzbY5IDym91LI4Z2+mPXy7Il7XbmxbR2HHU5OMgNQXLI5Gl6pFgoYgMQyLvfcM
iMW8QJ6gB/m/2q0QVGbvxWrK5zHE1y3tR32HW1jRpAjLhn5tj/IiXI86fDzVUOgL
wa341vy990LjHancYC1WpVrBpU8UAIFCHe3SY4irC+a27zXUc/o49AKHB+L3nanB
KFTqPRlHpJ44UFywqaV4dEvfMqKnNxjndRb/FFCnKsowMVNvNMuvIENJCL3CozIH
h5X9/7dvClNPV4KME/oTmejTauRh5ktlAiEVwzyOffH2/6D9D4hraV+SOqX9xFKU
IT+08z9f3RwTL+UZ94pKBAAM0C6PLXFOLP8ISeDmJVg0XoFFnC95yWS+q9LqTTek
rkuih6j8+uaV3h3n0AN610Qz0oKcUUR6E2CYAlnp8aDCbeMp/e5/F/HkZ4M0jqkH
p7SAQl+Z0snVVr0dk4zO0g+KccL4HOAB+dSCwFJ7rsxpmAp5S/hR6AuT3b4TkTtN
Iu477XRrhIoXGuRWuAMEor+ukxRImQRJkWwom0iYiMPP+7nZKdOnVK0K4S2AeEVT
3qtGOyapmYrHLVQVh2fXLfFrZ4f/K33CZ9AqyJL7XEg7HnDpDOqDQS0dj3OnJKOa
6vls1Pai/ES7Fo49wdv85t1Vaw4GWZufFMSFJ4oN+fOZSoMLchSqZODXTXUBVjfr
dm/lWCfDN/AuuhlHcQD36yCu7mIQe33RAWy3bA/21oBdliiATpeLBxxzhUyaDIPk
GVzcvXgqKF6anWK0MiehKB4ldE6JNUV09jMZSzDue7gPbVTkdx+bqXbWSklwM7mO
uc0ncIrn9Zu82C+F3xR0+AP2NLEAimlEKAXrVxbqF0CSPrT3qmyLkCgqiK/vq7nU
JElLzdQFAhIOBgRuqswHomZaD/uilJewpxSLPtj5PSYOJOljdrzAe+U1veppy0fd
Doxv+pf7KYo29mQV87BjoEEkZhVTzcS1fIfZWM2whTjdjBYupQy7kHpsIEaAl8M4
ggMUV8jRsL805VuJ+6FAHVOfE4s+8dDrm22TZ6474kq7YSzv8CstYJR/ktmUnKyl
CWj+scPhNgjQJoIAUasQigAcPb1N50ktBkVa4xSxd3iVFjRecnIp+4D4JICQnriO
gln1DrZe+ohBxc5STk6i57emuvNhL6qRYaSSbZTA4qBxmekaq6TyyMdjaYXHuRx1
Y8MIl0owsB/toG9Z7nKtlKnUdxYxrKSi0ja7p4fYbYVfsX3DmU8JDBcytqv5z0HR
+EMNsn/DBh8GHduTwoV+WoiW2KP/aJc6BufScG1KDQC/Wi7u3KXRfHsW6VxJ8rNu
yzj+wr7Ktlhn4bPttKTIn12Muj1vFWeiy/YkaVp6ohksYgd+spN0ZeCbOWFaS6dH
VWKzDqtDkcJuW4Uod4POrTFG8aKMBtQ1FS6dezo6d1kEMcSJXAh+6DLWN3ueGQLj
uemeJNlvk1QBpP8eOnvTvV5N5MMZILtFABidtIcSuNedX7AomeOHcY+LgbmbUDTA
nJpDzEGsjeTi5Ly4yc7qg0+DzytQ3Ec0D4aw4Zl9v2guDUk0F60Gc+czie7WVdx0
FRXJ+x3OQuhhwwbEDXGdqzwXOMF45BGISbL60000LjPxvNELGbtk5JzbiIaupCUi
2x43/cVvMEXuA3/5We4V7YRErX6AMybLB1LVcmiTq42ISRxD1QsiR1WQtzBmfS79
9iXK66VuEZRxE8sLY/jSprHkvcELgTogGuyb9AHOwaNjD8yWslorA2WXW3jZ7asi
o3MY83QOxy6L89+CbUbhmOkOpAovx3syw4Q2U46vT/VY3hPBTTBs08HnoT64EZUq
FlRv8Cyd8RVRNEnhYAQQdGW1ArvcPpw0Gn6uERDv6JGP9k/y/GUk2fI4v6jraiew
MEGC1ASh/llOwy3q1iobM4P6k6oY7UVmjkzYiiOW3mHAgch9kStWOgBDCV46hFu9
s3848ETwjcf1HY6ieSm/M8Eb0hWQhygc/CJso40jumIzmOoKpbBIoGsoKmyDl7j2
edUHbKgQIQhwkVMeAp/FO9RueFNvtDL/CU+scyNaRf+Ym284ioughKRhfO1np0ci
89pi/mjQyvNtgIskK49eWj1k3BwvwKL8i26YLe3C2HDdkNO8wKfOSvg1zhe2T5BD
HwY+IlEKqGU6NyglNI9PlqtL3WimtOnZ+oOcOwGnSStZ4Z5IMKf0QboROgLcEhzu
fMBtbjzQFucYvte7dIjYXqs1ESDCqlgpmGVTXx6sO7c2jWTZ+0n9g3QzkdO9zBad
yie4uphYSQZSxtFJ0OAFv5Z4IW/Fm98WeqAT4fRWN+uThuaKznE8CE+bXIjFV892
CBoFJLKdoBLyaG7jAQmtH/sQtDwj5NDxBKloWwPG4X72YUhMqoCUllSgH9uqa8cp
iTvEmrzBdnNuF4dkCFeKutatP+5hZzRY6L2gti3AVUNV9XiCHylGnLP03xAR2BUm
PiKigVE56uNkpDlxVOTUXTSO9RmfTJPwaIhoCM8+/HLbZqw1fXSBkHb+AMgImFQR
XLhOnR6xXCdlwGfR8DWi+zBgqeUvNCngk2KG/0yjJ/7Fkh6awW7Ru80tGFeud6OU
WRLbZRKJzDT2Bg7xjuEjH9/nGW/UlU9AADicRP3TinIoxYYnPL/Iq3ok8nZsF936
GDAve7WwHKVd2kz/4YGxZ2sFrWNHx+6CcRC7sVmDGOz3zkFptahAxeILqF7SSseC
Hx5/5X+VEoMbcljbQFT21iqnBc89Kyi0TnbOm4ta4kZrHrT6c4mNd04zcQMUObmG
pcXVCMdM4g8NCYSJUKsd9/HiKrh75eBiGbrZGE/RdicLY1nQJVsbWO9UWuL6akCH
igJObRsFJzQiBcGLVC2LVDiMS8TIi2tehQGL7+6+fPmTE//jpPoE1IhxRDr9QvCw
VWQAYOMidrKyyDtj8OG5sZrwH8PUlGG3v5lLgdzV9204V8bfNfeqtEuDhvIRyhO9
+F+mD0ZNz95V7FLcqMJrZRtEGwuvouRc/xDMpqA+GRN8hlgRgT0s8jeMOCzdzyYm
m4QTXPpHy45pXgeeG6OJFSnLonB1/ryV3P5lL73eg6TVqpIGEMhr1s9JBs8pO0Bd
Wdpxpy6+kXnjUjtzQ6mPiWwWA9SFaT1j4tlKRkkcvHgejSu63HaCwvfk7XkUOqr+
bTBHP5e6/mayBK1dpbI83KVsNT85CiMOUwD5fRd3hvVzG060Wk9EgLnOoWPnsUXY
4PZKVjtxOTvdsWPcySVzP+3Po4CP4N5PQzNqOZV9pwDzjAaJGro9t+8xEC2zJIde
Dz1B0No4mEJi5MBQ/WuV4hzlCeYkSaxfEIz4HFmwdccCMPStmiwQ3WP8WYYUiHwt
g++bKlRl+LsLHkXpP4WFnhb+Pvn6ASjvOhxjh+I/HjuWhHV43t5l6FNU27T974Y1
Q7MI4sC4itASf+mUE/hbBbHg21XpHZbxwWXtilPo1K3zBpnSdGgr6jcFORTfLOwn
WvUoeQwwhYw2tOf84znAmrGkzJ0dBXeIoXU9B1U1UOJENKdGCbHX3DoE36ybB3WJ
/klhp1tqKhFFutyfH3BXHvemwJrkyAc526i9HoFWCzrWbfiMix0/q7CINbO6AuH3
MC1WujF3JkxpkwH8aZKA5gHID0XpIeqAZFdf1O0YVZTBG+ZS5uSWyIBz/WxNH+Nu
RvcZsXwwX8OG95Z/2Pl+CsdqC1DXL5uIFLFV/1SN9oZPhsdWt1Q1hmtW20A29LvD
x+KcsY184YOVWq4IDWSodSjELWlraFCe/jgayj6e6/zuHvkNsPIzRI3GAekjN6tS
IPO3OvCEmqeIfNQkd97jn6Q/IMhMZYbf0Zt+85Ulpxby9kthYhuXTGBqFQs+avcM
0Q9mj9WR2KJ+8/yU33wTCzoWLc53tXnfTEGIpz0D7vTLzSMBjXZUjxaut1kinCXb
+NQ+LtXUAmhtubS1xoW21kGtBDbuQlJ6SnftxtQprvQK234i1Y7ANXVZ1ToKTeAj
sQSVBRqX8HhOESs6iNBcSzH7BVZT+XdtUpMd1Oa5HZ8LgwuPBbo/xjILbJ1AEH6D
2pIWh3BNB4WPJKSEx02uP0qnT+UEAkxqghiArUI2AIXJ9Syxn0ZGmW35EztSKeL0
q5QMBvxSb+uZZq7HWRRWYJuh/bCm7VF1VGN1vPeU90k/LHWlzCajA1QUrwHTuESc
WsikmbAmJhTItEkwVMiu3wWhUMZK0ycbNDBNB+aog5j+uWxZiYupXrnWTIkzX3CP
b97uBYwbZIz+0mWd0p6ji2fv2gILhbPDJjIcEiKK9Bs2/BnG0T48tULlmAU/htx3
Pf016G/LR2GZYuCSrUiN2ZDrgSg2BNGfqwnVmNcsQ14ebVDpSLCr9VoxE0mBwDQJ
HI0oOSd+UM/nbC7mLerMko1BXMu+22WcLxQ+IDYfMqOBtHJfKHh2xM7m1aCOq7ma
wZ5d4wWf8WKcZDxhlG31SUCVYUx2HdW+1lx0c7r2lUuJNh7lX5+jHjZzEEhqRN54
Y97FGdlpWf2BMg6d9QWzap8UbLC4n/3KY+qlM0vF7cfgfqI8+9oO0+gqrX4Gz5xQ
Lzn80FHdQHFrRqNq+l3Ud3wSf2NCF1WL1nMKcRpgBPNTBT6M/q2OXVkB7m4CE/P+
D09YW9b+J5efrYm9Z1HCduyMCwaophaILHf/Ahv/t/CiqkyzxDfy61QoVmkHJepN
Y/dAVQYMdI3wNvL1ootyCwk4hkQ/qQixDkoTuNbXZry3LRfctZZgCDcRsdqv57s9
PYPWbqaSHYKKhn+9FXNPMsjvyWlSzsFC3EY/F+6rxApCAOS02zA0fJ1F2yXvf+C7
uDCr0NQ0/NNqvmFLga/pzdhkMt7N2SidtjYJG3ejA6fa6fod5/4ksOAY0cYl8U8X
KvaotzwbAU9mCmNvscXONNXb36+BiudZYFX7fPPNtjwSkyaCu0HJVtKY/2rEr3Sk
dlAh4Y/3+Yz7JFwulp4dmdgvl6MVEaepYgr1VLAabBT1OSCXkx40Qe4zSsXC1bus
K0WLXuP63c73ER2/++N4yCwrTS56tQuvzQf+8sZGWO8tNHpkll5B3BBKTau7a81x
hAPaLIajSxEb/ASQmDTCd6t5gYY54qCXqKpL5RwMnCntZ4Ssr/Jg6XKp5x6bUhQ8
2EBuCLoZ+9ntBMJFeqWzYz9FEzHTqB0iihyn31OEMbWRCr9Bc8z45s6wpPKl6AxK
zV5qoTUFjdbA/Nag8bKbtJKQMI/7D+N30Jn/aJqeQUG4Y3M+CDZ3m/Q0UkBNyXad
nhAdAWww9PylmYN2F1IS3oy6cllQe3NRtpJ7Snn9QIrDY3tw80tfisWOo/cZLdca
JVS4kl2KV5mUj34lhx7Yy4jbMEyszjZF6fKUKfhTAjn7GTXWR7/B6RQH2+1neTMT
s3s93mUdkmFMC4eqRc2pdo8UINANGs99Dvhh+mjHZk75mSy2SQTJ7p0QbwQ5Lz+Q
o2nXHTUCpKWT2xehez/edbEHxm73ob5EEbKtkNhvPrhI45j17KQA0zMK+17UguvU
D7sW0nQcS2Zkq2rRTp9C0NGptXUxfb+pbeRAtwL0C0X4j2ADEF/w7xLhbF/PbrIT
/AO+OWt8Fp86ofGq+uBogh8a2HhgqbygZv+OXdRBX/HR5lTurBVZ/rruIAG/ibrO
GcBtU3r7rxmpKPfysVhXuw3SY+brMta/poUnpuGSEwMPYP9/v1zQmXGlYhZlKoHJ
ACuvUEXwHQnXQE8bCDeQekuvwp3oQtMd+e3ioPEZSkJjmILmFwa5Hx1e1YAajKQW
LhJ+r/YSJfnU3NnENvLPunQUN6SpsrferwE3iWgu/D98yC3eWiDkIMAEwu9cDTJj
HvzumqzAeBzgFCiPP8IErPm1NU7UdfKVwV181rdVPK0Va1MBoM5SncziRahDjFzM
g4Cg7Ocy6jfxKXkn1YD5dQ7w0i7NJGP+yQqeE/pGDVBGiTk3LMo6bwSxs9fTbRFu
dqiLth4+f+IHNNugizIbryRoCCtmI2gu64r4lydiuZTSx5xa0+yRB1B0sm9cPFVW
uTYuJ0+usRgpkLY50cZffFnx61+qQKJu+r+pca+Mjy4h5HZd/xKYOmu/3ed4+w6m
aG/90bkMEG4+3igt8wnmxg1dhSYpu2kzAtTyMQgA3R6mxGHZK57SfJLsj0j0jMBj
OF009y9zJdbzlmsngXPiofuJOCrq6HIvhs5InotzR4aEvMtcTLgKuosOmy0jrbpd
cSt6A6TyCtsBQwwXLBvO7YFuZbDpWlH0Jd6pGt+oBFA2TIuMO2KKpfiOdLepFDyx
y6ap6gslGZ/azNwlF8xgRG2hpf86AOk8dk600e27G5ZturxkYA3dRjrw1WAH098s
RtovyiBJBOcr7UisVV4VOGzaqF5lW+z6u2uRdX0y3D7SF72lzngeWKgMGzwU4c4v
vL3cWmxr58IhKg+C79P4gAufnLBkZzd3fmSod/sH0a8uTZeSXpk19wFX+BZrlVro
9DPC+6dMir9E3jHxAtXjKbSAgoAKr6hdNF7pDLAU1MpuA7t0teSTc9c2AhXN6owS
IKkkILoIGkb2/FLNdDgwTO6NNnIks8OFExkIpdIJzW0EpLtpJ0vlkpTgvKOvuSHv
mPocFAkxkoxL9qL2pNcR8IfwJ5V8KwbneqLILyQxCbJaYhpfum5vawl2ZXhAmsdx
6CZcVWGynzt0VWUrTnYpa+Obe9mlGJqSeQ995XTIFnknd76l8rAvVYENULip+4SM
V0Ro8pbhSJwz0naP9ml1YmxiESK08KZDNHRKoCa2/QwVwAuuwBckCskJt2HcbjhQ
m74kuEt/mBBaI3FQcZ+6vOBNp9vrww2SADIt6leWBjBlscMomQjTOl/eXh4QYhsA
8cyxfwrldgMOjm+KurvST+U27VBbD8+7It4ithEY7lnGXZpUEsdjWt0u78dkdVjf
/mmJaAYBVz7NGEsCQX48YS6I3SYKAm5nbrp8ZUTnoGWXPRT1N8Wi0w2ZSAI6zEpv
J5X+Ch3/vySIbnLLOIQdCWffDmHEJW7zWPWlUia0IVRUcWLMjbsGoD1GnA0WrmGU
FBBO9z8HvF4e/xv3SN192OedrtgrvonuBebmjK1x1o6ZKl8TVUPqqE4xul2wP6Aj
zNsXoI74yb8+v9SovGtZBAKxwrVG9wkaP17IO1UqnAdL5K/PWxMWrQbYW2kKfRhv
3ODnLhe5HEc8axxlcP+5xrrqT4wE/D4e0PKVf3T9582y6rRWCxSeSO48NiR4qfgb
OQdlC3T+mKWZQTaNHrAxT9fpNF4do6EU9VMIcC725674W0Eaob6LB1Ez2saCA9ep
tDZ6DdUdpfQdKaQakyAsd9kxrYqiWBfXBMFF3EpunEMkfTvKDyeFbzLbZHXCkZjf
F8Z/jc4u2rgTD+JL3LZ2Vso/SYtTs/m7wfqWAOc6Z2V8njAYNObT97pFS6tptN2F
xxFcKnNx+CHzA1ZKbQsOnGkYFaeQocPhnPn3mY5doDqJr3Cs3IA7O+gBbaw790ht
Z0TJt4EhdZZhox31tGc2foThgT80PurUo+VWGFFaK0AP+UdiSDNlzdnWiU4uJ2ax
IAxoPfUf8rPZcqjAPSaHTz/je4uKEBKuuNZNvKjWW+CLgi+3LLrdnf1uU55odmaI
P75Hi+/yezpza8VCjHRW0McK9k1aXQnPKVf/e7ajmb3qb3PrQ8U8onTDpJlTxEip
Vn4NMpCfuQdkqEAN08ob7EDZAFvDPj5SkQM++9g05xgpbXsou39driZdm0rIwlW7
nUpziqTq/OC8MsD4RJ0rJ215dVa19QgM/i7J3+So8/UrPNPnEW1N+zwkz4o/ZnAj
tVaSx2/oDbeTOZfZrua/YK4r3AdI/0HryjAStnD4tTzgvMw83WLyG3KwZXhtviBC
S3sfdeG3LyyT+v+4vqYQCNjZ1MfRSQQjbNVCrEOFpEoRJ9TcYFM9V/Qb9+7LQ8sU
U3xQfDQOVrDgWd7OG+JKp57p/didn2NfB48MZI0/wIbN2foU9y3GsH8kz5c5fbWG
6SL+YxjBZ3as8uEgszcU2QcowBf6nHxzcjpsx8LWju5Jjzl5f/+2hEaDZxKhzNph
LAPg78YqjAPwiHVwbETi0ZwF0QKN3O55v33Qqqv1t85zzeTmHqYIbq/PNu4lmJrg
hMXjmwmrJ5togFSLp5iavCOAVwrbhi7HCaA8LR3DI2cldrkrOdHyo0eDuwsB1buo
7aZHzMH79eK3x2yOD24va2fKZDlHyhHZhBR5QC7Uu4MB6ffNj8k1F3KDDBE8JGA6
wSnhQjfcJYpgNO6BxBJlJOSayEp8ATEDdE/UT/4AniOni7dfKU2axmvwnGYOn26S
e7lxK4z/o8GxenCq4VsZqAjKgkr0k69ooXAD9nWY2c/d0AnGnTSSGZvzKrKfslKi
XUqd/tKuFzA/IIEv1Z7OnRkeT1boUjc/erOG8th3Xu0qAmQeJrpJOW8jKV7ksd9s
L5RyiVNj41+5nsx47a/HgN6QnX70shHbBwpCpMSQB1VTLjSHTOAYL1Sr31tLALef
BM21aqQOzC11FLmcdlIuL67ryk0sJExY3UBpOrMitAo28ubCy8f0ir4F8bU/78wO
e/u0k9WeKvwkXrnO4HWwgdZEzCw2Qiy0s2UnFumj04uiKRqnjjtpq3aid8ZQlVyF
74TYGUz1KKO2Lcr3P2JPNDPR4CPBq4M/qhYq8Fonmv6VMd0/L+iUaVjyFSQ9x/GS
MoTnsFee28pOHVQhweau8df98El0dHFlDsV0UrUOwrxWOuPP4mbZ0ys0BDYQ9vC7
FYFnhRWgw4WaBJnNu8eRVE6pLplRKNRIPEBS0dfQDLQZymSf30f9DoGnJdxbszjf
v1DJc5XFSYk8dKD6TMqvm3CUoGUSasuMLwIxPjAzRdvArPQ8rRWgrYE+b33Rhkg3
BLT0oml+YCYYiB7db4YHa8jCUtYHIK7OWHXRmgaZBwHidgL6PVfkySBkx2cCfxCa
xQRN0S/F/3oJr7vsQx/lxXgJ8HfFrUeLCFuyu6gbL2QpIEJEyJj6cDt1cApoVqAr
2zBay3AX/bRvG2KLmNB5PBplhal2F+lFMSCrtTrHo0Uw4/Pf012Tdkbvnq3QfGmC
RF29WOjyUXnnOgfvtEJ7o1UNDp3/rc5NttHSHioNR/G4h84HUJFgJoPi966WT+OB
K3ll/5hDxXQlwVS85aHvIkicX15hID0YGGQ2oYrutd5RVo0hmyIcXjog5usxdTGU
qBcQwF+yvoM/8KmN9LHFQI3Z7KT1plL9aBlOJHQJas0sokW+ycxxgtEBBXJ7EXS/
BN5Svxta3+kyHkTPbHhjxzjPG41z6cA1g4nPA9daaF+nbhuBUN8SKInxmfXrPgvR
Hzpstq3OWfK2Ke+E94rVbVpzMcxFl7F4Kz7m3Jp7i4WhPKnNJdZDgBs5fahGM6Nw
MqBITAt7RR9EWthD33xZTw8qkUAS5Qm7SZLHd7IiZrBSzuygR4+hHXbp/7yevFLX
8+E6tRLIFGMS/x/GlmY0Nu/15qugqb1T1YcqAJ+I54EgmSSrdEyYUVdN2JcGT1O/
Io+22I23VmiyX7K4et0CO9afBOh5Prxf2SoAANYieqedKdJ5MfHPtYT+1aUo1hvf
+H8IFVmzFGaRM7WbziEAjkQ5599omnD7L7fIqxG7fQnJousqB/L3bmIJ1mti1/XY
2NypnmxKiyETuHBA/98wc3D9A2Bwq2vXF0wGBfVTRFt68VNKopYSYOkNbXqDww0a
8ghOTbjDJdEg9YKNkKO4ksijjK557+XalUlgZJCDVRRnWfqb+MFqcRK19AjHowkE
pH0ykymWl20zFhf12hpXwnbB3Ptw6MuXJ7YumCzfDy2DG0owGBIdB2wKipKNCnuc
b9p5IQo//zqy/cFrU+wI+Lk/EsqmvokgNErhi3ZN0y14AcfRzMR3fcnz3dZdL3kT
lQyYJjv012/E2NZVkayxh3RQZyAhbQej5p1HKskK5cLEGSay03aO3SPw4cHReOjm
pQzz7A0wJYhVjsU8P8mzXhc9nZIYkMPl3CFAavEYi+CwwLyD2LoVhySWJzUfGMwR
2GaimtU6674btJD5JBPPX9B8FIRKcneEMr8UUNYkKH08qpysahpsfkj8DjvEekhP
mWKpVCld3o3YkiuOKyeJho3uYkHXYLkqPLf3p7abBjrI6OU8TqrvCYpmWbXpNaaJ
VhErIaWsvcBzJwr0G7joL44XM+IBtTX9qrB4zzCLWajf0Z79wbFAn0jydGX6XjqC
glOHUMU2Xp4G2C1shd69S5EInG034BavkBevoO5RoYMobEZ3RXfyDwO/DOjSiJyV
uwCacRLJUbdnvG6yCZdkZdpzyTiHKUZnos9OMdX+Dg/yTZQtAxxYs9pISRqZ07tx
N80g0j+WmbhoxAsAQ8/cHX2Nk/oSHR8ZoOqQ/6RVZKCC3hHR3spyp5Rj4OtUVucR
3+xRi+3srhZTtS8+W0a1QVCLt0iBaUHoLWEXSTwKhCInApMk5N+7qTXoI335Vf2u
Io/9JLxX2121gmcC/X+RbVWJrqr7LVbo/lar+zFT/v0hTeReucKcK9kLljDp8wKe
k3cW7YCNdDSX6uOLdyBBV4BWoQcvNC6djLNW7VZCIwPepQsGEbyhSEAp9aXfjlnY
qTWxzLKFU9RVD0KMWzbSCQ5f/AhODRKLIycP0IWlF/uoSM6h8CshW1ARJzjS7hvF
yoBXPVz6JzSebUQU3a59W63eqSuS21oYIh2A0DTc1ewvSDdqqieO/ZxSzqryUX3X
bmblmnILZaL4nCEac9FfH4BiMRq3X0IUuURR6lxB4gwh/selv6SAeJfZV7bgoYEA
a+e1hIRDhjNhzmhAOIOxPCZiZpw2uG3bXxsfH61csfwBcSEJDUwPKI0jAHdiuI2b
vveI0TdOIwViDBXYaVRqbwzk/0Q+W06dkdcl8GWXuJ3QrYOH+awIuA1O81gyQKjr
ObVizYTXky6lCpLVyU7TMziHY1z9v8aJ0pjAtSqm9VHTrq9AR5chzGPpaG+sT0dY
0R2bREysn6OV5RF4jPOJKy9OnLl1KTBDiEoIVup6WCK6ytb+8B8Hr3AZH9vDO2ZW
ONGPipirCQBFf10o+UNBWYgSjc19LZeXBh5EjwAWDjm4ebsVm/+CnE7+ZpmhMNW6
r1zOgXxbv88IZ/GwoO1/l2fNB0jETqfxqHaAiiR2b9kd9MnkWAPRhhNgyilD6BOZ
2fT7SF37Sjn/OXijwoQ7WQMCHhjbjEss6Ercw7HoCZ9hl2MoL+Tpe3/ey0EI/WY2
CGBxkmCZesYxSDoP4rLROBzNCvXHmC6q0Ql7bLQTpy7Q4Z6Kyubvyu9TRfu9pCix
hj7QVOuZf93lJJ582l0nwGfwmIuXVJ3dT21J67U6YMnLq17dPFpGVjyI1EyIPjmn
sZms8BOkj6P0mFFny87j75HYEDMhZpKwpTyEpCdl6H90Ako0Eep8eUiDesAvb0oj
1uadgpNX3kYO+8gHgJdqEAf92vjC48y0FDXWD6me0l1bttr1azjHed4YywmUqQDg
EatBQtcD8jb/NdCSc07OIk5hpmTNjZus2E2ZBzRLkCiN51Pp2cgM6iUBCng6g+1I
9hhfbMHtm7RFJLHOeXdowDzz4lcJe0kesgDhb6n6jdRpyyYDZIqkyknUvyItwzr6
+yfTpDC+uDyTJHNFxh9X1OuBGYoIg3JSWe5Ye3NZPSmo4phA1OcX1xD4uaQtgT9f
/Ai76jkW52XWPplqA0pSZf8bkK8s7edWBqINbJkHQtOIz0jLNhnqqZVCzJlRBqO/
6QEGqAjmkbeezAbDafBzu6dPM4fXr8pd8mHs2rKnm2QP9CBL9EFS6WWUbf01kCKt
j1+sclttYOzkmZvPXYv5tnU/co/KOyQyIFF8mBdyoAXOvn/Ssa/SgV6mHGnsO7Ja
MT6Tg4K9MEOZEn9eAcpoVcQREHV9YjYiNJcZX+Se/Vke/nbnmn46Q4A4L5Fetv9F
3sm6PNXmaDCuinzwxqzJ9Dje9TJ+ZS8CtjPwSnYjMa7XqlGfhNVcwyQ2nIdQ1+ar
P9Jr8n4lwdTTVjfByC2MmQ3ODizBHfNEGSrK2Dcqans/ceok0ZT7s8shFPU9gbtK
uo96vvuN15B6oDedaa+1nmCB1nvH9WgmzFUE9BsCBY/2l6IjDVXqtZvgIY1rapN9
D33kxsPp0eNiEAIMW8MiMbn/AjN6nQVwp9+3ScNAndfw7wq7wYdnfdiZrjLFqnSg
YlJlIgFrqmwvIzx8tYC2KPTYfPRi8TmdluYz/I5dzlSq3OQxrstzEWq+xfd0gvge
Er2/+uyYW30Ibd2jdhnwTd5t7NGAdpZoJUUCanmWgaRXAm0F0AAaZfQHZrFHnM/h
INwjJ57qEHO044aXMfcoeTNSTdV45xOsSLHYIX2dCAvIWTIfonoxTJs4aZ0F6cYx
kbVKQnisMvQCPA94p3bc+k45fMVIMDsvdmr1WdASulXTsu5d1S25NXfaEuu47SCR
aFRBuKjzl/A4vBmLPo8K4B0Q1vw/YgiHn8ghLCLyks3mWfF7FOoQNtxUtIBn58Eh
oRYFqfeFpTSyfV1cpD9vVJRptu9mvLrN/k5p3X+EJy5AkyxCxyHDOvyLSjvJB8F9
1oS7hR//R0NaqG4fZ7nmev0JiFo+Ts5oU6HO/clEFdoux4nzfQCV4lky6doOuS7P
ZFzTYC3fVqYB4TX8Wp/bMQ2UZ++tORihahzH/DInoN4GJfghjRv1lWYLXpkN2URo
6MaWoIleQl45lhVz8n4YafzCvPfJkj+9rZ/hjTDwXWQ4AfrmGtMKnXdmdcpPjtDn
GQb2dx2NpcEisScxwqNVof+tJKZNBzQX+T3DTbnm9bSo6L8ARf56i/1BGHtv/nla
V4WD4TugSV98Ql9AgYRLRuSIAqSUdr/DutvOwRiR3Bq7sS1bt3IpkGPX/itMGT96
6nJhGrbG0yu5WolTZNoMziZ6TxwYQerTNumoQtQCUmh/maqUP4RUSVqQ7+ZBM38O
2HIdLL8z+j5fllCfJy2cVj2tE6JIb+6IFVA6xsOfTvQwuUc2eIiizS/l+ktPlWak
ZJDn9FZ6kRawmFsKJWfczJer633wDiw8nWXRPQrpywb8Y3DUlSQwXvTRjJQjvq40
7aUw9852GWaRfClfTscPU8fPhGL7fSq9dJHnbEgLS86wrEhOCY2omz1U+nwAXKoB
NMESiRW7NTCxuE9eGb4Ssax//ljA6R/cKh1ebGtNf8ig9Q7Cu4E2iD/vozjfMeul
hkFdzUdrkD62vVVuyxX9c1sgMue3fY0pGUGuA5VEkMk/m+xBHnvWp41xOrjBmWS5
HkJ7MgK1xugBMLr3ynX5BkqEmJJDUA4u3NlEMYL4jfUp+fPbp4wqFjZ9PMf2Q64j
EBEoBDw2G4hhpyWjCZfPe+QpByhFtF1mXLw8aLm/RcxMMN/riSSNP0znpbPMDVCM
inK0yyIXEOGkGbEY4y9NIkpH5XNdTzOuLYSqmPWTnzUNwJlgiKcPD7D2sOlzC1KF
Qkq2y5EXYeeCh01DJqbjf4KW980CBX90jTqM3WCf/6PwSm4rCC8/7YWTBrmPGA50
EOokl8Kn8JBv0ZZixFdD5Q0H3UaaxVk3PtZmK0eEBO8yZLeRSVCdHSlnPG0d19xz
wMWCo6j5Pxw+0jugPcDxD8snnH07T28f7MJ2ciUjWpibaPLqOHoLmykntlqA7F9u
x4mYSuxOxrgCBr4Lgjq0A158jxqAyG6D7VNcO3ADVorU2ORQNqLPl9HEISivka6m
wvT+VOpJ6OrwpZh5bl+Ts5nCQY5Cg4gKyoCio92/iH8YM1Ij9Mm+lITAUb5ynY6B
yl+2yI1HQCrOtOynQZMdlvXQ7AlH+bHIgp92fhkAMNUzvYkCU6oUAxVsUBIfQW+H
R4fj/9rpS/2NxzLKwry/kd1r4L/sckpC5rjqawMUzvB1ZaLqG0bcrzxNQDQ4ENsl
8cqfOZMx83ZIVi63amj3Ki8GkYtvUVXJeZu6dIucy5MCagz41YTEGyqKGb8BTL7o
nTJjOXfTOI4pI0KdQnSwbwGRez/cItV2hyCUF+urLY2yxooeNxLo6DABulovANKy
w1bNtcdLXPBO8k8PXe+BeSbY0tltCddaxq/abOarC6OG58/rMI4kbJjCyCULn5o3
qHQwMfwhmvxxH3ymNCYdTlofAtZD4KwbLHjY8j0JgFGARGWiDfIU9WKE6CJS/4T7
wy16CZF0rLyLlVRVqoYUvXkYUdyjlYGG5cCOE7TCGj1zpY3NXtY676bAl++eEs+H
TGpBDD1JUXzhIlUL1fz/KVf6PxuTyBSIVKKj9MJ6IJoDJhGvGq9jRzp2FY4oZO5j
fnd08/Y3Dlw2BTUzPesutD3SIid/SDxY7SX1h5oOIh+skzjni3kOj6RnqtFGkHAe
Hv1fmlfv+UpCLk3V9rL27aSIHEM0vxo2g51r8At6MFzCZkFWGbf/GBjagfuwpLyh
ppnfCCL2Axa/V1BBMwyLnLl9kcrqv3AgVcsTy5Jl1l/83pY/ZBjGJ63bcEfCOj7m
pem8s2KowRXudcgyBYyizQr60N5DL3m1nTRAYOhRRrbjl4B8o29ZE2G0CuOcTPzN
ntqSVXs1wIrnOMvyuLRCfIOUMqt03+TCklrGlYbeU8CcJ8VFeafO7VMOdbiUIRYK
oipnSReF0Kwdt/ZFWvUv9hGT7eIyguABkRdXQzbqgusvh9amFvi1OtsGieKHBNsv
b8qc3YcspKOUpumnzuyIzRq/WGn5/kcle6RIFy9bld/i/RfDFpfO9AuBtV+pPz3F
oO9KaJI3luIRGa/wZO3Cl/vQSRajlvZy2y5qL48LYyyFR4GKMGR2ku0C3DkVIMZh
tr0+BtSYXCvsAV8tH8QsduCwYnd0JUXOU0rpk61kvLh8ITT4G4cT3yN8uLfBdPnN
EQX31Jd/g8Q0CUEfovOpO3ZNviI35swiQ9zg/JPX8zeBFkizX/vpdPFpH82k7bsY
vfiZcHa1RHokn40rftZlHM3aH4F6ES8sZz+2Xw3u2wp55tQFDsrfPjtwWcPtfc4X
087VnNoHTJGdKBmTXIIvPbapWvuDZMJnHNtXUbZmUODBGwVZzLA4Kr/CpiXSTz85
wwA2z5Z+Gg4sjUdKj+tAzaurXIdkZ5Th9sym/KZNl0+gqiOD1tOvtzRXZpGYjF2X
mnLXZCEzvufgKqnl5jj8S5CdOiUkXZyk/jAi4Kb+p7E3ZCaAQIcVtU9ABfNw/4pG
tZ9zc1qi7lom4zSUxaoODCoz84kX1BYsSZuu3G5e7b9vl/zX2Uq9cr1tE/p1TG4s
i5iXjscre2pEeEtd5lk4OkJELcG5epc39aSMn00hmvtK560wX9N9i6VedxKFEJid
Da3EPosUMQ7nLHayDNtT2vD5JzPqh3DIB14fPunmvYpnSPrZcnXpxpjjxCcNxl+l
gmbL+bdVmv3MAAh/R5L29RxShlfFZXlztAQdIm51/fakivM3J6wmVouY//fNqABJ
zlsAC4751LgXKLani3UUADZgkYIH5PIE42u3kChKLcnSFWINoe+om84AroGl8BLe
PkFqzewMYRpFR3O2XclqajdWA8mXUZjaVDqKyj4zYTDMzMCTY35IFXB+eF7WzPYP
owtuioGAHp5eIF9qtk/Bqx6lP8iFMCl8sNsj+adESePhGV5tFicAxN1JzVQdHEyU
ugqEpvYgvZOv7/E2/hn9pyesgwBoHDAzq+QnX5NbYsQJkNtHPpJ69S/k4OREuRI/
9wIeuiC+3Kr9pOD6Oi7cLSecVUSFsiNklByzVkeE7fWIRatWtfsfvWsLCfiCTjn4
u+VCKaR0MpFUqPkPkHrSAPfNoj8aE4Wyuk7pfSNdQuQxbPNHYU4BMitnf2XkHENl
FecaaMrtkrXnnKalkppql6sAISbF4vrwpkKPSniPVSRboEoTo455JyTvSd0x8PMW
nIoiNeqdd1XKPooGmYBgHWIhkMm921vHmuckadiSb5EkvsLBOLONf8RdfbCoiy+O
5aZQ6VOVKqSJC0JB2HS21xOZvMSm4F//C4Ah1lwSVme77Y9IG19vq/On3LXk5ONn
IPZcZy6iRwOIz/PYUvm8qFuH3ei7ywKd4KZOEKD2JNKeK3SE9kJe5DwmNe6ZsAsk
QTEv3+/DaiNjnBuitPqlJxuxZ9VqKllVyXKPjTd7KkpXTbfkpRNBR2/8yoKi/isq
dJZQKvF8C5LuT/ZFpLl96EVn96bG2QF5Y6fL+Jene8vw+lUMYEPSoMk0E+cUHkkf
65c3irbQezzaCA7YJxKF3rIUbCl5XYKle2YOHcGH+7a9GMY0gdxhJEEYGOdlqsqv
gpUe3EI/IOuYjjlR1KJgYRUdKP/qM73PbvQiTMMvHJhjmo/YUtMFM80TwubNUKWW
qS/mm+IRPWdEWjQR/C6fYYr+oJo9Q7H9x67zwL2qkgoKU342YjbhIU6GhBBkhUBu
JfERlNRNT+IX+N+Lk7xewfavL6ezTHlbG39QMfNAVq0rM/gayEqSgChn3nW4MwVy
gLph+YIzXvPAUTZwDoFGU9DTghp6K6AnuV1WFD8NecbkaEKgVOw5mAXegDhS3j5/
fLVxJdStzmNKq9aeofvuGwFY0hyh4WFGIpuTS2SDzoq4t9+//Cx/gKGE3HbT0B78
ZFniJ16khptlAL/kHfHrubfQjlZQ+rz4u8uss9MHYelLVvxIoq1Rdk+4bkh4KzeP
upo5dij6g76GFbbp9gS3kVLszIdh0ZJ8ssQCpUSgAC5b8uWL3pfFnwecZMThHIx4
Uyg2VMUVGZHKFDGKwT72WHzUS29PjWQ6rH0T+VEhpZR/cFtUq3XV1jV9xNOw8x/7
t0BO5u+KztVjadKwmgZ+kX3TEH5OyBvzKKNI/wzdYS82qfb+sajXA5PkwyW45KkL
atLL8dQhnSDxhPPxuz4ClqVOWueS16BUQRniZgw5QvVzZgqEoDSHOvNAKhXz98aL
m7EnOnkSoi5QFeV22kL5jb3QIElCZPQYD95XE9TK839tXVGEeK/67apI/lrohGII
AKubxhb6w1eiykPFY0veUWK6u1sgDFJHJscyjfpWahAlzdUofEoGs5Cj50zLug51
m7Y00hHf9xXAPbCq7pdJbXkdLeOG4jobSsZj9JOXOtN2sX3lHsFgpCOHUEGHfm2p
2XJRPY2D4DAu5ZHqUXNGxPtr0mszhK0uXg2aUPrO4CUIeobeW3UX1tmYkpHuxSdm
tpeLUcmS/MyCQl6SUzrxhNbUVzhng2hTZExRZWTfH2KRaeJLYzDs4VZYkSLq1Dmd
V4V8rizHhubWi2GVxO2Wz2ohscbIkE9GrvDwYtoVHbPgkvUVTlztFyeZijfj9Swm
Ldg+gZ+M92hJ5HgdAMy7i9X/TUuupZqIdXWQVKDCHjyG0oYRqm1dxeZeGRwxGeFx
IhqO5oPy27OWixK5eI9IdoGxHeLokCMpEOhW95Aswuntx2Htsw303zqNsh3AxaAw
VD8HESTMJe56vgY+pP/UcYIdrbdpV+eaMxdqMjzs7GSRdA53wG/tzDPI1YY6wYhN
sv7/zG21e6iEPjep3NT+dm7GxayZLSQ8zc8Kt3Cy0KMGIA2qPdvG3KFTQYy7yAH+
Gwpqyyig+3NrwM+i8Fj5TE08LInyHL5iEfdoaDng17WLpOTj5/yfGu2pUzyAIFgD
BG6Jyh7n9eEEwibdRLQHmVXJB5YIzAnXXqn3xqEQSLVBpmItX3nPu7NNyiZtUY+j
MXf2s411QrY6Daj2w1DeNaC3gRppcS916bx7ntjZR7g88lH9UCdldAoEHoXJsalp
hACEjXoDRTWLwQwH94HAAC3z3pCkH+LrVbwwIRAL+iActQarKGnQI7k3VF9AhVo4
im+N804QvXDBx4RejLgBf7i0dn9aXySNJIWMxbhQZ4IRdqNcQRYqpSD2x0TZm0FY
OfRW3rCXD8aWQLuhpgmSH4gIt44ZEfT3DFG1Y7r4034dAc9FegZXAJe1QoDZzTiy
8hQ/hNWiQ7ocW3nG1P/By5n/uqT5+0d1xXI96AOG6dYoYQVBed9SSPSV2pAFKbXa
zEPU7xju9ASZaCtVxPZ37xrbOdfmLSC+hHng/D4JfsA7rawrP6K5NOfee2FSy6mR
Yp4al5xNj3toUmqGMzc8lTt2yUTEZxeZCqPSAKbXszbv1N0x7cM4XlDUF7mecBJj
1fB8R5Q2k1uzjBqgqsQMp4a4SIfK9QDJHGO039rPkB7Y2yj2Wbg9SC2pldcrGQko
7R4FbGI+nPb819ykGXWsJq4/7yRWfYwTBwl0WFKbplxqWI6EkJqtY78B5q/1zq7I
HSmQxuuutQWMMWVI5xsxYzmylowOebWVeFmjpQ2Ko5f8txH9J6on1FHg+hfc7+9K
EYacGKpsrXas3s915RaTtDu6hq1GRXPHRnU6NVv/wt/VP7OPWOPFBPl7mQyfpp12
INtwfG3XNx+U1jLRbDAXdjAQ5mjvgq62BMn82DPvLROej/s96TihOdgQiv8uaDU7
wOMNJNKlbE7UOEruIdrVpF8EwV2eb/HkB9PuJ2qUMOGx+KYLAImgAgTbfVEhI8/t
SNGtsVQCjEQPP9YoEsThjJr4CcQlJ0V1yQQNRAvaPAhzdz3v9po8QIGbplFlfFRj
7Si04UC/VVLUiUS8NwthEo3JRWhWRDk+2Tw/WU8yMlUU9iIPsffstD/6K2t/cv+1
lEwxT5aijB1QyRR27rKlhG5eykeZmIOcDlQq/ndNvdikanD6D7s3fNHXwDIxW9uO
FAM+v1kuEg9/Oe07sXhQ7/oxFPm/HxI+pmHIXfytdPshgFhiaRSeqYr08uUg9Vgl
EoOo4XvdWcIe7DgbDicWL4yY6PXlEzKuAJTiHmYdZ64+oI2+HwKbdrNU2dxlt9qA
sBEimrqd+v8d73YxTvXetHqD7sNz3rl004/gh7rh36rAv9hD8t1aP2KMxgwYIeoS
JDH5QnUb64NAIV5XAgjpRmMpT4X/EEA17/pjMc7YDeP0Mdwk7MYzv9LLKi7v/I9p
ohjERCsOLs7eBE95bg6zp+KglbQNLl5zu5tRNJ2gFSXEqc/FB1e3eZaDnMq3vHfR
N/vqMwhXMmmbAzliV4GWBQoksny6XN74Y7hCOP0Ci1fIiTa61J+I0yGTntHpOHOZ
wdc9FiDtogeg1vLlBqLvVLwCU9ZulDbYVqKpjA5WgKWIJVnYyVdO0G+124STHf6y
j1CKUjEGaPx09UDrewJjzH5U0uVFJ6KI5P2r/JGQ7MOhxblozdRLAtxOrg4BDUqL
SGuSoXeBfyxkwEk63ahpXVrEfSkmt50CCw7WP0nSLs9wNdtyeELno/8QPHPhAI1e
mHollP4M1llVEcyGZBIZTyalxrP7pmy8KbnCxK5AZqi3YksVSGqPcB4SVYKV8jxk
Zv0Mi4UjwSpOMRfrsLMF4RncYPMPw1QdT/LYBYVM/+gXJgrYXPvfQ20DjylTEapK
1xpiGMbtYNcuU5dAy+Th416E3ljiXKkw4LVlgk5lMz2ouZECxTYqMUqMkdGMxjOD
RGh44r8iy0ZXeylZH2RFwhvSSPwgaQmM1xQKYBO33UhCrOuJcaJQN/zah+O/ZN43
958ByiLdkRLyQlI/wRPBaIelv8+/aUjWozqKKRkEoU9fPA64xKNr1qnejnJQmdUO
D+DQzWrJ+NLq27Ne0X1IN7d8B/G7zCm8MDQJT5XK2+jFo2xu0J51j48AbRRDEV6d
+kOu620DQNfTc56D54yNeVAVMkHtsnP/b1pABzIIxKx81cbWICIB4XtukxbKZs7l
OjqrszkYlLURirupseI5p3kw5AQnjRUZUijemEugcbfEjYLmHB1LQ/aQW/Xg8M67
46JtefFmySXcRnmYQXDwRxMios5jn4sfuybMBi1DdpjZaK4KdTuQN4B2wHLgBy2U
5yf+327az1FzxYPfsqNDaDbzqkxd/04GMX56G7Z3BfzTWBu8ssw/KfO0id/JDx7M
9gSU0dE/8DCYI81VDGHz9DL5xYfKounmlSY+XE1nK7Oup6yJfHrHQezA5fzV014j
SXz86usk+36Pen7nEw4pg/gz+nGuqthdfdKcy9XhXoEcdYtqkTH0nvMba8LGSCQ8
77U5boEWPLAVjq+OLj4KwRyJaXvRIlv+i3ifKkOcCH20nonvVJzzv/MJRAXvKNFS
CS8OBYedk1g0KH9dEjDUF5ztcPZ8HRXD+IIsy0VdePxykTwz/K/53y1oBBnGEjso
UTD3srFlZagStWbihlJvJr8tAc9fk88byNJsIRRauC2qypCTG+IVeBBgiFNLMHA2
iISLjOh/CmS1QI1aD0PVbfqd+xklaOX3+vy4q+zb3SZ/Y+8r1RJ4DM7wqNHQRJAK
4/JzOXOFxdJPFRiE/F7mbEbsolO2QBNuIXcd66UthcE5S9uLNIzQBs2b6eU5u6XI
PuCTznxLE2Ulu61cGz4n5z9KU8QLtHJV0cV/whEsFNTRmH874b8cRNdbCJ/jMt0r
P3omtqorbzvnWr7rBRHfdstNLTg3t1M+Onb1EcdLt7WX22NbUzboP2tKX1J6OGJ0
3MogadKwWWYBDh24IMpUEsm8j2WvJ6M2xR2oGHiq5h+ubZDnpzYAtsF3j/IvL3Xf
eSMtzHvwc1hDJyE6AxEPrNPViCMaGGI5xZTlJ2idnaYbIlEQLRW8xPpkvqdrqzLD
v58C4KH2tY8fjG1XIUL27PqgJ1f2OjlcJeDCJBYCEmDojpofyNP/1Uz35GIqMuVy
JjLaIn5xnxrP4yRTC1O0k0/ORdOMA56I+YjoiLJjHqdp5CR9PwxqQH62Iew2V9Un
eug6TS7244C9m04yU7IZV14Dh51uMK9y+GcNtRqke2XAQ58MkKnN0d83spQ3qJW+
TxBWehzlITLFBfa3L31hkQB+IXHhcbNzBHSNpkWToPL3PvFXOmtU2+gC7a5dXdLg
NON1BFRproH/yKRr4ag+UBuhT/ro7O6+4LS2APWA5t8JRXSgEBNzJXDJcjKwX799
jTGaJy2yniX+haifawLlwSzu7k3UVpEUaOqPgMFyx/SRGWa9UAEQnQGQsPoJrMoo
4jdMUhTdPm0904b5eWEMnVhUXbCeYv/7Y58qma9x06hWXZiJQ/uRYGn6k2LGWzY3
sIl6tzXIGNW8uBIEgfDgweUZLVOlp0Ov3shpAz+fz690pcaM6yerXFyoBA+Kb/bd
q+1wGx88f7E+46NH6OLkgOfaZRihqZO45RlCYRryb/vkdJcRp3eAgU7eEBjGFGJP
fVXIUurxFtxlg41kUAYZFiJw+jYUUBbXJ4VQw87xNFVRTYMtcp3fWiNnra1VjF/D
+b99mDdlhWtoi92+g7kFgc0rFOwFcsxGlJNeXx2JyDOn3PZNS8qcy2iXJJRa2ASx
djqeXYbM0Bkas+BChj9nd/e+AQsLkZQrYe5s6JrvQ4yWhvR8FLX/J2CZhZrC01GG
wX1PRoYxpZzzsI/VVoFdDewffyq5mqrn55DWT73+0k5rxVpzjcFmYXJcOzx5Y7K2
3+bSsBqlT2FRpLwI+865VJOmdLnmKc7Ko2D9x9KhDfXTj+hGFn1jMFYj0ucqLsc0
rDSG/GZRub3whAxYosLkgMlOx4zRCnqkR1D3vC23j1D37y+qlkWKeOAwdGR4Kp8j
m1cc1IoKDN0fNspIFE6IsPPu26f+G2UTCq7z/q4Z6mxL/I41cubRu3ivszQb9gnB
GypImOFh1DL1Sscjvg1OZRWE2O3R6i2hfHodqfXj2neeuQMgUyQBn8Mw/kfFs9NH
KsrXv5ogfVIojtB0UpFImFvCgDbWuZIZvijIrKYMrpohkHl4YCOVm3KsGKid/ZFB
Yf8pxMbRVIo64TYlPGEKHfhnOC7vqgYfezNBm40Tl2y8NObs8NkL6Pj9ky6Cxrwd
yRxGxKwnk3Hz7xepdhXE6RsEBQU4C6B6qWYenApBRAF/GFIrM6OMjeoPMtzto9db
rYfZD7Nc5RBD/qRyLWlo+E/LJn52BP7mb8hAZyMbjr7jyYg0dRaC2QB/lkq69PPL
0YGi2yvhvtud1F4cvwSZ/g2uKGKN4YhZiPjeUcyMPheAcI18nWsuYt1gNi9/8tMU
7SaI4OiNZDIyNa89YhT9nchNEUpw4TH+JVvgQyLgC2XAYWXhZDDS7R7lr9FQPJU6
H/KxUSg+mQ2Fc4HAtqNhzuPB142GvwF15fV3Wz7YtR4GkJAZtaRdgMaggBQO0Qgh
G29t9tOHhHHxbvInPhLq6Fgxhpty68Vb6CFSb40yJuhwT+np3RK5ChFxbEm+tfUg
vdSVrmBAAmp1t0XiBkzIMMKINj+OiIyYTe1Y3nyYo60QeIInSwN8XEiVNmpF3lGu
cuN725G7UIcahJq8kR6RAchzDZEKRKx/meU3ieV0bR7xp1lQdh/ky0tZAWtVYL+M
fV1x7zLIAk6f6IAlbj9IqwzkLizSuqT2Ti3+uS7wXzvFv+zboNgqx4FfYVZmygM3
6DMh/Ft9qwWvJ6wqdPOR+ZMWcFzp109eMQKuR7tuF8Q764GuYEdg+YeaxDdZB6PG
HfjPmOPcRBI+db/BW6bReJPd+cIVWsnX+ro/Vew53FLLEC8ZfrRGwux9BzP0UXgI
bXJ/K3Fnx2IebI8yTrBAUm0BFVRsFhAdUOu21HafWSjdzwCWEDm5Vcot1SMTrmUx
RHAxQh1mtRiQafL5ur/ePy9X9n6KeRuomD3/L7/ZKKjCldNzSkPDBPnU/Csi8TTM
o5p41FHTBVp711pFJDBxIsZ1z3nSJVQ5SdX2qsTDXnep2WaTyrwbq6RkkfozX+ir
ejwAhsVP9/tnlQJx2Bx6VPUSuABidPQ8NAOvF52TWvNMzcB1LELj/Ze48Wlh4VHc
skkzTw1XZ+EliixSKA8rExOAr0GWB8DC9MiSZn70Ed1nIn0k8xtXb/hs4QPQs8s6
+3L7IoVHb9ht3zRz0t1f3Pv84DALlWNLxU2YAaFCgDfSBBKFTxyxzCV38Av1p+lf
MZEIrgtOn98KnG0ZULtmavnY45O36+scaYSW0aeWUjo4FMbMjAUgAY06bN2y1mJN
F8DQYo46TOthogdScOtFquMYikSWWQgI+vA7hmcEw2A4D7ORL47ZR4J4nQ5Ea0FO
AHFRivoPcc6SDT6cCAYJZbjICdD5+P2/KA/LYuZ0qWHUI35YB4NXLHrX0joU1758
3hdGJ6/cMLu3L4XchOpepYdJxEPA2C8rF3Aba8S1N4elvZ0OdDH1VYNaN6wyTvPc
pMRbbzlZr9WKrRuEKwgPoSj4dDOeqIxZJMxqQ4LBbxSJo46xSPzKgqvTvY04ENDL
wzA6fPw+gNs640+WnyJyBFkfdkIhvFW4qHuLOFb0sPYzfKfoody4V5TuSzNqnviu
F4vPsHzxFLc04BxuQ6phDV9JhevXa+x4XV5jVHYDpd+F2SobpSol2nFQr4mXjUug
QeIeWDH71hfPzTFJAK619PX49HT5ul7GZn98T3u4VQGkH0M8U0Z9BLwJ2OAbXHLK
S2Nm6Y4Kx1YJHIgDIr6Ca7a4KHtwYlZP4OMIZ+ts7a6xfSYYxyMV8SxAVWIm7s8D
tqK02vce4SVbMeORxrw63qdxL6tRw7mSlXW9Wuy9TbNa7ZK0PR3IwU7ofNwUT7NT
f1O1ZMu3i7XNa7ij2jvWDoXlnQTBa4yf8+SwEgzdh6LBY7LjQjaMJCDckqwoa5hD
UnilWCLeYqsFRetFgtuOhVZca6fQMAE7YVKCGzquPUdYLXgPNe4oLCPxIlf5v1iD
QtSGvLQ5eKYW3US+Kskrq3bfo8aF7fBHDjXyzOuumAu/sWzzh+JExdTweS5M3bo4
oUR3Xsz++iCOcQSSClzLrWXqbgpc0DodXOPVGWXubhuTt+hsRFRyVc7ceelBFzCJ
ZigtBHBmUO02o9HFBHhMwmUY8Atwh4aFid7vS3gah2P1keCXv1Cvmoq4+i4Q7z8c
iHIrIz5lovli4gWWwZpAELySoGy2889zkPq8RRMltXQHoId073l0ynw/wp6K+bHn
TPrl7biY9Syln8qdHmY64SuCJTZJu+6y95C2z6WbXBzfMKUdLJSSncO+M4ztWEyE
Fasdjln0G5StzaaEO49+zpjzc7XDFK+02Zbp5gsi8XgpMogASnJxcUj833Y5Dfsb
51XKiK7lypE0L+FJrGIMicgidSVP2Er8MYJaSCnBu42wbR0liTGJ5JrF0UvjRWAD
jQPG5lI7Zebu1F5gqqpivAvYj/0hAfxANV4WUv50xeAiGlKD5wCkn9zyb01spLwa
E15K296j3ysWQ9ipFZ7c7t9OPgZP8h7RG+uUnJGbnPnz4WmDz4hGfObOAiWayS6A
Cdd1ZpdWoMti4/N+BEdiqx0Ubdvfwym2+I7FEBGxdGS8UYBLgkLJuROThcjgpg6J
g6c6A3BarQ6u8fkMWatKUEepSN5vn9m1ADow74cdrhREwdH2sj5wSe+HOilrhIG9
PgMjrd0EYUbQA6uh+n7ZsMzEfgg7kxmUW1uTU11YEMaBCnAe08EzFfF9Y2eqKXYp
a9SmKH5sWxEZ+/wYmtzj5u6XwLEPO4nH4Bi5EQlah86Y1JrB910bCgnAjyjLhjKA
mv3JWEalW48sC97IDNj9JYCKsQ5s0NMGVFmvlZguIW7/MtdLn2nbg8nYxGDWEbql
xXaXW19OtCYiUIuw58Vu3f4hJppcfMkx/KY2KyYfFxA8FkakJwXybOZ2ixvUkmpx
lRqfvb40ZhGSe7cmvSt2WRAQb1iT0gWrdIIJ2LHnvoaXCbdkwqycwEDkjVXU3kMR
kXITIluj2e+ETATGkQ5DP7T9BF3qOBVM1smJL1KAtT6VQIbX52YopNwy3R19qThp
+z2VBj8eHV5BEn88UMINelBJml1Ej1N3Vs1gGSyUY8WOmtktgt+1hK6EcNoD0b8i
OtIJ2kVFOSVY3tXLk9KPXho2n7dvTfbrRXhxlb7aJO3fx8iv+EOfU3TPLQ3hC0UI
uNoPkYImH/l3usz4Qm1Tk6f8f5RliMoNygAG2dl9/fnxe5XbNmBFKr3hoyUOiZC5
mIK++sJQJnzZzNNK8VAX4m/Lfz/Xauw1v4BKPRjAVKCxaRILE8Se/3WbaCP298fT
sDnUY/lpjrnWJDrx7KMQYYcMXNwR0ssrrWO9VTxoLDOecLsnCVn0Hs+o36stCABE
jGpWhDV/cXtSX6NsaUs9TstKgqw2JZFeroNghBhEYQxhX08xSLGnj5g1WLAiJe3m
we3PpzH8LlZb/fBjl5HZG6+/mBDc+Q13bwPMbUFrB6loJrvI8BZgXC6hevpc155v
5yeX2WKLh79/RrmuuIXUhiXdr07N/SwJbDYW/zZhv9Zhc2NJCkR3UQAToMr1Hxy4
T+JylMBFkjAoC5b5R9soqP+0qztzUJ9tOP/u6C28sCmpayJkfbEn0RnGPh2Gja3p
0hER9UsbjjH8Pn5Pk4+UTY6naIqPf77qjuADWua24cbPl23R/4NIqjBzfy38uf8M
2gSgeK4KtVqjMNFlStzqB9zwdXwHq5rxNUXD/L0Z7JXk50pnwuDeue7i5C0Jef9u
Eqml8SJN25+MLYTJ4jJVyIOb97JnQPudushdkHawgFejgn2afafxDTwA1Omn4N+E
viwvHGdoPMQKTqwz91+SuPFfGvIHgi0LsCbo9Z08lsP833GBycpkRCmAqn1mK4dd
nh8PfQ5Q9ZmatvPJanjPsKe6idbmEh4+eHjBWFCaecaacDaKpzjSWVTcsYI67bVa
koENrIu01F8cGfWeqLqooK4ZfRLJks0JJQbnk3XhNGXb5Kr8gaETFYShKbKbQbn2
K40bZCNJ9toKL8HUgOZ4/U7+SRKMB5raxKBmBBpdNmDnOmAnIDahR95YqPOg+CfP
Luh8fvZ9bJGvYFt/FqB5lM+ieBiy3XLvMCPhvL09jR6v01efE49aKxabgcaaNutb
rsYSFeZDE4dG7RPHYQwjZdbYd6M4h1cQD8HQq4lcRy8jQALwcuVkPC6+le61/rjx
qP1DjTuHn/ZHyglditEvr4x8tvBppR+Q2J1BdD1WgWnVZA+VoppuQCsQsqIazZgg
pbUVDB0qxaGLx6s8O4eFz+69hunFtjyZnETH7Y13FFjIlZ0pRsJu6VWtofTM/L2G
VaD6zJRrHgTo2aEZlmzyTr1g2lD0rAFa4yIwStlflFalpu+YZeBueXS2Fpnq8wy0
PkixV2DCE0vDX2IXFFx3eBYuiwJZ8MMH0zUEFE3/OEOHGDfM+/NG/uMqukPiNoTy
CVFXXsdL4XPn0PTqM2lwxOubksG3CUO4ltE+mqmtjUBHzJKOIk7wzMG9pye/Cv/Q
4crKLyHx7nMNEsIh+mElmknUdrV3iB+ipf+H8yZh53cVOkDJY78UwntvdnhslrqN
2564IiR8C2o1FZJqq4/yXMqehDXu2hreikpSqSRbUACmPnCRF298Lw6j4XoYGx4a
C8lfjl8twpGBj8Y6dD77zGgnK5j0jjKgunso4MEWyVTEpeiYre6lBKIXk9d90o0/
Uw0n0JhCUn0dilEi+u4029tCaDprywy4JZ+FS4d//dWAMF/8MuT//r4DgI9deQHh
LC28izRmFtTWbWUwelboBmay3kpy2X1PyaeRPjD+/YQTqp6qYqcR62g1c+flVzPZ
+yMAyiikL8WdxEEdFmW6049q7IzC5zQdPqav3Oq1UewCpVPfD399mvx6KSTmnWP2
wmTmOo+Iey9qVY3GHHOwr1a5x+Agle9cOg6dUW3qtiakhJq+T6sX+mBQNxkVvZ2x
vozP7cdYCTjVKL6wfr3JJ6xUUhNQCOnWEkkTSVFRvPgv9vYGzMs7zqvov/bqhXtJ
oyfkqIiWdvGBGZIA2UAc67/7tLtGPR3L3pcq6ljpJLafnNUMz2WO1DXih4lrWKPL
4L139mnIQchoNccgiYW4TKrQ0FspngwZzW9X0nyYHRHDJ0AnftCVOGnlio1WpJxZ
3YDd3RNUKBvremhMWWp44ZFbkHJsaqeVJ6Sv++RQzpwEKyXi7ERQg3TavX6eg9jX
3dcqVHGK4rhHa/TND/poPhzIKDYHWtrsQgTETUCGcmrZ1Yu1cGDokeln7PjKTR4h
GMjyQ3OuZDdo5Xs6uAAzKrI2EYtb8CxudSqyM6uU5PBO3Qyh427J4hP9k+fIP7yC
dzt2kNxXBc5kuXHEGt7hiACk2/HoBCQ37mPKGQVgVnQYTb9zlYyGu+eTKM2E3mA0
vIrzGXAWZ+oJDYiWPXEcyr7fc9r23hiwWPN3vaWjFIfNV3V6P8/RZMpbyxj6c6rV
OfAvqLQYHaLblUCP57xkHg4yReqRf0FMrMIarHRSZPywAnkSDKpIx+5NlbiKxF9Z
xgxP0Rf/SWvyNyB9rTpqs7W+MRrThyUHnof8HG4xllFZaVetp/fNIssCUxTd5Lsq
5RcgYIJLs2MIfAByrhO8yLAE900e53xnFHDEDwvdNLlxK8G9dWzDr1iyg6aPnI46
M/+wDkwcd3qOZ7p9tyrtQFGPnKqrHPNOb6tBTw7iy+VijGm3AcES1qwi5yw3zeZy
GQaxJrQeczRmSBNnJKithqVF4KWwHwixQH4x3BUOEjKsw+1LmIJRrABjSC1H/gLU
HZShdD/zjShBlE7hCjIOCC1mkV1qxvoYYnz6d3eS78NuBpF4SZoDYLcR/GzdrynU
U/pWGihBKLsvM6/iqpIHkpi6bjMVVXNGbEbh8RZhMlxB2oimG0ZqMwF8nspk3vpS
qAvGhJn8l1zG3Dr+ihin8GaVDJ86yh43UTRvpoXTvOSKHI61q+zYSI2a9SPWusjW
90Jh8k0JsU2gF+T1fwCdO3DjAN84R0NfqNIoUUtApCFOGTiq26jUPcVbT0WTt7Pu
9T3Qdm1xPqCVrGSaX8865BNMSpjhibHkWjl3AjKNp7g6vMM6nnRlgc+x7B9P2L8R
AgWHm3VoGQ+YUX1zxenuZxOY+f/8qun4sB0n+K4cyCln3d+UaTrX5v+a9jWTuWCO
BfwJg8+PKXIHKBtki2CkX4S2471xUxY/wR82hXKTaQCXuftIH6O/A2QIHPJS2LY+
f39HIeKS+nH81FiCMdOzE5n6GgU8O0IgQ2GnCScHVlONbgtCyqr2KT2w6BqtdB8O
1QFNus2FB0+NmkQG1uaDN8UOxNCmmrI82GHo5b5iclGImxUgwnrIcBzhLpb/NRMd
CNgFe3s2hf0FM4aDQxINeCKgkMqup5MBYkZIUPenFUcanoRnEv75EGrSxCe0SBiJ
5jRuSu4oh52uS0V/93DxHYzvJLspd9si9egDDL75ivbNq3t7gaX92j5IlpiEhn4l
mygIEZGXN2hPJ/DO1mruNM2HvPiXeZcASIfML7TVqmcnkUjcu3Xbl7IcIJscTK7d
C0cgNdtpSNlPX1QFXCrk+ynnYld/gWGqDW6OmCnfUgIoxvRN3rzBLLPKEXk8RJ4w
t126VMQDQbqk2HehUrtCcpX/lQYCh+zSP0ovsq1CCainvVLjFTx+la1ciJ6FVGNK
XB1gw0VqNmqLVS9kFF6ywzAY7xaRXhVPje+8YHCLINisK3VXG08FXX04sagbYhDc
i1jTQvOl/Gpgi1wHyMayC2w9fmVcJsN1a4LHxGk6NrzEEpuat3IXqzIpJeRV86M2
0hFDaSyRu4UoiCOY6R+lTKkmk4rK4hap17dvERrZv+w9BTV5JCFS9CIIGsE/0XKk
5PqcLIROv+hiHs2f08ZJbU/8WJCENQM/xhoZw0rRTly9aqj2Jh7Mrc0NUwQJMRUV
SOtYg069DWOX2Opi9TviOLPDLr6UtOyeLzrB/YIWku/aRSkWT+YZKa55LX3NuBLk
+cVPH45cxHA7URjH18ANZ0MchHsaoVeCYScdg3USX5XMyTb3AKDnu/x0P5RPPqov
U4Qil4yjoLgE12VYIYp+2pB0/uckPG2043jSyKeyr0B9Wnw1X6NO4X3KR6rX04G2
zAD8zjNV09aYggQw4upKyR76n/6ltffYTE/YNh3xxcNT+gPhptcuWH2S4QNg+w3s
2jU0YD4+em66xQOw0EXCxkJRxMscpdAirTmU/1LnzWdd77tD4IRNsc/JuuzhkpHF
KE1D3aBVy3mu8M4Tp7EMe/xevg/k5FU7fKO0k18LNS8Htg1+LYPrw5/luwl0scQh
gENLnyyUnis1YoM15TTdvYViw0KV8yMm7uYCstje+kyafDDc3Qq1Tv+UlDFtRPMt
CpU7MQRolVvdtimaphPYsUiUamXY1U7pZwQzAJ1XfqlpwykBR5DsP6OyJK42+IcV
oPTnnwdSBVRfmEJ5UH+lj36nMOPkPR311OXtO7oNEwxudKUrIaQHRpV671h1plQ6
gkSUwA53SZ+yw6VVJf50m8NswTf8DlubFYlBMsWUnyFu9GCXwGkKYIUj8PkibUtH
+dKvnackQCBdvzT//n5ndKm2a6eEp2CCB0u0GtRoLgGA9SUIzUc27UZurKCgYCci
ibz6GmP0dpoJ7UbRs45zcq57dKAb0AxxCLS8OGG3MDoZnyMyu4fiGUzKGq1o4TgT
ZhlmqCgPhDcLymSo0Roc0QwKBBexS9gWADAcoiDbeJ0aPLOdC2DptqjtkT5cm7b5
kxVVKncdQR9ykVoTLVOi2XHSWfJqDm7VFq1FtEgwTPVWNNo60xUtuO/m2qJElEzL
S2VgFF34dmuwdM6y2Vgi3TpeUR6D01XPjBRsMogRwYc9C6NH6dBiSjwrPn6nMaFE
4adSoAfy42U32384Wl7yZOrDBL1yRkIC0mRHPXPUwM7QcghvtcUTcZk4BgEie+JZ
m6OqrwY9GANetWpINaed6jOvgienlRNOOxCrUozT2QBdA4ayHZ5IGA+CE4x9rVcv
XGlw1xWeaK8EkoKqJ++KDFKowWEW3iZDVS50lLf6ynteEycSBv3okIXWeAEtBaX/
gV4bTPNZWabJ8Wp+daM5RwEDzd436154MeIeVyIjSDIt4yIM7Fo8rIEZvYZNH7BJ
F4T11gqMUCL0c8SHTnmzPzZl4C1683bQ+EUziZvTk92KpOOSPoTxO1rr+bokzaac
wje2ZCcUVcvYb9DWyXNJWUM3gEIe9LlhjZuo6RnlBl5DdMuuz4EYQEDzdypUbCH0
zsmJdTGh+3Of/5qRInDvvmzpq6hNugfnoHHU4+vFMJKtOBCtt95mK32ezGNLOR9a
9X8OSem9T6mAKsoz4+mhvQsYxliXPiid4Ms54UQ4XIeH0/LuGBEqXW/IlGRXxugT
2Y8vDjnhheo7uvY7Sy7FsBxmmBlQdF5FcM4x7RfmRRR56GBmjY4UT4OH5yy3RSgG
wyt+CnJHNU89NgQuZIYhZYkKzEaBZkwBmTAcX9/AoJ6Mg87h/9ZY717E52JbHi/d
N7P0hXgJrE8dhdhX8Yc4Nv8zeuZG1xGeBY/xn8hQReFiyVst1sHvW7HbnkZUflsI
xnc7Cn7NuZdFGZqtz16t0GXJl41i2QMhIRDPwHXF2A6Oc9rwZ9f2pxXHCiCWH5iw
87hmgoAazu/1iTVAnSy40qevkuCC+SPKv4P3lCMemwe9EE1bQslTBESoXjmHiL1d
aQPxahMhpfBysYtFKGvEs5X8ARnPn80JbjaS1/7xUKfoX3WxYPT7O/zsVrtnogf5
IYUNagMLRwEr6EkozCGuhhfsKa7ONtVMLf7DUBCioPST4VTy9T+Gt9xdonn/wIkY
fm+16w9byucU2nObefQM+WAAQDCokaAfYtixHx4I+C9ZEC5EfN48GHFaB1qFCWU3
5d0lT7Y+vVBCRxOl7Q/IsfNv1bITTp3xRcJiERSnftYGSibwMeDSsd+xOSFgkmui
TRkaiETq5t9AxrKVUhkTZG0i7rGi9wjgSvCZCQ+mfyMwH6ELfvk4PM6nYGiP7nrI
/IGCLXt56hwpmtN9rIATXqCHz9iBxjk/px2MamWx5/EgF9qqQea82egOVQAk5Tpc
ZPmEd4Qln5C/Dtk2JQTKO2luipX491VQ7ZLSymI824AmqmtAsx1MiS9EdYxcy75f
gCoBRD2wre/ybvVT4AQmT4PPyBpif4DfybUovt7ITEksFY8kgAGaadeny9B6Hj31
OK/JdsgZhHAtro2cn+haY/yX7qNmTFK0+vv/6KvTfqaNakvyJrCp41+odBASxJMN
/IjLZySy2LAbkwITn+RHQTsdEvv4r6SFS7K6WnWhZ20cAesOgzcXH8AmeicmWgZI
2oC/7C3dQyWrVy/NJQkGZjKZHIbphC0ISU98XwY4W8E138jIwlgk4Fv+tsU2TcBD
YblJcui5tVh5Yv5SXoLwS8lsXrYN3cZKSXtbVuzE9ci4UFhT3OL9O+wa1xuw6ZQp
h+WnYQRBl3nC92zUPCe7xDe3Ee0SO9Y4anSPWKirNIouzBNls7Jp5rdJ8HbhPbR9
+xIV6EguP+YXIm8ixEHfo9gzKF20f9Rc0VRBnqZxirzGB9VofeV1kV+xK+tTm0+c
`pragma protect end_protected

`endif
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
liuVcxlVN3l+nAhVJCsNhe+lo3Vf8z68FnpcQH0pd/fuarSq9rZxcXUE/cE5emzi
sjYe7X7ywiUdeQspNW5ifC7ma8NeQeruNux5OmHkCOly2iL+2bvWm2nfhMrlPikU
uPotuXgietLAXRl7Xtny4jRh33Q1AilJtXleY1mcTcI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 64722     )
wHTUnJGFGr8slwpfq3jfOJDJLDkcCMmaHMeHmGKkoZwTwQbyLmHfrJMqRd33OCr4
4IwspKTPiBWSTfP1Ue05WPbSisniEsRQS9cz99fACrYxtudadDkYNpJsEq0mpuIG
`pragma protect end_protected
