// =============================================================================
/**
 * Class containing the events for scenario observed in svt_chi_transactions.
 */
`ifndef GUARD_SVT_CHI_SCENARIO_COVERAGE_DATABASE_SV
`define GUARD_SVT_CHI_SCENARIO_COVERAGE_DATABASE_SV

class svt_chi_scenario_coverage_database;

  /** CHI Node Configuration object */
  svt_chi_node_configuration  cfg;

  /** Array of pattern sequences that we wish to match against covered transactions*/
  svt_pattern_sequence  cov_scenario_seq[int];

  /** CHI transaction scenario coverage */
  svt_chi_transaction  xact = null;

  /**
   * When a cov_seq_match is triggered as part of a match, this variable contains
   * a list of the objects (i.e., strongly typed) matching the
   * pattern sequence.
   */
`ifdef SVT_VMM_TECHNOLOGY
  svt_data_queue_iter  cov_seq_iter[int];
`else
  svt_sequence_item_base_queue_iter  cov_seq_iter[int];
`endif

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
JXbC5MsMJJQwKp4Hd+0zL9ymcN8+f60QWynJtTXn+p6zBRL14MhszALcJUjI/nVc
3JRPC0yS8qaFFpPTiCzMHYOFrdaJvDVFZJQoUhFYffHIdw49rIRkPQPP9EUTT2f2
ji2oqlfDjoC3VlKJVOZHERsqfnggdKnqSWjcZl0wj0+irbeYtFUHdw==
//pragma protect end_key_block
//pragma protect digest_block
U2jf6fr2Exxxsg+GoGek5hajBNU=
//pragma protect end_digest_block
//pragma protect data_block
Lf0Vfy/3q4HdcCj0abz6i2r/H9fNN4Ik3JfiGtvHr1kiThBhJ594FXWyDWG/qZPX
U9FQhGp0MKnybSAFRZUAXnlLoP0lh+EOX5wr6F7s5RnXxdYxBKZriKVR8qDubYXl
IEXKGh/YJfr/UOc0NV5zwNPRoaTGwuJEAozTQ4yUgATUytLe9eJqVp/zaU0yQp5i
f4sFe4HQVHiFx2ejNK3X/XnwlIpENWERlkJYHkU/0eTeUlj8HNlAtI4nuCp6G+Mx
pHnGFRqvTdETzVI9D83cXrTtIeiKxY3lc1g8y/BhALuTcD3vmLZWR8SFXZZy2qC/
TfixTxhkzp1ODOQddTCaEsOPzqItEIS0A+vxApcneZ1U5jyaWNJTQUofHE36F5EI
/n7gFOUk5pUFWWp95Oe/6ESjwm83x6aLZXmA+4l9SN4yTHgmqYyz0cQHZLEJdEgT
MixjzIF4ajiWKm91qCae9pss9onYIwe3Oi1Y0Pdw5apLdCOsHI0cO+K+LDA6/HKx
aGx29FLMMEELA5no7w0u6N9edWwFzTV1H8EEB3LPdsIdPLmdtm03UmI3qGtzfmAj
/7OtTahrV0OJhPKZ6wDT3g==
//pragma protect end_data_block
//pragma protect digest_block
pAkkSqLmjFxCCnG9GHexwsn+NQs=
//pragma protect end_digest_block
//pragma protect end_protected

  /**
   * Table 2-9:: Order between Transactions
   * Applicable for only CHI Issue B Specificaiton
   */
  int  order_between_transaction_sequence = -1;

  /**
   * 4.2.3 Write transactions:: CopyBack Transactions
   */
  int  copyback_transaction_sequence = -1;

  /**
   * Retry/Cancel Transaction Sequence
   */
  int  retry_or_cancel_transaction_sequence = -1;

  /**
   * DVM Operation Transaction Sequence
   */
  int  dvm_operation_transaction_sequence = -1;

  /**
   * Exclusive Accesses Transaction Sequence
   */
  int  exclusive_accesses_pair_transaction_sequence = -1;


  // ****************************************************************************
  // Sampling Events
  // ****************************************************************************
  event  order_between_transaction_event;
  event  copyback_transaction_event;
  event  retry_or_cancel_transaction_event;
  event  dvm_operation_transaction_event;
  event  exclusive_accesses_transaction_event;

  `ifdef SVT_CHI_ISSUE_E_ENABLE
    event  memory_tagging_transaction_event;
  `endif


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new svt_chi_scenario_coverage_database instance.
   * @param cfg CHI Node Configuration handle.
  */
  extern function new(svt_chi_node_configuration cfg);

  //----------------------------------------------------------------------------
  /**
   * Method to kick off the dynamic pattern match processes. This forks off one
   * process for each pattern sequence in cov_scenario_seq. This function forks off processes
   * which will stay alive until halted by a the component which initiated the call to
   * this method.
   *
   */
  extern virtual function void activate_dynamic_pattern_match();

  extern virtual function void cover_xact(svt_chi_transaction xact);



endclass

// =============================================================================

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
OUvqEJ66Q3ud2fag7WhvVCtZoyVgvN9AIFDBUP7ySZxSNPvfEKiLhu3Ory/gp7Zn
tbc9dwjG/sIIs9oaFcJjVlNz61eSfE4CpIMLjH7gG9+6umIQjyz+VjAa9XRakAsF
IjirtwtOFEynZBDBHhoCmt7mO1y2lnntoGUnh8QH/ZtPAfe5bP/AWQ==
//pragma protect end_key_block
//pragma protect digest_block
ROzxArctHPgWdh6DXcqK3jLFdLo=
//pragma protect end_digest_block
//pragma protect data_block
tY2RIk1nH8MRW/qwVgBAc6v4jIy1/Wlm2HTWn31FW6OMIR68NVlqaRRvaXo7qUoY
g+j3rrrGnz9kPAAvv24gWxoo96GtIgMS6c0h9nfnWN2gdas1nuJSqCyN6fdMpAZc
DWOlrOI6AM+w6f5UMFTvQ8+L+rtG9ImKg5I8CY9uMQXM5aziINBSlTkXcDqFlckq
qZ7kYkh0bqRkaSGzFM7SNaMpyhmd0eLt27umcV4vd9jrBpWYwAgr9z89JQy6sY2U
0AIxaVgBraHlF9nAPsbt2Bgfa92rWpkhlLdKaJY+vo2W5NPIMXpBK+3BjDWydVmg
EkhpeC3hFR+ei02SkYiwKnwXiYO7fCEJRzMolQgb+jr/Rc9TP2r9VvAl/HAoyy5a
oRyWSajEB6F/TyPHXeJwY5JPBK5mtPKKVozqtkW3dagf8UaWa0VQc/5Y+uL406ut
kMwN4QRsuh+wD3Rz6a/8Jb2O0fOAc3N1xYhwacyT7CU4VeucXvLY30RL2q9nvAiS
StTXwhvQZhVPi9/cAG89i0CBEKwuGB86EMuR5c9lmg6ypAyU13b5RqN5E6RVlOvK
AyUxX5UXh9cXGgGW1f0pGzqvURtXqv944Dtlla/2+2KFoaxxB88NXFznf+0hI9O/
DVDtxV/+nQGllpO7wmqLTdQJXXiEL2tmyMIKPvRu6d9FSixm0w47H2wzElEM5Gc9
BbM9GsP4L5RpuBCxO3KY7xtnwwyPRHIUoP2yaDWHq1EztB8CSMLoHTCP60WBq3Ov
ha3DFnF4qRRKE60Yh0f79i6e4/FzvUDLt6B0txFzyW+u81KW+aYED3Ip8fvN1Lqd
HjMY24p0t89XS9tF2udFbfmBVi2aIZpWgQpIg8nbs7t7mh9jXB2DIGXy5YX3udtu
jaqz3oBZMONcWkIQdQhax1bIJj8hdtEwCduvicwnxS2m6R/dw1iQtS3idysD0TVX
QXR4r+MbGtHjLufQl4SG/jHvqmphWkwze4NTyLZLBJTlcwCHzQ6QIUJbkE7NGQPK
NIpaQU6oLgCsytAw8she03wyBA0DrkCOuUpuF+tnIC9OX2Ss6C85XbHp0GsLu9JM
2Y5cp20iCCUPqRXgoz2SDB6UpAfXjfhQqxkpBnjqF66UOLgxvOun8HlDpDgv1AwU
CPwOTGMgi2YxCGYn2FPh17i4mACHwXb/SRAqwD67BpuFnNWUJBgLWTrUJsUw+3Ae
xds8TgngJR+0ZyE4ow9mcX1I6P8RYKtVzjB6+IUoc+ihM7YHI2/stFCwDVv7D0X7
Zwb9IZ0Tko7jOaB08+Pj4pkwkXjq4x2HLOFOxwdcWdXcVnKINE93bJbzBRj022XR
YW7Tbl87lvNwjQiduu4b8UMC0A3YOQGWvsQ+YHHMHu6EfmNHb1W2dKDumDsXcXA1
CqvKHCv+cLxIfH0lJoxht4WdfyE3OUUHzy+3+jnfAz2sDUzFkyCRjzLzzX6s1sPQ
PYmT43oLvrWPnka55I9LaGDBofllLRmXSjQh3gFGR2oShBnnGlaZcYruVsOyASoU
i/MWJ189WZIYJrXIvhYUvwK8laQF9PqiaR0JHzWGLUDs0gTIwV+pE2m4YGI2jHbY
x6Wep8yUWzJlqoRpuA++YNwv4xsunF0DjQMGBov0GrNiS9pUPfNcU4KA/XcrvhTg
8WzhYaqodyMg1wUlTaDuDQkhy4+3MkqVikBOOlZZh9Q8JHdtXM3ZtUvcwMvAik1m
Mjlg/wVcZ8el5Ynx35GYYxC4libBx+v5QNYPSkcyhY3P0/yVdpzFiWUYJc+PS3GF
Ps2PjvV+bkde3/nf7AjvC9WV4N+DNseZBNsqhJYGhfz8q9WrIb6nHavHKwh0uCOg
cxCgCYceyLvPrl+yoAzXZkg3oHqj+8YuCf+0juF7m0soaj1tt6h54ek9LPcmwPfs
2TWB6JibJf6LDQSUHmUjxUy9p0vPoF7fSIHPhP+HntNTSSjdtXm52qZjZvOVTiGM
jj297LwwqpKR0Ud5QPkmJE9clLfNxunzKp06+t4gvvvgx4xxkzSOPu7oFbE97yRg
lbUcqt9YZRoZfeHz5T7mojZTnG8uX2CwPN4CY0ckjUsEFc0hPQ8JAHjpLpv11DBR
TNOobXp0pDLWHahBwC+O8qS9rXaeC/jWCFiLCRTSyQuTTP44gM/kKK+49l84kW30
YvupiwgnY9wdGWWGHTT7FcxVxj/N75/s+bWorXM0lutsc1vjQDGNsJnP9oob8Q8n
/aOZk9DsUZ+7Wjx8VNzR+JYurAcyq9MaL24JZ1X3CQlIkwlNhVIIqBrznczfZucm
lCgDIvj77Md7b1oG2esjHvOCUtEhhQE66WuqA8zLMNeZ1cq8hHciguwwCdop28BZ
fr30qRfzz9HCNPRWkgfB0I2tVj1pilWSgjA+POk+JSUnnGqRr5UiSQRhWVC/G8CQ
6fLQ9cS01calQCz5cWA2kWzNqRvz6qtbizx8T6P3fWZ46uQVIR6Zk1D8YmhUij98
d2CkyRopRXECHfze3VS2k22/bhHQnukcDFsMsetqVSW4CqJ89bjwHwsrb8z5uj5y
nygGX9tSgMkHyznKWk1/FBpnBbCNW0gWLymnVe8V21OJ6j/kgwZ1b2BM5VYJ4PUe
SVduI2AuHWLHZKq42OqQ5HZOzpwazh7SqJrQQiN8Z/qc8ggdA9Cik+eG2DfVoXXz
5s1bi5+9y9pQTXR0jWgxpJPYnjQuEUbleC0irgoN2vUysBnZ0N8HMlT6H4a28Cw8
IV/YYZhTny2hod905skpBM2AsxkEom95uL01BvhvdMDuJ4FbJcl2gOKE6RhyG9iB
LJ8Ju0BgPBn2CAaj3lTgbh5ty8I0BX1+XaN6ScV7/ltcWwHKxdM8viDMfP+xIZLU
jWDJ05tmHWuC65dTfV7WnQbWgU5kK1fSNTKnaCZbJpUZQBDrHyPG1AsTtf+IUDx8
DaHpArE63/swSosFDNuIZa0noR0jVEd8zUci6Ijon51arQG4SSyA3RE9qRy4ZrQp
mQ3CyTiUIU/QMcHs6lf6mnGlHOFmYQPTDuXkGQKicoYd+AHo2LskExily5sqim/F
o7vMeCVXPlxFi5AEsiFIjxi0mrsLmy1LjThrUWY59tasx2cOHzmzmB5jZ4ZlgOov
U6RjJ2HPHw2Oqq6+K3D/EY1flGYv8CMsI7yOx4IGqPzxYiyRXC5jS6GYczcA2th7
j+hso1MVqhrUFfjrNApc5+DWs87V247gygcq0WOKRjEnv4Yqb6Ssoiz1nWluLDgB
LAKJe9SIXas9OMVrrl72iGqJfq//dNDtGMM/mljAFqF2kLtbqkxFT8X+0GO+Hms4
CvaGZycjvZwwuRYYIRTXZjqcoEUiMVgd0nIN2u8B/h+r5y44D047E0zY9c1pMZNJ
QlxO4G8J/Z2L3vslJCEDyK+789512knbYR4sUlsUkahsMlwgu44MOasrNjS+rXOz
1Bh4OaELAjehCTM7yNI5neEH5rtqQXa1bzG+m/sJmD8SybnY2jbHALeuDTyMz3Y/
TZLg+kCPnvtPQeLj2wBTpq+GhMkDCtSpI1QnpFclMPE7egzp55QtaoTAla8ZyOa8
ZiIPMqnFJzlxlWM0f46DAPhM82DWvX3UNs2X+ePrHEbgaR2cbYBY6EEbrdvPRWnC
P1OIHX5DzuRYyscj7Qc8TV+xIbtfbAb2t3zwsh+H96fsGWLRgHVdNTwD9bNmYHPH
QfJiAvTWOxUr1Ociwu/t+ZeINyMVXPrVVzVSoRX1eXEmREczhyproaMNivYBaSxC
6r+eYze1iSgEymByT8oe8k2uRQuXx4V7VzhwXNFtvGwGrHVkGwI5CrtajcpZSLK9
r6LZ5CjtK/1nrEuvm1H6GBK3m2SRJ8YefZY7r6nA4LSXrZV5cVv4aAWhUHgW6zz2
ROrtgjOOIXwK0tIRj6Jt/Ph68y7jfW+uVpDnt0FsXBody5VYEb9y6N85/akbMwzb
G24C619/LT2GituwjpeHpIOOvzdd0qwWkRJaJSs69XwPh2ePskcqktRaOLlgBvWQ
86vbvF1TZmC2tA/31o8JUSfvewRHN4rBi2fGrshf50ORNTx9x4gYZWuqRx6XQfMy
FveH13FR2MXAiOhTc1ilNmaBSbVezttCJ5hN6Tyii8bfzqOrdg5s1+UBzP0jeAgg
Hq8Wja2KpMgGVGQWcmqOx/JakWCfCLwVqhFI93mEFZUY/2KPRSrvw0yDKDoCY6VH
9ZwJmEyUx4vJ4RDj6oJ5+q2u7zjmJ82yTcvBk5ZBGHyPYRM5KdnZaStoAzIT7tNx
xQXGQpXV5yqN2XjKhMwFNQDrHE2xWiwbzCgblXQzDR8yYfcYx4oOo4jsPZgac15K
edJ3ZHISB4Buo3GC9DX/+Jb+GeM2g6/iPk09cAQgWfCy9QPjSdetV9NFWrxNfN58
g/aSaXvuviBRHliUqAd3fgiH7wqlusgg7/v955UQAJxhZ4wvqiRPAQQsCF1g49cR
rexs2twWgo0+jN8fU2guqU8vhkTfJO/ZYR2ez5CxGhqpbFy2SFfmyd/TiClHpzQH
3rgvne5l1+xU1YXGSVrNAaZwv89QLQPEAexGQJVcaVV11trq+4LJZKBIU+wRNx2f
C8YCb0/+Nz7nHJiyo0LTc6hl9cRKKFwzp3jC9IzV6yBZzcM2LYVgVFRWRQddhY0e
lMsiNK/SEeaLV7XgSdyngZ5e3WrX+S8J0uj5HibjIVdSMZSAciGWkSHD3e/5trGv
pUrsk4xwSwLXI95PNrK73sWzMK/PQ5bOhnEAeGhfMj3uTOXRNOydpNU+OLPcNCmM
jJXMxO79g0prb/PHZB9BbZg7CyVLmicCm3/LNg/FPWTuNtfJ6i+3wLWVvlCNHlrJ
Z7evFbmc1ZTac0rCVLm6rVylYbHvSysELqSUfi7zhdsrWS+kTVYnI6fbDN8NxuiW
UjHd+90oBVWCtbjZZK3WnnfSi47YLxRJ4/djV7Lgxljic3+8BTpDfiUA3+NN3vim
xE2EKOJN5bY8H7vxqdxNJaAatmvKu621mBnB3QW7U9d0tjpbGwMIgiMyrc812u5z
KybGJGJxNm6I9FsduIXKBd4j+o2sClxJe22OzEIfBsb0YQheHxWKMGlLHKrfFZ6n
iDlsFm4T0nDoaExtSAc13y5iUDXZjcEx3f6vU09R9ne1gceEPEAvmbcIFvAEuEOK
3qOie/nSueSXh3rZl22Roy3r10dbQiao56NUiMLbPHiOBkhoa+PLi+OXxpm834tL
7bBbLfxAkLENqXm7F7XQLEuRN1Dmdp6dooNzQ5yodJTVEfFthFZsNS5XPekHi9v5
hb9Vg2ZiHw9YYCLgeJ8x/nvEzsD6bUCi1ySeXHN2Y8LzXvZ0Bh20enggyS3WeplF
FzSn9TYSSJxWLND2HQTauM9+b0rcnbpbPKRY0rG/r8tPPHetZOPqw7oMyCEvOmrh
00FRBIJ11ZnyHsTYo3zcFxjA+u7w5TMOk+vtONzlCu6V/ViFLHdLm34UNrNgMUJn
EDXiOvubrfLg7grkwzwO/8IOR1b+0IhhmNc/ySYVDWWU8SUGPO88OH9+8IQoJC53
Su4S9BunJlj9IUtCU7eV2RahI6efJ+8tyE6cJ80HSC9kfVo0aUSjunAa3/SmAxo9
GeC/JLvrU8xnzNWNSLk2PrpuDCJWvqtqqOHdQDnl6QuiN/gxmqqu/rZejzVNqas7
6c5sjzTh2jMwCalBlYqZXZH2ZBmmdkaQ/O0HzrjLQ4zckKR4c/Ccz7zcJ1negctX
MI6p/41IwqtSqcCxaeIpfylL4YE9kYvnGoywCagbWPWZFMS3dtSeq8ZAUGoigP8X
HadMh0PJtxRixL5E+TbkRZN44kfhHe4EwskaryDHCwpBqNdVeMcyeyN3q5ssk3OY
D7MrkQWKy3+3Pc+4jaXfFT6iijycYVbT9MOWnL5AhjQqoIKXaTIK5nL0YCAl687A
hnutw8hC61BZJ3Fu6oXIHZsB5mcJwIXHCyYoMllhIsOk/32a4+Nd32czuQlW/ixM
IUkG1XNWficQE1b8Y6FRNXhMMOA3gHDMvr+SraC4JgrCH44VQN2D+4PwHcXuu5fL
dExUdZhj3DZUaU8Wu8zQRYrDS6NSS7f5UnDOikmO5Zctg0X3jUXUe9P+cYbxyoKx
4Ff6LbFCcue1h8NeBCuvUCL/xHPgnmW3u6YTcAiHoSwx3k9AhQ90P06A0Lg719du
tnFmmWaIOGw10mnkryGO70ERGxSV559k2S4ZoYCN33Mr41aqTUt1XGWujKw8Y+l3
fELIAJjBI3kRUbF8MGsy5qYCD6pQiJNiO2mBIU607C721ktYK+46dNZAuBmQhTu8
GfkT+d+4Q92dKMA8oCKda6ypoH3JPShFKyhK4p8bIDZQRS+SGCNlnxu1xgsaD3RJ
a8OeXQ/F2nmIpzJnKaeWwuMDrWDwr4PgAV8JkPr8v8+ypRt+ubbDlF/xRneZl4nj
UVo6QZg06W2Rs/Q4PB4UOovezy1f33tT9Iudw+webz6QVl+0CshJluBXMbVZwJWI
fDTl0naY4SLOJ0KTnafHCxw2u5V6AYEMqlxx74jV7Z5ydNVrH7MaTCq3kA4Q3PYm
u+y/MbboHWI0QxjRWXENq+A6/M1pzhfVETU7g5Yfs8diWAABed3PgvGwCeaP1+cm
xMOcqJiMKSMpWQp0B2qp6m9TA1daWORpGVGCFq+R5urbSUEbbTMlHx4z9FI0IlMr
ugGyd0QIng3JLFlkttq1KA8TtnNo/z3H0wenPqzyCfnmG50wZ4XRcdx0ni58mgeu
GLCsLsHvuNJHqncY33xS62r/RbNEhoS+gOkQy787bZCbFso++lZzPkeLrvothEXS
67bG9XOjj5cRL9+bgBQIuNT5tYbwc+AhTBBARFz90Orz65BKJwpwPjwGEvSIL+v6
TeHzL5YWtqqNYiO3zluq7Rk/OjTb2uTLHKlP0k+fDULo8pnNSn/1W1187EmdVZkd
55TzHVkqAua0dLzzUUfzIKyCS3kB0c656L6lroTGRxx9yA61zcMjt9jO1vlmrGRE
d3IconGz9YrFD1dd1GvS8Zz448ZYRB4BSW6I6Siw9Q1wgZ7021KxKKsD5lwV0xlv
I7c98OhSAA8d7aHxWPQRS3IthD4NdiA8haHU8ksUvUNWPvWiTC7ouszg3FeVefYh
Y1jnPkghqOZmKSy+SD2mT1tI5Iq8MROf2ucB61GSLym83ILgCy0V+Z7tl/LxYs4k
L4aMd5HCUH6KTCGGuttW2Dg1LYlzAaNMHhres9iZ+Q8012omGxcwtV9Ozkcxe03/
GROEFsGQ96ZoA6QmJU4/5tggBzpCbidQMaAaMDM+e3LwYLShuTSQP/T/ZgcQEiaR
ngrN++6qtUHUP/ocs8TBSIHAdUHF+6NzvMt9MJuLDkVwdbjy6ZKjRIycX6Jpi7W0
p4x7toVucL2v7FBg+ppO6Wt54y4CSo9/y3FSs3h/SQtMtoo/d8sv5+WYTwFjNibd
/ltieqTM/XOA9rMhBolOz0nMwKd9tUDJrbLIExthpPMiBch7MSFhHsUJP6uijmB7
LW+YE6ZI4/edwggCNq75KPihp3hfMLKqFtEmWwSs5JRXl2zufKGxHkqxdkyTiPCG
JUafD7K/UjHUxLJCx1dRfzveiTd/PN1EBvYx9VX9tGIg2pXDWhx/3GXf1GArE1sd
GOnxR3PA9Y9zN2NCAfk1FvEskZJopCoUzZOglqRyLfkUVgV1LABrucN2QhHFvSNF
Yi3DlopV6fKfjdyBgbitegZSXh1WxK/J1myOGY5enQIS6AHlR3A0pgAKnmMFXxYA
W2NrLvr4T81KoTSt8xq202XTNTXSD8/m3Nxf+yaCKm1KGQcRJ7AkPOM1LrTl7nM1
sriP/g7xnZIMPo1Q4GjAH9XcBedNv3E5B5mOGSIYHq78x/TqYfOoaP25kGIEM/DZ
p+mjz/z3IaMpTVJI/ked5Vqn3kjXpjEG184K77z7R41eMdpmI0decL+vx4Yn/ZLy
VdVfd7cKLmsT3fe2PN50VYwTkiWz3fWuHYAN+hbryl8EFUPRiRQe9IG7nQ5xsJob
Aq8KLhNNKkVOWGYUQq1yCbo6mjKSXU2Jn6kyIKQ+4Ji4DYZ6lDVSnZYJUl/uswvd
jXHW0DyhPRbrxUa2rHgfrEDjFal3Ou+ymT4jM3Cq6FWLUYFsmZUlbj3Thkfl8xpI
lcKG1fMDIjUGBv+xGsAPMGfap+WIy0i58dLOFlQMEMK7TuvS5JOmCmB5p5Y9WRbj
P8uF7z8tKZnlLiHOJ0mK989NpnffgzbCvmqG8TpGYpX5XK6zRZ8LTRjAxwIWk6Og
XLS/QVlzu9G211FKgtkwonf1+rtvF/r7Q4S2jFfI1nFF0b4gJqSJHByJMsqfineD
7axGbUj9ytS+pwNBE3XaIDMA5LPJyZSCl3rbVRncnqxPN6yAkSbfK25RxVSa0f9Q
XPjdsn4kwiIjCOQBY7JxUfCr5xDMxVD8I8GwLMzoVhcYcoqQW8bjO6ESqYb71NF4
MsLNpQgZFdvroi6b50+l3Jdm3UJxTwQHEqI4yOzEJtY71uc+FCMDA2R3r4nYsVM1
t8p6SGDCIllNdgPYXtfC6r3y18qAqcz+i3cgclw5JZkZzL1+tM3qtGGn4uQV0PJg
HFw1m+EI5vWYLJzHsLP557c2B1jJrDJNwA50rdVOCLepsmKAdUsjwIFOU52fUpiO
ocBLcW0h3t82gKx1ju8jejZOuJTkhTbFpMJ5Hay+IOd5QmU22FjUIdzS16faAOyL
W05TITZX0+GHmBtom5JtvJE07YDPphLyzwhI9/wezDLPWfwuVMTxPu/JF0/X3qKn
Q5OIrJJrBvCnyauOEED4w81N+6Qu8ZWBJcyRrqjQseEtTFMCQXT8qMqAa20ktzca
EGgeU3mV3mTRldiErWvUuxedE3wDm/v6ChE3tYPFdHhzpoXCRd9EykjZflTh1fkA
Zr3yuSQATyUG4y9OiY3MoZUMzjGNd0AyanmGQl1QkqK8kK2/0+RTJc6+S7EvDEHV
2g15+QG607Rmip5ecGulOC8YunQsNPe15SWw8pO3pAREI5NretkEq7Sn3l5kKnzF
W4J0ZbtGqhUSnsSb/oVAnCxugisMZ1qccPrbA/U1ouUQ7Oli5r5kpXUhxXv8YC8X
m/zdS3A5ccdyL+nHXG3Owkxbm1v9pALkM5JlukGhmn+jfdgmh0KG0/zj119ifJRq
rEyRPYVo0QB6erR68mKacE3IyHdpzHbwl35H474DMrisbEr7KjPyjyPssQxbgqZR
F6qjuNICfs9cFRzE4opn1bGcfSJuop4D9b6MxpzGEwc2QNLlQhD+HgzD1hbfulGH
RnHsNbjCkZgxS6dZCItbaF0tUMIaDk440pCVK8DcLj+P7IpTgol+Bs0MwPwwPp/B
CJNvc6Dfciv+J8i7V0dYdoKqFjBi45elHMi4zzOP+4v6uvgXQ0SJWgagRoY/7OvK
29QoSZp285M3GyZl8SiPyufu4OqewKGD3fRDz4MnX0flOebfVsueW2WGM6uBI2LP
sO9/roKmWEdnWhztWOBQunh9Vxy6MCLGStx6YHU0CtPIxCEYwQKsFkPmLWTnB71R
9eSs5pFs59rJKL2WQffwyJH9V2jBTu0qy7XWqCFp42FpQMf+LyDIBWD5t/XFvWh/
oEa76z+Xz4XJKbkVSV1AkfzIx+CQsdHDD/mz7lgOMKj8rUguVCRuzNUy/XM9t3ZA
MNvs49FeWM4Ednpv1wnxurJ1F2/jeFvsEthu4XP+WjKMXJaElza1mVZYLS9HpcxK
VqJv3MynGZczdT89TcnbsYmClZFfvUoYLkT1ZbqpzUfFSIckst2UPEI6AgiHW3ya
2qd78hMUBJW5+URa7p0EzyOzfJtYgcPNVjh5gQEqadsWfFPOzo0xGQRU/pI9XxKu
gpM+e3mv+Wnbv/8/yduvc3urHhSqHExRfFjgBdFfvo05QV+fGAv1dMx8en+58Z2+
rfKKci8MnvbbOTj2gIR4YM1uubzlsgpUA6nSE947LFrznTcApXe3O9mW9lWtn08z
mZ3IWF+r5NY15cSQuFHq0Cd5mexOtwOdgSF5HgTDxZZDAGRQ4KPvuVPTVgH0LaFI
NuG2TZqjc3JlqHW2ThN8KmOsOQBqS0xWbiYVNr0TIHTI4+EcBZGvOm6I5EyAH9ek
UwQueXK0kWta7iWuXFmKMuKlJXqtoXu8JZa4ugrvPPgk+K0IoPRFuonZvCaDWIdS
9XBmOcqTO9ZEExxOaXYeHEnJqCBpI5nRrWPVJlv4E6WNjI3wCKgWnvQLcV1qKzPN
j5+3UNEqYy6IXZtENh/hhRQuxQeCltS+801vxhWfkynnFWjn1hhu9S27/X0lptvF
TnZgD/+KCtV1gKD1IzTb0Ytj0wxYUbFvS4ZJf6x3SVLVIJuL/3/lyVXElO4AmU4Z
YPv38Rs/ijA2TituY1NWz5R2aEe1pLCpb+9wRhbHZOu737PSTspu8oAK3pHbvMtP
QXOnL2gcvFLoIbVvQXsF1/fiFdvLCwMxniyNgGovxvIzf5bgwTa/hlR12V3r/CRc
je7QpQRRnJNEet5eMrLWtXQiW97ZIKEYywDrG40chg4oPXlwWrNJd15JoqlaF0uv
4ZZWJqHa9W/ybdKKQpz7NaxqnDDfGbgQCfGADvst+PtQkFUWB5bTulBfX8tzSjBI
ApUxrqukrNvzbfTiZSft/gvB3Hyc0qwCYKxetY8BFAt1CCR+CAlgFRpyc3mjp5N/
6nHhYarwnjoekFPc/g7SrtNzuCuVVAPo5y3K38LdCcGsdpOl127PfAriZL9c4tTI
3EeP++yalDlOiBpOPjySezSwvIL9mQhX6o9QLSe8vIakgXXsomlueWQu06HSB1lA
uc9B6DjtA9NVKNC8quGD6bfOih8hh4WnaIpOHnGPrA1e3nYwqu/y2lx3hqx2km3I
dbkZ+sBZibLtAjbVuWuT77IT/T/RLUjG1i1Q+bzqs+YVImYSBJtxKboqn6IeWvgs
PKDJKJSWK494kr9subSxTgbafQhv12dwM1d8WBuH2pibOV1rLyxSzTPGTcGMt+iQ
6Cgv3G1WppSFqVNrROC/mAIY8FIakVUa9yIGzpgZ5nWcWVHwsVkE2K4eRoB5opb4
xoo1JfcvQlyPBt9tpoZf1dAAzuh/uQcrtJmyivGp3fytI2XQbbB4lKBRxZqD5MyS
Y3RyhYIzLLGerDZCp9VFmD+ja272peesxMcjqQt1L3IOm2Ls+wozXQ6TLig91PhX
6vNF2UH67PbCEJZu/4dvZ7SowiuB9kwke7Hl6OiDQHdGTuVxwxs1d8h9KhRs3qFc
SBVb0GieNNGu8PrcY0bNQC5ss8wNpMb0sevIflYtl6VbNMpr16xiSDAX1n2lYVIP
LuEt10OoDTSYjhDTgN9dNsiLdTYsv08zjLio+4ZFj/emTzVPTiF9UEJrUNE4XXI+
Hxwlxy2nnMpqKjyrltHMyR/Fo10gv17OxWTU5rykMsPUswLM+rUh6x5+zyIGNddV
6XcxRPSfdy3pELKP08Go6oT1qtHQxqXbYMuGMBxxcUE578nTnDXByLf+1vrajasa
uS8Ix0BIfoqR9395w+4EyA7lyWHiUvK2bSO9nlw4X0ykvgOMRFdjpFNpVuIeZs7q
koJ8DcLl3htLfQPddqy3heLd0THYWU7HR/cDdT8hgSCOujUHzAqRdvGnwKOzLQpf
Gr+vO8+e4wvcYbMfonGxOZ/dTnsqWI4am835plMqNYEGAlwvaCe+LrxVPGPwD3Tr
mwiDBfpN/pficdirp5ROMH88l39Ugja6PEdOGpY6qaLF6GwxoYcL3JHUCyEZ5iuH
/iNZ+qZZV6fVWgcupdLkDto/+46R8IwwBmC5ymgbblOha7EekBlGNfGKvWnfUu56
nkKlETLg0Cqmzo7vpr14e7mW/T8FZt+wautmFRzsbQZdkYfQi1ZR9u2/mH+PaGz5
QROTLan3rnvBR/sFbbE1gby/pa+BXsyYxXDXrOxzrKyBcxCdcQu3/khTroENiq7v
vCoodWC58F7CkErRZqCBee403o64Q57JPmHTu4lgVuYVya2MiwoEJnooXPyKQPJS
AeUpUnOkJE4COe+IR6Dfp4XnIPOmIcouhHDXpHsta1G60/sIOlXKAPztghHe9rgt
xo193ourR+Uwe+KCro7PqBZuLOzoTfDGetBgpxVw+hB1uuY99Qj96VxYut/LTtWV
4TOnOWYAYGc/A9bVoOk/edcv5wUe5amdWTwWkwDKKgMShrZb9IGDE9yQWygP9ASj
8pGNM+TyC26Evs7l9UPKojdvzZT9qHRlyHQOZIhjlykaUxJHNZcV33xdNfP2IPl6
ZTNduBFAERKUq7LOT6DQnyHXiqxwDmuzRTtFYc4xXreeQcOAw69Ji/NBb8FX/E/h
SDETrSlPshkJrhu6ooo0BG89V9H330CV/gDBHWXKBlcd6muNYvjDRkCzx+A3RPjU
EqO5c5RCn5rzQpR3uHIRrUzRJxRoZnwwjguy9c5ORM7vBA7YmXaffxA3hoxxLSRE
FR2qRL7fgCTGxYiMgc4gmMfVP10dzhaJ37DJPL7mQNiaimIhxMZLZ+cESQqYnGV/
2nKK2HN+3dg38CxueS+uh9O9Li8XpYXrorXSTMLLdiUFB7QmWt34F8QaxzcMVobB
/22KTBp2B6mH6Wyr50EZnRxovBacFTRCbdz3Wpwn60f2S1ii7WOBz1Xz+3ZDjQ+h
xR5YUyVYmkEpQgtla5jgarTR0B5pSchLGci1LXHy6yzfu5lBt9E9MI/T7jDZwwv8
LJ1fweY6FgMZXzLTCv33NlpbTGLnWQ9g1RqqnzqHhYDJfbcJGBm5+KTYqt38tuzT
VHaPqtWtKNBQEQSG5lrOitmV3UVHWkGjUWtc3fHkCmjG86RvrbY7v37a70VUZkjP
xBcjjkJfoGSzGXpQ5OSZjbLwUoUP9E+2DAwWcoIbA/97M06rzzXmWS3A9a+dO/7R
SOYx/D9xu3tbGriRBjUMdJKS5+goQ7V3yTrq5IRPNi0r0XtbEnv1V9n30qbUQd7I
6BI2fJau/DPxaKQA81ITwxNNl9Pxs+2FGOlxHyn4Yv8fGSk3HQ66oA0loBHJ31dm
8mmcGt1sVUffCGtwrLUx0ztd9a3f89sFHwzMuCOjNpC5wzLkwnn/m/L7UQjPffT+
ZS/RKfGq65DGL3pucu6u8o2OW2OJ7lbcQyH/cApuuNEMORVa/AUaiuKmjLjEqzMj
78S4eSywiqc6BXsqG5pqmw/LCFryeDHJ43pqCQN5yEYXQjVVjmd7/xzxx+liliRd
c1Q2iS2MVSj7MXqMc6LozG1/nJzER0MP03Ge04v7F1JaPRRMJNWskmxbKsGixKCg
AS23ozyPbHvPbEBFnuTd/6MCl45tuSM0hklgtXy0tp5n2aetDABYurLG9gG9lu8H
tqnpTWEHw1bet8TKGKM3/d/GnWLhCKP/RFPQpFTMXVPmhEcgcuMQiFyyZ6Pjx38f
Gp7mzSOzyNxYvk+LdbfDgwaUF2UFksmEWKPmpaB/DAtNEKAkkYC70bjNLBvf1/sG
5EnhteOU09tr7HwZFf4AR4ZpoSt4P966KAR1n8VAg2tdrWe3+W0thTYuJ3ai5tvE
r2kCzwGy290IwPvCxyxdvZNVFEA5l+OFncXqSld49qGnpmk7C+VNFZXuoYaLXLAq
60xxr2U1Myul5fQpdlhyluCMP4m4XCrcSDjgs0qQyUgb1057BFePqD1L3fhpyeJG
lxdXKKPW/be1Hr9/9kPBxuzIpKX6qgnJsZ+IzHiBz87YcudCaXLooI8KdyP0/X78
fQw/ppB48W/WPp/4IlgTX4CVTCXaI+UW8bioBGpkfEiVIuVtd4k2w1aVORN+FzCN
l3qOcJY7wdPiLKH+YKhSF7BVAyS2FTsLGLDyOg6rV/mrn52FTEBNnfvVJcY23dZo
1G0TzrqGIhtF6WEPTpiY7wpewr777Ad0jxEh6h9ute5DB0ZOqdWgl2eJXJgJ8e7h
x6lQxUvu2jiFbF5H1qR7Iq+CNR2ia8h7ubuGStk0NJ4DuSX+37mntZ3J4RC8we+Y
Rf+z1dP8sf8TMSLktytUjs9GQiaYOVRf2U7avfWaIAFpcwkmM4LODKqi+Yi+5dQj
LCjxya1ivgU/o+82sDPobkWh1KhVLwgEzJ3pPJD+bgNoPHkVVf04SzggVrA3zNKR
fT5nmsuKvcdBE+mYgU6J9wSmLgxpLVdK2hXGSCd9bAo8rsebDjXl4yg/YsyEc/Xn
th1eUdm3SFqa9QZMjPAD4KppcevtI8NI2iHhU3H699oT/KStAon68S6OA9jXEG60
//kLncHavHh3pI//K9n2nm9DXGKeVz292bBp85aMJGuIKotcxm5Kp2xhlk1OsKWB
FT5tyuIHsEOfOx4Kt00ZP4QW32TIU8hTcZZY/fMzZCYf1vQ+7XWrC8ZmUM+M1Ch8
1AwtxP8i9IiRaMOXoj2gj2zmw34M/zHTkujaNYLt/9CiPVtaHeHblyvF5En1F7uD
Q1jse9VINJx6eJAuE1r6r3jS6reZzYlU91hj6ZUkVmERD5H68HNtjsS/lRjcRrk1
uJzxKNP+0E/miOkt3uQkqWi71G+Obyxa9/NHB2sHoClpowcjSKSx/zM4VL621u16
cd9R03tQh/zRJf+1wf7bDwyJRFBf24Aq6a0dlFZIUa+LljKhxrehGZJuYWbgPOAr
NStH6ILUVip4tCQ5CTGOBSzqHjHxcok8tb8tRyKxKHPhRmAZMHwy5k1nGLpdBxLa
7U72roK52P7UeBin8lpiwQoI2/4yWA4QqIVG3HlL57ZSRNntXk+BLrpHTLkHgslX
2HAWelYtF04Iasfe9gZQuJGBGOHvTF79lgNy2Z/m2rCZp7ch6qzm81S1deiNoJNO
7UWgscNvmsH1xvTatGBqfS+f4iNQtQbeODTPS8Iy5kd5t55oFOctXmg/yI3OItVE
rfbBIkF0HFAaVfQEciQ01ZekR6909wbY/PhAyi+ai3R3CQBMM9csP6Yk/gEfJ9AM
+/brw1N0EFLaO2y2o5rYgY9O0vIUe3ZjfB7mWawxk3m+Pw2abATfVx/Rd0Y6okdu
KsuNgWnmgJZrzOySMojHrXViP20arz300ZtXsJli2Xn8Z5MV07H43pekAqBXuhC5
0bvXTcBJKVuf1wBkUiUy6ZGE+v+n57w4D5GJRr85IlPoPJRguYw7K5DJpCLzuwSQ
l1m5zh26YNSX60gQ6CrGdsii5pRrdNy+O6vYPMGDIJfinrhG0x29srJubS3iNGWg
0kbmiTGB4O8oq+DdyX0R8c56lq/hu7m1xlMEoK3CWa/7Ek0LB3M6EiOzttGtIO4F
9+PyCkpALU2fwNFPkJr4zZDyIFip5IIP0tm7bTVBgvVLY5YoZ4YvNtifTFIWdl4Q
c7DAnoFBRFF0EUrPhNJCr9U4hbhD7r6F4s8231o1GwHEaCjeoTDMstYq6wzuoMN+
oAXVpauqLJr8YfnBCbvwDAClMgVFsOsKmQj8u5X/S8R/vgzAFx5iZgPP4/nkVkjq
8R58mfgpYJuS7YBCzpSWyZnBuhFFExROcLTXxH6cQDDuFQhMhyrIlDKEKun26rRK
VmjXoHZRR6Ja81YvpDP0o5S1QnA1lAIwNF/CvONQz2lOOvzlVwXhuyvtkHZ3K1B1
6fGqdJO0pv7J6RSn2VyBGUEU//0wnx4y1DyIvdviYEGQIb+dqAEzS38EtI5loqcy
4sDr3iHBLsizlE3/fwZbpCtzIIUM6GrVvmIvcUK+89SJovW6ktncniFnY4Jfo83P
9GylZGav5gmtabof4SZBcRFyHJCt6KWOh3nhXH5OVZ8IfgBk1IaTH4bRKBfdEkOk
1OtVzjoVAJ6fJvvTX7PgD1T8g/vR7wLM+6CA0mrVGAveCzzAPwpWpJKnaWzVARyK
4YIgEauiPgnDA2295NcBs3uttIOisOG2ObXUoR0GYCoAFe+lykwbPUkYwu8XBy2K
ckfcoYPpy7Wf5Qidp21D3s0pHXzsH+APZVwwGzfbPNltnG3mN0O9hYX2HJrNwOjR
Zr3a726WOxKmfHqTjO1+nPEWRBM6Vlv58Z3r9h3VpplTYxi3YHoh5aukVXEXLA4w
glNRCKM3kGoAqhj+sZcW3U6ufvWxn9jf4PBWmqXe0N9YJ32BiBBy485crStJLxy+
cM4PzqfCGZYLFa84ZZ4S9MXVL8tuZjnQNb1Gh5OuFczxFWgBKqti8cZ7Q/qfaDsX
iWhFzaSI2NGvhWvSdUnGT8utzbm2bjaQV/W/y2orHnTuKTZnPK5V7YPgjXhjU02H
qhJ/WqCBEjLlCAm5w7zNaaqDZ1JXkPqIXnOulCxKXGkv/YjV5cIzhd+cwQomyXY1
LD+7BRT/Y9WGHkRbp4NLFHdsrtAxSQynf86OyC/Z0FFjb7HZrYlNdQ9tnvheWbaZ
kVNUXi40KVJ1zJ8WnKajdc0bsh8gnH8gUtgemiJf8Ixs6EaQrdjLN529ikAGH7KY
0qZsIS3FIud7+g3WMUCXfuCm2WmhPq8FAasMjpbAdpsVDnyKSCfnvmUcvbYQNShc
bpGKihKFRhPzuq7cbtw3fGzVqGkWAjGQtwhQCXv02NOzUm2kWHaYllxEX1h5VMw6
pZZIndFBPfY7Y/tZP7BF8OUXSQOLmtvYmgqojuRMX6RdUvUqoHCMbTpVDsFMVC+f
96Vmcn4frqQbYEMucJ+3CU+t022r5x0IAspM7GURj6qSxMhMUZZpLvkjEj4bsn7z
ZQpRwLoDFam3UBwawn0xc19yDwhJJOBnGF85SAUCZ5fux35owulT2l+sAKklYbwC
A5TjoZL8NktMD4Y1TP9W8ocBJq8nrMIRW7yf9IP6nLGAD0x88AEQyfmer14kgxGs
obVkecVC1OYKfbFTsZla+I/KiAzNyrevIIMIgxl+4//BJRlVZPW/kFLzdPqaJ9cU
TS2cUmgp8Jn7t+VCRz5rGisdQEv1Ha0ciK7HM/UwEuV4fT5QeqPuJMymaqhPbh5G
zNhLQdfcBCCgxROGWuQRyEoimckpMSrzW3qC5+8G6bLcGUr3nmtYvNDz6tbYHwX2
1tVoOZ0bcQ3IC8Az5aoR332Yv7ZMdzwypZsiYn+3Hh3Kwlsu/DWbf3nKPt7i9XPw
teXVVENh9Qq6053RT+TtwS391obdq5ZIgFMiO6vteiyuXNr/tipXMFL/6JOL/W2s
r4ODPRdG3zLNRMItdwNg0D2IuKNv4/RKgTJ7vkIU+1mSjG/6bGsh8bGn6/merhpg
LNBOPy3/vxwxvAHHe557bzFQ7VXNING2GxTXobwNgbwfd8lFe/YD0VGxzMvPGllY
KqP/KUDmVGvcC3WhrEtIj8Ahhdp2kUxMu9czhJdvBxwvFLt4ZLI77x8mZysP4o40
IsHR7k4EJRUWEN91+KSOn9uEv1I8Oz4V0NDkVbVth5oTo6oEug8cHnAmzUI49VU7
KSohA6hDc7Ho/xoWkYrbmlXXGsi1brQk4156baWvYXwgo0SbrkRqJKiacGB+Vo5B
wQN17sNEbOCyh9tAK1hgcBixu7G+tsWzyS2eIXc+UZ56m1zCHyNXG2I7EyYqfU6J
fwRQtx12dji63x2rWIEcfqrWkz2L7PI9cVYJXizKQ2dtrM314ohrNJC/rm10H+sd
M4QFFc2rjPmWFEMg6l3olr2t3q/3RIJWAwWvqYkRK9gdXW6ZOUt3c9lAA8i+VM87
gdZwr5bdrCv7Ci0eKpjI21Y5HXd9PiGuqXWY+ps+pCvXzXqdcuZLkHs6plfamTJP
JD8I+R4li6KBtZxShVsyTbHAWRvsfE6VVHQgqrxOXhIwDvx8fblAQ2kYXqbsnEbe
kDNTFVLIfszZElHMUqHsGtMdTrh65ppOCkXruG/eKIfUqX0m8/Gv1vIWwMrLZdnc
loiBybCkFyBYuYUoWqXfh3EkKMq/ykyqiJAVy0IG4D59b//je5N/ZsJpuBoklVQS
8JTzR3fephYEnux73TjeaCW9bjQrNEcLZ3C8RAYPbwllTt2CLMDxPTEY/HcACakN
MFVUhgimPuyJskptGatj1Cet4tYQTvEHnm3WXlxCk130vemMGYKUUd2dJEdtg+Wa
pIhCZ8yRdPoX+pagf479SUmJ/0pmFdGUhcz9BoK0juFE+/gMED4fnlSNGdjli2w1
XIxPCXjih8TkeV6nHY9rh3XckTe08pERsAV0wl9iapDqenKx8x656o1pI2fnG3cW
p90zZ3jaeKnrf9Cdvc6rCSB4MBES3/vL8udzeAABCOmbnhYsEh0r0HtvUjoH+DmT
CMTJ+0krC3BRaD7MLZ4HBdT5Mwlx1BlAv6GfrF18I8pZEgI/+RFph6DqS+6aHtHD
NrYrGH5jfJkzWB5SrB1bnttUyPoabhyV8z5Oqi/1q6gd3EcF0SAhiAeMMQtuWwRv
1RwEarDkAi1opx0M2rh1N9ih98OXwmdpM5VPC3btW/h9+u4vvKZvpOgt7rWgvNIU
78oAjlF1N2kYOQ85iy1tfOfvlQHadA9UaZYsCAOuLe7gfQmL7pJydeN/m5krn3Tq
Fz65BFt7ncUMak2KDNqVHsLAkdBkHYKDQ+EBUnuSR/vXYBNoFitEeyFHjQ+OT+tv
ARjCOxQJjC4ttnV0y2Z+FLrQ7NgZWfE7uv4DL7Q0OR0O7qLFTbbfsndIKfsaiZO4
2AyDyzIQP+NSS+/XQPECEpaGPCr6uB6LbRPqp99VLVSV2z67uUXiMuCWBkPyLr6/
wG0SZ6fNdat+DHaUPzBYEfe8RCq0td3V0hGf3myt9HJNXBrDxLOfV7indGohJ4ko
a+OVYJTJehRtZgAk6le+BJtaYeYVpUEYm5C2ayze4P07JnrsJ4XPIzPG1UCkGJL3
5CwQ9+HxoV77ldByj50ac0eqqp9laaGXbcqBLhujDkYK0B2nPpNtSOxuZsbZEmfH
iUKP93IJMD/zfeeHkQ4BDERVLBx1A8azeqOKJbC0+6whUUEbDMtwQFUZqxMkV/IE
3C65YBDGTnZagWZVwO8zqmoAkyg465pV2hag689PGH6ggobZGyi1IWxIU5E0VseB
gW2BlyVs85UvHxsaPJ5nPaj63MINm/b5CoP85exbrTS/KC/UY4MVSWtlISDYyel5
z6QVPlIb/irageh9THk8q6juzr4e8y7CPzIrV5+O8F75fMj5R9cj36tphMZAPRL0
xmMoWFOUg41Z2IVJetw8nanVleA4qPamYAizfLvtnH6EY8D+fwF+09UfqYeFNzLF
pdf7ggYTykz+YNvreBWN690tD83YJePjjMskY+TCkM6hBupVdgF2qAx6uNh6jzQ5
QQBeclRTXYev/dCuLeZ53KksGNTUr8SpmAfMGMo26J4KK1JCBNiVEilvzyJuqSBJ
XTlXAjT6nHMmcOUzj/7wW9ORCJb51EssZbUbvC6Vu45E+VIVJ8J28yHtEd1Kkr4Q
RUwCZ2n+PZA+KRBOKg77jKSCE6O27qpoh3oD2WpVPXFDVEYuqCEA9VTK8k2n9hAu
N1565wapcJjy0OnPsFtl0jo2oXOo+BorO509NgQnqhjoinB6komjvIyuSjoc+Azr
x60fR/ZrCreIHZ6UXvfskcYKH06BqFYfmpCld1bsOXkbfOWEbh65kwfkSkQ9p/9i
OQRsEqcaUZGPSagtuT164fg4RzyVP/0G4DPFZruvFkkltUy+NRJsOhEA0swbco7f
UhB6fBY46KV4U86kvzCu4L5WUbJsFxq6b8jKpKslZvrk7LdMamFWqWu1nyVZycBT
/b/ZQylsueMKkj/cxf66xSxiLljNsCnJvF52SQm8u8ei1X13Nz3bKS85bDzGioIy
0ov6U7887YDsK5lS6IMir5gr3ddjPj4vIroynxx/EfaR3Iqy4S5HvOsgLLw0u7CA
+q0Mk3wNDOuHPzLzqFrMKDHvgDQsDDx0+SWMTyqneUznY29Zk23T5j/vNmded6Rn
6zbVYvmIkzU/Oki9bcrD2jRp5OhY8Cfz+9WLWZbItgS40W/3e0QpshIVcwAPXHov
ezB9He8nEVM6QTBinUaFscIbod7//vNmqGv+6K/e6x67m6YWccVOcAgVYEFXDZv2
ZwNQ87a8Is0popC3RYbKh9Po+liX9+YQHAUyzM25bldmj2NxWU5a5pUaQcmo4Gln
XifUDfBUtFlboqlPxeECadGo3GD594Ldct+zWdVbNra3cPaiFyUVhYgHlmiAKxXC
A6ot3YxMz0krWmtQ6TiGJGCiuAeiZtCtWjzVdIeXmlhuuu3iRezbhu2JX+geMUI/
4hTYiqMPSqpnN3CATBTJKF6CrioUjze1fexquUNosR7A0XVrpHXI8UKfBqhStS6u
XflWs4PoRyDF+AS3Q1xb7YsuswqEeLvCoqwuARXK0hx4yQFWeB5VNZ2qi08sj/pu
o0rvz4QRe1eoz4Sh4jh60J1YX4C3WrkuT+nXGgNk5zB+LTl2vRRUaROUNqyr+H1B
yPnupNmh076it9eSitvLLn8KeOrh7omZ9eWRAbiePOd/xoRjJiTXnwLUXJKBZpsM
VyvwfRGc1C5OslbFJvmX4cDDrg/0uhI5P39yoKaD4bmew7GEqzCDRuIuQHnx4Qjy
c43JhMx2pj8uSNZhP2mnWLgbepgn+MGOEjm2sIJYtCvLxMYILTwcy5KLwqIgt3uK
wkQQ1Z+I4RtjwNdGsojzF/O4I12UE2mr2ZKeP07spJ4rDDh2RhRadngKLz5gd+pp
SXunebVE/HxzsTpJF46Ms3kiAlUldL6WMKWZPgy8S9Yn4yloxgVFwMHdT2BuWkGv
ST3Rc8SKx98ICTeIcJE2etBXrL4aoyH+r0HSSfKfMDVF5CXwj22DkMYACfT/1zat
a3JyOh6F5xAnC7/Ov1dDWXv4raju01mRJwqOHDW/iIrU6uWF3+mkqN5HZKozqe2D
02ytL7sAGDKvktaJcjZE41qRg7XQaYi/q8pcvHQo2y4ToQ+qvvHtMDpEdT44cPMm
BHT+Af0cqTd0Xa5JpGeYza7/qrCVCSLksTXCy3DnXipLNbjPpkPCyQ8KePXdcvWj
c2auHsG1dBa2IVNjM2Ufmjf7lYqZq0FCLLNrXKFjQMRM6zHyz77/SddoKIaGH14E
WZeGWzjBPicrRKk7EVXLvScixF+5PE8IXu/dKVx16TieBwYt0/xfxXsod503Rujn
/lpi0SPoqIWH4K3o9W8Hvppy0/bJpjcZfb3+3dCLiBPXuqEAuaVQntBR1WugYZKp
oeiYGtUEAt1LH4rUr+4arx0f5cTBq/R4QzXEprGCM/tic2PvEeDCq0tb2eC/tr6J
zlpIMhuSwolmX2ncbkTDbEI6M5F8JoShRjvYGDxTtCl+rAAMRoBHJjSsLc12rxTM
9SX14wC+miBAu1x1+ZGAU9inXXIgbusuTvgj3zaaCt/7/NCSIZ8Erw29EYkkGSeB
ycKXyFS72qV1YR8HZ5jC4gTgaeAjyNvm3VL9NEcKjrz91mLAuOMEWxB5avSoNAR1
hnLbIM9FzKMEUyK5QH3APMeJjdoXFMTsHcJx++0kERkdLWGalq1jOLzx1CKXXe1U
JerYPiAi3+vV9SXBZtw2kiNAxwxljxAheFTaDdc4gHUl7C83KB4Iir9A7WIZPaUC
t+yadFSTagoF0FyiUR38Ip2zhr+Mj6KPDl6fh/IZf/xw0VIAoJ6UBniLtj/MMAAl
le7VpIjd/ohmoGPxk2YeigMEY114KnH2FXmgjTQCvOnvW7PydgQSgM3z2NvP0VSz
Jheux4ZkSsOR39Ap266294L4N7h4siWX/33E1w53MxIRNEYYq479aZobNvcH1xTI
sbNQTcr51+2/kcB0kPPVct6uFncutgxdPBnDSMLgoVZ6dKn44wYekc6uuZ5eyYCp
Dk0Urt1TvI/9S14BfZ4W9LG+a84SyyDTAL7W1sia9tTMCDZ+0sk1UTk6TE9V+zj/
rPLQNy9oDcpr+Pq+p08Q+nkPvxB3xYfVLo9OoYXz9HSoyaU+eLGahsZDMZbSZgcP
NWWocw6ZkzVAEvBhhnGixusXtqRRRQlSmOjCVa/DPAoUVLN/kE5ZbP2vjiiP0w6q
2QP8fVnF5xsi63DIffUeGUj/9qCMNpj8IFDGBqJzoxgNmCnlYBP5LG9w9BSMirCm
Bm0bgPA2+6QOGjTHjd1M6t85RdtmgDf853J+sIrFWsfxOztX6UeD/ljh4EcOyzzy
yuLP9m3YyUQoS0OHfU+0mUj9TGIyj+l021cnI0meVY/e/M3r525wYsdQR3Bb7lc7
AFW3aGJLzanVU0wuk0D6eMOKaldxJG9e+3s4KU+qmhLDfRvLbPDd71FJMwKDVMng
cmdu1CXmcxlkI6SN/ELs3B6zP3fmG8/aYV8CHm7lYXXXvCWlOULGIVLLPaLzj43Y
eB2GPgPdbxMfqE/qtlxFXQHCuTgi0Dp0sPAPyRsn0WJ1saa9vjECRq904z+TFNws
7SwaEVMUMnBXBaLvSladalm21ep/g7Y4lDWdnYQOay+Czg8FLXULzuPdpb53DAkb
vL6jJAysvMqiDYXadcZ7qk18pm4uvsZT3+TapmD0HXKZEi2xCJQNnFNYtepDlG8Z
P3k1CcPvbDsAWoyVNrBH5k2cGkEEFnBIzbRch/b6TOzzZp6CeVBZ+fhIpPbOQ4Bd
dtXxlmhy0Q/UUk6biM3lS6JOOAJ6iv+EvrDZ3shEG8ZlQfXZ8ZK+rHVqO75QzWYa
art05ZETw3W9K0eTl7dSp0YkhhVR4Ts7CPULVCmHNYJgEfA/7XWFGaYkj6iZelYD
55o65f7ioBFNHUZ351oOq1445w21r+7i7wE4Nu9xQyWn1fTMfAiKluKjZ8Jf9yyt
vo8LVLbh4CorO1JVzbdfwFhXWfrrMOcrwhwz+cYS3d2qFVz0/KjQenZXD3leOpby
lS4p4KCG6XIwxHdcBkCcZ7vGmklxtjCwRFBmyYjVqKguDknWz9q+O725BnubVuQp
kK2j6LDq2yV/233vi55wnZRBRdYBZ7YWdf2GmT4L9futXUTJUmqC2dpNuPje6Hoj
dOsHwaCvuzkMa6OQQ8uwp2VdGQLeARzzJq0E1AbILo5Fyeyrwmx2QXLbXzdRPoth
GFbDYt4NSvbyiThqUbMk48j8NgJA3pXdGlw3uw1YFVp1in/Ye8darsh3bemK00Wk
+ioliyjiQ4OrwNHIZPpoBLP6K5IBQgLj/3/PXaKfs7mOtL/Aw+y0J4ZMPrHlaipo
bEHbtioUMLiiRp5mLWq+6N+gxNWYDtI1PwL/0mXY4MFs/i6GURXE83G6wAxwDgUK
7Q4cG8ZZcMpPFUvMU5srwrzVRMrBhayYqfF7RDeHvkZXA4K05C/KpCbKAfkJoZJN
6lU8d77Dd7Jq4H7HOR4VyPCRPNuwfIH1UnkfcyGXuTLmfNLfPo2U5wUbJUsV59DW
6MqmUmEE+kpwlUY1gM+DegbRcaotFeYbE3tw7G/kdGfUuyMZ4lLD1UKec4UtLXiW
SrxAXuhjTPrLMBgISIujhs0tphuma5SuhiXI9bXqrYaEo9qgj2UgpLO4oUkicFce
3SC+ryCS5cfE+0HOU02Sp18MOCUeDoWpwKJf2B8ksZyvRn+BbMfIlpbpGqHOSXwk
MLVjS8AxQU2UkUrRJSQV0OBYddpf5WAINGJo0p+T/ziPWdSizh/9GhIJAUU/t98+
E/7z8q2grucgV2xnEkurriuK2KWK/QrN5l6owiUDgJ9ThOx/si+mutRpKwTI4NAF
FwFNA5sww26htMGkUyqwVTHO/yGyA93GlZuWs5an2gDnS2lJ0SrwtwS6oc3EAOHB
83a+TFhn6auw5VawPuRCD3S5P2XaXIIagWW+BXGVDYzFZY5UY13t/WZV3KZ5c76T
+hzGlrmTnR/kkhNmmIgoLL/YcHZk3mOvYtpaqP263leN+EnNEz7ZhE+vQ7QJavwa
kljfl8Q9+HP3R9tNyizv2nOCaxgTKGIJ89zsOIdFAGYyuOP+J/RcPBDDY/d7wIMY
y9iVKJNoQHkLTMOB6j1o0bSZr6vQOVle3PMNkvUTWODil8qmNrzOqj5lfI1TrOig
U3GBG2qc8g5UolbKMeEj/ZNyt/ZNgFPDgXyPUwpoAUhkzt5jxMz6kDlIwRUvmGp5
0IqB8aTXyKsO0znd9eYJPLmwO90DTNPFvBB4tCCkhkgGWhHL94vOn1CpFvkV7Qc1
+vRzTaYSDRa/1WMYpPikMYg1eqADB8cdk9ObIe/XVplZWmQMY1nGX/IVWp0dCHfi
8KlcST2JKoQlaI6l70z22Qe6GTl4oyFGXCgzYmPKo7ldtTE4qrCA2VhQ3lvQBsym
DHrqyQKxHYdW/Vp6yY1Lalukamwv32UG29rrafFKcOjlqUWl/PSp2pAhTN1pem6y
LLUCn3vg8VAU21TyrutpYG7NTjLctDi1ZxgtvUcMlni6D2ttMsIGswBOjNNCD0Cb
G9Nt1rOO2BgygqjD5A+BBUoqbG4w0fpouEtZ0tNkYAXu5imWVuST1E4QqPxT7p4t
NBi3X9dl859iW4wp/cY13M3JYPKSUyomWdn2VOu6B0oQ55M1uAt0A4V+1eTretdS
NJvmi5lVs7UOrGH8mcuNARLZG7GsTVEspHb5VaggCYZflz8JcrW7yKAmm3ZgeqZ2
YNB02jXydEtIWKTsmqD6Y0yUnjV/3a4DklkY+9RtCGXjsdcPr5nyIVApTeiYhQPv
OmKy6fbpR2z2+YLhCruKRv3AOzev2Vv54MjKgHnPHCWVVEMH4tFUVmvknWo1I/HE
Y7IxTTQ1/E4PtvUst2qfWqCzPpOd6mbLV+z04UTN1bs1+I12ixK+yErW/yYghlEM
5/m1YAIklbXGXHRzd/z8J95UjZhWfnVsctMdD3XrsJWdKomAwpQplhSNS9Cc17QQ
Z8NNGOkZ7CRMsLSfSbk5K7oUphyM+BxFtpllX0lbpFqTNTV8e+TzxQoVQMrnO9DX
Zctz2h1Hu3nMbvVpONreL40toMvpVNfw1iA+pIwNa8tHdQzQ9Pr8UIfqG6eF4E8J
oEoWzfgZC4DCcCjb4rdwd9HjEtlbJbNXxxmd3i4gUV8UjkFWopwC/HsI7jfeXevz
xWUBJRPunt5Sa1IhN3F0yp0kke8mXXD21FAcP9yAJaKAGdb9jNzAsSEmfbjlbnRW
aIRUSCBvdOEi3fVmy1TwY1CvGNznYnQa6so51c+Mw5ksRlq1nCEpU1SxIUdVeD61
zAaoKI3l3bOJvJzF7JMbv2otlWYVn7osenYgExXT/Xg3A+VWSm2UhM6FEtY/kfB+
P0uIXWyNZ4awuG6b0lgT36D3LlPSJdnjLcKhc4PP047+hrZ5NhS/QNG7JyIGxX6P
DQE2GfAoNuHzZsAyDhqCqPQSltiyA0mcf5QpesBUA9ylrgioBJ4UuqDSYOmYDnJM
m6zq6QNv059cX4JYp5Qi6ulvczn07A3+BftJKAseld2gj6nB2a+uo3DyTir3qAhi
PskFv2IznlUApZyVAEQTiWVmLA2Vtl2NwOKBk67yvs+1npDOopRGsy7Hs4qgOSYr
8yZ6+ABAc/agyQdEzExDlj1v1CLogRe3qrZjyDilLufXwFcSH8VuROmAp1b33gIj
rNIMZ8Wxekgtk45CHZ/DbOz2XLEApq0xfwKG1Uq08oAuS6C0I9ZlOEDQm40LMQn1
DriKe8Q/hTH8MGL2auebqtyl1NiUEkqplh0QXgNuXRcYyy7ywwN2zscjHf0uOpB7
JLB92pMAOtAeyPrGW9tgFiqd62b8doOD8a1ArCmptD+xO6JgBmJfpb5HyZAZKI9N
fdbmstc0MpIEzIzToPFPhRz7vXQpCG6XyDGw1dq5/dHiVmUW/fEkMlYH7G7qFb1G
x7Z/fht2zLpu1JOF5SChoB1KixZ93K0PdtGOfmU7dh4DevcxF/HQq0gOZ7cGRlEb
L5WkpnxXBWjpajNFJTlHIQSd1axUuIx6Hj7hJghgJBGZtO93/cfBAo2gaqrqbaat
pb+T2eCz+iH+Zw+5d6SbIMMDJYhT3zYi2UIgovTfEYhCKQcPOWYqsQX9SRtV2cNu
9He/TdZ5JrnJ2A0pkZQopKyZCB7iCRihAei/Qii5Vti1iucgqHo7ya5U+6hWpPtt
J5Sq/hig0eNLZ4S0TOjmG4ytDmmQfJ3mcjMiPmZRUoGs23ETKwAzAalGJOb0869d
NgmKay/plN514Lyj9QkiSrsqLCoahrbXvNpyZrZB92guZRrVJgoIsJC/oYZmgenr
adqCZsV6ozew3GyLqOjNWhN1LAFg1ZDZ2a0h8pR5Pf0tUB0u6A3A0Ivo89ZJPG0U
FurgqzPfMuLvb0XGoJqeCUKYm9WWxDZLkTFcWH2nd9rwnZVdrN2F52VBNd7G/LLm
jSbdemQbSQfQDgLPio7Px5guIQWyQEWMp7U7EfUp22tepgJACLhWWdriIQ/M6vvj
T3Cdi1FNtaXHutj9U3mUKXYQwe+c74cbPKAP+Y6bgN6SLSiJMoTxRvgBcpoSqMWO
rXhLre+THa6GGY+WHa1/Szl8iCfhnXqNSNiy0FyEcWjuu2QFWzUt32IIH3+YDMYc
DjHyQynXFjgbHvukXkKveYo4qqihlC0/Qa76luITab3n+Q7NwFYL8Jv5p7DeRTHe
SOEXfGmkTnGb7B/5e2WufWSYKEdZFCkZwSAwt4lRGLvQWVPWd6djPHyIxN9J0L5D
S9aDmVv22E5N2R+rM2oIdflOtmhzKoU4MS5R/HoKldNI182TF74n4KqQAiLWxKL0
afcdsnnKB1nbJmfAJxgxaV74dpaoagoxeIPcCJdPYVHHEJFfnuNs3/3ryG4Zy65G
LJYnPUCY476eXrDWmzL1VZc0+VlEPareQ4/wiJ1MrSXM+jAOWy+p2ce4jRix6YJH
htwP/QN+K6Hu0w/3oXX1rBJ1fV9m6Yo50bzksQrPyu6g1JTj/MAz/afiqu70snzD
cHavzybVrozhyXCBRCtdNKnas9tauLtMcGaTCxlyagBnJG6o7U4FtMqNC7SbehHc
8nR7zueeqsBrAV/WgRcZ5UD3dVkqRpqbnqec6E1MnzDpisQRHuJlb9oPxL4TuDZ5
VT+Nd9W99CB+GsZb/qUr3jwnpPjU5El1UCUSxlDKoT84c3OxhppKxRxLFSqHVVYH
B00bXM6mVPzFuWrOCHtvW2Sq0g+kqlZ4iIFyDfbGzLtf9Lk8gIhfNv298yIPOX+F
dHjmaaVWiUNqk8NT3092r/6D8GyyVYXlDQpfoK/isp0mQ2aeBLgtE+IYDv0yaoKr
5DYCqiwjhUFxgEUc9GMpUaKM0gyf1UXTiX5CtMOqzIF+63p/IVCY5tCu3lUTVr1G
620701JWRLuVAJGbmHlHFdCfWHlHDY2WftLxdI7uYqETn1IEUPg1QFYhyoDVNU7m
esh9c1HU6OnjzpXx2kmOSD3BSYd5TMn/z2lO4JLahWGcrbK/ZziG1kKrOI4pFlGr
YOP4WUrVD2aQCJyoYdsUhs9FxWHs2dNJj74HUWMBcPpMgmzmcEPikMG2AaEGAqHm
OBBCIRPPDrRZzyHcb5ZND2uyx/3/FNZQ4/hSyfaImRKZ0J1bhmTwIIbFVaqKVbA8
jqabfV1tZG4h2GLI5GzJ4662vIHokeUzm5Q5o12F/MYVswZyiDgpUFSHdvhsdbQp
1B020hCuhD2P78jtZnAZVcqe4vrQc2FI41ZFbdERdD6Y0mDOfVasemUhB89eTiSt
2DbWukq0nWYeP2YhGXaXk2Y4TnFowROzuUB1Z/SH99x1NyxFnfxYoM8CPeeGx5ta
n1LgDSzTEr8FPTRZbAiww8fw8h1Eri7+HjMJKJvrveMox8OXEbUfMVy18kM8/D0l
q53oC+kBbk2f/evyk8+G5QXA2ivYhsXN2OjEFhgFrWILpoY7G+WiST0SQ/00NwFL
2mgECnvYZxY55a08jkN0iEc6p1c25QC5665W562jW11F/CnVqiN8BCfTP5JnF07s
7dKrLdnEJ+Ac/0A7QFzR3T8z0/QAZGzQ0h0ckPPV8wW8ntrF+hwURKTKxqOlnGgV
aU1fHZ0yTBZqhliatDnPHb1qn+3jnWEPqrgagBUxyGTH8ocTYaA80e/ajGaYK/QJ
BjKva6yaNfa9EiV9bCdA4kP1aBaXvW0b46Chg0bj+pXwMed9ruVuw/n5lp8rHXlI
kZsU484fYLA8DEY1/wdQvZhr6QWKzaQ54LyhNLqvbZp1S/dbLDFomJuL1jNBqJ8j
63O2pQBHonk09qbTl9qppLoA9VYyMggJ8TyaTL68TYkEGBmfnr+VnCBmDksrSfYf
llYVmlHUBwRyk7Vb5yUaGWiriJftDtllYPuuaaZ4u9IHUHKSvyuIo/rv7LnByomb
Ve00zs5zn2mERXnXnVn5RJJYQVoxwQfd7GkZ5SO4cC847Op9fjBPDN0PTaIkgpy7
q1MBH/0sqCtEOMJaae5i+1ZXIk31DMAGWBrMJ8I3vwNpdfaCAHb21XGAarjjvdy3
QAP9F6y2vzPpKWzmiTKo/zRsigKBKnFtKEAZlm5PjJ8fGFzMs5NBxuxdrhHTtGsB
puk7geOgPE+BB9urf6QBx3lv8o66U0hD/ToQBxbLfAr+OokQz4Q5fq0GjTQz7K4c
1A2Tn00SgtJ1XO/H5H9Wssnkp4W8OQS34FamSKbnceUHaebn8db7qTt3tKBFSTre
8iSK3xBPdUVawxxNVwODypHu7yylHAG7qDmmQL3PRZPNp0szANQ8ptYCwNsAStMW
oWEbYhRk0lh2iTpY4drFKLFkEWtDjrtwhLqXEBQt8+oL4nOO5qQjbt3q2nQgY2f1
eX3ZTfmHg9Jfxtl+rnfxNSR4rxQKMDl16uf4Y3zASMBO+LRhB4Dmjamz1ubsvMm2
Nf8/e7ipHAOwXCENHwuVSRz0nfHhZtZhAyjO2NZxwPXKOXjt8MSXEJRSw+UwPfxr
xp8qGQTUJ4O4RDJn76MhcrMTBdJnb0FNc0IF76rebasGdPbEY8p4qhFAA0GdtlLt
QGbzq5xERmtCN3Xp2EPs9upVJKtXf3/v1/lFu6rURfUhM6C+DRLOXEBOiHfu/HZy
0G4k7xcqFogjAAls2PfnL6oOaW1EdqBjeuT9CNO4E7ip2LGfWYwutrnA5YaUGr8l
bj7FBhTAy1aIsmllYHs858L+GJr6HgZvuR2zGHwLoxPNHeKoXXiMIBHp2SQOSyk2
P8mr+FfTliQ1NVYCNToOMqOU8JNAgZrOj5cBjfWqhmqGTOhiNagns/eTIyWgxttx
xqmH4virLcZ/BihgrjD7NnZosdLNOCbkqBk8tc5Dk6WGchUlRYHAz6yE47xZiq3W
7jQV1LRC0QADAm1Wo/UkdswKAZb4AWqMwt1ngBvxiLcu94MECTSa11R0pexvpiHg
txSbMmTAiuhyDxhhqWsYJzstaoRiJc/GoebHXY+AJplgy1/Il5qZnyrAAPPoagb1
Ew7D1xpQB5JVzQbQE4G8dWS2obslAVShy/yggea/W2yDb5VPUv3Mp+K62xNeCTs+
HpxnM91XL0HhQmso/skxgITGG6y4gKGJ51iJHePfSTika7nkEJSPnPEidjW9wOvj
tzVWwwLXsfhTLI6we7x9bwcbtWy9M29iVxCtbSklUeSjHNyK896DuJ/lo0IKftKB
PELfvihSUk0KXBKrolmTmq0pQLrjFF/6pudr9bxyem/cS8IHn0LAF/5pEaRk6tUA
rBz+VyqzhhVA1BnVr4upaSwlXwgMq/+zUpEP0itctaLaujdF4dqbe+Y/aglbxHoZ
uyAKDYwJN2kTt1LL3Keb3ObpRk+BuvCSvkbW92g3/6gCaqCkCYwud4iB6CyVKvSX
Moc2+RYEe72Og0iWX85D6xew9iH2xYzxc/jmdIrjtxwYrRa0whHYZ2Cmjh8Wx55k
yHp8ubVmSwx982kWeEcYyG2w6rTrTzk4+NC4izB8x8kIBtQWhGFEhfKRVbMTl4dO
+oqeCp4GVdHx608muyl2sObzuSTaGvAo/10YYgvb8sn2NSHl5/85xa018QKK2AHH
tT5zZJnG3qYxS1CwKTGHJjxytL4/EMZ4Vs44vfzvIBjJy359U8zEm0OttbXsMwcp
a1P4Cvi0U0xlKj4gUVPL8RGpw/xKp9RK1nIeVjYVGrMsdicVVlroLLtZV8cKGJnV
GY2mp/QpcBOOF1RvVvRDWYOx4MatdZtYHLpO7N4vADfpIZbAMv2C+c+YPqMPFeWX
25R8NaZJT99aaTLq65CsY9x18mEoh0e8g2ORvMiHxpjHUUgrFfWua8195LWbT+xm
aPJQuJfyVZseAAIlG94dd3DQn0OCQCXEOM31eacLk8UbDvW6LUD+Ys0Sv5DP6oYq
Z2f/HlZ7cpXM3xR+bu/n7Z/xXwvUk0lfJJQBuJoMQ6ccPNju++eO0aUYebBjs1jV
1XZB+Z31IxpUWDIlZR+X5fyb+xeS93QzZAewFbdDlPyOq5UWl/6zzqyZGQ9Wrs1N
CZ/+dN3ISptYisnIpbq8eE15dDvVfgG7qj5ysebr80+/pCYfoLDFvVRZ0AVAXfWN
Q0A1G9VT4tzsVq/Rkuf8CRSOReadCYQ0tc29AwyjmcvK4E+1oFXCHxhTXWOt6jup
8qnUP3Mpixccxp38/SfiTl48DQFQNEthxeEkc823PBMpWIMG9105S+bpWDRjuW2d
NKQYlPQUSjxel4f31z4CRD6AVm3eDqF+yhAKnrxfqtlfNYk+xjmYP///9bZWLFXm
3T8DPdbvFxWrdEjdQfQMorvJ8GBLJcSZRtY3r+PRB0HAg4pspoC25JPkncW4NJjs
TN59w0IoYR//ikRNh+ZVOxW4sl8Ba1/hns72vUd4OawJ0vZdPW7cmJxLoxROUqo6
pwYElMAnB53IJZuIFQ2AgHCulC4mnzLVZhS6Xo8Vt/VYfTsVnA3Tb4c42AVUyl54
wzQUdYIwyu0LfPHtx1k0h0cxOyJnNJca+DLBkNnQaTM7UNTL0/Lyp09p+8PnqSXE
qhsuSn2JnDCBPja51uj1090KE2HXLskjsU+Jngv7ihc50hOKnPftk4YChRO5nYwm
fQWIkepwieEQ2RjMo9sGQ70PCEjejSClZJ8GR4u8yxwCBdA9qUQe9hNGPd2hPAf7
esynZvF2tFA6tPCxNkOPn8l8dd4zbst/SX2anolpWgRGD/UwQJ4synbv2MSM5sdr
iY0bRANNSeDn72xyvSg0T4qdiKLxD48TVZVTTZDu4E61/EEhb9wWTLXWIw17Aupu
XqQsjtZ8lPX5mCFtL/l8o9VoBdgtVQyEQYzNk4a/pMp3/Pr2dL+A2K7dvvxM/qjD
YbjoFo9TSw5bygZ7UPZvMGHuC5fgB0lvZc/Sp89YqKQ6uy3XiusHS0ygNST7cDzP
+09Nspjf4jO8bZuOQbNKWtDywU/EYxtrfHJQohHCUSo5ekMIFw+lCRLB1PfX1XZ9
CmMmgHgUQ7tUamrFRKMAWIpMZP+TNOQZCJh9Gqx1yC0jA1ndqT4YMbCmNK2r5l+J
LjMDI1xBvU10JHD7mODTJyiL5D1zc6xFpbyJEBccHTidcRlwXZRldZIiF0DESiCt
0dQL/O/gP5Q1AVwQubFe6Z1GCRrlcidIDDfwyVvu7HuD7twSl1rO7UyL/7XIWimp
o20WVqa5536T2sLWIlH3GORH3wGlxRT2LUL/lW59bmHLvfpyyRjiuvE/iS470bL5
zebDCPOQDPoYSKnB0/4GBJ8jrDbwgI61EXzhx9J18ERK0amRnHfBNw4FwpsqYXny
MwjQM0UEL1bFtvQDPdNYc2Y1hDoQ5AMBZR/6d3U2zkn3lAbyFz+h93pDo6wDixVA
zg6NGVih/8ECjmF6Lb+t/NwsGnKHUUG+ncT0S5NKuPyshvZsnL2qrT8S8wDNm9m0
eWMssP9kqloUwq911QW+Y1kK+oWe883mdHzJD0oBKfKFyeIJ22qQhZxLn1vR+/vl
04M0zyF9YBq/2r07/qDgtePFm1GAz/2qFk3aWNV5lTmL9eVlijZYT7ctbVLZGsZD
IxjzvGJVH1nKEeyaQ6qrgbo31JDOgGX3z28HToK7ZHAskv983rJCRVxyykiQw//f
AxntXAY+7kP4BUn8TAQpe+9ttsW8ix5wXPcsWtucaKPcTDQI/XbZDiVmjtkzwUjK
5zc+kv8WHkF1Y0KmiId5MxddCOu+mRRD0e10VXMu6pZbwor/ejtsQipY2axG+9CR
2jOtzvkInPLCsNVCbXRuQRwYXMmnQBkU0eKO8vN6o6WstAgGyrJz/wUB5OIvfXBz
j7ZxREU7Yp9Ov84u+vELLoKmFirU30LGGzo58wHTZm9mIj8XZycyA3GPJmw5/Xlk
EL01wf3XMZ8mmJHHWQeuwcS6h2e/1nIt70E3GnSccvEv4UzqpC/jCHB7geHH9h+B
XYJ0TBEFSiDoxnNZ+9jC+YEom+VclEiWNh50ZJiBmHb/LwqI9+1Xjz2BDksM34B2
Xyknfqaz3bhQB02qnQ3cZ+BkBaUa7TubtwsU2Npkrs5kBRkFS7IawTg1hqFfzcgL
0T6Cdrb/1Qv3nivTpQceybqRRf/INpP7xDQcPNmjOf8EBEqDRfazcrGbz7Zsxn5P
/42Zl1yrJvawSdY3s+hqzbJ1xsg14AZ8hVAkBZpV96qPUt2uKXW1V1Gd8/lTHVMd
TjIlxViVH0ggEGIYc13yQ55AWv4l8nbZgM8PVupC3DUaRpofO8tCj3WT9HMCcl+7
8Cc3+duta0XF68MugeBbsCd8v8fU1tX8Aa11+h4Rak8vs4kVGiv5oVCmnydLT1H+
1yorukLTTGBszjf273Z7N4HLRhkh78lPluc6DdKm7rDcJO2l2dam41Do4EkU/7HN
yd774N1N6Skf0Xb4JmgsrlbEPxb/Quh8GHqn0PnAUkSZUuUR9tmXwoa9g8u5ci7J
5YkSBGQfiZwRwtd6ZLWO6X7/Lt/TiNyKrJuS+YQXiMQQuKp5Frae0TWjUWhbmY1b
zlYUkknPYqYsECJ9/TYy5sKwMeSrDbTXog/myqIQQVFVDqxXrUTfuBV6PLPnaKci
DassIT6sSDNbOFHhgpo+xpdmkTDeGBA/x58f418TZrP13Ur+hOx+rno8W3ViZ1xY
/uFPanp63RbILB5Lhc2+DobEZpJos4t6FRBoFOqdz0VGB0O5/wWD3RDauWCwNkyw
q/CHue2WQTy645DmjW/8IcVEQO6bK409QsGDUUaG0/9po4WQ4SbjP2CNguZpnzem
UJfa2ChARkT0mK9FYfSv2MYMZT+YKUpPD9rVE+3mGdL2i3UBgLQkSuGWKtoY8IgL
PtzjRYZ92DFKzEilr2e1UN/feoeokCS/8SWXftfjb2OUpqbktYOEA/diezqqeGQv
lFiV/nStrwGKFv3jRMGAg4Vwu/M3++Mreiw7KAkeIqj+DmcB+qvhQlttNRA7Ejr2
FCaRTy7Lkakn2LMA66rhS4hdmBQWgNb6rwuM4cnPfqWcjOsYLBRRtowC+WxqLFPL
sz2gOAhVfNrSMzjgEGkkkr4hO6AmcVvxglO3gtCRZ402PnJp7U233YzbVBbROV65
lBNrzuyyTOAIS1o6kGlvMh4tYg69gGLj7CtyIxmHiD2Il5F6UGVWxY7c7tuXK/uo
EXgQENJ7Tv5Tg0vnFXSB6hC7Xf10bFytEZ+8iuznXeMvVlgHTXdii3adFhkrI5BZ
dOhXyGpbMElF6Wu27O2l5kAzabL1ZzGKUnLT3CVoJO9y4E8SHCLUjAAKn2V5NsnD
q6wE6j09MyT3a0oanwG28AHk0Z88dZNqjOfvLPeYkeGDVknxhRYaBql9kzQAHtWw
XcEzn47YprF71IfLhDYmFOO2bhlZ8oXHbMnBYCeT3Yr7SRh6M/Bh+v87Nlj6w+qu
Ne9nFqaAYWpbIZPf/W4aU8ApAynNwrIU3/VsPaIt6TkhgjqkRyYMLnqy+LNgXsyF
C9/qRDOs9nc/9RlFiRfkX84oyQM5iwZLICSbopi2OBMerMZAUn6qVuoIPS6MOZXw
pO3yqWNbrIMhhCrJv3NS12eXzIuK2PjviKDm9TnFydyyIdlsrnSNcSUXPEv0eG4j
zi9JUyjwMXuQaa2jUASSUe3jljRjqKO1KaTs5A9GoGjmxCo7/FG+RAaLWUDdrnTG
wkEbZUK1MspjuCdWdohXLhhZDFk/cnG1o7fZV5riLxGQBdk/MyPxpdH/Y02DTNJ7
5TUfpzJo65WmrdqXhPPkuZyfG8M965tWNuwzSy1P7H4XRwjrHBVKtUqy+TmnrT8I
yOamKSrOIgIO7yKs1uOeJhZtuHfZ+sGooURsfsWOpigjYCqa877ErR+CnqbTiBKK
BSDghSrclJvHctIXCXJrEE3oPuAPa9ANdWCStdzDwqwlzv9bbdBMzYJ7M6JwYL7s
AHnKIupDjwFYRNJSTOtsnKk+XvM9HN6ql6+dDyPQCP8fgSAWXVnKMgXhAxYFy3ZI
IN9SSZfmCUFi4wf8+WHn8QJcfWtkfF2f/nwm0pbzGTwr2AeU0P2Bz9ZiCfnjvw6r
r0y+gVfCDHSvier31vwTY0FqhlepsMB7j51qgdnFY0xlFoyiVziuKkHTCZ6JpSf/
5d2BM09OmVFSPQi7qMp9LX8NZFLEpILkLSeOErD5Wejk81hX+MRD8b8Y5UrwTYkH
/Zl8VaWK2Xlw6ZDKohlo8nXWVuBkQluasSNjgyICRorntPK/No2z/7w9AN/KgvG9
o0EOXwltbpLPYM7Jd+Bb+ql5ijjvbffz89Gr2qq9/mXgCz244aRyi5NZpLeWPem3
MJtxvE92Yijv6uknKvElJVmlD17qIKhXqgbSkNqt1rgksyEiJkblkr9YSbwQxjPT
cL20fSxb32VWHri+1TNYNx5DaFay+tpgN+i3945Wn9JeBLiCNLiFPCQ8FgM7kHAD
zIPSrY9CuOBjAPws5KotJwrswJaUbHFP581AI84GXbXx7Yb4OKcAvlB+phAzZ1rQ
qRoR/jo1DFeC5YuIlEdLerdLgd+O+HyzPCnG3IuA3UMMGPcqZDjFJCwrEBFIgQZJ
Z2prrINPqzJPKIcaPhJzhxGLT1Uj9Ky8QIhvK/O2bKDP4If5yO+vgiRPcKyxDsg+
Us6t0G4uKTXvzWHh6vBLsLI16ZkD/dpJkBHNfM2Q3+M9aVDHBCkew432CTrHO93g
NkKEPnXB8eQOIhtLNpLVLpDBrSP8XFMTKsvdhZYEaA89pC6bpDlNXf10d5viwdYG
MVcERj3j9IGje+V7b0W/q2UDLCBdYjmP5VGpUDGfYYkRS7xgT3S/ea9tNLArxhrq
3pY0aGQYpL2gWaf+iTFvJ+Sm1lQnzYlhfV7lH0vbPKfkWhfIqn4Nu1IELLTOOHam
kpjY5WLHFqo6dGUgYsGB05zLZ9IHaP/p82WbEv/9yEixWNZ632rlrfU+hrXDIxw1
78hOyAUBHvNMAHOgj29lM32BrQgcCtUhTyCRAzWSWTs9C+HDmQM2Pmj+s302w3px
R85hvzzk2suAPw+MLVwIBHtQXQJTKoaFsqol7YJgsUABHqTh240cj7q9nmzuMbCX
2FlhktSZzfWrKhoU60HE6Dn0i68GevsmvDR26BgBxRsWWGjjJqrUNsGAHHNsb/wg
t1kUJITKLhpwd6WIWBLhMMyPSWzJmPXaPmUUwWHw7mjj8bMYzFgELvUsXOwcvfND
kFyXblRhQwsrN0DjHeTlC5PiqiqvHQGM9PlYns0cVev3tn7myBSrhUgHH2v/wcmc
9yzIpNwjlZp+xc37je9CsN0jUfvC56NQUnlgQmQBDJ/w0QH8VjvcLJ8Jgo5vaA7o
8XpBydXC5/Jm955fNiEyLqWI65DOClwYGxxQBXsCaBFlPyaPK8j6m00A0J9DUSAa
fpgNPM/CH7pgxoahiLMiar7TYzJs9J/q9k3VeC+bYe/r8JgB4f/1rPLNLAlj8M9+
VONhAmybF6O7CodjwqgyH0Tofjd660zlr+CKSV1UT2ZeJ8ZHl4d/GK+9QCsOuMC2
8gkTeu6nBwNnhHjmg38omMa4Fbe4Oiy9ni6maNMXC7WhrUo/MqT8J0rG6LEmYVn/
oGF91QYy62ZKXvRZEo31xErqbkZlmoqLCCFcEqDyp489SZcOaWlw+Cxblc/T86Yn
eWIVGHJGLophnUNnajBjPe31sBA0ODGtNz8pyiygkdOmfP7/ZFAfxHbCjPOR3Eft
bYSvSeP50e7gSxBPYJitSuB9HOWb/FnOrw2eCTvM0JTp7Qz8cuFpkq8pqlzrJzYT
LnTa6V3sgiSLPWM2Kox70neLfach+OtDFAd/vfDfVt0dxv6OrvhiL8KpAeEfyawM
eFy2ImVoTYjXgumP7eLlLEQCN0x6R2IwtGeubNSS53juQzKvGTs/Rc48WQSApCpR
GiFFJXkksGkoIwxID/YKGJkgYTTwjHp5CJy0l6+IVqwCq33cDZRd4KtS7vYb+Crj
ssjM12QDuqzk58xPZiut1myX9rM7ZexSi+soZvRowO2v7bpS1ksITtPaLxzQg6dz
aAvuadxuMNTZ/bhaBCS8jU64+OBnkn7b/RIqvAk7tPAmkBN97phOLy8nV6FgyLOL
BNc1hlxNPWxC1JBiFjjH3vGe2zgwMLZZLFTzVqj14a40eZzndnzHb/3plNa1Gqm0
YnuPD2u9AvVu2fS/tuLm80x3EYzdGhhpTare7ycK97o65gUhE1/SvO2MiYOIPZ59
r2dDP9COmPZodsghkoQ6xdznYCHg93qf7dlB10EgtH1JHHv6oG6JXIihmLtFNgzl
xXjKmh+IOT3dPttUFs5YxPCQQUYv6CP7NfLFIVb/QsuFZU6wP2tzPW4hQWptUm48
eUjS21FLt3tnBkfcXJoGk0Q1hTVYZHJ5kdfKYxbMTe9j1p4FLCPTiW1EAyo6LJHx
Tq7PviEtUz+FB/LrvwgOjjq+WCMoBmaQD5xYsKs4RImolRb7HasGRPqwK84mib5v
FTZMQraL9cGnV+CdFrc5KuErfoBK08Rs1sEyrHe5VzZqesUGRgZICGEZM54icHPJ
RrXRsnlLV+uqWJ1BlclJON+OliL5Or6FiATmYnLLNmvz9i8XEWu7e3sN8Kdi7FTz
q1iil6kNeb5CjoRXIHhCSpdTjZkR5l4xP0HxhGLPPr2ZpwI+a2dlUvMsxBxfIXZj
5RCwnjNt21j4cZ1FEnqbtYf5vlyRoqwe1tHSxnmUo7Q+m6+1Qa2sF5ylox/wTDKX
pZ75vXYAm/cL7o+Br5xGC0mci9nUJqdEbheBZWt6HPNmnAp+DTjOzzAqWQWapl7h
WBSqfpIb5PS2P/FpUpNGWlfQDwhBrP/a5hyXmB/KC8nYROfiwE3Rhdk9xRZAlyC9
UVOyJy7OhRenvI7Bjr/KOxbQ37HPyi6oh+HIgJqRHNJjt/MNepgetGqwZcrxS9Uw
06o2RfrAUfnO3vuahTEyA53LumJyVv2JoXxTps9PZgJlzaL8m7S/zyH+ncOMUChl
sRiaeTHCuQShvMCCUXbcKqaXw0JWwaN2QkxhWhXQ7gt+b6uFtayskJd+70+Nsn6L
2ixfawnmXprs8YQwDOfL+EwvEjPJ1y2JKx9rudgMioxr0Q+rMWKKMVA1rBzIpnr0
3RAR7n7HxLlUQvW7v6ynKDUyoIQiRKOz60XU0czo/661TkAsEFDE0tjVqfHl2Uo5
krMft+vJWCqFdvSv/BD5tF35Fk09Yc0A2N7aKptQ/cxLcSQSZxmLDQT0c1Pd0JY7
jRlxNyyoBOs1uK9nBSAneh7gNc8aeERsTYE5wX8T4Ks3QGjZEiW6rUkqBkl+iJXn
YzuGTaL949Q1528vyPzFTj4Bbf3Z476KnHPeaOwl6UqSZitPhJV9f5jrLSiWPGI6
94K/OVVWc93IUXozbQjQ08r1fczfk4R5U67YuWFcDOGHzYAEWJx/rNz0SQ9ta3vy
vagBDiBMWrEhD2lFc44K5vY/dAeakKH8IUzXM7yjVnTSlGVghI0nmnUXSMWJUB+K
Crlqx4u/P0Cdq7E5Mbn8l508TesnVSXnhqYha5dp4IG4lwTdamN1Dj1wgSJj+ulC
QR9GTo77MUcIzTJ9jGiRsgpsd8i9sxn3BtyNhZye5Ymort2BA2lI/sXTHE09FM7Q
i4ubs9aSvqR8p1dtGoynuoO8z9lwAzETadxOvY84txYRrg8uZvF3L4nFMuuhEKiL
J/beMIWZhCy/heGLCenWUT00h71Ql4wQ9MSMCzgtzoyyiq0zkbZCM8QuQAQJyNck
QcpIrcdzXWrPxn8MuuhVHLazE1r9gQLOQgcZLW9Km1DhnZIQJPGFB2CjeUGk1FH4
mP57fOvtM1sWemnuOMT3Q3Iwz4E7NnlRpwQBpReNeQF4Ye50Is/tGv4l/n2gGoXE
nhNmXjDj2jJVwrjGNnFAMryyYlV6LDtcngMmXl9TMhdtmyzbxtwRV80a10Tuaua7
e7paBeyE2OIe4yCgL8LkhDdZt0rovtL7c3pEQ26f9xS6QiC/eTiE8UARUNKROZsM
spqLfoENkqWgE5LTdEmk8JJ4yR0MUyPSHuh7AKQCVnXEaf5MPRk/yoK1imqdzjGg
ui/GfRXXLpc2OyhLJy+VeZM1bdPzK/eviK6mc8+DNiSw15042eb00q+dOCabRS/H
fnW5ocT3WDJ1riELonxbnmtR3JpWbzBnCddJazCdOWJ0omePwCFgGllnlpw+A9Wf
06WV+b6NzSpxbZuzvmIxftEkHSA5w9kUO/lh6qIqBYFVi4+dc8Ycp2RIZANvvap1
ONJR3ItZ1xZm++2fxfaAWdWaIzSjJqLnphV7dJromht7YzWyAl4Xto/lKMDuUJMN
+M83p2QWdncV6RubQt8XBk9BhKX4s3pKq0Qbv1MNoRiz58cg+2NIMF6+SqWK7DCj
v6kvyU65McmdNZW2wwKGw5b6AgdGEWgDRDJU+Qs/NXh9avediVYWopG3DD+jhewJ
3xFsbhprdeOmkXG60G84VBaa7ezs6KIRgc5TbyvMKXLv1ZGd4UClAfZInUFoAjiI
P3Cw/GV/OAwZbE0+RW5zL31yuRGPKdBDrLAgdZCpBfBsgwz4R1NSHDyzk7IMPVVm
4m7eROwBvhhYsku4xy3SM1qSPhLBdR7LlS87HSur/xO0o6ioRjGs09FvJO7UVL16
HRR5JkggNo5STNLpBx+S2Yxgc17Fyka/EColBnMbWfIYQtIU7qN+Pj5Gm1p4MgMd
7nn3pBrL6s0dzKxqd6heylo5v+BNtEslaasSMor6aBLYX52eIg4mbjGEbOKszQNC
A2AaJxyhEvYSEDJjcsklNrToS9wLr8wiG4W8xEO4q3t+Ml22fO65HoqleEI1B0i4
B5b7JJMSEvh9ZEX9pT/OD7kp3rvmZdV5GJxZHow7VMldp2rVrmQGFduxUh65I68f
NSKrei4GYYWGc9kLssjc8grGtouGmKKjXpx4NTLZrl66lPFqHlE3JS93bjND1+pS
9Tl3Ggw7qQVhK0B0CCmb0NGwwmDo/PnQElml6rRuD3Hp/GxB3yJAlNXAl/iTcyL9
/Goz3nkJxxBSDGkINw42Uwpx9DutdHGnordH7dOJ7uorBCBX4VWkYd7C76esb5m0
E4qaSdYHzKOiSVwLuINRsVhitlhGgBOAMQkdzqwQT+yi98Lg6I7DkBoKNGA+oD7M
vZf12HDPVefTPUqPCukFyp3gpGkqU2fxhku7YV9t4g+2HwHqeVSZuQAkl5fixSeB
KGk4SzMEQYakewCSJiSbBA5ZkQ5zRBSAvUU5llOmVWdS9oR4JmwMWdmbHndSfFmK
nVLuWw4ap/z+2vsMbiuT2BRATfSyjhF/BMcNTVw3pWuNnGpWu1IHxi+xe8f/r1xt
cbWjTyQPD/oR0zvyeLiBTaObn69KvP9c+u7cQLyHBqI8FWyPE4abXwXac7EuclKx
3UTQg6YrobtK1BlCnlnk/uF9OZR7AEvWmlOdztkWY9zMgfEnMXKNtw/90b8kUVUi
Ma9FsvMEVNLb+9p4y7rRq8Kwvr7QjvnUfAqjkVln7ARuw/+VF1Skc4F0vaJjg+RM
8Taoz5Yif8RG0KUgZMuhu28BXJlJK2ktOYP3lRb9BYzOMEMsgQ7viPYFtZlQbR9w
g8A894+EJGn0Ss1qCEPEIjqoum9ykSh16Xoe1teVu61QNgmV0UVW90dCmBrwObH+
hdctNvh+ihoWww6vTHCctD8f75WXCJRqAlh9zs5OYZahHFhNHilrTZsYbxt/vQ+D
DxTo2EBZqYkGL0zXWUEP6naSStX4zMfFKIuuoaU/Owx5nTKq/XW0YVYZ8Fe8p/vX
lSSL2W206TOuaPnVsWo+R5Mdoq9KRJujTZJNvi2ceq6BBkfv4dhOfVpzH9Ni1Jl7
XgZPdVDvQKXG6CjyCdN7xEWe9wO63MwSglGeQZBsplDrii/B5bCXMJ0aUYgYvVnk
BHE7CfRuIC7kGbXdt5dzL+UdcY3+X8Aj/Vm8UAMgoXqMZkhLLaSjo+YxVjF7kWSG
4xLTeree+iVw5kgpu0ZwNhObn1vaWf6i5SYCR/hVUq5lKO/2pdQS0JBSNiRR8hWc
Fh92/tGCCdw6U2lRNm5LhVL1zxC2s23eM+Yf5gd/3yjzvXL5Ntc/gJzNxQ6Dhuvr
z5Ibj48myk6rGpdf1kGQedd2YsqGgB4C3kgbChcn40Amfy0zHzrJrmE6WbT7GJvv
N72kLew3qvGHdkvaCurt9eG6AmDGH3aoYRaongBcDc+DOvzoyzid7sapyrFDrIYg
CUXet7Ax8d+gpJ8E7pOpJ6mbqvahU+TZjSv4vsR/RFAvpZOoJjtGl+2UZWXje+mJ
W7rUTFvUT1BKea+OBPNFLNkxhISa8G0QPuQO7FAY+UG+jskK0p7jpjChl9ngcuOH
Wj3DJ2A96kVy3rrAtfgX6eqoutD5WvYONqnNbVjMZzF2ZsI3LW35z8w6MZZ0Rbfj
Xbwomz2tEFTg56vtIqs85dr0dJOaD2m8igle/wHI/FPlWu2ynxlwefRhaXJaEEfZ
rGmRI2zWd/WLJjVo15KRdaWgPmx99jZGVa1114KGrxsRF0QhlKobJO6X+Bw0/KmF
bZFMHuZydyoMu46K7Mvn6Lgh9lQDP5orZMCo7QfOzTLMfEDNeGaX1cF8l8SS5u4c
WmrcH3YMXHWXUc228zv1OHRahafFxJJrFWi7GnKuHzeR96e5iRuJKNEq7jP9d36/
uJW6qZai0Eso3uXBUWcLtlBZLQ6fqJewKMxsI3Z+/WtkloAmEfoBeuOy1149l/58
LahcSRCVDugZ78ttbRHvHjL7QRpB2Ed9cwAymNRICXm8a7NJvTeo4Zf07cNcTIi5
QRnB8iZWh2HMOsK28ErVOoTyKxNrZ9XKd0jUIBdNtC0A24Xg51qEm2BQZQ5xso4o
h7qfSHiGIzCRF6pvYrolawPIyvZv8kT7/aR1Splg1PUFwLyEHzfmNREnisifsvMd
PrlQ9FCq75XCD6pZVUyRVkaG8yMNo498zr4UZTxAGnZdg2xvSf1Mk4mCccYjtlOX
rOOvmEQTYWY1gELoO4MGCJvQH+e+QnudahjaPjlvHqg06jBpl57X6UbPKyOoL1WF
Hz+1J8jr7dcWLZitHLq3BAKsaIG0gax+vWRQFowi5iwhSo3GPvDnwMidiA/usb2E
tRVrRQGcTENgqhFa0Mq87dlkAvaEqBr/ERHelI83HLYsXMtRjNpkKbV+QIz3qaNy
sqx92hky7S/1HtLqejoO3f9RtzzOXnnZ2S7KKAtcuRnJIsCuuPnYfKNMX/9mMIv8
odbussc0u84L0t7rGJZh0M9MUWA/+ayeoBXo/N5hP1KOPeO78HjoObqzWwYfIVEs
pbUFa9MQ26+t645wQlg+ZpmVFtdr96/32YvlCqjhuLBUHCfUF5Fr+0HI6IxrknRf
b3IzkqdWa8/3azsYgf8Ay+u5VZH8OPWLLUBdYhnZBdHa+4B4g0966FSfI12O37Ke
eY5c9cQr8eKIeIp+RLIVf6aSoGchyy/9mmKJVUmCKs22tOeRZ49po22bARfvrSJG
AVB50uHJRvEuDBX5R00IBIhBekQ5MxeIdhhZMynOqsLmZCnaAb72d9iCfo0ySlsU
HUCS89r9I4t/+qgHmlLc9AmO3qXVUh22qyTH3mdnRpuzPnr6dANlDx816imBo1nw
gnlFfsRR7PKkbA7Pz+rfJinvxx5WXW/dyCldPR3zTVfEDWjdbaEuNw1zDdVlNqnK
5ikDDucWQefF11mg9pjK0UGsc8d2Yxz1ALIzm/a1N+4x4jO0mA6HqV7ecELQlJx+
tahqWjYVce4P4905tmbhYcsBCbLOf7VouBfbujGZJ7IvQxQcockcMTQALUlEXlnX
XmaziP9QHgLnlgeVYoq9Ql/tNI+XW9BPYdtg0cpVCurXiAvoX0//qSppjsvTbQRA
TcoTNjOsMRCsB46/yDmE/nkk4ZEQQ4RPvUfEAqTDzr05FjJs8IAQKLmwYlr3779Q
UNHcYRexswB3ZC/dLagiVSRI366ZbxM9tbcKQmxZPD2sWyZNzNDo7Shw85nIdrXe
mKKr+kWqs5wxbTcSP8BNei+VENpoLJltqwmEyULGn5iwDvoSgwm6pOc8VwgarS6q
CU1jmaBT+fE1sRcpvjESOy0R9E4mmkr2vz050dQR4geOnrrq79RFF8QJaPuVOiqN
mIFBxYw1rpSNCIQtBmt6STNZkFaLyi84jRK5E7jWagptdblWI6i9F//2fND7xqH9
/A+tkEmFHpumqFSOHnPuwegpzIP2aOxoF4Mp3hrOkNyzyLDJbbp1dgL4gaOsL5hJ
dfBwTnnq1neNoj+J7HkNec5YhooUKe/o2qVckJgApt8tpnyTVacW9FQ2PvqSWAx9
OZeXZNHzBuRFIHi+OGe9kHyR9IAkaPADDk1qvZSBwnRxEI6rN86NK8MIUlOFXjWK
OWBeHR9PPYHwiIyZ4MMdbk6G0U8YIJlReGJXKqvFq2NqiPq+dCt1/hanDiUis7Fy
+A0P4TV7AzVGyGBiMcoTSIU+MiZ4UjkSDEE8kxvjPevXff3F1rRTu46GuyJvh8oE
rMBoBRyVIzxjJwRbmPTwRnbq0VcIO0W/S6NrD/XSIbFDXAU8zYhlwJYIg9CyXH6y
qiM3ih023wIAZgu9pSR0zrERezLzlvogi/zH9Xxb3ku/qu7sVbrVR6TNwIkZH3EM
1rhLKwjUhDJOdu3bMTMEAoZA2ZYCZXix1EWqEN2toqcOZ5UUg1s1e1ULnny4RSBY
XYGdl0EmOsQnE5haBfKBBmyBHc1EKGh1UAMbT3Nv1ZYRSvV1BeVjhpjD7FaKQjOA
pMnU56GNCG0ILvXRE48f/BlPYQckgOIwB0BJTG/fKGtbrAE+NKHuRio0BLNHBhtI
rLphzQ5HnJO7L0YNdVe67OwbPD3ZpG1bV3z7Zbqc1bPAIJPtxvZxKwFPCfbiAcaC
Os1qrMTeUfCEg6MQeMhXQn2Ia0xQejHoFX6FuKS4Ez3BBtpDYtQ0C+Ma0/lHZQVQ
Xd9/8aofz24LHWaSdZEiVkS5eXwZUcYi+iuztrdcjdj0PvmMb2y3iBHTLegFOuGv
ypYABb4mfjs6rmXKi8I6mSUaMFkPp4LYFW6Cz31uwLLEkEmnBise7lAzPb0f5/5F
ldg8E6wN5FVAG6GDQ3R5FEG3EunjkBg+s2qKgQ4pThA2+Tn9UBfgC50NKqyK1JU+
7aTz3swUYnYkDL2LEp6gLqcvoi5zFAJx/yUK3drS9yVjtHGjHdUcz/eXT5nZ3pag
602FeSLjfvwV+/yvp04+7FCzAchsFWUR6jqFPjRY8qEAyOfFsZDSj8UTff03NEPx
747wMfFEKogpQoZKEICEci/zcH85lJ7jGbfT7nCkOt7xVa4GYDEh3OEMmKPO5Zx3
oUyhxCBPgqRAXqTA64l7TdEDqAFx3+QLgEck3lzGrergfZ+665XyPc2NqqKLeooK
W9M/yHNaRDIkavKLegsC+k/frzxXIzE+6yoTsgyVK8p9JaC2pfYpkiDyusf/hAZe
mo3mjWqZcHBfUjK0MfKsOcYdM9FQEaZk1zRBXdTrshsOjOAftpldGCufY9+YE2Ex
TxwIwnxHggPzMoceFPsZrtc/5id2RJeO8ZQxVhKzvWgMtzoMqz/n6Gui6G9/Kxgo
OwDVXQGQI5YfF2oWEQKNF2OXfnnDzIW6BE4p1vXIEB+JnVCWyLp3cc/rkxwGNE5F
SK7omhhZvVZ1iikNIaAMvHuk9iu11Z96SyneFkwO68CSJ0BSas5dXoaar1PXwOgC
G6Di1cWZv42jqECWgW7rErVdzCCOW90j3Rab82e/WcAob2GM2d8PxeA3Lgzqsles
EIh+WloDvpx2Qfx+JP8CT4v0k16hVRev9/6NOWOkyFh4qkLNrREWiL3zeXfx+q0k
7EdfDFX24yI+LQAVMvHvXLgtce1ng9k2acRCIb4+E/Sf3vcoUxh9HQ7rbLPOrWM3
wduT4ZzFoTfcLq3ZpOqkSX9IFZaaR/YKKdLoxZDlXJBPLIbWz7MZiieqKxGnxQjO
TeqbFUh1mYH+mvIPHZwsLHGc3sk6X/KujpwqxDo1lmlDGmkqUlhw0dPAjOidG15S
iYqq2Xo8YE1rsBWQ8pUReAS7CxXEubHGveZEvAcWBR+oNICYw5hrdK9L113oBTVQ
P8bF90bvjDpFrPDs/tsjLY9fs87ASNb5hwfnSuVoAwgV/O2ru/J4rypMb3ZRYmX0
gGDTCETC5SC2uBywAHgiHTpgbb7bgKRGl6eUuqnQioySK4mAOEVrDRG7ZUzKVJta
tocKyrxd5kUFqzPyFkU7IA1E5Muk9deNMnmFlKvA45rI+jZCM8OsQu9SyVSno0H8
XHppj1NAzmAJhN1g/WBglsQVQFy+00omyqomZ48B7gOMiJrLcPeRpGgkpYZsLzFX
4yDSo1DFKNJrB7p6DgDUoFefHBSks6M53DG7d2eW2k9DrhKsTqdXTDvIVWAGoB5L
FREzk8k3fA1/2FjHK+1e2iCkY8jjBxsJ+sNCu3v4TEAvOFoYDgPk2cazOr4+NaKv
SSIvvHrVjYKj8Kiitc+RqtHb5Zl8a4Ve348ruEiVhcRXrOnLNGYjq79O/4cP84vP
9xPZjAfxAhRs09qePA3RKp92wiooHbqb8H9NG3KbK9xa6u/hzkeOahcSylruhqC1
vKajit0D9y16vDL/iHgnXaBSUscyr8XdXvBLjerU1/uHc7+HlUzBW5PNkK8QpSXa
u6vu++iPWdHu6HQSV6tP/rDLVTvB7MrO0afoxVOuKdW/GcodprpEhhm35q6ZLlF5
waRV09mfyqSvtjF/F0U1bUyjgZVDekmFYQIUTH9jtHWfdh5uj5PpFqTLxKlI4r92
87asmY935U29XpGUZeJpQOXc56+sJyLBQKuTA/j7ZtNlYIH/duE1Tt8UKaeGT96i
y2QFC9890l1v5TZFbjRshor2lNKoD9dtRmNY4p88mV5GW1CgDu/K2SfblFNTd5V9
oXbiURjJJQIRMv+UhEsgO+Xt93GxUT9lW4bhcRM9wmGxZ2D6LwGaZAg9E9jg3k//
f8ckRCtnDZZWyNxW+VuaFYPMOw7kFyOhLsUB5NGrdFLbtghN7DZsjBso2Igjp8SK
UJcbASXfnbdg7d6MtmPr5vqNyjAjEWMjm4KTdvJJSzSeSy26H2YO3oJ3oeg8fsoa
IIuIt6/lt1bsYiH1aIzLLOiJg7w6zJuKSSDgb5pt5CRdD0A6XJvEdqvhNtMa/0co
3F3VEyTw277heBH1Bljd2UvgLym/F2QiwGgnfxkqCSfyboQKFScWgRfvG+p4yaL+
LXcm4EHOAot5MfBd+eNHqjCQVdsJu2Pg7E+NF4bt0vOkN1ayzrCA0jObKePAm9Im
O3hJNd/+thDSDJarPVT8U6ZYoWMY5ZDRzoCHb2cpz2oTxv4pF7TQCoZ7sdQy3/aM
P0Nloa3FbLFDZ++dhW4hIEN7FnS8R7fZS+0qqxUkSq99B0d8fDvWRJF5ysXlHfuM
t2DG/B1ttH6SOkJwku4RkCda0hlnUpsDkeEdZf1LBKBzrnkwGBOBhhN9feDw4lc0
nxLZvil1mbApWNrM103wHKYzjiqaQdo4039vOPwxHPOCrD4WpVPHI6z7EjHTwhI8
/v4dGREWwU/8YXgb80qo7h7zO5C5ADLeBVpi1mzn8GttS8INF9N6q5RSHllzraky
qaPRul+YUfezXUAAl3dZwcSgkAqsWsvGe2rclXVJwEi7V0twqYJEQadQ2nh0Oyxd
yoEiFPNefxbiIrv4lPUrbLo+JS5D118s+4QK/XlsYhCS6os4u0B7n7C9qdlbb41f
dDDL6goR01DJjwXT9PSQ+RziF/y70iX12dScag/hHu6V95+4+EggYFkhHrMVbs+I
7CA3w85fAXnrBwta2XpcFNFYsfDlVzdk2s0quX7r5V0eHj2W2jIsjfUO77uEy8PZ
3rX7ZP/cUjkz9m0GN2uPQ7kfAsGkNnKlhMjNdX0r7lsvXtV4j/UKxGv6OsBqeRGh
YoBQ4a2UKJK87y129eIsZBV6bV+a3Exu/Vkn1Fu4oxiibNToayXZdPlwfVvJsdDD
3o3ZbUzoW3vn5HsYee2lDgU+el93da7FVJa8GbDlts/uMoCN7PhTpU1eMeTCuL3W
G7jRZPxaEeiAlExtdhaYh3dNTs7zF3c/3AeR+2uAHtnJEUamZIUWwo5n0LwIv0lT
e4E3jd51ztyYW+7OZxP51jHHKLJoIBIaKKrkljaixBCyApb60MSVRe/usAOlwRXn
ktPrq5BsKG0azEgCw9fRkp7ZvJC/udhu53GtuCUYZX3HnB850GCUn3arXBnoiSQb
BFTaE4Te6wXSjW8Da4Y6CWP5hWlfRZi7g1hSVrvvILoY9Js1pZ5j+Y43LedFOfwy
xPRtT9TvMD78qjxogI7ZDcaJL1dEyKo9HwZC0aYLaX/KA6AO9c2BI+p554eD8FiC
7obOTsL70U1KRXQXYMLDAimcgH27evLa/bsFplrpl613uiRQHHQt+z0wMM63H3bo
Mqc1lY5pXqZ3fxJxuqGgn3M+fKox5dtJkULsva5/+s0dtpr/kIK+LUr6BoraMgux
DbGtpN+B+9RAZ8llVLT15aGt49DXL74dgKnXNp+1HfIkS10/UXw92Okyf0/YlYM/
rdLKqDtodjxy/pF1+RH5BuZV94PoOlDb5oI7iJg+4CB9ztYH8461H+T6QvgNsM6b
BVYaosDtRcu6eZnuVUach+iY7qcw/10rzvNXBc0l3ibVHk3oNBAdPrhG+zZzPEJ1
jyROwU+u0tQycMuH1z63gf7ZXi7O2pkTYy9GOTWocI4Z7+SsshKHFJ69fE8Va/Gi
dJw9yPMXbc4C6YngstGFfPOFV+oe8YFXkxng50FK2IFrTt3dr0BydicweIo5odmO
yAsPu7UjQ8miv3HNO0OrYTkT7pHfdTLh4WTj9ewWVAx4DrzDsBVFlx/4W473e/iY
qQCTG8SfBWazFv2TD9sIm/yXDuTRi7feyNTzOgiOL22w8X8VutRPzAPhEzC+y5i4
dKPIkzeCcUK8z5KlXbaSxMUGy5MYWpE7nznqZ850zViPV5UDZBBYomKYB4wO9zzk
wtyglTAF6vHntZbCvq3TYMVmk4ORM+AE/0xJzrqZyTyfpDZddfM1ctEdaQNmnPnp
3tDXVDJgY+k4HKAxjyyCd4eoLk3TzYJo6wAJK/8Bv0QTFaR9ZmWZJyz8uMLDlMWN
46+xRP+1ebZ9n5V0C9rFeeJjaRn11OrC05OTEtd12cGGVCo+GvNOatxgs+iLkgQa
9sXsE9QCPLtYqmnQ/23VPP/QEWyLtUj8tRnDJPnGtbVtdeOTAmXxjG4H991hg5B2
KrInlrPtO4Q4SjEj7qAPvs3ST3tNuOcbrW80mVfTjk4wy1wuLvcSC3gD081BSjr0
6GFMu2GOfQmYt4+lYMJQGaSjglwk8tE/Ayn/yzg8wF/SsBrsqsJ/mBXj6Ysb5F1N
suaIVoycXegudDabTmsBsBPkRN+tBI9BF0Zk2aULxcWZCkciXEC4Wp2XTEjPmV5x
uuk3+hOzFUscQbFXjV53MlCg2zNgCjLmhLxhGW4Ii7pBJg5mP81hsvq8PPac9qfF
2YBhJNi2ivO/1q3E7jnmqhTXdxtxJ8ZiDwkOrhxQKbNZz00VZzkG4qDLfsieqq2P
J5s1tJ6bQJH5wvXXzfiPg6s0qz6ky2xL0MaJszOoSIzoADid51wVxVK6ZlGDRbbA
ywh5R14RdK44YW6ZEi4ROuaS6lOt9FOv26fBF0mBpzeNklAw1h0brE68sf1zCABC
0v5FPxF2f3ClRm3zVP53qipKoL30Ox7tERjRnd5EeSnvurbU5+RvQfY/Xl77sgOb
hSs/qDT9KmDa2BZqnI5Iag+z3YdY0a/s9jWAmRSJywvbgjFF7GC1SKHuGGpynyT7
JzYRQzJxEOAkpzJXOXF8tqSb2KRVtxNmRUl4AR0ByjMHsPMoV3bytqF0uLL7EUwm
BGDR712m8rQpHMrhC7VDSnbEoAp+a9Lxr5QFwkdXMzh1R753gL985c/PT4N4zCzm
vOA3sdfQozzqewdWof6+Sj8Xdmpe/9Ifko7Uvlj8MWLe2JJXAkVBhLJY1+0PU3SU
RXcdj0kdgqrtC5gwVPUB49zR5ctDxRxdPSyefgF2+NsR5PONyPUoUG3gFMkj7B9V
01vCLYg9a3z22qENRM1Hbdt5yXL1EWI+iUq2arVrQHP7qMdWxhOuDR3r83jdmW6U
JZ1FBsgriFNWtToHQWVkNsajY7w7Sn/5aI3DP1umbpPCoaNNsWHxxWT4MPkBmQfh
aTweQy2YPho/qI6q590l5gb18rDKXbXgIEEuQ8bXG3xdKZmWdzsFXRA7XL01AjSY
xTeUTHb/aTPYnveKWQElsa/YmesQu1Ie7UqepOqW6VD+3LpZGL45d7p3M4nB+2zs
8oosY8PAvKqFHgwsLDtNzg2n/821p+tWiy0PCNJMvkukjlhqCQsHsP9gKr9RWSf8
am38r97Yw2ZMRfsnXoCmuAaJsVh0JXzbnPX1rSgaU5WVP+dD4wEC2W8eTXgadOIs
3l9iI/4kDTRyDrrcgiJRiw73S/vV83kMAR9n5aJBlteXKZ9z4KzoeTNT34VjXR0l
Dv2k5PmVqCDY/RuTO0wurp9cfOOOj86uDmdYMnzRl+y4ABPRsJa5BVvmtAJQE3hn
FNpShQkfH69j4AYwgjna/T7y6NbskEHOL/g8MW8to06G6IvwoLWL7VqZDUctVZUi
u21npAYUGxPw+LSfp4ViTeOZ7KcRZtwqOSQsHT6Dyg/9K3qepYZrfXDWAthisRL9
WWfeoK/g7OfU/lCIxEQyEjwHbg5f8pS6IZGqpjw/DcHtx+Vb9F0QSVJd6mj8ZekB
gn2Ty6tutamkt9Xp1wmUlCDGSu5Z46RBQz5slswc9TCw/zpBfIWe+yLPwC94ZKRg
S2hJETtEm1G2Oze4AvbyVK8FS9gS5yTn2CDjLoRchIvRQJ1cjmSobcILqpL+8luF
odnTCNv+dwOHGHqrlDqSdQpERDalQnhKQtmvqKoyk8fMn4JOrG79G+Zh/rwQM808
yLdxxq/OR5DLnkwmp2aPA2a6ckbp1UEwQ/O75mxQsCnprPsLlwc8BJfXvC4M1Xqe
/2LahY/yKbBxhrSpdHxcaT942u/N8E/h39VIcKmxtiM1eYuo1kbQmEiJkRyNdo+e
eCWJg6HbFNZHT+Lt3U3akLLQ4fFP5U3UDuZfwz7wrgNAghD1NMZI41FujA0p5dCE
t9CtZmdI1SRDiI9lqwlJalAhXXf+Tzy1UJr14HXJCD2M29dnCn7n1eaXuyr8eO0p
aaTzq7j61F3wqQDTwyeQo29qoAYg0JwhGpVOvQ0uIHkKMgoaaqp0D+Aw2621GKyp
w9A+KjqFUgjt+LU80WHvSvxeKisNbmYYZjUK+pcDQ+jl31E5dfks3JKqy03iM645
lcrenRvD8pySQP4vZOnGN/3OePXGXjSluBgg43C6jOON954CCkS9SCPL6tJSjhxi
zGgdRmze9gz2qvSwNSSg+H4k/D724ULCc1smNwOblJkWK2b6BK5640Igia+FW54r
iL7XdlYYzkFUbJllgglKAezCDvOiEfbxsBI77fjlhmLs9kzpK9QwEC3+IVH7zWTT
TucntIRE9dm1pKswVaqQUNnUymsgxFWP/54hUBCYgq0vbsLBsF+EfyXeuWSec3eP
quP0pV34mWL6ekhH60K9YkyGjqCUjBYlRf+Hgmr4gZfr7AJ6AVIg/eFy09lzM4of
9d1VwrCp7FyqWSVDXct4hvEUQ+BnpDlZaROVJ6biJh2KLedRDCWhjg063FATcPKq
OZduA/RATKf+nMPt6sOAZ625+sMYiqR91Gdrau626Bak06f88vujRTzi5Leh1DB1
cPCxFUPycr0UiOHeo495QYOZ+CfBp6VMFYQIJZR/ysZV/Goz9I3HxW2f8+PILAgQ
D0OICy9z0fnYIzuPot+I7Mwyw5rqfUb89KX5v8Kzxj3XVfx4NktbPNbmq4yX6RMV
jCDeqrdyTfBdJepjPLoY/87aHXl3Sq2GjA4tF5TuxeF8tkaP+D05i1Ktr/JD8fhT
GC4t4ep9fA0sPU733T80zwk3ySjjc6GocuDaCjDCXBbZs+TfFlbd8TG4kG4IRTvf
uRpbgIN4c4dgSAJv2113GOOHaOpmjBklilGXs3knlPyqF8VWFiXs6Pj47j8MneDD
lQVSm+uWoR/JLQb7Kz/OJ+pfNp/FjCVYBHsRuw/29gmdL5ZJXz2pxkS3NwOB7VV3
ESGqA9PSwdJJL89DaO39ARn/39ayoXsUGQgyVExnS0gBUtfMnO5RUMJ6QxvLCrlw
cO3O5zc8XMFtXrMB1tOW1JDWZI/oIF97eBU9tNEEefKnmGi8QgVOgbUzWmOMRbhV
2cDtY6QMpWqlXw8y8jiC9Oy1kbWOMSa8KPnLXOG09Jm0ctyUYJbxiEht2tRQZ7np
LBGT+YKdMX5nxRGDjYreHUVb1WNfmDinE1565nDtvPz680B2uUJZDs+W2UAP+LKU
7ZS4YBr/2+pMPncIpKsUVL4VPHuffGzOKx2Wior/7OnYi/H0l5vctuNFMU6QbhUY
3guFP2qU9ebazauCgXo8YGfVuUycp9a4M/f9KMtjArXCaEYuyHqrZUUeh6mXedlJ
CygWue4/GRP3QAUWM9dZnS1GLsYajAlEupl5yde4OFooAJWSU49/HMsWWf8w+CqV
hrlpIrVmMvnLpCRzVwSItTReQaIN5wsLmuUvlYbHVo0jsCgbhoZU+QCJiwnahnQG
5ZZGS3wI6p/D3xnlnSQMZrd/Bu87v//ezVriFBpu23KmXXzhQHFrDs+XbX2dTDk9
4mkktBqsirux6uN6Nj84LlQgwKMH+ry0qMDnZ/19MCGW3rz7Y7JHqp8bXO30jSC5
Lw5O4LOsi3YYj9jbRAQ+X6WA1wC1r1BSYN5WfTQn4fQ6ggjkPDby9uq/toI2v8qk
jckqcbaXrPKNWt2mixKqvGq2v76tmL6Z+TKSu2YqjmvqzIMsKp7jNs2/xhfy5Cx7
L26e71tcWYO241AkzMG/InOllB3UVsNwtQMu+DBTOFZQ1lPz0B9DZFbnuNRa4P4H
iSC0pSdL/wXoRoo5ezZJln9agEUxSp8eBzugVC6hts3w8rVGH5JndJbxUYMxjQu1
ysWf6qv+1e2PDkkOE/m9gGCgmTqFrrSx21yD3M1J4dcGlkHCYf9TpAV6ltGkE/En
T6zjyESBIZfvAA8TZgK2Wb6J1qityDIKXoTICfrrTdR7VNsRugPgg/VWufag6f+4
J+A3aOywyaiQY7v+vyaTqcsWEzvk+D4EgS7VKAdpkmcZef3QDb8FmAXUFahVkEhi
oSf4t5gqifKjX0qELs33VWFTJ9bmkWgV2+Uj8Imzk6txBYs6BhpODTkvyQyhPCQD
q2sIlMfXAs0z1tsljf5hwccLWb9ZGgqiBMP/hdNMrJzM30HM3EIpVkvB4VHCG3gn
T1Nh1r1760syVmR6/Q8K74tTrt9sLe3JrGNqeDugA8KPcvuWNeolhuWrF29uP5V+
zw3dkiSPLIptfx9ceUnGHT4ag+24bq2ymPNr+pIln1SuswPtIcn2f538+PJN/Y1r
0z5pA/AzIlb0c+ZrGF4C6zYRWIJpwmOYldLl+vx9+vlY1s4OYrx4A30U6wmI7D6v
tTWL8dwSk3F4KW11fxHzyyDKg+/MBKE+k41kbJcl6tt/GAIex45bnhvx+p0zDZFA
Cj3Zyc8plwklFSHVUYlSuLFTFRojiLSF+aCt+IP4AqnHrtoM33qm3GDapX6XaM8G
auRJyxshtHunN2xeE66n3ox907EIgjR7H5orHykdb2pZw+8giqGEgme0prJ506eT
npwMhQW6J6qSMSc8xWdkpm0eIZL7a4LYeAdaW/Srux6xZ495Zg/JvzfWWOQysg/r
Caxp7pPpkj2gYIEn0ep4Ks880aFN3rU0VNCq1wwlzzuhgkchHVZ0AtYWTzHcbsLP
X069ygXjDEFq3RiuwKoJoj5w9mkUrS3Tsg08s1ZpEIW5Fbk29634ms1OcNcafnY6
KjBa7XWZ9NuQdnXUgd2Qn90MAHImoxDmHawWwV+0qhkLvuZy/2v7NtMjPsNQ2u8g
d6RhvaAgrn/nRQMzLK6cBjDewbRGh7oSmzoDocszY2n6FIU9ab2otISvm9henrws
HbloAXvi3gwaH3J7gG4up+Gz2BbpKttNAYMcmomwkpFfWDvNSxM/5aT8PaIdmcC5
BfNkWzfdZjEE7XXlIip+fVtUZKk9EdWXV37gQN/UHNc0qhvSIITDqpRhgLHDDICX
HN8hm/jrJtXKA1y+kq4LnU9aUfE/GesnmVp6C46oByCfbLePbFQiubIZrodgM0bw
dfIwf0kFQPnnk7ebuUdCofm0K/gliNvSmMfJKTamoYA72j1vW5z0oo7KtM+OCvP6
jO/YYsuX3tv8aD8KOYOwM+SILy64TwOHX40cIkn7rmlP6NCGGifBZi5wemBVON1Q
HKLG+ii/760+OS7Iv+1akK+D7sS0V4GrluBOR3ts6qKVYYBFCg7BDDDt6cSHWTmF
d72stNAmGwd9HA5BHi2dxT4nndtLFNwYba/Pr5p9QTlbBwW0oR0tQlWija4vygFx
CVTEpONWa4+23n49j8FsFd5qNSblGn+v8z8gB9OLqpy4jIqRkvULpA5444gdKFKn
MhikY9QDaGjH38jt9vWyxm6F0HCZdbS8se2rG+cSQcbShsG906GZERzWD4AQn6+S
PAqlZ2rfY6dVcFgxtCOHZxrNm0+22FGGHK5O7p7RqvoZUd+UFsx/PJI/lFtF3uxs
Wxtk8F1JKuJgLSFcXBkRfmCLjB4ZIG0TM06Zz62FArTPA6TvIH9/HgoSM2tMH3Vp
RXbKA4yv5DjRGEx2+q8Hmefzqm0zcQdwIA7/HT6YMk8rs1nC1eJdFwWrYjmabd7u
QLiKzgh/OaPeZOQxUKv8ULJdgFVUnruqH1bsifLK6eUP4y/eJzMXzFBtdjB6ik/a
i4Gr/RquLq13qDBmj5Z2KxgLEfvUg5zcL/azSsYCmO5aA90Mzsii7VgG6gpWR2sX
tUGf4uHqhkNelXBPeZJnhR7EUjpNmcoarlA7ut727JJqnVrNT2sa8wnubdKzjojI
rwgBb+Afc/U9HHLieljFmY9GSxOrv/6D3+BLPttnFrogIyAykGsoGUpdVeOFNEza
VV2BxKJewOlAw75fd0T7cVkcZzO3JED/m5gHT66LOHaDJbCP4EsFu4hk2cNFTKxh
ALSkBsU44msXO7Spa1KP+AttpqWaSFfTApk4S4/aEKSaKZUx9TuLqzlzYwr/CyUH
792KJeG2AZYUn1WKaBVTCI6XsG2ciHggRgJcLJFD+5l1JMQ/Xal2SaSisbO1O4P4
c9qSnd72MLAJoryoouZydy3eKYhdxlqStLqAwFBY8QSvfKTE27hE/V6geC6+3omW
C7orlTacGxCQNk54uXlgIAbH1klnsXOiS9XTVSQ/jGOPLYQF2PF41BMs4JO+gyMC
neyXbqRsT26NBBo2VUEXS4fPmhf+6PlyP2UVoVDcOaAKqIoZglYkGNc6VSpoE8e8
o3jlN0CTKolkPJ+GPd/bfWz1zQ9gMJ/h4clgCCsdJMM9bBxAcV29vX8JXozF1SRI
/xrVMiuM/hqnM0svP4ar/v55Pw1ISdGLhZPH0j0Eax7Bu4lKy1KJonZ/ZEr9UCEG
5IxllD3jodqgbBCYzN3U/DV5rnGzlLC+FbbzrfmFhZUPZgPOuKYhLEiwIjOkQlMO
urXFtPL/+kiAEcxHFaYUoNHCXNu7++qIPF6uhTsR32V2DqqUICrRlhZE8DED0t9S
VBqCJQiJRA7RXIhcOd+GlCnBjr0oDieRBrkUJ8jCvs/1F8GKDhv5KQ90qC8I2gUe
vjYrvhLDhwN/w6AgJSx7B01OZuRM2eAXaR2qKM9OZzJgYqIh2QqT0IsgnxAgBkQV
AB4sxodgdwph1t3RtOX7Zn8wGzaGDm3/QMDV+8/LXvHofMBZswU45Z1g+RPlv97H
K+SIWBZbAxf33o5evSPncuQN6XDLRHaMWJPwZQIwVJQSxuDW4AVGaFl7DNBxAltV
iV+pz9pXj0pMJqtant3pwkAEdmtqR4WjXl6/jJXkbxUy0Q0wxsoqVBmgj5720Yc5
so4dGrJXc5TH4lBsITspkyeoRPQXr1tr3iq1U6goKZ+dQMwSIU2jIg73aWEJ9iyt
ZJiYe7XGAMjK4qWIrzT2xrTgmEs0pJ034wBUNM7xYr4i0JYo+iYITBXG1frrNrqW
1V5GDayEEgUjxsNFa37aoIUJO81M5RJUPTicqGlhXm5XXq+agu8coMiueB6KZlhI
r69Wia0qJOcGcZ6AGWJ+e0BzD6lnNiaRPuYRFFa7csZnD7f6cbAjPiwHQjT8BZkL
LrM459cFXV3GIGgmRFUizTI11kFbwbFsGMeMstBUlbpIAvZTQ8J0x8ABMbzAmswp
n/BUkrrm86GGgE6XkUo5tCF8gWXX9zWtGPFVspT2YMZU9FPd0OkNQ7iwsuyBJyWh
144Ps6e0prq/bdB93eX4egff8K6VdASYMQT1SUn50W9T8ZcYzFxQIhvHFBGVkL1K
tR61aXUCtud5er/gPcwh92OwdYvgzZmuG2/xio54+4yxMJa8lX4Wu5taD2qlFfrF
OYxekbRq5WTQq9CM0VfIJ5eRIke8/CGwwrxyCZkZmxzNHLJOLMuO27SHkXSZJgST
W96QE4RbtZywOzkMhejgBCCWyUHABhPeCb3X08DS9oV0kD1e5V/6NlnWHyuX8XSY
fzRa0xat/8rSSPqxT8Gt5LeUE5s+/WRryvu9OkJpfqfU+Nf4VX4vR5hsAWWPN+ti
Gt622Wp7397SDw4/ajM2Cd6RD7aZqj3yvCGeFZKraIAwcRUsRrFY2df3lf6PfhWL
WhxPuYSxyG6dTjh7Fquqv4prfx2R0wHPYmeuPQqw7eOLwedEOrn5GkHhUYyjM/BL
9+cMx6QaZVk5SIVDBqlumc0EU0UEqR5Q1OSb3n/OpziSItajqlTDO8ZsvZld/rln
h8LcTaLDfjp0Aw9PImZtRMVOs3AN+C3p4z+n2Zv7A+xbXs+8R24WQ20BIoeZ+RCf
jJsWhuIPqlex6NmYHgzjcHhg08BM9m8oZigPP6Dra2P4c7nqvOLwcECaZxFFFvfS
94LlSk7zwIeNl82UykTcgb3PgxMxK5EORmVVZ9+RkP0Nhudhl4+KwJMZYeMfMCET
FdT9VWp9emZgSj0eYjXbWOJRRn3gqiYMZI3BTDXDd230r4njoBrYNAgUH/zaSTew
ZeHs7johHrYTnPYIAVWlpeqAHCMemfVXYsgxTyJFF0SJfUAaX+F92bIAkd0bJQTK
BbPM6Q1dQTkUbagmM2fIlPAC00+PiqhZ9ShSC3Yahg8UUvc+zoSjGXHlFzo2Dfbh
Itwx+nsjGsT+4T51kPObZQ20kIy6lxC8QRD/j8Yy28NL4Qk5QIOi3ctV0oPSE0Wo
i5Kd/NT4bDHxl+S512q7P+fuwhH4y+hDTu17cEvNdCEYxZZnGpDEmqVPGkjOnulC
4L6Dylc+Y8VK1YGmRcZh2SQ/gPaZzu7iYdRu61/stkwRH/ugTo9FL4w3X+Fn0AYL
VUmv7MsYwdCYxWLFupIr4hhYoKGCEkvlUZidvrke8TLwMaNZUmW4Fpct6G+swx/P
0lkLPCfHb/9hBK1y+FH/OOR87fiZGEYMLDAMegX585TcWJwsMfIGzzzoF1Z3VPOu
wmbEJsHUFErTYcCRw4gCpAetO3NwYNcbercK0kxezkZKzgMxCOi8c3HSp7hSC6B7
29QAGK5I5260/dSp4HggBHZJ9QuKu4iHlJZn3D5bpQBgttQGzlCxXUJInA+/nhIf
fBUoaewcy6Bqua+MUvpimhnvDHZaZ20PYBCnJR2yQiw5rbdanj8/OYQbEuTWYAy8
huh69/CHYj7ue4g3AmMrYx97pTOb4v4yUmo8cj4Bw7VL3AU8a4fdFXkGZ6dCh7hL
koyUxlIvBWxkoO5HFvkWk1sFDK+xbwYN8wcn2G+jKyGjju24IxGcJdme2Z7KDQ31
agO8Bu59Id5VO1n/4A2I/RGsrn2uXV73aVZ0Rc32Djs/RuZsEWQSrusdrorxkcFq
NMwiAm/FPfDjHZ8P1nBcjMGmBu0xAFuHrunXCD7baNZH5y5cgh1AuyM90QB8CbZH
kxwlSbFs+AbOOMDK4vxrk3GwhRxTcYwENRi6JJ4WJ7gVXESR0HShPO9gz0sNm4J2
L2hdu9aP+uSjtgsruM3A6W4yx9Wk3vK+6Gw3+O84LgbLuL/Mu2XUs51F/FSjKs3r
E3uqlPHQfzOSWIPVg7BU78jJrmYMpedot6M+cgH66hKN6Rr650x6yelcfOTgjkRW
rS29NLHDiTBETnBLsCjcuXEcATsUl5/Etb21cq9YzFN5F/kxGGiCMEUzwari0b0U
oT+xYPtS+7kn5CyxZdwWUOF8ex4wfAjqik6Vlt7oyieb+pCMdDVCxAskRhx5iCEB
SEQZ0hjhA2iMBvohe7VSPc/+kpY6gf7u1ZZuBoVvg7risOknq3VO+fOMEXvu6JkD
XBDZdQLj63lLfRhoa+IGRHA7e2FeW02TNcqeTM5l6ArWnrL7fFyD/9IC7L3etXOu
9wn9UlNoQWGlVRUNIWow72QCaZRsXOhsRqCeQnCuzPoZQlbiUWr6Dv44ovrX1JwJ
hUhd0PsvTMAk8WMKAyYGwzocOOT6PHZkbT0luz1O9dzh/D4xCqohfTbC8jytEalE
myzwpvEMrwbkL3dmlGPhx2G6D3n3dIw3qonmQ9U17KAiv/14mZi1TwGAeC/1/WT3
8ClyDcAMoV8aqm3V1QfXW3Ol6Z8F1ASjjKo5iWyq0QgqAFbLhq0Wbzx22DIiVs/Z
Jpv+eP4TQkS3bAEaBTD3s+eWQJsAL5dnZhmWeuP2w7uB811O1zcSTLIpJZHaGigh
56u1JczIbccBm+fEWSJNBoqJuxMibeWaOuPuXIbkEsaUCRBGg8K72cTMxH/d4Vct
lop0QJ16bLbg/PzE1Ns0Ne1QteMB5KsA5H2TiZNckVjkpwFmqLuPML8hwL3RB8wc
irdOjgnsDaafl9g+TL5LyGkqRTu6Yo3cbGAAtWWvaxZGDXzPD+QFOqgi0Pq/jJRw
nTjxYGfRBw7CdypW0GDmsmHTSw3FMoGHuJ/qMiO2AulvcQTF1BKPwOD0cIReXRLg
X/LOgVWnxP5Q9eQemmh1ZuIrqOGz2CPJ2+bnWhAQ6PyGHEOypzZGuNYzVFa/8j3k
YWAmii2m3iM6KdInmpE86tPwKETy4G/pnSRrB2BYGrdOWreIYhCjWvCYtObkAcT1
MsQb5MZEiUzKM+oOPfzw84t4GdI/7auzyAElr4o2H2VW6M9+A129K1+SAkwjPNOI
QrjMgKK/uaKwiw9ydB9IVZ4Xc2nUa4NWWWkOjsR1qRCpJvAbPUOrEePE8HJ8l6rz
TDgtFkBPwrwPVi9mwbtfIHNXPWYK7DgITd7tItyuHrT9lODAESowL8izLZTAnBfS
k6y0SM/6hFtKxWo8LwyCTe5EEySRcVzuIaf0UcrBypsv+3RLtiZ4gKIJTzd2cf6i
4dZ953UDNcycKcN5+vdtLmUNU6GE4Xqmvzm3XBzA5jD3HtEqnYEvtx7BjELNbapm
QkuA3ObwI9FQHsfsrzrlvMdEkqKuL/2MRWqPv6nK8aQq46W1bfRpeK7JVBjr2Bdc
BQ6a9S8Ji7QbzJiNxNHYKa3dTI7jZX4k483xRxFsQPU1l1QCzx6tGOx528Btsqe2
r+SSTBQjGUYMOGS179QbUaWvVykCB9y9pn2RcbctloOjh2luJ4fMliGf8EXEOmn7
riF7ZIf/iwuR+bfyplf2NT+131FNwx4dR/dLZ92fEi+balBkENGi10ScqHVKioDG
Vwwzxd90S9xRWqa5qzLx3vW277mm8jb1pP7bKAXJnlpg6NeFlwph9WxQcboqy7Eo
/xH6mAwf1t6YGh7w6u56OwYDyJJLILNGIBEQ/KxmQwuPWCD94JU9LT3sksWA83WL
s0hxxZiQK1GJwqKZI87w+M5AkUhoOiHoykLGzae/SY3a9UTrT6o3yY3NwSEHgyl+
3voIhPxSUCqDxY1dDAArfSoc6UrVUZk0fUHL4AbIRWEKZGd82sML5N24o2e5y3QL
alDN0SlAtmpfngLBMN1Fjc1LXSX2brpYnFAIyCofBuvbFFczC9FmEShzl4/LX+qE
MDHCUCVolEuTvhUPjcPfex13cvEj1y5Cje90fYDNgaoZCpcKFV1oJkKCNA6JX4J4
RFQSdeJFAKnz+TO3fkIQYLiyr7lkklEDwJKCTTSlWUm2/5uqiXO7CWvABDGqUl3n
3lcU9rhkvHG5SWQJ0mZOUmfBr5cC/a5+DlCQLeWbTwetePteL23IOg95jZubMwVx
w6ooky80Av/06G0d/ZA7vOYemkb5+14qfA2jPwuZc0RwDESIzw5RZ398oyMX0oAt
ayVAVMfswSJq4qAnlPlV1Ev9KtpsSjVbqbWW/P00BvIYUJDp+FCyWyTP+OdkJ7wg
OizfDoR5T8fZgeGszInQvtVcSLI4ADffUFHf267kOb6enpcsMVIJRHSGJrtFEJKu
S7JO03KQdWoagp1TEYHrrOlidxZuG4CMecacQ0HXfKPaVcWHutPvKtRFnNGG8i6E
TMnCvGObK9WVOoy/v234a7lZiPJm9xc1zmVckyf/kYoQZkSECoJ/LGsPSyCuXzzV
kh3grsBJErS8lvmUtUiUlSxSJMOrm4ulOY2WyG0TEJeAYKP4CzxrdfJfm7rMe2PD
gcrKVoJFZm7af4+PQHxxCsKG/h7A2zVMdb74GnAeDyb7eRYW9s9SHNl9txn/78QQ
eGzQpDxKpzD9WvjmdszPac0lA7hqG+GmCvBnjwmjgRHNUHJugv/FZxER8iHMlKKG
W6jcW1lRude3T1Eu6fPxVzrdP7jA9q3x0nbeCz2mNECL8RXZ9stVgPFmrcaqmlAP
nGGO3keZgwDOmxiHOyAD4+TrJDBNhDiaSSsuqQwq0t8FTsH+s4VcY1Lth9a6dS3F
Zx6B436I+8rHEsma9xWCdevG9X2P7Ul9A4muor13d3+tsXdE8SDcL9glpM7cbZv6
MgcJxJwaccu0K5x7dqFJsOGGsBpJPGxBM8ZsohoJZECkz6EEN0nQTcbdLFUZ+oeU
TvPKAtD8eYpSegc+QWR/8InIsmxeG8WTT+Rv0Om2IooW6r3kMmmNq64HrfdHXQoJ
4DMUEn+f/oGJkNlRKr78HyIrHjrGDwcxuovZe0TbqDEWHkS2ACjz6rq6bw8VRT7t
y/co+091hOaf9CGBw1bfsVqR8Ib4MxEM8E4Ibq2G01lZXhZ5LP3gxUgAreKlteHN
h/2vYVqXd+3K2RrZgEGlvC0F2uDbmLvgk/wMyUrKP+IRM5Fd8bQPFEXVuPT6Kozi
8BQGm7aBSba3bchxkaW72+paxM7HcigIFvxQsUw+hxPlU+wZ/o5i69gh8JfBk9Uq
H2O/NpzN582oRrHOT2aWtpdXeL0S+oiJTBpz4I98+N2csohnEzDasxoA2I6rm57/
zby1qdv04L5wAzTkdM2ZlkllLx11HvVGcHCcAktTdYnVsDv9QVpuOxrPKUhaAHaO
f8N2tdktrL7ZvD5+Wbe3LrGj1xzHe6NA90Tc/lQbnfXQEZmXSJCknoTbMa/3vRu0
5pCamoep6IsDidA6loq2AkR6BgTQJsnkMs/4G2i279+MrcwiMs8Qabz8JQKvxI7E
HlYS2eUO2kXtxxzG2eAope4TqK2lKsh4xUP5+Qzej+pvtbDASvUVaZ8p32841613
9EH4CSJkXD9JT/OxzaIz2vR310rROdKFUlhwrifaUo9R6jJozO4Mnt6/Ivojwp4Q
avN2WFCsPkINNo0Fc6y6ru1mzs+860+dPL+Q9r63iDF1tFYP1PD+rHzHhUhhiUNG
z+cxa6MfGRD8/ql6luuzlLN5An0B/Mv40jK5LxErOB1saVcc8x8T6ExQI6Rt51cl
I2CSHF4wdbWovJulXUFPPcVh+9QIlK4sWd14WdMLgzus9fT1cizPYZ+tRdoxQzVY
lZNXB3VREHjZd32Q2upAN+2OR62AdopHJ8Ga05CupjZluI25UslamHHmNqibyPk1
ORRZcKsyu1KGzTMuj1cTodvevtEzZfH7HR0qQbOesEvBH+gV4ZYGwGX163PSF4IG
dA99kNBc8G9KMBdhmXeiugyV8sgbjGz0waG4/SiVfVIroqK3gOKT2RXkN9Nirra1
6+m1kiEXiozRuY/745xBXVV1ThJ3BvEEMc6PzL/qwJydMwAt8sXpYURDUjoWkSyI
9XR8KplXxwV/2Ay9yWdmLX3TcUjhnCFlxqHLANgXe23pdsdru9T1qai1nX5EbrDx
9GVMbtCDPVG3mnZ7wUMoD2xaI7qP1JlAjk/3+Y0xdNtdewWPFP39RdYV5WUUYKD3
6c6nCvH3UYMhSrrCkeDPZ/tDq19IBIbD+b527/yn2NkBGNOL7AZ61qbiYKzOsBQ1
I5imczMwhb1gl0Z8z6ZoFj09XYBCYOuwYAHZxoc/dj+6nFyAKoyGor1+UFM3s7Ub
Xn+5Uiwa9P1H7d6vY74plAeB9VkzIKpWCKFbIdBfCkfiOzjRjrq4+WnRD80CCUXG
erNyajct6RUaBSZs5LLyIdQLLWTqG0vMGyoqtD2TsvqH+JudwWiGQUHuzvhadM8G
v7TmiLyicnMHSpTQl1UUINgWrpH389Sjt1gewFu8Gkeklw33MzKmcDxgC0el2eBW
CwgG9bggxRVbxpUUQ9vw3RWK01ZHtQkNVGhQ23Q1xuN9w+FiEc4QPuSfHkSeLtLB
NctJ8/b07+OjYXEwxxYPZ+Ebv8ziAWLmlFN/4vUaVDhNK1mVc880LWPvh/HscKDb
hWaSbshOkQ4NQP+C64Z73AeeRF06Z3OoQJp5lAXghWNTKkqwZ0tGPps8LQUsmNXj
yGpUObDQH5Qqd9ZXgNaWGpzbVboJlfbJguj1cveT9sad4yTWZPvwFloCR7qHO/6f
tImsy2ZIwu77TgRvIblFdBGsY4e1SHlpsKXxQrXk8TEmVQxM6P5mFa0jxgytpvNe
b8QZiZM/CBmUmvPzl5GOVzY1Y4NQpfBKsCccXjqSM/K5yiUwd0OnTb/lzN5c6y5a
7yraHPZm80kh8hocguGO8XbXOivhDYLiYGVeH+d6FHj4sFjRmLxzPNZJ/eCObC7n
ANeRDR4s2rSs/SPP/cDQC6Lad6R7UGaVrKtNcm3osg9ySPQhsLamLvUHSyppO7J0
qyiUx1zL8DaSsvN5p/VBKTFe0t/eqZF4NPdF1xxMwTyftPu43taGljR8m/XNOXyI
1oYp6EpSoAD4nFISX4G4AFuiQT7EmTXCRYG7raq6hxowkVzA5rkh2tVJKokePr5v
BDAclB3MI4cPmrtwY0TQ8dBp23uxu5A4KXNZAvoFjl5NuYU5jhUxbtfrQsLAOfIP
gRQuwYQsYHB0B8/vsF7nPH16f+/DFg0ovzJ+/nMrYoLL7MH1h9YYBrDCjpaIxx3x
DI9jOzbiv1MI6kcaHdgSWc2q4aqCUEsKCuHUWh/3OwqCiaSD/FgiIqufPuiQ5euG
8Veh+reY+excgXXR5Mk40o5R5Xo8uJ5ERJ8xSd81dKlZ/3TeDCKh6tV75nA30lYZ
gT5WAuaecESLruc25rVEkZzg8Ln9C2wTbvpo5lfiwxxEbFcgRjBEPv+MtEOhtaGV
QBmpEfHFM9VCKH1LmbI11BxkYrmndlO5nEndrdr9Y/zCDNcAA2K7TfsrZxrRmKup
uS0D/2X6YSRG5e/hlVthZYzqmGyqgMJWKZkqkIDydJFSM8/lRrCgem0ZxXozwMpG
/nyLeTXb2DGDKiWKvHN4Zw15wtq1lh4piww+q4KF+vPkOIAJvH72fAzlA+DmNVfZ
nY//w96JK4a4lSHjTClS+0sp5xWPpf5zw1W5PxkzwM4K/sDFfe6oiqteOZXjIZxK
gC7lk+JYJ2Az6ZT+fs1tun5Zr5G8mtUpqgYBN3QB3iLHh3GWK/PCzxMEi+W5PFYZ
yfzzP1pfKQ2rsWEd1dQChmd1Fr6LJfR+DGw7wN5AMjS4BrbLPkBatOnz+L2bHMDj
/PGtUxfnuXRRbL0D1m+fCiKZ70quI3dtGl5zooauup7AvbfQr4wPpyLZGMotQGuX
4dfabyjecSxKgOqb4QcTnqpQ98cqOvTwf+qjlF00VC84UuMHLBWvypEDTazZMSb3
ROVn3t2XtF+nm3ukDCDWeJD4zuMbeJYfPNzqiFPWqe9ks3Qk9D5aN7P1OvIp5a3b
0UwRY61Pvt7U7z5erGPpfapoPaCT9/DNu8YJIzUx5nb7icFcUvW4ofS4OqIwY5W0
tBooi4tX2w7zCB97ORgembuvOq5jH4miLRcD9eMeBSfcK1EvxqE7vgV/mbQjKT3G
CGN2YmCCrs7kAd/Ayfh2B45r/z3Z3Z8FQPQL60SFd/dl5Pz12KeszQyjTSElCLc+
BhnsmOSJxSMWLZFlIsU+TgdUyWHC0YdkKFIPepMlXUXg+uj/KZLzgeX5IcQvOR1t
3y+cMfGcIvi67q9H/qDH0GAXnhPgt7gU1AYC8Ii4HGlXu4q68bVMNdFjLm6qmsdz
h1j2AU/ase5TeYS2Rp1YxFJWsJ9rPtFY4Mgi6zUxqiK/peAY7vb0HOwb5WYaDf3y
xvqCoAlE414BV89+Iv1AEcBvdLmTnAn75lPJ008lWgQJwWyXWJbY4evrokbOrFke
2DiAKig5CpnlKpLKH+CbxnUKz9j4OYPVV5IuHIToDMNjgeRk8Q4yC7ogvpr4fA8s
kIsx0wxUS7T5ysC1aOKtP1S0wEaQbk5NhHmpSATMrkkAuSW6QxYt+JAl3o0qW1t7
PodFoT8COiRCC72mMcj8TJUqTpte5tbkPyllQpE1QKKhUn7MbxHZ4U4qMymvy+cs
3A69d0xgQAUOGz8Sg9znjmXCSzXFTP8CCR3Vz83MciBD0RDnUB4v1jPMMK2KiLzy
gCZNxM5aPNKkdkp2JKyI2a/pTQtLQKYror0/V3gcYqnUcxwgKGy9qIJ/v4Moxtv1
8f7Cpn3+vVi8lxQk4G4vHRUlnlarCplKu6Tm2G63m5TlIEJPqZ8aTGkziaSRiMzJ
edjZXrm/g8ZDHCOdebFMY+CvO9A2/YwTUpQElJFpS4ovR091r+tJZMRewDScG0kJ
oDwH06cLI7l1PhI4rEjQzZX093pTfYiyc1Jr1uu6B6JB2qimKK1xswaAzgdOvo4g
CeNhJoDZuszJ2FGKwIAYH+7NDgz9LpA49nNHA5/0DFB5e060Mn6pwluFXyNxShZL
GFjA8WQeeGkaKEVuThQoBP0U0HRf9I3BQVDUVT5jdI2uZg2gc4ZWIONaWMUSvM2z
6BKuOZ1+NR5XiZIdfZcaFj7FZ6bBFoDISbvNA6ka/RCC1Rml3sGFfcZ3+JPv10k/
CUlYnuUTCknKNHRSeg8EhqS4QaqvCcB1Vujou7uelmiTFYJDEC1cHtV0dQq7Yz9A
mF0qNcSIlEv7BHMuGbQv/3+e8sPyjlduV0qwNTkoNOp2KdySq0GrgVDiUt+xBDGg
v+Rz93PaDNebc/g7sXk4sK2/BaH1OkIqVLspIKoNsZ2tO/HkrBVDIJGsmbs1JgsZ
XV9wsSSCznm4HzcCiQ2UzHlj3s4ireyimmnVmrWYbDucA+thzVpDwaFnf+QmG54G
il5+Om1TV1xlFy4d7/USkWLfMxCezK2p9B7eYSOiz5pxnsb9fDk/UGNVi9z3SyNz
q7xSC88fmoMENWMag2M/1B8FWBaH+5Skwp8ZsSgplNdcr6Dm3nH9FfYw+iXYf49n
q0R627fgyRnsv6fCGD4/+9S0WXOdRxw/f7kDAzaHD0WlzMxK448T2ezhsLnk74f+
jhrZxlrB77wYA5egp+AUvFSBwPL05eMlMfhwWWVVywYIcaSItzu46P65UW1Llaa/
BNMqFzdcLwn+3fhQDbENwv6MUWj1ioXA16bziR41ABU5mYBERY8yL0HYbJliwQy4
94tbkNOZcsknprp3wEAlAk6ulCdVIrYdRmlayoCzqwOl1fgAgQPUey2THBX7wV0C
SJBkCXGTVU3Um8F310/AUXilQd6DsiV2epGPbtRsJUL4UXmkfCZlI+UMjiX18rAY
82D+d/R6h1yM5XzBi6EGBIbjUjesYY+izSAOUET3Efe7PQ3u+yT9/RwcZKnp5gTi
ABVicyCsxTOjxpxa0jLZYik07ej5vOPCUa06eh6GnlYcCh0XsnrYqJRzGYDbo/lv
Gqar9de/X6KCo4hnWmuBWXeUOcaVs5TTHv488GppWzt4qJ8IPHz0Rr5klvjBlCPh
UmmpXmu02+8Vk044xlGeAOmosmCyhGxw5h617aiGBrJK+uLzf1mRxlvwYAmET1zU
LcLxpd1w2TQCPQRYTjX1nEs+gO2DonHd8hyQQrDf/moAwvlkhgoWi3l8yKoqdR3f
WWj2glpIdKNg0n3DtXqHEIowV9hjQe73KM2ZYF9IUO0Ts2OUUD/COPor/xKiBH3s
3OjA0LpTBVuamogOH1Yoh0e9/HCysz4uJYsJPPow+2eiegzyshlA/kE+7rRniaRt
POArZOYuUS2IAZ/ijxRMaAAmcJT4YbVlca9Fq02taZfDAB8l4ZO9GmdS6n/AFIg/
ZWvb5oaizIEdclfoty9VfjhHEf6zvx2GtsItQoOgdcrlWjS8c3YnwGYNI3vK6v3m
CpQrxH7wbT6mDbExoWFpn7aaez7kLzSEefvBeSK9xK/gOHUHDmC2ySdb0MNYRS1N
ViBlpwNzTi581qfzMVMenbZSKD3jsNhYoWtiQW1k0VXd1IFN1o9tyDMykn/6iZ6Z
/QCpSgfRuDb2z4gYOqzkUZYBAZ5XABdPXckaMQe64c24flBZnEC03g0RdfvMc2e0
DRMRdeX8VGixKhwuFMkLwZmcizGD/39RV6rKOXLHC8gGwjjkNfxsZMKhxZBQk6M5
as+h81xvjaPMvgRKbRNxUW9ApYLd4yNv+rQYyxjNgFTFUN2Mr//tey5TqHRsBKtq
GMOxr8ewxltxBdowTx1IPQxppQaxv7UMloIAA4CrT5C4/Lj+5xSniNjfZAnzngXk
uPjmOWZHy6G2jIVoCDROfmLn90eFeawJqLQ+KzEG2pTfi+6O2cDD1ygil21jcYum
+GGFSwGXlGHPJUAnSC316eRAav5XKp1uP+jeCaEtMILuBZZhk8P6fQOnX1IVzcnt
W4/yCnhqjkv7PjUfpjVAMQV5PsHOi6uwKUR5t8czk/nSLyNtSCbf2zFDEKTDCSnY
mLzf6bqczjO0PC39QxPrTPGtnBKaHMORSD2t7vVqetF+ulv5RS7kJX6Saq2UEA7p
vtNgVgEdi1IGdZPKF8x8OqUg2OA6kenqVxOCjsgAMxJgBes1i6lEv/Vbo4DmwC57
ZN8POJ0JxOcXGp+Cv6y/G6/PUon5gxjph59YO2PMYy8s+3QttLnVm0tLi2OPIuGj
xTdxGZEcghPPDOrzu9I9wL5ogIR/MfPfUsTVveG8ADs8BuJGZqPBlWUJntjXdlz9
k4hcUW3Ht/Hrq9psVH9RXWVJ2jtTzdyZlc8ow+0hTStkUmMwuyqzqSMG0LnsSNGp
vTeyZ2f1gN23nsXTKJxzP7hT0Ajpvo4mwMuZPcvEUsyvwJ0Za9cI+LBzcwjrGhCj
dHqsBr3g4GAEjRE5m3P1wwseylm1eLHFx5K7LcRGYvGwdOqskwoBgb84ojkJK+rG
0eU8VeZJPSnrye1Mysm2fz4FjOvZ0NFUlXC6lDQ2xYIQ1ZLPuiPsuMCv5eK0OxJh
ZxEbaP3VN1NHNvcYBNBY1/Z8CX3tPUxlYv4qbc+NUAtaRsx0WmzpEPCtbKlHeapD
AXgHB0qtpaRm07xjIQAFfDO3Ec5rq9rWN95bNs/nIqPdWJkg4nUQsmnlPl0TR53b
U2uVdGWlohAD/C4trJuSz2Jd6n13Phm6g68hyjlXchXFUsLn6/35s/ZeNRUF2Knr
yI/qDNAa+mP+O8viULF5w2JoDjSGYVeSLkQ0OMYkqwRoaBDyeH3CfphocBZz1eh0
1+DRom45BfyhN5G3zOaIHNvF/Uj7fVI+3V26dpCtEuXjhhhlt3CLj8EeC/OtYDQd
3oULRsld5qpzUrtauTSkBUMQoHqwIy+gHrBlf2OMk+V+UdHLu4N0BZAaPa5vMki0
vat6H5KWsd0YG8r3IRfgSPX1kWqrtsIvvfFMpRU6iRECbuXysIpSqNMeYkrizMTR
CqJtsb5mcFOQQ6Gb07hMVf82mNcLRa/j5v5Y/ZfMIjU4wxbwWjjV/h4F9BxWxPIi
NDocDng8HSyurgAWpV1yhwYpN5dD5Nm8h6cfBV1X4cy50xciUnLH2go+ih85vwAt
s48NvvOF9FBSUYpnIdkTdira/2yPfvbkLpC1m9v71D3OV0bMvrX1youBpgnFKRF7
vwiG3vyZE2/yAmsfEJNTnBxDKtCudqnBvAV4514b1UgFA+u8WetCgpAPch9zvxIY
HUdtNJxZURH2KMsVan8sCfabzrgqgR5K8Ulk4lrcKN0Pa54X9+NFDNwonHAS78ap
AxuhrdP6c2/WqxClrRabzIJmjQQDDAxqHaY1k9ui11M4oB24+OtWIah3eJJtxSnf
TKnCgyLLaAjri9YZnflfp0B6VFC/YAHD8HTeXjPN698YGhHWn7arMYdz9a9C6svV
iodsKVJ/lMId9sAZhOPJ+yJzsypeXFww2JvmUA5GT4J4Xxxyhxw8P183m8R9iOvC
nZncT4Gj3U9mBmm4kLQFWxARhs7tuAM+NMT/2M+SG/JUt/DSvYxxfg22eYKSVkbV
XKmeQRkwHT27/CnmzF+vxuAO9j9hQn51Rl6sBLoGED5Jnqj8chvQYRAzjKQE+n/q
7V9gA2Q44b7S3DM5vQDRQwVG+dwxmLQHGIT1Db5dQSh3JrtTTYVRm2tyxEdWH9rz
pJKi0lzjM3kIPy77ZqCoQEOwHscWMv+tD2A/xZDtFduJyi0jW/EcSm4yVciEmPZ5
puEoNH/ieRY29SDJXj70q7ronUy+2Py7uCBWc0747YJei04vESg1Ayj9Jxp+owKd
6Av81AVvRAIkJwf/Pd/x0kJqCaskzu7LQBHBLE6xsnVrqaL+b65UxUf0NHRdCHAm
LaVletVhMefjU4IjfPEULNR84WkEkUQeAgvj8ucicQ//veOhngG+BG8GfpQfzexJ
EnkmnG+RtI6/8CEq+J9ugOjGo7PVRU9/+vJmaJGhxRR38TxjOExL8it01l+FGcuh
qO7yU+gz9PBFAYnXvBorcHkopKpVKh0IhMKaZnMC0ghcHj6WDAhEpml1dC6zHj+O
hS5PHChsqn+ZkEt5p05FaOtXnizzJSJUFSbdBL6xbvQuo5QLt3DShhoMU31wUbPg
RHSVI2ujebgxt/wYByg+LBo6/jQw8v4YNSFo5yPDW0QvpayHKF+PuEA7JuTOSdWt
3lNrxqHjeYPxuBmZdpyzKV1Tda8YcpoTwYWUXsU/3P5J+mhnWDrESsuxaVSj8oCk
FGi1VFMdf/ah55FAq7H9o8cGMVE+NFJ0VaCtN4rlGSptL/eZiF61qj0/aXikGXnd
30pX8F3f/wO0ZBQcF3CAObgNIw7Z3xs9mfzhKFe+FCBRrqI+5W3DdC7OXUydITUa
le7igBoKoox8j5VRKfIg3V2Y572f9YBBPenq3lY5z+vo0uQwdkrinoIt6phTv7m5
ewDfwiEfr6v0YDlnhC8zSRfOaJKmqIW35l9KVBsh8Oe2jYXCbr8EwV+5p2364Rhc
jwt8cfiCPkvoMzIAH1VUc0DX5ezZTMKyY//WtWdWDOlPT4icAIM6/2UY7M2qH5JT
PMZw8PTfrUaV0EpHomT9fOOkbxJmpDAKSmkHX+TEA3vpIb+oVQEocMOAdQkVCTmP
xVm4+y8VA1XgFq2AgYL4vjt96kepwlOpTGoQEke9HsZxr6Spq/pAiwjHwNZad41r
sKVkhvqme9oQ2FVQTUpGujIYOKuUjkdqRj1VxssOFmEDeY2S4KNoFRUyeRLDJqcH
6exVyAImCrPZL48YAu5J1FAA6gcTkd/rFF0hwKhD1iFwGnZp7mmCn6vo8wuzExbP
gmAFtiZTgznno0TImiQW9XPY7istFJpVP8Drk7nKAmbm53heIc5FBG9rwtx9bjfD
Tszy4tvePYyf/OaYrVEJengrvaWK7VejnoVL+OJdK7tIaDCovOjmh7jHiif4Lx+f
dsnYRnJuj9S0PE4s1jQWaAwrVMU00jyl237t/CA/Zec7xs9XxfQjNo7XNQplqZut
pR7QoM2h0gkjFuOwHeEYMKXAVgXQHDV2ihfNPsPsmMLCyKCPIFtFzPjsr0tj3vt1
Yw6foMi92tQ8mbJ6qrSD8FWcjJG4CKxwhDlpD3IqfLRWYsSGMrXlW/cIenquFqaR
CZfNSw9bkpx7HQGnQANQaCBDKGkTSOIHwQpTbJMAGsR9Mj65y0kyrrYudUnXxICF
aBzRkOeaIHAJ7KBL/BO3fM0bSVC3VOwZIwCGvBjoTyeeuswzwwqc3KyfgkL/Vb0u
x7hVwBpGbOq1rysdrbY1w8we4U4rfunDqEjiDSfKnYm4Blb7lpDr0/zbCJi2YEGc
96R/VV6BPeb/wo3S1cmrZpY2Dt02xqJVna0JHmvdaysfHP8d9jsd5Apnevwme2iX
69Pg9xhWGXDH2nH29rzLhey+aql/nqJ3KL6C9mP+0LNx/qNMdxKT0vNPb1R71SUr
bU90dsJwaZQkLf3C/E5g/vj8vMijR65Aa+rG2ldRysTzKHHN/iJK6B6dgFOu8MRe
k+33AvWWFyjXHKOiPrxStRpA09A/06dyR6NPy+L6mk1v3tkhWNuofMx2hiWIeTVJ
4wZayZyTHSHyfr6pUyTwRuaj5OI2jkIdTetbY9Pkj88fZzeevdDaF4PNlHaog5sx
Nlz+NveDxmZM0wQfUZOBYXmEpi1RL7y3O09rL19qzEFFRgmzyK5gCn/N8N86omxO
0I88JCGrZWjSSz3xDC5xwcMYkoblJXmVbFYSjGNOjjfagSRF3IJg1QZOHuRppVPg
QUT+mahjNBlFo8pe/yfVwuE0CXumqPGKZeBBJsK8J9uafEPw14AJ7Gc1TY0BX5wF
PaidlpU2rwIYS4YItFqYUjp2rRXrQk998tIlQHHdvUgazSUZBExl+0cGTaVqlqky
wjyFIpIhxZxrmKegImu+N099flLLRb/Egt/pLL8H28t1Gdm7uop+jp5q7kGyJhfv
oXPnAE6RB0zx/iUHduLjEWzesW0JZ7CmxLTGUx45FLL6tRPFoRVfckVi4fsWWd/T
KWfZRg1MB24aNyUO9DfkDrnE64ce8irBKh2WirO3+EMYN4k1YVDcq2B8e8CPEmlk
GlhAKb9V1/KVOGUPcezzywxT8SvA9nS0vhf7QU6MD1PblEm0K1avXDBP1EJrydDM
xbcbpE//q9v33gN7x30/9SwS6bh10U6xbOavd3ylshU4b6YPafopp0mtXrijezKE
nGQnyY/hdJVVQqkZ7uWm40eTmeNJ3+7LGf9qDLw2oQQac1jTz0PR1KITgFS0YoXy
d2/vj6Wa9J2y+a2an0Y9zxrHcP3pZ8vkatyPKqR4ovYOsHdJtKVhRicRTyja9crZ
NHIDHnN81XZsc+9CJ1TmJS+rNipfRGwZ5vb5ZWf44E5ucIJA1MLNF4kGIvnXpqgR
l+AsBN3mBDLmRlelpXPtHqLfoQ9upfufoNrf+MJYargVC//RVNtBTiX3viMNdOMN
AY+AWVjEcqHRBzQVYGAm1w/BE6kq16iAZ4tbwJu7V+/r2FAdr9MZv4OFmXH//DfR
q4+ROC4LNw6/8b3xzQXx3V4vlhxW+2j9xTOXottP24VJFLdZPvq43PDm6yGRQ9a1
pje3X320oZ1HJIkj2Vmd4lEW4UDHCKByQqNU8CV8xPTOJ+52p3B1O8YjcB9R+9XP
Pj6qW7r5fESJGtET/nRAgA1384vLBFPNnCKDdQHjfuPnEDsfmRXQeQVOltnq5q2S
7ftE+oMRRXllr8CYlJbZMYm1jXcRhgu/6kHUTxMICWhmukRmDSNWoZ/Q4qSBvQVW
wXAmnn/XELdEyZ2+3eDVSFbkV+wrInYxvoAiXibm6Bx+i+BfbgvVIXtE5toRrVWT
hg03/9XD71AzEN0lIcyvqp0/MmOk2LEPsRuM9YRb6PQZQk3QuberJq0dBupKr9W2
ORhK2PVLHIpVCsMo8qfXlmTZNQToYTc3wNOdtdLK6Zp1If1pVLKt0dE47zErIbhX
HwNIfNBUFZu26t9rUZ/JM2GtXH+/QpXv64EQj/ZHsEhQXrV4cNIOqkjjq1j92syo
o6ukYifdbPQz4AT6zIFR2Wu+7cNGmSa53oL1rgMeQ7CxFuTLTr8r3barfyLQwz8S
JbXnbD1q6v8lBAsh70ZnyPQXCtqJ2TYLpEYg1axNQ0K09sxEtqimauSLP9NSZ6ev
3lerL8tlN2Kks2LXJLPDxCBAMBl2tWqEnZgZVsj7w/ViofROftEHQ3cTqxlJzUR8
yooQqMBtRIiP0XZsraIT4oNmcS+s6WJ1NBKw9m5fGLg7iC8xzJRm9mRsqCLcXxu0
1waL+HSV+S4rv4VKXO61afjkvLFHIunuE/1rR9wNj6B3UUMDsIIZlJNqUw0LxVF1
u/LkY60B4IXS7L32Rf0+NMZSzJ6cvPMp8Qdj0CXjMQxjCDXXHOkVOzcKNYDvREzZ
7CoYt3e0MBA8ShFh59dTlucl3Gav7sD3xG1u50ho9V5ZC3MptW4UsRhZek8J9hgi
dZd4oGqQuCShxas5+Lwinlgv/5WUR1JJenro7ZPmfiR3CMQMS8wXUfiABMQHuFES
+2Z4kzjN8AO7S9ZXFDHTH6GbzTCk3qPpuEuLud9o4W8KKmoo7HcWQSdaHFRdYbAo
3YlKPSpmFtYSiV56b9E5OgOQ0R4+Q1cnWebbLdAITxGku0K16QFHWwq8ImbS6Y1v
aKQcBfsVziMCDKOz9UHLYzi6Jr0CmPWn7q9z/Uobcz5OkdB/5Yp0g4uwsYumIKot
RpxDiJmk008ABg472w8s64QT/82c67PrRzxiik40BkGkxgjr+rjeRB4YEuKKZPXY
SmSwwyoG4Q37A3xOiV80KvdCJXfbi17Vfc1/KsvarLYzTPklNQHHvk5t1hK3/O8b
rVSbKkRacD6nyef7OU6BHEHbgn+qND9C6bUUkjW+NqAVtx7zjBEzv3cbY+yKBKGv
JXydqyvdL4xHGxnmCOZKo+FqjwRTCgbeJRVVF+rfcBaTW1SpDFGTmaMnPjJAcmgX
fRWMGy2zO8pNqB1QRy6QMzRPCjJnCjJ4IE/yL3vXEakF+d06nwZSFJn9wUC4B239
IBMRM6tbAY7prwymZH1p/fQVqIaDBs8NxemK8fEDrrcUwZ8MWD0Ofqjm9eCKUB51
I9v5Sn97j/Xk1PAofjUwl//twkKzQFPucPrHRlmCC129D1vdXwbgUxCveLS50tGY
/x3xH8PYwBXQkiM/mi3bhMJhqBqbN4czoZ/8cU9qh+dpcdFQcDxKzN9rjVuF8kha
D+IUJ7MWR8Rv0CPYvhVKZJXUn8wyO/KMFt/7o3/vLUP7Aj+LHghCKqfrnATLh0Un
sYnE30+qvCP4fSTu17yXZvRUCp9tRP4PA/8Nb532BghsZ202fISJTFnv1yJTWkiC
LIsD0eMImahXvZAuGB6IWkzQdsMMYJ22oNtQ2p+FHFxful40Mv8QQexvMcdt1OtL
e9Hy1pPAfLNZnO8WTLBL+ixWVZiQAPkiTV0wfZDPRRccdcIFLuMpOVlRC+pbdQEw
Ru9ZvemEObjC0t/6B9240M1uXoNmkIHSEwXD940g8PlKGJfOwUWeHlQg+wpleqli
B1U77rOYH9MoiYUApPx50dDgail8gWf9zkjRy/yj0TDY7j+59UyVSqcoPFHBhxH/
VUHzVVBmkDLsGklkAzm0JexDmjMpcMUdQ7eZyTA8OZpaGSuGd1P/WCM7s6gDwUtv
/EByB1TwRn9Nwy0hdExGdhyYr2UVAYCxu7Yr1QLiUe/9TOWXVVErOKNWOaOGUbNh
bYk4YRDp2QOCEIksLxEOkrVt7tKGSE2DqE0Bk7XOt19vDEty45BGGHO7t08iagGR
81jm78HIin+EQQ6xUDYFwI05jC+FrwqbHInstYH4SHxd9U9kIXm7qZSkolHnj0T3
JrQBEu4hqT8wfjEGidmILtdVjRST6+1L/Gt+eHml1+LiPSsO0R1JSoIk1CAgdUPs
b4dKxz9CW9ZLCybIkINt/dcJUU8EvtOWbQ15m1/fZj6Zbt0Frbx7scKVbWrHSX45
BPIw6+N3GKTT40ZKaLZmXudP28fzemuc+lMFcZd/uf9nF1Pyw9kWDOjehE04Dibb
2Z4Es+C38hDtJeyzzInQtJBgXin3+vy8uR2Ov8jvlXJT0N1gnGfjbK5xco0/ZVOt
vJu/5yHUOt6XDE+x+WxGIPEywVEHdM3xt0VE3BCL90on9fFX19I7tiEl8XRHMCVv
wyrhvF2YSA8KYDTk/zCfQRXnqhOTsgadv13jm6Oy9lvOWuYVBgK/43VnXrcRKo0D
kTWyhYOZhK19vl7PBJK8WcYtemJOvw3E7ZWQsuS1CVQMxS2ems5Y8+j0QWVQ7taD
wZpYANnJYDuruXu2CrEgZKA3hdVRmVW7itBUsiV6VR3G6hfIqHpF/nTpNdUC0K7a
nL4WO3a/cgtfma40LUZTHCIcFNqkjt1m0kxXYbw3TL8XoATLlJwfEfxgRfGrMDxe
+RPiWb7zvwsUPUxRlu6sr7AZU7T74WWTLgEqmuCvBiYVziFdLQijwPRipQs8tIaU
uJtVHV+vLR/yDFyfOfIONA1fjK0/lsf89f/aAhgoBKjOa9d4hmDDVFcWO9u0qJh2
k3LP5XoFFhn85sSx4Fnu2gwUn7sKmxkuiQXCgbvpKkKuhLY1LYYwqlJ7eo4VsQ9u
Ia1qpeNmICbUxYRlDg4Jpd9szWoQbTbZpGZot6n0kDtWTPISNpZZ+PyAWeaRxvhI
1najo11w2fxZvpYDBQgKl5KXpxzSgtm56jw0zIfGl0a6Snpcx4jqGFTziBNjQ8IP
WlmvdYW0FO5CBDPYrq457IPqaFCplj0PoF4f/iiUBA9l88p5kXJqeRYqqmOq4FPf
c2Q2p7ptFzvNzyNn4XaNFj/ogN54Sy+saAqH6u392kkL/Y1+A3B8AAEwkOY1lddF
V1F9xO1ZNKmGctkseKMVhifopFevzcuZM9wG4CUMbJASQmgmurw7fLHO1gbs+a0e
q0bO4J6Q1+TUDf7qNCtRhBaWJT0PZJhXOGFdw0zmWBqY76wDFLItraBPZ/zl+Vgt
l6YSVQBAA4hr0VC4d+bsQdo/HZ+3k0G90Eb+xdxJWtp+4MjNYhWBT3WaSmVyPVbz
nmh1MmNk1LKSgMiLDCDVAl0f80i7hulw8NT5p3op6BgXInELi4tDQbneJEk9hIVZ
iIcOWSLCSfrKS4OBD1Cnxzim/4qR4mX6kpqVV4EjOrxwVe96qAiQCbMefnT0/OuX
311qAq45ottUMKgeZZQ0nnnew/GbwtVNpHTbuo5snwwckmM4RWGhPkWZA5ZScyk0
9OLb/I8VURNCXi0srxLHEvsWc4FmmEEs2kMbKXliHcFJAuscxblum3a6GqOTpmGQ
Na3ocrWGQk0Lw96bERibGddln/CfLimps7qmg4ZNge0pX9KwHKRE8up0baPRhRQq
YI84kEsHk9jPSxcldlI97GJTNiwD0Rxk0iX4f9YBO2PT6sLcJVrJvg0XAQPz8aZW
eX5BmgMwh/d6+F1pdfWXO3CBaFd5BLQ24Lxlr2fnuWgLtLCjvzJr4pfbgCXU9Yhx
8Hs2qFDC00wYQyKArow0e7e5d6YbH44rF4WjEh4ywMIsn0GDG1cVXxbjNsQSgkWP
1WnUY4FIt0hMyIT3D0LO3TooczBdA6FtSkUvcClj6VmCI5Jv+6y04D1jP3fE5bj1
exftW3G8/WsoKI6woX3pc/xdECQvCaS7mKH5kkX03TdYSGRND4Qt2bGVdaoBBV+R
8EwAg3NbA/03UDZnTIAWPQwpWgem7JfWApIjsF9MVH7FD5Vq7+2x1PUGDAopsMG8
a4Qb4G0Gp/WmOjvvLBFgoIrD1B6ZDWPpNOVrC+0ujncCwlMZaMHS8gYHsYbCr6z5
XIW4bali0pCwMUc2esMLTx/8ekSHA/7Lcs8/LH8Am6qejz4oTTJ4pWVfGcjHo6MG
swUi1w3cnak1qs1NT5B/P/ADJOKH7Z5rKiG8V5B/WwQJeO1b29ZISb6RQe+JHEFE
fOUtpYCWVd+vIjhUkFqSMNorM5N/N6NoXa8PxX01UawkOdBXd/L+w3fWJ8mp59d1
djhSodeqMQ4/3Zsf8F1KrmK0ABG8jWHHIu6ao426E6AtTEu19fB0a892r8S8hh7q
1QHk6KduuNk1QpGnGm4Bgg32rDIqKEfRTh+KSB4z348KGaNJW8dMuhyuW1wDyCMx
ZDiALDcGm9JhRkJlU+FFd1ks9iKEM6P9zg6L4LysOFd9bsr8eXhaz2oYPakyFyYR
a3iHnKuz/wyZvdOBCvUyLujkeXEABwZT3S+4y5KfVwQtp4+9vU4KwpcZ1sSgPGMj
hjU/qfaqQvLGdF8n6S4Ba4KJfT9Cjjx0r/C6JW2OYrjc3r0Z9cnQvgDzuoh8rjnN
iyPQn30PuCnwjJUbZkaeuY6n/A2RJe7XYXcbg39OWVNFlwMx8U7k230h8dDaAE3M
iXoB4JYZcAIXNcnETUiT1aFl2tX5XdpPNvkeU170KQxxTvAXfAbdvVQDoEcPuVkW
lk7qKbx0MyrPNDW7IJsI7J/KvO8vqEGgY5Z0JYArQ1eXkyYlUYIv4K5V5NW/lalN
wBi9AUspUyP/2t15/ZOUy/dvfwFI5GUlQHRVG3RCMOK1UZZRbVC3vvxaTXGHkzUv
/rtgTbqohlosQEj1QdXRzjOk9ugRJixurL42mJwTIlukQW5e3FOBLetCLhxerVJ2
GdbczoJqNve/h8JLqjhDclGpxUU9DAO2VtsisWGrr3I2mKYUiF/EEHAS+gyRnKos
/2LJUe7QGmurmaVwvnKcQgZoKlJYYhqS9yos+rjv5zFeFvXefx2jYHnXbUBSG4dn
N6uJ8vlfB8o4v0fQ5MuNCN1WZ6cv+D+ChHC2wMu2P1/NTB+860MbSNst6yL3vnSn
WAnCQdebq6cVKqpS3UKEJrhc1Teg93izM5n2MIGo0poha/Kri5uI3GngBUCdayBz
G3IAQKIKQIFG5VkyGWe0j2sbghQCyynyRiHy/DRYbDd25MTe1JDW3KdHOc4q6JBF
Dr6/WlF+DC15Bk85a4bTkiiH0nhcYHEj4pw6MQe06qhiSppqYd1bZmUxkucAqdLb
2TTjKrNw/MGa8Gny6ZNuTLZdVs6RHZOWWwhqJXlCKOYeMOR4YXwKurHt2mNS5D7f
5L9ZtKn0wbm8Y5mwQgY26VUIRL4IxexH4CTM0TSy2DqiPaWGXW3F4zpUE+aMSZJX
4INrrWL6cZTWflLCpa3svsvnXooumg3knlDrIO0SVxOYezGYQDfR4ZLhWth8JRpi
VxYARlktAvZk4p2zZZxEniqmBjEolgFHGURb6oF/cm7/nuo7yoqrUyOau/909In+
VWQ7VntXtI2dK/Wjh+yOh9W4uGGdislawCkzx3+pzyJ0BaLo5sXbTk95WociXerq
Ca/E3Rlwv8+500sfZQL7i9BD+loFe+diQCqnbddfASVT2WXZE9Buk0+lCRct9ljH
aoQ6ojZiIp+u0cqDmBadobB0hwnviRvsLHrxwm78z70WGpGPEjshitjhP1dI9Xn6
BcttNBtaAhTD5SPdQ4ZCxvJwI8iA2P7LX2kcsmAb9Zey/cGig5IRTzINZUYWhUa1
gSRA9aBRSAOydKr9Tol/Wd/kAXRIbLVP+nm6tk9fftgL0krAScUXvPxPYjFP2Pzw
J0b7S1zM/gPFmM30ivuNdsOqVemTvwkkkJTin6TdLGTO7B3NpDEU9ZpAJRxRIEfy
ILfYgTZS6XGfravOrDdGfqpCaqMbyYU465Qmkuk3sdjmoryBrvwtr3u9UMoB0ETj
F1YN3XnZ+Jqjk/Sny5FVFIpPlzmEihL5Hnhn+UZrDBpj80PL1RvmsREPQSyV0Pf2
PqHt962g+anKxQU/szUL4E+oovU3vwhjZ0KLUVuMAa0/oeTIQjNMiYu92w2gH/7A
2Sz9ZlDowj/VzbUNtEaCIYdN2d2O/YEHR8BPuVsb9x+HobFo8smyOsl6OwCUdCEj
4R77Huo/FLea9iWqFf8Xrv9fgI2ZtOGi2Cn9oy44pH5KYUvpUoYDllEJNV8bsNNu
y0jCQGM6v7hBeBs8z6kjZaIKEX9Io47VYVajpU8IDNQ07+5uPD6tfyKWnSZHgaTl
Fe2sLyE+kZxJD4qDtIYUvil8RzYa5/BczC9PrgCbBLiuaisrrQDlCjUrmc4graDb
jCRQbYcaay0VikRvaNXedxqhM7iPwHH08UnIEmPC4QeRcxkUIYvhTAsdETqwB6LI
msH4xRxQYtov+UJeMAam5d9f01RMEttfc/NHvR3gleBNHDb+hHFVixaPVV6AbwVo
MCoRywMsqw07yArAbiGMNga2ZnhuVav0fWOpxz0o+yQovrvZxyZIndShU/6ilQeO
AmVbFdWI4wFfpBpCRwEoFe95zspvrfXiMl623RlMLSUZPAegedYRB6bek1hkrRF8
qmC+TNaZJF9eelaTTO0eC4tZDYxEIQCr3YLKBi9drjVKQDoU6GjuQpbywf5vDEU6
KdIOVbLtc57HmQ4DFkFpQiZgdTkEXUNiRfe100cQ+jlZrQ0ZCw8m56ag5Q7zDMaK
BkvY/+ulzZ6pKVoDBuF7DDonwBw243OLJv4pCxrbyfmFViSeh002Z3x3L6Tj4His
9V2t50ECJsGjAPTfx9d60+YBKQ9U/guKB5YdgqFaUewCw93PEGlOaGq+nDkuwzPI
27/Dzpko7+CU+TzEWoGlgoC4Wa05hupRL1XiS60K5RFP0RTfu1B7Iv9XD7p/XwQh
7xmanQMvGiN7pSwcaL1n4KKaaWJXRiHJgH+mWWb4hgkh0RRz8eSJQpZsw9kp68cs
nG07F1n4UqqDf1T3CNRgosbRvHDzDjHOQm45haVBTET8oJWNTDIwUqkcevt8OBl+
htgVq2RkhDS5HSZZwYAa9ijq550IFX6BNFuOc8sNRSNCEfN2KWViKN2hBdiUdJUZ
NcIHGgSBjflzh/ZlC+Do2lnmpS7d59P9/NCQYl9t12prHr0HNGHTcXIUxXsnO18H
jLf9Yhck8Q841GaY9rL2Y+YDCw74ELA/J+3iGkMdFplV2UKV8ccGMjhwHR6B0pMx
leOJSg7is1OKZkMGUjF2UH0u+hbFc5euD0BM3UHmJ9oPyM/qEG7GuXbGYwKvyclQ
Y8PQ5VNnhenA5725H7pncoB6VQsdGGhBTU3Cmo4dOy25RzV+iLCLuyipv2gpOAk+
gvUoo0Vzr/04qFxv4MCM/gKmvuZ+6MDlhV28lJY5IIwjTonTZlrpFpTrMo44tVF8
DtASSRdFKClo0MQUvDrt+IEt4vPhfnG2rd3hFOkClHA495lQDQ2jhHkNiRXWmhCC
S8kejzewyy4rR0D/c7SJDzK7JLVOXI4yFHHOMwMvcYRzStgUBaZ1NmMkrrWPchh8
ysL5/I70Llp9o0GOQg8EbRKy0qAU9n7V4fWGkLprTFTwYfs/idNcLyFPnDIaCWf0
GHxSgB7UEnYOCVLemqJFk4jXNWpYQnnnvbSoXWoVpEX0otWQg7Q6znHzp51OUI2W
3qx9g3QxrkdTVOWd7jXOXNo8WvVXHHuOnYCPD0ujm1qOlt63wXvDrzdaPaz7aiut
QzDH+gDg8cjvPJw32ODbWJrdvTHVQ3DarpMOlBE2nBrh5nl/vUTtFVVnz58PUs+f
qcALZfchRgCeAWkO+yEf2ND2AJ7h2EyNxKAJinO/BguGvaLAKs98AlPDqn03j/oQ
7dk1qusccEwH1v6PMw9nyDoCL2SakUCRGD3ubsHvQk9D68afrouOOjqGfK0jErFv
k79RO16ssMILIPOcbrj8lv7Cm4VzLpyfRX5kip1IY0BQQJzeRCjBZAym35mlH4Eg
aDjbb5y3CPO9iqthFfWXED2LILtPhyqPmw0D3g+u2tpTOkvRS/JHe+G+DDwiQj5A
a8BK68hgq0aH6TVTUu5bF269/QxuvqGfQe0Q0LuDtLLQm3x51psxEN8Vel6vX0dr
EVWyfGpHdp1aKcr+2SFMqeoQk19U4Q9YTVzkU1D7oDYnDkr0k1Wy7VjC335XI9xZ
T7V5wMchKt8+96hJJ3WqeVoD4R9h0Aqb0vS8frNbdCpwMk/DefmLppQA8eaoxlfO
ltQSM4LPpFpy7q3xkf8KBZJmZmVgY+l/8NKHVlgxjVMw/KqBkbUKpblR45zxDGnn
UfdCA1zZS0u3bWp066QW5+PifnO+HpWC+StFQZiDcafOQcgxXWPN/Mme1GIRq25o
55PLN/mDHFcYvCv+CBfiu4cFjdhuTc74i/XT9CHTivXadwT0bL/z8khVDqmpw2LD
3UeHULxs0GQiadQXEvTg88tYN9qmXhTDN0tkugFtZYCPtNB2L1LP4AD+aJ0vbKum
f4xMkynWGqM50FFnIx0j2bgTDZorzuRJsj9MWuoT9jzoEb0Hvcv3L161jH59gO4O
eRtDomA66Aw3sZbXEGmnc1bWhNvprJsZ7nVTeKD1U2+sIuZfnchyNh2oDUSvhLJB
0uPJ2Dv8w75rmcpFVpdGEgULfD1/fTXjoPA7L9VHkDxMvDGl7hD5fcKmzBSYcWyR
nv5+G02iqC+pcltcBXHtUndgRpseBW0uBgrQDoABtq+gwj/XRqVUZlyT/oajTL8t
P65+HCvGYW+aHj2zIWv7CAOto0Tv3qCJjWkptbtx3sdFLgiAo6qt4r+yolYmSiUf
7R3zvnaPMkbbefOloh/VHodaNxvb41KYvAK/c1lydXE4Xb3CUihxaZd9AKM9QhFt
UosICAP7wHkPnQMqqzSa+yMZePRF+39UjezXp9RX12yUdcTxh6QBU16Bpmp6rUKG
dny9xUqpMD6MAK/yCz1u4zxAPrKDo9ayvXhtWyDIE4RRoed44GC4E4bcmrQDLZeb
6QjzE1wV37RwNada8NP12sKtcQtOpCgTeKyb979qa94NTAuLZ2QXu6fSC0Bk5z/i
heETFzKufQco+Jz8CUhyUU3rffLOngXdKdt9R2TfhUEmHpIGF9L/i0qWHJSrUyRS
P4VXJA3xF4GMr0xyxObp1FovlMBlbPSw4gjoKT80mqQ/oI92K2DvTYmAIno8AdB1
5JPbUfurV63KAkJrBxYd+eK3X/4oZjXx9UgjRjG/K6PBNN7u790MoLI5ge+8JJoy
v9jpXin54xjRwxSsJZY0nAZB30B2dnPYR6EPTl+9wobqDCjs6nvPprxAxTfA1v8r
MmZRTsDCrMY3XOmhKl8dmmt0ocEw4dBMEmQ8l/7ie4XD2TxHGmDTHZUr6NFeAuxF
xmBRmx1j1DpNECqmm4oyv9NROKHXGh5DJCAFkj51t6vj8bas+iqEdemJ0DJRfFZN
/uP+G+XEloDhBnc/Ii7vXB8yrXNVrjTv/8ZwAKQ6o2l2PEDPER8oCiroLPiyepTw
tlEGCz7X01BZKgzf412U+G4re/qjgYopiCLUV7vDXcWbSWAo9M53QikWiWrAU60m
p6uoKVfkJ4se96tIyILXJflhoVqULTknCWd7neyiJj28YlDvSRvrMdiqe7RJFNjr
o9EvMh0rYL8yg4TRYl2VDQZUw3ySn43N5hoKfl6oOwvA5RDJ/Q1AyjVItvBUWS+0
E5yFzJMrRP/2ewCzXUk0NHQ1R9e4qv+D1a1Okb+uoaB0ycgEET1x3kZIMy3WltqH
KDHytsWlsykbyKvR3BpVto8XCBvjEAjvGHqR8EW1L3Fhj1JiSUpEvViQAydgQJCF
kH9Tpu2RlEPTjl9wcGwm23E+5tKYqYXLyfOlBdjVyGP1T5RKjwxzf2isxbqzYNR/
7+uCSzjQGBQYkRT9x7gr1N5Neksfr/DhtvBVqnHfxtMSxaJIELl6m/Bp22Nfj2xg
dhyRPLYFWIfXGwfth25HolmuzUgxgWHZOMu9kuFO9Xz46WBmY2Nw7lFT6UNhLP3J
4NP9NSXXpBKwpyFlA22tNhsTqnJpUcY8yFWgblDSXkVQ7jlpsYzYARg7+WsukOYg
8T7SN5G1sgKrjJ8JZ+VvbGthTyIc6xwzziBMf7IGD+++shW/DBvh7sdp2uUO1vFh
NGxEZrXb/qKBzQcW5eL6HBfL8rZDucTnhUDYDF5qfnKmpVQzbHaZykZNxsDf+ROg
sNIcW8VWjxcAnsMUisivxVl0WoJ/qQfeyNfAwLkXQcAqoPBw6Lk8ETz1P9EGAfDq
h8DgNQZPZRHGUvA2VaGbXJIB3iGHex3U9jRp9FI8xYvpYp4cwI7wNLC/CuWIH60c
jcl0VMoLUcUBUiPkyCNGI5SrT2fFYrtRQ0MtR+ZgLJUgBQUtmOp9mFSKLl/JAiKl
H47hBPcmv07A8ITSHZD9zOa4ZknMbvNY2wiGCI5oXrFlDoVJ0nzwdQ3ndAhfbUpA
Fpbzxse3Yv5jflUVTUxGm2B4zil+lj0fVztVwYxyeNL23Q9cCu4Rg5aHmQ55yd5+
bhrGY2At/nngBuYxnsKWrRUfZuvWaxfSQlHsb0Nw82j/CP38MT7iunYAl9JM1kAi
y0h4l6SWZuge8FORvc39UBK44P1e9ILZtURhVPTjmBwpjkL4eW4IycV4Ryip/uxK
8he2DeEa9nE3C27EC9EzdEt5CKlq0EjUb8Q83y+3FHso1PfJc4pmxZ4pEUjifju5
+BjuKA20n+n3UODMH+PtYYjq0zCajhphKd/3oXLUgXXh2G5dfkdr90hlTh2wUcpy
Zk5JZafeva0ZNwNhUR5p7J0CZL46EUTMQQc8lCrMpqOV0hdryXwM6pBrG2wnpzlH
SUPEyWuZ7HLDlQqcObubtYP4/HShpJ/vT4p14RiCRHJa7jDR+iHvzGNqwU2wIGVd
lQxGqtqMTau1/6HIzMLgB6aA0E6Y5mNCkxl4/6HNO+eX2HgM62tqNjD8bAGgvuu0
8kdRgOYd/AlDAmTtFIklsfCkyYeFP+fmtiPLgHCaOsO9ctQkVkdvMLrvtdFOxWz9
RWxHpVUr/jorSp1wCOFId2YbuL9/FK+4JZ8wEz4dYY1KGS64L15rJxxAejrRNQRs
eSs8anztWByQ48QLe1p50fK2G4Y2k/NfyfnwDqXJ/fkqrhQZEsugDW+XOZSINTpn
d4E4mLf05LtTfwlICvP26nJzm7jVoJf/3dVbBO6YrZdbgvgpdhA+yRJ+e4xLpmHd
5MQHYottG0Ku3kEnXTuF4b4wz152qLu9X1kNPswgZcPQCWpzdlg6eDYQfqI+Z2o+
REWF7Z/MzMzX1+yadF9Lb+cRj91peb6Qd2lkEL/EMv4ptgXBzK3NwVUVS9YleSeT
WVvH+66HhBaKtqIT9Q18mOtdOtQzZ+/g5hxXUm96SVrgwpYfKiIFn4mBKkJ+VNqb
fGVs+Z6EL/xizpUqCowPN0z9nWpV9aH4ipJAAgPl91x7yxSP/7s2RatN7yDyK+If
Vdym9If6gGmqfW2JNG6Wo+5kdLFIfI/C5vtd/f2C/glGTrs2fctzaH76+2UHbYGs
Y75F4bB+gabWWTUpyuDYNKRa80L46WJVd6uXsBhnIIJFvnqdnHsGyUHJC6CAf6WT
BUhD/jviSfKSEqqndiLOW85XKIqohSRGj8S2OYvKbm910VZ35pA2HxAmLMY/E2Ea
20yoYlPT7xihv9wRDl9co3WBFviPEFhaYLFeA+QQSI2fouDdfaT6n+63gTIiKNSq
msYVlvJ4Oem4m5slbttKa8znFvOB021PGUo2ER8fWpLd/JEKymh+HsHlqFjqkUmG
WcrllVJCxOX0zgaISpMYMYZHFf+9KLX7H6J6iNXHacQsvJ3V5jOHvbfuRlTsKRcT
LVQdwJGG33WBzCCoblJpgOw2QpAgAWMFSSJLogxgg0SkCeQWeqz7Do34RvJW2wtW
PkmtM7NiS1Ja9B8w3ZkNJR1ND/qwAkF+4UNxc4hkRjT3HhFbm3u8Es9uUj6SN/Zz
skxHjJIIYIBgFfdW9ivNIdjOA/xYSVu38D8S3Teo2FM+gltHoeFKN+GmOXwaADa4
Pe4CtoPY0x8Yn6F3FHz5IfR0DT4f3/RDEcnQ3XPakmQP48IqSC2Hf0/NouPEFzr2
e/ro6vomv03P0VWVAVxHhXSjTTHh7hHnjP1W1OWc3535fM3Kxzt08xyEDWoO9xpM
zSJJLhMFOy7EdpfSUKCurKyKUU1VWE5WSCuUdoRsZXP9h5rWaDlRyhqD6oiEif2P
7ZOuCnggc1uBpi3zoFpdacNQkqw6ysjF8P0ApmQvbLeZX90WFlrleCnWJhq1XlP1
LQLkuerYwEGP+QQEpgAmaAUiQEMZjhfrHSzAn3rxDl/3q8bNGOPYO+OUNTx1Q/Bi
Tls7WTNsdLcC/P/Dj5nM/yM0zP6Ol4JN19P0V1HmTFQj9oGXFs1n/LAXFLXzPHeM
k4ykO495qGHQv4rsC4hixG5oE0um0IJu8c6C0sdkCqMRT7+H7Cqc9zFGrkCKABG5
Swuz1IJknAqx7aYYcVAzVSB13N5RJZXphCEHr9e/QWHwAmIjro6XL5kTMmpL/IHK
xph3MB18eX/SPGVT/C1zB9isvHL+p3ivzXactuFMs9l3AwXVqIgS0vnLiY/HF79q
Rznyg0Ml8/Rzbyw9xe+knCr+TxRnxmeBCxz/zKoqJUaQeVQ5tJeZEdzwrUAslkzA
1WYWJ6aJ0BAfVuFOWAQUSCeM5cwkVPUBURITT4aHEn1NoO50A5i1KtbcDomaQZNS
den4C1keL/XC9pXlgFiTKZjazfF/LNaCzJIc4sAShLfQbWmgMQF4swS94sNpP0Fv
uhBHfPyaYHsLU33xxrk8O0LfCh1c2tUcw3F2wBnOOHSMsKvt847dOp3VeNt7zKfE
wh1oAqo8Qfs3eQj3M0ugfOVsKRfDYnSG1HBgIhlRjzMSN9Sd1PsrJeHD7P+e9/qn
Y0KC/G2vMUrg1cCGOj9IGJeW28Ec6t5o6cb0JuoUaWwwAo90oqtwwqaKoGl991uv
IrWC7Wz1Q+Nh+LzUVtp6e62tz8qYWUgMhgpg3Hy4WSo1UXxlccphM/SwsqIou2DX
KSpazxXubMZWEwpj2S+w28q8v1b+7si8mhskwFTXYMBDqgAJ0GYFmmZP9K7cVCM3
tDXr9Dfhcklt78/u/3qW70A2V5fdyv2k7U5zxWM6Zq0JnYp3jkRy6P0kc4zBlgeD
vZL+tJQcUFTcEqKitRhU5pt7XgOHEIS0o7kOGrAKasvpEfy29AjmV7tqP2/SmOn3
OyShssaXOoK1C7pX+2LWBGFgQpbGR+A/PilTHx2o51pY4wo12agTS5lBj4mWAcjQ
HjXteujEYpkmOLP3r/VxJSVLH8uvADImXgmWiuzXarZg2RwBtu2fHUMyyaGUlaMY
A3kp9Yegp2iYNSpUHq+sU5gVCiY6moHVwyKwQ7w4xNfk+ws/CnB/9aiRubiCAGeh
V0BiDcpLgfF1e0oMFcAa2CYNB4H7runPAhm/7SqOF2qiXVRuik2EjfxfXEhYpeHL
k8RKXbjtlZ08dD2Hp0cus0amZdOWjfzvOt37xivdwJsKLn0ZE1kXw+0AdLCwrXWq
8XST1VPEIO1aRZeNxSjcDNLq7jG6qOYdnFak8X5fVJibWIOIdACo3y5Vo6EDkxFE
W3HEiqT1EFwBoa3MkYx1X33L9Iu+huFYVEVi/hDD2Mo7pcaHNGcggDJa33nUy04a
nsBZJ0qfkR6tas3FEm82IpBz15AIqHhBydviRTsJW8yn43td67OYbzPGVEIq1bdq
NE5K4UuaJ/R69KEL04fPkAYKMFwindIi03XFiZfMX3D26tN6ymUjnKL9TLeNoYCH
N+PzZAmLigeOnjyLcntm0goVV6hWkXuNETUumsoysGUugGEHnn4b3lhEhSkuCVp6
KBeCQCaLhfOp3gLacKL/mMEKH6aXD6L97APYE3PF1KgoIa3TpQQAmqdmPcINPfQt
DxzoN2gn7TwinxE5rLmNOXpQbYuiaIxiiVLPODYp3wQPgcB9qEF68RUsC6hIyvkQ
RwrDHvp6KqsLIccIrn+ZnhE2MBtU1DlTead+gCuQlIO/ylv7QdYI9Mf7opLyWY8U
Da6fN02Jq8AKD9PAT4cpF8Tbgq12BnMmED6Iv9VAShetzQcAR+2Q10pa3KIoz4s6
+Eb3AgniLNTah6cknMfLSn1yWOGY+hJRlggNHHZZvv3gNkLYa1yby3bfyKkijkFz
0/vx8dVHLFumH/jn0n4MtJPyKySJNn7YxrbPQvWmUDlhY34BG24Fk1Ti+4tc2imf
/K6VOtocUJvz+d7vBPXoYXMNtJJRGCJk12OsqV+ZQqAiqnmESHBGIaafHwDtHRIl
z/WHYpi/raJ5kKsPt3JZWdMVtyw8VjNfN27abM5GcrbPn7/qutZ07uZvNYZghH0C
ZSV8aQacujuH6ejCv4TUUP2lKzMXKbuFp8K33q03XYhBMlz6EmbH2NDUrRCjT9Su
8nc3viTOL8hHfXnHbSpRbiaPOkqMfnhL7tASN6ylCYLYgkXkTIhrkTIenMZ5UT47
Ou6gSVyfkgiATLVMSP45MkZKdXl3vXiV6ENb/tmAg5+qyNPxyLPJC4AGEEBOb3Qx
kbtt0CAoxTNo+BYkoK2Xff5o4xfzYdsK/tN8R6AvBaj4n4+Z6grt1mXqMictYMqs
eDhToHfuznGLH8tNNl62LVBZr07h79F5KO+2XASzkAN55R+gx3qPCblXLfJ1BnSS
2TSurvGKTkko8s0cqznVZQVE7r2zT3i+tANae4w2JwvtZ9yyvD/ltaKiaEOA6iS/
luiU9Q4p7fgEk1c4pIKduv4hKTsMnQrdKWR7kbop7apzqyntvnlwUUcV/PYz4u+Y
PRIr+Bq9EKbLVExxmELTQLLEB/h5tqyyr0edEDgFLBTqNr5ynzsdWi8PLprBHhlq
uxUcIpY+05nlc/qZpwlWpx6qk4WzpeZa5awKgw9mIzEOwzMiMhFljJlLy2iSRlpW
yq+9xGxmoaA2QxQVIoT9iDnYFaocDCW/RHw04DTPtO5PEq/vNnOZbZJn2URQzNeP
5S0qpKxOqEmblnP+iZEMfNCchbA5l9pi6Vbq22wCcW/RRc25XFcvTU7jrncT3cfN
8DVALIaE/GWd0MM0GDCubHOwfbNd02EYyZDc47q5u6QW8UfhEOnfkPMgoatyucU3
WLUOqos82TP90AMuuMOS2iWLzH/6EdiAyK9QL1ElQtZaEC8SPmA7EBM/MjkIqyet
prl27P0dchgfQ9aRd9V+jSxEBUudxfu2ioFhXSGTmXl+iBqTN3cKthbEZzFOHQhb
VwCJYRadu9RF/z+MRHDMcnCzHkFHRjG6RidP9vwUWEaNflHPggFYsfOsz43yhyNR
9/mfgq52HevNjWVuCI2zd6yjTXvbqmwm9oro486oixiALjn+zbM52QVcYxKIj0j2
sKr3BoGjv2967qxUuqErdXofdc/LN55anqV+oj++GqeQwpVgm5QAf/PCgLgrirFe
j0MORBZqvFLLiVZWYkN3s6JzD/1oTv2lvyns3h7miMJq6LIC1KfCBsi6ij52soLi
n8ySP/0pDZ/sHxeXpAPNfx+JxUIamxdNrFKPP/ybeJPi29eJDoiQZHCj3SSQBdgE
Wk+Ms2pTtVabiWxzQYGk8oiFFec2WY34id0li+bBq+EgW8nLzlmVeRQctkfmZYBA
nH/CndTuZOMd5N+G39mIjo+Bh7GukYanr+rufpTqQMaxD38ZNUnC9GGUGtUytDSZ
HRsOMBkAtPGKYvyPwZ+jiDBtzeiQgK4ARzuasjikSTofRrPVVxKTo2bSdLW+4+CX
FfUIFpIkGtkOY/2znn9gnuj+omTJCWkKyQlZkpUmQ65ZweSuBObebtS5yhvp1Kkz
bmCAetF25I5tIsRo9Duncv5WpdZbnKA1diaPHOSUbALPfk/3V2CCGf9GDgoGefQL
oGBVdBL1eTF4D11N1TIagdcmI+16FTPp2SYTu8hfH/T4iycW7auJGGbUtnra1cpV
qkmK4q64TzqBvtGWVfgSdSrxw/n1Rh+vbX2+bl63DFirTxJkPApqvGQNbOsqthvb
cRnxm5k3AnfMWVVqrvWawxlAZsjfj+jKxoobps4dg0iJO8rTn9UxEPl4PQDUurcN
9Xo3cBibICrRJVMDHsooywbeE8KUN3BcX0B2jUEixGXKGu2akHpOB/JPDs6JdcwB
U25WJFSwdFFFVthkC7jzOv8c712vbGGkJbAD1EPlej4noFOChXzKp6pD985mmAWk
D9szSvnV8o0s45OO2s8mpoMkpdaHGXv/YxHvrCt8po6/eBxN6THwpMnYQ6bcpWbE
ch0vt99rOJ4/3Bde+nGOjTz2kMsvnbmWIiBZhOefhyfLQek8GWMfc/IoYfim33aU
9OpML32NkIsHk95clMQcoHung3UvzKHMOcP1DCFCI5lrHudhI1TTgTk+HETwxCSK
4hnYYQWj7e6unpCaQe1apEBZlx9Hf9t+Vq7zTtCmySd9gj7IBYaFokLqZgZ5ohuZ
4VHWPQ7L4anrteoTWAwfzLQacH3xgnwfq04lKvBSVBGj7sluOK5e9iTLEQS4m4FJ
Ar0LutZcaOmuoLpN+ILS/ux9eLpLatXKL/2932lmTxAH7A0StUF4FqNMwP+eQ5SM
LZevSBp27AcsFIjrkEBPZ09yiMhPrxNpwztuuviLSuiNceOI3gSw/a0pZ9APxYvb
PZhJe/xxYQ0WKYjBwi0NANxMDSkqGrdHoVV1NoB1S9SlAPQDoWKOIaD0vvCma+OU
zrn4/7wtVWPKBBJ8iqLx4a4tR3yAhi5trNCsE4TYmvECl8mB3NJx4jK09f13CcBO
PQ3VH83k+2JOfJdHriackzV20Y42qJPloUEoMe3vHPQz/AYPe0GT5f4VSYJ1l4K3
4z3SXC7lMpbBaDr0vxQtYLeTCl3L0C3Lill/OknwSXCS9FjXVnJE+WRv4zEXiNJh
VNpjwRbBVY2NsTdDhGORdtFx1Lf1KCUCqOQ2iq4WmohXBt44ASNv3yHrj4d7u8Wd
gCwyHxJXjXY+noCbqC2/O1O88fUoHMdFiiUsxnm/Fz1q6QaNvWYlseX4OHxFavY+
9nT2035Hbe/4KwE9EzXNVpQwDXt63A9BpPwLmazYnZ6yHTMKPSrxhaqfKi7T7NAu
P0NZIFg0wppDe+MZNUdKKww7UDzgZusQCLN1FjbuUZFCFSRA/W4Y9yB4oaMGn4xH
ZLGqGyzVRFlKIhf5tRHhgbsq5KhJX1Qau4pHef/5EKb9XDGXqMrGhu/NHiacmrTg
Wdu5E6aTxf1tRKbfLXab65k6DlZnwCELNGUSOc/aNpgAf3itvxDVMsmG9i1eQTee
Id0K+cPfNj2aaOQEQH5wSm9Dg5nyvj6Es9VuOdJoCJd+7fNyvS6yOGwW1AwfJCAm
a+QdKfzSgUeqFrucG8ktrFFfYxR2w14C20c+ZXkl2E7kTA2fBdYIuzz1jX57gAEr
Su+XjYbWNfFiyglVkyVHs54tO0X8KHzvoQ7Y/MQmz9a7XiKf34fORkCMmZRV9slk
RxxU1iqpR7KjQtj/tVldsEqMDw8zrL+FvES78xt40eq9N+7QxdFCd4XjRLqklo6t
bQnFjXZV2NXu2uJkg9qVQHH6drw00KmUJGC4x0/AoFHt5dIBuioM2/mOXM1MtcrJ
Q6E/pwgSvrPp1bxP9uP3MHupyUnjwQGWLG34pwDIzaCpobwGX5eImqGseMFgXZCN
9iWdGE0xKx4aDjeOpHCzVTbQK7wTwnJrkZQ/ijf6hSf4/tvXd9MnoHHjnM/0ZzVh
TYawKCw2Qk8C1YSMddQkRoPXobWeW/6wWiFtrjXYBd6urKrld7OcT/TWm6H8Tl6J
4A1wOg3OhS1DQysD8K3TUK5038IRRtBitgFZ0thnK3jSj87efN7chw6NgeBC5OSE
+ZGcCMrAHOxQJtLgCtWCavz8THg//IDnl/dmo830uv2n2MDHNMtrbwyOP+mdIcze
BYU8fvv/R1s8s4JZtWlGrcLHgkOdm0jxDrnPuQ2/H2FaHubp8J7Ywf7CiK7fnkR+
kM47G+N5O35N1zLroy95Lq9GpOmQJI0N2w71POjQY4kdUQMhFOcOnqW1/qmhTVYk
ydVSas0mFjcDMbNU1P6g71MWa/AyjEhCRYwcFhWnwRj7racoQrxtHI4QUPRlKenQ
ioSJp5tsxO0Hd6CHIGggi4S+fksmEDh4F3LtTYfn7QLWbmCaUVDndTif4dzUBTZt
IGEXI5uNLSoDUu5C00tOi3RGBrcfzauRZobVBvotDB/fEhV3aMHMefFCXOFGL0V5
n6ZnlZuvBCj7/aYVIrHFXkPGREl1sVCFt+xpTAqY5WazoL+OcXKsCTkn3ceupO2u
JAHjP6mc/TjUo26jPc6ATXvbyW0pbE2tBRUqKJ4SIfKLETqEUENFyrujYI5VjCIo
hpasvmfTqTC/DOmqM2Az1mhMTSdLniGz3BWTWAeIiMDYKKU02yY+Ue7m/vpIAC6O
JfIBbDyNqJAWcQ/n4qESjRU/2RxO2bWWdqBC9mb7v84+a56S7KJomgAHG4YzONGb
DWh9EQxLgjUFDqSfBALVr1pYZTJu9pFwIgSCZ1w1LX7Ox/Kfy0y0pF35n7udHmXz
QeumH2xJ1+s1u20CLRR7x45FA1k8BE3tDIPq1R3OR9CPt996pcw7hhlANDp7QZkM
dlaMktArc6woB8vjvCCU0+w3PGZv1H7w4fZ89vpRaEg1udYYZqs2GmQ4QRNlYUJI
t4m3gE5twN8BmdulkflTu8pojYSfiaHWL1wSCOVyFRwyzPh3fOaDPzkpKsHZAMEN
/zvKagiNGQo4v664s9FZzU+hweWzgXqyFM4PypkkraOoVxXCq8kbq4QT1tZpDIFE
DtB+HJMdvg5mQCC2zsOBpO6EQMCGsaMNdzdajJ0IkUxx7BZv2uXHWUR9fXJ6H5z0
yS/3QT+BhPuQYCi13Kf4gF4MYH33BsMOmujNrN8AxOcl48vPjYzU18z9A/MwLGom
PeIuVW8NfUHy734kUA/6LE5nTRHZd1uuuktdM4BFt6a/x1YORoy5xhrnWwz2lzB9
o4g42j0wV0vrZCe98SmV3MkhNy1uBaYMfjJ2/AJdT0Fh8VG3K2yP+cJ84bqCtk9O
wXHK3rdzX8I9TmWuCJHctra+RpyomZtk1HzbduHgFIrZfdAdnvFdKGO/LAiRQbff
LF10SDVsJsC/spIczjGferUroTW+F4oYX/mUQd98bog17UzME4tkwY3fFNNxo2Ue
UgcekFyJLs5aN8tclaUFz+YXyaJf/oFrmCPjUhi5w9g1kppGIqMM8RK+Np40WfFa
xiW3dfUmvBxXgAMlCvNtUtUiJGn8EUoe+AL/I1si+8UJgztVEk0SqHZKNd5jxDVv
aY0fasKlGXp+4gbdRwL91aDXIbGjKPnN6dZtfPTeTojBz4VtWcLYOZL5hpbEaRYP
xrAUwsi32bgaR1j5YEMxkcJNgFEfgxkZC3NZQSxjcK3q/zCXqRrtr6E5waTfOFM9
OU3vPUcTzJJ1ZBYYS29wkylf3jxsiensQ6q8+ZvRPpLHGQtxeF8I3s4qNArh2/Bq
D+jdLXbw7d4TAO9WtlDj5+SAbtpAzjcsMk5RtcsL9delyOLISzQH92wO2dokaByS
vFpsTSKQ+vch0sNAYKGy4ihYFNBvaqcPl4YftoElJTxjIEc8R9XM/wTlAAJiUMs8
5nNulDEe9rge+4dBf0gQjtYeEduMuR3mw9ydAYDKZ9R6WAQNQyT3RaG/uKOgaThm
CFDXnW1UdmixcPI+AcgjfsezPopn/guWL+xkRPd52LGkOz0TDWlTj7Cn2XOwdCAv
UnQo535Zq5rBP6tSAwzGDRc2EZHeRkB0c5smb5wge3FNr/Oeib34wNSupmBIEl7s
ip2eqcXkEiu4wwxBoeczDZTVtEKD0hTP7CzA7/5et7vTSQSjZWRXxQg1MD+UQgjA
1K3Fyi1GHxWBRDxoVK+OkHWWJ/GAw+5qF9V1GyfyZaEMessAFTUZiWGhTJlNgNnP
fn/y183u352GGWLABI+URmwKFNU83kah+WeYR//DsxIsAmpoCOSyZ+LYDgBunzxW
EFi8sUNcKYexckAFgKgyXK81Ss9TvLa4fGKYnXFkkDJ6M7M2lqpW6s1YDQ727QHF
IQT8BvOjWpVHUVQ1tDF0W3seblHhhCSCJgOw72K0PsJ9g2ymzfyOh7OluOzGE2lX
xhbi0vEKWnnAk2zjIqUGPzRgYFU6bNp7psyl9F8YM8TqvHL+NBGP9NZNRcr0zJKY
HXWkS4mqFkqAe6nn+xLFSq8oRN4r4HzFZ4TenektycuJeaRGytTV1OedvJn1G53K
9h6fubY00C41W2RTjRcHEznZuUtBF7/xZDcP1JwmYFLEZUy7EDJJQZ/MkpFcL/wx
jsj1j1eZ1zrEdcoab0aqedwfup0WlEnzfjMkwfhu39SEEpUMyYgo9+E1R6i4W+vV
alNFJbOjR0smdk50lk60SlHrIQ2oygiaRVuA786ay1knLpB5v4llEe213+KtqOON
83xgZJGN8V1Bw2sVKVEn5mtHpQvKEwgKpsf6cFnwqJzzSJJrU0XaZ5U66ZUDic/E
K6D47D/xVuqQU7FIJj9Fh/QlmUU2trcBPXK7Zo+UqJywW3GJY8pxCY3598OYO1zo
UXjNpB4EyMnjgLTlIvsrie31zZotw49qxLzj3Gq8gg2uZ9x0lir8Em1bf6B9A6Yu
Jm9x1Ti6XEwYyyX1D8Oflj+gBhO6jIR5sHxf8tLQRv7g+cw0LKZrv4d62cnHdN94
p+8iG2Jsl0T0CLNkk6Qcf8JYmo7iNeVBwG4r9pFy8MhPe9vqXDoWNxafd7LOjSVM
RIyheqaDk9dD6JDwmRbZSTljRlA164PaqPztT5k9zmzVrjbm9r1gLpLbgsPlK/z7
WnM3gqyrV7WiFGEwp65PCKvCklzP4/Hi5OzW1+2ZIvRHS6AVF2YVIUNEEbh+j29X
B/SSMe7hTeF9ASRlIM3w1obIpkAIPV0lNSztpL8yNs7NbBN2qHPStsXSJMV2WFXP
NLbvRPl+C/nKDqhqAMNgaUxafFSYIOMTB50IbRWBCPFZn0wKI9WA+eRForLtr+ct
ciD1jY6YrRrUDrAQfKelVph/Yc1oNZ/TVyXjrvXLpncPAH9kR0y4TlXD9Qvj3Z3c
/QuPBZMEDPjRjgtzPCzc4ez+t4Z4kVlKZ+7x4NZUMzYu84Sgyf7ftxWE4uEI5zGt
KNZJt82onlsMBEmSfM6xQP+N9rKdwBy0hh25R+dsNcmp8WHEdsve0UbFV3dD505t
efjyP8H9HvjHJdZoNhw3D1R0mTo8adbPwsjNcIrSSQ45bHw/STdkw3z3qWX1mvgo
c3/8pm8TPYg7KicIN6WONpA7HuT1CuiYxK0+/fq9uXGBZp5ds9A3Cwf47bsFkg6P
QeskQfWFLpTi9nY1l6T4P5o5jTcw9XQet/S/z26mwK9eWF7woBe8snun2xdlJepj
ZcCaMhDfaqWMzVQdzyyu9agndHXFyGJsZDL1JBLsgLOIyscG3CTMX4GCrPeVKhiv
5K14AvBCVvDMKfjabaC7uZzz0DVtooGmQ1aPFV+5KNWs66HzPKR2Usl5KQJ71oF5
J5IFhEOz4ekayj9/aDIfXvIWiUYZtbV8lmX4oJ5fHEfHC3+lOYP1R2zz+WZWTtDF
d8iB3pEahvSjXyAoWMtJREw0rrHQxd/U01BhtPDhMkiaj83IOFMc0ZHeWhyNjX/Q
GixZtyHkDjfK2aoIObN6GK/3IuWD6nrdMOJokBEwWX0AOroovL/0lXAPrTc+Ap50
IA7oZyEiz3lETWe1Tnweha0AvP6OVQ43tN+MxlL7knZOz9xuREm1kZgDta7pqB9Z
E4Ypk9QD5MyeSSCEXOuLQgHBUZkiMcBBdi/RxU9sONMhZhUgWc4552mLWJ6ZQsFZ
wMqwcvDs2SxdeNajxGlWmZTR7MI7MgnIf6b53WnQLwp4tWjioxux+gE8vZ1x5YxD
OkxlKOJ76CP89A8Io81Us2WQd5AHEZolqs13kr48opJUktSt+PloA28pbvWHNOxq
CykEc5E7L1gCrU9ieDOEuu7w9Q0ScSu/FYqjZ66nLol+lbJXd/msS6TJdsHIZTmA
WlLr6dcM38hAvbB33KfdrHRohAczZWk5FR23U6qNnt81kIjQncTXWSUp7MCK3qXe
vD3gW4tF0Zf9sR+ryy7DzorACvB1BTDlVN8NhBeRFnueE/Cbs5PIC2JP2m+LjJO4
alW53Zgx9plOtGUBHRam74b8QXNiuzFlahQqnU3JFgf57oxIuDJ1um92tBXs2KKg
32CN3oVejMpfhpBxiUnWeFGzIF1T4Xq8qLVguBaGOacLxL/N2NympsdNoh3bwcnC
sVWOe+nQWfPJriUEP3OYeKUIsWwic+iPOoAMGNH6efrkge5lbJmCwWlsjouW1/Ly
CAYxzMLu8D3jPSWBoOOWpE93cxRHQ6qo8ZLK/pHa71LNtSF67TZ6JyJLGpNb0WoR
rVbf3vqgCc3H4WOujsDQb156GVFPGnHaIVCEXJpOpVSC0Ib290I+rdHZ503rGfTN
jn17Jht7bPTBdAl4icYR5C8uxbZSn+rbA5EYRaHxPPPPoXiWk+bl185j7yVC5bJY
e1QyD1JzEUXwoYEI6NzP0QKLvKqhuNmtWrEZu1mxRLlI8OB1ODjNAm2r72tFjjW4
27J95o4p+PzkNKYTZc0wHSQ1s4rK3hafMTx8I7fqynZWvspb3is4JYvOZUiJiox8
+QXG8NVIbZO/fiOaJPBDLGJrNf29wM68UsiU4aU8TJpx7zV9JQN35dq0MYJ28Gx7
42SaPuMVCsTdoCqBBHcC2j9MNvSY/WApe15R5Vj0iRxzy7ExfTkf0Hdxx7yv6OwH
d5qlOHdDpRpJ2tr4h6iAs0b3d8pJAr9kDm1ymgSQxHyTv9BVF7x1oq1E66FB7URz
mUW5HbFvI0Im3oFO1J2B4G9q0G8HWHA1C2qYR+G8UJNYFXsoe833grUXEQJjsHJk
u9DAYWAhKBNDm637xPiFXQ4mI3JI3Z3N8r3aY8WohwRtY0rN1Zvvp5D6KNaaml78
MlpjJl5P9vPyjN9jv5xp4MCauXyuBuYUUFmtbJ4YtEnpmp7ag2k1hPIPABDvgQT/
NEQ8s3ZxuAV9utUogH65B+nscp67bAT2JcBi2NF2UdHCzuTFl+0lc4i7/unyChLG
YiJlElFTaedSrKppp7l2nlFVvG1juO7vaHP5WTWtq7ktaM6fFnNvJHdh96h5Wl9r
vrezMTDoamkEUmWv5t2Yk3x6iUaqjr5xBEKdkXJjDpRbfUtrj8em5y49mDyYirvy
lK1KeXiXnacHzflLE4wSFbLTdAYMlqpTbT8eA+IoU9GlUa7lpZ9FwusYgR0HDKd/
zqvG95tEfCCp7K8o9BnnHIGe+Uj4Yoafx84P2IhDj/RKuywoFP1VdKrhOYOTJINK
ybS0xDAWxLLUr0yHrv3a9k/MpmtU7/v451XteU2541bZcOfDeTVzlQpMeEEVs+A3
jYcIpw1xnRu37fwaZ8dMv7UxqTY6cMyQYvnc8bpMx6F2Jr4xn0ODXicvg9hFgnPJ
F9PHIJ6By12BLe1teNzvYrkW+EkNR76Fpgj42KwJfXi3jfXYtnkcB2H5TfkZF+Uh
VgY00oZ1l1o223Nt3zAisxYrkl/6/Tj6xdJJEQfvkVgd2DPbCXI1lHCl4KJuspdF
pzPngi9yVrNdSGj3YydFh9Xl0uwDXNNkXfUTUVNC1sPF9fisGPBj6CmDeocgcD8Y
eFLPA9GRipP12CnDrvmSIS5DJjyX3+y6iHtJbce2tVIH9g83QPbSRUkP8IWyMbSy
1puCJSMOEobbpPtaa1DOUWOiUMWbNsjSOffYy8dryi9EO9YfnsPjwsX0D4YH+vTJ
jIznmOXw0DYSwFWituq0OLEV7wQxD10/pmV2NZX84DQ7g3OfnmvmdB5LT9iJkqCa
Lm969CsFcT+6RclyGDQafCsTU/EELtZnCVOkNkhfcuM6FFDobry4o+asz+H/wfyP
RbPLi2162O/RON64aPJ482rPLjFBIHhiG6RXNsV6sgCOFGRxJjWcaLBZBg97l2ba
OCjfLLd8obfpu3IOTw8Mn7MkI7TzLJFP/UOy0HPCplk0cvDfWXGLtNxXasOTjSCw
VAp0lKFnMAQvHumJCM8k0MGOrkXW9VZp3U3sIFw6YowiQ5q2b6Nn87hKIJ8r/Luc
QdLnC5qpbi+OkOKVBBC4W2HCzotYjvlJhgj1Uh9ccYqDjJUiAoP+roajMg4pNoeb
2DeHyPl96mDPWLjhQFz4JBS5qR79Y+rjGuA5ONyQt/73VwYZDNayaPGklANLz20B
PLgnVGvyWhUQEHLSgnRf70GtIZDGQobQNwA/lXoGbZie0KfYE6aNnBc3KeFCGziA
u7mUI446Ia8J6ohi9Gx8MDEjEFZnGo7U0aSbrftiMcMJpE0p9ue1owmbwVRgkXAT
MAB74GFjugsgG+w0WPShSfVMBrCgJAuw0p+2uOCjrO+M6vhy9b8NJYy7Tk4HQdqg
bA6J89vKJLdCUEfDDIJMUrbEn23aXd9V7WoP7vL0RO2NLaXjJIT+ukZ9sCE+jW2P
4UO9BoouGk7ief6ynEHdcxaXiWYrYv6ryN10wM9mTNpCDk0tHXwruOT4Du7w/6Pj
ofwm/jublbnexCW0eUFcme6v/8V3/BtzJpOBENhsdTHod07TRr5UsWFRau/9/sTn
ueBBPKa6+ralZyuP6JnDXXQDKO7E07j8RZ7WzWde13cY2JOrzqWqQUSEJd33cREF
+8AO4A5YzskP4ek/LMa80UI4MXW0rVlgIUOr8aZ9c4piaQ/YAN4MpmjlgCvyf3we
KUDbgDXCakkC0ZlzNCzkmz0OTxJi/dv0sNP7zdIszR9fyE0pySMJ0QFCUO/OQ5Xe
5/JBMwlRUbuAgjMs+nLPo1UEl16L0Y1BG9ZIXIj7zLULQ0yclLxD1iKJNQ6agXH9
lkfdA98nccXS5nbrgS1lZOv0sxMkXXGISnbwBrqE6b0CObvpn9V4SKDL+KcYsv99
hCo9NbOR39CkgT31BA/5ZMZd1FBZO0wTwrjs8HrrMMQO5oi6pk8MpuWRHqNylSHq
5GHAB1pTLH7rh460tXUkVxSh5WLhVTkvmAIqL+xBjY+nut4oG6PDMN93Strtc9EX
vca25WZJM/YZ/ALYdEKR3O6X2ptX+z12vrD1BX4v9JfdACInVnilX4fp7+oif2z3
8/4A25oiLz5OeVoVSx74ijenYNA1HWGas+STS58zZFfT6+FBXLGDd9kTiGIdRIAR
KOk5OBVl19caQbEHyxkLcS2cUBY91FpxYB2aFExR7VOjLYZf6k6MDwtg4ov25p+b
a4Rk4EDXGzTdaAaQJwG1H0ICEMSi9ooishyrOVxNo5R4IZjZbFOS5PWiTvluXK01
d0G2lZ2V46CALFTKMniGRaDb6TC4HRAPEn1wHEfjdI+fSe0mrfnDls9BF/OnUuhR
ppoez1O/+VXd/p5wv/IRNtqrnSOEFNc78qG8wfx+qfPfY9yWJzSa/dIm2YkQwaxN
/L+/KZr6Da1jdNap5Y8Sf+p2SjzrhdMgo+DQsePA5xrXt7fkaWoPZvo4xHeulLST
cSKYtdyuelVaFjUa8pAQkkiPHUtq441RHA7Ptr0/Zsr7dqP6g5fURriBUTCSnei1
MRxikGS8tMwP5FF9wLpytDYwNwekubwqpwMfXNjc6EthXAVIec8/5VpqEzR85Tyy
7FvWF0MYGJntFLrdSqRClNd1paU8G9mNE7ZB6E3JY51656sO9gdbFgsKyvvsNVKj
hc+PoYm4t+hpJT70+9mtVZAUlGYMkAcpYnUhgc4SAfQ/S1y4eMaf0DCm4LWUYT4s
kauYB5embICllbLSc/tMsF0bKVMxECLwGezlzgpokRU80fJlqdc2MZolaS58dIYt
cpNDpYVpSDmlOwoFN3uvh9/5ZAys6OwYc2expF6B5kUhY1hdnRZmwo7QAX4r8jZS
BgWq7hOCiXMpsPdux7+QYMd4LRzgPQkwluqBTdxTCCZ8Bft3s4SDr3xIJST91H9Z
0DLIHeY0zOjjvvHO0yp9ibsdez2hdi4NwBr9OEzjRCCmusVVQ7cw9ynZlhDQSSUS
16p7NYYaDtw/lF1GTQ3JyuxCbIhORTHCoFM/ahyvb5YNl4kJ9FKKaoR5jHgOiy2H
iyT56Oa7hD4At/gk6b+zzpcSizSRwou3ZB4+a4DEC/iPR8V0nx/LqzHL/rJlSBRD
DW+yUQERg70K7KsMl9INPUozae37WyIfJiG2A1B7ApBoipM5rqYo6Xv22pCdrQiW
Io55YYgeK1UP+4wYSdd9IFkDxr82hUOBU4QGaNPg0IvbEivqTqPcqMgVYwiD8aC/
OawzkdxRtKEqabZOWlG3dJT1Hl4yzH+jXry+f/B56ZKzTrBt4AuEeDZdkOhsTKpu
q2KFFPqA4wezOTQoHeFiTANBisgtenl94EMwOFQ52T3lx1KTjL/rWCzmTywkGLYs
IpT8u8+wsFAiMiEiB+mhTcS/TgOLY9B8MxRYTWQ40LztJrPXpjxtB+UVJ4LCu7nU
yBS8PKeXgZ9Fhppkz9KO2JuxHyauWXU4NjRLF+qmNnbnMWMmo0bLv3V74BUL+96s
XNFAMUjtca6WH0JmeIEQ5s+tTmlSGnTPyxOYzYIxWoMn+RJ4BCVROLSNbRkgmCml
dmXyRE8jNRw5PVeMBlkmjtQ+KkX9QpfDfJDDQ/YPQ45vXOGFh3eFA2lHkPzbEfwY
rY/RQLh74HWVYNIEnS/5WI7jp6PDtsm2Ic0HKx1LPDX+oNnVJZSzHxhxaGA8igFj
pa9liA1po2VxHR5qjnruoqKwwd98De6hvhrbWqatPO96nxaVmS2Tz3rJ+PLECdAa
oH445hKsLtOWxivNkx9IA1Xksw+MtVJj0N491f7Y6/uxIyPrlFfxqCsY6QUr4Idg
7aYNa3bnFhAaAjCT9aNL7YVRqKO7ERvtaojlA544P+vXtI18V+NQBYCDp+xzoafS
EdPogDdr+un+ydRwRllK1aUAE7W9mpIgnj58mluU1nQsc7VtPGGEpeNuakKQ8rB0
+jWiNuagA7ZG8gcd0xybBxoAA62tWpoOMptO47nkNWK/QyrUn6GlsREURMGiezwU
ERg3cZBLM2xNBDGIFhQfc2d5o+22Abim1nJ3ZtrpKLQ0ay9MTyYw9Pm0/1rlvaSu
bWlSAq9itb5ghXcIuqTCyzbraoyt65IefKdtqaOvvPiGLpw/vs2J6LVruQpkL/xE
rzhlEs6q2fHsVImitk4EeJuI3PEGLRDOonnpfKAmbvYmC1+H9EejjqqPP8AUy2wn
t/noi0bgsd6hMtfmL9WCAGJhBnOvNDuNZKb/pIhpvbC86n16R5r7249Vsz5ZsP9/
ft5Y/BS8/3vPh+tkt4u1iwT1XwwZSFox/TbH3GQbq+sItxQdHi+Z6Dwyx1YRhtr2
zqTW1njUMvDpzBK+x38dWHhwNOhLIF2bGw8m/UC9xuikmMibcfTGyKvcDzQU2WR+
6MpOLPjZst/Lyotrk067qSrCXtzF2m7Ws3pIgphIqQOzvhL86LJEUUnZFCvz+RHA
Cid4ZPLzxa/6R54t5oTOw7N/uh8Wrh+Ptb79MPpdnr/PWRR++GzxjIp1VxrCVHN+
oVpz9g/xNU65zCoXLiAusa5AIrsI7vUw+2fxYPhZPh3S1JlM+P8vBt3hkmVMob6c
EgxdidBso7t1qgMn+6LlZibRum2KRujPFzhdzoUH+nfLcX3+GgyCfvIrh0B7Uh5D
eTLl46vTbYm3ygh+7boMvq23en7ft9XIbD6Hb42OmV1UZoxcWI0394KK5G9fAAYz
6PDQEFhUx7lUrjOjYrx4uKBt+I7OIkOu7iBYFbJR9EtQOT3xBC93M3sbBmTsuto+
1jCoq1KUcAHYsgDA9qmdzbhhQb8KDvNN00AuQjNcblN9JnFdbH953gw2QcTtZF1g
BbxlHmvwR03yn+5ATeMoRR65kizc4eVP5tS1IU7VsBveim0Hdx1MUrxOJE2zRsKS
L5fE3c+paYjoVJ7kwkgc5fDf0nT7NhfPwO4wBLjSuMmeuWVbH+W4SvySXMaOxL6j
lpmlBmx1AaxlhtxDI1woagMEcc/E/MxAjLnhrRYRXsCb1kU0hRAqhUfMuF9ccn9y
WvaX+T47b9s8PBwBznqktI2IJ8GWrNoxZ/OEkGbhyw5b28yZVf8PREJhZFao5yUz
T0lBa1LEU2+ZF0du6ATD8sv81vgnGYMZ/fSHGlGTpsYaUXgKpV5t3XXT6zR/qxxB
7658ns8DA4Jv8LZ13V+Jr/aGcl3JSVkLDC5n9LdGqfiTTNtbwcgTtptdZ2N3ycw7
oqNk2sAajXXlnx5ws0O+zRg7QQ/A87j+CbkYkfUHsCBAN2x6xc4IQAHuXTijOCok
6HGnc19GtN8gTORXFpdKTooRjdABaEAU3ZW726XWobF+PKLytaP/ixGWLai7s8zQ
v+JpPvW/h/PX13yvbPMvxy9h6/0ab6kqT7bcQH2tnSUK8Zd4bvWxDAUINx2tyHgR
3h/s17ffhpZlp7YXRKZKg6IJbbfdqTO3rAlyua8E0cq++KPufYTmZHZ+YZV7LjHg
RJOpP4ZzPTVMHLYK2C2ie2fIW0tKYG/oL5p/h/1XuVjcZOo0D3fSJL6IQ4Ic5tKg
8MALfDyYUwD75k58HcR3sUAHqYbZMe4RZmKXOsMGCec688veESm1tvY1lFELMnhB
+uLJpPaHmEXipD/rWfM9ZSNn9ClltOigTC4W04ua/DQ4L4Mb0je7XabDAyhwah9h
Dm+YuB3U91d8DT92dUpAwRYW+5/4EFY/eCkkNfiu3PzzLW/TFa35flaWzjV5kiX9
R0HcS0buhNbAwhfsJGIn/1gw5JrmwIEwR6dH2tQT7u3+EK1zgtj3OTBCIfZzOJcF
+3JW5nTJM4fnTUkbFGjWAFSmjDvSs6R5onvUOEOPbNCjHmZYP38LKiRD1FWWkbxc
SvQSpClThBsAPyoGkdj8dltlHK6fTgaHOBkbYcwl1tC7+6fcXzhgjycEICqAOtb4
XlkyxQFxr8YF5W5KWW51xZDdzX9cdSa90MVIBqAlb081jDOuEu8sX0xVgx0RwauQ
JIytMTTNVYIdqAAKx6Z05Dz/OVM+MN2lcwXwKyt+eH23pVRLNJuyXOM8FjB65Ryu
d/kOZ1neBLbKZlhHxRmxZy2dBMoN9ma4hBa2vgfOpCqiHS1Ztib5CInGkwcJiNjI
xvTsPUnLVzVGrYTIK12PzHSXJ0n15h8U214btFfQRo8kBagG3uB0cPSuQIWfdvDx
r0d23Tonprf/jIzTlHrGiH60uLbbZw3JXuG+Csnu171hNTa3Vmzaf8aevxz/SQrq
/RhUuPHDCF8/JZSCRNJoLFIQ5xg9OKEP/eKEep2hK581IusyJy4GPuEJ8PB44goU
Fx0zss0S5huY46fBktPB8B3e1pS9oUZzWfszh83miL5LsQcAe/X68Wr4MHetrkBq
smhGsB7CNwQnA1UB4v+rkt2zPL7pgZdQLh4L8S8ZqJdsQqRbmDGdgwJV6koTCXP8
n9pN+FZFlvUrir0Enyt0J3dspjzVhf4XrkrjN8A2MXWXR/2omil+1IgMB5fe6Pqr
arIP5CkFiBrqerRV/CEX8rmgpfljByLXx1Ohq3mtGGNsJ3z+hYrt+Ng2YjcXSCqn
xobBE/rOinUHr+jTYR5UpisrzycdGGthMGEEzD/h7nO6SQGg0caC+L8HoMlD07Wc
Z4zPI472rUKoLUtv5+96Q19nOrKleQ9P3LV1yPs/gTYy1jSykt0Euv3fofVmEBlE
Uh8R3zwaFSc02pLaFbTqmQx3k+adBdFVIXNrez4wL20IGNDCNlZJjXId5rZUnINq
fK5g29jcc5Tc2O1on7onPt17o3AJVJuJjp2hSyDcEa6NmIzLvyqYIYy2XXJw+D3+
BuxyAOKc2t5JtecqkISgSwuPeTpKZYzleHPrLET/1QOlZkQ/BPx9aXiqmEauJCw9
WLRPVyyXTLf7dRGyulvHrvYhU/9Bz/zmPnWhb3m3N5X4U4TV4zK3Hc5XehwJ0hdr
2zyEGPBE5rfajJ/08PPe5HzyE78xpBVuo4LNuQwolegElA0+U8hY4X6hn/wvP9nw
7SivQRVsPz3qMhS+Y5dLf24x2AwU6aKigku9wICFf6620uSE4oyw1KQ0D/ywZlZa
zzc4+rTKRsrrZCP0S4xnZZtvpyqn0rdf8Fcf7Ir7Zk3e2HvHKWKmpwpDc8vzR8Li
BHaQAsS2Sk6xBv2QJdlTEhnbNm4vROkM5nntCuQ25GmOgRVwkmgveD4ua3cGU/Dg
RrQ9mx140RyQ4Dc3GjbHUWiPy7E78fyCwY7E0LIa+6j1HIykM5ELtzjiOihElsTg
FWo1MtjrJCNjgsVcXVgylmfsu5GnMytxnJ9TJrTLD9urVGAJ+WH3PbtqDg9DxGqd
hGDkw4iqye3u3q+ANSOSm/Plv0sanoWHFRLEynZj0LMO5NZydSm2aOLRENB12Lqm
cpUGPCahI3A0FhMrvsHN/ow3CCyrheTzvOANxSSGVvbvW4ogZdT6bMCnEZO/2LQ9
mY0TN91+7hGSqpTzLfH/ybmpDA4YfrDfbQUhSF1g0rcPF9Hyxo3cnXFPXKuNQGD9
/n2j5e2aDX/x2to822NTIF/ZRv0buxVo3k9x/z2xi0hBBnJW03dZbdCb+4yT6NO5
Kr9uztHZAOrzTzwDDKdJj+Zk7WvGeoDoMsntpR/16fYf+8bpe6ikFJWgjx/sXlyz
T2QD4YBZpa9bBMIq/Y1wGmqPVW6oUvJKM/oK6QlRFB49BJjlz1RGE5hOkY6WQW9v
fPJGOtzK+1Lt6rGCnpXf4V2/VXPa1Drsq8fX20C8IUfe2IsY8XDetF4EGryw3ixB
enTBAT93HlzA16g3jlZcp+Tk7L+Hr5V12iVJVk2dfPw78OjXDuB/Gw4YzMMt3pCW
pws7WXLwkaMG9IK9FZosRPCSUY3rJwifB0BXnAD3osHF1aIs9S+AO0piqRPaPICT
ZjlfOOOi78F4S82EdpzXeAzzymxlRItPJn4XpIXH1FbzIltRi/vlKe0iQ8T2Z9rM
k1fryNdoTvF27bj7RrXeAxoqiRTzbSSBpprxLAJACrquMceZvzsEBeZlWrYGDMDD
NNBizkg8RG1fm1toFbTUXAV4EFeqP9bNLHjWc1tpW4H4SGWgmFO+zpExGhmOykKI
tEgtj43zTIlj7GyKyyBUloAdq/XTbcowQhbtZg00TMt4upYxjzJtaYXiZ1S31MA0
cLFnv3VkVVhNRRhE01C4XuhUjjzcCpCSx6MWBuMIhke8IKfSg2RZE/AdE814R8l7
sIRNq4k0tpT73jyzW3c/J5FnrheKJd3y8bruP2CPnm+woQ6nyltcggFVCerDCuCi
qqbAkMbIq0x6PMyPhlilPl5MA0xoiagfi7YT9qBmGMNlZe+XF8rczSSewB3YAfi8
M7+vMIhaYRJSmuRWSA5ct7eBelBvsDEJLwbtZMikeXFFzCOm6LqgDqQLvcrMwv9g
CqjNIkkeDobJqWfuTXIO9HS85HkmomQZqzqcyIEfwVyu3D6Hx8j6iosVqzPj6md7
cBaMF/xDLpX8FF9+7AMcIaAnINOssD9eDWmW+OmvVpfViFSvKsGicjNpv7NGjOjk
YumT664ywhx6sXSJ3yE/SRm7BuVfVWdQB7i9KYmaSUZAPOnbEWG4d90WZf8JsE0U
nKPRmlm908NOcNdvoZAv1DtHGXxvF6qQ/PALaUS9JkdyPvwv3qWUK4Y2IKqSiLLO
7/vI30AwcxFTWFCsgEuigbiF3uHzsts7Z6Y1Na6TLlqdpfS2ZYMUhK8wIiAMI2mB
/1LanwSacwQtygRIbrlzhhMLd64aoV7Fi/1FYe3tGv+oEJhC0qnttImezSlCs9Xp
dqVuVTUYSkku+jbNQyZkO8g3EEre1eEM8eYiBhmXYUxeskZFpML5p/AU+a3OF3fG
3NyCTZAm4rfOPqwHn/9om9JyfeZ2S2rNaw9h+ot4Et5DIIG7UEHVgSDvQyp+vXMa
bbfjfcodCFtuFEroB+mal+gbik+g4bSGIpZ1aL+S5gtWcBUrsfdNbxQVVfa3icS6
mblH5LrPCQgrXYRI3pFRllrzhxZHJOR56+cfHB9Y/73qlNe/rdkZb20az/CrmSqw
TM0k9tB6yI8RXMg1CjhKnKrqxMz8N7fO4OXvnCIeYQieGLXrNRsD37OS42NTKI1e
dl7iW6udK9JGmEF9L5sjniyTHjZioELrZ2F6t3ELDVwiMtyJiNTZp0WP6YTAexpX
imJxiH5r1Qkzw9rSFK4kYJ2M90IxcEyqQ/NH93MMKfrDWVRtf+Bfpf9haleFwKmS
v7XdAYLnlhUYDEZkp+OsbWkgv634vhPysGdXej+UPBcq+d8Un5Os5L+Ph7X3JAVh
bQ9DGLwQ6WN7gE0KJdqQoVa1CryPweZUZIHMN1BwkCghPfRx0GZNtzjRZZovHEk8
tPuZnFC3I/SLHDOFTLPtTSpeIatAGeuSW0z/AisytH9EZVHPoAKb5Wfa6bcIJxS8
MRkJXsg9VttR9oTKGNnno/B8FPoKND6uPfe+uJMmpaUoYszOAH2NAMYrkn/TI5W5
EUNx0hfDBXE2TVxJBIKk8XYf/PyEGcHq4coKetfRsKdku6VHFa6YEEHuHiI8LU8g
9qx6GELM8SvEfoCG26cDS+UBgcNHCJ4G1Ou86YYM7yr/e+sGKz9Y27trTksJSN8e
HbhgH+L6F8GxWIbkG/z6zkg4+4ULJVGkoWk64DALdqVRlSNEPEgB+PnULzVtv8S0
yeGs656CVcJCsHqKxUCd58lLGWGK4VZ/bmE0FdAkbcvWZRe54intjCDuAZU2WMUK
acnBWxZU/kKc98urYfjjGt0rMOdoN0euR0KMSFQXkA10SHKM2dI8WqM2K7wup5dR
E28DxZ+ZUxSRM4YdEuwie0V4Tqhy4uBfe12Dm3X0H2fm041B25w54zTn13m/tcXH
FNxArlu6yVJjwKOPy+ZYpEQz7pBnGElQQxT8jh8rf/KhqKFk5hXO90fs9MF+rO+F
rkPwAUxyODR1UQAy0yu/fgu0z2U4byZhz1rs22VB0786WkspHh7+bZA5rAyCKOBu
99j6nfXw3Bq5GfXbowX5im4vAdLDYtQSIkQN83XH5qBVmtTTuBx2nqaQip8WNdAF
Fp7dgARyJsWRUC3wq2BZI3MP3xOWFj0lHIa63ZroqeZ3fLkGhJpsdZmZyF4UQPD3
7V6ZAHu7AzSomeOnER2v8NAUL2N3KDghSeZTIXx1uhx6zK/2iExyNWfONe9zKYuM
36c4FPsa4ulS9WQxfzjXXQyWOC3d+pceF10V5vWOkiDGpQYWGUetA57uUKCW+wsQ
Xcs3eoziQRXy5aoY3EilsqfSMQYI9q0yXE5+oSGcWnTsp16cWpjkMqvr8okAQ5Va
zyuFMZtTd5hsrh85xBZe1y5s/0VI1er86ZH2f/S9HAPxfJtC8ZNF+LwrwPWVwBi6
hjmQ8YW+hHizGnbUxQ4a4k4EXECkiAtyTc7Gqe/B/sZ8EaGVt+StvRHjE/G3kT4+
uhUOeei+i6A9zDGW+oN5eNXiZcfoVhcAnJQ9PlQGOhW8kavQ6siWr4qzU07/E5D8
VrQ/ZrDqrMsFwaZjaDdVR5cI6dnZc3ZzZm/0a4BjkYJ6PGL24H5WSCcqRqKeHCyM
ucoJoQjfUsukUgPFizzNl3IwjmHyh2Y+uhZxPV5uhmAhwVRWWVXFmrQH6g+db0oG
iRjosueXiHGseD/mBftDG/WBuWVoWaItb2rVXzg1CpefN+rKTpNgAfoTAEQFRiLE
n+LJWcR7VEbMkhi64YVqOnFvG3nfS8edniSWLC87SU07LKaw/W22+QfqwBHF61am
wg7B5uZd0JH3myr20gdSXDRwsBvYnwEtr4+pg2R6ErNkpsnGrf/Q7BvtmAjKe/Tg
PGNJC8c2BSXCs5v4R8OSdkWsc/nTNg6VdhlRCTOKq4HnKMzdpGnT1wkbA67rJrzw
UeaI/yXpeIF4GrKk8C9BgZZUA8V/7yVPAs7d/6G4h7hcspWor8JO1jppjssam50Y
AaK1gYOsNdYd0xsKdnGQO7CAl4wSoeLnorTWFYhv28h0e/ILkRNwcECyByhpq4D0
tBPxDEpXHrjnR3wnd5OWy1qqfdw+6SQtiwUOn9QnAyCk0ahloLrHbKKMyRfYlymU
26+UjV4/ZHfEEzk5XIiQB59kDy7DMURmmyoAgIReoz48Q3l6BXKtw6uxR0EIDp51
8SNepXbjadOU6BDpFPu4V1D/2aZjtLY/zSweQGl5CqhHcs2Blm40fNmVawGkJiZR
MOZG9hVLOuxmrT1v5sfhiJvsfYMVYNMrqtSr4ggObe5w3PYTzHPAH3lTwwtAdZ6M
F3XimBp+TWlR2TIlh7+ncotRd0gyN7hROngBb963Obk7/mA9IO1P3MAb3jQVa2a6
tncjGAMpBGzKTEjTebiPWGkDHktwZtXe0VGsz+kAIZGsIGse8hWxWQ+0FzMlVzlw
tkeqb4JSD3la+43ji/DRB4OESolzFeiT1T3+8Fo0DoqJK6s29YdepypdkRuAB5Tr
51NuZNZ5Nv5SMSf6P5I/tP+sflQOoQTXWxpzgf3F+2tcyKy0I9bkJzfBJnaQ7se9
Omq+vBWAaYwuoh48KIYRnoYKCUtITe/SoEs26fxV3poHyNjpemYCEiKputv4H4YQ
8ix0ymRm4xaiyKmAlXIl4PXgFSs5121KumTVtTP+aNkxVqA87vlCTn2429QeYgVa
O8CppB0Toty/CCIG3ZzuPmZZsAjDBxPl9szbiU3d6EQ5Kcq0t8+660uii8RMAaaD
cdIbp8ZUq0dkv6QdLx93lUJAPtrQfEukHNfy+Kr8nCWopNYa6k89AVczYsJlXM1Q
EGDfm5ZziKQrks/V4PF7Vp64Ls1Pgb0gLpMY2+9zl+48BPTvnow5NszH209djW2K
65j7dx0p2+OAv3PKu4+kFdTZW+qsQNlGZFfR4ejFMEsQJDISdaPBlTziyBMcIU1Y
62iUAWU9//itMUoA+q7nTuy5y2Wi13prfjQCVBVgLjcoMTN94VAEm8O5n5y40u5+
S46iqMVmtgy1uW4uCYSktb+LgLy8N65L+gW+t4J0aBQfFzlmnKnQ2pt5ByZSYoLp
jZE+DqH+SqxQdCfnCVPV0sVOsPn+tPQvCa4EoHgjmltvUA4RafYigXyHmMvHWW0C
wVWhZNbQ5xOkK9+4N9GmPtowk8mSi57Z2otU19ymQMy2aO6DeXr4ElUq61mI6ud6
kAysPajIE+vh+WCQXOdGqrLoyNW0oiAJI6LpvT3an7Ri39JAfTXtqkMYDpPYEfOU
i1KLaajnq4T71DlZcVlbqahoOcI7OlpRrom44VcOrz6yhn7IV6fdXmRWADYhonku
G6pfmEUQVdP2f0RxropDqeeWyytK5BiSJHw0HbiAI9UDLkb0xxTk9j+0nlurhuoF
gt/ZCqys1Kkjy7ELuF1TAbLpT9GZY1trUTJzKlsqm8rP9YlQ658orSvZXsCdMUPs
v5uvirsJuXRzhtQtvO4OxS92t33HM2LL3DQb7pUHlvUCJGKBp46kyOfqeguZ9Ff6
Pljg/sJ4HoaITJyPWawH05EU/hZRdolDBdXlB0gnl32mbYoGmwAIk68rM/71+fHr
11eZn/wg1jkUgcuL/gE2IoI+n2FFna8NCQyTW+6AZ+/gAeN9iFb7yROtQq5MLS54
ahtFPbqlNdqudl2ZvKZAY9jOS4TWxkkO6b82etFRB7skejFmD8x+4IBL1Na6e8Zf
xt9I2WlwWRIxC+wfZxP6t9jc3lM/dnDezBMAqgZ2tiWzDT3BUA64pDsfFDnHDzIe
eNJlcBcJv+fGCuKI/S7UAMSOcNikSSqwW/VGbT2Ar1ZfPEBRhilUV7+mjq361XeI
6AnoaNibsAxoRBqu0h2ab/j9qjExVQcXgFHPGgS1Vob+y86kvikuiYJjBdvKXk1M
/4dU9K9uesJ0yEFR+ZH4/1yZiHhSuVagNXc9+Q6KA0QHd+t2fsxQ505N6l9Kt9wf
gy869a4jAHnRED4g2gSkGqv984Nnlt3D43fO6FbJ7VSq93Y0UZaAN6QJcuRx2CCA
Emlobh8rCXrX1En71KlfBD1m2+IMQGhB5NtUsGzn2mwoj1qqo6Z4t2Nf+x90SkGw
ob60UTZD1OP5SaguGhVa6wJfjoWkSkWQu9m+/YczUqMJob4R6lnbPs67s7tOqVFG
0HgPNSadpNOUY+Yboetz72YpVOtGLOwaO6HrOnl4jLvIepGnoXdCcfP6Sh1QsokZ
wYWknz0zt6NIPSOmdv3NKlym9nHNmxes149MclYMWUlnTpQmUAVYBDFuU7bAH2Wg
SCNl1NbkacVPH5ReBu6YA3liykgPbRyPdVscMMfKxvumVaGgzkxORtcuI/z6rd17
GI7xy1d2CvtIdG5vNBiGpRVAqolY3i3FIS7peJr93uYLGxlMEr0vEf2wRoksYVge
JnryQnGsE+TDEpNIJ5RxnuzTzD6O65PcEDXgiYx3nsekJGSNkOa8WGEyQUx+KvHo
0yaHOgxINIuiMeJ6c90BxocpQhbxwzlbyYJtgxzOxZGsorsWHYiUvjSc5Yn8kHfp
jf8zocWvm7AJMcPZi4A6rio1ptCjRfEpyxFIwtvtO8kNBqpq/Q9xMvfLf9gkDRCp
2lrpLys77RyijFou6LbONnC1Fcp51U9sLrG5hoyEwUgCoKa5kwLb06PpZ27lIjbl
6Us0SAZ5FRQDXD3VO2DNpwtIzQjlRHECoLoT+eZoijh2MM3qLEhyj9jmu+RmH9UM
wDSaAfXYrem+uua293lni4wL9VDDxJsVLWuSWlXsvSsJ/VYBrbU3TV2HDAdZ+PXk
2RPZkYH3Nyf/ZAtTW2bqeY/QDjTh5O6iazVQ/HbW5Nnv01/qPiS4cVOgVHufwCyE
5n5ItxDEYv5RTlsScPOAx1tmek7CGosH7owaCgm0tjLikDMd/Y7hwsNPjxUJ+12i
Mmgvq8pdaXJDWptmcztJ8LLRWRPzX7KrvbRjqgW1jYqBLYY0GgGkvZcllABQEK7G
xBFFKfK7z6yVeSaXCZkPZUI4t0rRm3Tz88JNFih8ep7dJwuenK0FQ1eDM8q4A3Mp
XVWyCWjM5Wfeuc5Na1qK5failaY8nP4FG1wNJs72mWxa6+4tMqZyoGbjbbv6pcTa
HgXEKd9WHwjXdC4f8xETKhOwk3BSvu90CRff9Axgwe8+mByOVfBayFw7muTaZmRD
X1Yss7wWr8nROF8LYeuq/gi8amxTVL3kZLzALN3AcPyDeVkXNkj/gXvyHRBNXjB/
/oLFRriwETTH+yNQpVH4WygI7cehMp7+R67qR5kCZdufSFzuTwmVjvesSpFkB6TP
FMiMXyxUANkPcHXYyK588K4+sMVpgVfEzpmixJyVRQY7HYGRqcAVVRGkkrlVyGcN
PbUhzJYC8rqI79KypZSUKJEB4aAfrlF1EnpZdIBixHMNMId/qcpJv9FqBH80IT7E
VMBi5XE9nUnzEMSWkGet3bdo0qqliVHzYn2o0hOdfUHLJwZnmoBVlKKuV2cw6H8W
eyu/swOeULT3Y0q6HQhnFYzBlcusEXt8/dbxWYkk/vXNKn6J+fgqrCRUbrnU75i2
KcYgSa2bq4yfFpuxu5DevZJ0mrdCN9orWRLoZWKZGEAyKt2/Fx+kohfMd9JYJAUH
hmoiYVzbDJ2XIHrPpGrqZHgQe/ZkzE+e6LgZeQYXjTN9pjskr55NvQZynIXRSluZ
s3prMtdtrfypMUidCZ8nbXfF7MdbT4eirwt49HWZ2fUn94ou8ZPHqiYN/zyLRp+k
QgO5AabWKbjH5P5p4nWCExovM7g7b/wcSvG8rJ2SLjs/VLY/lhs7RG6wIbqjw39z
ss6RvlyjoiTUPz0CQvQZm5BkNH4KWvvlpwk6Y9mXYDWV2WIR8UGthVvQAEBR2Tke
VCxurNH0VbGNmzzbQEvGz6i5tTF94Xb81qQbFckOMuIUXcTbHY5B0W92PwziRfNV
vgqu1RNOtn43jewq0OTJ9NBb/Fuo2Vru4sVUv8q1gPnU19v++jHMNKyKL47S9Ror
D7VTVr0FUwAU5EQDsP3c9W5cYHJFUpqID9b59x2eiM9R7KxjNx9lrmAcUAsJPgBN
0osXevLXYRWKqeGr7I1+HUbKUkPLPzPPfk5G04oxDIQhOwJEpJb9/67iUp3ylmdP
BM+nrQWf8sQ7yUO1CZDB7fZ6N2VgnCC6wKmKn6hE8Okvi3dfVic6rh7IXTP5FiYv
3GemrMZ/XIgFC4LR+4a6Cdc0TWfp1H6v0uz/rn+zYK2yggdlsamVFSpX7kQKBARX
jCePRGNcJ+xDChS957lY11asMdW/2gWnv9QB30OGw9KBF2FaG8vnUG0LP8IKKcY9
vrgLkFRIOWYMACI/Df8Zo+BmtahnoZytuZivI8QGG0eqsQi63DzRB1MHMUJ5Y/Wu
X4uzsg+Lyq2Sq3aoFh9LHb8N/jx8t3AVHTOEKcMb4w0E1K0EoS9aXowOhVodu1ud
N2nWWxdxd1SOd50wC1G/pzZpd2QHbBo3zD/0I0qRb3+8JUP5tqR3d00zamGSpLu+
tajjDUKO3CNwaV+aAVQftX7oSzJgONm6dwein2N87eaByBkGVU4z4Hnq2XejKXpe
k5J/Q926/ZDDZoaR7lNETb6BsGU5FNJ+Cdf2Vp1/fKy/Oi01F01N5NkN2ZC94JNI
Rdo8ykGR4A4BWOas1GApNkrbYFr0Abq/RevK1hlV+0l179NHpfG9ZOsjp0Va+zzN
ZzKEFbPSmaxBPI90mDawry+RvZcI8s8+BA+Y9x4zxANWItu+MMQCsLVTQ/N0q7vH
uMoL4zOxyakYG9YQEc0AzXmwyaVuIATQQQUmUxMRzODAfNTGQ6N3pqiT/AnMkHml
7+yfggp/+0TSoDcIS//s6iQ7xRNBiHW4gA1CkM6A3guXB7sG3G5tBP1tVhGseI3o
oneAOaf2qYyxX3i7h9wqZrpZa98Q/ATyiaTIek4YKkGFnqMSsqD1pWY+BqzwkWEo
ZZVQadp2kS9JVdKcWxRqSn0RWj1J1V4bhEMu5W8t9aHwY9uKIJ5Jhc2NWIclyrKw
fin9w/ZOieVgw2gzRKpp+ulSlxJ7EZtzKNobYdjo8m49e/mTtjfjGGCC5HEARYCe
z2dw9S0ElgpU6/JDautoQqn1+VyWEx2JdOSqcsXyMeZJleRLsjgvKojQDfi1sTIy
+kLvrfUuVulYZJn5hq5fGjlEXXhbnZLhSczGFPEvcqaeKC132PZ5bWp9tWn/0Z2J
Mn0VMgCyOtf7H36945qcXf/e9aOi6HEFR+J8HaQGurkXFcgs7NcgF8WLbLH5pwPc
i2DwWlhNjZ6bSHg1WQ8W8z9Y52v4LmmFSRB5r2Z0iRZan8QXorjoYAb/vVNlT5VY
Rb0Ks3VHLQRQSXm/K8gKaCM64EUmnDeNbHlG0M2pW1BuGi+QUqepfLFU0qJOlUkT
iO9lrj+bXzwEJ45YX1aA+L0RMn/cnyz/vAtPt7L5GdBYQ/EKa1L1QksMV0a4iZsd
A+TY79yOotu/aiKJA9Zfye5xYgRkvdgbRgpjeN7kfZ3uBoDYUaL83AsM/m38/9BW
NEHc5KJA+bNlPM2ZVHJeRz6VoOyiFMw15f+VOXaq68NRXdGEEl7iWMuOJBOt2vB+
MuglrS/ZyE9L/yZolTsaU4CJmvvYm8bEaKMDEJMRvdTaLajBgQfcn5yyS5vb9O8S
wKOfNvM68yPTn3qKwcj5BLDC7glkWF5f39hkZWh0ktNlnvljcXRwlESSjUjo/6Ue
6pZm98W8eYWI2yQKjQIkeECd1UMmjecpuKTm6fuEqA5rCyYeeX9I8GRxmVv5kMmU
Xz7FvQkd/5IQq1ZK9VGg5xPnDAoF00GzsrRa3Qb7QHmj7Newa6QHRqnjBZKUkrhq
Giv24ovNFIzq9Ra8RWDi9v+l8J/IhWBTVEZQzeNa5LZDe0GaPn9+QeRqZX0fGi+A
eOaWYpocOW2++YUt5ZZPj+LvRkn7oNQpS3v9nQut/GfbGFq2oJYLuBUIX+atQ5cJ
mnHFsZtsx7BCLM8A8xl0RR3TxyK/bL9lXX1C9mSPmH4NWyCgjCneunIGLiCk8YOT
haXrmLFBD2gaKOdsN5zGOPmhQ3XZgAEER+DOzXmCEfpmx9NDtBZiBcO18rhZMcwq
VUkKDOtlkvqTBHaYvzF5pwxO+EqvDRfad03OnbXZ6Oj6mNCi23zOfInR0gY9uBwC
xpprFV7K+VYcd+WzVh8aIG+3VyHC4D/N3yxOO4o2f8K+LUpTdOQpuPMs8MMeEnd2
P1LoQZFL3U/b/RZehITBy76yr3UGAULA8o8ccxbroiiK5lEmDLfqDogjlgdpM9cw
yHe/kI3ucm+B/EKcWEMV9BJP7AyVlkoXNwmagl9CVFY9AFtoNXGyr8qrjeP3hGXz
8FtbUKSArcmeNPPE0N9aclzd6PdolptEqqZNsEWPnJtrTCQCh/Jdyiw1+6Pr1u8J
DvRLumzsNYv5atu0+zXSdEcXmZuyhFMxaHnQ1aGod62VYsk51VEuLBHHmoOn2jrC
BMy42Y9yT3Ylun9dnqH5Lrfr7zLcoeUeH8lXF/WWnMA/MuUHM1/8N5N85dXzTHlO
4ENbswfsBwmR4eqAhOcea2y/ZcjXVJAzUo/+1nC5ikir2qecBjC5ty98GyEeeQ76
IsuReFF/YK9tgiYwHhEq3OmUrhbP/+MyTtk+qyWMX4JPnZpum1qCaVkfRf1O7gAn
fDZPtbIv+5VMi9+XT+7yk/Nc3IaL6nYvAempi9zq8Jp/J1mngKh1lrHUcgWhN1+K
43RsWXSIZwqT7UII4LzsTCY0ZXB5gyjhA1LX1GTdpck0nzTt6IIx7hsvOLrNRvKZ
Rc8ddBEVhM2yiL542+THeM+p1dquziURD1RIBmrd9ePfRWzs5HrYLAg7CjtiMzsB
CgqjBZ1EeXdtt9NbkhbJUj4U6VJprhReMu/bOd2fC5DoXCghaZtYRsQ3SuO2MBkG
FljkLdVHG6bM4yXcf3NFwLRx/BdgAtRsIqECue4GohDDSj8zsZwBUqw2cG6sJ1V+
TLvIOh5BzlDKCMsNvAfuVC//k1hUAv2I8jZWbx+ZXl8v8BgDQoAs/9r1OQCA44a6
iFLay9oEkmDYiX0qiyn0s62Oto7DWpEtmow4UNkAdQc3UhoYU3adk0EbRsTVPYgh
HiT0IMZLFuK1z1k5zi5EqlIvl+Xl4DjyObyPt/zoaPKRlqGYJ1ZkdWe40Vce7Muj
r8VVlJxxqI2OOFEbRV1lFfa3ZyR6Brr4AqyaUvHJMgxDok/twobPfYCWRSwqjzbH
mISjdcBJrFxhOhBiXqj/16ZFwEzVOGO7oAQjJDPkbOlbQMxb0k4Z0OAGhDAMOYmQ
LbxmqI0v2yxIPM4287d/CgsA+0zdMgezh6R6Kk8Ni/ZFmee2w07ukCsean37WVT/
DpEwunKVwvUpVCyr4gz0heyF6r9m9k3aRx9nI88m9NJWVtRQTYmBZDqnJPAKRa48
FheMrmASS4ctT7gMEGOOTFG8XWTmh5fJeNshtAQ/xLzRTqeNoLgSYZqjlNX7i2JV
cTlK6B7bkOPb3Uea7uBVnB8s++YzROIVP8/+oDQgn5p2TH1Jgqg9qJ1W/xedtb+v
JmT4qzCJ4T5N54hgGIHsmij+MhIeT3Q0A9FuI4dg5ihFpYQu6k2DHl36Pvj85kPd
/wUiecs9Y0ClrwKg+ryNhlyXAvOnnr9gNH3sRAKMqCZg+BleluXMbpx/SVg3hdOP
2FPOLXlwaDwjFqrp0Zo9cFmuN5v9dWdQN0AQhLeCJZvTIHlqJhdc0mq7ENcOXzY2
lJxYvUX7V4ZwAJoj6l9+D/2/aiQw6wnsaWZjHYFMMpBgAbOFFbiR1a0T9Kbd+5cj
aVTudiFFmvKMYTOLRKKDj495Doo7DpjR0NRcxaK3wCcBUgaBXRubhgE4WLZXnA7H
msyYJ/ZBvubvPDkyfgTXtPFw1TC/mDwUkipE1WI/RuumtnP++JLxw48ckJMI4IHs
CqV/0C7/6+LXLCf7lls8YnttYd6tmZvyGPTdnVOt+iK5P4zKo/VvrZ9tdrucphuh
kMBWg+leoLAVSfPuxd+veQXzm9fJ4For+zDbFG0uWYzgxIrP8BcHgDiygGgpMjnF
8THdceF/kHY41NXWVp04sNlzpgfjmV8EQXjF2Pdk16mwxTuZAopl0D0oEjdeRZ6O
Sdp4lxslTQJdjBhcPiVPCi12qJtvnYH05cQ9WT3svb7/U788/mFsf42FYf7eGTjB
bkJ6lnuGZxWNhNg6OMmFu3/8MCebjyUCCjkjOHzQACFQyjAowjjWq/vGqLspFXzN
5SlymIJIkhaTvdFdWmlQQHp3ScUUiD6Dp1jUc1XbtXuE+VqkqM3+OnBfpy8LoXrz
1luLIh2mXkOiAE0hD4msI9Onk2unTsa4ITabWhjrBOtCNcBsBOjt5gBYQhiVsqyY
Opr5wpmA7cJ4cVhu77ACnQO5SGUpcK/o++AcrB60TX5QDyDef4uTqMN4oG5B3zw4
9DPMyRYzCOFqp+8LKa2SP56UL1upyWJ50PVEI8o1ElpsNLyudlBkmVE+ES1Oia3O
uVHyyqpg2tbMSiEf2Pvb/mn4xs3Qp6csSnAjrtSBWBbZGCiyWChwOV34LaGDv4YK
4EEzUOQOxP5+c9otUXFZrqOE5SFvasWnd6IR/+uJ0TZp4wnKG/qLNFoZjODPL+/r
ViP93UMRwtWYC1GujRML3MxECsXjFoD3FGsLPkLTbBIVWX3gVpOHLkZU5DubMYaz
oBd5eKCLo3W28p5a6OCD0djl/Mz3R5ZwBnD6KTwPsa0v6z/yoYsRQBtMW8SLqPXl
y6sVtyX6e/uXPBqQPuCccEdnVTMxT5nAXt25+MXanveL9ARL+NJ97ncyAZNuoXyK
M6Uhw3c9CqUeksZ6ip4DOEGXT0QkYJlc4+uwVZiQWvesKbJPn33VugK+pU1r2bcy
excPIp1SfZm6gZMomkTmIiFEcvvS1QN1mNS7FZgl1SFdxpL8soO57JaVVQ4BBb30
/VKtl92J3oCkgp2FjXo1TEbNwfwl+s2zsmjPNANHZ/el6Z630m5yw3z2MT5SBG+e
t/bwqJc67rgy9d+1PKBSWLs9vwNbZb/0y+6VH2lucGevrhfTgi33lvQzpgOwOy8a
vjuS7jtIa30lIZW9Tecba+rqmtJAVR2LBWEfba4X5aEnfKnknwt/njhdkEEHNTGk
uXJHLVTBolmqSVelT+RxRm3p0OkZRVaL50tFQWQT5B/3qXWY7HVd26AawnKebEm6
oS/72mZkG6JdTzIV0hNPXqc7wRx0ncH2nU/faU2pTJyWI6U4ne535w3GNn8NOpfk
f6GW+q5T4bm6cUKe2n0AANWDIMmHxAWq2ta29W7IF1TjbnKL/0BpZxYLf1Wkf9Dr
NL+iTzicxcQWPsYG5EfMTluyAaZ30qalrbE4g7U0RCeuiGfURD1aSGizQ/0c5u9E
nJ11kfLI22XMYXnU61MV+Z7qtghYzbrrh/kiK5F5MvUINJ7brqvFKv6MD32LDXXi
rugGnJu5wnmomlRcXrZG/iK32cI4K3/IYIu57Dk8V04QwPRzNdu6qn0N0WdWq+Mk
G5WC3G54Wh0Flwf7iJGcVW5dzYBtBmVAyQ9g3hrZNNc39RR4KhMGjeYEAs25iaPk
tK0G27wzGRzy5a7OkZL2CKsLUfrq/vKoNNNrwv5Buys9QfKrXukov1KWJMMGMd6g
/h4fMB2zqp4pkXF2gY1FM5C7W1K96gtOD5p6PXYXsQ+sl00wdYUyS1c1vGfAyPKb
TVnfnFJbTc2nabNLJ0VHMfm4herZMYJ/SjXr99nG/0o6z5bgy8NH0nkWIL6O3eEq
0REhkQSGnV6rAL2227iX9fD9JdDWVomVOiZFS0cbyjIZEKj8B+Iqq8wlsWY2dwfA
bsoiH78sMQ3jG/9Pn2aklN4NtH7w7RTnnsrMwbsUIu7/UT0BvM1C3AcG73F4+1Y7
FmUMqqTcelLwRhWODUKFJSPgHtUVVEFtEaRn6VnygfG5sK9hAHa4IToipppsRHsa
odWS7RFRBewTSxNKmkMStO2trDGQ0GFZ5FViRXsDD/eDHHxPn3ZhD8dRs1zFHw9Y
Md9vwFNQbcEpjE9XANGCMAJQtg595WvL+d7uiR4yG1QcbgToKJ5qnNv7EMFef3P5
NLSQ1/G4anLgtp3phl/bpJeDmkIrl4pDUMKHDI0Lkab/RweZl9IhT02riSkf/JbE
whEwJjR6x9uHU0Ct7k5xuCtdlDVoD+rd/5TVokacGEjWEy43G1LZy9RCaDP/cObH
HxCToY4DEQgJ2DMnRavSjZh5i3SWbtl34sSLKcQRp4qgh2gAuNfp9DApqFQyfO2b
2SDhncpMFu4VCkViLB1LAx+2BGHWGL1Eg0ZBVgx0TisHvArgzf2xUSCklwnNcmgS
/xHT+rPW/fQDBLKZxub9ZMhPwcAXs4x3YtYuUbU3I7YY2BeIlFWE0BcX7CzGkzOW
e42KeBCeAhx8F++m6r+J/gJzPgPcYvSeb++qwq4sBr4ifABbT3b87PEytWTHxJIt
QworTt3IOTfBpuibkCHICbyqTDtvgYUe3uyBrnGQhLMoN4s6BEJZZJ6CUDYLPAwD
mi+MBjpcsUjKudeS3hec4c1XUxG4LM4pmnVddfyH2N3329ACq3n/ouGcrutPdgH1
QCcqFxAZXHLGob3JzZ4SrkmKmaQnk/sJ06erMVSISy1wvq2A1aZGAyBCSNFCviVO
DCwcUMuckyRbr912f/Qp6szOmCYie28a+L2WPDjNcp4N63u/k2vRXiy5nnkiExuT
Gh6CKIVODtglEmb9CZcRhjj0qjhlgBlFwQ2WrXgsrIeSoqH4QFGuNfbIEDU8BFUt
CqhbifIHJ2pC64FgFYCfdJ0wJz/UvsTXabawz/vOr4ZMT3Q0qpRpRtfZJ2pAnI0N
E59Ay+FnyYHjs0xeB1q0XCfTZtSGIMZAW577rtFgrQWDlRuN3vVZsS+2wb067we6
RZs3jCTMwbA4GAOCrwalexEfJsNms/1G/mcGmxKjkBCZ6WCjhhKKC4qLc8EulDXc
rdjLj9KyRPcpeqq9sC2uvlvG4jzrVAiQULhpQNgVOGGNTc/VXxeJwXcbWQFn9+fO
ybCGvTNUFmGTJomFHKgBCv15VQVf805eaPGI3dbkw05gKaRllLDAHfPPC79oZuRc
Rs9W9Du+F1AdPoLfq0dS1bRBEJcYYDXm3/K9wIOQhsAYF2eCFFyrRqd1lgA9MsrG
CL4QGJ7RBYXU+YdmnGhUy1DHPhMO8ow51rOJZc2+rPlDyn6wk9eUSYZX9T6Wu16F
K/vhFTzjO9WMiiQLEGpNIPPzsorJ4CR2hN2wyYVIYEizbsDz7BVgh/2IHS493UEM
wJKjb7MULOfpMcv8CEOel2p6QuF6HEYwfuPor3V8Z3MPNjTfTO4rhCSJz83IbGR2
vMWpJLwl/llh/RijvVLi+uHluSLCdjgxvJMXFfGcefDsD73uy4UvVr+MyBiYxlkH
c6EbQilk7uxgoTr7xfXZSE5n6AAX6C+A5Nsm9S+Q5wIYbuxwXGZ0+xx7klsYMvs0
PHxhHEVtSjU8X+s6Ln/eZxuDfU6+no3BpooqDEgJyujuO50aV1nlcRvh2IsiWI54
5+5qRh6u+5FPUSjL5puH8s/2/dWf02t7x2EWyD2lQOL+XTbS3uYmXrN8+xD5Zcmm
5i5vfxSWqeTxNaYlNW0Q/kYX7E5zOmQ4rha/FvebUVCsjD9+GT+r9yrWvOCN8bmC
aHEj5t2JAykm9niOCkAhU2LG+Gq+LyKL3b4TmvPAXYsp1ROKGJSR0mseEcLVgRig
z0JlDpNE3I6QMTatGoQusWMxMGtRHD2F6zeU+XJLIQ0zeIzco0hkfzrHPeNLhBWx
i3xzgPaRs/5T/+V62dMf9Fo+oGGGKxooykFx6ox7xyVr239rQax2SHnaZtidNJKM
hfBfqu81Iwlws9wWGovRUMSYCp9chBSCuhrmI0s6BNBK13SqBLvtDlHf4MB6SGaP
SewUU0XDAyyXr7LzKbSbsCT+MAuFCSMxnUG8dzfKBDY39QX5ztJZ0yt759qhEXSb
GywpJAL77mC73jk2dhnSII0r0JY3lt91519D6DqudwHT55TBDFrG0XZgdsXw1+6b
gDFj+4/nEmeOlyNWGV+Pwul4WvINiiAyBDtirLXxGZBlUdMSO/+qGAaUA3u5TwJZ
izVTo5B31Q3f3cRA5a5F/roaILrSHaGcrsu7Pi3LuAB2I1CzmWIOtrJ2V+XI0aOJ
J1N09ahmvhdQzA/QQAOBReRMSTvUup3pDJ2WDCGVKJy2qRFHoLRY59wUznUWWK2A
TvURzzDnkkMQWLrhj5NTZIrAP2c0pu8/ZVvII1WmS8fS/WC9zg4UXT1CCXOQ5hhr
DnfNkW62Hlm9SKd3WVZX3JNF9GjUzQy7JIz4sa7EQbx8CzERKadCousPd+HgofMh
0jFyC+3b0AOz9E/8FKc4P5cHfP6Y/r1tmKeIJYDrGgGYdJkBHRNOH+pFfk/4sXF6
NGADepAX2+nZCwhvDNagJc9FAQ/kmXJq8CPMThDuE7FK1iyr/TD3sNoBgHnTnoX3
XrRgVgEVBplKisKQavd7NAvsOK/rFA2xfrnPMj5fnyZGeRiihhGmFazrMfoJIBSU
L1vQPo/F3C3GZH4E00ltHd20QW8rki0p6QSrl4jCQJG2FP1ZVW44Jxq0J7JaB4hA
btxtLYNM1zYbWMzFrELsEyaxQo36xNzENSKuRDje/tmMoRMQQ+WqLIxJJYrZ7NnJ
lDJE0xCjq1/I5yvNlFzN6u6n/ZRqZpYEFxGDo4I0PXSqBYvcn9Ef1FP0qkarC1IU
nPXVIX98Q2tUVXbUIgSMNpTA7z+SgbSJVR2mJjUs2dj9c51na4arleJf0hoGQxXH
98UH3/aFnIYlhUFXIZtuFkMUBZJc7OxkdQCBBbu79JTVl5KXPLbe/vsp/5JBwD4H
kbCqqgXxeAVX56H6YVeiZ/c6PmyoO6Xq7D1MmtFAz8oaUkrmn7zAa5L8oj13Wywb
IzMZmqnVt/FdYSINjDQHZDgjWHa/Mn6SeAM9Yc4hmQxzOliaZGwT62R6IOVDBhCO
LpDWjHj4nnRub0J5x7cC8InJwLlfqqfL6sXAfNRaWd2ShNTxHcjK7YWcoq6k3cNt
fT1MLYzuiaAPeuU9BQevKAKJqZaXV3Ts2Tac+TwSvaslH0y1ML7385A5SHHFbNd5
et2nhuhSCp0+UYKWCG95FRqUbjnMv0hiq1i3GAYLXxE0sNoMHx+7EdhKUJfD8fB8
cjxxd4BGF/R5Wkg8OYHJS2StLg2JnIc+Gbu/6mpxud6UMEqHSrx7s3fVef+Bh6Uy
e3ftdcD3fAIF6FHXXygFa5hcJUIflkUEzbt7SbdwZux3mkikTlCTc80/s+sXHkFM
E7r5Vdpl8vhIrBetjV36ma9Jukmgg4+u2SXb8pE0rCKgoNUToCf54WCLdKb4Qw23
zkkw9aQYtaMGs5dZV1RvTNaOBthibzm3jQf3VrhzXEz15+pjgvoVyDcksWxhmZ24
pM08aG7UCdSj0F4x1oXonl2SzLi6BWgHGsDYOhmC1ocuKX4aALe+DJAZhJsh4QNZ
X2UTSoRmCuBcaN5JVU7B3AzsII1JYJIWgAhJUOe0doEgUKrQIODEQoGzbA0TMu1M
CSb8jk5rtVsj+zovSxoMs2cQVFRBWx1g5bMsCbyBzIlDyG40qhblQyRWzoTYHcAf
UzPWSU8PPKaGubwVjih98VX0ZrryFicOv2zj8t84gPrWAB5RrQPbuNPj9JDu/owa
EzoNPQHTwa0tWiuJcpjdodZxHUzyjIdtnfznypOD/QpflnesM0Ke2UhhKx95Lr7n
5+4H5KdfzsvGQnA6cJDuNGa0dMUJGSHtzxfh3i//F4j+Y54YeJQ7jfBE15qtkSPi
wUY3ZWz55dw6VW6RTCaVDMdBedkDDHwmIb5D0L26qmVAvwNNRqfO75bbxbhz8prH
gHx7o87lb2eE9foByXkWGmHWHTTHoFAfZzEghuzdkXW86N6qPZqLQ39zx20IeP7M
MU+NpFdimdONxxCwQjfU423saatelqayvxm1ghU3UGjPKap9vo400T8fKvPS+LQm
GNdKFxGg5RIzjYpE6LXKIrfom/sfQ0dnmX3fg+kEQ8mxBvok4ZP0w8EU23TppaA7
mzRE7rLp+SfknLigQgvlduW/6zNou7W4gp2pSfrORocYjhxtpOciP8gLfgaKhQC8
A25S7pLJb075ic2McMe+g/XlgKwfT8CQ26yRih0zuQFp5CrzBkLGuWUBRxZDDAg4
NkOIxi5fC84t+1sTKViV3m3C4/eMRX8JT6XK/7lkLK5dsXU6IfMVM4PYectXQIsS
RzS7SOdNXf+4OMvLwNZ+fFBWVVmtjGOfKg/HQVfs3AiklEsWt2uBtoYhQKcpbRzm
Lv1I8DD60ohzpKfOQTG7SoqzpXcNgl74+ziG6hKkU45fdiU7KrvUAxSu2xnf1GSc
p8xHNaXsejIeCOb1S5MFH7tUoj71fHN175mCUpGt/ZaRlGEXn45YaZSApTANit8l
U3NBqwJ3oSK54ZIuFrkxHG0/6hZo1ROLhyoUhyuVtIGQzMsjs0C94DhGQwRppI/5
GKeXH4waU5m3w3+Rrmg0uL3a3KSWNP4ZPnqOmVhiZvwir+RE+mDB1w/2mgLsTZKe
5gJ9FazOZVBjkrO3nubuQM0100t0IkOyyFGojdn8I0gG+XPv7caz84hsTBgUYTpt
CycyGgW2cKZ9lXDsulMntUheq+H0KKM0WvqRiPyX0fjK1UQKEPKwx3YGwjCr67yJ
2U7dS0PPU4+9tZex9mQ7edGgttsjp6WEiaHhpMHV1FSF7ZBgp0Z/KPABX+8oMtrQ
pkQ4PPOTi9mc3ZLGbwdGvgRJoUl8GDeEQUc1FCkxVqorumEdP/txdsyOYP0083MJ
xlQ8mkX/NFLjLS8KIOECdWYXFQrmH0lO9p1BZz3UDymfLaBAfDnFSzbxoCZif5IE
CTAd5Vn92tFwdGKslzQHOFqGF1WwBhgjl2qCbuOLz/Vwo3X1bFTljgryQbG3VLl7
XSW90YF+WyF8s09gcH9D2OeRhyOEhUswORX0YRcNU0BPPiFX3SyzPaXE6wEVHcRW
znm4GdZgsoDQfmeBsT4EdYS3kGhyqU2qMmJZ3K+bX3gp38Mq/5iFtyC+0avR7kEq
RjE981SpQNOyS1aGST2znWSk5yfzExrlaQ2uGikLyaRNuFVppiGPVoOFGAaM3zC6
Nqt+buEavzd2VUmb/Pxf+3vHuib4F6BMXGXKHtukBsfDjHd/HQ9p7qiAanYVSN1X
XU002JTVjKHiZH47U8J5icRlLoxFI9tc+4Uw1R4g96PHbD5MiFUtqR1I6J8ZqF9i
ngszroObQbe9wSJsVGzk0UWk20+f9acm2n2zBabNN5iwqPtvXQ9wOgfih9kgqNMe
K58vLXEsvz5ni+0OK7HCKm5kLF5lDs8DDZN/CDhHPdRpWweV78KsQVuvoLPQ1W9o
/gXrWy5YUCN1vYGh8MRMa5kZh+NPgeSQRk90DflaMBZfkQo5X5WkmLXDTGa0Ij3C
Mu+6IFMFtqThaIzjShEBK69ohzaNYklthUe7On7gF1KPxZb+j9c0dHZgRSm0t9qJ
GR3tfZvSqnKet/qhkPWRSck7bCasiIXh1IoOB0jHEvtqjnqpnG5TEdk7w9kT+Lbg
DG/p2vBaBJUbj3+gKYpdiSujEFpppG5fOW0+xwgSTlquqiZWiNopVuSA04z5IW1W
8gNpy+GfHc2bL8O0MoIiav+DShqdOd0OXBAFx6U9mvjLV3UbgAvMMOWVxoKozo6J
cBZqnBOL0ch+rKtHmBWL7WT9sq24fkikB2eVnZNsY4dgm6EjaSJbAzQX95ansgVp
aX7b1diTldU8bI1Jjhg+LWDmCtBhIi6IAB+pryLMXXGEsQ4F4oltOHjaedgXMv06
5jS1S72hr9F8INbjxxqAKXyELhVeeauroc5RFVJ7u5cUZYNlAlVKu7c7REy/dwSy
/uuB2uk4u2hEEFsSXbm8OBpBptElxAtSeASKfbqfIaqr6ywycgrFLdIcJhM4kLgj
psYcy4dEy8fpFKMuWuh6Yd0frxsDQwJ+5w5QG4TwQoCsCk3eJns6woAaatlYWb9G
ieuoEyeeDRpgucnqVL7HLzu0KA9KBXaMkO8JUQ4jw+oB9vzTOkqWOEnX99u7/D7E
5hdn2HmkG23mBG6bkHhBc3/MWpvvT72IgfSDcXargqFmdgWXlKkzzvvPbNy2lOh8
Q2DaxplkB640Da2KD7TP3jZKTmfoc1sUhmFrn9KoBwB+zdmVxdIH29Bdony8mh+4
ZOk4jVXkeP8SvVDtLKCaUPPBV9kIl1/JDIuAlYp/qnXdZaJlfCf+f7IBbUTazT8C
SI+Xez8MKPEyyCZY0W67kZjJAeAp7O1yBleiYg44zSa8Xn6c3sam3DoCMjOY5OBM
LG6hnu0LnBC+2abe4vp1h7B1lIKOWiCzmmiYkeQqVyFnsVjQVnHi2cBn6c4wJ0ag
M4YPQ/1PqLwMQDgdavSrVw2zACd4oRI/L+9J0X8ob5C6n1UXIjoQisGr6IyVmSO8
+byqVobCNBVH6QwJ2gkiiY7fEuHkXV9wBVzia4Nld6vCWVBXSUIxVSuq0W0D+LUE
9vPbjTV6ShnF4hqnjYtekfwQUWlJ+aoM3T6adRSQClv7LF4tP0GYE7azhtB5lNtN
r81I5uBb8+HDvxwxU4NixL00QuiLJb9cORD2g0lGYxIqRQaa/u/eb4LJq85XHU7v
W4VWjj28oRaXgeLrOjRHibnfcuNMVD32E7lXOBoyI4MoX1WxbkpVsYebQpTk44eM
nQH1ziHmeJOqfsTX283YgAoTBQATdu0//oYZEweKKt23PkXvbVs1VoZZZ9sAzvbJ
6v+Syvpl79JDqi98pzD0wHAKx218VQSAU4lDD3fCJPV5d/invSge6lPdbH5BPok4
RaxuseH/dPOl2cNMzZlOXqJMmzkHC64FPBe8n/kl3OraEZkaHB8WDGSeh8gcDMMw
w2kNKk7lpNJqghyd8CkPY3hmR0sHZEBd30lt66TT1O6v8+NIxsPt3lQKos49AXnd
wrHWgtRkdc/4eMmd3w2tmPE0DnWl4x3h++11nyx98YSeUT0/81vNuWPboZD/OSuC
pZU/2YBwqj/4rT3+VRfKq9ANCrYLyhJfpBtU6lwoty70h0U29VP75qG84hSfUfk5
GCcPA78kUKpnrtblvWHXvYR8edUtA0StAWHjICcAKIa/5eqllVRXmrimQ0hTxMnu
jIT22bfQZ4UueQVIdFAiiffHeLKnK1krZcv6mVZd+HY1sJd4glw3tsAbSYAmQLDM
ZHaw+0K+KQKVPktbrpbmYkAB/1prVkSlRpHDqBVdqx+U2ZBQJCG1A/OB01kcn43l
71z+XRZmuNpsabMChOI86B9yVGoE0SrxVSkSVUtEpz3YnmEA6uQBxXFImpWNRk3V
KgjCqXo9G8SFQgp35V9gQwFKU72yF4fMc/WxOx+Se0UhJwo3Dr78Kjtid5fKrKLd
2HnGfMNe9oo4OfaWP4c2w1y1naW90T1iYCEeqoGvDJqV/SXSrh6Gp2QlrlEwQ7uS
NFoQMZx7mU+rVfbY9H70fbnpxfl3QlC/0uP23qjvsSOLRpgyxPqWxa4jkUvk206H
xdrduxTiRCAkMB5vsroXGZroFSsHFwTAzoAvTUhuUceKeSFIKMrBk6lgg8hViWhr
eN6qvdfpWK6h88R/YIXkB8B9I59/h0du56KgtrtLJoswONao70hfxuBSK+I13J68
NkfEYOIQzSEZ1JBiarHgVJXpOXXIJZ2HplqW/8hzGtpPAjPuoxnEjPwpX2QtATOd
+cL+773nJbiXfw+/KDB0Px1Q0mUKYd2ZX0rdLnRQiY68BsQzONL/pR7hPkeGBDPv
n7prD1PZcq/nWkEgCMh0fp4UlpJnT9fpUSPSr9tYMznMR2tITtwH1W6/rqSkcRF4
AcRC8CJRKGzrMtRrLn4Ahx6I242p9rYZY/Xbc1CKLMkdfmz6qk6sjlyR/KkJYqLD
WZMGjN4cCudjcHAdF54WP2OSuMYoQ9LvF1G+wD3SmexzvIR3oIo59j3OcJg+wFrb
DPGn3uvxFnVVqNzkqjQ8fazptD6U3m7LCZ3EvRWwfeB8tRpAQLr6kVYe28iPMX4C
pgiglJzGnpbG5pRCAF/0BOPawx1WahMf9KnVsMhmO5K8iRNQ9nu8JdaMdUD+fBWr
El/ZEOQzw/8O3EzvXrLjQ7RihRVdr5UncZasQi+Dn/fR+1fUr3JWTkWuI9sYdjjj
MyXwjGCyx0g45+bPLDY8XX47Q9lUrJ28AAGdzGhXMYD35tjCv88dtdGuIxT8evc7
WCVcRl/ZSuDXDPm5N7iFVJLEAXTvgwdHHWX/BTVX1z5td1nZBOKfOrYYK0e5xlbv
kYVnmM5sLZFzsuGWQ5O1fSwsy7j+IfmZHLyRy95DgNM9lhM0fgTOD1OyUvwcNM6Y
XOSEGSaD4CWT4isAL9pNOi5Vog6A63RY0Qes2gv558v502JOhmNtZsKjZKSa3Twl
dxi2yEVLZcjWb2KiCTi5Rr3FNbO7wEwz4Cc4kMNKSJCxf5JsVJtLdvGBLvM2q1zX
cQ/kCg2sEZzVxg8EvrYYnf8qkE8FGuiA/2HjC7LbS0EunGqmI933hsfvvji/NyqH
D42FWw6liE/WoUz+QJ6YVUrOK5qvOV/9Q7p70oqRcCdEDLJNv/uai7RagAV2HMs/
JqzN/sNvq0cRFbfCztduPVTGoiC+/jX3WLqMLm3ArFLrbKMAc0VPBVAewldc/XfW
mxugI/rglHvTec1eRayjnnctx89qvjfoFYXfj9fWtPnbwRPgpsqPbP+4bu9bYI72
LkBta9CLK9eBLhSIWG1hAk+WKEvo5RwKomz391+dKm02jEY3dmkVbZQF780c8Z5H
5WBMiGURw/K3wE372etA8xpja4bsXxdocaPM4fBncjwIzTsyPH13QR9O1RxJTXu0
FPlbWVXDonRyKijhIykQCMSSkcgf51p2eHmym6gRVieru8Z4DOr0bUJVJULig6yS
w+3IuRfUj8/dEWWvNVJKq3jJCdjkVMJuQBowQqJHgEFcrkk7GjHQvVV5ZJsRwNML
3szVl/vomt1AUYyv/dn9DrudUsYlfYyR85IjTPbB9k/JtqbEpcN16izWusIo25lF
egbH0hQm5l4H064i4bmK4ZlDQTT8rTE3LZCoOhEeZmiGxh/68e8fm9sAkD7xNjX+
gVvF9ZUiWB5UQouQIo29gGPhh4HMLHX9ei3W0hUsmkfZT5N6Py9iwZDtnPsNxTgh
KeDxRk5uUeCRuPLGx1hJTyVGbNtK5kcR48l9VDFMWid7to+63c+X77bp/rgoPr5m
LYvQQPfvnJM2ghqmntxKfWLKXITW5nlSp5ilQJBv7qgX4qeiaA4cTj0TGkYIQZfc
6wz9Jkgm3pqazHCFMqzmhtr5zchUoIHtE/GxlRBrBoGxK/+YHz0vr2K41FeD64NO
pWlgMTbfhRP9HLcsR7zIAebatfGZKMWwG5JbwDnZ/9uyneP2ahcmPOLsY4Sfr4MR
c1+LL2j/N0dVyDX27GTZhydTmmsAbRomMRIX1R4joboEjd1fVgqby8KGZFZw4Qxi
m0iFQ4p4oxRIqdibtIG8iWLn6Jkjxfj2UGJP4mdZgQQ7K+8vepIPRWWUdSHDql+5
CTHeogyFdtjP0av1IrAd2l1dB26kcCvDI8+qxdeYQEZR5l8RKCiuWwdApWfYCCbE
s/HqYoLboPK3M5MRPkUulFCW85TOi8Jh1I3/GUrwWD2uoet15Ph1jacA9fE81poP
eQQvUbLxP/J64TsRNbuVhy3lS+kVdhjMXNUMEJS/WIkkQukObM++LCRKEnKCDuME
WvJxa4RMqiK1ZinEXKkkCGOBHK0cZYcsTqongy6R3MjjE6ZHkNL26pmXyUr0laPJ
PB+/D0BEAxw6jyOhhSKWb+3MgM4TUVl39h/2kGaNO26JLGOtvQm9Ri44MkvietLe
KW4HGqajJCQX7uZUZC12Dde3wnSgEwnxV3yekctXKj12RxCJXnUsM5oCLdXa4Sw/
/Xbpr93mZkhsgzWhDACqZFv6lvzFKTrBYeK92C9C+HL+8Bttngy/qtCYkmbyPElZ
m+V/ZwQBqp9h9D5DEofljU5hJfDk8qJFEqp4njcl5NoY36nDu22in/VDopRLBZ4j
8CMh4yIl5rtNGytZdI2XNaRsqfDOVa4/52KxLd0kj/KqGAI8DXQKTtBqMhr5ozU0
XrsJ0esptfor3VMfznQeo1hxYbRjT7D+cTpY5AXDzAavUoYF0K24DGWSt3oxAh4p
bL7Vzkqx2+aWPUR+zgmghMOzLUpw0BZPeTNmT2J9vAAkqnY4gtxmB9sTSOvj1AbL
ZzTJEn70GJe7uWug67pTqG0mZA4AMob7JDBV1JxHHE8G4IJXOcE98w/fqw1XI0uZ
tFZNA5gtoOfV9UAvPBZV9CfjPhQX1Y/OTm5An/E0LEZ2iq8UZ8B7XFw+HFlnr7Mt
reM13VUjr/pkzFLtcqjLHM2FfEwCNT5zIPgQVdOjFZYxy1Gxz09zBt64Hd6skoxd
aK52eK9MZrk5vaBFqiit2kzXc1utDsc78bcGQweaVGuO/gB+YabbmwXd8Srzw7w8
DReJ5qunhcK048pHROgw88/MgJPCu3Ukk+7ar2McScNZG0L9FzFF8CNWYjpN+iiH
pEFQY0vttD4gktG/eEzosngOcqd/Vuf40QjXdgILTJCzL6fnTuwNvETqbdbv9k8W
6keFODkOHxFs57v9upSnJ4FkJ7s5yoL/4znEidv8hlcLvdEnb2mHvQo2rX0Jw0gh
RboEGOwzGZyrzf3nOFfJMY79t7zg97zsOglnnBTQlc4O+kxbSIDRQ9L6ctP8MocA
rWfXqmqj/vxjneSQEeheSP2m/yZX1OSOfzeBFwXbbe9YgGORWzAeKTdqaYvXvWkR
WlGE8AUWcQLNqJHGfhXQL1VTRxf0TIlQOXgwy97pHskHOknwDqrZB+GMyuRHpkNG
VXnPpBAXhoqg+t1wHknKG3sTDKOgq5uI5k0GOo3x/6/FGPURhYpjuFrFbtxRp4cq
KpZ811FekbffZdZ/E38TjkkUcmBZmckBeA478ATUHFvmt6mwNXrDJteQ0h35XBzt
WnoBeR/WKU6mrbnj7P0V8JM5Z2ZvvtCU1n0VCrIaWhrlweTg0B6Vb6cmayID8Jag
03vuql3//yMSZkkBtTjgROmf+DqOpq5hWHm2qr7w2CRfBrQB0bRHgXUIBTTNR0yA
Tp8etbaRa4smuIbOIjxEshdk4+yFd0LUodAO7bVCX7zVNU7VQjtIGhGWNXT+ktlb
WnRtl737093YzckLKQIxnhIZ7X5HwTJuJswyTmmXSEH0u5pAIm4HJlVB9vrZy0YJ
IWnmYt2vPasunVZ6oFcopevAa9zgbDLB5hoeVhjds3Q4rvxSa2vVTLZU8QJm2i95
FW6er4wAMO/s296YddFArt52qiSk5mxx1x/lzbYZU4bvTYbCJdbfeHBUqI8U7FsX
qjTPZLiwX3H9u8o7M2d90j7GQH3Zw5thJbQGG9W8X4hR4I/ALfP1VWz8Nv5EdKtn
SEvRbx2Tw+XRobKinME1oZmTtba2py5FnW9bZ18iPlfZunMiG068XE/rkiUjWW+e
bBOE88Dg2se/1yCDUZeH4/J9hklqS2PvjTV0YA7vOBwGrDTf7dceP2JtFZes3FKp
R7BbvDmO6LQICVqhd723QvMUq3sP6suL/UBduqkVRUpHjAQ2F9GKDRCKe5Fi1Z+L
Ptp/mpEttWs164y4A6whGz9WFSOqadN2P6UfHJvHCRgLvGluDJ9D8ik+PdMeUkIZ
fBG2S18C68L0+mI1kkwfL1txf2IZhcgac2I8I/QZACl6qiQOQNwcAWV40Dn8WmgV
2PRppjZ/q/9EZA61XJY7+xkrL1+B1VR0vCdJU5ueT/B/wLzuFxKpQwsL7GWK3tyB
LS21VFDpCk6J8qGPXi0n6gptmAfHog5cNcObHIryGmjSvyHaUOfoq+7aJ0EvnTxx
xKpXB8s3uaX1sSi/8p16Jah+w8V5eLhVc+xA+wnKDo0J/y1Wnb5bcEliiNz85BDV
HORqMu25VqpRldVgSM/MWTibqwIVt+3Vt3I5p7HwphqUmGyTcJpcLT2ueu8fWaLh
DB1zLbWfajYHqJndQer8T1LjBgXbsc0nwwYugA1UcH2YwRe3Xgjn6EyduCGPEPlN
O8OwB3RxpMHENeGN5dbzmcLUTlnH7J7yVTapC244yBc4ShJHlWwwuyxOpy34TNVu
A5EVCSn5AAmQh03S6K/B6djwUlM8dtY2z7h5hRhShQ8I54kAnnM++qGlLNF0g3Zf
SVAzwOZjHgLUl/Uz37B6GD0dJEu8ysShCwDVjyD3D5mv9WmGKv1W34/1+8B6Ih+L
LyrMa1M8394k9mDPc7BGd/xxH2LwyiTV7L6sA4/gehYHAnP5HYvGQzVZPYodQwtk
4Mmf9y+kbzCDFJX6ZC0ny0oVzazWhxEmkuP/YiHdL/cgS4jBOFrI7gMGf7W2O/nN
VwtRB+0l241WbTNubDpxb6yJdVYq2uYYYssdY4AhO4PNtWkv8O20SxhCwUZUI8it
Ww1g/WpxJFzfCpiCV+yJdNUDG9iNG9TugQhR6xaNVLQgkKsW3hjK8EXtuZC85d74
brTNGnpX8+zykF7obbMUcd3l5q4UGyXsFNWhNs48TgMnBFAcGMLZRttJyMbL/gAt
88ZgMQcLwYREZMHuwiR/oRuoaBMtpoUhgBXLt596ueudvOv8aZa+fCABG56qgXxR
CGpoe3EMxv0jb1sEY5c7HkKR28G8cdlJwQcC4ovu/Xch6OMn1E7nQR2OmnqLERNP
/h7E3qYFFdnJfhvfzYhX5dMrIeAA6+fgxVEH4JmUUPJ4NDe71eg/gi5KU+rE62/L
YMQ+YBBevj62oQW0gLoZL1acYwqgUmUgg55JKSOpJV+TPXAaSFNn6071OrNi+0qU
GbOwRi9UnejDIXpDcF6R87mJD634dfWtmIey+/eBNu41v/UJK2eCKJDHmojvA+jM
Kk28OG5LiJphmDpYPXvca4wJwfEza0Q9TBQ+6ZdpfQEGdUj/EM/fa6zwOGT3RTYp
dpNdogJ+xgMkA4fUr7JZ0Q4k3v9I0aFMdMgi0eXGfHUozXsnk9EUVRyF/Z3kBKvn
ASWphs9drvD+3ch3GkUMAjx3rvvInk/61c3UmcGjXKJOdQLxxd5Sh0+zauv72xlh
gos3bZDvteD2z4oYgxJQe/B5AezDKVMXgN267coPGv3lYxMo/1Ay1R0FgBu/kwaI
oldGog38jguWPEfsCbuTkxmlzLCXzFYgmfzTBYb2fLSbs8xCnD2rDFuWo8UW1eV+
O0RlCGra4JoUh+HYPkzvKyqJN937SyszFUa9wpRzPpxZLE7he/YunAUrRDCfWZgD
eIU4HQeDtaUwJfoexs6bQzGJiW00Gj5Rj7lXk6yb3E0K2PxYy3uPhYtJ0C5fObsM
NHRYEkJ9vkcAYqaUgv/HgLUmv5k908/VO2oGhNN+d4bxGV4iN0YcUUE6XW9nWlXz
BamrkaMoPVW00+O1hoSLl3pBOOOYnFisGgWhpUz7bFnPuzMDiMSIOSbkbgCo8b33
II5EgTqxE2d6lRs62ic6JybTMuwlhFEhOm+w00L12GpKkkrLq9aRBLY1nZSWvwrh
hwAERREseCfBlQjSMQ8b7lYobHQXUs9xRl49bt7Co1dTNxWSzbLgJ7tofkbxcBFJ
+zX3Ws4hZTt+ngtZpMhcf6IRAN1VV/MDT9x9UIxiox3HXPi4y6May7AsOQSjbtJ4
7gPV2UIu64HRbMGe12cZSN0mmgVBYcexG6z8tdcrEs3XsxUBztoDUkoUw+WxwMc7
zKeP37jN95w16Rce2iaCm0g5dnp8JQvmh8E+so/ewqRX9R3x/PrGFlubfkwMgDQo
Yn15ukp13wgE+QdJx0IFybA+X1P7XfRLSiS/yqPtC+09clubdIBd5e2GNcVFxdOY
0q3ubJREkeDuWGC53rRl1T2jBlOiwp+mZMjCGOMvAoI7gJ+y+/RDqt9jusV937wJ
d3Of+imaD1BCVORnGtxt/iPpXtPxc/kZLn+gNRaSIi6NEg6NCodjYJh8frdo/SP+
gKMXS6KJKiNrZxlM5FSLhlIysK9jPCy1jwO8lHL3TkKUmpJGniKwnjY3yIWo6wV6
R8sDXAyx7I5TPDp7ZFAChZ9ZCxd8+SAl4yh7gwdH/Oq6VXUIwBcpmrjd5QASCiJb
1zW7sRJTcQAASqZHtmekBiZXhKg0yvW2BYhFVtfdfgihDz1Jmpbe6KHNmzbnAV9e
c2iMAmiLZw5x5de/MB0qZVRVNtyGLB6jUZitlz2JOsctkpN55h9fXNNJJQoG7X7H
oqxEwznn642WYpkN6YwtmQCTZTcv+VLH3qA5T4om6Z564KuK4QWRFm/sJNJbveIX
RTDklCFBJANfahmdXsNE8hp9Z/3ROaBWZ5GEBxmKy5OgJ/X8IDWKsbHTdT8qn33w
nPmS5E//AD0Xx9ZvXZkKnFDV66oqDvSDgylgFowo+uXNR2aPZhzBOroLibRlzIxC
z9Z2dzCcBB/J0Ch2yWM3gMk4awd7ZgdTTshwSJhppU2Xtr3JS/uRge3499GyXiRZ
mic1fjBptDCJcZ2jpe4j8fLgPDLABffyCX3yba99UWnvPXDk+n2aSH9ZM/B65J6Z
VRKekhs6pdeV19WzSSSOUSm0yIG618ZOtANs55LyNIfhhWbxDwTGaYL9u3jPvvh5
lXCdEMdoPYfVNYAQnJ5Na0skh8Z3nTtH29uZ0IyK/92qCFGEy59COu107LN7SS20
n5k+bXLoWfheZ1wJ3hiwk3wLdTDQeGUaZd1DcGOJlV+PA8u68mh8wvZRCS3bYcCU
DYdRW94JzV2eROMAzYHbUBBbQEORChx33M0XHrWQoDhhGJi3Y7Gal6iKjORdBRrk
Pk+Te/xhq87/XbyqKBqn+vMFX8mR0FzCrqJJjPuMznBt8Mq4nwfVVDhUhgdrmPMG
LhBI5EAjLSLp2puGjvaTE2UpaqWiKdz8f8d917nsLOYU3o2YhxTzhVDx/CKGaJsF
boVL0lqR/xTLOZcW0JMyrF8UWzhwR22QdCLMOT61SkaDnUBcNPiPta+fi1HGJ60W
ZCHlrFJhElcjsSgly98I/Od/ZpnOhj5S6p3ACzvaQHZxjmbEaMndV0uBPd2NjYDL
QcG0RPzjflbQ7OxB6Xz5pVxsmctqGncbG/2vNBVYSe3gZPCC5lHgqhanD8DINpse
k+PromFNy+2AJmIDNHNGUkxoSpSvDBQxzGG545sua6Ag1DHPvqLrRCeGNg+mBzKn
mrUha/TXXJMHthSZqeKjQ0Jz6Ykg5Ez/rP80c3skyl8bzRBwomvybMlt2i+q2qMJ
qwNSH0XQla043r0p5mO5iiGAQMzDHUd2n6SAwYVi6vAoQS1UshqimsiWc53W7Bqz
Qq7xeTmclEiaSSIhai1CWeaPAdhE4dbK4lueyOxWlHXsaqJpg0aniAZ9EUX6LaLu
frJbp8y0QBRZ22EkXmJtdp8Wd6S/kj7C7/fijy86NddApgc+/OOUM36rLwKPYRAP
IPNFfV96dE0egRQerXFSVjAyb+qlLL+66fQPXGHxL7FV8RIzlMnbq66W5kxiggMy
Zfly3tA6GFcMRDSDljOn2Gl7TZJbSWWJ6u3UXFmRcISo0OiiaojHkz4K7/q7+PLz
GgMQ364I2d6VWwh3veAkBYsViwejZ+u9OJAwvETq99RWvM3/KpusiL8x12SHuJZG
eylNRBc0pvza3quKS/qdzMBA7eOfOyMD63i+aEEhll+t+Ip3lTBxc+7pXQyZWTRW
F5T39MQZCfpuZWdJg2lAlEn6/qZ1xmRJTfxmwDiczzmDAvv3TWmcS+aB9U9cgbgh
qoiph96XPKLRXZVjcV8yKUifHzHAVk0sPg4v9LQxSIVFKNm2SxkW09jmxdmG6fyk
+Fasj3uAD6a3ni+ljBD4mb2fkrpXB1fB+9SP6EO0IbAu4tAnzv3i8mBRqBTXRNsn
vDFe+u8zFAyIFAAvKy9Ps/s1k5GLXvA8mPhm5xEIr+yOjsCATV4AtaLTukbwPtB/
NCIjeMwAErbrnV1mxXiqSn3OiUEk0Kv5rhF+SCTJWijqt9mQ3ysfUGFnFmmeov8Z
5SIW7jsWcyJijYJkfT3Srn7lZwC1S7r/BRoGytUR8HMR/RBWClvQpksNHrfQg6uY
+VMev9U19aBfOlgTSiBDXTBLnVp2GUtgvAeVJdwl0TKidxnEY9TKseUO9hYI1rUz
nYL6Fbd8MLvDYXm9/vyPmHXbqrv4/BRCaSuqFJ1uO3UM6S/VAeh2212gAj7CtkBU
Rr95nm9TtXbMSL7bR/im+VHgCMjjt1HWfp9cpJwTHCZeNZvWJYfbGTRJOofN7FaF
kItnJHfht0lGqtKvmWea5VHsK6J6VlldDNfOcWopbGbNp4J1GLnLBXnnlvyKp/HJ
+BRPHp9CLA8vwhTR/eoiQxv4/2qcPiUomXGjy+FDD+JmP5/WEw37xrlLvCGd+9+w
nL1+IxxQWXGkKuQ2qhnVAb6TYGk1tui4L3DhNGrhYeEs39jST+iR5hTfnZCagair
VEEwAnMfB483kyGteEFRdqstw6TPGG8nTXP+4LgXF+xNhKDEaosx2729PfVYTYbq
OVOJ87h0ILj1eE37k4iLDaKyCzr5YQNckCX6v/OfqOskYq6q7DuGYJxKsnWwLTCx
vLAD3cIcEbc0KX8aEjO51b4rMa/ltEIwTw8nKuSqL6KI+27DtzcAHoLAvKBWJ9QF
K96Nh20meQHH1HsIdHMoHqFE+7RF/pbdI8WsU15W77lo73A6oUDmMsAxjkQGBz+L
az0bq0snDkEAyskb42KI5/vo2xTYeGPtn+nR6hwV7FwPK3puOxtnipwSA13yo7Mz
mu/zV3cys2hCSkQ/n/MOWbTZUn2A1CD29/Zi+pkXII1cSpGueI/wvjbusb5dfTBC
5uI9gZlix+MwP21uBX1z1/MYwdziD0o/JHD8NRWjhwRhtmh6tEyrwCqUQHGAHrjB
YxLGGISyvtV65ZztVLVou3SOxCnVgGgxebp1Ytu0J5O/xbkC5eswnlrtLueN7wcR
1aBc0O2nCvDeisIJk/OKYri3VDqiOFJ12RP3qsH4ct/feAihqN4KNDRuh37cLuKL
z+9kfCBCwsTnl4rGjv16FynyU4QjIhzS0yFaQK/ptfM69o1faAly8GmHUDXOoBRn
aK6jZmLkwrp5sp5hwp0Amgw0JkLa6Q/zHjEVzMBffP5F6+qccm3Pu9PgKW65RDQj
3+ftNVLxbVeaajKbjW08FmEfGmT7q0FfttvcKDAqIwUwXltYuR1Jn7HcMUi6X9ZZ
jTUNLPkB90r9UvtPh5S/2tUvKxWuXBZrl/Sfsg+WxL6odo1BJ5GwoOQ/YudKkgNV
vfsS35HOWQBngLm1tzGj/1YjM15SXG1EK5NpG9pd2EYjtL0sJeyq8WwcuILswP93
pOcV28ZodfmdZim6yOSbUHFimuE1mEEUgkinG4OGsvcqPEByrONA6rz2lJq93I5G
ZikO/YvK81IUQSKM+NoLbyvG2eWbhVZX0OGgH0juYgivgIV9ILHo716yHiBvkJ1R
xBCY5R5juF5amlsc2idAGykfw1JomOi4ZzGG+uLyt2Ep6yDxkvSi7Dlnvu995qjI
7W0gPBgIyrwKqET0V7R3digcHYoop2EoSY6+ifpyOvYYLbpE/bCQlbjOXipvjw+w
q9seQ1fyo5Yg9a6Jx+enc/ZB57ufjkUbrN+9QshfjpDKxAqQfJlzsSpxOBHSN/S1
6JJ6seBVw9vcMYW/fe/i9vyiQ8ncsjGIljeYl70JB8zMTZsreqWnklYmiLPtbJZq
z8mEqAP1hKJm/x38F4Yee9PopaWV77spaKqqUpnCDh0U3nqTWfrJEpYszWe1YVyq
5AuRHiy+r03GxMtvjIZGdjFkLIhhjUdFE4kcdneNNhhZLcuaTAgT6mh2ZsF1Jh7M
Fd9VI0A16cpL7fgo9N95h3dp/gTg6MCveRJzUqSD6OwriCq6h7HF/QTlo1CXnC3y
L0YOPY4b57QgdFyPamQaO13pol9pwZCUrurPnm/aqtt1+OapMRciD2jtjjAPBX+p
c24oXdw/zKFSA3Vk85cHtFPfRMwGc5PIeeSsXNcDZWTPkRIZpqy1EM2lGj4sM+Ef
rHMVZED2YR3txe+yxddacejcP8nPqWly+MUPWL3RfoKbNrZsLIx9lSLICwIkaHnZ
n1RgL9QuvfysGLfT7b3A4hzgNSspWBxPqZ2wFX3yfp0X7qQlI4LpeYX66tF2kh9H
gu7FltQq99czHvEamlxWLNFFtm9PtuC/sz7FxYZ1sSDnHzH19YxPZEMJvT57Dqr/
AuNxP1lR7qeDTjxJ3fNRf7OSDex3/awOtgO/Cm/XsJbOeRQwK1AYVK9dG+r4XqFm
jJfTmD5hw4Nw7aSGXEC0xHmBn30wBW+XPGrCC271iXT2DF/DCqco08fZDh5olxf4
quyrnnQp8V+A6xDwlNU0ELvbb9n+b5dNzvZ98dS0fAPmbtLIVr0lv14CIwWQjn3g
nYPVxu2zyrjISah0TWSfyMR4tiuzLPhyrvVWWW16seiG9HX6Rr2/JWfrqjJqFXl9
akC6W02ssjizOap/ugqWXCM1HNaDAhqxVu4gaCS5rSH72LoTxd8gVKyU/1UHr7fo
wTZkDVeo57UEz4l7BnAQs+YfuM3k+mjVKQd5Yn9ZRMjAMHwfEmAGzsX7TVLkFmQR
fbdG80soMveOpoaO3JzpWBYoygFH2v0zh3cIjAYpz4R3/DSk77uCwPIYMRFJYKh6
QNMdk73zqNUKwTYPNr3gbyhxue6jBo5N/wpQoJkP5bPa2a/ZhN008mcboPMTSW5B
jKIENYB9jCKuYnmPOH1+E565qQwL0Ux3VxIxP1oW7wKxyJApze/W+MSDocw5mwVH
iPvuXFw+yCg+bhsqbcud6O2QRTFYPeMmf3TlHQEu+QuIpexgHcLGsHwO7+ip5tGd
aN3MAL9LEj37YbWlEJHgeAC2O8EOlsvDFWZI6i2gZCmYRmMVhUNNu9nea7mtut3I
B+rvBYbGDpCxZI9EdTLs8k5o6b8dqDlhUGl5TvnReoozN/IwQPvxl456gKstHPWD
TLGQHyQSzAr9dOlyek11V0FXOKlFxMlb+5d3XQejidN2TJsfNGIZ5c9P+pRQwiCR
vca6mU3q5MfKwfKW7YPEg5i5ZTMJGW+e9MxuRzjGpWHRbr2r+IetfcV8xfY8K9Zl
Y2EcpXza6VP/r41+Z6+rPQrX3nocxQRezr28ftqxNC08QBH9GhSSgg/8n5vd1C2Y
95w0xBnhz8V+6nGF+Nxjd9vrrzxZ5qrIyZqKv1iSsQTVDACE0pobfxbiRf6ewRp/
ILFN89SMKdVapsbmb6U6tSlowDz+qysdTlYAouR0TS4YyFnMeP3uoM08tXXOvbo/
TAg2oXTiJ9LiZLnZ3c0SQtKtiPjvY5KC1mR+Gda5AOHaWHlwZuyXk3EeV6CNZEXQ
UPpYMSHAA9HGeqWzffo+4qPZoWmXT2LlcK/uxUwxydwr5aV7whrT7gNB5sRZDkWp
s7JaVsO2kzfnD7EWL3wifK2oYedigXgxKSoarR9Z9RLBiZNi0Ha3ZOo7Q8ccGY3u
SZJXoTEquMLdeJNzoX+fG40V0foqpDdl3/aVbuXfDqdjlvDIseG72j1vqwiKL/F2
N286GQIeM8EG4UpfICWOaT1t/qLrl/Zgl2ME+ZYqe/EnAuxrBK+ufifiN7DFfg8w
txzRREuNMKhLt201yjVb9cQQetjqHXJreZncmUUzbxDItkTvLBND9XSckVxi3sCE
eWJBzQ/mVNO3Ev8cLGopsm5RZMX/sfHS7pWa89xk+DTNJ9xFIETorAevqQsbNNAm
9tAyt6/cebiSb5tIFyRXsiwpB3L3v3LGPkAY5KGe3aSxIG1EehSQ5DQquZ7gTr2o
TqtZ+K3XU0T95rVDoLcaGby+ClSR7L5q7A1L589+IuVhmgBBHThmaKFLKQkwAp3u
7AV3t0za3pivYQXGTQhKheZvkmncbGarPcAWBY5pQVsusIctM6bokOPJj/HYRlJv
Alw9bAyLva6vIpYWP4EM/ipCJWvYwCVJ2csk3zekdOArRfDynO/zGu6CPmbWAqPa
KnCJr6lo1LHbX4dUKkdFlLPjiVWj1ffM/RmJ9DNCTTRMcg/o+A79P7vLrzqKeRit
DwIxgQHKzPwK2da3lzZwMDWXW/bqm6NSsSkUY75NSucJC65FysuqTJHwPsUcLiRr
H6xIpFWKg7HNyigyvf2mfXXXG9whsvkf7CFr2yp/BKFU4rCUKvbjEmSo/KmaUFXk
F91yEKaysvXA0CMWcapsIcdHEUUlkdvvrmSwNTlaBzktCxj43HQyD7Ps2+U4pqJ5
q94OjYQVf7rhrFBfivS3dhPbCeEzotSHPD+Hfg4LA8Zx7UoskearloWQM85SpwXp
9kgkYGNX46QtnH2ADcZyWUSGc1f3xPubDtKcIY2i2in7V9EiMq0kxvc8bfaZKWD6
RW318VUaUj/ZXHEJ4rwF+Dz2WgAdkr75LN/kmLVSIftct7OakKJ1DMzUcBw6Nv7S
S6Zp1lo/TgIrrWalAJpEAbgWTWeDjGOOYBPTgt8wqYLBSafX0sQvVHZoesScjENu
Fh0J906nDPYj4XSVIF5+IauNrepnS7T2CX2o3y43KkU0eT0Kpr90YwpydrHJ5AZ7
fFwCJjC8TduzJJhDpIhewyjeOvxvkeEngqjEP0mo9232CUENvxyCrAJGSQKvH1MN
VMPOFH7a+O4IpMF2wVqYZ/9q8TU5rKM9HFL+luc5FVb/ALSmAr1kIHqcJilvGs06
Cb1S4Nslro+fbaOtekGBvJm7L+928U0BxSggS9yaLKV6FsvS2ZKKKXTZD8ByzoLi
aCXdQ5sDDKRcapEPWMy7xK2pb6E+DbfuQIIaHDIIAXkBt1qp3I51iUY2HXnWnR32
qsKqWIPknT7bGOqUx/2senSKPr1gXwAq7zXxW8FP8vjTlp44Z3ueBW7SjnyxAi3W
+Lx3tivtnK6YqPwODjoFLM6RUrQhzHjKj60GrKqOlqr4xCZOo5JuZMuMtwq5fE99
ZyMBiEyyrvn5rf47xoDBlGPEDE9FPMns1shHSuvSFXiI2BpeM1EpBBD6NOZrtuG0
6BQisGFvX6gu39o27lvy9LgRaKiLZSuJV4GWPju6jaokc/rDFFvWrm085VdSk800
h+G7n4KbscErXTxEavQkYS8KfuKDZap97ylJXiopbYPHBShP6TkGGOV9VRViMhkd
PYvTETCAmx9ZdAS+4JunmjwOq96Rjj7YKRtoi2Lw+4Nh4ySyWvyFL+J2LTBOOVKT
vo7pDsZhMIaghdBmvpJ1gLvYOqlHlzgsbDlHy8kCOn6VdW7TZKvdpq19g1+eZ1ZJ
XlucBxT7bPkGacVu73omuKWS/i4W3SxcxZZJr5As59jEke28un0i4lg/zxZGSUl1
9tutHKeY/m8zmNzRgEqdH55Uc+VJ05XmMPuB5LxjoB2XMEIOlUkoG4NAul00U0SP
5nkpaZ+n3wYtGDS9FxUUc8//yo0LcuW1FK7fjTE5Fqh3Qn8scZpQcgdxx7FMmgBS
3/mlq3uNNUudouY5QNvTZYJ5ZHhyVnu+UcJQOWtU+fNphW5G2JoqEQj3Q9c4MiWr
E12aVSxKxQIq9pTtKLZ5UCH4azrR5NS/lo18gkxT02rEBQ+FeutVd9e9iNNAHnWA
L4QKL9Or/ja0elu6E0Sc4hxl0qVGxa943JcLpyW05JVwx/EVmmk9AMD8P0TXQ7KY
uozR/LG0GaY5WQlNex5F9Kj7buCBObmE9Rx8zx9BtMYrW45c7zKCXaGdOr1Mw0TQ
m8l3+M7NAiUzui9tj4p5+n1U/r8fgxeM/XkTFnf3Icmvxw2W9YiHkCogBduoOMHM
9nQyFRoCD8U9gNO65MnZqLrZMeQWaC+m2gLyh/MxW/nYmLGS+yHiB75DKE0yHp6C
MGsOrijeDfEZeDUFtyOfvcT5NnWg7gfS/URq/VR9Wi0udZr7LZgGypsgKaLcetaf
h1a4ofDVzu/+f3z50Txa7i2N9+iNVt41yclB6L3KuGboBXDvYlryFH1/U3JPTz2q
yNFrhEOVcQOt7X8R6ECT+zMl+5dAb+C/aoSTS5U1TNLxdfDJv2S2+2VIn+Y1STfZ
dDMPO37iuwRQiDcvGbn9VIWdBQNi3AXsr7iQMDFrtBmo0Jh2UzeqCVrMO1tjkQpE
gT0FHwnzWB9PFrybj9CANGwTb4yBzB8G+YmsFSkhdE2/ca6a7hnHn7yvti+bk8EU
udXF9fRGzKE055RAr+noSWCyu99QmTrXC/OLrgac54+xfrteCr6rwlfpGh9f+9AD
3gANWWQpXju81lyIHhwzbzZKKWdV9RIgQRhbr/8tHTQvm8MwrSspf190XUVbM51w
s5ZGhsDv9lSUR+D2dPI+ZYra/SeXvagIRY6exr7XChGap9N2Eg0lCUBSmBkY8CPP
ZLiDZFUZeSg6eLjgToUigOBlwvHuwTyGrldNu4fFnKRdrOKj8FyGC4HKGxoCBoXo
5uvO5/A0XDFd1XYgWRfiNeT6qVc42cz6/GL9BOSTA2x8OM/YSQ5WNUrx8e5BAWB0
HlQ2o6R0YGTzSTwfxp+3waUOHf7mVMpJ0vjQeFWOthINWwugK+Menb0bG3EZYD9f
sBsTPkOiLYCCNcFf0zS6DnwAWGGrOTXwODCelErLjsKV4g5nwzKHZ6MNNGUhq+Z0
cJddWNa5gDvyoFy+ych8xVjm764uSWU5qCqxGYXMg254wsqTpQ/Ck9acKRje19c2
V6S4qqX13Sb9tdLlGY042qrn+kMdNirOQhbgksMDlgS4EKSHIdmQ6XrLeV6H292Q
HKOYQmJ6guoriOcyH17koxEVAO/qpBkMTeTTHpwFs3WkS1pW5UmxAxIPxIk4m+/l
YeMJX77Bao6G79nHP4g/bBWBp0k8Ub1QDULYgnnS7iow+v07IP0ZDsYLrTERKnBF
hAX40Y0k75f1Zjl9Gwc1AhOG1tLMNWQmu8AaFwFzGMxUFAez7BMpY/93H4hD+i8T
Z5B1pH3nYfhKsf2HN8h74z1duaQ3279b9swgidzPMgkEue2Q3e3+qrDhf0juNft1
aIvy1if3qXK9DIwZB6Rtfi4egZEgiPRXUK8u51DZjktLJZn+bzeug/oPhP9Kmntv
sEWS8RMc56x6yc+JQW9lg8TGN7FiYjqGM0p/hQ7cRFRUkHnrwLW/Udkn3kjpxDGu
ReL/W/o8/a/UnCOxbOGI39RN08wc+PqeA6i5uCflppc0BPsmkAZuB8g32XIY4yca
zjVoug65iMHZWGVHRnlkdvtnR+sTVvY+TcpXdlYRAU+FaOMNjFGfjJg0JALQDvdc
1hiSrVYZXn0iCV8XoMbHajNEfTf+ZxmTlMXwM2PCznmQu82x17Trmm2AQtjA8ita
haYIqyJ3qyUfiRFg1peQrfSEz/iXbcg6tDm6gM0TKQIPNZF/DHPFavKpEyrI488E
iWmsNL65vXOsIuzwQrSsE06c/jamgnYsME9kPyegICao0htXxSu1B3WJ35bSJsm1
YiWuTxbHEtP64p47l7wJ3TaiuUz7KMbCj+xSkRpuBnDOuRvnc2w/tOE6OcibxFMD
0cirPQ4YZt4LYmVPcTKDKr9TdMtxv8QVoMb7ThPp/gdFcQNoWBJBuD24sw+Ku6hq
JWCcTeXTNW6FFGSSDBpgRFNvGamBMmMK0EPFOsyzvs3IWHNYLjJMOYuxL/+tgbdf
CCRC2n8RJOGJhgTt28NgrSdoj4NzP8J6a6z2KZoiCySZBlJkSaNyr5GxjzvjjPQ3
KVg5QFtJiC9ukzv/8SI3ukQOW3TuU6IQ7DcL15BXQvmYKMCz6opanjBUOs+GkP6x
4/+bfuWwFfEN4O2zyOmnHJS7YAKC+XLZyeaxcAgMAYUruDiLw7zBVJADCll3LJ6z
yJT1Q9R78c9xT3raIed5n9vtEMF7aRNevCXw78wV8ahi8Uf1CW8Adi+tQYpkzP3G
y/ee50MAiPPoAtHkb3LwRYGxMgtPKln6GtokRfcu6/1EWd6Ex+EThxvl1EtbODJD
7O2TQCNIqitppm9xvtkipwOTLMezr8FFsaCH9xwpYB54pgkvQGWrQB/TvXE7ndQh
S9YoE0gDWmh8tO0NSL5gqBeY2QKcjvEd+cyX000CuT3FO5q3YxI2RPqAj9VZjA3+
YagYXCdWzvYZn9ibXolmbCwMDAUOJK6DB3zwX2u211xyUa2L3mLAksBvPhY3IOAP
RPWyUFxthqKkPpHc+4Hw0LG79WYqNV/D5arJp6TIoRScYFyGX0zoFVkhJwadKtse
EbSdvQBtr69O6Qaq1cB73lsEQ5ZJGqub1iAg1O/y8jdN7X7W120sz9ad3MfPFOjv
13wh6jhBVliIIwiPdjgGXXvWM9T9x6OpjXSqkevMvDcpSJ8BnHv9b8/8c5CldEpo
Pw32vJeBXrjBTupi5m8RLVFDyrTdy2Yq37rMgjcofUYmOy2rY/QElYZFci5mpzoG
mWzcNWWbTqD6w9kXwlbCEL/J/+o5gox5/ZeGWzXJa7F4O/sXcCviOX+s8uEPKlry
x5lk8KgESYuiaVDNFr6Ob+HtCVCVneX1gTeQ5dLT9kjCmYnitzrQ1WGt7mPAgZD0
0SxyAwT8C23qtSnAc3KDM/EBIsH9711vpxgwiRNlq9HO79K/7aExfq2sxke/fWAH
oVgTn8WQ2YBxzaJXU9pyXkwvGdLKamvh38hRGGWlP6/XrrIv1UaYZjyeck/xpgsG
boW+b6uvmd9LiLb7Cr0bKdIJhndsXM7vTZzVk8Kh1UX7VTQKdzztDxiwGSN2L3Gs
61KOIR2e2cj8/y3u2y5cvcBxyn1NwYummt1Pl4nvmJ5RvSplmZ9CA2/tT2Dy4r4m
+eMmizpcW8TlSWHAItTWVFM30RULwdGpZcYECSt0z8FUjd5r9DImOda3Ll6H4R7m
FShq7TdQdDSDz5snIVrXCdubdNeQ9SL4EJ02sQ2kSTroCn2dMZFruxKu1df5fQOh
nTof/yaSHfrYflWNSwh7nPlQbNJ3q/ecqZpV/tcVpUOzFoFCxaOqc4ys084NyaMK
8KPuFRPMkIjvTNlEeaUtTTr8iVHpcnnivdTm4eLzyDJG1MXjt4AfgWRb90nShYCo
A+SJxshKyJDH1UG7uQUnC88fjFpkzXSsC0bquVjt+pBv8juEbl+4AJWa0tYFXZLQ
vQu7XFBvrG7VUtdAjJ15x9M2H9+szI9pCrUhj37XENKml34h1jPxMaf6qsy+/iG3
JxGrTKRIOK64J+tx+JGLVXPMkDt7IMRJyD/4GT7zPTNMWhmykQA49868NR6mhWQb
EYn12CUcGUkgbhcdq3MduW1RgnWfzxMPW3H4H9l7pfElOIAr8BkJqXezd2zds+pd
COyaP2AvQhFGg0a29FW4sE4wkz65btELhCY3zlTQJVEmYBE7HaNu1vPUe4aI7iJg
bs+xje3KSLEkUj8M99DQVOyhv0o4RX2pJkmI2dqX9UUQYOoUvD/wu3WTqFh7mt3A
BO+IfL4i663u6js/tOUZ8ltwHGxkE4TNybeqFEY3eh8U5KJHkhZjW9ZOYQYX/uzM
/xuHnrV8Z1wse9riuICTgQ/WRaT3KMYAfRIq4/BLu3q5pp54iTzSij/ILUv4+3Ah
a0EJBd0a5FtqOIV8IhJCX0SHY7SghKO6B7HkEox+Fat4cv4HOFTJRa07KTG2lNre
od0Sal5q6+h7sC8y6LQHtXCDZ1mFBVcXQt6bDVw3BVc4Eyd0Ia26Yh04nahZUiPI
+umcMtZjOgzVktXvrgimhK5itC6NKfbrVsgn3T4/vY64VMldIeb3mjfSzXCafuak
/D6rPIx1d6reKVGkiP6j0XMR2CXB+5nh4tdUXM54d/ZaqSZzOicLOl4zvHO92T+H
nmImtFS8JgAyTQ2JYVWJLw1Yqz9j0ONq1C/cty/FsN8jddb7EHVjqC6STqCWt5Ge
hh1Q4rCC6o7ASFbb67bFt1EkdNBGQJSxJK9UUtJOo9bYsxN29HOuRACNqe6cNxra
TH1wTyNxNJkWQ3YGOo81AcBjNAuNx7aR+dMf2SCZ++faYon0zJh6WU/WsqB5Ceya
GsIEyf0535a3jQOm3z2Y5IxOZpj5+ba/v6Kl4yClbiPyW/jVC1jmcgKGZGXgEQXG
haKulT440UtVidHp8XwH5KLssD/iuL0KM2adpy4LhzP+GCmWiZFr6bCYQfR7dP9e
5zS+fXxtjtZ2S9Ym0qzOkrb3S0yEBn5uaKY9odG5sybjjS0bIE2b3jB9Ew2GOTT/
mEgfjrQFKF6vVIWZSrfywR1UP6Sz8F/uNhp76k1iS7f/6y4fY4M/Qi/RxuiKQIop
9ffYPk4Rd0pu/wx+JJVrH6XyD7t3zxYklI3J4YZ6To2WUkmJ2YcvVQMns/tS3Yq5
x+NiuS9tnn+wYDUXBqMCBoNl7glb4RIcR1fjdgEEPg30SQGi8/1ApYGglgCu4c2r
6jA1mLFcKsIsI2fJWQZF0qEgTd1RQPqK76HuLjsSLz/uozt6mre37RaZQ2v5OFPB
GOBvtF08/+w8VXsKBtYn68Mc/cJS1wKIkOhIIaz4mD2q6MGk5d6SBc/CcchUys7q
xHBRJPtdtyR8Bh+ckm/Cc4gEU7rUd0d92P9dXOzd0/T+F80OV+8BHHP3y18QEE2t
UgBkI/u+2T4JTvTEWFL24MafnnZg8q3Avr2OqNYn43U059jyeYitYJ2J3mxGBy3C
HtnB0xxEVag6xnHzi9g4xQIoSyHFT/UjVifRoTpqlP0a2RZOyJ/ExQwBEdbQuY7s
KfL7OGbOsILJ3AIb2sKGc+aRQHTMul2d2pOg+cl/y8/dIe1Nj9m7AqtUgqy4ltot
VjqAAEQmG7quzT6EcWco+mi0IhF8nwCldryL7UxTp5ihE/V3Rr9aU3GT7Zz28fC1
Z5DXHqinq1fDD3zSbz3dCLt+PCVk++RTGJVPThPd63EqymXLPJgY8PnkX9t3sP/d
MuX3kY7ij5MJCzaWpXgPM/dOD+pN2uUIIg+G4b+w9Nv7ifLzlbPJEevYHPxpCuI1
JjJIqkJyjkFFSOgVW2T1hkX6JioboqIKfNXla788fUVF3y2hZo4d6X9reg6AzOiP
MOhYDj25PnfmWRTYChe7n5bGX6aedBKz2dADzfGC0kU2qnpv+mvgxxq+t9ZuHv3a
y1p6/ERuQwWlEaZTgdsbuzeEVyP2okzgqY4FlG/U0scx8Eg1E0YJwfqLLFr7lMcu
yXww7aFzboWs0lJA4k18v1OjVK9ndSC8KaiyPoqzBHPteFRoysLATvOpl6cRCnT7
uXUjLSmvkxrMAoQ0yq1m12fK2rDblUWH8KNBjBThLgILHyxSwz/CgdoKHSskTLG8
I1WgedPW1PDtlZ+BR4Wy4GwJp6Lck3BJ7PTDxSr6fVuL58fWqI6QrBmkWrWrP/NE
JSd/aEIuSg7cU/qbwghgLHFePS6EaLZjC3CelFNSe+4utE6Tr6fagGKccElKm5Zv
ASJXN2zpMkJED+4BCK6JQLFedRno+k4qmJyFTma0jE4q51FSdI60ciyUuBUnVeQ0
wsjtddMEv8ZPp/iaXTUxnXsHvWoalGrSKJs47MKO4EQxL8MNPpWNMzx4VJflIJbi
rcedwmaqLvWgz5Op+Eva2BR5WoIvpKiAU9IYkRvMGND/w8srSpsY5D4AWFULexG4
fbq3ks34WVD75eT62+aOZtwAcj7FD7Wo0SO/MHQsIgGXzoBgA0F9VtB5PYWuusR0
Dx5sPGqEZzxRPuOrQ5pKkhK9CJxkUOEFt9atTGdtU+0wmzr3ijcEzBNjYxY+aiVj
pohYq0wR6hJUI1urV46DYL++i3TZBEJx9gHIQwGiGDsNCuEbVnjSjJfYfQETXy9l
0YkZ18GD+y8cklAkRpfvyVeWnZpqvKNM8eKgPW0vl6BE81gg5/MrSGdY8/p5TyuZ
G2j48IZrgEka00KzyHO8gMXE4EJNhJCureuJ9RU2gPwVQTw/x/MYQrXAlUY0eYyJ
OuILF1UIhgk+BvwWxgA5MJnaFhiunX/S5W4V8UJdeORh5cb65MKpNjXySnI8ctiX
ee8nfost1cCyC3Zx24B7Dc7imN8C3AKPEKVVCkrbcb9EtqXXkZA6BeWk+4KTJfEK
0+wd/W1ftmxGqf22GJZNci4VB51hl8tsf4y/pY/TSgdCme1qafArekGtCkJdTa73
+/8L+p0Cdujdseb2++ov6npopH9U1OTbBc1mGrssW9H8shgovrr7EN0jvKNfndiK
vjB23K+e2GFLwYDEyRACu+3LU0XrMwp2FEZwmJkWmPdtTBWgN1uE8k0iOuY7An7f
hMkL3oq+hspIpWxJHjOrvaVAAbyGCOVdfDfhI87L1M6CCCRfnIE2t8s3Z52c8TVZ
r6h1Rmt6xFyWkv+sKMUb6D7WlnE/fpLDZqm8LYGDq4boqF+nUjUob28VdQmTJBrd
ytcS1MNFF3Tt/+jTgB19XE3VfTi4Ep/1OZjgitK4tfFu5FEP+jDwian4AfUyG6dm
h+IxsuVMW0VIP6nICR0TZPJpodzU6hQzLnHf+xTpZ8reM9rsmS5/+p9ihUx4Nnzq
ztrGm2jqPdohlGa/BuguiHNE14dp5ZdolvQMzrsUWbkUVdR5fCm2HLq0CJKAT2Sq
Z/wmrxzQZCJP4m5amVcXvQW7GdLRr/kocPxFbBOKU9ggkQzwds/UEZcyYusNMXKJ
RfJXrXI7CDuXpcj3USfgoKoxsrBTZbii2bPzCvsO0Z4ywDkvae+RatUNOU4JHo7a
JXnE2tclTkolu4EadlD3C4E6s8ioyz9iwI8BGTfNvuomCemif2i9dAXw2IurcxOw
TRSwIc6UvvwJCpUX7wf58+mt6zJ/pF/X5vtBRMtjiF7PAfafzE8TNhcM/7xawGG+
tcqC8LXXuxJNrHOLpicXyp3cDBP1pV/c6E78w1wqsY0c0qaWUfOZrxLS9BjwN7U4
kT34922gvGFdeRUC/4DfR+DTVnZNltOycrY9uYWwA6ni+OMUYL5rC7koevTg7uFE
YhSQVsCioOypAP7iV8k9adHkgii5JZh947zM9ik9X0yrXCyFY5NIeVWkE5gHdszC
Zfrzj+rZfWzf1OTFie1EROxDOAQIJrJpPnxY8WjVX6J2IXfrzx8w5i5ML5nn3o/L
dWLFQY51+x5Y1UtcDJT5aFt2XLvVqxysb/Tv2/nReKlk+gs4WkejPg0e58Ssg51p
trj00MJnborKgH7dJjm6XAKspjk6sZ/53FCPwxSipeepOE32B7CnkMxQf8EzaJlC
nIIlKzUn3S44X8b00eOoEd0S7/2ElC6DX7OqTVsiGH2UdCwQa4XDzm0lO0nkVbcO
Lf1K+rkrwdSOvVrHF9/n/OnQRak0KHVJS3HyLd3zR1fWNeCrzdk6MGy6dyMDrpvm
g6zU2l4VsYBproq5E8HitUBS8En+OO28nKHM+D8dHAokl3gRTI+vpDk+O0DpdqyB
VINWfHtWqRfZnLMOigHuP4QOOildXb0yaJFNPCDSedt1lF1NpGoXRtCA6jPXgPHr
NMiAUHnnYZeyhVNQ8IqaT7hFhuY6evmkMZ7UmkeNe4s81CjlRiXHBM/weX2AQ4NO
jOJJUUQLVhd5VNc3xKzUHNcXmkJbwWUWTKOP9zi26gRqPz/wtmZbildHLndfR3jU
3HKn/eX4kJW0/uS+ihifzd4UDjVw0X97JUUITfXaaSwd+/+YjoTheH4JvDHYfd0O
xuaL46TBuv/NId6JcJlICtnzjZOwee3pRsDP4XFvi8YM/5yQ7J3hEF70T8LgPhqf
QcdzIZ9/L0LKZ9XAsinYtUB3HlnMI4vsrqAoQb2NGHDDiKXs4t7NPe8kEkVv1DKp
vryOZMiF8gWhnKoppeNEXQiOqKivDWRc+pAsZSJp49uVOxzuJbVdJScppkDTNm64
1zFXGSGwGY6Jy7x2OLGxT0r1TEo/M+r+5HxfLnjjh+r0xBKvq0VXuKEQOYraltUi
TdYCGjypLUqAy/fbGKFiwnpMfJLT0ZRJQ6VNFho6G2luCWBQiz/jj/aLwY+j5K94
2QCgMSmFAK5ZAJh2AZu1RJ6xgoWIR0sduy7CGu025wetjkLobmONw9H0agCTFcTT
YPSlNAAQ78SRg7YfJKhFHtL5O9whTSLRKo9IaCfowtlXu+8rPXK5CiU6OxiMu0b+
S8oPsJK7wzELvdY+mvBC3GyMT2MhT2IPphRM72+ZOqo1hKYSq0GGFAAukt9EwAPz
Iyqo9owKB/c+ESccXTTnqakSLFJV5NcNBuipTE52XeTLOAgTARpzjtOquhMIz4xM
m+qlogJqxJzicjUhczODl0EncwVqDSOnZpRZLZfcSnpZwXplzbkiTKYfnBbFp4S+
0gIBJ+4+9yRFpirSXTnD5TwrpvyU9UoHFKQgN+2KxvMBs0VGFdwZ9bG+y4jaJVgH
PSrtOgAFtubd60IR8H0M+QkfkwirV5dbttlGF7QO7t/jTAXhXiBZOtmjw/txGU6g
t+t28Ihnisp34LucQYM7RrKPeyTKF9cN2tB2DEPWet6BECLmISQVkxFQ/yJueKvs
QB8Moq5YuHB8ZijSjZjJEluPANHHoqQf7es44o6YW5IEzCu1VXNdCmwlT+OAHZKa
YnsCX9Gpw/C/3FYOAaRU4ccqfi+dNyUJqPrU3umvWJv0/bnCF/7srgHkRCroscjJ
bKaGZASu63jYCvuuiLSp+HHI1rbn9C8xcRTMlIK+lh2umBH0yHxpZGrRti7b8vri
m4NcLRyNWmh3OXqCchkunhkvGl5fKej5weT0s+B+dfTkV9+JzwFjTvgqsS0fNKFk
rEDTT/06BlZByYT4IUXTuUWbevV1sQFnFTGhIXaUz4j18oWRrghvJMFx7nHT09Sz
KAkVa4bUwitQPPfZF/upqD6jRDOCXb8lYmNqcq8CwemXt+ncW/Xq0/scSTNaysAU
oev2YCdq/jwUAGIzH7WzcBrHAHpz/nLSFP2vDfuaA3wv8bGupEXLLdd2Scn3gSnu
Gkx4vsL0XxX2LSbmV2/bS3yfip+IX2e0u4FXiNDKC2aAsDIcqVS5jerK2+vXb0Vk
xUjErKzx0rTljgLcbicfFyn7EP96k65ee2IMCC5Aqq/vZUcLusH16ZkJ9aVuaNW6
iZCG4hIYrU5oMnu+zP7AxauFH+zUBeK93OuOWP5IvBi4tDjxGrzYdm5il5nQ64Sm
BcxT38M4xvzQh/eA6C5sXYLS4hkKZPy/gXDU43VMiRUIA0cwsuSeZfbunWBlUDj0
Q80w/VezffjPskts04ovKelUi+i+fM+dFff3iiPTirAc0mF9UhFfi/l2EW6Arr1j
8ExIPRr5NjNJnnHGajklt+fwD6GEtsi30NeLZJ9D8tdWTcUIyXPFy/Ro8hjeJ8KK
ZmcV2NAp8j0mDd7Y8+ieX90OSHtscHBP0dZ1uEBPIXzem4okBBe2msSJDtqXWBXF
eRQ+2ZLH22rPN0tT17wrbdwLbK/Kqn1YKL4ibh9INAAZM2eju7rYeX82l730wIwv
R4GTEX5sDtZUc+Mip3CobJqjjcqU1Kewgnm8jTCq/Iskmq8JzGkRVMf5ugqOD5W8
CBA/xFNK+mghzKskSKJilhFJ9WxEVvBGkusXjLryOyf6rdhr8oRzOSGeX1kuC3uv
qElUdhg93f7hWuNES7G4aSK4MjQ1NlGs+wSRiFiD/xVCxI1pKh6QzfWudzgX8s+X
RQoFjAJG05A5VXHOWmtFEYm65jdtpOaA4yDze6hdo+4gQqaSFBthwTtC+b23eF/w
vG63z+V1XYujhJwVci2JLGdrsXVnnKHxgTqdbJJBWzk5qfugcFNcGly+SLyEKNtk
OKfYaUpk+Afys6Mm0FHJOraAOPznkhvCzTsEIi3zF8Fn1KK4mb0jh16ifL29Pmz8
dXQRGYeqowWmXwpmtrKYKNe39Vlnyl5RbnPaaAnOdTkiPhiDm9kaczbPI9R94qmS
2vhQFUuplkQtMB3vCoFwVnaOyNhuaxezQpRidBNJLaU1eboAHaXBNJMc7/QvDRuc
FHS3BeumQygQEDc53CBbExSdx4pw0ldnOkfviuub6A1fZMd1li9AbB56TMOg9osp
f+SNtK4g95SjvJr9rD70bku5dzPTOSAd/jTa57ym4AN62Bpjfm+95ha1IarJG0he
IdeIdGTZ1TbLO8sftkCCeGviexDFpU8NMl+llx0x5PdSRpiWIHFmC0d/sOuuTi/N
jFHhcq8vatKtDdPx0gwzt6m6YjVL/LFaV83BaKvhO9GyH5w/LmOfSHMpCjzTyqQZ
RWYrdtFIFCTaT57wNX1aaiVG19W/JzhBEIOH4Tniqf1LR7U7NOvGQV1bkJ/fDBBz
vHNhrXCI6V170Xzk18kVWUwmbvJpU04m6n0uujk11PPlD5EGFSPirxfLFtpUXXOW
xbSVq4dw9XGohIc26s3ylHyllN8UYf0w3LVZnmkVwW26DXSxY2zBAChBsdbnHxAn
7i2+XnEsPtWnIpB4DkAPeKDk7qv613E6NNPHqkLMNe7MNBNPi73yQo676+nm/Owq
1FBk/EFPEzDRtCHGNVIm/TMbKNsGD6moa9oUQaZj2UpYCfLb1Pohp3lzWv+ypFiZ
lEGlxg7uSoN/88NL2HtyVlXIxdx0bCapTpKRdQjnG/2s1fj06Q/MP/ptxkpQXfeF
IOlKaVcID1amNrENmd4Q8N0uTxnda0LKfL1qwm6u+ApZwjwsNfPnUgXlU3rTUHAM
Dy9y8MXQr/WKDwfnz0ykpOV+DAlJCilAXzbq4tTdL0GfA0iIBj5lhj06954dkPEp
5TlR5JSZHk6GiAZ8k5AKxk4+RwyeLqBDYd/RJIUQ5ZvlCrJcNZscW/NGd7OVLO75
J9cd7m6FAvD/xtdzBi0t180tVm97F+GISzQ3gKpzkxPzkGB7FG19rU3PjWaEGPNn
eQRBNHzlSKe1XEWZ45sCUsXWGe49f8ozv/1ifuRa16u7O6q4z3GlIK8BCH5S7KR7
m3vFZsw18n8QoqjqLdjgAR+k6zJar5kzox6iRkmCwanQVzz2S2waLBejlf4w4tRo
wUhoBwr5NNJGlZUc1ixRvmsQ5hqISokZiZJLSJezOskHQTpDP7kaJpVZSs7SEmOo
NUonkzcNrs7cexmPJVJmbCg5TeflO7IjPZ0vPMSdWhNvM6RGLyXVPAw/ZI+Xfmxn
vJDvYD2QKCSQbaGdBaI517oah8yZCtqPNM7jZ8k0z1YfHRiALWLqKJmP5AXpqzlL
X8lEhZzoZ+I0BGnjVT4A3qNrY0JZZlYROeqUnFbDdtuC4S4nTAXfLifGBj5PtbYw
9mHYG/e6+mSTg42BCNa+1NbGpz5QaU5FxXUS4CyNiPEU2qSiDFYkolzb8JW/x20s
GoU5Idbn3TSCPqx7LduW2++5gRXdfqeLncXA6AMuhltytla0EQtAaz5fnLFgfgEE
izORxg66VpGhrpYTGSCUki8b/D+7DgujXkJJbx/tdlggDy0Zyulwbfjq2ieEbPfv
vBVZeHOT3aoLyHGLVNzLIj7GC7yAEB0Sv5niWmgXJQIsTJ9mVVDtWlg1N5b4FTD3
J9rwLP1w/Rjqv8XVDwwBlLBFPocpzms6Fzhcy2L7L1dN9aptBzv4hcc7mS1WxDeX
lMVC9P/XceZorgVO6L1aUw8TDOl6qJOjL6+R0xdj6jpDV8fiz2P+/liTG8HbZTyA
mDk1n1ZWiOI377EXWj8hF9BP7Wvowmbr1Rpo0B3qkdMSntIGCZQsf76ixkCZngrG
qUM0Oc9K1gsmbI7siolsAeKRqQI6Q1iKuJobc7k3craDhLYqMwt5F8I3B00Pslbk
RundXB073ipH0VV3yFRNaYSAT1LoQTBDHZUbYCSSjJMItl7aEY16h8x1MpjgRWMF
czpNhZNnPV31T1ZtLkreviy2JZK1qTEvUIW+AtkoPvJcNoesZ1tKVM9k9WuTPcDo
A+ex7srnbU96hljc68thMOJf7Ns2z+HTPljRT4IYpNO6Ke/HuFJ3rYuZgpK+r1dk
PNavoS/wIrR/mOVXIEcylGSOxuhscJlRhbjRae4ZB4IIga7J7G7dIWlFOs7nfiM5
fqG2tHpEcyA6HKvkp5x5e/RA6JlFUe10d/BYuw6z3Y3YgvMEJBU+LZqNGxHiH+ho
KHf8BAmXLfc4sah8tIxGhaTT7KkBakFu8bchk5NJ3vwAxotjGv9Y8FNsQpDzAeg4
NiwCJWFqZTjzJWOgNMr77PLIDf17+nM/8ve1r47s9VCiidG335Pn1oGpl0bR9qAK
zOZLqwSyzzZdEM2Z0CWbv5ThJMi3q5aDO5ywlGoq5ZqPGGvjxJ2uA8uYKaxgEAVX
KGxoS9lA+8wWcMfTjLBmgIOnedZeRluPvKRRwDt69HK62nO59tsdfGnEtb6RkSse
J0v7lMOdLJGyDbBQw7xaGTvS+IP67vPpVPqWi4kSJ+zI+sRyxYvAhePAcX/lezAF
XqJhtjM3fFr6HIF86NE//NDfG8P8wiD7BrzqY9/72+kFLrT6jcNO4YNI1G2kEghE
7gLrNZfe+hb5kTd3LC6l7+vybbg/xOjcN7b4Y6pVEFhHFj0/N+APJ1XXJL4O3ox4
RyIMRiKRRfAxSeb7tyTVkWfycqSVxApfIwE5lAfzHR1m6EIar8KjpL9UnzpKid17
rYQXskoZlIkeP/ev9xqlEroyX3ujtMLdqYQqd880gBUriX9QbREU21Nq3QFD2xMU
CmJDEmFX/pZGHQgLcvSS14BFgrC2JCD6LlDYhOS+8c8ptLcLgDbFpiETfQZD9yee
C81qfcwwBkOv/M+rRqlmr6WCgpsyEQ2i4plB0J9nKimr6EaisH/yDPs7W0AhpjSZ
Wly2/AtrldEysoRnk54yFHoiWaaZXX8B4CjurcqiLmKkRE3s9a2VYW8SK+DNBuWD
CY0kV+nif/bwA5p9RLFiRI5YIvRFJoPVMl1Ln9oDWLHQfl5M5QPcMLRZFMAGovcB
gzNw4vvXHoHEr0B81HStVhh+Y6Rj4F0H34cKfpA1iKO94Vo3LYJGEAOfP1ZmrWIv
dtH2W9Ge0lVDAeNRh979MJEdDp2C7r5FY/R2dvlIX2k1QKxEHB9EghJJxDbfN1y7
BrGE3G1HUw1w8fTrlYZLbkOT8BXBumipwBe87PFU4Xt0KOzvcM6oq/bbqINAXaCD
kpWu9udnwEc5SgUS93mckR4TSO66npA13eAFLXrPInYIVFWUmv/t0o8qRltK+Ezu
WkMo7F+fs6boprQX5wbvXXlbkaaMM4jfUp2YIjtE0UtxcyeYcAAyJHXqaIzkgvwI
FUZPUb0jFOhzJBUfK6Aootnvx5E30CzqkL6GCRqTPY/XPjOA4YCZBdEZwLbfpzOx
Yrlwa/KiLINOvM6aj9nMSNQ9fmifDiON5XZRpGgfg0qQqCJ05ZZ6qfe/wrgeo5go
i+RjJzomaAcdWSu3DXh/nH2Sm32xt+6oiKAZIGyQSAJLNRXT852BbNOUC/6hZj12
BaVQYc/avD5gaysnrjUjVY3sVJTmIREZ+lD6GfB87poCSKQmlpsyUY6y6F8CkxOa
IcQfpTKg8xctuwiYhj2TCRr6GtKup7SYF+V2vstVi7eohAsnt7VvW+gyugUweAU5
3OQTDuSTBljHB+mCFXywpyB7X2i4zgVbtkNpvwvWuofjCU/i+zVfXONS60TRZJ6s
AaFTmq0IO3M8vVX+9wB/aHQSJfvCFG6nOO9DVbyfadY8g0XPDxlpon6+C0fsQvFG
cfNRcFQnE7FPL75KaO88XJrCS6PAB/QQFfOKri4CigPhtH8bk17WuA/2rSKTmT90
LRLyCLrOgZXCokMLMtCIUiI397oV/KJkoEMWBxuwXVs9UpUlt2KElukZaZMppGUx
mZiqX7D67ZIiKf4gtZUhBAbjfFCG3MVYppBow7AMbx7SuNxXiXEKSsc6BLrRLtJQ
imG0pcL/43ojAmJHrWDh8Sv0CYIn59cslpOT5txUeo5kUAC3b5X7WUlk2Izw0NxF
dOnIvg9NavJbzAPvVe3lDzooiJHGgKekTRluXgjgtsLkXojOO6fYwyXw4G/vIXa0
VLiV9sblucMrsjoBgXjuElG8VK4WoT9K/sWghL9UnZUgURB0Teduh6YICvIEE7hn
5CeDC1qpND3PeaI8NmG8+DLTQPrW3q/rDiwOpGgHwpeQl5nQxoSDgKTdBEBm3pK2
7kdsaC8Tu+ikLyWWnEYbCFQqzShT1Mk2rghmK6XPn1n+e0nGTwL33MG8hFIWbduM
BpgVqgY0x7bW5xeS2qM/PXpII85luhFcg73CFTiqkSnfVf7Dg5vB806RV0/fLL4/
veviJSMKrr0mUarN1zcd/BKXMZzWOYNM2NDTwD0jEergp2Otsr3spL/VAGjBWaiB
JDTPQmYwAmgHop/BkW+iC55sfDBO9JpV/pERQZcPRgnJhM1sIrS08gOW+vibsKcd
0Fs/+jQhwIxMAmkm2kaBC6bdmT9uJIlKKgQwqXnJpCDuskd479iYYpHEUSohk3i5
uHsdnhPY1kTIck6wmE4YzKBS56NyhHSb5pOLy9IHqhjnjm9QliTw0Pi++rKObylF
TjEitIA6yHdBnPEwV5MFXKyviCrWbPMzzD7L2z6Kwxf98UUI3f359r5425NjN1LC
CjwL5ITBjMv7qpc1mB8v9K8gXLgB5lFVgbIWDw6cfxIqw17L6+2UxSJkTHpue5g1
OKiYdXGPDVkmpjjUFKtPCj5v/0geqBzzsPUxEYXbNdc74Zpdcnu4pPpAsrJDP1ji
6NSvZtbTKGzxgq8IXqOaIDGEzRHzwXJbpsXpX3yVKaOW2b04dyKww4ACLuR12vMn
4V4lp2GdtUzCRwqwApPs5eDSJ4vmuFXrmScSu8y7d1OfBSWyv9Upj+QiJWXLtwJ+
joUu0qUx1xlDmAeSt4NDFOssV+YbT9z1AXzElZcGy4mTU6tNCjXIkXdlaw+9FoO+
55vXhDrEod/oozhbWqx677TGBt2WRCLJL51tkHCey3m/ZwJLU7sKDC+iXbTpsJFu
2kj+5CSkY6vAK+ZSCAMa4jcHyzgiwUuTu8NKS6neaOPA6ep4GDYQ4V9WCFusSG7s
8JHil62qU4/iNn5CGGJjWMt+R7u5+Di2dUFLHnMkNseHstwViKPiXvIOk4a9v6D1
jNJsPCx5Af3MpDipk3I4L+2AOn6TXk0K2xhvobiw5FO1ICfCz/qgcMN+iukQiHLc
C5CWT6kG8rbBhsHNsElrMSWSZUCH9L0U9IRn5cIUef4UL8WaOVTL05nr5OkWallx
8cwlKDeZk2uuWuwhlLqFu8StqN0xbCWeOYZk+Tf7W5cCp9MIkanawuQBohZdfyuT
064iIn5e5h5cu0hue4Ct0bYPU8t4ZzeN8Iih4GuGHsmiTtlxlmF0t+cCq0wIeHgX
bGXW7qqxVNpvbMRj29mFwB3TH76S1GVkmEKOtiGu3AWCkygziJIVbOcQ5e1Pghvb
I2yzLvsahvsWa7uJhM3RPmxiUdgzVcg6P0VCW3vyU4eFKf0bmIim4YZJuyr+mytU
hbpwImKu6W0skNF2Xm8SIG9qGen9hz2xhk6uOYzax4tMEXiZLSKbzl2iAoJdtjhH
ygamMgMHtSXOmADcLlW5zCfgYIcQsQPhwY5RPnHngm3wj6R6XsRmMMCv9vJ1EANl
1kbnQikTMPIftRKOAI+/JRCj4not0iBEb+zkJtSpWHnjTNbpwHyGPsO0uId6pTaA
Ul0dmu57v7CmXuLp/m/SRO6IzY7GftRTbYEqUgnLm1R6u/p9uAkUx3LLSmKisnk/
HcyJj/IoMnwWQe9ji6QusB+D33o8eZRHA3+KAZCbHe2+3foYIKs0cH8ZVVqhV2IC
mhA6fcAPeMBWxFhv2SHzqS7ONeekCssmODC6jtCIJn+WPLe/p3L9qBWvaw6gW8yq
YFsXwtwun+lDaa79xwUuFPdVZawfU54kvoSxoQqd0VAt5hN9BZ/oeRv7WsY9fFHP
CrsMPG2ns+ik1pilT+8Xr+h8uEwzdhHxZkUSg0u1e5DVdLY8yRWy8ZCi9w2NuWTe
vKegIzKLwgN4Z/0HveeQcCKzlH7wyURDB5oSfInkt70ZpylCC4f75iNg+hPQm0vi
YZ3DIGJB0j8ruiqCi6W6cCGo1c89gvL1aRaZSWWhSKedjgc/8ojwmENdJ32Hl08X
XyuIYHMYw3W13e0QItKy5m9GjbP11yMsTW55UM1XeM1eowVDtpp/19VoEPwwuGcq
S9EHYaXYtFwVNfXZbSOBU7RRILmeJuphYpUN/5se5Ft6iVs/A7ITuPWW+ufyL0FB
llIELiKbYOFs1l7Og4hQvs2ykJTIs/7ilvzw7iQoZtx6f0/wIlWa9/FErln7UOCs
bTH25YEMeB64KX++AALL42F9daaibqdfYoj5SgveVmSMQszFsYmyQ5/uYV+LBJU2
eC/HGPAsCM3vzL8gv0ViHqLlupaVEM/lE+enwQyZ5TyoTTcJncmHFHeNhau58XNc
TqJ5Vpd4XNk0DP0eRpU1ojv9LltvsBxdd8eI2XrM5HYTNOb1huOQ5lwQovnxUCss
kDgLo6JDvlMsZtivWE2M//JuNQw/u3WS+8KSB9/dWNNhfkyPx1qGMPMtNopqoO0h
fqO3eHrb1cuTDpuutRXrQtFGFf4CCfAJvWczzmxZtAoQ1Xriza7dZ67CfTpztLZD
P5yGYVSckIMUcctHRX87vswuO4jO2CW19hePhXLbDDVsfgDUDN9R0dCnQ+HPwVZ8
YAZKb9B7AQZBfxJMFQNyESj+4z9IJtVJgtBryDiMaWH0ro3KZzyA1Y+vYEPeYjqZ
7MbbwfsffwtbxOqknZvwytqYNKydMX9Qv+B3/rszORADIS2/rxMAkxqXUh0G7h82
SUaeaDGYAo6Acs9+0KCUOKiB9ITZLODK0L3Y10hckiydmBhbTU6lsqoiSztKtKCg
YgEs38BX/PD/EFRQvtfYWzwMWsuAjKzHMIOyOdskN8W/OeC+h+r4k6jP6FvkE244
F+4F7/+ujUz1hFqxHgIijvO6XLcQ+HEpdYaN7Nd7tugiDpbNhsNaWqucNfneI7hm
01jfdqDjax/hPFtBBQzFSuIuTW1DIb7PSdHNP+1nUkvnAD213ifWZR62upt0l/vs
fvNZp/oJvXtpVW/7ibPXKNFM97cRIugKi7ZheeTd2x3urRGYEKiI6hEEq8ycPzfb
wyiiXn0pCz1TMMq5Zuks8dr6xWsEf8JOlQnXBDAccmNAwLBnQN2ARhFWI6ZPMW+p
KwG3NJebj5V5BHOogQGk/Gtk43DI9NrO90lZ+sq7qx/+axj/qyCwGMLQvzlcHXPB
M3fq/JSNbWLQM+/zbUVkb2oKpgz7gXOZCaHD4tfPIwa/lrJsywYz21QcMm6YfDLZ
E7qlolERy8cmSOuXh0Ug8XIBJgRAZbqHHkroFkAQtwnsdzb+eNovveLj3mnr1Wj+
YY/OOq65Zp6lSV5sAzublM+WWb5SsadQiEjZvl93MjGR2w6hQi1aJIzyIJJKi0rc
AzhaxYurUDJB95pYK+gPTaQkCjrL/KOTLclrRrso3ZLsGwsiWhIJW0Vto7R0gDLf
Egbso+yc/ZasWU9DEQ5pMgRBJqSwShNR0frZMqDp9Yphp4Mhw+e5mOlNmH1BF28k
HuJaB5PxCTYNXKV5GqoGdkZT8QXUFu4OzajsEQD2Vnz/Gdf3CZW4pjC8LZIqNvlt
HjrFfnFCM02aFJ9MxN4otUeYwN8+AXG76rKHcMLh+q+lXN2pRwGWZ7pHzW6vcTGi
GcJvO3z3Hba1UwceJ7bEOLqDDs/FGVPBy2l6Fo63lDBniQ0Rf4LMqPFsmSjBxp4u
YaFAJUDPPx7t61oVQX1ZCYcTnt3NW4qRGL/6l4XrSI8Ce3ESFZOcdXigAj59Crwp
ClXkr1om5wFtHb7K5YtNBPETcNC8ZPQUa2GrwU8QMCnaa6eRLzCYlkZFEO69YWmE
l3ZVByKC5DtUXT0HqqOz6YC30bcGP1b7QLeAb81QlD97JfRkSQfWUQtJWYdeaap0
ZOhfBs9o0jpqXbRysOM7t1mxHM4E6h9fbCPuvq3S71KCuzxd1FiophqN3r68XY+6
Oz5t9WT8SXSVA3YSGBUroagX+3ksfydsX9+2aZ8kZGGdb8GH8kFWqG0+iREIQAFc
jbrkmg8+NJ/EIOSgO4z/1+SWejtrAzQkmCrYQchPc2C99R5TCW5w87pgTDcF711C
xPRrKw5y34/bKrm/tq+RgkRi1jHoHNygyo+DgXI0DSR5ntobeWOIqkF3+B+qihPe
kavrXIUCIJpb2i7CmPzPDJceN6uSRoDSVL4sJkdA4hyaoWgI8szdvLXvPtE0MgQb
jQiCQq6xIVbbqjJnCxhrQwsPuPOUThifPPdQP+DXch6BEUl74hR+xX0D7d2udUMG
yGZf1q1/CorJxnQ/fmDckPeRE9yRdPeof8D23Wbn6OTcL7ObnvlavvVPeVEUKKRJ
OS7crGh6F7o/T46ITg8HuhuI3y2l91CB7WKGf4nz37JNy3wnGW59/Sl/AUWymt4Y
jAZnGinPV6d/X4oXohbw3TgZx5dKF0wjwh6334KM5a06cohDMPx0VkDhrlozP5Je
q1Wotig5f5gYw+cxhy76z+w0Kj6A1DKD4pPLwK+l/vqmaVdZHyCILtdsDoQefXVu
XBy77PNOOnDGQ4XjCsqth+BwAIlbjSPhS7ggIqDEMoj+bWNQjDz3pE8W42JL0qb4
OuzXCsUHHtoyPvchbbDvkrnpbQa1+9dzOx8FjM/tzoxv3A5nBAAIH1mW/di3r215
IG7ZGGCEj4sueU1WLVWK5wsgApc+k3T85k7SEjCWRJtr17+pkVuvNCXlgKRLmew7
QzLlvUXdrakkORZ4wOr4+5d+mUWndFY5dMtDN6rbQhtHawnJV1YIUgypD89nvzQz
NrhGXtt06IoPg9W34DarRWjXwx25kShuYE+BrF1Bm2Yc+LbLEavs0SfBQCSuO95B
Mzzs4V7qwQvEywQkbhbXi3kahBjdOIPV3byeo335ZG/TEK5tYA/cs5ozPMOLgS/5
nnZ9AINj5QCRVfTfwzYOo6PYUJPwFGCl36oQvp3jE6QtHELgdeDmHGfdnWbyLryx
MOfdL3u91svoEL+ID6VsDqmEXCjI71xdfFIfV6B+hUuWNNtJpQ/TUGDi6igFVb34
B77AgBI7lkP0oHteVmJwR9IG0STyUrYi0G0YmyTmhUHzIrLD9WEee37s5+mSm3Pn
ywt0KehYRkIXft3J7YkX25PvFSv8WP6YoOQgbbwGk64NvHN26JRUZw4aTTTQWvgU
ARruTFksk466uLpUtUWPKBgxQNYmsroeapqTzJ8mPRhwfEnwuTTc2mV67fXbjU5R
s7HudfvW+aLqjiHpu9Zv5kwV5ld1Ah2/7Olqmc51u5Q0bmZaaz/abxbC/k3NL4l/
BLU5/MiFJXr9d3PROJPN0Ly7Dm37Ac1ROyPNQUEsWsjzQfgaLmw97CeNYKepxHA0
t/Dtzqs1cUNuILL0z811w9UfE2dvDlQsyfTD02LrU0bVEnrBslP0KXYtgW2YDK3g
ojlIO33eW41KWrL03uBG89H8DsE6cTBWcd2S8ycc84EIbjotI7h8/Ds74tWd4J1z
8ZDwY5ZEyNjVbdxLZ7K0nMjwScbg5p+7gSB6cmsCZJgXC3dRp6IivLlmfAD/Kq2j
yBh7cxr1+OFjMxf9gz40WHd3ckYW+P+w7jqF+j30kZoGtdKHCs3MgSakcspTulSX
PFnbzNic7J46ZSm3PcnosQ/+UyxYpLj3jsFHqUTZaBZqI+30Pi7QH+qawpD/Ya8I
leZPuc2YK/dtzu2avIDgCDYbFV8SYrFS3cqtrK61ZYWwNDfoJeTasCqRrqmys7ZX
zzePbxSpvPpN5N/KMsc58OMWXYnPFMkMI3LIpO+dG5YSNbch3ISvFDk23s6L7zyE
0XXU5rEbmWdcBCKaA3WhOpxEwkvB0ziEK/bumv+1ZmOdS7FtGTOWU5rX35tztzS+
xOncSNO+dzDb17CqpYoi0qw4SVuBLEewbWigzEVQTmWpgQzg1t3riRku6fQIJIO9
iiCwFBSv+qZBmzCykNqhVs97prp/yVjhy+cmHEz9yMJIWy3OhKcKFtJtAyHfBb5d
+nF3HDomUOJoAQpfg7oBT1sRPBrxdhXtCgNgZbx9MN0aTo3uKOcbGjYln1vU9KH2
qlBbtbCfUre5epPQSfJ9eJ9Qdu4DkFg7O5im1/N/8FGtFw5cLtsOIrYs6bkGWmqx
3wdubFUz4mdPouoiSPxYf9kzZTY83UY8Wc0d+25EY8gYV8cBTIZ+uXVPshR432C2
O79UubNSB2Av6PjRau458jljaz91n9h7Joq2JgCRDZ53Dn5ELRW0AdYBW6olqpxs
ebUe7DhtDzKU3Q0ez1kw61KPPc3AwD3cgg3O2/o2oehNu0xCBBBIKnaXfB/gIGr7
NEQLNkfHT8Y8nAz+guh7mF97V1t1E4gdasmxo7sVLjUnDUQGV25GKlAfAu0UlsoT
HkRMIawhmDaUwik3XkZd45aaISWg/MtxTRtbpQdfpeBwKgVgbz02GNmpc4elfNe1
g9RR0IHH2gEoW4xK45KhrTVwHoS0Dlpc2Ui45Zv5dDwI7GlEsCh/cURVbkcCtUGm
aBOmGf/BfrIMZr0jhuI557ftoRWSCderOs79A+ZP3AxXbV2x+9PJn76JYWc56X3E
qCosQfaeVch73S520rf7KW8oO5co21ImFyzrgONisn4ncKI7TCC9FpmvHSr5ocHW
GawhaZ8F9ENV8b7K9ocWcOxRY23AQ+3zvrLa+oloMEmXFmQ7Ygh6xSnc+uJ3Unm6
x1CTt6HbV11upaWsvWgC1hDEDjD2JgvU6QWebdYHUuDQvP+7UvMXL0XSfH5VaDsS
ZG9rFjf+pEyHvV3KWoakFL0ZGadfVOHVEyeZXQEZsqHAz+KXcPuDN3drSr/4VjQJ
x4RwheGWfwzOFrlD7issT0/kB7H6rjtGdH9oySQysosHnU9NHsWjmzzKPz8bjdp7
1GvcHRib72DGWf+MKj+64Eb5CTrmHYw6YVB8lUwLYGn468+2FNvduRpmGXDCEAek
Y07tkM4tvXxyBLL3QRuJyhuECWuNhxm9cVmc6MMh1GHXcY99k83k5ZBxL4X9sj9y
T5MxFNH8eR1IWMhOiiUnL9eIWWdPLPFsciIxPTmno9c/bRuXLeDOb06TPesGFEbE
qqX4r4H2Wq/VwF3XvDMNsJRAk+Svv/l/InRSOl8xuUWo6rT7PiROtBI6k4JbJiIz
jib3rBnqdPldbq/gNVYCEwcaBmsv+XTZYiz6EduVLyB6zH1KsdPQp6o3SkIxFMNt
qouiDmy1A/HATev8BENXUJxvKljQdKxoTLFzPhUWhV4a7G3mpqA5mBlGgxW9+Abd
TKX9fJdQwVGPERDbLiZ0fuyzqk7v7tu0mcKuhkdr8Dgp7A23NUFTJOXnmMcw5DIE
BuDNPuswAoOjJfcrTm4ZLYQK10hu0u4vOUBSojH+KfDxGHQT57OeAAsMclD8jc5e
jJIbSUN/n8D44NXPArwPPLO5H0IE+72NXSuS9N4w0VVt4B+2IFEG0oD30fOjDFeK
Kf/wKKRN87cOg7RYbvejnD9Avq+QDGMXBQYdGeYRvHkzMKtoA+hQx6vZtIy4MSit
0seK0L7JHvU7Vnt1g12CH43+sote+HH/3nIiQpHG1SKScn7TlduNgdgkg1uEUxFj
Y/HS5W/RjbJEai8vSyrth1GH6mOFujDFRGWT3nMV5LiqqS8fWbGSUgM1mro6Og0C
+qAPYnNg0DQhQQQbxicIJVRy7FcLd1+yRzzTbgBcWwYTqpPmBMX9gDZ4k1XbRmY7
uKYMQFZPUgR3tBiXt8cnadlAfx+KW7kRCYNOYHmUE9nml6CUSoyOb+IWg/EMOBnv
KyJsAlaK+BE0ed8OSyxRyyySbDLIGCnYcQUS6xLUMMzrgGpmz8O/wk9iFmv8t2G7
yQ6iVtHARuPNvhCivbyQ0XCo5KF/WqY/L277toSq7xdlj0fPd7s6ThtdivuEXWmt
6Olp5Vcfp/vSLpPjgpCHAF9aAfJH8/cNXIq4f16RTCEUSHXO0GX4JTe46QbgaBVq
PnjMZ8bE7Ro0h01/UwnHz4bWUSYw7x536iajUL9ABULq65fnJ7XtCJGvSBk6qxRg
v8ScL4pHhm1SosQDxInAIq3hL7M+2/EPBsRU/32FE/vTeSZBz5ZfzdYThDr9sH54
61q6Y96czM8zpm6qTHMSn2SxfNv/n2Fb6EaUQosvjsMCOUXI2RtU8Frdv3kPox+N
lRLzoLhrIWIBdLLmPJLbfb4IZTlNJ/6mroKrB187FXVEwuAukzc1uBVcB8SM8ean
RI/viXV7bHW+oSb+cK/t+8ddZ1NSlq1tYxIdYjuJZkyL7iGs0fzJYe1eIS+LWDFV
caOKIqyCNfQzllSZi6igYf66Ql0nW3B6iijk+q+RbobXw70lUm7v/aJbx7Ob0JUC
65YWD2BH9NtaufFqFddk0aIUIpY0cUs2UiqxdgD/V3mSKb7B/zGfs828201a+PCg
pFp8JwrbrmT2ny9zNgGORQ3P6jmGKrMq501jH5uKhu+F4+Ytk1TiZCIFkx03dCbZ
Op6f8r8bKEJcDZo7X1yneT6B/DqUey+nNeiBIgQvEJiw9jPg3ml7Sq62bKbpA1By
tP2Wl9QqelmF9mnQbk0/UpBASwBNV96lM3Z6HSxT0c0eAj+azkNTinC9H9WXTZmf
HRS/xkRjZlAa+tKCptNRLhshE+B8i7QlNXhMqzImkAA09t/yfVnGSuY+fQXoZKvc
2z3l3mtdS58lPxjEkwMOCMkZZT2/i6nh5/yCusJ4FiIghmt4oebARaXswxA33LHN
IkyBqymHUvt5UieDGnNC3nCwIQajSSOH+jzLhuPLlzCOrMmN67wYKke+0klEXbxE
hE4ptfJHODsSqmx0WPcfhvlqu4GdkDxdxFm7f5Rt922n2EoRg/OAWfkyLVlGGCyr
Sd/holxfPdK0xmBRbtevVlNREGCkzfBk7UFxFMNaJUVjFAluZlsXscUP8tcwjfoE
T4eWjoZ+puLzB+VU2U2v6fjQodkWSGr+d0KGi1q+erg6++BGC4Mt+4LZOuU0XSqg
t1yScW1G9zP26csnBB3zrAmYYxybL5kuIHA/W3xp5AOPsjPE2Z3g8VFOOUVfH3vo
NbVDeY8LsyJg29Hd9agFR/wxNiOkpi8lPvk3Oq3MVyzvZS4Zub/AqzdHHzyNTDDn
KHc5hf2YYkSRNmVtga+wGKOfP0mTcezaqQZUsQeSDdlmb2Hw81qw6Rcwqf71JiY4
wvlia8HzF6pSryofkTA2/+42F59YXBfD9JUOQYLJ4DfmvKO5fYL6+0G7gmtwxD0P
LBmMTYcPa1+vdhkPrp+Zf7zr1CYq3EEA88T79qAkq0nV9TYk6QvKteLHA5a7HYHJ
ZUtSpsYyKWTb07os+4vBgxXZuB3Nt8kuguUtk0Si+eLt3CYuyikDC1Q3pCQxt93N
mYsi9CYoISS94zehRAQ3HLMLoKogoYxVbcyl8e7CnM+xOq6EYvRK7tD8xRdI+QBK
oI7a62rAov7SqBA6ZBvb3FiqQH+pm8ySyhteK6VRLBfWn0+dIRRMza57J/V43H/m
/4SXoa0c1AFHUCxrcoCLKHEPOadlwgYqdevCyzY5E8aAqJyXCj3c1jl4qpsvV6Lg
Sp2wSj8zatN3O7U/Yamoa0HX6I/SC+oxhO1MuH/utUfDuDOtVuV05ubvUX0CxY1T
VZqNDtE2rVhAhdS6iUaCqcOgxYKT4akd7TEzFPaVF+xIEHoSS5XtBuMnAbkNdmwh
FkuxrpOqppRArfNLFJaIIgAheXERsDPQ2wIn4xRyZ3JIYVZurQcq2FZO5ePKp2uw
ygu80kSORXN+N4XgP9zQKEbPOTAYss3ZcQ8lCDVeeljWVMWqeDU98jP9cLMxgP77
UlV/O6+9bIJXn8Zmqzzuy3ZN/vmus4HLuJFLvVuu05ryNjD7lbIcJywbmN9oTwX7
4UX+ewpyvKC1/kADlWd7uXCSVppreooO5ie+WUMX9UwttP489Tpx/4lFhpH4J2Cg
fh0Q+EGSRybUymaVpWsIcK+zHgIQsc7jweoAC6K/+9NObbad6ilnwnGeBaiBWLyH
2X8hDWd6O9IETNovMHSglUr57//TV/tgOi11EXfH4yegorZXnH/0LGed+D67jGc3
/LgR4yh1U9EW/8zynlb30+ANIUMz/79pDiaD40izPHEoG3DDIWt8hqE3AMa+3D2q
GT9AnJUISeOe5iHX0KOEBs70pVdrK1YkBtXeSPSJA/6WB2GRbAuAtI2QEkiyx4MV
mDVY+LJKWb9lby55kySHLZEUysf0552iO0Hic/1CmQFOC0CiXcEiWBxKaUJyp8Qh
ERf1nR5d78j9cXOhNZHm7lv2b0j2e91028xdeSfbmLQnIyMnWf+RBrscVeMUFIBM
s5Px/Vu1j5YlsK+8vulkbQtYRx+YmGeaRYDHTktV+b6GZxZ/auVHAJ+91QHyB7ub
kmVZFGSy0Az9MQDFq3Cs4ckERegZTjR8ulIre5ZDeRD26/+OvJZu1XN7zsgWBdDn
f2JX51rljb+2EKasjGt/DuzxxkSTYqGyBeoSHrBkUO18KKPkJ9G95H3CpteSg3uF
LxBOB05AffTU0x4m610O/zCzJMnj4kNXkYSZDU/C1x6XVMB9QHNqDC7zPSkt+B7l
34faGYWQyFkgeV3slry0VkCSG+H7kvUAtcWptNfzeG6F+rRy9lLvIMdyFESizie4
bju1k9mq0fhPUrPdJfEGNqaEdjB+lLV9B/8BDhQVPyPLc/fUPRUxkjmwApoOIj6b
U7U+wokkwL6vjcL2oi8LYABoFFwgZIJMOncUp43TtrHbWNdtYgTP+c+ymH+y2pAk
d6EM5wBwGT3tPZCHoIy1dreLWkLCFSOp0sr0FA/pgCtXlqu8JugkHNeL/PVzIOyM
IuzQLbx3oQWsGaLGUykVFcTCqUC53X9PQTJ6UX1tbHlh5TIDYzRXlykcEgATAcWM
qu3OdZTuaxrzZ8WvGBVvwcvYJhFsnGLQx7lyu3cfKLYcFRYZ7e/lAUbapvsSa2Og
LdTmgw3IVkLrMYJJjQcUf8Uwnzrj0AWA32U9szEl7MVjyMan5pRdfUBw5XptccTt
KfUwgJOOBqobUmIPTP7ZxC3Xwljw9U3OSlFBbWLgQlBuyjRnJA85sPfORrQC8CmH
wNcAFgjlszfuVDXCxMraWCCqoxYmEAbLW5MpLy740wfa/Mek9rK++GvyRzOllCh2
i1DJ5n0IpxN44XMmWmId0GqIFEVY+IzfRh1I6VoMoSMsY4UmdM6e7kSoVtD6WoyD
dqEq8I6h+XPrMkzyWRziCQw078eNIWiIS1E/fTP5IHzdNqT62Tu4p3EHeahDxIdj
4UOhwpiHqY7C+ztYwaPoM3njVgb9uOm5MeO5hZ+4RZ/NJY5h9phlJO5QHw/qnryK
lLBne/KB7B16b2dR6jLFRi7NbHoEkVYJmour4COKL3B4PrNqH4+sRmAg6+ZJzn05
+JDu1I4Z5rBTRd1zwjrgfm/ge8d9FdfprVrSz3s+1Aqg6fFDFRkEhrIBmte5taTV
SceQLVAcpG6aJYJSvVpcMlHFMz5X7wcLlEwV11jz3mXlIjuyoxx9lVBZb0XZI9mn
+507K3kPUOUnl4UwqIBfyPDxsK6gkttv6YBOn4FlR+4lNhRElJwDIT6A6ASETiO8
4o1keB+D/GmYqZIXJzCxIjaVFwG+06FQ40E9mrNcNl9jgKnL+E/oqmi7Stw9UDTe
iDfG6kKMoRdXJ52mod7k28C4T59jdG9l8SHhFigXEH4VBNh8xxlzODFDx9XjtV+G
XaAvDWxvqldXu02mXn7QoSkoGEtPDAYBzDuqwtQZA7af9tEzNIw09lh0rg0QjYes
j5Y1BOj6Qeu3D7isfEkFH+ftTxujGIWX1RhwxPEuPw+aetRJ4+px477fz20FEPuE
AU2fh5zIaXAA1QRy59ePX/zpjmm3JUv2jvxMpTr0fHiDytQI7YmKOvHQf0j+45vK
uIUDvaJdxMMA4aoS50WyUee4bBWbCfwICKGiBU4tXdnw/e2yEymx0p2bpqBVLWG7
CWDBXLxbuWtG/lPdgrml8+jTHnKD/dBz1EsPtpnR+ddU9EkAhvkD9os3lJZ6/khV
tbVggAuR0sjhdyNT6YWywjmEfcR0Imu+0RRPfVhIhzelPg180puifWxADDPlEjDN
4Ko/YFDHrlqwd16Hg05F4RR0CtRJuDNrXp09Y2CyOVhgkS9IUpQ/HqgNxMD4lCzL
Te5OKs+oEu9T8QmZlj3YuGDuXqttqLChpkzwuhPtXfMes1oZzq338tDvhOhXzLvw
MW3LiIIHxj+IiJ0+im9Mx6Olao0a1eGID/j8HU59wz4ROcX5e+vsQ2itH/rywT1f
eY710v1A9qzTZqeDkNy9hZLvilmQkmK3agUUm3vkv1l3ymBlve+fO6tauPe5XrSu
aZEbOTeIwalyziKf5CWNkNu1eRDbio4wQyUk3X6sVQP33zMLy467twqifmKrG72B
dgK1y2uPgr6vxouha7uQVPjVwVLIuA9mro61bq28Xs8KX2zDIZn9RZCfsRk/HxW2
l0+eRIupVLNPE0IC4wpSKGGDkqoL3kLoX70P/5rauRLccUBi9psctZx/Hzuf849K
zAI8GsCdJKzXvn5V52OU88elHcG5asiUTRp1lxeEtP2102I7BefDfkoxAp0t+DVg
bH8RAd6mzNLpc5nMEVkuevP66Eay28tY3n16rdXj/+FlPR9chdohkRyeKv8fitqP
mQdAN/CKOOQ4gcFPEmSQyF8jDGTRw27kdr2m3Q4yGI1VNHJlSsomQRI2VcVlxTx7
QUvg5k/4kqWyvJRjtiE1pJvJ++o2YjGjPdn3vBbqVxIUCmAA9qO/I5ZPo+0KhT/C
DKQIPOXXfYKFbBNcPFVeiT0XrQOPq1t7amuXHurySs5TdHQn3+bwN+IBBzL7JpWJ
VV5ZJbG0IA5WBQpanvasdjhKrTQfBkfJgUnCDA2deKHN9qmgwzur1Y1ZtUlPYtyG
fV1Int86mi/aUVQG4CoWxrB71NO4+tBOT4sEMBSCoC9eTkHiAwa47yM/Z+H0iMMz
UxpATrA2T1OY6cHiNzB7ur2EXWYjdZ/5n8XfYJoA1rSoUzziAv2WOSrlOU2HJe6Q
9j4XLMR6ircj1i8yzbOLRYsmtP1uu/DEMvq7bc6yJ6tEShce2BXHgXwmTdkBg7wu
P4wd2zLutPdkY36xZjH/gp0dSb9IKzQ3hKDRV6Heqa4AXo6y4gwn/viMEY+7XECx
5B8s0u1NLEDGaVphoPjwUI4GstRG/03b4Pw5qS0p5g4hxfHYq2jZWKdmEkcFa/EK
jy7Y+XIExtQ75LJxzrE5kHauuG9JuLXDBrYgrHabfQJrLZJ/5lYqxA9KJASLO3rX
EUFfA3NlesHYM5yRBV98pSbVRHGbq6+TvWyo1y+6Y0X68jvXZEMrg9T0Tv0viE6c
ay5qYfEnGTMdlrJ7z/wZ65779qd6JlIsWlgNNfsjisIkMkwS4gYZw5gOYMOtgtT+
YBJfalMK3FKNqYNrJo3hRSUXsZYM9TAzjE/+wIQ2UfvKGCO2CuOVISus1PMnZv2u
3nmwv/exVOesLb58W+EVKMECMi4jgORaMm2AGwXVaZ7qbg80BGMGjsplHBmUrZu3
CJmEWIrN2ckomq2LUTknYobpmQf49SE146bhpv88zhgiR1nvZXOfERANkzL4viH4
LA0Nw2fqLTdmIdcWrkvpnYVYyvkPG6Ngz4+d8RVlAB2/Aa8OxYwNEycB5JXpJEwO
I4wUNf9VKHYOsiWRhw9P9YKx+C25ILJ82rtGAWFCcGU9i8Gc58Scn8Nh21+9mQwE
91fWtVbU9tCn9Rp/gR7XL6CIdI62iPCh3ZSq9IpzRePtty8l1JvzEDPcWdyI7ZHt
5NDmuYTPVGOAvx2QOWDrLYK6wj5LkEasLcBLkQPhjMmvAi1ft1EtPm1Tfmb+mJZj
NmDtC6zSxGbogmdXJ6OamWTB6lZUtMpA9HJbVzljgbcSsYEMHe7xdjj/mGKUFBkn
xwK1gxOLMczU2Q5OLTw6mfqUmCwCtvJEqDqa2Q01MCIEbKQf5I0BZhvRn5A9DEDz
zPznhUnWCeZJimRuq+OHrqkaB7IzP9z0eHYzQJccQWBcqzmoISr9HevyfUiULdRw
ar6769GB8mYXehRjL2DdVqIngjZIRU8SMGdAs1WVDUkTEorHOd6d2m20X1mRrYwd
/9LnfWxwNm++ARN5prlnOLAFYY02tdY/TDEtl+6lSwNr5dWJGoT0AhQLkyYQALHk
TCw9Udvuc0FBYO6063c0W9D1ThGBu2XBoUDbT17lD5gNroYTL05OSg1utPm7UzBK
GKgnPtzBYRNgjV5el/vzt7km4WEbKfSos6z/EkE+M7MH1T5pSK9ecrpEcxajg8+2
11P32p/G/xZdBUBvJCJtcMFF8Cw1mBRm+XRYDlWqRkz0bFcSm7fgUK2bcOfN03s3
jIKN+8pWvNY4CDPMimgnzFfFb6L3YdskIY06mXi3jDkMzCehORVIqFH0lS6eOPb2
tGvhbhi+I9B6nVfq3e/Kih9PfQKl7hee4WBk5hSJDhp9R2IK7d1x/U+yRMrkmkX0
xG9ce573tug46Ytx+d/9f/fxVbWvKJnO3kOnVqCFb7hPHx9yeGsHeWJrNOjQSPCT
nkNr5Zr3/bUrhLZnQzXWSLHTwmTzR+ekk8Hztsk6oERLJPsszTtl7MOEvE6NUT7m
Kb9/yVnZosrmJmEBxDxyAtErFyoBcOdE8ZO6YAatLVFbGl7xYOjX0YpMKijDY8rV
OqcK1NhOUSx/O0TmbqdSGX2y0aCvM1BxLf3vGyvVwM20nYG/9MKZV3Yljpj2U3wx
2KTm+oxSRct0qvecs3lvzoM9RThk/x2T0DLu1kl4lF4scP/8ma6r+1KkEqEXkMF/
USUNyUYYaQFMVY/UZNK5T8sVpSPY3lO+z/0vKhIBCZTMgGFcqyWWBfdEjqxbXOjn
DwD7cWcdj1mgXh2qrTqpTZE8U2i56nxdv2EAYBqKg8I9065ElKABVJymfzQK8L5q
ZN3atS49vNEk2kcDhNa+jGz1J+8RVoUrafBGfgTL5RfTt9/x7koj8pk7u82ozz6r
AX9si35eWBGmvToqEX9OxOZcmZQTRVZa5mKdZ4GYUFylHhuodOVSkCsJqPpncZX7
Btjisyt8ZQmPAF72XHMePEw1gE+wTKIBkahunuk9vzOUdq7sdDR9KwB63eJnqOZK
1cKo5LAMywgua7PhQ/n5yt39JQF6FJ4NZDM6gyQnMyqRGOlmzLNz+O8gGGfLAW6O
HU1RwuAAZLDIQkd3OozBTEKOScSIEQg8zQ9GESD/XTmpAbXszFPETyP8AXDazdSJ
q7BoPfDs9TqBuMPNogyOknVzOPbhKOR7ZE4wr+0SHDIDpqC/fZppVpz9VkTNNuz1
uclsWxuFF0bFsa1pK1nXN13qIciU/ZWo3r8nbwvdxpvKNp4p3MRcF6ycV41Lnuhp
XyiUqIqPPsssECiymHvuYRAmw1AhvrWM1B33BgpJEiK/JfzPZBl1PD/V+BDXEDqo
+Yy+mK5g7ayC0GBR+omW2jW4HtJ7ZAWJGaL10mjp2EGnT6UyrXn9rYsMGvlQXpps
KeqHSQQ3piWR5Q3DsuKpip95xUDHJnkah8pNAdSNXaGOicthldP5tpMgbIlBk1X5
3gwrD4I/TUkqlK3vyF4HQzmzxbsPbCjGOtpHJJdKX1td3S1PQ9QMVFAeWTmYX97r
0DWLOzcBAneMtcQ0YDsh7GlUT3ZG1mMVfB8tOStd1juV90SuWIf2G1IJzIusVy79
Z+nmI0kbAGAmQXzhnjoRGbeCUKWz7wfBtHzjnNWfcWFmFRIYqDpI4nLmqnfdHOm1
t124Jaa5BI7xmYaP65FZvo6Z3ageu4WuawHfkmayZxNVLtAzuorsk1EpN5nmVYBv
br7Vrc5GU07j3ZEmJa5ZewugiyqyVMBhhMgffRiiLY3GvJhSeFrGvQXoEwI7gZlP
qE0m6YAFj0hnEsXGtyQ6zqF5fRRVOin0y5E87T5AzlI7lWy+PohdChBDspDcgVGx
LHun41+hUBrltIuPBf2PMCTO+TptjQa1AMSFBu1sm/RERs1qrE4gdggZijeFqdaD
uFN+1OXuJUYStPKT5S3IAuBXCnCBHwM/p99uShU8uIYluWp2uVy2D0R+XBFkLrGh
u99Y9k9t6SWQDO8Z+KESzUwKfj8FjFWxM2Fpp2PbKUx5FeNi43BJWoy5oqo/IS5m
C3uLARTJpwjUgN6V9FlrRVcw9tLQ04l0fB8BKKXMLTNoUWPogXqS+10eb0Dl+Q/+
Dj7i5DLMD+uYJX/RMOF/tlw20Y2zLlJXPE8GvDNtjZNVLFvg9o1sBrV24Xe83d8v
FRR+L9zbPBd3DLc6Q2zvEGgWAx+CtOcg2NelOP7O+/td+SsdIzkKXHBa7/Amv+VM
kziJkTWylBO8P3ptZV6uAqcp4gogDp2s+BJL1mD0tHLpGfxUfj365veLEa5uIeR2
FL7rFAvueDbO8OUhiVP4j/5C5q1kfHK8zbintPjYz0z2pZRYllijwLXH51hJspi1
oFCI/N+0SZHLoPtdiTNxHCej9X9VC2woGLaTjaQMOhPm9TdANTb4rRLGiDNoCw0m
wve3uFBE3h2kEkTr/nNcD8PBY52YIUKS0RLVgl1RhAV2Rs6+vHd48mZbtbm+NY0I
ZdHct1s3hGth+IZSPNDaR8DQkVQa5rB8ZJKrU4mbm9CeaUJ9rgYaq/WxFNIELEAw
b5mkeF5v3lF04/9jKuEDohuHjJgw/KOHaSpR2zp01eZZAjY5X2rlJIPI5hDgMBuz
GggCOm8oJtjNRvAxYZjI346TATuSb6i5D1hjgsUzv6lhaym1SJDFXbmUyIEh+vmf
5FYrG1CWzznrdfi7S/R+PueADDsRCSz+Lr9jAf0N/lI30EOPLo7Ylst87DXTYeWU
0nFDRuGhVg0S+4AHocy9ahOwp4b6GbxRwScW6ukPib5ZT2yAGOt34c9Ty+vBat4a
SKfuXWpUa5sQnU8tRLQcBbWDstDzAWIBvdK5CCdztCw11/OnF6ifphJ0QTi/ORo6
IQw2cOPUER6v1v/X+0m1Ug5gRNsOyG5VGT3uRIZDUFu48WwwFIn0GdQWDkNSHav1
pkuyYnSUVfbLOE76XlNH1EXKPpN82lG4u+FubgxUTNRqQgyyvTTjpoY1QZNgJXVl
W2+ttMBckolA8LoghCOquZEj3zM9y5ZBr//p36lLqsNJoSEGx+G9eRvPyF35Pc0K
9FKazewmVjhCLcKRFrVHIxMlZpc9NA3hTJkZWqkXP9cI3KRNR+fVFCrE78HcO1qC
8ZLraUvO/UaHijth5lZNj9IZ2C9BAFGZjzxDXuhk25EgnCITUS15Cc+aulEBmVn+
AQgTjKD50AcJ2V9U+axNdmgLrLSevMUPViP/+j+wOytq+fpzvAImJ1DiGOjoczWf
sjXyIkQ7RmOnHqzboIA4jFzsPpk9zJNGk/p6DfpO7AXae/MQ3Paei6q3JpCoyu5x
K2smmlB37WYEIg2Opdw5mgueR3DTV6VBzk+xQ2ocOetn5K47qwTf+iIJc+hycafE
OzRanbBKUXBqphan2V/2RvgCKIZwPpTadxlRwycu9yhyNwPg780B+1pSQrJki1kt
W5U58YEPVpg0/YzGzHe7EDiBZSfk1sm/i6oGaiKkEhytZ/WjSm3Jt4wRrtR2cTDK
Na4S+D4BB02XzC/T4JmjVQZAfGpMlQZLpF8h5m1ttTKzi+bi9vU7nWVIgDhMZDo7
WB1Z9TESa/Y6rZsRT35ORK9w2LYww7CArM6lHeFHps9ihTpnH7T5V5YHYxJTkOFS
DMYLMXSZgOFHhWptBBxW1WZBEtuGuwSUDlBgbatDe0cUqGE/UvuIUe0F/9YcwgtA
URcpF02A0gONhTWs40h6lFgrW9a4mP97inV9cz0PRV+UySRaZ1rRNjbObwbCCGtC
ldZTyDFT7ansmsRLd2VicQjrd66yUDfBMI6CPCfAPXXiG8/MahPeZ73yhLdx8M2I
vccTOc/WeU+p35p3H7a7l527a/cQyu34yBaA5RwpaQAooGI2Lpel8PQB8cf3flTe
eEMfdGf1y5NyBX+fFsifTQej6bprGGOXZ2i33KQLze5g7xYujf84e91mbNQb5glR
eHz6b7WVO618mQuVH+zmmRU88CpMMOP2IyVhsFviPxhcU4pI8p6VR5sGGdY+voW8
mSJIIsLwRoZdjuItEBNFnTEK65zgOu16yAK3vz9sS2HlWS5HxXzAYlMnYEtraITB
KlG43LeCaBEshpo+dFj0MUZCZhYGJO3moUZ8+Er7XOjN2nJBYl0N+/oGEhi50xKF
KEJYIFawOVwQ85iUJUosvWbZN4hdGhZCY8sfDeKHcFsiv5K4XKCdjUmbDXDk7sna
+52V6IXBsGrtGoa0BYqFJaSiZvd2bnRWnFMtCOnNZlZzxBzxOaYIfKJTQ/NYldMe
+k8XqYzdvSZPLe3ZmmC3Po1ldjFGIErv6EwK61Dh+moc1KC14E+OV+MI5wdjLrBd
CUahpHcLh2aSX1BIFvJtkfTDM/4y1qhS9V4yXVkc/BOeUuE+nKJ1vvFAnuKRM7YL
GoX2DFo6D2PoKnI+5kE5voN6DKh/OvCHrguyp2a1iNCPeGsWeYiFanyhezIoC3ha
QCrnOOBG7iLfIxT8w2aoPgQQTPza8XEysvpXuDHdCk2eK1g0ZW8L02mTn+TgiWtd
cczwuE5XcrPS1u2IKMkVtlzHB65QIaKi9KePAajF/ypMNj+QAp2vA39o3IvPn3k6
QOj8XAfrAsEtVuPjilWkClp1vznYws09BtUn1cEcwHNfLjueRL5W9Ew0eXf52RKw
T5dZWgTAcjXckTEpnizJPj2fKuMD/DYPqPAfN/AcngO0igshYBdKjqb01nmbapnX
e6M252MRkkPyepWL1SIzDQ==
//pragma protect end_data_block
//pragma protect digest_block
rDQXPCvHnl1kPaI+JU0XmU9Qxmo=
//pragma protect end_digest_block
//pragma protect end_protected

`endif //GUARD_SVT_CHI_SCENARIO_COVERAGE_DATABASE_SV
