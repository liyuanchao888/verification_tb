
`ifndef GUARD_SVT_AXI_COMMON_SV
`define GUARD_SVT_AXI_COMMON_SV

`include "svt_axi_defines.svi"
typedef class svt_axi_checker;
typedef class svt_axi_port_monitor;
`ifndef SVT_EXCLUDE_VCAP
typedef class svt_axi_fifo_rate_control;
`endif

 /** @cond PRIVATE */

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif

class svt_axi_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** Analysis port makes observed tranactions available to the user */
`ifdef SVT_UVM_TECHNOLOGY
  uvm_analysis_port#(svt_axi_transaction) item_started_port;
  uvm_analysis_port#(svt_axi_transaction) item_observed_port;
  uvm_analysis_port#(uvm_tlm_generic_payload) tlm_generic_payload_observed_port;
  uvm_analysis_port#(svt_axi_snoop_transaction) snoop_item_started_port;
  uvm_analysis_port#(svt_axi_snoop_transaction) snoop_item_observed_port;
  svt_event_pool event_pool;
`elsif SVT_OVM_TECHNOLOGY
  ovm_analysis_port#(svt_axi_transaction) item_started_port;
  ovm_analysis_port#(svt_axi_transaction) item_observed_port;
  ovm_analysis_port#(svt_axi_snoop_transaction) snoop_item_started_port;
  ovm_analysis_port#(svt_axi_snoop_transaction) snoop_item_observed_port;
  svt_event_pool event_pool;
`else
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_transaction) item_started_port;
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_transaction) item_observed_port;
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_snoop_transaction) snoop_item_started_port;
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_snoop_transaction) snoop_item_observed_port;
`endif

  /** Report/log object */
`ifdef SVT_UVM_TECHNOLOGY
  protected uvm_report_object reporter; 
`elsif SVT_OVM_TECHNOLOGY
  protected ovm_report_object reporter; 
`else
  protected vmm_log log;
`endif

 /** Handle to the checker class */
 svt_axi_checker axi_checker;

 /** Handle to the port monitor */
 svt_axi_port_monitor port_monitor;

`ifndef SVT_EXCLUDE_VCAP
 /** Handle to the FIFO rate control class for WRITE xacts */
 svt_axi_fifo_rate_control write_xact_fifo_rate_control;

 /** Handle to the FIFO rate control class for READ xacts*/
 svt_axi_fifo_rate_control read_xact_fifo_rate_control; 

 /** FIFO rate control configuration for READ xacts*/
 svt_fifo_rate_control_configuration read_xact_fifo_rate_control_config; 

 /** FIFO rate control configuration for WRITE xacts*/
 svt_fifo_rate_control_configuration write_xact_fifo_rate_control_config; 
 `endif

 /** Sticky flag that indicates whether the monitor has entred run phase */
 bit is_running = 0;

 /** Sticky flag that gets set when a reset is asserted */
 bit reset_flag = 0;

 /** Flags that is set when a 0->1 transition of reset is observed */
 bit reset_transition_observed = 0;

 /** Indicates if reset is in progress */
 bit is_reset = 1;

 /** Indicates if synchronized reset is in progress */
 bit is_reset_sync = 1;

 /** Sampled value of reset */
 logic observed_reset = 0;
 
 /** Variable that stores the exclusive write transaction count */
 int excl_access_cnt = 0;

 /** expected exclusive read response */
 svt_axi_transaction::resp_type_enum expected_excl_rresp[*];

 /** expected exclusive write response */
 svt_axi_transaction::resp_type_enum expected_excl_bresp[*];

 /** flag for received exclusive read transaction error */
 protected bit excl_read_error;

 /** flag for received exclusive read transaction error */
 protected bit excl_write_error;

`ifndef SVT_EXCLUDE_VCAP
  /** The current fill level of the READ FIFO */
  protected int global_read_fifo_curr_fill_level = 0;

  /** The current fill level of the WRITE FIFO */
  protected int global_write_fifo_curr_fill_level = 0;

  /** The total number of bytes of all active write transactions in the queue */
  protected int global_total_expected_write_fill_level = 0;

  /** The total number of bytes of all active read transactions in the queue */
  protected int global_total_expected_read_fill_level = 0;
`endif


 /** Internal queue to buffer the incomming exclusive read transactions */
 svt_axi_transaction exclusive_read_queue[$];

 /** Internal queue to buffer the current exclusive read due to reset of 
   * address by incoming exclusive read transactions */
 svt_axi_transaction exclusive_read_reset_queue[$];

 /** It sets ID to 1 if exclusive access at any monitored read location
   * is failed due to current normal write transaction to same address */
 protected bit excl_fail[bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0]];

 /** * It sets ID to 1 when matching exclusive write transaction has been received */ 
 protected bit matching_excl_wr_id[*];

 /** Semaphore that controls access of exclusive_read_queue during read
  * operation. */
 protected semaphore exclusive_read_sema;

 /** Semaphore that controls access of exclusive_read_queue during write
  * operation. */
 protected semaphore exclusive_write_sema;
  
  
 /** Timer used to track exclusive write transaction followed by exclusive read */
 svt_timer excl_read_write_timer[*];

 /** Semaphore that controls access of perf_rec_queue during read and write
  * operation. */
 protected semaphore perf_rec_queue_sema;


 // ****************************************************************************
 // Protected Data Properties
 // ****************************************************************************
 /** 
   * Triggered when a reset is received 
   * If a reset in received, this event is triggered prior
   * to the is_sampled event to ensure that all threads are terminated 
   */
  protected event reset_received;
  
  /** Triggered when a new transaction is started */
  protected event new_transaction_started;
  
  /** Triggered when a new READ transaction is started */
  protected event new_read_transaction_started;
 
  /** Triggered when a new transaction is started */
  protected event new_write_transaction_started;
  
  /** Triggered when a READ element is deleted from active xact queue */
  protected event active_read_xact_queue_empty;
  /** Triggered when a WRITE element is deleted from active xact queue */
  protected event active_write_xact_queue_empty;

  /** port configuration */
  protected svt_axi_port_configuration cfg;

  /** clock period */ 
  protected real clock_period = -1;

  /** current cycle */
  protected longint curr_cycle = 0;

  /** current time */
  protected real curr_time;

  /** Async reset assertion time*/
   protected real reset_async_time;

  /** Stores the last sample time. Used for calculating clock period */
  protected real last_sample_time = -1;

  /** The cycle in which last arvalid was driven high*/
  protected int last_arvalid_cycle = 0;

  /** The cycle in which last arready was sampled high*/
  protected int last_arready_cycle = 0;

  /** The cycle in which last awvalid was driven high*/
  protected int last_awvalid_cycle = 0;

  /** The cycle in which last awready was sampled high*/
  protected int last_awready_cycle = 0;

  /** The cycle in which last wvalid was driven high*/
  protected int last_wvalid_cycle = 0;

  /** The cycle in which last wready was sampled high*/
  protected int last_wready_cycle = 0;

  /** The cycle in which last wlast, wvalid, wready was sampled high*/
  protected int last_wlast_wvalid_wready_cycle = 0;

  /** The cycle in which last rlast, rvalid, rready was sampled high*/
  protected int last_rlast_rvalid_rready_cycle = 0;

  /** The cycle in which last rvalid was sampled high*/
  protected int last_rvalid_cycle = 0;

  /** The cycle in which last rready was sampled high*/
  protected int last_rready_cycle = 0;

  /** The cycle in which last bvalid was sampled high*/
  protected int last_bvalid_cycle = 0;

  /** The cycle in which last bready was driven high*/
  protected int last_bready_cycle = 0;

  /** The cycle in which last acvalid was sampled high*/
  protected int last_acvalid_cycle = 0;

  /** The cycle in which last acready was driven high*/
  protected int last_acready_cycle = 0;

  /** The cycle in which last crvalid was sampled high*/
  protected int last_crvalid_cycle = 0;

  /** The cycle in which last crready was driven high*/
  protected int last_crready_cycle = 0;

  /** The cycle in which last cdvalid was sampled high*/
  protected int last_cdvalid_cycle = 0;

  /** The cycle in which last cdready was driven high*/
  protected int last_cdready_cycle = 0;

  /** The cycle in which last tvalid was sampled high*/
  protected int last_tvalid_cycle = 0;

  /** The cycle in which last tready was driven high*/
  protected int last_tready_cycle = 0;

  /** The cycle in which last arvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_arvalid_cycle = 0;

  /** The cycle in which last arready was sampled high - update is deferred by a clock*/
  protected int deferred_last_arready_cycle = 0;

  /** The cycle in which last awvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_awvalid_cycle = 0;

  /** The cycle in which last awready was sampled high - update is deferred by a clock*/
  protected int deferred_last_awready_cycle = 0;

  /** The cycle in which last wvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_wvalid_cycle = 0;

  /** The cycle in which last wready was sampled high - update is deferred by a clock*/
  protected int deferred_last_wready_cycle = 0;

  /** The cycle in which last wlast, wvalid, and wready was sampled high - update is deferred by a clock*/
  protected int deferred_last_wlast_wvalid_wready_cycle = 0;

  /** The cycle in which last rlast, rvalid, and rready was sampled high - update is deferred by a clock*/
  protected int deferred_last_rlast_rvalid_rready_cycle = 0;

  /** The cycle in which last rvalid was sampled high - update is deferred by a clock*/ 
  protected int deferred_last_rvalid_cycle = 0;

  /** The cycle in which last rready was sampled high - update is deferred by a clock*/
  protected int deferred_last_rready_cycle = 0;

  /** The cycle in which last bvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_bvalid_cycle = 0;

  /** The cycle in which last bready was driven high - update is deferred by a clock*/
  protected int deferred_last_bready_cycle = 0;

  /** The cycle in which last acvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_acvalid_cycle = 0;

  /** The cycle in which last acready was driven high - update is deferred by a clock*/
  protected int deferred_last_acready_cycle = 0;

  /** The cycle in which last crvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_crvalid_cycle = 0;

  /** The cycle in which last crready was driven high - update is deferred by a clock*/
  protected int deferred_last_crready_cycle = 0;

  /** The cycle in which last cdvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_cdvalid_cycle = 0;

  /** The cycle in which last cdready was driven high - update is deferred by a clock*/
  protected int deferred_last_cdready_cycle = 0;

  /** The cycle in which last tvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_tvalid_cycle = 0;

  /** The cycle in which last tready was sampled high - update is deferred by a clock*/
  protected int deferred_last_tready_cycle = 0;

  /**
    * The configuration that will be used for the current time interval
    */
  svt_axi_port_configuration curr_perf_config;

  /**
    * New configuration submitted by user which may have updated performance
    * constraints and which need to be used at the next time interval
    */
  svt_axi_port_configuration new_perf_config;
  
  /** Timer used for performance intervals */
  svt_timer perf_interval_timer;

  /** Timer to track periods of inactivity for READ on the interface */
  svt_timer perf_read_inactivity_timer;

  /** Timer to track periods of inactivity for WRITE on the interface */
  svt_timer perf_write_inactivity_timer;

  svt_amba_perf_rec_base  perf_rec_queue[$];

  bit stop_perf_timers = 0;

  svt_amba_perf_calc_base perf_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_write_throughput_calc;

  svt_amba_perf_calc_base perf_min_write_throughput_calc;

  svt_amba_perf_calc_base perf_max_read_throughput_calc;

  svt_amba_perf_calc_base perf_min_read_throughput_calc;

  svt_amba_perf_calc_base perf_max_write_bandwidth_calc;

  svt_amba_perf_calc_base perf_min_write_bandwidth_calc;

  svt_amba_perf_calc_base perf_max_read_bandwidth_calc;

  svt_amba_perf_calc_base perf_min_read_bandwidth_calc;

  //vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
EtoqtgWPYykRk1pNr2+z1scykJmWYZtbfjolzuuZ64p4icHkHnkFodbvE7D1MJXg
lyH/yn0ZQBJkIFLa5ZYe5Hmay9dbs0nE3p5q17q9zY4s7YDqI09k0+8eTar4k9KU
2RYpzY+ohZ2HP5wiUkPeF93qyX/klbzeobR6F5yVLfg6ZYv6YZ3Ezg==
//pragma protect end_key_block
//pragma protect digest_block
vT5AU9UMz3m4QPFna+Z51SfqbHM=
//pragma protect end_digest_block
//pragma protect data_block
sBZ/+j7B2t5Jh6fA2a9DdBJ0fHsXugWtVEUe7vts7S6JMFLyqOY0rcrNDV7MxxyO
j0/usJu6ezWkQyB3qQ3Z5X7c3n+QBgmUrRXaZGDbrjXsiOkv3gCSC878fmA8Q/qJ
NsCOYt2z3q/OrlRZ8ozjov28TVWBevDJDt8zophPjYkhli35zsARZe1BLp2QR9gY
5bOjC2Of9Hc5JwuCSPtFlvxr2rG33QQJMK8TG62H9ucVqNMD16Axa5wZAyamRNtt
M9c8rP2tKNSX7GC/QPPzW1yLP3ie9+MmkQHICATuTFDR3AwfY1uWtfUbUXRD/rH3
ucZPlT16kTUKDA+UXc/0j+KYK/Kq4R0lFyBe1TsTMy/eGWQnNRHDMN1LNPH3UA0D
fiAC9dqLCnidcJp7SRtKrqYt9tWcFap+rwzs61OAoB9yJapdudTkgm/qVdLtNFPS
w0cev0gQ7Iz7pKd6XQm2u5dWXvt3OhhykOd39308InfUaz9htXurMD2FoiEl9FTb
YSoDaxw7sflRPxzZclEDodUHWWhgB5kMWoo/roO50H+GBwS2c3UBT7YsXugzzj6M
ieDcV9qM/GvSSrim9DjbuxzLMG8Rjd82S3q6kWhR42I/XU9USwL434wpL/WazRxL
rkbOD+5DkDhDlmejxJHRkVJgF6qixmT4bUgHqvSKSU4=
//pragma protect end_data_block
//pragma protect digest_block
VL+F4i/R0DAoq9OH9rX2BykkPXo=
//pragma protect end_digest_block
//pragma protect end_protected

 /** @cond PRIVATE */
 // ****************************************************************************
 // Local Data Properties
 // ****************************************************************************
 int report_new_clock_period = -1;
 /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /** Variable that keeps count of number of DVM Syncs which are accepted and DVMCOMPLETEs
    * are yet to be added to the queue */
  int num_active_dvm_sync_xacts = 0;

    /**
    * Method that auto generates DVM complete transactions
    *
    * @ param snoop_xact Handle to the DVM SYNC transaction for which DVM complete must be generated
    * @ param phase UVM phase from which this task is called
    */
`ifdef SVT_VMM_TECHNOLOGY
  extern virtual task send_auto_gen_dvm_complete(svt_axi_master_snoop_transaction snoop_xact);
`else
  extern virtual task send_auto_gen_dvm_complete(svt_axi_master_snoop_transaction snoop_xact, svt_phase phase);
`endif

  /** Returns if all Snoop DVM COMPLETEs are received for coherent DVM Sync sent */
  extern virtual function bit is_dvm_snoop_sync_complete_done();

  /** Wait for conditions for DVM */
  extern virtual task check_and_wait_for_dvm_complete_conditions(svt_axi_transaction xact);



  /** @endcond */

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter UVM report object used for messaging
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter OVM report object used for messaging
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_xactor xactor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Detects reset async */
   extern virtual task sample_reset_async();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Initializes master I/F output signals to 0 at 0 simulation time */
  extern virtual task async_init_signals();
  
  extern virtual task suspend_signal(string signal_name = "");
  
  extern virtual task resume_signal(string signal_name = "");

  /** Initializes master I/F output signals to 0 at 0 simulation time */
  extern virtual task default_signal_values_async_reset();
  
  /** Initializes master I/F output signals to 0 after waiting for a clock cycle delay */
  extern virtual task initialize_during_dynamic_reset();

  /** Initializes signals */
  extern virtual task initialize_signals();

  /**Aborts the transactions and writes to analysis port if reset is in progress. */
  extern virtual task process_reset_for_new_transaction(svt_axi_transaction xact);

  /** Sets the configuration */
  extern virtual function void set_cfg(svt_axi_port_configuration cfg);

  /** Waits for a any transaction to end. */
  extern virtual task wait_for_any_transaction_ended();

   /** Sets the clock period */
  extern function void set_clock_period();

   /** Returns clock period value*/
  extern virtual function real get_clock_period();

   /** Returns current clock cycle value*/
  extern virtual function longint get_current_clock_cycle();

   /** Returns current time measured as (current clock cycle * clock period) */
  extern virtual function real get_current_time();

  /** Creates timers used in the model */
  extern virtual function void create_timers();

  /**
   * Sets the delays in the transaction based on observed values.
   * Calls to this function must be made before "set_deferred_event_cycles" 
   * (which updates the "deferred_last_*" variables) is called to reflect the
   * corresponding values in "last_*" in variables of this cycle. 
   * In the case of bvalid_delay, bvalid can be sent before the address
   * is received or after the address is received. In either case, the 
   * burst_length information is required to calculate the bvalid_delay.
   * If bvalid is sent before the address, the call to this function to
   * update bvalid_delay must happen only when the address is received 
   * If bvalid is sent after the address, the call can be
   * made when bvalid is sampled (as in the case of other signals)
   */
  extern function void set_observed_transaction_delay(svt_axi_transaction xact, string delay_type);

  /**
    * Sets the "deferred_" variables to the values passed through this function.
    * The set_observed_transaction_delay function works based on the "deferred_"
    * values of event cycles. This function needs to be called after the 
    * set_observed_transaction_delay function is called, so that the current
    * cycle information is propogated to the corresponding "deferred_*" variables.
    */ 
  extern function void set_deferred_event_cycles();

  /** Checks if the handle given matches any of those of the active transactions. */
  extern virtual function void check_xact_handle(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

   /** Checks coherent transaction. If data is available in cache it is retreived */ 
  extern virtual task process_coherent_transaction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Reserves an index in cache for allocation of this transaction */ 
  extern virtual task reserve_cache_allocation(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output `SVT_AXI_MASTER_TRANSACTION_TYPE lru_xact);

  /** Does the necessary processing to end a transaction */
  extern virtual task end_transaction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit is_removed=0);

  /** 
    * Updates the cache based on snoop response assigned by user after 
    * receiving a snoop transaction from the input channel 
    */
  extern virtual task post_snoop_cache_update(svt_axi_master_snoop_transaction snoop_xact);

  /** Waits for post_snoop_cache_update() method to complete if any activity
    * is observed on the SNOOP channel */
  extern virtual task is_post_snoop_cache_update_done(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit check_outstanding_queue= 0);

  /** Adds a new snoop transaction to the queue */
  extern virtual task add_to_master_snoop_active(svt_axi_master_snoop_transaction xact);

  /** Adds a new snoop transaction to the queue */
  extern virtual task add_to_ic_snoop_active(svt_axi_ic_snoop_transaction xact);

  /** Drives the awakeup signal during idle time period of addr channel */
  extern virtual task toggle_awakeup_signals_during_idle_channel( );
  
  /** Drives the acwakeup signal during idle time period of addr channel */
  extern virtual task toggle_acwakeup_signals_during_idle_snoop_channel( );
  /** 
    * Adds the transaction to the internal queue. 
    * Blocks when the  number of outstanding transactions is
    * the configured max. value.
    */
  extern virtual task add_to_master_active(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Notifies the slave that a new transaction is received from input port.
    */
  extern virtual task notify_slave_new_xact_received_from_input_port(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** 
    * Waits for a new snoop transaction. The monitor uses this task to get a 
    * handle to the new snoop transaction.
    */ 
  extern virtual task wait_for_acvalid(output svt_axi_master_snoop_transaction xact);

  /*
   * Returns the number of outstanding transactions
   */
  extern virtual function int get_number_of_outstanding_master_transactions(bit silent = 1, output `SVT_AXI_MASTER_TRANSACTION_TYPE actvQ[$]);

  /** Returns the number of outstanding transactions. */
  extern virtual function int get_number_of_outstanding_slave_transactions(bit silent = 1, output `SVT_AXI_SLAVE_TRANSACTION_TYPE actvQ[$]);

  /** Returns the number of auto-generated transactions. */
  extern virtual function int get_number_auto_generated_xacts();

  /** Returns the number of dropped coherent transactions. */
  extern virtual function int get_number_dropped_coherent_xacts();

  /** Advances clock by #num_clocks */
  extern virtual task advance_clock(int num_clocks);

  /** Steps one clock*/
  extern virtual task step_monitor_clock();

  /** Waits until a valid or handshake takes place on any channel*/
  extern virtual task wait_for_bus_activity();

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_arvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_awvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_first_data_before_addr_wvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_tvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Drive the idle values after initial reset */
  extern virtual task drive_idle_val_initial_reset();

  /** 
    * Adds the transaction to the active queue. 
    * Blocks when the  number of outstanding transactions is
    * the configured max. value.
    */
  extern virtual task load_active_from_master_buffer ();

  /** 
    * Adds the transaction to read_xact_buffer or write_xact_buffer 
    * depending on whether its a read or write transaction. 
    */
  extern virtual task add_to_master_buffer(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);
  /** Detects initial reset */
  extern virtual function void detect_initial_reset();

  // -----------------------------------------------------------------------------
  //                                EXCLUSIVE PROCESSING BEGIN
  // -----------------------------------------------------------------------------
  /** It returns 1 if there are pending exclusive read transactions in
   * exclusive_read_queue for which matching exclusive write has not come
   * */
  extern virtual function bit pending_exclusive_access_transactions();

  /** It checks the transaction with the same ID stored in the queue */
  extern virtual function void check_exclusive_sameid(svt_axi_transaction xact);

    /** Pushes the transaction into exclusive read queue after all the data beats
    * of exclusive read transaction is received
    */
  extern virtual function void push_exclusive_read_transactions(svt_axi_transaction xact, string kind="");
 
 /**  Removes  the transaction from exclusive read queue if any of the data beats recieves a erroneous response
    * of exclusive read transaction is received
    */
  extern virtual function void remove_exclusive_read_transactions(svt_axi_transaction xact);

  /** function that compares the expected and configured RRESP for exclusive
   * read transactions */
  extern virtual function void perform_exclusive_read_resp_checks(svt_axi_transaction excl_resp_xact);

  /** It returns 1 if transaction with AWID = ARID exist in the exclusive_read_queue queue */
  extern virtual function bit get_exclusive_read_index(input logic [`SVT_AXI_MAX_ID_WIDTH - 1 : 0] awid, 
                                                       logic [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,
                                                       output int ex_rd_idx);
  

  /** It monitors memory location for exclusive access */
  extern virtual function void check_exclusive_memory(svt_axi_transaction current_xact);
  
  /** It monitors the response for exclusive write transaction */
  //extern virtual function void process_exclusive_write_response(svt_axi_transaction excl_resp_xact, input bit excl_write_error);
  extern virtual function void process_exclusive_write_response(svt_axi_transaction excl_resp_xact, input bit excl_write_error, string kind="");
  // -----------------------------------------------------------------------------


  extern virtual task wait_for_cache_update_post_curr_snoop(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit is_snoop_to_same_cache_line);

  extern virtual task add_to_master_current_queue(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual function bit add_xact_with_same_id_to_queue(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,output bit[`SVT_AXI_MAX_ID_WIDTH-1:0]  unused_ids_by_active_master_transaction);

  extern virtual task update_current_snoop_xact_handle(svt_axi_master_snoop_transaction snoop_xact);

  /**
    * Creates the transaction inactivity timer
    */
  extern virtual function svt_timer create_xact_inactivity_timer();


  /** Tracks transaction inactivity */
  extern virtual task track_transaction_inactivity_timeout(svt_axi_transaction xact);

  /** Waits until the transaction ends */
  extern virtual task wait_for_transaction_ended(svt_axi_transaction xact);

  /**
    * Tracks suspended snoop xacts and triggers events when they are ready
    * to be added to the queue
    */
  extern virtual task track_suspended_snoop_xacts();

  /** Updates response parameters when supplied through delayed response port */
  extern virtual task update_delayed_response_parameters(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** returns a single unique number from xact ID and ADDRESS */
  extern function bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0] get_uniq_num_from_id_addr(svt_axi_transaction xact);

  /* returns address part of the unique address-id combinatorial number */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH -1 : 0] get_addr_from_num(bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0] num);

  /* returns id part of the unique address-id combinatorial number */
  extern function bit[`SVT_AXI_MAX_ID_WIDTH-1 : 0] get_id_from_num(bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0] num);

  //-------------------------------------------------------------------
  //                       PERFORMANCE ANALYSIS
  //------------------------------------------------------------------
  /** Main task that tracks performance parameters */
  extern task track_performance_parameters();

  /** updates the READ inactivity time performance parameters */
  extern task track_inactivity_time_for_reads(int perf_rec_index);

  /** updates the WRITE inactivity time performance parameters */
  extern task  track_inactivity_time_for_writes(int perf_rec_index);
  
  /** Updates performance parameters when a transaction ends */
  extern function void update_xact_performance_parameters(svt_axi_transaction xact);

  /** Updates performance configuration parameters based on a new configuration*/
  extern function void update_performance_config_parameters();

  /** Collects performance statistics when an interval ends */
  extern function void collect_perf_stats();

  /** Creates all the performance classes used for calculation of each metric */
  extern function void create_perf_calc_base(svt_axi_port_configuration cfg);

  /** Gets the performance report as a string */
  extern function string get_performance_report();

  /**
   * When invoked, indicates if the performance monitoring is in progress or not.
   * - This is applicable only when the svt_axi_port_configuration::perf_recording_interval is set to -1.
   * - Returns 1 if performance monitoring is in progress when this method is invoked
   * - Returns 0 if performance monitoring is not in progress when this method is invoked
   * .
   */
  extern function bit is_performance_monitoring_in_progress();

  /** Reports end-of-simulation summary report, checks etc */
  extern virtual function void report();

  /** format report string */
  extern function string format_report_str(string exp_str, real exp_val, string act_str, real act_val, string unit_str);

  /** Gets summary report based on values in perf_rec */
  extern function string get_summary_report(svt_amba_perf_rec_base perf_rec);

  /** Stops all performance monitoring and kills the thread that is tracking performance */
  extern function void stop_performance_monitoring();

  /**
   * When invoked, performance monitoring will be stopped if already the monitoring is in progress.
   * - This is applicable only when the svt_axi_port_configuration::perf_recording_interval is set to -1.
   * - Returns 1 if performance monitoring is stopped as a result of this method invocation
   * - Returns 0 if performance monitoring is not stopped as a result of this method invocation
   * - If the performance monitoring is in progress, that is is_performance_monitoring_in_progress() returns 1,
   *   but the axi_port_perf_stop_performance_monitoring() is not invoked, the port monitor invokes stop_performance_monitoring
   *   method during extract phase.
   * .
   */
  extern function bit axi_port_perf_stop_performance_monitoring();

`ifdef SVT_AMBA_ENABLE_C_BASED_MEM
  /** Converts an AXI transaction to memory transaction */
  extern function bit convert_axi_to_mem_transaction(svt_axi_transaction xact, int mem_data_width, bit convert_read_data, output svt_mem_transaction mem_xact[$]);

  /** Populates data in memory transaction into the given AXI transaction */
  extern function bit populate_mem_data_to_axi_xact(svt_mem_transaction mem_xact[$], int mem_data_width, svt_axi_transaction xact);
`endif  

  /** Enables/disables performance monitoring of each metric based on configuration*/
  extern function void check_performance_monitors(svt_axi_port_configuration cfg);

  /** Enables/disables of all performance monitors based on the argument */
  extern function void set_performance_monitoring(bit enable_monitoring = 1);

`ifdef SVT_UVM_TECHNOLOGY
  extern task write_to_tlm_generic_payload_analysis_port(svt_axi_transaction xact);
`endif

  `ifdef SVT_AXI_QVN_ENABLE
  extern virtual task qvn_process_token_request();
  `endif

  /** Tracks the timeout for the signal argument provided with its timeout value given
    * w.r.t to the event or status provided in the argument list. 
    * Mode will be changed to enum type as seperate activity. 
    */
  extern task track_timeout(svt_axi_transaction xact, 
                            longint timeout_val,
                            string timer_name, 
                            int mode, 
                            bit status_equal,
                            svt_axi_transaction::status_enum sts_val,
                            event timeout_event,
                            string port_mon_name=""
                           );

  /** Tracks the snoop channel timeout for the signal argument provided with its timeout value given
    * w.r.t to the event or status provided in the argument list 
    * Mode will be changed to enum type as seperate activity. 
    */
  extern task track_snoop_timeout(svt_axi_snoop_transaction xact, 
                            longint timeout_val,
                            string timer_name, 
                            int mode, 
                            bit status_equal,
                            svt_axi_transaction::status_enum sts_val,
                            event timeout_event,
                            string port_mon_name=""
                           );			   

  /** pushes an exernal coherent transaction into port monitor */
  extern virtual task push_external_coherent_xact(svt_axi_transaction xact);
  /** pushes an exernal snoop transaction into port monitor */
  extern virtual task push_external_snoop_xact(svt_axi_snoop_transaction xact);

  /** 
  * Returns the number of READ transcations that have started  and in 
  * active queue
  */
  extern virtual function int get_num_started_read_xacts();
  /** 
  * Returns the number of WRITE transcations that have started  and in 
  * active queue
  */
  extern virtual function int get_num_started_write_xacts();

  /**
    * This method is used to get list of all IDs which are currently under use by outstanding transactions. However, user
    * can choose the type of outstanding transactions this method should consider while extracting ID of active transactions.
    * "mode" and "rw_type" arguments should be used for this purpose.
    *
    * It returns '1' if total number of unique IDs currently used by active transactions, is less than all possible ID that can
    * be used by an AXI transaction. This helps in determining whether randomizing ID field of a new transaction which should
    * not be part of the all the IDs currently in use, is possible or not.
    * 
    * @param mode Type of outstanding transactions this method should consider while extracting ID of active transactions.
    *             Currently it supports following modes (defined as string) ::
    *               - "non_dvm_non_barrier" => all transactions which are neither DVM nor Barrier  (default)
    *               - "non_dvm"             => all transactions which are not DVM 
    *               - "non_barrier"         => all transactions which are not Barrier 
    *               - "dvm"                 => all transactions which are of DVM type 
    *               - "barrier"             => all transactions which are of Barrier type
    *               - "dvm_barrier"         => all transactions which are either DVM or Barrier type
    *               - Note: if "rw_type" is set to '0' then only read channel transactions will be considered for non-dvm
    *                       and non-barrier type
    *               .
    * 
    * @param rw_type Indicates which channel id width should be considered.
    *               - ' 0 ' => only read channel id width and transactions should be used
    *               - ' 1 ' => only write channel id width and transactions should be used
    *               - '-1 ' => common or either of read or write channel id width and transactions are used
    *               .
    * 
    * @param use_min_width If set to '1', minimum of read and write channel id width should be used otherwise maximum.
    *               This is applicable only if "rw_type == -1" i.e. no particular channel id width is specified.
    * 
    * @param silent Suppresses debug messages from this method if set to '1'
    */
  extern virtual function bit get_ids_used_by_active_master_transactions(output bit[`SVT_AXI_MAX_ID_WIDTH-1:0] id_list[$], input string mode="non_dvm_non_barrier", input int rw_type=-1, input bit use_min_width=1, input bit silent=1);

 /**
   * Method that randomizes DVM complete transaction
   *
   * @return A handle to the randomized DVM complete transaction 
   */
  extern virtual function `SVT_AXI_MASTER_TRANSACTION_TYPE randomize_dvm_complete_xact();
  extern virtual function bit is_in_reset();
  extern virtual task         wait_for_sampled();

  /** Checks if a WU/WLU transaction is received from the sequencer while
    * there is activity on the snoop channel. This is checked only when
    * snoop_response_data_transfer_mode is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC
    * Needs to be done so that the WL/WLU does not get ahead of an
    * auto-generated WRITEBACK/WRITECLEAN
    */
  extern virtual function bit is_wu_wlu_during_snoop_addr_activity(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /**
    * Waits for WRITEBACK/WRITECLEAN generated for snoops to be added
    * to queue. Applicable only when snoop_response_data_transfer_mode
    * is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC
    */
  extern virtual task wait_for_pending_wb_wc_for_snoop();

  /** Gets the time at which an address was invalidated due to a MAKEINVALID coherent transaction */
  extern virtual function real get_makeinvalid_invalidate_time(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
  /** waits for transaction which has been blocked by other transactions more than `SVT_AXI_NUM_BLOCKED_XACTS_ALLOWED number of times.
    * It wait for those blocked transaction to finish. This will avoid starvation of some type of transactions and will provide
    * more fair chance to all the transactions to proceed
    */
  extern virtual task wait_for_severly_blocked_transactions_to_make_progress(`SVT_AXI_MASTER_TRANSACTION_TYPE xact=null);

  /** waits until VIP is out of reset */
  extern virtual task wait_for_out_of_reset(int mode = 0);

  /** waits until VIP is in reset */
  extern virtual task wait_for_reset(int mode = 0);

  /** Wait for start event for performance monitoring */
  extern task wait_for_performance_monitoring_start_event();

  /** Wait for stop event for performance monitoring */
  extern task wait_for_performance_monitoring_stop_event();

 /** Perform master signal valid checks during reset*/
  extern virtual function void perform_master_signal_valid_checks_during_reset (
                                                                          logic  observed_awvalid,
                                                                          logic  observed_arvalid,
                                                                          logic  observed_wvalid);

/** Perform slave signal valid checks during reset*/
  extern virtual function void perform_slave_signal_valid_checks_during_reset (
                                                                          logic  observed_rvalid,
                                                                          logic  observed_bvalid);

endclass
  /** @endcond */

//----------------------------------------------------------------------------

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
PQQDvrG6hPYpuPnr5Mu9wW1WSsU6g5an9x+gIScnVas3PM33LZrebiA5wPkzKGOL
33EAXPyajrXaQKFAwUONbqU/Z3EZlVtB/z+yFj+WqLlmhB4Vv+Qt5zke3iaarjYw
24V0FOodYx/GBvMt85A2fMalUAPMjnGMPTw4ruWhYAESpeamwCYAVg==
//pragma protect end_key_block
//pragma protect digest_block
AUf3gN/uHCfqeAFdAl3FKaTRtrM=
//pragma protect end_digest_block
//pragma protect data_block
SosJ7JSYoLHwqMOrleaRPDpRT9fKavgVEuVECeznZ++42EcveZTKtvYi3EcIey+0
GEUUx/tPgigu4P98pU6qV+lA4cedeQxMoJFMsEqsWYuYm8eSC1GRwFzGGwll1k8Q
C4CfSm1/4PpZbTi5nCbJTt2yQpmlD7gpXphYM31kOiMbxM42Zg2fiM4EWGmWUYLM
Qw1RZW2K+afx8plA6zoX5v9iGrWq83SAA1SS2OH64oONe9OwjQ6tNdcYlMYifpX+
rijKWipXIRIywIHzPecO9K7YhwS/ObwhtubQPyqzG47UONqNNR4aLmCUNQV9AyqI
rt2c3YdrkUer/gH6d0n9ywS8h4wU8h0Ev2/HwoY6gasTKsp1Yf/e9AvXGjEbxSDP
WKJWtpp3JS1KLe/6G6p4hJJH73RiszXxN60FpoClHl6nqiJuUmab9Jy8+KL+NM7l
vZQzygpHLH/3eL6+5rVXJs/m/fcBAE2Vb2JlszEDrdKRzQ5SicxTLeHpGgiXuOVz
wHXFms6lfoD/BJJ2jUPpg/jm3lQjylwzQf67+/bc84wLXYtH0VNIETnchX7CU9gl
nZMJf+S/Rn24Gjs6IpXJRk4Lu5BR9+bNWnqkwmNN6ZGXWgo/A3RCqZRRRTpZ7rjS
uVO878BQ0XLsekWQRVi9Q4dwRWXcyD2PAQlHyVlD2HqtWbURlc3lTsyevg1i/RxI
K9Wq+ARUYZopFS3lFymY3LJoylsDY8gQ669DMZdJH+dgSG44ywnZCkziIacfx/Uz
F4qGDd0Bk1oKfbCF0rKctdfmhZB1ACuzfMMS+VtarY8V4SNHZvXzVkARXAapDmY2
cbg/LPOmgd9sW29OI/eG1Kg8RlgUG1NAuGkdFN4lcoLnp8hx7VNttrdIRvBjrqkz
pxmR+cu6kEACIrhHwKt5gI9xe308WC4bpyaEW7CbEa5SahUxdkrwHk3W1rcnX9KC
26ohMVea9dAFP7ePkx9zZn/QRwgl57dNGJz378H9WAtOnCxSIIt+PfdMA4jRDweW
OtGbliJZLhGHUpNsSc7NwXRNexVJjnQeQOqVBbpfe9RdqLlY7pdWWQMs1VrIzCiR
XAWZxpQmwlaqdSKZAm9ut3d3joQN/TqwuWXTYCChWfPRtqW+CLChh2YGY5c7Vb34
ort2WlkLSbJfUfcEEZ50SnlGzEkFuwWwVPUh8VKmov2TgAeFcCmHDGd+CymNdQ5i
eYCZmpgSOxgW31RWu0xoZN1VKwW8EBvvIWP6YzJV2iI4xpO2QXbY/e7zxNpiDix+
+rheNETM2Pn67qzPcjbE/ZSFS6NAcs0DrbS90D0FBCHxwuX6gDsrel92SXt7ytrS
bd+K/T6kLLvc6t2wLWMIZTqxfFWvVlGtAJRWyJP700eSQ74ynXy6jD2rXsgi6KWm
M02CqW1d5jqdeBTDeD16kLEevNGJKtm5jE7NBqX8IgGbRJwLYRN5kdsjLzoXV5Bu
W4F46okSgr9uKpXiHuCOU4pSrhTwMKdxdroZNBlz7h1HHdX+M+LkfkQXDutUBOj0
I/BWNjXndZxgIp/PQezCelRS+P7TyJi+9RUnatwHYVMAWxVdsj/GzNIOr33XjSzr
DV7ZqoiMKpD/aTVFuv7KugbQmJiVxHPKmgd5UxQchCkBngA/WLU7x2ILCQFB4/qx
GIDfmGVbnz/1M0h7J8W8axQT8n5vkchMQ5asc6xxWoiiUFTdeE9iuakGM+RzNfO1
2JKorhM4KEwjfeLuMM4hwFoJJz4AI0Fu91PgzWb39PWK9N0aGXWCsGTwLoOf4xUv
TVhKbjuEdPf/BZ7omXfGgHyHkNFgP3pVMFLbr7KwfgibAhURI8r2cDMVPmLrsvjy
GnW+SRkZlvg432otNdBdQooC1idJSshGqFSkZ+6hn3Dx5NBtYBMzgk9YwTrwkOnS
Ma5gDHF76DWO1hCgWWP8MsgCEKwX3kLmCMhqmIVSw7KKdkmXW5zFWSLJ/p/c+wyj
qbci9qdL+IsXzRC9153UcToZ7n4id8q743OCf0q4Ci1Y/QlL1XsRAEKkNk3uDagd
FBCItmCiCE7SNHzMg3QzBO+b7oqg+n7ucfoDBxxAfnpurMCxGSPFzNvxnXCiFRPl
pXJtN3g8MNjVVwRxYCfjg/D452UJjUUuNYJuRxzaZOFTQdzmkL1L99bj5lcBQYwH
6/aiS9n7+Ns80ZZrwfV0/pqX0Lvji+r7ej6Ft+WCw7d/LurtqGK7vFxWPdaAwXOL
IZFBtZov9EElTPuDILrZoMFW8Crn/n2ng+vnzcqgkezSJozpsczW764IEAjgHkJH
dB9kGexhkUwg2SBzbnqP+RW9b3yXRKydO5FC8LbZYVH6zPLMGWcktiUSXtDzplxb
6I7nT+U6U3YB10NLFcO4YzYglTaRkHIsmR362GUWnc1Vk6OxuJZxI7k4SThFIYTF
dYRNAMBP1Y9kQB9UvAO3+ntfpP+oe3sE0V9SCY2S9+PG+iXyPa7M+/Q1JrMpRTY1
PFoMxw6BDHkFUZkaSrgtiAp+DWH91efgxBP8Wj+0l5FEAFm7KGU0gFHEEq5kILgu
ANt5F8v4VTvVtKA+Z+YCYdlpC+92oCn9Q1CzHKiFC/Oh9D2G0xLBUi6R9XUlqsMC
ay1rrYHoL4xX+gE6pTzEBkeDd0yjvlj2492LXxbGAJQCqgivCDZZnGFs9f7nNLuj
bFU2J8SutrHDH3SwlUmvs5iZu2/OI6bS7ZyhGrC9p3hubQZC/rATHw21jDxedO50
jPzgXrNgk8ibvPJAzG7yGrXgkiuexS2KD3v6h2Z26dDBrBXVjQtPUhww0vqFswPb
m3yNb6a63PzkRALRqBjPH/v9bo+s0iuzSB2pXZLEYaXQVhdd5hXA78gGzdMJUZv4
6Zv+JXItE0LDvyDrU/13vg8RNNGZN/2GpNVw91dJO7HnMBaHoFuV+ZGa6+bVBvbX
QS1CxU2e5NnoWwk5RQ0QzKR5ULpQVSfyC5eTUbebeC7Y58tygztJCgooThzOpozh
rlKzUSRGF9qEcZqHpjQzANiyI5QpLwUqfDT8Qq7I4QIrVjAghYYVIggOscqLSzZo
RW4DMaV1L1eq4msyagvC/uGnNknOgvxN/DzRZsWyulLdvlBmBHmP25BI2Y7tNPGM
/v4sYBFFrUMY9Klg8AknhgU4LWXzCoOERyD3xm9DExk9pIMwnuZ6RU/6e9FWYPlV
mTVSTWSMTrF8V3ucFFJssQe6UB9sBstnbMEdKjKSOPaCTRhpNoVyC2vmMDgCq9kp
Kb/IC3v7W4rJ3irrICyvxYjSxqqnOJnbQBWVjt4zhrMzIKP5QqOrUjvcPRG0Im5+
5leonhz4cVxQw3ALw0yDXXAZHvAB5ndhqZwqKWBwaA1OvaLWGJzebvRAJ+lYD1zS
Y7eEoAHNDeVHXhG0DlNGc/xjT+GS/yjEFH8CRueoIb7CMkjY0AHsRsiKS4JIxcvG
85b5xbT5zbfDR2uqCBLvXcpi5LPouBjXmR24fCOawHv7b21FRzh7VXB+qTfF8PZb
cnqpldnuMD0Ac7QRXV+zUCPjFzuqZYl/lQraRLw1pbimO+prA7ufBtM8Brk0Zujc
TxDucX02bZN9jo/l8jL9r5/4xABkstwe1TOIycqVhnDwzzz6UPVMkRKA3l8sGYS7
rD4HpQa93GMCehOlMRbACGuPM8FLH0bUSxwPW6b2FJ2uR9jx90P/32ni5eAn1Vnt
cgQUmshfbockaXYd9ElJ7FeJ1VkcJFPx97+VmQQDliAJCHu6WhM3zYNPBemP5Zn0
JOQnMKv7r2A4ZLmrm0/1ozcDLpGSoBbYRy9I4Ck/I4AmYuCU8h+XaBSnTMKjzudW
r9nfLYT3PcViaWLj2MCjz2leFO2ctjkuUBzOWUxxj/zq3ayis06JwKHp/ICcvCa4
D4Euvx2sIzeObyMU3K5GVr1JmlOb+r/TdC/4kQu5wbtACoLECCacg9+WEAkiNl0N
y2JwiKYfflBmhZLkoMW2XGdoPJHjXKoELpHP9HiaR1hvFKzoyQRZqM5AEofKpjLx
eZIioVWwkeeKmxUy9v0JoQWR9GIewNPUB5M3gHk0MW32AIGdGC4hIzyfhCJXfdag
kZ0qmGna9hJ8T0Fs3vR7VLXEWb1SjeZ6YmQtyqqNJRxvw3ijRo2KqTO69a5Eyrxj
esqT3T2E1FgNuQr7PzsboPdrfrYcW3boht3w2xsWsSQ24kfnFqWHbN+TmAj45nm+
MNBE7OQE+aTzF6cmYO9Nn6Wbpf+cbCoCc/5N+fQiRk9BWGJ7Wr2/nCqhpKBYNRHf
Qad+miQuYgOU/QJk7x2fzoZXCohxLWjWsSIA/tF3FHg/slY7ND+vAI4g8ZjtaiEu
Dsxj/lLQT13FEpRmyGCOwuO2vO2C4KtWylpr5zGpvd+Dks+kBu34g4ewa8IurUtP
apnI+Bg8Hf+K8OvTnXpeGDeQuUs3PAuHEQwGEa/o2Snenchs7pZuPmUUTH4AP+dA
k0H9y2TzeZdiP/ZErLZ1WuAhgFwxFzzUQIbAa+HXu2KMYyeQaD8KSnE/qLDOueTF
PxuDGLDPrpiB4nQmEuIkFf/e/YfLk/LNJSYBVfl2RUQYp0lnLk9T2gKojxgMdGUp
KUg5LO3Vwbr6NQxaATcnD4SSBmhb0ynYhbztX9FF5BTQ+COJlok2JCn5xveqFAIk
/PL3cwHM1G/sFQxSL2kZ8BOENthdgR1rX2NroyW9TpqwAibKl1kQZfFw+31g736D
IVFvCnEiPoUW+VgoeDridCUGYj3cW7FYxA8qvBs4fr+XzxRblv5yRnbv9EgKA3xb
PqvDh8OaNwsQqRgHzuj7BZq7LZKgwWekvy1TkRSVrwHKADRKvD68qUVDIHA+yiwy
jFGLaWugNjQzBlmcllet5ATbGunttrHW867ptyYSaYgkSYXjx2bBGBFwbJ0GyvdO
FpIwOY98GiVzbEN3fOqWROVGQKeqgu5N2aNQ1u8AMpx9QWxGNEVBUp2cbgpE8fpo
45yK9k4mR4ohoe+iyuRjxIpn/ZuJ/U0WBlhXqg2/YRJO+ZQVBc/Zs4J7hnivGZ0w
Szzy1V/jeSpDFt+qcVEKFMATHVmMkUJTjUZmiaWl/4h2fAF4pONihg6tz/aT4LX3
bYzuPonaST52Ux7oaO4RmdAlxRyXJUZ06BbxRMch7YlM2nl019PbKa7dkKJzTUrW
WENVi48Ip09Y2y/e8OjsBgQqShkFSWbM2hdLIyhi7EXTC1AJWXwvL/0lP3Gu+Erp

//pragma protect end_data_block
//pragma protect digest_block
VTt9kCuwz8OiNdDYU/VUalkqPf0=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
1uQbidMgAxzuty5ttatQuG3V97Rj3PGJrfpVKkN42W4j4ezOFOPS39jbHuruHnkq
JKLPaVfegNmBlx3WOrvBCRHqE5ZsrZf88CV8GxZWv4VKfXRxAwiZnZUIg7hADxwZ
CkJfAQc263fc+Ynzes0L02pcqdK9K7vSrZNpZR+1i3CVtaXhqRHNOw==
//pragma protect end_key_block
//pragma protect digest_block
sctEV6pfNGYFrUHsrW8NN3KGZbQ=
//pragma protect end_digest_block
//pragma protect data_block
IxQlgkv8kH4Dv3ZT+NZk9C16n07wfnfhHRorARs/l+I6q/eHWTcZKlB8G3zSX2ZU
oixiZC6/r0/rswdP8Xi7Gz1AgXSMfU47Nqhkeg8e3CdoHrJKbmK7McbpoqtTH7nL
f9wVj9o3pYwIsKXE11Y8v04zPivzDxYxI6aCXQSa02dcWFcZ2IW57cmPJtAAqex7
/OTXZtjOOFM3XDtE9vrwkpQIxhcERMm9+gZcxGUY4NGYBGe6w1t7rgOVOsMTAmpR
UjuTwGlA/rNoQ6cALuj5ij7PdZDp0Zry8RfrIa4f1xKtjkmcDs+XZXTDwKRtcn7G
VPZU+RHtwv+eXn2+R0msK59sxjfwc5EeyeggrXdIYtOXzyt3gxzivoA1+3xUoz4+
qrDcU3nm802piNfa016gKoATjkrHeJUokhDMEkSnDWwTvdqLqa5UEpUP/s7LiMUF
EK2WR7dkpPqEaQEq6rBhEKfrlP94MBAZivGdQ5nk7ca18bJ1hOv6NYZZqkiWm6Ah
Uh9h25LxciTMPtznsgEG8aC3x1f0eAR6h4WKZnIbeaEAM+q/yngzRqyaHLQNZbab
zgw5urPo4amDaFdntMuq4NmS/0avYRCFZXmPcVzA8qVE+4o34ASepdEtpI6i1IER
8gEZTrT/knfdTQ8prL2hAi8pDVG5dStjzjHKRiw+rCBnorO6e7vKtys6bZv59koe
B4by2tD+z07DhHQeeB8ZaorI4S0hPwOhJFlw1mSZT8ydUx5X9Pc+DSBL3LP9PuOZ
0fKXXskBpllDV5BnYcnTy0TiGVrFDuUBUHsRqDw2jmwmyVS6nHGjtju9JdKLWg1E
/Ekg/4hIqn8As4urz1O3H822WXLc/rXVVdeBXn7O09zYQEggp3ULlwPCKQjG+O26
MkUMS5AxCn59aN5VcM3IqYbGpF2Vf44ujX5pYamVRVfKGOtu0CPbKz91fIotCxPq
HgancGCfFGs6cs8hYLTY7b9a7zvReuCPTdEBS45B6FH14uvbDuIIeMQp7slNhc9K
OcX4nGbhe+G0ZPCgdjlwP4J8T5VsQH06/pveO61m03EM7VzWa8OyS3kDHIHvcVDk
lw9NzPYTH13Bh+whuHbZk5swJnl+vBIUy3g1/ZAwfGbOevlVjkhNaH+fP5KgV+Nh
54woC5ymtEUGhJw8FXAGqLaobO9W/To1Yh2HV0RFVhvhyraZgsV4GbfZt6GzBDBZ
njHvF5NRvSGI1y94erRqN0h5bdf2JryEUnbbWfLhN3XfqXYGE1h14rGVxgJ5aJTJ
2ubCch2p+KeG4JBrtKLbYr+hVouDR8KBONgC7fJwR2R1IPBhHn3r2d0ZJdKp7Mlu
/WWCraQfkA0qeFJMSw3GoA+akeXOELrrc/RB4b2lieMa2Z6RtLJQSHnf1UV1RPav
ZPuZIQaeafr3JB78JNWYGaQ8MDOdJSIHpnNcJPFSO0+3bIVdM+t/Fc3MdpOMvp/+
9PMmbF57kE2kR8t6zy07ykUHhGHoqevO/yf9HBrWEjhNiUjpedHyYnDxdEVxbC20
shnqHeOS/WMn1GqZ3uNGT1Z/EFtQO425oZRcpk4q23SEB6CWocX1UMxA5gekU+Da
gQlNKxwqvGyNboghhchz6Xes51FCnj5k0mj5SSutBvZFDlTLbqrdj9F1YCLCw/fY
V4UU1WomG3/Ulg4RKylsS581SPOnkFoC6Am3jDf9KOQLmSKL6koGnvwZeoizEe/Q
Zcs6pm24XIoaPB5QPQg/qjLJh0gVAvZC99Sfo6ufgvJyMg3eGhrUmrmlnK8m/d6H
rOEapfUmvLNxaGIOsuE3vM2YDLlEig4zFEHzTvH8zlbgwR9GR4fbIb35cHaP3dP/
UPTlmJcOwrB7Pl15SmpzvlmcRGaBEGQdJ1GzyT5AY/BmN1rrHn1YzBokcbdIU3qb
SSMb8yoMQZfHnnoBuqRXhoEQnQjFAc/vbI1qHsJTwJ3wKjO10AZ7MrJeVabXVxs9
t2v/b3eRFhE3sTAwHiR8qaW65pqQ2nfMAzaTUgOPeryDQjhzdb8lhbmoWEXhUIOw
sTg8rCVQaK3b/sBPpnrHpvHYxTJei2GwvjdjdYtBD1nkBq/QdUvbSVaLq1E7iDD1
yo44L3obdHRErcH0oBDQqfXnr5OMBft8HMrSNZZixd7pik4cSbDbNwXHgApqbwCA
yal/6jkaCZBfNq+2jp+wapFDihupFG2Sl71sCOvozfUQiNhgdbqNbORSgrhm+z46
/rAqNSdexk1KyolY7BbBoh5zeg4+AdNW3LoCIvJxVy9pylCSzWzwSe+YoQqXrkXT
fRvioBHxU9XmsDbrkzXfUbTtxNzZRDHQAZ5ZG7GTyFUbbwQ53vslMkP59/xTTRfa
IkOEtAoHV71i33nmZbRNDcLCv7gazT3Xt9DKyNh36llf9YyhUo3dQVDmF53IYHFb
gK7QwEanRUJO4fepxEWi3z0dfh7hkCX26LTXDVTHzpiWsdySIKnEKINKMhWlJVza
K807myAspvhhw3ezNAs2onN4zRULztxoVFSIYnBkq7YWxNMbmooJxcQ/Ola28cqo
NPWopl3WFslt0p7raxXS+pibxvrV+2LsBaJN5O2rYDwd+xsswhtSKkXBOMX/SSFz
xIsBIjb3R5gDEpHUYGOeZHALe95tVxkU04hSaoKscQlEoOm9m9M4qAMASaL+0juw
pwoE/fhBcxrVHH8JlJqJe1sv2zrSliYrVDYaPBf/zMzBmRDoQl/VwQa8f3R0YNgr
dnyZ6qvbHCstnatwj3H+VXU+awXlQhx0chGq0xoZyEJcFYSsdZwAaiUtelzATvLV
YqfcwRoclvdkyWHSb06NjjLBpHVp6NbaJAJc7+Xmkq+3AqOtxNtGZv6/YuIez8M6
j93KImFgY7j21FYneTgJwvi5x0TINLzgRIGMvGiLZU3LH2SUlRuLyYeYkxljUwqR
xb2NEuQOdMh1dBSuU/R+pV1P+G1ip822BIdnM7ejKAkKV651pZeqPV7nmPV22+UL
GO4srLxy86aYG0TtVarF5zg9eBVfCSfX7YPOWPDR3UrVHTqt3C6+C+O/NI0ko4Nv
7cn50tPQ7ih3OmznQdlujHFmpohho1WaX5aQW9Z8SBoA2e3b2hRwaHCOuFhQTuFV
MIIq3pQVsd0QrQPuN/yYBY44dip8OgKSw1ibXvqrSFY+n+inKtl/JvXPJ0USyY+K
DWoAbHlrEMKyOiBueHidQWRkBmQ4poQ+8mqGCqGnWXKNEPwRxzabC7ICmyClVmbA
wGAyHpKwtM6wZi+emdGVRjr+fc1pXYVJVHPlr+e0xdt9tCc7E1d03xLsqklHCTYd
Sp2Zhl83sA6lnG8hzgKQAtxERn9B+3gRvJNqEeraniF7sN9OpJe8O9qqj5l0QAgR
99hVf3msvi9WPhVAa2CqUyZdqLbm798p0qJ/eB0R74eMGJhWVdCrmgNnaFQlsHwy
rpUFNgRNUT08Scyll09hVZuNlDq+DL2i/RUPxd4DY3SxCAYVGk37Q7Y2fm3PAVwZ
4HSuqFNKvlEhdQdfZ9SvHtUzHeUH/y1+mV+4Daabl1/CMNVLX3D6NnDKKTtv7Znn
1lPWhPUFxaxN7qf6MGolLuH6rnnmlsSnppUxld+35A5JO8flx32FTc53LxKQCtVr
0Q7iU1oZ4gPf0t8h3UKc0pFA/wE+gCmnz8aL2pXBsB4QWyyWiSz8RtPh+9yGaY/K
8aI7XijPa5fz1F9ejNG5OUP3RXIp2Z6oaYLDJIb+z1l65jAC8OqDs4xrv8lIKneX
SHWcLdfHp/4/it0MPR4aweQuhFCeQYM5g55Hk62O+zGbg6ReyCTJjNTEiuDjdHPT
Bjwz0vD2qv+7incQnBH/BtIVky14W8ZpoNmCNaEON8SAnIqINB5N64qNfwyT1D50
B+anpuAOdS4MtfDnoTwiIyfLccSP6KOJVMN+LG4g0ole4L5jgH6zhKr2OIYVKhmr
Q0QhihIKiGtXSfhRWVQbpK/yMSd5/4bIn+rAbL4y+L5QQ+VzIxg2F1Lw1eMosO1I
NN/hxnd0kS7ccuINzHwFI3TE8MJQcXQZjJ9aFBAzROBR4bs0L/13MAR3kiTOpw5F
vazsYl4a3ouadf7Mjzc6e31yW6kxvaLeIrqQBZ0a6pTFWg4Wq0nHAMWkGatFiCrV
1vp8zi0zNQZbDfwH6AqG1X7tQha4j4StrGhBSll6JArfQJJz1AkHLiK8ugtvf2py
w14fE9y/03EObyc1mr7siCAUPgqIYYgavFuUtlqCk81sZjuaaej0iQ7btSLRyt4E
4eSxtW/ZdPkpqi+FRQf3dbgq7oiCDY1cFBv97gEuzZijdeybKHum/XAMyzE0Toxa
xv/ONIdcJypVZJOwK4tGHqfuR/nhL7HviFp9Ccmw+Qoj7A72STtqaptf6Itk0Dzu
5mGrIEFxIeN55s4I0EQVN9YqskpMeSssXVsG79EW1Hyh3dRTWGjitQqaDIt2U/Qh
RRqyNgRSh7aibuQPTB4jKQEBRPRGPLzpVFraVHpl91w8DgEACTU2GKDW7Pj+IM3b
vVKVhS/AkLV2xIY/qCXmWAttnF2W+VUtHPxVWstZVgohCdGDpAAWdHhVF5JGWhRF
i8kffH+r8gE7535QX+2abkLZtMxRQA9S9E0lTURSuoQ0FVW8VPbdsC4s+qAxBIkX
PoAwNrtuygfMWnI0CSC/nEAL5yP/15m2WoLGAlBbT0h4sNdcwt85fmBEEJQNj2UM
SWgC0924HrrTR1EBhiWz7dqWKBOonl9HWV7nxYM3rypDIVN0X+p5pIy9WtU4t2b6
dG+Atx0ZyycVogZY3QY9Zqct4u/YTc5hl3CMtM6ScOTSwFsc0IRTXMOsnWHUTKLJ
4C/A5+3DF6RaGGum6Uk9G4b9iADziVn1aHOqmhSK1QcGsI6zbUMsyg+m3lKDA/sd
QTngLrHwzUqG8HOrdAQGvmel6s2U9QlqFtdkAHEHnCrQLVr7alwBFsrMXU9EoOoR
GtlJBrYSVA58LWsdawiTDpHqDdGgs09n/iAvZVkMZA822F1jrk+0jttLygsMsG10
I/p0uflFs0iuPYV1c+tr/x3p/cGWT1hEc/mp65JWZ1MdnOI4QTyE1TwiIz+Vnt9v
MUAxlXx5hOcWOg5iq8gtRIbjmmrZcD6AMBm1rUb9pUhoOUXwNlUkt3yIUM9IFVkF
/kppodkqxMRqVjrkm9buAC7g4SX+XFgOUa11VEtK7ajAbKozlrn6GydKu8I4boNz
oCFwbuCUla/LWzSBkFxL1Y1CimGr1xRdePwh5FrASh5nRtCgUAw0+ATCO5PziFti
o0fc7Lrs/9wRKcRdrp4JoKS07iPd7BeNfnR5IXmURm496yMFThoeq4eHmdY/dkZ/
U13MJpGuWXzIpiLVAO6YjpOh7x+9mcH7ie9eTtYJOJKvLex2y4KRaSZYOQRhGC9q
BDfZojUW7cAN9Q/DRGbspFoPlm25U+mYSp6UWwAR3YiyLxfgDqWYyM/2xJqmjmvQ
HQvsYRfVHXQb0GmNpfVmxTo7HJytkLYSCkwRC0ZN0oBlRySC53C/NLaBop6A7KYS
vsjpZZrtrzFJBFzJfMSs8/2DjO8zq/ecvmErF70cf6Njl/PLsLFJ1ctLO1kxFKBT
2ISI/RrP5boVyZhPIwoT9e7hkZA/4hzCmyiRiFZ6vCNiS8vMekDKNOG3jp1eM9SP
w2LyVBBi+m4HIYDX/FEPX7xlkRQ3KB/cZFZX8DALwh3HHLN8rFISr9Y4t7lE/Zey
FZUZMsQh52t65Xmlr9QpWVd3KbI6teNuPFxgkvLX+9zQw+1lL1Gt70jaG1xFQBAb
gKHarVXa9e9f/i31K3uh2Bb/9yHsBwqkh3jbT0yc7bK8T9146auqdWb020OyRXIS
DRODUjmWylHuxLV3gn7njjyqdWfwGHuhaAbG3NWi3BHFENRy53jPBTcm9UR61b3L
KUYX4Jzk5VhG47KJky1dL5jNedhyae7tja4Ml1BuZ1T6oiwcYomqH53z0puDGI/v
jBkVssEE4OosF55FQTtgHh7KhYZAZmpOc5KTFxOBOEiSUHEzM8h3qhKrMutfl6SF
6mbPugKx6wBG6dsZBS+HNXuQCP6WRC8kRws3Zf81q9oJnTzbPjR+3AviYRC0FeEJ
k4dbW7iSpOE9uvLO6GL3JHCA/ANc20gkA8Rmj1ajGBGddQ3VYcVvVHz5u6UkZB7P
NtNRfnJxeFJrrttzMaaKdtdfcdlr4OEj57dJRg1SGPTNTHgLfFoDf/7lYNQrXRni
MuBEvpW+ui2Q2a9vnMAZw4JUTsPfawvPRWqjTXRrkfVE8KwwSrCUee8iRlp1YMJm
KVWBXHMmkrQND7QEZ7eB5Wgi4NcmicBJqqAqwDchc1DfJyBJjs5quyEjFH5ebwVD
X/GZDyGV4aLi6N+wYDBbNauDbDlbSydeB3PenCcK/L1e6vViieNSM6tytay56dPZ
UwrtORKM36O4MM0CD3ED2wCdn+/OEncfLjMBE32xKTE9drqTU/swv5A4Gbfzk6Su
LtzxqqbHY0OGix2GELEqi7etVivqrUx3Ivk/JlNWgvS+N+9sTLZahi6qPHQDo1xA
B6+8PTQeevXGOHUoPBa5wpkRGQmTo3hsP30tf8iZa1PPyCEJg0ngqi0KGP+Hh8fP
GKgh4SlW7xZwUHyttkac7A8Ng8O+2RMedhHMJGKhnVX/yEjZyj/HgNiW1A61P4D3
VKHlCYoGnPVik+TSTjOmCbGtqQDwCPnlrBsbAeOukR4BNyfS5bZKaY8H7obgYqZU
jPgPbufuFkgnobjVtLdUaVVH6rvTzKn9grvuGKF9jKwSgF7P5EaDftRvxUAm8xFd
66k5QWYKcHMdYEPJhOa/pDllB/D9b2qJkxdnFkkLvwef5rXNQKL0s7uM6MMThSMu
gIFX5UWS4uzAWjQQ8AtlUtTKDi6jN4v0iB6fPA7CHj1BMyxy0RuL/Aku02GI+ZdT
wrWcotvPOzSp7wf1oeG8kr/dTM+nFGg/y4kBUh/WYd3uiqdI1kG8tZ9VDKRrZuQR
R0t2aGYIpU2zGXDbFXFRFV6XfULH2IJVxD+NLVDt4HFrEW/Fd7ZoY4DAIVXAr4OT
NiPYiMFMG+3vl3mN1B3BO4w+RmRe8JKxjJoQoMwlxkmb5UcokZ++WjeOqNcNoEAg
SOahBF9b8rlKyevcVIOcqMg6OgOy/qc5B2oOS6RmXecWPHKE3j4EFwKYGgEu3ACN
SCCpvj5sna/1aa8eGo3yyKhvtqhsRkgfip9mq/QTs56Wb9qr0JUsbrQh7/v1ph2E
NzyVF2Dz+P8p9vVx2m/KJVqM8SaSmdflaky7TRnkOWyrR9Q2QN7SxwaXNI0k9bNK
EVRddlkT77esfxvvsJa3sVG+X5aqS2Dans8KB+++aTTo8FLfn/IP9T6NUcumLK85
st9SOXPWd8DJuZ7Dc9q1QCMkLZQmjNgug2YSkA5VW4mUYMnKRf+P55dfeRXvH1/G
SobG+ezhqj8GZhukuSjy4t0wV2Maf1ejSyXNzcTl7MAsq5ULhZdbxyZ/ZLJSpRy4
IAJlnLcBh+h4/EG/MgxcpxAgA7qvB7TC6IvfG1ZQ3/Nl2aeYUIS4EJvojeVLub1j
C+u8TKLdPqdWRpr4mrkjQiZsc/ZSIekXVXpmD9S5hSkeOdEoDEVVXp3Bg0FqEF8s
7kLIkB6nwWy5vJUiG7IGovbsgVdiJTRs8vEpZxndYaoKjL3Cyz36zWdQhY3RrGCh
A3MB5tgypzf59YZKyXuXzO+hsWcVQu5sSOhetX1uHOsuQn3SGtnJJLr8ZDTyVz0D
sgcXt02LreB0dTUX8lKkmFwJYbu6LuwM1y9nOArB8Ckm/AJcN3DKUK9sTYagp9Q/
rzmcCpkZgo44NqPYYP+BBMIIVwEuO4Cl+jKGMDxo3zpo/SY6Jg1/cQgZn2l085pE
l0zOwcghcRg2AWinDOGxc2UoNIKk4EEmK488LIxeHxbU80Je7crFngimVBF1hNy2
RRWEZ6vTmy7puuPf79yZYeWhk1JYXUo4MsF9/v7yfJzAbxbT4fx+6SBg49VvgCZZ
gyUQvTPkq7qJPimx5ZdwF9gnDg7VSHERcNe60pIfndcjuc3yO/XkyB0rIdmLmBFs
go1GDBxN6V8kzDh8AAcC2gqV0a4sa/hN4+H73YDU4aortkhMtbCQP7MB/XIOD6Ot
HDGFBRFcrjNflTJ3T0Dticw0EiiBdF7EIet0dWyBt+42eDzZQXziFqBlD11BbI0B
16UBFmZIumz7vIglhAxPml+35yHk6I+n0j8OVBFbORuT4Miku7OFdRE26xgCCdxm
xc5C8vAaiwE5LfajENDRhr+MM9Hh+9jHYWkG8cxr9WsZKsr7uLr6qM8NDLsn4b+O
Vimu6AHEArhU3okMaOQq6em6NcvOd2Rn22f7SU7E8WGsRxcwrVKwKNc07YbNvM+U
MQ7vg0uROXd9R/I+MC/mo+lGX5hiuL0HKP5/4g6D61GfwD9zMlx5QbKDyoaf0AGo
LWQLQ/loVrGuGbR8acf9WI3f86Jo3f/gInVglIb1fjMI1/CWlA0d24PtN4hkmkJ/
6M0VTlWl4LXI5x+PTPXk1YENHu5SIBQq5fT4Y/hkT32lIyFKl4oVIb8ZZii8rNA/
5mu7ilwl+FCxZumKZkCN0uvnwtn2xLAUvzEircVS11rSBmCNP/7a7oAb+Czyt50L
GD+/Hh4fT/ptNq3PmdsitnVIaPq6rvN8kfXl5iTQmB6A/dySiS0bbVzdxiEZtez+
z6NQOhPwWIHQosrr6trO1gRqHhs939X509iNw2t1aYVaAjKcBK86EOueCeRmaF/h
VyFRbhTkxFJ9MIUxql1B8uJyj9MDEB8dvxuT2o389Ue6etdLhUVSzeUzSmzg0PAg
hEHSDpWj2ni423loSjCuEg722P+2EOdjFl4B5hW+TBnXhl62ZTXDWP+bHf+LVxSj
PvL0B2HMsRtpEc0miOZdqtD/GIHyIPm4vCvUHVgNTPoknl9RPsIaUtbz4Wg27P3H
Ziblf8hOkNXyK0jiULJ+x/9BsmkkFcyUWzE8VJvtLK9FkjpdZA6dOFKfYixih0c5
4zqQnu7hZcYjq42tC4aDYG1xdxA8WC8RoS/tpPfMANF7HEEq4rQtiND8/JPqOkdh
QcvWZRpWKQDTs6rQ0TUAlbQ9kB5JLv+bdf2bjV6e3HJ4fMg2cqW5FOXki/oZh6gO
vnAYHmeDsnLekrD8weGkR2EhGFoXUn6ku7l9UOxb8fbwRT6RCvYP7kT6B47yYZ/w
TSVj9JOiKnmPzRJ699UTl0LgoJ4MUwRLH7pAUtFRXfQzzQGFhI3twO5HDn/1uxRN
C56gvCSg1yo8M0MIw4q/zHNVXD3CUrCf11Wu4rSsFSCFCfhh23iPl5TXRuDdqD9D
JrnA0FuJKiW9cS6tYmD7B96l4xYF1npa+t9vfuKOqm7FYDyQX8VyEYIGa1HMzKb+
mXTBMAwogqOp3Ku7/hEKsds2og3rmSOLdaVIY+1QAumauZMOS2kkY6C/MZDPcjIG
89VcfwQAYp8xQXJZYahXNtbOehVHEYk6IDTrWEMjQzzO90ABGP5AC7AK6DLDlpGc
rqQTGhzHMzHxKRRHzwlDNTwb5XYbTqeWlTm8nTpNecgyGc7+uka17NTXV2CveStY
yQJrFqCrkuQiQM+RAUEFlbsU+C2X8IjDe2bOCP6Mbpdy6coDjXBVPDBE/TNs1QjV
dhDZxiWyi13NcuZz6oXhzs8wfRtdVhNNAgVFVn0vz1fppJ8VRvC8SUiXeCGJMbGD
UPmFEtPflaNcwA3Az6c/70cxcCFD/aXXQUgGyX6X8GMvuGKbBLzsygYxxLyEQUsc
6omaglyH4MPeZF6/jQhJe++/ckIWtK07R8x4mA1tcWgLQt3agzPhFojibvyFId9S
jPm8yZfplIOR9JZ0qgFmVq1GD8ru6+qMy2YoxZWiv1kzGI5PB7Mls/lOO2pNUqNW
2yXm84x1BjcSUI+9YbaBv+CnGKYLl+m+TMrc/OXZNWIEPr/sl1syPnjhpuQMQd7n
ErPqB+TwWi+ed3rTnysAON/4qbDmWCuAH3q7u1ShkBTwQwTDmYV6AoGJYQvQbaml
nGZiy5toxG3D0GuHV/UZo1mWwMl0Iivq0OUdykE558Lq5/uIyz3fC3+VyUkyUEjV
JmOeKprjokK64ZSYduP47q2PKTdaXQ98dNsdK7xieZG2K7ZoEbENLl9NlYMo4W5/
2QLA4Hv/xHFZ2HFVjS5ytDgfZ+CrP5uZkgTUPCKGK01xCHVtlGPAKOkgimDIQ17s
7BP7bOV1eeUO6aUQ+8EHkBVyBn7RBmTpsXVZzcuLi7sW736SATwGmi0N6nIOMFAg
tXjp15XIqt+Wr2fKtY2G+VEpezkRibXtiBFtC2q6HxagxtcbgBLEf4eHNv/pkqZX
zpc2xh+75Ww0MCQKhoCiBNBhpTFx+sZP6Aeg75GQyYdqjX3QZhpzk/I8gA3KnCZt
fgeuJdAgacKGwDwQN5ksmYCHLIhiqTp7RgMpU161nSZdTBqDRWQx27LKURANmHst
++WsXFDwycS5eSjdFUnaQOjmcffNzGOk1RgeqPb5GQCwc1q58gpbG/v/Sk0RyAFy
HTkzvwH6Gqmca9qS4sSxVlaz6go30UTX14P5kMZkNRHAkRPiEohaEKIY0kUjxYKv
8GTqNQJucjHKhstveRltZEMQBmOvlCW23skhcHstuPE1M6y6iPuR6NIuJJF5RA5Y
JwWYuiycWhSHvTUgiDpg0fDEbeH0B1oya8fnaO0bt9f8EgcQqBA5yyo+sun8l8U/
iWUOFkQBo5dIiVqom8XHuJlv6LVQj/TQancfsKMG44xmu17YmunCI6+5Kl93aTyk
C+wZcEGgf6FIA0pJCAo+gSxljsgGkowJJzagzNObnmYP5C5vdwZTMIwPeb4WB3bm
QQSi2t/CB6bIhGS8AH51+HP5QjIyOC6rsOnx2X6SQL9aqUAjnHCiRBc/YY8zSxBw
iZ3YHkjWAqc/79Y8SkDCWYdn7h69k5jU/h4Ob5RsIDUFL29c/Vc9EQY0DgAnnek+
mU9E89uJPKSe+Lr0iB9xHf3tGELztNudB7QSGJgs1MBEP74hGOeoyBUzKDFRZUxC
LCdce1jDVFuqDFJwFYAC8GuL1ALkMUmYIRVEfYOcaryDwE+WSsJDrRysYoYRAqbk
D/Lb9Yk1iMKaDwSAZdlqtHjcU8i+HvrOIM4so4IsDhI=
//pragma protect end_data_block
//pragma protect digest_block
4z+VFdnFdhK12pOC0jNjcAbRp/c=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
0nkFATW98QWl5VBRF+Y+iTS7qNszn9I+Hq87TN/IZxGb3vjX4vLbLlvMvE6kvu93
DUvlj8YJVDLzWreYnav1/2FDWFlsMkQfIcYfdcV/PFL/bu0eXcWJ7/pubgS9m/KF
cNgy1Fh3ybKjsw9JWM5h3P1ddz6drtBttcSuEHb2vAYWYH/6ly7Iog==
//pragma protect end_key_block
//pragma protect digest_block
yT1a0dLDWNFff/TV2xZ3x6+WAzE=
//pragma protect end_digest_block
//pragma protect data_block
USQG96Qdpl/k6Vh2j+OtkilQGfL3aTKrZZVNMpW1pxRgQhTsuwXVvSP9Bc8p3FKP
nZqP0sG17NqjXzUa+VVKzNKVMxe3gcWFKGn5KLTTIS54Oi9cCjnpfdK7TK6uBrqP
e/VXxHNru8dMfPKuT6NTRf1uTCIVJXM7aRHHQ6mF8Rz9QB0BKT7GPciDiSR6/y9f
7DbVsO4yiDYfTZvQIUVIjtEZ/GaVIIrfltqNS+zwsgAobM6UB840TYWQJX2MXrBp
TRa/kwEvPtzW72mjHwq9zpTkrCj2+9XYSgC0S7PywQHI1TVuCbp8o7JJsW0C0OM7
SZGVMrhC0CBgeElWuYYqpvgBlKmuntbKRlARhuuHh+VJMJfN62VobnJWQ11jF1V9
XJLAqmbctAuIXTHTUq/anXjDHKnJNRpXJdM7OXTxRO8=
//pragma protect end_data_block
//pragma protect digest_block
BWv2AKe521jvxqML1YHtSZQPG4Y=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8OJ2uhCLlqYsvQqSAtv53O4wuFBpXrB5R5kqwHflsKj/QFoaNghYr6cFtyKtmCaS
0pRZ12rpFa6cD8bxmPaICWAKhhd/ft+4K4aUA8JOsQBUazZhH4TCyNqKjTRB6wYo
k1J74qN0YzlYn6kx3c5d14qMPbyoFXXwe/NS/a9dM+NYwXYprmRIzw==
//pragma protect end_key_block
//pragma protect digest_block
oiruid5Eg9nhXcmuSbpkX1Qk/90=
//pragma protect end_digest_block
//pragma protect data_block
Pd1QoYFheVQxgj78KjX0A35pJ6TRFfVryS4bhsXEXZSZjBtwPEGHidauIgAdNvHE
eQ/aTerUMPC6C02+/NIcRgesR8cgGgkfkmZTpGc/QtjWAbP3xdq7loJcliCnY08n
IUK3RCu04nIQAXjkUol2Swb6QEREtnaLzZf77V1r8YFzAv/hFfjK6DLp89nujHRA
FDzLcZ63e3cqxbQKo0RFCiLWH+E2s3mSinmj88Rjp6VW3toVq+kzXSd0Qixcmtd3
wri8+IOdGwWqJ81Y6Jp8j4NI0wGnTMcNxUx5vby6PNhjcvmlLwzF92lejcFzjVyC
0PhFlxaP7/yNZ1S8ltJlVaRTGsbSAqOpvpxt9RZ5Hn9hE6dVSZpn62ij90E4nKRG
OtFBjLVSGTZe0aLMxLUTiSC+dirF19L6CtM/q5MW2oV0AZUFgNafZ5w0iuNMakRN
yJoBKyfRUKOyWCRJviE1DqQ1xDEF6YTzRlDiExbyN7Jvp35u62IM9EQC0zSmhAtM
XUMKsLasww8M1ucOmTmRRlE8n4ozAky5Rcr0ycyKkpYg/In+Go0b1qFBStbllura
a1UGvgGU9cB8/XH4h/b7P2amyMJxxdPKfC2jSqnn2NBjeZgOA6W2h4Tc3rdXxEiv
IL9PCZkSk0BKk1MvCgRVoh0kltroqt6Q8yl0qlWOwXHB+0TOxzvedt6ggyZII3ws
ciKdLXKAnRTpgyUFE/xRAQsoE/vF2IBxj1d45wTMYNbfJK8HIp8Oou+graoDjzfC
SrAknfOq9W3zevaxwpVcFIlZuzB1q7gOoSshliQOy70OjkCWVJVhnYMbyzna/k7S
g5x6Qk3VSjLtTo/jaD0fJ0v7IZmQp1A/CiDvl9xrwNkQiTr2YBwO/t/XR7mFDpx+
bGKbBCUPF2UHe2KoAGaiyG9jSIVbyac2gdhdd1CG1EWsuwyX1tKJzZmROjmo5u7X
J2zMBbtTxb/sym7uIGwx9SOCkKkWUcTWFxWK9NdojL9/ox81X+fTeyHk40jHnW/o
4p+FoeaOJIe+QFjB5kfzwIKYx7zOK+dTL8qDGDKrosruyE1XqJMPRnP8wmSD7N+y
nPvcRTU0TC6cq50MzGBubwITVc6z3zKyBerxdfMc3Ek0jAE1Mj0HYPH6oErOhLqt
pJcCIKMcSaxV8uwIFXYWelOZbTxeCcRDLFlapOF4OkzACV8gW85+97B2b7r07ami
9AblNF7GdcTjg9OMyjOCNpHrmlZIMclFzkbv5C/SjNkT7jy2VWrOMc6OngEtTEGd
GPteTRKYFk6Bt3IS5ZzLjFbZfMaK7v67Ok1qGW+K/+PYBguty9LsvvHZSi8DsFfj
ALCrRCIpG7s3jnpiGi2asCLSWCnYwyZ+5YtrxvOdyvY8DaD3NvL8iGF2sn4G1J0E
OMqjy00RWGgBoPqzWsYripU/Qn6izRjA61urmhHDnln6j9XO143VBPsfxvQRfQMZ
zBwMongQDeDQ7AcvADw7Jr6DBXXF52jqy+y8zgreUU2hfjU4UFLWfM+lp+3B53ZE
a2FmdJ71j6wv5JGdI5ezFe8BRogqB8XAGMY4QHq0+d49syb9dkruR1tQQl+Yzg0g
/iGl6uRDJXYHpnyVUNFFTW9iQyFAkcQ7aR4YbOkcWZRDY8FfMlzNyba0+VGiMq5G
CPN6bxeeX4Ng85TADuJvUef1GqW01aFt5goP257h+R6dZPZSdA/APsUrRUeXp1iC
fW45XScXm6rq/Z0+/igGteDyQuje0kcWz1XeWHrtf6IkPy0KiYygD12Qv3Mq57F2
pwznTbh7ozDl0kWfhyfcVEwHC6JinnR5x4RqVysRJuBoDu0Z51Qf8y9gWBhcoGKT
9+MZm7o8H8jobiwkDr2UB2PiQoLqvQk882sY2kdHDfU9gg9QHBC6nsPhmGVHVsag
HRcxPVGBu/sYjC3tDGkbgfe7hsM5GOTA9D4OXkcaOeIDUT2l1OEGTxwPD91VyTfW
Bns25tANQTc30SJOamsSIBpp8JlyZuD7qyWtj+00dQJv14b9LkUEZ2MsQ7xpEz4D
wVjOcOGRlf1DMSlzSdcqSz+3QiKHyYM95Z0FXEQZvTlH+I9ZTE9vuxuLOD1lkZCX
WeD3DeiRIQ8NhTlfyp90yWG3fRXQo6PZgkrXZsbAHSke8lFgQMF6/0M40QU3nlJB
sCO1b8iHx9N1NXwYYSiOcn+QYeSvFF2Df4qSYcPr7kHHMzAe6A5Tw1oVypIuuxRV
X7fib2bC80ETrXvSLeaEak1atZvZpnQxX8y6UHzJKmM4B/q8nfJyi6OoBW1Ylkq+
Bo7+PuRl0L0tqDy01/afwsx1I3FLLtYgCKvC1ELuOp+RHXDQvRpmaQ4BxaimQ9ZF
MjJJW1oBF5rPTGoZeM79yh/SjYcB2bLZ9FpermDfEtkusTGeVLmu+09VGxTHBhfn
MzAJxfyx5JCHcvDnIN8juk25dmn5JCDD3HBBCiBoxh4rWAB+C43JO0gUA/2jTcfz
dZ+9bEZOdGa7yC/xwZjGU7EbG3NgHpp94hDEkUKmHxCqTZ1sST4+Tvvo62fBSHNC
5fSyIRE/leC4noFtfOHeaqylpH7J4w4TosopxjI0athPinAxBvrLOzpPiYd2KOvn
7vbfJpI3kDI/XW/1ztbXuyAdBjXY+FE9h56eG1MRvlnmN/xHCHrKCeBvS5ODfAzq
8ZxspZiqGilBX42ydpzkJyAy3jcRRdteoBD7aa/2N703QRqntxok9rWeOJu3kDWm
4zFX3co2ooh+UMYDSbjObK3X8eBKEh6+Srg1uGeh1h2OaphuWPfr4ZQDAZhsyTQq
SRDoNMQBvezzYRFd3PJw/SSUP+fxnxAlNAsvQTxWf7V9JfawT4RoO7HAc4wfI0bB
+JpSBwkolJFoL03vfAVzbNGD0qhHhBgMJXy5WoPktOUW9cdro1GulvKLQktl+tXI
hddQkVpcA7KnRLAOCjAwlcGhRJxfcOpFowmJckMWrX7M8APCjXo6XINKPUiSIw9Q
pSw0l+izfF7RPaTARP5oXiaLhriQ4pP/tTSUFdrUQA8/z7QbUkxnTk+LyCuQdaqn
IEiH9lxA5Vq7LT/fuFS1AAFDsO+4lX2WyR5tJZ8sxQcmeKe3k2WnmDEQppzn403y
zDpT6bq206FAx3FYIIFNs8Bx+nNedFiEd66wGU3E8/eUQhNviNoRxonc8peD/i3H
ltgSyRB28AC8Wl3NoGMZOGZ1A/tPr108GS72vJw76k8pJbiPqbarVww9gagW++rR
GICz6Fs/vjG7VVACmkRWRnRzj7aw+GNeUWzBM+NYwYHuM11qd6EzkWZa7vvn60iJ
blcBD4XVmmp+SZbhRYC52zkaa1yLGV+mcJyFG/XuNPJoxnJxDnwlxFkxgvUt7jCe
vJxleQM/OWrNpUdAadeTVgA5AV/zKyGre+vUCOHCSWOV+ygpr147J157prqzIJnv
rHzcF4GJ5kuK97611iQbvzIiSlZ2B8C0h6Iw9AnFOH+D53nCllTlhUGlO2K+kYjV
IJ63Yo5VZ0itAeffvbWvoAqTj3wPdsT9MY2aRwysWRdcsH2bU+62+ODwlc0UMFEJ
Ejj0JaCMLDrvZb+R0pNIfeJ/+cfaubj7Mhrf1eSF5NVZAqeXCsIH69PrWNVquksK
4i1TEbtM0x9Tu9fdkzttr+frN1nsj5OwQaHGivBqqf1KOs2vrJAwQC/sct3RMrLf
UK+LPOKaELq/aaNt0SdNz3JT232EC+MWbNZjwNTPwTdu7XbzEXeQRChEcZoGvGwV
yln3EeIkWtHPl5SLosg5byd1NT638N4y2FJH3XsP2fnDmaeZg8+cs35R24tkfLNm
/cd6aw+RkYoGY+bdCR+m+zkvj1SZkHgBa5lkC/WBUUQ1j2S6mR1d/sOUoMOJioWy
DKHVuDhRbPXUJEZhMHRNa+yRHxxQrOZazKrQBO62j4MGpg+ptWD2uBzaDCesDukn
pMtUNJ2Z9+oHCoVytV8GvaywcSacNhUcA32Xt9nqqqA9YHFE/RYUSvviSmXhOwlF
Jg3W2VLmevquE/Yyd4Qvt485vFRosB5mUAexhJBRw8WtNALvJO0v6JT5ptls3fCc
7d4eInsCKLTnwqcLru5hKJyQHQXs6NehNTOXwwlaLzo6IvpUqu+AfhVEzRbN67g0
sPkVlIKxDi6T9IhljiahDXtLQwiHt76q1q7UHPKblAVHNEs4h01WXFMGf+w37wCJ
8sYlD+CFuGcJb+21CJGCjou8vxWg7v+umD4E8WH7JD5gZunJCzEpQoXwHfbrbGFH
XbISwhxT7DQBmJTPyd/5APJugYpHPrFciXsk8gafSCdloppzLU8qiyY34KvLM6JI
UAc5nrlPyj7rE1MKjt4TPLsWEk/tQGZq0U1gSLGb9ET+uxJUTXPvYQ3JSfnSUFs2
dTfylQZjGYRnKqwmH7EjjLM7OjDi3R++YeAQOJLTTk+JUj62AP+dKk21K4RdgXGZ
N+mVwK6FjZ/uTGqO9bHDJuv2g5Z6QLfQ0XUSSmDAQXVKBQmrA40yrjcYfxiehywF
v1z6rueRiBnlB69rapztE3/tSOXONM8Of8Kttf1jk7uh9aGKZ5I2CKqF4JsTiuWW
Cw2T3DqbGlIec7A3s3N93xk/WmstKLEvC6E+R5MZDLDp+cNCcCkUbQ+vOxRlBTxl
1i+jQzMaNHTofP/K23Jib7FG/PNNyGDfxoNJjRatRHADWIwkdnhSg50UjoJKcPsX
KjnFao5+8M4jxHqoT0csABWn8SciMhPHe0DLDYfEShkK4AOvDPdWr6BTlNXR0kkz
j4nVBopi14ECD4q79QIp0cHjaxNRHVE/78WfpAa/dOmAdUSxW1f9CmsLZRdXbV80
aQO4OKW2elR2Y/J8JTpVnpNvUo7ZST8EBKGDbnWjgs3/PJ+Ewi4iOTU907yaG8fU
dls1wGWB6sA05gTy90kJ3WD+OmLQK0e7AVTAm1hMdk9i7V/ZoiAF3LMX8IimIoyK
HA8gte3k/KaowKnuWbcnjNO/Dget46dRrTHKjzAV6gYlna5pbU1lXMJCCB851APG
ox8uq62J8s6MjUljO17bfJG3s2mWdHRxYLmeQRok7ioNeOgl+/3yb5BWImQamt4o
77xCrjvf4bIejtGFdsY9TCgrk8F7PP2VPQ9nkkVQpyR+loP90v3/A9hadInSR9Yc
R3gxyCjeg2pqtfr/bFbuMNt7H9nmyKP/lz976y076Xa5L8cqLG0VoFrCMOTpIDkt
PHmQWLCSx+nwxkW5GmSjdai2qUgrs75SdI/I95ny3TOutNTVTWXCkHrMnKkHRLFq
Q5Ds5K8Tf3mCVJBYNII6HdWrybUo/1DCtoHGO1CIbtrd4nhA/G2XNJGVZqYBr3Ja
EmCJEgq51VYEAl7yBp1LQOcNm8G+ESkBv5sEgXEqRYFtUCTNuPUIB6p+JPxPfhC+
qvQ+wAu9TBTS7i22wRYqqPK/F1WTpbRAlzhNE0BOgBSvQPzW3lPCd6pFXBcvz6gq
US8JOSfpZoBpSI1MgAm0Cqa+WbGpdw4w11LHsDG7+zAPn1srPok1Yzhoo63HxuAc
wzTWCOIS2y398ASWgTCiR/mNO+VLs+6xL8nBMPJWc04cT7Q5q0YVg1tgddIjlIPv
3vT4z6SiIUsBqYM4Dn8BFC/B4+7/T2g17tjxR0tWQCVLP7wLl3/o6nJUvyEP+z+W
naUtNs+9b1cQ0ABi3rpSim6okR7JgM6KGjGp102TAz9LHrKEIwC326LmfgOb7OST
t1j0NESFGu6kJIzjs4ITejwGSazhzPaRVpm+Wsg/PrdyM4bpVEiMM2A3qic+F6Ii
0ruoQD2PsdOKK8SDZpdt+HNYt7yvOQBy3OY8oS4lH5KPeREbqgCb7+/qHa8C5gA7
8iVlMS+6cCkgAfTIc2bSx6tf9ovrPkDdUFsQ/XxBEL40fR5CikSolYFkkB9078tn
If3c6grKr6Ls4l8F/bDMUveEoENV3ikK6mj12Tu6Hil4uVOFEyhM240YQetMY6Qd
47OeKH8+GvpEKzE4kxKrTyB+tRv5JjQIWKn/tV73ZR2LOEadhaqtXEmN8cVu4+nu
p1zHerEy8/eOTwV0lEzlCJIJ9SpPqy34uLaXqpVqtwXhAmBLA2+LriExEKoyv8KZ
h+KojYwNp1t3ZZIFHU1f9J36mORVD7I25jPSWWcwkWg1l3s7a60+4HHz+5eudaZq
7j8KyDTyYs1Rqg/jaUpVe8I6RJmSYjlb09YXp8AjkXD0wIclhaG5XahbhrhD3BBz
RNKTUnFTV93tmToy62hHGYaEVBl5UCSw6iD1Dj1Xl6Zc8dM4Lz/fSNFtb4PgsB8e
BJq6nW0jM1Ceu/yc53OIyXYEAxG4ldfmBjdzPuJrihAzXsYSWTZmRLIKXp3FVUGZ
eas2mnFiP8HtDHsP4Xrb0W7hihUwqNdR8muI6DVY9XivVEmmPI2NYPEyanCytV6z
onnfFK4Pg6I/hce6Tjb1apmNgQ5GDuoun04tp+cXEwDh+pG46T6zRELHGXNPM8t4
hnPs9a79xOXUPBhB7HZ7ODxo7BweuaWzkc4/qr9cIC2vVpl0YwxJCSPK/Adm1+87
AnzpW1tcMkkk5enOlsVHpO7eS1SWsd4bRkQ2Qy2cYt/ICwIZ+vZbWUDYKRGM7uAw
nGso5C8SC+jd0+mJvHzDlxNkyXiBEEhgHL+ZSs4BlKA1k7qYUaagMqEBfTsi5+f1
kJQcMLOBgfWP71b2E7mKdABdd3+KPv/xb+rJsS/n1Bz5IwQezRsXOn4LGkHgT5Ig
I4OUmyJEjyCuHcifSPbkfURO56pAqabLAf/cpy22azt9E6nn/IUdLLsu6Vvq2plH
jkbasaIR72TSWR/Trls2w065nEzlDHqXu4rZr5N214aanHAPRFcZpyJj1CqmCqdE
Px0r/rtq8xSya+bAfWsCyWGi+MHrlKKIcJxpxpJL1FH+3Md4W0cQyfZ+ZtKu1Oaa
HFwM4WYv1jMCCznUS33RtdvCUViAATN9dcdVLAYR+WPdt3B6c8l2QoIQd44i2yTg
51hqjSi2Wz0eLWefgcM2u/IysdveCr0gM8ruTNztQCLdCY3vlqzqvZWlEyLvzSoE
82qLDJKs8czNR6fW7PzAX2RJCZ0wVEYD1agogc8fnCA7Trzgu+z1VDsmd7k0G+Te
cWope2YUriyzkdOwbu3oOAMMXwnMTu92TbBv6z+0E4z4RfSlcOJAI90813zZ8L/F
G1mDgUzwQ20toPlbGLwztF+4MXM/1XlC4ngfJ6RwJM18Oz7BDmhMtJTGU9+Xt886
9vwZGvJs5cRoInNYZY1gwVc1iMiHtvA44ep25T1xAFSXIRCCf/+R/B9wGHnJJPL9
MYsL6D7Y5MNtBgpZgNhyYi9pGLZp2VnUgZX2j6/g0CyMSCZ4Yx1+BvTuAigrW06G
/2WRxfv5Q+K87JCKliJep1GjAU7z5w/3rcPH7tIdLL9qbVPcOda+cYUhyHLjdQJF
FTTFirlhBnAF1JUog8ZJ7eGCooWJ4NYrTWmWxe2SNFwxb/uoTBxwLe9lDjT4ZjfG
Y8iZVJLqewB9DR7xm7fUyFMVHNyitfCIqBjPEdyP4NCVZOrmFLBeiWYeVgEaWLVp
uupftIXBzio9VaCwRlQ+70M+tYd2Dr4jX65l4w+siTzn38yOXCuGK7RxQnoCZTBi
6ux0JcErCinllSnZygwhxaxyqlf+02gOVS1aMdcMsYZkpH4wBqavt+uICTt2le8J
7bmXqcXn8APrHhg6oS+JCiI9vzqH8axE/sHt2xMV6hIQP4nL5sjaPFSmwAA+yci0
QDCSM2EZvlQRm0evX6LiVKpEydfGjOelQtgVS8oGqf3spPUC8UODMRxxa88BBhNZ
wOFWXots3FLzlu5Is9Oo9jMVC1RBgT8dNSfJOU246WpRxRZnuBZb32LUa36YLwm/
BfJUHGl6xQ+L9s8Oc4Qw5TNM18Ud21r5yZt0Z2f6gq+LEqDspi7+mR3ezM240EWp
lusUJuFhuf7Mr0N+IKIUhADH/KL3Su61u86HUA44W2h8P2S/Bu4dEQJh85ygfMXr
UkM927V4r2mgRvzChyrPSLCopEgBn6eyOrGZrUDLvcPTue0KCwl3sX6pwnF1JALE
BCmnPnPUkBBqbzm7TmHKHH4/9Kq6z66jff747JrcTXZ18u0NGtDcSyhn3HB52K0f
cQPwXHONqox4ofY7oyljB3BD6Vjqc/4et5PnhTKst6lWgakJhP42knxaWNbPqrdz
5Y5BZWjP0jgwCaohBVpJM82rqjRbELJ3HN4804HPAE2NWvO3u8kcmTNykd5eU8g0
fkNtllioVPyqxDfUAhCl/6Ils9nTuFTTnn/IwG/rxerXqQyC752lSGpYOt4B/1yD
lEIQun5hjXXZxr2LihD+sbeCgVzuWMQBPCZMON3VNeNkxuVCdkaDgTR1+zGDX/GE
uumGWzn2ZzC4HeXesyyKMxA367tokw2n5I82cIJ4xJctPhBbs7bN43egaZ7dZIEI
sbw9hji2N7587IKW6POiQFNTBKIO35xsrRWU8J0XV5NKhI5C4dgrwVGMpDa2HGha
xP0QtYdEhE8RNNXDY9+UqVHFlfeQ3TBQiQIYzv/UHDDrfrQg8NPGXuSd+q2MoxVg
KWnwnTOS5A1CNhyvyKc0VzEZ0XFbzGtHXUk6e9mlfh8Zmcm2aTDln1dZFo72hdUY
DL+RDv+4xtQufK8wALG3NlT0DyuM377rCUAq7n41+IVwcnf90+JUDXcboCjDE1Ox
vWeGIYYM9RKHzrCYb+VJ31mVSnkthP2sOPDey6CPzyTiR5UhkNnb7KL4JKd6wIPV
6GxkUcQOJ+ewE16OsS/sTICWmpPjk0amNvEsRX8/VvfhTPe5f0mR9MPJBn9na4+1
Ot6pBn2IefgclmY5FBF2qK5Y3fXHu8k46YWtAjIES4FgNPrTrPPXfTI6jXPKRvib
lwminC2DcR/Vlt6LAcpNvcbCVMgLRSUpIyOPod0vEt5OyW+NsUBqFVnrwqVuEWpD
6nH5EQD4JF79W+b9rE4A0/REeRvXTuqkn30nMaKhYP8N/wbmB3gv0li0eM+mbJ3C
eoUPmYSX1dn4xV5ng+DEYqkGcgAh47oH+fjVAGkOvhN1EV7D1FwyR1X6n3Ci9Xwg
QVuSW7o+5lLUNe8ZUOL1yqf0trCBKcUnC3bgx+ZUi5uHDktyBrjrln/8pL1xn/dU
Mwe2RVAN3DTOuf4CLqP8UWp9XB3bLAMZrhdqqpGb2gx58jWicAEusCvJVSYJ83f4
EpQKDq/jLtXZCyIy9SMmzsjbiszV80OOY5GEhClH/m2L9OH4usWcq0jtqxw986ev
8Vy5CTDAADOJGRO3xBrqEjGUK3JY0ddYxtGo6LvcNxyl/c7L5zBs7DV1s67tPZjg
TsvLwkxbNG5o/jUdQZOK4aQ7pTaAmybT3N6LRp5d3Q5XQejCD++q/OXoFMz8iMW6
GJFxinsBfhHyTZOc3VvP8KmzLduMlhd4Mw+O4zltgZ7BSW2VmEMVuXVe3is67B1N
+b/brwtBJkpb1oKakwGoN0/CxutQ1H2Zdm6RQf8LZb6kayKhDcU54agpMtKwflLU
jgrAiNyKIc+GLbe8aIuDGt0kkGTsNKWGdogwe4OyVCt5/Lq0mkiUFyw5Z992QWM4
vp2t0JMh6bdj9PCqX1t59uuL2S7l3e/IllrR9l6nAn0rABhEoeW/gytNM/H56KDh
5J8tvy0yTj3M1uH87dlZgjaoTLS8vi8yIDg51I7VptLV2Yi/9i0e5uNmzTO5Pszs
ITjVjh6J5avfQhJCjE3TPolCORvtxizv1pX/x6dUNIzWgb/PeI1ArYCEUNvWwPG1
dfO2MAAG9iPJ0Cf5GrAAB8m8f0hN/29xkU8TswegOBTqJQwhKV0ty08Z7mjJrrFu
1Zlm2YC60YpY05wGR++13ao0+YOu5I5IabiVF+PJ0ovhlhZBeIFOTPZBbulmCmZa
2kXRY0+Ibm1IZLri9OdD1Xfrb32CCsqbpM6OHsdL7JQRKCtRpSYZSDkWopO1BJr+
K/fov4+w5VVc/3Cm4Q36ajAPWNVYPhfPSu9Kn3TqT9IlO8e/8c2jXPzMhdTdsUEJ
ZwUoyyfzfAA8DaHzi3El//GEQCKisdCGLy3KR/mbvvEsieKuVcnLsH1zJbea88aR
pLCNa9H5v+mfsyZRIEJSmxuu1EVi6Q62LYH1vO5ZmI8Z5U9IZc1HC6aEcAS136qL
yFp/EQC8kTx2jdR4ATNo2YV2/jKbi/CGHIjDe7qo5PhIETHRnHl3EqWiLp35TFP9
RCM1X4Td+RU6Uq6/4eh4rXW/VOE2RRS3ywTX16uhNa+bDpND11S+Hyi2oWagHQEA
ORkl/WkS6STJep83E5GjkcpbIW4SUBYgu+T0uyMaWWzCYbqniJQMOOYmfskPrwxT
EzsgdihiT103SZ3dGDevD17hHt1Oh+qJk1bKfepzbImNggIb5w624I62oVv9uyfA
3MBeTTfTwEqoj1Tqv5znCqW1ol2JfrW1A5Pa+Bp48r1x/Jpw2tAU+srB6vg+jT0z
S9tYyCs3GxdBVncGnpgsESeJfF1361lcO3jpguwAOBmg0J8R4fz1pLhjLafefFKS
ah2UhOhTBqeSIHSOqq072egLscWNVMiCdM2vPzB1Ay79/AiZVcdy8h84ZuK3uCVr
TpORAaSRhlzfByx0A//F3JvBdG7Rks7JxqSK8I2FbhjL8pVfbnWTIy5x0Jibd3gW
K1ItE7kGXIm2hEUYhZQpJkvE2INBDlsz7BR6YIAhoVe5Y1a2EabIUZVZD8VAQLxr
9BxDyrvdy+m5ZH5Hu5hjETwRO1foYR/mwdCvCVvCBz2Br6lPJXtOr7eBJsWxBjwQ
vMCMwx9Pn6JprKkE9F8nAN3E44IZ0tNyCzyHtamvukhxv8A8oI2Tm+0GiEZ/7KMo
yR0dvvxvjSDjZDgmGkA0n7bTyxH/twJJyXEwHjU7K/yT/AFS6XgqOVbUEr2gNpuE
hwMmZaAw0lXJ5Z6bCP7sbGEsOxS03/7BLJOtYx6bY1zcqINWeMgM4G1duCSTLjzN
J7PD5gRjJrDoe6U2y2GK2yUtDCYojnjtL53Nq6Y6Pi1f6vwg+ePYIe0bAjkYw/3i
Ty+4uIkyMKKhyS6339MgcV87/rGgeqfXYd/xOwjQyQzj9z3Ga1ykF2OOTfwo+/Og
gwrF2XmYuJUkWxqs7GTphkCcoVCOTs3U1BPbOm1FtseoZe24oGzN2qTnGutk22oO
UXxT+qIpYf1EAiMfqsMuF8nFccqR452RZ2emqWf0QpgMxzZFIhz9uzuyvIMJzo+e
KX4YOT0fN51RyQyRgRm/LjWAMHIagpShnA9NzovwfUlsEwu+tgwmxm8J5FcYCKwn
qAuQqe78NjuVvkp9cweloOCiVFT/N6PlydxG6fOOB56X8mRt4OAXXXL+sASBDPGY
R+YIid/h0tnfpalt/FRab6zFpPyW9UYPU9L2s6SE0qtn7qdqiWoPtBDuDFTH0IFB
H6fvWg4eSoTTxVkJKiyhPILtvadCUt6tvq3isq1MGqwgEN7PrngnsGOlmbiC1SCx
lVBceJ+4UFlecPnkqem/hdfpv1Vw22gY2oHfbuMVj0EVfAtB1OPAos/E0uVht5xD
QbzDqfQ1ozjKQzPPPdZklgEws3bacJCHUOMHX4KcEXsitGQ+OId8Jp7skK+f3Crw
bDnTl1HRyGOoPiqL4g/NlXqvHvW7GwWxkeRCvSHgSn6vo0pXjAILvNoNBZ/PyU2B
aqGxJnoskeD6l9iC2X/uPx2poTu5+V6fr/60IxuDJB5mJmDYz6pk1xTL7HEC7KYI
Vw/4DeMo+MppjPg9Ax6N1ewEVmuFdz9TcnP09AfR7fuTsE43iW06G8OMe1H3QyxK
wCtk50oyjHPDSVRylKSQ/nAqnGx+7SNpJv9oBkpkZCfvhislpDwDQ/n9eDj2Ny5U
TFLDf6ocCr4oM56C6EsMbPrsGk4Wio4tOHpGpEvyEmhPIstXVcLjPRz7H88/G1OK
Kbj0rBz8LQUZfyFNDUYam9qAf1MHD14Hhw8rYhSrmU9n2DEYMn5B2FGEVzvLLgBj
hbk0jUT7TQtB7YOZKb2Zck34MPEB1JoLXVnqbi0mihQrA9DIT2cMz5maklkpsYiT
zt5Y/AfmXq3isuPVl1zQjD5Y45MkXLGEbHWoCvaNXL2h3MCYAax8BTjQlcctLqnk
/UUwK+NKA45cd+u4hQOlChdiVGtcOYEv+hDFtNXkKkm3+Anz1TziecVNU0tVNaFw
cF7C/0ZUAyFzT/Z9yYskQlN8wCu4GYUY9rjhY1FbtUb1wj0EVqBVvaeo7HkIN3Jk
QL2korXmM5VHa0h1sICoW+y7Tvp+up9mIp+jta+rRKNHi3dUZPDI0Pjor3KM6OnN
yZyvxtgDN/6C4Qwrh115fklDJa/jTOy4ZwBXOh+/wWLzSWY2rj5/2J9KIwBEMebz
0bdnvI+e7OibmmMRZdhEuFUN/i7Tz9dNXPMsIVIkr8NPCIUw3GiO1GiDZHUn0n8B
6K0rjJR4AwdeDv+80KStlcdjkcTcYY23LESZAmZgJ7yP3JixptL2Mq6o9d8KPEgX
Ne9I6gfpyt0XcVYpalDYZQukrQbBAABii9THXyI0mY7ScKG/D3/xiczx60RrcBCK
vlxkmbiOaHWYhNtGS6ILEWajCxaCXPzCxlbqPr8ldBLakWZp4i2Z7b1qPhSVuP61
jy+sEHdErJL/4vVMpVf5jB+gaiNGv34goc0LJH4IovKT7PRqRS73YXQtvu2BweFt
S93vxGw9lK0gtKZA8VDPrh//f3q1bPJ5HD+1/Hoz8cjY9QT+dB7easGzDbJEQTBp
ILBNFMpnR3KAWO3GHD3hpQPkIDXP6KPAc+bDk2NGQ+i7lW4xUxgd6NVan3HiAvFI
/3gsXJcW2oUIipuje74uZ5wbMmbT9g+oG6CUmqlyNWNxjWc4Ybm0H9t7D7I97B20
RlpaVtCKJS0/Z9XUVF0RtiYZAf6T+45DcfBtirBUlS27tAPZOp+Y7iO4puclf6ty
uUFNjR9eGrUJinTVtTNejIot4z0dSdG28SrFWJhPkCJIjdmrh0KMog4z3zQDbz6q
eZAyAPqJmfIHW5sUrco4C79RoGwK0RFJaV68NHXUREqiYdZgI5w9uoSK9acz5dCq
N+/ttj89BWUI3fGFleOTqoeYQ1kRSlSDrV8ZlUdNdPJNd3A6/FKkDL4jbhVKs0CC
109T14ZC/0itEzJxQRq6dCcjgOcaFbQefbH14TaJYE20v4B1IAPdmMxZqbmYJRbr
YES0SmRtDNUY04P3gjE2F3Dfn27bu1lm11ujyHx1Qe2WGcz7OMFB6utWcdvInlym
yGGShxWJOADrF9ZBS83OrYJyds3VSliATCX5ABPRi03RmRVYfpGHk6ZPj1EPmQXs
49RXu957QY+VKAW2W5Zp7iYua8w+gxe9oW0Jyl01ct72VTWfxa8GvJcSYSjtB7ja
6eeEFBq74taJ0HuAsg1nXrouhXRvq0ii+pHnlk5RxDNcCn7+iOy8x4a0hyvJwwHh
pCVv8a27mPkw6wpZh3Tpa5Rlc38fj5YObrXSsXBGdFuFqYvtqtYyfy6fQTQaHksw
egrrf3PBLh9EdK/tnxTu9Mnza3bd1fEFSiPHzi7Sri4sYpLLpeLQMlskJ36aKFB1
rC4lTLCUzBBgejOYd4En/YNv4W+MHCOFKigtis17tCnGP61Y8PUdRHgGroyzNNa4
FspnqQQku7Y4CQqzVC/mgvgkkY1G/k4DIZupmCcD7g4hkFRnV0Xcz3ob2nvrNOHR
Mr2pmYmjLIMxFNZts93i7+1/Av9jNVSjPTlttk5yMrx5wwSp1Urtr4UD7wwFwQP7
yp8axw/EvNfXLqt4Ry/ID7DPpwCpfSvDrtdALM476O/eomuMTunmxoGfxyGBu9jd
rrlMWyI/uU1w+fTs5pHQZDrzZjZzL5d8nWHKg2K9V5ug5J0sQyMzW8+lvu6wYn7X
FZBKwbVnVSHHSpL3H6sECH5/UfJew/DH+iILw3yhI7z4kwWxt61124PO25JdpkJT
IhN/IONMmanrFHujFtRUR1ahaaxLbmUiOCC7M++Iv1hhGkvZVMtejsyQ6RrCtXNt
gjgc2I/krSuV59MbXd2PmSZZT5nEbaTv6r79wYUhTgUp2MR9Fq5N4PSzpBptSpYf
R6Z1ubGfbOiBQVD7fEFCtWMXa63d2REMtJgm2WNnbGcdIrj9qfsZndsdRCJ84/8E
+gG3/ZzAa6bT40kqAWMdI5i4VSkNefQVvxoW1qksKiXY4REBwTWyk1FnCF0aV0R7
fucnQPoN+KziFFRaLbT7B530Ppf6xcQIRSYaq+40Q/48x5veMKIGfCRhErPIti1M
NoCpSIwiPe5JeNInvRK0Mg3hJKReoG3JUzyk+hfDjYju2hj6oKuhTD9EqWX1lTRv
3vg2cfJpDTHtXn/0VKOLnszO/pjWe5towMrUYN1PsgUMW4S7Z3gytE0+wj5xKamb
lWiuTJmV5egUPfQhEhfHYHFOdOYUVVwAoih2cOPd38BnfHBTKncVvCnMMXwe1+Yg
KzEFk8OFqu3tbOyrvt/+1/6WNntmH3fQ4nM86Rhq/aLDROIqXFeCRowgov7ZdgF0
O3FKJwI9szBQhaAZCZ+ouSDZgUe39YYSXpJsZE0JaJwtOE96npOQ1aDutD0ctc23
TNIRb93eUXL2t0+8tJ1N0Y37Riaj7uk/cFHlKj+PByyNwu9HYufUqQ28QiI5ZAZY
fU3GEVjtNJCisvWZTwVxBPKwrCEayDjTMyTCSTOsvNzjQTrOgUqwq3O70iYH6pp7
lknTmidyr2cYrhSB15n5R5c9bspKN6OSmNP9UUF7hfGZwrf9Gbs4XhPvx3YQ4nPT
lL/qbgTu/XCZX2iWgnVTRerlzv5SMTlRhB4kQ0UQ8TH6vqphD0O8+ZKlFdOdtc8c
4ZVh62VcaxXn3O3fN+nv+uMvN81w4ieroKc7YO12oEhMlYr6ilTB6EGDl+deO0C5
L9fO61joMsPWZN/io++msDX5n+MdCNn/6gC9nwpB2BWRJjaNBMYPCDjNMblS9ysD
+CSqABufJMkhT+hAAbz8vs0rviO0YQubwChYY9eZU1k9ahkid+2OQU5vFGMyXe6q
wKVpf41Zbx1E6qzAUJ3q2e8eEpTUW1CaOnsaZ8YsYm1x43JVFX5GFb0E9ZROHBl8
Hnffy+L+nauGBEASpoMvOGjpBkhprm4v7WOrItNP/py8C4rW8Wtuwyr3X5HIY8rs
AbNZgDZXYHWaiojtC4mxpNiVXiOOnNTTW2PAZfQmx47LDCqU5WZ0LnlRumoUAbG9
ac69kLi0eBSU28hzzzxo2zVEA2v4UjcZ4QBilnVumzgLjQ56fPH0LNstEK0BvdvC
Myac7FxeAhAvV/gr7DIPyERaiyNc/wv7UvCKdEc99QEdARgiiqHsZ+b65rp9r4VO
mYvhJ7CRclzZj8L/5tSgDFGnSP5RZMwQBBL39I1ugVNm2c5o04tIBFSLZC0Olbux
j023iUZ7XsCKHphzrxypQGTlbKCNj9gR2CWWBMFHTHTY8/e/ObRa/ogj2Snel9Zr
WgnOi87nnMaCBiYRmVBzNd6Mkv5ip5jZX8L/xNo0oUxCjd9RABpb1YTs+msuI3MN
b2a+Z3csjFn5xiruf6VZrV3nbjhpe++bK/waP2iq/CRF/hg7BvF7vyuGqnIAjfxA
VYWw17MqxyInGXxZ3eYPjWZ2Ejvtp03CbjkTQ57wkW/YUjap6vu6ueIFhQr1Tk5y
6X9khc3OSHgIEtWL8ZgMj0Bi3yVQXoN7o6xdlJGIOfsHeKX1PHFGWNfwn+HBAt44
0P64YY+U16WsY+89yyiy8wMQ6YUSaN7YopslTwdup6bL6GJUZ2qf01ubvmDUPyP5
xtygiGzbgaSvSd/jUyUyQF0vBENwfS2nyaEBRiCzILsWE6CBdKVGtXQU0R56gtbK
N3AvWfLVUHZGcKp+ZwU9FqWrLNehi5+/bbGYHoEibhLh2hsasfbawnlL3xWxMAnL
bJBv3b3twxUZgCAn+MR3m5A9iMd26pxQZOiRqyHWXyKOpDZUgtaZI7/K1F1y4iG3
hL7ji2/CvfhViGNW0LEALNqTKvf4KRqsX/beNU4M+Z9k79F+LKwSpqpihXbcrTpM
sancNNUk2UXDV0UZXmeKsGHyulX/7tBIN6pXSkvBKc08WYQcJtC6IrQwl+5UcR30
M+D8InuVQMVHnXMI4QUGf2Eb6mTIoaJqtewKZX82c6fQ/0utn4148mHu6MQjl4Z3
kDq78zWS7KXrgcDtotFXSSAUh/MegXj4QdJj03Pqg0XcuRcSHjAJhYSb+K6qBWDk
QpKAom4MjC9MdesL/chGzcxlpqw2UpnX2GaLdDkDbOQzObGXmUGQ74SDLBCQA5bq
okxUXLHbIJObI7ZI8J/QmBbZQwCB/dgzVg2LQoPmr9RgQ5eUOPMRqG10ctKXPrHw
m8rLWr9bl6tIWr65YeBdvkwHikeZtnGKGV7r1gai7mLMqx/ESjc6xXeZSCQAJUqT
77MRIRgJq8XM5d4u0bNvbgmfPOTGfNK1Qhu8Mn20Xi1RPab3ets3bXhBgAx55SVz
vcnEOZ0UYLUM4YS4yMwmg2bGHxbX4J97NDf6YoOFhgmmChkrGptKPHhTpd/D0jmi
wJRdCV2D0z9zpRKahspfKiXA695w6SHj2KqPvq6fXyv5JZDRIXM0aTzFzBrgHiom
8prdHF7V6ZmNZQyvarCMKcgnOkh9fyJ5icy4xr0GdX9F1A7f3m8DiT1tNOegdCty
pmlFq2KQNjVozu2CfW80lo/3txuf4sdomuXYQQULXhfDyCVqMdWXthGk0mspGxjW
GqvFNR/pxFF2GNMZtPJaXGOCXy1hVOCKyO41aqQTWmZmPW3urixSLgAcWzSj5hR5
hsK7qDl+/p8a5w7IAKPqUoTcZgxrqqeUo2YWEFR2NhjEn6+IHaPQc5Y/pdFjy5GC
EzsD6pkdFINhhqTfXvbSRShTiWNfiPxfL6yvbaZwI05CK43Ukf6Sbi/5aq4u6dnc
T9DJIEeckz+ly27CHfAbZapd4gQVjnue5P6Qm/BnczWeiYMFJqC04BIR1WLvOnXj
dnPaAUfx1lCd6WKba6cXfYt7G59Ff4xjLLkewAIMr2hItMIuiENUWyUS/0j0f0uW
381Jibcs6ZV1zvNrhhUCuVHmlXKRjbcb25CeWS9gidXxEJkRQ2b99UH025XLjha2
tIxGtnq9EgIoK3QJHTm9hNZfXTu5KmFrTsXKZm/U6dsFtPAwCkAhGBiyVlECvgo8
OuidXuiClAliKt/JBx0XwdNcwkypE+4Ntq2BG5KtG7HfkshtW4fiOpzKwxabrNtB
jOm+2YjnPuKESxeAJldFlTdJSqLIwjDny2mXXmMks+iZxtX+8OMT9yQgFaFTlzZj
T/0pWiHYVUccT6V+30o9ExkjjEMCaMlWrQrZjCt4nd6KPhUshry0OhFfgwSs/mSd
cg6mXZM4U3Vjs32Tq5zJrodzyk3DcvKpA3WIl9OZKNMD7QhB3iYcaJQPQ0KexRZu
fVa9nYgCX451dv+yTrX1cmjAaTEi/DGIc1GB7fMBGNmOO4njmwVWIhgTwGCrrTpf
lZVSCeL+6noZUogUckPyDT1uYnRS+O7Ord0NN0lb0OQTNaVSRbVUy5vc6olrP35E
x3gtxSW2TkUk1/1vsov9y2wvF5RgFruiCNAgBVdvDobJTl35n74njvOdsxATllSx
/BSs+C5+K74QUfmJKksZLJ9nVyVAum+V5ipLz9XwKwY7QzgOfFWkjSSVXrRELZtn
F0DvM8MICNzrCfBtzT2lOSlPr+gK9r4MZgfogpBfJmIqYgAALZTXGTcTTeYoiYwK
1CYlaMUjbnF9K0ehGnza4k4Mk2p7fbipiRUbGE5ZYlx+C3NcZjyOAiZPg2SlPpEU
STHZVnhN8eIig3uzlOxihOH/IsaipaQVgf0a1b1j7pYuMBPSWHZU+QYNRaqM/HPr
Se6lbrXV2/GIiQcr8I079xL9WTYkfA6+5gcJzpehMkERKP5TFN0foKltaW2ZIiyr
mDCe0iH/Fp74em3HKDBp+JLeFngCpnNlex4Oie8mlMOEq3BH2GRNrtkD51/I9rSj
6soPLxakqZdnSKzR9z8QPZP8IyFxa1MI/S9yBO51F0qJwkfOn9HxswXuKg4LUAXm
DLd+f5EQzHoiEDKuF1xDLKJbUV09tqWjb6ggIxkLUfZLE1lkjsX5l9Sx5yQLw240
IykW0h+ZEereGuX4hN0cHC62Y9pNfAM9PnNMz+i3Y7n/ZHuh8SUu7xV42Pt0qh0X
rXm6ScE5LGczXQ8puAOQiH7lf1bKPezsFfc4nL89eu7Azzz2jYVpOP4nvUJIxNim
ot7pUUtVFH5GpuJ5WOHLUQbCqPsRaQzXwTsDvdfiPWL0L6yf7gADOAW7aK43Tj53
Vu+8BCyPoujgF2Im2+X+lvm2DBI5nqGo7FIAZ3FeILy3j3CsNGtj3D3Z8RRZGTh1
FVNfIz0RmQLLfrMyUIZC1EGG6e+BX91c6fzLRnDmrlO7cLiwSm7v/+GQklbm3LMW
k/aIx4K8QzklAmgN3ege/yyYk9h8NTZeno9NAkU9nsaHdnrGr0DrWefKJJd+yaxg
b665eKhUzKhVaG+f0IUtdeNZKtLeAEdL7eaYQryZXRSoZV1XB5g1qzxohv846KWW
Bo80Rf9JAAUKCXMP2O6zKZStgg8KftTDuB6xcJbUzpqPwd+Hy9mpG0D3uGuQK2oE
JCDNeR1auDjhQXRbyR8Q+PQX8FBEc8UX4Cq7t+2hjv/XIWXHPRWu5C4fEFjPYhDT
ozC+WuFV6bmDPauigMT4LRbDJD3HW5h6mv3hxxalvnOtj9/kmh5oidBcGYwPrsht
YLdVP3HTWs3WDU2CILeJsLAjH+IBIlnK9+evciFYbhRMCHzIn+3oyT9oSa2OMio+
66p8ysFtCL1fNacuqB2e+tBke51aFF3G0Q8enpsW8SFiPdZzWMOxZ7yEUjhTvHjw
/lS7CL3ZzK3Io9cBlgjPTxL6WBHEn/QQYug4KRhQB6z4JQV+i960ZnIJABdezZ2d
8H4MdZpMpJSzTHOTycbjQk14nZO9mugFCRLzx9K3/95Clgkd1ZrQNU6k/Umk/4H/
xZ8DKtj57ttVhDvVOGIthrnty5AXV1NZi3q/DiBEgmjQsEnkcom2vjF9TDMhEmDn
tLZp2OjhGzWTHJswCnrsJD0YVsMWR8WvaUKV4fagTxYqonSRH5Tuz5HD3xB5Qzbi
q9WJzXN1WbBvmduoVVf81Ule7cb8wicCaywmE3rQpi310PLkMBGykuStKGpjT197
PWmeXu6uxtCKgrXZTyA6RhLx9rNBDaQFIv0v3zkW9WV45nOs7cn+9voeGd+/8W2V
/d+WLxnzfEMumoHKfvIzklgZHCmW0u5P4Yj7SQoGXFuc1v9GAysNM4ogP2lFHTRx
YZ87thrJENLVtgL/LlBb91AEqu6w3cGJe2LUsi/8VTZbI4Ue9D1IY6amEi0cKCC6
edyme6/eSOAGm46MgNzcDO6jn8h87Q2cHmfOX1i4wH3SM23jriSE+wJ+BeUUr+R0
wnzboJ3ICuNIchS9crVw88Ql3sifGVM3SQiiMY8pJqZhE9Pun6foHzA26bO8z9uX
qyh92k6/+8lC5gkSLeFDR9pfXNIqsbtGrniLMMSaWQeXju/jongZ4ZUJ8pv5tYtP
5uTzycNxdDsTFiQxZSy6Q4f1opEC9/OchP0SqV27Q0sEvqJDZf8bCCXvhBelF/bm
j2pZsMWha8vUqK+yRqX4tBXyNwNu74E5mCIVoCY/8+XFoC2mJXl3my4zVDOA1skl
ViZONgjDKwxk28imFbMAMftc8qpNvWRksq6bPfCY5BAt4IIWRr/svclu7+IJeerr
YsfWRaf+sDGqZx9bJ8pacGEmAkBNxg30AVs6mHhw0m+mf7/Gl4Ve1efqOwqlIG5F
AXW0/W9/n/wrVCtBiGyKvsMkNoLvEj/jht/kbYtv58+ITatX/Issb/gfIAeTQOWC
/eEE34Qr8Q103HrQ/RyyZZu3+AoKpajsUSD5LWDborkOvtJypF2Bg1GfcnbWCGK+
BYgcZKylzu6j+VeKtqmTuG9uymfRoe2dW1oFTopNSWyWMpjJtiuqdm509dLCd3pD
Pla5cl3SwDeTcpDVpJ7naKSB/jlxQ4M5amNLXzQu564zU1DdBTk/KhWXXt1OB8/H
ju/r0SzdCFAcz9/vgGM3EtbQe/UMg/BhW+5ZOcIDrt0OMOMWKqE9gTvio41JdGEK
LZikKNzd98GciR5tacDLDbhyBZECjANVYwz/QFj1J5fBT9BE9mkuf//sDOj/YQIg
oF+DNyLa6RN6BYxwFjs0H/AjsnQB7P+EgfDimFntmbalZ+nA2S9I+Pcma3rhNX10
tGAKvP5+6BygR8zn05+wBFD0Rc3PK8VI8IreCLNmwqZNCjrXGHFfJ9UeUzUulKHE
4uUZQ+4zt/g1P7gqENehmaa4B2GQE6jJ6McJAYWSttq4W9UR6HlMuMYhzEzgBJcW
yW7ya9BVWMEoATS4Az2TC+C1hiDuZyyXHNPT6eCyh5E4/wdO304fEYDKFZia6atU
/k9rxcMX2+RpMKabUrpYqVr5wUDCz7rMQ57V+oBIYr1ngo+p3ydeRr116xI9tTjC
ry+vRCgXl2EOgL3YMvlSxj2DLKj38R7wIBQlyuMpLkDD+asJmUauQ+yHl/e/8hv/
N0S3mJpCOj35gyKO2tRgL8kh9IPqFeM5580YSy3UK9OrG4cAIWLqgrmE3L0xEijm
5YGdk/+dQ3b3c+BeJEpvP+bT/jtGevKGWsYRxjAzdV3axtQP8Jf1v9O0nVJOKrDI
CASSPnOKgp+Xh/3QKg4Joo7rFdxuCMkyprMzj8JwPwX+XkeTeSwwibEDHodqmym1
awkA9iIuOtmFgVaLftSpCeLh7oyrruNN2KPnytyqAGFzEwkDdOAvmKbnvrIpPoyT
P/iD756Htt6p461wcBT3yknVue3qwIuu8rVXINRSZKqs5guNbFkE9Sai18rTlaG/
keKyQXjSnGXXd+6+WwYtNPT3ZZCpJyqJlql1SxL847OfeKC1ty+r5sFxUTlZ3d0T
HcYADte0gLeDTUZOLYShJjSJaTDCaeLT7VpAI/j2XrV2xXwR5iDZBoqbxlOHc0dk
G8VI0L7ccjjJfipmfDYi9GiN5gsTKF94+P3A+nKr9J/5fgEcUyB1295Gof1guLAE
ozx5BZfupX06kbu+ML6tJeYcUjobQjc0oaI0jGcFTVT1WmTMbodOR+mUqwVpuWiF
pCKJqSobIW2UqkQm+mpKNG72G9ZeLw7Yy5O+f/H9fJE5/dM6HQqPTbDIjWuxlokP
c0GWW518k92TKyNlSckA7obtk5fP6Sf6yceIibGljMfVmUWps+t0Gv+V1417/AW8
mioChdYvZYm72VnYD1fIbg6FzJCesc/pgOJ+2ZlHwsCnjWKm28ZsX19dmjB4PNy5
2I76yumPokSaRUwJeYpOHPY64OjKLNnMtK5FgEcfEseVCLmcisaqtveS0zVmjVrm
D2mkdYjtDvnuKR9mW8fh54B6JQ6lTNQqwG1l64SXOoAjAJ1QzaeHLc8Qh/vG5VwG
gt7RnaCYbD8f8hgenaUw85CrNz+ed+74XAfjJWLrjqFLQyHUxbC6V+zelvI+xdDy
60zVF8cl9S/IGi8L5fVIQf/ifFCbOlIaViNTvqn080H0U9J9qVXw1d+S+u09PpXf
00G0Nwyj78pQa/P8X5+sDbHnKdQXnPFIZzSSZ15Mhr+QclqIMvegltGk8n/BtmYK
iZEhxn9r0g451P+yWWphbrpiB0jLaoSJ2kwA+XwPVuodrVHYh775LOHRhdXKxVBy
IegnCoWGgdoA5UZZF6BZzrunMB+u0oAN/zxuFrMIHIudFdeiSM57ue8130WrlH9N
P9ygM9Dcr+a/4xmjaCsikrnuCPgYlTEJQ9SxX9TuiskSvrKLxJVJPeGzcT74CFiP
MPzdKfMbLsVB8Aj6Kn7DG/ce37Ojzomu9EqLCZa1LmHR351xJpVu/d2HAnmnIvI/
quvDGfi8TitwckweyitkTMp4X30GWWxn26nA7ZqsGbDm7VcchGr3pZjESIHi1B82
ClAh57+Bn1mwkr41Wpv6qsBz2LJinZphhcUoLYdskEJCBQNDnQ/GlzdGJGH+4s0k
/OquZQGz02/2/YDHDklRyKqc6WOg5RWJHY9pGIVc7DqGdKdokAFH09oUhlZYGMs9
WERvY/i61PbLLK+MEJ/t1bMCKsFNmezPgc/+CptcTynvth/AJnEVrpQU6x7SRnt6
Q6s6p51a1z4nL0Jj5bVBKKVcxc2YJ9lzY9hPYc3qKYOrImqZlwfnbnXD2kdbiGIu
AEGrpG2Ek3lqfwRIr+3/wilX7D7bjCavqDVT9KfoOOZgZ3hxfYgN7A/nEU0/f2pF
OCdc6PORGY5kKhXAvEegZIApF5UhIuN4VbI6aqRXw/D28UbH44bElFYFWuUnGSeT
PzjKpCs5D5eLhubz2M5nVMt/jQKwKtewyuKY9hM7fQ4icaDKCaiWiG8Wh7N9zKnL
fnHKfsvpWL8CTfro0riXgDSHMCzXTNsZ6yHeeRmGfupTmxHAdUr7chlbM5Sm4scT
kAI9UowjKsfd2v6+/0ATPyug92DbJmaijBw6AMNxRfiF6wsLB13Y6claUvcb1eqt
DZVy066/ss1q8hVCBHg1T346wav10IMNfHSgGsShZTYwELQwlZDwPCaR9tMbEKza
c8/DG+JEbo3Qqxiz8dE33lVtouQl1W5W5nFeGy8JoodxW37jUOrbPNap5TeRMhdH
sjnOFF0aQ6cWowI1n23BpKpO18Iyp/u5WLqmg416w4UCz3yQ4LA+uzednBVCA/6+
c5cGxU4QL1mt83NdMZazjrXZFc0sLF3IZPT4lJkOS2K/t8TLI3NIbfK89hlhdZWK
kLZXqpGjtAePchar587k/D8kWD359c7R/40jqm1EN2lVrQCvIUJP9bU/tGwAteoG
9I7ov/bJUg93NuC2I4JyhI/OJ26SLvTL1LPsLJGjpP2s3xMPDGJ9sCTkhZQZwbHP
XfyRs7FW+Lrx8BbSIrIQ/5CtTZH/TI8//8B4lRest/hl1XdWjqrAcqN7aG9LcOlB
21y0x3ShamwHEdgWCFON6O+rLJVwCgEzmOPpu+YKD4V0NosxSesETz4fNVCjrGj2
blzDTAouNS8njIxADuZVQlUoB9TN899j1/FVe16vAHl9spVrZ20O6AumEbHKbkjY
zNcnW0BHaMCt97dXietLgH9WUNSJQrqnSYtrZFMw+ICR8JGI7/abAmEqJz7SCFbU
NGAs2whE4AL96VL+fE0QwjZsMBAS8YzAAKXQ/bkY/bf8eEE6Fa8ilQQCvywgCsrb
gP4fqjQfkWGoUms4Ge02fN0Cf7VmefeQrSrSIC+adRw0BRHpy6lGEXmk6EPTY/ej
Br/K2/sIX5mriEyInZwo2OrOzzMBJf2hXI/gKoC9JrSKPIpvAvxpozpqaVcuSNvd
FKJ16NLcHr6qnQXOd70FyZnO6cJyqvPdfm8y8hpAcVLiVhcOyT5EBx3RRKNpgmUa
FFIv00rVknvC4k0JZ9uC8yQSRuvo6v2uE1C+9KpYG2oFLRkVICYS7roqrGC5Arz5
ANqYga074NFNY6kGhxTe56uUwdixm7uCMgq8hueFfe7R2jZP1QEbSRHdkwP7dSCb
CV6rwV45ZfJUeqOksy8z2znHhZrP9jqgDY/7amW4fGO3DNyr36g1AU3aDZw58S96
UXVgt0m0BpB4zXcvC5R6Do+DJB+w90Imi6o46TlpCcBz4Ib58ypK4b4ZjBZy4tU/
4JltR1sIVZGqqgW/wdihxQy4XaS7BSdJbPYvG5b8YIpzLKNlkGQiy9185ITDNxCQ
t4DdnRgL55jpNDjRf+PVpRaqIAeHFBB7nwUb6SPCJSGvp9dxhqEu0zdufHVcHHS1
pRm0WjcHfyRvjla+6xIMKm7ioWi9ZnX+iAgiIRZBUVOIq8krrajBoC3bsKVVKnnR
u90ZbRz5bCDmvJD6d1iReGLUW9PkAr2I1e/7Y+Fm4dZ/PHp3PRAzOM0qL4vqf5Cl
gVVI5m4URgQUk2QqKusS6/fu55NH/IuWd3VxNLfHPoPfeR/6VEY5VFH0sIYX3YW5
Xc/qBby73lgHL+uOu/6Lm6/R06tdxJf+w8ENPOFXG2iUSW+0ctFLC1xmJbm+HrtN
TtpJ2KJ1rds4EaGGnkq9Vf6oSK8WkSIdHjhzyib3ee6l5HZenYc4UVXdju52IK+v
RWthVUbGEj4tJyqhs8iaiAQBJKPHN/kkl9zjMl/fGbFj+qWiAuRvsymejCW/m+12
PrgLyKOGHpfWFzzR8v6IbRav0mUsG4viFNYfwQx6XotXp1hIiK8LawSSbU7f8eBK
dfY7j3jQ/tGbz1gWJQ/BEpkpGJGawTqOnYqIpilPmKmv+rT4WWxRQHEBqvZAdyYw
r4+eulZtaQI7B2s4BG1WR1AEDViLOosB4Jt1q1F5b8ELEkE8cgJL0DF4N8hbBDIV
IFU5jLh8nhbByVwyeT5gUnViYIiRUIVHKPeHtTGCoiVz6GolsgP7EyvVrxmelXwC
pAdQQmQcj3oNx3CobXMn5tkMynl3QbCW1PflMUB4lF3tup15ODKErHBc8/miVycv
huE1peH6A7dnB+QvZx4WxWkiy1sels/VeG3urFwnyRw0iC3Gw6ReN6EV6TR4v2On
DKRv3RNqt3Zp/UwHcMTv2HrLJtrG/0fN6mj1eD9UyfY46Fbh2yWHpa54VYx1/OBY
fZNbSo4rc4PvaQ1U24GOxt509FBiwpdAVJIf5k4zDxkcTYfhyaHc/PdmokmzUDV1
9T9dRHCG5y9ycT2GXgkprNDdwa6igdgr1+VdYnKGsxS++R4evKQ1sT/XE/8BI6wS
bYEauHgabq8h9JyipQO34/+KMSWozsJdvT2OzkEo+R3b/Tu7EkeOIgaMZsl7BtVi
RE+PxLKQ0pI65S8sZCHmAbh9NV1gP0GRbBlFfrHh5Zlgm8eX3g6VlxUYDuf6VOEX
JLtm8mS0jtIvSdbSB6yhZAiTnxyo0AzrDIpTcrzXNZ9Kf4mo66+PAYbapEVq2tqu
tiR7T4XsFNnRwpy5WBdp14LWWFkozgrjUWYpj9bVnEMRzNt/M+SOIY3PVoJ7nlea
NqQDs9FZpBiyxgoDzRbWLSW43hcjmHH3Ublm0fLJ8l13sqvXtslfqtg4fa3qgNrj
prS4WWYrtJ/gBPzX9ifK5e6X443rsW0Mhjuj+BuZQxdSseg1l0ksqg2lHfX3kiBc
IdYQjpQF5Yp/OucaBQ16vpJPELJhwB45jxwII+cFDcvPTk3kBJqPuKtNZ6qu3bEe
oFne7SICsB2gZcmoMapiC5m2vInRHBAJpVqXujv4jZO69RRROD5k+HJHtcuLDZzq
IcXaZbzFIt3RAn/dNbW3mWE7xc5EnfPnH8FJ5DPbMlCFmClJerwqRq5Qo4KwG890
F4CcH8EU/fkF3D80+EUEASH1fZcYErTcNSa0F8STuWCw/MaM6vCzvEkY7Y8eG8rp
KuAiH37DRv/mz6hJTuHvCWXdhyKOmwOSkKlTgpcNVlUM9yP9DwEEINCktYZRWVTT
4/RnHjz+HxnlJd9JhWR+hPvQ/24qJdsPV6ru4VEbYmvTjS1aaZNaOzicUKwpUtBZ
Xq25y+wciwMR8vef7KpAa69Xjm0g3EaJw6ECSOsFTBhPl4qvdNuKtPaTV6BEu9Sg
yFQNUeo3jsoNrJFvXmur3TntTibFahQR2srDHTMudMIp4XJjZsV1sF+LjzLechSu
MQZQHSObUgr+i/nXz6fZbG/w5fJ3NLDrQdljwvuV2ABOY8X+yNn1pQ91cWGBBFor
PUwWEfN/uVAAHYpMqhG6LoShMaJ351REP3SWu85vLD9oMuzFG0xjo2wW8P88BRGZ
l4keKrGlxXnCRAP9P6kO4ngAYkD8nTzI6fZ41LXd0IdDk0lduoo+N6S+U8cj6feB
SdWzHOSP3a9pp5GrooSS4UcsJLio3JObP7JuekvNaXoT6N7xnw7XgfktZsxpuGfY
pN8jRhzLwlftTxzsK05/mCGLakOq1T76tCDaZGVgF2vKRkY5HmwH+7t9F7cHo/a5
0HmjHCZiVFLGb4cwfYN+4ioxjFk2I8KfqU0n1KnS7dsaLc9rRLtxrea14d2o+jq5
Nh+SR6ct0CfT5CWW31fy/fi92JZHFF449fRLIynZNuraLgRZxGDbaypy9gEXEeWF
QtUd11wmIRcpml/BcPGulWwWdn4n96+7YKTaovNFCI1Oj54S2nFYdBmnk+ZpctiE
sGdOCRKp59YhQA0Mh7a7fop0yzW/xeXggcF+5eRyoP9+ItwZAjS/cnHmiircxCL9
T8GA9qURxdXGZvKoSHRmb2FBnydYdPC5O7W1g/BBTRxSoKrbqkoLt54r96N2lIyy
/gbj/hZ/7QSgft98ehlW3TG+S+03JK1jVk1pTRl9l4Xzj2bM25J9TOtCyhDauorF
8xl1W/94vLKXQd+bdBFsjaFoPrtpRFnQ4npWs359lVvA9AHVkjN1niv3ZDNeHqX5
zO0TWGbzCXL4D5to3llW+ElUXAl97Bekmyuc8XzeeMd0popwtn3VSoamujx8+5xG
rTajxJAphlLSUY3YhdbCGPxSczSi/xhM6tKEuT4Fnhs2vAgzwD1bPnIzB2LuC4Bf
FUOJpmX/R+xK7zBUdm3npcP0up52JAtW24GL9imdISUeQcXzcYYKvUt2LZMAujnr
EDMeJl0gNNFGsdWzPEjq+Rl0djXxd2Q8pWPZoFoKOCGf0GWrsnHfz9S87cDkuQcL
KAy8VYJERKA/1wfrHXm55AIK1uZU8/0/U1J2/fqcxMNxQEFocsTst6INA9dCRtlT
kUiDCrD8jLXQwLe9QuUsMjdobmAgWmKkitro3/6iuES82v/g7I9Dt8qPH4S1NyhW
OlUFQp+HwzVjXJ+K62LH9WEt7xU9thwGDqMfVS9TMXonzswLut1gCAgAlaNCqeSk
g94pd7PJ1hAQNJbQdzxw2Rw5aznzO8RTmA3jzAPO009zkEN3tLIGLq+oXz2iTKgn
V9i0Q6r7CFOZAWOlPMhnM0cHlYGawVz+0gjGmHLM4I/76wL1isHI6FY0RetlPnLE
zn9KT1Eo0WRTdanT9pUtVboJuBnbytxpF0jgWapMD5GU0GhEIEDcL7743XXwkHOL
KnSDFX6SA2l/Z5ESSfd7X3CAcc7nwAq/Iw7zshOkjgRCuHSDQPieORMtegJt2o0w
v195alGjJbGjvk33XnEPOaKkkCcYLtvw8VVC0Hn5T48sNGWQZ0OIcO3B9Qt7PExq
0gN9/iWLTTedziMrL0wl68ena7yc+pGWfEv7e7v6e8CpF1gObsyImhH7tl+WvHB2
Tqexx8sQwhsOytd0b2okDazzhc3LUC64Iy6McoK+UfN/CAvJA7QtkNNTL7bhR+lL
vb+/2EWkx20caanTGk5KpUZFNx9PzHDPOEi0mNWgTggP+cHlwtBz4i0k7ZSNkClu
vQWX9RAHNjhYbj5nozAxkbsBLeWtOy/8Zihhg3a8CQiAnAIVuERPPxx0/cLr8Ps3
E3MGrrPR+7mW4idZ6fBCudErt9t7+Be1SBMm5YAjUa8PCs/Fq6SmX252zQNeOuqK
k9to/IVgcKyvTiYhMiz/3Shh4pfO5F3dNXA9V3luHL8yWcfuex/80rbfNNA1gwqU
CZfv1Fy+0sPFXzpsTEvoxRUaL+jlDPuUewmTPtIHSUGBsJJxdD57uZD9PzjtMlyQ
kvkBwhp+8eJa9w6WC9qFS2lDH9QE41PnG4i+BOIDocmEeS1RSvQ/vLy1iiv6U/QK
Gg/SkGA5Xr7iQUDjMxkIm5V8juLfp5gjgUtILiW8F2WvLNdQaiTeq/bU7iITmAqO
q3AEgA8qt0f8dCM8SEvNnGBXTGWJGlP3w4n2BvakNZOkP8FfkPYIqzzOY+T+SVRB
79behQJTxtXi2X5O4wPA2NnFfJ6yzPh+eDSq524YQ7RZ1vl3eqrJ0szjeXCdqFMs
50GMMaqmVJmbH26si9RpFrxn9eh4WxpxSB0F8V9p1kUGhwOb/lv4GHGbvh1Nkl0p
vdUdxNUFSriNXxK6Iumkv8/O2e8JdyH72+Xb2dJfiwEMDus+6nISvtomJzERyiyC
DR/QuhFEJcQ8mX6BkjKyxtcg6+V/WmQ9w0CTbXS/Ugl/PljMBYFL9aLBoyfQxbbb
LBb7tKfrnESnAZ+Jn+u3z183P75vI7C57k9urJczUvfi2g58g3rDuqJHTqkonu3+
bqMOT/ir5ExowpVHV+N2ZT1Vt9/XMgui+ZNQ5H4mI8yADS+ZkOxlAa3tAk/Gqyjh
7z7gfN4D7mDdj1Lhf/jw6E8lY0opfp3si07xkAG+9+h6TNK+cw7ez7bn3HzEk44E
et0oYqPCk1dD8V0kT3PE3WDbIcTyBZ/BPZ3A6wPBqwLueejQhkS34WWGK38Cj7Pu
p2o59FJcunfs/MM6D6aTVbgxZk6zXHXD/WOaEUpLGK7OVxyhLYof6mLmxFr4KoKO
gDhok6apLs2BK2KgOS2welCs2h8o/4UraoJVcR5i+XZg4pdB2txmzqyFGnTxiC5c
nTJNFUxD+hjqjIHbeT6OZ1tXhiteVN5XINUD8c2rz2AqcJ/0/PuatG0SfOrFpm1F
O1JtWmnPsL+jwxI4RIVIFmJv7oGr/ZOuMCcopGjXalyqrALbojfpGKAzsAsMsUuB
ZprTiREqZrwsqDn2aqrANvvIQz0oy3DuB4+xPI/7RpgERat0U64izarsRwrB02O2
MmDLCqRXpuI8OW2o+4p75iGr9ToBOPf+jqIZPTCfmiT0tCScILffrqMPkR6+YoIL
F0e0x51eFEym3IV5Ntg99s9DHrWq/kFdyUT9IbN0Ylzb53iU5TNqTu2Cm9RQuMYG
4xC0Z6ogmMwgNT0eQjc0NY7dzrWdyoPpW0HvQvjfrKe43ocS3htYZ9wY0Httge6H
jPlWLXaoVEdrxLRrowMND+FaLC3UG/ioDqYWgWKXGXQ36Q8Hf3Of2T//j705q4E9
reIJDJpipa8r6QprS84mu3rtPNz2PXxx6BvLmE/QSdp5Df85pt9xbZLOJumZIRE/
Gk7Neq91uIY2a7DOftae14mOCEA8pPKsWTRaszDs25P2LlSFP+SSg7N4yefZCJur
VuNE9Y5SRpAoZWIsvGog+u4XghF1ApGiA2KdpzAhV+0XHPmPbbYxU5aaWb2NAHhB
6vnvPmTAgDvjq/1hweGanHhXwtQMdo6eUYDyqxTPIzDcVTfgC15uspvUJu97i/qx
1Lj+IgSIMVjTwqDMapq6YRmlO6OBwImev2w7Z2UoAvG2nRomyJs7nm1vAPP/b7/H
Rwk/43UKcDOPCmI7VIjuNzszuEO2TNNggH+4Gy5ZIWZnUEc2jnz5HmPSHy87k8Q7
mwDTT9pVj4tx1GVGlaR3+/TMGRWK14JCNea5vVY5HTitGzqCckuSX9onKAiGM2em
+ZB1aPo0/2L0M+IPPCOz2OK623kp4PH+K2Gdb1HTBu8Us8j3/QyCMV65d+qbMBwT
rhnmjkumfC94RjISaI3MHz46ftFDdqJ5APtOlmBGoZMqG/KnbZhp63hW0vgOJDeQ
YE+PFKaJ0fAbfAVE394m0fe+8iek/dsv9lnkuc3cEdx+RbKvOCjalFkBNgXTvLrt
VluK7DM2EA9hu7oF8KZPl3/UUTVgSqU+GD4oPzZxYkdHcNouGozkkUrIKt7MoPWk
xK3A4PeW3bspvmxSPbERRMv7zbmp0/Nlr3BaUKFlnMrWLVLkYA+JUcTBy2bO9zVh
Ow3jmn+ovRxcfPun8Ccvj0a+t2xZ4D4wCjOSZozIf7N06MgiBEVT3ZAX76ZCAUXi
eQ6p0SmLvI26KeStKpYTL3ztupPfUikl/0mq0w+noFcN1MqbCOGOUjnWU38J/nua
J5GxWUM3uoULBxPSW8LIq8CrjL0R5rFJBMiOO3/+xly+ofML/tsUtHp//xHHkKJn
WBTWIx9sZpzpknm2lT2T5EQdIKcpDLxbSIEvSDNk8ETkJh0+2+zBnjLlv983zsgB
Ugig/kRvnWnH150O93iyYo89MpRrrcL797DHp6P7VOFfYTeGU3e8D3ga/bCg18SM
LvSBeJ7rTrET2Hxufx33qtl84u4RS9HY4+ERC1cVsTJvqhK/ud59MZiogpddBKEf
i9iM0k0DyL9AmQgm3PZi7sQVNYc8Mb5KDkuBqQITiEM7HAZtWDADEq+Jw0SAYei0
9Os9v/HZ0fjsENHKbLWrajByFUuzXXObPGG5QpWcB3hNAv61i5C5yeb03WtlQpl8
GpI0hgOAiIR4fIq6YL+DshMy12DLeBvgYkrv4N5ozjxaYFROACNcCqq10ekdUMqS
xStiZFIYa5v4Jd8u58rpdwZvYTKbz0PDI9TwFURnp3KSdvaj1MkKtdBh4/Jv/QoV
O5zR+rr5aquQzC3hHF8NHQHqECsAUMjBIjPUYU/LIgSh8EXr7tgPukhJbc18erGQ
B8cghfFCqXoJtmQE6rrHPloFjJEpo/AUYVz3cs8PvjeFon4KUffRjAEx+MDu1Cbk
+YZ27s+PQZ72hB27W09ChcfFriTLCwjuaAmUa9MyDbuj1ORokNLJghIJkv0jfVds
xpXGBqutIXN/wFYClCI8He0Q7n5EjRipJXWtFGCU6O/QWLNQCDuN0ps8OsDr+3p1
DhVejXpUJAkzihBlG07WHe1ccxE9zuNzHTkYxueJP6ftxwSUDD9EnYkq0fl8iEIq
eh1nCjTvlRt9IpD2Bu1nfCrHhzf6FLBPC3jcECHQwaG9E2CX6KTYhpzpz/isgWNw
dF84xm5aIRL4z1AoDdGxoU417SjiGZlzhQABkdNIURlpOgSCAOZnDrMR7ugvhGYW
ab8puOr3aTR1P9Ga5qjiD0+Z13ULDk7Lp7IFZAhHECQKtzPsm9ZcXNX/8fip7Hpt
+kO0ZNXuzBUgrJraeEYNJTGWDSVmoE5wgJNiZO63uID46xGy83qe0vdvzB6B/LHI
iAdOhU8BJBcCAdmKXnCp8laDskdzXYKOj0rP5ZuNaNG+b5SinnVaOiZl5TlywgGA
yWreExh2X/umr01tNTQbEmLHDBTSdyB/QIDQ5yTOgA2rC+P1z1w8x+WvIJwdYPz1
kq4k3M41a2vZDcyMp/rhrTzEqMFBYrtcKGXorgcUhNHHmSETqetkCJ8GKRclcXN+
OgAZw5HtS2OFArKacvBT3rQ/uRehKOApmIV/x+wXRlKz2QeGglL4XPGuwvnET3sm
C7TPR6IpE+BHc+FBlLemKSACRMIX5vpEbIsS6NWlH43I7+g28ECPOfD6kI4Qum35
nx2ACF4BQFK1kc5b0pkXCJ6DmXvyfXaP33KH/wuh6PgoSoE0y5IYKhBvoqfHpqMM
fqtBMcVfrZWLLXpIx5uaYm8ztSGr3dAhugV+EVPqoZGMnxtbQqJjkfQy808YEMTL
5na6MLHe1Ab9krqlmomPJdWSfi+06mo1pC+MFa/uDqGzu7QQzi4R9ZMFOdowE0II
bdPAm9dWDZN1MZRJptoaUue5SVlm6qh7lZmMH4MnvSv2QUbBV9ejZCCHigtwdUpP
2NG4G28JLCg83nk/9Hm75QqVwrIaAt+sgjHNuaIrp0HSqfXjAOYX7eUNZwVPsciA
jkfnzDwOGtFIHGhjopcU6vZqv8j1LqsVuAMgHODXQoTsQpTFy9aXpb4DKHB7IR3+
5ImCgP2HZ1Fa5HefB9DoNA1a1q1UqDYQxOwV6tlVuWsrNO8X7PAb7oz7oCUc7nRG
GGEJJGOO/m3RcfOHzQND0kwrpaJmepunI/AvPa86H2Z9khha5Gbl5XZWyAUnMP7g
qnGWKl473wCFuH93jNVyIYxnILSsnqrygSlVCWmYWlAktmIDdyLeCXYbyfko8hUW
yh9YYCHW8CfqKl35Yo2uyND8IIqtzuU4hMFsJmjZogMROgR/8rBls3cV7Y+IkuXa
HvqmuyyoMFd/Abtpu9gN7qIGh+sIaEN3T7zyCmD4LnNtAzp2rRh4efQqfrRXtcJr
bS3uJVMLVhselGzYTinxtpefveu4cMiHH3zosrBBr3iEiXnf49j+2ArAAD8/RoEP
sKc1TNtukqbh8jKTo6nWNcEZKdddeq5b8U8W44ytYUtJyIqfQI/s8CADy5Ebpq/y
XstdY7Xg+e4hCCCdiWxL7Hjhv9uXJWr8QIrxY2XCt3SHiz6fUpHJw2iixiX0zCTN
swggLMdmBM3bsj5GCAKYWd1yyNspnQltegxznPtcxszFUBWoMinbZo9At3inRAmT
2c9IktP5nV6TjIqIZatORPM+11bzaaKgKuAA7XBWKpHJz6+boH1a5DLabyI6yOlb
lC7lr29Cl4Jis2F7t56EW0nnN1WjDFFEHwr5NKmLgRlXCZtGDGH9MiT15aRG5oVc
7VpkCIDHOs2LON01xNhtBK0jSBeveTZu8GgxJ3/7/4UkQ9zd9VjNptdr/4qt9olM
Tlj8cdgUhJLIDZnrcYvINLxc85VzXrrNLRWtuT52Qi3mlNy0BUtPzLgFEFLok/0x
HL4JjZUeTYGYIF85ueQ2/RiI0cyKbsTzJOzpxm1/Z1SvYUc1HoGAb2fhZqpk5N/V
FAmc/M7UcCsUkSd8ynXBn0JNU+THH3JJOmFfUpvpZDQxQRzGfCwmG9i7sF3Nxzcd
lqsa88pFeBwd8mwRf2m24bxND4n4+EXPyk/sejgP+pIPzD9QeqotRBuUubvWbhrJ
hWsS0HYNQLBURraJv93dhuGVnXTNdAftpPoMnI6bITZG6XduH6DHZIMUwsrpsAeC
DRVIfmy3l+zMPR2Rjd2U+Fs3gAvCOomqhRt22QfqqIxvp1NZDgHbovMEg64yW7W/
70RB7W2tllphMtihDsuopx9JFTSZDJLi/3M2UIW2d8lBO/jKVNc1cuQiW7BKXSse
kT0ydXzdYKwqMDMyvIlbzZ/MXpmj9fJYDhgHDTSnc/IxUTGNCkRHfYEQv4LqYrIR
AG0umw/4HvwmlQYY2iuJWBhxT4g8zL0AWlF4slKFJo8V81OSAonxEWm+0SKTPMzJ
m05Rn8EqE6v4OIbLrvtCWUH20I1q1W9pPRGor+vIDgFG9cNuFuwPlPQcItwF5VlI
Q667kib5wQJLva1rRJHwwTP7K+UwsIhiRux8aUG57zHb5qbhyLGIAJu5+ai6HqiL
gbJ7cQUb/Z/vbjMsyDWNNB60gsYavFNfq8I6kIoLeX4SxH3FGu5ve+WbLLJ/L3Al
m/UEGyffpL/rL7YgvMJ1t1N4HFRAYOyLRQsmjI8SFkPsfc4YwgS180As0NY1OGHw
eJKtnWD/OpHSELhHRunESNb9IZ4F/WwSECNPtTG2nwntDMtrE0ZmQdwYNkXHH8GO
poRiuvSdygT6mDIaPY3hxHspufy8TPE4ZSQSlnNsIvPeSZTaBLgh5x5bcvAZp9Y/
kgE/L8QZEaXKpsNKss1SJb37PVDqzjc3IGq+4D8acvrOivJWQw7Ovl+FT/ZuabaG
oQHdI9cwPzfvOLzOp8kK0Gu+JUyOOQhThkGw2XjlcUwANuK+tPqAr2MM0uA+tIQc
ZEe/MHT4ileISrRIFhfKD4YrRmE8BlxBJv220nrFME1BqdAjTYyermC8O7yJqZ8V
fkjvCMk9Dw1jKs7wgXC3uEY9z5PH3uE/4e3R37OpuYHZhWpKxDEm/AP/2JzMzSIQ
vScthJNFBWAHIdu23MNrqB+pj1H8qvHys4mDCJwgItVrGpCoOqsc+/BANE8ZYu2E
gyerjyB3oQWIqIZP53sVFDuKzO4Xe8HQcR0x0X3QyNV7r7He8yu9bU8SDEuauUYp
plbH4N7iJTFpXSHYUskugVkpizjDIuNeLRl+BgVuu6ZBar3vGawKW3GNyDP8mg1A
63ak9/HP/w3md8bK0xAF29GkrMNE+ARPuUQYdvN/J5f9ffkvTd3zKOWEPjDLl6I8
671A3JRGtXfdoV5Reo6cmCg7AcQ6zhsrlMUPryyYmqSgJVUhbkLzTMxROZG2d51D
2mqkwt2c2DuDs+dlXI6kI+/ncMclXKV8e5TJWp/fEVf9CJwtQ4EGktxdP7/NvRJZ
AXqlWgi5Y/GAN0ozjgM3sJs/xzztPDaJcLwplM8fZLUzpi2oYSV1gD9wQ+DUgjz8
nD2sM4hrrx2T6BnGru1d2EypwUEuKpWlEp43NQ/sXz8Cvhr36dAUckEwo3465kcT
dP6RYS5loS/fXYVzyvKeRG0HiPmw/3KkYN5vedJ/UWlYi0MaYNSVBxZwLjNRLxXO
MYJsqFVdzOKeZTEaYDruOjmuRK0nMz2qtqCnMpdUXAcAgqz/JwWumAQFdebEarfK
dYT92F7ia9GY9bIfKn8Uey2mu2gGbMIU3+g2apqEdckVnU20U009HabB5k1IPGNP
fyA1t2Dd2KJxJbga1TAFg0dYbMp7vkE/SyXmcX3dONrGInYs9Gok9l0acL4+twjX
SD9MTT0+KdmX1zNPs0pea/PFhUpZaTh6CF3REj2EKa05obdQ+sdPs+kB3DWXLrW5
zE2ce84z49qMhpsIk2LfGmugoaf4qFWkkrqvkDsd6rUh7iFV8k5IHHMQCh0vDPzO
YelaILKjZEzlK5XBAzD/sXZvlziYpzhznGglkeFRbesjscPguG7j7I/RcpQ6BEV+
VJXBTfnnY6sifQwZeRA+knk1l/z5/0CP9FQrNcJGtruHzTTrhnY2dVWqMDFc4KL0
6nRr8k+t57L1/wbw/LQVFmcla3pa3RCJlm372Vjh2AQVBpqCMEJ2aDkeqzMZREg4
YCvrB04hYJCzPZfP5b6MQxwO25Lp5Qs+hIrhNav+/6Pb4jScqSHBpMPMfq3neHAK
V8WXB/kJ6lrLIErUyhfwaKiibGecFEvNEScwNAHKqxclu9Z33ZFaTQWEId5alQ68
dZaGzDqMaW9bnSSIx+6hNFtfXwNyMDnUZog62LrXiUj3T5gzgHU7kOrXqSJ1NVK2
NhSMdzUHkitS/X7v33e52vkLICfKPf4EggOsqPOdyHqbDYPRf2UweiCam8AUACq3
TMWhIsbG3OdEXitSaVRuguU5e8waMWfj0+pbvwmP+jMNpufXNmnLaHP9/KSSPZut
gCp97ug64uWtVNwS5L1dKsZIhEKw/tSdyE97Z2+Tcv7bg/hiT7109U3Tc8bfkCzm
++jDfbTPDi9YM7UbhZ69gwLCYUSYiGS6suWr7WLum9ri3WwqczyhGeyblXnpKnL5
j6V8RCiqGKe+OJP7Qz0jUe48UZp8XrSW+ijipgHplajTez48phiBgAkdlhnirbcV
eraR4FfvsiMuabd+zTog+361s0slaDOm/FK8bjMMq0YQvol9glQYD+m1p6P/dH9W
jhzYDmOVU2cC3qyA+2Kx/fQ6ebuQ/yC3nbkVn+A3T+9i4K2RDRssB01z26Q0O8F2
88R/MsG08+mm2zwxfg40gFuF/Nt3KBb4FilNPjMC4fjsSzsF1hU5GKugLpjp/xI9
IqKK4Y2FEioTrxkzoC4mTdCHQsJfpDJQCP2NfcAL29VuLHADusUPDEP9oC2zsxT+
B+HowmLQdxK5CKEDCLVnGqJBhsWgouodRhq0wMHUtl5Uybj65xU6yFY9w5nn0hYZ
aRMdAA4L8tbeniJ0VlOL2kzNfpWT6Ssm/wTfyQuH7IM4yMQq0BNWW6wT3G854+0B
+UzHLoKmSYuqALb2Toi0mOqyP8DVIwg3YpV5KV+R8eFaXSAJSEyQjAWi8S5HCLvh
pT+pxPpywD1uOh8Bh7+s0zcrnn8+KikrsGQ0bf0MRAGIfJOFfrRap4gGI8fY30wk
kf5i5W2fOrPjm5xZDpWGOGg+Q0JRVAB087YPZUBUZboETQuuNWk7FK5yZh2dnjFu
tsyInGAOnWwXKFlKk1YDWZ9gw1SILe0azNpHWR5nhFBwq2siJNAsEVAYJUGxl/bN
N2tEAlOVrhaidZVcR6WjTXLC12e7lVChV1eMcQVggz8EKTknVqQzaxchT4i/Dzxm
mJnv/t3H1PubjY0PJWow+fGRPjK4VXLNk7Y4685CKbVQOKjWG9rrPSqqmWizm6XD
cMQEeuO7eKdWjoLfnzM8uOXKB46sLWrtvlQ7qu7siq7+arDH63+L/veInGT32KjJ
JMwRnkhK6ErYB+FcqDH0U6M7ukBLlXR0YOBkV4fQneHLD/8OKPZgj3RB2AX4TTnk
oCIszdre8sQUrsflbvKF2e+T8oi4Katck15dQ9CUVoEe7HUm/nZyAjD8kZ0aiHue
D1+D7YNm59WD6FALbEFsyf/CVCsaMgYYLekCfJoYe35MuoIacu08XJ+HbR0GRBKG
gPvAT87lJRZ6tBrnN7Hwj6Bu9BIypbWoTEfX6zntNt6yp2Z5Q/sjRMDcQz9Ki20Q
CBAC6dvAaodcmQjflFhEHgq8FTa8jBUHXcZn1F+9dhqUYKyQhRw3iZaEdbcBhx//
sYUciWT3ad0mFYstCJoqL2DZJDvv4qUZ8zaOZWL85F0Iqi/wdynkLNYxaQTNGZGR
i4AIxhutEJDcEQtJSTNQ+DvHYDSuwOfwD+qrxMLUnCMlf9CFz8JE6Ofd/TLxq1rh
9KsdtA5MAy2SpVeYErLKUkOa0ft3HThF1q1UtSgiT3/WjxCZIorAtJSstbHpySrE
0MW4xq1VtHc94bQq513ZsBddfNLcFilfWX1BmoafhLbb6bh2NuFpeoV2ubj+xUEH
6tQitD8911OX3fQ5vMkEGRvxkLcrTQYv3QeXD6n7559zRLF0voDgn9nOcoQJde0U
3SDF9tfVJ/DhILLj0mMbDAJHozxFzZ20KfQhBtV0DVmxwCtypd7/60FRT85nB/dO
SZrbzcZ4xfJB9YgNC2zHX/u8iHgtJ2X3PySNNPtq6oYIf0CzHH9zaO+tbybTPha1
XnuRvntSD/q34qRjrALMhvnPK7SUWM+KxQ+EO1D9IQqwaavqXX1+Dp4jEkF4g3sP
Mk05qWlfXj6gLuW6oaNVqzwbxEKnZhbhfgJQBdjhc2ZEP/EOpT5cTfvn5Sn5YSRu
DMl57zAFytJzSeVaQl2XEXblXu7KRtclokL+MVSXRpgBoZsS6pvZQqD9vgsrlOpO
8UewzS0Y2lTbH7hfh2VFJ8nnUTvAtLU+JPxkW1qDEyB1qS31hnDxLj4LQa79mnBU
2Mni2HWBs8cKkZ6julRZWtpB7EEkbyBuwNB1fjIbRVoyqLOywLPvAJizBmal1Pgh
oSNiL32FokEXjBHjQPdr4lEwCJUNIEjDG+82NLf7PgvlKFjwvq1M5A8RnYnEuNtT
DNhSwUeZFogeqquOMyuY9xg2ZrlR+Qwor6DePwKcc45Ij2sf7ZZISp7b+sbJQZVX
frCfBfD0m3MoGEQB2tN2HoaPLjhCljV1yoB0JHyGtOc8Hl7gVK9+BdCcauyMMdjf
aBOU8nG9Y5cH5bUr4NCwX8onkCnfuZGfFGg6r0qHUmCc8A7updYDOMkZ7vaLgGSe
gj9PgSWV9eTpRvaOct4qc2XkIcj9gAry01yQwo7rfGx/lE5+XgaWSYDx0dMZic8V
jgqdsgVFSkIX4rxXi8X6+g0kQjYNdE4wq0uGaON4w5972HkYLdTgdkOXoMAPPIXx
KnpRPQrDeRWAOZ0ssl0DW8CqGdhxi+mytluLvAUZwmleQXxv2fpHK0oKUK86aSkj
8zj/JXzjuUD82LBh2Dq7lQG8ERdP5nO8/3nOqtJIVP3CPGclpDtQ/KLUoI3wCKV2
Z269+yHkGKwFfkWKI1iPYKKAJMptzPYh5OIOPYyZWYk0BHk23CM7HLuQ5zmAMrVm
cqJ7uBnrnSyQZCtJhxF2SQIY0g2HQA/926pCnHAAVz9WdefMi3OKOP5mx4EM9ATk
NGlwBT6Hhe5xeDpBSeKYwmYDLv2NaLYlYHQA2ic8VDs6YmkyuFa0wmZahAYVnmnr
9QFWm9/IKC9s08WPSVXrsWhadxToxk5HmrkAEGiwi8QF4GtOhNwttlQMx7wvgBMq
ae2HBffsq3ch+9IKydw/ngJwE2vxL293uRLDKQPiqyax79zR37nXXS+NIEMgHVuq
Y9orHh8+bhWs5Qh4Fj+xQE1HTAHrlnCOyccW8gLq6TVATwLwUK9plQ783TuGXdla
M6HsqSJHusSaA9S/cznNSoUfLSR+pbMrmwjTrYF1u2OwsLT/zo5w77S1nijVggae
1GnTMvHwV9rktR2Tko7i2I3FLck+kA+JtlxjYtgb2GbSxX8AFYXpCa21lsCZN9Xj
DzxkQz+1qDUM0sweExoA66wqDrm3qJeQ9ywjemGicxriQtoEOuLA+sMHbgbGHqzR
jWOGXY7w4uZWJNvJMs73XAf4KrpfP9vgyiXJtmHC017vXF2J6IwL6aLezz233tDO
J70h2BKO6fSi4G89aR+UYnWL1Ls8+xE+UQMgWfrTBdcwFVz2LNoE9FKtPQ9dFt15
jUOeO4jdbhVgh39jQeqiSjFYGcBQpdfEYAYWRzVGZqXXvve7AlRSQxGhw2jWRLL/
tqwdBwzrtTj/Rqx0AJ/+DnTmxl1qZ20uHoFnJmCljpCuU6fQUPhN3Z78sTMsZxDS
Ys1xm69bjeJIJC0gWhbTsKwXZnT0deaBFeqwpwQ0FW9laXz4LJBSxde7qfi5s+UK
q0hBo2lay+RtBXmO17nxOdSqebJW4njZojNxlRAHLfDtd661ujp/jtyeHSmDefh+
/N8UjVjjLFgUlub61iCw5SSoQSSidcl0pAcL7Djn1G0g0zrV4LCM6GYcrqpGKPvg
LE/X9CtDSI4R/pwr5blH6HoJza3KlR3PMJUSNNvnwWG/1kKIfXOmqj1tXHb5BHFl
PT1d9BQ4dogLEbwWmb+4dnlfw2a4GgtA7tr//t7F8XMV9AR4DnucBoCIrMwfMviv
MlUQru27KWIclS3qqLpS0P7sF6cfJdpQOA2750YRrYc/Itl7a2mOtKciUTzVWwS2
hvKLT5VvJdRfKq9EfsrPbZ5G9oLsaYFMXJlkFGWTw/6Q+TpT6xN2Ig/H7lhbYbFO
JqBVG0DOvI4f8BKHdAUfwqqs0tOIseJiqTXvUEpyn4suwE+Z4Dulpij9ad5/bUfQ
Qo7Crq8ATRSdbmUbhWh6kyQ/9aSGug8N3xwTIprpasiS3akIrNo07Weu6anbiZU+
bU5+d9JaOg1Fd4UP9QMGdWSm34Sdg/XsPOeqs3hkcGLCzE8HVbSA813h+6tkoF3S
5LSl221p4vc7+7pG3C3hJ7hbCynHjJbEg4yTvuz+d/Qe4mud9BDmW/3wqlaQB5K1
+f+e4aJtnLiN5jEYC23fc4F8z74mAFufORJtoAy3MxwPibWcugJJvgc2ukYjEGvc
v669m4Ghxq37zdkEnyiOskvU6/6HV5ejxs/El/LrA0vWS80Z33zGjarTsDANcS4S
DO5WGxzYPlC3yQfSayqt+nOHiC9NFrGMK2eJFOAwu1GKwb8LdFFHBdD5R8aMsImu
1AiHAP1aw0ceNQVA5BpH6jSK8sqIgADU0a8HI5nGhhcvAOjiTkK38WFLQWCuvfVC
arkFEB2X38DOn34oWCybVF0+l/pbGX3P62v3uyuMReh5kUEEdvi3GJrElFA93i/2
DhpmihNLELkm64/LLBbyRguydsMta07pO53H2zugp+dvpxhwdWPC6og0ng0uQZ19
KkEQr4vHchgh/7Ige/xZwAMQx9tgPtbjSovZkN1hHJx215nOZsmskDsbkPDCiZyL
wBb9pT7p0T4SiHEkVNbzQXE+ZD1FUQ2Khu/LO3nbJKxXWzS6IWnwxbHRJ0+WHhBP
MdvTFt5965awr0uBjHcd6hFslgwGGIqcDnKddhs2raObnZGWMD0emX5Ea1ElJKCq
9BcUdMOMEjMUNzLmfg9cEqhBbUQK/yXajQ5573ByK/J/dyLHG0uSjsliTH2s+N1l
wABrnpOj7pzt7htsIHRkJLUeHE4wSIepWFr9btEgF2yDeUD7JO9hkvPlpP6g5eyw
1/o6ULhm73mB9fIsAnWV2RWXlVEvsz/48EXv5KyW2ZlapFI07BHgULfE/pfBpGUG
xn2o1fPJMuyW9VoXJBejf3KMXCLfC8KLFusiG+XGAY4CrO/G/YJdUc61ZzA1eQVH
mdwqBVCABL0BJ5uczPA9rO9uKhCtKC8fUoFed+jwhIp0w13St8RvuMtzyd8QnTkb
uIgHimy6SCrcVu/FD9aTFjCxKDq4zzk9v+XBfkZVR0auS3wNCMRacmPWQlvFLoxG
Ea57RhZ6XjlbF9oifmXe984RcDp7rWxZjqXXeadV20LUoVG8R5CbCklUrawbxsRp
ZSiJlPNyXg9FEtoHN73QPH38dR0kHBfSafv5HePB+LpzRCWpU3DhEpaTpHUFXDL2
w54H11yoSC12HcytdUR54m3ZwHTVLpp39l8OhmaFiITuLCss+GNM/PlYLvwSebjQ
4viR1ZtbhGmR6iKOXKH32y8PY5yJtuG6gG8Xwc/prfjbVmTlZQiL5UdVtOkz2Gd4
hXwOGoF4eJonbdEWgw4OyaQE0BEElijdExNTpbkemucbbtZzUYM8P0i+/AiuFhuc
WtWL88QXoQsi5NUEkZ85Xmc4aG0Mzonnd6qzwreoH6ond1Bdu3cZ/o4HhiL9AqkS
eJ4sKGS+Qm8h2ViaIRZ4ZTBu3d4oPhSXAaypcC7xK425U3+QGqvZIl6BpEmA92nU
+I/OADeIn+sAAcI0nHTuKr60B5TSsGCYiNaKcMyLKti7PNG8a/anG58nX59m5Xrh
sMpD0P4bmq85r//BWNVAG2F/WgxGe68xBbrwkjoL0g3nN6HJQ0rYy0D8F9qMvF3a
uWXuxVmrPnTzmtZX5BAGzT14lovthfo8fzOf14K/D5CyEySFATAB8zQus7wtWJ7R
IHf+LIIiWCrwbVkTux9U/+iM3LbO+Ba/8YNAEQpd4s23GPPKM5jrsc8UAtyz+iTG
0ZD3ush/eVe/P8AWDvBvp01OE6Mu7TlswzNOyvZEaFwp9cR+dFUjhhQJopuWLtNW
O+miCkomMdPe0aiMG7mbN9TklqIqD21lqjkEnHBYw7oe2fHbDyv4+WC2uF6rL7yp
W6hvEzT9IsiuO/uMPNZKOwvhRYt/CsudCjxQcZzwKbSCmlAWY6MaTvzOPOmMegIE
B32tJopYNbL2UCwLIQNlOEeV5wFln4aytdT39cQuK2SuSXuH0TcuMyLx4GWh8iQI
7Bk8FNyHiKxYlQj5t/YGNhkMqIshtAbolymAuCa8reCmZmBwNBkR34VvjlKCmYoL
k89Af6sZ2r0TmenCzQrrHj9BwntJO0bX3Wzi7nJa6oXU47hhb5PERJoJWf4PlPdL
oZXWbNdX0NNm3O21eZGeFDYfM1Orj5rjmLT1Z6WrhJ7UU4R8aQ7lqZEyiQeN04Pb
WTZhy+Z1d8voMaLXZuzC5qTJ0U5oDb2lJR97FslHUSVx9fPx8/oFOVTja+m3BWbO
XlPx9BX80qjlT0cbWtvSD82/VXM38keUnKqjufpuAWr1ZtZPVGJpVylmhnGAICAN
7qBgUJ0TVEs7Xhw2UmuA8sB8l/4nzqVuf2+iloae+YB8vujtCkhIB1KBKfXYXNbD
xLx4ReSgWF/U5YfPKupRHG4EAfSv4qUJBG0uzT2ICnGfqwJwMSMKmgzREYvwRBF/
4Y/LXNCAKZ4qRUfgSlDdncPn+KypUTUJ1ejqKny0cYVVCBvqdafhEUXoKkBTQMdr
xBhpfoYdUYKpC2yqu0SzrpHOGoNwMxq18Bb/NgCH6TaCJ4WD6aOuPy+HE4wqEZGU
vZQunw7EknEHz4tTajnTKxKyAErsWm5SlLSBw6M3XxFZ8v+f+Mhcqk2GWjwdAEQ+
qp5O2FLURMvXduAdNXMOamW9gST1FC3/VnmCBVW3FEEqKjV+a+148PiQOiVxIot8
TUJ1tKPhQ7v/K3XeYQSx5ERHxR2dJ2dVUyFKiHC410kBWfHmSQhWl7GlkJAF6fkT
T6gbOPM4eL9RU43tmZbXUERFGYBwYu+roQO90X+bzUCrumaQV4O2IOust381g468
WtFUjCnnbEZCNjezvQYaidblmxSOD5Q5Lk7iem24NYoO2IYGtqoYTtqPbjGy8/dt
Lm+l/VOVRRqi8OB/WVLk5CLUpu2ym8LWTSiE8xlMtGH3l1U+TIKL4a+OIeUjH7aZ
D8goS04ahcbyMnx1pxtSf+Owz+4Z1dw0QdsdQ/eOLE69+DOKQ26Zcut+DiTwTD2r
jNSL6jOh3Lfy75EnjlnNUdebsDbI9Uzw/A/FlRTrt2g0TVEaWYlv4Ecl65OEC61g
yfjxNXcQGHgilanAdT6s0JLOUlOKx55i54CD1acdFeESKYdtwXorkxBu9a6Zy36Y
snDIH8g9jeAJyicI02JB8EziQTDg8JnJLwMCDIGOF0P9cPt1Vqrxy0yud7JcNv06
HBIWWJJL8FRTNdFd1vR96AkF77fdw+GhVIkj+/Oisb4R49OszUQKxcRVApvIiTP7
7pkwnWoGRyNrXhaMJBXe+LAltLu75ggGKwXeoaxgrdRRH8aEoxOdR1/u6knnhaMO
pi8MzdTTb2HW8mmC2Ntc6zq6uQgNtoNnvOS2ARhQn5HyR4mMDdM+2ov95V4g/8Z6
FF1irWCZInYrctQ1rUqXlTdVLJaz6A2z77jWp9JHwiIuLyzjVbAPMRtsIl4Er1ME
4KQA0VemOkWAK6sa2N1rUyufrL7mn2/gwy8bXfVR2roVT++gAmA56qE3jml7aBOd
SCny0ge/8Uewiw5eStblSxNJoi1WvKeUAod6vXFy/qmUd0ANIjy8GKaCKKyaX1si
o+eFdqO9hyQQWH9wZIAUk8TlTiIbx7QSVnE1JEyWkJi/+cZnmLywgut42nZ4SvwB
1vfZ01m6wKz7ZjJizAl1l+2jg8jFFHqSD6AwT8XeGqsc1GAIhVhnB2UBo45kHKR9
IHfReVSI4k3h55Dz8J/KenSiETtFDI3spZNXmcyDL4BKRsXFImG4D/R8LAbVv8EP
FZWdMnJuKaiHPA75rcgHYeuAx8vUsInHnd+bAHiXobDo+hdFjjOs5xvMZUCho7cK
tA2KLEppK+UfJA1jZDWR5ccdy1t36PNhfz8C87Wd7AbBjJX6BHXpZtgaW+rAG3B9
k+OQh9b18lVUE6llOEpBg0FjDR7kaG12Kkve0wqedMUreTSgdQ4nT8LSAxWvzMy8
YRAxkwtZm0kleDZdTzZ8Tn6JsHn+l0qMjy3In9/PRAVkPH0dJA4ry2F3q6Gc8AYO
tk9JK6PaSTSBFItHDiVyu/2GhhQsy9en+ted5zdxxo4JUu3pvRTd4YiRVmfRilpg
7llPJpPmCl19Ers2IeG1AfviyHqLc3tB5q27KWq589tNxdd5PVvITxsDxffznBf7
LTs+ZffvPzxIxRev6hU/3GiaH6XgvCsJ3m+OBMW8gR6qVovDBV0/edJpwJbdUHJ7
yX0iKwdkysB8mpVIGc6pzzqZMaDIoJE7IkhS9c1q2ncXJUnL7if3zJbLqTp5031D
ELPQKOsCanx3716bebSFMJ8F0CFYflh0TeUwSvNuzcq0VSgpkvpOgsa3Bcwkjww0
U0H9weX3d/tzKyk/af6c2CcT8o12jNTFdFBl6R1AQ6F3tBx9Fwu9JNjAcxKjP4Al
WnJEtSnv932HO7rsqtehNRe+8S70FuCfRDD5TAGuJUJLQrlesMrzyHxyyoTlhdlI
lKPd1rOvvK0UeUTw9mQWxjLdPiWvGpAF5vSYJUaGtT5Ko/qL9h3g53dW6rzfQU4n
GKq90iiNDZMQPRLPazQsX8Xoua6YVG4nefzHwGJXa9v5KpjBV9Bjt7B3vly9Tp16
RT65LzpgOe+/hdL2IztQ+9EZPieDqIZuRyZz4vWfljJ/rz+jccGMlbeBcVAeOa4U
uvhfUiXdcRBiBnXr8ny3tChSw1qBapa0xXh29Fb6ns1Qrpk547U2NEYwV4istXdm
4yn05chcFArrYmWMpKUvtVVTmbs1iw8yYITghUb2daBDrXrd0Ujcz3KG4GV08Ffk
rlY/V2OzeEmTYVUfEnsM0aPyAlyPDWFHW7Z1l2wTg99oPE7+Z5Ri3+xyk6l8QT1F
83tdrfBMf4YJWknRcxZ+tP6MPwhGPSBMuUmLk8dS8gtRSm8JGifiKiDg2jHdRAO6
XxCxidTy9TNLsTOgKpOa8vXQEgxFbva5JKCQkCE0+yAuhXLqZFb4LRGBf19lmvZf
LKIppBwGExQGYyatM5jm5jg/2NzfXY9+DWnMXPJ7VNAWhvAFAPa7UDYS1XRLQC9+
FYwjnXDE1Sf7z45+kp0j8+T/FkQvrsCFesJpaexb73e/SIkh+EwmHrRTs7q+yl1x
1AHoXnr/vbjkjCvP0Q/+je4/t1PqHwfOpklKo9Cw9eC5zLj4r3m9x4v4wbW9VLbq
VaGr5Zz+o3cMwsV+xtzcv2El/cvn8acjdu7Dvi6zHiT4rQAxRCmrUx4qO5mTj64A
HGJJlOhM90oky30JmYrS9M2BEF4fL2iRnsA7URASZue0aP8SZcSjyO+w8oqONHdX
2gxxpkz4Ec9zOPrnE56cvFW03fabZZNq1PhyuI8EmpVLdTRCIKumfR3gRtr5XdPh
MrocGyI6bl3bMocVsgcWGJbd4Pp/865ai6UEbbsBHDX9oEA4QZktS5EsIUKAjNc8
razAVxDTWOGdKFGprRFRM/7XcikJZC6H5/qAcj7aSY9+dA3z1pETLCZ+iNsQx8J7
TKiNXFDxVof2yU6TIRheZXZ8sEj1HPhu+pj4YT1tFff0fZWN6uROnMT2Aty55QPo
0N0EvcatLL5XyjgLFceG/4Bzh7De0Wm49Z/POVIgQ19mA7ab+vJzIuN6AiF3K1CH
gfcqpHTVScJPQ7IowrHdmtGo2CjVhb7As8Mp2juLlrZ3/EvxZCRa6GfCm5vtbf8v
cCBXBPXv5CzOu98Npx2B1vNQuWAhxeD2zUrz+fwVdwuReP819Gu/c0uKYft1icAL
uCC0xpHsmC8D711N03PLlPwcRFZ4Afc2GfaZLfJHjH5ogdm0YErd8t/lRvTheepS
LLo1yI7D3uFDC5UnZ4wIAm/HnqoCxrFDTmlta8awtvFuYX4nuELV1T62bbu3zop+
FuMRNcepW+rboygSBYkEeKLhNroGJoWyTheSwzo/8XT5W1Ese6Bibib6ZcZ9tAWk
o4RU1Re3oJlV6TPdbhAhvFG2xMZP38pi446Q71wO5GkiFs2QrcnRIbxXtSzQvxFA
7Hlyk6WLvRxkh2Th/K8P+6ct4IV7LIZ1NRY1w+EP8pOPG57nnddv9u6T4+j65zfv
LCZ1rrad2zEzN8zJB/5OZsV0i7KDEg0xfKM4vUx4/44LOJcMb0eCq2sbj3L4lrI6
/Z1kmIFbrbPzwFOlH/057dv74iyD1lJpz4ume+XrgDVWNuG2Tud8NRJEekqjh5Wd
V3bJ6dSE125xzbvjqIBApfdrHIGTRHTiLY29tcGQlzzQ5QEI8KAYytMmKcDn9JuT
Lf1VSjH19X5aTu5ljVcMHZbAy2qCUFZ/FfJZSy8gIWl0k7sHoKRa1B/QSyiHRbcL
iE4PWM3EaT3FxA5WchfPUIB5WPJDysS431H88dGWDePk5CKB78tUlFUu9/SD3Ow8
0JbXV/akBO1G2e+xzR+bV0tDj74Gp913sWmDPTj949MQD4NG/wjn4S85Qss9W7ZG
bVAzXTEpT/F8V2iAMIUHjbixOKupJhpyzYL8kMyRTD1T2ixA56gYGqqvHVNhsD8r
Kgr3ZyAE7MkjIg/awgcxcwzlngj4fzQZhS/5xSzpAE3/AaNW7UTWy/hgwZooor3L
vCJqfK/oLlAJL5locbq2RyY+ybFAkzGKl6Hr5LXGBHf7ViXuoRrZpLBpVKmNVk7n
bA7atM7oLORyfWNaft+M/S5muETy5HGIttQkoGXTEsMgx1eXkXkKMfnbSjTC2+5J
YYjepBLnvySl0dzfEoS6iQe6TCTP4LCgMgDmEKaK2TvSJqzdQQ6QD4T7wlZEbQhE
1Iz0IYiVXAgya4iqGME5yMR++IXajjqGnMvyA+xDjFGDzQg+0YMufYgC9x2uAS/z
eP/LWe4xqdzo2wkKcgyiP+xoxpqoloV6dwY5slOT4PICTrdXxaNfXfDKlzRWF7+j
cO/6UzmHBH+XnGy5QXzAKTvpt5BrJyA+bXCd9rifRQAYaaJ2+z5HNxJFGNr6NKy7
SwYTJaPZuX7ymn41OFpTpSQNw08cNcqZCkNXWKw4gQvRJM6IuPa8hKKi0tdBfgTb
scucJ2LbOBsv6kvbpva90D37DxGv8EJ+7JjPe/rS4hWn3KNEnBPX1B3a1n0MRf+H
mX2Xb93qxKGIaXJucaKiA8ta94PbfI9eSC5wg4I8YObzZWHh+POZZWAmRbsKSwfc
aZmxVE95hhoZTRIVMpXZoAoGNZzeKWoCjgPKyVnZZjQ67QqiRaVPgvTLl+7zxL3P
mTvDPVBwNS8x+RgkUqygLSDIbek8dSgliaoH2oAMfcTKHPTM+YlNZ2uudGK2vO2T
TI3i/XMiGSPYdG8+a6FIyJdtPRY/ST84QurXBoSsJgtOEGt0Wju3A3mbBtMGWBSy
gg43/6G9R/flCqd3Vek6S/A/jhL0nUQask5WTkpCSlgYiDlSCx15u0qRIzdGzVJK
v/z/BvMI1Pw+8btzpc0jqNOFhq8qAepiS2FeQm3lSkMRyrucQ+dcECge3afxSl4B
VJMycw86AAMDMgYlXOGiOwqIjHChuPbg14R428f7BzkyxC++KHTFqq/udVr5Qs37
N8w1sPMnLZGAS/B0BxvQtBhUaHf3EmOui7kVYJtgHi6fCtv87HFmOxrh/ePuLxBM
ujnBcjwL8T3HXwOXDLBetSAbGaqErJZMLknOhWpITIZ1vYT77TqbrBCM0OP1yYb2
FyiNMGLHE1Qz660a2B/YfQXsrIMtUaq0R5PIAqqMCCRhjHZ+5eAhKiDv0Rsc4SJt
jJ4YpWcBI7wn+WU/aGF0PajkXydVsQ2sva/upfBtS+g4zGgKrDxeJu4C7oGB0QOi
zNhYfkB/StifRLHDEWu+qoNZnhFetouTP9PI+67g07u4bUVfppoZ+V0Kpd0FP08h
DTfD9DuWfYBCxezLwnQgcJGRDQ6m5ctVXAi/Ayqe9ZDG6qp9TjjjHYUYpw0+EO7r
AYw8RJj5t4Ebuh5fLxpa4mZVszPnl9jPASc3T0MZxWCNY/hHtofDu6Ylst9Db+5Y
CmDyrgeevgxiWejvIcGlQEpt/mBrDv8t1vUrFTdTnAMAfS/VzIXyxvHS1TW4U3BF
YJACeEBfIcGsj9dvG7wF+CDb12cEVFHfgZAN7+zk+lPC4lcABNtpxQsj0fXZBeCy
n5/uyLEmls0p0EwJhv6qFSzO5t/HnlgBy6P4DB46eiSj609WT/vGBr4cFt9Fxhpx
cLpU9exYcyTRHaaK2pvJnVfE8zQlZnd9iVYROQJ6yYCD4R5bb5DFCkmBTwPIwHw2
l9B3CrTEY9MRG2Qj68XFoze4xD4ZdUlY7TDRr5sPYv5XoTpGh+soCjvxMzn0NCsA
KBl4e6O+2kkkb97oTW7uPnlESYo0+4JyFoIwXWCq2zQlVlYmrTnfsVeI5TVb7s/2
yXr3cEX8p03/fAsBhFXdBVhjC3bV6VPyCvzsB3iAmjwN8DdSNmWhjxpHZnAtWBm0
hQ0ntvr4Gt6DFzyJiw4MAyeflVziJmAiNKdOrZEF4towajLXhXJ0R1UVMW/gdy/N
01LwhPreqNxJK8I0XP1TTo1B6XxY6u/iKJvDDCIeSdy6p0XtuiNjt4Sry5taQ3Ul
3Pz0NjPsZ6+uhq3xLFt1uFZZBIn0rANPVquqc6OnKXJV11uLIbLZ750Zgmih/gon
f7gm0Wu+hjn0rquefKzeyHrHHmBd091FugCCawAZet28Eb+nUoNU0rBsOSrl/vuK
gX9aUihD3kyvBrZybRAxNg79lNxd8ivBrxvH0VkdHK8+AyoRYd6/QY8nKH9L3MPY
Io7+ZBgZQZxinStUnVEuYEQ5jhkC5h8TJ+3oV5jQ6ixIbUvOozVc7NQuCbpiV4ZW
ze7m0MWHaeRSRqGKh4BaOSOrgvkUrIBX0mA3qD+LLbTFY6jZ/Vi1oe4veR+GaB/+
q0OFKxe8FOylW538Z+Jylq0vNl0C3sfjU/NIN4lhO/TK2dtbKMwjIyNnCrFJPUUl
BdVhjZ5h2POErhmegpk1UgZLbCm6GzqwQTcOp4XviOGk6LF6de6Zbjqw/++FJ3l7
MQ+56AxdQFsa9Itf6w3LeCUSjOSWIfSkgH091pPj04QFgU1VcPC7NHx+VbpdcyWZ
fF/APYlpYIsWX/wLdLsohnG41i+yhdXjweCa/vO25yCWkuxHeHhspa+gPu67drsG
kaeW6u/mP9LZhLkWCzWN10qWaWci8UJZn59I8dXSuIub6qDoMho3j5MwGRtLACFJ
lkDEr7CBBA1HbXs6iZE+OZHb7XEhR2PwNpg2j9NcC828W5+e30ElXx5DmWRgiuV4
xY3zTfOSkVJwnBSx/exNG8spPsRM3rSoRetTK099zDuH9LeOm/CxqJ7LAsogOwPy
HVEngQS+ldWYTv9pWMso6sjM5rr9qQKanNaDS629tI9bimT/40m1WV9qI5DXRD2k
IsvpPzeW1Q4uLNmAviS9DW5p0jJAmi2uDbNaz9MTyBXrGgB09y1d1ay+Md82pLeT
TULofgyMOZa3t8b//ofUbibqycIEuX425n8YiQkrlDBy1KBJsqwPVOkUEb7r1aUf
eSS0DLov4nP3zco78zKaW0ChezIFCXOD2LovJvzMzGyxIydVHIRzRT9Cugx/y8NC
y1d/50DM+j7wBRugJyDxukbtvegdhJPTQd62g3GO3/TPscUhhvS1zVk+HzlLU8yO
wnDoHUdvkbIQOHLDr6GC2nzPX4pbZLNkNVhji8rjZWJDILnj3KlDu+/jblXCnzbr
VTdVziRs+fOZs5vRQNrEld5BFvfTlT0HlXcp7lDErmVQ8OJF5uBjCeuvRj8Iqqqw
bMmom/G3PthgRiZICSXqbZ0xJ/OG76kz4VmIetTXItE5Yv7LoqrNN5Y+qim3wPLD
3wTq97QgG/ZU+EBtmUdqtaHpfxwqTsxiuoqbMw6thteI8+kZix2CtKoljtI+1vy0
Db8rkYQi4J+lK9JDwR8r82PyzKcaGK2QweQCUQT6glJMGy6DcH7cqs/zY69vsufR
V7iu2C7BdA6yMT21Y+WMPyJqE3ZfPIHNbDY/Xuig6K6QYIgpLSPJZznWQaKsObQH
f2IWKBBf/avjCtLJUotk4H73lG27y821oNtsu2sFrkMErLc776a98Axrl7j/C91J
UxlfFWECQaW6yLxjvgyzTnbyYzvOJyBKpL5JUnj6grPeztQQwMO4ZJhDnXVqPlmW
uvpifL0AIeDqMA8Qm6+YUYDGsC114eGzavMGQsVlQfe6HIqcuSFfjwBdVBs/BXx4
5v49XEfOGoJCRazGzBt4de45ApO1fngR6fLtzVH3K4TUDpfUXa+yhd8MOJHNaciE
4tolpYbRwq7I8n+2dROlZOcHuE4+VuZuKDvb3byy1dWAnQ8tboOE9IVXDN3tCmU3
Q6aOFLawVhBPsFJH3buoFjduR/Jiho1JFQNF1wc8dIgJ3mVjZuRtrjOpopU5stJ5
0icRjDHgZvtB67qFCD+/JXIcG25fm3NLAPB/YylQ8WF9tcWo2DJBLSE8mKggqhl5
+5shfDUF75gWWUPEfteDZmB8XoJ1R7G/syVJq4qsoViGPd9B079JxKfAzA8kmQb4
YWTplutL1Zv7zd8QxE+vZoyeL+TCHO8JOjF9eTqxpPKaur9t3j/hDnkrBqIAunvp
6XyZhjq1i3wcRCyaTRwSb42M0ie3S1wLifhudah+k3pFh5VorQ3Bm/x9UQYEATed
x57/+PdWXt1UUomfzAtf+aKdxXqKMphFLTrS07s7Fe18jAavjMt2E5L7S9q60DNw
Cx+0bYqsTVuLsFl4wdfOmJ6v4mQz+jtT7OlwpmNo9s24wYXiR1nSNrY5xUZItnlG
dGsWrrE5+EQZ5PmY7hESJ3nKXigNcTqlLnK4vFf5t0rEs9s8ltOA6Fqvw7cTgXwH
IDo88VPY3Uall840ZyACKp7Gy1erH/GQlWYFD1T0RwgknEkEPaNHTNkCDicj28fV
kDTCLIrSsfvRk9uXGznLT+6OjngBJCyuyWBoPAR6Tu5XBpuQFTJMIRK6/taCGrBP
7ZZ94MKVP7PsqnMPD6nuYu/YgS/V9IcgfzyHfK8W/NbIp7BcKKSr+ZfiOqYTTdg9
IWy7MZe0IraaMeonrihexim/fePMovB+e6/J7x0EItUn1yOvpIrIldSVv+1tJhHc
a+bX561rb+LsTxKkvlGCFQQZOCEePzuDOLyPcbs+3Fd08xHqS7+WL2cx0VfToBaK
+zFRsAJnLhS/8rCyayewkMzj7odTmlqbP7MAqFOQhGs2TeHDMa1jEYn3LdPDI5TT
LF3812zx1RPz3+HPxHpPcL6S9yQsPcwwlA3o2rSoqMosimaiLAyXHd+OF4+fb3gc
wobcg44fqPXUgvBEGvkD18qIT9ZSnw32dnH/Pet+MStbQwUeoNWyTXBaG8d5NQk3
NEpsnnkVPwSVkrLPZj3qhTffWn51cfbUmGYhi9vDsf5SBUoCATtGFOL0F3SP8cCn
enKjcZE2PdBTDieYUNUaD2HrZ23wfAycAgtz0Pc5g9Eq5ag9+zNoXLiWK/OBEmGO
d73qMUUOS9H+YuEAoUT8X+/9UkXFpWJJ6Y7j4zC89+hDbDrF7zU/IPh4iAKQFslV
ZO1a3802/llH/cKtSHFk/+WHaPGieaOW9fviX3cIWXhWZiot5mvNWFMCH4Tr0McS
lkqNNHy1Y4pddXxEJEejzyavoBjkSjG0MaY4QKzKwLeppRNFfND8TjAlp20lU+nf
CGj+RQ/Tw0pgTWtkhWpEcVUxmouivo3p6lt0+eYMku93Ix2EZCEpbfuo9WWeNfTn
wTPhr9CNhntb5BIuLxLeulrxrgbAri0v+utMGdxa0/pT5R2HnLjz+UsVVNtJc3oa
/HlKFs2a4ORL2kHDrHfuRQwTf9mMnFyubC6KxFUoCmNw25Q+N8lE2uHPAqf5tNxM
RekzIKJj3LocTe71I1qvOeODJQpHK9Iryyn/DU9xKJeDOJQLLvg3dU54IWWnzahf
7J1+AzTEttwlGqizflhYevMt9kFMYzU9okgww4aYlW/vRvjUTSewiI0nKndnHn5J
gSivSCkLDQoeFjPDrjzNEpCRe0AXThZKqOACI1yM1h2OS+bWlf8oGTpmPw40DUG4
4zyzuj3+0r0ZCkOc7RwjN9Sze4bL9TK+zvS3M+NE21peS1qn4EQka02Ffm/ePdEj
g1pBqgCUSpVbuhl4J6trZKNboamWqmKgIz6jOcW2/9UaVOfHiKNgI6j/8dbyGESN
ENdUUy/wi1/l5JKdkFMYQ4aWERcWwG6zCPuLMca97qCjrG5mNHEonz19q4Ox+aye
wfHfo/BX3qD+R+2cBV8ABKQUyryhyjxvyzZPFrmBfHdiu8OZPq7/Mt3PrYj79PX1
KUnabnM/akXEbOgYiice5vwDMpx1cMceKdDGr81Ne2kOHn2HMAFmcWeVjIdfUj7X
ahyCMi/O1nMqaS4P/QsjAeKLGEL60hpVtzULBVxUbhLfah1Oep5j4euJqHvekh95
qdFDkppqVFP9M5Cv9KGz40RGnKxgLrmNr+Om9jYlaM9mf2ADLOCBxqJbihzXMY3z
6xVZifx9yMV8z593eR0kTskXk1BbC+S5fgGhqqosR6r67jkJ055CqjTMHZI9O0TP
zJNnyY4CTvqQhTjws0YNJlq5UAyFQI98ID09ZpKUe+6b2f4DTEzJ6QuKjM8XafJY
lcNt2IXYPUNwd2fpj016YV8+KIurylPKs/qJdFYmUnfIRTrSIn+/x+LB187dYFeZ
G85rezmt6fpbKwnZrFZxTc6NkQ0w3sKZdrVRtaD2tSamnzcKwj52xAUKR8S5hXlG
j/7n6My5keT5DvbaAeiswc18IwUj4QtP6vyCF79BPeEbcMpsHcqOJKe3PRlMY0Ma
yAgvsYD5IxjdyfsvqI+QyIaaS1jGfXuZ5YdEsQKYo1TY+UcXeYRdY6REuViT39cW
/Gv+fn5RTctPq0MizZ8yQXU0B/nkss93czJb480c9675DmSlDwZEq6QoxlnSjJEV
FhrPxvfXTSTVIJ2IdK3OUMNT72iyqgzOdvAJW8pKVNDqAcOo21i/cgIJ9cGG4jSW
RPBqpsna9UDJztGQAfW6qD4J/y4ODJ2C4wlM33BKouw+S3TDp3Pt3F80cJhcONZY
j/hZqe7SVgVaKMcc/co9dzH1hMp+XQ1uQrqRJqqFybOeRllfZgPZpmI7DcDZdEiI
6W+BJzkXIUScADN/dNUBdjE/VoFT9FCRP+30uw8uZnHPze5LA7BQo4ysPO9OTGhY
W5vfJN47OormyLvrA8so8sOg9KDY8DSkfpvy/XamsDl990394r38LfxFK7B7Pdfh
3/xzph5B6xMWVANn9CrFDdJZYmUN/mD03519K20vU2ACB+8BxuK1Uwxr5rN+I4jz
YoUHKFl5supyMRfGnYmmg8zvwpA76aMoDIVQjSO7KU6yew1bchRMFhoOPlKRxUNR
/UFDw3xVWKLZ5mU+neE4ki92+E2eGKmjrhx1wQhBr9GboO7vLI7x6qXDFn5Jl5oJ
MLzae6jEvyiVRN+R1ZttZOy+vAXixvJtJMNIFPBcxyBil8kqIbzV8FmF7WVTVrnb
CSgcUsL0p/P8pOtDBkLo4yLjaZdEyrmf3xcZuesFTSzePZrKxOg+NIH6IWK31COf
d4H6t+BNRLnBPwmob2wyqs97yARaakdDE3LzMPTYdzNU8CzvJX7SO5yZq1t9FDcQ
DIyD9/SlzLjc3DRsgB8BI544wDYF2GqTKR6krAlaESDI9ORjYiTcruKe6Lszh91F
KSLCJM6qntvuKOjVZA6zDmIpNqDzLHrtkb5SU7457/RzJailg9Nadi+aSvwBTFii
dvbujblHDTnkOSYbb+bVmySyPyUs0bzOtrGIhKmoLgmI07Qxdlh60s+wzmKtEZul
Hd3KFVrmiBrdLYG6neZ5ZMzP5KrieiyHX9BGODFlLqQRaML/s4Mlsyabe7okBi2J
nm3G/gW+O/AbLwOKT3GuzVB2y3tuzeUZc6JBHWoGwxPLos52or3ZhPDf+7Fiauit
2iPygre2YHqQe9zJsBnetqdhcxDgSz4K4CE4ae8+D6hiaHBbPfxuoNmCbdGQ7/G1
2OzkhYlsRwUOltsm3BvFyx4zgxfNKHbmpVxkRdILYRzdAsBOyEKCHGEujO/itxhP
LRBLsMOI4z2JM5Xtb833t+HKNOJSvDTKchyfw2iCJRhN6qmqgv8JrIpBmdINrHNl
nUNFIDhjOr2gmf7GBrY6qbkaM7ns4KUomdllNKWSQqEbxryZC2d+7X/yYVCs207k
N7LFSLqDPpTQmPwXVhMbo0jsV+PUezOrWhlg0e5zcAy9hFtBGLP2EZqb8r5bT/Bb
OI1r75/T5debKjf1poUfgsQvkaWHlRJvSAxHKB54vBmqbHuwcFJ9hn2B1OGNdVks
lVFFRpbK8xw2jn9EMbhyRHOXzu0YcsFrEp0xo5Kjq8/X1tFaq+qE0O3sBaOHQ+hv
9zFuIEnWeoBbfjfNG8hpaeHjewGiiMr4rMkP7ltWDsQhWjQj5Q5X7yhtMovcwbi+
ac5PEnUz0MKhEhg5e6YORFDduaG+5IEPd9I3W7os20SfKEAni5/e8E35MNNLVJru
EcQFaQydD8b4JPx5OgM7kF+c7xvp2IkgEsRV1nXqM+ql4ZEXC3lfIBLJU1woSLHN
xLaxLsprwvRoBbxnpqH10+oAH35IghVfjuUS92zZPZ7hHww3CNqYoYhziwPbIgw9
50FJE+v03izoi8l9KV0ipcsE4FfKyJtozxwvabId60J5dZS5n3YdOEQu/HwReQQy
wYw+gdYf5q5Nia4bMfwrzenJX9inuM/DZpvVee/35ibt0wDOgty384u7/THob0KC
vnlZuOIRi6/dvty+ibuTQAEkVNYFYdLyVnjLrPynOnkoQnz4XukcD1NR9jn3rzHm
+QqbSm+jhmjBFY+71VBmZ7RhAs28ikU6+0GgLujtX4eopzUglAabKKpjIg8OtYM6
cc6iyBxR53UGtPx9cEcGKgWRm2M1uymBmFLjJBrML2+9s/jT73k6JnWYKtg6IYe2
S+ZtqEj0PVKya08UcugRmsoj9P/Y4X+KIgBxKetclQVOKVM7W53DJ0DTAooGqBjZ
y9lOiVv8IHN3MMYy/3mziwjiiM5IZVG47TzL4ygrQos+cmujBWV+TICvqh3DJTBS
/+7TaeOS9ki8Pcw1cfUrxdiRWEeTkEyEpRkxgdQ3MdttEi5lwoM1/bLc9s09oDWC
nhb6taMGtWqiLKOU9hQlaLnau2dvbps0T9cSxVI6J0X6z+at8QFYEDQ34bSSGaKN
f4eaWt1HZp2GsojpqEnrKDxZOWj/XE54yLd5LaeLNYSzPRCTxmM+eXq16wGrWT2G
8c7nwCQ/Wv4fncMXjzhlk73ZwE/ybABIzTAKnVQYBsi8L08V/ot9dNAWjawnbJ2H
bfwzxXBQoj8gDPAtjjfhmF9/+kG9ETeebr2DV61wY0KCk3dkm4kuEY+GrYB1G8QX
ORhuL+Tg47iEFFUfTkd8wBk8TyaaAxl1Ca9vju3FsgKm2ucvJ81k+lSPGXwi2HpV
wyqPn8OCzUlpK8bG/eH/EmujBlvZztHgXrJjRJWLoz/ZeYtXGtbZxdrQLnr0lUqd
PCfRnnA9tXKLILAmwGLqgIwyHHWYJT1RlCxQmDONgU6dBchipZmxzvjEndXDJ0FI
Xrh9Xb5T9SMPzERM43tbuX+05OkvpAUN192R4rkoGb3IyBH5xbLNnB9Iu/DShJnr
QF1yQlSfYjUiO3GEnvKqXZkgrRrN99N+OfN3hHS8hAFQ6vobVnVwkOtWJMzANK0q
yAUd1wEfQihxFWEzw9RwHydGbcdmUzCweBXjL/X+bQ9Fb6t5t5I3KX1iiPK0qLXe
9NUeJEedr8hCaE/HMh7BlVuGUZKOi0E/RwtD9krcQK0NKeU1h4ENNNjVdPFX+LCh
KW+aURWFb6wMKLSVLUqegucwYXBQ96pPj/wmgwT4kVO4Srg7ngnNpPdEa8GiCgEj
DVtZYccQLfbignTrlQmSeEWgVzSeQW4rWNPb0d4AJlQwAgpyldQOvuTiCVNDms9j
OHOET4QrX4MzsE6h7dyuN+DnXkKqNQH4fJG5PdM7qQPmgSKqnECAyDzegdfH1Nkq
HDMB2LMdWNti+FnBUO3c8u3s3peogv7QFLQFdb9XfPezVJdbHsYkjZXe/lYd6vow
R6t9MkH25DTV8nE9Po9SQGkqZ4491783vLTS26JGJqYhdIma1noy57Qw+zSnWfrR
XOH55Obo3aIsxYzGYtCAjM+Y2Vb0nBQO3VYNUW56HhcqnwPmYEWMWmkZWlAz9e7W
fK10TY7XRHjfm6SgWhC1h7F6mruqt9QP3bqh1MWC+wnDDkrtQEkYS+GpIZsReK9w
HRFe6PzH68UQcCMTe+Axc6PiTGGvMz0NoHY5Hm1MM8v0c0WCMbo7EjP5sHJGfICv
RPEuycUZiVJxCY9kvVK1oK8FpwIf4Rvz2Su1o+5ngJOpZHgxYRlwfexUTwMHNyxC
nK/Rt6Oe136K1lHfC6En393ABNPJltk3POpoaGj28MyyXpOxKloeC+1ZbOTK5PY6
gbbXJvZqL/5wgWRbC4qcSKPu7CjiT2+pKGhiuXO9a6dh2RHh63014PFuJK6oXXUE
/X13ZsEGZ7KHIBPGkLOl9gignlVrCZHQMvqfUHJ+9ug66VxSmSbCM0HjowF23Uha
K73dWX61jXpNiEWt1J3bAlPQmunXGwT6o8YcB+pLpXaDQCyio6cOBzA5yZZmn5ia
fbY5aiipQivlvk2nesrJ0JDnznB/Vr+vn1RuHpf3mRlFUp9OjQrwwrcKU+wJLJrB
SiNB+vaJg3utpLspyffM58jBqJonbUBrDpMZMX4/wb5616ZhFyYqycY8iMT6DIKR
C11fy9QW4vyvCxsfGZnAVFy8Mp238bdzwJs9JIi+4hTACzrYL2N3gFNQ8XhNq7XQ
dGl2bVgQERbhMw0nTngGgeOaMgnzmLTGUOXKzo3XkqHchSdIVqq5k86sUosR6omG
ZRn3fTotGPJWw60N5xaPIUeTNlmwpdxUG/OEk1fLMs5EStWNDX4ajJ+J4WNefvwd
sPl+RKn65CLIsQyhQxRbNsU6VOJqLRCxXWiDBzOyoLd8tc7AXK9B/Vs3S1MxDG+3
6TdgvM6QlzEu/KCTZzXbqZCOyf7gSsWohcSpUAUgG+sVFMVDKsc8zFfmwDzNDbrp
3tFRSsIpoNnjWBkB2ZztgS62N23H83aXrbPzZFDyahLi5mzdTIbFwCmS1PvdjXM6
wSP5qqxRzON9jQnIt7f8qjxqT/iROoAIfQZthaOBPV5KVdxKLQX8IRojtC/4o5Oc
KnRpI11zpfgWcq6oM809H/VeRMSoSeUMBkV1Em4yTgTmjrFoV9JwE5cdDo4YINSU
6VT/JbQVBIOkvLGUUtH7+J9wpK3IjYGaXT4eL7B67JB+TnNn+U7hcKqd2HdOXUYw
Mie+7SYyu5ZY+U0JyUaaIAD758Wtsq4E3yR2Yw6wDOeiTkOSm7cIV6wqknfepNlV
pbw99JdtX1lEp1vEfQ8HgwTIBqclqjFAkh7TWau9D5nVyoe1BCFf2wRTHi2++ebg
6fAcgRBSiZsLg9Zub5doVSJH1i57OEgDMp25k29HHR9hXfZuITjwg7bI6fgjSym7
J1UmvG96PSpiP0ZXlJrT1ak1+dc3797bNyA+QWwohWrUAOhKr3NIiRGaZo2ReAnd
XB93Xpn+Mt1yKjofFMY6BJojasJ87UguHI44xtOHOIuPEVGZ2TzSsHgKYfMKVyZI
jmriWUDY3otMdBjNtAyUaXHZKjvKBw0iYam6B/MaHj95x7PN3M9m7uHPMl3d8t7f
6iooG8fD2WF7diOoVz5GUyYa+PVLg67VdijEElntRENV9AcTo+VqolDF+319f78s
udzxnjzpCc22Q/HC+heqYh1ft+nAh1KsItqsEsKGK6d02EmOAJxdf8LYEtXmUxXh
GrqKE3fZzQDvfpRFBUcNuOs0NEfRUmAKVvRNwmOxBMv16krZS/YVZxNH1FfoXsSN
4hAG28NmfuIF6JYzt//tFOC1Ap36lklqXe7xYr+5DBeMCWxA1hwbi2ih8CtOL3PW
YX/5Eu+CNwxVp5OB9Wwoa5MwqTelMN0i8E6CCcK7thgeEgOTWWJSw6Z8deHuNmZ+
pcZlBAZHb4CTHedUgyA1wS5rWzZ3GbVEYgjTYqJQzvi8cl+8Iyubrr0P1yyAOgZU
+htxcg3iEyqbrkLrFWtTcGCPasCv59uMCCqU47JqOV5+QPkTYn3iWXsO7PVospxd
SgHWTB1ipJ7WFttWc7dDLimftbnSYpw/riF4P3RhvC+YBylQ/cauJebTWH+2UCiG
DDfZJIouP6w24s+pe+0YNFlfaeq2L+aejCl8kSedDAg97tvYHAiOyEiQ/i3KAUI4
JuM13wzQeXvmXCV2TjPgc2IAWbbETgwMmwlvCNtijeKSSAPHdOSa2o+rpaF+aq4a
Ae2rvbkWqULpcD9K+Y17g3w1todESYM1OMYO0QSgbZTYOxCXX3nxammJkFddmiCZ
pbZkKdKlQ5GYBl11SfPwz8N2mFXwouxKDG9NeXItdiV4KEtsa4Ook1Pw+MJGa1Bl
z3HQ0lPsXqhuZ2g5bo5O6AgSnJZH+FK5XPWlJy5+r4eDY0/ujAaYjbBsMBCDO5Dw
djuiUN1JeuAOze2hxwRpfFoKbSvDOQPAGLU9aDh55Sb1weLk3l+xk/JyGesgnGiM
thNs0YPyACxaV/xrFKHipc4JHtKj+toEtqcdMUAQVEKUFhpRNbDb8pf4Y7E1pSMl
fh5/8+PHB9x2OkvUoW0Rv9Cl60iEDy9ZHWilRmG14XfK7+xsFWlxwA5tFGJLUHRS
H0jGCi/WStkmVVQYPos0XvkDa4ReeczwEH+x6mPBvOYknTS+/saJ6I+O4zrG/Jwx
M1WvpR+Td1YC+EciLpD/OPZLrA7bGMuUW2nhWcOxgRSjo/iDWh9x0GSOYpRjCgCL
ST6Dz52vyTLZZgmOY4CZP6T0RPb0HYjXtgWhTqqlbfSJ6dOCreeHlDBtqFp3eZGY
nM2i1gCqZW+rgic/mXyKOk1aGzbOwtVkhhfk+Wsepha8bdDuhUwd7WOA1k3B6I8j
8pGhr4jHWB3Dzf2R1OGDYXb7WgB88NRiF/YYyj+O2e4O31Tlgd6z1OZEPeefvrSi
WbxN20LyPDA+eSYnJsRrJvZq2HMl1FIR3uhRvL2Bs5GaPYdTO7aR1s2FrskLBtyF
Pq6k8VXCILdA+rsMsHUUZ38d+533JOQBm3kPdfGhJTqA1QJuB2JMZeeXEq1KJ9bb
KwYGnfXxASNO03hKyG4SBApPZVjdvPEQ+XPllmVOTidvdMmt8v+buPDvcGSnrGH2
ZVJlx1glNKBa1vOijouLaosp2PDekzgJq9OE3H4R8Fhb9viL+AK0Z11hPE/fqB/g
ooC/0LfSjVIpG8XUdw49aBZdFqgETUgrEL9exRMZxAuGF46+t3Pp0djWtM3AbM89
2bXoJ8TksZJxcT8suS9X9pEOrz1hvniCI0zwB21P7TnAkHnBfkSTIvjB81PfxQSY
e1/MQWndYSPuvt7GZG0YD9WTPN78HJOxgWoyIrzPHA5x+oMTQ3NZ+jCw0Nvj+but
TWdX8Pyg+/UUq/o2q9w4GlDHI62SykftO5Qinaie1IT7o6K8qeQOTNPJP8JTMEed
vy/Fj3d5McmglSR8kxnbPAhotI28PZEfCrjgsVwA4jpD27dYqi8E6SHAX4qN03H2
V57etQ2XCYN6uUDmC4kQKiNMC3be/xB6E+sQ2W0D5uXOC6cRC8AbZD6gYHqCHx/s
/4YmmKWTceTKMh8XB7Jmeq2nPtpCJZrXz8cUIC5S6sYMcGVNQlzJp7/H8k1BCzNq
HvMGp9fB7xFq8O6PAilL2/8xBNo8PpnL5gCEZL+sQ8g8IpvK6JyfOYyNNy42aplc
IFZm2bYYsswv3J51VsLT5Kxc4X6AXxD1W+dEcsaC2tKpIF2Pd06CgUmiHVpJPJk4
GgvVRraJ8+tL4eKI1hn10wQglRsLq3ez7weHWCj8D5Q2d4mwSVo+aGkdHD1E9Zci
XpYc5JWO6Gd5QGz1arSoMSkNsvooxTrvZVqcVz3yqZWCc0FYZD0uMOKoz2RbujXH
Mo2VHjtBWbBg84B7XNq396N+6itXh11hGOXUgVWImX7cEg0eBA33rgV/XqiMWWHf
QGTLe9FQuUiKhuT6/soBs5ndsMGdhEwz68OPyaXdyJFEAHekvsiU/wiTe6l9jmvK
yr9TSv3OMAQrTZrBKUTJs1gLV8UhF/RoOq+WP/K/NujWC+oUXslQ51Og4XZlgtEA
J9mXwI8Mn9KQ4Qo636dy3DBLPIcVRXuonl7hRDRjGE+i0Qcs5KEq5CApvayOd5zE
3AkbDQgTIL9V+EGRBHemEuTRH5JifIyvIfG5qsLdvOtti2YHjnsmabsOK3/mNIE+
AKjPitbWdb/2A6Ytne7oOsF2YN2xm9C6dNx5Rj+dwFawMqW3n5hGAPptswaZDjSC
Y7jpQEGNyR6pqG6L5Lf1T2Lc0bCJO+YfRPFrnpwNDm8uk514cgfIT2as94FMIdAH
NsBZyFbSDiw9LieffFBiIKajWqFQ9ivzx+EHydM6bJnGGqrRsj8vzISWMki1TG3U
8YnOkEHP3q9cyQaFvyZK/h3GpHXdFq08QFwaH/sRjq9S0rPCtugaFojYVJjQoNv/
TEZzZ0g0t+0B4GlNwpJVlZU2zQUNaqlAa0z1KEQYH6wUfAB6J4JS5Wg7L8lGdwmx
VL9PXOFDoz2Oz8jI+TPJ1hWPROeVXz2RUKK5B4QP6fQFIGgC0mB3dS9cO2+88hmM
iAZUtTJQC3jpN0ajeBXIgjUkUxQW6TaHBXLAJAEZ4rp2K5mWRNs4P2hCrHqD0Fno
nC/Q4rOhnEk5qfggZfikHuR6JUM//RmlpBzx1iuo2g1g2HXLW/t0mjR/UKNr7bDD
e/Ivkh95x4jJXYGMuPnci+oPZ8tt67MAoB4o2q2gjEFY4XJDO4dmJMolCxXwj2hu
TeGW8PqAES9y/SwcIutdIr4fScTSEd+/v99Xt04h25T3UafKBLd2+thFhDIFZfw5
hpbDO0dUydGzrIVLlxGtqmeXCxj4R5K071F8wgODmc9nymvXyQrtfbZu+L4CaZMd
SQadtrtRAikhpGNdWJ/7ztx5Tt46DT3B6zpOU9yAPY3AvXzoZMzW/8OBBgRrjJ+8
SMXzTdGSVoUpR41qSrdPrXrpzCHCmCcPQls7jkrPseMO18dyIQedw0uSMfhUyNnf
gwSTqNNuXw+m6VEHk1CbP4aOPPerV40yUx85tXriMzS6CfiEe48Xc9e/nS5UfbIy
uYkoTwfU0HrmvvfsPWrxnFvyHLbIU009M3k2QTpV8PdOln0ug3MBE/Ukj3iAQkXs
HaKRZlN25s2/YwhDl75ukGU+2PKf6VIEImVgQySApY4bi5FQu+Q4mthG+Gnnw+zR
qt6w8zn/FWVi3GDESzG2L0YK9S1GgO3zfJiErfsyOiY06u0ptPm2zoetfjhgO4zx
ASs9X47wpPGPCljRmFOOUVjYvZx50aLaKRXX/A04QoftUG7yNlT6/5sAR2GRr4O8
XL9CiCSgiAD7Ydw+FaJLimlVyHUUOPI7GmTptKZnlAy10txRowwmuG7egKzmcm9D
tI4M4iFDaxVE8d3G+3yVgWrBN30FyWn5cB2oAGzv0Tg+Xq8AUVdfPPWsSuvLKT7Q
9RBeq1GPu8vz6Zi95//uXongACo5TXhP5dACYut6BVJLEF9ZJ64dOCUwKUx+ynzK
VPmdwWnlT2JK2bv8wd3TR0vJ8srSf7SOsoRUXtWGFrWmxUEFUK+GWOmvbMK151h8
AYyAjITiOUJGcnSMuQOiZLw/uKt+RU6XJT3jofA/5LyDpiEfHEQvy74YpAqLKHU+
sdZ3d0ZI3Y+NFI6ElMKDZ7IpyVa41EeJc1kIeodygsAzfChNg/fbhexlIyBf6Uap
1FoAtTi1ymJk1wh0KP+cpCpY0DzRMUUyz7zsn0zuaA8Lu+LLwRIqgr38ptnWsqZ6
wHCRbYMGri+78sZo6HrhyDX8gI3yA79i1QiVwUAz+Yj5bPmTaCuBQFzYzgOUuBwB
obHxo83Qdinj0X7vBzVyqWa4cg8JMIKin4tGZORR8MXvJqse//53KYIn17oqVd4X
Tgk0vr5fKhQbeBAnX8aN+BRrFXW7pdLg5QsZnYtbXqSFoci+wlP2pqeyJydQqDk+
c4PJ+aCtxb2+ZGSyzGxkiY0VlrBLhA9w6nhqyySh9lYXedLrb/lQ4E/pqoVtiPoN
lmW4G7+gDRW7iPv1v+hp334k7DEIhWfeO4yui71xQQg/w4ruD4GnlMg1OTEbUeU+
Dk1dRgNdm+gJfekIclm8u6i3ux3hPBEf41dCyr6wDW3FEdc/pqR+QoSimZjXC9Fd
FuNEUoe2JWVzIr7pJ+B6be03WcKaTusCn42Jt3hStTv88vaYW2e/pNIK5oZ2oIjj
CH+bxrlT7ulsgE85e7vkPYO34u2o4295kYJr/Wj4UAhi3YPpotL3rmnSzfpJJ/xf
l36netXAWymCly+LfMCMD0AKh0TGvZOIpPI8wJ06+GF5eqclo3CdoMZFjtER07aQ
fLEa71Byc9yQJjFo/9mQxIbY0asZzPqfJ2JFNRf7k1+go0+POI9T72MATDgtGY6a
OidK3TzRyOZxUYHzABuYKDAl5lHjvPz462CC57h5r2RK8S2T4oq9tyo30Wq0JHHg
T1n7JDG74MhLNaWBkCRcJ2Cs3hpkAGXoqODp6o0Q1kDZo8uUt9LvwdqqzinPEbQ5
00+orbAm7NdAzBcGLBzA0yj3qUesP3m7ialSrZPqPtqu45DttKaBytRE8c9W3uJ2
SIGqoJa0mhlYiu4drg+A+7gL3x8n4kNticzv/yy6CyD7O5YdFeafKQiRVJjk0Ue8
KfgD/+zDuGtWyVGYueY8eVtqOaIGgjnHzhyZEju8S0Ki5GkdaN+ZQuKONFETOLQN
t/dCVW0osE6Hl9Zjkk576QzJFUDLPlJqe/m9NPzWPBskCvOHhbbdF2/Mgq+9sH5q
AYSq4xFDc9LuiQVKzzshPsASEOxa19t4vVIDZFtOPWExqebfZDVnqStJAONiNjry
PvLQkWFIOImLLz5DnJfb5/CoaYQiw1O0u4wVxpdaniGNubl2GSfl4pUeJydGEPX8
0ntp/0p0FpUlpiW1m6zuU94iFbxACemhyqSQQ2f3glj3r44b2qFf8hu19g+i48ij
57AVJuMi0fzQ/5Xg4tArbRvW3j23/PZYtsJwmsEP8g57ZmcJqSfEBb+ZrXqirND7
Vi/4AJGyYpKkB+k3IRpZeShjEkJuSg2kVUUNJB50OuJ2rxp+mTvAbyEQ6ZHsGv+7
pw2eJLsd1yKq85Baso8C2FwBJhX4M+gWutt3C/3uYZHGqitraJGygtyNQao8Uvxe
3W8HwGs7iMlLFTaOnNtNpT4TjE32uhD479fjMp1FZkyMqcJiJzzCwg3hpvG9wjUw
IkF8wLyozr2Ujpn00TxQdiMrIDjMLA6NqadlflVUKaK4DfwA9P+rjv2GYkwiMnHY
zFfBJrIsoabklm6Lbs4BGH+7EzMdoayqnrYMeH8aWevTA7io01BdD6cbs9CHoLqm
VMnNsK8dCf2iwofBKwYmGWXTqA05wL0ZLARqkqmKMUh9y94BABCyYkPExnfxoY4V
uWoIqAegHML63DyiI96fQpw0DKMKOQ+IXUR9IHI1W9mbyTzPmidvs8iQn4J2dcTO
F57wM0djckFHgkTuz305STtECMIFGt96DZULZo6auZoSe65s65oYPrteWEYplO+A
SYhzYgglhICznbRgr11dXAa90OX5gvZKj2xgHDkmkftZHqwcqCSmceorUBK7uAQn
eiPm//kPJKeZ2J9fzvy2GFJiebWGpLTi9gfRLYJO0Fl4y7veVx55fU1W0+SE2XPd
c1VUxqac8yOnJwQxsS5TnhXNhcse9Tt9YDbyNULrIEoU2XCqXOMm8g+NjbmQMeKq
N8ouiSTGYdjjO6GT2qxYzmGn9F6KPKamjhcdwunz/VPcovxQKUKnjcfmnsb/JEo2
iARopmT+t6D0oFCpprtCDw7BD8SeXPuPfIXy8RyIHiSEz0xhoGkpkALWaITs/g+h
haZfPBuwv9MtpuOM3/ig+6AHfCxtOs/KNbrEMWt27l91ItALEePgyX3DfvL0BLTs
lb4zjgEnk1ucw/3M5sH9lWcR+oFxXqdHko3lhEuJB958KmKjwyUm8NTKOOyoKLXs
+52zTr4F7/H9FO3LOV3Hf/7pnzq6EX9uHBWzOOyEfopP36qCcon3PLIa9R8iVavj
+FBekwd+/r2Db+3rARNdza7l1yczDUjH7dRSB5by74MSJiy6f/ZHRWkoIuUwHTLD
cX9O4m5oNCqKyfyuHCY19YB/UNT4dFS3o0326B6Y7dLefTu/DW/a655tmAnSaUvt
XR9ZXjiEYdJtUXZjp+8KRiVO42z9UUZaSGRKU5Pdl0sGkahNyvBMdO78ThuoZfo7
QG/CH0bIbFuWNuwRT8jyGockJByDUr5XPnTKx0DtR+Rnu3B5z50qtbecEm9ruial
AirH/rDcds/MRdPiMnd7mSNdTLvQ+L2CLEoypJ+v5TECBKMfSyFYMA5VX3K8Db3x
XsEcMjsDz87nTLqeV8yZ4DksZayXrAK4zXS74grlswLJhmC7dsKHYLz3l/dyJyXO
p0QINutA1OJfq8ndOJFZf5CuLBa13ey1MtigFNz3GtEZiEDn0xiGKReSQ5MtHUl7
VtvsT7ZkX4N5CcWt/mJaJatEg5P0AQZvG0tdyL+coakwDgynq0ZD3l6EG+HcliRQ
w70SNw0oRsXGuKMKIvpAEvR3M4riLInMEIM923nkxKVgeIAAafitn9qhuh+Hysfz
vp+98yI9xSa4lgXnZHARd9g11/5N2DrnSBSgTS8QUjHKQJQHTskRpZDnyKAE7V+q
y2K4S40MRqJvZ/+9uks8YQZP2+upxCm8ZdSgZWWeU5pCMZKRLoy0iqTdnuVH/g6C
Ek7ezXYxfIWdMmaY4A6ELWR0xworhdj9IKBhJsDFx4cFrDXFb8nP4EyvGPkJK5Sy
av5z7NdV/MqDILUVh+Kq2i2tdv3UHBgXsAZLXU9W9NSB7yAE+1QkODaOl7Vsook7
AlJ2tocbmTvMz+yEbW4iznmk3I936HzCE24/jc4VcY6EeeFO+JQRubdtdQAEkI1x
NwEybsXU1h+juX8l2R9eFg4nNnw/Yzo/KRPX7G1IVzk4LiWUDGwd/nlC4utj3YP2
sqX/O4vWKh8TW82ALALsGrSYbQ0BErsvNNkboi4aCqfBchEo1na8HLQtnVd/fpSx
3lNVZFAnrPz02siigJNyV0BubdIBYoKFmKS9dlti6mERnCAi2fGMxTr1Pa7b4PFl
8QORNoHH/N+W5cZjzIJ4M/csPguXEHUGZ7+n45xWtMSuTDeOJKDPgAcL0E3m78wn
DGQ4LlgqiE51m/ngmO9eBstOcaWV5o9dzS+gK9qgka3cMwdq+nlSkllp4erPDIn9
dmYfHVwmlB9TuwRqbeH85OTHdZRDWf0Ibqo/ZqTqQ1yEjwZtdVm+J9IdiHqdzNYX
QJJwKIFt381RKA8OGrmwiThc2/8Tll2JQv5LTJJzR0mbuNviHAEMaeFtZX1rLbPG
pJOAsi94Yk6JONZrFwjkjZMhDNuMIe7Cej0Cbuh5UeX72MaTBEOw03OEcwo0fct9
4J9a1+TTpMyDF971r7FUStpq7eQh6E0wjPVIuAE0DzIR4eg+GWzJGe1/GRq70OH4
+gwyrmFJpXPIr6YGIcnmA2b41FYisrlGNhOkRDYkDsZj3QON1YXtXiF5OGCOalfA
/W2xLiK75BlcKh8lHM6gHMZreB7BCvI4qQ2gkFh2EFRc8YuMRLa1nVKuK3y07BB7
vR6+aW04MdILIHymy6wO2ib4tDUZrJ9gKqFCy8QBNOzDEzAmwJPzNw/S+NM25Uwd
k3Fwh48MCH54x7bdvQ9mgGi8Qk9ihgKteui+X6q946ggxC9GgnFWvYAQVoNvw9UQ
F9JRldgxG96vS2V4mRHyilkZbtQXUDeNWXt8mtTNIgR5z/I2mjICcW2ZNv6karIZ
+JZ8X0ZvuJDLf+2Hqw6FwGEa1RaOscNe+Z7DqBURF5batGkpS5SMbgsrwgYNdcv+
V26M7cagafOsuW0xHhKcWogDnwSIQTh07Cjs5p7KSNGkgAtQiaxxtSDx+NED177N
zqeteKaTym2fEI44l+vbzlekFmPnLfAN/60fHiLcIVbiSMuDHyCIG3Cp1dS8QqbS
2cCU6r8LXmVU7E4gvrwyBkZJVEskq4mdzfkjsYuAbE8Xo9FevE+nvzrhDrudqwyM
RK8/tuLjptf7JjpfRtLfnXRrlIxwacu92TDNfSje1SC9rkpHNvwdUJyVz/SZz/1/
ZyYXt6id/aGj/oqg/b5sssN2HFakczLe9p+Oj3XxVC93ycAjv+eRktAqzYJID8Bl
6zq59rmTarrm3Uz31iDetnbwWNA9oEHkpb+ErAkWIhxnEmNqMks0vnt4TBtfm8WH
bJG9+ixXEGaL0Q9vbCV1yuNKOYaqgap1qZo2kFqNr2O8mPRU18eQ9Bou5P4O5aus
nuhoXurN0DQvPNYdIzux7QKNEDqTfkRr0EKK66MezY6LhcnR//PDgIlGKaqKTsET
dq3xxlU2WWhfJm6nGMn7ekozIwjFD523kS9/TIiAFanNgmm6MjKqVFgusUwSfwIq
gx4j63AZjHEBJEwt1uZVUB5Wkxte5diubHt+N097GY9/S6s/CIiwCnv7wzqEE7Nn
8TOfaFFa3Dmb6iu3/KNVNKKvAFjPy+9u2Yarfhdg5QzgVyOyTF6ZqmGoOXf3UWdS
8nnzP4iMo/metahXYm2EcEHTGlsn67qGo1mpXXco4uGcjIp/jPrSg9m/7TdV8Qz/
WnF6A1Z5T5BPSYN79lP8N0F/LkqxJq+i7DVuRrRvkdQkcAF7bl3ugZYWY0yRqtgA
UqU32vPH+WXtaSqGavTSnIBxVXKCSGGICAMKEx6Rcn8WKOm8JVRbkZUkX5sPzp2S
F72qTRJ2nPaaCiaDFkItQpohXGNO8iXhMagJd/RL+83eohVS0rhR02R1x8GB3+ga
qnmXoUp1u5xFHYcsZBsohLVAFutJaQYNKInrAMhf9uZFDkK5GJOQkiD4LVP3WbZv
YQzgu7j706V22mtsyL4hjQcc1eV8UUj9eiAZXghXV05m/qZgi32cZcBzjm2BmpwJ
oEdgMTQrOokd1p4j+oDRASmA2/wt/W/Lm7+y8kJ/80L4UihGUTUrC1QP+r6P2p3s
jF9xClEM/N74KkkIiXX1eIjZ/SvDRk9Untsym6tK2xJDpCacQO45pbs6xFjSHrZA
X6SfVgvXYXSGHC/8qfnAhm/LeLerWQ2Qga8bGWpcLoaCd/5S4Rg+RmUkXwwKX43R
SmxMbR8kjqXgY9x8MiTVFW0a1ZqQ2JXXeSnKY2XQ/Qa4AUL9iobGvkh7vAYz6F31
mb0KkcFxx8vK59S0vcGfGkwIr7Oq/XBzRu9PpLzu8k9uFCEsSPyEjIf1qBHRqGBA
jvpyktI1Yzu54t4reNZ9GPLn+r8JfU+60SqDp4eNXBDx3+oG3FZum1N4AlytKiJt
awr+EkwhQW7XaYNkT4NcxeCzfZSuDrk5+gqwpZtFt7Q38pagvVucbCAZdHTcqNML
RkBYGS83S6hP8OrEyCyrwZUCpzApYL/9c+4QX326gQpj7pHkBsrUF+9VvtOZAQ6P
WKXKG2DEAq4Bg9IQSZYaJu0BKqoEcovldPv84rZTSaNUAgTtS+NnNWYeoHLXXhdZ
PdKnmTZhdO2M99gEdYWjZQrkOIrfSzer+E5sSYubnZdmdMKnCSKIZveUbSloW36q
cpxssJzLB6vtyvF0TnXHO9oC5FyLriYto7nJptHB/+CwJOqYxG2rvyuf05TMlFbw
1P3G3hrjYHg5bVNzwQLb0KNGAMJj7P27KGd97QNaNjGMQo3UtDQhAFvpzCyAsRGe
aqR9fg8ZFdgZIwZH57oTwb7wJz5kSZb5O6Lxc2+Bdx/VVL+GhWK1AWUKD1hNqI+r
HKca0jsZx0xIVHkjtcYTUhtcSAMg+XZ2wZ28YDMeXe+YcgFiFVSIIklEb5ebbwNt
/SZKPnC0xQhRZ2uX1FohAWnZYdaS0g4l8AhXYi+22H34bC0P8BOJ4Jqk6m6rzxxb
K9pzUhLnf4Dzd30KSUX4PYt4/Crs9beZah7SoMYdNXW4WDYZtygAz6Dm8UmJhLzi
wy8brIeQzncMFdWS4A82l+OYEgF+JjvPVPEwHdu+gQggljGRiikyZmlslTmUvTq5
M0na3XWJNr1j4FCRk6vGAnf/u0m+GrgXW2MtUhWpnfJY2Fa8RHe3meXUgUJ1fGQm
PLzAtgheaSDbUnMvSxxAdXRw72JouRijqX0BrJqiL5YH6rKq06/8iObpDnpVSSAF
g3bFUj+JFpPznmGkZEX9RRlkCp6NF/4dxlKRr0x4IqunxqUJYOlDm2mbYuCZY8UD
w7jXawhMahntamz+YCBu0jz3LlgsJ+1zfK0ruQIrXZV9am69euH3UILgmauW/D0R
rTemAl1i5DFCJSyqVkUe6YOS3jl3yuwtJliFSNReApOF9bW7W2a4cq1fwjCtClSU
lj8X0FktrDGTlZTHjwr1U8wcHbkx6mW1Pda0Z/9YnMtKYBcFfeQots68dXRDQZNb
ELSW9kRicedXQZ+QjBwzDvpetzUbQud/LCgu4BU0JDAthTztH874W3uvMD3X+k0f
TISYgMrYSCdVGKlHE5/8qEKXEoicgSQq9oWmYV9b7WgWLyJAbZmhuJ53IiHaT1UQ
IWvYrF7WgzuqYiMrj+qAv8L/MKRqES3v3tqfjdBvfr8tfCHCWb0kPmE9ohE3TXqY
b9wa9/kwt09aXS2CNbOuYeioPpiscuP9gPt1W1rkqqtxbaZtPChSFYgrrQXpIODE
s/xpfacNSOlFMu9QFgW+s7O5mK3IcDahdse5rv73wzrD4iegwa4wKbisxw4l1Pvh
adhVlPc2Gd8iv9Jbl1HdGI0vbToqGYzvgLO1B+nrI8QdlZRg0uGIywXoB1BAYP/M
ValnFRyKS0c/PRcRHFhAu4XV5UwYhjNlehxSzXViRt8RugjfNoTZfSUDiX/GkRs9
Qp2ZOlNchnOuCgGMduA42lLSByxRSb7kyHI9DLxpeEfUE/+JY6IfMq8ALfaQeb9n
+SFoVScbpt/odom8tm4oW3isdlOBbQ5TFRPwVehb2FTbuFVQiMgHn1uy2aqRw8IB
Qw8YW4xQBOpbh7Diyw6dUSAqRbs1vCbrTKt01CKjXSrU9u2ept6GgHetKLTlaXSi
jxnGCQkV5s9FcQCB9+mYlhd3bOLtp1irN127DewcLfbvZygHh36PpwDef6SRC9x4
XaJqqxrkL/NYU9yvXUK+ij8mq+rkPEm2MAhuyKAWsoVTHwfAqc7ejl1sasdaTGoB
fvvpEpVC7LQQKF1yHVKTtzzaHLmDty/JDByG+Hfz8RqLXECf8yvjWS6uvaXvex/o
5ALoqhCvz0xTr6L4icVJ2jCnT6rZIYdLxk0JSaNMDZ6jUrq1BbjwEU4ahco2YrK5
LsFaKLX6O0Xnlu+Y4RZWR5tzexoD7A8qaLdqa11/uCbHas71wNx/Sq434GV3U0L/
qS8y/yU6EwnRBpv7velHxUb/IhEP7HshTA0xtvvlna46qctEHQbykKczUEW9gx10
3cgU3T89byHWdG7l928YZO05CCF8qm2C8UGnNGyFxcigo3xQwRlh+xPIxlV0S4hd
Rgpding+d2a+VBjPL00PY2otpeRkFOmk2qhOyWmiy6XcAMXRPkNKujRjVXEBiU3V
MmfcO3bYyASk7IkyhFfkRqsVWDMmFByV4IBbN6FtbGs64N0UFQox6MDMAsTyh6Wp
wFEzGkDK5C8+wk938nHVH7TM5Vx8tohm/hLjjFBhUORb/h955NipXOC6TNm7GGTh
wOa6vA/3+8Y/XjB5Rw5My6GLQe1ABQiwh6tMTpaokSY4XYh7o1iYp67TmHriVZkL
n7N4tvHZge1dwOWdJ8rUEr10VSJFAuocoGAf8s4lIZlk7DEXvUT9yVwUwUP3ubP9
lZwSyKwHdaSjhaIm6cXrnEa7O3b3dXCe33MPtP6qRQvigw3jiHJdah2XcuXu0woB
3LASsM7ObHlW3KPTR6Qde4dzfriRaewXTPQvJ9603X1JOa8J3rRDRzh8lLhnuq2I
ARoDdlv0GkKjkanW0wyyZEjJz35mdDCV7h3opDLKxpTapcEEQZx6qhgQZYcbaAmB
zfake4wZDylj5rsWc61nPh6zx0rFCsxxkgjpe/U9byAS2N8q1LFKg0ZWphmLao2X
e3wxAMzAz/ggO6wQcD7WT2KVRyK0sgdXpHb40fv0XQtsvHedD9fReu7JQVwqgM5G
VPb+zlBoeb5H8YUkRMNRveatQbHgx7l9mG01SQVadHajW86wxuCS3jTAwCPQo47/
qiPbfwitksrCrB+1yEFpZsr3RV1PaFrw3HxOXnlo20m0RNYBeKrRUX4EbMziAx1c
h3BeD2rtmeIpotj1LAe3XbD5jXn9VpssguHrHOW7kqUJgV+e3yC5/QD7+gx1MIgn
FstIAvtFmslRkvbWiFQWRRbyOGjG+n4/NncPuO4PFzbxXyZRmIexUdZiuDXMIb5+
xFimuuRFYOv0RgqzQ8vKk7RPQ2NvSWwd6a2H+6TOXK8yYw2Cy8BV0yXm7nAs9mxG
XtO/7nCSvARw/Ln78wz4yDLd8+WvR6EEEv3rIcXfFUDB6UT3hxXuRoTjB5Ve8tO6
3+qxTP1PJV8ly99hYnxjpvf9lyVv6px63PL8oIvD6kMXF/Dl24tbLWtihRvtgfc3
IIrSlIpcmuNMS4tN472XgcRGBdKzS2d5w4Z5uG9bNnMutQri5BZ5W1b0pZPPDUGZ
LPDQAz4Ov1ulv/LHVp3jnY7FUHVWr34fWU2rzLydI5Q8rh0QqQklT949Z5u39Fd5
qZGx3fWmABU++K1sfPfDmaoCkzdkcL3Q5wi1Kr96MfbsyPz8nddph9bfX5n3Uz+f
Ceoh0XSGtKDoWYVOHcaxTqraNc7l27y2369vC5p8LQAxn62e+r86nRmqpKQE4Vm5
SAegnc4VqgZJ/z1ijkqYlHQOAfIcBQ1TgQeqew+38saH4gpsmPPfUecciTTFouQ7
34XDeFJ4OpS0WbUNO4ojFtMZ4lZIbfxjrXpoJB6VDAlioKspPxfWopQgsmvD8GjV
Z7cWAvmQEWHAhMuvPSIOXBPGET3Y16AwbVIWIoZgkFZhClqCgcfm29m3CmsGv1Pa
ePRIoZc+tRAGyi0zub/R1mxGMLnVcbVKIpoxC0HCH5gyK9jrpiDkSRbxV1cMzUty
4RdU8yvAWBW2E5gNF9l5mPL8gkTzBe1hgCPZFJ3hQOfuYhuxkic2I0gMbtiDSwBh
+oCxumrO0Jkq95TUhBL0lxzSWkfVHu0zcI/vv8pZYrLqo29w5/K8InWOZIGlC0gD
GxGAjIUR9BBd5vqkSfCoVQsddI0dEoWAh8NlemlKzACtcI7OWmGZjspVCkMcdH9j
P11HXqeTK1qDAKwqLRun505je2I+y9Lp+QE+nXg3UvX4sq+qhnh0UTKkOxSTn+jr
qN/nQ0HJzwYwmR0C1dtVJGzAc7gm92b8iKydZA+w/VBrigT/8KbFjba4JRRtQq5J
PNxe6j9YibLGSY6hSNP8uSWDxG2QaFYPTTvbitnJERxjNlujvIVNB/FqpRYAfm4+
JgbF3jTyTV8NjlA1tji9RE1pwXvJhthEbXLK66q7a9zb9+5YM/gcmbB7xepyIH96
HYj7SOU0RtkrQuVzovUe/sj3rhHKmt8vmIs4FSnaJBnyCpeA3zmngaowvO7q6yiC
dEIk3JEX9aA8RgfFtbr0cgs1EfF6Td136ISCfJXRfF5WqpcXfYkMnC1tohhNKljj
A/5AGsKMpmUma/lUoKR97rLr+V/eO9oc78tzkpzWKZHvhVkBtN4G9XE/V3nixZJ6
Se/9EYOY+PxyokE6hSut8zPr8amhdApl+sMIhYt6fEWMfFDkA0A+7xhRBL1ta/IY
x+wfOHu3SpJ5XAcQT81xBgw8M2LcDygjfP2JxSXbu+nPT2KNYgcqkf0jj779+f75
5o1Mck1AhzNRZrvyn6Km/TV+ncPDEMwM+IW7GsZvnMhF5yW5iFwNC0i9M3Ngp3Or
SsVNhCz61oP24GteSnyL1HA2Vct3DxQP1bbfT1dpR4nIEbCc5uOpR4VPLSKSsM2N
JTYnZDE9NJqGNMwOCVYyDgB0s3vPlSOa8PWfMyPRVUXDLrviBBDixm8FzCP1Mbxm
jjeCVRIwefUAlVY24utsQux/VJwNgf6ir+od8c0P+fQUVHIvsc73H1EgKKtpp0YW
mFiHQZYPIDXwaU7JtnOJsbEGiNXngvthCHl3kOcb5MP+MVCpLFmCfSLsvJJpleDI
CDGTbP0UUDTq0LcAimtmHRw8BV12uqBdgFceS+VITfmC9NluXOEyWEeCBKpwYdvR
l87cFG1qu4646w0VcVfE9W6VxKKJDm0zHJruvgRml5MhQY/V62R2RsULK5M3cqA6
/u2ws1qIE1UnmxzHOZw2YxV2CEUxFNA0QkONn+BKOonxUCL8bU0ThDvSbNcH4CZl
BwcbNIIVXgak3/dJEChztGA7nZ4KHlu5LVnRRpHLSqrJVFcwZQcZHtMJU3kY8jEe
Moa/j1yytcCzD2wqYVMu8qDslrgCsk8Wudqv57Xa5+/8FF5Bu0y+msSnp+FqZ/mS
c4qTFgJfFeqhTbzKiwnLBefyTGHD6wjAD5XTbqwj+79+PBxt5MRi+Ufbnw88iK24
C+yxQw3tlpvQ89IIGuzEHgAB3bw78DjH5bbBqGuQADhUavV+X224SLuBqzI6Ehqx
xVWZ6xi6YJHvLGF02gECtw8byq0fSWo5cvya3vCBJXEePaaGGaqDQO7dlJEdUx7y
PxXZh4YHAY+DnTYfJLTztOnZOvkAJmGl+PkZ1/U4s0SfGpf/RDOLSfbfznPYUUiX
gYS+KPZP83BrPudYPdwDNcxmwDoURb8qRzIJ4x3dB/YgOBRCtAMuPOxSHXnwvFB+
PVSnzR11FCBtbSQoT0lwrJT/hRYzc0uYFQudjd6TFxOz+R8Qo0/FuOCs4FamDiVy
DwcrXMndACNsy6bzPb/3nBWMmZes77tBkyrZkvkty5xOhapUeHbcKxfg95QgMsmR
aQyeWfhv30OIqF92kbed5S70O+hc1Nst72fYyBuSVh1fExsFq2k70IC4D9p6l7ag
2R+siKjdq9xBtweFcH9Pe4uwI1mS4uRUyjPteYWHrrsXd61kOi9xYLs7fVcznE1G
zEtQ6jJ+KpfAchxCdTbnASfvgrtdRFPJRXyl7qkyNkNKFN3V2iM74UcSIAF+zspW
YUq8aaEKgFeodTV+ZuaxC2Ma94mJzhZ0AWdqfiSKnkPJIjfIM0RFrgtr9WRgxBFx
GNC3eWlOAzhqkBWs6Hnd0ZVgwDy0hNL6WDpoRXE9FAHBAIQ1L/tP9sC2wYzwZz7k
8VypKn706N7zVE1xtui5wRGzkwXesCID/gnjNTYQfVtjRaTvxc7rlEgaMT2utYgk
c00GuwmNSHiXf7DwP4llPDj58fzUihemCKOM31FHaDPRMGVopMCFQxZodoLsS5Jv
K3zBcQ30C6uqGZSSpYU0un5yO+hSnItAvlehw7mZUvnTdHh5RqPoT1c6dbWp7ygp
mKrD9miQilEDW9V997qj1kQXMOSoh9UeS0AVkLKcuE3irN8cb6GiOiMhhAC/4WIy
rWNKuJ927yGWoUGRNJ9Fo984GULj/xfE8KDA+u8KR72QR7aTl0ZMo6u1CxF5r2/4
rIc6p9wXXGEk7dSCeUeU6oCH2wOgglbcXoVrL4yNIaLEhgdM1e0lYTukLmx2Y9BG
feT0/IXPUk0GU8WCnrUBzCrxHo9GpJsUixbwQ3hinT7DlbCKLJ+a3XOfUtW+SoAp
OHUPWmsfq5KDdi/aqjLzF3yG+WOOCQF5KmZJg6xwxUjpJ8z7SgvAxXNQ0K4wJ6Vl
grhFliOxAOOGcbYjnjcGzvjrYz6u5M0mFo4NbvMt0T/jBh8mcyJxJCaGRH/WmuFQ
7AMKvPtYTsoweyKLHYDG3yYNTso6G7Q5a96RuAR8ZsdXOFAmAMjNSJvzKiUaiM9v
EwFPnJX//dL56B/UoG2tQfgP77MBYir5V4ADVHGHrNeYdxtXs+DXZnTU3s0RLNrS
M5wj4p07nGtdcSY73wCX3v1Pc82TZo3XMU+pdoy/lSnNC9QDFiW1jx47HM0+YURU
10rj97iSPeOtGEyTAkihkKc/W5DiXDkj5zxDrc7OST0BNV7dE3I01Cutut0XDRck
WSmE2NlPvimUUtVX1M9S8DzjtRtGTvLRTWwKHkbkW+7J1ys6uawoNLBnqH3bxlsX
/f1HeGRivOjQKoZEe091pKikOTrJOlvrj26Hk2kviyjPTiNmZqN3pBuNNtsX5o0t
6oxKBX8poTvATCINui2jWo+OIKldH3xKqTiuzK32m06mUTPlgVZFiYg0ekeFq8zK
pulMxyscLQfZtTpRnNHB0X5eY9YsqsZqf2WTlvAJcYZw8+mR/nDruL3E0kQAn3MS
9zmt8U5PUc+Btvut99pJBDPkGMZ9qEQG1DWufjORPCGV0a6e40mF8nY1bK7nYSLv
Uwj2xoDAWGALgpEEwkiPsIVAeoAYBQZYpZ6jBrNGFV1Ve40v9tLUWddM/PVa9H5M
s7W2LD2eunKQkzitAF0ofySzZvcolfCl5LPvQObbY24uOC7EQgHMOxkVo3T9k5qj
CCZN5oW2TCgiWoU2H0vKLMCXCaTUMlMP2SSM9c7dI/oMWTgnBekBWUpQXrma13xx
dIPmY8TVYHh41xWwZT3mn9QY88JcF2qbFPVoI7FKnFiYLRZPy3i2sOeliM3F99rI
8vzTYSn2Pd+GyNufsJQ5rMt5/kIZi7aJrzBE8dztAX74fh8GXO/bk21Ncq4iiXDr
1r2pBDMZUHw8P2kiwzuVAidNJnoFlWchKKxJMhKLz7y3Qyyvo8GwU9Pw2I8MvoLi
OXC5iU5LqJoQmYz23ZugQvNKydUNrsVVN3PZb5OV1JgEcf7OFiNScL92mKFaultm
UxQHnrZev0oQIb3jAlnHvpmY7QdQpJVukC4hBwrLfx/QiWIh3kK/fmmtlKe2V12i
OJNUU/MEJ0jyN2On+nq4H7WkM4zqfj5R7B1CFMIqoNauxLrmXbnRSI5V3o9V7nGz
ow6LrT1ZSnR0zsarYNzloLUlYjAzdOCSjdrbxUHSVvqoAF2N/TvpTUJa7XeCthfL
g9NPJPIW+98DW1aFNde8PRnGW/mbToIjsRYcN5FLIv0dQGwMyKHhsSsXfxwEhQx2
gs6KGhK96ZH5CYYBDe4YzqruYuK0sWBXiJole6o/KS5hWKLtBKn6S7oYBiPNIAtv
gE1MoPrSNV4VTV/XXYaZ57UK4QKWMNN6B68+8sU3I8xjV2145HRoJiDr74xiuQRK
oFvij4pSWzNlthN6BefuM9N3Qwi2EOYchQa07epT6WduWoi0W1vkV/QamYBdW2v/
HLaOWLV9aHmvpONZypJpjv6v7tPhKPgVeFXcbHJBt30w05bVmfPqliLD+hT1BP34
9mDjiEmF3u5Hlv+LL7ad0TsIfsg0KMzui9g8qSDgzHiAlWK63CZp7sfHSMxWxf8i
xJk2sVHjkQBaH98QXEBfHGHlL5yVg3fH59YY7DWGXhA+Eb00LtemtxC2gR4ff8h9
djSh/1fuK+QMZf6P5s2puugLKV70ky2nMJRhk3pJBeDzEaHS6qP4G5HGxg+Oyx3F
HQ3PJT5RgTbJXq23ImxcStEiIgaUnz+QrvtNKx7gSrXwQ4v5b6uZUgKzq80uLZSf
+b/8kHhhpuQOGklp9s+AF5onMdwc3JYqTCJjwNPxXU5Zk0AbDFXIOh2LzE78GOGQ
Z9D6QVfVNgsfAeK4yWwV8CqU+hMBey16/tIEyKZw755wOVWssUX7PubLf1Mn5DTd
Mf82NZrMdqsakC76LeOI/YzpbHbUm7vMXbKzm6Op/PwyCfsu+Q9uLHlKSBSwSIZ3
Sf/zkEMDjC4ib8iygFKQnaqumZl7FWLmPVZH6XMgg8zvhRGvLG3R6+O5kOtWV/Sd
5BcR3JOEn2xtUbsVlY2THC7x63v1CnGrTWeBnIh8oJv8ouF2kKOVN+X27irR+egX
amModfUKJ2y3ileixhokPbCFA+lp+GRl3iE9KYhCgUpV+ggheiI/UsHgjExdHrnv
5jpXjXsyFaXXKhACPlSrOCUFwG0MFzX34b6RADmCaM4o+EUFNGawcgAKKTKHfYd/
gGd6mVuhTFQAtHtQhZkOQBSoukXIfAJ0BsnbmOiOsGeL36qQXsrJCJHky3mRrt+k
xzp/B4eGtQReBivPQ9iKqrY4O01PjHxl3ibrNlOC7eFZZt1pKsxyvk4cQISv2Nym
i3oIHuEa4fLKQiw1tqnMlO8mLUESsVDNWlUxNcCLmu89eEHfmzXjt4PGMAdzQ/me
Woxl4qbcmuKRlX4vVpMKMy7ehDRGLvdg8LEvLzDIdZTes0N0RSnKWOCpbNpGig3G
U/Nb87NC8DLrc9/nMIvGRbKhJ+eY7UXSgMFSimu5Qitz4xDjAlxhhWBgoYGhtRwy
p15tebpeCO/YKI9ZlwKXbKVTXVqqVZtkJRqJXfENbNzxqQO+5AeusQVf4oV4vZdW
TD3c4LIT3uiUXXwReb7e/ZQfGjdQjtvm+/WykK5wuE6KnrUzlkkK33g6FBE5SoBz
ouKhyRCDl/VEY6YyasIcblneQ1jMIwHt1HbtRpWv+HTOtbTjV4jjnrKzk0GY89o4
Iq1JoPZuBDgtR5xsUSI22HJqTU+TwUuTi7lWkDHzGcC4e/K82b8i7Oou0xbPx7My
Fc67oMgo4VdU03gUM9oBJNjXgs7cMbQ2ZVVV/XXLfRSseyfj6wqCW45armu6FW0Z
rTmugzRGMXr/1IvLB+eCkfMPSZoI98E1fTNOVDsPeR65dW3zbQT3BNPoNHHs9BNu
2k13+NcNGVQype1xN6JiyO2oJxEOVX82O+WHn5GfIRs7pkqtk3OP7sSPBrAvNggO
o9b/ThRXSoZAM8FJA0nyAZXV1ikrEnKSty48RwIC/CweaxHFkIgcZ/t2TLZ5jh36
suZEOmUtXkdEkO/nfvYmYlPYQSCfEYgQ7BZdkxdoR1ho2x0EkAxmiZA+Ezt1ZquV
qjzIxHZE5EuxVtyvj0gERV7OIms/IEw/sfKE+ghQHrCBSfVRqrLeHz3dWJmEh+oA
IhX48KnTb1u6mS8m2PHWcGHCDnkjayKWZoh1QEuYelKy85DmqMIPIpp+7rlMzyzH
/USRCTIXt5K47PeI2J2dADthMFkBvm8vh1I1fHKCy/GUAzd62eQMDkYvsVH4ksX/
wTzIc56HFwIV4AoaLWw96aqwrWfQSzyfjUyenj9IWkYfgzD3iWt/qxNHtYC3VJDa
IKySKZRp7eRG7lCVTA1aqZFd1HOe84E6YpMXrqZhb8A/GZhiSj/BWdGaH7ZHb5WI
VR5GpD2o6Vym89ihxV1sBnj+NEShNrbyZULnYlk7nX7F7G68EFWBEySsZMzpSlvt
bBZB/JKcRrGJyCVoWqVp8pRkC+Cm5Yu0LGe5xH58vcWKaG67c6edcw4Ew2+pArmY
uE5npv6WTcBW0pOvdQ02q22xWOM9xQTYR1L6tZBuYJXTc7Y/Y6sYCqgtl2rWQHmF
ioLIkKJRe+Ns1hD+iqV5ChTE2paeXcCHrb8DqwxMfEnMqYyAOQDf7tEUJIVp6XTJ
Vordzu12udeL83TE00mNIj+3atiUQLkj2bDKYCQxci+3n593TxhSixqlMg4PL9gF
HwEbrqLnNl+jwZmQb+ZNhjgzK6ElYdyrJOs6R7zuhUSotUhVvQprDryQ1d2ndD9j
6gD0XTqNY0wuOCRV9jXmIEZxH8ao2AYS6vaDmw07/PHIebz6hUdNj4tCcKAW0yO1
Rdec1ka10hse+/XYjU8GNXOFJHa7FbWHK/t6jW2d9NYQ0ZN6Na4Mu/B6Nryvh59P
9B64S0stT9PQesQosqE/azoqfHT3imZKGD8xwTSSNWcOxNlaVrqgi/DpPs9ocKUD
Yn8/HjejRXR7Cn3GqzVTmQr3pGIbJ5jqm4enHp24Ry5igCM+yqHnJjtW2HVcR9nt
39BLuuXD5dlkdnL9OPpCcb5H9SmPNz8DstKrTjNZWRJ4PhcmNcgoSP0tsqouJWtS
qfjapsR3y0ZUuHvbtZ39A03uMUVmuPraDC8EFnGTGBvXB2kj5j25uzj738PuZsG5
Ax170+qqs2HmFlIvqCdbvo8IAdcJSszJQVVobghiIQo149NqYDNqg5c1rL2tiJzZ
NRAXliB2AGCf2iKvOFu1DUEzoB0oRNKK1xyX/60Bhs0wb5v/b1TJjWcd35CezzME
rBLoAbF3i2jFZgU/drjQWaY3x/lUZYZnYOSQKA2zLuVhdjfx09MbmbOSJBEc7fyr
gNcYnZuWmnIPpoleWVptVCbOGDvSIwrihmHbufGEvR1I0IEL+vlU8Y2TBWoMmhzF
DkgW4BkYfOOcYh0j6uK/+1481vTwAWUOEIiz4JA9DofQGaulwtOoGHhCnWx3eg7J
G1fpQ3RBZj8QJ5Q+wbFns458mXOSquaZVYXokSvZN7UQ8C7LeNIYns0YKl5ymwms
SnSbrNuMfEU9ipZnscI2d4qqsc/6LEEi0hbnZUbWq067eBc63bQWBVHY7UiOi4oK
GC8TSfPfTHv59HQ2KeKFQ4dNkt9j9Gcd6v5O0LePQX2R34xk1rvdia8ATckQtxDb
5sgbd4K92B7PP5WK2F2OgocfQ5aKBjY2usK4yzYxxAPZ4q3LFjxLnkEFKIsFcCmQ
mLaiF+PzGJq+08mYPJWnA6ne93L6r6l81dYJLtFGvabgIhvMEeIPq5F7c575xwPU
lGvYIXqyk+kIYyy9PmDO27MDVUZ8iRGGlrL43n15QaBurNiFzhPSbo94P6rW2wpD
Gx2hd3YFs6Bs9NLlHshp4wObynCD44xXM0zKbiDTO80yukBYu4YY9X1L0S64hUZY
3eMsdFvEY9RlA/h72yCGGfw4FVVMaqljLZZ6T0geJVru9CSBJpfSwlgW1AG3b3YK
GFRJ9lpUAhzarUVdiwCIJLoehvn2eFDYiWo1ZnW6rVkemgtXPgQMeh/vvI9FqXkE
70D7SzOYZHAi7ZAjgAl3qL5ScC8Wbuty9Mez48oq7IY1vJ9sPdY5IjA5azxzEN9X
6RXETq5inO3T3Ks+sv53mY9V8zd7vm2Eyy+H0Q0O9utD0hYppalf99JcFHHMaV8n
z2FiHfpDOBSu5c+NvZqHw2D8jJEmXfNPCG6Ad1COpg+T4zgr5nTbibF3GJzW4n4K
fxIy62xW0DfU60/p/Izo2zNPcquEk38C+rAwRz5e041cfnF7qGklcn1EZyv3uNuB
XtokzrnfcUwYw7GWrAbh5Fl9Z6fos0vvEdJrvbZ190BMFPg5c9UkH303Qgl9MEUI
2YtrQEwllBBPiP8MAZQynFxdR0AGTNJ+r9uUToliSC83wIje7h2Oa4bTNOW+mYUU
XfvN6/vo/CsJm3nLG2AZAPHYTXoQRSjwEpLejwqJhyl33LFj8HgqWVESdVtZtUIh
ZNuWxmRWgiFnDtbJIYoyUyC8zx8kL5PhSnDb9A44mb2iiGwwjRY5GFsVhLW9dIeu
v9GuxrRsj/GqSRhytHI+Dz1jyc0mtIf5S0VRtPCTMtq2fzCcBJ3QJ0khzfazKdee
Q+//gIMWG1AcPyskUiPwklU9f6eMvxFjBOPdEhp3it7dnO+BgnTXihrMnxTDPv0X
Oltz6w8l0irIWPefrtvUmlvFm4mQJ4i0cpCN2JC1gTYhyzMYgP9NrWn9n3FxTlsr
ZhkDYgu9IGNElm4UcRDk76AJCGVZ92zX1VdZxf0Id5dTwBHLwM2b/9HoB9KpkH+O
D4Cevl/fGPY8wyTWuI/hJOhrDG6GCJWSC+hhYG8vgNiQY9hIysYnWE3RAMMAQvH1
RZD1eNWJkDLupygsQOEIomGMD+pULbbbw1p4peQvjxKMAHYjSDBZaE7XbxKgNixY
pDRhQAtnmH1PFoStYr+xdvMFk7O8vZ1ApvE+GxaaM51yxNMbrK9Tw/GjYFkcnhyh
ctwuYKZW7BYNcdNQBbB8u4gu1LD9zosc+tjF02tFbAB0ZH8OmDlUIrBoQUy+rz02
lqSIjdEZ1t0B1E72/82qQZ+9rKa1rWsm4I5hEv14sdNyW68q1j9m4G1J3qbWeOLH
l/yBCRiaEKMsOFCp0Ww5QsDgtTqCbIrgVDnlxj0P79Zvmao2EDQh95fL/OaU1cIG
lTQ4A3c8Bf2C6sBsK14tpREgVR/rwQmJzbmSB7tToD9HjsvIFAZYbmqiiGCjW0+7
3cjmjW/CptJR1PIXv3D5hw4lnLP4XoFm+QiaqqD9NUWEIEjP/OW5tA2e5YuRoJOw
erQcyhndMvh+Z68D4vYDL/kfp3dTizT6Vzg3GFYm36ZG+suH6Ydho+2+N/YiTFaQ
WIOXghgphwQOiji3RVS1a1GGrBFS1lqZRYCVOw0/AOr8cnlggyo4XwP0NHfJ37H5
CG6kyNETYd1xB95a6wplgvgs2aat/FuwfEoZD0Ur7YRM9Yh+i2gc59tMab41TTCh
/Kxtqq4a3Rj8BcTjc9K3TWPw+trbQecWmKDXcknywGj4ceKrLr5Xok2WE8TdaiZR
6yQUX0T1cWFWfARuoDbE2y4DL29MPO/3lATHSJQey1zlZFj+nr9FL+0HZn6SCt5n
G5ekZ5SaJuvNxjsCZ4dQs03n5Tw9fEoRwzNSm7R+CWLOs8VD8TA4Ih+7d9UV331l
hPqqE+xKw4RG5fjTvV6X726Gn7DSmxc4wAmw6713GWvHPt/mW4oKDzW9O/d7pvQa
Dtp/rpui5zfLX0ct+UkONHQvNjWQPGVyBrYANv2WhYQBCcYKhtUaOMHvXP/KWteZ
8S4v6gdfiaqOPMuMTH6kZDgZVul6i9EadAbIF+2kALYRM8VzAXHqp3g4OD7JYPMW
RJY+/bp3LnUPRGvWknZokIwwEk7MAkf2C+Wa2gs1f1ZvydqjYu3mnOG1W4LAQGx8
WwetLh5mpP1YcKYBdCNKWryhD5uD+UICeQ2ARbEcuJUqW+LusRCals5t89oa3nn4
Sz1gX059lQ+wlSV/TV1lEMvm5Ur0LW/MeefLNP6vIK6fFdY5DoRiSbSjH8OdeySf
oULlPQPO8sBlNSAS5ES3m982AAD+/AmVgsMUi+g/AUqdwYKXdAoCns245qCwY5zV
hWZR4AnnmovnqloxG5gNdDgynm7ThdGQLL0RHtP6InoydkXZHG1GD6IbxviqAGn6
SGTtZqt9nEvZKYNNTPWRntLehcDS+s39iQDq8VTluJUN3/co4KEmYiGc2dsDOBhX
HJv46N3nd9zNccaWzIvdugGyZEyBaulbJdPeiehlu+CUBpdtThqZ+1KMSrbRAYDP
LrYk7fxWKH+/ujsxRt5pqtJP8Lx3WTCRfiDAgQf4JY/z4jxtsxdjgsifOkeawnQB
idgZa89/O9Rd/txd58A5T0Y492VhK8HHs83zdgOmaQhyJ//4QyCGDXYsY6ALi0mG
i/gkhqzHbErT0r3QDAQ5q7bc2ZkEDJz2RkmqFUOmqub5BQ70O7WmCGTwep/RHeep
89/9vNgb1QpgeDsm1OLUT8UsOqDGESFd3hRmW7tHTMw9vu0MDrVMK7ExqUlHwLDG
KgrvAYp9IZ0zLbjNGYgds25AiBuFer+kFVim0bRiqA26/9dJnV+pVKaqDVM7LqYu
t+nThgnLrXcNg8GgSTN2wyPc+NGz31nDV2r10ghKebujfoGTLxsJr900jIZPxS+a
ed6pC/wJvjngAT/SYHqwqzEXLpwpRKdMw7w8v4hU6OVDwxDJ59WzpMMVYHs6Hfii
jdFssbI1qQM3HQxocO80zZNbi4PAVkNTVdmcgU96PepGqKi5M0CY+DeFraXetC7F
Ul6Kb1he31cR5Wegurbj7DgAn5rTFjwFQ565kjqkIblaNszH6wkpBWJWjDQEXF9u
Y3tAUTXZ/OYecEqXk75KekfSAvvD+DQjbggsxNAoV3nshde1xlxQvoZYomm47y0x
Y3Eua3TB9ly7Jeh0Aps9zwf7iOpzqZWZBr30d1i0UfhPSHGVwNQZib9uTviGuM1d
aOKAK6V8fsTQEmsrbTFi+q1+ISpmMHo7OEJfppOczDPadarS6VFJV1Ma2i88k+kA
FcoGP6SbdhO9oYe3I4IcWNabsaFQIUNlToqwkgcVKOrDk4aGS09t0oGR5oPG9axB
kLL20tW5NlPiNMIxe4TBipaMXM5XtC4n8g0/EK10TKetnE34cji21eyGOhcPeRzM
wvA1een5ostNjfUS7/7AmlALJKMH4rs20IlRwUHgwHikaLisnM4A8oGpcBca/TYy
YU//dwZbFUN1krxdLZI5ffPteHNOhx9r7CLnUR3hKhxCo+K4+bApxbKHhZ0XwHix
HZjADnOO1OnB707AR5/aUipnT+t/QFaBr+gnXVRsHZ4xGkpWBSbNKIdkAPxH8+m2
dvV1OTBIPXVFqmOwphm0+YtBrd0FfRyelwvsQDhDd8GLrc2XlG0gq/BGH4Hi0tQ4
9B4aVOykixvqPf1o2d93jG5G+Oex0Jak5H6+sYk3Cfx0CcXrKyvqyV+u2OJOczEm
XjB24lomIT8UV35QpPeBJcOr+w0njzRyHHZqxCld+XD+88NznNjQwjxke4NeI3W+
7zqWESDr+xYXa8wir+StjYjjJgycHd4AFi/+nXvTwPzBHQo0MluMNSup3iA0A9cv
/2hLxnidmTjdpNSSKz1NcQkaSri6FDS4Wr7BTJivAZ/jCIoZ+IbtbCP6nKxEWRF+
kGlnQM4HdP7GWhH1gXgSO3IYrH84sDYvUKVBpsXmLL2oqMS4cO+Yb3kzNoZmLyeD
IrX4tRAfRuXRMhVxwn5T4vRsdKKgpL4W8bwrj1j1KmeBJhAOVZqWfESuvIdI7vmL
I1RmF5WmOpqALm0J3ILFyZ4Mjcw1CdoeSxIhRtG/vf1GlUeJ2Nf1+xiHLqzRrsXk
rH2ALRtusnC58UphPyW+6ENDoK+QH/GPAHGtwddqVEHE4ZYMu1rbsRZ+fHW0hpnO
+f8AllaFLEMOprcnKtSknJSUpyK/g137U1sLKiA36UloxPniP5txt1tcXJ36roIz
lYlfd0wnTevBO/UtOJYQZbnTKDidniKWcNU1gO+4uo0ykEjq4GLmSGi7nQdCp3AE
1yslth93p6XXQCmKWlOhHwNYo3PPV6qlWI6AQ3t/6kSQzWQq2m1QAfZblmUBbLel
BlVM1ZgDP/EdP/3+lzJMBqrCcYB+P497ZhydCvKoRIRPa4e8it6b7HcPJS3WCLqe
9T6LuMD9opfhwsYZg1eibofruZ9Fq4ELRjBGUKZstBZvsrEGmkAbH+zwkLnJiffa
IfA/76ttB30v6uWN3FFaYgUb7eGDwzrIEfn/1WGJC9rkz1GCltoktuxa+ciYUNFz
K06ybxnuOCllIISvSRhU+eZzbwyFoOvQJwM0Z1gzaHvlYQEvpJ+RZ/xSDZ62sv6w
UKHQ1eGNs84PE2RW/SrL9CaaITL97PTKRt/KstYM34AneAK5M1QbrFd8YN2/iXZa
MVJ0cBmpwdwQoOZpV6jiRRgfgjDI9LmvLZ5H+9h8ea5IzpH2ORIfKSFFZ4vF+jAd
sfjJGsj2j5J7vX0FfY/XEiUdYCjy4DoYvRybXD9dz0tZ826XodxbmZktYnlmd68a
Im2ay5Ha4MsvtGRnvuJX27PLI/hRd+mEeR5jOfk2boadvRW+Cj0QYQILaACTnbJr
qIqDFXpcT9PopD9QEY4dtLuiaBn88/Zxnw1VHyJ55wuT7XwHoZGLZRDznZFcv6wp
wZobHTfDON8+6U9ZvoeSIJaFgfqaORbiIFZ7y5YK5cbDcCdFYZnPepChYzigE8bs
0+zyVEolhAI59Bm902UDr7SA6t4JZSXOA7f+UwnomPpBk5200A2/nUOszHws/Ha3
oGltsJYFPdVLS6Kxl4kIOyPTYVxKMhUE9IljM/3Q1gi9p/V4YrSaQ2QjLMM5lgYQ
lAASOQ7F0zKVzJWTuQuHgXi58FOBYcZxIOZlr03GR7MQ06D/GupklKB0Lv5QGA7E
gvPkxrMzUEDF6e1bUVycNo1gK6OjesTiaBUpqREpe4epbM/5RVF1ARmbvFd8taAc
o2lgi2+NazyO0fgg8eBcNdUKcf1nTxaGNcCSAu/yEuqXyHOd8tSwYtbF9rH+yKwx
hdg3BkTUCF1V+LwrKn7XVYVJAnTKAWCg0rYS1SyfBpaAz/DeDQp3GnTp/l2YBNhe
nAhrlTAMOx5XfW8iXUtm91C6utLYQDDycs29rhjyari22AAxxRJrHK7poioicHEe
cVuRG0tPPDZgOTw739RPlrgp5BbLXSj9QwcngwU5DJUyUNHIw//WgAhn38VOjWnB
eXmvxz9s2zLjEzEOj+Jjnm3TP+R28QiPT0wi9ld9kQ/3SCm3jUJvr0fTaiZtjefN
d+Cub8pvZoS35SGwZg+POUG0SPTBvR5k0TZ4QlKPcJ+fpP3jYjRyy2siGMXZq4qj
t+xc0SKgws28+C0KRmwL8IZ4Au4Wf5N7lArVLcPXVVwNi7zYdBJb4Ra6xxhswpmf
dp14MhQzgpWbg36rlKPrmuqOqQixPnSnQTAA6/DCC/A5qXy9RDBSOx98HmZeHSDW
TatwXjZH/cd+HwKMnwDE5K45NCImbYbOZ5Ns0WKisd96E2vcWOK/vxCSq3r+HCiv
zTSPEtiHsMowTvGFA8QInXKFJzJz61LaZSljI9eqRsmlTUC+ktVi4DoYhJ/pJYJZ
YN+92fefsFvbO4T5T+mKKUWKwbJSaiZ34XCUBnW0KPZMcDrggyw8wdtufvsZ/XiS
c9cD08PRsxx9kddsAHQQSvY9RMFaupEPWevMSE51qcQ9gDj25fqTDyHgtHszrO76
q6DGxaB/X27CVIV3W8GGu1V4CfiefHB88lkonmo4FxhfuHMCc/9cUF4BLSCXLf3R
1L086I6qB1UKSC05Tyo7Fj+xFMU+0P9BYbqHflXMahjZlpT94GxfKS/z8c8aawZo
f34EunGZE3nnMoiV695e9NIN7WKD0CxBG4biCUrH8ZUvGLJ6XJbjywHqoyeG/THW
zqNfCPcNpmsawlMp42K6nmcBJJBLxA+aAjMdN4mRUJEa1JZSDySn6z/PdMdauu+F
m63ZCLNa3HkClE+2wzy8afbZaScW1fbAgcWhYwD/XM0A31b80S4PtzE7fnDSJyas
3xfjUF4loQDUL3kESf02lOYKq2tOfMu4FURE71QC2nJW1bzAV4N6Mr5r8id8T58F
yejbAjDCuw0K8BICeyOeuTgeCmY+ezh/gL6UliwdXOpFQTI+lf5QGeiCWesImuvs
r/6ndoT2UviN2tLgTUPr/FlT9Dc0s6BE21q40RhxLTfznemQdpdw6KnPQalyXYqq
bBfh5/nOgjfNaWIytPVO3OIOI0J+2UG9GkNPRSZJ0iT+9cJZXUJXgdj06mH9juLp
PIB8lNhIN2LsQWswAYdTAGQ/KFGDhn+EgpIt6wJ2fTUGKTf/2DhYbauUFaMAhrt7
Wm41JzNwWlW0WEWzeXkaEUUfNIaNfSES9Jfwe3RHb3lOK1a093ZAH+z3/PXcrfqN
3jjcrKm3Dmi4JLiTErAY+PsCWopP59jfDP/lYubVqgkBuamiGUUB/1cnEVesL2Qq
ipduT2PEWhVVm99TpNTcdDsZ9IUuGxw+KQHn4j35unI192M1ZG0besx3VLXsnvG4
PANQOvshl3j0Q7eHSdaXt75GJivolgPCxYvPlzdaAWO8W8f/hfBOSwSQKzlg+u3L
4IZO4tB+VueNcRmI0vAvz6/8UYkKv5gq3+E59f0zDR9W7ZWTkjj5S7z+NOWwQ5qZ
eVVeXr3p1+Ut+QKevBH+9UCh9U0MUyF/1Jhd17/dDTfXYYliZPHWGqei4qNz57Nj
+HLZMboEVRACYygdMZdNF8ljHyYvhb6SbTUMLxAXiomszs09/qRZ3bLRJKQcp3jg
kkR6ZVivygzLrv2i8/V46PAYv/mhmfnnsDP640Ls37paDNnUd2j8cSbrx58Xjar9
x0/N6Cksh+haDGRLkFCIoxQmr5tMfwWKQKzEsMh+GKhfS8t6sCwldArXa4/loRgZ
QDdr4eIFj+VUBCFQ2zaTeCkibu3WdLYpT6ZpfC+JUlQAKoIXKGurLDEBZWL3dxWw
4Zo4HzB7YST1yT47RFevYX5WurhOmTafw/Fbaiy5lOtha7G+kgAirTSftQdqpDmx
zJlOaHVKsNWZyipf0fmUbwFOMsdxqPs7yoKUdCKE4v8pMSEJ9Pfnkzg6vTLB7Az0
/qkfAn79jqg6VUgVk2pAsRrqp13rFCQK6Jh0F1TJf9PDB3JTEEXDPrGop2+QRdOq
1TQUr8bZ3PbksexIo7wgyUkXCr/PPg2/icA/hP7hfsNwWmGn2kVwN6vSqhbauyeZ
qjqen/kev/J7UHNPHrXvRd4ttVWwSPvD7GQupVRIWQ4cpICc9VV74LIc71SLo4Qm
A5ArDDwRCC4EtECPUakRfPpD7XaDNcCmkKeZeJN7u94d905RyRBW7Zn2iXWUnCNH
YDvZXq017LRjuNHlrqirt7ScfxEb2hr2k6mJskALqXxHS1vqfEv3RJbEtEVJlVxi
RpQwRrhVl2wz+hd9J0qU+4K/DKU4zQACAV9kbj++TimcH7cBpXeBa6stmDMyoA6/
KHl1p2xH2PTYM7GNPtGfJXdtNjxeDZ15OeWFlpw6EcP+dTM2nNtQENJU9/xEy6ha
Vynn3rWVCbGVMQ+2y3IaKCkcecO9qjs57vJtmRmNpswNxnqV9JjKQdLz+J9b5jxw
iL4ZwZUMsHAGqQn/tyLTZOe3kVYKN9M8kUBq4B6q4GXY6J6kcIibKlE/1alDXtQg
FWcBBu9n1rIM6L6CUi/6nIcO52N4zK5tYz5H/Kjq/SF9+etJYjx6AbaTz64xg5zV
z//DWV22aWR071mo0LAXrcV+malbO4tvYFIAhxs6NUZfg5Xcy9XG9h2WUZMpZKAK
32y0nOzF0t6+MfiOtcbkEcu7/57iv03OnqBMj3CA1uUchpbjVafaBxl9CD4iOu1I
wIJ+sYcTMVZYhvWXII8HQh4IpGL2FTKnmQiIvNMOXxSEfK+nVJKvDp2s0YkVWDq6
xaEGT/CurUew3/13MEV694dLQLYlPNBvFIyTOJZ/tlTDSj3U/29tiJGFfqTMCxtD
oF00IhbJLMO8+1ogub6zQ5Aoa1xdYSgmNvWerph6UiYQFwyuoW3NyHiya5twvU2S
5wh6mP0nQHKTdgpxSBYzxMR6YlZ1kYVPfEpMh6ejoj2EfvUfbfxnJ2d/zRLAcOEv
7Abf2xvU8/mQCivyiwJZ+plU8qjX13WEn0fyhs+N3e4p+z+LdLDP1vYo2ewdpmHf
UugHtro8i9JOVrqBOc+rWJc/iK1Z8gqy4/BRou/fYrtdMRVrOtymIMuXk6366qR5
ME1YDv1MNjn69MrSYz9XzJuiA2/9EeV2HHEh8W2nUCegRh4j2exELcB94/60uQ0R
YW/MMbT4C/aLH7tZ0te2EpZfF40y4I5xqrCi8Ofc+BYUE+pF2320srP4sNuF9L6s
ZkwXQuXtGfpz3lT23m95bPvwUUO7e23mAH2VyN9lTDo2NTPCzskSMoiHg1NtS4wc
cbRZhR6QV/9nl7kenGf23L0LT1gAHjywtTL0+AUjEEI0VCLX/mHH55eD+666ObkF
utRCNIMFvncFAlTRvl6D9StJGuGAQLryowalm6A/kl0q+iqQ4UyybJoBaA08r/Dp
kNAxQc16REXkRW15YVGUW2DA0/DLM+w3OPmkbgcrmvD1x2jRYra6IAaLb2RWtyzK
uWZoNKsSzXRuhUCnRzi6oBx744H7j9FYAWZEgpB+dUQMzIsnhXFsQsSyjnmJu5ep
03sBBk2kqTt5Ffrvm3y/JVYp0TZllYqeO8KWj8oytav2okzZoVzACOqjiz1yeXxl
FLF7UOPH//9L3vPaD7GWAwZZ4PrCnqTaUiVAPdj9zoTtVBGmG7QvqRcoMdnU1QBC
MgKI/qqVyFMtJEBRIx3GKx9YwmsNZtyhxtbrquu513zxK1od0Pnt/b+/KSY4nxIO
W5NYQ8zoGvjlwoyJhi6T6YHR0sf6/p71/ZCftNS1fL8s7iIntbM+4NQAyzDcDdXF
rw3w1lya1vTmW0+HpyRzu58r4Nm960FfBJZlapbnzrc2vzyx68uzNvRk1DuG8EF4
LxnQ3lrKcV44oDPXqMMizZvmQaVrSzvYhNWDvodIVERr92q41sfHLFh+xpj+MACh
RuqJOnIjVPGpAgYaTpLDNQvM4d4aYSgLBjlmlPXnIA7Wk6AqhcG2+GLRxVxBUXCN
r9kOB2tzbXgLKgBH2XAKqBW0zyfV4W9oOT3EJIz1YFv1vBa7279rDys42o+lLSDo
nwsh6RJLei2AnQC1e1mRnOl6Or9RXKdKYxZaD6LvS+mawN9ApH2sYGF9dlDFm5LZ
8uGNlzC8nUxrlyFAXVu6V5d+HilRDRqJAUaAklMQJZeZXHTX1ONJB4Fdz1pYXcFB
ROJlQ+kF3UMr17uyqEhx6jfJJM0RHa3noaZWYwHOwvku5oVl8GSSnPp6U4sfLL2N
pGA/1DS54Y517wZ21d6eAZGe2LOFvMXq1a+U2QvDOHbd6kwVYulbcsgLB8IJKshl
mcZi3KZTlcnGEnVqX320iNecHWNO/Op7OrWZXZuVPDEZle0MToc+F9dQ/pqTmec0
lKkOgGgbA9f/n8Y3eh/+YJE6kHJ1cpz6HMRQw/MtWczgz4AR+/9iKFnPsiAsN7ey
3UueXk+wRiiBgX6/6S8FBN/0DA5ZH7IEh7d7Eb4Y7Y/C7tmXWlnH2mpDGZKcSRIE
qnFayHmNLCK6Ni/ddxbFNj8RKS1+z6eC7oXdxzsjmTwU9fcOpJPZD84z4vPZ2U7l
m2DdnPhgHf6ZnnPx2Tm31Ui/KRgIO6iIqGVi3HzPA6y6HMhwjCNU8/X/MecQj4Dm
aMzPX6FnScDMRejlMAjc7kodBRXU+cDrb6NK6aa7buWAGtcdp7TO6bAM+74GvYOS
jl537gGhIAhcm08GXD1wmFY1/rPEAd88dRZ9kDfHbiQ1WRLOazUR/5V9kcP+3Ga7
FGZtc8gtnDtrWgVndO5oNYKsC+O8YhHT3LGZDKzttiCHxWEePp/4cc/KYZeVjCyE
BeBa0RRru7ypDqHxtlGY0DcS39EsxzlliLo6ZTu3v/UtIGeJIJnYqTFQG57L8Yss
6uP8rK01mxmI6d+XveR9HG6C5EAi6gIpViO9vG52L15XQw5OUuK0pA8yB9ugijCf
1O2Gdtevu+afTFkmFB1sbw93DELVOeP6qYvHzMsVmw5Q0N5ldnNDiZNIuHK6f4Fx
46TqCWrS7mNqJjCoAc7xtGWeFPxDTabxXKF2kvfLaVWleqzzCP4IDv8gsbFqBgtm
YsabQkgHDRrtYUyduOa4u4cKH4pM5pZaXQ/7aE9ljJegN1kcXuRWB5xig98xTmdg
eqPgOcpYvdfWMpy0FvGuNRYtc0jWu6zGhCeV4Xi8evqG2/rQu/uJ/gfMr//gp3kF
0WT82Eh+3jsSFDAFjLhvRpsrBKZ9O4LusMFyUmRHGQqobEJcmFKzSRqU+Blpk2UZ
Tflo7qYMPgG9AsJ6ddM2wumjbtforgSEXjYbZ/Sn8yTcntu9PULD4hiWIThL4dSD
Ba5RBeGX3wYgADCrFPklDwjVKGhnxmL8ugSGZswCOcdAZC+f2fbJCeMPvOa6wira
afAEOiUrv+W/MJTqwjyyzzNn5zOZFWQ+InJU6ZZWQnf2X0DRQhD8q3wce/UB5W5D
ixSsW+VVS4FSN2M3kC2UkbZpgczghFFjuPu2NelM2dupXDzbD0gCqRagfuisSF1a
PP0+fTqvEswlE4JRoSq8EBIfmEP2u3/HdylWeMBxFMRiXa+aH7Zek0lw3T3vRiqk
LyGfQlZKybOguRLq/HbF8rPIM1Nr38XIbJGUKlrOPRK5RXL2YB6zGVAJuGlL2vxp
40cpd2pJPzudKfppBjKUefH5xYal2HiaPElzcuPX18djeRueNhmcwk0MY1f8CVu2
07uGDHSA09hnSniHZmN3vYgUTpGf8BJ2XxEy6Ev6aifsfTBfznU560vmFkNfjRZH
iP+86uXUfjQeom6AZe+UhGo0KyQzDEFqf5B+G7GUSz/SyPX2dPmggEflj2BntKub

//pragma protect end_data_block
//pragma protect digest_block
lmsDAhqxUqCUev7YBwPtl5nue+c=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/4DREz5RggQfKwqmCWpWTBP2sR8AKyOoOPHDMOnj+lv94x+JliFTojUuhbWdThMN
4ZmKiq+U6ETij4bqnXa0h2ncO787eMrOXiaFZY2QZZdSQwT+0i9u2tyBIbA2Jw2+
3VA9GEunHfW5sqbIEPifP2DePaRPUMYxx6Y43vkne5HXICu0+ZvSsQ==
//pragma protect end_key_block
//pragma protect digest_block
tICW83LuEPIDHeOAhYuP4g0uKAg=
//pragma protect end_digest_block
//pragma protect data_block
r4dtHRrdBaINWt5YQyHD2l5lRwpbjltedPDfOek8uVbXE6/deUmvDHzwsUstc+/R
AGRDas3zHoRmJy5ZqKUgAK4t0e+mU4JrAkIv5AX5hLkDPUCAZBQPYjm2HSG6NIAO
fSKpTLdKES9JheIvQB6d3i/QYzYpVuWZ9AOd22uXGTWJp3ggMizJUV+xAF/uMdUr
IBrrfKtarVIdKvRXNQE/cKHgiJbcXp/UUV8yKOkRC6JVxV5Y2RCnw7N7Y/jX8DNl
jUWg49HO/ateQG5zQrRnJOaVH4h2awSXex1wMEV285pAPkMKbIKnJ1K6mvvQ2PkD
jNsHHvgzwQpDmkmaMk1XMtXcFD7mWpLiXtiBVxIgd3VOkgVp+mh9vGUQwPzNEswc
6tTYijWhKMKm9xn+OYAE2qnENQM3uZ/3Pi8jr4QypXTct1iwpwzK9zyXYfHN2gLJ

//pragma protect end_data_block
//pragma protect digest_block
ojva4afK91MhroT1iyqd221qews=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
qgoQEnQ1oO/JBKs+Rxf2MEM5PMCuCUqNMPz0mjEeJ15U4QviXd+gXd9qZIDMnTZ7
8q0077xRR93mPEtOtwIsjBJtMvkGr7P1Ln3f84LmrLtSEKzH+WVua3IC818OQS0Q
1yECrafhhvllXDwny7y6aNLT7qSNPK3uuVJEB6y3g55VuS1E0Rpb5g==
//pragma protect end_key_block
//pragma protect digest_block
eFynIsuX+LXsoE2IAj6rofOU6HQ=
//pragma protect end_digest_block
//pragma protect data_block
4/SZQwADuUwFIAh7nmo2ard8mKVJfkw9SS1U1aMwPtcnhEWNiaIgHahWbLU9mC0Q
id30hzBNDDobBiclblvCfu74PW3f6BrUXBjIec5YQfM8koPHsRTm84ybbYUejVU2
luGRfZau5HJ/apuVTZbZdAJuFsO6N7ZxJ6CPe5PSYhOrezuHCfbjN9lwqSnEtYLH
0MapqvJIIUczNk2stamon6NPTpnBUzieT34DroHnAo5lUFEE0rfPNPQnwY40DKDY
prHgLrx8is9jPRMHqSp3OXtxZ+T8MG0790cv8usCBITVsLCPRKMM3JwDb1LixFSu
yGZKlI0xPKou2sPQJtk7d0omf6/7OQHJFU8XXawCYXwLlzEKnKVv6i1tLnfFLLRv
Nd1nG2TPPzFU9MjQx7p8Qk0wz14i2p2EMK5Nid5McausraTNRpj1t+xT0QX1E1pN
9AVMwWX9/w/nAJ72xB6PEY4htzIGznZN2fIwA82ndA5nBq+4EPlM+5kScCPXkEDF
UX/R7enmXRqnckTLRxKxhzXvZGD52SRa/o5gIb7UNugD4+nQtipTJMOPbHkUujOX
FSQKcokpuHAXTBxLgwNYnygv+0ytoOI0KlajGYTA6dTKYt6FMfVQ9rJ5OiZ9Xj8P
SGYHpZndGpmsjw1OGP8vEomVvx+oLkNAxOIBMAbYB0k4c9lyUkpDJDRTVkOZayUd
AM+bZ4ghQ4WJwon/FH6f7MAtyhuiHGo/xH1JShje+t7ZkBcUIW1mZKUvdk9V7S6U
tNk7+lK64YQ328kxvV/5olvZIblsedOr1d50cG4FLfev59/VMUXJUVoNEGH3dZxQ
XF3z4+8qvhrblBJsGNsH+TM1taa6rkK20iM37bP1RsYwmFgZxYt+FMOpPGsQ+gKm
b/AcTETKopDkHkMwejvejQGObmXwe4d9I4r66Bmvi6QcOgVmmoDgt1u4IcDIG3IH
ILbAXFS5EFC9rVsiROQF/mwi6AEYt+Kn7NRbS9vQYSINwI4ws/MwFkdpEgEUHCnS
wr+659t06PyRffn8pBDaGvRpetMW7Ay9J2FzygpA9rLLUNNbuBQ+r2R0c+DwBSgq
p08Lfa74DzDRwkNENjPO2iAvffiOs1Gd7q4b3gitEErhhoSwak2unV1XP2KFQaYE
xdDwdIi621lL65TmOtUTlSBtHJc1ojsUuadOgYZNaFkj3GMaxpEPRlnoiuowVUGi
y1qCR2gE+t0iKjTMLsgew5bacZGKwXxSP8ga+SXYFCmHWxQUN3R/GXfoVGC0Ksjk
yyTK2N0n9P9OclcMsOBsDa2eP/ap3iHME8xnWj+iMLYG9Lb85ioHBkAOO/CamAiR
ncrO/ts1SbJUkU8niMp4NvfPf0FMcLAJ53rcyqXeI3K/LGrHCfoulXnNFny+pZaS
Tvn0PeDsNU3xkfOyolgs1Np4zFx8nwfUvGAXf5UOWNAp0msJy+zDgWcyo3PnwHuE
fNpPxZS06PYgxOwxaMBGgzM7MxutYLNmV855hQFtPQh5rbZd0j2Rb/V4l43SsM3T
cNSVr1Zr5NOFaffIHGwgQN7Hwn6Kv2AAiJLXjk2mDualN3WcMxsjoNIHkCpWHeb8
y7nY3/66Xsk0mCunrVNjsC6/+3IlaUMQ8cf9F2zzKniDEdr2OsWCRKM8J3jUoFYH
ZLEj8yh0kb+63w9FRt4tTyVtKY0ieibIA9oiNFtaMNZ1DHdUt9yk8II9zscoavjc
OeXec3Ja8tMeWvaYYo28BioQkCSBwhTOB6IpgB82Y6NRXoE0AJz51Aon5HG3QG9a
5uen5jesXSvkaCX8ol5d6CHbxja03Qi1hkng9bOs6vArEFPn4+QN0w4YnMp/Mob/
tPu7nOzyhnrr5yiupHli8S+UFdsb0VrprElZXYliqlo/ff8w/72gyrJztYVhT+h9
Dl4LZRkFMJ5nGCng5mXsTAahNFWQE9daLVfZGxiv1nEckwE8o+MC+3O/2p3MjoJr
E1jE24+FQv5guLDugaTQr6H/9q1r5EqZFdpJL6jMvn9Q+I4ww6juAcZP7j4kfNn8
siNi8BnjTluaIsnP9g4SYcX5qrRk8G2L3eEfD9xktjlriJAd3/CZPrbmxqOW2Fmh
UyY7zri2C313eZ5d4p+nWaW+cxeclyqMQJJwrP+v37YAFMCmftux7Ovi4tCrgHQH
cqVoHC7FjfHQk24pSf7PmmPSZoJHK6XziC2TmYxTPcoxpEnMVrvbL4APcDn7WfIs
yDuMhCSjG1atYuXZVIjQxmtMB3sj1vxJ00c/jkYqnsMd7mUhHUUV44RXx+lU6XWb
Rbs1nBScvDBt/C5qmPom5R3fwOMfZHmXhiMnSubGhabDN3LURqZqvr0AEzFopM+O
B6W9PCwnFvED7mJ80B7knFpdtLjkD/3PECvEA4HM2HzeKJtYjzt1zKtkDvD/l1n5
GrgHOmdufyn+y56gd8OnTxBNfeIcn3sgEUQKuhJ0Q7ekcaYD6TmFWsftvSgfNpJh
HlknSlNDxMwdd25FLarXwNjtjLjrG+Njo66aigcnz6f8K5vzAZKj8LRempJXxa55
XkqI8t+3Ps/dJu9c598zBW+CDTtYrP1xmXd4FojPoMODnXYdy4wgQLVvJq+2+liI
+lHh629iUpGtoDI2G9F+gEhIQVcax4FoZd0jqYs4OBbv2LE6plygh+qQiP0Spu+2
4nGJb6VpMQRMze9MUpn5EW6OE9wnjDdvmKtaCkkr3XhB8ptTFFDWEBjJqPf9SUYD
1TqPNJh0sMDXfMq39ge0TIOdF5rUUgZo6f/LhV4ryZqE//pK8JzZpxTWLBsZll0V
RzpI1zXyxEL7fwYXvsfPudOy8dgd+Ll0tEcP9vU9apylchvQ4EsmfjslU7WbZdhq
SF8adOQyEZKOYXvRcUIkvt6IrvWKVVDMFRTamkHldLiDQUPyKOM0m2C8TyGMZ0B4
r3DsVSxH4yjVOfXciNfxj1MkOJFqvlQle90Lz5tZamcYSNo1ugdLbgd4m0VUu/nT
iuccghAs0Lr7pGOdJ2RkzbIZojGP81YHECM1qnzr8RltcR/miPVDvHV9erDuYynf
U33eZy3+FVYfprATlln8ygVif72DsI1R3g0W4ZNMRaULd3VkhtI7+AOQUvbJM60W
AOxhXf0zkLJqgE0/0OC55YWoXBLk3dP2KVnqQP3W8eWmTptkAh4oxbn4N50yNHLa
+A3HVgw6TSQ4XyGtxRSRsJ3jHErlq9955afnlO31UfpH8+qqZi4JW/Vg2ZuEp/Ws
JE4iUZDGMxMFLRALhN9KSnk2d036pIuJefXaveVTi3lOFXvEk0Si9iJIYVuL+ViQ
OX9/tSIXllG6jGN0wkh1M93RE5ybi6mjrtdhJmPa2Lg9OEUF25y3aK3+NgeELQpg
oIhGa1NpAlEewduWFqvhhS96r5aYNUPcI3Wi8h3yavlU4hXYDcqFKA0xKOpd3cYa
E2ktGTZ2rIzgzBQ1BWzWcsTYmmEePiyX1JG9pSASeh3ltl1bon+KVxD7Dzpm1IML
g03ZwrllqF44JEP+roa2KIMh3Fs+23mFXGuRBSSGnahHQzsW8BIGeD+W/0hGW0db
pQrbZezpzkxbROfupGz1INtgFD52HbiA3jmHwV6K5uqeCRflbkiFIAtKkFlBUyZy
N7SVDfaDooZcRk7ccyZBT40xxuqsUy4EKBGyOvlEc497FtbZpgF6h9OezFzeDefu
zp9HFJqdjyWnMELB7hyQuagG1QHcGzRdzuPTyUjuh3oicz887HGehah8b3gcfTVJ
yfmmX/zff6zwOA/YbKsKbeKQMxxlB6Amz6Udv26XcIvXbZsZ0vz2AP/mRE9YZ/jh
HbkXjsHyM6zdhWWbzA9MTBshjdCLEIwTKgpVyOGo30vlwrfFup1EHtzCL7lW8Z0U
gTZ5fj51l6AEHbJIvdTx0gWiIfFGs2+N1GywlASQ35ZZ1+xs6au7r2svk9sJvLOG
VIqVACvKihed2HiU0ZlNxnPF0lO0JSDz39FqHRGcqD/My/1cN2XGV8SzFhb9nXbq
3iwwy9u2XgolCZRNImfk56CSnPs9rM8NLvn450vCPW9vauY6urJKZ2KUa+l5HdvU
JesRPiyM1ItPeUfCwBE4MHAjbmPewI7UPxRoYhrLl8lYSh0GDuj8EJ9/ua+GH/TI
La3/sAFhE3E0aGB1L2lMb2Kv+mwpG5HcA7GOCxaf/WezHM6F7W23Q0sUjtKJZimG
JGVFw1eA3WXMj0NOI4BS7PHLry+JWYCiZK7sni5M9+tce8dOjV3+aLv89dChvl8+
Wry+hudSsLthSEEQy5hHmVbyv4SEFLwiCDKX+s9xyV0ZL2UgyNgwMk43Kk9U+u/G
XjqgPFU9Z9gnaJ8LEgQ6cM9qro8IU3xkXyPeXMpRwcM+w1FhgLGbrtG2mw1ai1iq
b4CU4SOnWx7aHRl+11oB3K4Y+CwBAxWmSABmUCwrtk1y1nDLN7uOXUM1+8V2opyT
js0neyBgmBT3P0mgIMK/Na7Pt62v3ieQV8J/AjDxBOs78QLZPnXlyxrS8ssMNk0Y
p5cBODPuA+122Sp2Bsy1CsS92egO5C3F4riplZmyfTOY3VcL5FzM555/gkdcesab
rzSL8XD2Q+wr9+4VFRUyNJNbF6T/iyyWMaDAsKRFQz4zLoNIOrH0Jmg12m1pVz9A
FFSOS63k3Q7kiI67K5LEpFqddQk8Ey4bZJ3O2GxDyMootK57AWrhavXF/nvKhHKn
1nNWr3PED2bGiQ9gDEs39+vfwPyrFqJ6ilnzPB2blv0=
//pragma protect end_data_block
//pragma protect digest_block
dd5lVgvrM2zw51wysKRhLDrzy+M=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
JM/h5Z6D7b5mc969wa0mfMH9FjLmL7GNIIOBbSnFtskwCb+RdwCbc8tsD6SZagpr
7tSg5jZgDtyNH0ICZvDFu+WbTUFassp/v+/lXzuULAaS3Q2FharxGIs2RhiaUo6S
5K6yM7BCzbCUAhNiPGVY/SDeTWZbnle2xnPp9LSY7aX16UofWr5dyw==
//pragma protect end_key_block
//pragma protect digest_block
HWnK/rMQQts+oUD369ibq5rrySY=
//pragma protect end_digest_block
//pragma protect data_block
bh8F4n0x/W37HzykYDnIDWKKAPdbaJSeQl+9NKfrjvbL5xRY5t8RrPsbd5/4kabm
/OgVrThTf8cmwvavYDXh6c7dbBKACHx8/kCwOfhBrmFoMdyeLV/mdvGBdcQES6Fq
BL1MA/6ftHU765QKMfHvUapW5jvwFDJzX/+CkcKMLU0uXFIcNcPLNA/xOw2afzlA
AA+GsAh/Ki7KJsl0k7UxrHvNq3pysgj0VNJAPzwct1Y0Sui2QTL3TFrqoe/UafSN
wBe7kHLhKU3c00V0a9KJXiHFt7sN7mD7/kB37X1PyMbTn8B00Z3LTfj1jZMkM1Vq
2JKaPOPGo3CCglOaUDX9fg5SuwChTOTMNX7sYNWp2zBmn3CE2G0hcjLR3BEjpu+N
ZPV0p1hTdnhYfYzLy4ztEWiZzdfpVO2oK91wUvqqRM8yo7tsNEkkgPAYE/Dmx3+S
SWSZRHXF8NaIGqv7kCmOt8mS4XVws8jjj9tmmbYmpwM=
//pragma protect end_data_block
//pragma protect digest_block
0B1m/0rTbMBleL3mrSuByfoTQgs=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
A1eUSIGblLMit8VSpKjXEDZC7W3VGIt913ehKTWPWS+27asyVq7HOHNkbBgZazpn
IpFBVcE6KJ88UFOJikoLH9YIArYg6j424VC8PgHo938gM/IsNBze2msdBdIMsjCe
RqspXz8Fm5jhVE/Jx8h6CcFar/R7S8YKWxlmaPzuGaf2fQ2qW5zUVw==
//pragma protect end_key_block
//pragma protect digest_block
PNHcflbTqTv6dBId+L5lcUirXAM=
//pragma protect end_digest_block
//pragma protect data_block
42amr9RMH+dwEZOMx8yLzzQoqAo0pR2R0uTNZzrDWaiNkZMORuI03vXdjs5JniL/
D1JTZYQ/ZRLNCVgHF7YSrPTHLRS8o8h2k9BFwyDnwV2dQTqD9uVlJ9Uw81cH7pNU
aksfgPrPQxk+1ezJJ+crWi1+iJlh1VWKM7fA02T8fpJ5YHFtmuA4BQV+4UCftoSX
FjFeBbN5yJ1qOM14MOyyWQGLEBAX58EOr/K56jkV9qhWbxXgUDtS9Qco3XlGygpH
ziULxw9jNZ7j9IvBsYSdCLsIkavUB980X2WO/bltnlO3aje63eQ1UAklfkw2aQTu
aIKVWtUtDD4eH9pylMyiZtodUsaeXgK77BreU0Pdk5tmNSVeBZclOy2vlJjlVnYq
IMhBEFfhp6u8dSvyWtBp2B11Y4t9vJbcDh4r8MyWa6yUlMvRFA3uGzHhzXZasYFI
N9VtiDauMy+RFGW5Z7eQl4jo3AWK3wHHjYHQOEfGGnDV3fiWgLYa9AdlhpRP05CQ
6VQkh41k+x8A1zqdd9iuMaQuQWrN6tivZE2kLQxbGL2ovjMUATeEkcBRLGgno+7j
OjH148XjT0eqPjooZ6FotlboU+1WvkbIdZoCBqLT4gNjLhgG+7kvoEKpegsbLOck
ELhCOa0YPtghtF+IXpMmNcL+bviYOP0Q1lRBBfggC+5NoKAEC0bOqTWYX4UjSEWr
91r2ONo1c96fEXD6iSl7EZd+jQKG+mYOrZB2Lb02LM7BeLZHCMyCDNQ9e7lrCemW
4PSV+iwK4lCoOrevGGwUJjmV+5etZPNO3w7fMQtjaV2TgpR0yLUAD1/ldfqrOfTt
2sxB1EdXOCP+LgK5vR/+1KXWOY1T2Cemez30KTwajG9bNw7RACF69Q3OcxOW/XBw
0zbve2AqokFV3Azlw+MBMPd5I1AOZ97a0+9ysyczbwhcRQfc5PEHxpqNEsETjD67
TUBUPVLf3r4B3pQabN4sq9vgE/yzJPlfAdVahbR6uZjGlsqO3M1qQIgTkPIFouDt
Ox2c+6xL8bsHr0bMkcHvUfATQRu9/m4Btv7SfAa3H+EFyqCjydn3bIgbaTQYQy6F
u13ZIu37z7TXqeg7BmG7KiHJ6D3x6yCsW7XSyDNXOVc8Iw59STYE4aqpyvo9lj9r
7Eh49d3dmhWrkw+S2vX+moL4rgFWF0BmMm0cf05UDCUTqOL6sBrS8p5KyVq300y7
UgrFz43eHIU3puRPGDQkEXrVH7Lj5BX9i+JxMqYsd9LCqJTepa+eyHR7H/quMx5F
CrnUEBx+5zoiwRaienwTsy8i6Kt1s68LADFeu2fn3p9U6tTjrhyuAhHEcjQ7U1S1
MeWFWE3O40Jt+KwWTI55JMqS6B0+2jW8+43HN7+ZhYv8v0E9DiQtxJNJCBHagra4
qpLkGkldLipWBXTgxKMIU5r099Qh67203Cq04j2dna4Vrkvl4p7IZIGR/bPeZlde
3HJsmjEfnKQoupLt1s3/4m3IRSqYooDmDDlRBwa5/lXR/o7QtxRa5forFfde6vKD
GX8DnBCiwKN6kHIPpPW0H8Rj1X8axfsGGP0x63l2h3fVbsYSoTKwWaA/w8sfEhlZ
T2OWM4jr92iUYp4obgbrT7EgUzPs/YgmpehRPygmP+1HomQlTrxJogqjeQ+TDjIE
KjvG7qwKvnGTtTpnQ+Ran97ttvAaE9bX48hxDXkXQ+zmFgfnLNlT2PAollYZLZgU
7RaWmlQBn/O/M0gckJ+TyeFLjftPByUwsUndfXBIJtcPHmec5+pm0Rb8pTn0cev9
XmfA9QZdaN3bFUCbv2IMdhWfKJEE8o7wH2B3PvbnFiGP8f04lXRDyseXzLpteAOv
xXSZlb4ROXdBtaJVZdVqA2ZZ4uqRHNdVSS6bmHwAu9fbw1TjeEJ6Q4ALLQsvvbFx
Gqz6A/FPD7oT3eqDMG4Bjxz0n8uGCXbuyTxwFkCjeU2ZdjcjJ/Ht8ipQOaL2YM1y
K09tGlaIVD0DPjzon4SwgiNUkvst4uhpD0b5ZMMItEvjpdyay05iVFrujTcHCzhw
hEITWtptnZ4wRbzqSUreoo6/tW4eyerkt5Cu/K8hHW272fsf951Kqt5ux/0NKtne
D6J/4ybsNcaa0IuoYcZuZgNuqmCdN5C8dewaE0Xujn4rdgs3Q2L0qwiixfgHSaxP
ViLqk3x0T9yk2+VeTHvuN6C5bSFQxHkgAo5MIci0jMaukmySVnJTEZR1hwjTmzsj
eC5o1TQ8bRO29vCYUnpmafoj1yabyKlR2/1D21ziKNYywqmgNjmFoo8/dRrThZAn
WjLywJ+M/6jlZr7YFV/NfeRJUfXBunBkelbUIg9TGT8wAcFlYiV4DTpGuDq8kPr1
D62N/6xW0e1/BdpIPUweAuudkuYh2ETs3iSoVCtvNBpop/XtE5bBQWT+7g17Km2s
44fhN0lucggqtdeuwhkZZE1k0DphSBA9aeoA/0BTVxljy42OGh2p7M3V/ImO0xvE
ZouoAUImkpD7iVKl/dugeVYYTssrastVvaCeCdT/e6fUktTy+DMPteypfajw9i3j
RVMGG6fBvP/JQlmq53NSLKw+JkSxyeuPAtpCIHhebTHHLSEMXOEa7BG6/rCM+y21
WoiNrh+vNk/fXAUZ9rLRdkBjdxm6BNFT26zJpxWJAThyAQkz9bN/16OQq/eQ0H/i
ryus6pZnt+9P1CmvxgL81DlZq5uvNlsducrwz5QD/iKVf/5JYfWBv2sG29Hy3fra
jCtYPNKLpje3fhqY+X6otAnGpkPps6Rb363rUedzKZvq5A2yxBCCI4zUdR2nory2
WHZ/KpL2jquTzyrMJQz+NE1FpSlIzrG6esXvdiRFcOW0OwvYeFAaR8+uRTGptCID
vHWqYxL92+ODv/9Z6fBGg4kKjA4QztuF5fC94V5D/OFz6WzVGhfc0avOUggYPEoC
RzTSOjqgxX56QHfzxrZmxoC7ZQ/PajLkhhUaDvKNHD/1k/p/T4pW/upg7zXJGe2f
CmPoClQWu4fD8/1aD92IjkFxD35gFgUTW2iw84s9QlUoS7LZWh3MO5/bhtDyV+Wz
sOiqf9ijDmYodDU2CaT9/FGLOEsEcAAGxHK85q5sjfgJE2lPChf5+6syqEmCjkoY
54CCcTy2A9T5LMiKalN78VwLVigXWl23dlEpmY02r6zV5CMMvJmnrNxkv2Jml/Qn
V5EKgkByzQ3aAwR3zUps55qMayempi7WlljIEVog3A7ktkeDXbwGp+eT2gT6QcxC
22uE+MBxa176uiWTFPi+atQXoWxabRbLolxzD3qnZ8Bqb/p2Tn5pEnh63mdmAbnF
8oq5CZX6/tnhj6m9kfdQ11SJc92G3vfUcV0PkdTAqSlxEVHwYdQk1Rf+5g5+RQL+
tvk3rjl2Ndue0xWI9NqQc8RGXXv/X3eu/L324CSv9U5zv/fKWfRsBTTq+Y1a5enn
ATIVwNUqrUEoxlTbQmm1VyfBk8alCPCf2y4V0Y9I3IRZua/dKX9nAEKsONPm/plD
0i4eOoxoHO2kBCWmscdbr2iAPj51EQLas2aGmUC+5jjZuuz8zjYjroUtRToRsMtK
2CBdpFvqHJLe60OE09lphEblAQhh+jAy6UaKDC1o0lesQ2oNiZvhcM07R6ZjHMTE
R+Bkih7X/9q7YTmkztyBWfORx4m8HdRdCKKge7jQ9Gf3sklAeid9cLZyipJXDTGo
X7kAhsSD6i7PK8fCyWcwxqZDYvPMG5yC4wvpq4C5YoiT683Gtx0YzCYqOoqt9EwY
d1FVfDKowUjYEurA3A6FgmlZT5dUMN942OPMATjE/uJ79/wmrG2HkG1SlzuU93V+
HQMcEE/IC07oEo8Wj9hYlUpd4vBNakqtNtMCeSNrny24++O35lO2F+R6Fw1P5rNJ
tJe5J8N++1xrcacxUltWZtB0ihcqsaTRc24+Ty/8+B01lOJTVTIYkiun12L5Rc8u
vKBAi+y5Be4ybTrqBIRWgv7eIXrq/dwi1PITGlvTKn6lvgkeDrkpjEiiew1NppAd
x19o4uVLEsOHkMazPc9Ahk0YBopHmKEOccTVbzkJaQvH/MKFBvoElFRoxj9ROcWp
995MK+8CrL2he26f1E1kBuloJisQszwvxo5CVO54jqcgxtz2G8xJ3cP5IvJMKsTw
dmNg2q5XAPGvpQuzi2UWwmSm6U4bKU8y2qn1XuERVqmrv1hXB96hpZJeaDIy6yWN
BtzkOwe5fCszn4wQQKymYG3JVziS2ZdJWe0xYOdJfvLhkTP6eibTdVWEkiJStw9V
r+hRIf8l4nC2Mc+MY0J9aZqNVl7z3xqA9136zck3Murh3AaF5q/F4/d1nqJfeWQg
YEEbgiL2FdCiYjdVkYJWXTEtBlxOjQByd4BXLKHo65Wmos2hv6olci1SDl33HECS
FCQBcZ92T1iPMwSu7O3TnJVgsE0a4W2bwztSYbZrLYoiQeJf8wXUQGK51eulUYgG
LnK/q+T6FZJobqFQywp4YRgw/7jB6Zv+tjPrTefR+Jk4QqeOBIfiqmbfCQft6jM7
txUv+CvXxKP16zslNsXHlxaMxH07Zx/cAEjPfCNjyiKJ+Xiz0oLUI8Oqyd9gLpAk
uGYMR46F7sWBXxWD+wHvXCCHtZX0mfSrIw5eFuOz6Stgx3Ut1JaJM5RjwOKG+GEx
yIokszWuEfWLE97zi0dEOu0SIRPedwvQ03thjwZqAARsKFRDv3ctBVt9FDYgAGA+
AMGdGslkZz8y8EAaYMa7QOGE4bMApSvlO2o4ajx8T+9AoYl5rXQe4YB+dEmrotgi
0ULMzg1fjGrPLcK0aQjjvg4uAzIDZx8H06gCyo89PxM8g98U8MKD1FEcDAP9qKk3
DpwVBpJuMdfIIZ23qZQXvoBwrtAVNElw+pGRsm0eihBiytAo601fGvAjoDDOKN2I
QFDQh9FM7g8yloCUTvGslaqZF98K4MgeieMjX4qBWil0xyhVmx/bVKHbQ9oWSy2p
R363jNQPnx87NrMztgUnXJc5nQ7P/LP9jpiLZ0PLe4CW0XsAGd0R7cJTfpn+RqJY
cXL2530Y5njPSsxmkaDMj3XYEXo/Nuq39oK8SdPVaPfLlNwrJnecgH1j0p73fMtP
Q2XgQ8i7oi92x45i3UZhJmgBLgd7mZcg3rdNV62X5N3UhB0LIUPZ7R+OK1pFe0ty
HRuX6b7fkAOMG2EZpAr1oBaRdcKFj3ykTwJYTnNGjXEpE1NSq3RMgRWozwnQlZnr
WMlo09NS5OP5KFByA2sejFvT8usjRud92ddCHOCshDPghINemMRkoDmx7O0FzZ9D
YHET5m1kXtrIg5wom2dZ7rxdhEedlozTZWv/mDVAA2/vqPe8owNbLr/4p2R6VUyg
vbk7jVzPXt3enOBExXEbAXTW6NKIHH48I/h2+yu0B0KdRZaA1L0tDSVoJf4Zx8Ap
sBmmEoCFPSm8j2KCktKWz/+kJVnA8t25YVKrjWEUbf8g0a4GBhYUm9ALHAm7mDps
YZw1AlSUFabJ4FVVLAN1gsq9mh98UhIveVZ9sOmApgC/eazHI+xpOIOy0E4jwcbQ
jcs9N1PKj9w3fsEE/HZZkkPFLHkkwM5snwo0YPqHwY03F+6tki3hdtqbGqhmzkoU
TRxHn5jS43U0HdSHttf1SsLj0Xw9h0Z0O7wIVHAV/hxpbj2FnkuKAVd98NhjQfBu
eVE8h0XM23JGCa5Y/eKEMOm7yHYm/3SkYviByUvzsQKWfClqaximyFyWz7zb/RFc
Rrsu5IsxVIhE0k3oWyVDFC472L3GwuWzgrMFz5MPZjEBGWUCusbVCRzcu3FBbyyc
TF3RgeH5iJOIIRHJq/l5+w4OqXtWof4B2JA8BsIc4dBiX3+/PVd96Hr00DxFHKbp
zEi4uMMsO0ryy3KuniWC0CFCB2nyiwBnQPltFZYJw4Off4OBPZmSx/upzBaZBwCG
l4sJxhFZHRMFKe9ZdYEzJBMcbGbXjWDh2mzXtwo0znFXXGov8z66/5a4GYQQC4Sx
vKKw2m7aMgRK5/RCFVkYmAFFQCIZ37MEHGZBrtRadypPmJqz6brAu09E8w6+Ck5j
uXe/AfleDLpgQzBg0LebG73vSwCl0luTSLnBaLy3D7O9RkdmOwH9AcAu2vqMI7cB
PCg0y8jjFfO5L5H6xQuMegPqW/S3EBhGDEGH2wOHb366iB2wah3n01curc8fRvKV
svNckmLGJOGFqOahUsz3Ryro4qchNmOdl5LHLgcBOpa2WrSjMC2JTvDyLbNVPTtc
o80Pvxnn50DeCKc31X98Cefgzun9VY7tFiTGvqJBDphcYSfHm5KdmEguzhfCxp3b
t9tiBGBunNkba6v/TbV3wrzR7bRlWiO/GppY9s3q/qft8z811TggZAXY3eOGoZf1
TsOXHnqK/ZLCZXF9QcTslDLpdcVwUhSYHCpPNH0du5qiOL5EqGZ2HbRe/NPnO9v6
C61g8e8fzJWWmPh4umdOuKFZBQZSZsQjnSAGjfhulwBsPC6o2G9O3CRbbcNVJVoS
/blNP2IRkFB2uBKXjsO3c6/n7Q+vJlOBUDE1rpafPa8VkawzmOJNvCLjDc6Bg+Ns
3/3B0tfFBY2dMQ3aAObbjgmPBtCuWF7OkIGtEZNXiqZzRMsHwYVpF9p0VaYxQrtg
xSp7ve9f0CRh2QUJWKa2m7rJEKCJXevQNnEJsMO0evYTGqQ/QxtFTyb2nZZZm/Sv
rvT9nxDApGaOWuzMDjW6lzs19IpuRg2XOlyxK684DBcKYx5bK8pyL4fIWZKPbKWZ
k3BkL12dfGGL58gai6kep/ZGl2/VnqB9uUN/lfBoscCsuZyodkp5TnHM/IHX/9kl
Xlevc85hIUR4GUU2dGd1MDVuJgUok1UB7Vw5a8GlV6OBA9BNEWmdHVCLagtD49Qf
D72qe4ckcgIIKQF6XJcvP0OFvyiyBgNeM+FfonF04Kvyf5HshksPu/OIyRB9HVfi
12IpzAoeykBiM9MS1JtweSBpyeMnhFo01mgSN98kXnNlpAcY3R4lwqQgQoKjrO2v
KjvO6LfkD3B+Sqf0oIJ9Q+2fIC3nbQmMj+PAW/wgm5n92NqIQ5byFP6KcODLlFfP
uQWXbWqogTDXAsw/pPRd8Ug7G2wDshkc7DEFxFv0r0YHfSPg8hWURqd1QkWxpH17
sGJGGy1YZKZy6cZ96hYI8AN7fFvPNYv1rxsPqCdxQvOXp5F/LCO8M+YWYjizCS2j
Rz6DFk1qqfvbQECL0zidotDviNYSifyw18JYwKE5sOPAhmyjR+17CyRC22Ofw/vF
AeGkHzIiXw39bvZ7VUqzLpL6/WC0tJPk6mDtBos8O2UtRfIJ6ygz2K7Xm+oc0IFG
lJTuvVhaQNFhzxjk3zdXYx10+x2JnQ/uobBHhTqQI34ldGbNOxjCg6TjtlUbi+mt
b+AGOn/7GhSfYftmpa5PhPU3UIiZqZMdyZYxHNM7sgfIosVSZp0sopuIFmD4YgDG
nLEL64p92luBc1J4viXt7LAWdJmo7MasOEF0c7Yhp1Llv1IT+Ijb3DmLhYlaLEId
ydpw/AmCQ0x469Y3yBURadXuiAtVF/vTRRvyL1JowRa1I2Aj3RdLjiBzgHf2GCmA
A1dzQqNQR53jt53IMUSyrT/2fpLXUCRZwBygqsqkH9CyHeEeT41Ew0t+ev0kDAu9
+f5Scd9335xrg73DRGdlXpDtRnMW8gl0m6YhyRXFdT1NWbGdVPbtlqKD51YKt7Zi
PZvjI4r4M5Y6ILIFb72wfHcVYNAN7KWgI11RxTenAC0PQpmZJ8Hzhl22D2Wzgs3s
O1T8Du9wwiquQZsnXMXOMbrQ2nCt+TVCQmphNJdjeaL4p0z0jPhLFEorAc3D2mmc
ZlC6+WNBe0yuyGucdMlz+GJ+OmO/7bN47M3dVpKhQf78IPGbiN6zifH3OzLqI+bE
VEUA6zFhqQtVrfx/1yqvn9X66yXUjzJsH2O5rLpouVpqWMRLNnAw2fMTR4U7W2Aa
sMA55kIemkek/xK7pFoqF3kQvQWYPtQQAUZREump5QMMSlK+mgVCnp55Q2cKMSMW
8VcCiXkvXmJPvv8ZFMsp2NDBlGkJYSnhPk4qWZcgjKrNvhP0GAcYrf7rTAYw/zaE
7W5zw+WFoZqpx9fVQOuPRgPQhYMssE5Rlj0I/NNMOmNJuGqenOFDhtWseGvO8MBI
1jlXE6vQYWO/lM5pHoXnJGJ0WXHpbR6GjRFk2I+06RT4rouciA7R62+ckgUm8RaX
wrEf/OfHrC7K5PTD43CBRKXCORevo2tX3JfNfnXs0S4wv7YP6DiP9fEEWgYh6HqC
ggMcrXw+tO0TW/zwFF9hpkxKkPhYkw2rP0NgkT9dj08NvwF2O3rX8kYzwLukPjNr
jertt5YwZIvMp+HbLpmCL3XdorTpoZe2WMTS+N0JjKw4/QMH2pzGHEINsljyLIWD
KPEZi8EzYjC0b00uXEWVV2aPaqtlVHXj3WrWmEOX1Q4XJS9uZWl0fAtzf8qj14uv
bFX01hBunBbgd7rimb3kXIfGYNE3cJIff3GEFlR66d77NHjCzzv+cPUaQDalSCW7
Pz8IZ23NJB5u10TwdO6zpXJJn01X/4/OKnDClf+Su1/HAyDxWyJ4lKbCNpBvQgwb
aoCqQLG/pbYIRhwCIEeWKQTUDXkwkZj0cniZYq12/A3i5M98f36ojGn6DbB1U6g2
qhpGeK4BRjfVQTrIH7IPlUibA4Vdz3X5flSHpEj4fT3XfDlfXXaDJOwTOenCeUuB
dp008yT1MnzldLkbNUT5txt5aBCDqRX7FgJP5KvZfE5XF1a93HWtFA5vpUhREwG4
e0kNiyLyU5Gpmav5R9fvejIdPN8JNf4+DXnGr0A7eZNrw7ptPxbR+01Nld/nrHGq
unh/tEGTz5x7A/8KoGgTbNlHqlTKL6MmDccoteQJ4Qaq6xsHUKGcHATOCTpUZ3O/
PC9Kcq6p/2Vro+ntEzW8M3YOkeiz7ryGdn5E2h9olL/VpLxG4eFr2olJdkIly1/p
vYzLy2r1B3zQREHhr6SqFmT+sq6Jbf3TQhX360A8p2X0PZAbWaQzHHnIfI5UTV0X
3lE+hEbQAGIaOI1QwOjQ9z687azGbgXHCJtkPqoarIVFi3yLIGRVuKfSy3oaLH7z
9eoR/XJ8QabT0E/pCBPEwRZ3TngC3UoP1cz3qLQS0pfZ5zoY2kD6MoxshUOVZwbC
sj3R+cFuOEqkAaUDC9zwTHSILD6SrOrIYkcuqcJHwjiOlZQSws9LwPHDaDVTYRt0
aa1YWwHXOjDQL+1KN60TDA6BUplVRUJRe2/U+0u07QDCKkAJMwhDdlE+yeu2wezD
19gB6o3hVDXURRDctvYb62uVfNVMGGL7S39JyXKzaXmw9+HdC//HQ3e4flDyGm2Z
oUmJS74LIK1T8w6RBsjmaG4Yvi4wK6vxt3i8pAHVAco3c/9wV1lfjFWxEFWI50UT
qWdTC+4JV+irLg0XR/jcfKNQ0nkOMIJOxblfafprGxyeZlWevhrblKUqt0bq1/Ca
KTVQAnHfN2gxnk6uU7HHFanfrQ4O08vpqynmXamjtk9nZihWrZh/c3PMmQvh6G/E
oODpdLbxubeLxacs1g7KZwp548q37P/obO21Fzgme/yg7ek9jN2J6rWQcne0kZtB
nRq52OyA06V55dkYywV4PxTL6HNWmI6z41U8Lj7ykpMIMz/Ic4Yruq8S5Nzcwl93
6rrIbmLyORcCwsCbJ8Nu6VCCwJ02OkxUlY0yU06LARSEQvk64cZiOayT6BFLGr0Z
aK/SxYPALWwJK1Uy39BUp82ii6974NzDofvTr/EeMHNg2+Yrn5C09JK7asdyfYKB
GRaIgh+uSq46D//EDbsp/EziXu+I5tut9Y+Jlzc2rMQonMnZmsC+BDuxRmmXZnDY
BaOLn7EbP04z6G17NLbuVgs4SRNVCtKLMieh/NCrDKooVwTh2zhYMAdXA40PE2UD
n5guJ+BaWDNRosDDxSmtFAQvEYFHCmwDXMurjKZtGEYoffEPgX22Eh719R1u19JZ
LWf/uS1sEHdaknFYJ1qdrR//soccLbgrs9SG3Fw/28aPzMwq/RfhCcT3beSeEccD
SjFeDvPWYJd4mWVZk8BT4IvU9DjWWvnDdl8qIy+Ul/I8a+x+5UiyugpuvK/t+EKb
MOTTbs0RoJ/XocdcLbFTc4Zi49E9txtJcHoizcKjdJPTpSF3FT9EiAa8cnQqj6Kx
DC7GQGFAwJF5f86aSNF+ScuU7nduegWpQuD0Wvo50KgC6swCvkTv0he/KELn/q1x
sNa9lOD9Hk+g2rnXED09//Wi9ijRnE+P3K/PGBaDBFx8GP+HQS38yTJ0o7v4PdUJ
1J3+PDCn+HHD8nFdmvTzmvTXs2a5+jCIPA8TDi4Vv+Zab8Ek9c9MapDQ7aOWsdUH
lzS1IRIMeDmE3fxZoeD/vxDXwro8tkHAHLAjbSfVQP4tPFQhrVY4jIcZ1+Rm76TM
akrwz33r7NLmBDtgGPz/P6Pshd08Y4lXMeaRxwGl4YLD4sKkRaL3Mj3/CySAgted
oNuc+OAOvcCPstYf0bWmBfFftQ0cc69xyl4yIH1mO/VkelAUOav0pGHmLrkotyZs
MZT4Sh7Fj36enQcAfrYFdwO7eCioEU+t+/YOIQZM7GCT3Sj1Ph3AOM3Wm6jnOB0/
jpPBc0eWEAoXBolrMf88520BeMiCBy7MevtQLcwu6+kdzSvKt+xYbmWKwWbuqj5T
OPPxkAgEzVMgxQEEzlrCt+SCW1y9A19hi/x6DQ4mikJppPcjEmbwvaIV8s0zLtsI
dICNwFnjRYxIdKhL0qGqP7QLhWVZC3aFjr4K5BS1i4eaS8/6w2b+cUOki9R+HmJe
n9YFwoGiEnpMhqnc4poaa1dRP+GEKMsGhiJIHBfZFhcg773xYxVYvYYOoLM+6kPW
SN8w7MJ/KucfJxhrYcwTvHdNiM2QMt6QWV/p1T896avnHxF2F9XeikD07p8B1Asa
nw+CxDG3kwfqp0qtf6LO6wpCrfsAGxqaQDesyNFVrJPskXDaUgM02QMwVkZ2Lfb8
u39tTUMi79rAOGEjQBjMfVuXNFCQx8hjlL3b3aykTReQY821QbvG/LTKvdUgvOc0
cNC+ad5yjJI4Ej7+sfZfEx9amK6zqiTQz3VCX+8F1Efp9/TBjwQi9VD0UiTdR2RV
WYx0hCb67oet40FkkuJfJgTrzWz+xHXyNp/QGhaP1kb0dVveyPJ9YrqXqfa3Rqs9
yJY6kbyolprNk6mw4ClSK+NjNty6Cv+DZ1TpjG22IlQuFHqjLY7Hfa9CRsubUyTI
wkKp8i8+LT96G6wrBPePAry4cO7TjrqTwkjYjbSfPjvUdm1o4BkdpGL1vGYXkkfn
AOpJnh6vvKyDYDh7OQ/x7Ummfh5Hs6GDL29nHX9Gqu0yZlVxbri32xEilIyfI7pc
2ptBrrOaifVczXvJsj5UsK7DxZW3l34Nbpd8KOm7JJW4T2ilp3z+nIJMZ6la9b39
3xpvT/GU5C5JWcngL9W2p6n/i21TVQMHIWZ8SsbtzPALpJxyalaNTwa5n0gTdutI
KOXpBYK8TdftPLMfoSetGUPL9LWOoqqCG83nmypoWvxKgiPUKHe3aXcvA1jArnEe
nRVHi2tllNFmjIvk2r9qZHiktWF3Jetjd/l/bhVbXZ7feRQZGXtq8y/uJ7BLyqCi
KyDNvPBC7nrHt1eAyCXotOglHiTQf6i88+c/fYzGioHppz8TT46+bYn1iYcwCPSg
XBYBI+9ghYfLYEfsF3ZTwSQfoT/TMR3cismUhIysWxcvV1kttZsBOurkq7FJ6kK2
hzC7rKo6yNHWL12CfmJt8ii+I/Y9bTHe+iC12lEpmSjz1JR+Eo6LOuJEFU7RooXR
LmbSAtJvaixas7grxI038DPvThK/hMlcThWwCQJpf3RoxKCPkX7Ch+srEpIN5SSa
gPjcZgDZ3OPEzccbNNHKXH/8GWJ+Ssij5XLX7q0NKNyQaOL0Tq4lUtjCwHQF2fg6
owkRrkm1AJK8L+6ARsAtteSu04XgAOCV27DXmyMEA3vnnc2y5KAcMqUUyuSAZCx+
Ajpo2p50YELJvXxHfYkd/NY4zluJsxVIZBYuFA74FU87RdyTN472gp/+FQ9XTOfV
Qcgq5xIQ22Oxl7Er5o+Lupn49zXKuQSXCcxboasz00UoDPm/ykl57v8tXywbkk/c
wuD/OweRT5y4XNz/lG7eYB6UynXyFy3QZzWX+bjlNKrvHSJFoLXb5Zg+UQWqz2je
QCBqhNVzqI7dEuRUeUwoJmewBoE7fKnHJw174Pv32daWbMjIhIQCfnuZ2OU9Xxz2
EEcAs/tZmFGhbRDyTX3YROlKRohJtkF3w18wSsQscEVs5WwfitSlVBgPkJiWC2Um
7bOwO6xNqQaW+VYv9/Ar3SjdFJAW2e8rhtENfUT1VV4knOkJIifLw+aIsnln7zVa
Zpx3UzGIW4XzXeAxGO9SRBcBiBzRlsLZ6qM2HdF3Zc3MQMNuGAj6pEHxdYU3eotV
3O+D0LI35lyz2+hebEqZbpCQkKk1Tf/u1VwS5WUuZKUpxL8KbNv39ErHPT92Ou1b
mZAOsqedLlUwxC/3usjNjfHYKAtprfaLMEgi46adtqqiGkEuG53Hq3PMsRMlbTa6
Lqw2rBklJKvhILfZnpZalPPwbv7YiydxwxmbBOgca7lNoykCx36reuhj2lmeNm0N
YmhwKTkeVZvZ0udxJ0uRNu5saqokNV43TXzQw0JJMqHjUVuONSkYdK4WIHyF/2dh
JQjD2ASZ/dcv1LZ1iOUsvXf0EpxAFPj2PNDuKyNPLcOg3om5hYE2acAd9Ti4niEy
AG+8dogQyqX3BXEL53BFnJEkmjQyIXCWAAZBXWKuz54eOJIK6w/C3eCgQDmXjARz
ulEMWwNF+Mng7XKYuewOJ08lSRMzW8K3F8t2FpELIR4W49lLOJPSjs+wVhFz21ud
ujd2UJxNUq+5e7V9JhAFk1X6He0NqhJE3qHP9C45eDuAn32OqRDqwBeLxc55tiIU
XM3lSmuaVY7rRS6yNVco9xAnApNhpXy1iN04WJTDpKwg4NAbBEejqUL8XLs4tguT
y3y43y2idBjskL1pWX536bTJk5dth1h/+3evcCeAz4S+Hqnv75iZVHA97F0ijuCQ
YYYF86yewkBAc6SEjyudFdwhbN1yprFNTAiLEekVbSteV2iVgkzno5GMKSxjeQRT
XBl+k4/TBCZmBWUAcDx/XGORoFcdrhIwV7EhxkjR4WBzJvGi9ued7ehannWeCVBF
Api/INep2cES0fRdOJxhnCVTe+f6xJP4G4Z9A6iFmhSgXzHMoG5vbzNNy+bGQjDy
pBnfBxqi1+XMCWlEX3k8PftQJs59irbMvlt0az0K5Jshs7N9PPRxw7zoVfl2cecb
UwNFkZVxuQhxfPQkUOdVrDjtWtGWZnaO29Fii7N9oi2i6DmTb7YoztT3+lHlq641
9ZY/VRsDJXtxvZ61gDc46f8S+s/Rv2CRncwrKvdu5Afb2qsnBIMbxrUcD/VSGTpQ
LeorU/YR2a6ParyP6s3Vj+/ya0jWvdHOuLrRFWd9gJpIjKsMuEhLRvLByhCCm4UI
xm09UAjO0x9G+sRmnt5h/d/Am5thTHGWledUhbKRgr3aViqlq7dckNNY5R56mNs6
LYYo+NKINpPYCY9Mhfo3YfTKpGQM3RqC2U3y23tXdgQu4CGxb41QM0Kxayr1uUVM
mMBXbVFcNWRoufMXd4mGkoCQLy46ZUDebXpyWs2MBJG2v4AGjFtlFcVSDDTi6xCC
VkiJHSiY0L47m3SfH/HpLZPCsuUlWsxjV6ZXP3BaLhDIFZKXcHnrst2oHuKIhn+8
RIo4bpTSMet3RhrNGrE5Q1vJMKFsMDcXXjI//yJBUdzOAaAygApgrhqeNWURXEoc
D8nOJp2f0seZBlkq7KowcnSPjk5rRgIPa+nI2CB2Y57NWhWrW6PhK0NIw6QsopKX
J6WASJA9q/e+4yE5yo+vl2p1cusQKsa2UpLUSwh/l7gCNSkaizEDfqLolZBL1T1M
yKWmV+Uh2RtdgP6E9FYUe/ILD3aKmMIha38JaAFOs8kEeZZns01oWJCehVr0rbkd
S0v1J0yWP7WqasED431ecISdlvnQ/VZpOORDGY+bPVSfg/6Tbf/OjCLktoSpbvYS
NLoWEIZJ9iv9nyfDObYEMLwced/DF0SgthF3CLwEpF+AMVhfMmhdeF/tPdoBwD3r
yUrCgMzCUQUqN4hXaXh3G3u4DWZ5lOwVJ0OqONKYJH94sJlPU4Ks1p8TCKhZvLBL
oakAnDmHYrzNR/e2qB+t70GwKAeyZYRS84jQ8ub+0KdAKnM2wshTbd+itzslx187
HPw+ITUhRr/UTCBx1/y8dlehWlohdHxWGdO+SLBlMVPKd9yvXPi3W8HRpW4YCw2Y
/uAvc+iOndsGJVXVxAeTEGSERZUEzeN1q1qGXaw7mUygnLPAz6fYrs6xCJmvz/XN
+7e4tLH+BnM5z8gjB1JOzx1sqHxvBE6kVrxgn5Z42mweCv8g5x8ZJfnMQBe9e9w1
fKPZWQTAj7fK2HxGwIyiemvfD58JTsJviWRlzNlbLDXKeiPdfafchV3E+ttiustA
jHv44mGj6HENuFcARODqmdWYXJ6+UCbmCLMJb40DFvDG7OAPr02IrfxlSi+fRdTY
3nXxMCBSTT4qCw+LtHMpK3rHQMrni3mo0nJ+tHU15mBwAGadhuN7WhiEzvX6L+K1
oy2IUmwLLLtHjKvokQzeC1ZbVCQ8Y0goRmJsjaqJUxytO/nQq39cn9b/feggnKPe
a7HLG9SoPmy5owBQUQcr2qMpdmHENSjUGzcTnzxPjq/VX3XuuBP4gqEOvCGWbAP4
QMCeVReztsKTIkCHq5jXdr3qH16EFzLc7iLHCqqiQrGppEdhq4xJzMk0Dq13W9ND
ejt4O6WaWb6sRr5E3FoWGKwsu15w3K+uuGshOdrMUBS+IriSJUQ3ORCTqQLYGvHB
8ZWOfT6dKftVRMKbzT50n1nC5NoFAZn9D8fvaHUmkXiHT6bS9ND+L2VQZy87rNzN
TnWRySN+5iQku82kS6DmKk/1OBC1/r8MWRzBNzwXUBE6CDLYZjEsfRcE21wmhL0o
9qBUvlkheXQlazXo2/JHJD7qro2sxflq4T5PKXJONqilUSte0SCIbEiLmkK5XfSQ
U1h3NPK1Izy5VPe6O80ZqMmL4pefVcIoYU1hwpLQY451f0EX+A5xRIqSC6eDe81m
BCU/EGMmauhXJdHIf8UPybiPlkf+aJ6M+Rl0R4KArG9KmaUdzI6PF2ogNVIkxoJu
4JO6EsEG4gmtxL1egkSpYbDd5sgG3A+cTelaxrvDnzOEvr3KwnmGQfipzlwCl48E
IdcC7HYyGK5jOvI6fX2nfUbfS8MP6Qc5DlUbs264O9m1IwbkW+iODGLEbWXHmm5d
6R3HbC8QMDM3A6VuCU+sOtLGfFrIxfG0mY7aEhfmzaCOWCrR2svCf5yh/Ti9Eefr
ud5iUg9W7NoWU2OaoFZrUHaUuEWuWCfTm3PBt7Za3t9xdmKIlEgVHRfjS5xu7S7G
zxB9gzN/BC4FiAst+VKwPUo0Cae+xh2hL8IN317qmaydMuIkCkWG93f5u+FUKT+5
FgOBN95Zjxvza0gxLlIU8YIKm8fVPtXshE6/3Tfgp2YIace4XCpmywjqJBByCGQZ
sNC0Za01canhAefAFhe6iXbJdlOqMb/d2spIJC47wh0Mak8Y234hosLfH17+ZlMZ
7fjWuZzh82sRMG6LZisBUlRDAEjtYhZGyXlod7UCrFg1jpxQb8VGW7a1Xr183PLJ
A+7789r4Py104j+z/RM430ydgEcDYukY9raTkZGpb8IEct+ZdOjTCSCXZPdKbaJN
zGFHNrv4BTmz+ilho4ozODGYGt5Q/uYzx183V6jwVCsC6pX3dXEWvnr7mZcLbGiO
J40K6ZmGZjD8WAbK2k1W9SD0j2DvKJjrwM8EP9zRjFkc3yLt/VjMbh7DgFeG49No
KnCKICK78+pdaYfVkyGHZMKPoU5IIWnTMVsYa5UcSY28mgdJlI6qi4ifCaGyph0M
xCqZh/I1G3EfcsHx3oWGd9qQ1OVIBTYSN0jmd/t8qSYU53E044G7KsGn9l8DsU31
2an5romL1LtEKv+X7fDp4dI91x+SyPaZbHeYYEoWvYogOEjI98ZjhLEE2JGC+Gxi
VMlKnoRs2qsbm20CadCuM0XTD5UM9hyZzy4GmJTG5cwNdF+lZkYUSHBQ7KQseOFT
aiSbqaJFDrz/gQl4M8rlG0EryFj+dMGtajXH2YFERBbgq4lzJZ7oK29onngH3vc5
2QqN1Lb2Gns12Hwxksc/or/YeOVsocFQkYneM53JQMHOP0r0ONvR5AS98Xb3cbI9
H+qrznmyQdbW6lpaRbfQs76rkrqRdC/MqrG8zL+kG02hmDv7nyBDxG1dLpGwxE+e
g9cT4YsruSUjPbBTAZ2aE/qCvHVQKAaUyqb/RbLGaIJ/5cLvz1SnCNfyaslmDSLT
aQyFYjZBIWyG8Kg2Gg7Kzx3G/OEjcUuFKz87xlqBbvTb6/J0SCDgAaeZyYaActbu
6B7JHcbbyE2Dskw7YxGEayMKAiQIxqFmYUZXNd1oNDvRaqsvDrOBqsIFmjSgsdse
12ZTav7AwdyuImWCW7OLSuYuMsYVk+s2tMwtd0bXN/mcpLxAimr2kJX9uGTJe+BZ
1kNMExDpmj3hlbk3y+szASUeOCgBUrdnIId1DOs5ywoECCx/oy/yT1XlpBcZYj77
jXzowA9PAAfd+oK7KOsK/RSW2YfU8KyjSZ7paKJYuNoP0nch1HZnHxH5ILFu6geX
kKcvh11LW5pMc0sfhQOjISFsySEVipXVIc3kYipNSXR+lmJkNOdtxbdKd2Qm7M9j
/wj0gNP5y/cK9lMlBfHa1jlCdJ/OfXR5vVjN77UZKamcjORGZsMJjGDOAV1VFbRp
6FVQCWT+Ia0Ax7yAvtkSGk/ZQTxIBYJYIzzIECYutI1kSLP8d1x0dCFCfRAvlt2v
2xuJ38XdPLc43mfY8ALNc7TNhO28BhgWZAozLfLu6A/Nc8wyFZpFRHAwkREMeB5J
a4rtbe9pDtAKOPFcoWD7q+OeZYMiDCAixqB8NCDSPUUAA8UYL0TTCpRPYFCE9m8u
kAtzx9uvWxnNtyj3C4hKMZ2UjMzXKoeMVocI35TDUWKya34mtHyk1eJEOGPvma49
IyUxS3eusMd91AVvw3GxU1gqqtaZ0HUCIdp8YJVSSRv1AUARoK1/jJ3f3WrNrvMP
DyBemKIP9+t9XrWJaRY+bPRkjGP3ucbWJGp+TYELX9vGEnUQjlySBIX2Iy5YR9nY
4MwfQpHukgpSNoXIhvpW8koMgYek91UdMRZVb5FfN86SF6FW89swo6/O4It0PFN8
USJ7Xajx++QS8wrzqIEIuzf4diqrKNyUe/flsxQP0DHCyU4/LD6dDVZeeb93qTks
UZybkyajSf1JTmJRCHaP+wBpF7+rCJPN56J6vKWvkjx4BAtpnGL0/O2u+cB135G3
IMrq3QhIKfg6heDcluF4ZiWUdKC6nw3S+g1aSTB+XTXh7CN5xfNZxC1FRTfEua5m
RDOBAw6PCJRlQR/4gyOvsCfPh56p4Qx8KyjTI9oUKPAoDAfDFsftU69bfg5V813A
tHExbJnW69ToYxAKMwWlDLMEaYlkrow4ph1zOnjIPnvXscQJtxdu7Zi2G6yuvnYL
vpHWZShGjszS4ArjTKSUp0qaVfvH3SM5zLgb/I22YpJ9UnOChOnD3PUL5cwTR+1g
NE1INfyFi3+IF72sCPZOClqN+b+UR50Uft8QD2GEKnJZhC1bfdSNYyEp+RGqycIF
83yVaArUDf5iZOEPKBjm9dD7gAw6DMbsCMjs9Z6LMIkoVqkPGuwK9ONQGNTG0CvO
2Rxg4QgbDjNDWxJBf7/6ulTY0M3qoEQbDhM0M6I98mnT0s/oCnj4icH48oPtm8sR
CtD6IgqszXsXqzqVrOMHsPgmxrFtksITaY+EjpetVI9pZkti/F8tSLnlWTJpGZSU
Ds3encOnFc93Hz+1YlZsL+XRMj4St4/fV+RjtBFizuSivZ6C1ewolTTQhX4DHKkZ
akV1s65JyU0AgKt1A/hVuVJ3TNOfIvPcXhLMC3Q5Pb0ybEosRDeHd9sTlqmsOxos
tfirPW/93VQZRxCwn387vYg+TIXX85oKQcMVAXzAXNc7c4N9K10evp142ABewckc
Th+ZMYNHi0+DwLTczeo4d4HM/O2QD+aopLMjkusrFPL2WK56U8I6yKhCdfR7NTKf
RUYA8+RUAKlNodaGtwVJGCGPPEAYmC8ab040vljiYdvYmtyq8o4vQTjTdBcyzwAj
nCCrBFrai9tfSz/2kzvQXclF2lNXsaeZqilByNot0yuGpDXpbdL3KAnUJRousGaV
ZpE+I196Ko72P/dDZOretX6drlw0wEMZ3JqzFfd6ke6jEPUbrOFRd9EWhAUdjHoQ
V9oeicRqDGqSDX2xnii3Kn4H+sUxlHM0gQAj8QsdOqLRaupWNjlCOaQIxTdjtWDi
IU+LARajO/br0+1lGXIGsMVYCc2hBEz/HHHPho4/kpydkH/Rs85mhwTcwgDGEYBR
rIV6rxbH7P3BsrzcUMWOc17pA6T1p0or7dNKF7dRamsaM1PhPnlyVh2toh1A/MUW
oeu5RHWfBAmFsS8of3UoUDje0rd3qdh7crQYjwd3pHT1WUCAZ9oMevRuIXgcsjV0
s6vsrrBJU2kJjG6EbCheUCatbQs1f6W++GPNe9aqBjomRTsPOl/8rtJRWmNO1Zlq
YpAxJSoHYfAOkIztGQR0JLkQbmZsMDoUqpVRZ7gjgnAqBy7C7vZlLq/QlB5C0qFq
YxIS4byQ82fUkb9azzEzNkP5fA1+7DNsW2RjwL9HGjMYGNuKwBCETNEwbMKtQFL5
RHySWicHYuWGPtt8cWrlICZdGgfkotDrDgDDSiEHsi9QTzhOPwoM+MbDnNzNR7uK
sacmamPTifNS6FZyfz6xYtlKdoOFjhnVfXlq2SCuaIJ5jHHxRrwEhhoBC4YpiyT4
RLiFzeeZx2ZrUg5nQE1TEGvkuf7lNjQIfjmHN276TRQZn8NTKZlOkAr3YPBUAFFV
iIOgcVUm29BmQHOqxSPeNnFsbRkmTHRBMfGLtapdN8EkkLbbNwsSgpILwhstmTfl
FZT46wgqP6UjS6c8hlyiFYWgUbzxjCVxEhjRig9X/SUTxfipx60bvQCvPvCcyUSj
5RmVaX5c/IMvssZ2QT6kdfY5rb+q6SkX2MweQmPiBwTLBXhXH5i8d/eb8zMdBWgF
nYMHDZH3WpikUS2+9Jn5yfr+MJ3rDlOIW+sX32gldHkISr8q1zCz6wAn0iWmBlIS
hlA23G2OpW7oFobCZj1zsWb9uVDqgJ/lyCqyc4jwbhUoSf2ErL6M5L911ob2q8Hu
zzr0gppO8qYe5gaFZUabKwqj1yKVZ5tv+mD1KpS7nawTGjpMV2GJCotXlorVjmPl
sWaPFiTmIzpqPnLYh40bnu7ayCLbi3fZyeTqwvB++TQy+Ju6SjU2cpB1okg9mC/S
Lj+wRpUuVsg+DBCLbx/5bGlQGomzuP94umEhN8gTQYmxq9eW1AikgO/a/fVMsqSx
yIiUwFTU7WlpYS6StCrRbpG1Tq77OccfUz08ScEAMp5do6aXAlpG3vRxyTk5zp3d
FB/liebwbqoKvolb2i69eRplf6JbAfQziqaWHptqA0bFlDOCtIGUx3szfevRySOP
YemHcXbwZfoC/lYRk6oipwZ5jSI5WGaaltj5w8vItOWsPuxUXWW9/izwsGHV1cUb
PV2XTHxdaeOkiTyfaZNYrhEiFZe6SrvHI6O5tsNqbEPvbhBQGV7GBk3nKpPMlOuh
u11NZD8MFkXIPPCEQovm4Q4L6OryZVMFmC98K5uiBEUXCnlLDcOsY8ibuMwj62nY
/9Dvzt+8bpVqL+WijDv2tV2f1Scbj23a3Q5fM0J6RLPtZNk/ANoVvHFULPMomy/F
OsVngqAkFZ5KHvsCL8TYJgnaRuN7vO7EEZ2otih0GRT50gFITX3Jb9zq4TCmcJQ/
E0Vi1V7s8jpG6PPtqprPqXP4sET5ss6xQDsm3d6dnVFXNKw7EVNbOe59yJ0C5N/+
pqCXIu0Uk54QHawQm1lZYW2aBOjX2Of3MU914G2MHK3OuGCCcUWZCVwmfOw5Ddit
0nK3uRwnF+/3bZUWM2MH6Vh7itiVJ88arYPvS8+dbb5tYLg92H8boKbKjllE/eIf
CQ3BfT5zCmP/aqvnx4yzAK1YZrQLSBHAsZbYv2EpLvunWFvXqPb4ytwhrkfRwIo0
tuBnkB5dndOAuF6k6WHQi/igWisLugG7tH0eJ8UVCrCKnLX306QqqLGB58GTP6CU
Sw5tiSPkT5gT4S/b6N9BbhgGylAVw5vulQPfSC2fvrDTFRkATouUQePit8QxZQLM
e4PDzSD+HavDvgBbuSEfWw98g6jQ765Z0sWcMzYjLKn6/BwW3qDemL2XYdrrRY+Z
yyo+fBwnZihCwQ8x7496h/WgrgIWbic2i+ijxvQCbsNXXcnxo2/NyTwBDm9aoprn
vSRPIcBFkhYRn2RJ0S5w2S6va1+ZiEQcAXbvc+ntjAT9jjgGAJ5lRCPqo9MFOYAb
/StBbn7IUG25MZCgkyc192mQJGgdJ2Fpm/AhtvdGuD25BZBjrSKrWbZtEMAkTwLO
fsufrlvgAD+Y1/j1vRQg82ur43Tt4E25FlOHLlY3szXh3SmyX8CAdvC6HCznMzkj
0A9xbwQPooLbRQTTfYZQ6DXVep+Vd56+viki2c0wobUlKRoRHNbfZ8sJP07V81yr
Hkf7uvyXIImX0Oen1sBjPH47+FbuaTlUaoVG0T6XnF3zmJiJn6Qz5qgRCsGQ+u9N
spVoeeXZrZcgkWNxHXoYKpnq96xAZdMer5v2ViIetENsP0CNdjN8bGN0P0Opj9u1
iapD5FOSHmkk2XmqEs5ocuVHuP8btWLNZvvM2lyA71G7wVYGwDxL2NuhU1GFHNxn
MrWwupR9yakoyvh2En259jRG6JDAxb2kUNwti59QSNUeU835+9j1T4momHYXX6Jd
JmxaC65L1d9Sh8a1Xach56yOa86zRlkllJXi8ew8RYpQ4mm6iJ+5WWL6YMxSxie7
0RTBMjCK7EzbOyOyFAKRnq7gJJAIst1ELw6qZfoFOik9VSMydjrHXfQHVcf2yMX8
MZetK/7uCRAzeyE2JN8/bsSohRqF3gjdeLiuI5TIv6aTWXU4GeWqa/kDRbaGMhaI
4KsCliMYqZvbcSYMEAqK/qPBt7X/eIzZc9RJOfdqT9QSp58PgwABu9kI+LJS33An
i0HN3p3Vdz73sFM+fwTiXoXmlIiEohsW1+WhiCK9McOK2YHesLZ2ESnA5hrk1cQd
1onL+mjHtSgR7xTkunk+HDLhRMf4vDwTn+MD1+0obHRRjE8I04sNDBCwVF2L2Vmc
y1JNO4HGEHMMkALnPExMVWUSKF9GZDDmWMX09tcGf+4QZeg+vRuxNpteVnZBa/M+
T4+dNyycUzu6Ji2wW1y9Pi6EnQAfZOberEs2/2IsBa6PVB9GPkQgCJLgM68M5m2F
H8QgjRCRati8sjpe+nlaxoCJ67BCyFRdgnMXtqHDeRLeFln+tBAv7zPC6aYU+1p9
ZB2UkNWlDOgr8JCYdx8cxZNjgYWzAs8ZVs7QG7/mvdKj6jxGaobv1tblWHhwygBi
P0aN7k/5T/Luzblcpv+mGLMoPoc0ci9/2xlwdXGmtfxIHpUXuzeRtCaGl1YqXhZN
8s9xxkc54+EQRjieP7TzvScgaqaiyu3sMPwKm47mNfWVmMMx7muw9jE+h98xXKS1
mzfbDgkp3r5UBdDUg/HANWShdmn+PiDO8SCP22Ar6grMhS6D4LW66/FHYW0hd5Yb
3fdLgW9NZZsaCxuslCNIwG0bWb9zUI3OfTIZnqFndoWJqfR9M2qm+XQFh2zUY0Dr
d4dTa8FLWo5tcMZFhuoykI3yvHhe8uKq4LbDUcMT+X//VCrPk8YXW7eOQTEvguZc
yWhQ8CfWVo+Schc9JMBaE1e2BiAZkj+33GVIABaKAIAtsnQXZgau340U9oOoc2QQ
ML8DiN8joAq7zybIwG/mKvvSykNK89GvXBqeysjI0k4lNFcp/YqE25xfTCMVxlca
smIpgusKxYkN2cn/I3/gnSjZogReFyNdNSEvJO64B4mYp7NVZ9F2qJ3PSLAbn5gt
LsZQDBOAQXPNWEQcikRUWmh9tWgKSuCAXgbz5JUm1w5Rja2zN5+JfVOVz+4wfRHB
C1C/0SwSPR2shTHmo6Q1NeioYL1VgicSNWMR6An8bM2PkkF7WSUHmyj9OLNbKDtE
JGj4Db3QhSdPt/VRpbmHAGxHEYjzwgsxcrd8lROdsjNy5aAKvovXR2L3cZpsrUd+
jgnxa9dVwupirXZldnvgV2CLSXHSZmMdx5BNcCfMmIDtv/w5R7NHvNY2ESjSQDLj
6pQfHggoi0i0BQdAGQ+GwI13GhObzsKp6Jmey2te3SQ3HKn9KeQeLpuuIB+bMSd/
sp4jU//e8dESNocUkSBTBNH/iRZ4Wt419WiS0cM+pqMv4YA976VdeDOsKKUxuSR9
M464vJAho3AJ5LYca9UfxT1dKCRXIKYQc2/YcdjQazRh/DLCmYlY/OCKBYWU4bHl
jnvrJCu7eykKYHe9w5+reYqWYog71w2Jpzqvh4NTEg8IYS9mSu0nmm/3UQuk/f1K
nfuf8cH2RrcraLE1ygcaT3SdiMLk9fqDqNgMn5qJ2IfWYh6D+NlzzSNX23/pjKLB
UwMagAMc9swR9DxNcapCNKswgGGOdRdhX3KckhEMj5RP69tbpbytic9ABcP4mFdP
mLCjcNoLp4xqUoVQjn9xv/yLpDD5e59a7F7jkS83SbDtchyQRjkjlLQ0iqBA3umJ
+HWhu6UgoyFx6Xz55CneD0IquyspvQ3Z5XQmrbK3a4BG3aeynli8Q/4aMGI4lg33
Jin++sZqzfn/hI32dqMTAW1fR4fYyBpMoF+42vnqVtqwa/jza8IHqbO0Sm2sLjZS
0kzEcLedNcs977Ofib6aX63k5KW7eMQ+87mqj8XOLA2w7o7R3w/RCos/ciUsqDRa
cHVPnOcpQG1/w8ycsCATPL6jtGofwUmBxOTIpKDL5A3R/15PQBxHRT/oNu0kq6CT
RggX4byqMt86uwBhly6FS+KSPCRcnwpvw8MxP8+fDhEB7ODYh3PjbKLHh9mNK7B9
9acFuRwAzEAuu9n56Z5F7QI+h/wcI3dL6NATfL7pi3LW42CTjyuAj0lB6nZnvN4A
Gil0DOVUggcIuE4e8qqvIzIWLl2FLIIl7vi1gVHlPy9rGa2DkKPXzQZ3K21gikyO
VeS9977E6JjkE3IydDsY57NMceOgYoxc/GZazou4FoanZE3P8MIdZOHDOcieI3Vz
I6as2gor/uJPuw/lNER3OwNS9rBgsHySkqRPKcVyKWTRRZw98WhHAxZWdOwASYyN
Djfa+SYSm+ytW0v8f0fpOuETe3IcpALWclPtafYdLHYm+e3FTErCjHP3IcDUj3TW
JgJicBnyUlN6PgEZVydiJHoT/iwHLMiQddm+j+FrNzRcg2lra26zdE3LJ3hOgOs1
QL2VeGMvW6nciYx6St9CLsf+dhpBAUfhhEVSku38xCT9Iid7hUuv70K3EGrk8RuZ
tzPOuLIAZ7YXjAknMJhfVaqEVpkbCPvFq+KHvXzZoPTL97eFV42i98lcLp39Cccj
eRGrJAxGRsiDHLLOuRbdchATdWU8e/7hqVcFIGDghMVd6dFktgaskN8ksDQWCs3U
4jQeUPd+GBwfMnmvChNs0ZQhCvDQs5N8FwWAP8wJdoJReApC8sz6fjbfZ/Fh/Hg+
eiSZG+WZmHmpX2tNPxHqvzrvSoNkLv0ckS9RIQRdcGuSoE3iQenM7UOqxPhqzbgw
v6hMZTjLURxMSSaQpZqqbQB0okUyLeT2Wa8NzXFXpVcj2MVW1xRe8PQht5zuBnhe
s14VnNr/mIKwlUP0/+LmyNZwHJCzqmEgJYoHEqB21BpM1ao+V54xEmwMoq/67sl0
8SYYsvv+UsWrW4638ysBH8xfdRrDqCFoJRsteXiWZ4VmBymGvQPFbc6/dkrsXcq4
KPb2KvqWP7d14vBPl24ggE+b3HNklVqkTsNa9kiy506pc/gmurY7BiDqVs3CL8A0
bKtG6xSBZTqmzIpCBauthRMXhZ1RH0y/hzbDAu/gz/ZRkBWS504bTpHrHoIo8YYR
dhvopkYGjojkSNRukzQ+bu+w6KXimqNunDYjzksP+1tFaca70+QbPJ164yKRaGB2
aHkXTJpD62/EXtzGEmcQ+xRInnHiB41fnLZpRwPcxBsF8lkOOjm2w45O2E/fdARH
mm8x2NM6l6BYiNcDyqG1xzMi2LFDxuOa+oP3teqO3G8Qwx1h6fSwlV+h3e9b+X3G
npbvW/lUxl+hyIOseMPa9nLdw8yybVXzruWhD/tH7Cie1OLh+FdXyTwhaVW7HhNi
755Uw7BanofqdlLfPAi53XIrQuuFnqM2XQNc61Ht3Eo0Fvv1LgKyEHwnS9ZeSftd
mhCCA5LNfc0qi3yJ4gRjTgqSsT1IspvwzrGUBg3D83GewYG1YIIv9LYrHSys4UR1
f7/v3H/BZJ1BsmCPNAJxl86BUcVg/DZleHSaTAFGhgZfqCUCFWgQu+fzNpdAui3j
mKtvgFu0PPSJz2JiV90TQeHM4MqK8asUbfsaEjLPrWrX9/2k+Po83FGi/ZxONLiS
YOuOVLr5KvDB2nEZ1HI4Fprn2ltQoyBOtrgourDF/348j9nT7+LhLybJAilri/5Z
GgomXyQROTf06Nw6XuoqrCSW0JYhBdplMGnVVdgOU56+b5Z3HVbmN6DAtZwuheRx
1s33M4QIZABWzlA52bx4RGk3PF9Em+PIrkm0YC6I3ngouUKx2lRoKfWRNcao6r5e
Xkdbd04taC8+y/cnIxxOiSYxxmnkO/XJwzAk5Xrmm4kYUgn7hKaVvS2mSM6OsvGw
95skdYYJaQ79jQiHz7heVteJmYcaHH8H5gc9jQlertqlgB94wTuBBewQsF8B12K7
GPLgLQAjM/zsOL/rm49Mrkg9KOX+Urxk/ij92wxxObfeYTlHl6saZHAty+LyFvKH
0aXURyMWBkUFHzFUa9cz8S5hVdeVCS2zDaTB7ZyyIQL58Sjl5r6nGSglXvm70iIN
0iSBAYx7OKjJv+J5KRRrhkXiR8xWS0VXhLsuKcIhd3caYEJRHecDjOXdJus/rSQu
Fr9n5IFnrAhVDLjOvo+d0PmY+3BAmCHh5NLV5asa/owC+GRVBsx7Z9CfogJj0NlU
KwLzDbETCzzCBv825J3MLKrmii94oHJmJ5wnFNp48mICu9clkF4mBX7ti9l1HeIv
Eluctej2rDyH5wQGtws/zeCgCTS1PQ1aG1E5Bve5ehjj/DdPp6D5QJxxKtmdbHdv
EU7vis4lXlDeJlXzhXnkux/i4n9PqqOrs0xEJehCdgJ2r0rcwnitSeiT5xatokuu
izgdxjFLXuko3pteSfdIwcUKQc/i0q/zZLyGNhH0woZPgCChLrqEvNXCfWQSPIU2
Op6Tc/gUaiB77noes1Pj+Xo10gsnMIkd91+CtNLpwaWEUtKbzf0Ldx8mFWapoiiM
D8n4OFRpEXyT8Zp8xrkTH1sk9J5puFh+vK++mzZMsvyzSGai+isZ7yo2GFlBNj9e
RTtHF8Ifs/mT+WBgOGntGEMLIH1qozHn7Odfh9SmrLsLc6e3qha8PpP9G/pwKTXl
BWJK/hWfxKoBbcAgtS/FIV5pPWn43evxOlNnAms7sKmqtbVtCUCwoJ204Q8lVobu
i45dXMCYwcNLH2R3pCFghhWQYe5fosYF5EwQjLO4/iiio6PxpDJYcc+DDUKh90Pm
xzew3nXdHxYNd7XRgRyKgtwVvMJsXF+vaENVFvwc8JGxmvZH48KHiARIC47Y1UFe
5d37/ZfqIaD7clMu2+xL73HXRA0lRyalrQEzOJv/S9wiQnm6nHvvp94IwWabAkaL
IgSIksjVHeerWfsbsvVzhMKPbM0XrQNTq0Y52iatrQnduZ0S5+qaJMyoo+8pSWNy
ZMhyZQJHdmLRg5F1+nzd32zUwdxgCirpX8wZDxRusLQvslBonAryzyElet6OzvEG
vMUFgVp9v/qm+P9tD2qALcWQRf7zhQc4rqJI0/7VCoTmdYaUzf09rHTM3X8W7agG
wWbAhA6Y91NhIXPIhJGqicYkqfAfsllQF7zJ5mtTW+6+J8/g0XiCTDtYXs4vvqUv
bMvpOFtL0C1Vi5mbzGJ6oXWhIEAMw8cCAU5dYEy4dhb3upj5Qy4jBTGn282vf6kz
uCwLo3vmuqDP2+cfuUCBA3xqoBNfGvPSWnh0uYSG3rE0RktmoXaAiFBIyWtHpXc4
KowEYqwZfUtscSgGCkfaecLeLc0/ZVAGeIQgQKx/eYmLosuubYi9cpAsOV+abQcx
U5LE9gD6KV91E73SNyCK0Ju62ELsTfAqWsqDG8U5Xo1f3qOaaueijEWDep8MPGFl
UeFpl4eo5waz2FqTbMp8Sqbm9gjPu0+JYt7AsG8c6YTB5rr2go4m4/+96Rg29ooR
i1RqDj6wSOm5des67USUsZwSV22C5sH35J4lhVowY27ygY/peJ0JxyEnvjy7oEvd
cNel3zVlqyRg4vOUp+OuNhh9IyOonAaNJWID6vVAfQVW+Qvy1zt+3Sq4e2HvgIKI
B1QdnsXvT00q2RnptaozMf/VMoveZW1GUb7llnGBJWLcHeLyKnjWi+fr7fxMBRA4
2vE+1S6FJQpOgRhyDVzy/wbM9HDRJyO5I1eDoSC1EaxI3Vityif03fkM7xWLGcFE
URyNw9AJm1BLcWFO4kDpJ2YYU3qytLZKPqZiZVC7S0WVDd+GRdeg6TBspvUqUpAK
x7xa35bEgc1FBtZ8PFYJDaivlkJWPzzXiO8Jd49Tq/ybRb9tOC6yYOVC0OPio5DB
eRd2yaUdce2evffpZDTwDYXwZ2jHI2PaV89oyGTVdneVTwJ9I6VKRQSEITgCrlxv
mUlSRTZjXA6bkTw07rCr+7M/nO7Q5yE0amAStgATMR6+HzHgJVliI1YDotQloZN9
BwU5cXizt5ULQgnl2sH6eLG/MbX47csZUmuqBvUS3s14jiyfpSo1jlQUUIDzJaDm
Itiio8DiTf57S3Zk22srXBPud7veJJ0GgaD6JP9CnADFuzhdQPrwWoabNhvKLPkl
am4besX8uWz7Jl3uDjv85L6KoSzN2mCZBI0uBV4MYctwkw5g+QCzAQadPa4dTpJv
o7/QAdoniCKrABmhgo5b3+yVgnpoivcH+geDnm+cJ5BooJ+ABc/kCAxvsNbOotQM
KfHseV9gG+6ZzHEE/mrtdLCbeyqefmgnYrdsmpQm4iy/Pne10HIj7ckjL+7Eg9tn
bZN9YlBSL620ID4DZbT/oNE6ak5OtTfX4qcpbRAnuJZbphxWbGiuN370xs6HcpoH
IlKLvV1fVdY/sAEOfTzLNA3iU+EtTakcYCqR5kQA/bA5glrnOk0GQdfRLYoW6VxN
q3fC8bjnoW7hG+2HkEqUm4Sznd2NFdpc54CLzKeWa2GgDw73Cb2W56FPcXUzH/I6
OlpyJiWg4bJ3xn4fHbJ7IZS1fhOnlrfwPo7w6kNb/Hs+gongASDf+3aIaYuvpzLF
7laDH3asZozJ/+aCn2G6beGplCJ6E8wqyi9vT4x4mvDj7ZmSwkRO1DU/bKRI7zmv
Z/zaO17booCSUUP1NcWZ1SE0TDfJ0jxQxuMahuqTrAI9LwIGwYkKqprwdwAtrEkA
fZc5ApMZ7OZTsoNCNxyYO/uMQ7YHvdYFuX6gTscWifNUPTBEjOD0xHORxdkHJm7M
g7auVjLJrIOfcALaWZrc8QrN3vawX9Ig7WpVfWog9q58wVDHgPzs7Dao/bodq656
iaJwJj31zFnprlr48o0/bnJDOkOeYMtUJooiICUsApBOqUG7NDfxRrFRWtdJPnp+
OM1zxmMVxgZuFb/ZnfuWCGrgx4LGwHnghP10SUaSRqTioieg3hxunjWRLvxOKZGs
PVifd9TGw2YvEfAQXGiHEwwaGbYB85ZEgX9Xi8BgpWop7is8P9fq6KX5lIZSl+uK
GjxJt/ZoOXXCvqsscrdPN8Q19RWOTwx/BCjQteiSvEe8I6/GuCruYzAeDneNaMwA
g+8HuykD2JSgTwqbs/lddW7pNa17q/Mmgar45R6XcwWyu6JRgi3vUaDsR6it2+tU
yWlxDKj2jr/9xmenuGHjDkwe8gbylgEaIfa0Fry/ZRRXfjuHt550UUPn6addYqJl
Dq7+oN2aIhprNpukhpzTe8XOfsU+czLtYK2DiC9gi5NC+v6vE8eg+3PXMTnx+qF+
ndRoua8vAsa9ZeQ+ZIUpIGk+IbvBZspY0rHsP2UitzBiNJ9t8s6ir/tUPQsosoYa
WFeYlyIFWg1QtirMaCp0Yd5fR1/RT9+BxGrFrMxGFWT7/0JaBr1CMVAvNN5B39Vc
kBiJYgAbO9E+UKN9rFcLI/ukuBdkznB6vQLgfeoBkBM6gqh/Y+fHSVepsF+4TBle
Rqo/1voQmB2v8YJn15Yxk+q5ImduN/XWbLaPt4yihakQiuZhzynyu2jYLLH5SUR9
cbVw4HxxV27RvsTdq/u6vVCkfu7KNQpsPnwWGYUVhTMYRPrckrOtsRTnc66K4gQx
xmUITbBfIzGalijfIOvOrje2/L5mPAj/ZNj3/WMoYWUUXusYFg475qounagrRPro
B7eWduC1kcEajpBWccYqV8WL7MxgvOZ9mJk+Bkk5ugLowIlaa+04EyyWmIN7g/42
jsX89t6+K7zMs1UJqq0XYkqmDpm1faxGe3p2YPMuPR0ly2pJJxJ/MwQ5+r9bLJFZ
bxAhTs/n9zdo6Apvr3zXye64HHKOyU1w8fCQmIsIqcFmjHzKZUC1XvelRVutiKPj
xOUk+7bgg8aOEoaIl34gETs2Rh1t2IWTg6RXQ1RFdg7c5/Nsox+cGT5UGo2GCKaL
fO5iq3aw441ETD0Trcgmh2wGVfv+AvNxIGi4YUfhDuxfG2H5+wgbxINUp/AHSofb
WAD5cH9PIul9NlOc9Bjv72eC7t5Bi71FUHS2qwmd+Rcm1rJA6Lg/C2iGGn5n06SZ
o6geh0vIoXCMkQ43s5bpZA+fOQCeEiorFkS2E5eycsjyr4IU3n4XFWhO1OTg9QU4
jYfL2vsGGhlWw26thikJt/Pb2LvSqgZvFphpzutfJ5jJK3wcBcLzQRrhqT9HK2dS
79zYp4JQna3daVT6UQ6drEaLvBVoAq2cTZmfZLiCQCtJQhnvOWi/dZBl50YrnNGs
8NIjSx8Hu7d5TcS18thAy1KF6VxXArLgasZrrwXBpXnNu8MelW7GKTpSwiaekKj2
1fu7w6lLKu0mSjrvw4kcKJnUApI3DNM06/KHdgNLWJLlqCGxDhtB6al5d9Z4e00V
IP3fmtUuhptmJFPx683WKNuOtFOXRivQkPoRQUSQPXMLuHxWRdOFoUlar/wQPe2K
PW+ePkkyafjPN8NWZWNm5IHpPsZhRH8CRVo4DVm64wLR538D8d9c37ZFfsXIUuka
5jf/b7mefuQVxoCWzIqUkwm/KVbBNDaDZStFylKTuqExSQQ4Pp+oWFHGdYfKlYj9
ghtJvESgukrLxGerfd4EymQFwyC9/pyNmgSYu9Y8HAI66rw0Hgp+Gx1NNsWhcJSm
mmRioH8QXglAY/FVHvtXEzBKrVj9xCyFhXTdoDNLhviF2dlEOvcf8ioe5+OHm3kX
fF1zjeA1uThrnitWgca6W75r1n42vGNmTOC/XIIQNXcNjwROH4B+xEAV9SqdKtiY
hHmFOsjCZsgoadWaa2GiSikDWCKH9yGoYnWV1gX8cpEv2ppsUdRk/x/wlXLP0670
FPnchhoHPqbUJxRwMwkw0l9eDiV0bdh2Hke7Fc04cgCELjQ4rP4S2zJn0sNKdwWh
f+W+miepmdP8IY2BoE7I2rAuDULZarYX6P9RsQR1SQsmtLC5+ESYIj5SLu1teHKB
4ObtOPGEELACKDN5+wfOAA1d1j/QWp9wJb4LmPZPuKmzSZeE5Qrc96gdC8qLmwQP
9yAhibblI7y6wY+aD73SlGfOmzi9a1B82nWHvICFhHahcMra3aj1AFA5+tODsuIa
RJEua8REd4UP7dy4ZquH3Yp0bgtn9ooB3C8ydGUYPPbrLgBgfUTA1LblRsyuqmkh
KxlAS19C7wkyTeoROqqOqF32vUTynJn/9Rc2KVevrEtuafo5owRFnpUijzMLBnBf
yAicwxRbsXlKwrVe1jXQ7JxZXSsAugxkm7JOmB/esVySiesucYnvwWI30U0QObYh
l067WybLzjTfxt9+X4dXgkfoFqNiy9TytA7qNt0Xm6ZbM+yp5pUStFBW7SwghJTn
ShJnHxJLNB1Vs7mFgYMotIOA25p9ftN5nRzxMmwrrbz6BE6V5h4yqAFkIGezIg8J
98KfPsdOHYQRz8OYTGO4rvNMF7QFOUXyvH6B66NzrUlLTkKkyeyEYPyaRyMVpQAV
BUGp41e80rvyGZrAdoA1xl5Jc1vqb9jpK1z4ytOfRvAf+SC27A9A+/2X/lL39Axa
zLyL6Gp9qskxqyG2SbMy+Nz34/hbNjI5x5pqTZu8xYCDYjOAz8FAxBxerWzeyblN
7byQG02eHs6CT+ltY+iYaoRsGZ5wi+GQGp11KuvhyjVDDGDF7vTh61YK+TmokuAt
0QGGOoluQeALXj93tbZy1LOntYK8pDgtIeyEAZiApyRsHvYi3yqjktOhPd5flwRO
T0e59dEWMYoy2dpu2ZjWaWUWrVoZGqkxnfEyCz0aDnJkrPou+KFBqo3zJjtvL/g2
5cLAYVcuSkBEQ3J3CGt7T+tRI82z3csRVB6FWoJM6mPVQFXW1IJVSYpkFoaIGAFC
Ols80YZLpbl2eGz37CeXMfcLzdoQkf8iiBIwqjLUngDJtfYYqi9JSeKS+jCio6s8
mK2hcKYpba0pq61cAzcRYAoPreURYLK49a/VzhIZYWUlAuR5evhSMd+2LYbtaNS6
7swLqct/UvzRWcEwdz3BZS35jHMnzbxlwpxfbcF8ZhhIgAmtW0n+805k2eEmNICU
Jwq2iO1m5mQ4Avk27kCPolJbQfFtXQ0wo5HBS6I4SV0p4YBWaUtcy52o84k08QWJ
1lA1sLMrwfVCBy5/9W5BhDTAmYFk14KNZaRW9kryFm/xnw/X3RkZWT8ZZ2mQVK9e
ayEV83xynnpGfddLR6ztQgVCO1p79rYCfNk1IC8no0kkO5SHbIFEphO5QFINLsfi
hjDT+fsjLGRNc8x/s+LWHhkrG6CnFjdfFQpGF9/1gswQVKS3vblNmn3da1P6zpf/
SxWUW7EOEgXhNxlM9OAeNvLg60dtv9qhAuqNlXjxM0uctZOX/uD4DHk09Gth20Es
9KOx0EU2nGAx8CGElOyQlM8W1K6vM8RzTl7GP/HwO5qsPifp1RKQsOze91MdkAE5
LPg/fOmj8DZZ5SH41XXW0pCYBgXVPXvUhNivLPDw6sWksXiuIWm3k31uZF8yDBMh
3HDWD5UgkhBkvle9dM1/gMhGpBFbmdwYSPgz7vs4xR4oOcc4EJpMmEPdctmBU6hJ
KpsS4U5vzP288RnLihTcVj42CAJ7vvnQgGp6IR+CDcbD5afKiBuftdIGATmSVU3x
M/5g9h2ownBY67XtIbyiJ9Uxpr+6kidriFQoHcUiTuLZR5QHjj3Z//rLtmS0eBeg
j1IH6WTlqHabBRqlqb5ujwmr6tRMa/iu5zv7RAu6+snyE7SqHkFF92+yN3M1F0h5
wi/7jNaO/m4+N9orK+a72GGq44BsZ+lYOmImiCSAwfrUzM8brql0aIMf5aZ6ti+I
VNILP1cqGwNg0yNubGQl1pWeeOPqY973ddMAxb8o4KxoOvQpB/Dv68KVO14xB6gf
qa1skaFuJWqeoNXDGaZePCeKsmKlrIoA70Zbk1mOIzBCbn1UBNE1hmaBUJDXCSi+
PgUVkbG3xkeQgMNASA3jKOTtuvbrCoIwKDnS9d2mPpEMnkJXMRCCIo+rpabOCwgq
yjCcESsfuE4rUzgBXPtsmrcKFCj5QM2UWLAd53xGJjWVliCX9hYt6uoAgGDA0tCs
ecjyY7LL6qhyANe6e4dFEXnQSZW8XtbRPU0bJBS8WqGoER0zYquO7btoRQkfQmqP
f8s1tOkVzPMDVKv+S23nirAhd+yRN+6329Ff27OJigilQ4U2Vec/mtrCP+vkOaeH
HTn/KlbJj5k0Ue3WUemCeguNZo4P+pj3PkNRQ2Puqj2/7wKm5Mw2Ms5Hy/LLsCdX
Rsc+k2LMLGSePpKMi6m9x+LdAl7WjbscWkfvoDW1GtibJXpYjZp3DDk5GLq7N16f
+fKrSn/EiZUI0ntovCiv53+2iQddgXkl6xxec0hEPVePTFi8GIqLd6Qmdhx42WGS
h3JeURSD6XcdUlfbEVkdndK2g3gKGadnuOeSoxH/lsPlUB61TKQbWUYzDi5d7niM
x99ruuIhu16+P7MaJQRKWXOJ8CexC0llWXoRrJLB8tGdDoNrgt5MsSview4fSSmj
YhsE5h8U6av3l1ONvwS303x9JWanXbZ1cLT0CXqUNYu9SKIF7DtQ5RSN0yWAT9dn
IVDfyUtMth1MBoz1iSx92kYRrD7WKhZIp8y7dDxdbYhyKRsDEq1xvSVYySBR5Xhu
wBeD9+VdaXfClOG5IWC0IAvmvzEB7wIUMTFdbWUwBtHxflrK+1l236NoyKx3rcrk
0F/LHqJf3UVgTeT2Vq6BYQ21bY2tGjoZzppaPAayJWqpM/ikOfsnGkFrRBY8aPY+
4OKq67Ns2M+49J9Puj1fNnAfX1DEAIyG5Tnp0lFnA0Ul1zM0d7JKFzIv17I4rG/w
dwpK9salyLNHOxOOoMJazNOe4C7dJ4svyoKELBllr7g42X9pxcQ2vdZ3NcOG+6MK
RsqPj4vYi+B0fICcE9+IdOifX+t0u7C8aEeFmyu0S/nM4v0q17U5gMoMRvoHuuHv
Zbzb/UnlRK8cC85IMfjvTyhfEgTKUWT3zJNkfKKiD60v/ZmCCVpxmiZ6XpS+Jdjh
6HwY62maLOl6hHj5ra5fx4Pgmhh1RAlGo2q7FYIUvShpDc3BrKYpmuZD10UePchE
A/lRUkuIufdYTPjPqRuLeA0NaRdbGFdUaQvT+XSuNaEkiemIvFk6LQipl31UOn9U
wtzJ37ZWwgMWFmRWG9RKdCozr4Pj8Co1uwOIhiBpzrV7WvB5yGloL7r3A83o1uFX
vcIGCZx5F5nCIFB8Nm4BcUo+zjNOlqy14WHpOPTMYYpLVYiy67i89eaGG+IOhEfA
wo8kh3n5tiulDBrPMZR1bpsdu0isKFHqN+4l8CdCJOpLdPP37+sHz4HW2g8bPtsO
vVDB4zGSTJWoH8ZRzetYSWKH8SdzfACRkLLFGXz2cK2ybtmNFQmijxMnKZN66ozL
o+YblbfnBF70QGUSBB1jdSJRlkekrmYP1U6n32zndHeVWbmiAEayG5x9GVCbWyQU
DdDWinXACpg9uBYTUGjxA405eRJ/salb3iy9xToB7o1fZ3TxISosmA7NjfN3MVNg
UipM1vnD7VCm+5vZqpu4BUy4tjOYkEZFWMi86mxxFPI6I4/1r4rU3eGj8bwYb3CQ
P9saqemBY+2zZ8EjmlkJssNMyqIv52Dk36Pc1lckNOtM9rC8eL2A30ClgsMhAbMw
oFer3SLJoQKsMXauPNWDiWP2OPD5n8ngOsNe5tJCMpMd58GYqSn/o8itcKnDgNIj
kWAgS/Wrey0jg4c1EQy80uxd7n6dOkcxEFkKRQmr5UnpZtfv8Rsl5UdfEnbhkgD4
Tt+JgH3ylM5/QMbgeHmP+Gbi6TOi5XsHhRjnjCwdUOLvkeMd4vpof9Am3+re8BuS
PJLL/V4ldJ2Aav8i1aXGCbZ8I9f8+R+Jn4a0QBWwMa6SGEmetq2IQ3RHlJTabamE
MM/DJ9r/rSNBr2aR5HMnBJHgBNIRhs3kbLZFwDVLYu9os+RWtszvaz0RQdqyptov
aJZcYIHlSfQLEQU2uIzmSsA2/gq5DCL5uOZplZwnNh0HO3YMznCOPpcwodhaS7hF
ZpDq0k92odx2eT+MObVmvntdCXsAj+6t2GcTtuLHtctTZzgVqCe4r52VlCXpkWQn
Y+OwKCUluZm88aPGMqWRdX6Ov2hn5SnjdnVGm1N4fIE2jbmzusvVbdFVMDbd08Js
E7oc5OJu02eiw1ek9MTVak7U5S536uXzWD1QHCN1S43Uyavi4x/wAeDavfnjVFUd
Kl5x0avwskqd4TdTrRcfC9NrZYJdfZ8Mhon+N1fBn4/gMtmztZ6wIQb199WzE29K
79DMpNZIVlysawYOV1QNeCu1LKUPXlmjRiv2kfjF2oXld5fJJYLYmfbdjyJ6ypWn
y8KOrKJb77BKzwZWjaUaPbFaSSqPQgRs3L0tUpTjRBcT02DUEELTNDdIMQEjg19u
eZqPtCACD0otQYrtM84ERQJ2rvxhTq6FEiIa5h5kNwGGTeVR2QB8SXOU1fDvTiII
WI5Qn1ibk8di/GOzRmFHILudB/o/AQAqI22qEPmMHTjmbXCb6L5I0ivPvCkXPkVO
PhBPlvfc6WPZcgf0BQPLrD3GRiL0+vn/ckxGlYWQV9KPc0ovg4vtfN4fVKpQANEZ
PX3eiPlFCr/IpKTiSP3wG6x89x4+JAwBM79Ja8iTt0Xz9+Wltd1Xsksx/LR8GWO1
r15m1AcNd66U/Asi/IgTvGDuODIl2Ho45FHwR+udyf83iHYe2669oxUEvW+KBzgt
80j4Kw3vLursch761JivG+1K09CR4xFoLVK+KP0IAhO0B0NjyjysJjMQ/HNVlGRU
+pj75Hg3IdtwHxwccK0ELi0b0f9HnsSqlVPkG/GZMIyfrlHaKygwQ0SsfTGe+d5o
wxesYtvTmDJ49Hm/Bps41nrIeqDEf7cK43W8ngf7Y2gpIAgN+0HM89U8EUCuLDQV
JvFD1/FWYNXH5wgjBw/0r7A2Q5XI/b+v31kfSRIcEqSGCWbYDiBNLWYbNS/WJWkN
w3NGUPDlpcx/cZeR7N916kHbxWPtDR7ErbfqCH6W96yVMewl6OQ3PpkV4HUntmqP
6HOmYSHY2b7Go9uTv50XKDI+aEHiG/u4AOIzXTyxNCc/wp1uWiN5xNlKkKIodVX9
TawuBCg9tGg7wp9k974TD5SU+tbccfO78RvLToxvUvRf/KzX9xO0a7A5yvSDRsET
OPkL8pGsU9y3stU/3rGRYW6VFQqavIyVU9bCJyh9QJWvSySsL+2gmIsZHkQKKleA
QqoAUq1SpCbgjGeaQPpNGjLYoCIy2DhgfJpwsxfvRsCxHwccypDtA1Wo53+za9g6
EqTdNlpiagS2JFjaijns/dlHtuloUSgfMsQwQOwqvukb408ojbpBxK6ljaDdBSRC
XiKDk9W+2fyqQYug+uPMPVhsEGPkxFstoWIbjpY565VVrN5r5xWZ2tHW7TkCx0nS
HhVwNZVG/yuVQv/ExaTyU3qrOECrJCykFDIFT4NeRKLUBzFGfYX4T67tdHUsf4gr
noFACUbTtiKgGmH5TLvd9uo/hXZt0vxBltInaDzx/XrKRk5x9z+l+HguOxNMWVAl
AHPW60pFY25oNl+yDY/RZyrmdh1nv0WKJIwp5nY8eNOnNsfWbg9t23hZVeFJmoBM
AnNoXcsut3rAGSHOAxjQwfM466OAgEV7pNMlnCdOL3J0jlrdbiMNLlOC2LQHdRqV
IlJj8Fu2npt3kJhgiWEUA7TRAvzkHxzpJX9BGFJSmIdFlgtIPnb4d9YEAr18y79Q
p19NzQnFfaX5Aw3Pa7ioJtjQ5Sv05HI2vDb4Wl0FsP4r5bQ6wo3xvs9LV0HIf0q3
VuJC4vDTWsoBBSK8D0PVcLKIvzqJ40+WGWB79eRc913SnZYIDrJAQ8oGMmk+Rzi4
Ub51Xm1XgIcTDmCo3+8maLycJr9/XkTpYY7X152jxvDROVkkApSteSOaGSCUAPK7
6/4uoENrrjPPxs+RTy1IFEzZNxByVSODIG9Lkeo67wGKrBTl98OGM+ZPeBXFMMHJ
QvhGl1PXWiEbVoXlec29sWoNCix8WdQXco7V16WP5p4GAEughWnIyV8V8XiWQFZl
mj27uNy0JJBkgU9B8v0DVkaOS5+9Zt3qcXiRFMnD+Kyvchb0Xj+2wfNIsrlkyuZw
XGGr3SoGRKNpZAzwS/Vu3YGLstARd4TkRDpoC0l8HG0/X9m/DzYA/IMql5nIqKV8
XjgUUYiyqM+ljm9vko/T2sf6+9hLYJCBW11B/yI/vbKst049tRodb34Ag/MCOjKB
5ebSYpbtQOdTCorqTct3rFFd93B3zr6wPv4UCkpuIN66xnaRNeu9nTPcOWlF+gEg
+cr51/UnMLi/C8juM7wC91bid1x8Ut8pScQd1tTX9nXT9xTcjhuT8sA/ucQ/bFiW
FPEuqxgN0XM4ta5ulO5IE2JCH1t7FHqIS3r4tiEB3voB1YP2TVCYUbHrUqgptXJn
4G1+xh4Asy+cZIlWP7bX8gTG70bkos3LyJYV2KXsx189oVLVLvKL8VPyCBlMxXIU
nzngGL1qPSWVmHfDwTDbk5m341v6Ltug5lH0HDfYGEwwNjkUmmlH6rCd799oIb4v
OYH8Uq4fN+AnAY5ISJzQjfWLYzTkREbyiH71/AWWm4k4N0k00Bt5KjEgGQLiZKl1
5++eKZBMDmi8uU3NwAPWklxoGY9hhzlk2dY5MwgDfl2l7+Rn0RjPcCCCz/7Oj8YO
HSy5ZuwSLDl/9VsNATIYjJKQ0dfligV0zxVJuDFZlT/T5r59JlLxefUSTtXiiZQw
A/dUAc9ZD6PNfiFsYFDm/ZYJsyojyodCFPRtS4luDvAuO+u1PYd7vU0r6FCD8BFl
VwAyW21Cw+gRfwxXSAsqbQVu4T4ZiGsqoMxHVHvovZFl8RexM1918fyzyBz80vWS
EMTY42FM/oPc63pGz5TzmFH2636hB1yZK4yyJs7iAGSOEPahH8REjTySIr3uR6+q
zRpg99wWsg6thk52pf+yk4PgERd8fPa5481lNPZepShBJ6NmN5/Mcc4YiWFc7Dy3
iyk1D/pzX8kGQqHGk+/Zayz4pYDlMNrv8B2wHJSdaw0ThHLX2mMtT6UxWbSCI/pm
c5IlSMQmfo8L03aoL0eCixH7z/Ej0PY9qHyUYj4AuDel/94rbNJHjsdTr+ex7S2z
pH/LXqeXjFsYzX8yCzcWhZKgcfLrrDJ53BGfwvODIeBMTp8Yhg8x00SqnsJ/SCNd
YHFQ20fP/8cGrc0SaBtt+wpxmn5oRoTdUz1jKUyI1Lx3hEoi6lgsRqGC8H+5oD6E
NoG2nRBaSVl7owNEl09H+QXAnSTdfyPezsLOfjbUxjSfOcXENvGTPt899oidko4D
VNdXjD9RGksR3mmHIVcG9NtCf70B0650L4hQTvBDzt1rV6yX2TXSlZqhymlddzAM
Ql3LIRIALXEjthjoQR1L8jgTViRqoTfHdWTq6cGCnnTCftvgkhPd3TsiJOkqS+98
Rh+kj0N4IJYDmmJDgI+eeXj0Y1OCpHOjPLsR/cf0L8MaSb6Gejmb2Ads7cVZAVVy
UcVXYdvQgQReqxAEXbYYVLlQgTKYkBpGAjdxUV68/Ou5oDP/l4gzyE9gEMMEqi2B
pNllWKJ4PDqrTE6lfUeViOjeIBPN3QUZOKuKUxh6JceD4iQojfGbHHBVSFO0ue5y
/ITrpfgy8yIgAxoaQApZzb5DyzcyhNFrq8/4jVvzWDIPJ26qMhHyuH3NjYygDX+H
j71KtiiLOZxIiJ1bh1KXo86MtWVXOETDAnCWT56jntJTtZCUPqgNivQPoIPcDvKI
uXm/MrkRHLd5raYoJ1v4TZJCGPZtFiqhyDi4olFDs1yt7g4BU3smGkdFPww81RqG
1Wi6sxwtlR/wLak8OZZNWcyTTTj+kaDcl/JBwnxqBKh70giD41TmBk+CyIyAaCF3
FotCqmaugYHx/3si2E5QQagWebeZ6WZNpLS+llR5/E/b7QwTnGS9wyuG7bGzw6+R
S/55gsNLsP+cy4vbfrKJ3feDEgkLtBSIlj2Dba1oH4A1HhxGYy8drnYSWnNKOPfO
UijnDbRTMngJnWode3EPxe1BFwRCFNqJhzn/wTgLY9Z+pnPoRAKtPbyQ1B702Sjr
ozWm/9Nrg5Pn0Yjvyp7c0clvdK80kM3x1dbxryj1TKwM//bXL3AJJeWsGpa16Xb0
+7G4Cf5AnPuiTNugrFchMC3QifEVHvJO59wxlGohYQfZ8adyV8GOb1XRbFhCL6AK
GCuw3oa/hj+GFU8dAftA+wYCTynm356k14EWeWPHTj7P8vUie6Zpizt7qGXk7r49
v9U6KDS7FZYXWTQoS/pkdrYNVfXEnGivAQ0oDZOtvavmhHy/gyquLXQ54jzkGj/L
+R8lcdjDjKERFcwmoudwpn0rbSu4FnMJ5IrsHnoRE8qGLOgGNYD1H/sEr2LqgloV
g+O9oedg/ugi9VU0ZQcQKoZps/o+dRCp2L+tdCt6r5cIl2oOui9MeXEKEB034zqk
E73H41pbKO/UnO2iPcBN8otqZ22J3wo511Yb0at5NMq5snV0DZaEiAve6IKkk/Bi
8ds0FRMrUlkoFg4KrZODLXxc2wyz3NlXlTi/TOEO+5pMCsR+rsG/M0nFXOYRSFZG
zrg+yCp11mRc9GNCQOB4fQvPIG1Ykmr1x6Tkx9ENYQscnOL1qwvUBLM0YI07e7CX
AOEIlrb4iXkxesNoVtgBRGgJ8jsDV1O6KImgJb5vqFUp7a3zQdb2xPvOi3tCSAuy
TetJ7xfgVopImv8bhjgEZO1PIgTY+7RlGQZMPboD9UFh2wOlJ7cHcZ69jPWh2uyA
C4GvD4eDVJWQcN84ss9v5pMyP4DsS/9rncmKvSqOR/fQT7XdOl4PZlS5z9a9pwSW
/igqMnmFQMuhta19E41DVA6QVl5aESvJgFGHwK9/dDdDSp2tw0lVCMEms4a4eGbm
XQO+2WoK11AQq4LiEJ95KpJPe7kw1NFgwOhang4/Ij7KzcVNqjxdxn/PtUwH77wW
RagGohwik/3oKsqBg4iB4wyX2oxeTTL+9xF9UeFQ+VPt4sdrlljj07NU0fIBb2LZ
ssyHIxR26ukUU0J/Gxw5McgcglpDiirn+ddPsyv0fgXpvF8zADj+SfsBm0WM4Qlg
vAxf9Ic63czfmjRZYbRSZqeX4AUYlfcH9pal6CZVGZoD30ghHncgzZDAeKWYUt4A
qRNjK7gh1xn7/D+jq8trUNct8Q0mlZ2I3DBWH7AesIC39+4xWOc/dvjaGhgosFXG
q0jV/Iybi11Uzp+8leWiMzfiXB8SpGOnW6WwHpb93IjyFddPwCQynMGES4IYQLcu
z3WrB7LNtOZanua40lTXA9S0nweeRsKgFBUp2/EXML1t7xQQvpY+lPTJGEa5EQ3E
nM/VDoHo4gMWu2TlS5q34CUJBU6QlrVEsQOHBbhS6EsyeM6Tonx8KwIL95Iu+OAN
JFvyh4JoDTjRejpTIZAOwtUUy42HYubHSGjOI8h19LvLJsMAjDptzr7KTFTihYsk
e8WWA2uTw9sifMsn3ytCnmQHFEJZJZHiYXyUbONI3Ge6kXk+/ZM+Yw9Ab0CVNiPI
DGPGavlT5uW+I9j0p+mWidOk3w1C0c0a0V2eKXgp557GAxKdjww8tM3qx5NuXYYW
DcBmJN9kO2i+Aa8fMUAT0cGkZM9zQLpUiCZnB+BVJPFtYuFtt2mTAg6fJXNlrO5f
OgYKeCrHd+vfavxMwJADLWIQwu0S+LZ0iyzU7L5NbQgmj9VcQ5GxCum/X9eFUYWt
ooxw4BzJJgzoPHGupKS8rpoxHn7TzxAYZM7ls77vQiXlWEl6FTx1Rjj3J7GOKw69
csVKm2qCJr61ebbAyqTC2N4ykPXsUrocADs0ifrB7dXwMHeWtZVGG9dGNYbj2A++
hSx05BqKvckvCK3laxbBd/no5MUsy+itzdNxkDPlA2lp3RIGrKcn++FMTBR5C+QX
fad1S5zl0RXCm6e5IInJXex4MwG6Hv9eDGnztQ1iKP0v2gD272tmZL8+hgdTwm8d
K5X9Jk2jJKJe+AGINC4l54HMuXiD+mEGHJRybZUXoSt9S9VQCx1cB1Lp0dVIRxJ3
5ufjbREgeCLQ9D3xJlYki32n3deiXbw/bLqoXKRy3yZjtIhUzOzuiDq96FdtFR02
X7NJrMcYdMRalcXrGFDsMuERY25QOIJhK9JjL9+zqbZ9stlg5WmeOrPnTr+4LpMc
acsSO99K7r2YyZGsb9MofhZz2uM4chH9jIjPczovyBG2HVuhJjrQajSHdc6djmIN
LurJMTd8cHLlk5xeGQ9vWaVCs6EUW52VLrNu5OgwtuYCgV/IeIZQikSO7FNlqZvL
EZeVa5M/EdbYNWcWsv0bZA8qoKSQr54BEBs7cXntbCaNV16V5c8RGn/QR8Zu9fLK
2rXnTJwfWBk2OE1y3t0l67yCVQqY9bi3w7XSDvcrBgH4ClCV29YMdKWh1Z/zXcE/
mcO6tlbYpI9aTUAL9OaYLp0tRHmuExQgvnjxa3CfHjZ0KnlkyNlFUk8HOCO4eImA
O89fG0tEImrekNBQ60wKNrAvKdOMXKEEPPvrFeJmOa63VNF140Uaj6wklNqKYH7J
J3RYjH4Jl1+n96s204D84seRbm2Qx82wWhsThmhf3gdSTPJUthOqOGHXKN58/11L
LyN77ZotnmT5IU+zE1BzNHG5u92cVIxYKa1EJOVxDy9csMY5TVIv+b2TCJUES+FF
bveuoL3cnNs0L+OkLtoa6i5Pe+zEO6pk8XBn6JhIgNRuy8gun9AIR6IfsaM+sSOy
nMogboKD5ml/I7e/6Lem7TQa9/+eLIMzuRQctHQGo6p1cxBZYbP/LihIjN1rd5Qg
E/Dm/eTTFTkGnXx8+qLwUTo2haPtO1zqrenzKxba7K4YR/Rm31nxAzdwK8ZM9zN0
CGXfXPPOH2FUUPltWWzXupIpgnb3L+stlivvkcnBgssnbLNaTCEV4K193naBwIuD
v9Zk6etxnfufZRNCuoGjLeSpWDA51KJjzxX9oYl5/xLG159ve0A5o16k9Q1FJFv1
LybdVmdoIiD1abizX+RoJ9hp1Rm/kdD1TfOKXW3iCa5lsrA0OPGLFMMhEs3AcGFc
81PEsvAGoplxjsD23bWvpqpq7p1waozOP3srZPP4+lTMyzJGvOh1FQdEGHXY2x7M
mMmMbEs8X3aiXT0iA3C9X5iNp1LM2tNGltpXeSyQxOP13BGvtzOI10WqhykZdT7x
E2i056hw0BA8CNuatda8X5ZMQbnLcwYijOIO5YOdR88u3xCg7sOFLXe2wzdhg4BT
Z1bBOtmTEPcdL15+Y0zz1pZjdfJolf5VW/ddBfIvSKpkICw4HLwuatKUxdg+Oyae
W0BbvXnJCBCTgTEKOkjVRo45lIcGZ9R/KazPm33pSbppC2MXSXPpvb4rshnGkKz8
r1DZxxBBhlOh65OZ3IcpvHriIpIBSWhtwtDBmifJob37VYHC/f/vp7HpdUD1GWzM
qCUYM3vwNoxFajTU9nEFFS1kq57lX70vtSz9IMlL/pv+FEXYF6ArdriEpE8GDbTy
5rVf+MqzGvRZEmVcgm1IiYNPXOMzfY1HWy0pOT4FZbBac18TzikftfW0RNeohWyA
P89D6m6+xkWfe8azjEQyvMEFcyvl78Yy3fMFzNMSbB/wEjM62wWkffZCiI4kyJPg
Ewsore3tTsAQ9BVW+UkTxMaKAJrZkkwhCR5eiRns3j6vbPLn1jtZ8P8WNVbCngZ1
j+jdqTM5rdXxBvOi3hrNOyhVrwuN5ujkxKDoE14RzEcW6YVmrF5f8pMGmtBl9Awn
9d/VvD05m5Mhvnu8/S11mgK3DecILycSaXIGwZjLwpoyttviyzS0MtS7RleVp4ZL
eixs7HHGffwAD5IzcmlJRkljBX7gh/+7INTE9Nr3BoiShKkOUZCUMhi6W2LzUR5m
o0AZlQYKw0FdzEa0sKE8eS0oOC9UnZuQGML0aTnyCeDuDPC4JHQQIGkRUQ3JyNx/
EUT4ryPjT3Ag9Ba6wLo4naUvihe3qDQkRKJi2cbpBoN7ewbgvagepyy/qjpgnaKC
+LHkUPRsj0jklQ73ZxQ9iaw6EuxrNBCBkeXeICIXin3jFkATwG8BES/pBIPtuea7
azUevHLGfCCEtvgJ6vlaDSBJM69Wi9FteCiL1o8kwQCxKnpcIg/FBYdzs5iBF6xA
3abJVIuiF7xWxjz5RYGWHHkpQB9jcfdracuFbhUoc/O9rmWMrB1Db0xlJdCyTrmE
EIXC/v03mZNnVCtTMFZZBmW3xvVQMdMOyODJoSf5u74zVAtFMgigm9WmxH4OHRCD
tnE1+DUTHHPwCjX0oF6SzJ4ZB+w1OFuU48Re6Ke8uvW8pSEXkl//PVVaU+k0K+5Z
xQ6eWq59VgbtIw3GA+Jx7RMDO9bBj5mWiTN2OjMk4A5Sjqp+i3zH+uZFLuoaijOy
3bI1RP9y3ObE5eFNVuhDlJFhEygsI9bJ/iaMfGAkhIZzHupS2/wM9Gn9bcAzXx1k
BCZrDY9nih2WrLfECvOGHdWUDP2y9/tySLnDada4OBMVkyCOT4BC1f4lVMLaUWSX
DrEco3ecJGWeGRwYI9r/GTRT8VuNQzxG+VPuQjuiw0Wqe3LEJ20L/ZhKRoE0Y33j
q9D7ms1+tWyBsvgjF45gQ0lO8Y6KrLECm+wXL0ssCVhk9ty1HSD1Et4zM5YFt8CJ
tRw8bzOc2qVgDCZ5WwsNx0xG4elfpa3tyseuY1Il5PU2ui9acPuC67LqMKLgPKnT
f7Qjl2u2920cW6cwh8Uq9LoVGZsG9AvBQGETIZ21X1a9xSF//3Ppm7vovP/mg8xq
JiNPl07FUNotbpv4HJv13KKM1cMhuL0Dc7NTnpcL22AxXPakFyFCinXyA9Dyy7/i
3Ui4d++b96qpiNkTYN9jGdJepNS719y7Gd2PtV8OQ/C0Z0Np3lHWkyftbhXbD4Ou
m+k7hsYOukwcxsdN0GDC4TGlDp8dH3FG27W6l5XKwBltVzz3mj5SknUF/rvFetZF
O6KhVRX08dr4Kdt5YRHO0ET34Wo5T6WuOh7dK9N/lj9u/KCRMOZT+kqqddW+JYIn
GYhTkRh5aVTycf7oNskNsbzwcNSdTDZkRjk/137kwx/46fNhyKFQFN7Bz9f5L4/2
N8+YkyNc5trDe+ZTll5AMLSXZaBWek5QT9Bphk61MfmGoD63Ig4s/Uqp8gj5d8Qi
fNZhNP/QcrbmvmhLKEcDwIeqS6EhNmOyVW+HkcuXQgAYcbV/dTZ1WfNmAC1ei+KF
wp2GOkG9klZPuKUP4gOVtbVtZv/EOtPbZVfA0VvmAbJi5PVlo7iwI9wILyFCiHyk
XCymK6G6d3Gxq8Pr+3ih3hDsrhNAxV+tA9YvTAiRw6ODqbhDc17VNNHBoRF02ZUV
Jc830BBgDnTpBTXHh1vf94K2QsWbM7B0q1W3/tZ96Cp/DDF3dAW8G3IrMMU24+4t
duZAWPl0R6RO6dZtQogRL3Yr51h35es3XBQ/3IJFDAG0+pUbZ5m/WBPVartmOkmk
d2pxsVf1r3YumoSUwwwwwYWbgmscuFFJ+zMAtRjw94N3ftuahxyoCTNFhHaLvMeZ
/+xjuT6gCThJwoi3YuW49houwxiXj70IL3AQHiENgMuIxmen3ZV0IkniTq/6vbUR
Xsw43zQsjCp+4KDcV/8jogx1Hk7khHsrkNf1yhRLNs+jAHbsuNICLgsBA74iOeV0
8L4LfGk1Bgb15Mp9qKZfY1oiB3M44Fj6XQRXeFB1orYm8CUUaq09apsPCVDwqrzm
rRKFmfQ9U6Ew0LxsX0CSZXSh9jYivX+XThjmqkL4mlo5CfdJ43FARXadT57/uM+P
MqcFyWI0MENy1umq8EYnadwH7agoidS/gyc1wIbVvCj1suuYGTcevZumfdqxBUmg
jcoxlhvDrg+z2EluX9rbCEEH7wjtI+3K4LCL7oPjKniOTb4vNQFuzXcHhADuUzVY
OdEueP2HVsNz7r0NzTFGhQ4xDpQM+Ad0W/ZcNRN7koLgzkrU/NiINs6tshPjgmP8
tFFFQfYSqo+0tLTrP2zLeM6fYoGVlMgq/QltiJzLJMzxjNDOBaBFgFUNecFBx5s6
Dc9NJjsjB3ILhZvEdiD61nY6Tw5GymwNwPxBvUllhDjBbddCyGpv18vgUhGud1JM
2cDfXGYbk+MzKfP49RoGrjf2SdFnf/MmgwriKC3BuSmDWFg+NfoAXSoCC5pFk3uV
M7R37+Mm8fhQlI1Fw9sP3kUvUCmRI+c8DyL9Q9bZdtovWJujFXsJaZjqnOcVK+uD
zvqKLWQmz9AhZv3IlQXoEzpMTmB6FwgTtnGg/d166G/Eg2JU2MNJ0ups5fQFlSSl
7HPkZRmh3UQ8g1ryTDB1zynZsnGfSDi+JDk1UMtJM241O3Tz1vSLiitwoEIvI8lZ
ob5hMpsCvmftQf+pFHks0TQAp/l2KaajBeB8Za/YELXHnOYy75EUhEg7gkZvdoig
HkiDJt2FOb6LN9Q98UW39jmJNMC5B69JbkSb7ZPtmEbZbUo6jZXtvwQaMYMyFYnH
oLTzJyqljjSzcKg91/4lbToq4Ceay1AAOldBNPPGdzDzOTFq6in/iIBN2kUS5AWX
34r2o28ZlLBSg84kp6FLFQPtprfVClO3fxOJxdBVYEknMV708x9ksl1LfsQ3/qsk
cg77cTqXB/VD6/tD1g9pSLGqR+9sR4rd2Ll9G20OINFmnhrHMQDHbrJxMuTVmJBR
dPkZM/KHrpGZ0ecxwwnaFgZK/Cv4Skn41xlIWAujRs2ue+PU2iKV7F4ABE1maDP+
4gxbKvHmM2G9bm+JzWRIBJgQUWbPPptICuvROy9xT5zjAQMrSFNbcK7iDOLFM2rA
NUcaYqEbeXf9CV6iTBvVrexscgf/P/h21JBIqH7p8e0IDvVOe02wmmzaRZmhSEey
UIAeNGt0S2mjTZp9UtevAIBYPHfv0vb3JSvB560gU8H6Y4112ajDnbMWPSBvnbf7
ab+679V9Q4sGP9DwWYfJkhKwpKKPdLiXXrvTkcauUgCJf7XLNd22T1djJKaBvJz6
yBSYU+pxqbMvafReAgDzWevI5Whly3LJEcGkqHwbCw+bciTmANCZKj+9KSG0bMvC
R5D5MrlcwaChnB2SVO8tLcZkvJOlVYF/D/wacXLWhew7VRyOG2ycg45SXeVvqelk
81i7fzrwGhTeDSg1XR1b81qls9l1cw6EvlOr9dPwdoYL3xlRPs7HqlwS8CDYpNYI
ZmKGNFuHNmMWyq6/4UhQp9M3cf9IFrv/r0+zH2dMx8CHIzuzA005tEz6mchQ5lFl
bPTnVhOs3k6GtU1lCb9KVAcG/bNrMR9acX7K9cMOjgohxkK0+WyPfasiAwQ+JtGc
lUWaMveToEr+c3uSHYxOuxCl1YNu52N5Ydil7iDxxKRuOfpdvH+AXRKbsoG833qW
KYMz6bgNIIgZvR3SYHM1ACNm8R7SzsBTpN5Byoo+XI9a2cMORHEPeuwcb305kg+B
oLvlO8G3QigeoP/s2dDKHAUZkPFtVuaCroI8VHFNCqLtEjAv8ZQzJIYFGn1BdNaJ
4NLFTL278lLFVjgmqZhi2ya1ZI4Hs+eYE3fc2mQ1xtyAD33zTO975gSfwGzX2W0Y
CUwVQsvU7irju4TmxEl+juh/4D54TLCa4lKhmLbxXJdKz3L+7O9mpXElYqW85jWp
vR326MhP5kI0Bpn9haevopiPFg/O264KpdOhJ7rXlCn1mDWOhyrKVqhSwe5smVKe
ElKteEE0BxfW4m2YT/7LY0uA0PRrxAibPuc5zGLiEIIC+23KNtQkLS4UCPcyx3V9
5R/VmP1by8NRhIzU8HS+w4Tcy3MWTFlTyTaHom5EOeNzTnuUeRBgMktMlAd+D3tq
yIlziQBfrw7BNzXzyVS7baDJ1mH0DKM52LcEGqFSghcQd6U7VcnD34weGR0Grwh5
GObl4iRsHdUtZu6o7dxd0ouOmLsEAy9QNV6rt+jOd33huQyLTiUH/1mpAGVPJRf2
Z+uw7vJYSKhNfJSAFtwimBgiha2TrdQq+Ezxq2T/jkJh4AkoQd7ukiMIUJAAIALb
T2mBkCImQHiftn1DBZPyw+4d844K4kB24pcwiZfuNqZWBwjxrFYNugLAIP+lCCPZ
5xF5gd4B3DEu3w19qLh+uplh27/3WondANvcYXH8hX5vzCq+2WIEd6gH+OjdFd8i
XCqSmfGG0n09wswcCnSFmSc0DYactyDAcpZgCwZdfCKk9cM6VUzx7NOy1DyZ4hqK
Jyv6NmpANTQ4+dQZZV6vYVQi2OvmNwSh9IR+4cwaOidgeigkIYyfiizbDZ85qFAJ
cxht1S6QWxkgVNC9n41QFLD7sChdXFUM54yOntKIB4lTQStEyTljtoJJOw/bYhDm
uVKrRw7K+6ve3OAa4VQoOJrwVyCyjwaEge9NPIM0+PsCzAWISJiBCH/Kc/4jiOO6
0BQEPML+AJ2UQ8XQCQk6TiQhabaAlSihHvv4nDg8M6Ax7wuXlrJeJBReVlSO5kxE
pZ/OA37FfT+37k352J9A0r4ENpEmTFSSCAQJVWLiXdYnPAJnPewijC/Cqu+GuIzn
1t3juKSu4vztoDFUSWWD4pEjbnTNl069uYdAIt3GX3loRvce/KoM6oYmrRPaGjhe
kNmeA2UHRzq0/LVqOmEATBQvfYTny8n6JGkGL5/+3C/zHxtXDSWgEr43Hc9cMx69
M9akpYOaZ2tOGQIsHPZ7STaOw9Ao0cfQ0ZKmxXLG+tN8/ApEtGP3cJjWpJz/fXrS
/CvAZY43Nv0Vi+Pj0H2jgh/p0+XNA0PS/s7ALbtJKLY2DMilhLOke3waLqNJ8qbL
ohHgauIAv5uHQgcThnjiva4LjSxkx9OixGf/hIPB1clBoMWoN6pIUpJo7DxlIVwn
IdJ6ArZs/413q1mOaQXGG94RZfsJJkwzdjZsRaP3+wEiEhvVAwcQsg89tz2hilv6
LjzxDJ24czSCYHcHB+1aIiuf85mb4CPF1ZldY9YpILJXPiQLcZkLPjHsx+RIQG+o
camhuIapgwy2/SsmmG1eQDEOrUoYOH0vLD25w0sPBvGwRKEouIyHCItGrJW986sE
LMS+0VQPMN0ct45vbdCEdsufgl1uCi2fHQavcH1qJVXNGz7p/yETpntBmlgfTWmr
mMiWLlfQin/EdJy/kWunMW6KkpyZHupAq+EdyKf58SQ1ek6DPJAYpc2YewlUAWSI
oDX86LMO6UFmsw0WrvDQ5Vu2sJLuoyKU6Ofy9AOp1Il3BuPRpr1ASJ86YjBjnw/C
84uQ5+w2gO4RYCNhBIHZy1uuI0Gcz9ldjVQbVmQ68S4nBDsInnYQNbK2Ay6I6bDQ
BT3ruCE4Oi+cKAPErb45YeDbIMjt4w5FVmqzGOF4QuAH0YxZRQKiTun+5aazq6H/
cWYdGH9aUWQ05ME0H51YBiX5wzqjhxX+uU/uqamPc9UF9+bnt+Q1QjbC7+s2/3h9
JYnEsHVoEswP2injwhDACBiGVzy9HJyhEgnHP2M6d2JeGtAK5NaaA3jhgvlz7jTG
S1IWDdAZQJD1rLoLqWG+L6r4fW2jrpDz48CzzYIVX4Xb+lmATbEWddpdyPGKSzwu
RkqDrEtgFo5iS8J5uNCpt+6sj6cN7R+WwWU+Z57dII1LEPH7eH5U7E86txZOWWtI
vq3pAQxxkW7b+Pg8jH7HSKJkJU2wpFy1Ni/MMUV9GmIbo6Tc63+gnoGgD0XBDAnb
6NrE3/xwwz2FGsiUYkM5JqT9TYiYiX6cYfRdRgZhKAU6MeT8VyWdBDMFI/W3/laA
ST7ARxQv92AFRsgGCy3bxFRId5Ex3nxaen/eT3bEbkNs3hRFGILcUeFgYTCn4i3o
jFnaQYkJOPUB4inKbZaoLHV0M2/MmFI0CcOt0baiZVkthKVzv9VuKG3Xisqf1kWp
N/oK+RC/vbptCNlfOy35Pfa7zL6PQBC/Xr/wWY2jsHcZ3Jf3ZacCdy0jqKjmAxTO
C/MfpquvO2UrJNR9v00xZT08bA/ssKBwE0wFjvP/qfqt85YYerh4gG/qLF3fvGyt
kPphelrOy9WXPt/1ZP8uJQrR1biLtiQflRyGfN3xuFMQt8pBGZnxB5OWgF3C4YON
ULpVdP7YT9B83wtktCpE1e/3gn+FY5/OobmwDiswIw9nkDE3Q1uqWMNNmhhgzUT2
ApRFJrYhQwNARNxv1nuTFvWgWU73YTuwYlWfGuvJmW7zmQkq9qXbttpZDDBUgBpi
S+cmfsU2YtY5VTyibwgWmdtOp06w/JiDzTJbyvrMju46XhZoyxl/wLAByuG1cAfs
hUr7SuaIs20Ukd5hVp1qK16XjwPrin6zg4L27uh6dRgKBQR0GEJus+CDRDBpPDAo
bdIc3yUItlwvkyoTLc+Hl/sssDeyLo/nx3+/TReZPgSIYhsKd4QIDr9AC2ZyhEKw
RNrNj3x+UmC1XRTuGr/I08w5qkwtTR1yJZJvgbMd6Zx3ndRJYVxRdT9U43LG9cbe
yPvIck1kSrwsIFEMvX6O40oZXMj75geDBbFTpX15ue2mFkOGs9JFu8TcfZg3Z8G5
FfNzQRWGuj6v5Uhyj5gfclTV0DNnMT6FTMPYoBnl0HzAgUSeEV9VvKyPvspZUOfL
3s1tm0x8lKIiojw6aQDP1A+gCH7d/H2T9JWIE3o9rTzpUTIFr8Urs0KqQCsN0SgB
lBdZjT4mueC6wY8U0tjzHbrUMXnVuQ0ajBC/OlYV5eRqXMAppPgAZmt7t2DuEhUn
55tFKhlUJbMe0EETCvIxhgTB/a6pymf6+b7tPfcb44iZihv6nbu3V6kR4FujvqUK
+fA+SWNsIT8K6MbxlII2yR9NnVDIimevbJUEl/gnR6mtrIKFZUJYckYUaZbbGrrz
vGY1ZW+tvs2iBPvX/X15w4zswBK/ly2kxRCwSCk4CEeBR8AXS7GcTru6fTK3dOgQ
BYoj72a8KGdVg9RKIJzpqE3qSUOQMDg9lpSOn6KToUwdXXY3L6AsYLlwS0DiycRh
CtsztA8Bi63oAOOT5cnemtwIOBFTwReZoIbDSLsUbMKJc0Li2EiD/WIVjG0iFFmK
xAPS4R7V1OBJXw86LzZ4t+cIaMlOLWHZDtKT0+T6nMdYcMdlzINhbaNX8d7Dt5sA
kTPWdZQAE7Bw19SkuD+Ac0XLPYzso8jSkFK7dDTXepBkQirl0mjwkY2iZiYhuEoG
r55QjedCdZ7OMFvxkoOQ4dwLnQYgSup2hV0Cuv0rea5NUEAumemPSCAZ5PBWQunZ
/TwbV2VBKBLibZTILy5KGkY42f3ELfpnb/UwlqqrQnkUE6rYQpd/esu/6BRpzFhi
UnBzV/roH68YOymdJwtq/MTHb6Et8iJI9j3bB2yg7vFu5D8V/j3G0NGG78cuf+YQ
RtHTT8iIZB7l4Xh2doPLTZ79rmLRQgZbShfSwNjk9nEzJA5yOD15Y7z/FDhTNgTw
iHuZnHsxL2i/3e8HfIwLYYwEHcpPtyXzAcdO04vJ9mRqd2N44zbqNhqbXGdVpHLS
K92TR2hylBUxRSHNqKceI+5slhiR0sENI40lqoqBcsdun0jKJcQxPT7Qgv3ZOYFM
7SxjezZsPmRFhwERZTAKjZeAvbRBLW5NTlRicdPgqyMsGK+aAKNqeaq3na1nnCOp
xfs/5fCrbOWu419ut9vAKlgSUZ1hrGda6P71kbO9dYUE97X8c4pjzD4R9VuyLVgH
V27sJVNggF1Vce2R03BFduTnh0BcZQQ0U9N2XppzewpjswhHghTNBjjzoJ422wlm
F1SRcQOvyCbSRde3Dmm6TwtoUECt0RcTq1g6wApPhB9jV2J/63fjfUtC0LR5VmEi
OTpcQoUtlxDEC1UsVgKz1PARW8wbnEwMqqX2yBtReO11ZkO0bCoaGH/fVUJjnnxO
8lBSZzM7TpFd/JrqcJymk5Nk7lpyimpmEhtuWlSFAEPBZso9aE421CUNFehjnFUp
evipn5kufYQKhLemgNADm5dtbRiNvHMnkb5Nv1gglluwq/wzEUXyhnYvyoxscbZe
lBSJQF0Xbwm9ZYB6DtUNHjQsAOBCjR1VeKrvysBnDj5zlLL5hzlrUKT4SDoRhONd
npCtrSZ6G3rIl6QjmYDK5muXig6cLM32ut9Cg9K1tncZF7J5DYrlofs9fLH2GvOY
Wc8fTTER7zvPFGsTE/cp9+H6NQ+piu4127fqQnNePprc5eUVIBPA7Ifluxn2gL27
OrUX2SMZ7BUJYB7BGDJAMjBND6//X46DRqWBLIGsiR8PLfQOT0MGnfeuWV9a5Knw
X5CGgYTkgMSixKIstykLs2H8f9md17djiafT9zyHySQ58yp01BiVIp7n2U1LSbb4
Mn1M3cep9K5XO1+irlS6TRxJDQX6s2eQm0ijWnZGUFY1wNiAn34Z+Ttl3Frobyqe
pLJEV4eHbp+8irThLGcjpby3ZgMqs57k0ZQg8XSEx1PtulE0f7b6nXeT8o+OdTUt
MOBWPggq+nRZp8RgaKgPZn0ub1alJT2zL2KaTuy7uuk2/3RzMliem8PI5KFB/RFF
/RUWViZGWG2nCoRoliLcjAeQQSdtRlNu8hvY1rqxd4jwaQ8tshdrh1uCfCixL1WG
2egsK6ujB6ZiEEZO/pp0rOiXvsZuvBqxP6TKRrdhrbQYPwxr0WHmnxLM4R4S2i/r
Kf5ZFmR42xExcQzD+5kFJsdHZe39UAZ4AmEMTqc9aepoDCC6xFkuf9m0dYp/wzMN
oE0n2Li+UKP8DPDKa4nwSyTPe4kg3QZkeQIxkKzFhSZeU11emszrHAY/MQET0rD0
1FHxsW3dHB0YZIWS0hg2WHDWGwuLVg7AFYNSwPExT8RfaU5yWl592gYZathWqs2U
EzzBm8mGZQya+kwrzCDjkKsUm06kc3ZhLDOZiNYMw3StRSfvcYlntvCbx6ORIRna
RqUqF2rlPg3bL50xbRaw7icMGLUfEFdFze4TX+H3sRTG8OgS2qALUe6YZyxrm0NN
7gvXMuCWj9z4d8seG2Kxc02pfaG8rOec8sCclLAYs2ZdtAa80MXln1wFSArhPbPZ
QxgpdeANdtE30bdOQJWqIRcgkMoPyckBFBBuBOsCUSV174RBbH/mRa4YIymTQ0Pc
Jq/rVSMGsA+JBtvdmZT8GZh+CQohAr43w04TWZVQGcHHHCCHS1gZEykn1FDROt8O
BqZ5CQ4mS0KUQscOMcW/kOPT+n3RsvzKARYqdM+hRxi32VqBD/Y29IGWGRPVdUdA
84w563ftcQL1bQvb/I/s0gxhq71NRBOBNqOXdMuHTE560YU63zgHthVvOIwz3ds2
ydLxt/KiywYcb357PlSxVTWLrC3GtFJJ/vby2Lz7MZkQPiZ/de3woCVp5bX4AFiM
e8UlbETH92OiR0ZlKBddMg3iUKZzwa0LidxkWInPADXLMpC6BEiJRzHHN1pHlN9J
HGu9789zVVzTCNSTCV27b3jxUxUeg1EBZ/lXELkIst97DpeG+pJ6qWWNIA8Lqe+6
vq0ZSy5pHCBKwboECrRX09vsTQRE4sErObSZy0Ej6NoAJdh/2yPeeXrssSAg5Efw
0/3kaslAFmimMNsJeMMOjhxnEab2j3xm/w1twHm3EwELOaXOjls61PXRUczuPLca
v8j30ln3BDdDOgsRc41pqR3tnne9MWEsffDSRnqQlVlzpzG5F43VGq0Yp0bj80fJ
5fjpVWTbkYurAM48bRPfzcG270qN2dpdoaZhixL5PkGCcG4HZG9BdGz+HVhHkS0H
/PSrsaA8Du+x49t9Yio3DLTtI+S4FhTv77y8Q/SwhJJKuEy3uCurZk0kxMyCpNCl
9Okmbsx5I7pgMuiBMT+F1Wu/+0mO6+xGLphPRC9RrAu6ni+8khQ0awAUj6io2p6L
CX/YFGa+EfwMY9w0LeJ8Lt6n3nSSDe7vCY4TyXOOgupYZ1MXDtfNB5kGGUva23Cw
zrUfDFqFuvwtk9E7NCURvzaSbUbhAu7XQ/t8h7E/4tv3x+03XVUWJ6HWCc6Toeyw
0vAJkkKu0lJezr6PBAXoKBSjXbC5DfSQ5CmVqP4kXgRrdPLext5TGTUTVYaLj7FC
xQTSrzaDMlsl352W8xT95uFw7iFdTHimVryDHNl1z7ms61oQS6ISYDFelo1/Fn7R
aaZaC1sUnq4zEeXrdV2C0HQJKhjcMXcp3qE9vyZzyoJ+i57X+omPniLPAKv1FEiv
xXjUs0McAFo2VSpUW+y4Bj4joJowJxFiMoMyzx9g3TcPJD+QjHjEJsaaX2Op1amg
rDXaULNFZcfJxHCvdhU3olEAZAAV3BJJgr1zv9WloFQQwrC/0kx29qDl/aSEVcsu
BHyQoorGmA4Vx+jKJn9/njp/gsivg1gtR4FfOtV0Gd7JslzIxjBCJtMgxkt3EzBp
n6O4dRJwa4CjUzO76ToPPhrNSp+DQSqL4LBxDFYbNKjyNHsA4qCz84O6FcOOTzBN
S4VgUvn+JoGI+HDZ3rY+tj7U+qJs4yZPXvlkqVcRAbn0rpJ0MYNgztQPQgyu37Zc
MMk4KRlM3Hy98Hk+fx7sSTyKz+/tGbDfrAjIdhW8EY9y3mmddNmUcEolHn11Qo/4
/piCSRNKR33AzV3cqlDofjSR0sM/l/DcSdvERQLocvnsEVsIVEObdRsI5TsZX0/c
VWfkZl+4TGYlx7MHgJJHkU3gky9whgh5aDjgd6OZ/SdXr8c5Z0kburmBrE7UQeks
QEdthVTQUWgrWFLzjiKD3Yq42EXOWrrVe6qWzjPlx+FLSvRwcXLeQLpaTUtnI62Z
Dc+95BV+qAkKDV6R3DwDVZ10Exc0cG3kbkz5Ij7EVTFyDULunlWZPqNosH/h6lCU
EQzoTVd9B0Y+/Vo12RVPLr28zi6Uk6IFb4WbINt8hANyVRZWdx2rZ1klcHThnE+p
2D5p7iaVjHkzke9UOyulKHl1fIzVhbvT0NbGxj/4y22a7p39vIKq9xZrNixqX9Ur
H2jxrsvgSd7FLz77pU/PCKwYIGbxKPbVLkSQA4eP+iYvDtlQ6HZO7B1A35gIyX3q
3tdpxtrpRgWGqfUwoURnVH6d3tFIvv+c5Dr+E74pez2OIXwvVemDfyaIsqq8qNLZ
T5Owdqecze31huVoXZc9ulYtWMeyTI61jayWhpMZ06jMus18BmdXlE/FqCKcjMNN
itDYxtm1PYUAw6uNvvb5kHHdNqFd0QcBAPQbqe4ipBq6Pkg0LxyEEq/2a+DUf/35
F1oPSITlKDLJuDf88g30KXVD5F489gWe2D3kZW1JVvg48HJBqpSpn2DPHi/cdqaC
jpDFxfF+5S8lq1mH7xPDflz8025ZFzAVTCIPoJITWYMKxq0H3mHxYDRDZBKGEreK
GVrKkF0ueYX9/+WW8fn//E3RQbwkkqev3GAgZC7xLQcEeMqCQPTNsKkumQ45L8KB
36d4FrIO512iEeNhui5ZF3ah3Mz16tODbgpX6b4e0WqWDFKNjotBH9JomE4p3iVV
luHkccTN5scaNijqFwVUi+1N2QKlHPCbwdC3HEyNT0bIH8a9iWb6KyfVmcT9pP69
r0AlQTb5vBEELZeb1Gr6KN3aJxsc/j67PqbgDrHUe3tOgFXNw5dJGszog80Ip+V1
Em5S9Nauf3ZeqRON/vty5NS08fVRQXSUyFxSzoNyuZzOIJ7YEBu9QKPYMwFxzdIE
7feOuUWzmFUFljzZojXE3fF5LN2eLAhWAbynS+5d9KiQFBDO6XqVJcI/081QofSj
4yYEy3D1N8xbmUXmHtSM6WxROQUrna9GWxJl+eWexJE6NMjnTMpY3W8nHGQrwqPD
SFRIokNFUzZ7QHKo4uSrAoh+S25JdoSv6Jz/K6wdfDLfJX2szuBk3mTOIyalAGHu
umAH3+I9v3n2x5YDzfP3Xf8X3f56M6UVISMZc7BNae0dLXWG+HWR3g73zLdd5s6u
FxeYHT9IcTjIn7n0x/U4BGB7yFDAIhbeiZKtEKtnCgT2wkyNTe683HzRZWxFE/s4
2F6hdD8GNVFPljjsPxZ2ea/U1KJqQRnueH93pGgtVzdIKVvSuerHvsLo5y/XxLYw
yRzSWT/bcsXQVSTFcKxfOTvNg4V1Wwynm6/vvzfJJwIKtyyBN18aezmGroK23xbX
lLYZESJ4TGDYBPuv7T2ofrrgdCmT4M/YP9k9H3c+4LClRKjke/Ms7itikKonaYOY
7ToJEPQvGMb/HEoYHYnGJJqYUgbjJIsfZXfnENNF6XDbOUQ+5mdE428irOF9c2Nd
n6pyVmk22+iuEaWfqmQCaLzI4DoGYF0EOmBgecEJizKwrM/xyYjtAmf2alXKibo5
GBYYa7+EX4hQc/xUniNW8zH7ka4ICrBKkFW/X+A8BYz0zu6mjhtOOPYwdn+xg4Re
DUo80EvfzuuD4/t3rsd8AHlOj1zT+XA7tnbR8QiQ2UIb+NEJOuAcsN1s5KWhtDCW
bYfOJ79RpSIEiGmjjVfG9OFqer+lmTSegJGyclcUPcbG1GTGLCc/RNUX2m65tJwG
bOW6QeQU5TWifFdUmIQlcmrx7DaC1CO69lnKPbbbsrvc3PY9BH6W1HRD44xN1ivJ
DD4/0zoDW25Svatwjg/epsCpE7EnPkSI/uhKb8kBjc0kRN9YepuolJUlcejOqOxc
joY3ToqLw+nBz2PkHqbVAzDCFUrXWldQfucQeyI0EP7fKK+/SYv+I4aSa6/lSMy1
fySIeNwfQW+NYd88NFYHEo+uxn35MeyaH+Eh7nQEi0392asnmAykDFHrTYRaefek
fVA0ezLKX2TGxmAiK65dxutlzjBg9ijsQXxorU8jPpt2/4kvV3CpyByk8BQjPd2T
Ej/+BVjOjGjU+iThL5io/Upd2fY7Kg1ee8XgIKcZJ9gFheAcIkI4C7SBtokxkhHI
qeemSGBWCCDGf06DWz5iH28noBPCIndFgv4lsf8bgxMf7YoiatNVNx2GAT3OHM0A
g3IZY1jRpajy5C0sI+/wIzBXnEJyQ5ugPwqsZOsswh6BLW1m3mTl/B4m7XVkL+L/
nJHMCFtm/CT4F0QcsaEpB0PNQQkCgE4d0Duyn+XicjS0PQRhOwLfxCVmv54tsuLN
lnoLWEqBKRzqvvTqXQCSgbYRMnyYIkCBGFU8buKS2ga68aN1MR1nJc8LeyC2jHXT
lY3Yxfe7eykzlM4wpv9WUnPEHlzay43GOtIM6/0xTAwOiygSInA57aME2v7QezpF
6eIBTfbPt3xDnBaU1jL4HDtGNuKR0+Or7gbkgJO/w+hv+fKXnZZ08DLDY7Yh/mHi
dJP46LUGfteYbz7OIVKoyoPbaKNikH6U6FAKWlsP7rs/tYgR5bD9UIl2qf31WYG8
LzVzb03nOdbHLm/1yKpUSPI+Jy2lFq4HeViaBiCK4ycjoCy9pYoAmLl421WdZ9DW
JKKM38VSDT7KWOQLdxbLW5v/wbptIE0zw0pyoY5bXcGRAmJDwNuQw2NanVfRyU2x
v1v8hEzJTE6MijCeuAZfKYNDwoleiliP1Gz+f/YRHHUQHPx1heIFbYHSo6e52Zjn
g6WODM11Hbx1Ya1I3ZrUz0ALmI8kQH9BGC0+md3OAbSprfYQygReEcqGQEl672xP
rzeY3eE4f5OZYo+0x3UfMxWCh/CQx+DmhxONUOoaizsb0W8DjCigKWB+I5513+oV
2hYmUzL+eV9eG9db7x7Aj6EABC6D/JbamyyTdiCCjl5t2zCTITgPDfvwQwL8+TOF
kIf88KRgWszCfmRr3OlWdiLamMgA3y9ZtNIxOPLapJZRt+5DDwLR0sfXh6c/mCbX
N6w7n1FX7cOy7OziE2LKoCeNPJvTeY1MNxfNByGGlt4yHLXxJLhr9GQpLu1UNYOx
KiOe3KJLeuNUmRCc4yq7JSuzmOYRZHeeWz0YzrpIjgsrDziWm3GfjSVJ7orcHXsb
NKMMfW6TvLLQeoHdgfWrb1b8ph52g+rcMggtAN4lDWqH7FM5C7i8IMOk5Lf8AcV7
8F2f+WFhi/74LQnDmIdqjpextlc+ku91GWjY/jCNR+rTEQNZNa9wWsovGHgtl42D
YoPXY47RE3rBnOCpeV82mKUtn62YATcadC9plNBnM9wcsjAMZx/wldlN7YgGn9ro
XtxL+RziFNonFlcxGE0d6MHFeO2OYfKYa/68wgKuartmRX8teEuwrygomGu28NNZ
Tv1Ly5Lti3q8pGr9fsUhU1BB+TWQBXK5dcIBjXO7vhg/oZPXpzewFbrhxoD7oNBX
CSlBcFqYoweaNaVZgdxaIvULyH5BtNKR27d6G7nwvJjut3kkI6EsxouwY6FaoyT3
eTVRmKfBtHjoRKbKA6PEL/wzM8cSCzkrS9gDVK6OE5b9HVTfkBF8F0i6rvMra4hF
cY3eSeMZNpTWEQd52OQlJBVzfCRPi9Ujc1/4FgOog8+/lbhhZ30K+NXp5RkRwcGb
eqjCSt9Ffcq0esmtUqedE8bbhYe5MJ95eDjjtmZ+jm9tZx1XfxpUl6iQDHHWMQa3
sIQ36juL59foFoil25fJvw+HRrBuF+aBtaPG2O45Oio8XVjytykHYnMrNH3bMA6f
vSpxLlr+x0DlSOxJ7CvDo6b8tZt4c051oqH5E6mQd94UViCPWDAP3xxVk/ti2TZP
misoixZdwbxp+VCNe2P0iCimI0AaAZKJXQGYw+6K8k9pKfIa30JBmZgfg2TlGxbg
bBfTzf714ZZ/GKnc23vMy5iS3WroY7atOj/uJ03oo6j6Kp+1azbRCkeJ1RpHiQno
F7zCxaq8wOa3Ko1DkpPj7WNyjVAb11ULmEMpg2FY2DZTPxNVlasnRyy/lch0Nnvn
Crzr5cnHmVYhntPRFE6OMcr3UeTioidRrWWUxUuEXRLXK7cOVUrX0y28aL2yCUg8
wb8lG5mVesdQhRGN2cEb2DvNBPDBiKj08Gj6TIwKoE6sZ/voA230qVj1mztBDslg
uBeADKiksLbLQE+2rSjThYvTtHk0X8nUwYDeMreO9VXcbOJ5QSEG+twmHUUgiPRp
lorJ/S5L3Ihy9hHJTzhTGF2rps1488Pwza48wKFZReNQpQJ0jiIK1ox9buJbmEYy
KXGq3ZKGsVrwaL3LhdUfdWTW3b8wGu7029RWDYs4fLjreRXh+FiQyAYZC+QWSwnM
aNs6VaS64vwpOt8ZLR6lzOTDhe9729e8QzXmC7An8iesr9x0ZFCuUgZZPRhtNh+8
bt0tXbF/F4l9miJbn/ke2scaSYyhkMf3CQikBb8tCYoewo/TesCHodt1BwbxHBF0
iKGgwDYQaBi15q36IA/d6srgJ7oqrJkt7y4MzsohMBsQXeg2DAX1KLkj78+Y8E3C
kSq1UzxTfOXvvHWmzwf44Mnn5SyQmQHRn2SblcPBXd3Awa25b/tbS70lGGS30AZk
Z/RKyKMSULql6zSNIEkb+9EZDnFLLh/1D7rKvs+hvSJMRxlqIpMtGAY6v2xn9wrB
uSnEx33BbfXGPLEa4Qj92wyOMAnJtO+ET413n5xPRqo+OdAt0hs7NByd38TO9YjS
pmG9xzGikmM6C05Kz0cb+Oa/0FU+VAjBRdlP/rYngzG9JlC7g9QJBrqghyU5S3Ud
yWEM5S99dy6QKOZdIow3LfOxEfQ2nj30k8Mfy5WFNdiK9H61fOnRpuTNQMfx0Gbb
Y2C7e6atlPaP9e8c1VqQtp+ukpn5oWiw7TJvTTox6Qaby2/h9K9PSBy3VYDq/w5E
XlhsbdyFI+UfxYwUHduGAT5iRSVGeRhniVztORuA7I3AZ15kPx223kPJfP2NwnGx
3opPlfsVwUqlvnLTLnfQUxzWu5HzbF4AssuuOZO0VOz56vmhmC2YbW0fi+tuPsB7
u8Xw9fJjSxd8754bA6jkiIvOJoLPxWx0FGKZ6W6n0970SswuonzjyLKIxsItwy6e
1lHYEcFphQfVRu39VhxKJYw8QcOMmbtG9+3QFAyTHbmpJ9WKv+PWQuRgDfve9Wb6
dOdC/UVCM5a2CooousqN1lopJF2AGmO7+6Ghp5m0DBrm7QPQNhKiV06v8flmDrUj
7TPXPntUPs8CCEKeYEvLwfkxBWzQwCa7kReuFGespwT+5WNV83SkI8SzckZ5XK+5
z05krmrh0/oe3SSlWJKQ8HESQHdTztOPUGoQDzhmAAjzfIpGIfHEL9JHPJICMg5J
DcVZHlPKSn04BtniJDVhAQo2GZfmF3dQnoTvDhnbLwQUppIExYBrbqbjOZWIk6Lw
rTl/ZqmpfStnRd3KlLdd/YJsKRSjcEw/RWr8kKJyq2PvjNF2wNbLJU2pLBT3tNXs
g9UOHKfiAnX7mS++BMbYehUtEtWzalkpt0jg9hH7ZZB9u3uZoRAIXDLAh7gBQLan
3X7hQhI+yn4XGQ8r4C8lVYR1CTNS1oSPipbZDMAVY3DiPuK3YpwLfnzOEFc/uCel
UNaEpXPMEInFwetQbArmErJK4CGOcsCh/UDnAmptW2+lFczTa+GXzc2mSi+sYbdw
OyHNoezgsg31G83WckbMvpN0sC8zUOS+ZIIN1SyJAcXleifh4oc6X4dv94TkGBCw
xYHiqwTWrsckLOKg9mp1WHOcyU1ru9IxLHXQwfnctvDaliSJG9zT/tCo3fWDySlP
IeQx27fu501lssWEzR0dmF19UYK2f/7jXYXDb46qL6ioPmnCQ99EcsvVVBgGOOto
cokUfYDuftp0PPKvY/oOffA9knuwrBlcQBI7Ty2a8iFJgO5NtuZGz8dTwJ56GaHP
jumaMbv/qPJQs4a86Cr6xk1VoFvSV7wnISIpEO4/T01Q7jbrj/pualYjkAjAwXOj
57xTj4WqZfCGp3Kj9Whbc8nQePa51XioQfbMs11540p6Gc1XJkCrFqmDc9InoJFS
bMc3yFiLq4o321CCOJ9jxHCL85/DA5f0dqqm+n3M3pL5pgfJXbV1pnyqU9ezlaNA
p2DaQpQ8ZkHDAIIh1GOHez3xEludBr/c4OKSz2oqozTrYySjmgK/lre/RLPqJaoq
fPdhty9sDgRdyvfowmTnNAbvvWKBAT5vdnYJL9T0bwdbH4uzTcXRoYnTwPxYWasr
NpcWawxeIdmvvUlzN4J3pS0tbrClCsXbXal5YCdRHb7A6TQOE2TgN3oiy5hPZhzX
8iX2Rpq2Z4Jxa6Bzl4ZcmhwjiZ1zYpK2PXmhdMTqU0ExhN0WMGZplbUt+5d9yJkn
vzm5C42yMmDtz2CiFVpV6wNS3XUM29rU+/03S6fq3gJ7WNl3aFEYTi6SBQBciNHc
HIPOcYwUG8QyRTgpmEIx9BA7HGGSf0iRPwQOWfhFCTRATT/ZQe1y3VI0DcGMpZbj
Rj9qzx26sjzkuohHQ0g3nXliKp9A4ygFB4gH5hZaaSwvFEgF2Q5Uas2QwopWvrOy
3BOlaafsM0rW29qqgX6mb/fJp35QTJ67Pwj5G2IO+TPLXr2i7W+7rOoY5Wgof8hm
tp/HeUArCROBqLQVJwHKMB+KlnS2fLa5IxHDi2iriKc2+xLh3dxVm9MS+F7vWroL
x09ssr724NhYXUrZOy1Vuct0vvOfn0NkEOJe/FJPl1a3RTUNuAPjg8uWS754TU9M
iukP/eW7h5tSUpX9L9m3DFuA1EBDb++BjHsov5hnJ4E/LWVey8szXLx6lm52ihey
xQaHekGbOQXpyfZRLwrCwpx8U8uHFihBW/YDazA3Sff5+yciKvg9ETJrLlN32k1t
ASqqcgLb7YMZVUiBygSiVliJfvXs5InW3BwdXDox2l7cWOp1ZCIWwmVwdSNiSoWw
UPDvVPDiWFtAH9XP/fvQlMA+NdeAR3xlu5o6MoTcKQJHwxiToRR9WVu4rJEGDlmn
Fcm9jWrWiDHQnDSY3VrNzWPVsi6Cwu5+dn9/m+jVimVl4/8uM5kDqkPV6OtkyuYb
5KPrAm6bNhspNfNlPDPXuV9qDbeks39RzMkuy5SWxL5vVOjJuLAlrhgKUGDR1hpp
HG8vaL0L1CsWfdMzaexzI6f+mKldeE+Cnp25NkeRQk8Uq7Y32ADSaYusCH3pNodR
nHrGZEGEKEF/Hluk6WPDqK4CYag9uOD2KCe3OxgNZtEogAuWa6u7gnm0nBAdZ0IG
IrXl+w3L4YtHE8mF38ZLDd1S/EwEwZisBdXT1gnN8wtAv4p08IsMnHk2O1LVyy8+
M/0jMgKSmEpCio/ehMvedqULCsWbmektKnClxmWhNSr+a9M6tDR8/EiOCDKTNbdC
0ktZdUUs41cLpSPSZGlO7IyO9W9qWfcw6Y3PcUa1ZLnFwSiBsCLhMmQANVkDkiIK
fxkXcuJMsnxQEQXUwBKrt41UFfMQIqxuqoVdVng0T3kHc8VtDAz4dbFfa2bAFlR1
V8h2Zi9P/7TAr7tPllfOZ/y2uG7Pi7GH1phYu7w2QsXCyH52UPCOV4y0AaFc23ZU
yx1n+G1yyvzwHn3iXuIMPjJMvMghQdGbTSRX41bJvzrFQcECaFlWuWkROX8mC32z
JfqDclcOQI6yH8l5owXHxkltUh/2ML/zX/DV8SLfp20ow1m+/jnYVUZKYHRHc8ym
YjsyjpIex85PnL3HDpDpVU3hlJcXMIPp/JipxMAqCIGCBwC5ON2byZnXUxkI3798
9f50dfMNz6cnigfbw1GM+zqGPwzedmQ14SgGS9G0Nxxzl6bb78Cq2fC6ExZTzkxS
pZOgGNVeuHZDwMZ0+d0AVY2mpfr3Dl7mqb7QiiW7gZTkEOpUB1K8DLzr1q9oRRrw
eSj4Efu52e4t/waoV/2hoyttMXnVgdaOiFSBxw2XSI0ErECVeTthWL65RR1aTrV8
n/lClNU1HfwD1NPVY3wA0doRDBOTbMSnPwr0XUspM4ZxOwDDPT8WHbx3dhpkFImL
oCe71VBULRXVNm825YC6e9mkWy9njex/nPLBjrw71gZU+Nb/n/sYSOPgct2uyvlA
aIjTYL6QBkxqAl0RaKb6LXjRpeBSqRTwXmZ+81fTONUNqNHmkgt/ruSV2RiWJ6Kq
v+5jM1ZQzCN5MPNbhiH3HSyiO5qcm7vk9td8OJbojcufXK5hcm6eQGRSFW6ZgshP
fY9EAf5LhJMwCTjz8I9U4UIcRR2U+NGmgzk/ESSC9q74OZtDpwZ7kRQ+tiIAKhKz
J0msU/GHrNCoOEdD71LNuwPz1GfEAa1Stpxlpf86LOPGdZSyz17x8HkDpZ34PIcD
ZFj0YbthGf9Mu6iaS1IDz+chzojcdFQ/7Z4Mbbb2Fos+LAS0FV6F4EEDait7sq9S
5S511wcEJCht0HahnTE+hw031FIqHIAzLB6LoT9hxp+tOXK/boVbLduYKvKLuq3i
W6+VcQfZQPoeWLWEkOQ6GVcxnK5Sy/di6tZjRT3VwPCPhGxN96FyX6a1COeGdJjV
MCsVPo3OCaFchfuc5KJOy4E01PfpYwIn0/X+G1Z7ukt2qWWMnU1I3DVw0WgPqdmx
cF2oycx77ifZYJrMvv3fWziqdiAqAYT4fqMRcWnl5F/mY8Jf/O/TImmvD+QlRiCP
TuPxCsMKV6RHnaPC8IKVdvq7QVH+mDMRQ/NaNbzXpf8LVmuU+ude2n1qRZ5NRPm6
QeVUGct2boXK7XF+LvRqUUaTnFEDyqYEa+j7ON0aPsdnxd2U9QWA5wpyGeyjZ8wW
jak64OkH4BQoUvHGu2qhMvSrRHgBS5xwEl/Vt14Za9Py2XhmssU+t0eUXlQrrep5
QowzrAdjDu0Zd35AIrzrIUNKd3ydDW8jfaLrYD+WwPiI0fyMwL8dkY7zhzJYyci2
wMJHpoHfCUe8GmXw9apuqw51fsCuOgXryyfckA9dxbC6lkoCLkikPOsk5b4oQM80
m/QvdoaxMVPZTEonPWrut+NHvpjDr7CtMqnzCSyVbtD1hOEytQxP+3SWgIgBbWa9
4E8CIPvvFHa3Ciq9GgHD/w22x7rPSg7e7IvggUtZIhNXkIsZYZASoC28YJvpXZm4
aRKYIN5BoV7+3heZ7BXSIkkLG5+GTy93o1ZdMZerfugMzHsk6r9kOQoII+d+BK0n
+hj4lQ+8lrX7S7Qb+Bm0I0VQm0TiHM5as3RWGvgXzRwtgezf8P4fU0OovSlp9bku
j+f3BmS3PxI6PyBk7ai/6shsRVle9NHxACLn0p7WObEfer6cjYO0rYJzlRbIRFFb
huYpWR2uJIeMum/+Isf2fX7/Z+XoUuUiVuWYEDUUWspk2IEi2Hyr9dssUHDiFJun
PEnk2M/Q+b16wiRcVspTe+6NPKI+uxr5ZsQzLYiLA2P1dQSHyYZzR5TXsBVdTgXJ
Ra0PnJr5XiTMIUkotvpehHVluhoVzicNVMSaoTd2ko2+tG4FBYAxKQKUvoiMwVRy
GJspIttZaDVUi20GjZUSRz21cRPLNU4TN8a8A4BUp9Tzq/Gu1+D4B2FzgFVQvLfJ
4nq1k/QqQchZAa0x8uU4rJc6ehF4GI4Ik0mmH0Xavrc/yGW96CEM8skbNBHU30EF
7LZ8Bu2X6f4i5EO5+l8GNVbk/apd2qRTHGTWBRrcFCKobG6MZs115NkoojMygyN/
ACp6dcLFTFKwx4J7mz45mkWOEBFzYD81t3VY2aiaEj2TQzYjeLvR581q00HB05u7
LFHNzkXkrNeuVxjdUrT6OPwv9FMr8SILfaHNOZnnaV90qWBcooCI5NvzlDe8W+tv
36kH9TrhdUEQbwzNxckX2G0MOYLE6MreYTjj6SvQCdmEKXWWbOjiw2q8zBgcVcZZ
r/mK+RK+9RYIytDU03EfcLOT74sHyCST+hde71CopfmLPmfZVy1GhYGHlkcCziLv
Vcv7ap3ELwjQVktmANUaVqlC5nTgk4nlYaEII68/Z2zIsLK1vu6WXGQ1FjO2C79V
9Umv16Af9AbHyQHiv4WM/vnkdorF+k4JSXxtso2xqGX0Z4ZfOuF8+NRChVqHzf9p
n4kx9dKXJoocB6XXtZcLNIt+g60t8Hb7/mjMfxGn+Yfy360SsLPQ9Ic2cQpV8NNN
9grif53QVR1UnT8SsIcPjbNrAlsgZgdRsg0JvBKOqZ8ttAFfWRNeLs8L8a8tTtjq
l4HvO1Xh6LL0HaEWNvpF/3l5p9cvhxee0c0HEM2uw+Kl9BKQyUGnU3bFzDSPnFW0
oCRd4hUyS2eTJELGYimiPV66woZc2dF788STFWkVva40XLlGFooHvWccLNTPvAlF
fekyIxZ/trLM5hKqGWpmATIsJvocFV6JfgKOobLWxXCrbuhB7ohLiM1o7C7ttAZB
Tjb/6vEEmE7hcGlLBHGtoGLQ0Pu4/EqFzk1Mji60KJsPI+LdubiO7tMeaxbGJMvj
M3DDAyNKZjMTMlijIL9AKUS5pdH7j15+B6gYopNUA+U8sua2qwv+GkB+haDEyPZ0
XaHYmt5ljfkb49wvImf/4w0MXRXDyPYfAkZ6+BzcUCRNjcnaFCo4+HEaj5gJe0lU
vNgW0jDh+RD6uuWJ/MtIKd+bWk1FAPVbdpfvYP0xOdZAv2oRv4qArJuVEDtpRO2G
u0r5Tr8bknJzbaxyR+7g9342Nys5Bvhh/6Cg56f8qMkgTGQ16ip20q4MmjdyJgJ6
T2nBE6BorYPeqE+9xg8ALEYW0DFKNZ/LqSudIG9jFaYt3JLXlNxsp7ZGHDSPwmWr
3RxTKSmMpIVB1udJOjxCAzv4yM73EyIr99L8RzTQiGWCnzPmeOhRWG9oMm8NJxye
hBKe2uSPAgbvf28uWExc9kAklt93VdSsohQPMRVvBIS/EkYlMohaJrWO8PQs4kXf
GV4BuX/aL4cLwqc1M3PyOiivMIMpnTaYGnftDZo4Bi6HTnP0k4MW+h7uD7wIPaNs
cO0gE069zHJq94meFICoW/TthZxlGGLjptcjzQ+hl8NL2dg+hsiQGzu8gan/MXdw
V3UMF8AmnozFyArlQ9/fkIPy6BXbGE4Ln3YQGHXHcYVyV8Asy5vbN0g9ITLC23w1
006JXcUm0r9c5a95TVa6+bRBcIANFriZPTPZjF0Hfb6PpAsPyuqFJegfrrMC1fgy
GNC24inSnNBfIPrkcn4S/dbhJ06XUICSIL57YWeMdiEuNAgSU7/MVtzL8CekCldH
ATwfbE4LUYCG8lWRdGdICuAlCuijIYGqBlHh7R5Jy4ETbrPWbfSOV/s8S9p1N8LK
CYP8i2fj+LsC5hy5GoBFOfEXvPly4gyTpNeb2nWQq1ERwX39vvol77UEz5NF2a30
qaoi2NuDT8gJJsv60sJMhPfNC9UpYvE86j0BVwQYfI8sI+lIjsoStYylqlF5Da+E
r8Ol0jxqCKJeUdqq50G8vbBjdo4eI7NdibLblC5SjFERR0rrlzDSW20HPtHIo4eV
3ckaYx7rq/K1wv36Vc9oz75uMhVkWilpD0L1wrqalo7VJ8YxL3QkExjY/m7E9ilC
2WcSB4YHIPAlrmj++ZLH3rkIfzTLTPeem5M5l8p2swEd9v9g7iIGmSVLLZ69CDH5
XIWGWpfqFU1zVmiuch5/OuJ2JZnxX+PBmHogfO7WMw+s+PGTYfYaRF8nGyhhbbVJ
FlaYt6bgT38aUGwOgQF+nfvG1Cu1hm8nPtoIxUimOx7Bb8Zv1COZntNk4hHmZ0Ae
NLIWfCMDJwLLDIUcz7PABEtmu6WuTyCUkGM1PyM5v6oEQ21bNAxj6iwbLQLN4FgY
adJ/obxk2PSTJAJE1L8uIN6EgPpq9uE/Z4+R733hNepvBysB/fUaVb0WS1s2UQ9x
/LYTFN6S2sshEYWbpq//3q2y0X31x0DwgQFvf/ICvcitCiI7DHupGd4txgfkjPt7
nvQhTFv32GYcJZ9XO7rxlc99b+NDckUXlRHRbppxyDRbeg2itCk82ByU7jyW6ufl
dW2mEctMftZBEx+uC+8p7OVz3NIGAOb6jNPd18n8PuHqDUEZUMfwdUH3049o8IuU
xiakg97V3WqEhBT1aiZIcGms1MtnGQvzJ1f5MjylSUEqnODb9eEyzTd2WA04DF0M
bIHHGfJ6ZRwIkuSGS8rKM2gxPKpBjeCaiAmssSOjEXJU3JDre6oEHqogJI1AOoCn
/N4vPcftbQNccwYW11owzZA4t1BLoG+1IgFkWlLNxD8ETIrdbCOfiaXGRX6VYP2Z
rfb9blSYeTBPTBPEYWlHwTYmnGf60sExMQ9kR1wTNqADkKw/trPYAtps9K01M2fO
ghmtf04a5kly7lemjzF3uAqDFJQ0CXT0yrBIAFL0T0sfGjFGQ3q4uNZTWi6SYDQB
jpU+CgC1QHM2I0seYGxNQ6SkxOj9CkW1bjLLmcBa83JczmRJAiFH3kxY8ulavfMa
6SUOW6mn1V55X+oq1TTb5lh0IgjxrcYXnWueutHxHCK3EN7WEJRy0OoXHcGgnx8x
TL1K0AGQf0nMZprLxJDI58zlsOiQMPPj01bIqDea1gQvW8anxdew7ascPAjZFigf
wIhEWjIQuLjU/f1s3xUacyDwxJYUNkZ7rml9rrvNH1bsI2jBFfG0xbEHGEnASysJ
ML4XMDnHn9XkqDgHMMfo6ELA7a3IImWLNwKGy4bTBssr87EZRsiunxxaL1Pv3zjO
s4aAdaOkdhp6/NpvwHUBheYDKFzVuJL1X5NVqGo2m2xBoNXrj4TE5arbe6XhHhUV
/UNDOhoZT0jKUupSROFlFz/bDOx5OkkvArlLsAlor61YleBG5U+m2zvAfTDQA5kl
3RL+GqpkrdEIUGOYDHVK7mme184AmegCAZfagzo555WukAgkagAUYAzXgz496Y5j
Mqb8QWVJxl6+nd/XrmbGe0xaY7OGd5c6GlC1vwpRushY1AQRewL22QtAgR5z1qVJ
mxrm/As247D0kECBI1UnqoirHBDSkBf4GMwxYSlEJNgiirZiVIpbq4OnTS6fgDxX
Z7uQdoU8GMj/5UdbfkS22DeJ0owi/Vqdl6xulz3L1ak4vzSDj+gvmyCIoXaJ6tUc
TdsymUyPAMsghAaKMoYTHwYklou+n6kdQoluLuBEva736pqyNm9aPkZLvpPNfG1u
jNEHcGGxvjMyZz3ATGt9azyrUSUGi1qr5L08Kf3+lzt0uBzToqcBALP/Bsy+aP0D
4MJHpb4lsHxhPCWVNIWfSV6Qut1/Bf233Ek1heZ8PYGhtj3TltWgwWiccdUVPAB1
kMcp7Z8YWmqdKYw+6046bf2MS6QZgOqU4l9dZVG/GD8u5ZkAO8mHJni85jB3VOK7
TQRiS3XKmKGEvNJdt3sL8hmw9/HssHHy9PUhd7unjwAf57B63stMdHOnazpMfm/y
y6+kXogqZENM7bTcYBv9pPwDU6Te+fW0mRIBaequnKL1OUPCUmZX8T2PZLWuE90G
IfbVAoz56lWD6Gow8SwL8jamZZDXTWQlQu+L+UfuZbadqCBFecRTz2ObJqnIPIn4
S/hWPhAYD0/5Y5qXIJgfSHmWvIQ2X+dObsOPNUDii3NJe22FphqUPzevYjCsO9m/
BWHHP8g1F81EfIWGfYhz6DToCFOQ6gVGr72BcfC2FCGZtKvW9F7xcqTN34dk8Tob
tK1xTIR1IUqyUesUWTpY8IK6N2Myxn+2Ym7eXmHkT07MwUTdDNStWRrClOI8ITw1
ih9JkAwGetTORcpYEGfUcRyt8yxT7vYLn5QwBj3z6j35luZT4ewqPIJWL4PYlshY
qqrS4HDQAahKX9GpMILoNOEqoyPiKo8d3LcHj1JVsVy6qEv2D26q33bsy14cVQn3
cIG9L2kNQ108TwEEljDiuq2K7W/PlZoyANlK9tHFtILYGkZB1sLvqlWlnGNVsnV/
DzKjIPNco5zm1eDAcKhMxNmcxxr1MASw7BYpN1P9Z+T3RwoJXpuTqW6PYSVkOMhf
OGjd9n1hre9gk9g9CVhcC3EA7mblnHr8G2KJ0Q3iJ3aiEWpgvxdYIjbR5xjlVumf
INsPjAK6C9+VP2dOIqEfSmj6YC/d7FNBRQ1eGl00Z902/X0OK1aqD41PvrG3aJuO
3t7j3rwz66BNsYu3a3xK1gMzV/2PCDmT8020CKLPcGbvA7+iNLTFZ1OUcOWUiUUu
PPysQJAvQ/Dfggf/xJ1MC54K6FSldIl3a19PYD6Y78w7kv2P3S3LCDG8u5DJ6mkP
7e7bKCYXC4lw2J0/V+LbxRNOS8U1d4IMXRLlC88zsKlEXc96/Wrw3AiALzcZB56N
6k8959j7wfXQ95r6IJBWKdZyjE06EIBGbVsIsU+xOt5KoqW58T+UnAd+riBJ1QqE
vUjbr31L2aVKyBXJmILCKPG4TKU9MVkziGnB4zClFmDIQiLowHS8/IzhF8GZI1Gb
L0xr1/JdOJBVABiYIQStJaTMfhh0udaSxDkxhrBFwQOCVGpljVjI1FjzUDVZI2SC
xKBBhlT2YwprOTC2OM6VjP/bRKS+sFY8JDKlmSGsSgNbmvhwJiKC8xjRBxz+g5B0
hTeybxo9lHCbT2xVRPl+Zctx6MT6gWj9DCM+vc+ud49hinSvO/yqDCK17qgffTNS
AEz3q6+7HO2lyK9Qmyndzvfic+DI5JxRGd8pqE0UYL1CPXudHG+utqh/bZSt/Npr
lSuQnX+TdqPtu1TCL5fONcrzQkbh3fPRM0MWO5OPx4Y5a+eg+OHsh8FnZwwmkbw0
WP25+tLZCFBhZc1VNKZIEOgKq8D7DYIfxbi6pyy/hHUT5fOzWjnTdKMTsHPr519Q
TC0WCJAWDxKeDdJ5W+10XdrgADBeb9EiY71cyzpiwQtacmMgnZRarN314GTNql9W
hXVI83CeWDt4rB3vMD55lvS0bbM50DwA/GApv0Mn1u+X5GXPi7UFHJ6MxEzlg+qL
1rX+xOgj8OoVJv4cHCQFVZ6GYdxa8b8h7xD9WIWP3JcGQJ6gzaMdDl4AxGHYrVVe
RjFl51juZCcm4DLvLR8rz0OWW641cqz8chy8wR9uMpibCXHZQw3+0TbEwjcqPX0W
SDIMdo33BMfFS0p66z8Z47hZP2lbALwknL8KcR31SNMr/EV43+lR9ScfPErZJrtc
trhVy8Lf8lwW+SqwPEkoGW6eV6UjuucvyHXwHvGS8nHhIHY/vFayCoi9W4amfvSA
ZWjfM1qcBSf5GHg78EmW4iMC3c+4ygPOKID0SB4sIlfBQVm4bezW+jzKfxGnDjzt
RN0628UpNmM7RKlahqpAvAvsN6JnbVh/1RAZIpZYBhd8oPAXqVsrm1aposKseAHf
+06i7ZCMVqDQiiwEGr3slOrayv6ADFAZimFu+ptLN/FY0c56+kUBkVJtZbt30oDT
B823fBFlahrUsfaiLLTqHGNo1v73LEeL+28bhbLqfD4J3UVJAE+U7muPPnq//j4S
YSxcjFGCW3RZu3pAp3RJiPXqA2zUanr9eD+c97MsvTXd3D6OTJJ/OTeREHHgETjj
e5SRiW9zNtsn3e57uDYNCusNj8RpJi+ph12R+3xY+hKI+arjzFUHACPZ4KFiEPr9
LQJbdIHYuwfY+FvTap5DaGU94IOLodWBqm22r5+Ssh024js54HDwBTBLnpEWwo2m
+06JvbL5Avdu6EJ28xyjf+w2Cj593SaApMT9lb6I6k+P/EZvskzhqyrnBmj/tUoI
fRdsIh3aO8El1n6SkMfPh+uJNDbfhPHuHiiypeM1Q22secO0n0zq8I0YKeaz+f6r
ls/inGN8u0+rnLciuwpmPbBt4cIxVjZ2ae67AfBSQ2JNPVYJSozi1TkobysHixMJ
5lWZi5lWfH7vcKmrprZH5QrHoEPSUYUfpsZ5fMFCtVclLKLdyU6HtIyMadg5KGXa
D11hyiN7aFAZhXMKUaUz98LBUDEew2MnGeA52AoJxJaeVFmyZOTnyl3Iu+gdMhVN
0hgi0eKcPZYP6MRxAG3M4u3l2GC6ZxdSm3icp1uylygfehEV8MOcJW9KwYiG6777
GSqJEW6GFNAtMIiUNLykWeEFlv4tbofomzXb69+thWuVSSpPJLL5KwwjPZORS0vf
Q8rKLIFzQPV8V/2K1ZE9/llirsSvFj3U3SyHMrCbL7b01vte8zfFMCHpy5VYvqCw
nvaGZxiU8N/t8PQK6hMXdm8AsKTEqzkdzZm5HklSJcBvIm3KEYeTes2VP4W0rOtO
H9U9swtX0WuSyr0rXL4JxFK0avxUad07Ig9n7Ho3PjCKITCJivpQ0ZXFTYBpLxnj
dI4RC1V3zlkXR5xD7maDNgBIuKQ9ahCNTW7+PBWSiIbUsookYFkhZNTo4TFhf1Vi
iwzf7JENl/td2ireD3dvMFh5QXyaNfQkx/y22TvYHAk/dHTdIpL3FL4NTpvCb3bM
1GqeUPyRFCDTi2QIi8YyvCN7I7Rl1goCMDZcAwyGU5+xkWOpec8mJdVZXV7d3nqp
sGrvGUJio4nj2S+pYdm1oKd2NEPoHVwZf9493CLLsn5aQjW6GY54KQdgO3VDX/Mr
8+C7fP0999NpBDch8LMyWKqW1EPbUGrHZp3UDVU2ySfyA+FtJTV971sKWHkF3WLV
a15KUaShXJa8iBM6+JSJ3+0tgLAURlyxbyN4RMnbySIq5mYBO3yqOiQQ1ssaV2F6
I/WzqxlXt/tgv72izf/ysqRymO/sQz6/1tY8r7axiYne7p9l5gy5V04vKktqXOal
AKn31rXBbMMfhJCSytvvNIXUzSjpEps5OYxF12bck0eryYP6G9aOQlFlpKRzc4AO
W0ehIGP9QVrPI2O0BkP8kGXLzMvuTLYX17Opmg4VKSUQRZE2k5VVHlJBSh/ZSgbF
QZYwHS+GUNAsdYyXCaz1kxBfr6fXEOgN7G9xO6lDIsiIuyEgsy2eootDuNHIR28I
+pDpHLoTAKY324rD/PN7ISzLzi5y8w9/UJpX9gbsblWjcVP7Lz2TVA9A/9s5hX5t
ZVNWWexKZHFYU0/nOq33P5qJbAdJZp+kDSv3h9kdFQzlMI8ELgt5u6rzR9WtnxeE
V9RhpQ7//ZGfmlz9CEb07TT5n8mOgvgaSAGqr+kle6bqbFisv4yfHuB88UPr/wv3
ZQFDOUFiQ7H8UqbNz7mhJu7ue0JcsE7yqiHHyfqzXEeOY+/M9uqAzT405aVqbiDH
/1tLiUSBNlxHt9eXm0uB+zvc2wIKRXPS2CazRAVB7JwzF74tnfv0MLt6iL5HATOG
7lso08B1XZHuis5lPhlQak1K6wmYwKlkkuQkuU13jntcSf3ysCWPkAFmeNl3BcjF
VYbphHeq+OlpZs7MtiCtPQA5UAC6lz5yMOhdtLQao1H6BRlzniB8WJwSbDTxKHIA
ROHzglM2qYHNNuvzMVHSZth+3rFbova8IP/yQUKKUl+HwTiFHBvmFWnpZYXfBnDV
zYKt6KGjUTYARI9PoDbgHyCUKiMrS+rf5K7ucEXGEXzp5S0FGZ68B0B1tXREfgdg
wGJmlQcNa2aP2J7js1LohiYRzRZTz5ms556tGDU2vjy39tDaQRo9Gdqj0eoikKy5
jSKOpZCRpEXx8dtz4d1Frak1DBAGCOGXLMej2KiMBJ80J/wwODSFjgXPuR48dcHf
a1FhIFg1GotoM2mFU8m0xrNvN1c7G15bsIuvag3p2m27S5aF1nrLazI6tlyu//xE
arKysMLgRz/SEpRFh4VDdF0jvM3x1XcJ2oi0XMSG3WZjoBxGP277hQuEJ1XqX20u
zCy4b2S+XbQKQisN9UyGjHY/A2jMYcqo1pHT/1xJAkJY6Yov+3+2hGuN2MrwGv1P
1cgiQWnnXX2UQaih4tQX0XIzxLJwtdZuFsgcRCAwZFqyt52ahB1p2VGN5yBWrtHz
FNsob+sNSwjuX2Qt/cGt5Y0vn87cQY4zAxDHI+3CKvM5TJeDh9vzUCV0d5cI5+J3
leQVZVOWCJ+6AxT0Vh1fssCcylup4PT1MMNd9eFjFkpqmyJDwnFRBmdPMrzXYV5/
KljSPc64jpAARd1VNV8wNhWemcUyRq6WweA+A9O1Ohdh79VcNzONM3K5sOsMBiH6
dCkhzMCfYzkywWXKxoqMDhWw4G5xHkmSx3MuDaABOU1fgn/Dxwe3hpO63A6YFOkn
Qh2qLrtwxyOO8NXjqNk/lQIf8xK0pfr7rSS9xcmT0PMy9+r2wTRqYJNCWfhLdCQZ
zCm/t5UORnpMvvMuJjpvdow7NdYVbKrpNHoZx2MK2n6wIXCtL+dV8MIShNJ8q36e
2S1agdgtjWoV9aLgQGPd2GY6tTI5RCjf3JJVccsmV2YNwwyCIn92P+yK8r0r+to6
7VmGB4myX8yJIT9fEm/1V23nTis47sVcslCw3ja2FDu4AkjxMVfEqwFOFGTAuLmz
H/VFo4FphLpAiAtK0tpaxhOCQ8wSeKIOCdGP23eEjqFyc+fjmFptr17yaay7J7Vz
/YzX4hKQBH2F4oGQ0VcC3vRrJeTIt5h3dsoapICubOhfmkWAVYfmG4+kxqWzHQF4
znUlGU9m4AJzo76EXtd+4n9sQsJZEqMPgZK94V5ynLWakTempOFuCjE5neMw5GPW
oMybRe4OQ3lCeV6Gx5lJK4i/jCJ5O9fcIppFoFy7Z6N9riTwCEo42uoVDsCjMUVV
mVu8RYZjbQpTbf8/Jf8BGVQhf/oxNy4i6Ol/g2fr0Lz3CQoe3d1zOT2fE9VCh8lx
OVUUUGrMIFdl/m5/XZYau/uxkGTE3hMRu7Sj9GWfkRUX5ZSHSbb5Su0ERH9FPKAy
vGNCqXo1gq4TWcrJzsMlk73wlnsbR6Vr/bYKaYNiJ84UxnVKx8AtvPkVjGXoCNrs
5wejpu5rZGW1QySj7aS+8hPYIoSHCO18gfadwK8JiyzGsEhjov039GnrXlav+sGR
+yKGyc0jdFYTgitCiAZjIdWszdSZMMfD+uYKADXm0khFZ1ATL/wMwEcUT9SJ5YR4
0WxZOC5cCL8d55vaXNLrrCM+NybM6fLa3EL/XjbuqS2Hq3gvxLaDOLVWgHQcI0i/
o7DrguPzHnrClyx+ObPP+xUQrLUWVNa4jtldgIebQngKlqmIz7EyZzEjd47Xx2YJ
THg65JLfZljizGX1SeZZbENYkKcvSxn3BlL60I8ooCn1daDItPbi/XcfS1xRpsZ8
89Hm618/yqQmBxMcaqSLWuSnix77TH8Krh9tggcbHzAdGw/NUoK6s4NR6/N7eFYj
Pywk7FjFfThhzaGDbeYX22LFvCv3+bwqQ4MGfQ0RFdVKnV/FnAnzhRmQp013SAVJ
qGJQRSjLfYURRAQ941ZsmIuvMd0BJHL+kh9uzaCExC+KlEMzCZ+9o90MuDl195Il
eseKCDImxl+1HrSesIIn/UZUyF/cLdIh9JcC1hg5T2nQzHzwUjJp0JW7C7JxpbIS
DOv9lnrDLW7rlXQjnJb7u5cq6yTVqrXMtw05M7Bs5Kt1b6XVlBFRFPmgtrEDkKUd
by/HqMtqpopT083+9yN6J5Ps8ugl3FMn4Zt27yiPhlTOXZVXatQjCZnehW/OmYjn
HUqGiyj479yDEfsbEU7CqSaNgs1uHuEPRasE2yGA2JvVYf/GqXGIwK+LXI/PDleA
bgMdaNNnKUM01GLvYUz8f0PWFq6Hye3FC7p2jt1FuhYp1EKVEORGnMONzXTD7wQY
qbqWVe2sTe+VmEW/ybU9eYaV3C55jrvLxHKAu3dv1zZ9PQBjJmmrT7JBRY1ASYae
BjKMxE/1MiRXQSxs19k5DeOakbBX1KS5JDMoIXCxU1TSA9NrZHKgSsG0p7oLmf3a
ZtZlV8V3fEd+G1pg73YhcQ26BzmEteyoAD+22SP7nfXrb1fhgA0tEfNym5IcFRlF
50zrZuZBfQKee8yd1oH+iyxdt+wg8yGJthKvw8s6jj8Gkitau2+dr4DNoh0e0jDz
8cdNvh+FoBQ91fG0P7diIgrVRM3bRaJJz7fvAparHBOgSCct0SlHW7HCtoa6NiQD
TXdb7JH1+z7RWfJ7lhgKUoUTEY5jyzRq9Gvez6Ptq7nmZsoKWYmghBDR7cGEmp5b
CnQvbzMrkeHD2ijL+HAxgWnrTJ+nGj3LD3i0WUYPfKgfCnrx0EcH0CPA60zOMSTW
bgwbjAZlo8ojjrxDOrCcOE4HWCWlxwl496sd8LN5Gk9wEvN8y2KkjNYBPpM1DUgA
Frgs7d+NFCQ11XtkaA3R6BJoawtLjPU9dGT647WXz13xU5o8yp1FFITM865pb9Ly
ZetiC3A3dHpv+VLhQwhcGxsejUdN3dxowu/ruQw/lbuhIml3Uscn+nnS3AFNdm7w
Nx/cAvF8JZbYc2NvhL5ITCmx5zvVHiMDiCkM3uwINu37f/y/12biz+Oe6SiyOrXG
ynTLC38g7Wd+/no7BLi9rPCnicAT8pXprkQRrfbpEpaHyUdj4pavuWz5/LOy8YJ+
XvLMkZvd0db7xGlpRCyJsRem8sbnaFRalaGhbcZIgwJfKEgtUXO52jHsFMJqdf2z
v+GrfIihsI6Bq9pR56CcoAd6DDDkifVqOI7VAbKkwnAU+JgtIHowaNm+PQ53VIXn
ZIKkGkLmz9DiLMuWxBZZGf2HPm1OzXa6aOXb4G5fwiZwTeEK6AKh0IzdG9EiIWti
cHf/7OjJDPVSWsLpz5Crwi+QLex8wf3ng+6OJ4ZloNg0RWsodSLp0kJ8rvoiO6+3
7s9szWIFuaGwWuXf6q1cNESWIqyMtXAyctmOohY7eHczRWx+bORwPnqig1vOXNla
tTnuYYnKNYgitp5KDueWu132RulA90dJb1QmiQLYGbcL3JGo3vzHsAnJozB0zASF
jR+sSBCqTKQQ1PVkB/vlNb0DB2ICPw5B9SmOYoTLnBd9+V0rgmqaR0yp3drIpaHh
vtC/89kTltkwR1P+AqNV+x7yoBgf0pyM+ezE3kgXMKP4whxGZaqN35tMPPOOuasB
6evffqz4bv7Cfjar78VdGwgqiq7yOsa9r6aYO5zckv3iwHoW54hur3dkDUrNBh19
f56DOzCHyoKO49imqS6LsFxjPfMnHTob2fFzlUk7cLWgSeDeixuZCFx5SvMuWyJb
vxNNQYU0uCwtroN7EJKprkIymFFZImRpDUZN8VfInBcgJ19rBYmM8gYSdFBgsfKc
n+P2K2e4mNywcjKbPjKJ8Tbtebf+s8Y/cgm8oKm+ZhM40oIhWg6Vi6OPL9BYfOOt
DS1TcH3UPPPdCKliDO+YOkbu6uJAjqjQHgW5BiLpvLEXiWi8tN6cM8+WPE8mNZlR
EarnTFYzSsUS0XqWcP58xYtSKZBqOgonaOJ+WH+qOT9/fIs042+5g/xjcaMA84nB
EnYiBw4AOtlRzO03NPT+oGLAVpXixndYpqDecH1tTXRz8mOp25wKuPjcKnCnhEP0
lJZuGEd8kMiXuMFXy9DBtVEUVQLtfaFI5ZYuI5OkzcqMx2zcbXb2tV6RpgVdmGBh
yMMFxLfYbdFIKxJLPOY/W9xEM+w4MfO9OXpuipM5bKouyNPatNIRQWXTxBiZ3LyK
la++ceeN4ZqsxgCb/pl8c6OgU5zVYzGbj6Ghr47ZmXq8wl+TKIPYtHGraDwFG7O1
oaPOD0Jpq2B8MUXjal6HSqXgfUBMg4Ttm1os8oEUajfeFh5ryDhgWI+35m+nLg+q
lO3rW+QOPY5BIWj+XrHlK74njNLtS5PSUws9+kSEWmfDGmiJd8ifJbA78V9qkICf
5kqJ6fFvvOcnbhJNmAHfcb9OMak6aykH2jJdn0Lgx4AYQ/3OTq9DPb6MPpMcq0a7
Xnff8ePGCtCt+S1mDVJy1FzyyI5AJOPk8yjAlhIY1eEgfNaeHfCrDHMWEA8hPiNI
56FciLfWtDgcmafsEA4AWU1ySrh7hLNze6nE/QMsW6OCGdvsesVdbdemqLkcQIYq
F75k7lr5Z92SPutpH2zh4BYiCN+idCrYQLmemw6DfMxHgwYNVIcMzYzbjrJ+GrMy
teQbNRXAvFrSVbWVDXM8sMmTmqOcEPMzxgs+8TeFMRYvUkEe+XOTYI5oC2BhOYBE
NhXiiwl1+DSwtdFXX3lQuHXMOVaK0TWrrR+2uTCpRXwJlI8c3ktATFKJWwlHKlPy
joaPnYHFpqEDdk8j+d/RfgIXw02isOe3JQGt3cK1K1UZre2mv1wZYpdc3rPWmu58
4wWaPMngfdEO7fyC7FAStqIGcwPwroWLuC0DfOvGZC4Lrc/eupTUAfvWH/uzmx+P
QdL8JLnovIqPbPQzzfguQ3EP4dt/glEIXAxEkh2INWP6Y8tXoGbLO6WXfhxre4az
QHEG6WTYIAaFcVv9JjRsdpE9YuUqMMXKjmz1ArCuxzflWHO9SqiTCHdPHY3t5NOs
IibvGfwDryZks2OCEA9zAvLZoO3Dio3sLULbQInr/kJUV7Wp6JmP824BJagd7Yon
lEb+7FB0Web9rGB9IHXvYsZYgzDsz0A4shkH3uhdZ7m6+/2WPEYDoAV8ETd0Qnwj
L4RdB598B4OzVqR+wd9wKcg2GhcutHZGylpojpzHn0VK5fJuQoP6kpdgVrEqWwLz
h6pc/pibtfuM/6Zaxrl5LJ2KTje88vWPah0OvF/2ot6L0x1E7Ch7jNYKSX4fqoxo
476aGiCLxMAJIgbQanjBk6/4nQye/iO+TcbpBgOMEM7/zrL14KopOkoejUaPscoU
Kz156AEArbUOQ6g0CEk+eDjAKN6ML/6Q3kYYxZokXweIUpVJahlPgXFfOkJUrvts
h889n9YS063DTuNKLA9itZW4WVR0M31q56lc04ABxxeUwKd/k35KUPfJ1EHRdjdy
4dZSKWFuRgg4BPAHfoxOygJpWvPobZLHb8sHNNo/F9pikC51qrLxo+BZ9eNq+oVz
hokHf5a8euY3DZeP8zdgUhqJPsPnp5JSxUX8D0Zwy3k4z0CHFltB9o8RTZt6ycTA
24U9QdZSs+jFPkDKoTqU1RobZ/NR+76NsqAl/HjwWHERAL/7BjmpGD4cLBOR8Kma
1+KeWsEbP5DH8/yC2V+nbbbrxCwsXG/tYvbsO6z5j1P+ujn0k8IVSnL8BNSs9z8I
w+mooCJ9Wtn8UCPD7XwuYf/rswEBpTN9Ids9oz7cYi5LOcHDzgIbNaKqmLf3kOyp
XCyqsniaO4GfbcwyWrnT9VwyedB71xC5LzsuwHXVmKW5HPfS4DxJgqMUOsJ8EmCD
LlMmMMUk5oxnYPZ0K3GmHDgHUENYO//qtk++bdTGdcK+Ekerv04K00OCGTVNsxep
BqchqXXVnTXeROvtx5/LRKLZz3gRtqgKa/fGBcdjtITnJChqcXc34anWdQ6MOrVR
hTVTiMQjRIoFVBQw5E417Lp0ZW4faXpAB1nO9AVZXQlrmH7AAQXPoPc+wtSpdayg
5o/bPtvhiSAkiAvf1tfFqzv+XylqnGBHz8E6tYeQmnV1ey31sk9ndpO4utgyqGJ6
5JjJnQYBn7cfX7b2utCSVhAyHw9RePf+o+JjHPC2XQ/B2amuXeipLsk220BvXYtQ
ylXxoYvOjTE2x/2nQ/MsKXo5sFd8fS5WPzfngxOpYTWq5zZWYw0gZWruaefUGUkr
+Z0xe09rqZlAI115C0K3MEv5YPu0AGIFBQAPa/RJ0ysdSLCbqrDyS5VZSmabjBU4
BFf7BCpZAY/9OTzHaz+fq+KGXX/x2IIwi8SgLpnKCXculTIcHoIu+f3akujRakzv
KlN6CvKZYNM7XwcX7f0TqasU9yHbCnV+VbGw+HLHbCC7YfwfopnRAB755wyjWEMC
KXMNoWM0Ak9svCCqLVI17x/iBi5WNg5qOpQW4kMACOjeegWF6Ly8xyGhHoQx4ZD+
oiMyn1Meq35WMj6iWI5eU6JngxElQ72eQWuOnIum/dQkxQ+lSW82GzYTaZ8xsSZ0
je7zjeECQxGMbEIQbMJfAWb5a8r4S5qQzHf5Ilf8uXbN3QSC2A73UpF757DwF3of
C1q4YMyfL6oNjDwU8gdCNsoIZTsq1oxzhEwHHBx5P9JcxbmTj99hdfd+I+p68/KC
5Yc4vgYbKpxX3VtnH/rz5uLElgUbTksYPCagy1Rg0WDrfLzLBClRcWHgt5yKSi5P
yH732l1lAz22s4hDzNqe0ZJxUWzamE1jGAMfstGG6WjW32QyaKUr866u7Zn1eoqK
qzz7tRjcDE9AR4RgKzyRrkHu/XOj4xtdqb8HIQAbq1stUbXRjGva1FoSVrHTpW55
HqiHn+fXWRg9GANTwKvnnAtzvCZ5+1ZVnzCxR4mWs//OMMs7IHD01Lbk7c4XhZ7f
DYvrKcWLgy+KAG8rUv315aO1lJZmPI4aUU923EQd7P8N51urQljTO8WJA1CQnklc
D5/lcv9li92ThR74ylxrI7q5hMyQYNa5pwEzoiIlfCG9AfiNKStrizC71NdGoC19
3Q4OD7ntI5vFrt+SBHbQOhxQeM1rcpUtpzuvt04iQWZETUi+MlMHJpExVafo6lpF
MaCqEZ2iqC69t3kjUwigWtdLxOynjg51AWuQ2YJkF7TyYCczFunxlbZ64rcHgRS/
iBWTYgbgZFu97bM+80x4PkK8wExuVooCDeF4pe5hnetEzBd3L52VWuuDPfkS5nig
uKrFVLhhY+zOIR9g/bzZeM+knSVi9NkZRh3mLzs8twGm3wPd8ZCYYSKi70jmtYPE
DN1Ahts7CYg6aOu+eJ9GNGOVRzGPQ64q6fSDwMRoCDLE3ZfR6MHWuxGh5GraQNLd
+9veRHKZKy2YIt/tzDNu+tJBFOFVw3F+mCMXLdW5sEfwKTL+pZQYRjvpgtgd4HMm
DY78umfXTONwPPBp7f5wl28lE8h/4ijVbqJA0JttQObMniQPoRvZGqbkI+tZDtgJ
SQ97DCCKx7AV4j5KWGUsKKLWWqjUKc9mimKZj89iSIMtiH+K2DRbspanNzIQCdQV
ZJPbaPrMCsJR73OckdymS243qiVZpoz5u3D4zSzC3M75QzB6JCekBQInKBFHqa5e
dnY1BdKm3QTbVdUjI6sLzQb5frM1ctqMjdiwXqI+o0JHUBhFvE86syH++AFryQrJ
MoVP079mPMCIPaaLq6gtOE10dsFSyw5NEu6g5y0nmPsT1L2JkQecMy5b+WMhvBns
+saJykZOfRFaxboUAEPbnUPYWjul89XdfKZFKAIkfGX48mn/NTRDyATkAhGHTX9c
aSKvPtWMWBlSJKPgpvAiP/Em/0+n3LpCUgLBC2SpGczABOKux8YyKjMVBpP6jsAm
qXp6AOOJCkL9BnpPjgqUdkY1W5UH6OsPHlFfsQRy5daGv+sdg5VouzDLj8abElFd
d+7WLu/gED6tg1QiAyVN8jg+H4/X+E+fspl3CGR4Yf6c0922UXjvGsI67mnHAlEX
GjwZ2EzxpEZNqgvClYOxz2bjUNNN3DBGxMrFWdjVsvr+vSRXj1GAWcXYv/LZnHPK
6DXILaAN4mfQkSlLSZ2mp3iJVniiRfeo86DDn/C2YGxqBUJSQ2RXFUvxCmbMpuh8
xA3CNCrajqXvULqbCnRyNT3PNTspd/WjWReATAdBB0KIXsfnCQk/xfxiGI16pOrq
nTqdwJDJcqo34fzJsY0tJKhdwubEaXt662Q9zgtkLejQfop0BrdSxjbR0ZQheK97
eKoS7AQ/+r8as8szPq5MWGnZC/68nCQ0jywgtI9W/e+2svH+tEsBFotVj7mb1JwM
0E8FdZJx8A7HEoXUfzvjt67GY4rxsdYS42lMaXcHjPTumc4GikUKXuLiYgK/lrER
KPxvnMLL2MceUsh419pCY7KTQUu9WfUDS9mY7UFpc/eW++6msvj+iEIn/HYWPpH3
JOgSGZBGSxhWdmHMJDsf+W/q1F41q6/oEoy1DBou5L9QGKThnIh4yPDCczevOMVe
+9fTo6bUejyOpwgwFQkyGpq2jyqcSW9f+fxtR9SpVYRP7oKC1hknV9IRG/6MDu64
qyvPUNlqAEt98WEP/visiyNerGXGgUJZYZmOI5G00Iy4ucGvJWFiG5PnR8Uwqu9F
XlTuc+OboMmDJNym/BxznT5LqGw4lzEidnXjiqepvt5Ihkp3JLfTyOzO05T+vA5Y
6avqZ2b5ooE/dLzKIdMb53gUhri9IH+1fmfo8Trx+7Dz6Y2vmS74UZcvlGwbODOS
oQbEikTQaU3+YRGnKUD/xGsy4cbf2Vr7BE7LC6biUYvOPilrQ05cJgM5cR16r/tC
rRIWw9DB+VJ4QcUGxbpm/HG5E2Tyzc5Qh4obghurzikQGvO2yEutNplRWQxjvn2m
OstY2ZlV8BjcugUVldZRi14FjeuzwQdlN06RET5KtzTz7XeVu39CsD0bG+4kxNMD
snuEPuoO9tqhzdYzB+BXYfS0Z0H7bYAcTDhv5YbRZVL2xFPu6IUkTNSP91qY2TT8
Z2l8awn1xPbrAemv/OdLAaDO9MCEzIGWsv2gzR986Wq3iR5o45KYOFPy436zpiZ8
D5nLwBfRqBpAM7rA066Ohp38tyo+OgtHDDIZiIOrj/SVUjdk/Dmy1PGrbHRyVIor
0AESypbGuAr34SRWIK4kI1xFq74BzxtIH+5KviJ2L3JWYDvT2PsJiAsK62Kx6wll
VWVAm8+yiuKhC3QHK0Q+QnxmjuOjsD2OtvI969mdbU4l+PlYAy674q/4bOuMW/bD
7oLfuu59v9zR9e5yfOl85qWmRdPpzuRnULNsZjwNnlEICbRTOC5gFNfD4rk680Wt
p7pgBPAsUrT7/SZUGlowQM04K9TJE6n/4R4OSb4ImOXqd9shqbCOkRwjcGk3wCcH
Nobv5X4Y3xHH6AEC0Puq593RCAgKGvXjheVuPg/vf5rrTEO4sVtB46I4qnwbrb2u
yT2ksneeuaRfnLnmtIQMCFk12dBfh+A5MJcgwekpuTAFTP1woLNVK8cT8iqC7ZKW
AE4HCWz4aDsWilrr7gnN4CmiR8c/lvmKK37J4pqulDvQNQQFL1NykoFJG1Q3sSMY
8CAed2ZHbaeXJq+LA7kM27cJmTEhog9rEfu9fHed8B40o91+RAK/eu5EWAWISrjj
a3QY9AIxC1iBCUI12vvcvieXHOCebYGWftElu7zchj3oh4gmARf9t681/pHVwh2o
6cUPyiTU6viX0LFmFpKYvxZna5Hd8RuyL9BwfMdoFeEE6HSEorKoR5PItQ/82bCC
PkjkOt08NygGUvBubnY4xpZ8l3bN6L+bVSPi5rhoI/1jXcs9CkxyVZyfiVO45uck
iW0mwzuLI+lXEd2RcJpljQifim2iao1q5P88PR6lWLDQfBO6cK5oDo1XkY5gZgg3
DEKf2aCUxJUMrzjzop+7dfHXcK5kd/799HwwLwDlZ5kI56WmWb9VlIddDrGj9M4E
gr82HIfLGmDxeFq6sCj+DkYlTk4dvatfhV1L3gZl9SnK+qKpKTrAkUQ5/nOze9bn
oFwVd4Kdmhn5c6DCs3Hw7kJAvIA3/IPjc4vgHXyd209vqW3yx3ENrGxsu74E9dMq
WqRIk23x0t+UxILjcn7oFe6c/UgUp7O7iJO7ROqhVclNLy4xIeqTvmNOGJkAeKPA
eLvHMwe7i+7odiKyfL4zpk1G3GcibfqSeLkOhBMW8QaiefG5Ha0u9/xYiWF0Wikn
xJsagQ2YjiXgbm7S212S7dnG/0COsuaJcI207HGM8YCuOV3PYCmn8j6nxEKC2vO0
9n7xkXkJd7vD7zHuHjGEPIngNZWJCwx95myaNp8wXP/jPJnDyqO63M3Q+PSYmaG4
beWC9jRJr0DlQCnrwM40AxSDIMEs2FQoBPyLO2aa4q8FmScEcSIaDt3ENLAQHdFG
IBIHpVZSLkAFpCOyufOaNfs1yhHRFzPjmzoJHhWzouJsh7c+L7QbTbaz33UYiMU4
5pmeEFHURlToGWcPRbuTMPzENHbjYZzbEtdDKXDhuiAgjPqLxBxOqLOBg42qc4jd
CMvMkVk4Yp9okMHAc0p4R1ng7xWXFMJ5OzBh08jkx1CSH3CmDZlMnVyX+wed9ROH
CuzXKilVTp4dsXBdZ2TtcQBJH1YXS7gk9YHpbtuyZgFal/Hg8h39aeHwW9MYfsbI
uvqop93KKUFr6fFyi8ajwHyDnlaxezLUUXqnfGWqihekE/If7dEpyiJCZKTVMPYr
XBlfuo5JxC05VZrW2LB83mfqKJdzcQn3VDnrwVwidnnqy3e/YyzA8fCLXLziP3EK
9V3R2mzQxZ9fYHnWX/UBcC+7U+zsAasMmRmy/SerL+tkHlUvB09oEAt14M7McHXn
OrBTvnihw0cIVwNGGS07aHtk8squW2JKK8gOS9FSSmPk8/kwjxDEkOk6wh9bWNEo
fIoEJmQjZZRv3+sYdzdvMkrW9OD2JJdTHXGGYlU2L7DcftjvsIXDhUGyJJEJhxii
vxQ9UaRHRt1dcLMFOL1CqV8RQ7txFjMPWXySOiru/EcFjkFdYWTSXT3k39anGZwG
tFp7D2eFzo1upGyi2s4inRBsBGMv5lNo859EdrhRdtSqGk9QCc0i120av+yp8NiQ
KX0wbyeAWcwMpzjpi+RW9a5lcMTSQiNO2NZEatP4MuonyJ0WrxJxQVnu1STXvJfP
hcDqWk5llAql3YtBuc6vATiLxG+lUURlbzUpki2nJRbZW9ymEoJ59USuAA/Kw8Bm
6wL6c+gIRRF6k9R0lFqz1yDP6xtlr0M7IhUrHvkhLFeBP1iXsbpg4j/LmYo6+F4w
5K3G4DtzRgquWhZ4/Br15yVdTnxPcIVXFNKfuxR0xvtP+bcOT+5yiO/rdUSTr+hz
vmaXPw4hpqTkd5zPF/k72ffqVhZ2nj1ttW0IhVhDxSA8bIRY8ueceG2HH7G7jeQ5
R3uehLnkoY+BSvTwJSCpgymqSKa0dWFAjwJmrFQOhsh+htlzNtf5EtbxWFdEsa8x
I5TYgiWQaMqGpef7x2xZGHkKuZAUY8p3uWrpX5Ah+7hlIemlNcti6WAcMYuSU9px
LQ6MO8/yE7QKIr3pR1FTJ9dcfsknIX3UQAcivUxR/ioLA3JV0ZM67qT6Q676iATF
bh/6OQZG7T+jGb6A5ILbJ+b4SFyH6nzKYTuFmxM2LMHnr5exTMHoC30mUAc1QQib
emBbaNGaWX4nghGoRdCeQCPRJihsjh1p7gN1R1fQ4S/zV5ViOta2t/WUycWIljHl
qwh8ndhJtlC/bkLcDcVQOpvTb2/KDAt+YfPy3J9Qp6tgyBMTyUico/uk1RDnYb54
cFX3YNan5XIZ7YyoZ3+cORL/stTTN8EK52gaPurJlGzK5UaZhDWPWwpB2CiD3Obl
lBGpiTqsiQwaTSquZctM1ZMMfkwiu+Z/CpaOWT2KaDZbJ67kMc8/qmKxBv/pgGZz
O1JdFnFqGt4H0ZgYIbkFrP2k0ViyeNGZXRF5QPkiuoqicFOr+hVvTnrNt8sMnlpz
oYNW516ZLJPMpnH084cSLQpLj/0mPTvbIUpO6wsX77RXifPdU8y+xA4Hl0FYhj7p
EmpAgdwbnwJfKA/sqh5l/0s7ZTrZqiPQ/92+DnJaMmO38GEyiLfPApGhLRDjYRaF
PzN4hsvTTe2R3xD29IjQmykzvO8vCmAVnJkrlr5YIbdQcUNWY3hMYKSw73kkZ30D
IkyFoJlKe9uN8TQFpYCIHiGOu6sFm5hgEOGpiqoqTcycaZyfpwEC/TWgc5o43zDr
Ax8GWjacNYq9ZEfBgaQlIxbQWhcoPHt9vLZigmcUirjBTWMLWSSSaxrk8GlBcTxv
jJeeR3xs3x8gq2JoqVYUrs72EN0BXBtU68cn8Hrpjk7qnipDK/xs4O75tdlsMOaM
ich5awvxYAsD4m3spkIj/g4gQRyax/54YeDCbAgt097q7Wv9TlNP4GGeYNBblKNM
Jwb0HThAltI/nZk/EgAzT3gyV17OUaKGpq0iB71DsfRoz+2doUxcUl5yLQylAb3S
NsMYB0y5KKMg9L0dEcsjzmNQbaLxm5XZgjsQehjh4hvV5ukQqIxW2gzQdh2pwEfK
8+4Z7WtUz2EOdnpZPggoVGkc5BkigFoRxHbrPzOYEwu0RICWnqh8i0qBANd1dDyb
Dio3oRs0brp8mUm4JcO+bN2ALGHL3MHw3IM5AEyDE9nepYikH2YOqBzRacLJgmd3
l5V4DTCDGEgKfcy9M6RWtZc3U8QF7FMJiHYqNh6kRcGqvK1w1pGDmPuawA4h1ZMH
XhUIIiC5JjXS6i5M9u1BsX8PVazLm0iiKT+s8xZrECSNaQipMd8y6D2JnqWWVA+U
RLbbHBtfhH9msynX+JuFteH8xiD03ofzj7T0Ir7albi/AH0NuRezZDUa0OF5148V
4XBcQ1faJ4KRM4bzvaPfAa0RJB6qmttG3Ddd8pAQjj2Lkp+OCbG6hzDrysXPTkx7
S+6wpx7p/fYgTsUWrlwuI2pQveE6WSYuksqLs76+N/jHjYzPfklP+DTXd/r4Y3OK
vjdA3TSDYmuA7hprLfSST3mnNqzJHAZXWdS2yr9K34ntIj1nfKYqOCUJ+npTB+cn
YIaij+rVkFR88ISoZQhoQ2Af4tGwGKovY/6wmNacT1MNcsuoi6Tdgao7ESU5R2Ys
DMBZ7wMNV+s5WarezR+tztivYbM0AgYAAyiQuSzJ2O2NjSEL9Oi18FiveHcXx2wr
dzuMEBZeDFAyW4E2rv9aINGibMTjGCFihDMh4SBrLSxrBVb0u9HKK6thDVaX/H8h
En9xWoIRqJcfHLywmUyN7kK3Ne5mpSy2HKOBp8FDMUAtxroZsA7g/FYjQookvb0K
0NZnY85wHu+ZN+G63g9dmA/FfGrgAOp4zyaPkRbeuXyNek25m2o9eNCOcx/WNkdg
oIf3ULHtXkrWp6Qxau+7O0cewAqsPOp6aXG4l/xRzUH/ztdzn2RKS1NUsiLeX1cU
f7Dh/qzeemH5p1NdS8LkztKXyjssu0MornGijjoFc0iUmLIfgHBi2w9qqyxy9ssO
fHZFrIUgPivsdvuHCrhvZ33Im9Ub4/v1UMxHjvlITZPu0MaRDSda5uaGVsnAlbx+
FXYWRXTyWX1KPr+XnIjlkHVcd8XiBKHAbeG5nPJV3DI+4Q3WmVa1JTJzextjSi1S
rKpASjBz/WwLu27eExIeB/GHwndwnOa+o6xqWcQ6xhRBi5bmTf1weeg2ihNzADH+
allBZkcFDtVceAFTNwrE7LJ9724GfkOTdKFFoeYVfkbP29/9swLL1AbuNAdS0veS
ucHqJ7yPGjiM3GUDxj+gOBdVzc0fJgR0A5sSBlMcJdUbdfZSs41OA8RCzyR8Sw60
D3P6SPJCxwoaddLuWyUh9ANAqIG1Znt9RU+BHvPvpSqoyJ/KxgQRKe6AOwM99uao
1lIBDFnvuCFtbU+LVH/DTNKtYWPhpNt2VK+4sBotxl/mOl01QKBKPZe9rH6X9hKN
2wlKh51UIXuKYXpHYTl5huylxzKpzbG5g2G/RzHXaSpBTWQdAmcjwxzPfB0KKaJg
bP7Vq3cMAPi5VuM7iFGcL1rl37rAtFMTjwwILOMsaFl4HR82wUA18UgssXFqUFwO
ugHlQG2lF9fyG+DQdar3VWqNyyOdfwOL3H9XCsLRpu72zv7zjO108xKjSbE3siWx
UpxUTc2vj3StHHYpprhjybaTQyuHWX0Q6akGu+hqXuHqBqttZd338iMA6rH76svE
qoPr8nt0kQZ5xf96CB0FTxHhkrwvgjlMnWAb9uW2M/ZBbLS2LGZpk7i53Xf4bw4m
JL3Wd8knKEMq5WZICJ4JCxQ/BtAvrDbi1fSkQVGvnfDrANUzQ1vsP7HpaL24mXl7
FGCb3+rRZyMLFBixkqdplZWP3HrjCZJJquErEBckZRqF5c4o0lJog3KVOBYhbSqN
Dk0kLdvXzGoXUJotlkWAkmAW+BikFvwvVdxk69cmBeWYJJjnbRZGyLAyB/TKv4Nt
NchoaF0FD+0DIElwOLJ+9xM0DDuszvAqEUEcMgsHpDHS09CE+mInT/PVawkamzF8
pCcvxWJzlojshGU3TMqKJdEWAJmsuzIMcHSFC1wwt7lo3lRrcMw7bewjAkXaly/H
VEEm568+9kcfzDpODVM6bkloX1AUrFMqTRGYZ3glqcidKDcPynaB65DuJ9iAzzkw
pfiNkQf0j+xEkzmr/FZK5z4CekFRNe6q7ZufQ2oDBpzZY9SaHt19rH13X2+GYoa1
9R0rlGt5mBCjb9AmmaH6HODK+nx1mqJosCh/UJPrJVeQi4vkEmqZEqnQ2NJteAXC
5buRb4EWSyFDLmq/cuFiAoZisXJ03yd8xBat7WtkwXhwHgGDMLj9bnKnzO0/wKNu
A9UfQcCrP3HMwVvfPsoxTAJLNOUGZOtyJcoFFUUCi30OJQgOAg/oLS9kHbcUmgUj
sdWycqUGDyEIMUYocgObT7tNvZ9782HRsuRFmn4IOc5flq1OPevjgjbhrRdE6H5d
C2WIfpH9/TzoEMhtfNeqY/A/w3O56yaR8okZ6Brhi2h/pxCOsel5RbRCU26UyMoF
EzSLq/KfAF8NF8lFZR4dhVmkP0FJYcJtLmNGRGs/IV7QTonJo2ed9At4/CyuN1JG
tiAcvRKvLgOJ7BxDjgN0OvcYAkDywD5eSTR72COZnZO0b3COKFu6SXKw4BnHPwZs
NI7hJMZ3JonQsAJ+8sRAbYI2BtKKovRmnk/Lkhv4ivdhDAELsk975W4DoxXz9FUI
04eCdks641IR6GKKL2RywrLN2VRHqhMERrPJqZMs6umAf5F8EWQJAab1ZE1dkk4R
IU4c6E4QrcyL11Lfe+ngi7O7u67VBaHC0koD/CxpPtnphZwjXnU6qla59fppBu9G
NknGKEON0AZIfEy/b10v8ot+Vk7TU+1YZa3wLKqdss91iLOdXrsNzbJ3I5g8wTi7
qWEY5QR565HyNjZiL73hBJH6/b7mnlFuVEdq/84bmunoxX1LDAdWA6SuYTJtXXfT
nBdnNOVFwAElspi4Kjuc9olNq1B5jwOtxb8JVXAOPRzmPiTXRKsOgGsLdRo0+g9D
gqLNCch/UlW5/tTHHpm533FD3r32xY+j39wEzWFlJ2oVuByK+cr5eLPSE+zw365k
XUz+xR+PpiOjTylLzwud1JNe31aBCcRMiabVYyDdxHV+/tq2Zov6qYA3lyqVxf3v
hnCx47GZcSJmdp6Lst7ykFTRFZxqu7yiNIPLt7A6G+faqCKgfiDiSp7TFpLxvMFc
PyZWwUolSChsASDqQU9rP1vFpxenq9a8yjbRUi7XQssVq7WXcqaOaNfIL6yIjZ+H
/9sNlpaeJSJsL3EhFZJha17nc9MPyono5aUe5QYa+LouFzdcQDPuHlEdWXW8mRCV
N17hxDlcRD1Yy98wlEbLUXItkCRXN8LZmz2POk+YK/WaGAI/LI/e3rPvI5zb9yth
rbcKbRCkK4QZwdqA7R75e/Pk+BrbrHMlXBtsqcURj92s/pNmvQyqvCg40IdzydSa
h8WQYL51xB0lKkgA0GfNIIwMD/Oe/D59MHntlpuHDKs14gi6gq5bRbQm0FtdezlR
5DL5EylNI1rOVFxr2aqdoMdGA63FP4E5emKJAD2bd0KxU5aqUGb4uKWdW1Vg/YD1
77xLlJbPsxqh/Uf4/PLMo4hWVgC8+fAk61cszgsLe9cLwzdrvr78OJgmtpF0PzKK
2gU3RkpupBMOKyib9WJXO2aiJK4124ujZ4/+T8z6aaWRHMfNWJ7ob/4GjdWsQxfT
jZ4WXBph+mAi0DGhW7PTqRDPe99Q83G/YyuT9RmgdOgsN85KyJfWnGJll+ioRRep
D1g0psSfTgG8w5091wwCI/eKnZdNkRpIGp6Nut1z/bRT54HJbgzxXV6VXHZG9+mZ
n8+8mimfqyvfZERElMCu7Xn2kycD6F2xLATeOGyViNDsVJ6NUcooX1qt6X/g9gNb
l/kMZH/x33XkrrUXj7sHADVf0lrGvr1DwD40d1ezCWLNtoi3hG15Zo0FX5xKaC9j
OKWgmkOohzDtc+MIM1AsshTuj27Cd6rcrIvOym4PzYn154rmJJkVHg4xY/ZYxlDc
2PWFxnmNtG8COiLKMFZyLYD/hm/+P9nNdMJADLL6XulmoSw7JtLWG+8FuBg/Sk10
C5NUI3TO4wp2cnryxQ+Be3jtFivJEfPCK4+buxu0++Btwt/2qvoM9Nq1pHZJL34/
/q99TVbFIRdZIFfmMHq6pjW5vUlRw4zRKFTBTancRTUiCX1/UC1c2LDaCBO6OD0p
ZryuJRbqHPtwNXFAe8ru8LW168mq5naIt6HpsTISB6/RfOjf+28nhvGKSALUCRQs
lTUcqmxuCv7bOt5Nn/yeRsQU7l0762K4O5Q+utqTjnNWiBFZxUM6MHEJdQboFmxo
LCpgWf+QxSa6N8FN6hkSwmI6iujr+T7mbRiTX0fA4V7mfCZDbZgWQUnFSicXBQIl
KpdvTCSBuQHAz4myVjp3VigLIfLXgyyVouKthjgnWtGfW5hvRKcq49PkBSEoDqlG
Ip1+c7Ds858YYRtRRgJE1y0MYoocaGnqfTmYJDMn62qXusXnG6VMK7aIpIgMnEyg
S/l1ZLpLwXgXQgBHTdWsqtUUJ/+40qUh4QxpIGWyaROhFhZWqCRDypffzMR/Swqz
pzCG0QKHiPDjQeuemkjz8leqYa6aCmVQsA8YOQ7jPbP3gch4Ev9cKxc6fVCW1j49
vq8hsaCwYwlPqv7fQH4QRZb52BwIDWooGEDOnr4T/ly7JWrT6iJIlyrWWjCijyZ1
jc1qm3/1ehskRMD4KuHfF2onxD7V7kU4HyN00xNEEGZVky9xfrZkacpNkstg+v04
ADjVhTZ8ta9tFkXuU0AsBsLLS7WqHn+aExgFbnIkd8I7+uqhlx0757EB7q1BwlHs
CQHAcMg0QnJyEY7K4Iu9am2dlYADCspADuirKHaPgxDAkiRppw062Ik+a5JHWFD6
e4OJBdVeiqxvedG5811vHVcYVjFa2zlkuP3wWACVbh0oDwkh4Kd3jQA2k/oWmC70
SJiyPKZewY3A3JrZHmyB/AmtiQnieK8KpJ+Ec4ciof55XZWJU9JnyRljD7LQV3s/
dL3ZRZIJpkIpz1Uxobe8/yoUTGxj4hoLRwN640Hrdf5pbgpwNbu7wjIK3qL3UjoP
jgEJ3zhf9P/AuE3zuB2rzJZq8QO40eXBQRLA5hrLJHekkwZ9fDjaiv4Emx/UntRT
TQ9WFn/CLi9jA0tlszDmnXD/mT0qnhp1y+aBs9k0Z21W3Cu5Cploxq4dQ1vqY6FV
FWp00lBPpfc5/ft0w5asFLX4pIxmBOGaIiv0hutfWH0FUvnawGEYEDYX9wP514Lx
/l66T0YjwQlirvkE4tJFwOssbZxxiKkNJwBcefXFRmK3p182wPKkQcQPWtwNACFt
/nOupYF33IXKWzei15k7r5CcjXBgpXycI+2VcThi5hvBNI2NBaZW86DIALNHdhI0
PKrv21oSqcJbtjcLSjpmm9Pk8jTtI5qQfUuqrCLj+R6YYR7BADenC2WKzpSNUgTU
UnRQV+1Z2WPriFnr60wUYy2PjNT4AXKC07nsha+DdrYHPbGfum30Xi+DOecufN0e
IyJ4XvIz5BMWL4UcRKJecX+974+zA2c9UGsAOpWjb5FwT/nfeOTZmrGP1mlycMAv
U56XjXD3eFMPgI7L3cC0Du6FUKMZAVNgK0qI/OFpwtU4WASz9yKp1u7CIHnXYxuY
+sa+JqSevXPZHl9+kdfC/HTf7L9LbtEZJFdzu2ZfIMQek8RlesmZQXblRz9cEVwa
xuqXc4Uney6uPANK56tbqADxyHjDrSi1J5zM5cOz3Ox/n9eUHWfez8Y8vDZCsgdJ
6xfZx3MdJ+QRimtgfIjBY3ORuihvK18o5mRkScLjPUd/1geL4PDI+0wGw5O+NQHu
nv3rqEfyFr48epFL+o7FLcZDrsvl/r8S+nqQwyOKciK8Mv+TAWSsBX5IFciKL1Nk
clDx/VoAZ01ORBM2NV8LUT8UhGXj0UC6lw4v5uH3i5wmSx8bEVbZxtKH02nX+sCT
IrZfNZSZ5aP1OT58kN9qsL7xz/LuSQ7ENpAYKcUdGJMeZ6/ImrYFKXcHyHo0c5ey
ok3js9c8CptVSKiOsEwuzs3K1UEwgAeP5MrJd3CborohoEKxVaNBznq3VuK0fiNH
klUez/VkBj+RI6Aclsa9tuuXaTnEfnttXMgbIs+4S+r0myUPJId8sFW5KHeN8bmc
8fYvfmsVfMkNRfXV2U33+r07oT+xkLK/gADUq2YvwgpgMILd2hkIYVp5unKJaXRZ
cxp3NP3OXK2CZnmhkodcHrdAbkiLR3sExwYFUSdoSAwVAfHM76ep7JEaIzjsgHfJ
NuBQJfwQGW6DY4OiqrD8yXV+QCmrYJcqDlNBul2pbNF4VKQ5KtH6+bRAglAnIxq+
INIY4pWfnoOWtU5H0tcWzBB/rbORTCRynw4F7t7UPhHDNEPbUoH1uBHiLg5NOr1Q
i6DtyaH3oUd0VK/0qMqmL/QaUs6BmmCub5sd+gn33/9hQa6GhQmcm1XXzs6yGg5R
cNR8qSfUwDDCKiYvKL75Tt0oPD/sGmQVzO9GhPEvCy4HbKL5fZetdNltyxbO4Xua
RFQDXq+mCD6nc9XOQ07snTHqa6h7pF/zV1/YSDWozsw/CGUXgDI3g3AjQdtbYqNO
qA25kUZYYe+mocd38+LVBB7nhpaubpRhGEkVUTwHDbQpD46TmmJQtUm2QzCfxqoo
Ic28CFOxVvxdydw/CK1l29bC8ipg/8WaHDRraBisE4XR0K2KHEZ5jPADJ6OtVaTX
e1SKDc89xkJJhBeXUt8NyP3Uw9hO050gmoKVhRItIjuWm2iLV5iX/you22LtjtPs
ea4cwgYHHKPCZJXnWMcrUBXvqZinmm6pc9NBg3nYF2eSePzAqmZ2VV4U9Y+HhGfU
KdxH+m+4Mj4/uWkvcE7Ic0I2yGF5BzHAjVXvMtWYU3E6qiRipDL2/oJ5aWuZhlbZ
dqkjidoWZVqijvs9YEH0FoqyqjWF22mf9Glrsx/nz7oCJHjTDVd4Tn3hLady9TAf
QykaMEJP4VZePajokykUiiFLqyW+UdDEtxsrPqss6ruWZV8MShzU/Jlpi7TRnz8C
U1IWZWc0AsfnejcNWR0Ttdrs4sXBmNOuO7z+BMzm0LHdy9WjAGabUUJUVAYM5Ss/
EUpfdFG6Wy5K/0P0WDvpKh3dmMpdQRR3az5zdjCsTYlXkcEA1o7I8NWQxFzy+k/H
FBEfflY5iK6r7B8psN9lv1K6LXiL9naYF2G0UgA97G8cRje3lKhUl570j5Z2pruX
Bk2OD5HN+x92x4BRJgsJpkt9N+bretQ46S2BIqygXdozwZWdueqeeVLDwD0mCz2y
WqzwjICyRW6wlj+grPtF/rea9nkOTN+u/jr8Df0CPFQQla/ez5h/mwfTVc/teCJf
U+nqgDTi/ICoHFFaCDLvRqj+IAoJOhCa/gmvWawp9hZvIz025UQsF75LXpW04Hap
Yjfabwiaxqi5BsM/XTf7mXv0Pm4JGN0v+YGrJ1iBATYWR5SLLpBWOfxzkNd6wVKL
sTWFLBFppKAqJISBzyxGn8B6CMSCihAPFLvHooln0cTMDhRPb+/TOF7AKNAN1Zvg
k8unEctvGrFHzaud4/5mDFkWXGpf9c8hA4c43RTKu05aJOS2iTYPAOFIGLfOMqwW
3yHIbbew6e2YpqRq0P47Fqmqk8OtPw5XEJ3ZN0t8KG3/T3NbPnGrHACHxbYc8ZAh
Gsc9koP0oeVxcF4qe8S0t4OkSkeL1PZIpxrDXm6nKPSqvl3R3MJ71gRFQao3LsHC
TuCNJJbEJ3HbIZ+AfPNpmlOLaJqGLER+xYk6y2B7JrRJT/L/lbutJhpW8RuS8XSU
jVWBZpb4xgn3HWj+dD7bhSkn+5AvlWKMnBIyLoToLa2eKLB8rvKYWH0+Wv4SQ95p
3Jp6D/3ha7BPXteeV5mWGf9pT/uV9Z1ZJ06y8bSua0MGyl43tI4T7hPi5oIASuvb
enLhJDX/ZXnzmQ4rGCIVBrEyv/jrc3AhD4ffAJH8QTI5cSkyqD4k/BVQ/u4nshl0
mYNOlWMb+G0IqtofmCe9nY4Saw6cFpqXEmaLhHCyTHxrxPuVq2xO7q9fGQPbPIYE
GSit3qajqi5xXE1339X2EPsxgCMiYv8g4nOz1QGBHZihQgooIfoLfSSqCX+RP8Jq
fo9AOzFbSEY8uWgxTXhQN29++3iSbcnU1YF8Aa0IMEDrrSscZLexAW/ZgVgx1x0i
quetqRBJ5XH1pixtFwAV+w0mOLH73VPjwJ6QTzZB2i4gcgWJ+yMmxSNBHEcUru4N
PwK8BAKqia8JbYx8Kg97OsEUJZZICJCFu3yXTX/tTRu68QiHbhGOZ2Mc+nbSC9TL
+Y69GujzsysnpoW2fWVNLzVSYHB/jADU5S+g/OYAAdlFFlY0zngdq8QFHz6kdEM7
HPQs0JedIZpEwigH22/AtpB0Ubc266TDZryNxp3kXbSqzS1hHbbMkjzcNPoV3+WR
SHCJRYathDUSTfzg8CZN9y+Fq006xKOHe/c6pp+RepKLrwS18hko0AXCj21WuNgz
65+FBiMGAPCIEJTUDFzRoXTpW6hBm9AZaFmGJMtKxeI9BVxHHT12nIhW0nAlOnkm
YgO24qn7TGOWb4Dzi7uiUbPcmaxr9oSkJ6iRBNazvqWILoC5hq1rLOzNmaLGhFMs
m7YcJuEiFZxob19RJWm4+aMJsWaRrrjxkdygQxxOxFKhSYKN0SOoLe9rBoKLA+ck
D4LMnokuPfsTiRHe1yv4UqGljpH/csSCVstL0RiemxTARL9XvcmJSJyHL/SmhFry
xC/SbCknOM4DPeiYfqPq4VPHPG3n/NBx5BSJdr6DN3+LNlluAiFSad+Fxvx6+Acr
ATnEBQu4BuQEWqMzPHY3FM5XMDXHqTgoq7G3eCVABdTftY5ZsvJytq72eNCcvfeB
wY7Ai5l6BxcDjLITMbvenGGpOFI0fn4Bx1ovvXCs7qK9O3Jbt7PE+LM+QWYQ2ZPJ
wAOyppi7TOxX7ZTgNXkJcFief/CysJBu44vuvwo9U56z2XiYRAcKLCYoCZtoNUJv
DRjwcOVlXnfvIJYerEXOw8r+zBhuHfenfb6AD+g4sELG9aj0BzC+02C8ViYyjBlY
pENaghMV0upESgGHnUtx2kspcEpVYTe7YyC83jkVjqClg4n3dGG/RsLVbCGXXTLO
FfTzw87flxxdHdLYdIks6YGeF+TrYwmy6SJwRHZhJ6Blsjj10fmnCFT30scgbIiu
Nte5ZV0mQmD2RpmvNI9Ii6UN8T7+CjSqdkqpQEQc8bd+zSD+SsGr5NOsrEoBaaFP
AKCsaHMR3eT5VJF13qBr55e8c4CtQ+aeRdljWsRX8LG7mHMVzLxdzLOMdgqOE9Fz
0oon7LDmIxfBJDbXCykyau4acFRicxrC9VebsYUx3fbHQ1wPgIdDuF2TiFUFeMq2
YcHSBe75I3v33N8l0ssFWOvR/heiGIdiaw5yaX3vSUbulS+eHi0UGQ+JLySyjTJF
Br6BYxQcto9/rBHUj+MF/4YdvFBtwgVyQxMjT6wp/wl1fQFka3AK4bc/pGNH+dzn
qKNRm0azIMF7Le4kNhWgonlghKNHnBjm5yfgz9H7MGbR3+P8/5Adrlr6lzD3dm6+
qmeiZ1Rs9sjWJp40qdBq6TLPPAHtUbiPaA2mF4aT/xLaOv6m1jF+7MBFCEio9lYx
Xk8eYvw50kI/Nbezfqvcg/go8icrOeo7pVWNE5lWvpstbTeUZkdGSwkuJfAl2ug3
+cnPlUjDGg1N9LSDja0urWcCMYGjyB2tS0DEAb1gbEgB2mbCq8k2ClH97iTAIfX6
5OFdNLpD3KerfLdihzMeqFY232ritDzpNZ7RA4DJhzr1Kg/TnxAoOOqd2wyMOAyU
X6hb8yH0OoQLMYcaHeCGpUL7VwcTZGegcuoONEch7h/v+4fCBBNVeoMUewc3VB6a
lhKDDhzBEID8Y9uZiW6Mp+TfPGOWPqIpFNEwaMgOhK3jn4yL2qZsnx7DHv1tM5Ls
raWGbUfdTMmZPTW0858AnISOtyn/aYxKWu8mfZTWSzgnd+hQfszRZvEMVjUsR/Hg
kKBDHROxwMlamTufNq7ia3vhkhwgoFR63sLaPcq5MDxMaYUBwQc7+JTFa6JRtv1O
rAZEwZkzWpVfCfB06KEfbbsBVlSHJ4S89KAgnBwsWA0uPt2eYLhrLzZApvYK+6DL
0nSjSnT8941CD4IG5KtfkF+3rWLmFW3XQFjaHOlsh7LzE7uVAxEOWE8nvTPerVpQ
iK3wUHuNxXETQgei7GJFJCT0l2hMX7qs9iNfFMFShgGdVTV7dOzyrkTeH8q5OKaY
CRvI9dsO6ciX/YGoVjw1M8cCjJ2Bp8lqwko082DE0vSA0woFbulTFUGNYzSbtbQ+
06AJtfVmppmmymOKkBTzgw19SgU06T9mM92m9RE+KC4CcsPPqj/NuD9gQ4dLEzdB
kU65v7KWCSvjxoFUYaJLwiUDtjcPFDhnOcZkGa1Q8aF3ustxA4h706dXRyyBIYjB
o7Hqa6uE528ES+HRk218K7dKcPDoUKak2+cpzFPs8YNOIkdtz32vWROPgnzdPVOw
TXMal5hBEtUiG0LwB0QHFoDdDqBgMBAbslpq5nJ0+B6u3qq75BpUFSjUppYMp7WN
6yxVn8Fgt89QeAeIlYt3Oa9EXQKtu0kNTnmGgi9v3W0ujAlLAMQItT60pY7JqeMY
aJ2YboafKjFsnIfPk5Zw4Sj/GP5pohQ9hdK5PYRCth1sFrMNRfwgjHH4q7oUHsks
sdZQoLhVU9lKG/+9o+uI6c8jNsKIKFx7yPOzxt0fxy2U3kWqTsSCqcIJe5jLTCoi
illsKPbV7jw1606Elq5c7DC497UMdfeIqMClefK0WwBwyEQCO6JnIyO5FsspHDmd
RwFXWkan76ITvdMrP3mxQ5tserZJCKkGv404/tVvgSS6frpXQ0sbeY6r+vwklgd6
ssbMMKMo/RCPhTSPpieBiBB7yzkpdg3qq88l1u8rQL2Nc2MwDr0X/owLy9TllHfn
qwRSsydBlVanSEnf3hZ+2bRL3b8btzy8TPXrVxBuY8sE085AcqsxYh1ZEbUej6tQ
cUHXnAJ7Hq3yU8/MBG4qBRJH/xsPXnRwpQRDC6R+fM8jDKCp6jUx9HmNWIA/aVlV
h4BbCwfD/iREUx4X+KA9r3udt4k2mm+DA+BFAHvelNIE9gHyDG0zqFnVe/VqpwCm
geNHcWRi0ioUvnjo7wl0esm9C/Xjik7p1A1rVUUfQgcqsb1vwHkK++WXJIm1SDnH
KWhgHoXKHObAZ6KdoshlF3o8ZKGDiMtiUpnhagAvy3aQaG5nT/d3MYeXH+ro2njk
40gyrNHOz8glFdNgCQPSSBMIdP3fKgVDW39WHmwCtTHj9RBRJEcoOwNSUJvVLO21
PzigNn6ZfX7xKO5QMtzMUp8lLmZjG1VS9s1KQg93YHfmwUCCyLbaTopKT+dTJP0e
DneysqeVoglmSY75gqt9Lg955CYlCfZ3Vfeu4x4FQ6TqhhEH77eIPaE1U7qbtfdl
qZXO7AqP3Am7hvjkGZinriAu8Pskzof5wDPQ8fRIZXKcMwTy+qdTMfMpgU872//q
VQhDLavAIeg+x0Iyj8ig5oAQDLcjOF/PIxCGbx0asJYKoa0FrlqX5wOdcabcFbeA
uTJCej7P8iSlMyEC/fin6a5uQ61Ja5m6E/1xqRO2RARHpsCqCuCkg/EvoknhQ2Z2
GcXRRQGN0lyU+FAAU1AQkp2F8INeehIcW9XylXo1uqEIbjL03da9sy6HdVxHNzeo
ZIxDVmAl1HJ+uUZ+PIGRQ6aw0ojmt2cs5Dczx15fRxVr2r3F2UUQjajbj9Vl/B0W
TX8ItQGspgBasw4UgdpIF3txlFbs4xLASZqAoV6OmuUFCagCvUT4cEsLDEiH13Jv
kb/AIUc1uJ4KbrTmLDO7klLwTjM81E+ZEL0fxFLhbTLtIqQ0umt/UFWV31YCLXVH
02qkby0LSOmu1xLexztSaNVUMIsRj52KAzpk797PeOZP+aM3aHyh4qB1UOFkSNAh
Q3sC4sX5ZyPsHsskGoDkoara6EITOTkJpTsoZipWOQ5Nw+ekZ7Exrpv8yk8COeWW
J3RN2RQoqqdvsxjcessyrSZMPW8vvVJMZg0KdG/lrSvggnzqBAPOLkvj3DU9L61g
3jWntQspU3EzGkih/eIbZgaC25D0tlcQijkWLotXqJw3NXWhZcoyXmZQBBPlOULJ
z2IFNQxS0AqZS8RCI+gbfzlbEY4uDfCik/4Nb1xuWPVRofLrDJf0jnQqUXbLAiCm
wG2aK8Emm55rZcMtR6fThsDS1krPHyrk/8ZgAgvzjdlG4TD4qyy0b7EXp9/QZCX/
L7ynA1kIA4R1ukItVhhdy9dLr5RjGAF06i4sfBKzjDuRW/paPz0nJ0rzzmtoaJII
uD7sYjYF1WbnuJX54RKo/T4WWXlg9zXqXdW3rELYsmT6T9CsLVBU0STwyxRuijl9
1OvSeaP3hJvb3VnXQztaCjtC+i0GEx3js9GLaiaWe8JRsHRQrKxMaVN8O2RvpUl6
suSTZY33akqjz7ef9Twxt0s5qb6MCspEIoFZKrkTiHvUHaXt8K4al1YaPWctwT+0
PiI5gEj25XP4zAjqG24snz3oAXep8xKWUtrVWQOG7YhINQZpw1h/VZc0cAGI/YOB
LUkIMRnWLuLm40Sad02YyiK+pR2ab/VYuoAbez27xsVoiaduXCFVTlmykz1zp5XZ
wP/iwy05XOolsOtulmn6+B86jVLcSJKBxfJA/BIDV8s+aGnaGZU4fxK6uyK9BeWo
Rpi2FLRYNplbx/80SXURzoa0vrZULcFLyb8RBF1LY5b7UbZ2ftIAgSClKV62j/Dp
KyqR8w3eel+YkBhWc3q01QyWCAVc4fO7K+PFi3TiUJcCkOUm83nZntkB9qsWsTdz
DIVwSkYyzMAc/TXrv4NpDvQkpIbJD+0eLdyyzPdaB8s+FFfSo6iM2ARHNlg2P9y0
lKMb7lkJ91WTrRcN97gnWy2LxYSWEkhkdGa9rUVW9NEqcU7c1NSx2F3DBJzm1tMV
67iEPmWcVo7rTrkTVHDYvK/j7j7Rb3eaz+MczjGC2uAYeyJ+PHZmCrVop9bCdwlP
LDGyTXeGiG9MREZiztCnxsc0GW5INN8KwIJOODcCZQik/d+ch2CroIZ/pOcpf6IM
S6peQdESCocwoWmtyyavbjuDH8Bg3Sblvy3MRxPERcymzEY3f0Y0HNBpcuok+3Sv
vzgWIN1y80urr5tjK5WAJRXnWpkb3kMC7cecj/dqawFZzF1Y9QTeSpsNS2qQst04
E9Xo38hm6Czi4/SPYZq1YPSu/q7/JXvoIUfr5zu4HZGuzCYmsHkV7uq6IXlFAlh9
ZvSVNEj9klduKEqxO2LygIs2Sy0mJyLUiIsFvj1m0dv9s4v32IOQq5rh4JPrKxb5
Reai7+fNR/QRqmZLbknLY9f6+BZ4M0ORjRZTiHZ1wa29pk3SjX+1jdA+/3LXYUv2
qCwZVDfjPhXfCTwuH3remoBVPqcdPDWKcy2wRgiVoa0Tha63icXdhN5dWRgnv1OS
UL/UZMWRLO3Vlj26UwsNseTljPFJDCVOyjvvlmR8nLnSUssk40JdLWbg5HIruT2R
f0JuvB3SUEoEaA+bVrncjq8mP0hYa1T4nsDH4rIhWRC3piNPt4I1U0kdkoOiTKRC
zcXuPM4d0ZWsMEZSF0xbhud9bLEFiMR4W/p7CInQrDtVn7+e7aObvjZRfMYw+0Y+
X0fHFTQqm3GjDngwJZ7LWo0sN0ohn1Epxh4wEZI2/7TdxZ6KKmp/W8zRQAHm6E8X
3F+FivAH0NO648vkrPt2o4p5ZbnqUtIZNRFz/Y30OiBhojeCWiK51xlzMnpJxQ+U
ux7W1ZlcEHlM69oqPTNG2QsR9uLg6wOMkAhBL41Ce8jS/qwouaGzCkJD1WeFJ/LM
1YvkPmTWFLFHsFUqj4d36TlubraPuMi9y3sEppaX5Ss71sjC+Vb2gI53OC2W40/8
mjomt2CH1v/oz7IkyUg6QR87a+Rat+tkSl/80znGPcFuq7yFbMCAgL0OzZRZGUGH
NWUNmW+MiWsg+4lOCmmMVWn55ahp0eygM11MoUZhIjdUndZ7iIWYmiF/HdCHyhVs
bXvVUOhx1BYLC3SzqfkgKe3AYCM1aRtyDaOjcl/NsEMrQjARiHFFa13Kjjc0Y2ec
OjR2Anv/qq909jCarXeTjhTYbCsPl+Zv/KcBZuBb+VEMvDUJH5yLlnSIUdF6sa5Y
uUTjQzrNOl9BCmIFKqxCM5GJJTPZnS6LdrVsXC3vjxP59HkXqfFe3BlE322KBBWe
Wqy6QMhpfGH3USidnNdwevl6DQmN2BrZ20MQ0qKXtFbrIppEH5cfk8to6Y4lOaY5
YNikotYYkIqHUXuycFdUWjJL1EH2u2bNQ6RD6Im5aQx2QAUFhBpfxftxrt1Kn+QB
ND+DW05U83cm7jrUIwEGkOTZBLxKuZKFkmR2+H/HYbK2/IBxMSyhL+lE/3vgOaaS
+17qv1i9xRA67URgIwAj/Ubdbwg+DJE7RQcxSZ4LZM1QfKNS6SOxAvWLll0Ij/PT
MPaOksaa9EbHGxzcTOyV3gO68Iy203HStjEl7qKEJOiCFk6pIDn6VYIyrbOyjvSH
ZsN7BlKF915MsGZ5MsBS4F5H+LRcd1kIk/dFUCDsFPrV9Nes5fuA2Uwk0GAJ4h8Q
OsbtN5IFByrzXRWX9qERUtS10D+tHSyjjI33dd7k/kTJ2HcgKLiDXqn7kuc9Z7Xv
/f/qdSnld6sNlBiJzlkgWmSLlJ05Yh5S94pZCVvUPj6NsXUYaPd7N6ECsuyD1zRu
rpvvXjfI1O70dQcj1IdceFME8bJXy2ng5oVVfabe6u/iD5ZJOtgDabrbfhYD3uEf
Io0d8mUPGTUhzzPM29gagAFF1MCGhB4c8sdkMfZyBLWoFhDc3TAGMq9qDbUU5pnB
rsceGXCyZ3pFkXjD/asndd3ywGOcR/Wq+FOb6O5iKxJq4EJw2WuHT6fWXn/1d9/y
1qdURb3KADzQ3HQhEbc65Jp+ZaJhkJ8HPzajQzEDTvON/amXoGckJIh2QG2ad0Fv
P6QcGOe1qQgLxvjjGWgeeLzQSmdAkH6ZHxyJ/rLM0Ztobz7/vliUoxeZI90888x6
68yPJzVp9KaIw4SpQIddBqeI9H3ANYu1oQNYc4QK47XnioybwAK20hXOQSp7aDNs
7/W3vYByhMZV/z+mV4IPbA8vzdBg6O8TAvD3b9Tq/1uCIQJw6RDESh3AkQqhh7gi
yPsw170Cueuw5ey5pGaLxRgjCfXDJXoMhSZNzwQg/xqLvEsJpp/2rKhByScsX/Ed
WMW2rpRvQgOO75y8D2AFlGnicalxwJB05D/u7vn1ojjf6zmgEvE5GyW9ZLYYj/SC
FIhUTBO+RZWPx4TT0lNM+tjIU4WCFOzpSUbEIXr2cZ/zEErSCCcdFBd0JqcM8OLM
YO8bK5XOZK3YsDT1hfHPARstKzOdSM/CsWtm9JDQtzxbWIPBOpn81SsGU2+My2ik
61fJLJyqPwnb6YkedwnIvMHAJjTU/SmQGEDBklpGtfp2Vtm8/thI01kfo54+WLfP
paEAD7UUNJWBCq0GemnPphUa595ghFgviKUltcR2u4W+EDJXquVvHtKeOt0j+Sp4
byAr2YOsGzDM0QU23YGbB+66fLDFZO+rhCEWH2f4I79gzG0162dSNs5p6o2KWZJW
XycQdmMe/ZF0OhSmk4QvLPkxKiSIU11uhKEorbEtsMb0zPWeHjbboz/JLhaM1Qic
/Jc5RXVtdWl3zzazli9Xg+C7yS6oiPlXccSmFxbMaGELxBDL44ZFjc4fpXgrSxcE
POyosmtUKGXIVYRVRMQnKQlGLb6ZtMFPogbzr7DCWBYohKXaxGT9A5DL114tZ2ha
v9wEaK4wjoqqTxmaa/cYNwoQxoIhPmooKRIkxh8Gbsr6BwEfgXjfiCzihnmLhP+M
RzK2pU3fJH6dnCmYq9JsD6IMf6awo1AiaHj/hWOPrSxSfDGCcIcnzytJ8IiRd7BA
ARqDhuVYDgaw9Yc442IGOKFF7V0BrpdkH0mmJGeY6RMCra2pdfCrIxQf5Un1XucC
8gdJOth0M6AWytSWQXl9RhPnTT71mlCHhVuiVrgjI3hEcS/XxVMHjOu8oB7qEvAv
aX6X3RfeInb0LbzJVZCPoDqTR0ugxPlc8ICNIRY064z2+xS59+eKisIyr0r++OQO
blYpygXtrDT2OVLopAIGmSCAIv60OndvzXMBqlgXMLyUAFzurCT50mLDue1KIMO0
207znBHAqdVSmW1lTIZ4N6wNK5dASHRlE8jO0a710hYa/FvpQkbSTuCiX+MN4ii5
/UXT3wuPrleD7g9PMwccurWxbVuyVwpneK3lsh4dOq1g26LoGdcbvd3BDTAxa9Jq
vwT1K8wG5qVvx8VOyKrm04jQYJF8JiRBSTvPj8EjHqafnvVkOk7qlLUWvg/7gHEj
4Ksyah0aSisgG90rPvO88UuT840u6nTA/0se7riA56fOpYYIwF0FQKaflmiagHL1
4eKHeFyS9qalhjitrQUSLs9wOY7DRHiXNztwiUKY2OM/n1bBMs1/IR+HZS35akZQ
+pPZ3+TQ1a5/XkbJDV1KOvR4Vpmx4pcWoNQSuSgrU6md3s1Ay1ZBOKVYii5EcJ5o
ZyCI67CkBhHF380dUTXfiEh+JBokNibekf80Dz/beEW78JRLejhTEFDUXQrAoFJs
a0IK2qik8QOaAfud3JSj28OVwSzFtXCW/8wje44YMPILDXUZnIEHUz4ZmZ+FFj1g
H4HD9N6h1ewQUIKlwodPjB5ugAyq2YQZd2S4T998RMaSGaPeRfgCLzZHtRLKjXTk
uGpJzebK5bDUxbbjC03GpxT1uSrbU47OAetfcc50snusK0crVevC8U6Uq+EEUoEB
NpPuANTlOt6mKtwgq2a631JPNG7oH93hiuFP2iisXC6qSrCitxlTbues3o5pxAp/
R3m7DfKz976QUWNzlG3hLg/XOJz6cyxG1qmvrTVLnh4af2PSBkm6BZn+3qdka99Q
Zs8x8Xk1KEdNLYsyqtfrhkmTLw/OPV+DuRvOPsZVw3AhUU5jAp07cvrGp+9E3KAe
Z5n+kWDPDT5Xqdr9u1r0yvpkMQ02+s6fY/rhkYfgbAQ0dVtjJUzkBoEUe7obRVqo
O717zN57D3G6Qi35HEL+0auEAWhdmWL3YPspGFFVd41kwedif5z9nJAZqSDwWgt7
ObfQOiOYdtnCdDMjnpwvb672jDmiRpVyEJBeWdHLW5d4MgCRECON5NkUlIkV9LZ+
uJrYhF4c11dUlidEnavWoLv0gn+jdaXr+1KqecOKrdmuVabOA2xybOEXqi732Ne2
1ZAk08tciL2eTarBFcISyETr2CX9+Up/2x3X5ewF4Y/gPgnmifNf4V0SjoEKTwt1
nWCM+tFhVYUyWqoEYTce9CpKhlenaFlWbnwNrV5bNk2JtE2E7TH5S+k5y/LenAO4
qljQ5N4QCr/MrPckxyUyx9aAIZycgTCynnUpLNCfx+IE5jbXUGdX4IIFVL5n3H1b
w//W4+35I/iMR9g+L9PTxL8wzAX4GxwWzmP2lPKqzfJj1z9ZXL/0qnfl4VIjoLGx
9dO2R6X/udE7ujTN6lqiPBn0XUeFI3/JF5WExFD23VFEI4CfaosvEpFmiSEGUVmV
viwSp1Y8X0uXmJRt9FqoRX8VgsE5wK2NbcDL2mH4eE/BkMa4sArFWEJi1YSJSUkK
zRyr+WvmDyTBA7uHZLE2yrBKOcXYd3Q5S82b7q4yQnc+31JhpH17JzlTE/bkmwlB
luYybGkgGcHKubs0X5ZDKF5P+PspacnnabaPwvd3ktzYy/SFUMMy7Sg3P8PAtyRy
tQDcWWadYm8YbB805P/0NuILbAO8VjmnFFU2LcbPqXMl26c6W5dBP2Hk73eZ3hWo
bL+y+xJuhDHQnZ2YqTUzwa2ga47wR3aH+nEJnvi0HGlFdlVuWmLLWE9kFYCmPX+4
WhrcldVCl2SBCUWO9XqRHmfk+two8xNoqZ8jFouCh3EaxkJZPZL30PyoIxOAbgXr
Q1TaBJY4TUGcEc0Z1DrG89yz2rFzKQrBXc8OSFrTxWArjNPlCwE5bZI0VQRR5wBm
RGZWZIDlfEnfGTyiKAysxhWcUD9eLdQqf5xCKQUvaF5MF+cIPgSnNU9TPJiOsm44
viSN2XpUpPZtgh6KU4KKbsfYLJ/TfC8PPE4oUleM8oXHLyr1zi1cKytUNQpwWX/T
Jor91QLkHNDRD7SnlINvshCi3wrVgMTJOeg2a6ac3NvhmzPrvAHD1G5DZAuz7ZWf
ANL6QC40ePYbtaWE7GKe+A/UnYkjjjhu3NotuAcjD2NL/pRkYJ5rnQMG/IWvnFq7
BDTdWhn4JykKLoR6Rcb3pexWWZFsTw14u0ZAjpPf4QVZKIVq5RZLzo6AsmugHHRz
BGSVBihxbyus7IoEAvnm21MRVxt8M0M7lSQpauFlL77Mqonwrp7GtiBmn6YO7/PX
ki48bwawSH2XG78grmUj9H+enUcoCS9maj80n2vi+/qa9poTYk8tIM610Nwxi+sw
rgA6B1av4SeV9sq6cws+/sTCP5cogBVAXBiiptMxpLa8ZcMqqcCGsJ1hXLapbedn
Gg49pJFPU5aqGag2IRDEODpRZB7WUfbCDJXAr2i4+X+PAPKSob7wgCWojG+O6Ohl
RctuvUYj8bZ63gRLJiYvyaATzaJlOSB9gaHohF7Fx5EDGlcqLXN1UsLEoxVb6LTN
qLNQAdcBsRaqNfnzPpAZuN5Oy1mwTPPQh8LnbKemV0lcebYyLI29mBzsxS9aiH1r
v8qJcJitlVmslsWtlM8+U/9UKTJFNWVkiv1nj/MvMKfsV4HZ3242qTZhvSKj8rtq
DLZBwM6qDUu9uGbJ97jj0pK8EBvNzeCejKOR5v0BewWZkHPN8Yhf3uexyRRDXpTk
EVp/g1ra6kAjrCg1L/Qvh66E1z0sTZLd/84/dJF5kIxmHyQvGmcdZOdzz2uQKuMJ
yf4bvQDFkeoFSE8VSNWET5ODx6z+2dzvk8iAepZr7gL1qZv9qGSj80995vMDnV6O
sSnF9u2R9vA3y/U/OfK/Eyx3EjtxLZ++FVBd1KTdxXUp6fP3uTRDmRPgI/Dtq4Zj
e052wGTZQ5JGC3KH6Y603a/Xv+HlLF0z3CIEdWTG7bOCpBWEg3Jvh1HJBHSpEuKZ
BV3D4ZocWxLDeJA8CLljz3AY+XM3gq6PxN2jb1OFbeHvswMya9iLMqMKGcriTIw3
yPT/YyioTyCIx+ODCutgynpUpuTSmAWNUag6pBBIMoiL6yX2JRjzmxi9qpcqlP3Q
6aC8G/YsdOxsx1IwTgnfM95KT5H3uj5QuTR+jci8FZpA3wzy7OYX4xg/7UUXORNi
m8tCbteqDt6nofBAiq1hznV64e4jRd9HpacXMqrkViEkKz9jOhWSi4KrCZWE1sug
IIP8loAfYbUpBppHtmL+fNRkxr7OIX4n6LoP6nIky85pTavGUCfh34SjpZT4mddM
bW9ctqFkzqx1oe2MhIHrHFdbn/Pu0oAQJXp2ycdyqKNVQkOlpciSB0yHJ1vAxqfc
vQHOxhPOQsXfZW9YTPWJB4ShpcRfo6wza5ghSQoWr8MS7Co4PrsBQ6wn3iQBZYck
0/AvDD6DR+1j/UityFXTzA4PXrfLl1eweSb7Nf6UcyeJH+PlCaWr2ERLkCXhiP/7
iFtNaXOsI3DLx5SncjxrHk9wOg/T0f+cDBBDvPFFYlgOKw0K6HRi+WkRXoC2kMRZ
UPYZcEd6d+plWcTGzC8tpgq+LJuZAy6i+T63I6rVtLN7YXuOB1iJESHlDumHbMvi
muQyOZBr0tQWg1D8Whr9Gf08uzkWw8oZNSR7NIOTye6UOvHvWnMVFQ8Gd3nt6NYZ
QXmJPIWjiHBIJdbviMZ2xN6DxskyigjdfwdPInpUvMZRve/5xWgFr6e9oM9jcInj
JWUt7d4mdttXjoID75vYjQlYv7MZMHiqnwgEw+pRMk0hQwq/GHpBW1faFtOSGCbj
DqqWX/C+r2xue4HN67jnvnNNgmEvm4kM1AKZmBx/OmuXO3gfPYi9nESUt0iHc0IV
4Ec1Ki3gNcwhEg9d0Yon5MnmHts04JXbYS29eqd4W5CeU7/hKoTj9ztNgI/LrdJM
uI2sVAYUn26yLE4sI4t2VSt3qsMC/XRM14tS5TI1bJJAmR59V65DM51ShGWOi1J9
IzbsCYcIGhuNziuBZLDnKg8PR4n5j1QpDz1wtu4Y+o8gOAnAKY33aMfslLFvLQYJ
S05oAyyIuiPKWO4lutYiKcmGegb5o8i8i8Q8+fla52YUrTODxj0GfPmZKi/Ry42B
Keibeag7uia9NW36v4J9rKvZnmrkStO6S7NEAeSm6qoUUjh3j5ukFsnLCae1p2wA
1FMu6a44SAjCutuBzhtTdBJfKlElWlw9OlMAxA94shU6UlkUP58821QTAUt791Sv
Q48O0FxRAysUy1Crqu1BhGS64HJ+hmm63wIVvfqYl9V7j7yLxwz1m3dwPHi6NszD
8mmuLLSQsk80ksu4PLkQyhfAjrqZPdxf1mFgQss76pqgrgOQXzSeOqNah7IsVM5y
lTIIW4Umi7GuNyAAQco5rTPLkP45NYkZQTwsAVRsbdg6bAHpqg02iMY5hzYw0un+
A+o5+W5AEb8I6LuctY5yS8kUIalfG32LN+xGu8ljYRs5SSRac0c58cvXiVKWg6gy
PNX/CgHl1PwWGlNEz11ZErQdrgQeNBoFx0+yonAnd4qUuL7jkiWLviwZ7UyJAJqX
9NycFuh/qzBnxn0Woy1JXolEfGgE1FRINmSHEkxg9d0JT19/lxq1bemnqrIdlxzG
fNs9WtTg0bdBdGRv4HiLzEWY5My5+QXFbbe2BxnHkSyQzp/yRE9cDw9xfUZJ6MmR
98myBnZpS9aWEp53vNigqKT0Gg4T3JCf1fYo2rNSQ8rp8jjitN131axQSXQqLSSw
NAz52wNAbkmCYjb94VTwBp6vcIZ6d2QAFAT8lfJdv+5/ogfMyC0vsReHFKUi8jBF
NGJWZ8yaWJuQhU+tkoKtcNt0GEHyJj3/N+XbCXnwhGZNFV+7WUEiwHS3PJKE4AjY
BBKJz3nWmAzrV0OT5HjXPw37EvW1HKZCSnEQJvy4syAm9f5HyD0fETHHoQsrdUpw
2cGKn2zTtyii3aNymXSESyBUYGSW/iW6OkaUOVLvUaxsevZkgbYtoYvr+UUQeael
csmLr+JwtVIrGlhwj/5VMh49ukJ0Oitq2qypg1AquTODUUM+EnX0VTTLe4Q2RC5e
UzP1mtcaSW8Ds7/DC3PqIdi0JGB4gg3ODaWPb8ZZnrHQGkZkQScVbyFShE0TCmqP
ctJJIHAWkHVU+1vjX5lTIaeKzZLPVDTr3UbzT1/ceBJOy6ZeGqaWyI7qS8zSFnu8
iLfl+Zbmh0q9SFfuxAHubWRoVl04nj8P6uizOTAkRYflShR8xAofGnfkMIUR16pn
JxSONZzdI6k8Bm0SmPZDQTYwUjFCuJYKBxVoZO4qvAjrM5HMjNN384v0wi/4OCOT
ybSKnOKXJz18k23jmTN+wqUaeXP+b6H8VbIXnckdLlR//OyDgPWl8Uck1TMaPUmr
oNwqcn4JaSqy7SqXmREzikAA2EJQ5rfq7kNjQKA0jQY2x+xMyKU/mD8/k8Xjv7C4
VGue8sp8pjMuxcWvkBGludCocpfioeycRxeCoiHvNxfc+rfRKZs8OdCjvN5sn9c7
E1En47Kava7e6N1iOHBHn4ioJPOyQbm4lJ21yepHAE45cZhsqqaHw2F7G2L+pzHg
gqwyAARbv29NQ579bZDJ+XGp4osGZnPlW9f33ornBY7abJSI8XzY9uv6H6f6bJIK
uEnf4VKfX9aaUZtQjMSUMjcOdHmejpS5RGCtID87QU/wcanq1dnwxCXb4FoDdttr
V3xvJIkryXTU4nCzpuHgGtlOMFA8jwNBqguZAwVeC9g5ulJgJcWczuWnCyg2WKn7
H6okXpPzFoW25JacbEp2vT8FYgUBiOVeNBEk/2s/yAq1bm1+xTJGITBF/SA6E1KF
zM/M046la22s2KRWKVCKykUrqt3EWX3jWaWJgnRYtKx9sEC3ymMLrKuxBFr9u+hl
TPhJ+s2v2bnviJUFm/F1AzGUfgZ+JR/sUz1Qq5H3g8aamiypMBb9JSLCaAVOg0CE
Km5XeaH+QbmW6qdO67NSazIdkzjR/J7S4vfGUOg4qN4WqJEVN0fbO+PN1V+dJlmR
XFsOlH95swfdsu82LES4nKLapM++pqL9lROONZw2xJs1Cx8QsUKP6OOy4AFEr+kZ
+nw0iUWNFAss2CsjhXezu9PFURtm8jvQaNJsatl5vew7YYpuTay94lF7pwDgLSDP
gFGhbCPw1fw6oWVL9ehO2mRxMhSQwri7z3Nn4n21S0mQzGxd8x2PihzczcfNKffF
xhjrFksU6+9hvr190oS5GuCX2XIxseplnvm8IRWgOVY8TdL5/lwt7cZCza7ORtYw
qes5NHemg8LMGMIVTYLm0D9P+zTUMcydi7wyZSI30rVXz2VKWqOf5hr50NzNzjvY
D2y6ANXu7MTGlv1T6ExOJ89o+RHeAeCnq/bOI5Kk2rgMhkjG/TAI+psz3PMUqR/r
FKMuPcxzsXkTehiac/lx1TbAiSZ9U7KAXv4UgLjaSifCxcOBF1L6AigPGbYqMp5Q
MuW78/evU2/PWYS+GHo5fv0I4z27BlE5VxX3N35lc2KMAu0qo3BI/Seko9Gmlznf
w3fm0lKvjc0cwINmrWEXD8IeELdOOsbjnvEmi1bTLZ6kxVabFK3EozcvRl8oS7T2
6TOYHlO2a3gYkA7abxUnbZfza80Ll7yJO9z9LOusAImv/0FifDo4aRjtuN4UTmZd
67TRu2+yIcKNWR3KEJNpDhKiI/2O7OF35UGEcm/v880Ldgbt87/xQxne1YVUTr1/
7B1hfX7fxAuPH3wiONQntICY1VqLj7FsrLPY5w5qOqWeWgXxQuD5hcc+LgLIETn/
Nwt6jLH5z3Ud2aune3jGSSMdxIdScFg5CnvWZ0lCTE4ps+pjAsYsjwkFv7cThCMU
Zn3zSeRpd6heguLzKzDBEJb0bO3zbhQ4TpV49ch0RJGG0Rrb0+8hLl0U72r3y1GP
YEIef5xHQrSQtM9olJfBeADzDjt+uLlKYU3RPK1gqalDZo4+ATiFAlXL6am4JRDw
azTr6Ev92xYlsQv5P8Pglp2YL3zBj3L2lIKlcgQmbr2vQRmgrbMZVzMzLeYgLEvd
nxHop0r7p0xthddRBmW+6dJzT+1NUmfKDHFBRZohaWxLVjVsne2KE6Gt+AlYffRb
lD+bKo4JdybkTV4hfy07nHD4P/iHSyI09rTbEhyXTqDOdzbZV0Ikiz42vrZ8mEj6
+G76w8DidnGg91Fy6dlnGWPOcS5P3ttryWATtI2aUWqv59HGerEVfKnp2TO+m4CD
uarSpNWBp1E9NobSwnI7/UlQwkeEuQHHO8fyFXXVBOzAfY0+IKhXaiSeHfIRXVbK
35mniBbfu3eTs+bAWIsxf9tH2a9DAbGJ+jUF3HnR98pH0gQx7pbvJStj/nDgmtNj
ooSiSUHoEtPYx4R0AQIajru2AVRPmvbjMk9OtY2Kn8UyqopQ28aRs+1kdyCAFvOL
u9zXPFf1Vx+IxSApcoZ9TVVhXpitKu8X5+htvjzJ2sRNvE/NuTJINy4/lvu8Whwd
pWwgrh+lGASxuG2QXbtqtchn9faTnOggDHxu38FhEaubdDdUm2qCij1IlisWeZPC
5yvbgPUINjhF81ItIKBmmI8GzpgOy2pzVE62MmgWWEpdwXHyOeNDxSTSQbM4wyL0
Zo1fFgiNnTHKhI/cQKSsDis+b7PGIJ8mjpNLqghYgTz9gzEgQzRrddJfPhjs/Cwh
5gDy1QqEVb2MvPfTSp7YNpjQmUyNx3VNil499/3Mxx+HTSVhBWrtCNMIX/BRX/aB
pPLa+63vurUr/ec/0Py/1Mv7FxZfJCo+QtpDq0IES8N9Ez5JraDktVmZHTLYloRg
xKfUy9ulTuw5aSGDvsem0xGOprS8LYtcU6/tgwqu/68NsrhqAAiuojYCNqky5C7v
8wCygu6owRF82YdHBu6f4923XaqmEIDZOILKBmfbULe/Kdndb5zG5OhsBwynF37V
kfsDujMQwnhdrIzEoTpRJW5aJ7giuEU6WABYn2pYRWsbXfgQ28pDRd7cx0xrvEfc
Ud5IgHvU4bYcKLs1++5r5gFBooNfh07nEl+wAv0GtVVzQ5o0Wams/aZJhcDYU6A9
8Sy390cyLgdceiqtPCFgPed1m6NEaFRCNzJ7k0q+btlADfL9pBsnRH5sxIAEnw7J
t9Dt7TBaFI8LE/2Fzk4Wlt5S+oXqq26JLd+jBRYY+zmMdpvd2dbyhtazMTmECClr
m9gIKaNrZ6ZvuvhbUHk1cgIWJBlVL4MiKNbqND3clYkfSf7eZYLxpMRXXTRRtI/M
tsElwVoBdGEvdEq0KODDavH2X72TDVDiuSZ/6RW5U8dQdgASXyjhN93335OGbo2+
ZOebok8T1WRQLvFNA1MsxE7DMGKxDUy4zZ3CzSEsWxHxcWyMRyugEM0QAH4MlGNk
4dj1ki10TD7DtqXg23nVWDM6MXZdQA/cJbkk6FW0UkxA84VbBs/Kb1YVyz0N2EN4
oHIDSNf8g+YujlREn56vgLO54vQu3kEE79PdBI1pVOUScV7lHZ+d74/qWf0ptMZa
yx1dGmRgL1IVNRo2xQjNhOpNmThNwJ7ounVNwLgGzDg+yOCI4/4XzpKTEOaB8zZK
PsjIvI1jE0ZcITEVDXuUYYV21x7HT4EnuP1kiqWrfHMZ/E0epPLwVaq59+sDbV3W
iFDx92x+9luhJya9Vj6jGHtRXO40pMhiogCD0sJxHsD86b3Y1saDAN7UnEc40Px/
h9sQkzzheGyudz6je+eGrJ0c5IUBXa/o+bcbY7mlyhqQWiUb9sYwfC/EjaFxrQSp
tZ3qjoWhP2+aCQFGEDzksT3VPd40l2vhplks3yf8gi55bLgwYNJLdQP33CTrkfCH
U9PCb4yyaRT14Ymjq1iGym7c7hr2SV+pL7ky8cLqs7BFJ1PDw1gcyuxQ5Avvp4wa
TPhzx7aiQLhqJGGMmbQmF3cMaRi3Enkzde6LScsGazLyRRGtvMAX+TIAU86PEVfr
rp3L7f5lMUm5RUfq4EOyLXs9yRXRoIWnUJXLT7d7rr4GYCcuAhlFCUH33asrjy+i
0S614IiJPFXxGFMDhR8CE8mOaCu8JDnrUEWCmTrX3yJYcsgUtj4BBPXDditFm9f2
kcf0mxqLpGTPe23vmTSozvZA13P+zyFcKOgYKupmmv8ev2baKfO12PInO5SQJbng
mTuVcMLhlYeAJDoaTzWnxlBp1JNupmF91EuvnKpTrB5ouaUSkTjAE4F+QPgR//uY
9f61xLkT2GyAwFZCzBgPtoXbUgzn7Tu4dd89gfSD/RTs1xKrxXb0PpnmHUaZ4wGK
UgDmOF+O8iq1jxjjuFfzgV3Yiksl29AqqwcCWXvF/uKrqQQ/JP00NdE6GMlzMfgx
AbBIFP61mTGlSPlXa0gTAzO4e7qYy647EbK3p0Fs5YFmc33vfI0j5VijOE16MwWS
oXHvjRL0ezpF9q/LIrltu/DHURpstssq5UFLy18uwIzTTltbmS3nvhLCBgA3FoYo
Wn9i6XPGnRhCfckWchulA9vfVRVBNoHJW4599HLvkDudYO6jWhmfdqZEUtpArID9
ip+M6Gt0JKfcuNC1UTsCbzQyI0wewpo0Yd4fmi5v3F+rLd3l29W/ycRq0Vdit7iO
L/uf2QnnkP2iJyqWISVva6naoEfCKlTF4U8DLXS/Xy2J4z3KxB14xYa9RKTBIAE7
vhGvhF3SKvUX2GZDPvYvfhXS1dpiOLLL3nnjYa1ep1NMYre4pkpU3qDi/uOZs6Xg
g4rNUAnilQYiUYftt/EoBptrLEmLl5hHmdrz1/2rW3sl9h/1VTmGRXk/8fEQUdGo
kjC8hYK9U9JhDMb1nPUil36sU1zuRUy730LdX4Ko/lIBsquH2fRt11p428RCVlzi
lHOcyYG9TeonrvJc5g3FF9YpQcETiN0Y6yj4AVc5A9EdLQGpKdpr7ZVYv2lhvhpH
uVXrLnZ78OThUD6gwPpPCc4tRisPutFxtzF1kXTfUu6aQUuMhWdjOjpb37Wr1Awb
iRZrZY9JLOsbC+OrbxO87z6EMX90I7yWs4uS3NK9QA3ozMQiNr6j0UY7gZSMG2p0
XTLYUVD2zTLJLoLjR0EdVVkudMP3oaszEFhGFNu55MEl9nmKL8MDng309rOis+Lr
SnOVjjiZ3SEBU5O0IoDt/HmsBcKt8xDPGpbG6Plcdtc4i+7ub2R+aGQI8RomvsNU
VDz1qV8FXutmNhbYv/fEChyrRdZAA8yVh/Fhl9t/dbpcKEe1Yoy3HMHgGEB5cOMN
SRMEcZL7elIjNVBsAjFnwgFKhC1sMbZdQOgPae26athy09+wvz1CZEvAqCKEpwHD
7n9ovkIZPi1eiERI9xxZvlg4JFq8OKGv4Wna91J2GFQHShwNQPsv3+NKUEFaa35x
BOgmaIjSNlLxAm+hIgbQh86hkL/blLqIPtySYyjnOdYHHKAK9NdjscOVctaeKuHJ
UGmIgfvW3EUzrNpL55DW0go4WTTodfAS+Ddsx0Wh/Ch/ROQLDJb1S8bljRCCgZid
OoiRf1Gir/qpTSuIX3DREHxQvwiylBQ0rA615V/Kf2WyA5ouCHM9sJL49yBavPun
0txcnp3eilEjnahu6Ukx1L6pCY91tDR+L5mEc5jYN/y7vWdNgrJess9iN/zTRNq5
Sl+PHnoixgoqz3svDzBeJ/6gO/u+18wvMqprQdAw80mQYKdfjuNJOIiSt0TeN8NZ
uH8Yud052bbDl8XfvV2rnRVVY6Edxfh50gObsWRqlBsltR0KJDGlFA5RJ6UCqGak
NxqdSm3ZtRBNXNGd87Y4EznmfjB+ow2wi76IPCo+ZYFypQdaMj1mdtjXtJveyuJP
7KDbFwvV5AHkvdeaxf9zMYZYhMoM9V7YpN2AK5vZVO8xAKD+P8l84gJX+8rzLEGF
TrvBMt/aotnW+kn4gpdsSUwdnJJEKtFOkB62FAOn9MK0rHBt6APBZ8qP1OV5LtMQ
XG9Ec9HzIvW4TCL7fOA/bvbFZKugJUM8azPTetlUEAfuCuZrjsxufB9FseybcSW6
46Tc3liCG5ZC/+pHhpI9Nj1sLB2b34QcBQblkdadhR03HRfgHY5Yzw1T27J0SS/B
oNNEbihAjvHcG7duA49/dxU08siDQ9xGVu/JvNcYAoaWGXYKTv/pCj33+z8X3C6r
oOyEfLxiZgROtQL9lf0Qdbhee+LkQfiBKgZ6hFsQo6F/PxkjUmz8RlBB+fiQlC4j
oAIlNLCf+6RUy2Qpn52N+uCzyXC3i+frp+cmFKhvH8C2prZ9VlxtIbLtE7xoVAUN
ej2CYgV0Ub6JFTT7fS5htH9IuRZc+7lfjJ13JIPS5Puh+wG5UQdmey0Z0CeBUn9d
UlT1pm1rnp6IoHIT94M0GQHrDwY4gGtxTY3hxqeQtC2neoKa+1ep1nRUNrstRDsz
nsYAGzukH7jb5ulpA2X11DAvgprJPB52fkNW4K6EqXsGbI7HpHvO2Q6b5NtpCIqm
Mw+t1hyp0cehYcldYMM5V/w6/GNhXEqIJWaJVCmwvXst5vqTNZ7vDj7O+oW9B++j
i48/VF6R0NmPvb9Z6zYqS2UEuxSWGGMut4jH2/0SLMj6VmCN793CMnhalFC3aawP
7Ng2cLgj3UOvI544R08dIDCjWiMQQH7EU+LIAabed8eEYUCPNE5wC5LWGsjkJr+k
8Td5/QCpjmBhTQtZXys+EC/nnfPurV1sBgtvOcj47iNMQir3b6fzrQgdDu9VSS9K
OWyiUdYR0E6u8/T7W3nTK5CTvu8byp8ixfXp9jUhIC+Cnc75OipExm3hMVV5Yh29
JlVVryIvl9yAuB9ntFl6xEMVU/qjEn7a+UP8edI6sSve3dALZMMm2qnkVIGMJ5aP
f0EiumboPU38w4OLbV8TukjhbQg2Wtmo2b35ZqnzjOyuopNOf6smdEeOwURpoL1m
jG4LIUcKw72RCUEuJpTGsHkPIe+65BSU0AGbjeAMOv+Iiuv1DupDlSifPtuY8ZDf
ZjGVE/Ea629Rm8xTPiiLgTfUgWW7zkjhpgrGTtAQmcN1doGZaY9nCut3n6452aKi
uasmZ7Fwo4i9visepW9SI6UErC9aaUOwjGgJLrY4rDbdc7n0x6MCyGrwDSkKqx/i
hYdwDkh61fhAmJ5rQcmP2rab5XHGr3vSaIluB12iVzkbPyI9IlUn0vK73GgEkAlA
IeMiOdTSdeTL0V3bJ9FQ4aAmD39lbQ2PLRegBUZRmVynI37jkS5sNT41K56MFyKu
ywRHuIwhYrD99RstAchHYiATegjT7hVR7IXCV+2rrTxstPPWk9J0LueZ3pRHwM6x
6hVmIuHWNq22MGm7Bk7qEo+k3PMfONl0T22r1AxCe77+dTX9qjjyBxpiXIRGf7Zs
JcoHFxNg7rB0x05GL8awV2wM3pWiYxiyoD9xjHkV+xej22Sl1ZUsFNwXUDVF+0GC
YPz+vKyRtGe+dUQBJSAtxffFejsJSNBlKLcHGxvXVJ+1vnEo9LfszUQyC+USWmBJ
IScfvSCHN1ThS+wui2SNiFizRCDeF+NN8uyRTeQ8utRtgtllnhqo71hN3zV15U2n
1MOKBhLS5SVrfSh82aAmbqRg/UNFfsZ2rUhhobJDpAfARZOb3aji/fLje9qgVv/f
zGjJNf3amohlngCiRfyXNtEA5oxIcPIZGX3vJturt+Fkpe5gFNaa6WUu6gp/AbbC
t4F6Uz6AMTINDezOEmeyB8BM7zw3P15nkhj/+VyK7iruRynTxN0WFZYybErxxrc+
WiEZ6lo7QaXAhkAUjMxlWYSuhJgVaULYBMLhf3+prPZHiOQg+wmvApftKPEA68WM
FdtDrxfP4edPsMDWWd5XDYwLNZCp1/DItJY8eK5NrXta8vJDkGU+eVRwWJgA6VfN
9Tu69q/7e2aNieW++9hdkW5P2znZpNi/ixlDbcmo33eIuNW96XoTco3MIsz4GeSr
Lk44w6OpOvp+Y8D6y5+n7OrmCdE8yMBNRiAnb44HUuW1oJ4ge94Sorr0frKM2OIH
c0pq7gPFl68qI185UIfS/ljnS3Ka28PzKE6tNA1lI6Xip6aqhS6jIga9B/DgoYHz
xmkpq/K3FRHkez/mPEYRsysStLhkyQXBdvALUXA2fZx9CHtFUmKMhQZTrvhCFPHQ
ilM+W9c5imfVxzosRCoJiZXeVxVfxVoi7vuSiylaZqUpopjUuKjdQpefJx7d02Cc
wwxGfKgHfP1Qh2AJ/SrNrMNHBsWzKY0r1mXtaTatgwqB8p3XKeiSAxARXwsdjUE4
K5Oc6dR0P6KrXy8OzlypbsG7tiyMB9Bn7wbu+0KYSSyGfTfJpQFrJOF8wOJAJKGU
NBZ/iGTbW3TDevpEi1zuNvKIWJuh2Kvgfi8K8QsR7Mag0zSQUO9qd7eKlvQSz+Wo
9X+MnbRB+BYfhGDUTKIDSCQB6paM2/wv/Wnz4O2wk8aYHwzmRvE0slgQCJbAbjly
Lo9pworxb8VZkvBjVxjIZrCZcWlFY229Q/6Bmkj84iWmD43AH4TCX/Yiy5AxfAPA
md4VGnjX6Pyx9r7n/orAppmSKrUJn6Q2ubhXUMM8LKv/Rv1TXMKE3ATon9yVkle9
P9CPAHAEJaIxJ3KoGnGaYlAuGDQG/TWcnCQCncx1bS5yH3GN77j96evAIznqK9WJ
VxK8T+Of3tWVTNiD5ZFLgpY4Ca2wct9ODaO9XQAl2JNKPJ/7DXu6Ext0nxIZVwfl
wsNB72o5A8uuTZDsEI4LYBHJCGu+kfxO1/LdC6C1olsrIcP/xNsgQ1PIX22qS3iI
7XKHE8SOzeWuZPE1MG/JWqmJDKhKBhUdccGDVvqIsBoFyy/vVovXwv8on6jcncpk
BZ6r9ve9ztdLUawnMCAqgoslbHaWcOYPOsUE6l/H9QvGlClqrAAymUELM0wUDIGg
7z2cKkHOslq8g4x6r6or2qmM+GCq41gPkpDsVYGKadD7H7d20X/F80IiDpJIBBbe
FZNYv69bYVftqYqMWxoXq25aK/sijGsds9cslXUV1Wx5eL/MQCfnGSE7NnPyQcw7
55YVGqGHTUFgkFiqsS/Z1DRuqHuK6IrffidYUQ/saW8c+IzGBh3hArH+tnh9FgTl
7Yz/I28So6SLQf3bQlia1cFOZB+sbp9ePQcODV/Ts3f2OOVlDjH+AoQmBd4kq6Tu
63ZHFUtk5NMdPIdXYYQePGOV9ZN4Jb0twmznlwrM0yRLl21R+VTgESEkNCAFuDtk
uKnpQaGKlPKLVuYFDneSmTRSO+XzodCnqef8kumuD6aTdAmWIzAQWlZGPI9aCHbT
uwzOFNrRgCEjWhpVh5qIn9BlRGutYSjYk9XHSOP1q6HCPvfHQIlJV/g22dWg01JY
JGIwaNiatcCHy5pBgaBpQZDTtKwj1XoLIMg5cZ8lyuqzQNjCFBmqQNyW2QPelmSc
064lCyu6bB6uywWWAdGiX2nMXKj6P5Fa9HFm8gjHqwF9Vl/en03e31ufA4DniREB
VU9/Q7A2WEPcwe0Nws9T3+J8WmD1kugTWoxbRif/msv4toDmvovoc57OjDRUi8r8
CoYKeLR16O3lxUBQCV6d6GEMwP8bGislc4qq4/YTEys/QL+gIMLLTjKWMVVXZrTB
HUsuka5X/Wqf2mEjMTqnL+duz22s1Ou4VPFNd3NHi2OZJxtCfrZRsPXrNt1II00I
QpTPGox18ZIdeGjUIk8Gg/NnJoZ16hN7fsuI3rSEZug4EIWVrZb1wL2l2/myjXyp
618DtxIGeG2YVZjz5JAHvqHzBl/yFYLavrtiGCQgMrHJM3G2KfKVZty/tNEVogko
Pqd03af5r8Ja8e609eLfWwP0tYGhBTgEVPJXnXsrjTeJ/xb0TQOHwf3iHWe6x/rd
uddVIc/NXQ+z7H/pNK39Jvl/wGSJvzu3CciSpzMvYjnaDbfzoyzOAYCHNVp4vwxz
I/AklYxnY1NZVPacFNh8k996fh1sBCswr4U9og0yO8ButKPb/IXzVjF6wD87zoBB
7T+X/u6kNhyMGjUxP+kL1K/8oCprbWCotBkpSxfU85/7NbanH6+T0Nz5kKOh7c95
VXA/bqVsDuphT431vm8vqc/AY6jBSI8QkzTReUhZVNItbOL2TBy/RTDTY2c17UH6
RU6jvzmr/9yD7bUEZPAPxcs0lMfhzBkqS/VPyNQF34PL55pAY1tJcszVhpVQ6U/I
NgpfIEJ2uu1D+Jc2tXnYjy82ixQglZXXfzpbrrXDoCkk75Nch3WC0vXMycBEyMyL
jDyfMvG7oYjRlLnqaPCC/OH7WP+/WjLzwL/y3qBBUU04xuSYH+Gc0SethJ91L8R9
cXUyk3mb4cs0dSe1yqk3nY6kg9MeYUcQscIWKEgeG/YwI2pX2BefcoKgePoDNofB
XFiU8GM9RlXLqh8a/PtCF0VEsZ1znA61QSdiEgDzna+4OFQv4qO0WGm/Obcgbvlg
cC8P4ybav09NuEJw9YvS2LqZQ3fpFaUX6bvvmXIwmSLrJY1SgKRBaiQbZaU2+cnE
9h+0cJr7RQtL8fBNEksxSkFwdAJ4tUVJ0U3v2JIdPLMCHJwETNn+QHaYOF4At1aC
gOSHClRmqu6My1Sl/EcccQHUcI4O9gxb7Nvu3dfac7QXdMiTbcvymFDkstjrcAMf
Atfe11Z3EcORKO6hDxBhdtl6KH+k42oZhgxaOiDIjrFxXKkDjWi3t1T0plJK7hAb
KIwA+9Glh6mWU93x8+NgdCvik0N3TYhL1ilHGrx8vWpxTtPKTSIlzfT9xce1A1u3
H1RDN4eRmGtP9v5/SjXi9PnY060zZQYVda0KkI5Qa90niI0ckAMGNsnhPSckUmr+
TDwYREU0NkfhOkPDXU9jCMQpyRBcc+7dO9vUclyRyo3TXWxFzcI1gD1Jw4so6zfg
7yrLhk+rlvRrSA5R3jD1uK0VBc4xNd/sijB9hvOfBmYYxREEaog8k5jzsKEcSXes
L/B+ikoGxCRmD2+7K/JZtBZ0onPG6b2MNvax/EmLtk6QY4YzgLHautJjBv9k7PQZ
9AmpM++WGZ0pKkDwXEBxYiUi3mBlroNDh8wenqYtSi70mbBApm0Re+knJfDfCPQj
OPOHPaNVWz7xrAwXCRx/E3ndk6ru40fP0XTaJFE00allZtgVh51hIP6ExSwLW/Cx
gkkkO+BwDtH9vL61HtzoQmLuLgYprVK7D8VraOoM5zAljyMi2aTwfngdey2/tbq8
tJPzjKk5ifGSsx26J7G6bUvF8aYRj7GZ1u9KbOb/XkNzh4av947DSjv5LacwdDVb
g4Ul25SVesBI+F+dOzaboXR8u3mupIMW0um8z6QAt81NC0qVn20mNXaQJHoK+zBu
pDfUuEmnU95FNPAmBg0RkFH3K1FP2L2lt8VFJ3zzmge4PrqppaGSdPej8eN0is/f
ORJO7pO95iSY7ltEMM2OPH3Xfsgc/qpCOWHMIAAbSqX4uXqwsy5SuhlI8H53SUGF
pSGrBIpFL8RT1nv1B36xF+dAlln5T/YpTzKwXKRg9GihZfJl8CGxW2MZXzlNNxWr
j2iChYoVSdL53/bvEAHFvbp77VrE7JvPIsyTwrisSKMhuud6RwrZSSLEHyApDtY1
R1Dc5R3dJ/3JCrB0Eedy0WKk5WVumu113qTTnMlEUJa4HvZGSQr03jMxp5X62zM4
/nzxfmbwJdRG4LshT1XPqdbBpZOwMSTrI6Y5DpzInlVZeHFuN+XUXctxuix3Ms5S
vI3qB2UgcuXf9jhCZgAIW7bl3X5maQw9dGnc2ONlPv8pW5Px0JVhxExfGwUYQy9A
xb2jySFbb6FjzMw/ukazD9M+oTwElbBxPoHYJWHpLoHOnFrgPcS94fRDjW3TYS5U
w7cl5fSlArlPP+EzJ9M6I1LPCAeiAfssxKvwO/cL4jATwZW/IpztpHYXSME+s5i7
8rXrcgGCIlbik2vT0di6e4wWPaN5HRb47lHCu1V6sEcuzHUQDYUvjoVnlkJV/qnb
R96pUuYEpoCLeIlccb2Bb8ew8uL5ijcnOqEY8N7GRPE9C27Ebvzvq5sYnCC8BwGX
lBVLcmA/bgm4UH/yQjuyCfd8JGnPC5HSUP0vKf6fknrbke+d3xAyDZCH/GEEL8Et
dz2TM9NkNpYtLQzTv9XLAUDSBd7WkgFcyGHF3MLRc053nIzBXBXgBqtsXCnCeRJi
J778MQ0s1R/wYEgkiQWDnDX5Fza3jgYr+/TKRg6XnuKe7qAT+1250BFEKKcN6cV4
zaR2R1vXk3a9WWLRqdNBDi+CMNNjaXW4w7P7QAAUbCgHeAJhgENZ6QICbctDJC3Z
CBVuFUAXn2QLdGnSblslqrn+GnZJCwYFGF9Mg35FeiblCkfqQcir8xNcRRgz2TqB
iEzHPQTv+ISpD6aGmTgkICYA0sEa6EAHkc7EyQYxmWyDw6Uvgn7dyaby/6IGmBMQ
vFWATrIp0KZDZfiitPFzNXN4N06ufzQdHW4r//fe6nMsEDdhBJ0zhcGHjSG/fQ6C
90cVyiXrIhVESXK4PYMLexDM3TpXf/ReduBqyr+zHZ/V5S1sN4FA+mpawwXRF5YE
A/usikXgByXa8I/GstExX3l97uGIY4jhFgDGK8FQP2/7b9uu4+w9h4EZWpRZsiHK
xNauTo6D4LhO0hLi7ASW6ipS6+YK6wyhk0HikFdcetQnqBa5gIBFW+WpWHTM6IBd
/IGKI6U9SBJvLCLxeD6pItzmcSgnVuZdju8EsCouhPJeCbgDjqzHjMN8CGrLe0ST
IEt+e0c3mfxHp3dreBKkITU7OrMjtIiiDa2cb6pSIPhum8zeW3AXbg097RBm30EN
TZbrG5pHkbWxsDKiOQVsC0z+FSpqtVzDb4wEwwCxpnscb8aApf0bcdYuQOIiwvOj
OrbgqvexmFEAR62OwdZ89ttyGpF9680LRUE9fOMV8HTb5Brg8JxyB/YFep3tfCkO
HAceQ7Kpl5u5Ar8SeZTFSEeeT916nrzLF3HjGS1rnXU8xd6Xn86cuBGmWJLZpEpg
PSbEhYNl98ehXbAmekYHCIhP40nckkaC/QAkxjDkrzdptGSejx4tI3anxqTFzltE
10xk6pxjVlii99NTre4bQLWwHk24yOLDJFDZ19Hh+3yws8/0Q4Wq4Cud7Xki9M5h
ZeplSsjdsPAxjxB8yrLECy4XBTVm2pLeO1kgA3IO4vjh0LNz59yTZvz3O5KRu1hs
TCm1mmUHXaUHw6lj4TxH0vUGqcDBgyRsHEIrHmam9QLILdC+ZbCvpgraDmE4pTR8
p4cQ9LbtbEn0UL76JrSBrEq8ovLGkorMouLYQD/A/W9bwoMyI/bNkZKYbu2rTS6f
pPy2GN4nz+FOgz9i142pKm7EIfiFjTNHQWG9xz6rDy2dyetejV40wHVlj5R/V5KF
x8oLSC493Kf9fAcmw3SqlQZ9/MWfxNOIMpk3DVhrbQHYSImOgl9nPwm1FyOilyq0
EP8HmgDyFWBwNww8zrcgNdXF2XZGqr+239eoCYUnjDiV7GMfYppC5VjJ5kN6W5dV
7SbXoNOOOgkN0xij2AiPz2Fvhr6wxLK8Y96wcz8BqBKpRYMxG8bXZkwol60Ty8HP
FFG1IDTa00sa6W6httttP2JfpV4l5OQI1hfzdPvWEvlmZ3v4aegW2HWVM6jsHHCE
/hKDWQctyKujbRQkyR4jZDGhILONu4A+qRkovrDxRCpHI7T7ShuC5K8i67vCo/TJ
v+Q0TXdxWn1AuCQCYVptEmm7jIph/Dnpn0hEmCVARk+nCJW5LhUxJJEsSwnxzxCU
/wI5+IgCeqfHR/Vs0wv9ruUJgC1afakrPLxDE3WnZPMIRdw0eovQPkksrJbk1abX
qsHwryVphkrMfMIHGA9CSVme09Tg+hPDvcZefo/MlTctRIP0P6L8KZvQ+9aXF4td
JmRlyBQwcpTOzcc7zADVJhF5ZNSqXQC5114NGji4BRSTRSkmYAEY3nO6F60vCunD
92yEMcztEKjPKOGXomlGvqWPlFZi6j1cpL7y4bBtqGxNySfPbyNeeuiQJPYbtX2R
uneAVQ2k/UI5XgOJj/wzaIAGyuE5IlmKk40hP4NFBKuObLS4d0DJ+9QbKZvUN7QB

//pragma protect end_data_block
//pragma protect digest_block
sjpVWeFJXmJinfm1bPMp9y+uDs0=
//pragma protect end_digest_block
//pragma protect end_protected

`endif
