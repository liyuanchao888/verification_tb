
`ifndef GUARD_SVT_AHB_SLAVE_CALLBACK_UVM_SV
`define GUARD_SVT_AHB_SLAVE_CALLBACK_UVM_SV

/**
  *  Slave callback class contains the callback methods called by the slave component.
  */
`ifdef SVT_VMM_TECHNOLOGY
class svt_ahb_slave_callback extends svt_xactor_callbacks;
`else
class svt_ahb_slave_callback extends svt_callback;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_ahb_slave_callback");
`endif

  //----------------------------------------------------------------------------
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
4yFQC9WyrRQh20WoTf2bypnDOhuX41UJxfHmhKdgbF3j148EQsrLWprUWZ3Jy5Xp
w78+fWY+u1bD1qRMxce6DBoEdL/lUNH1u582p40bM374jyYRy6R/fGRLLFZHzMt5
P89Jh3W9QunaHv8LiAV8BRorgl1lhupp9JQpQcJaJgfmLV7ClVlhmQ==
//pragma protect end_key_block
//pragma protect digest_block
KSdfCrZNkfBUifd4o86RDTGHVIM=
//pragma protect end_digest_block
//pragma protect data_block
N3r1jC0HaeaSDasHKe6qq9LsO+KFej2s0zuuChClxf4SWdem0iwc7Ek4vRSAyjHB
WzBN+FSnQR8nppK5gCT3V8stY8/FrdI2aXtvTZjISsDLn/+ntUkzEVkUsfZtgJIS
wazXV0tGp15YWbmEW2SeB9BfsWfqoNsaww85v2NZ+NfgAZjO2pIlaE/ZdhUyMXhl
jxyemWFaTdTveENosZKH9wsPwYM0hcG/vsuXKx00ffzzZUkHRBcmQZLxcFnSXwKY
4y22RLZBcBybSevieefz1Pw0+1I+DuK4bwqmEq57kX6W9liyO9reenegqzB+SJdw
8ouyXsuk+rDqcrJN19X+/vSlXZvwwbJvvwij7r0WtJuTxmYonERR6hhGcjR+4C5U
596nup/dbk6PEiFEVinZCJqmwSU/nxLIx1Knhg0D6DPbhPtTxVEheUojMYPwkvVP
HBAllBVSgd+c7Vuct+nDm78z2HIsMpTHWmHR+4qUJHkPj0b7nAbFKPXWUvZb9r4G
J7hBmBA2FEHfFU1Dwx5AzAvbRSu2SIBHEec4EZ2BuvpxRf+/3t1stvo5nuI32ZYk
Re8CFns3bx0uLiSk1mpaBnwNiPt613jvOlDfeem7+0B0JoDaI/9NCFejcmuIdfUO
814Z3Y/e3/dTX0njZlHXtwL7wJnan906kmryp347/Xw/2s9NajueBtKJMM7S0fGa
5Vh4TWCLHkwC6wronVnoxwsNlkLrJjLefa9gpQoSywpIF6EbsJBOQ4sL7iooioRT
RKtx7SaYBAh8Vt3LM+d0XGh52HMPfCUdraiqrWLlrZLPGSHg5pgeM8bjpFyIbv3h
C/p/RmGouZSGnvY2dtFG3vKxI0g4tCyWjBCI+CI2GcgJWRD1WV+x2RAQqs8HQM9m
N7aC3jm3THLe3ffof7CX641j0bXftcRA7o2MchKNgMAlTQ3Qor8kXKU7tuiOnLBD
pVG/BY/VWq9L02NAQISSOfgBIW2Xf5+q8IZOvxi1cxl60eqX4RxXjkRH1XVcao+7
M5IdSCcOaj0CizxZNljckNj9RAfDFyPqnimtl5BXrlpPOkTxDK9vw0f8st77gWqL
8IeaxzpF/0+0D+btZ1xSTTlJvK3d9bDrShnciteuFogEiqDIdPeb03zpJi0+ng7b
PCFsOhlxpmueuifhoBEpVShexewoKCdX0T0djaai0RwZkB1hIGQeN1MC4MzdFgWv
2jfgayLXahgjsXn1cdcespbDVCQQQfGhIMSrNX2jwsjr3XXcUFD31toCelcEnqm1
KNa+Xlq5Pfzd9dtUdiXlEf/OafPw7+h2AY45q77JKBw7k0BvFJT/DxIGeD9vV5kX
GZnYusLwhps3VE/RPuGJ1y7zbl1m17/Smqs34RoevAB6CXxShNgcjLrhhXQBoqPf
NhwA6wmTUQmD4iBZjVJuGDI8tSg9mPjjRDkqodXmBcPxOl2PZ1rR978xuVeYliI3
Mj0IwkLRpB8s1KvuKD2DLGL+ZAjR6JK6hvKxrzTj8H0J/PMu+yT3jtEzy8q/jmd+
yYAc1WP/6JhT4jwdDwhiBSsr1EYcCM3jWjvBN2bPEd6RxD8SgqxU3tYJMQXw9Qch
Okb4rXETL0Q2spZwW5+NN4Tg3RsB0k/PjEHbBaSsXDGyeXYbfJjp1AOtgIkp5w4j
E1ECReI6nuWz5Q5SpmCFHA1hZ+Ymk/Ix9qOujYpHAcS8Gx3AwRLAlYJkzBKGMtRu
4kABDEvwGaGjpcmUNci9S5IIDPbTHuKeRwNHi5CJiggih1G2i7o7iijyA/mzpnKu
L4DL96NsA7nmDk8IGlieELQDBS26iEY39zju88ykDMzn0WJz3Z5no7UND0hPpJtP
akoVI5BgzpOHkb4LUWDVnVEbNaoi+mNYKEzC6Ndz1MNdCMWETF0VrwV1SJN+SGIp
YfuV2PSN4nA3KXJGh4MWx7DS3G33Snyor0cfyrj+Su6csdpOaMUYiGzNGoS4WjZs
d4O2ZW3GXN7btZSF1UnPIgLlGSEUmzMhGwlUmpGBmn/+/QPfxMOSw9F9F972IOWF
V9Y1SoOVjrxmSYoc1Sj62iOr5fSU1lBC1Ie6mB1Q8TjtTSo73E6dfx1bHjUgdnE8
0R4lKFG2l/ajzgHI67plpZrUJZABtOfmwf/BtxLlKegrJckjHTXCH7f078xZRIbD
FhG5WGigyH1Yh66yI0sykye1lIpt9Oi+qSxt5U2/v743sczqjLrBOlPsDLD1oN2e
GXCBIVoV54Ek895f9fWHzGVWTe15dhWv9gotJ1nIccagBLcX7JdUkpsAn4Y4Xb1v
pQ2MgShrtXlo5jj0op0OURDU+GMEPb3U+teD16LUPDHCDrID2w5yI271NtO/dRTI
Qps6sKsAdeT1KvTGlveesWFio8PaJkDEaB7QfCIAG4xU6kflw5PCCqQDnSKM7RhK
sFeiFKnWhsQZ4v/ynaiNEG7ZtGlSWb4XfkogsJz9NfgkeayFHpROBjbPHXcoBgjv
UM0Z2ipSRexqGxVb5GpP7iBOG85OdLkS9G2NhrFH3qvuStpdM2D8oGHAY5v18H32
tIBZh0U3OZcxZzSCUY9fxg==
//pragma protect end_data_block
//pragma protect digest_block
CAIvXnC87cBJw/kC74cViuUFSKk=
//pragma protect end_digest_block
//pragma protect end_protected
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
h/anozODbV1mVdYxivTvLkhW6k4EVSoccXYROcoGcEOiKxmbPWXig2IwAKsqDUKX
FHo032uz7FWfAN67REYN02LgjAVhr4AEGHhmQDTFQL0XwF1FTrVCMhKyZijHOydT
rFTVDGCXxaVEZbUYxCfthFUtW0V04yQbObSNUKgmCyj0fm/n2wnX3w==
//pragma protect end_key_block
//pragma protect digest_block
wOAbelkXeMto2XIkJVuaIHlHMNo=
//pragma protect end_digest_block
//pragma protect data_block
DJYR5ZPRjJfqMD9kEty+y8Nani2x5cDSpFq+6xS+JX4TrixTSruPp9Em1y10LWv6
xExO/MC/oDD0wLOLIz+iLrWjQO/YJPIvkMvjgVrWzU3Q8Cv7ydwKMTzoSLkMuHP5
dHSWqbwk1R3yEah80Efvfi18OoyC5abGLx7ZNnSiTTKDEsPfso3nKJp2kDKBXoAo
R1mE9t2td01UwtDQGrb3SwhJ6zxogeMCK94oZe9fOxJZk+8jq0SrA4/y4fKFnWkz
oCHPD8P0PSVkwdrmXm42OwhsqnHMOVHsc1078x+mdk3+2BINWO+/cnq3MION4404
3bN14fa4Ug1EZc/AZZeh4JCprbdpvj8OvcheBP6F3J2UMiDibQjsp1gjHXwboy0P
mrcfWKcd6C4yoY0j5gusGhkf1xHjp1/ST3wmEbiMQJcHyMxv0nvraUb5vwrDds78
DolOOQdGQWV3Tigg6vb97HwVuEIeo073+Kj1zBVd2y9k28IVgMVIvpLhy8kmFOCD
l8wUdgq13Cku4PZ7sVVFMwBn7RH4+66caKMJq8//ES7j9puVvQV+GXLv+JZe5cWM
GyMiTrXL+L84LM0cG27YqxF9FPOioXvQLlZ9PxnnztjaV7DrhBO3lRIMPUTquWaY
p/StHoT1DnmtUtzCpbuMcJNOigadGpvowfdgh7hlfbvT46+eW/MD6kl68VtzmAt8
Z089RVz7xpO1TpUn01NvfQ==
//pragma protect end_data_block
//pragma protect digest_block
WtSKG1YI0yKPSIP0g3OdIQDec50=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_SLAVE_CALLBACK_UVM_SV
