
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
FqB/LMQOmtHI40Uuye/b29DZ4Xh+955q94BFNIoRa3q/TZImk+/AwECPH072V8FM
DYa//Xbi08uglTOOnehfOfrKnsFM9yULh4sudkXV94CdC3W66Te3/1+6aedsKocU
YUPPYrvpa8+qkww1JXE/fNaIF5TPPMoAYlIoBsV0QOCDM/SBaGU8xA==
//pragma protect end_key_block
//pragma protect digest_block
IhVC0u/FBB2zuug31aADREmFL5E=
//pragma protect end_digest_block
//pragma protect data_block
8GgxI58hZKOkPnofQ05o973weXEdCqkjraZMihmKX7zRJzCMqhCHC5xLyui/ydJ5
0QhFfrUeopylLwgxdYVieGRuDn0dZhM8urhM2c110N7mBDp7GWrNI21RevysGUCw
ZNh1wfLd8y+dq/yNE6zAljiTrAKaSmunc8jpX7NHeuKG+c2cB/4aZXXlsuGj4D7E
VKVODlEbQmVIrmsbBCt08SjdA1Xm3QxmXtMBdxeLkPWRDFz7TlLFD4Ji9vtJXZRj
t8He/8gKg5/gSX2CqXVeth0oUcEVcrU+5DZks2CQ8aq18omw7bTDenjOe8TV0qfs
krmesaJjPj960LEh7P7eoZb60BqHBTGwy1Iu9S0oRAM8BeKSs8tom6DuYQF0OxOS
eiysY1BydARQhm1LQVYCa3Njibuap4WNMYTP1ZqZIVI=
//pragma protect end_data_block
//pragma protect digest_block
S3PBzbCzEHRAViBLus/luwjRh7s=
//pragma protect end_digest_block
//pragma protect end_protected
`include "svt_axi_defines.svi"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
7DVoNxiuQF+JjaEUoAyvUgIM2p+amj+lxM9oKnaPof3o0Oz8QzZHdA1lsgVMnFLO
WLN3Z5OUZybmrddffLxq06CI89+b7JAHcpUA9NEXTGohDHrfNY/kH/aEcC6mKpT6
c2BK6IOuHWzXJW8jCVCMqj42y3gNM5g+Fcx3OBvjnwpCSdkwY6VPEQ==
//pragma protect end_key_block
//pragma protect digest_block
0iYIg9KOZ5H5WkH8v2nxgJhmrUQ=
//pragma protect end_digest_block
//pragma protect data_block
Yje1F7Ah+cqUty9tY/seO17ue1762dQeQjZFvoLjkiDDNgZ8ARZvxc60sVinlo8R
Uk1ZFsVUwVHzETs17HNUn4qvHsQNFSqZhchTmcuZaFrY4TXG9euWxJPyULPKmNOa
y1H7y3MkayD0p/5NiZR/jpP00OXH52lnFro/oqtAxKpLg8gFxidOodwE6ATB3Ci/
NkXM1g0bqMVoPMdZKfkMdCQE2zHRtmROtBLGNXbCs217RRStUjXCZ4WG+8zLxAkk
sq3Oh9WAS7JDzPOaELRQyUHH+ZjBgteVMIndIUit1G9kIlSI3UGFaQ83zXjTjf5/
sSpKDN/bEfypJmT5pBDty7b/jjX0nG3hTgwj2s9Pj1QH3I0rk8Q4IE+VlRuykcA5
wLPX4qV9jErepzvoiQ3pGoEDsE9xONqZTj3d3zsLOMfdHwCfWlbCtEkaXtlJDW99
Fc4QDPttbMHlgsbOAGsjhNzPVJ2Xs3vOcoXVObX8UabZvZH8qhkGQsFpYTCKAveE
NSQ00NRFkxVFPjYRotRLumuRMHhL0MN0KeY1SXGZ3Fk2ndOw65GE/jjqQmYV5Qxd
LIqFtkz2BhY0hUwsHg931gS/1sMdiSpyP2bhfp/G5+5DM4UqLYLsOQ7N8ALtbNP+
Z6leqQ1TO3dJfJzBDPSefXQc/218B6t8hgQvJyWtBIv2Y9vxbmtd3TVoWzuBZN60
2ay0DS62key2TAAOJMCK/5GpoNBZKkUR/UYFEksVqvj/LcFSKxqO7k79r4zmN+hQ
RTTlVj2bdkHaU2LqWvsx1YPDUNvpQOI+V2yCeQuwSWQGUdoZt29JmwgBl70VLCP9
OjFPPEsUDEq8u09DvmV1jG9QITR5HJ8vjcM52GNh9WRwYuv9Y1a/8rdQyDSOS2yh
cMqiYJp64YzBKmNsqL2MVhxygUiTNTP+E09ncf9uIn600Iw2zLIbVL78gofgrkhg
UF+M3XuSP99vF70wZCiESfx8Lwzd1korbLz5kwU85rUdn3NrlfI1cu927uzpAB6A
GVW5jjaSZeGR+UCaOVk0rn860Yu/o5vWCpaCCWywe4rTMV7fMNuFDy75f43v0XCN
rWbDT5iBeb9QtrCzULGfBx1jOvl1sMvH8f0gPN/kCwSE1ni+zB/KQKzaJQUQmJln
DlfYCM2mVLDYd+O0O/5NuJH/l6NYr8Xqd3vzoVFfVgz9Y6IbRi0j7N8EnqwWXNga
7jI0HarwefNaq1xLj7SZiNPZW2oSz5ZAfkgCuG/Pcxf6aprw64JIGH7+X+GKg/pB
Pfpxz7Ev7bk7Mf7XPPeMwr9o+/A3eeq9LPgNA+CnLG2nBQm3+zcruE2p7nFodmrr
yDg0/UHykJKhNejqVFmY/dYw68CinDc1uluuVaBu/m0FOM6rQ73wKKn8mbLvCxCj
olfr5uXhKbqXBYcUF2QWnUJEOFbe3i9ATCs5/HI1MnaBcn6Nf0EFN+StxabpZzxE
QSDwz0/B2/AKJONjRJ1j5rOzKSaK8P4SQW4yrRTaQ6fFuvfsMS974tztXUj1jQ7z
BJd3DPVFrXVjdXHfGgJnI//jc70MGVASfyV6CwAh3DBsU5IEOtzZcLVW+VoUQdff
coiW2R1LLVyIt8eX6Od4RtWJ7Hy9zcbhbd3rohwy4l4sdpuI4mrKjryYaQup+zJo
DW96x4vt/iaFZsAmdXFV8SGTK7jkQCOXoE6CsvLlod1AHrBjiMRos40DVb4+eLXJ
v37Gn5nqy+FQNWBXgjPLiLTsHRBIGY8Bsx4MirM0CfzrrbT/e30KakfnN5ai38B0
Bc/z444Lhab2AC70cfyeobxwWEpBP9yGP6lAA5iAuKCekH4lfekDk4/uW30Y7n+n
evmjPMU0pG0F2IGVmBivpl+dCw2pVw4Zpy+caDxlY15t60qm+9GtPlm1MO9naqwL
oRA3IdOYIUqxwpAYqcw98/RntNINFlbCXuWnSHoVNMByWF8a/FaiYX1QWBaSL4M9
tn7HvY3CqX05MVzaQxmBiZcsV92JDPtYYTaqxrnxweldSr5lOFc2uTPB8Y0oi1OM
PytkRfCTl0oxUNS+g25KATTKnySH+DANg5+0bg47CZL04hPXei2mJrx5sWlFjYw1
g6SAmPBtJQzR5aVTnAsyzXBsluf1YhewuFuYqMnt9iS0fVY6HU/Rbg7S3DiJMpJ8
0oAs8c3NwIDHBzopobNN7bnZOhTMKbvG7fmobk62XXFYznKBYjw6flmCemK9TpY4
GYZ22rroJEXZKUGEBxpDoDJ9s9UxmgVKGwiKYwy91VLJBBxJRAmE5txIJJbM3lG8
A2X3o9gKQONF10JUXKHhOfqblV2h3EFO3F3jxJTXpist7Swg1na+8w3AwoTHz+7e
zUhx5dxA/HbTYnM6d1W/mkDgQjwlr2Yy3BxiV6nJe9PLTtJh+tpJBFOPP9zZ3h42
+ubLpHeYyrOpv3Z8w0psmJ1WP60+1jgSssuJt69cFFzX2xBXlaCfz9yKm1nB2hu3
++/EIh/+DT68ucby9+W+Zu+RlkS+hLsa2Zlbm4WSUGSAUHkf1SalVlmNI2kD0EJ8
3KXUXBGW5m4xwrE1SKhSgFTd/0r9Fx45CeJeQWGnbXEVBqUqnJ6/Ljb9d8SISRk9
bndJ3ZlYCAPMcvF9tNebEz1k9pzopWiqPczVg2zp63KvR6v7XQYhJHSCsyR26uTF
WFif519zJG5YXxGfplIkdSeFkkAZOfwmW0wId3NswLygyFXIqRITySK0lF0jnRwR
PEKzpiW8zdJPejwlGKr0Xh9TI1CC+YLDtAmFmHnX6exPzuKt/AJy5dnPaq0m7Ccp
P1ASniLtXm4cOjdeUiQz79aYyu7vmlhl3Cc0nRu3J4GnLFcaPd3mbt6qoc1jF2H3
JOOr78F5pc2q3lZ5hAZUCOAHKgkJdUvHJnm2ZoPS+2PZnTUb4e63qL4MPqu2w20Z
TCgJF9FlsDcQ6RfI7KXqCvalXqp0BzxXgl+z8pbFiSADgYjJtehbHwsAxacwPjHs
q37RHBRLX8sQIJRkby5C3eIRJ3IjZc0gijKu3XcSYzd7rjkrrBRHc/shuRLmEThM
dYcITlliM7QxAwe8NN3MQdHrIDdphaXEo05rAXR4utYbFYn64AsbB2wwghaHJTHR
4kjLEPGdNTGMzeX6dVaNC3Ig0VI0bG2XxeTYpLbi3+6IUJPGeslyBRdnSfFXDuPU
Xa42pc2vr8cRhh0vo36d8v77xAkEfA1bExou0ASoE2weQL0zMPi+QiTP6+6S7zcJ
e0kqaHwXVzie6H0Q9M2Fghwmn3C3nOqMz9tC3n6lB/Spb3sub7etTozlFhhEpCdK
RMCzCtAmgaqStUmIbDKdhLrPJa06tZxZPz0CkPN9f30C17iAOimhnvw43vLhJdlw
hpKvH7M3xY8BNDGW3JJfjaJDN+AJingV08KewDOApaBRs7Afq2PPT4aqzI9O0vbg
R2zsB1F+LKgoMEWkdZdfdQ2VdxBtKmk769p77PQfcJKCwQ1Ysj4MKSEPg1VaMYG2
u7Ou5kdnOjORm7DGJ1Et5dWyUwqVp+bJB687A3DpCQxEED0PiKT9D7t8lRDEIlxY
7ZQ7MY8/W2/ITc/87mmQUaDd+gTF7gtC4IQUwG0qEyw7nPcxJY7zU5G16yqq5nnf
GpVDWvYBlc3qVyaKi2jcf7TKsDZ3lqjx8W4usAhuF1ZmWKb955XFH4eUal7sjehl
M6NXv68GKhLgVWfEGlhGD9xhhoEDPccLuKYL8sMrIsr5bfBi0ppJ2dxxQO2Ntk9n
/WpctSpu0UKhq0neDWq5IsdJ5/fh0VJxFWXtEz8xJHgRnLTqqmNWpkJeXR+53RvW
mJXMXCY+JtNAyi8+1CgKueozroB3HAgofAkIaewYsSyG9U+sFKF+8ps0ALmUgoyT
sb+SH2pxhCbEKuIC2xfERIz17wmWbrWQEirDfvrmVDjbET1bFnMPpx+3a5xBB/+V
YFIzYhysRlpKTsgJWujsNasnwANd2u4jF14w9xK+BqygyUh8pcJX1DDfRSsZBD5/
HvB/D7tTwKTlH/CcfyFHzZ1vsuiJzikJYMsWTaJ8/U6vBAB7udLNqy/2h4RbPZZY
72pTdPef08gEd0hMGSyu2glJ6isdrwYDrxZQRUbFgjahsBk6vXL0VATwEd5ndugI
wgTlKecLPlJgemvvy2v7j8xqOkhljQlLqD3wBp2YGBJjJL0L+6Cg2SixRfJ4emE8
gn+jo+mtbMMkng7koBPYoMyVKz4/7ia0emcI7qZMcANJLsZ7scH/IlDDuf+sYQ20
LHilVgdQf7PONnI0iQk0q67RSmPlUxxoQq/YAZgpfB+Z6lmZFzRXdV8BLqMdOpdq
wgdsFRtR3kvOrMqyg8RntxMbFbDSBf/HdpHLztW0iYgsoTf2ywsS7HdpC4VbIX8l
jpI7Tovb1ug103rsfoEL6dfQdETflrcLJYLfXmMf7WU3EAn+rGeo8w7Nw/modbFV
KTi/ODNn6NqPYCjmTPnkroi9U/xDd/U/KadvLco9herUfC3c9fFOK8ZCH9F/7KKM
0FahoVrqEYVZw0PgRig2imcK+zWhOt4fgfb3tIGmbXacvhsrkMIMrSAnhQ/rHwgh
OMIsac4I/cO4h9N98CLwS/pegMAyyPHrnq7630PgJFswsLbnEBrQAQOFgupqIh2s
2O76cyvIw0ygJqFYK2z/2ymM4aMH3Oi6BePJZbg8QNtSueeBh7AlvbNaD9oJBqVJ
l+96NeU+tH7qcDIgVGna/VJwy+X5JwaQguOzVzPFoMLJtyELgE6mTbkXm2eWCrC7
ppKhz1ldrC7YmZLCYy3Neg86Omfd+b7JjIBR6VoekqUaDH3Emtkw1PNZLBMZjnit
qcdP6cG8VjJfm2Mg8GzojmXSU0Ytk3LnlQ+n/y8UyWB26HFGVlJKvf31U9a0i+MI
zLSi3GslvG68fMKyHIPL4gxXzhP8TkHN4nvVAIZla74oIQb1Zo1mCyEIdL3sgoC/
tCq27+HxEHAR/VV3q31s47efFiJTRrEozy73VXtZHko43w9qLEXPyQUPVtc4MFcA
ZusXfxzB6N1n0C9r+OgybZHMy8v0zLpFGgFYJb/3VJfZP49924Vbat4j7lCeydoN
21P53J/ja0WSB61416AfHyFLYZduaiX852XcTBECsmkQ/rEbyTllhBU5xZSERQmq
JP5u+gPgEQUmQdeIVy5apgbWX+Nni8bfijwC3oh5Un4mV2j5Dk+oSuQoy5cK2yzj
rzya8pbadqVdQl+DM0I6hUYBGgPgNdlCPOfQuPKpKDPWMCXQ9v1KmQiBomaffEGE
/l5Y0IqjUxorhFRBFOu/O83djUs20bofThortTmQ/TCim2PQw6Z6pODDl0HVZakx
CpN5kxq3lpMRM+qGFKXwGqplMb7WZLjCwloqC4qAKEPHMxZfj8RGne1UpToSNzdK
YtAy5M+EDSaKDomm4I1fS2EPgXWvnaYVtgWnpGQ7FNfocKEFTjuawG4NU+t/xwsM
cX6/P1Xn1JDeRnya4v6pErO69U0zsCSC4LsBiR4VkQMkUVVN3/gCQkMZ7kNdmDs6
Xv8sQ3te/5mI75uFV8wbnyk4MhT6ZH7x5XsfbwKNQkH83ozLXqsQDF0R6tKIhy1U
4k4nZAffVLXd07QOoFGyS/imrjqNk3Rcg1GzKfwOrQ+Kv+ZhszZO4aPoWRhr6L4z
aj/tM/Es5Sh32rDGkCcR6vqCmywBhuAdpny32rIqZxFO1fozPq+BnfZrrvcFvWRZ
RU7ijjeygC0n69dzAKh6AAnvOWb05oZTjWTyHcWZYK7k7RbQWCmOzFjwWMuhEmb+
ePhYihtryV8EZY+aaNkh5oJJFAqrwFWWB7ENvCOpy2NoLY0qY52Xve91PjrlssuC
SButmIlKxiUIZKOTRrOiu3P3sBlOf7ND78VVyP+ShyuQYo+HsFcTdmaMzkM+zDJ4
2Znl+cFzegDAkBcPuLspPRgycqYNaor5dLqEITJUcT1RDGQ3mjzqosDEp4BW+Dgb
FuNJIBiZyXEU7yUZk2ju40VtuqsOh+VJlJ297UDalKdEUAXy0zk0WEntLWiOWtuj
mjR1d6kLkTGFMGi0wKRHaQ/WDqRpsDbF8z5pDRWbA3YKXfsNfcKGC6cqTQpbAbBC
5y3hMz6R8B2Scpsdn7GtYQIzdN+P/kJyl9D7pSZuchQj+WSXGALP8rWhpe9UM1Mj
1N2gzKoOkcCQSeOUXxt3leMpB9wIB6a/C+j82ZHwXDTjC9ryskih2CSvOkFGS/H1
rGYD+2tR/Xu+t3CZyyu3/8AAf8DbmqgUiD6zWCwmJ/T2XYjY1JQm/4CNz4wDUjFw
F74NmnQrkE+QcPqdanAnDWLl/iKXoc+4cVKPuJ1EipxBYyxMkpjdUzNMcKskDLbK
OVbXH6kyYZvuiB4Fb63vl33odn8bSLTgRYAfqcP76kkKaBR1zi2zSYFr+cqTD93T
cXwewXXsPp/7gXVCPFD2LELt4QxENypVko7jFMVO2+JGCtnf2J+X7XU/Q2X4eGSq
4Ja84JYafq1wdzkSbNFhblTdSWWnQ6F4E9flLPiE+TgAEEw3qtk2WAZYGjh7QQim
RpI+nZr1qQEUqcGkdTnSaglkiKgNtSugX8U7acuuOTgzlMrqes+I4b8m/DV2+Poy
+4Q+GWqIDBbzXmq1qfY7SwwWQANmzPVkFv8K+EcyQGikBJMhwetsyV1v5x5LvAUn
msqNOMJKV30pEgUEAOYSUAa/FdWeva4GAqbYToEHtW1qnOButC+Y7DecUP5LpvnR
A16YY4C9cgWVUsoGb/bDIE4tsz+kapsAIYAedv1Sl4eGbXyXhtXGt8gL9AGyzQy4
cu7erMS0fJvqYv+QFXoBIHZ6nW4ZymRM3xTmwL5Wvqh0VryyRNVlfsvOANqOdA8V
s6hklOxsStV1LiuyEJuzSL+tO4raNk5Fba0FNkWAh3+rOQiMxDShcWSbpMn7Tfpi
9sWPhYUk+CQGbENKmoVosZXb1BEpaLxH+3yJrfszSZqGdwnG/x8tCfGLHxa53rTu
6bGpLN3GHmLymLfuqipZrGFvyiD7gLHix5teGpq41fcKw0Q/tu07NuhD8ZjBFOh0
bQ/ZwvuWb278hOdjhe44OMupclcO372oy/wvV0YkbKSVhITKiGYjQ/DrtPcbKE6L
ziDuJ8mlpnq05NNYUbmXa/G1pFdMozz4Wq5Kri/rGQTQwvKheXc3V/yQekIdAsW6
jjASjnv4Kl9Nb0O4M9j3+KJfPsRIy9YfxWxIEXpGNLfQRmBh7fNpBZ8r6rmsS8ep
uQhetnewkNBaVpw2TQP5LzqmrNvzxNRXC8REUjRTpKg3hb6FZ1CHg5cx8+97JaUA
GMoJLrlN28PwjR84mQXE0+bWcN+URuGG7jGA/FOLpesPtKQ/QyIWeWNrTxxG3okP
eCyPQXvRT0pne4FuHe+708ONYwUTsaVyrtBDKxF+NBvbRZ1tnmRdAgrUC7q9X3t1
glgYTQ3cWTjNc0Tl5UuoKUS7bgvs79lMxI0vYzXkTBfCBvm084lLL4tSUZ3aGEJq
DEOb+vOfz53XFn2S+vrzJhb1ojKpqfVkkLac7RpjBImn+ZZ1iYZlWBNY0pSkzh3x
cQEvVrznzaT5aKzoMppN6xnclWwnfuMOY+zLKGpgijIVXPHcRrDrKAL3ZC+q+MYj
JCHB745VPXh14vBNvmexZJVMiLcSZh5b6xtEM6/e66dkQ8BFBfQtlaM8V9Uf94Mi
fygtN2sL2mIOW2kmPFn/Mb8uO/mSxarw3IlCu7X6O6wMKP12sWPhiDpauoM0Tims
9JnUCuoaro0Se49NmET9t47fk03JnpFIRWPr6v212kZJs1KE6gDljPsuXg5K15gX
yei2FFDp/hVuwKsG5g55J4A2LuExUjcwRjauQ1MHlNbQKLlI4sZRMtVtZYm76k7r
VYdfKahUY7+lpaSZ/9+OEDN50HYquZ/sz1AHWmD1oUR+rbjDi+zl0jF5gt7zblcB
+zLDOE6oWM/t0VZ03dAfhsFEqVtCdoBPt2L5fS9U9Ngy9nN6a/R3T1ozPutNc985
bbnYVBFAKcnW/9ADjYazdc0isDaSoeFMB9vr/zqS1ra7qOOIJK4s2ValaKm+7wjb
7e0BBiqGcVdlvkIydfhc4HTkZxq5dKUJt9z+3xGm0rjGsKcdHEsBQyzLeCoi6+Yg
WmbsjLtU11TitBy0Ot+BrgZuSoi4b0ws2/CcaM1tSbSNCLhCj8PQheBJnTA4bVke
LWtdJdoWJjcBEh3XMcf7KEiYuAYRtjuGqVW/Nau9Q6sn8XJqBEoN6HpEYc+jdRzZ
SarC17S0APoAiRf3ETTuEimyke3xncal1RSKsI3sEOkSbMsvurS3dQCUoTO/K9HN
Ke8lncKbENymy/cNSnY3MFUC5KxQQe+0lu9tZkXoWHrDQ4LLY60+9f+XnPPEGenn
dyUAkH40D4M8xUDKp0BgQZz+28K40dnQXmsA26FlRpBIT6uxMEY35NwQEIKKp0Sa
vYOSOaqarQduqkX7xCCbtr+Mk1aD4MHP7vRV5ifHdLnj7+Fd06EXbwfMrXlcqIUT
cqH5T0nmkAdJDkupvZkKNi7OTPlCoBavGiA0+n3MCX4hJfX8GGpQ8eNZNKi+r7LR
Sk3w+1UQO9HedMRnZJTc60UYixxCx8P+n6jn++AzRtFpGHbqh+dkpFUmublBacUs
qwyV4arseeqDamk+y6Ot94ipBqKohtlXOs2ads+h1Lb3Gsp2XOwAFUGfcG7m8E3L
MNHSXHwUfymsPk8Lthdt89Dsk+DYCb0hql/TYdbLP+iG3XjJ/HFRjD37r7FOHZjd
Ds4/VeKzbHYKlu2X+hMQ7Oifsgmvbk+Y7fqe6PQljGmcN5y4cldQGzDyb+X2C0Ck
SQXO0OzYFpNgo3JK3WBFzhTIdXCU+4nvsAxBt9EXe1JhfIBWpKb6aofN38xJ0rjG
C9RDXASJDvAiVyilOHm5tPLqJePy5XO47nOxACGOJy4MIXZz5wo1xJaZK+hX4UxY
mT1wxmg2qvXjj0UNjgO9aKE6SMbm8oQK66hY9NIKyABL01nKg9uh7I0jN3HJHEhg
C2WFZdeVvQr/Ddoy7Fhjq+FpO4+kW3VEXcbVh6mp6BhcRHZcKua+Ejlae6MNsQpS
LtowsdL9U7gHcTSUKLl9k0ZXHiqqLHecx3OdY2J0WmdP9fC1jl/VahJBUQ8+9xpY
v55hQZDQTsVFa9BIKm8G4IOFuF+ikI0Fg0UE7s3j0IKAqNPCCO8yyjVqrh2soM+F
mgcURLeCgHWD6CSu0aICZQMZqQ0AIqhJsjCIysYy77ZdyUaAoqkdGRJ2ItXvVUWA
BojTcgN8S41cAysbKCBJOg/szHUkD8cSHxrzjRCCa2lY2LsO9uDz/kKVgzeeBxYy
ug9iOfEBYL/DwDWuHmxtoJmtTW6VE2XbVqp6JxccnYA09LRsGA9zUhbv+aVEIk82
dekjxDrk02um3DCW2HruH7peo1nQ4/B+uMSny63+h47bq1FGBt9NZ3kGu6aZJBuu
2kx/5dCJKc25fRMJmfuST1xANio6I2U0Eao4/vdBFFHygzOzwZxGtoH5RGOBGmCJ
f6P7QIHKqLSaqTbDrUcyqUDCfsrld6jwewgAEwP5k9Ch2tOuFcwh0PQ9WQBGt9rI
Wd7w0CKtGiXntbGKgEIYI6LGY45zfZBiCMYfiR1HkC7b6pvbyPvPN3zXuEiKTCQ4
2VWcNFW/8JC4C1LGlxwWme9TBRFT3evt2BAQ64NR7o2TO+uoWXQPrtbiPXTSxYKQ
VPzIHTHIO+UmR/TUlgr6G+FlfW5pLwDCTmrxttpDeqvkYr2ECR/k7wwLCHvXrY8f
mRNc2YZyXPych2lRav6k1FepQSFCIlj1vmpuBvjDy49xh0EtW9Gxb0sz+Tv77dCY
frniwKkGZ6UMYk/eiBhzd9M0mBKFReZ+vuGryHBAHnXDDBJNdES8HUSYPoanHAyn
0mOnRFHdxEWqzY9SLaA7KmfsRSvbBgY6uxQ3AgWnHaKiyjcE9amTkKU/McBUBg7G
bjFo3UPbjpjqYx330twOoHoFXy9gvaD9gloAzHSYD5hHMHV8GwxTarNWVBbzsMjJ
7n02ofC7VgR4Iq8j7PMz+N76Kuvnj0yia5R+hEAyJyRwRgzTuWYXRZcDQuXoiF2u
kEPEEItA0B10b3Angs4mhmSnIbZ5WLVGM/egzPB6w/bojNEtgfjJf+4IyobIzs/9
su2iHUZ532skICSu89gZNUM5BKLaQFfU/lbUakvOyiEtqk28ZhNQq+qBzGui/UdG
en8OStB4bCMkTujggNcVIQ2sxE4uP2+Ec3ABfVP6IDWmy4qjGo2ZQ/Z81PLPIoJ4
2VUwsGXJtAWncprhxZAsVUt2mz6I5dVM3E96XIW93ZAC/jCPVaAnK6DTIdHmhje1
j0Scjpv1gXHWwtbZwRJ1L9qLJk55xFMTFpvYL2BuE696tcXLcBs3leEyDeMQe5BF
dy6EaZ1z8iPqcNnKXKIY664BrTMJjFVJ7FbkXX5cN456j084QXIN75xfIqBnPPPJ
LH0QIxHXZRRC9bht6Ef0wPYz3WTSNU3mjoHXLqOhjONwu3X6Hk+gmsqKgfJJQejc
u4ag1o/a391rU8sbB6sfZyl1U2Ex/Z/yzyb4RUgmSUatDjlO8wHgYNcPRjzRew7a
CHZHdA950CKzANuQKdw1jliWcQxfM1VjgNCGjXi0fSw1EufRYvYaC0Jefi4SC035
OtDbdSHx/+507hAhWGaD4bHDtadcmZXVjTm5df2jDdc4jcNrfeFZa/xo4q3VAxvK
V6AbjfR2S3LH4qe/YTQX9liUGJlJV8JBs8L6evJws81mn4Ffiop65p3M1IbqvYnG
wXJHAxZswE34zFeZedWcSDJ8hLtl5iwOdZYGWXgghrfqLCu6Byqh21Z5gaByh5DF
K5NY/kxSbzmbH9caq0O0Sg5BlHNITS6ZmV0oJ0Yl7mn/5hbtL4LIDu7njh5hwcjN
cEKHutYrnBB26q2qRUd77X7GkN1WDuCzb8lX0IqldxM5tvdKRwwl0cMUOZlF+G2h
QdxbXakhWIbJKK5cP7oLDaKBkTjgLvVogY935uxBatuhfV3zKYLySz+G5+KaNC+g
m3Q60JOSPip/SGBlQxtirPgW0nREe41pefLMJv7Vq7Kdj++l1he0O8RJU0ZcT/Vn
lWa7fIKLG0verMfATRUcNPmhbTac0axccqGjQbVJKXFDL/tGk4m1F+NhSV578Ctw
yvhrjyo0NEo7naAGnKudoKPCYvfQuiYciuwcKRL6EhUdDQO9tHH5T165Oq/aKufJ
/oqgExkju5tfNwAcgJ3MpyyY7jUvRN4koERM60qUf3cbpmft+zApRev0D/c+n9lv
MfOQ3YmW3rPR9lTRB7+HdvLQlXbJeefHy6feXXpoxODr8+wOs8w52gdqGT6w6mvD
8o92HpxHQLGbwzaVTzOymTm2knFritRFh8x48+LUIEXVM1bCzKLl4XBu3Fhdb/8P
KTLltpMzvq1GE7mz83sn44q/AFRnm8OymdE51udMRIugp3mV253baKhH2xBuXiqD
SCq+SjQKJX6cpaKCrIqCjt0ILkfknCnmZeh1oHJeF9gf56diFZXbCIUJuu2y37tp
ugU1ZLxa7i4Tfn8/gu1bbPomnopypt7uhNBPeVAc3FEtUhSfgzvTiogcPrF4jHqF
hPhcu5JoXsDBQ/4L8frtvX3pj8mTvsbU2NLJMAMWSZ3FjrIWf+eGTptF+MADQ7vm
8xnOkiM9/+xGJfT3yTjV7q94TUjMfaeDdepdCDsZcdywH2sdV8e2IEGaw/euySsS
WiyBGMUogZigoZ0i63rKc6JSTFip23tsROMsF6t2IYucFAId652wLeSj492mE5gV
+WylS/i+p3QbDWRnTd1t6W9IJ/fA8OcncsXVuhR4uoU5QRA2ODjz1Sqjk7+QATLR
7nWUd1p+76qKEfToSafYfq4v3wWFM2KmLd4j2FdYX6O3bnbyAq4QJMrLjhjwl6yw
u8i6JovlUfWdXYmGBXbqQo4UU+k7zH3dJRnBpU4WmANQrX42zM9+s+2tQZHDJp+4
kvSRY7BnoTjZE0LrRJ6pPe7gSuOV0lTAIjZ1QnKY4LD5mXuIRCD11vCRIuRxHErj
4MPRRX487+PZmnXB4N1a+IA6YDpjcg+K8SAyA56Kc5QLurpjqx9c+hfFRw5G6p2L
i37tM0BCaECastLeQ2xCATqpAEubErFHc0k3UfLwGm8EtixkhL6F0K0MEYYtGtc0
8jkAo+xamSK1NJloWA5+Pf3wTp1k/+VDuKzhn1r1HVuMBV5P7pp6/nVWEI3F7rXf
4kTBRykxyWU3kETQ17HFnOzjrf/P7dX/f9mC1qt+AkOYqDXds+lYymUiFqbj16k8
EA9D1MXYy4Z9oBPqSSyD68Z4/PhHi8xPPg26nnr+MmZYUHVpjokQEcYukZoQsvGc
7jcHzybJJZyE+DBl8jpNJalcenL+cquZUFocPHPDczjKqRzbRTNrq1itVKRM/OkL
WQ2Ml4xjwn/KXYoUI0MxOVzrKwAM/CjhpfF1BEiNqlFknhAhDoF1y4ybBzcOanCO
nI97PbTda+jvD/k4zldmSwYYkHFm7aYPeLX5qC3Cqb1TffvFwkvUmBRc5MMd509x
zBM38+PVT4IPl+RWvfhU9vq7oZ31Wr2Y45O4qdmWdgsC68ESvZfgNQWuwdjkY3l/
Wq+xsXq9eeb6kLdSGmU9TcTOGKtgOjQw3bMUBNEuJUfCMaFHEVscvIT6yUb/wr8v
QAmZNg47zIfGndESPh1hNT1BzdTqzbYcAQfPUhWy6M06K/wvdT+Ddt4u+zs2dJH9
q8VMlW8RMnhgzosLpgUzsIz58rH3GD3jQnWUIINc+m3DFR5GhZa0AQUPtgJo4eHg
0ljePC8sG3rbUbqla2vkjF8NcuuUI83ZlZsKV8aUwVmuv0zXefD4wHN7FLRyDnXH
oGhsV/rql2q86T/9ZCgGWB4L1wxmPiFzmJjmmKMpQGR6y5I/Fdl439b0L7FmSjy9
8Oh9eLCvWXsm7nPPiluKQD1LojhFm/NePjD9xmmjmkCfBVwinqM/B9dIylqHt1yA
WfJxKDAUSBwgJxrnnMMZrlE6+W3PfIflaKORTkkm0L0LT+N6xSu00RYNQkt6Q/Sn
TwUSEnscNo7tIz1NtvW2+c0mackVxyH7Aldi1kSYJlHYKIAJLUItJGR/xclUytUe
I5tTVmoH8K6p10WbXiDpvrF/2z533qv+vJ2aFCUh10D8JRnFIJNcB+vmS+HuqHDT
SG1q5pzZhLmPDkkMKDAvBw2tHviQdwuMVjGclLVgzqZDaRff/TW63RlvdNWmQhv/
M9LD8wtjt+FV9e+l3ujNj1E5wXH+qzQd7yU87EERBke8gJemeKU7KKSP26T3Bqrn
qrGKGeplvcROA2v7AjPSDE1r2JiCoxqpTU0e6JkX+vT7PE1UQGVG9ibO0Y03hE+S
9TqkwQWbcpu9IrJ0pwo5wpjRVFSNWdF96clkmHcRnCpn5SY7eXSjzg+OGImhLSsN
PeJq4qxaxO45Rcu532+fnaJX8kQ2KuxRH0t9yweextASqGHybOHFYOX5fZCMPrxC
oQFwQCK38JDRQ4VSeZ5RCn/daZkeqpYYWuSm2Po+QusRmHl0VpJIrPDlGX8nO+mm
HNv81K749mNwciliBSI6YfX8nb+L9d7sS8aJ+SyC0jDv6GpfiSKWZdVPs9UwzFoB
LOgb12/x+S4UVnwUjDXwR+dXlW0lcpBwiidB7RcFUlq/MJge5zQm7aHqvL++Bx9A
c4IvcuGUVpiJXbZH22P2HOY8tQDOFnpteVTm+nVwMh0yITN/Y6zCYJiRNvkxTkUn
8RXXZXuh7CaLLUxoD3r0Ufa3lSAyDdUp+4m3yF/FbsYrPDlydGPuNPAAP5527g3a
+L7RFMBw1Ka+hJ6ReCPzfG3d1Nbf3skbm1rCJKF06ezm14yp9ra1mP4M1Tg6f0CG
jlTbcJj8dtV2Q0KNEVYZBJWILQqJrMtu3ajKdHZ0aRbwBwrUml3dbmT5Jn5woQVf
yNtJSf56OHrn+yvgdsGLOjre2Hkdco7XammJwrSwoHOnGIqHzfSatMrooYFXBAu1
tgPnyN5PefhsacVoOvstQwnD5wtHgxx/Pp2RtUqa+HtSEOKt1xUzQ/8DLNt2y220
3w9JQpsGceiaDIX4+z79rDHEZaUVFfGHxM4DXFhrSs7cak6oTQV71ji/uaHNG1kw
hYbfe/ptTHXQMjHyguok00l7PJ8CDT9v8rQMjmw/MtrtDQpA65PHTlPAcBkjuD6g
4b+QRJzCAfEkuZxB6C1ycgtsZh5L6gAtZRfETfTkOAOfydrGhjYp+QPr9gGwrRLD
4w9fG2u25r3NrWYif/bJwt09G6fGXw1ib/Z1pBG0z9cQU5BLe+m3GgrK/JTqeuLK
PJleUhAAh1IMkE2VdNYwQ/YHZUETIGUhBS8xM1ZcYdM9SrpAiGE2zLCijSCvaPTf
r3/WtNu2u8S6+LEPiWXJ9aPp9T7fSF9qtACm2r9vFsmoU8n5W0jTDYkBJbO2jjbj
tWf6ebx2SM5Lk0e9EnUMbJfsf4+xSkBQLFfx5SuFs8P95wmgKvIlgMOxlEkIwsGS
wuK/Jk2x+47iBqhukCPrxlt7NWnasuQiwGLpO1gCskw8jxU7kUpBqqpwVI1KTXsR
G4tPI0uCelrlCiXqp8b3yLDbFucHLLjuJSWDrl7tZDAHAgOlr3K50f8nv7yJg46y
zf5X2ayH0nw1dNadMqc9UpTwce7h4Xq5JLqoo0EGlxo45+bXwV1i0Q1oHEUnuroy
jsTmCVCv6xgoFN18UoyO1lNOx0eMte+ns4w4xtLHWkTBLP9vR7v5ht6SjiA5OH82
vK+yA91TORIqbWOm7y8+Sk7CcqCtJPoSSo0RZy/ZQZb7U9z2lMtXkfBwtjRf9cAi
zsRcauDJRBruPTarffMGAoRIQxtp/d+TCvRPgA8v2YdfQfcHGOwQoutKKm1Gj+nm
wnm65WAR8cP8bjlNiAaNLPvLdM/2G4wLR5DO73n0f8buZM1iN5cnU1IxJYm82dw1
PH+bcvXUS/sGbt57wpNG1B3CmJ/j2ya37mFPzwLPFFkiaDpplyzZ08fYxvtJEWpT
o2sxnHddh5PP0m3D3dTwWpAFKGcGBL52E7w+htI0Yv2cRFw8AiV73pG2M3N1XLeO
JOGS6SzpROVfD/7H7+dxg6HOjp8+UMqsAQYelONmo6NPo+C8O+qzoWym/fjKukCV
fZ0z0MJVUg8Xgm8Yuaf32gzBQJBgnmV7DdnzFbwlhjtpXA8PXA9arlRQ+Li9tdda
Mz/2NB7zRJfwMCWdEpYxBtVrNLcbdkW2hSq1qKRuG344F6XJ3cTo4RNALaMnZJUk
Q0gL0hRV2BDLR0KK2+sxlqHX07cqR7jlJqYx+7msmQozCBLGVUBflzYl7x16Odqq
9qESlin2gaErrdF+y0tirbzS1Amrw/9h9jYFuRlFNI25Fh+1txFyu3mBeoTkLD5d
aLQHsoz5M4urYbSDX/ej+K7PeJkf4zYUQ+NCFbWm8mG+neV+BExjJE8Dxi/hFMme
sBN7jxJbbVr7ehCnVzxD4n2yPyD+9HoPJhujY3hKis9/PVzSo1cXTRnbBT0CScgm
pHb6I7lLfL1q/lFTbvpeYapicvdBbN6RUt8O3C352IgfNX+2VRiFfu3tDe6a6Mkk
1fOi8NjB/CWqnw+jveDhsvYrl9ffCFoNM0q6O4H0yzqBlrAfuUqrZKvKO4j5H45Z
pL1Dd7SNRTNzMlTeJ8qXpzZEGfwlenfaNN2mZBgwvNT04QI7ud2sqnW5qvj2/xK5
l5yBAYhbv4BkcGu0xQFrRLWoZnsJDrjPgPzietYmn/CS2Jjc5PxYpZXQrqRsqPNn
ke6fmeEV3ZM+lR5zvBTQtVhoILFF4xAaJAzb9D3gM/AUmdVDd62R3zCShnw7BJYO
8VwKnjGhC/UQCPH33yE0RECoxgW7vK3zmjPKb9M750E2JkQWPfHPcOaeyqY98BCG
3sPbtaDtYLzZUcR1j0xfLW/drvTaXTx/qLIYvgiXvqsr03rNa8IS/SIpdsXIvcub
xKlRQIxxWaM5uu2gPw281W3pPALiy+Vzhwq28poSvakmn15Lz4tG+yZYQySKuITx
8P688RaSOy2iq3kH82tN8cw7OIJ+iEqp6BZ20ac6VzDslcX4SNg6C8eVKMQuxgjm
CeddUZW8/k22PHCP6ZThr0twW5rfdAjtOXdfsytsF64jdmRWI7UBKEgyi8YQLDMD
U2nu+ZW5yJKTO+d5yFpaAYvGn0fkOZ+X//JPObpvgIwc1UjuEO+9YQwcdhJpkeTZ
5/8OzPymel/0asa7W1h8lqB0bYfLU7wLnSJDYZ3xTgS0m2OvFYUukXFSAxdZP9H1
qz4JHYdGWCra519LYu04NKpqKDmeQpTleUjVW7nYcIm39KCExDRMXHFv1bEp1qtd
Nga4Bhqpqew5vBXQCNGzwBW+d+UA4fdi6fv9NwNa//pFXcN33v+bZ3sCtbp5MR2L
T4PnhjtdDV1n/GS9nyWK9aQpSW2DBVENTWzhX7s6sKR/OQqv9xGHNHqUnSnnrm9J
1CFz4sYz6qWvfIhDLuTEqL6YiFYGB0HdhViZd6AsNXtwJgQUiQYmLmkRDjmmr7/t
Hdnl8xki4RcBjljApqtsupCLnXlDWB5tQClmgf2agKRRExg3eCigBcZvpkZzRVwb
qf4mz4DtEbJmQtxkP/JMOrpSnAhMDzBND0GVh6V7iefdM+Z7cXpy6JQ8SFGAs1Nv
/F8ActoSjXpeReS999QsCFKxHOe4Kopf6Qzq0prMuXnp0lAyyKYyiPzc+HFOzu29
WWS1jP76L+quUiXY/lR6tQrrJNLdoijKYYYFHl5yI7CzY8f2+YxegxNdYIgypTgX
nwID0yRW8VNj2tl/NoVCfW+qjT3XtqBeNIGJI2ParTBYqhkuD0M7eZZwfTKL8Brq
cNoYnLX3uNF5Yrh4Ii/HKW9rWCqu3gDsy/c4oZvcVprxMZxxeeGg4UsLFLP9Rbl1
NsDYgSEjXPFmo+sJXYV8OgLQ0LGgWAG2zdgvIL/GrqaZPTqmhtVDR3rRygvaZn/9
gpooizIC5bbuV3OyDkiMXoRDlesVtJItBpNH2qjQpZGx2B9XCkj65Lye0Cm4tdS9
YOmFIkX1Cd9IHi48xcrEbFXjf5f295lm8uVapTvEX4NCS+sDIvSMpx2PI+OX4aZ+
TeELAQASCwEVfXjFxqqAr+3pZAym2OCIw4vmI1LUWJ9UkgBsi9wqaSSI4HJxqT1I
wihZAdW4Vw2B11EKh1rNlWGEMpV4EXd6ih3oVMZeT7xFQzESAZNkB+FvoGPA5/2W
r+8j4kYJbdrUeKVcb53kaNqQtUXRsTLphN/r5SZjFCFSF21hh/JMEhZO3pfQHHiQ
hxPrpzLzS0+I9FIxIP5172tZmwC2gJmVWD6a0AonH5LqG/Mm8b6kx40QQadx5pld
GiDhV8ec4iIYp/PBBeNQvg0Fq3YdRhbdRLeN2a9ZatITj55F4OUZaEMNRXNA6fhc
ocah5t0Qkwf1zII5o23AZNVv4jRmFZ0Jqs0u4sr++dMNNpPmQ6kEm9qyUA0NwPOk
vcj2idx/kwXDgQKW/0tEDa5KCdHyWnsBISnaXRo2Xfptto8F7ajk9MpaEkttJ5+S
d07Vhoqepx0k550/1CLq15YGpxywaGMAJ/+afasol3PvQqOibH8uWUGMjgby2KVz
CazBVT+FKXZQO508b4xhswQMsPkGA+mYZIVgTWG85KR7WgsmyT8z8m/M7LjaHk3N
DqPa36cdCmiJN8+c4Aiy1bCny2voeOvOE2koDtIy/MNvf8a393URzk3NktRwYUwS
8zERbW4z9Y5JYvSE7EgtyESyHkOI8kdqQJez88CZxi5wzOfYFH5Pp6doZ4imbUmY
FO9oqCdeJCzekU1ZzVQfNJW/rDUSZCE6xTOO6puoSHcHa9LS44SXtrOwaPeMPnJL
TNCGyF0tnZM/zgBS4TIFnLqAVlRzHEVDEqWOcnk8AZHzq7xMv1rXnaTqah6evPqQ
1OMSolN6I+QB5zFA1zicb4P10UXiMztTNOdeSXRjGdQuhyEWX1ibgYgmqQTcbd1A
eSy0IUI0QQCb91FWJmnfjpXqz9ublzyc2YvHNn8OM30+098aZdbEOCeLOWcybwY2
QqkCUAS+N9poUIkx1znuq3RCGU7vpqlTJ0fBEsWW4hzXMo7l+KR74Wj08EA8opSQ
xiSNND13EsSSw0dQLwndmTtGqxMj7y07SYWLMrvrMDPB7bNkQKYuueBk0a0/oJMa
93W0uxlbzDcepETKTrYkvQ/Gz9SsR8EITmJwReOA066x44k08qDJOdoWJn/1Ph6Q
B2VnHxGtRz8J/hcN45gcQyx3gWKTs6cSv1NwUNfXUUwx9KMyL4dWKxVkzfOTaebt
TblqcWaXLVTJixbZJWmSy0hWmIGpuME9qtDcevyoVzaHErE6BUx1N4PvTHRDjZTo
j7GozKzwQRXxLA+dgT646UPwUUuOlj/O0fhuAc2JVVeVIqQ1IuRKxzvHj7hto0DP
cVekBpStmJ9FDEJpFZf1Yo+LnParwlYVBD/vuptT1vcp5oRmmDhts5jgRQrr0ukQ
yAbh2ltnbCeuuP3zvk6YPKchIXZEN39RFUoLBVzIT6usCiNC286nIG9r9CeQf4qA
TZERycf0PjdK6FRbxYtAkPS14eYMXiXy85zzG84QlQupITM0Tl9lGchBK0YjT9BR
Q/b+qtNchNPrYmrPOU8vU49zGZoxTbG3eBTH3vRfEMYoN8d49Qic1YX5gpIF8EUm
ucacQWh/Ye/6fYailZ5RMIOXj2YgqQDvyPUDxtnwsmA=
//pragma protect end_data_block
//pragma protect digest_block
i/ZccyJ5N9GdaqCDnYqg5k0Yt2I=
//pragma protect end_digest_block
//pragma protect end_protected
