
`ifndef GUARD_SVT_AXI_MASTER_SV
`define GUARD_SVT_AXI_MASTER_SV

typedef class svt_axi_master_callback;
typedef svt_callbacks#(svt_axi_master,svt_axi_master_callback) svt_axi_master_callback_pool;
// =============================================================================
/**
 * This class is OVM Driver that implements an AXI Master component.
 */
class svt_axi_master extends svt_driver #(`SVT_AXI_MASTER_TRANSACTION_TYPE);

  ovm_blocking_put_port #(`SVT_AXI_MASTER_TRANSACTION_TYPE) vlog_cmd_put_port;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  /**
   * Request port provided to get the snoop requests
   */
  ovm_seq_item_pull_port #(svt_axi_master_snoop_transaction, svt_axi_master_snoop_transaction) snoop_seq_item_port;

  /**
    * A reference to the cache of the master
    */
  svt_axi_cache axi_cache;

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  /** Common features of AXI Master components */
  protected svt_axi_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_axi_port_configuration cfg_snapshot;

  //vcs_lic_vip_protect
    `protected
&4F-MOB]OU>5Y,@-C78TEO.Wg(.C<dLJ-PD59_^[5XeY;e.,RGHU4(#7DW.F;CUL
CW-VKKD(\9VgESdO[C#6K]fE\YWf\V+Ff=O2Wf/.#CU>#]WBCMT5YdKON3JRU=A@
.Hd/X#,&BW0?<ZI=2^YQWDfS<EM;<W_fLQ@2,TG#=OQ7T,[PVcdSg2>Q+4AR=W+M
.Fd1N9-05+>Kg)3F-YRO9F-f.d91+Ycga_>3:fRK](\R;I@Z9[fIeH394[D5<_+L
\I:;.[TD7SD\3,a[UCWFAB1Df78,2S^8VO=a,?M4OU2O^SSBV]#gR_.8P4BF/RBD
Za?_39A&GLdPgBXadbfgG3Y:JPY-::bd@aRGD@?I_ZM?e8J(@T5Lb[HTJ3VZf0A6
_ZK_8RF3I8/Me&=)XJ/ILDd&[DZS:b@-\c.]Be[A^,3-#cCV9VS-==PX8+9BQ[L+
UD>6BQ/YS=:PaP,fT&Sc-P<_CG)e2FRN_K<7bcW5<V,GJ6@HNg1T(/=eZV(dcP#-
4NAW0>5A04>#B.V-FFYJX30eP/+8DKZ\Y,QU=8eW-/,=J/;8338ReA5Y/9^[<8N(
gb3LZ:8/d7+E?de1X5[/RJ8e&I91.I,e4AMV^Y7N/2cHI>F,T>?53(D&a/<,H=eC
,=J/.2GT;f[N1W5Q_MC+W=bfV\U<e11P-fJGg#)GV2bcR5OH:\_fW_K<g3f;67[5
I)5@@;]AAZH76658[NS1[OYV<P4#G:f:6RA>;&EAC]1JM^)@OF7]XUJ992L?B)?6
-?OX(<_F(.AN3cZg?+2HZ:X6OF==ICK9e=@GB&b0Q\.AcA_2ADTFb6PGIOHFgFZJ
^+eUa(bJCJWA9N[PI3Q\MR3b.M<EUO5eGg1J+X;0.P7=2.>9d5;9.#4Xcegc4M_P
8)7Oa\G#F@BeWR?EGLfEGY(e_+f0@TPXTPAdc,)<@[eE^&4KH@5_XaC9;YSIb;4a
f)Z5)V&EY,^B9EZC-HPM82E8b]fC0P;g9=Dg4e+P=D\R+CLR8a<.d>#c7(5#Hb([
=c)Y:;3IFQ(SKMAMaeL_.6dK;FOTMT&]Na9a+4IM^2/Z49b<a9O?6+7F9DfPX.7]
M:I>>@(9GHWRD.KUS#)4R_#7a-=5c_-^I1\GUgVI[+/0&SSc4NQYdB)91#SSaP0<
C>Y\JMM7+aE[T\>Ce_E1BA#74$
`endprotected


  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_axi_port_configuration cfg;

  /** A semaphore that helps to determine if add_to_active is currently blocked */ 
  local semaphore add_to_active_sema = new(1);

  /** A semaphore that helps to determine if add_to_snoop_active is currently blocked */ 
  local semaphore add_to_snoop_active_sema = new(1);

  /** The process that runs consume_from_seq_item_port */ 
  local process consume_from_seq_item_port_process;  

  /** Variable to indicate if the consume_from_seq_item_port is blocked waiting
   * for a transaction from sequencer */
  local bit is_waiting_on_seq_item_port = 0;


  /** The process that runs consume_from_seq_item_port */ 
  local process consume_from_snoop_seq_item_port_process;  

 /** Event that is triggered when snoop is added to queue */
  local event ev_add_to_master_snoop_active;


  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `ovm_component_utils(svt_axi_master)

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new driver instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, ovm_component parent);

  // ---------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
  extern virtual function void build();

  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads like consume_from_seq_item_port()
   */
  extern virtual task run();
  
  /** Report phase execution of the OVM component*/
  extern virtual function void report();

/** @cond PRIVATE */
    /** Gets the active semaphore */
  extern task get_active_semaphore();

  /** Puts the active semaphore */
  extern task put_active_semaphore();

  /** Uses try_get to get the active semaphore */
  extern function int try_get_active_semaphore();

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** 
   * Method which manages seq_item_port. Sequence items are taken
   * from the port and added to an internal queue.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_from_seq_item_port(svt_phase phase);

  /** 
   * Method which manages snoop_seq_item_port. Sequence items are taken
   * from the port and added to an internal queue.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_from_snoop_seq_item_port(svt_phase phase);

  // ---------------------------------------------------------------------------
  /**
   * Task to drop al objections if there is a bus inactivity timeout
   * 
   * @param phase Phase reference from the phase that this method is started from
   */ 
  extern local task manage_objections(svt_phase phase);
/** @endcond */

  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_axi_common common);

   //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void post_input_port_get(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param device_id_queue A reference to the ID's of device type
   * transactions which are currently beeing processed by the master.
   * 
   * @param non_device_id_queue A reference to the ID's of non device type
   * transactions which are currently beeing processed by the master.
   */
  extern virtual protected function void post_vip_randomized_xact_id_update(ref int device_id_queue[$], ref int non_device_id_queue[$]);
  // ---------------------------------------------------------------------------
  /** 
   * Called before driving the address phase of a transaction.
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void pre_address_phase_started(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving a data beat of a write transaction.
   *  
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void pre_write_data_phase_started(svt_axi_transaction xact);
  
  // ---------------------------------------------------------------------------
  /** 
   * Called before driving the first transfer of a data stream transaction.
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void pre_data_stream_started(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after randomizing memory update transaction.
   *  
   * @param xact A reference to the memory update descriptor object of interest.
   */
  extern virtual protected function void post_memory_update_xact_gen(svt_axi_transaction xact);

  /**
   * Called after pulling a snoop transaction descriptor out of the input channel which
   * is connected to the generator, but before acting on the transaction descriptor
   * in any way.  
   *
   * @param xact A reference to the transaction descriptor object of interest.
   * 
   * @param drop A <i>ref</i> argument, which if set by the user's callback
   * implementation causes the transactor to discard the transaction descriptor
   * without further action.
   */
  extern virtual protected function void post_snoop_input_port_get(svt_axi_master_snoop_transaction xact, ref bit drop);

  /** 
   * Called before driving the snoop data phase of a transaction
   * 
   * @param xact A reference to the data descriptor object of interest.
   */

  extern virtual protected function void pre_snoop_data_phase_started(svt_axi_master_snoop_transaction xact);

  /**
   * Called before driving a response to a snoop transaction. 
   * 
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual protected function void pre_snoop_resp_phase_started(svt_axi_master_snoop_transaction xact);

  /** 
   * Called before writing into the cache. 
   * 
   * @param xact A reference to the data descriptor object of interest.
   */

  extern virtual protected function void pre_cache_update(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
   * Called when there is change in the state of the cache. 
   * 
   * @param xact A reference to the data descriptor object of interest.
   */

  extern virtual protected function void post_cache_update(`SVT_TRANSACTION_BASE_TYPE xact);

  /**
   * Called when barrier_enable is set to 1 in svt_axi_port_configuration and
   * associate_barrier_xact bit is set in `SVT_AXI_MASTER_TRANSACTION_TYPE class.
   * 
   * @param xact reference to the data descriptor object of interest.
   * 
   * @param barrier_pair_xact Barrier pair associated with this transaction
   */
  extern virtual protected function void associate_xact_to_barrier_pair(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, svt_axi_barrier_pair_transaction barrier_pair_xact[$]);

/** @cond PRIVATE */
  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_input_port_get</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task post_input_port_get_cb_exec(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_vip_randomized_xact_id_update</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param device_id_queue A reference to the ID's of device type
   * transactions which are currently beeing processed by the master.
   * 
   * @param non_device_id_queue A reference to the ID's of non device type
   * transactions which are currently beeing processed by the master.
   */
  extern virtual task post_vip_randomized_xact_id_update_cb_exec(ref int device_id_queue[$], ref int non_device_id_queue[$]);
  // ---------------------------------------------------------------------------
  /** 
   * Called before driving the address phase of a transaction.
   * 
   * This method issues the <i>pre_address_phase_started</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_address_phase_started_cb_exec(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving a data beat of a write transaction.
   *  
   * This method issues the <i>pre_write_data_phase_started</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_write_data_phase_started_cb_exec(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called before driving the first transfer of a data stream transaction.
   * 
   * This method issues the <i>pre_data_stream_started</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_data_stream_started_cb_exec(svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after randomizing memory update transaction.
   *  
   * This method issues the <i>post_memory_update_xact_gen</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the memory update descriptor object of interest.
   */
  extern virtual task post_memory_update_xact_gen_cb_exec(svt_axi_transaction xact);

  /**
   * Called after pulling a snoop transaction descriptor out of the input channel which
   * is connected to the generator, but before acting on the transaction descriptor
   * in any way.  
   *
   * This method issues the <i>post_snoop_input_port_get</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must call the super version of
   * this method.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   * 
   * @param drop A <i>ref</i> argument, which if set by the user's callback
   * implementation causes the transactor to discard the transaction descriptor
   * without further action.
   */
  extern virtual protected task post_snoop_input_port_get_cb_exec(svt_axi_master_snoop_transaction xact, ref bit drop);

  /** 
   * Called before driving the snoop data phase of a transaction
   * 
   * This method issues the <i>pre_snoop_data_phase_started</i> callback
   * using the `ovm_do_callbacks macro.
   *
   * @param xact A reference to the data descriptor object of interest.
   */

  extern virtual task pre_snoop_data_phase_started_cb_exec(svt_axi_master_snoop_transaction xact);

  /**
   * Called before driving a response to a snoop transaction. 
   * 
   * This method issues the <i>pre_snoop_resp_phase_started</i> callback using the
   * `ovm_do_callbacks macro.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_snoop_resp_phase_started_cb_exec(svt_axi_master_snoop_transaction xact);

  /** 
   * Called before writing into the cache. 
   * 
   * This method issues the <i>pre_cache_update</i> callback using the
   * `ovm_do_callbacks macro.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task pre_cache_update_cb_exec(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
   * Called when there is change in the state of the cache. 
   * 
   * This method issues the <i>post_cache_update</i> callback using the
   * `ovm_do_callbacks macro.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task post_cache_update_cb_exec(`SVT_TRANSACTION_BASE_TYPE xact);

  /**
   * Called when barrier_enable is set to 1 in svt_axi_port_configuration and
   * associate_barrier_xact bit is set in `SVT_AXI_MASTER_TRANSACTION_TYPE class.
   * 
   * This method issues the <i>associate_xact_to_barrier_pair</i> callback using
   * the `ovm_do_callbacks macro.
   * 
   * @param xact reference to the data descriptor object of interest.
   * 
   * @param barrier_pair_xact Barrier pair associated with this transaction
   */
  extern virtual task associate_xact_to_barrier_pair_cb_exec(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, svt_axi_barrier_pair_transaction barrier_pair_xact[$]);
  

  /** Gets the time at which an address was invalidated due to a MAKEINVALID coherent transaction */
  extern virtual function real get_makeinvalid_invalidate_time(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
/** @endcond */

  /*
   * Returns the number of outstanding transactions
   */
  extern virtual function int get_number_of_outstanding_master_transactions(bit silent = 1);
  /**
    * This method is used to get list of all IDs which are currently under use by outstanding transactions. However, user
    * can choose the type of outstanding transactions this method should consider while extracting ID of active transactions.
    * "mode" and "rw_type" arguments should be used for this purpose.
    *
    * It returns '1' if total number of unique IDs currently used by active transactions, is less than all possible ID that can
    * be used by an AXI transaction. This helps in determining whether randomizing ID field of a new transaction which should
    * not be part of the all the IDs currently in use, is possible or not.
    * 
    * @param mode Type of outstanding transactions this method should consider while extracting ID of active transactions.
    *             Currently it supports following modes (defined as string) ::
    *               - "non_dvm_non_barrier" => all transactions which are neither DVM nor Barrier  (default)
    *               - "non_dvm"             => all transactions which are not DVM 
    *               - "non_barrier"         => all transactions which are not Barrier 
    *               - "dvm"                 => all transactions which are of DVM type 
    *               - "barrier"             => all transactions which are of Barrier type
    *               - "dvm_barrier"         => all transactions which are either DVM or Barrier type
    *               - Note: if "rw_type" is set to '0' then only read channel transactions will be considered for non-dvm
    *                       and non-barrier type
    *               .
    * 
    * @param rw_type Indicates which channel id width should be considered.
    *               - ' 0 ' => only read channel id width and transactions should be used
    *               - ' 1 ' => only write channel id width and transactions should be used
    *               - '-1 ' => common or either of read or write channel id width and transactions are used
    *               .
    * 
    * @param use_min_width If set to '1', minimum of read and write channel id width should be used otherwise maximum.
    *               This is applicable only if "rw_type == -1" i.e. no particular channel id width is specified.
    * 
    * @param silent Suppresses debug messages from this method if set to '1'
    */
  extern virtual function bit get_ids_used_by_active_master_transactions(output bit[`SVT_AXI_MAX_ID_WIDTH-1:0] id_list[$], input string mode="non_dvm_non_barrier", input int rw_type=-1, input bit use_min_width=1, input bit silent=1);

  /** waits until master is out of reset state 
      @param mode if set to '1' then it waits for 1 clock cycle after reset is detected deasserted.
                  otherwise,         it waits for reset to be sampled as deasserted and comes out of reset
                  after waiting for the negedge of the same sampling clock that detected reset de-assertion
                  to avoid any race condition.
                  values greater than 1 shouldn't be used.
    */
  extern virtual task wait_for_out_of_reset(int mode = 0);

  /**
    * This method returns list of transactions which are currently active and pending inside master agent.
    * 
    * @param silent Suppresses debug messages from this method if set to '1'. Default value is '1'.
    */
  extern virtual function int get_outstanding_master_transactions(bit silent=1, output `SVT_AXI_MASTER_TRANSACTION_TYPE actvQ[$]);

endclass

`protected
BN&^JGcO/88Q0;/G3-_A06\WaU8K;McBZZQH)8,5C\6RW+A,U>Y[,)3a-\8WL4EK
/E2E3;3b)UeADOGBK_TRgfB:FQdN:Z>W5<X,AL230==dbU)3/4VMY&XQ/<?C7F>4
_UB44R8XI3A\.Z>U&=aVbD<[L:9,TLO).GfERJG@YUZNYV.F)?0TY_=cPf+fZ/ac
_@H?H1-C5d(;V^XG0//X_g,-Jb?1I8I#<2NC,a,3,F=T#B&\H.@)aa^O^IINf?<(
DV_@-cSXgPd@.XEeTfX9NEG3dIV7>_[)^8G(^L_D>fWQ+7H)#aUN+.W2@A86=M&Y
Re-CaWS;EV:I82MgRfIX>_\NKb(8W,E[4(6\#52RR?G8RTWXTFbgGYbE>f&Vaa\X
cO^#e.JT1?.R7DWFI=1\1C&-Q#@#P08FJ-,[]HUg(g9O-dWa2e5G=C+-3AW[KbM_
(WYf\]8^dGL69AG;]30)eOGW>AE(2eHF<4VTf#]2?N[eA4>RECR6Ng_TNgc8GIOe
/RFagYW\+eJ[=T_)ZJ+V8dR1C9UF9S=NU?\?Y9.<X<5/,5(JTMfd4DfST8N9YaJS
+R.D<.D832)[0$
`endprotected

// -----------------------------------------------------------------------------
// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
B^D(MW/=V9+>2?WBYKLO7D)ALeU:AV&ERO]T.>&1V_@bM[8Y(WAA1(O:3/2\BVN]
=4I]fE8C?)dGC9@E3ACTGO(,#]+VdV8L)UX3.2HIAd3+c3Q=@[SB.Sc)I5SNC>cN
UTdQ48E9&DO38XVMBFb9fc)H;/K_G;0\3fdDc;7KG.^SK2bXEa&^gWMcSaLY?D?+
G/AH&4TDOGa@ID.IMBZ#,<78NGP]eKK/=9OH7LZ,Z](B[JC\bO;4B]S&F1B+=//@
G4DT)]R,I6,fF1T:NYF(D>X:G=TBR6E^gPHTI4E,BAQ=#bbY7gTea6d,#=&MQ2c0
)PH>1S-TDG]>L=&2-HLA6I2GaI\/K56D\R[/W1[JE,N13-+5WRC\@-(d?2EZO1)=
_eQXYfIR=1Bg_0[@+1I=[ZJAMZ:Y#3JV^IF,I3A33Fg:&UGbdg+3T.d;8c(dS-JP
)>ab4IDC;JJM665eUACbZ;/?=&D8=9I\?F/7UMT++3@/K66Q)6Q&;D?24H_OM71S
8=DEF#,;c26<?&a_&:;GgKbGV53/&M-dVL-Ad&?Aa.4JD^?V6G?U\X>K+/Z\cdP5
757A]D\&GHNMTK5>)#2aDLY9M#,IHAdS9NTZdbJ(JKWNJ;T]2YJF5T<Vga14DdQ.
ZZ,\?9N8=IKBCAX4QDU3UCX91,1+W0IX7/>\0f8/4ZZUBdE(IQEO46#L)(-dLVAD
9?YMc7H?dJ7_Z]_S(T3c+8:R1X5JEc\UBA>;ORLXDHJV9U-XZ?&)HLU2+^MDUdZX
])[=01-8R6Y,fST5U5J7Deg?LF.KLO&7]S(72TO)KN]G;G.GMU.#K9N,;ET4.d\b
3JRLD01UIV?9f9_X59IY&0=b[:fKD/EAc-<gUf+SKdH)A^AFBH_B88DC->1Le5:I
ML/a<X=H]OfI3:GP3E^LDSJRdSRQ>3G;2ae;.KDB#&.L:ecb[>UbCMTF6RD/M=(^
A+BdZ,Xd97;:Gg6?\bP6H85M^5PX8XH(UG=RUg711b-N/;J,E6E;H>a)aVT3H,Rf
L:5YQW-P[O.&1@ZMWK+18F6<FSQP;V/.GdCG)A^I[B81,5a#W(9-:E^YU]J_?P@5
H556eL&QK^FeHaV\EACKb-ZfK\TGJNe+;1X0b9Tace_3(XK)55;TBXW4])X6</J>
EX>OdSUDfDMPW;]OEIL<3@WA1&LZPXTH6]EDB,MT8/6c80/(dJeY@W1@C2L&U&\7
\XEL#W/8>66\cb0X@3c;Y[)U_AEG(W.DgP,FN47Q\.(cg35\CgR#f^e)M)JK@AI1
gM^Z1TCJCW-P-:[4QR/S3=/?8G;/=6O(GDWSN.=\.D0BZE?UGc?OSB@VeL]]a+/5
GM1fQE+^d9#C6=+CDLdU>O^(TKA_#U5SP_LI\#d;@6H1<EV(;Q&cM+Sbc_.P3=:E
.V]]GVKKVdTZN#RNX[,=Y]Ee)::ce@Nc0,CYP,5;c=##[7=@-S61KVELUf_<cYX&
:KTc0/<]2Bd[L[FQe?HBN+8BdZR5V:HH32(KJ/\X.bAXTM0;e/3/B[]/,?<c6).P
R7;cbQU-TJ>3(YWMWI9?eaX+>O8JC]a.S@0Eb0T7+^8[E(gFO84WIGf>bJa.79P1
dG5-X3-ZY+7g05U^O>]Ka@V^O</.9UbX\]A)R5dH;\Qf1HbS4P8]V^CDc;TX[Gc#
TP@;N(T8-YELFF)b(1^4GKaDPJ;?-0J0M.[W+.MKNV3SA@/DFZ5,R37&3O1:5:SI
5FV??(ZAd=#3?3PNDQdeG8dJ(1?C6\,8Xf>T.R9C#S&B8-J<f45T@(MJ60R3-bJJ
@IQDa?G&b^e8I4[c=O4]T-H]U]b=gKA_#LDWG+,7RfP_:gA4d8gfJYa=Ba,G6(<[
EEceSf4A#_(-IHWRDGL)<A8cZF:Tc3FBd?Tc]6aCZJ;G0U\]580b>N&a0XSX(U\S
C4A89GZSe(;NFW[MgEK;UJALI[789OTK-ILRDF5VJ78:=IXgb8NI&]U47]QN^;RR
2g,\3eKZb2;KH+(AFB/gQ0b0&E.EL8F3IQVC+5CBdBBU.g+3ZCD_W4EIECI6Z,Re
_,NJO1\ZBe@?G01cM=]];SX^#;RD;WWfLb3(]:1(DOX&IOdK,3MaEEgT12C3QGOF
N4K5:]IN=:C988LD[#_;0.(fBJ-#M_b0;&</@1)US4@];50R#8:^8&;]IDb/1U,8
@;cdT4cc8&3@1gH1>^_7O/F2H=,O;J@:a6Odb?/g5<97OJe];cMEW&a:R[Y2Lc_U
JgDa.0cIS9B2H99RPfbBTd/Z@)I7T&g4QK:@6EHO7Cg0N=./N2f_04S[Gf1_&(Kb
\O=E,IY&U.3AA14>[E9cJ03;_8:+F/IDTUd7HB7ECP2B3UP3fK@#a#)=L#\1;H5Y
Ka5.eKHHPFZE2aOHK]F1VHCc\9McCZ@0:gW?N:#5A>>[4ENYT]LM#A7B&O)GEfKL
eOLO4FgC4U5I6IB^@bfF;=VQe+P^&A/L3a4L=@#W8PW,1KHOYSE_W-B164)g:^fD
<:cBbES)C80d6VOP)gW,IOWceH1G,/]bS2DB4aa;QV[#8FI,_&fRc3JGOR4TMd,:
??MHVOS2ST..F<=ILaZ0>S+XOHG\P:;FS.[LP^04,6RRLFU1[1e)Fc)H.0R4FbG5
RcO>DN1Q^1HN6VHFAL+cXKR8@HLK]XT/#-AcH3ggf9U@-U_R=8\>:S0(_X/@a6F1
6RYO8)[7V;a-#R,e_P@-KLZ6N2d)[gX=0GG+D2>VVHD0c:2cbcgZ&,53+3.XG#0M
UfFd0SA95Vf[S.)+,CQ@4P[TcT7&OPPaV0Fe,HNF;:<-KOG1,/I_6()BXZ-NVWe[
XY[]+)M:WK]JZ15ID>>HV58V+ecUgTVK@8\;R:]aW?&>X=_0391)4>1aE-[cK?[I
4af5IM3CA;HJAG4?/V.3SdAfE[HN18dZA[+=B04OWY)M>SL&DdfSS&(J#T5FZ+=8
V(]Q_Ud@-D\U[EJM-6#eF<.PA>CV08W\(-(OWB(X8@e.\XXA1Y.;I\IYWg-L6SH\
f.c.&6gXQKcLWHS>E/1eIWV1TA.5bA/UY;f,1f>cM^a3XBSQS_aRfD0YTUc()&O:
M2R.Z9)fS\gY>HB#9edg2F3.eI<7&Ea+VQa3>QSP8\0)TfFaEQ;]?7Q,S#UC^@Lc
b]4?>fZ0(^F?V6e]9bO8DBHaQ<?2/68d42\,PAaAR94,K\BW8X>^O?\E(QZLT7:4
5;G(05H/&_9:R96TMeb4;_7c]V]aL/NAIS>UU\_]=>WUHZQ0[-=Y@:FN^P:Wc+6^
5[RZ/]I-dR@5[]/^=d9,:aN>>KNSLLXR(f;5]+F?.Q3-@^<A8[;R/5/?76D_9+f7
(28))30=[&?-L7U&[[]1T&E>Z)NO6#KJ<LGZg:^/QdEWU^I4#N,g_YgFT?NGQaN>
Q;S?+J]L;XO#GJ0>-R>8Y]EM3Rg68&;;-MO)DY05CW;Q]N+H.eG;_,e:CEVH@N&5
/eed^V;^>(a5T/PZ:@61_UU?C+8([]&CV^a+989FEeNP:VQU[Q@34f?SY<NC:93X
S7#-dFG8_(=aHM22?2Xb5TR?Qa(d=J]f]_X#+P;[TSc?B\]/Z7e1Q1HA,QbZ@S3;
X]/&+D]I)O3L9;0OJ=c65>/)V-G-=acHQ6,V2Va#H]UIU+>gR\F(4YR3f-=UHSMB
0)+#T.><+K<^&fBE[V&KS2]^>9SDB:O:Rd&MB6g#P6LeCf9Fa2L)9g2b_[,eO2Of
7-,NDB9TPXdC&XQ8SY[T<Jc9>V_9P9(.:<R];KZY8Lg0X/M/,dC;aRBLQ>1#3aKX
ZZHSSQ5S:g\3f^A2_g2P+ERE>,>7=JUS?[/NK]Xe=S<([@P952+[4.T8:SVW;V&H
G?4]JJdYd\#OgccNQH1AdD2S6;[-.&GJCbCRR?]U:bDT&d7YE/fM0XfBD[#[Wd46
AJ[YWMIX4)M(M-R2JGD43L5,Qe1A.XITIHS2PKJ/QX5,4g3+:VRPC^3)R?d7Z-(2
L6\R-.UH3J&AYZ8(\L^5Ab.C;5ZUG_L-EKUa,#]AN/9RJa5O8Hd=/RE&PM<XaK5X
:IR3SD,FVI^A8<2b/99HdScN@_.7PNJQMJ<_87?-C=V]C2E(0VUG>1VgG<:.[ZSa
4:Bc?1K8:\#>b&[:A2AKBIdc[^<@c]5EVUgOAO?2+\/BF24&-IB/4?E/(2O;RT>D
b8^ZOD+)1Y?U_U5<F_@J761N.9G,E)d^:(N\2ZS?TFPSGdAV\KK8?72gf>U\e458
Mc+4UaPO)_/0:;3PO_J^F.W>F1E)<PA=?F,YcWZAU.&=C>2J\CDWDPM[?H3TNE^L
VXa>QT2;CX2&P+\/,We?9EBN36,<OdNe,af;&QUUIg2V5acN:/6ME8W^\DMJ]40W
DS2Q@9U:6X+9c_Q9NOT?VegBPMQcNO4e.YQ2L4-BTg];fSbe0B-X94Q-)IgF1LHK
UEee&D-^A.M&2IL2_[CM#e]YXR->dMCd)HRE2.b-9DNO=FM&1^=#_a@:\BcbY55V
F0E1/,39Nb9FX]A=77H6-4SUSCf(>U/W(8A9>N#.]?#)g/.^N.L.d]\?.aLZS:V3
((#6[.TX3LH?K]>T7YGMP/.4J,KH]-\-/Yef[cU1R4D#XX:QMeEIFI+A-^KA6UN[
I.L0fe_7,Z#<AgN62&eN.VNQZeW_;=49-&J/a/LeQ1bZ4Z2SZUFg+K=AF_]>d41g
\F1>FdVSc2a\=NdF1-JXg:7U^E;QO0#V@;UZgTP/MW253e(4c\YZHT,9Yb&]Ged^
DMVS,+K68/ZAeWFQ,]eKA,EdP>b+b1-J?E___0<32DCE/3JWAP#,]a:BQ5WW=97;
X1(&ee2B:ZY16b..1382XS)260/>T<ANSN:WL^O7KCdH]KF/_LDH]7WNgCDL&.=#
A[bX@=UE&6/NX4U[O<71QZ+GM_M3YL<+>?8BM?1_f;<O9)K&O0=^?O0d+K?GZa&?
76LQKVdH[K&Z,5-/>>ff6P29f#I:^@Y51=_^IF(Q0:1U86;X?Ge/9.L.e#2L2-6d
TEEC5+SaZ(9#L0S8PSCBe7UVUCD64VdR#,AB)bHc67)f8\;C0PZ69?CNB<JLL32,
00\YgH7C]K],fG9V:O8NQ;CeS85aZR2e^Ie?T;2NQQJb,=,XJJXLQ]I4+R(B1e.?
NJLF,GNAU>#.VIC#X7ae&KCLCW31)e)5+Gc><SA,RedM8MM)a5\8b-OTUI<.5_>8
1G_PI0#U753ZWVF+NV-.3AGI)Q8WNg&Rae_=e>dQgL?7A#M7;ZFTb9a:+Z&W^8Y(
VYUSYOK9?JO2V[:LTJZE8]S+,\U&Xb+;8N#OfDHL,K^6N6PM<6PcL(/=S]gB:bgJ
,2QOT8S#N<XI-d^T;&0YOXLD9NY-1X/B?/)XaKdTO17PF:;H]Q=JG[>Z(>8a0X/1
9a6#g2Z#H,e+S^)RcM5^C/-eP[Q/&&AAX?EEdI5eFB:d=0b=,K2@.C@I;;[+)E3c
.H?G&c:E.Qfd640Dg=HA#T-:8X@=N-M3O\EbQLKPJbML(+^.BNa3\SZTLQBS5=P^
BQc4,d.feVZd?88\G+WZ?L^WH^36#M0/F0-T^=T?3+A8&83Bbe@ceZ6Hg]<B940S
I[G>/f/9)eI=>8+?aDP?LE2&YA8:9QfV[dA?OKJ5IKO/+IXV\-2^#71PFS<WHC8S
M4#,ML_QKFYeYIGcXQ;:];5/^9O,/c:_.,46YT50Cb:W@K)\b+05]=ALHfHR#c.J
MAV1S#KET&)5d0SXOIN,[303KLKM2IZK[,fL?0C\]])FfXeW>f6HaQ<<M#]=11M1
N^8ad6B,GL+fOLRd=OU-(Lf-,gKXM7gaN8fBe=J<6P+]b#(KTJ;</-0gI9N=+7[Y
]9;E#?3=;R#g&JVK=0B;W?R9aZ69?Y85/[_e01OE<9V/N+3#9a@U:9.:#/J#.MH5
^-\Zc.;,dBVA;:)V(?0N7(ZQN-(@cM6PU2S-JRUS_]RH>]NM8f+KF40^I+AY.0TW
TAc,H7IUNE6a7D,?<0\O59:7R#XWUDHe<UW\C.C_-(bIQbNND;<56S>.7U61IT8\
NS[D@M=]2NF]:cAgdGKfWW)H@6Qg>N&Y(_40[W\aLH;=JSE)VcgQWVV=5d650<@<
](J0C1[.KQ)J7,?#[YGJ10:-,gB?-NUg)dA10Kg[A4_(J:,3XMM@@[QQg.+bPd1-
(++I]:>E&[,AC&,88)+VgF3cV[^\6.;IKA+-YPM&bJ@1?aaK-N4;@]B@N?3Ze+BP
FMMag+B<E/.D?@F6;GIW\/K7,6UGe,Z[D]AG@f>EOgKW0[VNcb4Q2\2>X1)c#W6N
V8V-RAcT:^@73OYB90L#>?=9/QUEO1JYf<V(/6RgDV6KVVC\E#<<S@GV?#M>N3D(
B+;L;PGG)9^08R+R>ZS;/BfV4#dMUXYFVE8cBBX<N/d\(d[)3N)ON4;3:SAOPP^X
UZD85GaQX_9aDcEGg6/M5[gSd3YZ2bIb/aQGdc&7V><TY&D[ID=?T.b89Uf/V=Wa
\#?B&0]6[RM:OYa9:]G7.HL<>V(Q,D7(,g0a73,R.521V.R/g_^?B[T##2cYQR>N
@dE@(&:]-6PT7UV&)\9.S3^0LE@VG.Q;d/\+a6f/2(5ZR8MYAD9<e6HgL@EBY4aL
]0Oe=]@J70=5@]^IbCUZK+fHBF[A?MBI^9?aG1V/)Dc(0WbDUS+eK075bSLUNWLR
.5_HIdRHB2a\&)OO-LT-&5BFF3,#cVJ.8?]YeNaEH/0#>\6H:MfSP]7([I0T?-P#
;bEAH#@GC]1U.#DE6PVT3bCa#M-2,5[:LK3LI/.L8TH80QSMS;,;SJbGCDP@8WG4
@4Bc64P+=QW2M2^A?a8Dc3K@ILL/+WY:S\C0+);0[NDSBdY>NHHdeYc4X,Qc7-HK
.UXQ.<S_KNK5U35G53&We^T1:336:3#OcGDBLVHL;&KEVO1;1Z_].a]GO1IS82g@
?AG&\B&[QJ4fM.cPV92@:f;^P76=X^<#(@G?IB3R>&CRdCC_d>.Y6gL-NY;TG)<Q
6&=R<4XJfcIEL6/UWR4gZaCgO[@bJ.BYgLcG#<UMPST?^a7Ee>]ZdZA>.WS.c0L9
9SZ[++f8Nd[I)\1d6df36FN@R],.LM,eUc[#L<.aM^5XHV+Wa;XS0[#<+<dZHC0?
4:[VdR1)EGT2EC)Oc4B/&eGO_M&]UHP=9YGC,RJYBX#KE/6;8^TQ0=9^8,U8?9F8
8fGBdK()>7D&W][D]S:#XTM#99=+1^\<=4U7E[9P5)dOZVQ1PfRd53ZQd8f9V4#@
/2e9O9<cDeH8_Y;P<(1\f5eHUU:V-0@^fNC(f3Ue[:U/<R/H2GZ.&=N5WAN=@aZR
c]?NDENJW[U-806FQHRA/E)V\4]B,76Sd[g@-cE;J4dEAW(1;?cM^@0a-O2)5_HY
2>&Ie1NcR#2YQ[f7BX))NeRDA2,7Ge?R,ega]TMDa5OHb(DM[aEJec(E)KgILO7F
LE_+R<CbH\FbY97]+)56eB=fFM@392BS<17gII?RV\6<4dX8+=.]CgQ6KHW4]Q[?
ZZ0a.V,1@BC_EYR1W^L,#f5c)_K069P(37fJ]7eZNU0K?HGGHFVOHN90WSY#V][B
>J)&I&]GJT&IS+-AfV>U>+:[ZV>bgOC8:d28KdR,):-9U3W_YXIO<<VV3KgNCdCF
]66E(6<DCUb1,/b&3+&e:,L@FRV1W5g^@5>F@acHA:FCIQZ>K:_c8Z-U(H02PAV>
Z6Y:2Z7IR&dHe/c/1OC2/&_MD=8O=/>dQ\,+<S[Sd^TH^7C3-9#510VH6:(<Y?BE
>X=f;RBI1X76g7P4T.XF?ND.bEN2GFg^RRNAT?d0_SAT:;gaX\HZDc[V=N5J70\A
4-&5JJaX?,VN?[+]&9G:JRL2P\Sc^KacCR(9U4+e-G41eKW^UXY#3/e7CM+D;T=N
TV8B\8.E_bG;GI_MXD.N(1#[SE?.AfX9[)F+Y<\+J:\(RVdC@e@_gK2@T(J]&WCd
_:f(c416>efYE]FV9&/7(TQR5\HO4cOSe0E7Y2WGL_1)D]>7f4<+NW&\_3+U>X):
QF.dRSe=#4D@e866]=M^<L<baKO4EBW@.&]N@34N:d_=V[-/FeE#C,BFEB<8fUD1
=Y];=1.R5gC^9)DWe<]/+;4\G]UaSNOGKZYIUMfg,B1__8ET@PA5YRZd^C#aO+WP
.:2@<N(SfT9O:X?-K+/b+=T:aF2=bK=+1#:AS9I5]Y[9N_PLcN#.48,ZC:QNUOI7
RDfg2\b)K?,SGV50b,OLB/fG,;H<>YZ6g@5N./N>\<OB3QXN8OSA046/7-?[E&0[
@:/:N99JYY2bMP8(^R)^&g78WB/fLD/+A6YN-VKW5g/-c^+AE=XR<Dg@EZ9=YgO8
PQ>g58:EUa1b,$
`endprotected

  
`protected
@9ZC2J8Ca=EA#J5B^S->HfWXb(.g]I\OM[cXLOQ>gD@;44WY9)DY+)I7H;4<OQ2&
M6\>\@_=3S-3OD7NHcgW8>WX5$
`endprotected


  
//vcs_lic_vip_protect
  `protected
d.=DC6eH@D0^>V.F+,K6YdI?<.&>J0c^_>6)DR_3(T)V#:e,L9NO-(<K4,>->::L
5@PdL+BO(/PCIYR+;Tb(:;UD<U:6G8LZ\]e]-[3#\51a[5E<G6_CE)RG,.GX1.>9
1b<;/\?Q[A);XR#9@JL;YB,)-J>/#V8&<7K4W8SR&&Nc&L1d==<Qb17DMR)1,f3b
K\RM:?8JMb06ebG+7+J1XGc@gM[aO4KIR&Q2R,0GPX?cVZXdDVKMA\(;Q=YH7ZQX
5MB>>2K5^&9LO4^V^#^X7O#6IKUO[?cK.9fc.\N]GOAe?G2B/NM+C\H7bc6QU.8@
aKSAH-]3=d2:fL9Jf,U>-AL6Y\9+JEWd=L+bH?EA<3<cW9dcA1_G?3Zc<1XK__Q3
(?.3[&->eb8N0?g^P8],@DOC.1^0K0JON4#TDbL@,PMWX5:,Jg(]c/&R;XgWMQ,;
KM]=g+9d[ZB[_Q.66:EG4(IeXJDZWE@V2VCg\,KgIAWP+/(.HaDZ>JTP6J(_cE(A
/[T=4ZXYegB=JXNE4.^WIccOf;Lb0^L7;I-9ZE-6e<0AJ)0REH\e_&]-cQ&Mf1gU
>.=N_1ZR52:\eN,PY]6&O)>c<7b[&S?a+/=.Q/K.7\&_VZH^ZfgY^YJ/1.(;HIaS
;_);e&^-8g^_XW6C+C@F(@;f3-J+EA)1K\[DUQ;?K\2KNB)C8A3Dc-b5/PAfR9LS
,<A(=O@O+V@Zgd^G2P=R?RP8:J]TX3/,^S)HL2.]GbQPZ-LJ_XEBgSW13+b\O25D
QTSVEVCTWQ>K?HC7aNc>\bMf=Q..6D0bTaMZC(F4+EVL6fP8BDF>@9?cT<f8RV1(
T=0/;^>\@B1,ed&-3bH>bO7fKJgX^5gd4[&=9RWEA>\+S_XYQL<W3a;)ODI?<EeK
YJC1\>47/ZMWYf\\VKb<Y<J#U.H1RZaPT=Q/LOL2X72ZHfZLfR/<?b\M6J)RO[M7
C:(0Q2=M5@VebN?T?+7&9WeY>@>KI++_KS;(3-&B)L[XOBeDe??I(/,K^L+_=\WK
)4>B=g#UA=05)@gC/<XR+_\GATE,9EFJ;G+c]N5.^WNcB\A>=8GT<N8bA3bA:82S
8SF6YMJQ0(K@:L;NQ&L61ACW.31fYT9IZ-@Y+NXD8Ze=+CLb2\P\U2J92/FQ8cdR
eOdLD4ZN&b7GP@5SE#O)(72?3fB7TD&#KQT29#W?RDXB@^f^LWG(f=\;8+)_+26D
:<IBgb[b._&<>::QGD/bQ5FX^+6V&(8Ng,c\-C4RSf:M9:T=P=\5634eR7UX62eC
,?eIbZ+J+T<B-_.]AGOdSIHVRE;>Hc51d2_,f<&(Vc^UYGHF316g[a/>..HaR?dB
B;OF(X@M;\9(@]K_Z@^DYDMXRNA91:+URWE0+b:1:ODc2Z+^c[GdI>85YYHUe)(J
L-[PV@?D0b#9M@:0[ZWA6;7FH@W^)3Q+E]1M-)+KS>YVT_YN0CcF2cEO#\^>Q(3:
Vc?IW?>ZXQ107^RY,[LJQO=25S2De[IZf:Ng<dV[J,0PC<&P>VF>]TS=df6d[-Yd
BN@MdV#ETWfD#4RbcO/JR-I17=@c/CX[\FAAaaQ>?2=#^.^XIO=^+>9&Y-Vg.=SV
-AV-gM:PR:4(_bFH2(\BFOHD5_C]LJ(6NJHUZcc\VV,O4PeUN4YT>0:B^B<I(1H5
ZN\&+7UQKH/_ZF9.M,\&3H^@-_O)9GKOF?\>&MM#6^2\@JB#+e,M+DF@]f7-Vd=U
Oe5..814>dLJ3[48>6)6C)25L0Y#]WUKdDLW6=&K539F#XY]#JHK8=fO/Z4TI,PW
X0-=cJ)eVM7V6)XaK_Kc,(?]RZ\(@#M4[F[5BPAOV68@b=SZU)bXEY6@B^_B.HPQ
eJM>3OA_9Hd2W&+U3b;dbVOJF(3E8e]1Nd-_B[3;F11(&,5>bO1@fTA#5T+MG4@,
+Q]N3)]9dfI-F+>g@Q4LL+fQ_6gg/NNS?\2[f5(QY7ZT#>RA<6O2Y6HK#ZbC&ED1
Q]X[?:ScdW(E.;04K>A@cM;/Y90=Z[4TH\FQDQ?]V8[#/YS3g]MA6f=_4]Z<)/G@
K(VKe)#IS;4^Pf/TDRd1^6D^?XUI?M46LSN=ZSg\U3A2Z@,dY1(?:@;+XA(IF)f]
EFA4f.[K&+JO&HQNF2e:4egJK7M6IeQ?FC1>TW=b9@5.a.ff=e(QYO#3DF[N?TTf
Z>5+W-2eM=SQVQ:aN>-PK:=[d7L4MA5TdT;XW30TgaTe6#-B?;OY6IVW]5.3b<&6
8K&MZ^bGU<.-3@..__M;>LAIU3_e@OUdB-I#<-WfCdB;U_15/g.D<.VEY#C=GI8[
\G>+_J9N+\W7BdTId[VOQ:3^e68YM2a3G/JDS471AU4ZSZKM?g,;b1H<#(Z04f#I
^U+KX]:eLVY2.aA_J;.:JTO,f7TMbZ?-B#J,)ODGgS6YD72V&EMD#F/,=:H9L6#T
5(;P]>d(>.g]bVKN&\#+DXO<_[#\TG@=+.U7B7#PPI6b,)0DfJZP1PDbNSgO-cZd
2@f:1-e586eC4>8EWFIJ3Jdf-[95/S16]1U+;YEfEG]^2a]gDD6J:e^];>OdcZ2J
EUS04eU?KKL33:C=T.B_2VR>PJIX8cY0-X?3@Y-2&)4TeD@f\-/MNeKZXM7gGWZ@
>8ES=S9_GRDA2#1AW(e[+X>28ZA[54#SIYS]Xc5L).2gPdJSMW^<:.V+H=BJ=dB@
CZ?L;Kb8I7_>_)Jb#)H1MC0^Y,W+O&PcOJOFbEVR[(BSeeNga@\f6M]?,EVAK>1f
QZ_=[(+RV5-PQ(_Q63,FYYgb=]Wc>b#C_/cH--1&CH^0YE?60YBPKX9@D+@\f^.e
(]:7GVYgUF.L_c/2FC2UZdH>.?6(W4LOB//(L5J\@\0QO=>I>J-5(,RcFaCG](.f
BbGVJ[0Q9afYG8C,3DTf\b[Z#L^=>BDT?V8VM4eO(+FfdeG]\.05^AGN_(dLLK^V
6F,56EQA<@BTY3bCGVL^/R>BM-?J#ZM6dEX84E=:)973]7>Cg]^@eb3NL,5.+D\=
:OL7E2X[?N6]FFfR1S/.gHHdffK<g2:ff/JTefF8]#D\EIf=9TVFOf?Wb4M9W@WF
[\HOEIUC\;,&?@KHV;2LVSaX[>)P9OPPEMHe@R_=OX/2M#7<,:2:;f]DELA3;f3D
DHS6<bP+;;JGD)OJ;JY.A:H6G0CUJ,@JHBS?Ge_>FYbWP<KE;X7SJDM^eX86-HF(
I:dO3,HSX8ZcB0d1^(L)<d4:c]BM7_)@G:P-<QK:GBE>P28.J70AP/>44cI=CRTX
_U)]cXR(&TTU#VgNY38I.Z+[0KUS_B-E@Xg(V.Jd5QGQ/S4?@GT.[9;54:)#[WA1
^H74]1F/,)KbH\P.VgSXKOeOSV)EdHgD_de4B33Hc\\NXV#eP;&4@RaGF1^B=D-J
JNWff51USE2M7O-O^DDJE:I1D=Cb:SSdJG8@1D>^2&UP@O(K,NJ3;D+I@2.DdfAJ
RbL5UPQM;&aUV;@?,dJUY=OI=BPWD)Y^g,E[:OZAd>3HdNAPa7NT#J8gT#B4P<IE
4d-b2aeG-OS:J9@IOgggREXab62JQ3UaC(MXMYbL_I#&I+b^M\;.C_CYCIT,068V
L[dgHH]ac3&.H+4eSaO5[)OI;>.PRdfFKcW\JTA.N2+,?91-O6@K3g;#TUKCNK\>
6[YIfE<B:?8TEgPX?=2V9DG>LFRf-:We7M;=I=V<cH=:/8:1YRaQWC14ZM?>IZ9T
ag\/IM/G@0W>>df+,,Gc2eM#NV;X2)/HLYRNCT32S_Y2[N>N^XU&g+K36Y,_A:L)
[.I)Z^_.D7\57fXdDS;^8X3-(gaNRFB&b2?D.-YJ[<#B4.XLC4IVfd3aUXa2-).[
I<KVYSEUDMgJg(FKQ3^77U.[U?K]P#T/Me,4KY&JHWFU1WTZ[9&^#;SUB310[^BY
8P=RXYS;QeEB@7dI8FA:FI5Ug>QgH#R8AF4Q1?=H3J)P^,CQ13QI1eE?_,#]&KHV
I)XJSf,K\7>RbNFHZ-W0/2dP,^9Kd#K)RU=VeDcaCeD8L:<F_^F0a?_JODf/UCT-
HQ/.(L6W\VegLfD=+WV_gOaZHef=6/(R?Nf3JO]RP:8MSQMaV51A;Da]/?g[24e&
XVW;RQ:M<I#2A816)fXKWU;=bJKJAG3Lb0;M;+9788+IPdP&bPYK^)KFPgO^=BT]
e106LJ4)1>aW_dXCXIeUcGcTQ>eMb[-:fT,P)N(YV8Y6?f<A(N3Lc9T^//aeL6D/
AFe+]\?](IUeH_#5B(B6H[;#XcEZ:ZH?N1F]B4YYeKA=9CMA8F#f2I?d)4?KP-:&
X4?<1T);I[JN=SZ]]0X/-e<UR0W+=4FX)&(:[KFJ[C@-WRg387W,CFFW95NOCb,[
f<a]^E_e/g:D&fU-,=F^bUgBY3Y/LaAY86?NOH1ZP/5/Q9XFT?D>FA#:IJN]6=@P
dRP._UV@1G=,18&_eBY/8I(X(_g61JP@8TfHF3;8//Y,bP<]BK+>MTSP&:_Z/5=Q
S=]T6RL,f<O#C&PP;<b9ZX]>N]c,5>6N92AGbSJ#RI(.fPUTfP6&^&X2-6O;eP=T
;AMJ<^P&>13:9Q6PHA]+S5AS2J+]7]_?LgbGYBB:V:T.AWSXZ/M3-#\)\.gGO]/>
XFB6-(LaAPG^IZG6JSF3OZP_5Q/HJPJEeOa0HLJ/RN\/_:LT;@TD(F;^)V>6YZ86
YHPQ,.aP<A.O1M>gU,@&(b(UB416SOg8@#<C1V3PRAT&#OQ8K>Rf/Zg8/A>f.Ta:
QPVJ(^34KT+6fEK47@XYP;1HRD34,ATcWZM64Q/]@+>;Z6=c)9)&UXK];Jc:I:>D
(0&CX\a)OMB);(D_:;>T07?#df^&bH]J556@(@\VdAF[CL\D[[f),fZABc)OML\_
;O5NNN/JH^<9,e+P_e/_\g]#5UL09?5]VaE-P8Y<:TRXPO0T:63fAOSF6KMIC.B0
2_Z0gQ7g+Ag_A#-,[WT#8T\.^[;Z,+5VT2T<CCOAL5N5)aZDH.g)^>66F;)8cZ-8
72/DMIT?.A1]dQGJCSF9S&(f;:W,,:(@Z7[A:+Ie>MgVbe8B@?8J#DeJ)F;I(H:a
QI+RfAKLNePZ8#(<6Y:071caONYIH#(5Pc?9[U\TV3a@Ig_D,6SL-K#^Sgd@F]6g
2E_X5X<LN;PF::6M8D\#c(b?UIB5I:bZ]fBg]4fTP/fX8?WSg2(6F]=CY]]5(WP5
f3,X8_X\=@=1.;d6E-6Q7c-bC+>aST&.)Oc1(a8JacYPXN(TN;d3N=BG-W&cN^WE
3^QO1MM&SH8-c6bLX_8-5DR#Z:AA+(6W/HCNO^M^D7J:,YQeQ(d&C=U4MS,F09<^
?6A#M8cb)a[[BVfLT^;5.eW&+)BMKgTP-XfP@/41L2aE]U2\D8/+>NOZ)=S]Z#IT
U8R44QK>PPJ[\(\eVQOO0RdeZ^VB(3U;XO+L^e=?YQ/TZUeV#-V@fR,gG1LgU#W1
IA6G6(J5HNG7Z]SIRY/):=2_0UB;e6R3Z7#EISC=dH+Z1aU)M8L4Eg/S)dE)eOVW
RX[9JZ<:@Z?I3(N>>_839_g9KA&Ie@.CF[(RS]_E)Pe/aZCF>#3e-BXR<KKH&6Y)
B2H0M[d)Z3<M6W&cK.JL7,VS:CEU3@+]VGG.Q(V&M;gC]L,)U>cg=g&Zb8@BA71Z
0#a\e-\?372(>G,UFY[/]1A9R49G]G95HLZKdM?NVd6<;/5NWVF_9)BL)=-Wbe.f
FVG<)2B##(945JTTgO@aHT0NgbE\&cJ]#92af[MV0HLYGXN8?-^/5-WMCO(ZO[/&
^1(dH_PZH-fCCI>GVV<c[V_SU\T&:8M&T.THI9Hc+,]&:>05^+Ec>BBF7M<^>W7W
]AJE9+@a3,SScFbNY&gXFc@_6.[YO?W6^K1[S(3OdONDE49,VfW?,8Zb&bE.gT,C
/N&@M[=>?H<7HF_=J8DI+YfD1.6_^L52)^&]=)^\F>AV\KA+Xf;[G(eD,C5QJ[3;
4gc7-:Z\b-T^=^J;OaIILe7fJ5Z]D.[YGY2Z.?.HV;AM_=F@]R#->ZH(GLDF3@C;
JQ/OBFd.EOPGOH_Vfd?0>3\3TG#N5>U)4/J;[=4Cd.100[)]X7\_Z(41A[.9,a7b
^>5cf;MDE9H0Z&6J-dd<3]5[BGg]gL&L8,2cYRHW67X71W.I4?6:8U&//5fK06V\
8g_K&X5_e+Q2FOF+0faA8\#O5.J3B5egM])?:RES[)HKDe7^1F>/YCHJD9XgX88g
VSCK.N63NTL_0eBXd>KO:X&XQ_QM/O,,-26,([aGY#gddaY[NHA&d0XQY,]J+R#Q
Z]B/f09\@,;VfU(^ET2+SaQgWJ6?IA2FNKIX77a?5B#9d(S]).H-+>WT_&8278;5
0@b1;)^b@FV>=LZW([4O;+AU&I?AH4^1.5:4PXCDJ9K@/aKUV5&L/1;R_L+#F]Eg
>8#0)c0.;AC8H_NdfD_[d<a14393<Ec3aICY4OXD]SM^_ZIfB=)O<=H@^?H.IY7M
V:3HM:YdY8NC1B6cC16N4RD3g8bGd3V^:Dfd&TPYSMYYQGSQ^FIN))<5(YJBc9FC
ecdgQ.>C_H)O02,P1X]F_H)dd\OYT#(MZc;Y5WX(AMOd?/E5OJ75F&;;[/P9b&;e
FML:T#^UEB2e6K9d.>LXAM-.NM)I9U;c35TbDE(fP+Q]7RQ.^V57T^)P1V7><?6f
2;(4G1&-H--A,^Cb1790_B(?LeE2RTZ1[:+J0.XPH0#3<@N8[]\&Yed0<KWQ)MNb
C^gC@BO=:COBd_1TKQPL_(e?5>]?^U[I]X8(18)OAa2VHND9M51H2Qg39dNJ<+D-
)FVD4gQ&a^VONaf@Jd\,[Of?XTQQNE^K0fEINDXFXbc\8)bJDDI.cgWCfG6N\Z(d
[=eJJ7IOZ\2ED:;E)BGOS_<ZI1=>cI17&_(#CL\0]8fWb1Y9/EM7;aJ>)R0Y1.P7
5-@YH5Z9/?Xe6NIJbe141b=4>F^]]H.F^bX);cWZJ.8O9-aCA59RMcI\=a-0L8VF
>YSS:b)Z7__f_;fS1-0]]R[+&LRG[#ACC,YQGUYX-IN2J[H12#L[1b\+<4;_)KZa
,T9I?I\V=@VU<HdH>).3J\>#f;I;[BYNDK9.4:JG(:V6VE@LBDK1aEe;;S)f(.4e
g>M/f3L@4K.3&(HZ;YLHY(fNG7B;)1=^),Z\+T64ZHg;>R[]?QQ[,.643f?-WP1:
TgeUUdG666KI^(#aFO7QMa9S/935a#-JLLU]Y30g]SW(X;AE]b0Y1U8Z/87L2L?>
.@R44X4gQFXf1bb^E<V7M,J#2=7YcQV3>bgR<S0(]2K5)dJ4I?Kc4(S(9-N#>H^J
6M)BCU)VJ4fa8a6D)W7EFE<3F_@5R5Y1W[S1(:7-6IG]5J8-#9FJ<S7\;aQVVC#5
M(L?fUe)KO+8\H5dQM7-f@R,,FM);+&?9De<J._#+86(W#QMaA,=]Qc,L]85_RKN
CT9<B[TeT8aR,O^a@c&;c),P3TI(-FE#=Y;gdg/FfC[a52GA85Kf@O4d:G_<7OSQ
:1LXZ<#Q;N3^(L=2G&79DY[78C:OM[C7D)I[K&a5Fe[6.Ub^.V46S[WM=^bQH,1(
C^ADc9EDK1-QO&ZfXeg3ZWO_DBB?X_?OEDS_]0D_PJ#E//M+O=a5@SSX0(B;])@]
BT)];XK3bO/8&L,<4)40WJE[F,EUB)Q^YA/I;a[\G_5>^(A([HWa_?]P[+V,\3-R
SXF&P-/LY1C5&Pg7^dBD4WR1M[H;R3(92P=4=I6>PeC8b1UbU6NZKS\2GSKFf-.L
NEM.c90aF8@SM^DV)9J5S;VDU;ONGZ2TH6W7^f1X#gacgO;/e<aE\70[0)(?Q:N6
,+C;FE>[02c838g289A]XCY]YUXC1P?D#G[8gT;&Y?ObFZAM00_0MCYVdIc.3(c/
KW+6X0EHS/\AU[:K+OcRN-<[dS8+S5CH865(fE>>@=)(9Kdd/;<4^-fgaK17WOCD
<N;e:g-U-ab^F=O&]aP:S)[-R@6GU1dZ/fRc#QT0]0eNW^@M.^:619<Q;6aF5OIS
YgEf^MRZ7GdU^D(a&Z7][S^,bQZT2MK1?#1X[^[UV@WgK>S#<6F#IWIBTa(;HM13
ESc_),(5\+AI/IF;Q9N7_f=_U8aFYY5:IR+KC=?22e3Y)9D5a14,UGC6_(BPUb)2
IKJGCV?T@EHMU8G6<1NWaf-@-U02IVgCZDfaBLH)]WDbc/?09LICb,S_S:b=,I\T
Y6&e:0K/He>O;QP@dAb[C=NP<1&11LLA&0.HbG=-gJ\a7J2=64:,(X1-XNAgb=&@
^#&=_@+4Y+YH?EGdXHQ3+0bg&./<b.f^5aF9bF6C,d.NYMdG[VO@16OKP./O+T+Q
L,8,IE_G@DU:Q8MI+,6B:CHX+VRMO?,@B,>>\F+D<Le[(JNX7W:c2_4Z224b>3F;
RR:6U^L4bBd#3+;N8C1[SZFQ+_77BBAW2BgRf#U]@0R5K2L_4c?1=>@/R6E=KgRP
U7#eCXT9;TWU47I46A0I66^]X#D:4:R-FRX91U?,GPM=FaU+fMW3B=0b59]=aJF]
b[R)dD6&b?1b-L\]B-5bD3#E8)bWRFDS=U[L+Z&UX^=N[7GO#CIceYc.>e=3&+DA
\GMFe69dEJGB&E#I_Ac^@9_Z;Z<&_1+571BbIOM@[28#+F^6-GE25&X-18;b/:&_
b[QOa1KV[@Y@8NY02<1TNLD_9fZU:ADE\;fXM]S6^UVH0-3>;>E;(J]TJT1963);
#BC..T?Cc>LT2EGC,8W.a[:-LVDUN12\L.I+<6?II=KJ@Te.AHL^U>0BDX^6^?=K
_VNJ<A-,bCPK59W2+N0d&1CgFT?e(T=#)S7@=5U?SC&Z6U.:U4SSQS^4D\F5W([J
RQ5V1:Z]C\L?A]e8PHCC,K&JM]M.6V\gMM8DXe0JPO31c)@=-dVbZZ@2>68B[=2b
fE7;f&SCIC;5KNEeTcb,8BRfI^;CZ;0K&C1=DJDCNEXI.EEaD)YE1\-gX3UKZG94
]&.26F91]:6J#X;KD;XG<X&;MK0g.S556PP4:RFPIW[VKb-DKP6;^-6BJ>4AeLd6
)PXe(H&cPD-cZWU:Cg1dCH<,=K6KA\;>2f#]TRTBD3[#_VcR^6,Q<4;e,Ie:LHb&
:A6O.&D6<^KC(\T+)[09S&W8CMJ.X_#a+_?QILF],V;7F7Z81U2.#=2CacfZCCI4
5A1H\RGD>4,#YGZFf?ZPKU-TU^F2RMZ1-fR+#.X>_46X:)GN5>Gd=VbD[J9/O1=V
>AX@?,Q@GMaBS8AV0d6QY_))6<YQR,[NeI1:]O4N<[bCCg_A/VdSYXU6Mb0O@)5d
=EK@D11<27#=Eab05CNTPK;BHAc2C-I>Nc:?U,HQd,LAJd(KX58#JH[[,YMP(A#R
4X.@N/eFDd1R_ZgL&M5&@N7&+0AFZECaL8K[M;gaK,.CHWJT@c-6E;^FT^YNBIe1
@HQFGFFRS2Z48T/]@1bR[]dbRF4EYB?[U/Hfb@@I>#1T-SOa:6GGB1U,fL;:DCF5
&<B;QY4>N>FJ/\3-8K-[)2fSC,\\FAdad[b\0g=dP4ZIAMS&dG6X(K-7CcSX,V7G
-cY.(GCXe1B\03_FD;6/+_c9edF\;UeYMD^^Tb.AZ&f=<aFa,8L@D7^&11>UadeS
gUOG/WZ8^_5a9fKf\-GZD9+68E36--0P+XV:?UFAQb,)/U2R:&TKN&.#NR8]d+;1
W5@?2?YT=>_dA/4_&HO4?BefEXX1ccc-U&d(bE=a6?]c&KF)/V6JGH3JE(SB4@AC
[G,-36=Y<e3gD13XZUGWI5b,&S.SDfOUB[Y/ATUO4\7#agR^<<?\JYMXOZ;+Lc3E
MEWJ?#@,4G^5\3Y,DVW?3?FN^9Y/E,g3Gbd63-_FE2O#T(e8&@TT@QRWKa1PRg;;
Kf\J36K=]K]D-U5<BK6g.TXDVA7#8?NU-#:]F-4E;[0YSaEF^0RC-^\]2gcH&]K&
Ie2:2PD52aC[?3gUaa6#E?bH>GaS-HFg(^_fK6ZJT;:;Q<?gf=1@(0c8b[Og)9,L
5b,ZFE&80NWB7=:]<?+2fZ2KE+_M?TABA6]E78Pc0UKgR@^Ka_[aEZ-7(HSF;A\M
/ET#0ATcP1O>N-Y2F=X[Y>.W96GfZ>-&7b,M\^AI97gKTZI-L[;&M^NJ:QQ[:Q7:
JMggPU/J=?I?DU];C[/?4U/RPHO,KBfegd<&YJ(/^EcdB0(A\YI>2dB\&@Ob/MU,
6f5&34G/Q9?D)2#6HQ=#8_-UC1f4#;986YY:X#REeWY2-6;&),,aJVZZcKA5U.QF
U](MF\f2F;CP^edBR=[@N&8/.KYMc(aXX=8aAg=I3c&N35,)OgEE3C3\<I2Q,6e2
1,La64S/L3=N9GGgT/TX0,]@gH60-GPF^-\&2UC=VMeLPA?ff6IdN6,aWD^0b\e@
.DCBbCH+a=Ca0LN(.<5J5&7_E=TL]U>N8PXOPNN5\R4P=G(bD:CI_#P]d)S[T?TT
eA##AGA70/8NQ),aRg3XR?,,L>Q2+:[6A,4:=DI=>4/K2JL;.P\S[M6-:D_6]O&_
PPEDge,bUTPDS8Pa-@,LJ9^F0X9@^bU6[G]T&I,\5#718(eDLS7I?<63gQ2Z>F.D
94fd\Q(/RC+g=cW><b33OgX@dR>;:<RQ0&Z]9.3aLgRg?2PU_MLT[>=U/YR@XEcT
gN_:;O3[d0^8O3ac6,YOG+3GPDNf(DacSKJP]1c\S.E>-,-3aG9-M392?O8[ZMUE
S089]+-QC&U>>GA8aFD/Y56R#H.=>RXQ&);;&WV@;OH05?HC,TKI4T#PYVGdPU1K
Z^8.<;S1F#1>Ma#E?LYed@E3C8<W1S:9G42U,(LfT)11[YD_J.\.)8XE7XTDY9H4
.9FJK4X]Z/,YIN.DOGQYAZ-c#3b)MU=[12C)2-8La@/MB+JZd+OgB<6HCWAb@,O0
M+J@6<<QBCK>DdYDF\SSTgdBF1ACVTc,N<&N;10QR)<N3X)9L?OEPE]&f^acNKFd
cH-\QLg+4WUb2UO-g:5<.N+\2AD,Y<M3B6QQPM-&ZaB73[-L5=\NVA\LT>B(dL]C
+<(]&VZ.N8HCZACfT_]IdES=52/#-c9IJDR>.FN(HL&BDADIG&;1:IbM@@@Q[[19
N[-]gH/[8;\Z;#WN)=8/E>+N:4NCLER/LI5@H6V<7d:bX:[Y>^CF;=)31)]CZN\5
HW#KDRXdHP/6,+QY.VD8SaY)2cXc/PZVNFgH@R,aPDdVCDeS#S93c:OMS3Y[EN(V
]K&2Be7.N#]fJBZQ+\ffR.0c1H2[Wb1LOOT<WcK.&URK^)#MB9^HFXbA)V6Q&>VZ
:42QC6\M-/HXQXZCGH+_Y/H\M;H=b-NK8&X/#EfC=6V^:^J&UNV[Y#gT\+OY61#a
a5Q^8&I\E/H8b3(YQ.#).DA8EKVH@b_]Q4T,C(JM<F)?XKV0g@aC=P9F7f;9TQOK
eV@26-4[/N7DQC\Fac;4MeU0[Y4TcgbTf8ZDM\Xg.1d[TU\HXbQ]Oc4:_fY@G:Eg
:&(ccM_bLJ;A/ab<QgbKSFcOC.aU0C<4354d<GHa9a>W3IV.431[Q@<6\0OSD0AV
N9);7XCBX:e),dL1IH/4XQKH8;bT8_@gD9OH.dY4(=\?QTF<]<9<6;AVE-dB9\SH
P,ECW,]C\]]TRJX;W>YGO-,COF0QQe+16SKcbZdeN6F?1D?:dDO5gE&JZ>(D<SJ]
9KH9?0N)K,EW/TH^5OGPa)MD&1/.CBHg)X=76;8Q0&LYVc#/@AbR.[0g490L9:#M
Y8fSO(.dS/8V<IObf\D?P@4)6[bc:37K-:+CJNeSfZHK1cZeND,DL>LOeM[&>cB)
?b2,,D:4.D5YaRB0SUDgXQB4F8S8N#KAIcgT9L//MPTC?OUO;(7PU#V]OdQN&]<-
]&0\_bL3bb)RL[=F,bOaX],1ES^O-QC0:1()]T+HR2+Y-7IOM#WgbX+QTUg<>X3V
G@;9=7GVMIR=a64>TeB0Q4YQZ?TJ(E0(\R)POSV)=-b10IP4?gQZ[f0NL@8KTA11
??FQFf6R_A;1HC:d\LA/eTRH<7T6>adTOeb[78FW0:XZG/B#U/#8PdSZ9S-)4>XO
AU8V?&)MY4,^D(N<4_E0b><TRgVI+KgE.XZ=RU/^0N_]_7PeZ(KHab8f_J?cC56S
=>Q?f@MX^fb&d2_OURD(NJZ2.aK-gH@Zdf5#7Db\^JMO]Kgg5I=OPdO&+9C7SRT=
7KR@c6URMPM+B.=@C695,^9b#)N9>950/aM(=(3S\<J:.4.29->D4HQF-T75B(2I
\gYBDR-LA+d>,P]fe4a;)/R;R834P\I?AAgZgRc=9BR_DN=\0-LJ0CO4<R=]WbcZ
W3QFA-B=T_LC\>1N[(0CHaAR+)eN4S)8,[aUFecKa/5(fI(^_\K\=OD5B76;g,Nc
@E_1E@1HW>FZ<K5T^KS218KDc+QSa#HZU\=I)5\[[,1[[3;X8QCe<PF:_5M#Na#@
,^b=aYOf]7XUc]CDMb;H@JH&)IV7#^VL@B9:Y6&c28?)c@FO>LQPA/P40VACg4>=
bcQg@:V4e&d#4OTbHX/6T5NKb1(HLQ3,QPg0-9Q7;-RL>ZK:.I]W.OEdVSLUBL]H
WHO8QXf7)</97F&DCb_Z&e7F0a(fA<b8gFYTf&KVFJ=?909/E^\FN&3(L/gQ06C^
IJ7CK5)?OHd:cGR_gJN4W1L1^fS>2gT=/9>NJY_]K8FcJD_0>5e<SX=I7((Pf6G/
B_8U#Ue;#OEXF+H7L@g>+daeI^^[V(a)gSH3^/F//=W[IH(B?dE7_IJ?afV76dBC
OQ9=>cX@7]gB>9/8a)FY5X4R<CB<1_>@ZDUF4=Z[:-\40,#_?8@g[0=Ab?KSJba:
I&M>^3CP32METGI/UCDGa5cE:O:]8D&397HCE84P2O#dPeB^A^SG\_E>GIJdWCX,
[D#)OL;J,OK#@I^baFc/2F>Ddb.:C1U(aB-X-0,JZFe:].f_D)DR&NNFCS)fYVeD
KcafA4Da=/g\Uf<Yca&Y^N:_BJ[Y0e62f1IL?:FB+W.X<d.-(gSN?:e_D<Ea1ELP
e#30;[_5K,FRBY9L(63^W,/4f#&a2DIC&E02^J5\\b>/2.M5A&8fX:+U?.;9P1[X
cCQ<-MN:TWY+JXU,Zb6>&#^CP[724.Ac<E[F\ZPdb?GH9:HeQd0;EA4Q8P,B:FK?
/-(aNdLTVUZ=5GU(,SBcH&9(QTH#:ARQ,17ETdS(1<O8aTDJT/[?6YF4CG&4-D@c
/d<5K?PV4[(:ebedb\g/Q<(\\aDXb_YR#f9;3g-c-[W#(g[@EL\5f4ZWBSUbc:.X
adA1CWg[7+H)0;CCU@<[K@[VaG<6>J(&3/ET21>>#XW+R#_dYM?Y-HS;:)(IZH>I
9=HXZP3&P:ZPF/8GK5AA0b5)I),ZEO5]-Q#BYeIFG6\,_D-9LeE\U=c8bCR^)gIB
;b:3f=VI?gR1HeF6@H9U2cC+e>[8Y:a5^L#c3Z\[U(WX6&+<Db&R@J(Pa9BVW1F)
(Z>W8\,MRGTIc@-6-MN;]C&NMEZS,V\7MfN(BdXP?.V34H+K5;7#Na5E;^GDbLJQ
\cTH]:ZA6>D?.R,HW?-c5(gDeGCEY.PU/5-Z9BW,bZWe3+E<@L7S\JF\gU=^>OYG
X6g,JT^c]a[6G/;7O&Od7D.L[I=dJc7F_U2DNL\@Y@_WY#]c[HZ(PFScY-5V7@ad
AZ9O24A4bQ:YH=8^N@:>/IaL;?BHRgQ#X8IPNT0C]S,HeE?FF=-cGIB1TUX98.35
Z,^SGL<;#3\1>LLTUKc6,bINSV0YJ6(+UXe^U]<VY[<HVL[5gFGcDQXYT<;(I1,H
MINfNbU<E;[JcJ^SJ^&fRT?G#DG5GK/7M:AV+V2LWD_;V?49.N_e\fT8W<)2;L2\
=e]OL4bV2NeTFF9b/BDE?[OdS94DBcV(<B&bW>(FW&TF1cZS.cLF]CE(#eZ4U+A1
.^gCG=];]R#+B@84K]HeEJ)^B<[KIEd8&BUZX2JRP[8feV6AQ])Z(TH/e&LR9^\/
[WU?eJ?,T6f<OLVOPX&I#:]E@WBBHDdAXfVdXdeS.=4/>T(#DUA#7(SF2ETg-6.b
\G)O263P,>f<^aCOSV.d80IR^^e\7I[5c4-&#>0Q3V1R@bU_@=bc[1KY2ET?]W7I
GCR/7b2#e\?L<Z>-EbNCQ3_SEd9C-\NZ?a.X:7ZJ(\cDVSCKRc@/XKBZ:<5W0)WX
Jg+Q584De,D6-e-9D3&C2d](^7L/(Q\?@4Le(+_-f1OIgR.,76_G63OL\T+IB0XJ
Q(dPYOaF#Z)ZSS)6f:)V9?3DF>3SX;=I@JJ9ATI=aC5&c=[2g;_V#QI[J/Q]IRDA
JNR,14P8/4GaP,&1=?N&[9:0O,S-^<=<9d=9S;<,+06#&efc>PA&g\)d-(UHQ692
MKJ&)aVb)W2E#VVT>DL=E:5O6c3&(YBY@4JDJ4=05:S[6/\g(W&K^a_&>NUA3O=9
5=+.EH)_8IO_P(d25\,,;.W\O,Ac&O>R^5^GZ0Id?e)0a6K]HZd)@&>,1=&UDe>_
Q8JF)BW:RGPQdaeYTNaH\(9U+&FCD2H7NFYU61:)LbgCW2.6-5X\-)E+?D?HgECD
-(5T[=gVO5?-2L.7/AaC=>G)e6B[K[FRMV8QY]1dFJ(cK>&[<=A;EbfCb/)8B^X&
:d.dDJd4Q^LWUL0O;gG+eT)86T81f(O\8C1K,M?)-W^Y;(R63Gd0_[Gg@[H4XD^A
NV69D1?dQLJT>aXTL.H=0V^6K.56^\[5>\J<XE:0f#CWfgC+5^72fV)::Ge1F_gG
1D^KM?32M3e55YKTNOV_(bM,CfK^1_((]dZA-@1;?(/-E+&2CZ0Q[U9&GIae49(2
?,A2aY<?e-@2GWIK:B)6@X@/_b58X.a/I2N)=CB)Ue^W@9>/R6bc#f7(dNU)[8gV
.+[RX_[PR\QBZB-K2,C_CU/g)<RMe^1:g&O51F7F0/9V&>I&F[K85C.+Q.:PS4?T
]W(0VH9UK2NQ,,eR>ASY?+-F^cLOKQN+Kf?MAB:,@,,SJKOG9#.>],13f7Q0:VdX
eP].WW\GZA29C5<+>]7=JN+0<DSYET4VIE6QB>Oa(>#@YCBN\/_eG&,KKQ_;cf6P
<DQ):?PW2WRM435,[WQP)PAK>(7LOKXbHZ[8OC94A\4F:J(-<a<^3YKNBec8/=(>
bKCa=0Xc+-RZb;aY.EH>B)efO3P_6FRV2P[V_63^0EP?32J])^R(^6C2d]bYCI9]
(GZ?@WLa(cQ?,1IV1Y0]=)R004L#7)2PWU\W59+<WS#gCA(0PK)c>JWUBLH[QfQD
g-HRcc#6L]5QH@(665_=XZaeW-Wce7RJMc9/F&GKXSH:3IM&=0e\:CO84Q+0NOQ-
5H,)MCdB8ZgKX,V@0>JS=T9-SXfE=XN>C,PL.PE=9,9#8C0a-36aKdOOP4;;Pb_D
8#D#P,DK1L]?,8Ud]/[[f62d/UC8,/>7OGS6TOLVg(6Ha=+b]Jb;(Cab&b^(PU=(
f\MLDeS0>N]?dJQIFVHag\044[E8Cf#/<]@JTQaE>d4GfL9\TTHQ==6RG80)+0T)
R(=.#d?W)eH4OD8:=XaN63..3\U\e;X.e.:c)J[PI=b6[C5[I@1bF;^V.9H<WBAg
5._CD.4SZS_5JKAFGJ;V]H9NQ#[RA3ZaM7(#5=VT>[N1=HUW0d#WOaDJYf&HO-I?
.PM(eVAb?OJ^L.8V.D,L0MS(>LOeNIK#Q<2a\8Yb&?NJ=6>JS8W9O.QM]AMLbP39
;KTW9d@B6\LcEH.1WYHBXc1c4+UJ3gU8+cTWR_ULN?>b>@4,#<Mb>FGQgbGOR&3Q
:NYXTME1?8A)&cR&TeZf4C>,-NFUX5e<KAJ2aaHWZ94]K1N#]9A^5M)+3<X?Y.<U
R-NXcdH-OT?V>_\TELG-,J5-;\6dV)<_d<2d@KKYdS(U_8F/M7;XKN/c9e#-LZ\4
7H9I(AEZ+_>D,L?O>]d,&+g?+10O1S&e@IFS8DT#NKYG+QD7[a&PHWE<=55&U795
f?56:AEHA]VJ.R901-]19gc-/:1],Tb?V;c#f10\AA&)X/)2XD(a3\e9B-F@1(-P
@Oe>N@5:(L.4gIL7A4<Be0C6T@B7<:R0L/C8d8[BgRF+/ea._4_7d41O4@(O?5OO
Q0ba[I;6HQcFF3=<]W6P_10[S)/X?SV2V]Wb&(4#)YS>P30>Q(([1XA2GR&Y]&5N
OTDY:O&IINbSIaQ-\\\0\V3&7J8V]Q8\V_QZ<_@B>bSMS8eA#OPC4UU&#T#=9]Q3
/\.10cDX0g1KdN+HGQI7D??7FAH?IQ<=FAOH7M/b;V4PBZfI_:F7??Mf6R56EG^_
:01SME7eQCU^(DF^Y>Cf.:E50&\ccB8U>Ca6/[G=PE3?DHU99XM_]ZP+;[TW8;TF
K:4/Y[eb.0Na=ZO/]]((;J#I[SR816:0EBUdgeOGW+<gfO<\KIS36ff1+B#/CE9@
#e#_gD_^5UNJ&]b6>VABE#]FA^ffJ.ef;Hf=?-g-e8^WUCGNaAS2/,JEec;0(6X@
(X6eSW,-\b/2LDLSeAH83WM)cWQ?&Q^WH.&IFY>@W6(7&-be]bb#8D+\eS)X6c18
[822Vd652N>cKEfg0XP&a<:D;P+72gA6dB>.VJ?4SD.@V)0>\C,=?f-D-@R87A73
H@(N=>M80(/#@e,6^Jdd32JQUH+](JENg^))8:;XS5Jd2=4g2=\_GRBeeO7E)3MU
bf^UUAC+J4F67E(^-FT:?E=;ZPY?AQ>?^WM>&+/dSdWIT(?^,#GQH(a70#-,Rg29
2Qf7)0&NK5O^EGe<PI70;5,TDCeX5cdF??EHgR6TG@dK)R\IYAHNJgf(Me&:.2KT
HQ:O&UU;cO&+RKE?-KG\g__K\TQQdWV4IH_XgA+&U#f>ZZ+#G;Re\Z1=E6_)4)W\
OHX:;0[7A[9d;fQH5PWLA?(5N4Df-#9DegAdMHcM-C<f1Eb1Z,D=-Z=^g^31Q-;[
?=70N;U[O>RD+P5T1D=_CT=31Y3\<^da-EZ,8JLe1?ZG#9f[@<Yca8E8f<\(66>#
J@dAdS)+X6_+GB6We1S8#aO&Z4/)IXaQI<W=Q;c[WW/Y?\N]d:9Fg0@XA\Y\S(4C
A0J+R5X-5@SEHV]YbFK>AX(5D<J\eU>D+J56A;ga(,8X?3O^C<b])+,E29gOfO^K
c&9H+V31DbLT@P/L>eT_=>:C8AeQ,_TA(RDBVY2XQ)W,>ZVS;XA.UQ;_[0S&G;4O
W9+.[d/&2_N/&>Q7GNZ_TZcDWaZYY+]O@ATH(\F)[ZBMR,AA=5P.-]L2Kc)C7=^,
GcTYEABU-\U=4FNIWX[dUE6_8^OQTF7S2F)?bMLe4gg)cE9RAFLBX8&ZQ^#N=P^&
ULV<)[IM;V_fOF^WaH0:.EUPSJOR)/L.I3>O56:,7=MIQDa&H#1HO4BW7M6GM/M:
YY]g0e986[c7>Rca;P1@)S0:[>#WCJFEa[]g.ZPQSOfD]Y_/<?eH41[WA-[+d^;J
-]If6L@NP:a:JSFdW]_LX3-FbMbaL_0_Fc:OQ3BJ[DPJRI7E7(W&CbJ9OU=I8a5&
c;S=([@YMGc/W5H0-CW)&U?Lc5f4Bf_>JRRa,M_9+0cf[V-0K?.A4T3VeF.c9D+d
2Ng]Kd&:fJ?c;8/HNPWW@cL3F/T#,_2c3@aGX/&/a]aB:>P+9S4<c0=0/R1Q5Q/e
Y5-T07^]Rdb]2MHUe;g0YA-Y(3E#=/Nf<6<^I.cMW,IK\1\X,.L/,K4W9@Zg,I4,
4?O61IM[-VY7.)KMOHZa#QJ81.Zf58L685MQZ.f/GJI;?8=Pba;B\TKeXPD^?;X;
=A4082^+Y#Sd:P(80dLMI;a@.3b1&&&^@PI[aaCcLU0B>?dYc6R\e#=b]M,55dJM
cSC65H25C2=@KHD.FTb-6G)XF5]f<WFb68X@NZ@Ae4.86#;YbK7KB#7+8fU#2)-&
I3KbJQ\\/5M4A:G?Vd4_T:X#JbZX&0/DDgSb(8+bec8:#-8@-Z+a076WX<L1&JL[
@VF6F,AT.D;aDU<BH9-?W<AE&(Ce-Ge1g+UP?]&VU7EOC.I==XY\f/+C,FLG:F;H
0JeHebT=Pf18EfZfMZ.0P0d8D8J^/VdLWRc</)gB<[KgPN<<#,Y9aQEAXO;P_[5>
)?VIeZ-3;((0SZbcE9#@#WQa@N<-d(?5gUG=,^)3\H7ee-N\>@DFQ8810P]8.d][
Q[5a?#f,>BCC][FHP6Q2O(d]1a>_=4)G.Q2b<XTZ^Pb-YJ8W[^K99T2C?\NL5UHD
2BT(:7INe7ZX0\;(^LPF)f\I4][<E-DC_M;Z?3CJH<fEF9L5+@EG;34UF?@/&N.Z
_7(-Xd0;\/cZb\e0FI.>8S@B8N,\5NI4a>X?>+O=,;KU8^;OWUbZ>^:4,#;XV7IG
BXeDADGf.8^-0G),dB?CMP:CZW8XbRR.R]2?OW8.QY4FeYOE82WM472U:CK2F?61
#&5(cJ+.c]P^c.:PWX5g+:L_G6(Z>(ZW9##_^:E=FB,4ZVV3,E]-JO65+BKJBaB+
Gc.=WBI8dG7GM^RZE=eT=aAFW5X(,0B+a=YQ3RI]C,AX<fYfY7-IAMOUaTU-&<fL
8[?^fG.WBGPfF;208d)bR^).Y,WW9b-^_2g1/14X_X0:F0bI-J-/ZWdBHTQ=T2,S
#U\Q)eP<D[V<3KBa)3A(XCaU&IQHE>4X#f7FSXIG#9)LS3<6NV32]6S1?SPQ)KJD
W,_FWX8K6^Mc9XEMDaW87\8<,5BYF+f/#Gff3)6T:eZO@gdZN)V:H:LW9dO+YK+)
[0_:A&<ST<WDYOT;[FbTFVY9bYAb975cI/d)&W7(c6&dS0N9WYVG5RHD(FO(^2.I
Y?^(N>Cd&/QH1@NY9fXNL?<WBgP?,/(#Uc&HeQ<.aBHXURZ?G3,ccT/Fg2HJcgW\
7XQ2B]IU5V9:6,g+2^:<W:[UP-5^a<S-J]\?FZ\(X3VE2(<E?eV):/f=WX]g^)V>
1FQbTb(BBD\b,#Ta#I.,bVT,d/SH?T_>R<V&3:bZ7N;[R)+FUgf\8DMP:H:[;beJ
1A[+WC/T3<6Uc#^YRIHD;f>#<KGdMC9SaC/S,9eA>+<P8fN.0f)]caQL,,]A+QaX
MX8Wd9TZE,Q/PeS(B[K@dgV@YF2;/02aIQ<f.1)&0BYDF1NTX7W>/W_H8PHX4_[&
V^B:+B9HgS]eCHVfN<JbA.FefV]Y,S\L-aZ=Q2CPRF8:2c5^V^<UOGC/Xg,eHUYD
PMDL0b.bF:WXY(0):Y9^6JN\=RPK/&@QZ4c7ba3\,cea,J)W:L,/AW2E(5-UKFU]
R=0MOU2[e6aY@,+)BcTZ0>W6fH5/][>3FKYcL0:[;G=BIG0)>;RPGIL),4EE/423
^:\#BgeDa,AP)bJW(_[(T)Z2PFT++\O-95211d;8#S\V9.&^f_75d9C(IUA=)C-D
PeBFT]]:#+gKf&Yb,-<Yb<3:^a,?3Kd&+E#>\+Ie_Z^LAf7)H3GMWb23R:B7_+#T
f_F/Pf][HO_+Tg^@:UXcDE8LLN;:WOB&E+)4/NabG4XRM8#aL,UN[-Tb(&]P(5U2
::G)(1Gf001RNM0\dBf7_22^LITXfc,1B?C2M516Za=&-0Q]/-cdPC\UP&B/4#Ae
R#QBb)4<dW]]=cgYYU,8>6F#Y&G(TWD.0WI81G(V6KR?O:^SZQ/cJaJB/eSWa>@:
H30.AH/<37Rd[+NXC/\\MCb0PV]HTHQb7a&V-,K3SM>=1H\3FF^I.;.^-RS]O:Va
fAQEc]&UV9:B:BA7P<Y]VEW&>P?)UI:e\YJ6V+OYb5<M5CS5+4).BZ^^2_)G,JeS
;e9#..Z]@R_?,4@A[>6JbEWg=+be@g<V1[6B6A&f0bOb[eH07A_-[C5,^J.>EK,5
LS^G>>V+Hg?e]MMBd4)Y@VN2[@[60fXg/-@)CVUBW2QdYI,f<(X5,UUb9eNWCY.,
H)]LVQ,W1--F.A7V3IH-PD(++2Hb3.#;[/\;XOKLF+SD90(,A[_[1/g;CdT7_f5T
5QZUaRLZ?E#ZOH8(8X<#dD=fd?JcGG,bNQO5eabC428&K,J]a/@S;a5,D(5g.#<c
EP\?-ZY>5D1Z;&T[5@8;G4BPF-I/QZ;bUGTdJEVON^;+;V6IM?]7d_e)VG&Y/IOe
T,W15XYMI_O.;1/I[_Yf^C([U]B8L5NQE\6f6XGPVV)Ra04.H&)=OU[N@?b_Gb.A
.SSHMdIJ7[6MZ;IDYS<d\X=YU>7IF24SJ\]E7QH+cD-[-.^3-IgOX+QfLQ3Ad1<Z
aLWAHY:4MZ\<U&@fR3D=NeBC\TJR-B8-fSOQF9Q9>c;Sb@(3#REKWg?#MRU?81KR
/_PWb)B>;Wc5I2_bXHb<#EfK-EfVd1VK[@&G?RW-5QV_9][0I[9RM4:QWH71a55V
9eY7X=-^.Ub4M/NWbCB?2IJ-XU<7gg>MFB8D]1e;I]@7QL7aH<9YC<@;6V=+O&3^
MbUB<)2Yb;[>;ITJV[8da;-1_;Z7+#&Q.]T2Dab5PV(PE2W5\N=GK)a50WP.f(Z9
EQC_</[[(60@X]FS>-YcWd;B6cP<Q.Q.Z[F)eRVH/34e30Z0I]SW]UIE]3S]ET(N
?I?0H)YdQQJf=@I2R8/Q0d&DgYJX@CG5^^NAZGK2;F_7U/7@I=DU+JSAWZL2IW;<
]F<cc9FOE->Z<YDIJ(0I3LAZ\A\0TX^>NLI,HTQ#M5(.A&U8eLOYbYUD)ZZ3&L(Y
\7#<Y?V(;#(JW^1SU^Ge:?Q__HI7HZ55OZ\3a&DTVX>QR0a-KMP:&_[T/](_:Zeb
R#b8N\H1f-PIUeXY-g<JJ4dI8LX;SAC8G@\I,8&K?V7(K5=K03f4I3O9Q=Y?SaJ.
T:B.]H8Ae5>9YH=U7</R2-GeBL91BY+\I<R2&^2O(M@8C6:aRe>g=cDF8DUJ>HZ+
.X#XTe5K.MD87MUG91\2E^>#.72_/R6V#E]1SAKM-QSCR-Ba@T?4A;QY+eM#TCXf
P6[aV;\c<_13g2=@#eW-E4ZH59Bf1]QIB/b1&LR(b#dH,I[&O.gHJce.W],YRF?0
BNF?-0JTL-9>aOUTL]=E0:/:+Q;/c[-eW8d[M-a@OG@HU+^_K7Yf#,5TVCIHPZf^
d=U8cPSYD.K-8RI;KDA1]A9]Kg]JYc_LQdeg\OWG[YA=>Pb_:OG&L88([=+M>bB[
0EFE;@@-I.P8H<7OTNJeBZKU)G/68-5a1/(MVHTa07c_,&X6<Ha>5_OVIU;@8CZ_
eGK.feX#L[^\^0NC78<OA9YcW.?UL2\7R\[,YO3A:LMT(S^9+LP:cY^5K.T>]S(L
C]QHXdGN-@OB>#3XO]0c0bc<cHFa3(:1c5C7^[bJR/Fe2N8KIDMR1fB\Q_@3,2]b
Z/LR?5dHf.eFdQ_7BJC40Ab=P7U]&4OPXXCA;@ULLOP9T9\H3X2Jaab1N))AVCe2
JO<K>S0/0?+[X>KR@/CVRX(.M5/;BgC2?8fS.PXZN:a]WUD&GSV\^?2ec7?IC.f@
Ya.FO)MT0N)cRVZ2Ze0C9&F?&G9LTeZI)g1P2Z\-1I+04SZWaG.>gS^EQ^e<P97a
VJ7Wb6\b.75PV8:J9OATX?K#_X/=/f3@5>&:M5QB.?DO@FQ4d70I,EV(KYHM_K(O
:[/_c:f.J\_Nb7N,#@QCATUT&9>+K\#U/5KeP)D7\Ra=e/-;(g#NNIMZb)gX7,VU
LRLE1Z4-RHB3/0,Sf.fD60GIEZX^\-8H[ZT)/-@OUS)FAe?_E#4]GE)c-S1HUWDF
6A\6.XQEgE#c,5g=4]W)0YV:SPX1fXd71MHX_@R/e#P5@dV8S(PD7#Pcfe6V(gA,
E(.12=_X?[>I^CECf\[a:?.,Z__)R\[O/b[L3RM#gO-GR3X++G&2)]7=>085gWAS
Gd=6[+/V;?]@GXS2L(fSe+da0)WL:dbP3b6:6>R5E7-N_A4c0QEK3FP:S]A,O1T,
>W#T^W(c4F,cJd4a:cIRPDZF.M=5C]X?BM09a,TB/0FO?TXM7U)ePd9+71A@E7NV
SdYff^(SPg&\gM)HfEEA0KXPgAaG5Vd>?HMbX/?6=fE;W/WKe>:MCS-f=G/,eU1P
Z/7^Z_(SGB/2[+b7;].CRI3J8=#Z+8g372-gRP@>SRJ8dOI]Y=T\7M?He[\XM=W,
)(dCTW]9c[^:G=/6(1.G3BQ4(,T2L:U>6.#8;g2-XWOL1GG\=:#UDN5ZER7CgWG/
a_LY9>DG;@(V4@fc?F&&9G=CSG,&3XEgBH&3c:,,.ZeU&Nf/cB)YKC)g\E=fZ:KA
2E6DTB=MF7-gd,/.\@L_E4[C#38MA5+3^SQVUCfXUD0g2I]F=;eRM4?S/W1fQLG)
\X^ZX)ggVEfYBA=e[bP+&\dW9Sd[XU/+87G-@&cgBX\A_eF[dGA3Xa+/+?BBXLBT
D&\9F[7Q7<6ECKO&W:5dg(4Xb@]ZJ.H0Wa67W41WQ@e=H+PfY[WS2(^]1FV=#4^,
D9/]]XA#aD:(/3NL/LF)_]Y-9E>769,UL-1,a7>L@7,Z#VT]#T\4KeA#DVM)K/3S
Q_PQaF0UIN4(]0.Z6C;ZcaX<[EV\+0[T6<\b=8V?=8#Z:W^N4@<D;dF5)D<0_U[M
VcgD81EALZ5HC2gDdWd__5<))S;(O6O(M^[^R;:>\XPM2&eSdd07JRRC2G<?_2;D
a4=RP0?MbG^[FY&,&+;B/HFXHVFOVVMQ(bD3a8[QQ.Md5TC]K.\gZU/3EYC-E.9O
aWWNDVeQG?cTaBY9b5UQ>22c/F_dU8TS/\#<DbCgUVY6fg6COL>7#89ZIG&:PH2.
>J#=0Y>eGB6e6d6d/):N))cafRd6L_dL,A:ea-?_KC&^6eNQ=e)60VRM=b5J1eH4
WYBR61(d)T41AHY=>NV45e5Z0RR;7KMeF3cdd;#:bX/\.L-J<ABF9>Y+T&JM]L=7
5QUa,]300,))@TX5F&ROE+a9.\ZS@3CJP4GXd;DS&B2E3fa:M_EDV6H1+>@d:PC]
\[5<eI1(R-Y)aW@#Q\a[G1C^N7WIIPE)C669#NIB3BgW3M89d#H@#\],_.\JW.U8
<ATI\>e03Q\P/O-X8-FbMW]b&dCb2ONT?[B3Rc,@NPZM;0Qe2KgX8eCTS9JFJE=]
\LC6ae/G4GdW:dbY&<\aa]A;AAQ_(7H)V)V>PAWC/4[4)-dMX:?cSLYQ+:)B#2PE
:OA?<FJe[64gCJJWT7W==,@\=D.SA/Oa(550XK)J+>3JS6]YES=><AWUW(:fI_=.
Be1&O__6Tf<Pe-+bfG93IIXWOg^d5ULJZ3QPHO6C_8GQb_AA)H.M34:B[Y(1IA^D
.VS0V(V:7U54_a5FJBN?MP1NQ(SZ]IZH/=aJV&-(VFMP85L1O(^ENF<0K,g^8[>;
QKe^;O>?g)a\bIW-Q)b,/DL(<L+IgUX41OQ(V_cT9[H+#KE>ZBO:0BKCYdN89\4S
MX3GKbAbTA-61G_McV\Y<=aZeI_-;)6UP(Z6aZR\[JY(@4VO+YGZ&MM\/8cBTg3c
7>()DGJ5Q9M4fT(_+<A-1:.4Z:2_Q_Mg/W/U6/YS_=\H/<bX2X@A2^K?WL&b,QEd
FNUbPJ:1Dd@]7VH5OPFXP-M^M0^@\^>]J#g<+eRPI&?QO:I3g^<]K;b\U0dc.M#4
S3,1Z>VXJ79L<2cWdeMDIFQ(I[BKA#/_4</0;e?JbMVdQG\Ja:bK;Q-K]gT72#A;
&\#.S^UF]\\WR/)040X>;11:PS-WPg&TK^FKa_Zd<YSB;Y0:,0JBAQO4?D//B\@6
9U>^Q39\/R#3DQM5XQ)G<VA4a=O<EV?B3^0NM-P)<_^ZA5(@RgY\L+I^>2^a1+c1
Gg4F#FfEZFYcc_:<,4V1[AA-U,>R723D7WS1QRY=^,DBHg]0a^,\Ce[K6[9ODD2/
IL6^O1>83RXS5,^22;4>eFCIfF2Kc=?NF[ZC2A</SUc+/^,d^;]G@4S4;/PO@f,T
WDC,B:b-0E>E8]Ud8,PgBf0FcA(-FL082S.I=,]a#_8MKUB+=>CSLd@ge73&;849
1R^#?_;.f1Z:FOMZ;V+.#L\I>,UMMc,XG>BY4gCQ-9G_@T66BKe#>TV[KJCW6e&F
IgTY/]?GA6gMJ.5OBcQXeI0;FZK7NL6Te=72EOZ1K1Eg5MHP.Ha+R]&-(MDb/,E#
(?V(\eO-S-geJ6I0:b+O.HVJ7:Qf_72/V,O)AMB4\a6ASLSSD6[WBRKQMU.YQ0^U
LAAZ0G_M3LJ19+=7aHE1abK)3&2T_082@NR,f4PAHAIV13S-7d_]N3.2)6[ONORC
B0_N/#>X6FIS/eU^+AB5M>&B)OT13Z:;]Jc2BL,BaLG0<F@^I+CW9<f^46=3Ib5P
V>O-:S>BKYbAed94+BEI=H9NY27.ea+&@C<957_9W7=_Gf\F\(7a6SA/B:e&K8MZ
+K7X,d<aDG5d(^P,c:;L#2FQ]-OEEKO38E-XLA8T/9KWV&S7T0E6Z5)8WN,BS5+V
.)XT[+0RBJ>N;12A(ge7AHcM)+A?4d[/W_e>Y(KgRcRIHe]DM^MATG6V,NPQ.XME
:[^.L9D;,d<9Nc@OIcG]gE/\0B;+CNZW\DBHWEI,[TNFM;b=Rf>aSWZ=-<a3C;EU
1(.AA&a&OI4gO:ZZ1UdLJ0-IN\ILQV>GIWebD/cH+ON;O;4CB^e-#J[^R-fY?dZI
B;0>5-S5@<<+T_B1PK@D>eEgZ2d5V@M50BIJ-FB5>b-RcgH@]>[P?Qa47S+,;Nc<
aSS7]:aH&93<^a8#gJYKX3/D2JUa[fA/ZE^)A<COCO.ff#)c-B^I--eg.PN(<c9B
CgdE=_&/bSQ:-F&:->d:RODGF<W3Re-<&Kg:JU0(48T)FC,A]12F,I2;<VF5\.YH
cG=+XKYTe^@US63E(2V55TXbCK^)[]C5VGT@)Z[^=:M.0Ze)TV#>NZ.Q=MK,YMFK
g-:[:?P^5RXQ[7LH)eYU/&eQVeQ\A(\[b1NG&_K7P=(+7K2Ug39eNN](@fRFaOH#
U@]8EdY7Q@7]B:XD)_RWa;43,O#g,G,)#CC/E31:b>4+B3Z3([Z10&+V^B487Fb^
-QKQb9LGBZ0)RMS-[SeAY)b]_F9&H[&,X32DVd[Y&8X.a_0>cR+Kc^[JDf//K09f
\;^IEUDXHH\UHX#O]_8<eLH9C4A.T3K)SKJ5VfcW1,++@7?=g@eC+YWIM;C>AV6X
D0>]dg4)EEJfEag2bV>CVN@XGW@Z6S3N+I\TK7U<SL4FSM_;=3[5CYRFCce8OSQ_
05Z:AWA48\.KMeEeXQ1).:-f<PT@/+d4\>7WNH<KcZ;T(WF]&gM/0^gAD=:PXANX
GgPH&_;.8/dKZcN)CW2P[8[P;HM(A^L_W1M2+PVW]@YX06.BeS#XL?9UMUb_R]C1
80,0X:I&IJ?55bgB5RIgEEV62c_<QSH]X[S8ZH#6;Q2PB\Z@JAUI7],@:K3[B@6,
-#VV:3,41D@aM@7BgCK]=Q^Pdd(?L:3W\(#T.JJ4]DG\gF-5ST>V2Q.U@BB?D(IG
/:3Va4WM7G1;V/;/F-A1fWKO4]2d]XKRRXK3/+#YD9VUW_59\XO+U<T/2FGC?RZ<
Y[RSM(a6B-.(bGOQ6,+_^EE;d8P1A+A6S)PQ^T-O&_O?S<+GEcdNG40L<PPDX)A+
U^W@+NOA-AdO]7NM\CJ3X]<I4V<^9/]-49Y[:8-b[?,&-#T0dWO\QRJ,cD:)MVZM
ZHU^HINcMJ8(:GcED9.c[-S>(YLE=US2fY\2dKdB^AbRPGf;2^BTBbULX?L+.(<?
CEJ<(6VB@HGMCfWO.B7ZF_>32]7[,Y<=/S+_(G&-V]7#NYcQ2VTJ1QF#K+E6-\RK
GYE<WM=:,2879a&D_Y)]3Rc(/DHUb-A]MO,a:ReGb;<]B5XEa=<MK0LgeF6QQI-c
9)AMba-Q2]Q#FcY1B+#:HSQ:8O;]9(I&CU5a=40[OI2UJVU/3F&f#X-T]9>88P;N
RW0E;1H^LVD]Q4JO-NI-_:gd<2(K?1+6[_U4d8(@PdNEd5OY6)PP/3XBV1?D?#Sa
)_(03RVcJ0SNCgW56.G9,:J][0f27OSK-?J.;0(C9:N=V<\U80(3MM,P\3P6bcTU
:C/0_E&3<:2&H1Q<9QF:)de=@4^PC@EFT5SO1R)a)455-94[_:K]1I88\6_=JZ:6
/Q<=]?/[KYI3Q#/ELAb[)T(ZaESOa6]Lf.HYP1YBTaJ>88W>_[UIBSF]7F]b<XJA
eEgg67ZA;U;R@(.+U5Qg-9.^&aVB]9?UHabg5bRgA7RPT8;<EQA?=,_V[N5/?DYF
G+EL2=T_?>7d1[2M+5[)\[T.;<)f_\)5V@332BYZ@fcZMVbY7M1=059WSY12?<[\
2dUbL1OLc;^^?GIJ9]1X3QH64>1=\>:B.N=U7-W_IdKN5Hb+4B<_2CAdf5^,O7V-
K<(9gM=5151U<4/QcO1e(9/QO6J@QYBc(),#<a=N7c<)>W5bFTc\RbNP,[>gB2T?
:Z\8KLO)VC+V>d7F]#BUL@<^cH&9#C>#JFc2aG9-Df9@>K7OIPf]>BG:g8M+]E-/
T0ebW/YH1MJ/>ZJ^^-F8@M<]RTR)C\Fc\a#F1U<M9V>:P8,eV3?Q&@&L-g[#O3DA
[7b?_BLQZKU?)N:][e+O3[MN:FKC#L1R>Tg1@]^(:9>UCKe9EYY=P,RK?5bbAX)0
.&F+3GZdAJ_I7&+J@^##Z3H5U^W1H[Sg4:NO+^Kf4N8b]PSQ&9CD[I;a3.F()1f\
2@]+/S,-Nf/:YJ/VD6Kc)E]\-,_@:#@D#P+7L_]\Y8=54[C8PA:d^O<IR;Y@:P=@
2)Z?3><NPeQW5:33Fad\GPN6Q89H<M,M3.=@&)9P^^aK6_C6HCUa?QRS1g?]Sb,3
5g+VS02FKWfM\Y#\R99.0LY/SW1N@JXB-LW],P0:FL>X=]9=AQ^3[.>a2R>L5EGK
XV,Za6?#;_]Z(LK1;2I-A<Cb+beX)UUIe,@.BR009PP)&VN[Q?4_9bg?J1aC];dQ
.;5_L(5b58(RT>AXL7<_E,AW\Lfb83D89;8Q6E8;NB)LM@J1TVI=064>[2Q;8GDc
)3]^09-UPJ71=c.dY,8G)&OU;e3R)LQS/G?RgST3e;W2<\1EE+g<67)(Cd3S1Pb(
<F2N93YNIgZAaX):bAg?7U^V-B#[2<6@QOJ8]c0A0R0&6MG)TW49@PZ9cg(_C1ba
ZNPZEg2A[(2INRf5GBM93,,=@3P;cQK[_<5+,SMQGV^#KU>,4cU)APEC,9N)(2RU
&8efE[Ja&I?PE9d-F6HVBCbaVV6CB(I^_IH>LA,S4W=S^;F;RLQ;,fH\D<U03,g-
=Y,.<ab&IYU(-V,I[V/TC;R&6H_AaK=4R)WE01>Y8_:0#\+)f/UV^QY&-=_.IL0.
L]a_IS\&/9gL@^8/LYQDb9(g]VBCYd[FQd]EcPZ_LBYE_RabET7)dbT9cb5/33/1
MI9QF?7a;-A//P-Scef/K5b]dIQH<#I#43H+dcS6L>,IYLXI4N>PZ01DJ>6JQ<e\
)#2FALW:>c<)H1@7OFdFXEf=+_]A>0]VI.C[V[<??2b@;),T<GEQ?c@bB-H#R3G1
7L#@P<,9=)6E0MOCbSG90F6a4aLdZ)c^-BeSK^;0##&XV7CGDaA_N)_]CDFYZeX;
SMNQ8.-Z=T_-C0N78Bc<R2YJ^1-M&<V(@R5M->0#)S3O:GI?5_P)NVR1UD<L+B(N
U>&OOeFc0PNVTZ2_G@SAcV#&JKg21(0&4E5#4(ff]31BIaIg9HW=[51#;]+eA#LC
<0+OO@HCTZ=AgG\:2[)&L93,T6MJd4QWBILgcfOOaV6.7/bPCTY2/4LUSHN;_/8B
@^(N)5(V5V:89(0=b2S1@a:P;1fD6QU;<P_Z>I27?eXZ6VA7B-?WA(SQ=.fO[-<5
]X;38?L.-g@eCJ^CF^3dTbJ]65Y..4WS#\e/)3?#fEbQ;eeAI,BWNQ37JYa>@=V]
aGWW@HRDa26,]-)D8NE]P&UCW9@.9AVaUc^]@gSC-F3fQ&A,BWc#&?AW[SB2<b?H
A(Sb;6R&VKOXT95+A0.?_,8_BfF3f\#C_Q?83;QRC5Q.\MG.gL4.&,DIA:;DHII-
ZS>c8?BZ8).OgC,]Te/I.^I9aIf,0^[fa@;C<W2cBRI1VFHfTFL7>]V(ATa#N#0G
7O#Qd]U9d,KMP^:,_AUXfCeb?]/^Eb9:JBe6g4/?X\@S.g7R-^<:40QISe[?^G=9
7[R[-E:g=;2OBGfXcG_9];5T6JWOE#Q-Sb,7ag&),<D5#400-&0Kc67XN9Y.db)W
&4dgY]-fKc2NKFBDPW=;fe[AYFA94/:Z]UGF<U(GDDY;7)IcK,ULQg>@T8R@3EGT
/Y/=+OT]Y@?bWPQ8D_VMc<3=:4SUO<g0\LaeZAH#CJ>K^3Y@R2+VB_.c_V4D_^DG
4[[.P1YaFa3H6[9-b6;^U^\B>dT\:0J&7TMK;T8+,Pgb+R/W\]bOdW9Y/Y>.JE6N
<H1^2)J>B?6&a&RbDc4K6AJW#g;F_\(+166-J34).#8A]bJP01R;cFa0-YeRT<<7
=-;GHO664>+MZa/G8L[>M?QP>6C[]CQ;.cag6^.gRAS/&+M?(VW/FVGg8X@WR\Mg
U>9gPgRSN1F3&c0VcA)eCEO6L)fWHdNV9-.4fJ;d3ddN<VKb0VN#.D)GDTKM_Ta[
._8CN@H_)O2O0.^J.9@5NV,BAU9?9T0GP4O_Uc5J52:&ULfB5R7;7Sa7G9YY-GJW
?@?\(g-Z7JT2_5;TG+_DU0J9_5[DQ1d^BXH]e^9MD7AQO;(D;bHYB9W\5f(L=;db
gA7N9@0cVgH^@GYQ,Y-YT1PU#2=3L#gUXG4SBeD@T:@Wd/8>O+@E_,<7\dZB:d1D
FYW8?#8A]7G[O3d_9R:8Mc+JMH3&30C9GOB84RR]8B\_FPDfIMd:K5DX_)f5@5IY
S28RT&WC[3NfMM8L\81cC19:W.2c-]DbPCDTE/2L89;+O<CgJ4-]:I@DXa]0P;dR
U2FI]+U1E-P)b4K9(_^Z9W,&3,?<B/>fAF>RR7EBD-X/d4@WE#[\PHBa,=&U2ccJ
6;M:L(?-QNZ:S0U0CV/SW((.6c;fI_9;I^/3UJB-f&?.G:DR)M@QWE2c3D&,&&+g
3ZVP\Q3B8fLR@VJ&G/8P&6?3UU&b?7?4(gc2EQQ__U[^gB?:=<eS1N5^AO>\T+fB
-\99)MVBHed<cF.4fE56Z\@1H37@C_9S<[a_/D0LSP,#c84JNX:Bc25E5WDKK.[2
+bP>6WM=6F9P\<?8I#&0LK]F-R87b);Y61?3Y;5-EEB#>-,a4D/0.E(?GDacN:XK
Wba/U[87-2HS]0/,0W2S0NK[]WSDMNI;VBZJ#&7@=aAO-9SF6F9_dEPS7E+UG3&I
-)S3H5Q;b;5>>IK_T82CR8_H0](AYD?,LE/\,7^HD#BU_BU+LR2&aCLX3K@0>/[F
M/5=g.^<f&#]]-E]I,I<A83]_1d.C,CY:YXD2II0@gS;_GaXVgbfeVF4QeE_L]<N
-U^>PUJ0_E>]#5bS8+6M/2I]YIPS4[bBF:I9c?EE-<[=W5SR^(</cSGO/MP0OB58
)I5+P)3fVNddKeN)W4[(2;cPW)SIDe,S9(;_A[ecQ#Mc8Nc0bI=WUU28R/656Q,9
4,;_f5^Dd,UDa&P^#MRT6faEL46:VbT=G+67UV?Xg2\@eFb)IG(I6_-[)c6#RfS\
G-I_dc5\N\VW&O;IMgF@#g@bVJJg4_ZbDC9^9IS<H4dEG\AABbLQV-T>HW0cc6F&
,9QI-e<b7f1ICJ)M(UUAe=PV[6PH:O<I48]6WXQ2\0]\M6Eg2BYd0=<>aOd&.6B5
):LNOV8OO?dU/)DbW9\CU7:g\5B02P_IE=5)<_A[5P7<0^eU<RYD:J;FW/?KJ>bC
g8D]9CAN@TRE3_)0gD3a:B59S3<UK^&Oe7HI0Hd(LXXfB?6W;<d+\,#\[\8.g2.&
QR/DUEFU3?OJ-3Ea/.=,a5P)63#-6LG.5@Ud8<H;O1=ZTKdI87OIUbZS4fA&/_E(
g,R]=ITMHO_7#0L<575F5A^^Yaf-f9EL:KPF60,]JQGdE3]BR=A+,3E5eM#KN()A
be?RZ?ZQ\6X>C4)_WQ(<1KZ9KLWGL9Q^Y3D:48MKTdeSP],UaBQW2@df^bK#9\S8
C-MD(.e&?X)#O=F24F27J5R5Tb2SXRB8]<WE.G8JW+Z(-@7APcH4W-Va@IXVWSfZ
QKQT\\I-@;fe)8E\#2D\.3UZL)5,THN?ZT.45@,T&5G6Z9ggY+2bR(<9A2MePED?
P,,C3NM9H?Z445U6gPE9;\7#Y7WI>ABRUNQW_H0GURUC5gVL8(&P,6=GaA&@)bN)
@gbQYg0IPEJ>U2^6^,O>Ic#S&7,0#W46]MTVeW.fKTaJC#F#U2^J?J;ca+;F?[<e
^2B422NY[A+:B^]R&J+>EXU,^Y\#C9cK6]12T7F8_>Ne4C>><;JW8[@(@e_(3f#?
0^&>(C)<33DRVO^b\L.2S3T]<FS1>4g(GGW+O6>QEZYWP^BSe[RHFd55XJZQ75LB
Y3>0@248IE)9a(d&SYPTE8a64=&]1;HbOQKIeRS@JA_G?.05+47<P@dGC]Q/b;U>
^XgSUM)J+-[H&[FI/JS3)?TC059W?013I])FIf0,H5:P2?WZa^<(TdaJX&a1daRg
U-;TY&9Y5)^RHbZXP[RGGJ?7X^\4S0O0NaR9GKTPYbAQ@7R4^CX.MXSbNg81>XUe
fZ(F,a@UWY/:WT>T^J-8ZVCP,9K9UA,.aAOW4TDeN+@@4=K\\Y@dE&^0YT0BF;:F
8_D&<#1&>f>E-cdK=8d\dL/P6QbGT,G_44aW9bO4\-fe)VG\X[/9DJBK+K>3N>@.
2O3IVGRZ3W9LI#:QGXA2Rf>]F1C=<I7C,H@C@E\b0-?N;L07JINaI#:\UCV+Q3aF
GA;FTERH]QWK<d[4Yd#X2RQW]@?NWe-RWB,67ENV:S@O3_X;IFcR\2)b)gX,9KXE
,/H6_3?Q_>f^\<#BX]0GCdd3)ZM@SRdGNS5f(JPe)Y_#Hf,eL;2Z;0Q>-_LO4]=5
ITK<Fdb:b=^,Z\c8N(:5\[7D<,Vbc/ZP-39Q_TNCRYR_RQcIU5[E31@34>,/e.H.
12XZ[>fgBPJY/RC7g>P7_9.J@c1I]FGGA@?e^NO]Q-<(=AH34BYGe4E2KOaSaZ&>
UC\S#0SA4JcDOZ.WEDDEH8Z\C0E:KDB-#,#<B;a[K2YZN#/5dM)aLD2KQK.4IQ+U
eG6#V,d3<HPXfC?O(BcYXNd]5RCf(Bg-b_//7VbeSRETDXBEUU8BJ4gE^)83-,5G
:8WNMf>PLD((:,]#<YEa,1=0?5\(NAQ-e9RRERDSXM0=aSFOV-9[P<6[V<Y3B[VT
,LF@DZY5<A0ZX5C9^B7C?I^B^)a34OMV_cg0a=)E/a2+H\W2e<.bLd?5.R8;KJ(6
e<8Z:DdX/Ib8bR97\?9PP6;7T-/R?W-0+(\W-Df^83X@0\c]2g2#c1FSQTWEZB^]
:80T7OS)\-#Wa+dC8I#1^[BXLAT\KMZ=)3_@P-JY.LLI_9M;e&Q@^OB./eMQT9O:
O(M=g(]UeIP+2VJ0Zb&a8G-KCT[04f[U0J\>Cb31&3SgI\2OKR./Y;#[<dgM54;4
8[2H^0BeZSK5aAQH:K.(PAb5YQ)(M#JD+X+9AL5UJGd.:bg3G\#aJ@cN]>eZ\H,V
>]=;<OfXLELa>@C[=\3cdMPN,U-+g8LWe+X+_f=c<V7=;F#:3,bg\64Q\Y1.S@Qd
,;@4H^OH1K-f\,T-)#)V1)YaR.fZ.89\,Eb:6HZE+9.QSOIeIR83IM[,=U?)6L0Q
TdSGG(&^)[ZL9,]3D_<MbDHL^a9X:H8CcMSf:PL+d@LKOCO:,NLR818,]KH3<L-D
EdA_8-[1<N<8&1-SOT&Q>(U(\I+fYR/,c>fL9W.HF&BRZF-C/;<R(=G8XfQ93Sgg
d)TR2N&Xe/[.5L]<HX6W<W)8=HGN;[+EZ:Z:=E@06@-IYX9X?J?H/1f)AF.cb_>W
7L;4FOXefE[7c:+IWZf3GYUYB?KKCB&?[QHQ?,K/I)/U9EY95daAaGe;#&Sc3e0C
YgA-;G>H,?;0FT(3cM,.g#XV8B7AVagETU).S>B][24ZJIP=(fA7R.Pa=D50Z:OI
c7OP,gC,,:De]b?dTa5Jg)K&,<2JS0MP8T<Kf,,?d=2>--SQa_6dc@HIPZ0LSa.(
-NZ:/f]Q/cQ<2@_F7+SN>bWfW<F_@8^b6]Ob++VY<Y:OJ^f0JdUf_XPbR3L/gSH3
+FeED2N-P5K=FB<QRML<^;W.5FE;4G1\3B#CO(HKP(JFM@?2fU9gLBZWFRRV(^+^
I8\MBaS9^2&ZNGa4AWB#25U4gZ/2;;Dg<XGMF2.>3/&3AN-)KZYRR#+XJ=@5;Y>g
<U,C5MgF<1276[1b<VO-a@Z_A=@8HD5dJL_:^+(^eXE?PUFAXY^c_-,W;#X3S#9+
<4\S/#S<CO4H]FB+aJ[<>3;5WPcd;2EdCXM3ZUe_+^EFfH[>]6B:=-W9_.@=Y-3V
5PC8e_N.@AKN8KR_Yf4U23bH3(BDDT:B>=VS^f/D7P;K2R]:(UZR4&XLXVHeSGdP
c:0F^2f:7Z,U5)I,:bHe\c]U&CZ&)[B6O@T?XQKSG;RUfc]F4743bAK_V7dXD[?:
.+=I9OMEYcA66\V)E7E76G&XFQ5X>g<fc)VPG^H5dL&3KSf;;./&AOTA@.a9XG&M
:I--O,OLR9@4QJ6a:MN=ELEV+M]feD<:OXFT4S-^f/+?RDE.f[X\[9=-1JW)-Ofa
D2fP@2URda5JLcJe+7S_>8T17F,[Y=b68gEGfH&\+66/RZbPY6A,05G-,B8f\QaI
7[]/S:bI@ZgI]OE0WL_LPb+_GUKd;FZg32=3gGZI>Q;cAS@/[+12eFANcP:J1[>)
LF9J-=R),U5SR7&=X@1^Q:8Z.(+2c3(e=VJ^,gR\^C3R5[Z\Nb:)T.2bD1R^aJX0
&2VCbSW;_O)eZ\e1R4G5gY+0K,fbB,[F;K:LETPRL-O2J(84@>U;LFcdE?(3-@RL
XBM<ZJ3XAMTRc+6bZTZ;aWaa0^DbP\7>dPK6T-L8OCL=-N-K.a3?=HJ[cD=;3G=,
FLF)fJE,0e],)/O1:Y[_A04QKUCP-a5>Wg#K^3ZXa73NV&b(3)P&57\_WadBK[dc
O/.O:Kc&ZVAFHBe,OcR\-5I8JX(N=c&-7S<e76GB]]2DdD^T8#e(4I\#I5G@(@/a
We.;UQM7LPDfE:-cC23RWeW\EIbf.KGSHX6O:_/eeHJ>2N8fGZgeTbaUfKJag#ZE
5a.\@.[ZfK]_fCHR[6_OPNR/9\WLS&-dGATYPCe0..Z:N=(/G3GCf2Zc-<d7A8dI
?]8>d(EeWNVVaI0b3,=J5>3M5RNWg0&;]VG2gcK[FIe9Y>;:b^c:a:^g+O\#]<7e
SeAH^8+CIg3PP,EbUQ=:7W\;EY)6:RI3,1W8Z25K]WIJI+PUZ]f#B(P0&HWe-CY6
(\2I(+R1ED:aF_2XJ/NYU_,Q(>\<(DE@=OZ1@,AHaL<?]ccHC=\EQe:]<5e?/R[c
g..14Jf3-ab?6KR)]R.\C^b=NA&L,aL)M>D<OO&>a6)8S<VcIQ(.[^QcICL8-9cP
U4EXF7f/SEAXI4IR@Tbge+3>88D()<-(.[(NX#JR6,57B57.\O?)GXaL)6K<D/10
,^dN:c\b:&Q?H3DP;A(B5a?aX@6[<_c2_,<FA]LA<IKRPI97&LEf0Q>H:R4HT-Q6
6T5[JA4HLJWVIVI[I^O&<LEd,R-OOIG-[V&0K?\R\SbV:>ASXJ-A5263(V&J9H.A
2IAfb,X?Y2H/1/#]]U)NMWg])@6UVY]RQY+LE;.;8Q<VC$
`endprotected


`endif // GUARD_SVT_AXI_MASTER_SV



