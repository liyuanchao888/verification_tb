top dut(
.clk (clk),
.rst_n (rst_n),
.paddr (paddr),
.pprot (pprot),
.psel (psel),
.penable (penable),
.pwrite (pwrite),
.pwdata (pwdata),
.pstrb (pstrb),
.pready (pready),
.prdata (prdata),
.pslverr (pslverr),
.reg_sys_rst_ext (reg_sys_rst_ext),
.reg_lines_num_ext (reg_lines_num_ext),
.reg_rows_num_ext (reg_rows_num_ext),
.reg_channels_num_ext (reg_channels_num_ext),
.reg_filters_num_ext (reg_filters_num_ext),
.reg_layers_num_ext (reg_layers_num_ext),
.reg_kh_ext (reg_kh_ext),
.reg_kw_ext (reg_kw_ext),
.reg_stride_h_ext (reg_stride_h_ext),
.reg_stride_w_ext (reg_stride_w_ext),
.reg_dilate_rate_ext (reg_dilate_rate_ext),
.reg_bias_en_ext (reg_bias_en_ext),
.reg_relu_a_en_ext (reg_relu_a_en_ext),
.reg_lrelu_a_en_ext (reg_lrelu_a_en_ext),
.reg_relu_b_en_ext (reg_relu_b_en_ext),
.reg_lrelu_b_en_ext (reg_lrelu_b_en_ext),
.reg_pool_a_en_ext (reg_pool_a_en_ext),
.reg_avg_pool_a_en_ext (reg_avg_pool_a_en_ext),
.reg_pool_b_en_ext (reg_pool_b_en_ext),
.reg_avg_pool_b_en_ext (reg_avg_pool_b_en_ext),
.reg_gap_en_ext (reg_gap_en_ext),
.reg_sc_en_ext (reg_sc_en_ext),
.reg_sc_add_en_ext (reg_sc_add_en_ext),
.reg_scut_mult (reg_scut_mult),
.reg_scut_add (reg_scut_add),
.reg_scut_sub0 (reg_scut_sub0),
.reg_scut_sub1 (reg_scut_sub1),
.reg_in_bypass_en_ext (reg_in_bypass_en_ext),
.reg_upsam_en_ext (reg_upsam_en_ext),
.reg_upsam_input_size_ext (reg_upsam_input_size_ext),
.reg_upsam_table_rw_ext (reg_upsam_table_rw_ext),
.reg_upsam_table_rr_ext (reg_upsam_table_rr_ext),
.reg_op_ext (reg_op_ext),
.reg_op_next_ext (reg_op_next_ext),
.db_size_input_ext (db_size_input_ext),
.reg_relu_a_ratio (reg_relu_a_ratio),
.reg_relu_a_A (reg_relu_a_A),
.reg_relu_a_B (reg_relu_a_B),
.reg_relu_a_C (reg_relu_a_C),
.reg_relu_a_D (reg_relu_a_D),
.reg_relu_b_ratio (reg_relu_b_ratio),
.reg_relu_b_A (reg_relu_b_A),
.reg_relu_b_B (reg_relu_b_B),
.reg_relu_b_C (reg_relu_b_C),
.reg_relu_b_D (reg_relu_b_D),
.relu_a_zp (relu_a_zp),
.relu_b_zp (relu_b_zp),
.reg_gap_ratio (reg_gap_ratio),
.pool_a_kernel (pool_a_kernel),
.pool_a_stride (pool_a_stride),
.pool_a_ratio (pool_a_ratio),
.pool_a_div_nomal (pool_a_div_nomal),
.pool_a_div_pixel (pool_a_div_pixel),
.pool_a_div_line (pool_a_div_line),
.pool_a_div_last (pool_a_div_last),
.pool_a_pad_up (pool_a_pad_up),
.pool_a_pad_down (pool_a_pad_down),
.pool_a_pad_left (pool_a_pad_left),
.pool_a_pad_right (pool_a_pad_right),
.pool_a_start_ext (pool_a_start_ext),
.pool_a_data_type_ext (pool_a_data_type_ext),
.pool_a_cut_down_ext (pool_a_cut_down_ext),
.pool_a_cut_right_ext (pool_a_cut_right_ext),
.pool_a_result_line_ext (pool_a_result_line_ext),
.pool_a_result_row_ext (pool_a_result_row_ext),
.pool_b_start_ext (pool_b_start_ext),
.pool_b_data_type_ext (pool_b_data_type_ext),
.pool_b_cut_down_ext (pool_b_cut_down_ext),
.pool_b_cut_right_ext (pool_b_cut_right_ext),
.pool_b_result_line_ext (pool_b_result_line_ext),
.pool_b_result_row_ext (pool_b_result_row_ext),
.pool_b_kernel (pool_b_kernel),
.pool_b_stride (pool_b_stride),
.pool_b_ratio (pool_b_ratio),
.pool_b_div_nomal (pool_b_div_nomal),
.pool_b_div_pixel (pool_b_div_pixel),
.pool_b_div_line (pool_b_div_line),
.pool_b_div_last (pool_b_div_last),
.pool_b_pad_up (pool_b_pad_up),
.pool_b_pad_down (pool_b_pad_down),
.pool_b_pad_left (pool_b_pad_left),
.pool_b_pad_right (pool_b_pad_right),
.reg_width_wrb_ext (reg_width_wrb_ext),
.reg_height_wrb_ext (reg_height_wrb_ext),
.db_group_ext (db_group_ext),
.db_pad_wra_left (db_pad_wra_left),
.db_pad_wra_right (db_pad_wra_right),
.db_pad_wra_up (db_pad_wra_up),
.db_pad_wra_down (db_pad_wra_down),
.db_rd_ram_sel (db_rd_ram_sel),
.db_wr_start_wra_ext (db_wr_start_wra_ext),
.db_addr_initial_wra_ext (db_addr_initial_wra_ext),
.db_wr_finish_wra_ext (db_wr_finish_wra_ext),
.db_i_cnt (db_i_cnt),
.db_o_cnt (db_o_cnt),
.db_sys_st (db_sys_st),
.db_width_wra_cnt (db_width_wra_cnt),
.db_height_wra_cnt (db_height_wra_cnt),
.db_channels_wra_cnt (db_channels_wra_cnt),
.db_filters_wra_cnt (db_filters_wra_cnt),
.coef_i_cnt (coef_i_cnt),
.coef_o_cnt (coef_o_cnt),
.coef_sys_st (coef_sys_st),
.cb_mux_en (cb_mux_en),
.cb_rd_mode (cb_rd_mode),
.cb_update_coef (cb_update_coef),
.cb_in_line_cnt (cb_in_line_cnt),
.cb_in_row_cnt (cb_in_row_cnt),
.cb_in_channel_cnt (cb_in_channel_cnt),
.cb_in_filter_cnt (cb_in_filter_cnt),
.cb_in_kw_cnt (cb_in_kw_cnt),
.cb_in_kh_cnt (cb_in_kh_cnt),
.cb_out_line_cnt (cb_out_line_cnt),
.cb_out_row_cnt (cb_out_row_cnt),
.cb_out_channel_cnt (cb_out_channel_cnt),
.cb_out_filter_cnt (cb_out_filter_cnt),
.cb_out_kh_cnt (cb_out_kh_cnt),
.cb_out_kw_cnt (cb_out_kw_cnt),
.kn_i_cnt (kn_i_cnt),
.kn_o_cnt (kn_o_cnt),
.kn_sys_st (kn_sys_st),
.quan_a_i_cnt (quan_a_i_cnt),
.quan_a_o_cnt (quan_a_o_cnt),
.quan_a_sys_st (quan_a_sys_st),
.quan_a_m_val (quan_a_m_val),
.quan_b_m_val (quan_b_m_val),
.kn_zp_out (kn_zp_out),
.quan_a_zp_out (quan_a_zp_out),
.quan_b_zp_out (quan_b_zp_out),
.relu_a_i_cnt (relu_a_i_cnt),
.relu_a_o_cnt (relu_a_o_cnt),
.relu_a_sys_st (relu_a_sys_st),
.relu_b_i_cnt (relu_b_i_cnt),
.relu_b_o_cnt (relu_b_o_cnt),
.relu_b_sys_st (relu_b_sys_st),
.upsam_i_cnt (upsam_i_cnt),
.upsam_o_cnt (upsam_o_cnt),
.upsam_sys_st (upsam_sys_st),
.pool_a_i_cnt (pool_a_i_cnt),
.pool_a_o_cnt (pool_a_o_cnt),
.pool_a_sys_st (pool_a_sys_st),
.gap_i_cnt (gap_i_cnt),
.gap_o_cnt (gap_o_cnt),
.gap_sys_st (gap_sys_st),
.sc_i_cnt (sc_i_cnt),
.sc_i_curr_cnt (sc_i_curr_cnt),
.sc_o_curr_cnt (sc_o_curr_cnt),
.sc_sys_st (sc_sys_st),
.quan_b_i_cnt (quan_b_i_cnt),
.quan_b_o_cnt (quan_b_o_cnt),
.quan_b_sys_st (quan_b_sys_st),
.pool_b_i_cnt (pool_b_i_cnt),
.pool_b_o_cnt (pool_b_o_cnt),
.pool_b_sys_st (pool_b_sys_st),
.reg_channel_wrb_ext (reg_channel_wrb_ext),
.reg_filter_wrb_ext (reg_filter_wrb_ext),
.reg_db_width_out_ext (reg_db_width_out_ext),
.reg_db_height_out_ext (reg_db_height_out_ext),
.reg_db_channel_num_ext (reg_db_channel_num_ext),
.reg_db_filter_num_ext (reg_db_filter_num_ext),
.reg_group_channel_ext (reg_group_channel_ext),
.db_pad_wrb_left (db_pad_wrb_left),
.db_pad_wrb_right (db_pad_wrb_right),
.db_pad_wrb_up (db_pad_wrb_up),
.db_pad_wrb_down (db_pad_wrb_down),
.db_wr_ram_sel (db_wr_ram_sel),
.db_wr_start_wrb_ext (db_wr_start_wrb_ext),
.db_addr_initial_wrb_ext (db_addr_initial_wrb_ext),
.db_wr_finish_wrb_ext (db_wr_finish_wrb_ext),
.reg_data_zp_ext (reg_data_zp_ext),
.reg_para_vld (reg_para_vld),
.sif_0_debug (sif_0_debug),
.sif_1_debug (sif_1_debug),
.csr_r_baddr (csr_r_baddr),
.csr_r_len (csr_r_len),
.csr_r_loop (csr_r_loop),
.csr_r_stride (csr_r_stride),
.csr_r_chnl (csr_r_chnl),
.csr_r_run (csr_r_run),
.csr_r_irq_clr (csr_r_irq_clr),
.csr_r_ready (csr_r_ready),
.csr_r_done (csr_r_done),
.csr_r_error (csr_r_error),
.csr_req_strb (csr_req_strb),
.csr_r_auto_ptr (csr_r_auto_ptr),
.csr_r_auto_req (csr_r_auto_req),
.csr_r_auto_ack (csr_r_auto_ack),
.csr_w_baddr (csr_w_baddr),
.csr_w_len (csr_w_len),
.csr_w_loop (csr_w_loop),
.csr_w_stride (csr_w_stride),
.csr_w_chnl (csr_w_chnl),
.csr_w_run (csr_w_run),
.csr_w_irq_clr (csr_w_irq_clr),
.csr_w_ready (csr_w_ready),
.csr_w_done (csr_w_done),
.csr_w_error (csr_w_error),
.csr_w_auto_ptr (csr_w_auto_ptr),
.csr_w_auto_req (csr_w_auto_req),
.csr_w_auto_ack (csr_w_auto_ack)
);
