
`ifndef GUARD_SVT_AHB_MASTER_TRANSACTION_SV
`define GUARD_SVT_AHB_MASTER_TRANSACTION_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_data_util.svi"
`endif

/**
 *  The master transaction class extends from the AHB transaction base class
 *  svt_ahb_transaction. The master transaction class contains the constraints
 *  for master specific members in the base transaction class.  At the end of
 *  each transaction, the master VIP component provides object of type
 *  svt_ahb_master_transaction from its analysis port and callbacks in active as
 *  well as in passive mode.
 */
class svt_ahb_master_transaction extends svt_ahb_transaction ;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

  /**
   * Reference to master configuration
   */
  svt_ahb_master_configuration cfg;

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------
  /** 
   * Number of Idle cycles to be issued for a IDLE transaction
   */
  rand int num_idle_cycles = 1;
  
  /** @cond PRIVATE */
  /**
   * This variable is applicable to a fixed-length burst. 
   * When the value is 1'b1, every transfer in the fixed-length burst 
   * will assert the request pin. When this value is 0, the request 
   * pin is only asserted for the first beat of the fixed-length burst. For INCR burst, 
   * the request pin is asserted for every transfer regardless of this value.
   */
  rand bit assert_req_on_each_beat = 1'b0;
  /** @endcond */

  //----------------------------------------------------------------------------
  /** Non-randomizable variables */
  // ---------------------------------------------------------------------------
 /**
  * Local String variable to store the transaction object type for Protocol Analyzer
  */ 
  local string object_typ;

 /**
  * Local integer variable to store the current beat number which is 
  * used to created unique id required for Protocol Analyzer
  */ 

  local int beat_count_num = -1 ;

 /**
  * Local String variable store transaction uid which is associated to beat transactions,
  * required forfor Protocol Analyzer
  */ 
  local string parent_uid = "";

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
H3JDzlSDT/uZ5IRbPKcMmifCjYRPX4+U5jdQLT/0ZjNKpmf/QnCRRb5k/1sWTx7t
CJBCxEUqYPjplxnDyEAMj/vKRmvYLE+JgcLJYznAiui6OrQ0ZdlBEMchT+PTuOOl
5tXSxX0YTJfbYM07ramkvIMSwobzRMR6ZlaTvccD22U=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 8648      )
K2p+L/tqPCOpsJJFwmmbbyADvR04JwEMc9z9/djVYrWqAlZ/UlXG/TgzmqfM9hbR
FY8ecNiTgLRs74kK7ZvwJmFb6Bnceiz/9aIxZykqUj96/qdbp3dm96rSV+Ha+We/
sXZ1wyuHCnT+0kO0BCdj2fgR3GBBFnK7+w+zsavgopxPHV5bOGt0WbaRgFSEmW77
MDQbpbKoCxaduEFtfPVlihrvWU15UPNbgdjYiq6XAPnd0ZMoVOk+W0lKQr/U+7Uu
WajROPOsbYZ1SElbaC+roGAmLli7Xl+TJbfZqtBMouHM7Lj89jT+CrWD/JaQjw/b
aH4AoG8RLNXKjkZbMQIRYHjn1ipzNolsfaBsqs2UCa7SfNgFkuoiXLlFTRUBgqkM
bKCgQBLMx9KOoyHnREdpulWS4mUWSQ2A7/xfWz/NrePdI2ekAG4CoD21tAB32lyX
ELBHGa4NN6at+qSwnhk5e1+ysU48j+7iy2l9FjReRHThSN+9nscp1TaGvswcf/u6
ppqEBrC2VsjLxFPex18KPnAd8Q+F0dVMieVlVY/0sJ50pq/5nphVWdwF7PrkmZZj
c5lb05Jla3JvWJEgCTeRqzWmFmrXg39vKy0eOrutXzJFz48RR5lFdSCT14mAriW6
OdwjTjDro17aj6gdLiN/lmcmkJjTZBIqShXazMsKJX6MtA9eW1/DVOP9OEvm6X0+
MyL0lBC0QKeOyrhMLjN13sGOKc7MZIuW6X0MrAHgkd9ZXuNr/q/ZVUKc8MxckDGV
4nllpDnkMXIDvGs84qu/dOOxesXWE604tdGPoiSZCPuhQlSFQN3TC1iYKkTfyJxu
S3za7HQ3/LVwgs31WMNfWHVJ20s2fqfnPFVL8DSbSCwtdsEO39LBSPsSjCvgjB6C
PxrDPMyoQ2Ui3F5m8G70Ts0Gi03haunjRE/i7/xIzmlzfqtOJJW3VWEsm9l8dw0h
fJltPNDeeCc1SNFVRQwkXOP6kJb7KJKq1khLfK1y2nuB6qypWUI6Cy172zpHqTTQ
7emcGtmYG31ax+cOM1tMAoO7Kq8UYhkO7SUS2yXAjOQfAvpwhYEdEIb1LjmotJHe
NGIbm23E0J+EiYQWIBCO5fnVZj32ziS6ln2I0yfKZ05hgQOQrBkePoJ845Q+cs2b
3b1Qbf4s8U9LbJUzw/ntBTNG3lLy3M6FrkkJHzWUUf3hh2kZj4BULd5ZQ1hP3DWA
BQJTMDPP/Xvz1/Gx/OY3Irn4vqKygXLsq/xMCSUGqlLZ/CxIT3KO2kpADgmVR6eO
LYMx4iAwMeBnjMvtAxlTRiEvLhp5xc72Rx7xjyo/cNyJ2bUzZxTVUlm4sLanC3BF
6vc7BWDhgKP9iZl8Zo9IeGOGvwNkcfPAHG0qeb3WU7sp3zVEkPmbrUBVhVk5ozUq
o2P9m00SA2ItUvXwlihZN7rrAnOHFLJ2aIVGqEoiVcIWc/wmTpk/xW6VZhVQ8H1Z
lsYE34upfVsUbqRi/1/dO7hrCt/vwHZQqaJpUQIlAG3JzSHxmU2Ov2GCW1QGs6+i
+0RtcGL02A0clBSPxaphEI549j6OR1URlhBTah5ac/m3sOQV0kEIAmY705UfR4vf
hOKeL1jqNjdugFSC1jurmrNZ6doKhalnsM5faCiTPZ5MMpCPSlHBZQRr6v7CTwbt
kOdTw9G/OqRfiLxh6gFVNYRAyMq74WglA7f8QlR3Ppkoy3Y4hVcjDWbXx7df7GiG
G+fucUzClMKMuDGA72jw2Ew7JNFnPMwEB74QHXOKTKuf2T8OuFVUxW5oXxtE+TYM
vQVNjS0NmNItuXE0J0UX8uF+TsWzylwC21hhtCWj2/BW8JJnJP9xOw+oCaoVxA6Y
MeOHlIKanv6wrM8ifKsYRv9FQZUGpDKK5LmnZ6TxYFw4WAzybd1PzH4Hl39VOPGz
UefV9oofgdnzrN38ZyeIC0p0rYObHRghPLrtpGHwJjW1L6M9Gy4Kp+3kibagrH04
P4ig8TKJLYcALqkYAikzXPllCpTA8iX3xD/BeFdoVNN9QnnwiWtEvkiWdKc8WJ2M
N9xRY/YmsM1BspHCPF7lH5ZTEqWCVjAD7dOPjNzKcEULyRnWY2JQydJolgL9gfLB
a8VARUIr2XeHWUDmkP/RWhbnJly4JgqTRXp09+BmxoAbhgo1NMf38OuPZyojT2DG
0BbqRK/DaN3MObWA16otwJJuQvQTfwXdENJU/YFe8DHwmzcO8z8AnPJfqofV/zW3
xWjHtw1oeoWvCI+21C3GAOUukzaN94cnNGpyypaffx8/rfKHX12ZmPrifIpqbo+G
OjszhOBC93SR1kCQchNR1WhQdx1t8ZQX3OLKYyagDfHCV599271j8M8SN66uAWRY
oU2UFtn6R3qY0yK8h4qr9oAD61F8PUe5pxFHhsMjvSxxruCMOkLPjDxIB8P2OTlc
MfCg/NPra/DdM3JCYmx6uf7klww+zBYdg1i4D3FlbrYO7R5Ccu+pCn61aO4QLHNh
ZuK4Eb3ff7t8CRLQXLFG1elbnYl6rgvzg0VvbDmb7tkc1L/GHX74wXJ7vWobGOpu
+aFWP1ymPyj5i90bCC+w38SujD5yzY9oUToU+43Hd3qCEa8/PU2SJL/5bRs1iv9U
UnPo03rxrE6wgT6DEt576AvFfkJ0a7LW3dvxEa4xTAM6kVyJeu/+llaIUuaUbJzZ
h7lJxE8xa6sbQwU1d97y05eJSjECfO3wu8iPO3U3rObjDm29B4w2T5jI67vAaOAx
qN18AEssr0YL5u+UGruPwM2ZewxN6ADU8+R10BNOCW1zRSHvpDTTzeQTKbberZec
/PsG4ZaNqW8wmUxeL2fwe0f3KJYbZv+gt9O0IGiQANSEP9ZsInYBsMtvQYDEsPwE
Pul5isU7l9IOuXTwcvvfDOKo4tLwV8tdQXpy6AVHHEWp1zAnRJDVLOCC+Spqm/JE
RF1LEPEClVxIRj8fXB9oUXvvuIB2ZfbdHvuiFu9VknpzRcZC+IydFvEqmsoN00mv
7yWMXGOtay8TPBClWGyiwNPe/FtlCNrSqBnxiD/xicJhdbo7QBVJWpmaPCYXFi61
BY6XDuOtISnf8Unw6AIJYY9R2mnVe3B/bbvfi96UDB3abD4l+aPjxsZKbT7pbCq0
H7u1CmYTB8AnMbAwrG1wLVeJMsE1fSVR2Bz7z83lzsV/eEVBR+U+fEXTWcpo/tvr
G71XKL45VglBHLyo+vLQtDLKyVeFlpHlWVSqPeHc1uBnkfh9afgey/V8XNEMlHFE
tcgJj2GR5aeMl2E99gT9WoJcvE336kxJ91xqPdBlEbpQBt+/7lbTaC6kLh/ay4RJ
paxBWG0kRhxKNlZF9Qw5kO5IEK9X0FnnTOtnPR5Zi0yqdsvx/wXbE2MFZKjsqJV7
Tqtn62oYYq5BbnXFbLZrnDaiYRq54r6SWZWXnqzvMiT7yXGT6pe40sL4fAd3ey5y
vMiffuyHiaM3CWCGmEtB03x9fvGUvzuc3yYUyhQu9m9zX63E6Jas23fpmCR+twUo
FJ2ikDM8aVANn5m1tXzr/C3gmeONF+U7aimojMlwFT32HBAyRBV7w1eIIdhjFBw8
HE5rWnqzTzw5twenu+QZOBGc24g3LmMaNUJhdEUTLRzyZcfWuSHsUzJ1QDUK/xQj
jGxUeos89X0W3r6dW1jiK87+JgOUCpG/6HspR/4W5nQ8t1R69OFtqay4TsehODqN
2yC7i5jlQSpLGM5v2PSgwKs4/qQ4RDD6an9Dvt/9PD0rm1F3YpkQR/0avAEFRZwK
vrTujUS7SlBYGKhQ9T7F4Q0Yjunlz0zfHFHa7D9bldU509BykrZBRgstRAXGViuN
o0iFgF9jX0L7UpFcHdI2gASHpkgcD6plhnJlsb5If9WKZm+sX9o8W9X0PmKTgBh5
B1trLmUyU0rBGqoBrJ63rFMx8T8f5ALBxoFV6dXDB8Fz4eye8S8mnKgyNzy2zy9Z
ZLYAykUIGfngRRecQjQinxV1y0HNYt6x2jih3IBy3c5smUzHj1TtfxomFMNDFl8I
/Gjsv9ibcvQdB6uhdAuEG8Uiqcu9gdwl9tNUxdAySSiehowrF9cWPmUamWNWKNvI
Rn/Uxr+4j8UIIlDXgexYCbyhAHroERO9D8WfWpzImXWHoDo2lxvhdjNZuB/alsw0
Wif+F5pwLSgMHWRyl73DNhvFeswN2PiRzzFUnREn0OpD/Sxqkfycq5Gv3TR9R+Bj
lIl5O6wgZ0W49tKIhDpu0HfMXp27qpaJ+88EoGlcXNtkObCohK2a5j79F1J8eOxC
nOztIK1LPSVEBXQ8TkQX2BJqRk1NXSsgpijk8p8+7fpQuhjWortNAm8IVZZUR/41
l8bVBHE8SG1zxJuVLPh3xzRgH1q5Ix9DFsf28NgK6s0jf2CqOziVXeZJwIzZrwzt
2CsqR//a/GafYKO2s4st8G131dMv+WePnmMseyo2iTcpZd3ZlJWNqM32jZJPnjd6
rLdENzEBryEmWS5pRZyPWUAP+LsXyQMJOEZvjGDPzzFI71yadF4gYxZP/bebXGOJ
3FxFujgRMpVDQzdl3LlbQg3ALdB9k5abYBHvaFH4hoMbXyVJ+r2rnhawL0pU6mD3
xa/FyOaStKl5WmfaWVKLdo06S/B1rKQn8h7HTQdT3YfVNafJDljBlWIYmU8MnPhh
0YyXI1GG4o2F2KJmrGkWN955bCSSscv2tqxutS8mulkznj64Ovge+NnmImFU+/Xy
Bwo01hGVXAw5FXnHi73q01ERPkPGUh7OFJ43dP5Zq8m0sd3yqotcF2M8pifVXPev
k2tst0Ak5JVmdSdUoUUHDd5h9TTIk1DoN79v7HOEXoQ1TdbN5v97trmxJVv58+VQ
tMH8VfMQu4toX3siMMl0unabb23NFfPD19s4CC5xJDc1wYnkPYJJblf3Fqfwl+gZ
Ciu8qJqDi5b3lM6/9fte0bJm+PZTCU6aMianxM87//aRHZYKfCYCSiznwdEmQYMI
ImdEvlhAVqlUOc7A+aqE6iOAON23GkP52IFxqPwzOGnQjq4zxlXRXyy6Io1sLMhQ
yjYRDhIDXj/Zw6MEHfn0YTzkNdtjb1p2MYDOqnyP/xKhjX1SqBJJcAB99wzjakRh
gKSEokTyLVTWBuldcu33LXVvMqf4A7CxfOP+fuwVLDGgcYcAlQX0qArsSmlJVUEf
s083fDLMlIEM/jJQu71sposaLsPt52zui6PLecnu1hDLwuCHiseT+YNbDyhN1Nc0
fg3j6PqmQVKi9EM34cV15D72JbuPYpYrkOwxLFMrKuJLwmK4Q2dwzPCUGUSfvvKk
bJll+lhHY+W7kW4aBrQJQhHAmdvv/1ljoi7kipA+aMKyjlOTODKf3aqeg/IciGkB
CsHQox4B90KvUHJL5yQ+eyJ1Hb3JeDwUhX/1qHgLDpRVQNpdJZfLonJUvGjLKdmy
d11LlbeRY4Osh2Gfwb98Hl8s4z/3vpU5/28zL0hVSoQdMkEHCPcZdHUfzRaD1ZJj
gWjvxR3kEAieYSRgwT0plQ0Q77sx5ksHUskSLLLgfbAkw3GQgi5TQzWmYfYVuw3u
8aGIx1JRKJZEIq4yIgA05wOcw2FjY4K4ywS/ZklqvJYGidMon/UCUF4HqOBcyg9V
MVTwP7aZhzXDvJk4/4kt80G7zOxDUBwBcy+S2UE/ch7gP/I5Um0318lQk22dlXkx
ven8XTgi3v54qlk0C1B5lZQb1rQS5jlbnbwQo83F48sHSSUMCi6K2SWweKNjxiie
dHgZPKcDUlm9zNmu8ptVQAp0Ju1U1ra/fX2Kp5matxVwZzyElZob3xKqP3j32Im2
mcOUVbhjuTkSnNqLKMf+Y954G5n7eNIEfpAcf4CTP+ApHw4tInsUpCdQfnj9aNU3
QmMf/4aRhhpUvin2yBrMDMJhCDUrFuWjNafxbvRlqiqF2IqSYFPZm3QI16kGZLcY
8j+IS9gKIDIA1Fh6NJNrbKbkWpjPBJ0W5ykgoXnOwSekzmj/aTMxkDVvppFHgKrb
dlSwNWPWtDEaDoECgbsMsNpfqXxVwkP8Lo86+nVERAFNhvFPlznHzMt3uFdjNDpy
Zsf/GwsWCnxWrTdy7Paygg46/rVX63ZH/OUyZTlq0EaaN4QbuCMLn9FykRN9maI/
UvWzI6yvnbzXMUH/3Wpz/NMrUGO7IiY8L9U/ZyluXDJyWoLFeEMKSyN+TOKsClPg
ibuj3pPTNTIAzN76OWgNmmllmBPqqRR+gYhylLhtRvJtwx9RtgS1eHRaatPWMsyE
7USTPEf3V+woVWev0g0bsDV0lySs0F/+RvBd/OdlQp1v/+OgjU64FsnR6KsBiaM2
Ep6UPb70RLABllMd1vWVp6JZ8fMgzwJmMsmDPUydjK87zK2ZGjR5woC1MSmZS82s
Z9ywLO98tS98Y1S5cENbDsre9Eevh0dLhvQNTQifBvuirsSWQdp1rSwT3MoaJTp4
X3rVTRk7Af9NMybjTw4Jq2ugiV6JUd3x42IlkbwtSf1mC3hFprusjQULGGz2Jz6X
saNGZekdq1Q2ynEo0vrOO0nzRA0jAPx3mM1iKz0/udYba8xTHo2KRFZjQGdN4B4y
bDI4V9aVy0ip/DTB5lA8Zn40RdCnhci/n96QenCFtRuZjKp+WjNomYwn9BnkCaLN
/8pwfyLrjgdGBzUSUf+aCOGDEwlqyRnKJcZ4bIYCOcHlxyog6bnbhTRdpcelfx4x
s83Ik69iECDZ85XVtUqgmWk+JIa3IPDQ+okC+MdCVZ8SJuQzmYUychJHwPOM5fTh
0OzPjowQJ9XkXQZosgeKNwu3NsH1cS3fF9jyOZDfjm9lmLDnsN2vk1oyWleHlGAI
sJxvftZUcO3Xc/ktRxO7nArPilGOEeLFY+n6cvF7vEOklLNYZGStZx/K0adJJY9t
62MpuoV8gxNQOi0K0W5jk7NY0jlDNHiKu3Iy7I1wPWNN5p0bGIrpRhP2ybWyiNjp
MNS+coAKLnD1zQaCciou4mwKYBC1NxbcC7bAN+20qPK9BJ61o7bSTCCNCtC1yZ2v
/GSwvgLGSEDGk1LenOX2Ew5rF1SIQ4hFarn5i6tnPU6AzO30NG9w0FgeHdsB7YH4
Vg76DhT+f/R2rnXXwSfeEq7KtAEP7apj2bKFMJxz+wAyvR8GgkvWSgg1AmpN4xFs
wPMiDYYQZQ1iAiX+m1dqbQpbePdeFmieNU6g+jhQ5HAPAhVUGpEveijzj2dOiGbn
kXKb8n2ojo8jzDNBUSJMeoNj2zOPbzWEXzN143lpllf/pCAMTZ8HX0qrvXSwqQmQ
COLSCB9IutBMC379ZYe6xQ2SkTVvTAKLy7TnD/n+LdVeoij3QAs3j9p5fSKGofx2
2c87DsJH+yThIRIO9zwCMWfmAHRRQXh5MZehGCuT7yGClmdQtnS/bwxhHAXugk8n
3gNLPqLTqpWISRC5Je+x4A65pMGkIGqpbPZt5h3DBCD9i1XAV/JfPE1P1euW9hQZ
/8vYIYDCKW64jsqSAdgk8ald2khyepu1cSAGLMWDqEYhxmnPhDaYCSnYyhtw7CdD
WWbyO4xw3paOZDhdudFXWeqt5OP3dUIcJGbuplDtUrAGkcdpp++F9AGsXlLYZPl8
4VXLO5cUsJ+BjllKAyXrL8MFMvFSZIVLo66+yayF6qVgTOwFYYxOOcERy2pCiidB
S4U1BfuKTFyy0T8fWWB9QPWZh4HYw7HFUJYQ3eRGW4fvigZhxuKTH/jhVRiGeQ8A
qRw3sNfq99PzIX7jAZYdsIxvHCQFr1RUrUK2OmQgUXMD5lDLbNHZJWNIAABhPrrc
i5m12vjgpdxKHAFVnbI3ElUBQJqcjY+cDZ7OXBivYZNchGOJEIHClXzGT+BunbgL
i25XD8zfXB+NETYr6YBXeAq4sYSqDZ8oS8Cb/Ew9AQ2ZbVhEy4SAWXcu8Sa4ms86
pDSTqhVpctIQ2nPTkGS3Df2Ny+JHql/t3EQdpEHU88HkVCa6ysOPPlJDKYNxevE3
CESC38CR9GoOPuHqVhDTrrYGEH55n/34BV9c2jB75iIvuIqSJ4ACKIOTUvQ9rZMD
ZHVVbftD2o8UoYxL58CWT5HFhNAixGmWex0tFnQs4KvRzN1DBIXvZpr3tBmmQZxl
uEDc/w1I0UajYPjAw3kBsXQa7d7Ofv7RBV9OBkPz/iyI+57i7d+JkoWhdejox3l6
ZJ/uj76zsesRxWN6KevCLVaYZ3wwwRhty6u37+1AA2vSREZ0OvOW/iQa3TeO6Qrh
qExhgL0SNKc15bJLnV4Z3+iUkchGFm0HDeOvvFwncchvKJicIPLKRNKi47SGIMtI
yXUw//1d66X1wsbzTSaBdw2DTY/iegjqLQibE6lXEta28qPK0D5XEJH4Y+SnJSna
OLOmRDzyWuRz3hbN9Bs07hoHnchzoDNQgkCI/A+q6v7OuMajfqnz5MYGaqpH/lC2
XQhhoF1T5dDrOS8e0G2+yjRFfQruyE1QBmk4ciTAmdkHujCGZNrRDWUPWffpx76R
BDlNrTPhvxS5oQkbc4jyVWkFAzSNcaHZeqAVPsDMVDOcw6QDwR2apF8tOFekLbnu
tGdfCS8XmDiDg9phZtGm0lZwlXzqih1GeAsd3JvemTy0tU4BgJVhXWvG5mxqSeOZ
GklpQhJsjJNyQIMAPdy9j3/I7nUon32s2xM+mGQAo3h8Lnp2u5TeQFxrqkzOGwkq
ugbUUOBg3XQk1rSR7twCQ4PCtuLH4mnElZ03BJJqb3DbKGvbXyXydtFdEQEB9ZFT
s9X5q1U5a4SZe+GuGQttSQ+Mz3HaHqK+CHps7x1SZbWF2nT/3Gi7qoguZEBOCeI9
VXQ6bTlYFr7h17rKo3ViKeSgsHBQ8ygACErYszkQ+PVU8yzf6UHKdqA+pDDx2Gkf
I/9C7x7cmqyfIRCpoggPgTNln09QdcH+DQH3Gd1zWfHgT2h+GkKRGMOpyTKiPUFk
/B+WlrSvuZPCgNqmk41LpZfnuYyMyAklhdoN3cShRsDpc9JkdBDTYRNP0NcKr3e+
AGD7taLBeva3/QIcrmQgzBj3aIb+VuTGjBMNDi8/Nz3cD8YqwHejk1k6o15xqDWj
E8ANOnTsT21apa8jXEWEha1CWLuFcj6NqUtvLtmzgMmMUZtTzcPA7m2alLDmRRD6
75fjKkY62cn+/OKtQiT9+zB2Ht/5ydfPXwQQEhPlSe76qDprDVCdPuwFoLDUSZuF
LjvXF5Xc5lLFE1hC/IUmlzZuWgmhjFlKSha7YW7m6JPdIpVhBUi9uOFdOQWmqsA0
pUPQjmDEIhX5W84BX0TtJzweoQcY4IOUEudC/n/2fInWb9AyvQQRlZ6010TE58MS
GEqeBvwPC2vY509HYctY+R//N7YMj92pn50kMoGUyxuBFjykxInIYdVfyYzhzlEu
epdZzgU1ZbUcVfXTxqLqjamWyZ2RX+oGt64IunffrEnsGX9z5x/9+mfaZ3mN4HSs
vKj6QNBJ2l/EZBX0ZbD2lHUgvYhoo40C6gfML53KE3UtdPR24UT+cB4VjkqJ+C2e
heZlb621S90kdfuVTc/ii2cJIgn72zdeUvUmnkaBdKZlGblgqI3Pf6x75xbld+tw
s8J3TS6Lasii4qIp7taagbfbreCajZY8Ex3V7SPkKeSzUBzuM2oLT125GAEP3ZVc
TIVliiXbO0FBAj89mCz53Eo9oaNMVTwRBS/4181Eg3Rmm7B2CAyExyqFb7hjRrse
ggsh4gBNSratSpZD2ZfxIPgPz5tzh1OR44dx0C9ZDvU/Bfpei5qG9E1vUy0N3SEk
fb4wWcFk5eN30/0btuJTFoYhrC5GfZrxz4jpg3bNuhorVMogTqH4XFQu8vJMZG2F
75GNs0JbtlSFyFQpvvWdVBEmkJRxijGTs74Tjn+Sk1wIK7HTFS+lgdEkRkdriDQr
9DxpC3llyzMHAeM7jVs85NptnjpBE1k9vUEzuLlPN8FrPQarJqRLS2TwqP6pU5Se
d6whqiiOLSOXJZTVgghsemJ9iDLbj1T8V1jtxEerLgB5tMhLD22CcWYft/8sv7we
iyxZd2cGS7XdpdNK7Aif0GfIyI8TB5yo1GsJekckwG2deVFqXJC4/3F4ULNlB9SM
SY7s2Ot37lf3lltSLfl1PfPyVEYmMsZXGuBctrHxNJCc9zbbXmxJCKp+jgnhdmv9
vUB+YvtGXC1m5ZePHyQAnBibWanTwoKxS0XAh3QlSxl6PA9g5BcccOdVygMUTest
pHDHxzk8YXzYdRrbwUud1cLTPcc2aCdakuFAMNO6C4yss/qcui06g22GwaNAkW9A
i3cRDzv2vZVEQ5hXqj5ixOC1ILTsJeFQF7dCCDzU42aWMsh3lAca+pu/XZ2N8o7l
wBHtUBkUN4mEtJbOM/xNqtugIqJnV8aaZg/2WNna2/8Ho0prN774DaY8rQ+8bJft
/tSGXwlBwTXJoJnJtQD5cAhnomvJ6DFaSv2WSmJnKjj75S0OnFvMlCq+3d7Hq2Ax
2izan997pe5IBq3qeMdTPhChGV9HmAjo+njj6xhSEEOLWm9p7Mykyob7bgI8I4W1
OB/c/W1V4nngbOWgQ8vvMB7hfIaqoZC1q6ZSFrLVf4WdjdP4WOyDuUIgahAYBVXr
sfxkIsXgrgM1XMWnPcXp6wPJj8kg//zB8CdV+PAoInJPjY4EuXwzut5iY7V0nhOy
PlUZrcPs9apag4b2wT3OTS+vjtCP1GT2l89SaJqI0JtuKzr4FXX4rrY9GHOaSExx
7BYtLU7jvttgBnB+Ymi1Kw6EOcVO3w63zU9s9WnKvMKAzPFzja5VKZDIt5Nbfgzb
nHcmBvAyylMD7QoLQoEeYPzHVQxlqCcE0fuwo7pxUhbwptxt92uDpYobRvzj8Lot
PvFwiToipw8o+16aLx0/X9PRiqvcuLmltIKH8iEcEiERLa0zztGVSaypI+KRw5Zw
vhqr9WAtgPMiybweCU5x6tDjPG9DgJrPj/xhvRA/NjbxgnqatT+nST3zFzS0+CYI
aw1iuPJ45JHDG36m1ZjXvx0RHyS7uC/cODutl83iYxGDxk6YQrVDdknn1yA+D64V
DdXH6D+VPBdSMoLnVTq0ltC5rPMqd/6uzG1lwQJf2gIgPNufO3ZM5C5ux58Gj1us
QoymajH3cBjCkm580Ze9Nc8QUpA4IIn2+CpmG4/nPyjzzDNyMifa1WvQucbAV1+e
P/7npgx43yZWjsGLGUs45WNYzRyVHVF2lOmr23ohudwrHey75hHEtnXLq2d/iew1
kPykgaXUAxD9cNQ9iUmxpBOsqYUYr9t4Ljya8Q/a4rTGEkvyedZILWQqKF0GZiER
vg/SxMOGDYNgjZ1mSSfKFd06ifPsmreHrcOU4YrVTq8bqnSE/1U2VHYDGcwKZHYD
Y2bgfmVodYTN7Xtf9HOiKko59lHpQTWwnbnY+9G0n6TXLApFC8ov+U0bznDHfmZR
m6SqUWjCjr5QWb74YSh9988Dj26uf+5GW583rlPgo3Oms5stymYp5rKSOtJWG5Nn
PIbCFQmZrNjN7yBrkHGEdw==
`pragma protect end_protected  


  // ****************************************************************************
  // Methods
  // ****************************************************************************
`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_ahb_master_transaction)
  extern function new (vmm_log log = null);
`else
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   */
  extern function new (string name = "svt_ahb_master_transaction");
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
  `svt_data_member_begin(svt_ahb_master_transaction)
    `svt_field_int(assert_req_on_each_beat, `SVT_ALL_ON|`SVT_NOCOMPARE)
    `svt_field_int(num_idle_cycles, `SVT_ALL_ON|`SVT_DEC|`SVT_NOCOMPARE)
  `svt_data_member_end(svt_ahb_master_transaction)

 //----------------------------------------------------------------------------
 /**
  * Check the configuration, and if the configuration isn't valid then
  * attempt to obtain it from the sequencer before attempting to randomize the 
  * transaction.
  */
 extern function void pre_randomize ();

 //----------------------------------------------------------------------------
 /**
  * Method to turn reasonable constraints on/off as a block.
  */
 extern virtual function int reasonable_constraint_mode ( bit on_off );

 //----------------------------------------------------------------------------
 /**
  * Returns the class name for the object.
  */
 extern virtual function string get_class_name ();


 //----------------------------------------------------------------------------
 /**
  * Checks to see that the data field values are valid, focusing mainly on
  * checking/enforcing valid_ranges constraint. 
  
  * @param silent If 1, no messages are issued by this method. If 0, error
  * messages are issued by this method.  
  * @param kind Supported kind values are `SVT_DATA_TYPE::RELEVANT and
  * `SVT_TRANSACTION_TYPE::COMPLETE. If kind is set to
  * `SVT_DATA_TYPE::RELEVANT, this method performs validity checks only on
  * relevant fields. Typically, these fields represent the physical attributes
  * of the protocol. If kind is set to `SVT_TRANSACTION_TYPE::COMPLETE, this
  * method performs validity checks on all fields of the class. 
  */
 extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);

 //----------------------------------------------------------------------------
`ifndef SVT_VMM_TECHNOLOGY
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   */
  extern virtual function bit do_compare(`SVT_XVM(object) rhs, `SVT_XVM(comparer) comparer);
`else
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare ( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );

  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_ahb_master_transaction.
   */
  extern virtual function vmm_data do_allocate ();

  //----------------------------------------------------------------------------
  /**                         
   * Returns the size (in bytes) required by the byte_pack operation.
   *
   * @param kind This int indicates the type of byte_size being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in a size calculation based on the
   * non-static fields. All other kind values result in a return value of 0.
   */
  extern virtual function int unsigned byte_size ( int kind = -1 );

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset, based on the
   * requested byte_pack kind.
   *
   * @param bytes Buffer that will contain the packed bytes at the end of the operation.
   * @param offset Offset into bytes where the packing is to begin.
   * @param kind This int indicates the type of byte_pack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being packed and the return of an integer indicating the number of
   * packed bytes. All other kind values result in no change to the buffer contents, and a
   * return value of 0.
   */
  extern virtual function int unsigned do_byte_pack ( ref logic [7:0] bytes[],
                                                      input int unsigned offset = 0,
                                                      input int kind = -1 );
  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset, based on
   * the requested byte_unpack kind.
   *
   * @param bytes Buffer containing the bytes to be unpacked.
   * @param offset Offset into bytes where the unpacking is to begin.
   * @param len Number of bytes to be unpacked.
   * @param kind This int indicates the type of byte_unpack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being unpacked and the return of an integer indicating the number of
   * unpacked bytes. All other kind values result in no change to the exception contents,
   * and a return value of 0.
   */
  extern virtual function int unsigned do_byte_unpack ( const ref logic [7:0] bytes[],
                                                        input int unsigned    offset = 0,
                                                        input int             len    = -1,
                                                        input int             kind   = -1 );
`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>read</i> access to public data members of this class.
   */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, 
                                           input int array_ix, ref `SVT_DATA_TYPE data_obj);
  
  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  
  // ---------------------------------------------------------------------------
  /**
   * This method allocates a pattern containing svt_pattern_data instances for
   * all of the primitive data fields in the object. The svt_pattern_data::name
   * is set to the corresponding field name, the svt_pattern_data::value is set
   * to 0.
   *
   * @return An svt_pattern instance containing entries for all of the data fields.
   */
  extern virtual function svt_pattern allocate_pattern();

  // ---------------------------------------------------------------------------
  /**
   * allocate_xml_pattern() method collects all the fields which are primitive data fields of the transaction and
   * filters the filelds to get only the fileds to be displayed in the PA. 
   *
   * @return An svt_pattern instance containing entries for required fields to be dispalyed in PA
   */
   extern virtual function svt_pattern allocate_xml_pattern();
  // ---------------------------------------------------------------------------

  /**
   * This method is used to drop the transaction if it crosses the slave address boundary
   *
   */
  extern virtual function void is_transaction_valid(bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] min_byte_addr,bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] max_byte_addr, output bit drop_xact);
  // ---------------------------------------------------------------------------
  /**
   * Called when rebuilding of a transaction is required
   * @param start_addr Starting address for the rebuild transaction
   */
  extern virtual function void rebuild_transaction(bit [`SVT_AHB_MAX_ADDR_WIDTH - 1 : 0] start_addr,
                                                   int beat_num,
                                                   bit ebt_due_to_loss_of_grant = 'b0,
                                                   bit rebuild_using_wrap_boundary_as_start_addr = 'b0,
                                                   output bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] wrap_boundary,
                                                   output beat_addr_wrt_wrap_boundary_enum addr_wrt_wrap_boundary,
                                                   input svt_ahb_transaction rebuild_xact);
 // -------------------------------------------------------------------------------
  /**
   * This method returns PA object which contains the PA header information for XML or FSDB.
   *
   * @param uid Optional string indicating the unique identification value for object. If not 
   * provided uses the 'get_uid()' method  to retrieve the value. 
   * @param typ Optional string indicating the 'type' of the object. If not provided
   * uses the type name for the class.
   * @param parent_uid Optional string indicating the UID of the object's parent. If not provided
   * the method assumes there is no parent.
   * @param channel Optional string indicating an object channel. If not provided
   * the method assumes there is no channel.
   *
   * @return The requested object block description.
   */
  extern virtual function svt_pa_object_data get_pa_obj_data(string uid="", string typ="", string parent_uid="", string channel="");

 //------------------------------------------------------------------------------------
 /** This method is used in setting the unique identification id for the
  * objects of bus activity
  * This method returns  a  string which holds uid of bus activity object
  * This is used by pa writer class in generating XML/FSDB
  */
  extern virtual function string get_uid();

 //------------------------------------------------------------------------------------
 /** This method is used in appending the transaction count at the end of
  * object_type to get the a unique uid for each object that is getting
  * stored through PA 
  */
 extern virtual function void  set_pa_data( int beat_count, bit transaction, string parent_uid);
    
 //------------------------------------------------------------------------------------
 /** This method is used to clear the the object_type set in set_pa_data()
  * method to avoid any overriding of the object_type of bus activity and
  * transaction types
  */
 extern virtual function void clear_pa_data();

 //-----------------------------------------------------------------------------------  
   `ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_ahb_master_transaction)
  `vmm_class_factory(svt_ahb_master_transaction)
`endif
  
endclass


`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
gMjSraJDHTETms0RseJJ8EYuBw+v/cnWWDPi4dyckY+m64G5GjOgVLr4sTe8HLxY
6tpUfr9Pvrvi0tvZx+hXhuC9k45l5botP+11vUE/eE2KlDBzctE87/fmxeKDMzx8
QmkUUWG7XcEpybAv7lNhbSkus+rMjGPvJ2zq46gxP1A=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 9703      )
xseTgp1lsm/yzuSmyNySv7mkvmRsLRUovuoH2VeGxo2PxHHuwKC+l5OTEM/hXZYu
ACEeMnQZx2zBH8WBjISylcrstVsYFfbBW8tuYc0c1OSsUeAseE2PuN38JBpHbB3G
Mn6qWNosdfTS/VD2FeynkF/IFUP2J2wiE5X3YqNaNaeroIyedD5785cbV6PxApoO
r3JtsJB9N26Oio2zqKhSSUD7l6t1RMDt4utZWkV30M5cWzfEKhbKuh6IgjHXEZ0X
ZXnBLmd+wzN472awMz9N4jvOlmVG/hTAceQfKNdO/PS/XdnAV6jGYs2HjdJJvekM
aB8zFLMo62JqyxBSOvmHIKt+1JehiyQClxHGxqjmvqqUhwFcdECckVf8LvHA1rBF
725ooDlgzDME2567PCLn6aepYI0qC23O7H7Y2slo8zK4WSRWto3pmAkqOQv8tiVX
y74waikoOaIUa6ysMNiZYKKia74z61Ovf+2xjtiyzUm+e+zuY41gGTYFaL3pkJfJ
9b0nDVuX4eSkFK8yvPFstk7tmRMTKmuAHKAZZxPU3D3EmpUuEuT0Cxp2gwuSKd0r
8bL/n1no0gu5fsccQ4Q6peSXireOzRxuXpYuq4swApgJ59gK2OlEXvXWSnBJ5J3C
2MLvWnf7jyLOlzDSSCzcTxahcXp5gIg34qrfo+W4YqHUPxkjZNfCTXH+Iz1ikIEZ
S8i7RK+MnhIl9lK6n8TaeH5rUKq+7D2N8ZWhwdRvi1VWgQ7PuAgs7LvpwI3EwWE8
xPatCeBBlqbCzPgxBWQm2x7QK+rbWeKvfAszJIRnCMx8PckRtS/Jvw7+YGjnTjYN
csEDaxyagSX59KiEm+3Jlp4RJR7Z5+p8WMVt1O+gnA36Zaz1OuODEOO2y3okcMB/
35VKJrvhe5t9O+0Gh4dWLzS6HJVjImcWXSBBsL35gCDaD4AZETJBaImSPV+akt7I
H5hXWOt7S0CD1zceBU6J6bGaKc/wZ+C7aXTMNSXiyXLohYMoYfd1yzbJTWNmpMx7
3zQthUxv4hjWc523ggHv9zQc5PJVvTNWbEE3ClxP4SR2uepGK0OB4IfIGReb6cvs
cdXK2LecsjAKIsmvi8xowOOHIRlrq5UzsFL0ZFYlMHyiB5YDgFyp2FBAruDhO09n
1Sn/nL6sebzvD6cvVivw6VeUmcaQ6CqmLxQ08908c6UrCufnLDFfdVfrNvIcWNcL
CFeRUfE8+OnCYXoIlhB0PizX49vZZO1kYa0i02rL5CDwEBOZPqPe9rGwNPuOUIK8
pCi7v8WM55RtbEQ+VA4iufzaSwSNyKTRySm6qlw8xQnzUe4Kq5mRrkqRS5bbyZtu
zMhx7zalLSmQt57Rty0qcvf2UTB/BekY7UB1nNDQ3ZjI4Pmehlx/Ylq9AkPnDdyJ
`pragma protect end_protected
function void svt_ahb_master_transaction::pre_randomize();
`pragma protect begin_protected  
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
b2fbrAwPLPG30oxUnkLDYEPSLh4tNKes0D32aGMjyplLZCNBjHc6tFsiTi0D4CYv
jUomPYqkE30Wny59YDDaXqXxAmiJPrWApfgTv7Q9rb3ULuwTDlpHPUaBOYNIH9gy
bsOt5u4eT/NU1KwQ/+HbscS0VFvhDKTb5CA5RVVAzXE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 10348     )
EeOxIX8fGZjtU489IJFeWhf3ez/dATsDKdrLTB8WYJryvZNGt0OPvSAQxrKgwwi3
r1HxGoEXg9LqAyaC2yxaFIngak7nPVgWP27sPXGscXu7L+0UhWV1KPoe4vgFgxbW
K69bwxC1g6/5cL/M2s7M7VUIrskVL6jm5RiaF2dJzgujEoFr99RnoR/xowrKvSvu
tDR4wOiqq/bWk2eC9kKmgF3ZeXxN0d1/f1sxv2gKCyxhunj7MYm6XQp300iWNYSA
RVoIQWMTMec56F+PeherThgsPLaE5edRZZVa6nM5Y9qVkhy4SGdHu7pLeTwAGgML
oFrUGRBFYn9FOgufpboQOKrn15U7YbWuQXESd4jHO5DJxDsWq1MxRKl54H8j+kOc
DzX9IE8NlvABH1c9AC+pNhJbDxMQyzZBbYtrOY7SdlSO5n5D9chYc7gjZBCgRFuf
+CXZu3DXahTrHa+Qz0/gTccNiqc/jnYK1Nmgt1zA7WFxXnE2YFwWuvMrrTOyD8Mu
riyodpGVCPXRPbugN7hkP3vO2xFzdUerccr+VAs3ZI4q/bUsyertiM403F92egin
BZ6CLB/64nAcyRpIGYHKmrOgy2lYXCVKXaMU4KZl0SzUTgR8zuWx0NmH78+es9QD
65bRCbl1nLK34seyVuJYrORPlUg68dBbaSK+UvG6swRLoA7HAeHp35Xuroya5wKo
lmO3pQqBWw78LRoufSfmULiXyL9ydyh575CdBBrQhqrvk+1QLvM0zklWzjOSmLUE
Xus6MPPSUXuOBBLfXcWpPAYY9hhckgLBZlyKjTkNUIbIkBc/x6V8Q8nMBTZUsBVn
Bt4dbDgfYF87zF4uBRH+kMI4F8c8qJI2EJLQ7Yrob6g=
`pragma protect end_protected
endfunction: pre_randomize
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
WI7ygjsO4BFtdXbk+wKxUui7PKtGlE9d5Bo4KXPVa1IjvLYQwyi9YPFnh21i2LiW
ORXEVnfdbCbvgx5/2k7fRCFD94w9KgS+SKlSZaoTJVxvj3qMc6INyqx/Vi0cxIgQ
0RHW/F8jZrethveyp8sXkvHTlFYqVLsAQrIPoT8Daww=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 33843     )
lzmvZcDm11csZMp+c+Fq9b5twr4mi9xXWoGNpch2f5ulPMWbPClplvL+cu5ZxzRT
bAuAdap0E+KnP25J/1pyY/f0BqzifdV0XSB4uh+PMbF9slR3Uaq2WCjXBeNTndOD
no3HrxcLwpOONvxG3JWZao4nvcwMNPx0tjOip5EiSlgo9Yuj2Jgg03ZZPnRnCUu4
1UTzjjQx2zDnQYqH+d5q3CwUBQHOrq0lSjFNQ+ozN+C4ZIOC55Lyjb+UQ+gZM1+8
73yadOe7StSRsOKjWKMsJM7Mq7UwonOeBwYrO2a5NFRi/mnwujfBtPSqE+weX607
6DLo56LwlgGloFn6Id5fgowALMwIH0HZJomEpwWAF/FkkriKfO9EwygafR8/hpI9
gv9MS4Wzxi1Xz7LEG6yLEkB2rUOVkqtToEH6uTMp/oH9MoxnNINL7DrHsgPmOscM
HKdjM4q22MS/TunxwQ64hkPyZZo/fqz+yHzVDnAO0Mefi5W3ke98bt+xVPEnnejs
YPNBO+qVl/13Tfqt2P6dcBN0bblGeJjXpno1loHpJn0jYgwcKAIGMXZq6h9Zb5LG
tklfjdW8Hc9hD0PJVRKqGAW8Hq48r3zn89KG3N1bR5OrsALPfb0Z8BGkAIpbAesO
Jjh1LxkrOc4UAhWCvvAY7DwV16aPe3uYCMx+kdvNcGoJ09MfKvzF+mZhzV0TEnUM
M48YfbKjo4AosY3JUiF0Tfs67e7h7XQPqHvhDdY7wnSTmYk7DnZNbHjH/xfE9C0p
m7OaKzsdouWidpAmb6pXVCLw1MZbSRFCQo3XxcTxkcFDuxvhwObGLnAeuRp1eFJd
ONMDyfqTLSObRuUqgm39nWr78PoDUCzuep0yeKiBTVDQHSHMhNH1qXMaIDeS48eZ
fkW8l6f4YABuTZqip9JteRAeFhNyQ2+dpoovb9OvJmBvablZvaleIZsgOLXzo8sz
R938/pnP0iRC6yv83nDBPCqYrn5aFBFcFRpmthpfj0dCxY3EhNZA31aVu3T/oGGI
he0S5cp/mO6oDz0UXcUU3nNTu9Umhx49XbROh/4fKd9OYJMZpT2basF/aTONBjxC
Ioak23qICrbBknK0Q5TWFMNERCkXl5esr1MnEVIRYHhb0HiMIUvlWeTlt5JhaMKh
vFKsIfH+Tfmk9f4G0YVJGava7O7gNawbzhBH5rcSd+51nzyEDUWt3JPpsXwrVMF5
PrKE5UxEBz7HMCTiaRRfC9Q1jm8Xjiqne0N3+Gz6dykhfDAhIzqnUnWS6bIyo96L
N1HgNz1E6+dNBJ+8Mj5Doo8g7CYp7iP4D7ZFXH1Xwac1+5pcQq4qT6s0r9RSEE/4
BuTNuHjGdhnhWWJK9QDObGZBHlyXSWjl0pg5GpA9Q2lh42R5HcPG3XEEC48cTLnM
NUS5viid3K+PwQ2p3K3JZWN9NTozOvtWw3AWi/H1/Tp8I6C9r/QUnel8yDoGV1B/
hMxJFHTAYJZSVogBZ8lclCeby6rqCxtbmMa6oBhljkS8I9zvXvd6ebbynYuaLe8w
vFat5mey8JEMPkx6qHtcqQoLZiuKWaR98uWAWUEfNDYN8abC9UjkySSWB8uxYoc5
hr8IH1FTMsdmsNT3PzHhs1Xndfszo9ZWSEoS2dTe8J7NXIPF1mEhCGeMjJJYxa7x
vX50rb1377QJY+plKgaKth2YbyKd2sSagdBNohzm0lPuxyxG53/ZWoNzTtsTilBh
3zhBlKjSgyJpK/O9Bxic4kpMXvVgXi/NwvyCbzzmEd6CJqc9qI2qeF/4p4oP8LSb
y7kUJ24fnmx52lX9JIiHWSrZw6Qz/7jLcvk3fjvAHDX4bymjF5KXXotSE6XLqzaN
cF3bhSComvCq9OUUz5pDTrtE6SIYZJuaxXFhCggFks9ONCv9LJPtExPsAuVj+fQF
XMxNlM14lrlhwzUNw3xMowweWljJ4ujA87vAmXsCRYy0BDgkwu1vHfYyAn4ifWND
NDa+OasTGq731DfVPKkHCEoC5BXWZzm6upeAAx72/jMmae7h6dJ9CuR365AGbMmE
a8mfsoPheszjeLtoKCsGi1OqvjV84BAUruy8fF/iJ3rT9h6hCHBrFzhSeGb+R0H6
nFjXimoNsfiENyxYd/KMen9Ibq9SZpZ2zkqgx/TUX1XqZ5EP8afCXf/nIrW1LjkI
H4XagGZDGD8Wr21cqDVA78zv7XwQ1VDjw0G8wzz/DOGQhroU/lXQlm33DiT2GSwi
Ane20UvHpjaMVluHSsLs6gnPfTcg1SO6ZMB3VrrYaJrZVGgo3NxzKHoqYW+7kmus
qpzAMWrNk+pwQt6IfyldXUyIsIlAEehZOklkHUHF9C2vcPdUdlmCIOJy6dSy7FRi
DA9XN5lK+Jg59xw2G0rBDXpT9S21YGKyei+Ii3l88FfNOJ2N8a1tvUylpwZWhJMF
5COq0FaGJO4NtR69yswfnDwNlauP7Lk1MfCJc0MZb+GjhJsN7+DbCNNiHpqjehQa
FPsSqBXa9CrPXFqnDWcXSrdzZ1YpIiVhY7bReylrtJEt+xKdfDAFGFRM3i9QcvYR
eSHoHYQc9JiBA6TsZbm0eqHoqkYZKJpTdLXYtyTBGewT+auvopiooq9mHrB8pEn4
pB2LXp/i54+8e2MkrxyiU5GoIuPVtZ0913tCpQXS+kSRE1n0h0wSM4T2v4mRsDv5
u9M87qYnQzf8rds0ucRGQtvPS9eleorxKHBVJWObRq/8ViRnjWETp/5bxKuouyzn
VX5fclo1RaS+Vct5AkkN0iOSXy7doOh2HsMnguIFSh30GYtL/F6zwSDk+hociwta
CxzTRjof6bOiXuYa8jU6ha3tQx5mKNF96Q0PV5ovHdLJo7HW96IXaKkqnhmOy4BM
DIWtHrTkgtZMr9A3cy2ql5Z9vc7UVvvC7WUEAmN9mO89thHWMsE9VXjASFA/ALzw
h9XiapVDPhjd38SWHofJVyHaSGP+/fpyD0AtyYrGQhpa1Ta/OUp6PJTQsyt8SLIi
lP5rT+KpcP9qVk/eqAGrM1zA7vuqeR1O8EW5j1PkePJA+D9Df51R5e8reee2YFEy
4DSOEVpdhZTDjQbDJDNFnIYHX6z4H8QoZQ4qm8jsz6IQvxKfq6EY7yPE2vUCDWMk
87PuwJ215l8vHjwNQkRg4tffoTy+ul9myc9QU9gOENdgO0E5wIbfvE/S/2LeHB3U
RrdpFwezBiChLJk5yjOa4asLHpxNKTDkBwXL4MFvvJCPGqQIkGvx11hfIe/YxAvj
3hAJ9wWgMRJ3eiK+jAUgIFSnrmZhbnf3ieFo+09fxIEMt0Jj6jTPLgjqrPhnmWkf
a4bgj+Ud6oWlCb0Nn/gQcbXxI1eAX5rnyfrAa3uNG2MAf4fGXlzI7Qp8Z//+9FT5
dd3e5jS4KDge/MTTxA3QAugkCnX4CwnOfZHb4QNggr2UgEsowZZutPkqrhPs5e7Z
Pb+Q5glpEl0GLiIxl7PxaeOM/k/CqLOqcsb7BGE6bBjU468QlPjPIynYxt77D+zw
uBxOQn5fysdMfXLRpNRZKUw7ceSxXlOYp4zW4oFJhVbjLclufSkwaNccCPrWN78d
F9p0FkVP/jVfTzGzX/eLXFBLAIdpyUIV9RJUJjKp01zoAkQkCuSfrtp0+J0OZldh
sITq8DCDsAqAV/uJR9qXfFKdx5aXomyIgUT3h+qZ4+4M4NtBNCYYGlGsdc6N5dlO
slzXt7zRQ/k86sQW0Y79V58zjfOSwdIxhjAmtJREzvQtnFp9TnzgkaU/d+0c2Hto
JRtzmwrXiAz0ol694C0YG4Vv0vUdso8H53llA7sU8bx/y+BzldaUOlYn1hKUSOyf
VnryCg5ePL33RensPEdpob+8tqGT1UiwAonP2h5wJHAOI6meB6x37XtovPI73LA4
AmHFFyFbdoQXQDhTWWYIMD/Y9hh9Do5pkc/jHIbca9dTWcC7diAA2g5SWedemV7O
JIxMS3gAv+3hyO7iDDDJa6ZWAE+KHz6Eas6W654FdI9lnby2VqiAjCUA0a1GHARp
/L+rFPXNvcO0KgG64L61zQ1hJ9xZKZXrn5nt4gGAb8PhKW/ODti19S24t2I6t6tQ
vWPDl0/uEBeAnCAYlJ5H0/b0KwrnmLpl0MTpfaOkveubLwvBlUmcKSK9eNmkL3ZX
Yu6ARbRvgGfGXq/4eqb/QIPyj4tbHUK/9mA5utI9mqOKFNJESLczDdqnYnlnO2hV
LgaZZ8ZidFtupeLkl+uQoJKQsFK4hmBlU8uIhcdL8qGOh7IAzyYdA6i93iEKcqHh
9LCOWDGAOy4y47+wbxTYYZXxt6pznaabhm3X6rflikGUHKFm1X5E4Of32XfNrhdL
OIFD1cOYFng+mycjxrWRHDKeT78/gfewzUyEsJcpZqNNgd5VFj+eSygusGz5/oba
WNQm034Q1Nyd4GNMDKzRgTX+r3tN228ZF6wPhL/8zmkCyj2pa0g/aP5eA8S0FiNf
OGbb/elKNF1SHXk7X75VBqOIsdmMG4iwQwJLfQfMVeiTFLxIwTKqGIC3CBUjL705
hoqbog4f9aG2e85O62vwLsOI336Sq+xbtQsSdjVGgs7n10G5IBCuqKe5R5h4WmLi
KGxnMYhInp7of8yDYz7/krO02nIdnFfSVjT4VpFNOJ1T0OLi3/ls5tCL5WC2cFQJ
5VtO6MgrR3KTnjxLpIkl5bvstXiNynlOdNVWOBtUeq3sRoUGG+geQkc7FS0WN+Ut
o9hIec/stO0sey7CtbSid4kMo2Zr/bPwgc/OWsTbbokA6PM3sgl2+f4odKhkulfZ
evlRxY+V9iPvM+tZsv6BgSoKRZ3kh0/nKodqzC2J+Ylz/K91ZHh1aMmVW4KwGAh9
rNObDRJCg3aPPmn44vHGkfYVmecdqLUfBGymzNcYmRLzcmZ8k7qIhT0USDYXS09J
qUx74NjtrHSWY4VNpbGVLyXE0zyZpQX9pLLrvPck+L9tvsExE3PWpJoiZJ3xo2/v
Wdg3tVrsDPwpd+IxbrhaBZcp6bO6TcbIdiG9ohJywJuMw0G8hXLiKuEjAxpKs6Jk
CHwOmGAxASI7LHa9QaHjtTT6F/TmYVGYiFGtXqHB2frEIjsfml6XlRUGXtP6Rnt0
IM8btINj9MlQsw2IFjeR4zBDizWeYBxuWi4tJDoGFnUg9CRzqqvIh2S0TrXl7J/V
f+Qnz1IyTV5BqkWE9UU2J3y1yT5sTIjTpq0wTApsF0iEYcCvQm5VQt5Li/bCZT7F
wQEbh1S6qE/7ek+aeGC38k+kcL9LeWvykSVtPzcO6LSVP3LDtH6yG8vn5XSDfg0+
ojwX6B0+0I/RFCybusjdNuNjqm4rswtkWGMlntBwJCIDVGNxHxn9rRhCTMH+7VGx
lkAPPNbJGGQLNulVHgWBLfqiRzzVH/2tGBWE8svuR0eREwrsFeNUmBnGRZgwm02F
UcZhd4lXOyO+mKXK7Lb67S+KHD8Rt+cy37jrCgaMGv3pwo/Yj4L+xdJinisTzzQS
p8u/hDIcwIdFWp7dPMr0IB1CKjy+DXc430X1isGQUIw7rouw3yyCzU8jeN4vp/OP
alkdeD4lb7ZHjrRTxwD3VnTTfMKJUg4c9OAP8cwPgMhr8IL0+IFH4eMIQCkFY+D4
NVu389pltlOQsfX0KW0d07hv8E2k35oQ7JDRiRTOajtpMoyBBJRKBHWHqOd2JFEs
yej1IMQH7xZyDlE5u/faWvQdcERFaJUYasG4sMrU7I5J3PX2gMbrAFg9J78KX1ag
lM8X1V4pzVeircVrbFePCUl69IYIIsHqwNsRr9LJP5BzCRFSlGMLNLzPF7CrdVvp
rTPmKvqC+dQKBt1ZgqCsiYGijkYB2W8hpH3QZkGe6yH4VG4vsR+pjmOID813V+D0
w58Y5c7e25CnFA/2MvOADIEj9+e0CQvFotBAAO4F0ltZvyfYMPn3nu8Xx89cY2MI
GIa9LKtkCUcOh+FG6GEcBKjBP9l1mzDMImnSife8zQYo/1v4KNhUuvQBRUz7kqic
/7Q5g3rOR+6vupqusRpniXpAmNNYSl811zdcCkHAkBiRfda9lFnZAgDAi6U9FiH3
7u7unm9sC8Y2faetldT0rfq8NRVZ0TmAeKZFdU4qf9UHYV9BbYQ8NtduaJiVlIyd
XgRfQfimbV6IYifd+2R+G/mHn8TXRvNJxSxf4EiezQh3QyUlFB1X8akyUB/lWni1
HBk9TPPCi2LG7g5+dV3pPArwGxOqFW2E4AmqhUaHnRi57QFtxWnO9AslLtR5Bwt1
NwltFrQ1TMuIR1d2Z6Cxju/TDoeggIT9X1BeCo6N7GmWiM6HIrIbj3JupMAaYN8F
YDuCdREBBcg1x73ANafObwlNXVadJnMtKCKvYgvZPMTqOy6McK5R6z2D40Yq/zDx
HeV7HElKAPTsJRG0584+BMpI/jng2jm02xtzjqARABABmNUZwaNs6H7N2I8zg0pH
CigvIs2oD0EdviRjb7wLNz47r4iI9TqxmqwAbL3+IF65Hu9IhZ8vUwtk5NgJdXGF
HYMRmrrDgLAC6mVoCZvjSabpIoo1zsaL3olF1El3LgmGqcd+EoAwxpGBCgdcZXva
SqPi8P0KMW67Tx6xInInodt+9AXSGJMIoxWlj3JMGGLIXwhEXuHWwEfVujOj7cTH
yJ51nuYF2iTft1aC7LwSCtH8M9I46qYwT8gkij1u8sucxrF1dppBlJ5b5mIJ7mck
M5221qljgwvz9LHMdmeU6HKSNqV5hJnFCm/tJiEFQZbcSSxZgM6nkqsGb2iZD/t+
D8BEEdub0oYvEyhcoJEWoWyJYNseCAlv515N+3qXM6AhWMh7qwCRJM1De50cSBl+
HjG4aYz+oWc4cPmalHcD7eSBCUy9THC6AEQW9y053dmkx39ydlV4f0XiNB+OtG49
HOHOdGsXMz5ZHuw+yz/NwfKcxJtu+sqTVwzTBzw7TBWLTNUBBKIHSLuQ3R3kEt4a
rpXAn1kv2zNDj3SzRozWIL3gcKRoeMRCTT67nw9pL1P7hUdfzatWCCFCNzJqVnec
3XBRjR0UOE7Hit9cTpdcVBF6293EEBYGzDJIMVeB/vpn/90rGFJrxyUZjTuxSCbM
WUeouj2G/dY3xueWMLi5iBBHQv5k+qjLnIMMf59k3LUeAFKAqlG7/YV3dYFP0BXW
8FHXfM3vy1RZ8HXsJY5F10Yb424aWD6UGzwK3VJqSiiOEYujDSIIFygOi1Rt8n/x
J8Ohu6sOOaNvrfsff2UiG+j/KbyMuiA8bR3lx6xzi+eWDCglHhnyK5NRCX+M9NJB
zlLdonkSmi3mvJRYfegjffQ1WhYaSJTP0uhSDbx2CpCuZ3+BpLroViQkYluZoq1q
vyOb1FyeXfyO2CYK7+tkR4CmQ0bf6GA7XnZV6fWm86D00C8sleOoofR8gb6ojakY
3CfoiyspYJllVRf2ePCvTGIDnNsB8sMqyFugSVS0LTTSQU6iPuu0/on7sbue09s+
AQbfkph2Y0xdhezDeJGl+X78ZBOdzkm8pDe5A16m4jm5P1h02fXj6/0R+LU/nkX4
uOcoeWvyhjUtB+BHx07T6DWDj/PxXzb+QzkoF0g8yfd4nIyUTImlTZSoFbXU2p7E
43SmyrkvjYAsp0o/mkqKng/2CmhvsUXREpFgzI+6BLcJLxapTQkU7uJcbROjZb7C
FLVTFV2ICaUd6anE5F0JbNp/iHcPZ8tdfn1sS1/D5/Ez4CTz/zCagZdnkZaqVk/e
I5kzt1azr6/VANGTswYf3PM5lzuvJ8EkWDmhEk33y6m5fry3ZdpBLWwP1f0mxiqI
9zZ/pnsoZAsTMBfLq/JxQKZj8diKGrEH5ByFeSnTYqu52bt1msayi8m5rav4ZuU1
7SlRA0vJC0CBnykGyOiiKRg7Bl+JSBiv3pT7vi8vLpSQRpU7rWs9Bs2XvtgfZJpN
Q8XcalTkn3n5ABRQWLINBrxlnGzNHsHoRMbxTsNXvaSlQmlZHWy/lui9xVCHzG8F
OWT4IiBGuxCLQMLfWACPfHmGgLOfTq5Fd9OzOzfWyDk5e73Ktrqbkba5BWuuj6SB
cE5ioFBPX28IumEu3NUWfaE+zdd03VXjyfOOrrix7pLCNlY2Sz/ORfCgit/8aVLe
7s8TcRGuti1c1YWL3WwhcDBLd/DfTPQODPw1mS7KQHaS2feERlVyXhBqXrlMAxlk
viI7eOUmN3SpATJDKRkNpLoSMOH8XpYuGjI4tFPqE3B2L4U1TQzqeqw0j9Sozn1P
FCNpV4XkjKU1YGExVa+fyWQmTgGBMvdwI+DuAacxuVo3edt+jKDtjatCTUw8J4Yn
OgJpUu7fOhJII/MFgwc7uLhQV5AuA0UTKU6W5jTo7f00ctBcWrYU3tnGl49KBody
IW0pT6nPWp1JKxjP55paMcvvvS2BjY+ij3s3v6Xn1vkmEZRbdFX4RO+CnRt1gajC
2ICX10W/yTzna/5dWZFVpZ7NsEfEGbPJklFRoe0BMdaPEZVsHqYXY+iq4R4WCrap
/5Q5j7F7yhTF7aEa0kedn4zLm9fQrwGJ7NUFWlJYiTBwnpHgfTISgF6ZU4sgh9OO
3U6V2llW1Wnt7agOYPqEs/stSQWZn/JeZnNJjrEhnol/NszimC0ItkJ3a1zIVSkC
7G8NTjMt2k9hfavOrdpibDPSb0HD8pEA/WZ8aWEX/wOcf1jUQ21BAGFh6u/gcPz/
/vviml02SmDFHyzZn0XG58gAUv7dWpYVUqCjaay9BJ6CLnP8707RGnnOQz+L0jof
XmdXY+9dh2gIgdtCpxvPjR8xGFxhOqKIuU5//heWLJ8+UEed0I3ZO0iMSsorL2aY
DIBxIXabUSbDV2eMe4HGAVBBfQDVD7IUZmBp6Cxm8LIhiqGj+QyhPaI+8s03kLof
r0c9Iti3R7oBT0+xAWkEEyZiRiSkRfwViuWFvR6Y7xNupbz1QSIop/l2GFXtIgEv
JBeHxtFX4qw0gg/BySfAwFw4VWP4dtQetgSsP778idTreqgsw+R5CXn3uGFgQbZo
/R8n2rM+6l8xlHB6opF0VONBCL7YAOs5kfCAge+2Ox81X/pLBS2KKu9nkCGv4sNp
Frqet39pP6G9+SJeKVKb9DbSU7f7+eIykm6ZASum3KRdssGg/9NKLXFatCuKEdTh
enjd2oC296wioS3yuFByNX+bC/HfbbM9321j/G9uoQi+30ITqK5CVwmEELQ3TCKu
VfNjY31EIiv/a5tZoTU/J13xGUWGZ2Yd0SmvMRWpzhQh4uZUKJ7guN6cnR9LVlTX
F1kUsQJZEAOCF8RiKAz5ebsW7cwZTDKkKr/zfmfhYpdnaI+WK7y+1k5Q/kMHxMLK
724sEcXL3MA7Oq1I6wIUU85mFnU4MbFJvlT1fS5KNzAZGpOZR9a/UApC04r3Q44N
MFsqXCsLDTEVUeUJOedMUF1idoARP1oX1fyVhAn6X+9eAEhkEgGiWy1B920YvbYe
tlBninpatXnXzTuBBc3Sl82BJwnap9RH0V5ZZ7WoDFoYXcRmCHkPnL4YFqkjau94
7EKAC/3k2qvBwIAp/VMBTOt/v4MSHGZO8hA+B24gSsyM4yPRcGzw75ZtVdAV835D
AgMuAYXlKorz0YAXqEYKDk1107ghegjrCP5csnLWEwOQ9QLewf6qgCclk+g/BXrJ
Y0qWCIhWCZ7GWQA34GM4uaDD4LUKyFSmhWe8HqfcGZNP+S27qDrJIi+ycA2j7LAw
Uyd+6ZrEyKLg0+hSDnY+RDzqHGsVjoZucdnHXGcifLlHJXRpbyFw5DYiiPdU+hYs
JQDGItiKceQl5TgA/QSJrwFBcHOs4jcTwb7SO9ZLDQbxIzZz9na5hDiiWtrYcFAn
qtcrpxp6Ks86pjZZQL8lejHdEhKR6O7lnpq+R/jLzvm0UV61EGycN0Yn9YLP4W0g
ps5bOzvCgkk4uHSbn1NvOUGdWMn0k7nt69AU8WNDvgPZRYCvciwpsoSwTfldr0tu
0UxOf3mdZkGRjb21EbcdQ9rqU6qur8GIYkcW5KLjR45JRWNnirCbUJUlkADNeSPF
bUoI67qPSE17NBfosi4a2mxlCbHktPelzgVhMM1O/uCWWxRW1lzJJu//bnryXNSu
CtxUEntDhQXtWNYUEYThIGKaNdmsN5dzgXYE4wBHdcH+d0iw84LJl6ZKERuCFRMu
EZzoIkOQavHmQqi/cdi63BlBZt0+hSnQXgy+0twaaWovSwd161CvgXkGrl39fgvK
brMGQjK93+DCBURJPdSfQCuSU9S0YHrnCBeb6xstoaNlFCBSj4atjCa4MQkghAVq
JqyUnv8W3cpJ+uxJq79xBc18eHOx0LSfBn7lAu337A6gNzJIXj8vc7gstWjKmMM2
bbmqSgcyLy2htmoH1KFqhcByIU+A9+nRVzxofB5fejGz1taXd3tgBxtAZG7X87OD
ux3fmsp8G3O59dxongLzhSGfSkwe7jcMbuEfXoyFWrK922/qyd4XYNGJ0zLD6m+h
8MIepjijPqbJ2a7RXELy89BsTAM66ftEHYamCusExPNQgKu6Ab1rvOUbxsGzQpmb
HQKCqbkNfzWEoAkA2T7mIEkf+gwQO+BPLWntG17B2spVtPJjw5GnlRnKABzs9LP3
bVIcg7eOTwl0o13tydMKF9acL6P4pEu41NPnsIudr1uNElUAG+Jg2ydBvcRJsQ4l
NexeMgExHiCFZYxwBYoO9GrZqJKUgZs0qbnjW4FkWxITfApfs37HGh7GcxWL3SVv
enyGdsenU0OWGxeWaw7ufu1ybS0w1vLI4aP3Le1oE5ob5jOEn+swX3LNcYTfp7u7
r/2Dz7DMMx3y7SOr+bHRC5isNn0SNZfWStSxTUaFSb8K3Rx5rag1hIfgSJ62Lnsh
kjwX1WOQ3p17pOtUdzzTCBO7Ytkd2AAue8kR+PuAXF6yJ38+gaiZz70iqmdCxyVE
6S7OB1a3M7QACgtkXqw19KvZjPjPuuiFViKcHsizsckRtntQRRnu7fkLtw1igz/J
jaUljQpRL7zFdwSsGdf89jlkA7y0ILoye2VSNmECuQb/yAmFR7ehdaFFyHF6u/S/
KOLfpKSEfgeXguYaZ4s9iZucyJkgBUBbgRONYrSsH3OQ2sB3WOSt+vzPyIGB7NdQ
nsp/StBrDiAX9fkolLaSaUlZUOvkrwN0mrxlbiiHcZkegQfwLS+yFW5V3kooHNif
ndN/VohafEmFJaEY+i1JyRC30M7aaBga3svRhyY7rPOXdUE86McQINbEKwFdlCGY
kHXjc6olGoB3ofYlxBdmrCS5d07lYrTd5sbhzJmPyMViA0OpUlIW2jV164NVkXwx
Td1srI0ZUDbf5yoDgUMSh73WlgNpJZRSmd5RIyW8j9n2VDg2SL2CKO0+lHC0Jqr+
VKoIy8Eg4Q/w9GUFXP8Jy1d4AJF3V2IvcY16r0wlo2A84zA4wdNKh7xtdMh29MtL
ElSLrWfOcoW0iU1SUM3Fkc7Zt6gf4hscSDK0IsIffRATslw7veCiNfOGreg/E8PN
BR4/94jKLn3sSISE/VRccxuJqc5MKKW9nyxCSnERhVdP2MAKGCV0Id2XZtkbK0XL
37VtawiFkHRn70hm5F4L96Zf434tDYZSjc5lysFfrEUIddZ6eu4QYSuL9Fdeiihl
a9FYDQcuDNzQ0Mss2lZc0EzsO8E1uivCysgH9N+962sTWgCyR4wNGSvw8NFzlz5L
1iVCSBoMyBo4MPliz/cQqR3Pkw0tP58TbzNQ5Nna7dAvTzYfiW3JjssOCI30fvhv
InwHchzdfX7WE51ZdKG3Y8yEYH0Yea8VuJGg+0zecieeJBfFkuK2gB/9xiKQIpqI
YFuJU5qMyZUFZhX/cMy2Lp0VM1D+owsOINDEQvmIt4fSJeJb/6j6FpLJeYzx3/62
sf/9QT6W6qoQSSMf02M0OQJc3c0exRLpGpyaUL/n9BlbGioqobkr8E8HWRI9FhpO
EgSfqKWPHcu3W9gPaegxyc99FJVfwXde2ByS8mrJOGjaPFdVWIic10WWidzB50VO
UofPrS+LUGuKQ9dCqT3E91hS+JWe+2kSvxrv8LvN+6btlewUJ64W8UjzoFCDGaoz
GOi4aCLd5r8Qq03yvX4vxv13J56BE5GRv2mlDhdvSOmbYu915UIgZcbSNliwGJrk
t9+FxEO/+iu42KnTYmVbFBxyLQ/44nLm7NIBqdvzM4es1Ntr30JNnQIIr6B6+bmU
UvDeVRiDDk9ncAybw2KStkJhNCadsemhZF86HFR2LGESlQ6gjzeFv+RukmJWdISv
3bmeKcrvVsSfS8zLFteyGeMy273C65X0Ik5y4jTn9plME51jf5OoKtyp6EnD/wmG
bLj4mt1x8YI4VbeMcs8s82zZxTcrmHeJ6HlQdGYw4+h/TLnpFhe3TiB9CZIg7RgB
xiC29VxToxzvGMGhuJktS1xgv34d8h1sJ9bJaNzZKmzZD9PZqPOmcxHxeZxSpL9S
mRAjg44eTwAG8qFDNkogQKAmiekTjqY6cwlXLjMIFYAIZRUgEa1ISy3kU+wOq5bm
rATu8h+grWnzqJ5jSMDTZnSeAlxHNs2RUSQUb7BYZ6wufeW+UVsdge8Bi9kLxwPP
I3ibg/3lD3JSqrmi7yFUiWxL//lQYf0z2ZOhdCmjM7HSavxFHoCUrSYGAWDR+XJO
CE3wHCMIi78ARZ5OSWow1q6EZ7Ygo5jO8RdKOafnGyvEdSFG6iADqlPMkye/tBN1
zl/UrNDRcxuFZML+PbTpJGs3CaF+Jz+34QHACzBs+Eo/2I5SnWrUbYH4o3rwXIcb
MwJbRkADtlJBbwXyPDLbGKQDMz+4WBoijotUl9sqsfN4fmwL4RwVwxyGLZf6y8vP
kRzkUml6KTu5H7Iusv40dFb9fxorrFgw8m+Mn05uNOP7jEtLLMFueNssZs6X4Cmm
LyECK9k4i5uuUYnmyg2s+se2zZxWwvY1NwliMA6qKq4XgNQ4M/YqI7Irli5ChSC8
lBdFJHeu+R6eyiRELWVmfM/R6rqGC18ZModOTmgfzbbIahKHMKv/pnzBuCOvjsTG
CrTJ1xP2lTvTJJJ+GC716eZcj3KFGqxsR/ZDfVOr4P1XFCi+E+4ls/v+jgWjEpnD
5ZNO5GQPalHJuTeIhu/BCvDBR6tFB4SxK2xrWV7Mj5fLvH9/5MsJdfecpjMOTqpn
d+TXGncN7o4KlmHxW8QKc3GHgGPRILYugPdVrWNCBYZUlwA5Hz4yzfsHtNirgFxL
C51+FBtkaf0aSAWz/E5Y7CFF+KuhQ4i492j6BKeUQKA7IaH7PaJsrPmZ1d9wJtSo
r+WDwJy7EJQezx4c95LnznFW/YY75v52s5IM/Ny79vYMZoexaCOKb1F669ozmdd6
cdhuwWiIzJcZ+9h4t3i7dqBIgQgJPl9obz3FSWLQwLxPuaLlXaWDs0xsFmpBY5+M
cHiLsMvVAr8LCVQijxHevCb4JwO4OIncs+2i+RzxqIFrhO4V5nha/Yvc0aHIYBRE
Ax3T/ddlfZq76X5RsjdUOgfW/BgI80wCzNYVIRT2eaHzv70k7WwbthhLqdIGz6Gp
DYOgNcM3ZmYIlBvaaxwAPxI8RjJMgT5AhhUBcmKtZEwfePYSRe2rnhg8YUECjJXs
GmVC953hN2Y/o1sE4UVw04PrxgDgd+r4gdeH5yOiq5MQJ52tVQ2dutRyPsnS5azq
+LYb1R/FbYEASpyIiD2NfB4KMuvH+x0wc0ch0qNUP6WOSj2Xo5oX7Nix2YjHdjwt
mROkPY8MEddgv8jFgNKMs3l5cBPf6cmSFlRC5KF5jZmWT7dnGDArleFF/eqCnp/y
LqhjifjuHGNJO3Q2ZD5FTNgRJPW7sQbnm3WykgHwVUp+BPeae1gaZxNi737QANNi
mnjYocLvoSHI0d9xS3B6nb0vol5Njo9ySsg9ni0bZPUnruSRgv9S2N8JH9tCADmD
gP5T/FwtyaaY4rC+69AcF5c44TbJdiy0RNjgdZDYLFnuSMiNCDcWL10c8k3Sff+E
FFR+qd6MNRhn22APktVdh9eeB0t5vapTCQGOa1+YFXLpvhWG6+JqauJOg+h5VhSL
EVWbmOISwSJmPLtZLnEeMsJ55hr4B4hHN+frN7GKPQnU9UuoKl8yuNaqustspywB
LVPb2PPPAoHvhsvF2NcOoEmv2DnanvbOX/KR805BPrbSVoxlLcTY1O8NM2Hf2lf3
keAuxxtyG8fkwVHL0V5sFTLqYz77zLEenWHNW5s4+7gpcc00q/kKpcVUR/U1y4yy
//rfRwPlP5KxfkRX/6bCTXbtOrEM9Wo/ay3SGAAyuUwmnBlNGuzsZ8i/5jEUREFn
bWaXpeGSgiexnOuBc4+6WN7VTBEV4jEcHC5gUkixUsryHdXMnlDA3lhIkCgn13Uq
kRYwPkB40MdpreDjPr7GQpdnVijpLbzWE2+N7KlaJmCG1QqoS+4ZwfuL/tb3xOSz
uMYP6/AWJmgHQBKzmJ8idkpAMxMbbrtSRklpOr4eRCFxp0Ugkz70yQYGPewQ4Mdg
49khbSSEiWriIb+25/ilBHxo7oxZ7DeKgUVLT4293mpv9rX6So11im7XaxDaSKQ3
7NAQ/RWPDiShb53ePjX2k3tVqvOZuuL4IMou/EZCTINy/+crD5CTnpJFcjFmXbOV
fTTFtHscmuEwD4hYOT42dSE1ztc5Ki44Uua5qgfw43ymw2FFmoWpBjc/eqxXbkCm
tN1MoscoryuIQUfs/G2K/7dQL24HjfHik7TPo0mvKYbuI/43s2quQqhmyQjaKh9G
Dz3UbvxQ8CYG50AhJ1hrdnXJnI7jihT14dB8MsfPiaijukflk/EcN76UaZXBvyQm
H3I5GaOfqaFzYp4bliYuu3ffVnZ23EoUeS+G5n9vXIQCGxySgx0Gp82JSVakgWK5
O3/HG94RW86VdRnyp4CNmE7vxs1E4UhveykZ4R423TlBSAZuOLRh9d+qLWyTLdKX
8rnLG51zlgdRg2Tl6ecYs+M1Ew/MAjgk6sNoerK7zepv6MV7J62v14zgumNCzR3S
NI5ANETFTv3P7+7vNWzMhuqMLoDaugS6hLfi6v1z6z2LpFZ4B1sXQTo7EpeW8vA2
SWYIoubHLKw1FFPqOUVF6ryeSewjdmBUTodIoIxpxqEtiyRqUHuIdbDVNLFmRXgZ
z4O2YaKudTBTHNx5J7BPHRXzDFy75LvTFnei4gu61tZ4uzxiBqGHD/onY8btjTGt
6DUrWw6/wDZtABB8MdA7lDlQz7ZGloTfIS424SHn6pP+Ysv6xi8Cc6zjgMlNUrPH
vizQIgw0QD6XkqLHIlUiX5t32RH/rS5johYRGEo6HBkDrAYEKSEQKdN5yqLdoOjw
mSdOrT23rygsZsw4KfAoR/1M7jnTDk4oAQee3a4AleNsMetAsWFj45i7M3CfGvKz
ZzLrYnuTxjOB8HmtYzQ0F/Z5/c9BVxz49E1eh1fr8RK/JO828I4w2xuaF7zRXriF
wNa/4+vvLowwhYcDsyk1eQi6aCpS/+QB9HFbDvfDJkWuPg6YT1PZgGbb6xFUrqz+
FflJ7Lj67uiCRIPsLbhXO+bH2ltRWOW2/jm4t4ewzXkVBdqok3G/hZSZb0e4t09V
7g9X5x4QZ7CaPFgj7jesjt4jCmK1TTcm1vp96KutDz8EdtXiAlRdJOeNPRrVDvZz
RnkhMJyO2ry1baeHfwOSL0GheO028bV72e/GiDR2G5bBZ2I3dx+aummQqyYfacPK
SUwLGyFpVH4QfciyFa+ES9h6m1x+x3H12ejCfB+GBOy5VBkpUtz572APUave5mbu
yxiDRFnVn5yowFmRvg2rOG8pLK2plhzxyebR9/Dk0Q0hE+xg+2LfFADTbEowpcpI
QwIrDx3oRBMchERB9/NBmmNSZn6QB/N3SbMwsIIpA+K/8jemXLqAViPKjDeFi+xW
UpTqzAKMabiNSrMxsay2+dvaQ62B3iJvvwl/IWC6FWAe/ixOt41llYF0Esrnx+mU
oKlITcgQLRYBYldAZXlXYWhAoNA01eBDJhJEtHwcrFzTVK9ptOiB8atiJhuh+u7K
QwX4JU44SSlkA9LruHNwLBmIWX9NZwkAJEkL9bWFnOmMqfL6NUDE90GS3NBXvOW5
XVYnGh9QoFuAwlYGMpdT5u7ULF+58T8AZULU1K4vmgBpVpaNCTCrRTgC7p18MpLx
XA89zDkAQ3i6HMuXDX4ZqWS5phzXu1avPzrgNt4JDzsWKmIlyMNeHVSjU9i9BPez
z8AsrDYFCm06wnT1gBobdaDOoeEd0Dl/iBtMOxOJaViJWbzaR3EAiEsJtQBA8BR3
sLMAWtRazyAEv5iDF+BmN0fSKsScJ9uk4P1FrKr3vxHgaGaw8fT8HIjmLnJTDjom
J1KMk5dNIyMr6GMibeU+s0wXLlKuaal3ZeBXqfbJR5dJ1WsN6Qy4KATswnU8k9pO
YmuazVEo/5KeEe9Qh2xNGX3+G88e84kalP3x8wBQQixjqCJbVQhwtJ7tsmbxybW4
BA5gYDJ0jUQVPG8XtVEk0fJf4nlFJMELMBTjzVgfA9TQvgkikCdVPrlSeRV1N386
cmclYa1TtpA4M5LbAVEqx+Z7H9NbRcJsh0QaTxBSJKE3Y8d8PMMNUVZug736ucVx
HwKM64b4pgQFgUW5kXPTAX70JPr4c7NwFN7RF6HLRUwxMBWZXNuG2MNIwXojFd55
D6geQXIeiss9DbOyrSAknvxKDTIpRWhnKTxPd9Jmr4WOgnHIrbPveSbBTx/nfGkR
4AB2Mem0TVbV+kpTpPm8i6xaaknvz9PYIom/xMvvyeiZyC2xT8wA81Kavivkrpvl
W6+8DLVtkp92Rk6CxDQB26dFa/PzRRbQ6jzt69eDlHptIPF0ngvFX5l9hjZkm7h2
qAZ9r/YkK9oGmGtoND6SpGvARa8dLG6ReJppmSLHEJtBkCS57hy6nL+AqzvYcGXw
FOlLDPeTwszWyD4mSFUmPhTkF7OyKO5YCNj+kjL3u8fj9diMy46CwvWUp+5PAW9G
etKGtAilQ7CgWYRzAsMi3RMDC8vmuI0FKckd1UlkJPE0Fdn+5lgJlpDgcZ8H4NJU
Suz5H41aZ3KK79mVJ/cu8bUYFV5H8OzI9jeH7+vuOdThEopJ3wAM7JTejTzVVWma
fMXvnNZvR8VVoFFgEfhePbg3jWrWeizBDpvtKOY9zYHSTaL59LaQdb1w+pUDvI4A
yCaqQB+MPwQX/xQk/3SdB0Ko+PaHCfXW3Bt+uKou2X2VHLKzedPb/N+0MKO91WNM
wz6AfjovpzQ3virajtYNpmfC3Xu3QxuPTs6GCnr/pp03URWdWN7wqdXE1YBzfp73
3DzdkghT5Cj6wj042wideVtqiOtJn4aQ9bYcHG+6iZ4zK2oeN77JFIihDOyFjer3
/kT/QK5VsbsZ56q7nw96Cbz5U6vdhKznWYXUR7PdPEFrBjFvEKIMxQExwCGUXCb0
oGh8ezGcYJkh54WwtMXO7pLYs2gob8X1FIzddpx9GMDBIffWmjjGgSo4xgxEOt5p
THfB9kc8kIGq2DMr6/DA+UfOIn8pPKXxBbwFk6OV3wLtCZj72/JxQWS9ZeBZaOJ3
4vwvk1n710lRxl4P++FJepqXFaekVnxKYux2HaDx08Cg7ViuV+emzsVQe+2m/6FM
I8JkzLVOpU4d9MTr7+vTX70bZ5tAx0VkgF+ZgjxWzv7ws0uB9iSMBoQTeU4zFK6G
MxQCUPFPo8bY/JIsrHSrPGbiu3+or5yapCkNxHDl+1AlEX1L+kuMuDEhSM7Vhork
6uO/r//pdWZXdlvZRYUrBEfWutxpXg18OSkbtYkMziFPxaMSoxq9aFF1z3WW+PGJ
ssMeVwBA4ewRO8g2Mxk4K9EpXGsvM58rMsii/I7D+bNb98rA7exPfNvpzDucGsMC
oC1ZukkKBI0vSp373GBlhVPpENGuH4eAyeKH148ucM+11Jg2pqusRVCvBh+6nkIm
980xswHMBZMxiICWo7tzcJTGixV5WFt0GJZNAd1hfzO36oV1773KViZywankXVZ/
7PqVFiB5WPuS/HXaLhfiV+kPoIkm5xhprGsw+Qlh44SVHXSCkTTz/Z6ICWaR5Usd
F4YPXtate3gCUggEjNSeBxt9bwz15LjcK5BXIdm+LkBGdRieQiI1/27ezx4HZNwn
rjiODb8sjz8hvbgfKQXCrUbROhpjcGjtnW5vQRWn2hgRKHMR3x/YNOXA67k/Hmy4
LCmsn3IwNSRgsYjeN3iyYs6BY1i9h6uTVgOFJfDG521NUHgkKswrMbUJ/RvfziXU
QUHVIkG7ffsRYMIxZqdu/sx7JC/Yx/7ELsuRTv3b9UtdgbDk09VLzmxy3DvjTuTZ
bGTFNPT7uhh+H0JaqfZ3Jd38MDL/w3STMjakgkFrSl5OWNjZ7/XL9/U/EkWBSJqC
5NufgYhKX4NZDK2/iLiblY6Oe/R78KvxTPFYyTRzPrdV88BB6zTTkihD33H7ejYs
+POZlWaidIHOspbGLC5dAS7CDm30m/lJHRgoqgzLCirdTTn5X75CTHvcQjJygapW
mhoeQMKcS1Iv2GrmaQ2xbzGUWZW02G3SdgcjJgGNZOvu35IIg7tWvAaBS1hS1yOT
h21n1EsDt96m6ifHwgA8ZhFEfS/Hvm9P413glq5n2cEPEa4ABJRGXmxAl2VdQauz
7ffrmtta8DFR+/WQxQEYui0oEcaUlYIoBCQvkwMgGA2lns1mqS5k923fGv0CNZgd
amb0HRt0fT7V25qVSJYT5MjqOt0pBM+KUGj+BCDBZyPzPeWF+WS+UvZJq1V9A/1l
CoZ3vLOQaAUYofn7ubLanKs9G4qmsVYCDbTIrG2+JiPYJIu0iaD19Cfm1kyRMCoj
og05uzLTR5KEVsyiaR3ECpcB1ePGOUVd70pjn5PTlXFOdzcbHI5D7zsA/Vef1JIc
ZSgNu2fXctoGkbbHMoCpVlhzO1Nfy1hxMwNvXhctsxJvBBvtHlSSWtOKnN7d33gK
fIAwGRmWXyD5FVhB27eBhBmnbkYK4mqKc/kDRQvSAcHZE4s2ZFVm8P4pb7WChv3s
YtiB6fN13uyvgGaMCvRjNGsbDFoTzeXxabCJOhLhPgMPR96B6Sumjxvr3AL//h8y
Vnpf1Bduv0adVAXRtwqw85z3TLiUr+OPtZBTPQPquLKNkVRL41yh5wELXpkCYu2W
HZRS4o4G/yQ1b40yEGnb86oQFXya4DOfbkS/40aEnSxiLnaNb7+f4BnBdF7X3DCM
PD8p+ISB6KGnNCcavnJyUD6gRp/ff57FVmRqJsB6wa1yvDOr0QB2RIGUQXGShidH
t9k6GB9/usaJpiv85pdSTpf2WA7aJdYgToHziELAIRTF7M3/gHNMdAjsR9Uzrpgt
Yk5G6SeeFhxTK3CW2LOPEBTqxajqu5TgZ9ctw8/pGevZZ6miAgZgTo5dRxq56OkR
EdKLRZBUkVv2ketWjuawDFuoY3NXRklgldODzGeie3pp1oiu2H4xdK9430gF+75+
96lpFEuBCyt32jeEuDUQf/6kuGKfmga4mvwPDA6SH2ZVZSUXX0nNF8vxTgK20FPT
/ygipAAO7uwMdBmvF/JP9r3Sd5AL8qQuE3mFly827+xS8U0m4+F5Rkf0OxfRbtJI
Tq0N+oMKa+/DoBN4QPqe76gD52oPFbasModwX0MTnF6CyEiuFF656xj0u7SUOXVu
FB+XLVOUq/bO3cb1G/+6bRG6RrsDV2LLjlp9Hvm3P57ktUflpaFsOuVuqbyuCx7O
Rpo8Jjen7p2zSrU58fy+wytUiDT4FraCSuwFZdraU6A4q8JxxU62aPagHw2cPguJ
Q6HLGg6Tlfpg9g108rzuKy22NeISiRP4PJOIbOSBolDI2ePYGEYXUbeXBCJOhoow
7S9k5hKnDzt6Sfj6eLa9DiLk7WUKhSrxrbbAmKJQxwaQfBTHFMQK/KlVZh837YVs
4J4MiGw8VIJjS4wG0qbLB7dXUnbezyW1eqOWj6cbKbMOaHzWT1a0+1tZ14zvnF/1
qkZFjyJ/O/4nuBSuM7kuYKC9VeelqQhCSisDt48AZba/O7r1PoKl7CAvzdDkNKBa
jb9t3xqLs370KRSUNaBLaiQGY90sGxJZvcmmEfgDegKHx+DbwqqWcWCSKBx6yjOa
ZDPIL8c3hH32rQLroJahsgU+zHojGEXZuNI4KIwANW8EQYGQHZ+lJAmzq5hIQ0t6
D7ZsiFuK4zpPV0NzUHnqi6yAYogsHN3YFAcAgTSN54gfcWQCBGUhTLQOT9iOB/ma
OX8wtvgfz0TExXQsS43sxDwM8/NVPoOtF012TKN1WhEcQ0A2eHQUi9GvdM95nhqX
mUIvIs4NesFSTH5uUK3pBbyV8vxM4PEtNO64gbPpaqQRxGR0tlAzThydA8BKnQJm
W/A2oD9nZ+XDON3lE6SN3zOoDRw7lCFq21DrOEB/4/lYH4WmdAmEjNIJW72SD+UH
AUvFAt+PZwOBLliwDphNZa1Zv2bt5hlejoJ1SOCE6jf7gasvQygdMViEQHYAQ7ex
5Dnbu2E2hjbo+MJslNf4eJwMWC+lK3QpxXQs0HFErNP1MzZ2N/9jrtkG+m+IDrMc
fbdXjJZ9mcJsh+j+LLXnaAAxj38cs+4GJN2bBA7CqlD5BpVimgPjKz+31aUKSkgY
/J7FglSryyFdE1/j8k9g9Bg6vH1phsF4ldQzdQZlSnS5zSji1YDl1KXNqfVV/WRj
vTzc0vIo08iGfUQtriUzol4gXQnQvdbD65ZXs7nyil3aNIe/+5aRhirxRVm8je7d
nZsmbzWtAXHmORNzzNOy9tV6ZDLcqej5TdOMEGH/Fb+JnPIdv0quo5kKD+6bzYSf
fMOM77egYIDXCO7yUKC6T/9qr6jdJVjnSakWyQwRjvrNGGbe5LMRMln92TE0kOBN
UwOwoy0gmvQcP4eKzrB2rg4xdQjRbJB4MfGxJvUarDqSWeVO0/ArqIM0MvFpmHsE
149jTdqXjEizyzR1oNbuBmGPgYszDJ5gnXs+WdW8pzKbiCSKnvc1bUichaV7U/K7
6XOihCXkbxWwYiM19plu5qAxJJYAnoMFIcBhs3C+F1ZI3KuG7HIESpogzkRNAOQ3
wzXG8Uou+vVCUbZbYDeiIgb4+O6J/LK0pqtnW5p1a9fuvZiIhzfVUDcsgYsdv1Fb
BXy1WxjUzVJbubM8mKndMqdKgsfCW1qdO1+5lz2VYp88uVpUVlauQRa4bpXoUOtL
aFJzb1W93NV6DAsTsDFr005degc7svYfJAJOHLuHkr6PvY7LfRGR6BJHR5at+4ef
YdjnLqLGe8HvMsJS28Ph54CShCN8SxjbxFmsttvBig+Ze84grSNl77KKkmVQsE1Z
H7MqCxNgwb1ORIqwoNG7HfgIWwadFpozDFHFFdKiUlJQYEgg8cDQoTzdqAkqBdEB
dU0vToL+pQV6TWgYwkBH3H2y/ZovaPh9eaaPjkU5xUuV2Qd7qq747N5qxmQoDVhi
Q2jB2heWN2OrEvQDgNPOQp65T2VQFy2r2kKJUjDqBiUyxcfDinkUZ+FOptmcpHMe
5HktikNYZhn23rMYSFiYfT/KSc+RV4q6CVHkA2CAOCvAtJcr+ovmziw32OXxUDKQ
gChGWV8kRcUZ2AmL/V8rOSnCgnW4ZlWt4fRRJirojpH4EYc3jkByxoT8tLyV05hl
wc3ximxQSEGLBY8lGZSAL4kCW2AnqSGrcP9sXJ4z0N2VrIuo2usNVx3BXoq5IL+k
QHLttmpHO82JDwOld/ojc/cGDNcsuDeIMHqjFgEX+C+l7wY6mU6SokzfmcvlJsV+
sN1lQaqKcK/rZsujbE4doM6pSGXWleQfZ/jACRBXPGgyzJXCaMKbk2ajwToleozc
D1B3SD4hgF6w0bMh9IObBljx8u3boTrLEqJ1UctCUlpWggwEAepD2tMpsM9dPlwX
Opi3WzR6XasTvt7mfvCH4a8ouZE6/8SoMYjS4g7Xp/bJlg6m/Gt279es365kyCwD
8TnfJLovsaBKJwOihwUeGKiZ/Jlx2vxipYNXBH/mSXjjz3+OkXBelL/MqiJLZQPR
weqxRb83iwVeXOfX8o41TgDYXWOYYysSPGQZRaMF4MLr1Y0okXZJALwpM5e77gAA
J0weahijYh01roWtHEt+lf5+ty9Yvb5F1ddEIbm0hcXtg3/CzHD1lkntN3kz1zgr
oqEAXuJM2/vw1KdsiBZRnRWJH4/DMJxeiVaogYBo+cmueRM6l04WTXS8QcbTil6u
lvQ5/3W19zTYJS37w6zdh5UA/ta8Sj2q6IcEjN5MNbCPnrE8NCRCFklhuZtLOHip
yLE00CYvZCyMupUImmO3/3pdhzBGXDoEkIV6FlTbNmu9XUVlcx970DiR6HH1s02T
bfLrobudIQB/A59ejOdh1yO9HfHZLBp5N8+M7DAjxYN52/T1xk0+HvGLDwcPvp1R
TASKl59vmbp9aCYn2x2WuOa4mEqxyUJDZdggvBYUtrVojyLVd0qGleWWZqXxbJUX
7mhLPfQUHF9JecD6uuXZFEs5LU0zirijbUECwT8E9dB395wmVdDltQe6oifjiGUu
CtswhHnVcnTnj58KFXgR/Yd4hxmaT6uaH7sbhNcGCOdPDL4zs3ncmFnMeTlv66NZ
vVRCX2Mgi7mNUucsV1+QGk8UUkQLiBfMmAmoKQlwXAG/KDuqE8KS+qLzUbBtaJtT
FzaiKyNKzxeCp3f5DcUxsukhrJ4IeS9cSb3CqCmWTARTvkAm5MX94oCDj4/AeFdy
7R5Z3+o9nMIsJpiDak3rMy/OniPICxuMoOmLLrLI30dMSvG5yFxDbfjihvwaQLZe
f5Zfv7fEu4Jvno8+N1h1tYxdU3lGrYsdf4jB5lhWA8pofgSapFGXSu3/Jn2/VVW3
iz3UA0Gyy3E7zCAyO3gKDpo1bPY/93r5akMReM2nyZzco103QapHCqnsa/Vl3Qqk
TThu/g/1s/1FiKaQJe4Nmrjg7vg7zTebMx9kW11Y1xPf59Np1dHviKUAbkJ7nIU5
b1IfUiGsGtqyLMzXhIn7TyLw8EqeQ0h8lYvGfd5bBh4SpLiNH1x81ndzWC9uLT15
c9SApeZJO4iArecbD0TSg/OtvJ8b+T7+umMAJiLOLvMzMj/O44Mt06XWpynvmkUq
zmZo8OoeyD9j4RQGOnqFgH7JRVEYQgKj8ZG4VGTgfNT0U+3Qjqaet4M8KWp1Q/69
Rb7ETf2ri5fjbg0yPDh3fibDY9KlTXQp1FWgtCDmcL9IuZUffZPC2L40VlEBBoO0
LVJMEMltsKlXLkWtTN1Ivfd8yyE3abwhfEjUAtAEvQ14A7Vnko1HyMwIR5CRCSgb
UyM9cwaKknMTD1P9KkEASY4Vr1WG0oYfrBLLYI8YEVxYF4TS7iIB36X3/y7jO9mY
9bH4LJboF/yJ3WTBgQYkrfY5trlu8/1aJharK8DXR5bJGXu7RuiauyFyYeMmixkX
pu23LxAGvze82IT1usnFpQnRekHt5teiJw1Bljg4osSBppYLxTf83L/Hwz4YtjZK
stGAm5AXsXtdlpoXDX7zgVRPo6ebgzf+7kqjnL0suD9rhE0EWRp+7r8pBRh6SPTS
Yl+39TAtAf8jwW5Vp5s5YNB6wEO2v7HDl9xbWbTsqnZDGVXrWq6TYOlDfEiKB9uz
ob7jjbPicKnQ/duulsYpiFVjUKUu5zZqLbjVdn7Gz+/vGwfaTtyoChkPm3tIXpln
OsblI0EFuNSr4yWQylxBGoQtOIGmu27kDXnTGIVpXDnSKtAtNXUJ2blcDjMrBVed
FnpOEyHFpzX52NTS116hIukTHw6X5parwYjxzHwt5TupCz6eobeczHRhH7qKeBAV
rX8qn28P9FVPOXI/eTBl12pNWAcNnv/HXKCKzGoQ7LmO4Sk14SpuskqtwlgX0zPl
LsgMDklMa9dSkxfTZvP2wicIOEOQqEwrgFjGhuRPGiL9jDPIhGijnV9Fg+dl4GNG
QjEeGVS+e90zj/kvqApwiuZ6ni+VSyz2ZTxUUxj46Bm1B9+FmmMAfFK3K/CUUB6Y
RYClil1loW+Q2TuWw6Wm7g8YGEtlVDNg9DFme+DWSFqqHI1dfBzn9lKQe29raeL8
rH2luxKgsIqaxh3mqSevq+m9jeXriqe/PEsGx0o7WSrC3xjbX5cI36dlFPGg/iYR
vWktnDVaCkGCj9CtEMV68yk89o10WF1d2hupE3V4/UHZ+wrgk7qdcqk4t2jEQ0u+
+TA18gr40xaiGNFA9oGI7PKp9pnXYNCbeYwDW/4zDMf66ErMUjWlXJw61UzMs3Qq
FlFUdiP9TxtK0VgbPtru8wTzGMgfDpYAU0z8IISOBHpf1J53lrvfd8+6EbooXDdY
re6eOQ3GTaEyHDjkGBFd1j21kSjKezPgkTbTrJyDCOe101frWzLddL9DkMAGJ2BJ
0EP+jDJoXwj1alYVws47EGq2YwyI0wuLXqmBcSSa9/rceLYw3FowPhonp/vyyJSK
spXEppQq+pjuQ7JnQzx6FU+xONf1aebjWUHGrdXLbud98/RNgIGqcAVeCrySOxTq
9gdb04oPvTJvFl15/V9JycWNwOAVGJlSdQynQCXqBXZws+t+xIfQxI0T9I0WDFdV
3ad012vLMkhaAkkw9dsKXnXeYsh8XO/U8d1bboxQwbMvwdlIdKtWm7MRoT3Y9pkJ
K9I+xj/QABWW5NPe5Go5xD8l3amD3F9dY+JU4SRB4TvifHDw1qR7f48EDbhYhAys
6+jPBNEEtxVWaJLosk+OnTjpjCh/4hmPXqGDkLVfokjxU4gRMmoPY802cjtH5+j4
7hgeQWEF+WaSwpfLc6V/5mPU0J+SQzRT6OXtXf1WPomSrioyJb+1xuHTjJoNnxh+
VKL1XZuB7pDEs8a78jX2QRxuC+0ByeUSNoYkY0yQaDDAuRTo9FKfzPxuhi1GYeZ7
zxOwzTI7/13/4+TCwH4HUtfjDlXbs46hTRIY9GPkSKMvuBirAmN6idC0to0jxQKU
MjUC7yXE6SK2mdcfHTYfcPtIwHvrA7auG4ASXpoZxrAUSc+En7QOMc9goSxdA+S5
uoHsRNWJHcA1ETMa/H5lWkOLjilYI21IkjEDz+ae1oHoUT/eUqykQB6VJyVWoBLM
lAXdGu3CPfY9rrRtyW1wiRT+Ybn0zN/8mUmg3/EKOvgsyLkzrS/Rse3tNxr6CGhx
mdwneX6mybG+qs/l83wyRBCy1dpzfWRVK0MdBcl1UwJtdqfC33DWJfhV668f1jwp
qoWkw0qbvU9QAeFHzYb3SzyHJZP1uwHxIUWmY3J/N8O/0g5GERMnELvCJLMdIVz3
UR/4XkxDSG4cttsDPwJp3ihYMVTnpIN6ZGw/jmTsiyeVbDfqZZN5/tMq6YdqK/fl
ioEPDGQd6rJ3ZJMHDaj0qwEMh3H7QZ8wGwS4lHlkKIM3hU5aQoE4d0138Tze6IC3
5KX7MaoYgEu7FbvAezX74EwI0yazfcbhgOAoLsLTthty0FW5X/+u9TGqpfs6QyiL
0trN/oj0Z9OXqKItiARotPLNBy8pVCmSexB4zczTQdWSE+lOz54ZaWIRIlyoeGqH
NOLZpkVAs33tnlJGvR9wEuOTvyYGsTdbxFRMJCPzvLvlzhMNCCjq6bi74O142uqV
i14aFZyYWnpas8zLjOiAKSicn5Cf97OsvfHuNWcglRqU8Xo4eT0TZb92ZGwRIxtz
9Sh/ChKpKfgViWFN0yan7nKZ4OpBJlE91Ik3Wq4rkGG9g9Sd3SWkVBLF0tqy8n8I
PfLko7jQZj5VtEMFJ/nJPTr9rXlmRkYZJEgXqrUoOp2zqjLO2BWb31kAZSBFw16W
scjbbBe25a0kM6UdgWk8I5DkJH3cfjK/noll+DzA3XC2GCqWd2/pMYdoK8SIIBtY
P8yamlv6VxLHiI/zVhQWITHqmqbbwLVNsY+kuJ/3qCD1tmItsLdNoYs3ehHMYYmk
4d+Q6/psgDslLnPnRwdn+9U1WvU9YoHmUm+imRhGG0qiTpEVm/bVvj6IG6c9f0iQ
fxtpS407U1J5EjeDA3h08Q5IDW3mK/7pa8IXtLfU5eAqnKVr0jidX5LH2ToTNwiQ
bbbUUTekPqnmWXZhgbphe3QvcUJpBhHfOcDRm5UGEmgz5scwOQdKGdltRA8g49Zh
SnhI4K7gdWv6Ot+6GjepKwz049PESSioxNXAutJpvOUHMbaNVJCcvIrwuQqcBl2Z
kkMCT2UyeU4zohN9UKU4Gw+pdh76zYKyQTeWMMcmd0wBav3RGWfrCUyhi9g2henC
YDPGwO4SagFRrmGN4buGttW3sjw/5NTZlZCS64c2kfLYrjVE56I5bXxCi1vhhdIl
GBehOhAFXVqBJM9gZrunFbUkkgxPs/2LrtJXr5t/WCejhoe2Uh7vGvrAOKLN7z2o
vGeC9GN4zz9RfUtyH5CsqIPWaPFF9CjNXfW3E0M48V8FXNi2in/dHjXx7tmCssgW
sarzvCOwi8mJ9jKXVAmy64AJUYXB1nN4pNyCB8tcwRDul7aLDzpCdqV5oGwmOyIC
TenVzbLKwC5nYs2G7DrTvx66tvpspNgU3IiTeXoXT7SCRdb9Duqc/xiP2tW17ilM
b7f3Eb2pNsnDw66gBEHWnLIwgV3BOhRxmKGkzmzgEQDp7ATDhWv4c7AU2XFmIeqj
TR8ON2w5Z/vqbH5hQS9GI+DluhTdcnDSKv8Kz0wiDhXoqnn7ZeeszYCuBZjebg67
nnKXZT7or7pU7/6qm3zBb2wegT11LKrbNojZJu2S4fIPFqFrKp/Q0ukqK/w9NxZR
RDWi+jg22NnHm2KNR19JRiDZUNAW0oXl7H81MK13q2ZrvApoGan200xElKK5IVHA
ta7OV7l7GQVq+3G6qarQKgiKPfhDHcaJSIJMgHjo9MCFb6+7dc6ZoMfT5lA/AdCm
X+Ydhf5XOa8spS8NX+NJ1QU4K3Kdd0NwI5ROpYGZ1pLrtOfjk7h3c/JNzoNj8tyZ
/Efh2nkIJoz+h/KxzARbs4pzXP2EB0ucDbahl1tK/WE6ioOsPZNUhHiJe1y0Gs/u
gEij6ZO0dMV5+PFahq5sxMy/6y6yTXg46KRAbIaUMdYDaZBs/OoyE3mqY9krDHNR
lmxher9WjB7jpvf2HwaKWXKOuVSzV0GHgKYpZPcJjKIAtuMKjSNkFs9+kIDP7eIE
HQWbE1JftAPAiNgoRcWyrMukrdDL+LFPtXOrbmQi0hbYusA8XvAYTYf6jPUYQG/6
v69bm4koGRfpRQXJPEP6v7nJXshiXnm6H8F00U0gpwXK88rCLD/nSQMlvLxnCbIz
oD4VR9wJJlOcG4MXQ/v2i2+sXzDTkOcqrukJgxfnMdNra2H9tzL28JAQltWGQ9mN
mWQfHQBN2UXQ9E6tZuw5TC06/WmNLVaPJCtT3KbHM0Z4Gdo96QLAakKRpcjKxWHc
DB08eU64Iv0Bw3tG6JmEDNc3OpfiPFWYXUoy3gwNTHaJWfrFKy93UP52CUkQGkp3
EbcrUtMBH8PFAj59MdXXaDPvpDyn1wDccCJrscozy4Yk4yAAbJcHi549mN/dR/aB
Al5lPaGGoriHNVxRnb3o4n4apynaLdUMGPre5ya2puUupuP1jv7B2HKJ739qWLWJ
pydwuDTqWgwFSURWAwE7i/CpYb0GL27Z+qo8+kD9621adNNujQUrfZbE3fnau9jc
1fjv9suyFnhShYACLpgx+DADGAr3p6Ifr4Ooo8XzvlY20aEvIkjMTEFTvBdjAZFs
mKhr4qYzJejFehzgTN/Sy4YGn5RFcZxqtYniaHIEPOM/py2jL2Rjt4unDSY5kol6
hHIlQeZNWurdfJvVSFwP+xh3eT7MoI8ln2fwAKry5YJRyosClyBWcc09HzXoKwcY
SwLvom4MPh8cRrOn3CHSw98cGYaMKDTI5PYZ5uBj/cmDr8V+R25HAVJrTKMTl1DW
MVTzLIYc8XD5cxN0zK9xB8iEcIWF2HNE2n7o2Doq07p9IC+2o8jpaIVOEd5OhvCI
QEh5gbk7lHdQfc6gE00emqTpDJ8mJcLjQIaB0w2miCbk7oJc1IBgmjSUIlQAwTaU
ymIB+pPGCJv+u+IwGZOmkWGwkrcwkvOzQLDR05r5buexCTaf9WeCDT5rSdo2b+V+
XiNMFmwJ+CPYhqApw1vDSOLqLzwvMIX3cIs8PalJ56HuPD12t2H7iW9Eo45fB+NO
8RN+0m6C/Rzw7SPwhruILurcouLfRmKkwO+sjPoIBypcLjKJElnApLp7PZUIesQ2
48ZprYeIjDH09cJNKSZI5kcoqBHNTtj88RRQY00QETIo+1ES9MpQT0Yxe4ukiZSs
1CHh9QSde91NHM+TY7G44rxK9RWs+xt7wU67LTwQqPkauXWTD1k1Cp8e50sEjnJU
8IdgIQjNNc/i0QOhWjYUMfCeRNMnyJ4kPdoN90BumGXHqsqufsLCge9vG427JiBM
icBUhnUhparGOwUxGwdKue4kUck7ZfkYwkyB52gqfDybPVrm2YfHPgR7yH4KjBaH
oRxp5X39pg3xn6zQPEO84kxlYc70c3rWRjWdCDV8toVj6Rw2+om6R3905uiBAoKs
/bNZpL34i8FFb2LuhyHX6OjV/w+XaWA0Fa/ZrjXwWEteVbhIXrtJAQQ4OTxlFvXx
FCrBL6+xVOdVXHVr1/sjKE9pCN8QbqTEf/ZS1WLdDQ8n5FcngAqIe9F4X8XkgaMT
55JaIs9Vwqqv/abeS9AahxHF7ucF7+oVEfF01CWQCvUvK101huNGl3G7VerFPvZ4
Hab0BGJVyLIi4Zs8FZT/X/L+MlRVWTVs+MtKOl6RdROJ4ach0+Hmm9NQ/d2/T/AG
d9C65Bo0t82cD10Jxzoq3cDDAtLA3bRck3JPlOXb8mt2Dc8PQQUnGrVJ2RCXgIXm
CNU5Ld4vkIkhSjCdERV7G+QLTgmWbVLgWbKbesbxe+ooCMCwIfJU2dGNLaZfb58Q
2hfvo1ynm0a46jfL7JQ5t7f01e1nU86KODG7WB3XZz2TUA0obFg1opKnK4Xrd2mR
TiC9nOqNiW6IwrCNzqP/GTchXZRvd0Qx/w+PaUm/SecweOMc04JRC8H43+c+Uld5
ZoNVHWVMOTMlNFlcfvW0LBXsxU1WS8E44VGY47uM7FeCp1BFtCloarR70pbs4CXj
vtujHe94GEYWmJ4cocdEC8jk4X3CSc6saJrvZh+ayA786Q6M0eqOY6lfNIU/aamV
zGPV1NGLcBvWoH8SNsBjGBew/BBlt4pvNmx8T7A/Qf9eNJMkEb4njuSzA7Od9Lu2
4sawwMfYvb0N/dg256cih6sD4ec/lYMGIfY7IK+A8aK9bS3WHI5atnG1tp6bqd1c
k7Ak8bel/iQT0llbdcVp1fNNNRcWRU6GkSWsGd9bwEugHNXIM3vsArdc40/2JQIu
h1ICT1MkH2gJecOlB8dgZbOHfbzFa5a6nQVQIHHAXt7/L3/5ZetHRATBHVKiGHco
FjC5QWXY3WmOd/zo6OP2AdD/8/sQArS56bSKWpqbdmIPGYVhkbjXCzE1MyqWIK0d
DwL99PXMYmd0+9ku4JtEICCn625TjqGTfj9heby62zbODO695EMRQwHUN3Spavuq
IiowmwJ3pX5TaNtZi5NJSts5qkZXpX2oFplB3k+1jVswIsF2cV7CGJWK4VR/WUlN
GAyrtx3aH9u8wN0PwPn+InhLtBzhdTV/ex85tcK92I1n0A8yPIGJBFFGOgcW5SOw
ha3rSSrp8lWuEJTkzDz35+KOmFPWd6fSy4vkyfBmiyvlLAZvj34XRYkWX8j/bpFK
WMg9Gv3fT6e2kMjyXNj9HwnMoxjLoU26X9U5mbyXv77iX35d2TcwAmtQ19a+covf
7jkvVoaN99SoS+ojrCu+lb+0cvX0N3rHXO/ROLdT6oQxVZxsheJp0wLh69AiJHeh
7QJF7eGmukEKMPT82PS3SN8v+h5oijllhFN9X2GtXPpBsEJfxyvL9/jikoyGTDg6
CJn2TQRD2+uB2NnJBvUwySm6+SqYbhrq4YEPhYq6AJm+eqAaqVweHToqHIe7Cbc6
q9QOB0FV9fJEgNrp0NbMZF2wERiNUMbqOjNPkqaOLSi7AaBrI1uEkvhqj7Zi1pgC
ObEU7SUmvs44wdhsIBbTsmmWX6Z4U75JBbk+5uJoBc1cZua1dlhkn3sx+zbOKBVL
L8QWniddRl1RYcxxBe/ya4hJB64V75CrbxCcUCHyXsetvXC4dD/0qBWVDmgapPM5
xOFB/gEzB0pCa5k0DEhO/XDoqg91H2UYgBSzoK4HWZ2WHzSbgxlGbvhwISP5T1NL
08DTyzwkERqBeKep1HgYAcQ4+8u6ikz4AfMiBCMYwpP64IVhFtQzEFIUKs+27Of/
J0zVKv1uFxDmy73GQ9C18514UVOpmZzDRRugIn8v/NTWLzYFoTaLNJTSRLUbxuTc
lmbY8tK1QmjFWYW/0bKZQfD4taj2KNLj600HrTB57egLx+CJlVUdRvs0GiAvEDgV
S7VwoTX8Q7ruK89Tx06kRlp9mCg4bwrnV5Ay9SMbl1xveocWjBbrp81kcT+vMWV5
3CtPUYYuc2alxKMlj15E34NrF4ErE70WIRdPSsDEmnJe9vYisQULWfCSK2mDKemM
N3MLcqAFSoaghgg54WyjEVi2tsbyOGDcdstOorhS44HSvKcjfDDWRyLreptBcWSr
llav4JRPSs27cHBnuEXCcdZLTmmNaiJwyAh7Hc5e0a+5ER/hw5ee5MlHWJSBlM3/
4+dVlOxZ5J3bsZMWuz6Tj8AlDFvDNAR4cp7Xu4fnhUpBSNtL6Vkm5MUeS22Ko8WX
WRVEEZYmCNc8zaIKID38enG7x+8Cj+OrwXnd31wM89L5glGR6WhMmYMe1PeUmxcx
bZXuz/DiymT9kLIbiOGgZa5+PawwRZ7uyPfHsWgWyDfGSA76/EqvSwZjtajbIqRM
jf/oeTXNnL21nXhn956Tg5IexdQsylS7k82k4qgypIFjk4q54ZIdtA/lWuUzTnz4
lhAel1SXk6bfQADEJf1WUIZT2xSwBrigDB3hXxNUpzqUBDNY1QKxT09A4ICglDsO
DLkxHt+hWs8joUvErfvURlQj0oXOKt74RA8RTyhz1KQN6BuiCCrH85r1+I0XbTlr
zf0fT49kBa730de6FsP67QsKpQVNF5CXFVsCGdeEsyNL7Qo9Xod9MzWX2KgzUduE
WXP22iLreJRBv1jV8E8ewAOD7e24ng5qdzkD8NaYtiL5rZRdU+Kf42A+laR7Hrny
IS1/DCucnWgYBxerllEDVToTOsiBOcoitixWTWAaAvI=
`pragma protect end_protected    
  
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ZXPmc5pIRQJ7Cg/LpXx5lP1NePAaYiaL0RZCl9xr6zotKp8Nd9eRrvSd3nTFO03K
M9YnIo+0Ddilb+4bCWhIHXoj4P6kOaK1L71nrfKAsP9z1lVyRjd/acZFRjbd5BSP
NsHpi7F1IuSu29ZQ2eOKKKxX/p9JdmTOPD0f/yr0qy4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 34028     )
elRo3vgLuAUEWm7bAV4hVmHpiaxgu3bsKwB2THBSE7dJY9kOm2JiJPC2z9jMd1Qu
avy+OXWEU3dY/n3WUkzQaQHzVoxt0EiWY8824ZSRH6FtZToaYHtOp6C5ra3Unjug
e1y3u6tokDPTtMVXWz4n0XLYoRUTWxOue+1soKGIecef0VxouzP8pBmvxxTheUe/
nAlFowtTJ0d36+Kak7aXWFPR+TQoqZ/y/I7t0n05FfAvVV4hh4++9ewcLVYIvSaA
`pragma protect end_protected    
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Zw5qTPB3l4KvmbQLUDdLovEKOshdtwnRA4ajCOjTmdsJw6RVoo+4aoCmdaAZQy0N
HVRK8N4gbufGYsU6l5icN2HD0O+YewSnReMdOlpn0TwOgP5f0/YluuxI8NP+W1E/
Lj7dQTKNDCsB1MTIuz5LwInAN/9hMXBVuPXgiT/zlf0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 37015     )
0a1BYVROhdCUg31LsS1Td3vbqClQbq6dcTdQkWXz1y9Tuunj6R/ybra3SYap1xpS
CXiJPRAx17iT232a4R+5x377s4Ct+Lq++a2vJViL9jy0dJsw534gE+wss66cYx8X
I89jYUQvxqE4IBjKIoSaFDnGAKnzE3tjRauWvbFXN5Z2Ku05hutxc4rp8d6ZQRkn
5zmvyFD9byHT0QImERznkfdZWu5l4T3oTut2bw4/ZVUUBsCBePz6tUHWFPBEUIWQ
x24KH5J3pfxUvLoo/+U61kH8uADyfU+mqU7EDJkK89LqmhwdU/ksSsA9TmdH3YgX
01XJC2piuPFnDAcsLKBnmdMf3IRNY5BZFNs2Z0IJ1gPuatOh2VV5EnzDOpxqN87f
wRj337HW+IyVLNhVgOteSKmsxekdX4de/c5iU2xULV536WS8ISZ0kJU94DTwgK1f
2MVpGExV+IhGuR8lOckoOeioP1JkgZyQJfgGuNKTGsjwoMfrJ8gdJKtRXjd0zW4P
mANf1e4WcAFdgbt6pYiQBWz3pjT+ylU3hsVOllelRoyHT9/2b2Wa8MygW5MgPDx6
7GjyX9Q8yei/h+DilwIp4tRaXs/nvvYEtBQ5rf/UQ0GRvK6dHL2pgyJIGGyDBBLz
MTV9HN3GqKIIeCF1QN7zc3Rx4SVnMC3CR1W3BupgNn7zTycg2Zcjr51nPtigPlUc
WCp8FgUhCVQrEHru/DiIj+ABX2NuI4wG6JTu/9XG88tt7X1iYAGHQaKDwk/9KfL1
IF+20YINgq1LjAPKGEnTUASp31j1AFnHBrsvRk/2kpedeXUukvHr+dHoeO4WOU9F
el2V9h5P/Yk2JcrbkAluCq2yFs8S0yr3cotE91KGX4Nqni1mv0anVNv+Iw8hZOW7
LmjhEmTkha1aZBPkEWlLqA/dCBr4rI9F4357zJMZ9IRADZteWWezOkAMqlvCaYmM
Uy7vkq9TI0NT/g+PJzqrDot3rtn94mlXKslaJ3noQbBhrzCoRe1OCLPeE4YNn3pz
OWDOPcLnrn21CUWUaRrnx0GldvJt6gxufzP09VQtBkGG51atel7saZUKeGI5/oFB
kz0a3k00ED3uRiHSu5Eq0CV5v313VzQ5+GlOBbFa8RkbkaXEVzaCpC19oBA5DN5Q
krJUwqL/odmq6RAhzML9e/H001bdJT9j9PUT+Q5ZMFuUM2RCtir7p/XUT99jD546
BY508Oj+EQT7ZODm/xFe96/iFQy73nVPMGsd3L+KdvUtQ7FQvEtctg538G7G55l3
NWtooymaLu4tgv7Ixz5VtzyCPPETEgBhL02/s8fB9nG5bJtGp16mFEZzT0M2QkQj
ClTmxunZ3KuAFbhuF8thYdtTWEexClF7RFW1owrug45UeYFwDv2AzC4R4ZlrDumC
C55s+J891LPM6tMN/NmAkK3Z/U+0LbVOdMaz+Qqxmt6hPyiYkqWV39CtnusoUisE
kIxe03DpV9gOPozQ3HnJRMue0ycaUCOyR5pRfUTNWjdTtSAQMyeo6jXICT/ND3qW
x/eTBD9ZxgxmlajrQJz/jFnIeXivwa/WBT7bONpB0nezpwWV8+KJnjKmlYVzHvHs
34gy9v209rrbl61V7zasxp+KfQspE//VwB7lRn23CWPuTL8WqZUaNYmbbdAdwtbt
xgw97TN+aVCE1JdcJRTLP8BagvU/FJTHqvUMETM33uzMDxEYkpSUshNbkOKi63Jg
YlnVoKteny3J6wW51rXb2tew81jn4lQ1PUN/G09Y43H7oOqaUYDz8UGtQbinuEi2
9KzoT+ch3Fgr5/5hgDdglMgIQ59X7Aw1zfFAS+DffTrzaS23liPRXQ62DVq6N05i
9SIYNNqSC8OgnXRJWZqaWc4fCIOH+Z5/EzK9pORJjZhd2hrwU240jGpYp9zwzl+2
XBOGCfMkEU8YIoVA3lyM8upG8nwClNHSBfs6pXHGJGT0aYD6MFY1YFq6NMj4TKz7
YCDS5mvJ7ywLme8eflr5qFgbLmEDz7QGlDYnanAqhDQ6fNUog/R4mYvcenMXAb9j
SDcGRO2i7FCDK+nfh83dPUZeZyXwgd7qozcIiea+Bu2QgacXHULKb9YkEtur6vjx
TcVb5P41KH3IHeJv60IH+wqlDO3k7jVMiEaBxgvSM2GcsoOSAyHcM5R4GAhffeC2
FyVXIAUKfDqRkviWZztB2L7FNm1dmtK+s0KJmrdMJlU6sVVVAsk/To+re9QSwK0N
V6AFp3yXqxnOG/7l2ft8EjpVlgxisNtuhH5xGSHL1elzmzHTe/1xNCENKD0rJZHb
w3UbDvdsFfQGhRsKjumVsxPzJJxSzDiK33iEMYJQt3HWNv/ZoO0mroOsINBLmKaI
f73BlHzSkciZGsV1HocSiDUS4+WrJyep5YZ8UGH8yK22TznK3aMoAphac4MnX4Bt
I7VdSK6EkW67CWmv1B8qGvqysRYGnFtkK+CzvApK876Ks9DnU0SXxrnXN8cy0Z7N
1PD+CnqWJE0BMu8lFXiZ2ctEG4wIYJ1CGBZAWdCbOo1oet7aLWyjc3cS5dSmUNqs
uzoumqqRWOBQxic64BLzZpkeBAX63OqcOWVAXV4zeduklMoWfdTMlQ4oWMEa4/Xd
RM4Aw+Ie7idBxeqp0/eESRkU/0UUEWRLkCQFawrezx4CjO/5t5tsx+mroa4eoz6C
AgAIIyOjspbHHp1epcVZuMDgY9sc+8mR/7c6DKdKS9ggG6k7t38NstSqSymxJCH6
10+/BrtX+sre9ijF7O2xVzNjwxR8CLFbukMxJVFFgSDg2isTCqidHQGQA/CdjMLB
SJ+fmROzFFoGPKSoUqtvyWYz1UnPVfJg+nriu2Jo9Edl+yiDRTI3eczkJZg7GPYY
VlTdYyIBlf82UgEq/jdNcQeS4yQtm5G7BAZMbSAh3y2w3sBXWcO1IncZ4km5xn+M
NsaDPKpx2XZgUTJFVei1yYG/sYgtLSDFEF63wtj9aAH2hrrXZTq6oWUWC6cSi82W
F8dM2ZRJpZSadrjMNsU3EwfEzNSOF3MJGsJ4KYywNAdYAdIY78l4u+ESY8Q9vuQ6
wdKldM7BIZc1M5f8UGnmgNz7N3csm2eihdY7exSIG8eXMSG9LepgqXFYT0J2BF/7
w3Gf7GAICqFLJunBs0X/N6twHl/iit2qRwMiTBqvJc9yJnFPULZUHndxWkRh0GE5
41/OHD9l2ZmCxfwHaV51rVJw/kFK4CgGxN9Ai7Hfo919f4e7LP+GPxuep2omr72e
A9ejCpeL7rfOcFUkHQmTmeGsjSQnoLMh8AGJ7W5shg4iqaIqEmORf/rk5M2ThKzm
yhnAM6D8iA2wZIo5HMTWnLsYA9IbnnXrqrXGCIod+7qV5nmNYhn3ny+qklUEf1SZ
wnY7EbARuHIxJTpdw1R6CI2tHFEUv/GKseNmZnKVN6OCuf25puAU3hHFrLZ49iEI
xsUSi05MOvAAgUjfXt7LVq9o//VGSy5hfGIp/pIEa0PcOUtPEJiYPFqt8uDnMI2Q
dwjbq41+w5fbyBuDFpnX/zXmaJqJztil6vG/MJYWwzQ8aZbLNpc7VOw4kRpqksmc
AtVlL5qk1lV1om9q1Q4pgy0pUa2gR1ad7lNwIeBi9sHgCQ7EEzBuw9PzckSA2cmu
kwApRlJ18kXjWD1ea1W2Tq3d+axEvd0YqoBjrWQyl/SqlAQcRgl7Se9ootm1ZY9e
fNAC4pf/4x09+xGsEcnPzxtFWB/IE9u3sn8y5rS2sRk5By2t4hCURaFz8hGmXTpF
hyYkkrVE4tQpplZSjQP/Wj+vFlvvsf93Lv/07iFPF+vQxXEdapJ/iGzxEhRI0X9E
TtPyjh0BW7BpnKZpEiWkn33BAha5G0mbmYuC5b7km/mQoreo6TKUZMN7dO5oUjJr
4CcnhkB0I6r5la3eYKQ+16QWxJ9vM+nXHSfbESSRvV7cLFhC1oK0xMW8uoEAUi7T
l8WVj0nxuR7Hm1U4nl2PgQ==
`pragma protect end_protected    

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
fsSGMUGYzrg7QgQcMo1jovYVrYmNTswWzTO9wWlPV1Zb+10Y80o+s+DwG28fMoQK
rmTGlUqJOOSABtLgyRXrRyMlRkI/OrZQ5AMiu6v+HeiYIpWzWGLa5EOY+5BIm7Bh
otZZmp2hpISGbqKYQyD1Ppz3dS2RJaM5rkSeVwp7Vnw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 37200     )
36UyrGcTCVlxQBD8WnQDUjtEKh2YhaBbX9cQ9aMWz8t3Np8Q6ckSGH/jVuV7UGtD
7A9lZtn5/OfIhK+CurX/7hjbgcyOKPxaloRViIlKhYoZ8S+hTD/MakGBV6naV9HM
1FmG3LhjsgkZ298JNhcCVKVGRFajHs7x5f72rFd8FTSkk7kyPT3/886spor6a3qx
vtD/zs/STJYlD2UHoBY3rd0jci1e9Ceua2w2VQwQ6qJNapmhN5y06+y2iYrDQBm0
`pragma protect end_protected    
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
GACqHPiuJ8mPYdJzpxJ6YL4jRZE5Mll3B+LieDveCbs00skMkHGyQY5+wuuUNdY+
FaCz0+Kf3WJh4IMn1pqSTqsRnphWGpIMzQuxTuf2AaXwXivD9rnyMX95sZt5vsF5
+IuiiY2WwgwqbDXcArxByzYpNTNzXHg0xwuPDdKnEV8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 50528     )
umWlYHA3Gwa6zQn9Dav4a8yhSE7b7qwYfuW/GFoj7vbogXoQx959oCYxgTAdTuFn
MKXjAtn28OGCqCwJoc/OouATG63woae3yE+cUoTbjKAr7YKb6TB+1PsbOBYFjAbN
H6NYq64Euwy6LksCmoHnheiqC4Xv9pRH2tDSedAj4VHYPJBkYZvZUdLgO+zDMoDP
FtI2JTY4yodrAxeFRL13yfYb4g1cqeYDiijiADQh7F0JRqACAzfTqMqFsXfEsvC/
qVixGHmkrAXX1UQTa907i3sUlqrbmcKEU4JxI6QOQqsD1ZdyXaBVZ9VaIWXc0cba
FwH7aFyTSOQYSRDjEPMpPgXuj7vxVIkz6C0WySEmdutYD2J+fld+kp4Zp9rAk/tu
BIEJBC3cTgxPAkzxDJxGwubkS61pD2b5/W4dhziBRkIsIp0WEmM3METzZ/p/DMNi
Xt9zF1jmX7sdsOnDEJUOy9PzjKA/aen2Q30tVubrMKdgHAstqqwuNqdXKFp9rsXJ
EUFu0rbo5uyvCzJfu3BBtGo7SFBsn+XU2U8Q1bfYaaQobTMQRTKE2Ma/K9p95lpe
alSv36MGfgtEXa2SJhR/FR+ZL1Jq0ZoO9PZ5D7VcWjMR5ZcxpjFOVSKFwA+j6Udc
E3vyepDB+zzWW6APV/qWvudqJYbY44ueLUPfB5vy5BBRJVVxkv/TaGiMxSYdrmvq
5QNV7lsf/ImDeFReHdxgcMJ+3Nf4A8rd9BJiR6Gca/x+HMBSuplqF+RO+UnHqi0H
8UkIt4MDavhbZ6i2FshCdomaN0csQWd68SR1+33LUdzftoD/c17ONDYUYQ5GDWHe
MFJSL26gNBTyAI/fC9ahdLGchuWI8TZ0672fnb/MUfBBzehGQs1KNpkNmlQpplZg
xAMCg0FFvC8scepichpcBAoyofx9enfbXRZ1R6qWuO4NleAuhTQ8D4MI828Poyyd
cPzZ6Qpbu4w31W9K5jml227soiqicC3qOcRybf3a81v31l29SAcf/Gli9Y6tDGI1
9t78mNIBwnj728sIwliSB117ZiAY23QXzZKwC2yabrN2h/Fw1arY9ef6fj+6OAM5
xX4Y8q1/wFcWlR6bLsLiScvDqu/nm8WmNgjo7Rc4NUOFHLIceKCod7rlqv6pXLVN
UtgzYl8McAeE8nLxuh+mc1yxm4Nrkpvho5jQXa4G/KECJtQsE1K5Fbm/F4ebPOnE
+cuFg5pzoIPQ1GSOZVseufjxmo/VaUYgYaN46/9xV/y6yZhjARiZazvyUic1NtbP
0KtZP2CwVmgR5ShhLPpp1zfczQeyIytOSGX2zSRqAIt04appLI/0EuS4sy+/S3Kz
+aUb9Gjsx1n9Maovk5cqQRkZT6heXZDtvoofWC+gSeIo8766RV/8w9sOqtiiA2Lh
DwCzYOzi6VHullxdoo/JFGobpaXYbHcksNamsmYg3OoQXgzCG259ZsOU4fiFVqG6
aJ8/kn+w5Krtt6HUBO1OoCNqoSMfjWCxg9jmYoAvJNY2AsAQimeHkMpbtNijXMWl
OBwup4cvBBXT5Rodz5GXu8tDi9zLWqy9L5oIA2v1kDj9iQYARcYx9grZT2DLO5ak
E46dU2sdSsm7oJpb6uHa86BzdCbWL94qC4q6vSV+4bQnWcdcnonOdqBlTSNzQ8Hf
0ISVgsSCku+Y/dOz8KWgbww4K8452CzHDbg16PSizaQDhEsPH9f5iU4MYG6TGyOM
KSxVKAVD6sGvpsrAOc+lWxcslNK4wUG26r0TwQKqwCLIgMERc092WiP2Vb3URnUH
cK3/uHeoxEZ9jW7Rj6iVnDp9jwI8VU+fdHOQtEunaX1jHBKFao9ypuassyD7t+gc
BTJqev6OsB2mlP5b6KINfZmORj/MOQV3l8zWcqELhNskNWt4L34JPSkFASQEYvZS
Zhsu+fxyKihaF1XZxsYmhIJnoSKtMXuKJu6PFULgQdEngxFt7w+/TqkdeRFxR5iT
z96QLbVv6+NcgoojebJWc/uX+vv+IixgQxVnyBFrO2u2/dm+V5Rx4lWUx5D0Zk7e
ThINpIl4wTcl4/8tJYLevM9F94s/Met5SXR4IegU0mDadMOL1+V05IbDscTRwLUp
wsxMeLXHC2PF/TwAkAJWPTvon7z2spU1BICHLdsjG6lnBkW75/3aKzMdJPZS/hRt
F197z+uFN8MFno9dk9Zn69OYaJCI2AJFdtR5gxwCEXdFqg30jHj0NU9tonI/yaEC
yoQEucJRRgm3jYLEOCsISYDK1nj3AH1d0ln3zQlpZETZHjlXkz4Y4JJtTxjuKHYa
l8xIYNQj1EyE+pK5OSm/FzxxdqlVwZy/3zfa/DRKL03UQt6T+iA6yg4v8ya6N047
Vzam/PxsycRQ3TvoUx4KKZy3x+d5lo7ocX5QtC2w+KABGTlPjtsbdBo+8IsiTsTk
yy2A0X3u2+fCdaPtcB8s2yUc8ekPY8UrCfz4GRm43+qMI74GrWWYaub9j9mavaJz
OY5zq42lXeui8amITYLH7YJED89cZU7Xt8RV21IKJzph+bY6zgnK80rJemSVw1Ki
8dLSImdC8cJyJkQ0YXab7ffQgTe5tmDtpu6r6VSk9m4srNTkZvA/7CR5MgtTF01r
exvG0tvS4vPVxpgl0A1pZO1tm5ScZu7M+hzie8yF6KrxMgkbGhpBmyNfNTWkoN1c
eD45JOE3KiyUr1vjo/E0stOKjUQLlG0M27h8pppJH+swDyxo1nVqQu25f7DHHk+i
EfhIk8zERC1/at2TEzUc8tU3sqpqYZqfAxG/wXh6dEog/AGfVEHCDcnQq3+fRDgO
XwhJi4pllsYDcn6IeDB26CYn7rrpPXKySSBBawMAVxHFiwAfVcpqcjTR86bysaEN
TRvqdt5F9KrC7bsXcXwelWDsQPRy0aFRQFKuz2n/ywScl0JKE5zrW0e08p0tK2+3
MwV6TJFXzxQlLhz2VB+YJLksHRpik/2oW5Ashf/MOJGhAPKya+vLSIl7ljIJ9o+t
tu8l7aRHncKO6DnO9y62Ju7LqjT3nAR1+Mm4rtmh0eWG2E9NLHZiutLmoplJLCEV
CIAPSN8Sj7pYh7NafjmeuCJvrhuey7kwz3L/TMG9KFl9gh+FpSrf3vBmjx9F5rrO
SLPMELtRt8eLzcSqn+evCyWKY4MbWFbKMb6Bf2BbkuEWgKWzpswLXaQbQC84+oka
5XFCD2uTaNbMCg67JoCsE1m/MV/HotZsACU11X/852/t6O625Z3pgXedo0n0rbEA
J+MLGf6d1lwvPX6BQxYxIVCHDzLJmyU27QpbnBb1rKtkLFu65oEpQzl46Hl7b3Ad
iqtGc10h2PVU2FEl2reJX2QihGqL8v2ULemPfAiDJYlPuZxruRkflhEe7eu3rBRQ
1zRbO5IP9+/WpnN6gcx+Qqbdgl/5fklmqX2eaEGDQ9/jUgI1eW1V6hvwnmA2Zxpx
2wdAWQGMGQ5qt4dJEciivc6996xSaGw3NsJr5OuGk6if3ICiIXPKGV6HcM/gojm5
oz3VbdHdXXaP92T9jm0OXPccn+0/im4nNJbDHWiGC4VhUWdKjWpwXTe9+JAKMoZZ
WJRYI0/aWqBFmDsrfVWkPIQcw2AJ+LlllHYbrtbO4QFK6oDAxlgw2RH510qSNGPF
YKkKjLuqDVpsLMAutSrk9GTSFR7ueStIaIs8pyuvLJlyiiJrU2kctecitrZ0UdUO
bb5G8Uav4oCt+2/cjp6SuP9B4oTSv5RScpLSZCsueEsUA4sFxuIaMZ+SRIGiA4Yv
ssmI2wQs+iZ8xR9XZffNAp4cyglMQJ15/RBY48qFNqtVH/LBdbyPQVB8cl66RZe5
E/H13TbixSzeGp3cOL/fNwGq3TVXhxWRfV1Bex2T9Ai3A8xPmVXUpnwajI0IU+V/
DXmqfY8docXmQerf6aPnV/T8m8NSbcx3brJi8w3nuWrBZ0H6pG8Z2sSJUzJtXKH6
lelB9Agng1vZwbXROtFKlKb4cqlE7kh1m3dBMS98Qlj3i5EcVwLX6/8Ek7gbtjZC
N/O7LOErU/toHLABUWg9PEIqQIntXQJwuz9sA0Cv7l9A7XLTS2/uVUptElPWw0vS
cFZoW+a/kLyRtR/8c5GnWoD3bqPgE2We52idVq8BNZyCKezzrZrfyDHMR8VpAoZL
4Sfi8GTTsa+Tf7teJAnWkACUaRE0sgbRKQezdLsfMJpN6XQ/a+mQFeONTOjZddNY
0x5G4rvZaFiAGQvUOO2HBEVyn+Vs7hzuGFlu0iCJplCRv0iNdkqM8CZ6BAjvsXO7
1cDGk2qSIMq7769d7xkZivbKuRLM+2ntNUhC018e28+25/Qyi+VPgSki1ffhns3m
7tuTF3VUlkcKvzyysSbqPnImC6guPD7fo3ah/OCq/pYvOm1L9hutYuP2fk3P14eA
Uad/6N5VrdUP091VAZZsgTmF22DulMbewUCLuF59eINXHejkkwANexIbxj4SnJ1A
9wp77cnMQCRRitfeD0h7cHe0h4UFnnc4LesGk1R/Zsdz3qrLJAtJqBj4rKKm7lxG
o5q7qHnaX+K9lHEaHZh5oLbtaf9ZC967E5g2g6TwdRgeOb5Zp49c8v9EgP0+Juky
7JK/sDVxRKDTuABUK/8xJuUc/pdu4JZTdmwAeHKPLfko8m024X+RT2M/O+Goe+P3
MUl+Cfhw/ScKTMeebawn7MCHNBTiHzKoj8dEI3JyQU8OjRBMC6RzbqEaBchxojmS
o8x9byt0ngEBFPUAe28OwZ1zoDbve2GS0TrLPBFM/QbUjpOQcUpVC8tUC2Z7kYeL
bbphHkDomKM9vZU1No1QJL/Mn6DEwHcfdiEqfqWipi++a+OTHf1x7oeExl4K9r6y
2fLkq7TOttqtic21vTMbCFO0a7Fm/0w4/2AQpIgkp+uw1sXpv2SkTnTPV1IQqa24
x0sWMwjsfELuVazto+qa2hlB3VjGISt5fScfRXT8oNuPPlWTe24qoJclkJAfPedC
Sef6AnPTAh8CbeMNENPM8zy+OTWKdlrZVnP4LH9T5gSva/KPjVviZwQv+YRIHYu0
U58ZR1Mvz/d8mTPDM5V7wnAzpgvwt7PW8zrb/RKsbigWeybbjPKEhV/V2dn4etZb
5pPT1OP5UI05XKmLG9+dACQjx19JJoaEbK6HpZzsNhx2yiVpRhbj4MuNGF83+C/s
2qJVFVOE0Xz5SFXr2Xz/IpBGpBwUeGTL5E9OcrBX5Afc75R+p3TOtXm4FvljBvpZ
M+knvcQuEhZN/QNkabc69ITSCteiobG9PmSiWof4eR1353SpWN7EkLRkgjj1zU1o
PMkJsRbOb9wioOKTPcpurUuRYgqSykufcR8QKcaKhTFBZKw+KfVAXkC4f4Pck7l9
bZHfXmfWfMLPTUBhrc9MXlJzVgiqSFnTH/Ja4ZvJiQ+39sEA5KGKs/txuBP1OuDz
Q8JWbEdvtlSqNMjVDqNPVbCKEciJtavuVC/75eW2iOHElrY5GIGoO6ndYGloZgdQ
EEptbm061zcTKPNR5QH1bX14lz9SB6FMMTN9yDU50zcmJjhPYdAp6z3sy5NET0N0
gnbUUXvM3OMAriCCrjBaZGcaWCkEx+N46ApNMT8hEUtN98mR4Usx3yEaAzCLORwz
KX2UEq0l8WoBsVkdhAZZ/qgciUUnl/QqDPQbqKLTeo2BkzBNfD1rTP6sxk43bh9w
97qLlHXm2GI8SQZOkI0sOxYDe3HokXhbpX6TINRJuIusejc001R8f1On2+q+Oo2y
Va0/OXK2qPnugfL4WiwbuyCq3MN7m79MY6ar+8GSGTbc4vyhbjkRA0M2uGS3oxpf
y2jsQ7dRMHsVYLEC4wOs6woe+4eZi/3FccbfYlmS+IB63ftWb2bF24OtZCoYCRWK
VU4fdseMdwBcKcUWrNcBR6gRz+Z0ITDqWh246230UEohOL5o8duWzfQyqw010mrY
mSeC44H0hbRxqBHpWTrOjnp7r7IdC2K3Tym/CsM0XDe6kwPh+UkWsyP8r76S0AdJ
w8i/l7ty6nmqTTvEBjaJnZL8IF+afQHT4mqKQSmcJenX8VFdsLDu6EyJomrlrHMq
CfuC1QJp4ltHH4ATohJojzW2+9n54vgr7Zt1gADZvRB9iy1wSyPLH5u0FkhuUuwx
Bj8j8ow2bDks4d1LI2D9DFYxHl0PBQ8Z7LChlztOxu792i6HAKom9Ljgbimm8+kq
UCXVBvvnYkHyE6rfZbCflJu74rr9DpBw6UWCIhgMzQDDR/U4JGiZ9TcZ83fBojlY
yPSN7ThlKGZJer6bdDZ6KDob7RGY5F89CSo81gWYDQUr4R5R0oHilRg9QbvD8emk
P4iX/6+zH+av9zK5ROrxylolqGzKLc9d9LM+YbobAA8xHJ6sxATi1fmjq5PK7s0d
2jzF7t2W3oPqtqBoVmdlfh3Fr2ao/Zsj1XstvZDH90LYCJAaqm83grOIJ34NHIlQ
I1r95W5v+l58I+U44BDL0OfGGT294NMnrE7+89ytvdr4B10wa+obl2Tq2mC8Jqpq
BsQw8963nwooWn05QMv1kw+PTZi0BpgseIupuf/s0xWErLtA/Uj9T53kfhdKiuqc
rvb7tqTk585+2rOpMsOkM5kG/ThD63AfjlWeiSek4HqMmcXOa9phw75sVp0q+1GJ
sjEYuxtotNsW/FlUGCow9M0rXNTD20sXBY4ZHWrrzr3QArcatAkM4YkD/dvjBAEa
2eFxkAsw9/fUsAyT0pRT8KWUfpWzf63odA+CZ3l1HAeWonTwJTRdPfZjNJja4cNW
DNAlilLR6x+efLnAv+4w5p1p/Jocja3EgfvhxT33gGbp1QEB1UH7SvnH6hIJqsqr
jYBTUxxpm02n7jMFpL6qhC23U6pv1z9i0Hy2XaO9BSKKXl4HoJu2JMAnhfwuqtYv
V3Hbp1gaXluo/6cz8xmL91yTYshPCO5CoQvT+TDbwmQ9ciQsOch/Vc4kVu3vg0IE
BJTvEI97BiuAqL6slfC1CMoKSKo1B1yjCWX5EIjPBgEJns5Y9UreNhhK9vS8Ith8
rq/M2GN44+CfrpzxQflwQi5d+k+8yqzs92jkNKmqwPZi3Rl66CXWVUmt7LSlLYzN
JPONtd7WFFAwZm7bUdQc/KewDEpvnuzt3SXKvbgpJrjeVNVEYFrZeoB3+Z/0m8Zf
7DhJGIGSBbLqorzVJg2Ry5SmXudsio+t9btW2wDQNtBnO6dOhQEpqns2r3sdN20k
pXP69f9qu9TrQ45HUXyoIO1NnN/uL6Hkhx0eXgBQkBy/mKpGIU08cxdrZbi/KTDy
TTX4TBmOEKA07T2AXZb7ESTrObbwyerYKPAijtLnytDtoel3YFLSMRsRsGD5OhtM
yCU4qUajQZVcsZ6N15z6MImlYGteowHtCCyoncp8WjrQETiy74h1PY9V53R2lnip
bMQoKPxyFxEYSFetcNvGVGkuJRxMc9utfhi9wiNQ+9If94+kVmIURxvbpZ8+fHb0
xng6Bgf+eeAyyzCyny1finl6WLw5p3odPSoxBXS/y4PaQD/mKlTy7peWtCjb1swQ
kuXugRUR4kmVF5ePBaQVVrjeExPwj4vJEAvlRcmBWijrj6OD+B4gRQTmNW6W1spa
PJQIwxkS1Eu3melQYb0RpNCx2K/H4FZyxOP4GMP5OoAasQ9+fkxi/Pi+hV+YDwnc
B5JfEUqwCCFR1ca9qGhCqsji/wFmEXLW5MKltf0SJ23p1lv2u7On4A/OxhID+6En
QUgwn64Lygs4OSsBAHUYuNs8CCrbneIaQvsY1GxxYDNO0lPTSJlSBfkhGFk8RcR/
UHggaHHtnn7MuTlZKx9UapDa5pBRzafGih1jik3IRUZu1ebnizUzBJdUhyO6XaWK
XI/H5u91tCumrUn3RLnDHMjwyaZub9CnQKpgMCWcOR8sP4J49PmuKk49xJnyjdqG
Tuqp1wz/gX9wjZQkosjfyl3y1osKfOR2a/O/XuOJXzPxo9tPh6GkCq/W4WwoNE49
s+WZ5gg276LINRQcCC0p4WniWGlH9j9sFThIyKLTlooLUfYN06xU2bbG2OkfrIwp
DI3MrLMucWWtPZTm6ASNjnIKFHlTkEFroSeC561d99aeJuJp7gqWKrPVX5Dr32Tu
MWx2D5wlBTICk5vVsslExg6GOMDupFuXLa1Sr1A5GIE76NkZtOpq6APeRwRi9wp3
8057fY5QrlZI94Ixo9AR34VlI4p45LNU+uaI6ryBWDe6P3nL+UKGme1I7LNkvgFp
xnF4ghQjEHV5GzwUAzXj7e9oDgxSM8wpO35bJI3sFFGtbztn2lPtRTOWiarC5Zvf
aYB/ScjoXwc0IScEwhdF9wVE/jVplLJJuRcSsJKnQwLtNT9Vxc1jBusb3wccKQqz
1RSaZyuWoEsX6Bzm9+wdQSMgULcRmPR/UDSvLa+Gm1md6ri98kGltrc7oYCCpERx
vTGOkKSltD1JCzB241+Ux9mnnzYVBEbp+EZc7QPjQCu+m0EzbNNak80LkeKXa/jg
WMdiQqoAiyW/hz0a2QDHW+D+XXNCyzPu1F9fb288j3Zn/R3nqdf7eHdyHU9/ttsI
RzjMO+4xE25I3w1jwVtjX5VZIsFE7ReQV3xHUvGylb/mcFqMTYk0hA/pdAYiEBqE
OHsczQStTr7QaCCcIooKm8cuYFVD+iCHFbIIgQM7OVI3Cgrau1z+fhd47mzPgdNG
0FO6LCb56Vt5MOCrEack7GYJ++mQi9cgZo9xI2MA5TyaxXhgbhK75lTqz88KHEX/
ZlhZzA4mXcMNJG3a1c9j87XFj+pICVhddxi3B1kr6t1uyvIgDBej9QHex/ErJezp
mjp7PaKix3slw6qOFV4Ff/gpr6GzcsXTlvRLKDNszWRm0qbiQuCHFvAF4gYvfxQ3
ErXS/t+2KUOlSHxPME9JX/ZnnO4SgLFo7zzS0/fPmI+ya8uive1AITZOg6UDSrqD
OWDyfCu2DoxtxuTNxZSk3dWk8Kahzrf2yvORZNCp8d5Pmssk4YB5dss2pT51PTEo
JMco+r850zMsEvQEJH74mx0TwrQTs35ts0XmpwbsexOyRjN2Sl2Sv/E2DMjGzePZ
srCgoPO14ag4B5TSik/pRHATe7O5MtDM/8pXKQOov83e9IaJUQCY8nBD4bi8Am5y
BIHJkLD6VF2RtK+L48SFNJgqtvbHpvQBwrOTdZPn8lYfDdnjApYaX8yIT2sLh7KG
5ZzkFV5SYaW1NApzlW4Ztj8xTvR79QzJ9JZ14YpeYdCBGSOMRZPJqfXILAHpAYjZ
UBmdcKJ+lCbF7fedNy/4We+v9BCUTA0pa1auCKbKiB+Fee3EoUWzGTIFgxMRHcIO
2iF90NtnUOd1La/LbBCdUIZgu/OTCxgN864k2jZi3k1/DdEyAoQNH0p2zfV3BCew
IR4spD5I/a8z+lpNSzqDP+S+gm5z+YI3eCZwaLiag3AP9aMfMC0aSvBHFKiYXgGe
2AozT+v9ZwZz6wFFY+HG3xvikwweQO9p82294oZa+ilShv4/K7jQWFW5Y/0hYzPP
+9oKBKfWJAmWmzYiJ1xKLoKidSUKi8+RdfDDzyoKMw4RwobVLF27eOsb6IhKBtgE
jEEc8mktewjGZ15hPhnSAM96CWQDIN2LDVlxHCSh/QgOeW+4+4ELuwE5/V30cpvW
qlrK3tarOSAe41DG0ziqgulmNwhAj07K/n7c1u6yNGn9lr3dYLvhkvpzT/MRwHuu
tAfwfQJRsolCdxDcIAjNOACi6RbbeTTyFde2E4BQttD81mZhMxD0QBEfDMy/piC2
PsvrrSmQFKMKXl4cPPJ1mimkevbeoLVwHbqGfxKknxO3Ck7iaHRYTX8raNhis1GA
xKeIviWFT9XPtfqgTeeqlje5PosnUu3acMfZvfElBXWjQpPL1H1yAYnulr6dxkdx
c6pQfIWt1TNKzeyosf/EHH3KcugUPEinFb5F/wnQ2W3kUBGrsiIGi2ouCXktIP+f
mCVYm96c09m0FBk9ATzvKlwH474aVXNu7Sgi/qIUIaPL5TDWVqbM4rOii0OZ0fs1
1ixHWBMhwLt3/wzW0smKpF9bzx8bG068xVgqSmi2m6SjVDI2Mm+pkh/38xgNCkfH
FJvW92UbjoTnF1TUXIZNZrLO5ZenN9Hv4LVpY1iKAuj15Ddu0aFs4GmP+yg63ZXN
DEWuZQngMopgGXhltE7NWZWwKrpSYQVxP/5BNxH4AtE88SeFyXRb12QXxkUMUDnF
gVRO0FQNywcKSX7V/LUL5uUuyhG2IHRTtHheO9dOF3noIraiPib6Z709PNj8bpmw
3l3gRuGak2lpcKisAkzbgXg51bLwU0hf5DHSYddCrUapgWnzecMX/SXYHKHHXJ/K
bKpK/U7uBkM2zsgKWeAy7MG85pmbRiUt32d4mwbjAFC9ZF5Qsgsw+AUVxL/L8b+8
0FVd9cYfewMhNtIEKrkTcvCqSESKBIjWc61EdNLSMtuDBfQ/dv31SaX3BvMe8Yxs
8w0KAQuEd4X2MdJju98TQysbpNYIiyPEw/aVAvBv6W+MENaLTgNp+LPv9+mevhyp
O6x8Wg4rpz7B797KX4m4VzAxA0WWe4tIYS3N6hNJzSpBYogjtsm2Oh75PAbQ6VBB
k6InO83oKuosOK30L3cOgJO3PE+uD1TltbEkdMNn4R5eLstRbzmixBjan+8OHIYa
iyUZYgfAroOT2+V7uGTBEMaifqelKSvw338sd/cENqoK2SPxg1pQLuqaG+NgfIx6
Bx3fbFhTp5VguqRxdjMTHz0KSA1QTeyx66R76r3qaFUc/he/20LXWzN6c1scFmHp
7sD17dWVNhT6wEhNVTJrE7VJsbwwmy6R5aZpDicLnHNMeFIqtzxZRMp2eIeyoxkd
d0MqAYBfX6xLx3MG/biYmlMd/6ofUV9FPFjd+RW3PH1w05Zt1hgGk9E6IPdQJikz
eOVV4qYoHzlSVQPFCOZKSOGvuc7f4dE7GHNX4BCiZhoETN3MIHgUlucjiLOmyONa
pgDFfTFQ60784INIVhHw1I1nPOXKbmrdlDU+Fo27mECjJcjaaJVd+ZY79jMoIgTZ
2/jeoNiWrxx4vflXGQwI8VgHd1Pa+VuFtiZElhjITXnWRgBgijSuuNBGHM3/GHCm
x9N4UhG+JExfKEpbYhqe1UY+H2QVriONyJrHh5oQx4bbkUlTwcJGaBFDX0gndMNg
Ykok8juGgv4iKW0AFsI8rWhkC8u18lGA1eeZ72EcIiyOCavxD0hnTlNAM1pK1Jtg
MXWtDVKKnETB+e49Sl2e3KFGSI/B0GoNVEnOrD82n5p+w6xVbxDCSxXMBQz4B75u
bgzr7BWhO81//DVsEXDlt5RIec+1tN//P/d5wBGKxLYelcyMuA9Evm01qiDA1Ga3
nA8wsfLdxpo2IE5scvrP0ODuPVIgISYQ/SNgasguydCmNj1t89ug/7/oPh8DZRZ3
m0w4UW9bsXJ2zZvPxdFNiqkHMRSJSQ7BCnUdPjfmgwVhu0MkNR7YPQYb7R3dHNUh
5vm1XD7+HU65cj/JEsbb4umKn6NnYxaw5p693Zkl/2OwFPONIcLZhRxL6dN4T8U2
4wqEg6Z8WS1Na7/+bny7gXKgnSl8tBEUET33kUJyCL1dBUQ3R9I1lJUt6yIFrC2r
rVK1Fs54F6nknd4efLAa4AVqu/JedEcWcA5rlWW/1D5weklFCy0JmGDCfKYt+bIi
KD9kBbN6RnWznUwaUQ4mUl5ME/VT34VjoD6jdoZdu3Nn8sfPjIvS2JfGB9qjWhgU
M/5H0Q8XHk/1nSZo0YnFGUMCsQPJYtnSGm5cqcP7YmOIF8v806tmAShtr8B8iAnv
5AbUewkgNElrdxvVs/STKunkP6sFD72B0NozhfGsENiMxasozsLgY9rQXg5s/Ecl
HAYECEfuy36kJ+DP1Z065j9uxeIzlq96VtPf6l18KZ/qFKyqnIH8eK29aqJAFwVP
nLLRJZFv8tzwDxBeUGD4uxIFWKoDiMDqGx4CzSWdEqiaP9ywq9/O0vvyDTcrNJUz
0WQv8yfJbsV/wnN5V/1EAwDC93uylOm0xKQi3THY2/BoKUYYQEkAii+mRh02rbqr
PH5Zs2I2XFXRvX1wQlI/x2fiQcMd85fxv3qd27ANxupAUZXR3IxgZ0sER/UnJ2Si
ivQE5OWLB5YV2BN6o4hzXw1E0pUm128i6VW76eZHS8/ZmA3SxMe9WuifOk/DbPuh
gZQDQlMWO3YraC/vzNFUw+oAZ2z7nosQmY9dvY0GjhDn5imOEuUbzKlAVDaGpfFy
QlWI+CwIm8i84IhIbZXAVHyrgRYq+uQRmS6zn9zfECOnlPq2Zk5LLX/LEru94Dkp
Osp5F/mm2PBtsU4b3JO+6r5ihfl9LESDbXaWMmXZh/oUaNgKtSRbk/96jl/PT9e5
Z4dkUPXAVHFkV5q+Qy/k5E1O9UnR9bsRsreKrtpuTVTBJWID6Cw1TBG+jGnaV9tn
2XLwSHvk9BGLWK3DBQt0fUosEMJ/qL2SjUAovpwM54sb4hriT3PFqyNbXZE77Fo2
KlRpogReOyqwAu3gII7eBZ4yQ0Jbn67MPVsizjvfLvptrcDnfb5Ypb1d2KnnkClz
TPwr4np5gLrMMSftkzDl+8faUGzb43mJF1nKkCgUzoJdc4kXaEmnAfig5k3pKiak
gcKVrSGxMnSptESUu2K2ordfVOW9PRjVihzJD4WR036U1SLM/7FoVJWzpNPjkcfY
YNR4gO3YAfGnvDmcIE2mhEhpw2S+N9MWqxeof8BOegNhBt4IL8D3wqXmlRVsTGx5
H174Qw8ZL5hXKsUus7XkovUw/liC/2A4MgEMRUSdf1zMaAq/8izG+5zbXUKX26QX
KIY0gJmBhUIlp5X3HoX4iVoYvXUkRUg7WlhJYkaHvxI7vv1I+jUvYgOhcib9lNaf
q0uLfqC8QzK6PtyxDbQWCE9BpBprfc26dpInFROvc3UcA6XovEmU1urMlHbjAnaN
M8jlJmlNM7H3ARLMhjBxUAhiJ701p0e/SlgOD29pNLjANWaVBCtx6dSR1/oZSBEV
v8cap9tZ13UxagP0K/Y6S7Y5HgHLrAltjv9nEHUYn0bc7MBv8+W3Q85IEjc09qx4
nMKYGk6BTniQW7H6OEL4zsazEK+DA5JHta/Y56bBl1Sc1sTtNfg5cdxpDSYFkLUJ
4GG1i/saxbXunoZvq7MpaVpt2TVCaIKj0sIJmV5SbKbK/ZRT/E/qhxtwQnlr9wgY
czQbSkpW5YOJyHm3uZXHqBCQiVdTTROLRi0KYdEjXsnuqg+fEGk7Z8R/prsTSTg4
pbLGfBIgfRDZ+OpovdGKjUxhFmi5kzGGkw1NnjNFHVHDwSj1JW4pnL5F5K5kJJY1
uck2o5mE14YbOn8a8Ctz96rEh3ISJU/KGwIMSJoBIs27Yg0yPrMKVsl2X2Rx+Wji
ZUAkEOwtG84czWG1ncGeFNfj+ahGR6CZtgeuHH0wxPLQrU3SzqrViK0Zb/16WwZb
TxYo4bf/X9NUjckNi9iSzejqbP2+ghUidcPP7gg0P6/VMMgmPh4/UPEKkpf84YRo
WpPqLuL7L5e44UVjzRF/+CoKRL6uSpkts1CRuDsO1Ilo1prolLJQEdYFiXxoRpYF
VUEPUO/+U3ZntsqK6jMP3b5SmXmOgK7jx+PbgQU2m6P5V7bl/o8ZHzYLcNdhvXgx
zkm3FeRCg9n3m3xLqDSi3yQng0zh7A2jLkE1ttV6KVRizvjzUJJy9553nuxb92wS
2puKk4YpanMq1tDEnZtUvjQ2m9eNUBpu6dYGMLik7gDhQzF6/PVIUjBNcQbHElrw
0y6/9yux57L4j4t/s7EOrN5OZ03zupuk16DfU/JFFPtL7DwnEzFt2g2iK6XDN4Cu
iyQmMyiNkENiTEerhq2T/3Nadr5HjEWml1NXcbX6xSYgVoffjipkjEo/dY+UJ7uI
KgflV0scIkm5030xGlhznExmuS0BguqceZOS9rF7XcqHiqQd0lBkMRFudBtkx7yG
nMv0PvXpICDslN1szVGFURtW7Pm9JxlCwwK6f8tGOyDTo0rrbEk0qtgwPK5ARZW9
L+Xyd8mk77yPPU2RdgFOFHL+WvtyxJ74SnkORzsHXRIOAg/61EuRJI8KtBjsc0Vu
lEQAPJnpRSpxZ2PWALvsVIU+ADssZtE9nLtD5Lb+mKDwg2M1Kow7cmYvvUWzQweI
9tBGeXP1Q9MjywLvpHYJ778jIolsD0Htc8qySLfV4Ro9aVAwwivN0mJp39U2JKtP
Y+lasBB62sKpMcU6iKAht4d3n9JpzX6TqjIq9cv6zHLbEVU7w/LEMbny7jCbffdJ
NobBg+lAiB15BwScyDYeVGoTmJ3fLToblt1qhV24/zJrp1yz9sGXMvN0Ka8ifV8p
F/SSw9+/+bnJsJTibc+J0TaipMWC6S2sgup7XM2rQ9eU3AuqZFze/X96wzsyXWgk
cqAPVan36wrjq6p6N9qb0UN7i3a5z1GGBUObaXVS6ofkYTdHQBTk12HKYWUqaJJB
PzX9LSZKIQlgXBftqjyp9VVyBKvSIBaGm2vZacxpTI8P3Va0NWGlir0/f1YBGa0I
AMgpKYaZGZ+Sw6tQG0tRy8IIVD1uDAEZ8C1Uziy4K9LUN9r2Efyqtg89RXeOvtCX
TnjpltyOiTxQviLUcEEN7aYMngU4XpjezqrjSFO/1XwAaQ7JoEYYLLwlUXH2ve7B
rylSs/OopQNOBByawzCVu+l7g/YJ+oaq3UPxPSra43uX0dHRpp5V4RLaB74YnQdn
c+GHu3H17iffleDT6/KIwImX9ZY6PMBjBwqgM3SxU/ummuWAo71qBxpNp9uQOXiX
gxX65kQwKvY9jRMi/EP7qNNCY0u7ms/jiDmhKTuBZenspu8ZtB9qmax00odX5nhf
Qdkto807NBteCYi///FRwcq63KzZcEXMo9RuqWno+eISuNX8pTExCGz2At/xy0EE
vYW+9PxT8CWeADzLW8M9pT8iyP08ZVIscy+8L+ZMxh8ZI22kNyLpuPLcKaVfs2HI
xP+8QPZ7XaSh7pfFAQr6C5wPeII0Xk3h9OcbzTWXyzyJPkuQk7L8XMzdlo742jgr
tbInwQymCcI2DHjH7xRu8GO86iapR/pD4onvrxS9yA5ArE9S5NkI8aLg7gtwU9d0
Rojn9tL8qXIdKmB30Y6tX8tSP60xo1ylzKUW8AfKnqp1B2Imo98Z3cD3Qu5EAFRT
eCu5dn5daCQwH3iV9ltFoo8aDmQfdMnegOixnPPrTIONUSaGc95itosGrB7po7q5
q9DWhfD4dqE0dsyEpsBS7P4tRbh7EktI9liF5SZ5GgrY1eBzXaShF+asb7NBueg7
G8YRRLAktVG4jg6ILM6TMbuC1mMOBN9Ex4b/DC2aAiHtRxZJQDtAVfw9+LCKjfwu
itcq49doEUF7guPSzDQGgffm+3gJUy7OSdxSSJ/jk1+E+nXmhut0yPcLzxX63vO2
rrw2or165QR2hXkd8z4u87Fx8qIYGL/qRjmHPWc81EtFpcy5vuvx57ntjo2CdZe9
TnJxTq32aoHiOy419mjq7xi14DByTaMwAeX0S3zGgrFuuGV5voMQy3NMx0Jhvngq
BvTfet4sMJx0Vh0IDgcKIUsBWh42FNaxfLhUZ6d2Tzv8Ayhmpp8KNZF8JJqc4lgH
cniWu8VVF31EWZKsz5I7hnY9NVOM/wENnMqULYCbLIYnK8y1VH9lzpZRGJvXA8T8
DkRoIFwSA3hRtYYPWZvyEXf8de9QSsAcWTQYby0MXuZO5/yXycSToi6yHEcJg2kh
K9CC5Mw0hiaeJDmYa3ylHVI3bAo/07qC0ViSZlJi8R7em37YkqVUmH2QxGFh5gbs
/8OKs6w66ttVuYvA5uZAn/Y7EF6hsndQOMMSRbZtuF+Jo5FP8387Igli1kv2TD2T
5qrOAuIItFrpHO2HT4Jda0rV0RzVa8SKmPb2yjR5x7CBbxv8yyUSU5ggtOHM1LlQ
Runk/Ws2phQQ2sCO1gt5Re67i7Jyf0djFjJyFpw9zBZsGsxhL64cr9O8BQLzOvtH
WseoAuGvOQ5zqO9c1C6P07AuXHHViBA8BLAKtqiUt4e4CxbdS/OfynSR2KEJQxFr
jMKIWILNCJpct1qii8VI6TvrNRVZPtRDkDoopQMRSPo4ACeLb4/mkBwxT0kF4f8t
mogMaHQaVA5n5P636YR4TkVuk1YB2mFnLQEnmUKFfRwN/qCf2CPKeU+dAtCUVgL5
FDmzyKvk5hG4tZvxofHebBMI9Y0LABH6xzQ8AoYSvVTGiDdJ64Ii80rxNtVI2NnG
PS+vMoyy0uB+ed2m4DkxhYtK3fTS8pMhiC3WRMcD/10R51qO7k5ZPIP2e+BN2Ykf
S4YSOm5CkEye35Zi0RIUMVmKtllgRBBK2yjJMrTMLofcuqpuORGA8Da7VSDCEAZS
GlUraQJdoX+cTHPIhN9g5+nq9oFK43Q3jE+A9CFKs/AqCkG+GWeaxtgc0VgV59wz
y0buOSAFzmkSeXLrXI1oStz0LvWHLHOhDtpQYUdK53cm/xrqRmVmorTnxVaf0DQj
BzvYPENHJoecM1nRwW0T33umP/kBm4qYRelgv/YWOl8t+ekd2mXv7GgeXO8lYZxD
f5lob1X/xAa2xtl1gl9/hnzy0N7FLqGUpF2ZmjgP7cxFEGcprpUPGon5B/lR/eHk
NP0/xPsUJiVDY2BB9hP2BmvWg1+Spx38YkOaA2bLP1jJHrxluATe2KKFKq3zBqpC
ImNybcskAyJyYSnGKXF6JP522DOcpvNX+ZcdpgLIQ/YMZDHo0jA3B12GQTqx0h3X
xO56SEizXYI+pR3cR5Bg+m59p+Ctz9iXPrPnL0joLSQ4NTEcv4LM+T2dBgDi+Mgd
9RlMMEYefxHxhVxCVffA505vMGJ/jqWX8MsDUYUlSaVaT0ePzRxZMoYaBtgfwyA6
kNLAiMoPjrZx0oEPOnm1d4Er3WEe3H66lKThPM4evOLN/pjeDTMResZ47QN3zsyZ
vajECLNwmmJg6g1nro2RUQ7AutXr7ccQFY1o1ZVrC44IOykPrpOydGDgXck8ougy
3Yxv4BCzlRGgNjqM51id12417w9DgD1qgv0HJ0f6nygvXvZXRJdXy7lwCEm1c+JF
3wq5cdIlFgYr0CsMJ40FElfW5af9X6kPKliZRQEBdzab7eqwpVGSQED36QTE7QCN
3O8U9HCkXxZgRnRcjSmdhmNpQRgj8fHOG+u0mBOVxLPAR5SPDN0xQz9WW0kUHP26
A907pCNfXRBR7f4cPbYLK4W+kY/Izke0frIByMHVO8eRWhvbxMmUD7i9TyhSVwSy
essbwKom9OX8+nkn/nh1CSAF0aAbfdSJPYpN+WUyQs2lC8SCiLhfrEdkHg5e0p+G
2ddfme3QqtUfAKsUWxp07DGKET9/zPjK+sE6ILJkfLH7JvvwUa0/1Sk49lSZgrV6
Y+aE9E5eqJ7dyaxEjSqs1SJUz4tRXoeARLJZ+KRJUp/pxjIZZCX94GFcF0XKL0uY
xuTfZagocK+jEwX3YhNqlZYa6/3v2HtgEvfauUrPgGJQxFugywnYuRmzTk7pfVYw
zze4x61XppnfQdYxCbPA7riGOwd7Ji615CVoPksoTOUAjTfoNFi9IxvGueES7dU/
/Z0p3vco1W0uW2xOLxr180AFK4CNabo3KCFjkn7eFpn78LdF7xF8ClZ++ahqfY+2
bHk9dI16ZFM8GWA9fagpA5ZafxOg22KHx0NM3KLU6h6RohxpH6yirkk78bHPW+Rf
`pragma protect end_protected
    
`ifdef SVT_UVM_TECHNOLOGY
   typedef uvm_tlm_fifo#(svt_ahb_master_transaction) svt_ahb_master_input_port_type;
`elsif SVT_OVM_TECHNOLOGY
   typedef tlm_fifo#(svt_ahb_master_transaction) svt_ahb_master_input_port_type;
`elsif SVT_VMM_TECHNOLOGY
  typedef vmm_channel_typed#(svt_ahb_master_transaction) svt_ahb_master_transaction_channel;
  typedef vmm_channel_typed#(svt_ahb_master_transaction) svt_ahb_master_input_port_type;
  `vmm_atomic_gen(svt_ahb_master_transaction, "VMM (Atomic) Generator for svt_ahb_master_transaction data objects")
  `vmm_scenario_gen(svt_ahb_master_transaction, "VMM (Scenario) Generator for svt_ahb_master_transaction data objects")
`endif 

`endif // GUARD_SVT_AHB_MASTER_TRANSACTION_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Rzpzkb5xuoJNt0s4uR0Ah0WfgKIiKEN96bFbkLgl7+HEluB98S7PVUPxBZiyLgUY
k17Ka5ibPi57LX3j2omj4tWB47O0NfiqLBUK+VCb4OMDmiTlzcxqy4z9QXHjtHh+
W/59KxFdreF+EUwA/c177iVDbeIjU8RQeQYpHGug82E=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 50611     )
uJWGiTrYjZgpS++GCvRDKy6VqAEE43ebIxCQGBzMsvufNbOSRoJ4PAiKFgwrcznL
ExkHFcvLwjPNpLn6HCFA4CGwxkdK1LcD3/c1qNlZc13Vh8GMQQ4e/lIx7f+UJGiZ
`pragma protect end_protected
