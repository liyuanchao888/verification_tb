
`ifndef GUARD_SVT_AXI_SLAVE_TRANSACTION_SV
`define GUARD_SVT_AXI_SLAVE_TRANSACTION_SV

`include "svt_axi_defines.svi"
/**
    The slave transaction class extends from the AXI transaction base class
    svt_axi_transaction. The slave transaction class contains the constraints
    for slave specific members in the base transaction class.
    svt_axi_slave_transaction is used for specifying slave response to the
    slave component. In addition to this, at the end of each transaction on the
    AXI port, the slave VIP component provides object of type
    svt_axi_slave_transaction from its analysis ports, in active and passive
    mode.
 */

typedef class svt_axi_port_configuration;

class svt_axi_slave_transaction extends svt_axi_transaction;
 
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  `ifdef SVT_VMM_TECHNOLOGY
    local static vmm_log shared_log = new("svt_axi_slave_transaction", "class" );
  `endif

  rand coherent_resp_type_enum coh_rresp_tmp;

  `ifdef INCA
  local rand svt_axi_port_configuration::axi_interface_type_enum slave_interface_type;
  local rand coherent_xact_type_enum slave_coherent_xact_type;
  local rand xact_type_enum slave_xact_type;
  `endif
 
  // ****************************************************************************
  // Constraints
  // ****************************************************************************
    
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
P5REtRpMZ3h7PiCB6KeAGAEbfVeY5rLvlOYD6ogvgatzvrgtA7+iedkEIO/Ue9fI
BT7diIqrMvtxtha5wGOnrsu+4mswdrjhWJ6tyK8coAoIs1u+viGN332B+14rRF91
YYcxzJLs7Me6Bko9hQOTZq4Q8NhHYhggIpoRlh+QtL92Gn8/unWpVg==
//pragma protect end_key_block
//pragma protect digest_block
Usd2GFjCKiUaZ0yVuUT2iWqPIeg=
//pragma protect end_digest_block
//pragma protect data_block
AtTCRX2OMNZgSttVXnri03HRx4seuVV+Lulw9eemc/ywRGNTvkmzb04tNzD+jWG4
r2/yXusyrgfjs4upsWioJL9EWMolXf8uhuiHiRS4esxVLbJAqMu6nATMOOM9/iwo
c7LlL+/VSxyfnqbDmX0r3aWRF3SbywQ3ESGQiX/g9asuEnNpHT0wsSAJK9F+t8RT
4LM8WxiIU/bUpBnbHtdcun/hXuiO0d3YcUwoakRscXwv3nFLCDPX7pYMs+JyaUiG
NBPuapKXrWdRj6Es8V8Tzbk96QdtMdtyivmI3S2xHpIm+b2Y8B0S/723Eydd+BmA
k+bXF2e1aMbjzDZQ519WDfCocDZH9anvSb2PDroKR1IbAUDdBg+LjX2FCv/UquMy
rjLXhTIHzwG7G4oyaWrh35+CyrHU+0AFo54xPwavBNaB79J0LXNFPokg/f9d43Wx
8hKgXXWZKLHmBT8dNF4nds8LsWEaoOTZXKXFEht9fv6PLu1NyWznU2Z5GRIqbKAM
wfo9UgVdvqIvlsd42K3mvlCTzIJDifAs9cC3XD2NwPY5MAB/nk54ZCUcg6TrGqvR
YxmacdCa3VPepVY1SrI/88+gkkIz/pG8c4QYxmAOg+KJWMcxRDFIrZYIdNLbrefZ
MG4VuO4GVjN+ijNANzbeJw==
//pragma protect end_data_block
//pragma protect digest_block
rq1iANNCUeXNCOt721p/DbJBEzY=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
DRZDa6esn0Os5YrNfi9JzXFbx1PrKot/xnuWaPkDkTcOblZkGFRJGfjUj0A5ONuw
npVw/KIrvl2iPxt426KZ72yE4fu7hTZ2/r7g5UZs+OCf4COuwZYWhZg+xo+xBAVY
wiJAcezcR0jnzP8874ni+BCp0bV44N/8lAIpiAHwngm29KJF6MDaPg==
//pragma protect end_key_block
//pragma protect digest_block
P6i0wlMYPmQrhiX6nISSzb0N1w4=
//pragma protect end_digest_block
//pragma protect data_block
C5ZB4gKpgUlSilR3ubI/5sq3rde4f/46+QwOHHSGzRG4Q4rlAqlBhM1pOfareFFy
+b+5MNdeF3+yfl/jlQH3qhHhHZfBTPU3YcySRFNf8b78xT+vEbXqC1vbBxgDygcR
oD5YS7yTc/fNRzl5gpraaQRPq0RfUVNxt8OElc/lQ8jm+CDfwPI+cKWaSktMc1xe
oPGxRpqG4VAZaOonuTcAJhoNWqjBI7wn7ebyS1fZcxtIjIarqwQc/ZrTW2JtrYKA
odv1gtmFNcNiZsetlbofCAfDa/SxrCGIwzCoIdEp793m/9jmq9N1XBwZq0Mk0d6c
o2szYo8xQ8YT1NfyUi0wIa7NruS2DAdhzMUpklmB4UzqDb/+2E7StQNMUqT8bxif
3qxKdPRa8HdfsNu9INdLrbb1Jz0GY/alyrRBxm9NToqcDYNxRyy4hxh+8tlDXOWK
dgTZ4FzQ9pZxXpAgtVBmCL57JFT2zVoVLhzapzNX+b9omRfjO3XQUPvvhKyYM3+a
2T0vseft8IfSqar0kVKpJaNiYb5gp0llhZkr/TBPZpjignOENATACRuqDc0AEFaa
bYs1RCz4eIgJUtoeJcPRO4wCI/YAOMpX7h2M1c2JWcopDKhtSO0WyJrAw/CNESHe
Qck8dV/r9TVt52HQtDJjgPuAnveWBnMoRO++mT/6gEu4tArGn4lmc+ZF2YUOwMfN
RKYYrB334l8iqnRbwrHEm8RvkIi/WNHhuxYXflYFjaznQHmHlowqZhF9b76C8Bus
Xj9LR3MZqloPZzXWrpL5qqHqWOHTipV52RBb2IakUSQchmeqaPyXwArWWEn+9fhX
zC1LyQYOb9yYZF21sqxJivUfEgfNiRqJyZaNTGYiMPyBeF+B4hHnUJRyvwpCdjjh
tdCzxU4/uUs46tMrZMWkWBe8rpnU5F+OW41IM7BE0aq/scjKRnwmh4Rzuje3TjEy
Er4UC28QWunpCBt6ryZ8SyEVY/rQw9SR8UTNumBdmgL57aHPhXMg3Ujys7fI9IgI
H/cXN/BPPzLlRxtGhm39Xg5T9MDVqDVfNJRkstkq4q48IdPsT/mGQfu4pMHDC7eg
j7LTChdmz0jRxtUHdk80rQGYUXxVV1psve+dwA5o46DQmqQZE08upRe4mEREmtTB
LneQv1nD3MbrkevELAxGFmzFStTVG/ZyKrQ0WEF/08b98udTMQ7TCsNUCvgqtPW4
XoYbSVXp9yVzgrxmV1iogpu5siNe9nyVtSVO2hX1p2jjOKeG08b2KksuoHnWyAHl
crnzBUXzcIKZQFzc4y++M8siRt/cdvFiOu9FYXxrHwSUn+LEUb8HG1i021CmbK4o
mzvBf95BsgVuckPLnjTxcraVtR3bd7SVK7rhGfm38trVJVk9G9mxpeZAAk0bLwoz
nsHxJ7UXZWg/jNtFRBwngf3NNtqEFOo0yUFUnzvucju84xFotzI6+CtCGVZK3H4v
3zQZYP8MsICTtQdQfjUdGKS4+G7BMpnjq7WqNasCfPYu1PVEQFtLDaJyKG9RLfck
cwG3MTvdGNbcWWjIe9q3wNCdqe63MoJgvJDawNkRuQhzxboBY+wgAVTE9cneUm1g
SFS4nWlUdCOe17bbS7fZHyjksRnbtd84yqv81LPQOIbyHaQ3yQiFArOj6XqYAlup
bjtnkytOKMBYG1E/Z//gN37vrJDdnNaET5ZpbCrdwRDTuNGQjzTi7Bm1O7obrrud
L7xMQNa3tsAe6FoDB763h7gXUdfzEbQI5eeH9OwgZ0FM9C4aTmexQY1nNmYqqQTq
FhLNTxn9+bk2RbUn47xo8tWEYxo2AU9BprQDm+lbZA38a+QMg2lyE5dhtZHa4qdT
EVSKMiBwd1Wn5eP8s7zSQBbS5Z0P4BETycWd5IM/sG3k9yu8aZdcDdwc4jNNUPCP
eWQQMLJHAQDln+GwR6HQToVm66nWgKDtQEWYx5sej3r+opeL+a7j6HLh0vXIZ8VS
WtGOO8kI2VEuJ8qsGghtDSgOHIwwM8V1OF8H9KE7jlZX+PVie7PIHxeUQL3we3zT
EdePyt5QuidUk2P7MAjVHZcc16avpXKe/ILe0WPi7w8ayySjsBWHS/6rms6id2Jj
I4fKpwvCpPK6IAd555aNS3pIwArAqcy27PArlVtcFx/yfgMVy2CvvHqE8tev7Ajh
tcBPJByLckwQCZsC5iHGn3AtpOH6AS1s8GKz+Eg64YYPLvmYilKzXHTzpMtt4a+a
u2rcTONO5dI761klcp+SpZFYGWZzcsd9E39IKdxelAfwVwgoT4rCrSpwgw5sLBH9
flgw+nGTXjShuiL4N2EIbQi8ufVp76N3MWm9S6v4CcRrDe5CUNfZdsqiSYW7TqyF
5mA6ITn6cc4eVTad5zpB/5+imGtDXkijYXK4gl3IrumNwrsBnHtiUSA9aatg1ud7
luocOdETnQH7M+cXBePJ+LxGDvacA8wULOuspblSY0BZU+4uf4/t563mPNS6289Q
tviIB5D0XTwWsV90GA8QTBwkwALI9L0O1LWgjIvMYroElcJpknpR/Du7q7/A5hY/
geL+LxggSz72r8MaORgON6SELeT3tH8UfyHGh5Jd9wEd1lJdu9mvDPF6edD3umYa
NUDf5gRwIfQfACgIz1XM3O8stdYD9oxMlhopqMXv8O+/6MzijgAVJIsRu8SqTWpt
IvT1TD4O84Puu+rffnkpMsuMyvba6O6CFuPV4x6oy3TTtbGieC320pl7/3/9+EJD
iKo9jML5Z5/cN6+yAd6o+aVa8ju2Y1hvCZ+P7eTPXKvj/dvNnpSd/l88xFOBhI4A
o9ba4hsW+ex7WLVUZLGirMN6AqLaAqLnO0zgVO7rvmDaK7xOiidjBUCn9pC/QFll
h2PIdMVxo9646b/rHtKRYKOXIla7FZIvCmbCaLE6/nt/yDyCaw4iQjUKv7A8zeBu
+/c9W7Uc7D2SRWtH5yJCqp8QktOUxD7GSU07WBidXoNhC98p00jDGKva0ylGz1sZ
93klr1M1ntujg7gWdq4ERewQPFRzbXVLjTqfkpgt98dljMjMFYTQuuAmLrZo9JZy
PNJKAQkjyUL/2YKcjtRnne6zTXn17D1B4G4T56N6y5EtyW9KWSBa4TJAD+nHJTyp
SPauEBKquEVLVP+QnZt6GA9hrnnZ6cCqqzPFmY6LPVxNGsNkzLmEJHRNdxaX2ddW
OtTm471Hd0oiO1ek0Gb4y2ida0lZyPykclOQlZtI8Er82lMmO0RNpT5+RdRIrhIm
tflY+ESRvd3sQ6mFwikLZXWMizPJ8o2ZB5i0PL+qeb1T+sGK9K+ixrBe5lYodlgM
LELvaigq0F8TGn6r3iMl3ijy/tX6vgQJ7A1yKHTXNJsyBUeNfSTqLw1O6ksPiXbf
+85QiJT7qOE74YlBsWSq3QJ5NkgLFarOEUTxMkWmVnjvYzCJHVU9du+1Da8YQSyG
DuZTJ9GEmb89CFswhzz6nEaawRiSrTmFqmDuDfYmxbqM/H8a4WGseZbmYAlhD6Ne
8gqzjXVx33TJbUf2R3DvCXpu4SVmkUiip+ahIBeizalfnh/04Ab/ur6S95Hs8KuC
wfCDVwgijIdu3M7LjmlBZ3gjB2XeKTP0m1zVui3q0q3RK/7wPrnJkuX/ANubjiFf
AGMvfb48briill93C4GBYUFRMkR3CLyr+s3wRYh1vayDXN0KdVkaJCxAPdB739mP
mRRbGgdTYrG5xlWTpbHWeZK9qlyXVvCqySj2z6HqeMRpsXPwGtWZqWR74Al+YdAh
kN5LEiPtJMOhy5yS8wHWN+knVGRs8IqxCVevQ3RZns8bi74UVbj6OvWQtPcH84HM
cpnaIrtrR+aw6wOrKNY4X5vvNZ6NEJN75GbtmQ0FnIlMU7lerQ3n93RPKbNnGHmA
bv2z+uEo5dynHtNqdO2WhAzOdm2kACL3TGLJAiV6MlY6gVqUoOH7aQB62fdKF68n
G1nnRZqAEyk5vB7j+GC0SBhNnL+2tZn1M32yBcMgXsUCK/qU9gwcGt8UE5yjd+ph
hIxj4QpLiPAN5+ODtG/qx4J7AG1NRpo6ofahkvbCCGStRsnx/bZDlyjgCrAyZ2Dp
GWqozemPdlbyXMG+Rs4qpjpLvESPGl3H+lDlE4m1WyU/h+Pp1ah5UNlm+Eu4jV45
hxVm8iQuBTvWUyP5vZselr5gPUnL1BLREoktPwMO8xNhZ2oJg0pUV0D+iPQ/uJpi
Bu0jK5F4/h5LPGeNlg/IbXM1nXyEfORLCVH+4+3xDkSqlg0MhF4QNAcnvqwBQRHm
FyGODnp+ZZJqckaigcVffoD9mkKbSFWnBVLQdRtQJzWi9uiPmLQc0IFYQcMxK3os
IboFZVRnzjFpTpLYtcGDAXkCkVmpnP/tXPYH/zNHbIAYius+1SHs5NQeknLyuMqq
/ovWZt0A0dC6mQT3jgpC0c1m0wtSFqGDt8KXciASrFJ1LKAWV2/ACrPRXU2v3mq5
kBNJFaIDweMWUP8WemsOPLJ4PcFlfkwqAzRcqDiH6Sg420nQBBQdcVMhZQKzu4AN
Ylt6QsriiISO2PYoW6jipvydMtw/U5BwjnJonipkAwA0BtJHc3U5CJtKMFkXKSGo
Tz3CYfCAp4lEXyJqClc2T9AtAExGw9jC+s+Tvp/ACvipItqn8UxonaE+kzIspwg0
d1OtSU7uOXTZgXK1q9hogD9IYEehxiNbj2VCu7idAyOxSFXQIXTzEAvZadUtTsvB
/idKujyA12twkmi8Vz5eKPqIU2MnjurV+HI9GHAc4YUfezUlSBnzfazW0Lk9Gdju
nQnl0k7WTMfQtJLKSvLZG8huNwj4yUnBOmMIqP4mzTgUL2UL4mKBThT83vvEBvSZ
jdV5LQN0bx2x9D01JPuysBGbOrpgkMIBb681UYTH5/5zdRfCKmN3cKpW4Q4R/Sdv
JZ7J2txgqyoYBrscYcbhy238QRw6eqx8fWJUTFCkX6731/VCTI8WSOCWC7V3ywEs
pFOIY8X2058o4hgEtI/cUgFvmr6RmjYdiGjsO8VizT9tvlEAaM/XwN25biCwYFyt
HAp8M90iecnPALmdY3GebCJsQnh6BogUmg1FYRpJTuuHz4uakPdH7pEz6Q1m+NvQ
zzmyaLq354BdzkZL/Y3M3u3cUtVEBMxWg8EfK+lmt55bhN+u2bCilxyJFr3hCeHU
T0cLhV1NgEI1OLNMwLm+JDlAI/bPKIqRhGc3pqnJ4oRAp6I2Uc/VxX5FnaeEIvnZ
XtVgNFsXhjnv/moNxwd9jrXFijsAz2vbyQ/Y+6J1KGxfy9L/ycFzV7o7oCSNaL2Y
9u7/jBBWMOkCRbEV8zF+0jsbfrA8iU4i2/lOx5e6V7cYLe3RjDExR/FCksdr2wdh
B/TNkwYRbnm3OSYN9+//esNuIrdtjAaFx8vN9kH5q8JlxM41R/HZMFJIcXA033tr
2B0EpNM4cy2voqqPLcax9DyFvNP2O243teOxtcUsCAR+lmZQrZn3cxGt+32zdBqH
v6qwGv7Lw5+kZsgcQohimomNCcb8tgDR1Q73xK6il1gy2KxQtavkNWT3uTQDTPdD
XxgfOG75GOdQe/UDjh0R+iAc/U5u15SCW7EyUkvpDdD/UWVLT0BZp5Ov3ruTZ7Ww
NdJcX6ymES4sZdBBbWPYTv23tYjpGLZEbHXcbYonx13gULWWk/YSt4nOU+xR5IOu
XsEoDNdFRL2An8mvyfLzmHtvR2fM0z4hcSlAkmpoND4MPcSEKKudXtzZeNaFMFc1
pFI6oJT5pesQcPvujXtO/wss9iI7JSaaokacNPb3LLkTB9rpICP6Aigkn2YocNWr
wyaEB4JmW1lkxJLsCVOvcf1FIqXl50FKtHys0FclpBfGpy20KFJJuNsb8T2ROCxi
i5KPeym6casmp14mtt7XkDaEKQTgPuAHcaygpzR+WaYPR1Fq8ZUnB3M3GVPUqNMi
JBddbhpGB1aUBiIj++jR6V1SN2HQUnIYNWDvSRUGomVrrWU2jJBQ4DWIS4oHSB2w
0xnHRa3mgmmnxnQLbWidGLm70yFz/Jk+ou3oZYUB5Gul7Xny6KJOXJ1hUqSp84aH
R1OOSjebS5RqKV1NLYb4KnvfrxUrYKnJiL2rw57dmiNqfpfa/cHENPqDEusQ28ry
m834ZMUt4mt2n22T/5JxXVnb5RvUYZ/DWXZyv/GDvesr8BTvr4raC+jEeOnV5o4L
CB8zcgAECSUr3w4aYucplI0PH2pNqPlGFLB9zTJObsWFIGuODgNzySdLb+7YJLyl
OAfzbmb8W9fNk7/7OsGuqNUX6byVRG+jTgmg19D0oDcm0VrSJb2O4BGuJqp1is8E
KUvxBiBex1HGcWShwjfIfMcds4AeIkIiu2WKffGdLVtkM2h6IPq3md76BPB2u7Hj
k7dcNVpWW23+qC40dWo9htzGx5mOkxA1+dQ5YIRHQuXdOa115GYt6GfWA+J+gef3
7s5ID8T2J3oAWCooMhzTq0ijvhiiWrkoFVD7Ieyn2KkBrf+Vkj6ej6Z3tY7vgsMA
VcD4O5OrCQczcep+DmW7w4SARusgwJDEGAM3ZKT3kd/L4trMLToclOFr8OzFxFw3
VCMb4UL5qWyX7zOT7HL5XK9ujNtEu/N9Gpi4TlbWv8nR7wscCoZxRUJgES2lu41V
QXkRuxbwOOtZdCZ72QbBjEI6DZhSg6U6x7hVWIandDNefpVpx1gR+mDNoRZVqDaH
uPSQjl5rBe2CIKs/TrccAqzqOKsiwNB37MpvYj0t/xz/MibWaQ2PHrF4ncdLJiiQ
TtFBYezY0b97gB94h7M3Nnxa42zu1TEhCkZ17NasJ4aZ2MNizBnUof0GgS6kEZj/
nTg70bGvoHIQ/6fV74DLtQrfhqSndxPT6U8wb2i4UNUGf9BCu3RxPh1rpv1S+4a4
ItrrVSUbDkG3pOH1rxmHzXThAksvqNw8skOsVmCJpdlwGyNEo/bFakVh+FaNdmmc
7QohKiLkhEdEpklqrK2PuSqWokjoedZ8YyZGcOI9VxKEno3zXc1/xbEZ4PBDKyF+
5xkTBveysPWWWC4PkEfZS/+8wtt31jtzJGQ26hTR4KGNFKaY67IVaJrOgP3bdPoW
qCNFNKSZ348n3ZA4WeKDkVxeQ94ZX8Wi7jCrWIVRyj5zscmVSN95Rh76qvcdzdkH
wLnUOWZCghQT0QNB21hEiiU7UF208L1TViExOsoaMKcwNra3JJbHwW6dd6yYUcvt
tq+cCfWOSFDP2+qHFoimgXuv6o6fGa/qG8oSOrcmQTSASvDKFtsi3K+RMC89wJQi
72wuaekTmwnZf9317Eojr+xkAyDe73Jldmwif8QhfCUMfKymN9nWs4JKPeDL+Xrl
WMBk8MR7YjVXmQhc5R7j/KF6lup85Nle+8UTxglUign/skpVGZvdUAqItNXKjEnM
BPm5VTC3rXNFyS9Fk7ryOq36jksKAhsAhWpQwqWeGXVXllaAxXoU7WviXqva8qBJ
Rc8ExvChGZGJ/lQKVrB/hcCfpJsq23oBfiPVfUUgpSpt7fSFqUx55u0EU6acmPlH
NcCHfrgvkf5lgeFt9/u5qx09lmSo1uloeuLxHZ6KP9phIPYa9098WEt9jsgnOnDC
3pPGG5qqiTeATgMgk2rohVfWl5X6TqHwNthqBdN567iYhbMDBLnkdpDjnKTfvaCr
fW32SgN+00/V0weILHND0FyKLCtsNIXe0F34Vnfi/NRk8Q2siVyvEcRcjPCHLxEP
PACvs2gPyStQ0uqH8o5exqRiiFrydF3rYghyg5s7XJ1+r80Ay7NwHJV01l9/8Rz+
EqVkVqdlPPFjS1sle8yVcWchi9XICtvy5hZlBUokskOerq5NdsVLQXkiMYkR+iOH
xH94nYmO0+AEvJzNilQ2WtJvA8Vry2znLulSYdWbvDVpPqP0mtCMbS79zQwwljT+
bZaJOnNp1JqLE/om+dZaCWpD/tEG0623BjYwBwpSbXhCyJIPSo+PRM8hkdDQpOLM
+nPdZ3BMpyPhsukeFZ2rTTl8Jy66GrR8qs+FAgF83O9uOmrP6Dj/tDHXj3e3oiI/
n/zOGNj3MalGtAkgYDVpSadtJbkvn72JguIdeLU9XsDxTqURAufTHaXHPrTSyg8o
ixk4qtm1YphS6xCE+JANzwQ2QVOfWEbBxxn1iVI4uVjOo6jJuPqBZQ+7tYOJDV0z
y8D8BkYje9y2GVgy2kWNjHsasX1O/jcvCxSKJZejDfCIc3cLigeOt+ByAmzdbgue
1wU4LTbmOrG/gTcQLuJpVvIb8DUjpPOGGjvjWmikou9f1hKjfBX5j1bK04wgPIzb
lNl499fjTzcye5h0j+Oa0ZJYjyT1YHq3q8x09d5G9s1fAuWHE4yX0io08Z9aalJE
BDk7qL3Ed7mzc4ztBg2R3kixhVCy4QQg583fUN2s/tEnDVUbtPNhjNGp+efxE1TR
88xlEOX/dcG8QQTeu/QRK9uIGUSw4u5i/+4oiXaWtlZoeqKd1qGhK5Io8ZANFjzG
xSSkJqJCWv6+7s41BP4DOJxNZz/EHE/K7YiEcZr1akgqicxejU7nER1VBA6r1x0H
PTShk43S7Cq3i5UePxUhLaLp7LU1sDIWieAZZ5k97+SYnUc7/tu4eL5A4SV3m/hu
4MzU0prVjJccLctzOh+ySpmKK57D+L+6sZKs/iOcFjusm20qTYcbZwJC0eaRNVAZ
wflqc2444bEfo1Q7cZ7eD+PHPiX8yDYNaitE1W6mkWhNRc9jlLrruAHvKKzwCSkO
mN667q649NLJb0ecb5Dq+/1/54T8UY99EpHWiGAdKgYCAwfGQkXNVc2HHJh3Py2Q
uzqwz576cSGLecDGLWPMsrE7mm7bzqi7wiM0OoxsIBCLuwDpAbS+PWJBnpkRt130
tAVY6K93GpTdUSBdOtQlJgcKGATL7gN1hhDQKZEdbOddR9Ch2YH0LLmpUQhPRmkX
m1PA9aJq6G3uNJy0HQy9sZVgx4z9Z8I/Wms1gz6lPEGE9qogITs5t71qCASuHVpp
oRstu2oMwZ2cN4IRGKwrasQvTe5upSQlWJl5JK9UIkGs9pOJGODr97N4Fp+YsVEL
+/y0613KTqOL2wUaikybaxug3H0o7ZOcRJQYNxqa1onmSjun2ZFeANnQ9g9mP+2L
TgvzCegisioId/lAnoTL5aoeDJ3eXXdfk8lXdKPazDPMR4Ek/LqGQ8M3ibXVSiP7
3qqTmSvaAaLh+LIsrZ6szrvTNTI5cA0tzGLAQRueQ6RhKW73aro/Dybgc9sE3098
2uoypRjxw4T1PllOYqVbchQXVrgRRwgczssicf3Me9svZGS8be7aeBNbIb66+8Lz
eudbiCH/SAP+YNbJlsbO02+ecIGUbzlT6QUq7OPD3dKVgODPNzdVW+PJNuSc0+Pa
7zuiN6SDvjdNhkdWEYTObcDlpjhOZD8iLefTm2pid0adh4ohHy9m5T2UEwWSSXkO
DeaWp/oAXEWxQ7JrBWcByjhuqNXcygP01iAfz/sx8qvTjuFqaUXarcDJruoOLfjx
x5e44cFS8xRK+Hzl31y56kVjf2iSxKZyh7z9Sy31BkKRDyvBAbUSoN3pdaBMtVqs
NPLoHGboGhCAcVby0pPxmQ/c5JfxVNehnS49IGx3qVy+8rsB+iET0P+g4YFeZFqz
R4A6ltiil43jw06OwVn/biYstl1ZMd7c7w7JVKPx8c56DHyDMG4PCSN4AyzVlgbV
n2vaGBnTcLc4SBk2Id/a+3r1DGmOaVCw8SkBKdICbjeanwYKP2C/ombm6WpdBwLv
XcDWOuZpfFa6vaLox0LPcWjaYu/qC38kQSLyj3MocOX6YWmabzKjOJx4j8LIdgRS
vC7vHQxNCYQ553rCA37blfLgeRN+thSQ4vvcCiElISxdsTiRuP6Ta9Fx7oYOks6J
DaRE8yQ7lP6x7Xz7jDSvdvdKqh5v5oMDuJEI7cX4EUeciMafGJPsaiPQAOyeC/nj
PO6Bn5iTde2rX4IBtkYpio0n3lqn+9lk5JQgSDsRIZX3U93zGHRSydVu1yvFo4th
SYelwC9ixgdgpRLbOJg3jtYy/K/Jw1RLgusYUmMDxXqBPMDCrsT9R9BJFWeSQsQ+
DF2lzJ2/G9NSK0pYfAat5noAPgnsUFDyGdSfLAdbmBfdyCLIdXQmxwM8GyV4MbJ3
Vd5ly1ZIYVj2NY2QShJ6nhcWtT7UAdxjUd7adcg1VkddkZYw0RCU89Ty0If6XvVx
fIZ/J8HN8na1dH5iOSVzdTlb3e1BEe2H8gPuHOZe59qKgInrBIpt7Yigr+a7eRJ7
JC5k/Z7qBZU15ZXjnT+hkvI5023IJZpKH8qZUoeNKJQrtARNsQrAj8sk7PJE3AF/
qabf4xfXNsxnYN9YSx6/DYZPd8kttNXCaDmgbcbRGaQI1uhYuNfo+o8rx/ecQ1Ay
XnRwbdyVMlZOqmuiUDhXqkbCpNpRNuaafFWEyscJJatwhgS96miq9z6+Ni5178An
d88zTqcK9cQ0SM0sOtw3e1iJfwJDlMvCOjiatk6Tf9JoVwJHia5aHnOhzAjfN1vS
NsS6//ixXlR+5nF6Cht0e35PA2b0/tMl2Flpr5C5gmQSONYfrqFChv3RFXjITZ9W
tWx1YCItssBax1XDtMzVhnTADW1PfyyRVAP118k/q3xuJC9EhZhTdRn9+U97kBJ2
tL875DQFgUeQuSScsZFjjfNYNn8timCla4zGl9ZgoSS/vqIlehl4qXJN2wTvN5Od
D4WtSoWKhBevUq5rprbq/Cwbu8LCbSSte7I6nP1Wrfhpt2JPuUgIKCsoF4QlS5LN
R4mCzTt2gRzpgfu0pDUnT/vaqZhVDH8Ig8lHavdttnKDuscgCJGh+RMNajYhtapU
Au+dZ5C4fK1tQ8FPXHQJfqWAjHb84NQq+fstYIUhZiYNHkkyj5dnrPWVbnVtp6Ae
XNVVDA/OuyeBDIuWrffthC2GyjmTX9HbzBHQHlb+VgJJSh8Q4nMsBR94UUuYR7CB
/+yodHfIh6KBukB/5y/U6N6E3I8GQ7jOUBEfdvVKXKmBD0zceveCWDQzZSj3eXr7
rnULrZyYE/CC1p9F0CZ+thNTVLLTNzBPcVDEEqE4V0VFl9l0JJalWM1DfwA/OfZi
2PaAjduYQirW2/TAM6pmbYiHfYNQ418oeNWg1ZYJ9gE5WGkpuyB6qwr8N/eBlisH
KkfuQE0jCx/hb/OVaf8krPXtsCp7eS4UjEFMppVzoiCMWTTWNFI48K83zZ4g+Ksy
h4KsJwGcYQEZ/LTd9ZNg3ykQPg9yVgLfeXxVUPI0i+/XTwcMkZwoJ2cd+sguROIR
EGs1UjKc/QVmgJYiDzmE9ZNmymEHwxiXYGJDGVAKBr4L4LAUPvbF30paIcN19Wjp
ujIWuP3Ooy/zb57ONs4CNxQFXpZdca0GrltOf+RWM5eMFUCVmMS4cIkAMgYW8Ymj
oGC3uKyODo3a8Jc6/nl/HlKM8SLcXqSC1lPxOygMcWWBBqCWqTiRBOqr1zbNwwWz
MtjzC58q3aanTeQM1f9up++c5kvQMYme/VdkIymBJ5HqkVeOE6N15McLCxWrEjzP
y+PMGxfA2ZEocKcMtIFHzuXdD7QqaLPMm79u4e/iYJraw/7Efdf4DZzx+cebDH80
hGokVIr0ULn4xrRQqVDOmJsxVJU1QDsSiMwsoaUbxoaN2uEBvunxS3tpsbF3KPue
ggA7Rblm4PZNS2mbqqhvAlcLBKIJp3YYxFpregNFzhsPgLXlF+RUAawf7hgQpvIh
DDlpdghiN/dopCipIDM6rmKlSfvnEEdpoQ7KIRAhSFC7veLfWq6G14toP9Joz6Tt
ZVLCzbpqRfuMFIzkomkpKJj7XisRVXpTw/wEf4AuUnmwxusmX8UsocDhTNdnJMSN
N9jiegGs1gNrLmydQhif+n0AJuAhRzGP1smCD0VZUr33vFzZzWm8tLoqxZCavooS
yEXjS685tXI/8MIdi1QATA5XAM+cheL2EHoE9lZ7AHnjJbkt+Y/fjpxRW4Z1qV30
/yfKvinLuJXO+6cIlBywzA51xq+PryStY67y4F5SpENrQ51obyglDGw5jrOSSUj3
XVKC/lqiM74aufv3HQjdAoe7ewJTbWus3q6A6hzVyunU0OoHlVAx1ybHm98oX3/t
ThDmfB9FJ4jF0qi/UIq8mOGQLxOjgu4vOrkBt3G89z5WYIX7bMSK0zTlpAqPO/Q+
ZBKZh1CjQXY+31wUxQzwIPPJo9BecY/fFlYpYbXZfai7WQpX9ABe08QjoETPQLUb
8GyZpryJ/560+A8EXKr7Z0hK4nyNk9OtU/vADI64rsUojBen1MbKEwLrJwS5radz
nTZOnLYeCSvfYcWRrX3dB4VtKqPl6ti0LoceOSUO6LQo9LGHmI1t2NpRttwtNvKr
8zqEapLOANQ4cJ0vOA/I3aJRq/tXO+/u0nwdh6PKLE6Oo7VBDXP6ie6aWlOejGub
Lsph1ae1Sk7Em+hfyobdbWR+pWOmvgmTEdrXPfRSpBs5rHs+fudDhDiv73FVd1Zn
TaXHCey+6iqZ/+K4NUkElkgD1zi2oOGjYiP2MJm4yPgrD25DenAcrGxrix8NmpRc
4sZryM6Eo3bLxx53LRLzbiM/tJDW2ljYJVIJwtbTH4PsXT/W+IkUjHdsMTyjAeL8
NVKd5H23aAT4yYFBm5UBlUsKQuTvc38FMbFPoDr9lw0SR2ObRPtn5SNrj1waZpnl
nTpTCdxzkc8h0eaw9h57/lzpmhIzxkwonOIBBuptEY6PXYUfworiYtboBkK7d2qT
St++KgboH9nFXJE4//LdYtT12rg/YCgOhodCfFcU8+BiiZqVmXJfeyw0AbwnwMdm
/3lvoJoepOFhhnEvfi9Ktotdr9iPMeMJ4a6iaRMQeXV9CE+sOcVuQUnGc8CP/yS6
RSY3sUg6fMJciL5xBZYIzqEI1A+GZ+sQd56nucLtSjmb2GdBrTVqxk1TWdT2UOrL
cZh6aM4/dGbD+dT/F/bAp0sW+J+HA4QE0VYP9guudzeNrM5yQtR1IfGouX0oc2u0
FQC5w50MtGEWeWZd3mD6tlfeynRSQ3PLSaatzinyAr6xSVCO1MtE3EiyUYqjE2aE
gxzSvgYgkfbLBsw1RfCaurxkhCszT8f4yTj6Y+5bcX06BqWwLb7OCthGbgt4cpbR
Gck79JFfN6Zd36HuXY3AM+rHfsvfnh3lVWz6dQTUaxQHqZamo1/7bL95vsHyn3k1
71CbYhcbI2oFbNXOnKh9MIHqSqdFzendQf/s/yPjnSBFpm2XzX1wWr931mTL2+1X
zUfIdI4yiZtQ25gCVDt4USsMS6skS2GRgiTYFoMSYN41v2PNfUzDBoym0Sb417KA
CYGwmods3zVCqMxmk1tmR+9btrYZ1YZAFz9bfVkFmjwhHWrJ7Ul39gTRPFj0W4PG
3vEYgi6Pgpy+L6NsjEO9k9eRAT1We/o7bAE0peuLhvG0oyjeNgl2ne0T+yrT5t5J
AD15wOdN6ZDivMmV4PriP6Vr017EZdAwuYotmeimf4a88Sq/465qRqOmdXw+sLjp
zMuWSzDjEF4jCUXZsWi4ec1I+AvImn+oE3MoeTVBiULPd+f1ou0vQenari7NXjz3
d2NrELQIQy4LVQw+YZhk7IWUCVS5RtD2a80r8/mgZsS5VkOrJ4osphSzykOIFaen
BEyP2GRpOfpxDrck7Sf4C6SWmi5Gi/C67qE4eHAHQYa7MqD4Ct0JCK/5SLjYIyAf
XRW5fXoUmlFBEEFAnPGRcQsSkqgSsAv0TSuWkNlKm851asPmZQ4wPRWVt14TCf4U
C6ISfiV3MWgM9e8vHl0R8aWLNxkjv3jW/lwNyIz819cJQJpB+qEibOGUZ00T9caz
WYXKLex0ZFvv6OmFhRbsc5v8zGc/ABENhwfXVyJOciS7OpfPYY4GolHMX6yC57iB
YacNaElHDIA+/yBbrpcQlZ1UB19iPoHHa6Hfq0bP0e9uLSXeS8PLpFFZRNqF1gik
Zy/2nrZs9LbTLHYPygwnr/DepXRz7xn9jJuxKRWE5VeaI/2qfAm3/ph+Yn8zXo6h
as9dvZIArFTu5+wZSV/ftjLN1BFDVaiqCA8d/n5KVUninHUcjAvtmuciBCyDlYI2
J3c5BkmajFIdUaqPGguH3XTVAPp3RNZrmc2p2l9UDKfdjFALf/rVOq4lxvyIi9BB
wk5/ZR2Gk4HzwNahclEcPbtU5sYOcw5kzfWCLxBD7y54vlrGawjAd2XycUJrZQ4y
PPWsZiSEdg7oc+omsEDHiO/yQ+FUigYom+fJD+/9bt0xEXe/Q3DuYr2WQ6iP1xhs
kLXnNDlyY5KeVVvPPzRhVC0/jNBhcMyqRtBRYrOH6lBeggAvcpLmCv8M2dapLK77
gQ2Fk2RUE/Ex1Iu+3l70tbMkpJzkNjkcq5MdSWkYcnnRB0Se47kqjpNSbUd0TAsy
b4ax/KyPIgGNoNKMOy5qHoDHCcO4s41um5x1k0mgE2LMOPoSBFA2Hl0dTQ61s5Pi
1Th37eKvrxc1om8hSiTVQMesJMSWbuhcZSmVxYuCoPcJXeo0bEeuVNGYYvNMFO3v
1ncLwAs6D/7mkTQfNIOQDyLdEtdtfXZso46J2bSJUuN948spRYz5SYokDi42f3H1
6ExafJa6hw94gtfPBHybCL4EhmKgos/wYOjk0sRebwkM/LopsnP+YWtNpe9mQsqk
CONBsffoicsFp3M2RgqL3JCsaSWf8wu+ZV0TH1/s8BHyHazDrgXAuhrhtYbezZpo
V024Y5BrU6Go+zmzUTj1atOyo5eUn1TsvTY60RZjbyGucnbqx9Wur12xtVKZHfv/
MMyZG4DcMFTApNBihFrbUTD1B/+1k6HKxDXUHTDEoVrC22jsxI+IW13FOUDw2Oih
X6VyVguLZUmMtUZmD8ULd97lgr8MGyeU1x9qF7LB2Iqd0OKqnfe27pn40OtpFgHl
ufsXo5UE4twDmlXk2KYCzxhBLT7hqRGuOlDHbBxGbmGOFBUS+u2uoPjiZGDyHmZ+
85++Vp7RT0UMLfE3qTLnxf8w6QS6qg4ERPfzMBJDLBlo16QucBdw889ij4mzSmjZ
ROeNd5nIYtsOmCiNw7hAFCHtkmeKQBxkgNFGz8B3Nyw3LbVhUOZRH0uEsyPDH9NW
O25uB2I1BShkHhp7IgZpP9D83lC7vM2cSZzkncYrAlv21VoYsbQQoam5jLhClxEI
7e4q2wosKVTuhtBy+9RDMILoLCCVkEfx/OmNU5BJ1kfxJu62arQEAtlFrXFaXX5z
uxZ/sGXDJG4obbYwtePQ6SDfTCEfx9C75gYMnZjqYIJr3e2Ug5rT5ZYptNtVrMLF
Z+PuDbTFWEWdlmHESd4CAJRe0AGd5ViXruOHK/8yyTn4qRTN3dA/SK630ON4da6W
K6AmjYdSVdfpdnoshsdCVCKwkOSgM2+DjzQjAJQynSTKZOrfK5VxHRu1ALq1f2Q0
AlolvnWjgv+wFuqCaU5YygnfkJIfsOD8rBZ8E/BC5kiiqilJoRGp+XVF8mcCGgMI
gJdVIodZLfw9cLpUk0iMWh6YZPBdhJrPbAsH3RbikzYQZUkox7MrwEqHdB59bicU
XjJ6Mncdtjw4PPRI2d7UHL1tROGic9j+VMwOwwBwVGFU6FvV38FDmfLt7hYgEC5y
CMV/wyJ+ftrfTEwe+Smx4/HhBfg6U61vrT1SQyRrQjO3r3lBZR7AEGJnS0tc3ELS
T3yNDWdk3PmCThIh/YH44q93Ws5omtYX4ebrrJjPn/OhaSpHfiLUkpwr8VqsumEb
XjdshUaQ0WVV0A4dVD8H8+s3Hxshm6aMUc7bXVZmC5VXDV7HLRv5Ehwbvfg+iCYY
I8Pw8qx+BxzSXL8fVIbDmzFS1blRprfak2qevRFZOOX11Op3jqJQrK5ubk4YrRwV
ROEe81+O6/nXvazn8fdrHtJN/mO/vWUqZjsYMCGwmb3akAMMtUwVeXN1YYkP2WDY
KYxCsynO76MdiC6wmMFI77kSqnRTuZAjLuddsS4elRQzs36v3WiY2pEzjbh2x1yI
6MA15phF3E8aznfX+jpZRzPdOw9zGju3oyLZslvC+gQSQcH6UrbP47WoMAykaSiY
NDFKBgxXZi1UAmYdYOb3W2l8WZz7DGcNOylQxAFdtzsXN8cQA5yGzEJfUnuFKNsn
pb5Y/c2/gQbM4nbvaanipDjZ2HR32MW3Fbo/KwuUqN3Vko5hb0I0Ub/PGZgZpJUa
E/hLYRIcQIS+tR7sReMfsNxwh7mHcG2KiShdraks3l1f9XSmjcT0azvysNAkc8Vn
fo2/CVFqN1noXz9zFtEERDWspeGmGwDgOQ/LF3AOzmhkENaknHfhBqolG9CNXai0
HtM7rKiY6HL1WxdmowfMKIlFjqMVuggr+P5L6hY+EnFkP+ezm6dhtnx67hhLn2pu
p4ugdzKlR9R/sl8lo/nOvJRbosJUHR0EhLMbXxgURUY/fZKKWbVcnL1z06pCZNgq
v/qjBOqeXX0iY0Zw6RIOz7Wmh5jhfajGOe0ssC4dQ0uEcezsFy0W5Hg6txW0ub0z
RoJzuCh9VyJG9nngZM0SY9HdoJwj+fvhgILuGBWjnFqVOyg+RouPb60yZLqLubhG
mp90dAEYIszJIf2HCWY5ehyY9b8AkiHb8YCYzRXk8tyKji4/YVaOzZ1IFMDdB2/A
rVg59ueEBrRBvpHhFemW8YcBo1bYS7HwMdK7pYhdKz9wLDxIOmQLigoBwIS+FqGY
QJp3xoIRQbR5YfVaz2+FAN9d0yk/RcfW9Xf/fzdqBmC5dt/i0k4fCu1fCgC214TT
heE76Pa0oJD5JXS4hOopwmYHssBbr92xeozNzBgK1rD88/P2fGOsppiAEJqbesPD
UVLe5DKq1PK6XOxy2JhOR9p7bU4MR2glrZaHUg1tlyGh/Y847ZWmA7gpvmWsK3RE
8cUceegvthM+H16r6DTlcg2mmTD9GyFxDrmK7wdkz9/2k6ZPPKHjE+cxXTW3PMXh
HJNOFYoPtPC+gQTzwr0cnrPMgoAttpc+iZYianfh2m97Ybpej8kmuFbVqCzvWESb
ULgMc5f9573ucpQ7dfhOrHHz2aVhGtETd5UXkKX2L0PeaO2nHMYBm3QMj3/Cyr2R
i6MXjQS3y4o4ngxF0aDIehwZk/kHwQ1y9co8+WlJ52JSWM8xk2oozzV3BoVscOCv
rLhgBF5LnAwydhXkKcspRI+V4LJnEKkhrBAiA+snlH30BxVqWqFCBPe7frpmZd1H
R99yH5nhA/Oz1uvUHhdC7UBl+ZLmwLpctPFLGTrKz1DkuuM8hmzs9dGTuOEDp0HV
szrJVEK6DDvl0Lk8AI6WQPq1S69O8OwMBj/ixo8TzhCZ9etQQJhXm52OA/at4HL7
VwZnEXcSf0N9GH9a/87nNjJD60hkTdbQuYLS5bNN9VMNZjz9Xtuf7h1YguuVzitX
sZ/6unDCBVDXtNKUZ8CVvd4bwjI9i0tUe64ClEcxy2MlaUXdS6ZbSMW3KbGY3Qwf
hp1A3MhiTYeCsIF9g+k/5i6GXQMPprP99+GV0jAHCUxxOp4q6o347YIf+xyKIzXn
SwuKwwk2TMSrCscfEIOHQ1xfT6T1gRJALxdv+eoLqwtOt74Nz4mPnfeujuVfASDP
JNCeN0ksuLQSLTap0iLIaCFuphjp8IZHFPaqIfjtE+h/PBttfU6MHywymdlxSwpv
BSpg9BL4FdJgEgCL48C4MG36Vlbr2Lu8j2iRyqXesSUT+pF/ygvANasKfiKUa/u6
MGaTHRJPIFyYCqlelJ7nsOO975EYIuprmlYJ5uXZojmfQKAh/7B4g9n7nHyrgN63
qbmupzZWdrLcKheHp9y2iPrrGdDjDp3UGmMag5CZLld+T+uwbYgm7VVVgUDX2l5k
M8K5Gs2CSrZbUcRYNCRhDEMYF+DXlLeovW5uhftEf8yYTOKFRibqawd8znY1Nx3D
xwCKrW35nZGJ3r9YKPsVlaYi/SaUPXkXN55qY5aijkXUX1YZMaY++5S7XXAIigyI
eEYSMvXgp80sQygICnMwsZ9VZxPZZr88Q4voDZZFns4/NoFb7eeptIXDDhH3KMqX
RG0nwMO7U8bdzdpd8/EUm4a+dQo/ktvxcmHSRRoYWRgiPcd5s4QEC5CoGvbjo3Cf
Aqzi8fOpPkvBkdv9nV0BKJoX0fSPBiSPMH1hF2pju323BAEvGX1iM/iCK2RBYa/z
+lW2cjUYIEX7DSLBLLUirTlwZGobMByyypdRpnr9rE9nRgtkA5MPgS+hQZ0Pk3p5
wOXnEykIwVI82nZmAJR0csnhBHmUdV9ocTqD2jWi4hKlulxY1z8Sb3UASqJTrsz4
vI1HKUTjD8Y5PT7eCPwTaYSvBJ3EcFmbJPUWYsm5RvMnsFtJU2dYlWzVXXHYHg+S
lyNLr2vpg8QgZNTqySvhG9nnVVzJc5Z+/gaKNuTNgVHlufPX6d1ZvYoup32BqVXM
8dPOmOuXYt+wjyfC67iC3SiL4wCSgtmlWJltNks6PXFuzvT8fhLyAIR7W4swaSNH
c/13MqIEJzC60qsf4tp/cINJCUpKAaA5bsyBG45sPde9HFL5suD5vE1ZXu5twbU7
ats4cWZ0Uow6yt/vUVGB53Swx9swMrw9frJIFv8VzfWL0F+K82J++Pm5Af2K65kI
UEQDGkuQA8kATbZW59KAA/Tss/zyw4POIRBrArRSevIkbYLmlwevK3/ztUIu0pFn
jd/bG7tpurOkjPOAxUB1bRtey3Yy6F//yFYrnl/el8/JjJPJTQahrFXx5mKy5eOn
UFvch+OOYrob3gsTkii/727WJ7pMdKv5CYa54rCCexOtyfk6oTOFEsAh7i1UXikc
k9lJ/tZYH8uH4Q3PRHzX34EXdopl9hDhyuP/S9PeLts6j74x3N5nMaAxl1+ZolVZ
iYHnG5i1tk8dq5OPKA7pKDCwoODZOH6XtI7m5x2Vj7pJbnvQI/F4dy7EihY3Ylus
h6qlm4wxlHGe/aW9o37h3SYDooKuz0qoyt6rjv5Nxlgi7k1Uw5rWdto16xqR3EdS
WhycMFNffS25D9AywNSUg9WIr/9u5/tiigeoOVSHVnzvjTekkbg/RXFjlGcXMP/0
ipxB0fmnzaxqCwpU+dRtLqF1srj4989kk8QgB9T9gaaVDZByFcoI3uq7Kp19y4mT
kqArf2ZEqJijpsvt4pp7WdLF0mjniOUjWE85wNwMfZE7NGNzF4SQpDnlzxeJ3NUl
K1ldGPD9zB/plWnaYGU/EIG8TJc6g1vYjScARN4/adT4EegQUgIj607PW1nRypvR
wOqcFyngrGfF4vKhf6N4glhUP8BuTvFKFW3yKOvaycd8IM6ZZ4DKss9DSfaamUPY
c94Cl4ZYkReHZQYjpZmfmu4i4lFzMgFXMErQ2SFuh6B2IQr0EORkg0239erZTdUG
QEjl8eHtVf1e+CeOdLI4ZDCllchdAwnaOICAi+ngnv8YJ47ssA2zG89CYD0zni/j
YOz8p5CzPZc88Ap6r4jRtl7fjH0h2QRwx0CPfEMrEtAiOUzUnH79C7xcfSZ3uZ91
VD2soUaxzEoqOlK9oWlFtZotq8sOO8gEyF/bLugf4hxQ1Q/lTSEkjixUic0iefiv
FR+H6Ouas+kzdO8ebBJqCRNi/aOsXDgZIt+Vohobxkz5rIi48yfXjFM9yckZLzOj
6mUZ89bmDluhqWjTDNa/iZAJkzRRFoHmfnpI5bC+o83moEEwQp+hMzxZl7BNey4B
tsr1w4OCzPWQDq+gBBXGmjNlULZXZ/0bR9x/JWBuCC5cIhMpc18FqbBfiyEKxL38
gJJFg36Ytghqtp4P1P8XSM4E4r2V4uGDyaI6tVXyLiJNkO5rFO53WO+ONLcIKhCz
DTqe4ZJGUERlMXBv5OFMTLH6e/RjYrAgfWeZrIRAkSSKrDYwF1L+pEHytKO8wJqH
al8uQt9OYFghBTFcjPAmFM5L9pzct07vz1xPU/Ml7b3QU4ZgMDeW1lA2aFI6lnJ8
saNgiBKvDXB7Or8N61u+8YemTMdfZPGD0jbLW9dOXxE3hO5z506guIbKSSjFGPaH
6ciWgzv5ZHtML58L+v+HDnfXxKCMxP7wvkCI5122QDMo796VAI7nVRgkUWcuYSjZ
7zv4MlQq518kUmBND113j372+SgD6L/DVUcUbHgwkU4aPg9Y/YhRKh2twN7In7g/
4Sa0D1uDXo9ijzbYzJLjFfJXbw/mmug2io8CRqGHLtyDsyGtScvhaMRPokMeTzSV
2h9TnJQiuslChnxR2cEveAip9PGE1eeR3DS4ZV5FQFklpKry/yU+vmc1E4ybOn9b
4SgN3Xw7Mtj3/VIOxJiU48B3MqwY5tcj3/EmZcVEW4dykJUh0Lm2Y8+/WgsGbJ7T
vuJ4SN7nPOeb+Ba3iYGjA2qATGvn3UH5O0lRLHDVXnacFIfxWkdvbAAZenh6XQcF
CB8WWMh+h11GojIjzfqzE+1GpF+9QXyiqc3eZjGCVUXlhgaPzM5Gbg/ONK9sZ+NF
SegtppmsuDMAhIfrHIprV9q4NO5UM/7SIgXqr3Mxs05kgQ/39TrBrpderQ8dpMoO
7I13ajDyxiqjxeaLeRFRup28RSU2iMitbDtmjjtqlbIKsJAXN+WeFxE9C8hF3mo9
siJLNB2rW3Hbd9WqZraUtFw7x9HdHuGdjaoVsECu6hp7AjMujb0VIJuaNiD6AVwD
pSisrqAk7C7S14n83jBDRIA0vhz1exFnO+8pnv6NBsW0Kcdh1cSQY/reDuAN4dcQ
JaiRWKb075vjJncjSV0g5ZKzh1zt/JE6Fr1oQGv7Ij3AjvhMNNEnvRfThGges047
WHrM7KVlbY/4/jeIQg5aLK3Cu4QBJZqVzY4EJjk8x6j+V/Pf+vONA2EvaTF42yqz
/xvBs1I6pUX9ibmeF5QpNUaDJBIzY2kaaOmNVFzGm4LoSecCPmNGPBzIAdxFDG3C
BrkqltPpljtoY0f2veihfSCFeu0qTFtd5RfTyX9IlAo1HkPQj9ONnxquAnOWeIma
VzuHiB3g5OEldXhvFsgobQqWvT25WISQobdhjPar7joLliPNqWPEKoHaAAdjBV4L
Eh+GHtJVGxrz9baEfDwCUt6fbA7toW/CVsLdDQhORUIouljy+ECbqbFU/wbWEQSJ
o+MsdkgupyOPAtP5XWApqm5/asM3LGYsESPtDIIr234xJoZPbZ8B6bXlNUCXwwMc
dd5H4ghLTgzzDIaal3dTZ0w59R4Y3WInAysmvKmhOi6Ql63QI3la7ppcXX6krFof
4nFSzTZ4Ur5/p4xaIOyQAr31RzHuZkdbqFF3ibKY5QmlZisQ4VvtI3i6ajEWMO/+
Sg8GEesvcY903uzn0PO514SQKoiXwmuhSjLCBusTNvt6gY2rawmVnASPC1xVUjeh
B11JqTJFxcQmltf2ELbMAfO0zOZsfWWi5+g5jSlQ/H8pBRdVTFZmdJAVOalyquFE
TU96ESe+8ylYOBfR/E2cIbseRGgu0tOwfhH7hBZSarBSPDUkoulc1jlYR7WLpXpL
wm4wRnm/SBBeSK5v2isQmuklsEHA0xnoJW4GCqxEGjIWgCx0nKqMy8KYejtaeLVD
M+f9nccRzow72ecRVmYJsjQfBlGmsE67810NrFzD4G+FpRcK1K0CG31+iJg1pCt0
rWTcSsqB1oBZqB3q4CIfrOF0tqB34OvQxbxxZH9Waxtm2oZflngsVJPfifLzry8L
CR4Dh3ezVLvaEG+o+SpJls/JmYSmjxiIVtGZP2viSMpJMXrOUuAqzBLuKC3cv/Mi
mAxtYIDOVM0xryFD9UAHV+WMh3f5NS4Tlahc6oU40cxD8MKgTV4R15MWqqeAoCio
K1/UybajEu7Z4Ovxb6FRk5rDn+aKnRqWkchEW5c93sIHoEyprAt4x67yhoK0Z3CI
aaC7PidzAeumucil/9wljtswANmrjBhlT+atOWu1pItFzCTjaUsExM2WKQ2nN4yx
4o7WXqdxFLTY9b8APgkbLiGF4Zo640phupj/FL/vHkXbtGw+4l0pnkRO6g/ooDKf
WeZ6HKollI+5wQZXxTInY+T/IrTmyotkxbA8EJB9zhtzbXHDGbAPehb55eI1ULmV
EgIQdASnIZ5vHjRSe6bIT3FPqmzD4nKfhtl8s47XZnDEO3l5MxcxKk3bR5sJvkbq
ipyINJUVhepB3HNCYjWxc45+c21Ps1eDFbx+pzXMou/ibLM0GwEcmiGkYx+y+8js
LvAvCyWTEFZiuKFg/lqqnCyCJVt89Z653tRjzJMZLxNw59iaWUOQ5DpxhJIjVn3g
uX/Mj9h6JWRvDtNx9G+++8A6KqVBB9CbczbtD6kMK6SWy/UvpldCWBTTN7MdfAv2
FTt1yq9Ehdw6Y1KOj0yKCk+7G5os+6d5XRGIrki7cc1ohoaBbferJkAb6gDRCYAb
hVdZHuOuEnHPGntA23zrP4TZdr1+Q6DLzeygCtR+zmlbcPRjz1EfFJH1gfK7Gbt1
7WTfGJaoVbJEEgQAX98zP2Nlyn9oHycaXyBo4XMpqthjgIeh7SXM62CoIZYjOUgr
0SYs1nVPzdkWUteOD682dWfc6XIvOdaXmiJfRi3wNwgdpLiklbyY5u+njOe6d+il
Pwt3Qq07e9kUE2t1yQQw8wSIVy3Ec1TLxc5LkMX0MJcBTX6gvALNalevOMAUK2rz
YbNisJYTTfULSjtdM//ZgBtlkKqPuX9Foqd6IUmxrNRB6t4KYCMza27K/gKSVZ9q
YMqzZx7r52HRJnUccEsCEFRBuZoxM/wpeY4AgB5AZb8TOZFEOqIeoLw92M+tCm0k
1lYC2J/zFL/sOP6pjyV3ccXVKsrsYyNVkQV9Y1/3ZuoskQfipzxNlkqIu2GlrPNq
yT+cO7AS4MOweRy2cNyEFvxWmhfdxPa+D5o7VOSosblI/yomHzE+ithpPo87mznk
/f5RBo4dWVDXIkUTet6XeGImwlDfmLHYazawlE6QTZn2MPBI8LCC1yJAyztAmur+
dPN/zUN+FVOTBJP2EztvQ46GoAN81UmvuTKbX9M2owMsRV31JBdmg45UUifastZW
tQp6iVdwJrOo3H89pm6nU4AedH23cullq3t8aRgoABAOI+O2xPHou0YHerFii5nQ
U5WNp3saVl8/H2Sv2pIQ1wEOpUdA3EDuQZVnbk+XyqV2YsIIPrFt23gE3KTDWjo/
NwvBrzPM/yBj08AINP/OVZgnJUqTFMtbvjcE8Fv61Puy8seS91qaNs4R68xfqOAn
bCGNcebDXjEd+RLzMGu7nKOSWMIjTp8ecmLTv/mNdHPQyL0lFbf2FgxzLGvOqg1c
Jp/xg91WTX6RCb/GeYSRcKGm/MX/kPoNrdA7Gt3yUe5wEhZLa3+R/aNhnl3fzQ4y
Qrw6evEDPo+cEzdhgC1QpcJLnGGdFuljw2rSwNeJ9Z7Fw/8aosz85hH/Eqe6fpPW
W2YMS7f3pIeE+fV2CHccSNXVL7CvOnHwhfEHowU9QdkvQCWJJsJUuOvGcjLdKs6m
RmQJQ8Fq3smSwPCEhiTADIyZZLJ/HaMukR3CogTib+BlgMDqTZ6JzvElxowTggHY
kWBvJd3E/5SJ2Odg0vT1czSAURZ+0jWDdv3HV88nPIICWlN5WhVQuYDy835QtufC
HBNUFcLBUY030PKH3jMoNhEiO9yJZtk2gn7YcdINBjgZv24a3hVO10ECGSk/2FkJ
zhz2XYq5HCW81yLR7AS/LkP06Ov/kUoC2sEUIU5XkRiMndPeqO23WGnOUvnSPYAd
QLpNAeSfyL2d0icvdXeOLmteJ2uPBkRGz9cTvJ0TirGcI4HsHwJL1xVYvW82Z6Gf
+JQQoM+SD9ZiLTCCZXLo0WOu4RChxCxxAJGC88wd9odXSqEJ6f482zWCnxWRu5DV
vVKPsrONorQMSMlImZnf5cxUy1mgB9qnLVESMg9LGG5fPf/eac8RYsBJV3XeWLmN
YAZwey73fifXsNv2b+JJ9AU/PdFNSID4SuaPuNp2MM00m16/xEqVqm0jWGCn/1gb
DNdC/uMUypd4xVO+E8+ukT+ERsjvNyEH/zm68M9LOC3OASsqEXonPXEp+W7iNDEk
j3Y1u8cmDbhCt7CRT0hQXGTFUQn1CC7IvpeDQPpxgeaGjQ36xSx42aBbdcsoZxr6
cGxszpQcjmJbjvTqVROFhwRFkLCCGmBD3LA2CunDXxeattqrZznzAXOk9VoRslWm
YIy9G7JYCugE2Yv9CJ4aEAVx46k/NQJDf1j+sQD+0vSR1+9JwlUvkMHiTIGoEcmd
vrNw3tcgC6bmzpF/Ein1ILCMNri5XMC+zRIb7r2Ufjkl1C/d4y95natzGBL9Eph9
B7IONkBFxJxWsqEQjPdcyo+2is88BXBIRUnDbe2H8ICHiwYiW/ZDz2t0tETlBasL
2g6RZ+5wHTqvT88lnm3mE0bPpnroAgl2UOFp7kJr0mNil653ZUABT1MHZFZNAh39
kmA6RCcPWTiMAfdohBSRUQq53WhDqfWfnrgnyv/CmBfLb5NMG8BWu5dVgin8KVS0
dXm/2wF1iHH+WEcmw9dJUfb2MzfvXGGcmLVA9uiP4KU3xMIiALYDsZy0VUWbzpDR
pB2xN9wxkdEgZTfx7dq4xNeSBSN0lq+bl18aNF2lmmCURQ6ieILsZfWNVXaU238V
WcJ46EBQaLI1Ffnrjs/L5NcL5tiUR7XUi4eV9nxXDxCnQ+QiyFcETB+4C63qzMZp
IjRpk2dIO+o8hgvRoN3uoeC+yPrMo3w2ZrZ+51g3Du7YG8YdO97xUyhU/4pN8yt/
EMkhNGc+AQ6I2X+uW1/DkvVFcfy5/CoqPWPi59Toc3ThS/37IuSpjYHkwS5nQY8K
QdUlGsLCpP9hllY4syqjD5NwA9reVld3qkaAGoy2HllunmUK3xZoig6wA9KUwuc0
GYo7PuqxZ2FBiz0ahh9B0xAARzlCk9D09MisagUVF91XEC2Q/dv23oMILI8b6fnq
FGJrqWq+OltyuecfukTySad5OciZEvvQZHexxQIlcqre5yGNqlin/yDUq3DiHIvu
Us+txzdPbn4UlAqmAX3Vpi4/Za5rKl5wr+2rz8Ky2iS/lNPHz7Y3utyRLSZTwvnl
/sDJpM6R55oLby105ZSHNmI0UdIP6RVlp5oNSdakOQqiAJMChwlesCW51alf/byb
ji5dFAEhyQN4XuxYL776zDcwM05fb8LKe817qEEcUn9HEQML8PvKdUHcsVCZKi6i
HgMyvEUVBfKj9w/YmwFm7Db6J/dmQNBkcQiROdC3IX0PuOQd2ybFY+XPGD7ocN69
FTxzzCN/CV8SL8GpgLGMSAq93p589RFXab5YX5+rf5zJ4kyj8Oak2FO0Zmo+3zOC
nep61x0b+TiccDsdO4H77QLv/TFJgXD58bHJp0RaLnPaRX1a+S0HhgIVMLLyvPLZ
ZEkSjG8rLnWr1U+1EyykdNdyE/m4j/VOIA1TioL2MNInKbznspSRXC2cn3bFn2b5
v5PGRHM7PsXyxS6xugf2TiVAipmpKy8ofwtIg34rP4qaGSYVrzrpXBu2YtKvPjLh
M2KJbH/Sf4RxIqydAn6EiEonXYcEN5O+ysMtK98p82zwfpujTiwVXfkgI3rDj7eM
KVhLtd/pjZqujbVaNpF/HyVs6uMk9cdDFr7UW1dZtYum1vR9yX0zRZFpVIWXRmY5
YT93rkYz1A++JijolHFCnYw/EK4iHBG1tkEosnnBke6C3QHcezZltt+oy/LXuaHo
F/MCGVWivtCFGsvYP8m+GFi6gKutm9W0u2APevSInT3UNqUE4f89ck+4kzTP2f4F
X/qvQzy6uWi4864wMal8wz7fp0wHsumwz+atdZwJVGqGGm18BqWmYJwbGNS+fvCF
6Ko8Ikz5hlw/HZzfmIxKsYGWkUzu03jWhnpGo1n2zPj3gNuGIsqFm0tTVlfwcywj
slhDR/SvUpK9n9kP+u8N7eU7Jxmby8ODi5ScqabG67vAdLOffO/whYmClkpHflX/
sXSFV17bU3wWUnDrsu7dcnF7s/I6MOWT//JK/XxYoTO+q6heZxH+C/GKaIzO7U3U
QvHj1vcYFdaVhZu55qYCAhLp6ibFI3FMQ8jJN18pIHTCdtcwjoMlc51PLChfvpxd
6rGGFfyrZB7V1a8TUewcziNb7IgHHCTu08B7f8GjZGH01yjOtL34DuOfvgDFgfDu
6gSuKk03/49VINEwaIVbd7VtmFo/mcjMPPXS1V1KFkuvM9oXgQK24l7YZiywWP/5
fY9xSicX+0A9r4W6TFdv97TLbXLUig98SUrX62turZyN1WRh6VKJHzufX8mWo4nN
SxciWuYwRixMe7bOzfLqxAcM4bojzQtq3gpIgbQHVLu57DI29lf+0t5OeZY/65Cw
XECQ2MmjqXv3JnKrDvaPRUQHTDK4kBywACCDVHJckhoihEW+LZxRTh773/k2xcx8
9obO0TlHxYzNpmBqUEpNt1aU1IwQfOEMLxj71YVsnn4QDRX3HxuPtSf8hjWCGgsY
R7Mau2aCU0Ho8AxyhlRSLTbOJ1x0rmw5gO7Kl1uAK5ZMf9imTTnNTUdEOO1nC3ur
mO89U+uBhVyWTJlAOMPkCYbsG5lsdhy7gsmhEMqLrMv43WtpLQh3AwqWNpNkWT/b
yzkRmaalcjEa/viWZb5E0jUa2YcIXNhLuI9GYT1ElEfnGWu/BIELgTQBBR3mIdx6
5FmrjdLm+AhlPLO/whoM6qLRm0UT69Xlz6E3ti1+uhoIWUEU03ttoQknPkwEBhiO
GTJ/MqCBPrtxGEGGpctA1fZVNqSrZUti2omOg7WNKVkVWghnTuf7jfsDZlpUIFeG
lguA4AU4KmJD0uXN7AbEl5lorKESz4i+ergHwb9sTVIEZ7XseNOH8rFhnwwIx4Ul
n2iXsCjrx12qHPp9EUV486OyhqaEKMIAftXqEnFGpQM3eOwDh8eoHdXE818r5wWb
tQtl3fU+Rh+B87BC10rtNdJEWxBrLR/xmE4EN1fZUvDlqVAmpfcS4PNnnhA2Gk1x
KMAqp29NUfCvGTYZPAVMu1VEbVZbXlIG2YHYp+60YCN4AtwX7fYtNDEhGkqRKvwu
zisvS59mc6aslHTuqQHzR0Q7uLKBE2Mn7qAaEIOThC34ypzzeW48Zyi6v1hiEYSb
4Uv7TBgkkHnfBMqKKahsqzNGVoukjGNfo2FWhEddXopeVRGfKzbbVUp9meTCIS2D
kq7yY3ixs6ORBBwKR/XUvDTuZjdOZ9bkFrJZV1+J6MB8qamDg6cwrsqwCP0agQjy
ZrtEQpcbD0ELTEoE6c9YFMeZlqD6jccYC84RaJjNmYDC530nlCJK0etW75bC5+11
XOPpIET2GaegMJSuVy6+6ExOPZXK73kLHqtcRm1pbOnkB9ihPpoMMR8XgbCC9Oq3
14fzKyWDPyzz80BWPZ8E18l1zffSIIO+y/2f2zJwqWeu1ZdYT6yimXAL+9MJ9or5
y8mxMhdybTDNkrh8rQw8WItg0jZzlIMwa+gHMtqmrZT1ztWLFchdQ0DcprSUsTQm
dH4v15n+ntpVaaw+rBB9XqOtIqwx2Fg6rqncw8ANHgcjF1iiYNxrPpyuoLjcv2Ge
TMiNZS0OAtnRcx8sFOgH10uaT7zObH3lrq29KpvRSe4c8upuKRpdZSjS/Wfn4lQ7
yxcx2XTpmgix9Yj/anVII8bbKyMj1sD7iCSTAS3Xd5ngStFWOUAIaN4NmDt2KIqP
G6YIDM0FwIipOkyF4vDgycxEgYjWnRfBFSy0LSswIEU6ziNytHwzvwD/lfMONhVs
44Boxc9f1113yYh80HGh5PNUxK+dRy32pnj7xu/Wxm3etTT04Z4/clzMF49W63n7
qPTSNMGOJ62lGhA6FM5MeB7mfZ6IKuyiVr7MLHcnkz3wVQrnJjIK3D7r4sdenope
O63UreiKPNWO8AhxLEo6xqsMoVqxdK7cnzQPWEUshkLffKNxAs5bj0RwONDG4ex+
T9KeBwEMG2kAf14NNTzafvSH5EOjxH/8tvS9tnU3FUDY6tVYIdSLxKbmO+ZYRTsl
tXR9Zq5fdaUsrEUE0yrseSutR2eCO2AUUcD4WVPvS1oX4GInr1yIGjLVTVIA/4z8
qmzdUbqdSWJGgYrpN8FO7e+DgeBjWGefQwq5TEK3iGaaK+9UBsAVPWcVmYJ+loZj
RQQWyVVF91J2msTHvqRuwPSeQDYl7N45wSHlIy+QvdMFEXWo+YB0hFM7eCach9EF
2+AHWob/hC+12Jt+8kZLQdnAPVBJFhcpsRPu4HttMtG8w/7ksQMOBIcDFqljBler
lLeV41wxzwGo1bPqTCc8JPi/PwntDhm/JOHJxrc8BlW2VPcsSQqfSqpWWYT37jZh
AqcZfXUKsW4eqLuk7cv1RNqwfbEczhohQ1wOaJx7HQHQCISHK93Go6GSx8NVTSKP
1GVZfTMkuNiA3M9zlwp5XqLWSrTpCkXS4CT0Z44SRdQDQW5GFIwrq9FTwLmXgJQ8
rPiVPm8vXw+F6zicqgFoZy99CsW9sYRalZPjx5lOkyG4ybhWUB5cRtLJq8wNb2/a
VeNlxMpOdfCWP7rh2Bg96vhA1dzt56xhDkXFVuxsyllgMuooqAQjclMQo3wMCbGj
EiQ5i6SpoCDZ6EiWE1uxe4rv2CBTJwLMcfRMdonOSN7Aei/9XcGRLxcbSwlI4mgc
knBHBUfOvCj1PPi8HNsvwVkDc6dFulqOHWEL3b9onhJ+w+HWFQCKyk/sS2o54x0A
Qfn6yTBu2oX8kLtNYL3swgu62/ozxxRslnQG8P89meyFTkstNVG/J5z4SKnEd4Ea
cRc07pK6LZTeT65hAWsPRQSAYwwoW/2Chz5fHOpKfln3bYz8NrDuv9s3KCgQvjbl
asLqtnUdYbwoVdKXbSxNRk/Ik1PRAjPCvwm6yjYknAlFR6qZV1fi2bo39X/D8c9t
t/wAfE3mAZsd7gre9/bZxXeFb/6AB1N5E9b4UfJpLwIT2klQHpVsErtofpROF/AW
zZ4Vb+4OqhIY82scu8WtvHV8WbhaXssYycE1tmlOHC/XOwifOU4hTUg36Cse346A
Ibhd3VSuLr1pioZ02EDtDTvxxw9UsdrQeBrXgrro53flVeSErhbRgPEMHotbdgrK
ugmj12STDVlGQM6eRH0i+xe+2cwXv7z54d+e8v3HFUnUzcOVBp+DYeyim5bNJ2+V
gTiUD9EZOWfnAB4QdCr9LHgoLJsjdTfvFkOpFbq109nk1yq/L6LNB0Zf/omuuebr
lQK8hjnvwz4mJ76EGZ31f7Sn1sanffMXpG+9f29xxvc36b9D9qNuQ67pJ/003fe5
bEKwjKX8Q6UioSPFYt3X7Ax6ce+6juIfhIxbhaqN7GPorIj8qa7a5FMbFVSOMUGt
lYeBARgY9HpYKLs/BzppfNerGdGqo/YrIBrmACsvZnuj/DLs9en5HxbM1mYiiO9k
y0F+DYThB0IeyJUJ1PGpAKUgMasZPJM8yQEAgbe+862mbNVnSemH+IaIOVCL4zGq
H19my2jZxkqiXJJZdCIxLwB/+nl5PMBXvk7DPE0Ofraah0mFEVTxTVXfFS/aCaKN
ogu4Wef2r2uZr6u++RRw2fjZJNjiLaY8vJQ+ndlZ8sjE+Ne2dRUTYBwkDDqgcD7e
VWSbne1omIx25ilO65TVyS6ADiWZ2dUtzpCjWU/oBox1CXbFm/1UKY9lXlMU9QZ8
1WOdmiG39WgvYJZwEvs7KxeUFFNW0+gslQ9qlPIHwTKdr3XREIl4aGbrdF/QiXkH
736pmj57SFeGTiMMLP2dT4lH0Bk5hKMnHHfhtjG8cwrT+hGaCLbTVLc6Ci4W78mF
rEJyCADdKPDL8juMWmEv1sNfan6qlM4ZJrlAHQN5JVfPL/arHafHinGNC+hzxdQ0
7AauMEwRFpXzKCEo57UpuOS6vwPPZugcOCtII7pBQR0Vd6DLG8yOIqqjBOFLHS98
/I/LnOU4MHQzeqf3MTkJ7Vcr4lsnzY5alYhx678z4+7HDNrdMq2h8XA4mC7a0+lA
pwfVIeOr00Ta0J0qDNeVDxTh64AQ6ZLjFwLvlttjyYBLBTUzQQCOOsqVCsRO7sbG
vAwZQohFA2q2GpkFhwCePH2oCTJ/yiIHJuESFCvLmysUrMcC9ovS8Oad8d/gte5Z
1zXY5bjymZnNYdXR0kVAHECao19+SX18x3k/3/exKH0bubkT6hHFO7/2WFcCBH5K
vTn+H7pq5Bt5Ku57RqZn2jMofN9gbh5qGtp5O2U85sDjNAZEnfylsxdDgHMxbK9P
BZHF91EsOkVfFiYnyJFBJ6THHbPH+VAXFWA6i7CS19Ref0bX0uNWjLV0UTFEjJ6h
oQI+YwkKpR/iHfaHgHwgM53+Zg31ilaFdZxt3Huamgsk+tK1lm4MvTVocZu/PO38
elMYjW5EsvaCqY5nAh/Ab/HlMAmAfxrFzmm5xuDpfoVJTywvu+ijfSBwJ8TwU/AT
dqnDiifenWMI5NzwA06jEevG9SS1aVLiTHZwAeAdUMCXLkg8OVUz9WrtM5AgBJAM
V+OQm0lq5W1w3kzkHNQ2QjJAfB45qRLUbGK8a1NSST8c/XgCr1Fdp/JBQJ1x/mw6
udiBVCOfS7B8MbE6fsKqNJM8TcOFj0YACKqFsNFb5JZIgJpOnlgq6JQfm6Hj8V3r
ONnenyf7Tahl+2Qgphjvfd8GnyShRzGluYdRARiqyP9o8SQzt6UXAj0VxCqlKr/e
uvoGe4O4CpzjpY3Hg7XTTpvcGWIpZhhWRVqdrPM9itF18Jsi3gCDK/awLU6W80am
81F155nvOEt5XYWWY1dkl11BlvfLHKfVaV6rTziDwvrgOelkDQ1Pg36+ZmaeprD2
fvhbrpwoL5Ye4CEKMfoZbolaSNh9joOR4JB0H+nPlW2R6wONToiGmFf3tRDAk4DG
JR2ra1kwUhDlk1zRzx0XzZYHh2RAWmoPkiD1OcollDTaG8/b8fIugeXdT0xIc9pl
doywd6Lf4N9+uVaBuAaXKjQaq/p8XBX9yxs4Qv9UEhQYfuH2ql4dTMOSxL5+saT3
uHMytJObTrcge4S6BCDdezCHSaoxQYsgUm/1HhKpHohEeqvzN5kmumxzz6IftLpw
xAwr5jlEulnt+InZipCnVNHZesLqqO0vYz3ltGfRQ6dmbIL37bWtzzkE59wfeyRP
KNTPrInEEiyxSEcy3y5Wha2hiWi+4v2x8lGOggZ/9QpUBh2FRrpv0O4/+h5UJVsU
SxCnRaSf+ljMNwVt7eV2pIe1CLLRnkZf6eR2+5IsUtymm7PxAzXYhcHb5K8XtriZ
gcA79D2vge3y+cDBIlAJXlEQcOJoab96nQYG3Vw0npiDbpYReOY9Cjdh6vIpS/D8
ZAvAnnaW3Bo9kRsE1OMCK//1/IY2sNQ0Tzi5kTVWE33F/zK78pt+kAUSADCyrcBZ
SkZAey1S8bP+I6zwMXYeq/SeY3/kcnoP8Tw0GxHXm38p4JrPgU+2K4yc/fxtrMz+
T9cgAf5i7g15JaSWJJ9ytPXZzmqHWuF4ReWkV882ECXaeIp8FSktc6z+1AYdeySZ
LIexcPgvABTAU6bgYu5sUrP8xVlNN8qpRobg6fc/d3WmsqKzgZiMYXG6Dz431wxl
kBh8U8lLQUGFEnCHsG3T2Am41Ry7jZIaLvlKDWuTavr7++fOideQTnCmWeCaNqN8
2PhMsIKoRFY3avscZti0CUAI1+fBBjaUv6YOAmlbibj/UOt9l9wlYzF5dogDhh10
1X+BaGLfjjL7K71MyPRgTmrC+kyYoLAORmiHzaeRgywZvRQdZAXZsOCj63+DnPbH
ABHR6ycW1++KtPVgol1wKCkTIWI5spmimTroMCPJJygcQk5bFl3Ixa+GEUqGfXP/
F2//ca5Q4Zs04c1CDiSs/vfbx57VMNKbr0l0zaXZZHdKkR36w0tpJX3txExktb9Z
nJw0UAwI7I5IDL8XzGe5ZagAYTlu+i2TjOzy8VELhTMyq81VSZ9frlGLkUYgSizX
jphL3eTUGYSUjWAGbIZ96V60M+/hbQX0I5mk9sHKNkrjwYR5TYcQj77Nj81Yctjr
4cnw2hO7S/ksArYGz2XbSi05rO8mc3XHxIgWssWVWv+iCXdtBQSuyAzFbq4Lp2CB
5kTt06EAOq1yOMigqRyw3P+6UlGqR5gmprXSNFEIV197NikV7yvcrIz8aZavcjq1
a359guZ1dD6ytB79gbxZnpQLuDWQwiqEl8+0qGvtLsiBSsjSGQbpHuBL8jPY/i/7
4s0+I3sLmK87/d209kaDzNdNAhodA6XN1iDrtk7Dpdg8+Zdd1wzTR05pjvJ9hBx3
UHZpljqkq3sNXMcGGBaqjfhlt9kWZcyYeZ/ssjLSLr1XOHAxIRw1OcDVN0vHgdND
ZjKqrO7ZIQsJrqDQsJqz8Cw2AG4oyKdE3gyO+DJA9LEf2jit11WuKlEiAhBczZMB
WM6/rkfC7WTvq1ho6D6jnCz/AQvllwW7gxluswfdJ8ZFfuOraHG7A/AucpKLhia9
00TC1ovNFAvdpcwQIe12tR9tR3EKfYecNAWmS4orq+BiIj71s0RKDrNAI8c5l+eH
v7YBpjcQUC01aBekV5sxynbODFtlk6Tkw+sS4mPhOtLqmajrG3parAAgzQ7T3xMW
1GCTSiQ6BHvPLI1VPrGkJtWV/LNH+PjApDalNZxZmjFlMJYDcO8yENAxBJnzVoqO
/ZKCy5zpg4u4NDGl2PMiIABStIjEX7RAKhnWiccACr5DhGsG5mSZwB0FF/mVERwW
arZGS7n7Ar28xlsdZ5npGs+fuO7smYyChcIg5IhW9iWTV/rGY5UskHfCXby67UhA
XursoViiOKdzfOOBaPX04LJAqwKYS5GaKsywLqNMDil4eOAGjPCLlxe/bPDlpX5v
QZmQ2LuzIrGYBPePnZKgEGVyLA2ZfLyst/95mXUSQ6KHHZcLz6PicTMval0nvGmU
S4veWa8KR3p5kCZ1bUmZTTVUWaFpwDToY0kH1+BH4396z0n/KUbjSECe3LS8DoWv
pwgdXCDZ3oFUsCXtcAXQZRJ0eHnqNo55QeTribJFIMb11hrh5cpQ8IJRDf9jWevU
S1jshFR8FkFhAKAzF/9uZ77FU15DJ6RwWG2kqE1nyVwofDp8sd+W6XL84yhspRXy
PRswa0AJmqrKa5IIaPKj9+WGCilbhSZBgKBJkX7HRRdaxZ9HF2K5ewTaNzsfIRA8
yt+ZIoj9A+khlcI/ZiHxxoZqXa7LM7YfHjEy7YlublR7RoV1VOQF9P/xjVR7hL9M
93RTd7LCBKuZxDW0c1NNKx/oojyeoxsLUwHiTCaDOl8Lmgr+2Wik9Hr3YTPFKAEE
Rs68Um6CBdtkfyzzjSr24oEGPU28e37krxcR32/+AUFVencGHbLoar6VujT/VSEz
C709MgtRbiCVJ/9xPkRTfiMQVfppUYMy5lT36ezOkV1+/M/FFPyL2zjmC7BCMDxr
dGdg+IFW4Vxz0xmckj1PWACd8y/p2oA1XZLT3ip/DHEr44Tf3nxQwu1nyiP0Sy+N
sR0IGD2TvEMRxf6tc2QuumfREnMUuUQ/xhL8X29Xp3p25FDGfwDl0jzYpcQot+3X
o3H8cyr8l6MmnML2zNIHs8jnRf0bDnlrwvrSMB9sRkwxQTb8c2AxCgtMRkgTijN9
ifB19a29kJXBTyKxPs0T+Qtyuu41WZ+AgqyAqA4xWbCJQ7G+Fqodlfl0bEr2wXK9
HmgoSuWW228QACN3eHsq6p5xe2BV2h7gYpoVQWkF3FesqUEWoYSfIF0r5T/HawDb
dhMJBp2iq9i/UBKihr1OPMqFPmtrMoPMmiwEMWf2j2wAr8ucfSpSaYUi94/TFwWX
pN0OP4N2v/gj+h3n+7MPhEfoN6cT45EhiFPV0UvoGR/UoWNAp+w+KmfmgE+Dn+tL
HVqKbp5JyZ5T+V8nZLaz87zjDOtxdHXlpjUYFiVhm0hZqwxhbwRqKrhZut/+oF4P
d7Qy41yRRjTugwEyCkk3N6c6ifg7uB80pj4xVsrkFYfzZ5S1tY4c+tXivd5nloic
84FNeNu5elZ6BXcxFkvnpF7evaIe4GhoDVqp82J+MaaUSqoD9MSS54ncohQ9YaJ9
mPdJctsqnkdM7nXNEa8t25iDR6oj7+0WIzifknOQ3Ui77fV9Rw6QfFP0xNhDEXGA
/1/v2TKmQLcKkfZ1wpSZTeXrWAiWExKhOyCSjXKDxwXrkvhNij8ss0sRKwzr5Dze
MJZ5+U8gKLCWqUIdUB6kblnaMS17GpGgkfXX9ZGQppaBqZsFr8TBVeOT4bmyS/tq
WrlYNWf0EeNuJ3pffTgmwZGrOPhvkPP3BcmzEwb1QvMoM/pvqXWx294uE6X2Omat
BZRgsTQMgelXbMy+ARDH1MHOZg5nCAlJUNan+KxEGEvPhvmxxfMQSJV8wv0it+tq
11IaadtAbjhid5ZkKlT3X/kDPRUwDNqbpaLWAApiEWvSscd5QULttzymgO0WHHCV
OORxYvoQji+On7sVYdoQGywTAu/uN6nTQbrKSgWZDKErPfW7+GY2RNjB1i96n/6E
Mc71JQbhHKpINAk1CjVTEi3YRXrnFFPLkFMgBdNRfhyE7vhZKxOn8GsrxVQrwCWO
21TVGMADsvfMrLuK9flnlw3B8kZ7RKIDptmqSny3e2TBsRMUEYrt/S5Pk5QAQZ2g
VICVU+O+eLuktLHn3jhclUFc67cqvhQ9JJKivKqpeLqBun7SvHN+WjKYr5AX0Sor
dEfKbeL98aNUPXG7ANByu4VyGm4tAk05R+0m+1pcP6rawwq30x4qypH8vaJN/GUW
FGjYFmAfgeIyi2q9bQruBu92br8R0uhMIhzx3BSx1ut681BNa7Vghz/Kide3/hGW
b+h1HF1x1G2VE/vNrqNrIE+U3i6meyJLufmsuhHgss6Ns/hpsxUtq13KB1DJDRtB
PqdF2q1Vz1MakX0FvtSo8oD9I2T4wnJ/bSiby5Ywaxj0ZuGTCJTJRv/DeiB2idFB
LtIxSM+zlY0ziHLX4eSI8A10noU9I1Z7G3LD/ItY8lmXuxxciJ6ZEk8zxgP+kRWN
WS63r2A3cIiwht8WKM8U/nMNa1zgropz1JOM+zVyjvnKqbVO1FELNCDw1kbmbsDZ
0qe8zZDYLBOzp80n04MlQMQSCkA6V7MCk93mGg9FHIQZwqTiygnn2N5yVGREkrWa
VgNhxr9YN4UvvWj0U1b+FXL/TueGaG2ial25dIBQ0V0uPcCDC8QHRbn+4xx7/Frn
g1kjmOoQFdXra89s++EiQ1InJxnr4UW8O7rmt8uc4P3KpH/eATO3G2IX8aL0fgyu
PjWg0GntvhY2ehBt1n8klzURKWF2TqrCMJjHMgN4c366yoT/x0Ft9ALAHQsl/d5+
CrBnuxD8DYXPeWRzHTArx3JCjHHSvyN3ovzxqy0wOEb1RYY5mufgs6J1lFACli+P
RXIdks0NniX2WD++MEcLd8j29X2WkPeLN9GkLjzdFO/19mlpZPdpwATK/+KzamDM
XMTjGA1/ta3qcTSJdE9EVt++/kH5xLP1QgSnFhUs/sy8p+6l2IBG6d+Yha6VMciG
jz7dLzrUAHSvE7I39BcYtj5BQqrFMNLRdaYSpsdshTP1s37l2xSDmTZBQH49PRpu
XShKQFloWRL5Ls9JJd3on2/VCXciLXOV80VCXHxH6SnQLLXeMWezyWGM2vDOEnQt
Ldh4YPa0dY/F6NnDIJFFNFMYgAiZFgOynGSDseP4Gtf6X8xCJbeCv8LVJfKH6iB9
wddVdVhPj52e3V7HGgosNjCJWb7ky+61c2Q14UKEKYIkIC8W1RPp7TlCUYhbMujS
vFtH413xQkW5cfw8/jzkoTqZr3iC+852g1ZIprYag7I3nSYLktz0VYGEreaZhA3/
RIbiDi5YNCs5NghCvh/QEo8fObG15rQJBPuRePmb8GhTNmQzFR2b0iL3tEzCv7wm
hOOouGIHM32KBFx1R444gRhiTf69XtWH6cLmE3s/9xQTtYGBaiVMvCOWEI8NETkP
Jr+xa3cRq6oJoYx7l7+Pa3ggTx7iA9uyKNA9pht+3PnYSP0vQZwhFNpA/ai4XBSo
4Nc5KUFzDnXMRI1fjGbHUW45gq52BjNWpnB5N+Nk/NEZgV10CiAJobNeLXakMC6A
aOfuSYHblYQ/a73zoj7Yvab2/22Y4G+xlk+a3NCo2ApZgJSFHDTaUNBKkxGLUkCM
noD2WBAq0qCGjRalEchJM3l4vMqOA7XxjJDZeXruFiBNbR8uwbZG8J/SbN1bEome
V0AQcyo+PfTlvDXYT2t21um5g4OMCdEFMrAp40hyMS3R6OYBfjEMhsM+2iDZhhMn
rxir7orVChZq3VGk5/7Iuz+gKJzOuuCY8zkkjtMOOBoDgXSOy+PZiuImFEs3k6M2
t/zevJbQZsC91OYlbjelm3j4HswRNLw9+m03rMLPJSY85VhyGpyYbtqMryKhBVM2
ahRLQgHuWdLP0t7PJsNzP2oJlKQCKW+8EMgmQzcYaTpFq5Z/VhimC9pU6qCi+c16
l0NWHc33Q5GXDsxPWKA6xkHExgKKNRP1TnwKmLXbb7rYgCFwZfi1/sV8VXnHRbub
tf9zx6/pAR46p0sqiNYhMcN/NjHH1E9Nk1cIkbItA5pSIct7BjcALMUbdI2NArt0
wRl/akx/EA1iIbEBzR4ehFdiBseEvRFcfj1f5wauII9TOk3tTGmf9wuLF+NJ+UOj
T8Sy3ueRSlyfC0/W6786Qh5HMkLJeyO/c61niK81r8awVPEU21E/SR4Z3g4UxmcZ
JjhpRiu+QE35dOawYZSenarV2S+Q4ffZzvet2ZROSn/psXfnr26gWWv5d2TGFRI7
O1uhdm1L0ILjWPxPUWiYad3diTHQ+wWnzFMzvjEAsBbxKegbN06X2vrJESxf/3TU
0DYn68JgWVRXNfvALR+zcdMW8BYfUIubOiyz41ryOy330RH6DevMqj/Y9Iymwlsp
Lb+duSf8hTZikzv9cVPiEHZVKfAby1FXKEr+vCgUfjnHEJYioXCc1HX71KvfuZoA
L6lEcA1PGYoPziSbq2lHvUX45t83GG64O3LQl9nWawRW+j5SxTo5AaZUc5Cexos+
6ssdiLg0FNi5SQ67YiB2rItX+933inWyxSsP84WYM+mGMwP9qYg+ycO3mL1g0LCG
U6x7Q12sEdeeMlMiuJFGJWe1ykm613B6mN7RHW5JXSij3uAn5+IwqPLx8rK+3jBk
l/Wp6pulBGEcxBpUhGAhUOJLBjqs69D66j2c3AMnYXU15HpTx+oUSJzw5GTdMyqQ
5noUlRWWfxupQ+T3ALCrpq9SiPkKK2HXX/YGAMU/8sjvWnF8dZIzY232/OXhdYtD
Z1o7gB2/jSPn3AjoaepLAWa6yEDKLv/8ofxCOnqPQWszPKE6VBFy6ZdpKbtcrS+I
f0p3Jufctjy4lmGd9uiDbExXHSoQusUHK5W/dVXYqWaN0jjHMj623XL8jflzgPks
hkprEyLSVKXOzLyaTwcpdHwNsA9h3nXXdz6avoclSvVWstsIBaHBiNFsfNNbO8lV
iKwRori+BNvsJkFfZLHaSKVKP6GIgAGTsLavId4W9E0jhhvYPL6H6bSPtk5sFB73
UFCbY2Zvfa3php005CPkd+wcKN6Lkhh8YMhXXdCeJY620lk/p6fTHukTv2KTNiRh
kkrhOZALaeXyg02zMoxNFhoVJJmkK2EmIsj5We49LEgKVvTpBVXCrPeHgpTMqHxD
tNFureL0rMSOSWChm6KgqIyCcO95ixYnLKmvPhGYDf1FMCCNNnzqerWAcKt2iKLh
Ezod1rUfDO7nwtsZzicL/EtfD2wma4ck1voY0aszI3z+bmiA3RGmlc3a1lgqPncJ
0m1bVLBpGWOXMb3A1rlysLjD6wMoO70eUyd1AXfv/Pqfu7dfZ0IGB+Xgu93a6DzS
1g+HXXxMirWe4VIRJIAdW7eZKxwVd1CeGCqYxBCLh2KS+SPrDUG/ZAbsotJiJAnr
mWcue0R4iZk21UgaDk4Ll9+KadKPMsylGnrE/+DsPLsGGnQc56g22dI+p9Tc6rlp
i2tUVfKtE6+dkIM45vG2pd8/O9Up52T7JtEYE8l3aLsxyuBFvVPbRNQZr7dLnhf7
YusSR9ljJSdlhhO2GjSlakl/s0gvH25fhDelO8TNloDFh+q1qaum9MwbQmzGtH1z
PFrRlzqHaf8N06hB6B0JdXGrZ+XC5u9nYI1aYzioMEIL2FYZVnnW9iNoBA3jlHfw
iTAY+foH1Wv8Lyo7RkVpokvdmXuiZjrnJhLwEh2YPlTsafUQX82TaCQ4PIqN+6TT
p9UpwHC4CjDp5BkJlGdm/bfBCwS10NCK8mdVI5oQbFu/D7DMWW3iIzfuMctq4f7R
q5gEi7NZAIZcW8+/L8PAK6/1XwzV8eMUSJtvr7/1CCUS/PGvf2h9ODqAnb3AJu0F
ckwas3vxuCFaD+VyohuU/i4Rd4Ad+KfZLL+bAcRltTMMdqhFyL1aeRbahoD1RFSt
7AJuPH1w+1eQiUSKYVR6Y9wGd5AQxW8DNcz50MheFHUv1BiqMPAHzuyulnjHkoKX
yti2FoiF50Le/wc0TPGiZ6TCZTQ3BlUBA/Ujofst7roPuTbOTyeXFoj5j5aqOIbQ
MXPRLrheufojA2vrdUxzUA==
//pragma protect end_data_block
//pragma protect digest_block
Q7+gK5a0PUyWyxz+JfRTwSlnEuM=
//pragma protect end_digest_block
//pragma protect end_protected


`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_slave_transaction", svt_axi_port_configuration port_cfg_handle = null);

`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_slave_transaction", svt_axi_port_configuration port_cfg_handle = null);

`else
 `svt_vmm_data_new(svt_axi_slave_transaction)
  extern function new (vmm_log log = null, svt_axi_port_configuration port_cfg_handle = null);
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
  `svt_data_member_begin(svt_axi_slave_transaction)
  `svt_data_member_end(svt_axi_slave_transaction)


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) Tests the validity of the configuration
   */
  extern function void pre_randomize ();

  //----------------------------------------------------------------------------
  /**
   * post_randomize. 
   * Calls super.
   */
  extern function void post_randomize ();

  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode (bit on_off);

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();

`ifdef SVT_UVM_TECHNOLOGY
  extern function bit do_compare(uvm_object rhs, uvm_comparer comparer);
`elsif SVT_OVM_TECHNOLOGY
  extern function bit do_compare(ovm_object rhs, ovm_comparer comparer);
`else

  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_axi_slave_transaction.
   */
  extern virtual function vmm_data do_allocate ();

  // ---------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare (vmm_data to, output string diff, input int kind = -1);

  //----------------------------------------------------------------------------
  /**                         
   * Returns the size (in bytes) required by the byte_pack operation.
   *
   * @param kind This int indicates the type of byte_size being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in a size calculation based on the
   * non-static fields. All other kind values result in a return value of 0.
   */
  extern virtual function int unsigned byte_size (int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset, based on the
   * requested byte_pack kind.
   *
   * @param bytes Buffer that will contain the packed bytes at the end of the operation.
   * @param offset Offset into bytes where the packing is to begin.
   * @param kind This int indicates the type of byte_pack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being packed and the return of an integer indicating the number of
   * packed bytes. All other kind values result in no change to the buffer contents, and a
   * return value of 0.
   */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset, based on
   * the requested byte_unpack kind.
   *
   * @param bytes Buffer containing the bytes to be unpacked.
   * @param offset Offset into bytes where the unpacking is to begin.
   * @param len Number of bytes to be unpacked.
   * @param kind This int indicates the type of byte_unpack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being unpacked and the return of an integer indicating the number of
   * unpacked bytes. All other kind values result in no change to the exception contents,
   * and a return value of 0.
   */
  extern virtual function int unsigned do_byte_unpack (const ref logic [7:0]
  bytes[], input int unsigned offset = 0, input int len = -1, input int kind = -1);

`endif // SVT_UVM_TECHNOLOGY

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>read</i> access to public data members of this class.
   */
  extern virtual function bit get_prop_val (string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val (string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
   * Does basic validation of the object contents.
   */
  extern virtual function bit do_is_valid (bit silent = 1, int kind = RELEVANT);
 
// ---------------------------------------------------------------------------
  /**
   * This method returns PA object which contains the PA header information for XML or FSDB.
   *
   * @param uid Optional string indicating the unique identification value for object. If not 
   * provided uses the 'get_uid()' method  to retrieve the value. 
   * @param typ Optional string indicating the 'type' of the object. If not provided
   * uses the type name for the class.
   * @param parent_uid Optional string indicating the UID of the object's parent. If not provided
   * the method assumes there is no parent.
   * @param channel Optional string indicating an object channel. If not provided
   * the method assumes there is no channel.
   *
   * @return The requested object block description.
   */
 extern virtual function svt_pa_object_data get_pa_obj_data(string uid = "", string typ = "", string parent_uid = "", string channel = "" );

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB.  The pattern is customized to contain only the fields necessary for
   * the application and tranaction type.
   * 
   * Note:
   * As a performance enhancement, property values in the pattern are pre-populated when
   * the pattern is created.  This allows the FSDB writer infrastructure to skip the
   * get_prop_val_via_pattern step.
   *
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
  extern virtual function svt_pattern allocate_xml_pattern();

 //---------------------------------------------------------------------------------
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+gUlNlPYTynZaAQk6dRXh5g14b/1p9BWF94jR80pFKQqyjYozBlccryBiRqs+lp3
3Iw9fsYWyZLwOJj7mHahgyd+GPFPQraUHG5Zu42G9TC1Va5COorI18HMXpLTkwcw
QGMw1yyoTCDyQabXM1wg+R/mEYHDbkDHhWN8fbuXRagxoav2Pae9rQ==
//pragma protect end_key_block
//pragma protect digest_block
ax/hT2ypBOqeDvDASp3XwlKYeuM=
//pragma protect end_digest_block
//pragma protect data_block
zeih9cydj+y2ASqXskvn3oxNzLw0iXwjgfUfOwZUkMFRXoOF00WuBLr8JjWfiKUx
4T0vHV7kwxWH3unpv1Hm869cM7XFXHNQdPlahoiZXNnrHR9F7c7lHbcu3oaWu6wd
S9W12Z38txCgop5pKShDteXKMuZvj41KWmCmSbhtofq1GP3moPb2/2HKJ5KAGkzL
oz7FkWlTTU4tES788Z6gZ+z2jCQIAP0JK+bUrdwpvMQ5qgrJWRZwwmxVHI/MbHYn
ITrYVjmOY5HdiyZUQ9DYuY7eVaicL3mEYyFrBb7aXDTrtSuvhxLVR9MO4CyDBSC8
KX5fEFuJL4Qi006F64Yq92jYHvVHNpxhw42h8befWe2+oXaE0CDxymNSsJpJQFBd

//pragma protect end_data_block
//pragma protect digest_block
VT+ljgME2GJOQwlY9GlKEPiZqY8=
//pragma protect end_digest_block
//pragma protect end_protected
  `ifdef SVT_VMM_TECHNOLOGY
    `vmm_class_factory(svt_axi_slave_transaction)      
  `endif  

endclass

`ifdef SVT_UVM_TECHNOLOGY
// Declare a sequence library for this transaction
// -----------------------------------------------------------------------------
`SVT_SEQUENCE_LIBRARY_DECL(svt_axi_slave_transaction)
`elsif SVT_OVM_TECHNOLOGY
// Declare a sequence library for this transaction
// -----------------------------------------------------------------------------
`SVT_SEQUENCE_LIBRARY_DECL(svt_axi_slave_transaction)
`endif

// =============================================================================
/**

Unitlity Methods for the svt_axi_slave_transaction class
*/

//vcs_vip_protect

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3eT6xcYqBLJKpuxDP261KIHkqQ6dPU3VBsm46vzqcixkGp0wSGT1rR90TqEwXZvs
0tNdoHfeNeUOQsA9VSEhB9tM4w2Alv4qrqUD6BB5R47eXLIXI+JGi3y+6WWpidsa
jcJ4JuuEl20z8yKwo+VeswjHS53oXNu+1wk1vYMr+sayAwykkYkTGQ==
//pragma protect end_key_block
//pragma protect digest_block
wBOCbwILWGcqdK+61WgeByfBagY=
//pragma protect end_digest_block
//pragma protect data_block
HlcsndmE5X8w/B0OcfKhUxo3GJibEyho2i/Y3gS3ZoeKdAI2I5cXJmg7bTiTT1Cn
JOY3FDyuoywP0lJD8C8WxdhzA5Emitw91otgwyHmYOZQngbplj31yyyxoKWTV/CN
TH1TRuIuxtaHNd+8w3hSee92w2kuVL4Nwvg8u+dAHEzgpXWvYeQ0YQZd5lBCXPkb
Gl1lI9MYWyS2TFJ6TdH5DuCPyOprETrxSQHSZySPFEeR8YkdSliTVdAhPMzdwWg1
cVcZBQgFVuPCQDInA3VTrWkjEZA60PpK57G/hpJQpJGrgUXtLuyn02sTlFBNUhes
ooTWIpFqqrWhgFCOIjaY1Gs5lSO6MrKbiOl5a79GTXB6kP59mMgomnPcEXPS3UnY
W58++cBNF8EJinzjsp4ZLl4/JcVrH30lbgosZP0u9eHO6N0NXWeKSBD2M+wMQttw
Xm1TkVQyR8WgCQScFZKso9g2ay12U04ZaYoOb3LUbhoqxPqVbkMIymC9X1LaWjft
6eLDBWYs2zPH+xwwOMlgw/hPEASHn3EThs9eAgyernRac/tPvJJRAZgGsgiqjJi/
M/gH0A91ke+rnl5z/5qsOgP7c79Sh4Ly+nyAck8ZWbbWOzUx+R1dWXfSJ/Xppa1k
aCRrdszbCNf14RWzb2vu9c38EkLnK5bp0U4z4PP2Yob26zCD6dLaOa1zNJ2lmwIE
kTKPT6cyVW4LAQ3MBT4VFqQMrGnBXRxhqmxD2NcQbSDF1WakpQ8JvlFC8E5UwIQY
ekVtsCNYp7ig9YhGvXNHg48xpoNPuT69mCktBEhaNUypdYu4VANH76FP3bJhIpJp
3z+J+ocNI7dej0EyunaOOE61kTiuHd8lID1PvhnhOyY5aYoJk4GsvhU/CPq6LFVx
R3RiyRu7trcBgI8egtH98bLaUiPXCI2Uwd/476SDDU4=
//pragma protect end_data_block
//pragma protect digest_block
+/ReAasx9f5BGhw4pbhokj2mGIY=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
i/3KQtQMc1qhLFxCmG62vaQKnT1k1CkGaaQNH1Ss2LgplifhwaVZL/YR6TFxQsoA
LytH2+WapPrd2fkLCWzvumM+X5tY5N4Ae++wHJ5M6pWrvFZKQFn3RvGoOfvJ1kXs
LwxLAnIe4HOAHgLn3XCWXJq5XOh92VeBpGKVsHZSuSV4gifbIah4VQ==
//pragma protect end_key_block
//pragma protect digest_block
Xaw3D65NQCyY0iMSyusNMYR/TPw=
//pragma protect end_digest_block
//pragma protect data_block
miZziys3qkWQxcHuETx7/NrN4Y0lQTK5uABVbT6AxzJX9ZVNANhpd/2rQCgGRNEX
JA5Ot874iNZrBwhcZ0h75nJtP1GDy8W8op3SFGKAe7WO+QU+3HiEPNcsYXz1CzKB
0YdZqvAZRVAKyzN9nHFtls8QJXURsjE7vd4lv6cqmR5PsFhYru4NQzfvtDqYqx0H
jSh5+Ad7tbNDOTwJeK0mlepR4WJNmK7lqqKAhMXgjHUr7bkHPmJEC5mFgDuesUEt
4kmRyKa3CnzWuEuw+LU+jp1y6UUv/047A1xe8jJAoF6JZEIwi2pNsHMg/NIeIi9S
BYCazC/dol0caxdyNtJvlpKHw0YJ2EK2+eo92KfdrA193mZGbiLQgs9/G23RrF51
Z3qf69VTCojilALleh0CWwDQK+TA0H8pfrP0b6LsortCbrpu77/RzuSZfO48XDX3
G9Vv2bXsHvpIrvSZg+zZHWkGByCO2SzJYbZgXeqdEb24rRnCHNG0Yox6aqBVBrfw
v+EzapFkN2wcLkKMaCD2yFLJEBuHK5wqM6Z8MTAN+vemqOgxvQTeFF0OWOQpF3m7
Iy65aQYBqlvGLbe+DUetwExxCJrLs9Xb4h6DTlXYW7jlxmo9DDynXJ9q6BYB4Pya
557k8nzkhQ8a2rsjePHsDbJPybuT/SxvSGc3T/xfcSYxu+bCZ3qFG0JutFY7U0in
YB/8suFnrMjSJnp5331BHhsf+v0DNQs6ONHvYbBo4XAWk5f3X/ZL9lhv3bxaqkfu
OllBYuGjkHNSsuka7z5d63MnIM4E3RJgyD9LrX6pfm+D5Gg+uwgSJqAzHuXPTRqW
zbMUEqeJFY93BR6gNMfEnG8ela2r7zaOw+1ISOqSl9Djm39Gxf2Pb3XHwLQ8sx1m
MD0GTX8g886rdNtoxg6nZqZwb3juHo2QDvKY1vYTa5RM1vUnDgJ6hJHBUwBNPfr1
g8rWHH2YkDdWVdlyEGQWX/vzyFLSM5N38DlvYvYFAoS7d0kt2ZyntyjKOkCS023j
mx6bRPpC+2i1TfqLoZNo7Ep4BcjZ3GTlxHR6L0KjufxP4XCBNulP0KsMrRnAzxMc
oFyy9Wvg7w8Gtrc+xoMhbbVTSk9qV7V3dwXP8ylpFZcz7zQB/W+tGAYRFt28yl0a
Uad1U2apFs4Li2Y80kmxxKNl8JseQ1KnPugXc9lSx7B0UvKYmWcjiHU7wbggkvDb
8xfxYdLU3RKo3SLTnggqsvoJ4oUv/jWYsv7BO8GouP2zaPU74tEjbwlvNBcZ6Zfq
DkEOWIS9hvv2kQOA6hreUEhXZDHSyuQWpZd3xDoyIjASYXObsNjE1zvf4Hd5q+eR
cat10YEngajvQKncVoAc02zmlYuynfo+74V0nRnVHxiIgLiyH4Tm2RHi3E8Bm0Ex
3OtNowZhBSrhx6nEgIjLpvXBlCg1k1170nGy/FbKM0EsqqITAkjhcOpXYrPn7TqM
5+RsPGF95BNihoasU5RHGwwFj7w0yn791THMU+X8DmQS7dCE4rse8wo6oFljmPN7
2XnLmcQ8NQuBo7UjNEwe1CDqWwvGiRsHz+ucNVZN0OcDNU9agLpLnVjUtXelNiJ2
+Xc1PDpLB7iR/WqwcW47OKdb2rB1B1/wAFskL11FUzHhjlxFhv1im8V7gGympR/C
sqzF/Ny3bojseySSE5KZuWE7c/dyU/9Dz/OWRgq6XfzujsomLD5EQ/rnTfYYWZ54
9veKBJZ92odaT5mSbK73hbAOGzbnA3fA2ghn3/UsA8TpdQwf0cTGs2p5LiPYilPg
E1RgOL4HwvfuziUeHVBYS+2oL7qMZ/laJv4dgzTpLoh9fLLqldryeKz8diWKJZrQ
48QLjW3XldFvUDf23Az2yeyp3MsvyXXVTIos93yeOvD5RfqocOkmbFDOdhRB5oHn
HqRGU073c6Jb5KN7nSq8Jca48Bfc7QhRBYl1OD0Y+NYMO9+bycNh0irUnHKyeGuX
PVixsKhx6brf+POqSe+6g+Pn5m8iZxb+45BKMlX4tkHn1CyF5n2eja2TDGKKzA6P
53C0hifE7FcVbkqPDoZ859EXCKI0YeYJ+PJNDRAuUqixFFiPQRLbBoXNm9z7baTG
YsYVcB51CazDYDuDVz/XOT1QDPOKwwqRGabI4g/A7UlLZ3QUpFBvy94c/AtaE1wV
ke5KOgL4lDgIQG0lm876DkdGLTD5425pvsMSY64NaR+uXksf7Qni9WUX2DQmw3zM
e0rTqAs5RN9M1LjhwacA6Kcbz0YTDOCVL2n7gVB1diNIE0KImiXFOC5dBVq/UR6e
hcWpMbgvr37v3GqOdeph9BMQ4DmEc0AV+wPk2iC7ZvrYAgnwEWogMEhTuwB0dG+o
rJmT0SqweJ6UOS6JGBP3w3oxtu//MXrTGEoJzq3BaHtCSaYiIWQnevu6B1kCAwVt
qSuyQDVdqkpJzOIiJbAFTiLm7haYF3g25HVsRmUkunI59X6sfQly17g69W+TBK22
oN6Gv97mroxLF2XKUJmIpv8z6UCSxStQT+dpVL8WsJbzjgFtkmRNRS7YQjDT8QJE
KXantH2GuchTDQ3W3hVQjmhQp7qAWnavSBFf+F6A/kvWoQjrGVsos33ZVg4hpSgw
irFLpVr4pZOPkGtCf0AAMORFfBt73FNftmzxBoM/GOUGgHNM3MLryuz69rTK37Mb
tGNLTZdwXWsrLJQrsI8GDzb/OEP4LpSlwUFLK+aDm7dk9OPbl0Sd7MgAd//nNz4Q
GAGD/9/DIsy9rzU63KNk1ZsmyG/W1gi4oo/DQQjvxFONPfWTr+jSIBvRyc+Y/0sP
eVAfrIKJ3LTi+sad8fMgRLtXo77o6Fg/bpXoi3ff1aiFxVy69Vk2chnvRCH79gFH
8+CPTyt7kx4y7rVTPgvLEk4GjW68JIqmg7iysA716ufjmI/TmW7L/HgKxzCMQobs
pp1YA4eIsYQ/CR2AN3stkmFLvxHm231cOWLjmsiWEj1c87fJZT2ZobhH7fD+uPu3
4gQSFXN7COAZSCWdKdTKyCmAdc3BHJ7m5Hf2NYlqcC1PhesSEWti0OhLON9x6y76
OUhsNZXNqmcFYZqRXHMOZ8DThMVzDmJR3+xIa9de1b30FHOabjJpe0sr1b4lsEzl
wm8sTqJBCjqR6anCEmYelKFxsK/eu+kz88TkYUWNxq/GCYgK0IWmR1dw+GBOMd8B
ZzP0zxkd/69zPH3wuGp6/FYRk74ddNKMN1xlWmJcy7v6YMfYy+M3kYkubMnGi+FM
cDppc0r7nsOe7DLqx6t7/Uy8M7v8CjpSjcO0AHF+bKwSraCizGz7PfuBcOWDA7lC
qd1xsx+ppMSszCJyfkmvXBIwY3mPxYiw7oKEX40NFFgPdwc8ieLsILha1Qs+44O5
KM6CSOTJMqJiob2bFvXiYiKWzw5DN1y4N5dtmJPD7bwDiOYAtpkM5um//a4DY9fJ
s/uKHg/LS+1IBVl10ll6xklOhz7F7KJijpo2no4Lb7YXCqpyJ6EX7Y9+GO6LqJha
NVikwfy35UCZP5VYxmxJo/yQnNLwd+zaKlvOP2/JmhVEjLd6a1BdYrMuQgX4p3p0
iCd+CQwEAzwTrjIRpVgyTm51xtzz8dmkldmB6ZcH+3Y=
//pragma protect end_data_block
//pragma protect digest_block
WyK4+RDjlrsxzQRFGYO+kRQ7kTI=
//pragma protect end_digest_block
//pragma protect end_protected
// -----------------------------------------------------------------------------
function void svt_axi_slave_transaction::pre_randomize ();
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
FRRlLRwANpKVxnMGvDfWajgX6hyhzEJg1RrJ6wUuNUHP2YbgM6O3y5SO0f9IJaPI
tyHEEoMIAxkOcjzee7HWfUUG48v7m/4sa0MvmDWpXJ7yxTb4DsPAiZ9xd3yWV5w5
zCfKYCzoXey8n1ewlbz3AnPAXlSvlVLgF305gJLvYJcn/WHqg2Kf8w==
//pragma protect end_key_block
//pragma protect digest_block
w6jxVCIRYurXdV+p4k/gWoiJtds=
//pragma protect end_digest_block
//pragma protect data_block
WWHlv1N5+nRIcbs+/ktc8t7rKmUrZ6FjtSECv/UE7RxdXTnxL/KaneFfiykLv8k+
/x3ZWSe9kddvNISwYr/9DyXtzM+ENHl543txPTktZY1JWonSBfQWrqs1MsKSw433
LZyQSp5+OSaurKuZtVvUEi5YG4gQVo/i4UmsLoVd/Z5vRCgn5r9O2GiKs1XYwR5J
5jRftQ9gWA1gEL6TX5W5dBxN4MbM2jP4WOpHHfxoAKOrxx0dzTAbZ/oWWRdHgKjh
YmUGMiSBrUL79+B7wYCb1apKcUPmM1B8LdBilAB3wmj6n/Rels6dJNj2C8zBdaXJ
QYmAVIuQmopwGB3ONIMxq8BhbM3rhYJmyDb6NGi0LRjCPoARImrx0SCI/XP7zVXu
oU9FgZKrN3hEQ+Mq0sWWwVXA8tc9lr4HBmgfD9+xzHxXSl2bX5yQ+UDLoQJ4TdHu
W6Em1K0RlaRZv+4pJxVvFqwg3USUOcjIavqfXnNJTvUdIlxeZThFlLUyFelWsVMU
y4sFoVYYlm4Q60k4K8acJlFWhgNozrDWVQdUHFW5JYerk+N3QKkBP0COyP7lIImq
PDhOfnuSkfW8sru7p93JZxwglKtFtZpZyasJ/wocrb+45HAu3SWX/P2XorbGvGbw
EH5nr+gsldcOGj6Kmd4Fl5686m/emLUE5tn+gKm93vNOmfU/7FCQobVureLpFuTx
m6VkWReq1NajKALo6UzQ+q3+hEhodxTuWOPctNtjTh5Y5thonBQyLjQmNUtt//Z+
eAh1YCVmccc06vI8pwPqo4/JBX58HJ//8V1J7uuT11WFePiukmefTWJQ5L2SX5oa
0852rSjbKjPBm0DQN971XMkvcnfpU5CGFQhsbLfMmzV+Pyc3jmDi0DBPAx+hmh92
d/yuJz6DAFr7NX4Ivmrth4vRAH1dS8IRKJUFLBxjpBC8hUzlkBodZVnptoJUuUSQ
h6axy5U4nSPa2dBJw0LVeIdmmSfSjbY6bs1lcOCYILo3O39BkYoAP/I6llFgC/GW
fYs6CJWRoUAEQchFUIeJ8lkHMsvRsCN4D7mNVEpwSOZYE1fGOAF1Opl0uobcBDw/
JNxa3+ZDsHXyiFQ+688b4NIjrrDMU8S5vTV7hZkiZ4nHnAHOCpHS4rRTpf+gMveB
VZFqRC1bc+lV/8hYrnuBxa7VUDcGWrpsNJU/zEs9f9LTZvYPtzPOBgk4/57123vV
zJuHXE86or2enqH4B//Pv65nTSx/WnxNtM9dWiHoStrZ0jQRrZGg5SDX6gmabpwM
J0rHqoc2V3hnO8LdFJ+n/Jesh1f4g8COvn3afjV/yZzxFixYMqcfUYGEIUlGQpM8
YzbMhExajLYl9EFKMgSf+/EW7mVExBv55G+v6LRljTQR5955SdHbmmxdGzeUCcWO
ijl3BELRQ2c7awOEGZHBN5bTrWRKwKklPix5G5jQvvZA0wYgR6B0ae+FhBNeDawN
IUWt/GHcf5tNHpfovPCO6M39MDIWbMCKgyhl5f9boq9yUrsOaj5jMSG3nOsMJhld
b3udT6sQmYbcrZgZgPhHhYpr4doINEzv+H3+PbcNLbgYnF1JeYu5+G3F+MlvNB6c
qmYhdZruaBaknkwfuVa6AEnIdQxAWBEpUp0UHa1xkEZhWjHF7LjPZPAPA0pUxmiZ
Gp8x2G+pnvlZpej7YwxbpQ1VTF8mbiUev9huxvF3shA+RkqVcGztVLrNXm36HHJV
/Q53S4T3LvUZgotsdFDDGEDYH7zyyBd4vEZAjwz5yfYWsbbXEPF47VeC2tqOnc12

//pragma protect end_data_block
//pragma protect digest_block
Zsdw2k60UXl0uxaDks0USR+QnFA=
//pragma protect end_digest_block
//pragma protect end_protected
endfunction: pre_randomize


  // -----------------------------------------------------------------------------
function void svt_axi_slave_transaction :: post_randomize();
  bit data_only = 1;
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
IHZv9u3pgFv2IKvM1tR7PA1Vj+8yaksSrgqU/OLAGrc361RzIMJEj6ubeoSTa7LD
0EM36jBgRQLoG0cU3bqfwZUike6BePYst54XxcHnMHJeoyfqvi9BCKAun8mVdEFW
7QMnBuwumg+mx2ozS/bBWM6t+aqRYM+WcW6FdWkCWx0g8/CeXWZzgg==
//pragma protect end_key_block
//pragma protect digest_block
0WlS3mPeqfyjfgv1ghpWfFzx5Wg=
//pragma protect end_digest_block
//pragma protect data_block
+m4EQFJ/Wtz5McFvgb+fi3ECndLK32PfXvdsA/vcaaXs1szN9/KOYr9l3tHK3HbZ
D1DW+7DDSZUejGds4FYzmA6Xt1ZM/PQ6Wip3DhCTBaRBi38jHnu7B1JOdiuZufZB
ZFNTK7OjMipFQ5yMqeqNY18aY73K0VUwTilUo4MJPkarmHRG4Xfq4m/WYAxBM1fh
iSeXlc21nxN2Gwv36HwsxTff1By+kvpzSSNPODPUN/S13JiB464ak1nylFE0RdKD
oEtUnUx7WpYFnfGpEmnKJKDEIvKpl7nMCYnhL6s49Qzw4UF4f9I9oTyunNxRVPAu
kgMM6DJxLp8u0pPgzlKdA/cUciA+wBfWpy52JW96qu04G+ir3z4sRn9BJQq+IWCT

//pragma protect end_data_block
//pragma protect digest_block
hrly84v3MCYXbkk/7HV34NNUoQE=
//pragma protect end_digest_block
//pragma protect end_protected
endfunction

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+8klnsttAir58Ze0fXiiWyOtqt1kdtDyDrrYDBWqhDer8keQyyD49xMkOQTa/ovK
O/kjmFbv3TlCDKdZXglSmffcFJovceEgUKpe6VBAel0JD0CpKUAMdvxjVkFN35Px
g76DDr41peGA5dl65lzWuWzXfRaWn9X3GjpMlmHkVNHLcRvdxWD5gQ==
//pragma protect end_key_block
//pragma protect digest_block
jGUA/eFi5Tz4lbT7eOlmjVIipO0=
//pragma protect end_digest_block
//pragma protect data_block
JRrB5bzzrClN395kywBj0dkykLPbd70a6m4A4ZEiEtDQz2kSZAfldSVnm0IKQwaB
36JZI10tENtf3zSL3PNoZZbv9uT9rQZwA5V5ClIIbaXGSlYQxaRzneO+IsruGEjA
J1IcAa9xGbjj+ln1O2ck1hfzShbUEN3qLxkCR88lNhlOriCUppLhFvV9UEjwygSW
8QJnKsOP4wFp3L1/WflWMQytpbiKde6YH2QbbDlh+63pJ3HL7x1S7oGPbUpVnSaN
+dBYgBvBY4rUuCLLar4Xk5BTngYG4Y7c1tYgf4Le8JFsR5bkCTN3osvRtbS/AjVW
oOHwcWABmK1Q7MEkRNb4s8UZENj8CvvzvOU0cB+ROD1AU9CoXuHbSnQUP+MiFgdk
uAeM3Sk15+H0UjoN2wmrwjaa900WPWaCJYkL08aTwn97NsZJv11KGQAZfr2XD4Bs
UrIVLLYWY7eTL3jlGvI4vl77lQ6K2LFfg3Q+D7uGBEx3NHnAeOAqFnKmAQFkqEnJ
oLnRG3ZjwyiRItYEqNJDbZtlmA3epRv2G8abVdSdv8TDVMfGiJTYKww1kiipAa1v
KWSbiL4MHxnNgksY9OfLZDQNCnih98+uNSrvSUCaBnIjzJ4Ubg+89XbJQCdHN7cr
lcIbpL3oT7eHDvfhkO72OR1XzP+BWakmBy5jAZW9UM3XHyRWGlPyjaflFE4RTbbV
KYfWjUGdG6zVRwIhzhBCjiT+ciu+CFR8s8cpsO8nYpVXiv/0ZRXv3ENun5C8IGGO
5GZfis0BW85CQbq8LcIS/Rmyh3H7mspNq9r2URrC5/23NQDstM/qPglS1AtT6E28
nUv8dxFnZgaGg50aVGFsZsTrGkltTAfwPeIAwexfoICcSnrN5paGzVnZu9b1BKLm
F/f58Q0b+gIPIgxprXNwO0T3T01QfLLVo5onmmCkuqVWXW8U146aotsoAyX9qxkC
CQRN06slGwssAVjhOQuzM12AQdJ3dtffHQdcG4Pp9JvNB1ySpZcUUcHyWKtgKIii
xB7rkVw43mo3JnXQ7vaGDyXwozDd1QrRiilW4qUWD0+wiHXfSLK5RfTAlu0+5/KC
/ySXoMW+z2GQNObsm685B6n2U0J4Mmab7DbEKc5lf6Hpz8o7Yx5nWt8xZHZ7u1VQ
DgcZ77STz3depz7tVWJEhAJTvmLI4PwmCeZNHIKD9AFGjzK4iYC+uAAq882EZguv
5gzDhpRLsVWMd6VQWb4+5E0OiqhEHRRehqJn8Q2Vvo9Vf2i5IXqLcJ0C2yehszwp
LFcZ8TqJ7H57q0WUvCIsH/UMsZh9nJAJdFYmYTR5VrV3wWOnjBS7I7netQVaY/ie
B4e6jBXr9FMhGTUcxFoo4LT+vNKMyqvdmDTCiyPI88oyk1++PBMSlpdUWRFL/giH
kLJP0v4JK5ydtpEeTDo80E2kYCJ6fnXlXblldutv/pFNwPpJxx6kTrlreWz7EPrd
qKS3y7l5eSKCeluo95c3bWB4Xkje1E6H+nwdtGGeSLtO3uSMun+j3SJbbV/n0fwt
WZ3H8dbo5YuXwoEI+sXah8JArvwt8z+xBhbDwl5n2IdzfzLHEnI4x5HvOysLY1WR
NdUDaP2B7G66CyxY1jjLnRLZIS4RWC+gvj+B0lGWSA98Qq5xy+rElIyAVqvJ6PRX
TDfIf6JmuZAlaMylg6brk7kXlz074yq9oZUd9QmFwalLxMRDBWA/6XoMNGXNFjJY
o6noClfQN0ITNs2Iia9PElTbiOxwD9nYOwwJ6ZxKDDKtS6z9BvwPnDaIntYrkLBY
/UEwRNZaF0wd/6h39dhtZs6CDov+17PJpdwXSF4Zabht7tMW+n5pBbaXTzDWhmPK
Gslt2sTww/MAnTcw+I2xhLKKbHSh9Mjb7QBw/c7/JQetL9Otb1NcKtOiWYt6mCFX
HR02JDFkkOO3hCz8nWoyCbGxOnp7OY4nEnDBhbPOYjuwT7RRkoBq+xUh1qHyu1mb
jHoyPMGmUEwHj99LBm3WVDcFh0L2nSHaImXLvmyPkxDhpPBIaN8nAqsyLRKAnnuA
B3TedJIYd0aHSKBNV62iwjn+PgkixrkMG8Aok6mnS3+uEzSy5ZjWjxL8vGeZI95T
r3K56/ODJVofzfvZh+9+3/lsmxGpM75MunDn5OlJaVteBMW8D6lzV2M90wYNze4n
Y+NdnodMbaXxnwgGzPrGnjaGiqoeXO+bT7XBscZ0B4mamq1QEZkZD60TkTRIx6N2
HIOt4FVy6xBnmIhz6qSRbBMGNdHyRgwqZcEnqrGYO7I5myJNRVtUir4NhvxX3ooY
4C0q5YrbfJbCo1Q9+6yhwCZ1DCqtuTQbXj1r+j1nDNdAJ7F+bTRoxzumpSj7MPZZ
wPHn2QgWG4h2USmPWjA6Ne6aXhP9WuHvGTbS+qb89AEoJK8xw6LA7A7d3Gqu3me/
+5oc1X4kMFz/mw88kKeQ9bbLlRPzr6dp4fDg66X9DL5sYYbhkMyRLWgdSC8h3BwT
T5EPNU6ouyzMg3V5z5JrJ3mIyQ0ULmh5dsGaJzaCwWOJsVC0byhKZzFFwAHb1O5h
dascq8HnxrZuux5P1E6U/JtXWTI+9rDK+D5FiwvKodb1EhKmbnxjZHtnBBEDeAeF
PDRsalTE5E2s0ZCwPRCka5HaPZCK3h6aFvT0ltbn9eqExqnvdo4JgtO3C0E+C9aa
4ZAsmVhupLQDeUyC8cw+AysB7v2JqxgVP3/y/De/LxbxmnrOuY+sf+4dc4oOby5d
RpfJcSLh3F86gZnMb5DAOL1oWZWfYBLv/IZzaJTySfx1oSxH14x5wQizGS11bnsB
lCAz82YNJqwjZK8NcteB0/nq+NmuSnoPtSQdh5Vyq26E4nJf1zaTfqHLUzSySmBp
bn8JMcVnHlLNimLLFyf0C7ZeZm0DnpVwWtiK8XR8mAe5FltPJB1p7pW0miUhWbcA
rpBqoMge1vj8TtSbW5AAxxvXQIvjYfWJL+aH/AwhaofOm3j4aHsG60eRcakVirMy
YAkGN2jnCG0EeRc0WSIT9Q3TnbhLT50jGmzid67l5cfb1PAcdkR8Z6vilL/IgS//
2AaFRdXSjn7Whe0HDe1smNQgTaUzshxo1RByJupayDyAZQ0HAOreIX+C3rn39ypk
+so13oR7DbyBMreQO2kr9O250oyAzhgSQJwKgogi/mHDZvztDVYXpp6hvD7MtXmt
+XOrXIqjncQzpBWF7/zq4/EROq9fibqdMk6nEwUR4CYFxOdk5Qj5NAHDn9fCJ+5+
ZXQ/gLWlTFUB9Y3aOBFEIdkFSCGv6LMvxowbYNyy9jlCMMu/Wy+9WSCuoVoTEplG
5V/6qr6QlWjzJXNtl5SX+FxLP1LouU5/mhGlMWwy6ZVaxXkrr/C5jyHhg3PrpCl5
hdbwGVy3Lz3E6rnTAAMn1FO69Hr3tE/oAf2wolKrvEITWbSPH/6ImIksHg7G8pIC
4tOyhIdaetat+0tXeGImOJL//pVIYuVYs6ft8JM9OdGir8FOZvbqCKRd2H4KGZO0
4W5ikmNs/FKBgoKt4XiWfIs8OYRAUJXmnjceMXWnxVv8Qc46fP7x2iPAonfalnlA
yOS+MNccOQkbmHoMPU/8VfKevO133AhQmNyDP1InpeVrxoI3jQr1V3ZgPL057VBv
hPZypd/NzhlTGW9CJSPDxsj3mKItsY5cox48PYLBjF1OgnNIeZKULR9+555XmHDy
uUCaPK+wvrY7eiU0fHqGkgMA5mRQ9SaTqa4NGosGBWjObnSPSTGDpu/ZnWLt/CZf
aJkBfc1OR84eAxnFosWouwyo2WzLobu7flQQ12AXsF/QecwpY8mRHK8uxKfaj/e6
mUTwRbG58g5ePYTpuCwYdVPwAhwQFv6pJQcHsnxlgOQ3rqvJbKUHEwd3QatqG7fG
dab6Kuba84qFyqmJEL45xanroXQhs6G6zOWnMCrZis17U2Wt+lDUFXXxgwSQVOL8
/mfHQvwYuIlTF/deXVCp6chD/zwaezpq9pmyqKhvdmC1D8QpQC49MlkCb7hNiynK
9TaQNLtz6IdmzWQ/xhTZam5HntE602tLpJhJd7a2l8P2jU7kVGHVxecSP/GvF241
LdkRz5edsiZl5o80qdCBMhAVBovaIZ4BkbOPDGvDC9gg4XNQvvm5DCpXaq6H+o3L
lOwXj7XTLraeSyRd46mwj9CkNEkn38OGA88ls356I67ApY8OxXACV5Irp/S88Leq
Sg2MMfJSYAKeJbPkWHB6lnCUzmNa1bn40VwKyYWU3LJLHl1SPVJL0ksEP9E3ufMP
ciScll7jKaIlsGXkvi62YM0OBh7dNuLdzAPXcwsthyGtOuuCpRYjCVUJNCO3RTY0
CHj4+YRf7b3fgqpw5eG3CWcYVCrwzWAU4FRpEqe2R5edO2i8/KcGwr70v0IvWgZY
vqZY6Rag/nb+kr8g2FbBttyXLoex1S23lQYXjEcbwkG+XhDkYXnjSG6ARoinNb8R
/jSm86wo2G9im/JTMHrB6dodPvBM0Qeifuo3EWitOnCX/DGtd4EzbzPQoID/ZTAG
OEVJG5LyRlrvXqKIvWicc3q/+oRdbns2PrxunwlikT3H32TwWbydYVW5M23eUz4F
dGR6tjUge65AcORJUgBfgvcBAOXP7P/q6y+jg93rYCV5A6W431Mo/dOl/V8XDwYR
FcelGONpyTVd0z6qP6Ioh2bu/X7hQ/3zXCpfTtneHXx2MQyL3VQmxtDDXWk53uyM
29h0OH/ZShVHGYhGwAXZNZXTT0WDAGyZn+z3LwHX/M9E78vMDhYrI5SKiDI2sixU
CZm8g2NB73/EH5NuKx9S0+u+Ai6PGB9Kr74wGzpWdqNnOh19MRnVwXmBTEUDlDWq
rOyL1q02lsUipmIUxLb6dBTXKnCeVw2Ysk7PXibxJkLLeGil4w0QH5df4A3s0EoC
EqR7OjZIs8gWEPHubOUOdaZcALgYinyC6NnUT2zReBa882zFqOYghMHAA8SGoIz6
KwSynltC1rY+Sac2b+Mpa9IXN5KGK6VsKJ9kJa+Ad/c71RI1tyuBYOw5wuK6eVgc
Nd7j7w9tkGpelFKAEgkLv3Lrqwib1mXZabo4lyc/+NI2hiqEUEKgDM+Q2gICtesO
bxmOrBGuakSJwFEeZ8fl+JcZBwhhZ+R4Gm0wmXkg/wPpJQ72StG/30VSB/so/Mu5
QxIgFhhxrOEwwWkJ4HdGuxtkZGnzZLu4+dw5tRAFrVWDYpI4wChEsj29rBvKfLFv
y4pMpS+gbADlV/UfAMnoNtDMwVJq0p+6X4vKpIKINigYcCscCLQAlaBhRDB6qQA2
X7BKEw/R7y7LsDBAKzAkPQ+72hDdSO/KJMunGd2LsUZXd2Aq4tj2vFTx34fv22Cp
ZdtotcGxsE7KSTXMSJA/51sLaspIwvIRX4eO4A5WamgOyqf3t9Yiv+ro4G8PBO7Z
2shlyWVD7IeFYzZHKGqs94wav0mPl24XjyIf4dQrSjBOouEvaP2xKnvs+1DCzJBI
TGhLQycZ1ibYcXrxnOKzMofKvEgh0XatzoO+fG2fMb/mYmcV+tSGiu+VsekGai5q
eSEAMlRIar7Cr31r0Z0/OTg+BlZ1fz1JVpNFlVp4SJom93/g4/GvGZv3JRwI3PAs
dJbef3nleZanRhrSEh40ExXD7gaaen1oIbPs4sGfeptsiJmkghHU6+C5MQ2whQVZ
Wu1t5Z5OkxkGhfSy3qOxsoe9wHoEqILjANguqmyAchY5CJnz9LWFoEgW13eYWCz3
R6Fi9CE6dIMRCLoKQjKrsgKbgGlVreK6+ATWA+usP1Ng7F9Czsbx2dXb25rXPaJB
tL94iWgCx2LfHxN6FYFj8RhgWuT5Swh9sgVXj1bA7hEoW69MdTEukMGQZSHbFQBC
tLl/PIpffAEoNC0kKTgENEDcUjtnIwELkizDkFmbZff37JnMohnbFb6byozdxakx
FwgD5xhLG8uT2sKDAgSH7ya9Y5yHw8jn5trVdroT/YZSN/Sh2k2q95dkWxsl70xW
pEzm7uvoE+SM8pKVSGO3d7W2TOuRM+rtcPZAv6klCS64b51JJL+19YSigeAMYz9U
W27erAQSCBlYb+vokIyzXAxniiCDiQWEihSAeGm2aqpHXSSIS8wTBid2V/cs2hl2
YfM2HO2Iqu5336dtRSzrQYuhHVXbCeU51q2Cbrs+c3UEq1oAqBZxp9Tv9hNNQ7WL
0KcHPP6XHjVr8+ctTX1vkXHVFfBnLJ/PxJRETayGFIBl3r09R857nI7a2uH0bs+J
rI70Wo7tO9b6zU+1vcTdTDZKrHIyJJ2cmyPCpUb5oU1djRLtQFoKbvpZU4Um9shl
iruYGQKj+85WPrXaUrJxA+ElW5d5oQwPV7+Kz4Y4VKZgENhFW/btHH7kRG2XFBB+
tfUZNDhq91DzJQQWo+ftXdphuvADcVCkbnblqGIS/5MFwEKObfVGKY9NqXeh3IDd
IbXUZdzvbTaTFJFJ+lyLnHSXpIWYTsspvxwb6R0Frhb5D8PwTc+PBVbVD0a4YoR5
NCulUzjiMl/wPbEePhORzXU4mABxjN/iR/D/p+vnYeIfOKjGnQ1S73Vz8Rb1E/Wr
j/G6pICCNzyIem3CZmOyGmjr4Zahrpa9E14XAIbMnXavj1LFCi91dxiOAsNnP0tL
nKO4xGwcPgJ1NcJd0y4DKRZAmGPvEyFn5wVyLFp4690JYs0VIWHJSMSMJhwWOo+U
7m4UfuxyU5oaVwBwS1BbfT2BjLsAF46kQ0OEUdF5EaCnqGKYLsLynLZPR71tPyBt
KtD4LjqQRwjNbPsZ06ZKytBLk5IpGJbSpMGOfRQkrKjXOEHGS8AnJWI6+E3zbxFP
Q4rcEzi+P2WEuiu9AnCC91hBtIKvuWe+xeT4CzXMqTeGllpy75gxQTcPjbo3GUhj
nf6WHi/YjUow5ShIrb76WpWedRdW5xQWH5LJ67Zewi5gG19b/7iTferGQhswKX6s
lXkDKaRPY2bWOdzrUCx3goT9qKMmD2Yvi6GB9QRCubqeZnllbMAxM1IieO/l+Xyg
NP/LTPhfyLSekGndtb9waBMa/QYUU+AbSi1ll59S++pp5VeS7lzdOU9yZ5yIhxKw
GW25hfCBO+87x4MRhwDjug3vZju60L1UchnM3ZQzg3x3wv89D+krMDrAPZ8bnZv8
Vs782ibXY5Qxm07P2RPCSS6tXCe4KcdRtfN0rzh6rzStM0nfbV4J4euuQSNrNpLg
t9Ljo6QsqgH4ApRxiFbwbi/t6d2Optyelo/BsteG03euqPJzduLbpaKaecMBaANw
KmV5IBQS8uUE+TEu5uJzHhzfN7YGis8wvVJLUYbZgwNPB37BaIQcu59J6LZECvlP
5x5ABbzRC3tUW3g/FUFhYvG+0py/jw320oEOxs9e3ITYn62Hl/SfW6pSXjW1MBUj
A+wfmv0pdUCjsOqBau2e5V/g35GfbBebiM8bTzc2aRFxBSI33A3/mqWB/K8kzidB
3zMshNYxBbjX7g78ba5a/6GXQlxyreUCFLw1V3UiGy3JaFL7bie53UwQWl53iSb9
sAQ3FAosfx29kNDEkGbPXJT4/YepdR46+KZQcm8P6t3+WHurETdGjX7z800PiCtq
BhEo0aYohuatX/EhmVk3X5U8GoapsbcL3D1zlHliCovSq0mK2+odC3HaXnzgNj3s
3Wg5il05hzLl1/mvRIzNtzKV0iCT7cZpoihsnFYs2fcILFjW5sLzN5m+IZ5ATOpU
TCNwi45MP5ygTinHAy4I7FEEscch85O+JpiZ8C/IjpY8uEVh6Htp++XK9u2DinU3
6wV5nUmsA4lGOLDC1tsAivc09X5RHONk0yZZ1BDt/P1PsqtzUTC26U8tJAxSLhz2
OiIpxaJh/g+AZPckyLTFtaONPxZZL7wH+36zQsJZLMNt2+9QQlB+bmUd9S0oHHik
QiACbkd1WQgu5zI4OUMiiM/cRx8cjfMfOG+L6dpNRliBjiwy07pXLlpLb0zSK0cT
bzsBhYUYXjKwV5Tmh3F3hUVB7QqaN/2l3F455k0X9ufocf1/txsqxK6VKSDeAOYB
qCXZNsf4YJfvfFspw0idO98TENbfjCK3Fj86mkXYYXYb9802qgdKxIYdd/0DwVcj
dk5DEBU/z9HjBiKCgjlv8sKT+mTjeHZGWRmad8TAaJ5/r7RVo7T5vj3jES88S0ZH
6vFf+iACl3x2u+8BOmBqzNVqIkj3HGdQGHFma9+bPKGHcNlkU+rg4tWv2aNc7+M4
whOHdFd1O+b0VE2Z9Nzmhw28Dvr76VxA+4+hEwNYYUwE+vz/4PnKR27DDNxKKWis
eGBV2nF95UeRTBfv/0TnRkeWgKTbgr7oM7EQY+3GbGzJt0+nOiD4Rl23cFsHB5Qo
NMjA7BTwC+WjU9tz4gUUWchJcR5piWEERsoa0cPwEcdWOxNqjbcWK9SSE5GnOYCJ
r+mQNehOUmmvkPC7ZdShes6JtJtSAgPQlJFOqvJEK4ONcrS4iEOSA5pniHIG/Ket
wva7dK+6MVHe2w+KksDOIPkD4tLkFUP8c6xGQS6eeHlMZl26oW0A2tFOzoOvv34S
JqV0xqGkeVDe7XJjMZTkUVfdaP23uYlWCK0si7GxUyVxxHcCTMGXj+5Il2ad90pG
3OXd/tge5/ize2XjkYA42XgSuVNIk1k+kZkZoEoFDgqARiuqDR+cCzUtqlOHzLWy
b9CYo8nwjHBxYuG5ieL098kxq/djstf94LqnxVTWMPcm2clMvykKNM+QIVCPra7j
gu+TLE2Rux5uB1ea7FtA2QoXg5BHCCn4+a/C2rB0rheRq/MWTnuYCmZRqTgari9d
wtNCBXxsv2De9wnPtTsdhrH/GVjl4RwXgKqfVcC/l52KdiF1xT8suiBu4rRK7k5k
Oj7HjmebyUbSED1i6Ax/Phuq8uqsTpEWvk+bSmIxu5fY6Pl4Ql350pgLm8Dhvto1
9y541rpCAOwKOwfPvW4wziT9EYc1EG6Lsn7IQg8uPNoqXBoszyewcxIBtemD3kHg
pNgaQ3sM9dyxwZf1bSCc/CnYGqkD56jtHcUgWmerffBOA1MSANOrfHHBEKRpiys1
e7dvZY4RHlp1E81eH5/gOAf+EZQ/kS3P8nmkmVvhK77HzXhcitoZ6TTn99qqjkjk
AEXNosm1KqUHq6jfS1WF27wv12T92yI4Mz/RG2ZRElcYZCyDSujBjqQy+qWMzOZn
EHIzAbbD/86ZvZVIDglzn5zMSvEU1iMoVp3aDnSwSPJXKAB4vzlEoWW6RTmkXleP
LR1Xq0cMkZU2IVkkKtQcQg5MXw2HxhtiFu2yWne8xv3QBhsZt1r5EXgWBXrt2/vM
cOP6YbhMyuy5/VoCVdZ+JWk3akexPYMMccvWeCQZ7Se3WmymcYNdVlNweB8fqZAo
fhs9/as/sXLVR7TiDE35ffuXbzBkAqxfN2VBKwTq2VG0P/pH6n5u84JrDcczl8+7
CQVtlXUlSFoN/J98W8sSKSutUYylFGhBpun8fw2KAxLnLTGlGC+jnvAoeMQraybN
ZRG2u6e/AOWz2rfz6aQfa8jvDSzXcMKc9nReE//mtoaBkFQD7kQ5VIEuNgTEZ9Lz
wNXvRpORBWkQ+3p4e//83/uqWhAc0c+2QqwlCaj/ml67Sxc32nGbLj9JshY5GZCJ
oEJfQGHqzMxR6PYa6f63+LGB2Px7t5M+AQv76P2cSxP9gHlryDrsY/FdixCvtLAz
EoihVfUP6B5xZvnBO1uNSp1S9n1cALhk51VZyO5T+jQsdaVYh/9WKuLUbMVbLLzV
GiTnsb5YJ9+sXDP7g3n4ZHb/jlefJMn7YrAqV8ve7hkxSRR6Vs1jKo8IZcDszaDq
yAVBtEpsFsC8HZ6Rss0f9Gkz7hT/Sw0TGZ2L+2JJjTJpZkp68orhFlNDz2DY9N4K
vTT7yKesyrlvLmr4OPEI04r6QnQvd7/y1rVSdfA+hpE1hoq6q6ki1y+ges44PbdS
3PXlDX6lxs+78TQiJEkhKpfCNjYvWjmA3pCOO0oxecTvNLQxzMYnL7ys2WPgBK+S
GyyemN1cgtHPaRURCTg2ge+ucs6Lrqi//aw+SGNfxNCmq5eCNEc27QrjjuaEjDaA
R3fYYaaC0cV4ksOnKjmrmyOlXiS4UumLUXtY8Nz9mkiywO87dMgVPVklLw2yGYIW
1hIMNeBjVEluufO1VYiBbn1z0x+WRHv43c4ejME3JntswBwyayyMybUr7MKEN806
HwzcLLBxr7jtZcCNCmWdU53V9xhJ9GqWi+DwpQkx4bCXYW8m7YketHL+2gd3B9l5
LuddwaBJO+3pLhYdp58N6LPormgKvnY9AHCgkEpdMJribTiWAWDhzOxiBRHE5GWp
0SG9mnoqCC2RnnEb+VbZh7MJ9v6quxL4Tnup465r/sZ6ernI2r9Z1a/8TD07AWZf
SGHBzU3IcMFKG9W+jQrPXR0eNY/+WhhopG13fNWrTFnfRkptbkOFk6pT00W/L6TF
5bXMG/QE64prFbLH1pnfVkv5jGvG0qdXY5zHyL75ekIsIZ6HQX/ob30AmLfSufM+
yRNiIBVMLHYGPMDKhbDrAH/lZ3G6mbGKHHG7Ck7YbKnauVkBAO8lE1+5Bfcy5fLD
VbEvICLuLc3m2rViRVZaMhNhNpB/+RCmvJtuNvIioltk4CuOrJqEVhRHCauBPYot
rMTaNxfSDt2XUhYLxHG8HbTJTDWhu9F9jsq//ywUM1uU4Nphmaf0GLI1dAn/VEkk
9TA9XgiZo9CvczBm460Swzo9bEnl3glSoohgs8uWsojKym3UdE9p0mlXAFGWRoJM
/1cXiy56Ezuy6o77le0JirfbJwVqrIwcKquf68QQAHh3ouBiTkPw+tr8nM8+se6a
33xXnI4T3zFQ0mYn7VYa52P/sbTwU77zgUHRFK2eAFUhx65i6MWQQs8fElDiW2ZZ
HhH/PwDBU0Dzs2BuV7BhdQlgcsKPs6VbnyjtRLLnsHCKmNK2EImG8DoCZC1pUvbn
Z8eu4cw4vunonzX2tBcsxVlGAk6x6YoVs4yHoS0sFCFksL1jL2hCIINYiSM9RjrW
EZaUY6d8H8E2PFIUFloMA7jWb6YcsMPY6QUr3CmDsTGYeVPEWUbKLdSxaM9a3LOB
AdmEv/Lujl7APMcWfAtQQrnmFJaVOpBvg7ahYj0xYpS34rNA1nvPF+g+bySyo3dJ
fxz+aOAULtlHonxkNsPv7BEiflJkoa+G77MBelr3CfYjyQ/jy64qr2EHKFMXKZCH
1gZC5fZfQugPSmqTf1GMUJVFirfpayC2wlp5C8pNg9PFyi7sv703v0724jIm09bq
kUzVKnO7v3Zg9tccb9J3zFA5JYvnNhnBZ9EIBbsYQoZufuYv6bQJRL7fhT402/Iz
QmIOQGbs7ZCZpFaRkvoFLUjThhf3ifbI7H7mU6m6XqSNWlMp16tgRPNWr6dQ20cR
o89asmeu+hssHS6SEGcaAqbwku9l86WwKdFGOsQpVybJIn2S3B5Q2WrhHQ4kWdBB
3flMnliiDkmT0aj9LOaoT5rfXSDf7CeDbqVWGQxMg5C93qTFa3NQkiCtvFnHJb2q
kvUqC9MG7HUenIaR+gImPDEUjoMNG1cYD2BgKfNLQw4pDruf4+n73J/IrfxFkLUq
sw79x4tNaNBgkeHIuYv+Hd+4bxpaTv40yeCg+ALfyYF9GBRjr0RHBTKDhbFW/++U
yhdyNeZQUUTJxLwLBBIbkyo8rJEitijy8jVqowobzrWOI/e1iy7I19VQPZUbN3SI
/l75PZZDwkOZaWc5zhexCKA8jx4aHnSMhgvomjIQ5K0YxFCB5qb08pJDdzMoDdBt
gq5VMv39dp4H+2bj1wDHF8c4cGQZLP5kPVrnWKgNu1JQ2ElNOJkcGjyAAFBUJEl0
kBTEe3HrZO+WYhbueyVzcajA+nuM1dkBHUAeUMd4oZo0jS/uCmVD26by2mSWW1NH
n3qal6bSTrXdQ1Ve6f22a+sN6SzEGbnYQFex7C3w53KUse6+6K1wg0Mr8Arzzsjr
6zFRgTaF43dhX3DssaJMXFp32QN9Ti3+1kFSSVAelHs+RL0fHGu1qCWIX9YLMX2e
vuZvKCvyJGrBpNoxWyrcoQkpnopRgdlF6hCIp+nZiRWF6jXAQNOczTTDgu9S8+xR
v6Wgl5UkW9g/OkPag6jxP8T5ux4mvI6CD430pTvmoxSNOHIHTY7Vuz6ZAjcYPJWn
6DrovLD3PgAyytPVnmpO1skzVV+xLWsS5eivrJ31LGWv/mcjRqIbY+VEQ/oH/iOK
NXYWndM/q/YxMdvHiE5lglFUIsJdHXKi9S/S8IBQ2xluQB8sk5RCcgeB45hfbxUs
d+Fxqe9+2linmaBe+Iyvf7wSDC+h4sAb5fMbkpyU1spiohrRgUHhxMMcseW8bcvd
UVKsr8P24JfVJ1PYOgl16JROj8tAS8SwyKK13Vw6+m9pmWVNHlm1Bg7HFGPK5qwR
ffY6PSR32JtEERv784BnacdaohqmPNGUi85FMOeSnxDjpUb235q4AM4hOUOJb4PG
Kf1kzE+ZxUYpiTjXdrSs0rDh2/p05zkU5Op9O8lhySTtmE9t9R6ZUfgOC8CTc8iY
aH3mNwAV4qooc84FhZLCYNa23bj1+B0Ax6zFzM3ksaNjNkt1lFZ6XOS2POiBJ6Hc
3cft9Npkjk3X+Y2iZg0ECYX1nC0L9jpXNYqJ5gEa/DAhs4eM1TF6Y4SU3ItM/atJ
2mzEr9XZ00mQ5JkktR1gLFOjN7YEWJ/vx74LC2tx0LNsMUU12vsjgW6le3j4iQes
IexWuyXj1zbftCNWZhWZERaYMA7MKcZIiVkazJt2lPpyeEMltxogFWcUhpxDo6KF
rJYdCas2cF1Dm+pXNiG05p8Rj/UQPFrBwqgDNn6zPaMeXlVTR5PLLsaKzPfNTiDD
PF3l06yQ5V+D5mEurNMhQ/mPhpEfFSYYjEX+pw+EVMfCUrDH7NcPLGelU/FgQdT7
rNem7Ou2wo6pGF7XAeahwSaphLmvMUfccuxKNcoXfXSH1onuKwtUyXxWhj219EAD
2qzu1QgERh83Oia0PXtgv/OLiwHT4lNYI5zmfLd57sIKK/LygnomS4Qa2jqkHwNV
VkU+sshVOA2xuJA7Yp2GNHwdkFs1fLoN5qlQPDL6i27bTKhVGRFjYWE6kR7HVkiS
63lavItrJ9tLbQ2NV+TxJNpWbSI2u4/ZTgFDG1EQqDXLVQmNjwFVjYbubIj4PfQJ
Kle7w+Tfxf9n3hZ9PGhFdyZVrsapBQ93bZrgCBJYy3EjVfDid/5GgP5XWCgUNpxE
SsSHCaT5pHz+c9RITODdMez9GX9i0O1vIdXsxZuBFdXm3vYDGZ+hFnnAWhkRcolB
9n024m4kpSVAjM7PGtROKSp6lGqsx7hCr0gEr0sbzAbuXsocpiXlXUqI1xtimMwb
+4OmqrHxdK50+9XuVUf9U/ZnNC/UrIIrF4i+X5757EyY1TK1MgvlAWeUD0gGbSE+
cEsra6Y6BTLDRZQR0KYhabESAfz8iBqwsEAF4UEsuxnT61a4cX8F76oKdAiJJ/Lx
4A5faCdmUx+bC8IssDW4Mywe1dCKs83Hz/B1i7eyiuNyqufRovGbmxT+OyD5hXjU
e9V9ywom8Ol9y4dW2XcSCgib3UQhpsaAf/JQeGmhxj9zOzIJDdAs30au3o+jXwh4
uJYiIFlt/gwg+C+m3Se9w9P8tDzNJ5S5idLrPjnkv2Mpo85wxFvPlZ8znaKAv5uJ
3rEhW2VZ6oIYeCkqZDaqU+n6gnVGVI7ytYIEMayGR0Jbe62UKs/3j9v/tgQJQq5C
jnkleOXukkh993gI8fyPVBVnX5+RXxUPf2wVMdbBMiw3FDQyL1qsUudz434yBMHO
DXXfq8jRWHX2jXspsKIkC+LWz8YBhzPSHjl3lNO4xrfRI2OX/bLzb3ug0VV8BnXX
Ln+mx8bY2IRLxH5rlni2MwQf35HOgv8rSmQTQAcIxXO/8k0/AVvRj1EgH9QS2DmE
bT6rBD4tA9ExQRkCnflO3g2/PsLMBnB9xWkAva80+8PC4/VfiCW+0q/2+2INa2eB
DYmPRE+XpQ+neBJ4JTpdUTJIvkGPEVkMfxMBE5mAU0AHcY7W5qVB5foM6BF+lDgO
a/DaOFtBs/li+kQo+SlGVVh76UB/kuJ7U/qMvhURhon70mIlXJYvvpXj8dRvfQoT
1kmLmMQlGGZqtM2hEHEZhGF6TNt5JFnvZ+HBIdjzAphdRVaEVqFrvyDFD56fxMsE
2vonVdPvYeOw/M6jFyDw9euOZQchDpXjY0w5lEGLpKXvTam6AHR7Kaicf/2KsM3b
xdSmdy/EfFyVK8a8BfsLl7sBnl/vieem/IVzihcJ2vZWEerSsBQXDl68yWY7SQLE
FSjIfvs/Ep/HkVK/go7Zmc9niImUDqUUzmM40ATIOE1HJyDnhjrPp3cw0kjC+73r
8D5oZmFtnXGP1d5EuxiHHvBTanuTpTm5mHUl4OvzwLjQMbfViCya8guXf3yn2YXk
Cw16l9j6vxysfvQbKpvoajEIH4QF+ghCuGoMbxGCmcmnusRqUuPMAIMRDVJbZKbZ
uQFjOhRMqKBb5vyVdF2hjRKOf7gtc165d6QRnlH/nWNLCmMv1MYKWqXXXzdVpTBx
jS3NcfoC4WYGHTeY31ZpzQ3i/VTSkeM+YAGce78AxGhzpZmmSXhOiENkIZCh1m5G
hII8MA8CuDyhYPUeuG3/jyF7cwMeaTY1yFiEZmiI3XEnDDmnV9K1STEZUYhUOh9X
ig1GWAC1SQmg4+jhEPZzmtBOi9lRdUJCOqx6dcKzmQ47dBG639VEenw5KacPrgiU
XMU7h2GoPjc+6OrfUrd5QiDp4RMhNCxF4jM1i1bqEzXoACC3GsK2tzheDek7Qsor
CTJK0qHMeXiApUQuFJEUeV5bqQHb/HDjG+B3sfJWmPFT0HxPEg6yxS++EFhK1RQo
kBsp4nRQmoJ/FtycTEcL0GAtpoVVWOwWWyiKFHjPP08ja0h+CTaTToOOe1mBmMrx
4g/f1q+7jRMDjiAq90vSxApN9wnJq9ZfKRuNHRGeHAI5uSZIOGJCrZt2WCpugEcM
d11mOKcVsNzgpUc3CjltpFsG1OVZM859xDS6JNTBxWRbN2Z+c64mYm4+i53cdXZu
KHKwERzNph2496hHrIrKOXjdPK0jECr9y1/0ymf0u9Avjqm9azIMgABzipRdcR1m
ZMiyv9TgJFd9Hrfquo3zrt3Nt23ZzyTEDC5Z3qRNWXC9Bmxttcy3XqINRLExApG8
ai1rnQa5an0UM7Kt/bnmJ4ftD+Ew5XGns2Bdvwmuo77+rJmDVSlfmD/hswM7pszD
ax81Z9Ifc6LS0KcLC1cdYicQ846k4DYO/B0GFIWHpdFCPEeooco7c0DpDEAw9tKo
fy8xDdD0k6MCv1xBXQ1LI4FMNMzuzF0qOHrW/OO2LZhGBKjy/Bf6T1OsrXooxvww
haWfCWnPCK12wUvn/ac7b/YTPj+SmzhJYQP+vkRW0xHzFPWz5y3l2KmruH41GVlK
Eg/4uLhAGUNMiqOweklq1bqRl4X3PEZMFx5N8xOnm7FY7qBfyfbyxgbEpA0v5DU9
odezUysgJxUUJnmZAFUXnonrfbiOzdd7dm5M+UoLrwCU11viLooBmlSdJgOxS9io
jPxUDN5FjLC59FQ1xDamSORsMDqm9YdLqw8kyCxZgbh4jmMMkTaJVObIohvYpnY5
CCKVajjERNUcLD+SweClq0M60b4OK2aefnMD+kBjG0vJrfcxhb6S/9fPxP2dsIa+
+2ky5IUG9iSb0yloaw5kaGEr13jB7BWRWeiB5+pZDzx4p9sfLCeVIV4460Pmpr3c
veAioJIxfbUIHodzs4Wobh7zNxAlbYvdQBRQ79Rg77xHcXmw0kCh8IfrKf82tFYc
VftYJwTUiA4i7oB6Fny0Qds8iQ6VEHh2m9461hf4O0SqFnPZGvn0DNFDOUp7/e36
AA5b4pdwDX8Y1y3bSTzrYmEDE1ezmy2MuWdz53X57Jq7vHVsHNkjF4LWjeuJzpCp
IQNuJ7jeW1v0Zw8h3dcHOkCfN8PwBKlhkXn1Vo6hSXQHI3Vqr2e9YuTZ7Wrto11s
uieeYxnLcucbFq8XY0uhqcK6RUKy3bxKrATPwf24qkqhPr45HdyZpdlEqa0BvPP1
Wa49ev2rwlg/RzboHRkxGcrqpL2WWWX/Zv/1GfFX7tOhbk2QsAJ1FbuXUN+sFI6n
YC+IWxkFp429pTwVQG0D+371QAEoNq7XePl0ZF3Ck7u16VLpR0+k+BTt57INMUUD
LR9oBlWFgM97poNVDdYFMZngL1Ax4UFajUl4icpcwtd6ThTyHpogLsir/IXartfL
GN+S5TLX29jul6vz4ujJrSKOYNl7ScsT3m1PqX0jfd1XH7rBzmtlzxAhKwdLonq9
RgIzA4uUKGimbJU6px2vPDmw/lxO33tiJsHow1t57g2+uVmlY+IZw41AHPdk8Xiz
qPyOc/ryxE4ZFH5w684iNJG6gC6LshdTEwGIkjfFTC83VRUYNI1R0qe9e/Nnk7eh
vW5eWS4JOn891DegxGPdSZyh9utbi3cziom48RCotq8x/AntajKCRRynqcXPHxEY
rsx69qCoY22hb9OSr07UED8+lmymK2uETBCTEf3kD4o7JjiN7iYcu3/rMGefNWS9
AHbJFaW7Yaaj8rRQHp0OjBqSriYhFMYINi9nGQ0zENqjNj83//sHTIXrlwkajRzQ
EeBjmiAQk5b0/4DlE61AJ+a8DVe6pCC3x10b/ro9ToH9+FQyADLn8DATAM92gUaq
NydKDCYCY+SqWpyHZDQoC1wpDkdo5kBTTVX4BtwwaF/0aifRylFy7gkBDr8YOCKD
8qH9x7nn7lHTXFrkz7Q1Ezmi/GgGETEg0ud5lsywZ6j2HZ3sZVeejGckJ16iju8d
JDlmg6HfL6uNOynmseca8aj/TMdSmPo94QP/hOQ15EM5Ow/l8QVuuCTWlhM3Qfkf
jZkBZWLSgUKlazX621Eti7xT16lcSrJpL/7z3T5lSUEyxpJcui6V+A8PMN5T2Y42
ctxbv0Cx8GifCMBT5DUdnKCHj4IjLTnHCK3U8RxzJZWg4FsOmkJx5bygK/l3qB0b
2xCGVgO/2ergxyEp+usDojwQsf7Zb6eqHpvJgg4V/2YXxoAh3BQ8qexwrvMiHk3u
VT8JRlDIFvOmNWBZCPUdcl4vsQN4bFYgmzt0g93pnseV2i/NC4s1gS5IzurdSbYg
GORZ7QcWKqnAOlVEKwW8kY/3/3cH6NVGiUwNUU1imxPeUtIsHbCYCAWKszzKTl1a
9Qt/BkOWj+js+nRhInVIXcN7451sw7JT1EL332PNt5+yax+6jK72w2mNhrTjSZ9q
Qw3oTsN6yMIKovF5RwBbt2CA/GAUnuswM2yGNW8XGMk8UQ4phoYNuzSKrAN87soh
bnVXdP/XLIbQjcVj1Qwpmi/BVpbB+V448xSOtPQa/NhhU6FXiOStYVGIHS8tZTBn
BHhf3SFJZuY25VoRT5cdrJE05t6OgiXQduE24XQJ0Txm4fSxiCj+qFbOzpETtZIA
Z1VijL/SxkHPK/OOz/siIiZqpeTJU6j0BIKJALU95EFLe/Z08AXx15eOgUetBvO1
ezKogakA6as8GgCXUZ+NLKKVjuHo2Tx5ah5nSazioiv8vsXM56apMFzUAfRvWqk3
xqvNM4j38MJMZfEnnkZuiLXulb/vK0t1CUIkNbKm6W5PsPRs+8y1CeSHaxlICe2q
k/FhhJ7esSZ9hAspM08UQfUJBuJYUNbn218b9Wj/8wjqqQr/Wn6Pe3QWEWj0N7UG
PnglzPIv7qhLQriyMEhShOkaWud2XbeastBDVlZCBtVsiEcAsapENejvFvIxAQhI
XVFK+bCebsWkjGaQcxq8sDyBVf6B3RSZVyq0Zk4P3PQC/mo3DDroiMMVAPt2fD0P
JISxAvKsWySE3WxlGqmdrkjFSuI9n02Yb9/hkG96Cy10igaJAF8zA4GtmI/bUvdo
FhV3xRiRs34n5isoG7jEWbfC/Ttfi1GL1RbTi/jEnbIldFYuhMFMjtCmUTwWH7Vr
lV8RsHYWF3oH7kWkKjZ9Jz63aSS4bnmIxKqF0kcuaWIIdjIBVUdg21fVa0dCBKPS
Idd5XLdOB4TyFMjSWMaH/fk5aUyXdw1dgU29xcx4crNFZI7aXflpyZJFw+QvVyY6
iy1UNrl2sBN67SFkBaOHy0qtsRYYT6zUeW7bkM95LPAiLNl4gW95kOGP/8nBRnHf
e76W88hOZ8QUYVBq+ijsFfJE/sPg06Ip3QKqy3pLCZshB80zYuHhD99P+6EmS4IV
KnVpVBrm85RMZJXYuHDvOla4tzWS59fLv+5h/E/s1216L1sD61/qdq2i8c1mo04i
hst/OV5OzkNgN9OyRPAnIJBu1nZEQN8o7qmCi/1g556PGUKYCetGbUIuxfzsmynf
y4hiQW1dZnJUxKFJDgq5ILRcFuxOJnyVU2FRF8HenUr2J+AuabzyZ41ZfU0AxrIV
A4FGkROrJA2qOKfBqN5+y/pH/5H2TMaeYP1ZlBobMMwuTDwGHfMnk+4D4v6EFMWx
wyPXBDeaCP06goAXlugziCQrNQyRBP1eRlq8rS345TDxdtqLLv2DkoqTeZmGgwVX
Yp3U2k4bw3R+9/f9+7WWVZCTIsuxHacaPCtc98jz99Bxjkfq8e3f6c2zl3gX0vOl
7Fn4U7iCmdQB5uxXunodBRaDv5it6gaDh1cebmqkNWycoxyR7NLyC61rdsQq0OGz
WCM/q2MKwNQKeYbh1vjv5ZVfvCB0hW3Z7D/oDZjyeWAMDvxjh01gVGR+i7Wa/5I9
eGTay0bn9D970WVLdMWy9Fd/BWJyHgiRj7bUOdG8FaD2cBkakvuMlxf/wdbp7eFW
a3pMfFkdptmTTUNRJ6Py8rHPQtEs+9iiUmBjDigs2wz8VVYUmuCIndhfA++d7OdY
bkoBD5002mcN0j7Ahlp8Pj+ynggTia9OxnpMcVuMROFC1++1jILBoRmPby3xjSCr
KSrv5G14wQNq6Sf6mZM/gxGzQuIRyHM3BqgRpiIhkyLocxC2FjxltGatMJow3Pe0
5UEoISPCFh0OpCuHY3Yg2zhZi6n/yhAKpKa9OSr4e+cSfgaOHGb++RyT2t400gCY
SKjrXlru21a4uQ3X39E3moMElLh+d9fT0a+/yXRtOW/4txP3OVygkiYkEaudWeX5
h60ZGgv9+6bd2k2b6DVpKwEgWzOv1PtDTm2gUOrl2i1MitjJskwGJSLZAUkcube2
GBVDFTaMZDU5cFW2B9nBq3g9gOhE+0dyuC2ao9KhfaOfcf+VGVW2FJcLR6hTjYkS
eA+vzf+hCAUN/XCMBP4db5qT6pnxPcnWE6i0ltfcOBwvcRXhkLFyE9z2CYc1bIUj
cLLpQhPQIzgscCnPcZsohE+b2brOmRCAulNwlcNdtqHph5l+gUUP2FaYkoNFp2Le
AkY7Rkb0JOOkue8/fIWPbdB15B18EBv0HQDlc0PokxNhk6STBFoIGSZTFopx9XZn
k61VtwumPYRDtlotGNBMLsl+9k1OeuHjtkvvEsXB0yBwCyb+YNETy7PTNkrpH0bO
Pf45e0NbfOKfPeQpd+ZNEKlZLcriqs8NbjlEM17fDlYQpc9OMrDuyMRJpTt/cn0M
yUlby+SfGXqSC0JIG8DtPPB4eg9NrHMxXbrFXLbbDYcDgWIfcUG2ekdIXu27a5kj
KChV0e1cG/8ip8B2THLfZAQ3Y9bOWpLvcyVPe2vtDk+2BGGiIa+s1uXA/WGRG41Q
koeT9rLkjadgQJAAGtPB9YeCITatyPTSNt844r3nfoggxjWEQb/8yXB2fRKIA/1P
Rne9pvI/tKkF8Cd0wsfa6V+eWzClBqKp/ZpDZfvGJu3VcTgWU25/f9P9OI5HR8WB
pQE9f7OqsRPNnALakZzVqCwDSvSlCAtuAblWhZ/kcc1wyFpZXiTCoj4yMRXiPey0
/muv5jETixwhxtsMSr0H0kC706D6nmzdNkqmmByQ/qgOevoGXb8M5ItiD4XJMfNV
idx7XrxjXs2J+i2I0Jo9eH7nkiEBYC/f+5Z2gpO1ZvXeFwTKU4E12Vp/WdA0S39g
5G3RKAF1gR/20VpvmDgV3s4OIdJwLhMIy1ZZQuOJ/xkTY869FvORWIfgGCVYEQVk
1G7TngcM2JDUipQ1imevKl7w5BL9WbQ6DscR4NGRNb1e8DDfDnIdVZ2dzSIK623S
/zbSysb0hLjoIaDB1OXc5P79rU6NmxNwRIFx4C5mJPc6TZq4vFqESqEkp9QsR5Hb
GlIu6FQbAs2vsdWRMozq4yhepoLIkQ5dY+dSOCvRBo2ZaEiMFoIKd2B6QaBLnnCL
JpreJT3avlTNMxt283c/9dW/YctUz9pCOzAJsuG/zCM8R8KsPImJlVvYlKl5Kz0p
koTJauBlfKW2wBDdTMyQFzblkq37vOQ2rn42yGM3qXhMMx/Yt2Rj03D+64s7rfk1
I1icc4zAYl+sANbyD0DsYOn1rHpWA6UJUmvg7zLiAzN6yqImDJU6kSqPF8CSsOpK
ayTrzQR9Lnsu8U5crR3d+f5O3IN2uIfUm0Noch89HrhBJvL8T4yVljTDk6TL99+V
lDdaYFvHmGAf2X8cftt+8s2uB0ugKy/yux2146vFpO81ayYCo4IknDdVtxWWbZTO
4YqVBEBr7fXUUghQKSavllC34uC4pLmveox3jPdpr86CVTq45YDINDXTwno5jbvG
vApXE7qLtyCh6+8Z44yndQsfezT25Rbi7+yaIJOlJYM2hc8tYUPCKQiMNQ2OHjFL
s+OLNXhOQGCFp2lFA0h63IdLhHGnk9SfWS8+uMOJBHPJv5cwx77TMLRFI6ez5x4C
s/x96pe5QVJc2Qx5tsWj0Mr8lpMlo0SMY2d8pukR1FALd3iziBKvii4nI64tpVoh
GICFDR5ILgUz153sZDIo64Enb0+9Rm7d7ZC3mj2Q1zBALepr5AIvIBrYlZZ53hzP
f7fA6SD97VTE7BAWNr9+4sSTGT1IMGOxSXCO6GhrmgRS8pjPptzoXgrUMwGnjlwG
+MG/C8358Qt0qsl0cE0Wt3/dOUlqjUAUjr8/e0eH/QChGLAetJD3FSxyOGBKuHwT
Kluv+Fwgp+LaJJXlVQs97VHow0rAvM3SfOty+hGTHat2ez9r1Tskhs7emiBgZZj7
JWRsk/2Ta2XNYyh85huntt9L1DLkcEjKzgz5ZdB7mHXTJ2Dagttjr9oy3SLCkSzW
rv8hwxcukVe6xdUcCtabXvpz1LBN+kX7RCbAAjdMMD6F3WSnhb80BmWDF6yDr+r1
dhN++7ykwtaXO6B6TML5CrEMoXhnJ6QfKoA9plnxofS2DNRS6eJ/WCobkmA1YP/P
yLG/HmQg71a6aVtga/PF50pNLfUADir+fAL7qrD6ZK0B7wajg4Oktkf2ecC4IdJQ
6yjEthgFCHji7DMQjjf6bQdE2ZrHorrMQb+02H//e7sZ/5k6/VGZj0S27yFoBvMP
5OE39yDAO4/Ss1REpo7YUXqou6hr0RyajF1aEGNb3M5Akwvkmj6QBmb4IeI/Gwfn
AiT71F2ipWBht1/YzyWz087VObO3BG95Kqqow5kCsOVtiUOCstjgjMyNhe8AdIrO
EsE+eKHG0B+0XwUpxxFfsCxCP9WFTQHYohu/tCpZwWOzdobtf/G7oSSs0rS4csSR
/N4JFfvHyk+lwLOXgKHBPpyK7sglWXCVCiwtbMTYqrXsPERcRXLEZ6Pn4SRodNtw
0Vk9RymeqvIz49wMHV1B98BLQ7bxKayYdkvp1g5fGKzd+/1bsH72WZ5r1K6c32em
Bf4Hfz2o0/GvcZtbou0Jfci7ncr+th7RFIynoQoPsEIS7+HaNVMSPdmpUEs2ydlU
Jn5qgUsjj1w7hqqInXsr1DST3hwwXEdR8/DwrKjPgcCrGkJo/eJDQirHgdime+q+
Ygwvfm91CzqQ8e3U7o3BYyh4463F2m/wYIHBXVZ0eqG7gFIYGqduN5NZ259+69uO
ZVwkhHTp/rLRFiHMmTve56PMi9JaP1YQE+PMkEAPBQmMZoAPpVh6lRU+x1wL1M/s
onC24c37Ti6v/eO4FeFy3UyteeFdgntZAwpAmkhg/jForL6vV6obU8YNGcNCqQCs
Mxv91OjIlmLhUEMJxIzpBVIrx3Iria0x+6uar0QJhwipFCIKrcDeHtmQPvMyYUe2
MtH6+XZ5yPlDv902gFXjx34rmPWrRCC0YCi9q1vZGRh6KCO++KuiDNviVJUCh3Wr
ynEaaCC2wX3x7kmQzbtILqnonpX3qSeE0X0M6m1wgEFlHyGPQQhH8Srr0tPObnSz
B4edXew6O7ZHTEdSx1ZtRGLRLqXRDaaXu27ViA4TqgvbSu3Sd7INGiDs6+Wjth1R
pANl+oaxBgRNP04NTkw94w7rHeLZzVKw2wZq+z79XZhHiWlyF8BnzXIPfi6HtEEw
6dAv1hHwc6PKQfddxXtOKAVAgcQqj+LTEnRVxSSmQIVxjzQDHgsbwZUll9b5XFxn
757jb87Mppwg/1iVBK9vKUBZS3vum66PZbCr9V0iD584LuXkmhFT05lDRih0kyXt
xJVYsiN1Lhm7hkjxLK+ATawbOibXjeFpCVmPUrSeUQq/yH4ieX3NhA1dAsBJYr51
daUQMzTHpWGTNjEj2sajfGMAl41UkZ4TjKZh8vHS1hvHmfSGfjx4odDYvVxMpJxV
hyzPDbZlvCF/RiDxICNfKsdrzTcJBAa2tMLyQK/r/jMu/cow2ZEYYkgFn+VHvzTp
Z9sKe0fB4D1wg0zmyU0cEmEKVs+XH5I2ISnwBvLpU6viaUf4e6qQulo99NpoO6i2
Y1aO43n5ZowNRuzpG4XdcRxjjKBKv186vGId9DbLp5+FTZcbx4ov00ngCB4C/AOo
NFlXDXYSBFLPoc67nckq2T2vF8U//k7KIkeCQ0V4v2+iFOi25aw3tlsFbFzAV+kf
xI417WlOBTp69C/0at4S+im25ed4viXUxVmhls+KyDdWQocyA4nTqVl31S98NRki
vXM8aMiROCCBVxJvLiCbN3pzfWJW5g6sP7ZmM1LbvqzLRVbQo+D66ZIj/tiT/2EE
zvEB0dKBiU4jgSoJ1EmuOfrOfwG1KTsYet2+DFriy8ABoU8takDYFFjUS/1xHNGp
Rfb9LeitLi1sLx2kagZGP38aVAebI2nHFzxlYBPUPP2IShavdNcyRJHs81n0LSim
UJqS42H0qivC2PQMTF/5m/F00Kqn1VpxechxHEevmu5i8ttkxKA7XPLENpGK6B9w
DmagfTpOejKwPTNYBcKhgkPTEZv+jd6FqRcvBcohZ6uRV+xQcMYGWThXREvgyXqt
zhphm24CwTJrZQ1tN+CQP0Xq2ujjncOmqewaNz7r7fVvIGXhaz5pjta3pXMTxQsX
0Yf0htUMb+mdjZiTVBNGUkqDQ1u5Chz+r8psJ60TvkMZZiArvTNnQNYjOvNLASb4
c+sKKgZHEfigStYEsls6Vqgd3oG/it0khdKpTNzWRm0BAO/UbnyxV6oovw604aqQ
UCNj8b3MnJ3U568UHVoXdqxcFRIHYqGuJIAOkivErW01b80vL3Q/6tneFFoNdhm4
NGNRrc43DmqM2+ofn3AKSaImw34xTpX3ebAckIi8kzfgdvaFTQi481J/Tr5CyPpV
baSivKtlu4LjYrq7wy6DOVcZlud4dzreg/uezX03bA0AmlNItF5YWWc+l+oNEYjT
Ia/qjb8owb39g5iSmA20zkz9Z8jMmunp2Gp/0arFqCPkylYh9PyEm5PfNIacIh60
NnaoHqT11bREFfd8J9wJuf67GeXtOQ3ooMqJ2/NGXeT9VVOk4rQcP876yChN7bIS
7GzfT/zeU/5CnxwI0imjiLwUBogkdCGANYEi4nOHWOog6X7w8XgDpWi66GERkydU
AIb7vYLhy03PNArclk7fbuh5+CICtfGfBoPva25Ki4ufYG5PMTZcl8KlV3sAJZJr
Ctv+vGXsAIRekCcpjvrmxJjP6N6dHAr+/E0PDWk3jJxTtqaC2hWX/rkkPOJin8lt
rMpaw0eZzNeCXT+3D+5NOoHRtmn4KrxlKjfu98iBYUaN/HY32mliK6M3jcvEfXsp
2Ba2PSvBi+gM3z8r3aDex56dtluSXL1K9N7bHXzKQJXM0q6Dqtc+rN3H77wpPg/u
FtEDXf5Xagq7PQeTxWiIk/dgg7SHqQGXLALI0wsnecI+5aVDJ9paJGArS5fmD10N
gtRoCofBPW4NSzQfdC4/gEpXAvTDPtLkEWZOIUsSW6wQE/xSHybawmQ3+TyraDH0
16vMuJ2dp9AlrY7XrZKIf2dQI5Qg3pGrNhGtxQMSp8Mg1byXyeR7MoPy6R3xPJ+o
bGoSxTK031AEgDZj0gtxjSTX29KOobFNCtyaP1w8kwe/LM727Wg3gA2hLflBNinE
Oz3rsFdu5Xayhtse+DRl7FpoM0293XKmRNn5/f/Vk2mSA1Bggl/m6I8wsElHE3qb
76bzcdcyevb75WSCLFSAH8a602KQ+KdMeJdhehbyu6GuzXMjphu/IGHv1ncik8iM
UOYPg0F/0ra3wPSSjKlToRmg9Y1aY5LdYDw9Iz4qSBmlpnhG6iEA9fkBUT4ygifp
dlNdHgSsUpW/93bSzCs25eue0QBr7LrKSXy+7dy5WkvN4iNJcoXkEFuzN1DCdWFe
jnWT3bizUqm9LKOTn9vjzKCKiKo0y+9ZYCTcEgRgyna7RNnQCCOY0qci3BQHtAUJ
wL0nAqLeIgHKyHME2+zuAXFJWGHfsFy7j3HASqsRtugBDYHQUw3VT0zl/W+H8ASx
toRuCTzAn3iObfn2/iij1Q43nRCNk585CS4uExVFEW7V8KDKbwnSm47jMPfT+NIF
ysAavMpoKsyKAa5slDQHKmU+/Qs0ZOWpPGvbDwmyjkrGPO5bHN9YkFlD2ZsavOhh
yBhpuPS5n5lv9q6A6qR0Qo3A6Zyp1u1VBWLoaz5cYWlKKN33480YwuOLChun7gvv
201zseH4Xm5uuI4LBSuLLJixvHHBw9W3cRXJ0YTw5P8cvCe5nux9Lm6oyGGbBrg2
ljIVOFEeX2ytcv1EHHgCR8fIfSR5cvvTH+bQ4VMqOFaOEamSHPL37NWud+HQBRc8
FZNYH8cl409lO3zDM2x4SN7h75TJaOyP3rpMbRvCNAPzXWM5YOrLHwnXiUCSc+JC
hqaSToNGLtvPhwkWtc/dS0bprT4mQm9hrZ5QG8MRl41qlXV8tVZTE/VS+oY7OLrc
6ha1k4rn0e+DODGm9U8BV0hnr7sQd+R3vqsPFUDUfYBEWWx5e3I1dSyJG5mYA2MF
t57aA98zNBZ+mOosyPyLEp4kxCSAVqv2cwFXD5IWDBJG7re8OtvL5uI5K9L/likD
/kZo9auZGLM9XiXMcx/gdTu4bCsmcNPUJovCcC3LdcmfSfPwMX530Q/S9OPUPzq6
xEK52VFW8hfmNj0vSCbSpQpUH3W45kqeCU0jgZzbF1s5KfHhOMPJsbMW6ZQ3jTV7
fqtiE5Gh4zeScfm2IJFFc36XDQexF56Q1OMDr2R39AKcyAb0NLjVWHIa/DiUbasW
AYf9RQyspXfKoF0g1z0z4e8pLzhvWFV13L4GGmym+gKFQX+QYaWXfjXnkbrAUKjN
Cu6x2La9frmM5t8jNr6H6a5Qr8b0s9X24s5V3di3RlNqf1uP+urzV7hqEwKuyxD+
zX7JlMLTtTLNjbxgqr2lw77R61u75YZU3j7o3Gs1fOYlU1HiCAQwNVs8Z8WftX10
ESndY1h2pImS2KJdYwz7E45aOCSMzIo0AYLiWuOzsa8weLOomb+XB016tI4MvduK
fnBQ8toRT8AQaRJwYcx/VWUmB95aGdUEITiQCa9DnH5bBfOSwE1ppqJ4EcfPrUoX
h+IPVJp1Rq7heC1Icsat/cYqoKuFfWskxMyxmyNgZQ+iUiXVVL+Pl+JgzCQCniOr
dUJQEvQlgHhWTx9XvzOC7shBYn4K+o0/58vEKJ8EOAaeFzbGk6YLq8Y3QmC0+Fm4
wx9r0mgEil2ljRP8OZ9N4AZ6/z68Q+TY0xAfm4YkHIeo7sgkVVn/uKPhHr5iPdNp
OKSeGfL6wjotTq09uLGw+RO+bfqeHmAQLpjUF/DoqhChD5QlzrpAMYKtPHE0XSAD
3/YylFtdJNV8wI/TnYjUz35m7aKKKxvUZrRG2X+ZxvtbdVgvxIZgaaQWWmcUUXZV
byqDvFIktXtlUDuHzMha8LHZ12dOZOjY/zGRYeV5+kItN7bWGPLcXVQxlcGcdT05
rc90F5DLVH2qyJsbSzXckJRrrBSv+I30yCPEH0tv2lZjwJvzZC9V/jJ9S4VfvQQM
CWfAIhBEemtlj6Ps4Pkr9ZYz1LwLIf6lUi0STh8bu0oeA9qsieNYcqNanARhtzgC
R0woufLaGok7Z1y3D54Abnk0JvMfA+97tDqvhjk1ep9EEr3cZ6bGjpg4O0Uf1OKN
QmPk4pLaU+xX54FRN4ImeooTRodeWTfbuuguoJ5+X+3HH3n4LUv8naQNiqaPcvB6
7akp/w1BmBAJNnP5jaqyEDRFNshqq8DF7Xv6L9+6aHckG5IUlt4IIAB10PsfVopJ
XO89MbvhH5gapo8vch65x4Wr+1fqVGq27Cri4YV4WoRYjRF8KEmkfofGr6Ltr081
2ImuDgouLvDl0tdJIXRwU2sz6Cg8I0mFXjdtw9W2pOAPIaw9fP6ZdMELxn8uHlcF
zs66SYg9Ehw4clYGwSW+VW9wa6v47ARVnTkvQFpmgdan6mXzJ9ms6Yg7Tfs+vhC8
XeyeI435yvJvbO3NEqF+eyTJmefRUBMYdzhsfET3mDaDIFwnFyyyc+3pf4hUudw6
tLbl2MzJjlL70I77+lgDuk/iM8BECpFf+2k3k2k4FUKBL+HWvNmSLAmju9GKdxx3
jnWKiqy8Qh/g78MircROSaC/fUuuQy0LyEyklvq95jwIKOK/+VJfcRhjayHuLOry
6m0kX6aD2gXExL3R38mDtE06s9GZaie/kVTycqrZM+CEkKtJYf8lShDpLJAugnkI
JMOBTQSwRgpH59bdjf3MkeaeA1L8wNLjWNYiSYNkmpeaubPGa5drbisRtNKbYE8/
SNQnPPg2e88mZ7R/HDaM6FIbmojN+JXL5qG98ENmpgZMMb9S/kzXe30KwypvOivc
1EofUi6WfIbnGyHT5Hp6uQAWe35EmkfJwNBTYZqnqB+h2//MTf3sPxIEGwMitRGE
vXtXuM+m95te2SMgO7WJiDjL7KLJuBRcDnGE30bvXgwkK24KnXxaG4aSBAFp41aN
23FgRoKoSDXuWOlqn38s7r3w6D4paFRU5yrCGHPk+Pwkwp4O1YRCDi/4rFZhUOAd
RsXiWrGIBHJBWxx1gnOGBlRbi3IXkzGwqExVsLMKgGalg3zVLsPu9b4xSarHQ5Il
RIg/YwMffaXjjjJ42k84ZouO0CAotObc/l7u8lrr4tYaWGLmTrzV4I3jYUzVh9Pb
seZqek4kEPpbn/81qxW1Wrq4675yUyjsJzol7zNdIyk7BDVUqxKPReFibrDh3mrP
/+74hFztNiNnSgdK7hTpXGGMpnaPSvLsl2R49XnFx7YB+2QaDJKMXnp3dLgxlVUb
OPIJGx/qKBLAYDagcdVY0JTka70N+v0GbHeoZhOgRyXJtQVj5LBEEW/F+qByn6AT
qEKtC77zZV30f3aoec9qAat5ubKySuowtN/6G7pIMS8H6ZWz2q6J1WRGvWIfi6Fq
4B13IoGcjg52iEWAlEU9ZcQolHDUTdkwEtS9yGja1DGysFEQ8sRyKHgcf3EL3s2w
Ph9HKZXTuKX7DadVA7hAlMcvBoLZw6KpZCg+QZOf8cRg3G+cO4rsna7r4yHApzIs
/NgZvpyDYZsN9zei07To9Dsx7074yLoQo2ptfnMxxFCeKEPbEFo6wPRVQkJlzV7+
Iz8lnigF/VBuLdeD6w/XcfpuHYR9olnwtbfVRiDsgpOGBEq5zTaUWNX3RGmpt3K6
VE1LHr5PNtaJJl1St+AwoDC7kTZRWl+oDe1+2DcSu3JLyHTA+6hxzS58B7tB2/sB
2VX/zs9f6khbTe2QrcV/6GUR85mrRlM6G/f1/QrV+BOvlF5jvXvlCNjZAi4FRKJI
VsPli/oID4rcyj2e03qnreepppfk23lJaM0WMwjazHqhizgEPSHDQvo2FGffhmib
cnW6O4SsYgvNW+nMXeTqvVlph81Gm8CpCXTpLBO++z/SRnxksFXAKMsgiQ8dVolF
N6uacx7BiudOjzBTsI2gqB8/6kFIc6LOQaTbykZS5svXjaRhg/LooU4RW/r50ymZ
EWXEMYYar8dmNvet9nDhl6hA4B4IhISOkSZQKQmCmwbSa+dY6+rCZL3uNtEbzHM7
HoEZVN7Koy6aBhalLgw+o20q31ogQL8lzpBs+jLFcfnvSXKL+dfnkz62al4nhH6F
w5O6RcU7WJPc/EfR3hlJ4CB8bSL7bTygTHIBOJANfw7tjGM9gC+OCO4cHbdh6a/+
gSR5TwDTPVCtT05d1BXQi6Q04y01ttPvDEdXifl/dGV6/cdkhRO87ruHurqROS+8
mzccPs/XBqVcKKS6PbSHLagAGXMnsTMVmmTqVRIBd9J3h81CjKTh0X84pQ/IozSa
/9NMz54RF2ACYyAFdPDmp0wcExxUWVN4ZwWbPthJTyZ6JHqCg+t93+/j6sA//Wej
3u7pp2aWTSFeXWipZhNlc6ORC5XN67b5vFV7GAI5jmAK0YOOVFCBE87Bjc8LcF1y
U6R2fEzhiGfZ3lFesyvtL3AgtJd/9IyxT5cEeircDQv9A8PduyMqHeFHPqEgIlMJ
Q3jrDiBvYm+kYgl4C17jrv98TsuYyfTZnq2Z6WwbjPsg1zd3lfk2Eioj6u67EbUx
c5zFVcFoLUyjpsPitde08NnYImFcFlY/lB1dYOO9yv+hgYJHzfzWpywynSlVahIS
E7SEIpeFGeorkmUz63mMQZCnp0xdUsAY1eKFWXOHdnXVJil97Cxh6aNA4MseXylL
PF4JpkMiCaSb1Bw6uDG7kzLBUB7MBPrCgmXBsARq0Da1MCQ5ezseNDZEqwneSHta
JHfy22+XYLia9CBU45ccggdukwbTkFP45LpPu+NjnUFtMK1SXKYd3JFbg/zygj+E
f7ZazzhnGbG7QOFfclBK3QJKOCnT2iDJX8h6oN4rKIIcMrhpsHC/TKYiz3eMN/Si
EkRC8a2INt3ZM02v500hxotRvC/2xYk4QsUrG/+mYL2QIU6HYQdf6lwbVE/ZeB08
ntSOXvHLVKEVLZ++4s/jVIKSc37uSxOAay+iD9kdnV7SectmXgEx8cZEiBavS/vU
exIONE3uxNJtr0dUaMYJWzn/bE42L2+WR2rDKk5FIt8yRC+p+6dyPoglsz8eCOvB
FBAhdN5tsRQUVZC2BJ0cPMdADYEo7Ft3+ixFf1ry4lfoXTJwVwj8kUpaYeNyWGWW
ZvH6GrDLylcZF+Ll1RSbnCLeujaUGdbrsSHR7eM0PZmtlbD5pwbkA9GvwVKpFjhM
ALp//i5yv2KNOoG3qBXL3x7eI0f049SvsGKE6FWmelxODPMBuJsihYoOE8gIljCj
HLkPEY3V/cGi3gpXQvDQDdKvAntOZxDwPD+gt0uxyWWSxV9C/KSyquI7DM1sZ1oo
/qcXlZ87unFrbq8S78G0feEvuMpfmDTBnW+YQZmNxAKFQXHjI+ULqkqz0pjxcaMt
UCh6Da6Abo34dbWZJyweQXadYIRXBxLJECOO6L9+E5hRSW0RKYmVJsBGQ6OZByCL
i3ghUYUiL0lUHaNKnlZOpgz2+KO5h30MRsWyFlQ4Jj59vr2O7DVaDuPKi+loKuOZ
aCmFKMTnke2oUjf6hix8twUnhFCUawkly3S7t4sxmO/0j+65ZjhevUohh2pAsDfD
P3sLkfNQ6syGebMH4A3Q537fx/KmA8njLOM+Ebz+gvQfXdZzust2npqOvuUtBJdm
ITM2C3EVC0cVJC5cZUs+fBUuClokpEuSuLoauG2u66Xjc9lHGgm42f4qffFxZPtW
uj4PPLSrrX5ajMVrJfHtZhvcOfqDiU2BKuo+zGQ1qbYxbc6ooxPR9+ZvuWTuJI4r
WyOEYhIDv2SctCj0vVOB8qBx1qCHUB4nQq07MIURhN1CtnexsalNaqQDmtK8z5gi
EzVt0BVRtiSZdqTNH6RV6xBGGgTsfGRvnA4DVtSA9g2Y7pkVISFI9hQ4Zl28aWRH
W100hEMA+ZBnwJ0i6WZBT80asA4jiznQAXucH46k/wtWKt6CKk6LXRPpYqL0wmPP
sm7G2WsmCNkG/2VUkKDd/XEEjCQ8CTqOJjzlwy+w3OWEMGy17FYTRzkh3rHH8pgN
fVIgPvAdeTqLYSipAZw544Tr/Uksl9WqD59lYE290udwWBjRmTYGHFJfBdae1pPG
/R6onNY9D0q7EwEJERGBuu4dG71QUxmskqbgNMzwHjpRiRdxixpPpfbHEfUC6VLY
ZGdz5yhcl/m6oFcrrhYT+5LnL/UbkjEJP2P7Y7XtIIBp0SDwhuwCTWiWdHMo9xuM
BzdD1G59D41EKsnVrKSz481E2Y6oSzEkrD830Wulcu1trWJaaCDj1UUFXZY9ECp1
jzOlbqVqcvqJDtSAuyPTaSqAnnw1PTUla5R9ZITbVzNygAkdKFNG9mK275G5J60H
TsKyNUObfYNCW6vTNt6tEqpNlcwZYPdJyZmQQ8oAEyORb7nP+BxZXg9suOQPlY2s
qFbwxbv7CnxIWwOgefTXOrEBHTqWtDigsD5VZtI0Oy/T9/UyGTguU8xlABDPefh4
0pcstgc4GzDkfQw4g4zYI1ebrwCEedi8sU3jFCwWqm9J6zcxY7u4Eqz0n3F951li
alTmHd/duBw0kTzFk2zlhl+8VWUESeYIBVyOi36WKlSKRwTZjiataHylOYJ46lCw
oHJzCvw43Kp5zFJV9HsBR+cdP3Q6/+pu3zB3YvGfnEtLsAH/+7d/CKvos0UuP1Ds
JD8qlWZ0qLOtbLnAWJDwQ3IUROKL1zHqzldJdMgaNY8mx9/CjyQTcdapeWocy3bL
tRuPajoRG7GTjC/HlX11O81gKv1USFUCq1/Lb86Ndo2hijvkr6qONy7cS+LgfNfP
9C+cGu7A8aGa4Vozli4qg8n44JQ55zn4feQdX+yUsNNUf8en12ZIyd07kWIOLvPD
Npr2lrFparNUexhtIGwsbfORjU9hFvKw03VUjTh5jF6HubWXywiQBWsRI/LsQeYn
MizXq4d2WMdK9F1hNUnVKBnb53SHc4zw5J5E5uN7l/YalQQoXX+kK7+sjDIxArPw
DtTDk6cb/3RDrFhaC0QOtNSDohUFzMOVMsFHirDVXuPkd/uOtkSYD4zEpRUWJavm
8RQGjoo91ewA1qLMast7xxsjGGTKWk3/0geoYeZzst4C7cl77Hq8g09LehstH2e7
zwfLwCEp+vtsRtuhcRhtXl1la6XMWBQdNMppSoWC3JfeoNS9wyE6auhJHTncoSFi
GVduF8hCe4c76TQ2b6FRPgeV5znBRIrQGprw9wiOaoaNhEpAXmBotGd9A3qgsyAr
uAKcWs7eEZ97mW6U7i82GTtUbvWwB5oDcEfMn1+VgAvFg6FJkaqL1Bi7jzpqBMeR
e9mlphhMImtI71gWO/xKV6BnG2dJkY+qmABRhTb3B4Mb0FWM4PAKqmx4gWGdcPcL
VQ2LBTeoNrkQH2HaY9wbArtNnyejH4mVac3bCzlr4um6v9jVG0cn79DJVICrxNTu
pXUCS0pSeCoHc3CTg2ZGiNf7ma63PcPt8hBhuPtoKM0tmaijW7mLVXBqXpkAN/OT
IX67HSfJE5ItfVLxtOkXxWNYo8g4RcfVsJurkt41duAlPxOAhkJyrNHMtHUAvDG1
MSKxamGXTkjsOwsBUlZrxN6+8cbc7DAQAW7SyBiigaxDb6LM8//Q9/LICp/PY+RQ
qLsLUkifQa87LXQbpCbPOo2roFf4KlXyLJM16UmjmY+xqSqTNodPEzEEhDO93bbH
DYaCr/5aYU90r223ULqWtPG549EJY21mb00dJC2HzHDDSgNncSZaNv/Ul31gc/OC
A01zNL+9C+YUukBNSYubfBkVZV7H5jdLiVxZ8tyHSA9JEMHVZV4AfsZkpczSWQde
i5arwrhb8NtTGK20f8++3FTvU8c21lrJs/xxccvpyhtkv/v7GBgr10h/D2BPbqZt
WNNk7Dexx/H/zv/x7vbOW174FEq7Pgva3k0BtFxCK5uYuUToV5f8etvdjZssioSg
WxGyTG3l/0uZSRm224LbViX/K0S7eaQqrdSpaPo93QoYq5WeRExAxNJbRHaZHZ/j
qXMoG6t9BD/E/R3EhEvYPbrMiUu41tOBN/J9JQmSSto10ZnV0O8+nKiMTJ8M9V1Q
DRlGQDZrZEoR131xmowtMcvID/yJmvoFkjBkF+YNDtH9I/vqe+fr5lWJvEo71N0U
RuaL4btN9lBXvTGiHOBCQx5k64LTlP242fTIQlEDpmflxHzQ/+OIDBGO6DM3luGj
LUGlJ3iiZRgCOb7CxEr1A8ffeZknGSP0XF5eUPRC0CHtG6K82Yq0STylvvZKmqoz
lkEebq2gLs1oTkn8fmwWumEgijEA9VSZ0Ny97oxKxJQYqMjHFFVUGTaGSvfW0PBW
yY08qKgchQKAfntEgV95tIQHUnw7FmvBvisJ6iD/rMCgaq4XFyi5lUPcP+kVfRvs
HXw6aMpIMX3qcm2rnNXsVJZveX5VjrjdnRW8IdLmqBQWyeytqHXqPfOjHUfs9u2S
NnOrQKLO3baFS4tmBm2rSWUKfaBCfd7dMdJdzpGzDqDVX1IZ5K/C5gImuhSkkFcb
Jov2MZ00JVmapjPmIklKs6DskuMcP4kypBOvrAus/elkg5YZmkZlwlQE/EvbA/d8
rgc4CtWh7g63eu1dur1h82bIaEKRTPgEc4IAMH+uyDTVReTXcuL+u3SzHdjmy5Kz
BOGQT7hKga3vPxFCWzz+de7Egrv+ilvgj+mlFCcUUmujlt3Dys9haY3QRczKTvtd
GbdG24SuZYLuEYanTal3xNkvnJsrV/P1TXTdwkdi6kxemrK2KdVZyEAcdAtHmMc6
nFYU3Z6Z1Tp/lcUXLGJFIT3M3dqWaAd1v6dnymh+iPBKxeSCPsqI48baz9C0/kxl
e+kl54x5F6qkGzzm50aCW6EI7FIinZr8nc79BnVDrGY5sRarIHgglpDAHVEf3rx9
NqKBXXH5GjfF3TvrPMzBKG1hfvMV892iopVLnX1UwpwE3vppBFQIhzT+PrTvfu8l
nrN3P8tuIrOB3rqA2AM2SrPp0hHWIJwIgaB8nndoKh7ePg6RbEYzawVfYscDrTep
Y6hODzaDx0aEJmepoUiz5CICwtMeW3AZw7NE1dd/WwZZzv/AIEOL2JzDiUo/qjyR
pv1V3N0eBcCcBWapXr7DJQRVg3yDv2tATBGVCno+VLjU2cZE5eo1O18GpfwHGNVp
iR6+fbwuJwcX65Yef4BlB9LsMMFdFfPPcCQewVjgSP+2uvuaGXTMMJb9RSexknTt
9l6IkQ+YovtsYlRapNi1SZGb2qqmOjuRUmK7XtcE4bEOgb7einybGH7cONow4X0W
tCnaWAW69UCCs85AGQ5ARjht+xu+Gdha9/EMLz9vG23ZpyVWDlDmdpAwrioZAP4N
FJ8n3TLKHWKGtYjqzEpHrj9G2c5SVVgEunbhMP2siUa/4ZYI0wF0iZno5EMQe8uz
aV5vNqNK/2SF363PACakNe8Vjb6BQ4d7NYQOQQyKMCgyLyry2BCzi2IJtnOUJ7mm
13Mu3hARKHMThqRSlnGDmJ2kncsc7QYm1DE/vUFrFMmsiC/eV7ZLlCXxwpGyNA/z
/Io0aRaR7oJbiDxZIWFdtx0XD1JOn7JxBzcsUPpOJ1FpE1jwYwjBesfawD8bZMak
ZO8+ufAHcsYSa9EbP9Jw1boa67ZrsKnu/EJjJHHOwzk9YPQseWQUAytiQ/0zyHOi
WqgvZctrBCrZ4Rgw2mXdHMIr1JX2R1202Y7s0R1ArtUv9/Xam3ZoogyNMBu1h8X0
kW5TvRv3yY+FCJU9qo64S+YR/583vImAUM0f/huJ8HQuQ9/DeVqSLUAGpJ6ydnIR
W0PHgM72WmEs1W7qjBcDoQIsvVBCE8tUxnZwqFahngoSG2qeC/t6Lh2lVC4ohFwM
YWkUQ4YdeanV39jKgF++jtA+B4NsWwUe0d3rXQw3/5jdZ9IxJla3cA3FIoJmH46z
plHMcr9Ag4RLAUSBuGspdRXD5OOClOdqlXNZl1VehejIIhk0Z6HwPnKANyKFV25Z
SOkVuvgbPeTPbWbHgpx80Omcexoycf7CdR9e8Wdmi7SMhZgvwcmsOo9VeJJVz+MZ
EWFR43q1wRA2uQbj+g8wq69tPBuvHHdFp6NwK3Cb8kUmsmOWKQwmsvoTvOKNZqWr
d7TPc43fnLzw+JPCm93/D9xh2ZhoOKsHLhLz4qMWyg9qHY0FCkvey2rjuIGvzZ+3
m3Cxen2d85aSwhbX3slLyglAQ6AvEBkwoSHq3ATFRcNg/YZ4I5BEW4K8yooJX+3k
b9X5BCzRCEgCmDf/saZ9nJam59iRJChSI710EUpvqYD9jSCgOaLrxL4hw6G25udL
7FotbnYkNLq9GYs3Wc7khrVlyw6oBJWRO6w/2cNculQSZPNxkLkBL7pbdfIUZyUf
xuiwqbiHfSWV3srPBGaB4Hpms97HWrkA5Y8ny1CjjeNJoBmHNOEvHzpoblaLbv9M
VUnBpSgVP4VFZNihvQ10svtR/YYhG1QsZypXBA5i1x86fUexLGVt3E/3rBEUf6Vr
rBseQx8wYW9W1ACI9crDASpW10kYWGGjvSuDF9AXs5Ng7DmOFdyCIZ317JbGo3Vh
gs3NZ1U9aElYN2ZiadYtdvh7Eg4hhNCEXvJ1w0Q0sPvOM7vTXhGA7nR8ajKULeaG
MLIlDK8CyrmYn151bR3Rf8C/ysb6sj76ecE3hJ2YPJo1n0SM7gRKRrJyV35JnBmj
VSCHtu/ERks/pM1SThOj6TU2E9XWuEpq0KofUSJf1RkqK3It+usisUQhxcbipDDi
t3QoHJdySK6sXg2b7iZd9rBnCjqg0tzVVhIxNDOnAuLtVFfTFyNtcvEZm4yyu9iK
lpsBFt0DOlGfM7Y6hdiuw9byd634jmzpkVVl54OvllWBPV/oUHLcS+iyLZW9y837
wplVYHvt25UzGewxnIXtf2xa5ls3u2HBME0tDnb2kaefVDlwv23h80ifZxqH9TTb
mg1kF4mdSyTZFPr4UbpYX2gvxn5AiGUKDAnQZSZaoiZBAsuSoD85ckb9K6ubNk22
1QNdaOItImRB7/vsBXMvFqBZFlvjmGuwtmW0mKehY8hXh5RZCqFwhjL1NT5q1bcl
QHQlcfdrtGd7ROVSc2ot5C0/l22FdzBU40UD20fhSpkxV/BMBVnNYD4M4vDk3hQ+
gm+eLPrwliBQMjgj5AU3993lkJ21J9qus9UC9TOYAUCOrxF7iHKYfp5Ho32afton
e9zPKPf36LC3KPXykzkWvf49HO32sbMYGSDLQWCfyzU4CfbqbFXZtyVdYgwkoAaR
VHOKo9nSvftzvJwu//H9CKeOvF8OmNyUvCk887Xq1S630EiXIxUwFaano1YxdHlY
WQ33DcnMWKMqfPd+QUcdRsXjYi4LKGHKSMQXcXmKJJExfXlLOuyuG5VxQ+QXSWa8
9k31p0H80h9HKK+16J3gzzH75ZErAKRn0JPbVFujEPQwUlaNfqdx4BUvWF2IxyGO
V5jULHFuGE7v+tauDhhVF664PtOEtVL2SrgHyld852ZVZdOFa3RWD6SMm9Mxbg/2
If/wOsyOqRnNM2jrfKVsTs/WSK0YUVcGh/WxLDUAxlgfvdi/4KOYLJlpfu6hhWP8
f9oqQsRQbD+nocnkcgbPOyE82+cpI3M89RZhjRjiFUgKwETk5zR9AeEjxbwVoqtM
Spy9gm78UKuaPh1HwHC+0sJdVvv+uWwIBncOQajZ99Kimq3KxqRxKBl/OGd+x3Bs
wbUd0H2kRWQp5j0zzoI+fb6Us2/BmZbEXXr12atOir1HPomWN92Ed3inMqWpwQ+O
uR4gZCcvOxPqJc5iIFk7YHymJByQ9mU92HnqLfBsi54dHTBJPSIak10Vd183NXXX
gV6Q/I5ku7r9K8Pw8S+4GlmmPcTezggWMK0yKSOyVzy5qQihSQXhdKHAUCRVXbmB
zY5hARzB7IgfD3VKikyiKj8i+vs8+KSo2su8HxekrqCOi79pEwRhtrchxAjnhr/D
GlFkzjWg/62URKb1TJwG1wwNB/W3+1RpGxM1YNmk6uL/9WcAjhemc5NLat3e9JJa
QYEFJv1p6xGj2+q3c5CVj1PRlkTC6bX7BoqYHuQIufYaASy7E5e6NoJkskrSC1Bg
WdySxCsSLHI08T4gQKTRDhAWZ2OTZ2LqdmLlTpcBGpsqHr/1PTV3+OGw560EkJwC
ZqaWn0RQ85yXo75lpM5CQ+m7QD8ivS3viZ0YhbyXXucsjS3Ob1KLl/7vRLLrhtnq
QZmuAvk50tMRw2hCTkfMLc5CzKrJo3YozDE7cibNVH6j56eqtPimjY3wK+levKXm
VDN/s1FF+1+OwdU8fppbjsMXW0sySK7lfniEljsunQ9zeXidvXDMg22Qn1elQBJb
qmTI1KzWChmO1uJs0mZtqoEc2utUEFnP9Ri+cybpIs6tO1VJT5O9KlznDep7W5xx
kwrkxTQ/vo4tdHlOeok0YkdZ0ueo2yWAX9ntb5/qrKS2Qo0n58BVs0LUSKFgyFnC
TbuNfhMuPmwGw5COAq0gpZGrX5WzZA0jvGhF68AqubuRV80nwnlX3wfpo8ZtEpAj
6a7cceNuTCqC89ER2KkZr8zu4cav+isgkFgIydMEyAXREWwHTMi+2NlhbnMUjZXj
P8mm/T0FPiw5O1yXmE0tlBF/q7ntk9lQGDy5qMpxjLXDkuaLFbltoo52tjj0zyMY
VYoBG1zG8l00zi41S/4e5VtPt6XJFY7+K9/wV3B+Deoamy7camCXiLwHBm3UFKtc
PPl9qPo7UGTPBQsoQpMUidctQLPPiCzcExKJ6GNLKG7uSPZs9xNV2SvMsg7HfTiy
SfXKq9RM8xoC+EvFnLqwfJF8CcAvVTPVpoC7rnGl1WICVqjygmRnXLYMZobdUpuu
OYKL5LYVgyqsmPXsRjWshnaEX4a0d2D0o2xLTGr3Ea9StmTvM9kZBx7ZyKHn35pY
7vfggnHonMBNdJ+KFiEJxxcr37gBHeFpAnE9Fs/nyuvKA8D+sPHe3AP68zRbAg+6
2rzpMZStsKjl67TlhT92s0j8Y+CHn+Q4QenGtT3Q+RWeTPjnt6hV5fi6476tU0jx
GpehNlckMTphoqfo1EjVjFNZXUnJGb2NJFWFN7Og08eAafUdbWoEKIyLpEXtzISV
dI4C39n1SN8IlId9c5Nx1StvuT8r26JhmdyuBN3Ucz0o5b+5mTpvXTPHpwafYrew
n9uHNDkpHRhPodvD+cn1OPF/V7lws1tH2EorFTUPoQM6zUVvNhH1deYdJjxGauzY
XnIzWlICUJV04KE/yiZd+virl4FMxZk+dG7Zvfi81M0K2P/qujlaH1xwwEGEQwvY
yAfNJ3aG0bWIi7LEFomEIfVf4/nxiAwNzBFJVxzNjxRK72Qopz/Wa8xX4b+0jdvY
bmvuSiYwe+GMkjnijh0bs8DomsBbkfRcE5HM18UL23dyQ96awfA3JCggkfVEBZmL
Qs1NR+en+rh9KAgzeB/+lpv4LeQyZlyw6USdD0CNh0mUk+6uV3yt8mJM0EKVn5a9
W32+GRpWA7S1xnFZuPdRHm+mh41Hgo949ttXPuEXkV/IsCu2ii31LHPij57tfAM/
ex1v9OAHnT7bmvTQn9e5DdhXGUKQMYIT15QJXPYmnv+FRSZfgYv+vkqJHv4idkK5
RpeT+3Ry6pzgqIkioeLTgmhHnd9p7aTHkluMKGHOvI6bDdxg2OAZKINK09Ty58KN
VPZDuIyX6gYGyg+Ii1OnKhYC/62TyGhiB1X9FT9xzjYZYGk+PBLyjX08LmJ0wGSc
BjDJ8uMMp6OvzaYYB65V6jEdsl1nJ+ZD0Km8N8+ymIJf8cIC+wVP6s+gU+IiBDHp
2fdYL70sfv38IuNGsFrZuBYdSD1gNWXDcE9Aqw4GQNi8xJ42d1LCQxq4uyHlvZYZ
ee70GuPVF2FLooh1NcnLhvbcw0UvEBm65j5RTQk+EOge1a0xehYIuo78AZe9flEt
7oeQlYmHXicYY8WyG6fvhQL4VITTRdh5R3tAgdFm/GdXCrKPzPeHS4kVc4hjntwj
wrD1UgMHG8ifENeQ1vIiJ/wOMIL0WfsOxxxDMAQ5oUXwV3UAxZIbQpWN4CmWVD0Z
ECJq/bmdN3rbKwS0dpC1CoGIDkaw7Hfzp6KVyADqzDwcx/w3F4GlZ0/pBqKv0p/x
7UKPlph4mIAEcuIjh66I/Y12T+TREAgIhuplgJFv0J4V8VgSCfO5eQSPjA9IHdam
5Y0ujE5IrSI93Y3z8N7U/8JZsk0OQDg86v8VSC7Wfj4kTroSM2IQBmFhKjuD2Piy
zaj1iBzluKKPCGzdy1dnIo28wRGnv+6nmWCYYFSoPvt+GtZ3vxdstVB36n5kYSjH
dIRmAyTlLu2mPJinqae9MQO8v4chY7MEvFzjWB4IgdZ3so2Z941hpMuEe7lbqhit
s+XtVFQr8XzBeM2xR+LPC28xS4veGAAc1urtOng0CLUjK91iJiD+KLb2K2lu+Jkq
eC1S7qDcI74kNUA7eAQsWuR0HPGp0tLkt/G+TuBOZzYT2jOuIuUhS1xjr8axBvYd
lZRhDqOaD/n58fJdxjPzoOi7gDKestnPG2/LfBJwlD6EDUAm+ADZhqzoyN8IC7rg
SUF3GUAtLlTZoaxLdCf04LRJhIYiOfzbYmEytdCNAF3diSOYkanWKvGqOYqJAE3c
aSgmcCrjSGws3CfEhyqro4FCpW3PldKnUg+E3n+WI04IBNBMpc2+1wDfVbJgjtpY
+fE7UajjWmi87+iTEPmfkIVwdcBP2VX4RqKJgcs+zaAwueMrSWqfuHB7x2i5HJ1F
DWB7TaD5EW2qs2dNS7/yu5MUqPEKidNUeEui5kNltEJfPSI3CQaNiYsA/l754CjI
XN1UvUXR0HkdPgm7y9zrbSM0NwE8nuXMgcwWwV2t5q2lHwnbmFOK+H5gwdwDTeJq
5oAY6VIIi3pE+daWRLtrUxG0CytIj+Y13Ys4taW6gx3D/L6G/O1SDe+IPExEmvUD
7f1+TxB+/ggVL87nNuqxVz5O7ZrZ+kBLAmUcQrDj2NoEVwZj7lpmhi3EhpTYAc2W
RUHkNuWul5nmSNN7A7iS9sRVgJfwaKFINmpC24nYU60gNlYJWkMKWyvsjBkEgLNp
PhdauoPmr+7OVxnscMv5R7TI+2mZIlZYMfmOgHFbKhLsrOSscDTEKzLZax8JzPWb
CSjosHOcatAkuZ7eOEHumf/0Tv0zhAhR7LuWfe4AeBW7N6UTuilrusc2F6Sm9lgE
UBayjQPNBom4eXpOgsRoymLgw8eMfYJl6R4W1MRrSqzfMHPlZq+OmmfFNP1jOpuz
CmxUT3lRvt8Z1qq1Rd9CIX8M4mCtPKYnqRWrenq4cg11VYAyc7JNzVJb8tagQF7V
X+INNq2n8tMjLVxAjXhVroJYlbK2fxNshiDgMctTlhwCvoNC5/kfVABMXuqxa9Lc
zyZC1A5kTCw5qVdTuJQ5Nv43nQp1Ci4g6kwTA1wWHnHYo/jhENCCNp7mahq6EgxY
5TKKPIMx7C1rCwm5QYpPLQ0bZ/lOdgALusiqR+7YGI6IyTZm3TRPMyU3BcGMWnZt
E3jy4Irb3ATe8YgMXHhvfk4RVy6AbhkffxWYMg30VDE8wA4VPoRQUyKxJF8Q9vzQ
0Tyl3L+y4ZJ6+FeWekj7WaspbwGC3TMEPoXFx07vSaGmIGyifqF2YD4qy8Y00iNI
+CK/bG1To8fL+yfLMHOpAYKbqD560DFNFYWTbC1G6SEnFJ4NKV/PfyYtqwEklmu2
ZmKR8KjV50HBZBaKbQDvbPb/GVPl66uonuHdLjGem46Le9+BtO5eW2mXAg5RoCsg
9aW07PBqMsji+FT68iezl4zAWDlh6PYP0dwXytjjIFSGCICXYlf4zz8SQF5n/Zs1
kthSyCFJ1ISygjqit0tXO5Rft2lIG5KIzqDYy7iGmZBjOKI+JfmudlVUX0WBNkap
ukF62d0IlflaXbolwXZE9odeA+vKUhHmsPumMMk4vgNop9vvy7f/RnBPtES3dd0b
xKNxFf22CobABqYrrbDXKYsBS3P50V1gdigj6sQzEwL6Wb8NkkZcqzc9wPG8FdmW
UsIlEfMKsEGgYJe3fzrdLjXHTmpl9wQMHjPjCiOwF9oU9+RhwSIR3J2qdWisLGoQ
hzlB81+67FcmeqMSdNUTYRg32txIpUVCZNCIVgS0aM6cUCpUjyhGlNW/zk3ojwd4
67IKatAxKJologYUPh5FeAcsJLBts/plQJUs5zMOu0Vi+Q3F8g4p05cCOhL22LKd
f9beuw9OeDQgIZVXG6v7VPBFiQ+paQLvm8sSKl5MvyhSSBt6fw/K0RjHCW3gqDjZ
dB6GEzLYVFxuQYNR4qMtXeevuO2j1toH+4N93OWr+9NhzddoOS0jQ4iciYWpWPoI
ssn5qokJ3Evu2AkQjkWUfkgf5CcEdKgBcluW78ZKujUXWIgsO4IsIx/+RwBcsX0c
1zniUnP9lNWZb9AJsQnRznyQa12RBFxghKaKE0y0sG0yWo1wpjCE9gpa3TsXqoCc
fITMpsrhQ1eV9sfgPdLZTLb3UlI/CYF61tpPhBgVEuVilesoMvwCqBcRkh+/gDQC
qS4BrWugH3qmkhXQ1QS8WQ==
//pragma protect end_data_block
//pragma protect digest_block
yj3AipNdrGVbkyMFW/UZ1KVbq50=
//pragma protect end_digest_block
//pragma protect end_protected


`ifdef SVT_VMM_TECHNOLOGY
  typedef vmm_channel_typed#(svt_axi_slave_transaction) svt_axi_slave_transaction_channel;
  typedef vmm_channel_typed#(svt_axi_slave_transaction) svt_axi_slave_input_port_type;
  `vmm_atomic_gen(svt_axi_slave_transaction, "VMM (Atomic) Generator for svt_axi_slave_transaction data objects")
  `vmm_scenario_gen(svt_axi_slave_transaction, "VMM (Scenario) Generator for svt_axi_slave_transaction data objects")
`endif 


`endif // GUARD_SVT_AXI_SLAVE_TRANSACTION_SV
