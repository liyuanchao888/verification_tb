// =============================================================================
/**
 * Class containing the events for scenario observed in svt_chi_transactions.
 */
`ifndef GUARD_SVT_CHI_SCENARIO_COVERAGE_DATABASE_SV
`define GUARD_SVT_CHI_SCENARIO_COVERAGE_DATABASE_SV

class svt_chi_scenario_coverage_database;

  /** CHI Node Configuration object */
  svt_chi_node_configuration  cfg;

  /** Array of pattern sequences that we wish to match against covered transactions*/
  svt_pattern_sequence  cov_scenario_seq[int];

  /** CHI transaction scenario coverage */
  svt_chi_transaction  xact = null;

  /**
   * When a cov_seq_match is triggered as part of a match, this variable contains
   * a list of the objects (i.e., strongly typed) matching the
   * pattern sequence.
   */
`ifdef SVT_VMM_TECHNOLOGY
  svt_data_queue_iter  cov_seq_iter[int];
`else
  svt_sequence_item_base_queue_iter  cov_seq_iter[int];
`endif

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
A47coDCJauFYdmi909CSscMFt4V9PtH1WfiFzH0DcsqDbn7/9iHz1mfXnJS1EE+4
Qi2ooC/3hsK6wnJMp1tZTzx9VVzyPjCB12oI4cm9J2ek/+rAeY5a1hJTGXcl9PJK
Gmt11CvS1+5faW6s3/V6FkTSFcwAyHI4i9SHsJ2E+dY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 276       )
FH8w3QwaWqch7ZJUHQqHUCMWnA/nTqe4W6mUoh4su8uTIFeu2MLE0AU6Mzj5d7eB
7aX5T9acuMpndztCRFm+LgG+stG0xC9jo3/Mwpu7qwKuU+t0XlbMYhZjXeq/BvkI
ksD2nj0zj14W+9iHgkEQMGxVDmu2z04RISslogEwJwBvv4z4HX7u1Yyk1oI6lyVj
b9z4qk4/werLJzkKDvJwpc5YP1Ng2WHSKDmpWWN9M1zsS5vabbrP00qE66N2lZZu
f8Zp46e667cFBJAsRAfKmnV5HCPihLI6t2PB94Em1KeaSI6c3ZcYfwi9b0qYPNrr
nJMjVxPGJulyKTaIzYUJ5ULJKPXJ9+wZIsoMIt4snqLy6arFpsom2TKZoDNju4Nh
`pragma protect end_protected  

  /**
   * Table 2-9:: Order between Transactions
   * Applicable for only CHI Issue B Specificaiton
   */
  int  order_between_transaction_sequence = -1;

  /**
   * 4.2.3 Write transactions:: CopyBack Transactions
   */
  int  copyback_transaction_sequence = -1;

  /**
   * Retry/Cancel Transaction Sequence
   */
  int  retry_or_cancel_transaction_sequence = -1;

  /**
   * DVM Operation Transaction Sequence
   */
  int  dvm_operation_transaction_sequence = -1;

  /**
   * Exclusive Accesses Transaction Sequence
   */
  int  exclusive_accesses_pair_transaction_sequence = -1;


  // ****************************************************************************
  // Sampling Events
  // ****************************************************************************
  event  order_between_transaction_event;
  event  copyback_transaction_event;
  event  retry_or_cancel_transaction_event;
  event  dvm_operation_transaction_event;
  event  exclusive_accesses_transaction_event;

  `ifdef SVT_CHI_ISSUE_E_ENABLE
    event  memory_tagging_transaction_event;
  `endif


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new svt_chi_scenario_coverage_database instance.
   * @param cfg CHI Node Configuration handle.
  */
  extern function new(svt_chi_node_configuration cfg);

  //----------------------------------------------------------------------------
  /**
   * Method to kick off the dynamic pattern match processes. This forks off one
   * process for each pattern sequence in cov_scenario_seq. This function forks off processes
   * which will stay alive until halted by a the component which initiated the call to
   * this method.
   *
   */
  extern virtual function void activate_dynamic_pattern_match();

  extern virtual function void cover_xact(svt_chi_transaction xact);



endclass

// =============================================================================

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
YQJ35UoTLMLJieTfDGqfAJkR2jMqI3j2rK8Q+Z1gecCigM3tp1g+BS/oVZ8c8yGd
ia90RhDGwB65g+YSXSoAp+5yoRVwdqTKN77j3uK/vV0oGzoHjt18zB1LY7GOTw6Q
SNDVmKZtbhWv57NAcodGGrBEmFcrZ5nWBFPjWHIDpkw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 127840    )
mw7tjsDpj0lI7AkQbGGLZ/dJoSfUqcR1zHfsHV1+S1EeV/1UIYR2rKZTO7RZK/uy
prb9ozAOYFwi14Y37cnTTtNt5kKqQ7gY+k3TyOrsYHPCttBIqj0op2+ba0DsRU4y
xgk5iXpoBJKBnTJ8MJi1Ffs82WQBxJvm5v9QDJkLCrtZOslHhLnYx5zz1kf6rQ8u
DMm8TuWQM42TAZ/PnrkXNGOV4AqXSi6GrgZwWqRArr6oVa96Z0utTn2cturqQeP3
L84BKhHBxMmyutV8L/rqujkXp6a5H2DNFmOGlMjl/28Jx1XuFe3oWMgCDcaZvh/1
PMV90a4/bzVXCynEWXwftD6nM3MX8kGk5XIGSO0T38ylJ/32pONQ84Fpk2FCxN8j
gAw0VPw/jcRGVBBDENL6wCIUfpSDrvxqytfEnfIychM6Sf83ngz0h2vkX5xdUomF
Y1K/ruF3ksjo7RuTGWGmDoY4gzuoWsizC0vZCu0aEhdsF4ShAXuWv94eeaLlRlOE
FcRNzuX2TY+CPCgrjRX2Eh9eOIpgQOfY97vx6MuUoz4wCEb/JOB+8sLke9MiiG0n
MoWHskj0gpUYiiDzmWJ+giUwXnpz1zpH/56PZiAFFpo/9d7KJFEObmh1VYYp6UDP
ZC6HVMyl6dDPV5jlmelV5Dkpq20jzyjkUnqZ54FZ0CTa6NYTbxuHOMfI3tFGNbIO
pMYtZhn6S1NHLJSHFVg2MCrYsIZDsy2LxdjVAeqnliSU9isq53Z+zIMoS7Ix0phh
afarvj7yAwWGtgCT7PiEPCMZv0+pHhVZk01zicmWHw0Qxc0EelFVK3IbyBYJASZS
x+jT40kSG8jEFW1aTlb5esf1k8cktZIUY9pFHMQIERy5GmXxeBZcXGYPBJXfm/Sh
C0KGxfX9QhgzEZVW1bracd8HXfH48vDsH4+ZWUsYx8efWkJwlUOoAolcBIgYLq4w
veX+53gcnTsSZSbN3iZbWHicRJbxe8nri8hiACohDhvQnktFi7ejd1ZqSun5nWxQ
AEmlNeN03CP6AJYKRUSb+Y3xuI19Xz8NuZ8SsV9pkTj5pwPhMS3YIYKBu6tcOjtb
lJzrnxRVoM0UsVxbuR+JjmovWO12LiGCbShPcjHKNHeY3Kv+ukvqrZJl9zZirKxx
FGiG4wCVAp2b0aboo6Ky8PfLOE1BoM/gzEV/5O/Z0qZYYhwoKmGC8Y0WHjSElb8d
b8pDxCJZ6J6Nl93HinsbS1IXRvsJqQbSZzgldddwr/Z6F5sMFfIq4o64MlcZBobq
q+Bx1Xy+LIhuDAMgnCK9K0GKiT8qVGZZEDkUS5lj9kig5QRE/CX+VZGd96EMv+od
PrUwEopIc/pHbW/M8GNI9Us06gGpv50TfVeaSlzULz460nZBS1exwGIXBWIjGI0h
Cl5ORG/sQpXg48kk8Da0D8SDag1jMucskr9Xkf9cngES9ml+0Wl0vJSL66X0s1GR
NjWma7k+gFIEW3vDJesmbN5dMBLUnAfmvvW0NXl+eOmXRcqGuNCKJxzLgm41gICq
D0JGxoKrGKjWx/E7GKuhOaEU+T22kIR/D5HpR2oQXlG6mdh0xNiEKmly5igRJVhw
hAUIVu+3gZhJPPFuSVIHioviLq05WBvv+fHEyYQzs5gxWjwRdHbwg2pIR2KNGUTn
86iMMBvK00xOKjJIN5Jeanr1x4u29N08MTxUfixMWQDUjgzg+u9CcGV3XClXvbMc
AET89YpRDV4qMMoKdGdVKNBZffnEVYHqIicc4nS3cPC9SO59kY9HPBc00+vvPKbx
Rt0YLWe6YIQP7drjqgQe2zFfOkAQmjbX6TKyt/HTeL1/rm7SlYTH+XMd9Pnbnvbg
ZGjF1EagSLToRE8C+wvnyH6MCvVtPtqbfbwIdm2ueL/G0HYiMvw9CWE8+BpX6gRh
jRKztA489B3Rn7AmxCMHQ6JiPFkRRdZI4VkzRisjNSPh7sw0nPNN6Uip26jwA40z
nXV9IEv+vegbRBOJAo1sV/dq99S7vq6w4Q49/jOHfycBESrq1INR1a9V8ElAExgA
CvvGrazXSjT4zr4Kisj9ykIZaJ35TkYdF8eFAtOY3brmSy9GGaI878KVJ8be0Ugc
JMqfKMovsZpc/u5uEeGrVE8PM1LTE9KT5LYxtOEVpXvyAYdHzjaZTn7ZzA4/0xLD
f7pfpElJpGZeb3QhX++21a5YUZmbhQtzHkRyBwDKUxwc2YPF/ytSKn2I5MiOgrI1
I25aiETewb7sifbuWHNXBfHVXj4jSTGTR9ttf+6NBBsBYLaqRV8lVJepVKqNeLiU
ItixG8XZNh8lRRdC/tO65qti/b4BxHVkbEQCUXcL4SvYohF+hszN4Tc342h8sa2q
AGsRTH01Opufj3PtWAQjbhmgJOLqzpbSOpivgaGYSPnbX7nx4VGH/dGywMA2TNS4
xmhDHIoLjNdz2DcmvRjZ2nxzhSBGhySiA2eJ/92uhukTyZaPjT2sn59oU+BKgq+r
nv+EwZDHcoiBq5J5nJibnL+NG2d1RPssqkAKrWR6iEfEgKro14FHqa2MnYIgXaLK
bM0sIhwB3/po9o0Dc6wXsGZZmBaob2G3WlSI+LH9R99GoeJdSHN4whEEL7OzDSbk
c1YnOlBI7jROCg8iiikuGb+Pol/UAcbjPTOiiU4gBLOc7FOlkhqWQpFlfB2jkjZ9
v3zK1FU5qK9pvqhIAVRgGuL3/Wxqbh9fQ55c5HPXPamnsrbiOkfDghHPCiiC2fq1
46pQ1290swlHxSaM3P32C96iO/G3UmGpRQZN90CUMfzrgwUMhpZt4c58++7S4Zqh
YR3XlztJOULZBN/8LgUuDW/AAXzPviJP17++NPOXfHk4VaIvFVim7wGQIKOX9IU7
dR06yV6ZHVukThIqYkIy7bx8nvxELjnIcOOI2ANJ96D8iFl8Gu46LwHQSwvQq4q4
fxbgUI9PY+fZIOREG2kQQM2N1chrSluqwRv1ac+uTwfncSQL+Ipyn+OZAQjSlmGS
+FfiTi5ieqb6+VCXeqmnCc4ZW2rn2SX+ls0hiJCrphP/gSwgqmfDhnuqTyy3peIP
xEiJHTmlK5w0syxWQdNFxvdf56R9v7oZN42As7qDmEvY9KGiyy7LnKFOEyCLA5tG
xdyFMrw+A83PRes4ZrlsfSQj3Y6hRqJk9+fupRzeiBT4qPt/m5pwP2z/BBIDjS1o
gHBkYTXs0dU3qKxAbZL5Yg0UI4pJrcf6vKWiH3tHfPyAkdiiIfLgcKHvhHVp47YK
8RTPBruA/YVCnw17rr+HZMpgxhtgDfo/CoNMkCuH80QZm1xoFzDdIhB8ZulUu90p
rc33xIyU1juSGN6ipoPXWf22iXz2XOGR6eejtV+W/CrKh80bRmrO9fonzRI5xUdE
EVFq2+z0wIog9sHGK7D4SklqrXBPdx1KSRjss5T3M4GXDIer4X0f1M3K8jVlDcC0
hJ/hn4qI9iv2G0WqPY/xBQILZgjYDaC4lGjy4SUjGsNaiSA38biCIUHg1qGbLezK
5e7kd8OsjYOcoawhytAvuxUYgeOFMwKl3nIGAOAZQXMARl4zKpDFQgFlQg2VcLlX
IMi2pPopCwzvidX23HWsiGwtd9D4gdduJbjQkzRjcqtHviTMDQOVAtdM60mf6Px+
ONi9yMEDjtuypBVOj4pjdj9Jt59HEVaWpD9sSK29tmx3EuFAkBRD+MdilYBrXbAl
jxEg5XJxBPm5wbL1dDQcPSfhYLj+P8T8jW/uQ+j34y8eLbyLFYayemM2f5LcvK7K
w/MZyr/6aLXt7TF+5KnbC964JJBrP/9z1QsiLfyQvQnFnH93phaJXe8wJZsSZhHD
IeUoizGDRdc3tZfivo48vKnCLRsI/elW7wnDtgVpusKyH3xjla05zAjuHbNpHYvf
Apz0+5ssA+qLNPl45XLei1oQWNBfM77Zvme9Chfk/+Qra9gh3zqwyzCoFFbQDCfT
gWZm07usoOh7rviUlVF6Uar97aj+hQ9PSj0RXrf/6l9xbW1KJTZkaqkPVDr9CjuQ
99CcwAVNVJJC9axmZBSq5AGqmAhlMcTqfh/gePw/ij8z97kWHRFCWUh9jGUgJZH9
4HJ6RhlGmO+DEzyCBjFCAL+NNpj2+Hwz/+4klZhRZAy4H9gVILVdobsf5RJ90319
mtypvxRjWyhRKHSL3qWQK99QfPbUwKRh6h34zDpHoeLGuYMCzhVBtgGViQJsoMM9
ynRk85+kH8sSzHYeyfZf0ojYoc7sel/txqmcyDSpD1Zgw28HEwVNFK7Z4pdRcWV7
ThYOY1zt7BFeAo8SlfHxlsenKEx3QuVZtWbRaHBYhcxzdto4AzXXCvC7kbx+AfY8
21Z1xkn/3k16bQZNSFVOWxujGd9ga0Uf4Z1s/NAYXiB/sYIKN1gMgA0doa2T0aiQ
3HLfjzNpkvST9bYmHFqB+mcRxucsmPesQYkXLIF/3ayJ1oo99F8wZX9SToYnYY6L
dbh4MfpWjIbPLwL0EitkULVJAEvyaJmwd9LOBFWHqbho+VbyMkYdbaBxeQHp3ne4
BshOSNDcS2WiQtpwCaIrVMN0IRmLRMO+uR1tS7/oeYIB5T8t2/j6mg1bg4PNSb7T
IJTU+OJWcDTDgxVlJ+7kwChd6mxoPaIqPJHHDq2otkhAdpU5uKrF6QpdcZSm6QkK
YPG9ZB4T4Y5AFqP51BMRtaR1UUMilOjeQA+HGMEdF+GB6Otc7EXRm1YRpRPUD7ki
iXgFUaHiZtD0gEH9d/DXDouCumIaD31ac2lAUxDgsOjnIjUuKQ9J7vqCZ4eOgMJk
Psy0ba4+EGULbZyaQV0xwmPzE9KhQk7H8HU0zVmOhLBwjrPmAqGi0ztuyEBk4zEC
ETmNmZ4wsrJDz9H/b+8ucLqdV53t7Xvcj5hlklH1JyAIGG6RA4on+I0tOlwMm5dR
NPi+ojnmxdHi2nefYd+g8NStj5kL+SgVNfRtoKTzuuEyNIahs6LNyelpb2yZ11v1
vgEMwdU99K3GjiyC3Zinl5p300D9RghsNN1hfs2RTyriwSDA4SwccpMbqW9PvHOD
sv/XlnTj7QGH5IarqJEBXw2I+W1U3OgzG2gGQIjuGjKvOKh+TiKJwJ7L0IgEWu1E
f/hQrHH4SLJz2of5Wm1Z/UxcvIy76mR/b+2q3GsxTYM3HHFCvgxW0BxjYz5M+LxP
KnmXAOm6BjwDQpmBWEghLWdfmlfosr1uBNps6bvFJAafEpZGUyEaK6fCmXWDtYiD
/PTkdydO7hC74TJVFtbVT3AooqqY7LIzet6DJ/sZRJbSD5C/rCwo3uOJh3fyzi0m
lbZXgVnDlx73jFtvRG7Lnr7ce5u+zET6ttToags9XH7gxV6S53n16trBldjyp4Xp
6Zr2NCwqkURwjM/Qe1ryi9DKtcNF62Wo2L2qIDkvEvUe47sJ7bYniAzWQVBpBXiG
cAFokIqCvDJDDdVVmcv3xFVq5PG6vI5DfOzbEAlk1JKN5LrUkDQpWmSzCF+dGUH+
Hh7uoopjAEw1xJZTKoFqQyX3qLq3SSmuQ2iLAPMsjcye0YZLi96URTooYUPTK2G3
pU2SH1qPuba6A08n/erKcZiRRSGgSe4fNHPJN8vZm7yFmcrzE6CAcPzY1tFyky5D
RY4YRnKDQH/U5VZGHHcEXYuWe/tJh4e8lUERE+yHiGLLLAZdDxiNTTXGl4UQ7zTd
x+6YOLM7mTtQEzCnpN85KdSyn9sblbIPUdejNWat4uui/63wE+F1LCdBVR7ZZZf6
Fkw4a168tV/LXDnHy83APctBkTq5bG5++XkgHAgiqUeoxTPYO/teUKO3xpT6mLsh
dgXcGhN4cnET2C0IET+khL5uA/jS4v6bSxtGjIIZzTssIi7/XTjcDTimdCKzRgX9
uh1yDp8KbaAS9OkvtendiRcV0ug4G+9H1GS+c+IdyB1EuTTfLVoNYMncTsTBrYXk
NkKK0jkRL1jPmCngzwaBJ1HyafDXk7+DKvj0mJTVjB3AOzMSTsVLx/kVBiCdLjez
UxF2d/45j8I5Il5INWb3+if8hJ3kUwI5Dx/kqywQr5IqPLgcxX4a0Sp/aj4Rg4Nu
cgEB6NXy4N0tGyJyfTC9xuTfjIb7+xbzidauiyVsYtaxsRCnLajy3p8VCZwiESiO
epxgQnF3K3otFUQ1lpmkosjIMy/6Dupup95o/2tQXbBduBkj1g+OFlMxei/Ymk4w
RphnL6/Lz8nehZjYcOvDHgdruQwp6WugfzZXd815IjkWnnyBOCcZNj55yGIfsrKh
EGC0xMO6FrIzfDnAtrfrPNteDFZt0wgg5QKR5hQMRHzK7MlK4aiTLIxmoYla4LxB
UpgKyiThe4qVkGUmaZ3oHKo2EEQH2+U0Y1I6ep7jDdRQl7ImlJ2UmXGzd33guRiS
8S79y7kvJfYk1O7R3kyUABebMl4rpsE8ykg63SEKt88gvmJnrebf0Hnv2sB35Uq4
4xjOzR4s/bnFMACBFVDckDAq9KET2aJx1egIcaBSLPRlPt9bmrwOa+kqb+gh0iRo
E+5MyCsGRPk/RJ2ADEoNN29kGRYDNNOIBsM6eowGGFCSkqIIYvHMtOJSKppZe61N
LCdhJJeezuUQuAF2vvZlhjPT0myzjpY/oiYtw3vpZr2YfxnN+EM/JrseKRowu9lx
3bA1tCYqpaLZEGpGbQH2LQP7ec056G7xIobtIxi/SyYbNzwFGrVLZ6sBR/Kdibvk
72eKaQvJkSQWeZZI4R1GxQRbDBp9qSGC0PgKMttiTAzbG9FAc2Cu5/DWG5Zz8Azs
EgKhr00XVB2grIVH14HV4XKm2pNOw4rxnWA1xH7kkX8p7oC1uY/M23q3HmWJypjJ
r/UNO2IO+IZ8dtO69h0hezumzyYdSmxuAUG2DTQZk9GmTYJsLDjWaB9q0Vt/kRmq
8DXdf/JWt5kTvqIMozAMJXRK3R65SpK6zwGUpLbZGSUbqsmiHZWrb2TSlV0tIydw
NA2pJZT+Xtr0uGT1kbv4HHKjzd2iNVN4bNBaEqkuDoFwU7cfrgmWQk6B5Marm7CW
zyI86WMTjzBunU8dAr3iA0vGXPa/fLrXC8bbuHsrSFbToQ+kd8r8Ea5C57VLjWIB
wefLBuaXrBQv9CUzeCwe7Yw3B7Rf3gwFVwUPpN9RVR7Ok6GhIWjgwFZUFtTyZYBR
+Cz+ohWeEvkVNAhEWGZuMqBz1m8kDvzUNpdRvxUxCt5d0aYjVIlyYE71FrF4DdVE
tyOJuWvanWMLWqxSNwxLChHdTigv4orv6uzrkQ++sLH0vqIVz/80G65lOYuih7Ay
NelTyulQjOfPXI5372LBnhZAlmJctiO4AHMIFagHPY0BBAcYLx1206eZKKy+5ftH
56i/FvyuxPDc5cuOQC2SPIWoSq5C/nAHTMFLtX1LWi3FAN2+MOmgoy9WIcZUrBCx
awVTw4T96hhIjoG2fPmWXlMVYY7vV1WI1hwebY49CstImeUW1lkmvPbWbuExxpfA
8K6b/uFfUFHtI/vNadfJ5mddxwNvsOo5dU72M0OXFwRhILN/1QUS4akawuQ3ES5C
nK5F9AcD3LBgp/0QqQhK8buC3AiM6yKvs18rkH2/6H8OifPv103hOQRz15cnxxNZ
+u0z6dLRI+0eA0dT4P60xmJbKr2ATv1SokvAU5gyl1rVoH+5K3YiQeFpdvUp6OEP
TOqqzqcbI6qGzwtWtOMal+rIrxlNj9fCoObc3cTs36iIvKKn33gl+VdgPrwH76zT
P222l9aqHgMDfI7yd44thAfyj7KQjyohhBRsY24SmPahcXrcAVeGGKr0ksgndd3s
K0MlLV+H1TIgf4KQwOWQxw2BGXPUMYGDImN18kfl+eFqu3HpeZuWyOPfD4h1Avqb
AgC+u1fV5K+t5KI4uJRGI1aaQy8fGD5egRDOh2cRAbpqLAfXencD2R2AyBmaMOjo
oSduriF+J841Iujkk94atN+74ae/XChp4MpilvQy6vktpgg+77tW/Lc0LNU7aZzM
L6qruE45NtTBxxbrGD/bbDoPbIHpXIBgLCh35dv/tUn+hg6w2V3BBfKKQk2VlTgm
TuLrIbZkKi71R0cKwBCQk4d5r37lCFqKtzD0a7khZm+eOctmE2WFRSE2KTl6ari/
mlNAnrDRzYv1lLABxSmDlVMvK41VihQ3LyzVEUZltOd0NRzgEFYRNSx6tc56Y2/g
fumVrjIXOkneP1zRbmX1JIJPw5hEcUYA4kG2ybJl8LAvP0Sudg7HE06JOhPjpOFT
XPu0hw1lklVWrQfimhMGzzCRBCFXk+BbvbzqcfmQEOjH7XdmqFeEoLnuwNaNn19D
mJwZl4sWqGLf0Xo4K34rfaENhKcKYI29tRUp5K7kT4qxfZXsXwC20tQIqfVvnBXp
0Tv0cST0y4gzp1F53LYe6BCwHr7ISt2e38yCUioacsKFoN0/h9441m14S3KcM94T
BmYFTprlmaAT28Cz5hoyo5TgNByqEd6h8EJfYIcFma7KjEhgHZDQLGrOE9gYxqhw
FR47rg9iM4jiYIH4YB7mhnKMl671h9vsKTVFOR5sOLwEpbgIft8hNpmwDnU1kWYb
Mb/Nnz9HafbEBKsL5IMORAAYvxQ6uX7NSNNQe8v2zkG+j3mO1G5oqDtAi1YBAOwa
rtu8txIbVF4l5ujkS+PARqOOkjOpQ2kh97QHkWnaVBp+grlVvE6i+AnxQSsPp6sv
PL5YNsSW2Rwev4yOI+UuYf69f5Jm6/5R0992cKXAwEp8SnCulyue9I45WvV8kI1e
yvpyZl66HPoX16PvJPM/jWYLU4vLXSXlAwmITlFxgeMIlZ4YSFAc38IG1ILENuAM
QTWtfViw0u62Sf6zS0lYATena6BhvHQ8Hy/YKhgRTUEcZtMoESouIokQrY3Ab75S
GVsNnVTf4yeRyHjx619A1QvqGh3QLZu85fUtT132+QGcvcrDuhqQsUrN1S55k4J0
LZMKgrRcAcrMTb+0bMeuf61pNNVlK4rieEPEyuWr3fFuVuus9TASxPyEJKmK3orc
rGCdQ38Os7aHF1AaUfPDJea6lpjgoNwtJ7ey+Rxk5WUT/+9P56WqSiPLLjt7yXke
u7Cltsh0Gtl5pRjtypZ/Nff1rkCl1NQodLoq2ZkjyUhkySUuWJgh2yxa1AA1dx9k
ztPzuEz8USch7Udp8PgQZvYx5f7EoloPCPg93D57dRhUIRoNVBEM3yfZrEFhlGzC
SJk7WUh26dp8WMWMT5daC6/B2wYdXxWcTK6k7ulyTkNYB1IqxqF7NXwxjDhNFka2
J41mo5WWiAhoyg91pD20CEcW7xEVH9G1/D7gCbF/2UbwXLmmw0NGnenilNP0umXz
4MvNj7Ivh2XRoIppsrKHfkp+dLoJgD9wDeHguMyO+iSPDs/xkbarJlta+GBC0JoM
QGKX9Mdm/CHRjivJnmBjvrC6EYRXzyL97NYPytn07KVzl4TYM9wuDacR/8ejl4EL
Hj92vsyAGQOXzNKwAvQ0mhl1KC0PlWSHrxvs6wU7hp5rjEwqg2ib0TrTbZvOSAb5
L6QL7NzqWyrY4OtgtBsc9o/YWZkAtR8rGom4ise83+dFfc1AdyxyqC/F8MoPXMsg
9s+phkp8YNzUnTuOaWvelTXyzZxK7ulf4YS6ydoQvCDb44VnVlPp4a/rtw1wtCpT
qeyzrP253dtKtG18uUt7BWhcwuSNxWHlK3TvNWtQ84Do7ROL4Jn3QRIBPszVkbLS
XmJ9XSZ05pGAfxLLMPrH7pyMKw5JvDh5SQ8T/kQaXH/lP8KqCbxQrebUkKgYj02B
RFJm1YPB4Ea5YWewiN+2h6brb7m8RXYlWs12PYc6s7wHk72BTx6itDV0zF8rOoxP
iEj5RuyZmhblpfxCpI1Sj0IMCY1/jrrkZ4FzPD7yEFn5XZ2VYVWjtzoKOCnQ9viq
1dx+RNoUL8LdBYCc8fvBh9uFmm/+470i+5JfBNihE1u8p9X3086fTO2/q/vdfLPf
A+r2xhTktFReMGD6B8jRCPofzKPTKWAoaXJq3PkJLMHBWPWeanCiSmEk9tVAPhLI
8IB7tcB0yuROjbNwXskWmxbcX3Vp5gHZC4TQCabWYyzJxZE8vRILQ+2aitPhs3vn
u0b9hJaPoNQWC+AI+3UesPlJKggRKWJflFQgk7J089bZxZ8ngGaQpT5S9U/QgQf8
79uiic7+F7TWWZNNZvApk1rhQNG1/wcIyR911Ww6DFa9SMIPyPdEWmldcAd4yRHH
abm1/2+cDLjZZfot9RuwCxLjaTtcBfPBVGJlohvrfgxdPASrFHXZYwgABAQWcWl+
PdB7Pe3rUT6lo6czQyF/xvp5qVaFCS3cj+1O7N+RTYZsLTHT6e94qZqOWCQTpZ3P
Z0SLKz9upDI1IzxuaCF3voz08FmcrO0ETlna8MEqZLJZfCfoJMSfP6g5JvhaEREb
GZsqJiRhRlIqUJeZGmblmW57pvxX07wo+zRP9DAiVjwTCqtF2MxAaH0Mwynd8VKJ
EDPBTjq1ub07hJhHozTn/yI7WUCa7uH2NMP20EqoM7ogZ5NUdCrQdNrFga8w9fOE
uy9KidIGAY6oAPpNZ1nffqiboe0VuD1ADVDIp6NnJfL0U/iuVXnUA8A0+0OrWgWw
dvby62Lxr7l1HWkbkvhBEXcxw21/p056cfGVAzjNYW4C6bDJhRsLEQque4CkuIt4
AxqKvhHt2TEs0TyEYKEpfTon+AYMlnhK7u5i88s1HtJ3tGbNXUfbFnFxt53axBFb
w5i6lnPgHc0kJ8+x6HUUD04h9zsYpx7ZnzAnWcU5zSP94FqfM5XKx8RvL7QWCCXj
/I10sBeHOt+nttbCTnN00yc5DfmlhUtOgs6y2UoQIiAwLE6+6QX5nS4TyqZSOMXg
dMWGLEsECb//sMcnss8qDK5CVwowfAhCDWG1UPDaDMJ0PMOici7T+i8LFRYDtZxo
E4fLempqTwd4c3k+JkhnaPa5oE85Hl4AxGuaxMlhOUja2kdUkyriiXt0Ij1vw5HY
ZkJm/AQRELbdF1xnZvNAb3aPxiTDef9A9vmANRYIu/QQ0/S/j2vL7l1tSpcWzC+P
lvBrHhA6b/YTrFm2vlhXNUEu61UWbKtc2UtU8YTcDc+Jz0cIMFRVxukoRZGS66el
ecut2BG82XC6yoLcGo/kRcdJ2OMrBfuEFQnOUDb3lspDwG8Z1yJiplDuCFbi1ULW
tNM+6B3+LNmIgUd2dsQkbQ92D1XXj0Wkkm7Fn99F71KyBO6xIgH9tLgw98Pw46P6
dNf2rvk5912SmVcTMCfc/7zkNHh2Gbe7U9nGRZEOwdcUlYHXYTuePgvxQsN0B/PT
LY8GgDmLGyYfkf+KmH1KhP7oz9rwhKapfkFrV4nkQh/gs8SV7w3YgzXaSkgNnZSK
CoKF3Vh+dAJjvrhSTlgqGchEenncH73aHj8Jkc/n/5L1tQuDr6GXFDuxB8CqBQcP
uPhxBPiHEPLL5kYw8oVi2u0SgSatCeuHRnyHrm8GE+zTDiJDE+H1ZACzfom6bh3K
jekZOWEb1iG5XOxRdCJJCqxT2hMqgIs5SX81gll9/pLR8v9NsOx0I5Sb/I5NAo6W
R4HghbGbwleXWd5HXm7OpTSXl7iL7pw6LADQa1S/4QixkADOwPFyky5OZnMSgqaX
Rwu/k4zjlvyFrNUVoYqah+FI68rZdoUXfwDuXAyxP1UW+dwhVavSjlYc7WDp7yAm
Zew/oDMUs2YxtWnsziytAJK2XLrDaYTAx5s7OOOC+DM+JtPgdmU8eXQ1YmejEQpf
4VoUqVyEGBQdVk1MY3sM8rXwRlIU2oST3IWMMCZ1tNWyVeHc3yNhxnjoipIxQN+t
cyyjB+tS/Vvel11pIl+uY2xoVx8eInixdrbYZwnbx6fGiEgTsCjMOmcDfm8tpOPU
GnFMOQTjeIqmq1Io3Wq1LRZS0Mqyf39bs+0w9erV6+SdiTFA++UT3tA7mgp+HdfH
RlLNEY682wLG2Ygap8yoigDv/5sp5kiQw3weT/6kvxjRYazIBg0Fz8CZVWegJ82g
dd/bODagB4jet4T5od1a8nHGrAxeOBH+FS1rRxILxlJU+1poQelzD1SBF2Gdfeuy
1Jc5C6Ltq/IWswcjO4Q/Qp9mJAHozvCdnLYt8ktUivJLfRdJgAreyh0W6QSp/MPE
F0H2HKZ9gCBvj5t0gGscSVsbic6rcpDt8Eu44kU7zG27VmvCP3pktI0iiwYsv+AT
JL2KDUPzkYohTIqIy8J3qd6FqPr5dgEPJ5yG/uChd0y4fNRHiwHAvCD8OWQ2ppzC
kAcUq/I7h66s17og9WO5EV5+loLKigdGJRWsH97SXqxj1PQJ/hsKj2ur21wGbmNV
pqUbUaQojTZj99jFEskrxKFjk+OEuv/mX551HDR30pRp7p4PvX/YaREFRx8ARS5p
EdjJJTQSvL5lMqRwS8ot4B6B2Sgks3SPWCuT3VxuYdhQADnDGScUowDYjy+CrmOd
xpnDc33hEgZsIEYk7OYOG1OnThGZBvNGhadgUIy7msvHHhNPQK4blm8IXULqSlox
SR1um1+A5NQ7oguqT4jqaoNpu35mgUXGHbRy/LCiNOVHqxf5/BZfeBg8YR5EvRtK
k20TCdWaoVTk6HMGJl2gZlLw0ubdH6HgHoPoVQg8XXfZQySJK5xAc4pd7tyALecH
v7OIzfK2YL05OkH3wNIR07m34/M1y2yv7X3W4tRj2l7WrWJ0dKYmM/BLyV+1uJOj
mWgyz6519/PZfwQxJpZo7DttYiSBlAaDopknKUGBcckcf/x0yPRQ57PVT14jrbrs
O17f7ulPQ89aEbLz8XeyE39ICafcWONorLJj9pDzFhnoc1TeG295K3+sxJEiPKLM
VQCnkA6gtzsyjEkjm00+Tv/zmIQourpAAee2ReAT2hbdUtBa6ik7b8lYA1uTufYR
MIPTAYY6oZeCmx5F7Pbtta8AvP0Ik7uL0s8ISYmNgKxykMEjbu3OgJW6ZALH3zF+
61iJrjtgbPUz3Dtgd+X36hCKDgCHFZEJW29+a/5cJJ3rhTneak9PEYzTr3M0S50+
X6oOZm/uks8HsbvwdIkev/jWe+7xVrq8NuQq5Kk/1mxtLOgNBiCcSP7f0N+v52HY
6/q+Ia36x2RToMlmUzNvokjQpApi83DxhVVxW1EpwWtWWILWRYryBDqniXuTr3ur
mSKwkTp+uk884Z3zwc6TfugmqdS7672Hcw/XKR9yZextMZg4gslxgCwHF47FdNZ4
6ixd6qvmH0JFmPSvnVZJ4X/jYGj73bSGztWwiNbjEY0UmkUwHrtIRK9Bf/0b98Wh
IkKSE9fZV5Nz5kOD+W4qVa9HadjnYiPUrrwJvCMvULj/cwNjr3ikjhh0Tzeqrlef
3yetC8vI6Br7u5wvpmEt0G7GDaKGWJdhY584yliK7NGuqsdKviZmwTA4phwpDNmY
QYCnhHkLRvYmyRA/Y+oJ/stKU2DrrX6ESiHkyvBFcfC6sRz8k0U1UhkvEJ8iXtce
0LxFofRRKrfyKA4cKa5ZrbuOfE9BOhxVeWruiRKgarSUmO3UaQq5GKXiEdZk8obL
0QrjxHH/1eGvhimL4ZHsl4b3UvbH/BNu8SgYrHwlLIHJM9XKv6KK6PUveM5f7gPD
BZWL1ZXg6Gh/wZZ+sDX2i9hiFmqrnWuy5UM+8oM4yS+P9syOnAV2atDyZO1dVFMZ
oEIe8Zq1AjsT+0xcmK0Wsp0v5R5sXVfLHdx1IeIHBKIKedKG6zFCyhWWFiYKUKdc
M3v7K3f0LBLLBNGM4KugrJcyUZzUbRMZd1GTnvEQhGodS8247mbBbLLG6JRT+klO
KORJiW6OrYrSF6ZyTVO/FHpuY6uGfiGLbm3J11ipH/Zt4xz42O69ZD+7jUSMKiiH
IzJkFxeHHdyHo8RQmm29tsYTsU059ryAPcbjfVlmk4dHEkyI5RTMOmW3wo60zL3w
gCGglm7c356F8eOXzOY327xCSagtf5+6yKx6RsKk6Hj9C4JAXJMMeUIkcawccc73
7Opj3cnDd0f8sgWL3YeiXGRgSlSROvymH68rEYyiIn+vEnwsZXYkJhbm/Jk0sQcd
htZYXZxoQc9u7B/duC8TosQxTePPW9HVhhFmQXjzM+U+/+MUMochCD1wC+yyFUOY
LX4ghfX80V4W+Fs4icQPPezw2z72aEhGKaxzVRbWjkLvc6IG8SEH3mUsX+Fv2EF0
Knk8NkvtPHneVEs1ezn6u3hFi0AEdtFbAfvznWgG7p3SbZOGMoI9myR++gKoa8JU
CWW9X1GhovFCrT2C6BIM6oTEBHqWsa1emNuk/nCVIhmszcvv8CNbxPzaV2+AB0J6
6mnYOo9E8T54M+gRzbzNHxVJcL9fQl4v7TnK+HW75Z9DpP2/lB0aJowQ33YL+pN3
p7mqK74puolt10tfjTpPbK2lygvMUecB79/dX/ZpepVOxc9tW2dFR/OuCKQ9JD+p
PWYtxdEmxPOZteoEmeRWwfv25+SfpaK8mTV4iPxQx/U8y9PNCWo3sEoWF93gvvHl
Wrz9Oowf8iXHzzNrqM8XJhmUeNRt1eY30gy3C68Zld3OkPSckjPVnzfstL76FU0l
19dKpUgxVLfTMD8YNI8drN0YsmTQFdflsmd1yXdv1Yrkale3ckp4bEIZh+Yx9Xlg
LxmWAUM7MNHgHR0600WEOdsIHFEnBwxHK+teZdvEOO3xYsLwBZzlg8rKWedFGVrH
VzF58H6/kVIjuI4u1dQ+AmCsx40IoUjGm4bbYibORBVhDBovfTbj3tTYEEQeSDRs
PzEgNnmP+LvLlm3QSlOBq96IBoRaxz005Pix9Ta+wyfIoCU4+jWLAeaJale7vBIw
7AQsHuPFYuYoFiovTvaWoFz/lwLitgCEu97UOxk60w4TqqX4ApabqtYQ4iTPtlx1
ZAhRi2s9YSR8GeAwMXX9u6rKW+q90xMNwjjTO8HYnn3s1uwv8YS5RruEjjaGdu1u
+zCf0zWHt/TiC8DNOOU/lOySACZzmQzbnmPxgdBV8/UwfFq63wQMm/6YaD6ck892
VOXPwUNJNMhlkcArURi+1lDPDMv/Obm0BmtOWyUJ6alCO9ijTi7k0urX4ObdykCh
7+yw8JjygTLxtPrT3wyXZQUjzYqn+lox5+wK6NVJv3++pgr/bNz2OVNBboDsw/sm
kgTKBgFJQ7PQ70QFd8tX/1z+MPvkjI2QXe2ZS7naJqueiNtF2bW9JmoxSKY3h843
xbpVWpWQxqKJO64xzZRZGNScn6VnwW9svsXPUKkUzQzR/XAzMUkyvyf4ezHmrcZH
lTW+7klrY5iD/Z2T2/g0jsyg4/QdpmA5VfupyLvaz8eNtPZ8zumZXMvc5mX4mMlU
Ik/QZisdCAzfEXF2PyjSeXRhuhc9CX0c7LJbFLvs3yr65SUDxSAW+ylI0w/i1SYf
aEORl71i5yKVX3Wdfl8yyj2l/F9tY/Q/CLAqASu93L/PXV3DL48+c2ssh+va6Q+p
PGKuTrFbxPNEGMJS3HwoZsBhJS+OEIpUgvCmCRw6JFyXaM2ktzYmG3dvdvrMEubR
o36r2+iclZRRgLX7/Lop6Lkg6mT9CIv6IfWjpjUhWUjf3Tq3nkflQ7/VfrBL39yq
kOqJycfiNi3FyTdX+BNABaXRRtppUYRwyuHytXDM80RckZTPkT1XiQ2D/8nSGqiP
BpcQuT5+Uwt/4nMfSOxsifthwdFhYMPKU5oyOvd9bO5QWVLhZgNEUDqvUlWr/tWt
fdNOA9nhk9Bk3sEtmgGEH790NGfJhUewROUibFurqqIwUHNrwND+d8YNTKFaasfe
2T2hSF+VwKgQiHkZxkIsdB+NdieCW6cMYUhTwAll0QiUt09BJUwB8czDvp93EAnm
AtKQWhzSpIzfa2kNsYR9oCjUca0jlm5E8HC26+k3LnIodyFMkkd6kgbwTZHGfXKC
6v4hLq1vQEirva0c/8e2iLZ2eakoD6co/nK1lGipNdcazcIwj1w7/bCXbE8PocAL
SGphwJGTkq3zDmG8oVLmS5rhtEnL7JIlwfeaoKB37Ju5ZfCcc0HA2AKuEbvRY2ys
K7qZVIdn/WCALBPutlBN39TmbgcQIW6ovPphVZurKm194vg3egjMBd66D8RurRKH
R5rPd7FpJsXdNjwfBKBb35UeMwWrCI4hBFltJwJKvLighGRpJZi/PHLV63TYQCQW
zhiTqL3u77AyTFImhaXBsNZaHaWNhI1j6nqeHnbkig7Hij+l48Em/04uLW+ABZWq
gxvsVUdz6oHEuMTFzX5MFwo+O0XIDO6W1tHGF/Vw4NMy2qPej8aQrr+X1Yw9udbx
wjoNv+KKPgWJgQXht++udJE4bL3SbJdUe6oUgx8YpfyybA2tUegGnwnNgWHnQZrC
2JukBmYlOWbqIbwD/RCArZsGCjvVm6+dlXHzogUFXJi6TJErcqqP2V5xSYmHHQSi
UDyZBv1Qu7qYD9eHFR94viwZa+i7b9C+s3RRO74bpZF5RGO76OPPyZPEJAQyk3ea
VJwzcsCjbgtKxDINx3gKmzUkuv7Zq7f+fAoPA9uWijc02TUPFgFYSGlCezSCwED6
+NtBl04GwnMj0VE19BAHfwIBiHiffnXcXhNRcPl+W5OR34AE/IVF3/SC1dPy0f5z
9p9tqFJmH6/k9ym8OIWmst9iPZD2WML50DXogk0R74nqtTRTKRNfbo3WZizd7ft6
hf9zo0YEou/yCEHANXvMivXbuV+9WXP/1l1rsDfzcqF/XMbD1cKZG7e1dVJjNG9v
2TBcA5tOKUdwodb/3G6nq0pqFXHgf50gqXpVGyi58AvI2ZWdBGT50W2adn94lnCu
anM5qNiDZuObLgr/xAX9CI79V1sNHmG/qdjPaGfYcsIhh8uW2Etw0EJyCOAjRIiJ
s9evYet341PF+XE0VxjrlQEj0OqSH/fVnvp/T6O+Fx5WaaL8+OCNJF3JjX23ZVn5
UmN5n+a0801pJ09LC3WddvVO3tYDaL9eF45cMZV11BVszcYkgLM1hxVnFGRuT+le
2yxjSQksHkPO1zcRD6HCtqQM7ghJQTFlJ9AT8OusX/5mwWgYaJ/PYp59T3WQLM1y
y8w9mnDIZBwpp0P+xpV9t50k007LpkJW+rXrAEcYcNhz/RUWOdZUJDWSFS1QPexg
pLUFRUmJDKk0b9NRt772P13bKvivC9CkbvZ3gq/FZBqJP0S6spMGqIcKWxIrdT76
hzZsNgcu1TmwkHauJV9TCgZ6eC5yYf15JHIw74WDMUGpSxmBIhdzCcAZnObnxk6p
sKoAwhdetFGE1LON+vDEfmDhrxgjJD83CcsNunw5BLz7hxaA742XdC+2MapZSC4x
VsnXQ5AC8aedEMA5PUuXZy9gcLR7IHpoz4Fg7TyKYURzEcTgAq37btSpQ9wHgeS6
NaTwkST3TxZWzIvnjfGLkDbdfv+chZi0nM98AG+Kmq4gArXCL/guEdjyWc8V+lAL
n4jIY/ExszcFqhi+yaRoYrqY5P5965k9tDs4BS2G8vu42gZtdzlBONL85JLpKQtW
sYweR0LiCxXdVZnoQ0LoaCJ93FzdOqForAvcmVJkEd5bwPDSC6wA5xIHhvLDnegR
D2etNeXijHS9gwf7v6ehB2vi8PS7HAEW5WO54mRpFrlT5Q6oWEs8eRpztHOc7D3U
v+00GWH4bRco0V7PiBPUF+HOfwkteXXl2UcJyo3AjfnRmkJmumboaTu49PgB3xcV
IubZS6YxFUrtDli8z9KoFungITslOEr6cjAtQIb5i1IRdIsQ8473jI2RuzytwXTN
QSo/xv5tiJCQzouRoO473nws87zQNemsxUFUo7qMhGRA7zbPEAQ7uw+6qAlhogW+
+CaYb5i1+S1C9+eYr5CD9bKr2huR2cqbbicTDegpj9zw/1W1sPhGgwn9F9mxNkfZ
jwL4vlEHLmHDFo9wGd4JGLO35nHQ3dlZ5MIowHMGEILNB00wBUWj4QpOkmP0TAep
zlW4qsbw+e6zAamuAmjseLzKsV0nt9wwwa5veevgboS2sQeeZ2YexzqfKVKyJZsR
+gjdr985FJ9u6HYG1Ey0L77pSBheU6991RZFVZPWeINUBZBAbqPqblS1QorvG1mY
AeJzJda2S7KjqAxQGtSShk3O1bZKp0Eog7PpErHPpfBKtRFbBSsvXu4smXTZl1NK
4/b1an2gDWi5sLBxOCkj61jc2A+3f87RXzNpdPNlKSWyyo4SktR5HkXYyqVjtrgI
Vimj6fp5tGb4MYk4nnSJ/IDWzJOriqm5tE0Y954i+4hwdoNOy7zeorE0o/nhjoos
4xTeYHQpQkV5gWyoMWkYDpGI+eTBRn89q6RpgtkbINphb5iGIq5V1+6/i/Ht+nmX
a78E418aj29D47jtHf7mdzwyvK9OzGpaNUlqOZRFGmsosaPKrIjZ7iTvVsXXRAgf
AeWEmKAFFoHviSN5RE742GHQJXHWif9QpZnNFfpL8acqvBOS9TiQkw9RFVNMcyK+
CSOO1jhXEttMQsEgeLoCSR/eJ7+xmPHaK9FFSG0nbdpAC4TrQIQhNgMadr+qUoyU
/Ppfh/2i5yUXo9xKtfGEAsbv/LrfDbD4q1oFd153+SShz6aNgF1xKnImM73CuIGM
hwUtPc4f2ulByg6SamtYyCpqHmc4JRENKZSkthO/ZwtB9v5KJLz6bm15Tn4hwAjj
9aZL4sIItbJYDzSuB56lNFQ4tvtyqyB+Dty+8nhStmlSHmW1aOpHFYiFyNDqrJI0
0efAdh/BbLyWksoHATe5g1msc9LZsJ6S96sfwpOXQXB3ti6wKz2Qoruhw+B+FoUN
9y00i8Xq0TaWBFUNpi2+/tk8M6ZMWgq9cmkb27i65HcHRnVOmAOlYMnYHeA72UOT
zCf/919y/1IM3h17vNVPk23YAtmHq8XTflB+wpKeW2dE0NTBYnbPa2DxhKeY7ENw
O5TNbHEhO3de+ilGgmBPTG1lG+TIiR6XBe/8Sx9b+ORuLZB3I1rEcoV4VL0QYu3a
SiwN8JmLQejBjctNSRJOIHA7BMOzuNRxN4Tnn3oTlGib6OnPqHvWRUY/1/5b1iSp
5PaconSD1E38g6ZDmhkg7JLzCLdzBx1pwuuBjnu2MoQS2EpKBIfCzOmF6gplvbex
9ry3eTP3A43Tn0ojh3SwYVLqkAe9czPKxdKotcub2676WJ7hB1ux7hijNsyVaHXz
/VE7oMgUqzujzGzs/zIFMI4D+arrW1D5zeuK/cUtbbl6FyI8YL1oFGy+vO+MUhpO
E1mcLCtvT8r5ZOOHTKavjws16O3A53sjjb2rba1fAjSsfyqmb83dqeYY+b48PVEl
acsLgKOs8wHzAxH4SKoE3yIBAJ9sIat9q5oem4oG3lM+ahFMZMufmvKQcdkAU6lQ
Nd65VOfNWgifPXrR6t+sn3BieKYlUQs5nNpzNEhRmNps/u5g99LuwOHorCk/q89p
H3C58YjPDUZoVRSGT3jGkKMkI3SFalA1QbYwCJ/ocrrRE6aY3U2MHY2MGVOrLFWH
0R3L/dY0Fn7EmIgrUIIDhS09Jcvfxr5Udnnc0Y7+fgc02T6GjBap7zRgnCN/PqD1
wACUCTotYtVp86rrJc0XY4XDCB/M5X9hMbZI577rwQWveku3mdujnV1GFIvTJ0rr
UVtbjKEtaW0RQJxnvZH7M7U4NuxThEAEQzH3XkIAI3N2n3Vne23sW3jj4gk7qfZH
Vc0K06p9W4d3lci6vZFWrsqDVyBdazKXtOG6NPIzbag1b4NhHpQQKgGbSX86USWr
Qj4IlbYD63uHHeQMuPUE99FHemzYfstuv6xCZI7UuorCbNkqCb+FNHnI8RKISHxW
ohzs+Xlijs+dbhttGGSageI4WjLZBGtJGKSrRyNyYUjVjqfQ+NDSFTBfg04OYZLq
JUQXndIoU06lMBQCMcIFbO9UPWQR4ydwjgSeA3xTwRg+XD+Dw2Py2bf5yUHL/fjO
aorlAFTOVXHebK12f4W9rwJ/LxdUmsZJptu1nplj6j7UwRuLzt8dHN1xdLAgClqm
uktsmgR+za5RsRgDy3ODZaKFzSPp30nfBWx5tWSBtqjLMpIaAFdn5ApgVykcMTT/
08UbRWiyeCI23p5GbtMHm9w8KtVmcS7cixO6i2YiOZ6LTTwHbkXOt25D4aX8cL6y
/8K/0caTK18w0ajaqXlisfPZ255TViRxsQTbuxp3ebVPHoqbDsI5zunosSYmiN/1
xmaKZCPYM9BkpSdrnsRoYZHBWmLhc0tyYYAdCRUU/AOJ1xbScyAZthGa3rJkMy31
vew09uPUeZ+buTJx6NY1Rp+GuldeUglGQNBDLTqoXndkG1LW7U++6lsAmOz+rP53
QT1Q0rOb2Ljy66NN2UpmVPORkJv598xtPrTHl0GF/fn6zGmQkOwqKeKgWPyh9rDk
x4NDBPbymkMsHYBIhpmjpGFlVYVQtSSVY/h62lb+CWmm0vD4yWHGcF+N9taSSpy/
IUX4lftAS2zXMuDjB7r0jJzdqB26pzk8vMzUBq18k7WhBPzy/a/oGxsg3xZr+zZz
zEMi332tI85K+oDapA9mJwZzvDKvuxZGWZkr3O0ZNooe1GOfytNJsV5S0pF8ONMM
D3C1dW9BBLH0FMemYuYGK4DYQK0uy5EjZcsvZyN/QcDexXBZYO/Y5Wcdx569Rjyd
OOzFBqjTJOAa/brDmxbs0y22IJq5XHhtBJ8T9ZFr2NKD1djM+Q9OGzB86G5ZqNI6
iYnAGAyHzi2l/LUlpGULTsrgAat0TkslkEEmOcfBrFbPWRoK3hVKprivPB7B0se0
2SWEcrcfBw/jlta9UXb1NFl5oCxkOdgtCn+eGFj+pSVxFMNJbLPuE2HIk5kH1fCM
gnAlDwBb17bcG0RxMskF8aeDi5SYWvIKk7p9EEj6owMPNdAOpKLI8YPAdeWaoDLK
A1hk25cUdOuvA8ZCIKCj7dny0/Tk01hIHlYcDIrVNMiZjl1c22Hij5PiXYOuoElu
W6sRf2JmaYeLqTUaD8tkZ/7S0I/+DQEE922jmWr1/jAzLBv5rTEWcn+9g+1/t6h4
4QDk1QhFWNkhVFFvsdCm8G00mMC+I1Srt08x0o0CcOpotFlY+c3tFINr2mzye3GB
UuI3k3pE3iGv1Em69rYzUaUSpFA0UXJNodX5eYgYRYj2LS5tW30G/zGeob3lnzOE
3T42avif4gkZ5GL0/C/v+Ypd2cBwJEXViXsewlUbjNFGm6jJFP8WixtapWoTheFC
UTJwULSsid83//OjJ0/56xLjVTcymEpxYXzy7Pbu+4D1fARwnGwpOEKFbDGOoAXG
cRcf2/3bW2Hzpg+H0XOLVtcsojXKkdeNKm5Y9KELlDbaoz4+iiB0/EU2mL7RpGyT
HSsJKOJxy6yTb9IuNZXK7TAJ28M7XGGRz8OvoqWGRdfzw95wfU7JuemqkBRqRz4f
PhnsSfr9XEYx0mK/VCNF7LRY3U5nPhko+DqkcXKkafzFECzJXGrjRKIP+aKYqxLL
SC5llhnbXgGJjR0ACIrDjCGjk9tIWz2/Teu9ZBgyzKqGScBMh37wL3GJedRRCJFC
oR0gudk3m7WbY5Cj/q+I+s5IXq9nmyNXvnSHTPiV81SI3xMM1YxijAgfWCqZb2R7
I0YpEN1/zCMpFzwLz/Ez1pFhCEcX5vaM+zwi5RrYGuVYi6u4cdThHTkNJzsIp8GI
e1aVm3hD8nqrl7KWdI3gNL+cM/wyUosLzBFEKOPDbVnhh+oQGB+2OvbhtA5ZitA1
uYhj3N65hxLcm7mmjb4XjC7QDnvocDg9Xcczvg08OWH35VeTJVVv4X1x7y9Vwy8t
LJCebNJgpFsb8GUT9V40JwEFTpuhW51xgMOsOiW9EtwDY+8/eisvhO5NOtSBuNjI
eWdElSo9we1s7kNNgvS1LuPNim1bvF7ShmSJ7MBh/BqbuS+wzCj54ONIgnUZiomA
FYfpJTlx28dGDVHtOXHY5CgrabHXVYFU+Irt5mo2zdJ8ZYhWJTDPSgR9gpAmTpBu
fqopDUZdDwUQO8CKR3j8gwVfMRJIProuc9+BmoTzUj4PQQz/hlJZNtAoJxij1/B+
ZahfITQUY5cNfS6skb/yQkAyPFhduz6tIzcI8b5loLiAri+AX7ZIV5Kn7T9/t5zK
3w9mIIEJJDVKhJgH04yGVVvO3HdUpZMKMt+1tZw/bIMg+SSWXwZDkr/RiAhYoG/a
Xvy5fiWoyslTEF0LIgWPeL9lPBakOjHA3kGnJckmqYtZjgj+lU5akTAQI/D1Bp6Y
Auv2Jo8qxazip/49GFcbvkjKXJU5epgL5qCtDXw3oMepegHiF8kClGSPRwOJ6K3Z
242SkWXxPiI1e6l1UsQbhnKx/RKc79ePMaNX6BW+SrjyQ5T0bF0/Bfog7A4njMBS
W/3/Xqagk4kdz6d5GeIXRNXgr1irte+DqxcqAAZh4YDozH7w1VuAZFRAdlx55fmI
XMjufT4dAHl7bN/N7a/C7hemSyASnmBIwfG0gq9VJ9TgLYznbPGb7zhlpLxdR/It
MHc5hyydWw+aGGJqATvX4Hhm3TDYoZx7cwiRX7toC66OKOkm5gGf/sPJRbvM94JI
HiUFhvZWjrq+qEyvdPiM6JRPbJ+xG2Wd9hxIj4ooatIK7KrfzVhKEGGddDc5+niy
5FU0LLsrHPELxUdHoWA7nurHNMCvtGOA+7pMUNzoFGqElNJmPOEKYNlM8z1B5Bwx
DHcYp0pv5+AxxVF14BfYEQ+8WIkUSzNmmwBol2nh2fHSNqNJ+AalBl69+UuIWOqQ
nwjZVpuot0CTWtif0cIHRlDzlLA00ZKkFkFaw4kDg6AbsP8TWbQONj2K1MRuSBcA
e172qcNjZQfP1JzNr1eb3RuZHBN8ZEjHm1xYuPqLXJ7WrRU6Dbn9rHp1AR+BosQx
rArkxo80HFmv0hW7OAZVR8cTXqBuiDIB335PXGDExcTaEcP4LnGCRxKMHpCc/5Pj
wf0YBoCBzGy99c3Qy7zZBXABLa+I7X4fI12OOLzw8gt+/kp36OcyS34OMp1K2Vt4
8iHsU4pfuIovuTVtf4js1dVn6p8xTOjHHHSVtnZSKakLc2tKPBHIhrPGaiUkcKuV
2BL3yfBBv+BuSNDAuOx07S8AbhwCWNcWZ0ugNWAOlShGO41HU471h6F01VhSwgBG
FmtjulSg40uoItnvfn6HfabRBeJ+hWYMo5zJwhQVLu3qtWQS6rkgW5fwJNm5vmp6
quLeR+vP4BRvbJkJsJMBu4sy3MZAsLHmhuJ/SWyTduqboR3z/DR9lCCNFvUfNe9W
Kv8TfCr6XJo/DSMkndXx6Gd/HHEMdWFVf43jjQtAq8ySj9Phh/ya4MRI+Chq0VZw
yJSGYWgOdeUXiklEfqrc3NV15uYcxFEeuOhIYlaQKgRarpRT+sWPk345yUhtB7An
V+7xjS1GGXwXeSAX60mw2dsUBLslp/TLHIlnE06VU2bjXM6wylUJTTlSgumF5G0q
1wFId4FVDgcUAMKWmxlMjeO5Qhl6uQpsPCIW4Rnotkggka4F0frtdSDXuit3u6kC
mHcsAj5OFGDdoXxwb/sIuKHxe1JfwiH1jEP1dr6ows+gAhCVQiXuSYPor9BzaoDl
CawqpMBbD76F/VMpWbX1vGd+8aWW64T7el2vULv1r5iny53vzJOc9f4NFWOdM3rS
I3ukrWa0EyIuQAY7CWm4Rik65zs4UIeet1kVHt0kMcI4DHit8u+8aTIHQ9OBq66y
UjwRc4hRPnju9PD2LTfBf/qmvhaMdaJafcZw3hu0ibSM6XTf5/h5D1D9YsySCyHM
E0BxiKADZv79clNkwTY8TBLBO6DQGYlNcoavN2gA2izx8whKDQKfLOX2UgYLuiry
nhEI7jBct5aCyQpf10R64Zoc+wvBijuALsc+fnyTVy0j6wVcDHgylrbHHwAVqjPE
/+w2j62LRFWXaUynW4GClisp+piccnpt1MIs7mNhxUg+Fk1ynJ5PtsPG9AJEbfje
zKW8E/dSdW3sgQrZXMxtnvBbDkNASEVbrT4tDpPz11f8TBbtQCa/nvwNrDx0mQGn
unxb5z/y864qfiDz+ababmqq1wWI460fO6aH7WgB2ZB9s+ECMPjnr11EP67SeZHw
87UefGEGDpHnqdRRRQi+tWBVAaTsC2Nexlw5/eJHIaQMU7H6skfottmfEbbnb9Mz
hQMf7U/mVq0bhZegVE4kkgwQVBKliWUMhmkd7URJ6Y+2j7JVKgu+DDIRZAmP295j
/IJKDWosME1RVbstS+LO3QsL7k5jm9Qmi+enn9w+Xs/vKc853ihS+RFcRLa7g/rl
vsS5EXS9O8GoCk0aOPNIkXTaDyf8BibBx0Zj+MhlolIGkhce+tJqlVwvLkBoflUK
vwZFzmkT+8aDwZ9SCDRxWSdsg+rdDeRD2yHxVgxdWR3XkchrQJNNkwbjwq4pdDTs
4PxprnMWnlMb4DIj6taZJkhAvcomQ2jdH4e8iqbN+XRvGS07kaVGeyzHaTfC5CKd
CGCEyrTIsAAjVogOVqKBTrMvNmVf2zMFK1QLKTjoBhU/rmUrFHAAODWYcTkAuaCj
qrvNVQvTdwC5Enf5Qho8y0C20rmnhUc9E5lvDZ/iYbl2X3il602cDbhuyedI4PPJ
3CrkSlwfStjRQaW1hYo1SLQz+jntgc6J6cQpTPAEFg05xyXcU2tQtoMoO9wcZ62W
onA8pVH7APaN4RmfvxP4lWxkq2BjtwCRe3Pm44xu2vnzOfblGeNTPw66mnA5++f1
c12zvGW1qbMhu03FGwiajn3yYwS74Lwgpcka0OfX8UboCyObh/BW4WQ8N343XbVd
KLpo0+viEeVUHmTO6fQNPO2iijUAaMbccmjt4VBtobk+o0g9vB0/8lihWVoLBsD7
dtHTtbF4BCwHnnIr7wJbetslolhezFlLJ0BHkLMYqbin0YCq9gEsEfq2yz+RfkhD
qLKaanQAvpruiO49FVWIjWkXrVT226tUP9VwOvBf/8edeWCnY7IvqtnXRlOMydbf
M1pLEjJHnfHvOgH1m8p7KEQw7sLaNSbeprpTd0VnKxn1SJEXnfLXzLJziG1jpBr3
NojtrvHyN49Y4TN5tSy+cyd69sDQouTgwEHvJRuK/3Xqrm7pbbkRyca0e/tQaaI1
dPwYrSWjvOzxODb2QzOO7ZJbowgdmGVLH17cccPZ4VyDuX8tkqc/+2srxFPE/CzG
nCeL5U6qjTfQOlQEVkHTLjQXwZ0guUFtUhauWwBPEYHyYCo8FJyQSVYTMJOSxrl5
5/6rPxUvYzmW67Mxn+ZipvPBN3yXeyEyC8sllkUmP5yU8U3ehD1ggQUf56aA8g4q
lp5DberVRl1KVj0cntchZos0Q/EhgYWf3wI/9arZTNMKpt+z4uT3RQuaEPnMTox+
9kqJPYhh4D0LFplPjZ5n9ucYMW1Pv3iP9JSgRAWihXH23GEQNQNDJCtuN1UMNfWT
Je7WllXVHwHJcfokkSBTKR+kI1C6+FYqTU9luFRAai5f+Rbf7GKb/Z8m4iFiN3L0
UACO4Qmvn6TOP8r6OmuhtHQXq11eYZPrgoqrxU970hnEmMlCQRoOIvyz0SkQnts0
CCf1Yl20GxeAYz7cPwyGIMBp70p9O2zLySTpEyx+VgSI+eC9GKJS59vf9v+h8mA4
fjVO2/BGi1kiTbCba/8V1l16BYqmD6vG+4umP2qVqb6El3HiZfn9FJcA+NSNOwq+
X7oOOTY4XKW7IA96euVCrl60T4/5JZ93cSUYt6Ljs2y7Dd5YTFn/NydgVPMI4/AY
cZtwkFb/mrJLwmaFz+f4jJwIJPNWYKCsBqTNJCUEK91PIqB8Q9WBH+nPV+Eauw1n
W5I2UOBBVvpfk9Q2rMzI/i2grVorLVA+bOKTU1OmrogbxEP4XEiUmpI6KDl8qHJz
eXd7RyMCBgx15w8XzJ76B6ydcD/fM6qJvcBcyjtduDOQKumk/tnGjIvaPMvTFESc
mZsS/AVahuDfN9o9QSc6HPn0KAVFMhQpW5TsLhYMLbNmDmSVvvrc9u8K8LV3cy5l
B/GhaUCnfjdfBKrn27oINYHrQhAoJaQ2d+MeQ+MtdizCA0GWd8jObUPqGGU0qhxu
440fxZVdP1a1+RzjdODWI3PH04kkRy58WDrt2obG+iATXsS5+ZKBju3LQ+q7TZ35
hEJGJzldT2XhngfHsAceF29n+XA56rkzjd86QziwzX2sad0Vzjh1Wc4NAYa9jjvU
ZYEQYHgZMIG4sUWfSwFfDVol0mPQn0yJ9CkCsDaLzB6RF3ia4lfssep2CVyuHQ9v
PYWVmsdZ5/D6Zix79PNqbIyhID1DcoejFADpHgTbrMM47ZoTEgQJAptSq75+A+MW
DQCZVx682Xct2NXkqgRYJvKAivB5z6h2VgJwkPloY8Lg/leXRwwV9ADDIYxr1b2H
F2Mtmd8p8egB6ij44Ae4bRO4xPI3mi7KJJbd7Jmarwjae4f9cEms8XSd8Nc9pxAu
fWS/U7Oyo1kL4YM1eSAk1VxM3xmNDOl6gHvHSFrf0VB/558u+SZqTDQge0ejlaqh
Ozpyiy90aZdEDuR/s9MQ4I+o6TQxdb6Js+8BmcuTdirKYpcAUPEP0b5U0fROKhnS
njZYdjUw0v/MOl5ThnEqnA38s+cMjJeUuf2S9FVNvZ05TAWYX6UdPS2RNVR6Pz3D
8fU0dalbvE8QOOg/uN8XN2ZSA6/VezO75oTGO7+4vF40ekR85dLzXv8Qkij7HO5M
jgIAIPU9hs+e8YrpQlWTc4NN1JymHFEX1Qyj1hEHKz6LZyS1rjDtBOnQlqXUq9vX
VSGZ1tavoalpmaW6Pzf6L7hKJhaKyge+rifzyk/9PXSjz73XbrIo69ZYNxHmwJyZ
RI2CAWDuaa4WXf4C6VC7H7NFysPuN/pMbtasKd08BXRGb92EbUC5SUyAjZHP3X2y
EZAIVBfRNbPVRY2+oQSfmOMXRJGMZgWo3ASkffq2orCwiHKyx4T6wg553jAc2wP2
5zGa7+FdAbju+YeqOu+p2p8tkC/TU7dyUKClhdCfeeVTbdWbCCVVYVV+l71sGHIW
ahJbPni6HqW6PN2ClZUTq66KaVWLOf/vgR/wICHLdmh4zpcoq7WE38joQnW15KQ7
fZjchGSFo6MFvDx0MsaEWiIzWGD7S0U31BCuxu5rn/bwDSe5IYuGSTtAwZVdepFO
a92b8enS2s0YjyiuPKVpvcZ0dJQ+X6FW2XMwzyWVSnjjoZz6Y4POVFeLF7WaG3fE
daKlpGFLWEHwa7mUQq73kK4kk81f0XSWBQNrFIb8B5oOybf0dZI50VoiTBw1D7LC
+jpjoruwbhTwnFWF466rd4Fh8kuxP6B6pA2Hp5rXerSCFp2iyrxQ0pe5O6rMYKKZ
e4N7mi0kRt10CguVaKlmzqQVh9uLp6gj4H/eUX8Y86MLYHrn8geFg9V4RzKd/CFm
QCrMSv4euE4wuvhCG8+nxSQVSz2s6EiuKuTOq5IFJ+8lH/7trjOJXCVBPUYkWmz6
Efv/noKSjJ00+zp1PCWbgHtohJ7JBHi7SagckFZo+sV8bsP/00VytRo91Aru9BGM
fo3xCSciM4MeTDibHeAhbqef6foPh65MS2r/iqRiWPynZoPqdQxZ1BWlPeyAsgfm
V8UJm6kreLDmCChSXaThn/MzA9qyg0EAEPMxCPIIDzd8vriwp23JzLNVcJpJTncG
OQkn3I5CWAv/uBHsh5hecmtpNIpA7uuGZlfcKcPVxmBd+Qgd2H1/QHruiK7KtCQd
Kt0coDqHf8slsfqmcT2BYTWjIYuUMFqf0bYPuihDorvuiFyvAzVwanpA3zqwg6nh
v2zuHGRx4cSRYNBkYq+jh5du8eiaP5fq7FgbQrf5epI98v4c37/6L34LTRZ523at
kk4AISF1JZnX+b/1dKYy4Lt86tDKCJyg5wMENf1DIsiPJNReyx19YFAnt7lMP2Q/
qgLWlZ40DMQ9lQgYIru1mxGXNB35X/kKqVuMfTEC+WtxvSl5+y3j8VQk1XMdhj3Q
TjOygSBdGyxMyYbHbJmgqRmMhaY/9B3+7Rs8BAToI4fO0XgZqIWaH1ykdixvGtUX
rusp05K35WsHpfp+OwRKze6zEap0XHPcSXxycc2CU8cS5wJ5Ll6feH9YYl53myJg
oUtrijOPxmBAE1kaWOfmT8T+WFVq7qQ1sWtwf5pyanOiMVw0GEVpW+31StP0HB2M
MbnSKhWL0G0blq++yZB3ImTKHRvXXscvrijA7ZQXXA68JU487tr3c+Z3e6wGnJ6h
Dc1YR2HvZZgAiKpRm5H+98Qp0Yj0l8WKiIu92Y8f1joyGVyathNY6pPcw8FM26b4
CIXK31qNQMpopveS4nwXU16B7fbi8HYuIjFkQ/B8g590dd8LrxxSpYU0IG0EDEO/
WklZg42gz+Q9n/rwg3PPZtDJyPjdO+8nzVtE05E+D4IUH+Ylq8HMi2YU7m/U+kuO
LkRBbQHZNe37CY43xUtGajW96LHjLFBsrNEiOj1XaCSM1FDr7T1Kz3KErmeYwIFq
balgBMfrNpWvyNvd6rdXWpTMUdpZEfwWR6EB4fmY9qCMzBK+whDyJDzNdTUzi19L
7ty1KfjHotiOiT2H2EdSvryFs7I6/0Gz7j475JsTwJKuNbFS95Gd9+ihtphQReL6
pnVpjtzQtYLgXaaoL77jZF9F+q470Sp9235233g11SRMwBtkFHFQwsSJzrbdt8iq
3ObhW+o8h0tNRMMxDKX4keoFkTzRwqsr1P6y20Y+AmT7nmRBOaaBnOQoP9xcKWU0
ArG8EKI4N3E4p469GjZZj8cc42QXf3hBqYxIIwfxRH2uufkGsSa1Nl1d1vuzhnQr
GZT6xCfA9mRIgiq8nrWBh6yLJ5sLr8mtradB6lYLGWaL6I4I+Lq48Q5Ozn3goBCa
WWXL45M1E0RHp9bufSwlONADeB29RjSZKbGhJ0fgQvz5HMycrDtIrRWqXFl5KV2m
L7BVPwHCuoeNbsawvcQ9OJqUvFq67DsEslHUYuERyBMKcN/pU9JY9yvSCZNrMfdz
DAr2eTMfC4a3hYI0V1E31SgUvJbTYAfH2813MNO5NY4yh3XjwKqjrC/LEVHekUWP
7GMPpol6Wvu5bBmwfgaej6ZaGYqxbYfUBi44ZlReNCwznQA/QghiPSIVmJSLiAwJ
KbdvJh/elnpqdT1DfhfwcIP4G+eQOHwYdSsVpuzN2f1MEya8rG2j65lz+jn5C5VU
d0zx0/WH9VGorjGHasPYKZh2CDd/XbsAyX+5pEQzszgxuV2BD+Vua58YvpwfP79D
E02AFMDL6nm1AzGvDWSvu2x/8zNvIadUuuei+Z6q7STNh7f3cUz9c+ChdIRZomgt
dDoVz4W51/ig1sg7Edi73Ieu6qzwCIaS7rRsDHdzmkXuEpwqQqe53tfs1m+VlB0P
HxC1GLmeFFjSpi+7H8JV1qrWQ/r+bdL05ecgzhCktdBPKDvzRXSYiL5awohrPqK0
ONnrcjP45H46GVzTm/ZmnlioGISKv00tkpDWxy/1a8gK6oRFBZdZMg7vfUaSG78W
ZyxrhyCmIuq1shzhwNboShwmXcZuXCG0vE/9yC17760Lj1JxoYZB2nP6aizIN1JM
Cx8UsAY5GIkMbC+lalJrcMXePqR2x4UI6ZPba4DQPWhpiJeAVigWa1WoKSHERU5p
eXAk56dn79CDrkiuiOm//M0G7nF6Z7/AGmqZlbnK9Ya5+ovvV9eJPPtEOrxMetY3
kAhQ+oO+zE3ngJGj0d/VCaBDAxvHabnGksVFjZ7x8nIhSBQDf+AzGk8BlHtrllie
MDHLykINk1+OoyPnHewFse2tDJ1kSq6eRfOGDZg62ADFhGuBwmDjz90dldPk4Hr/
1KvEDl2tZCvBe5XMf76e0aOsN/2GusXfI7S56BD8rEFJFov0ops16g3FuawKS6aT
NWU3zvkgPbR9euBflTfyIc+JeTtidEEzSRGlmVnkgBPeaynRhnHxCP6B6IHsVNIJ
/Sk3tDQtKV0lnNJqDFXuTJhyvd9Iw+8mqxbBRNTVKSm5wiy2FfTOBgoJhQfmaXYA
sgThhxzuk0cdFpGz0X25OdV9Yo9/9++daPmz+bBtDUmFBdxl/GeEuZ/BUr1zVUXq
cNWxc6t8tW4HYi1bxQQ+Z0g9NYQUUQcVPZkbTRX2EKXRe0ODwmVZHznrq3Zj58U8
LLXytGw7B4to5KdGmW7LvYr/KCvlopKH3fqhmScpZYeDuPbRPZmYwtLaHCr+XLUu
R9uyPPUmKlJwVFzvjAnti4G1Gt0ri2GBHn2E3mjLs2EIIXWcsA/YQ/a+hNLcrCKZ
0PZ0mlxarwv0GuWRHZBMbXKNHmwNf4LmYUB35/+T88AYgJLX2ewUxvbBbbH5p5dS
NT5lFiveHTkEOqjqnyq2WPdjgpb7s4tgzDxJ+z1CA6R850XzwFbewjqDFXkqj0tO
ZkFj8nW5TMvFZE5t4hqHX0mFRD8KYt9ECrKMq26voVPSXEU7X0LqQn52FL0UiX50
P6hSP8b1lTGCj4fbybGrORmG0Y6H91rJLROVToTYBRMKrk9CrTQIjn1rESXKUhFS
iziQNbsrOI8D16qOXyJk5582hAX/kuRJRxXaD/+uCRpZ36BURPVWjZ5Ymz869U0I
A2QB+/605yynEmSHnof7R42RRMZQkFcBzkM3iNbhXNlYWxPL3+njcJ+YPIzmdLtv
7AR5O3yqkIj0+Kc9OnYC2ohGWGcBh4ZUDbrRcqVRf8etYAKneDqkIa6A7lN0FeD0
kkiB97rEDv8fxUxmTDt6enBGMWwj2qWIxlmaDX1oMBirI8nZaWcvwvXOpbYdi/R2
B4sbFx6nyekIpF7cxq+VcOPC0qcpbdbxS3cgxUoCB3LahkOho6VK9QIYLer9M0MB
B2xML7TazwTRcIBIwOpsccEjkMHeXciD3eVobCR3iVpXIpMpTD9zLfXYWntnksJ+
EIG//YRZSG0TkNl9uBj9x4SmHDH0QQ+ACOet2h3VgxlGpmPdOOfOEMPkMgiK3cOX
AMxxhBcVGvbUsjaergK8sqvh9XHbSQg27TftgsFdiRs93pK8z9Legeuiuaysug/T
UJHJ9g1uVWxu1hsc7fNOTDivAIk2SZgfKPvM3I4ybCO2eTTBn+1IaJsOxrIkUteA
jxuIAV4GhoxHkEgm0sHmMAW0fQnt+BDcRINSBo8rS28vE/aSOdItqHa7hCSa1341
nzyGozGCN98ekjxZzPLEIguiDP9YDpkBElOx39ED+b0bjQzFJmCMxgvJGLUkWkv/
9OepI5EjaVxxs4O1QwNHYd0wDqg4iEs/n4/1LBSkLWjEyXh1MwLqCIkE6/5W/V+W
WNdlml34NYs+98ORgNHh4fytv3qBXaxYmfR42XBFDiVR1ylUG5T7JqBs2+7UB2/0
/ZALDFdbnMZrPJFxX+6MvpMtevaLcxotPkuqXolfswquoa4u5rj6UIm2kJw7tWBu
yqow5b9VRj5qk6e4GdRJj/ylokj1KwfglIDzPFILxG7cmUSxRnVS+QP+NwV6pjc+
ob1HfCzz7A9qfTej+4p8in47+acImlMgkpoJUwgCNE1hnwbIxziKyE0NJDU29t5H
50OvBK5KWrecvqwQwxhAbYE+gyuXExwRh0A04PjA/e0V00oId+DdhAtT5EtH5HEG
1y11wfdOtZ8gy83ypfGNHRAybMfTdbxkmLlSdtPkklGrhP4JU9Xz0K+TenOzhrUF
sRpYdSIeVs8+V+Y4x+28coTJRBJLJlIdhHX6eHmposQ1rtyIPgOyI4EDcgAFgqs3
O6UO4tK4eGSVaJ2iv3RafY415Yyzrjov4scdgMok2Tv6lcrTDP48FjUEDifTOvsh
zTYdGvqHHiZsQ0T0+qFNNa1JcM0wdmKdjn0w672QHs7DRTWl5zgmvwd5SIzXhfqs
pC76VWzShX83X7kFQ6RsgK+AOW76ft6gIf88DJGqm3DMM1d55jS8iinzhTm4ywGT
uwEdsw5XhL38a8o4NxxB24nhMA9to7p/9BcO3EG38jsEIuFtiShHnCbo2OmTYLOr
e6rp7ZSi9Ysx/vugxmvV/aUDJgBFYn98403ANYTVC6+zJ3SrhyW0vqAPtcxItRCU
ABedYIkbKppDUldfsKcaFo7aaSg7JUZTYtFhq8kgsCP1SAPzxvE1pR1fGcsh0tTF
t/Nca5LxxP+6gHXytI2sDHU1vqsjH/nC2jfFd04ty4XOGSfzF9DzGYr1fEYFEvTB
NMWbuTFzHq3Y4+LrLuPLTa7KvpN+vpkfMf19KC7FiPipHIG7fUidCzNqbxwILQn4
8GylzL/684FBBmQkDUlDMkNOpGqVigSPQLQ7biqDyl5c8Z+bYzM2bRTDFy/jLQPV
v+L1Tx3psO9/+LRjDzRYLyF7XRK2sMC6ZiBVSjBh2w68e3StvGNnBg7RdHeElZld
7KtzBfrQS2vgchT8mXNo88FuzVPbJc8o14rZ8BtMHTkivz9aH0miAXM7f1hMacjd
EhOTdILcuvx22jseyMzemIruLcFXF/q5yRK5O3ll+4LRFMC0lHP1JfX7YikpbLwj
rtCeE04FBiq3CY65mt2+PWXaJi6YlRavujg6BxAPID03PrYR4HPe5xp91YB6hayx
TztN8jgU19QVI1EW5wrnsON0tQwT/vExslRP/IBDpnDpTr+L019lslYTXGM0YrkR
7vhMWeyH4i/zJJ8daci2iEvMkWZNceo63ZHDFP0Bra8+MByjweZdzxMirxeUDkEv
mmLBESTE1QaGC+miHEPvUFwKGuTxQMVNLQOV7wodMXqzBHdpxn6uARDr+Z+AxOnc
0oEC9mesvxagayRElTK0yJ8l216hZsg+m6vd83gTGR6Hsy+8jUIfQCJNLXiVNvwq
maOa6XA2eMxp+Ne3whO4yEt41GlxiBE4lMPUYGiVb7nQmSY7xCD/+tUzaE694hnp
UTKODbb5pHRK6g3au8kov0KdvZBbl/psObnjovx/tVAvyl/ZqV6Z5mWnFgvlmo8S
5LPtw74ljK02Xkv5E76ENUFioi3C+l60D+059/68q5p1V5z1EOPU9agW3MwbCYe7
33pNN/aRI0LkzKe174GCdJ3hbPmnYTYcuyIXXOcrWRvDcioZsSVlT0k76xDxbaQO
L7MGAAMNJpatnuEQcnRfaWcoueWuWT1qgFZ7J2L2nLU+JLg80FC8VpAxuNnSf3Yx
e8+M3cVid3VXtlYI7Mq86VLo5+YV416eHtHAlAt2pVJ1GNBllie9nSNDwNmPKJ75
rxKbzta/A+CfHv6e7tQbtmk0HZ0+RTypnNHph/zUrsOqCztTPVWWleIPtEYmaIAK
BreHh8NgSOCvW+EXGIMlrMsb9oi7pL8oebYh6peigEsrw/R3SX4EDJMUKvzf3wEu
8uNp5O4FzgegzhsMVxTVUjg2EoSkXORyMd03hM/8Eg7RDLKmKkQkZbeuqMLU5lWM
ZC5VWrrFNOQC2HFKyfBXLsOsajSl+RCKiPmKeVHnbx0prIzeDqJQ+VqpXJv7jWxG
hy3fj775J3Z+NqL8DEdPZSjZC+dkigwRGJ/qcXOzjRvJHjW0cyoODK4ENnpddM1l
1P1+LxUuM7VwmUNBewobVhbQp8VgyRiqfP+GEEFUJRWEFjRbbQI7BrD7f0Qgugeb
gzwqbzk++dM0u2bmtNWM/Qn5l1Yh53IUQHSaBdPzXipM+hkYNEaJv61os9TH0cCV
U5hVzQJgXJ6CmHTdSOFTW9CvOmrNv7ERDKu6Uxwfi6mMTqsCabboxhkn/R4AXxFZ
M0uO4caepLGyzA5UXOnK95dCsmhrM25EWhiDNvXQl/m/L1SIaFPrqUB25zXyKGGk
dJsDVBNtp1fKqlLV5upV/OlwN+gyUteWAv4++L05LTQIkG0exxaW4T0S07GUCxO2
hntA1F+g8O/cNIImkAFX305SL+jHA4mHJ1MOWDgAaXy42qFjyD7087jTUoStKMng
bbeAebCIqMrN3PBefKLhTHFNkHp9b1a70MwmIdliCdoEfjT/+E1sIVys9ntmhRfL
4C/qaRdw+qISjUTBP63Gqp3Yo8DpUc5FIUWRQU6TQgG558aJpLsDew2GFFCrNk+9
EccWPByjW3RRY3n0bzuuaj2eFGqe2l0Ebqcgtfap2GAZdXVvXEnBxaKZJxxtjX65
SKJzzwHC17CZYlPoCMtfnIAP5Umq612pjQv87H4qz+USrvL+c7t9bU+TJo17q1Kj
gnprf+mMb4vOI2WW86ouuXdEOSPvCW6yDa/JaAzl/K0qBuFxPLIaeCOBmXtrf1JU
siqSsQXuI4d9vhDGtoyGY1S4NnlBqXntCCcZbX0ojUF1J72ZUw5vWldSlwKeh7wR
euQHhoFdU0cJXaNnszVhROuZH5oFvmMmRiSoMJ8lklyHBoEZ9uqoFIl0NmXNIaKW
3EcHrkqGAP/hcmzdnPTz1emcj6xwORSihnj/xV24cNjiCrl75R9L0CTsC2KG6HHs
UAdheLCblyR+AZXCRnLYq3rxY3OETV7p+jFIS9Si38QJLnQ+qTVCLXILlEmHvpVR
Bqh2tzXJvvthslOW1fqnYnuyvM9e4dlqqINawv2p3GDGyzYk8ZtytnQtUiyPL9QZ
xaEDsFfTgCEAuvy9McfHyJYWzeFmoPI1aRhwu6IPIytFTZoOpqYiCVYy6q/fSxAV
OThR2tELLvRfTuNhI8q3pxxLbB4CH5nxsPyCW2Q85FspbizP1A8HeA9tzAwmJeGf
91e4wwTZ9aOXtofy31ZqwJ7wRJjE0Ubmoo4WJqB0QKEXRgQdB3OblFT9ftwHJGUx
MNkhEoN0ik7ofB5ryY/6KvbU8XkIX505xkRtQoGBLLAsB3h1quiv5VwyK2u2YN3q
zYMW+z4LnAOsmO6CpGHEGwdMCEDiXj9kGxBzOSxRZbzOpejorFbABY1QXSnUboht
xHQR8BEByedrvLJZFOD/vgV5FIxt9aZ+pxTf9pGfp9uT/bFuJUns8Q2cS/CWLR0P
sCBAyDhhKwRwy4a751WSTNiZFRfp6tTP2oGX5Pio0pQekJITCzNaiLmyu40Enhrb
nYUne3pS2CjlVDnMfDvrBeXpd2cIESgO/5AmVv2qZaUoJ7LzR12ahi34yxZXruXb
+l7vo+JBqKDmfeK3DFxUAjAZOF7fjYFhHMnIC8yloDrB4uP27j4IMd5nQ96l7KL9
CH8TGazPwIt34Njcsr9rJ84uvwo5NwhzEHFFlOT0GWEIMR9Bv3MBGNzB5kFx1m26
ITxsQr0vBqHgMUQ41z62dfxKnk0ncBecN6034Jkkes7XZCcXxBlZ+boThXJ3GWE7
thfu142DtTG2srZHdE3LSCNCtvsUkRHKXqXoryx6ab6NCjX+heFsaTurQnLZCA8x
HigfIEAQci/n7kYYgZGNs5y7wheLAXF+2/G3H8Ez7Ray66dlR4tilgMl/FkHGvsH
BsJjeO24M9f7jGEhBEZXYseCTjhLNd5EaX+kglbnLUpB51Wu21/yBO8v0OuxzvCx
dnRjB0MK3G9D7olIyZUgDuelk4lqrw7k3TX8dbx0ps0L0fbIp+B2J77K17tonOEj
Vat258hXb9krvTenKMy7mf/1YqEZYoLdUVMVGynnHfBtSGPPpZwsRux2ClSUX6QZ
BimkO+r6KoyuioXf0SWY+88BLhDh2I0OO7vw8DBtZue7qDQMNouVXEOnWIahGw3f
0pD8Wtr6oiW/H/yV5ZazWCzW76W9kc8enuywJGUat0kLk53RVoYG9NJOB79qR9C/
yR8WuQ83QFEGwyPR759pa2y3MAEwG/tQFa7prr2ZGlbH0e2PUMpTC68aEPqV2a3O
BT7S91emmj3VKup4vUDVJlrmgzYQi7Kr0et5A41oFS4pIcweGIirn1tIuZrnoyde
Zcv1fh7hNJnRGhqdVjjw4tAvmnktuAcLkfV6kIb4bxvHvn4W9qt7QbhXhPjPr8LM
5BLH0qnfdaUg/1VFPYC+UVIxu5RTC3svHyR1p4jbnJ3lFbcha4OnDNk+hPfXBC6O
7RAEn5lUKP+guAOJFyIl51Skexg20mrLdHyKeJgf7McUWQKZQTt8DqGD8W/qVjI5
CoF/yv8Rp52fbcAB/FD44yjLIDXEBSfotY2qMpn0qU+CU7vC91WKMirrSEw7VVSt
ieQr7kmWZ6trGQt+bGq9qAF7RNafpUa4lfVcN+ZPm0/nxvpgYdR04BPEoIEqSvuJ
kze8FaBv61ozCp7LkRu+YAf5tIqYE7RgGLGAHy8fPdzMqF/xWzu686Ve07YsxxSF
a1wzUwqyHOUwjR6+kmOPtfs/gZ+8fYOBkkgn9zRac4ejpMsfscKfmlkrPM7+C3yt
roqZD23h9K1VvO4o0XqFNgrkv7vYJoSQLxTLqBlehUmjaidMfLa2y1UTXF2YDmeM
raTmqgYEz/gi49twodI3ULoJkEN5fXVUPbACzeTmtTjMr75c8n76CdTtcbaZQKAc
nni4v/4se9zvGDIcWiKTktj6WZbmKQkt7OIoH9tHFUrnbAzjcLA9XEpR18LTKGAk
8CkAwFCf3g+S7FPg7QnjmMhKVT5vCV85T70BfQxPCGvqr5NTHH0iFVSJ8+dDGe4H
pWI26MSOBjN4nsZiN7exQMHT8cdAD26CbqTyIxzkgaWbDIPfiFBaE7VuV4hvOL+1
aI7ikgyvloI8U9qBPjpvdtjGCqImJjAUx0rKR3Obe1IJmkE2fylDwOI4VXR9MmoZ
bMGovjhU4nxYXeoBDzk1Oid5+gltW6NOuirXywBWdOYN66yyPKwRIfDgqttPQzG+
POgMeVUogcSnMu2z3aQTxTQvznH1asX1jXnayTZT97+b23RDIOFTlv9Ar9W8UHY+
wzfK8TKvk9zuVksoisJB/QGEkkH8KI+Zo3PS3V9kWLwhcJohGuTu1n3IoXZczhFx
x/HPN+wJ8bm76cZqAzJEKdeAM7bA6hLYmyJMQbNOkx+YVNsvEYSz62shAs3fLrEC
XE5x7RDFH6KRvp8J0x9QUlD5zf6kbAY6uFM8CK8+kJxpec9NixU0aICX7iRqXipI
PkOiDqCNxvpa6MTuDsiOZhmDNP4UCO7OSYZj/jcKtNVhv0WP5cbmF1afo2z/Ae2G
GlVHibIUaQTXx6IT71/+I2Ceup0dudut4oZF/SsnrE43sLZtxp6VSaNFIG1ifCcB
E0OI/DrngwJ1X2pxYd4kv4a2C2DhCjLNYHsCPPvNZ817de2iSS2s5NKdkIewX66u
t6jVJgeqtB4FPY3/6b0UbR6BumB2cX9aY0VBH1+XOgZ1nXe9ISRja65n8ZXWWUpV
F/FpnbPmcLZKDaOvAmJidGsFWDYShz0XV8ieAsiY+RZPwUhsfHvvALyubXn/lwFi
p5/cSerg2A400n6bdj1xMqaJlb7cJWx6nSYru1p1I8t9ssFPcLjzAmWZOl1SPSZm
x5g1zYDuZyIAIV0c68N2hXlrpf9FIOYKYhrIq4JzNPaLMD61s6gROrFj77xBoCTx
4pUa9Lc/bgGrOjMMVubtRKUs00V+qgfHbZUW+qQSK67BxMIxjnfFIu4eLonki6oR
RJBN3dlXx2GbmIaQMFXz6FnlJjvAOO4II98YO7KvOH0GGUCVySa/aRpFm/YdjkIb
sncy6Xiy89b7A8h5ZEXOREclk3LA9lymlf/lWFxvZU+NEok2kyJMcOsAdhRaWsgR
2Oxz8kk+P3M9Yl1xhMN6urBdOQ3YkBHCtti/uqoFMe2Q6hiuDNTrG2Y9XHXA13kq
vZCYCt4HG0R/6PDZns+WUDxhezWqiiXTmNCXX6PDj53RHN6wzzFWA6sXdRkr2Mfw
ZXuW+7PjLOqlyBSqfZt8ZWuOVNiGClB3mHlryYXjs+R3Y3PJD6Y+ZpqlYd429Fx4
esAKltKqzjC1PsHSFG+zgMpU547bHbWuTOP/ENDbtQqA9MYEf2ERnBU540JjAfdh
YtS+dt0lN/aNtrz+rtSU7/N0Vn7cMH0L3QhDOToof3t2ZLt97piSS95quvanAEJV
UVL/OPJ/Vn7c2MmzzNObHVAKOysDklutttfvrdp/sF9nICaXvy/BW7GVgyVc2yYk
uLS/l2B450PQbAzeCbk54sDsZ1xwcutIwnc2dX++Z/zhJ3ZljC6ANU0OgysNzV7v
HPhrWQUysw/PlCwRLYqn1/xuQLOLJ1wvVSNxoqT0gXdhTPuxwtC59Oa14sbT94zz
yM1n2DTy3Cw6n5iWfVm6vtBpoQO57wJn42cBG13iHZPSvqHym2cJ8l0GoN4WoiKn
rLzUJatOvFNtvHmrvCRb/KMrdHYHE0TWMMX5x8D5cyqcsm1PGSK/Kesl/1x7lm/F
DzOrhDwTL6ehsLuUA+vVR27dJBgOf/iIWFM8VDY535vDX9Kd8kONgt0+iZ8SYLv2
Rf0Dj9BTS6NC8mOcNXdeZRz7pgM0hs0JnKDytpUp+rlEVvKujrt3+GybzXlZz+Cq
x8bqommGuMZ37bHxQcpcU4axwIXZ6IsG2F1pefW3JXa0iIZ4GUplcNKuOGYC+UVv
AksM1m3IasGkSwgGt5Fc7iISjqRzhGrCDNsHdSKwXsGQ0UfCpOHz9DOKcrD2dVRe
DX2CM40xNFPIdjjdU6eyk6FFccdXM0Y/JIRctOWkK8Ke9YWXuanr/M8ZPQZr/1qW
hsECyg9/QWLe6y8Zcynws2uunQ25KsD0cgEx89ZA3/hkpmyLkuH0xSLdjI7zenr9
wMNfiO0fADzJVeZN0k66iUKF2zKiI/KRL1/Gr0aM2XzHSaQ7QDvkHEkQpg3oaGSN
dxRh+tEPbAHWaPs+LWJMwKxGq+tF6QWFn0skjTSN1MKYcX6QLVJemudF5Cdh7A4k
iREwxGBl9pEXiWZGKG6vPkinWuNo6jCiivlJC3sq+UKerfzO12o3sLTQcf+W/zTv
Ir4aJ7c3lBmiXexk7IfOP+qEk+OaOc9xwl4eKKNrCzzBqJQ4Hhv/tNx90IB6tFP0
agOPkDoycE4DWkdNrXOX36wEivCF2+VRYN3LBYu1GwUWF+pTII1ixdvpI4TCapyI
0k7DfcDzRMVE8geQ920TICEkFAd/B6dNxg3CYP4AxKPV7l+WIGCbUdvI1iHBZa09
ld93PUz6ZPp03E6fIrcfaDi1Q/5b6USfWjALOca7Fil7gzNOCewwscFMzbbs+Ilo
gASZjg2Yqzo1FPgIyHkX/Z3hiIH1Zf+fuWEYgpLBCfjnPnJdLHa3byejfUrp6D3C
T2pb5EABywUqGXlMkvnMwMRQyYXAZ20vXgKLiaxnBrLsQ93G3Gz1zGr48IWjOT4A
ujv4HhVZnpYOM8t+9eTQCPJeVdgNhkaIsTwEQRUZ+scuqNJT2OeIlNs9zoSzF0Xn
iPRWvxbP1a5QooeyWPcFIS9NTErSYoQFHPgk256ttzj+1FPfBSq3Oeubf+0ANhob
l/S/sRGtDlQ1/9zcc1Ea1E1VOW+eW16YoolBderz+b6YVb3AjKuxagGu+Sag+AcP
5sXBnJnJcQoJejIeAsVEI/v8/yvwNabItBWt64RMuyvnFHC2fHC2lqNifZzb9zPF
X/LpX0qPPS6944+z6t7Kdzy7GoExYCKhPL4hADCESwZGlVmVrylRsbZWmnO1Nyl4
P8ggL56zRUoS1H4mWdJ86aE0LLpOeCQSqDhi59VtP9+K+xpVnMHDCkRnOMQVRaKd
hGVUPfTbsAHtMn/vAe9zRHfB8lR4aZHaea3bON4MHJC3yPNuDejBJP5czrLydQ/Q
oARjoGL/NA3UjlcqTzEikRNGQN23iUMxf91JafjousBy4SwIMIPaa5lMkDPu0Ik4
y2ILqJr/VZ0poeETL2Hsd/0TlI+pIc5D2MArUnSiivL8mJ73zBcCeuMkWyA/ol9x
EmYJgNa9QVCZmJgqlNgHEBxoNUbfZZ980AFRgI3skAOkezBKYz+jsm58MTkQ9TT8
8BdH5nZHIhFcAXQFCrLSmnzo0D2hHyJVM9ArWCXIANy5Qf/UWIA3hTpXsyePbtAv
wAG3BFPKVa1ha4Ydr91T+uCa4wEmvZ97irvcvB9aElrJYMBKkaaDhyhnbhO52iW8
4w1CxzoYpUUUPCyuqv28Xn0LQFU0wD+/FoPU/iPkWXyUFJZj62kmZgi6ToIjm4qk
3ka6EUO2KBTpHvzIqMMLzgdZk5/Sn1+sOHRS6u349KXftd4rPpideaKeeuZuhV/0
8ZS/I4BMNSm5D6DrKpv5KhLH1Hmdu0OOnq0Ux9XdPGYYeb0wj5AZMK94g2VbHlze
chu2KTLXdriQyqngtoMoCgaemRL+QhfrygUCEtn4GrX97N/LJUqU+s7S8JQLc4gQ
xP8kZckvk7qC5TtR99w8mgZMwzod07Q+I7YEZaDFT0C3ZkAE4fzj+Ija5r1RV3ov
VhPYUxxKkkOR+IcA81Gy0x6+Ut8eMAS+AhFjFeBaO9IYiZCjCc3bF8HhVSdvv5Cv
v3qCgZd/TzgnNdo6D5PjvyN3Vs3yCvqPF3GBFJgzF2xOcQeFmv6TbxdmqGj70piH
4VCfPE2VE+VPsTQOHC6SbHnyUd2XvijSmAkSCug24KxCq+McqC0DQn4pm2L6KS92
FuafnndyRRfmjQKLgpJ67iNpqTwx7c2X2Cz0Fc0MN+ZVe034FtrMfWIXFw6XHGKv
tY0bJi5f2yQ9tkmsVytMb0y/6DwJpXxpO1j0kkKV09c4mSUFi3bvoABV1fm636XD
L1vaSw+NwxKIQzFWAtuKRbCjbUohtfU6tjxojBTF/AEeU/CkCbDH0gSFUCiaJ+zA
tRdr0DrsOLOo3OhJo/nkLgGHKgxrkCA0pDJE36smwH0dJMt8ucQlLjtOMobPmvIu
nre2s2P+VHM7TKereGJLdrNsAb6NzxofhuUcfcdDsr6JrnSuAc8k0K48wl+V7iZW
5IF8lm0XPlqRv/i0i2WvodlagXnKdp2Bf62acxmNoayC7CTT4tGHOvhByfM6MqKm
dififr9EF2GRPQhMiRHP8Ft7/3aPrafq6PB9pIwoWFe9OLteU+JQxTFc2zPPIIXT
iv9Fwe0ozTfy3MQgIiK0ksN6KrjvNCF83d6XnhuvR7UqgFteHi/u0DD3viqqEFdt
6ZXTYCFhr9zKyqbDP0UiV4aCaeXYjjdirh56nTmZVZIjP6b6QhtNmPZqyfRkPkfx
lB5+9KhQt19OLDYaYTZrm4wTDImRyDe7k7yJiPKKS6rF9L16V9qCAtRXdZQiAJVP
EbVIzqX1SBblMpNAZG5cxYbEa88C/+knYlK+k3KxEZllEyIViFgmHSpEqKTxchXP
d4RE/22nEn7r8oSibznLMoWGxBSMbIdSOJr7/qQXwQKnNJNVlnBtUyc4wmFxc8N1
WoV2jx56M85z4YeG0UgpMpcoj/G1YNlBlwyTatnYC4cVz5Icc+K8TPtqE4v/h9N6
KvY6niuHVhRrgXuYLbkCKCo7qeV7Ag4eon1Hmxz1a/1cmivOLoa6YmeJRJIE9M2R
1Px4i0/ONiYhFVHFjBawQVig3xFb2kWZCwJ4GQYFaq+frbhD8GHlEg3c1eK79EcI
EJq54BFe6QtHkVzBDxMIbZeeZ13vA/jQ9cn/MFXJD3C+uCCDYZhBxqP/ieIus221
DZcM+Kf02cZE8YtT3Ljzg02I2ydFmHQYqy3wioATaBi76j9tffpvFGlpbJF56niC
Srftvyr4cziIR3zmlMFlY90by7sDlcFdED4JhafFnY1rmZrEkj5wqgdUpDGNuCaF
G+uEUCfV9IeoAazoFfGngCIFOM4SULERW5LagliVWt/tH/uqu/vcX73wcQ0HIt9N
GNImSneXl6znJUKKDjDjfi3+vzqn8xhD/8vYkgxULWDuzP16uRATWS2YBvoTQSqn
5cC+vqr36dD/rTqE38oyuSMhBMrGyaCs8u/J8504bm9ZFRXtY8g211VPw50tzp/0
fTTVx4JNDxwTZDPLSR2llo/4ODCtGBum0MpYl6BWqe2URFaXom7uzbT9POru/AD/
gH3Ex9Onrq4OcWd9xdQO0WZ5A6SoAdQjljVzSkySz3AYtPkuZyO2mF0tuY963CCI
r0wQxCDcYLxT1P8TdVF1QeNsTsIaIwRa7yaWlCjE7BQZ8n6GIImyjihK4Hb070vd
d1z4tCvQyLMtp5JpC3ptfRKRoy/XJoRH8zHgDkfeKXizi940bmZZcS3tdNTT/mzg
YuHI0XzGyPZN0TbCbdzItBzas2fNdg6Yhr2SlVapao0Jwt2yc5ymQhBXCpSxLUNp
8TboaS7KSR5UssewgMj/N+LUcAdn0kOz1eSCP8OxoW2iLINd3HFclQSoAnVb+MeE
CjcSjUHIYaHW9koJKXuuVapgUYK6DMRhOnQTYP3ryh6eV21d4X7FcxXho6g47U5n
Rr3jZkDBvaqTWvQiX39DA1qX29sPEb9sqQZ2hiNIPzvpSIt0m7GBzcMxtMm9tv7i
03X/1QX8W+faSWehbkETgvF0Q7dSAdHOKadlEKKGFYkVbdqNCJsijZ9ywtlk/Wma
eFZUWGEzeKGIse2PXGcE974REldjDHTHWjlR+ugy5C+Vj2lvFpcxRSiJgq7xXvWC
nIs+oc2HijG84KXYlgFdhhQPDvgy79SZt9YZJiOkHmidMdoDeCHk0WSM02uyJB/D
lzHxDJSyiJi/7+fMsIId3MmAk7EJPTMK0/HOUOj2RCdQM0Dt1tn48f58TxK7nD/r
YMBrg4IHl4GrIAK2VqQiSJxSevrcXydbKZk9cyEJF9KEa+xyKXXttbn+Eqr8PbEV
N1a+OfeyX0T0f0AKO0Mw3C22YQ+xo6T2cgJfEJDct9WggYB2TKREOBKiPfw95I10
BZG2jY1UlgnHZ5hhdDHZSj/HouY2IEtYm+7uRVYWz1S/2jg6dw+uGfjMcQ3H2KH9
lckYhcfCfWaoZSMfZE+TISvHKXlfv6oM55wrxiHjDznVuxGo8fYeg0O8Oe2LR/k3
4VE+Sn2SDeglKLpcJm6skGskPi8OfdCH9p/2DSBA6mGu0VQdQhgwipiAMOqWLs6S
OlkOoO/WTBKnEvFdNJbAt3EhCtAnIb4IyK8J+ho6kBJ7xYI7djU6XDmaTLQ2RiQr
BMCR7NaPZ8O8Lfd6tDzFEZSJ7+HbX+8v5YsH5YSSP+lc/ux+A1hYGx+dTsMMw8Pa
rnYCQVpigOUKR54qoSd+Oj20nDx5abJ7laGxCuZ4NmuJBa+S3jnnTScFZSBMynWr
Dn+PiT/GlNcrRnrCnkh7sdVUJkfTs602TQFb/QgN7QvpQ0smJ7ESmEnV5/RDueM9
cqQUQSfAhEGxeg5s8OmpbPF/2FBTTKxS0HCsfP7D47uCjafMKNu+ERfLjKA3AFgo
ZotNtEhbS4+kZvx0n6H23LC01Oxyrk55iu4JHfJvdt+ODB4ZM/2XlCuJ7aXQ+GpH
lbslQwn01hjhnP5KncWPrQaG2ls2glTXAmpDPUwKr5v29SmspqLn/6xiLtw6yPeU
ZlFPkbeK9BbNHx0uPDYnl7/DN2iG1sjaZHiHJreJ3qA0gyoQefUuoYkYMzNgWF89
F07cqhqrrIrypsfIgekGU0ml45xbgYcyycDzgsXrsbec6P/wkiA8uKCXgRKHzIYX
/07KixHlnoL6wNEAkzoWOsN/GgKcoDQ2U7f5BeuofoEENNemhUN79r0+/f/8S192
fpTl37g2W8ZbB3P2evNqYCOdDT80NZ/h2RzgH+LAlyGPDzbf6VMLdyomqt5bw1TY
Rq32DpTfJApUEzbT0xRAcrNvNIHG6oJKLY7jAJwyE+cz2hFBEeZJBDxdDjmiWw7L
xiTYNWqLcqS8o74yGWfhmDltCM4oJpWkuOwxpdg56wXikzsV403G2gJQFZZiA+NG
1q3r8K63XOwArWFn6JccKjanmgpQl4rR/1ajJ0NP3/fLKoAB6WAiT+tslC+WFoT2
pZOewUc3Jd9GRQwmEd4aZAFgnNoxAOHWyP0mjEJI6J+JkTg0bE0GUXbQmAOuZAs8
K7D2alzaX8cYUkHfRXYZOlPPGpoMk6fd+QLxwqq5x9EpLb6ltSBjl9gOJ18BB/LX
eMQMN62udMcmGe1m5bj03/POb+WW3vgPSFZlliuoivgTmtL5Pnz4m/TZM0/wBAWY
0eU9DtAp03NYhBiaDY8gpj73t3qHCSs93i7fhnBSmTqOXwiSn9wNG4oA2cVQG4Ad
oD4NYzL+2uzhwVbhYQcx+26SLNghQRXPK3lsKS0O7rsUrCxpkgu1kDgQ8hnx+D23
YSWGJKqXRE+nvd7wAXHE8Zajh3IaI/MoTN4RAfV4vBd5ffvqWoRZJIB7YOJcm22/
O0lQu1FCb8nbh50WRPts5vwCz3XSYT3aJqYIrza8TnaT6JEH613g3sp8iW8UWI/x
qV/6j/PyHq1b4SgRe1tRqei9zmBDlRGyPTNdR5m7pyqn30XJSnxur7re9BckCggR
ng+L268FXKDJOrRuWZ8c5jrhX9vyW9fNrJntXVtSv/XMviII6mFWSGWr1zoWHuOk
M6dZ71RiukQOkkbOi7ZJk6+fnlONtxN/12RXMEul+4T7WYaArynpVB4KcK1CWuqG
U8KbodsJAzRP22I6uUbXN9rRCWWFtJBRGhR3rT/wxMqb1af8+P2oeuX9w/khNpJN
r4fFVEzaT0JtFNu9k4Ncpgdl9P5M3s9axOg13nUK7uiDwu+O3uS9gvyyAwDXleTY
q6TaCTEtkUe5DDlHJTSx/tUkbSb24xRIFmwF1pU0ABCAaZ77Urs7io5KgqWhwT65
0evldEtR9VAnxiPCJZ6B+Sp3bywve12fK60Z/w8EpL/FrdubnZ1goHVQ0xfeLNHC
hU0mUF6mlKSM369wpNe63ND0znDYF991ipTXxe+LH7yeIQvJinNUK6+Lb0bKWB6w
7mb578BsB9Hapn2u1rIFORAxncZiKadzeu0OX1MvossakoKU6tGXPR4hDPZzFWFI
jh13cNxRrTWIYhfawBWBN7/jZkTQsBJhJJcNTV8cypeonLkK1vMm5lIb8ZMwO1ms
mx2iPizINCL0G9hlyQZRgI4AfaCi7Bh/2X/HV/rZlZW2LPG1Gv9eaGP/5ylf5Twa
z9Wxu0hyOlBork1XD1nor/DOvtiPixIKjf2xz5cQ1vfqKQt640J9F2DnRy4sBB8Q
lMvnT3tY6AmdutXHoYgDYq8zPY4YGAWsjRaOoR/OfqE/2c6alTHKlvSbQseAy9TZ
jpmhExU7FO5+37pGB5phxjjYiYR660tC5Sq30ovPLMgm56JpHKNe/WevwyFBqR6p
ngn8CxvgJP89gRj5scFfgkIfdgIY3WIi5xqsBKBxcp0QyvM+/aH+0sDHByQtTmTZ
iJQ0k7B+aRAB2mKQM4onOyitRNjTHhZcFcvbPxfI2IwwBX/iPYcM/phjQp3WBL1m
tatsDZZUWE25Q1Lkk9lApVC3yf1Oc9jKlBdH6URWaj/0HyHmzp4m+oqrh835zg9K
s3w4sbg0Rp+ZEeuj/cfgfFJ+p8wZ3kwAsTvhSNEgZgRnuJuhwsbJEl3JTfYsoBe5
3qV7FuDsEB8xbLXOGqOUeZzRtgZbT1jHbLv7+ItwW9i2vuc5KZraTztq9t6uhT6G
n6IBLxG2u7/r9SQl68uvvRibKCO2DtXh4wckzTEk63Vgg/oUdSux/tLcLNAIFwkI
ArCjWz9XsLWnYPobe5SiOldD+5gmi3moFjA6lWR8nTO/K0r3SaW6NH5j1gndo4IV
tUIkXd37fuuWZXG1r3tkugZUj9UWPrCU+Z8ywT5OPiD2giEU2uix1MDu1SYOfjbV
afiBCdvTdSg0mNFbpNxcZlRJMbW4E4QVxVESb9Iwotf+9xPe3/WeL80bbXURCV3A
TC6r55bqwlej2PDJ4XwNq2WnC0so1CmpG8U3phcmCh1l3zCBGeECf3POxov5Aw+M
NBBBEWFT42+qSuBhxcCSC7xnAHjqR7/E9I6eu7ie8Rjl+SGYdFJwLlUTWOc/F40A
SIRAwtqhqu/6XriihYHFih1tnQ/iCOpMCP0qY3AfhPuQFP8HlecYIA8xhPE7SlFj
9KNQy5h0sVNRquyq+nBhqP/1DQEK9ypMajQD+x11gf6t98ZpTGDTyIqEhjkdH0w8
ap5s90vD/+dhxc++uZPFjdKhFwzTQe4GtNm84/CTsbMXM2phZGqiotYzvrusP/hz
OmxWFkjZnK/7OvD1nfpmhinfvuVWd2zWuxReebteiZSfiYgsEL6wMK33ElJ5FU0N
YMHLzHvQM3JXnqa5215TijEmyFHYejwzOsTiYWRvEHrcWtay6haFYtutuCyuzzNp
GmDc9qDLWTCSzSrp3pYo0/6+cp0ihRMD4FU7+U0MUFcMfgLz2exYTbGsGujSwKfM
89KCRqwbUf3eZzCVhONuzCSSyVFZvc8E1pI2QxV3tYJuh5s3CB4a9nFhRFJRa66E
XYhfMxzQLKn4vgaimF0y76xqmFLErcPPusFaP5imqk1KwFYG3+znUgrUT+XnAWXb
VUmWYLl7fwbkZJmEr0T8iNQV/L9CaqIBxOLuM7owt8vLk2ZPECaCk8EjOhE4agXh
osnkoGhDY9H1XLBLgyxAMcfWqkQaHQsHaFxjCYgH2FlTbZMRBhsiBbqrGH33a90n
JHoK7CgWL0te9ifjlmW4p9zhxfbha+6VkULVd+2vs3INqX7mZW5oC8rGuVovSCBo
SdBJ1jM94YENd2wa3oCvaScpcbc1B54ubcX1faPQe8DMvRjb6pz4P1oasnUDzAf/
Y7PMAbzPZAXNuzf3qbK9OIl4UmNR0QVJnmU8I1/Hlexd54lVSiO1TbZbjIoljG1l
9tIAnZEkayB5ZDwM/P3LkOohMVvPUw1ecG0nmadqaQN3uozo3N4h6Z55VPI/HOWZ
thVodugFGf/Gjre10i5s46DFtT1FyvjE8dAdb13o1xQGrcMTF9FYyCxLyQ7hdFdt
YkEZlf8+yM2u5gGkdMzUMKnVZipLsR/zAt8RB99d38kfqGkpD8HeDZGC1v/yYjZp
zkFrOhT3yozTN6vu250oxeG/9sWjDkaYszA6Jx+9X24XtYpMU6AGbATpv3u+TpEF
a4Zxa+aLN5be27aZKztTJOhu9dN3Uv2TnAnwT3x0cPk9zPxCz6ovdJkfPPTGXj7V
Outpge1qdkanUOARm4/kYmgLIdpVjnSBGY6pufMtenwiyGjdVPSnQxlxfZeXMpoG
bCATTa6OX2buIS38EvgeGNwud8m/YpLeR63da6M6uEvh19t0gRwoUYYVP9KlokoU
xk9JIlTUaCTDB8x8uaoYoHrFWnw7ji1IKWulqRTkI9BKHuIuW0yGzzVgDbeVMkNH
5GXZEn8YlyiJdv2Hitp5R3ynIyRglPZeNKsODs0E4p+QQqv/ATzGxpz394DgQ6qT
RQv+RsAMtYfriHJWDNdJSaLYuUvxRN/Ua00Y6JSdqMJWUMRV3ZEVpLS3+aA9j519
YlYYGNDVbdQ/EAd48d3yYhElC1Ew9aWqVwjc8uUfcW8+/UE4qvmfSucI4tvpqZSw
5RBVwxPA0Wkf3ro/3aQSQswVQnMnHNycy6TrgqrVPooTN9N8RcQ/JqCIm97fRowz
9wK6m/6Dr7ZYoLriVj1d4Hit2I6OtW4Hq8bc+Z0z+R8y3GlbI89i70Uqriq7gBfG
bb6NbUz49L421L7JoXIDeQcOVuhVlsbdNhRpsRaeWF9DRdWhPwMoSUtmRv6ofldV
2byZ3VP0uFF4D4aKUecja5wk1V7dTf0x67/Uj+u8PFb9CjRJ7DOYIMtqA8LI10uZ
cfI+11fPQj4epmaJbANzQ5zBxVIm+6JUdURNOVO7I4opr28dcB7DpjUfcgdU6jX1
o/bPg7D26MvUpVn2kRfuT+7RAz+XRIu9Xx9x9YZgzIF/cInu4UZjG+fPvnacFmtC
Q0rnyeHSKvPWq7UGb+KwPjiPy3m/t+Z+Aa069iv6/r6K6risN5boYg+1NiuGzVEf
orRTqWgy3U/D6RcLD0o42czP4D2g3E5y3WW9bFnSYC/IdRVukUSPJw16cXA4hBnC
9lXco5Z//AEdPeq74MEux7j9lI2VKlhYWXHtvgtomHiJSKqWCPNx/H43579H4O5d
3Hr9f0RCHlwMJbYv2bp+3Hqtdwrfgt1BgdMlEK0aaX7aaAJ3K/tHp2pNNFtCxTR2
4Q/BwEfwnYiuhy/w7KQFq8PO3l7hqRYGB3OOPg6bDxDcymB84DIH4T/Cx7jT9kc5
srcb5un6e374/uje2/yAOzTL0/Ge0yKSKa56UeVxDzL80bqE/N/C6o0gIeITBnXK
w/0d8RkGwYmhSjCTNRpIHMJUtWm+jkxQyTOD6pF3JUA5MMsjX0a4mWK3+AoNHIJ+
J9lZc9pDNqf/6nWPuIgiZHHwhY6w/yRNtV5amXe04wZekReDqaI1ufwiZUljmN/f
0FeM9e5x0WKDjZrLitKMqoe/FR0mQFTkLlS6Ozr7BUvvovgrqPf2Ll6VpWO91Guv
kJHsIIYBMOUiy8BaBSXsKEP43JTjZIEpxaznkEo+dAg8JW4MucEK3xKabiGBiY+t
cHtMsxG7tLN3Qj4uXyCWHG/+4aWzyKufwLflfDHmdgyBZ/2x1EaVFbj/reXZFZBp
XIL5xK9oxtL32Rm2xE5SXTYo1xdPGKCUcmALjXunOwh5eRwmK6dRNivOJ3e21Bdt
ZXkxbR7WkcjSeJPIxQTSNpK2apOaJ+uqi8cURtE0i0Towcs3PU/CzO89w5igINuN
hDBntN4j4nw9nW5v9yzXQPlSsyrlbJKOSCEv2Gx0sabHC42M5GoI/bkP27CETrd/
9Rddm1nzcgcto7pSW4kuHBsYM14FiVejlwPNyytfDBtbiw+BLvckDTSJeKa4F1Ub
6q85pMVyf1g9vGZJnVS+bDxFuH55ogyMItNGMEPlXX1Uuzd3PiAntWVNkx3KpRxY
YnHCFNRoKfNZXJMlY1ddNMPejFuzXYa/MzBl2FKers274QFscPucZOdfYCt9wY2T
EvZ68cY9NbFJJOqU9wFImIxoKKzme9vGUpVtEdex6TvdvUtUDCqvspquB8HI6h/L
vHCaCrayX7MSNJL6EC8xXRpbDEisJctF2CILn6Was5iNFfR7sbT2k9VLBlND/2kA
6iuuTNQVzTUUmYSGH4EymomOUdkXfvSbEbmJNIs+96MeDskz4Hw+IM2xaRruLfdY
dMMCLsUdFTQGX+An8UPJ47rDo9veNZHCTpaq9jlIMYbhUwtyqBXS7rQwaLel0E3v
c6jaO0lGY6QK3DV3HsIszveP6/ZT8H6lZ1Aj51+sb+PcjgZjK5UBC3mDapYx/8zb
A4rMY75sE8Mfqcch6Z6YL6YaUUek7ghtq7HMDknQi6rhEDkj7zfAYXlwek40kZgf
nOomMB4FY3r+LNDQXdyAZRCOW1QGX4rZdh3z6oF8z/5i5MWnX1iEprQ/IU3ILmHS
qYrosXS1E4MLWEATnuEETcf/9FLyt1nbYxAV8V4M7nT+4WciFmxLOgHMWyyRxIQ6
PMREmAep8qQ6ffMtVWW0nmmPaIcYzfsalbfI0dn4gHGPRK08pWqEteIkG7Iiwsvy
Vewi14ke5IphWFZ6I6z1bscXro68dylhkFV/l09kkwCdOohgHLuUlVXKOopcYUSz
aSpYFPb5DsxeNijT8/GnnfJmVmP5ycJlC3XGsoHeU5QtXpjOP1mrYSgnyBcA//XN
4NDuH0a2Dc2WFM7YYL4ZJyYvBTOidLghChnH5/rtKVHegx73n32VFMOLPBQyq1Vz
viGacc4ZL9yuu8HWCcYrHKXvMM7dT3A9UcjuqyEq0WknbjIOzyaPrDg6r5oBcBWp
zPAOyoABSYDhilbyLtsJLDMtxkeIm//xSRleP9HvP4vB7yp+XsWNIb0dBjyH9drr
W8tLkcUfyksrJtec079MOWA005k0LnZGUPHnc+wFs3Tdk0X2uLx02Ux8tkqbuWxd
y7PRjjAUBzstv22HyhM2ETa8s57cqphswE4qcVjat6PpJlCV78MS6kqWJsjdTNIl
qSZOVq8okE17yXhB0bocdEsC1cIqn+eIQbrE7WLkuK3TfJk0ZtJkXpab+1o079nk
xzVZf7J5TFktVmwi34NfobyIkk3IQRLrWgGBId4tu0ALyC8im4wYmMzL1bKPSbxP
ocophMMVxURZLEAtgeHEy7coQpvHpUo1L0ezOUNOaTY6SfA3j6TIdaxOYl934XZl
QNcYyNitVTtBwSrSf9c9/lMisrXgWBaZDM1viO1XHiYpwfBnZNdOMm8oLZHqtn/4
3i5MJPBeFGL7b21S6KZVXsY59XhVZbd21jHRxIqSrTj1w2oyY3OaK5+XWDder1eM
GSSMD9tlEcpWZB9366/spR8MfMrRiYkD31Kh8Lo3OfOQWok0OBEPY/MIw3Ogby14
r79JLJ/ew2GIdHdGzNMmoYV0uzxmGE5rB/S3AN2rA/WZlszN2Y0Ka1M4OEx7VijV
r0bUUlaTzmOD1yZEjqhjuQo/31j8q33cWzSlecEBUowXLjvQZFd4OM72r1rMdV9z
ZSxW0/Aj4D88aw8lv1zkTfsad+82FlK51jUSCwPlMckfHcbWTmUQTARljKEGTjj1
orShRnE2G6NxYWUKPT8hr+fcMgr2vsVyYjMnDGMqABRRk0vnpcQvPLObua3AnhJ2
rYJ7CiB+JOn4NVcPMyNBqA0yx54PZyle/Q+eLkXZ89eJezh5K6DSdJrdd3Pfd5IS
7qXx3GVHmc6L7Pes2lT3PNYn0Wn0CGK5MXpiEcO3USdaGYLQT1rdTagIIoynNt3J
lTLSqTXYBegWD/QYEon5VN8gsU3psbIVKalI+Ko/FsX3FFJRvQ5jJ/9+LG+GDIsS
AdtMyDKLepfRdXs+FTut2PDWVckcrCquAcXLzWjY3xbnMVlzY7PfPOCi++W7JkzL
KwJjyZVJEQziXFqMdNBJW1tP81J3QdlLUcyqGU/DZnp6gCpYy/9FNaeriihZ2u6+
9Pfg96VKa+qOcVuEi42cGS8c7UoZb/iMGrWiecQv45SEfEaohcdUzNROuaWuGrV9
9tGoFxV7R4jAoHKr1iTe0UiFoSG4DY3NpK7aZwMQULYS2rt86mOVD941LmCr9Uhf
RRmB20zX8VXSsOPWZxabr+NlaeWnhZcTcaB3gb5h6G18nAkJv6Z81ZuaAg0XFAlN
V29z/AOZpbatb1FzfwUlzBw9/vrHfNIgra0GyOn5QCjPCUAwi0AeaFeTJWrvkovm
W+5g1qixEL4SktenSwwck6I0BCCIyJ4Is4rVzzFOubvUApRDgMxfohnhQIoZ1u+Q
UJe4N1V1/rGU2uICAYh24iKDdkohPgKMEhKRULxbwcKkRpL0k2ok0cC8q8WzMpy6
SYnRCngvbOPG/tvu9Yw3tJewTqgX93byUoClF3+38/2pyIjxD5PWGlzTDm9RQKuC
eqwO4x1ejQ3BJo1iPwvMWzJMLxn8sSRRlhM7BfmZZYMdFuNbF2fRXja1CJU522i1
cOV8J6CmCjNw3aVQnDSMD4WD40ttFVdammdv/l5G2N1tBU88pYKkgwLzUTU1DwI9
h1v/inWlvj9c6XFM/9XiSGdGRDLIuGymmQsglCjKBwXSxJZmXf4GSuZpAi4eMhCj
YQ0l+UshLLpOO5TgTPnxp5mjWNhN0KwlLU+ysC0QitcEaZ/AvtFo+Jn0JbFoEYLo
xACo24D3BIpYvj+X39xjL9urq1yGZMfoKIxnCBpi+k3jcMM1Z3erwTjQKZRFpkQX
qn/VUYl9DY27UbzokOBW//sxXksfYRP9riodOlnqg6w2Lwcp+QqvLW/ZzXDiT82o
+s9JPfuH4p1mvA8zzUG5A0dH7cj+FNaSUC5vj5pa44wza/f+Ska8NHI5Axz/B+Q/
jD0I4oBDPaGbE/zNZTc0Z+g5E5FqmUGVX9qTGMarlUJuzHXHxLCupx/bKHkjg74Q
7QCm42Zms/NiyZ+5XyASvJQOWJXmJAnPG/8vb6eKHqXSPwhZOXDRavlMscHUe51L
DnG/x+dYELPwEQ5ApgXdZlBYIh5qZP+zmRpasQSljIJQNCKdif0Asf9Kwgp27gpu
vSjH2c919Ssrh4bgHDg/BoTTfvYXkAiN0MiIgA0O4bxDWnMEaVFhtDqzJyx/UeKQ
w1mJQnOsrzoTMGRgVMmvc5yOE4Uzy5M9KELCoHqFigfe/k4XXiW1E7tVcDu4csDe
WlgCYlfIrD3zKOuSE1KdC/PCDmy2PHPS+GNgHCTuB3fhiIxWj8BcUssdiG2HdxDw
byow0vXqepjcdDPkwGUz83k2iiGGDpVOsQH/l9P5W0pJnnSetK1dfPK2pr6sMdm0
U1tsRqKz9a/LCCzvFkCHa3y/wkE0OHRsRKh9v23CdPm+5A1HTRZNxuMJwFNQRvxf
rMvOJ+KmjBuXAXP0SBiqZj0SDjcgp3uBRG1e92/fmYR/VJkBepYkAHMmaANczILU
/qR5uS93/jW8JvgUCINOjjO7whAvQsLSXgRqD9j4GD9t1z+ZiIcjujoBzh5owu2G
YsOB+5w2EXvsAC1E9EQyxRy0QxQGkfk0E3F9d+NXZ9xuiAShpWoEMtsiB94/bIkW
F1583Z3r4HpVKBbBHP5Lc4BfyZJk4LvXiPKN1xO0ZbBS6A1oWYE9HfIMu2SKcJHY
a+qvAov2ulWCrW7ZkMbTKdQe0HGcfYhT4H4GISgR3pP7vm0Bop6T2BSKVSsRUqc4
w/JZM/NRrRW3Nj5AZMZInamlvXvGHJU6/NjlnO9WHTMoqM9PSLowd1JEuMK12QjB
7C1c0tsJukzG778i4GXDHggn9bflwJRJuvrz9bWwQLWrS/vAsruRYVNa3KK8/g02
heaBU2zqSCCRHmqnr6bQBPEI9TpLiCAnu9I0I+yWEXv+dXFpJ4w5qy9BFSWN5NQw
YQFtWEcwoeo8jWW7trx7f0HdqulZZeFxC/HayRHBavPOkI5lSx5PVLWificS6gH4
Tof8XOsDJl1/jGJBCodJySpQ2m1/Tw0ybAebgFM7ACWibsGqkQ0ojTQDjfb0J4Te
5fN/DvCL0DyUg9M8FRo02B5aptFYafV3KBPaIISdsfy2Qt10sPoLFeGcLwZ/LR2P
tjRkiBVMxpbNuwAcZS9Ys8jOAo1Mefztv47BxQnhjy3TVq6qCJKhkY/rwOfAdIi1
PsL7hc3qX7evF7ZIQfIhP/5OEGSkIEzGrya+oXyLKsD44vPp6pS9D2GKhC/gJulH
3r+aF0GTOUh+gJ9RzulX0fQ8EV2Sp8DYMg4DN3wkwwAxXM845zWTmPb7w0A8yLCf
md+awZXPII5flgcwJAaJ4RYnhrO2oGQBOhccmNcFjcHuis9GBq6QJUc8fGNa/I7x
aLIg6DiR/f4aiq3HJ3dd/BgV7cUumzf4p6/BKLvz7k+yFzlTvho9c/8soMIqk9M0
53JdLheNHdaGMKWklOM2n/KK+iBq69w5XEJe4UbWdAlglgOlOnoIixfQbSpcTiMV
dewjqjZDaxJmkxW1defWyUcfvMsZ8mmeqYckgQXuxXW+9OPqOfGkzycVcw4gnhsL
76SZg8PhWDpTm2ojXYUuCRALRTGMgOOsEl/eyza/VYYsv7jbFjlZe7PM0uTVjVnK
KS+t8s+jJ/G15Pz44xkZ9P13Ctdy4hzxCTYXwsUuC1HwPaYYGyhFKKAaZ54VOa5i
SY0GSLiM9/+ybC2XSb3Ryb1rveHdLb+XXNey2v41VckLOsAoFgyaHxI68O2S/mur
9rd61H8VpNZlkk1dibRcOe8G3lKCICLrULEt9PzlcJ8OYLM3YGJ631QYO8daRxrV
mQffj1exLn/4A7H31bWh6N4R+cLKJ/6GBYpM2fhz7d7QPsBlSio0ZxAUrdD4xowq
nDs8VL1/dSktd+zL1YEttzMejOz1cxufnZ+ohn66spTc0ykkIrrohsKcWu2DYNqy
A/lXV634gKIvimJxsNK1quo7QqygiZCVhTixk8IL19Dw7ytpnkOq2yCwqO3OFxym
5toNhSMdGLC3avlnNlIR8iePAdSQYdHnA9a3SfxI279JuSkQegrnuLtmNcfLc4wt
brgVjej9yXNRa5nvwwypwprbvhIU0SvLFTJ1/fIukMDxzsVMT8GScgvkRxQIZ0PT
w8WK7pIlsrDVoA8+cX26kKrrBe1lTyexb0P2XyHh6/J6NZfMtuo1RRXvvrqBs8HD
edMv57uPiYJr+YK8/TDq+BfDdm5edndlRKwV5fg8nHZ0oQ00TTjSKcFVQK3OdwlV
cJfv7yxTh9Pl7obhrc/Gflp03DQKqlKoSUMMiJmgU7AzytcT+dBx1k0MRhwmuwXG
hBObMuLX7u2zhXMzKMRX+ULovqQzry2CzdUoIMc0x/X4QU+fv3sySvlOdJnXNvGL
6JaYy2RfOWyYaVa4GqRukfys2ynpU/o3Rr8dVfbrVnZszZjlLOaWMqFGPKMwiJG/
h45LM32W2/c8QfJdzXFhC3qa+trwJ/Gg3r7vgUlpb9373B+GrHYRIw44cAZwdiUp
drn7yBbTQIYw72Lzx24Fcr+LowCm9PvQkURBdLgt5EoHFwOlML4jgZ0GGkIKcfrI
HRdWihi0J7YRvHoVFvOB61RR5rhthPrjjXuZ3CPMkp5pGi2bMCvMShFhTgGolyDd
7/TMys6VgtKE0Kb2QhkMc643uRmR6rPgIy4Q8yB96Z8QibEOgTWBDfXQXEu8/5ZC
2CpGDR//OzoxKspXgHSpmDQ3wv/zgl9gonYDqncqdT2llHDjCc7glLK9DEaQwcKQ
CF0gwdEqKkflnAeMbA9rOshtP861Ppu1XIk/7H+pNaaFFc5g2w0G7yzuy5Z6oCnm
pLHwBkKFo6Wf+r4eCazb5WqY7d1McfMxmAI+Rz3JKqvcnLNhfkqXkBaYGY8ouIqQ
J/FvnhUZ1cLquz/VXE60ZOanU9PRW0I1QMljVLbnrQMelia02hCOsTMvRnLd/4Lj
AGGNdorNZR81PpRswbo+gjL3jabFLPaiN6d+iw0GGE2Lc5aOPTdRGNr7Lt7hwNKV
DXVnLjV2jGY4nCxRXizDmlAlcK/YMWkc/s3Y8pxrWdiBOWrClKoOoUmPj7cTBbsg
hdkc8MPYoxgMohNzwTxy0R1WugwlcQ/7Q3fYWsfLdVJXR1HajNAfcF4i2AJZmXEG
65S2bGO7kxW19VfHPuBYtIynAj03YRFfU/YmNXoD3rCOsm1bGgGztayxmEp8q8ti
If0HLeZfbsA2bkBEPRiha4zs7tJARY5duGHLnIkb1jD+VouDU7ifMdIAEnjkgLS7
YcP3ueJ1TCZm0m3hWMaPwUf/9inUWKXoHbqtlfr7N+C3lemdOzlWI4IPj3co+lGw
VUYp9bRwlPtZpgNKRU5PhESXAsebQ29FjrQxjQo4ZlnjxHvbj205FJnMbKMgVQaT
OvKLkV0IgA4jLN0MsCnQV102vwOR6Nw6sbZxXDdh8wRUK0/b6ajcHR0UiWxx6P6k
EZb4qkOmXXi8n7VmB2M9eCRzudJ/rMZ7D7//6Fp01CpuE31AqdVCRl1oYYvheixU
CsEkkPd+oVFLIc3e45jxzw3yfIPC4B2bcohR7Xg2R0T2QeHLNv5jzL4MWzHcth4A
StB3vbETAYOB7SIqjd9HOVxX34YpOrlMyX6rZmqdqTvcQArfsuhRY0Jb4Xw6KAfl
03akewsYWBlk7i1t/Uu7RHKzWgAXaKT6Whh71K4Ex5nPLCul5Q1UQrsUw6iOcpcp
o4lH/gewV5McU9VITXln3MQPhIAqTqtKy5JZFM+PUTw1PbtbMVSZAmZ6vLpYhzCC
fT4j+bEbUgyg+msGTRYaxWANtWZ22oubCwZT3zjNiLZ4qMwJqmaJzkfTOQKCAZvU
svG6MBncD6283LeHhxKCI3i3dfJ+6AQ9tdpwfd0diovZJHYVLktRoqZ6D+ha2b/k
f8yvzxqmM0v2MKYge67slxNOCYpbVMLFqg6DJiH8GwksTkW30HThJZ3SJTZUOGkO
d0HFsZre6VdeQRw/Tu5sma3JY6Pg3WCVarz6mgstsvfyWinAy37RP3pikQCh2Bww
ncz40ZRGRW1EsC6qXs+Z4TCV9SLPD321LNiNxUIHNZvYFXorm66/HOP3dezmwE2X
sfhZZtXyc1YgDE8WKVJb33a0WhpScWlT/LPKJAEAzk7lTTqXPwcI9Q9NO5cKIRal
oDwBt/ENlNBajGZhNaCn1UlRHI1im9NYYhTc/6cspD0G79ulfdskWm2pdD4NbnFn
SuYUn5Z+470tvFz+JcPOJ68Ad0KlJTgseIfzFOa+f5CpDmu85dvVa2dQ43cPKWlc
EIlJHs1PgSlJagWYpujiBYr5sdUwbvvY1v+xZCYyLVFgSagHbXqlXjb7CCzGAoRO
ZfClzwWllnZUSjF2Pqq0+khnFofbON2NS5c+8O34meNNW1yL5rLJimjufcCNxYG8
ftUN5nJwwUyAE6n/v/rf1IibgRMLK3TDsH2QvJk0rAZZyiUsk5SfV1FYEEauLptd
vBrtZY339S2Bf2Px0K2WM+hX/28Yh8ezcDSJtwXPy3ZMPUnCMeJqcRqUlJAxoCH4
3mZe4ZsBhlAgyTRjSPAyxArLyKK5/hPGtRNizeeMbR7X37PsCka54geg05M3jVuV
qXAYrsTEhVbPY/+OVRrYJzj0iOk6Tvqk0n9oZrS+SsKvbra1Cnz2d0eWvFU54g3g
C4nhK+wEC8VCRRBwMbBu/1c2Orj1bzb7TBwY+4GOwnvu8dW7CJykRsCY6DkKhL3o
vJC5PKgfcLalFzx97xvcJ7iuqO0myO5UshAfwDZHPccBnyuQGkJdHQYyu2Ji7EMn
j7ssaEjPLVZAmucqXrwtAbbajHyGDAnB2ef5tK2aALE0AqWwn4240kPRXSU8fvjF
QE8PP9BHS+p9YrrvuCPEg0My9KeTFBRpNnfAKowBVZccLcFC1Kz/vl7KRCwQIeZ8
v/ZV+VszRypPPeH2Uo6vo+wO0HhMMQqpdPWfPGJ3hqCWdhGokCv2oLvBz1R1k0e7
2j++AApcNI9XYI6dEtrpxJKHqw3hFX8QV26lXt3EQteTUPcFwylUjNgi7Vj+iswZ
flIfILpI6IvT1t+h4nHwwn4rBeKvoeBPp/g4P8nvh9LzPyQ9uTXqNknjrGdY3mHN
WKyqsga/WnkaqVa4t+x+0IExakbCv0HYXPiE8bYHrFXJ/mpps/+CI12jvtrF6g+1
ARDOD5w0J07OCsydBujV+TunxtP6U6REXgGwAuINVF8YFIi3EfXmg8TwjqkZvoKr
Sd9TkfkBfW4q0hAxuNwKcC/stuXtPMa3gC1xrHauX9SJA9H7z1dssWuApbudTD0G
Xcw45yOOlwo0AwhiqRKA31Oj1Phl4z8DGSOQi11VWtzocpPDlf9oS95ZgKNJ+AAP
KKIhrljjUPZG4nnzOeES48H1NqdgknwbN8iFJ0BqCpqZ7Yy/Z7mehVOVS/0ITxGC
SANP4XNVXK4OT7v56zHthYuTd/0B+OEoBnWWqD0B5M0dJwaaiCMfN0pq2NQUuhMj
S0Enhd5CXWxQG540LsJoZJ7iPRcGGeuFhPBfD/f+0wgVEn4qqJaMMRbjZpJhNZtT
pR55bGL8F+Y5z+VMTalJO60T3swkCoRwei47Z7n4gsNVRgzVSUCC1d0yDV/Ufbri
QO8lfjimhpqRZKF47uXGqftde/afltkLuaB2FoJn9sH/Dv/+nZ+0sfisfwzvxOmY
ea4iuphBw8zjFVO1hkKFW389cYa7+kc2iGBn8UfCe67TtHzLsSC2QSi+PaJsII3D
2tyQpvyEq8a017fPHtJQQk8jbcaybGpMHl4dnKWse0svbb0cnnUIgyoVgmlkhDyk
lhJrDzgMvjX+2wAAL6SzdtDFBO3eZC5HL28IFJogIu+kOBNHhN4NuS5mZ9yr+kTt
NbcnPxBQ/Yzkrh2LgGOXeCeuv8ee7sPScoh5pBfT6HhKXN++iwtsrh5Qo4yHMkpm
FhKLXZnKwH74EEdmb3Cd15FUoRb51OurOr1mbFGht6UAUviXxEzOZYYLsZ+RfS2H
uyZa3FAS0S8xF3eJ41tYy/nRb4bhs+n3w9zWJvnFUuuzB7ZLoNt3HKrzJjsmU/id
w8M1jZNbxwnRJxpOEuw6RG2lyjW+PT5r8oN3jyCxeSOLSAt3mH1x71OHOtk8M0M1
3YJg84PDT0STAeq9Xys29LASp2DlVew8YnjiOK7JcNH6Ob7OL18/PFy93ySlVpsa
kG3VcoC2EhQc7uGZjdBGU8B9vpi1TeAEZRDJctHeCdAi+tNSM0DpyLO8Z4D7RbBz
6kg48FgiHAyC8nmMoR/t6SjK+17RbUMpqqpZBKoP35a661q5nAfnneblSs7i37Bp
e53/jodfx8CZTBQ+mIvJa3sE/ms8hbmiCwCVdKK6dc2YCJPoAf11E6IfgZg02hN5
07LdYX55/ATg2pBcjoQUVK9SiLW41ib/Al2ckVCiQiFGGPnW2Kdxm3sPqRzVGRlg
foXmScZxe0ZORI84r88XlXH8dahk7jUGdjcbUVuUt5VHo+j2O2KlwZ4TV8PkZgRm
mV1cqVr4a0RVIGxKtZUp6CiBW+HAPDvpg+FMWAqHlWG6+8O9OEBS+ZPI6NEFHpEl
oTT1Xc6z8Yrdc8g3nzWhd8eVgHmZx9MXF+VPx42J8J2wondV4G01BvcIDItEelaw
w/pSzX6y2SqFYXGkiVqcZ+zgkzBqv0rhuL+5XdoWDbSN2pzJ0lCIPYlE42+RUmZF
RvHgUobEerYIR/YGOK/X1C5F2ij8jZwCqKVAejYYyABpA6G0j9BPrhA5EZpnGKaO
iPS0RmpRoUt21rSf2oPlgSa4FVpOXcQVvTNVVEZneyOF7Yzl6z3h1sVFn6kIstu7
GJTAIoI+0WrJW2g7NgZxl8xzCm6yGmLsSfFzAzN+j7c4m1cLDTlYoR7LEkK6M0JB
YLZ1WDvqY7nLL4ABS+WeFvzrUpdE1Vm2+qTG7GWPbhXoCTZSowBVmE6g4vVZMM2U
bQP3m6l2ZUaNhUuLWjAfSt31BOjV7X/uugZwEDkXUW+WhQtgIGFjwzKSuCPRtmG+
KYfHlWnvFNrraTNax8LXYs9e4s8Wt4u+cFq4L3aQVatBQejIfHL2BmRY6X6SKkq1
Grxkh4wjeILV5GILMRIpzEbmSJNFuSK6GPWYrjN7Hnf+KaQ/F7//higwe9Gv1tIc
kn/MyG/K4ylcZ9l0DAKoLSeVQriP1kaE9hSMqvh1K9VrUDPkuT6wPmcqAKD28Oxf
liN3MGSMl7bnoVPbkozHHnmoyR0gY0B135RoVLdI/vXG/x18q4y2FN2c2XJDAuUw
fdXK7Yeqr1M6zeM31WZygt7X2TS4/6iZwwUeu1wx3z3KQjupqOZ92TQi5xogTwca
8fn5HGUs7VeNncLh4pKxZ2YB2osZfIeon2NXsy9H49k/lYty02DVwBWTk1fKUpoF
eB7Mm/Z39S+PtowpIDLn1VibFcyNmVW4eSx4i/4GtG3Rfl1gskLrNJbuBnw30+zL
5MuRnoAO7R/pm+AyV29howMJq+yrLQ70X6tog0mPlzDhnAdtzIKBO8dmg26ITY4l
+bspefuKwFeLmJhhB+cu1rsMvAQ987W6bxvVQYKbrkwhFHuH0FTcVUUwEIhh+1Zg
+3DOl71qF1mZvAe6Zp92MM+hFagZiwKcjFPalvhSJFDbBbcEHiczC04pPgq5ExPE
/69Pp7duj7Uw37L+ilNm3A5UmB4qnJLdeIV91RVZw9gSdn/NXmK8yJTNkXKUSFXZ
pNWHjg67snlHum3scjcxn+OOEgv/GdOwJuV1cBu8FEWqg4HGJMwnk2T0Ow04veNb
sHDwdw4OGzvb+5MwisOYWEyrhAa6s+L6AlhfIwDg/kNz+S4F3BMxZ0zL2jMkw/5b
gqBlkC2QaLo3P16piwQM+eFM8oQoz/1ablM12BUmrYNo8xxqiK7nBFqWIsiMTPDs
83xXRVsXByb0ExFgl6auGeRF5btzbPE9kh3AkAn2OcCCZCF92tvqFEnpTHbgPFgL
6LopXRR0WsZk1ptCt0YS3aOJDna4Km6EskBX+qpJgYhUFACAJCty0UOUfuj7icZ/
NSyaehmemxkFnKfLY8FPwh1p4wWvgal59N+S22x3TvxhDOqLH1ntsvhI/eKkT+36
/ydq0Af6SwQNR+DFhqt3lqHlHGDqCe03ccQqdLCouo1nhC5lRQYmetLHEsxO9Z4H
JSBd/GmMiXHXxB8GmZTNqgRvLRHV7LE3W00CLVSqz78z9k8vpEEcDqhiRNrkfJz1
dw0QSTSRBas93ehjkUfR74QBs5G57s5fQTudB91rAjcw02td8f1+WrGpukhdHGWb
PPWftnOmd2hEQjvzI1Ynh8qAgF4bd/RqsbAqIpcoSCr2SNnxf2sBtuChxcqoqY/K
DAdcsqwyAsTVMm3TYW92fF5muDjz2hgz7Lmt8w6dAVJmH260srrpM3hVO/wR+qya
wVg0p1EYF+i+UGZXOyqXSieM0d31zAHrDDtIobIPepwwe9JmNk1AjORKXkd6pp0E
+Wz9gzA51fKIhjqs09YLI5kCetQiriDsboICNgqvDjbbzNbx5nj9PLi5xeZj8T3k
rmFxKOrM/f+KRjuUTF6kc0hOoRvBU8mdp57wD49hKRPV6SIA0Uwjz4IgrDjc3eFU
KHn09q4JbYsjt5hPmCifACIFQLvwHPFuvJKj4KJQ4kXnZ3Gt9Jau9opF4Wigio+2
iWRH9++jw9A0lfWUYobPhFPJPRjtCC/mKGv9nHqbMaQQnVK2dq+IpUyUntShGy8g
tSeunHnjz+Uq3tfJ4Y6xoubNzvTpfI+/3MWwcXJjI3X0ED2Bni2EBIwOKQc73XFh
tma7bNV0hfNlGUBBOqCbr1dVX/D4RClxZF/ZlykpRJl0hiP/r02kHwI1TKNQ+YjP
D7FPpgaiIqXbqxx309iLnrxNdhdhyL5AEeYHhnaJmvGzVct5MuLilDWKqRGbyJHo
xi+5LPKWI2Z3wT2O3RaWZHEjr/y40eQ0LcBhZHu3D0atJGTRpB0ppO5cR9kyRqn/
JuCkK34gPOzlPNJWxPI0tVjPPYgfuEMSkN9LYvA/xFeAP6y07MCvwKI8LzYdTpjM
2qw66QrFTD3rhOSBqH4v89t6gMExo1JNk2gJ/m1luP2prDYIJBn/ianGFRw9ZWMR
nV8W+3z3Jv7Kk8eLaq4ufVNSrSyiFBldWrTpp2pWI6lp8ofvVfYzDFOO/P3coTQK
DOdaw193WLxtUvzR18Uv5kSCuyCjQePU0Fft0yDivFOW73+BH1yi6Xj6+fSWUs5o
gtiDd0g0Apnd80QGX+rBQQms8whvzrKJnUHHkesS7t7/qLAXsenmKFKUH8onjUmK
3quok5BS6zSxuRNz6fQWUEZAqMABVLeLIMFi5UZnq7zwze3b/7XaTJmjvDmA9jGr
eUPVntoJyoBtTn7KIaK3DSaq402jtvUCLA1e5kJDMiRZ3+EgCimOOBc6vMbwZeS0
T/3eKntbsNK6kXTCGYZje0i5+YQ6S/r+DeSpnXIrnyFkyvLwc5f0y+Sy1FOQQU46
zP7G7hEK0lBp89xcmn56rAAn8XA07U+/aXl9FAI7e+DB3mmHvYg+Bw1XxLIp0fYb
JnlBePjJlYU+bUzNk6xxJVK/YOBH8B9ntmRn966GxY2fLAalRcA1gcC3wVukMZGk
1h4S4HEkffkVf/wVfPq2/TdKC77ZT9j7/2PUxR/qvYzDbShntteqrnNgFKOMbDGd
zUQBEt8r+c3u5SsCf/pg2Q/9peQwMBVGoA+9Sh1Sw56WEFRGQAYWG3nKwx4WGpxa
lngyWZgDnFovY5cG4ZTMGtYtx3PX174tkAtYYjAQVX4R7KNAclbSnvIKblE/h7bE
o4/ysrn3VPxs/LsNcFSBCkdL6CIsmCl3/HDo5yvP2cr/RbQ5i9Wy5Lhwqi7CDPo8
S69ha2qciPm0LkGIfldLX4gPcP0WdmmaQlZ4uXpsXFSr6rK5vZsiV3oKL8l226Mp
KrU7r+WWdqF+9kv0lKbJKPaptiHxs+3gbudXiz6EMVgtMoKhvTc8UYAFjiQypJfi
p7s9InGhqIBRnEJ7GGMKW2eUn1IK9IdmSCJ+UffGMoSj0AWEJche+LyUhJXZzCl4
7cyMMfxP1Pu4alzFOSkPtBi6znT1g8atfTYlQumOnIYQa3RmThlQyzS3icUbQP8w
fznzWPw7q83zTIbIw7/ty+GjpoFNVe2EmLef+PuPjPifnK8JqiI6SK0c/FmBv/sE
niq9FnqIHy2kRmXCHjoh1XIu/JmuXTSiW+nq+9bxdmqd77hb3fbxIFYfZ/ZUh0ow
oh8jt+oP8T7Qh6LdRS75mwnXMk3hNGplyJiOoVh90kS6tAanMw4vUijd0ThIjzLv
QJlMEVnWGVCVLq5Kl50qLy/is+qPldV61fCJIH51J57/XJcHdGyH6/gq2/eEMK6x
wOa9tXytOuyPyZzXznIOmCHVNqgM9Rt87IAZQf20g4PPLVjOJKIlX9b25xYjffvd
4ubrKwqHiQWLU+Ec3GlSdNyFeGkNTGPORS4tA2aSs+HXIubpjAlIXdDJ6ToUNF/r
3jfg4vQl4/ew2PX+Hk2/GnUouMP8lfntRffINP1QAfR9wYyVbn5bmgSsVG2kq88B
Rk4HqzdMqRbxkeFtaVFmlEkOV1Y0sw5k0JD/yYFOTWFVWa+1ZpGk3zc6COLderON
a7djuwHJQfzbnBVaf1FpE6zLKMUvkq0B/aG/Dnlxy6b/JrNqQ3u1EFLB8+G2AJhk
kSs6yar4t7VvQQ8KP+cLQJIrBuDSpG4UI5JAXyIC/U6DAAhskGQzz5g3do5z2jzG
lXDH9fI15Pgry/yaP6Wx904UPzxbQfAT344jwAVz71o+thEXyGu9xLEYr4h2lYZ1
Yox/yC3aUJ4sFQueeO0+5iQAGGBvzFupEOcI/gdNf+sBhB2Xxo0UIUZV/yn2USZR
7fgfucCO+Q+hElT8zHYED5dJsUEP4LwPDmKKwIbNjMzm+A2o7kiG4L/KFniq+RT2
1txFo18zGRYUJMpmGprqKuYVGuni6LXH/qTUoWNXc99hnDWgGoMr9vmURTlJvK1J
MHj3avYWdzW2SYyb3s6H/1w6zRNVp3i+lM+eiDNOaIc/lnp4j8+OhLzfWZrlNm1r
xpkwTkF+cahcOjc3gFUsUkQ36E95/CwLhDZz95yPprJ9mhPBcw9gRQIsgd1+LChU
zpLZQ9m8qteCMbKVdlTnJ3tfj3Sd7t8B7IPVI1uOQ5Pnl18rGszal82XBt8snV60
Gc2Gu3VMeoOh1eSMejUDOay7qmrbZ5aXUPuWpoY0aKzIBxtZlfJSyxqR6OMdyFtz
6fEPp3wHi8l4TWRDX80dDQxDFbD9jzXhMxuZnVsJjyJyOtzjcyRcU5ZhHDcPKkn9
EClZmPOJlNsWwfLM+rAgZaNWiHwr+MJhWTChoihJGz7vTGI9pataC3RjzfraPQkn
x+KuGGogVBLgRWKsSTeccOZp31SObIu1T/9XF8VhjCvJL0r+/kG9wz2T2oOybqKJ
71wtU+RImy6Gf87/iNKlI7xJrWn18eOmzE2pyO5NKZELBzcGEzRf8wa5poWA1ZbV
3ovPn/5PYs21KeQAKh2CDpL1Par6f8Ni8G8TPJmkRzyhTf3GlZ/1qrYcqX+cYwoc
e9fyb+tP/9xb5CO9l0gZRudHFUeQmm6CnF+ZzrZ3c3sYNeq91QpPlnxNOXuiqEZy
nSOGk5YpcEQL+UqPzW9vx3h/kigpr7D5IAmDJHVsjAKG0WBqpqOj/GW7QBt/Jbfq
bn4bU1p857Ez7etF9Qdqt2NjYZK6C6n1O4W6rl0EnXR0AEgdLZVl8K7pqmfeedMi
+wFYqdL4Ly3oKyuoFjsuMclKuBy0qMjElBuzLV6Sh56SVLTLublH/k5krO51nfRL
A0t/mqs1s8Ojy3472R51YciDLtILtOpt0DIxsC4Gyn3No3pGXtWx6+C5C9sZY6dV
eGYb7MjYUFM7/Lh9XKwoCTntjbQqaZS94kG/xepYmKkudQ3YKph2TQqXJoGUzZw8
O032tFfSw/ZSREbPkXmfOM+whLcU2A9YTqs41I7ZBbH9QCc8+TmTLF1uOOg0Dw+I
KKl1iM3lvNDkIrzcO48PSM1Smrkb046yIS8i2XeTJRpeh4MUSzBT5ZdMgMjEGszI
Q3XCSMb5MfezSGPTay8InqCgL+Z39mvF0tT2WWGu4R2R6T8Blje/TNgRVpfeqEWm
lW/0E1EIaLTLoPTBFWZGVVpx6+gAwRHCTzXFfuZWbBd3Mjr3hvZkSrAukNErUIVr
eRm1D5svM75j4dgSHzp8xDxJZKvUeBV6rLyjybCC0P+dLjeWXjvU53q5rG2pcZeb
taBDkiTXJY4bcYmVmzwOR7XzmkpVa/IVCFVA/BkPx2G3M5/LYEg4FpN8k5k6F76E
s68NKQUob+/b6sJWRa0Jv3iw9h7KTK2L6t/0K0Z67BevHv8efSGjHGw5w/5tNkw/
CfT6e7+yL58H7ynFvdx9XYpF09/zf8MT8YN2S0fqabszJOJq1WHgZEeYf44H1rIg
xdspO9WR2nkcd3qcGHk01eMNncJBArBzGJpkjVRVP34c+jGMjbJgesfj1U/eU8ti
bSiJ2UEkrogfnxoB063TOLa8bqglWLP+C9OzMfLmNBiqCF6X5fb6Qgc4Cb8FneCm
DqgQkd8TzbQhdgoa1EeMbHiBlpSQvnr/dsUdH5zRm9E9GMuR2sWFHEMhuYtOkEAT
R/DANNCVZr9Q54Iv/Q58Ru1tuii1m1/+ZH8GJHmv6sgxzbEoU1U2MkzPF3LJ7zMN
jbBAbWWq417yQYAUcSa9Zm8cPnA0Ybd8h1X3CGufDoOURtb28dJA5HIAPLNdN03V
whglKhZWGRq0SwcCAdg50DHcIvSJl8mup0L7DeV1W80vgs0taKjqnTGMVlxIk3n0
G4bU8soKXgnMO04nBVlMdySGNAfnYU7DAufd6yipgrpw5On8ysfuIRlVKA9q3f9e
qx8d5B8SAjCaF4rPCjxnm9mxj2O2Z6vSvQqValJV77iYkqEi6YxGJWp3cowIcSJy
cZrnoNu/wymz2JmCywuJl+u+OrN6djX0wSJE0O7i0evCR8mRZO4scvKn89Rj0Gjx
0kcm2iKNKZ4CMEDrgXpX3v+Y4x7qy2rUKpl8yHhzC4nB4cxgIsA35axOYfjHxSOC
HUZUsw5KzT7kSB4Ur84llpKoFtchjVo/GbyG/yZ9uo8lV5NLwjIl2IKkOsaCA0VS
ar8Gk5ZsUCO8lSUoV3mnnMwMF5s7qxNR5ScANLpjSZpdTAGloLrjl0GwULBLP1iH
eg4FVEoRaj1dSotf5Sbg8jLqLeeffSNZMnp+1iwgmQiVm7J9SdUJm6ngGX0qyrgG
mZ8tGtMvOuRGUKrsHrpT5Z27Nz947i4kV/Jb8S/1R46GrLcM7NeTPtqGtOG8+JDf
Z9s+DmWJp9L5MKoRYECo47Lt3CqiPJsEDrKPwXas5HB1OXcYoSPHQ96JhwiYuRdJ
V1w8KKg1BYz4js+WxtDWPZGd8Rq26kW+JfLf6cKoBr9h3q2ydJMQJAHzvGu32l15
O5WCx6ezC8g1SamrlWENEXsUvf0NW34Oj6t4GpoihVCmKUpXlmKTY9k6qpuJQcTS
b+0VP2k5Rt5sesncDknCf4D+VZs0k48jYDgSvWpgxPRAelhR0CAGm/+W1DA4maVs
ymobBaqwdKRdCQ/vnEa2egNzw56o+GYph0A86g/Ba9LVmoWI6lz7RuCDQGWXI+d8
SFqHyqlknrHYz+z1jKZ3o3isdwGOqx6hQRmM1x1ZNGO/zEJrY2UEAjiUlRXkO9xp
MEis0pjGbdoqxH44jd5wJceQZiT5iYVmuwWBsjpDTlTSDCI5DfVhhll6fBGbVk0L
iLB/H2u3gCabBouGbrMtK3NDI2odtHzFkXkxaBecHsi+4iNlvrLobMhUnZgWipEc
AvglW+PrCMkX5tqj+mweq0M6K0ENrt4n+TELtEWKUIwJ90WI+lJWTCO8DNX5IbXa
UP3txmEHQ7szs6E3RUOxromf5yT+RbdLgGsHcCwIi0I7XYfEVTSY4cMRZw9nZGbF
L/dlGNR4DN63LqEMdKa0A7xIx8Z7n0YJ4UcNtY0J5//MNCxvY/OFwktlL0C5qzTj
+G4QDboK6Bw+zy/+ZKqmaeV6CSYpy0VpJi6eV8GNLcG5GrjZLPEqH5HwtRlYohfR
Omzv+Pd7xB51UgA/XauMytDDCke/tuQHKXtl25amkk3R3Tx1udWHF8QUCAxzvbYu
u5I6f9P8hwXrT3JoOJT6T/YZQhBBU7C/0bgQR1UKSOLYkb/AhbZaia/6vFz/mW7z
cTQ+C1EHHLAkoX/yWavaxrmhsV4GfIVI8A/nmevWV+UuuNtUXgL/IIW0O2ZfbnWk
b3+wqJLkZSQtTmKbOuRuPQnbjWzM3V6NMiS0JBBZbFczgSM6J+EyKP+iaZeXm3Nc
1h7H8/zszLJw0LUquZ4nEo8cwdMTX3y5ie+7rAJgQEDSraic9bXYi1Rbq3G449h+
mi8qpTLlIY/flx6zaWjBn8OGDDFKumvcwwjEIS7iOMyuF/a76ZylsejpKk+ZkDjL
XPa+Bmc4biCpTxvfccyAQPEUmfx8T36CpAbyUlhPhypqpIg/+uFhkwxFGgzXuizV
VRoevxxP4yEexzEwq5aEUfRf3tSEGgDWE43qTeYCULltFj0JegQCjXJgfAmizzdU
+o1Zd1hOOrd/F1JxPuAdewS6y8TBq3fpH6JiIJJH1MOU+z+/JX53DJ/ImPb1vk9Q
4B0SwLRRXOGiSqB1vLCyQL1fBRLNd0Mqzbj0kFRz36TBGRuiH6EzjMgPUQvSlwCv
pCFt0Du7nrH70SKrxDkThR03RQfgCEj+Dam35Ps3ZNAtqrSNO9sIicjlQqgfTa8n
BNaCgFUMXaDgl8G8aqQOzoX/oGev0q1oKR0sugubb7hHciYjKZwXYrgFO1T3uwjP
nXhdsLriOGO5Fn3J5dle+jnTN8a+36LjI+D3gom/pyM8wO8ddaAp3HlfNaHWZztO
t0jnuL6uPVOMiBC44QyxTVyA3W+gdEvfATJKEiFooagGWn31HGsuAMT6Sgax3ou5
NPW8WV2CEz+5z7l4YIfam2c5RvYIv0yPUnJ5VAN7aL+u+/7jzVFIgOgZpEtqJTcr
9pPAhpe8PCaL54BR2OnxvjnkyayTlgZYL5t6hmOx1xfDkkKlp5q0Sdwhe6/DtXX7
U9aLZtt9MLAJpeucDhcbBj5VAn4lL2H9N6a8CKgmuAfAUC2mYTThJBLOjC+n/4Dq
UEjD9p39yxgOosHBjegPZG8KRKs852afIk0cQe/wM3xa97f/uD72FgMxXjZ/SEcS
HB+WQXzvXZjKkMs3AAzPfDoQlhnEVPfY6SS4ZQIcXhBfJDxoP6bOBTGa5srOdsKt
VjxJWdVhuaS7smdxyffgypOD89T3mb8PRiXYw2S04oLeWcjtt6kOu+i495ezVhlA
sWlTXhOZ2448lMFMYAR+Wgl71gFnpQc6RCS+UN5zklWSkPRSKabMQvIDHrdZ1w7/
A6HPdMvAx1ctpKKmor3YfO5tjctVf6ZQDnYVgQ+VLLGkgVn1xVEeiLusKlt6qQCB
OH/IkIRQrt3ifdUZ85C/VL/hkz2wKegP3DpWO042lwMr9IKyBK7ltpbqNJB58VQb
ih1VRBHMIjppJGGUJFNu2Hzi45MfN9t41Amr4WwPt0v9ACCoo61r3CvW9/3EJhZg
457Dp0QJWz+CYPXBGosI9qzXPut1EQQJgqhjZ3iJUUJeJU98RXoArri3u6YGFW74
IMBXcgx+aIEJyNV2smcBNkH3+Pwbm9KLnWz7dDEVlVyYOm0bFcXb9GXuRzVbmJMx
jhIvOsWPyLaldyHU3in6CZOF6avrRjyu4/Za3JwomK5GPqCvzMQfY/sOZ/fh1wQZ
alOkf51swzeA9oBzvs06GkWXqzp+8P/3v1fYW07xAWm5qWV0YNARtyij5eKnIqGh
pRBA6NxW8mET1kGedlwcYfdafPaWRyG28QDQROuiTCkbikvtZJbCtMzFFDfZJRmZ
XCLbtvYeWWjCOOmbY67Gi3QabZf8AtJNab/4FBb+UHieMeQ8pCCAu6xhCDbiYGKS
Zi8lKlS/xn172wmnraZyCB4ca9HtV74e9PUvaWkBRloTH62MxJjUNSTIzAmLIYsu
v8weFnLSOOs54AUrQaBkt5JmfTcYMmU8/zVUQyCT88GEbPgTD0AgB5WvOwyuC+yY
rOpm6E4zDgPgdRu0wz5dx9j34w4hmVRMWDKDpTW/vb5QrJWultL2w+BliIFBgBur
OEK38xCHu8dqIZIZVQQ1goLrKjJ9kNt09UydXfYq+ZmHdyvB/pi/9Ybj9fhDn8Tj
e2mPPhd9STuDnvcU20YcYEknW6EHJTV9KewbC8IH9z0TL1FmF+rtwgCer5ZXGI83
KUzob6njvwOHHs8rcf56y6rckyJ+TOUfywbdRHEJgQEEZuEzZu7k1ZAq7h0rYgo8
+KdLFE+VCKRuFTEnIMHthwAfWocDl8kdK9POlQNQORGCUn5pRddY/i3lAwwgKDz9
7I9BEJ9OWKe9r69vH+fkJQRreUwxS5NPiaTG0CN1qBVlqTtUBPufKuMJkN3Os/Bk
FIyLal/kYWJZAW7S5TCzMhv5/s8ol0XIxwEPzEPdp6bqVbv/3XcPi5zkk15R2hpJ
f+c0znOj+DzoOGdr8ewPvfjWlFbDHjpJ9l+za/vKoKWKl3Llx1L2r45QXx1An1Fs
5VPZGhSpjC8JXLDF8MT9A7BQB0ub1zuJgfz5bHYpKMSc0D335tGlqXpv6D5a41kR
Q1vhde0eoJ95zXIzuHsm/ufvEB9FLrEeabSPuhSUQd6SnuT363YE9SL1xgPcKm2j
qf1TtsUcW1mmJ/2dmBaA2peIiYNLysjdFd39rpystI/4vhXNxPZzOlkJCxjxa6k8
PtTWdbFLn1PSX3z/WjnKP0Q1kO7tOBDMq3NWDOVELSJh+ew5V8+Aq8Fv6ByUcSGi
oGD5YakUw4eccRklAzDGoXESEk9q3FD5e16oXz1G7co7OtGEq4q7hf9xmlmXXYcH
K4zjpgNuh8KTIsP+lMTpEh88TE31KzEdit1BjMFh0ufsrhmntG8SfnAcnKIEYCpg
yAy9Pji1Xa+F+4a7h8LxNbctwUj0kU4tJqwzMa6N/bBuXRtUXEHqwmtmg+zFnFU1
itUFc97Pv2FDMmNKvB4nI+kvGJE4IbbTi6zahJ8ABWVlI0eeuxzjpy7vOMZhmg8x
s18I0WpigHXpsVALQDHevd7j+52plPNJtb4GOihWW93OvgNB6mnQ1bG8VUWGy8AW
XEeCR6Hu7nyyaI2hAPinBS7am7WzIOZzgKvxQRL/z//bw8+hu3k+UI7EMBVez+LZ
dK6MKUk4CnjBkcdfM9SYsbu84JZaceN9cf6XWFkiB7GEXM6msbtTDOfAjT92WZlO
dVX+H2O1SG6TwLSbEWjBHjtTBR1Pk1MQD0s5aQZhvP8YGt1JpIOK90E8wfhtRsUL
GEAPBCT7o+8YSEqKu8K67hZPQNv06xmIyykZfvIFySy3t9v+cUm8AMvwJAQiGX3W
ynfQGO/J7ecq4e9RVB+rDo3UG26RbWsAI7Fi7N8uNh1miqEhmlogA6TPqd4rY565
kFrM9KDiIaFA0WAkw9N/AakeDzFZyBrYiIEdU3fZKdk441c/1jUZvmLF0l8R2Izs
d2PG8ipG46FLC+x3hjoxbJVY+RR/JUdEfdOm5fMoZBg253vjt4sU0VIfkjnrRLSa
nZE8Ga1GZeQUY3EFV87bZnG39tqXtq3rl/0GPEj/jpw4qsecvkHtDrxrtYas5YgT
wFZbXLVvyKSa2Oy5b+IzC0dqUTllJ26H4yvXgGiXxbmGhmXj1sGi5kaze7qRrqio
nV5eWzkWNerJhY+zFK/+FvFYQXV8yal03mWEj1KGMQP/XKbx/VjrVNACKbQq35R8
299MTidD0vZmGPqKVgszES7124YKdDwuM5ax6EO/7+XzlqrF2TdLpORcn5xzJ7+f
k49q5tHV2gI4Jxrw1FFUZjBae/5zXyZ/dwTfvu1gxAVF2CHN74OFQ4v4OIJadkgO
tEmCxJ0vozH0nGWOAV8RlyrOZ2FcoOA6JTYTH69oGijSI1NPavi5jERHgtE/QwO6
jFzPcbgot9q4yL6ZihtDOfswPhcYPZHazZfvy7CyOO81rN1Dv9LbY9LRYmITkC2N
syZ5wbkkd0jH0tegEevN3E4JkoyLJpIZbuIzEfATRJWu0Quo9yJTIj4YBQbcV9nE
8ctAoX25L0HBx3Xkxs3RUPnonmBxnxFoczGInbz9geuLzmCFdIn3YhV5IUM34ILR
JcNWxBXV56GRNJW12RI8tP5Z12ziSnoM5GC3JvR0IeYnAfXR8f5enH3YGil7sR9x
WpEgqA8SNBbElIdYIaq6rRy/7wg/Ql6htWVaye+uvz7NmRDZn/wpKNlQVETkMyX1
xB8RQ7F8g19sN1jntJZqDGnZWELT7xOZ2FbkB7IWKPBzN5WkTPM1J08f+BsV8HKN
kizr6Q1gm5URLKhFN8cEBail03DP1TcXhsB/hMCLm7ckYckX9SG8UxFeKpfyhg2o
XUYw88xCXPwtpaJd2nl7lP/yDCCc00MXsLOJTngUmMkiMExPDfKy+bj4VNmVNTdH
r6Ozy2jdT0Kjv02RFGE0+SegGjuWNe28BIYP8P1537j+zVEFxOMDKk3xaDeAm2ia
wa+6mVvqyR5m2AWe6hPWGrvqqWNuZiErSIz8W100HO1rISjjazxLz3QLQJzHVxL1
RjElxfUIYILp8P18poW/bGcPZj7/QlCUg6o26XkfVXwbawIB1RfjgwsKZ+In54wu
yiQA5Y5vDZlyPr1uezBnHoYsD+SC+QvZX2OBDdkuuGea6xsQteP+y4PrkQ95aulJ
20LFr2WRm7J+gpsA/sjvMUQ+ssE41uTa7kx3OihcpSokonpuIvjoevokPr40KuGr
8VUXU5l719HIKgeugLliZhCp7hrZHv371P082F0wgys3y9JRL3vpC6tTrxk/rJG7
XYNSbjxa9AXTmgGP65uvG8wlhg265cBSTzkrVzWlbp/INar1XoDDkTQvVMz5v0x+
XnDM5iiWok3/1h5W/udqBPLEM4uPIs62gkOc3Jv7fG/3Wpy7OvhvLskUhvlblUX/
Bv55HzJLlOGj0N1eJj/trU+rxqlDzurx78SY6+FQ4SSzvEap17Qv4bH1fatIEShy
ZT7479TFXLEB3XoakgoFuo3dbi8xFRvZTKkQDIPwNtzvU0mkREuusci9C7OMh6UH
kUS5HLA7FBKFKk8zmdIhP+mAv6XeYxGchr8Z6L9d4fLg8nmwtVO+BhGOTRnXldyR
dSR8BTL64PnGpJOmWsCjuq/hsuC5PKzL0Ih5Z7PF9Lqf8A2cdcpSdxfEvZS/Bzjc
SlnI3b5lrvYDSjZoAtzMPXlzAo5m9/+90XW6S8lcro2uuW4yGUlpwnG8lIF1x/aU
1Qsw9MiLvZGSLjYMyhcYflncOZBpcuSDCY5aDUlZcX+NR8Og/QPMCS3yGSMy9FbJ
nWPqMZDKN4LRfY8AgycNcbAwTE+Egun1wPS0M7k+xqLj/84LNG5T0e+HNKXhNk9L
OtjvHoq3GS65psL6sERJNXLyAimnwsk6vWFKeIt3r9nHB4PepdH2tRmeXzd4AyV6
UG0eD9e8cnMLGgaDnm3Ve1tMP5JFyhC3b8ZV7VfItKgQAcPYVRxPItzXy9iWD0Mg
m4HilxP2NR6F4ZmhuDfSfNS3an4iiX6k9dR84qC5f13Q/4/m7TY5tha/zTTDuRzx
uP08he8md71EcBrA6fAHYR5q6QeZolKY9wnwOO4jKi9CjIz7RV6rUc8v5otxVIoe
l1kLd75h8Slrlfpqi56bZ2dtwCM94NKcJk7A7dtcflLhtMfUBzz1+22t70lpys+o
1oZjL/fk3mvScqjUD4nnhvJ8mRJzEQxXVQ0JYsamjGpdIcAlxLPjCO0oPzpCuI6G
zH8lizOIxTDga7isyfHMuhqbPE6A31NZ5jOwWXUw/Tq3l4FAbHv25IcWxhkFIm0t
XlTEWpCK7KRJDZ1hXEnedZnr+iNuOJofe1mKsstAwHWyTNxlX20XHKdaoPO00snB
rCk1chYo/g1M2IZg2fOGS1NFEM4VEbYwrMHeJp9vbxogKHjMsrNWD8r4x5VOhxsr
CNw85do//At3gKaxbJ2dSEsDgo5y49f8Qqp5wM0S2zoPbXGIbN6Elr4e6Q+AKq1f
8EOMM+r4jQFwwjS716YitoXwqHYjiImi2elSqur2JmKpuoc+rpz9pfLeXxZC8nvS
KYY3akJdNSBhgsPLpS0qlyRKUGWNVb9pRuM8H0joYNXcgUlWfpSewaGqrZD0l0uO
GSZbZeMR/4b4cH/FgyoY1UGX4iFxMNBTRbUqyifkMvA+MokGIHP1EVILXn0adXWP
GZzB7npUAosnMj8MDyWTsWOtT9eVMPS+YEJAcBZeN4I9r1zGLym0xQBTLRfs3toQ
EDutcsOmDBzjfAqo1Q7soonNu/OSqzTPyq5GWJhikK/XXPvgdP6MVG+IJlgpcVne
Sx97D/p3U+40w4RJWAFwqiuSR5P2JkV63X+wwwUZ/Qt8nCjB3TWR034Mw5KQafeH
WwMaYDybgXb83UFRLJBV4Mn2FQeBurdYqea+FmanNxMEx6Cmlgfk5u4Jw9zkfTu/
QZFKJrEXx49qpnGRki3Du8RDZxPSuMN+pAqlQXIylqjRidCn0NqSOtrPCyk6vmWU
kJsi0IqrqlhzhV2xNvGoGWIN1kPbowFw2FZCOCKuL/zeI/i72BV4mPG4bqeYyyH8
xLxgpudSID5gLwJtvnZaw2mpHiZUMq5eWn4GkwLMw3L9cbeyX8xoYmmLOa9gmybx
/xwE6NerWmaf+HxIck7XjTzkizZvKCvpzzR/KDgYkzP+3vMBznkXQDQX/Y3nsqZE
vmy4yFg+Wns0hLVRAGBkdiRZYBW/AsFMXxLdbtX0w+j+Kgtb1m9EA3b4tVY0dHwR
KwO/jbEFJB271UgqxrNerN0CftYsmWRFEuK2g9vhGCJPoWFZzq3NGQHRapMF9btR
r9pODkhP4wpIBbQdNywjGeuDYBlyYuN8EaOqOnRgFD/kTDH/vRGkWLBj2XAJ07oK
/3V73EUEJ178sf9+RSsSbOAXBKRGMdIVaq+5BKKyPmUgeHQ7QnZJd/WTva4r01lt
ZSDWBHolFm8+Jqmkjlzzkeg688FI0nRYsW89DdNX7+RXj/vp0PdOmI9jkFq4PcBv
RABC/uhSuXWUSkSrhO0NesIsBYs469DYylPWtPH7zxxRuAQB66Bb6PyqdvJHbUdi
IpsZoR13i1x3SkwVqRwUPmfJVOObNCqs6RmA0BUmb1+L3oLsrdpdnrlffIVbK1NR
R/L3wMKZkAgh8H4738I1SleN0z/n7PS0blEYXdL8EDDlWMC6chxb6aKgzEpEo7cl
MyTaihIyCMfcNMiz/U3QVx8xLiE5xf0ssLwaFl+VznCVQix0KRHmvRPkIXGrWt6e
ZLdsTQJqM5OGWGSj8QFbWg61xt00E8irsbeRYhMwa3PgBznxOrBJBcbgvM0rPXdJ
enhAVCYpovPDEF6/0kKwgesgw7iMxJNuo0vJ0PzUfUfVJ540GG+tmzteayutrkxg
4Zh7JbnaFRjKDlnw9OgE5mj+V73Gcu0FLqk03NuteWbRVb3WNq2jZ7Ake9/7WAB8
uYd4gqgvU8xHsi+lvpIgHAOlCNogcRopanrGguGGpWbH4ECHqxbJUhAZVypoVkPt
7PelUs27yuBQ/c7njzo//UK9JZqOgFLk8OcksNohh+AVC7BGkZIAT894qIscql35
3wJZWg2Q2QY3+kBI9jnsPS7eg/+4AQiAxZ8i77qCNYql+dLtMMYr/HEZOTbmge2Q
1btCmcqLTp6ND5DkK4G4UZLxt1sJJ/2A3g6FQilL9BQCn1n+sl7S+AcbRoU973iY
AoYs7WS50y4Lc9vpLB5XLfxT+m+RQr4g1nK3gAdD2NkU2blBn45vjJBN6+qRdH4j
603g7kfzAJnqZeAeVe+Y5GsXDsTG7s2vMLnqWIUMsbN4ajMb4Kp4LUxZNl/jmK69
9w+A+QQ+eZhqhZz/QfwaP3RLK+uGKCwOcMQfWYPpEhI1vTDaDuA8iU0U99ATnlbo
Z69NgwDH57uzjjEgI7551DjiesBnIN28Zu1E4tp4o/AKLECI/SiE2x88wUc+aKrH
+NjwAh++02fLzc+Ie+moeRCfaudJ8auEKYJ2fF32K/FFGtBro+2R1cnkvCY7vpF/
SrsfkWP+rFta+MakkFqoRt0ZnbQS+ianldA2ZmsjAgcwgRdWuEI3JT5ILUwxt+aD
XK5h2iMX6HimDF+VO74yITagsec43cSUdRBS51q0gPwh/oa5TzaTbO6ZAyZtGNmV
Ud7EfLRIB0/fdV5ZkAspkt70xYJImE+5GyqB1nCd3GmdpcyjlTzEPC+rXbG8+SNc
ICMRWBC2xnjjEsL+UIOmPG3GNXX2HXOcs/3SBhpK23gVreL4vzhgy6nagoKzFh8B
KxTL9mqElzqwg7G/E/kR3C+aj64L4E6wwVRti0SNR52NVdqGM2lQxAVjg616F4OF
aN0w6yjz+YNFxc9aW+t5+N1sk8o66MT4uCjL896a2+LdT7iGDqAAfTQ78nhlfiKU
NjXeU5qkM1IG18ZGWdhP1DQjsHtjuR2gov9DjGCtshvdkAYmGS/x67SdWIYfbEX8
yow90FkH6tLE5RwJQaykJYXvHHz8cJKkuir//TOnsRMYjwMSSYJJj9z5rZqWVKkU
Z2hCxH9guNAZzuk4V42lTpOMIM3iNhFsIczgbnBI7ldlKmd342A61KMNZszbrX6U
YOzhYV9+2d0/Kiny0i7O1g6zg4jB4zgXn4UxuTC73ZuwjWUu1glszDa0APe0S64X
luyLlwDyu9JSno8OVRftaf39EdybALZTYZsgygdPOumJRSsq9+B36DNdgbmucPlY
Uj6UkiDwaOw9WOBsfJhGKyL1UJmjRqcJRipWZOqaxciW+Ykw7BbVWxyEukVdycsR
/wngqCv9KirhEIM8wF/VVsAxtDt5DxoOeWkt+SZuS989kbbz+PAWTngsMpnJ2TY/
X0xIcOu05DVKSUD8h6wkK2EB72JmCpFIH0bDygC+BU60bduhzj6ciXK1wrf2cKfB
PjmprcK02sA6ZQHndjuIfeezZbnMHB0i4vM4qaWsclK/Lkf0QplraPMaE/M0qJwg
TE+dr+mfvpX9/QBtN9ZNgQD1SAlNppccOKI9zV5VejKDZ0WKSVoQ9+P4SSUtrFfv
iu/uzeB/y1E7WJAieEAcoaeHejVWFjfjVB7LZTqOKJCvUHdglLUJLaeS8vEBluIr
sbC2u4ANlSH/FwFOoT0J1HEA64UxjCcxHvmxaEVbje+GGhm/mI9LJnWjJtrXnY4M
oJcQOmJSUY32gG2u9KvI79Fq5Kojjikl5/lAn5E5nMLf4MFK/BGHZAA8vdOA+/lP
LwvCzpAo7M0Bl8U7Pl4cqbVtVUq7/Fa+bOGAyI9VETuqWcz73NJkIG44U9GhSit6
UX9KtMHx1/lvWotaIzrgeEgYSkoI8xMWg8rAzfhx36d+gZpV0TQg1Rp1btOmY5dL
0qJ5OUDor/Vd3O0zC1Csn7C/rNl0CUjLD0hwK5otLlle/CdKs3j6oowZHAnNAOr0
4kbxDCFixw3p0yb4UA9EuMBtZU4xHN1SGL5ainG/d+KSkTjTEVkT7oi4U/9XuHhM
8bLzn1Zg4YlkQn/THbXP7sHauuJ/CBfurT7gGiKyyxpihf8C+C5I5q2qugUIMkOj
ldUFWZiAx17bN42bneQeFTUNJ1D/AylUOr0fTN6PBis02PIBvxGsdj4EyWQJj+dl
/Ebj1SRuZE8OfJ6AAqOnUiup/OvNBY98IDm9F/KFmPeTX8mg3shQO/063kjMDagL
H0fDAw3Z+Q1Od/0yvE3f/Q/NqzmdBjhk2pfBaC1HGzQAOfBVzeBVPzsbVIf5E1a3
uKKe/9XYaXKHIWdLVrp+zN8woYiODAcKGN1eMnoVCh0DTLuJzIeQ80QLYVhkakzw
1ukyz2NztEy9NCr+FakhnV2j4/TnG1vh2laJLIzVilwyhgQNNOfcV7VStqbKo7W9
P+mGQRLVJoskOnxn57gBTXQWMm8yU4VPHPjSecorTD+OzmPEDtJEvMuhOkf3XNLU
cUk84qiV2u3Dpa0je62vpRT5uVFaT+eknJgqVjak6oSXgFVqWG99LOAaO6Io9aF7
c5Lrn+vhtCLNmA9IK9nqYBTLoEfTSUdPDKUSNZnkn5JFL5mv5eq4yYOQEr1+7RFS
U0OwFqrK9q/s6VBalxLha8p79qIMF6A3zP15bmukapiYPctKSdhla9+WsPfXjEU7
cg6MmO4/u+AmrAP0ZbZGbA1qb93Ll5hclviRKoI0IUsHrzGdBtgfILYID8gUwf/U
DUnKjViMt8M2cOyt0diMFM4H9bAlRGylYouB2NE+x5ahIKl7okYp+HmkOfx1pxEF
KjdHoM/sNmQTPQlLB+QHvTurHs3CrCUD7olCjtTYYJNE8uMMzJTu73wB0YDn4Xod
QNLO364fEdp3Z3sg1zkNfd0Poz+hKg2rXbZo09COg6gajTPkv/MFoHtcGQGMM2i8
RDoHNNG7x0DlB0K+kP6lBiXzLiLid6ky0r6vtAHHLpeUlAbLaKNW4ywSa4Px+Sdx
v4178oFUkSmrN8/xcfxjjzTDL7TLV0m6ytNBP7BjjXFYzpQVhdYDo13vJm9/MG+C
im2t97eycpU7XWf5w229yS9E2w8Qjy7uS6gnoShItOXXPlMcTxvkLlyztgdSIAw1
zbGKhbCMhrG/k7gvSyAzkiJzCOwyaCNKnYkzMHtOvJKJUw1GoYVPEUY+/RiQJAfm
tnRpE4kGPWNfMrZ9eXz0dRxRYK0hgxn1Q56YNQm5KdjP4z0Ecev6VZ9Z+DuI8Xr8
MlTQy4PEfkrBbyld6kr+EMRmGbXAq5do8Q4EsGPVHSSEJtB8FjBDUPl8nh3JHV87
0qEoxgJhEz30m++hvIyyTEkjw7NcjtVydgncmS/dsTpeOgyOuSPiundN53pLNEFA
wMZA0whe9EcNVw5RtJ+S/razXExWKI+Dt/+k/KkBLaHepW6F95GlI3+g/TmM+C4d
Emp2VpB2+sYi898KSiB66MdxkNz9gnYrRhoyk9cCUWGhRrPzNi24PW992F0ch3ks
iaDdkkA8to0CDNCH5/lQISqZk3SMpHSrpV2MbvBWQzjK1eS1DJ9tpWubM/cc1ik3
4OIdW/kyKx+7Z/SK1u2kKJz5JD6bNpDJ3mIZf8IiHFLMdmpOcKzr7WPWmj5umEF5
IrKAC4NT+s5LOFc4AYH/nWQ8M7FSeVOycFCsrx2iJKQeUASXPQ+Q6pYhG3WVUTjr
NkNWM40l3+IFid7kdFWm3v0ByczaHvuCPHwV3zrQscB6wOGEOZE/8UEXvyTY3DrX
rSmK6hoMbOoSfhPdmXkBirgHlw2Ls7qRMgef6XwX/YOUUPQAvuce6J8L9ZX00fIe
x1UzdkyXe34S8/lBCBg3xjGCnBmYrIGjR/94DyrYwKhZZX1qBLCWAZftVDBoqvrW
sKTphmNrNFaZwKheJJolk8CTjm+nXR9vKuUPruMWndo37D26oKeF7ALyw9n3NVvC
jKJpisBXm9vEGsJpfJuQGwXQ3KWQ2rmDjTRyehz22Yti3NT8lsUg9FYkuOjqu3ME
9qi47IXFMLR1CNOERreTWU6pP9RmhhAVP7tHogZX7AVAHwPslZVn7U+O4yIeK2wp
pRKQzHPa4OTuDhjHSUinHGUKkSul+DNfRexSTZvS/pL9JlEwo99trU9yoq7TbmqS
SrvkNwhEg03gcz1HmFsz6u58ZEHMIKhhAorSKILuNSd40884PgVIZxKjoUu5uUyY
4i3JZ3tct20hv5U4A2i/oJe+g/K7zHvfWZ4At9Er1/NOOkDgnUQ1tbsg0R/PU4Yo
4LMj6YtDpsXmvmOKXWX7I0n5WZbEObgpOufE+uWbaJDS48BQ0MYBSE5V5LVPb39s
jECvASdIccW7WOYbfmjJHLX3NvkLNNZZrYFRfh8ImFKlPFN+4oRAxQc83JGNZpD6
QoztwCk3VZTwnb+FUxIbjAkWcDhKtMG11NO3LOcoYyMkif1AnhHkxGf9uUvI25/0
DDgVDASabPi/rWnTmnr5EMkl55M0nc4BDBxgJvavlq8Fyz2MZ4k6uOue9rst5L3r
FMx/6aaccY3eSPwgKXInCbMJ63tGi+yQiXkqTOjjezmTHHKIRPtnPxFlOwlmBNiq
6Q1U/Dhhv4VhQunhlR5hrNuZM3dxorPEO0sEwsqWmOSsEyC7s96A8OKNlmm2LFXC
4d9uf8xjiIYbSqIEUCDloJhmbxYa8I2rIRBumAUkfEFYn/7KERBUNoCkQBcJqv99
HHF/tr35yUwe7MP0EuSPpYGpxqVDjLXrvoweGAOgu2DMoWTEdUCJvfYEKBetxjQH
4w6ilUJItT0uQO2EB6jGi0rUbDDWvN1beK7ywRhCWEyX3xiUHmS+qn6hS1HPAXxn
UCmwx2G4PG+EZBv+Gbt+E680sE5GGUXR9wcX5LTfdIBaAAdd6ag5h8DIlrHENUsG
WTFnhR/jBNrUJY+7nGFNqog6AJVYMWNz11AVb0m4d5g8jrrnYsu0cVEmxmrvjhP6
QaZEIWjF6Pt4uq0ZKtLxYAPX2SBpmIlFZw9j8ShU0MvF++9k1hFFqOyAgrbCZ2ex
njZGbJXVrlMh1N+scDq5yKSBtD90WQYNVJ/rwlGluKU7E+6tkTG+fGIczT9BNmLm
nN1S6SF08P+9efzwsxX28wj5bHG1jDmTefz0bpNemVH46Qw+1RCItdOH8En4PjKY
NlS065J+241ptk8GQ+RWIvhOMCdbGNnF4wbvuGexfwYnDRoxgvIFIKTfxHZunzIA
BaRq2PuJVDyPmhC8XJ8fcYmoYcE7iCaWJ96vm7aNOhhpe85OztkVSJD0A7wKNUfI
sem0qXf9cOMINXb/a88yYIhFCHUToGyY7LK2ue/wEaNJDX82wdvM8hkkZOpwLV3R
zlxB+Ukh2arkvPBQEPbuehYtWsBAGdonqVzHBbnS9Bmw+bRSreGydqc2ehyagRJg
5tDZF3+hlKZhGuXTYZE98RitOwMNo8/p4ImzygBYi8DDYDTzCL9XMmfVrA/ftmzd
ogtIwQsweN32BbV7AqpQDErTJCRzcGpyLTXHu/5gXdVVVf4J4FgAM52U9BcuN0Jd
6yNRVFuAZsooyuwGstEmwFwJFVqx7mQ/WcBCAPRMI7ghN6KKGFhcMHUEzmgvDd1i
3UrkuvTyutlCx/AAA4IRm6pxSBYDJbaN2wFSoXiKj51hTG13VpZdLQ540Pni5heR
HKfvt2LAkYcVmVSOBg3uGd42tl9PcrJAWmS/1itQ4mAdHnV9RR3KNh/BBfg5jB7J
alTciqwYOu1YXh2a6ctaaweRaz7hxydHPpAjI6QRQTlqDTZIfSluqrjs/4CPSh+Z
awWUjNH3m+HNgfdjhWwwnQ7RxhtJCRihTN5YuUoju1riBZ8reNeUzL7FbnJUmXAj
xqLN3f1SHhev6Ec4fviCeR9aLdo789v+L7pRVmcINH8RGpy3z8J8ECYxmF0bukpl
LyVlVVzgEO49/PIiBUcQwlsvz86vZovD9Iw0n6PLmnZMLIuNzrs68DzKfdj/3toI
MMSGnlCFUJinOtcyJXiN1F5yc4HLE3hfoBiMHCwvbTQqZIkcLdr8TGNReNpx/6Ne
wBA6KXtLCNhsFEoRgveHI3n5vnvsCW9VBGSYbMasXc3p/hQzwrKyqAugqzlnrgnE
rj3F5N8wytnZQxEWUXOfgGxz7P+VrRPEmk5amy/f45S3Osj35CR/PsatXaBq6Zjx
60gzY2Hjvp8yCfN/m3LsBTeykH++HMDRPneep/28RueXduDt6Yruk4YkzJQrI6+J
3mngpYrPnT3k6N5Koi14cVOcg+9YYRm94t5MQ2GwALjd/8er15VdUuCyE7mnvcqk
jHSoaHRSidxFzIXgWZYF+JygyaK2bVbrapVS2R/PZwICRLAWH2Xr1R1C1SmjsL7v
IXjDFZfD7KWuB9KzP1NCDZpaptwjsUK1cyUoCIsveD9HVJPZcPj771x++wHuw+gq
4Mu+D/ocfibU6F4k2HbWxcfAbK0TT+GxSLMTJXzOBY8apdKH/W128E8I2btJfZ1G
+dZTWnMqRUPpJBLRSTgW8xCIS3yBMm+WOlWHRc/LWvzggnRTvBU+3Cks499smndl
TT4TY3xoRLkb7ege7VBkd+bdZC66T3TbUqUal/+S0QJ2wdOLEoyIJttcZIcfgBuB
gJd2kKy8+s7R1dtZNNRibUFiROV0nu5ePBzbjunPsjxiGsEp26fPPAKBE/4YRLWP
sP+6bX23LiCrsJC8rbYwven76IaUdBpCQIQLkzsiVag/F1J3xKVAMNWjZaLKEIzs
LAHt5A+bXKleHRApM0HZTgTWWV37MaXyt1x44jX+xYn3bzDIBqO2qDoX4C4SQ6zF
je2BUb+qt0z07b0ESDqQnotzZKfTH47/zprItlOmBbrDWTyM2t9NL2xZgCyOM3Q6
T1HDJ9TOGYItaWkoSF+2S5cYxu4TwRDtbn0aXpkB/bciLIyCPzhtP8tGH79M7ULR
Yv/jCHidVxg5ia3vgIsMwCwy+xe13Kc2bpgkofQcxgjTjBn7PpA9C6wrA3F6i90J
MO4BDoSGmVWem4t0yQ4Yy/K116+ZBjDjycyYGu8hiZiJFT3SSmhZ+AQR5BFQf3f3
0mHuPI7mIct5dF9giBLk2pkQMYLuFYszIyy+DmCBk59RdxZuL+OM2YgCvIa5Sv7p
rTbgoDiielvflbyT2tE1a/hZvEOk1KTj7MLgzdXXb6QZYU4XImnpDTRh0jHfuSFk
OidF44/Ep1XucJQ77qYdXSS+jxLyJckMfb0HZA9jxmjAjPqcx1EYEqtsm17oUB9X
Zi5EDas+6QI9us+TxkOb4vkUM9OFMKf79N4FUUZZ6Pzfwschpm+y6o1EtZlHzGZU
qblmikoj0TENpPe13gVzi9omk32Wxw3N8WMqtReWz0fvJ77nWtXPUnyYqbTng/DX
dDkwuuX43VQgZ8aei+mYbyD20eD6HFHXXmAog1jJNe+CG/I+dZBsAmKLUjFY9e0a
YmGpBZ+vqNXQfmGnCDN3ktqtTgWmCb1NF4DSXWaoqp8/+4wvPAF9NonZpf98jTYg
DD/aGyj40jJzq9LJIMlj718xDT6M19l73UcHxRPDFrd7ttXq9ZLvIBo1/iiA/M/h
Zakle14LKDu897Uk6b0dp9lvi9WW5vikgwiRwWOk9ll/AW2H4SxP3m/dtIgIRAhw
WTUt7RMpw/Zh9bdiE93nnxrcdMZwZcGuwICRdNxrmanyjcVXQPN02v1vzew9+pwk
LoWLeeXUj/Dzc6cbD7jTuK4tUWCtrh4u6SiqTkvrWITspI7DLBTRud6XgVU2pm6h
rA3uol/wNrCZqZJB7SBOXdCEz1qbiLXaBR2yvW79Gk9wR6kAabSywHLqn+fdS2bS
eXKcfufKSU6s8Tre6qUY3ygGLiV4FHDhoYuluLSLEb8mO7Tg6HS3rKeRc4BLBerh
2bOA0ckLe390ob3MxqWmzY5XyUD03Fv+0ZPx62Ao0oEpkWKEhC1Shur3ASqTNKiX
/39WLHgJLAlS1obx0y8BhUTCAfu1qBt4+KENw96A9eNX0Czyibn8gWP77jDRbKs2
1xIWYuoMZWNKVWx7VN25yp/KCf7yblWVXKwfrHN4pGB99Apeil/poIJLmKr524YF
Os+2IN9bWkPrnuDnOHPAUDD0CKeY0XiTM8Dvr9Kfk86abt1TQlUpdKV5dOQ6FdAZ
0cZqsksuZYFAgFY/jadj2a9MsDQpVOUUGlji5T0Q8tbNWGkAuD+Tc0IGjpZT8Y33
X0MahfGb+3PLk/L6afqhurTq1jgqSHAYa52i/yovAt/w5ZHYqal6Ptw4XiI6Gymp
SQLXe3/U1Uwr8NZvCWOAo4FNbSZhRak0zviCAhrqQO2qMqI1TBo1TBonPzU2h/ne
FcgJETPHHG5r7P1eodeTUlBws9/SrReE3bfWUaPudFmro8VnrT9Q10PE21LeepOc
7Vr0x5JATGaEH0PFew27yq6QzLYnxMo7lJ9bumVB1yk1De1EtLC56biBvQ4TP679
IkuAFT9Bs1+RjAO8zM1O878ovtdXKOfy9wSmB4Ed9smjUmrjGbycJ6hYUScIylKa
fdOYLhrSShXyPMEyyJnowayFnp6xubHXWrCJoTPsouEiBUGcilUJryE8dKvsnkPk
ztdEceou/nvLYwlMOpkf4CK3MTbBHI5e9srJXm7oLPik+HmBd7YPaljvLc0X25gU
IWjW16VtY5zsnCH7qFO4Tx3+CR0H3UqsgnsVM86e+oNZ3qwfGfrF0ZMsnIyUkK7m
IAOjdpvlqf6+A8XnybhLKCYYFPCTkH/1Nap9Xf3PBIx/Dxqg+zHEfwQoJmfoMNJe
DzX7Uv+Ck1GhDBuqQSoonpaEBLIqPkXb73RbI2yzhWoNznEc8N0WCxetDuIRZjpW
FWwc2RA0H0deZzT++ylxHycpx1fUSi5TFLywitCX8Ux3agPDgavQNgJqKykoh04s
lghXY4xTOyPAiF6JJo17cBPBfkFkUdYsMZ/fjjYhAvUPqeKVoCLUy31//QXVsayc
lVIwwgRHvCPphjfdV/I49E9EbjJB78dzUyPTwGDQI5T5NXP8nrA/CYA2kxg3fWT5
VkEJHk/3x68JDogmpQDfs28Jk7nqc8RnAjtifoICPQVaMUxhDCR2/sanJbB+Qiy+
gPAQ07ExP/P5GyrOG92WLJgkIt9nrZfEwuTK1bMKpwZOroRMis/czVEndFOT52Dl
+w94jaVH4F6LW/298H6LNozoqnBUYa6yeRVyxfdaOMcx/nxyD7vOtkK8EyCCZpT8
1ivKUa5kK4MpKagoCrs9Fbrl9bdRquQ1lAAXxuqYF1eO9fV7t8icy5k5oehr8Lfl
4R2B32lZ9Ki+DNgYNttgJOapyEEiuH+DiEWBBhFRD0TTpYuwq2xRXhlkrKDMLd4v
bQtoZcJqr4CLj83jeh88l+OBchtPDfa/5e40FQ95HmFTnQcBBJufsnPP7DEQyy8x
+0/K3GgxTPZnvleFJtHzApgScvxGzOaiPTGOzRhVIsPmVOb9i41Oz1Q9VyAcsuP1
fJJcN0lsW72bXNoHxHXOBi5c9SYQJjZdLOUZci0vEL8e3nv1NeGBVy+5MZDJtelg
8GngVnw+60O2kgSv0z7Qk/OnveQqUiRnx56MbbAXIr/6+IzF+wXFsRJBGvKdUPaS
fAjQvEVRjXeHorqaUQzCKo7ap6SepyKnmThYL4dxjcJqC2nlywdUUyPkyANH0g4I
9sKHJIqAeVw2kS/HUci/HOLjma+0r0QTOMtGr5iuEqc8xU5adsv8vS10WgdKCsqX
zz8XmSf2Z8G+m3/6P4/PsjnZNxbZ/3DJ0VVLtJGeXTzbTRLMJSoT8zrWAURSS0h2
hcg/yWktznv3Fegt0AeYiq3aQQG2ozz0Ojf/+P1jGntPBathuDIFA/vnKpwgSwjo
5dnuJLZ0XgEMPLJk2m94AV8WEL73qT85uPnvSQiYIG0NcPNf1Izx02mkG0Fqhoev
O6Kg47eP8wMEn23Tic3shQFYciyCl1BanJob3FKWD5sk+feS/4yLodOUcovN/hgL
M3qgVcKYpyFgq4qsNT/Xz8XtYrmcCO4L3bnv/fNW32AepMe1qbJbvE48a1OWHRgH
qaIDYTihKEKkNUkONmVE54y4D+6Iton0V7FaH75IZwoABjjxXLi693kfNbw9Ocgt
MFo3e4tBYoEO7wVMtgVvquLYWlWrDQnKNbkFqItEWMi5m7gMNkapjaHzVDuNp+8h
aakKwPj+YvmXx1l6tde7T4Cm733FUDc7MMHKUTRbu6crB9Sc0mQClEnhryG7q7LP
UECLJVhlsBl/PR4t6rdue7dw4HqmDRnHc9k920oci+uPNiulfqX68NWoornW02I2
nYN7HbBC4qZ4JKvYxuAlfeJuJJooK1VdnP42c+Gu/pCJVb88u6MdF7LEs4I8e3JL
pcaUW21wvq4rZnUINxj7s5WJHWi/z203KDyPQBdR+WWr2reoKVqag65LldtkDKA3
ijGOYd4ErhdjapC4Fw6nOTcOibiQsjGDvfwDrz2YAz2hcelrVjbP5wmJ5L+kSkgl
t4F/vUG+CucpTHQxtlUUlizUqZOZamg7RhzZ9U9rOHAr3mOCJVFTyYi7x141DWVJ
Bn3xmukqNZPuDU4lm1gxn/NfyHczDeKlwicB8ww73rPNtgULQ5mUqsLUjnSzoYS5
GIcF9M7l/kLcq72TA7n2Kh2hxnbqgRCabXEKc/m9j/TDtVqjokqVI1wSf682ocNk
BJML9eDC0xuL6uSYYdV+2uIMePEfECTsbjReJcoC36/0Cyu/+04m72eTcqooIEns
27a7XZ3ImYTdJmooRU3WNkMQt9pdaClf8RF0VhDXuUVgmMxmHW0EwIc9ZZSHJu+y
aHS/nr7xtjpVnVaRoYvCiTtGknnSl1c1NZqr4mUqNnTSY10T+IG4HJWBpNC/EQ7/
36tUcgu3SBqkbKIvsGBRDyhiSqNXAEMnUGwdJOrUxNaeNuldF4nZsHvXlrnW63nJ
HhhCWcTywQZ9iH4aJCoWUrw1Qs+pkGhGWbAaNfASnhwH4UCoIbOqpS52B7o5PzVY
Aq2C7TApsqUK5JV3wrasI689moMIxa3F2CKndeUiBxISJImqxGR2pNuEjHBvGZUP
1J4OrFQd/hM9rM7uezTID+e2VA/ob7H2x/mWzpe/9eMoOI5UbGBnnailDh/hV/XV
sUF924QmVBXPtHmVpSI7dxNMetXWatvkWIZynjng78PfF8gj9aUkCr9NQenHmANF
qrJfLTDQFhQeJWfONv5IvST1II4bRWZWsvsMMZWtrACs6Aj10O99/2dV66Bqv4PZ
QDESr4EFuVXQbZKRR58JEklW/y1EPrCRsX6Z1HZWn0fr6Ee6f0sb9S236PDuqKsf
q7fzPRxwrW2kSfiB1B/Gemq6zP4iLNGm3nIN7Rdy2YNDES2yLG3nP+33JaAwSRY6
sy8a4NLlKsKD4q4ox3uG1c/SKMiQTjXLgrIVZS0T94dQV678vvsC7B2HCChU8BKW
RtSZ6rrxRbK/x3QBg6ZBu7Gi41oPfbqhsEwF/KDhT7SH90h1lwUNp5G0U4J4ZTGF
TAcOOnaVEH+dlggTmfY4HFxG28Erq0AOfXoD+8kHElopUMDTb7vA7450tH4TXBcl
pkqkIyeWdKERnVtG9R47P8nrCO7qwDRWFWWCZLjc/d9fyfAI8Iu+NWyPi6zeuRA8
NuexWkj9wDsrylKzqEkDCckPWA9FZPKaXGTFwJRBRAmOkLzHVwyq8g+nHhW7p6BI
PVHvILWlnusei6HFbSUWUAdRlWptbNehsCq9ycEgptVl2CHR1Gr3Sz73Fr9sB89G
kbukDYS8i2SYA3hwEDe7XcGXzgjsfDixpCs5VJgFgoaclIka4ijkRhU5Ax4cShlM
EQ24B8AoOKXA87AXOAfKvFihNvgjehHuiOhrKth6WfTYgMeFNy+qwvIFA/FbOepa
yEctD30aTW8skAWp32vDO0ksWJra0EZApKYykJofkpNqrkFtwkoZbeYu+bNDh+7P
SLk4aSxAqHWsFJE2qf0KHIO3ll4lWRts7MAm4PjQLQ2bZcHuNsVTKcawKlCXfxiV
ykO+e3eJjcyxIF19vGouhCyTI9HbwZSGvw2DGJRgtyzDFKmoplSlxkYlA7ISa6Pg
mRYdO9lc5dj6m+U4GhHpklrgAsDi4b3HTYAL68A9Q1g/2gVnrMar61RQEBLH8n4w
H81xN8wJFtlWGFNWp8o0wpgVzdZdy6YdWkrIe/q3IliDI3g0zBcBJ+eoix/qOC5m
SpuDUJ8gWz5+JIuIAGNVanbWqEPEQGECkC/2vSmZ8Xs22nIXrHkZljZEs8ZLAnUC
qLbiEsmci3D/kWKvBZZYG+w8DHu3QG7iHFqHw6RaagSVfnIIBq3FpDciaBb2rKDq
HAFKZzjyQTYGabCjR3YefXVFghnXAmr2uTgr6gkO5qVBsEfbx0SqiK2x7HVHRmO9
qwehVq2QHTJAwP8TPzkrQWECZPeD5QOGNxw7as5N1iiAplglSqQXPEhb/a9B4hgR
qDhV0/sn50uJPYhl3yBjBI0KfkDooijO/fXazkiWggArmQBFAnbZxAZy/Clmn2M9
eh6Uv2smwMm9M6iePWMW1fwluNWOiSyfEjstIi6TxgTPDoi2NFf5Ob+GYUo7t+1X
zI1v/4dgkZ//GIfoLbN8Be60NwAgDgmBy/M3z9483a/yP128ryt8Gqroj1exB/VQ
mzuq4SFewsK6JVCTDkNFOFE8/VIv+umw1Yj83VkJJ4phANhSpVtWcBZBUBHiOsKY
Xgny+8+wjz0dvr7AlZizEBXHVRj/+oDCMruf+hn9lpwwRgGWv2BlJ7XmSUdubytY
f/TKaoBPKe6SXb82TCFQ1oEvflgcqH5beFJQWAlKqAMJfJ6H+cREb2yitquGbmgv
WjmGn/JpmqIYXC5LUjdcPkAaPxxj3G7QlKrqHATWtClCEZsIKiGPW4Fuonz68dc6
Ap1ix65SqOGvBC8xDIqzes+5zD+mNTBviFO3GrR0l46fK8sLh3bNPhOg9ZpBclsS
MeiaEE/AMCs+QNTskf9WsYa2Qq0hKmLeqWVZ8SsKCdvYWCILV7Mv3EqvGnV1bPbP
55AF9EHMvoRprSpMFsQH+l4Y7WQG/OFH1cuZLkSrl0tW4coj+1zZi8rixQueCsJs
TtGQv8duPpZfQXz7q4h2DPT7yWjARonc/mejCDiAAIZ3yP0inis7/9I3DPCUhSki
F7PM2KBCJnVssP1CTR67LWoyY4DGGW9ceXrq5ys7flIpXvE9xGcdcGyN+yYqnbWc
4g3U9x2Xz9ZRzwqGUNGQEoncgIlYYjT+fjO9bb1BPyLZAsntdZKtp3lKsRuIt4aC
vJNbhB9SMUH2GX8ynNieQUxXjQff5S8fiSzrgFuT1z8r8FWkgFWNxwKfq53vTHEg
Bvt+L1MNCfvcjG5nRK1WLxlkr8vx6rGqAnvvpXKVUP4OL0OSPoViZazlC/mrwQxM
+cWpM+JkTUC4Em88pZ2u7kZ7JsF0dvs2npg6370hY+YQ8vtTwnWU40KT7W89N3M4
p64eaoSjABiORpo5Wg742DWTaVFdg1jDN021v556sSUxzqF8muf2wcA6b1VdyRgF
Qm8f1y9irwi8fHyb9wPJIgp36wgZlbgMSWiTvyVFEXJkG1Ih45nbri7/VCDBydCg
4jrVIOjaKQjWJe39cSXLoEarPxi1O2Xc5XcJIMKktoGMBUbmrs5lJCll6S3bNw5x
HIuGm9XbEZ19EikBWOickNChdD/B7g7rY/1irBL3Na2Tsc3HJkJfvVeiATB9/jcJ
tzYi2PqK0Cflb3oFePgSQ1OtqLwqIGT9nKwK+KKsG4/qM5m1v7bnQlAeYkfqFwjR
i11kmJ1l34r+BIh7aliVx0Mj1flOTj/RYkhQ3F5vZmuwxefANO9EJSKlUqIZGkfR
BtHKzNV3/VgcnLYvpoJgj3tvYFfHFNHoBt7xSflrlyao3enRzMNLr5FmLTh60WkS
KU3XTBFLXRnNxibpzsCGRpbiwOD5A+qX5XxAt/OwLP/b8+Nzd0uc0wiaFO1Z6THp
I96WjRbmvOHdVzSWJg/Z7hpbz45FS5WX1TaQIPQo4zglc7MLyDY5pd1sGGdz5uW3
aU5AUo+fqdfRCqZkjj7Wk1g2oj/V2VXqK26K7GfWDpRwpUbRL9xAcZbbk4z93W8c
eTjA/Qu0xxYPp2igkLNN7RYMPfzgC8VH1AttozSa1rD1iugNcGHDXmXyqkht7qbQ
jotZiT565y1gW6WFlq7kDxrQ1ocbsMMTG+Fq1s3EqvSrXcIwuUXqhmDlhOaelQBi
9aJ6hVSztLbRxZ19AJvF5PR1UUg8vuUBRU/auHo/VNPG0WM9LLi8Z1Kv4Yrwodod
vdpQRrrJUKB9IQhlwE3VeU1xRK3G0/JKU3Yvbt6AYVuHHES3/VlfQqqyL0cDCWSa
oVKTwggKTiCYQBw61Y7UIc9ceHmeSY72Ac1v3f0OWASyczl/EnKRUbmM9hnfDTz+
oeH7Ewkwy1dpf/Bu4Z91NJ+cyGJN5Nf8MWZUQuo2XetQdQJ7ZqXgFdDTVbJDrs9O
R5lHF+y0F+BwGmY2YN3jUCV5QVHgXzTS/M6gp0MgGQTryxEYq+gDmuZtR73o0naW
LEgt7V2nC6KWaNds9j8DvEmwhPPgvCaAqtM9/VWrvuMc4kCbtd2DRcIKeBto84E8
k9XHMTbdoOeN6O+rAO/ciK55pL/vbs3g4UedoVxF406ian/rK+w40n28y2BTEjFP
yfDgXLysA57kYOMD5ssR0KCfuB0E7mDD8A0Vj9O95tameK0aWj5C7UDHRr+s60Y2
742QG61rgXU/HexERuAqFo2T8L2fcKk7Y7it/f7XaSdycgk5FjWcxelwmVr8UASN
EI9Nw9CZUAtua0UbTXptbR9R6Ozg9VnF8GeFgh6EwqLxToSZS9yIBdvJqof2AbnL
I2igdSc+eY4Rm6Kvc365qSLDuKrV6QE+6S35+qL+9Kfl21rmrn5mY1vYi2+XO0Od
foDgWkjAsNWR2JlWHXl/Lff3OH0VQ+FAzDw8h70i34T08VbwPZIJQwFuSwwGcg44
dCHyPtVynJbqU44YMhWoMHHVSBkq1WbabcLDoWULYBMvvje8vEe1jlEfIpTchN6c
st/0bUPhLU9Ba2+/8IzAEhH/vJszh+Qd9refy7c34P724z/ODkEU2t5tPoNk3cG+
U4DH2grkyO9ebbnUqrh/U1wkgcACjKUWHu0DjQTESAq6G5AkU/3zZO6znNSrWVuT
+WKCuFjsn6xdOrnF5xFedRr7tFtJp11Y0tKq+IBPt2DQwd7bvC/2nOzb12ZJyxVs
1DEfGIr4bMo4vObpqWaQlnyOX2EMAxab2Nj7F3xPnuSyucK9dWVLsgf/ZAGkz2kZ
8h/TrN7SUnzIiBO8O0OlsqOJwT5m92Q7bQhlZ9q9Fd4hBGGPMDe16mf7fGSknXfQ
ggeq8O77/VdFYBcMIi0waeaAD9x01Ybbfhxzr78/g/YI5NMwU7ftW14sdaLMnHyv
8dtlxMlYDa032nuPSnYyVpP5V83aDvkIZ2jSEMIwMqxEVskipvB1VH16g2AJSWSC
UgaAH64OcxZbLUjQDcGW24WOeK+q0/2wPHm8139UcdGsZB3320/iURUxVWo1QlPo
eRo90LhBZKq8jd4xJr3ArwRz3Czn9mSMtWVKOp3+qH5zR7ZjetbfCUiG1fwMOebg
3493/YTJ16oUrrNc+rqZ7vNKhija2e4/4+yk2RGE2glv/QDdcVcwAjNDl1lIIqi6
tjeALUdQcZjfAwOryPm23snVnyzFd2wDtqHrRTXvxZ+JoBiQgeceh7debRQTi7nI
rRjVPf5NMR3euorBwmKjvqTHCdCCsdZpJcXcbC3iNKGfrK+e+Vkl7Qk66EXuvdw9
SjAK9Yc2z5IFf4hP5rDMNp1ynwwMlNx41Q38wA0NXu/IR1UyhkO8JGaJceKkiKdw
nV1fPZrScKzq86gIHoWj8vHYHJbxrVMKEjTDjgTQrPC3OlYMW/iyDiLHcSl/foY3
6zN+Pwf4UaZC+U9QrkiPBq7aAzp+IO70Gf6BHYlU3Q/dahyU2mWoiK08hzeb7foq
rPgWNBn+/TqEbW/Kh/EsQO5Feafo8hWC4Dqr0EVOqgwit5+s/ED6sOPHjmyGW3E1
QouhP3uW8L3VVFycCxuPiB9CLu/BcVD7BeTigB6kM+piYUdSGf9dYQUyVJRsHawc
ceSAiS+nEsAuSQD5NlZdl7wY4w4F3ClcyKlRNN8xe+57NaINmAgEU8wR063d6raL
IJ8IP1g8HlY1RGi4aCL64/qARAd7UjIXgBwzDHb57I33ORFC3G11dwRyZ+fkvSkF
7O9tDXljrhGdsvcZuv+a/g4LoQUudmwCoBuLbqrgs2Ur5zawVkiuKvp9rdtvjrRJ
t4y8Wj7p5l82WkxLyZ8fIoMT83T6wYvkSRqbQU2roo9Q3Zkr55D6+jlWLBD8ktQh
iRc0l7W1qCYqU09Wg5wG5swkMaURgq9ztdHN5oObfcEXsHhpfIhnffHeuFLZP48f
TtDWBV2tTzfBOgahU+WoHKUfiRHi34mYXAFxZ2sfe+KjCfL7YROPpFhaQ4rUQV08
wSr4W46GIEHUvqs++Gcuc8NYIZ5H9pTkZzKOXWxM18Pl9SD6WLU7s4I5HzKxW/C1
jy1lnbtclGKW3uIZ7haIA2Bx00MZurAcQ6SnDVZhUjFxS6+XkUP6fjt2tBAFjZU7
uojT4zmW9r2xo8d35fuTMhLg79VP38oRZkO2kYmaPYacznjJJTIGzCZUnzOtEpTq
NqyCNQD4SD35ImIrC5FmFF8NnB3pmrFNmPWHyCyoPzE1zlaCmcqukbVMZgpvI4uT
+Noi1WoOMe+DJ8eyBdF3zeJ6FDQFbyrVVx5t1HkVTCJ+/LrGpn1D+1UHSY5vem70
gBrsCuNUZlYhRt7qm9YaduE1qHmW4QaU/oCWk0d/xykiCOz8XRuVl5pkbnpUPbRc
9q5FfFWY6zEMg8cJ8cFR7XRv3SIVV8uwSGVMwsegGc+ZLoWBc/0E1DeOc8xyOrtm
hYygtzpLECjfaJoAAF2oeEN2KGhUHIXKCBHgR3ZFV8S76pDOLmindA/qs+n5HvSK
15ild6C6sRNF8WzOMjl52J6WnoK5Hz8fHt/wtZQcVgKlPH7hdYNOUkbH0V44uzE0
gYoW1HKosswCl8YeBluy20vwC6Oac6hUmyeHa2SqJE+0K5jM9bcdt/bc9IoQGat7
4eFzmIwmB7RKqxRxW3rHvwuhItT6wg0OudXvVSpo1I9I7qw8mx4jw4HnqLOj8jWm
HrEF91jLcG5jZFkTo9lwlPFa9XlLg3cHwvZQUpEjniJKPOTz8FcE+QywTV85jAn2
x0UZKnhVU9081/uLGeKkNarjXMbI9MNrxYK3HeIvb78KDI7RCAI30EsJQ+dLoAv2
tcOHM9EWjXpZWgYFIMnStf1nQgg6/B2B7rd6uM06FBRBeLkc6u/KALRpwZYzRh73
0U+fleJOD1XKmt84LqpTatZ2AWLbZkJ3ad65gzQ4ihInRH9WJe9IIBY6HXDOmQvS
MSFi6M6O8rk35AuhIMaee+4srcdIiJLVzsXQYQIcpUTsTBf1ZrAZShL6idIBcBdj
qspuT5aFtsIabzU2UKbxBbKC+17DRMFVJfHZmEBHsroo4GRVjF2mc0tpcaZ9xCpl
D7gcvJni/gyCo0TX37gyPr8tXA3zw1Z84b04tN4agapE6RBy7UTzpc9dOkYzh3J6
vSpQvDXIajW5VtNhq2pSoZmIh3b5jaEnmONLzBr71Hu1ZcF4eCDe6J2Xpel0Za+f
NgfrOnkHonZ9U/C5Wog2RjgQQCJuD4W+7reJxHmOcoJTe/ygLHB9VrA1VU8XEJBg
Q2oXEgvqZNdQ9BhLapnrCs69h+qPjPfqn2U63MtEoAyqjd2xTrTVa3k1Ife4xuPt
UqlgbmmuSqvwATrPwgqH2958OtTG30a/hmoZYpauMJTOaRBXQvEmPjpROa39UEFB
LukZJ6KPd3CalkP//7FwAy7jwuFzShTFmvTweWWiFsXmQCj6qX9N0uE0Zr2ugULa
PuBVqZEG0Kn5906EKKoLtmQ2cWyvxkBP/KfUU5rG+9TphN0lXOxa88PCqFMxwyCf
ZArQ3tZ6AL2VpkkyvX3Z9UuHw+qXl+HizOkRHbbeukiVDTLt1qAyCZCU5NilExzB
ugNR0gmu0Ew1744R1Q5DJDIxjJp724aidxcExL1D8U+jFzHHqTI8obEfSQgYLc6q
Nu0/N17/Lx1tZXo5mIoZkYeq0TpaDn5MvPy7Ghr1UWDtnc+jqghUfHDL8pigZF0t
+bNbGR8RA1X5XD0/+C+F+h3N6Hin6VCsKO8Nmhg98fX+PZH/xv5/w9z37lBKfC3R
ZMLkMBu6N9aiBXGLlj7N4xq6vq79KbLn6k9UrmmkMDTDUMsGdC/UDiaNeuExiqkK
OlDFCiFghCyl7RR8LoEAGNlWzG57XqfVY2e49CHJeo25Jf3p1T4dgj645oe31hnB
KWpiMCNXh0oSixypcpUA4CjbZasERZzI3v5iasT7wxa1vPk6zxFWMeHfLvsXIW4X
TPQpFQG0jTk1XChoLefkeaegyNXJbF1NHXJPvBW0RLvHd4XQCnXGzjEXLq82NBcV
jI1l3GCk6nryrEbKz9Gg7aOp68fh4avoYLl4yCwVU1YjUwavKsObz9MfoHwt7qiB
H2M0duOBg43YB3/rqws84useQkUFRPs2qTZ2xqF3sSG24lKvRFQueCdoK7cgTk/l
iYmP1FU0IZpaUSc8v8dU/LmGjEQ8VUV1vF39LRtZ/DcWhk7Jeob72d3BbxOtu+va
/8NA/9StybFRfmekhjXS5HV6/+LXsw68AF/ZtYSLPjmhECpXETfcqVa5NunXIpYp
NCR98FmxQjRT9GrirIQDaTlnXOwxj/Gk9+pGjwbsJLrMoobEEzXR22Jzz8DGIiOh
xbQiIBXVtfJp92KOyue4mjcp24fEHs5xRjYVvxxPWv0jNCyEoyD4rs+AEaoPC0Ty
iK76MJGHGUJ4fwMIlrhZSGk4d+sCd/QGenpu39A1T/WJEHcoRmoNO1tuXajiQgK3
+lrPTzwB4NEqrHfuSK7NOaByZeHgbDvl2UdcWVqwShvBMjlyD7eZD30IeOw3M5dp
vhGH6kF2VcdbbHfkM7RjyF26IrQbg21pDvXD7/ay3qyNZ9C4Q/y0yPB1x1r7cDAt
FQKFkv9gf1oEN+47k/lm4vRtgLxTIiQuc8OsVX7ra+j57SMDzjCqClvqdaFzuW/d
X/CqXb+aDad8MhiMKk0+ZfuGu/GITcZs1yG5srdBdBe+qrXUPX8kdH0RHQqzCtaW
JteOjuUHAEltvIh+WseXLDesV0OqHK3P8Bp5hrAPeDM5UNl60n8j4LwBCIlg0Fsk
z98LPRWij5twWYIpWV4K+0RRUV4fSicUNgDwU9oEnGXpyOvTIhiww12qYc3abHff
OSeZiGcsoscUmVI3yqlb0V37LJjZHP1RCqj4tSvxEVVV9isHqGrGVDjXdce8nNL5
4iVbGjIiTl0ZIipd+DoD7uVQ1PIj5u1PQAeKhLJKhION8SwTRolYh3t+Kbpb8lXG
PLn5B32LkKXmU18a7KTLSrn2i9z3DAf38AWUr6cklBG1s9jP2X2NdDGHDkVoBPQP
Ulo7XTS9OeESVowIGum5D0kbSG11ICDL2MlUYpxiWo1I+BtiMHyz3FQMaL2r6z6A
LmnLG6HijOr49etbNNdlWa3OP2EKqSvPLz9Re9VViEL8FxsbDZTex/FSjFKlh0GM
xnf284//w6MgmjU2o7B6iIzOxIwKLgv5dKsgWSOTD8B8Y8sLJKMxorOGPx8wPE/9
bsYn+jOXFuHkDzMPJyo6JS46j9UcTlxIMYirzk9Fhxn1EbU1rpyau2BzqdTLkxlp
XvMK+NEhmzX+EOpGju2w3/+mzI0tmvxlEqWHoZWV4oY3s4RmYQj7inbOD+6JDDRU
VkFJ7L5+VpPhmyY3QB7WqcbazUKx6hQnsWzvPJK4XQLBNZYqdOttjXg4akcvfrqy
KueAwPEaISQSmclEkteXtoPwrFuedVO7T0S9QwfeZIeRtLwPob9MkzAeu6j1XrVk
JyHNbL+tOUHGIE2YCPZU9Q1gJXwk9DTwB6hW3pUqzLnEAH1kWBiUIw+gR0YODoh7
KXjI2eAvpj/SIe6WQrRhA+en6KQBH6q698oCqgrhGy3TH5xPMRvCrmIXlckNTDx8
hFAMwCLIM+ruxyyXinUdyoBcubjLAh/SnZsvDGI3Y10Yzh6rohZvAvwQZ+TmxHGt
b4gOzo6AIK/tyFZZSj65Qx6IjsETT3ZL74SGC97eJKvq+xkRJemYOF0TqwKmI4ap
eRR0UtsXFTKC66lpZFp9z9P8qDAwnyKLIBCppm1oTGzr94NLT6Bg4yHVGX/FLyGr
Z5iOrBF4unPxX2cyInCfmQkGDuCGqeZUBf35NQ2JBzOmz4T93jbb3HIJyfz4JE90
IWGlWkY8SIlEaQKJzU0cmr7LeT33BjJIug12Q+1VQQY6TaLHsbH8HWC6JAPVFCGA
Emxrcfh8wMRyVwzE8GY+6sWRZc+p88TzezCP+fkosxRK9xDVoecgPRG2uy4mJ7ne
axRzazhk9YJL0LF+iRQ3w1i+PmBZrRNgFSw7klzabOc/pmt+7iU+b/kKo3ljubQm
J2NLPePjbtTqzhn1IIkXOpEIFYtlPNmmk6cHP9PFeEWwbTFWiZYRzc8QTWralv4/
MEiZw4HMLeS36iixdGvb2nsBfRR1bUP+zuGBUP7JelgfG+H80KO3NqO6Lhrhx+Jr
+aiGRa1BwnaN+RTy0F+HACR9oMv+ULX5YKJqQ/YfaFNB+7rnDI/+REEUHIZ72IHn
Axz80ofCm/LZ/A2uLsHewJBYc2fd5sxr/oSTQNJp15lMiYR/990QvOX0U9JFfc/a
FSBy9p4evqbGvhPcBMb8o5Mg2LKqzBiE3QU8UKA6kFuKFfxaOKsSuES8HprXFlWM
qPsYGzoenfxjTGfA30G8WAnUXVrVW/yUx+xoA0EkvGkM4xwNHBr8SgOVlpeLcggi
y1NRVCDN/fTBkh6a7z9saYg4IizG+kqk/JDQ+Yxr9E6CEwxO95OmHC4JCvXOaXFp
fSDq+LNKH3Xu218eTlmfvjB2RvaR+R+sJYKVnM+heYSP6QZwbnXINJpfDkysER+p
CLRM326WM/kX2geiuzebqrt6odIpTqmBsrO4Tijt4adHn7gLYcaDhwIh7S7K2yCR
EEd6f1XtSZ0nBQztIBwHl/xx5N47+x3UfCJqEZFtHOASDC9EPHXoYG9uqpa7i0Ov
V33NUuKy2Rc0Q6efWWIfYws9Qq9CMKDfuyUw4A7SRWDcunVi8MH3NQDD56Vir5yh
pa3jsi88+dqk51OMTtfo7q9R8MDdRXzYJjgI48GJlk5PvBoceKaUsJySZe17Nk2b
5s7HdZrXmlEM3i3aIXxavC2ujt1Lye3Cn6aYhG+vy88wqBIsix6ExU9QAkrqkWMn
rfPpmGqgeAqOEqHXZUewXv+EriBCkpo55/MZeBuG2yknNsiFgkdN7QwujJ1daohH
KcQBPD3QKGlHQAVekCOCw9c08/9XuqwNMREVebvmKpDNGex5sw4gHh8WzVGgKVlZ
2GfdXX4GM9RfuP1XzKmvdabFZMPP1bYMKv3RKlNhT4ym6ZH4WjD9AOC+Diw16t5Z
YVU5D6s7r/Q8Q0tZDnCn5HpdYNwjNa26mmG+FFDAGP53xamF8+CdH6NHbVRLQFMC
ZNrImWPH7qVyVGM9sfcg1o8ZZGxFk91caKiunM9GDCi6k/lGFO+nLOwjts/SZyiF
exSTEzq4bCxTFcv9lJfpYSQ/MfT4CFTeuTm3zVh7uTZ6gRkVjdSljYJK9GX8GhND
UE6ycIZ1v5NITGAr6s0DgwYJkFg7UCOFD5GHwtfrP+W0aw0wVRcXQLMpljSv/AZP
hmy3gVjxwHwb1Yw8JfoJ5cvOGljgJncRhXohaX4PKMR2s0mGCiwt0qGUeiQgHSP2
JYnMfXZ3RnKYDoSjKQxhuESNUpLOy3Uw6Tjlft1MPCSr2mEBA21vam7QQ2EB5Y+0
EnDckOpxyaj83m/k9VDflA27XmS1pX2+OxbhDmu5ANo0kkHB+uu2mHEck9l+t4yc
U5bjZFUhFe6X6OL+o1DBBvwFLT8hQAaNhlQnmYQg7b3tqo8ofT/hjl7t93eL6dsJ
fcaApV9NTSs9H6z9fnZjkxwWqRC3SD1ap3mQV7jjbprHK/hJByuWDzQQbkaNwH1S
XCOsqxUpLImDy2bqvd98b7dj9FQ5WE0GdLguEf03yaUOAqLXJcwoAQWvrKwT2N1b
o17nHCG2jUDS5RgYAfmnfaPrHD5OJICKM7yfK/3l5m2vYUIEyNt8RlRZRmbjX44h
hrEogWUirOGdutsfpTAbaQHRKYIbJbPy8BsecmqKViqS3Y7tu2108QwzROMZg28t
2hpafS/ELtL2UY/XnTfNBenU4vftHIPbtiBZDh+8o2VHCrD2bcJyRiJU1pPMEaTf
y/JL3YOoQE+bApUTLBa829PtIguBJtiR5ips8/O3LUxmJfDwvy0pwWMqKQwP+C2M
plmx1om07Y/4rLvHtM9PqpuOEKNkJFw86L0SIT80bcHY9EOFIPhc7AqXUteIzwyT
u0oo8DcQbZS6XZUd5YiW529o3FI6Vakp2fCVg0bks0tyMSRomgA1903MzojofITq
Kvn6DY/fFb2NjXOKKnsQSE8ycpUQ50mgFmX9zzoGX5hbiUxrwgOK4FEYE7yZOYns
5RIz+gC33qDNHYJdP7C41t6aN5t5XqQPjUkePsMlAumMy/zMb6Ok6FAUIwSSzr9E
z5ySzGZe070t5fUWF4vmseP0W9wd+OqroSrxub6BLr2R+DCJ3842af/nJIP+Oz40
K8qqZAs+RzTkD7uMGj82rITz4kJncrCnnPFPBWz4W9N9Hgsiuwr5YYzLORTs96iA
drYvcsZTYOEcXuInDqGpGUJ6ZQkFPQTo0BQgnTEt7/71pIWw41WJMvobK5QBU8fw
yP6PKWwMbTdxe67L1dXi6okqgBRama1a3hJ0Ch57E31gXGxUCwnsiYFwgO1vO0u2
NOtedWH/MFjPBD+QDfBBxIWmtfqVLcDoeACNCHX57vqg7d4zAXFf+IyGgS4/whtx
5OGxr6ieOmeZI1NGQDReS57iezeAL/6QYrSekmnMZ9496HCdf06k+OhWsHPnAg3x
qKKcnpEYThnCNBRIejVp0oMfhUhPQV5AWvwsE+00NMATviQIwRqlNjvtWkp+ZJe6
EOTIKIYLpxlJEVOLsZfqOvmZXAdYXJmKkyufsEWcS4uBvpZVo3JRxMSfZBLTXyL4
X6iWS42gHnbI95m3CAKGYoBb3NiKzJcXxKt2Y4lpSD0dzQ+Fb0neHxBEM/1jyWNg
XS3s2WuuEUWER+miV9FYjUoNJoY9EztCCrz/AvHJXFgpeGeEtU5L4hwlTyNbeh5u
7PIIi+sDj+nss6Iryh+3IVqMVaH0V9gIiO0kRY861RCCEAZrAtjp8BuF4TuEuxCB
ez9t4u+qODIajkIjAv5eopZMOWsebIZj0v1Y6e9ldXzgP+05h/wkeQSQU+wz+uUY
cRJyb3ccoEotAC+p5oesr37vrX3JUco3Yz9pFxEqq9TGab/O2dv1mk8aG5pJZrz4
4tsjB+m2s37mV8mHZp4terQhf2JVorwzOXt/DJlC7BCIEEsLTgqcu+4WLs84GrED
4NhHKqRkDxbBolAKSOHbdiL2yBoI6XxpIHaf7jxHJi6uTaszan4x4cnwUtPHMU9P
R/OeYUVW7Sy8320Xi9mhIly0yvwG3ibBsyMFPJQNIvlqn2m92VC3CH1zIVRGfTiJ
QlQfOFtLn2OxnO8W9i+ockB30y3Ap9JHWraUFLy+L/zh8KAH56x/yF5QJQAm2jT+
Z26oKrH3+Mkki19bs2t21MxhyiNziVRfDwgR9bBx3TJZLCMsVZg5kTfJNA9j3fPf
AK/armBeZ0ahT40/Hmcep3S3E5G7W0I0H92l0KKn+EZCzkY6nDAXnl/rmm4QNU+I
AjxA0aYwLO8S8nz9IU2KCwuAKldYgUPa4niAedYEEtodV4THNIUvXdysZ9EruNTu
SEt2VDMyxtW5PP1U6eZ1O1ZX5K5XWD6lVIf/cdpW+93DAuAZ06Rl9d5WRxp0DB1U
9VLAKjfJJoWRNeYheVVHJawk+0xZzYCv9csyWHJrAVE5/h99vFMonFa+VL+OLyyj
KrR0Uzxk+e9t4c3Gq6XcIek+MqCurvVBepHvdAT78mxhdvSZpxami6errie19QKG
6FtXRpH6gxGPDOfAlGiv1u85494Q+aTbmQwILve73y4IB9faKwDSgX14HbrcjWjQ
zCXS159MZP3EyD8uCCwI2Cm8CaUJ/LprRkd6HHqBA9u5Oh7tk44a97Uee990JRz3
e2KTDn08YZfjGcfJuBFznsLCcHFHQlQn3miDoEHFpX7AVJCnu3GB3Jh1FEcYLybO
q3tR4WNWroU6ljY4LrgdoMuZ87SUWTsrG2s4ZOa5WsNTZuf+9j58y4WbJoSdED8V
roCK/QmD/B0XLNkh0iYPO/BV2NKmtg4vytj7nk4YpTRwKOC4YCnxE7tw8ASGGQQL
imqe8tNLd1VZUbgIfP7YeNZ1WVuwgkhUIATOsPCRoxaOXsujryla4IzMJyHs+Yoq
g82pozW9/WzbpFPGfc4Edhivw3KMZQhJr/uXme201pxK0yWHhQ7pPEqJF29n8WdL
nN3J+cjw/3JS7QcAEcFulCh8dVIYNGYFMCvloacW7YSuLnZSPtoO9rA+kS0jhbEC
Xhqn2KzDiRVq0vFqxjG7mD4u8wtcULgjIpUJDYYs4GMSMlBDSLSV3rgGMYbyC+/s
6tSFNQw4siWVEpWClSprUkzq7D4SZSVWZBJ8D8HGbL5QcTSboyXw50eTDG0Pit+v
V9HhkT8uv2/uojPF8kfO2KSf/bBQpxeVXn3xTcv9uTGMJ8mffexsWY6ztDuYZieF
O31q3KqlWsS8VDKWe/VNBgp/5H/J9P7qTCnqaqx6ZMH0WN9cQNccIxhWZNXzxcT/
bf5PGPaDnvAUPI26Q43RpeldPEUM8LaldMUH0GO99ooUfUTCJxKdUvy8tKOv1BPZ
ulc1NxcjWJ2NoISlamd8bcEvierrm8XLisJf3D/V5l4+649H0oCpgPK7dSaAUJxf
pf5VF5n6Q3412xL0otlU5aEPGFVLh3VlweWq9hB70r7I9DqleNUpNXxiPt3Ke7YJ
Jk2riU/x04dhNON1SG0G03fGGO9iDbX2jAf28tkemkvHQlCKdE6xnk5LP/Zd8lTa
Qw33o4adbzX0ZOVH6ve3pa5ZG2iBxtjL+N/QKsuux7pykTTIeC14zOxHg8cH66NK
0OOGTIlZo/KU4Ompr+YJgXGJwfN8mM26vOOLxvaWesRw/qzl3V2/f5T1wj/pClJp
QMp7z2kHU6X0Y/wSINnTVj1bNMDkwN5inIDD8+8oFvbdJLoJHd0tPGIyI49WmV5L
+BRImEnvZ5gbsjvf8xgA5LgeNEQ/73Lq/0e9ws1DD11WfpDsBJG9kQ2DcT5QNj52
303tUa0Gw+v9dqvbWoTXTL/ZmlPg85YWBRozgio/dBssnoNiOzw9sOyHJD0/LcRO
25/pK7ESbvLWr2p+vuWiG7tN8T8jVamSIkypZ8IDIoVGNUJ0BnL40NE8KJsQuLOt
msHAyVQ02bbj3j9IjhJ+il6kALK4TRX373yFhcccbjH9Jvibw87i9j/k0v2caq59
kVXmveYU3hg2zacw8HRCqxJTr1iwMtoQvN2Tz+HqtgOWdTcNtfFAuJ+yluCvfUwk
FfM2JG53wL4W0BnTEP7xCHIUnGtvD0Cj4JoOsqiOykI/iCiVZ+t9hO7OosbC6J4k
RUp4/oID7YMGQw3H1buXtesb4/Tx+FZ8R1lNGbXHo8dgeaQ2lqO2S+wS3Sk9kf1x
jNx50YkJTUiF8s/iVPTs2Pp8ZreyLAasEiQ1jBzr/s87o81kD7XTuU7bKGIazv+G
JREWQtSm3JkJO+aDkcck40C8hq/IdtgQ0TC47sIhY4Fd4MdIVYD52NOBwt0+bRrT
AQgjH9izVrC06GrBD8vCH3zKFwger5pDIItzmecswGIEsa1LWJdGj0+UyypSsuqK
RRNaoYm/J/CUcDIBnjXL1PpXR8Uke+chdZ/jaf/TvUZzV555i9dVUq4i8UJiCfep
gmt3cEgz0FRxH4yKPiPDHH3tT9sg3GAkvbTK4vCCIH2wMO9VQKIzi9DXSqmoldis
w/CPno3uyq30rIY0DfvnM+A/PFG7kvHkIZFxxIEqf0+g4Bx7aIk0IHRwvk+P81xh
rSqm+nFnv2gd06n2zDxh3HChB6dPgVjzJHvimEt4ZZtfq8mXDYUH0JC0aARyfNGl
60FMuWxuPDhHK7keTUiSsRku+0OR2OGBlo458v2bU6aXQiwZEiyVg0ID7YvvrJ6D
Sg0+zzZcP5HdpHf8FD10MEonQ/O39ecr2FkbI9MZAwdxZOYrlkdLkAGrgBq0TgVo
3h/lykGcI/GbTQY55cO0i048s40ijSpRrLAMY9c0v7U2IAX9zz6Kq0MHBfEyfne2
NNryUEXYmoqw4VhREqTapmYzsDdRWJ/IF4GuenhYa6ZOSW+RZ55jyq25wFzZxTN6
K9iCLt2LbPKufRzHctvoDlWlubNgdYJDRRNDt39RS5HxGZ6erQxNfU5zDsVkIbSt
oTE6pqS4euDRS12jGDd8+0dhRCG3vxqrD5ie683UipiLesQ393fIdT/+85KOAE2l
gvV/4GmZIbnc4St6jDm190eDEOSKpR/bAOedL7gBkRMio5WDNgirucG8UCpNi3sH
wuam488nhwxGrcPjhW3AvOGdryNKOyAs6tA8qDatPueiD73MsQpMoWksOlWdZoFc
KZBM4sIUTcPAzzZ9RsQoNeQA6n1H8ttrnx12rHUpVZDhqxy5WQbUFjLEOSCN33xK
40EwakfFTC8XNJrjqeVjSlBOBslf0KvRTIZWb4WQlXNi1YYz88vf4RHg872C70+4
y20kOpplDy27MVYJUajfcZQhlTJE4lqQuGIf5EiHdb/Dznb6BpqllVsYI4BTE4UD
FW18E6ji//R/2VyzDv6yi8CdcPxq/K8nkcxjqsWnIyJXvsuyye3cwE3nj4qI/23Y
2lzRIJEcvVGzkKvSHyKrvkJAHAQTUAw8I20JvUaO70G8BJw1cTyJ3E9m4RlaUKo+
thEmILhPgHftCsba448AzSvsknluG/tDRbSXsd2zs6UeL8+ZbtBwS+scDGP5dfG6
WS3X5efisfR+ITIG7NGgGUzOVWSVoGYq3+M64Fz+zeUNwvqMTDXTqS0CWwcgwSqO
31x8R1Q1vCyZ6FgApejwdl+NLP5D/rEXu+CuKvw1aQMXLk8paGS8rC9jA6BS2uhu
LrHQVgm3+JkcIGJMKSfVa+EVhJSMB3JeX5X4RRDhnS1rIAeCVBaOKD3AaA34ENll
V+sWWo+hwzC/PtqXOzUxkNivtb8XHrOt2kFczjBUOBqLEJZYAATHJfga6b5nbuzc
NxVVd2CMPd+mqC/5ZEo5Q5lAjcyvoEezb4uYcot0MywCHqTgmhaUkCxbZlE7hiAe
KXQ8peB3jGZlhjso0ggmVbzVQXstU6hPKOamZ1KIKLz/e4ZmpgdmykAWPreFXJH4
m9PHD4eOj7zPvY5EsFRdBfBRyup4uGPe3Z/SZ0jj6WSLQqkSwQ8dvEohqMQfrBh8
u10m8qGFyEE2e69VxTyN6rYIGXdnIW0l3wpPH0Qj+VrBFzo7xy+awJPcS1ucbhlJ
xpRh9D7Qsd3tgxoCbeUrMS7rsx1rJgtn568d20iLmKIv8hrJG5jNLjdq25ZHsRL1
eJ5s3s8lXfsRQu9xAoIPqmo2Ohsc9CWA/K88Hgf/TbDVfhB9Wlwte7s25FWeVuLa
aXC9okXsW0FmKX30dYweSpEgs55RMBqNMePslicB8TQHKAYBW8bSSf6vjz0RC7ir
UlMgPSWpR8+2KIKRNQAkj2mAaG/8bY3ruVe5zXl34lLAHHVL5CZTFIw33HhFnG7W
09K8x8Mb2a3g53CaufCBiiFSkDd0Yuyt0Yq8bNnJS+yvuKTYuCth/dTzYJ407cs3
hPwTw6Hkv1AX/CV7u6gsbWBLB5u+tpJ6yMl2cQKZkgPtX/iGEuhDF8JgshzfjEdw
ZEFC7DQ3rCFWnD0J3chNVW/wTh4lwkamWPFjFQcPNCA9G2x/tB2urM3X6luwtHS+
jhiRmjKsuqoPyD1ybdHLe0xKFQRoq2UFHtJ0+la6HIEb+uFQFIh1oRw68idexkeg
EOnVTHiDJl4IDVQ2gy9xY+cUBKXGfFdcLlPYH7T+5vmlrqGVFtgX7lMfnehh0yee
7mejKR3yL2V32DT7Y1tPf0E51R9KBlCPS3iycidzE1fiosL5Jf+yCOELeADTmej/
And5z6V/I5vNza8oTSRN0xDIX+0Xs7Hd5HqUc/jdELFez29NQR+peL2GaRw9pg85
09yXqPJeTPc6LTUjRpnULWhbKP4ZaWth9faUSQSWn5Bb7ffdKoFiq/UhlGoYQstG
7z9TIny/vxi1EB4tIJDy+qjTTtyHTB6zoPYbtgkwegGRLIjRwIWDhIaoX0C41aBm
l9eTXSZaUaAigJaumDVPQAaGCVcWpEw2wD7jhjVeFboViScLIPWDeJoYSBTDyQme
uCcN4PK3jVnWqVS8rG4nsky7cagPA7WgMstTy32sik/1qcdK67vF6NJFuUvRfjzs
cPsDeiLHLXDt+15yZ2oeqVFYfMG9NvYMUfQIVopCNMaSssEFnxqkzSoyOqUPtuuH
fzLXqd3OfxGZERAyQqw7fcAUBX87nrpvDJGzWfRFkhoSFFA5WIpkX5vgI7WAYrFT
NtxkbPsF1CAvqvMz+AOLXMkb6RSgk94WvIN11E1dH5CXQ9/4Y3ctZfu7W7lR6kzR
CmsZKmH6nL0g88NPpqFLepwh9EaXUfk45q/rov90cbFkumX2xwdlbT3xJ2F15iY1
MnrOWAsTNrc7kKNlv6FKn4moZsu/jJkXvBS1Sipzc4M4Hl438V6vFEgNRwW3lkbj
omK9qUFkLz4qeKK5I7FS2Oz2ZNpEkewL78ployNxJZKLwMwUH4junLw4yAcYSl9M
txn4nK/wvltz/+46Z2nOHzu6LuVBugbdBJUhyiaNujLEOmKZy2oM1zuHMempAYXn
bvhkjlbuAaOu9pi+K09fbpqWLuM7Gg0Qe32dHZdU5APsebwjIp3j2vzWTEPZ+L+K
W/G0RjzHDqdsWtdQamcD2ThwCxD1lHlzamFNqOVNcN16aUXD1cJ5WMt8EQl4ooTH
TxCbvM3X6qsCa82CJXbmvjimknqfJNv7gTHYEwHZ/4uLxusRjjDCtkvQyTEegI0Y
MLiY13GSWFGrCwT9s00VCQfs0vQLYbas+s5inzcPGOFBiB8u4Ex/QZ8dXKSShg2K
j3V4PNbPeH+mu8V8s66mxg8Ix1gz2crHrZOTLAegV4v9OXqZR4dm/pgkNBW2U3D5
IIoWa6c5CrV6aI/Aui3YciMQZUq8fretyZUyPvN/1OZS01EV7UxsuRPIG+55UAQ7
fBULwgyeAxcZAjwp4lMfQJ/2KXcUELunKjcWPgmXoJz9gm1i8svWBC9a08aUNh8g
4kiwOAV2iPtPyx34qImKTREJ9E+Vyib9XAyaBOLsFrWbGRxGLxkYMZ0KvvVlhrdX
QCMGvG3GovIgVJ5OeGk5s8x7owJsbf63vauE8DXKY0jioVCw4lo69OeYLQlfmh6W
YaRVat05DUOiqXgIIcP0ap9jwqRf/Kkk6J4I9B/IK7D6KSos30e27GAZhh8VfwQp
5thOpCFA6mlCHdR/BKnbUFhBw/alo+/SHloh/DZB1J2XI5LRwCn2zEIw5xZ1OLVG
kUKTCUWcHkb4LwRRYqqyniTfpvy0N+2P/G6vb4ea1kFSWkS+mEC6RTUsxIHCxE53
/G3HJYirFRiGxzSyJ7esW8uRKZvBmjAhTIqO3yuE4vyfgG3iMQSmxDp3MTYOW7Vo
tZBvJwmUvmxp3KNhA92jC56y6KBHhoHsXwyiC90GBpSvGJ/KnKKrVKohBppUXu9N
/Ffn4B7z0Cdh8z8XiUMtXKjIw0Qjk2fGdA0f2ULw+4LfR77qAcUZpIROfMZIRbsc
Fu0wQGg5EqsV3ujbQJGxadG8FLCt1gM5UzpZmZDczNOUYgnc8K4dkbZsvvaBd6UL
loIKpIMvYrR9XrSMFWlZPcRXPkm3zYkNlw9/BD/bmQMGIzy8mMk5HSalLrgoSvwu
7Vt/Mk+oWo6y5t7YHWR8qotUYivtg9+gfR1CIXJmOip2YlsY3YoI+8Su7I6UcE6j
/H4+GR5BjG+JMR6knnzHGTJAG4Q3BTfTGuxrsz4xJ1eThHWysfMAFpjJa4kDp/u6
uXlTMztfhl+BebMivY5tFiY9tgsU+PL/uCpOtJwYJSO4K2h7gn1e5VMFeSA64CfQ
5msyfmoNI9VtYfdNue+bjWmXY/pTTaUTOBGo4IGM7OPnYKCUDorx00kxRyQK5HZO
Ju1/i0GPtgGtHm8AV6dgEvp5rxFAjBc0nZuT6ltYSeefFqTGNvFuQ6ezWTxqw1Yb
d1km0/SHyCzTxWfeHzTL8T4S297v7nrri1Naa7iTGtB7YoUut9HLratJwMWBerlT
t4UZPX1O1XcQVYm3aC6JdDWVdccy2YHYF2/8yGkJigmhNcIG3+a1wm+zAR8VywzD
Sx5Q9t/U91s666SUidAUBrAnuTMuygYgTKKGjFOV7++34fq8LZDcOuiEMlOuklkJ
K/xzTuidh9+s+ybgmmQpBzUdHuUm0h6AFtuOREVsdjJJJ6MtZrqJ5XboBft+q6vu
Dq633F3LQo4JdZC07UT1ZJLGpNAMYBwNi83C/dFYcUjDiOunBlF6VjyulXhayVDc
QSYFboeDJ3uvna72jem6dJoFAZo2yj684xQHmV9HJYW0HjEZFfGygEfvGpUIbtPg
dQ5OGMVI3lfUXlc9gIOqPB6qonOZjOzKihOMuyO+5D2GPd2rzpSX8jyQyimwYFxC
gVi0ZXyhOFzEemztuVsC7HgoTVD3v4+xcJY028u1W5C0w6QKgTO/195khbdqycsh
G1QJigK9YoKQAuCgBh5fsCVrinYoYM/Vt0w5Xg9OggVeEA6bhhH0Nd9QC2Y//VhJ
WlD9Pi7/+Na8O19SJF5Fk4hu0XBGGCmJRTFUMg5y9TW2kF39DL/JxuF/uPRFyG6u
DPL75/OACprrrESiAjwp1FbQnZHETzdZz+p60qrpacZn+vusItV7yDuEW62QrPnc
dj3UwS1gdX2DUv22Byxz09VPQSNELkI5kfm6gDfSt+RDldLujWiqTSxO/P35KTVO
d2AQiEtXhOyJF49wIrK4u+1LJ4wXAz/L8rYuVdQm8liyganeFUcSSCaTVDCmuAdR
1w5FuKdgsD8th7zpDXcdEvInNZ973lTpVsAFfEhPQnjGP49zDDgkZy1jGDNHSSQP
6RpnkVB8AnrkJGyLctTPADrsaJyIrJF4S6BR3oOJUxk7zTyyiXE4aZVSrpDaQi6x
FggZ/RK4PAHZVsICzint6KYmlDrItwtSWO6msDVmj8DnN5mawc/g6eTwG9X8ol7l
al37UXLfXC6SKffp/WV66KahnxMIVZA5JrPJ7D7QffB/PrYKgqlnJiEl1tH3uUL3
tD2dw4ohmw/V9VBRj5gX4+ndrm9fwoi7b/uY/S9BjH5rTf2dNqJ8KGjHQS66XTXJ
IBD46s3arMseZvLMEMheo1/WCldIOufzYX3VznDtb1uaTIF2yNUhmdCC3brq2XV6
xSsSKK4aej+JveSq5KMTbykjzizepa71STGqMhTXmAk8hi+JFtGrmoX+Spfc6K7H
pZxvS/L8moSZElD9Dy1MlcQ8+1YcqGek51Ol/CCxQNSkmqbdMHG09BDN/tegc0+7
DIVTX+E9lAXQwjoj9hHZPbwe709rJWzYOY5HcfnfV1YH3IKMZ3l8gsXxztzbXlo7
ja1mxv0zovBTWuEiqtDW33MdiWfKZ8T7mFM3s7MQCzPo0nHaNQYoZw+KINnp9v6H
UkCE+xnMCYLRXXPS7/wnfWoml0/lkk1qRtoGWWNixxP2yKdoVFtexYuk9oCHxyhr
ZElV0bTF/FtEhtX5iWYlmuLSNVbovZJ5FJ5sBWqu/28ibWNCfBru6ui8iqhzMPvh
BiJ50kV7Sp34uONUbxiH2ECdUT13gHdFYKTMNYyMfmKvD6jZigMkW1jp3rwcNw+f
TW6YhPRzwAml+ZLgc2q9bLIhlZRuwqIoir5NcWNCgvkiagH2x8ViP7xsv2ejW81k
aj568BH3j/SD09elSxtz217dYuA7ej+vKibMJFsnm/p7PNn2IS+z0f4VsoyHk3zu
PDE509ixXYI7+LyyqUqOO7cm3ZoNrwz95z840fxrWtqNTTEz3pD7MhV0+yoLVsiW
V/TxfJFujI1mR3p3VquUjDgxgy8BXJ0OxjGcXhL77KRgsgVRjzJbo+Lr66FRLQB7
5N+Z38qhyUZPKKYNUbAJqkQvVHqWiRzJtOBpo8wQHpAbiOdO9RGBbWw8Wf4ORGEg
d+p4Olf2iQmc6tphl0jO2TB8+eOYbN2mTABG39diRKjunAYlfxx47/wT1rTwbQKi
j3qTKruQEr/ZxJyYQZ1+7SHbnTAqa6mrqJzIOgViliCZlzt43rFMC2gaRRX/Dxaf
E5o6p1HwcDwG1nZF83ckj+mRAGc9Venk8FevbrQlfcT95Qcs9N3L+al1SNI/TLAd
h7P+pFYJp8/7u4hXHOsiJWGguNzLqtgiD4LTXWYEhFYBHXhnXjm0p1gbJaQNOvrM
pJM5yC62vxmcZa51Zupf038OhRCzAVRHLF1XYwoOL2i2j2NNJrtbVBJa/jlbU49F
Ocko8+MQmLYr7r6a98Du5amz722zOLpPTleXkwg/s+IjRFtC9OPqRYLV+fJHUYg0
vcpB0PSZ1T5FUpc0twZFa9Gz3Pl8yoGzS0tZL6RbCqIMFy/n31IAvRH7oPLJNZ6g
9zT+El1OqcSiWN2Le2whd56mgE9qO8Epr1Fs2uIpF2cqIxskkmfQBg4tehwYzkfE
oSaIjf7s/cflcAXaQTQIKC3EeKLO3w2k3xq0JuEUl1fRqaCYh7aJ8wL3cZCOhu7A
1VG0b9GSF/x64CDwG27AIIzKwduUY5rlbdgszeRvgNGBZP0ZYt/IXHvaKcMAwKk8
zSzZ7/Ycs5e15P6MjcO2OEpCaFbWIjsRyTWcHooIvgOXRmDfKT/2aFvVl0yrcqW1
rRjqF3pQnHdOhRC/8L1wVUdo32Wp4/TbYyKiGyFiTfwiD38HhlFyTOPa7IlgNwqL
DvYPRbX47PPG2jfWZArLVABJL9MqeIH/UD8aT9whOZ6+wShKh3txN3vs/nscx1SL
0lTAaQ1Huma2JLTg6F14aucXiacWmGoRQ8PRnkFPuStDDKPUprUxz99OrGEMWVh1
Kbq7ApLjmTAWCmus0oXKK+35JD5BV6VbHIGlitpVLDp7DGdG967862cEUjkTAc+u
PPyZBNVZ/1qKBf1hJRKs2bT9L3IqkIW9k+qkc2VFKM5+G5J05s1MsU8aYSMRUP56
mnKIaXWZevb837e7tx6zrtz2pKuETEmmgYHDDe0lf44Cp2V6BLvOeabtbBG6JXIP
ebSRqqpvfSMsuq6pt8N8rTfvA6b2TvqBYbtn67HWRCusGe/LyDJDsl4tPGHZeqDs
BCQ8gVbSoJEBIXZfRdKY6bFis3BMeukDKPkAsba/mxtt72Zwq25ViCwET3hXsVMA
htCoGadvAYPb9ejx3jsJqBTToQ1vOZGnO+fFlcgYbAbv+ds1Rtcuw1rjHTDcuUu4
wqYE/cy+8ruAna5WiFtPeNqheTh6s5wXqHBVORVkTAgknTsVIpjUKQH4R8WFr1Ms
m4p6lGOHLRqcQt5Fa6Nm+bOuzT8g8rWZODwpVpoaysqART2tinEZjJ46yrJDImt0
3gKbPqPB9t41KiKJwO311e0auuIcXX7P09ewCT4GwHYdyDeY0k8Ysl8/prUIeGBw
q1fYUzC1wEolXjpWKhm+wJYv298mlwNi1RhUwNkT7Hh+POuNh6h2+jBoRkWDRHYf
Ef4doaZy4qsb8Xe2sGrm6S3C/1tDUYfYZryNZX/FyPjXnD+6dXRJJUIxO6BHLw8i
5pBvHt2RV3Gv3TtkURSODlGr79NS85IR2FYQBLTdOEzdheXFX16E3Ng9jyu13Voc
omBYY5a7eFVoIQdVo9MRO1EhoEmOnQ36dhZGfsE/mi0b3I4xisx1nKHb9G9PgHWq
eVAeV+IKPgO1Ko4Jv0YTm0WfruJXlwkeMC8Y3fBYE2wgdsNunsEwAS+E++vT23qb
HW3rn6WNir9YpLSHq7Wwdjnu88MR8g+GSrAUARGbuwGMA8WE6rrT5gUxc4F/C6Wa
+wYLpA3R/opzL7kJL3WJd0XU8+ayT8BUhr/LP2PjsyyJ6BRCylsDLrR+TMuDzBZ3
Gj02kqagFtbkrQEfF46ZpabWMGe6aF0Uoabcc0z5MheMRStgslpvoEbEPJtXVeYE
Ah2tVWbyECG/AyM4FCZfRiBJNkxhWoiNg6GnA2NmGkaPvsBJzT2AAEe92rVdPb++
G84MeDWdiDkxxuEbYN3D2/BI4zuHsvhCvMcFaEesEyADpB3h/hZjVkAk8qEc34K0
CpdZ0bcPq9nc2Gbi61Rpj/CDNHGQOZzLM8+sZJN3DKx1YmaTc9nnpl4Oqvp0mR5d
CCt3O4moD9lOpQ1hsEc/HasfxHOamp0NPWM0qxADjIyC2OvMWbF56EjFcJJ2/dQ/
5CiwgI4UGdsiarR1P4wthecZV50FG2WAUkwPgQ6dKkFgvCFMfn8GdW7MhzzupjZA
b9+PC8HKUvP0RIGYVfHrz39pfZQrqA0GttWMgMvu2ObLvmYZl5gjXdx2isnN5K2X
o9tFRwiQQMwnL/fF8X7EDzIvU7qstfYWTAmteDSa1W3F0Vqywg5AzPJOks13PYjm
1Ci+bUPGi1fiRfbAtEYgtNiRNso6MwJFT+PlhvgmlopA1KqyQmLq/kV/Kj4k+cUU
MbRWmysoybnLtt0LjHTC8xLJNnn3VCtvAKQH4Cax8b2EUqoh9nYtHDSPlKMeHezv
ZVSz9ph42C6yq/1cmRMG97KuAJAhcydr9316lIkpAb8c4DYcI7rUgso4HdzDVekG
6aqcpY0T+2FNKppDJ7EmyDjS0nSzm9eb4Zgu7C2dyBAj3U8+6b0ajAc4lGhxgxC5
aGb3zABy6yK35zaKHaMZyuIakVDal2W68XVtGFV6ZKLKCxNY2DcG20ZRb/Vvt15j
mAVi/pUVq81fjZTVfUQdxnWLDEk5KFJHLcPvRCHqr5/pSiIamjRMBlueIP889djM
i/ZIfUY3AsDn1DYMdoP2ffTdAoskd8UOFPJzcgKldnFnoHyqE7LCja+WEQugqU44
dW2J9D81rCC0DggpaO5m2deOepMEeYbjb4XYLZrgJBD4OVTXSZ16usg4ng0yZ9gT
ZzOsfRq5p9/PKJsyOufb9DS9MR/nA97/LjfpHTSP6tC9nbXxmeyanBHy8KtVmppV
OsIj2Qn6qziEh1LjhPc7bnG0Od9NbNEigRSBxxXNC/lFrNbVz9bMVqgQtRAX1hcw
n3+3RbCyNyUgoYWNAymoyvE7TwQuXsXfTw7btvicPcXEFEEpch+HnMvdxelUa4CG
TJyWMewAYnyOiloMuglVq9Bnfupe+YUOZ3GCaqqnba9+03bw+9HZl7uvQzTrgX0E
5oBSBjj1smxfrjcdtVXfNub1yVwUhKSAO7hkAFy+tBTuf0ninCQbzQubilDeSbNb
Lge2asI+7ziuCXDaIOVrBJ9NMiAs83GRDx8wVZAMmA+wxarAyp7jyIIEF9ReDQCB
y7k+W7Y4NrhXjL3TC5avOjjK38DoHdwxMg2pMvxPu1LAPm1BKCtMkrW46aB8/dZ4
e6mFesIcBlf6YGegS3J1OKc7yRZwXYvq4uUU8iuAtYnSfh5MTtjpHzD9VOc/61QY
K8tPokJXduqnS0d9oISUT9p3QrgMkOQgsD3Nf3o+qpoM2pTb/QxyMfap9F3rkIdk
13uu0veiPK+2EtoWd8vBllliPtHkKyGrD1aWb88Mng6kww8AQ4BRv70j9AZ/kcov
ea63pFv2lDw+IuJh0qpi+kQNyoYmhQBSQB0wSgsUq2k+AhjvcmgGDM7qB1KXbw+9
nIaEyudm9TNhXpIEsoESnizb319D5HYC8MJi9lQwQleTUoETJLXFuNCvG1dVxazi
ffx+shKhYOpldvDFMpGYHNpyNF0IgbtYiw7aJvPeoH4WiCSHNMAeYdkaaicLi3pK
SPHpb72ly8f1LfpN23T/wQxiGri7xcecFTFi6QHmBQIs7wbp3PDSfb4piKjtyvSo
MlSSOoUrIWERJ9LUXAD+4GLUsPNN2hqxhQ7yWeLA+zduha9vGQp6jXW4E9JycPVp
28SXChC4kEaDGWaSWjQlfVnnddIeufMgYBUWcqEy7xO4tNscHxSpHeLgmUMiE5iS
e5LPnDo0fzi3FCL6xdreaIYZ4cenTRrWCDKUgN0HptKhcJIsJJGU8XRj8iZAxkPv
2ECgL5SAfG9snPbU6EjrAvywyTUi3V5MIAh70huvgChEYZ2JP1xGSu7FStwQ+MNV
BiXup8hFc65NZlUHZvHY4dZKBWiBEXWDRBZ8JV2cOtXfA8jCV0SAf3s8rYRoG22R
M/4vRBaKWkdkcAcW+nzVVibub0jTABYx0HXdF3tzA5/GK+od+u+SKcruuJ3bR+8M
1KynXyDri+yk7VecrJoNbzjtoKz/2HX4/YQjJKlxsK4iYYXDE/pQiQkqYptekeXb
R5CIn8dCDIdUYejABD/tuQewsG2iaGK04aoLU5uaFM7Qw2HSIdveo3QGQz9M6p9m
GrW7OIi7UyYcXFfeDvWlQ+WgNOE2JqXrRyGLTvwHForVxqDjjAA2LtEN4eavGRSI
RgpkcUVxqxlI+fhZGqJAJX0huILbihWVtZ7KhEjEneiHlnnPOXkH8h2QVQqCAGS/
fTnrHSb1yb2fYVOjaUZdqKJHNgh7+I3Of26w0Uqe2ALooNVHQR60cLuMsbvph3K/
s+amAd7A8WgGnBN5KtZYHcD1sqMhlPp4QQCX0G8Pe3qoDAcQJr9bbYTM4+fbyDwg
5E9wVUMs/0iM5gFaXOrvbyjPm5C5cCi8nvepQzN541lpHztDV8Bqw+KWZsYui/3c
7RKyHGIYM7mvf0xKtrDxp/6XDeL6cotWty++9ttTXaoPI2dnGUQRaZcUrLJ65jQR
km/k2c0npXggRT5QSanRnU3cROt9OEjpldSFohDI/GJ0ta7mYMitZIR15QIp7LeR
H7W+eIOzA1LO578wX7rujyF8nHVOiM6t3qk3heiWv+AXXFJKvSUylvuQLESuSDOt
F3b0Fi91zwOeTImeS4fnTL5b/4DvTGwipRPyDNcBpMAR4hwN7o00SCUGIQLUAMnX
bFkIFmQXkTH2jyExM8qV486f4pVkJy3Qd/oMReFx4+Ogv8rgAysdurdbCVADaWZ8
D/CtrnPzbSxsx6tL8hFtoXULw4UZvMJtTQ529LR+KbbRXVHy3w7N+Wir4p7qGWcK
yc9O47UAWsNOPe5wulY2U4tH5WT9KOXBtSE7s++j9PCTzyZhCtlAb+dFcOmeF7xL
fp6MJc5ZK9bwPBAVWtJCwyOMnDjAlEyR3YvovF7vTdBMd0QGSe/shd9eU2WXvDlS
tjGSGysVQyC1qFLVBvMRu5lnV0tzfcmpvVT/8n2H1HMQiau1jcgMAr/LbrdCPU0M
cGBU0FkCQYcEJ+k0xzqEm7ILaxvwDYyKmV7kgDIC/g+t+cZCiSW7I6S6j9k056M1
Dq/3shrZ/V61qKhCGPy4RS7O8hnePm7A7skXkaF1ksDOs1kzfWxFsIEh0jXpPBuv
ITmA5u0k22YMg+cDfaIXNg9XbqmcZhjncTga+NBEm5oIuodD68r6VTwcDyL4upS0
8+pg0LOJw+cIEDH6LspwQEkr7OjG44Hthu7zYKeyKfCPuhx5C4OV6o8MM/npObTA
nF4zCl2VUynzU8BmETP1qNNVD7QE4VoYl80k/fOdy75i9XDdOf38c8DUKP+HqtQ3
yrb49sXcBBMCnoiE7urDGuuRNMWpY1wtgw3IPcuzz0e3MhKTN3d67hj0BiqS2fSb
R0bc1DYUkHsXwe8tD9y++O5nA+jDugKeRxXwh/ceREiJmkJmWjHDKeJGuKyB8TLx
/TT0hx32h4HnT5F/hJ7CIhsFNr1KVGooQ6cBedf0M4dqRxOyNYPwZCId90mtBuwW
tI7brSsrMsgA1b7NbwYQL679ggWSOrIfyICgcgQU9/qapDpTwFVzXL2Uf+FZR7T7
zHLhNSMrzAxyKY7Ug0rkmGTBVl5E/aRIhmwvy5ctMzGlczN02x+S9r7GHLHrowrq
cPdg8rZo2tYKs+mgC9OfUM9HgdQGz2+5gplQPDL4snfXKskvzCX4MO/xawP6PcAQ
yQZDMetQ45ZcZI4eNAgtrlGbZvw8RxXxGvjawcR9bJoyuYgJ88i5d8uvGB7sLzlU
X2YsluqfgDK0JP08cBVfx8Lb/7zLHwWSyDjNV1Whae8vpVxFoC0Wg0ZD5bETJxKJ
ECBNQknCeVCyep22pC6iFsS+SgmCxZtvgSE8ii7k9e/jrXMOsn7lk7B2FBt8ITxL
bXxdvjnruDa4UuMSPU6LXSif8pcbbC1Y6eTZ+UyaEBAHS9zKxP/2GUBknnO8GDoc
K1Ten7hojGDy+Qetb3rQkKZsavm1hg/IX+PxMmZAK9ymTr6KsbBkAkXcaITs0j8L
pK4qCNTS0A7DJq/clC9TY26jnzXAygQ2CFVS3VLQxqoZVXGcFYsH2V6YR9JGA1co
camlQPhZrNuXxWOBwDKFCr+04MyecCG3z1cWbs1KBzZOIxnbNQeJuxbccnSm249E
lhP/Q+4dS/+j7b5uSY64NL2BNRd+EpaKCqYbKKs7ksGMRSAY+mF1U3P48Ru9mv60
V/YNvJfj8qLGWXgrqwawpGHZlWbOdvIqMjm1SbfVUdshR1GrlwXFYNbgZizf/+aZ
RaZ8bbclT+HBm2nx6kbFjXoXTjvSpBqg7Km+Bdzp7PRoSNRZbXKy3zWDYJKa3F/Y
65rK9G2+b3W+8Oi8ssSil0bV081y8Ha4UAq6c2IIdmm4Zt5DteZ4Ebyfoixt0o/Z
DV8Ip9ngZlAhEUZFHAKZhx25iq58YGZcickJY3sBNQSR42cA4j+lrQSogNlFjVSL
xYiKzodhbo1Leat7/OX97gVgZedJ49mmleb8e4NxkFhwnUDkIKEAzPaA6GkusMsQ
jEGt4veIhsq+qD3Kk6zvGWZYm+XtLaPOexovWB1psV2C2d7yoK7uCKJ/0fvdCB+A
1nC7iD7NHuVajSSUaE3FE4MThLDKc404P8cf9wI0g6FbtZQ+7z1xNLQCLu5e5E0c
SSFhML7hxC1dOIZrAwK50/XhiJIGxIhc8G374l4gPkMQKUGCaVFR4Rq2kUqLKuj7
mGNcBOVNn1vyKT9uWVzcXFWt9KRLEXZng0CN7WZgsYSzESrE4KmR+k+wO5y0l5cr
lueTqWiofzKF4vVksz2RNAnzSOC8I4utr3cO70pZtclxFsKDrCm9+3eaZfK4OqNH
xp3Wqgdx8JtNZH2GbN0RcEW3PzBpwomPQam2pCke3Q+0zlVJAum9FV2uVQJeoRXp
w6Sf8+r90qPrucOJz2iRvHtWAk+3qQnCHH5sPAZnRvG9dz22L+Y34hornk7diYeT
/i0R/aqWN9LAobciHH938IPxxTU9FVDxdwMMoAoNXb+OhWbvyGBnev3PCPcwSVME
wOowknu+BN7fmhnqDCbuzbO8FY/gCt+Uwrf216q0rRlnp/K87V4jhLrGB2KL6RJq
NRWPV9/djKXOp6VXXYcd7NZ+9wNPniwFQGUpi3rt46yFnU2mEPGt0joPNlDP71rl
mFTbktYi0F4ChkYZO8HErBubIZf1ZN4tO0FEXtiBm63K74pfOLsUvofRmpvzMPZ8
dzF6hRYeLZygEGdBG6rVzHrYEAv7T5DXf6FKAKbdTI5h4QgcJxTMOSXqI5b/dU3k
wE4+lAokKH3/SseMZkUCGUcCragpjoCk2ZOHZdm6NPthAoUkplublfDrWAW72ZEu
YnNp/LI0XPj1QhDNji2XZzf+QrbZHLm/VhYqQ6RoEBn8xg2G8uY2F2rJPkp2Ijr8
rZparpaDhpzOmnbrPUX9GFAIYT6Vou9rDfbayYQVI2OBZLfFg5w+RbzoeINyO3lU
utrATGVu004cwvy08vNgBVr21604ZPXDBb6c6xMsKtURQkcOKeL1T3N3Y7bJmNCV
ub5mETzCYfbIZPLFUYLweaHPLFcnGTsVkl4TVbGU182eZ8PVSxu9IO1K3sEKgp0n
2kxKfDelcw+mz68cA3KJyl9ytvDBMJVgF/cJFturerxn/o15q3N4WMz7nPa0pglU
9BhO6WZbxg1WWu1EP77BO1L3JX/i66J0t91nZae2rbg8xWt504XuCAOsLwS1/5wL
2S4D5SSRt3AJ0X7d3k3VVa8IGeIeaBBig9i38J+ek8KXYGdUfeSg6yweVToLVEIn
WAXiug+uOW1O+JQeOlDbhckh4K+R8+Nk/IzEhB4ms6zssKDR0wipEjF0mpmHt7QX
eZhk1CophLJvMyMyoi6ttLRvVb6PKoi6NjhaXYg97u61fPPdQrfKxZj6CrMd5KaQ
9M59Prq9Ib6ODqoilLuKoptjLm18FmHCNK+CUl1y5KYUGcPQuz2B+SmaaGFfbmZX
CQxRUIYDAIzr9uJbeWC3c5zr0rqZGrAKgC4TUI/CJv0CrtGQSqR8hAsN8XWHn8IC
MezXObmMSnzqsSVyTABSVa4Iv8ANAosWtMOSxvxj90+2CsF/iT6IOCTCWYccfOyv
46aEFq4FTnFH9O2r713Ra7lkPWbCJXtiKecr9FuR2H8Y/s7NDMfQ3Ihn0YsYyjMT
GGs5v0+GGpiIzBplhLW4bNr4aTvLi+pBv5xlV1gqf/v6quCh8kG1JIhL2V31QeDs
rBJX/WxCjy/MzDR39dfqviDyRB03FZDv+TUdwvx6ByH3drplYlgbMvJAIzM/E1/H
QV1aP5k2gp4akT6lHOb6I6v+l02KUK0R/Np/CElD/wJewQnHKT/6+BInj6naf8N/
iv1M0C8HlI+xD9b0zBIL0YYegcd2rNcCMTrfdg2WNbq0io+0T1+CpeX5Zw5W1YXO
T251u551geAQih1XKKF9DUjphHmP7AJ3nlZBbT4WTnJ0pF2RYC76HM60Ijahyxu6
DpxEY3YlBve8ZCqYk52dIWFFY/Uzc+jzn1H2wXq7Lm3aKNYldlfaJ1JrSnwDN/Dg
kpZnDsMfxUjE2mNyljlfuxj2QDDIdnn4vXsN0uLP53NKMFLPGZZ5/1OeCovbhbgi
75G69Yyh5bEl4q3VbidmsfZ/XTSCtMrRaWB4nuWJwe93lAoVHNxB58JU3acPouMJ
fwbOIuanRqRek6bTyfETGWzTHUDEnyP3+CM6GGwyNW+o5pt7+YywPFnFxzv+pORt
4Rvc7GFN2zjAwKbR6NNXlWvZX3I1zVkzQNXEsWJAc82EZ0bOTUwyM8nZxe0X4OT1
7gMVz2WJL5qSHwWJ5WtM31bc+PLMq+ZjdfC/gWTAdZ6FZJ7Fd0b2rEfAAOKai3rV
qiL699QudajDGmVvdwDU78XdWketZgFEgWrcVZtVUb+ii6YoAb61Azi1J6rh6oou
PDAqEhT0Lzd+6ge98vD8ZzrQrDFRQmtlnr1ZfUIky8d+mhPPAmDnuOfIVR1WlNrf
iu6KWCB66FvRYqPXG634gC4jg0RXGaND8LO+97KO8yu5olyELD5GT1hCdzDDP22s
Lz1OjKpUWA2usaCsDIE2FubBgnEWYm1wD+TJy7x/AtPVDLx0lSBqN4VtRRId5x/g
7iISqLwnQPVuoI1hFg+mOW1Fuenj+KC0dhC/CPPQ3R9I5mFLzNHMT909snE1PObg
kC4Vc4+KYn59c2QbjCpEJ2h9MnB2ScP5WnuLfcuUTnWNudMEEiRL7c3jrrcdQvOU
+UOZHEGdPI9ii4vkBi3FhZzsa+3MAl7noR0krI+01Udsg1OVW5E1NiVGQFPkuJQJ
a7+daxT5DogLyJ6+doX5mOZc7DRv2Gzcke/xMoB7RggSof1ngWCv3zly2TdSGE61
dDfW90/ui3JP8XnEHmvfrntUXpoYSGkUnPwStxbR0qq/1jYTC6jpqU6dbrROSKvY
9h5MlQyZtwHUOa/xOXYll3jKsIJoxdIO8sjtTWh+NGPZirwgwl+wAEybFLvkMAMs
qsgenYZH89klp+bqKmgq95KD8cVC2cEOCS2Ytfq6q6SY3HVBdEi9Tg4Yxr2E6aMK
bcJC4bhSESo6aSnx0It0Ryrl7QTt0GbJF1fZ04fApUEXbG1pDscnjd5ybx0Qvmr1
kaUwCijfZm/VNB3wO6TFRJ/psVhcfz5DnC2wzHrvWX7uY+cDLsnm3C/wnxmNW3cA
O7zFV/Bl/Gd6N6qybdNp/uGvjAD/n1QYihypaoUAVyCQJ2lduz5wxRQLIaexhaQI
EuWL5KnXNDBsXlJ+fj+ImK14Z3niy7+Oz0OoyeYXID5xmQwHGDtYQvIPeJTcCIrK
S4ivjlfTJh9rqgkmMtWjauAVhn2y+OrV2XUXHzwqZ6/cWIdq7VozMcHVGXVUnDyc
I29dT3G4nMldUIOtzuuhxsYDElToi2U2mGHSt7KUfmCJ4suMXrY6KGQ10tpnU/ry
LYHV6if0CLJ+sExFX01q/w85+NDodi7qaCLiJtAdRGhvZMzcDHMmQ1L//my64TbZ
tuaTpYGAlMU0tyx+UkFmkqNO66ue65lNeWjY3fPtHQDJiOkXcWg8jFOR+6Uatm1f
vIJcpj1F6u+9CowAAIIQuCn2PtX9PkkcBhEDfptNSAK35qzYQ+TAGz1VkcBseeg6
S6qBKgNBlC5xmaNbttjiLrLN9XOVJb+VQGD25KLg90Yet4r7WTsx5UlSiqoapMGy
tEaGtUgkxcjlu8D0aBMCpdd1jX9/v0dJ2LU0ROlBXiK7smNAhRLbfWIvfAw+gXkg
6whKiVqluoehzUJRFY7v2F3brTVGidY3Mxcm5rAyC1SVCwYzQq9h3frXv9rMfk3d
tLRX4HDd5INPk9ZPo35Y66kZzl58QVGzDto25X5yFgoMm/IAWwKnuW2p0tZVZolU
8NPyXADEVwM1GAI2cdLve6N8DK333RRpRwmCg17zvNa/aA8+F73KPdlMaMSFwNMg
FBSyV/YHBmdEb0/mg7BglabIVkOZ4inpAQueg5w4KZb/ErxQN7uyA4hqdMlsUuPL
TXnuU+mETgnf6x0ciojU4pxol3vOJwSgc1Tab9rGyb8SfDvl6c2QZkr0L8C1cqfC
o45VYm5RhmxGyi0sZxYVqJxJAddOiRR6dVHoulMec9YQY7Os6Vb+F6Ztwdfj8xpG
bkOJXrwFONbPotW7SvyNCZNW2/NZIV2TCxSEyWKIXQ0Z0W1ljWw8lstBdGcrAt3b
tXj1N/1uZHa0WP+9xUkTBknzxDAWJG7Z2nubq33hKTziZ9P1kP8det669+5+7ZtZ
nl+d3RstFgkPYak6YUuX956Q6jOxDEgDoAdtIzz5CXWemEwXUZK+E4DXV4eKw8EV
ZVVET3VMGgHTESzBsuV9amI7XRUuOBwt9pv9gMv1QApM2aSt1tUiNVSJ1yEpLcx0
shr9jnOUBJKTOtLmMDdo9AufS8GuhPrrtwpqyN29TKtPx67bfOMU8EgXOVL05VHC
CD8MUHtLqksz+vhrXVmc3R+afkX3bYyHN2LLuWW6WjtGzWzHviX9apO8SrlVp1is
3L7BCguwAWrBBgnTUvvwIL+/U3VEqaF2TWqifygVlEWEiG3ok1wyAbgBEGazgAyJ
ychMyeZsDR80yoYAMm9fprWVwA3EiznHgr6dF69W7wySY7+H0JylCCzeG8kppobb
IO4gs3MhFH7WIo+EjAdF7Tbh61gX/6PRbcazN/gHV99+fGKw23JvyNQmr4xdw8I/
epuJfDuY90sJ3kGV8qcfLht3NUmVn03webwoLTqkVlJs9VhBKXiiqu0kQ1XZcd2f
wzHjRAkmed1j9uLFmKU8K5j+Z0BXjkmDvn2m7rmMg3trpBrkFTQpzhdVVze5VCfW
ApD9DCNkg2e+MTlqDmtJUW359wqrPb/s0Kbj7eVWbuSnvLZeEsMYgKjJ19lvVWV7
A8ACkEXciKdq4nTAN6LsC6cuQn1RrYRTORBUS6KOExMwyBtBE+Fjxnpzm4CtCPTQ
I5jjFMMkLiSYcjmt2F/Inty1xcgEf9HljZugOYIDketsZJxvjvKJvLmPJmrhruhq
Q5nMfdovvA4N6cp0bKLes9RrR3Ignysdl7aks+/am1aPhDpqKl3S7Wj1BEdAGxDP
UB8j7vadve3Wbo/6KwnbG2JfjaJyAMPDlkcn+66uFnLb46kDHhw66zve/Miz21Dy
QP5QYdwQDmu6FEWLqDtXBkwLFvAquZGbOUkttRHPDU1WUGCSi5zbXnFwnx9kwrl0
b2nEcDqBXyqHPtP1zSqvRttBzR0FS7Jv8TSb72GLQPgr13GEwjSyRU7/dGMy1hiA
/1oW9gj4NnZT1PQw+iWEvUgFVdP312/a5cz2L0/ZIg66/16TZe/kzgSX0xrSXiBh
3ro8QA3RAO1MZv9LZfmVhp556JAJkarj6y4dI5kD1ZjfjSSYdzxx/cKrr5gHHrM4
JurfFbqvROQgQ0Chi1IT2fNo2wMh8yJFcdUekjBGrls+OY5QHQQwgL80juIat6xL
m+NUhHmZ/fRL46tY0SfZ2idyizdDsAsV2sNks9kRNuiIjW715DuL3V5krGwdM/lw
z1QHSNOZYsuibtxn4kZoB9wFOA5i5j+cQrpesBztLk2Y4AZneN8rK737I5s4nnFz
NHPTLHyGtvoXayM0ehGRT64jZHuMdyKjMl29n2LaJmpPUOhArKlYTAp/CBJtoLaA
NT9w6UAaiHxbLPHW37svqLoeDEhbNFJyyZdZr4/q3tZ0RoYz5M8XWqYbI/6/IvnD
0S8LRNzUFirmM7u47q9yy7Tiief854ceJB/rXdpx6tE98fGHAzVf/jorkk7TALJj
xLIdwbQ9v3trf3vmEMmQZQYTD0ZMfi1j1EcBKwmH0EPc0RG2CI5RuxrncWVf6W3X
BLkeh/SGIuaXv4EiRvtW6unyuEFWYVEmdjxbcgCwOlRfrqlICgvYS4OFhfNZRS9A
7JXwxaI9mAduMO3f90MZYI6qxp5ThtlwcmtX/Bz2VHKywZ14mQDYPun5Wc7XOPpJ
2WUMin5WDbZJ5kBAjjOkbskD6W17bJbUJ/iCUTSEv/qTt89iPtYbWrigarIhqKA4
mt5t6NCVnVdQVuva+kKk3kh8mSVI/HzICI87zdMrFlDJcUmq2ChDsEAOPZqKxtAj
7+1nY5pwl5MzmhLUbHEwWep425e04pob7tTPMFlahuKYHByDVTdJLdhmKJrikAcu
hm71Jrt3Qp7iWoG0UHSUctRq9NKf9fqCRei1MGyKuoaqerPN8TKnjllibe42eoOw
7/QuSxNun8NpXGXxqPy0bwpTHKdduaCDMSZ6DPDXXcG0WqYeeojRA0GHvQnwmiBd
woRssfn/wVbn7uPBHPgSIEHHoUNGY3FoYrpxL4FQi4L3wmZMcRcT7z3kWYqkOYUr
XqvHQgA2j7KchTzhcNsdYOM7EQv99TeJ6ZdegywNkHj+lj+aUtcJvCGuKjMGwOop
eIZA/5Zz0VorDpcg2UTFomjg2QxeaB7nJSsRACVPWccqF+AzFeTctEm1GVxVsbDA
CQP4gykDqt/SDOq8CpGH9Hsq/7j5N14EV0xaipyFYE09Dynm8dcPau4Ign5snS+5
KwvTS85//SDecVte4/NL3usbBYZN8t/zsViz7V8Bt83gaRRPu5oGBBfAACFUrI11
iH8rf5S8KiVgSpDj1pN50SknADT0aR0duMEx2NaNT+1AcqKjXRLwuLatbgcvg02O
KQDLBPxrf5/Em1f8ZD+7ISFWJHmCE/sqEv7/6/dga81Y5OxwubGFj/9Yu9gLVM0I
fijIX030CR+lq06q/oB+rZnrNRge4+2gNRsqC84ciTfu6H4kiqg5skNr2zeINHwY
341rAvYC36lOCmuhGkdUUfpeik1aLDiPXoes4QEId4+siN8LT8+qk/uHy/Xgdxr9
WuM2564aj+culwAVB4F6aw1RDJr8wSOFDP3oQAVm4I6irsqu1Th182BkpHwCi/op
V6MDHLxL1mkf+COjxRkFUoszMibMtUeILBwyQhKVJvulFPLUoX1dDs6YZSKvaPLi
A+y2JsoWpcjYEeNpvA9ALXZJiJoNb/q10inu5LDUyonwZDLeUffpMApOd7wLgwX0
nzfbjAGSFenqPMFhU7u0Oz+JulFoyxK93Y5joBmUvoZ8azXWGFHautbWZpeCZh5v
6AT/HcHk4empHUlIUAPXPOm1V+ZbqsBPFkoepg6uRM+V3BH+kAmFS6WO9fGpcOoF
ls+TI9saunf59jGwNffTPGmoMuK9y0pdHaUw9fok0EBO7MbP0JuF92iBVKNr/+YW
gBL/K7eL3ac5/PcfhDHv3ZFQ29dKx6koa8zKfICP/gHD/9HjveYhPP6NHEdjV/eD
TwOuFUXlW0WYotILa9D6qStPuJ32Gr8+L6kt7rIhfDJlPw/Ta53nIPdnCAf6ekhn
KVz7JXcTI64U2z3y2J+jqj5oIl1EwNNmExFwUjh3477RCF6W1r35isfc5FIr9FzV
KKl6eJ5GwDIj43kz0p1HUDm8nMHiQ0aYJ1/1yqFQSQU/HomjMdWBGk9bPifDHwG2
N57BNJ9rkqxofAHMA65yPlzhEjHa8xe8WGrZSTpqm7UXpCeWTpRiEv/TilKFW7RV
oNoHPHbg3Id0jWj+NZEbga002HaPGOkXoQwkiLPQevp+Wl5q3zRXqFp5Dxl8Dmll
aSQ6Qf+A3bRzEiZVzFHErgc5bLpD5UU8I2JpXH6CweMfMMlwNA423+TLuhIuNnjs
Yg+RPoDohpzW2Xy1bDeQRBYUfasQNN8co4h0jG5AnN7hwL8AZXjLS+4C9/n+Y26u
SbqL+ymzPwhKGdHcsF5WEiaHIGtRWZnzYlslUvVpM8FnAUC8+hBqKB0PvZdWB9iR
Bm4jBJ5vD4nnnWbUhFUdsFb7G75IlE+mqPT9g+2QerT7XwbFzEgSAtTHp1Ad6X7U
fNdhopNiAlucwScqhRh7ffOoQbkO9MXJsrF6b3gKvuBErphlyuAqgdymjlJPS+KD
94uWV193bJDC15SkI1GK13Cog4NZygCQac4q5XQQwLupUcXb/C3TXUmG6pwABFqi
HuJ4zxO8p9fIz37RLxj1wzWna2l3Xm6QK/pHqaRxFo7pyzP5e3N2qRw552PgPbVx
8Htet/SlufhO1UZPr62yMtAsqa1fIG0mUFKE3stuzMLvD7o364ZGurJNOHCaJQCU
wwuU54fIHLox6Qk+6/3kUJQtuMfXHy4u4aCBV2U4TljvS8YMhehcI2S+ra9tobnO
U5g91PpTY3guJ7+9bfhM3Tel9rNbBiPvydL+7wxDSs7R4T9IgtK5A9AyEXQ+m4gz
P5HgxOvjNdGNzYs8/ETFNKtZQAxtRaAcfh+aDw8QDVWjVMPxuZGIhxyhMSp8w801
iy1qvxdFj5VNei4jj/UxRHKOXrZK+4Ck98y6Lnp5bHRXtMZVKAqq4FlDcQpNNLNI
0tgIuaHGUGK1RjO6JI0lW81LZoJJ+HgY+nN1iSzsSA56jdOxxMwlTEtzT5F+3/Yz
Wonumnu1x2diUctNqMewXKIrJJrMWZrf58uSZsHttg5wkiaGiYAljHk+77Bb9KZi
Xfohky8b6YGPQhXt2VNZUf9pDJPsBDAMSPzEdPxzPlWkLQ4by4Ek05F5vNshPKFY
coyN29nDO+K7cvze1R1rTu25MFIManKRzJiJVNS+pd8McKSFWt2Pn52eQ+uXkRoB
HarSZe+cm27zlV7hGW0sgmIvd+0UA6jjywNHjLWQK9KjtPcsmeA9vVawwQM4cYa+
mSKQlMBUrXmC/LkL8PWJL0rkCJoZoUjAx+1jtnoLpvkQn772ICRneCVLaj1Mlikr
JbMgqlwKArCcsFhRo4sBqdKZxcFBpUGEQIUeXBdQt+fNeTrEpchcaEyjUeKjwElH
uRb2vKiFhcdZ4qzR+YlB4C0Awfyl4cOxTRuhvG90UDiUTfokUxewPVvehgveb/l5
IvL5lvEfw5m6Y90xPxMI3+OMO5q7J7QegaIggIatZTR7OjY9ENqZ/NxfX1F1/TtR
Zx7/62NqgEqrdKCOIPbpuby9g6UBk53HDXGdsT2zqjALQ7OHU6EedpY5EuOgTlrE
P6HJIgHcWAtT5/967ddQlhzNUiCGt6iAjn4FsgFWoL9ZIZML9f5sfXz1p55axLR1
6g016UNVNl+ajE9HLKaU+nG+OBxpO07lq985Y40sMDFWCwfrTr3uhUIpkv8Vhdjk
+DcOibS7cVhDeiB/d2fHaurXOHEprvQ3ICOPUNuArqZT4+uGzLwZ8fZigj3+XV+u
n1HAaA86zCL5eTUNE8UGC+636uN8lOohAlvZsUFyPvW8GocLuPdYatOlb+5fMTHJ
uNKBftnYOgzd12I5+3hs45npuRXfkPQ42xoH1ntANSU6uWAeFzHREnx+Ldj4abHS
erw5x3TDinMUFQ6DMfVRK/zwj99dfdlaQx6HhPSzaYLE0ffM0qT1TjF1ed4OXDQq
hJlFVQwqhvJZTRVZ/abp2lcp5BZSZBwU4nFtmustWpzgx3oFumxsDFwNacfZUrtH
x706hZleN1pRP9gayyiDm/Gm5iS0OTxUXCt6W+kGfjzbAC4DKOatYja7tD0AgwBh
NNvOC0PzM2/oRuwQ+kb1CrfHIvMIEldkp1cZBVSJWmofFhtwcXw8b/ZNxoexUy6c
bo/X047uotPtAIuZ+jrT1thAiPmz3mpPkQlKRxjgwexSJoBcRDgHiCra7ghbzbA9
c1Cof6dL6BbCg4l31Oy/u9a381YvnWWLw7O4p39qFUiQBhUil4fG0v8x+LkcOoC3
TgQuateM2nGuLgaJBvgJyWpxVYp5eWHNcHK8WkdkuPtwkDMizWBS9FgztPVndXFu
lOgzelcqFJBI8aoDv1Au4N1G/9rcxjqm+kTotDoBAwLrVJcyCDxHRhOc1iobcJZj
LGde1se+gXgSWaHBcaR9tm/puh0G6sM5Br6GQElQMcT8hKVYtzKtE0pTW4Mq8aYj
H9avM4tZh+EEqzqW7LsXtjRSF43VEf2m2Gv9tSjn8VNz4BJUkvN7HrgAijFyTAYJ
6U5YUINLyyxeE3OzYJ4E+dbJLItMadGy3H9FFMwRHCfAzuR8MWe9zsojdPsSDVEM
XE4gO4zS8iUj7GGn57f59ZZMYy9bUwXKTyrOsADKEJcLR8Iv8Z8TwVJ2t4/AMpiz
fF5TpSBAua/jcIb3qw94O2HfPK8U06SIvLXGFJCpCeN/7kOSeWsSi6NFW5ba0GDY
Gly3UEL0nHKNfJX47ZH9XsrPfRhTKVSHSZEvOolwwUhZxKcdlmQiUu6TR8W8qyZk
F1NWjSp+wJkWKec3pVoD2GgK+zRQ43Jq7jQrBcUmGbSdjrAUBat5TE7u9xOcAehF
OLvI5z5c6jG7zXhqvuWbVpaUrs5Wh7rUCaWRi0LLxv4CgfXsMQs0c+1a9pAzruqC
8RFoZuNIq3ZXWlK/Hsb7hkbL1G5FBdLhShxpL+nHC3J1N2+L2jYtCQjNAT7C7O5X
mX4uxQJLm2Gmhxnar8dGYJIRh3hlq6tlhDqkRjJ7Fbn8Je8xUucHDjZ6THuelBdm
BlKWb4U99KHk837tohxA0DCuSSPv3b7G4Js4KKl9fcJwdeQEdIJKF5BEX3d93D2e
zmRRBrXOQitnIc0L2h0kEx48U2nAlljkeJFH+bKquAllWTMOFHC3gVnUKmdtKEK0
bujRPxNys8zFpXZCvOKwKFZ3PTV0wPAwI9tuuMAC+eo36q7CQ7cVpll0XoweaGLP
2oBdlYXX3ev2iJCwAhfkmiAAwHSLCBXiYEf6OxL6oThGzw/lnMoD1F35gh/+ttF1
gBZpRqEXwBn3kqaLdIdkDqkj11pgyAOuFfQb+c2ROIExilaLm6bYIIQ4XGkvYj5i
zcVOA3I4SF/IY7BmdBboC7tmq0kpbioUySD1m3z9Y5TXrcJuwcLD5aIwaa7lrtrT
1Af3nUvZugLYYoE6EV9TV87uN0/C/wG1dClf64IFqT3Z+SCW3KoGrTIG227rzxm1
7nYbfngBAKHBec+wPMgKfzXJh7z5R6JVk7A0nfAgigXtMM9vAXq8jLupIbDb8rpU
7CUPhW/bh0dvCYSQYhmCGaBjS7cl/IrSTt7Xfl2FdJealvRYbDNApEryydXloj12
IxQTRMYCSXyRmDDkHCzC9UXnuCOp4EMWB+KSxMBiEdt/pPoL6Uf7ZgRuYBwHXOqc
e/dk17lJrrej2z5FSQ6zuRqaRWEQaftIMt9zGdh8udar8Rx3CNQZvLoX0RMapflN
RF53IU28tAKBjaK/37TTyrNBTVR+DBWAsiXLizfno4oSuWCPeaE1gWk6TiKwt/+B
X4Vi1QOn+YH3pCdfH26J4oww8kv/4nlWXyhNAchfUmovqt6jjXNji9harmEAHYBc
dRaNWWzQwnEx/KNAvNkX25eOucR8CEsdjgEG7mj41n4f4AZJTYOWplqWKGWJLAXe
LZFBn+gnDJku/SUBXjeLMgOW1EajHStUN2Ii68DUQ0p1i6idBAssoa0XE1rKfHcO
vgV9kqIqnl5log2kYs+eqAyjpYWizNfJHEMVjRGFqDu39uvwqAiVoiQ0Tikx0Rg4
uSDgvE22Q61mnLm23Rzg5ieOahNCHjgjZkxLf9DdBKk9TnVEZxdEhHvOX4QdwxMp
gozKHbkOI6gSSdj9FCMBrv1y2oThxsky+NJyP+ZWxfpjvohuQZUVoMD+g+eU+9hz
ELYwj6U3w3EYW5GVD9PoS5n42OJbo0AVzzNh9VylT4vI2o93mMfZ3+DIie30pCrZ
GLqzmz0Zs8px9o6oXWIVZerMFSrGbnsQlDgfQ7Q9SSp4nCf0kpN7Hm+XCFQJwhwr
LVzGYeoLq5hekYL9Qv1hMSDZTPzpIlZTNZa2IIWFSUgPjZt6UXzhVQUrkgwI5Yr5
24IM3CpCHVl29aIZs+12TaLbWz9KV99BiQitiKjr/dJhbsvH7oh9E9NIKMBrABZC
pwIgLVRgvDbPpGZ3HjcZFMN7sPKJt9A1ORKRa9rCdJrr+pMtEg7F8J2L9aG/F4/k
8rPevkeq/Gl9fgPS2B5Csg8N2nmhJ/fDFz6Fi4JPljv3UXQjwWMBMQ284ylEbdSW
i96f4QQ2ScSmiNgy+CMJtF6KR3GtLuU3KmqwYf3kBWHXLWor2yZFYz9XDKvsirf+
bN5XHgIdoRaaUJjP9IZjf3+NW59y7ceZbYJ5vaFqjlqtkbE2+NpSdvqcGXW1RGoe
nW/7P6Lr1Z9qaeI8AsEaKrf/LiFC01JlUxcw11fd7a6ph2p18b0AAkIi7L4v3Ojn
YHHdmBwac1dzEOd4mchL36zZvW5s+jvfUgQrPhqiJSQcLim2mI8TVfmtIXCu9NcD
PGLtKiRNxd4wOd9blDmYHRgKKeRr29y8QXdI9qR7w7gDlB1c5XMjEdNO3bMoh7Xr
nGyvsP04cR7DlfgpzN1tW5ubZuoI50v1IDXk4FTAN1D77pXmteBHkTD9uOZg20p0
m4h/pWrOjC9g3dEU0x5cj7hjHZsUEvMEPWTuApb0BV2qnRBY1b53hRjLcJmsiBsf
4B3tBBqQ61dmtoPhjpMB1U9RVWrNT4IOViA4r7KJUkYqTOaGM9dd07HuHqd5FE2c
ICvhVNF0QfBwbqGJB0ZmDDp7KQuaPgbNqZHS1i8W4hFEXxrewg44y/+QQbGb8hrK
LQt6rCve9ZpYw4PnrsqCEJopDDxL+q3oi8V4Oi31qOtk1OWBRWGFqhFzdSzOwpLF
WCP2LKa3q7oyP2I/9AXkp00FJt3f6aEnNEoCCGVq6EMO6sh0VTg/lIVo4DEBN+uJ
g+eVEP36DIPPRkh3Z1i0eQK3EQ+k0kpAqQi/wnGCJEZCLwvYvTQfM1B5d21ZrZ7l
l0GgpT80Ns6o66maRJLJZb3NceI6G4qgefzoN2JRoqB6l1hUnzvDsVg0fI4AjugO
UbMTlW3xJpaye5GMHfPSvihyp9jGB6YG17FRLI/jRX/zYcRZiVPjqWwrmmeC0d6g
TJ+Thr+sZfLpgGAN1vbcS18+knUxKITchihMVHDLPsZx+zn1ZQSa+HzKbVSjh6ht
rl7RU26n3Cf2nv2srZjyZ9yTquUDsN+x8jwJ36/Lte3qwjsgpZN++YZeD/N6PV5D
ErTP2WuYE3QN0XUB+g23SgJkjr+uAVu6AYotAMpIWoJTzi+WzkgRt5KvvpY6a6gV
3vRr5MAlA8HJdYd0Gdmj9Zl2JeW8KBshhmkEgHTGveZT93i9xNeQIM+28M21V7DO
Q7uL2i96WWjmJDrKzeVpyD1CU+fBo1sjA2NzIYUgqSai0iGZHzyeQZbZlLwBrm84
HIpgXXF+wQO+hRdhotDw5x9ze87c8N6U64qLuwqxzmbX+byo0AE/9mxM41AqhpYt
0BioqZYKdCJQ20N5aktW43vZB81jS7kxzD6RzaTBxJJvpwcQvVcim3m+su3iHIMm
p/TR3KAKKkaFXxJzg4Z10e01V2uGn3+DZRm7X17ppLK+zhbG+bmW7PXAWPmDDoyj
dRnExX5jZkrkhq8TuAakd12FrRja4ymfY3Rl3F24frhSFxl3NPrlqSuNU+I8TgBn
awLZCk4Q8pGuIt+Fxl957A8Ky26GDeh04sCkoIY2//H4PfUmoJdUNYVHVeyXWZNy
JvBBshyN1ogTBNz+Txmu7A/Hcu91tT1Llk8AD0Ic2zx3CHZpMbFE0A1IVxzTq3dM
571sxKdGWROBhKMZIBkR/u7Wg65vIfcub6xDZvEbBePyAO9NBlEB7WNJl4R4oHWd
86LZwtJICZ0EZCH7uuYkQvH6lh4TUZZ3ZHF66FnHUu9NOW00TlDizhEhJ3SCtbDF
QEOIsKRTJvp0Uhq9eAIsKEOdOZeoIYz6jmMuioi+PpwXtMEaZ+bznfSv8D0Y6its
suY6l1z8dq8DQ9+bC0gapBcry80vICZzjPiQzi53YjPu4zDY5MYNw10thlGr92lp
tdTyhyc1KRd0hlsjvKXVsk7kxV/DV4xfHVhSaiIbue9VEJORsIHWHo6noQNDjqph
BSlzw37ZpzcTBuHkyGMKkA8cNTdmEbVn5ABpHMhZVctHky9G3+kCdo4LNVTlTpQu
aPc6cKhS+6/3hN3xmZeqmE3EHOXkC9cygufoRxsXUkvwbb7sC1UBO+NMqvBKP9y7
XZL9H63KVjqDG5zRHJMhnns4NRObYA3P2+lgYAppYgGEeNkjR6jqYF8zHbyoMqzH
XFkTUApJSHozc2/LcXD/cljP8p5FcX/8gEUdW6EukNTjJhcfC6ZrO1hdUnaJPRuR
Si8ME7iY+1BHidX7B5iu+DF7ASR5kkGqmMwKbNQv8EWAbyUbVvx0edi3gV3PYf+Z
l7akSTZNeJobA0O9uRnWiGk68CDDpKkRcF34K1qSnPHixHvasOe/FJbawHStLBsH
0UGwAMogYKrqOwfVq5QD7cpT8a1LdLtpKlXzQfc+Qk2aZyzzwMBvN+fpS/KGm00Y
pkyLFmZJdAps87/swbV6UqGux6qwdSZEFNxddSWxvIdxeibq6JP8myt4Juu8GI71
8GHjHSchuu0ycH1rOZg60Z8C9KJtSiu8vAp8KxhGk1ERIAtgChT+J84ARtwqGL+W
2rAq4IMND6XuJfBxCn3P3IXqFxLVNrKEwai+6aDxt+N88tP7AX7+M6no50ukCFdu
yfpGW/ilbkuk5ic00qPYhnhF8Ag+aK9kscHrPMd7N4AZUWE4QX/onJKV56XHPpmD
bIe3ljpCFw7hxoar+ow8kcLhXPh1fa1RtMwAD0+f8OLN+N7E58iQCXHRiKkJe/tY
78C0nuiXSk8MwMK1OxMeK49rwqxrORBWUCy2dFf9sC7e3iBoSLSIJxN2/FmPec6u
HOtvWR8Ci6CM29YrKaZA3LW6+oyWkTi1jyzQedS1+d59mwyRtLr+POiQz5mUAIq5
uDeCQqCmqiiISjhLvgHyLzRCpvGn9V0FKX9OVrhD53/Ubkq2XMy321U0GDiiAx+p
bQI3uLogUT/BhZKePVdtRdYzD+tApZelhe4n0Sig3m1v8VDp35ucpzvWWPZSvuiY
i+4xiljlfS1CARQUDeRsI2JRwG6alRBFj2IEmaUmTiDUP0IJeZTBn9ERmFMatYG/
NKXZ/CVp7clKi9jAKZ972YxTT89k6hHjV/tk5wSWUJBt/k0LFvpKim5nawunPiaV
TG9bgGaE5bpjdGpgr7lRvtJqDT+AUlHeR1a3ga8OGKvOc3AbV65K4aIDjp/ZoH2y
GbJ42pNf5oUeFbxJmhm9aozI2B4RFVOKJ529vF8KP9w1PpbLU3uJseLvlpdwfzr0
ArY2KnGwc0yUeInxZN5pdgua/8qJohJ58ym64uWfj+Z/LS1Gg7L7xz33PWs4TWnE
sXnctLXpQcK5H/e9+y9d3+PZPUvKdcvtMJUATraYeRQdfCURpECYuCl14NUjr9zv
C67QIkFjYXv/fvsiWK579D3xrIzpUfDWupExtIB1G4tDiQlUlfS70xLxDZUecG5+
B5QW7hyC1VD+bP6+Ge5hS5gxR1V2kOIFJFGWDKzgZLNPtKGvroeokSkicJoDlV8c
mEKFxuHu/xLDPDwzvwWRNqXuVwUrKu6d/xPscyqsi7CajwPtVwVBCxBBsBVSdmCH
u5D4dN/gQ1uaLuWd5fUt1yXsHSuCtMWN05I3UH3kCcXbrlT8uQl4FJ9DPRXe+44I
ODTdjxAiTLxCD2fhfkI1n/fiXERdpfwMsU5ZIy5HNBPALA/S6eroIan/Xdqy64yv
bIhN6p0P6xGCb8m4GFRbB4BMtSZF6qUQsGRTn75UyYIWAEkAXwP27GGr422NMjrJ
iGVjyi9SGbXmGXiyJ+gE7NITz/IX26Y2CASA+JIKQDTFk4X2Z1MVHIVNeiv1hGGL
ELnMrGcC9qopSxWGQmtpFuctLmhzheOa4Fa8VjfALWmr11qh+oHW4goeOHYbDTJ3
9J9hUbuK4XM+uhmv70qZ52mX93C/Mg/0GgPBo93cob7pgb9hNJz538ZeNbDMVdXc
UjABHXuh82Md8M1sxqgq4SyuFm7rmM+kAuVF4OFc21hW0EbfSKDTJ+1LFsq3WDVC
nAqgiXsB8QYkiMYs40W1a/NxokXQMEK2FXVo4s/n8DBzXCQ3aoIFSQdIQ8OvSpS2
CKgPkPbZ1L3dj2SaPvEf8W3xYvYCZrJ7+VVQaPRhomJNahpcp7dIAixVAjzxqRdV
IEDfjqJYhRh2/KHV0RiV2tyDNHiUDS+K6VznSQOl9IxLIsuQZ2rGCwVT7w8pIdaz
LU1r+cdWZILSAddHo5wGc/ndNN+NK6uY7VE7SKXkGjQbyKnNrRXp8HgGUTvaI70i
qx3x+NPtvjyIIs13n9iizPmFoxzoBs/8SSvB1ozzX2NkNsjXvFFXKRXQcmi1rWux
Joq0kPBp7rg5uGGJ9IUWqLKzItPohnTgt1Qh4/sE99/9gzrQ2yt795ElOn0Exry+
qSd60+BsAM5d7QR1JLiYV0rH4ot28YnRuycRZYxJ0xwk06fDSml4wudTWQDX5+KR
xgMKRv8w7U9tJOyAfeTzilkX1j/1axJKzurTrPJD91PHuH3v4VQlz+QAiko1/zE9
LeCmCszvmaacAw5oaUgNjoJZJ2jFw7eXXh1KYEZsre4QwUSsNNmrwxZERqPPCDuF
P88pGy7N9YUyPk4xxrYSntW/oewy4/X1x+rWlhygnahE7IxW7Z88Db5IryKS/FgA
JaAzb+Jp5uGp6Tctb7veGu//PeqzF1FhV0kmea6Ju8PsUhb1g0E0xf/CqoOM06KE
N+clnpYhTbMHSk+lwOIPvIvRi+UWBtj8aWVRFYLoq98/zIv0FUr6mZLvMKctGHK9
8OkfN0pqssbLNCKd0BCrSyksAWQpgN1/5IZAdLkoPmD7cZHdbnsgahsEP9/l5+aL
fVoiu6QfI16MGU7r5ULBuLBA9oKQs7SJOJD4F8C11mOBYDYkyuRKmgJsha0HfTqU
hgU4AOcMn88Yuut4lzobeqDck+Ln62J82cYhd4p34D9GBPnJrhIZmFu9WJurJbWO
910fzC0ONVdw/uUwzTsecCkHZV4qxm63JDyJvhKktHYxikfDeBAdW1uh5fzajTKo
56+ztLEJcQmoyGT7AtYTRTeRjDjMtH78av/hUv2WcuMsWs+F3F+J+MCVU7puqnKm
s2zB8GfwE1e/A/kidxFBjscOMspdzgj7azWlfDe7HCUznBi3bz+DZdaIHFGuKwXF
d+PNlRcviyO6imdR72tJgtRDDJGvWzHzdeQlCw0z1goKsYwSicetNInOffTDSl05
KCic2kmO9XXoT0h4Wu5QjaZUiYitXH4Gso/c8J/Ba/IrXW5Geh2J6aYTGp/ioetk
FARWiPJ1q5n2GNBsru73xLrbZFCR5x515COl++19pQKSqHBoNWFddSspJ/51lk5z
vkUxApUXxYV2MY8THeTtJe9t8aKErsgvpHVAvh6rjhE8qQw/3vXbabcDSU4myf3m
EXbGMbo7ivPpTqVzIv49MR0HQ5X3wPKm3XiDvU5GIRAIN3dwERdXg1JWEw54/mGO
hcRCFM2tkTb9mw+MoeQfpncptFlSX6nAd9XFn39o1U+tNFGP32Gd48NtW4VCoMgr
Fnx6DGEnUDhB/9xW1y5i60s0Oi/FTZQ5RLF3yUZgyuEjWGUT6QwpwulNn/7Fzceg
1Wg8BtQQwzeJ7U62Hhg/+eIHaTDX9I4Y2Y240WBHYJIW6HtcGacR11rlNbyxu+3m
fNS4It36lXIBM074DKN3zkrEnFwI/H3KCzSJpkHMWsODIusZ2+hb0Jnl6eLeIbjQ
PIV7PRHrX7fPgpNDS1+Hmozvv3SojEb9vaFDg0eRK7zOMyM3OwOF7Z6LRMG18+jF
FT6leoDvOzkbJomqHehSOZVyAMo1a02IVYVHAdpz9Vfh/Pq/GZ/9HXpE/fv+KGmU
uTaNA0oAG6plfcoIV0Lvy6TWk58E46/NydcCCeAYLqUwloyPLyVr/AIRrwh1kI6d
L7ZnSyuSMmI/CugketoXgzaFLKU8dlUSZY8J3a4UA683mL7Jcsd6Q5INY2ywHnSH
jFwMTdvEAorgjLFlMnJpfIELUEM6G5Dl5s9/zynckF2rJCu5Wh0YJ1az+GjimDba
cpfaN8G9Iad8kgYcOd89+h33TNkwGzYtk51aRrZ9TQlSCZQUXiJv67OuKZa3nBk3
uDPCVQLK5izJjHZLaAtzs9QXQsz0MF84VlSn9n9C4KRRVztF9kOc5cjkrAYQbsck
sBlqm29GqgSS/cXbwXAZHYp99O6EsVuSVrmsMIdzcmsCRb2WI8b9iVihsX89Gr+f
OfUWnywTJShUdz9BVCXVaGCjAqt5UXhlll945UQv3/zw4y+WiBQosCG9Oqr8g7IF
EH2+K2miKssdsgifCr7ite/3ziikbTrZtYjLei0KvZ5VnZROmp+wUFbnKNSwguzQ
5Z2sbZWbRCwmlYw4Wr/ad+U3Rwx2VA8AP3kumDTAuYeGhJlzUYTMzC5skTnVePpC
2DPrNyzGYMeL7agkDxPr8JONlz8Ac580rGK9CTm9oYwZJU3wX18zMvATFdbuwxzy
BdgoCnoCxa/wHQB6tqebNuC3Dpm2z9ds7HIgJTsfeo+Rld4zuSQRHA9eOtkID2yK
WIUf739K33+5cht4k4sYgHgv45xDc/uPx4JG36zI4jsqbT6b4tFF7DXPao+iN7ZB
LpQDhoDstif8fLASiqY9nioqRuGC86tttd+gTBAgtY/7uiF2yodxwHCk6jLtvP24
IWNJ6vN9KHKm5yOnhK/pAy83er6UJVHCeTWDEzzfuJPJhXwSpQaESNzJv9xsU2jq
DkB9nCPBtwaE5RzMZpOTxzJbDREQ6FERTqNZ3UuuXNy6xdztHcMFsi77HGDcF+Yd
2/4YkEVVJjRD37NXs6aUKkYLkMD4UhNURdzd0zSBrNX3H8XtBzLZnZBG3z85eRqn
W7t0InCeezTDPVfSsw7sXR6qvZIWNPrdYOqI6/MghFTij448PkcNKi6cmBLY0q8G
EWdyQ7ZxRfEsvIZQJO0Dc3k/YvJvJ5ASFA8H7cmFutcGMqRdWmzEUIHwXsIs0lGh
P4I7J9Izo8sgrWX+qsE6HCA+bxSTZFS/lrr5l6JlUFkiWv1NSqq4Ofz+65q0y/x3
ZP5MddPL3jWk2DlUdY7gNe/xMrU4usOErVEfQ0KU0X/uN9nViPB+/xhGOaNPfB41
j1kQLB1KflShRGy82kjHDq6VhJO+KPTkvwE6W+OgMn0YIJX7z3z7fu1xhd3ZdhGz
4etRomCrk7MtpMwNVs21I4VCV36Jk+9Q3dO3C129T8GpjhtpgkYrJxzGabIvy40Y
v44yigd3jtpEDwNeyDoxveIncQ+/NDwW24qaXkmjQuIPQ0YBwUDi1x7nzh7+wNbv
giv2kz90by37PEJYTWCG+frLQRiA8Nqg/FhFXUWyMBfsWMcTiBRNe9KlYMFPUzg3
6R68sDD9pveT6QlwBn4a3Obi2M0voU56M9XqljQ4Krq5JMAH19QyJUituJEa9cwO
LNXkuPK+NC2UVypWI9TsYrJcPpMKRhehcjA81a7TaaW0vaoIo6Hi6ozN8DD8kWK2
I1/h9NxMJqv4GUD3X3fB678MUx82NDLZSeqHsZF3ppZ11E/PdrlDR7Ikfgn+QG+6
XLS+YnhmaA6K2PZT2BIIRw/VEJiU3/ubKC6R2ThdmIWmHL35IBdD3TLaikWELRz6
QwFcErrZ3P3l1KBjitBbxHgqCjPHRQJ6HuJK534FQ/wKS66FLUKObAlPntb2qtk+
Myobu+/Hu11y3k6ZQjbkP1cNpi8b1GI8o4rXP3DZyLaipge76Z16knAhbwsOAyWS
RcHtkf3Z7G1ZoGAoA8RAyoavGM8kB4guGi0p7xpk1cgCsSfu8B3cHtnYzgXnLFsK
lG2z1bmocTjqsEZTvP8ii5ZHSyUpl2tNBglYg0Q3rcfFelV6iidvUFyBfCQsKOVc
BAmKSOFFCBzGofVUfb5MYPNYn19jmbySLp6Oqw/LZhVzgsML3gi3YrNO1lFMMEJ9
+A3xH4/FYojn5Pl1kaafKrXm4Sq8b1HoQBNpls6JTVP12bvJicsKjzANy42a/MNv
mivImR/pDxPGQLClJ9x1aAFxFURWNurphzEN9pCOQwYmUZ7bzMUWUX552jhZFluE
Ftwynv6d0Uw2x3pnJyKirvp+i3ypYdQqog05DVQpkmdYWknpKM1NyUbQmMesQp0M
jn5HU9EzdaqjPrIu0GkYJHUkvTYNR0ibtqWolF86GUCtC68IICWdrvPQ0wBkQZfM
gTfPXIBGdG6JHstuzeFTZeadgdrAjw4McXmMCp8cXM1UPY99oqlw2XjaywYzvI4M
kWo4siUmZ5R1E2Gl4p0Ib3hhwa9tYKQ4lQ25GKwu8dlQ11GQdcT9pJx8K3BiuQa1
kQxB2hrU1E738996I1jmu2klMPo1ZUUmdLP08GqcBfimXN7mx5l8kReAjJM62DrV
3DFeCflU4nQgDpsa2PeWn77JFjeVc2/BHORS+oeLn2bw79NBkXYhVeQuTSYmm9mD
MOVD2riowvuXTnQNJCUHhSXMsG9osOyQYy/8gZ7G4+ZnmQfZAeGbHmH3KC02FVAP
1s2tgf2p0u1q7a+V+yqumoNME2iN5bk7GKyDCoIS/hXtoyTDdB2OS8HCZw/eguyc
0Vqe1jWpondgHGjCQWMU9rIBlrFjafkFkv6YxRk78eDQsZoayO4AasYHEzZisRWm
md3jPvRs3Vxe9E0XgD61U/xMUjLrJeL4OutM+mDymjpndXdC5MfP3D9zQm/ewGf9
7zwODy9BZPLVjWgq7BMgaQeyoy4b7bXz70U+5YDJCm8k4fyDX0BnD0X8Jajl3o7h
V0kD3K2rAZZ5G5laNy1FsV2Ufu9vEtSHgJVM2OO/kNSmLL33EcbAm7EN6ALBl+QU
EXXgXFf9BlWfvcIbWh+vBN8DJg1Oj7Sjp3NlO+FCyBYNaK838939V5YkgCmPiv1C
JSSuTz0iMmz5Fao/3+10H9Ht183ngs4DjqgHT+TRokyIoZ5RO+tnnVVYN8lQaOaC
Rb5l+kEHOpYshnfN6p3MDkDhscjTL6Ba/dVvgS8ENeg6tEyHSWL374HztYu3q/3J
X7NyrmfXOrRvh3A+8NFZvgiSnHZts4M6GybF7BEYTM+l+cJzf91zu/PJqbEuFg0d
Or2yunMUEW6VRZX+wSgD2K6U09smGdVV/X1wGzL0qjQ+01vY2X3S/tyqtEr8y3jM
NpIWB76Gm2W2hDnjv3/tujdqJ+/KZw8Bx38dQ2aNFI03X8kGug3NYWPjQ6s83IF4
WZjpJ6/Tgj/gUvhs/+B3M6EoQ3iuHuO0zz5Cm8FNikiQ6KIhIhXC1w9VVi3ywEiJ
0PetjXl1iFlo41ponuCsHNLEt6eDq9Qv+aoH7Xk5SQ1xTlLnT90aGzhVBDC7cNIb
huJdEK1BwGUBJnH4USqBTCmkrl/fn8V3ZukiXLtdEv1NhvcvaquxBAfM4jXqf1Ju
ExJsNLvqPuSn2TO2PpvFnkZ+h7ZxDWRgPgRWovBQ+AhlY1wiI0nBomuKWLZWj8DF
wROW5r0JNj1ArNHYVCp9Pku6DAo/vBTtFFB3L9lwLyYD3lsE/ply6gBxKDydObr3
GU2WA+H6TUSb1zUDeQ5mEmyGFXAHzRPTPJB8aavFivjfRS5tV4eVHKf3lnHeJeht
iP++sS4ntFAk8X8H+AUYdaYUD6lH5u7c6NRIHIBVRkXoLIQoDQi5XzWS5KFcUvkF
vnBYaEE60YuOlM4LdNJ+CdZYApTOeZ/wzWsirsJQW/6he9RZMdamLfgCclAjOHdj
kpPlg5EsqB+QOhP2l7HRrNah8uHMGpisRhSc31EhhdAbptn6zFOs3M1/lXgVjkay
3WkO3x08Pf5V/zRlp3Zjp3dbpXQwHajzcXTgXrlmwylla/RPyQ5BK7EaHAIbgR+q
k71vyTNvgtL/mUnvgOlIMZppbqN0c9faYNCxtwRE3QiOrppYY2vfvFCOJM78jO1w
3S8pAGgG107bW9cX0At1X4BhMYfJR1UWVHd4Nd0oUK2zkfecQ3hd0NNieVjS66XM
KCWeLiBEk28rUhyQWcmtJD1tSLx3kGdS21wYaiOXKoT3ZNa5wdLOsTplNWOT9C76
AVrJeDv8CgnN50HNLEQV66+ZOc2CJxXUS84XdCqCV1UpdauOqqKsO+yCF30vzDWB
BODezN1Whu1WRhLdDVDGIWYVkcsgw0Jc+ymI7EHbmWIvCBz30pTJ91VsKF3QIqFO
5Uw2Nd/uBH4nV1aq6q4VQvzCNVtG2GMOCiiVWCIVppFOFWi1IAuQP3nea22GYAAo
59+ecxNN97NhDdZTQ1IveMu2I7aG32H825Mc5zZG3/jv57hRd4/pOkJsR78ETfnz
l7n4BcVysq87wwuJiLzvTYpQYuRfT5UgbX9gDdaPMab+J75emMiYD3CMx14sWrTW
nwzeYOCMc0fedWC6QTWv07dWlu8T/8NNaIWhyI6RCm5746ObgiBzHpgb0fucsX+7
6qb0JkAU+xyJZEMSrlnLkpxo0jdJaaMHKvQ74nQ8S3ZiTmT8Q4wn2jJVMQ30ffMY
DcXQtjf2rwwkFGWBTcrr4179ool769F2l/XxwOsIW6sYz31G1SahrdBpLnjY/Vre
KSJn9kXI7RZbUGSkthGdC6TxAJhq6n8P92V4ibd9AwDq1jeh9eDGLG4ZEKORTM88
6ICjfFhtZk/HJ9EjrtYuMe0ePCjLlQRkyBfIs+1EF/yk3N4MmvXsD1/yA2aSsyoS
D0lpkBBNtfBweartLeUK7N1FTxy0+FmXV4p0Mu/USUPXL7zy5/LwvO42GyokfE/x
nqfmKPrn/ugU16yCLqgDMvislYBp0OauVqKYjOA2cvNgoKlU9egu+pWwQCloxJ8H
g9CE9JsLHI5SKl4roeL5kEStNI6EE/Xpf28h0RJvArehjcGs7vD+CFJjGYcYMeJq
izdDPgd5w458Ng+Cscc50ViW+QnVD3Ea5nwNUWWE2ZNq3xULP/2VaoFT+aNsOltM
1W9bZxo/6jf1iSvqo4f6SG4NPesLZpMqn/if5nbXeyp57ysQg7e3RTtU86N+i6rq
vZNNO/h1o79CsUJUabO9ZEheEi1/JsLbHMAXI8wkVul4QJ5mEb+bRh2uOnQeCMU2
vHPoNKKxJWn1THULyNRh5tmvNfOE8jHUnMmCUAxjVBPxZ0GNim1LFo/TqvZHtlxB
CWyh0tDT2oT8peKzLFe20egn7u6qm7pGvgCl7HM+XoJJn+WcRajpg7KDbiwPDcHL
FHsOAkUfXsef8oJYkiYePtoIAh5I8I5hBAlYYTLEIq201y7ADBXU0oK7XVzeHI6g
fgBcupZTnI6D1ba1NBPdO5oscNTS95oSl+FPktra52MzhpMDu8ochcqqBAxYcQOm
4SHWxe4ObkcjIXmyFAa8nz2LjFhEqTRMbr9z5d1fQaugDJs9cqzcV50Xk6jUCiOT
B5LFHJnq9nddjOasHOrdWdxXJ5hGBR99CJQgxaiKLKG3VbDuSKoDjggpt9pXCbNr
dH5ePjaspE7xCiCjBnMKN0SmWnwjru8Pl13UdoKp2g4xjHVtWEk6ZkL2Ree59ian
FNKHfZWrXQvMsLZveKTMsZKcon/ifXn+YW5IFf0LIkP7NetXFQSsKjEqqOvFvq40
VwSNenfgCexJ6pXslp0TSLiBOXFx9QAyLAoDv/16zBU92tFNPYiRU775jHFXTk/I
LIJVnxJnvEezJXjv6oT5LFiEuEgKWIEoz1EHxbBXWK7Hls/6SIxj/nrkkDpNl+oW
xaaDR/LoBTAVvPMTl8IitCniEg+ChajF37OgpW9mHOa8TRxUFBwSjr4pK6vB1IAX
limD5MR2J5rops6yF/echww9APl9BWADlKYPrudQpgArMGZdc0oIB28Dt9OGam9O
1rwAgQl5Yf6EG40RMTUe+if5s/lvF+1cyewtgk9Qdw5ZjZz9LAcKeNjbZ+Acuous
/gEEtvFLeBlRBZ8gAOon9VrlgNeGvgDKkEYIhOO6eUyc3c4US24n59+BpszMZfNW
7911rqj/fwF/VXY9mqIvnLDXLQlt8rQijT/xVyUwnkWAQAzPmoqNSImMxBBcoTlw
dGhIsh/rCvRq81XE9NJu3HeuNA1cg5mRwEZwIDVxgIdbBmlPqCNye2kArJfgK9Sl
+Y9MzCsdaBYkGl1Sn3b6QYyP1T9TynTpSO2Faae/OfqbNnBOIKPWGBW7F0MR/tjW
MNcqlk0c2r3jmNVSMmYezBN9jqy0eDDJzVmauz2+l1QX9JRyswU0DUjoOfL3u5Uy
XdL7thHOaUbCn6ubPUpa99vDeVFfNt1yZZeaTUQJI4Ww673QEozZoKORme7g20WX
0r27e7XF37UV63AfsSY5VuauLNfsxAsvxJ0Qe0Ce1EHfB2g2DWlap0ghiJkiGhHC
j9YK1aLVmarMRvIS7n+yZa5zgPnzQ0YncIvKpZohlM+SbVSvLFJ8h/X0FF67CSsE
ycZyCEJY9WLSqpIaerBZax0MxLBNvrQNjdVxuTwzPySVLcPOCrB0o3sNhyIE3fo/
e0zpEOnIDr1oyW2WC5a2Of3CZ9fnAeTt6HvveSGs2nr1KuR1L2/TYDAtJ98iNCCB
eLT35TsP2p+rZsLIAvUOkEfELtQUsa5f/MkU70VUrxOPewUDu69gbCcdnMDsGams
8ge9AHh0iqKOK6fSJUemiOiheh2fdvaM9M7/qOyoCGnx/znoI6hcslDbRvkqLmrE
dLll6CunFl2qH9svqHFaFBcEU6/OfJsZ6Hy4+8Mj5DAHjDl7rlaQYneBypAVZZWT
TmkvoS/c/VOfQOPWfxh1oKaDXSfzNKxP9jjTRMeSWUm+XjsS8H0ZYV7herQw3gPJ
z5XU7Ozg98i2qYfGBqWVCQDJ1EDUFDp0NRgZynMeQsGwCA8jr9fv06rHGsglFhcS
9QuiZXe8rMjoNY1FNRsmmmTGlsodWLkLmJV7WCNp1YhNaV984SvIZtFL/JdJjrj6
i4hoiP0EJSGR4euf/H5ZrzJK68vxGovdlU40Cj6QFTqDh2jgzbroQjvD2+9SPSA/
KW9c07i9I1B8xbyVBhuiHF5NfuLyujNjJbflsUNs9HCYQVTeTnZ/vzY/zTnm3OLM
JYcsSQEJCTFHiX+BPYcM9+mWZTOiWV012QRrNrRDXOoIPDLBcaM8tInzZj00nlHc
sfrS59UIIWmWXLUuWKdW7uOYGbpGMQrH0hKBggP0OpAQE8qiU5/aRr4jQcmU0gPq
UVrgPu8zW3Nx63dpZMLmAbmNIYenjE2QZ3h/43223unjWI6XZ0jT1obW59KPYQdP
5d4EoZO99bTuoryu41sC66Sx0+NHC0b8k2/yzPghn1d0iFUQNxAJX/Y1JRaXKRIT
LKjFy6OSjeeXtOrx+Cmhq87oQ9NJpDbHjlaQtVirBO96IGEi8ZNJMgxQBdM0jYSW
SmZ3dtDZgqmMT1K2kJwr1FaCMX4EMa9U63ALJmyLA56l/w7M37wpmJ6XicttAx86
S5mjowZtH+U1SS69Vzstg2DfXJxrBidb+bHAWHSFS6wPlHSeVL1vG8lRJoQGP3by
leU6eDzkSnyP3JA0wwb2C49mxYwqNHlO+vsneaWwGW5I+cv62h3Al0izY+x5IJ3r
RAE5pMAmWk+VPBF0IHbsBKjbj8E4zbL6RxOhAoAfFPidYK2RzN4Xz3Cn911EDMXb
VRWE/ChNlLiOzXhzpnEOtZewk4/L/za5Q5FN/62BIIQAU2CHhqSHO1MtsWmFSb3Q
vvKWTfycGoHrs6ua9E+fwjLXA6i2VwqzS9tX2izFshsHoQVemiHVg7GRRuAzrulB
H3oOBlpN2uWyyuD0y+tWuciIb99tXBYBI+PNli387F4/FzE3kY7FMTpJjoHtnPZL
pm8ndLfGFli5VbUQNeOGWugVKRSim2PBfkONzk0/LcZg7Lg4j5Yu8EnfC2BEwT2R
CcE23iNnUgnM2K+q/GCD5fb/xZbFWkuky6ulRZrLL+RVw9easaZqtSXYxnf69kH2
Ly3RFvsrsELUea6+79PJf+4e/YKNIfnTyCsIGlF4Zxdgl4pkTXsMjOjxIoz5XqhQ
uETiEx5NCpnaPcurtw+cvHgpccDPoQrkByUARj/uSPrSQ1ywjIcZm/irkRXdwNEb
3enwptG18BnbihLEBAxeaCdILDc6q+0DM+DVaA0/asI+G4fMf0yD02OCUQhL6fMb
utj4/pPpCMVmT08qlLKhBSeqG3zNM9H1N0TpEZDKsz87rX/BIzL8Qjdh+pi1dgf+
Jx8l7ZXldAwGJQsMWS6jHqBPAA1S3secYYarJm2wYvmz1qR1guQ3MA8dv4XOEVJv
kXgOxTCgXPGfwcRCdao9rVvycfvf+jZ41OUiwqboyGONJ+yFcYHDSvwzDTPWoBMB
ENsoz62c0ifs3RaikexI6o26noD8aMKK4lIMEHofLdivDfeQU2tz1RtJ5rWalOul
cdZmzeooNubTndJcA/esMxJQqYrADTW+OIolOqP9V8eAhpymbceo+0AGcqjqgwH6
xfaPm/XOAh1asTQkwW9GifQtnEl6l4yJ4hqlI/nm8JEfxVDfRH8QMR7UYsBE0E8Q
XabYlc65krrPRu+vWSNjUf66rtwY+qaIqnchUPyj/T8+bSgJO3yhSFiZGqMjQRRm
VRR1WIqcJtOYbQLdDAi880bN95UlUjdVScVUuRX4hdQVV9P7+a6bAAuIZKuprXQj
SM/EL4Wc8YmM0Nbr29s67cC5Nn/33pJ/thl5W7GLq0MKcCUugLF9P+qcEeuw8nVc
BevTB8ULsyS+jSJdBESTFtt8bDRhCgfJLf7XLmCaoBLO5NVYCdMtgy3F+0rGJq29
8A6ZxPHVqi5AEJEYBPVa3gIj+4CF0ctTitLdpReZfK3JBGsk9oovqC+1hkDi6BW9
seXUbAuNG23zgRK4EFf/SYtwhfvLe1v0IJn25AjK6sJyL1DmBR6N4e0WQHd4sgaG
DOa1gbgntJNYIUG5vStXCFOIwR/oAwr/6R/FExig5QkBYpAPJmTtPgR7b50ZgnPH
UMhYWPtlHDhe7Wkkg7tOOXUo4mRe8XDL5uEGVnEJDUdYqsWfBNwOfRfCfgF9nqGu
ihrOn+1+UtOh66YVyWgI8Xp3xh1vLVKrC52DfdRpvT0ryt257hItFSsZJE4HXkWu
gZY0qdCOyTF6wkQBiNJCvkpa1Y8uzgOs9DH0Jn2jf2HEmOiyNtSRDLe+GAk9GTdz
KyJAx4+V0W0iHDXfaLEOeepzr01TC3b8ZcsZQFybPCCC2dzA3UIIKLUYrkzUI4CZ
b/1/kpbE8urAXZ6WF39LbhUt62cDTMUjKHFHgyRJlVD5r/BFkNujeVpnkAoMRk6T
jZgsW9nSZZX7DKsFVEyKVuGaXK0zhvuDRhHzLIDgP5tfH8BXn8ssK8czsS4nPcl/
LKG4Omy1n5HkCo9WVHocL0K+sHo3YslHV0PagKvGK+HYxt87vzRcPj9gHRJ+5Bp6
H+t8thSq/y9OC7Pdy8CsA6F/kH8FfSQLR94d22C9L8jtI38lEk0vg5N6+EsHrR8v
5Ldre0ZjAjTrg2L0lxnMuTcEW7qtj3rrifjHDwJJAfsWCUwwC+JECA/VbvOYS+AY
KuClRXXztFZfb9x6hmsxv5nbw6rnQaz4Yt8/6xPqU+V6SamH52mErCz25WK3c48R
g1Tbsd8teZt+l5PreNavQN+7DXhgwDt4avJT2zxAh0Dp8oOJ39B8vMrqJ3Vvgikk
O9FvGG7Y4usedHb+DWYMut9XufoQnaPkkmQBZD/y1G3Oa3xLHSxvDJICTA+CIBzK
dU124DVus9kW9icyER2+wriRbyyVA+a1P4pHVHY7iB08v+8sSJTNTcMBW6UZKzZ6
zYoaxSzuZ37rtuhNpyQcrUXBy16Flj2NrejygtDKNUszZee7jcAdMAdXAQ/vn7nI
W5Ih3yEhkgIvar5CTtOwMQ0Vfw357DYDzOLj+wnv5iKJTwOEXcpI4CYSfUyrB5MU
k3Po4hI2hWipeIeGreVEp1z7Z2XqSMslK8q34idxT09HHAk30CpvvvzVEqQZvNpZ
IchOAptjebz8oAlUQ0M/MYU8dubalptnh1+1+y/I45Nm6rvWIMoguRau+4GzD1Vv
KwdglApwM8KFifRRyQ6AaIYgWVtVYADxBN3pbNfQDqtwcMnRUL5pdPOmH8Z8/o7N
4dL1HhjTk7pLosCYmFv2CrRpPP5T5j7bBCNs0JR+dcq31r+XIjmcs+d07oN1z30r
YHhBYidTBxSNBV+xz4du/nNYVOeQwCgazice6JbzN7QpJbWljQEwi7THHGCI7rQ1
2fon4szSycWNTLMC5YCptKc12JWcB7gf/uYCWLDRoDRDmY4sERDoIoMrlB6f3657
A2SDBxVA1KLIfPpywXl5wRNrmNxxWsJQQRjMeNq1eBhJaZeNNSnSfZtqva1xxY9s
DrK6cBs9prLJEP5g8G3SL5UX+TqFjiC/xEkywL5rbOCm2EZoL1XPe3OYEZKUZF+K
q4pe1NqkcivUko9SLmA45/0U3TzyvE9WqVajH/HN1+UE/yuRgPzicinlfVRCH+oa
jKj7W+GxGWg9/Tk/CqN69qYKUsnLsDPM1lc97xzDIOP2Mko/cuSZs9wWEep5t+Ok
DBxTYsu3EaPJMDwdZeVJgP+wisCB1py4IL8O7l/1ZWM7g0052jatjCsApFduXKLC
szoKHKVyNruTUSQVTvkg2fBGENX6GRAijf+cefbekDcseqen9bMuJqbBURqc6sIj
9QToZlXGbXZr6enX3jkqaoBigxPl84NTHPYXKIypef47i6ALxzS3pi5vHNpyDyJA
vIWqrIE9/YLW//lyjWOWnrmZoKZzp4k6N/qPxggvg5Y8dtxd/nxpm5t7AG4lWnea
yyiICIVHHjl/Kfgmh6dEIwxu4mb5eSzKFC9FGe88kIyza4kf1RekF+VLcWSGFtJ+
8B8VRLsQZVYRtywC6rpUY5qArY7EA59SBHJHT49uyfkQRyHJaQ1PnDd3rc0m85nT
o+39a7nKYGUXful99kHsC8Y2srBSmpbDndmjpOSvNi16GTOWnKWeE57ywTyQsq9J
uRXQ2ROiNXlcRvt+FFDz+SZxyzN2sIlnD1M4wSZuw6e97Ngpzh271v+pPdTJqVc6
WBOHvIrRodVsmZ+qCqftBPCLboGrOJzAb78ATEaOjNjUO/lpdmQG8Yv/AOZEz5C1
jKRbcz9vvC5jxq7EK/V9S+e8HfYSOS+kkMnWBZtF4nqaH8bBrKG95hgr2d3nFRO2
zY53Hc3Ix5oNoGcbl568UL+xsTpjWIFjnhlY1j0Ac/4vf9hqLtSeB5J1cGxXNpes
JddaPguadWhhqSS4E/nBGPn1hHsYm/nceyvwhZ8pmAxrwjZEPic/lSEhAZi5eocu
bQxZHpCPQh+Sj03+DPLCI/n18l/Cl7eblOp2Dlz4ip1VKSzX08ULUMJ91bA/VUz8
EHOCk8xqjX2stvRjyP8fZtL2qbz1qayIJTR8Ymw5U7arJFENfywVL0wguU6JHyBM
TUo/P2YGaAGeT3M34ZRy2fCkdPHk6s7skTw9P/jZCz+JamUE7/tGmeQznBj7Sf9K
Yx0b7maRCpa+6r8vH3uiQIcWPLR416F3ldcDSgVHzlquh2SNll+76pcj2WYLbeQd
TmIqk5uZeS/e+G+axiXURONFKod9pkgcEqiKLaq5OCknvrmSgSLWcD1pVTYtZtZz
VlsphzIO08Ue8SbrHY70hiVPRsUdT+EOdph31CasoNDDFOPsN9bbPZfW1VkmRAot
NPpjGr5ya5p42xDLnrvtt+7WIn0MLWUiO6lwDs72ouhxcVKLQzRgjEVg+ldTl1/d
Mr/dI7FOUtxykoUm2Lq582cB28YNp+4wlLVuk4uBWOs+Y/ObmtZ+oR/FgpQDewa7
rODZaSdTVRJZju0iEk/EqhZLcWYZPbtBR6goba+XfZ5HfBV3JiwtsP0Tq9dsk5K8
DKiqQg2kx3/AU4zAEGJ3hvBg/hz8rDu08pJOkHeOAab/tlVWcRmwgH1UWetm4aly
H8V61DneezrJOV2YIRJVgnWCjCGvVWxcNoMFSZ2jMJ4ToFu8VQ7BebyxOF1GB9Ss
mGdVUoaJKqWVDk8efA75NxKbzX/Q6Tf9uUQDVpLjXu/hYhlpGlZvnhvWFWt4QsEP
rKjQG5mR9eFyvZx6do5g5seBcF8CFHTjQE0w7G9FaROFZ653Q9x78hj/IbKZcUA/
MlzWRvZOx6B0rrEVnZXEtPj9FduvCaWZbGXS1Gbeu9DYEP+Cwf+wk36Jwz/dNfqe
dMyxwVlh9rOK98xiD9hdUntyHApRGy2rhovNvdkfUI4Mf4Kuobfqkr2RhpnUN721
BX0njJFDhb0BKZZXI7/ACco7NeBWF0xYpqxG0a/VF5emufgS0/scNN8bjHLqr0UL
WSPHhlyDC+aODj3EMlY4OHxqV6f9IfgvsyuFyszVS4lwtgyIVlOyTyQuvobma6Gh
P6SJ+Lvl1j0gRYS1WLTow6/KvybPwj1+ikE6wehB7CkrOmaA3gLEH7gcE33zUwCp
C9hTGSC8nqPWJ3+7SjXHZgbs/gTmSSQ/u2f5aA4hMtVpcFIVz5xaWfnM/eWECRxL
7M3AkdltDrrEknp15ypwFqzs+qhBHTwr2SMT3W2jDzSuHb/eVD62Gkx+8fiV4Epw
RWGtE+i1no2K3Evs419xLMFhJjf/mjX0qNPnxkIgqLNtOQTXdiGPtA2UcVFVIi13
fH5sTDDOre5u/3syE/n4HlmPKyZWxYMCfIz09OuOSQUn7Ae3WbzqRGCyaf5+iBWh
WnT+dHoaHE1MMAyX33ynshxp9hgOh9TXb+/qH3sdlfQtc/OVnS0eoheY2F31jTvz
8HXQuLlUj6oowlDpniimqrHY6LQrGR1AlufcNJuH3/nT4Kv7Ko0T4woxlqtQXWZX
3VdcKhSYIRVx7BnLRi/acStWErf0VoBESVTU7Ocm4UmOUwJ6W3KoWsPWAM54MqF4
80GcdYuig/hzTv0D2aHb6hBxMEmQwZ81DezQ7/qTdbZpglN++PqS4y5Yk7+V7gNR
ajkvcT9c/Okpv2auF/YrpF1xZ0Mithy105J013y9uoSSaQUPPDbIwYh0SLCWRJUh
S+geRYr23xRKocMrvvZbHDFuINqJszH42OcWNTa4RiAQEoRRBVrLGR4k46y03KLY
XgtPNHTickRR5jqE3wPCIlLYDQoiEa0WPDfEKYs+/j5IYp2QXCUahSh6gYy3NBlD
38oZHyn4cr0ktAc3emRY152+vc6kGwKc237JxeRivpgVFjLttFuozOzaRY9WRAB2
gnLQCRzUC2MSk5fGU0W2oC7GJnLdK0L3LbIJmpqJjBjOr3HCNTLsRzUvp2szyLMu
LSljoIWTj3+i7keYbU0D2mWRWbwUPqiiV8wjwpJFyftLAIpdmrAQ07TCUZvkrW0T
I8QZaia/0U73YZJ1ADZkJC+Nqf0atq626RQDugM/oZ3Vgyyv5T9+EsAJ+ZtR1TxK
L+n7AQ3A59LCZk5QhENU62t9Pl/A8IVrhOlMBv5T4bCGVFBDmr/TyIPbde9Tr5sp
V73HBS7ZDOiKBNM2sI00tK0k/simJz2Byk1s5X6fkMFTRRfTyK7+0syh/uSIaJWM
lrcKw+6GpbzAfqCW+SnYLqae9tlZol2YttcXq5h20tbkQjK48czrIKLllSf6IVMB
lKe+T3dNRpylygurn7BQT/uM7J+IGoj0VfzDCLCXwIeCQBdTe5/RW9yblk2K8j+g
S0R+XONWx4F4i843JlX9vpWzaZewx57m4gWcjOUVxjVGMyH8k4P8IHN8IP1qLQDG
wbz/3yciNJwkCyoANZv7gj+QG/UcvN7dUmzwgflynjpKLsp1byf0yhKRQTJCPBXJ
n8/X6Qud3OqjZoP3YKhs+DJ3WLmWNPOKFMJCF41h/I7NEBUADTwTUAcRZt7OQ43y
dYPOhQbFC8EBFpqgdLyQiKiz6FcxaVjWiW54LYYEm4UucvO+4JXAGr7SKQ8CBjR4
M9UL8Hd8qpDGtRrmtOJwUctU6KBz3gGBS5pBN5O9KAR8ffPjL66ag0nQRv/F88un
j1tCVTFI4zWGeoEVEhK2ZzGNtV4cOWiHUOywm6glZpw1zamGbeQ6MKvy0osqp32Z
y1ipmT0NNFzSSMe8MqRcI4UNNrvkMkyjsEGtE3ASmpoTgBaTVlXOILT/Y/e4gQZ/
tai9nknp1iEVUTakzGdWEnd7NaZz+BqNwIRRTaFCHndqcywL87Nhv9bQpA6WQl2k
uRHOZtNtiELAsIm8ayFPfLgH1f3xnYPaa5W6wC5BgRaAzaZb5JLSRUbw+i/cpmnJ
LPw+P0x9c3DijYbadMdgXTG2wEjuWKBiJEwonmjIzVvqjNQm64gYt7EEgU2Ze/16
yHO1IokQKV/FerAxF7JV9vbmwpiz2Ti0caZxFhGny6KFskr14JPj0nTmv8SHBZ80
BpVPt6KyOC9ZTVJ1W6ceLOK/C4yyDWbLi9D6T8h/SWX/2UtaSl8l26hb29ZhZqEe
Rs0tMUGrLVP1bajLwIhUKI1G73NyNqq3RZafT0TiYduL3CeV64v/v0CapghgXJsk
+xhm/ojl6WXo0QBTDP7U2Trsk/Relr1LxNXUAMfMpM4v7UwheM75oyPP14qzPqcB
B0AJR5Kkwxm8FfGkZYpyjRe/rVxMHtddoGjzYshThEtEvW+QRPV1UwhZd53A+7KE
Iak3TUUm14gI1ZYpx9mV55WOQeRj+EnaF8ZjNygEJuVacb6vxwbIXSJOC+dMYUtW
LJpLjEjyEPxthWFEXimyoouQ+jFvQZLV7D93+q3Gf8G0mXVdRUGADHLzPuSk/IrX
0Trkf+caKN0zJCW+wDAIYnhQNU5VqpCDQgqsPldgSUu7PeRrZTaAjGpR6GrbD2DJ
bv3zR381m7wxDntmLSYVOtJg7ziBtW5JBkNn8L4vyhTyKT2okNO0ANNdmFTghvnf
QchCjWYt4mj2YgC2CuJ2hWWGlnZw11Ip/eZOXt1ZZORD3LeCuQO53lr2NZfsgdGH
XKnYxpel2enRFGdSLnf2lwg+tl7QkZc0IJF80R8iFxmiGQ6Xt9MPHV/jVw1vYgDw
XFyOs3JdqBuvA3f7m0hC21NCi7z0aB4wNBFX8O0e0VCp9V5P2fnmeISpPcuyD/7J
eAXAte/Ze9tiMvmPHXC0supTWBjVmywPbQtvoKPCJ6gTRBLESQhkGa9LUIjHTzO2
LcNywpw5ZBrk2hV8hAYhTXEPoNpHGj2BxQBpJ8GM8AjvZiHMde1/wEI0htY4dFMQ
FyodG/5lPLvurzPwfZhya/xzgY7ogxVOedbPQgHuddcSbXaX+aeYzwuj7F1oDfCJ
sJgk0UaP5iDqKD8ZMlGXzObqe01sldr80ujYfa4t5xPsIkeB3m9Uyjo5tNvMgGJd
kf4avBRCVpsab5c8wM73p3DqmVX7JyvFy2MCU+RlZpoH9mRfRK5506E5gQ0J04NT
uOfng0/ybO+zBz+OjVvsiJc9QLiydGSWqaLRqqfR0GoPqH/48KgoiActKCm6Gjxe
4gQMju5VbJ+QfbU3e7ycnwIcp8hRZ5ace9H115iUNDAVw9apUvzJE1/9pPb67YZN
XgA/gjSO1BoZplg2qvwu12EDSwgGmzBbZiED5UEBYBWz5L/IIZkX1UdrKgiXZdJz
WiyK9qHayA0pmoEO99YDppk6juTrz386yyxST99NVTDIJr2uwwl0j4g52jLgrpPE
SU3WyLMygGIzpLL1uGlw3zZzdcUYSXcWaBY4UtVt2kBE4c8YYkHwzTiwD451itNm
t7pb2DK1Z4Ro6spEhXsH9W8o2h5HXF3Zz9cKUhKYWjAlvzGYMPbVEjJhWXd5ISm5
Kb68Mb38xU0fV7YSTE27Wrx1Qm6Rh9ozkEcDEmBlRALTHN+3gcryH+wkRM+idmzn
jD1oBtEELNLkNvOVLDBn0o+dkzs5LTV5/W/e3BtEzXkQ+3fPheVrqR0w12QsgDP4
g3UePFOKpIZKHvpZf3JECgpJnpmOBfvWGnldBfIBFFiaoWGmHh6pMPhZkDbCLdXa
Ij47TRxWtssKym1reZQhpGyhLL5ttZ2CNiC91bZS5p6uwruVEuAsUUeHg/uib150
ZOv7zNaLNcsntehpMSqeKIuVSHvvrpcfHmSWqZnFEuvYm5OSeyFD4PHIZVOVb4my
z3lMjX0+qFHH3TkqxtBQwhI2WcvE2vflnDXOeIHjxXVABNCWCqdDdpubGRWbguUf
pFmvJR2BzICw7Pz2WyY5IwP0+DMcO5ZqBuBR31dvVB6t5t5GTcapuA1PBD/Lv3l8
WBqcGurHTBTcX/dqxctYaA+xVOWeVjR8K3qT3+rOTMizNB0QL1Fe1pF86CYgVsyH
YCNZv4M49eTxYs8r5qwRiatQBodGbhtl+WBi8NO3JExRxvYC5cm8GKOMDtF3oO/N
Bxy/BoeDmIcRciNg+s/PEH4iW6uLNlPWHptzzsMNxZ+eTLPyp528rtgIbWAFFt0O
vZW2UMDXNCULjmy7YAzyxgsYbLsFlY30qU+xeXdFDrvAchCC0Ar7FFjJ2Hi6Gww5
PrX388wiD5ulZY69OFjOXcRTpJholHUhr/nVv2jMrGmp7JgLxcglQ+9XZau2/9HQ
5RUcSWID45DiYCuSQ6mDvUEce7x4fjVsVM9aXdKmrIOhE5i05712T7gzN2YYqb8D
AZwfFJ/1asFOOzOnQLR1Uyeb8AKpwfppi+IFG0b3MU9b7fM8HQyr08IDavVv1JQI
xdq0ZfgG+eonTuRkzjNymm5GHfEdgVFui7+RmHLozZs6z6p1Z/Ihlw+VJ6O4TMqp
+hUE1tUln6Y7snUYnXsRuZVvnIczaUtDtup6WW760xGK8YUqHhiRj1XoOyfo9RiU
X9qHMG1eQad1vMOPD8QBEvqAu7jLE+Nci+MtGs8Riw3rnLxzm/qf4X0CMCzXGOPB
ugYT+PEr9Ai0kg04z2zqsVn1bHgm1sh/A+Bg+KZHKFEqeMOpDtTxQJB7JiTQnOA5
o/E8FpI+2TroxSn09jACOMAAvjARi0Czze4XSoedmLoDFLBt1WeTXubhAF1+IGVa
4CveLv+WaM9MgZMvg5beF4KqIPsxy2FfKkyQ45YgyRgIxjAFNVKvkEfxoaBcdoBL
fN4ix9Wi9IJqCEH4xmLxaeEyF2WLiW2eJ2YFTYKSowvxDdoCdPDexpngsLvrIEMU
AUvDk9oCLUSBoA8m7e7GA8guDZhQB/gRBOHkq+DV16nNu/YOFnuJGUaJ6VRUBKY/
qFI3pPAgxwMgHx4fPmZ7WZVrRtcFtgbxt9Eib1sO1hpu22knWU+BWwRnlS8GZdGw
g7mvz0ZHvVBHq4JrGmbRCiHoX0xntKJP1AxvgPCkl5DFuh20hNgQ/9KSaib1Hxn4
vC9XBUY00CDxUN5ER0RGN533mdcSb1LLiGLjQKo2zti+BXJfhxs9TPrcqWBwUeVz
U3SQ/D3wu1ZnKSUQNLI0AwQb8sIFaac86/rjoK35HbZ4UUA59FcNCXvFQexln/+u
kdUyeNkixi+lqJFaFNLr2cVln7MYzWUzxnZrT/ynjDoyBLTHG0+f0TOZMw54NPtz
BR9R0EDi27656tjm3hMJZWUhUFwdjJ9rIDW8cbtGiWL4Mo2EgXRZAs1QNLYfo7Xj
lVkcgvno8FIi9zaeiYtk2nKV3efUtlZ5wRhOHETm7vnsSgLReuf0E+RNo+RWRA1s
EOOr8XC4M8aRj//+70u8v17iVOB5hTS/WVXcV9q6TkK5XlkeSZGIc3NxP8jnOR7m
I61m7EgofXD3EThYpU/w7SfJtU1+s25lIzQz+WWfPxEPVDI2GF+czVhkk2bqGgNe
trWTkZ7Zjy7Gpc9ICrhCSiJjqBfL8WWtXxsQrPsmorNAYF+HTh08nHphkQDxYHC4
K0fsIjMul/N8uFJmJ+x9ZdsMM3Zw9DfKGCkvUWBpYK/d/2zXGDdhw7GYftBSHIL3
dFJ0/GFyBtE0YAqXbR3jQahGLJZnK8StDd79CDOnxwcgqm3poblASMkVroBUdd04
Zb9WFYpQCJhJwOssIQJWqCsQLm+q+CNDAST6E5Qd2M4x/27MLVrYlU4K60CU0SYn
PPK7o04d/cVBHC4Ulg2vHVv1k4Ye1UsgEY1S3u0iZPmoQrGAfQiev20DmbTanAT8
cfS2Ry+vzaJ4tplFb82tBZnjhy071ys2Txk0/p5gsPe0Y2js52VyI5nPgJCJVpRc
pM9I/ldBpuIGOiCN+0mYYdXIyZsmyaJIgBvLR5tcuTwrkQYmiNz6MTejHoBeLorU
shPsaVI1ta9m7XIeQ9encO8gCVPWbZc+9H3wuSeIUf4KIJVZt+U921n27W9cu8H3
HjdnoN/kNktkXUQpBSYy626KmU8UB6mxImMPgArw8NcMdSaoWody/h10J27sSFgZ
sx1wkkb2K1F3c0XNrNr2LvEqpOldHKC3+fJlzIphkK7eWmtQJopAQPVJZ2qsBvm0
KQL4leDeb78JaSBPwM7mNz/q9I2kKw9PoRpMO5KeoiNpbc2HHzbKJylp7j09OgMo
u+8uBX084dhRI65bGDkJTEhl/G36eFeHOE+nAVt7ymDXBzuNLqLlWzGFFfIKt2y4
JCbnNWHXqLfj2CexM4UZ3vHa/l2mia9lgYACHcK9haFK/s3egh+RaWuf4O3RwWs5
xaQ9TZawrBwF9aCRKMGrFkIbXkddnOi0E5nD6GqQN4RNUOZtBv6QMx/fbWMbU3vD
Q3GeL0gZNZl+R1HC/R+IHtm0KlH5YQftTgF45Mh04Sy4lPc+nOSoFNScAiXICvJC
R8nIgiS1ttGFi6FlxjXmul/DMbQ8MZAC8bPg0LukX55JVS+Q6fAwYo05Mqs9IdfS
d5boQakcOznFiSzUGJ9hcTGasTZMc57ruwMp7hLgmu84zHkFENLzbR5fTNaD7hBQ
wRGMHGjGzKJS0CevkcpsLEZHn8G0vDA3HDHhRfxLCc+1Srw7eqSJ4zDPASG8LLVb
NG14HDRZXYtkQffDfGP25C0fI3vDQQIJMCc2O1/cJv0sfV7DrsbSodta8jcAa3l5
whmZE/obT2Zkn+TSg9WtqlpzbXw8q4+mA9e4tyfjgtPJZytBm9hFyDZjKnES5nCd
qiPRQkP3YpDeI5kse3RTMHavoO6JwMDP0iNWggLt/AwgGPk4x+5tkv7woHeMVN0D
JoVtyTrmQ2Zs3AUpIcPqvHlDKvcS4HsHH1WQSxX5d1sWohxeYDGxAHVR6dMPE6Mh
jcNfHHwvK+qmgmdQ81OYXafnnXSIASQBHK1BNbcG3sm5CLHuMAPimVdw9BXcdQZu
5BQ0A7uzmab7CHz2qlhiUX/YoUE+Xz4MG6tFnMxOK4NGOt3tTDDy+OaLBui9d3IK
cDDhDdAyAt3EQqR5bjedq8G2EOwbDSCdKz8WfjNdHNvG8a3obXR/GVx55YQzRt4j
LjlSoGCpNvw2ojOJOp2WpHHmtNrwH/7Gd/0pv7nXzXiXU2Xt3bHP8/CWVfamYGf1
MDuIUqR8Jep+QtBFWV8fJroHuBdcBTjhdQ1tHkRZk6DDA5WLJ7tu4VsF5Ew20C1K
L6YpEJX2PTGzGHsmLrNwzvVMADLA5Upxv3rCflzTqg7Q+B1a10h0DGZBF/q8XQux
ZuLDY4Zx6z/rXSqurHpALRMF9y1qebbicV5P3hp1o8IrPvt6PLLV2iN7XmDDCcpc
Kr6QHnFsXZhmLJJKfV3CBfsyb8HBPkWskGpW40mr/scjSd6RHBc8lB2vjM00s1Lv
wHopmIMBNcMVWpSEJnFNN8JtbrMSmIjhWhw3lviBvWUYzCrh3Z6DOFnrquojpdcC
qX1AEVQ/1MmRDLCvMLeYspY1kmF/Z2gPBj0D15AzJ+um6FdHngvRdOuFb/SGqFIR
1cb4TQSIVooQH00aBsjhimfCPKw+4isn1wMCH0cG4DTSI1V2saZxtdz9ONaarLnw
gqEWrPy5EY4bYS5ePL2sXUdbu89Pm4ETAsgG9cUhDomWyTymk4/leGD2yEQxhwYn
7fnKXPjFcL0NRxeW+6W2x/gF38AeJLY7yD2WMkEs5Br2xK0saDwC98bpSM3wNFGM
N6asd0GlhfcFTD8uae6zriYpJvk6PYrNBZkJY8/IfiVXMSUktwMp18i91E6EI0HZ
N/ooz7nVdCC1zPtXK+s/Ry88rd4UI3zDKPh1qraLGuhdqkb/w8g94S74F5xpgpXq
Q+TIkN74gQn5C/mdAhFbVPfJFyZS0RU/K371c1NNIcFl3wuDm4wDIAtNufmp4ZCR
ZGIFJxNt6x+DzKbx/4pC4UDJLMrbjXh9ABx29wW9fgTS4AF5fjp/VfcnkTT8R70k
YjViScR2eLOpChd1hdtqZQmioqueTUp/AUWJ780YwhH17juX+5TaZpbRDCgCQG4t
QByenVaVB31l6gxILxd+iKWwPV49cUguVGovR4Qpi7igsP07QfIB/ZqwIOyCZ0Mk
Gf6LPTpIc8DdMzbLaFbZIAEK3HnLr1oZnrETC+NpueKv5/B+l3dTQDjrK/0i82Ty
1lD24iW363Yh9ZArxadKQV24Ku631nqqS6FWsVk8lDUVYlOJXcwGgmoXb2gnco9O
5lwENWerUETYyYmw93xdUB9aWlsnK9eV2I1itwu1pL6UNY1m0xLfEPfXlzclHQua
Php6tCTb0AnR5pgr+Bhs8FkNjUeDDXwHbsoDsY5pKK2VODFoKfvHFiMRlT6vPGRo
aueAo4P0Q0FsjQ1nsghCGVDjUCSrnG32WJ3PcxufW2Eca6X/NfMoTff84ypWmB3r
p95uHkAq3moMCmrCdULUvbkr7HoKQk7zXaxaNPfjqbk5N7m6k1m/sEk/7D03IOBy
Xk3hrp5V/zT9gmhkJD4qluJVnp/BkwGfWjzGJXPpeX9pYzbKJhOM0XaErUsinwH/
4t4TetzenZ643d5pddQKtmsrcEmBHE1DXQuTMGFRWTvcn917N41VUFY0G24yBeg4
iFm7tPOXf8c3JdTHSVWB/zvk37QX/p31NXEgN6bSOf/QQTfIFaxsiznOHXJhULXY
Wkm+TDEzW2RDanh5wpjmF5aUcthaTDjoDcqHDq+xzBgr8S4+eD73piOWJ9Thvr+T
pegD9aLPSuq4PgWUUKzRdBs+rnaB+7ghXj/EVSwRl73Bf3/P3z1Hxmzb/Gdgftz2
KoyDpeB+mExOGjS8EsFrNtvuPGiNjqD/TbUFhlGy6MizgL/snGt4V3ronat8Ehl7
rri3+thBv/As6VwcSi3emQmyoO+wNN9FWllkXtvfQzZJMSgx2Skm8SO/wGFdeCLx
R6FKLj1ACrsDmsWifih4R0JwwMGBzgP4wjbEoYv6PUB1aALmnNKt3q4+4eMXWMRe
KpYuhrXN8VPgqjvhYHuqZrrZDN3B/2FSTlXk6PtMxbv61m8baqcBdmAc8XV0Eq5r
OypdNUlSalmQqZAsBuiK/q6X4lH4OgtbiiRp8E7BJ5KrK7XEc+wugnOKSZsV+nyH
djqwqni/1EcMRjky0k/hCBCUMZT1EIpKlgcJjyBXpEbmD9pFUIn+B3lhVr22f1ZZ
/wxdAGyShYJvvHPUE8qOKp1puZ8DlQthqgpleUeHbrh+HBeOBXPsahNmiiq5oogK
/b1Db4ToVhBIkusoZW4Mw+b4r5Wvokl8vs+89+apc+spg9ma/Nr1aCEbzQwZo5LW
JglwcfCJnEh6s1sy3Cq6nFfpPIpUCq0FnZSyDclPXj9y+Ah4r9djjRckvA+lUZ2D
jx2E7TC/jx4tUu7DZeOd7q20M6a4EQkqB7/x5WDlFtJ+IfBIrhnKr+KndbynwYdf
HTM8xr6rUde+scQKQimjd36gowfQcj1Mskqiozw0Lvui7IwzWx7x4W6qaMZUKzoI
pm1OY7OFTmGl2B1V4RfZXJx2WTbYPVT4NGNF4ATuIzu71CGYG5N9AV5zgDKP5N5d
i9j5XPKzG3yTZHbKnSQOQmAjba+aCbs6pWW0Rd6CXu4Qc9iCBUnfwTJsB9ixAsiS
/YSvo6QaehEA3rNdEiTiVjBb5rfTFZKYl2Nz/uha9XkiLSUUif2foukYFxgWXxEM
p6S/CqsAHUqpR3LXBnvOEvEZ3IgXPdwYtULo/quz+EeCkS6Yzfk5nN/fUap924zH
XENLd2yv6Wr7V6oSjsJS0vpDSOYWPE7S57JAi/k0eWuR6Mbi66/qgigjP7XMK6pb
A5cIR2ETvWtmynv4My+FMpoLX7NtsSPN+jkml+417WC5jxCRb2kewE5qgu4LqUWG
1Hgjur3fxUU0irluFKdPi4PhY0FsrEbnU+1kQzlC+i1Rfpx/3bQim6jCp0IS6CzB
mQsRyvbN9/P+IdPGyaYvqsMja9wozeJIxd+AB/osH01bMrMuoEBZ5Eoji04slHUT
aMqjEAUaI6mg4lYrs65zNk5HVDjOsEvQMNNJq3Tyo6jkDdSnFsZhMpXpvoKpjwCc
Raey6QIXQvdOyYBz2LfY8rJUr1+hAu8SkRMnlvq1W03MBCxdcEY48oCnhriL2ReA
BqfppXmm9q2plWidAlH8KT4EvtCq++4vFQg+6zQwUcsj0NYqLqzuOIfJP/fldLUY
N4zbjaXzThf5ydOA/aanXw11GWPr3JVnJr/tImV18mYZW5eVyyHSeBT7XLpcsaJU
h6TCw6acb8jJ6ZIGaWSRBTGD2LQjkuzzPJiJ4AGY+MjKvqD2SmGFFrvPENRABu+x
hWx3nXUDYeo1SLqXoarlshZRis7/anjnnW8QZw+5Kzum7oyfUzPOzJq7s39j66Fr
7PtxEdOwZYOAI94VOmmEaZSdI3QeXKZ2IKZsVe8d1MmwTl7kgqm0l0kz/M2rnjmh
pR2DE6cg/uA3tgHK9YIBPELoZpNr/dfop7ee3YlBfjT0eAQS8BZUQgNoFQhw2xXP
/IogjMzIx5KMrlvY13dOYLn6OOT/ZfaU7iN1a+tlLBh+c8JSNCtdxpu/Ms+9Efta
DBlLGsayN8yI+C9JBkHqCbE1hm7wNfr7u+wkQjDWnxk1vWz+s+eBKRaJVaPxwqFw
v82TArCzEEhBifZJMybTPbGYG2Cf5vrKiczbCzgILmemFBf7mK8KChxn8GLZ2TqT
GxZgcDF3tSN6H5h1IakqtIe2F03j6crr3/wTwvZgG3r52KK0tURND+JTevQrtMdd
wPrfOvl+ApGsLzwwE/oAW3M54fbS8tvDwL2SKAjlrI2gmBTc74hW+Wsie21VYfvL
N+I3q0F1lIKDr+Tq4SHpWqnIuM+TMJmODDTSPepuH4jSqAD0C7GzZVPRPIOZ62Zh
Ps2//OJh9UXJDh6sH8TxmLjy5u1jC0mL9o5QAQ2UKCoG1MWcXHYbtETOP+8kIPln
ooUen1rZGLGd1tovGrbv6idzfo/sZgiZVIedG1SqdKJb+tLDq/xsIV1b0CogMgOz
TJBlWAwe+sATyv3TDTT+xTIGr7IxZ1NqC2ZvK1g+W5rTRCrg5IRJURgmW8HHtNkD
jW0Ft/o1/T6yZLq4UXC/8Uizw5FqRAov5+i7oJ5ELDIYwT+bC7V1avf0a379760l
vkurQ5s89S4a/znKBgosItyxWwv7JZ4IsnUNv3IIa+NdHbBga4EoJvWYADoW1aas
WKoE8/1aB6J7j14JH5gsf+HPrlRqXUylIWjExrDlvkgESRUu8qVUlC+UZy3JtqAV
RFo6Sn8sBQumeBpDnblC+Ptjm+rqeWkPsjzVnTknQ+dZhrWTSGFWuvkPdL7+qNMH
msRpZQATRA8m8Zb1Y0moqMJqYRGv51LkJbSrNZIzMEah9QOnIquyE2Qz9rwiW2hA
g16Cj10ZF7BPOSs9IcoWwDPuyImhjS2Qy2w0nuxk75Gxo2Wqw3Zpl5AbqBJi+w2K
E8/s4Etsogi2dHDI2V2YKpIIS+cw5Cmnxza7iyb6dy821bTnc4L7/tVNbJxQdDTh
ANJBH2iu5v4JnpE/sW3c8mqQYVUMiEc0ykmplpnzW8Cvp/WRTMBGwgtitygzDUtS
8oIWUYTEFLQg0JBrO7x8wvnFdrNFlP32qvZRmvE1OkCbdkHmNI3/7GACnTpTkaQb
0AHVZWVVjIPrzCX2SQTl9Pd9POP+tln8NxXgySVM1XmUFZzn2ZN+wyqH+aIGj9ZM
Jt1MZsrJMee01aAnv0ShJ9XQbVBtxcy13CY8GDfgKyEcNYR3DOHaA8jaeuedLWLJ
km8ggx6MB2RlBOcRf5/Hu4Z0/R3NLQt0rGpZhxOgyVozt1C56c8wk6i75jvmeZcE
fWQ/jM0mQwMORXibyIvl/WLrDaEAFVRHK7lO68GhAQbHfZkpkXanEAECxFfYP9ez
35lFTJSq2buTJZh3cWazQXsAxMCjlPl2GrcO7lQF3yczROdf4D9xwye5sB/Kms4K
W0huGdZWxpjqcmHdtoRci7KK8VTNINFkDn5sYi9EHxIVrsJRHVpOAKyXb7ZdLTgZ
OhtU/OwvuC3qP0xYkGGqqiRMccMXfHhEtf4VB6SLI2H7jiOQ/eRtprXoH80mVQ69
Kjp7sM0ay7gzJWNHn8v80xVdlrqlZ8WrftIDKQrBGAw4T5mGTZsZrBZtF+iPKgI+
sipngq2cGYdTM7fmQxCEnQaizstdJJR8K973jcSwerFzMUvsKSYVK1a9+6QyXUET
9lBJlXpxz8zyyn9aqnD0Dr79AlVJfl4uPVCdjfyIsGAPA0yaTRr2czY9zJRDh+tt
OPnQQDtdtEThSCA67VR68Wd+usmWD7+mgS+ZYdv0sbRal+o+szpZT2Dp4/geatRk
sEndaUutMUJyeMaxK1qRhhAITjHNKMmqgDQHUyxGiqG4wu3KUuGp4K0qgO/2VcEv
2AKWWJGnyL15Q80HxmYB8iyyi32ozkh36unRsKJ/vaw6AUnrAeTvEWSHaXEuYjY0
58WImKz9pUlGaCqmGg9sHa9BK/pR/FsYlFU2k1XHm4ykAWavAXtg6QgruDUR2KGu
vXx7Y8JtORY9UU6nFyoBC4b+Vr/x5xh3mSiiM5PT5Yav6qGt80IKwLB3++fsrfDw
qnaZHk4miNdASYyMJqEsNsTrwhqumcNWuMw+w8VlqZZh+qCCaNOCemW9y3HXADy6
OHoBiucTDiYUM3ttd0U9dsLDTFbu4xxalUuOiATn/QNinaupCkHx/b38JHx/8W7s
FgLgDw20N4opPxwoGQjRVOW0FOJTo4J7K4+RZ8b/C1Yxi4tHJXy3tjxnU8s5iBvq
3WsFV7IP1kAaTqOBs7zI51F7phF+gvURtkhDKfgQuJIvOsuR/tOGqKHJMGzP79ew
1VLigW8vy8bt69+okQOHYdQLglDlkvQ8/n7DlvCX6OgQGK7GxOm/rdB9tSkOkUrp
ssoNq2jCcWdFGgyG0gMtoEd4BB7T51j0SndjR3UBt6D0mB9ujCaRew4HISik7I2V
oujrv/+HZVD9bTWufOiwdgDWw7CnZEZXuvVpcq+bTd0U4TeI85XkT4ot4U+h0mN+
8mXXSDge/jzxYh8cC1E5PsB4uvqDwxwJ9k+hteaIgsOmnp2ITbG7GY38ak5fU/3K
zEJUw/gu5FLxvvETMcqxbPBMzdBenBnupCkhz8Pu2HIdK87KJLpsHYz/UHyeqxPR
JyFivDLCKnPmpBM/daojdboF6kLy7fjY1epwgT0ToXH8yOv9roPc3sNs2VRmQ9zM
mrmSGbdTdlTq97y3fsdZ3MrgXyIBMbY2fCVhHbBdSEcSxF1d0lu58Osu3XkNC6Xc
rhCMH4d/mL1I8Hl9IHMhT2yvWJ2TBiY3rmqGa0PWxXCoIttPbEAJZkxzOBgsuo7N
mygHuDGzDy5xnDNtvs50TTSK9XN2CTQ68S5lH0ZNBsaN2zg4phODfHZ0ozTwVAzi
vQ3SCNULeEGHQ8fCElLI1DYn7RPe0lgockw+j4S1rqWeLOSnJIgO8vMMGDUw6PP/
iHu3fI8+9EqEFmV1ocT6i4dz9gS3RdjRle59y9st/UkGh5Mi4OpsA2r9igN3gLzb
WbeZQsChHPq5V/DkNsKrl+aeANBCJnbrSY4NHo8QQqA3qLcd1bfNuBQJnoTF0GeI
dvAWFpgTyHangQH1WGAGkA0EUzYlx3fvP+vtuXuGSpbaKUpIP6VGJ7lvy51/aZgd
w1tXbPgBtVCat/7E1QjvQKIov7z8PoWUgAwG9eoyRxASWE3N51yXtKA/viLXv/qM
XF4VsVpOHQydeZEYlbUOLv81NUMzOK+Yqpi1YtH9erXq6UpJeSscaCWgXFIaawu5
eF05+pPVWW/0xqWBhA9DA/bbKOECjR4vIcFNff/AMhubXpBxCdiyxXBxtSCZrj+h
Jy1UEkQC2oQLjRHN/ql265/zEXgEkHSzU7CB2txw3ldq25BZ+GG6uPzoMRuhpwzB
+mAVxu6W0yt7kw43OsUXVd5K/uKDeiAajlBVN3zY6iTu4xBHTsF4zpqQX4GgRPG2
KHUluJKfp7VZa5LboVoLRjFE4SIjTOUMH7wVREO7CWkloTtrYtFIvgQI1qeTMUKh
XcoJAIetCx4klv8ZPrxhIytouGphwQnOquaCn0l7QjsQ0am3qmlbSHB+PoqZXxXh
xJq1+TVtzOVv18+GYgzemZ+BWowlcKwIfG6J4e7I9R8zdXhRRCjLA5j/49Mp04IH
SnIm2CiikwWssNuN/avVl80PCs324hAwb2XfpAsGjFO5HhaX/ZUmWKZbkXqQDF+H
ygzpWnrHGJlfa1wMoY6TbPSFFnDkeFBWCY+IRu2l7/oS9BwHf4PXqlF6taAvnku0
Qwoqw/isBGJbPnXSq50yuiv8o8vNOzABvATHkHFNX9tIaJmxnaD7KyLG8J9VNK8d
YVnl8r/ggfJVqe8dVZC9LwfLO9/+4WYAo8LKN3p5XptqA2TWgqkMTbfSJZyPhLij
7tGG3YdAjAeATvew8swlUWDDshWLdfrFgXob9hBBzaPWigD8vi/rT4qtm8Xvtw4A
qHjKtyKAIZUq/8PSGhYDAYFaflil9oJsHrVRfmwL/NYs1pd8X1ybZgveLQZ8EQKG
yStpl91mIb1xI5XGAZb5tCvQbLKP8VG2QH+w+EOUvOhCnm5oU2JKHShYAMnYHBd4
4JlAfCAcNtC6bjFWRAfLJnGwzX3PgJbm80KyOfWrmGWEIzbcV2BMENqv4gAt2tmx
NJywPUrn7EsdhOVAPdSjNpsfoc6LKgQllKVrdLlbSw9LXKDQrUQ3vi5kmPGKMLRe
PPlcQgN2TGzcAm+63LLbHS0vGLcRw5r4uHlqJWFhrwIwSq3eQ2vMbY7A09ClOiiG
/qt2i8920ohQGcnG5AlRdS4xKOsDktdKcwQXZJL82WMqnPqsqn956C8qsP04Yp31
E0dNSnI5Mg0aDRs+igL97EfYXsnGp6dbfX0isSuSJCZg/SBNINNo9epmPIN7QjSR
eYWpAQn2mFxtPhyNWpYaJ4AZTVnf3XfQN4AlKEJ/Lsm3rBP4IGtREnReElI4Lh25
4YDtXBuM2QfxbIcSiGSV243KdZhZ7W5FG4kUjnrQdQFzBu17BYPNDHPpIRh2GDJk
O4185/n5wfaE3CTF9mY5IT8UmcG0eRKW/hXrhmR4Lzb6tCP8DutIxfuFmJFuLheG
BV9rVOyMhO5Q9bf1LWC87XPunZWDCzCOyjWivN8B+hbZvUWaYG0PVJ/3wN3rSzjS
oB8Glqy2Um6f06WXgxQ3YmkrJRlL9p3NEgT9DArU21mnB+cWmZsXluYWAtQVFf6V
s7rH1wZLfBDeji6nzVl0p1eHeLn9NnItFbDsfKtfQJ2dR9QaIRam978CJxU15L8d
NzGpWcnAil7Pz0678OYOVwCARxqbvA+5TH6RSAcPSKqZvh3UsGspBuR8qaDqf9uw
VnszmRGX/XbNY+vMCNpYyKerlw8INuob3zYfTn/rFYORPdpoRNZR0/Eb9kMkpqYU
hPCfo790tkVb9v1BUlvY4zC4il5e7f6WBhfaQgHaY8CdJz2ptOYiO7ggm60RPWDU
JsOisq/WREPIpY/L7uF9YfxQYqcxo7VsKbNbBUobqRSD/54jPI2UfxB1uPJRJQ0B
hZX+TvEou4M6UUGYASHB5R9bGZSALWh54iwYLfwo49+SoWwbD6K5t4N3nUlpvX5Y
AXAJacLMvUxj2aGK9aEIz90FNkH07v43AUEi0v0eKB/k/woq0J0eqSDQrHo9FRpi
ptPuJUWeQLH5C2oIn9YQrN25D4uDh3/sjDjPR3duXbqd7/qCmGpSYs+UmhliroFt
WXmcPCT6CuHQK/+V3J9GxNq10BysZ1vzGqAjtD3ZjzWZTn23/ZXP5/j2kNFR8+aT
Swo4ihs7Ar9Cvl0xEzYGe6ecmcbQTEw7hl0xDgiDa8axr1ra77nw3WHVI0V1IE1s
Qk5Ho6GBUj1d7Q/3HoedNNRyiBaz2TuAYLzXurZuzhZeK6DxWnYx+sRpcCjHBqIT
PHoPZoXxx5qZ0buJ8CZdYnTA7/DFSV/HUvCpLi90tzxxfJVd+Y203dMJVD9g6pIV
UnNdpWnO3ppfzUKpDdYf/5O3+sU0Jc5mRXNejLsySbb5sgaZsP6xbQtEVfSFytvH
v7+516BJMqg7Kq3ec2wfjrm7MdT2oVSQ4vkEFmvh13iDCTCLXVPNaLCC4DphSBGW
VuUJkyB4T4zKORdFFqHE5mnJHXUvoaldNX0l6zJwVZAgZPu5YCymCSxmTrq6N7Cs
bqUDOL9/cVmyzZn2gDa6H8qb1dbj6Y2AE64DIK9bspKi0tigD8qehPgnXF9zevsg
jF40yo/Fv9OusZmpd5YkcVdEyCYR6RTjNFPNEA9ytHBeHwePDt5R5Efgxdkwcd1O
dgLF6ngRUMYAsS87MNhxUp4v3zuevenvtl/tBJ6+1jL4d43knPQ76SDIH4mr8OTq
2a/NyniIItMAbQQFYiUnk28ZGXXgYAt6u/B2hrZK3cYfKNBI/Gyhc2nrDNZtvpYK
X9FC2yn8DME3cB3Vm2iADUEcSiStjX2dsDBEhQc+lkJfDeW1IJMYXtM7fh9nOGqS
zbnBqjf2Otv9lj6djIY+AmkjcHifdl/0K5Xns6aYQFSQVVjff29UGSOIDFd9/FuQ
GTNPewB2HHQTrIeQq0OHQ1LWwKr769VUb145xhoWowPdRpVzVVLz0B7ppJzPy89x
1Dtm5autgO6do8+/z4+ZA+e9jXUNn6FrNAinoygbKMGxOpndeUngikUPzXmroP/L
PMy04v7azymPi5IpN+XlY1oEPYKq11NvkR/TraL7x+hlL9mAMOE2OWgJM/qWCQQ6
ppIN/4wGaaWGtlgf5vf8dh5cReQvUPqyhlNRqv+8PH/xKo6TEdMOEYRZnD33F0Da
xKxlrZ13ZqC8k3FiWeTLtV30iU0/QKBZkUaTQIxJlHx6kFybxBm4XlxGNcx+Qxnj
1CDMBbLWsjcshthHzk8HzYNEQzkQoqaGnnA96br6SHseQhIMElu/W27I9Q29K3Hm
0OHluSzmPjl/QVtDTeY67NRgHvHIMG4HKdnujXQdaNorTXU2FQ77cT5w2VibwxjK
oKYUigZUlxEV+7OHIJNfO97vaM87ZHI6Z6SFI9oc7yYCjnxANhmlUMshpigU3eS+
NJNHfVlmPzLiJaZR2UpYcAyYT4kJ28wjhqnO0fhTkjVrSGtqog5LEAIirqWksFQi
fi7cNDyPF9+SEjL/pQYz56FVvlW7pb9FfK4PekQfTKkQcDXNstnjc1tdz3OmZEIf
7vEvGUitTkfJ/RCYCvfg4fuoGxc/DE1Y6rbvcw1HOXo8zKA1qGBxRW+I9WuhumUK
iaT3ZCIdt3Kw7fL8vwB3NorECOS1Bf5qWPOAOTUGGZvlL4wGWQuuW4G8C5qjXJ/m
cCMNT23XAKIMleIbweAj+bxVj0SYljOPox1RiQfA4X0zGx0+nsLLMAi1IC3v5Hvx
9sefzHeGe8sOrPHWqmM0tr/efy8l45JvwQSS5JknNc6TiXLnZKfTOB1fUNAjLWLZ
2bHOOPK4kpk0UMJIsqJNQGjoydmos6kbUgxu0LSN2k/848iCdpYZyyfZtIu+gzKN
scMciHyGQ8yNdSZTSe9AHmg0IJXgTZlnXECIj6sTrZBSplPpKTN7pZDjEwung1Xt
fcewXIoZsWlj/nYIVYbZvpKxFMQnkhXg1N+Dc278kOgMoMZb0Od8/YggvUkfnnY/
CCKFbb1WaQmZ6rNd6EWScpBe23ldL41a8zt5K7yg4xtAQDgl3b9VOJhHgJr8tW04
bkgF0aJfABeQ9YLrSiyTHfeeI7R+5F6s7SR3xFoUVLY7TBli1sSVw0viN4OLjELT
uTlr0Q4sl+GR+xaILxjYVUeCBZT67CqOX8YZ2k+Sj8udMGjFiFXOH9sw+I7OPc5G
XqO71RF+xemUZPva0qJDchaG1IQcdtEZEvdek5RVDOJqoqpbIPWpIUAACAejrWQj
QyCcnbAtGEKO0n46tr31QuIx4oC/g7Z8sVm0jVvnFwiay9UxdAdfOriT7chtr1pP
wIGrBVwyhUbahGmzIHTQmBZ89S3+Lx+CFk2bYpBt/+xgWF8qz2230mKzOORfUy/k
bsWIcA7rauo36rZ+qUyPEEW1dZCFhRgfnpo7TjONDw8yhda1Z4SrDxNfK1Wp+cmR
10oiHui9Uw9BMbr5WlP4afdAZ729+Iuw7dgj6PBEn49aJsV81cplyOadB83HUncg
NIqWiFNdQVlxGfXFvO6Ott2wNlVKdh3ylBXzcXd85ZC6nNwR3S5sQrKWP9rEd8zV
xumzZWJOUHfPAqKXv+HZJpSpGGR+VZgWKmF9T1dQ8iyYnVO/psa8UhSc7k+bDAH+
ApdhCownF7prNSiRiw8/CqMBevrCUDizhKDZD5lwf9QQbFgUnBQvTI2uxOwYMlUv
kl0BIeJ5pZ4FOhBY4zkh2eNf5tr7X9leAEjDmsJe77/wpn9dUW9mXvfwDF3bA1fn
V4b1L6GOxv6j86TLt1OthoeiuRkmdFTXeXkev03AWqxymKG4TlBp3d3G1/xazFAJ
BvE/Bx3epEJIk8QHGYuwo8AJJTvC4Oehv+p+nabNXWHZsYcgvSW7tT2gIkih7gNv
If8QKrCMibInuS+3kU/rIzV2k7IVG0axUOgsPjQYnzp/A7F74Nmop36Sz1N0KwJb
Wdflw1luE6BOHh1vGBojSwIvwWVVrnu5vUuBrsvax3zMmV5hekFUFJkwg4pS6+6n
wn8wehGHdfuNTSdBFXNIjtEbL5tHaqkCCSAzOiR0W4blSrfb6NuRd6EcKn4PFWKQ
IZO4KtKzJ6ysjsbiybQM1klxjRktAElD5BCyNgS16yrYXFROISZQz0ZdLWwjc+dS
IyH9ZUA5i/yDg/09YvdFmT/Mgm7jdpg8PO/s0kB/Hu66HkYdYrDYWOLc9IFBkBkE
axTQu1OFi+o9nxWhqwT4o1QiarqGzXQ0+BfzHK3jsKGyZVJIeKr7udD1Cxw0MppE
FKZcXkJX8mp+JpuPOxJUz62KAlJZZhsinqQ1Vd0LixTOpR6YLs2iHbojVwIG0Bvx
z1t48kzjSGavEt24oCQsyC25uMpyPw7JaPXPZUDR/q/RNh1UyFtJFxBUl1j+G8T3
hdVI0UzkviWBqsuWSdJuBOY4CLePSo8V3XmLgKe1gZOmjFGxjPTT9HC9nzcWllP0
Nl1uxjJJgAzem5SJ14nLLN6TJ/+H0NqWeMZ/+i2UAW05n6ro7kW+0nfQ4+qI2FQ7
eN16KztPe3D+N04n6woCqO+YYC7URzzJ7Mt/keS/skMEhVNuO9VPQeOK3UNZ9bxK
jUDKQUPWzyGn78MdmiTAXOCFn7QU2AXHQ6qhzCU16DwWbytdnajHhrdc5HokKos4
R1DD0RTA+ub2uYKHUepUCiZzH2ojqC9zTZUQvZPEiF1u8XbiJqB/9zae5ZEd0ozi
P//pwKjY4UBloBS6i6Zc2rSxSBGu36Op/EC9Ko8LgNkk4tdLOk+i1syZMQWqDK90
0rqbSUBoTHVRd43kYWakyRcQQ7c3rbC9Zt+TbR5llJOdJ6+Bb/4e52HrRq0uC6Dl
zfDD8TSk0NWs+0ES93Neu1HCtzVkI8qq4zG8/xYUeEOac5aZst40XBU7On8MbzUF
Q+Soo0BCnXdUDVR4Y+Tn6YK0jG+atqiQMcQMKT8rNVLLBjr0EWytuUz38Po3J3GW
lFmLY41VY7zh/BEPZEWOLFjXnM3pxpE6ZS2KIMs13fm+sMhCCh4YNj+cgWGWdXD2
CsQU/45wLGDvsSUppNM0CZR9iYnOFwanmg+0aiUVeMwfj8lCDr1TyJEPME+txbkZ
oSfIhMgNVnh/Z4oCyoIu7iudRGOy2ha5V/yyv9CKssM8nX3Ssv6XY61FPqHongYn
2xzYVaWp4U2NKl/VPgmIN2xtWGclIJK2JsMEvSWy5b2aolAK25fk3zSlhpzY4PdF
458kUlYwZxCfWXAAOBgI9pRJWJhcx1OnL7VU8LjeO+FejgXuo6Ss0jeG5qxTOHdn
SMXQ6Lp+Ozw06mBAeZFBUM0bPANaTVmHhFMCQ4FU86qY/dvHdic/LakYz+PQx0iT
Gtvz1/YRJKT6ncwcBxHgacLQ1VjgWug2ZOW2FmuTebSXh8QXrrISZxkUHSZK9dxF
IGJCsXnczBqMD8vLaML0/XSouxLd1MDUBielMOFoEWN9nia8h7jMkUDeieNBOisq
BEs8zK1C2r9Pmz6ROSmw3SPIx/DDsHpeocBf8O+Gf/kw+q7Uwm/1pcH32rBr5SPo
zn2AYC2E7LXGwRIIWyFuaq7uNjpSHYqzZyOA5LbPg11ks0inC6tonu0+qhMA89j/
Rmb4+Que5ahO1K4Ad4EYq+CkgNqxAIG/7Hzu1TaACZNaHJJXkKw3YqvaSdatBlht
aQ1qQ/GrUbNZStQF9jWljCn3VjPIRyeWQiO3UXGII2S81sHSGIcDKSuDo2VOSRBU
PmWdC4tXKrZ8CQPUjfaWv6alGJdgIvimlKg7cm/Prj+GOyBe32hSTAUm81vCSrqZ
jAYoYQiYSP908iowhW1kh6ZAzLBqDhTlgqomN5b8Q+h2FIhKabM1IzmNAiv/cl0P
dIXqorPDuu+jH/5UQ5pKzRH3qt4yctDfDfswDqJ1ks899l81MeMfzxAR61M2q0U7
rvm8doQVyMtrIj1F8E7X+EzTB/pmdzteqQkMpuKBipU5OyOZuI8l0fUhsA2LulLj
Rq+r2Cdi1pGsTwQcMTFNX3jukJzGOUAN5gt693fnIrx038Ugt97+3WNJBbxiPCHM
hOIOvLa4yaJxX5YBPtBehhji4h7YOuKm1Xhum5BIt/WiMSS2VfzI4wGofENsedCc
8ubE3Hm/tELf2f+IfIaufgJ4JiqG9mclIddcjo0328nIXm3SM/dxFn3srSR3yJ4q
Lw39VPz/K4xR46pRP1QSKvH6THFenLhjQLq6sObohEMQXaBXtSjFPaL/Nr+DH6LM
OPxM9SfpItauWlPbLc9VKA+CXgKOFabjjpYdUmRJxhU0py6+ZBJVrJegmfdE5/Uo
sn7YLYGtxnThvC8CsJUCp5P1ui/P7UfnGB4RHYM/ueV1VTrDgo3J5yk6v9N1F/ez
rtkHck2EiugkJ75fX1/BpOyFvtTjZJz5iqgy0goqd3OFjsTKa5UrdqW95k6Tl8Ca
0k07yBeiciKNopkUSb6jiHq2tLYHdxNItktwEKFCd+5sCUrpnuNlFbikfSMvp1L/
+4uuOPAvU52Xr5/z8Pbk3mhYV00cUUSR7b3H7rTjLl18dEn6I5VZzvK3tpSvbbJ7
uHnyCVJKnGOqvm8BuW/Tm75q3U8rU4sbdLWDZyAPrpMpE06TKb6x9cfwyN36PuX5
MmbmDYUluqzzCcy3rxFuePF4x4iHej7f9eFCfK6ABr7FHgO7csUAK2uiSe4OVuVb
zEHHcdgD5HgAX8qimzDMhNtZ5Rh84a1jwiDENEG4VLiWCeX0Sm6K/DhTHseiopqV
qIwyp8g76jhQHIvowpeKlAfHAUkue4hRB8jnSs/AvIL0WCV/weFqbjG7sSr8p8qN
Tt6oAG0RcKF7oHFItZDDG60XN9VgdALOn+M26BDJ2l56Q6DcJIH3T0lwnriUkOCm
el83WjFMAOnY3AwHvBWGg0f+SKAWvPX6YJy6z+59cpCvy46kI9hcmSWj/Q0jaDoo
VtRBJSl+hZyhi4LsKdZMZRUrGi6IaItAZ9SXZ3ZCytjJo6ZKDBj4tWEveitROH/M
PyunBoXCM18OjoLieF9XZDModrkmKi9+B5XiqnLBgEA5YMUZK6E+q2gQDkGB3o0U
W7gkDW+2hMheM6KNVcjAvJh/tuJu5fzyygVkM637wZACdnGKuhezHpKm3fPFk28X
LAod+LzjZ8TOaGlNDeyjEg1ZFBXthsujK0SSPlCyhIqZLDsYXf7zKQiKE50t2El1
gEEk7QhKIF4z4kY3iTU0DbGXyA8dzz109KNvB1RZO+uxkO453vb4p2aVyTPdvK0w
zWM6nbrajqACtQ8y/GGgt603dNQsgXEKFraGcdHQsHwuSihQTVCnjCsYAsWotbHM
ROsgR3sLBE+AHmMLDL4LiNnciFU76IkaBtkh8QdYO7fWK82JlflFqG2wHivf2Ln6
wp0uaDNR4K5jxeww63FgdBJKYv7dkWte1L8f1Nu3txfqz8AEf+jE63wPnmWBOgv1
7+5dsBIPwJwg6Kfz5zCNKbP0604Pm4qXy3uS0xIxy2dbimXshi52wp1fCfUptHAT
cpC21uzr+Wn4woSILMjG4KMNPP2EKc82j/59l/IIVluw3FBZnRPVBCD9SmJJWiyB
dZ20QJhiCekEJY9zCHTRBXnBYs9Qo76DOpA4L6o9IXYujWS2mhl/AshP/knmWuB7
GZqcM7MDSimj9AAuI/z4LlFU+fehI4fwwkMmTT0XKv2uAnxP958tJWpoiUYlmQXS
CxPLdXwoMnct5IsrfYdnUtrG48SvgPF1JiWPrvYgFCymn/3SiQEBAx1pkR+wEZce
jbFziqAfjESokxz8v7HJhXFqrfCfSZ6oirx74Ik9MbMBeBwOMZnVhkjeVizaaydo
PjxGhd/Rzqtp5odXJ4khxqvsf6e4b7cAE/JlPN8oT8u7qQK1XVsr75ldnl8mVYu/
R7Z2M87dK0slTvV805WcjQ6+67GZl1K/1P2pT5Mc0NSjPjSn3Ln9X5Y46zlZ033q
0/yp4+FHgzVF9EQs24Wy3hFszh72GQxHB7wnrQcCGqmhlQmloMT6E3f7XUiSd0OT
aWtET9UOGio3jWiuwDTO4wYuvLRpIJdjRVaHwX4Bugv6RyvGFYjRV4XiDqniD4xu
gHKPp3HeuRnYkVMyfqVkeI7bT0bNDA1vM5rheBN52x0MXGNr5nXUoj4ayv5RHhJl
KWEeJHa0B6Vcashpy435P7yhtpW10y4hGz62erm8WlY/y0+5XZfF/igiMvPGViSx
zxZ9EM3q9QhfH5kqknsfiaUpAsQ6eAJU5H8scOlyA5wjUfVFdxjOEf6Zeei3PM04
odFB1KN2sGxdK7brJ/3A6HlWcKSMON8ShRmsvIOfJztQtAtIf5qkElYwwHs8oLOs
3jBfDHbLIQnsRUtp/isDp79Phkhdt+BRDoXjaWaZO+U6TmrXHay8niRybu2MlgTa
9R5mb3ftFTa7Atw73Yqpg5FzAVzB9/SUtmBi/QxoZZyM/U84Ry3xewJL+0rAaTDV
B/O2ewPaJHSgSzN79MEs4rZjUtIlVKss+a0PPsvVSzo2zZoFk5YKWgAX0N34vEhH
YUp1T3ZX90FALWwinQ1UJWDSB05OKr69wHSYMgepbDpUh0Wvq3+m859zkQRrTB4b
5bGh8XNHNnp4eNtqO86A/lgtSm8Vzctxo6pkJlw7C9EqNtEOzA49apxyuEuCoeJP
91QMA+4lyEDMMx+Mum4s0FXEy0UG3aU9bJZIyodobI+FGDGwFqQmmAR3mQ0QDNT7
1Fsl7bRy3kjYb7EDK6/n1tx6XbwWMcLjTz/6XPulisK5ci74+WTbShMYOi7veeSA
zFryiUtEKOJsuRVvxTmWWH2JO3+xkf6otvk85A16BBmNjHEi3QF8qExp/qZGyoWg
57UXOecOFyq2ycPlkz/76fcTz9HfRUfmC3Bz8wTy2m0qGgTwHsRPAbhT8ikbdSVx
3WY4bRS83aUdoGl/cVPcolEHWIjq1KBeNYmTmn1n+RGvI1xYryVN+19oIfiU4qNT
styFKPdOvNULiObtMR7AZNA0hLaYRmaaIMoD3h8zjMmkBt1qgGWx4xTH9l5a7DJl
f73j4QBHQKvrb36mm6JiSRx6dhecuP87XlMD/8FSJqGtiY8apv8+Uya59UNTt7oz
Tg7PrY2Rs1H6Q2Jzy9EzfmsWor3cqphTBE7yKDNK7REcXCBnN45BTSTpufsyLg+M
vDjeLXBQ/nM3h40MoMDdIKwisUlQN0qWB3lJrML9KxBe/Ndf6pC1/c4mFct5gRqP
eQjK+8qzF0iu2Sy95EBTVRkYzpMvwzcrRiDA8bg1nYUwPzsf9FTvTb9ygtqG9N3/
6Oq7koEbqQAAk78LGytOSf65IA9cGfYyHOPJCfPfVCtLQwxsFx0iXqyh7j0bDs6l
rkBUmeg8hzY4AIKkyaDjGmNoRVpGkMW4749WPOBh1kYTMqLRFbJx1NtAVgMR5TSe
nCMYKq27viuycOisgyZqMSChy/qlH+xa8EVRFCT42rZNuOwrvV8RtYu3psxT1sQ5
28NJluPOOzTW0JJ470V8XBjyQ0Bw6+bDhjgSB87VPKOtTblNNy1SBugSiKrtnivc
dqxjRTwoQdOJ68cTqqEHVvuCNzVj+ucE7Ql1x/QZwvL0aYJOgGYImqaNSUKqyiqs
EmjJ8txTUV5Z3fqnD0k3AA76Z+ZlXqdrmNcYUaw0aKa701EZPBvUB+DokectkN/z
SoP7I3KF6KYUe2SvJ0r70V+REwI2AJepgHc+5mG2857GSNRPjRmOg5tw5eLeVxIV
poLKo7hwDs26K7RW6iOumS5ZJwO9CTWeNdAyfBPPoSgppY/plQbseY+XKO6cfJGX
VCTboTCHSPg13F7lyV75bJ94msU6pWsMaLzh4AawQdWGavp8F2lRdl1/+uwqX0cb
nSFygElHqcV5HFrgBgNpGgii+CKI8CLj6bMjeipMpA0ULPjdmQwCSnHY5GZIq8wL
SlbC+s51kjYi2xuQjjNwoeJdpqL0cV+OaitCJzRbaLmfPHGEU7LCNcq6VV1AsZSR
n+r3Gz9CmtESI6gCJX576Q6AKPeHO5EqU0TSqrCDUSQ5Zox2OeAwLlMgFJfDEQGg
gOZN6J6YqkDDULpcLVJdLiWM49omIKsRcGuPaQaL+w4lfvAnoI8pZlSWSISl7Ey1
1me5sEVhtkuuUNoGwgzaTjv0plsQ7IxDrIWcNtm8BtCQMy3Nm9sKfNpDJEuJztIN
pxPnV0FylAueVtEaAcX62WIQhQByqbD3RQRRKA6GfxiF/OmIDHP/FHdvwTuCYjMB
UGSGjlkAMjwJlBZiFM3q/nLhzgJo3EoIB9c5PoF6BIbky3VGgkX1kEwycUEZcsFT
bHPcjG8xMv/g+9H1OddXLyddgiKc/eJwUbuezQCGzqeR0Pfm5lTAlQ87JyBscmlR
5LsFP5w9YiQwh7Zfcat8dZO7Uga0rvT9j82u2lPxqYV5eyaDFveAXGfp400HTGv+
yMl+WVCpRCFqSNMiqHcQJ6lY52hvT6dCDbMOd9FzQ01qs/TtyD1quGq0C79PmT/P
GAggQy9CS5ISiSr7/uoVgCOtBYmeUDg1pvjTzAgXLBMimrDoQmhiedmuUFk/Llih
GwLads/J6xa++OMqQ63BW7hd2x1TIHZtrIyt6wuob5QDBUDKsswOBp1dRdb0Um6I
jHz8saN4YwzCzl/qmnt0toQSyB+oqXHJpP6YhY1SdbGWH7hpknRgULtmMHW//gxO
YizayTHFQPTYsWOUSn1Cs1E0YLe2pACfh8l3FgVBbNT59KklpkDdJmYC/9ykrc7N
qZXZvU0b0UtZ1VRdeHDmw9e1/pT9CBFkEMMB6sClQU5c8FcLeRsyDXoZ66HaukyI
xobdvIG00+VskYmF4ZJC3Fv7XZAK40paiwv+7zzJOfrZzK+32xBG0Qun1mRCmwUc
OScTwE5HayIKPm7q5r39vMcz8a0INJIzjdomFU6v3byEkvRrQH23F+fPHQcUFndS
0dhVpYNQ7QEtWU1iqXo4ONobuZA0KHPOzdF4YxmtEb8uRtvI7V/6tCvpAgDlU37p
aisCcUz8ideXu9ohWYK8iIN2YXTLpxhX2u+H8eDNx1wpwvKE4H5oBe/LYS0z5VAb
h4crABQNmAbkzByidbB3yINL61ZyT2SPDBLTJ6sZ6x/wiAWW7BUtxeb6EYhJ/RdK
eqliHsS147G9mxVWf+pj3498g4smn48HLj8IRy9W6TVgzzm1d/1h7LFNkIXKXtey
/wBP+pKkYMaQZmxMxS/N/9Hcllu5puVG9A2RAsZ6mg4LnSKyMZY386nagLDmIIPV
blM9cwIrJyePdVb6QTS8ulXb6qi04tQCPlsvk/UWJEtSrTe2cuSrUAUsgKG460Rx
G93wPP5QtHis3GJfy3kwoqPmKLZAGcavaTUVUmM65nzTeYzM9x+zYxG5vqBzBu1m
J/uHXRY286lO4ADwHLlOaS5UrfSu+Hc0KSxn1BiIZVZdof+0yHEnDH/8WjYQ3El1
QxZU2b74pX02YN6Xas87jHlj/9MsUoeYvsJcOpewEfHy04o2XUF82uqEPohRMofj
ZpfqTdS1/dns7w8icPEyVLhHV6AumaGmcsJO4CM8K7neeozYLr813sT1jGZymkt4
Ht+0+MPyX7RAO2LNu3oDj1ejDnvVzZoPFrCzvfM7g+M=
`pragma protect end_protected

`endif //GUARD_SVT_CHI_SCENARIO_COVERAGE_DATABASE_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
KlGKPBzQOxsDON8pZ/hGY/hR8J/YIcx5OVDrqm4x3w6GMg6tKupNxqI8l7LXBvAI
5sX40NI6J30ivq/d9acrmHCFbuXcWMw1dcYsQPFSyv2YaGd75H2HEHEUnBhF9zI/
xz3HMUjogLIStGHfZkLrG40IUY9cJ1v9hygsaGT6Drk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 127923    )
7c9HFXybtupC+Yfv0u4MdvUTqBeFEsWd/LbUoeE/tU+KyqumXjHJOLBQ19SfwNbs
MHT/R584XeadC1TQXAsoZwUnkZMWeUn65VAfjYlc7w87R0sI5fO2S8cV9DM+XDqI
`pragma protect end_protected
