
`ifndef GUARD_SVT_AHB_SYSTEM_ENV_SV
`define GUARD_SVT_AHB_SYSTEM_ENV_SV

// =============================================================================
/** This class is the System ENV class which contains all of the elements of an
 * AHB System. The AHB System ENV encapsulates master agents, slave agents,
 * system sequencer, system monitor and the system configuration.
 * 
 * The number of master and slave agents is configured based on the system
 * configuration provided by the user. In the build phase, the System ENV
 * builds the master and slave agents. After the master & slave agents are
 * built, the System ENV configures them using the configuration information
 * available in the system configuration.
 */
class svt_ahb_system_env extends svt_env;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual svt_ahb_if svt_ahb_vif;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AHB System virtual interface */
  svt_ahb_vif vif;

  /* AHB Master components */
  svt_ahb_master_agent master[$];

  /* AHB Slave components */
  svt_ahb_slave_agent slave[$];

  /* AHB System sequencer is a virtual sequencer with references to each master
   * and slave sequencers in the system.
   */
  svt_ahb_system_sequencer sequencer;

  /** AHB System Level Monitor */
  svt_ahb_system_monitor system_monitor;
  
  /** AHB System Level Checker whose checks are called from system_monitor */
  svt_ahb_system_checker system_checker;

  /** AHB System Level Transaction Coverage Callback */
  svt_ahb_system_monitor_def_cov_callback sys_mon_trans_cov_cb;

  /** The AHB Bus component. 
   */
  svt_ahb_bus_env bus;

  
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
/** @cond PRIVATE */
  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_system_configuration cfg_snapshot;

`ifdef SVT_UVM_TECHNOLOGY
  /** Fifo into which transactions from master to BUS are put when system checker is enabled */ 
  uvm_tlm_fifo#(svt_ahb_master_transaction)  ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from master to BUS are put when system checker is enabled 
    * Used by AMBA System Monitor 
    */ 
  uvm_tlm_fifo#(svt_ahb_master_transaction)  amba_ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled */ 
  uvm_tlm_fifo#(svt_ahb_transaction)  ahb_bus_to_slv_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled 
    * Used by AMBA System Monitor */ 
  uvm_tlm_fifo#(svt_ahb_transaction)  amba_ahb_bus_to_slv_transaction_fifo;
`elsif SVT_OVM_TECHNOLOGY
  /** Fifo into which transactions from master to BUS are put when system checker is enabled */ 
  tlm_fifo#(svt_ahb_master_transaction)  ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled */ 
  tlm_fifo#(svt_ahb_transaction)  ahb_bus_to_slv_transaction_fifo;

  /** Fifo into which transactions from master to BUS are put when system checker is enabled 
    * Used by AMBA System Monitor 
    */ 
  tlm_fifo#(svt_ahb_master_transaction)  amba_ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled 
    * Used by AMBA System Monitor 
    */ 
  tlm_fifo#(svt_ahb_transaction)  amba_ahb_bus_to_slv_transaction_fifo;
`endif


  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
 /* External AHB Master components */
  local svt_ahb_master_agent external_ahb_master_agent[int];

  /* External AHB Slave components */
  local svt_ahb_slave_agent external_ahb_slave_agent[int];

  /* External AHB Master component Port Configuraiton */
  local svt_ahb_master_configuration external_master_agent_cfg[int];

  /* External AHB Slave component Port Configuraiton */
  local svt_ahb_slave_configuration external_slave_agent_cfg[int];

  /** Configuration object for this ENV. */
  local svt_ahb_system_configuration cfg;

  /** Address mapper for the AHB system */
  local svt_mem_address_mapper mem_addr_mapper;

  /** MEM System Backdoor class which provides a system level view of the memory map */
  local svt_ahb_mem_system_backdoor mem_system_backdoor;

  /** MEM System Backdoor class which provides the global view of the memory map */
  local svt_ahb_mem_system_backdoor global_mem_system_backdoor;

/** @endcond */

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `svt_xvm_component_utils_begin(svt_ahb_system_env)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE);
  `svt_xvm_component_utils_end

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new ENV instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name = "svt_ahb_system_env", `SVT_XVM(component) parent = null);

  /** Obtains the System Memory Manager system backdoor class for this AHB system */
  extern function svt_ahb_mem_system_backdoor get_mem_system_backdoor();

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the sub-agent components.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif

  /**
  * Report Phase
  * Reports performance statistics
  */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void report_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void report();
`endif


  // ---------------------------------------------------------------------------
  /**
   * Connect Phase:
   * Connects the virtual sequencer to the sub-sequencers
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  // ---------------------------------------------------------------------------
  /**
   * End of elaboration Phase
   * Displays the environment configuration.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void end_of_elaboration_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void end_of_elaboration();
`endif  
  
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the ENV configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

/** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  /**
   * Obtain the address mapper for the AHB System
   */
  extern function svt_mem_address_mapper get_mem_address_mapper();

  /** Obtains the Global System Memory Manager system backdoor class for this AHB system */
  extern function svt_ahb_mem_system_backdoor get_global_mem_system_backdoor();
/** @endcond */

  /**
    * Enables AHB System Env class svt_ahb_system_env to use external master
    * agent which is already created outside svt_ahb_system_env.  User needs to
    * provide external master agent handle and its corresponding master index
    * number. It is important that user creates System Configuration including
    * the port configuration which is supposed to be used by the external
    * master agent.
    * 
    * If system env doesn't find any external master agent for a specific index
    * then it creates one on its own. So, it is important for user to set system
    * configuration with correct number of master agents considering external
    * master agents and set specific master index for which external agent needs
    * to be used. It is allowed to instantiate some master agents within the
    * svt_ahb_system_env, and some master agents externally. User needs to take
    * care of correctly specifying the indices of external master agents to this
    * method.
    *
    * @param index Index of the master agent which is external to the AHB System Env
    *
    * @param mstr Handle of the master agent which is external to the AHB System Env
    *
    * @param mstr_cfg This parameter is not yet supported.
    *
    * Example:  for(int i=0; i<5; i++) ahb_system_env.set_external_master_agent(i,ahb_master_agent[i]);
    *
    */
  extern function void set_external_master_agent(int index, svt_ahb_master_agent mstr, svt_ahb_master_configuration mstr_cfg=null);

  /**
    * Enables AHB System Env class svt_ahb_system_env to use external slave
    * agent which is already created outside svt_ahb_system_env.  User needs to
    * provide external slave agent handle and its corresponding slave index
    * number. It is important that user creates System Configuration including
    * the port configuration which is supposed to be used by the external
    * slave agent.
    * 
    * If system env doesn't find any external slave agent for a specific index
    * then it creates one on its own. So, it is important for user to set system
    * configuration with correct number of slave agents considering external
    * slave agents and set specific slave index for which external agent needs
    * to be used. It is allowed to instantiate some slave agents within the
    * svt_ahb_system_env, and some slave agents externally. User needs to take
    * care of correctly specifying the indices of external slave agents to this
    * method.
    *
    * @param index Index of the slave agent which is external to the AHB System Env
    *
    * @param slv Handle of the slave agent which is external to the AHB System Env
    *
    * @param slv_cfg This parameter is not yet supported.
    *
    * Example:  for(int i=0; i<5; i++) ahb_system_env.set_external_slave_agent(i,ahb_slave_agent[i]);
    */
  extern function void set_external_slave_agent(int index, svt_ahb_slave_agent slv, svt_ahb_slave_configuration slv_cfg=null);

  /** @cond PRIVATE */
  extern function void set_external_master_agent_array(svt_ahb_master_agent mstr[int], svt_ahb_master_configuration mstr_cfg[int]);
  extern function void set_external_slave_agent_array(svt_ahb_slave_agent slv[int], svt_ahb_slave_configuration slv_cfg[int]);
  /** @endcond */

endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
xuhFBAabV8mf2WNpeNfhz6XVz845tOComaSY7i7WS1SdpSTU8azG8N7Q6u15er2r
0WZDKjxJdnqweaNvimwijP/dmfq57Sf2bhQ0HjQaGHpZ8lhqYutsuCyUuXe8Pslp
vzwWAtexk6YWJk/35nyrjkWDWd49wChwUR9CmQDEf9qlIFtRIDRmYw==
//pragma protect end_key_block
//pragma protect digest_block
nWCHT2Qlcm8gsU2Hb/PLOZss0Ao=
//pragma protect end_digest_block
//pragma protect data_block
V7Wc5Q3eZ8Uf87ivN5diT+KDBmxxVsUv6encFz63YNNmqbo3i9zImD8gts6n1yzI
+L6LZ3QDLtdMDLIsHfLZBLiF5y4AGjJxXJVIIa3h66fNBQ1KKL+gZYIDP1qy2wUW
TAVe0P+vI1GZ08wtN3nZhaNeoQGOE1UrScRbYQt5EJ/oZ7BWS5rzz9d3pC2I4ij5
vc3JLm5uQHRF4vLvw45W1O4N1uKirj/PVucRAnAWha9rG71Lk2H0/FdA2hsztVYR
8ccovXT5sk6l/D581KZ70Zt+lKnK84rHSI04WT+RqnBjB65r3eBkNiD+BJd33xVl
Z3INff0Rg0G7Bnl2Q6HzsstmfMT9eC2Jm/rkSX4dUEgkcA0S4a4O0Lg0WTcofY/5
kygLpCI3ZmaLH43zIy1Jg+akMh3mVsMtdAXp0gv8MMrX7CJJWyB366CoWkE//yhI
vTf7Nm5v4I5I759TaONCcHbHYVkrjtDip4N4891lV04G23BMlqc/ymxmzCyxbG6r
/E/wrsw9RwaCAoFaZBedgHmCN21Xcp4HW1Sb18q1zpQ6IaszOfLLzyiXG7YzEaLV
rsv38ZPc+TnWsnCECzHDG7T0MRfC/3plaBfsGwbUlN7Xk8aaPFQSkuyxR16BW2YZ
j6CeszE9OfYdZTYYeCcbm+OZngGjiS+jC94WzcKPDMlIeSFBipfG1Sd0O0oI3L68

//pragma protect end_data_block
//pragma protect digest_block
UTB1tc3VWStfWUYtuT+xuFhCkns=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
jB/szjAQB9bY5JDW7+148ep9NS/LFaoLmzWl0NOVw8DlDWz/1Z1LtbOIfWir4pmJ
lHzvcEVbL+jI1XM/zJSgTqOORqYKg1It+Bz09wJklZziepvyqf9X46lCilyLaYa4
+efXJjDWX5VpkUCMM+J1KyyuOwk7n+SiNxQwmb9AWvxgCSDhNd8slQ==
//pragma protect end_key_block
//pragma protect digest_block
WQoZtXCLtS5/gzJv6iLXdgXHL84=
//pragma protect end_digest_block
//pragma protect data_block
60wWq+nnZaDQ7sV8lr0RAGWNS3zDyIZn5Qe1yB2qNMh5HLPlSLcgVxNt9E8IeC+/
ZwjJIwu/nxx+yw3nkNCfkdMsKqzG6YhwWYOfHEq3Bbg/sd2dj/F4WD+GYrMWVGjS
LwsA+fuZClwlTn55N9qewnUcuLUM2sMjW1eqNOBJZGZ2v59KeewBahIZazcWcLNv
nuMtaLiOEHVkTWLtQu6szbO1RyVdzPHpCdc262ThCMiE4oXCxKuzVHiQm78zpO5Z
swgkxA5pAwkX0LTfLeEHrWZG4YahXXVWqcGpEaB6+R8Q+CzbSH0UEADGMsIPsNDz
RVUOmwixiRNyyZYDYPgPlgWqHIUtNcYWwJTTZzwMoDYuIZWye+Kj1J/lsxpHz4Oj
i17HeOObYYfEicibcIheU10/eGAo0r+eXxfI184CehYL82o0+ddFYWSrNvT+RhSB
+xM76RZyp867lrO1Am7pqp08zUginhtGaFnpZAxjKNlHpXLq9/FLjl/Ep37XxUMx
FvnzlSI8j5Qzfjgxqczou4aGInvlF+MPlD4Ftez0ELEsCkpv9x6hBZBArW2wdT6y
XMtXdAjjIqvxCG4HtMNUlHp2nY/jXgyDoGY+chMbvmzS6Ut1UJQJXFpMsYvQhLK9
35NqTBisO0YdCr1S9Ep6A2jd3RxaKw0QzNjy7/AeAJ2dQ2h4hLwgxMsUtskP0Yiw
/1lsdZ1a3I+kJxeByPezdBiYtWbq7HFG+gnmGpeZvZM5cMkyUFSUQIyahnMmqhps
LA9KPhAKIWL/3iVJgXCMgQvJ6hoM7L4xlNyt+3FjK5kqJf5AU1Zxl54kJdrrQXEF
p9H0OMqMM1Gi3oRmQ/j+M19ItitFsvPuUbrMrBjM44XNyCfrzKjY65GtOOGi8U7g
bplRshrymt7Y8Ze8cvG9jSMFfCjbkL8brKH5x69pjOC9ILEDdN5Y0+WXVRFJjdDu
UFtf2kwJlNCFC0wYAUUrCi9hsA7eqW4hrOXYvmAjSOOfLLHE9xG2GBt09OMHLp7J
U1iWST7Kk9g7kYSoSimJm3jNbq6wP3kcj7Em+b05BJffdzyt9KuRjyrhGV1sLhT4
p+1vl5bWuPClYAKy8r6cB8i3mitxngMQwu/QRyU8qeTkqpjLS+roizJDVQr7/xHs
g3mJtG+E+1OefD1a9EW4FtUKMfr9r+vzf7M4WX548FVISg7makqnuZjrME1cUNmD
1JzHgBSv6tCsJsuLrH7t6NR6BZDJ5QsdXcqjR7ALN97nkYpwDTKtgWYoCkGedCP3
0UOlyJFRXRruIP5bArU7MxI137esctO5gKdm+eVuNQdS9CXQhlkT/AQwc01SvkxT
adbvaclHaLeIBjUlCoqdCbJXCppj3Jb0HuEm2Oy6EYeBT4lD9zb+8MCJuIfTCPb2
BI58brS7S836nZRFbu21Pm8t8UQZAHTJTTcTjnLxgPCtl+kp38w2M8lQtIbiGWiu
IFRM8jQyCc5PKAEPOgCwtrLfJyoGz2onF7Z/OBeNS1vI2mF9zShTvFxqQKY5VBU9
1/Fs6Rp8AvrmnbZ3tGv9ern+Glsjw0fA4OAc4olIfK8dYgX0A9C5gsXLGyhfaUdc
6RLZAjvPCgR6dIh+YSXJXvV/iJ5OecSNzQc1BQXdnl4GtUsMQf47KIDsq1bY49KF
q/oyPZJQwR8vfC6ETb7JqFm5fOGjxU7/wlukftHLMVKTQl/d/e1kTHrBaCz3Npa7
59Jp5zvoZnasecENRBwzfthz1ubUFJ2+YKIqJAfD+P5kqLytPt6jj54508XhsLLF
TwDs8vUF/azEjMkZ5Evdez/whPTM5MGVdAinM+OUmEy+8JlyR3/VDGpaT5y/NZuz
w3QWtL5Yfkz/gMgguSDC44BiYot5/n1qzJYYvXCAISqzR68P4cYOU6AoO9NfcYrK
ZdwQjSQUdCcc1qfdYWrhu+cMmrllmtzMvCUQ2IRbD07s6Upf4D3/TLaHXOgOq9bK
y8XRhIjPiMY+sOkWetdvWVRA7Vx4wd//YdZD7R6SblaRHqxwHenu9w9IQ/u8rubP
hiveNJ3T9S1cP2WA/8aAj3k396R3F/L04H0UOo3C2Ow3NcATGfukK7W3f6CZadFm
XLLsvHe3zcr4QIGcgXTMJJCfzBHmd/o03fNmpGfanzHN9LgJDLrclTIq5XEXyuu9
pGDGvE101o2EJ9hPXCZInw6F7a+9d2gb/kHP0dHuJLMZFPjxh3YkpupS9IhaJ44W
+6gDooPsfKgi/+dFQnpE91EXV/tHxxlfcGuj45jzOU15Zy82yluWIzN6UAI55gYT
qVYBHDii3iE8M8oPxcFZciQYnEudUEscTi8jlAeBNKF7uSQkzB0whgmIehfabfCl
yrPTkxMBDp+FP/21cj5yDpJVSWJ46cfKYDYobRY8rG79/aktWuMQBeN0v40a567z
Rz2pmu0UMgY52UOsWzkKDDeh2qLNvDTcNOSbiEcpt1TwO1SfvwdnXzkfIeRUjPh+
9huBhu33GcNPeVvVn7p9Km5zCUXgjaVhDvHaQ5glOLNIUevz4FFwCRDR44bWLtD3
j61TfU312OIm+jOLqlbq1UZckzdF1x+vdAyuJ3oEy82HhlLSWHP0IRi65Ac1WkdA
PLTndg7PoxsyhWIzH0XQZoTcqOzYpW+5myDbYtA4IzWk0fwkQL+s7HxZw/scNYal
1AUOgZUEtBZwzScDlqdBz0vhLiUA1xr5a+49xDZarN9rfjqtHKCxx29skfKY42kE
hPd9j/kGbHM2rYjGApUSsW6zYGY6WBYrqiLUSVu8PWH7N0h5mzdMKKlV0084JOV/
M0A93msGw7C7krq4rOJNQD09EImItoNqTO2ix15ejr4st4gUj2YdTnm0zISK/zwe
+YrrkZjMzX95QPqQw6uEq493NhuKmGmj/z20yPVPcQix3aZr7iwih+4DqAKyp6gd
oZSJYMWB2p8EBxpuTsNCo+L5cduDHXjAmrpqTqJQ1NgmaBmqIFLQsdbI5vY8RJM6
1b0Bc+TPxm7j6vWJ27JZodJ/v/F46UZV7MhZsRwKP4VJxFvhJlUqFICbxtBAm/D6
FYG1CgxHGZT83SVOBO5UAiHluRUzcNirLTTubZn7C5ONmuzN//0LzUI0Fmw1gY9Q
L2MeQnH9nvQdIb3KlfJ1Us4at8B1o2sFu232z6b9yuTwnmxe6UgPWFR2iqEQzGvA
Yda3dxrbRuHciVEnPjdB8vTL1x9zVPDDOPh0yWITp7gOcastic5BzdKVTT8WDdtg
Ehnz5Okv8bTkC+uGfud8L65aMtMY2NzYYuKfdv7Yqi7H5pE4p3a+SOhjvvvlkqB/
jQi29WLZRHyXnsY4zUnt/FOjQbQ2cuvDEByona8H75xTe3ZXq5mn2GNsn/U6fATH
YCJXf/mZVcoUCtLS36mkZFKCtkpxBjZ6hBju9mUaOGzSMhD5I93Knxxs3F5H53hB
VA6J0AGq7r+0tOW5R5goNK1pyP9UxExCzgnDm14nP9io3ZmK/7JxHiTKpcPxNa5n
WKt0gauJYynqOnR6AaWwnvNHirGbo0bna1z4rnQxOrG/HvEX/eLB0VpXhLBxoqfJ
mXJQOnjObm1iFK3wj4MlG6RrbfxkYhqx97Z3o6uXw489C8HrBF1O+aHJDkQ8i16p
p43oLE074EhmufCotblEepLHVqEeufbGtJER7TCcUxVgG8yd2lOIEOxHdBHgbL7P
YKzortYIXVLGsFgx7CMe//i9BZqsTIp32s/UXAkXb6QoMZluWrASTkGdVNipRz5/
bKMx7LvRGwyedOsE7GE63gIFmFiiOuYA6KEvVj55ykN3eJNcuuDTlPfrOg6+qknl
tLLTHoEpn6MGAdZb28lF+Xul+kIwUpJ8+fJt0503b/0bdYNeJ8XoBk1CirVPK4u9
6xwdOWUQ6yaKPvIiBP/ix9Evl8IuiaosqYcFLJuLAgK3UWw9uZpTLlums8iDVrcv
5bKtITDZjjRFD2kTgGbIE+1SOh3lf0PQCKVIOjBDhCKCK01a+F2eO6Z3yNGzQu8a
FuaBeHF6pAFrgkVkEqtGXY1133DCHYSB6PQOLMebUkGIw6vjAPtBKpW4qZPixL1n
EPKVo350vZJkalQOAyLNbBAOQfujOmz6IYxxH1nt618lONfmJX2XTm+OTCnCyf1i
aD26uYCN6Ch1OxRZO/7X1H8JtqgnNSxCFGp8W04sOlZR+50c/GNw+xQTBz7GaQfI
y36ulbM7hWoMnjQORekXKB8ZEHiQZtBF7odRK7B00Z4nOhBHtaQIqEuI8BMskILb
WCiIuvj2sKcLCEtYt+FA58PiW6ZbB9ZwP6XnlBJmP/EY8kpiahZUrg/X4TsCxZfV
G6OnpswHRauYlQ24xuEMWmaJdbBFUOaNYcaLh+RGH35WQSHhMcJmOR2Nx7/cHHuu
BHdzRLRzEavQKPcW6CBejXKLNr4k/vl2JadXcDyFDoaPGjQ+8ZCm1liEIL5nnS14
beq5prxDLdoxNM1OrdLVA7o8EJ/qiXQrEqLLc1EL2Xs4rSYxQd0KUgcXG8Q8OwLi
OlrvRnWjlhe8YmFoEJO1cBMWbQTlAr0PR9aMtkeBqQ/5YKZJqtkgxb018A7oj7vU
udFQBB4r9qsA0mUMbCrixoQC7TtZsRUoRan/grWnwnzSO72flqcLF6xF79rZLbh5
khlBBFwj5RX3TJ8wKxf0OEiEJi++VpnjCOln1Y6uZNU592cjDgomuVe4YIir86mB
OcaeOjRPxy8csP9VauBJEmLWfHEDdkEHhBSge5ICqBPcRX7YVq8xbHDxm4DjQ1Bk
3xJExTnYmhbkOJIWaZvEJ1E18p8GPnDATJlN5k5mDPZqV0GFQGQFxEUL1+0uh61q
Cge2z2apLNORokPGZT0qRtmRaJ9x0ftyaYMcQcaS1nbKwSd6GBFPKhHna2aDzCWu
ed37wnOy9f3fMehk0n3qriAKutciD3ZMJRIEIXfOGbd3w7ybdyU/3ROqfwLMuL3I
Uka/LkzFBPkVpMmFF47dohS01rg0IGnU9O3Fj297KtEAyN0tKXJuXvLOri9VGPx0
/W20eX8lG3vTGQkH7PWAt0RuZ5n7vV3FjGRJEcVEhH0eIsI0Yy7Zezm0xDb5l/bB
Md+chwgSIg8qaUbLBDMwLUktVePaVtoz9GJNreXbELoT2yD1pSigBRgrf1prhM5b
l6erS6NR2Yy0PIzzT/g5k0Jc7ZXluYg6lPkr3aV2Jn3hhVu21GcPjOXhZ2wvqR5a
x11X+30veSkbOajIYEXD46+Wp9Ty++VcQ3TGhgJSI1YhZaAYb/nWC7RHZATb3u3v
rwPnKAfBlwQGnrFmuEn7FTa1emOAbBFm+CcgAbrF9T6yI14Xn40+iV4OPJUQcdvW
0aL0rGBfCujRpzmQ12th/DqyZk6L3y7dMjvH9pJwZuMjLZ5c/KzJdm+f1purSi1U
ipLs1z6p0TOy0/EikTYpC871yapPHneOG4lwqm7xCB5+Uy9LR0wUQE72gR3q30PY
x6/jDwvIsGcrUAPsxojtQP3Na73Rf4VU885mbz8aSvoZ0o6l8+fIjrXhILVZL2XV
EyfhMKD+MRUeZZPFg6iMcGInDO2z4xRiLLP+4O8JWGMzEOOUK1eq3brCIkmclBLM
y1DCO2IitaGIYxWvC1WSM4FJlzEQRn7V78uh1mPL0pgCIHIVzfjnFHpPA0HsRunQ
rQH8v285R4+JHd8TEemsrVM7dRNYWL221D1vzecahJ1tZcH3BNjqUb1aiJ6eS4kt
aWCAoWGlbx87Xyao95q3KvR7ejEPEkAFYzqYJpNzANHDvr80/5wOS9DnHTIaleOn
XM9FpS0XlBF3DRvzT1OiYSZoHdkWlRbUkAZZSu4dLdlsJPEa+5NDxd1ovC0RyaR/
ZV/XwPCujgGTAWUrUt4JRAhBaEcb4QoHx+C/HtxoR8QOzn0ExqqFVHo0uvBBrqYI
Ua4ap2+/5nCHwfT0fXr8z9aPmWNVMHFH2gs9B83mRiRvLmPQYdEXIgB3nAF457B9
qSGougTswzchrbWxmkCl1ASXDsBNuETyBmf1w2baAwYNvsVE6diirFpl51YXZT2Z
TMKfPP4pH61wkbqE4JPiWUNhEJUKUajYyLH4iGlLNIOkqJAxRYT2Lo2ymHRSy5z9
buMSjC7YINIoPXDdrl5pg1o/J2ZxyQ5GvOjzzqgGgbt3uDNvy4qAHg0A9LVcWubW
TIZzd3TscpSMLepcvv4c2Mc2on+o9BN9UiMndKtOY2smQN+IVmIz+cMiCexig7Nf
e0RaFqfUwQuaOU9fbBZwqrOoqCWFD5fpcTf6L23/Nr3ugbgDK8Z1HLhpLYdu54Qb
bgiKlqFe+boTl1EY15z+lCRubSy4nB7YQgfTBXWcPZP+H5Eb9lJh1Xj9hrhtHO7h
jZNl9KuhpKfczb0Gyk7UCwYbxK6LFcQT1ACpmtx0xNhLeY9rg7RDf+xCW6OBTcoC
7lLgpQxvrjxfdEWg0f8+Ln0F6qZobmygaOjlL865kz+aDW39vywHYsQVAb01wWi/
MiJPprgg/7jOn/osKR3rDSHmzPru6hC5BOkNccK32hc4YJZHhqBo5QNdbEaY6BQZ
j55P421OYlY+7qHxLP4ecAYjtcNqHZNnWX2WfTxAIHl4GDBsZE94OW5hKegqgX+u
gQifivjox1EF/B/qB4r/GLombOfq6wXclQlSpnmVQohyejVBR1P8pQi9rvNx8nw5
2nup9vmokhwNMoa5oW8uxn9EsVqAfCxLajnUZhQh9ecq0P905Z2rUDJwsnhTjNQ3
buwKa11vn0Wx20Rrjgqttm8nl6C+Im+daWQNQs8R1A51V4le8alASz8UEfSoA++L
YlTICJqOfTf786D3gaWCeu2c2lviRSn8O7HDRqitPJWk45hFtg/pp0zDKfBUq+4e
2ldcmd7C0DeFop1r86umdPiFGg2Bd8DbNxnLkd8UihUdhc6S7WfMVGZqAL46+bgI
GP2aiALBimQtctPwqbEqdvwTZSVNhTdELvhpy+YoQZfZ7noOCzebYOX5w82y1mbM
fwqjkKBhpJOoCg60otKfFDOof77x2cV/JzeXZDTa04md0cxHOZSpmGoTvcA9SPYa
+cmUiyEZ2jzagTuZo9FizfTsa2wFbeA5UfwY4K51/kPwgmRxTmZECNoUpkBZplG6
fVpshQy4DokJpjutFwhSFf+Qn1UrDxAg4CTDoyHzqCisFLko6sGgVDmumsw7R8Et
psOfrPBQaOe2an4QCzVSIhQaFvsGE8EgLFtFSquVcRO4xOcBt7cvzBhW5Iw/OOpj
Rs0eFCiCrX9iS5URpcusupaJ2VhYJm/jmvbJVuAKdfdK6HxGkbYrsSzA3AS1qYHM
10FZm7L/WryzJdGxwIXFXRUsX9eLQJ7pGttYwZ7pQpFLZLEvaO9Nzvj5seLPrFol
j9wGVCzs8/vhT27LFOZVqc7qai7nyZ+g93vy+W5biDBSsZV2to9eWO99YUVHwzpt
BRV+E6L1gprn6lKbWdjrlB0eiyXMlNHqIaEj3eHSdSidGBx6d7IeqgAjqTtV72PC
cmYZa4rR+EkM2WHNCqSpkU3BFSyN6sca6Xtrqp+2d9d6oHdhVroDH08Ps4Djgj9h
xToGCY4jV5Yt2ZXM14/ZzGp8kp2v0hUDan+oWgJZLejoohiiQ7l0snd46FEXv7bT
LdGNpmdOIx7q24KTE/VBPvkEE2BU7WmSL2DklIdb1bSLmFf2RRtRc869E/6T3qxy
7H9y8aRapjJyeQZa+nqIg5Or52EXeI+s4GR9718Jfc38fY1PRbNdfrpxDP116xxs
BzjMdZKorwNr/kpGswF4TJ91zSzWYQbtUbcRScVOXTmnblDapDi7OLSJ74M3rQAt
hhWkhEIYmvo2dgHUqYt+3L1ghRaCR5RtqcFiAvCjTTR0/c4U4HsmMCU0pcwRfCf1
bvRBtwNJWGcYZrmxfqXrXUPr66T8ObVFcB6varwJf2Z2id4sybs1CS9GcPzXCUO0
0+zo1M7qmrG1zFdXnoX5PQXqV2gABCwBwR8ngr6BU6j82tkdQ0UPqBUWlj0of4qG
c2r0q1dtGKffkY/iJHFY+zTMsduq5xrOWislXmz5+DLYaJeCFDb8+OKpebpT1fj/
cc8Y1bpPMFdtmnqd64vgYYq8ql2L1dkNf7FV2HgbRxLXnqb+WKKDDrxH7H8gaR1D
9ltkRJALyjf5mLyFbPg+cmmzSEutP7iYKcxxtG3c+9J2/6oXG/tWyV/UGvJuQCvl
Lb1p3S8XCQGSzs0sjAZ5dDC3sOdYE0llgPqG74ICvGncofKSDfhvbaWZ2Q/s4Keg
JFY865g9KKv9IvTs6RQftK4JbT9fl+bkTznEEGGctfvkKM7TTu1/y+LSGgJ4Gh1s
VNXHyrMHvaafpH7F3UTugUo0+yAGuXoI6AKMCYq2QFpol4cdvP4kwu7qOsNrvhYq
IbdI4Je/cNN27rBfTSLUSxzZR51KTGwAuHN4ZoJfup//Sj8eUeTMtpijy7CABuSv
PRvrneUafOmY2FGamEHTq+RwezhRbrCihb9UxgzgpSo/y788Af1FCcztIOQ/5WEx
516X4KN088DbzaKTtrG9+LcG7DhqzUrXu0QV63gL7H2ighA3hOQzOto9ZJ+Y7kUd
CFRzaAhOA8ahwaXKzfFU1ilAVmSyXOQMfSlV+o5G5PyXoilvQJEpZuesjXLltJ4B
BHPlPzzZZjkPQ29NRXVzrQCYciECQIZfG8t5HNEY8I1bBiPVk8zlSzLd9xm3goY4
4y3A/NCE81UClgMCizT9ABDRi8WXYPf+6Na8gPnxow0sawYlu1h10rxzuHqMMQsd
BJZ9F32JY63+Cxc+3vmkDbI1uo4LcpuGlWovml4Slk+DFb9ktLvYKJXReJICVTzT
N0OmhCZyA2Ge69maUuVWieW23gtVzJtLY60DXsEP5KWPDwmOT1Jb3CBB3dK0+IpP
/r6U4ME75Yt//+sc9gNV8Pn2GrZo421B3CaxaD9RlYZSIzIB3B2/NGOwksuin8jX
jhuX5Jdpgri8YWDPyFM8ackQeMe1quAPZ/nB6SRcd/MjXTxwBD8OiWZRmqC6Sixo
HQRwpUUK4Q7kAD6RuI5PpMfMgMeYrCN3h1a1o0N4+qHsqeOa6Wc0LuxRL0P+7Kd1
kC71iacNYzyzfgPTo/l6PRCKwPBdU1UfHjyZhyzMLF9mSVh5vEvkVVq5FmYzBgHL
W2jhe8q/eMSj5eeQWtS0GQlAlq9EHQ9/Y7mbWvR5AqeLBCSIff4sfKzYp9iuZIm+
M9SaY72Saf0CjaiJ7/8PjMqZIHN7BBvZZXRpGgTcYv31jjNSZtIf9VwJm6HBb8jc
ZZa9sbG77lk2fNwmAzNrN7u6iXxnRot+826Ny3w0Pe/K4yAGaG+kaZHRzXbEkhsS
t8zLLFfgPtVS6kWwC/KB/w5KxRQWa6K8NRjG1ykcFYmJVB7OYqbSJLizcJ97KSrN
//aBl/pUuy4S3IzKeEF/Xqa6x6bdXSI9iqxeQxXJ+dXBKj3GNplRXMNRvCVzK4pM
3iDKvApuBNAlV3CItRS9F7BjG62P69Fk0j8mGzqopYgS85IfmxHM4ivBqlLVAgSM
29Lr2QY2WThfeC4NoPd3j9nl3UuNby7D7dXNPlL1o+ALB2tFHejmtqMgiL/x7RQZ
3QBQ3jDDOcy0dgpupzXS3Ll6Ix5TAdsbLIdKx3v2c7U7mbzMxC3su1UnklEXr02e
gxHoyhiHLXZuEh6Ht8unxNIDRTRzQs5L9Mov90U6VOBzpergQ2raUNBuR3kwMP1a
zbcyMHAW8J531J+uv6zxNoCE8QSXWlN1HUtcT2RusgYvA2whYp6okttGyzq8O2zi
1NQOH9R8RIWSGYBE2p1+66e0GUKkpJi0+Kn6UZuLJ03iMjIKrVZxH6tyDuoDLIak
e+P6bw1gSpLSP+i2Wj88ofm+g1RSzA5giNcPW1ExsemMkesq2eOBv9Ii8XSiSuNh
mZE276CzLd9TSr21uRsEfWpB1yneNJRqaupjt803gwBC4Z/ug41ClgC/PUCxszCf
W0Di/mlJCoMH0MUl0bJuM7b/9CjhYnKDtv2dOQ+l74pDO5yTkQhJGwqPrZkRuPcG
eBtq2Ydc+vfwaywUepsKkOhXs8NdQGNE0pwfaGQVkr/nT+BHot8lh3vp/dS4eahh
Y9CDmuYJxSLxHPsTn2jCJ/5vbo4P5bisJK99Rdup6t/cHqneF5ohw886VJdB2I/M
tsvVwKq/6M5dbm8zI3m07YqwtuMR+p2G2w5KINyeUSSub5KKjzc4rJgq+41kWEpy
CLyy/yvqnJeq4pltuit5+kcwFvVaFmQO/sV0gQKseLnpM0oQpeXv9Lfz5jBaxRP9
cPikyGthQNvToZU0t2/TxwtHPg9Pm8uH9RbdELfWaioYDdNQDw1oFEYhWGVuZKWm
bG6UA4UHq1dk2qgn59Mmho8H+H3v2l41V0NY7VpENnhHYLmi5fSq6tD7HLnP7hJa
1Xuc6f4d+jxbx65IcV1cl3tMKshRsDqJsQZEt0SOEP8Yz3DHE6eb1Rb3IxUTVB72
Pl7EccHdsYGDLbws/PNTksi6DVfX3RtEhdSxJHIwHGbeRjRjl1ENThzw4/Jgas8f
OikFKlFopMa1Kvknzt+Og8K2SxU6yRrMnRqldMFkKJYUuHpTV3kNXTMZStUDXj0M
G50cvCdG50aEzSZDo/z60Zc2QU9vS6Ij/pKs/bzXk7dBzlZmb2HzdS5SgG/0BFGq
wMPADiPZEsqX/wI6z8Fr4uX2+0UlN+QNyebWmGlsjFL2BWbOE4aprA4HNWCP2Mb1
unWU/+gkDziS8EyM8RAXSCcGBeHF5D3IvPGi5x4ii92UGiVrf66fEa8oiKFfvzep
+aAyePAqGQUl/9yXLPfPwa+P7SCskSgFrMd8o5TKuHClfUsi6kflkXckZHOVCbtH
nrh77jHhgOhyzR2GunJi7KVPd+HUPY3ZPWSf4SbSVSLjSH2LT+5Md0zBip5RwgfX
J+5Lrg9PB13ClBneheq7ieQnJabA2THyenIJy9aafTtKE1elEP5F3nAT6M36NErR
wAokDNpoWXB4AVllLAt95+Veuoi0LQAvHyWeeUPZIYN+5P4mbrIVB+af0BqI8Cma
XBRQEtiwt1suj0HQ5MCLf45ase5aSonvD0Hk4BKsy17Wagvdsr3fH4a+Eo6KlBoS
om0rpGjBDSsDWPzZ64p+e37Rp154YJRHpPIkHLNMTPGr2H5Zbb0j9ElqO2zQDLAP
imrHXnDhrdHblKU5hwE89GiYrXL7EqRLhI0vaHUe4YIxb3lF7D/D9/l1PrXKIWXv
aGoshpgCcUHZNIN1weooqBee1qmxb8laOanUsDJsa747mfsIUx+MKmA/4UpiLSgp
9JTMzCthZPT4glZvjCrWeJ0ZVb6hKTwC4j8QHuEB6dsrEIujWnXG3dcDxclk9iDN
nBV1mLdj0XQNz6nG+0HsxmUt9sbt/pzuZr6tzk0gAhRbGiOK+/Y0mzvewzQOBe4S
ehKn8mLSMDtT3NEEfStvh80B4bKP1AcLneOmaG8irloZrkW+52WvNq/DRbnODNlf
mkhA35U1+8B85PyTJSmkRScl/1cQdodNPeAWmSCwftuEU+TbkW6otjvgeHYLmZ/u
cN2GnR40/A4AcnWu7aP4MNtCKbZfTcze7Vq8bj96lesEGNEjQNv0exJ4hxTyPGBG
CY4Hh9dLUOyXjmSb01dczYKPPtGsdsRo7CsIdOQXY4KrJQGr02TU2Xusah/jcNaJ
RCReLAuIbv4ya1o2vl1CQPxa1Mkqo6Q9GA+brRLmdDRG+MfLR7Wr3oSG5OUxP3wB
AaPIhzCcNPAJjbpr0/v1JrwkqS0uSnCkVFkhraqPf7fb6Hw9OTiFbdZkYuc5eFXR
L4kW7VOq+oC7he99S6TSG0tw73wonr8QOkIMqLvHTWxlV8EnStCXgGnQtM/IjoKI
+wr6CSKCOYK1k0W5j50dWxpJ6roJjQVkuqJObpHV4KErxXpBq84vU62NT/uGYDN8
7NXjPg34hIEUGVvb9iY7iiGiLyyqWqC0Lgtede+JN9fVj36FMCLYxRxVc5xH9afP
U0n+Cp85P5mMabapBefNmgIUcIlgO5YPSW0mVKQofwULaTnVPl69zEo+2wj81HuZ
KS3BbPDDRqds9BAQnMqZ4l6VHnm/zBWe88HWTebBterXl0mr9WVcUaw+CwKbYQUF
N+xwlkjyaSGE640qXxrYV3SV1E3LPKjNgfyiiX1oJslSBAK1wqHFcwZqBh8OQIQy
g1juTl4kb5WoqSDCSvC+XSdOhfvLcR0S6cybf/iMUIQK6+otxx92vMr1/uhsQ1MP
881xGIJSP5gyp1c+d3tiCH0y4tpbDp674TNJTjqmuRXVvkGRArWeEkUzNdNO4bh9
tXcGD1KmPI70bhNRpYVfNm8lM2TayG0QsjYzz5GUGBHSbumo5SmsjUstwQzWQ062
P4Y626s4/2fe6T9Du7RTpVCOGntzRpQj1KkfaZvdYK989HsMVjS3JqbXtWgJO6Bw
wGoVKDu2duxWLY+xMTLsFUIxkqwEoOk1VBzOFEUZSJ1MdP3p+6oKSXRviSrtX95t
P4zoccrFEBoP1/geE2KnWoIWcUTVvyGHo5TdQMMHQ4dXDU585tjm6b/kYlHf7xCG
EvgEQOsJRn0VZ9xLqCDPPLY2xKXmGVD1VGG9lqO2JIGGRpLSA0sOOI7CnN0GlTD1
yq6ySMfNT/iJe3vrL2TcxwpCa3uk5bie6giyRkx6CVEVmzs0h83GkH5dHLRdRIOb
1lUKZItsBEB9iqO19T/B8ZVYEByNR9ke47tM+3iLNr2D64HHvO0h4DklhhAV8BqO
k6JwSxqQ6Xpa10j8N4eDQE1OAupUcNeGIMxR1hHbHomnTbJAknaK3XbW8mdWdQ9o
nX1wmOsCXsF88lxfWxxP8lzL0KyXHCjsIrjaVSb/70IPXjkqnjxv3dDYENbcxUAF
dtPec4lyLKejO/ncRUDt0PqatKZ5x3pPCchkZYXnsPpBV+gTOKclHmSYQsvbcRSd
OopRwzPkYC3O9ZosM7K8u9BFWlCgyW67FbhtkKo2oOwJFI4QuZDDb0dgAoBMyPDi
SnTn52jE/H6v/BNTdlg+eoODf0NhLPswyt8X0C7F4VStsYXFEgrW7vby+htoEGZo
EL2NtigXP5ZP/ouFQBLRYZXNVCxXdQDbgKGrBUZAXeD7tAO3aXhvzb6w5+bYeHWi
JwOkzHLVvYmV0xk4F2MWnNMdpyapZLkz4rpqWLuhgPdxSjBVQGeGIYR+0Z2SWXeK
lciyukfKWn0OBwisBTz7u1sdDkJ52V5MzYDR1LNiKm47jStxveb/k1eJAS2Gy5jH
VeC8D92H9M28QMxEJ/6ogeiCGHqtnIY6u9KuECx+vTa+yr14C0UTtCvG+SfS+Zoc
JsV1nG4COr3JqAeRzaq4Sdsad/SluAoIhGe3Bs8syRATqkrRsDz3xlrvu+St/avY
in/Gt63/jjyHHCOakcojqy5QP34gr5pJebJeHf6QMyMq/va545vlt4bJVzw0N3cH
0eLNETm67w2UXmRC6fVPwmowUszmFyc+QhRE0ynJyvAPAUNGqibIDMh73bcqs2yN
WPMHruKbhfLw3hHW+j02M2VIAQOLUwTzVzm8zO8B5i8JHEDKfq+pt3RHu/AIeCGb
5Sb992aAGmm0pXpQd2WVycfB/qWsWt143tp9aoIG+iU7ZLv5ooXllFk4qQ8Q9vdI
7KDBsUlvl6d/dC7Ss0B2QACFabw4FGqCAy+SMephYVBn9l9clrP6H+ZFNiXC6zGY
0C0qbkKWQCEmVJa9XfLuHirZI1ghFkOdDQl2TBCt8b+PRIl25US4O53qUJsw/LWK
tKiGLLawfA6Kc8DtzykLMzrTrbKia8JGr5RrByAndLJudOFiwQW2JKraDRx/k2ij
EUdHBbGY+3DHLG7vOIjup28C7nl6uAasqNxXx9NqiJ3j0JaBnhCJ3GRLssLSJ5yg
pquWMMhtBZPH9T0RHTJ5gs4THqzi3i4Xqyb3/fv7bkfL6YUYzckhp2xZfnIDfRn7
pSWMvvBihscriAE7G7clKJvEaOR6IsK4gX10GTdxU5luHO+pfIdWzX55Q4YQE59u
7mfE5Et/Z+Jh7QD3w8MIgclDg3MxAG0J8do/AzHO3DZZzw8IujARSfQT11XjgBDd
DaTtgHmIjGEYJD9xJshgow3yyFNXgOgMbMSa8xbJoNPbxHm5EF9CfTbHvBNAxsHJ
SkIyv6nGVZXrh/IHOQEafWidwXNGdVHeLc9Dh9LAZS+sgoW+CRIu0Ed0TewyMJiK
kmSvSKKWuIeRZEm81RnaPzBypxh9tzg98zDktsq09QhxNh2F0cMFu+2kxZxbZDdS
F6OpyAz1MLrN6OupOYR8gdvL6gYPH1MV1R8hKvRhQ9y4ZX6uygkYSaJELEwh1l13
jfpFRB9wDmMEMeCePXYEb+jthoRgEz5g8RM3e8fTaYA28aEa908rZklylkXzRc/i
6fW3wM1aW1Wtuz0tzKHIMMQiLg53v5mYVokWoe52eG/DWu1f8tenaXX8O+2CeWF+
LHH8CGUUqdx/xKA1K/otrXuSKEAt6X3I3bAwOyT0AWtI8eJd3xXoXJBJZDqgX/cZ
a3FA/TYmqYZghWyPo7nh+3KloyH7bp/fWn4K7YR18p74BXeSPAwCXNUpOK9V3zoV
Y914dJduoh7pqNyKCRy7jbEs/iLzzYN6uxjQFSGkN8s335SdGVYjKjTvDbLwcsQ8
gTccUNex5ATQ/4xQO/QpUgkkqJjyLDMPRCD3BeprYMnu7W+c2SSNqi90HsCKunux
iSFe/9gjvEGewiAxbzP+1PI2yuziVXnt213Jr3+Na4tA3o2hoYVAHPQdybfXUEhk
CF5B2EGKBA49BRXxED4lWeEyLzOMvQ7sMILyrT3n/oPKzyXpWP3aXiHJ0qh7/SsS
c4cX6XzjM30BAArPhuOvebe17b16kVVsDGmT/oDwXdSWlZfiayeLR1hFdTISOPgw
K/Nk1xboaVe4IvnFLcwxGCM8+Y2mlkUdPiVSuUWPPZNL0n8r9yayKIK5OniH+kR6
ixQW6zQ84uhOB+RpLUylEw0PT6phrjfz28yeJFCEuHHJgmhY8XSDV45OSisq7zd3
bzAWXQdaW66Fj5TPdyVNNpC20/udTvS4zr0nSENbgcWk4n0uYXrBpL5qMUIVJfCJ
h/d4x8FXWUaHaPa2cW9QOI8W/nNu1U7+P2bk1bu0keD/EQlG/LwJX+H+DNaN5Mby
TXDUVG6Eu/O0QcHS5v3XttM+QunavHanRwxbywRjFZugw26DK0+FTuxhuva1CqRX
cBAXOGVZRc38T+WCO/1rZAK/o57p6N8rVnTR+MDkU1eo+yzNJZWkWA7G7kZuz8Nz
tjuKiXcqr366MYTTYSGznc8Jpl9tkL6jZFjkKo8lg20gisnpM1MkNLHZNpSafJYl
DhTQHJnO/OJARuhS0esI/wXNs06VpOxg9G90hkUOANwjOTUdt04DCbdA85OYws3d
qRgz76gqObuA4K21IgqkgOrv8V0Z53yLtz1CJVoZzxVb78NPtslciWznAmJFmAsb
fqXAxW2mHn9aHE3OG+99iw00khp7h9fj8I4WiTWiPz760XJiiYDYW5B+GjCU/2cV
d+Hiyo6g+c7rU8RAjv/rPnOPBL55Hn8xfkcWkr3QI2nYkpTL/nOXihvFZZ3LXQfp
J4L281vNILxtAWSLa/UBk5T7VZlv0h0sG0vDIn4pRi/uIyM6N+ZJud+l4ly5AXcO
MiOUoPC3WN25tWENUiQR9Lh9TtyOO43yfncuc5REizhQrwh7hc2IU3VP9BOYcPVM
iFJZKCTdmVibM/wGH/HlbjDNeRQUzxI2PVokGl6GRidp0PjqTRjLhDrRFU8u4gCg
atUHtSGbzZksaFsBnCvRUZAzDdESkRU3M9q7gGDSdr2HhnyL/Snfy/3aoWqBahsW
h4lylB5EJ177nGH2BrzKjbJic3XJzpBDt0tCtb+r8VtAS9I1yJZGkWA9/KSXgPXQ
JEmdJrXe4D1iQrdAP5OcPf+yx57BRTB6fpbEsPpdDER6piM2cQ80qA0DPs+MN5fj
MI9Yep6O5NbQeJsaW0q6cOcaO8CXmbmIsxFPFesrRwJm91vRaMZNm2HwKzoEnGTy
19TDL89fEInUZQX5jnseCkJXh/AQqZLdATNoHRxvW1et9JSOOV+8tGe6Cdp2sNd0
7rpNlZ48KRyhzUeiTIRbrWah7UjmjmxVw04U9SNEhNZYb4YNsmXyPEx66WUnHW7b
sncqrWDGL4ARHb6LXnoGbm7XtCZkRYi6hWQlLbKIvKBnwFs6j5f7HYhbW8QJLieq
7CxDS1wm8VzXMtoPVm8oNbTPEMNJbqBAq09H306wGIPlihU5Gil9Z4rEBJj6BGNH
GiIMPYoYFXeiosZpcbrhh+vZPcT5XUdmy9rJ14pzBwA8gRv43ZbuQa3Fh1hvnUBZ
X88oqmn8qd7u5pHkTi7DJDTEFE9TRQjLew0194z3EJ3ebvjIiQ/Cj/Hf8PYeMVGc
4Mgy1cDcRU10oTf6V0aVRFEkULPKNTr9aFrqrFiz3Z1952Wy686vEWGNe2I9TgUg
BykXAA4F3LEGh4DH3p9sf5HJ3MJng0duFZnnPCyNoXMy99rUU0BzJjex+Pag1p+E
hts6SwjALmpqeNLOVRdN8UNT4/hylmfMJiUKF6w5JUgNAwLfMmjGbpJkz04hSJ1d
wViyq7rARdL2K9PHkftNntRTJa2IBAUFOs0NbGooTwLnTRlRHI190OBMMlzspgFw
U70zORQMWTDjI37UleFTI5PYjHt6phpGtZ+Kv1BVWyd3RGdkP5YG/nfiK1qCwqXN
18JJxhNZB2vmPMiL7NMyKOj6/1Xm2keOEYd+pTlYXbNAz95NZBMQ+3dJAdzN8iaD
6LQJaqY/K8nCYn3BzRtnUXsm/Xc9vgr6IztyPu2Z2IJMMopbF9nB2ABlX5zxeeGO
Jqai707gXLg7ZpkscwjoChnnRwN4W0LNtSErZpEV2vReskSLIsk1Te1QtpyvN8ne
1x+kG9UWOma19lGAEDKszOIyBjQy8VI1rr+Z5zEWMGx/sD1ssZAraU5dDwCtIMcx
WBKtilTK0R40F8xlTW68ELDHFKt5Wcq22qd2Z4X3sFqykJ8Mr6npjdyVuIg6bQZP
vP79FXKJFLjEQXmZJi8C4pXu8UXtULObMTug5YH/yFnJPI4Rj3wzgp3UDp3gIWxT
uOrz34DIDQRCwceIZKWjA171m+DLs6mXVwXRsYxempcNzUYOsC3yT2kMr4xqzazM
YQfWSite6dhZTMAe6gcuONBvA9e/YP0KXUZHX9CAq/UXwyZ4x6f3S101ATIuqv1Z
rBTF63rS5I6ee0CDaL1qvKpw2yZl2EyB1o16qGwV1R+pmNG7c6ddvK1FCkHeURGc
nHFVmj9kc5a1b/po7puRG8cT5K2BmkH8simVFhN57ZjIN3B7/pxsQvCRuTeg1cpR
ozksogXnhVTa3QCFwnti9Iq7q60GW0Y4BICSG+oFI+aJS5tnkcZEWXZpcTUkVBcU
8qhYkxvD/APGgyu81A55WdAYuSuE1j/jXqkjHV+MrnFaG0H3z9SHnrLCbWZdIzlT
c9nK8UUEStWeFnoPs77L1/f+cbhe+Io/Thh2xKxOoXjc3QG6so7NEzhN05xOVY4e
zfiVWjUIp8Nh3x00mqudhE3WDx1gsL2//zHGlva6MMc2tdBvnb+pT5padSGNLO36
+zF1pCpiPxKTbEllibpjOX3xIuZjqjqfU2kfa2T/C4UztCWcwYkMl6KgkixOW73n
1LaAYV6y+pXHlV4WgzO9rMoyccHY5ip/hOx/fL2tAutsmmoUig00+JukjuBXrPem
ajjmx1K3msehM8T9T/whm5twbziBz8yVskKzv/aatZ1n83Og2vOSLNJJB+Nlt3e0
iKUTr+0jAMTmcEF4T9tGKsU75zPxbT4mUUNdsdcc9Q88yGgtYkd01OwIIn8yikLL
RNQ8ImjbCsRWDA7Mf/0VOfCWnNVqvMqqXSjH6Y9rvTe4crpzLVAU9vJJPXrbWekT
xh18irJ6YOzwXkMbhtm4FcTO4oTyzSijBtAFg6riNyff8Z5hXFLKqVet1scEKgGG
RX3GwL4jcMf+ZyuHTbWpB/fLlXmwgRlIDIGSiAEXMRJo6jLorprwVxOM/2hTuK3d
MmzPRDmOQjGXrOVK0sDFjTpv9UdXWFy381Gxxw/DEJLuZaxVMbRfRigGG+HflSgu
3eE8hr1HQOamIQYM4Nu2Q2ieMOfplExcIipMPi0FCfMK/SoonGWF2dwIg/CN+LKJ
KhfwM75zojAhe5PA2pj16cXZc5sQFd7CupbUkrNewrKIG2cNKR92iFl6+C9m9coY
QsI4m+4P+xqnRZzAQjrUxt+RXLh4Cpqc9OVNa9jbK5xkL8z8vwkHzclAW12qwSx+
dx6bJ3mTcI6AWbVapg9fzlrIli99gn3rEXUXFbnSRlNiJfjW2oYBt1gqtsu4vYEL
tx0ypXehGkN96ggqapevc6W6Gq30t5LPygCSVz69ZzK/tIokhxIefG8VbXHDmbwV
10pBS7q/gUkXFh0vFnXhAIxbT0fG/QzezU1EAFqcadGUYdcMalpE6kxSsshkSZvF
rRR/ylH11oSuS58K912VYXfy11pxwBvKh9BGh0PppzCuWUQHrp5nCG+gGHCCRAmG
pzMYL3SkuQnG/dRQ/cZDuyScDkInzwHj6WWv66mQbNX5tM3ECDKC61f37KoTHEwF
RqyNcMvNeDAC5uwdiXiaZPo71/nU4gpj/UePmUtqosXs46MPfdR92PKrJlQQ86ny
0GmBh/s98kEhmFLERi7r5Ohawg+fVFBLoGPkQA3w4gTe26KJgj86Eux+upGKSNLo
B9/9z+0wOrDd98q6civ58aSpTCnvB17MQFD9Ieg/CKhl0a3ejkikd4ZLJQSqi87G
kCR0YwKzoroJyStxL3zXe/qfORzc5cVhOGDBo13rYwzE/Ao5GKkNSY8egsgteRCF
qJ3THIuwbbwD6y8qAkB5GJermRBYvsgWguyFEbjUMNjjqOY1sNPFpZvP/Kbu6Lp2
HmEXsb4lAI1pxJRNk3QW3N2QfFGFcJSHMwpYp5GNSL4uPkK73bWIobwSpnv7nEmI
VJUVWdJ02k9WcxwJ49kxsdUtOFr/Os7iA1EClDsc7/c8JW61ti6CeJAJvR8C0ApG
1AY4K07J/+DtWdhgzhZOPQzny+5lj1tnLfOet4chXiLynQkX7NKrRXB/1nkcUDRo
FgeN4DEqPqhSfEWc9sBtnQhOIMOoi6oQPDCGrbYoI9D+BNgfdHmGLLs/zwibIHfv
IGstkqSUZc7Eiazew86Yz9qOOqaLRbs4Vkpez7DDU2UvFhK5RVY7x888+ybXWBtS
FzO0H8KTyVJL+cSUl14kb+V5uJsEy/0ZPISUjOPO91huxD5GKgLBDKObKWO5c+H2
+qINAtK0wXoZjIm1hlN7B9YV2m2SVQoanO+PvKojl0GxcuzBVH8nsxmz/garGlnv
YtMDTMQsCOA2LJ6ZOMaelyYqDeAaQOQOinS6+NlYYhgEfQd8sSw7v8ypvYpFuEwc
4PfmD7tNVaQeTg5S31nF6O1QESC5xNLggZf2obbSdKqvPBkHc4FBZZmko17Z4+FI
Nj0GX6TaSMQUr4105ZIKBjpGkkq7nzhy1rQjr7VdsmmbFr63WMju7J/VYOjWarvd
DZTDAjiBK7QUEJil9LS0KN3VUxHPCMrtVICD7YgqgikXevN86SKDA2EvGZ8tTYCi
KKs9UBrbvHPTajyLRsjYjto/I735wH6G7ZMwxuIjXiVn9x1PGpSlLOr7uV6tIrHx
jkB/QG6JXDfvJELoL+yMVP+LAna8Wj+/s42Y2jNVWqDBu/nv60mFKR+RABUSf0Zz
L6C9oIsx6KUc6PSlKcm4dc3cDUFkfECEEDya8NHjuksg7KpfcszbpaMAwMenytQU
SlfhBDD3b16Rt0CDpKYd/h+LmhWn0jxKk6T52ZNF43O6IBbW3iLtSbwCTpVDxXoI
/bryb9cp2qpencITdq7x0LVj1hjo5SiJfII2CuwwK2xf5E7mO+bEu6UuTpB82uEN
XtxWq4pgVZLX3B6nN98HF1gd3jevlnVvx/G874IlqY4CnLfPz/Ha5u73hf4BV+P/
XIdpndzTriRaXWMVMsj6qQ5ODycKmwhgUvAic4+rPAmaUscX/jBC3kRboNxOcUP0
GYkjKIKNE3fdmkWiRHzAN2nIo5b6Yq6g0YfDVMia3JsZdn0svKF3gorMRFpnnmgR
GMPsM4XdsY74+Wm70HWvr4BOjbzoB0obAcCV32thj7+zU98Zes3gC1gHhVprDhhw
InzlNKBytdR3CgM74GFSv4REQBYlsrp6JRJ+pa1mzufFHyCAfU8cfi8mPGLnAA/V
qu3v7WEepzaggT/L3cN31lEjQX1/VLD+hLR31Ykf1BwbiFQ029ZVK1ZcVyt+txDP
hDeFTrXAifzMYk3ajyhe3uRZI+aoTAFqqfaSG99rWzqq2sKfqR25ompUBQwDoU3o
doTgwFsvb++SN8nMbqwvgFRU0Ew9c+k16/xmpGvXZG/aUQ3ss3/hMK6VePsnRg1L
tvwKod2ErbA3rMsEnEDEKH8jULmGtlSlNwlu32Y2+hR3izwf+HqUHlOZrAZjzpz3
RfrfCJMIQ+pS6Zw1y8zdR2yHahJlZJpd5pTjJVTHA5VxaBo5p+SFYmbIBiBF9rWW
QH20Y9iHaidJqJtYg5vhUb1JnWJxnQzr0pznL5th1aGAtDVGZ+WSe4VePKBiZ96j
G+xlNI1D9UJ2uJ+cGh4qhQgybJtAqep5qQ+XHJjFIaOQZYsyK8X1SLH3wcLexv8g
bgk9M2HJWldUzS7jbxc0STAnaJILamaYgWOtGzAa0RPkbUOo/QFLFIc1DMTtUM1b
CXeGSF78XANN5bEBk5KtZfT5QbVfdBKU7rMpIlQ3MXcY24TJ2JxJYTXektEFE6ub
AUcgnnKQTCPDNKyGWdb2VFRJfggj3COiVya/YTJgsrH4my3p2hqsosmW4KaGnQtp
q74hgKui0Rl76l2VqyPzdRnTeLklMhPWrxvQojdhZ0tzj4aF2ZUWW0LTr/ZtP/sw
EpHe22VcfEk65Gln7RBpS+DaJ8bwFLAKWqj7EtCH3fet8hSEe5IbCV5OueDi9KHs
PPTApRgcE3cy8lvNnGFr+n/Fe+Z0Byq2FQNQSnEAUcj9YD574uxu+gesvaIwT34Q
shWUnK2qjjKpp4hqAS/sLBdnBESz8B6xgbFzXR/oQ8b1+XxJvN7KGUOrJd4XHiZf
ADqMknvYWPZ3//yuj6GySZKIJcdTaBu+RPqvLHM0ufNe5UokbeqLHFKXiBSyDGMS
jjoYvUoSK8tI45wICgpr7pibCZ7tF9qYD8gj69mtmYuJdzuWjAA+3/VTYkbW/YxL
CzBOxheqjCAfWnG//zxNqfRQ18uVQw1nkk56oIguuaj+JVCI7ybBnTntzPnKV+3n
l+JUySmUNAogc2AGQraxRVM9g55jPhwhodzmdZgRlZzlWSmorXDWYzGcw7npkIwx
Yl0E9waBt7eodS3h8A3jxXqTjLRNZyC/PQA5DLdhVOA7z/s9HR/0tF5mOKuqlHTL
8eQViuAVPTulzFHc7ac55wDo4AVnMCyKFdttG6Io2Hm6w9i9KTKWWwzmAKCAEs5U
85DIuywsOXdRP9TU/Pzoi/V1x9dJP0IUkFEGvuIZXuQd51PJTr6WbAO+4MG3cb9B
IbdGS5+KYz0OoF/0P8AB0di4ueTTE2NhXqT1KADhmEJAMOgijtgFYjpGkrR8oop4
qqYCJOCq1/zc7SsY/QFtFAC9PCneREPtdhWX5Kvmp45rB/QjgyjOPsY40G9VN/gH
2tI91I0oUf+BhOVRL1ULSwkgif3kaM3J8aM0B3XVjV8RB03G5JFMZ/HMEz51ojeW
JHTvVwtcLiL4DCrduue04/xXTlOyELwd1izGbitzLq5c0+A45epkTaSB+ViR7Kmy
U50eNXGLgdXJJegMGF1/+LEJAOn+gUnNSp+I3ldnzB1gD0Cul3mfJHxj/kxIBWAh
K4JXqnduOqTACC5K9p5Ps537xruG0MVlsypb5a9AnJNml/5jtMwa8sGcJJ+9kxOZ
eUXzFVw/GpSLW76Rvg900dmrspbd73ieJiH5NJZuCmeNXbFMUu3CaLdMSzAxBUy5
FRb0l4jbAwRlrlEBcZwIbyDV87CnbUjfdxZ0bH1sQ9x52T0ICHT/AzaEvoAGYho0
SVlMFCwADx26haFuU2ijEljwDuy4uXuxopXt6nGbDAvD9H3KYAuxPimFe2Z6nTZz
NOIks6DpukwV+UUrNbz3hu5RWglzdWGU8WZP1GzPASGjadEkocwoOgJtrBtZVCvt
P2XXe/wmriLhqXgYFdwFWLOUPT6HoM/PSZEh2qrewS2PUogdMPCZmZa8lyfC3oWn
0Y/93PcuzhLTa9oTQDehCRrBq43OEhy2kdtG7Dt88d6eo1Odmwy6GZojRLbyildE
iyKnH9P0inl63HBYh63tVwCu0lpx4iCoMRHuW0S3eg5FUMPXLAiMS8ugENSuRHSy
7zzOVIHkZEHZm4VNe+kHAH+q1gIELrDF4AYgfBHNQgFk3p41HVUu9srYKJGi6Eh+
hMY7Dw7e50zMxyAw30DXmUrC3DSL9aGfwoCrbKwF7LQCK2azfNkESbLM3gT8eMUP
s7fX3voWSytsyYfJF6plp6DB5NtAoun6hnTwBIZ5bxiHBjZsPekWiHhtBordFAYw
b36SWZh0mW6xVORpk0zwk7gcv3gYp+LbrpHCx+vRH/fDkIdmhCxpPbowfRjE1tTj
ogGBiyiSikH6g9vMZq0SCObXfuu/vWUOcBUcsCNErLf9+6xmAM4Rx38aduigSgeu
vLgqs/7UqHrRFj+/HNVOuef2u2HwRA3o53W05fHXwgIQ9BJVFxq+85kHhdIJhGm1
imG8IUf6XIOTzqkPDm4t3s7AIWtu8bjaAmgpCg1kzinbjpX1goitjBBtoaWpGWsL
JbN1QRBjQWFaPRIkCRXiEzF1vjKnULwh6V0nQN3rQ0F13NUuaTJTMSXVFu3oBUdT
jNAbj532R3wAYLhw1ApzeMCGWEqxTog2mNgdw9csIH+rnUqlxnRZoT75GOaIFNpP
WwWqEmFp5gBIVQ9kgViyWlVEtVRoO/NrHNxpkbscluel1+AOxW3+AaTjw617FKDG
C9R7wymxB/Ie3xgNRLrgwjHcteTKyxxCXAqftm2RczvOxovrimb2CvxjoOAoXAYL
rQTIevrU6Ws79xe0gcaDo6UhxFZDKHJQcy8SNsCEDnfLq68ot5WDfwgzZ5RwWde+
aKbOlHM7IVrkOQrnfTJEQ936jhjkIsRnFkUbxt7OHzRAIM7KJ6tZ02FfVPm/Mljg
353uyw8gZmvMjNb6V8NrfvSz1zxc18NiMrTNOs15CZNvRBgWaQrJI8aIfTSpp8xW
KyX7nE2VVF7Hig8Ag7ySdNu7Rz+scVyMSPWIWWfC18B7EbSVqRtNJY9yi3UPWAsN
OA9MRSnb/24o/iA4qI1uRmD018AS0ngJysXNIweuT6TZ4MOdz/oA1HSEGaBAgtwB
q+TUueSieMs45HgdUowlh0arp8X0OHYrn3VUL43QYYfWEmkfORtayT8IEYUts3Jr
G8ZimiiLxjJF0/vWu4YOYMkmgDt0LXkAky/aEtWHoaVL7sBxFH/rSsWonET+WSN+
Jc43NIc/5yUzH0z3oQi/LpVRI4W7orJvBuhPwial53uo8sMLJIqeZhIEcqSPUriF
QLSTMcRmx8tjRZGBoBHJYH0EU9jiIT1Q8OZ4mwMSNpfvsDa16SURfgvbAFVOLq7q
ORNNLiXe+itCjYD3rDyg3Hu5MJRzAElLwJ6H5usu7D8iA0lYNvg6P9Ms4ZV/X0N5
4aQaYVDeVNmtPQUDZV+eiWCEY4gMvgM/41pmLDjYmSRfPtefuh3xDnATRXaPEIi6
O/pLYZK7lE40w9H6Jh81UbcWJCvtXQuQ1TiVmizKkfivIfKatpO1Rbaa+IaRP5KL
EiqSYttJPMBv6D50NXmtdLU2Yu+b6vKHo0qAs34kCffv5/w7hhEBdN90x48l82YE
t1FuijPpNOEMUFehfGVjyBkDrqwwsbDJBqEyEgiDEx7QiJ/uP6hrwyooWpsA4sdR
f7ha7M471Z5XbhhyF30YGwnzvm1v2PSYDosKTSFBwq0uuJx3ng1Qn8MAJIjSzzh7
BeGVMhS0mJ9xjpZlalMzBUQLGXOlnYinFBhr3aFJqG41iqluaXRmel30Nw3CxRxm
RKjQTwRffybzSfV8F35Rbn6UkzvC/tx4Ev4ZS7mk0KrBp+5Hv/GbJO33OsBPXb30
nO77IJa6ZwWbYYsh6Q0NoqY/PvJZHl25A26BRA0k55dsXrSDgWh1aQ9Ipyb0RkFK
o7qK7qoZw27TtsPdLZMofLBZli+ZXJcPHG/ZiQuG2CoWKJaBZYib1FdMVGP/ge//
2BdT60M8skMjn6FYhWtlEwS88STrdgyPvn7jkQC2GRKf35OdalrSXX35h4a5Nd+F
x5Rg+rA9qbj716XQqua3zwKufiQp0vPKFp0czKLE1a1OklKXQjUCvO0K0oJjsm9d
rXahTDY0LsCtnjaP5ygDqG/fN4W6SM95sEYdSds9E1KWFHLcahrKlNvH5AcTn4eQ
BOyoGzc5lGLG6W+wuCaErjPI+MNavu/2FCnBVoLTF4DhKbwJTIxwR3bM3UaJ4ytv
/nzV8Ku0gtpIZ3sYnbERwLiWAotzbXBM3hvZLgQaIzbooG8AXHBuSN5HICHrobHl
FbhAfCim0MGFhGLKZj9e9sJ52MS0jk8rsFQ6N16t4IpjZdMyxDfJrmJDnlkRTv1+
nNkPo2V7sYWvMIlipOt8UAhLSHG7eZTq8USzuUvVTUN+mmPcvFmxPYhlTyS9YtW/
6ioUnYN+cRhjG4BYyDwa3sy2tsqG/8rOO2imVqM/q3IES90KFL2cH2q1ZSrhVu4j
9dPY/qlYpK3MPhyP/KNTs3tC6uwmxnD/aWeBVhxGtSFbmIXTxJERZQ7BRcHt6RkN
5xxQqec+t5P6GKElj2C6PtNpDMStCv3GSUFlEIrOjeyL+RFeWvygyoo8oYmn7lja
ypyW9WE8WWQm61Ozf6vdPPSzyjyo2FUHUNE8C+aHhe/qod3AiQeQNDjIwLz2IzSY
OEgKzHi4jciTBsBfXPmythc23cmQ2tCkp6IGK64u55Kv71eoXD2Qs92ylhbE4PJg
aw21R6hvqU7RTzfkxdKIn495pOGMMNtrhkAKjMHtBSdqk8GFeNq1ej1iPkAPjy+c
4QI+wdUI/FRHQvjtCPaoUJyRbzcKtdTFPOQ1gByYPJAzfvFCPG4LW25lx/K7H/dp
ILAJD/czgRxvP0i787H9dPaNRqmF3K6Y6eYsv/BpszDOugBpkoR3v1xwxbopp5MA
bojNahhORAO3XAiaMkEaR78YWwGcuT2FfJq1rkztcb/uXld4sSzoSbA9phW+0JGF
pvXlC1w6XZ6Hp8CH1QdwykVc7tf5H9P/0ZG63J3+NQlbdYIZ8fLxiP59s4yQ1OKP
mGBTyxWqsTPrXME7QcU2HbFxLFwAu0BjQw2JYKBEO20Wkx36zkUkCbSfkpKdZOzy
YAi3zS2y1Yht0BxRz5M8N9a1t/b/w5rOPkrEMmpnsXkvWz65pXzLEft8T5zmToy5
cVoFt2zgyAtRAx8cvwRWTOIthdOqRGfY55gH8gjnaiGJjfhY6AvITgMw4Z7qEUiI
SugqPwaPd1LE7SG0WcfiJG0zYDrv7/iP2oAO/dbZExNVTzSTgGZvvkNDf+plpXgR
9wg0uDfgHrR9swuxc2ziosXgLPn/TtHw1IcUIx6nsd6PpO+oipL1389dPIiIVkYW
okfUSKqvDFLL8SchQznQoLIpw8cEluYLkWpB4P4MEUStYn5+34c6+y40mxlQ38M3
6P6Fwy3mgBEelhZ6DRwx3itJ8GRSaRLNtbUWBO8/dqrabc6sSLXrONOIq3iOzAQP
vEqFCQJXXprn/soUaSu2vVnTA4Uw0hmxJhyNOwZxRe+AWePkMJucdkARRVwsA4US
wdcBJq2J1APz1FvHspD2iz6sOjcYRBq5+JzovfUCYHs+Ou6i4bADz6XYUmYRKfrB
lNdzzkBbxXbWpYvvJCWOuJLA/CTvUZyEF7oYfJwyKl/3BTOnTtrPXBtb/l2Udgx0
haIUE3zPtTG2NsIxugULlPJMjStFkFeuPMN5w5FxiRZ2qqkSudM2yu9y74ieZcx7
phHJFbPZZ55JblyDifXJBLQuFKdVpV3nG1Gz29UbAtRZgn69MxNuk9+nOUrHlB+E
E0LahO4zJibmEUK+hmLsLmqWD2tfaQ3mlRdzr/YMKHUxVqkgz63ZLP0Sflid1oOs
IQy7oAGqy5zgk2wByE46ww==
//pragma protect end_data_block
//pragma protect digest_block
Y8mYOFzsHhI7Uyi4GNiazNkhle0=
//pragma protect end_digest_block
//pragma protect end_protected
  
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
NsHQOp4Bzvdvl5Rxt06zE4RgvK74GKsOEqBqlfm0StM+AOtT/ibjVSvZmjHd61Yt
MYBTm32ICl9SpVByMrKfOvA23ty6TWA6hJoGJ78dvrUWeZmiIQLYLhgo706v9b/L
9w9QGY2/lhe0O7ANJiG05+LZ3rbLlBbcXuz+E2RBovN7xDM1Ytf8iA==
//pragma protect end_key_block
//pragma protect digest_block
ayCypvDR4KWtSe6wNirS79G8qRI=
//pragma protect end_digest_block
//pragma protect data_block
3T35EuCUoQOqdVsNdGf0B6AAIPMYVyl/tkgdRfbc/DEXUxYm0AsSGxc9V1NLAiUs
3VBOnuPcC1nQzdlkT9L5hFMf4r9gZgD9Qeq7FVVWBnmh5AuJPIQuLYMEcdQqG3iM
lw7EGXd6beS91ZV5YZnmn8m8b98bT8dY8pxbdcKdla2O+1lY2KXe2eVqkYmjeBKz
hSa5m4LMfOn4UOS2oJf2s9RjLd+HMlmQPmWriCRrK9vlyo21r3T8HNG+5BK1evml
q72kH7IaUgXD+9fayBqN93MgC4GUE/WxmbckFwVSqCZxQUQj6J/aJD7vo9MVW8Qx
jJyxB1Fhv9f5TaIPOCN/FhDJ0W6fcodjKkP2fSqAK0fqsnS8OY1x1wR3OrkExt3i
xZNmQ3DVquG/nkX43zmewq+figwqIYKZT7+ORDkCHeHVjfZj86ZRcyOqwPbrrlNv
MHe/c+dIxAbJVeYciBUtc1ulJWcrs4mKJVsxLghUozdb03kcDcEvOGhXAlPoea0A
zhFP++BpTPuHY/c6P9SnsBDzRnI4z4Rc6c+kZHLv9jGEfrI8VIFYu0Nv/3k7G7Eu
yoUKIansgizAiofsDPNAoEfb4PNyxcX1wFa2HFieZuO3HIcrrTr8iPoJMUorlOGJ
kBaoS5XNk8ZT9xjvHElvIxUZZHn7QR63JDuEZRIFFPGBbhbQW4V9Ww1WlrIti9qw
SS0n1CFFbGjUNAxSyPe9jnZ1exXZXDxGgNuErERUNl3JsBXtfhnNP6Hmtjl96NM7
8ztG++OM83m6c4pAgmgglf1JTXC6qdFXl8X8S4g/hjMAeEkw9lFcInzLR+wW2PZk
NPHPhZ141UTArCmKEb1ukN6z22kbvIsWA3SnoCm+EIYFDqz8S2Hiw86iSFSaCVa0
ehc4Bow9iUXTHAQyzVGzSfF1QzoLgdyG/ceFSbtTDDblUIYoSP88gtlmtk+uHLtV
HcAj+CtyS3R3tVX4YIau3IKoWUAZ6s7/tonuGoQTdiARto4rrN70RfLC2zXOniGc
Tw6UmqhQA22ghIzHKdM8O0mVRTm5YFQRHB04UZvg+/TZYyCKoCYk86KHbduxugYQ
TBEwINIbv+Bgpp0NQ4n0qa5jumpJWpDIqcb0OYSTmIEJ+f5JL3+oncehHpDlr/56
mQgiQFl/HyI3jlDYJVbUPWWU/rzTwusDYuAzzl9w4QEn73hkmFLlLow2++MnTVFE
6rt8xY6rwVu9llDxLPm1eFhoCpKlbJXJW93g6xBtJ3wRE4ZJUU6sJ0qS23AaEZ+I
7pUWSa27H1w5w2JeDq+P3L43JJLLmdbGc+pTR1G/oo2qSQGtiPfWNjQdhr5aAl9z
uzRwTAFo7MpduNCg8aFCeH1VetX7PNbpFV+jf7Zoe9e5OTg2EjzEE2VCa1eSx39E
oeaPRIMpTy4Q4pZFS5/FShgbs2EFnCrjLqgonrXArbbEsL/+iY+FyqDVWJ9cOJj7
QxcPfDjIVxV7Xjt+cfI7rMRTXWpBWvXX+AHIUOMxkJHvVsFSrGpIVTptgALh4WBT
7x5Ft41HUNscCgkFYFcWisdGuXbuAi77CEYqPbm6AgI/O5Jphf4x3JKB8sZabhrJ
rc4sJS9i9WHSuA1Htvo6mbCxEw+LiJISxabcpbA8D6zK3yYSQmEj5WOcRtl/1ezP
jXlO7jh5/73l1F5Wvd2zRfAyHie1AZbULn5lpGN43mur+gJ5q71JXcIzXS6jyHBN
bDDO995oExZ4uxhhWXNmL9K8iKNDJAPuAEjYKwc4npt3z7+tavAWmY890WQSR6JB
kHbe8IVzDNLSuSWSOY+knIn/7iNPOABONW5LLab6Hpg=
//pragma protect end_data_block
//pragma protect digest_block
we8KlzslVLmApdQGVnUYR1IiyKk=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
nj92bBnqvrF/CfL9dIehPj0bR0bCSFC7sLV0mNj8q5uQsvBmaN5Du9no/wLyWmsu
mnbHG4TYBaR6DxzsmtthKPJMG1u8k21sAmOlhmqaqQt4AYu2y4cBWNP+J1vcUVVr
HEnUg4HyPAMYzLFrP4LGktrO74sTxhuh7HuQHFeZRq5QwZ7N/OvRow==
//pragma protect end_key_block
//pragma protect digest_block
HdJmrngQ5uFG+hFQb2gQ5oKzYmE=
//pragma protect end_digest_block
//pragma protect data_block
/OmMpADnIvSki0jYV9F/hmJVRJWYwA/Uq5FiDmq9P8iXDOfZyM97mX6jAIALwpA9
EPDikPsyQ8JlodScDH8lwLmjdkmpUTMIFzsq9OQvBBmwZKrmKZyhjZ45YAIBE3uX
K1Tua37D0cOMf1gOfD5sgc0IPst+u/Z8MFjYlDykiaqbqkTt15RA6EEl++gf9ceZ
/uaTN9iGWaIG3p6pfYJe7aPngxYbdgo9tIJCbR3rMjWdm2/JwEQD/o7AcCqS/k4/
f67RQi9/6w2+HVBoDDK9d9d4EjpggCx86aRI5RjMcKGoXMw22NEqComjros4Jj4/
CrLuNQWvMuXh8eOaEnn3BP4AXHZw1GR6F8was4XQ+Q8STvqObR3iEKjoJ+udSMOw
WpK6RnLvSuNhKdsHKCLzIwXu4lUi/valSnxqRemy0UHWJ0itg6WYEhkfJy3jgyJe
4Y0ncGJzeryODzrtyerc+YDCCz0vJMpbt4rQX5vL0Fwp9QYqjtbG29jlp4lTeGZe
IdMnn0rHGgsyoXBlkRvWQShW8geY7AQp/ldMysWTXsuvLUeGrZuUItDzC1wPXg3Y
bCqZnmrUsQtzeGZGsFIh23xHIYu7oyx/hGEQ+fabPwUl3D0xLqEe97uMjfW+fy7I
L9OY0ZOMnwLdb46s0Ou9Zvf/Y9FeZ9mNWaHzDNrQiuqGkbD7UjtX4CNR8KlcxmmG
HTMUjCvkymNqH7hsvZp6Fi8cXLodemu8B64oEU5z3kdzrCy+BG1iIYCrKhisQ3Cu
Qm2CRzrp07liQvHGErZro1Q5hjXViordY2rlDf2xLqjJ5rhEd3+ycUFCTbFrvUsM
RJybblxYTbpXKQQZBXbkrpMatgEC9h8CDzJUA1x11HrqCv/fjN5pCYcMU13C0O9p
dEu3PidLfZGBhke64YQ37XydSdAr04vS+KNBMayr5jcbAUzTPF6cI1gLJETQCDCL
r5JUagoUwRU3eDrg0DuzUoJF/zozvb4Ay5pX+XDfB7Oz4gcr/CDGN4MHUWlWIL+t
cSJekbkwOAQYyxcbc/JvgVjC3RlUtnVI1mJhyPVvkUUgjmBeXUpjtXCHEmdQKOEl
sCtB1AXKnmjAjzIQDxU4hcwoUgJXA/oryl3sklfYxH5gZWtpQEULfm0DU6uKFHKD
97fehPJolvp5kVab93KpoF0rgPxo57bWzNFuWFCJotWRItX5qg5NWwfGfyIXKBQC
yV2N1rfh9Lrueu/GFrYtMccYSB414kGUilaXBpHOOo/J/J2IO68gJzKB2qEoQV6d
IatGBezdmdcUh4PMU+hCm2fzoEmS+ZFqT5k3/e5Vv1yYCl/4cXn4A+NIq2EKEFg+
Ibukd7SzIDJE9LS5CAyuxJST4e0vcguhUY8epXQMfOfQazHubReVxRErtgkhCahE
XGJLv/5F1FPVoyq9Z/eHMH2f4SyTW9kUGYgi+L8JM89vWcv9fz9aJqDZQ/TDZolv
sp9mFXmW8kUkr6TuurtUbCAYDT2vBjN3SdPRR7u9rg3vS67WIhqikItOY74s6PMW
QmNr5f4CMCJti5OG1Y7fxH7yTK9Qjsvc2p9noCx9bLzO07/63tO0KNAf1T7aIhao
ppS11nvwK0SNbOALwiJNMmqFtKFXAzzJPDiuPTX3xYyYhQbypBRPAdqZ4YFY+zuS
l2z+QOVAr3ChT7Fpzkeq/Org2YR+nZ/3Dd6JiRuxTF909WXfsyfT8Dnwr6lqgAM+
z6/zsIQiQ9O8TzvOwidNmmgQ3gqjaZdwpyZzIba20oYA3Oq5A1xOCt/+zJPYoavy
C7CBsGu7ef4iZOeOkUN2gUongD03KLA2VxrZccxah2K3Y3NUgztyxo4vGL+sUxvq
8DrmNiEtk1qenOAyjLiqQkKuWPmoItF6D49Q0dAqXx+Ss63l7+nSJaQskk3SYnxR
iKVa9g/hNtDXxwwmIhHBrOWTWbWfTx/UXPOSeYnsvGTAzXo3W2IEZdYBmD+x9xCI
UWW+KswTy1q03xsr5/rRgXN+kLw0NsnktUN7B9spctc7aruBu4bQGc3bviMAgF2Z
TlkdmKJxOPH/qP+L0NU/SnVXTeJXdHiaG99/jzKC34Egl3YSE0TSzCwuGR6todwG
AV6lXmdPklN9decn9ZT7moax26ap4AwC3lpJBzzizLtliQH/4o9wRW/LRf9ou4pA
Q6hZDHfP92TnDMx5gmkTZ4X5Qmjf/VvG+62Jz4BcSR1XQTn5cSgoY0aN8aRdXzll
knJzbQFSTJ/im93eIQx8TC6ipyTz/Idksayy3P0nlYXBaW/VK6thtdd/UcQE2UCa
tju7j/hL28qc+ZfLU7pVYlmCfergTBPTnCItsloHBBZ45QmeIrCMzPCMEePcouo/
twcDos6d6aphLa72ToGDwF6TScrHDffkZDhp+sPIKl1XyPAPCvDFk3MkS2iDi+V7
GZDiVkWNIOmTdO4KFU2HahA5lKDrDfrhqbC+va8BdkD70FkKDNRGEeT2KiZiSVAd
wiKRGuupKKrpQ7jeKwZ2T06m5nB92Whu3V007bC61qG+wu6D083Fdb8vVxWI9A9t
Tmd7P7RuYsLkj8K9ldQ4eeVGCn9zGX/rwY1uUl969Rw41FWB7cGv4Y/nl+ZPI9zX
H4wv2ZVsC4JilaK3Te6hiHksgXTgn+GMEQC5GpMqlNUkJ+pM0BwJO4xkVZA0FXHs
6uqzN+jzemUxeliuAARTiHdbWpWuMVa0u9eT8pmkkV54c+R2e+mkqNwLKTkCZFGz
oDpXJ7HoVxBeJjbMx/JCGWVrPVFPLthbiaGSEf45arK3nQvGs8bWSbs/eXPF+ZY6
6XRBDrhRVu8nduLu9aWOSRcKYFJZsHvaVzscPkBo+U/QeFuNGoERBdJT2tXCsP1J
qzS2VaCXS+hakx0O357SvGHrjpbz3fzv4InBCyEWiJwtFK7EnHuV6eXj+c/l3RZb
BT8O0HrdYWFy0xasCEljsYMf7zPIcgBaTAowx9MpydWCODQ1FpghFKRwVY8DcKTI
6J9uW3U2ZH8QiIMTaMtGlH17fu+4vxicwHzBMow9xfPtV2OTiLrItabO3+MgojLV
TgN0QZlJhUCIV5ME1jbF9JZhJyh/6jSF94GzAihXxFt3whh1jATi+aPi2BIYdlPj
XxMy9EcWjfEJYMNToWvtWB7ZBbeaZ6odyl6ghoEC0Td/Fv2vugz9jGSnNOk2oJDg
H80sbigOW0cGhmihBjAbRt/KEnw52bkrKFd0dE4FO2ehFORVGJEHgInjf8Qice01
bJ8HkngxISOZzWGwEL3jolFls0Uue5i+xGTpgKYjlr3myXMKPZFOkhPELke+l3oM
iwoAigrSqU7bIOHk53DMWYkjfvletStJ35jMY/YXIfAWKpKFHwrGhtPlsBFCuGD4
49Nm7f3AObWYQ2IZ/0jS0LiuY3DQARUA0G/QfeGbq8WqPGd9aRRs0U9nRfbLQUWD
MdWzHI1F19AUW4SmPKhbVa9gghuZFQ1G3bRxT8+M3sl/JkNiuIkuisP5SRFEF7/V
jZk/nW7XGA5MfuYNVj6xOXoNvl/cBHYhMAkQgoYXyUYK65rKDFVwqJXXOXZZeZkm
gtYrU9fet/hF8i7DJX9bEpv9mN2jhhklVzyTXXpbr18RB3go7whona5Rzg6EsLSQ
0TndaqRuICN/Nfi16UhdBI2gowspt0U3hyeCovQQPfBfENfDcYihFpEGJoT7ubw+
QV5scUfbZWemdIzdTOl3/JwLKlu4DN4wmObeEavIEcccG7xgcnutFpqZ0SDkRBIE
c5mqb6ZFjTVkcMgH0viL0MDnJld7yeuL0vlbQEPg30nEdlENGujGChbCuCeBuQHt
7bqCFC1Bg4DZT1NLSDb4Ci/x5uDuXH0AfEQXfa3eXkO4iYikikoA6EA6Tp08NBTI
u/5+yEpbI1Duo5vpWJ3Oq/dYy7hboTjBk8FrzhxVv/NCHYXo8Ologue7A78yz1Ok
8C/UJZHRGEA+wRtIMFCEsqVdpnxBIp4sKKF515XPoAGZjKqBNkCfFcFmEoCnrt6v
EWodly3G7qKkEpM3/FCcDPPeoGd4QI5ilzT2P+k0feUvr45ztdU5X825vTnIMtWS
73pHOjfq9uWfyuCZuG0cLyjFcDDMm0dZrVwBQcrH7K1x4rNM5E3qO7ssHpHDdNqD
b+Qi7jv8E6qOAbmeNDrt72PP4kYkOp1SsZBhhxUjZniA9TQkfs5gTUhQ64XmHaqS
JqFval5i6a1skRCmqr209/7WnTV7kIM5vaQLVYpXwhWG0OGzHaRLv0gU58JFfqCY
SZhRMGP5/87SvyIzrTigBHg65hJuQ9GGsOjAfhPev6WZJDg8TsahparU0j1M5zyV
/SPiJhg/qmAFK7r6dOMCb4jtgRT8b3sAn0mL4zX/6poftgG6JRTNKtZ38ybflU4A
KLOwG+wvl+JSIu6ox7NT7r7ni8gJu5V3m+LUu1sEI2Rl3h5oPg3NYEauAwYMhO8V
19kdqKe0TDFVHugLM3kXkZgw/A58qeuSI+TOtQFYCEZ06zfdpzwui6pgaQdJ+reE
ePXRmhxv+ceOpA6zr6Gr1/mfPkaAFIBCeUHW3icviOVn8ak2ephOWLFL3NIuHKRx
x7d0Y+6U54G0KARKDJkGhTBhwdZIwNLbjiVzOGSZr4EFbtgp1D6840Nos65oOFIL
gcH90QnDtXyYWNyedUWmCJTq5HDKJ/v702ZWpKNkLhRvvMfdHjnrVp0vwb8TgAhG
UXyN8PWHSOMdSSsHObemFy44pxMPM+M4zHjhJkAs0D784yGQs18t9THIfvzHhSXz
GV3G/94WHAteIWZ2s+HAraNRuzuE/dU13ox6zdEZ5JIe+JpBmLSXE5PAayC3h45S
QFfyJ7w7QUSqLKEtrupIOc6BypDgaoQuTR3ii1Z+hGRZjYN5+h5IVRxrIQTWfffx
FsHsy2AUgPW994c+iCgt/IBe0FuzRCh1QXTzGhu/CT4ya129XH96EWS1jqRdtBMF
f41H7hzjfE23GwN9ajAInfWGtOdxLWZPtXDhG4lTEo/oFT1TWDIqYKP2l6Bxbx1w
S2mNYNgPYtDhsjeGGhMLzhYp3wFQwOl42s66IS3KbWWxNLOtf2LeBkT+chDIAspH
sOTfnptF1kNUMIpPeui/YtQPcIYpu7+X6WSZNIny+f3KE3iCHTj4nTizOep1pA7e
pM23CXS94CTlUYQJ204eque1C3SBv/3eq5HHWBFWMR4lfvXmANmKbDeddb+S4Ar2
wRxxuU7OOl1XLjag9IiJvzUoM1LPSIjUNpj3Wq2kLaah/fXC6LIpfNTS7oHncj0s
uDhv/keUW4YsDQPyUPDB3qaIUPlipADfbnh154LCELqI4rWa7qKs3M7yDD2Q+OWs
hR9dF3T0ALoPhhrbbvrZBnIXjhUXYfJp3K/heeDMaFiDO0qKAbEkxEsaTo7t+Ymd
EKeLZKxti/qRqRP+BuvL+YxstwEEAjUgDKE0BJ5xrBr5CWYPsASOB96oxAiu9faq
77FptCpEZ4YU8Z1XGucE49e1Tovf8NKMH48/o0OkYpAC0NA41GsDhA+6iEBfuKvl
MAd/i+uS+0uwFb16ooEXH0NSZz9X4g3HGEur8bYmhAWa/o59Pg+ou3w4eYqbNieo
cJnlhwxVlueS1X9XqUx+2xyvYDrKmpRlzYtTb8BwcW2V0BXqVyyRt+ue12/jYjrl
T/d7Q7l809vSG32LXcj2EPJS0J8tWn7B6MXSZbjdwRkuifVJ+IZl00v/L17AQHoF
H6RSGhUT6+qAhPc4f27/RMPMwVdLtXiQ0/RanWYdWgRHcZYgsUCmsDeWAXlEEC/n
nwf2hy5iTYKXII0rRhy5JbPH6uEnnmoBVp5/lYIkqGAd6QhwQI04+l1hYFo09kWC
6fzA2hadJ3vSqPmODGCX8GKRgcvR+5EV/mk6EpkSzn59H9eFVTzwVuX8Kt/caUb9
kwFRsU+dAWjdh6//Nl/1JemaBlrSFhTJ4hlJFqeLkfD6R+aBu+NTBKcjcqUqFaZj
VJnxW0bjKuTKdWK1p6w8Uwr+Dk5xI+4Cx87Ebbk/hvAT7qijILAOpOXoN/B49z0K
40nGNWe5ZMvgfIwqFjfX3+zb82lFWqYxxyo4e31ebZK1+wuimMB6tHW4ZMn4Ah45
2zgt/sU6omQ6B/XZJRtHWAlgSfK0bujrUu45tve/JfEP/XuPvk5BfoWL/xbvvoiq
n91vxChk/4QLMKxIzj2MarvVHlHnveL8NmvSPzL1C+UykNdeWcIwUfZYIWX4XdHA
NyigB2SHYArYzA88A+cTY9xev8DS6MqE7yMtnt/ViTVEkWHreaHR//0xuw3J2tWk
C8RCebYS+40KOVhkI3qcCOrvoU4PNbviAhh1igtmBiNLCr7wV60kH3fKzPaXkgOY
IeazE+h8ZYO8TlJ/orKHfG12Ak37NYWsn8e9Te0YacmFSkdUDW+OaF/4F+wROfeM
mY0b463HdEYj9u9Ta+RAD5iI8iS6Ts3iv10ck3LD+vdSaqCtByGrjqMvkYaRCM6I
mC/PUAdOpdPmcv8EFyh+HgxhOOUYeu583CHRDrSuADHMXw6n9GICJOWd0aPvInAw
ccicquE30frJRVLH3FWJKAl/Ir5rqtOrrOEGVoHCWzJKqXdF54PBUVSL4jlDuU5y
aFqLQEcbMz0LF6PIbmQPvTzXSNsxz6b+3WLZrcY7r67sp+W2NXfDRGoTWOPAMe6g
u6JSFtvhJqtv4wKrOIvVEDtV7AMg+ZKA1FxLby6XPYxYZuC1/qbzoqvgUq9xoyMe
jpR5A+bK6kRugbbSS2wExhWV4YMmhRZBKfAcXJSiwSY6G5sLOU8ug5aduH2fXUwA
st+e+QgJaYpDxDNM6F5LbB0hUinqc92CADWWG6914F6enw3uptzrQw4bciP88qEh
w6jx7jq3l8YizB1wZtbgMtuOsObS75FA7MSFpKJHdTpj5gBoauwQYBkg++Dc6h37
zCp/Ch3mOuAAPhDHIS7NvHPTsaXvr3K9ieObH4bfkDYKQUUxsn8i2Uam+B46FEtS
zST29idr3XBPYix4L5Ue0coJADlMpf7rUChTghxWADz8wJu3xRoYWKzkSJ0xyD9y
5e5owpHpNSHqFb1qwaCQJvSqeYc1jLHoLY+l/WCBjGEXAIlqfrpW/E2JVF7gYBIR
vBn5lK20UFXxRyYljxwYJFn6VBwc8kPOWU2V3/J8gv2si3FxPm4EZPoUfZjLJ5xm
sWmo8Ans1GzTiH3Z6HLPXkD97e8NiN0upWvudDbQ7d02QoHRrOlIY1s11tmm3heb
kWwTWBsQS8G9dNffPbsCbGdpbnGEgyJNI2FG3RXsl4OWx7yP1s94wvz184ECXhGd
1icy3RESKUZ+04zLmpIeLM8K1UHCFSslHpxMQs5XdGDgw7jC4jMfCOQxwmYiZZwE
ur2iVz6RWBA+UbOwAqBRZA9jGE/QjEHPIdhZSG8ju0RaXYWQvkOaIiLA54G9X+px
his/jjfxvKyHBySjRWAkrXT4p5TMbrShEMUmLqLeluP6SXtyG+tYbmUOxNEctAiQ
gUB1iwPuLaNhkKs9jk3ojkmD4kiBooKGM3pNQ8Yy9iDkEALILhzxELWdY75Q1JIw
MAhaFCCsYWhRj9ee84n89iOEktu0H0Tg6Bpze5SH2eg1zAbIXTezJSa3OAslAEvE
eB18UTjbiN2He8R0KJ9BxKU9hdhTL7hqyr4vmljHaNdcO140p373sCJrtJG7viUU
JE6jbw0TQnTjtpEGLtg6oRZ3XLhrw7qAvzhF+vDwsGHHRYmo738VVW60ew54OS6S
r9DPR1qZqpHbnMhjlYS+3JvVLoQrRJtTQMR/opg5Gt8V987XQz/nOSrbNqDKoTbL
LXdcX/4RT1fJOnfKjpD5LbLWo3NXWwLeKcHWvNBbNmkYGMXLrtErdIL3Etjh+LMa
/5Iajqt8/DRgFpTARqR2DeGDAkVvo/fnecmYIVIT8nZWrgO1TJULdQmOVO1C0x/Q
CpajS6uj9//fE1WS9CLEdSTz0RdsUnzzyaWD6SufkTHP+Cwc4X4zR8oFi1vUfvZ+
wJ8xuNftIHMRUW5nJiRzwv0GGP1aD9WsREbbXxbuarCffIdanBPWGB0r3iw+0mQX
aBU6VjOtlV0J4rzdnDNeXUQ5K2FZnJDJ4kZwDXSwnRJ4qL8sBvrd8ep8+2f3lUoI
pTHIHXiWTfLF0vJ6s3YXw4ZUWuiFSj3+b7YItSy3HwJpnGjFyKVCaL6v1606bvuz
LfF7vMSUljqh8ZpkVaXo6mXq9/L5RtAQTmUWgsFJ6lDBWUZDPLwpGeHgfODPvjpZ
+uFNNrk9XjZcIUGaTttULyY+oAhVyTX5DT+eiLxeq+PhdFQbRRPec8rEttveO2hd
pvvpeHqCeP99Y4h0e5iX0hMmRNbvY+7wzQnz9D2Fx8noQ1INLfaI3g3VWZyMhKE6
AsF7adzuAUHoHrouPt2tMtwEIL39QTVfrcu11W1Knzn6rGQVtv2iLpmrhORb9Whg
0Y13nFFAVh5BsTTJgvj2MbwasyyRg+5i2s/kMNHa6AgvzqaQVFZgzyFLqmmSEbwB
9d6X/tpP4b5FEc338YhGD1L8Mhaj8bOE6mf84A2WGrKMVJ0KYawnoHgdMraUoTOp
7Sqqy8twttwH4rk7GCFu/CLhOjbgyTIk2BQCQh1Eppost25NyEjumSCGIJbu2Ri4
lu0jVJIBp7bfxVEj7aXCFxU9spk3aeHJM58xTeU5DkOMtIbURJA4eDVIOOcDfEw5
YsXBMe7tu4AN+1th+esJMDwUWh+0awUn2yve/uXpjib5FXO0/t6zNxlAC9TSTSiI
v3zz11J87OpH9s5ws4YbADfRxd5oHqON3os9p6m5rVmtOrjJwfusGhDsflxEs5nR
S1xlfvwntNpoXqehNkeLvOCQ1G8p1PbK2umf6wZWALof2ci9Z+zwl5Hdkmf2NlQg
qkADUiEnfRkS+A65hYk5E3lQLcHFaVGZ6g0x0T+s33Q7que2vPRq07Apm1ld5Oi4
Qvz9NyzG2egkOJ3anb1thadymE/0AxVR/US73HB9/7wvLoe9taRapbKs+a1sjodp
i+/eFlKBX7ILaPF4OUF22WdRiEuVKPmZaQObYF9IsnTopxfAqVFPo9DihJuSEyYV
Gy+iMp+awHJ4fW73cuNM+a6nnEa537G6bQRRSd3Ra/kLUbjnnFk6xLlNQJI4vB/b
EOFAQFrWOaLp3JKY6PQxfvbH+RV9LG4f1qEe9/KMaXs3srRR9QoAAPIeIgUgCQ+p
8wm2sr/XvPnWkK33gPntMiqKTWO8piXiwNHPjmhFB+08hgwP2mT7AwBie7FlYNxd
z0yqV+HS+YD6Zp55KOKQ8dEvidAxyZfJaGFs504E2zQWjJlh683k++Vl9Y30ccmm
tUo90+y6y+oRTCqnyFMn6iowDcETY0PoVNpqqT/usXZERnbHnSv9LF5aLBkljjma
YJtlLdPAGc+MSTBIW1A5eIziXool9nWstrwX2xwF5P/dVmwAzgFSV4m2M2Hlc9A6
2bgnYsSaJbGEine8ttGmDDYsrkQA1uaHKkHMHHD8PPMlY7DyBzE2ayEeSqTD097Q
L7LhAbNxgDKuNDA14ygENJiDqWImLuWxfg8xbI46fG/ho6p9Gzk91GsrbshlFs4I
PwNagZTPHuL6XOzuVVhXQTARE9fLsk7LHrFCJhtUPIV5+UkPdjhlgidA3qqu2igk
d+B0Vu0CqXBz9Gn9QHGxTGT515ffI1KmerB2BpItCpEN+YTItF9njLvm+7jTlyMM
q0Df+q+0/GjcUMqmaMnxEYhXpGzoeTu0I2Y+92fbKMVvbkJX7GFW2uuxNtRsFzKi
EvxVxrhWHMHJfYJkab4W+qFuwcxzw2DthgIxjeftMgEIsOaya4Y37qvVNnSsl9vl
mdIZWJJeiqTu5xipc2OplH+aDqJnJWbZQkvdwKNKUQ/OSrrdl44tn4rvdaOEZrCa
bIGKWh3Nm70Ko85jSXBKSVGYXQ/tG9ZFhUENSwYPmOmwXzJ2GskJ/XS1Ws9IjHfK
tHTWoA1K8iejLy57Dg0Jkkff28SDJjpqz/JFfCn1ky9EDrwPUk9vkDb+U2wI+//Z
i9jr+tGyZIMMRO0wMsnV7WRfyMEO6MDKsU5F+1w006lHIGJRB86BvfdBq3K96g8J
ZokoG2m/SQO1djtmr1BHKs1K1saAQ0jcJk/DnOGSaYjtuw4TWU1dfzv7B6nOFwT4
+s0KznWJvCwpvAlRYgOou0mrpHlA+mvkm2uuHP4+I5AZdQN+A6GN3fGMQ+35PVUF
Pd7ihuN3PZcFCfHFciDlkXJuF6YDrrkdH+TAye0yg7s+gmAxF8Jb8msWr2U6fGK6
8INCy8AvfGuAcp7y/KT1vsXtM0JPSUiDAJawc9MkEU1ZXLuH4b222ldtx+HRtaj6
wr+D5lHuk6I24rEKmdHYcCIVzdBFW3NWF+5oCQ5sqFd9e8C2t8Ydn5KgS+m/fPbq
04WAaHSq1KAPoo6Ya39WpfGdh9kNP/CNC7xSDSTvdpzyIqhgcTEZXDSb6InFM3HB
UJnUaXtj3OlAWy5w9GAoZ401h5Hu8vHTO88ztOu66Vepemq9lzEDEORR5s4z0gax
mHARKXh1RgE+YLGNfhiwcVp9i455hnE+IQVD8sIB1nUzVP2blHzoyA74erdND9jg
kZBUGZM0kOlkPzGsVgXxRpSr6nz3pyx6PPHqnU+l+skyAVS1Kzwfp8z+Pn6NK/yt
UE8U73wn8k6KcEK0qmitPNkE5rqXYeVUjTS31jqm76/fHXwDwgeTnjptBmUT3wt1
o/SyqLTLjX6sklsAMmXKDcXvE4dz/6RAfZ2p7kPHIKvdc0BwSzOVGsce3pk1I6a7
cHEEKsUvwGI6XUA3o/Mct+wFKuPajG1GIB2Zt9AYM404ETfGqL0hcmDEEEqFZgzY
f67ZNXi0ssCQtoLGzX64K6bm9Vqj/yfbkPb12TlCafHjVjzjRuNiPWioOtnUFMvj
egoSoi2OGQAjcdKh7sVXElmwoyMi0IoauAyrYpZNomLbhwBuZJR2LSGSdQ/ShfUp
I2MEpUObRFqpkPmQbu5sIe5u1O2HT4vDMddwhT6r2b4TclHt49+q3eK8uD9YAvry
0MvUs6bZRfdj93HSeuIHYvzLAPAFn3/ariuQFcA8C1yKbOITzXE7t7d+qlVH5c6z
6B+dSTplqTQ7gk5o0z/Zj7+nHZGg4ptDCFZ6fKRscjRCIpp+CxW7iz9Dd09qVjdq
2tE7hv5CT0A9773wdi1kgE8UESTYuJeJKnz+66L+XWZLcCEgQ0H4WIm1cg/HtUji
LL7nHcGoRgOz5/EHDlhEHC2Tjuc54O9leYOpj/TQmYJPOfNHwu9XDNVBiF26lyhQ
oBp14Mcc822Ib/uUFOIwAF85UxFzwGSGT6x18bdmKZuDRRqx8Q/YxGs76WjWNdTV
mbwXmUXXoZClivFs6TP5i6QT8R2fi+6fVuEBsH+WlP6W/rXRdFuinZH+76FfInLY
P3xwMAry8i2mZijJPBTh8UGLCbxFtInxVKXIyqQVBX1jjRf1tYFR/MnmIwQb8J6/
z8jhxUqLvnOTgSz11a25DqSuTx4iYCZh6MP32szuyLHnL5ZE14D3lroo9oeB34OQ
yRwzfVhsCLlN4BHHz3SP/s3uSHZ24gR7MxiW/1SZxe2irLTMjTSakC1kH6B3lm7m
PiIND7WkXIgwGxxDafLGQRUkSyC4gQm4NLkCYCt5ny1RkeVjkUcyOC+qEV6XcmXi
B78o//xchQgIzQOMJcmEjAMuTqPUyrl+qju/xiVVguslZTncXrVYKbCY04QQVkrJ
yS5ycJRAjp+iKRdj1xdnmmtKs/LnMGGWxcLYVG9mOukmrql8K7sqUvVDaX7HQmQw
OyODhIteilkW3Th3BOLl/IL9ZjLN1zZRUfgflOo9P05o3/lhsEDaPizHdKsgQyoa
5+iYLziD6MVDdkJTpCeGQ6kUeCXMZEArHzppE3uPEm3LfKzSfJhHVut7rDSAAJte
9BnNVgmAvDQJRFxIe+uL/6nqCCDg6RxIP9o5KpC9pBjZzME8WBDyLjuxfLSQNRDz
MrkjsK2SL3tYTgWfXOtgaTEwoJQEcxebfPC6IxrM7RX9KB4XB4YXNMT+jZOrFcca
Cv1IUNfEOvPJLihUl8rpzG5KKnc/1xF3Y8PkXAYOCDj1y+otnvpJ2Ty9spxTFAo2
oLJvxM+S3Y/FKBUQWn+ko0il6krcFTo+6vuWXCMVFNoJwMw7cWxfcrSEXNq0JDWM
rI1+vR1OsWGs+lyBhrt9x5Zj0AmUG2EjisVX3PIGmeTq0tgK8gtHk95/FzkP3RDE
VJ/MZQk0WGjiYJSDFQCL7gOfJdpoXAFKUBOP17tmXeSRn4u+Rl2xX6v2wQRZt965
o4Z8tzemXrPzF3/QinCX0a8xbiGYmGlJedqZf96Ue2DM/5pNbYkddngjHb/pP50H
MEBWHwhZwuOiYjtyBMxs5OZpu4fet+XMDmVODtYcLepkTwDW+q1jgVZeMqfXcdIj
KoVJ8Ypimxa9ECc3TtA/mOzcxoMHB5SQCLXchDX1QjhqY1ngddkmXMOKPNpC4XWa
w2HS8Wq9yDbKqMpVh/mzUPgHcb7suDPaQNV4Ef6e63PfIwvUPg+mFynSnTaDzPwV
JnNh9pl069ZeKn1apaOehoRQyLCrdVwGhNgscnb+4BLz3grehvT/XWxHcw1NbHt9
YWEd9spmSxdRGj7zow6Sg+JACxjgaPlhZj2lo6JKagvwkYHtmrGV3rAa0UAFUygP
x3h1LEjlFCAxBzwPnKu9sBRa0+SZlFrVcXMTpovJKvLiuJfAHa4iyhCrmLzVXoRy
MGeNnzDmvJLPkQLhb1ZqST1l5GwUHger66qU6zEJ0B/Gj6w9vK2i5cFUbpxAA22K
ijUxTcM6QIUdsfrxaHVvdJvumCixWwoV5lvZN1QHBmWC+ZCyvStO6Axm3wZtLnCv
AcY2j0LSlneuK4oEf1x3CHpi3Auugh/pX3zjauHTMXl9LdvkfV9XYImGjntzrLKY
nuZAtNRF3D/PljcZtofcPaVhpyDExA8jHDT1/iq5jJZY/LqW7CXR8lD3YJz7Ib3H
5Ps2OK8FSqIiqpS6jCjVrIyhR83DHdNxH4bxZFTX8/Q6hAVY5+YGsYYZH8GR2AVR
K0RZmEm82a9u9KJuNoUr7cbXKOoWkY49QagNq9kGGP0XqWKUIGD4B2TOg35X6EDu
V2a24GoO0DFVfZrYR7VcQ+fYboQbX7mIm20spJIPKYmywaRZUHv1cQnlQAWAfy5I
9Q8nmEZzRAK1bZFs6gYQLyvQTM03OXvHP4jqTrJ8ZW/00hXZR43MvlQjwxCOLS8P

//pragma protect end_data_block
//pragma protect digest_block
ouswO3q5jTTDLsr5irE8X4nmZRE=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_SYSTEM_ENV_SV
