
`ifndef GUARD_SVT_AXI_SYSTEM_COMMON_SV
`define GUARD_SVT_AXI_SYSTEM_COMMON_SV


`include "svt_axi_defines.svi"

`ifndef SVT_AMBA_MAX_ADDR_WIDTH
  `define SVT_AMBA_MAX_ADDR_WIDTH `SVT_AXI_MAX_ADDR_WIDTH
 `endif

//`define _SVT_AXI_TEMP_DEBUG_MSASSOC
//`define _SVT_AXI_TEMP_DEBUG_MSASSOC_L1
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
I4silBWw2pQddMeK/WVjr9Z9FW0tuoOUKk5KNHVzl1t/qFDGz6Oh43M59G0MHZmH
qiGRTMvx6fhONC8cx+p8eU+PGwog6rNIal0CDYecSVmgOHbC4czZbgd+9RRK1xqq
FS1YZBaQV2vVRUES/Z9tuh7ul5Z3Y2b3GySV5xfkg51ilRXBVTGXgQ==
//pragma protect end_key_block
//pragma protect digest_block
IRDV3hdBBAdp2sUbrsMSsLz6Pwg=
//pragma protect end_digest_block
//pragma protect data_block
yOfhwNeboCd2WHM0LPue1VCu5a/ofgbm3rNULluZuWQf3r/OP5fJtliI/Ych15vc
vxP5ENkUiq2BY3BafLtvFHdBY4UqY7Hs7qrlCE2pKp9yAd7KIk67qnBTpET41BFt
4MmuxiUxkPNTZcfyDkfcphR56SDG2d3RqPUtiYZ0/MuOHwMD91qQJU81PqIQVcu2
hjKNws0bmuNvB0conM9ZQQr9TTs5rKYgoZUkvfyZoXmuJp5fB+JtegCW/Ru5lwf9
SFNKUyWdDL0rn6QwrPHtDmsIN/JA0Dv/lMiZMiadjdAwtvZWy28xmE1vD7MtMeb/
T1Bc0GyTRrcG+TWTQy2dM4ANGlSBlBkIaM2Gq/oeZm00zsK8oWrPxIbom8gKOLZ2
Rmo9FkeTNahaiP7dtpGJb/oizEj1AZ8Sr5DA1OQVODTep0lKyWZHpDtmsejtiRPE
OBMEwrB1Xnjz04ZnPQKNQ/0D8jyIy7JhUCMLwnKPtnWOMz98MRP4XuynCT/rRuLL
GOqs10x7QX5PWPhit9fcNIyoqdvmJ+W4s5F9jH4sSU21tsS0eOEsLO7OLbBvTM69
jaQb+9XWw29cf9Oc97EedLnJFiQyzys4bStkottDjVOAz/XulRpwttw2XaqUKwtW
AwlbCzjg7j3WtdtoFowSuemvayBXzW3VHmfQUkDukhuMqQJHF8Rc7b6RcX7qUxot
nT7GRIT1ASD7Ve5FWeVEYyokQwHYSgdpGiYcs8IgBSjlCHXmii82I+DY9/SknF5G
po+JjMst3nC8n1ejFgl1WCJCx85L7cJlxbYTuGN5t1uxPAZcYdxDB3FbPsrnAJNj
nE4McwTnWGRrYs5gU2iDJfT5pDQtVeDZLd4nPqmqf9Ksn+q6m1B/3FqW0uvsaaxO
CoMdvmS53Vf9AFbWRd1ydEkLwJBV2n/ycScFhiZk0w925HtVP94xoFpMs54WlRJ5
L1JglchkojjsbfKhiTq1br++E5x7/cCv9sLKkhS7We72Z3Di8LYh+yn2GKm8osn7
a2IqVnLA0uPI9slQygTpTx5NfOcH3LONA958Cgt2xK+Jrr1dtgsb0dRJjOQGojl1
iIp3fEmlYAJaepvF8mQz3DIrWzQl4YGxy82Mic0OPrxoihOgHCLzB7BViWljjxnV
RHP1GRXaQBUIgqh3bzYhzgZJHQ51S0WIADcR5dC8RWyhyUX1GydbDMVXTkDt/Ps7
5xr0Iozgj1VGP/N9bSnOIvzl/k9Or+n/wdz/tTgzEJQPHsT2PCb8qt1/YA3ivEES
mH7OE+WSwsh/WJ+T6JKT9URO8wbyokICAO40qvJR+Y4HCGBLi0/sFZd0VUXYbpx6
/3NLZKo1NEZBU6WRQQpIYBSkzJ/bXkGVP25JEXNjMDkZ+6dKFAwEfFvS1QzSiFo9
XPP3epkk4w86nU0nr7v61/+vsXbZFtrOPc49GkOSRnP8NZ4eCE/CkNkMEpp2ksZY
W1bIsRfuhXmq0mN83Vaa3szfyMzoHhE62m0NEwgbl+d8V3xl3dgHcPbpYb5bP/H8
HQxHrkHDHIHNZYxcjZ1/RdikhpMf3QKbxdGx2uHvAmHpSBgApNStFJBNmD9arWU4
eoKu07ph06XQVHWsCGO4NPdyXUOmaOlG/upY7apkDrOO7gZ7IvU/4pdrWBdimG9e
gJYecA7nDM/1O+513Yive8SYB2q0380oU5F30HYEBLrppi1pPtipw+dwWR5ObRkS
WBL57Y0SEueklk5ONHuvw4nidzKy3PZ00bxeyYWMi+kyDnI8NF3q8ELBjPaNOcqQ
QqZZBSLcpehoZhbz7MTKxT9YW3N9yCISDriO6Z7jg87ryWJ50lWf8uM5jNTGxMP2
X9tHlSOIxCNp9pCd7pwBki12gx3TCFSVhZZ7gxvx7O1m+o3d8xXg+C7aahqJwEeU
CesXyQHyx+eo/bmVOrDhf72NjnRW7uBKt6a08Y7hbPjuEVO9uel37HX2VnOc0Z9q
POmlCo2Q6dVAPC9rP/SS5MPS6CwbfDmtRh9zj6q3oJ0yMIV6VYqS8dL3ltDUOzDK
J8nqIkuoXXlws3iMYliE6kmcwo9e2SZIhSepPEofTllvcrPd8/6BG9G/2oYPGP3p
nIL65nTsBtksuNnl9nJbDrMr8vzZvfE0DlzXTM/RB+Cah3W1SIhHAjMBOR/FgCT7
jciD01Di2XWd8LrObMM8USK6vqBlFQIsd33prwguiEccw2qWZKlO+C9+jYpZE08M
3u7bPh26Pc/97kOLBvP9WGf/2xqofX7sT5rk18F8sYQwhUSd04fdCJXA6ypS0lLV
IqvYQhni1WSe89RQOHU4sl9HpdgPhKE6CDJNqm+10eiNAJlj3081+usUaQLO5uIz
mG5naph8ELtzMWEW23/JUf0t1IhxC+kHD0hKA+Vw91Zyt4LH+y3js5IfreySb+/r
tBiFL+z/229VDiowDe1FO9miOWrFbZOIOjRufe/KcYsPO4nzYX8gxHrYzMP/OgLu
nyxNNplj8by+FmBluveCANwMQZfO3M5sUCO63dtvcWym4ZNiuHgxqJTdYBOAl4SE
rJzGuiJ/Krml4Ds2azehEiljbmgNZNVtCRZupRx4+y4Jf5zpPn4NZ0gY85SkiP13
+meztaVdtyjoF8v2JkHRcANTOenmHJo9HgAA/eWhe2vimBSGbp1tAnpcJhjNHfAN
z1QL8GUjZ0BgHZv52A1FmS2dxdQK3gDkpOTrTcKpRAMPEMP8gb7MZtNtHOijHsFh
rcGnwkJuJLE1aL9JlwnSR/qGRahRXjdWODZiqSNYDY48XBfnTVfdG5l4M849Cbsd
AYEYLy92O5D2ZuGNBw5w5t6ETwyErxYtMVE6FIB93h3ERUfR17sow0zGXyenfcmZ
WMoFiB3sMpBZr2TxrainOHZCs29KU4LcTf4o1clZ5aNPYJSod3i5Z82W/gY4rcjK
EJ6lYohijwM2j1/AqDLAmg9jeJWJN/R3mf1gl2m/HwaKfrQh+AA8gQduaD+zwAST
c4GAA6DfnmRq3nZEWN66Kl37Sx0R0ny9rKbvSQjQMUHYAjS1wq8LOKBs5yzfumcv
SO5Q9/7S5SxNYcggPPL7YLIiWW3sZ62IJ40qztsvWCCBffGjr0Qnw+ySZf12IdvN
Iaod/+tV5dt2p0m8G1y+xb2k8VlFnUaB0cJx2wQWucnASzIFiIcuryVkSfCQ99mA
DcR8WWQFSRWEhsqBL+STgyw09q6afwAgImeXkTCGYkWqyxC0EPBqTeAuzcq6aO+6
UA7rvy2dJ4lRWwWo+DupazCm0giLWztWOrHHMXVG4HQziZjB9PLooU89ofVAYfEm
jCYzWlVqrN5JLx6bjzk2sht5c6WLmmugAOPc5oXVKD4ZsDLKkr3TsrQWrhLnyOzj
lhkunFi0AIRSi0afAGIcCs+9YtXX1us3PE1Z9XXBabRVhbELTMx9gPiQIhxJA+uZ
kEdozy49syd113DjIqYyaQDBwcuXQc3dnrAxgEhisesX6J5diIZVeKVGzipL5JMu
NizfZUk2+/rrIFGllUv1EtLa107UkhzK28RiqOeQGCVhvopO1JGeFfNkT0sU0P6T
T00g+C67H89k6GL97xEzPhBfyudH8+mGPVvO0DvYNY72TP0oBrqC3rV54cJPj8cM
lASItmouQUyHo/7FWl9ilYwm4U7uzsOQi0Q6d3LriMsVmwMB6HheAdlMG7QM7Ei1
YGHx0oIQjCJiRCI6pmWckP0OsLmDjeZc1lsRFrdq9rGrS/JFbX5zAYXDKUrYThLJ
eDXu6h6iA72m1BkQvoNT3PZBFKM95rLOKo4pCQzI/zr90TjOatln+5QN3xUSMmHF
rtoTssSWYHDuql2QGocCxFnM4gZ5ekELzMHf9tTa+LkhlmA16m1DR7ePGYuSjO6C
bdrOfMugjcNOmrsEr3RNRuIM+xv0K4GFd3jlz8y4K+OY45zKzEnhImog7UE13OSy
jSRflu7gsj6JzJOOZw3w/J2HKskQA8+rBFCSeRLC4/sEb16TsC6gPG1dft5K2lq8
1Y8H1xmVD4mF57kwZibCYAOacAeF/8GVtkC5myrhebIDLqzHNgkXL5bBdGpR5d8U
LZLbffK10TYk+TZb1sztjeuUKtnKfhAaAGfWwOVcp9PHLZMHzMb6VLtKqYLrd4/i
JxU+KSMf8XiL3u9uiH5iT17CiuWfyEOiil9NWwM2lo1OiBDSygvWYIRXK6DZiVJh
yf6Ps2xCGuWbfl+PAfujbPcn+Ai6PNikGd7/iARW+Knz7F9927yuhBdACLhtO6VS
XwVPcR52X0GAFVLvfoxuJRzm5KnymJp8QvwzcP0rjNo92UEQ84UDrxaa6pF63yO8
qqv55DAjUott67e9a5rHqCl7oi9U11eEVkM12Wx0VrnHpTRMrknuELlfgFlDzOLh
Es9ELT/gtPby22A/QLI/6eiKIxwKfpm/rBX//jf1LIrzxChQc8zMiPg17equdHir
69wSMfm14xEUv2brbO/mFfRB2PcazI9Kwzk9jIAc2g1IFbcZ2efbHzhSHQS6OA0Z
XE2SWDKkvStfOu3au0OYukS82m2x4HfUi5qf92Ei0GJfRhS6eOP80dz1YLcIYqQv
W212eH3ZShivklca7gfB34pNiwomdXUEzfrVIp3XObJ2xap4pmEVRyfNXVuCwcP0
714oqLo7NwA5btJ5GNrc/YANavAg3nnPYjRmIB7uKWxXv+T5/y49L3XYttJQ2r2P
gpr9H4v2jwwANBOpI+PK4fhdQv9BYW8IEYbRymWYtxg/OVQBp2PPf7VuW0DTmYgB
zYHjQMFdYsRs8EFF3WxbBkxXOLjVAT625s3YbwG0txbBNFLAfMVvTJYa/K8j/fE2
gQMed4qezSBVhkH7Ck6YKqaOjSHH/MvJ9PwKzPNt4tShjGsn/VK/Jzw+R21feQXI
7whp4BEiJDY0ICuFBjpGZVFxysgXHSOb0htCfNwqbLlIH6njy7pwTneJYGuuHW7f
EsMoG6M6ao90tLq9oidwL2AmK5mqrMEMgYuxFyyqB5c033vs+7iKX7b68uPJ48B6
15B8UtXu2TaadXDFnKp9GMd59/dVwuop26oH7iZIrJId38XnGXj1hL5U5QiTaF80
3k2ukd9dl7mimh+XWmQgxY9yT+2+1VYy+Q/8Cxyepk3H4OyqZpiCXDMvpK4RVlVY
qLVlYZcJFFwnTIugndEaQU2epFvl1Ab8wxo1tMinCiMHAGE50A/nXPE689bFDxBZ
GiBLeIJZ1cg/Oy/p25Kz98h1Y0qH69a3BX3XdDl1j/LqT2hQRuDWujjencbMn1cc
Vm3ptRYk+MyGGjopc+FtoN/2uKw4/R6oHem7wPb5NHNoh5ruDXceEXSzUJREJT90
ms8jydTb9RyNHsHT8tFtnIc7p0MetLG19//50ra8RHg5Q7OnHTuCKJz+mhJEf9wH
E5uFlVFVNTCQru1Ucj17u2t/Ok7NGs0epJ7pSV064Sws3Jk4bvUBk5ai1TsPKFCI
FIyoW+m/o5e8gWwCgcwuVYbyFX1b9kZb58wSNxLPB64qW/5uC7at763DRVURKzy4
2JcuGpxRUGiFM16yDCSi/LYl6qEGNcyG7q2sNSVeeYZ9tRsHRhNGGnGKfRYIdtTG
tzSRrgNRTjDNWDeJf7Ydo0N2Ms7WL3AjQ8y7OkAidBtnY5JC2HsL3Uqc6tP+Ra7T
FDSX74yJwm7/PaqfIrF7bc/PA1iQI6NdVv1VTtwdFnuEy2or+03+wFW6BDS/7TrT
VuS/yW3/ZHHMDfjsUpjUeAMtRx3sJSiK0WTT8z5xmhCkQu1u7xxsd2iX2MPBM0TK
wOBrmD1da2q4y9ZIYKBaqgCe9EB6AYLOLc7Srq1Nm4EApIZdhcahsXBhdk1vIA/A
Lhczcf+5EIKktp8KsNYZvTxFoDn/6W46ufaUMgCC25SFe+T1lhVsve5uaqbQ6oAJ
1djm+a3Nfa+aNP4i8yUvlXhRY4AgQM6LeCW4eqiICsExxODLYhNhPh5ZjqPELSC6
DqXqmKtm/OCyJaAoKJjhQcBk1UwsnWl67KOGUycfLv/JwooRfjvc52BSpVCrJZHv
usyVR3em2AYzeknH/hvLjyU1W5aRSLWIf8rm5k94bHG+EpN0ZGXf8+qHksqtfnyp
ktBY9gQj755/lJ1EQyYw0dvk6Wi8Tr9TUcppkaTm8JgLslI1K4MXH+ID8RRi8FCA
tMugtNnM64Hsqwnu7sf4p+yy1jlcoFO+fzIhzQJLH5n87bM+QujnqHPC7OdRueBq
JcLYPYmhgIsALSeF75Ep//MBbX8vLkCS9mwBO5u5EZNfb0gzFpY7JxN/HKssqF9D
FtYlEI8eXSYUrSpaJyn/dLLJOOQuw2JUFMiUEpXZ7AHrtW7aF8A0GmXEhwIiaTee
4jmn5X4ARWktwL0+eksEg6HU+JAhG3Fak1qRUM6Ikl/F+M2F0FDzblrlpzJhZUz4
5ESv8NPQKxwseF4FinOJTDOonTqutyy8z9la/2GY+IO4s4nzQGfgIZ5loA7rvF0T
jWo4mCuOSTIdizzHnLl0S5gyw2DUt/0LBuWUA3Zj1LUgT2Pm2My5zweoasW0ot52
5CT9GcLehjHHzXyEa1k6VetUtOFKpF/DDyYHYKyibHF9zJHnUdLlMVEPMcBXgi0f
QGjFNBBzSGQwrL0cY4V0fFJdpfZIPzcy+UigvbB8RXAgoINCtVKCu69B8h5JCFqm
i1VFDnVb5hxHbD1MEcFE4mgo66EPgvn7KG4YSnuHARUL34KQjgjVGW1je/VaJ6hX
MLKOlhEJ0xCBcbciGmFuIAPbGbEFOuv6UwQlxEsMjQNBAD1wSLrXqGzDZTLAfsoF
5Nc/bnlXDD02GuK+XO/IV/RqI00yNSDvhQrx0DptOOSB6Em85ApLbcizt5dnQwCG
MWoM3zG25yjQGn0q4CEg+4wZ47LQBHllZPUMEZn47I3hBN2MdkJqsgdOim0QRRoo
WazOpA5oSJ36FedZKs03H9WBUiOSq9hqvIbzVfQO9hDZKhkHvc1X9uOsxux4rwY5
+lP16OKryH+4UoUA3lCmpMdxOmltmswGF2L3LG22keGOQgOoRLuQlLTqshNH7cqZ
c6PlkJ9QR6WGwqQZ21sgKrEEwlRTTLYHUihl1SlT27WFxIxP1czQ6By3u33GGhlZ
dcsfk/ncWY2G89GnVwrIhJoK3Gx4zElkSnK9QKo7ZcJo9B+URQFr5OOfsNkObmdF
wCZhMDeUlQaWfFfpRJm1VgjOmzopcFEbCzNqzPtmjYrnSparfe/nyrXVs+0KK2KQ
ofgu9XpvDT7RqdL/+9NQmS+qgWJEb8y/91OHkWt3c5XZaI6VIjbm0jeUsJU3mdcZ
FCjs+TY5WTKtCQq/htT4XoZtcseA5H1hg8VpzqO0/4NcVW3OV4GHnJRKjkKQ88+d
RbCoohjSER7RQxbuzGxTGnyzPLgFE3ufTB7oPjQA2ZdjY1PA3aaRQRJJgo4pjwLA
vdtE7I1Ga//AE0QAZT1/keI719UT9H9XwcIbQiIm2N6UxatR9lgpKmRUPQkAq092
hemy45fsPiCVdl7IE3DbMVRi+jtiXJhvvlvOPO648xfMieL1j1uT2DHlQPQZPw83
366zA7gJ9QM2mNptBh/GuZklbujbIlO65vCXFbD+ZKMyiRAHEqQxjGBLDN6NgmG1
RxYqW8EFZRl2cm/nh5hxnqrHOt3Gt6+weolD65md/LzCREK/fRos77uq/U1bb/pX
WrsWWFyjW4TNNydIRgK2oRW9eLAUXOqzolYWHtkjKAlugu7Ain24ZgSkFS95R7hc
QNijwof6pq4qqS3OtGn6tYMtbGtO9iCn4G+nbOE9yzTmDfBXuWI3JMu3aqfu2E5L
xMM0nifnG6jWMLazsGZtazkszSH/v0RStIjekzKW0E+OvovjU3MXKcsd5lOnF7MK
1yk0ANHAVJ9TAJwt+RrfvmYrY57o3QXOtdqaiRQlAOIpJdh0Bwl2+Oupz/i9ToB+
nsnnYIY+eHniXgT/zkLSI/sN4EusqzF6IogNOgcKpU0HqA8rEleIybeHIIgSJq81
mTF99FE9RJr4x/zkR9haHOaDD2meJrJfN7VUBbjv/1wpcTb+ishpfFKeYKQs6+YQ
lRdvDT9nA2Fnr495/ZoDAmKtHNfLpEU3d9Sch57Pq9CZkoAy5LqE3vSH+S1/FY3z
ErPE4UeZeaqNBcOtCE080eg1BHrl8FaoDiEp6XzkPhj7uda0YBBbVkg2P0RBwqbg
VRrVRDFjqJ6S/gesa4PLKGnlI+t5MPc5lzvVovw1A1CxiJxWwwuAOFrCozPz1jP5
9JMjSFYevVUnUnaaK3a6tKeCmZhZW8kpFRu5QkX0lCjzSjpVYxjfXgghzjjrmeYY
5OKH+JPf9wNfGG61bFR7Tb18IKI3QLHveqT/XlD43ZJ9ohY5oAhOCX8+05Uh5Xsi
wr54+tIgfJ8WbZLqzYi679mXvl01lyx7uo527l0RMrH/jFi4BbkGKwDQAKHp1gG/
v/mn9HaNSGGBFTGYkINRpwoZKt8mpZEeS4XqCigN0nNlsdcGu6DboI8Cb0ndvUWv
07hpXP30ElH7wqW/cw2+cLRspnURPWrJhRasp+nfyUT5X63r9rf8ROizy5H0ziss
aONIHIwu5LRAmREj226XR3YiyRj8KhnUyIvX4/YBmRPybPisTxGF/4sdA/GqY/s8
3IXZLsnx/TZUmOiS43SFRaRELU6shn6o6DxxkpEkfIkOTz2BhW4UPWM0azg56W4g
iK935YTZJ2e8a1NkF4eFB03Og6eQAq9kKQkd5JZHKAkIL+XLjneEkPX7wBySgmw5
Nok5f0eOtelVevfvldRneHbaTj2ghbMNFxpoh3IW4dAFvnEbZHuOmP0LmIPFxFP8
dpZ22DPQNRJ41GVyQ6LtmJx+9/EF1GREDb7nwaVzhQbGE8LRP7RpR42SsnBY1utu
wHffgoJmkQpl4PNDOgNb7sivUkgvM5OtweIBAp9UG4CTMF7CPyPgaoU0z2qxvzHB
G4ZJOU7/oxsCMtol3YUMrk6XCuv1noqHeRDGXRj+pRAZvxceddwUd92ReR6OqNsU
mNqbu8UnAXsZV9WLeYaMK9lj/4Eo97AsLKF+Ejylu7PCskhIfdzdoIdOujtqEVLv
9O0B659b3yi3HO8QQOn3BN7m8G/ha74pTIIVKNXtaiPRrkJT5DLhMGqe/v5rskwI
qxgJlb2ySBjYfbLQT2IWCPit4HBsZ0K2pYd2EdcvWLVZE29l0qtYlNJxsqSEtfPa
RWFNiJ0EsPaFtV0DsUUCckU+IWuJ2ss+Vn2kaHrvhj0ALIRJjLliEyYS21FxsjIS
7D+ji4LW4K/BNXJhESaHw9rND7JzZ4ooPO4tyoVSA1o8LwvVVPX7lAL7SnHwMMkW
Ovv+EQhSML4nTpkA8mq28m2XtvlXGzoar6mtjiWGGBKC7og1pyFftG7/e2wvlXlJ
XRoyyTuy1oT6ejFLoeyJPDFCDeXx8SpQXyEj84AOIhP3S1b4+/xuTK45z90/gblz
zchZUd0A7wmJyM6PRbboPXUigz89JZxzoVy1R8zUW7R2F+MnANM+/duAoyfjaZFD
9KqB74+TyNz0BoR3YYRnIIHhIw/A/YtE3qsbbsyJIMK/ee+esu4mmcaVBxNyCp2V
cWTqmrTNQ/kWeQ3Dzn7llINLhh6B069BikbpO1sEyB2qj6UHylSvro/LDCunBFPG
3bJEOLWOaFn4rU6aUDt8/agJ22hAFeRzhIsUHJIHXdWOUoz8h9my6+HT/3PloD/X
8J7xwxXVgTIYfX/cP4REwB2EVQrPDeObVkUJGQiKTg7q0MOr3Rs0BuW45eAchdX0
heHu9rcmnawov9Y4TUd8EWci4P1B7G+EWGNU+i1ehslT3f1a7HwhLlSOA0crpqFM
w9XujlohSmSPXNfbZ8+Adfp1lOw85Zd7Hb//4060lamXZya7VxeKiN16i21fLdPZ
1N9rF6OmfO6RxAc4h4CdRrw315qu94CPJRRrOYRnn2yrcKOnvyqgiP4hFNKQas92
PubdGDist5Tryd06uyxZgqPMMzVHTtPu1c/GEjaGi1cKxOBUoTzwxT7Vx2lRbqSE
vUJqsOqKNguHJ8FP4lgFAbmx6zoCSMgdJheosreQDIz3WVcjqVtoS2v+qjEQ7hex
6f1stH/6bJSpe/CnymXPvlPGsdl1C6n0tx18+Q5IX5Exi/iHsHyXN1XVSButmLhZ
mnjoBTrPAkTStjvGJ3CBMpiYSxHCJnboTz0w/cCsa6l1COl/1AXMUtwuvpqn3MBi
kO8nBCFopCQOhEnxB/8zL2s2BE0ZjJKYZaa+QKkvK8F89kQGzcnDVVg96K7hIuaU
0jgBPf6pkWr9sFRxB/6f3JCFy97CgfumlRa39PUwZpNXsfF/44JiQk7Rwpa4tuYV
nFu4+FMhP96OJwofNwnkCrsz6uvoaRpeK9L4O0s0TQiZ0bUEMYW5i9k2IBgHG99a
wvoCotFJ74gcus8FptV7iQqUAU/3fi6Oar78oEe6rWPKFi5N/W+9jsdVdlg3NINR
U/N9ugNP7uJJmcPi365l664ER9bb3Pb8xsU/awbg1TI06ezv6SERINlz4KxXjwBD
rzVaIALF/yZtvQlBhUmrEgAqz25+gf+r1t4h9k3y1bjuqF9xkDiKqMqFAYDoQAry
jUFcv8IaUDjfW6RfryR9/4EtDmYxoHS0LZBBTCeQ8XFPmDGnFI3eiTkO7oPUqth0
Au6cHP9w+T/wd0nkb69+V8+YHziJ7ankNvuui8gKlvyLzsR7je4LJHugV+lSJhBe
Oflk6oUnaPCnqwftuVAY3lYDA4ip4I/MF/ICgZNlBFvTH0qL9JrmkRxQL+oCKd5T
nJk5wuIrHc0WkG0h6ZbIrpi5BRMdKYEfTXj1UX5jI5g6xZ91zdkjOm8x3UENWFZW
Q6zD89gXMpD8nU7iyGx1j56C7B+n8TrqloDIAg1sbmFHiepnu6mV2vMddAkJwju5
i4sNxQsP5eiyOpBW6ZV+pRznQWZUWOfwExQIC2fG0iGJEfALxPoC4sggIhg8t3Qr
2/CCysIcjnD/3/DGVhSFuIupDK7geNIFZdz1fhY/yjud4rhvqJfVB9QpoWO5SKRs
lCPT3QweXYIwOtJwsVCVhr3d7v9uomCDHAYArpuaRpxHBHcHd+2412CCLdn8rmjb
ixg8bgvpKbJRuCfO5n+TcejjTEPmXAFLmjfb1ksNlMDzg1a7Ny4q69ikD4CQuuX7
NpNFRygDmow8aWXjXqA3kaYa5SmGsGnwvVLYlh1lP/bmmNa4gGoTKRL6NUIaVHim
vNJgbEkIkcf4y3wrA9MjbvpkmjMBDIPUKXSC/9g3YkSG+VltwMpSNh4RWlJoxFqF
3lMvYAh58oeDCwiT5RIkmjrx1t1TNZ5QUz9s5eBUD+ynOjQMR+iiVFRsyZIGr8H8
2GSIw1rbyRw6zKtaWMz/PfCmlTjrPHlnv6F5DkC18kF/AdgFWMugp6NveyATUfLB
q0/Srq+GtuqxbNavPBh8P6L9btRuq5hw0xA31UG+bD0myDjRpgCPZizSrzONHZjp
uDEYD3sRssGAiihf3SlwL1Jv2ZhvyYKsICmn8h80kLE8UvS3Zt2x4H9p+GLqNHkw
fWsUO+cSgTQXBYIv2BsxvJagYpKuah5oH9/RDlYftBde1SrEqzme54FpyIIhjDXE
EzJGq2npZDV+O9UVm3+lV0ECI2d7F4LytuEB+0TAHWuIFmQNvx5iRlOwZc8mxfsw
qPC9y60LamqN+aAntGrnxxmUCDKmveOJLO+lP+opvePkm1dqjq3jinrllxxBIk/I
m2/7PxxnhAxqlGd+UxXw9EaDuYzpylIA3VP6zVCAo1EegHvdjbz8fCbPygm7Msa+
CQ+0vRYPWSpbHBE1znxStGYoya5p253IiF+Ia97qz3hk2xETwmYrK/0eImureG9i
0HtPwzgr/GH2gbb6Zhm3lw3LCEqMnn1gc4ch50nncXUYn9zoBp55cyrOKtrX8uQy
l02vBpRmF77ZcNLKTA19Asn6PhXqSCsw5uVhg6txq5XfdtVdAFkJ4aoZA8vhO0Ku
i0Gx0VUFUO9fq6O0rhafqfoJUzSlMteZPhtf9hYicbGpEMsLds/vNuh96bNMK5/3
/w/x0++RfEfeK3nTezKl98kWTopKtvYHng+8m7DrL6sLl7ssbP02z2rlPTmMvdBC
l00yAtfz8QUf3maox3vcLMgsogQQk5EypxWwpx+6YMfR93AXxiyPgLIQlzm4R3fo
VcQT/q3mq3cv8CMLdANMdhbI651OoJGEJbggYSnjxhb5WSdIv0alF3ftiqB2eF5w
ynOg7aed1LEhhn4vm6+C090laz6zEDZ1kukfG7VdRTh8lyc/ksx3tKiUcvVQP/5V
iVlfcw1TXnb4tJg4lNrkxHBUM3XHCkq6MFUHr5H+oXcfPMMc4PvjytTjHmGaJIjh
qa3ZbE/58kA6hxUhMZfShHew0+/kFCrGWD4U51c6f/11yzLwgQ8iIsJz8WTKI8pz
3wu0lUbflMsC8ucIen4gZIJUN0iEkFu91f9ba+HPYXEFhw3rSQ3yy0uAJjulUF74
DxDFhPCHOZTaIHZJcXJrPGm9hpIbrXt4wkuAJfVRWHWL2vdgxvgZLZXOjBKb6R/Z
8dP7KuPdzmqf7Cwm6XRSlPBrZOwLCTlzk2AZUt/kBypFiJ6B7N0onl0t+C/sdNWU
6nYTUr+NXXnLu9TG7VYFuD+OZQjCXfgeetoLxYz5SctheZBWuNC6Tu5qS4GcHQNE
ubp7YYeSjt5BOdPKPNTwOpaj373XN/i3vuDk4ECmiNungTuKThNL0tqGObe8oyjU
yVzoD50Mf7NmPECCuvsfCXR+fcQhwPSCx/aJNdMsgi/LQpr1zkINaBoGJXYCGHEQ
BVL6BR+NpuM8OFkBLetHHlVdhbLIF4Bk8pX2/90ikfDsOjbM2GZ8oCAVEk7eqklc
Wi9+I5vN5h6ta+3szFhNLwmLNUJ4tyQryMlDU6tQNWsITFvA5UWScX+tpel0B2Ye
v/5268IMdXEZNSbs9UlLXgbY4iaCdrniZQGy6mjL8YyNFKKU2NfmUy7/Igj3rOXj
dntmJScrTgYJBJOJ7C9RkWgm8vjgdFl5Hoys8tlgUlJDdgUvXLA8X1QgfN6SqNwv
CAFs9z88soqBypCZnGNrKbwStBqsjzquq6klq/BAIny51zpfhR+KlbBhqGaePydX
1gQK562FKVShyyNhSI4RORcbhC2CKWQLhISG7SN3vI9EalXn0GhCqUJGJhXay4Xf
FV1NzfxOw/IC6b2rfgamh/Sin8dRJffTqiN84hHESQOQI9m6ndIBYPqz5GFOyUxy
J31Hu4QW5L9VpPlG3jJtPYLmnEw/EAcAp2aJphZCMMcOXO6Nz0q8d473p7hjKbba
iHeog5j58rEojWFqGFIQpCcoX/jStLlZsTmNCNuOOqk4WgLxz9UwC7a4YpfKIcOM
sI4YtB6Ftg2//baY5+LKrTEgmHdAzYgpWw3QV4oPie3SCUPrCLJku72Z8QFOBdSK
KQmkNr/DUfL0GvJ7Jtd/tvbueWHSNiNhDOQcFkl+bpgZxMSgkLIgu4/n7zi2RRjj
++DV1kS7jQhRqmn2gZeP0WxFAeKzBjuv+jgvK+6ETGDvhMDCWtJdXkby7CSl6+rh
a+KtAbtg36I3rsA90BvvYBOoZP+CMMMYgYGCLM3RUSPiJMinf05O5/Zh47fg+8GH
5eo4SNPs9ddJpPYhwtL8K0soEJurYlNxYXffv1euOTbSupDvE8yD6atm6XB6d9/M
oKpJVxmbM5mkahbTim9D6ThOjXs5/g5K1Tmxf5MiypFDP4wi/DGEaDiz93lBexkD
mAwVKnqtK7TvoI6ulOKOIDdf2Nqf/E08vOiW/q9+vvg87zBjsnOCVU6kDUMn53aw
tKb4+pXmZQkjXdzI9KlwF+cxXI2iQN4ChdF3F8woHZL5V8KEOV565zQsFvhwyqv5
ZXhcTjL8Owzw62G+5Lnb4NDUwC4X5E8wSr0yT9eA0rtdVfK7HddL9Ncx/hkYzkpc
9FuecGt62GNCtBCku2/LQqLkT5MNXVh/AXe/FXPvzkZh+9q2Fk+tkQVk8KOpBJTj
DrGBSf9BzQXNZlXVxrcWjqqGmg4fQf+KFn9eU+lHp7XaomLmBwaRUvQwaT6fjGZi
G3NK1AljREF2faA2oizv0n1KFvGYjhkIHXwcb/HGjED+SGl8EnQDs7voVu21N+YS
DOwfyvivA9tfRhRNUe/ldpomn/vFdRNiz1OovmtoJ0ldQGuZdiZkwnJ74WGyln7P
HEfX7QuuJv7XsY+rdZd0TxhGt1Pctb/zAX4Os0PAi6t3V+2vcNEiTlDUVhCvysPr
Shp3HdCVpnFmZwihVj7GTuaABfsAx8eqD7gh81uL0quqExWzxGdSmCghFT5PtnyE
8pde5Nbm4I14CdUO4T8NmA==
//pragma protect end_data_block
//pragma protect digest_block
It+C5g+/CFaZzyZnALbshA55AHw=
//pragma protect end_digest_block
//pragma protect end_protected

/** @cond PRIVATE */
class svt_axi_system_common;

  /** Report/log object */
`ifdef SVT_UVM_TECHNOLOGY
  protected uvm_report_object reporter; 
`elsif SVT_OVM_TECHNOLOGY
  protected ovm_report_object reporter; 
`else
  protected vmm_log log;
`endif

  protected svt_axi_system_configuration axi_sys_common_cfg;

  protected `SVT_AXI_MASTER_TRANSACTION_TYPE active_master_xact_queue[$];

  /** Internal queue where coherent transactions to slaves are stored */
  protected svt_axi_transaction active_slave_xact_queue[$];

  /** Internal queue of slave transactions that got an error response */
  protected svt_axi_transaction slave_xact_err_queue[$];

  protected semaphore sys_xact_assoc_queue_sema;

  protected semaphore slave_xact_queue_sema;

  /** Semaphore to control access to active_xact_queue */
  protected semaphore active_xact_queue_sema;


  /** A list of system transactions used for mapping master transactions to slave transactions */
  svt_axi_system_transaction sys_xact_assoc_queue[$];

   /** Internal queue where snoop transactions are stored */
  svt_axi_snoop_transaction active_snoop_xact_queue[$];

  /** Internal queue of snoop transactions to be deleted */
  svt_axi_snoop_transaction delete_snoop_xact_queue[$];

  /** Queue of transactions that were a result of back-invalidation */
  svt_axi_snoop_transaction back_invalidation_snoop_xacts[$];

  /** Reads which have an overlapping write during its life time */
  svt_axi_transaction reads_with_overlapping_writes_at_slave[$];

  protected int log_base_2_cache_line_sizes[];

  protected int log_base_2_slave_data_widths[];

  protected int log_base_2_snoop_aligned_sizes[];

  protected bit is_amba_system_monitor;

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param axi_sys_common_cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter UVM report object used for messaging
   */
  extern function new (svt_axi_system_configuration axi_sys_common_cfg, uvm_report_object reporter);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param axi_sys_common_cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter OVM report object used for messaging
   */
  extern function new (svt_axi_system_configuration axi_sys_common_cfg, ovm_report_object reporter);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param axi_sys_common_cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param axi_group transactor instance
   */
  extern function new (svt_axi_system_configuration axi_sys_common_cfg, svt_group axi_group, svt_xactor axi_system_monitor = null);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE
    /**
    * Checks if the address of the given transaction overlaps with any previous 
    * transaction. If there is an overlap the transaction is suspended. It is resumed
    * only after all the previous transactions to overlapping address is complete
    */
  extern task check_addr_overlap(`SVT_AXI_MASTER_TRANSACTION_TYPE master_xact, string master_requester_name="");
`endif

  /**
    * Waits for all transctions in overlapping_xacts to complete. Once complete,
    * the suspended transaction is resumed
    */
  extern task track_suspended_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE suspended_xact,
                                   `SVT_AXI_MASTER_TRANSACTION_TYPE overlapping_xacts[$]);

  /** Indicates if there are any full AXI_ACE master ports */
  extern virtual function bit has_ace_ports();

  /** Gets list of system transactions where master xact is not fully mapped to a slave transaction */
  extern function void get_unmapped_system_transactions(output svt_axi_system_transaction unmapped_xacts[$]);

  /** Gets the list of aborted system transactions where master xact is not mapped to a slave transaction */
  extern function void get_unmapped_aborted_system_transactions(output svt_axi_system_transaction unmapped_xacts[$]);

  /** Checks read transaction timing relative to the last posted write transaction */
  extern virtual task check_read_timing_wrt_last_posted_write(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  extern virtual task do_master_slave_xact_association(svt_axi_transaction slave_xact); 

  /** Deletes transactions from sys_xact_assoc_queue */
  extern virtual task delete_from_sys_xact_assoc_queue(svt_axi_system_transaction sys_xact_map_queue[$]);

  /** Checks protocol restrictions for non modifiable transactions */
  extern virtual task check_non_modifiable_transaction_properties(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Checks data consistency between master transaction and slave transaction */
  extern virtual function bit check_master_slave_xact_data_consistency(svt_axi_system_transaction sys_xact, svt_axi_transaction xact, svt_axi_transaction slave_xact, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id, bit check_one_to_one_mapping, output bit is_resp_mismatch, output bit is_dirty_data_match,
                                             ref string master_data_str, ref string slave_data_str, 
                                             ref string master_wstrb_str, ref string slave_wstrb_str);

  /** Checks data consistency between dirty data of snoop and slave transaction */
  extern virtual function bit check_master_slave_xact_dirty_data_consistency(
                                  svt_axi_transaction xact,
                                  svt_axi_transaction slave_xact,
                                  svt_axi_snoop_transaction snoop_xacts[$], 
                                  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] snoop_slave_addr[$],
                                  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_effective_min_addr,
                                  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_effective_max_addr,
                                  bit[7:0] slave_xact_data[],
                                  bit slave_xact_wstrb[]
         );
 
  /** Checks if the given slave transaction could be a duplicate speculative read transaction
    * This behaviour is seen in CCI-400 where two transactions are sent for speculative reads
    * one before the snoop starts and one after the snoop ends (if the snoop does not return data)
    */
  extern function bit is_duplicate_speculative_read(svt_axi_transaction slave_xact);

  /**
    * Checks if a duplicate read is expected 
    */
  extern function bit is_duplicate_read_due_to_overlapping_write_expected(svt_axi_transaction curr_slave_xact);

  /** Gets reads with overlapping writes at slave */
  extern function bit get_reads_with_overlapping_writes_at_slave(svt_axi_transaction slave_xact, output svt_axi_transaction xact_reads_with_overlapping_writes_at_slave[$]);
  
  /** In case of WRITE transaction, gets the number of bytes written into slave memory based on WSTRB */
  extern function int get_effective_write_bytes_using_wstrb (svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact, bit slave_xact_wstrb[]);

  /** Updates the number of expected dirty data bytes for the transaction */
  extern task update_expected_num_dirty_data_bytes(svt_axi_system_transaction sys_xact);

  /** Gets the associated snoop transactions' data as a byte stream */
  extern virtual function void get_associated_snoop_data_as_byte_stream(svt_axi_transaction xact, svt_axi_system_transaction sys_xact, bit use_dirty_data_only, 
                                             output bit[7:0] snoop_data_as_byte_stream[], output bit is_snoop_has_data[]);

  /** Waits for all the conditions before a master-slave xact data integrity check can be done */
  extern virtual task wait_for_pre_master_slave_xact_data_integrity_conditions(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact, output skip_data_integrity);

  /** Waits for slave transactions with overlapping address and which have started earlier to be correlated first */
  extern virtual task wait_for_other_slave_xact_correlation(svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact);

 /** Waits for slave transactions with overlapping address and which have started just after this transaction to be correlated first */
  extern virtual task wait_for_later_slave_xact_correlation(svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact);

  /** Waits for transaction to be accepted */
  extern virtual task wait_for_transaction_accept(`SVT_TRANSACTION_TYPE xact);

  /** Waits for the address related control information of 
    * transactions in the system transaction queue
    * which were started before xact to be received
    */
  extern virtual task wait_for_master_xacts_addr(svt_axi_transaction xact);

  /** Executes the master_slave_xact_data_integrity_check */
  extern virtual task execute_master_slave_xact_data_integrity_check(svt_axi_transaction xact, bit is_pass = 1,string desc);

  /** Executes the interconnect_generated_write_xact_to_update_main_memory_check*/
  extern virtual function void execute_interconnect_generated_write_xact_to_update_main_memory_check(svt_axi_transaction xact, bit is_pass = 1,string desc);

  /** Checks if CMOs were forwarded to the correct slaves */ 
  extern virtual function void check_cmo_forwarding_to_slaves(svt_axi_system_transaction sys_xact);

  /** Executes the interconnect_generated_dirty_data_write_detected callback */
  extern virtual task interconnect_generated_dirty_data_write_detected_cb_exec(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Executes the master_xact_fully_associated_to_slave_xacts callback */
  extern virtual task master_xact_fully_associated_to_slave_xacts_cb_exec(svt_axi_system_transaction sys_xact);

  /** Gets a string with short xact display based on provided transaction 
    * An extended class can append context information (ie, the source
    *  of a particular transaction
    */
  extern virtual function string get_xact_context_str(svt_axi_transaction xact);

  /**
   * Returns the requester name for the supplied master transaction
   * 
   * Note: This method must be implemented by extended classes
   * 
   * @param xact Transaction for which to return the requester ID
   * @return The component name that generated the request
   */
  extern virtual function string get_master_xact_requester_name(svt_axi_transaction xact);

  /** Indicates if a given transaction generates a snoop or not */
  extern virtual function bit has_snoop(svt_axi_transaction xact, svt_axi_system_transaction sys_xact=null);
 
  extern function void print_debug_info(svt_axi_transaction slave_xact, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_xact_id);

  /** Gets split transactions, which are split at cacheline boundary */
  extern function void get_split_xacts(svt_axi_transaction xact, output svt_axi_transaction split_xacts[$]);

  /** Populate resp and data in split transactions after transaction completion */
  extern function bit populate_resp_in_split_xacts(svt_axi_transaction xact, svt_axi_transaction split_xacts[$]);

  /**
   * If complex address mapping is enabled, this method translates the supplied master
   * address in the transaction to a global address, and then uses that global address to
   * determine the slave address and active slave port ids.
   * 
   * If complex address mapping is not enabled then the address is converted to a slave
   * address and then the port ids are obtained using the legacy methods.
   * 
   * @param master_addr Master address to be converted (can be tagged or non-tagged)
   * @param system_id AXI System ID
   * @param is_ic_port Determines if the address originated from a port on the interconnect
   * @param xact_type Transaction type (read or write)
   * @param is_tagged_addr Determines if address tags are present within the address
   * @param is_register_addr_space Returns 1 if this address targets the register address
   *   space of a component
   * @param slave_addr Local slave address
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @return Returns 1 if a matching slave address was found, otherwise returns 0
   */
  extern virtual function bit get_slave_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] master_addr,
                                             int system_id,
                                             bit is_ic_port,
                                             bit master_port_id,
                                             svt_axi_transaction::xact_type_enum xact_type,
                                             bit is_tagged_addr,
                                             output bit is_register_addr_space,
                                             output bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr,
                                             output int slave_port_ids[$],
                                             input svt_axi_transaction xact);

  /** Gets number of snoop transactions that returned passdirty */
  extern function int get_num_snoop_with_data_xacts(svt_axi_system_transaction sys_xact, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr, bit is_pass_dirty, output svt_axi_snoop_transaction snoop_xacts[$], output bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] snoop_slave_addr[$]);

  /** Gets the number of slave transactions associated with a dirty data write by interconnect */
  extern virtual function int get_num_slave_dirty_data_xacts(svt_axi_system_transaction sys_xact, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr);

  /** Sets a variable indicating if id based correlation matched */
  extern function void set_id_based_correlation_match(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_xact_id);

  /** Sets parameters used for sorting transactions */
  extern function void set_sorting_params(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Sets parameters used for sorting transactions where both master and slave xacts have slverr response*/
  extern function void set_sorting_params_slverr(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  extern virtual function string get_ms_assoc_dbg_str(string dbg_str[string][$]);
  extern virtual function void set_ms_assoc_dbg_str(string key_str, string desc_str);

  /** Utility methods needed for correlations  */ 
  /**
   * Gets the minimum byte address which is addressed by transaction
   * 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Minimum byte address addressed by this transaction
   */
   extern virtual function bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] get_amba_min_byte_address(`SVT_TRANSACTION_TYPE xact,bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = ""); 

  /** Gets the max_byte_address for the given transaction */
   extern virtual function bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] get_amba_max_byte_address(`SVT_TRANSACTION_TYPE xact,bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");  


  /** 
   * Checks if the given address range overlaps with the address range of this transaction
   * 
   * @param min_addr The minimum address of the address range be checked 
   * @param max_addr The maximum address of the address range be checked 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Returns 1 if there is an address overlap, else returns 0.
   */
 extern virtual function bit is_amba_address_overlap(`SVT_TRANSACTION_TYPE xact,bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] min_addr, bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] max_addr, bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

endclass
/** @endcond */
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
oSTVYJLr0kZUC9AvKzaCecH7UQVPiQRj0eM9bf8zXVThYshAsY2AoIH9Ri29CCCv
wGXnx7BKkAfJyF5J3ZaXu1XHh1oy70knG9+hd5ZzGD21S792ww//xFfw7HRiJVFu
nguJLrlDCjyrkDDVmo05zULltKmqWSy/MWFWyE5sNImFDJ1Z8EiqQQ==
//pragma protect end_key_block
//pragma protect digest_block
qndinRa9wO2/Myk29HrJGKC0wv4=
//pragma protect end_digest_block
//pragma protect data_block
BX66gpuWuowFCNrQjAWZ0CvxIA/wHr0gHCvMpWuSc86QH0tWgWhXQsG72nAX66yy
2m6kQ7wSWufLmKsL5jKn6H3vJC9Z2OBfaiADLzmR9QtkEb6b1B82PfJNOijJP0CF
BDgkdtSUX6zBSAbPr47BSfxvPW249F03i0TLHudQtLi+2dAlH5ARx4UI3TRinegk
4KkIiBqcpBZfyK4CTzEuzAfwBHbCDrkEODkItWDr7afdQVo42s/BIFYKcTZkryJ0
HGYktO7Rohl16YxSgyu/xJfjfgeT1WM0TIRM5RWcuPLrA2HSb7nEfHZRMlxCSogD
exsNElh3hmesvJD0ixOmOHwt3OEnTHIrKvJYZ3W4WcWZy/CrbUuuL7ZflFEkEkzV
ezJ2a0pLnRSkcrhv8NFyn9I3xh4ADLCqH2YdANKTimnpZFHsGx/XyS+fzjiWqBxD
7OTpPPb8Z4OMCU8vQyPsdW27xFvTBrLJXAx+hELbLERQhyRjgjTiGP+CjPtsBBVL
eRMuGbTJd6Fsqls8xhix43MAQsPx33tZqxYupgjl0EOi3q+lOx6doMK2ozENnt8t
nSL0Uzu6fo24srvYkHbpv1ixMKCqOOrThDShXb5VfPeygipJGQ4mTl9dMcZ2JGdJ
kza66DmZalGImXsuritIqCsnILz+z/TRU/nmN2fSbxwqyWjWg0R/ImmXGYRrsxIT
OSRA8UQz6nnETxYlAlL09uZtaXgKHjsjb5kyFxSKbddoxPe3QQXDK8lOrofNj+xZ
owSI6arstIRoVJBWEN75x99fio67hG3HDhkBgYB4XNwg52XFz+YGNWNRbHbR7joI
RhG0m40ctxZKmyJgFiC/NJfM0kJOvPysTi3sZsN7BPCNNaQNoV+q2kYLnywqecwB
+OcN/Sam9mase6Sdfx+jqH/tzVJMJm4SqjG0aqx5626JRXIBD8Q0TYC+6rh8q0TJ
DQh8ymLjvCKrnVXPkrmr/9awNcI4Kh+Y+gRrdrZ5LiFkcFaBmrkMOSqCcE9PDeow
mccOF5VgPgWt3y18bxkNzazDeIFRGwABtMSw9F3mI8dVCMMX0RvLkmiMhS6vi/z2
YIvDwejo7Od5Bk5QmgLhTbD4Xc/TFszcE5tjGg1bRCCg9RK2ufaYvOXc4Ivt1llC
Ehr/QOLyKgezPqf82IdzMUuJP454HjNGp4PkAQZ8TRO6c3srwNfGNAWONgpEoOCw
XKTjiqoay+/pomNmTExkVOWfQIhaiXIjykzIt8n0zhHsc17MPGSsU/NRD5uXeUze
be8dE1MaoojQKA7D04naMPquRA5jAIwrI0MjYfzMfpxEsC19gas4flvBIn7PBMKs
v6F2dlsOynjxopXrsZlMNtMq0mynDVmNGC+6s4K5TfaYnFB0jvkISgcHVI7535DB
GNOyu8N6HsMytdmdZKcFZwBpcZGmidpVTL8fIeD9b0+GQ4LqcwvgCIcJ8NrWkYwB
+RhXRlz3fZ0JTOhoFzpmve3oj49k6shix1D0EA4jgkGtytwtxW6B/QpmbKqV56KC
SWGx+xeWcoUBq+Gcqa5qUkZvb+CQj9TxfktLlUOxlArOITUaF2SdMFH+V3msH1AI
HnYzcP94Cd7M1kucQ7/N8jWtrzWRH/0huAl5Ks85pVqGSRZRtd4XE8+acCApI7ZD
MWeShJ1/8afMk+O0BcsY5JfZe13Uer2bgrPbHYp/VXVYiVQhdnMlDFdSEg26w4rh

//pragma protect end_data_block
//pragma protect digest_block
oBQrxWhMNuAcaQuCgQJhY3olym0=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
z3+/db15jE9E5PwVtKwaGkIoqiS9ISICow9WgDfrn9Vma1ecsDoqdT9PC65YixrC
BMaCTZNQItXZoqF6+pBNyfO57OIKbAMMmI0d2XJNaCqz7432jqMcVzCoI6+w+Wow
WfNKuV6y+q93RCirVq28IVKRxzvKY5AZx8oiUjPVst2HZsNJ7XyG1A==
//pragma protect end_key_block
//pragma protect digest_block
EWnSu1dSa1lEF+eU4HZGFFMJHNE=
//pragma protect end_digest_block
//pragma protect data_block
USep8rzWXgvM8eXzmliTUkmS4BRD5VXG5HSzkTgL/7oWe7eqxx8eSVmLsUif6mI+
lpKwK88ZrKUBrzeJ8WWDAKyoCoiT3B3FKZWmuTzm4nbeybFoEtnSKvRJ0gaYj+UU
FP08fsMh8s6b39bFypo2xNJSzd44jFLZD1bslWZF2JwHtqAqwGqeEgC1lz4cd9Om
ZP9hxji4N10QncIx4glts4xUuN7yrqXRKmJPNa64HdNa+XPSUPkzEGFh0xvOc8/V
OuqVfDMqzX3U/RFb9I6wmh/qLHRlTAJKCtgFOTXQfKFqMZa7i5j5iPkkQ4jGu33v
NMux3VY4QrIAKoa7OITEeu5kGpaS+znKnpw4DTmY8sjYkFHp0/kRcN/HaLFbk2XW
xv7B+KsvdzZO646XVwiP+KDSN1MtVxNJVYNaw0sIypv/WYGbe5So+6xZ84c0zp4Y
NLpdUXZe48HD3VAMkTo9CRVEhPj5iZP8nGKMHbidEfFvSWYsrBHg66yskTiOKmcv
RapLD5SCHTiOWGsEuQwTCMYV7BR6GTaT1ML8s7I11IizceLcUuVrfnox/cAED4IZ
NNzYlef6+oY6RzfTI6iO6A90T1vswr/HIrty8sS9YINksMGuP1Zaed/stDHPMKCc
LWtw3ZUcpQTwopWHndnN41BRGvgLLWi1UX+eEEkaxABV0iStVtoBaMHSJ3d0Neol
FPzyieQ5ctLy9cucUQkiRzzhKDZty+fHtIWnWyD98dbTWVcZOiGjV+SEwv2nOA6i
WPzX0FLhECypl/A3f2OBZEx4po6kbf56BpfBLeKz3XwZiXUpGu0GSoYih2XgZf0m
4KGCYrFRKSaseBA1MiPc4cWXzK6InYoYe6fQTXtTycex47GQ2oVgZBUinulztjRL
ghy+U12OO2868w7Nq6HT5K2xZtd3ZQZfg6BobcjKPV+Lf2ucA3GzgTAAyz4yExU/
82zOOwUBlXixkeuvlUx+rXaZKCsmDktdrnZXmYcJ/W9s9l14kCM1QnG8Dy13QT89
CeHDyo5MVMT5hPbvwU4xAzS9Do/3NYY31SujIwXlTmBOR+0NC8J5ODNhAvNbXYzX
2OrA7eLW/s7fMotv5yiJFY+UhnCepuT6SUrb2nHF1w1wEYbjGkU8YaL4jK2ki9oP
PVb9UT7Pq2sz9LVbJO8lnV84tG5K984fDYhucVNlsK+aOjzpEb9iZQGXe1DbStW0
huInFUM8BojcvUKoAGKp5xH7kKVzBna5cw+6MpPC5I4pG6trkc9mPpYaBdGPGKko
Pz6mHLTrYC6A7+j+5M/7UTdcbVGr1Ii0VEG2JbMWP1Vc2S2hSGmLA9w0t3Vv923K
F4dS5aCZtichwt4YTEcvks12a8DJUD4uRTcN9yembk7xFv/HnygEYmz375U2uSt0
tMAs7bW3zKhjBnvIIejzSmPmlA6bpwqWLXikWpbASw1NeGK2tVXnHlMTpzYP+SCR
0+8Ppy4OOs6QEPowSt/8NGRMOSSE2dJwGjfHc5SKw5OR8pLnq2PH6fjTWxChAIUB
vcf9ZM17LfLHy0R4qHasRJ4/HYrHnMa8Mby9vcpKkzVOIzEz3G3LALhD9CImV5/T
0ZB9xlVYsPQ0MNMIc/2mWDl6qxutwqlZ9By2gDpb3VYEz8LBHT1uGSrYMWz8JGaT
9IE7Zmn3VOjJmMLH9hk8ug07XxW0CXxGEPqHJLdC/MRmpH6UFxeFTZZysuT8z1h2
AuJpOFGdthkZPMH6tiOwUWWGatL5in8dgaoRga1S917V+rPZEazxTLOEOgk6GfGd
Nbes8hXXvw4bMHvcCmfAZIeD1/Hz+0N0s2S/ub2GXqPRlh9PuI9nKYL0Ora/G1z+
R7IYyEDI97LviVy6VdKom4fqzq4mov3J8W/eMAV38A3l3Y+Nmd2cHlxe6Ng2XpNf
Qt0+Pl9GhGTN4A4ih70/n+lU7VmSu+FxQ5m0Q1J6Iy1AuR1dz2BNLFJdlCwR3w8z
zVsXdHg5qqksOwAJx7N9SDtsbxYllMtXae5KrPHZcqEbGUa8RdSPBrV1Lla/NCVA
H1RF+BTVfQ3kshjmVXlqyGF7nb3mRK7ZCqD8oDoyBv0AYj48djjQg7h+QjPXf7kO
pgJtjApHop+PlFH5NCVQ1hvgpYqZg1lWFpWkJrC0gBTJuDNAcbR3r5vNpQjA1Ww0
ERL6qb+P7l0dg6JwuPr1NCNGhWiMSVvnC+1cIHAMG9DyFkdJU+U+VQhCmkHDhMjj
EeE9yVSnbrafns/arvf9lpfdsBpJIRUjnaP6vRVbw1sTxPWojzNVPvd12fks5W/Y
hpBZ/xbeDEZYvCvoocjQECuKP1M3ft6GJx+c0PMI9fYh5FJa/YH3xOgUXLW4MnCB
aYoSWkBsQNDwohTcZT6HCjIAjmbjsQm7S0bzCheZHhX96+mBzeAnlrBxgRqy5hgc
0PTihsEuX1vKaidFzVHukEzlmDcOequWtDvOSWJljjAYuh148IF8+cOA9lgQG9bk
sUFlwMdxv+D/efSbm95T6QNDgsGDZc0HV2d5KYBqwHEbB24a4HEyaSK4O2lXBWwi
g6tfGUJaHB689OpxFjnTClVo5la/eFPn9hXMBX/7NrYCQ1CJA8Eccx7s7vn0uNfY
UB2JrlOsxPn6v1MyBcirmujM0HYD8F/dqvYtseP+LGI9R2yJdiC18C+he1nV4HXO
fAXlJiA2eYCGb+OWNcXjMQCWJbc9fQ6bVOQVP7d0g20s+HZXrXwtSO8rJjJeSAXe
msITOEgz0yvE0AuPyiblYaT+kAtDULpnnntpuV9Q22JHrd6bNX/hEITShhiQvS+W
rIkc5HBq3gp6Lt9imYsh9DWCU+1j76c+Bu786nltl6en6U8LJcHvVseF5/xkz8r4
joVYLS2gfRiH38JPffdSsrqeukaHbyFEYJtd4TIXoiQdp10CF6LGlBlhzxkkvgFw
JrrsEOurRd2jwU3pAeBb6rtxPk2+XxGH0bt2Vvb8MUqmUFBoPSBO+ooauJCpzZQn
OdQ21aMxYz1gz5LG90zDyk0jdbCqXYA/wyiXXHpi/6ndX7Rci9/Ck75LMa6bpz/Y
/qKZwR6GXsG6f8flRK6XPTzjimI2DzmBOEL6H3uGHuC5Az9N0V4Kpn7dbH6vBCcm
7TtEpt/INHyvSUPo50X4dGV3m4ESPrPLHkfCsg1rAcKbGf3ejK8Qd7meQUOiQjj5
0u/iPBgMOGd/T8oH/8CjLrPHD8yA9hchVVfE7XTX0ZH9J2ZYWz2WQHog/AmNe3sP
jO8cfGwga1Wt3k7utA/hvIq+VAiqlrkODqjALqmOlu7Tdiw6Ug9gqaeV6NgZsHBi
/OPhrFruyoOC5YUDBijsivumIl7iAeD4slknzsQiybyuWN+C4Pv3G70eT0Hm7Gq8
GrKFeWYJ5oW1fuQpPsPw4ldp79TSSs8p0F30fCPakr7pNWrBONJ9XKqsCnbQSm9e
kFD2iDeLeutuXfReq2yTHDi0i8V2PBW5GDaV1/XPj6bplemQs9NEBKX4DUQS+JR+
WGnEE2SxTjeosYbyr3nS3dQ4yznOY1YfNtPDQEmrjSQfEYuXWGVv1V76ExNzXQWH
4feSutW9D7U1cBxXYD9cwwrA4RRFSr1kQtD6as2pNieZnbA1sn+/eUCqH9lLcOxw
R4cj9iFwWj755DURAOUssQlqVzn+7+cRfScoiYdU/Q3IQ137IjiMo71nomSiUj7b
Wzd9iQQypBGnkCwlE25C5Rvtpf8Iltoahah371y5CDCN3XGnPWZnZb1OF8H2MiE5
zViMb3caOSqfz52PNW1SUqTIMS2BXW/ZVu/rmJngs/r9b+YKxc0PqzVuG2t+1pyO
czCF9tFeBlPWU0pyZKDI5ug3BPiZK0SBnovimv6x5hKAW2ssQttkXzshh0pODh5R
izmkakaf13M9F0mLH/w+5AsGkTvDeFE3z52QdMGaiDGlFIU4DoHvYwQZnPcvOE6q
NSJs6XM20LzGRWLtVnPJhhVAbljSvnwWRB4e56Me6m2Oppa2AqinFwLmkaIfNLEC
7k/854Uh0Ngn8/fx+9vt2TxgGKJJsJhhsM5vm3ROC5ke6qENTGcdr79dha7PYJlP
WYzn3WQrOJTb/P4zm79xeh6dsph6/3ihBqIGv0G9EFIlOqBo3T1U7zV1YOyvC8eO
XguXR+eX85rrtJBjvP76KyHFFigdDccTMTgiC71scswhKvUwt+n3BDDOxC69sylZ
+hj/tVr91mv9Hm72yfGI+q5rGHLU3YAx9+cOP8ewtebymFRgobuF0mY511ahU7k3
KLxvXIuWJHqmmcxAeB5EtdAPlIeKlJwUmNmEGo+jFiuR50rucSLCdtStfkS8HE3N
dqcrBClZs5J8JHaa7xHuyIEd+J0/pBuBcGFuVRSLIPnKNlbPXDSI1Z8uPA7LSbGT
vbqzDxciMt1s9zqpPqRcmFjsWewsB1g4rR8W/IDp8eq/rP9RjFF9LSwM6CS4UhBB
pvSSUG0yVCuhJSSSoIO32HJcn+OjubkT1uKY7ArkNjJcePjNukx9GFtK5OFBmFnu
2SVFU7RL07g3/hurXXK/rMPEPPcXU0qldjs108w3XxsbYygIw2UBKTSWt1EgxSrF
373/f0sHia7k6MmEaZBY5JZftSLBonmkSoX29icwwzHmeC6g6qXw87qlfpPiD++w
Bg0/z99x9geMEwe4gIJIgd+e6mF/RSx4Vjj7k36XrnkqYpae0Nj1W/vcZM0Kdmj+
yLxlr3VOLFeWDRmrqFpV8kGhEOZl7Mu7YqwhYavNQbBxp6A2xZ7xi2oAhm4VhHTR
NCwe/Pp4GnKy0aQmBqXWLzTn2rgFKGm9nyePy/g5j8L8A76BmXRkGrtocS4ksYEL
61JSTzNqGA4ufK2aFEEBLWmTE20vHTGeC6hhesTlspYBjn3pnfp+Wje3LUkeiMJ3
OmiEmQD4D1S1W1HQ2awar4d6rRC96fY+Ff+pvlQSwSOD6OARf6j8rnuOmKFiR6mU
BQsY6lUjt/q2mQvROa9Yjj1ANyQ1Xq70OLqzJIHAIa9Z3Xv4JGO5wWY2h9mRtb1f
SD9592XrJ61RrEBuZdSnDim2yYThsS3YIiwpjZ/WpfUyO8wwL0Pl+W8ZP7/8d1A1
BYaTqJLLZ9TVCxEMWBdAoINjDQnvPuIjhRqkuF+IkEzaCEcskkYxBwQigN6wR4+R
IW5yUNPT32J2izCxtFlbYd/wia/Jn/jgLRinFmIo6adNjxdgCRv+J6MVnQz/G5G9
qlGrZAu9mK60JzKdw7A06i7rdREBUz3eX2kpUBbqj6LKxcsmMJ2mmA++QOQbgm99
RSGfdUPl/EemTIiVFLQsJ5m4G1kmIMYjUqGAclcehLs51uOBZb4ClZEDJNX6hwsz
3a3+DairNlF/BqCIlskYCCwkEdOmxdCbltmPFOpbl362HTthZwN/HF9ztKZuSmsg
jlDNxFjXE27qW3GIwH1BPZ8jOw75wew4fnasIz089CQx71EFBsEYnFmrqMyd7xe8
yaZwlCPJS7NJgdp4IbVol0dye+CWiW+jhVwhYw0b3xkhEF04nTVcVKI2PjVCGcUS
WMnzbET8hwJuwoACE+gD8BbdHiV3iN505akia3RlBBoeVuRfjxD1ACcJgui9t5bx
ZuJvb8ShaRPMamGRqpysIY33VplrErUxraFpsaLbkS/GGX43mQ4U27sqneCkGP+I
e8qcf2ZbzS1hIpgDNCPUzCdBuT65z5pj0EHs9990ozvgfSDExjTTm1/X+jKXg4SS
FxmBfAu1Ud36Qonk6ha3JXuxZUn9+2kI0oGNaI94DcwS6uDMJCzMwqxZDEafkaus
HSh17XDWKPwXvqm/EhG8j8x1RZ4Mg24adDyQnxC7xWnHfWDs5VVeHaXC2SaByD52
LlkR8FZnYTa3D8lHhmfYFftTynHPemgHFmNUKsL4do3Fv+8ANKCs55g4xglJvRfy
EFE1gFlgjEJDGjSwm8yKCyOLrpCnTeZBLgDTwS2tJonNXEc+6xTA5bwfiejGEN4k
Jeqy+rQ762ost2sKxmpTNRLKexqZ9DM1cyphtiWErQcwMCPmIdkl88oovNExzhON
8rvrBIY0v+IB6E8Co8A1BUMEAU+7HJZaIaoaPDW/KFZEMInjIA3DDvGx+S3/JuFh
nVNixaF69Qe5PxccYDlEUU06dyiyG9ApWI6jJGVIVmZ/dfH8GV8bhnvnInll4woY
mkNDN87d492nXsV7/OOq8t4Ff7/AT4+0McMbrHK0kn0sy1aoOEGi5POWrKYGvJoB
rxd46oVmePqvJreuRwHGT6dT6Suh+WOgdlmfiwjoN7YgNJVQAENqutQo1RU8tMCo
bwRGVoI4Eu/U8vjXwMKSaGirfnn9eytYgBTsv4Jpy5SYpmJU0E5E2UItH/hyEfLF
wMT7GijuF39ZgavvbzbKQRXt6wjjZjKeUOrI/cgA6905l+XNKB+8hhtGnMx0hksp
Amq/8D80/1YDMCBfsUDNrmSQwOFk1mV5yrx/ZzzfQ7vhILEFPz8s7x2C4cE+rwMm
1fqTe/qZ7XZhirXAHCfAFGQnr/nD100t5wCr6HXRTr9t3D9C2eb2+7/a30xau0WC
v0GMgDH4GBSvjql0DWkz/15amXwRUiMjowbQ8kmXmw54B9bNu/2nB4jP925KaSx2
ERPbAOsrowtb8BxeaVyxTCPM+blohvhcfGmOcJYDRtUFDeZlMwNGX0NH1VzN1Ybn
5RLFvKpGi0/dmsAOZuhzuT/Njid0jkS2JgNBVNk9wDexXTZcmZpEPdFURvx113WT
dMUx0IH9YXFUl5ZETyWDIFyFSgwG3q54ZGMcRBAgESHCl75KDcePqLsWCi15xm1o
ioryaBwI12CQQuxJG4lRCvcZXTygQ9crMGRIUOwBOoyy3X61CUOIPu6zbPNW/X5l
qV02paZwAnrEqm74snH+0SOqg+cmnVcnW3F8Y8dDQ2RjvE058sicoQtaOJS2lYej
TmZFmInv8Bxmy1MOjMYmO/uaHGEquu3izDoYPglOiq6IK03R8/xq8yIqMOgWgJa1
JNqKm2oBAz8HKIDe5MOpbsskvMlhiUnS2mFttjfq+DB/i74b8DKSltgB5o09eRsE
sPz/pxHoTXwqByr+aQ3+J5tA3yNqHIFTxpq5Awr+psSmzOKOJlPMGteYpj0qzBc9
CIpvEdkaXKkBeQ/ZKMjrlt2/Mu4hj0+oWNk03iE9Wq4XdxoLqo8NZWuyMhPD376b
yp6DZKtkL5fNIZiML1SxFa6X+R8p0ZSDgrVD4IMjPXI7SmoFLt/VAMOOq1eQTpv9
Qp7azee7tocHm2dBrtxq6FU5aTHSlK/uPycehBbDFHZLnDdi9ea0ZVGfWIcngfLb
5bdN3ACm7JS7/q5du9Q8gkBSwRNgA6Ipr+1iOsyWWrMJaWLZzfXJ3qzNQNfB3hVL
/m5YphugudgfepFLCqwT/JU/mUvSkY8UMv7ZClJ4sl2jnV+4SRIi1+BXPhf3WVIS
qosEsoGmiSCJa3cJxfdl/jL/ZXU3abAo8ddt3s3KFv2Am97yqGFJLtq9UdBf0ovH
cGyQPsPso75LmAy2j0J1JtfrRjz/J6JFVX714bxxJq6FNFUmvCATeBrduaP1szA7
ti0LYDXBMmJ4O0r4rCQLx/BmCDGC/bw+TFb4aKlQd2x9EXzKW0A6jHFbkbexemCx
y42IzA1jYXEBEJZSVg2adbl+xYZVAQ14i0PMr5ghVUeOHuJtGHmXvdNUSgdkOIxO
kd5OmQODBKylt1Ti7xJuCVEx5875YWXPOOqQQbRT0c2NKiFjGZ/kZ3/4p8tLJhuH
kT2qWvc+Q4DQ3EkshOoiP8zp4pRObt+uVXlq0AXkEf7B7B+4Wi51JD2v6tpXr0+c
fucipSIqzi/L/vF1uW/+pneRMChGwKSs2HyRcifCERh/KkgKFK4QRU5Xid4HukBN
W4FXbm2BopwoYza8tdwR6pC7Gl9YEhG0u5cAVtSt+Pmy7TFXBa4bP3c/UxZ1f3kC
fbyTBKOJ9v6uMSTxNZk5IIShEBg++WiSWUfl1bqrBgDfiv/vR4xYOeTCil/ACUR0
ACQ+aZOC7VBm7Vfck/Wzu9ZDerN5swom4A/b85Ih/UYY0UfA+PG3zNwM4mLhUrt0
NFT+j2RCx4axM4+fl7JF/QffaJalKNBWtQ2/Uuwu1CMTa1fHa7oxSt9Omsk1Ynmf
ssVkBoVx9OKI0T7j9gp89ToxtL8CI0obmRVgRgFjwW0u0qtEYL+963PYNhzsurCb
cnj9SnfYagWlWAwEy5TicReJY3B11FDvvT1v/Y+hKn1QbtmVrMM24znnqKOHLIAo
YwnNmnQQDJXXMi7Y4n7sJSOtRFCP5tadZvoYciaPsN5SEZ5AVIKli1ncV+q8L1EQ
1A+rxkKo2SSoaAaR4yEG2X4xfamamnG/jKU+37PCGg13bES/eE9bVN+gGgwmRCWB
3xvPlgy+HfWtL3MDfx7HcCDKEUHH79c7PWUbfclJ2CwzjYi1LWkpG0P1kz/KcT7f
DEDoFecnBnZW/2ioAbuj+w1l36GJMGM8daEdAu4H/Sommbk2tP7MFe4FSoNUvh8l
zsDZx9vRSOK7QNafKLvjsfXFvkrtFhv+QoAAP865KtZwsHKGAqp4xBftyIbMjbXd
PMq72oIJza0pnJQUTe4KLB1Gz1Pb3CG0XdkRbpjrjRjh1zgsdmlgI9lZWJbmZ/NL
IvxIDrZq3j/SESuYTYRp0CYNZVMjJQLq+EZBfIOaomhIEipR4E4nih70jdRh84t7
IaN1IRNWjkviePp/kb6qp9RAWIq9dSNxU6cLHr8s9io1EVIo87iI3IFY2A6dL05Z
kBO638yqml8OQoQCJQex+KYSsfnopenDJRrCeM8jB3pbPs0+cqmtV7wf/jJBFTdS
quYFDZLhS6THRoLdMg6zfUxcgKWLijSj+GrkTn8yIYvSqjdVrGzBlfoBgGBBHLrh
sSY07AnS3SxHtEdbVTzdr1PcnvmXyFy6bo1/TAoy08i3vshj+E/8LJ9gECcVxYsN
2DAumfSkcXNYK3FvXommxiw7uubsNI20S6RXccoosZCdS4yaGyQQLlNb5nlr15vP
X0k5e8XHLbzJQxrNtfcg67wbIs5Vz3+7rltOnJs+r8UKnZ4L8GMLJuWbgqW6YBDv
BWxyfYjJ65aa+dXUVKLCbC7KywPlNTe/ndk0T9mNZD3o1raqbf5AVKeOhCEHR4m0
H31BOAf/d1FxlKOnnkoRRHw27NDj7nGd61PihgW4KIbzot0vwzCLUpgJKqCx04Tz
QBQkC3Ubx/dwZZhKPXGMnNUDRCNbzpL6wd0uR69WCTnMhhtDsyw5D6RJrmIe3aAW
4MUs1ESgGdzqlK5kgEf/0dAY1dkBP0+cD4aXW04evC63cq31XXWJu3HVzOXwQoYU
S0JoYOQRUcvP00GesgPNV/5PNuNfnQpBCN+zPNV2X3IJ18qVqjLIh34N/emvusxF
vsjSQrFG2Qs55SFq+ah410yfjdhA3RbpXiiB6NUIu5iP947Qwf6+sYVr7I1CtCJ1
1R3ilMJhUp4ms55eVC59iK5x2qQ7sY2TLOstqR/+nqu+TpZ6AsUMBUJjvfzwjMpr
W8sbmP46FGS01Wd/aAMuqGGAuw80lY45L2L6vrA00FEhQoI9vJ2j9oasxB6BLBT0
ajZpQdsOERbegEK8uNQQkKDMqIIEwvbLYTCVl+QLcGAOnuUZSEuR5tqW3EPrlE3R
oP+2taX7hZ6Gb9FlOrXRssViOrW65oWMa602GN/HqG4Z1a4gaFqxzFAIDv2w+LTk
xq+N4G2AsCEMq+t8T4MU5ab7fWO7o5JoqUSfvNneoqVK4+nJbEj4OT3XHJCFwA3M
DTtn6c0bhRLmZD0dhh+9CtXWk8Hiv+TBaE1kNyjY2BWzlbbtaiQXIv2KqZleUhPA
Y3UKMsC/dJOKR+DaML/fvqo4PGCT4ZSKCa8jFsGpoIJefDUQVIrEQ3XN4ezfo6OJ
9sNt+WaUhuHkc9qINeeoYWVvqeJLdKauq0LA2F20wqRg8pyD69vINmHIAvR33HVK
IQVEc+iPxAlr4XcxPXl4zotPUGK3d6AdrXlq5+rDPFIwX43nXBUcL2+QF2pwv6hY
GZhvvaQFGMb78dEFYy1hDc/MR7/jgy1gh8xwVdsqHmhYLHc1+P3bhajCRQJ8bFor
2j8rGNTZpwArVZhLM4ivA3byfi24TVQhzQedcrIxWRq7Hr6CtbhS3mbNOLfdL1AG
7Btzp9nmzzdNbkC46XOmm2K/mA1or9bJB4Vo6Svn+3uRMk51VbkvW3IbRT4TYepQ
ksyrbeegAuDgMg6FNNj/NFcnIpdfLp721yXp1lx+HoBiqx9DTo9pQPFpYuRjxjKe
On0GjSQImv+SkHsyX5Sr9vfLBnk6+POv5zqjifX4C9Wl5s3sCW0A3az1spm+YdX1
5SwjW01pJFf8Dh+iKipByqqzTArM8u3U4NqzPmwVP35Nox8idv8WVBWPlC8o22Ji
pDjs/+G+QlaBqKFgWTJ8HyxPtVLmkfMPzS8CWDMQV3NpLuFm/O8C701J/B2ZvNsw
Emufa3QbmyMJ9zjdlyNWrFWcphL+6PIa6U/PY00ZgobrUX8bT/v0C35QgvU6ha4T
tAag4zylm1jeMWbEIPvL3RkWRTL8PGDgju9Sjbi/5hfLxhlybVq8cPhYE5Kpmhcw
XYHAowMpXQ1ygmonIMY7VELucu46qw/A64jnxwReuEJDu1YN+JndcXhMsLudhM7f
bjQ52J5Ad5NnJpUmvJk5gbATdpqVn5Ypjp1ccdk9839KYSxC5ddy/I6LMU4eFLw6
b2SOzn6NaljOPZLVH6MR76N36Dh+sUZuU991IAyIOnQgYPA5f6OQjG7+GIXzMDRd
zuXQTRDfHV4LCSBUQaxNmunkZKlQSvfhyxtisMTGFqYk8JXK2kER+n7oWGfd3rjl
DOwxlnZA/sVdZZqHgl1Cj5Dl1gFSDWm6ydWouKo7dfPMeKnhS50GbawvPcPsvfHM
1illz1AAjfupYMV50hZBJyEFf2MYlqdfaNOta6o/1ADwybOmmK8ZJiE/busYGzMG
anI5rkDtzPgjcnkpPd7yOcu7qwLs3fvuMvaLrWrPsaiVbpQlKjH0ZMGMrOkW/R+K
qSDIbDcmCiDOG25YAcn8v4OrPoVY+LysCnxtivNjyMu1ZHYTOx1uQMJUxQKIhN3n
yOZjwT6TMKvc1Sd8w0DJRAsRhNy/dDQDd8fruU8QJV736aQe554qgavsL9n/eh+3
ErIph7CBHFDIRdI+LWG+hA+Z9Q7yScxZHfuOxFrRsnRYxgqAUU32Rx0wth+gwjK7
gRrvMOfSQJvm/0wEXeagZsTFxIFh2mMxHz1qbHn7vfjKpiq0uAB8aUEK8A9fPlwJ
uBC3oz0XT9tO5wYAq4cGA0nNlJWdI3hvSkiFxMvZJORzH3mt4nPPSL3LPsZYh8Oy
fU2Wlf/f1apYRdfmBOTF6vqjIZnN4E48CBdSp3DBismibdzwKkwGoDXxGQ+o6YhL
RKtZhCmlXIRKmQJLmFXvYEGB09Ne3AnrOS0bxm3Ezbwf0OjNFRd4XuLjWngiqa1o
mRf3ykEGLoO6mKl5QuNvoi9Y5n0mdN/uN/IkyMBou6VxHkFkNHF2XjjD/jzms2+z
oqBqMUfGFq2GIvJgzx/NuyYQr3Wc+rwI7Lq00fb36pa42ZP5UVQlBJTrTvUMvnVa
iu0G2AcQaJKCidr6jlU8h9nTNMBDwUBfUzibpm0TCxm7TFLX8TgqfYIpbCpgt+vI
2uLExbHxFFy7OG25BcBOtm1O3T/sAAS576d6V7Ec5GytMb0wPhWi2eWZDL+4/oZP
WD3sQtsu4bSW8RaaKcbahjzWsSI3zjXHFD6FLIKzW5E6TB//O2RkKxRfbu0qG8Xu
BEAYYIlsFmrScV3LgVSEl0yNaMUn2QdTaBtSS0rpiLp2p96m44uu15QPxjFayE6S
xM8Lqgiv5LkT2i5XSkP8h94OEpqmSe5C6PfFqvCjSUJpOsBpLkPEOAi3xdtGL5v1
JlXrtNc9LI1XDKT2aeH9WXGtdlvr8Hh2fS6UTYTCIzuCJbMeNT06OdUBOjOyVJKD
x3Dse96Tz+4tChYa1S4jCzAMWBDJ/0SD3VAHzjxRQH5Ul5TPOmcuqD/ffi6tzbJ8
YxfIPl/FT540zjRiewgEI/5a7dxVDVNxne4UxkBOdDcCz0WzusN7dav6MNVnFbP1
101kcZY4rZ806xawfyTIyWA8C72V73ut056hlsPX1yX6cbW4qeLgw5R23nz9wnat
RHZ1hzTIwqgNsp2p9ZYQazXyMfvrQUJIgTe+mlqN4d+EHc6apkYwnr6Pun/b2AWT
GqsvzoFqeXm7EWtxiur4x5RjOspYLiTH3oBBwhj/3o1MuAx+YTFNFetiX9EohcoG
6eK5xZLFML2EcuN+Krylh1bpyrmzEvBMB7kUGmZSidEuKIMmwYm4KePR58VbVg2E
HZw/Y1IQE4pG4Da7XKs38bPZZDh5aqIsqiNENKcutRpAQ0wyLRd9N5XTCfv+V4nD
GHCgPufI4D87xDv/sXjKFyxyxM5wQ1TbJhRD/hPhdprdQpHT8/Ez1JPLdiy7AHjO
/1Yo+IEniMjtqFCNAhrp7q4V/9hus+fuMuMrSxJBk34t4PluxQa+xCNg6RSQJ4t4
805eLoZTpMj3Z+fIC2YhKX8ZQUUiIivZW7FYtw2ZlQv2IIC8sTPTdx0JAHyj6YGm
PcVWnmyPyeOY+i0V8iM4kxJE1RsiVVFwGNWJSEbKSAjJflXCRj5pI/NJODYzNQ/w
mtZaY+pl2oVmtxXd8MPcjKmF+o6QipJTtkIxASbOeuOxsw58OWKDsMl+YYMZsQw7
IvLHKAoHYJ23N0q+BZq4D3jY/8c658F0J3wk+jkwtVVtbbcxj3qXdcb/sxejFQsT
TnHOs276wfWy/p0DsFJhp2mt/lmymXEGUznHVMXtDdw6+Gzfpbd7bCxhdK8QNa40
x2vrTgWRE2v5i1Gbt7ivP3offZVT7s2ztMYufUzRUQq8SM6RWzQs6wzN2vGSblcf
mOULCZs8toKf1cXBnlwtIxHeJqitcXWnmhYiU/rfIt7TDjjQ2hVBrELli8xE+/BA
ox2OSYF0L4cxVkC6xLnjQ6a/ISJFNCxuv+3wrRxmzrjMoDll7Jq8TdK+owhFRjNI
V9SarhIN7kfY2rKbDrkLdfLt/fgDlwQ80+eTm+pucbMcXA7OAbPd8x57l8k4xV4i
zkUupJUlxAvPPmilNXuY+ymtOhjWEGMv6QU2cC4IYIfERr/xLboULvEFml8qA5MZ
Q0gj1nMT3PyhlSr59tWItGAV7ECZOUAaS24OHS5PS32a3GrbkFyyA1VPdGyWM3te
9vlM7PiXqOSTPSqP9edxAqugDfqS2wS1YnWOiLZfd0l4CR6XygsGscNPgNPo/JUo
KcxCEK8Y+XXw1Lqb3ZI1pzGkLFZY2lwBl6yY4iNACgD7eXZtuyhQnex6YKhm0lzQ
QQewAuKyFdNEVNO45zCyrt5Z078K6Xe5no02xbJSihxU0ktZNfEv/j0geI/SrBHn
e3N0U5dXWBNPD+8nLvg33pdimJ2JZMkD1Z+k2IAV//B2sqztdG2qRRHIi54bxmEl
n6O2AifeRuf/vCINcskOvhaVb9W+SPep+FCnz8lsWTuGevpHZ7vHCQKd5joFNuyS
5gROZPX3sIYD1Ow5znC7BZcUGiWNQW6ep7YsjhwPxldvkcWx2MU/VEn68PLLwjc9
pN1EDrwFgkLYVbqlBrnW18PhPiyMK3MCZItlt/GBoAynyRVbb6adq8GNCt6mSNUa
mFD+sWFnQ4n380FLIamEgq1Uc73MG7Q75Ez6BLXawLJLsK6RagtO2AdW9/kHqbBH
OwlV6/ThmhQDFTZ5JQJmu6UDuOXGJf4sxKXnI/QWH7b1YGR5xRvO3X5MEyWu26rU
JNgZzbBnWbsKsjVPyGX5uKuwzbPMi17r9ScDuGPsVe9V4AkBn5PABwYxu9iaYJNS
pjq1CZXI9WYzbDuzFCldnsz8FNXoBSGuA5W7u5HeOewO1RXfMApMjuBoejHibxvF
mbkAZOMU6a7R4qp9nxZyT6cxVfmDd18WvC7lmVnw48HL6NKOz14oINJHR/lVMdco
ZD4u4i81g84RF6MPyTNXMv58sarW/oeqQltkANXerCL6p5xG3zD0K+JeO1w0/mNP
KcuyIcAQzd2n1dwkbznsP+eyPWxYvv3pbRNX436ijMAsOiLUcd5dzQwYhwgALXzb
oNV+HcGUNwbNDynlZM7xWS0BrmyQ3/lzBct5kAEPSD9+ZLjNFB+Hmh9KMacjnsMP
0CQ1pjZoeqJ7ONVHRNe7gwlR4bmaVV+2qWfwND2JzdGQvJ2wKPg0srsF/YsGA5al
5jS2uaU5Tl99kurJXmXX6CmQb6XaQkaROwiAl9uXEdhxqLLMVW+vXl8xQnlXPc03
pOM1eGEHLpEH3emi3VFRsb6Hc/l7FYH13qcF31pkUZSCR+Di4gojFa9ubGY7HcvC
jh+d9QjHiWjtiRC8M0FVyRz7vLPeh6Ej11XOg8TE3uoQOXOjeXUgzL5FP1UuMkn8
SDUHOWvlxp0LE7iRa3rzAy7AMBLKSJsnFOy3ywAM/+mitSnx30xva9eaFafWAwei
Sl9dJJmRrABU/OHB1J0h9lgKeIbcIZM2piHNSvF6eISgC0CdXg3ipvtafFjvktbA
zb+H0OrDz9uGZ2cCpQ79J2I2aDY8a0lDR4v7qaC1bCNzTgVI4wLrwZaU18+8QNEU
0llh4EVSP2T0d9tnnv1h/Yzajrwd1nC5f5B4JnrPxNoR5HiPiYsUaVVmCizoIJgp
LZGlPSLpzOB65WYZUE6wQciyeCzGI4BLuKIvS2Rh9yzjNsET6EHUeIEzbvv9uKLe
UVa4Q6uGOgaVDQxzA1StWh/YCCMI7nW3AXaqGZRUPgtDio07rNYfjG6jaYLAD2gm
jxJZljHrFU1faoPZWAOhhabZEfGUZvipaR4UvilJSn2UewBvizKRZAbLmv5386vl
DOQHrG64Awa/DdhUaKJH8cg5/NFgezfLRzRvUecge4IKaz6uTrRqiPDdOG73x9v9
+mH90mQSGMyaqgCNcXAix95J7hOnG9XY4ITZYg5nd4C5xAQEBxu5LxQn/67/EAdx
kGKsc20AwviV8pZLYSOyc+RlXuBbTRNH0FeS1kdEjKLb/IcWgB+DOhTTiMJ4pXew
XcP+5UEq8XbFktM0c9hfq+5Dhp5KJ5tbg6VX8eqKEKZNABrT++9A4g5TKps8+iV5
pEUPcv44Fjyx9uNUSojl6IVGqcPY+EO7L5pRUaW+QUHmcw0KRPlI97kgi9XGvrDo
VhVN2gBwLuXIVSSuogxkno2Xn3do3tD9kI52CqzLXQjqQmfYQG4v9gkrZ1KmVmpX
FUe/L9m1vVklBPg33ZdnGxoEjJJxd6ybtKz675/FZenqY9r0LdTUqJMbEa+NYsX2
KSdYmQLTtY+4jgDN1xDYKnTpwCk/H6eHcMXxU7OKaPUSBt8XFV/tx3u+hFhbApQM
dRlAaTeHZ++Dih/PP5Tl1o57xBAO4d/BKhb2CSDZTz9gGev5REWGRb1QAul1X5p8
0e5f/ro0vQr3xqbKes8vjSElUmRxoV4OiYXCCVKfe6HwHUT+B9kOHA8CkaGzjks2
OPvU5QUb076Eg896VdYDkYd+LtZMX7YaSlATmax14LisGvZ2t4hT+Xz3lyah1nN0
37TrHHW0nfCWeo44DI3iGgRVRzNMWIHvQr3VW6++XZtrPsiT3ZigggU1/dUPPmBL
r6FSO/KZRP10n8QXS7/B5CN45W5q0yQ4T3OXQTPSvs6Gr8+aca43j0BjwqJUfP+2
2CPkUp6aHkOGJvV03ZtCTm2rl77ArkHRLL+RQZxKcOyRb1huz3TQM2A/kpk4LbkC
h7hOtGFI9P3/F+F6H3MFXwiSDmD+5kxv7d6HXuaCFT5wPTPCGGTnAQGCi6FAjItg
gnHcjjP3Qp4+ECcoXrqeWMR1zInPnj7Iogqh4cY4lvXBZUxst2nRFEkTEs5FKoeB
KkzhZOcfOxEdySNwqwiXc1Y+Xyrmd9JOIbjBpof5jspdQhrJDFZ3cbdjZm3ba9Pv
CQjrhT2QWQNcNduwtXHb0Sa3/UW8Kw18LaBz/BJukUOvJXo3ZOSylpUqiYX0i33+
R1mUDjbHC9cq6y7wawrGTf+BTjcyHu+Car39Kfy+eAzhO66CyJ7qmA+6qkWinpvU
PY15jueuZPeSUJN/rOooEiSaM/x8ytQZ03ksKudNyx2r/GiM4peuYpHQwr/8HhQT
sVO4TnVajIpdaVpNAgBLfFGGKHhIjqJgSrWvA8oj8Lxi3kDa1S1xLT9RtPntS5RO
z6ZsXCmg36RuL3J4W/RiqBsIeqvh8UVaP52X2JUqghzD4KnG8kEJLRon/h9lmYJP
Gyi5qWyr1cGt7xYVXlVxdZAUbX06cGV8KhAjH4vagA+RSi+T92L9POyp4+QxmM1V
EpEMiR2+YjNxpF2WFJmIan1q2W7NUfjurbsLevuY4AxIXxUH5iG5cxNB6Fay7ja9
1/avr5vMmdzL2Y1uW0uQ75PbLOB5FLFtPIiQG/NFGfzsFjwnoornd3sGL7DWoKg0
ZbaforTwAOakGjJ8I/jBQzakr3XwJS8rpF9vEsnSLyy/O0sV/lpbvp85iOYp+tpq
gnO+JBC9AG/1aIuawjaSAmryfeYZMkxn+jtb5xk8HYUmR7WmHQUYy3zTMNE2lViK
Sn2jMMgxq6iaezdTak9td+E1BeHgUaghL/yAO007PKv4WDO10jhO0eBkwgGyVvxT
v6qGTU8hkF5XC+4SUHthUvv6ue3hQ0TBzc+Y7XBwFO4Lc2BNxsL9o446pX3o48nW
3baUZPdRDXhuTyiTEBE5YEoJ+xEECJ3H612+b0342QAcI0f+y81fMUweG0wa/+H3
kuzFMAQ0dSoijeCKXt1NoVHOcC0ZKRXDpReicaztWixWG5rVXM4pMqHRYHJ4ZMx+
bnmqRQVTrHc2RzYjk4VujvE+UymPo6adr2lToFtHAOtQueLUahup7KREMN2lgbzE
nb2DDNtIHe/ozb6pu87xMZIGcRmREiMqQDogm8f0WYr7FJyc1MtW2mMCcA71wpol
/rCVj95c/qUfBUZGm0IHL5YOFdwtSdh0zHWfw8NWEmebZ6aW0bUTtYTYhbzuoUyM
H2CabhwnnP06eSmZsS5eauuLJuBgktpclfwfBE9xhp8tQFlnq/Eh6W+A004laXwT
ZuoUbnnYWCIM6Ghs6JE8aOxHVc/jgfeYpgDHvco+Jn+XxXGoKeYP+wKghtrlyBEB
LJVahbK3QP0Y/h2BW9nxZkUZgdFdLQfCRvez4mD27fVit9VHkOt5a7iScb4ZnlWr
vTqxCRHsDPJnopGsSDS6MIhxPISlAl0b6m3LBDdjCg9+w1pIJt1K3hJC8paq7PJ9
ilmeIuZ4h3HAIzJX+Wsp0eV7MZrsTm4y5XLJbKb5tP+vj+5CtWBnoJHg5V/RQ0xI
4MtkXNiFWFioO72S1xGgRuGBeJiy6Dhj5PtszKbUsQn01Sxxryq9V+5oZb4farAU
b57DAdKLaGpLLgcdjq//JQNFw1kiKCDoBT9ehE9Y4j2iaDAMPde2Efjjd+pvC7Do
f8UdQ4TS8DM5aaqhgmkSW/CSiRHf1FKhHopsBwC3VBXu4I+NVDR/RI0ZGfNPopd7
44q7+IN/fLDdMrx0m6Tl0ynKuSZNyentF8y96f7SGFfnSf8evKnDb/hGEiI08glT
9HawxKJ5QRzRl1oQfzGzyxnhpkFw5uLHMxT/bB967n6Uism4C4E26b4uhVKwZKd1
NpxlBhDieudI/kloTu7QOmwCxA0ecKCiHmnIt2RA0qaQhuZdLACfbbarHDNUOOJC
Xk2C936fqOWH8xSdmzUclYyVrzJU8PqKha9V6ggGrp1NpWK/QIVoJ0DhSEWKtp9c
bM1THwbXvsvf5zoMsp1cUnddSUFYV01yVat75OvHlEH1g5nqWQ3EfAViWhG6I9dQ
kFvvGrU7KKVEF2ZSnBwqCRI4fkWV8PDJXbLVY+MS0iqJ04Oy1Ccfx4KPWFprwtyY
6Dt9dPcMHDaeF6hvQQmjUIod1JGmjV59fci5NeG/jOe+BcvaLk23OepSQq/WZa1N
4lNpNN8aaHcyMRVKdjpi0yg1MSkfjS5/LS79mBJnMB8QQZRH1L8MaWtnRmFa4Jcb
1/VNkQS4LF/dOelBZdEOqTo5UtTHJ12iFDUXp0/xCpC7617Ocyv4IxrcfD1EVqAE
ZMUMRvHB8SXgCGm5T62tVawwWqycx2jZTPwW+UILdlroqJWlRWO2Dk6nGmiwh32K
NLztZu5cvQY+q5M9Emrlk3u/RDARnAlOgvP/lREsslKk5a66vOG0YjALVTeqNYAq
Al6cm4tbpqay5aLtQ7nlrzT8CtTeQGz7+4Sqdrgarjxlv3CVhV9Id3NUAR9d4w5c
43o+dwBGqFCv+MeUigneGa5FZELwD3rXnh+8t/h+fIUUBW8gfMkL5MVNDqpCUS9n
uxxqzKO73F55gLkkzKSFZeNv+jHu+cY/9+qhF+a7s1Ot3TCOv4MPNADX3k9Ztsz2
0U6vs/jgiqyZ+4Il16soZFM3I2HNLfGjXDoMrxJgiVp+XhJRDpaRTuHCCuNI0hAC
zCTHpP4YBfkKqJuLRnC3AeriFul4it1CIyfgIGBdCS/E9VUL7gYpj+faE3adfEoi
ttj5Iia5TdY5mdrQYMUWcBrS3i1VIiVKS7ymeLSf+mvnnkWDlwG7e1eDqEEc/udq
jU3qG2BrtcTWOl+olCGU6KjsH5R5o59MRQdSe2D6v6ft1BXeFvsgztdVnd1s3F0V
Qe3DmMk7CkIrs5VdfQUO6B8u4aly/sjyqFLi9q2ysp3YJm8V1/pNwc22wQZoOgW2
BmJovM4T3L0OTcJeRdRQpsTpvbpq8KnoPfy5c0wZqXfeyZOjKoyWB+8vW92ST7tN
YO/UJqXwb5KGy4PZHIxCp9VMSk3iHRMCob/aqPAeUXNsxrp6Sp9DSC48eXyfRaXY
fDtOc+4x8+Ew3VuarupoLlC7r/6pQuiF2OY+Ja6Ukme7ztKPDjWSJXZFTZcM2e9o
PWI+afv90QalF/x4ABE8C/QkBhwL0cmVg93lzxTiZgALhjhow6TTDL1YslaPi7Am
9gjkOIbovburvNkKic2toR4tjefyS4li56jckBls18Ko9RbltQ170mt6TlyMxdVa
KmJMXR18obc/Neai7NIJ580H4uM3MVlLoCifeGBs6C3yiPH53+k45r4INSixTcfu
IwsS9b5BCGHn0+2c17AR2/oGc0p8aMh/MFlz4mb7/uw8+37TQiWfQSgdgJ2p/vHi
EAA6Yf6LWkJ/sj3XH2XCdqadkviP+blE0+E0IOi+Qn9TW8GvDYH/uUS+OMcddnJK
b40ezOp3cdLZfkUrClI+XEIgxct6U8gxvbz/Ag/gjB1ky5Rr+5EeSvvL6g8eCoJK
UwlHu9PaZWLmYUG9EukshGpx7fB4gdWn2tAT0+w8azSiyTjDO0OzYkzr4f8TAopc
ijiLxhUfsz06Tg8EgMmsqfSzh/QdCpdgu19ApJy3I1KlBdQeTt2+Dqh7rX22im25
/nBCkFry2Melq1z+v8EbSrXBqKeIOTSxvmtJTkXasvS/YSlxzJBUB2N48zolMnck
EmMNaSAxpfFP6folL1s7P6PgdmR0tgmL9DDhvGe5TdufbO6GV61tjPuUfqMo2Z7Y
0xVObrGkPb7MKN3lEoVOkuWqZy+cjDvhdj6xhsnZTPttRjxrW9/JkkEI+lZVWnda
pLrFTjZnA4rJ8+CdE7pHiZcsVAzMfqBZFG4aYglCV+G3n5EmWsNkAA3q9rhm0LRP
AeKzoOiRDOTWb9GBbnr5t/bhGwtJCCdFqBqOMGXe3NdgLo/uhLbpfaLd/aKHGS4y
bQY4F+LM3POKskVKcX8A/jPZyoiFRl1Ul3Bod0oeN6zaLIqfX1ajc7+j62Kn8YKj
/KdmBb+d8y44VdLDZl7dgZ4cJAU1XZlH9WCCyPJ3m3ugyemi4ZBtXhY25Lgh18EO
GGgm1yjsJsFL7aZQTcT/nXe3wArR5TEIKWnM2K2bJY7/6bFeLEXyvME54q4CVSL/
CBRfMol5SjOn8vgJ0HvZJjam4XNOVi35QalM8qg2QL15brL5SgHROtFrp2gEUwFN
UyK694b076V4labXQA2qY1Sd9WtTITCzJ1b1HK5mZOeTB0w0ZT8+sTy51HnmC6pF
gOUDCGo+Rnh/7d7OXSS+begPewYWkwwOK3zkzWOOQRZWqJTW3wYUXKiegdeGSXbL
Ixlp+ZiH/3JbS6MB6Vwvk540UNvc1mjouVEinQfjOPAgkJDvDt49ZfBhX/0tswfb
mDxiOS1V3yquWr5tK7Kbjpj9zTTyoeTbflPp26Co2CHWBzjF6EqLkC4TICuJHsl0
8g9gDVhs+WpFilltC4o10d1dtor1sHmX0AFdE14SpUdYTlZ55KRCZ0cdM2AigDlt
uWqJqxrah9R1gvQ+Dxbu0sHdARNwO41XppSQpIRwqnLnTr+XplVX6CDrBx5JFbZQ
yFv8Vu0/krqNVeHoIZZTGSzE2o9FTI5Fyi9iKfE8rKYUbc6y4xKkr+URFlsuO0lF
+nC88gOfOe6vVIlYDMvUHtLIzCnZSmde75Y5SkweDBvz//49mNnfR9oVTb96FkNR
4N5TbkNXuUEpnTQBzhsFNQ20U7Wha+S9vVGhpvKTEvNDwBsooZGvTv0gBp6N1sCb
LLDwADRwuP122noYhThVGsWb7AQryBDM3NXLUcvSwGce0RsXuHy2C3GDFKB70WNj
/fO305yuGIedBWDBm4lwxDJPZVm4bLHVVmVu4XZECcjFmbjJrOKAAdJXfhSdkdWx
UCaoE3mhHwZM0JVdh0QWWe4eHPR/pm2Cw+suaPMca3O35qSjgBlHXqHGhstBn4of
yXlq+smkbH47nT/e685pW4K8bRXw1PhXuZ/nUoXzUEbpLPoONL7ayP2pLITp7vJA
1TQ0MKNBkUGxJk6CbyS36pqV7JTS9WMHk6TTS4zsABgUwZH8Q8UJUdWLJJiUWqGR
wLnnUm5sgVfe74LWzjDEWcLJYBOPnn/382LCB7sNq6Joyj2XF2no/kN/oEN3JdRQ
RUuOGA2ebqLhq2j+Q4bBc75s6W0t+ErkCL5SygrMjbVBzwbaVYv9ODuquLz34eQx
LSCLEGYTEZmg2+kHAQDze6KEZyFsnga0XdfODgD2K0lfNhq7HrMf5L+4iUcablam
MUzScpJGwVNm5lrrI2uQEQnyHYxPVB8v4fZk7ukcio/H6tTmk4UwexS32RQ3ximt
fyflIo+wJIhj3vktUCsFiCiPeQBz0rAmwX2QYnjHpIF6VaAwUP2kmSiBDIYEmWW8
GAhdYuM4HcNTkfvkaBxxSVa2iDhF6Qb9HM+UGR73QYiIG3jUiCcOhU/fX/LpkDHX
F1mpcuFgoRmJ2qCvow2Iad2P3Z84rdVbDxUXk1r/jT+4mtlPdQ+CbunAxkTNV6gA
HDMZNyNrYMOlx0EQHnO9fzcfk8e1qflV8BRLHUbwxlOAy9qnvoLbJJBqPYGDQ9zb
9U+YkofdUi3nKUmMKE1+DpsdV7gZL6/9XcPB7CBnhH2VCryFwTA9E78WcNogDK1P
TkMs5eSIyZuf56ngzW6eC0G0NkL5VUqnQzFHa2RphWBR7YPpBF2wxDsnUM7vFjNQ
7PfT+JqthVrum6VDFB8rNSItjV9eSR9APbUjBDNI2NM1LbpAem+tPM2eNp2/kGf7
gmaHKj9mPkYpMbNbk+blmfFFLuqeFdlfMjkHyuVBVmUHnTvn/PLGTuQJyDsg/SHZ
Y46JyRl5s2qmV5CjMX2kfzZ9aHcoANDWPtRrYxK5sWnLEIpkrbmpIVSPo2s6y3fU
Xmx+MSrNXleU6Axj1cyu/ndvrHLoXRZjCD8PUvbIruUoFWNqoJ7SS8BInZW+FX9q
V7BEJ0s9j2M8S5vWU394dlf+5FlcMFZ6QfJ3DzT3a+Tajpg6CvY3n6/ujDx8eElt
/M9rFfUZwLNcZNlYrRxS3Cpbmyp/5SXasdPOCrbTmPb2JkJme9zXl4sdXMSSn64w
+DxGeWwO4WtPdN/XSrEOrebzNYfLiqwDlEopmtoD6oUmilp+Jpyic8AtO81Z62Ii
NeNC5nS2mQAAayM5woXSkdZ8fHn0UCMV3XA/FagJfKIlv5qCzitHm2+OXydqurLX
L68/BZZRaVm/Wcf6MOqCq+Fa7BJQ90A3G8EsNVtYTQQ/kENJ6gGRwcopfR6Vm+St
uOdcaZQMUtzbSisIW9AhoqbWFIiXYbBwm+qnKp3oqP+B57Tuh+WNjlA7Izy5RLjb
1DujCHwyAl0z23nnck9Ub4NUavtHNZKFXc3k6C6SVSJqz5xE2wnCos0e4S9VHBed
wvxKfuslIt/7gKNwO3SY0YTn87CYEiP7FFBPT4HLjzvcZfpRRByC3fdsE1f4yRXi
fN6kWTumcde9sA4M3swSEIh4ldSovCt1qvwFe/nGkjWi4BUNPo716FWsEv40soUG
TNt/o4k7QvmzMg5s5+oMkQwKE7MmyjmyFJhXTYHAP1NnhVM5y4ZIwJLNrnBi0G9d
iJI8vpCcuGiZW7nIYraytrBU8cAPoa9dkYznRU8fXE9ywPrpw2DMbTyKA1DIjn7T
slDzxOAv4sboFrTGx3PUVAlXQnDU4Nb8DNNwooD2sTBcll85fS6TD6eUgKCUTruZ
4bRofstmQGq9s/0JKeyUPW+ctwgrwqwik4cFbO4JrihmKUJeHZyN0VwP9m0Lk32l
zrBa7NX0+uSgSQx6EOxnt9RxWphGSFaiozL15ci9j+WSVkdnTqYqADQ3komzKMV0
xpUrfXtA5RBtGGioSKTOu0kcJzerNlW37p222UvxMclmJ5V0qD1Kd2RzZ/rLUhzA
jQTnkIfUoRPIQ2OVyORXDCUzrxAsbxbJnaeitAfx8VTgeFubIGcE+BjAZEdpkmGH
m46oVFqqrcOYYOJ9lZaUbSSANWdwU7Rv31lTrFdtmlyBNwPQbIaRyrXYNODVDqr6
0g6e0m2inOd9Ph6D4Cpf3hP0P7pN4FbyvH9bhxpEM5oaZJNESVc6zWaVFAeNn+UW
hkcPnzLyt7CtQz4BrldS7Tlxcljlw4jSPfV6HsHzUx2Vlsd9jDEPR9olyU9J5kzj
DsJTIh3RsmolgyhTUvLmUdG9I/kcsu8+NJ0I3jfvgwCJ9hv3R3MW0zujkAmsYEJn
/tNtOerGuG62LCzREnPqD4FS2I0/twCsxv7pQ8XmUKmzRqyABEV6/2vSC4TM7yVH
qsSfftzSeZqhgQpsNmRNaa+Fwl2XbhRKuBV+aIYNwM8fyS9JY/zJqZaBwtNRKdcc
hL5uhD4h5XL5NbJSs1medPasnpTu/LthAMpICgelKzirLfuuMe2SWQX+aj9NIIi9
gm33SU+Z/9vTgFOwNUglzLnynaEo8odV+2QW1lcIyViIB4GCyn4KYUq27pktOV+i
qyORA2lJc13G8fw4HdlgcHaYUGasiOesfsHVeQuWveiuPni4yi0jQ+HRI/FIO6mX
4tS9NbHarT+ujIrRpX2ANwe7lpOJCiR2OM21THawKUn39GG9WdN4vyu79neIyAH1
NkmHMvWGumiHPiwrKHgP8yi5/IGjxuETxnlkmVpKErF2sHN8npZZSUslQtCgTbsK
u9IVT4yMGXvPBNtdp9drsfE+e7KesPw8xpdclfUahhZIfRSMYCNkqQ9aQoYgEVAN
x1b2DevZBsisYmpC3hqNpsOngisrHlneJf+VbvmoSdp7gzSC7haMiCio2V+YC67n
bVgyUsXiOaoeyQOoll66kAUR5tfhdl/YryjteqSGGXZuXWXiJIfNoI86OptAmSYI
epgdRy0Y4YYo4lEdRmPsZUI/60Tjydjz4G/BiqCsBs69IAXT6cgF/xjw8/o0gneG
Yaysf5LrqKBcRQ0ZvFFWAATc99HyplX9NbuZtN4yl5DEd4oTLnGha/jWjuTVks2V
tmuUVW1vAq6HfiV9LsLMHHpRfiSYPURduW8V7/29HhvKimLqiNLo7vaW20u9OOUO
Gm+UFP3rEbTyTjPYvblhiYE8UVsXD2OIFMNLnme7/gqJSV4CbuFE+oP7rV/duP1u
rk0ppyDTUikFqpkZc27sngPaZqFhv/srQ41fNEqsr0K1o+jhg0wBJ6tshPxSQ1Qv
sTeEcWW4Ub3FcmRWS0218mg7sVq4kKMqMPilptssE9W+r+Ek3c4n0JbUasn/Yos3
NAg20ks/W6rXr9NEsU5uOmH3DFdZwM4zxFqjLsNdwD1agjS0OOZhQ2CTazXt5Zpu
ZHU9pFpPwE04vE/GaGwZyOHCboLE0lNcW+vk7JCgluFgpKnZc1BawT7vY3zRSsim
dT9yDfNW/uc/95eVKSK9j/Il2wisMGz9p91+ElhnODSmsCJJKjWLey422ytKJH2p
KwZZOUBOX+Ex5eqD3q/dab9uyEKv2i/40hbHD1jVkHrMTzvxJjqLnVNzM300yIeT
XOWGKCSDpbqRarG+eyI4Ew1ymqyYV8yPWUkLquJSLFYtWO2/YiV3fKnggI5OaRVg
rNk41TDRxdV4U0/xOqlR1mffinVe27tGE2/M2hWHh7p0S8yzezJUHFqfp7diL2rh
mfcbVT/ig0Iz2U6duqs1fheQhakZkzb4kMENd3wZe2LCj66Idn7j/NA0B8fD5Kzv
Fy6BQvYR4kws21Fswhil1dRZMyLe1FyoqNjLjNAhVcNU+eJ+D4boJIZuJTW3ATQ4
ywSmuAtLaFKUt/oN7FQ1482BE/xn9hKHgJJghBfcdpYTydDDsv2HDMzbkD5j2gQV
QhjigXk2rdmoqtzZpB5uIv3WjqBqOPL7k7U5p1/+iRnsIcefKweAF1lCQ78/J8UA
klIp8ZVfK6YmeaD/MfsQzd7SRm9eARoEnj9JFj8VKJ1I/f12mMUzrrQpSSdH6lfZ
umXNeziH0hruCozRz7IXNApJzAdSB2pwE2tyxNRRTPfZy6Pm7rhXsmmGc4QKn6Gn
g/23vMLRfSiTwiGgPrLv0DEp93tAK+2ypJWlF4vri6HzmD0J8tbdnTuNmPmlxrex
TvfgP2/7TB/SBeQRkHRi2WedpOwDxKwSW0BAYhqsMdBJaX4ts4YV6AmNxYbybALz
nvV4RRmT8vbG5ycGlts/7weLLS4M+t+g0YajKtDwC69XPSxGmfJsZ73tPwfbLxJD
L45Qa9R9vvBc0SWwi4bV5GIbggaYcmew5cbWeIfL+uPMBNNJysYuGQo6lmw006TL
FPBsB0G4MnX8OTjGO+i4XSDypmfr1mubf6s1JuhyOXs8tpf6eg9basZtu6C0uSRO
WkLy76dLcUP6FG1UjALI26xwxQH634Jku5IujrZNXQ+A/wT703Fgc1ZuA4YYX5Jl
E4rLFo1FukCPMaeUE1jtWh8QgWHHUXfFGblS5EHtYlpQlMtZRLdED8vzYSUlh8IQ
Vm6ICuTd5395obn67VYf/t9ciuZun/dVAskHsGzINYj7LFwq679EsEKZv8/AJdLP
sAsvMa05KVKlCZJB8/IeSgekSZMIDniCW6pqXFdirfjzqWH0SNg4yl8+K/c16xAl
jrsHLu2Ad8SfpocQXl17WlKWrM/LeHOtxNPVmUYu+b5phyBKvJdUMynrwdzg8vwg
9ilC8IX8capZLzUfmUprsnmKkU/tpozJZtNJs+psgbrVgbAGQWm/8KUXVxfYvgDB
Pk19N02/lX82XQbN2p6ymhevdx9jN50tF3JKdJLRZ+iumGr/HQtk3iiYWACWEbv2
WDn5rNDC/59+0Yc0OxpWz6n6sU9nEq6UscccJ+hhY5vB8iserxgYxCyv5OCreaua
/DKHbzz66IfaoSuHsvHGOHGODoyYvcul3FC/0PBDtbFd/D++KpjoKuYWqbVh/PJB
YqHJnchWoOg/4VvhTl/4pocjs0Ua8ZRnE35UvwnhdaW6U0ZAXrIdBswEqOD9C0Te
eU3jXoo/GB26QP9kWqGXr17EYWdm6tpSuTrgTq73Vwm1ab/5oC7ywgkUwrO4pTHv
IR5rbHVnU/P8EL6E/QDhnw==
//pragma protect end_data_block
//pragma protect digest_block
pTkARI2tyA2JLyeWjzCZiTzrWDs=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Pf+P3/FprdN/+I33u+chj4MxwqGFhIN47R6Gg9iaurRMYn5ygVmxjoerS+aZimkh
ja+PELS9zDIWD6q9SlNJDamcY3gLXanXPwM7sQn8zM/z78Q5upd6AhHKq/aT3alV
gHeCHreWlcfs6MIvV3M1HxrxXxvtcKaA4K5ljne3zJpcEdC6Gb8rRw==
//pragma protect end_key_block
//pragma protect digest_block
gtAyBjI8bFQl7LQDPJpy9lrd2B8=
//pragma protect end_digest_block
//pragma protect data_block
1NY3rs0sav5cuJicWcwezW5T0BcKAWSO00wGoRzB7Og4RNjuvqyQBvwZblV021E2
wqWprkh5hBc2RVSdu3oYNkB9nupUc0xCykQReTD5ZDB5iC+l1g0cHJAJiJBzjWxj
8AO0ip570/fiw5YLDwK1YZdeVD0Dar5oyFiEirWGcekPM8emPMlMTTAaBV4uTIge
BlHlrIxVODrjhdv6R7NS9n2ivB6KO2Hc3Z4cRsTfVqXMP9awnPt8j+YOjQ9lxKo0
6Cgx9AqtmSIv7k5/kqBSGHDyqyx8dh18LlwYLK8wO9YSwuvTGKU/rdyvthy2I67p
JFCAG94aInDSfEKRIVNtiZMemIZc/SJr0/LvDqOLO7zKAQgCoqwbIUURqU2japBs
rmHO7DOFRXa3xqSr4N9OVEdpbVZPkiCfknXttjrvPdtGYN/26o9XfW0+reWtxfS0
4xj9W2auRqfS/NEGHJsqTOPE1r8mJ6E5JfQRcncdvunnVgApwMaRhTmBjdDM4kVR
cS/gtFBwKoGI7wtKU3V3bn3YAcJn932+ByJTPEsZye7sHnZQLTM2qHsaUoGFQT8j
qc2NRkacJmiTiZEbpsO8oi+YzRk5V5xjR/Z6pmZRVIWAsOdcAcZA2PPjyXgnzx+O
Q6q/Br1+i4TsqmWRyB2FkiOdC3KqmtwOtgqmCZll/xJtBiMLE9WI03oKfe3M87pv
z7+61C54opRc43orcKX37DMySabklQljoJg/eSuHZaPzcJ16oosK6IX+JH7fu7zB
sJGvFHqaQqgdQsYwkgY/r3aid+X9LlVU1yREeDqiFc5zNI1b4OFRiZfE78tL3JDq
KOYG9Pn/8kSJodb9YFWwL4rv/qalpIEoFjgr+7OKQO5wIFgTd37KAmB0LDLr2hdS
sLBurit0WvTCf3d4rpeu4slDeSEE4k16TCFWcNwljupwyjyZS2nyLJpZmczqhs4K
z6Xh2RF8rVunzeBu5P2NRzTVCjXKc02Ap5XPAexXKAaJJyTCDy8TXTNxDiLtSi0k
FMOVVXoCLhvjlPTohvaLYqXh7ZztKcgST7EvcKsus5MkLPYX+WwkZgHWvvbmVbcH
ubAYX7Oe8rS4hnwzRtOvpNLXVA7V25tfc2FmsGqRcoeaSuDoR76piVWOFs1N4ceA
eEXu6wU/7Dfyl0t04hlYWTyaJKGD0hgwAAEeHWD+wj2cEfWJWHpbuvpuh1mlMhf1
8LaOkYC/EhKg73aqrR3+cbQUvRunakUlFp9UOsN9MICk3DVzKlxuHYPIHQetRVlO
t/al9bF4Y+vMDTt5ZRdN4nc44GEELCc9/WXxaVAvW6dOHRDDMjc2OxSVxRt/dZX5
5mcRRfJvUA9XyGGLLdMOahJkIDaWANGOZVJRr6qCF1IHyyxsOjAABUFt7uqfbONN
FnMP++nLHZG2/VIijzVl3UPOQqLazOvHL8y1XpoUOP551uJHZXJWl/eDdWynVh6v
Ed5OWJzxH05T8wcfdiSjsq+XHa3TkvAZUylEv+qrSGHI+zJDD9UYDt9ctzqdHB9N
P5CMQtpAXcoBI+o+EnB6JEKzxlAWUC2dKN3FhyhR2ZMx8bsWQmWT8j1mjx4GqWpd
M9eejbJ8C+1QyQ2lEwXihRoSc9I02Z0KpKlF19V9ofsyu6fIYoCfnswg5FzKqoV2
C8/RufwsiuooOpzUS/A31DA/217W5PllKEIa5MS8xJzzz6E11tSmi6QerbPhpquv
rlr5jeoxE1XSYNyEmjPw+FLHkg8W8MUwxXfgofa/qft/RwWICvd/z4SKBIpr4ZaS
pL1Nw5dm+HR4/Ky3FLbjkw==
//pragma protect end_data_block
//pragma protect digest_block
4kiCT6uutoiqTo683UCfhMj3V6U=
//pragma protect end_digest_block
//pragma protect end_protected
//  vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
zqxiqY3juOFuRd13wY+CpEI/E1qwlYgvFqjMYC3CMGWl4B2NqTQXi1VH3sGAY6jX
9PsupbVhFUR3PDp6knDlG1EDyNm98tl87fHXZ2hG+nZ7jqcKizOgOj+g9diC041v
pLMlxyxfIv8oQoXM4vuyJYIp+oThZomhSC5TC7CILFKJh+Sn0KkLSg==
//pragma protect end_key_block
//pragma protect digest_block
saheLDrR7nL6jJhUFziTWgG5MCg=
//pragma protect end_digest_block
//pragma protect data_block
j6WgP7jG/LRmkImmqV9+jYZw8gZUF6HwtjP4KxEphdnm2irWjFmkeuAdrvl1hEGr
9AqPL46T4hMBj6ioPALhoS87uDsj+lyIdr9oqlKDTdUtTKIyr7O/82eN/7XhFRnH
ydt6C72NFTZ9nb8VwtqQ2u86iHLt9Wbbc+4jtky4l8JEYN81fmsnXEzlepB9vdY7
wQSFdLqjgfeCPQIrICXesGEAep1yM0lTbWja5VOgr31XkLOnvdMLDXTs6o73nglz
O/JbqivlJHns1QtHafDzYjo1/goiEXY1YYLxFfRSA8BSEmcj9oNkuXypKEv4EPGh
K7XbV9cUe75SZZY9VW56NcyF+hNQKWE85zaG/AKuUIwzW2EXT0kbYrncpolvn+8T
vG6koxulKo5dgtylOx0J7s08sGxz4Pov076POSxGNHe0MYCikNn6RotV1Jmh6KJT
acnqvxrcDeWWmy/8kio2qWlccJhWD18TY55Ix3lN2xeXQCRP7D/4Oz4Hc/x1aw4I
wnrVtH/Yt5JH6v2tzMRb1ElNRa64pXDvSOU+KH7FPFlG499nLMfJeD9PhYzr0LS0
pOppfV2rxlLt4NceBy415ZPJz0zRAXG5iJi0nDidnEPFp40eBNsgInSiUqyQm4YM
+ewe6o9TMsRSwlJRC3TrVshUd3UaDlkH/QPG3SAlasPDjN+ccRZOSgKBS/U/BPx1
MU4S0Lple68AzyL6GP3dPDr6NkcODm1+jPRvX3oEV+uJcxAU6/+/lWhd04PN99Hp
1zIljZi+0+RQ2o5fZlVSAR00cd5MHWUfWCGgaNE9qk4A2s1OL42gyq1tCZPm7VWM
7WwQlzLawg5APfxzzfmdch/rxLwa1y6YrZiQIu19aEV/6cI7ZV4QAs4c2mWTTbUk
3AdFeRl9a3ltM/af6mTTLXWbkhZiK12zAncp6EXF5G0OeUGFlnm1+N1NKnLgKdHc
rR4O3FNoLp6GQ+xBORqFXA1b9joDunFPrYeRsTzhCxjxKNS05W56AAehEzCBZEa3
m2vAZZdAfy0XbhDP3lYPQDaztfSQR/+ManMWETyTOk6ZzVlA874YIXaPysLeHEnZ
qoybsHm4h4lcdz/EC3COJIQNI7YBcT85IvVousqQs8NsG6IEMDXBF+PHQgCcc4nP
lRXUB1p6Qke3/HV7ScYTbn7R5ZbvsTG9KPXrTOw5hZWb7zY8qH8x7yp8koZItq8P
2bBsQzktR2KzSYAcYRGYR9BAX6A9UR0UGf1VUV29/RuGqEYshgf7TzeRtHN5Ndce
DeqzQYvHgJiUXtU9C87mnH4vP1OKslWwvCuZ5ZEzlErPlgfhAeORnpMkVzJmc9it
LGfbsXFA10xPyqC+DJhafWu9BapL20LAn6F6TagNCJiD59u7M2k56MImvIjxE74A
VqywodUUXyGMb3JS1GeeyJfkiXLQqBIYspJ24QXJIlfHfq12ULnavFFQTVwBL4cw
FD3Jgn0ezoPhWFkxB5sugQQKlD5fFDr9oWS1kS+/A3DminO2UwiSr+rtboyydzF9
LMfconkZJzsdNOjScKREzFPeZXbjeY6RsUm7ppbwz81cMZIAn7ByFIeLlXwnis+G
Lt0vZq54gEuOnbuo5tv67C9jicZoScnxFgAuD/IIcAWHl0+l2MX6cVj///DpQ75F
n9JzrFzIFqU9tTctcmTSE8wM0din9GKPSR9qcK7K0A0jtbXco/fCpqH16rYOgQtm
QMMy6YZqprTfG3WDJjATHT/Sf7hUYr7E2V1h8zUqW2qTede28FynpliBQSElKqFW
XVREG1CATFWzn85by7rBzE9nRvcISTa7UmzPFsExM7UtycsaiCwA3me9tioTWXj1
WvBUcR+87VDZSXxAeNZpNUe1ki3Qqt/LIlTbvjh+08yZWLGDYQFI4ELqUImUVkEQ
ipnviLxtW2zp9AvpsFVOEMWOZmOSG00xZMdbyW9v6/1RCTRi9japV15GtjBVQpLC
6E8fp5Y/JWil9DY1sMvxR79siWnghtTIBFVggsF5gMk0fPC/ITsydaUiSOkjrX/8
wgICewO9PGs7Z1mnk/mTj1zGCPJ8UgTgTQ4wZVNSHZyPHb8LvA2G2jYPXpUa6zyN
Mh2jObtr7oe8GerAJkjrKtowTK8I6JLmgxL32U5V3ZcQCnxplDRWxEVNpKB3s4XM
bXcQCWux6NAt90dUmjxcvhRZ0yVVNr7gqE+XeLxeHKwgRvmqpW6SKmLXoUsCj6MA
ldoBwpq14mQcAYZ5GbHE1uOcuugkbqEFFAGyYw9J0ngXwkfiVFMQKgVDHG2naPJC
N+Y6nQD5LJXW5IWyZDB+USKGdQjAD/32a2J7GAIMDG8dg7h2N4cg1+aVF8p66ViP
OCQBDbynvsIUyRL4N9uZPykXoNbmzh1RBpKmWP/ojLob62IVnnf8Xz4WHYaJeuKj
8kwZ8uTOJ9L27mw2vp5g2KA+hxTQyqNlkPvVEo9S73jFivloJ9pzYZgbEzq9qj0A
QooZ2uh1auY8Tr5JaZUImbs8zo5UFaJiBs+Nm/U5A5e1eOlID2s1i2O6ml/sc0Bx
9whzSyg9B9U9mIgbxXk+ReBEJJohgkQ3Ru6ZHwwuY2GL0HzaRk5WuonegUMpBGNQ
8KWIzrzxTMCZsIw1gWifHbmGabh0v3J2aVpE+TkVJMxF2Z9sYBwXv99f4hqkApXd
i7YLhGKEDwrzc0x6cqzDExiipej5h2xdjvAWOd/LV6pUGzlUQ046dIcWXHelva0k
pjnYcEl23xLgoePKPP5naZ4Gh33JKZ91E8LsVMFga+sSgGqZ7fRy16y8dfYvVAHA
bVLsWypUi6AdJY4EzKr3K5igatG7fDKiPPjpwYudCl/2N3wtmiVySDGoxRofLhhM
yQ0pHBiL7Sl42/rjcg5K3bea5ZKcLrk5ENofeEBnO3QxK1ZHL2yNykD5wWcp1dld
YHPeKbxDFmLnNOaKFJl0/8p6iTdovuQBMppa85jTxsRBpvJeXqohOFvIIEkEf8qa
HNgIOPUo18FeCYvPRvYyL8tYDf/ZPbMZjmnICxur2Scm+Gh1NrxCCQS+3Gy6Tg8G
jxyxq3duvBselplUGgoyo7FS+UfbfVYe/Qv2Wp/2jLtBTmswD/oYlKOfi7ahNyCD
nMO863pTm46y5QUMb88ExT6nikAHGG66rmlAYci+RnzZk4N+Wg9lKoAsb4m9P+xI
MOv6tfrGX4LclsIgrjdMjOyLyL/EEEzp6Ce3+GqWDT9BvhQFyy3++sIg4oo1sKEt
lJKqSyT6pV6Sf0HxrC8UMursDoaCxtzMJUOgDHulJ+Cxqx/yyiLB2trcBszlCFTy
nTY+KzealjfLZrn98bj6ULO/Dq3knWZAaheKdqIRtAlo5WtDONIQcGNHITn+2rlO
cm95fi9c7g2KEwnIlMUpYNw2MyuCOBzXa5dqYjSioLtImDUmigqubxCZfpYEL2K+
Ae9iXr0MjKndnKsx6nk9PQXcTfG8QEosWipI26ch+Hblj79DKzHwiSiUQmeCW4Te
swvvrX9s43BdwU7VWGJEccc4TbyL0r6Ug4owISAruxx8qGFG/aHnvGrvxV0LPrrA
UW8bSZwjv4ZQXb48GzVWs5ciZjWDJVj0fsTPuOIjPqsyneRxf14x3x8AdmZpNZJj
xAG1WBbc7AgvXhuO6hToZNWmdX4A9jPYyOakxHbut6NWdYOMU5BPArfzlHMvqDBc
N4CHJ5Qmz4q8wn0zthg2lriKH8yQLHZz++DvJnGMMI7mKLK5dO67jK3LizDoX1uO
Pu39L54rvjlUbPIZs3shZCl//nuHhWjov3K9myMd7AxOAy7wbWmwUg9cpW5yYpXw
amgmNU3eerbfmPSCBuRmLdy3GQFzCMsny1fgl38qkVDrAWklTXT+kIL1Hb0eYNw0
YL9mJgS5QWI2Zt+8h/Uz0PZLTa6OUzPBjV9AMRKsJTERRNUh0/cO0KHpqBhj731K
Z1orUvDPT8A0nbtD5UznY5/+y55SY56ogXsiQmYDcYqcWR+abjxX6plFB1kN7fet
i/BceRmOpoqeOLOecYxt0aksITgUq+ZDyegNROuKVmbNG1+dJ2RxYpn4Z8HFLEQZ
yw5HWNckF6aliYQnSYL8WXN4I32m52XqEv4WSQSh17aECvXD1PMNw7K+H3lhjSh2
590CUoLZSAQNV/6d+tqT8IOW2I8urKrBdXhXTfF87IzjuxB6psg88FNjgi5fD55v
M2Vh9L3QKVETXnqlibZpALStDJR3DVSdxJWIMN7pkXxHId+gRqpDUARIN0IaozJW
1k9txm5uMTsukRhI8Rx8mC1SSOsmHdZoDLWD6uSyXWEDa14ODq53epthGovyNw5n
jmdvmB9RLk8wpw3mRaGgti6kHisg3kWx4Q5a+UiuTdl9luTHS/QVLMbw17sZ/qyq
c3rfmMhmo2tCiTkRSd4cSbVDZE4WbM35yEy3B36rR9gzKb0O3poZrB4fbl/jnyay
TpM95MoC7ZJ3MbHnCuhVWPL7XEs72hxRe9J+a8W2zzSwHVBUMmvfgRyLObu4BAJY
sTt9lLDa/g8hER7jZQHCAcaRvZgZFvSpj+J3z9r7E9NN281nB9r0aH2AiKK8s6e0
6/z7jla0PPPmRKMCrZ/BFBCadxpMU+dQp3KPM7dRi1xLmxaQXbiQL3hvGsvOcwB5
ITaRU+MOZj/KOJoDIDQUvspaaH2mGa3OHvovw8xE+jNRht2bX8Eth7nRfFNk/7Ff
2R2uX5ffqE2MKyri+N8TMd8t4kxpUOo1NKk/Z+bP4dj6Yx2TKQ52tYosC0C9VNEQ
HbknBRkEmjKtagp1MwBKevClDYL37MF3qtEFcfI6pEMXPywVJ+c3pOA0+sqXSyp9
u5DJgJYDkSWhoi4NQB+r78kWJpiLr/LH0tWx2oe4wiiWA1B81J/Q5lyoy0xtqVm6
fSL01ili23yvqu72fcvMnIJAq9W7VCikNkKMKgFyAtc6GCO8ojQXlFdxmr7FQDpm
4a4i8GQAKxkdvxxyEDWEIGEnes+dM6gr3O1mCZeWM9xkeDsuIxq9HMSIV+jDNSEs
9c2+/gqqdv8r60HW1e1I2VBD4QZqP8ACuRIEpJGK+nUwLx/uGj0z9PPxeysOyUVV
VjGPaBylNQbe44MuBMbsXsmV3pPG4YmWfBIuxGLFkzZ6t8hHpg5rgV3WVihQBaZl
yfkdTnVxD5ZPyXe03y6DyFVwE7URTKq9o0jmZUgzznGf647tJaVM556KZCLsJ4Sz
i7h4/A/qaoFJvMVbe8biX5f0OHxSimbQ9zlxKF6Evw565oVSYLksJ6E11QWKtU+n
IsA2RvBptoitE6t6RRe+NfkEdRlQFa6FzVvYQZWSRpU31qk4MJyGp67aKkmZK6Vk
8Wr2iya71a6UDxtPtlqs8tESQVq984vtmb4DAtwU/27IFKV8gXADg4Ekt9m6JIOu
LWRQOLtQF7+E/jsLSrBSxIKHQJMa3ZgeyPuWg09lRSg0RS6EMdg/FsUSR/zsuDmA
xzoDLvJJFkhgZsxz8lH/z+47wgk45JJbSh1JeYHMuz1Jr9GNPFwvrh08N0uCLVvr
F3n66P8Mf+i+RcuANLr3bATKmSGf3KxswXUsDSzOsg2Pc36L2HYrrfYFVEwFFiqQ
GTHf45fUxstk+rE/b0DZFDwpaRc1IsfqRV23AdF43FbblcdJz/LFf9ebHM52c4qR
XKJXrIq4VLr/33k2j9k+usq7SghnmcDexDG/M5DXg68gtjqajNjRxfmYJLaDJKpS
wE+l+02FMZhCkX4yeIba+tx2SluEL0tevcaTiTJBIYUjroBiim/u2mlkFv+F0rcD
7GtLTqm8nhhf+mqaqdfBEi0mShmercSIHkvQCx3gY67rxqgL/WNKkB2DVN30gqIx
HUlBjzj/5PKi6xAA5EFfGfq665UcVOIf1tE26Qi74pmsd2ZMRpexCWDuRfkibG+F
/DyLqUCA/TF2mdkbmobo7pn9Regr2gOYLxNDK3ph8on3+s2W+V+dJZOJny1K/tI4
DUbV/AsZU0tcsbNQKnw1/G4V5GqhZPVrFCHcXKa+22KPO3QhqjHkjjePyslslnYP
Jbv3iXaVTxAZWZYsRIG62gUZZbY9735h1L7uWH2cSajCC6SY461axrfn3BxjyZ87
HOHorWiDNEK79KQmH+aghhykriZGHycWaS7HgGsOp6vyIWX8LlMZp7ArB/Cjkygh
PzmHqNS4q2wn/Rta+y/63HSFeULJJwS0Xaou6u49pHbUYT0CwN1S2NVbfIXm+2qh
mfEZjPKLfWyItGWrYDZdNcYzAM45GhbaAGxo3hkmgs73Vh7ub2k4BNeKNogvBfS/
JyVMMY68+yvIEx8XXOCu4ItpmtdRcQ58VnHBNEcP52vectvjdkfxbopEDsp6ZKki
2zS7iPvGFNxW/GimgJ2BucLtVw4SkewaI+UALZ05VG6bzY+//uzJl/vriksyhBW8
YiKkrq6VZw9TnVKGFiAcNxbWLIfrQ6Q6pvu3w1mEoTDTw/C35LdGX3UW1EFkS6YS
xtx8zYzDUtiAyXcf21yQzIFCn+JrYfEaSQRHzGihty37LN1J/ODNobLSA4AEq9xn
tuPbW3TNfXkBAmHj6AnidYSbd9taJ2CnbQvuPVVwK3BAHoePPcFBoNNliV9LbLvN
1pevbg76OqMhmmkgyJybZcvRPDAwNSksCfS1eNDK29qOaS+XTRGz4W3S/3muQ1Hw
FnYRo3yB512LNK6P/ICjZFjTyjfr4WRyDR0CPaS8vBhF1Xi/o5DRA2FG29otrioW
YpN4ypDTwyvD/UxCIr+PeR5sAK0TLzfB5P3BBhtv1rrxVKfYyuwQpEAOomJIAKea
2r2Gr4iVQzMcnqGDoA4M2nwFhBsoacY+15XuAFX5gnEDYd/60huronhoJm50s6E/
bsSC/BDKIsCmDkbFcSMEr+OrCcEYi/WE90ZPrAKKsRZ5DUcbbHT6YfRhE9FU+CA8
h4fZ9cbnS0mGDqBggWxtdEKNL1bt7poTplK6q/iWnDPw0/d7EPRq8JG/9bY0nrUr
RGxGK8FhTAVZah6e8+iGQKYWq1PTXznFi9w2fXqa5hE48K/L2feL4G3q65shQUPx
VfToUD1uN1dxSqVqVyolcGHl6PpRleIgjM8YpfVUI2uqwR4zvQj/ilKPu3Rhu2u5
xaGe9IVMlYOZ06p8Ed7fXHtDOnji5Udz69m4ubYOLwffIybC4r0cteZKCuF6nRAA
vnmj0yZlpn8SLLxzkgQtr6WEwQppq4Ya9J2DRcwFOk1CVhCRcqO/KkQwmk9JexvA
nZNpEBPEepqX4AzLM86I03iEvmia7Oj0Xx2RWIF0Jos4/pBnyV3Jaz5TheU91P2x
RRnJG7/wAaQlbeUe2cFnfDKsI5sunExel92cP5vf7mTF0ArZgyp/MTVNUvxABBhZ
EHayXKrqECIM0cqglGOIGkSqCtSnXxT32TDpKoyvbrfYK6DcI3JVLFuahMUJVKqD
JBC5gfNo20X80RJTSOGNnnCvgtDkv21vNM6P4jtRX8RIn6bXwOfi3N1/W/k14H2P
wkibZSzo+I+9PlSBAp3GkLAbQN2dYLPdaMn/HVVNgrxIh1ehKgUKJKgW3lAzcbqK
ZAXtWO4o9V+5UA2EjslkZczxZGKtL4FjF8mqtltDnjt2iRFHW5IK1aQTSP6fu0Yz
OatTZqDaXpfGfBd2uRqk/KNBtltq9L42LXECYHmWP2ihfKoC+5BN/qH6gx9bfodO
KWkzpWCC0BVHwVplsqXqWc5sEl0n7rc55z8uyBn2Nrv5Zs+RWi/zbHqI4sWnLpaL
HkN2jFDiIcUHen4wGzTA8S6dquM6NKGAVt5Va+UII9C1y1OY/y65h9kkjxZbG2UG
qx+48sO92GjEhcwhN0N3aJVi8FBtdAQpREbeXbhLuJit/STkkE7M9e6oHvud8/ej
bH84ssLRgTxu6CAPpSw+OLFLKOYWKtH8y37mZpcBeMQw6W6AWsQeOIaKPonUy2Z5
qav9Pi6AcJ4x1dP0hRwGKRhgqlSSO2xGWna7YnLmYRqZAwUtkRvVBFTn1PxKQmLY
8z/jzn39Nj8PxRcTc2P9UyTfEvVqvx9nIX3NXdHXZjS0FnoK5hXdyGI2CWo5tP28
WAIvB0mpB28EwFydfjsKnFQ3YC7bbs06QByyopAX9+05DbwB7vD2+1OjoJmuz6X7
Mg2iGO6vmeOF11huKA7RByZcEbq2w2VpEfU/0HOYNGgMLQTbTrgM2g+VjQonQ9Ki
ftcZIDvbcMmY02DfOmM/zqES8nFnuqrk+aSJ5QORmk1P+1+d0UJlEJ7rzbLZ71T0
FKBMFIOvcjkPJoDmIckQbRlOUzW3zkI4YWdx94mQy+P8fWetmL58VxMHz4eiCH3Z
6nJX127zEnSl7qS0nZSGhd19bNrOKo4mxrx767ZlRW6P4B+gsNVwyln91gUw1v1D
t83nY8FS+XEc7Ax47cT9eluOqcCHd4IcNg6h0++kS5aBXlt+AXJj4oW0m1Fcc2Pi
XlrSXQfM4cSXQJPXxzVPNk84jdI9iJst73vbt78jU+mFllYK0IKrkJcJAe8z6jK0
lnY7JCqae5D2TTO15G4UVsOAuv93svN02Ezjh8x4MzuaBmrbS6ud3w99pzIFlL5k
iToVqhiVmvv1WsF5hvUy0gnZVQ9mQtjMm4ODquMgIU484x7MW5DK1R1nQ6fEUtaO
oorK1K942xMTAzA9Xmh8zhiWCwuUm5jmAzZsEMbzKC259sFpITEm+YtSSY0yYc3P
orNkCp0QUdo15qT2wqydMQnrAsqPR/qPgFAPWasvZE2rQOuE2RnGsasGnQaI8yPV
62XOu5EABmrL9Tg73cLcgInutgNRX16DRVPs4/wZ3Qgz6krcorvdsSz5A8DYOWMc
hwW/92OFqdm5DYEiqeMtJ9Yu6Ysjk3/h6piNdAyrYsvIJ9G3LoYrn+eeksOHbHsa
dkQsRwV4G752aJikeqAwcMfOR2kcrr1/sITsMtksV0Fq2nK453uYMv5UBUHAXK7+
lrtWse1foSClXLLu70utJIjgJbsdtd4DMcvBUoqsHj26t3faOZhw7jIwGpsuL30b
9Ly8fUGNTU3wg3gw8TnWAIEQURhixwL59n8vzcxinHWCT/ebKb+DDDEVuWWxG8E9
T5YkvGW+LkRpwnGfcGgVASLyxAuccMiP42N8Xd8xrOHYj28nAw3dyY/X/L3nCZTC
6ft27vQPgfsZGa6PcBp4NnnpZLSd0h8+S5TdsWH1ybetwYr50Cmq97j9wUCEVASQ
+1WyA/rkiK5NjQZrYlytPqN0+xgyj3iJfSM9iGUR/1vapcAedhELxIf9mTYj2E8r
OMoMTl37CDQ2uT2iN6s9Dvo1bB5uW9VLctcjy7yK63oB4iUnHzxDFc++LevKVDQL
pitDz0hu6gxGEYQ+v1DuR71dCLA2m+TWJbkTh2KD1GvgF4qXf8JuM2JfY6ekzFW0
a7jI0Isj/wqm6xRF1IVB6uYc2tUK0QC8irOWQS5Y8PxgWfOz65MlSYUlhYlZbpFX
xWSsoqCh4P6sJNNcmKtTryUPCwSRmfWcqThy3e+jzKSlhVCuryKGVQdOsbqLcjwS
9mfe8Ne1XRXJlH2a8k0AZVhVRkTbYFM0m8nXB3Do1MyXM2jBNEuSI7G+beOjiLMl
rvLNcP7aqKVdTSFK4BAMbMGltQwLbwa6JYrGe4qND17x+Itulcl/x4DTsbtk+CZ3
6gTKNXbFczJuKtK7VgrmmQ0LWxxaVYjlNhI5T1wbb2n9XJYsv68QoxZVvqyB8CAD
7yBZTzbdMG6RB4GitoHmFP2xDV4u9xeLksNqCL/QpeJdHcoy0FDMEA1TI3RS6jia
+nMQ+bqGstKmihv4Xy3gXj/FqdKRjd0ncjie/RD9g/GjDbj3mxM4IYKinnUW9Pqu
FOz9yXbmnK5jOvYN1qGaK+ZJZg5yeu3DdGIhaVwWKe5vICSI9DZWA/cA34+AX8lR
MuszdHBC9eM25zM+UM4COh/37RT/fvCOo6dcHwVfGVrQ6ZJaOsSZTYeyiJu9J8KQ
7wRNYeF7+YqnBPzOISNjFVdjyu4SWCImoOrYydfeOVdTW+Ofsb/O12niAstRqMq3
ogk7Mq6g820N4MedK/313ppt3WM3eIVdGENeZxo+RrG6y3oUOKSqrzQiq7qjPArv
+FC9YN3RHnpt4P1Vtm4Yne8sX5m4pQ0cJ44OBv3s0l/7KQczStzRdomB9igb4eSr
zQWiEeOYUbbU4uKw6rQ+2DGpwoeYLiXkDhxFJGOxIFJXWQdGgbXNR6eXMJ9j9q0c
Dhvpz7IBsqCmWcK8DfXUwtjG1J7tdVeMn48yJcM8DrTqq1en6VpQNUdxL5zn8bD3
gwyGdUdfmo+ozpSxWW6kSchCYmdldtxW+XKX+v5Gh++ZcTX0BXhna2yHQO509sGX
tppANZcZHu0s6bJAGVcDoS31dPYdhWD/hAVvcvNeroeRqE0Cwt8gLC4/wYS4aztC
idZmxNwBD53v5HRY2tEOLEQCK2aMDjtWBDXdOzHDkIyEBxiy+LzfcYvgKA1TvFhn
pHejGJyhB36tKNnr4k1lxLoyB0Z63VbX8oEcFjkpVpsX4gzBTdmRJ/ZwDQPOiDmU
aH02tWlX26kkkvCug/FyQNx6/c6nwhJXYIHjtTA+UBXZmTNVSx+r0OJSbMMhJDY8
ntvZ9kgPErinjQXhwhiF7hrlIGPB/12YTHWS93TJl7046Qv0BOA1yp8+5o1/aa1D
STlQzhKDOWNnbvBr9FrY5kf5C689jmNfmK2141oXic/vCNlNUqX0+f+mLS+WxS6P
XXwM5S3UEyVAhGAn6dCUj6s8taLmG3AX4T/xv/vHXZBFPo7Yi4LMCZURxcmHh0zb
wsZ9l7twfIblc6VGY+4as6iN7ClmNNheDa8kLc94ZLLOxTx5WXMi3o8e/T1JYGfe
+gCt0560bx/JBcicgh+xg6yCMlTV6k/lcmSjcVeHxbpzaxOG+xOlYdiFRPhreFIm
fNfeuA7N1EW1I020lC+45HHvM6t2GyVP+thcALaDVeDNvX0PtVhO2xBXmSvxabdY
GNVv5eXNteDYUfhkCye1XPjLoTxvGbBLlEYcm8hF0hdc+OgpgLOQpZi6HM1Ve92s
lfzTbFzdiamp+VgEUUfMHo1pJvIEkwjjW4vLeVNw0VO5Fwnd7WYK1qmF3iqe+8Zz
nN3psmbxlXUbn9sObCEPYPKf2sQyA8LafCdECXPqT0TVRAzrc244xAL9DC3Pewhb
1TRjjM1jRqUos340r/9qx1CZX8t9C1YG4LhI6BABfeE0pE+g+ClCMPzaQANrKDPH
ZG2Irx03hjWKuJZdLrl9BkQntdq/sjQ2ypfriugXdzFwAb0EwOWp5pxnVkH8wf3l
yswgHutaYPEKmJ+NQptFAFwiRIQI4PuWbdQkPiZwFsac0LCrcjkDUxOKIWxa1I5j
rAVHEBckK+gCCBwW3HhEkfzI343rGMTyNAqs3GKDlFcYj7frdEq13G/9MhpF2yYD
miOSurhbOzpvV7rxxKHZQiN2X9HT0zTrIsm6TrMH8IUy/zxEgiQbZDm5USlN4uio
VU/YkkAlKcJUmO4cepgHJjYU6oknsYlOE0hVnjw7DQI9NUnGp1G3ePGWkmCBQR0T
+zelb70+ZT2YrhlmJ0WLoAUcvlVdeiPncy8AfJeR9NUlVFcttSrtsriLUWElTxPX
sG0/Xjjtew2HPcNMRjLCWJay9IlltILfVXIIQJK5O2eNFbop08iJWFhC9GxVnZ5u
sRnn5FnadENKT9y3JGpjSRGtilg3mk9exsAhYQVa6yK6Etub4FNPP1I60BwJ6FWQ
YXDS4dTSnByQId1Y44/+LpY45GWmKhTTEVoCQeV84MTzR7CH/CLRZKufE080NXhb
/kzjz8QKXhY8YJZSrgCMOr8jGkNLEFvXko2BKENK8fJFQ+2Egtsbzx7Blm8Q0PJB
GktoWX6XwYhX0Fn26KMJhVEOweCQicyltJ3GKfd6x1S/g5KyB6m6A81hAzX6oSAm
tCFZxfx8ocCQRdIcXuYV3pvmuh3i+Pb9ZXXNj1HAPkVyr8zKL6PzF4AkUasi7Do0
c/HvGHrYr7tE0xX+q1oLlXuWnRbAH95t/4PSc5TuwsOqm99JPbNun0Yv1y/snW7S
cS6JZ5L+RGzk+2ldqk5OjjVa7Xq0RxZ9YWDwpyS2A861i9y5X3QCEVr1jccjRGPo
gzE+UOZZy40O0MADlPSqd3irgYkaSnWowD6M//tg/PS1weT4AFnNTb0M09G8Pnxi
FWd4yJLU6lFrFrPPUNi350HnfeMB3MRJgNXhBlxU3XtZvCTVhkYYw7ZU78oAAJGD
lBIPlxJs2cQb5L4cxgOqk7W99MgHIzL4askezKuCurWULm2UEijrjI6QlksfV4XK
ryevjvNyPYHfmlAsGmqDlIleooEhvzKbxsNf5rFYdMB+hR6XZ1FlG4UMYtkVSy2G
jUPSxzy2eXLiTMdEJ0L/bdED9MvavrWx+90aF8YJqc2sDk5St9HsQ/nHVjp7phzG
aSsBl0iJnDsU5Cw1nG7WVHDGc/es44Issd5XVFzpcWNekKcCVtx16N4AGs+klhjD
vgLz8Wa/ei2C2RoDMiJD4Z24P0jSf67pIBMMprpItFdRAhYeFr6Lf1R1G0D77AuS
pVnLNmlo2DD3mESRGFq+xZJ4cgfq3iwslrRJUSk/bkB8nyX5vkBp9I5ExaOXI8Vu
+SwKYKOZ5jEOAo1QlZWtnLEn8gAfMYezrc2bkwAF8D8XI3X13lnBZMkVzBAVSGa9
860hophzEy9OjelJYxvBa1udB2N5zYbuwUOJw/Tf7xSTt7I/dFSnAUOEiLE1MyuB
a2opj/suPtWXQEJaE7z4tuctJhfICDb87yNscsildMTLGACSIxoGZ4AkNImXfBWN
pFzuI4GmeNdvd3XtSNxfQoWkJghM5AF3+QeX6y+LZ5g+8zWO//TGn/1Qudftvelq
6bTm2f6R/xKKlgafIFO58SfqvAHaK/DGKHwQAFshFayp2NxYzKmZP5OPWgRz0jdv
ZPgoI+EoB6yeyE23G62ALC0zUTwdvIa1RX8SKhdmBwHJkM3FMiBhc5hx71KKGiY8
1rxW9MyMTRSEkQXoiFHw0ggEsINtmcP5Fb3j2bhxLcgPILhsEb0l9o6kdLdhpHQL
4ZmKWNKecOieXmvugyUWYOUszQChh8wY9ITcXUk7+0x8PEiETpbZsxuigxNWZeMX
B6GaEXz7ES801dpYpzkA8cjmCUqHW+jEVnn8rtg/DgFhyAnjR2n7k77HOBwf7tiQ
5H8ag5DFt9/0EvTorthCd9cDyDNh4BsjcemWTdMsXgkDAYLvZVP5N0qHTJ1GNi+B
tbWBhalADe7oJGUFDwH2T+hCwQ5PQPHX5ScJVqGQQ4S/L3Nz4A+KMOzHZoBobPvO
IQtqS1NBochiY3NlyaQ2djcJEDs16jeEpc0CVOIQfxxMYtR5BawSO4DYmvxPgSjR
4duAqRIR8bXK8NOfFo10/WlZloCFCiY+mVr1qux0cBna1Dze1DQk//5WN40GvrB2
HdpMHsTB83Ad0GaI6ViWHe4m+NZy3PQlAv54AiwlwbKb8yVHyodJ3otZmi2Cb/aq
mVeUU1hFN8OvCxgp2o8rrVF4IJJhK3b/MPEpvdtttgtl5gQ2vxyB/Gr4DKHiYM/O
AvQserNOBG/rsQvM8MhwJfpe9B9Z8jmaV2sDWsDl4VbkXf0so9jlVI/XuLZlKROG
xNbO1PrHLLCpLKVjG9v3sP8NotnYtEdt+4PIUzou3mMxzDqNzV28RVvxrbgELIDB
QPRSRSrzuhu1gLY7KGDL/1QJbjELhSp/XvLGvgW3BhIQVcgTRArYPA6nN1xdNwbW
etMlu+aRxCD/hSLgS7r/Klg+II9crozzubRvV9sAEd5qPB17X6Ht+mBsADMe+uO9
b86ZIiP9G/G0dct7Kpnat4B7L3fmYID2/LaG1vUHDqD0frwqLq5NbAHXc4T0szbz
0x3QEMG6hn5iCYTjMB38OfpsJCI0b6xQU9HkuBTfQAHQlsZMfoO0aG2RDLEN5LoX
5ACI70iOsNCJrG3IS6tnKKiWQphkLpmao4tCQg68FT5KJAY5gZyHsNB97NB5BnNI
znAYZuUf1t/v+SmVSzHcDqpuODdOGknQtU9ptcSTJ+wcHTB/DkULypR7RIVevqA+
ejjIYqo7p3NKm5y7mAcuQ61YziIhhvvt+bBt0+PPB/f0x+3qMLOYaqAu3RXQFybF
uB/ptXsNic6SPHBYvxMkky8joanIM8J8OomKk4vZ6BlMYGxVTjBmZbC7OsMvwai1
CxkA6WdpeGJlu18/5F2JuLVbItVbOJejtOHpunyZc8r9gFbzQsOZ00ZPXjL3tkMX
g0c+3nuG44utPZtzRSnrofVm6qlUAGnCp3N0RtpoQGAPyAKs7ezSMYphWY/UEEFz
lrr/W+IURNWWBdPkB4egA8DKnK/6AeHGsKI5iZ+VNW7LGm+9S8+UpnPfOKfw2bbI
fpJWvd4uZJtW5lMvJ5Ao3u3cdCra34soisS19o0dAzdZrhPd0C4VIY4KBDx7yh6V
BkRQlvejvO3c8mWVeWhe3aqBaBbJ5BbEDfMoAw19jhOo6C+KyWiOaBnRVNOTD6RD
V5V9f1+vOrJBgnl2or+TwTTEklOJ0Xjge1ActwTLFUSWf4lGOg6hcIzZYIZZsB6C
zDwrERX3tyFZ4/G6k1nG9eOgvEzxH6DsRQI9VisACnkil5HVY5ENPjMG7uvX5wgO
CM1H0uLtK7nIx/vgeVFDpReCP767h3VY0v5eQMtXBGmprnz5UBXyL3GdhDrJenLe
G8dHzjun1CJ/YaxtM/+VHMdLyHrOPbsDI3GXPacS8oNyjz/5JoL1kZu7JP3K2pHt
QQwYgYxGYoIbolZab8AruLcoU7wlDs4kxuNiQoerP+izzVckV9uJMLhiVldtvApQ
ck6BfVdH3yWB+CqHn97vhZ+3X/sXI/SGXR0YRvE3uuJ0j1j4nwOaRiMSKnff/t6b
4VOOqi6S2MdF4o2xfKyc4QfAsw7TBgF8NVzJwnvE1/g1lz1p5A742qbmCv8cTZNN
+0rxg6NMBNOz03OJNiyikd0JB4FykYrzSNei+A07EvJ/PkPUwro/cPV6hT8lgmIi
tKpWdiGxXoMlGOaMzxhJM5oNRF65okOVjp7wM2MxozjYMIxqaHA4LYJWY2VGHxQb
7/QAcob/RQzfjLISeO+ra2XQHFDVHFv6KoOZnKPAyMQMZT5h0vYcDDA8fmikzzvl
7i1y9aEVG45AWrmPKpH9Hxr3NYXrQtwmUqhQ2uHyh4cnwNTJ2TVXGZ3PpG+JHsZp
vL8Y80YP+hTT7gIwNQuAQbSl0cwqPe7a+xhL21OD9fpHEL8PABMvWlh3JPPF0ihu
wmWcVyhOgtMtta22ElctxzV2HCmg13m2giaKqB3bpyEiozFH9hDKrYiVD8zFjp79
TQLAqlvaOf9vCvdSOABOLbMwDcijeLHqCe2hXcUi0ZPzpOw/d2PU0/Rzeuq4riQ2
e4uwy3T6NmgFa/oft9bud8YkV5pbWTURg1x4nbG5YbqPHWH2BoaZ/iVjRV7ftE3D
5k0E0sQ9zIzI+uQazZuY+sX29BfU9tR/6fNS+8cJtkXgpRd9I1r/ky9tGziQSR8G
JYWELq3XVaWpqELcWB8v28QJ8mx/nh1cTXK34wwbQFZlSJGtMnpiYKiagsaIwnOQ
wh8J3hjwq6MQMiyETuIeVmZeZa6OtpENjf5ALKF2MH4yeGjBzqrFDGC4QU32jGka
r4dDcXUL56vFc5nRZeKKNAcJHinfWikbhryDgn4NWbihm2kl1iw55pUulguHh2Ba
yu1AaLCA7WNTjuyYjHpgBiIAfAxC5Dvung9wkUCKWfeSA9yICDX2fpvLWkkYbP6i
A8VwGSg0oNS9pDIbylxWdGVD6xpRZFUy3ni+e9k0Wm3Vxaz+0h+J/lTuS4R737Wy
o2XKdJMEi+eauRmwas6BCnic4HZ1GEijG5fAZMt0h9394W/j7xDQuB+CHhn8hRfr
IWvEsxB0LE8SOfeB4JjaFfO+Dl1h0kZDSufGTAL+vccBbGsJG1Xdc53aE32fvx3C
yMe9EZ/vslYkcsv2mwGdW598jBDBDs8VdY4S83prgnD/MifM5eWc7qnlkNoGUIHd
Wy+p1OgBQkOXiGixOhEIb2dRjyrFCYRSn0HVHTosWyJzJ70gdWEu+DLCBmoeh1/i
RPX04+Lx3fal5EJNvRSVUTaELimZGduz0eKfrlLSnoRjcENL7gC8ZTFkIZCxtGdO
t8mE/Aa9oDzPhH0DbD6Xpv9+9GPB5ol17E3lEfqhqu/Iy4n83K9wzcG3mrtJMC8g
Vh+ahpx9VOAOoFXpZJ7LV7emdmLaDaFSUPFRcBaiq9GvUNDhLeOEbizyIy5GoaNZ
ajG0DI7Ku34JGaboTB4CINqx7EDjkZ0PfLdE9huAgagY2yFEH2CYiyuj3KhPbI1j
zy//mkK02hN+5Of+x9XcaOZVUTvVLvKF5FR0WEtmDmwQ/rZcr87EzZV+2F/aRTnv
3D9qTxyLLpl0PGeHM/v/blpc+OZkUPqWoS9h1soZCUJ6FKM2WS0J9uK6Bfzgu91q
qiwng0zledfajlCsvLasaxmPQF0JJgIkbHc1MPqvRwsmxfCLlTNjIL86ZUTvco/x
HKVwh9PGnIOrODnDD9lF7S9Cah0y503wqJvKFTcBVEeKUGgFLwYafPdb3Nj6Zwgl
SQo613b/SKJIMODokkis82qxG20Fro5gQ9y+rJXZmy1TUtNFxP0vIjkbiKd3jLWk
Pv50zN3ApC65/927xnvSrEtDfteLQJOv+1t+kT7RERBaEgD+lJT+qrgqSC8xYtgM
KnGKQCfo3ouo12tB8fEfl/jRVZ+qi7ns783DRqaOevMdfQ+stny/mqopHomWiQHr
fYzewcghai58R18cTbxv9u6Urh38mbuHp4TTTyvIO3FTwN0xT5zP6HmNNTgy12uD
aA1Ubs7ZFzVJcErDxVjGTOrFkPlDIbd1Zn5EaXlxv9LLrEt8cOkNrbyB+ECeoKDL
8/wZcmSPwAG5eDcohW8StQvW5UttgMhX3zbYyshTAA/yqp4eeh6nrRGX6SrvN9O6
4BLZiq3SQttNnBT3+Yfd7K2WlgXg3wMZY/f8/iXFb3A9uAmZ3dMDkGlkmu/1qzKf
dn6U0/RSD/BBQfIBg0rQWG4cwCZ5lAga9DHYCgqa2D5b4KOQJuTIRAsO4THGRMlr
nne39S3P5kDdMszcCscywpcOQ7S+4atAh9Vw8UY+gjNQtElQAR2tjjX8pvq1oYiW
mcYVvKHjKGxmeSoJIY5WlxnvMviFZ07tQ0/LRXO5a/sspMHEmDxVb3xDoBW8iZvo
/Sw817IfAMjkK0ZZRp1T4sMhWMp0wWY0FmqYBuGwdh80+srlZi57kAITKjo1fp0A
NiyGwOwq/eZfUDcpq0g6ksyAOpNt0HbESL2KhExJZK66yWJfPRKSS/3QWI12Iisa
BMCw4ADJABldLKswChnQYBcADTRm1wOn71M+4wtrNhJiDyGW2JQGyWFeyp+Z0upb
NudMcjtQd2mOuZp0NCt318rVyXPEGmlskGgke7cm8S1Vvy+44Ey9Jj4ERAkIFphd
zfCOqn2nggX5cvrocYSJChnIE6UtFKrmZB8FVKBiU+Fk+ZwUbYdtwZy/scFq0nhf
1I6IbB/WpQ94SmQNJfWBZxmHFn/NJJCy1j/ly3nunn038IOcYHSuGO4NfNeFeq/Y
z4C+7YBrpWZ15rLlkVrkn6W5vnio/sBmmF/g8m2MZrPliwuW/r8F6Dp/n205bPpw
rMg34W9iyD5w29t/XkGOqthxFH/5bxoFZ1qfpMwdnpCRsD2mDgeXRosQLS3WiKrV
di+X9vYK+SxGGUC/AZp7MP7av4XF9m0/0gYbBzJwGk/pThOeNq4VWR8cslUAu1Z4
0ATn/zA0ilJYvWhH+itSuLRQaGmQq8/opndr3Lf2NKyuE490XQ8WYzl5o3dILRCJ
kIxVQyqiSJ072wut5uKwom5MGgR9Yk2jLdnD7dcw5+N4S7+6CT4yIEMHMDlZMTGo
4jFC2zdgHDiavzWi0bT6wpzGSXlR0oIJM9L8PdjSXz0RQ/bn+d4gk9MLBrN9iTEX
UhVISZFr/OrudEFw24k6aPziRz9EEkcawuNSyb6Zj6Ou6AH9mD6AgaXraz0qSJZU
ez+XVJe6eJwPtm8Bz/j1slDXHtvuwUmqhViIn8BENecrbJntKOt6mFbnfVOtu5mO
dvUhE6+F/jHXF4sawUrpNJOAcupLM8BVdXxL0drQJA2rRFi/vcynjMpjop6KVLHe
69rIxgVVSCRU2DSgDsD3Iz7AsPnMaeWVahnbJO7TDof168V9VGPIFuLQXz36Mbq9
NrHByc6UCTlcDPmDIh1bwYsSgClO5dlxNku1CPhXrVxSxgJEX/1K3lGMK8av5jmm
w5dTfoc3qbdbccG4rmrW+R31ZK+bBr0HMKOiMmPJqYZMZ0HojzWLGurk9N9C31wF
vcoyX5UuLBCYi9yHmmQH/zT2bu62hm4kWr38M6tS2yBCfZgWV9lb569daNIE//g1
VkeOaxZjR6XQbTyAUaoERBq7KWk1YYxL6XjVD0q1ECjoDm5k3/p81LpZ8eb+nUCA
RfWIvCn71usx7q6CnTWeK5tT/KfvbpPN//NNAamdKZeaClolAaI3Mp82XvVfHzTp
nzgBDrwwXNeFKpfU4UUn8MeND7q68Kv3RhEs3G4bI6LuEVaosGW5gSasQW30nLAV
p6i4P3ZvZsZ+NB6s42SvkqW6H6U4FnyTGOYS2rS5YKIGqp2MB41N91ZsCXJEYq0u
EuSJlS7Y+Ry9cqBuoe8BQ5oKkX39LYBd/JSyxhXdbG5I8DrPN026Hqfh9KQAqh+5
7Bw4RLAbV8n2lrlyBQPIs0qoK2+1Uu24IVFd+vYnFjy/Z88MY9dL8hw7F0yxqp78
unfiBASu2UJGGU9k6ENadLynqTVZboDuck2Qn5Z42DC4jLeb2j5cImZWJoIDNTCl
BXKzEWG4CifFldR7lRrFRl2LoHyLJrZJqbISnxzCvT9Ye1DH/Rw7qiGfEPpSLE4X
/Q29qxPZv50tQPsTUS23ngBtVg4jEg2ZnBHBQVjCxXMsWcbkBvu3du5I30yw176m
QdPhS9pHVnvr/3PaXq8v5ABT2NP9KJacjiL0FcvxWrVPgR4QYH2n7ba8107qL1Ft
oOJNSG4Ei15S+XJ24ezvGQIBz6gWMwhJRaIvxsfGn1eyDPP6KpqWMQEvO371RPXg
CmGApfZxAyzFTGyzusm9SVu8joHil6CCsC4u0vl/DUJyDNP02atTaw+hAi7Awtn2
pxtKQZhkyYrX61TYZO1E/1qoVo/UfvNTUAXdKt3nHcywLEwWDekZu96jTyyManeM
IsOiaU048oU1/aIZB8rbjGtzgumDBD5VZ4W36BS/62K7zyoXvSlvXs14rq6dn+jL
pP4pwoJXeAif0vnSfKtgwNlwtfMG8+nkb6bX2oDlk3mLWFVQoQ2eIoacpmcdtyzo
O2Z6trwNXLZQjw+DPiPqVjchpQf0JHqtDreCqxTFdfBlpFSzxHvodctUkDZrdq0E
PcY6LaE9Y9M5t9zCB9Q4sX3nxLgBy38L+otiQpDrzFLRcf4jcm2nqVnw2QK1YLOv
ISxxyD3X77p2cgIXJCGTW+F3z3CFcNFkkImpsf35ddWR1AyrJQex/7esjQqspJiL
XmpOcbU1LaIpHsuyoNwoFOhtovtBNPhoHYR4V0XzVYrG9lkfeVIs7mPppkul/RRe
p3+yg6JdzH8iyxnh6bFwKKSatG2EHbrwuHJC9H1ealBOOdnl2uCoZOdSkSJUiMzE
TuN1nl/sw4rOxMO7Fpgf1xivPP0iIvonXKAGevhKrKXMSFRiGdvaq28SFN7uAUw/
US0JeMaILzUgOzcXfSXY4VxF5FxPRUvUuxUX6eD3o/gthdZuNY6wTNfYXQScpKCF
n9kwqbHm/AYSHJunefo3qh3O9GYfeuV/VpMKS6JmR40mlvuR1/KoxCO7IP9J68+7
vInzJYe20DE7MSvN7DHjxuLvzlI8+Q6XuRPpMD5WnsFQrGyBYIMSOFwWTNUtNG9M
TX6J7eV/EnTGBNKrj889eDhQp9y7GnEtrwp+q8daokUYo2Oa/QsuVVd65hE6iB+C
bNRQdVfOlcvFSWCzwXPj73RXaVHLCh25TC6OoC041BQoe1Q476Dw7U8OvvCB0hVG
KqNKnO7eJVOZRVKip28A+NMVJcxBHWwhsj0dJjns0op6syKlfF2CRSJYuWn9xh9k
L8kDc21Hm9TzhVzZOcis7IceAkohIn7NvT5Y2EabkUiU8xLGa+559BE3b6CQZcTB
8Dssz+ULynzw/rUqSwYT3gM9ieJDwBKhfHIq2TVWN4JntWB6L93GuRFZY9T3Eeyb
j0AIXImJbvtA9DtfOz4LJJw28BcN6ftBtc4+ZBXxg5gbusSS07Mpp9VCFT84rDXF
G5cSTZCKlFgCNdFeUZuE03BciBAdTsmcH+t3fCQx8Pde3KCbHfAgTVNzWGLrSwlo
/RyUYNAY3DbeFLtmNlaPKeMhziHyT2fivabVEd+y0ihrZRdvHJ0LDcvesWFx62CM
5OIiuo196kZv940k/p9hzd4x3JbbyHVIC04wSdZOfUJGCgKWiwsbvL4uPAoR9NNB
gy/HtWPGO0MpM74wJDTdD0ZxYxB3yNY9jxIqO+NVMR0i46ZUlRYpW9UvZdm9JNFF
bpy2ckjkQCwJf+2hJGwHfpA0uxfAngxHnjRbRJ3j91nDcJd6kQWTB/p+l6+5LvKg
Hwj9hsb7Pqki2do7V6jgMC5TdVLdXcCCdVDfXOmeCvJoRC0ECS83dbw19Rs939pW
Zc5Y11vOBaWGE8tbQe5MYsVf2BMk86tLnM5TYQrtWxyjwl0O08jBsfX/ihu/ftpD
1vssohQiIvAPky9+QLog5DIdm8dkRAr9xKJ4Aie79lvwzEu9r8rMCTUVkJtyXqB7
dJNCKpM12GQWHh19Zyc2dQqpQQH5Tp/hFTlYAn0o3/FJo+lCK10N3H5lqnDLd2bj
2vKRw7eRpWqR5MhawwV2kDOppxv56JwtDNWpXcsliyrOcTL3IJpBbEMh704REaWI
D92IjwxNtbTq41A5pyF+gWnQtFymvmDyWKjN4c1Z2HnIqFBB8Ssm0Ruy7J/R2/MR
WEpCIkYoDhLuJEipxEoeUgK284HW6KTimvBokJqXGyF/IV4yvVnbt0veFJ4z8j0c
jUts9ycMO7U4NK89KXE6xHZ3QVf5gXyXhi3VEComqGxYpVGX9AyDtv4YdRvOmmkg
NHKqBKdwmBEaUaOpLlugAwH5Ojyq+MwntvW+FdGclwEL7ahS8QY+Laqd7ckAm0yz
GIQ+CbKdp7S8vZSTjUbvsipJBY1WXUbwq6rvT+ArB/f00Ldt3RE8lo75t1Zngtv2
22KLtbZ3rSjNflo51lMTSfZ8zMNAv9XG02gjuuJ4/Qtask3d5JaCQVHcWDV5qkag
zCB3D7Udy58W1TH8In5d6m/Is+AzKw3mO1C0Ps0zBsk0m8zAJ26EpdALOln9kKJE
F/CJ+kL0HJPDCUAIKM9frAN/2Fi665/wdKmkc7tG5d/+xmPqHD3SvpLFVe22Lp2t
oRSyoMw36CoQTjge42ggi91TwfTkNEP6wM45MNLSaCduGVINL3qvVeCfpQ4jtqQl
WKksSCKBtyY1u6V5vp1JxzWMmfOEh1LSwqhVtS9nl5v8WNQulGuMeklhm/GSdxiU
YTfdTlkNV2kaHVrg4bwiDR9ZdPAHPOEGU5WiOwpDuHFm1Hn1TKVo+gCdpRbN18A4
C2PSRhJQM/OQR9vDMbAEupiq1UPid1lrIHFyL4BpHWb8FZPhXuLFcGOCuXEkfzwd
VwLne0+o8xM4UAIm8CB2aFFZHSdMrADGqDn7cHeYzBf8EBmfnnVNSJ5o9Kk1OQSq
sZFAXFrrC98ZMPQyG5r+B77xOFoAJBkk1MdfSfNtx4C6lnykWTbpq6zPia641ogk
h4EcyLiigBrYeoCVTitRX4sU0/swL5DOX1DTUJYCjVhxB+hIs2LqEBbSsRqfXJTQ
FcFBwEw8YM1RNlNDs+UhVEL7KLmYEIthalWCm9yeqaYxWgpeXCjEyLt4ksBM5aH0
2EgjZAQwfbqHkaQ+fbWp60RzYP/9zCQhH2f/ouPI99GXtmi4OzMsOfDmTzLUKbk1
QKo7gpwvcl5GQk+OQNkEQdvu3xogVoP2BcNEzlcffbRFXU8Qm2cUzJo0HEu1zLHU
Ow0IxbVUkZYy4u08a/CaH48fhH+X3aAlWn9DUYvxSE8lS3z9rFODvGJcxuMRdJom
Qlh9L1rlCz/nfK+4KO4fi12V5HOAPcVWZzGIf3DL/1NKSKrggxsT++jZgWwSEVUR
Xaj1PXy5dV7LceZwgn5Vw87Lz15p5vJYw5oRc4/f0995TGRUHDUYBUeX6rjq5wJH
YLe9ca+Row756lhZKNzbUG98DNfGlJ8FTSTq5TfxTAX14TDz7TOL/gBcSzSPZah8
CsREYi8Ipe29rrKzicbVWLSbv0PYl7cS9BoMpC5Vn9vWAxFQKquchbD41EHjDcUA
SSzO47xv2e0B7r+swqG2SXGDWEbtaGsxSWDtpiiIdRBkNkN0EDym2nCV0L2vSlJH
QON1rei4ylN87btHlYKM/j2TWaE4jFbcC8yfiB8AEFvQ+ojluYGAVGTH9ITCwQhI
mk9Mm/ycjwNj4+/zbsWWEMnMITVLylFkaSabW3LpRWnGDWvSneURsuBsoKkBvNCR
+sJvOfMWBrXy1MWNc+vzZNoq2saj8iVbeiN7tT9cZ77YDGAjPwhEFU70kCIW54Js
p8/IVbv/ulVTWRfQcTuMvh2ZQegdMupHY0tXffpHlWWGHQdil+vf24W0hXhFavv5
FzwxGAh2Ns9vEMnUb1VPUCPdpcQsly2BYIX8yytS7NJVg+W3bRIhIkpIX4fxbk9n
MURfeoxkKpsuoAyNiOXKwS6aNHkMGSm/ghmWzfBRvMFI27Gv9T08hYkVJCngHdP8
jnkuKJVxv+EUkgCeT+cEG8buVaKr+dcdQCcTJ5pId8JOay7qyfF3QrWiD4ZGYg3K
rOj9w2EM8pQb2DsTi5NjTcuhz31MIwxg3hTk7U9KHcin2cnRHQVVgoaUN+Ttbsui
zFWiAL+t4MlAETWwXS9tvdpeBdEtT8AlJg+e/taYp3UR/pOvGpatDpk3GIGFcnH1
nHemXrb/kO0hVg7nJaKdczLLGrw3lyDxqmygpLFPD3tqFzH5irRpbwr0XfLZaQCy
VB8KxiFg5usFISQCGYFD6QYR9Rng6cJ/Vfhph3WaE3Rk3Cdx9bbhIX3blHOGBlmm
Y4Ha84cPrLisdWIToiTDk6nDCaa/rCFcQw2jspPzFXJzd9h07/UK0qRgw9zfOb2N
GMirlmKSwsO+LTqSMfXX0G4KKgOL70vbCg+L8PNdjk+YdbakPD91/IPtR5vRA+bR
4y4ud3uG3z6uh/3jFkfE+7k9vr5jsZpfOZi0vTK1Ari+8hue+bOiMEoQCxSZztEu
AGZY2Ttqft7x2hldTCASdvzMGETNzaCmwnKoOlvtELPGSj31hDaNBBi7cjy05mH+
GhOU4I3eVns4PxkTGSoIVE4gM9YjV4EoDw23hz8XyMvYwMacUfQ0X4HEcyP8wR6n
qbhu9io5bLBxMoelwW0oez61GjmTGU/0S9wfhLm4vmMlcJkjPQpV2mNeJ3VJP2vy
cH9wrnsSxfOenXrwggWZOEHtVllH5KuCyUHHw7DWJr+A5yvFKnOv7cbrD1Oc/Q+Y
O/YX9to+vOd9tJnedDSnYz3UVUxUYtqUQfXEc2fNieSQDukSlpeHlmfhJQP1XwW3
/guF6EvqXr9dyuRCs+xHjh+ojhf+uzi6dO6Bn23/iXyefBTzTsYd5G4HkCxF6j4R
bpnFtz8nctuc8Hry5UaVeIXuFOQ/8D24ShSLSPDKHahaIU+MWnX+AWGCHG1DXQoN
px5EO1SqFWGPTCR+8DDpSHyEvbLmBoG8SrQ7ZzKDgEOfmvh8DXUBRgAGw/vCyEBv
D9C03Dkop7GBjf9y4Ej7vCRNEF7wvUMtZa8f8mUrgOfRHUqCbLqaSdPWmb9xeqhU
fFz7nsvxhlQ7OPhaGwV8XM3HFyKUxLy0rn0SgxWwlRunJXPEe/5+65c/XovgugiJ
gPGZD1pyKg7kG2ipzBWvrefkgTTQ4FSJjUBYO0LfCyxuiAPDudEMsT1dFx9v9y+B
h9F2GlPQ8C+CArW8xI922NBlp9MCIX0k1mz2ILXSQmzGYWCEGPe3aWxfGVqjnfJE
+kg1gc3rDMIHG6a95y0g5nzdzXdBUXKl7IE9jhm40hIEOyugQLufUDoSRa5ZxgIS
1g4gdE0BOKCP8k5gxSCHq7FoBbffDuuTDvbuTyLNn4rCySR0rG8SVP9c5Xl197G/
4Wkyb1e2xtZw8rcUAvCt8iKukUnmnagsn6RCIfmK4ywiwm5GGGxoC9w2kzhrAhDg
V+oC3YTkHkQpW0h7uBtL8oOynV3F4nUo9JE1jAExn9K6JX0+pgb6N+wszt0Q2G8Q
VMuiPhJqX/utrxnf7Q5GnTjI1xl1QUP0h5kr4QZeEfgppEdF3PTNgbO6luKPFI+M
tongxbifJQe7ZMA8l5kh8Ujk+d2ecIRUq/WmHl1olry+CsCV+tOIrGa0IPrkfWeE
1rgYDGBP2O9VgtRAvsxEroRqEpYTnKNiH+6niRXhVdmudD0qUNkObiSP44ruGT5e
90CsB3WibTvJHf8QIyDtPDN4W8TZfeC0aIZZoRC7XEhZoCv2HGZ3O8dw0AQjqT6H
/J7knhty/gT/lWBUtRHv2zSg6iwSWMXdMU5TZd34n4iOM1nvzJU3V1kUgymPKXAX
YfRrS9x5WM7dwqKdSB7BZNE1ErxEAPLzTt5iaQiBrTXyRIW7iIwXZ+NhtgfglBYe
soeEcD/ZKnfujViRYwCpCDWAgNSJiOnt+4zpyYdBJUW3Qta7y6BdyEapxdfhmZbe
KqvRU/GUMg+Hk6alLmg+n0SYMt478aLcVH1EIy3xOJK1w3GEMGjdC/YwO7o/trDa
ivE0JVoC8lTXUYStKCuSM1jfJqAhRr0IXrHduSCN1BtXrNzIe+xvFlfiIHFGgquY
K/BOtF5zI3ei7YQvpeakticVPD80T5wQIH7qg+i2GFAwsUDp9hHZHMBivQdn/IuF
Rrf6W/74JuJ+PEHnMvCPlYBM9E1PoE+9mAeMVkC+NUJW8H8nalolLbYh0jiN9Hqs
bdsVc17xuyL5PJe7qNXorBxohLdMz6jfb7zwGqZ9E6go4Eoqsj6mdrnX4CFHH9+0
5sssyZodEu7xJ6U6I658rzFrFfe2rmG482fq9lWUEKHbdl35RAtiQiSdx9kLRq+E
QdM5NZofaMtT9V3W8dfV7KehrYqPBRHooOUkNZDJSHEsqCZCAchCVFa1oQZuaYH6
8LuzDYOnNXltKWobpdeGTDzj8O5rpUtGlCwJ788qzznBKf/zv2XuPzu5BdOzCUh2
EihkJrLOhE7ahgoFTFQ6W8nn5PfTPz/yV5XfMkt6Svig0pqc1OwTkL0iHWF7i1ez
kAdLBzYfkyAnd3u03pbGs8OjRQcKE5EarwV5wcT9Th4Qgvm8Sg7YsawPHCBCvmMb
uBKQF1TNEXaz70hUR2wv3fHmKIxNNsjR1ZYVgSTfbw0OnMdX1ZQ7wHSl3qJvZVJu
r4ncax/DzBwiy1fsg5V5I9WMatH56h7HhIqCn7XREaILihH8QeVXgVChy8NkmJq+
SFREXdACqcqHiJ/vRbbcKBMF7P5KByxOHP36WkdMxOWiDF6fvpUwifVbKaYsQUG8
Glf3Y0EddWX+UQV0oQE9BALRia19t7fg6KNDVt18Szoixas5u2WHlE69x/Kp2Zxx
IDhHXGVw8rQ1CX0t8z12jYi8iCISdjgj/unhitqzGdLCIQAq3WCPtYhzM2GqTqBB
BG5KS4/b2xdR4h01j/FUcnlLdQ0Rcuc+Z1cBuM2lhsN/04YTCU3njTwJ9DRMGbbQ
qY5++xAWYIkYg9wOiUbqYEBgIqqQpVMIFMfQROsceSVAE+ojqenoXeNivgHD6sId
D4Zhorm7Rka+MPDfslaN0e+WXmm/oDM12e7L1c+JBblEpmPbvF4Znt+uBL0MAG/j
nmojTgQaVN+dd/Afou/bShvktjiUmq+NsB2phgyWc70dFqCWu4kURbpj2gMZfKT3
zPdOf5isu3kWc9DjIGnQyHcpvYyi1kTWvA8eTcgVppC2OjTKoTO0SLw2fVTo1rXs
IjGHdfTMJO7n7zoMxSBO+Xla4Edhj3nBgCHYqeedKyvrgMkM9zb1CLWwhV7PM4Kl
H9mKcgQnphNQnevdAr8GECNu3ZTC9oex/++34dLnS3I9t+irxSpnoll8Oz/S3xZq
x8KFQBQ1zanc74XrOyQiQjalgd7V1w2hHDRFudQliryjTbhmk0u/DIaTvMot61aN
HuaR9A8EgkdqzWhtrOYKxODOSzNeAGh06vTO2rOXVEgSEJm/cokH06hcv5gfIgeE
SRlVH9mNiIv4hOVU17y+GBT7T9jDwmjK3fOLt6Mv3eciUlYdxiNxFnqMYfC8JZsV
Qm8IdDxmJJaaN84mGmr469ZzlAsKnGzJr1TA4muspvAvI+jKBvK9BkR6N3G0qKmp
nlPTia//GhfPS96Ul1XrYsx/NIoH5a/MMskFcuw79sLHBJ1Uy7zmsj8S7rY56Gfz
XPOvLPbgeH8LUDuyTdZMKP2Tf2QM09qbAgwWtYHWUPGOMsKK7r2HcpnHesyDTR3+
xSj79Gz9k3J/6ta4Y/1TGvoZHaPqwNAsUdQ4d3CJrdf4flP8egTG9f7s9NxJKt1z
UbXBhcrGRda5T1Kbbimc4CzH5j6o12PgUYxExccZ458DSOhmabEcdKQeqjzK3bqY
hY2znrpv8WN5kwmKwmhmbsTPo+gGjDHoa1yzcPPmddeQfagY2GzgYW89QfRikFzR
c5ifN1e7viS6QS/9ubx4UHDouQCeSN4qz61xzf4vyzQfx278t3hoqR9s4IBGc6b2
TjSzfZtK2wLGwJWVKDFKVjDxWbdgAWGIunRPAQ1ohW7a3qMwdPVQjyplIicUly72
ddpvoIyWm73stDOwRgqh9o6uVUCNQNa3AOMafAs+Smwud/vtKPtT5CPIFowDNlZ9
auSPdGo+bCzyOkFrCk575TsFh9VxHZeTq1maf5OOqc1B3yEM5um2bCqiVyeuYoof
2cbDlKgycZmzCGGYttijBgvKIn1kRL216SvqYrYroALitNPzAa2YRqA+xcIbHhHQ
P1OI1fjdgbHoYLeQ3smYiQma+ohnmKj0YfOUb8i0NSFeGB47yZNpp2/i9ePBY9l2
VgrDKS7g85gtf+G9yXdzFWzcGAbHjusfIy+xUgeE/ER4jwvG5QEQMZTr+jm6JO11
RclqlogfZ+yKNJPvSo8Oby3dT7jVsZPsnDBxQMO2k6ILR83ZaDUbYAVpXoOYdycB
12kkEQwqUjPWowc5HLB8ivaADBs8SuJi5i7Un+wxbjDVBHcJNz1CgiEEUg5kovNh
T1BKez9k9cCaH1Jekc1ivRzKnZxhdCQzvPvONBYUvgcgPFFEnDbt3SEf7JJ61MVl
IqjJtwyqHejwcyo1XTDZfvui5gUbWcM/oRCVWrU713vN2tzEVU6BEPRI0GzETX8m
XctIN4acA/bF08bSVCE7xb8TZ9IfMzkcfoeuprBuXg+xFG4ZP3wImuyRYPI4hLZp
mY7Tp4HRKYYnA6ETut40awIn1G3ziHEjOJs5+Ukl2akDCfpaK+iN19s8QoADPgr+
5wDb3tITpg0H8XBsJlbE0fbR1mNammnIKOQzoIYJfh6plkag9aawGCnbG4e4Q1go
xh9/Hti94c1h2PpRzDr4FgnzsQ9xGgEYq8aegYgNubxVh3tc2BQumrEv6BugOmdG
Q3lPoshApXcVKKU66QfBUjHr8A56ieFDEy3pHKnzEDfCZmm6Khywe3/XrvUhbfVG
gD7+Q0eLwsIsPZhrC7Ko2codq9q1d1ZKW1B4BVE9ZyiMdXtRZocQx9qcKg4P33Jf
72+k+jfeiyfQ2sHwS27Efvpr7LcUGCRur7oZD9juvRUv3EXl9KolIDGgrKpKLd3W
5QakPHdGxtZBosn1mCKBcD33xKjb4JPLrFD6Blcuve14KDc8r40G16gP9UAQcS5c
cPa94+dbgQ9X0XzjBOM0FY6T6ufbjIFEBNMw3rlmtHEsHU0E2dMMDIutctFqTVOh
2Z50naaiADlZktNxzK9fz9j9JyKPv+2bVSKnM/b+UPkzweNBz04GZnUZ9cS4BKV8
K0lxdEID3LtOHenKjfzIgE1S38yNvu+8PWEYBY+SZGp+NK6HclP36iRqD55cHcZ5
MdsXDoCB9YQFcbEk+DTOmsIAxpuaaBrnuv891Ur1Ml3ZzlP6ZzQaTUmLOG1GsZ5s
ArGX+ta7/c93AwEpcLGPnum7RjIuQzsTOlWdgO7NWRf+MJ+8FToZobkseYdU9VxU
8U2B7lYJF1n5TIj+ZRP2Vfa49J7jJ3vRkgWxtyiK9le1Jo20BlmJ6ai3qU9fKotY
blg3vSyg7B3yYlm6nq5eTqwhovD5fMGQG2IvWawNOwjiBbNiYVOH/FLNXRhlxBcZ
HDg7RnhPGDiFSP60srE154Nf3X9WiOXL0iTTWIqXLfsnOPcLZx5SAZM2Hg13GZr0
m3gL48JwKiuZeZwN77iYtmLe2JhTJ++rnpsXDzcKfQBZmlafePpIWpn0484HZrJf
fSoNZrJbqvBX38JgCo/vvjupEAwDBKPHrpW1RUxdyqwxHodTO3VeDtc2fecsnFkq
LjFjO9gGiti6lFvFIxNvmEOKN3clxODYnQiJv1UACK5KK6yMeiyl/l5RJnuHxUJJ
UZuTZEE4P0y/EAiUexcmf+wMwzw25X16dvmTFkUfu7J+L+KyGk2JJTE1yO01Ll80
AWiCePiuuEc345XqJ0pxtg1IfgQBcqi/F+ghOLhEO7UOuGwCJj8opTNIPMimE3kS
0fVts0DMywqJuYlDnZyNIO5tQ8ffKraJJT3293mmhhF9dMLgn8AazCv4oDBMjO4A
KV2FclQbP5wKpw4bxv6DJVB/ObsLWCR/qmaVn+ZGA8OlZ0d4fKj42Umg30950VjU
7NtA5JSnacL6iFiz9dObGZp34LgfFLn5TjlqiV2R+MMffqSsB0EIlOKnTCxPkHBu
lh3hFaPFkygkltBvmpENfOKQ1XkZwEzfBO5aQR6oQTtdJFEqYKsWqX937whzObsD
SFXQ5SI3noCMZxvvoKX+nTh9POn8rsdMk5d1w9BUFMbh/7UoWqlo+Yogbd1bkPN9
n9/vV34PsRy/vTuxE7vRYE6bYMs7QhHIKvFfBWkv12jyq/Od8yUPR9RPSgcAw6FX
8EBr8P3xU7sKmwwQqFlsl6N5dK/ltw9MGG7nX+Orynhn6aq54YjC/n+8cbDqo73d
aDuWL30QUYwQZgDgJOpagDY0wzBXjml90DEA7eeTIfymK9y2abnFZhyDE1p547Fh
jAezNbxYKv5YUQdI5Hl3cvQjMGVbUP0XInEW4Tz/I01/hgKEHfba7wOrVzgy6PvJ
58/QbhwrFYmiAU2pZX2v6+cVZxE0pmbvN3xFetdqtCHd78Uupq4M5vDsmhgPc47C
qRYsflDqzXA6bbZVKqlSc+P73RF7pE0wbIBl6xeYXE5+ln3Gm40oLIe5AqfL+ds5
qmc1XPE6DP7QSVVyTsAhFWTTqfVji1JaKlP7D2xZY7QU2mo/4XQdki06tuKoDpSh
Y1VN+si42BspFdXqKyBZkEAVCNNDZNZOjui+Oj3mdwwSBmwQbZ3X7Wamz8kBxnj2
rHV4YJfvOnhb3lZA4Pyj+zSQlzXXb7P6dmKqXBoY/KFT69hLRPk6SBak5LAgtVZQ
s8x6U4ffdY3x+eltFTsKMvGM62SvUWsUxkbzHTWQH8Zuw7uMe3xFZUfSGpqvIFxy
nF6GyOfho7ui7qACTQ+LcEDXrO4w3DsD8jDLBPVLXlgC2EwWEngz0JQvv4PxcZyN
mlLfvF0n44bwMbeosKaOPuWWeV+pwCM3gmxKsK1YAnwOq41nbqdBJu3Z99KwuCii
2kaAqH0P3IW0lXIwxBiVRDTDLEspCdFyNjEk6bBPLd3Tqhf8nnwbohHJqj6feNPA
E1razXYur0hPrPvwcLk3q5dDxkkae0J50w7P2DeFdLmHFIdEWaxjHR9xHiWarf+H
vizRARnDEt2gK1hqRBoVIy3OVp4Ms2qATCbwaoPyZyJIQS1KL3zz7PmTEIADIn5Y
FNswDsh2PnyXOjy2dOdc/jjWFX1I0LMN7AvoIYtJMimvctfdqkTEHeqgs/cJ0cX7
Sy3e6Be2o1ga72SAof97I2kS5lU8MpWqQYW7y5reP8z/HYN0jD/h3I8Y6+p/UUFi
ulVrfCgOW1FNWVN2snWUUuiIBpHzxjMstGfEiTG9AwqL6pKJMI7BbTz77TXsv4h4
sMWStJWlTziii8QubPwsJrVHNzXMjgl5mfEvFU7dJxWsLxmCwT64PGDDhbk1y3MY
KrpB/3AsHPJRNpy1EN/B4BTxZKcltCfuJ3wZ4imsGsay+vVoOatt6z2wGgcy4dad
YLfzujJIECj1WRsUrdUrdz0OueouDKXxQ+zUPHbwQ2EsXrgDj74fZsPDmvkwRdz3
58clWHgmWFWyNhBH7xtVZCYKO5GiTUF4S3RAwwHyhCHMBSNYWs9Eevz5jlcoUnw2
yHQpO0QUfLaxn0zeDtBOLB66nKXbdQ0zOPYAyBLi+ymkpKNzVPe7SQxNFTMvfs98
yhXQ24LQh4ehKZfwdsyhKFOReWxa9GiTKFn2SeZqvmZTQe2UNySZcNFqgV+77Qup
mCRs6fMaZyqEMWMVdImEIeUnKAx9bmu/E3BdL4pD2HYUUx/5fw+SGRGPeQKM/85Y
PujBnWz/7G06ukSYIryEXXAySl2DKvHd/TFmR63Q0hgCHKNT8eTOPQWAn29lhYMl
nRtd3j7hPyMglnCBsVqqfmeUkPM8+ZJti9fglZ3HkKTWSDWeTej7KP5EMoo42vaK
IoW1yWoXmtwfWoaIu8lT/4qWc0fV8J+InPhPb92tqMiz6za9bgghO21Q3f80f59+
GB3Jjj2qEznncQYt5MDnFpC/G1nrTfN3Ef0KcEraAaFJrCn0jmqqIiUZ75wAUWnq
eXKnKlhIt5d85Rf2wb8xnEKr4hQFB+ldQbznjWcWTHlGMVfXV5BwfIV+t8pe8kBl
kz/D9c9StKo4G7fFbSwHdgyED9CgGsbTTPMZtFeEoZiRExjXIcDoqQvvHQpzoBOy
31N7JDJztLKBm0LLzUMLJ3uVvz4/9J36/nCIYof7zpvGZcaAQniCxVAhjMFTQdnL
8LFPFVMNW4K3gec0zqcA/jYUgJ6QRe7pDYQoEkqXuigAhGc/7JwXp/+MnmURGFYu
5AMFzp4Na2a6f+zGfUdHU1MWM+P9uTxlfB8j+btagAIed727vRg6ptAG2Uzo8W+1
DVDUfJCh/kfxQwMSnmRyeJM1hXFpOKs/t29NhGmh2ReTn+RJipU4GrByF65gIDRu
yotk5l1hdonBjNRzsdxXQIcDnJAMJSX0bzjEJV6OUCHpzbg5Y8UNuoqPtH7xEbLy
PdhskmCznSL9FlCh78zbGVlTuUHl/J5t4vtSe06zrQBxJ0dAV2nR4RZggeCzgHoT
vYLiQEuLvkuBQThwHglh4ABtSliAMWkwlN8gsGL0FJ8NYKs8DNbCZCpQxLbnWmZq
uxznTE1FSHokpOlgUKcWjYzEmaOxn3aXMvZOV4C+W6Qs7l7mPzP9OAU8ti12/GkT
k4mU166Xgtdz8c9d8yg/JZ55DTYMPdUVolZhdGwMrjIPlVY489rn56RgLSMWhSv6
E8daVZ8CrAeGVwOkSM0Rm4yiC0q6RkVRODJDpOFKCn8Uch7Tn9at6Pd6gPWNhaql
WKIpDnsZaKoGMIHZ+tOzDPSwVk83VZ2RzW606ATXlJyKq5eb5gaYTmwo98zOCP5I
7vBcLJZv+R2Zy5XwWwz3NKpaDiEfdGQ2v0RU9wiCl28Qwabe/rdt4HJ5DcmNhO3V
b384YDC0qxL/Pjqw+hd89Qg7L64dmBgX0rMGTRMpcJFo3oPsiVixe1b6QIiJVTKK
C/JXePA+EVlFj8HFhThgsYTCa5JUgu9KGY1TaILJQoNIDcxJouiMk4rFgab4WusH
PyWfqm+2klf6QNp7TH+FkyOh99YWaXhz71FOBbUSYPGSTUT79D5imsqWEe7IEqcg
ZaXBrwFQLeRmzKFEpKnj8MxCfE59fPrxuETy03PpQXlloNrGPF9jTIvW3RcN6ocR
RzhwwRvqW/sJ2FlV+41Vp4X7dezGkUX1dCF6t0f8JrFfxdAjIq9qVKNkzVBnAt3o
GXF94mexy7NW50puvudjcW8kJykfaS0jTFKe2NAkJmbNVNqn3jb5uL1S96HZUp8z
lOryaMlf/pfEvOOBY33ghPtggig3CtnlEx7uaOjEbpJzX0xoDP6c/6sE0C+88uX+
FaCGtqcPzdhycjGj0XNWBRauEwx6QjIg0obgkSTl7rfIinIV++HtVzSwlW3Mt8Mh
VRbOJCIpuA+EHEvROHD2VXa1bVG497OMtYoyeYWcR6fHpuRcB74RvXZloLaRdFII
kisKlabmWkQG0VrmJCZ1fEfVffZ1tAMIUQk0TgZzpK3rS1aoH2j7Ue9ZPB/YS3he
W9EZH2WpYTT7dDEHXLK7d105WN5hUQ9kIf1Wik+Lhc6Ajj2feLAKVKBRIHKOpX8M
PQwJJEEvTTRHml3ZuUt08Rkd2VBnat0iXfdDMgB5RHZ0Hj45Dn/2c7RkFBh8IMWC
JVz+zVASC+RsXVLqm8vq9kxhdJoROjyONkJxDJ9lakUfRR2bBC/XTfv4Ioxu6sfd
lmnxTtXggWVk5yfWaDIt/O/ESss6fFnfJwkbc6/vFUFFHCBMd1qd8H6MgVZdSGyi
plyLBUGqihU01zborlWWN5gDH2pT7HVzxnRLCyFT+tbWy/woKcsmQxqUkxl4s4Ss
0v4XVshP589H847zmKy16t+dtCAn35wgtfIGM4KHvNfw5BNxBOF+QwxRnrq6yhhU
yzSaTfV3J7cExgDrXziyKCki5fSacN91uxhwGwRdG40rSERyvELWVdNDTkkJRYnb
M0EMPLJebMc2Am4GNNOAP/Ks87bBemPlD88Z0iCtN9fFR3PnGPxwJQMRhop4URwL
h0tiy6+P+O4zsRGD+hxelFE43QlLu9PpLI21WUNOA3g1K5t6v7yv0MUz6jxTWYZK
acZtHxRWP17f4zKanvUlHmDjA/8qwbqI5DM6n7gaen+ru83pBEkcV6SL0Wokp+P7
+nhpYphkvyrndTzivpIImAdCuQjytw940+ZFRcSlXBQRdNyVwna1Qpknx8ENEcsT
D+qV9hEOoEpmvHpmh/AHZeJvcreZXtjtxcfJkJAK0xdY5yoRDHY/oMzt/hN+tzJ3
LN51v6MdPCg3mK3gEjCpg+ALAPoQcxvIMmqZxO3xYekvPKwMjDwKOoo/xdjHcH9g
SN3xLZQLWJVP4lUlH0dZ27zWVSsMLRBg7y+2WYNzwzZIKhISBo8u1Z/gWXVgbl5i
/lcnTQZZ0ycMC/+o8me6N3o2Z4i73isvq7JwdUVGbDbtAPKR5q/i19yNpUFmmauc
CndHYmwdlEiuh1bc2YeVoS1F3b4CG9z8f7uzH4XEq02BZW8C8PHkdxG+Bys9hVO/
/vLEpjd4SRiEZ+mBRzGcgRRkxc5/cljWZa9KojLVIl2BVsDSXBEIw/t7A8+NdMae
ng0DQBtDEfB9Hm+iFx3F4g8GrHHny4v24E8/AcHC09d+ddqMxQehG4aXDnjxocD9
Xio5gDJDNIxyTiKry/t4BnMb2sIqKaUUO0CfUsK2XbcihngogAFt0Za9zVmYfsSQ
GwpfY2t4D/20q8Vz8wWIJvgji1QuEI1n8S4KCGrlv/5ewifx7lUqFklykTzcMYse
Y4GxqQS2pKTujpyFJI+nzSiOYo16pNDNEf3a1eH2WS+x6nSITgNOgZEoVnFv0BWw
NibMabWygSVkhxO+cu0PyAArtsLCJ/kMoDsqowQfMoYP/pD5YWuyqnJocMlmbPId
FfChWeT70lQpIb0a94AulLGHJVxyRenH9+Md7mLJ6vFHIh303IOrCsw8Dk42KIx4
AFpDgDsv32Gq54GHevceoLEoP88sL9KOUKkiCT7PmyqW0z9ZhcFf1/h62HCJAui+
cSIgnRtZoS11AksfZDf1S3ISsRf6kIFJcDptbKSbRjZ/8crL2EIKM1uu6q8ZUvVT
QJj8KGkPpVjNy47ifJO1gPvyrmcUrbWgbFuKfkIx/0Jf8kiILca+3g9YVPtWf2XL
snMAOv0ZT0WCGMdXVYrMaMYOC9YnN4SdBnuRtos20MWRj5cNFXg1S54uYXSPU9EJ
dq3maKrKO5lNFDRz6wZIcc0kIQ64drxJD6EPF+XFcOPuy0E/Au9uWgXcXDh+yKK1
aOrH9wZWQ65KOCRI9xfHM5Zu8Zp9fswcBxAqe+fLoUHN7htqx9NMdA8RfhHDl6io
wIMpvUwM1NzXTVL7b/143NilDJJlxR93hUBoXlrBsr1/GtKu5S0NB2HTYTfih07g
4An/dtJydkg6hfPNCNjPe3e8yF83rzIusxsnHUR7/3/UOmaxqMWb3NLF9GusVBWq
YhK9c2L0nXATVWRrhIE07Lu5/2DKSlNVkDq+tXSi08Ktw6XYU9RT26cxSLVG7COv
HB4lTg+lY/EgY7qsIrkfuAVBhZHpW41fRSYJ0/IXxckhdmPBSASNGDlLxkMVOdUZ
8nkUjFAiJqBWbdx5Im1SBbMmyTAS/LOYear1OywBJPCsTYCRPpCkEfVXb4uijVEA
kHBjpmdpCXsOT3MxNQLpTmWAcR2S0C5F8D/ThzyHfmrA+QJ3FucRdb1hT8GEM+Va
U6PPjN/xrF9oR9aWOpYmfsYP0Clucumi7aMoSdU35aJVe3FNAuQnb6NSGY7UNu3O
hJ/99eyDDiY5zGPQXs7cIsIRSp3rD64Z1riuUEhVvWxzhTIRAG1iMC4itLyqeU/S
kAbfIw8Ccif7/BgofDWMiOo1C52VSzDS/shYATOmuFO84+gE7DkUiffPB1/yr6WF
pdrXPTYfiTBZdsrGWThUK0eHXrbfDSd1nuA8uXmzFyh4stGaJ0iwb2QwNL0u0rlK
2b9wpHbaMrrV1JnwcfW41RuGVSGWR7/s63gweWPsQq81qqYK4SdRv8I7qsa0J7+Y
+OBRD1u0cJVPEuSSY3wHXi5EJ0I3mhdS5AHtaA0biveMugCpC5FDS14cT7IHy6pq
gOtLeG0ETMJPSNHpn+dh5d7GjDAe3NggMh+xbV0OuxiS3svYsd0vKGJ/pQ/dHj+S
33FXHFoQgf7UpngOYZnM15wCuy3oK6bnIO+YTxgPKDNO3ESGLfuwNkoSoKdpwWwM
NPwurJFH8S1VVLhdGI5Q7pXrqSPus5ciAH1QArOmg9DOQkEJdIkEsRBljMABB2W6
Oyy8ZJl/4tp6wsx4dCFoEHPQbOufukW/QBnsdAdQL9j5HLZafxawoIs1F0VZoSuB
Bi0MPDlxIrXw/4If6Edpc8L7+KeyeCkiNjEmTD26A73UNK2XNm0R6diO558naouc
Gqjp22ZQ+L5CnSa6dsVQIzQ9+9ngzCjxI3ll8Vk9Y/IEhM1/4maEjTfMGvqfWTdG
NxO9JE6yROtdogHwkCUkFhb5hCJdKELzFJ7B5cAsT6+5/qGpKfw/sCrrS9vcWIk1
JYk4fP1KfIgFIhoWp1iRM3cINLJwaX6TXjn1YJndhPNKtmsjuJrXZSYZGvxsUXWG
uVUNFn6WE5lqdKlB9Hb8In9wRIHc1XnGFCmXMQrpEwdJ+Q7tX870D7qs8Yb2rrXs
T0K/ByBc1YG1LpKpewve7FVVC+ebUaH89I3LcDArs+5ZB873TUBMOuFA7ek4veIy
bBCgjbZu5W8XeSxKVOm1Kn6PbYjxkpDOyO80iCm/na40XHNVlSLKmwx3HKboj8nr
7iD8URD7VliToLutd9bPl+O76jZWr9PKgcY+VP8mVo67fxp3nNkFFMTZCc2Drp27
sAHyrVxm5n4XzhBxUIstxg/xcxVKUS4GlqZCLZK0ug1x77wsdkUcRgGK1/4JE4Q6
dY/GDVcCR1Q1woDEe1u1SyxtbAFW0Lwv6TUp54CT5ov19GWTam9OjtFStuClQhWH
N3v16fPH8nCGfACtK1qyQqH5vYbqBQ19xTkqVjYTw9Yp9C7c7y/gNmL40Cdghn51
Hr17m8bpg1Dfn3Gg+P5IumF5XvOnKefBDYWgFx5LVFJg58hX+0ScKfWiC2WPnMxu
OE67Bv5sIv0fOuW6p0KZApLzFrswbWZn6yzr2NbZKbzWaHlQdpcYXEfueUBgztf8
i3p8MYJGiqrDbaUCENYmc8vjkAL9qug5QLPEgh8USpFYw9/GqGbQp0hiKQ9HGT6e
HCkyalbFtD3Zvl6fDHVpuy8EbtcO5DFbklgtSOWyobx7D+OBfs91B/9BYf7eiF0M
F4CoL7Bhr4+TGtkGgMeZfjtVA+3l/CGZ9rN4QSy92sBN5VLVSlk6lhq8X5bUQqMk
YSmgVUfxIv4ejR9WJLdZB6PoQ4J5dnjvZmbiA88Cj8+8lWHmnpi1ambFxbzMAgkr
Z1redjqZdr5Ii5afVP5vyr8fg9zJ86kJBRWu29A5R5dY0sGUN40YKRHbj/DUVyiL
V3Z2+i8Gaj/vBITpQg/T5DZ0kEM61kUmaCpgI6ByyYom3f/e82fVVo7wd2gRCIzs
2IVVn1uLEJD0rg45HzzAsISTey9YtqiK8il5glUoankN/XVnfUhIQGNJK6SS3XBN
/yj6+nloI/ldaXfHxkXtrkSLb6GTqYdv/YKIp8BFYysTmiZVBGDbeTwKcb2HyXSM
DCsIzH5tYm9R0DUAKnMUO8EbCt7ypcK0a4rz4wdV8cLbIJuSMbCHK/zaFPmD5Y6i
mmFw9l8c9UaqacZcQR5+4BQxmy9GpD6SxNcbS6szf0WHQAS2D8i5zmo4g2ILPrjg
whmCtRAkmecmujwl1K/4fSfk94vOK8Ok+0i15v8UAsn4Ngny5flqcLBfjGxncx+m
Qfe8gnCs01ksNpN011J4Z0FxLzZ3Gq/cu8oZfhpha0Ytow4kXfurI+VHjc/LQ8n9
gRnNQgRAbCA++9ksfO3q8mKcsj008YMd3yOSPdsplzw+1aGXXgr9xHhBr+QADt0t
WQppq97f9iBEf5XXZKyXWr2k5/SQawYK1G//khudNhBAO8LRyVT22fdju8JKgb09
hYescGjevvEs8XJlVttrZuVtO7/woNriH6MIGvSK8B+CUzc8U2LT7srbMLL8PY7o
Fu+yrhXQI31SKKv07ZDWlPT4eoeV42TNU6b7ww+mtYKwTZpDvYWQtvihbuA7xSgX
LSLTroAHb5339s6OgorZyukUgBDbYh7vOxTXpr2wOOJuRhcIGB1str2kO0xOIadc
6/BWbwzfEd1B3NDp6yBu2xk61IZ8j2TXykaUQuY1b44zAH+LEcplHFWivTfQtHi6
yjnwUcWkMXqhzY/l/AI3KDqyO6u+6Ztl50RmYG6+oKxK6NpA8UJsHdPxI7pSzB8T
h8kLECGQKg39IbZtAbawO5PitQ5tSDDqXLA4Irlj/7YeHvmIaxRjchPjOgK8eh6z
/rZjq6wYocY4/McW5VW+Nvhu4lpnBoq94b9+GHHUhhprffdOZ+jsGxb9QYpE2ULM
fgfDjWJZ6MSevmGWz2frPUeOo08qE5P7IZ1FtkEthx5/XSGo639UOY4Hg+NPZeyf
495FXbsDg9DM1YW3o/eeIUxBU2rHxJ+wgpCLUc6rRiwMsWltutAf14fZuj2D7Ubc
S5RmJIXqfit/ea2ikkpdYk2nNx4DYd+i4yrnbR3f60ueBuLTJuiKs7yuLQrG1TIv
wfo/2G/NMPbmW2FvyPCOjOzJEKWLKb5eTbeDhg6Nmti2UzkT0y5r1/PLWqJq3aCz
lrctXzIEtVUFwsMjIFzY2bOTsn3cfPuq41k0lrLh2vpTFBAzAXzvXightkEV1NCK
eS7hFnj+8afta8ftiK/swf4/+MAxu42qalEnXdd5DQJkRovlpJe+LwLI3Gt5nyd8
wawWGFXafOVg4Rr2rM0dPRrJXfdXzZoUaVzgnyUSrIEROPmw9xfRpX6BBeQ8lIjP
rM2mYEUb2IvtLjvwCiAOrQt+SFXBi28LqjZ+Nx37LDeZ7FXLkv6k4TwPq7Ki5upl
+cW+O+Pkd/TgKrnh+8/uosPcQ5kCX6eMv8vua3oGlvuf9FWOuawElpt3Y9/UIVO1
WQzR3nyShqz0ZalMt3dmRvDtpEU7o4e7sKMLQYxQeSLgWXxKFQDezzk1eIoLTqdl
J4pMML984iUZSHaC7So6MRG24UNUWwnPGiuMa2755zUayKcw5NXR2nR0dZU7uumg
iuK4LeuI0dycFdQVuXbHxN6x6tTVJftwRNX+REWiqd8bymXux7JOwmJa8eMXN9Yw
fvbC3cHSwQm7Yz5F1GOPXCzIe+TdovJaBSeO64GOwioiYw2MmSOFnV89UOUURLKb
St1FIBaaQbtzv9arfSXZuuvICgTDhDrbLJ4HJ8ab61hkgzG7usIUsvfzGsWdbQYB
ztYpFBkXli54C+hjJecZ0XoWypFVrhtXnAyCRd1CJvH9wRpeZm3D5O95oOCGwdo6
C27R5cFZyHvJvcw7LdW3dAMxnPexNI2cRh/xik8PccSEMShV52oj5S5ZmqAGQH2h
NigcX/9+0EFJ1OpNhm81zDr1VNhPZZj9FOkBYoCRII7GSxPrdutrZDkfCkR+KCQ8
WxdddvarIZ6s4/BFjJWKIHWHxg9Jhy8AUhHkh7OyJIuLCrQDr0YUQW+Gl8X2xOWD
LYIaqd9E9LtA0kIcC8X7q4iSQaNsGEN1XD+O8f5qYu7oCPze/VdO0fJX/hVEJNLE
lXJN/q3ZxLkfUij0kPxDreMbWFI30K6Qu/4m0qEIlB/Tejcr4NKatcupU6u1JrdG
TDaXBl4TlEECVI3PswYBPlsq6kjxDcs16ZRbGNFskFvAJNouZGXeJzHg9n3QBjOC
gSMaawolmpN8Ypm/hAtylMDj7o4di2vrEMRHMDTTU/OlzWwHBTuGf3MzrpbAZQGd
P5+wUHeBvu/shnQf6L84PNz41yXh47aTovCv44aOYyYc/3+74gJXxNZmzriqDmuJ
GMtVNsFo+lYrc9rlGcBgV/LuqqRcNuyaeVk4QM4AC+iRLkMhfsiO/U/PsS2VK4dE
4SfXf6c7IbfiTaRRO4FJ5UhxquID6JfohLBiJp9n/k3bnz8gCoiY+pSdowasUTkT
qAOCAksJJQxeIjlRwvfCrPYr/3ZfNjxd2E1LIIFeUZSl1QSXn/pAwjJAW7anG1pL
b30b58EM5IS2tPOTUA1oPm1M+O5z0s+Luk+YuLMnIjsgx0I3RUvxgW9RQpPetsII
fhF5VvKd4CNIOWbuzNmaCviA2SFJzJZ7yN22/hpS48YYZQtA7GG6Yf99R39C/MM5
/fw2l1Kzy0J6prurtixEELIxsiVVFPKml/ZGPXRi5Rp2bcp/eiA0fOpm+4kT/2It
QWe5YGW2tFj53azXQI8Jjh4P9zc+EgEVQcDMlohY2sMe0attZMg4989Vzu7QXXPa
hwj0icHnd7Bx5Ne8V2kADSwr8KJNRvFoX1T6b9brIxCrmgfnkI7fLUknXsSUAIM7
Gc+H1eIU8Ws6mnN63F/veWMmF4ecmASL8HphCSNX5vntmU17ZHZ70qK8+E4yLx2j
PR8b4t5+W582MUTVO2GswU8dfvvozoPwJD1YABZe7Yc21yZt0t74CF1NtaJiWjw5
SSGDxhCZF4uxOWi/PVD266cAfRhvLg5Ge8aQzZo63+mwByo0hqKSwQokRB7HKtlB
H7aHuCHT98dcQDcwmO9jqAK+lRoxqxJhjJ3HXqzmMLgcvjrvmLu+ciK1oJaYiLeO
5JpbPd+YKFMYCnkcR1jvz45ZRzvPWjMIyx4eaUc/uyvTfpS7XZ97LH9fbYdoKYM5
C7M2XEk8kLKciR6Ex9JYopOwMsjfS8AcjKqhWNLqBQiITAh1Ldz6WQM0Gpqby8If
8MEe+NQoD2Yl6qnY2cz9zKHM3GU7wlF/iCUcJ5uWoLNP26u1E4Qwn2jXv7rj1Ohz
9IXp1N4BjQwbxAs7cd87fZr9c29Q4SR2sNnqCY+eLha6doH7w/NdRb4SArOByl3R
lSbvg1a7Ns+AcQ2Oa9yJw40RcRdV6bBLl9tRVOMRSzehaQsOPL/UiIg7IpEhsCvy
e17IAUmbu12K7cdF8rXcxvMcN5nDuhFeuf4W/tx7zVy6xkCN4oB5/cwmdQzs+4GP
SiK02+clPV4sGf3IC7Re/empecuI6xs1fxU2zYc/mfAZYrFftRs3Ut22STFhvy67
UHcX2GgGy+TNwnE4yEzZ3DH7Tz2zOFedGrsX/VRrUR2ZlB32lKFcB46D1+GReB7T
GIk03HUZlSsLQm9Suh2A7HNTU0I9axceLmkOaxqrD6det1c5xMweks5nzGi8K2Iv
r6KHInsNOqkJU0HfXXsLW76qn+sXjurA/vC9xQoOeIHg6knTRs7s8R32Lc0yPj0+
omyI7E0ASvDON1qxI0+NUnzutLCLgJ7tafgvkKHj6foFWroqZl7Mx5E0MZ4uMKNg
y99G3YJe81pg7FRAGALRKHDRbVw7MD123fQP9Y/iQqff1zzlHJ5PHpM44raBEP/j
b1zazHFjOValhztHr8huxVpc4GjFLMmW+cWQNUnF1ETJfiwd+Tck9SiXK5T3SDyh
E7DRQ4XX0lN4K82QHLA2qSijDH+Y8PlbrydPtTbDhxD0sF/FRwnaLgaUho/wxQdW
Dvv/Fg2sTa/92DhbMRmhSotUGl8zI59aMk2AGOFVWDrU2KPMwMu80LWK5dtm6iXC
YCq6hxHZ+SAaHuFTBp4e5wgDZ0hjFmXpveD36dK+eT6404p8beCI0BF6zmv2iuNE
T8q4dDSu5L7j3ywS5MOQqr5dqIdqUvofGN/qTVxvKRBB+l9bCqPaMkBTl3CdZ8/k
IBBk5s1lDSTGf0qq3JieTicTsX9kl6QVXv8iNu9WD+84510wJrwhCW7mFaAS4Vzr
6LQ1++sDel7QvhG7vUt485M7C4yoNQ5saPHEAmd9FqYEEJKFau7gjSehmhs1WgrK
9VTiFDTX1owlufjPNc2Qodew4UUEBUV1kh9v9M6j54XmUY3wJQ0tUhK6FCFTjOHa
4iyC1Y9udF4EUMDJirZ+FdEsydB9HXC4CELlySc0g5ZJcwuRhL9OjlqGWIExTkHd
KFUlPPe3lGnPVuNyXwKW+xkQH5NjOtUROiOG7dKIq2+vzRNGfXVEgR83mRRXkGwa
PJ+z//mQP20dA2j5Cff4hJJ4uv41KpVtM4iUcvNDvZgAxik2W8zura26IoWAiglw
GoT6xrsZCNJNFWQD4c/4Efzr43KIVdigWQl2xwtGM6B9VL6nXUN4pHZ1WNbBFd1J
W2LSLR0b6JR0NLpwGitSvDzPTxq9Oh0RLY2ismYEy9xtyBPSlD34f0NAKrJo0OxD
g5pwKy0nQybgSU+JQIiyMvqEjp4W+LjbwetKkXLjwHL2AK97qaJFutjtcRC4UqQn
vuOvg9wb4UPPsRqjM2p5Z3k9rzT+L1suKbiz2czJoPZplO9X46Hr4MN0N5WIAZhJ
qToj0HHptiR85+J2IJCsrYJT13al5spJ6yvPZZ5olBr7Nlvz5LTS6atAK0AXIoY3
mrC625DSOx+qVT9mMg4wky7Adaidu1AYOsieJa0IRYPoURrByJZNz1+jtTJt7sKl
aE3LFp/i14MtP6rf/GDaiRpwXv0uYLAB3ZSh7s7A/eh3ubceUjmRNsx/8SM+L/CT
qdsYEGT7WZnOcRisOsfRk5V6C0j1K76gFyp1PvzovOoVjycCvbA0kXNVPA+yEYbm
4TkuicWptU/hAGNsSN2OBxAPscVmDTbNsFK24kyTxjATcCK9rnVLcKLxniWWTLGF
6SocptX8oEU2A69bFELtzNAK3f+uWg71VoLlF7bywTljP9GYFA1oHEiEjsDzsG4O
QdirV8xybYWFs/0hBTum8z3eukeNIdfTxcXdfq8KFnX7ycl2en6T32JGkR9Xvn2r
e4np5xnKrpqXiYJRO+hrB27EAdbjwFaBv5Sxg1b0dtPrQzjArATSzAJClJUXXhob
9Q4mCEJDzAMlBiXxPjMlvoM0YV8CDsBZf0CUiHRuCGRckMZGLoRqGAOB1GQMDKLQ
ElVXav0NxNMEwCHg4HX4Y42jy5quOudg0aVU5BVvU16jiymjlsmTzEillzJr/kuT
5M+XiTFjbkiMzPyVN5SrG+OwFGC+BZljXko7jwhqfaKzK4O417KpqNCT9QUjdTCw
/ab2cqOUsTdIlLrJKi2qsDCod8lIJKxuDgcF+dlm44WsOmxptvL1StknkCsrjOXz
+VhwdGnPY1S047WkMR6Sm+mkyGO1jDbV7cVxFqucUDBdccNTImIWbkKegK1y5zEt
+HmbzFXCEQPSyGIp6W6F6hqXh6yBBDuhsb2BBdyCvEOFrbJ0nUCeEKn0zsKWwNDh
mEPfW5FnaJPJ+JjcV7YsZc2cGpwiaMHYlJw+40dS3IcyBzP9NDekAYlPF7QoD8TG
eRTSlCvWuM2IqPTdbmBIZw9emt1vRNQdjyeDbGklm0r/V62B11fx/2Uo6WR7T9DD
Mf7T91EDyMAw0XZ0WW7DJYKRYE3Q997Qpe8u91hXatLtqbMMA6l6ver00kxTAyVH
TGxHx9FF+0ZuGyIm9tUzrCC2Ofgo60Hk+2Y2ba3OSkud7f5KzpjB7nnzPx/UoRB3
TmzeNsoWpxeEiy5vQLdWAlxHOxaLh/E9HRGwNlnBdzgKO9uq2eXOu4kK3bduU3OR
DDjkCNCz6VtPO5luEsLNk8JkEHcVx+Fwi6r1QEuU/izAqLMT1ZfgU1cdbnawXbmd
IrP4PvN+tl9aT+Xw9zvoaVoI7yosh14Xs2Z5xn6NpX0mv3RWQn7Ui5guJDGNbUCB
xqJK/B12AQ9o+a8cz8cb1uO8F8QHf+nIBEv2NLjqkbSdDO23ZFsBaz6pOxKJY+pE
tr+GN4drnV013RjGJFs8Hwo2gHhxWkM/TumaqUXCVJmYGj7oHVXyZ57e289gEwNl
0RQ/K0WVQCEOQbNaEHv88jx0b7NV9/HEpDI6JOZBgKHBAe00lLZY+isHXX/YpvhY
E0jZGYnMt/zJAa/7amYY6oNI38q9RjN4aJZssKuWFuq84PfZDEaMCWIBVHhDT8D0
9484I36VdFY0x/n1F2bSainMtuMlhsmUivn0KW7BBMS/XqdoGF6Q7H7CNy9CilGK
f+S+PZXK8dQcjDgnin+ZkM7qFX5rmz7YO6YwGM3BdfG0Aq/NqGc4igYsKtKyTLCL
ehkLVClYIukckGZfKrIym0hZ+Rq3dv4BF8knkhgcaVyX5IJ6z28jbpJMp+MkOl1j
CMUonEE3/7AuBHIOhAitJzW/MPM9kzRya9LqEruFrIRtiB0diGEAL0lY8umfBkxg
lY6ioaVEP8J/fpn7a+cbBP8+R+LT5vfgGb2TZD20yLcxi5G/tIe7c1HyrZZeSMdT
c7HSeEhINSPyg0sCdjJVN2nMXW6GjtibQEBf0FRO5cOcfC75kdqSAOL6C9vhs5R+
0Fc3IVSl2S4loOSsMukrP9o0cG1YgNP8ltx9R+cw+1XNJmCx22dw/p19wcXrsFfs
7g3PlHcHAvA5JcvOh3Crr8ZoEYwbJUagZVnizHPo5gpyenZDJ6fbhw2vLPKnJ+ve
/LwqkiANkCN3/MP9pk38Zj4rAdCgH/04NiM01WJ2Vt+FpSCJowke94MfqWFgc4R2
+aXstnEfXR+SD2oBHv+aJG090ssh+bTCX115yGgDqzORSUhRBDQYM16qPK70LxGh
pcvv1tmdV+mx3Vm4MbL3f13UIUaMZRz/N+Q2ffrFNRR/rZbeq+20efenwHECiMsx
p0tpSyzRY5HuS2U+aK9Q5uzdqHwhg4qkmY5kEAUXlQQtDSm9Vf7pf8Q/t+CkmuDG
MhTiUF2TwWTZMbRnw+/75hGC58c1G0PsQFembYd6+mBIZxHM+E11j78MHmqcOFR0
EGr5In+Jjl5ed42FayUgTNNxxOSKmSYs+BnS2R6+PhITxPT8wpvfyxE1qNZ8XUvl
5mTQtR6fyowmJ3pRkWtRUaF+P/kYqJmfvPKJh6rlXVABrtu1kj3ndgfCVGZ2AoPF
p2JC916ff9UDOOnK1eIKuJ0hJYkMR8l06IOSlB3rmJse6kSyqtWhJoE5T2EGGLM3
6t/FEM6yMvpNe44qjCcIaIxrTuFsXJ7NLXx0VZnKqQVcjreZAFHiTzuklKKMK1pw
wAvhfTto78papuqcWYg6hu/aDdDQm5biIETfKt6gwJa2YjR8Gda8eFE/mXoAdcm1
aehs7X7IduQlNtFO9CLDKJS7GJZBaU1vZPD4DP6/S6UvK16d+q9H2yNzDAZNzlae
Io9lOEK5vHhJUIpgswNLsKjK2y5rQBseX/jUpdrLXW1/s9upupCC0YCCMIYqwrt9
9Dwz/doTyo854qcGfOUlFOtMIFjS8vQ04MWqEhcK5VWfJUDSE0bDV5I7CG5zUbK2
6IQC7oR2ix6g+19G9SmTbuN9cyhGDttoSruPrFPhgo82Jijz2BMfs+EI+dIqq2Pk
JhdEWxudqvt+LfMXtOTLA++HyNj3Zya25hqmsZkQFzOisvwztIDx28yzya97GRuA
I63OsNzaPVZYLoYz2hVO7fjAZUM8zCRpdpEAzwwlsxnhuGajZnOh1x5hjoW9J5ES
3REWfEHXABHAFM/OnWN1do9Uc6rlSzHzcttqViAbIHUKIK5NsjZh+zjKUjgJMzqG
UeWm8K9szO5ov6PmkvZH2JXQezUHlk6634xJjz5lcPdMAwn+YL2q9kKlw4fqU4fI
PxoLfo/BEQ9s2id2o7DcmO9SMCdhefD6r7NL2Tr69wUe+mA8rkr1vzQmQSwOA49i
PZawBLKfXO3TUuU/uz9flj3pdpur7hhfJ3I65eqgJRvDwJN3D7vxoFga9/kwgum8
gbK94UOTNeLSjXyXUk7nQmhrEn2B1ZzYDwS0t1tGBmqUrnx9kkdxf7/Q0TgIGDGM
KVP8v/ID0dmHSuIABe5SDNEsUwfomnCv0G5At8ELBLW3REl9CyaWoZP+Qc4ihC5I
pHYX/TBE0q1hPdtEaJiKJ7hN3qAV2UgqUn/zacwEXKp7306HcpwRQD3HQIJNp7Vz
Osa5f97riUn0aUEILoBCLKovxGWZ3ByZp6tt3waJCMGOGbSQ4VSOZAh2mcW2CrMU
9U+j1jo6XJMyufeJwBgsH92m2/7SWNT09w2fF/C9gEIQln5lxKB+fXv8VbapPRyY
3QwYhENv/3yE06kdx57Vr0qnP3nHCHft4SP7hqwkHrb+YY4nz/v/IVs9ly1INKQu
OGQfwTKXXTMsbzu9wZV8BoLmBvgpkN6V6GLZNxKrFO2gKJL4Ej6ejQE/Zqx2/xHP
QezfQTOe5n2y9NQiskIwSTLusSg196DcsVe/2l9T6v9Lq3xQNtTUz6CAxbqqvrY/
f8HHpA/aXJBcxpMZkmZjntEUMpRM+qT1GeQBS/GAUnU9lJFjt9PkSIVKtw6AJ/QP
rtaNZXyMmQS7TLpCV8B2ptjSl7tU+UGMv761DDfCxXbpBtKrJaS3U77zy7O5KBmH
UWFIfdY66G4cG5VVSG73cTvYKPWQNRhIq1tDF8+82hB/c9EoTr9qRzBA2maV20Wi
gX4OthaoW6ifK+uA3vu5lmp5pIWcRjtE0MjVVegVVL6mop6ptzWx6SJZI5Vo6Lpe
IiEecDPlgdpLRAab/xKM8d2j6V+M9oojXuaLJ5uDwb/89ZBNzZq2peqtHbS918dw
0eEJ9wS0+R2dXYV5FI6sCCbZcDl0MA1tcvdrfZu2o8KV0TqJGzZoCqKBHq9EeYOe
nQDa9Fq3SMMvGMt/uJ+k+t84cdxZm0acodQReKnax4ydOFF0o+AGerwzw8riFpqS
DYipFq6O7Ts8F1sH1uIutvClbACYM4XPcPoIL+7hhyjGpPjz70PhsOipaeG7icUK
csmvMOec7th93LwZIeexkurE1wHKIUBWODYiMaQHQCCVjnXX/NzCKwes7SNrUl1M
3mNmXq1MeQIsRaLbEgxqizMFLtrEMPB22GgJihpJ2lY8jtv8D358deSAkselhyO9
dHkHv9UovnlM77mLgHmu5W1RMYrY5cH/q7DQ1hJXqyP9btwbenOnzZZMrcS5bzJ8
8KvBkTdU4KQtr058kx5l82pGBdlXSY1aVHFzmn76gIZVx9XEZvf2zkeNmYvdNsBw
11bid3hZ6DBnNLA0v7rTV5tO37xBxAvXrvXxBnYKRyaF2bNM0+aO9gIupZJFBdAl
XcOp46w0U90/lBIqMlnQJ6KG5Qi4Ag0F8MkCYSS9fUmqnSIu7JrWSsNPqL7iBE/O
/cdh+Uvz7eow5oQxfwGrBJVmqJhG+GaqrhRskBgZ4JCeqaQCh8mOO1BlHy7xnqJA
5ovxhv1JYuZO0XgYqgOaW7quGI2KECfHxf2aJHF0zoeu4xlygETjNDEbiMU5kqC5
op3jaOl5iyBtYF2yua12OyZWpAqEuowS6Mple7bsqvIE+eMcYyisvV/9Sa2uA05s
TrY90ZoLgu0IkTQDLeR60p9fQKhMaoMrr0CG7niI1vUOhS9pezrQqsULqa1v4jRZ
f4mK9h/bR3g8BnPn6Jr6YiHJ/9j3bZOtM4E1Hp6QtvKHRkIodi8VIXGAsum6xC2U
92cCx8+A2jS2lhS8sCV2/d/7NOrtOnXuXVlBWfL5RdfIxB1cOYCOpa/Rvo8fnuYi
+jmsq8gubZ1Qbf1qh4lU7Z0PDGSvVpIdpdPplDNs9CB/SezQH3rXFlpEn50XeCdR
HZG+EJcCo6LV8VfXi6Aoj4xL+kFwtJ0dOkJlawn81Jc9szd5aQylHywgPEKX5Bso
PGVBGLaoWIWxNz0tiPPKuqP7FKXCHFpScfJp8HDq82O4AEqqrFZBvszsQ9vRujaA
hLfG+PXn6R6bY0JY/NFe/OP5k3SDQtqOwSyJOrHjbdOtlzouYFQ62/NiwiXZQjCE
RmhO6lXRh7zax7E0DqlwIrxcUdguqmh8PTtPrT0CubMedG/fy5kublFrYxefhQGl
Hw4SbEC/qyTmNZ/WabG555cmgjYYH/ChOelQIZqeeLXuQMutpm+o7BTPYmDkD5/L
dhW78723fzZfL5fla7x15v4aVzb6IQ4i/fqc9gv2j5Yrz4c60BA7oiT2qU7bPvvn
coNwPF0E6Ku8YEoVhUl8yS2Cdj6tuSpmJotFUTox8xOllb+9qtyRC6iBF++I52b9
DxM6+BqznhUBLe/b41nio8mUxX8kQyVrOuM3KvtAS08JKt3Ne1Rq9RfVF0/uJtsx
L3qYho5wohLpjPDDjZvlwq+FSIJOhNZFkUnhBmvQkhhmO8BPvKQ82RfDJcxOjTpB
bH3pnLAQ0GnU/Rr+BqbB9M4UeurxEjK7LtfZ+CzQRA5Em4/xd5D2FqktFYBm3FFp
kxgC/R9GJygknHjeaZGRncRP+fCLgrxTf0Kaf9/+SVbJ6REq9h6zIqyb5zRA3IBC
g/TPvTHGIFhSxhvvS1yZyWh5DvWkgP7dTFlYgSGMfnSgXo8ViwU6SpMsZ9wUGQ8C
LMmN/b5RNsoZfJE+poW4o91ewY4KJY/sKmkD3lInrMOlCqgxVsZSirImdiS7V+ct
KnSkotTsga22xJPhPeAdYwPcC5F9NepSlV7vgYRX2NZ9ZXPoGQ76GWSIDMzYqLNL
lBRK2ljxZ9zakGdC2/R2tux9Tywb2Bl72MNEIOQxRiLleDnQSlnLNon41l0IDe5L
S6Zh1cIEzG+O/FtHAokjMp5YUcXDMczh4oQ7VbbhGo+P+n0eYMkyt9UxqqmJLLl9
yjA3ruHUa8/Nwv4K0t/dOmluSNehS3Y2JK9vX5x2Y10K8x3lKF2lqw1HZFkX4TXf
i4CpCGfLJHskot0PesF+5Xc+McleNCz84ErdNCzcKb4D3s93V5zJjwTvDp/EGPoA
1xVN8hetiLuEc87zveHp3fQinq8dZpw4NqTgBuyIGuCIhg3bYPK8Yzu/8H7MU4cB
/gwQ+rSzoKeuKp6vwcfn87XJyK/oW+uOiUXXTB95TBPkdNSr6JOEcNpxyCdFBB/A
+uo7Qrvzjwp+7pKk/N0RU5cfaZTuAfy6bXeMJjglefGxiUvxicCn40KFiLyavgIc
qoCaPSGPTsvZfA2YuPcCQXyJNNb9M8rKhGQ/nGIkRKoLQ5HW78hJ0MHCAYC5xzPQ
CWCaQimxZoSlmhtOh2qUFO428vAIOa17bvzcPnPygWmdL5aTfel/dIEJ0qstxHIm
3Zkq7n/lj0HNoUgbFzWLz8lZpufFw068HyPTUxxzSoT58oYe9/Idd2KHp27VwqJh
M4+NOCQj5UuWsQHJ9NjiQUIgmYM6h/9EGyc9VVX0195Tjm7Y2LXBrGwbNcSMkdKL
AhSWnV9hqSVZj9LuKRXiOYqX7xNTp3X4A3G1gyPi9dzJlVp6DJ1+9hfkgjbsth6t
A+0neM5uOcLFbeQzN84SfmKGzhsiuYkefozqKcDcjtlWs1yTQyZQ9kCOx+F6X7P7
4/7vSKFkwbt7rrt7IVzIqOJKOCA+LPe9uVFzfFMOVwU+lbc2cdFxrW2NDlYYXCZv
vwW3gROLuCAdfEEWHBtCNFr+gn9Qf7kWMmoHsO2E6+fW3HNcKfWLmMxka5abB37j
fL+kXOZtvkJnz9xkCOoRcvggbxoqabCgypt429iOc4tHGZpjvkpQnf7Kcm4Fgn4E
TfdEkOKIqYo3GnkPVbqE75JUoyKywnt+qFwXFYIp+7qHwQpMVMblLuzdm45n5NvI
6LH20WfxAinmTNq82Qg5KdlUmLbS7JVx68ltjy2cLsxDkvbJJVBceZiY4BsSS5N5
XNjdNH+d2gSOC9DKpmJVLOBVuNLzZtA8jGVa+qz5mqUsdqbrA0kLlVqO1NdCaCEo
evTNzZE9+cKYDETw4A9SjTH31OKhUh/Mmr6LcUF15bdWF0DSMTtbRKZW9Vnnt0pz
8Cx8ztYjeyTPh56Sa/1cF5qplkAXeBk47Bcxa2vXjwsS9QOO+odzEcVtvVM4Kmi7
9noW+EoVc00XOCpaHUomhSNWXtathuw2KVYOHxR5XB0ZVuQEH+PmShWj8dW+Vwu2
ERbttOdlMmhhH+rvW6eqO/nIxwh1B70/dk0xtXWhHa+xu1XZbJi9yUlM7AXOsdDj
aOssqaXl3Vw9ZbwWoseuTYZzR+IrxJl/fG+aY70bmlN/GMe0nAAso1IO2jSF+3/U
acjbvIF5Ru1IbccAIvbWQq5h8JdJ4rs/W1JMpV+8Mx5TjTnokX5Fuoj3dz0c+xPr
QagIHaxRnv766x4xHJTakXQ9yLE+9L43ImAqG5LteePiptYtCEhIP3RwjGXEufJP
9mLOTBrDV2Z+cei9SL7mMvcZbnMCMCp2j1eSYiSSpPrMvQGbYMYyoXrvLELuFJ9Z
hPNtda8iuVIvneWbbSj5IOwntNC0AAizabYtb0mHyOy+xsVhgmaemJneQNYqIU+9
7PqAlkHzkR2UWReF1yFayIIQaljxSeRpZl0Wx7SqJ6golQ1P03VwoldTiv5/fCxR
naDm2ljhId75UIBN31BPvGbGRz4qj6pxr5MvBq2Vi+i8V73Eg2UiNPIvcOk1U4lq
6Fbd/Fl7+k8U3IW+N+QLsKMavAoNYljCxH4XWGFsGmVdmzPb5wtQ6M4dCKMgR4yO
18/1qWNS1QKq2PwAohheYRv71noL4AxFJZ6ncyByVUI5WWi3qfAqxwEvv2e9Tq2T
RkQCswyX1Bx4cXZ/sMQ/8ps585hTbqTrjZHad5g1AZsyOtRKNbsRXncwAKUeiUcl
ohyYdEyGgPI7cPkqF1pvFWBeus+ln4pUu5twT+TfcXsDnprhP3j3a1ImJfS3elj/
jCy00A2JDU2F/khRrudjm1FKX3RsxCdD0r+l+9RxgyxyL0aI2J1tmX1avkT5oJfv
Hs2WZA3HrnICVADajZZnTlchlnHlWsgHUGd7Ks22dZr9QglJX5+IXjS4Tz+UZx4X
kBRhHlTTHPoIrk1xFXfpvMDNp4GKwUEeA3xmJrh5dX2Uhsl/LUgTkZfqyMcQe8SV
bnxexbKvKlNIbeooRTunNJm8aebJhg4xevL/PSeRQQ31fqMtO+ezku6ijKOd+atZ
0griPW2T+nXe6A7X38Dm8ihQdtNHkfrGca/FYPFf6+CiXLjuip5T8aM/fyoz6kYf
npqdL+RPZxMpi9+D71A8UovMSTl69p2z7E5LNq4Ury6D9+fy+6YZ20iK0er9ek2t
w6icfvhHq8T++mLMKX7+Z4GI3goKyzJECD5q78Uv6kOV2MqtiLgL7r1ORj5JFrQS
V+6jYN44v+AnslpjGs0f0XPugWWP9JVVnb6CviF5kBbb8OA4Ko0t9LvBHPtWzGn3
IFchLqSCsBrp6wM83rnSybnfA7qR1YYll8Nv6nxlJoRtrAi0R3YfXTosgELzOKtG
kPCg0iOKOOEQurBCEpPajmTLru1uKW2TERrsETUjrLwEbGRw3PcRpy6zezCtTdSS
BKF1/OhdtD+n5JS1U6qSXIV4+3MEaH8tjOr/1XAuNQEs1SLIzE6Akw4utigSF5Au
ONsuldUqaKe8r1OGKosZX4MSyMQj1ggar1bpIkqGj3DNJMQ4YgX6kwe0c5z9grY3
wRQYTp3AL7saqPoacpZw/7GPA+TXCpKRS8+61MhS6YmMkl0NFxm0b3A6aIWTm8Ze
GGxNK1D2OnYsVFa4fC54X2Reqruf4sG0uf3N6eqLZK4pXAJ4g7WCS58SIZhWg3gz
QupI1zUReZJQ7I/ZROWEk1TtJ7hO3bNQ0Nm7EEShRW7Dsdgnk1ER/VEKKVtqagoX
M5A8JRemMcEbr4zA2LL49ywqGRvr7LLUbqRUsIKZ490ujn9hfVY2HqePmOLUDofo
a9AF/cQHtUA4os5Kjv76fkVVmqCfRR5nE0Tx8fszKacq3/jHw7yqwNg50DKq4xUC
yvjZnpfETt0Ad0DXpLrqFKTtnNqcwsPmlBblp4Snt1g+w+Zx+QRPsKoVnpbT6X1J
ffAit6BUc9O1H1P8WofktpX2KIvdczUPHff29SeqpgQtkWCRgf+cVL6D9LlYpf2f
CScYYo/Myd+f26kVlhYGFHzohd1tz7O/AD0RezPKPgL3FE8o4TqSsUnhTYrK4+6v
bj2GKuQW8DZjoZqRp9HWsfPZJp+5AiHvaMnMjhYqWNEnpTDdxnYX7m2wWRjaYGAV
qncepsiATHyC2D+kCdBLoKA+OBlzkelVooi15MSYE6QUctpQzP/q7Cg7Ik5NolNG
Dz2Qzrvhb44Q2gB6Eto7aLByPilLliWy8ewXnc6SMz2LJ8ENDtuj6FzdpCzKYBK1
cP9YXho5YGEypb6LMUsC8CYP16TCLTWsBVKksMCTds7L+Sn57rtrEljfDcHm0b84
7bjl8NMmrq+7U6LBXqDv4WqjpIwCmwa5nrwPKW9YA31CmS3KJC6T5x7Ch2j9bAQK
jZBRHpkeNa06OA4reJRtROyRyBxYiSOOOp83iIot1I+YIGmlv9Vyjz/vUXb3gJaq
qUzXx2RK2PSTwLQ2zmZNH8IPLdp6CnNG6ENiK8EfGae0TPVwYjDV28YvSXs52b07
nyJVZXYbK4eNdpB1fIwWF8holyxNd5Lz3r/SQLTll0qcAcqS+8y/KtN27uzrfgq2
x91tvrXWTXYMJFhnXBb7YgDxgBoquVQ3EOwJ0PqXSWAOQJ1pz91MXopss3dbKeLE
X6rFZE2fV9GH0ofGrmV57e2Hduk+8eijCI1nC9lbmfO1vWh3GHLwIEioPe0L37dC
5b6iI4Bi6+blCv9Ml6rWmql+FvtaJsO+dQjO34nOWhxBaI8EBRbqRXoJE7LMxGXp
NYeehTfAh+Htk7HyzsU/d/Pp/Lm17FLqkuyE8MZYzcDrEvYf4gPYfBGx0BZoCadN
D+LWVSTIWW6MB0Y94vMVXDCP1LG4RDDP378rAHGM6VeSZ5BP3oX6wTbMpaRTWBCN
OxB2sge9soDSMPnHbz08i55gue8MAzgWKoYHDZSyArJ3YbUebP0FY1I8996SjJH/
plE3l2F8AInsOIDoWyS0CDv2c9dEyDcqzMPHTahY+xwWgPvEdeiliEEIkzxAz+k7
isVukho6iUTFhQhA7DDShMgxsT7CKldxKzriJ+bHa78y30T/urN3Fg7fNVEpJkj8
C3dSGzvK/Y6lderPGLGDYk8PSiopV0mG25pKr0ooSrbeJQb3V9e/nlypasx/w3m0
HzC5L7tl75dfRXNU/u/5xIa9G6juZtsx/oeEvqczaGevLRk7VopkBocbnTr88WO3
wDVd07EA2k6pZuhjxhb4FO5jfl26sOMlrXlmN8WmW+1yVI6FzZRL3ECIHLVHxyXM
RNI3i5kEL+MOF8DtsueG2NcEW5MScfs7YEf46qXWzil7zuUNw0D0alDnTUl2pfVk
f+c39xYlx0Q1CHzZi+WPVhVZ1l/MNFjCgtoGYXqTLQzCm+Z9gHwLZczAeIHSnm61
b9cyBlc5u5/jlT5tq773pvAOgpvXsVWmCfKX6E1bRBnYzhe7LifuPI4BCeUFLWYn
rqR1mXzA177+Wmm2B+siIiWH/177jD8iDtQYuMUUSygxRBjvrLQfq7F7UMnfQF49
oTBvqGJ8DCu8xL+axUcefXDYGNw9q3TwepVfJ4XDM9e9EQA8jFcmz1tferDSvH0g
QoCzp0Pu6iGHLEsxVOfcoYgxfQXhEx8wkeExQpg9EgLg/rCKKKV57vPZwYVg/6rk
UNvzDQw7nArcHefTbqliMfC8yPjGId6YqGeaax21soOkFgwmcSE6yzubUmmxi+SO
oDH8ZjeDsMa4VG60Qgli5DLwfWxLUKZZ8kecYNOWe9tJs6NaKoNVA3ufCH0gbFPu
4DwPncrBhzT3IVFK43FzduF8lan42xCWu6Mn8jHiLw94Y0j2OUp40OKETaof7hgm
keaTIPOJs7n6g/tCfZb8q/sYzbo0ufcTWTHy4qw0yaFW8+tTWInKoCIyBC8yTyWe
GGh5YQ1NnU4iqwDBTDDAJJQ1UIW+BX6hi0qnf9OFwTDSomt6RyBgZGQIzrLoKK4g
w7F1vDSDRVRccaVAmgIDFA7coA5PXU3RyVNBeFHl3TD8FClbrqdDp5DhLtsXHcDw
yr1SGIKbgx4s/n/8Wfs1kYnWTOScjUZLXyr3s2B8D2JOcql6UhwAhh8rM10u0LyU
2LzxCxPy3dRqoRGrk/8x8IEibNH29LJsBGdqBbSddwLO06PYJsq01jU41oBbGXV4
heg+PSQqyVkQmuCJOD9KqwqX3KZXHMb+oyR4yWMKXMxKM15b6mXQYeDbWGd+KdF5
FVVzW6s4qvFlnKmP/Dw/eByhtcezT2IkX7Pc4sF7S17aV8U6NkOrGliPvZRGdvc5
eTmZnUfrYVLuvlwmPhNjFXJ0nZXcWUqPwAf2eg5LwkzyVpigGMNXRI2ceHTulC0M
BXLfOR/Mo+RBeoGBJNSXq+4tw8hGseljjfc5KPCD0B0URdXxvX83FdKLu89YEtq9
6mBkQq3FwxIKbtLBrpcEG1mUDwfQvkUuhdq/bQKOWGZZAYCoOOfTrs7cnvib+AtR
/BDbcLV5Z+HAjrZnJwaSDH4Z1bEnfYTJCqtSwVIqx6x8Lmk+OB5aRMlNWI2wEbgz
QUmqQqpRqbqxmax+5u6ZNzondCKPXoL4OMXQ0wqPVpqWrTNCzXxwlg0l+5q0QhQn
cKipxWcrS7bI++wbl/5H7WkyZAnedMlotgcyLJZUNRwfBNVToyGB8CHYV0LkGoM8
PahkjMQyGi0UXnPaf4gBe+nxwGH1L8/mzrdv+u5PxrtXp0dOu7/uss8dysWulknr
WiQizd2rP6MwaoS74I3y9NDY2g4apGHlDNQEZ27D2Jkt4TrU0Iaws5tojpZnxnob
4gk8kYV705k/aw5uV58Uo6fr29NGi62EmsAI9+grQz2MNRjkNkfD7fr/XDg1ny6m
r4E1nOjgm+a+8OlOdBHzJyQestpvKb+MPhyB9Kldc3G2P3/jnyE0VNtx//VzYKZg
pQmgxm4UpE5tRFGcSw5Oe6iQi4k7VHTuT+DvkF68FMhcISz/i2VEwFJs+MYopOMM
m6S4y26Pd6qu472lQO9u1dsf8UO8vPTsHDhNDsGAWQQa1hGDYQ9DH7ClB01pQK2E
iNiDB4bmQNr4XO8x2WFC2a10FxQe6H/WKjPyz5GVbakKYotTTTod0NN2mgtBJjf2
eVZs9xx5Bc9sbJ9S7CmXSP3r7FReNvrpe9iDacWgeHeikYf3tmiQWMQMw3T5g/Dd
HfzFfQ0cHBq2UaxPpxtt8Ez1ZiG1hMbfS6c4K6wsxCqro3uiCo+1GNJfxLKvFPIK
JexHTlboW+GtTkm8SDyrBtltq6LN/EnGY3zFIpMn19mls9M9K7aKaYk4XhrQit9f
IK6x3juByPqOy1EK8d/xP6smt3a1fLsSbQPXliSnOEjoc1UTLOKghJQwhrtqiBW3
WSFVAOBIQ5p5vTwBXkiPNH+YUYDiMYjUfAksQu1MDbH5FelCvrY5iMjVpTQM8IPT
/T9XTUxNWpjgcOWVkK7NNHpHFUHotL4P2OhQ/mvLgaPzS0SiTRYVGKy2sQaHl7uq
BWFfZLeqsN55RGncNOFzSNde8TqXY9Ktrjk5Oe3RWJszxiaIYgwOC/2vAiWufsnQ
RSMmsrETig++1jkzO/4frfbxIdG7au0F0KM64MMX3BPjl5w3qHPySoJDRj1Iuqje
26dpKPL2ccZ8dREQIUz7/Fa9xvf99SrAzUQfU0sUd38gUj2IMpDitLoFq8bmEGW1
GVehCEC0y2JEQoSJzRp4oQNQsLne07KG9vJrHQv8Ty7A+kWx4776f2u7Imy3EfgP
X1dJ5bp8uyl+P2yvlYHmInYEc9Y9quU3SIKjCZlxgUQwtYCDrt6Cqv6TGfKgd5Op
FrAn+ZSuzezKDlmXsYSM6JJPLLcxdAWzSosiw/sAnQkUwUkwZL5o9cMX7OFYlzvT
RJ5Wk5iUX0/NJ9WYrssapl7IvdxAgHEzRAeC5ENvqv2WGKOlj0HvbtyYWi+tB82p
pyG9syuL7thUG0qG4cSeghzRLu56HLQLBh58LFyX/nSk+4iI17uWRL7jcoHCYNQQ
f/J9ZKkQg2VToJ4aHYpb7pgrNhBOvkTQz3qw9UnF84CZWE2QqBejjI2uLhdp9aJs
Cmod0doI92YlCuhiRcouA+0RDKIRQDuwsPM6OPlZW2VU0jY2+3fyEqrfMCyVXNLC
RfUAAmCGMJhsi2yrH8GHkmhCDYTy0E/sh6GHx9Qgt9xFTSu3KWX2tBsj8glsh1o3
jvzLNYVwANYHSRcivswDhcq662Ln1K9aHRFpvcFdhiU4rcOJV4hpr8BK3YzNtLGE
PRsjxB+mWSi1gQSPLpQCYWJr1q0gfhUYkZBJVDc5a24A6PIehaMoyIISEYNsLkm9
1mRM6MXTIzxzKeLj0078sFd5Le5ZVg2J2raobZVGQQmVpdOMr4lCwUXLiI/QlXtX
aMtwm5hZZgbF5cb8k+niLqy3/oedQtTllI3QCPh7q4XUpltyqcYuRwT7rWzWrzVX
4BlJuwI0BqEx7EOTimv7p+YKExuXATu6XIXFoV4If4fhtKhCCKDwexjgSRbaa1Tv
gaBiM6CirVhbBW/v1MCLn7ehQ7/C5a1l3M5+TRHo1fXdFxrj+VgPgsXGVZDgrvYo
VlfoaPojzZQcHPNBdU1YSaf+1TP105n98U+w5RQMIzizKfnUqmvsJC5hMY4JZiep
w667v13hvvOV0ScG6OaZsasnHFM+LUzi/wWw95cBy1/fotHNa5UvdDLZ+zihCFm9
QIca1RvK/q5HP+EnAxKjKwoKaN3koZgrnhC/IbAgnv/T995Xo3JYyLNwbMkY6lhv
vAorWOa0Yn2+I23A2gsyaTSZ7U6Fx15VmjTkU3+hxvfwDCY5KdWiJIYO8m1dAF7e
feZyAVUejvcALE5slpdWLF27b5qFcITtH8M9+kFiL5Pm5E8PjtVrVTGwFEb9xaTw
2zb2DzxSTetUUYSHCHCMgG/R9Abp1QTBjZPXjwlQ7cQbjreoBZJpnu6Wq877roxc
GMKZTqkUxKj3X7xOv6TwttnuGmKJHaCdCY6RhOxbgnHPBVCkI5YiLuActn1EjlfO
YmJHS/Pwh96wUVNDjQf5qqq538mzWYy9890wMboT2wH2ZLljMp3Aow/dA+oTZLS4
5f8nTpQnT5HaFKqJNUeO6KH9+b4+dRaW4jz57A7j2kaJriRs7KW0LFtVug8+XNb8
ROJ1Y5Xu0g4iYGesDzkwkLsv6FQYmKQ58xPv8g2OsuY70ygAX+k8NPTcTny7/ygm
eiR9+NBaAFuusXI9gsTxYTDo6DhK1B0wpCj2yswI8LGXqazOTgIH9xsW2jA8AWZE
xP51rMDkDLWbcuu8AHian5CRjt7y3+C+Kt2n3Y3ojyOUs9zPHhkCQwN8UpLS27oc
F/wscejGyTlxkE0mOXTLYUNBTt9tHoh0zd9zfiEPNX6IDSIgwOUuJNHfvPucuTwz
hPftkfMm28pr/e1gfQZ6HAeMEFUDAJsWHXasivMMrMGfjMDp4HUTye+vQsTTuj+H
qhY2HeC4ls0eyLQq2RevZM6kMQ9Pi/vCzsuBt8E81aNIIPwN9K5D95NCKEyKHY48
AcEqVA3E6SiWh8uL9rv9HoeYDYyX8syL2YZO2pUxaThl5sd5QVTZA5ogyqz6tNLi
omWz3dIRW2x3EdFP+ffm77E3/ezhfuCIDWVtIsQ5+3nBjkYa1hJk2gnN0XC/cQcR
9szcOhQs/739evLsSqKQVHTeDN6VObJrxa22nLIq6GvmhIGYh1h2hE9cnXataG9Z
Hp8hTrmSl7K18+5e3l3Jfsu6uO3zQrLae1wafrxkYH3graGWvBbItkE6hj+p62Pk
/bnm1apU5eS5AlEoRFwm0rqoY9NjC7PuZ/193mzIXWAHqUri+L5uL2JKVNSccc0e
I9G3rNxmpnta3aFU+OgS0dMqYqK9qojAAXFRE5c6X8qZdh4zDinIdqxtU+YhUtmI
Zadv7jd/baU5FXYvQejTYKWOCFTPUDfLDC9c29Q99z4mKmrTGGiQ/8+Nl3/zGA6u
HGrsew81umBzAIbourIcqi7B9nKHiEoAQ5kBlPFynQiiIMXExGt7rb1NQ4bk5Cqm
29dhDJTAs7kTgUiFRoUyW02oEGbJW50woQAZsUxYHbaAC1B7bibHmJeRy/P/LRIJ
NKLiGa/8DXoPeQr3Br8mLJcVkQvPT+WQsc3YwsXrPpJEVMNRTt9bRLQXYOdx0JQx
yPLL3DFfilWzMpW/J7fbWl/yiJn/jyrxjnD15SgnI3tXt4bx+U6TfWD8755viajO
D/BWa6eFjjWG6qtWaI/zNWY4SZvNAYStz3Ch254fsScpoA2L3cTDbu4dJnTS5101
CkDHRqlXNbFSsVqfTcULazPXcfgc/WE0oBkPCXIzg/czqso0WcQjbKCMGjXIFPEj
T9kQvTYO9FPzrNPEvUMdeUKJ0ZuL5xl/WJIwOf7U0cHqjeOF+01qQm8A1VtXELPn
aAMYru/sD2jg2LYe3ljutqB0YkQ+Ku0o3F9SovIRoRWKEtpHIR1eO7aLRDvgYL5B
ieMEgRrsm2aK/d1Pbq4Nx28b7rMmb37hBhP9rZyVNHjatzWnXr58P915JexKW924
sSex5S8mYr9adgcHphSHHUhGcBanOxVRUYLiRYwy/hak7TQkKK0ISuZ8QwSBpmIW
X7q/WMhsLFCNisdo4xvo6cadopcR5YdmMnWtsETYaNaxWaQFumfvVVGtDIsEgbw/
QXAm64dg/VqvsFFBVui2WJLeC5WRU1PjfQXf0ZZ7+XIuUrnonG85H8eD3K0067MV
e3uFaUw34Qdb7rzoaZuYrHahwhntqfQwwKPUQN5+xf7AboEwUjeyC+vPUiIknzMq
lgi8gLyiwC7iC5ATU+fWuIHmYldIzrMlMH921mkAyX8OXw9RDTHgvp3qEtaMFwxT
TaN5qahJy+shHZm17qfk+Y2eedWSUoJ1hyvH1btUSKgsNLvfwwVteNtXVhwANNVI
VGiyu8eadgU6/OEDOzfKhyeV9JTmMBYOjEPZpk+GF7di3e0m5I5se2xKkSfdzwpG
wzvJPPOlRA4IIKuj0L9b87Vrd3SpkU2Ocvr0TtSo+5EGkMOkus3qTNCFpBI/pdQJ
uLeMozAMO1CpR4z2LTatBFrw6AqV1aLPXi3oldKjvEWQE70lUfvt3ZuKjZGXcW82
GNIWzvRI/Wn9ub/t0GutO/Gf+zXcoyndENek2IwZkGuuYBN+XwdtDqLC5qSXub9M
UmzW1cWNtxEDFKDwEBJNXANMIz9Opc3d/8Dfk0EkebTqrdAuwqoSHBy73A5okgS0
Bhe0JUW58THGbSKBNhJ9XOlix/iFrbwp4ITtgfI6lm35yidvPQeu203yybS4a7Wj
qZ2U5aixgKALgirRxqdl7424yUIHzpSBlCt9RKqqVQvuZq06mL4F9nU9dudTyu1e
bfS40TD7bN9ly3NehKZcaQH23V2hsBwISM0FE/rrVTeYu/o9RWfGqRXEqz/JN2j1
siPq8W/iENV4vBULef3kizqQryj6g3DssSn3V+By9fn4hMwTPQUemWYc1shYBvyM
25ftcq4Z1VBLxyKWMxBdSaUXvfMP84RmTWzuc5luvIRnbqVVKsy/wkbyRqsGiee5
Vo03c3bzZ+69dX2WaIwddIJHMfuWVXfJXd/I2+uhyF63xmATOgV8OnjO3h5yH4Iq
CXla8m7LsEXbsKEivMj4kP0rDUhICNeEz7in8DvepJwSnUmGJxrRoZDwYgv91Mbx
FDw6pADeghMYalMWwagC/LtykTP4UUTfXp0nI/QMLTO6SO2K6n3Srh+wMwl0/4Oq
CDph9yYm81WYyffkKjN/xCbTuZH2LX6zvXBirHacw4C+DVnKRFua+RuFWYDnWPtM
0vNXwGgoQ1sp/39pOhSclGsI/FlUwZz9w0jdTI+BOfLOEsUIGPiwrs3BxYc1VF2O
baJqyYsyNs0BIOyas7ZeZ9EfJdLyvb+HKgrUDZ7t30MARzcrljIp7xiI2Qk4IzbH
dOZqrJmmcy8vrfDuwYi5ZI/tNEmQPIyfLmRdzYkaL8wxOftGdmnx8yRwCwaVYhTr
lB5mFRi5FOpdNcVhtAl3+IWfbZ9YZyrslN4xbPEVUmcip7qbHd3i+LZsyGk8VZGH
g9Gaof+2YbN+QzOSmTMEJdZpikL+PjzZG/Kw6i3lH00I+I1WyFuE0OJoU1BOy5t9
/EgUeNTi10UU7OcEMhNuo+1SXHg3gdrtGk0SCGwDpzwOWdQ7JsZq/eO0m+IgJ+B8
TiV6fs4YLijmcWH9zMeRcRedZCLx7KKocG7oOSdE5hqwRvH0EzfD97rv2LqkyTvA
sUW/LVU2N/ePRAr5PapfaH3bO8KtfSe4PeRdFuccDhympGLpJU2WbF6rVDwWctzq
1XVfTvkw9689q9dCtObkaHj4Bjf9fSixokRHLretvY+uN53J0MrNDRS2BU5w2GGH
wvUcuH9HXJkhM/BvY2k7UYO8AgiJO6XoFRibG9rXIkU4wHuXHOwKcm9/Ar1F6fT5
Jn4qDvppwAOdbgSg63BnsjybB1GrsZZSrAtwg65bBcMQNLAsq6naxMp1lgE8Sd86
BMiRCro9Ew31pF9mOQUGURvn9JJ9kgXWxBZMhw7tMEl/rGMHlLM9NVyA1eYqX8kn
9ZtpL+AFUURU3bHCL9DC3mVdbTKvaVv+D9H39ilr+lxa3QtmulJPWzAtVSxeQrdX
aIjJVaA/5fkqqNCrq45w8+LyE13eix+bAqf2ZPInLayh3sdGgdWWd87T7mfO5nPR
2PqpbMeWPu1uC/cgMUSnLJq9DKq1w8tj+ss7x/lM7HCcp+FdJX69K/cmdfPQ964g
ZyVO4xd9ZO9wlrsWfyMFBcf6zuqb3nK3Q4yPpaOniybgBcH9W2gOA++gFhRYKdDP
Cb1eftzzc/wHHPVANU5uhyQPh9P8W9C9LMc+vNyTY0lwTeR/c7a9if7rRFP/74zQ
440qpGY3sTa7NDBSqRtp6WJCLX2M21RVb3uzFN1ArL2g9JxWue9p2tf3AVLIn3RY
bvzpjERPOE4t9MRFzPykKGSIQdG1eNspgAPrGIL1TPvGvINfVHlDJuPzmgBECpbQ
iv0UJCdO0S1T2FhPl9jjRRfTjx64YXqV1sqoNneTH4jIgyuloIts5sVioejoYnP0
IPA2RkOijUln4lWV88QBhxl0SgceZMMtOfVOjG8K56V9LXSeiYyMkYJPIleWIA3y
kEAUM5FuSuUI5WBlQw+Uvz2Uv17nrMroNQwhAFNCWeLknYvB5WaaMh21MP94k0yo
X2Lu/IhW22Po6nXuHSVO5QkJe4KNpRkb+q+HmjbUuwHJD6ARfXaLY+msm4mgsUZI
rPmjlnFx11Tu0YGfBVC9W2Ku/PbqWIHq0K69jJ3ei9WlcPHynXPANqhmKHHiitKJ
EXZmFjbMDwGUqNRTJyYk914wQPFd+0XhtSjdSg8WG4u2K39lAPGvDyA73Sk/WV5l
bbmBvSevFvXumELlheaRzy6cfbiyEM+65LFMDxomnNlBqMUyFUXpvOwE0xm0nbyi
Bq+m7KQqbnaB5CKIv8futdRAKQHrmSVJWoFQ2LQXAGJznZSakdSRMw7Cn4T9gxBC
fyrSSFslPlXTu0rZKYTWgyU05A0iExsGaX9zuJfSGyUJ8p6uyNhsGIQq9ar6Lba1
BRz4OPwdbRhlYFk6jU62e/Xm/Tdd3iMphv2PvEAH+R6M5ozq+0GrPilPa9IXDnL/
zPUhKI9CyT0KBdHxOE4gF/h+X5nbgBCNuFellWyPd3mqxPLT6vDYem3hevySqh32
sdV8vI5gcr0pjboIcieKec7xIPHh8mvjwSmh+yDO3N4Drxbv8aEifpIqqoLvxz+w
tfpnmwHaPRfchtPczKppyl9uKkuOReVjurWEm6PdMxIXeo3hsmI8uGPoNMsK7nE5
7o+DkIqFeWCn7765/JBIsJd7eCiI8ZDEI31xChsmrHvv7qb7v1PeGGhssE4PsJyj
Y6rIxucorDwcgFPk4FEZh/q2tBcldrZ61EFtXKKnKumOhvZAgNdz7wDuIYEP1Wrp
NCnA7PcQhCLxJa6zs3zA2xuVzyJxQJr9VcX6p6qTtpgDT/IPNJMdReOKLEKvDnd2
4NT8Z4e7SsD/TkqHlWmBklb7QY0sf9y/gsb8hNrNVYHrnyVd8pBmzAt94k6xSt7n
b9p/Vn3V740l1hKLnh8LGbxxwrFABTeV6oSTOXfLcvMmgeh1VFwy4pg1py+OCHo4
zMGjXUar+hiBCD/8pPb9byLbPp99T5QAv+KHMJuFsP1GM4EwttdaQFdEfXKm38d2
B9BG2jUu6pt6p0ASiTvNvK5TYNDfo9mDAbAT6KPO2x8rmaYWJlPfLTiBuGrvy68L
E+fjZPXEeSn/Gsf39mxM4g26QLfcByv/7s6UKoDe6r8NqSGUwzCWjbrWsl9bZqCa
4lp1im56XSQSn8xviWJpPMoCbxdv7fW0fIKDsxFu7Gs0bb2miFxcKlrKUi9YcLnM
r0A0MASzbSh45QLUT10/FXXdvCPe9hR8yp29oCBK0Aw85xJU4t+Q7v0OLA5dubD3
kIn3JsbWYtOzfJ8oYVXIJlb7ZM7Xs2ldmmUXo3Ifpjf5EAucZB7osZmUe5g4y6i5
WABnckwSC5w9EKhYqpOZ5b2pjJFAhG7F/JME/J8bWI/Wt9+LHwZm+22uNBNkTfOu
NqrHR+OLbWFjSQ5u/+trq4AYSOFUJNMlitvu+A1KLTKJZwkqTm4+gbHZ8Svie2aK
Js1wdnkABKJSLrVPWOIXtJaY7m9kdEdPjqkKOssd23mW6wUTIwikuXrGxemlf1dL
7C6Lj97MBN0C192/WjvajHZSQVcINfu1CyIvIC2xmVpbR8cL1Jeb16uC3jhDH9eY
nYfRoRD6NGMMNqMs3b8N2mENz04a994pcHg22xf59MWeT003VZxQM0Lo/GUoSiIu
ciQydOveeaVw2EsmAzPkRUrpBtW4//7HCotwhaVGF65j8PwJdH7QSx3C0EaM9xje
r+Vm7I9yZVadIaHVpY9j/MZGvxjP7VeOHTKpjhlHqL5EEuwgJfF1/r9YRnqZj0cf
EBZUjB7C3PtLJTu4fGOY4gu4AQZK2F4bGKTKsu77vi8e4unfQxZ2B2B20uwioS3K
JnLls8eLeIm+bmZUvZfP3mI09DwFnAh+R2wSRrIkci471uKkvcvoijUdINehT3W5
7c1pq3CcSqrAG5kKLqjNXm4CFCC9CzEsbiiaPj/A+9TD4e8iOSMmxO336SScRSbD
99w67FVqr82HDOesuw4lYiP+2c8WzGHgyPhEvdeL2d9RKBUfvsiZIG5gtnJl0tPc
imEp/cqJjo13ROOU1/Q4ywh1MfLZmF5eDBNNovlDtOY1294+jUPKoRicdXXJNGun
T1VtQsTJ6QYOy49QZnOLlPP4/vNkau0APadrSYWMJcw52ug/d+NXRAmV2llOnwFZ
zDDsGLlVbTR0+NV7SeuE3X1RqYX/S4+ivPpBPi5Jg+xCpLGFN1CNHf1n3Sq4qtrW
mU1gv1IRMqJlVSkbK/e25tMJVLqBa2PlC8UNmOu1wB93s1C+7jdTUUnsIBD0RSx4
jCCfmu/VPgdOUo9tGE4q6Y7tsNX0xR9BiLI5NXaSd4Wq+ne/k7y7VKyl+QWuAePm
HrS/i++puRyYmqmmZNHHLSTT336YdaOtqRMstVD5SFmS/TP01QaPNAtn6AkU/ADa
LTLJmmpTZ7orKJ8z0JxnfqqSJU7rY3jyZlln2plAcZJZ4oVwoL2eb2Lpv4gZbLbI
6IRemkSPJtYX5hC2aDgT878A+ju0IeUYASgtdCD8o9IF4GMwnn43QXlTdI7808yE
MVJxs9jDr5uUzoYW7VT98bI/jiKhffkduGLzCpncnjtYZStxSL9ls5e+IBL2IP5w
XaocgMiyzgacqrn+5icjzbQ1rENKsWqVHJtgAzz6Q0rNDMpNjszZ8ajGgoI/MW+M
p2JSQMSg73iIL4AtnnFRc8jyC/pt0cgc61Vls9JmYDsi6uzS+kJJ3fleDV8TeHVg
8Q9LXvRvLiR/UJfnskF6yzyKEZ01zPGVYFh7P2K0+g7/ePggiTOUJUowBQvZoJ7Y
hl3S8kXEtt14nzsY1C5W0GwAHDxMQxW90YjfmBhkEq4R89XvbqEDthSzpvk7D3XU
Y9VI0XIeA6GRzl9V1nKopOisKGzlg8CppNVtI04uCuyltibcRCkAQWR54kcGnDlB
bZPK3j+nt0r5hQsMjoblU3uT7isFW+73VGEGJWL8yS4v4RQavgt7fnFxkHxiJqVP
QHL2LNFWTDepQH1vB72QaRnkLc1qcT4o9/5NsVkoTBbN7uwlgPwp71pIafNm8Dyw
2F1ZYdR+y3bHR7PEuBEyOHNH75sQf09XZErfsm4h2URI9cusD2+dOskLDSCfh99C
W6yQwpDVkDExbwJQdsi2B/TRbvtNTID1KMKsL0rDImQgIWvYrcJUlbeZYt0rpjGh
3CBLiUPrHcd6fTtGBcdR6MVsy+V83Ymszz/9DB6hm8AEoJhY1y769sD/2xeHL79Y
vpW1nLni0Ii5+fVCNQRTal/mXK5Oy24YA0FKKD3JkRjkcWGpnmOAbs8tJ30VCzbJ
7Mcc/Ct0ocJVXssIExT6s0vb+lhDuOpybBTst7m7dHTzZ0Uu0M1wvG7rKC1Cm5mM
lpi6B+Fmjj5dPlpkKzrKUULEXqv6hmARenyx470s5B6lr6OuMRlaZdnwgl+W4ZFi
1kyd1ImMiyKCufdIR+R2e9NOC8GA1NX0GmeaGYdoEETG0ElLUfnoW7Lfa6UDfeYE
jawD3pwxjM55Vndc+twHomVVdi6xsny4LVzIJ+uFDPFEhQGIDEhX6ak0Ta1V49Qv
FYVyXbsmU8GUWmHSjcfCcS+ltohregwrPK8kIn82KkIZPYYOYYV3k1Vmu0h+nBp9
Sbfm+aodCWzUa1Kt9RuO3jDZet35KhAydolaJEAytT5PeY3ghGwyS7FN6UtMCFQr
mnuG57yZtwYFpK4cd03P6aImuxzvGAqrXKXDgba4XExSLw+ZpCx3n/3l9yQHgOvY
POmgdx2KWdpCDYNmWINEVoHQlf8ylww7/z8jMLEwBJK/1eR4FjB/8b+5bqUgAr8g
Z0QveAzy4EyS00ojiWdWUARi87g+MJ/V3EWfz4kJZCaxTGWcvZyxql+SvjRsyymD
87PANqbVxz8SCiQSsHZjN+AyxM3LyvFe2q0v4SKetvDS3ZiVXtYMGoKQkc2mtXER
XnPZo0Z+cUZaDndS30WSmoKl5zSo8ICB+mpFwB2cDawnrxaAhB9pxCuD92bBUWzV
lwYpkdMq7AfNuSPODAenblghaDNfXH3H9V61v8zC8GDXt48SUaM5df9bMTC69kf6
8dYqKhsRkCp06DiObptgreMoWjJnRKw6we4I6T+3ShyHhPHIXM/4h9UYCfoCNGW1
Rh+SPzftdw7Nt7f9cS3R+qdN3IcJgLen0xJsWNP3ov+Gle6eJyrGMLSKO/rtu8++
+VWhYk6orsegRAXXJ424G/mPLbSngs9EICpZEap0z1Qvv/pabW0uGbEaV7Ea6jSk
hTCY1Ar1N8Ok8PVHG8G4NSpJseuQEDRY6Ga2xu6qv/XIzhWON+YR9kzljeTOn8ym
4mSzbe2D+ar3Z8SROQPW9hhibfRJlu7RA8xMiQ0MHA+i+XkyJzhbhc+AE1zUL+lL
j4+Eb0wnZSx2R2fDaX8vBB8SkmkIlkwQ2EJnS4VS9G1le+zl6+7uuRAU8CsghHA+
MXkBCDCfV9XbW/a0ZCMVBk+6ctJCDhNyR7+LLKdzKz4JeN/XCxpTM9ZfS4kW3cRg
GZLmeM3OATebhmFVlvBU93d9U4pwTX+HWwWJV+FIh8gV+lnqOW8shJlanRIEwE0A
Psa6apTPDQGRC7wkxQdDjWrzkj7DsmYhF0C2rx275f8p9r38gsufxz+Mh31d2S44
7wP8ztI9TpUKQp3KRa+Xtf3jQm5fpgpm6eS7q7COEGC4pxeMExDLVuKnVDFmxLu4
C/2HKJJR+YEUGJUXAl6dlRv6sdF9EXWMM1xAG+INtzGvB9axuPEDpmS7kqsGPxRR
2cd/u96FDGhuQaFtA3KFRPJZJlECnifUPeM9m3M40ZbUw2bhS+zNW2YftRMfpRTe
OoV2EY5pH0dWnWoQhbM6X/RJ9DXdTywNcEKRDtKh/JjMiP+1/9N8UbN/fSI3MokO
+bDEBMJImM8+t5Mc6kLL3vAfKjlzd/WPeD77G2tulMFBe1vff0bS6Hl5K24C59Ez
08Wk6MVdmYDWqVJ1/iMEAmfWYXfuk+g4xan0xBHIzs+D2E2VOevwlCIWp6Rarwiq
Y2GZkk3i3lqTMGnol1IgepZEVko9Ra8Q7b9gozG0qnpmNbCUy5yloqv9ft+elXsn
6FY7YM0bY2g4DzLPz5Og266EmSOFVFVPGiUDeAHx3t6T5jaXcDMWWphv3Xvf0eWH
K/Uqcl3Ts1opnXompv/S3LFvZvBgy5hUT/cw+uT+QGI/y8THlEn+D1UAdMNs0bqa
SBp48nFhXeK8mSGhgr5uyFzyuYILkMPeLBO6HnatY/jmA3O2ukWnTU2Wgxo8jtM/
CKf7z938F2HGaRtT4o/QPsYTShanRKHDVDsLMStMFTpFHt1JCCYLhohDPhLYCxth
hkXrggzlNoiU8tc2kh/ntW/oLtfJgwvTQOnSIZYRgwIE5ivq9HcjMin67knhIoNd
Q1gvHzATlZEpxnjBpYByWO8i1WniRoJ08CDdlwWZWP3fv+5pDMqO25X6rkAt8xgR
HHBCIM8hZ/9dpYWpZv0wAnUZBf9rhCQf319P2OSyZYvWeto/q+K5yiAz9o9X8AZ6
VoCUvoM3TTvaZ/FtZ4arjfa/xhVwxSYo4ctAdc+cZcrl/gNkC04UUfy49aQqNBLU
EkBXpQKWa4SMzlwuF8zENsa7WnYyJlsZa6X5zyrH0pheXbjJnaoUtz2KVzc4FL90
wOh6SmF3dUi0LGcMVDMN7X+3duMLwNBWaVfiX2iPFHn7I6HpIMMj5+kwvExIteUF
4rpBMNaDXutLOpXRvtZnxCFyXA/Hbq/9kALxd0+bCjYZ8XlMEUfb5feldfPYYQo5
2ud7erZvC/MARQjMZjUnjGcAFmFdC8K2erxovfGvkWaw5obavH3xBPGKxylR+6O2
QYdyrFJ3jjJbg/A4/sCnjY7eYvxsKFgmcnZ/rek5XxQ93LWlzG865SKSNPNq5q1i
JVXZAt/yBNTePdhE/ijK/V727uJFupOjxzbDSEpXXgblkcakA1rej2KfLYXwq8r1
jNtPEGx32kj10eSvJwg9Y+6RnROA4Hgrpvyt63PYtKpWTkvno30vJ4kXz2+2+P1I
fmKrCI0w7BvNYqFschOcFHZH3XmMgYM1Azfx7WJj/LHiQVUtAQgwSYHHdCz7+ZUi
/4xOfMF0U0JjPXnOyJ7+t/TO2m9jukbjLocKy4NJV0ecjAwNQchdfAVDGFduJe6s
+WqogmuyCEL6tqb5jn1QYchHIYkTam0nofXUc289TVJl6XetdbMi04NMvldjWncr
D17iYpWj9ZabJzPLKlhiC7Mma9a6mA245ptMg3JPO8KtFP6nqz3pQfI+V9NWFAwI
DbaD5zzQH52/c/89ULsmrA5lxU7+GRcT7rVlYH1pKCA06sTSUWI2x/Wsh1TyEDWn
AepJ7EEjyAAx5KBT6fWO4FgBaRPl9vSQQ14/pl7sHXHeFd/VgRKosvTZxECYRqOG
BjYjqjU+jstBrqQR7uhB1doVEJy1R1mG3U7TJjzsYGDVklJy4T9cODH2qSkTCFNg
DF7KNyRIw5zbOtSzy82hALLAIqBCmW6R06hMMuKKp0F0YkG4eiOuYNty+zBWq3MM
5xskuLJplhhVPLZ86CvVivtJDFUvIGy6ozl8ZTysreh09g1F8yNmQHuLXNAbaTnZ
7H6QaJX3xgWbSSwdRVoEAr2+S8E9smK3hlyklCVEzI+N5pzqWHlnbIXxINK2Fn+p
kM043cm+B+LvOLVtRX6c+/+PqOepKwu2k7dZwPkKjRAM+TGsyxfyBhgqkDu15m5G
wq8f91bqq25SQJjVziScUMoHvlNhE6zTDf6LcUaLVvTHTSNRsu7VefIczdhbWOvn
PwSTw0Soa/MqItPk5/IhwpuwoJvwdGXhSlvezStt7MTKi+XRnZ2uLgmWEvUklWtd
p0F+4eNAn+cgkU9kFq7lTQo5NUgfI8TOcxss06tdoiNaaEUATqjAvQlVc+cE8uHw
IUoKZtwtusjV6Mz+/2IjBZWBfs7tGsFhXhsNPe8s9+5mugoRyQ3NeW39BcKPJTlR
nMwmPRXkqNMUSdj6GUv2geMg0G7br2FnAeG/jN3DVSNoL/3e5AnIaZpr5ZCOsXqQ
RpXRBelMuoD9Ov/3RYhmly2DIQDdP8rjyAvdpno8jeoP5NN3ip4h7Se7LewaKMaL
ewJgZ1NWU7ww8Edy+M0IeArScTaK3Ij0RmZ3hXDZoDmsFp6izRcczWMctISzdPJh
H9dMc2i3A9Wpf0gTdh8jgSA7tKXQmNDIyfFoWNhrBGI1b7rHyJyqp8GRWB+ulghB
BrN3M9uWKylTiiAOTMxmZ1e1mFxMdPPgt4yKHxNIE5IB95wt4qVatLCU8L1RLGV6
oSmjKmtk1wLgCw7WFTr+8JKpUHYkRY9JnnGq95B31Z6ouKwprntviRGfqfEvLsrs
auFklbs980cMgkzXfzhO+drIcgNyY/ExuCdXSgzyFpfatyoK95PoGP42e5yYzEL0
8UfKFBQURoneomvAgpuXHfJoyPELA0RMMUuLRtUkIWBuhNofoL+diJgxuX6/L2VP
VLE6Q6B3E+ERarmunTZE7DWsPzTWk1QuCYcYnsw7CLL64FThPlbnEtq4Q6/HXCax
lxK5UM0fk5Sm7Bsbt3xtFYLZCSg9kAQjuQKZomxUYad/CVYkuSw95DYqV+kOvqg8
xoU9r/wLD8FpdLkkFxe2UJ6lbCVPIxqYgbgYWva13LqRu73l5hNjMqhgjbHy1ko2
8RRiRVP6HwrKEm9dTiDFTu9f9KuEtqMfTZ+ixxTshK+bh4647pxalG1qZmbtc8iP
Rbwry4EC1lpfw51j7v7KZLp9tJCza1XzAxSosOQ0+WOHh9fANmTF6QZxYswxZ23k
r33psuOTYDcbzFymB7N8U47hlB+qktt6H1sRo0gk0LH24jsIQhotNFslkMxklx8w
wWHQ16rbpsQoHKOwbe6007y6EWWrwxKd0+BL9oAfr6SMRtCd17hn+kBCxgd4Q2Hl
y0wlEBZR8jTvAokc1VvgdSoHN7kok+gUBWEYqkqZvmJchSJ2NFohHq1GO6LswbCX
vtyWNMaTo8dFssA7kMPhlXmNIDF3LNJWcTXMktdAjAhde0tzJiXSnjQkKC8pzcpm
iHexTCNtUf6fwNGcfZaZwjG6Vv7YgIaVlFSb1qMRZp4I7kNA4zMY766Z0KuNxpiR
wFQnkq3QCTfrFMzGzjsuOLaJKUhPmf93KlS5C9L61+Su7KIwpnYCRhqT4Pls9CV/
ycbEDo3m0F0HBban8CxSHjejRWTM9ZUwJWo4taypfq6FtjB8bLGFMOeKFXnQAacX
xlwziJMj7JaLAqWj61h0O/WbZZB0guXKHLJc7g3aiDNJmsV083ipNkpMiGnwNmU2
tWuZhpG4/BHKhUzr5elrSsXWd96qhbs5IsgwHI+olmu9ZEGO0YAcaVf/mdU/swQD
I6RytHXOuVCpAO3PxFqZ7WuKPwe4p/4sW/sYxKy4BmjbC+Z5TX1S1w8aGdVJVIpK
IxLTtG809wY19BLtHg3OM/P8zz2Vb5+cvnPmDWhQqCHIiIRS9sYBGf3S2cFzuQ+e
CysFnpyyrlnQ2Rqk1s9tIhJSI8AlolV1EwGKm88CKeJtA4XgFm402BwgmSPALUSX
ymS77phxOcHxrSG9WWHbDOTf3qbysID7zoR12PWEqNgosJlnz7jHkRAIxpOpLzof
waxMxnOBWApiuVjkgXR7tVDY/j4Fg6JLtotY/8ebgpz9mx20bjspSw6PsG76uGJa
0pO+AuyvMXOZhfZ4t68FGJXTS0XRTKc7povEHCND44cuq95itefL2vchgK2PvtQm
YPG7Q3M7XdbIi/0e/SrFJDZfZAAycSE1ruZDCPel10Q6+RZJ5K9mw+6eTp3UX8fP
mV2xcKoR0XqbMxN7r4TGRDh4Ln5b+yHEtBboe6TuAE72nlBDsjjJwY8Maenufsrc
jBrTCQY7L/p8ULfRCpGUSchlp4hn3jX8KX9e0tx7m0mpp1dt8zmo8xFQFAVfRLEr
OH228UkL/nolqocUF9mAiKHpSLBBaQLK+l5GDdo9JKQIwGFn2cDKjQ+k+XNwYBuz
5X4Fc9x1LC6rS5qrXnvwLFq9p9yCNb0cMAewsBha6Mhl5RBDSTy2OQkyUGTMNdMJ
qMekj2tb06xIDTmjjsIQ2xUGcsiCZdI0fRi2ShHJ/0W3eNmayA3zm3eiYwiKXkv7
av5XceRVbOOcEE8hEyRKYVuwhdXlRrPeu/Yqul0PHRoIaRguQu1y/qJFZFezsNVg
aZT7S4mjYW12bv3dzT7Z3qJSnTDmGhk9C1vjWeYaYp4FR8K65LNeO/0IukbhZ2sn
AAH0QSp2lVkpAiQtZTdZFLfxISJX9KAGdltPv1HOQQer5nWxrAkOkh9lp5IcgvVK
pH+jmG6ESNXOf+XdMisLF0qYlg0q0MbikHTBHVQiT04p2283Bix5qhkM72PTfBlA
lkhjgyiOcQVfqw73oKRHrMFUWgRnc2wmmnyVNRkgC7Mk9TKPCYF6DRHH1gCv0BcU
/1lfq1L3teTX8Fen2cQoy3cjzfbPeVj99kca6TjrEhblWTqoYZUzZuwhNiD8QG8O
Ow9tjBUzXYbdK+JpUFazgBsd4VoZ9Yvw8iMX7Ojim6i4i24ID/0XCuhpPV+IiNCi
uGHDWmK/79oqeGl6XMB9d1q0MyZrxE4DcmnfoqRxIQtzCQThkuIE/FcP8Y4lnsxL
RWds4JEH50+PYEqao8DNxlGnwuxzWdz7BaAdQy/WSWMmusCTRTLVlGgcUv9n7OS5
UG8InUNN5CYF0rHbByGF7kJlhbRYjqtS3a34xxfGnTYCyc24HHA4ETbR6LgMAa7p
HOkUYJGyI4tml1bi3M5Lc7lHLxbt0jeGvniB/YIliCXzPUlErjgFuk9om1mapVI7
ubiohSEo7qwYfCFfXfYHdm3t53sC7V94kWSFmUvsZRv49wPg7wblVgSGbGCg2AJ1
yqARoD4fSvmqNSyhmwzObVpwKckBPdjFQk0mt7R+90GPaSCet5PgxD2XKnL5RJvF
y7qzQnhtaGVLvxTOvQmQSijBToV5iqjfSR2fWPC89/sTJbt1U4MzyFpimbAQS4GR
NuumbFNM+zp8GN1uEBdLExLAS2xplEP4Y3rTQKuViIW9eSga8PQKJXLmhU3FMZLM
l3iRuFkcoM7sPb0wVNqu4EYkrKSrXDWW9ziPWwcTJOWxvqal7+GXW0WEv+CDK2hM
/qNo68BvZhr2aiZaOkLObykwVBifhh9gwEBXdWYHcgwB/Br8vMMwvSxm0kXHE2Fm
nFKO/fu40wGnE4x3tDEhfq+vSgLmR1fJtV4jiY1Ir8IVC5T0wl2TBqn3KU1VzcNB
BTVIQoHNCukI8PA2dR8v2l6ETL1KQEfBndvGn4bPmleuiMh7SlfNtYLWFH0OVPza
IMwoz+W18Vj/jn6r7u5/vfS2pP/G46XRvdB5EcrqC9a7toHTRdaS6X0aLKhC0kek
WJoVUV0Fnixhtz+XVst5s6mYWuW8fgCYkdWiYnhneRZmapLWn4UuQLvZJ0KgmGCK
pDjtZ1VaFe8C7KknRoF1Ojsrwv/KpN5Ug2tW9mJfioGDSYMvOr+Jd5BdCPX0jxxo
1wg9X/fcT5kzZsYaPP71QuCSvmcptxvU2nWit+orqJRHAha1SLL9RvJIjoYLWe4t
5McmBtcuYcmX5pQ2dvfQzN/FDtj4PB7VAP51qy1vDp4ttD66BIOzh/pTRm4Tu0k+
0wx0EhjSrKqav6RVNUJLEmtpgm5KgQ+Q2KJ+wBrjLyM1N9kaCiDYN00k9b7hp2eK
t25Xkd7RxPsRqWG8IDsKjded9FxOBceyrtm/b18OrlJgJXU2cIK2RRDcDinX9JIM
EmHf1nQVk12jsYF3JN4g6oHG4Ff0o/l+t44ISbt8wDRaDXnlStIhuYcnXOyRVbMW
rIqdmFB5BGvV9PUcdnsrn4sLQx1vNXq6DnAqzML78PctUOJjvhuRxG1jHbajhEia
sdjdiz0/DoB1HZ0Sp/MEydAY6Axke8JdA7hjuZF/7R4DZn/aSiVCacPdMm64xO+p
ySGhLk9ZZbKh6Mk9WvyCaiq1XeiT1e/MlKW6SfU4wgZ5dT1XkgXXB+D4YWQvfRBg
WYU3MV0LtjxCDdJ3oSmtSWx2lFzsumedt6o6+q9Uc+++n24qjFN0NGNdhziERijf
T5luDqnsXt0Zwd5I0F9wrLWyG5ym50ynaVqJANvYKIm/1jnWmhFWMmcrew3OTbfo
2wMljAgbh5dV4bfe76iN+hUT3Du4sQWA3BZoo27Uv9DEPqXGICC7MsKNAE5XNcuL
yWcZk0I7mqBerOfocPHbmsvaAIPd+3L6P1vjtsMNQyjod6xsRJ9eiTnd1qZ0KWD9
DhsZV0QKKDvjKfDtEncmGSeODrhIB9BFDlTj9sYPtZmbIflWPSFJmq6Aa8S3L2cu
BcknlRtN/f7Dgjn+gASgrlfZGY24aZiBG3x/KlJUOaJI7DSBarPb9g+Uk0/oAVZN
9KDa9TrZMpgRcTddDSqKc7hK4AgcZ5bwlTFuNViN7zhEpabn06Hc0GYEZBV7kFeG
st42YWfAI6+LURAR1t6uynKCxW0JQGMUuaXDKa6xBZNBKhkToP3I5xc4xg+CUyTW
lvMD8SI2mJ5G5ufS/5NF/nAxbfENjVbPSlYdbP+mFK8Tux28YrXd5Q3lg9+Gq5yI
wCCDnkVmtGr6kOifsCetPvlfbAfC3jU/SHf/Gu9OiYXOiHbGG1D9OQcIt3x0vPzb
dZTXLRFn7YGVYlQkRDvuEmt1UuvMrfiXqzOMVPnnqveARt8CpW9tCGfzmTVYxQLU
g6FpdMSbo07FQVza2wCHN5vjf4Uqwxd1oSQ++C9YxxSCcmFKC6010625FIypiUw2
3Lsj2qag3+SNK2xGXxDUXY2N3DjMXJby1fQXrmOYEMhTp9OvwRVME6+E8f+35EM4
MPEKBVsS+6LhSsbl9nPm4nf7fNKRDyHy2c7UqyXGFs8EV/Ht/Jn6hCwzBOsRSTAw
2BbjEmjK7N2yYqYij5xQxvlXT3XvjYmhLlmTzsjgaezszSurEWXHsz22TKcscqT6
HjHlITYnJhm2LREJ4qnl1SGwfVjWQLVjHx0x4kUzmcfx0FVAEDpdFSEBN8/S4+Mu
WyOKUPFiUAawVMIA+PsotGN0I+MhlXa4HlTcnTOagZ8uc4jCp91hiI6q/DQajqEa
rLfjgoRJFqY7AFTPhYEw7cU66680MNYvzt9BYHXGRGci0uG2XaIXhJ9h8JaDjUfz
sYmYr70XC0TK6oy5kA91Y2sp9frE3ZP4uc57GFhKKg28GEiOO/U4hi1bGT2N0Gvq
+StgIvhzjOfQSk5g7cBsRKMoFILxGX3giSryEdwIOmNCKjWkDQB1TUp58S+aciTq
zyPl94t2RDi8IXkERnVVZhjnU8EPZWUN/pxiULUPiMevLRCAQLC5/x1U5NK/ihzW
P+/JmnC8YoUPJL5Fo60fylrWbsSsGRBtRQ7hvWPLli9Rz2SD2shCgez/1e+15KC2
2e4G5xCcdydOpV6iWDR5LJhIh9orCyyPB3bv62ELwdsXOW52BGhJhSuRLEVi6ifP
3kol0sArO4Yfrb12rvUhk1cKQCTw+x0/xeelcWApZcaq+Z/NfUZj2Ce979xOtGDI
Mj/E12OK/bZ5uHn4vBD0S0+VhfiriMJbRdRi9c61BU41D4xCsDe2mI8u+sjcUwUx
9hJ3GEAeUB+s3HpAfwahttCJLHKT8JCFyJHsNptDtPTQn4Y9epBa5SqRk+3janiy
UVHBOXCHQXSACDji2+0wn7KzHBbPA+i5I0H51I4XcNw+Tes3ZuMWaVplAaVDu+XL
WE5J+V7V4ZxT5Qu0cR4WDPqJ0s5Ug+8I/h+sL6gLf1EtPitB19LpsxWeReDI0PLV
Eps8pyol2BB818cPMftFiFbGGKEo78MI77KCMHzB6LdaiPOn9dL6XVnqNnXob9iU
PsvT5IUxCB44uPLifMwswdWDSMu8syGRTwyI3SLM/S3Z4cgeK2anLtoxrYYzbgOb
xqGQ+21UeJmWaIJiS+0vq5yqRVztCNrcnCn6RfAspgZwT2tBNGOwEnoB+cZZJnvj
C5gIuYMeAZZ35w5ThZuwVnpVR2PKgU6rncCI0X4JXxl/rHo3NC2eYktJ8hdbPWpa
WiTw9tJuPsCceBhNjSjytWMdGlijo5E+EMDwdEQiMQi1mVm6X++BKrR1IAV6sQmh
Veu97BdxMryCQW4v/bN06O3M8Q8lbSMjdn6B03exxs0gP9I55SPaR9vKaXjhPd0V
/C47R+qVtcE7lkkmedwj+GwovtEOrnZjAKrMXQMKg0RBTfmK+7nxaDm/ijRGaT03
j6T/IjHMZLoliuZuNb2WdIu7+mh9DWRN1W9oIJXyrlXm7QEQLxV0MY6AmP4srexi
2WA4R0TSGhwTXXGZrDOoYMvT+d4bDHyin7vPDVZhv6vo6UnOmbHHDm71OhV9mmeh
a/Cva5AAuXKsw3wTYhoS6mcB1749dqgCeZSpSqKD2w+FE8AyfwUKItyszPVp6oIY
4Nw4Y5ntb9VdBYd2Rm/qFWwF+TTgeeVSp39bxW7/Q0UI0YvIs5SWnzIWtl6m65yq
2GLc66/eVfTZrNxlIUNz19uR6ie9MD55RGhs67gm4SvHasKe4WdHSwx9tHbMOepX
1sFfykfy3Ope5GsPnypeMTRZ2PbvxRr49qDBkpS9YKwOUfPbqEKyIvbzsCjyNvtt
caJy4FMVzcZah2gjuwR9cDXM5cyWFrz43T3YeiU/Nlm60hHMuu6qhfWf0J5w2Uli
DCeu7ucyOGAacDTQchyOYHPiEwvtxeIT4ea/EkG8E4b/B8KIn/QD5qZfushSQloI
hCrxE5drpkXcNouaHS9sUiAKuK3mBWPu1x+AN2/YM7i0CWhW4o9sU8BZgBqjvEjz
bcSXmAhS7MYzDJBwmsG/t3vTsF6Y8NPaqL/vn/YRen8vuKg/Q+BD3stWypvVPGXG
kBSUc8wfYnp9qyKlhidyu2wAk+up15T8dQPPwX9BGEWT5RthJcReMJ4pTBT3Bp89
W92bySGFTRJp8KlRa894Hx4JEmMaGYTT0WO2PNA9dY258X3Sxvhik7tdi4dY3BHE
tKoGpvdg5uC6tlsYFEcDcH1CfYG6TcdacYIZNvVj0Od8DV/krIyFCrB4UVtuyRiw
Vl8+2RjBHGkfi+gJtIx21ZVNDNa6s+cE48Ocq8gb6eonAt9Tc2TzhOxFLHgYKqRT
MxUfeHM7OJnEoscPS2sfTei+pEZ50BEfxYHfI/UF/KZgHJ6hhUQT4t4HGfREJtq0
0cR39yxfptJYvQ/Kl13w6wpvqQ+Tpl1Kosw/doC8xRU8plxUIbcSLxS30B/GU12x
gNhmWjeHdgkHwz5aC5lOMOqLm7pxS1LWjCeOd4/YEXu/XUK06J/jgB9G5kKF7JwJ
QhMhqU/2tQq1fEREu32ws6/xnupjJWbzNuFgjYHzJAj5EF4C/ixz4SGful6zsF3L
pzToRZSjpf3MpzW9HVvUDh/GKSLOVT3IakTCKfcyf/y8V+F4/hAkDIa6J608l1cX
SfJ1xAoQuNKlDEOD2yqxApcrqtFT1XYp9PpIjrVz3qftVC1MEFIvxza6+kCFKSq/
iGF7W/CSEyOn3lU18dqb5iS2oluKy3Sx76SleZ7PRVPQevl4vNBa1vzU38GSa6t0
3CeTbu6xo5B9OHHZyHHG4ZJ3iTERvifw8PuPsYWZyORlVvYiiJ5zEXLcYjkV8m9O
WzSqRfLS4q5YZ3mtp2oksK84xyX7MH+IR6wiE7WvTeSVEwMV20G6HaFWkHDdgFyi
mkLXA/h1kPkRK837502QOnIq2G9irpYob002/rqlCFkyGsPRzEaT2ibRGtEgomvw
+E7p5yCj1ThHGxucqIuZj7m+AEE6Cg6qTGMW/vyrWHxxAivjiPS/s2wl16e+jXyR
pVO2BB3T3VzpvMWjt9IDlNL2E9kXKiCJxR3wwFJV9Y5/VmOqDa1CZCrkb3DFeavn
7sA8iHoNMqqrYOieN5WBiaJWx6la7l47JIDuTJ17Re+Tjn1aV0DqvBv+7ElhhOTd
wt0XkewrDpUYcOpL+63/mmCaWLwgdlsfGPqOuoI/hT43Gh/HCKfigiVSVXy8qrbn
kKlzUJgl/vcmGeH4i+j+HvvJG5V0BHn3i4/jKzSAviAV8v3qxPMqcAXhKIRWrNGF
OoOztzYcr+RF/EjqpBwf1OEqkovx+dNVvTPyxq/BZaJkJ8XOXzgR0GzthTqTQP2P
FULqzUAYn26r8puc5+ROmPyExw7tOyjei6mMfwfQ9MRfU4sNknX8TbxelFgu+qEG
9mVWQ8QL0yk0BOzq/mSxZ6Lgre+rwyIv2LcVYhdVoselpfwubXkqmOSc9i0cK3q0
tZ4LpiwTWJesntBIqPV1WZdB2Cv7jsWulaeQwuqHfXRM9F0wxiv38kTLSZOvKhRt
7+vnA2wsWNnkGpHHHciFpq6fCdsqLOhFqvIcrHnZ+09kz8CsTSSmUB0tVhbStKC8
t1qsWJsoOFtLobuPrNdBC3XyUaaHBZ51Gy6dgIYYygNPeHVbjRaeTT1OWcsoAJHu
x6OwDWAcAQ7JoKgeghsXGsIeRmBwwqJFEHGUkebWbWyl6ATNHssds8GI09FvTF/V
RU6BGSXfiMNUE8TOVrgJJ1SPfUssvSGSU02OWZBAPNyGlPpHhWougJDIhEydEmAs
Yclvl9c3kg36pO1X/GtSmuFs6uCeDDs+E7O5l+nR38cm8AN2ViZpw5kVnmk8A2h/
s4dqhhBDCU4xtEpGoqC7tIa1Hl63iEl5X+f4cMns2xzeG9r8beN9k8S+BB+EOeAt
U3W/90MxRQ91+ZHqoekZR0Wpv2DF95yxwYF1PPBsPvzAyIyIgvn8a1IXDwpT0c/G
jclEsRKOEEjm0RjDddU9e6w7ixA/orIp8xdMgYMlVajcqzEdhvQGagaD2ZFnjPtW
3n8d4SgfqFIGD/SW5gJGhALIFzwUmVktD9u1+TZmwtjva96aXwsKYME/rmLvvo6f
xKLCDgqtFsBXtz5uAa1algh1VmmCIap+SSFxoo3Jeehuygy3k6tcfJRvB+qRTNd0
JE0Wa/Svlgln6ePsvZqEnMx9y55BOcebjSTXB/AHehTBZTNvhkBdk53oVrz3QJZd
o4WXHnD0vY3KfrZUd2egvX5hwzTdxPrEGfvltqw2b319dM4twbBA6axBBVdtN0jr
UuuO05SULOCcFUrKEVbcGeZPkAp9YQT4z/kzrnP+Kbx+YIX2UKMt135NVWITel7Y
Ya/3HGzig68ujfc3iagI42ThRCsmrzGaGRXOvW4auJ0nDCxLoReU8f5a8c02r5v7
wZBEAOlS1Z6wwH+jxOgIYPXfGJdHb5Lplwd2LwiOtroa9s60W7KtHgpVM3s9lmg3
oabxuc2A9sOUbVNB+v8+s1nWgYhfjToqpOsS2nG4wUKj3tjh3ucrYg2h1FpJj4Gk
qizfYXs6874qqgUy/d+zTSftHFFo83mtAGQ05Uoy0iDAtd1vmNSUUGDDlorZLKBj
i5clPKbr/PhLIP6p5EXmyl+jPWLXFvoHJOqI1GNNN2W5CMPXqsWUA8as9udMdGgy
H3YhRj8G8WzLRe4ScVK64Sx0rlP6HAG1XnesP6CqFkcceuwKMPeO1VcikFrislWE
Cf4+oI821WTaMS9wqnpZd8TV7NQZYN2lq43V2/zh6ILzHOuQqNscgErRfoANLu2T
fldOa7f8sHsuiiLXC5qKaZUDaE8BYZO4c+hkXaoQU/TLH6qkyP/OT6AMiHSZGeAk
XbAe/i/oxHeHDO6F4f+j5B98Uj1iDuPW4U8xE8gKCfT8myslmcRjNV2YQ/mL2VVC
o7sZWk0v0XmtwnAHbPhwen9zUK9rc5s8ggf3irYRdOyM886npxT0rjVhU0slVVm/
y2YZui6da52O+ZcgByeVFzuyN6CWJF1yzfL9T3P5aWAPctJK+MvxE9ScPXog7/+3
8aSZbF9l5xK0e9Hwi4y+fohP3ujqbqXv7+4dC5xKOfFAcTMaDDhR7mwt1dPplfci
PJAKVMHGCsrA2jNGOjjM9os4UwNd67SkZHPvMoFkvSz9nYOiIsVX9G3eGaJndrOs
MeXVMeudb1y60DV2na90GZ+gVjObqK+5G2GSwuyT/SmMeyf82YV4YL+Wsm1Rz9rl
N5T+hYx2NDRMuvCt2fD5Zpn8eICti7Wm4J+6oaH5MBfXvWHgkrQQ++HZmwZxyVUO
Y1lgBNTuBBqpSfrQ+T/7uuIwoBDs0r6C+oFxs4QWElWb+7II+jcQUrXIiJBffnh3
lYn3RdspRq6WY7z2g7/UwdvbHNvdfii7ldFNWc9wl/GYtiuzKx5xwxvvqBzt8Dql
tCwzvWGMyqvIFCCbf5/V70BmvxPY9ACFBa2Rhqi5aw+YcCmo0PX69Q63ma08ZtFZ
U2bYARQSMhLS6sK2YLAp5JhHMneqvX7UyIID+Ut/gQYBxLaISkGzgg0oSEGhfbQd
WafeQa5hmQZvtDdih70h4G8z0Of7/aOkzI1zLwixbbdGx0FYHJNagpgzAiJs2RC+
jpqXww436ktKGBZgmfz6jIPveuFS5q1KP7VQsLPhYf13Z8gk3yPIll1TIveIQtKP
gqNPDyBPm4uY72JxZ4kFL++66lUwrVPKSXhFnZBPOoC7JdhzbqHdHBAG5HGz0xyU
pqK1P3Tm8m6tvpL0yVlT4wAjzy6W5eM38wikx+dOC46xqmdem0YEa8tMstumsgc1
grognurwwBsTPnvGvd71ob+ZYc8Yphw+BGK028ErSePE/mfj8kd+jIl4btkRtFdp
oviFMbwNavwdlfMlCCF4GxsXUvnqq/fNyiGzi8yO6yY2/si0A6m6E7WgSilf5x2k
GyF8rKpPwGgqIP3tu4RjUPVL/sim4hjyLSQ9aPFBMgst9vx4A/oA5LRAYmu4PAe7
4RDDppQDXVnL3a+La1XBVLGC5qvlRr7srT38qlvsPhQDhtDbysAM2g7ZWWtpq9JC
mv/PVYSLHg8DjlbWtG9PanX3woSCyw2zq07PNM2QUt8E8jLNcNMcG88IK0kkc2Qa
hAvVsc5YzBDIusspXky/C/fJ8xqnUSlPYboKKgOchEkeOIKdT9YRLv1kXgovzeOy
BHP77bvOFLODAbXIyTy1skfcos6q1xFz5JRQtm0o7wHoD94BKFEz6WOozbnku34M
KUeJcqDYzrrOFqqEpVmQI0JGrkisKVtXkdgC/3xHkWpaCHBVOCMz1G4IV6Y9/Kp9
XTFQd6txviioP0bdynr3DzXtFKW4wULRSsTVUEBU9RLjM9nMktZgoueO+k+XHS48
r9Xlt6V3G5nGO7QSGT8RYBE3k4n77RkegC8FH6yV3p6AMCyPuuDTrWCO2k7Okh1u
+qSUZLuGfSuJp9N0dwLSgroo8GScwCIkej62BK8lNn2EOHm5AKKuE8YUItWOnBsy
71ePqwa0dMppdOkdhRcnGjTP+gFLNE/RA7a1Hp3l4TEUYoiHgV+Zr1S92zwRVtEf
djREdMyeylXRqbH95hrOJn+RJk9Pzz9nmYCY6ec3vyeCekDYMul95ABQWoLM1vyZ
Hw3mLF4jDkQ+RO34cNpzgskU6Yt40fRNjOGgzfforBENwfIUAV4QtVgCGZw29Sex
0++hxdpf2GmRKove1c80MOFEkhro7q/0MSI51evNjggvnWpGMxviS4SBIpSRvXPR
+CsEtnmhrfo9Q52MGV+zxvBkhzrOhsifKLRLTUC5W2ZdCXWn8tYawTu9quH0drxz
+AfGWnTtJ0491Wp01N2EEWMfTj8EDQutRoHDc7+hLex/4ou/2NY1Ptz7FLb4O4zZ
eis1bQRvTLYTTNAuwNb7sRY/8ipVHG4da5adlikERw3dVMTtGrsTP0aPiHqVps9N
Y/vT5IkR2gh1ulb0fdfBGw8ME8tRBV5x9FFmeLXv3JivImKyqphcGjwXijDSOUr9
7Lw4nv2gOddqwO6z2MQ4w2E7el7qW/FnaN20e9NAM0hofhPP8XOXX1u8fvGc6B28
/Mf6VSPNw8p7kyu8Qmr/5sIIK5vo4NqpLhL5dzC6fuSm6ltBXpvbY/PkQAkn/G61
8it8N9qd76XuNxKr1Ou0zXCinXDP/D5DHblZL6HPxuTJRVdrPQRDW2N3B3AK3Hv9
qitW5RlHZJwbLtfSRD7CXu13DfJRTLU7VYoIoelC7pUGAzmQZAjEXaVryT7w8Dy8
KBqELEVyNAF4AHhtpqw/3OC4Qr8GsyYN6wqLvfuM+ek+GuxOR395Xw0SsNs9KiXs
GXAivgFVeUS1FZL4FUl2FnfPXFAQjsnUVibbDJHZty51o8HWYwJYM89of1Be6by+
/iaNBr/n3OsmV5gwiLavEYYBYfXWI1erjAXI66RCr8TVnufnn5fREU5xkHm/pbFR
JoX2ZtHAjQeD2s2bI+m4zVRgHwHKJnrB7NTKs/mtFYSRbnxeq7iw0lQ6YjEsWv+x
mdMAh8QSiw5YeWuzH0tfZeuscM6hr+gfB1LnZOJIP7qfz0EERkOImzTGkyKlVet5
RgJhcSzJVnMSChlzSkrLTyzZEUa8xlswItpv1blKv6tuRo1yJHTHGdGKzAMZGhbG
yeWoYfQ8jfGt896qSE5eMwu48ROYP2jiWretOWq+l49iAsnUgzaG8qBEXjy2Zb2F
n3oJ1jGa1wLmgbeAYPdWyxr+klApbKjT7Y2QM6ymLcZ8f0pb0YymC74DbujXUXRr
9mM/JV42B7YpZmakqjCQ61jhMuhIVsuiXDKM/t3ynVrtKZ2EdpnwgT6jX3c+bTck
9JNDt+v3av0PZnnC3WJx+SWAWAbr65R0TMKjdsnYuZqzH1FWge+vrr1/iAhJyebU
wAwcEBk+Ma9/HZN3FgQ/deirFE9TafcO8RH99hQ9arhpzBnM9e6v/4d9FVkBf5we
2gao1jMpdzJ/ksdjPJS5RIg0x31z9aAGH+4rdczK3u+gYYb8mF5we7xzl1jzKQ1+
ojcX2bC/XBo8il0msNDyN1q74OcBH7JSfwlTrL7lvWHil1IFlK6SYpRhRC0sTPah
0a16Fh48uPvd9Hi63VIeTEe3ycq3xWWA/cIp0MW7eRzIyTm9XwSgg4mT+Ma0zkcP
IRtCWqzuzhvwe5Mz0VGcC7p1fNKAloH9OaaN3vrAMsxD4HHNIKDt1zCNJJIou6lw
ecniEqcDXGnm3lgS1lx5oihlul+as3KsiJhfUb2jBpiBxluprBcbXky9YlZTCc9i
CL5tKf+VgXCZgRji4APztEbdChBtzMAMB0sMYOZ11zg6zX+EU2x0BEf1qLDPm62C
4l6Em3WMHu5BjwilLY4UarNZSfApK0a8mwZPd5LXheGpf1CNoFBO5CkuJneIEZ/u
QySzvs7fg3V3XbPLd4Kle7BiqswXRm/LCNay11CibPydsgbm5Z4XC3BltbTWbhXJ
5P5mDhk020ZxWjY+RCfDmK4M3DyEPdG2Dhwd4Zo75UAThbjvc41Uf1K+WoFqfYTY
4lY9xePXq/ZkXX47yn77EO1x8r+jvSpVLXtIkIfA8A5Cuw5qsnHKpcxCS9dvh4zs
bAVexnztxCZLsmIL+2j9PJ20PoyoxFK3izNAeDp6qBL8XlcHe/+DihCbumiW3GhQ
rbpoJprxBMBDYvI3oiZEvyhJf5mZd72JJpLax5RRE7F4ueyQv1jUFyHVJftyFYX9
de8J0IZtVp75a7bHEsjVtTWTZYfxC6doAsdTLGZuDHG3WnV9b9jHS8wxaK8LibC4
F0d7TlI3NoEc/FNtaZw5vvV8FUpjgKQYxrHaJ411W5Mn9fx5EjNgI661gOgrnDkO
/m184dSAVd9sakGhf2b8XbnbhOZ5UEdAAyaaybE6PVqf1KLh/TlyauWaRwEcSTa2
BESZyjpkLMBFiBRPMiHHZTyeTly2PGU6hDDFqkoFFAt28/3luKBr/JwC/FGxIOW8
eJqaM60sgUronUq5RxCL/OzznNxGcfptff2erRf32jyOhZKQhBKiLuHa45w2s7KH
uvE03J7WgnSL7fOtopBzLWKma8kmx4Lmx5be73o+jvXqOdo/JNLoNdJfGoDBbSqe
2eFff5x6KvHRAgNCDSogExigx+YN2celvwM524Fkq/yuYeklMymTVn80cZIlzLCQ
OxXKt4heE5z6ZK7BDThPFE2csEMtszHo2RocZQl5BGY5S+DeVBNwhh5THuT4qEKm
cKDoJfMZNC2ijjmt7d0YUEQblkWSi6Q9aFhLBCO5PBDi5rBS6DqWIxdW4IWNw76v
DB5MsqqnGzVIrrFcoS/vYefbl2z/8JggyfcCgSjd5aoSdW1qaCbTQZ09TR5GStUq
lrV/b2AcwePJMHa6mll6FDeLtFWJTNDuPOIRJfnJ4IWa2NlqaXa3QXsZvdmSi8s3
wbY3zgkPLnqkWdK1OvjSP4j6NhFOOR3KC8LFrzvxB/Uqy3CFr1AU4UQ/K94S8U1j
1HXy5HetJnr4Y9ZyXy6EvvDB2xSb2KoftC6gKHn7q0ViC4kyRvm/ld1WAAw30XVg
5VFPZ5GuYZuJaijOA4BKTmuA8E3bRar0GpM54zvT4OmLZ6Dao/E6hfHmPRw543DE
wbrQ2QJqcJknjnnH9+HnMAxb/wtqY6JzpE5eSceDWOEaIDq9nWisEXeK5+22oARi
HJvRshmeNWN3isiZT77LG+259USg6NRvTpPicUvvYD/KVKkM3vOyv/XsdUY54CBW
eHkzc8dY7Loy4CxoJvgELsJG6KK9VVpraWo/TETtiO4epMZaIECC0MXKEO2qHOd7
g2B54QrfamqR2ryFO1BSB6N/YnGRjOO+uNEC2IggbaopIdeTMtVprwodvztGgj8b
DKFUvvPCmbOQikGfOQZnsgYQgr9C9sRvdeNYDMd8NyzEiVMiBkdW5b8NRwtV70m4
/48rjotsY3fqwzLFlMcc3hn6d9qzDfDimyV1bUSndIBqrcL5X0dFHHys+acPa9Gx
8wHI5+iYszbpHGFEPKHOOJ2o/3MNeq/8fWdxUbI67QpgM7XZ4F9yHxe6LndVfVZl
ZaQuI98mGx2uFaOjW7cnJPAl7SeWAb5Hgy8zP+B/kdENEl47gJfuyQhDNnnCbHbC
e9V7H2dtvB0DZs8onUyMI1C9JfClvgz5Bb8xSzJwFfH37bFxiwNAb3XG26f8AISL
L9otc0d2oslQKpE8hCAgk/PCo8ks4Gvh1Rhnv/rbA/2ym8PDdvy5rn8C6/oDYPrz
Xp/n4nmU+uCQJSe2Y/0702kpa116Z8PLBpLVeCymCoWWuzH4DPjoh5DTWN6Z/4us
XdSxT+iGsuPRNsrkatpeLSA8/Jzp+Xc7F4VGI4bMUhD7UtekyG2IcinrIXHevfXT
blrE9ZYXdsV9tEVEspvQu+gjbWky/NurY8IG7Uq6B2rduugguBJMsHgZysPRHzXi
Nvk46GB2pvqtIINY5w5X/2oiT4f5AFj/qPabw4icL3umBQF8uCP1vuDVpEL6OwrN
WcK6klKR2q8qC2WaOzYE1s98/oDOVzhyetczySw2G4NqLdlLW1H5aau6Dj0x3lZh
YiXrYWz9AQObQr+gMMMjHHkQi43zdbxhUNtZn9yRePIhoAiM1amgr7fU5Kkn0oqj
eg0sxGNq5UKkXTuEN/rz3nxv5K2toTWBLUF61b8/DjCtVIwuf+yD4ynSkp0ASqnZ
l1sHTRmVOISAV3PEHPsoOCTIg/nvVRvBMwPfY/OEmLd2U9gbqVl4p6WtnYS7CsrB
w5ijF3u1zoN9SeptVA0DOcchvw77SeLYAEiM7KKEkI9m4TcmPhYpjce9aB90yMF+
Uz/du0Op46oplYdg/RMETAPqJ1+2fZzMorJWjPU/iX01Y+HTH168hWZmWiaieRf3
u1ZlTcyT0pyO43QtdVvk01ZAaFchEed8rKloffkkmqO54I3MKFdvqSVoczpNjHN0
sq/gUOvjXQPSkAsQp7UnhG1Pj4CZShzEAIWSBLxRWU81uOM9IB2LgNMbyUbeEFEu
oy4sZsxFHPdva2t5BY+oYI6GuGW4NUSqjdNcO72KtCm2NEioIuSrEKzFlKFY3VOw
F5ec08jogll4WywsH+uPNf6Oac+Px579n62LNLjForWOkC9oNf4Vnl4f2oe6Fu2d
d4J1osDdaBXDEc5IMWxWPKyyZAF8iLwhftSDbmjkj7AxtTfPWlDyWWfd5oKPOQnG
JNLM+AjN74t9pUDcCJzSedzHNHTFmB4JmP3hgRsGg4AYoxK5QpEfd1eWQ/LIvOXi
AyVZjWRghJHHwQ3ux/2w92V/tw26o+CTNlIBfJIq5k3c7hjIIIng1T/J+rEFCI2u
Gb8Bw4vxRqLb0gE6h/n6iGHlPYQdDSKYq+BIP4LgMdtLwyu4iXGz8uiwChJcJcie
BzFPCUl1B1Ho24vwcRrZ8SHP3jvfJ4GyPXMuTcbh9nBDijSSax0ldx8Lzu9+N+K0
Hc1xHWcDEDRTudIfYslkpS+1ogkd7ybAPiqpG3/Icteyx5fLORzHD3/QbLF7Vway
G0WcFbowNE0BmuGMRMVFoiHy5xt0zm1ZOcUDKcryKCYmUgbcHK5yXTLhfBL1pxmg
Pw7jP2ay2R7MdatsV6iNZLn65rIjeARcABO3W0UtpydzswekSW0DgxljSco5z793
spda9APPnVYkiW29PYdEiFqn7esiGWPUxKllmvu4l67Cy1WaIWqWHdlpdJMaYnwC
nVAx557HKSEZ+YBQ8e61Nz3pEkE13onTcjxk+EA4HYNdyVn9mjWIVTP7ATR5jhX4
Bm46NIcI+fHmS6uZ/XWmpHZf5zLQ6VvkQxhEsuEAPX8cb0x8yujMtq+5A88ug5EK
1+U9qBOIs/xfvSxDRFSBKDWEjWBubvavp0MckbUGFcb/onuIVoGtrvTmI//1eQKw
ESgeeFCEnz9KWFysNZxp2plP2VzInrGBw4MT0C4HgrZMH0HfKNqx9MMyxcnSc1+0
cKZM0T3wJP5HfHx2CjAQ1YSJaNAELppW3W19o/T7WGZmS1NZDVtHCIZN9sU2/6xK
rwSI/44QP61opBrKlfBq5lFDGtVaiA7DMVMItaHM62MM8HOtuK2vbAHqDMzZQard
wsK1F3VMDnmWXG9h2z2nOZh3WuD/ZDkPLEdPLfgeivRIZqgi1Vz2AeUHhSblwV1o
SWb3Rr9SOoYNpSE2Cffngc/LH+tFJjPZbRzGEL+mQnmQoAIZdYWyRMqVjfGO+9oP
JepW/ZPhCB7XfCRvOcT5JioHglfpJ3xCySeCvBNcnQ5oLqrFD+3ZZVwmPeYiWnNh
FrPGV0DUW2bKJjipjWEnnN5CqO0e4OIm/KeUJq5/asrTqN9V9SQyD6dk+QGVPRFq
GCoTnhlkt9Yj/TzdQA5BeO3cBLqYvVvslO+F7xJqN6IBQ0xq8lgc+aHbHMYQ5ie/
VBaeNQmBDAagjnG+cPqgHlVmIhhmvFpsaOmhlUgfhY0W7Zm9jSuGGtDsbbcS8NLO
CbcNj9I1afwfcol0edH8RnAl2kq9VHAGebe5V/uB9Q04RrWt0fEXvW0NwQFNh65n
3UVZRjSZrp/rASnPP1c0cfkBsuU2dPs7g0Ywuy4f7nGxL6krsP+s62KiDOJn6xvb
VDC7RTJXo57bQxwY2BS/iYvDOZF5sOx7PU5RcgYuHCryyC5qdKSyhffsCnlF8dh5
xt3ndT4fDKxaYkdlPVxrqAj0XUHmdF61WKoUNO3L3Fkyel6HwPe/qZJyS5/iAWUN
KcbtWHG2os3yvuHGzd4e2Xhe9qHq0Y7E18CvA1U2NwQPsFc3jkU0Dc9Oxj/+qJzk
yN3e2ddplTAw/HQcySaRhCpICSwqPcV8nfdsBa4mdo799FlT1YHwPL5ZRMn/xSRg
bKetNCJdMjpA77dLfcQ39cJxJz3DEHRX5KDoGfbDckjVX3vwakFcwhwAOukSpVeu
GmARJ7nCliL9B4DiwLOzQQO+cca+WjvFu1kGeB3yrFoQ4qm5oy3OBhH0mzG9ZJlW
Lydko0P60xcQrh9KS+LV567/e+OChOZpgO5YBK0fNKGxmWIbadpUBNjLfbwoWQJc
iOy421KL2vp597cESFbIOW2hFnkmzpWfywZBeB8E6vVzQbxjjb9SIkEtz3tWVkh5
xe5hZTuWhfvS0RxKqnbNiN3ULqecpOqJB3CqtZDz+iITno7vNLBkf9Y9wkSfPbo5
DregonmwYn2W+rVBpXW7y8gpFsTSaOv5E3jwMYNGD+35PPGcHcjjNdZlQNQe9PmF
cEEIKMrdGk4QmJsOpnSF9gEUWWVHTCpMKUw6PSDbB4CxEICUenUNu/Cz4KqVoUPC
tity+C9B18w2iVpDlR7lDQ4xexXrFTYophnM/pgQ4KmuX7N8mkv5htABFHx06VUN
qu0djfkKNe0YwUdQyLfhr3CYvkIJ2kMt5igGhT4RBNzd/4RSWd2UV/M3beVQG0Hp
HIh6o/XoqKIOaJyHDk21RnbalruKkOMSyIFd3sqpGa/9VCr6wskyXfdmFfmm1a1n
klokhBDs33vlJ131WO4inFSVYcpVQGipgIozf4mHZtFgWd+g7h+uU8TeIw8l30gV
Vlz/o187XWg3xYVKq5QxOAYC4mofVfQwKaJepbSR2OxCp7UXLNVPQ6tTKduGogll
xxe3inROLE7bwG454pZ03chDO2k2MBNazIJMCOi35SbYcu1d7AwwZYLjFr6FX+NH
AAiFWknPfsBO6fL3ln6r8LrlD6t7h0BAFgF5xNH69z1NbDv9nnBQh46cPmHvhUa6
3+jXj4AkSS6fnAjrV/JGi/qJen0nlGy6OKYOtLVESGYIt8cwUrwNexC+12Q8Ti/1
NQuQt+YP3cT3gnu/7J73RTD3+JefACecjRlXxetd4z5kE9BnYXJrBvw3zqvPuEAR
HDCdYtR0G0YaVsin3G1q19AHi83uN6E7XPeFO4bHipp5sBRaQ+t0qJVkfV7UHm4b
dFrgfTBynBWNOf0Uum2yhR4mSBH7mVK7v28h7Oo7bH5G78VbXXVLOVEwHk6otl+b
8Y6D3DxnjBy7sDsxZ1zMx8JPJcP+v+VcY0CepGpQPy8TBXgCyNxw4InCrSCRWV6C
zFbD7egiX/3DBkKDGob7+6Apwii41r53zZmqmpgahcICg7ps++9IwA1vzWBBjE++
FeczI0V9o5IcbG4tpSJn+RuuxrqR3JVPfW9YKyy4ZSHeXgDhvUVDZlp/KuTpCvTC
qe7oUJ05inT2l2fevb846Ul07BGpt7YAk5vydpzvKPwTtm/JVC4agWcNJy/SnGV5
AQqL2vFb/CNOsJQhzAA8ScrV+g3WRcKjQDQ9Zx/oUQ4SXrNxCBCEkU1zOSfKc59R
1vRx/MZyYUMFvFLSHo8w7Hg1UE969xM4OF6HhbIok/8yO/MFsfobO41y1tgmcBx8
hF+5c6gie9ItCdvsSIbXSsFJ4NczGo88CX4amdFElc1lq2OV+LIVyBdD/adsvZU8
lXbpIZOFAHPiTtTIy1iPES60MTzXnzjSW0YY9qeOWvVlJySEf13p1qpvdaY5xVw+
byLC1RJ2YkYuzJD8kyoSeBfiJ7zgl3Pp6sDIKSU9fjklYaegXsZMvTi88LvDTFt1
Xd+AjSD1PZOwdNoWUZBgZvEA8aQbYpfGz6QnsqkFzh5FGg2uUO0l83Gc1EOexXaE
qWkL8Zo7X2B3OTdFt4uhjZuIrI8PXhXYVqK3I7edIC8/L7z5T+f9QHxTR3ultCc1
0AyADLX6u5KsBDwyt4qsOxl/OY+UCpHmVYXEzBmfijYfweDXKfofeCUb4LkxMLqt
XaanCLxTr5Eq4c3zYv1CzHRiCDjWQfY2JZhCL8RWzhhzopbSxGr4YklTpOcebpCa
RTdbMp36e5kqQtWVexLpa+OZyZjTOj5JFLy+aI61A8eb9mJ+yfa/2lzyDGvquUzI
0qDhM9KOlr3nhrVEAeo5jFc/PpQfdDnfa8WsmsU/Y+dvjj493Cu5p+deypR+b212
iUJPRS6IDuEyFCUzPjuc+BnBwWtMiLlZonML9TbDo9I6RApbz4jfGfkDIk82da4B
bBqvGh+95dhE62g18nRogwTMSdOUzjAYvjwhxoJtaJwfxC9zF144o0ZHERb4lcFA
Ysh3BFASO4KbWHeoGw4mNd6KYH2dqzEnBt4GMaV8Fkp7PPAXwJekJu6dFhxbFvoW
yWryZn/qclnMK6dtP7vaDfuKp+ygsT44GVKIDg49LM+95BGnIVoilOeVt1kmpF6s
U4dv4fOQRzNhBlBgPvto8uEMXTMVdNMTr4LCiljhVJixThNDKdK3nbbZga9waayK
4dpgGEGMmCoBHZEiTQ5gBvbpceIj1b6w285ZYFaSv6toi0DVXkByFeoz6L4y4SWi
U4DDIwuI+ElZ7IJnSZE6ZXM52Zi1EK4W1BgD47FouyeVihoIPQcx4uMlbWSZs/xC
iL6ODBySZjcpdwx2BK9Cnd1MVnvHI20UCiO+27vQmaw+zqmFWoqgv3QNOq/Qh6t2
8s8vIrN9oeFdW+mWRGY7gtkOh0L5U80xy+h0fWiEBwthmZD+u9mBXs2KjXpxXjUj
tn4LPDzftcxOf8r0ClVNvfylE7wmI+1St1lavDhn3WPIMv7jfucw+Cn8hM8Oe5pa
rVoJJk/RdSWVRFvougFFifAiXTu0iSF9SRRGIezsnTqLxD1S1EYdVHLuBuuh5Gip
piQOzUMZ+VfkF6SXcCadJLj3Dcak9ShGq++UaWVHk1yp8COqBXXnF4N8RfzTgxSA
MinJGCOFj7lJ1UiKzn+/mYWdWmpeg6WxJAhJ0PGTRHthMu+MsarqiXk/BZpsRFfA
9ppVW0VQlIHRwMsjOKG5OQ1MSSn9a1ryQBpb8VucPsmHec+/dzRj8FbKevjrG+w1
XV6GUiXov9gGaYCuAxhH84+HHXUyiTIqlQIKqfUrccJIr5cgA26YAbmZ2GaS7Cp9
bn0J7e/tGBmS+xNdIrItW0CXXQqi1oUqhL4m7ZsjW1vkklK/wQ9OBSIZLdE5P5Mo
suHeqvIZP1312/N4wWDs8iywEQ378HItHiIZtcc423HHUKaxl1s89jvjbaAMhovd
I92E+MGXY4EjzFj+rRQz9p72u1Ejld33HhlNhW7FnX+AXX3gDWmnQG2aIJCQEmrx
ecfDIjvZgIC8NmglyJoNqSUaOrWIJiCTIXr0X3c41Kd0uN3bYJ3C4aRmOooVWKqX
817TEvlQglYxrQgJhX98AYe5iT730dOUrKas1WsqAirSHG78fdZxA4LXOzIZ7vOo
hU9ByssK7TqAfQ/OyvuGjkiHEFXfsZrsrfdibba7iu28vj8NDB8geiBm9isDj0dS
D70pWyX2xQlUU1t12S855WGpZ9+WR34D5eS2wgXWVWb5tDjSg1nSDNYNTkfqDKnw
v34eQ7MRz709/lFVLa4LGIQA5tOx3drjLDD47kBscB9HL1+L/B3g1vqEWstYKQKZ
Jti+n6OEikB3w0dei16zmE6bLuWWtPAdPa/Js6pzXoNh2O9p0EedNAJ1Y3+IZlhK
UzE8p+qJSLoQwpetX8jZfWlpyvnBVc1/cPiDDKLWL4oY+w7G0Y3v8mw9VI7kAHRL
rRjPSrltH2qkOXbXjAQfnbqRu1p9lnq/RwTIOk61e6xCYMv9mBly5RsTF1uwBqeQ
LHgm/30Q0T19kpeHMSb7ijRSbd23rwbaoVoe+eGc4zsl600VV9duuquFIjpgmV8K
m/W2Au4d0uLDVIaC5aaKwKyaXIud0To5ymjCnM6GwrVQXqqgGFLZCBhU9gp9oNp3
EiS0OV8hvL1M/5fUnJaqzNo+4eQf+DSGJQAPNPQh/bxc+nTKulNrBKqvJw35pkyM
HP8zYw/14eM+xSOy9dK8LpPLdXNDWeo+ZZlf9t2Om75rr4RlBlPs/IfsESAjly8K
BeGjp56cix2gJbjeaOlaGHEX+/YSzVhrAn3oLhnm00UHSK9mo2jUgoSjXDgapCHP
WwZGmhuH6DudIN8uahWqE0zwJAVsQ/SqRkmAxCKqxGP+WsOK+L6EymGAzhs1TOB9
63xAxxFX1o1X+hbJZkYNB+13AI9epnoWhaZHs47IZqSX7oOGWtDvKZQpkEIVj+sn
WKJOIU6xKCCX/nFUgo93GcK4kfpJbtXd+cmCFYubF8gJfjspLdYsKTcOLfaKqixV
WXpUcLp1oNTcglTkoKrekPC1A05/rR7WIu+fZZm5aJmn+g63UhcUIvTeWWewg4ID
zKVnkBIUl5CLYrk3VKp+0jDr0D/GWBoWSE5p5Y3br9nqRC6zy+Ba/nDl9OLg3867
wbeu5jDO2icNsXq6fPqyt5sod9Wd7iEbYfn7DXChy+1U7g8MdWyUl1SGwA2Sizgp
AcWwAf3UWVrUfjdDHie91IbBo8qKUXUqhVwSD3JVx39NbVoFFVUBFHM3eP7ATTEf
hX8pcdC39hxVQpQAReeYjyd2wu5D+SugMtJkiaN82sEHGAK1vOwyQUTTRxxGaAwQ
2tEMj2SQFKWI4S8yRaD2WxekElCq6WY9Uid779Xl/0aeVRBSdn4vRmqhnypXmfu/
oaUpNRyIuD3WM3hT968OwF7SwrlPalb0/WNmHDqg8Pz/m/sg/JUEJiMzG9Nqie0S
QxQyIQacZJYOF3jA72vuPB/mfS5ayyscSbONuT/qt5XPzU5GpRWq6JrEMq/EnTo1
8rtKThw9vyTniu+dn7aqELiA1khV61i9mBzpuCCcCOBjfH5lwosjsvsmgCgHIYrR
L1NDU0fvHZwHCha8B9ymV1EC9dr3miSCR9SRk7k4Wqy3r3r7A94qnYxOmJP64bl9
SuuweHajjQDqvFEDcv4zTCHYdyw92/nalYmADyx2upuNod5qoxq8rinTEzyeImfO
u1if2hXb0omMAhr+CUVG2mMLeEj9lgtAez4oHnUMo/1JZGMZaqXJ08qLpyWALiKG
XENbUkA4GL76RkE1AdLTvOS7tzW2xo9rHG4Iha9GDJ/+02rDt3uGJ7m1s3JwDI5r
7QYtgJUGlQTo7SmEVU4nVvGxd6kysLQsLj2Ea0ZBH0FKryb8aasCzo1d7Pqyux/B
g2gZBjvehqhS8kbsLPATu9N/NgcIYUHp44GK4kJXxwibI8zHTNw12Jp9tbaqFRt8
r5pZrfBJpZy0qHs4tSlGEl2NZBAUbCm4r74Al5qwJwy4FKxyfqpQjBfabKg6YJDV
9AHA8lNdm0lZzBTumRkzz/vohtKwyrgIsPa1grcZGHipTYNOhmSWczDbr+fdRqyC
z99AITfEbBwl/xzZmW5TQ6coTpcUi9TciVnKbKVbCuW2j7PK3Vo3SRRZLH9awFvo
LcVaDInj/fdaojhi2CGlDXLPwx4NhzQDYuDV7oxMNTC9AaNPQItDXA4QyoQ5V7Jt
0PW64nI9vO+z3votr/jsuNtUUb3x99+C6h9LYgBW/oAMYhlpywJ4sgah43A8Zz4p
cmysybdbNiiG/v2LUV4gLucbVRreWgIoFPA2XhIQB4jhAXh4uiSxfj+7XB45Fgp5
kWYXwKWlPsL0aybSdPCaZ5V07hd9dcjVg0+AVmfyr3ahvf4PaPcmkuobCa2S4S/y
U7V0qOl6fp8lRZTxEKz9/0CCXLsD5SteYgBlh7DVQ/5anJ5R1jt2MtdjGaPseAiz
Nxzi4w+lcw6thNeCZE/nA/jsljNwzzVJxmCv8pAB4Zp0dOcxg671TUTUue/m9jt/
BtSCZ7sjGkUmc/vYvYfSdIjo+MRrw/S2IPyr0zBup2nxhUvPanPgrwbJ4IaXnmf1
aQhGzzLvq3icYMA82AimY4vrPI8mkkXMQSHr4Ul23SYUvYDTKc8FKjApqTQ1L2S+
0J7/YlRi0GNXDuMxU03HdywRv+K0tSNroPy3b9fj7xqIr0UtcoCd16N3GPkOembs
bOtL+ct0ubuNhlVDqJ+7mBGQPxWmIbCJr+F5OOt8VbCKZHGKIMecJGcdrDumYi8o
R1fmzJnP3bgJ+04xNJaNvWAs8WWCJOuNsfxwyACyiIKezoSE0Vdu9sVm0ERa+txX
sjYBL6yEJidPUwYk42KuXroce4GxvA9xKSLV7yomRg0YoNdUl9K9tJ2hx2fKhukA
hd7/ZMhGYGP8xR1mYFDSA84X6skPx6ySLLNLi0IZk46R6ywlqLyZSKWP7zdJhG1t
ZREOrR0rhE1bew+upu/ng8UlFSodYKTwJjspAk5snpeFAuaZ0oROleSWxEHzo6tf
thkiMXPPvAqj1syMLcWiLlSjvRlS2wwkNgtuXw9N/zR+a5rknX16/zeTJ9FMfRmW
Os6Idp1MvPZR2cEXXndC55Z0fj5rmZOmf3wlMu0MpsfjSpb+tmzYKi+q6txrSAy8
9RpiHePfbGL50v0rwOgZWuSnCXSARadOUjbQcUYhJ6/kzLv52oyGBNiDx5IlufPU
EdeU+S6XLMeYyjl2C6b1KjWxnwJejWrR36Jwtz8sSCEnCC3NbBbyv4ZUC71Er4k0
ZaKbDJQPzggyxkuls0tWIgF+HB2MXTWlqrTmFy1cZv5NcK3eMn8H9QGb5b72ooxo
UuFklP11vmGbZyaMz4MNsxO1qr9/kZxfe+yPvd28NrMsaABTct4aGkK9qgKifX33
NW8PjRWDNXTJoNbdzDq5TxC6r9On41Eo3lLQPulwGGCdVB+5TuDc4IfBTlS/FbOK
Dghlj9a4zh4oiaDxsA7PVUTbNruva9DzVhMAwJzWrlEOubHo4A2VbjnPgEGjuKYi
s1QpZHJbOP4NuAFUMZhGOpLhGAY36XOeRp64yazX8fSvuq5Gpe7eWHfrWRefM2Tl
t3zJfg7El6qol2sFPgtUomoJ3G5UJiA6qvqAejCXInqWEGCI8R/AUxj+G7mdl22a
xvNiRoY+lZqx2qIwSCfdan2F/dGwy8VEHEKClrtS4qO7lHd9AJxtqmwlr32th8ek
PosVEd6IByRxCIXCbhQOCo89A/wjjn0TqlNnDez/ykWldbCmNtTw33JLPWDary5Q
dBmEES6uQWqqp6cfiPSy/KEBQO61U4zXIZVmAsnme8upGSt3nfiH35YzA8LMW3fe
GBKMJLoujpcqRorrcKVscpwk/Vu4nq/AvwA1ess2FupL2HenqIiOUv9Zy22cQCZg
ZcA35FyiAPLbHqT5LfrNS5fVxVmYdZL7eppunw29LEDD/WvEB29rF0u+5XJ5e+/d
zSes246n7Jzpv9E3tKb563QgxBfgjddm4L9Bz9c4RzPE4lmtHAZvCQjD5B7K4sqc
Asu9Vg8uuLipMgyqInWCgoVeF31xr/Vuq72N7+6kojjw88c/gulmYSjb/pr2qdHh
ZPCTAtPuJCbtq14N7ROq6L0VAMxbbrezixevEQfbuysYenMSwu8a4qjgw5V5Mke3
LRCTbvqkugg0VfYtDPSqoCCLU0/sheuXbvbiZ7H4gNT/txT6Au9CXFT4E51LgZNz
UjEiHDg17tr9tZ8kK6Jh2hFIx6ioJK2qyrtZFEiR7XpaVw3GKAm3RIyyzA1zO7Ct
G606ItqH7XmEwPsjWbh3VnduFMyGFcnhGKewvTrwMBVyWxQiMdfOf3f3VT+Ezlrp
iAQSnic0LxcaCvN6pUrYnNellzFTffGwzGbg1ngT1ijpKu4B6Zmt3WNHIK7oN9hp
lhFBG5GciHU6xhn5Knsfe6RqtMvPqbtTHmmgkRuGQQe9D6H/Bm/C9W8EfDtmNtfb
NduVBFu4ON0P7/CAIEOFQ+kp9t3rULdfXkwmdwthGQhFiwwaWOEt9lsnGplmd7gx
Dgj/Ztad9cQK7TmRCN8lz7MygLhC0Yjnoa4z6bIAm4ywqjogUCnh1Ief9QH/n8A4
Kb0ljyPr9fjFxE60NU8EZctlEECmKIc/NrKL/6O1rq+FCAZOOg24vd9FjocTEY3L
ixbd5Uo+HRdPV4CpEJNIloKrmls+YaCPlwxFuDf09cMLLHDRiZOZ6JKc71EsMCWN
4zduz4/Ze898i/4tdbE5h4OwAZyIN0HJG4/9PpHGm21xgS/cmV2aCrmQwvBUwzOz
+tG6x1bTbegkK/kQGZQu2c4ZlrlZ8IjSou/VSKvVv1W6n3W3EkdpAcl9sfDynPMn
A7ObXkXbV0BJXToqy3ddm6/5nJbVzYuL9NH4h+WN2KHTj485VSsPILt5CdduKIww
DZhLOlaFnEUJ85VuKlAR1S89Jkq04kP+c1h2YLIvg6QHIMyMI9Y6jFmXsA/TZ2A+
DtX+hlH2J3W0uxxU2HOH8xGczJuSgr8RniMDacS75x6ftosrrEINMAWldiOKW9KF
Qa+cgH33DP0MZ1L0GZFoWmsQQC/TOy/GdvOKadOzwdPpV3Uz44kZ8xQTFTy/C6EH
LNxtzStw9znlgzeBXtvvSG765lT6wmNByU/3Njk3FGqshsLFPsneZcRgvtuW7uEt
b4GgTMCbz+ruXbjjmvYYSYoRnSK1V/E2SFzrpJkE1hjyWaSO4e1O66GRKvKRv+QI
FI/wCaY6FWkyiw90zA4wEnIsbHW3U1XAj/seIJHZwPoMI+Jz0J+weWmz9oC9YQpB
iqW1Z7tG2env72Ji5p8FPKkbQM8rYOBy5I+gbk8E/Uz4VtdNedLoRmsaAJhEbgHr
0XakJ5nhfbcJJn/NPK/irJSZEDvlhlVwVk9rdRIE4Yan0+xLkTpPsLZb3UHaE0OR
QSasKeWsqPGvF5QgTF7oujQfXKGK/b281PWn49dcRoJtmx3ep6xWv2rNFke1g+as
0Zs7lEQYke3bWQxoKlXuKH0LMcaKp0KYxzvabuJAqTrEvDivAq7yJSgUERjcHs+4
bgex/FgC2aY9736Dh4Oy1+rn9xTUGX7Q2/GYuw09H0jA2TAcKCugqrppovio0akK
67dtzpZLKoHSaBCHyOnCCCjQAKPB7MW3U3I6ZHctChhVDTt6nR8iKWEJCAQ1ezuc
n/z2+TbNMOg/HpaROLUSWlPE6nZYhpiZXI6AUVlMIn0nWVqU47ZQJsrA680J95c6
KtJaAsKxQMcPx5gkG4hQexo3dy8uS2x3w9ff/K+5Hu+NKTJwh6ySh3IynAH00JHY
N30FcBIG5tTMmYcW6/U9shDQDFs28LGUiqh9jGhtY3QruktaWHpSzK5ty5awOdoe
mYhw4gUusZus6l5oRc3V0oHrTiDVxFKS0HXJYyJc/KSkZlNZ6KRsLedvNH92egSv
+Z/yxeryODuT8xCzWY00YHbVtnqkqWgNSVJ0OHwN07RPk8zEtwkUsQB5engEhpTC
aY9D/WFOZDzeTEVtdkHH+Fof13my1smRvdPDL0Oa0CfCfYJQ5KV16fAEQ/+07b3q
v1AJ5XyhwC3bgCWmXwrSofgCHBqce/I0z4kfGGDZCEdlbrkKXkSN6F8NI5SadJZi
yvJxIAXFvFluSyweUtSRVPB5u0GZt8HQp64tZJSTihVRZ/0W11gYrNx7+Cj1oE8E
he5lbsdDkKDoTnAmXMPteF7fNXMr2JZcI0qyD7vFE4FmSrG+/Zi0UyRd5zhSeRvf
CucTXi2XDQCNzE63mpybBkYAdadA6y9gfo9QrNRdBH8FtUlHpk08USgsZHgOKpYo
amFEpNIxlAzywy2dj7LLMkpXhmnoSOkmvSzghuV0JnN0icC9CrK1FmDLoYmcAaD8
uPmXq93NsQHBo371yHjIawYBs5ePtDPD3gQtfhxSiNR/BtKDgxB8NaOr7fZLtZKE
A4og0G10XQ4GhayOatmRIbzN+ip+HxbYEXzrkdJHH8/14PQNmG2aF1IJ+8w6jRoE
BdBPOpzvH9WCUe4mPTSauOid+H/LlmKtu8eFZEo63CFXJuEt6G1yFswC2CHruBzP
sfXsEFkVweps2/D9HKrcCXFVvybG2aldrNXSRA3jPAyk/zXJBr2ZlXyPZtnW0ueP
6xcmld8SKDR6B8UVQYyYgYABMiXB9VLeBwgi8Inbvhp9gR0OIPgGWzgAZRbKo6KL
9bZI2gaUsN1hPyIiEpFmzESo+DwDXoS8iuGWu3J3+Zckt9c+MsuPNG3EzaYCoZLr
TuYmv2AJhp//KeW9SWavtYhsRTxZLW/Sx766MW+Sy45/i8BeVipFfODw5+DxsqYC
l/1NlU+9HKua7slk6tXXeX+7eiwYAusNgymZ2OZH1QN+Xgx0ATyCVKnq4zt5jnxQ
CgfuTe+yKCQkxJhiVrsv7EV6iNeZgw4Ani6dpNHLAEh/KUm1XIubzTgq/icOESRC
Wrg8wZWe89rMJKO6lGJKIeVFjUbbqW6KVVtKcUarKxkFZHBT0kijnhoX6oyDLieS
hB02KxcJIPpFr6V+QLO9XoynbJD5Y2em2Ufe2QctizAPj5PjqxCY5lNWaHImsvfy
yMuW9Ujuzb9KR/uMyy6t598G+0jVoxDiCRu+2XvHzaX112uSMcCjPgXFjugdUZEH
+TCQtqZl/tLyeL6LEetzvXLb8SEcz7WCy2+EX67sHwYDA3ferJUBe9o3zHkWnNYO
CMPsP22QgSVtsT7thTs3bbfpgeYfYKOzF0mj1yhGIvVA64cDDw39a6as6fE8bveE
s/eyHtxq1Wy4qLH2T6ikQNwbcBhbkdcasrQnbhSz5zYySeFoeSMFGpckcGHcHGAq
gZGE9fCXHbiHTTqk7+gOePcZeoREuI6gD2EXBBIwy3cEcl8w6HLHtVlweFZUdBBq
tI7NMSrilv8YEOfRvSAZ1rmPPEJRrmXspZOvSYVlhHvRe+vhsUIaS9RXnl8BDvGc
cH9BBNFpvQYyeuj//Ocq+AD5tKk7nZETsK8ZQri6NFHaH5fXngkKDARI98k10tO6
fd2zbUwuUFMh/3Fd8v6JAUYs7t0FkDkAmA905Edw/XAC0QAss6RNH2IK9hOAaStL
D+3cBTGoHPO1JlUzQ0XFr3SDBavU3X5PN5dSgxUGYpWNCzVJOLW5caQrv6lfwZ/6
Rxa8P76e3A0++At+W70a/wi7zynqk7Up4RPQgdGbfWZUno7XqoP7B9cl3sExv7hY
1DT+Uc6ybMBZg53ULncXEKSa2ZlqAOzrRvQ//kNuX1IJyF2WSeZ4JWijeJfuKS2c
NxVp9hKlu51/C/o2ExLyIyWTIrnTpb+tnJ4ZaAIR5nJkAr1ZuR8y+nc+wj93gO0V
W2ZR2Xsdr/NFzij0F7cBt54RtVZSf73d+/tD8w8pPV0DXa3d8veAn45EuN0u48Ng
ub+eV4ViLVC+EgGvOfnQO4gPQSrrr6AupwBL1crHBjZzem+5TYZNT2WpIZEYveF/
hv+FABWbbHQakIr1db7ODIXrKAG3N9WbEtVDnk0eYL+IuHJehmTAvfhc4Hs3+VAf
d6skUtV8wBEB+IhJRZ7xiwU2YinMyrvsbMIFgLILQ+0+UHtQxv2Q+pPgrdOfc+/U
d2JiI2itJ4+mkw2AMvwtP6mkO4tJHIsa7640DEDh5uC2rFgPwf6ne0xNPGyOh5Y+
skQE2/ONo7C/F/ajKnw23ehUyipYFnbk+87CIvihGA/H8rc5g0oI2ULfNmITr5Ur
AkHIjjc+yc1c3WTR3J5ldw2QwPFVa49/Oobel7uIGFYK58n+8T65r/H13kaqQuic
J+tmzuIgBJZf+ekPW5B4L+ow4FGi8flVwe42dVpJv+Dpgdbax8omTMGDtKqRMJW+
XKjx4r8Jv0SXz5kAiXg6EDyf9Pha7R/bIdySwkQ47G/rukQnLzqJTo/qEcaA5H8v
47qKObi+F4PqZdDeYl84ZTQyfL31ES1/47eJobNEFE54TqplKYZ1rmGdxRqL3IML
U4DJ8U5m6jIh7+NIvdnha5aRtEkue/XshHNNrPEakszqdrAG2FJDmKW54jk0dh6G
Rem0Q6E6aZYU39v30LxXQEhgfazyTm64cP/65dV9FzyORxFcEZ5i0nAzoWFbHdTs
habFG3QKXXbCptlzmEFPw1NsNqS+8RETfEFDOd0r7Lhznc/DJW9pBiOw6cj/6G1G
G1thO2HK4pT+C05lRpYbcIrdOQzfmOSe9s72zq3gWraWwGRwkUkNqVOn/BMV0a3L
y7sfo45mGcj62LMfhpRDHx4i47ZcBTfWCh4kbKHp+G+Yqqs1mWvGPHuZXNmWa3/a
KKSjI25nq7gZ/a190Edi+2xySisJAjpfGjJ88JtSpcCLrWBR2EAnATseud/ifYqF
GCP0Yd78OyaV2h65Ug9WL9CRXKYNz0jnRsoq6RX1OB6sMbLAEu+1wNr1Y3d/wzVy
9FEZlDE0HN7AGcBpESffyocSnhF7VliOApIv4X5icRca3zzsj6asJA04oIppWHmT
FcAhvzxqOoeJeQh1SyYZSGfr32oiOlLcR1/hvyOLYTfTHv+gwGjeu4faMciDDsF/
IyTsqOwVwy4qTsYmZe9MuSxvIPloDLb9bA5cW9w2xHqDz8cAOTflhaGtxTSUTflb
c9+001NlhLUxLYGpzJNCl8VCcZKynMSxXybHJqghr6rxF6N88VrZ6ZiPX4azDm7V
Hz4UnMTYPx+xsD8IJfEy6tDrJKrSKa0YiM0gTw+Fs8nBztiTRNUd1AEkD8PG6H3U
TrqV8cjVQ6PF6L9sQWmztq6K1g5gtXlV69rptnXIOellDoWMO9pOZBHwmKRM2wWm
XGRxJHTFJPkzQ1Qmg1VE6MGE+5mlCCcc+tDKOlVuh/uXjpVCozTZpJzoMV6rAdGK
yDldhzmb1N+08xuAE45bmMvOx1u7PDUSyKNMYIpgDvh5WwCKPmiO28H3s/ZYmWs9
ubXIaUiuh6VxgQuuaWkiyU2ssqmMQYtnyHfGmXW8hgnM71cpA7BiW2jpUl40MNUz
nnSWYJDMgubi20hRYaS5zWvrMXZJkNNtbVV9IROTT+N/OWOqOJEpUjCJb1z0bOHk
/GDSbcu1KSHsSeW3cNrCIk2bL9aK6+KeCfj+E50sk4LZuD9JrOTboZ1rtTprbztT
UtzgfqKRgh0CCfuwYnzfuLZUbX6n1AA+QGUzlFGyfAH1HgXXc0HZtwS5bClnVMv6
l3aAVzjU9L8xpsPMqtt5Ob0K6N1/NvbhsyJxB7Mp5BijGJ8J08C7wc9GGMI4z2Di
sR0tylvCykEEGXhu/x5f3XvEAZF0iE+ag5b2d3FmnX5alzloqhGNd+UznuzSUVqK
/5HQBAW4t3d1mR0E52K6sezrFXkTct7Ko3h4J/pcWuZ25l03tJRwBKAwhCLEGYoS
LECnOJ0TEJFT08S3nD755iEATkZr7JMUjjDJzslNwDT6xUjuJBEZQay0y6aULCDP
HUIxeG+XfqKE/Iu1oxwdzq0XeIhEM9pC3BReacHJ6kJs46Szt2SEqyxFj/1Gk0Y/
J5UKMF7L3uKQxn8hNgDnSKd+LMSCxuz463k4mu7Mjh8URQg64p1TKhkyaj0vTpTE
lEw8VLmeiWSctNcCne5oklWQ9yDNALyQAjxQNrwHoAgP8daByQFfDEOG01DvVaAr
f7a4NQhDGMj5iYueGyCPWjKzTkhLWX2u655cKM2XnRlS9ZnD/P2did4CO0ugGfVj
Nt5m9MaZXKniIoS7cIYy96LpQ1Lol3oXceJniBk8TR+/XTrW5/BQb9/NgO7Fvgdv
JIXXGmCVJwcstl6nYzd2O1gRb8olLGjfRg6Kstqx2kScNGMkgu++Zlh4U0OwLeyu
sxmkyT0mUHiVYd3fV7xCwoIn3cdBbwukRrYGC5RwhnT9vuyU8f5xIKuLyLAmZs3j
+51Abmk2fGLteDuTrNCs+tekPtRvoy/UdR38DhesOW89vWAV5KCdD5Z9chPzsR9i
qdOvZWJC3zf14jluYt6r8otb3fe1OA4OVY1atbu5K9CdUzviGxdMnxWeKInyOpni
+NwGXtIJKf83eTjGwCz+lVqhvHRedHCyZz0Ztv09UBqveSewzYh7COFcWPIU45K+
jC8e2rvTgVGXT30VlANon0HIutwNrn6ymhYG9tx0poh4Hy2vN7YuW/HTPRtf4Vdq
U+PhKFM2V58FGj55dCK9wIkQTggqPtP8tmdgqWlgOJuaxZbu5TRqJPTHUHXWjlhz
QloWAjFezeRXl3ycTEOf79LUAspntvl6qdSkyJ0vvvsA/PVDAivsNGFvv6jOH9mA
NuIwjwOtHxTAtsZm6KYSvb4Jagjk0IsyuVizUj8vAHt0kdAD3lUNThIIeXuz0ZPu
Ibr/X1x045/ih1fSt+mB8JDAyDdsi28JZFb8U9GiBkz5WCxcbnW+wROXjXSM4XCO
mdpXz3CuZcVyHPH/34PAAy81gK9ARIR6RqUAX371rk/1y2tUKLhQ5LLWsY1WsOqJ
yKk07dIVPl8+6UrZgPl90k4AHwzwonzQlJreWw59CorRcmnPL+pzTIQh9M2iJSOC
j8h3niIHYFHYaLNq5KKaYGlui29OEFaYmOu2lXOgEZekTHcWFGvju/nr//mNEFFm
vvNVeUITBa1V17sXRY74o9n5qz53Nv1x2wPk/btkTEQd5i3ZKp0SSqqh7y4lbM5i
kw0FY5xd90gJLP8yui7eg6tI+Sf6XfM52XEUDxGMlNLwTWsnHdH5Aw4vvhhtWH3b
xCPBT+a+463wZ4zi7p8AOaT6R9eTsSf0AFZI6Ekb/JI+TzLyvMAGshXLGa58XqQq
SHmrjSVByZTBNORulpaKZmMrisHrowh9Gb78hRBfvh/YNIT60Ef5caTCQcd62CnM
cBG1Nn1cfTrOUFl7PdvCEJIcSXRsIV5vUHMaIp4ts9J0rOFRBmZxz9JOkUKjL4+g
RnMMVAMPzaMtdBhK53KPx5etR+NcsdBgYUeFLx/sCaQarEJk7HHFZp7tQPqVeBK8
7hIgR1Hp/yjYDhw3fDRqZIRuhdb2gp+FsPr7yAg0Xhm0k65q/WtIqRealdIc3LtB
bgPrlnSEBEQ+cGxYjllRj4Ib5/uFpq8NgG3f5ZE2+zHbGmTNvtld3y8fK/bLrrjt
NvfX86f3dA6Tjpt6fSm160ekGF3ltfu2uyR7tpTiLaYuqhIz7bniqEAKn6jEHpKE
hgM14kAys2KUt1rrHlcO+UlmqMwDuIN2iGE0OPVoxpqQmrgVmvbxGXA/6c0U4FBb
Rvcu894xJ60sKVlvRH/DURuTq1QTo3OuLbl6KtGU3FbssPkLBcOOFErtfrecHr5J
6JlTXay42qQF4bn5Lr5ykBRrGSu/NP6e62sDboHpyzUOoDeDT4FVloMOAjULRqgr
WEb2GgpGLUqsQjU2s7KlNdH3REei31xkMtBksZypbw4VkEJv1FsyP+9sGkSWq4DR
NpMthLmWo3xBQTbfRllg5RQP32O/+RkLNGXf8lbhZQULQXX6WAQxSx6kAO4Jhc9S
xs6d/JT8C1VtDqi2LDVIMGpSeonHROqbEV8sfO1Yrpvfu3DI2pjyX2GytVOvzf9v
1jZJ0vFUDcsPfBSXZAgItpf625hj82FLyQde/oFoi/0PVj8Uw2/5Z4MN7og3EhcG
RJ/JnXJIcrZibay92r0uKJuBEihRH2Qjtyx4yuQyLM9B5K7TWTYmj3Z6yeWLw6Fj
w445gjHU8dDkIb8hqHENoYSm8q8VU1YZIKlOqfq+1VGQsdYceAVvdwNYMOlj26LN
zui1aE6QLcFlRFbtoSGYUAtPw/SI42cD+yH+v/Dx+YrNgXhPB/79C/gd1xfOpn2c
9l4utyK3rXMZFDmYl9/Wd9PEk5Y8cO31dfE8ps6vQetgQxb2MP0WyUNdzazuUNJq
OZedSfqFRLlzvQiT31Bcc4JfU43SzsSxCit9O27/B4OuJOZ9NvINGVsISxxadRDo
PR1MSvxXIRwgC7Wr2m6bEijtgk62fhNSH92kyC3kmaB6xgzD5S5RSwmf0W5+AjPl
xj9vVkRK8/i82qobVN2t8xUcpQtKx8IbTy2YsZLT0oN5YccIM35I+NYRleI+4/p4
z0BJskERncQIeujacySjc9y1omlNRyAz6JbreGGRFNXoj5B/FLmT3PXGS6rVFdv7
ZoCi+rg2vl9rgO/xOCSlK8gV/oajvCuIqf//DyFOCwf3R5gTdIGTZfeljVE89ZWb
pIl4VHq3pOlehkPS4Dez2MKcBJed58RjbGC80mcaCeod8H+IvFtyQO+BjKQ9Pm6t
I9MLi6DyT7UOyBW84/3wtWr00dxVW8jeViEU6K0jGJaF+lu98jA/OC2B0V254P9s
medpfTfSrDPmI7JMLd3mKtxwfTS24Fam2j6tMGv/CoV0y2ueIDrSJMpKA7mW8JB5
AI87yzM561pm3I/Vfk0HIZHT2h7PUKzkCMmb39v0M5yc44zhkYT90z+n5DsJqgyl
cEZWTdIJD7nDae4n1tMnjpv6xufTjB0+of14DSi/xfWy6wDlDsOc1NIDxzYNK+y9
NkUa1R2lj1P5HvnEGTNhsJZwR0PnleQZAFnY6e8XlKrwUEsJhq2+OAKqT01xBHrM
mQmnVcCbZ6ye8hcdO7a6U1Nh2dLQizqIwMvq0OIuCPsZCw8DprU8f1ZmG069vtzI
BkLDiTkjgiAfvastftUXiC7I3JeU2zCEBrsuzbqbR+0j3vCF14EGOvy05ueoReFE
DkiE+f+Vrxi/7VBbNONGdX5rtdJC9A0jR4GrvyHCl6X0fNI0SyqmE42yIf+a9jOs
s6oLyT+5JzKUoJfsGphMUeIjexoHMpRxGkJoGMroLT8p75ryB+rLBqzeMcAGO40b
ZGX8Z8jJBrGQsopfY+5/swdOW14OQfb6TCGQJ+/Ssy/qbkESPSxUMy0njtFjJD1v
P+LM9+l0R+QIlwWrGTGve/fZUYHMnxsEw4Vew3/BCa12I4WWjO2Uy8kzxp1UUsfB
HWBYgXOs6+3X8EcacucWbysVw6A95j4FDXaIxGUjX1kyyGvOLqnHlrEN+P9aNte6
+B6oXrsrqs7bA0DCTp3zIY8H72AkHw5rYhmC8paJpADU/hVG03+X3ii1nU20dss/
q6wdObcFIHTpfzYtpP30rb0eel40L8EEdUACpOKlNIm6aReyMWQ5Xe8OAoZp6vHi
Qy42sGrp2Mxh0dESK62GCnxfZh0RxDhy4KaaB2fNUr06DLaxm40NqOyCM9q8iyqr
h60WUnrjEAN11yLMCtvrw83VjMJPbUDgAou32NOsfTYrZQ8Ea8cMvgHthcW6tefH
TFVudT9opPUGPr8LAmBgzeFkakjgzBVvtBxOlI/ziFtZ8WoaaIoOMEvV/PNOTJie
qHiQfHSLkDz2BEB816F/i4HMSnLdxU2MU2OGITl2OUbGCkvM6MdU5OLQ35HROr82
WhnZiMyobKQV5XaLoCZ4uA4ik2x0DuuZF0XBwmw77UDPi1Qyi3ddsv3yUrAfkcsG
DZtU8+cvpBAd6YcaFEli/fSF8BSO+F+ymUvn0Rq4CV4KiLC7rAOqkX33+7kDBG+M
bClik6PVNqzzMoig6lvEgHqj7EM7zpLj3nSf6v/JqjJq5xKPRLNVb9YlFUvfttT5
RC6qJ0BadydjBP96Nb6hwJtXh54v5OXZyXUF2rBIImy5s4y+tjhc1+91mNGu6HDE
OI0eAbB8zyKEMN1a3SdSlu0i5eh8Z1CGk88/bDktfu8G+9NulQY9fYnzAg2loyFE
TYaWL1qRXGCMK23g3bMAiG+VgBQTQC5FhTCJlEDzKZNobeMVEWe9RhBZtPQoDGRz
2+SgW3VGTg0f+tUzORHssfLFFvfNxTn/LM+9OpsDxgbZBXRPKK/ERVwRk68oVPV0
tmZMXc6Idzs3lVLNlK/HPmZoUtoVwLWDFqlMVBcvXZwLbGza3ORE8r3mSU254DOs
Vn/6GaU1RCU1BzMJfGvEHVoUlIzUMk/usGpMXypLN9oYfxyNIWMyjRiF9mFBEaMP
7k3KBjlE8BxfmfaL22/Ow7Ih0yamZo1qku/tY4oDl86ffbLX3P3S/vQCv0IMKaJb
agM8bx1xmIuyJpfxT4goiB0OiLXyCRCAyyfZ/UzTuvSzFm8n7ubpoE1P6acyZCxJ
2nmYUsIIJkq7xcF36Jy8R8fBc8VIJOKA0MnLdbTbQv213tSSFIgp4Pyzk8e3rJ9E
ySLepdoCv+Q8Zk5PdcP/Cr1WcyAPvkpGm5tpg4EBmh4W+bOhAttYyXR26UxT8NOR
PrYq7qrugu3cYNgH+tg5eluM6+WrDyjL9clhKbhGlGVOvX1QBVbpHR3Peqx/Swff
G02y+czgP2tDBEwdvBdIlgCokQjc6zPnK9p+pRpsdQCXo9MggbPA4oMwvj6ZudTK
xOv2jZYCIScRT1WSUZe7ttrurNzXCj3uhXMSW+KVPRh+JahwtVFNvzttFXFQKZqO
E8EQHcxbG91awQz4+uKjzoQKyMlPUqYI7YNFxQS8hrQ+Wqig5gg4x7kMkwda0u7v
Ogpl74RjOVKXbL9QHDkoTcflhpXvXoQjJwvPgv4t3eNXSH8E2Du9mPAr7MBibkjX
Q+g1O/gJfBXv7J5fQtNXBk12mRodUCY1wc074zgP46l4gsaft+OHI3Y0I25/XxxX
RYrEyyNucHt/kQsF3ZAaX3v2Y9eaIpMvL2OUHkGjc35jZeraFPPgJEwDW4TCrNsF
2T24YjtxX7ZRxfVCmtl5RX0ubeV8uBfDwvft5PhobZ6UApIT++PTJ08yKG3CNdeq
esCdmOkDd7i/QzpEBjhah6VwY2TYowkHfEjRI9k1qyUHmGDMYuKlC3FCX8JWYEjg
R7mtNaUh0mI0BQfk336WhxmIkc1zML+nPxt6BmrqNc8FvvbJVxNLnVyvgDxDyPkW
EVguMT6Psarx/9Jf4752FTXJko5f/U2h+c3F8ZbMJMinGwXUX21PZEEJET/eOSdB
4DQsnPKRUCw/ibUVJRczacZPqKj6fr9vzdJOz3VUgsyw4RBL/3vq6ArK9oucfnto
X0CfCqDCsZX7j4hEHK6OncGrNERYrHL7UxWotvLnWszIgApavs0uxkKP60NmumUA
jlLMlhKIEP4tEDEPSYUpAaGHesQEX84kFat/ItqN44MNy9CnpXvFiu9alwRcN0l+
RdDvszjbDqw8Ik+xazCCoBd4jI7F9JI9YntRHLahqufv+BjodRAF1pJapWvmVwHx
8DMbNbTUjH1aGFjQnXblNwHbdrqVTWhgP2r+oV2UTNaejevUc0GHko9g+tvNxX1u
SYs9+8Fj9zG52t+nXDS1cQkJUHnYAeFBlS7KgSY25uJjHA/05BN1ivdJB5XKTpo6
ay9CvQrIhVGLZ5iak8n3z0EnvmcXZyyFdjRPDQHNkAxnk27vl2+m0u9EYzXoSqvF
nAxIUv6IRF62b5BNipwQpOQs2qARSM9l+toxPtz0OGD1xqf7bZOrq6wSqV+rTEua
5WzKyBxJ2EQ2uDfTScIhOHHITCVC9FE7VlxrDNWI93zJLiA4M6IiDSuRKD6Exuqq
kbmvUTmoTFW7lR6elQIF1fIDvrK/ApjLWPSqK+Z3FJ3rtg4kB1N3irQVKjUJ5Yw1
nFd6ph/kmRlKjxmyV1uxTkFUjCxYzFMQei6XVgaIZpLMRW2hpkvBnSWTxjaMGXOu
aJyZJMKEAMb+3YDrwRbh2yBsK0n8/Z0ScKrIafJzI1pLtelekvHbLuEYv+5pI6uz
J1NzkbYKHTR1bqs2nWaMSwtcbqOuT+1e2J+5/rt9UKh16Q2MTSZaI79iqsOZ6luC
6zwJgd7xuez22H1qKU4Zj5dSkGNMN081wLyRR1yyKeOgz4Z8GTmY5y0rNBuPaNvx
pNRJqEyB5L54bJQmsw95yNNjBt76sFuTxoip+S3Ys4Dwj2kJ+Kyd/PU4T9UeBfC1
FdecVy/4FQx6ieS3sz0rSn70eJ33tYvQ3EnBXMVCTrumxQXgKKe8AYJYDkZewTYo
xm9pC1uBz6cB7Coaipi3oguLnAR7+EchoJ96xmD+Pug4qFj7KZrJ0RzQYYqi95TD
TdViFkmfSDgkV3tiFF7Yq/pHBOY5ER5AQj16QCuFy5PuafX2su80JzZrZ0GcPZat
+SUM2Q60KAwzENsVZBBnYqQ3xe52vhUCkYnGG7Id/rhXC/vgyNYU9zmKahATFIeU
duj1rtQ8O+G1gT/J5WHDfPHicEufZ69wH1pRkx2Q4xv2qhQ+jCheT96DpSoV4Cca
NGmFZ+IPTQEZDpyX0wiKi37WF5R8SScUazhdyJqzMOUfMGYrrQKLc6l64KJVmv5e
/STmD0bsVv1WPulqvsb0YRNPQ607hSnHwcBXoxmgFKh1jPAB56ZKBcNn9Mc41W0Z
5u/6sTSI4JPiPNPj/b2+masIUqvV9o9TDQWeYSxzNSdDX+uOeGtGfHg8hZY8bDjN
0RSL1nUn5nQpS9UI2zvlTDVxJS45CdJuSb7QvaCwgd/AnGr0t954wSb6MKok0Eha
C1ryqnhLS5QK3fK3xkJcwfK0T7RXfsQ0l4Qjde7H063Zn6eJnFfma7oInJJ5OKXv
wujHcaTGkUz08nG0qwzwlSadtXN/BJYIdJJxCShhxzvHhWJ0Cv1p+a9kk0seNLp7
g1T2VJsL5mcHtWc9szVcTbQCdRR7IZJjY1KqW68FzAtUabmjgg5ul873tfkFrX1U
11RyyarbB/r+dqVQtC0l6T8LU+mLUXt9BDOLPm8KgQ2PXwxsVn7RbUguF0S7+KaN
scy1CXCQyVOxi8g191qNJ8x01TC7/5G992pnPSquMoHIBuLdf7EpHCwdW/9J9vlF
RQ9tB421fyEKctU3t+NuTM12sNP/UPK4Sry8Yc3ExSxQ1r3I/l7KQr+8uocPloTz
pymx3JA69yozpTmOCJxou/o5YPLPweuGOJAaaUFWz5eyraNRqyARIpz7Iab61nCv
fLRSwjvhg84D5NuLa4Cu0eRd9+KMFHmClpIqOXq8wBmJUOUbcRB6ngCfxWIBQ621
TWChJcsB7qtfvgkoC3Or1ef+5c895TtlhYaKUoVMbuxQqkZB3/iKJdVrxlWykoK/
8fSvqtzpBJUUIW2PlYIT0cJVZ6JvUUxz4eR1Py1VrmvqA8vFGKEaz6tJ7Wr41hx4
5vJN+IWrlKaZCWKjDakXZUxaj3iyQZ0FLl09ARgcv9F1pk4dt05y9NQQ1UPVx5qY
ilpW6FS5rCB4HuYKs9FyGFjGxUXPSp9MwGCZIfe/Qm295v3XTSTqGwwJQjQzqcV+
UbSJNylAP4/rUDcEGQfEb0Mlic5yKU4WZ/DjmB7bqupynKoqqgGjhIjXqKQBPGoC
ukm7RXwpKt3/TsD8H9FdEOnB1k4LBoYaEzIgw8WPwJqzIWX68TOP0mZ4+oVjdMRO
ltwDtaZkh2nh8BjYxPVO+tl0rKQvEm4672AlhHdQsZXuUeOWHUeW5RO3shZFZuNa
1mafu5+7w/fAlBM1BG1c6pieG1YiLiFJdr503Fwik1WlDQ8mopmUx733qG/slFbs
fYf8MtwSk7zhr7zOLJmzMDdb007TaE5RdYnEL/HUf00vj5EBSA+W8visqqn0P9VX
lBuSyi3iboZpkF7x6nv5LSryh9K81cCDilpi3vQsgW2D+AsBxXlyOK8GCdNKdvs7
mNEF3CIp2pmzG8NpKkz6Zz0gTWnBWWU16R6I37uk8ESHg7e2U6mIcde+/1LofCd7
yhOuAUFM5+QbPaBHoOj0OrmI3IPrCNrU9dme/Hp2o6x2Akx89Az3teEVZ07caYA9
uFmok1SY0UGIZjoJqAKOxHR6yIhI1pBPmiOs70+C/uOhmOVbDdSCXsdBXY8Nff9i
j8qiTtfA5pfvhXl5sNeg2ABLpWhOT1OejsQCMn3viiJ4jeNS0S4MsTzv+uPwfkC6
qnA7sP5hDiR1Sk1DgiYWmSxCGxJditS9laoK9soAo/JfFl1HxkxvCRW+cXUebaqi
THhSg+b77vud/lxFQKdtB4il/R8Dmu0kMhpr8RGlMyMhPvg5+fJdAUO/3y5z5M54
QtadVqpRfnvXI/O6RI/cOVo+gXbFGik2Im3sIh1g2PBiseV7D8zMBg5HLs5BFyEO
xefHdG+788khew8kB1RuzE+XHNw6MDkNYNsHiCAyTwIkITMJnx0zKZmdNzc7fIOy
IzmKFjKd/h+IWwinSID+k6ga44zf17gHprz4XXbU3ZF8u3X2YIhRfPmJdmwYvJqD
hGTz9ovSQhYmvuwNs4CJcDOgK8WGEQy4vOW2WwPCaeyiKUKKekzc5SS0Qeyahc3E
aUjqzfk41b0zxkFKx/ytXfx3ShM8A6Xq6ysXY3M07aZ5XHyMLGQ2oClp/8+iiZNM
PST/e3ahhzteSM8ZBNzU4f9z1eVTKaDY8CVYkiJ0QWdKFkXOJXaftF8huR4sLjZo
w2NemycpJ+1aFM9GGDe4CmK/LNOt8HKS7Lur4E5HcXY72hPMdhGZLIGen5nZgGli
ehvHoPS2/RoGpaGPgl1PToChiwhm/BIBCyzxDcLcIr9deOHeAq9rjQljSVOoWDqm
Nu6tbCCgWUTu3Ibn5sfjzRyXMGJMj2rkmjEQQkm0o81zM4xBN0xWOjfgAK9LTwXm
sBN4crdYPHUlIvVOp/dagOdZ4/avMeejZtgFbUa1WQFfXWdM0FEcWWkHQN4dunmS
Vv9j83s4NGpw2PG6UzrKig28+wKaF/Mcz/QkQGP58OzP1SfCX/ogEibi2JJ1F+wA
qysMHzWaxSY/HFBzTPPKukneoal9DfcErR53ebtmartJ3fvygNp5lA44xk7ouXjq
L4qohwXX4dY1TgTT9t8XKHxmtHn3DxSkK8pcwQnoK1SJRQFnSCgHRCYBoucyQJsY
6nY3wRISCv2cpMf871s00G3eCGkXbUZxgZUfJ6xKzXX2gFUlFGyTurGlv0Wi4I1z
KFbbxb2s8YLACe2Z9sejqRLgilvjhjOitLHXs3kQfRMzP84fHmbfbJ9vO4fJSucF
tblt2uIjwymU8Wr0X05p9yXrhBVEhpxtHmu85Q9zvBHhUvguT3O2fIeYwBsQSSdm
dqaR3JeEGQEMaMVy74xem/CzGzX8VZUaH2CnQVGj00Fp9Jk9vRm+TLKcddweEE7a
RuD7YW7mZoiXNkS42HyQEmGyEZ+cF//LX5FRCEqoo4FcI9jRBo2rRLp4yvHFz8SX
BMMOBHpkMAPuSYPpLczHLEM57ldTPnnqN0jKrptDD9pqKvEanQUXPIGhplwjqbT/
UkEz2OqwKMXjUZ6sug+VBzktW4Nm/jhfxzLakrkdu/3psBkTgg+FGRiY8fGkv3gX
E6Pss5Ht/VjsSL6zz1WgAD2/rRkbBVLf1Zc8QJ9RZJPCCOAdeLz3KcPPjsN7ttJe
4UxiTOsMhwYfKCF6BvgsFxtf4lCoDeF97/Zd/8Ytm1E6XGBnvjenJBBdswCli8fF
4cE5/anoQQ/uoHhgExFYoWuzOc48Ge3lPKfw/YLIgLiusuql+asFN/y/O+Kuj38n
BC1wL3FZyvkRhi59cFKCuqqtE5LhIOuqVKYaKr5gQRheZM9Y3zZn+tKuPbznVlhY
2iDEGEUkwg3KpAZRmolmWOanWCh0q0SEHagNqTXZs4kKdR1XYd4gBlfQY5c5UVkD
od8d+EfA69D3N5jk3f+znfSRLQWZiDZ3s9nx8pWEHydXCLP8ZHwSJQarVy1VRp2j
XSwhzzx//0GFCKyAeGhE5wgezFwwDHjd6X+huQppZc2CxIO7L3LdwtGVMmdBIi05
1tMkWTNQPbTeL0Mzcp33msWoT8IhX27Tpu8kvnQC22ciJCSPXaT/WjsR4v+o/AQ5
Tsn2ymi08OJt5J9nnchw8ptmi8QgstE6WlcsC6zpg/niXqPaqQ44VpEQBOTdp260
whPoU03gfus1Eh2ivzwtsiGNVcqIdnRVpyYRJ8xpaI+6G01Q7VZpueRR8J+Nd1CD
JZm1+A4GbC3S795lji3F4pLAXUxSDTpuXQWky06d7MKIbFbBzyBUR69dBoG5Jzcb
cYehQ3zph+TJiv145L1flPtqy2F7no3s0il5G2EVVASfSfv7qZlTdkrFdUcvSePD
j/N4KgzZh58Ek7a2r37ptyrU45GKr5oe0/9Ej0dhI+1MLD59k1jO+6oNvX6sCyy2
eJO9MXolg7rXSX0hPOi5Mft2vnFYpJf4SAzbyGxeWkhs1kCbaGdXF8YyMV9MuPGA
7WhEBxs6cOszfe9JFI6UCNYfVe7Gc48P8O/xnkr+98GlTzLG2bDAkB4qKzpsGLLU
ZHg3kOTxotYWrSurcu6R66oVxZNBEcoNZF7c9InoyXrgC6D6+P1A/ujX6KAVTZ3N
8V5vgSgNjSQWaZcli+TtrWOl6Rd0DIrfgjOOey6j3HdQg8xYrPx8QKH6jj82rULu
rvcuZYoaLB+HLWwjrLgi6ZIOGvHpAspAF7oqdd8Ubmc3LiiyYif7LBxzfokvismw
BLb4hKvJSBstyNussTJ4aJCIkVrNK1pKuCPdde6d2IdoCkj7S1MmyXLbzcmd2dn7
u5rp74AqIN8vseYMTeAwmvjhgRRG6qYHV5JT69ZMiEiL8aVAAsRPwDQ7h6PumDgW
oiltMnSMBMzHSO1S6rInGExdzlF1SHPmLEhv2YjD75CAdk3A6dyJQWmZZiw5VuP3
4dw/6yGy0HZuds1qUAHiA3sdjP4FWktUz69D+b/wt1eCENgtN1RR7IZElFWUCSLP
RB6ojMkSUBNcEJCEDv+N2sweee+midE2k2cKkA1QPALjxQ0CupsOsBcqTXu/hyK9
DCj5rL213399JFHEB6cPd0KxYCuzHse4uvEnK82gXfbprngGfEo+gQTKwTRrufGJ
ha2O6SgwCTQB+1nUDjAdlhZic64gQSwDbq5ROAesDQulN9CEZoiLvRCL/GG/YVC9
kB7RVPy2imZVaT0RCeya8lE2BOcRCoRA3mTR57ZX6BNZKaT1datJaacPsVmEfvPQ
bob3kYElXJRHfI4JMQ0y5sHf2ddDhKRb412k4YUnBxlhrF7i1uEXbLOrNrC+Xu/C
fSxK59ag4EzTk5rO19Fx9wz/KGQj1JzwowYq4lc+nM7J5ntM1UOTHQEoA/mgXuob
v2E2ZIwma1qMmAQ0bzfOiPNQlkyqvyDC4hkpGP2hAu1Q8Y7oTFT5bKvrxHoxahhD
9eSvdX4bNwIiVGz0vdKYmKzOtyCJ2IUnenleOipNnT5pA+Rgj26NjrBYJhYUdPjs
NVETksES7Fm3w9lDeg1ScFo2k4znNF91SJfHQiYfOIywnILhylNwN2fGBBqfoujX
As7mdc3pobKZs4UNgXVUSORpU3YgeSs8zy41+oo0xA2A4MB9QcsvU6Exun2QLFFo
Bj4qLkAtyOledlpmg0eYsRs/rJQ4R5A56/IAUON3PEmcqNZU5oOrP5cGQx6FlavN
w7CcYnMMmt4u9bG/MkZWbD/qDBEsWZnS0dMVz+RNnroXiNpEdjQEh6+2fsPCjnru
3Fg3S6oHyV4TgxPzi2+18nY64TuORWp3iOxLsrUEyJ9J/jeOYU/yvLIVHiQh2BBm
i8747GWAcwrFzHBuMlQOydxNDdSrnHa5ct2XchBA5YVlQ5ync0cQs/5M2rtVmttb
a/+f4AUqTANu0VdDLNd+VTOsTCfXOVazgsFipW8S1SpGnQ0eja5RqH1c/xM0HkqI
TMkUAMx0b3iAIW+xXRGIEO70RhN0ehFXgfMldE2oI6/vkn86/0nzxGhG5quWac2R
9HoGSgf3YwTjLigd2fRqekscs/oKyqXeHk0XPrFFVf1nGCqkisrJ5a4jyi2he+al
GrMpTdRgThpwtxe11sMpEftqXOGOdPhmYKKlVltl//BRQ6x9y8ofAaNKOn2wKXO0
6GpvuDGRzHGYBJ2NwmPq5eFPTIkK7I0MMdl5mDLxn1imhEAjVEcgpHF/pZNDo9rE
Q1ygULhfIFQdFyIDX0bCzbq3PPKqBDoUf5Oa/vr9eTTg2iY3MutDp5lOLYp3QuQk
zans+z8Wb552tFr51ud1wqIt9QtBk+9QND4hjE8U932EOR3VIZQeJGp+hK6AJiPE
Sd9Jym9LBonysaZA95EPRIq3UEMKhSK8wiXsI+FYlvsTIoE49/tYp76d7Hxlw6Vy
/+HtZk8hCrIYoIa0qnsiZVwdipa4qKpza9z5QW4hSfAqv1mCifgiXlGScoAjklfV
pZ2Uhgbb4JLVz9YOjo9Il3Vw/pWlorRmGrul9KkyifdSXzkSsepiksbzAU9pPefS
KkO/mMwyXV1fgW/m3p5RMgbvqoPRXDOvBKp7qyZhTF+0a7I2pOWp0I137V6Geg47
9oOvl/43uqknmTlOYJbM96ih8IihkZrGdxfOluYc2xGs00FbQPYHm2kc+zZqLxSL
wf5t4L2WUi+uSQ62uSVRZQThY22iGawRpBV1vy6NQjD2JOsWmtOD6FSGGtUjnCYQ
gVwIqBO/7fiOOVowwcOy8sXJ+d0KBDHA/zIa4rPQEg1kPQRiO/mqzmtg0Q6//Ggz
1Rqj9IPWR2haBS8sYXS63cidCfQLU9X0GakE8itexmETwnquwC++Kbmmqmo28+bs
3lFLZD9JNvzAN2reMmDwryCQ+bQOxirUv+9rgp/t7jcx8WkCa73J9J1k2N4pPXlb
tx5VzIbk0/3sZDOSb+9E3jB107p5u1nWE02cdwtAoG4xR2FH+rq9T2EHOg7GxZwY
KZpi8jOnJhxcGiT1v8iwCwfYQAU4zTeVrS7IKq72T0DrZjTJzAaV404KPzhGLuwj
vYf//HS2Qr4J5c7UmM6rBR0XRZ75VmzyNOYoFaHRwTVUEQTse9FQ+3c1r9tD+4x9
oYoywXobeHllIcB+hiCQvfwbktZy7wflp54DaJvmT1lUwRiWCUBj8dFl1m4xlTXj
Bq2k6y38FhAP6yjmUsEZw6bI6/Ot02Fl9ghumpUHGdrCLMa7W7Ez+yrsHqRnNhul
Na2eb2luEjm2ZQi4+Efrhn02YKAHl/RcQTYXZYlmF+TVfUr3bE6ywzboiLwVhCDe
/xUku2Wz5SNyjFrc2MfIeaCYkgKJd6xFsMjODbqnYGSS5DmffovYIYgffogX3Qit
ImeVSYjXG+wIW0wxVdmJc2JnPcQAXzoErHZSnqHPjj/LClWGW+eVEYPwOV7nmRWP
1X29DBZybrmW7rON7yQFsj9SWI0Kj58F2+0KrSO3YJDbyJtA3T3PLPlScyYe5NFH
yinDBIiEvZTj8OOt45VuUa2Af/sp8rxr4VfQiSed80YMTzjis+UG9xr9feiiDhO1
vjZIq55QmhrXhWKoIRKZyLb+rGIV/hB+UtdYISiF7n1WR5Lzld6qoFxI3D49syIO
OKW64eHxEX5TeTbmFGFM2Ddw+uRajcgUJ2EZhFxhqVSg9iALkRTFRCMnrMdpXyLR
zqKU2QnKutoL8DfIrlxmR4x1ts6sEGJrtbZz7Pa1/eDmpaVTANWztVmLNMyExUg7
iP965H74IYnMMMuTsSi4I4Sz+HMWhgu+aAPTVanEgPWyFrMYTBMtEuZaUO034YU/
6/J0CcKGPg/ilaqZ62C5NiaXsZvhxqQwrIn9983/8Jh1usdgY8skCJMQnqDm26uV
iZjFjX8qL+uiIiTseccHvJI8MEOeJFcdcxg5kArifav90pECIckLiviuflATNC9V
AWoAHki+u30/tuMv6fJSVjs6UbAA4OAkkO5y78CE2I4GrsoMMTHkRnnRS9s86cVc
5tRZB5ie5nk98Rjxm+YJ/IttLq3PdNaOMR5DtGpH56MZL0ihMWNwRShVoRPcxLip
fI5coH3bpCJ0dHR0HcCJ+U690IOfS4mMrr6QJDVuuh/LWzcRyl1ETUdm0lvA4U9O
LdNiIXKHoz+INVh7q0F7N39PLtsBx/AMD+dBVTaDQ41zhswZ0AwADVQH8fvU7d9w
gPabbjV6uXyLlS6/rV7BOYu+wRL77eNtoJ2EI+nlHirCMzWXNweIFppL/a3clr19
Euh5V6gjH3yWXY4i5g7h6BBi0uWH71XCvwehwz/s+3KZfh3QZex58PNvUkzVkBlk
9dgrcCaxnwJSlPKFya/P4De677FRG+E0LQTWUQD/fZOmjTWAqaynEfj+Mnr5V12G
jhfTteqdWhl2xrl3MOfJ+0sE33ZOqtcQgy3cyJi60JDgGJlGstAaIRjzdBMBcVGs
ASfBLQQPMdWP1+NyOucqqowbqyZcntOJ5bu28PVEYVCFgK/ymZdygqEA95uIROoe
6bqUFMg0sNDn+/AvYVfyGfyoYG9gfgj9muh/ldtl7k8hRBb2Uo09aA1Czk4uruM8
XnBu6QXu7JPK4oImetkky7CZYS4XZiFXnWK4bW6u2vXMJ7Xd2aRWoc0kJP6HEq+j
DH2FEw3GrN2oNVae2tEmIKYbmVcykApsyaD2fLK8Ye58d3QcT9oZ7PY3aJNQW/Fc
Wb1YA/6BloIhMWX2CGDOyDtNz4Qdujyqp0cpuJPIexYi6OKq3fgRRReK/zrdX0RB
YMg6Gw4SLHbkSDnpcbF6V8SABPl6FfmzobFYJAVIenQqRcmi19gvbRHyCJ70SPkK
uAfAUoj/f5zGTM/btXk82VUWEZ01SqjtJYYG4IYROaenOmG+M+AILFLm6EspofIC
Qn5Gi+8lKna3pk2uPgkh2FgG45dcklfuhlMgzwy7nHhY/Si2MjJuUg/sZVHDohIg
5HFnvP6My8esW1WOUAYsnfOds7LVh0v1l4RDmu+NxzyzyXHAEQkNZypcPUdhZ+uY
0HBas7GVE8XgA/1fZ2VFfRlyMw/jYS29iRrI6+0+eSnT54YjSkowNhRo2rSCUAhr
AgYLFEWa2K+2Y2iXt87IuDswlCw7Jx9C5q8gazW3L6I+1C5FEnBvaED0UAX3yED6
CznYtG59J2vrIVUdS17//SOOPFANyFEuRoDnk5cwNK8AMytG8sjoNVONOtwi5TAl
OE+2+e9ot5MRGZXW4eRp07kz8rkPtxL+oYJC/7Jpcc8jSaAi+rVe4a8a5j21RoMn
A1a0t1OB/HXwdBx1nBubb3ELgFN8D/11VRo3Lh3Ju6hi51/BsOKqb//vL5S9RFOe
JKtd2E9Ni+zmUxqdFuzaW6qfOYva6IOYDD2+Ct1Es9DRU6FUP6tKZ+04ZoPAmSnf
5Z6PMLJZK3hKXRmDrdXCqWiDwSRMASP6Yec2l0sYRANSk28qt/qjWXRlQ3pjZXvM
eXhTyLL+3ywt850Dm4/HwcQBSVqDAeVxihRhZAUVkmgKVSff++3SsKipMTC0fzUb
X38syRy5sa4fc5QGm/IOHPSS+L088peT0ylPvWB0mx4SEXlD+8Wh/XqpbvHH5f6E
VOPQWBsvL3lyGf4CocilYsrCkNLCWcU05N4CYTmSaRbLY5SGPZjDjR7Z9goKb9fK
O5OOIVamq/l9+vpFdbNecfjNMMUOH5a36rw2eGLdqCdNQS3hOg86NPky+FzEetP8
RudciU3/yj7RqtbWK8PaM9jsljKhjH5v7ef9syxGUTT3fBY3Ml19TNJ8BBDhG/mr
QgdUrPkUeDN5GELrv/yXcRMf7QWEVGi4YVciAuS8fNtrYk6E8x/wykdWe4EGWI9k
MYSoIEKwXwBoZoXsGcgEmQFA5j2IdqE92IBE/WXY+gNRMcrNJf6RUTJGGLoqGATs
OkI12iAF6Y9Cbt+EqfAq8d1u5j9JzUMDPpDaSnic/kmsjzEQpjuGQONa9hk3n3ny
OGRI2OMm7NlyYHKXPwpjmvidOOufiIadwOBH8oHR3IrdhfyNJBmiu3cLprYAqPLt
pYLGE9k50qns12XDiGeW0wqVlqOlyvES8LcJGZ1z5S8zxcUOFwhtpIIIQhhRMp0x
zCdF0Jzeh19HB5HoADfgXson0rWNf6MQKk/KcwKMnlH0/LHJmQPZLqpPQCxGTxJS
1MyZCXP0QiJh203Nf4cfvN/jtP4et/j5uRcS9K5+GdrSkRcXfUdUwiXPAxFkOfYn
w5G+NhDr2Q2FS19IMDa1dHcRa4TU6no0BGf2/Nn+Mimc/iOp2SjSle1KT+vTW3th
9445JKlFdS0bdYyqPEf76AMG2lbgqK1z8ZfogcnDJzDorPVxJcjcPOMYYmDVrNaE
Hlb5SSHmzPGxsTQe6wV2Ic4fB6qs0Vwyvb/oLBNMneD2sjja9sxNRFk+t8IVmRsz
8EWrLNScQs0f5XMMogikVaUu36Bvhrkh2ugFxwYAZf+8GN88u9vqjabdasMvmX1S
JVMJeJxsM1rfs4m1fAFLrgGOgsk8izcZP0OKBexnC33/HHUBQ9N6Crbior/NklZ6
Z65ahdVGJOydhU33025eBRGu0Hb4YN9CSSmoQLkeZTKhe2rVRRqu90TDcW815UPt
JOACrxlyYlv4jktTvAsKEjEKM8q7hvxnFnb0X2DgcmxHINMOFB8olJwTIbX7FjX3
GmcP1Khh6CkmmIM7Ip5N1ZGIqnPktWQGu4YuEhuKSWvCJLUt/srlE3eawDuAQdBa
XWB7nGmZP9N77cxE5TJhYVB2i7KRgZDcCSk5d0A9Z3CpWell2fLYnWctHEHWgC1b
Me9/jNX1yxniA/TT4UzQU1X5hG6JyqdQDfBHhXy3ZQUGeDhsVLkn5tjj1Mbvyr+1
66m6lFTnwUzeYuebC/Q+XNEA6aVzFzpIBahvf3E1H1avKgx831H6MnQYElGRQsw1
rcugGxCPoqERtZ8J5IKHWi1yhybl3YAEdr8F8hZffiT1gEGiZJN/uZK+Mpp/dCpX
8GW7ERPlpC9i+5WMNTjt6p7TJ8Uw2HersZFpfBcmEU2D/6iUlwXfLwZOxkzwPcoA
geHmEkqL2LqhhARr+rxh2ZPHm6OjZkt/elHCNJrj8w3bgeESVVMUz4IWYlx4g1z0
qObdaPZ21Qub4PZ31sFjHi2SV60klZs2bBdKvs9cyUnK50rmd81CUm2KZ/OVaCHv
RJ6kzohpI8FYPT5C2m9rRjzBeJfJZxjSgI6WpsJXsJ6R2avzYnKD9lQ9kwXQ73a1
UQecbS3sRQybN7OuWf5uNfnKaF4Idk7vr2k8f8GVIlbY70L5KBaJnLrODjYbncjX
zjylEMLV4JM6t9XBD9HO8b7H+Wpej4D08BkF1UEXTDOOu9jXJeM/9P1CuyAkAvMM
ci0NZYnKseBNQfCFZMEsBBDsnFWeUXXFDZ5eZuiWaKTcJjoUAtLf1+jRKAsxr9Od
WaoVCjJZ1ce21jBSbvE+Fo+IfH4RRJvsBlHp6vPvFPnyydS0J/pemZqW5xU9cf++
mmvoQvRQxsxwhav+5i+8DB1H4i+CJk4SxyQJdgBHJVi24xQA/EBl4JsF5Lk+4KPx
UsDJm/U4+uLTBIWtT19m4YLbz1Qb75UW1zVABG0R1yG+i3oWzc0vdQB/HWEVtc5l
yj4w85hHW324V6RVAge+hhWbAgxGrVHuLkvyExO7FmgI+93Oxy/QH/3Gt+nqDFdY
knqgzqt25PpTi6Xj4sB9Dr9jsR9d/SN/BQjFpz8szEQJrU+OkPDRFfwhD5iTmChO
p5t/gfjvewW4W7z6guGMC0pTESnMPG9lM++ErkFJt1uHr03CHNJHwbp+GOkzxAcj
rBmIUMRka5mBdChYq62+MsOz5Sc72nFnmy6kv0Q1VZau0DtMe08xloHIdy6BlysG
+8c5NwHjQXe1uCSDYeQo+6HfeqW2XGZ/ZavBEBstIJ6zVeR5oX2SDdf0MwLFTuIO
21Fj2zqORIgboUpe1IwheZmTkFIdT+McOYC+I0YbcKluGrHvP/yPwZXAj2A1Ykmf
dRfvTXaxcDBsiad2GzITSWIsZ4NfievdaXMeyQFxtqCXfiBR8eb8/77lPdX34byE
0zzzbGLptGEnjjR4Z2S7XsO6MvaS1wcgqldkOa17FeWIQTjxYaKpOHqb7lDC1geb
jRGaLR2lVf8dhkKuM5gl12tv9uvKT/KW+BXbURVmWqiIzFwE7T66FbBvzOhhIjx7
+jLhjlMJK0vAUZUd81vxdoaSqMshdK27mSK+SzFAIM9ObxtGscoT9rHCX/MqBo2V
3UUwrI5lThSou8FuhatmNztIHzg2wE3xNkihsYiFHyiKMKXiOrkXowm0pH/6i8kN
FTWllBnQw4B0bJJpPO0JUaqRaU/y+YHr7jvh00Z2XcnlDHMhowXx5Pdgmf4UUuvN
PE/Jz/EAjusmI6dccasoQ4/i6Yz+cL5KRifXE5d8P7xthgYA7bQnjqwjsiIKXcCR
oSph0VlEpx+OzbqDa1TjbLsekgYMkn1vngvkU0nhmAoe4xH9YiejTj9OOJ66Nw/l
z4O8sM6WP0PKSH8nImFDOwnBs9gBas9tPNecX1Jdlh5MvOubEn0YXbeNjnpj7gbf
WyYpA2xCifkDfh4wIp5Y5N7xOYZaxoO+csVKWA6dZiiuFXVVxmwPGqlU0co1dLjX
v7yqEk6iVEsPJY7mXu2890U9fMmgP27Yk31o6qCPVn9kAfEAHfXsmKAXhCI5BlCJ
jUMfxMiX/MG8KS4nJT7hMI5ulybnfmoiZ1kx/1iFBL428g8NQWthN5h63jWeycS9
VmoG+fiD49NqZRCk5+QmH3oah6pJoBvliPWB7I5Jf4TU3F/wIU93voW9bskPp39j
IQnet0VGrRdawlhesZoNHF7S+f8ce8K5Ef4s2DXcvxBVh0YZ5cYyopAE/nANf5jm
Z/NSREXuXmA7/6Fs0dhNepL+2JmInWBXFVebgxOrWC+JExwuLuRRAEPCV91H8zbK
1eFNpMgsUuvyI6ZEcIt5cu8MRNcnLb9l//W+RMmYB9Wfn4P9GXRdMtC5aEv7LZIF
lwc3l9nph8qz3fkJy5/V+CDsQHQyCnGCb6GJ6kYAMMaPgZvBDzKxHwSNaUV1g5aU
iB7qExU2L3Tp2VKQxX0OOhROLDqGx1kY7iuyYLsR6QhbjrNc7rnjR0L9zIbUVt5X
UNv+IGT1mRA2QSoDRRen8mcq6kRdmFGwIO4vfu3KeWi3JrTVci0lF+WJqIewUCLH
1/NLApPQr73l86rJBsPoRiXwLqMr4Yxmka34ic/YAZPkpsP0HLF5CFvv8ANckJfs
NXGDfLjHI3DInhG9/uHCG3HlYk5e+kKISkSAtTEnJqFaZ/OkD0BP7UcrBSv3y3pH
q0YpHch2p3Q0orxszWsi0FmwIzkWcbdKoTCS0cYxU0j0aA+LnA+IC+7M0FJ9W8KO
BCPcFPXo4IAYOKirB2fKaMAYSdJrpUSm9qG84Hn+uNmj85vkNNGwOVwkoan7XcPJ
CkMKgM2Jkr0gEr3k0IrPi3LylEbBGillgKTUl4gJAsX04+89oNrOGbWhKG11Qedm
4CGHNQjE+o7wTUBhY35kTUFP4OD2Ln2yCC6uknM/uD16JM7flZvn/uQIGbunUC4e
iezbznGEsPvZtqsdT3h9NODIixgYDSbSxP9oEO6/FG1tpvlZzDgCrYh4q61TuWmA
9XRs8cNK0u/j3SGVYADEaWbdW2lEFyR12b4t3pMGh7F3bwKmVljIa1IStzoGARa1
/42P/xZpMgM/yoORnvRNNnNayc2bsMdoSyxcBKyi3tm/3uVA95EVCFnfJwSYYu3z
oDNf/XE4LMfTYmSFnzVkscBEJIAY2BCELPGCpJb0OWUFitRKyYzw903vZyYlbl7h
eNHifGapb8rJ+MsUn8GaQ20owz+QzffXYZp+4Ty3cNegV76G9ms0F5w35OzybpJw
GJTKVfVZiGE6eC5LPqLOtldgMzwwq6o7kMG/g+7rdsp8C8JZoeA2Cd+o/omal/o9
GKZnaWQFvxPH6NCyDWaayXEA+0xMFVv+xR9HIv9oFrXVO2PGKNK2XxfeEjl+RiJA
IpfmKs2MiC/tXaHkVW30mPYuNNHG8fvVTXAKnDo+WDZAj7DI1wt5BTpXkuDXrR5u
vpisl5D24VJTqxVWNktSIMiyZyGYtBmpnRpDJ2Wbvht1AwEWZd5q2Qp/am30xlHR
brYBvyfFesL5l8ZnkZ9CmAzvBaGMnijaXbuYB8e3i8Eve06uP7MhLSoYTXyZY+i4
1vKlX/KHxwfWrlRuzFi7pwgr2Xa+05Kxxd71gZuIoUYM9HbfaP2zw3RBbc9nglGU
isfLByFf1p70hRZUstVka7EUf1/RHPk+6cxb+v7aCZ+zzQc+g18J1AiQ7V8q5uZk
vxECv65TNkQH+mLIpjINhpglVcVPYI6nLxBgU1XL4d43XGjojOl7FPahLoPgtAQ4
sITkK/+TlVEmTzZeLC2dKc+j+dMvXUmhd4p8KsnKj7tw5Qiyn1B6DO98qItunF14
E37MgEqZILI2iPuTaeHoVs0vc/eGgX8Qnzxgq1V5AS8Uxporr5tac5h58hekByvu
vDZVOaS/CTJYldyqPSBx85Vo2uO8hyl0ZaAoZDs0rlV0CUBTGB8Hr2Mh+W99ew+e
Tc3TfT4EEQ4AtQq8gZ+qGFA9TLClVXKrRS78257VOpCfWxAVxLj4/ne9eStv6l47
AlbuEPf+8ow9gHGS7Sju7EWb0K/KgWSeDG1KdQRfnQ4R2X0/qMZxglTnE9xse9Wk
DZyEUMpMPlDVCKM+M3jXtfSoZ088GwU1chYGOlYjV89J/38exGMg0AaIFhfpCWsg
iNlF+xzwQtfiqvJLKFgagEKVXJiffPvjagx09aWcObPT9mPNa93hGrgLSYU7P3au
duldoAnpxVAjPzJ80W8xQp3Qtv80O25G/gexd9yuWp8bieVDwKHIBM96liDsv9PP
+xpyV+OFiQolYMWfMsPmOSGubCkSl8Mss8mTNkX6JhxI0xUK4HjyAN5yn0cOKEF8
J9p05wf6klnR5ZtOHRXiJAQHq3Ne5SPTzbI77WLctgIl1NpVlD56SI7ZqkywAkr0
wQTVEjbx8M6Wn61b+0syvz7vdKd6E4l1nPL4lnTwB/A8OvK/6BeUBpS+RBkpg5F0
G65bitzLOgyxbHbm3/PPozlFf4YX8Vbo5f0GN4WdpaDbJzuzsUS4SOqQiuUIY1GH
B1K8Mp0fbVuYlKIUsnLaqWUIUbGxFBnziEC317GJLADcXI4VppalLYo5RmvT20mI
WV4yzhCqBzAgqbE3YI7P7Aeuw60rX+dKjgCvTiVv7BhwcTKNHkym8WD7tzCP5xHG
NDsJpNizyM4Up+bEGPSoMdibohZiPl6DpyyjBd0zhvVwXWGTBUt8SMhvxz8P54XY
8DyG4qnmakk0j5DOkGj4ljJHlqIYjbm/aSWBbDZ9QGVtCj5gu8/nM5VN9RKYmYBc
RiXo2JzZ6Z7XJJYr4njIPifhovFrDUVXegYkMC48JAN+/p3kYidhoE8R/jni5WqE
TTXSPerQXtgq2yhbb6OPxM//N/+/6RnvJ/702mLkYIBIenBL6iZgixBsa+NSBkw5
+DYxZUZmCtRR+1BOufp1a+x/ZGAMS1ol2o5YPsgyanDozzaD+8QJFHzrAwIyyUbS
+jXso/Fga94Cxts+nohKh7KvK0nzb67Nz352ZxBMsn8nDUIozr8AdbK/MWj7J0mo
HdO0W0g1634ffW+mmAyXfmuoECsERtecoi5rYSUQEeviKNuwH50mBVz5I4XOjZK8
+lvDcF8NJuTRErCgsdAlV3/GyDK0XEc5T6T5sllEK3N3JSraUK5a8F7vNOmK2kZy
r3+9FePQ4pbuqsS9zE8Fknfc2vjd1MVwCjsiQO9jlLM7oJmYiDirrttcyRKD1JzL
uCwBUVeI91lRQzw8mMHaasjvz94mveHUHfMoRRn8TSzCaetsETNTyBte/DAsL9Na
zdcFeJ58hfRlCzhwLfjF5u4wGIMgRJpyKhnlNO6EEdEtXhvABZU7a/IRsNGgqmqe
usO44CkOIx3R4E0SL+/UsHTP1GMlfIOwbFJYlTEOMMWQsi7awx0z4CL8Hj3D4sVP
l5rb40oEHutTN9HAqkgF7lgO+I385EIjiZ1Yr+oK7Q61BFsWDJWinQXnyvsff6Q+
51O12vMkzKonRB16fvMjxrHjJfzF2VS2vEmoeQSjV9CQjJk6DzWU4GsNWLkLSNbj
McHWkxne5Oi0P35HLUwCGvwTDOA46wWWu+YlxxbKM5z6yy6VjW7U1YBeSsVwntLu
lgzVZ9x/IBd5YurwFLpgrDVPy//mLxHQiKXjBM3Q/giJorwWKyhdpApNvXs+981E
8TFPC4ooUhs3oQdo/ZnOXyTp7XAJ5EVFhPL8PeP8Uq44XcLWFLAR/gKBemJlroYc
4Xg5zgHtaN9NTUxr/tnl7efSdy2eDCUk5S5b9fZI7JEYPq07tjczTagu3ps/iNlI
fGPl8Ui1GIgjRcBE9WQ21C+eeIlvkfN1iKVws/iK6KcDJ0ASEMKECX6ApmI4h/n3
2PR2ldoDPaKMKqEu5xBAFpJX9/EX8mfK3aCRYurVTZmG+QUMzw3gjdup3y68TkDM
OhecW6DgKATxMvuWPQaesfoL7hlObR2uR+QhdJlAh1djVuFdCkS8DLreB+boNS5j
wjxzqh7ug1QKkrMe22GdxkRbnc2GTzg1YRxbCvXhkh77T4xh4s6U9VYsQemqwOPe
62g8Jh6mVflzz3XNSDQz06Du1BULaIgr4eP+nFKZk0XZrwD76K3jetHF4EF2RhoY
UnIZqsFd2iAxsJLetWfYQAqE9Pv6yCnGBw5eQ0snRQ2QBMuy2DppZvC1sdZV3FxN
UXY291WXUbi7OD+WqJ7zPdB7ImxnZdCklLcdg4cC7R68nqVRUOHvDdeGOB0izz3b
Hx2zdtqeAY4uEUbeoWfSB8R7810YSHKgLfEE6aTZI5D9lq8dcK/M0BCBBjYt260K
lSz8OoUVAU0SJZo7M1KUeSoGp0CQgrnMXgyTpuH7hKhgAyQ99DvcQvpZaTC3+vPg
B6gRph8MwKfrudra7Hp1/JZE/4OLFw0DB+DCpsFLPj6sSfULrV14PwyZBi/A9DLL
66qKDZLAC2Q763aRjquYXh/Yl9jMJuzQXCqW1S94IkFwyLCAqzeofPv4gkRxTUqO
dt7W+AlaMuqrSIGRzjOLA89BgFTjNTpkuF1+ofR3CBs6UzWAiXDz/Q782uk0rzzD
53OFWwojYuP8lnXMBrlJKnumsqQO97pewIUnhFHenyOJxFoBY0lvzEuEsJtqqutb
Fn060WHWcJt7RM5+sZQVKeRcM+83pJqfe3SaJh1WXzUUFOqivUj5jZPLhwVwClTe
pQYKrX+/MzdA/MQk8zwInTXvo3Phck88Uc9gQXw6r8MVQDRiP95YJKK5mBiATQTC
6HLveICrLVOz67pAlAlS9zai7g3N/3tBBi5hKOvcXXaFuEDmw34jjEozY8gwdK+Z
OwzD3T8oq1Rp/Fmy6ssSj/m89YFBYZnzP/NH3yQzGofSrjKoNp1weKLXzz1r2+42
rF+US/lnrwvH8SAGROPaLxixd3v8pDdYy+JoTGRmfmrdm2sQ5mylTiw/xDfQf75u
7WYZfWzkgjosju3PLT3cmXI+K5NNV74DT9/VfTqcwhvSGh7HRA1FqqZPIa6exbHA
pVvGK1W5Ueqo8esOA/kJYenFFTfpG0I546NnVLSpCHjt+ObrkMA1RT1yjei1+1f0
JNyRpz/371aM/YqYjVDRuRYfGEkfo9Kj15BgrWNtrK57wCLglLx1fJU/jZcV9jaN
cGSMrES19EvQ1RX9CjhkEGkop/4ARS3ICpEc9wVEdm/rd5ZYB+dBC8lU8QdxsU9L
dam50nKqrgHfwOSOF188q4QRd3ZCCnxugkxgHrA/rlyNXQT6SXVNNhFesCx9NAvx
hmPJ+WJwMGw8PX0t1yfPtQVtsdb6T1ehKIciEKwtqMJ14hX7WeBFi1G3AjSiT9kg
RDJ/sEgsB4LOEwJrNktekez+lWBnKFC+l0zcyCB0yD6JtJugq88tYylvUnmt+VsN
tR3ocrVQ7y8/u8/tOjQVlAqv9SRJbZ250CuVXE8RToCW9310t8h+EyFH2jMcRduY
SlSkmxWAiXk+Y4FQj8zTDpzTaU0ARMLXfjYo9BVkdvwgM9ZctqXGwMS2unDNXPtN
BcfuHjG9T6ndi965KZhxrxuBaL0jC8mAZ8ri0tTdlwZJI16mAFbSaeO4K4us2Gc9
viBJyNXejj9cmYgdRbZyAhmJbpJQP6hQIFa59Q4UZjL85zAmyzKzCxGbQ70XDD/2
9UwInwoyqLQSp6mLWSM+eXYMv9RhgSqYuGn296yF2FLm7aFvur1NwrniqcZwxzqj
AAcTb6lZbx2xQKifiPysTwhK1KMh+UorWT+lU7tGg52xWGG1XBgubvECwL98rG5h
WjyVLsMXnhVD1VL7O8wpVjpLILN+dogbqqwlZnYsZbTvvudfXB5zrtt0JSeBCrrF
eYyoKfe9YzlHWPTKg0bCV2KYeDNmCKXTdl2JrZ8/T1WEYkQn87bAMTzOuwQhAk3m
s3LWiO0jinzcNx4Dg83gjlB7h2lpj/GrcTkjgEkKDaeRNtAJ6t3YhpPmWnhSy9jl
WOkr4hcknkM5BwY63V8BIykemLMrudNz9lQ318U+LWatgWWdXshM4a226Ey8NxiB
wG1EsnU1rsW+UzOpRV9rY/uY+IkfNVhc3hqRaoPR1HYcsTtR05xN0AoePS4n7oGh
apUtU/asFlOrY5yV71OLXWY2ESZRm1+XChMAIF/AWu1cIw9M7DPZmYVzHuXuRjCS
P+7Xoy9Vi7Vpc/8JC9QUkHnSH7MU6F6YhahwhNbsdhMFPddell3SIB2eCvMMY38a
Zohh2Ym/15aAEvJYmwWBhhSXnUowD09zk7aukxayP3J22bj7tVrPyM6o3Qsz8UXe
B0jeecku6CMVyxjDIZXz3BD/oZfmXSGulPO47EhRM0eAJHkYs/1cqOmaxNJGhk7O
93A1xdLQ7gtmdwPG7G7MPqfDlEtk0DDi9Yd6TYi/lgF/fySrjDsAT9hPWmjh6rx/
5/5MioIRw36yeeWG1yWLaLwkWZls+7qbx7txysXq45q/1L3OkrZdKWPHLeGZooRa
zGkhrs2VFCbofl0RUJg6NIVjfInK/0Zh3oIa6ew6ntEP7hxPT0MySCyvnAdUAPvk
6T+43/DbZPZIsFaUs47jgeBch+NPqBb/FRKKnUfPUppAWLdkDnoIby/exlI/FanL
Gontb1mxzPYE7z9Jd9sQx5R4JxwHFN0fjVoqHKN6G3CjRQ271FtF511UsYvwJYjW
f5KU4jyXWLXqQ/y2zUFFsay3k/xnOPdVfhE/kxdhDbox+h737j53scLdNy5IFGbu
ePBWHjoMJ3RtxxyX8O0fOZkb0GMRH8ULxqtWqfGGQHVZDF9eWZVK+HdXHjwrciME
hX5y/Iug2IA0pKKs7ziS1ceEg+teeIqwolhlrcobKqhY9GXVBdS65wBZwtc1mBJr
/k1sVkPa7AdMznej7RFgSCdABWsPfW5zhYeJTBouNECFwdIjbo3q1Wi0PJOtplSh
yj/Dil45PqZ+ZB7aCrrzxgQxbUZlq4e3/pSQInfUluK0iEmITlGcQ7rS2nsG3pTn
bDRNEoP8tFuICCDqDIOhmp+9vLPrwVdG0z9jo2YPkFHpIrS1Ybn2bdr3IAnEBEIc
nV7o0SeCC4LvPbfwd+Pt6eZ6GohyXI+enVomyYnDsvdzaE4mtZNDVaO8kfYIqkqv
63x+cBwmdMX9YS4SIp9/23JZ81caQWYuHFm0XFRbxKRw4n5XJa3m6fI9DTzZTENp
6R6bFf/ozB78XHRXJgi2tqszwEwbtw91t8nO9biL9m9nhDnh3NTbBb/cjz4fNwqC
wtRxFpCH7iB0nSZ8fo1E339JIrXloK4CuyQ35XeQgK8ZthUj6J6q8Hes453A2Nxv
h1cthoCt5tFI6gsn2kWo1LlnvspRC1Z/oziIa5s7w8PeehhDMbX6A8mV7oeSdNOU
oLlt5B1Cx7KVPY/dTOrP+cyw13IEa6B+A8i0j9vtzay2LCpXPS8Z6dJ77D/EQ7B+
NtYr9fS6HD2S4zmo9Zcpzv691ea8zu58Mmtvgnw7BrqwEW6nviXgr3t22Rp7JwqV
Zkw4/ymN3SVPPXX0XEvCryyJ15LMnO7kGGANNMQTDtR8Iq9S/GbDqImHRNGNLV03
9sQcUyMtsEDszkP23jeTGCj14TzPbhKpsN1urY8O3Mk3Uy+14Ell79ZGnBKbfMpD
uO35fa+GhhTIw+bfWBBkmWq/qOZBIIWVv1s60L1UaTMkWMNcvSK0A5+m1D/6vxtc
2l0JuoCSqjshjdmdqvTQL+N+CsVp94MQvZCzkq4erb4rDKsTWNlUESz0WOOSbudb
jn0mkoAWiz6aDYnyox0YVHnIZbzhEFOO1W4MU7SdjlluDvZSwDDjWvq5oEdy3jTJ
UXWL6HepOg51l6QudP2JyKvM28iWXOJx+Yr+CuqlBKmdWLqEk4WKrUZc2Yy/JJyy
8kQsZ7o3O3bvsxtaPYq8/rowwPqt2UZ3Y4ZVmbs3pEKsOKL09zm4A0j3rQrsiIgJ
VbkvaecCHVjLHcqwNyavgCoDFnxmcC16xShvUqmAMKVFEF4HEMTSbvIrFgenpttb
WDPProTioOVOORBYX8JsnmJIHkbmDITG763FY64wFaiT+bdD3DrEqTEoeMrYQMQR
Z1PjMOMni/cQw1MIAic+cKNKbMSA4IHy84zCChZHcm19LY9Ojeov26pOjjZRNY+h
Ow5Fqz1XNa8fYo7Ld0bVXpKQBZYwVsla+a3Yl24hhrCuR0S4c/6IxJbkIbN5R3Ci
bMMr1+LQlSBBucyG45mcwfwwhqiJe2YTs9snqhBb5ClxeunvX10cN2PGnp8QJoVy
uP6kl47a1OHLvSuIehFxmKFkLkkEe9gRrvzCvPt8MAofvGBIGyEs9/ftYMs40sIM
cB9rP9NZxkvEtF1PEKr2qRQ+7ec9oslCKiOxQ6yHNXNRnFIA+7MSZJVrOCKKDjBl
rFNUmmtPzZJhHVFM3l3LuZJ3RggA5WtLNCJ3r55PI8bZqHALJmAwQVvIXFLTE+g7
3Rx5Rx8KP2+945fgPJOQWaBJF4SztTgSQR7lmr6860t669/JKGcgt4m3paMsIY4s
vMx4nV1DZW/rCOVmdUIaSTcIXm6VWO7P/7DoS93GUmdKiS0TOX+1XIISZSvteOTO
faVHpNaoJ4eqKqsGbEfcKWqFzekYgcMm2E57+a0Xm6MT3zpWKh/hJv7faqFZ7dpf
5h0nNcaMW6r5gkvvGG+F2FJjki3PhWlD0qjkr0VBaNd6DyKvObFtOqO/f5nozJxu
oQeSQ2qJYfXKko4voJmFy55G42mNwUYt523MMkl6hrDI/ZrhC2Luz2s2fAFn0nCZ
mlyO2TcQ3jQ1WTNf1/9TgN74flxs4v8wNOqsKlICmnWafsf/qALfeACQVUdG180F
2wTYwjE3UE3yvUN+LhSwhBwZ/VLGJnXdPy+6ocsTW1Hx4NP4rZ2pPzhj3zSnrLfz
2e7KgY+hfJBrEfdFN6evjKTyqRfIkmKSvQNFbKnAcDodTi/fDACjPS9H7H5UlGcy
KPE1JBwCzFeRH78eeqjOjZqsFYsq20coG/cvwqJfnjyWnM42204XrE2Wpd3GBNJ8
AekoYbDMBUy4ggTxqKxz28FxNet1IbuhuC/GwwaGhtC7swioSAfoEtYbdT720anp
8Ku+hsNVi24WaxdgGPNt7RpbuAwvCzMbOg01tJNRzDNqUcnXAobcOpIFY5Hu9snq
nP+rbfcxpegHITVtnZ59icrnGUEGMpPjHDZfW3JhtsqqBOR+S+GmGR/4c62LCVlG
HjamxqDBMwR0V/t+Aa2HVTwvdF6ID6hmfx7mpBZiO/oiKHH8lBm/tFMJWgzMo7cn
hXiE3exunYnYUOqGn91GN38CVdjT3uaXKNour2ARo5RKLYAQbQ6ja9W9BAOVrjwk
Vrj2D5V3c4d1sPnsMi5UqmJx/NmJEkdMu0PJYp3WQ6stG/wEXw2g+eV8DMYwLaey
LhYdcwiJ9cSOYoGsg2925UrFlQY98vJXNvJvT1nVvAAe5IEP4nTf29X/7WJBIqZl
0MFxfEcSq9Mi/vq0akg88zQarEsggioeN6e9Yk3XL0nhXjAR7hmg7MN/Fm2PYVSq
6R0dzWbUYCxXkfOaR21RXh1SyEbVqZJ85bGPNjBiVpeYkVjVfBI1wEcpwn22nweh
dr2kmMiMrG1W+nK02fKCwdN2ntWMsAFUqtyc0KS5EO8ay0Gg+FlWt+Ia7gfVUfXi
CiREo6c4wZZOAbCHl/DD+f3c6M9K3RVQImKBCQWpwCJ94L+P5mkubXKmcMDgN9nk
PMxtqaD972KsbqAef8k3V20+UT9eOCJZ88Ny+ochhthb2cQNyXNjEHQw9o/FTzqe
Oxz3vWTDNgllj2elK3XIQdLSLEHHQAA46NJo8d4NTrGdNTIHhUvGeUqBiioHQPxU
YUNQcGpr/BMXl04TRarcysB+0+9NR2KRzXxVx4/fbYZyKMvXua3lkmAaDumMhnCU
6AVYmcRMbv+02ur2ERYYb/2eUs26Ywy0W8cfw76x4RJwOj6o4ulUhryNP1J+c6UL
AkV/H/L1f/Pu2qNmRUkBwDAUUjBuIIaxH8PWcKjZKc9jbQyeq8loyNAN5qWZKrg4
zJawZwwzqhqaMPPj3LD8eqW3EJ7upvQoK4feSqeBAwh4BuspJMAU275fEQQkQ+28
t0/qMG29YWzlqS5FfEvEZnK2EOAJ5DTr5bo3TqZpMkPC1s7s4Kn4ARoDlZcmCvFz
3kyGyMjNFwrhmAONmk8aMWuvpZMdYzAidLFlwj/p47K3wMixKVpSMNhCa3rjiyfX
jolTvRXy42dPylBTCD1JYnbQOsljavN+B3HzqhOhaxBkj6XZpFZL5cuSMiauUaB7
Di6Sg0Al4AJLk7PKnDHvV1DsNqm5MTheE2PlMW8MBohkIkdQ8umeLEEwtIeCj+Xp
qq5qDkQL5jhZZ1TArl9xFQm0QzWII285ZPynBLpMQojYk6jcxyzvGwLde3TZ/VPv
TdpQarEWpPW2L9JVDMWtOVcbHRrNQ92yqslaaClIIjEzY/8AsDlgMxVDLafC4kQ8
BoIjVrW9LxOqJPToqjAqmnSDX7Hv2KuP2yjG+nz20yhJHn0WAEez1XT1pyx7Lnub
8GsvrBAojOItbBANuwjgf+T5ftqpI8usYOX1J2pgyhBGjydXxtu901zhzUc+6Jik
65vBt4zVSGueGhPq0c5U20Xn2ddHDM8EFoopFJPVdD0eRlyyCBImb8E51YKuVCwA
TZf4BENpOUtZg/om8Ubud077BIx9xIc21Fx4o6SBSvMs41mmMKPNqT7P1xVfRE+m
9v6BTGCMZs9DytNbPmeChHNnSQaFqL6yYMlmoy4bYvg79M5g+zMOolcJVmpYkr0d
rZTj3XMoWbSj5RgoMZygQta9fAyVMRUqfCUrOBevyeR+0MEian6fv5RNVpZR/iAu
hM0QMueJas4cBipNpev4E67/d6SExGuvhK5cgd4uQRP1251wl/smuUV4bcVsT7sI
ahDgGnPqYJegp4Wn3Mf1a8HCST+eG6gGtU5MYECr75YtulKJQ3HfLmWQyAUa3F6d
g10pnNHppNKxdpUx52Szx1+GyYQONCUaIyUDWGQJGNIZdPTTzi5fak7Slnd+jiK7
9ZXaVT69wrmuYSWsVlaQxe0x1NHVaapQ86lkow0JeyMKJLu/fWv1j8a4rM93Y6nc
WLL8U8web5NXMia7K5VHhzUQ/csYry4JVNTBHz7Fs8oOskZbAqy8w7Qev5/HQg15
T0QD+7ckswPxAmCt3metiJMQrjCS+OK+pf43lYWG5kG7Kz9J7p/wqCYSIIex0UI2
+Mgt5xBtiTq6zxF/0eaSTHbwtl+iXRGP7ZIXNyjpYUgUXv79zsAfx3YJPyUg0aNV
C0+iId1mBlRoiPrwXRh3QVd6r2D0BdaIGSapbbKHUxew0BvQwE6seGIvijbO+hce
RVWCBK8iEhRQFd5QbSwDZ0G84gkljmyMbwsngCE2h1d4K8MLFmtTSd65cwhI7/d4
digtYnJlvRljdFieNQsYIVWw67g/Bt01+MZxC86z0vr68aPYZ5Jo7Ik/uPMc3ZDj
Bd2OW0AsrT/uuqZ1UrLDLCQkNkfagRndTaeYjDlKNJtLne27ugwT/R8MipWeJLAI
Z53x+4/Wd1dshIFwSynuBp9ZiRHSeMHiRSb4+9y/6CquQ7yOmc//9pMlMINvTaNl
Tf2E6I1LTPAdOjBri4pa7yJ1lP3nzU/lzV0SjJ1toa1JcSzYbaa9i26hEFYsqR5I
sFw7wMsPFXM/kj95RIJ5AhZuU0nkZhvj28tZLUtTYgTC9WiNB5wnHCiy9ULkPWWV
IcdPndi7DTbWKTPJ1NW1bVHMd1dxQmTaLeeEnX+C6xlrEzaR+kYx03gYtkD1NixI
evr55wa7xL1McN/pqM+BJT/pnTQ3FQDm+EoF/mlKcCcdbTw9PwcXhApjuX/0NfUc
H/JLo2LhTXYgar78H2f8TckivJu2CSKI4o0vP+n1BdMuEt+zz1dcDLN0dHio2fp1
Ucc3+Fqbw1isLTEHeoWCBC1fS5Jg7wH7ELSUwanRbHd4Lfb0ODH07rSOsg7UV0lO
ioYH3LvCoBu+H4O8DVrEp/jldCKz6CgXAlMEdztesR9iKUe+TZEEfR2FhlQS7B7c
BZ1bh2cHb3V69FrxaQs47VRB21bRzpUVpWV14WNB9kQc48o2oqfbF7uCTW4/dPXZ
AUnP5I/u/tIM8avld2Da5GF0bVP3JndENivO2EcfpDkNLIkh1RFDEtwnQIi3BHqp
H4ebWFA2rnC+Npi4coQoij1mLGGSG0qMPhRj6DRNJE4SfnU2unJt2kiE2WfpBskY
KktF7Vp5F+ems7gUvX7IAFUglz0ToVrMefSrc3d3x/bXhj4t/5igvEX79CdbLUXr
UqafXEnmFa2OwlsfednZVn/IfAFAHro2aKMFdRSRka/jDO4dIolofQpYtg9KKS5z
HyV2Lbes4yQM8CDiRBJQ49WF7zVdGCn+kgcR+DyFqmgJ+2/+CUXzWJo0qG5EGc5S
MLhYf9V6VgmMJapJ90KVSCJOyBRHSHhCerGq9y/dzlQU9L24sGVTcg/u8CsN10FV
NrWbpFr/xizZ5TIOhyBsnZ8+fYPkNu27cQOigIGLYYAlCcSX9lGv6sm06kWvjI8C
PDLts/gAv+SvF8FgPzNkz7rJYwwC0i8K+PF5Zh7f8ge+/grWYVtvidSUyeK7xwE4
7TYE9mQDkVz1GGQYzogL9EMACfiUkta3iskk/SSt5ImiFGaYugEjbAVPqMxZJaSO
dq4vBADlWZ3wasKqvX7a5/sEpkwMLIxa4CsbHEzyhWalP4kwARDcaize7StuctRo
r07kUBW7tFuYIlLzcxyJBuxCAFLpxpdAc1zxGLr074gKixWTWHuGIn4plrDz/B7n
Lqa/uJdt7TfnRSETBhIYM2AnGn8ko43s3CopjgopXqMrMOXk1qSWkkBZOdi6PtOA
2eksTlmWgL1QKF94kIDmZOQx066rR6G4V34NyAmOsfq88NaG937UFloE1+c4WmnS
CaxZL5cv7D3vNM+8tWh+VmV8T9HR3D/urdQIR+sCuYKbCfs0gdqHmtfvarpvsUl6
O3F27PIpP5cNY9+rgjYATqsZF+61iRYwp/x0K4QG/pHMKnbpDwnodt+yzJKHB4Yz
KPaxKV6bMCZ9pdOZk6uOznx2qKoyn79oEBsvhnZxYRf3l2mbTLsHK58ymFmkLPvz
DaFcB8xq+tbfDxHrbhwmK74FMv+B596WCObng59B8yTzcvch5Wtq1+OHj0zRU7ok
kYxcwppdYGy+hzHZS7kGJw/tzfWfmUqxpnikulfquOFHZ5wxT7NIq4Wbtz80O8yO
xjQhJ+RQp8qQzOChMrfRZkKG6uf+9cfBiqrWScuguOqqvjLug0/Xb2jnD26CqlGF
dDsbpBrpMr9Oi1vGaYpvLUfCtBpCHjP4EXVqdM8/fGkNS8OO4FTKklAmsLbPlPXn
UvwnHZjIvtbYIGE+mEoViL7J48Okbqu1a9bAmziye2xJ+elgXsal0JUN+TkO8ygR
42dCxBzkz+Iww6UDxTdGDbhnKOgU5BYLFJ7iPhrQlB1KoM7iR+7x176EG9OvL8Mv
EGXZ2ZCMR5hjHYuNyvqV1WSthCq+AdbD99taUAjLDYy3ectDOAU7GiO42hWWzaZK
uq6hRkm6IYwDtyNLIChvmt4BF8mUDHapQEep7kicXXOHhOCFBLqR1ZjSZFATjVzm
e03XIYIF6JnVYv2gyXLmToxEP1rm+zrlKf45AZvhIPwo3EshOoQ1o7jGlKmWo7vU
Rw20K/fcx77aotIvyPZa0p5Ccs2GcTkYGaJ65d+0thLn7lP4jce2s9rHHcu34zMs
rh/mWaiU22GdsktJr5YydZGDWOWYJki5e/tohS5Vy57eAKHZjllMGGqiznwh54Js
R7vLZuB6bQSu/2Epwg8TLKEz/2tQkFNrMfTU+DCuBT0kW35En9rnabU2Laxp8yCY
HEZ18IT8kQZtNt4TQ9xx5s/rpxqZUkeDhsCDaB3LKmSSFKlcKfARYTL3Yxxp5Prl
qsUAPMIUx0Ij6OAlCDgLchck4R/03zXYeOczw+Kc1mztX7jBNmSjvSCxF+57hhaB
jYow80JFGcDsvxzBToYi5qbQmOHzo1/cmvWABSNd3qQmKBsWT5ThrhJORK/aQIxZ
9KG3bwPPTSTqdFBanFzB0QoRmoKxL8OjxcdXvHh3GmIzhmdLKTdu7AhfXHSZGKMf
joiki+nUpdps9S9FT6H4f/IBd/MzXIjSwHlvZUTLGMQ3VnruLw0uJPSkvoe9ZnnJ
vb3mgp3MbbhaxsZLMNAWZE8Zx6xeqk2wnpRDBAOUeWfi8aIqMjZViD0AtY+hj3lT
K8n5danCOJFLGQg4FtthjKx05lNrtQRMRph1odDkRh/mfObghvWskCqy71Zdzxh8
AjuK4q3yrRpxqMgL4MhRpfjE5ClL0cxf2zAf4CYI/MIrKfByBWmLY+eEmAUkgerj
Qa7FPP7Mf1pnFWzHFfXIbLv6tZGxaC7y1Vw0oX1bOrTFYbn9/Sik3TzYO2Kq054L
myhAiN76CCdCHJP4gMUYq5ZAKNnPB8R2TuOfHq8EHsgufUZoRvpRCepRvloOM9FK
Pnv+N0fSJn/t05QQDc2KUQcgoiZtZoBbPv7PKLtGOyhneuzscurBp5irvAkB2dis
jSFFQscjjqJ+sq7y9puaQC/VajKcHbSuZs60KQ4zfomQBSL0A8R0nSzbSuq4oEVm
jEueVcPKA013EIqbuUDa4aYrzwQRDvWm4vVvzfUwWb90ubfxKoBhFRDjMSDizDs2
HcTky4tnr3S8bjMZFOrcYqGNzFu5zc8ce/0wDZNvnXNiwNj6sLZq86ZnW0ARyM9C
CIxgwtSgklYEzUpV4oWqMnRUmO1DnI9qp/ykv228SIykCdMeHOLGnItRepFQERQK
KpARoX5+Hl1VQ2zUeIsNOl/jMZbir0i0VFO4hWmWANpavEhp5ETnPx0W+uY6Nh6u
4TM3bX6SGxzsYPBXEWUJUiG+u0Syd94lmLTxyLDdTgkpfp7HaOmP4fY96bc/YtqU
08cSWdlm4WK5qYnEPiMzFUTt6eWgEBUEZff5d+FBhG6y24kjx8KR7EfqrGjAIJqJ
zIMF28b1lZSUaTKUuf35lV/p2XXqRqb0/ybWioG/UVASOIqL8XAmo7JprGt9y1oW
CY9YAgNhqB6o5WCi5xEdrME+x3KFQdbRyxXAc7eExoNg9ZMazVZr25DJvpQChNdQ
kKzxNCVSbpuEXJhlXH28pjGL7ltOF3PAA+7rBkraNbWsDwPpFpNRIj/H9zzx+l/a
EAPFZ+f2B6Ew/nGVutCOpN6Xn9uJiZKH/ydZc+vI+V8CjlCDcW/UxZs+9qJqEcd1
WpRZhAupifFcwgF8uoHE9Rw/DzFoEE4TE4eSMKvzzRtvyllo1B14brBg/FQs4xVm
TH6Ifby/vF+l3abUN7g4CAO31KHPhPaXb4J8ucEQnVGz7o4eTsnjEv6mhgINnKHA
k3xSQeCmzdL/LbZoQtu5TbAd4khtkmKhYFhzNUlWfZzJhrF3XfHTkV04+pIYwFUp
kwduLChuPqAVfdwjzn9QHZG7n61+IK+vYzOkYac560t8+3cWY8j326ImV45Kt5oo
xW2OrFwb0fQkpRAbLyVcKR4xQgeJYzaOozqiW4VJDWyOHkle0a4oOes/mD23mCW6
EjbzkQq+Cx7SztgaMJGTW74qy4xWO51kzlz7byzj1GFPWQFl2zS09fJnzy8vtVR6
WTJrUYcJz/TTdwy2a+IO3ni08uKl/uQmJYnXe/0cCNGZ7vD0M710GQgFW1Fci1vQ
kA0k90J/gu84aNLONEXow++o91fg96y88RmbhCFVqSZOOvcctwq4YFMS57JtYx9d
Z+xuXESeLDnGwfXFK40m1swysO05VktHi/AlFOrcb4rjGFM87Rs+BJdLMtDkHsD1
caJQtTMFuhfOVuHAqtxazRJG9hzvFgfA60KK4hnaFVguuY2zPcHRqRzj6DcNR/lM
TDKtJAbx/qETI7sdFTpO2OrWucsdYaC+L38HoOi6OVdl9ySVflWaN2cwjjY5Zidh
ghjFn8sYzzeozW9gMZL8ClTdMEjBi6rwTZbph+WOGe7o+PBnPKu82Pwx9Y8FKumg
TVIhlK74ZJesj2bnaf5WI4Abir3HTkgBYm4peCf+hh0ZZNY4fSXFKmzvgS2JR8EY
BIAmSXBBA+I/vdN9X0kMxJOHa8mqcbkkro9Vas1hhc6WmIH4/8PVM43xxoVrLsr1
xbb8oNo0z+eDpRwnzD9q6Wlu4r6/TPIPFJIjpeCFjtDxn0Ma12QiEICGxVVOIWcF
xxj7uAUoJ19o7eCB4+u0/gwgpf6PmJe+FkX//zM5qLvJONrcIddeTpA7dQu9hT+H
E11niyXVu+YjZyOMXuYHGOBPmMcceXtsp3spm/GRkBSSkvv0PrS6RGJXJUyJCEjx
tzVdAM/WYAYF7Ut4rhEEJXigJHXtynw2VGu9WusQ1pJ/gFZZRTEBH82GvloXzFbR
K8rdzCeGyiiWXEsP5H6GKHWdK+6HfqUyBhT14AijAvXf52FdjV0aU8igIr5cOPOF
U3+SCk9Pr0sEpoMWPcG4c4nLpV18TEKDww31Z0r3DFnaBuo1swcICm1mJ0a+DJZ2
Jur7+pyKv3EiPJvVM2Jxlqqj1CPqD4Ea17/6D6n/kBw+BENtugSYC+iU9cagVLtS
5PAFb0vCLhuYg/NPdE58gUv8N6J1LKsfvjAXEs2gZFiaHkCAuL2zciGLHSBU2MnG
NWgksCyuC2MIgBNvHzOGesc+bntpjijBV2Ka7LQ0FvTxWa0zJ5YjHBbrj23WkglI
OrW3whPJPFV9ClfAMTMkYTSlO3UGJZjOXcuA9nVClSwJCGNBz1+H8UydHNprHpJp
Nk2bXcwknTkxOTdlpGdlQRj8faFgFI9i0zpq+eEhXz5pKpTAliVp1lHFIEe3yrXI
sqDenWIQNVbc8gV+i1dK9YUAiOchkDUW15i3DWSwdqUAR4jTRJKSusUVo1bK+xA4
AD1X86JjAxvNHJPXtvKDQbZWT0ru9hZMJDp3Kr/k2DTecxFuMdQd/gh/DUq5NVTN
5u/v01RQSHaSLto2BncwXbsLd3IcuE3pKWwusGKM6dbYaZiBF09PdAHcd5hQwiTF
DGozCMiP7yBfxaZK8GGMLxrTU1jkk7GAS2Nn1SiiuV5n3iUJKqh4yoMD0JMUK+vt
vL/eMgS2azp3pJ+hzPFwJFAGJF1ZXlK5e+2ttePayau8293xtDLZ60o6q6NnpUSN
FqKvi24DVfbN1FzFu9OCsdfIlNqm7blhyI0pyao7B/IgBBpBL11HLW5rsSzogGqX
kZV1dhPClbi5k3DVawDpA7z+d+UH9JEXib5LW9YKkthE01gH4cnzEO82P2etTZPO
cWlnKXujRD38X5bSyc1QUJMIAXUiK0dM79JMQbrpT1pAN2hkDkDMskKE7TviSFpX
+mkDF+jerwSWDGxnP8uLSii7HuLO5aV+3lAYHloj1GaHW8zD3rRQtslGpeuPDdOt
8TQO/YnpwRe0Y1k2VVuX1TQXq9pSGhEbd47guj9U7i1BMLYRctWhlJmT/nYuuAMs
Siu2IUAW3spuoGCxTtotil3xyh+scTTJkoOTeF2N01klpbelDyEHFx7w0tZ6yOFB
9N4Zcg8OMLVw2YZegYMY6I/5T6QvRSkNQDttcg+Dp0nQlMH5lKlEW87cRSjRzwBM
BubqgvXDLf9sxNYZ8JtN2PEFxzChui8ViOIyPZdSpsdJznK7SbLuyik1rghDXMQI
9o4427bOVIi8Mo4ybJNRe+wJkhz0+CYY2VnyvQNCvoBM6E3Nmj7qO5ICufDr29E0
i0EiyWbQJoEwRQRILd5vFjYBKYJ0dNOw3g2/i9qqhpVvgAJHvdBBzyIQjWliSk7s
3177j1y1PHKOi+qaU64r6HdfFcxRN94VirOcfpnesHrXJvSyWv3XW9KdXirNDCBO
kmwZZSXONpmi/3nq9fxZzKS1voRxZUt19oq2x2N/EZNKfB0RKu3w5ab282v1AIyc
8ddOMSNKk05eHv97Jq/hpSmqe+DsByLpmUlmhK2uPBjDPG2yXgyWFqljNrC+NgkA
07h5qEkjlGxzdzgapVV2O1jpP++aCHzMvnQt47dFT8jF+brW+NntfoYB0CKhetUn
z4FqTiq6qalogRZmTqiXyOnm5tyPmV41nr1YMoMVjPg4nCgTF19gkj3Be2K54oBz
/QsFjt3+2dbwWtIW/hiHZVZ81209h2nnFXhM8kp54OBWFkBIGh6V3ou3r/ufWi+q
ZvOIuKWey1xgiPAZx6YDwqlYKwpS6UsnlWtuWq7ADpPlcrnJbLsgnxRCMY7bsjV9
P9C5AgkF8RF5pmWNOYdo9m+KldCbebmuCot5HJUq80YR+XiR1qHu4rpz4iFlCHPA
vH73tVgIn/+x5Nyb+jDVBHTstcTbm6bBWZ+661mOKQGk+E2JblJafg8tlkM5QAfn
D12pwVum2E0UDQ77Z+wHTVJulBDCoAQ7q+R2FmUDdgYta3StHQiQGrAfbCjjZhA6
7eJO33fHli9zDMGDBrE9r3IOvC/Vz6zkdDx3umAGFtT1hWjSnWXpmL406CS+JCIC
kiP3JnflN7q0XoR4Pkn/MCFwrkWF3DqhDVNR/EgirA1GZfETPsXBdBUheuMP6WoK
vOBbQdkCAPaTeDGkii/4//JZ7r+vhVn9xCI0P84ca8WKaGZfoRhsBZOKfhKNDE2z
6+q4RVT0FqSUS/g3RVEVs21B3VvW/+BnSydctuI+jov7sf9w6Dy8Gn8UHY8jTWux
ueFPGjgFIKBYjt8FjuxPqPoD33jjgKKoWjvMDDKNLOmU+30PiPWWeWlgznKBGlQH
ElBS/pHTJfrzhxuWADEkclD3Whe3JDmVb2gXJtSDqp+3CsRGWc/TxzaOcG8jRDPr
1tCoN6QyLh4/wfmYe5R2IdKaKATSgPvcpsWsFGccQ4tqFSZFZK2TvpTKQHK0DCIb
g8UhEX3r0EEU8HkKg3Fg55KG3jCF26ecA/6CaSBm7B1QLTiAT7VupQbOVejKioHd
WTv5BhkYwG1VVpdj+Qi6GL+5OZ5aBMdjFUYoTgV7HEv24ubqjI0sqqlyH992Abrt
CstFjkDu7VIKW+UnPg9sABqXTWFWKGlJ4EbHg3PU4BWyqhY1zTuuwKfOHO3kK+zS
DbiGFqjFlJvRKXrRaAlMmV9FZKqpkGqjUYrxMcU1UHyJ72CNB02TL6+N0vqSjQv4
XJvH6+J46o9pzRU3QvVCPQdq6i4r7YbvG1C0O1mnT78j06cehuvluIvm8ii+JUKk
sI9AohBVXBgyDxivtSITv/7LmycN2k8iQXuuOwEnO93BLQ+VSXA9MYZJW4BgNC7G
J9HUqMncZF2JnFtFUNd6t9IZlGoY0mjmvP9cNhhRFHpUdUxY7THGREH9lmf1RSP3
9z4di4yEiw1G4g+ih6B0cDJpfJXwt6c1RmeOuOtrvhVTHae/9QZfUInhCxyTJkb4
iBpsyI/FCJZbVujLUzqificbOL1xyD+pT+jzC2VbPZlybNqjdG4aKx8y0BRDWvmw
2oEx8lJhv+x5zZzVduXXWAnfuVD2NSAYcpOhffaBF1zpC4wk02kEawDddj/WoPcK
86wD+DSe3uEUs/YmTDgskB7BcKrC0AW+unbAkNxBZszjyf+jV/rp62nd22yC2Xjs
slfNV+cby1le0vk/CxGEnRYpZDGDYTr0QkQH3tH8BY5eteTY7yhCSekCV6Op+i+o
BFytgCDMowtUlXxk1oQjTqdVniDqj3CaQ7Otijm+JX81b6viOIB3VQ00DwSXZzdq
xtoPpgp5c6lUIEsOClBZUz6+gP+u+cBl6ZIXDSF7YMFj3HvdNtV3lRxRN8OOhfqD
w53IgVNFlK+BiDkG8uRwznNBOQfZjMRQJ34BYKl3pleOjfd7QkIT8xg37hqrXAIA
hzpd7GMXij0aRiEqnrsgaBmBFln0MdAJmUS1jovsSoQQSjmKQKzocHtPckk34Czz
jmFbsFP9WT0BD7iW5c+f8sK8m0uKVo0Sw50tzUHb4XXEV388joBOdQ9A/9Ktitup
XbjYQR8Oo00Z0/sa5nkLmKsEPeY9G2QKhfzp/twuHX+rt5Sfde/YrxzzQo4CRNcy
2uYC57tmYhzmppHLYMjzJNjCMtEb/o6zAHWYL4ni2GpKJnqp3I4cjhZvCZ2uEB3/
/m3sEkww4dwTleh7mbRfQTmKu447rlNKZGZQgZNk0XwmW6e3d3IY+09lqSt7DEMJ
GuF6fk5XasVvy6Ma1DV+s9HMuu0JvL9CHk7rHmzvMa1rMi0EFwhE2wGBIikHTlr9
TttOVKewH0BHWfkAqaIiZDKAaHce3gJeTT0qd0bstW5dzAAb2RCa70ZuJFqIGMXe
2r4YLjBPEB9fdsE/g3dYHVSMOvRxH9ubuzzdPm3Y3CaHuINQ7+bg5ugdp5lTcE1n
sbiKwpfz9WbLLSP9zJgwKRURrwWFstuWGEKxCTRLR35bDiy5enwboOE/9r1lBAEr
hMmsfNbTfcRZeDcp1aS0i5J3hZJy/gMi0XJvtjPmdoBEVPFMkC6stuUsk+mTWqq/
AUJlNM9o5Qe4dz7dQjps/whsHDRPxSn24AqGJzYAtFl6x+UaNF01Fh9FrTBFjI+v
sLpKcwkxsJeYf00o+K4JprLok4B+DtsGyS67zQFCUsv1QWNiUtLeLfLsBS6iSZBW
MvhSEjVdtHTDvT922lmFL/SFZuozneuoQgqGQf5zrshauVpCsWyeFKoowlt3l1d9
S5p7GaXcjM90qpjtekqfwhyMXZOXJ4nwRApO+Zt2HDJD3Q22kk2x+cCJ2Jc+ttti
Em/nepLZ/Y1rdtzq0TlFtEVBAIPL3BwhxtgjdlN7sVqL1dLkn6XvVwDB6/qVeL0h
woyrSWlPLh8wFn7I5AwJ96bm3+OS32EE0Dy8j9zRnddJTnttx7iVrZV1g1mpgZR/
IL9j6d/wNkzrvfEaBMOQ+enTQJVzw6o+qPAcKCdiMsijDylBwoatEsrei/MAmbB2
EsvKmYySPrd0MKMznsxnFihz5dpimavgQsXqvsNaQq+b8blk3VAUJ7Evg/z9KayN
IRrzxgbBANXOeuRu8f5Sev6RjoYHrmMzYLD9ldvPNvir6Y5lBkfvbqBYuaZ35TV4
/osa0eDyzx0h/ldxsWYI7OFwdk0uzg1LpZflD9NIyJH1lINcGolW9p8h14kZaeGW
4fiVJyggHHZ26IrQAJY0DZDhRhz52SPZ7LH2X43kWQQCz2BSd6tV+CIK191ariQP
G4zeniDOfVIAzAumPLblhiEogyCVkriH6cXVxcEMzv4ulNslChyiiyCB2L5iYz7C
cBwBaSC3Z1WmYjEeBcCBdlQ/NWnExsz4/rlR73bgB0kf2oNs/3KNvDa8wzGe6C8d
TFfe8FbCnBKi9T/mw6gu3K+lR33i3gowSmnd2QQj4KmHm66Ly/Mdys/pKRgvgz+v
bvrd7MtGoUBCeqN3QDcjT7eeNERCUjhZrvpwxGVYfltom1B86ZRnfBY+4OqJHyYx
G/MB7Op+t384rYdSDMPI0NLcBGPATKo/74GNd04wNL4c0hm4n1p2ekvBkK5lxt+e
9ST8h2uU/359Pk6qkjTir73CNTzKINJbJU3Eg0+G8nhrTvQQBu8tlRjSaATqyE3t
4RlR2w0l4ScjP7ce4NQRMvEtwzGncELxu2/V/U6bk75z54p1vqFhnGSuFo3riJOs
mE8faJX9fuagdfybKljsYkaVrVzCzIXiR2y7Il6JnCgFzU4MYq1++K3gaBIvP280
oIufzvBeNFXue3aXD43I9c+kl4uWl7NIMf9HExtO3yCnALZOW2QSIZZq+oTc3MOR
ZVTk6rEBUbV020ZYX8p7TsldbOberkkR6vr71Hue4BJq97ptE7gKdDeccsTJhKZ6
HiskHcLD/m25Dlh45JoJYBO45i+DDFKKBZqd2R421l9B6TUh4d68ptK6qmACM7wo
3EZR83qDMiJYAFqV9KHRQWhUZKNl5fA6xzALLRlalBL8wiwUDzlCNWKFOrB7WO6E
rvX/0u3Yf2zZjZ7NY8+DHv5JJhB5ZThUYJPKP4iFSeKVcPHxyvTMMj2GG1szVK7l
9wdgko60kXdCmuAVKXPzaE6ACTrUf7/YmBSRVkRI0WYiEf/sGo8lPJhMr5aidKhy
s38N8B3kPDBGFzgZLOk4SYPMjQv5Fvr/wMuKnqzGAUBUgalZ/leTMgPgTSjv2ooV
A6sCp2tlw+zHuQzuLE3mkMRa91siD9xUrNcDE9Xqi/e/br/Xk0FS8TFz9/5d5jDC
Qc4aUAEBcsk3yRtAuOqVQrBN1RPuBHJ0QumDqCIVhOp5vN8D0CMn2PSs2Hn11Dy4
lFhuYY+haPhqEk0v3x8byxxtCF/O9eXuPo5dT1T3H7P0S78gVvzkChBzIh0P+vqj
AdHr833zRPJKAaA0STUlOzGH2rFH8iDgzpwXR1BPrwCfYyX8/IFzksZuVDpno5VK
9DZnbFjURTSowO0T+LI/FRfDxp2IY9mOTZT1WZkZ09hoCBXdtmnJJQPltjlUyH+x
Q0uwaBfrk8XmaMApvDAcdzbAWdvqBwM7kosFmw2jRrYPig3C9OxsIUyATS9TtjXQ
k2hrxDprTw6cTFKcu0w11wZo7htQOtcYGmJJ1EzW49fv1oVkqpAuuPcH/fnDYwy2
RoiWuBTbNtJPsHBxOQQcQ6oPn4YQRLNdkuhfQ63s7INjGN1oVbpqxiBO0NhZJOTi
KZLsVmA+vB1INewnyTiRHdAb9exp7IJPKdSsNrubiMv3ZkohQ2gSRF4hUVxxmqPU
UE54Rrc8IwQKMZC+AVKrNAPBvoAo3eOneTt/1owK6MDj4Wo5ykszabP07PM38iVh
4a1sydvahEXoke2IA5G6xcUzErog9fsZwHSHAPfFmkXqQxQwlN/bQXuwbMXxYwsd
c4pBZiJZNofrVVCjTYf5Zfp6bj3UZqiyS2pcMutDsOx8zdZCYF0C70+qJQflRYP6
NICWji+vrlfp96WD+ecWWY4bq5hbOY/opDChpioXVCBEYcTMN1ToewSsaYfoVLmL
NTqyEOMtqgbcwRiCR6u+mSTNhVBVyrnqYflS/JSCvH0xIl5Id3xjFI6Q7/dtz8ko
t9Ai6cou48rO4hQPvWH2QU2CA8BDc+pR+CwdIyqAE17j+m1lp6HcogrUIwMO3tVV
6AR8z4FYJWSyk+qPVU5tvHCtUN/AsHVtjMVZlvzZ4d9evBx8luzhED3yZ97CGTcn
mvTtVelZqqZyNoycoIY67MFzDXlmBA7TOcQx4cjLJA06icOnvbkO3qVo5ub2XJZw
NkK8atDng5yWcIWqXCi6APtGZBwVWBNhYaeVCcwX5clYH2T8qEA27/M2juXDnvL1
7xFquAKzppqvtXTJGo1/KOdrK1aQsNgRd+nY4egRa0pJkQ9dglZX5kGu+Yjkio7v
zPToKB/Hl5rpBFyIXB+TUw+lqold/be+W0JoSrZXwSYciKyt9gi0LB7fCulCp8Li
pIxpkB/iBRztAMXGoWSPBA6IOsh59859dCaEy1VuiyAhAmSwbZKzYA9n0tnmMZoW
cDrPXyX9F7bjbem+p8OpViZKDfbkbhNZBHJY6QUkZkxw0CWX5MUl/O5p0ehXcMvF
0egfAvnbXhnQewXJ43wDgtRO3DYUsgoz7aWBdvHrRUN5+rE5YlGijWICkYLVP7cX
trR3PaSCMznh0aDd/hPcRDiTacknjp8qVrGFY4fpi065r1+SjRuK0hoTA1zXJt47
qs4Pb0KBwgEWCtsgsMlk+DU/NNViKIFgPjUUIRLF6aHamePV6JEFWBjxp87oJpVw
NiHu4+PHNJTgEZCOrNFpkqaImPs3wi+/DgNlTa8bqpto509spQp16HW3QGbg4ZCu
3efw0SbO2jegqaiiY8m+ABBc4U8FNd4Wz3ymAtJliAeB4m/zHjlF4h/k1UuTxKip
gCDovGTevvEKgZr651bnqAU+wMR5PjQ3gryadJM48XumRT0RcU4j8GR4PGVucou9
UrLWCXKoGV3gRHLM/pzKA4MDorcU9EZCgapgntiAUA39PxofOYq+vsbnbox5fGqw
s0gBwvLTXdzZkxzplkV44ODbb2de9fpuRCuIm+/E0wmjXHt3YIXTkMw1Nt56T4K+
/ECsMvzUrsNiPUbyYcJIkUwYI58e5xmbkk84sd+4XPPVsPNWE8IOU8gan47GSz6k
57s66XHC43K6kaOSyRnD6hcYBg07f8uiqlN0A4K3opKKb6tkynuFR6A3REhpCsA/
+iizxbs70rYtjvEQnddsvsKlGAkoFaQWwwRn1+APTG73+D9ccXdqO29FzSW/XtK2
4HCOjo4uSYegigA1IsuO1XY4Y7y3r8+CvSzL7hTwm809qeRL6r7/Mi9j0LPai/xx
/OmyZdAuFe8ARVWcX9OMbpU2IcjCE4/1DGjfWshiioi3vkZRHNwJFsJIWUfkbe5P
8bBFnFZ+am2242ht2++D2Ktkkf4YWutX0R65CerCoE04KivtauJQ2XsHr+DEqHML
i32xjm8aXnbPcTUSmpJ9XBwjcE5CjxFC36AUMAIw4drp/ggKZZqpmzJQ1Vf3sokJ
E4ZR2qaQvoHOWb3NTIAqENlGQT32Med5bwoQdUbAU2hYE2gGMLwKfRWOg9P8nUre
H6g9Dj0PKh4bMqmLiGQeMPRMoKq6Q7qs1Oj8TcnBYW0tLebWUYFdzZd4p6MvPPvk
OHofYNR1HhChn8VJPqqCilTNWDn7TmtPl1tr9TKF8L1lr1mYHkcwvF3bJ3rISqxH
GUZ8oVN1kkV3CNji6/do/fYnk9RTUveSmUfEL0ouu3jl6a1c/2KvvGT7kP2YFkpd
fOiwWlMSjx4dzb6oHIFlAiWDqr3x3JDsb+ZUkyAfuRtLsy9vEFmarnNRVCM34z6S
2JIDgrJH4auOYfmy3sk/z+f1bOy+kqT2qOaUFVUS6bvv1/m5tgWTQQLO/T+PtuA1
yuQCEYTjbQvzdAJCh1oyRZC8zagNt1JeG7Zr/jHIsUtzMR5qzXgPTqFVfzC3OWB+
CSipLx+bdscLjGifEe8HR7C2QbMIokkNdxZryhVsxjZ2O3NfnUrjjx6voud1Kx0h
bl5s74oXKlJKtOy+NfIGIiQF1Vu/gCnLZPPmVCidB1H1nGPW39cg80k7F3I469B5
FLz05CykNP56amV40xqJGAv9taAfJXFCrv96BlCJewBg9mwOYv9onU4jZi39OiOY
YTgxYGlrjF7HSCtqQyJoexz77rXuv+BA089NuiEzgOPpPTh8lDrWAvQGEptQUpCY
QOHEmMG3eOwiGvjN2u8P7orFyhLA5a0g9CJaFemAZTD0wCAE485zlbS/64W0uUXy
VBslW31qfc/gyMuXxHa/7FVv5DPwyPBOZZaj3UPgFRnNYVksUt85dLwWu2WfJAfg
FrHsklye/abzORK9TCI9C4kGy9siUG+eXqKuoXZnbFryaeULXPRype5smbjnmduY
iFMrJx7nR7gHjhtmRJqFAYf3ExmNAOUAu78YEMtyQPEhWEqlnRvmIZJx/fGvbUO6
AAluUzZfBur435utOWzg6M0/mfp5Y8xqEF747thWu+A3R4bDSaD/RjlpD6haSikF
au5WxFaOYcDMxIpGImQRQgTyfII79UboVBwAUhB85cwB9MTIsuKqkEibhH2Tm/r2
H//1fdLiAzkw0gDcpiGVmsoW57YLxGIjO96AbpiUaR3mbwaW9xoT9fNyIsBiFTrm
//z9+eynsw2jEitjO+/ipGlQc7PtIvAbqx4iIYhsIhD0EBkbbLXbS63T/LYa4tTV
L45l34KSv1Gx3e95054a3HBUxU6elAti+rLB2g4fsnXnW6EewSCGRgVAUMwyxXV2
bgF1yC02oAER0gJkzBeURk8+zYXvsrHnKqOnCMDDvRGCt/oKhRbmmU2TG5guYQgD
Yqkpzz0F8pGupqbklNWAwIuEFIjsmwJNwZUzERmFQ4v0frEfw5sAZvKjgaWL8emf
dEhbNylXJaWcLNuZ/a+nGXPjaSzBMX75+52YN3NjQAouS25cInzXzxUuMy81ueLo
L/i7Aa/yzKF6nbCCN3I1Lr0Y/dh8sFpN1IT7Mok+CknbzjwZIJswkqO/vA/XNoEp
iu7XI+YRir/ly2MedKtvhr3P6FuBSadhc01vQ4f8KDMTAlQt/Wtq9lyKvoe2tF7v
XfnwW74qDaJ3Obbrixo/++ZH1g5auqXLyTdvLX+2MgCVLbqifOe5eQlwB1OgJPOF
bdHA1uIXQLTOWgdtE9dr64C1npOjF/BqqHq1R85YGUhivZR9QyD1Itm/PBOItPSf
40F2rbzmU1qIUFcxNru9KeYfqhA7H71wZ505RJWHkmskO7KqMBdSHF4hYBJJI6M/
3aFnEh+RuKAG+cA9plm4nvhsdLXoXdzqB1n0bDD1LQTNtmUWB+djb5zezLTEJkih
3FBCRSCxRoY6PB2cGZ+d7t5bRAHsgu5C7CW99xlADKco+BeiobFVbc7km+L2NuD3
e6ozf64fq750pZWrTK39KtwsPkdbPvNJE2IlmOkWmekicJE95yPyhv4xxrrWl1us
NlCFBjZ9LszvOlBUgHHAOl8wDI2t0f08aBF355DgXztvCiE40vv6v2/d1elDGaZW
L3iUyOJJ5TTdBO5gyt1e3l2wZPC28boTbdVhZLIEpEdIqwGAZgEnYLI0BRI/xALy
vUVK9QgBcNTO9OicQdGFErqiAIFmOqEtEGv8pQP3G3oyH8CnTXvqUstWzxgqQ9gL
3XBeI0Cf054BKJZMeaxmU61MMdz3jXRdB1wonUnsqBHAA7U3nhJ0+iRHpKGc/zsZ
vEHHDjnJ9hvFaVXXE2y7htVG7vHqeCm+Lgo1rBQXNXbnuZLf0pF+4Zhj31WnchQH
C3zV90Qa105g+05BSIscy8L5mjEyHTBNuMeJxPV6Ej7R0SiS9zlQ552rjn1C+qrP
SbvYgpsP7mRba/YDMQUpYp2OpU+l7WURXVV2/PhM6foRnZxGUaK2tc4GaXEDkWoM
iMfg+fWZjjNMwar2BHSXnncmOJyQQZThUkeoMvPCsX3fu/J876cuiLfMAfWQYUvT
61tWOCtWt/kgQarbOswMqulUPn1kZSlw/glOpmb1tfZAaerj7nAxGaaf81TYO+8x
PoYPX9bU1BnsSfxae5956sgwyEHpsffGPME6Hyprsd0rbFNWbqNFEjWgDkUnuBCf
aPVQJSbBQc1fRZrvB1yyfVtO/o6EJgwsJCCdKUVXb1N0GUaCUICpO1L+wtsYQvAa
uCDuo+Llkobxj6U8hTA7wEoE5pjW2QedxUVGMG5hsREdQwQrv1Vss5A6yIiUtTZx
aX8wFMKR+M3hGasFYAMRBwfDWNnUPrizUmCncZtSb2iNwM7Lt1MHEJFfaiDp4FaY
Hgu7ZQFvMeGikmIWB2VhmpirkBbMq+P3sY2Wp8tlCOjT5QM3XHe7DEjflys0i19g
cuVEXFlUgR5id+KJgfCgKFPYUJUec6Z/HTOnGNqmqQrhte+QA0xSNkt4iCKTWodv
GowuLEkghorhbuG8E5j0LNKW7t7WFa9S/GFwt4INN9HeECzqPJl0gxLcu7u4+q+E
+h1I7lSbog0P9bPE9Ee59IyoMWeF2fqR0mNF73MzJWqZz3wkNOgJUuRsFD6s3Tkz
/b5RoHGAsTZSiVGLY7HgCt5/jLzAuuc8Ooys1ztBimvx7EpAyXosnmvufkeaibKP
5eKgW6txXAUqPM/LcigJ4W6sJRFDcye3i5jqtOPe2mSEIDpAv6yyYuEDLsx+Ur6Z
/X7sapSXnh95ugMQMV+iWNGLmC7hFE5NbK4xXlev0aCvdZQ6nuxgYiF5g4KgV+vt
YSm0xWzWYHBmVCEoGpytHxrnzUrYa7vFtpCYnUdPoK15pmZoYeENoOBqvMkHPOJC
PD6TuXJhumfHaCDtMwKI0h7KvIJzFTc0Xa4U+pvH/j7gNVwTqxb+t2XWsChv18DS
sL5V8unZ/Kje6BJodykoSVB6ZawIwnGb68bfLfWBd4y3FwSTdnhLXd6XbpjlnzIK
0fA3fDMtqh9+rboaP/qxO9+SZVsv/GBtolTrOdo2LPBsh9pfIpjLlPumbdlf1TMy
VftFydUGyh0sb1a6cp1trBr1BkLFataEz92r/cr+QeqQFULOV/+wC+53FoFcKCpw
wuxDSE4XO7yVTgHxRC1KLc915orSw/8Z6e1zNVDYY9wObyLzKeBHv1mKfErGa7y+
u1NKiyNi+BT70ceSQPR3qazlGkDsp+XLUk3YrclozvzR/AuObuAAX5NtY8RV6vId
bxBfVSUyo2Jenwws7Ms/0F6ivs1YsbRmkewPDZ3yow+/BFXxo4hlbrTQxvKNPiN4
YaBB4NK2+ppVF4cxrk/fwTJMsjjnguXtcalc53EKKLz3sxnTBkoXlBDICOj1S0EL
whkn/szbKQZLGWyZEMR9ira4cI8XhkC68lgDnXeuK8KYg7Zitr0ULT82w+xFgL6D
6r8NF+JHnXeWtoCOmQ7RlYvCgKufq1QO8MZrD2kkBQknEqFRzPey/LWrlUXkgrfy
qYNTwprXlUd059sLc4rZVRh+w3HE0ow8ZoBeT9LS7GMQVvTlWI2IQZLHKgnsY0hU
e9t2Nb2h8lazGlukcIxVU4wTBDM02zuwlBix4eXupkbIXwYwGFMhVL66RBsfBko4
KHqka2le21leoj3WR+GiOgWl+Y7bYtGymUxGaFd7i8KuaxPE02aanhubwr+ZAvjw
ibwtUvWX9LRHwWJTbth60bCzBp7dp77InNabQdw1+sLS+GlehmqjN+YpW7QzmP+C
t55fSCrRnsSdscats/w9pklJroLh7mpV2uLDU5oaoCt2zy5BS4tKymsWvvO38kaM
00WmH3rmU0dz11V1iDZIAF/S7kd+CAZZfWnU1u7lhwgYZpDnrUzWqknp5EoB6ldX
sh9JpXkAbKn14bxmXy4MpwZXxxWjqlNo5V+uc5OUuiEzEv//xnO38/6UvwUzFN0x
X7ve4A+ASaaMTUVVtsobzmWRmQLsKk+p+JiKHzj9e70OG6dyJ0vSMiWCD2jxQ7OK
xFj+SOd7oy98jrtp4EacHYNNggijeIUPsAp6SnrwKbmb/oCyRV9opVQb8Ilsy/0e
GeZgkIoS1wBDGnyj/GhsZ4bwScM7qkYbpo1OCUiaiGL2OAInu+n9jkPeZVEb+3HL
lr8T639EYwlUA7fjfW14QeVzzjpJlNw4J8HLEL8BLLRjGfV/tKAcs/pY5aJwrs9A
Swpt6ySNXugZLtYc2wgPx7qoSmJLgDMH/dNbQzvtY4jcVriLuqCAZM74GMrqhDxw
g2TfkzvoLzcYi4ab50TOtRFn5YjyES8WW3hvTWDoqQvpdQReYpIP/itkWdtQr5Lm
0DL32bf8xjaujh4O61aRdMCOiTZN3ifrEqvjBu+1ojK3HzbrIxXU51WEsVz2iBBn
LxBbekErdgEBJXbdUlZvFx2CofNWNJkYYFhTOIBfciuQiBFStXZzrTuj4ozuQNrT
AXMHASzfa9c9crtqs7KRe+XYS58WGBTsBfpdjY20c4/yPzySuTJ6o3Ig31eHg/ia
HPf0Ay0M4wYok6n8Q/E5oqRzlCd2eRhCaturLEqLjuFs8Df0voggDSYQPjfNk3U3
sc+gqufmRYax4x121oi8Bu+J+SSMgNnrmwNcIMf3e4LLpznKYfHtSt9XGIV7NKKg
4kWFiGxsGAmSPnTMFUbNM/OM2N0DoZs8maDb19CB/HzgPT6yGFfqDDGnpqNmGFPt
hNRRsa2Hn5hbZ3gXWVNZGH5Modvu+2/30WJI2sZxlIpGPxOzBFvlVbNZ98CHmZSZ
Eghx6DXIYC4P1kgSkNiiCr024L0eKSZG5cO3fSP/1Oo4rmx6ivT7RXOvEl/NPb/B
nPrABqtg1zLU0rI0/lkYqWyr5LbS4ajk2GoCQjpXOnSIHRLT1p/cTe+t7oHdGagT
V+K/xwqWNQnz28pO5NoWdwcxwyo5ptA9xB4Ku+zIdVsyI6SPfNmFfatLtLdmrl5G
fsG9kCibFMvQb8kXX5a1PTCzUw/dx5JQJbZuegr3Nk+akgBTTR8GCTtOPOYlWiim
sx5SltzcEbTegoHle6kDMinQbuv4hhR1WVU9Pi6i6qQH1n+X3Vr1h6tahAnWmFC4
PtDtHDA7TZp7AdLPdr47CqH9JsK64wwz2j0CIWfF0RU9zApTEN2c+ZbwSMd8n2wd
eOOGEfntXSkvU6cQ/yzr5sPxLv72qrUE4MWapd4wf0/3ms61GSrXgvAqbw1vqEvj
c7MDRH5xCQcXcXJJEx1HmzcOMY6Trd06agv0i3X3v0Pky1qCyEdgrtdGUYFki0wY
T6Gi/TWnm92WYNg1/yfGuvUqhcvYXRScgsGk++F3k3YH+DWm02ZVEAGHrgiBCeXX
WZoW9I41X+I5ODHBmQXaAnAFDOtwI4dF4so1SQ4lGnNSQg/zi49SUufmDaQ5wK9+
T1/PwWKrbC4YWA4SMxQWNWBelG9p7GLgSpTO7kybPY+RWyWlQaoCAfm/xXSD5iJM
yGdN4v1mNnNyzsM1n+wtj+KureWTqvkWR1Jsp+SS1J74a/lcy3fM5RsmpM7eSBIo
VhCIgpZMFycrom6AnpaAQd0eB3+hvujMB+sENvf/a73nNRAs2e0an2oKfKzWDcrD
fJDJJxYM/PZzFv7856UB88Tb32EY/NHNbSDpWU1NFx31EupEXQSVSZ6HG8/eZMJ2
+g/EuweIECWCkW2xCJ9nxt0k3BAaSzZIqiulr4tvPlDcQWUA8Ek+8Viq1Xrh/j4L
IRORt5d6iIe6LbNLsHuKG6enD8uSTiiDLkCDxkgczFMDjhl7wAnRcRKCatPjWncf
JcmBexfXn4JIzC53AS57BQjqFpKT+9wZgECgQfLcg6CHoz96FjY7FV+jUxGnNLH/
g9aGurZR0CWrOnw3X0PnPu74HbS2MaUCs+bmzDXJXg5KpErgizXEBndIrC9SNSZh
/WQ08+XcApPG8wDvFvM9TstxsMTxcJ4lgapi4/ae6/7b1yijz1iphuHztaMkw9oJ
j3A/jmS/aEyAn4astDnWcVYwDy9a3zXIAbsFnwdF120g75COGB4yARY8IY0ddJgB
G1G/Mm4yvCfOEkMXVrHl1FbFai572PnV6Y1DuDq4gyx+Tm8ew6L0RB9yu+R6u+pw
MlRMMSQjfZpMAI038tzwzHO3X9YAfzwHPHPjMQGe6qjgdgfQ14VHMPnma+mNfB6k
ZeTTZNeJJIsNsDR1H7SkWt1BoH7JAImc7vvwqDifzhY2WbRjCHtGRgGz3XOO2SpI
QE6aVdpENBM+8s+SCYfvx9WfQd+T9Tc/NWDAWJ+Q07e0niFkdV6Z5OQ1amV9WMkT
aV1UnzAMlcY3oCMiWNBeMyK852rItWN7iz9hzM3C5B0OpJEXFaNzY+JbkILTUR5u
pWvhtswu6ciV09cK5W9136SS9wQv0KCqgF7bc5uuP+ymYD8g1bcL9aqZfNi5aZwh
pWw+wfwypoIYgMz6GSkchmBlRmrJv2MPipG1pE5IzpCsZPlLQQ/na2vwZEMfIjzk
+D/REL+OFafmV9D5TiLM7TOXSxSHgrAc0FM9Bt684Uuxm5aABe0hH2GHFj4rTX6j
P6NOYFQdV82u2tTfveLaY78iOk0DsLOjI8gH1CgKq/b0qeSZIA2IExlX15EUTi9V
/nOQjXwKbQESDEYgOy++jCZ8CWW5xmsaKiKU3ZdjdGVa2AG2YnzM0VknZFyBn6Zc
X/eVCWjp8BAU3Cfmww6++LNCCZu68+bz8AnAWVXgJfQC7wLydO/Fvg0GBNBh8ONH
+Pjai7jjXAOundoR4S8ma0gFuClx8UDc/yGcsQu7Z11FzeZ+OR2lkxP+ROD8b8Au
SlF3ctxrnOBqvvDOe8d7kOAh4gSCrMrbcpoklGE5byRxwCUm7Lv4fv1M/isQ26eb
/XKhb5sr9l+Qehb2M9h8k/c3uWSmpbe5mcvS5Qgp4yj5ULc+Rw1+AI47vAeg5JtT
vxtydP2qfUOngDu+VSFsTluQMwS91Y5P36uOgQLc2UFaPsOu5Ysz7CtQ9knpc2cm
LypIN2bDAhcg9bFq+8AbX6ufCzU6bnhITbnwPVcR74wg77c4rlL5CNj9D6hGkVGl
AhT7b7VEaj9guI4E2sKkQT1Xy24NEtB0X2UvY+Ujq/0amybiV0b1W7pIOku4wK7F
jNDrs8B1Z+8v0e7PtsMrYXTy/TgtJ/FpUE+hahfAC5eqC2jOKw6zEHuKURpLr8Hl
zaCHe75zLYffZxVx4nxbbew60PRdUaBjUHh39S/NHGMdDntpXyaR8SsdOABNqWaR
NxzhyEQxC1O7olxjwjMFdRL/v5NuM3DLEMEurpabyzb4FukOQcvam52f9h+AwYF7
/2hMb3pnWlcH6UdTO+LpfcYsaIfjP2aE/Y7KJSZqIA5DsVnrSeLgFBsfazWtP3+H
b7lnM6VSKKH39uHTe2ZsCWhcRaXLv4W5SK5TMAh/ThaOuS7nw0thYuyN93OK3y6+
Hnu2DRj3BBd9/LTYuCAT6XwXBXsxQtRQelUKzF7m20M07YlkBxEKHtbzlcpqNBJQ
6O4/Rh15dMy/WKNp3ANtXMYep7XTm9bbnMufLjNQrsrxAxAOTPg0W979yxVwoH8u
Q4ErHkLn11bvE/z5waAYJaRbfhPEkVxi34D4aQmfeB3TwKR+b6GvQ6cYVINnVj2t
OTnKJdlTu2+nGc0Rvw/URl4O0uMC5NvARPveuJi98QNpegQXfzOjVWv11INtq85e
qaxXSJdNNx/QQobx7juRcUedVwJnJEscHRsABiUFRotFJekX2EzUlWoQZbes2bVc
pTQpKklg4UrpW247SQVCve92bL1Z77dJmX51XyhK7sBumgvG/hDXGS9D5Lo6ryL/
2pGzpoOqvz6ZMpWS8Jq3ANmMvLHg9VWxLs2faj50RCDwTv0iz8XWyb1LhsznqiES
j8iRFtq7hsMsmd3qgrC3E9eyog+S6pjwfjfdFfw88ejPQcIDypQk57DOL9oXbgPi
O6m2rCQosYsT0b0kP8DKIayLsAsT9hY0LOhiswArXvahFB9/A4zEWHwP9wIfBosP
S/QMf4vT1a5C3HpOuZycmBlAsP8gaFb1gZ2U+iP8WCxW+oXYyrvuLLQMIBxtDPMt
LB654jD2QH65re/hGN+NUzcA6+iyjsc0t+ILYmqKjXPI8xGkuwv0Ya/aXzhvmgsK
yiXL+VzeTpJ3OUp/BAndSKlSTbW0RZw3ouVp+xM6ezBCLv9k2D4SAhU9vm9Zv6SH
FPx1GZl064lTTlhEQonfrFe+w9g/hqBgVQDehYlbiUScJcrePl+OYisy64YgoGIc
IPTJ99s036JJGlaccaVNrS3S1FYaJcA2Zx4yj8DyhwL4iiAeyBIHBrvZ0JjNbdJL
yW+ASTwNToB45IsZtc4ueFkDOqk0v3SPABW8TCF5RpuC+1lrqMDRkmwy4C2yOYEB
fukBeWjxuaC3iehqDxih5ncQTW05WoyZDSNx4F1eiBw+qVkKb3ryhaKW3ZGidzOw
9H43J5HCMZR7S//rpivtUJrG980LD6F7GO8aDpVTMDB3SNRHVc78B0KT5404GgEl
qflVnzutsXSPafpbvw3PXWVxpvrM4Pc/xxhzQ6+N1iqqH1R6Xi+P3NspBfEW/MdP
xjQ6xeNZL9yn3Br8B7JbEppsEejfgjscPWZoGF4rXcVa05LNDiaB7YOaUsSP1XM8
h1VLboaXggrCM8DM8PoJg73Zv9ZdXN1ZZmp+01Uw76xCIPhikGPWsT0tRab+1MMG
StOj4qNplMQrkKR0uuoq6xiY2MwzQu7hzu6lS2cUDw6ocLjQ9NdSHyF0Kds7kF+p
2/Sbyyt1Kmv30IZMu6/pHUmufRv1/T8kFKSLnlt5t8NCDlyec/G6rUJkglKMcYri
UJjeXeYyKHaNOeTCjhnCINIxKm2dBVksoGUjcyurAS+kd4yFD7eojSDrfLV7Df6y
pFKwyREMcWPVALxNnsA9X+jLHwMjfKCYq8SPcVEhSKG7j2IiDWkRBnczZB8FqWOt
HCwgvsE6g5Nn8cy81g+vWM6RfFV3PVDiK6rQeC1NkrK/DMWG7nCBrkHACxSjMNMe
GA3WXfnqXhaIzRuRU0zkKMhYchY9toe4iYO5I/Cm7WCxZjucOcJ/BuYMrkf/NH8l
QJlSi3O1Xb+ElQh7xWuqxusWLR1HtgFrD6pZYujtIHYLp0YZm+BG8w0gsSf7FLKR
1kz/sQBMO/2Ld0WviDUS49YmSXnDDOj5o9YNVC05SzLkKREIiBFd7F9P0YPlUqGZ
2IcnmFHW1vJT7rWAXR8LH4CCROHuKQUw7XvlJmCLpmL+LOa5v4cZ/5gXxclrZTdM
9TUbH8xsEGQwRf0NVwzgTmZo6WryFG1Lw3a8lABBFBZyZTMjlOdKGoMGk2OmyTCA
+28ukjI0hLVRHXkhi5TDYr2xwXQnkWjaQfTcl4Y48cqe4p33XWSDO+/GEk6RXAVI
mPI+CpxD9aytUD9hUcmmfjEo+vHGm1nEN3M75g+SrzzyEFTdK8tU3rqKBZ6VUzI9
u9x+nok4bIfVMYJT2SLB7TwI3AozOODJpMSjFURMueqepwjA7VBObpYSIv+dXeBL
VsO/AU6n98WB8o+mHkMy2Tgf5FfLU/F6ZcGlj35Uc+J0bWQxbZYE+bk/vSBi1Lle
ZtU3MHEhHuSR5Mjd6+1UumLZP4SsCzhfIaSJAgOS2CRYS68U+xEqrTKPzX2xyo/9
M2XdnNoTQFDhZGFf6vxmCba3P6RMNPA9WvEknPmIO16KCuGCFc5ZCFvt6111mG+x
cr6QFTdi5hxEtUVaOptcpcYK6iDh0coOkbBTU9vnG7lDrT7wBEPXUIimV2m68WFn
bei90ovW1Kk3LhgLC232B9UtoRGbQ/fVKo6jerH8ZlrVIffe8bZvfvtEzAhOp7Xy
6ugEaScUqTFgffb8wiozZUTvdF0TLgwH4kLrJNqB1+7HsmkbdY7uA+ZTNFPAAkNb
wg1CfhIIkB/lWAs//rejWCGEyapecqZMWbIp1HNH2KuxaRirbR9tcofkDEcgjS3W
rgBNP2DKa5q5xXoZ5XSsxKsPscnvZ+SMBEqt7qqKrW8ZgAX1VvORzgyFlWtRRmlP
p5v+yBxBfKT0DnlpT0PjLupx0HOlC5VDREB6y/wJ57gnyWb9SqD/rm7JzaNbqdvc
e5LKtbs8vmNa2z83xy35ANP37Jt7B8Lkr2bAYEr4y4on9rC9N0Bnb58unXv07ddJ
cIn5JjL1M0rYKtYwnpl4F5Qa1y8nJCca+CzivC094dG1uGuBTIRdQ8Y4cLoAIdXS
PeLFMF4EVexojyqMcVoPKLTAFgYzjGrlsVGoN/5c8BF+y8QcSHQB6EenQqQhauJs
Y8Svr5uvG4+gfxpLu0kvisu4DNf0c/EmwIESewk6EykHC4KBR9IY38Qc4UABy0Ls
sacJNR6+c4KV9pkdRZWIzP7qwpJlnoE8yQ7IjdAqoLc9uUzMRni0y/LjdNOpIm3d
/Lchwug4tZhgWtUYb4IXepEtm4mluiP3MVNkkz02xaHSiFl8DKhStwdItOphYnqA
vrsCUPk8airz+oJ/Q+yi37cU1BHqVTC8wjFeaP4IFDXHrwYDypQOVsxBsnXhl8dn
UfWy7UNfcpcHR3jUH9mbaEuIoosmhFunC1guoGCaFJLO78C9aCHLc/NBuO3P1Ib5
Tum2F/VSpxxjUBjiOU+VnG9lPL5E+LgiZGZ0AxdeDjXAW8is6XkIu9i49qbDe6Kb
oXTztpJtLK0HG2NNua6ArhU4Hi8zk/+sH8m3NCygaillW7PNyf6cKVNpjjcys8d7
jbL47/L/VRSprEMHoZky1qF9iDsobuKudbY72z4oE17KlFeBVZ062MnfILf+S+p6
xu6yx/BSJUu3d6eXU32k67kNCuiPCwkTFDNOo0g20KsVhhg7CJ9/cGDiUqR8yWPu
x8xc93fo/EPtxOu2xGjtNjlBZ2m3z5MHDY9IRq0x3AsyuPmShooLEz8BqLDY8FoN
2fzh1JovlCNyXF7uDuCQKBTEFrVm7YItdqg+LptKePAmlwxM8V3iJfe1G5DdwQZk
9aqgK6EO/s4jjhkC00O88twIYOX9YNnuW/xqm+m864JWLSbs2dS+1gQF0OGPCI9h
PwQ7R0TebcLxaRDt09x3KMYspb3/9tg62Gi1kQdrVY8aO3AKAibWAT6Sz0cux/Qq
52E9Yn8IKQW4iJOpZbIxocIApSMjW1EW/azoo3aYQ+MDcQOD9DduGE8T3xvRgd2E
ymLItxLA23lznctD50ntzFKD2deN++IpDYPxVEaGlKG7YVjrEyhLpNhHHaxNnwqq
XYZGN8Qs1KYN1Zsbu2tROAzVgpCcUiH7iMhJbSOBBTDTrb41FL4iIg9Ho0VKwmUD
kLoVUdxr8Z3b8FFhAt13czkvB73c3dZj9VPNahuVQI2RMCeK8gW75icUWHPK3pwI
JOD6t4NEVURDh/JH5WBm4NRb/drS02cmGoiYJh2c1tXY+fjvBSniuOZHdVNDQ4KF
j7G2cvqVdaSztmUgqWDYbMAa7rourqEvx7h1cdI9NYH+fKW61xuV2B15ZO6i+qas
Qe8qsn1Vdet8LN8zpJ9cYDiY9GsvMbtUv429tmsnhaXAJ5qHVzYku7tbhfxwJQAj
ac704TJ/CYkth5bSXFYqQLZxR2//9hhYHvBCPTI/fTnAKm/shwHBlZcpemcN10YG
RwVLuqh7Uikjk6X7zqBF6W0N7jcOQPs+HZrChdh6GDq2YaScdvzf2+03YCnWXVrA
H0jRqvCocfseRSr+Kj4zJNYh3/pHaE6XGhxidWmxiY25p62ZyEBhhkVzJ6TYNs3x
pr276PV2zIXxZpEUpeWEpLR8IdgzHm05/xf06XqSMIkLQNPx0rSqYl2xp85pxmgf
/mrVnLh1P32t5Drdhgy6eMqnBmK5gk9jMKF35PTIwVC9nqRY98CYuupg07K19HJY
wDu4IUFQL1VbVMn/K4MNcP/pWtMQeqlI2gOH6PWWFvLwD50aIvKgCieIJgj1eYhp
179bkevUNcDT67Tup3WMXxtk14AjjQMUABNMwms9Q4KjzJi90gUu+kuTNEQ42enY
6UefKVk7Eh1HZ8zogaK8GqaRHArczZgFoLTbBxW5fzs4ywXQOeLprT/Xt2qlxcg/
b8+O9WQgi/zhR/WmGPWm34hgQHr107EvsxZevWdED09wQAgG2C1SW0bhW7qq9x6W
e1ygRt7vtHqk0Z+VpsHqEuNXLxpsPBFkm72nVB43hUsEYZaC4nWOQ1b18K9wxwro
6+A+uRh0dTWH7Tsg7aXMpZWytlilXQLyhKRSLq7SbQxKm856uYLDx6gCHbIh06Jr
uwtvLt+UVc7UtqlWFd/vGUxSnYlsoCpiwelzEqx+5nqOD+Q/WP6vRP1cpPz1FLiZ
CE6qtElwp+Bm8bO+EtnqBTy/yCehMMZJP1KbXtqXeZceExkorVn/BpcvoRsjphMH
bAhbUKPCWmP3onl4s7ouNrNqwtktrYyrTgbRDTSjdl3L2Bo+/UsbtHEdR/xWH/7m
2Pks25PpteTI1g7NOePAvAJ09+SRgDNa0Bq90uEcYu2/OGUivPToMcB8eARgKy0w
t5Eg3QT1+xNpMwdbvbKQ8ddBjuk7MXYbhtlUefNihZoEP5ka/0wapCnpPFV/u/Ro
mHitgvkxuRA1uIoB8P4/IUBVzLNovjvbTFKfILwD+5GBBO02d4vvBykLX9SkgKl8
AqMLLuBbKwEKeURL24yBkhrLv2dp0hMob4t8gWzx7i8KK2chSNdkfarTmEJ9zsnD
XMZOCdvCV1SkQHVykNPq7x0AF8aczcnJc0TBb6DAvDlVWefAUt4yJ/A2oAKSPIKf
x1FnEDHP+Htfkdq3JFT28SPVck+KMd2e5uvrbdWtm1qWbkf+hyFC+tifj28TYHXs
MRW8/xt1fzpA9rU+Ik461nvNPfU8Br4m5bISQlLA0zT1BVzTmx5/btj46v2m2h0r
5+dX+djvTM2niLSsKwfAvu0AK7+AEQ7M/nfnbjDnCt2d+xWoiGNs4xjyes1oMx7a
29CMy8YMKMADGzVXNfChklchVCLCr/1tM9yV1SKqS+Cr9LYIPgMYQr6TYCTuTzIT
HZ1nWHNLjMEg4o0SMJGm0GBDpF8qUifkQ/rAkO3idni0JbvBzMF4/9X8tSIXsbIG
1hapRosSU2ROK9CFqufsqvwWO64qL3soG1B+pTvpNioJzr0GGAbiCIpulq+d1KPF
lXC2afdqudvTM2YNpJs8FqXy/mz/2NGjbwKz9+m5yEYxczbgelDV+an91tiPOhH3
qV/7GdEhCPQiWABGqjwusem99xFG78T35kOebnfuT+zwMLIFiZ1KPjel1g/gVq6R
sUB9UD0DAePnfZb8XI5ZOHUf5LYQfPcIo2RT2y5Q8YiFds2o4PdfR5EHRNhzoeWU
AAnoY11c7FgWgRevzax7vcQxiBBSZktPQ+w4nMaDyWVW6B+9WCzRpy460SvkhgAG
fMaMgpLG+5LvclzkjLl9neCfCvIrsMClljsE/X69hLvWUSOFFoRyyJ4k5q491SUM
3zPilbeDBHX5EIOt5Rlocuxobc9flQCMeaSBQHcgeH9w00jkjiPV1AkeEWEaTlUf
MONvbm4uDKhJvGuKhPctvvTBqnX/DedNyeZ7Gfvp5IdFoN22hgAC2mJ/vdZF/eyg
7PEuHZ7bCkMIufnL9SJD2fznLNFPGLYdX6A7T+sV04fcJNRVu79hJjVTPqlgjQKR
XJi0sO0c+Es4eQmsEodQzBJbjPMO4ZOWr5uUNnYWx3kVtYp53MPKj7ykI8XiW90q
o3kurCJheKuxXxJy9aMh0EP83ZGxzncMNO1NFwfc9P2T2ePHb8sgJ5SmSiV55it+
oQj9xVVl9ZYcZTc2AwlImlR0GMZDLSz4wTiNUh9mQFmNKCTTzWIlKV4lwhPuWSz6
jbv5+nRDeD/p+jPyou9cK+O7EalLRUoIWe5Di2rseypXWLFCuu/Ly4zXTF3J9drB
/Xk1r6XIWiRa9+8Kh5iZN6O0lTD/HQLAzh7wUYUJaENVo9onv/yMAdZVXdA2lMv+
q5ElYQp+gVEg4o7dEkCCvL7lI90y3YVRpg8vh13etc9VAlGYQmzESep7DrTPyytx
wG0fM0Vvp4OJUhSO3HtOWkdYE0wBQ1CbroJ7liNxEKCf2JDXuhzvwL76aezQQvpN
hBRwFMmSu4PS0AdwTF2yL16TqhA//Zud4Zh6H27/jNkXxGEZdrGIA5nqlFF7swUp
nXewbEJY50IkTMVsJur0W8xrATWHRdh/ksT3KP2vrS3Mo4Ypfz11tJYHFzS2miNI
srxQ73yxKmelWDReV4X+3blza5C6YmafWaV2zcwaUfjDz+nnWEURFMiuUo7aXQM1
s97yibHg2c78a3YAlfWTFI4HnKslYZ7KFASthb8iWfBW34RmZc18b//cmU9hxXXa
T3ydTlXBjxLCim0UHYtA26sAoHzjHv54SFqdKR/4W1dV8SFM7w5xDSDl1lFS3BJV
2sfQJ4M7gdIu6L42KzFQr9GIy3EeI+MTfFpNarJvfDjsPFWBPF2x+ZrvsoKMro+3
NWYq44/I/BNnjGJCXUBo35+6AS6qY9eydRNbXQZT6S/P+zHbuwQlVupZkC1LORk5
d5B3pSKR2IEYbg4f13w3RXxJMfXumAU/pm09U07y6eupK3nJI9GxH4hlnMqbRw/F
K3/PeZ9Hn0yZD8xFl6+6BPL7we8Mzwahqe6AqLrp59rMrfGp2nFwYcLVhRt9tF+Z
DdRbjoDtOgEQeGM4q3KJIGqogW4MFFSkmxcXKrEPkzO6izZ6CTl+yxzwI/OQwxlT
EAVgbbAGyF4q3IhcYO9zyxdBw+pc4h942XbJfS18ouOf1iilYv3cewhTVSv04nDU
HULYZDGpP9W9GDi2o1FrxLcG1dj9N8su2nLegNs66U6pYGwHdQWV2Km5CG8P3j0q
rxENmC1VndjZPDFJ9KiYggb39REQ7q+1xGJwofAP32AnE3vPbJaKVroJQYLsrjQU
LwIA5t5H9uLGglMXUdVOA1EmfBFSjoh2Ko9nNo08pw6i5tGI5cvXJvudn0yuZEgD
oRA/v2wgDIfJe0CjAWGARY2evEcMKQk2tqXt72PNe1AC50Q0VjOVtkoQyP3eDqG2
VjJehnXeING9vNWEhSLy72RxHwUdaJJkxthNKqd39JAFmDYrEZt3FfwVoSNBHA07
smli7HnqfxuXh7ZOUo2Nta3rEzPU173FJQBQB/3gRZrtp+j/G5JA2n1/FGWZE26a
wasgxjWiFHGBiGVck5mpo5OtHeSr95BRyz7BH++Q9w5x6lxs+Z3Ce+qh9Y4Ya3SU
6SdkG8pgqYCpiLQ1Ig/9fkREHk9KChCig7jVW8xk6bbotfkVTL5OJ/I6EStShvMy
QcJSpgr3bPpEwtD1ZO+yJJ8TAkR07F3J+NumO6UdMx29Vxji7vK2ZyTqBmVvxF2F
odcizJCNchJE4fp79kvB/sdvXK/GOjXs644imu2q7movpglAmaPf0RmlsYRcUc/H
lOM6PK+DZ9/9dr9H5WPHHbFdgtBsC8GLCU5gMlqULdUofHL1F+h2AVknWLbGMcfb
s4TlPgrZS2kX9+mRNPFl9c/K7FxgponKIR6uQ1QICZJx4AO10Htuv5u3SMaWlZGV
sDsJz7axDtP8ZmkEMINEqWc2VXuWaVIHPf4ONS5PS4Rc/O83xY6ng5dqqXjTlnwx
3wjYtm/8uVYEj1ZWr2vNVmtUeyYMaUXiSko2R+u3Q+008ljtBW2osuO505Qod9Z5
zXMTQrZo9VKlT3sMxPEIJLyUnAyRkZusn6v8Xak3ndH7rNQ41YOfZ6v0BpRR4Vig
eUl7LYKaB852vigllGLXDmUIG1A9xYQome4Vs5oKl+7Sc8TPoERvlqSVEmrcgllC
W9Fm2joQM9B5eWC419vKaAvEnNKCM2nld4OYPuvMcfU4k57xiZs+NUSlil2CCVqP
t4tL2zsV6txd3ghTV6QfFTHDCNY5YEIDMtyP8wYEak9U+MNsdt/zW7HQLoay02fM
5NMyEtetIvWalPNfoaC6c/QKPbWIpvyDTQrTOLk133s8OppfpHggcVFuw54kNVg3
ab89eZJ7HBaxf8lEm+jaTBRqRky64JnLXsQIRa/Ku+bxhNaIPH67v0FbWFca0YDv
JCOT2cgaICG4pqEyw7FY0kg64WqvoPMU8i5OZDBzgdAzkLo8Srgh53/ZYQgOgk3+
80bKUmc+kYYetg5dZn4hcw8oEh6FiREnka9hMS3Jk2mvxQgC4FMO9axR1eygsMTm
UdzsqH402YSBP70VrwuAdsWt9GB8ThV/JeL0HZPeTcgko19AcV6jzU5uJLiSUVFi
BnT0oVjf0IY1i2gZI6vLt/OxvJ3cGFS46npM2xQFHgEiN+FiHNaGn7pC295RzcT3
l2o/mfGiqNbYcVNz5VsYSW6us3CwLSbcC7gRwGoB+tvncxJQEVTjRiG+HCB2lL9r
xSw2c1xZRNfbXyEXlue84VChBt1uutwDCzV+B/B6Ee2RNPwVuXGvTM/kbqlaMYRB
7srkDaAkgdf1IBGYt4lyGjlcQZ4KuLL3j1VzKS2Llj4CqoEeMu2kt2yF3CqbFoAl
zf10JA/hgaL79IaOoSbGhJO8Do8XsEpkgrLFDq7lJA396eLBUtCons1wQGkSLyop
47R6+SYXzqGWdfSvm5DTqWleE0ySVaJdXZuZAnSfMPk8h89cwnBDXsqgqlweb7nx
6RZ0jxMo8PyDmLe9VNUE6cX+UJ2w/X8vIBVe44Q/d8cTp/26t61tZ30qzPTCHxmD
yDLqyo5SZSEcdMg9zE3+K1pz/ZhAZ0fJrfBcJBkA8mp/67hIWLRMFfETZQDRhZwI
zCx+7/JStl2JKe/twj9ub8tJ8DKTZschpehXuKDkSs+ewjl0urlc4gzaNflVEc5X
VW0lbB4McYWXM08qcrZYsUcorP7IKQd5rmKaNFGmjpfX5161uMz144aOXdYuDTJJ
ZLdTGKeTf3gIZqs7KoSdwNRkyi4FVo6VH1QeY0dzC2ZFXB17+QIevP1OeDAI7CML
zy9wYwzlV4JewKq0ZH1LgdPtKF0HwdBIcjU2Fq9MP5IthveFn/ZJUo4+MN13b8BR
CKvE1nWj5pG6CejHGT1y7KBL7ODX9CqxGv0KXYheImV2Tle0gwvk8bLhdzvhdvmg
CNcbQ/4ab1Vbqs9BiO9hWk1FDdvjZqhbC3uEMZtL/3yq5RF5lpawDCa0gmTE9qwE
ALA8maYHtOuOdJDwkH7JGxUynY0PY19yf5ddkrr0zp4paKBdLbWuMS2Gxr45a3cx
X5qjZqNzFW7wE1Bh3u8Gt1chnJ54HWLqaE4IqoYAKsOWCgkJvifC+pr/ngrMkdtj
3e584aLU7MwH1j4770uPS8856vfQXQQXxBnJmWulehMphRYgDIJW45use20qkf5N
yqEntAQY9tLJkHIt8ScMm7oMuK55gT+epDMLEWX4zpVJZRrCHB/31GLtRhUQrheG
JC2C7B7ta97RHu2jKxO92ZM8GgX0QoB9HkJDsiYMq5UfV7RndkYHUMWka3Ct5Nj5
wgmiHnJ2x7kZEJ8LqSHvS0+9bQKuCQfuvszdiBMm02aGFaHMTABnybX8oXrOigXd
MYpDUdO0fHJ28zI1KJkrT8QN+gdfCpslhP7xY9sAVs2DxdraSM/4bVlA4K5o8DAd
0JNOoYyjkTgpjTi09RmriQ3M5OkHx3ometvbgXWS6C9XNo8uu+4EsulFrEw4evXT
VqsVzftf4IwCQUFzCDfJVGZ70o7HZ4ztigtcFKnwoxYSzHhIPBtZ1mfMZQc3/FCj
cz8Y2Z/grcDD3VrjdEyPdKmeC8PCiEtM1MViKcyvQ5z0mdPfsIAZpsooDZ5G9s6E
fwloHIBA6FWP6VDT/TQyTmoFyvrp7Kok98HxopnNXJoNsHftKFgKdMVZZINJ5nGc
N2blHfg5BQYwBYOz7uU+Or4oHkqWIVU3Kk0YPiIqYjAoqIRuEypBmNTThPKSVOlf
igrVDnPMG8N4mtK4MsC6c1pykuWCw5TFQ4vMFA7mFsZ9wCoz3vgMUf5VQPZkb5cF
2mF9RVsvHnfFEXXi6GJ8gWeIeuhzkadDHwgtr+TGqeiiSXgLjas6wJproOZVPY9K
ZrAUdW0v7oDPhT2E9/UgpO5JiwgALQg96FriP17vAk686cIdWypYgApxXwWuM6EX
BT0rcgjpDwgPq0Kqwh3NnAfA5A89fNQZCJj5D6SFHxs32gl4bToNpwqGRlTwdlQd
Ye0HXTMMBwBcJgXc0mrW6WK0AP+0f5PS/7fnVvCQI3LHg4bToKiNq0E9ocvcioNK
ql1CDTM0AUDHQ5F2RwB/SK54xv/XcwZ8/M73s5xflSRwpcEqEvJauYWNX3BfbvNK
yJE9JBfK/bDr1zXAdxZ7R5d4umRLfk14xcYjKvcN5GuqXq/472mn043Uw/088e2e
dH/thm/YVvUMBr4KoOKTtLRlCXayTqmjGMerq5WbneoC59MQuz8JO51HIFSm4acr
Bd3PY4FeOuevt8iPbE4OOIybXIuL0KXU9y+SLIob74E7mgkXLxz3AUSp+vYUHCKe
XIcA3xX6gfZ1lRUd5GH9aPzo+JZI9WhSxXTcmByfmHGhMOmLsFgWvZwuhGt5YTzn
9CvgusZhIMojCbZbrD5n9nq8Ji1Lm+BUSUQ8wq+YkeEUEndmosSswNNUChD/WE1r
t5+6Wjpgbmu/deoh23rAQAzCF+ErUQEohsNUfBbfafSXavV8CBRCAnLjFZhKbD8X
dbKFXLVuXeJlR80RilM/fErE/KR12xyLz8jh6JmEAx2g6vP5sSNWwpk/+JrKK6gu
jfJJHbUCmtti6LZRg4VfpmN+hTaEv3d5QHjTTxQWVudW2alCfk+znRXHf/fd3HQH
Cc3hgzBo1M6trSDJprCqKN3Ulqiz5fqoXBOaKCwflwHs1cW88bxwuGsqglQI8vMy
Dgti4AZkd2m4du+BNODMHQOLuaHAcu9OXuNQH51lms22CgA9j+QJ0YA+2B4CTr5P
gQ2XvwigOLEkAZ5SkjKqEH7B4XHkfJ/6a6S5FMXAdo9Ai1JmRNym1GHlhCiskxkr
tdu5fVs9H/WIva/oDYtWHuXSsz9G4ojfm9sUcEHS9fllZ0G84XAMnni6kL/gCwDm
U4bjYR0mG2XN106j893z8RaWvUdcHFqIbxth0l4/A4qfTW5A9PV4ZDQ70tB7TF5F
3c/MtgZUjeQTJJEwLCtWgy2CxK1DThXeAEumd6OWmMuB8FPq7mx7TPM9udnLMKfx
Jjux4Z4VHGW7Jz9+AyHR7goHEhJIYzVV1bQHMaT3wwdbmXldxjKmOaNZct6OgFpQ
ZzJ3cWHZEFV3LPkY3kX23dlNtZ2MqOeIWzNlDG5/3lPV+d73aklpgh3MBqd97gyT
NovAqd55Rh0u6bUihBlNgqCTYggYZN0X+xHfwi3M6/gNW6PiLySZl7RnA+pMynSP
CFnfzrK9HO7V7r3fBcKB3m++DC/Ezw9An7COabsweid0boOrwqxXtO8JEVP8O8es
8xxMxmWGIkp8YfpLY8RtRvOlFGQX2Fd0SP3G7G1dUUCENV/rTBZ6g4dQulmks/Wd
r7wy5/WK3VaBxkXakFVmd4Nx4N5M1G1jPL2ztCh79pwCo4XdSnGOX4R1JrVqkqUo
3woLDIbUrzh/Gi9tBqCIxag+Kz9vWrKLXYScf+GPi5tl7W4T6nlMc3M3UDNEfy4z
ANXVn2eBojkzZ5FtB3ecqt7IlvKnIjF6xFmDMX8nta/EHhBD9XO9jDxFr/Rljduw
dd67B96B23y7tFBQjY9d+C9jgyfuRKpY8B8iVzYXA9Mj02YQHD4Xid89ipOZAO1m
/8eSUqtQzjjPziUa3Bb9tcDDf1boW7Jyt2C3aX1j2msAEUraSA1mpFN0px1I5Xp5
rroP+obpRGKy4xDJSYdyHKYyTwwYkah7z2M89lczH2WvtXJTR5PTjGv1uyzC09iq
+XqA649qaPtFrqJ4w00WlvoRewEbw3VzYNLx17zHm0GYxaui+sMcs1ErZMO1bViv
4XuQRVgOqtco2F2VpAkjKD3xWI471a4fk4gj7+1V2HHoCWIjtLx5XKAzH3UXPeD7
HDLriBuDk3jlvmy13EcHB4ZpV5JMiIEcf3qMOeaboXulC/+joweDoj5NRj7DmNQJ
/nyXfUVdEmS5ekU1+PEM5q6lXkAckk4T4otu8xl2C3qf1/seI37R+Bu+FyXsXqZ3
VxZSeNLCICI96lvDGcfH+3BTnzHm2MCMCf4Kn/nwEN/vgfKVAHTPjPOlCZ2WQUME
JoqXFBIts/5UBvuynWpcK4b56ueiOAjTJ3mQK975AwH01whNPgVZ/Be1VvZWTpdM
tgW5QH0ikL0yrOiI/9RcdibDmgVjiv2UK/U6geTx0AAlGt0fFjlyJXCBiYjHOAmS
jBUP++hYnc8GZsMZM1ItniuZ8kumY7RAXWZqAsmasAncY6enljmiIHd7osVLo9eA
vV21j9OvY3ICMvhKXGTmEaQ52RcgrNIJlW13/jqiPTv62vmTywy50yltBH1rFT/4
EKsC69FGvymuKBFDiZ3gAqJzRqSDoHX1vzERM42f4KiAXhbXb/rt34NMf6lP+dTl
Hmddi7413IMWVR1G/t5UJm0tHVnIdyd7Jz7jLAJT5kAtT9LqyAT8xOp3h2/wAi0X
GjSSf2cmF4IevQXrPCj9lisqg+4w/lIHMWyMsrk+zieXb+GItrDB17wFq876YALV
aTru+1TQzV0j7w3rUAhYl/M5iConUkEE/xcpTzp6pse1/66fdbR+OAs8xZANSbSs
enjKWM8T5laH9h8LVewSwy8HN4MNJ2TfRdWlRe52WwSqXF8SaO9dEFWDjYch/807
z4J8/waoB4z5BKpNgtYCpKy78P8pzGPnkBo6on5J1GIZ8+M0QvJ7/NwbobvWli2E
Pp2q+UnURyPL0kdENaN7CkmzNZd0ix8UaeH3B662um6H28mJVQzXcv8fCGXZ65Od
m7iPfjlgANFbzzQM/11NvnJa+DSee08865Z31Q0Swu85cl3LIbGnaPFhi4eNgbX7
00aZRVUSQxjjRr/m5oBxwxQDAFajJ/hY8VQTYwWyUqP6/2JLNZsgwmLecl7ewVVn
jnF+RifOBC2M+4zmxfv5wWV6/8sO9oQIv1mCZkaI873/7+wEQL6cEdt8aRJyVBsJ
/aigY7iwH95bVr2b/TtRUjgXibcNp7YiZcCfCDbJ/WMAHXsttXvlgFrtFqN9JMW5
UvEcelnm4WbHGMKXmO9Ca9k6ura0dIwWuQ3ju9srWU0ovG4DYP8ygqewyitFV/Ps
iGjMx5vVH/AVxs5Vh1qg5pc3RJKgK05k62lfGOrJpiLrbcM4D6ZQDzWRiZ5leNVn
UqG/spny/o9T/hOzsBAGpOU2lcrgrAvtHwfVGc0eK30vcHV5ilRZf06E54ht3qBB
XfHrqES1jHC5wOwBfU5N8ZaTOmhlFRaMQPSIJDrqdJLFFOEgbjBJu5PTThfEFB7E
9zIcv87QuEmsovXlrzz0Lg968X1i+6QtDLgLbAjLp+MYjOYyjZp/QqhaeptoIJtB
fOKtotQ2K+7uVbVSCV/M42YbKrEchCSKaNGXRDxNLdckHi8VbKYNiO1kUsHvuRyP
HUJJ4P6Luz2WUyWdiCYGklprgy2UkuGE74DEvubd40qFACai7es/OBB0dnbs96D+
j89GjshJdNzEx0OtYYlnwCvZunrAzaMiPjws5OTcf4BYIN0silqVf1SEG9g1Hhrq
bHB+Z8wPRlZZWIdXqda2cwjebhlqBnxWmn29zc8ShDoa5uE0W3SWSAGtT3qkUFQ0
6lgLm+KhG86GRsR3WaP37yRy3T3LzVeeyta8v/Yrg2HvblgUPbdn3TDhz2bU1vW5
68/tOPbKCBhxq11P/en/vRcMH0dJN8z/7aWHH7I/gDzWEgnb0F5udJCfQo9dQ2zQ
4/93l0Lzec9smMG0bGO686d/rkeCvVF3qvVMIW6KwJMBs/Wr2hSZTnumVVFgwdwA
GC33y3FopZTBmVbxYC4ttFvRh0QEps95uuQqCVZwmyCObO4igS2h6Gy5RcXL2pJB
BSLDkEfE6FPD4upufx6InPhC3q7xC5UvAFKfidYwCYFs+GM9xL9sB5KR5/JgcMA0
MS5BNRTaJ0HGU33GFsaY+m/Q4biRDu5SBAaku7yc3B2sX6KlAgzRfKvdefqC5rlk
G2E3TPtdXDelJsP5amp7dQb1/KzlOfN0JWXuGzFvQ7qYbC/nwJVEynikTTGgaebR
HLy7ngkYk3a46GMpWwqdOQ/1NRWmS01tg/1SluaAWR1i7dKHSO16Ky8X54JmiD6T
MHu1CcI0PxPwH0sd4dpOHrIjySHvH1AfAvnopbD4+eF2RLk9nlWVmbiZSPE89p/M
wh2kd33CsrnU2AWMDUA5Nv0izGOd3PxMoizdh3QNzfNi53v4TxZ6e9jstG5kBxJ+
4cfJn/jGXt25ejN/qR6dwM1AzTHXOWMAHxs1x4g0xnZF4dxfzLa0PWtxvFjsblQI
oJ8fendEPW8C78IAJHjeJtn4N4W8qV0/kAPKmFbTdCFRjzTzKyDMSKEIL//uKGiG
g2+kLz2tIIZLr5v2pT4tzopxXCMlf7Mw9+/JOSemZjuMOGBf69I5kBsHJQUuoZCo
H9uu0h2D9+yA/EUNwzQDNn77P8koAAjo2L2Yty0cMjaMwDDyk76DcZQxdkolMnfQ
eRwddEmj0rb1M6X4RO8F4zO7EHPKm+y/tfbOHokRBaqmtG3/aXzCBHFjS+gEYzkd
CNO4EcoPZYoMwwNQa2/PdSwLBnOiURcP6kMozILWzWd+23XwlvhH7exwScjVQL9y
5gjsh0qttYnrESdCUUIrhmtWmHZ3PcblY8GGy8+3zOgI+45Po4ZVnryCGwbizZ8f
FMz88LdEewS7n3v09lU+7kty5GThmJEEaJ+YmU9d0105D/TvKvdiZfhDo3P8IcVN
VLDrEvld5X2ay0gEif6pBkjhut8Cl7QFF19/kp6+COu5fNlQmZzM/fwBCgcAgROJ
gvBUzXeNK+Wjf6RCicu/x3Me3h2DzrvRT1iAySidm8s4RsqOEXq94dSOjHSC3rco
s5Ir3UlX69HV/iEQoWnoPb45nDLansByDqTVooLytXGFV0fdLZwpXy65SVM00FYw
HhkhPhm4ANbLMNhck61/IM+WdcqL7Os3aGakZALDS4AJ5F81qNb+gtqXBYO+/RKA
r+P1Y/pre/SeNVagLNBINylVzFbjcGRLgKO8VZ+uHarKcktpRkz7yOT0u83bEtKn
jT4aIrSP2yfiLk45yTIrSQmkyRhlu/mc0agFYH9rOdxMeAv8KP98bttXfGEqMUqd
XjWAgFBMWju0aTooA03LivFt4kSA8PgQ7icRzej0JhwNOz9iIM+XRsJeyNyxRM2q
W5nNhoMXHrb26gwWXDa12LNwodXppdc0zgxuSry6P2sRyta0roQDKEuXHAcWfcuS
QKfV21x1UvBMuwc7Fx7EXKI1EgJfFih5TG39KmVeyxXcCFkbo+m2qhdR1OUD80lN
mnMgyejg8yrTmr0r7p9oqn/NMDi6yknxyOHcPgF+fxgQPKIx8Hwy0YLgvQxwwVaE
gs97Mh7hMgkQ6HAQ8T0ZjW4e4RLsmYon7zIlHpPEzy78vT2HM67ncO5axR/rpwJx
sg+ilf/DLxmZbzZqVe6okEY60U8T8GR6fjkzkFprL+7NcpOw8iX+s3UfZD6f0gN4
51dMzvTjaQggUgsCavnvkrHp/wK2NgJJZ9cEkrn4eWqsZpn/5MxqckdKOScsUl/E
MwNYN14TRW02kdqHJSqcqa8ZYmum7ygoh9r956G67mXS23BeD4jYVd/DiBt7sZI6
/E0T11581HF9ZoqIlZVTya5ostDcDQGmnHQRJsitCmTFWZmv89QWF5FCxREJ+J/E
ZcMIfnh40KNa/zAFqKSiKc1JsePSyCMST1Tu2fJQ8svhGGuSBJ06WkkcdKrstvHo
vxBWwdUNc4So9UKOqNNpYu77I+pgnQMqGG4DppQ3EcAsEn5mJhfmLVu0Ikf7nPfO
tYb2X1tl8GYufMpssiWnGVG+JrFxOztJe53YO67hte35uikGUoKFvxYdldnvfczF
tARjdDztBtYujfZvsTyZIw+c7TBBApKpuiMkQ47WmHnZE+xvdsK2WLIaWq7XY6GW
Aoc7KCJG9BhNXFjw9kmVc5LKgTfHs9mJWkk1+9zkIpuRmkBtX9VbDukyhGqMeNEm
6aDDeWyS78SUGfJDpg8IG9kXYD+Z/bunV/jC87QY2PBz3tVYSB+fa9wVSA+iRltw
mXeVAdw05dXZ/HJnbDJeFHBS22cHdZZWSjRZmA5JnUedbE5QAMtjAobDIi1DQ9/0
demd725SiwQCktaJS08wWhZBboMEmD/kMH1UlPI0o7QAmVJa8xzsfc4Wt94bX6aU
FVMIwTZEviGcBO/9PVyMl4BsxgDm33s/BTWwjJ6COfx3qb3N8FgxxGbJSnUc6HuN
uGJHLEbAFIruH0NMX80e0mu/jshfVQ4scQZ5us/3CeXvV9t250WeaeS8ax53e8QR
UTg1Zk/Njea27afRIaHAZ3BgG2bM5/1PefRquUuIuRo6AC8ke8cxOntJWT1v9E8s
1IAsKgsNII4qDnDN/aTEBzkeTsBE1w9Ezf8ts10TYCDrjKq0y4K1dItyhrTZagph
NerKVg9DavGnXLM8Cdppv1+sP6YjFSEHr2fsHNWfNKU4xZwspuEJf9taZ4VnEpzH
3PSUXwHW6G9VaESTE5V6clw0fcJH8LZp5KGX4sKsCHL9rhlDkbFJAs5eGHdlihQR
mPM9+D1/5QG4eEOTl3Dc63tEKXyPDcFW5pbJmZDMdmHH9zkyYpHB77eQQGndTPI9
SrNDs86Je6gIvf1bt72//Y2/MdA0Ko0c6WUpt762LbUf3GNUOdhg6OGbYWTnxEPb
xspqHH5bgLW5AzDLEvcfSRJwBcozW6K5nj9Etaj0DJ2j48LVDYt7TPjTqWx9NZoH
M1FsBgkuXkT+MxwsJ2zpVaLd+ePamk1FiMjpTQIqt/5bd3pp8rIqNS94wbP+YPvc
82K5hmC7q/ygzbfbzhxNd6ff78j0lq7x2IAVN4I1gnmi7Q6OqC18sYyVrUMqLdl/
4v3aOZxgQMymkM2iyt+UWcp1LaWU2gGxcIFg/Clr6MlWAbBvt+x39SbbrwTfmoge
7HrQlxNSVFmv+40vDNCAqX7A0V8zKGT7jIJuKXcRDsxKCI8m1VjnEYbxlxQOv3pR
KLINYikEm2ac15wqKp26mj97a2zwCu4C6E95HL3Fu8l4QDGUQiWAo79iZ+cB3lt9
jFIuF1IRna0lGJWNVW6fZufinU+CT5A3xCELwQN+EqMqvRonX7UgSN/sfLklQ3DY
zGrv5+Fq1jZkcS+Q3PcMZaFDUhH7zmgtfJ1l6kE45V7+X+lpyND/eCqGJ9wZM7NY
zsxW1uEI2tlStmVACu+iEjZ1UQlo7XIqZwJT2NkdL6/BX6aAQ2w8OSB6n/l9jICw
jYUn2JlGbrBtiA2q/a7nstc2NZysEBH82LMpXLZnfj7iroty6r7bMyZuV6Xi0tfx
5CQF/4YeFCYlG+0/TSeLSsowQCuOgGUYrC6xW6rbpw0f0Rvowsn9aPGHa9DOILVp
QNu0FvZqR3DvIPddfse0moNVYZb/ycWOLWr4vuLrRH9eZMRX+JwvmgW7jBk/vsz0
vVMtsHReIdpIKpnFbDsaT2S7IlA2xthnX/A5UfJoUyWW4U/VBGDdEEwkvdZ/2NU1
lIS7QXJH3tCR5NMIVgDo1wK4KEHOsSRH1Bq4wcHd56LKzzfHTcJJLpYGNcC1eL8w
PIMeYg+QEhynlwH2Ml9TrxaHJNr7h32JKc28OtiwfXLijXzMvwCfEYRNsprVlqKu
D6+OxqZu26OzWCAZkJOLaJXyK8yICQiuXhQ7GwyVkxA0J9OFOb+6CQRGw9sdDTnV
afY0svGiVAkVDU8FXQ/5LwR8KKZXq6b2Sxgpoo4eupAX3h040qKAWkifvqZJe1y7
m94/oofVS01/1bSU2rLxHzKdGRgVnT649JasMtHWCa5/upd7K8n9Bm49mfR8KH7u
hVmLwWtfy+yuf/aWqAhLaiBWIoUJggDVg0EImBMxtJj6ry7BwRYu8/rSF9TouYdm
n6zYpyamBpktgMCe5V+wO1lIXEby/Hj6uYFo9SHwF7uP2v6rbRBrKLpVgkX+6HNi
3BCgP8dFEqnE9iOKeJv7zZw1EexEWRkaim+uafyqXFbwW18b141DYw3VOqsy4muD
KN2LpFmc5dlfN85UvOTCzchojFZEdvlHzjMEWiXAuRoJ8jS3IXvt+t1ICxjO8zV8
+8RgbHdDk9M7dqtKEY15aidbU2SzEtozMuh/CEY6ZYcArbui3N3pmECnPlWr2HUs
HsQHOL/rASNQqjlUgf1AFavTcBI5PTJpAuZHrOJHpRVtfHujegQbaXJxvB/S2Tc/
X21riij8Lw6/8vYddEPfCuwj9ND3IdMO7FlYuHvrY3P+yVPvVi3IpxBZCO0dhB7i
rDgmQjdoNP3ZyK06EkNCLzjgLLC4DWBoTfu1avKxaOMVQZ1S6h1ykKM0qT6CYnF4
4KHxiC+qHjoxPvA/YInF9ECWFOHLaW8Rjhkv6KwuA0FEQCcEFfxx+mECPgQWlwWJ
2gd+R/CZRj9VwSKSN3onDbRwzR1hDavluHGY9mSLTPUc2yLI/7ZDlAQKJP46Ra0H
ykQe2EIM+jPrvUbzYrtPrJ7QWtlRd37HEQLfncyuxpR3T/35NEg2znKfF7a8sRVy
KJM46umMPz4n9qim1O1JAh3SnGPN3wwH1b1lC19ya+TkDpJJan2FpQXovemgmCns
PabYCnX2oko5XDFfRxB187vURbxET5DEAaq99lsy1XJuc6bfLvPCqGLOGoxwee5t
3KD/AKJSJQsdd2wpkBp4h+uYDKThCrMt3VbctwJGzYhgq9UcD0skXx9nMSa2oZNF
JLaBvQTDEZ2QdGyWeg1NM4mu3GCURgaeA4jtbXD0C1UywgskfpXmiXOA9Ky06w5D
KJFrlUxaEgH5KuVlVPDyjESkM9LNYV7AhuH1zJqfBSNHPqES5b2B8FW8xxRj68Cs
csDqdrNs7uBj+mpBitcSf9qO7zBqciql7RA2PeVyppyBLyR36Mi6NUxhdFaOlxh5
iIiYO2m3Gjb+6DPuzd+iEiFTkbosENyYG+CdBLVp/z5hNLd384RYT1IgmBbCmitT
ICF2iXTfN1BXp9JCan+s9zFZB1K5zUQaXiGb4N/3jDkVQvLAEtsMlg7vW85z4bm/
de8m8QZri2VW6gY5kBZ6gCsqkhErs5E9sfd5unuE95tuQUHIOuTCt5X/CVc3tj3w
wXWB/q9YCa30eNJdHrKTkjgzChUYGPMhJ81GmOTS4v9wHlOR3kVDHV3XdCtp3knu
n7GQA0KOf5B/VvUbFdzW2MXvwgF2rvaIipr44k5Ga0qTAmgZWjg0gdoHq+d2HUWg
ODp1hz9sy1AP/CoA14433sNIx0dIBVn/V4VsBGqW2Bo8zh4mjtOtzJYmuPTLvdB7
cfUHnk3ehEwB0gKeKGiJvgfE/eVjWvoPOJtX0XP3NiEIOW8bnYkJvn6YNFIeOM1Y
hsGwyjfMcfwhkC0WqeVMbxyx0jG0dUzTLsRmuHUCtqCOn1XL35M3cb6uQ7dztOG/
WIsMJaNwBWsIynZk1d/MOjTxSIsBm+JqrhwNZ/njn82QRIVrGYVbX9Tpi+aJSNGX
4/KfeNPXUmbgTIpJcKH7/5GSEslUKDuEXP6oHmok4fLcua+kN4HlVquuicIUGzHt
NDU3XJ5Gn6TaiRjrg3ka78DVI/RQKJDEEOK14gTW6IGvo1SdnwQMBcv2cxfxtDKp
tASjw7WU8YfeSSVvel2N692oPlSFu6b0jPutiEr25utLGVYwF56Hm/0nwSqY3lXx
/PHBeMx6QdVrBJPPLk8ZUJ3iPecBGI/rFkK4tfv2C1JBGrQuFvd7o8lv2GNm/rJA
vH6cDeQf4i7cQCsMeFGm7O5LzdM61OTn0THWJSVb9s+3MiZ7mn1giDwfAEJpyI+8
eBsK83eVeAVfmsFifNxhCmI0QFeytDjwkC+zj19vY0B5SNR6MBgSuctPYXpJdtOG
BZQXxBAn5xDynMVF55F8xZR0cYFR7hQcR0yVh3zEtbNnuJBY1ePAGiqkw1QbpR7g
6qB7BmcM23fso7B5VqQac+6Z19pmjAKqNugfJir4K9CiZZ7dnC7j4wtzACotdGSw
yNkdY+HgfzulFXMbI9pTlqYxESVCLZqwyYLxK/lzEzUtdb0V+Xn+hJ3gs/uaSsiG
iLfHPH8RmXnyOooOsyf6+aAL0DNfiTSZPzzsP89A2sHGahai9sj+5qBDR6FU0mZp
LidDMxlus0fhyXcMfko/pehC/+ofk9G9pMv3KltCIcBUiIutP60aJ5fPIjLBKfEM
7UiHomOeMnBNKtpAjJkbOlXRetjvfd8s5LsBA9OXYKawkj5S+dQbCLgYwEmxfyPm
WKp2Smd+G1EWajuVPTDVP0hsaH9IPwTg65rnYYo2oZFrYjWT+gW5Vz1oJO73gZH8
klQ0i/kcf0toljo/N6TuKpKVD6nkpAGzBmE5F4vUjafX+hC1nWG8gv5xdTJxh2bc
mYK1EEtrc056YDWlOzDiKlkd5vUMO+j+3bwFEcK5i8P8Ty7GiuDhCGzNTXBbrwYC
FLfPwbB7FdubE6eBjMuIXH9ulfOBPaIixyylHBvydU8RcetpJ1Km/gcZ/FSVQK7m
JxmU+wSF5VmQ3uRGbaJ642BKzieBoKoE7PkuZ2NCGDQqbdwPEm1ym+bQ4Bn6/blT
HfSXu0vvnD4jlQPNJHz7RFPWN57YOYOPqAq1WiGBNpzS3ZI4tjuL2oBauw8O2IML
U7p6OZq9/ccPvJ6UZoCu2tydoDQtudQHqWCTGn5Q16986aQWDdJhOvQN+m+5ZOB8
qRXL5P+QfozzHvsPbSjPRV916yWeM8CEE+1ISsSi5/ydhwsuu5yq/SYmWrG8bXmd
LIfmUJrix7QulWqz8kO8oQhjzQ9pQWf4gHMxCTV1khnrPpZRnkB9XJv6Ld0u/7yC
oBZqzv8YsevJFbCTzYACRJgHR6mQCPWPVCdFCVR5iLUEs5ORhIr+1zrskdxXkpno
skuIvzLW2NMph2xk5P0xSKBiJsLWdiUOZFMsknm0MIf7eg1y11L6GkttUZYyP5gU
/oqOo/v2MHU3ey6M1mPw1p2F+DO+8b1RtRQ/+8AzEXX6dwNNmCjywpFzM+YVg6G+
DhWorqoBDe31S9KjaxY5gUFufeEl45hc+TDqe2FtPnI4TVBDXCpS/zWPBv06UdQ+
b9BnOLeVT/NbIiZkCrGvwbu77TdhkbFYir1zt+Rw7I4LHOei+3WZWQeEcsIAuSir
H2FGDG/xIIirfUZgfGq2JJKD+jFa7auOVwgUujfk5StLkK6fqT6n3OD5pFO3KBm7
N9bi8KXqrkj520vJHq66DTyhgRVH1hvnbXnySaroKRUdZ3tqT6s++VeliZAxLni5
vwzJBFqn6V2JXz1PBlJG+C5vI/rt4jdwpRIEpZSFMxNGvSrgna2YIo98m1ofZu63
0A6REv2VANKmuAXIHlkGmxEX6EferGHw8SIRl6qsA7sQg7hDRY40YylBdnt/NFKj
pg3MIs7XB/zFX+oE0QyhxtOUVnI411AZFcDnjQe04/chb8DaIUsv7wBnsQBlclIg
5gUIAfYI855JUKdhE3ZosC7vZbuN6Qp/qTITr7X3SXpAhiIHSJ4AGyjzG+wO6MTT
3IbYHkI0DgP8MgpllKiHIRZHQCBB/htZWVlI8g/JrCTISD3VFiYfwAyNrgZH4wbo
fPUTm3VZa+PxAFBrrH6y0Z0N2DvOyAjAMQAdBz+WVqrOsdYisG/yJwZHQKwQIuiJ
XpHwG5QJLiICewPZ5El+LC9G9U/U033nX5hQF2LwZodqOw4dN0CT1XkfFUPPOHb/
PFiUr6HLhqexSqB60PRw4cdZhsQxgV4aRZdWj5K2AWP5NIxBd8xxtCnQ3sOP27wD
m7xaMcGJ2pUhDE5mNRWe5A8nMzxZ7C5c6yFMBlDvefVtFDtqLn0eq0w2u0pbLj4t
G1EUOA7nhqiFEPc84dMIbdQDH9Ay0CnhzyL9aLyfG5M+JM8maMZefoH5CrNBaV1C
/ombs4MxR2qLRZXQ+DS+OVm3BytgrGcva+Vq7oxHgwU8iK7XWIen81ljS+TZ8ygd
H0DL+fjZdVhFC1ef1NrsK/qkB8x4Hj4a8t+0It0wn/W6MqEVgOCmGHq9pNMTtPuC
gQ+6QhFqwAiq1kgIylbnDAga8Dcz8N56tHGgsnEkDb+vhyeC7bHZlU1pjoxkl8CV
DtEsfnUoKPz6rLeorDJZdzM8aKZzDNA44S8b12qT3FiUE6I5/H4mQ2oo6Z64W39t
0hFuB3xLhDY3Et/PpnX1IdDvzMRrxBxc7WxW8XAhEj5M1/MXHIsL8y1UQRVuQM5j
GYmq/RiibSbANMWizWvP9AHt54IPrkmDRokk4UNRyKzfDsIIsp0YCYztKya3valx
EGkDPzlnZof56dqsHVhnIouYv7yQy13+o2Dtc88ybw6pbFhV7reVexj94D5QI/Cy
iQzf/nYKVpehnJOmbQpnBuj2ZBA/cFlgGKoN/l30jsJZf5gYQh+jtMe3AEzy2K3E
tMgHgkd7CAYE1MBgWtZNLYX5ct0GXKoHPiogulmQ9C1VXMfw07ABxXQJT21+tZl7
tOX7zs9wq/fxTBfLVWHB5BfTv8lO0/Ca5OTFNulaa869xfdjwmws5A1uSKTDESUN
pD4i0P5wLvPBooTToIShP48793DF6he33tCGqAbVoY3fIT6wMwHO3PUZpFGRFE1l
yXuL6Cudj/yVqav4HHchMYP02oNyPFnK5pbxvTRgzaY8KJ4cgAHwu/585Yxs5eD6
9LLIqLQ6NmPqLxViXWxcCSy1gmcDuQ28LDGJKmYl1Qo7UAhjK3TQsC7EfU8dJJQ/
vxqgfLOZZv8GjLhOIB7NLyeWhE2JC7S0yZuhDYjaeP4fTZj2phQpA/3VHh5vlgmW
uMF3GM85PrIVFm0VSapGVNULsVFXFpCnIGMBqmbc+e0FGRk/+3CluQdwXUBiEpaO
IbMhS35Fa6trxmkWnCHhjZ40tBp5cuaprg1A70JOUC1CY7Wjo/QWF0+8Feh7Qq7R
3+51fev2O0BbFUzIh/Kzotr/pU7t1caAN6x0gMmLtNHu+FzqrMRzJtoP0LvRGE7o
avnQBY1CsrTzOPbaONq4wboM/5SuMmSvLPr59QUM+742z5zwLUGw6Rsjt4U+23D2
754OfV+au/FT5tX/E+sEqzXGFgPwj+ta7IRkPljZorNN8eV8ltBxIfJ8QhZRJf0I
T01o1oZIYknosAhUVJzI0u4Zlx1UDYPT+1H2BVRHvA9Twb3vwfTheZrjssZxmPwq
XaBr8dfDqhLqeo7BLZkH8c7rWZWWhcBjRRQo1/8O6SiC+R00Q0c9gReXqRcVGnQX
jqzXrhENky51QfJvhcgDyHFY8YFl4GpX13+omPT9hO9BWHlFbtMNGrfRCRjB7SSk
AnA8rfK7cQN+uEHAryxtPDMdG3vVHse1A2NVDN+ojdkcrOzskqX8HQ9sqHSuurHN
6eaY0g1HIzdwJ63bL+H58WSZbit/UHx8oX5hBiwe4YjRioa3FBaB1CzdWVXBin2T
adpM6rPAa0cHx8eC/wc+h9YWEJFnNOji+Y3sjeL/T+ftF35zrHPZW7NKCOVPkP0X
JWJeHu4n99wE+yHSRpQCgZBFBH/4nOipq12uMhNUlt1nZXDBR9nSkZ1QIVaNrevl
r06jiUVRN5Xq0cJ05Dtvi1mUJ/MgMYOaeV5tk+OXRslkb+KhDWJk5C4X2WUwmvKh
r8/64Fqkz4r2TLs+ftn/3Nng2+ajaHlPdVIjDWL74Lx8GI7CY4bPXv6IzJzLhaa4
fMh8d9nmYLN9lryHGysEhsuxTFtqN/GEL2wse5wmjm1eR26sTA4bstXVsMHbGgfv
fufA664qtiku/hP0uwXQ9rg5L751Hkb6UmSK8KOOu/tk0dBZJNeKAqpvZjQLjv+p
L9KryuZ1QkK+6vVAmIPprN9VcyUDtJA2YpUdrt0XVoEuEnk9DVMK6nzJKKwOWrxJ
lL17HlXXsy32bqqb9QZV9xI2KJRSh2tCaNfdagCed9CNBBUHLInAl5mXhT5nrNbK
iqdKQUlR9yc5oFgFWAD/5uvRM/uQmPFaNv4QzVdyX3z070NneLNXswd4sjek9h0k
tqtMWYewQ7dNUOr33W1LbuyFRXNFb6gpQaweP+atx0u2iMwuWuvjFmFjjNxFzQ/f
QpfIJu4/bhvWmhzfRW1XmGdzXU2VY6EpPABeirdT4toOIoIcWEM8hpQmba4F8tof
u/fBow15ZaySkDNvjLrbuOxHY0EITqICmixbVnziVA5xpj32nhRJAU7/33jckgpo
NhXldZwZbyrprSxJcdO+9A450nQjQGPoYtEAWbQ10oypX7RgveWfQrCFVQVy4VBT
/9egzBRZkTK3rPP32lrqlHhktGxczj0JpNpyTFzGsdJvKD/EHbxrxNOGEHGYjvPu
Ss6sOidASOP2xf5bNW6ws81fGcmqZ9sSZLN6SOjy1Si/nQuj3/uCEQx0KO7RICdf
AGc1naHyoJLIGOhiTv2pWbXwLgBEQlC9NWaylVFk0WQ1MQjPx+EBNSYhchsJiRIL
q8XMe7j32WDRZ6qJixXjm+ODh/AzieFHwyRmQyg/ZG3GB0kmUQXV98fUjIX8wxI/
mWlN+bh+HThg6nyOkWwZlJIClfDR0tZr+rp0xtVrGQ8e/6fRPKu3Szyh3iIZPXc3
GmFC7CDFxtFp+m2to0IuoxL4Bj9xbd1k/wiz+LjjUgu7SftYdb9nu77CEbwGAga9
9cJlKGwPdqkF4larhD0I89Hm3XQIid6ZCGIrhahl+xDOfHfJAhHY6k3P5eyQOaqs
1rMmJk7p2LKT59hZ024uYiNeiRKiNClVdGDjJJzxLbtiQ7yUcNKHgJHSjBXIEtRN
inqpvEeP9oDMzqEzuvf0k58U+yE3l02lV6f6KuJ1lwce01+hMm/MAuvfLTYwdcI9
guZd8KkWYIUOubzPX3C3GupK1IqcHTf2u2gDqy3Kc8iVsUyLRHftXrt9azyoAmFH
PGAaZDVmCrw54zvzN4z60NgAOoHZuvXpEDic5XuUPhFLBiej5g+8jrLYKUD2o5mO
Sj/rYrFTS6txAT3lYLUC1v4rL9KIqI5Gt4zaLwgjcUkgNABc7oKfOZLM/IxLWoQk
QvOggU5aaDbelcPT2Cj+XS+tDpINx/jot0bxek9YKgP9EwiTH0/e5M8btJ9fE9+/
LT8sFAzWYFrOL22XR2II59te8iiElp6pkhO/JIDAtOP8wpCP9Vzf3W1GvtiJp8CX
f+01sQfqmxPkShCcnyQahR44UubZqUU83XjmRQXyBZNwFFzp2gU51rd9Xp9o9Zmq
O7HHqv1epX2Po22rYlti5U/srDeVBT7lI1FyOGMHzdI1w17N+ZtLGi3YD9upoOha
kiY82e/kNTr/1f8PUyrgS7bDXLFysmYseXS+3zpXuZAtLXMhLGeWr4Rtwjiflmta
NXlBIxuxj88a1eim8dc6BeG9moT8JSnRXobDWxrWr0W22s6HLwk3KjnhaHo/NiuO
fNHAMumOhLRRMUo3oo/91uL9LxnPR/5QoNwjoPM7geTLoUEooVwXOSzxEPVOw2F+
TPnCTlm5Ms6acdAMCCLAwnqNrD5082qCIFIyxVP8JVf3IHd/n7S2/xCh5zWQB3Eu
yPrYXKwb7kJ5ZVxjiGEVTuxLbquLF0SsaZ6eUh5KANEEH47Y1hvzbhnGHn4aE6Wr
CPW7U1lAkMA+/GaD7v6iCl49Rqt5WWWeAY1qxE2/BrFnmjgDplbWmxCzMBYbch80
l9fM8QMzwefDQZOF3FrJynCoSsvg1dZT9TgRwpU2yXqvj9pQemXqnHcmPtyqG9Sl
waYGcY+mpciaJ9SXuuujmmJkGMod7Xx6++Bi0F0vxvzRjdTIzx+GRAZQTE2bNoI6
IDOLThDnjeJFwVnhpOj+XLLq5QaaXid6a/+gdoj4C5Gi9L1ONMOYHxTO8oruf2hh
WK38s/+BqWObZS+/KrC80UYHHj4g63f9WGimKHe4UGMY8L37DAJbgG+O8o6C7eWI
q2Zj2rNtF4hRnNmsa/ejJo6q6lKx47aQG6RGF4gbbgD28Si5W62q30b1DuLWNqbv
+Hj1xbmCfVMu/Eao4L+0VQmtFRF4flzSi4qOPuyQanKgbSZd66TNw/YZ7Q6+wdw7
r2Ab+WAUEoZXww5ZVsZ0hEEIs8c5DMPqr5LVKJ9EeblXocJEBjJ2pcup2CeUEPen
OLsyvIncq34gphcBG0w0gyqCxTZbAkshNZsYBkdEOWtdLUwDd+XO1L+lbLuZIc+8
2KmBL15xG7sICQ1JlGdv4lK3GI8O1uiJCnXW6qmJK+dWfs4Kekyjl0+0iIG5ezvR
RMQ1391cYUcZtBg0/8/CcE6oVLjaD9f+KRH5duz4rB8vWnrxnTSa+jfQ4q0dFUMP
YqhXZt3eox+4HD9qyVSGHU+r1HcGipeoOcNs5X/x1SjcpacKBV5HmjTxXxVYbIRs
80rB6CExNJeW2fiwI7DrfGy0Rhi0vW/o8jwlbin6UT844FbcfCd+wPlCviBAPbIv
x0r2ZAElTBiYeSqw0gwz5+hY/3Co+FeeIqT0gLWoiILEPbhKHN8ni7dXkDv3PAuC
aBE42EWH6Sq7hSyzJjYbPy7hZ6nDDJT7SSXIcJa8CTOHzZrpgo/i9uyh9cCvOJTq
wKV3EeL7KZWrQ8FjNBjGI8Zy2vmRM7sV++NLTL5Pk0DxNsgsHWN31d6BH/OuLNu0
y3Axu8lzYS6yQn70Pl3lnwslqJvaiKELYlLiT/X7z10BldG1vELKs9hfWPCjhYQT
m1YshJkoYG51pHukh1okFHSrMNHztiD1lEgFLuZN9k6ij3PmkzfF6XjUqEWbzVO3
pxORB5F7mRNln/iL81OEjLIcQNFpxcnxoDGFh/V2piyKVZtpZISABO0xyUeqwN5x
ScwylVFU5azIJtlrVEQ5E5BgOcwO4DtKDCjcBanfMR2UqXsx3EvRZTCmgsk/urCV
b7JN/GTcNwVc1gW12gzh6BY4D40kbMCH+PTZs3B3K6w6uMWKIIIdNhbwUMFl+FR4
saAPjplr1hwxqi47Xo/+tPpulSaU/LNlwyoYOQiiFoImy2msyDYRJMGSX5yzwJys
xdGufTWU0YYM2nk/7SjpnJqFOS9U6R5bFBWx+wgh7uBRfTxgmswRpNdjXT2aXeI2
j53rDpUZcU4hRoucXL1OsWnVx84m+9zeQqF/MgFbKAap3ltjitFDgGLWCzvkv/V4
R5YQGerfwsPojiq4KNjnXvqZQCLkW6zkhmeAeCgM5IqOgIfxaAkhnC/c4h6K0n9c
abHCOcUxBnnB+2OWRiUmW2IF/rHIxtWShvh4pTMfg/ffnWcFN92GZHgqa4w7meNy
M9KSjB2eIgMTEd+NHKQKEE/wVhEDGK9MYAne12II7RzYE1YJ1jFIDek6RGkMJcLL
Yw50+YVTIQc6eo0T7mtkagY8Y8hMP4k5Pch2de6sxuK3AybCiGjwRO/Ikpz1Vlf7
RpcGwzRHWlkbhCKV/L5dFdNudAg6D6oIjPMrx3A8+8tYaDs2RDqIRhBlvClJTxb4
aKArlCncuLLpj2vJSP86ruSbOeIYyirfJxsV3D8goby3NGhBUeI1BMsCsDzyI2oB
DQ1Lj5Lz4SVmWcFp0fdDbshOwHEHtMCdd5Hww77Dvhu35dGy8rKYIlLvo9C17/Py
mxJzzeAKv/oL1lb1ldc7QCFZcXpHgo4aiQ4r64294U3amJHeyIc1UVcY9+lDbyB5
Tm9zSqmk95cv9bTTxNCz1cwtRIMe9KyJq5nWS25FNewNXqVmbRMB/n45k5gn5Fd9
IeDUsCNSeXHqxoFaY8qlNehTR179IwCSMUhnWZGiMOWicNGYz1cpHMCJy00DhbKf
MUcXEpzhNDupgZkAtNMYrD8d1Ydq4VRLj1YMbJ/sXCwQAfAajNuR5TsikZsGYkEc
7DD/RRtvf7BOJtbP64XPWc6271ElbfDQleLsGz70Y154v2fS6DHOVdQ8H64n5GZ1
EL9jedmsO4iuiQzBa2YOflLrKmP3gqXWBkKbtrqY4lK9s1j8qPVGlNOO7e/rdcCd
SKc8w7S07Ln0nVy8Tv7+XpUK3u9/9ssIRDQ8PGP7JnNd6m4XfhgeSw9YToHJC1jh
L5e3/J85bebodnfEhPAI+KDYYY5rBpE+qT3fghQPWwkBONjGthE4I+zXHKoeodFp
pgHvasB+xNsgVp09VrQkTJEfQuCGsWH1MOl4rgu7fJRa2zdT2nhSR3GTm6xTnrke
nWpv4IeXL6k1hqq5hP+quogSTjNDsHF8cNusfyv6r3x8pfaN9KNm2QoI0BuskvfD
Y+ZjaEbbd8ellTlUfGIfiQobdRZbLj4EGEJo2zqfTdQTH8pZODByzfW+QpW2uUht
zxl/y66fPrkMJwxomEMFF7l38EoxSM0dbNRWdf8yNtTGFnjyC6eQlbsGja3iAxqk
1ne/ZuDfIdW9OnQMFN65kTxTdOvQsfXYhr6/TEFRze46Ig5XZAyHsJIGH5r3LUhm
B29uXV9YI4BpypX1UQE2n/iRW2T1dBZG/OZZBw8YdVy7Ia2lSmtME0hbR92ruN+N
pnOHoYqqRbZ0K/UMF84QG11Fzb/WlIaH+qLaY1/sMO8q9QJ/f9ri3j71LxKXYYZS
D7lSVYt7RbToH5xT+PE3RrfYzg14zemLxCm0EMWO9eySpR8QPHOUmLjdTMmPbwBy
m8QXEyJMLIKXHPLX6tEyGHlrjbDftFK1sgr/XqKd1o/SR7p9hj5Tx4amIkKYYhcB
QJsCubnJeRDZ63SD90GCVHlSVahm78ksRRwKhc7oIAuZBMWPUUc7v3UHzoh+74Ab
GNS3rxUki93EBIWoUBMVTtBPZi5gOJWJQiO/zgQYjyES5mYwcpUYYBUVRxxuK+lL
mrBeMnBtdGXQSTFaNJ/+v1irKWXmwJqiSX+iQodVoMJCMnAJpFCtzkvdQZHDFryJ
mdhZxcHsbSSDSI6HYkDT3YXWg8YeZk1u8TPFcRG7nFAbou3iyLb2goY8R71YiT0W
JWUB0teCtrq7fHlwB0xh7hVYKk5mhSi2bQ8jzyuwPWk6m4VoKca9RZqs07MaBi6s
/Ew5cR4VCrRA09jx+tRUlUtt3m04SQ7hVkUe3nl1zP0IVt2AllfETArWQ1fTrU/w
fN1DDpNPFuMbQB1sLfaDZ4lYWbWPIcXG7DLrbGrzXzw+SHnG3Qvy5qjIcIvWuzdA
UKEdF5D2iSSGBVAjpmLPBKKaCgPbFs55gvil+elqxMzoWOTPriC3jS0acAIwuNX/
HiBfXuAblgYq3KqZgtfbnCnSYBQbDaEgM8wBlGTbS2d8iAZzsbMOdyAoUbk/Kzm2
ASY+SP1RbaM3M+XmyhVJblJ3PW9FemH8l1JFgDpnV5ZOXJ38Wnfwzp1YpyWGiykQ
NiYPWtm/T7wnyykOmw7+oxbqk8pXjuGPDG1cCfU/st5aw9irxByILDVdh+jPIlcX
otoayi+VuLwtQ13OqlNR1PSYeC5eGzO0nH+DmiWnVTsoKJVLuLIo/LMrVciEveIn
xtemFX/hkYDfpg/7jgaLv3jjQO/n/YXDXrq0lvdNI1PIdDud6DeSkM3lBDCMthwO
uauorEst+8Ob3V3lh3SXFyyvUtnGUej9KYKWGihiIafW648gN8F8Iv3sLNlSZ736
o6ppkc2XGoq2HrXDiRSV72N32Uf4p3pRecbaNE64tKdhgfw2l5COV+qtZzQs3SWL
f/wzn76pLYB7vVRbiiKAKdpPaZIg7Im+Fb4qhAKMpr1cdVPz64iwWu6MVWJWgI0M
EfPkmbtNb3111307qMWTTbuOh1flk9XmBIxA/cAl032e9MNBXjZzU6KcZJcgK71g
O0w3e/aTF4Hs7UePX7QcOIupqkry3VACPLWnEfbWB51cFdXNHVZpPDHx7pYZdnLi
V68I8SdfU9Q6Dyvwfc+as7qixX1cDJNJioKGVhGVUV3lB7umy2kKLTHCiicgaFx1
V9SfhCAHqX90yKHxCHLB17q16O+YLYDznl9MytdN1ifrNBYQYSr0WE6ymfBcmsNt
AFVpDvx4fpxs9Kj9Ah4ATNPLu3Qf33IE38zW4fr45BYC0AZFMyegwUgNXq1tTdcR
9XZ4wQyB2K8Vg5JOG6sdJA3cpMKSyU0rZkV3Mu5BoeNNknvCF7TtSfwt8DqF2tGj
AybMTiDywx4bfZ/wiyzTXo0qUzdkIac8PqiASN2F1DbLWCPtqBZhbuXiMWBHpPAS
W/jWU8MN+kc6FGuMEZ1hIWdk0yfxHEoQigUBjdkYTQv7KMPkODo/RInLAzxSLtQy
PJBHtIoyR8owONKfKmZ6W455B1XfEfqjxRtii4Z+2ENxSnytjvHZ0cXAvm6TqbMN
3GvKBee4fpB+LNE0+TSggogGoWzcWWgbNPrFZnlp0pUqqQGRPLUlquW/mnq7YDjT
WGw4hvpqyspjBO9Mm5vrFCw4DuZWMotfHOHg3+5Cy3VjZl2BOmv32h1YamuVA/Ud
V2CiCr1J8Jajk/C+zJClby9agWzG8u0FABCr/I8rllNXss3BR6t0045FTT+r211B
SS9E2FCQpz0MBmdsrRSGBZ/HA5/EZV+gytNutNh9x2yuRdH/ErKFvTtVg2gpUomU
zCuOfOFqAEJxmk9SoGVqoMif17DV5fW7HS65hzbZinEDrQ9J+ouuS3amT4gCj+0N
+pp7viVroxo8q/ICtmH0j2P3hlttzbPkErFrTggccmr+lnUndzVeRe5s3KoFk16F
REh6yiXMyqLk7obDqgSE93dT98nKvqhkH9hRB0VCSlZrLgx8Nl14b1OU7GxX2kyN
180v+munmeL9+RnchC5LsCaQMkVH4Coiv2RakvlVftEkECNdLncsxRilKHY4qJK2
m6TNvkxSPfjmd+cCfQ1Q9uzkF3+qgQoebVBm/OMO3B4OU2adRVz/CyBDH9ZbEY2F
ISCJyxbYHvnJj73he+vQ5uR+6cP/kOJ0O1K5gCuovAUqlPhzGp8KwZjG2OGHO74o
nQ3jPrmJkmFnC7UXWimtu8ydvpZuXjhOs+O9UtSHM8195GW84/m4Ll0I4cjpXD1J
Hh1Og0Yd11bjEMWSJEoweIZ1H7Su2FhBOeqGSlpdfOAhdAvb9RR1lVgoJjEcc2Mm
/08y92b9wueach6CRWZhIi+vXm2o+iCLA0JkCRp4+q9M6YbdDkhRc+R+arET3K7s
9WsO0ZPLrmKTzK/kuRhL8BLX6K9vkENsPQlqzQHFQ6iCNKy8WnYOX74Nsg9PoHM9
GQQmPZSOS2gvfVCIU/MdvN3E76sIr5cEkj44q2t4Uxnw08/9L4d0wEyGnnj+Yf0J
lpcWwonvNiITECjFOFuXna2kSl76iWecCOdOMt38PubP+wzQDguWbqj8PpLmMLOy
GiwBsCPMZI1K1TF0Nz/50xS92sbGJLdT3034hYsCJWjka4fphPI9fM0tS5UQlhsu
Bhg+tCC/VPj4RJcMEjgErQN+w+r+iRZC96Ewz+RdGKFPZY1pSMRSQ/hLtjysb4tw
ofvRA/5PWqrTQUWKnsT204BhCuC+Owf06TVjG7Gdf+6DclcNISg3s2SwjvearjfJ
SdB3dxrF2JmHNjcoip+TaNDh37wVznv/fJ6PpGkSKL9iu4Xj1eWc+Bk+Rlf4AZzt
CxgPGypiKsWxFoh+tHc6NcSkOBA0cCMTOJ6EjBYJ6FbAEdiPaScgEVvnNWZhrUXS
Bak3dvUTou/KwcDpvzO+M4qcDKB/o6WpWx/RexfJYzM5ohcLKpf68yYQ3Ya7Aabl
alqTJj05T4xauaB2oI0t2/jLjUjUsQmdrmImcD9zDoRoBx5q+SrTr6d3D8iFUyiu
MQVRR6bGJnnX61wX+DiFv2w2hyBBu4MInTG4Juh37iKyPC/ypohJIwC3YjuaOpK8
bFT7J7rO8l3ZFV4PWRVKIrV4hLuBEruwwvWYglf/NkrRs/7R6mwv7FF8rN4rDPLA
iTNZKbEEbOd9ghgSVBJDIh3KAzz7mGd9FeBwzVgbpGJHdqddtO1XTCiaCJKGqerT
HDR7oX+nTaiSQwcTOdq7pgbzvZo2wPsIOjwyQ54o4H33b2smK9eI8hscn+WHz46/
QLw/B8YYF9vOhY5qQFpp9ve73Fusp4u0Dom+rbvhFqStPw+Zjh3uaUlQ6BcyHbKm
yAjVs8hT4jV/ddLX3X7S0nf4r2cva6vav/yoWGTf4bsSu9S/7T5DokBrzE49EorA
ErYvku2lYxpQyAIk2F8EOWbRLkiB0x+wPIeY0JdLFnPJZgTzj0zhbmFUpISyk0zd
10yQsNFS+MV/4N1ZcfbK0sELeBZU6HEysjFySn8nDieJ/nZueCd19ZZoX4F2hTd6
04nboQ6bjFSG4cx0pvkesOCb9A0eFySoYPLZxVSi6E+Y6PfGkYCfRUWAWPZMHVPI
ry8Oyy26lxfRlCqalVDBZ9cv4+SQXrN+0yCu9TREue9RtEbJV8ZlMuDY121kPQdH
tFLGFH5PyZHh8/wbQZH9fe3nZZBCjF8aY2CHmJgA6NZNJgX9qwp5Jmqa9IlQkRJY
qOgv6iiGC/ScciXr3wNv/akIAD2yGTr43N7vhpAE46kw5qF0ofq+wiY1B6b7GADU
hD0ZdnTtjSmVyAcqGzc88RJsfrXkkYCswlkLQJQRby6d5DVrurBk4uS7mgRXQ1gI
NyqjF9JrWvTH4E+7VUU9nPLMSF4M0lHZUaxRSEcAc/mNWsvv5jMwiwSloOE97cRg
rZUr4DycH+xswMx2RvYvsN/TfyYYTdiGrzDW8pQJSGKBI4DFKGv/IvFPCxxSehY/
fYMmp22uN1mKMw2J4CbnWN+cXRMFe1i3HIEaQzPOr/ziJuentwQmwYgViOtd9lFE
f4ozGB3IquKofcsMCy/MRoMwRPO3+bPqgE0wLU3nTehx9BteSNFfxnKuwht1binJ
eDnWAtibW4hpdN1+8osJFpRuQBxiuDYtoVQBkbM077FqGOfomgbQUwDW4BzWiVZZ
9NhVNMnR1g46YhiXhSC+BDqLjWKh7plO/g9aTf5PnyI1byiNGMT+ftCq5fqzncx4
hRXs+4a0HSrvy0Pxh1HLiXA35Tcg+bPxbTqrxI72vY4CgIhSmBH2Jh5eQmhVSSE4
UWRJvAFaQY3KL22mnpc8RMFRXiRNaV6ZCqsm8re3+rvTc6rn/0X1E6RKwdf8QtJO
d5XyOrxkVUXpmlyaHzXIlsSqcL2CYjLXXb7veS/vXrFjM9Y9AUJk2Z7hjF7zLs+v
Oyi6Qm2ohq8hHL+77snopHZL7P5/Zc4f0eFcojM4Wlw9ogw3h4zS9lufof98andH
9X8k6Hk6Wg/lnpdYKvhb+SSKkMxWOCk5S+YPOq6t6bhcd2IyTrB7oWRtNsDLAG62
jWpJXJNv82nJLAYgwyLIjllxNv0H6d67/V5oLqyMOvPJNLTWTP2l93+GWp0GgJfA
NrsiB0ah7cuELUaqQFwrN2q83W0wEL08KhTysfYwTjZ1jx/CfJzLNEQi0I4tjgUY
Cd9obXYJp5lWgocsDAJRtA47E32VRNtbA8sV0ouSS3Y7NByOgDRsvoIV/5pGs2TL
r9iNS5FGqWwXennKuIAkZ8RIMqCQm9AhdAwvLYZ85Dax0dX5Dfqrj4U2LgpQVfII
qqZnG6GBtsTdV9auujrUKdOkEZhgs9kZP4FVs+zDlEiFbjVfiH6x6qDgBZ43rdi7
2QdciJfc4VaVF9/V6UFSnywiyWDRAKitt+uZLUgi5/BX4Y3zsx3x+oMXwwTkeqsk
+ILnH9h6RVq+UK4P8st54XZ3jAx+ENGsXmzi2HYsLAbpOj8i1GtivHb2xJSX8Gzf
YpcEnhuspL7fAEn9XtWa3XI3WIwCSzvmcZof9O8Kg8FlO3X4+dQCOPjugbIv11iD
xIHTwOOiJHfd+F9Aau8L+BwN8ButsndLY6gr/9zsEmV740swg8taUMlmBFS/uon8
NWhdt/ZbKTXlMV3MpDLYiGj8a06q2JhvCsa+rK0q+g48T8+DCYfm2VEibfGgZz6U
+k3jgj2pUFvCR/AfTGbb9QjKArWI7/0Bk8tS7AeDcmkU0Gj94iOqHZOMwxFrrpvq
f8n4ml0FyxP3WXpT1uNzOs/Klg+Q8KwDtVswEQOfQ+A+IO6ZAPgpPNqQHnsMglEF
Abf1tSDluNzRgaRzAODpl19Llf+xrM4Hn6Ye8IBjLhswhaPT3lreItfpLPR74/Bj
hfYwBiiOs+gh5qhsFMDDLK11ITGOTDJB8ev4wP1JicYoXi4QynwspWoqQjssxIfm
Jmndi49VCGhELxtQfIHW3jQrQmhOgzuFcUanXSQxoKxAVzX2cF2suoEFLcaz/9r2
PZ1V8sj6YeklAB7wjWkgic8/Cx0c08b71wfmh/5o+P7Ywed3q9ZbS4ZXOhVRtzQb
UNWHypLAgLTJ6vaPt3W+Chz/gWHxvFg9zckck7uqtjFDAPHGXWlHMLTAhxCt6PHO
lNQd03S0kxyGfRVWGvq46Ocpc00f6GDVaI9XSnxQkFgspSMi+B06w0V0sMP/kbYM
enU/D0xCT2bgci2adV5SAGs06nQTlIUM1g9ov8dYJKEwUsZ0eK5tkuLc7YfdhzDO
46vKh8x0vPmdcOD71tkrIeXzFEPgMWzKYJYmGo4STRra11G0Q8bZCWXJv55ep8bg
zI5nKPFXy2fQ7jcxD41vmzEXhLz7WjeLI5KQkAN3XxUjTNHOtpetgf+ErD3g591m
msCm3sFW0w3zCSxKdk9w6+JmLmoTFQFoasRuLHKzhMNcjxdl2+/wq+JSfraKgXRS
659oBKiCvHvpHTMQ2go18s6A3nzuu3oaq/V66sbanmY03uZCI3CknKdv9R5SWEJU
v/F7mwLwDVYdeEoLkKsI2w5HrbGAEqnE8AnOfONEUPk8+znfuhVU6joWYe9GbuZT
IDrYfSGcHtjd9F9w4xr3lqt2toOjdvavFIzku2Pz065vkULIs2iJJjf1z2k4twh0
kd/3XN/tHVaIw9yOjRUqk8MIKMMIOPKeU3pNN/XdO0kCF5sgQXJkUHw+XDDd2kwU
jcj4ulKHZiF8cJmYeSu+3iktHYl+YeTMDxUQz40e2/lrwZDRoPpCA49eu3AAXPi/
4vWFPVynS14mCmrqWRO9hGoedncBGdeG/8wLt0L37vqjU7vPU1o1EwOw1O161JV8
/H4eOFDKJjBMXy/EPw33gBGM03IsmOKXQBhw1i1onQs/5PjiS80qt/aSXEI7Mppp
K8ReZyqwkCzpiuVHC2qL6t6cMVeub1xefHv638zTQaJGd3l3/G6rbgKZXjfsmU7Z
HwAokJxCattq/0vUget4gI/4ZgIRiDexQ0gcadcz/se7QMME5iZ7VGYeclIh0+T8
GbbcPPOF8gDSVmkJnAeKhjn/Qf3+W1NXbcQ7eOC7GdDletHAYNjVd/DjiSQ5Bj20
+NJkU8oqUNpxUAtu+51EKM6zsx9q2ZUazASqm/oXxS0wFSz7PrG8QQsG1m3mBQWs
Zjq4EzxLvyKATgnF0N+g0VNALX5F2Lw0QahcLDwRgA27nz7cRuo1roUMDdpmAYPs
ECeQfxEie2rCqT9uLZwxGnbBOa01FxLPw0/s7htTZiblTgxCxAnBhfzth/p24WkC
LjgTnmpqEa+bRnJcs+Ezaxs18Dfv75QkspulDoPtmh+aBpDsMae8CqrDiC22CT0q
ZVbU5SE0Jr1JDsdzKdDOiXflLF7D5BKVdxhWnFBPDUo3ET8k+knRTxwbFrR6V/xN
XFbBWOodG/fY6Nev+5KR7WEVhBYTjg/4Aol/DPcHnP8/tTYvrxfiB58CuQMmEOuj
BK2n1RrnCrC7E/lGFHR0m0eQGq6Ja9doIyz62JYIGyYLQ0xcM2d0O28qgErnKSV8
GCuRCgt2qx/wh+SD1FC22KF0jijxkylfQk80Dh4XY7B2kuC+rG8NzUBv4Eza5cN8
kVS3mI9mla9VFeZ1b3AR3mEY4QxnSii8lFFJZhvaD/phz+0hziJmIyfBhrsFLN0I
j6lcveqeJgPtYLreb09snn5V2e/ouoc1DEtohStltDtNpJMn89411kuxmRmutCX7
nB4Bqu/n6hT7El1kbKe8Z3oc2vrylG/BrV28uFS8xL+KwwFcT8iZ3sP9HJXo/HyY
MxfjAkptq+SuLHq/i0hVRHD0peX1SEG8DzTnHAeHNhxrQbOjcVUDRrQvc1OfVL1h
9rQteSV4Z4LAfb0M+FIkiraFwftt1eIhZEgcmiYvWfnzh80XSe6eH1T9YXpjHqdB
xtQcWePDizUoS5ZbQ218JF9vRZhCdQWux7NWzfFJqRqzmJcgOdZ0wP7aV0ErbcMr
yW8nrEm+mK4vcZSFmcCU6xdGSzt98CAhCyRXB2K2U+129JpydUDPNZF2eRIss81x
od/5/bTuXE6aI4jg2d/XpxoxoxhSunJtIQSaWHgOL+M9ShRlsufLjPAp89ob5AcD
h7y8uwhSm5sXy9GgnJuEUEBmA5kTc2UcEvOsUj3vvR09ksj+eS/pT4z2FRz4Ub8O
vmCIfLbaSZ9r3g67NmIyGfzUFO3+z3+Y0QP5eqmv8AXhn438JqENiFywiIPQJuqL
E/0MhWfz87s6rjKSU4H6u1EQfRlTiw1+OuyOJBlI406MOVNeiT5pxCEWAS+dXg+Z
S9T7n9GvUmWn2HH/+k1OPh288owu7pVZ6wbFzpGorznPatCtSiiMchVWQ7IQT/PI
Uh1+HdQU50JR521zIPoIZBcShm+7MBsdWGpww/hFDH5qV0p+ovpEADzyxcycC3Sr
Ymr6uiwxefaizCnJG8meDo0P5DJ1Q6PicmMGjwNdMyy7Cf3SN7PDuqdfNIYB8cWA
TB1uX6ejQKssfl3z9QObZSvFmZ+iH1t0rQzWfDITaHW/WxBzJj9qCep1w4XXTKII
703R4GAsKtRofX9/P++KPbKAzy1Q5rO5HvtfpZzgHj6/wx/FQ4zl84s+e+ZHo7eW
IK6Cj8elXb7r0AOb3SGFQsbQzmByXhyDEuktgS9qmZv2Hqz5oO0BC1rYRhMUIGbH
Wo9TYlRtWsQws2pCixyGvE3d4IUvLCf8TAI/QIHY6EW3/dG8lCjhBP8T7uURr1YO
o3Lug04bK326m2LQ7XWFkvTsNoeIs2y4hLyHi0tusWY8sX4t/bA70W+ve7XSLHJ4
IYDq3ZbCk2lqeWhPTY490tWR1rrI0jiWJV2lnEcG3G0eBwFgjoAkfv8LhnkPLOLJ
RIjtato6PEufeTJ92ebdIqU4h2nCT+nCmCKJPIo7Zw0geFEEqjnoeOJQWoWYkQct
GQzO6U8SySDn2HyPmMQFns0JeQM4+BRbVa5GF0ntuXgAxvC/bUudPRJ6czdORWzq
8UEFeCmlpvRh2LR53UjFMyLrBvl0liBTZOOse4vIsPNtLFbYlVu2nTrXJTk9zHD9
wZLXKNYq1r3xBI+LDRj476qX2FF9nHhBRxEc1N1aIXWL9TnkdCyOoPGlIcpzQo3y
03oX5WsDV6NX+COMLYhRzrDAkZnuF/7ZpCwB1REiT0aIEc1mXcY28OiFTVgFvXTK
isxz6mkECsqAOTuxW+UmUC1Z+XwvdVN1YR4RHW3iTo1CFtqv4/99uJU3mqIDBX3y
lXhXIK/+PbqBJmkCTgL6TqZKP8ZFdO/5nL2LL0b1qLV2kZLjeb1YaFdPrm3I6GWC
BzQ4tg9/aIKDErHBI1NGe4Oo/dw6L1mQVoOZRQa2Vg7N7hL/aZXN3vOf3dLvdtkv
k9JAgHrnLVeqXqL2Yn8gtleIMZIMiFQTsFjddJKnibQXyB/1dobhRYCW+JVwTvKN
GEQXVKayr7UxLOFMSTjlIaTYLoB2aaNdzgjlmG+NddT3udDvgL2TijTd2ImaPV9U
U5bMF+7y6Lzla9eVt+KL+y1L163SQYh7lV5vTPmKNWrHxNT9E4pXe2ZoruZalonw
e6zj8RKyTLWdgVCoD7ErxsX93NCHApPcsL4PUicQIKt0nvAmkT4NSi3sLXSJTMzq
eQrsN3AWVXyrHLqCRpYP1Dt7XqJkNZn58ICojR9wkaoAMPhL2LIRIMtUH/Erstx7
EZdf8ce2Mvm5SPYfyPL5pMZBmJzNs+XceEwAK+0WjWXnXuu81+OtJQN/BQ+BFjJK
CJpU3G2hetRPqQLLCIAyq5ROPB0NCtcmI/PVZ/G8HgpvyrVII//zGSsPw4hdKAzW
jP5vc/26ffKLD/CQPIFl58ZV6PUJ+IycfR3XUOsI/G1Xkt0xnid5zJ6Rcms5bNBo
jjBbNmQjcmTJwbSoWwuMxBvPzNPNGPGMHnIYmSD01zkERgVETNemcc5q8zxO1ZsQ
j0WpFo0WX+AB6ivLffjlu8a/gD0BrEgUGRDZSZPL1qJWR1fHXDKylZekMDzpKVG7
owZ6aXkUPKYXc6CLwpVknAzx+dSvgQHzQwIsfeegAKHsox6gRyIGNswvlkAn9JXf
nO1z6mRC5ioOKSpai/YO4imgMqZX1DF08CDrYJMVy0H8hQXqzWq4dPcDnrO5hG+i
86vP1dPg6OGZy1/6YFSiieoN/O7rvqt+rZGC4jAB0rbTnpdDryn5tKdlKpuRN23d
MxxubMPJ9ABJpVsKxbczBF1GsSmvDPTVvXPVUJLydS3UkOxnlFR4lYiIY9A9UAbs
61uhpfQAJoeFv5GZTVktKbIywqRqbx7B7yXOcfUWyP7Ys26HfiBkzZhMBW/f9Rf9
6LpjRava4EEZvKfK4w597tFssmaHRjqZepLHMrrvvxcDO2lSj5l9kOJA6Gwli7jy
kPgLtnL+LjYPxGmauz1vE9bjVud3hE2NMiYJsK4ZCVMLEYgrcLlECQNydVXD41JQ
FeBo0zfh9kNvsX3wnaDCOFxaUBkBS20gFURQWWUaRb6RWBc8IqIp4ngz5rIP4/T4
Dmjr1/4Uv+jASBrmauOjdv0nOZ5aXdMkB21B4KzRq2Y8iC/B+DHQQv5Ksekj+AJ7
tp9l+q7sV1Mnq18HJ2hx8idDrr9j0d08V1ZXJXUs0raDw8wEGPe/AixCDBtNiHA+
3aI2Ly/abhvILeYjW1F98s/ntAARLKLlevXcCdZeuSC0zv1jnpAj1FzR/osDPJae
0rU7sgf3HqES+UzktoKRpmKo0u/gz28M3kWtb9kbtsgnJa5b3rzJBhNa97Lc3xgu
PinAkBZzM0g60RTrW8qa28EYhG2seZFhglpWTw2YaJ/9Dvdd7JgDlshLuJ1W1kuc
ECyxaRL2zT+/lpxGunBS0cJi4J9vjk4Eed161wRp7kHSCbJETTGYVmW8kCQZwY5C
2IiActhluhcn8clyv17hrzFbajuSp9lB0OpdOeUB0PpDfmTtk5SRyZavwYyP5vm6
wFcWJHeUpZEu2L3vpNKr5GGmMjBqTeDSyrdGqerghs6CBmNUuwNEkS0M3gqum9j7
xB6V/ftz9o5mR5kjYy1GEx2EmINjjDMe/x2yuVtxNmF2x55Kv0Zo0iUXPaJsI9DZ
Qom8fNRuhmbX6xIt04fxOv8jnE2w9TQcmYujHslA0ccmRTdhi459U5llboZVJjRj
KlICJUpOwxaOqNB6ilUtG/Iy0f5v/EKHPTV+WrmuDXbCo2TjDP/rDLP5KiW5GUim
+Dnxvww5Y8hWl7/wViGM9hygHpF3AeEE/pnRf//hcbnYn/1LfOmKSwGYgeN7FwjO
UHNBjEmj5kMUvV+c/YF1ZDy+al0qpsrD6xYku3ha/USV12EeEqJ26hjtmpxLoXK9
EBODcJuFzR0dgGvBYH/axNYQuYN5E+zlWjExeBZ5pFQ1bu0jCZIFIqe5ClCelSw3
8p2bj7op5VQVQNsG3cb6G73GioZOStc/sGpW1tch9QQ49NCgILzRWicRM1n2TQkz
AL7BR3E/L2DkBtXsZcx4a8GUmruFju14oEjiLHFNUMfxRAMUosgUyw0Lws1SeLlp
fpuLkl9OAZF+tKDUTNyILO+SF5CoxJlJ/q80z2KBf1CuHr3mt+wpAsFGlENETPgd
CtrnyYVjH0UlXGpthYM4K5cDoB3evNzuzpppsYpzYtz0ci8sp4ZwZq7dCmoYc1E4
IJfeSKFWPuToVkRTesgBYyHy9yMefsalMp4fLZ+/icsIRI7IxQRXm3aPQnFrOmMr
fIqKSiI0Q7ggh5gr+PdGJzwL4YEfMGCqNb1K7mzb8OJrno2+YKCMbW1DDlqTSNTM
Pyn0AO+mczasrDM87KgSRfUdfbkIb94nmwoPaXXIHaBKKcSv8Dj4zdxqM0A+aBvM
nx/q8nUf9WPV1dx0RIsaRcwND2Qh+MtLCvGtN76xRxptM/6NmXLp3DUho1kV6G2y
GsMoptHi/uRqzumUXbxho4XKRA0SILcVMwQJOXmzq+uoz9qwybE0GaDACMjBzfQP
C8x7O3Rb1tpD2FBE8+u35L5c4oIxswkQmmQlhHqGJElzxDCbgETZBWF/9yGoJphU
rZvrw/Y7LQaP/f6tLBCaxR7CR3MM7Y/Niu/NinjvjZ26nuvG9TjLZ6JULyD2lfUD
TCmHokeYqPoNhgM0IzZMumTIXJA3vGJ/LUA3ymfLl9QTGPJI81hDo37TdTD5KWGX
FWtsIqQTfHnwsP99lqmCRI8qV5KZl3aB5QOEYIoXbkyOsO+58BBOIdHJwyhWXtRp
1LZFUljBYzChzTjDs40trFzRTyVBfhQwcxsueTJCZd6o5JjEZOJsSavIt0/JHtaI
A94BNcfiFg85QS2oMMid7vToeJYqXClP7myJFYst2Y80Y845Tf/uILsN5JvIdOjA
b6J+eaomqO5Dsti5bIpVIgnYCRe6wM2ajt0oFQEAVWDUsyfwYiPZj1GA5WGC3dru
5JefAMCUk52TDmqvYr+BIiW7cX6EvKJTpnHldn0eWVrMRsWafC57sxV5vBzwaptm
Lq2UrClT5kLaaZNlYmrI6JefkKWQly2K+T7eWjNsM9Zgfmzk+DvcSsvZ9bfVp5zu
pKYitnqDc36adtjTstOBOHeebTEIM9fv1eQrvZZltpSO5jm4ccsjgpWw2reMAPQg
kmORQU9AJdp7JgayB3ujMALkZBXoFWYM9E+GK8/uubBbITKRyJpScqHC7xWkGXLN
witt/cop1jf62bkxXlgo+0bQaaV2TsVKznnRyE1uc62wegr0vkjco64H7vDI9zbE
GD4vZv9dW431x4O7vRdz4kHdwpoGu2icc1oIAwadq+qlgWSthek1goxedBTbbU5t
BLsJ9cn3CD8toekV/SgXDBfVpVuNAsv4Lks87BXT4I9BgOzny4Vial02/aHn4xyM
LeUjMqGubKeKRjEl8tgGwzYg3j4ehQfyqhd3UCTmewInrO/Mupys7B8CddrH+IbJ
uBTaiAGfuuji4EkpSOa0a/MQKk/I5gia4G9tgCbh34WudT27/yFsMi0FIS21vp9x
JqP9YrWT+9ORuIaiXwCaXzWRmtxvQiRZdSfZ3V8l+ylPrUS5P+MNDh6TW7oydp1B
DCl9hstyNvm2vtpglmwhiTquxhdqkIt1Il374h5BOaGN0h1uaeOBQaRSlw5p2q0b
T5A+E/nyMiWpcKhl5+4DKjkkN09h+Sc15n86wVsH2z6eG8DjT3C8RJ5EAzGQoEOA
nYrXaMUsIcmZZFIIv6cr0sgcOrH2OGOtfTnk6FRXuQw0T2yplc8kRHJMD/bhIeOr
QishFMBHWaMmf2W+xGHwB05f0vnzS0d+quT12fd5d+btzI85qMI0ySRs/niCAQIL
N0Z0LJwjxDtAbcVxb9eSIdTVi79P3i8GKlLYYxB56Mo2s4gkBG0W7yh3ghsRRPjH
Z7c5pGz5tFd0gu9wWC2mDPLYvt6pVBhbZTnsmQ1v1sqIZ569lEj0bxfxXhi9QZec
0Spq+rcDsID/zYiJc9gO7p4houj5fjDsezN30WDXL7LUH1hRCASj2NqfgZ9XWXEx
43B8Jl1hSOF8jwY/VZcwEIlcj5q6LSoD7aQuqGaBdkuPsmTQNblpIBniFc0u8tyw
N4rOpf6HFxpNvTgF90izfuSsUAuLuEEK/dosHuVVBrOD7d4IJNfnbPPlIcDlhK+j
jDsaLOgHKNaXrvp4iGRoO/NoElv0u35KlaCLSvDUEo+WvFGgX3JE8WSvdzn4f7Ot
DJl2RrNH7X31kQEhIAvf1+MlFD+ZKECX9T1KHaAHrdrTcSp+CrJ5lhMP+opZIR0w
R0XuPZZZMqky+kPEcshK1CcfoXzj8rsRsPlr0dktMbBsR205c1SC9tare89TUfhk
maovNFxm2Q5foaGHvYHTRbz6R3bUqSt1lOZiOtRj8xZdj4wzeNywa3FvqG4QFKw5
WTrnrd+7zp+uHt7fc/HgzG0xZJLQJdwtX03B2zcgRyPtAaJxoTIRHVBv1MwyuUdc
9Xi+M9WPsAo32zEWOcEsdCiMNOXHkLFPXHJLH5pCNPqibsh7Tfv7w/KwMKOByvfZ
GOMclHlf/kCZ7rNv+zQNUixQ/if2PusDw/t01+0JsU5VtkWPhu9FpuStbBpNRApP
b+U6w1GNwq5vlZvizQNkWkSw7zgwNYemZOZ7pARMnfmIiM8Z+cax58EsHCvCbxCr
fU26QVqvF3vJGUBrteHijT+7kpxeRzE1k39SqO39P3h+0jU86Ce+haTRb/3SdNI9
9mBtwzCstw6pDr9U9JzsGkQb7dHzCkieDcDGMHHwf2/HOP93DieSuvNp6/PD3jE4
mXO2SXtuCSnMWKRFvlOmccZxTMmSTDoakurYn5HkP33g0MFynr8u+Wxki3dX8rli
EtTF8yNhH0rmE5YW2+3LHzPT18qS87T/Duh1IZ0nLAmalE61wPTrILtCGZj4L6g7
IxaqVgBy0kT3iMQsX3NvLjM35XpszVG1zKsKBITyLR7XdlvqW+6j5ks0Dxn7m7Nb
0hVshREXcIvf9/9OxZAVEAXKb6iYszXKpWJIMn1zhD/9ULQPjILcioP2sT4LIM1Q
QOHM3aQ3BX9MaRtH3wfd684pcuf4S6q94uLX4OONOBSYiabV1IaOfK8AqS2GxxAi
IVY9AlGrwJqI+MLJjIaP2cWTEbwB6+9uV8nL5JIPXEexIWsKVU2yF/yHzUBASImY
ddK8LfjqdhEnOgvyCE0McJtVBji5j7dCMOyzkeOvz2tDlN1StvasG+bsNSzetJbR
sqNeQPp26QZan5kuTIh/5xgRFD9Wx53q0cp5qP0f26FEhONKwDOwPz1paG/IcMhI
GsWaX+tJFzBd9ai46NFCTebWU0L05PPdkduDXqK/4iNa9k5K8UtGbjSHGHTterW7
E1xdgJdAs2gToHSk5ZuzyZzigaTbPbpdT2tLGJPpEwS2x2QhJxwRSS3fwDk5kzm0
CQ26S5OJwF/XVTVNs45jUa/wY8HfqOEmDdpJL2ZpxcMUgbB1wGXdEdx6V0iV+tZR
0Q8mSUjMPGdZUEdGqsVPHsTSjIP4JaBZLdQ7WSg9GS67ygYSgRndt9rGa59BkIh4
Wk8/HOBwS99D8YJj8MuPPUGDiV3yii5MZdt8NqKWE7YNbLaNueddbKQF54b4Ul6q
I8oCe1sc2u5VYSiYA2ux25MhF77iWSJ8HaGYZJLrEEWuo3v074w22nh1FVtnh+PN
8AoHpE2oan79N6TpNrZReV46aWJv3IU7mYuCzI1OR3uNCLCkiz6XVqxGMh14Mre8
T7sarOxaHbvyEMIOq7pL/XQ4zUiIITMRdTheKwK2CXP2e12eG/ACJNkZb0/cezmy
jFDGJ3GMMx8VfjUtfkk40tnTm/hvMi+Wgr4B7mWlYkjUcmNKVp/d550J2jZIT44J
c3TbqL8fGDjlaOHsRnN/UZtH5EyiXScKXhAhelKl7+NDxdzTpfVKAZQttuAKbCTY
8hN3nPh1ZgSn9K131VmT1gk7r6BRoUloTF5l7cpYzJ62+fAtuWJtXkmqJevlx3zz
GQVIe7nHn1P4LZl68CgEjl8SCriwBmiOtpOl+HbwEWRELtvi3HYrZBlANetZS6Yb
i9te3ls6bbZ3BvkZa8RpPcN5lVL3waW6ezdGJBDv888HGO7bECkZ4F4wCGcNeWFb
SmhzEKKBQ0DDe1qBXq/a/zvXCMkIaFWH8LMtHrLBf5j3VVsOBuBpRGHoWQO+peWx
JGcnVyHPyoLyju4anQQ867lP8gCc2L8KoLn9U8I2bEGgENgSlsfE7S+kBWKuqtic
2YigEqoObgIMNv8/rJv898gQy3yE7yFLTk+S+dfPhAVrxcGH4/tZFeLDBd7XQbfu
VcE4LCpoQqC5dALFMMY5H2u8NoFe7d/YaJRoXdZQ6P08gAxXet8T3GukSSxJQ7Y/
UgbXUJUtYJw6zkFPWOgKPvtbGPFYI8xc5kBsvyaMWFK3N3iDlwogdlTkrC8enzRF
7/+Ys+E/WBiyO2sLkFa7dzIwwIQuyLVt9WnP4wjsGiES1FVhFY6/NLM2CWhupfZ0
i1/fIiVpHYx2WUk2BIFiciEstD619ZRmE4YBw34pRaYVm9D3aWojcxFLn2NJQx0z
XCECf2HUMj3/7E1I6hbNS8nqT2RKIs75jRNy8h6q3MZWygZTa/Tbz2QnbuCeunJM
NfMUz5KnsKN22Gjg4ehW2XFXkyksRZS9Q3tRJkZQwggYWQ5sirPvydWcgzeLq5a4
tVTnyqASMokU9Q0z/JoNnph3WME4/3i7GoD+6g0DIUviYYO1znrikv+pTYF8g1LX
Ic5CWlW26ZWuXoe8y9/KUXWKfYbies4qiVDEjMJByQAQk2m6QSMgRCewZwGHYIE4
1ttrR2IkW9NcnGlfQ2s4cEtEa0SJnFIuVOtKwlG8FnnW7A0Nsvz/tTJ6BTKry+2W
HbOyhSiCQfkPw2nlJQPhgZjkIugGa63htSvnt1DIkX/RDQ/hr5w5B3Mg3/x/RqFE
DKkg4MQJ98qHuchDW3dCh/YDaafUziS2elj18lL60izyR6JFKHS284EtwaK65tl4
xMTorriG+581j7EWW9aaHw7RKE+CTEEzsTVTO95roFIhImWLR9sJK6CVnH2wCuRM
bVA/vQ+k3YA6KHBlJ4gV4v8p06XS5uBVYgEdEgJs8m+Q4JtmAWVdLw26bw5duCuA
2HHJ/ZnLC3HNCu61U1zVjzZwo1/wHKHy074CeGOcs3tQvhZZ9NmgXhkitdWMItdt
Bf2mEQR7waawImsi2aMwHnPfClQK2tg0VrYIgpnuXW8Z+pwgB6WDtzAGb0pH6FTQ
JuL9sZ1WfsSBn9h3e62UlsegK25z0ZDDxyPm4hUXuT3xASQlfxhotRLTJHBb790S
3q/1f9cYWd9UqHtpb1LsXaRaAapAv56RA7F/abwGRb385DTK6LyEJNM/RKh1Q9kV
dMKRHaR7uF0s54gMKNaZm2M374Vk8O/BxXVjkugmZ279D4b5qc5QZEaMMlxbMBjo
2yjWB6MkkgeNKD9MtmwfLfdBzoDWHdy99uezTEHZt8iDDtvnkjgp00kUnoQRjY6A
9sIvI/aKl/V4UcRIcIE2akVWoLM2XM9lmqRaJb/WQFcQ2qlqOXk++6lryK0mrFb4
0Qcrt4hCC8Lo31ZYwjAy84cDmK+B+TXoTrRkX7OftXOlk1wz3Tt0lcfDo67N+866
9IH80ZS9vfxzGJe7E/VJ7LFrmgLHZrZrKKYUBwg3gOdAtlz2cWy+Ys7vLgIT2tF+
NOqa/7BEpfw2CBmo2BXjfDdepIPsVN+3dUiDY86EK3A+gfUC3T2sJgUs8ldQU5mY
Qo5yV/l/h0vVWOQttu+W7IPUnm/T2acirbP/7Qf0ReWLv69ONAOEoX/tYCuvd04Q
9sCr8YqkxPZVSCrT2OwiBkC3qfaVm0RxXmJTmFgkF2AJF0BR2qrMt5WdC0AcwNP7
nCyjFVcf2yS2Q2agWDqr6ECuX3FJhbeFH0tdIsudDgYsFMFcfitKfXdVBvOGmwiS
PYwuC8pyUGgoUtfS+Z7YDXdrjMREmLofsaEKwxoFCl6tUezVbNarrjD7xqhl/hNm
rLTCSsi/vEkXP9HN9RMZN6Oks3J4GvyDMCnEoMFEkIkB2pvro1SERcUvAg/YR3MU
N0ftYiF/nQ5QIjQPWYKyubes5/x4XSrfEungiKO2rvwERouzKnUx0c6b/uDyllP7
nLXUyN4jAV2kDko56ll80R/9c8sQGsoAet9WegEC/mkL9acqbktJNo/PRcI1WUMp
MwuJrKAYeWVEzezLV9I8E7AyFH7L4+4VDWyzXEVsUKVRQ3Htv7I29otoaYYLPARj
ct9hCAylWlf2b2qNd0NSeVBB2JXD+K/C94a7XDf9fsxm039gLC4JR/uWlEkRQN5W
6OatDKpck6NjbOqweMTamB5Hm0i93A3HZh9AwaQ9OOVzHpIMSyWGJIphF6f1q0Bm
kL6FcV+PgXhIgdB0Z0c7YNu4Dkb7sh5buuZZuN1lHg0vZDLNvtStL5ZV9kApI1v+
t6bOdJRa26GpJ/Wj0WJgoS/sNxew61e1ScZonmnPdC2/6it/Ri9O3rxIUrRfXrD7
ZdjdYeGjaTlobS6+4Yg2xu75EVq1qSycvmNFFaXSDfyNT4s01odlOTNU3epP8ro8
SzLCkiqzBpXsq0DbCjPbj6ap+arQaI368fs4OgEoM2v3xCVxWqiEvafFs0Vu0o1I
e330qJiapEzqrCIOHoByclAELl5sKBVAjB4mT+KbF+poQ8eA7gTiqcZxPBMlBW15
pjUQGijc7frMKjQ64rsZGvoYJvma8prBZiO/rsYXn6DTdAbslj8DLq+LQLoeDTnZ
Cp45UFLrw+TOmRim6wE5AOzor7AqwwL9WHNw7aEVmba9dnqAjk2dWYfmMuWF9ads
7rdLt/LLHDwP+zg2FOYZTkwq4QZYbA42YHbrEn/OmKkgo+AZQoCqcOBGAZuWhGVe
mPQnmPiDKNTADOdFQMfQNzqggZjURC3iRu5cx/QXz+XuLdepm0GQQpm8+NZTiGZo
N+Gcvl5w/WyCGgrxhue6eZW5TGk+qiDpEPVCv2Nv5bjTpY1By7uB4P+0/8q9Fep+
7rbFPJT0FCaF6xXioJ6x6AtVQ5YdPmrTU+Mm8fEL9Yl4keu6Os48e2PGEC6OVSWa
fkQLeDK4xIKKwoGwp19zamW8W0W9/CL/DAf++3zhS2r4J2jDRpsF/4NyQR49CbGu
kLr1DbB+a5RubEyJL+a90DRlMj3fSeBIYyRFJlygoK4mPyxCZA4eWEmnuFKJLGyk
Ie/iFj49hR1PKUP2dG+MoWTzGOaMFrFworxKaqFzKvNIPJGwakyJtOnzxPmAqF8o
eWeHtYVePFJHVIuseG25axKg4RxELmTxP4M/mBe915ejmxJN/CvldRMgar85/Irk
IERSFyyyZ0+Np3xCoV5C6hdZezu6n3LNXjDnRNVb0hWD9lgkFZGnrWAKh1zl+MTY
qjpvdXfvaydagLdHTqTIxVJ47qYlUwdyWVCAwijBbRR10Sgqsw0yX92bg4lDMhs3
yQ/KxeI0vsTCNXDGOt+9bhcf5vfPqK0V/7dw1XVydfe9a3OEVjwpfTvUzJKowrMj
3UBG28M2TNh/K8KH5ibjKBBeIESOOathJvQpccB2eakLjmhbAonz3wchkVwS9dX0
N/IL2HkfMqqE+cr5khVTKTbZS4euEvU2pp2pOLqkjEq8y6REAT2vC2ZDhZ8rBO2k
k/9Q/BS10VRHiHgQwpOjKPAjRBb6eGoYUNmFAB6hrK6HMFH/T5fiPWnW+0D3dEtj
Vizna1h9vXanxhZh/fswIvpDICS1qxav9iWlgZRgHlVMX5OR5liTplOySCXpGgcM
LH9+DFsB2/lGsB9oJoHYwbziRQTDp86aDA8sBxQ0Z+GxeKbj20yGBgzv2RPife3f
f/pWA5RHz7AhDbuVa7iQX1xWdXqK7UIWurVqMeoim3k6NT4FypjUajH5b4cEnuDZ
wNE1VBLlxEDyz10luxVAW3ciDx3B1m7s8KOb6xR172H6YNw6jf1lyoaYuG5tUgLT
wLjThPYoGwlB9sOI2TryI6sg4pWirAWmj0/h8xFg643npRo+iM47MSdPS6WvP7jT
1k20+1ADrlFGzmdz7nj0GDxp90XexVsmQnYPUJYpkmj0dCNH5mhdLRsyIG2jbEAp
0RUj+wz+0wwtpeidU4bsisUZ60PghK4IypSBaSr0esVX+x+KZ085C8MEfddpR3i0
rgDv7+hOR6Pt9ouVAJti3c4NJnR1uUBc96EbA6ajhFrr6EjgGuFBYLoXf3ChS5WP
3PdeKiAb7+w9Avf9qt2IPYG4LhzBM1DU9NaFr77HQCBFemlJaWJnur705BPc48E5
tEzuaV9VYyJctqXkd7XT6x5uhKWagfcZDXOmGy+YFIlMzcFtjESWqmm8T5FDqqlf
SR2g89hjxro2kRJP+TIj/pdnXTdLmNoWUJJl8IBbX4fr1nuGs5/gVPp+BrCa4PDx
MA56XCcunKOBnTSZ84ED4vGmyiQ0j4SmtHaixVvRrTC6AYcTI0RZ8V5NKpX3ZpVR
Xnf4/0Xj/lSNZOU0vriHlwxtX2q6on02bAvHahHrDLXQVh9Z1je33ytyIcwzduJ8
Q48BFctS055UP2EuCzOA/mI/rC2XVPRYGUlixHxXwZYCRDt8oAiqXpEMc723+Mgn
gCdoYSVw9Ed3WsKuUAu37WdnR++zHF0+em8y8QXa3068XtSc1/R8wJBGjzdtKSIS
cg+h5gGtJRX7LjW1+7HypqGp10lGZKeGMoyIqjHu7umGoYy8NG+xtLACK3T8J+j/
DIokT4aKy1+8QvgYlKLmoUwaG4781abElsUkeebADfISBD1Z52qntpFpqQcMUQJJ
0V57mJCeyxydkXiBqr2EHp6/qSfqHXD4VQxqTGR9Q7uOeInwsQOD+eZgfSb8PsEp
0dHcBC3Klcih5bZ6GF2+rj5CcmkBoFofSKwtGf8jCvJX8qKwV2aiy1+SVZuzcjXK
Zagn9aDARc7kMUdY065yTXkdN4J06qygme/dUb9GZb/u/ewYmhXslu2cfzxTPCLF
UUTD4DYMGoXv+pw+fiTQOJrL9ESIvr51eW3bw+Y367zDVOmL5bh9/u6z377T2BGU
uUvI58ziqaMsG22exxpzx2UWoMqVUTqa1AbWE36X4+xcGgUNlPspzPbtq57B8O3p
XN3585rdMaaw2WRXqKx/8GpfYUdk3WPT6OlUU0sPGJBKP1LC+T/csFzPc6nDCp1e
XiRxQlZHyTMQwpmqSV6GjaJJrIx9tRhV8vnFfzp3xFHER+LKXRaA+UkSlR1WkZqb
PPY6oMNPJ3+mR+nmrsYOhzfwZA+fff6iwrQ80+2Stv3Wl4JhnkLxkfqsnVVuqzKj
0fVRs5ZhAQ4fU0bY7CnVlmZXbTY20vfmsn8aXlk1JvH7FzAkZ+F5/Mu5xZjcMS+9
XqsxQbZWgOfFhkpTZTK6N0jjaoD0Br0OhPiUSlsOgjTNSoH5RUbvhJ41Ib1BT6NG
CEdJxz6q8yNl1uJZMRMElYNNm/b1OYNUonpVkF+s9eMLrCbc7XuoYNTew5R1IVLd
jskg5f+1M0jVTwjKstsumqfc3ARpy3wJfWySvkKT6WExUiIBSZlH2Vo9yhs1E94w
PTce/ktIZoa9WD8gQgZmNMEKTaWAIdTz4C9aXpVAc39u963OPy/ogR5Fct3ZnPLa
AvbvYxNyDfNR27doBuGco6uJXaahoILBkKeZL9tQSp5lQ1U0/aPNTmEexrZiBWx0
j6MkWn6KUGcnfY1v1IpbqDzRO1TryFa7CtnzV2aesjT3wacbD+cQjdOiF6lxu5mu
lHurlCVh/pu1olFws9nISU7OTqk+zAOVteKV15M9MnCTleM1CPTD0vYNbHk5wGYH
7WbwwXaa85OacKWSCkzG3fDPlLUezH7u2sglsMn8554TtwDi58OJeJmvpjmt4Y1X
xFVoK6laI3dvWFNcMqKUPnKVsa8+WRyqPk3jFhhVQDu//Uxg7pvP1+bJvRbJLSMP
E+L3cs3izJY+hPducnSkopRLE6O3/Njuh3RPtDGdhjfZ+eWLaW9nFMtpVVbisY4c
Fotsy8V1XR1Ggz/AJiLXFVdK4uHX+eyAdVCvdwP0iXV2uTK/Zz83sgCqkriSTRSC
TB2DL4bhuC5OnNwmsHVaYhnk0EjfQKrXl4ZVI6Hat8bu66gBljv3TbwFNF6nE2fY
gffc4peNDqEdIiYpPaG8Ca50DgTZz1bCrtoq/ahYwzJObcmNr0mUFBa8Jlw/x8dq
GSRg2dugnWTv0XYZ99whZZGhx72RUXwu0V1odyPVb89qIqWoWNBDvkwjmJKdCKqR
Fz3XfUj7PBhyBxP5FBM3ITZuxCj02Ae5eEQyGOv8OeKIlVNT6CqU5aU7WgNWHFZc
efF6ZqeLytEuhAz9sMhPxle+L4NOcVw5O03cyWreV+h4Ve4KjP6LQix7AzrIs8VA
yFY8A0/YbuChl5kqofQ4cwKMhZybX2xCvuHmo8hziumXBoM2/e19XUp97J8V1+bN
uKMkfQYGNsV8YlPOl2I5kdc25EjIWTOqndyUkqVHUZrEVk/LBSghemNpd4nuW6/e
3wX/vnEfl6pBd2P1YZ+l7ZGt9S85AUgYU3D9WV+wpD+Fe8jX2+mxOYNro7132gGa
u/K2I64pRR9csQJQ+GvjyMH7wEr/6dNF8Y9MyeBJO4r9nijLuY3lKX+2aGV+S3u/
KCwzoKGc3dGwGNHNrLhxA6jycKQuzEDucWqa0F3D0cXVHmaiuS1PceQlipR34HAO
2ajMtc5okEvvPHdtDQDMGjIAfaMd/evQfcs4r97mAz2waudyVyRAKCMY0dsDFHb/
4dKNJ5a2wA/Yo3mMJ/uk54J/iiZVJ8wm/92m2PM9enFulmUjx+LBgQFtDWIWingC
3kkg7MbFJcTBv4eVvgPAp5KwifKF0IHiAsYiKkqm0Fou/Fq640+4pEQ3m0bC8Zwc
HGrBAPlTfPTlfbaGKVDOU3QyYUDSymlh7hX15rjNT0S9YVbf2N2QpScgAp2nvph8
uAYf78kB4aH//aZYqTBI0ZXsjzKKmKSovAyL75nuoacbCZQmcBeuBuJkcjwrL3bm
ifxImnh0BE6MkMWfXjj7oUdx/6niC5BdPTV9nfGd04hvNyKBXamxhx1MPKGcsHL/
mIchhTVsuSPuA+XbGEArgDLu9TmTfB+VA/4+styb4Z35nPXn4Sa2V7Xdr+QoUFv8
8Mzlewye6SBdEM/NVJ6xnF0YdxwjBsMOvoESDHAmVE5qfP4+y5rjDUOYXSiCeUD0
5SMhOLGLTbU+WhrL31K+ORYX0ICSTGMtnuyYbHq50KpuVMBqCWMTWh6uMTsGqTIE
9OHsA9NPrwWaztS16SMIH8rBzuWxHZSBeto4c/bmJDMBddSY1OEvWQGtiC0eOFLv
8ntMQnfiIpGP1B+KCPpbzEKZeQnUGcfUKPNJHyQ/l+O/2WRU9fxesEELN2ZTCDug
f3R+rrbMibIDJHl+xhar0on1K0Pk3G5knYBuDquaBbBYoNn7u0cbR0asmTnzsDGa
qbsQM/6/9jFeAV6ohvQeqnpFtP8U7E55ZYgumsjlfXZuui/0DxIiB9P1KClwLTnH
KVKvxpUHBvjIqMh/4nP8d0Veg9MMgB8q9mcetd/laOKcBkzLxzFzLjLafDjYwotC
kOeP4BmTPe7ql36vL4p5NzTMrnxBFsdA1aLl3Wome2gQyJydQikiQf0Tkt6xKd+j
1eo3tpasJSvSLRXaM45SMFGlnruc/aFbzJguhuR+PzZYzftB9bjdrtN67rqYVnFR
sGm/TULqy9PRdseLfKZRdnzh+9EJk0vxaL4B1qN9/JgsnfmzQmjU4iJOG+m9YGDU
B9h4MKV6Cbd5fOVFQ6SiHdsv1KWGpMjtJ0yWuJ5LArw0GLWeR5tGhd24R6cXG7g2
dttdZ9cVnYLgn1cLKCt8LLgj9eygR4iPpAdyOTAudfh0XH843ROYeF1ZqXB0YTXF
7ndU+Gc0RdG5R71vQUVAI6HmjyvYJN6+BKoO9Ffk5sAeHyhwDJjGliC7LqYq2i08
tZvcGQMffdLhRNqWQIKygzWhAMtLJdb5YOH2ESVA+GlbkHuzymcuiqXQvrKtObBS
sfvdmprqerFf8a0ckZFS4AnWdkLkuxTNzn1pwEnYNNTWCZ51sJkKLkZsNtkOYhLt
aFabF/Yfpl/GtFYz4rXJ3Eolza3mfesfMXST+MDdszGk3qMwxv/T20ogXqNoCwGI
+Tue9Km7qg2P+hqsi6VFadqM+MIoH42Y7enfVdMxPwBfQNrIIfsnt+PP16qYsjt/
WFpLm+iG0pnZXOqjlnbuKBQj7sfyKgjUfDyejVxre8RE4GCMeZE0Fvgj5gy4KftY
SkEJFWgGUIx7V5RrZg9/EuGZPngswYojbtaEw9cZEOeRDuLz8Woc3w5e6NvTSSZV
frwrRCzgySEponuIko76zBhEmS+qKzqJeNH2HOkgIJrle62i76L4D0bTD5tFWD60
phnH7Vn1TJZ2LhEGfztLJzY6CE8RoeYl64BBP5nUgRvBTfORyHDTI9TnCXUjLLAc
ptPTjF5hJJcJu4x4CMlQr8xA9LExieDFmnACWrL4purWfdhybmw2QOfsyDNs0AMA
ZYlSTxyEtYtn7ne5g/MjdswUCFGpXfIhpwcKrrARBRPrkLUpX5g0unB6HWqvmce+
j45F7RsExnTs8qyviLyUuUIQVVeZlCfOJ3xRqA1tMVt8XOjOyaDJ/31UqRyX0tdJ
276M6wjUPcXPdZOX6ci9L6Bjo7jlsHwvmlwjk8eDD9jNgFdCHnkGcw4Z40Ktbw1J
r/cxX5mYOB9i0XOXaviWgYgj7vAA7nxXOPn/fMIgibhYye3tPgVeD3fMqivGjJ/8
PpE7KTkpye7TCB2jqrxd0lu2vs15Ofyi0xsqLLypwnJ7ffDRNxb10u0mEpSecgR4
zhHzOr3CHmKk9uCxAu+kh8ZFXlzmiJQ0k9AZE7aRX5zXBYKU9xh5tFgkroOCKAYo
QXAGGbB8co2LU4I1JxSjiEdFLMoIeuf7dPicyqgvTEm79THCz+VZZYjhtNaUuiUQ
2TVxVIBY4Myhz2H9wVyQP/cKAzjmToEwi7rP2H1A4bEuw8pwKUKf5WzBJ8PM/Ppm
0MfuLgx5Uvx4BGCdEzv2POouNF2tBT5ArDrYZl0UkOVGzASEHwGkDroLUMByjh+O
xzrtZriMQdzIJeCxfl+FgXeOm2zHRKI0J9XJZOb7J0+/8GbM4mDfUJ3vBzpOuZ1x
p1Ld9I+/6/AK2sC7c2+pdrfHsr1dTQNIeeqF3qzyakL1aRCaX1Jp0c5ADVoUiQbS
QeaHj1gc/AS0dJk64/uGoY8Wkot1eGOA9G0mQTBnOZRLuhB1vO5c9fGNQYAMqyOS
bKDiPcCLG7jiga/tsp8cIJemf4tUQJsVeIeXXyi/KZ8iUZbu3VOMoC2QPJtRKZXW
4dvsronE2xeAISbIeEzR4tmhw9TX1YH9TWMwAC2l1dLJw2/M6r2HM7lX7Gi0WfXw
IOMiS4GWI0SzT1A6iFhmeYeGgjbK0c/T3dUwSB/mAWhb5Yf/m5+7T5Hm28vFHwAO
X1y6yoJ5VfS13HJ2qs47l9Dde9ds7GBsAubnmlz0OsOWwGzTohkM7YPC4k0jxs3U
XgfEMaKqwVUwvnGH2R3A4BcxyTUe96+wKgbu5uj0X7mbxOrDtPA3natmyh6z9ANJ
X/eeUR78WaGgTyGqqtczVxfI7TaFWzbunSmehCClbUcxE/mNoWGKmcc1uFRydE6p
pufFNDjNBkTpqvfhLkja5Kq4pCoBOHs/Rjds+LNZKmHfdNmyaWykx86MM6L8sxnY
ZkvuiiyGEDBfA+Gz0oOccok+yxv5mD/f4MbqitmdWLQzF4g5Px9/XXz9XX7cuqBL
s/BakeLruaF5ZXb+wwhIRiKOb6wK9VqW90USUOyny/OH5WJgOufSftzxqO7vp+0P
7EQYtsRjZ913avgSRADZVYVvU5kfzPz5awiaqdVL+PIFByxnKixi5GAEO4vpNkZT
zTE9K3zc1WXFBxzHlNLgGCcwEdmXNuVPBO12XCjMvd/PlXBfxgayXIORPLp5k14Q
mugT6l0Eb1l7bXB255i/kQdCGIlUARdxAw4xfXFZSyVeJgwy2+8VCRH2bMTPWMHJ
5isUV6MwUke02KJut4hYwmsXWfKtQ6eWXDCpu/e6yentbODgS2gPk3/PqJ54dY/V
w3y0Ry0BCV5HEl/gnjHzpISqeVMRpajRrXbJrj+Xwn4qPK0/jwJfUgjQV1q5H9Rc
dczonTkYZHoX4iJ1ON9IcJ5AlXYuUChrmBJgL0kjbmVpS5nexhdAj+dVCOXGyQ9k
IIiRFwKX0U5uRI+YM43psMHrLBOCx4dL7m+a9FZ1tDKbV7xZd+lSiPskJHATtZvl
HsegXHK1Hpn2iAs0a0REdVSmzZwv7TmyasLCkTYpK71sDVv/zirpLRLHGKGEn0F8
fGMykLSY0kUN3E45xG6SWfcZT69pfyZZ/h2Df6rm3qO2RLQS+sPPKeVv6YNP51zJ
z8O6BbilimIDmNO6Q8gMQRXOCcpv63mcPiZZ9SvM1TRDrIlHPKbBIYIF5eniHlK4
3SWQAv1S/q7z0eTHWdDn3H+PMaym+ytGnbu8GXThYMhPh6xRrTlWgUuN8YAxZ6xx
SZfI/YBMzKX//S5hN7sr10RB9twgk8OwBJ/dx4mPAxeA6P6PtRL5SOq+s8CkhiR+
LzGdOamLB6LjllxLmSgsLd6l2Yznpj7Y7kcws2UbRNNTSIvzX8NxucK7nxBeCOLT
RaOvqLjIyU0VIXKXXinJw3SnP6z5WZ6m/j4gupsKo7KUz00czxneQvCQ1w5gtWBV
idk27hFoTp5MkDvFw2G1labteTRlaHBKPMOLgp0vNP00lFj1SUF1rGpjD7/OH4o2
vD/e+t6SEkDmF5FT9BM8zxxjYZPE5mpjMhtgdNciiy+Wn8yKrn4j1xPQYr8npUSu
eGYYHOuDEBFwEiL7+fHzxtYgIG/lFt/3VgecIukMW2jLbRnDqANjy17Lw1leI3ko
qNRKcSzXrcR7sAROnSJcoQyZyFnL7lk8XuIBvlyz4n2EC2gtEXaaseLAuUtsDn7z
PgS3rosfMp+A3ytf7jchSx76DCxjjsxM4CV1mQFPUBLuvj1rL1OyGjSLCml2FiK8
WstiaDHV3pQl9vVvlHEVKxVOlXe7g74vdZ5bNK4ZURxpf3IQVAhI16nn1gCPeXQr
/S7ij7Q1zVcXQ9koAOMDEyTyBaS+0CfBk2KW9Y1JihY0rYn03qga+LV/gq+FrFKS
qluC6crsR8DTgebsYCDUKP1QSPvPQolRMBBt1MxpabD2a9FRUgpTWxaui7dszcaI
xiSRueQniPbDeIDTjR5lvZyjvnb3hE29s/I+ygxIF1AOuOEpEG+ZodPFRLv32R4Z
6cUqjrZTEdiOaal7ZLP4cZA7zzvieFuN3O0HPIgpOqFksGGr0FKeAxyJeBHxH+3A
LVHou/DsPdQY5FVeZudxpgee6YiDu32JsyIqgWP/krG2kr4MZfLnUXJAQB1jxFTQ
cVj0IVGuJWE7YH/+s1LCI4zTUTOLj8v30LQKEd5etpV/o4brLb74CMe/zxa0nCdu
9sfNJrmW7WF/W4IDGs+VNpM8kPy06NnueCF6l+bWcxVcEZdrQF3vwKQVNYvsGBcO
WKO2jQwaA7zMcMwjsb9o4UvL/gpPDFlRabntZy6Z4NyHOksovd4LNVKf9WhoN1WN
OqFwb2yPSHQ6Ltez7vHdKiMY7pI0w1e21hzzTfGiSHAG9w/zlxf5Qp3cw5AMoAj0
6cWT9x+YKKAP+D5SS5ql5wf7evPWWY2yO95Kff7pv0Eb3v+TDSn1OBsOHXe66+tg
aOGm+mulYmrAygD8bt+OPYRWQRwiiI0RAwI9oNHL0NEXJpnJh7JnpZUhGUHDvP3E
2+OFtDsVZUyE4j0cI8iUpBCANY4SdykcqWs1ubM7aGJTTlet1szC9TUMFL90cSF9
gFXLT+Gr/zcNVcBPFw6XFg6ygcJXvorem697Z3So34qeAxnV+t40Y0cz/hzSWrlj
2FQyl1NLt6Bx1uilTJnMrzVEgBinZw8A4brIBSHWpB3qNENBMdzY1TG4bBp5ZhiP
eVKbjeVrw3j/YbZ2ggcU1B7tZT/LgPn/ljwvRVB4B0QEDO3CJijUjQiJqHCT1Yek
x33EoWPuMab4+ZS9jmKzmosvKrGPFWfinsocps+c7hwBeZGLMdrt1idedc7b/Umh
Zne8UBCkItrKr8dfoAL6YIgI7ce1AKkevX7A/QhjjcranG5K4KKjg5+PqPuBbfr8
3poZPR0/y+5686+KhBe3NCnT+LroNN1uVMXXWBxjFQtbDNNPG8DoIlwbWcRU+bsi
FxKywXdJyW6vb8DG+cbH9AlEsA3U/+GpqK6v+TMBlFc+rgQq/5+A3xaloXocnHEZ
qaJknziHctrXbl0ppkexAqrKWSuGQbAsFEh2FAIP4BqjuCkoFpCqEamjy7EmRDCt
xgyIjWfthlynFST1tiw7cWOGIIAH2Hg5poxb1Lm8kUWOzzB944WNo4f872WQoxfE
iblXIVHYU8rlUgFIwtTZ7qhjbAZYbvyjDVuDdLDQR6TJEcLGb/rnTLGKGxUCjPEo
0SWIbwB6krmWBNM5vlilvy3g5+honUUvMXh6ieEE7Oq3cOofYhek9AKlF/6OSEgb
p5b64e2pOAA0S4+Q8137hM0pl0Hx/71c5Hf48ZCKX5CqU2qu3W4JcdsdQ869o/dv
pqvMdSZVmUd36rHsgO6Up3c5yK2U+VIBXaWlUxqb7BHUHxdOzkCjnUOBp9ZTteXF
RLnK3lONse5Xw2epb/OPxWdIEj6KbHk3KwNnmVqWXvMZjGFdyNWt4M9dRHCo+5/9
f5obHwcdQ1SaISyoN3ZFP132qTqbQ9kRFaeYlCQz1q1Hsi7Na82FnR+kdvJE00u9
s6/0Xa5fPYHFoGlP1NaDOyrkrIn7k3UuV0YBxNaaMnxeO+5TjRsOQiUgOb7VpGWt
MXiguMcMBReJP6JgKDczLwdJy5eCfAuap2x5qDHUq1PzJ+uugI54bJnKBfL/fnRU
GjWDPLadyqj7SBGrn9ZMbQUViAc6voogL3Ra162eYRQEl21ots8BahTVsfhbCkEw
uM2QQnNMGJAYAE1wYrcOHCLOohLpJMZhVC5yqf0pLuifjTL2F84FHK1jKLlINSJS
ig/wm54+SHZYFAfOLzSdouNFDSBUgZVKWWrR7MMbo2DXDhXsvmGA2fbRLtpkhSsY
/GMijG1awKkrncOQJJ5GYjmusLn3famzcpvacZ/2teHIr/XjIHgh8IcZTPWe3SdA
A1TFqQ0T+MzskrU0RNEu3g+UysVYmXhgRUbtXdkiH3G6Z0oEOZKN4FEKqDvlM5fA
eunbi2pPeDchFszqqsGwfCo1ayvpIgRRNZLY7LfxAk298HQLH+g36NhWE6EoQM4u
uLWjlGwJpepmyEI9SwDj2Oer7TtcUeZ+BcmpDjquvDcLRd+Vn4NBV0DHxpRxruZ0
jnZ0N4sHUc3sznTbWmMW0lMsfBHIfdT8KuyMY2n7dxLhvxi5vD1aLxLdWvTPLonS
OtbQbkU2pdyly3OtzL9TUqfY3IXvJ30V0VdmAIiUsCJAEkOXwZW3eUbIaNpU4mzE
beUSWxg68+O4aeXzxhugnU/WYc/13rbarsWsyoKDiVRPw8TQhaol5zfXMLy2wpL5
Gu8i4PQISA/w8KLGVCFkjTFz5jqkHJqKCC3VPB2mGmGnrQKVIbuBOgin6HoFknkd
Vs4UKTEHOFiCdYSBI7/ECtuEw/rcX/2/40APwIypu9CyZuAp8ZiwUG+elaFqh7s3
lB3+au8DriGRiIuA7MQ7n98EAcNEKk3+fdnfqxWdRheg4M9+/Kg+7L8asB+0JVc6
Il48naOqmTtYyDuETcSrOfgplmTZlj145KScRopivQ6nv2o53HOxESONHIXeTWf1
OX4yZnagJoF7RoZlKIo5jMTvbkZtJLaOF/6nhrEILGb4/VOvYh3+nR/KGcwzYlVO
nBCk8BfCvBSuFg7l005Zmca5jNzQk+lfzwD0U7RT99pcQ5FPO+WGZbGwtfc6hBFE
IsguX6da9gD9gAT0mKSPo0rQaohnWK+CcPijM2AWu1gSx6737SCuO31ixyDjKV/l
/0O3q5jlvE1kvnqLwhOCLFp9zp3fLr0g5bSQTEc+nMjfYA0RWBiRef2KyCLGrJBw
hqfnkD0CTViQGtrosiqg8a5SK+tbyfam8mQ25j9DnXJB5LDYFQY1EgYrx6PpYitr
GBeMzBsMVbpBuh/hMAtquNX1TEkzvws3yLf81PcyFNAts8rb6TAZK4sOWiml6Hlp
wkkl2t6clR11LlGuVbb1yrytCJmIHhfP5nx0zayeFj0IfH5IghG+huCtIjrWwvpy
FTehJMF1G9xGmkEawZ9DhQPV+35croCHLXR+ddZLLZV3JieRBS9TLw0GSwbPEzlB
SE8kkxjsSI2PTUGR0GuyvyXXk7nphbeg6jNpS7bv0PBBqHBDkl4WI8o2QZx1yu2Z
YqJ9YbyZjN/WoGF/ReJJdxjcqYj48Gm7U/IKlWwXwLG9xypAPaKbQeH1opr7ouRS
JZOP4TgURSvcWXeVJ0ZMT9I4WmfL6JNCyMI7LT7fmeTyfDaHgrf75anyhszpoKsP
nuylp9mspYj4UfDV4j40OSMPQyLoqWxtOD2vvl23k3vAoDqGR10BjFPaeForz31D
0wXZmreslpgIxDIY0W732Ip0U1ukGXSRlDYlNq3/wPA6aDxiyFU6GyMY/W6rhTDR
9XhY+UPrGfVlrRQQ1hJMo/kaV/6Lwc1RRHCtf2YfSzOEYqnm7nrDAKt9G0mmoKO3
3rjU2qXzly+164rbyeJ2XrVe4d7ak8WBoGrNszkUXJvpYwzpSa5a4xX7wW10izCK
gh7PdPWmnc+4nPetMDeAuZtSvQXYIteEiA9DgPsATZdObiovDdJcTRteK0756/DV
kUnRDLxp15IcSYyiRHO7anjpzmZB9hY3fs7f5FiyDmo2zZYS4TC/QKJfc/LIshO2
KJ6WuZNWkbGw1gGsbCmZ2+dsic7XUsvNgjKy5xIyf+0Eqogdlvko587g/ZIaSTIy
nh6+6fixe7RQVWJICbnDFlE2KNjtmCW27r42CKCR8ROKnILMQTBUCzLPyOIoP4SQ
N+94fSsuKimsny5TpHNwFddM403t9soBw7qITmMEuRQcvbEwC0vxuJOZ+8dh7cje
pBt9ZbM8eG2IR9dkCvpQyYngFqxpRpxzNnoPR1Hv55HGPD5gWDdV2wqViWUt2Ahz
PCQA3gx2APueVIbI7M/JbuuYpGoFXg/j+vpZ7uscb9ciNOJXJ1NnnCT1v83ORe4V
/P0GbenldbaekUivmcyNjiKX6GBn9FQycqTpvo8keeFqWwd8g2VmkcPNmAL9JRUk
YMYGgwkhfe7JQBr78VnXNMGj+5iIyTqnlX/nMIaZv1DOyZW3BrnWbbYSkG0r4HRq
Og5+3rrGO0a/DGcjAoNlnQqD5X8hN2r4fSdbCO6VR5RtAqdkoIEl0URlsFVNmbTc
hH4tNPAY+1eX2m2EwWWgQXzJnS4P83lZrpdT5oRjrU4AlyEie3LDyoHKEcvKBy79
ZKn3xX6EvThYAbUKpBOTS21aVkpBOT/6vLMQV0FmirQS+RDgbWnDkMojpNw6OxN0
x8K7Jx8hvgUztGBsBp5ViCPYkfAgAla+I+BnaZDhMX0OC8kHqPTqIntPv1RhTjsq
Bus4lgTV2Z/oMHUD81bDQGg7JfHUVGuX8qF4hx1+hlwzU9VBuCn41cR0zhcxnHTH
iMi4d2LRbNupG4BpnKc9qRHtiSCLRfOFCTF9WLbCY6L07KWqYmezZqsQbcS9zmBQ
QEc5drxTqxqLjTsLlRuBSXYqDZyhuPu6W0w5fBIjwuY1BEUe4IrcW671GrE1E6LV
luDFRVXn/0eJ16lr4rmTachMzxEgRhzuBXXIp9jzhk21vWMK1phfAd0KZqIuYj+r
dDxQQUtkHuT4T+zGfp2sClbleUBjN5JZWJP4KQePu/Q++RLf34ahHwslv2hPo8Cn
zegW68AglNiqUW+sENYRVvL/mkfNpjGIxjBsGflgXXFm2ii9NaFVrz7CealmSDZF
UOPV8fyns3ZOyeiqmc48zGov9isJnGtdy6UnEqB0zzMCxEri+zCTl8LEhjRqh+7n
bHPER/OIp9jJ8+PdsbHrGkBmfVirkCCWellsoCgngUfL8MCSbuJyA+bEeCBKWUIv
BXWFIdViQbP7o2bWN2MNsq5pM8xi99TatQ4rMoMxjoD1SD99tLnE4ai48eX1xtDc
Jq8rfAquxpfgxI6J/he5pw/CNgFZ7IRE5MQSqwbUzct5rXQpd1Uo+YeuATSDTQ+L
WnhlUPqbSnWvK+yQ1NN5xzVBobgFH7j5wcq/5LeDVFXFq4VuveQWyl9F0hpW/eYs
2NJ+1+pmgCy7GLj0mvfXgjNBWv7YQM+HM1E7M6b7FmFyRS/sixk++l3v8V/onj0J
H5+6bOjPJGvgq4EtjRT2YhOSvLLNFWUQJchozdplvgslXMO2NcXF0e2E0ouVtCtc
tYJFBwpWTQOGIbKBanzmzdFUkaW91vnxoydSknLo7Zk6113ZHR+mXp0v0ZdCRg54
S3O+KydUeE8s//Gdr2r7wU++3NeLtY851mweLOKucNTcjcnYXCqEZBo3mwTGqwvZ
ppMHQ6WhYsgYAfvxICfIbiS8i1Z7Bl1CycB5RvcR8+DPrEgdKENg8FjPHq2/o4jF
kkqAYYdiFBCh89OxTJwnL2mnZfEUwjoRAABs/Dk5Az2pGD5sbNtThtK2jYWhJZ4e
gibml1jFeGPa2l6weGiYbQ4Q8ZW9yZeD5VDW2VBVmqm0RkdJfytudUpbNQyebjeH
HBaZvTKDeQkX3B5Wflth24kpj+HW2bYdp0TB5P2NzrzMepOrpKRfn0BiNJXm6Vnu
uj06lBPyOqKB/mibFgNFflnWjh13wkNEccirwBbk0hYRrzFJq6epGE2+WrTrSjr1
HezkdGu42+WVt+7TFcuFwSUH7q8jL/8pM8XuOeSkvGhf511RfQXmD3B0sEteav8R
AE2LcGNkFs08pc3De1adH0Fa183T7iDJnadA3txjxCxAXSkajDOzHVIZI502Frma
+e84rvts9pCdjbR7ccSQyICfvag8O3F04NDVGbB1WVHmhmaVPprhxAyx+M+Fa+vE
oNJUbJgR3m7UKlamRDdNESlT4yjDNjTwbv7pszbpHRo27XLD3hgTm5dJ2v1qg+gA
xepzBLHDULW41rojkQ6+vgG7NbuQMVmp5rBupNLo5zzdYTSTs7BqSXvAeTAsrKrl
2TMYh6p1g2ZjUYwwpzhOVn9uGbLTW0+NQN80yjwfvSYuITMmCsWrSEmPwqOMGRJ+
XO317rL/RN5G5IN1HpIGLSGXRAAnNYm5YY64RfXBNvwXB61Qh4RUym1/Uqk4deHX
m2SxX08AkKQjEQRuyruVNu8RTMeww3pLSN112P0PwvL4uO+5QhDqnDYKqphkvehQ
8gbBCeQZzbDWmxVTAhg5f1gfaBeSpgVwSbeCLf/0kPzR047qZy6kmZbFrw9LRe0O
oGSBTv8Gbs5zos7cbeLBQzL6jgVX4vMYJb05PBAKaGGcWyz66RxPY8rsO8UjNIDR
Ap2SbCKx5ue3yZnG4v9ZiD23GrpamfHJQEIRFIMKqXQr5Y89wk0vGGQOsRIVDI7F
A9h5vcckVZyYyBbNfx7Wjx5Dni/TK9N6ly2bAIKfmpUJZIkEScOs717+R5QeKP/p
9A1Ke7ek19gTfyXPHW+7sR7RDum9U03qc4byrWc7Tl4N1TwIbYE8QY6ZUkvIbYXx
uON5AgEIDnP7eog/x3pN+gEX4vzoeWoFdn/SPiDMH7QZSMpkwnCG7LLY+CIVb7Y8
brXalI5AkZkRVUonk9+nI6sbFOEQZQzfXTwE3FPUSMcMsyR/N0JDy5w1gms71oe+
hvLyRXXkUifrA5m9CCyAJxWIXbtwCeqUzxtF2biFuIbtnTVH1jsdCTOvpp/6vJPf
kR1718P3ydQgHbAVHyaPDpJG9PdZsgJwkgEAjbYhzx45qFLi4xsA+FID2le/C9PL
3JCAZ/rNkpshjRxTavPhb8yXXoiMOEGCHL5vr9Jaoy8MEfC0aOjjzR5wD3btit0n
FtOeW5NMjVL0hdtA4vGyzSucTLoZbfLNuDz3rtYLfr1hOKeJ9gsuKrc19eLvLqVQ
Uu+9KIll8U5xHcfQYj0wjXv5gkgU+5fh8/NKYqEqKNeIA+86m6yWbYng1bkSoik2
5YNqIYDHcNteO3c4QZlmnH2sNDGRwgI7nLgoiHrV38XAnbYn4FwA/L477jgU9K4f
7Msg9KgT663mD1U7dF0l4OdYe8F5AcZNZh9R7UNqsWwAzOo4JuQ1gosSmyAqwcX8
P5sY6tLWr150XZvr0Dd0/ekGjUazJtGPWD/JBfv+DCuSJZy7vc2JLEymY2zSgNy6
Vb3pkm5U3vpRs/ScqBWximtadTO9B6N+LNQCFRVnrzzybN2tCE2lSt1WPaFJLhrm
9TNuYw5RdnFYu8lBIqfVFjTlc0eItDTdeHxUwXLYq01FHO23gC1Q7VHTgcqbT75H
orBBzwogaLj7tOG+UjLVTShfcnQMmBRUCcWmO2GlEJ5eSxtYLYrGH+jHSboowBpG
lEJtqnADJwbwzD+OvC4O2iDhIkL8BBp3ab1tYGyRts6DYS3o5LRHry1i73o34yda
pWkuU2rEAzYkQBMe9IpP6CFysKfgKtdLsaWZEwIbF8dqxBvAyDqh9+EOs8y+qLpX
rB17MrPctfumf/yb/WG74slOvLzmfGeWIyfvAFL17fSRrFk65NNghaSsozYBm/ow
R9rDO110p4ZYiAbVBWuD2QZjMczMgP+wnIjDItfrZHIpN9t58eYAJarOJ03WwZ0C
I23SxbRGNTokO/J3pz8un2av/h3sfLFnKzyn2kH6YtTlrrxUHhzLH5CWSMQ21559
nVsnW7d/8m84u6k7j5mOA5kXtQjAfPo0o6Q78g/k/PC8puclJQnZ0S8jtSboP0Jx
F6isa7r6eW9h67VtU4gRJZ9hjNu34j+Iuhz6uLdsikfKkh/AKDb1YcYSpg7AZKZm
FC82lfjGwYXd22JXgBVGTdlREHTZDZ9eEw1UrdgYBzGK/U7bkAw6mqPqqyCVYlv7
BhEpq5CVQ2fQL6sxb93HX9RR2zl0+9WJRno+OvCXJDvVAUGi9BKfqgruMDPzVebc
BKvyrmkqaSmTFM5LyeCw7TpLPb5pF8fzzgIsxdVYYOlqB9lQF+X8u61lntXKfA2m
xy68luA1Wmybr1wgdZccR+PChE12tjXKDearpxj5PYi2XbHUOTIFXc9FPVC9FPym
FCm346OfYXRukEVOcre1/oyZ2Md1LfAW2UKH9RGW93TNdofGBaVh+SiCwDAfbRLj
NfgF0KSYh0Yp6xLbwNEXnK51cVf7USl1UwVziWFUtdvyVVyGK3ekgjlRf3VVCld3
Rnb5TYsoTb0aSQ+o+tDzzSWOZ9Ju2Hb1FWQUiAwNGbaK1YmMNGoy9ojHhzg+Y0H7
24cCx6s0eYOAFaQoA4/4lHP8VNZU5XoaLN6SXP6vSpNNvWNu5nJYUMSv0hXp4xtj
Gw1fwoaVA4iLOM7SkOlSpJr/owBFeirOYgZqPnYkR0rVevN/Gom4Nkpq+q+9lcDz
gZDVuJOHDMO2mm9CCpJo8tkK73cS3OsH219U+73g8hEJO1T4iphbzLUxEcMY9eg1
0voxVzXvHKzytSPAYxr41HgNsByMzpUUK6XBlri+2efZuUXrTNppL3Uxk571lA6c
isqxoeu8Tq3CRuw2167kQRMPat1U+2ALJya1yFqgGsMsdBNi1UA+bLTRE7I3bYcO
yueqP/PQmnUc0+8yi8p1LwcdI513JabvCTg5TiyrS4lU9CIIHZoNpPFW5dbGn25y
DO2hCsnaoG1hfFpdEkt3Ff7tRW0yuILzbDTZizWUaTQh2PLxpBzBG2zz35c0NroK
fetR0DkxDRfAgqu7bJSjXHB1sDhF5Anl5emkP4vOcn/753Y223GeHIwET/QC2zYc
EiNtwCQpt0wL/AHCNs75Y5DWeX2uF8f8p1uXWQifRVBII06hgx/UmA1RihGBq/87
0fPW9BmqdhwyFltEdmL7qHaasB+Hn2a42+rY/3B4Mut6louIyuaAoG7bPQa98Ecs
FunPAsQ7d0N5bgusl2n/j+xeT1zAD7aEhFYqqM/1IC+ZKHXG++c+nNz99ag60uge
rA0htXePGfC1fGcA38hgkpRYw/Ep1hgxTpyS0+gQ/bKZshEBPJr469WUY26Egr8Q
tMqBZvNKvy+fBm8f1EQ2+zs8nfn3DGUZlNn+160EWTFvLyY54NqnqBQQURroefN6
bmMuXILwmwlxdLObn04+JWHv3X175yf9uhR8o3jBjXBG1JI0jkD2kOCBvjVU26LK
htXA24rLrfC49SLtZjCe+M9qyxbja6RVps9P3NhpRio0Kb4bJy9DTW1AMcKqgSWM
dPxNJ1q8rz5hT/SiVknx9TnhGSNy/unrZVD9kWxeFSno+we0/E3xsGOqbwE6BBYI
Idwc044CVijJt72m791mdsD0f7xFzcPyKOkleJ+8KRedXKtF8TuVCPCdLjgy9dxn
7FCemc8TxCKVE6DmPPXCUqiToy5rn1i6MIm1zsAzZjHz2o/2sk4jeFFS9NZfQ5H0
goxBczxgsrlx3I3UTHMgcpTaAIPH+nI1QUD/UeU1t1zr7z//XQxTNj7PK7hdGuph
Os5M9Anw1Nc8Zdc79//iqo0MdLxBL4UPVlKP+a/30JHjzmf0WYQlOA7D7/7SSo8u
RtVxomQNYrJT2MQqFM4E1XAchoMWwUQOqpaIn13S7A1xn13SHP0nQ5is5hz7G3Wl
AtAgtkQLClYwGU4lm+42WGmkmOX7B+XF7AzwU+Eo2QdVCqX8CHwb4LdO1wSs6OIe
N99TLcQhYpZ9JbNSixsnYdEJAaSpBtY67Dhb2ZX+prIOkSPfSn2lLUf43NbGWdXQ
2qUXAGma5yj4hOidLUyzeyngPVtov04y9zpVGZ/CPbcBupdZUwAeeJrN0oWauoLq
7LgHMJ9FrEAgpJe4kOKS93PBWjvR66nwsWBQvB9Otsx/OOZ+TRfb6bdYgBv+/ASK
gd0Xp1nOsPYJc0rQ7sl1CJ0opOB852Opb1F5u8I90KKP+0LqAuNfgE817kOYQF9c
T4ssO8AiTD2KQCd+mjOyhHqI6KnEf2I1H+5uoZMy/Xe0nFGkphRMi+32yT3BKQKK
SoBSZuAg1EtABqYr5eACpRaBedebeJ2kwF+hAKaa19CXXbx4gbKcfqHaYs2xBzdF
QZ4TX6KmoZyqNX7H0bxrys6350l5uNizCh8Zc422Ef7sBx2BvwvlVeP2f0kJ+Kbe
ZZEaaR43WZ/uveg6TAn6sN3bHPdnnCjy9MRRb1MGEya0YgHhjmPME6pahsLs0AZ4
+/DuzH8+iORmPLyb2qKOSCiBIF0Qyl4lVA1nspScZb0msxwZ2ht6r6Rsdro/aNXd
gQtgMZjlYqouZJJ8UWadUUXub8Zq5UTbIrunZTrjiJgbDQOK7OMQ0MMqJIReNDIt
yemwvq7NFNEHi1Ui0hpyIWIVGIF69Jkd77zgISQM3nHGpVCpVGngRlUAhPkHlwXh
i+knM2R3hC++tUQBcdE0wtZUt9aT9bPF4EwTY5OTS3qnlMndE3RFwwliHA1FxXnP
lLCOEd+OCa5SiN8/6ScmUFhcCUZO43npyFsuG4Leg1iE2/1gBD7t9qX0C1YL+1P6
RoPNwUrs3RRsx7d0Kmll3NkeTsMp74aSdCnjmpY1THvce3G30pdIo0Ps+m5Qrma5
SF5kFBZ2Na27GVimYLDln/O+BNwPuP5Wr9sLafoQqMQQnXFWH6y4UEFpqTuXq+uE
Xdwy76Qi8VFmzb95HBuSrb+auctmbRBCIdNw7i+LAba/r0CUnN1CUNSERa3LyN4U
ddUzTUISCgPo1k7tyaUB+8cFvJ7Rza/960CNP1idGaG3g33qg5p8/NY94Iuv+SZa
JD8hIkvgyfwkS/QWppQUBPAvBoORg4XITNlSk6slNnHQPaU/DtpZZz4kSZY1APVP
vRCQVkLeBroOonYPDXHyQN+0oafLV6M9+GgK1rpU0n2OyqR16yqmWBlTiy253eJ3
c9YUsU7VYQaJzSGm/lzIZ68x11KwAEuDubyAs6u6NERiLiK1xoIlZETADV83ttE6
t9YVx/uee2KbxDZ3rBaQMMwnx8pjKmbk7111ILR7YZ4drqdqHbswrnL8ofF8n027
+InQfUYSApIveVgUWj0Rp/m5Ru7v5C9dnjs0eLwH2CgXIvhL3PD7XJaWgI6Cl8lb
KF2LQwyzsczHrBtLwOG+2MiVOHSO0JodnCG4ENGl5wtGr3ff/fH1jV5ML2//GeKW
+Dfa2GRuvuxpF23abeEKt1bF1LQyjGVNHw4P4DWz6IvCwCG42bmmZQsJ2uqlnqZp
qTwGFm8L0dubK3nQIBFQLL3N4piYkXaDqVkeOfPh77U1DbHLFePow5CDwb7UIyY1
MmP5g0Z3Onrgq7km8sSJ+ulfHBWH8gwnUYbrAjbEFsKdRfKmHGeXz+udZktoDPmD
KpkD8mv6RotvCxQ+H5uzv+TVBa1jVbgCw4q37MhhA8+HI2zmSfpWkKGtMERiADoN
vExd1WQA0zFTH+qVIgfPj7XoKyiGGRWRCEfiaCFL3mPbipDONJ59ZTvrTtE5/Twr
S7aVF/q7fxPXypMoNBmNpDDALGHzi6oy6SNu/o3A3gsi6aDqXkUOL7Lk/Z1IuTcf
3kLBDobbKzGdbISXtJMMm7WznTgKxZGVyS5QHXR72IzaVfY8t8ha8xBgUahTveE9
GoUjes5HQdqlL7VcbCkB2+NtHYQPjoWkuVQRGHikzoYHKH67yBYqbkFuk0Ig72qw
i4f2VVE7AdDVNtHER6h767p1WYcmpwALX6cAWR/Behke4qbLhrdJ/lj4VDD2UOE+
46bQXcG5OaEWFMZ2E+a1mHAnQsFizLOJdLfFtMlEqS7i8rycYapTpkoW+IRjdNk2
gDEwiscUb6DL9L9vp2sUIxV4cJhpvE1yEo3qtGUa21mt/FXZnq+EIxvxccrGLD0o
yNIHdBY1abKvI4Orq9P5AClv6cqdVaWo3SXTU6NaFEVrgolY2rTR/OXoyDfHXeCg
/z/IKlLyu5+BflJnZ17SLiXzddHSXTuh65tBOEO2Ng/fVlkvUi+2vR0DAsims5Ih
roTz6L+pgQWwpdq/npMTB4ZoyKumt3U0QQ6/9gW6WGQRYt0WixOxamfWD3QF+hhB
uyGQDw2t/4pVBIHg/ZiW1snOZtqwG1sZ/TEL33JIz2xdyij03JrbxMOJollyAoXG
ukTaxDTsNgR7oOB8fnO1177vTfDgGh04aTNa00QbXRBvczUBP+lVxMMn8RI8KYhe
/zWeTDf9zLK8Hq6LELgXXZbXGosf41Qndl+E935+pjrJWgW7gNZOMeeSY2E1znU6
Km9aKEgKRi61b12N30M/fBnzsJ5hdNUSgzB6RPKh3L++deVpvQi+XKgKvMFuEaFT
ios89ZbsgF5ZVLCJFVxYWgZA7ghMcpdr07lgOAOBucDh/MXuIBOssuSUvxQXC/iX
vUL/SkfI1meL9OENvXjRmSG5icqMddDBIDb7uulKIzn+0wib9PSGD3q0D0Scu8t0
i5FyAlKn+VcPWxYNmG15bt82ZITj/csxeoJBUfpu/cc+z7n1XG38tCGEnhQepjZt
3qAdz4hdl5L0KeBOT52i934CRVjYEuqJE2VXauBshmyNwt5ibNFMQZDfrT0seoPf
XYNWQzBceAjE+MYCc7YXJJhr1SbSuLjXcq7MBbcUK6MernpvuoOuYiXfBhj2vxN3
hV37U3UzUGNeQik8lxliMNAj24B8e6YsRDuceDah13c+abVD+jtWK1GYlF7QfNtU
35bXpMpfe7Zix1za8gWyQgHk8nKOnzl3Om+VhO4ntplSx/ChJWpCgCBE51/yjwH4
sxhedjIuu00UrZwmWrxTI4nbVxVC3a2/vLbVnig8AFp8+jCgL7OfpvuBcnvCL+t9
6c5vccOPZVWfzyZ9IQTRgGAPINX7praPEm3sjTA+y/4x2HwtHu9CmwKoCYogAyFs
nbmbAZVjibO9/CJ4bz2vGaip1nVCw6Y+I7fa9IOalY4R2EiWxoLc1+sfZsxscMk0
R08gAGRQh+771Uhp8V58NOh7gXH+Ap5Ef1FxgucAekXFrTMVKLt19mrIhti6y14p
Pkh2OLzROYQqmWnTHSgVpcDLA6JH25FTj/vOkTOP4GiKbK4AHPe3q+CnNW525ec8
3BWriHa7uJf6I82ZPMMeJUPQihGTfxPCzDiHlYRvoakyNG7PC9TvRa0ahlDL2Rjl
4pS6LeG/LGqeDw/38KwC1TA5e1RLvwF/7D4IzrNinMLYimvQJbYWTlA65vYTgltb
5okMcGMl2297yv5N4Kg+lEGS5UX+ziQ1dHkGF77E94lT5t0nJqJ9DkOHtG/4keFK
PHLxxBJW/5IchFlGq8rClF5PUCRG68RyssMhnw+hua17BcBpLNkeFPQ1nH9H3cw0
JOUhK9du10EluaOuUnE9/WvrSBSXhBIEfTHI12LEuJNl3+bj+aurwNIQ59KA/7uV
0xfmW1Ih1qARVG7qsgYjDzNWuHWcnQczMNniMX9uUnPcItQdBXZTbSAeNWVKdfMq
CE+70G7bH0RDoecCmbgD8Tgaba2FVk5FWeZaJuvagl7KAuHhkAXIQsY5CaKxkNTn
WMw+aQTN1HAtGbb8M4we8HzNYNKDYk+1LBMHwXm7INq/rNy9XuIi80WsmzR/K0qL
sEDp7IGUkSLSIW+HX63OIW3lNJPGge1DEkn6PYS9mcKRT34ipq9915qtAFmFBy4P
mHwFyge1w99qX70GcO6SUSTzVeOrpb1UtZQpYTnn/j8Sg94/PT0KIr+UNAgCUQ9+
BRBUq6biV8RoLB8kzZcGGYRVNbi+j7wgO213kbsGFyR4sCs/SarPoOcP/hqJSpfJ
OhD/psIzRbsIcCIFzRCClG8SelookysS7fHGnkdRgYibVG0tbj3DPU7mS3S+ePMP
YT9H8EzvunrRPmpfaarqrXc+wi2n0ukDkrp5et78N31qZxJ4JATsemL3oxyKjn2J
EkCp9Jt0QEVAfEzqA+WlxKUs6+wUROVoGxaAVoB2A57SRNhRRi61stvPl2p8NDVD
eJwLauSV2gbY9mKmxzsxYmgEA5HbpoHdqQjj6ZEMM3FtuJKFcguHRVfxtqByWTu0
L7b+bSkECiSfCjd66yMXy8gr1HxHqa9iBltbmevhkUW1No8lH+ULlT9LT8Bh2InD
Z5/Uk5QIrTfZM5/SPSBVy2e2Hkre4aqPsThvkMaPeOpxzEk8QwYPduAAdxPwJuUC
6gngpy3ZcHkdmPBjpIQQ6xm/fMMMDQgQUooQS/1dSO8kldoTIvHZwLctT2rpqSZ3
KVkLbynS7D79QBxsBk5vOJ6khYy6Zn+WpT4e+9zg5K0yQVvmYTywcC5jK24VpS+9
2gzHAEmsvSw5vfG4VsZ68ILXLUeJ3/UWgV8EbiWmVvJvDlUn45xtlgLVy0YJN/iN
C3FzloU2jYC8bYo/9P05ADD6FP1dIqUKiVlVy/TupHLdxNiEh7CtsfHLanzcdZ4r
0BrjoWZT32H2xnKehBKccfGDG42DbQW0Bcwp+WbvEoLF9g+ZX9yh5RMuQL1T1BNr
O189Rav2XVAPIj6NnUO4ffjXPcP3GjWM6VLNKlX/PZkw2jiimWuoPZnXD8FdhCH2
qeUZ+RInroStL18jOtGv3/ByLLydAirUZfYOcys0glJNgHAzhqT5HJSDoY/Ny/h6
ua3Z0jwbtV7U9lgG8RoHPRLGQBxjmJcUtMrg2xbjIzghQzfNNXI7IqeWNLioCgWd
tmoRf6UGbwQQgSkmh9R2x9/HZyrvxaqbbw7GBYJdCGNtGgto8FX43Z8sycDqeFIO
cSH0pUsD3skBSfAdTp/zE/If7Pbc6bqP/e0NLZR+eAZr0K+3wKdBo/AYg8Y5s1Ob
8CNWtoXjr4eymWJG5OtKSN81OUPmY8q7BLolZ0Vf021jX38+OmUQagDCjrb2RAUD
i+qqxi7iwMI5KP46y6/TIghQvN9ZsDVUZUQRFMHR8VThe7Lpxqnls2RHWi+qXW2j
ADQuYqhYSfhv4+zH2bVk4uQBe8Mjx+9PALham71BaW6w0s2o6pQGtYN4w3D8oK5s
Q78uVLIz3kD5PyoS6lJv50JCVBUsZYatsTcKOHfLMCuC5wbg0LH1ZRTrp0Eaf1MZ
fP+WXhTsYU52aWHbmuZ4tkuzwSWKcgxR7cZq1CGkA3YfvDD2rrdqrmTPKFE81M12
svEVjBtIQnfXRtUO3nQB6p8qckqfV80k3pK/q3xREr8TeWjTrBcpSZnrnHfqyxZb
1PY4ns3TuhXFPQvoiv59LVjRTQk2BNULboYdP+3QTZHUUUMKjXAEuNWxf6vh6HqI
l7IcbahlVPtfDixbhAqRiUq2BPz1q3ZfazROsRkU8LIMQLbhIhS4SIrjDRI38c1J
rei7J2/QxYNQC2iGtI/1oU0WLsWQMU4XA0SNm6rDFXT4kM4x2IJA9Ljo9fwGRGwm
1OkyLfN1QMe6gYJawkHGa/J1D4aw0KqcvxPWH1kOVmU5INTpaTiHyp4dHiNBFrNF
dM6IpKTziSelDwoOtp7AWfe2wIE4NlopAwmdQ3ZUJkpJ8rfYAMSyOedp0M8BDNIj
sPFegUGS9Kyq84lGjdl3JlbFzYgTRyF5QDULOfJ0lstF2S5TlCxJ2iPqfJm73NuS
KBGmZX/jBy1Q+xBKgty1maXYe2oQes3AW9LVHZg55ESRvqktqAGXjl7L2acrXZ1F
xwENd6Mzz7k9vv8lkXCoIsUDE8Q1W1YWAcfq4c/oP3eKPvxiUL9l0nAAilj7bwbz
4u54RN1E9BaGHVd0MeRulvbOXvcfRItWBqz2RghbYOQLrLS5kMXF6wVvUHq8eUx9
mxa32DSe/7Q7mYoEFXVQm+66BlpisfHnxTaKCcxRkpryZiBOxgr/0jamMczAXsBD
56pxrp4Wi4ayLllnrSz5Zn67nCwXf6Ca8K7RCLU9OQp1w4cz3s2Bj4m2lcRdyay6
j96DIOtR4LyZIQAIvX7LbqsGhddmpTfCAMF5D+QEdXcUOQL2jiUoUHIXalwXgN5+
PP/pG3J6usLbhS1Z9Yb3cnHaAyL1C9RPmxtfdfDYI7iS4JTvvefYYpUl+MZEVPXR
uJ9ahcf0FHNuB6Q2JCrl3/B6o28B787eZvaEgzwXKuU3a5IbClc5BE5sMquO3w9i
2LUuUX7kRl4StNuzTcjJwLGmbhx138DV6EzHafXuCXo0Yu1KMY+lcyZWSDMp69r+
/oxHCYpFVavXt2t05OBWUfhrNwOGVIxDEV1DS2e0UQMgss9XqfqbuqXmZOk9J9cd
QKoZXp0CZpR6URoxkCOOOxDyJTqYbNEgw8Z8UfZtgOqLa1IvGHzRwuUCMLeiY7eL
gpEhmXl9WK11vn7/hlNnXEy3l88db79mdNQBLtX+kZaNJpbvKwXoa4RT7gouV2kT
9H7UPCJmKc41hdB9ytGlUcrtBTLddvXNpJHIoJrkK/2M291ojFXwkS2zmvmQkK0y
IoCBTZZb1eHm7Innzwc9r6CZ/Q8UMT6YPOSf9bvHMVbbiSeOMQ9dEt7C97WvzOvJ
9JHELe0Vg+vZbTMTUx4ExUH/0XE6R+QJ5xPxx39ts++ibQOctqAbsifDy8kzwP/b
uySoT/Zwg3Yz1yZ2E3kWsbLItJZASuH8Z8pWnF7/O34j/SxDPkWyvBDrTp1d3KZ5
Br+JMHkwobsujCEKzRKnevesVx5LLOWPUKfm2XuFjx3zFI2tawICVgd17B/m/HLo
63PGc6swyRTuVXT337lg/rlWNP236ndGa0IhPxqBi5uL7gcimVR5L/g7EJqOGuqi
mKSxJ5Ok22Wb5NZCpI8v6ZJJNQfs9RqnCg/BFAZBTl+Hl2878Z3GmWoewEmBzJOT
609NOLIF+GZP1uBnGcmAgXmdIR85vfxA3K2qU9oTcZUGHvF0bDboJkEmKYwsKcxU
ofLF7nXiZd83Fchgx+fg6R3XRR1Gnq+v8D7ZIjVoExYqXcyi0hwEchuVeVXDGNjN
y+yYHn2v8rx3uDd6oW0uleA1UUKmlu+cHZvGEpuxtQ/zaP9HN1abWl4LbsnpR6yi
4m9e06hkCgiAzvkS4WH92OGHpT40zf579RqFth2j+mEeDtENWn8B+mA/5VHeME41
67bgLsc0MGzbkF1Hk93SovNfT1/dTGnzDn1qe2fNwx93CmmYNNoY+kZxNdRksS6K
tBDQsZueO7bvEAh6QuYEgAfb60b9IaRTIjU0Q9lB1ULP09HLpga9wvUDO1HTgQCj
uqLumifzoIOAE5KfF2/GAe132CHO71F+IWVWK8YVXeAJ1EnRlGAUHvs5nMVSRE3e
NdmXIbYG0cctBod7bSmz/HAgBZFi6jPC7BjSpcV9b5bhMi7WcbiClCN/EGjwpsDI
iGUsVaRGTtEizmFPWEsdAU5sEr5vON9Mu5SbN2ioBVZOyJv8shKoxSH3MMLeHvNx
IoaMq28thrTYjJgFWv1bfOC9pCGWSvmyr/kKqr3HNWQCsryzEFBQ8xKHshwTulNf
/fOGxj5WNBT3mc1iMgaqEtHJpnIgDMevZ/71y6VDp62DVG1YTdLE+R8GSgZFrhZY
+I0Za0LzMYD7RTgpn2p2R3t9nJiZhO+GKIevSwYAAaBfaZgIWfRcIrpxVEK/+496
Y/ozhNtX7IGAG5jn4qfvMdMM5/YkWZAGulWnhkADKgHLkLXtbxbOEc4FB+jlqNCI
/Lk0NdE5vwEI8UIabLg3vSG2XKPVGFHgXRuwW/Ca5m91ZKcZg+yRf/lgwFg3E9Da
y7lS2/dKPjCghwN6fFgN1VZRI8JWmAukQb2Cx4i0GHpF3reTJaxDtPKLvo4pFgF2
DYujIHWSqfvlxcuXEU0L1O2zrAgwgfUJh/Ad3QY3QkNyW8WURADUqBkVYb8fRSs6
yeJlZU+bjN0TwNvVgzt/+vmEBjYhUiq9LBDcJiL8HBNHZR/VBTj8OiFnvQhcbWFe
ACVrP4PLBpOmmXJjaab8N+1Nd5I8SYYfZyFNo/QSfunUs4tNwssMVzplmpN8uzGL
CF4uk4cKVAhM+hIGNrN/nzv5GCRfE4TQ3SNoYI3TvqPfgv+kUVfPeoAGj51vYKdX
09DeYTbEnpn/kRfRA2HPBpu0Fa9mXQSmEYulzkKCqERj42T5CiQ2asOiGDybL5yN
S/eZDtNDOJkgPoae24pSKxppZsxbCaCZHVFnpwgKDg6PTjqvWvCHsTBuFh7WsYEe
ltH1nkBWuEz7Oj+HbIqeGCZVIn/y1pPorecCWQggK3anAYHIgfxgvqMhx4co6sTu
bwZBKfPIENeHDBlAdC+HlgIIdqfRKu69oOVcw4KtyWNJJ5n9WkONwyMIPnyhpfIC
EPRiBBJynLt+c2CmPUuNmMsLWSuge8zZDBeKol3ORt3DkLoGz2Vg0HHcHtBTrbec
3gAKEHd6BE/3eIL8013J3zqqWh+eAKXc/+6UnGncBmUAtKQ4J9K9/GHoR23PQ1ym
Zus43uUbPgvkk1Yf9uSAw3ZTTqMbyYAFaSIsjWcQFJr9Br5fwMu5D28iUOVqdqeP
umpdCvbMFyDDf7qJNauSypYCOrP382S1gWrTNqvW4OAXlc2+ToLT2jl3CX0zxgyX
TYZXfM6gt8HVxLO1SM4wftkxNJLIN2jmU/2wmXY/kcsmGKNCxYoRZN+VCVa1xpqp
Iv8AxPEjZEwoCcTAKobZ3V3eECX5rAbxhGbut8CEQ6Qh+AB++Vt2VXaTU2v7qniD
5yxmaHYv97tf29ev0saXJ/lOljN3pSFI4bJLOaBl4HsZAJwisih4Aj1CXCY8PFN6
dFfeL17sbJSekWypuKbd5/7G3kKaK+H4HPfHFuEkIp2Fg340O+p+wb+gqLLXICTO
HGAOi0jPAXyucwNc/v8mDfUNsoWPTVTo/Jiu7R5bBQsa3x4qiXcIu6UJH0nEqqTN
3/6jFolqUPtDL7npb7cNckIyUNYQ1lCeW5AqlRL7Gb8jLYbAOAM6lH36Db8cloRe
ketV4gbjW/clFS1ReXsJoVRPkXOHokeHTz3Dz/jVTuKZAuSN5Y+s9FaWcQ+dE3gx
EQZSTCtxgHUNaNS+7zi2Ef0LCQ5klrnU1XzSMxxjPGoDFmZ/t0SuJ51D+KS1/Y/X
wF1maKeGqwI1Bx3HD3bjwAKv+ozZ2UiXnJsdSF7VP74eXts1fIxAFlVDWqINtRLO
5bY/m0hlQBvsoWtfMJsBIQeGD1V7kQtZYsD9guYigG3SYFL4ZYW8QzfNTQaYJoQK
bPlXX4PnHMzHBDkrkRb8TpdZh3wFZgWxn7gKGG5GxpJSYaFWhI1U7YVGZaHFE51A
ANVzAuewfWz+XhctlU0FXkXsn2uAHz+1rMMOtiYIPUzjN5y6Q2BbfxNKJCouJdwp
3C4xJK86An3YsonEHrsWfxzo4/LTRHmKDS8QySToJBx/MD+w5TJYKbj9oGB1zgWu
j1ZzIP1XKuRIwu7r0RD76I2NQZwnivyOrhI+EYquAN3bKxR1q16F6XqbWtM4Hqv0
oIuugNA/pvZGYmr50xx10C8vWxJUQf0F58YWJDT1OJm5LYB1kIhp6vWn7pmBuP5h
YwS6wfUPNDNmx6lEVBnnRI3zb6nqvmE9piiG4kRb52S+qa/aPerBPWZXad4e42E2
C0Aj0H/mAqrNRLvGwEn5BiNOa4vYd01EStLT42TFkUjVaERPnu42xdTxCbNTIXCy
aEFu3KQk9fho5adQ0zKxI5HReQcAGRB47c1vGIEcAGH14oDJSYsv1L7XDVAZlAKJ
YZIYgNXbKHkIOu/M6zkjvaJW5K/GXrGAasDfiQr3OBgkqx4ROqxp5A8SSbt898GW
4tj5VjUPr0V4HSshLCxhL7k3etk9veHUL45mt6156pbJRg9sE9FYm2/j/XKUmEDV
vwqK2MbPzkgSj6QALUujHeXzvQISDXI1Q+Tfso5VfJo2nnxvmwDwuL2GUOlhS+qi
eQRXciaGonoBBYreZafwl30Qqnh4vT/UeLjtzxCf2PdVRg8V5E2NJfZpYl2+kezt
gp76TiBF4LV/5d4i2UCHoL6js/uOrrqTn+eTLIRbbnbcj5SJN/5enzbcJsJJ4ryO
4LKb/isXTuHRPaaPxG9okO1B+/fiEn5V0IAootryYc3Yl7z5npf6BgqVVWd+VfxW
9mmYmHBaVISXmABo3031A/0mhqTQ/yt4ljE15RMvT+hkl6tkmi7ob/zx5HNnGK2v
soRBR4dZBGdAV1sHJAPTs8iFKhsILYvGpwMcOQeP8rlCfS9pOSYLPehFWviWIzJF
EmT1NbqMHPrg7kT3mlt6+KOSaOfrfmjabdGGx2GEWOcf6DUKwRuk3FWAHcqVND1I
WzUNcdepVCcCIeDQnZACIS+T/PDv8eljgpqW8y0cUFZ2LHOWXjOcfWAwzdzWjijv
LrDOS37ZksSPqc2CUqxVvvHNPEtVBq2ROd/bRAZsbMDULUVCodGBeQfu+b2259FU
1iJzK5Njxy8x/fX4wGsR7qnjbuL1z/5SrJAwjf+hUqw6mmhYrpqy8rbr+KcjSdhZ
j3lLxg63fzwchMrdjYUOPw1VcgX5isu8OskpdiUC9iiQOSFgDdjgu97FLLxByWSN
MCoRwFFNJZUSpe3xlHiInzjH1GoSnrf3jSS3MC8WEcLEAqhgjBPlM0+664xjeliG
X8WaMoh+x65y8Tce5fuU7OWlFqsZtMNMkbZ02DwmVgSYaJqVGWCW+m0xFOzTlcVb
6O5i6ShdZ7jWf7c85/iV7wuThgnEdDqQbeGjeCM5Gy55oWs0hS59bcKBLPxCz0N3
7w+URQ2wT3HmtTXdsoo8gf8X74pnPzFLXX4MAHQqwQ8R+n0m4iooJJ92GV4j39aG
ji5BrClGoXKj3IOfXvfE/8cPLVb2dCi+OKArDzRCeqp88xwkdHm5u38X2LRRY+EI
+dz9usHSCF7VxP5IQtwaxomCA0KH+mo0AzU6Ylr55RGmpAln11SkjzXAlbrsReZl
t9xY9Pj6GsODsTQeEvad46f0T/earS2bnQsEqLLnm6KQpB704InICZLLLe/JLNBP
3Ag0Ppv/YvOI3tciMp0q1FdlG908oG9+aCViWi+qZAwFDcq1a9+E+GuL6f34kFxc
uTUAqpHFsfVxwrIV68ictm3rCvGEu/qAtFcxvv0fPUSGpHAax+jHup+UZ+Ye8hYc
eVjaKyEp0QDyGt5aDRZXJ7ZCIocOCAKMrSMVKdhF5EUM85+9YQx3Mqjs1cr5rmso
nKOScy9WgWDRj4GITKnO7QDMMNRc/H9JunOpivzmw7eA5OQkriOK5YGT/EKR+Jkz
FjWawuVfdTrHiXlQulcB4z2iCpyxuSWvRqR1H1eGIZo9YQdMnAJ1up1cxL6NY1hg
qq+r8m0z3Ak5ufkc6yN+A9TKmJbFJLAKTet0cfgr0YknPUXrolyMw6HfvMPjEjSr
0I3CxxTn4O4BjiVo1IrdOROiLSOXwAAZfIKGQ9coWjn1G78NNHY9HFvYVpEb8vf9
BkYci+yfFTGxhY06BcK9rxnXOQ1zm7MXDw5GBdLgnAmyrbTvW1VY6Os4F8PZq0hv
TpWi5yI/6qlmvwIHpT110UE/2fTNHu1Xqxy9FhwxYZ4pWKL9PPy+GvQU2rbxEJdx
HV2hJR3xGgJMb3YucdCTbMoPmpuI5iBh7Z3btCaIUZOrKLC0JxrJuTYITuj5rdC+
9BcmrzBwdQSEdI1QLnpS3PxpIJzkZSKKxH1YP71sldWUeEZaR/ocfF5/IGHbUxKO
7c0uqc1OYoGzaJ89kvjBtZQvrQQa/DG692xH3R9qrmGcbNr5dTMXZo4mdYzA7qta
E5LiK4z4nEC2NTifYHrD25UNmOk2h9jWO5HRxnrgOLTwE56sD+zknuupMfU800M4
i55191Gwh0x/U5SAsIESDGrwV7RT+yOaGjoYim9U/bSmyct2d4YSyx+NZDUcuAKv
BDt0Y0vDBEmmkHJiHADDxEyMJZEFYHO42sMMF5rvSCcvOBAnPOrzGbvNbZNxSfei
WuE+bCYSNr61Ira9yjFoQnmy7GeXtPEuQjf6Mn9Z8pOw1G/5qaGMAhIx8K5Df0HL
2Tf+ywtybA06N8PqAltJIwy4Tz7P3Q6LzKCfuaH6JbAEOwff9JSyRbap7GtyHi/E
tcdJAhdgr+4PKt1V5cR9X5zGFc1M15mlRuTFnnwMicVgtoHqMPhl1Xg3/nfkU95E
JmnN3fW0TuVCtMiwXRfEWP6Ht3BSaQ20Okrb2rhsMK4bcmPjGpyAyZ6kasoDlhzd
3phaY87BOfnfmqy/KYHLJZB0nfKWpFe1ugxaRlbLbKxi3soYGNNFrhVFv/ufZqX/
U7PLK4z/CaadTQh+JzDrP38kUKbalieBSpEyAkTrvpjzym6grnUo+0nzj0w5wxM7
DHsQMQANJaWJOw853K9tk3IUIf7Bzi9JmSnwLMRo9gHMGjXvPbYjouCjOWkzILGH
KlQ9qqhc/xhrxYJ6z8FyffuYdCKp4rHf6uCiSLmKBM5qA5ykbGuW8kMEAReF8zjC
36qmNMZo5IMGMAsPnvjEFpMEREKlBX2IZd7lqvkPXJQuTBb8rrvdn7suUSWZReTj
fOsRe+6rL206Gaw03kERVmPr0JTIV2de5sP5L+KaXZ+zjv2Jsb6gjZIRrTK2CEob
UlO+io8+Vs139MpIYuIthDlPVu/uS0jyt/O5yJPa6gjvnOv6N5/dYl9xGxiiJ/XY
veIJipzEnFuOxwJJ++LGAfbhlEDPOsdA3/V1//iPGzX/OHXva53euvtrziqrzf/b
JrBkEMFdKPWxqQ4DVyE7HLDT1SSxqmwvu6Xt/7fLIjC9YhKTls229K7F7sso6H50
iYu8t6ya1p56K3nBnD8GJrPl6KZxutowOk1t0MsqcshUHAKI5YT3mxEUEaQizAFU
BFqcXxHbv3oLiRS0qxr/xruCVQRdw1wsGtpzjRig/hCaY9bJuOedkpuMGIJHVJYX
TBb1PCMEkIbKb3n9ZnYKaamIMxGSCNE7f/9FpnBDkvBg8Kba9RBgWuwPM/wyHQu/
+/N74TV0lxoQC61qvzVfb8qQTnUl9K6sbyfH4OLllTfAGompiufIkrypfke8HfVn
Vqg0+Pu7rJggeXZFZ6TZtYikZ41tTFTj6issRKAjfbY9kx5iSRtjLLmyf2Lcaa7k
lZLSjJw4+mYEG8HGAMPTvTnF5TSxarIWAYlsQOGi3sVnZT+lg0sq+Kqn3Ll86Tkn
azR9WPhEZUvTp90+P6urS5bsEJFw5FJtMuvW0owxP0VvWs390VgX/app+nSmKm3v
zPunmaow02EDcmJrANn9LCmECWHRNeBLKtGs0aX4Lf29dzrmE2XS84JBgwvGIsK2
QEQSZD68OHonuXc1fO/uzXRCooKLRLwMMc5gp4vRzZc5DgdsuB55OzQhWZuNfWNm
mSgo4QT6Tf8ot2UELHZnvN5dpgYoicUFzOUEFUFqKFldPu3NE/pufjnphXTT7n8Q
oygaH6bbV3P5h75LtfnoLC4p+4qFA9seoHqupM44pAfSuJoELKiLwYhe3xcGHQCe
UU8IlTOAv1AXj+crpd7CVbwgnK3I+N+H+c+FKFgX1wSe1tHRQlVTnst+jJwDeOC6
usUpHvDCJHXrvQ9sanq+VbEZcQXIlk+uxm0NTPVZ8icCy1Jcqi2ckkENzxM5bbtE
JmCk+rU5nmOwkShXXXSO7+fgRfqt57PqL9dbAC6mXaBRfMHJSOJJzhMNr5ZvsUVs
P3SaZgSm5Bht0M7gvTnWk5QD5ihqRb0AJrPrDLs9yqZdxSWynoMAccoVOHdmJpio
gvsO9Un4KZAxJegaIVmOe679K1tZio9xTBk1DoSps0MYPKQuZlK/BOmPF2vXDefo
H/qvTRhqk5q+R1P5hoaoa6t7CVl+dvIPiJqsIadf/B0BGAbiFfnrx9t8WuUWZFaA
jZKzSKITpJg7Qi53bsnMv1sTu3jFWEIdYYCUGHXLLbWIte3KfYgG1F/xuJk0M0wd
DZxPmK2ZUUqLRFYTL5vlQgCV+vB/40Afu2wqyOcCylLIw82V85/CtJhQuTG3yRxh
rH4jwXEQbEMlecFwMQdL5W+0nBoUr2xxz4fRh+1hDU9DcRFw1PlSLUdh3eCbpn92
90tqAMzmgy0RXbQKZcD918kXPA9h7liU8KSKMULdVMAWPwRZuOEBckiDPXxlD8yG
PngJGz2Z7hqAFc8zCuSZw2WTXiBzOfdxo4wagdnV7HmdSsvalKzxEryDhThIzMze
Xbiyt2VcPW2PGwjODqWK8pzq7KP1EYiewyXYzAnIgfwH0OjzTisKw8Ybb2g0pmaX
dXy81NYpMd4XdnvJcFwwZtbYT3vYZQAL5Yr2wZrBppxLWwHFAR7ugmjbCeCHWBIc
0dm0ouQh25Sjs+HFjW5yF24ApnIKAjU0dNjaTrvHCI0ubxcBl1Qlk43gnywIEjlj
x7jQw20BcirU9JnzvFPPOVofjt1CxmVU4gBCqP3MhNC8qRXm8gv+Lc6AGWL9xHy5
XzsV2nr8JpbJGRa+UAvdXoHoukUOQldUgd12g5R9i7ynQxdFuemgUVXmO0m/vnLF
eFmklBql1dwJbPYpPR2fSUEDH1R4YNJtymypFrNPfyX6J1CFP+ULkts52wFBSzF9
3LhyvAtJ0lgBQ5xHNeAkZJEAmzTws7FTmu9l9bLg10wdijkzwt9KBXmtcSDnJowT
UN8B2829iR82RSS692BCexWu6fmf+ZZv+6dNFrxV0dHZ90OfPv7WZLwbXduNJXha
IPEmwkaID9cZupaBXRQVqEkpCb75phRW5LiX1Hyz4ojTeMD1fE3oPCju5BuZWQgG
qf0pvnNwEWWZa+vGwFIIo7e4QMoS5sWA6vFCLDPizctLcNNMM3GCozXnGldVm/l0
8Ms5nGhkMppkUy87mYrdGbnXZL3nbM6zLZz2xAbUMpvaPH1kdBLsp2TdxLamRY97
h62b9vj/kfYoVKsUudm5tEG/h4gwmylWyhWLLkRXS/av/xB/1WJuQAlG9OmMSxii
fthjb+0/UHilGnu+rYJSn8mpeVkb74c2g9aQk4A3SQ8B24lSVTu5Lfltzg0DadxP
eGAjBXjEUTN9BiKkmeQOQp9U7bckuYPjcJEIXaBcGTXlgxtGkp5wE68qOAgD7ydK
ds4Gj9Sqvab33id6bqTskdubrjWDc3YbTe8O1kKS48bwGKeif83fub9z1iA+h/gV
NRuGpxqXMsVWoqvr1hNeDxuP45oVucjSeBJjSgTqJQFev4/IOB/TelNxB0gKyAI4
GxXg4VFSRahP7oz62Yw64nWPl4Aln8DRgEH0XeJttKe4rvrvz+MNlGi6jO0DgULu
umzhNX84QsHFFSdpfMlyNnUTaU+IHGmk8TYU+20kt1yQC1ZiNCzkDjUmlatbEz9u
oMyoLU5yq3l4+mCJWtntI2h1OKowzAJKR1qIEV//iDCKg8OJeJRzNAAocLUf3N9+
+6wgNDXQ2vjFt6RpFR0b0I6t6oqsVL++iaQyboTOaxrYwoaBZSLwyjuJc8lUpdYF
aCh/XqptQQ0kmFVWxTg4K+7Osn2kzVKtbrqk39ov4AEBLOzfyw1CALynMQipqPKd
XEo7gmqHgTkd/B9Hruu70j0HEfGB+364VDSGoSx0kLH+56Mno07kUzxqs7hpY/fo
kc8+kZ3z5s6aP/13YGVfbF3H42sKPg3VJZZWqRhEuCLIlB0o5U3nIAPMOvuEaapy
x519sbyJvuGUiE22XX10aDXqxoSVjPdB8KPO/ZYrRaDL4VwqH6VknVUfntlHBGZE
jMAOIhIWbtjn63iuhXqh2FfOfA3fAkXTmBp+kznZY53YvumEUp81smN8S9REYTiD
zs7QXhxoOwKzstJktEO8ENt5/Bt2biiquMiDQA/RcKHRrhkDgQ0JYiZ0UgCY1QeX
OUAJ97csKIon0rSyIhETfOHb3bPD+Y7aw3cHrtZlwsSl1KsZerj+GDADMR2qtT9q
MK5iK/t7JfUdrBEtRqEph1iyJRAIEsUvIfnnVQ7tvKeDRRqhycqGHJQowgwkji+z
Y9byVExwAP3mwk/tjS04L24rFa//jBGRbc3ALQT98WDiApRXt+/y3WX33hk34cMS
WF3PmWgbgm8E33lCLIlkM+GckisN+r0dKZGwJL9fW1NysQ0r0fF+utUJOujJmXNY
SjSi50+i7IsrSJfb4fCq9cGzMl6iLUTFL+TR98Cv1zvaffWJUN2x2iEB5JCvStoZ
JIlxD7U5eQdgwXhZaM35NAJrj/BUtETejFapbyW7CnddKUp5R+55Y+CaqFgKbVa8
Thl/QhjqwtXiEi0jttOnyjZ+S0CLoFrLLqdFqcxMW54ZnXz94ifI/CHoxdK1EkBW
w5d/r4v6BVKvh65acV9hO8lC02PS2vehbqEJVVz6NxhPRoh2xm90PGc7nLNf1m0W
jTyxQ+SeCqUkQhOvSSKSMx358/u/0TZ5M/YaPPP58PJDLNVGFFCzmvztOKJEM52u
ueL3VJ4li6EtED3D4nP1pnJEmqvxOROOhKdTbvlZX3kDBz2CPWVi7fCpHsXZoSMR
xVmzzZBwD/wILi0lMwLFnZv7s4I82X/UCcCpczCtp0+M9v6J/kWjtqkcbCShktMt
NH1AhymqL0TEtBCEFIu9KbeiR7z2rahEEH0j0oY3mXDcy6wrW9FPe7nyLnEmyrLt
WgSdY0KR7Y/HqARrrE/h+EtnUAS3tBMjRruBSsUQfFIvC5AJnsWJQt67SEZ2XA4z
3HrsGvnBziST7ksac7yZxD3IKT0oi4IGUREkZN6RcY7IBVNOeenZJwMA0GCpfuwX
NHigkmyX2gefTQodKK+pExJ3Ev65+zHJQvf1vhvRhknxN5Du+QLQyM7+YGG2MrMe
jxwqGtJwykB6exJGW/YhFCOURxSdRzPRyPMDB2VV1Da8Mh4rhkX29Tdj7h4Sb0Km
+cyUJ9Pky+KjZqgZcR+M8ITJ95OIfqRUFL0NOurytkP/GPXS+7ZbZM2zeG76tBom
fYymRJGVBZ43EQYS9WZh3BNOeH5a/ANLV9V6A8SWtdrEQJwA8BeygZ0+XCVHvjaW
Fw+SB3XlPGk5WbJCAbJcDS9npvj85CKD4D/YbS0+a2BVonqGxK1v1757XQx4VmPg
WSpUCw56KqlDrHzu4XQA3CeDOyG0Y+/iLp7J25fwuJ0pqxxskF7LcNAXOTbPIb89
5Ken23FxbrRS9gZ0ynRo1wreiGxsBifsTHSBGirBPrm8gnAs2gU9tDOEsPvsLOmN
AlyCc0ugYFo81gyDH83JOLHoQlim7vakuls+urbOs2CJ0Q+7JknPdz33aR9HiwC0
PiHT1DsfwCNW4nbOciHREywizNGdgMqP5bydewrMHXPFpL9/Wk6SVDElOeitjsoO
7QN68bw0szydk+UtgoytCkwfsAQcb1o+Bhrn70EU8aQANOUFvcJR+rBV9dSh/g42
fpKnxh9qWvJ2wG68FRYjm3MgVINnR2OJ+uKI7+8YI/BV08IDwx7o5zIlyLwzs5WS
njfYS8dz1BV49nY5v0J0jZJeiR573jyMz+Bn5QoeuNcHk0YsWs/yNUBX+3BKXV8R
+LArKmq2QVSZmIpB9vdC++xF6iVxK53e1B6vp9setVo7QcEF1dvUm6UeUXDrfAyY
Wq7CE4BrHyedLN1bu5c8L9sLqsWzdC12EqpbcBrwn5pz1akQcPwsqqIg3lHxFH9d
NKoTynf4sfKi6uz1CFvw9Egp1JyhA6quy1djjKUQ7k05SCsUXSpAtF1nK5u9Lq1P
HwRXeENzpEI8NkCdB2sUyNZx2GUOBd9DKN9IhvcigQUv8/U1/iAp91etSEeBqxnn
sg0eFV7sAOMgRAoCFygKcKY6tG6G6FIiuMyByHZIho6A6siPvmWbR1kmqK8A6mX9
zYxJkPKn5tB1T2g0BKdxgVUxLgCudfHdCy/QeJYF1rRQAN7jAK0ct9FAgMaW7MLX
SXjezJvkGXJmciJQjRA4dqRTRB6myj+nvfJq3YvfNMw42EvweDMW5zeOPl4wztWB
jdFxmPB0iDcKC8d3D2auOBVP8zsyV+B7vV51xg6PpdGrEE0zlnOodXQIP3x73g4F
EyMOQH7N6kmuAgUfMarPCS2mA20lnpwjYu1IyCeD6uhPPPmEk0wzZtqpPOn6EHf+
ZS1hcg/67hteKB2VRcBp0uCghZciGu9G05I0y9h44aam8ebvKw6kCufbfU8+Khwa
xLXcp2qOWyJt5/b6jI2tOYH6xcA2cHAGOC5+BokiTdXzdZ9wray7RuxbmM+vM9G9
S0qQc4JqTCj32zu6g/vhKPma7XL6VxFtb44LwFGaOxYqFgrBzV78VYLoQHgnu03f
9NWVFN+/NbC5cWwnrWUDJ/SYN67UDlhvV1a5Hz/ilTatWSX8p7JraT1wXdGRY9M5
TvXrwsp8mJSWhDBIWt3NCRvr3hKzy2cjgzUgqOeJk7v+08nJf5hE8YvPyAW6mgLN
K4gen62GYXMPnlDKHTdJEZ/H+rWxks09HlQ8nr9rcbnUtigB/PdAcBMgSzBPG0Pp
ZVGSWGmLAz3S6H8aBvRva7wJu4ZiKlAD8szmAIYbXNBOGIwC0Yuk5LOk3CUOOTqa
ODHXOyfFAfGw4SJtkODsmwaG4t1B9kJQFlF1ToH+XMw8My5Wvh4UL8vw4MPvzYDu
d4xoFChTCcqWy9XQF8Af8MVl/wFq/Jnj8gIzgbRa41TwA6c9/MWNCypquyCyfad4
TpAc20ZZGjI8rnj22KmZRo9Gn459bCSEsO9bK0bk6a6BhyoE/IbikDaa/5Ffb0fa
TnAPYPjqkcFSnoBwmmCTwkA/cQabMfnrbB7vkQWRQVGxl8M5shRCqxRQ2tpmBQHF
+aJ8k5XFLMLjVKSOZQYP1selKraPPGUGulinxySw3HLVRnx5CT8VjSZ5j45+NQfd
a92cBhor+4D7dK/QHwbJo36chWDM7L5W82LvvrQQcXumSEUEchrHgiQemGg05dxs
kq6TSNIwV/SnVVo6q1gAAd4HHYC7nNP7abSbUOp+x4VYZ8n/cNZWuHMvHFpqL0kp
m7btZU9kwqsZjiNB5BfLK0PEMZ6jFzuuftM3VM3c4Mijbc7qi7ischg/ZkMBhWVU
1BOJxgA4Lg8RrcYQWDgFb4bK5lfn6WT8PjuK27W6eekneeWg/R1m7SLuMvIXXUWp
TDqWQrlEV7nNLdU+ayCiRq+ppzEsRAjpSweXKMHlRxp3/2FxDiRBhISOVKGFPZF1
XIwYkyijpuF1vpe1FjAvlsTyuOq/Ws9Rc9dwVMAodjPLf44pSYrQGhs69Yfaxb/q
TUsYTtGuQTx0q3smepuxHPphtCoa6+TYGqENMaP6b0TLQs94gnCCCQPYEjai0L+Q
fDcRcpiUr4Q5/jDjvPMOEGezrfLsGwSq8QiP9ujVHo0Xkt5yNRXy0WokMgLkmOa2
6gPuYekpruyl9ukb98B3jq2nszxb75m5S1kOkG0yaZCEz6n2cqYR4nCTwx8jIBTP
JPnBfxLxQRRPUu19OOE7LQOc+jovlKW91i0ZW0EM5k1usdU0QrbdDf0cc7vV3P7O
kjAEcDuudxoxObxR4NOKHbwvnEMofJaQR1cNIsBi3bbctcPU0LVoIZ5czNQdfmqM
ZwOVlFlZVNVDKgGwoM2uwhimR1zwqJQ0v1uTFAbP0+lh4NBF7SkFbGsEAJIjCoIk
K3xZaApVKEsQuJPmOY2uYqNHj1xKTFBFK805CUJDDOPXPg4hjXIP0oQWH02dDNWN
77Q3ZVGBnMl/8bZP15KcNy5H+AVS04g+pjcFPYAAXWT5jIj0qfhgt2GVMOuwvfYq
SKZ+o5Z6mIfMPDggR2zGF7JHug+eVUuJFPM0gBKE3HkN4Myy00iytthXdcdJjRG9
Gm6/VUey7KsnaygWC2Tj7gcerlB/VRssS4G+XRxtCuYEFgi6TuCf4RH/cZt4Y10x
f9A6wJWLjTiPquQhKOBo3mvKNZoEQH8xtvUPJJJ+an+ZjO6UEONbNLpO0PWOpn4+
RRY8Q4WwDpH+aeL7SBXqqfX52AIszRxMQQwwkJFGzPeiQEk3fDJ6RhIregg5CT+w
6KD1xxm457C0UE98QtrJKfZLdIVMj9X8pqrSnIAyX1jjYk1Mwgqwt+4SCTaBmbbQ
C8PHGSJFgncEtAk4xyUoI207Qo2NMUkp4ntJG6MkfTpkz0dFPvMbaOGD8Q+6dh1F
ZcRS+YQm59e2rYKyGYDaJZDX+EH4XWB+kFX1QLEtLFTS4VYcgWbqix1CHYxPH75b
5xbDNWBQgrg/p1t2ldjUTNNQnyIIpGfVqK2d1mOlC7cKeKCtcENeEE18tfVMKgH2
b/EtALa7WqH3lyymQsB405tHRBepGh95LMxNhwCfvdrI+UkcZzHwdWSZxQ+ijxyt
5V4xVFk4Js1oR3qMY9sC2eGFj/8rjPnAKCYdfAdEV/fww6JfVt23R94vwn4Yedpe
8zP+8NVfJHXiPdEdXXS+q+uxoddhAHKGMIa9OKowS+iNkMjKPMWbm0Uy6lFHdkWe
JxkJb3BBf1sNKfjPCAqkVuXp1csbT7k9TZFwWsO6pwDWvU/vmNBslsaJc9xjp+xa
eXudvyJ/6sWvTI+JI9QItORUTCOA462nFL27hyoaEQMCDd/3JNmnIOETbvowFVQd
VBQ60/JcYNnYC+mJQUfUEixyWYrQXF2aRsn+6FgqwXbE3aw7GYCggE79divU7ct1
Yu5H03e/u1PvGtm1mmIvsrPe5vlMOVeRr3IlhS9Sm3noCVEHtzG87gF1lUZaF4qZ
AnJACVI7op5V+B3CGzKxeJQP23gm51gU0GarLS44xEyiSheEkuuUjTvFkmPf9S9d
3kFjMuHkPb3cDZk77x+u8+ouEyVaWFwJzZxbQ0dXO2RYvAMIPgpEoOsfYATqPd09
4dt66FC98mB2RbV5WHL/MK4og8WBERJiRPf/iOQW9+zu8JyMF8L3uVfSqpgqpoH1
XXzyr/RaH/cecsxhzIc7oQhDLW6ou/DeSa8nko+emrOz8n1Rgk1ftq6pFCki0zjm
HPg0REk+roeXzdN1fVTY2qeVCqFU5Q3Y5Khr6794SwWmDJmLvOmP/amgJTLyoMMW
rLn7Qgd0knuNad/Wcb+XBhiajRuFNWgaYXP8J++nAHwjT8r4+a65eYlEfjghmryF
vMx7K5HYExWlr3z0ucgJph3+xmicvLwcCX6Ywq/zZaWo60PkzU2I0xBjJki2gyjg
qa9PugnqR3M6cdyzNndvho8IEJWrQJ/+whPdtrKRUmAwatCWsId+YWi6C99tvRg9
XCCLEqDPR0aLhfaZksY6Fj+xx6f6BcHaQXQqgfoSA5bI+u7g4pEWzPt+7oKEhKTG
OnHU6e/Kw0ljh6WSvzfLIoWuwLC7zSM9N0d/5l3l6WFKAjWwtkt/Zeb3+9cro9ji
RXu77OW4PXRvlSeVvMFIuD3kgPECD3Q2qyz2to/g1SU2jTVvzEXOIJkIU8cDaBFy
rhNNTHd6YVFCvJPy1q1RTMhuamRGSfG9WQwjtTE5x/YqvwCuckRKEHqJ6XXgbPzQ
PbHWpFqQF2ME24Lo17RDeto2JQtSHY45LhfJ+DztFku1z5Osm2q4EEgjMFF8DtSP
y5aScR0nnlAuZtRQB5t1GL1OHxZvDshXMASnT6vqMh9X4Uk5PvMY5HG860Kl5on8
xnOAxek8yOMWlKsyUKU9oVdC/HiSzCBAF0MMDjqS7hDfqyCjwQjd3ymWH4yWhhNA
edAoPyFWg4whXVj3Le7mQPJAeHKA7gF7N6lbJPKWOTBHO/AhjtWbATMtj59Gz59j
BYyJYuJMqCGyDxDYQP8iVxwdORUOOS9OTzx4/npUF/YRkq896NY+NGDN/Y8g2WJd
a4IkJPZPCnUIgmG+Ot6Bmjpi/95msVGpH2WPLPHt1QQfNvOdJIvsZ+pJheRuGm7Q
4CV/0i8gUlYeVpCepDkovpzW+DGktSzwmjx1sQAiwA17gH8b35y7Xc1+YEfUGYpD
Su/f9ZGqjMF8ZHZmdFLhDTOyKjjbJWTDWPjFG0w4k4JbKP/p8JVa4UEKXrPF3X8E
2GKQJcUgLd8XfII/UM1KlS6Gc6jvm4RAXuscwYpZEk2qHqSDu/IRAial3ngj6SDw
MXaswiz1sYoewomQWJIqkmb2iWDw2vUp4iR+9Avnn0XQ8VvRBrw0HXGJAOSM2Xzy
+bBgJk6EIk5bEuhIPDPhOxQXUPNN5XlDN+rRuP0Et7SHlQdF5h+y+uGKdajKFS1/
YYbTHRxsHO7pmRBzgAkV5vrNFWR6Q+mMHLU8oRFI1JDsDc8MZw1TLVw3rNSa3UcT
CTK0PuQnXAbeMP+k8nXHvxtUzkUnB3pg/jHC4pv2YNeOKGzcno9bAJZv7nIoNtwH
5noupzQtAAcqcx/BmwXThtmcDfLJrjJSN4KpnyGaEho0qVgvZXMaE3yAIK6G6igc
LcaZ40aLyWvw1+I6ZXZ/qHWNp+vWpZSjp0NWer8GT2PLM1yCydZtwy+NSii/BqP0
yPTAIPbZ9EnR1rQQnG73mSGLcoQiUbNmQfyFxgzfy2t/uEanyYzW5tUe+lCOExA7
hwDUovJ1T91PloBV4Gr0yG1kbhUCMt4JAFTrFwoV08aq+kkbNCOml84cblvVLHyv
GNugmW19kLGwltTr45tMywE/QZMyXZr6QbzYvNqsoFgQ8OoySETdkt/07e4m0mdR
p07kPfV/MBGmNbPFrqks1nOCwxwWtEvmrdLP+LhW2nwHska2DAhhNDuIGZpw+1Th
edmdR5JeQNohpz6DEwuP5MSFPmyKdepPQPV0TuU7yAR+Uk7ijno3fNMjyMsRG2BB
kvUHaVR+PtLmxe8zSSrQs1HsYJAhyIHmK708rsWy1vAaybNHvW05Z7TojCSvEOap
mZD0mP5M+0xG9hjASJEf03qkWV2q8Q1PDFJiCw3Xpm/haS4isSU2rX7laIFQ0a+c
55jUwtus3BtE9i/zxDBuuxDSGbvQSicocA30uhKR/rFAY5OjFmV/tnUK8S5f5fDG
p5yDh38ujHUUrYzde/OLhK3RPwyYK9cCAn+Ma37qoCmEyAn+x+W50oXMiEa83mU2
+11UtTUAc4NABVdWPTyzpfpPoAx5JXcyqo7CnNoNOUqc6eUbzVcLbPrqWLh0THmR
DfEYkWiHoHNhpFT5PobIp7BkxlaP40tWehbGu5QlcISvfsdEL9SbrrXndVosFM/e
YV+gEQW99rYlS6oh/G7SWULty+D8wepjco46GLUveNKgFcQfrNl7bdqrf9NFmNzC
dy0QZ5gG8cHyoE4izzxa+q9zcOqFjldJl9ZP6aNs9kpjxWWLMDQdPsQxVm2MUq4V
JRzog2NTx9tEEisVpppPRnEiQz5b85OxurWsHn8mTZ+Ivwpqzrl0Jmrc1wvZpePc
Nqh1q5cSe6MVEAkcZYBoMhQBJ8D+25ejlxR6vStT9gyECDyhdKbgGrWY6NuxFN8M
VXaLiRMRx9lc2d5uKrQItz4JLJU545bw1L012MAu8S1CvZDyKh3SW9UxnIzfePtM
5soeqNW57HK3YzziYac93qQ+wLq5e8CMocKiewyvSo7iXvtlKpqggmtqXkC1rj7d
BXT3MmbS/by0B5zs4z5TaCit/E/7x05T2VDVQQembrg=
//pragma protect end_data_block
//pragma protect digest_block
LFzEWuhWFjhZxpkjiszxoXLpqmU=
//pragma protect end_digest_block
//pragma protect end_protected
`endif
       
