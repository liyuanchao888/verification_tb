
`ifndef GUARD_SVT_AHB_SYSTEM_ENV_SV
`define GUARD_SVT_AHB_SYSTEM_ENV_SV

// =============================================================================
/** This class is the System ENV class which contains all of the elements of an
 * AHB System. The AHB System ENV encapsulates master agents, slave agents,
 * system sequencer, system monitor and the system configuration.
 * 
 * The number of master and slave agents is configured based on the system
 * configuration provided by the user. In the build phase, the System ENV
 * builds the master and slave agents. After the master & slave agents are
 * built, the System ENV configures them using the configuration information
 * available in the system configuration.
 */
class svt_ahb_system_env extends svt_env;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual svt_ahb_if svt_ahb_vif;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AHB System virtual interface */
  svt_ahb_vif vif;

  /* AHB Master components */
  svt_ahb_master_agent master[$];

  /* AHB Slave components */
  svt_ahb_slave_agent slave[$];

  /* AHB System sequencer is a virtual sequencer with references to each master
   * and slave sequencers in the system.
   */
  svt_ahb_system_sequencer sequencer;

  /** AHB System Level Monitor */
  svt_ahb_system_monitor system_monitor;
  
  /** AHB System Level Checker whose checks are called from system_monitor */
  svt_ahb_system_checker system_checker;

  /** AHB System Level Transaction Coverage Callback */
  svt_ahb_system_monitor_def_cov_callback sys_mon_trans_cov_cb;

  /** The AHB Bus component. 
   */
  svt_ahb_bus_env bus;

  
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
/** @cond PRIVATE */
  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_system_configuration cfg_snapshot;

`ifdef SVT_UVM_TECHNOLOGY
  /** Fifo into which transactions from master to BUS are put when system checker is enabled */ 
  uvm_tlm_fifo#(svt_ahb_master_transaction)  ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from master to BUS are put when system checker is enabled 
    * Used by AMBA System Monitor 
    */ 
  uvm_tlm_fifo#(svt_ahb_master_transaction)  amba_ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled */ 
  uvm_tlm_fifo#(svt_ahb_transaction)  ahb_bus_to_slv_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled 
    * Used by AMBA System Monitor */ 
  uvm_tlm_fifo#(svt_ahb_transaction)  amba_ahb_bus_to_slv_transaction_fifo;
`elsif SVT_OVM_TECHNOLOGY
  /** Fifo into which transactions from master to BUS are put when system checker is enabled */ 
  tlm_fifo#(svt_ahb_master_transaction)  ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled */ 
  tlm_fifo#(svt_ahb_transaction)  ahb_bus_to_slv_transaction_fifo;

  /** Fifo into which transactions from master to BUS are put when system checker is enabled 
    * Used by AMBA System Monitor 
    */ 
  tlm_fifo#(svt_ahb_master_transaction)  amba_ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled 
    * Used by AMBA System Monitor 
    */ 
  tlm_fifo#(svt_ahb_transaction)  amba_ahb_bus_to_slv_transaction_fifo;
`endif


  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
 /* External AHB Master components */
  local svt_ahb_master_agent external_ahb_master_agent[int];

  /* External AHB Slave components */
  local svt_ahb_slave_agent external_ahb_slave_agent[int];

  /* External AHB Master component Port Configuraiton */
  local svt_ahb_master_configuration external_master_agent_cfg[int];

  /* External AHB Slave component Port Configuraiton */
  local svt_ahb_slave_configuration external_slave_agent_cfg[int];

  /** Configuration object for this ENV. */
  local svt_ahb_system_configuration cfg;

  /** Address mapper for the AHB system */
  local svt_mem_address_mapper mem_addr_mapper;

  /** MEM System Backdoor class which provides a system level view of the memory map */
  local svt_ahb_mem_system_backdoor mem_system_backdoor;

  /** MEM System Backdoor class which provides the global view of the memory map */
  local svt_ahb_mem_system_backdoor global_mem_system_backdoor;

/** @endcond */

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `svt_xvm_component_utils_begin(svt_ahb_system_env)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE);
  `svt_xvm_component_utils_end

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new ENV instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name = "svt_ahb_system_env", `SVT_XVM(component) parent = null);

  /** Obtains the System Memory Manager system backdoor class for this AHB system */
  extern function svt_ahb_mem_system_backdoor get_mem_system_backdoor();

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the sub-agent components.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif

  /**
  * Report Phase
  * Reports performance statistics
  */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void report_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void report();
`endif


  // ---------------------------------------------------------------------------
  /**
   * Connect Phase:
   * Connects the virtual sequencer to the sub-sequencers
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  // ---------------------------------------------------------------------------
  /**
   * End of elaboration Phase
   * Displays the environment configuration.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void end_of_elaboration_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void end_of_elaboration();
`endif  
  
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the ENV configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

/** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  /**
   * Obtain the address mapper for the AHB System
   */
  extern function svt_mem_address_mapper get_mem_address_mapper();

  /** Obtains the Global System Memory Manager system backdoor class for this AHB system */
  extern function svt_ahb_mem_system_backdoor get_global_mem_system_backdoor();
/** @endcond */

  /**
    * Enables AHB System Env class svt_ahb_system_env to use external master
    * agent which is already created outside svt_ahb_system_env.  User needs to
    * provide external master agent handle and its corresponding master index
    * number. It is important that user creates System Configuration including
    * the port configuration which is supposed to be used by the external
    * master agent.
    * 
    * If system env doesn't find any external master agent for a specific index
    * then it creates one on its own. So, it is important for user to set system
    * configuration with correct number of master agents considering external
    * master agents and set specific master index for which external agent needs
    * to be used. It is allowed to instantiate some master agents within the
    * svt_ahb_system_env, and some master agents externally. User needs to take
    * care of correctly specifying the indices of external master agents to this
    * method.
    *
    * @param index Index of the master agent which is external to the AHB System Env
    *
    * @param mstr Handle of the master agent which is external to the AHB System Env
    *
    * @param mstr_cfg This parameter is not yet supported.
    *
    * Example:  for(int i=0; i<5; i++) ahb_system_env.set_external_master_agent(i,ahb_master_agent[i]);
    *
    */
  extern function void set_external_master_agent(int index, svt_ahb_master_agent mstr, svt_ahb_master_configuration mstr_cfg=null);

  /**
    * Enables AHB System Env class svt_ahb_system_env to use external slave
    * agent which is already created outside svt_ahb_system_env.  User needs to
    * provide external slave agent handle and its corresponding slave index
    * number. It is important that user creates System Configuration including
    * the port configuration which is supposed to be used by the external
    * slave agent.
    * 
    * If system env doesn't find any external slave agent for a specific index
    * then it creates one on its own. So, it is important for user to set system
    * configuration with correct number of slave agents considering external
    * slave agents and set specific slave index for which external agent needs
    * to be used. It is allowed to instantiate some slave agents within the
    * svt_ahb_system_env, and some slave agents externally. User needs to take
    * care of correctly specifying the indices of external slave agents to this
    * method.
    *
    * @param index Index of the slave agent which is external to the AHB System Env
    *
    * @param slv Handle of the slave agent which is external to the AHB System Env
    *
    * @param slv_cfg This parameter is not yet supported.
    *
    * Example:  for(int i=0; i<5; i++) ahb_system_env.set_external_slave_agent(i,ahb_slave_agent[i]);
    */
  extern function void set_external_slave_agent(int index, svt_ahb_slave_agent slv, svt_ahb_slave_configuration slv_cfg=null);

  /** @cond PRIVATE */
  extern function void set_external_master_agent_array(svt_ahb_master_agent mstr[int], svt_ahb_master_configuration mstr_cfg[int]);
  extern function void set_external_slave_agent_array(svt_ahb_slave_agent slv[int], svt_ahb_slave_configuration slv_cfg[int]);
  /** @endcond */

endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ZSL7Nmcr8KEDt/0ddEK/2TODKpAGK1x/0vpBambKAFGIMcNXfl9+z6kVhM5f67nl
60BHksA1dmTM6M3ljgVGyNhQd5p2CKHQhJaY+wjg2kzx/P089+EineJlfp0MJ4YV
dpc8D3SJU2e94nqpn0R+qUD6T3huTyZhHcT5luJEUgM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 361       )
7IJwJksLuzdpJoUv5IRr3oEnHpCQ/a8pQl3OMr3mpLhdYOwKCtTfF5HkvziEdGqa
A2EfP98K70dKMIh7tBOrZCqYyyoGBsdPhP7X+iC6Jcl+E+ANqL9dhtXtUXUTV3vx
naSpfxguuQsy1smUkxL7U/Qb2JEAJJWmQJ9ugZjuPBr32pyLEomHClecXyQJFmEN
9JLPI6mXgWEnaa05iwWWrWda/g21fnIdiHcd+G7fUwPlSeSptDFuRqeeNeS7RZLP
4D3XqHRIwd4YTPrJMwYeyxVeT7V52IbFstnuEncSdlpoG3H1LC5msefYPk8C+hvP
YplGiRauFj1tnmx2Sv10c54/YPXEVNgDcIq7KLzXcm2IC2OZhVgtlDwci30G8LiN
Kjos/18Lx2ftXSW1Ynd46ojYVR3P3gpYHMSBWTBbNFBydaexHoihWSybkiDmOBKZ
7YfMIPzUeUJOxRkbgMpLQNSnGU4ZMb7FdJP0+R1p2fM=
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RUua8D/JFQBteRHo1RT9nuGDpHSCb4BQctfnqDyTkUNYkaRP+RE1aEXWppD3UriI
3b6hyn38fx6QAhRYVgjWUIHWRBLFaHS2R5W6yIJ51oCqYwzER2LhWndwFG6tkEmv
tcAW7FhTNG9CgO8ABhAfJvFx0T3tglrPPXd5FExaG2c=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 20070     )
H9jdBIIjGV9VoZ6uqQfkdypztl5n4r4xlDaONY+QgKNonWtceqpipifokjU5NmGW
2Te7+fmJHAMrksW75RlBYpkfAKolivIvOUnggC2U89KWIPpvou3SNeXK0o9Z8NsJ
KxM9RrIPlVclj0090zM51yxcoBhx4IdZuIRMvqXV2bOoQh9xQEkPw806Oih3ekDP
YPPIlzmWv/3RKsEfym8nkP/anU2weN0GBpPkH+jYWcSDaUR8u3GCJVHn8RaQOS3j
Fz2wBhjFX2RzV2dZPtQeNl+xNwEVZNyAnYPU10N7LqxID6WLQauEfE/cqVUGi+4X
X3vOAIBI+o2rqqf9DgVHlg8IqpugBUOpMm0O6sfaIT8djqw91UxqEUjQGUuSIDuQ
RXrrM1bkgkvZ/EAqQTshcYYTrFdEWk9BfnOirEUBoJn2Jw7Vem6Bu2IXDsw3x/An
Us99OunNxceSoe3mf7AK8vIELDkSNzrX955CH+9z2FJkJ6Mka8eAwRPXBCyHWFpD
yDtl46T0LdiqYcBrULyDW8LQt63ALMGNn1b/sKW3ngO1ln5p0y/ObXQulxIvmA0U
50XZjh4cAm60pEa771rEbum1L4lZE5kwjvQkPDWUUQLFsHhHkdFKjBTSDp8RqsY8
Us7f9oyOGiduIgYUMqVhtP26rUWgfBbRZgDszcpk/Ojr6BtuE+IttjHQcZhHOGBr
iojUTXEZdFwy/KqzG8ZGPxUSNoxmGYF6ilBgqVkLKzninZH7ezJH9u/28DPNCxGa
sA8TUJ9XF9zHKkrvVWBmwGY0pIkxiDTxu62xI4F6g0nHI/yqeyDE4lKfoH/uX5mv
eZpOJVWfW22WUaxc/91TqawT6yMDdO4w3fVg/pnSYhb1CK2zEKD98u0yaC2Xb0XI
q4Nzx5gDVeLE/7hvPBgdzIuiXAfat0g9D2k/dZeqrW0BHhbfYyAGT7spTbsK/LQn
8it0pn+xx/2cfXBygrRGMMYBldn560mq6GiR0FAjEYHEdffpx25O1mpurCcNHuZY
usXEt+B4OBtU2M0HmeKaksKtlaVJpa7QgzHC2JhdnNDo1HJ2tu71mCTKt4R0hTBw
8Qi7sZwJA349zYdFz07aXpGAklVlo3BVYlvwtg2fUszvSMrYxNEh31lgLd3nRcDN
KlGfj+XPN8mKE9rTwGLDolLQmE9+ufAOmWhubqIsc3F4TLCHUNRdC2V6AcvNGj9b
w7ywsBR8uXHTST0At0urdHnUblKKYdLQCrmx00MMPPQru95ZLc2HjjahklQR/nE3
ZKVBoG0rDbSxcLoTbzXj/Bix+YQNmSwqL4NZXN7csS64e8drHGRJ5A0KPmUrA4RI
3rBjukmX4jRuQjdGiPj1wEsKE85SSgzzYiyOZ4a0Kaz3E5NxmeGs/KktEYNy4yS7
m2+0ODC2FFZ+N0cDhNhXRa/axdJG/AdLwKWlK2G0tJkH4pMNoQSqD4M2sfJGk+3r
3wSODnFhqJ1pF9jTINROHdrRbr+9853U4XEvi5Kyc9FU/masvN4Pi+FpOiR90u9F
kfG/8yy3RsjJU1FEQri/RPz6bhYOe2VfLIdCG5Fzmz/h4tvV2J39uuaao05q3re2
H0bp9oLhRy4wMmBysMh6fc7rzaxkJ6A1RDtJqHY+c1QNAPFTXpu+P6L4l5mr5NZY
WRZvVx04TvcPPMURzXvrAqFh9xo7yPccz+PuQkABEgzPgU/9sdr28wF6R36bL16g
IB+xbmLhP8NunZN1AllT5eI45kU+8NaLzuXdGfSme3SaI1PZdDUJ5lwFN7rfFt48
dApYhcwFnDwSjY+zWjIBU+9ebDmw8+M/YO6hSdrId0+TB8QukIk4VzddkPB/SPXV
D40c12MLDSZLxJuA6D+6glX3VQjxRx8NqIKSmOl8mhRxA/R22BCPVJ8PihIHGMOd
cWzzeQah0B0F1X93HdKdlKIuKLeH19k/SCDfeEn5Y6dWdfRxCmSi09cpfJJUUHBJ
ObSlg1dTV3RdPDb1f46St/q8JgClzvjg1FF3/2guHi16NZE/3NbBubPSFIJuuD8C
S4woy42c4yfvuj9lnPAjPgjw4A5jTXVwdjM9d6D2r3TImkMnPBPDFlFN7TXKBe4z
/6RRLbBbwbS63GdKJxlkAZt/D70ykMedrmPpzrJC3D77t2QHLeJIRAjRg9tgTWAb
QQw3UkqPJXYuD6qQSpCAhAn5sUSY6zLbsPTeZIeRybGRhGks+85+nHQXRlHO5E1v
HL2RBTAJ9Mnlj6k5SAHagChUoNXo2AgV9hEL5qogFY5AHwIMNgHqIjy9yK9r4Iq6
WyrK4vm7cfQ8hIVKkEfyQBJCV2PKO73KzA7bGioxt/mWiCvXGHF65bRIC1uwjXYk
CaPr/JeOiRJ43kXLF2zvVAhCX22lPEW1WF7KRGj2CK17ovndBSyz++IbThauOtNk
Ob1lA51EHCb7BI9nt6yFRZvmzvrCyV1d5gRUDhgZgV4UE3a0MuraOcmMdJrT3xjg
qXGWHLuiJP/cYJbxsO366iCO3xYP5xVw1jdeS2rWugfajMlZY0zRilXLyYY6iOpi
Ha+sz8PF9qpcMKPNVaZDuE3ORuQNY620QmmbW8MgxpmeXUQ43Xk4BD7f8ziEumDb
MxynNvBHOFO/TVCQ+uhnB6MaFHIrhJ4u9VzmjV8ToE6Db7IDolbLjH6osUtm3Bck
C+hQ5t0lJgXunYgUtaBx1JjUlgEYbuo4hw8N6P9jYAAC1F9KXJy10Q20Dp9Sx2C0
fyIV4FY1EcVJYBYdhkHXHBfaqIwcEoWl1bVH+JOIAv6r7IcjXd79L/r7sdL1JYfK
cI9mZ49cEXu8P9/Nn9+uwS6r6JAc7qRFyg6RDhAHtaWU9LoTTFP/7WrWR3mtnGKo
ZiPKIK2F2aNmqwXb1SAuUvHZwUvC6KIMQIMIdaWP01jOtLNo8u/zvDPt21yCzUrZ
17h0X1htg5FvUuegzjxUiOQwqHOhAtYLXh8JwqQRxGGVplFtBGYCweULX+yb/R9t
S9G8qu3y1gZJIQg4dMuPmYkohbGpPHOUvYbxMNK7Mlzz0bLlzLJ8z3xZI3CaO803
Lx2ickUo5Upn37JCN7zQm9qqc9jJo82z/eyk3wXyLlBq/hnBwmSRyB/QvXCiEo9l
xF6JS7f8QC5PkIkGTwWT85zwYuRFOblSb70coc8L61yavrR+UjRUBzv3rf5F+x45
26NMHU9zZbAemTG3ejngzCXDPpNgHYVhKb9GId7ARPZ0THJ5ut+gGWZ/AFK6cKiC
4+COvIG+Kuu4TgQnIUEVw4/RZ8fW1uQwHSMiAGA/FIOyEO8emQJCEWKCsnB668kS
PbRC6K4egAHpmgWignm9uskzX0Eexhj40ezDhjaY7Q4QyTZn8uOMKXEzSwJwSdJ0
AygnKRyf4Y2XPiEjDqHhSXBeE9AC7qFqrfZJ+adXP7aIRCIFQM5ycJjSFi9/Maoe
Q+fC7Sz+uIknxgSEZwdm7EzXTG7M/nqevzjRLXscarjAt1amRZ0nYvpX8mnqP7NI
wsKbo5qW2m+F3/xkJkbYsPc3++TDV4eQvVllNzRPDDdI6JeqDMIfBTMyXroflFbk
w05T5yTTIqsI+Qad3o+MZt8M3uSqzfF7c8auNafaYPXzTv1wJPIGvSvgjl2ngAwl
m5fTPpDlU6ffjUURcRxjiwG86AdB6zXGWSnnbQo3NO3VikZC0EfN4IOhSrGA2o7J
v5/Fj8o8fvDFjs/fchDlAygbRQ+N8+0XCZdcKuOcZgRG49U8JSn6yFxiVQqv4uTU
YK0s81eR1LWSFqJRN6PBIL1PoKah05kzs0hwI4KAOxIaXSOFa9TI60GCUBMUjejD
w6dS2sNsT7/wS509ppTOSQL5Xya8IvcQF3kNqoXqJOU7dPmxdFeBSoWD0X5ND81z
8z2mq8JDsd8k/SaLJW0FqpLtjkq5uWOvOOciN+Jbubx0Mj4FO3GvzK3F5Ag81Il+
JaQ331CRinnsQ3/JcAhluq10kxiyKH0UUsHMHAMziBpxKQ66pZL6f2FVnX6mSgpc
gQfMQQ6RuoDECBn7h+VfOgljXIK4zLaRf9azJ8+9gMxBJ+Cc8tWiP4uvABmfoZ56
DrtK1QOXUGdGyc5HXHB3Cf0ETWgKGGUEZ9GFH/Koforymz+vnaXAgO3Nx4L6UY93
UBsLXCfQdoTESvd/bdFuOjXNccuyC/ONe+SX81aZX8mGQlbV2EShQ2BYt2wF8RA9
W3yk4nJoE1m+0O2c7JD32UFcsLwxnG7QhwyJbPRRaVkWI82BxUl4arrz6cXqRHox
LRLjQXcFBWfKvSKxgh/c4k5NqaBJIaMksm+4zICC3+hUnjKMTwb7aeKVXJQzKsS5
fqJl3doh60IBXKNt7KV7QL820BwdtCtleH8vDgzitjOxVBuKi9QN4nJ/9f/LBEbm
xqm7j+F4ZzFVrkOY7RPQBUbuRSrdqHlJoNz9k+icWPX1/0pAmDwj5O7gHkfRbogu
uViMtozx7tK1aarnMreWaJWOL7vHZnUT8cNY/Ecnl8SF8g3Y1ikk2dAOkfZbEbKL
bK6V1PQcVf+rVwpSnh2XM+bxpmCqAPo0Hd6TeLr+EUHN3ymA675YwcuU/j4cIKVW
CFm3bZxKqe7YdeXj90tW2JHm0iyFilkdn32H5j2mceKj1SSuVXoFa2n4tZ3UDFKV
BGlpq051HJq3+oC1eIWvnrNlHAHqILAA812+bpAKQZ1ta5QNcJVhMCHco95WkIOp
YKJsITE/mqwH4HpRQBVkWHkxFjT2YVnmzvmnhUazJCpuWpWcmx9nDxGDjQa+ge57
GL43hF8JTHglEmUj+ZrJWhKYxbaYxhSOrWLtSjsAb7Yx6rLsEi71i3hcO8ENrj8J
dGOeM5poA+kv52qIEraDaUlrJcsgOerWDikGlkQz8hJ5pgE5lcywsKKusDaBr+Fb
M5p8oBeCyqGRslwwpYoni+tKSQoAvglauWwi/jTeYRCG6NLzWz6RrbInxZWYojwq
QUjlaIbQeBIYlSM6/2e3m4apeelpcWhiDdHMLtwWMyCP+NHcDUybkgY+Lz3FQnfj
2347M7eWda6FHhpFFhugcNu3TgMRwVn1GMVF3vbHvL79cMkg7cVBbwlhoJZv3LSt
jUtWadfR3ZJ9mVI5x9D1LIuYObxr23u53nJw3IGQKSgKSS3EOw/pbnE7kT4J1yPA
nmdFeEA8I77AfVJ60ov9VEhz8Imq0+pw+z3kLfaBxN5iOFw/lSlpxQYs60JnyMOt
w6F7MHWHSJs7+FQ1PiRftoxt/RA4ioBoYs0L1OxMt6AAVOYJnbZWeIf0qbcf1K5t
jYR7UUlKtSCKo1w72heP6B1Io8nPRiwidoD7f724zpxViF6gAxDH/cxU1NlSF5Ek
F/O2qaEQPFhiWKzNCjOr5Flr9UOepxkC7JRNLCm+7qPXRZlb9rm7PrIRQacsh2nO
RQiiMlol+H8OC0rfgawzLhocmP9i/HzAOSBl6J7zbEtEknQNAIPUuuEjeIaWztMn
HEZWLqgqDulKe/3jjkrP/cQ0s+PW0SVoS+mhhggd8yKZASO0GNvUCXQc+ZNMwZUw
Xhi95b5prJHhUEtsf+2T7jRxEXaG/tjgjA++avfclE7qwBLYUSKSlr8f0GHRokqJ
wFc82YXM2t8JY7A+vyzufVnY9tO63KwWl05ySTu4n6tTdBY5PncjPh2PeOUaYFiz
8uuvnWr3Gan2A5/+vHxMbJf1P3YZhqwBr5yxyVmTJF1O/HQWKLH5oiYjKA/iTpwo
t95oXPxd1qHDmz3heu2NEHMvMeEcOQJ7HUR/an6ly14sfiKODHbHCZhhp+GdyLHc
YeK7+2a8NufHytPWjsa0M2Q6v2htGObRTAXjrOh/SiS548dDSFT+9R4+ZF3Y8obg
OUK2vxROtEzgJ+4h4ANkZSvwvtWwDSPGVS06VWQmYqglDufPNERrjxw40SXwj5zI
/o1ycFomOH5evHKgbaRo5LlEaXx7LFl6DKXqjaTQ/UcnD/S41I3dS5y6YGAC23kf
r+wNqeqlakJQcoQLTqpHtfAM/L133MMEIapdvaL/ztM7E/BJ8FAwG8pWhy4tjvEM
SzDAvlLwTUmtMur2Oa3oBvV01Xy/yLOpXcV58UodUPS2Yee00C1a5/e4chtUSwKo
PV2E+a6VKMW5D0mK8hrB0oyabSaulzCN+uqRW4h26Z4ZwBdyt65dv896IkNuqzI4
OWwj6Df1svXNGoMLTPxDnedNx7UyCZ3V9xOHe+vkOF39LMABHMqRo3Ig6UPLSJ1t
1wBbd4+UJFCMLsDucohTC4oJjHnv86/b6LUhOd6spxPGVeLBcUG1uWTZsOYtlXN8
L+k0yNx9rf5cmDvBQQc/lrCqRh9Ay28ljukzWh/1K2plx6VajsYTi9RZ8ujgiBU0
w6UzdlcPn8X6H+lv2SihedF06Yeyvo4q4nwI6QKTkEM83bdU5jx2c1m14Wf/4f6p
f5R2qvxzL1UOSro0ll/iIUGDrXFeJ1CNB6Nw70YLEdu54eIxNEaMhL+CTeq7iDuA
t4/sCPJEtSd8K31dakN6c1fQgI1qjJWW3E2bOOWdtiqqErhPCxdyfCyNGiMGS1xt
K6e2j3/18w4d83Ds1FeiqbFGXQtr+zS2GddjxBWK+SOFe4PIaDdgZHUyf0E4Xhg1
CttNHH2Bjmmf8OJ83pFZm0F231nmJYkQ/nIuLEnbD2Id2l1gGeskH9hm58cdx/lK
Qb9HVZxLK2/t6zYOG1QbATpPHjdENKEGgTAOmr9SowLZtYi6MljurA92RL1k05JO
uk1k2byWbl3MBEuwo8u5NPy2zLjYhfxKJiGZC5FDqk3WAZrH8Hd2tn7w1+PRaCVm
0ItIljL5n6RXFxHOHtxw9sxHH9VujF8Whtm4ZxvLjxqITlv4tWnNiMbu83kgHevf
mRhJ+/nNizCvbmq9foBfXfQPvH2owS4OEKs5SO1eZxfgH4W2YuyrySHjeyXM1lti
ZGtaDBAHiyOVtaqT5uFSToTDFXz/ayUAa5ZqJFhSjjQOATfVi3I+jrYpUwakL7Xp
MtDRsY1uL90TtNkgNzmpeo8gTHeDe6q9t8v+AHVTpfxKGLXbWQquxrsVkmqZat66
UPX3zJzNI5EAEAIEZ1x86iM45quPmaNhuyL4XYTzOtIYty5asIiRk9nB8h1zqhF0
6OVw0kvPWxlyZKZayF9KvoziXdNLmgJk2vjwh8WTr6ZFfgV/FA8iREzW5SH5I5ci
t2jgjIedtENmoab712YiQ4M62U2RlgmTgyqUPOl9xP9uZ1KJ2VCtja8R23uY3UtT
rWxdB4EYtMRKMuV4yyMN32MjaQ6Y2s8btscuUpmu+N6aA9cuylYKWtd803qauH7v
hdPfnjh0xZhuICihaOfrn4RlJoxm3L7DBeti8ystAGdwuoiN9lovdhStjkjmqEs5
Zeq87j30K6TFsxQcqRPvKXXh5TVPjDhVe5Pv0bIgCB64g7eiVnAwnBcPjhKD+mix
FnZ8NkD6MyvSnNq1qHZTMnv9FOaU0ZidbLCWDrxHgDrEuDVpbS7PPmVpxvEhzWym
ymtDybnbCt6+flpS4gl8PrJVvKNvL+h48rEbsbdYMdyDXIHjObMafpMZCO0QWrCH
qe27FmjAWq6cLjHH0rdz/Nxy+GyNfdQ2LAJQkte0RHhEUuskpI+W7nLGNUJUzihe
17EJuheKiWkihFBRWmj3qlCHC1VxoFgDuMiGfoOMihqoPFkiN3Jmn0UzOZTh9HXz
D9JVlwER5ukL3HCejnvT+VYsUvKLb02a6DA69Wt/RCGh5N5moLLBR1fpHrfg1vCv
q+XhwaVjDcmUeGEbql/t8a9rVGcy/lOWRZ0S/dh0mZ7tOtGVE2ZQ7oFCWXeqMEya
J0AZb8D8ugRNwfPd8Ni69AO7gd258InKptmr4G7X0KFml57T4X21WJACVOtMkEix
eXkxclpjyYutFPlzOE17nORlJAizBOLoptXWjBshhKbM9996Ts1S0z2yU7SP+7Oy
F2S2n7pkpc4WpLubNu0jgwephH53NlAxfFqpa8frFjOBkR0gXYhjGOeVSnIYb0/9
bK7Z5EwER0zXOp901G/ObA4ABbrAraNvleRC/XcLlItW6flnNYc79uHKSaCqtuL0
fOqoLWXqE8crgFxzbnDrVLR2QeUi1tBY0h4txpyAmN7jEx+uqxz/9/fHjjLzJuuK
RMCOwSo3G5Ibc4rwWxrFIULWLVQOz8jb458yHEbN+X8O9UxezFfLQL87XKT35/QB
bC0XhcdZuVduydYlh6FAHp+Dkgs43bt+33Gn4Of7ncvvmuZskwf0OEd+2E9nnP3R
sLz+AqR6YCXdoyGWn5c4+grOWaIy8NW7nNnky9DhCajlQ489DQF3YAq4GW5s83eq
2j7nhkZ3b36F6TKmih8oxbNiQ+3MFnWlTDgl9Gs4i9kcDvi4avkm3VlaiuGgsKFC
FRKRnmXa35u4ZxF8EZJdy/xEbPlfn0WbC3bd4gtXUjziM/ytH8ytSU2enNcRlTcQ
n5ReSyJ9/au6Sa9XrJ7cwdfFQMQYq4aayoX+UjiY0CN1W6V9H6ZBIOebFt7MHOcL
EzPFFGI/0hw5eSAOyYRZC4eaFinPDDYVXdYC02QbA80JTJQRxqtniHdG9JNGqIh6
4eVHeNh3ZVW1LOwvjulnPMAamUDalXAIQv4AULjGkNGSjqJq1VrGZHUSQ+N1ExEw
GR7fN8ecBeB3uXkN0mHAQhWArlUAPtHb6DvlLWlPjxrB8x2ZO1tHTS/k0860HmOu
SGU0nWYB1Mpwz8rN0hu7HoXiDa4R+ekh9RPfFPwL3SKh9dHDO1anlZ4Bh+d8Bq4l
GstH9FN1wJ9UuUbZLVZvADxoPwhEGSFt3iDjmkf53Urg4xEFZ0C9rhaC5PF9fykE
jI8s3qt9UXcVsqpIJlWxLwSBKePFL6f58/3j4+cK/S8Dmq0GCOOLrkJc7co6FIvN
oTGOghLAUKKH7uqJfKWQTu+bioiMPXWbrFAHnC1lDw5JY1D4HVtD8zMj4/CnNgvF
q/ibYZK9PsYiAKgF+aNHddhDAdqAY7RccNhICSTGTPhd23JIAta/YjRORESgK1Ve
XD1RbK2ALFOMY3FAQDwKI9M60jHguYwbrORt9EhHTFiZ/RzONUAn+z6JJ+XosOWo
HRRmbQMeSd84oJ9ubWljIy4/97ce8ac8OeE0kBasjT3TCRYfeLzLGdzt7PXAHhus
RAKcupiyQXAigSFGAVVzQcEpAzDw8LcmsasKBe24K4C4R8sgel9oP9/mP7pZH5oX
m3DWJO3sL7lb8GobnPoUUbEkuJf7v9pveehVGRXC3H0mMe9LNpjJAoPRxdDzF6Jw
TJuIGRCFOZ6ZezEXsoScF7RYswOs6ItqLv0raEjSwQPeDyPeM2Xutv7SZAPO2Iy2
il7B1+yRd8DDlbXXOpVIMvFLEgRkSumJp41ZLiOv5dg2XUZxqsniV88QIrCU+Msi
yHJHbVuV97OtrhnsHn1jLVPqKkHNEofR0hy4UurLwlGNT0P9U07dRm5jsCDPwwVx
nOGXV41HWKr0kGjFq/KdzeUYKbo8V3tQd/ZfnYsYVTB0dpmTP/vwZtT0mGW0IexH
5UBtu5HmMU1caYPPL3pTA59M34o8u9xrgY48pWOLz2a1QUdDgIR8Yi0lLJqmuA2N
iVdKaltDIuqCqydHtTQ4oavL7Y7gZZw4YkWNSmgLhstm/cG2z5wzCAUGLpzOduJA
rJa+S+T8bXFZGlO+7c7S4yX8nbrmN0IGGNSA4zaB59CXL0nnxKYd5GwaiZB54h5m
PV7/+qvhpQ5lI8ILHqk8glRhe+dGqImUTcXZ+RtsA2qtchA9OFeHoKtGUAGedSFi
NpgPWhf+QT7wHMWc521hmZXT8AMTngcN/l9XWFuT0X7CKbpUvzT7bM/8owQ0j8XO
VRGI7e1+mwVpdp0IlbsGcoswbyNfyFUmZObGHRv6CIpvhke2xziLNLmmMIkMhOca
T6sS82dTyqRqFlaFGOxO7uYRG4wrle4yuXgQgUB7cItreLWTOQmjTj7mDBYyY4RQ
Bx8Y713/QQyuG8gJEEH5VVVBm6f6035SBRracgUQ6v2v/FFjeES3DLU1fvoo1Yh/
kDrpZ35JxX4K4rWJ93Iz5hg9sDf3KwWVGYt3fXMnjZOO3q3l0w1MJ2012SPWHffh
mE33T1BZHDFn71lgXgqzBcDs04KxvM4SvbppDBxwAvoOKVftwHrUBNwMPDRYBbUE
kETBU2FDrnJazp4BAzGIpe7vvw44Ow22i2+7/3JLy35ihceMfctTl1ARPfL2GGc/
9U9+NMsNx5I8lgT/wp6E0CZBkJC0G3BPgdRuRDLoDq1roShXGCb2bwrY8U77m93a
0+wuWxpYOg8kk+Cb7bbGefBIkXfl+mVLlu6CrnfqS1j48meHNEqUsjF4s8Yele9l
MaxO+oFMLMw/NcYNMXfvrjmN1/+AHx36fMB1LuC4tkxyEre3igrfWIVgt3tuDSuJ
mSVdObIti7TWeLH9NujSQ4VFOZ0P+3xAy8rjqFIO7YRPJYSwRS2d2JVfDQufMd3H
53Lg/iL9/7TVhixgp8MXVPGhUJouQZLFurGsqnvjLHOPHZqL2BA7wVG2sqG33VAQ
5/NDVmp6Q8rN35XzaFkZqHAWaJFh8Wo1lUR9gMcHUO1xx2q3J8yGFilARA6a4lJx
LXi57ne09S8pozMi7fqu8SYDcQk2PoArZFF0jDt8yDNB5tRWl7tTY6QLZEU+VxPg
ojBowtEqVqKgghXEYBd4A98BIraYpQpLdCwImbNaRWHvGzKauz6OOKT1kVwZjvmb
vB1tIUkCXgYt+RemlzlbtvKX5XBwrhuAYz0ZPfv7dreo1XBFiPl0NESfcJoha5wf
1dYW0RvVSLnDsH9O/5+AQ/ZhPLCCcBveMkZBkLPPPbR+P1fZPINdTe7Uu70tXv3h
+TLbt6iejtVq96FpNNpklc+o34MlxH0i9wuJnzWDAnyLrh8Agg9IuUl+HOzuMcGQ
CB65ffHawp1K9yRSFWGxPqVdY8bE9N4m/GsKuEPgWpDKXuG+Z8eUV2Z7di6rBMuf
jt+rYIWaMYnFq8CnCb4S2WTOaJkHeOuw76H12vAU+psv/zoYk0kNMrdMfoDLiXeS
RhB9hvySMhuboy+h3YHXnFxNuYqaDM2mhA2eThLGrwu66kRGUqVM+rDWKEH/8P6C
E+uts4w22m7fom2yM+A3FqPj/sVC9AnyA4TbTJao8ntTLCaijpXJr9tRKfBZxM/z
c2r3DlKLKUDpzWtILk7d2pzEf8rJbe15HN4I8WCNQySMQnY+fWun5uz4sknVPQe8
5yDi0ezmDGpmnlEjJ2IMIZ5dxcpGy08VXrFAmTnNd2TFQ/zyWYAAo5Ff4BsKVAZq
d5BNeCIQHaQo1RozEHhI5QpZ8TkGh67wYZ3NVbkfzkMTZFpsfnd+IPdx/M9CCQOx
LfzUWwp46l4BAIRrqE2TP1mrLkKn9wBUrL9URIFUAtuYi/EzBs57bDDrZbuHZqgf
2oX6tOEGc9yDS7csfqsLIoUHeVa9QoY1oVp8vOLvWXEi8/voo+Yf7qbKCCLhTlk/
3BTgw5WjimX14TbKOls4uF6A3GbnKgOZsjDdB7eC4Fr+Bv4l3JuUt+S23E4cACsm
4QNf8rr1UFRQnWLAvaJQxw07B5/cgJNdfGkjPrRRt5qX/IpUjzdjQA7ruCPU7iMU
0ZBE+M5Ag9+CBdwFd00cXlfyoXD3p5vNu3wYEMoXu1dKRLgpF0FCFxKzqVbyf4k/
K9q9FOYsImSsdThms12JkWm0Eatyy3TtGX4tXtiZUAWuQDnDevqfWQgTBDJ346to
IeRm6Hwe1TOpPz6cMMteUhBgUL5pFF02Eha92BJSbLPtBus7rC0ayp/ODQ7zc3GD
5eonx1FIrbgJC1Vr4TSuWpJGBl7o1m3RPuKxzbtzepFHZt2iQImxYC/RYAVkdWV5
rLIfQ9y7mNlW3I0XYONghAkZxlpW5mqgCEKU/EvdmbOGFUtVFdOymc4HKuZfuvuG
roKba5Z6DgFBxENgEap8+ScDTBJmtg3DnTOzw4V/+Jfp14hUVuSF2/YyRzvXDYa/
0sHudjXKjBkjiCJhNw2LR3ElwPgx4PdzgzUojihF++qWGWKy8gqM5ocgojOXNokx
8KC/TeQIKpesE4PnDdkwn2WP0U4np+IlS+IgOkWvcs+BlHNgQBQ2dGMEFyljI+iX
hsvWv2J49SnLjhBq4PqM1Kf6XUGouLttJWGoeTBLw6o5hXEU+qcQ8LwrczPRREAF
qYhCyubO9ETyNAmfXMXZmddsFv9MDJBf6rlwH1ieXNK1PeLW63fJRJq2ICXxKicM
AVeTyUb2c6dju9Rlo4u6l5BQntwHpJnXxI7MnUrPSTwJETiRaKpTcuM6Tz/e9UHb
JIJ6D40NOzBQ4KDq/defs1ubhloVBHuexiCXrE0o4zEjC0fzYPpawRQl/Sobfszi
u6q3lS2spbWTYDK1GW0GKjKCbHDv9J6TbagXjnJxWBnCPkCwmTqY5KcIhD46NQWw
HiLzoZdkOsBhdSgJW4pZbY6043SPuY8G80cEglyWiD/RzGwyywIvo/YYZQXDaDFO
SIAZkBMwKvodWRsGUErXCTqOPVoC1koz1dW/9Tk1uZZlY8g2ekZfLhTKb9D+p+OI
y+4yjtOXYG+iRO5jmumk/a8knFZf5BjIUNtO0S6uOvYXuo2RT55JP4Rsayj2oOd6
xpOmHwENqMGjeucshmdGDlX4cpaQJxbqFhJk/Bb8aSyxPuw4XOZwYYUiRtAqslGV
voOoSbZiSFmrkVmNd1G+WbSW8pEUaqlX2j/yT+JOA1OKdzyv6Otj3lodaLhRSVva
AER+Hz9ctO5fSxXCbGDSALijvmsysPCwZW9+6mZFUOryj6/uqT7kjWvmnleLGLMM
u457L1tZ18E9XzTfvevrHclke4PVBtPlIn33qFdCMPeY8sXUzxkdDJPl7kR1ctNb
4M65CThJTEsaaIAQJ78/93UGj87sQHn2/p2DFAGwG5tkbCLY82XoF1+01vHTPkC1
/ZEoDYvTRhCIITmH1klKs1FdEpc+9NQT5zi15MuZGWJbastmSciF9of8GCTRYzIe
IeXPah5o66ORavTIyd8zYIHm27JzVS2I053snBvLVIApfV2PxR05nF2Imfwwb4WM
TN8gMYkyJ5iAWSmxJKUGRTxdHQzwMdiW2HyqyvLcjhcDmnuXLsrannte+2UHTfZ+
dtgvO4vnbCViy9JEyw1Z1k3+HHzWKDtYn3vFJy+dnBq+LZz8KlaFJudi9vPN7vze
BL9rBkhsWae3pEGE+jbckv8yrOodTunrbo8uTEB9ZxsttE72TegcntTwWUwgLsN6
aH2iJgK3iSE+LTI1en4BfFI+Ew3DwPM8yg24eEJPJ+fnqmbtiCf17rzf2i0UFNce
Zr9rthPk+38egDgBuLQY5ccxEaOQLs3rGrpy7gldm7P7iykooP9Zy8mEJkTKdldC
2j2pNi8YtwZ3hRu07DBIVjTCrFuzL6aWdT6AQtftQ102DmT0tK4WsreU+anNjqz8
LN5Gp+fzRm7sVje7XSqjQtP4D0cDfwSVtDqx+SAFk3ujJ1VS1nokaazmM6pJu7L6
nF5xIK6zictOqQYYIUqzS6toK3Ao7wzukAcViLYOGOT4/qd11uHmau3Nt6RaIXFk
SplZw+nMM12UyqKZWkyP/uh+xoEDc5jdCjR7PcT8PzVnk6vJf0LCEH7gfcCkY67n
SCuub57jgD2PAMNAKID4af0r0H14aqAuP6D99NbR52NPKdpdP3e1Jlkm8xUS+irk
Rv5V5zYjV30Teb6OQkMlHQ6M7N1As/vwtDGHt+tgeHdHjCs908hVo9G5iNHYCPXL
SYydviUnXT2Z8HDeNZVCYCfjuEv6PnY1T2kkQfqER5/AWZ0l4ElZ7oR1mEKxC5bp
QPpb+rsA3ykmRu9oEZE/vmDPYHUSDtXrXIdq8nTXj9lIDGnPyvkZapl/zL6OcYDY
spWWKGvG9u1Yv6DlWP1RvxANJWaeD0nWrkwwaDbNFiuPmpDdDNpznRA2jE2Ay4HT
MNHc3RXnkfO3o5IqWf45CfOMdhpBkmoKYshVRg3sG4MyEf6j/6duHtuSTqoT4Uku
mY7+XJbqU+r6Xv+xYsaIOexDKM/dLEuMqR9yNWybIvHnF4JLTAuniL1ZDTHQeWNJ
mbI6x6dFbaWsCFQXgquNQ3zSEEApd19I6xkFR9GRebq7YpOmebXj2AcFrSif92aD
3XzTnRpgwK2JzIr5gbld0XRNr/7EfwyFIC4x70x5Yfqu5ILOVKd6Fi+ySuGB+bEb
eoV9HXbI4iJfTGBGjhv00E3gEFnWsWZwA1eTWo9hZZkIMFfKAwB3EI6vStLhbzzT
IGqPFYCGL8g2haob3xKg5jDjiHUw0JNU0Ulm3E1a/Sd3R8Hp7EGPwgtb4usToLDT
1jcLbrDGdKAYy5P481vWkPullz3HXY7j162j5a3F2kXjurQwP3XyZlUqfbYJl2/6
uoEjgZntEvVJ/ClABq9gYxUt04mt1x2zPZuKOV8WbM3qdmm8tMwonwKNw+YwBg4q
qgY6W48Ux28HZfo05y8qGu9yeJGWXbljngZ6z/GwwbOqKnR6nAlFz2VqPU0rQ2zx
SDCadGWJZGv9M+DYXjfNZE1KzbVbwL3Lsgli20pV9hhccGrdIb28GsCuy1cEHl76
pKMNdu+EqeTbnPGJ5J1hpZpff1ffbomYqq72cYqk4Kcf0j4TSKDl3mrvs99RAz9s
Kk7JR5aM/5qkNm5WX6GN81yNwIwv09OqdCcQ7clrPN2ieEI7zK6HtFUYlJ0ub6FZ
IdnMDJy5kRaLkrr8PGMW76wPqV92Vn7mI3azc7gSKba/YQvNUksDYFRDKXADkpMv
4BRKLg5PQtG8j8s/t/DaP39jXlB2pJ1QHKxFsjORHqdDd6HL5Mq9S+co3LrAuc1w
V2bu2bFPs6FvtaPFDWc9tgczxNJ1coQSGVVh3ASiQpPjwoiQ0puArLMjTFfQVQjq
mK9RehHGZfXFXXd6e4hMlCAM5bMSb0jMuxOMLFfD7pbUbJBqXvsHYiWCf30MpCl+
u5Nfc+Az2pEtAQ4hjwIFLhUHmSWRBgDFKbo7rLTje4Vxa563EMputq3l8QCkZWr/
XrQztYJO5Z7PZWCWjy6rJu+UUWwMZ2S4O8+L2L7nuNmr13iVinlFDZ4oDWeiOs6l
6QnTwPOvy7KMypgHokZznlhA3MnIKUpKmhEhPwUqwJve1M9LsLvyFAkToPaQ61XD
zI34P0kxXfWGP6bhlgsjf/IfbTnOhByWHow76N5YzUkknm+WTekRsYsQMInWAjxj
tU5BY4JVVfhGUA3yGJYrktNX1J7VKSlYFr25aDx8o3VmACUb6qG2d/XL7/rYVx9v
eR+rU8LSrsAsJL8VF5pugpuAZTqaBLEY3JR5x6kQB3Ar42gPfoGAJi4ze4ZufDAL
8xBlwsjuVXZhVz6ZzQbQkvdi3uD4ZxVn2uuOcr+onaZeWuxLG6GJBGUnhLg8igAo
/BTuSxPstueBn9NzsVIYsHpfxPf9NYcc6HrblxFoeeO+d5vXw87MGSXPcwPhELX9
Kc3GEDn9UQ8A+dwWP87TlwoSqN96bcjHGvZ54VrsMN3kOgOwEnNZnb6YvAHjGLf0
EEGvXAvWrHcLOtNy4ZaSbvPT5TI119TcpcX5TdZj8azi6lli0LMbJpaiBs+DkeUP
reECIVHst+YQsqWDZ8SCow9weKi6Y5H/Lv8tNYUUw3OLDJz9vXggjNOoQjml22yK
4JkjRLL7EEVEQy/1tWI+GmLhXxlG+Gg9SQyFPEZZohCQbS/Ix2NqG+nENS8DM1uL
jIrz03S5uLVnr8ovQZLuy0qt/M40G7gCyHcjK4rU2OYBUJ+NSD8mLYYu+NC8JdlI
anZUfHMt6kDDA5qVXpQKVvU71FEyw3TWOkJPA1/ddDLjiE1fxQmOtIF3D/z0pKR1
nRUuEQUbGLlYTbsHc5QERJfXY1U40eve/B+wLG+Tvr2t7pWDrwZbuE3XJzm65+bu
7BNvmHQ59T2YaCsNTvFmcb1ciIH+v/afy5HMsrICZGl0jE+ikLHklj4HqwhroPwI
kjRZPjWs2/zn0HmIwOrvZKyUI9BXx3CHhYLBviMprk71JA8hfF27c8V4hFxWz6Re
ze3I0Z87DCorMNYAjtkZGhoyhwNtfycUBSASqXuUIA2dFUqrx9t4pjnArqFA0DSj
2Qw7Y2ufhRGvQXhHrrPGrn7DdI8X5bnFURWxVo2Oy05rAvh3C11J8yTyuiwnzhT3
y/t/Z5Ne4hCIJCGMLYvewSXbL32H8EOCndrtIQWRGp5l+XKWHcTWg/d3AGFPUjy0
KilvAKMnxVVsOFqxKGjP2FAFpuQT3FzYNqraS5XIwdc2dTZAjwrstOOANVLePOBo
OrxjDbD0zACP2MY5OO11K/MbmLfU/WCjF16shZ6yng4axhN6IawXFVbrYn9rQ8Fn
ArrnzgM9XubDCdYRqtfDp9CykA8PcLaC4huukgsB6H6pFRaR5JOjI6t64kjL0o1C
W0ZZ9qwcksrCGOmUSriuMnpbr4rsw6sylbFSODpDXPgWnk49QxFbp2CciKzuCVG+
VfdJMSNPa5CNuAG3X6Sr6tf66irEmEKXt/SCGaF5y7lrjk7jEAHLjNILjWAX+NHX
e6IZr0opcNOwwhnUCIeTJHv4tVIWI3DbmALUfvPo4s7yVLJMM65efDRxKg7hkgyS
KjnYyijMFq4d1FHzFO8M08zvxnP22zxKh6O+lq9xhf8RLRn0kntQjHbcaGOTTNMr
Sk+lzoiEPRY1E83KWVUKbhE+l5Y+zDVikj2GliVq1/Ke9m9B8TwS1aCS9nqoFCnu
azWCoAAQ/UlKZXbmB7FEmLxYfAEsy6OhBbKo5GT3jXFQdwlKmdkCMFDAs5k+6HKi
Clj0LvIeyJUV404qFKGeOWmAmsNfqv1DLgrKz7LLM87m1wcsYl0mh6L2s5oUZs76
dIeEval0EykdaA3rVqcTAJ2ubbARbJz09i1NzO2LnEjaVuGj+Vk0rIwYSb6QZe3M
hArqC5S0baMAwJUhDxHcZy7WFjDpvQ8tpM2//pvvRZrUEJmKsI5e9QT2CaelzBf5
EXyl515FfrqoS9p1h6Gq3brMhXQaqixOgcyrnDY3/hLkzkoVdhuU0VHuATda61oT
37+tDQH1+5U50Pd5JiYKhpuT7dRYbbyXewKB/FhRZWSwY3Jw6ik/RzATENURGtdE
u0hH0uk0mMB3vbUsJh++aItEkjQ2a0ZascuV7aGbn+pZxsvODVUvUCyT3EaBjgZZ
F2+HdeWFNAjFJ/1AX7rpojvUF5tqvXgbw6JE7jjchkFW1hGosbDf5UmE6lvxBLb6
ayK7ZaX/I9IEZRBDPuBrdf0IiL1Rt8l8ZHSk85yZ4pFAD94emNxBWnSUIqUAxZBK
ju6gDcUjnqC1Ve0ElT5uh0P3CE85QPRZ8qlyW/70esLoPqPaC49X5Ni4GDxQpVlM
PgOFiHA4h1jaWsIhy+Dqg/4BZLixXaUKpqS64T2+UrNI2FrWUH+5Zsw6Si1548AG
foLMF2VCk1d/eh5nblfndFGoWKSe0PfBj68FNBg9LDKvJsOkxoHDq99bx/bxMgcB
386G+JuoaKgZU+F/DX15WOlqJH+i2caHauIc/RPovGPv988DxRp65yAyWoXrqp24
acmOPfKECZrPF19Ug64NITP8xcwIS01HZpwuxlHvv9ZdvM8RE0y3ZylOw0qudGg7
2AGCP+WOhj800pZN0cc+3JDoPPgUH/gQGsQJZuxeUaLOzkI097xAOQqgDHDFiuBV
WtADOUIcWu5pFVJvyQtUxg3qrdxmEcXHf/X8USGTBdoLeDio4uWUN6g1BikgygUU
pDXhGY5aHvJFkjEL4Rtkk0WJZ+ANd4z83qa96OZtRNLemjchSjz382QiKYVoswge
MQeJvL+DND05N6Yb8YTL5z+OzteeLTKDjcJmSMRTX6pCfgpOaSgCW626gFpE1siB
plQ2knQr6ixpQlqtpuaHo96+drviR513MwlzxoqwpIdVd1o5Lb4ap1t4V52NORm6
iWgJki/6exXz+atWJ3tH6Th4dUyp2kjNfF1DY0SuEUycIQZhxjB4KRryWjpUAtDy
55TjdKSuhC1OC4tfekhHVnofXgL1BotSFIi+u5+DwXYHXqNBvpnB/w92QKPbYi87
QMaIW/HPtRaOLYjR30CCkFBzFJOCSQO0goVFRUOLV/KeFwoZeLwRC4f5YnUoE1Hd
uY8kD5wjE8g+BxheU96VG4qoieSdA3o5zMCl+CDQ++rUQ62UtBuaTEw5afNGDn3s
ItPM/OWcewLBHbc38j6jBX8Dz2kYtDV6sCONc/9Xai//3quJqV1p883Uwe+9BbG/
PAnTQ5VvrfTRAaC4L1oAWvD3amWitd7P+Ri5ukRqdtjr5kNfLrYVKfAtpCKk/D9S
RVPY1jYnjrWhMqKrb16JMjlFyH9IfuFy2hPZchPguozb9VVRxIxqCNUgFpqhLObY
5UYgQkGeBg38fgqzIGrcKKTlaouRHZ6pRA03nk7lPhn50ZhiHFW5FpcSzaPuPLnO
GI0lx6d2+AjsKP8GSYf0RMSu3vniQWp0//deh/bsbIotXGCvxsiMZ/7FEVr6LIKX
z2TrkxHklUzeUbQ0oP6YmSkQ9mQE9rD3ghl27DJfDen0aWFxD1Qg0O+sZTNCGdp0
Fgr3NCnwEljPrzUrNvfF3BH2y0un+6aK7/t/GyLTuG/oBnHWumFhhqtuTlHADiyj
hmdN+rC4hpiGxIvLajWHvvGOP38yGweoN0QnqQO0vC9xVZiF8NKKzwrUt58vMpgi
nNkMwX3jeQlEMS8CJ4iLrQFpbcLK3O4QOsI4bbImMAvu9h2OEwEBUXduYZ2G9rvr
HPf9TBXLJsySwoqkg1CQR8kWzEhl6QqIIBZ8JlDm2304k6q0IFFbH4wYUUF6mIEm
GPJNiuEHY1DrAKNVLusduYYuKQ1lLrkZ6Cu/5w6oE4Dxvv4J+Zlk9kdHCDq8Rh5M
eeB5aAQskpETeqZ+n3Dcah98unbcOeb/cMpSwsAygvgeFz+D8AD755k4Fc8PrjPt
btayIGuhXmSqlEqBntyu4T6FxfOHIAF7Sz1ThFpkd7IpRkPWoHt8BrJWqpab7OPg
z3FdnjqaxOn95qi3ishF2pSGuLrtT3ksI2oMvFlsPZv+3oM+O4h8p8jFM8x+PVNu
xdULMvvrma9LpjVJTq9bEkna3wJdnGiEiHr7Jo/1WZ3X82lXtPNDwgvaAXlJVzkE
tJqxPZk1REJNJ/2hkBWXCHsjT57YThJxggkOAADbI4ccMKBGILQUZdgPrfPBoyql
EipphXtDgrg8i8xslABfHis50QGW8nwToIHDKJ/HUzPSUuCTuV2SEH/jowN0nxCf
mkw4O9NPucTtbqfSYPgmwsHdPyU1rU8usGbSb6iKNtN8BGtITT2VP6HggtFZQNCl
xMk09O1RqvPYBQWED72Hsm14W+mmvHVYAbU9o3Mqc1SyuR9ZCdjv2k+rP3pqv7Jt
1Kkp32GJD57i3mekMyhMoSuXTGcpVBX/A2LrZGWlaSfhtW2ZLSL5E8mWd1uvtYKF
sgrAeXjmWj+dEtzKLkChQCd9i+jekREVT43hVNEOxEkDX3WY2Yk7rbVRdGXWQGwg
/NB2Se79L2UKf3zJdlcdvUcqD2P6T2ghjDEtHHpBZLhElUHBCJXDaNV/u/5yxPjd
79nVzE1VDPCDYwjIgYFFxU+9FUADmOlXvm7ramW9g8jEhZEPXb10eT1RQY+1SM40
OzdesUxP9zmjzjEhWwGIoAd64+cuXh4WceMZhG6B27ZOoZy6MHZNBvDDpQrFfk+A
hLhg+23J55hlmKpOGD6yaYmpskAMN1iiIuE7HrK+S7umIwaEwlO+xIKQiJggjuWy
8EFVajzJy9OarqYkfu1WiZQLrHDt6o+xqwkh8WDNLBDXsD7LLafpOvvUHW1tDB3i
eTryoPQHHjrp2w66ntt/sTwzex/t2hQXjfO08Ba/mTyresegWQvQX6lybx+6y12x
Esj8s/oZHflXe1VVf0uKO9CYspZ4XbNtk0un/EAsNyXYRAQTGnKXpZYufRDpBHme
IHnuz1xPZQbl+RLxTO2qoMJbdKtXxzjSE/wnZTnblPNpEsCRabcVFqZWulilQrnJ
nf0JFpcmPZP1wAWbfQNZ3sjH6kH6fHUzy5UpbRP+IW6IQJQlewJRnZWQ9QKYkIg+
YJLV5NKx5FmUo1agmds5OmYb16tvoEMxSOK7x2+HOJCFp6IGhgRgdXrumcCaKydp
apw0xbjjWrgY7L0WVBldXl5NBMhmw60e3Pc3744G8vJ4Ul5bmI6RbQWGvhejgftl
k/09KJb+M88DgJtFoSBEPXMCb67833L1tDdnmNqjLp3S/mZOVRrbyu9PrUIJhjTL
QO+aG4P7iyEKdVDhY5Il01xXBGKcMizHUBYB8hwS8dIhK+pAqRndhAVqifN7qX9a
41Sna5g9LGmO0gI/+gXAsz796IBmhOhddS9TCOY5GqJ2J00ca1/fo6o3+aFJLsNr
g4e7cg/6newPCG6R3VuTqMstYKCR0qNKGi97+STiAciUX0m6QIrh530ueKS4L4FC
0cfCwKvMQ2hArVyJxTfnV28E1gM8ozw/Lb3+UdKOAh3xR2rXOlkh6msDv3arXD8+
lldVdfH5t2sj4EaM2Buo3odE6YxyrQymrEuu7QkyIfPzRt1PSSvyqdml0Ufg+1rA
0Guu6NZ08AiA8QD0fFHrcbve8P16z0R7YaUwbNgjzyovNiV6gwveAL7PdMuim9S+
cfEezinHG5aXa5Ra7iIq9DIRVd/ks/S7o++9PHzCBtrRlsLxX8Nq1siDZGsD21bA
x78KkYAmmVSm2tMHxpGTQa/Bi8ZvKJkpFBGGSdrmCFpc8fp9/2hLIAT17AQSS4rh
STGHcNJ5/GLA6aegwZDaspnAyNkj4BmZLtWCbLnE/gLoQFml8q+qwf6tmkwV8Ti6
wAzVEmbFe8RAutlDbZQRNmc+Jhelz7rKl04i6xBCcEIVjm7iCQVdEJR4pUROUDXY
bZ8n7Pt4SRlreSq8bFfLhXNlMP+u9b3WB7+XoNLPXFuqGvEkc9sJG2nf6imkkkCt
XceLcc7TFWPxcBEfcD/z0NqhFFtDBMv2viRemLwmuX5/tW3mjSzI9MYLa4/ilL+A
RXIULAcNJ8Zz71/rrYaTFymhr0CL2LDTVMqvVIrkn5UcUm+4u8OGUhSuhQ6wWxoN
pD61N5Mzvtfo8Bjh7q15TGgeYPAx9IFtU2Nfq8hfjSe2bUv9YQtXJe0edyA/BDOx
VcgdXhzBzUC5fAt4wMfkveMKe6boxiryTmowddTp5/K4187n8YAbFDmrAGoaUJEI
qZrcpQ8Cg0JHeAON98WIdAEHAi5XpVqpyzPDxCSRfGB1qAYnU1fErWS82R/m0DYD
2EEKjES6km93oIJzu/9M+D704Jef2ulpK2DSO9q+EKqdP45rTKgB3bcoJakyYYnx
ts6WEoBIXsc7DTZQGtrWflqVOgm0b6zEJZ2JJdRUBgGnLCofdwMpgsQxjFrHLlSS
1vzTMMpcL/Jx8TxlqfQeM36IOPS173puwqyqaowzX1lUww1WxHP3t33SWW/2e5UB
Oj5IoRM8MfKpprvPOB+dm1WTJQ3veL3bg3jZvkRQMQcwLKQfADiikyMx7Ocsp2UE
kv071z03tz+IXmPiAs5tiX6AmjKDNTNMg/xHEeiUmpWYvzn0ADnb47cLfI+mnQ38
ywzM4139rm7DqvGEdd4dqcAraFNyKutA/HaiUydYDE4BYtvq+iJoCHSlwHhzlNIk
sTG2Wf3cGXF90bMfNA+jXT65BYVSEcTD4MAcMoNTZCeNYLXVBMVkd2+uciruWYhW
Qng20jzpxde3hOTcXUsPqvIsBb2TX6LUC8yDlbnazC+ofTPCBQomkkfcaVMnQPNE
djxSKUusgJVsp+NFtfs0tC3GN3WW2P/tbZc+6Xx40HteNZspM/Js5D8uxmXqbEa9
s0jZEIHWvj4Ds/rjNWHq5jGEpnr4BO1+Z4BE4kwTe51EY/lZ1zc6el+DyNR9lSEI
3CSnNU71qYFmhGTMW96kWdfuESsnSAIgbMrOaMmmcrpeeG1zM5CT7hGFx7ZK5jl1
6FqtJD3Q2iVdVuJNbgeOtwDW5GGwrtTpCNmjU5zP6Q2t8tz2qiNM7XGPL/Qi+v9n
9aO00HASjxjZ52UCRw4ku1pHZ08AUAkAB9Lz2VXDie1fjOLxfdvmiO5Ms5EFRzqf
wFfSTbesMo8cZmIKj+FVpHl7TAheZ1GzJk6RCi4dHzMg8FHISJPmVjrOqh3dfGV3
WAdJcwTMvWhC9VBUgklk3q3M1CfODdxjO1OWxfk+N4dLRf7tmFbUhOK9Vr7eabb/
3cWkWF7/DIaQhyU4rtvtBZNW5qYEUW7KHcfGQEu+M/YvwFEnTJqls/SWYwzSh83V
07Kj00mfr/skIC1ck5tsM3JpPeYB1xhqQfDxLM8rOSLaAruXNloib8X01KqCmC7f
s9jWjKVwAypqLBARGWlDbdm65zlblfbrzoA/c4oAbV4yHHTR56hLmOAi1pW8A9HF
0Fu0gDR1jMy+BKlCbpgKE4cS2R6IY+01mRT61QfwBjjcIY6FSuVB+CsrNZbDEs/w
aogezTuwglSRl13ZhDLT1vz9Et0ABARXSkLw99x5y3TH1RnbqzEXOJcw+mUQEGNV
D9vbdkZcNX1PED5apcr3u/IwjhjgSengzRir4FO8scjOGrVwnvY1mH4R5iJG7LqB
zKRFLA2MEnaus0oDXMXdjCcXlD3p1vr2nPJiurxeOVnr2ABvGavsTarNS2wOi1Et
PY3PqyVIxTsBm1V+47aba3KWcLOkxJIxessH1CKgmYJqATsBN04H/61UGhwppmBy
+r5SBds0aplq+6QIirmGUpUiAGMhjg2eTUZKH9QHe+2qxhkaX3q7mY60HauwU/TJ
0PRDUeFYJ9jLWQek5OSUfvy3W2g7AaAV941un3P10TcimMIHRLXbu8rM2l9TOpJQ
wW4fXGLsOQgTcwIsaCxnqHmm046I0zoC/Pi48SsEvkxQ7pBKqWkHVlj5IZpNwC1i
wPanIdCFYie7f78ULwirU9/ZAXmMSafl4L04seX4laqtL9tO9DvoOXfLQlsYesFX
JEvtbj1UURxVUjBHspG+sMrVmDCi/x2y027weY0izGtlQ6nGD7aoXXdTv54WHV+x
8YSldeAXmnXFXNecCrr7XotvWydEEDRZ/NAx/rKjXrpWY3btrr1yV7TemFKrsn1o
oO6MZN/es2/VWeQYyzMQDsRpaIulpPGgFPo0OOEfTccmBOEzhp9vf0C1uGkiAGRK
/S8TTLoIGRDPKZRyK64kgVD0+hv/u1/hSnnNjspNsn4VYnvof446cd7vb/dEJlAj
rQSJUI1k+SfE0MAxdJVDDn9jJm2ChEaJsq8I21YgA9S8KeKywSovk4EtkdN0p1KU
Pw8HKZ/TKMazwE7ROocwGqNDaW7KKaUPZS3h4h1tcGbG9Sf+1A89TC1Su/NqOPC3
FUSIFH7cxpkPGL7PIaOJ9oirMbCWLC9DunvW+BECRmCsNvaaq+LldC6WB/tLMD0P
kUGWTTWWNtSsvFEwZ7PiFAEQi+E0KS5tjkpRoobB8o+W6OXhWd+RWLN8fE0eRQKz
K6vuGw12Z+2iun0zva3EjLfsK7WfBGsWVvQXlaPvrf6fQSatAcAH367vscLNaaXg
aJjRlcUj1/7/dUxB4R4M2wQ0ksLzfWtv9+37sHevpoNAxgdOMpbI2Fo9qq3u1S5Q
6pW96zUUGwayjfLfR721Khnlfw5OTLjQNroFprd4XGdLNmW2gsmtjXl/gQ4x1Ow7
t7gxGTHSuFXddY2zBoEuRkvULXX3yDDQCI4nddz4bfoPl3O+KzoH/KEfjb5yzVxc
zPGM5AbaWmOaeDhj/+klG7D7pjikcmzOIVABuCU/IvEzqo6doyG0ak9ZDXfdNsIz
lYiBc2SCOg7fO9TtiKRgSjndgaD9fUQs47542e5TwoZWyxYno2QiOEuVOsz0/30T
OLAZahp3feJi7csjy0wpTJBXdS2YHxH2R+snITNqtj2XdS4HWnOn1PfpB9eevwoy
G1jf/swtQB9+g6HncIZyusVIw++muWPywPdKvd0DCxQRQacpFLOU8uC3uC/iUfdm
CvKgRkVQX9KZcQJaVTeforbCfJD80j4HPL7+b9brSgWtaRzkdVE5/Bf52+fkN358
kZ5i9UP2BHxA7vqYbZPhksGTRMGsIJRDMTCWyFrqtMQNJ3ACRA4kupAYdmIjKsIq
5C+wxih3Xgp+y4MYny8wQXn36ErABiJiFxznmrVJ5bHmErnCubcOFAs+3tbxqWJb
JrvwiaCB+ZB+/mBUXhYQd4Yokmgf0OzzUsLxwf+WJTDmPCe1BIZPTjhgVus+/o1G
Awv+W2eenlQ8BjNazL16l3Gc4iKoVE3kMu0JLiOoSXyHmAVph3A2SktpU7toyJQa
6DnXgz515nezZZflj2YF/NYQoJNdBxfO4dsfhfIFX2qkiSTCbMeTg2TX5FjR3qTC
CnuzP2AK9WG9773ODunKNlwoBfZkjBscSrXGG/YsBHDfgFr4xT8MOnW9ujkNU+Vf
qLDwxGOknMJF0TdzeEP5nvVKeNBc+KV0AwpcC4iZD1DrRGgAn+cqRs6f2xBlAnlN
euKzZZft7pHqqgObGrJXFbPz4zFdVrwF+ChPqD5jOJaLMoeq4CQtcv/uUecqjmwJ
wQGFIm46ke194k0NP9vN3aDwjoMbl9Q0S0nbfU+IPvhxD6rzPIogIpgJBJUlwZh7
Mgxg2VJlcHwhtjdCtwrqJNVtLJE75jTSS9f5ftL9rn+4bmo+ZEXa1CV1b0PV8Gxx
sra+5YsSlHbomU0L6OY8MlLADQKupwdXCbDBjgMoZl2+6aKAhjOqRfI3F84OpuXi
u6jQuW28k/GnAF5hGwDll6tasvkA4EHQDGW5fhueW8aOvkoBir/tCsNioH6b6G/U
KqyX5MfhvHzre0tTVt4Ukq/i/5mLgVjHlaa6P2UhTHmaP5mEoSgFDnf7zFctxuz9
cF9CvLbtbak/94bsx/DK8ERaQT7ZK/VKF2F4CSFsKjeRT2Lw1cMfqYrmoPedRkH7
G21QYeVdfOAmfbSshjHJDbaByAXDIbXvBDieZjVQbNhIr8L3waYaCBVostM4kyNB
ClJniKP38ENDVn1gITM8vvME+TuWvCHbYERYmjzSLDeh9qiEwfWUsUeoNmx3Tynu
O1Jw0H2e46wLc40mNyYxmGMr5P3GtvzyB7biW8JLIhFK1exX5XzZxoa0ZK1SPa8g
kjXDdLZWICcGkcvS0Mbd0RJv7n/81FnbGaCy368X0htnmj48cYvDFOO3nI7ceUui
CHY31o3BjOITR24TQbLu6kPAyO+IVbFTwIMduhEMG9OjB3Uf5tkEmh1opXeSfnpi
yQh+p+Q1QSCLhtywUC8AYJW+u0yDI2ljVGBWX0B1avgBiyQuwnX/lMo7X/YKqbx8
jSLc4yZn4vBj3Gk9dmAbVuFoK9qV5ZvG4kYrVryhecaA4WIOEfKr65b3YUDloEXw
nVvBRTn5R2sTnRKcfYmGAivplqI5Mgy1eWkurYcl14P1+c6JmIL1xqOGN+oTdUZ1
UY4J6puAVvAz+f5GapNXqub0IzK9X+J6THrgDqWWoVwX+UU+jp/anvVPyQHjiyex
sjwFk6/uwuvzJhDAHs+AGZyDkatrah3ol8og333AESgUpMad+IGKMC5oZNlTMrG7
38CCvsOYJ9xeRiMSSwh3R+oLhA4M4xfJWJrdq1aPTjH512WRyMJCdFZHGHq9W43J
QSPqRvVqh3WWNHK6w79+sg3Dlx6jGz/mm8eefit52NWxlcZIBY4594ke+fFqZAvj
9gggFvMocMw0b2Yvf5jpEX0YC3uXJNIf57ghdaUciuGnRvKzfVKzXqzJDuBleCU2
pjOl3P+CRCtVORrmzwALmrtBt1cmsPE+tNnE9OLUrsPhyEtck0q9rxinhle4gCpD
8/gcIoYmwNbEQySYl9misZjmo9OsEAbYwlAR89xgQCeEU2MUZGwLueLaDHs/IH3m
8OwkuUMvAiR8ARXEO4nIQGo5Q2xt7GPyVVeSk7eRYbS2Oe3JlxjlzNlX7CQA8cTF
97JwKJpuuhpRGFcrJcC+cr7dUJaDxXSd4fc5ZDA+mHA=
`pragma protect end_protected  
  
`pragma protect begin_protected  
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
VVL1A8owqqdRp4y4IBDBHr+vTWgbTbd3u8zfMs1FfbFhApbGiXnk7eZdF9vN5X2J
kcGcopWmhy7KqL0xOLVPxTl+l5j6PEtlj26nc7mdXujxbWAbgQ0MrnehMN3pEDLb
qfsgCyfzFqLGx+xXs3hykxyqEP8xvbAXmA1kr5DKTSU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 21268     )
sZeacAOMmo0rADvrjSTUi7pMKA7r9pVGKjHEGLWgCFExcrPyga5Qu4B1TSiCF9cm
YeUfIuPdfHrxqJh7/TWCmUnOp1xU2oKkV995c4Y84RqjnMIYC97VIbwcFqCVP2VF
QOT0P/ZbvWcT4teFBSNt4NsDJgGpxP//xzXYS6gO/l7cgIqsc4ab9+jMOma3AmmO
wPoQV8xqRi2yFQ4EEWCsV7JxoZqYxULxts8wvIOerIPSCcjd7HQ0D6tUutz+LIsb
+9rArPWolQ9tm8uzTmC/DJb5EfkhmH6k+9AbdedbYurq73+R0Ai3ff2g1gjODMgD
ss4c6zyEfrFglbcy1hOg80mOphsKGZ1LWlIt6fcjrRZG+6ilPHqzTn5RT9eDsfsv
vUWpfH+KPcfOGgxSd0TApOHL6+bB6/iKI6d+FgDJgAIL6A2au0cVe0iZ5bv7XSOx
yGvCy4vWkAB1eZ+7/G2u2Q02lrgOvdFkxhULpbKE65gfzSNzWvdHC4w7/kG+KXql
refFVHLi+H8Nj5gbDmPNh8A789r5htBkr2P+kNQ98ng7hNjmyCxkw/VttLyq971+
UFIvp6ujH9cwhxtB6GcLJr1uVjiVPMKDsQSVjM9HVFIRv17quILIzUFyO6eI3+Kg
3qBXQ2w6V+9QiCCBBFT9u2qD+hDnrhT6g9rvGvFRk+aWLcjnEsFRgQ2kQWn9gQwk
THAy5cyZlHD/Sc7TZ0gaVMIMdedscIaTXdNCGmlZVj8blfhaIkJnaNnGBhUOjmup
Lc8V6+gkwihtikI+LdfHMWtKk/k1MDKOzxZ7lVnVwI9H3UiutDMFz/z3wFrsQjsK
P0ED1t/iAJIQOk2ejTeUFqZ605mpoYVcSEFr78a53Uucp6wG6zWVWYPeWnthVDLZ
dlZNjRp2h2UolmXvCCZyhEXplc5chZfEsP+AxTBM9gdDUkCi22KCvpYVhW1MWKCW
7vg/3O49zmScA4VB7hJK2WkhPXqoelR7zZ/jk1TMgEUKL8ip6MWDaHWzmlNeEHq9
Ubg0Bu2mQyhSqTMBB7H7BsD5HfXIYGa/00t3mUla0WlRYyrIWmbPK7ye/zbpD1w+
b1oZMJpWZ37yocFUT3cO7BK0c0oDGWUAXWK1tJE2/2Ubpt0pwf+oAlPdvd+7SnvK
qhbEEdHO7IrtSsKdEQFmRBv9j9YmS8dT11LS7YzOjEgVFQaovIQSpjmryji0hlEV
C4GPIKuAmHs2ghsFSJRbyZfyUVKGSwdMNZk2sYSGwyXG/Iq9FDG68p4xfCKAABa6
9YHRfcBxybapKEbpn1PGwoJIgwUVZ75ukKhGvJ3MNlqzMb9WAR9Htpbmm/JTJfEy
ELZm+YltpHPDxCE8mwXV6BbqLhpFSRxxRaHcadEUWOqdDIwEAMIiQZPGQB3kpDO4
DRMrk3a/dIJtOVj4NtYCQz+LKHw16MO6T6nK3AQeffdw4wOr+LD26W3GPj214ku2
bFVmxqDOt3oPU6ydWfyyxmoRtJehoa7u+m61/WD+pQmP3pJfcxLm2ZLGPBni6ggA
+N/CuntJM8YC8bEmLRoHuBNA2Kj2Ja8TmEyRjGrZUZFnw0yLmi0mAsDyODzTPKxw
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
HQxEs5uxfKOyUYtcgGu0uoZOBDFS3qgW2/9cTZZZO0T9BLE2Tedm12puHEOdVuDe
7rbz/+BqqUMvyyjQ1YE12k1lZ/wb9snxtcbPFdcwlPZ/ZcGk0K3NWX+SZsUSsksg
cTe3vzxEj9H0A8xPimmfvhTY9Zvm8ch3/UEzgLvZ1NY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 31124     )
kh1qt2/kJKiowjgRXyZIM7yJwFa0FyOza3Y09qFjY68v/VLwPaGmXytPaKD6Xl8P
H3ymg8Lz2aUGy5b4nQ83xyEDvMOrgmghEJVzIaO1oxTZ9Lav3snp+dT2WxwnQeTf
s7/yy9cWqFQvhCnTyMDhmle14fSO/m12Q8VghUvaLNoQw/HxlBc+5vcJ1XNqaVC5
1u7vhYsm0rEKfSMxIHb98+rP4s7DLZre00Un+c11LKIZ7FgutGG06PVbKns5b0UW
T8g/XH9uSNu6a+kn04PyweBS1+hD6EkfZV5DbsHb8qJiYXEAevEV59g0o7Mbc0/x
+xnKTHHYk/nERRb0e5tyBHbiZrTml5lotdkN0FphpyA3EODNMnMhwFKbZeCfht0E
RDjbxTR9LjnRfKl1Dn9uxqOiSeo4BCvR9HNXgJWyVqupEbqdqGpy6ldgu6cZplJ2
C+GVvOZhjXGil1RDyI19o2Yth14BSlV8pvOv6KTyQmvwg1x0sQ3OgBEOD2hrBEHr
CAz7DuvKaTniq93gOFuQgbd0FKmb5xmMm93XFOYVkCk81ommQMP9ianAqXyEbjEm
eqVU9rBBSqz/UtlGQVZcO6g7lRbFw8FD5+rHJeFB4nb0qLx7c0MFMXLBfbfvJ+0e
fCPJajdwA5VPdd3VPQabNLlyPPRpyC1Rmn/Tfbdt/4zZOVM7HgcQodPiut2gt763
U/cUmioSdiPSWWRRSRqyFHoKnDOalvUCiZFt4cPCOjwcx63TW3DFiVwA2SA12+al
nNG8TUH+Oc4cqKWpi5cF+vSeAJH3c6fY1DyH9VDxOHRP/NEbtBSenZNE9c02CEr1
PJIUg7T79T6pwJrKr0EkYRbv+XrVsEmRicIrqX/e4BOxLZ/EA1bcENpaz9WI7Zmg
OHBKUCZa52bCWZpOZDYOKWGcvQ/677Veaa/BplQKFtu9s8HbOdNb1/48bfWjAdDb
K2VzROfKTmapIRa43XOnXN7pyWSnJeYrVB3sEEmRWyzBHyRFYVfKLKn28HL1Rw3b
Sq2fz+xhGjL01/EZP7eJO/eV/LHsHw0FseYdySsXKj0sMEggRm217ZkUEDgqPucJ
FZoXDDYZGKSSviTFGYQeW797vfZsbR+a8PMf8GsVYQpDe3269URfJdOrBvlqbTBv
7YnzXpzgNaPZupONmptx2Rb/blnBg00ZMSywslYr8CgPNlvSZFcI8trgjSkyFJAn
P6RMoMYDxHTsA7gWHZH4Sl+bqsbZI4kLWsJVQDYue63NqmGkg7JDsGSLs20188RP
kmM7q8pnngQbdUMm+e6piGd6xngxZAD9+p96pPW7boUblNjHLHwLyAR9sN8t5yQ/
S1xB4vgGi3tTQYdvm1h/PXvAxNVuDNcTDLqUV1YY2DWkKFiX5t0DKH+6bBDndmwV
nNAkC8ZEU7OUsMyopJJVXsmaPjuHL1Qc2gABnInunIMq/DNcwCALlrNEP6gB75iZ
ZMCPAFjXG23gt+blMBhvJH6i11/Uwp7XXxGr1P5f77xPgJ72qM6UY8eGVkQP5oW8
uc1NhCBxzORJkG9/ULC5mekrZHvATkWQHfL1agMivOr2NgwOUi3k6lsdzcmc1rO+
kHnh5ZyT3+5Sw1ZmsvP2nZdUdhdbJW49gBa2XgMn85rcZdiEnrhvYm6ZdWdsrqNk
upQ2kQQDAHnYBv+6vkSnXbxUfFFJfVKCQESAEDj4BAMv70lg38I7g84N+muvgOAM
IrHYAM6GEPnqrQVyOi+BoZfHEoshyV8VOB6/VRBovemunOGjbmByfdazVXk4PiRg
f/MLerVRs/yihfXrrFu4c/Rjg5zhp7l/mPRkpvn7JlphmJNUvrSXPdYP/hW1dGV7
WmfTpuCcpoM/Zq9ArYE/YL/8BRE2P8ZGLXeupvnIlhuKMjsCxq5MP+b/EY6jXjjl
Ftd2d4EMXJ2eGoNLFXTuwVnW8g99jMy59Mv253dDT0aM8RVdTEkSQj2GsK594MWL
i1qriSjrFzDCA+skpOxJNX1wYVtGaJF140fIaQ6aotMDJ20MTCaPz/glPU3yOFON
PonYgPCfeYlLYIvBHR9Bt/Mo3VG+VkvK1xoF275qrSvAZp6TT8mlwCbUrao5yDU1
wTQqWiFeCbgIKA4kEA3A9LjVVC7Eqx7W76dTeiPRIky3UEh5bxdSEiQw4sMbf6et
+KRKj7sXXk9KlfzsJu1/jbXypfNZL/PR97zNUNyn6X4DAUS/t5qH43BDjcB3m5lI
xiJDt2AkRKPHi09B1ONLGiRzvl/q3DeU2FrMOwP/5oRFcDm//ategPHHalcBp2ch
oxp52T8aOc3uey1ciRC+QyeFEBaVgCQmvIhFOmmMF7iJR6w0K+8ot9mqSGCb98M+
0yGIAvHyA41sTX8zLGJn2En99O/+vJDGhG9lciSX4x1Ui4vMaAU+dfQnPWPQ10E2
6ZahZ3OzSX6InKqUKG/m7i9uU+g2GIUh5F8LyMEw8mTmPC1rgbDJ4dIt1Tj3//1I
Dhj2F6mC6ytxT7ixXJtCFCfiaf9sdJlL4mp11prQ/l56ln3qSQwquuUlABxJ6wKt
Ti9jgQojLnNuGsTvcpn9QdRBKl9EepikCamJfNLwGd5hh12k6KrYnzAGUFjZ/SOP
2sHr9Cy7NDhwPiHPC3NHAFT9idmilIgEWJDfbph4YiJMFbhFFltqv7I2y896jUeX
JYZHiSbcUdUvyHYYbeeeehGaU4dws9pGyAHu8RtxBMTohh3W+rLvgKiaSifptSmr
2Qd41Kt+0mYWFwrt0rZFXzKZVwLwk2h6dxDoJSg/VT1Lwi/ZUFCZ4YfXT4kPR/iO
IQXnpaeEw1cq2WPwmhJhIWWb2IzKV6Og8rALCsw+6S7BxYxJ5rbE8/zfjY2C/Sok
ys7k+j1YavcpHkReMQbVFpk54shKXiCBnOQq3Q7CnGp1uqIvFf8/7XDtCvHadpWq
qhPspGvIex15zmWoN9Ifzm7ZUW1GWytJ8d27utTWHO3gNYVRm1dXSFkvRBR3RPGw
twYRpUUB/sf34hWPS8VxiCBJqURHOz4JthwMBUGuZOW6M1s+UwFxsv85PdCvfyzh
SkdOf14yZAwhwvYunSR5XCnFwDv8+34NcZ0ocUr/gr30rImKJU0GTq1qvnthyfy6
aJ42Zm5oyUyG2OQO16253YpPBs2Kp9XzNSIjRmsjKnVIafkoWNWwa9PUnYMQ/CKb
NBn2nbBfE8KFSl2+udrXqfKCMe2ezXWA75rHeqHSlU7ghQ5blvsGAPo/MBNaQm3A
+rKh7A0n4d41g3uUT20iUJxSCXm9L07/mxd4/iIus7ig9rVEsXX8DYyaZJPXBYQZ
t3bUKFIspowiuq1C46n8mBP8vhHEssKVHMIYaDRDZa2Jx80GKmGPzIp3LXNcFHs1
x93DIRsOdDmDsA5kuX0+5fKSPmNWu+RI3mHDo1N91o5vO4Lfe56fQlEqnsq9fAH7
zniztwxmU7Xn/qsgFdYqFEmPi9zvrAZ389ENsp7NV0WTeySKgEPniBmrJ+linsLf
4oFCKXnYFRC9+hTuyGVv3P2Wuet8cs8ZPsmLRKEcdqnYt7z5zDRl7yA4AGsL1qB4
52s69T/gDF7UlS83wpKtKKBQcpG8dPRXrVLyOi6m16QnmwPPw6bMeZNr89i2JnOw
I+yvPPHEMHiI67qulBi4XA1NA6e3SaXBvonGylvznOhM4vY0UVrTrchem9OaHMBA
/mbEnv0RGJJqBOP30vTfxIlxO94pWBk9XN4Vxzrp60kdk1XVnoyyyDrUD0fPR6vo
xW50beMHymkaxLzvXfcz2jkHNRwsmitExc18YU1+/WLYKrXcXnPosbg2l3DVHYBr
/SMf9lgF76gFkQk3hGMSNJ+TvkRciQoScUyyVN7D/54jWPh0L4BoKM6Q7xW3N6am
OOLAqf4fd2CVPoECo1w7rVvimt4xqhI6ePIOe65oh7LddZCpHzcKnjN0kiqU49Vz
aVBXR1WqXRUStZjzTaQXbGuGrtPsku5+M34Hx3FPfPS5yXfcnuiTj/90DAXMWnuB
udp4wYRGOoLU0geTyki7XkVH5ph1fBO8meceWyc2dJU+EJnDwhz4mZVQQrLx6SVA
mGQsSW5F3zUgwjKy8gPy2jR2vvhuO2icW1/qi23GM09bxm+c/G7tA68dWe6NuBmP
Y6h7sxZRqgImIfb+y8SDNKmK0y9jzFbJPOLyX8icGEVdCnXameAFrnx8ygngPPLM
vHTTBpb8F1sVtr2jcTuvZKiNOwX+PL8WHvlen0hDxplX8zfFOqeGPTkiREuQn1Bc
hvOy/ZfIUlHY1jUMMjz2ofpSHQG2zbef1iaMuBhqdDLR9nEksPlNWFrdP3tB6MsM
peZCCb7nLB1THQTjks4aCNyI/QUzoZDwAH2vzOeUN5WbAIbJ6EP43mGg/WrxqVrh
rWBFZUcY9kj1Lz2ikbdn49gEDeCsPNjS8f5GK8cDJ9lOUC43FWDl997K0a/Q2amz
qI/2aJtPHeVeLZ90nnm5ssSZZW6MOV5cbqSdJo6XHqUehBWJUB2wdpcV/fhIZ5dE
KoaOwhjojmjP8WpHXgLATCHpv9xs3MX67HXwuO0zIMtJ45qiekiZ0MZ8MjjCSJHc
Yu9ufJ+f+SM00uVoH6Csosb6YqaZ8mFNbYlLvBIoDw7jZ7APFdN/wtFIYf6dz/3z
Ix93TX5FHCFyDbgD+LPizK/GHi/VuBa746UTEjgA+u13xCNowzTL+ZIm2eDleYx3
i5XXLYE3riOuXy0fsrTiuPs4EHEzxwsvRkxnwKQ1JvIwqShCOS9ow+k6s7V8dOTW
7zsHdn6RwoHqiHCqjrVtNZmlvn7+SYBjQfthv7vyg4RJLyCg538B8vD6WJBlv+9z
4OdJPqiMcQRVOLZW4j9aldh6tPN5R+rir08cAkzycB+tO/3ZRReU6Ndvwyss14rz
SC4b+XABuv16sxqiWiYrzQUiCVYI7s5fQsUkBGi4yYA1bcTegrOjBHCHb8zqMAJL
uG8ar9QnDkQmc4eCHkpZ+0NuGB+HuqCrMVWuA1rGzcvQUqUi+OOfdbyHJovXKo5b
wfbZo+XzK+75FN6qKCw/86nSZ5ouJ3tDgUKe6WeN3SgbCvnCcKCpPdP/NmAzBFwQ
xMRi2uiHgLi1plZ6YZq0oToNSlzXIT6C1JHCvqQ1Pd3qDhncj8chbFeiHVvsvsbn
qGaYkty7agsisAjISTg/r/ENs8HUKjrlMR6OmvpLveNc1vFDNNcvBFtd1oHaeehT
pI2BQwbetJK8WSm8aTlUBcb3ZMJMCcgsVQ7DWkIYKFgnilJYHSnLeqzEY5DZZ/8w
XNvdlWqBQAgXUT5a+Iy6lUb3r/lLr2buqU7UVnhZYtu0LGKArJJMClpyQAz89qq9
OlLIiTeFpNzi4KdwtujSikYC8A5k8gfIwFTSR8JIFbA4pDHfMwkci2jKo2Ygt7uY
x49uwTp1zMtBTHGOZhQVxtgJYfMNXR4RRmF4ZC4FLR34A76M1EkuGzw6OR6MbanK
zbkfzzl28e7Mz3oBbsug6fx0qWaOiY1FItBEXSFMHhpeFyJ8fn+E4996BjpS3edf
Tpt33CgfNeN1elV502vQrB0TgYnPpqduDsCisdgTt8BaSw16Fvh+1sSUw6Kb8Eaj
lzpnp+YNuIR4Uwl7Z75i09cy4/DZ8Sry2L2A6uBkYY4sHUc4k4Z2y0bSv63E96XR
NW3JMNXCWy+tH2jpNSlVoHg453xEmXVPCQjGQEKs0zPwN/z1uEIuzljggRDgzD9J
J8VobVNv7TDLKIrgKRGn7zynSZTucw20vdBRSt+Ae1PXq4WoQ+lxD2kApWQ+Kt7/
9yoaNNVHQfiQ6uac1q6cWJyG/IbC/Iylum1cxWG5z+oL8i3/fjb+eP83264GJEd6
WCGy2LpualVezBolnqb0LZ1scYYqNYhJMaDOdPCpQY9AlnDliQXAjtVkP4v8ONdn
v3ZDFtQYEV5R7DRnM1kUpFCb9pJYeh99p3cIVXGtYIC0MQdz9f//Oy47WM8igAVc
oZO7smGkEyvGcQ8aJE0SCOHSDB520zMQNLi9vDRHkcBphn3YSGUqnzr0dEUw30Gp
Aj5lhF+IKyz5Y0xuF5UZ1xKsbx+SwzZLEPngkpx+3PYOPYJ1f8q2UGRJGZpyedPr
XHqGNWVv08Imw6vMhkXTbgh0uPO+lVCuJAa4H165P5nDYX1QueSmHaf0av/2fbi+
SKMzY0My7CmvYalYt1i/bxxEMbzbbvUN18+vWVRBYHQGfSAzKbDGFcOD9HhasYH+
4AntZvonvMXSSpaZBkBpim8tY1CdCg9fN9Z0tXJKBzM7nNv3ksSXbFqMqPep79Rw
lVpVbe3uAhH2ySolf/70Vf2aGYFb0EBwoz0UOilMkxP1c/Tb11IHaD7WPNF9cuMz
jpsvhcTcGj/4ImyFv8mqWuwvSNil6ewdI9WzCezhjRTI/chXMiXmpDGvnXlG8r4t
Ta4dTHUBl3yQOztqdOxH5gaHCIeJ4q9A1DolVPV9pX/2VgUjld2Wh/rjPyNQiois
gGUcIRHFwpEgzJi+RIoeslJNDCByrTMSPLlIPhwfFORD2abjCF8sPVyGaUcV6m6o
KDQ0MmyxIPPr3DrGMmeQnfjNWXZnybZPc/yOrTyViHq9IKGGjlfS9aQtrVgTd0QK
CI8XlMfdKfQ3td3xzInHcMQFdTOO7lPXTYRYJtDCxLMVSAMB7vm9F7YP6S+Xon6h
qpc5ztEaR4Kf4g2WKdsmU9cv4GOiotm3r13kKgYie0lknuP6mK2PLSdrRxOBJ2us
wdlDrcSMK9LTfZEoucggqbf4C2DMI13w4pxTKRhyt2gn745ADoIjxJlVTnrfHwyS
pOvf22HZyptbFWUABvyAmICc8cu/YSVkV62m8I3WNM7rd6jJmCK42X9u0zB3SicW
y9u4ktY5Rnz3l31ryACdFCYWrGYO3AmiFdMNrXSSJsW1r2yJfGfT9o3r/7ROJJpb
wnzxwsNdBTHTMBADVmyjwgMOarSeb7VDPYgWb2w79Cs1GKBCR3TNYfaQCFwSIjvF
+v/YsznPSFkDrLLMfcXX+bB/XRTJ2WSqaQNDVNT+MBZWU9ITDRK1qIECTQexBpMV
bofXcyK/Sy/RwTkLQhP0sw4r2uAFpUIyc6dlsvG7l3WxQnqunYu30lae26CAnTT+
4wixuDKNoj9J2AQY7Bw0IYnRP/fa0UPOJSAKjR2AvzJUlorctOvpOp+iqqSEjuSq
FpECdvhFgfDZxMp7dKYbJpeaPDWdpWZ/g3/QRuhJTVo4GKrI9pWh4dg5etBQDUET
hw6hWfjJHh7bvxezrartOt2cwJzV2GNxFbXQ8o1c9QzwGSP6nhjhQExsIPUiC6Wx
JWpo/891HkezOqrQXi1zZKWWibV0PnFH5+0Vx7u+3FxTI4GB3SGkKWXVxbBlIvIc
yBzbxptQSXtspwUwIfIHfl/nEzflmLI5nNmZjsmISran/t3Hjy4OCWKTm4lf1sjr
l8rehXdmXqYtgWKgxRPEP/ZBE+v2eXcNHpoTVY1cPj2Mvq/HGR0yOzpeMNkgvj40
YV8GVKZT2PudVp8Lo74kIRYW0Zzox/93cCGD2JjRNXADeBDVMNghnC7AoMndkNOS
tP9/F6EZlnS6jVmg3RHIrUh69TxqP1z5USa8bRzDMNRVriHmMjfYmANb6a1yk7BP
vjKihqF4iFkPvKahLkSCOSxM0hkABHUa9NIG+Emet0Y8++O3sOWRPZp8xykDcWxs
to9HcnyInrK6NzoS5cyBfgKCM+M1ET/SiZMfvqNRxs4HZkG8IVu0NXqPUWMVGBbB
Y/hRqAh78Y3dsYD5N9p6BxPavLFG0lyeJcM8RR0EM/4QSZ0MFF4UGaEvO6b6XCwg
q9bxqIAZCwL5MjMB/KdoO5nVx5AQ1+Xfv+uyOJZtlf2Cpa1Zz6drvYUYH4WkVVG0
80W7cnTdgT3D1Ztj9OoalJMt/YpEvirDTFMxsbZ80lWcaHM4ttcbQUbkutD+XQSQ
hFxBPuMU6XHW8SLO8Ic4UwQr1DK12sVIZ9BRg0kV/S3UMwXYKAszhjwLAZ+7VwJF
pSjw12xqy6UmPy1hTRwfw9LBIK4KOyqjpVvXor5eGra3P6WtOOJ4o7nk8u3aKzl4
q2oa1LcVxiOIDc3VV7gzCnFMqxzM6VQGEcvWeDvoukRUDhfHvI7wdXdvppk6toqw
3UwHIQ/vaAL8CK3JWQeE+W49xtjMG+nIxvNmI0DY1OnpeL+TC6M/qlnH8WibKJIM
qWzNp8NtSxQhI98NlviK/qc2oSWRL7hE1LeREbAFYuDk37mgvrq12q2xg/jFkGkt
YLyybwT7ZCU9iO0rM6cBTcYon7+dkdeP1p3Cesacf2N1BPn4s1Koj1SKPFRTjidV
Fo4sHWM0oXugpPhCpbZ7WVLpIjNWQHe8wVNpPBXydT6Dlg7OiR0XQhjjWvO2iOL9
eynBt0xwiwflRB1yI5jXd5TekexoUhh81dijkONpiT3YsCpIilJQucWv7CMsOoUC
aVAAGi2Jk5iMnl5i3rdAF7ZiDrTc8W71jvKDEOf+igz6BYkFTlBYFi40KRpeLYIq
qgEXaCocNXNGYO6b1nfenL/x3f9aQnXWF3WwwHrHtymheiOMq6hnyVVAU6TXzyZt
MlNTKV7gzyUQQof3kZNG0l7op3k3+B6JkHVYf5ZSFs9uYy9QhSEmopwJMrjfZ4fp
HhDEL1DBUGH05sxnHai+2sSbKMf6sUcwegP9VDZVicWFQaHEUERwwY3n9gwo+nNW
khT6MOhJ2Qt7d9AyY3GEmQPil3dXSD+5kk2JyShhk8C86Y/pgteC1463683GsnpI
VSofcTilf8W/QIBJjNf+UJS2LkUOUNeGCOLeMZdgSFJ5B9jpQD9KRkzxLk4Hu7Qu
8U6U6HEixIR+sVyHXcHJyF7tTwjEVL0scWEblyOLosbslhc4Q3YdmwCYo0b82jD0
f2QTFxoGhNphxF3gHdCMwXvKm8UPS+l658mUNrkMT/jYX3pTDk+7WtP6w2ECs/25
fDWtD7llSqHvuXIze2j0w+eymlBKkhJ5Fgn6J846qCj8tifSBkF1JdTWzRO/Cfhd
7rnij1DfaWLoq0c+f/rFX0xFh+OnDuaUMXCmx6LiOuTeIbZbsEi2i705L9P+DSjH
WDKUpqjcY7e3kfmunW2SYZghqyQ2Wb7rCDyzHc3QLFphQ3RIX4jW6BmOACPcR1dY
ymcYYiay5RGX5xCoIxF8fKrICZR6fPERjLkH+YODjIHRqELUJqp5hfcdSAqc6byD
zmMeNUeFfMf0tg1ic5CMzePzdcif1MO5cM7g8NSZlWb7qgmuUTt2tebsqS0+5T7Q
BaOYBkMlG2Tk8BHuV2wFzXlWWn3nkWsh6BxvY6bViPGeglQ5Phx0Q9baZHCLOC61
I+wFEvl8Xk/z5NRQ26NT6V4H/63wfMCk0530V8IEHnRLRk5pfVlzOWj7Wj8cU57L
gzQElLZDvNFc49xUMDSoWoAd4n+YCgA3hbsNKsfOB3CuG39in2aXspPkzHm2xqFw
NKjWsfYUxxXXxTjbNHUKpyLvOPlHumEBGxT7me9gtfSkuU12S9boEey0vDQeLaat
8grsvew41Zq+ixtRrMPhSa5wE05DhkRl5NRH4jsZ68LZwojsCaaGoMKEVvTRqIyU
R83AFA9LBZMt89wNrBhME0TMJG/nChcVMxlSi+VI0fskMFXVDM+8mn245dmX1l3u
d+SC8ELRJMd+zzHLKu/iNjDtmg11BRaAy97SdmKWABSWIo23Sr84LMAfh3diLDz/
kGwX/KheFnsJLL0K/BiDlTp5OKU+wBQjS9BGXeOa5Ae3XxNa8K+NQrDAVSdpA/57
PX6/NrHobjQK8XaJSszkG1kxrW7kS8+UBpS3SRI3RfVXMT/SKDZs06A5gdBz/DkX
Ve5xSZ+ySmEe2cnj+cc7dmFWIBaJGnNcdErEFD/mh6tiRjXUBbvaTqhR7m74L1L4
tN62VN4PawXuhEtZSnetqQAFgGqaTt+PeUUt/r1z4alsJ6N4z3yulOUCSOkA50ZN
NK97FNBfxh8/KyJftU+A43bJRPEYMlPGA42RkB5sx6zbEJ7LrUAxjAZb3oboV5VT
QBjpd+Cuxtzgd6E2BemyDSzyavUW0X/19NADdfkS2xhK7wOag+1ipj503d4Ep58o
KJadHomHVfQEhfCsrcgyOJHTeJ6K3u89WUjbt6vQybyz0u194XGuie1syoZyQfhs
JvhbOmDSvz7m8AicOHIlXS/FYwgBFiQIw0BvZlf7I0pSBfcrdcBnOVZlcVZ1QXkx
scpbYaaqbDYD4i1IVvGnz2Pt/YfjRpv5reiFyILIH6aFN/6Z7jNLrQJkcoqo5F0+
w8MgbsqD1x6XMqZO0Mo7ZH6KaBw9c3SDiQgf8rExsWqG4ZaDyABN/5HolISbrp9I
3+nEThYPJrqmt9xA6Ae66OEWPkkBtqxihrHZeOc6aXdsKjpjeZCPDpKzKwwkmLmq
W/0DC4vmA//U/XoqXDaP0yj8+D/i4/kBlUK4VLOyXjhoD396zd1GaRSZvZJE6vlg
7w2piCRioAVsm7+uVrjyAz/ClKOYz6xWwAl3p1bYG2Bg8QSlMl414GY+cHXHRvcw
VO5lBiJlkBcSKFn7N+I4NFVK8XRrYrOjZcnE+j8gTPYTksg7KUwuldjXV/JI2CEz
+iABmt7pfCsckBEAJ5f9hKIryAimQxhWPbXPVZvy7mTiabYymyRCf5LWbUGbce2i
7ZobFoMzzfVgbXZar1/3F71wBNNOFcaNN0aiwDXEYdYVer+svU/FP/H38Q5XFw+f
bsV4To0OcpGetpTliNJ2WC/ETyhCh8NKIHxKdeNdqRGgkjh1Rx7FylcRlEzV7/gR
9DOTE4sIKCqBiaIjFuWBaSEAvc4iS6N1n26JzqkVgiWq2R9n0/CCeu2DRZp8jZUn
skDFkGIblRQajZNjLFl9+IPu68VLQYUqaCiD15OP4KXsQzzVmXLpcv4LA7qqZuD8
c9d7BMJ6QUWuCoHN6/G+JI904rvM+Q3SGTI7Zh9XNGL2V3I+V8bBsK3MXqkapTcq
wH+MDjYrYqB831eU+rPEKm6B4NLqNZawo6MxoTQfP+IKUHWIxnd2WXLnvkLOF0kN
6DpL/hZ/Vd4HCF4rVRNsT0iz0p3UX7J4f6er25b99zA8UI3XprJz3P3by500+2Bq
6ff//fSaFoUjOPu09/fY7iBnOzjOxg2VfYPI7vho3EfpT844LYYfFpNyZ28CA91q
INUekDLFfNEJ6q8PDqdwZIznQRg+llyxMr17j15zsKYkgKux3cYVng0ASzM9Yuoz
t1wS9L37L8UO4owMG56/M/g/92DqktqtCbiK3uBnfmJq5vh//H7SbUlfXhbT4cjK
1wYFe4O53i8ghu8Vie7+8PmC5WIX9S8WevC2Uifp5yiCIGKzRhwSoS1USw448f/h
5EClZmlDOfTrRJ4mZi/EukqkE9avDWKeOsADjBTpnGCzI8covskhD4QIo0jKShML
UZxKKTMFW5fAP5cm6a5D6A8vLUKcMHSyS3p3n/AVAevcancO7Sa63/dCCQ9GH2L6
npJT4cs+48lAHXpYFgDEpZ/XIFL3oxq3T8rBUtxu26j78pLr1bzIEs+mdaIkXet/
N7uMJosJhfPMqcz338gG+4kApQ6pPnGzZM8t+n5T6drHCR76HleOQai/ifOa1L0O
GHcn7vgMvCjOTJY9eeE1Gsv3VnTVWJJlDJw8fmdjqjYClrR3qeEEIpEN68E54Sko
iq/WstLG4vodOL0D+jxRo7DzrQft1FOoZptqae0lvbch3Fuioi1QbE3V+7h7+0gl
u3p3G6lmx5wLMqhIc/N+NGJMdcTehMB5mWBh584bKuJtzYB6ZuNgyNPgrEzeYidF
VeB5YOJX7l7A07xA/bOyGsQo4cS0yLU9me7MEGpKaATZu08/SuPQSS/WMljd4TR6
nhOxnj/mZuGqYC+i3ih/yBiqWP3AvIhIbB6tLPjyI++ZUeHhry7GZW7D5rwMy42c
eFyowD6oVGHwUo5ho9Im9+pp6vbJo0X58wf38J1zsrAYHcQgi2pehaxsu8tcSLnM
fFPX7MfPtVfb7qhIYXbV2IMsCw3cVVG3rm9MJdzNRprXVQ6QEhGGSzNgqbmFyzuT
1qRqg6jhmxTz9esUw6+W0GbqjkKII4iDQeL1uBoTdPUCxjmxDhOeub7bjQTZzJtp
P47wIHuWSH1MYnBVUUAhQqu1Hwp49I4AbLaNVo2PR1+DkI2oih0HLoQ1s3lU2qWb
evHE9OQD/Pcoh9u93ITsSa9tEpJlnbp6WFcp0Uoq9v9PkhYHTIbyQuUW9laEtj59
Nu0BnS06Wi2/E+bpzLCmYBZphaRYuNWDTKBNeOP82Ep4dJ8zNCBC5l3/84K4p/2+
Srkk8AjFC4BwHuKh5CqXeH756zR11eV3sVgjqL0Gzv+BQh2StUspYrU+3ECC4zop
d5L2EBRhplhoVvkgXDDgB7hcwa5GAHQDO86DgPy5TnnD1iqrg4xLrIWvm6vXR9nb
sSNoRyJ2CaE/mnZQc15TPmuzDCCk4d/jGHvJO3SFWu1rZisZjlr8HFDUJCb+x1Pd
cgg59mEhePpFNhD5aLJkwLSRoM7sUV2sjhK9guN16YfzWe7QUpEVgK63JiewGTLa
pig6bDPB4N545mRhQ78izSMR5Y5/p+cbkAmi2mJi/UuNDHpqFPV6CCfCq4C2df3t
fjKlNlkMV1bQlHG8iK1NrYhA4WFT9CHLYVIa1yiLFTF4aUjmKa48rWDp96XONr5z
Wb08ID/aAk+RqvMCmVOIwkszuvL1PaZ7WzWqxYvLiISrNVI8YhlWBiRC6A9OIyEZ
khqCcImOq5Kb9XYBzUOoD9OGJZdzvHJXNKTL0DOjSaO2LqobIU7AzEVBg2hZsFIU
4xkai2QbqhfT2NB4lWcYsyPxZJPLIfpTy+zRCkumXmS2riuOH7J2V4YnPaRSkzgE
l4NIW5coCAQ6aJ5JKSmARQG/D6MRpjfa4c3BJe/+TvUIRozhK0AgzuC9tAfSSOP5
vfW7o8Q+p/YMZahvfgHTlMxOlwZU5rhafcIF3V3sPZpRMYnGCp1HMKShwCHrHAUK
RAgBVfRgt+YH9mmDTFmdkIE90YKZnXO0lISb5mz7p4A=
`pragma protect end_protected

`endif // GUARD_SVT_AHB_SYSTEM_ENV_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
REwijLHo/Sk2KEy6YWrMFcpvjTNNBbrdKOm444pfMdaw7wik4z4g8zpq2SKDNtzf
q9jy0dLoCjhlrA1lk+XoXj0GDNr8Z5PM1LyZtPely3i//JUauAI4rMi57vXbcjSQ
Izd3InQZJtPtL5wTFqoKSDh6XYMijsVQfOsdabTWfec=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 31207     )
ahA3B8BmPhWMdpgnn9knwo6kgyar9ZaO+2N7xxyqvenPcg/S/VyzcQCpY8TKcKZw
BYyXsHopOis/Y1hbz/1wKCj+ZNQ4Ol1EKhs3vig97lJ+r+thKPTimF+WPaEBExRz
`pragma protect end_protected
