
`ifndef GUARD_SVT_APB_MASTER_AGENT_SV
`define GUARD_SVT_APB_MASTER_AGENT_SV

// =============================================================================
/** The master agent encapsulates master sequencer, master driver, and system
 * monitor. The master agent can be configured to operate in active mode and
 * passive mode. The user can provide APB sequences to the master sequencer.
 * The master agent is configured using system configuration
 * #svt_apb_system_configuration. The system configuration should be provided to
 * the master agent in the build phase of the test.  Within the master agent,
 * the master driver gets sequences from the master sequencer. The master
 * driver then drives the APB transactions on the APB port. The master driver
 * and system monitor components within master agent call callback methods at
 * various phases of execution of the APB transaction. After the APB
 * transaction on the bus is complete, the completed sequence item is provided
 * to the analysis port of port monitor, which can be used by the testbench.
 */
class svt_apb_master_agent extends svt_agent;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual svt_apb_if svt_apb_vif;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** APB Master virtual interface */
  svt_apb_vif vif;

  /** APB Master Driver */
  svt_apb_master driver;

  /** APB System Monitor */
  svt_apb_master_monitor monitor; 

  /** APB Master Sequencer */
  svt_apb_master_sequencer sequencer;

  /** APB External Master Index ;not supported yet */ 
  int apb_external_port_id = -1;

  /** APB External Master Agent Configuration */ 
  svt_apb_system_configuration apb_external_sys_cfg;
   
  /** Callback which implements transaction reporting and tracing */
  svt_apb_master_monitor_transaction_report_callback xact_report_cb;

  /** Reference to the system wide sequence item report. */
  svt_sequence_item_report sys_seq_item_report;

/** @cond PRIVATE */
  /** APB master coverage callback handle*/
  svt_apb_master_monitor_def_cov_callback master_trans_cov_cb;

  /** APB Signal coverage callbacks */
  svt_apb_master_monitor_def_toggle_cov_callback #(virtual svt_apb_if.svt_apb_monitor_modport) master_toggle_cov_cb;
  svt_apb_master_monitor_def_state_cov_callback #(virtual svt_apb_if.svt_apb_monitor_modport)  master_state_cov_cb;

  /** Callback which implements XML generation for Protocol Analyzer */
  svt_apb_master_monitor_pa_writer_callback master_xml_writer_cb;
  
  /** Writer used in callbacks to generate XML/FSDB output for pa */
  protected svt_xml_writer xml_writer = null;

`ifdef SVT_UVM_TECHNOLOGY
  /** Handle for uvm_reg_block, which will created and passed by the user from the env or test during the build_phase, when the uvm_reg_enable is set to 1.
 */
  uvm_reg_block    apb_regmodel;

 /** Handle for svt_ahb_reg_adapter, which will get created if the uvm_reg_enable is set to 1 during the build_phase */
  svt_apb_reg_adapter reg2apb_adapter;
`endif


  /** APB Port Monitor Callback Instance for System Checker */
//  svt_apb_master_monitor_system_checker_callback system_checker_cb;

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Configuration object copy to be used in set/get operations. */
  protected svt_apb_system_configuration cfg_snapshot;

  /** APB Master Monitor Callback Instance for System Checker */
  svt_apb_master_monitor_system_checker_callback system_checker_cb;
  /** System Memory Manager backdoor */
  protected svt_apb_mem_system_backdoor mem_system_backdoor;


  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Configuration object for this transactor. */
  local svt_apb_system_configuration cfg; 

  /** Address mapper for this master component */
  local svt_apb_mem_address_mapper mem_addr_mapper;
/** @endcond */

  // ****************************************************************************
  // Field Macros
  // ****************************************************************************

  `svt_xvm_component_utils_begin(svt_apb_master_agent)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE);
  `svt_xvm_component_utils_end

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new agent instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the #driver and #sequencer components if configured as an
   * active component.
   * Costructs the #monitor component if configured as active or passive component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   * Connects the #driver and #sequencer TLM ports if configured as a ACTIVE
   * component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Extract Phase
   * Close out the XML file if it is enabled
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void extract_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void extract();
`endif

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the agent configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);
  /** @endcond */

/** @cond PRIVATE */
  /**
   * Obtain the address mapper for this slave
   */
  extern function svt_apb_mem_address_mapper get_mem_address_mapper();

  /** Gets the name of this agent */
  extern function string get_requester_name();
/** @endcond */

  extern function svt_apb_mem_system_backdoor get_mem_system_backdoor();

  /**
   * Function to set the port configuration and port index for an external agent. 
   */
  extern function set_external_agents_props(input int port_idx= -1, input svt_apb_system_configuration sys_cfg);

endclass

`protected
0]VTfK+-Y:0-/]>aPD110bG98WbP\[8RM7FA1P,W9UVW+K9#E&IK4)9G4+TP34M.
&WY[(VC#4ET.Nb-Ab3aPJ2-EHg2(,.UH>#^/47POX0ZRgAKCc0=N5Eb=4OfZVQ/-
6=(3]4F([PX@9H\,dN[7L#3c?.RNRHKdKc1_QaENJeSC:M0/Cf8;_+IQ_](ATe]?
^C/Sg1B3D<cY9+9c_EN-DKYTYY3XT@]V9/?(DX]e#1cALZ0^IU];3L^CE_BP09d_
89ALQVVA44\;_YXY,^\#bZZR]Jg1-V&@.J]]ZYD4dYdAC$
`endprotected


//vcs_lic_vip_protect
  `protected
N7\+I=e^:g>Tb-fX3]S7[&M)5+PF<5ZX\S]E+;)&B@IbMKDA-3Z2&(9ZM,.E#;/)
b4ZF/1L]0N+_N=dHf\KfK=XdV@FD>:F=I-;d0(-&dV7A_-I-fE9;f>06Z)D/gW7I
X:XQ@UXU@J<\W_;,),[K0MJOcFG-)1bY;<7+JgNC:\/gD@D_R.D0Ba4c/@bM:52.
LD8K[,#A+XP#Z=#aY?2c&>T09ZBDXT(3e7=?dJ>GMTeUWae3CXB_ZZ[98B]>&eA>
dCEZ1^bcCVQ.2I+X1d7LgPA6RI/B;7#^fDAOSCd_cC(<Q;aC<#H96e)=ODcTIKG7
P4AbgOIN?d>S;d:#AEgA]#OX6=3gg27bIF_68[A8Wd1B[?H<G;fL\#;Ub,7?7MT1
K70V78g5?M;QAH]E6P/ZHHU_c6G;I-.BbV5-]eS+eFAbT#O^<?N@f?0P+Wc449bU
D1?_)R=[PaA-5+LWdVa??PHRb)CD]X]gX]c7:,eU9[e__ST<a80V8(0CWH<6S^2+
Z;;/,=8#acH4.CT1A5MA]JX::>95OL7BIU)N5]&d585Jg?58Qc.UV6MO4(7cdO\3
A=Ta6gKG2VBJb/VTaccDFg&BL&#2TNY8G#C[#DG06CN7<4f&8U)YII&[F:S0PJ41
<Sc<(6C<[(FS4DWdAPI2]gNS?8Vc.J#1P@R9]:82ZOOFB-S7(,U_YgE:B74V_/g5
XE\K73,&R6bCDgfF(7^DP<HgdYA6_gV/8HaVHN-#[X_0V,V2a.\I\c_M-OU2?WZ@
_,^C3<9@Ue9[/V8]Q6_dIB=E_+bYRF.3Y)/88P#C+)3-e)E5A^O4DfEP@<[If0DX
^82faXH6=-+6I50C)[6);CB[\=0HFAQ[YN-1A(#@M627?0()FDCJ<^Tg(S3729Nb
-<X/dd.=-JeaL].g0=5Kc-bdU\^J=2)J;ABOT0Y]+\f:,@;c8W0?IVDSI-6aB3#=
L@0W]MV@4J=LcS)#a@S8>_WZL@(AZX0M3>[NLLa25Ad14S5E1[UY+7aY&+U@=NIG
M(LbG.(1\HW;GW8e3).0\6bCHI\04Wb978V[bKLbN3)?Mb6([K9Y-I;_NTF#EZL6
fZ,2fAdAT#ZI=?fS,)D+?K;gRgf6<Z.:F[TH\dY?&#/)(<Z5SL8YF-O.>>X:+ONd
2c8Z\^N?:8[(MEJ.@L=4HD<;a[aPH<;d:b7(JfbeaO^IbF:gffadU,4<CU)^VR+>
;[B_D;A]-_OfETQV4BNEH/[-C&A-cIPB/7W:P>0+4G\&]J28c5ScgO<d;I;cT<YL
HM.,4b_.I=[&cJ<(gC_TJ0b(D[,#cXKID+XH8\Kdf/aA2:B:8?a[W(e4>8dIV0PX
L:b_;WC08ZVeG1_TFK:#^X#(F.09DRF>250cGNZKd>&\.c>=fGaF[]BI5eRdS1Jd
+11D<+4HC:T^OQ.+D-^<O1H\a^9O+W<YH>WcO]S9g5=bX6]X/8GbQTP^I;d@9S\R
CRde=BIK]=9ID6JIAGN.Q.1N4efP+6;(P:.)J\2&7e8U2-ZV;VC#G2(0EZ6W#aTe
eVdI3?b<d:L<I6d9/4L<g\5f3T[E+WR>[V)-OcT34Qdg7I<3@=U3FII6;Od?P95&
;f,<:IQg;PVD&KWK3DLH\B-B9G#^Id?=L9_BS&3CKagO2g3:>])&Y;AXBPL((AOX
#EgC2\3e#RE6)eQfB166XKdRLGQK--4U1W2K-1Q,:654B<&0Q-]b(I?OA+126b<U
+Wg-C1,?9WWB_@<C04[T@ZS^+B/;dZ)O<;?DSD.9U.gMD=B>D35g)NH34Q)Y3VEY
TK>(DA<V1[W20+fL@R==W39)HNXEX19OOH8IH6QJV?PcVV;10N)3Kf,+KDY8f:^)
7E01;+)MYLSNBBe]7C,4Td_;4_?+,8,5HdFG6Xc5TIHFO1,@3de+Wf?\-B6H5eJ-
/6f6X5X;\TPE:3^0=G]7:aEB8VV/Y]TW&TLO@TTF@Q8/88YgX4WI3fA75&YK:1&M
6?,KGBEH7HC3?D,NV=gGO]VHF,O[1<L]PP<8_80BVc&?B+MW6W[f276M1XNDF?0#
U3\(G74^RP0O#cTN1<:+c9]U)T&JdDe&1)WE:N9E)JA;OFe(3F6>KTKR4__HDgOV
LF>>NX/FIK0/JYXGK1\5V0d2(I(><>,=6HQQB>f<b-e.)Yb\5>7LBG8d-Bd=P#gE
^QF&O)@-<<+[f[=>MM]b@T0fA1_eLM]<ZPS6LcdI^Za>HeAH&&84gP9324IQ/.gA
V\Va,?NVT=:::\\e@1DcNFN1S78+BT1:B<a1dI20@NcU?[))3dHHU[=>;@g.\V\A
R.]N8&Y(A@]ENZC0b1UHC>QY(8EF3@JdaLGS/(JTB@RT.VYV5>8,2AV\c[[cZ&Y<
/@?]USSW7a=+)BK)W/J#ZI,JZXd7T9gHVL[8)7(-9#[F80\RL>YDZPGJFd11+DJ,
g_NN(5-VD69MX714a[\5(dB59IV@Y1+7c@&?G8NE/:c=-HHe.WeD0AGX5+_K3:4>
=]JO:RbSQRaDJ09A)1YT)]KZ(67FX=,30gS^Z>g:aUG-G:40V2\\6,7]^eXCg;QD
7^YS3>,YQK3I)e22HT91;A(,\#I9-Uc5a.^bR]M[57)Z8Nda-LAS[LJ#E+QK3&g>
BN1J=P#;I+G_).G87;>Occ[Pg>Zg_Q]D[\bXT]EKE/V?4>>_&6I_RF0-L7.OGWTA
Hg4b/9[]G/;(P\ef;B6cdHf:<5<6LKMaBE1DcHc-_c:#R3Y&U-Ob&d:O.-OK\,_O
(.b6&]bG;P\,MWYcZ(?_aM=B9]C=_MFF@3_eO/.1U>a42-#_JWJL84^1&COCS#O<
U:<8PG1G>7II].]VcZ-H;N@KQ3]G^EB>@[eNL#ZU<1LXe-BQZYV0(,L\=3(bHDHQ
DWA,b?N@WcU_ZI=TOJ:\]A)Q+<Rc>5+QcQBaU3>@-R&JVBIFHePe#5[Y6(/PO;-K
)3#]dFJN#?4BV:]_L1aWO=XBGH\(=N+HBPWFM?#4cdZ@@I,:K3=IJFKG4/NQ@CRE
TX5O_fc)\;=0&eTK<=<[?038/Oeb./d>c>O>0#C=-<C7c@S^BK^4GF>bcT^6L4_V
cS65(g;1)61UeI]L/&gP:f(QV;aIM=f;=<;YNdA3T1U=fHO1;5=XfCL0NFF92\K[
>8PcWZ;7R13,=6g>GE;[GYI;<I3:J\6B7BI3efcW&DN>K6.XdK/Y#CYL@D[R,;fG
U&Y<\I@0XX@9]\(3eXG0])R(-faZDbO_7VZA:3dZVfXSEV(8PSg-8]S&fN\O\YK?
N9E,&9B+8^G>_8K&L,=c4R/?+2-gQb>I;7#Y>/H_T<T]e_&B]I_3--(38@J]_eCA
Wb_5ZRBR.4,6@Q+7,0?)UV1^54N@-3MS-O[EQT__M;93:X46:d@4:]fMB-OD.5A6
La@]^UP=CB4C#4#,XT1OCLTg8LHZX@5#cB61O=X\P4C&]>eDD-YK84_/R60=.<6W
ITV+g3-7>F?gJ4HQ;^SG[_PeCP1caFG_^CdWS4BdeL#M0e#>,#a5LIa9<AW#=;,D
MGTNCS1&3M7gO<)P>H6EZfeT5:2&3VC[Pc6S6-S.B+W&F]bR#L86UA.^fC-<]8T9
(W=3R&6NSg@)/M[L[1g7\LLC#L&_g6^+b3PNI&dZb4EgE#TA)^FS&IAIE1OQ^EgL
WSPMMV1cfM.G^]IQH<aUTUdY@Sc[fZ9F(4gNJ4#,BG^I+D;,3PK>XD9Q1=[Q1[:g
7R=9.aUgPHB5OF/e;,.LX,ag&7YWF&D15eH;0_VQZ)949YR@NG=)W&1^0J[1B)3B
O7d;aQQN^B=UaLGNYX/^PFJGEHM.:ROXC+0?\\W<>M#R\2,2#[P2]fX/&5HGLA2D
K3a6#fcbZKNF&Af?8F,?E2<,TDH>WVf#<^^:Z,EW(2)V4IXJ)8A-:_C/0M&VK/Y/
/M_be[69(1;93:Oa6)Y6RYR-?AM6f<d?/90=F(@.:c[663<8?f\KKIB_H/XWU[;)
XL^]0,2@P=532gT+a92((_\;C=d^3QRZ=\^SV&,a7Y?TB2/9:_1_JaLH4T\;MMN/
^,0b-N<R8f&.O,-L6D0ce+OP@-3;]H),?P&/NDQ#B[YJ:_3Q50UYQTUUC&8:8-MD
CAeS3W1136fY@c;eFH^ZgAg2d2]gE[_AH=eA39-??E).BMC6^8eA.g/\_;a?=e@L
f\f4D<;:Z9AcZc/TeOQVRB0VM>^=ZaeFW;907cLE#ZP_&K[BWK3[]P68&OO&KVP_
9+0E.NYO<Y<d)/bYUQ10eA<KF+F##^TgZ7E.(T&PP8-Q)7RQ:++1a6=^V:CL=4JB
Cg5aAD\]J3[OO=W1R#gcDD)4;JDEA;0QZ6[7eY6gW\;M^HY5AS^P^WKdQVC]g>N.
LE8]cKFf[F^K>\;;P;@7E;>\N4HC_K05WAFfE8DbF3.8dcc;eOMAA<g0^eV+W<<3
9f/T@f7H^;\f:9&D2F#0aeN@2B-c277TOVH7fZP6K2_WLXYfK_Lfb4V1=g\95O4(
K#I-H-8SH[+S1M(5^S+a&bA1)A,WL+V^a3V++6Y&Eb(2074AO55b,(;Q\9@F3K31
)S/15B04^gH#H+MFT-VC<0<7FV4@@3B-E+BaBI.@\UPF;UC]Z,<:@gB1@gWZ,D[d
KJ@J:4<TN.=cM-,7=_^]\5Y#ZJ\O60/-KJ3N.GP7T#UcPR>RA9@LFgaJ_d,Q@HdF
(PA_AP-M61YO>:;\F^KH\_5Nd4Z[6f/;QZE;A#K1&Z_E3L67,&_D3>Y;)VbVJA)W
dRIXNX3(LB.d9?;I;-E[cg??4I_]:JKV/];W:=#JZV&MB6U>f4W[QDaX5V+GD.LM
[H6RF5,-MX)/c[0gV64(2O.KC<^W@KE->2_XP#-4e[Ace6QPfeLeW;A-FM_0P?:2
8g34I;&PC\c2JX1R-/&;CO[NXcf7KH.ePU6T7gW,,-a<1La?RFBe[ESF:+K(fa(b
N\S(H<b;?&_K\S+dKbQICaAU6e/L()WZ&G+&XJBDf,d=8FbT:0<ZcZYc5/CDSM,D
.KO)db+?I3bYd<BWDRPU5RB8Q0:U<U<A(7R[\VB8W4D]FAFeAN)Pg7EJKL,ZDT3F
E4J2+d(V(M&>,03_2c5LNLb7/#2615JAb[#4)@1/MJ0JP5eF6WDcRCNd/X,UPLQE
;H)1J6@-I#c,B\.N/E=_H(YIP8O5IK<;+PE??,X38DYJ.+LC/?d.@\A1g9LQ^Q.g
W[(3fSAP+G5FOUQM(F1Dg5bVgd-^ZWT]8Z9DE(F:]#Z(fYNYRV8TdL&@Tg8eAbHP
:+cK0[bTF\,Ya&,188?J#1/<SSJ6XfT].Pc.YccNQEeYA&237+0,b5MRGY7HUHM1
X\#c(OEb-bF0L(CWVRA,Y^bA<.JQ&#RB-AE2=_HD9\)aM&16AgbZH&c[O3SXg4AQ
:/=-LOUNE@E/:.bM4;LG3&f(>;(]60C-LAL5,RL>a4L9V+M^c4cSX-0NZHX-UPB?
^.PdN)&AJE>d(-JXS+/O.HUQ)M;WXcQ-X:UeBG1MRMKQ9URdW3YbXOQ0>>@^_+6<
]IEY<30BcL9#7CHBJM,IZ)X/9PH4aBR+)):I)[G&3ec6<F\X?MVATg.,<X,CT-/^
U):4BX^5,H-=B>^P\RFIS<f58SZ,,U(Z9T7ggec0e_UCdXI,BgZAGYMDA4OZ.R\d
INEUMB+[6#B4;K9VQ;\1GIFc;^E0N1UY&02S,ZR,VfcS9=_/U_T:EJBU;;=_L)8D
LV+@dTKW)b==7c=_Q/[J467+:>_a)P@PS^5RGPS9EaN5@A(6<]Z;[SO_(dY.<:]D
L2/E05]E)Q<:3XW[dTW/TH2N,U5RR3Pf)0V&48N:=K@SY6Q5V@X)/Z;LZcS:ZYGK
,/L2CBK^(HcHAI5?#>be[0HQ8G#:T)QD\9\0:/[Fd:(1TJCM_<6:;Iff>Q=0E=.?
3gV]1#&aW)^EUBOQW;OgLD:dCNQ\U#Y(:_NMD3f2GR6PZ+0=Rd5M\dOHW.@4cK^Y
)U@1-MDVOF1,;ON1F[d,B_9&0&_ES;BPG=?ac5Z4KE:I7W4V9C:)F3P(<]@&I@Ta
,1Pg\Qad#&W9NF4D@TLY^?A:aU]9SFU_SG&=CX4f@KT03Vdb\b\YD+gBYG4B1cZa
^JQ)3KJHcaH4_J9#b-f\IMKFKfLg]+=)[b(P2\LHXTMe.H]9FO8\O-/X0g.3QJON
bcRD&18Q-gB.B\,][D-<d08ZQ,/+a6B9H/c5WSEZO_A(GgPPdB[;)KBRJ-C2(c?H
OLBDacD3=Y8bU\DG_/<6L#I>dPN68>2I>&Q@TEKQ7=0=YJgO5@=/>=Ra+.PABOb5
+O#ZRD19WfES>(d?_73827.>1YQ)7=e5P;(1;&Y0Ng6,.]Gf3?WAOL\b])L.^.8(
DMbL:YWGW3OFO.bBUB94c(2339D=<6XeGUGI/Z90&XIQ84.E<\))[;D@Z^@Q&Z>S
4C,]I(W2=A6,4X795d,1;?O]E=-XV1.EFRe=/gNe4M3;afCPfH&a,/Eg#eF_WC@(
fVN[FE8<N1T\K]9e=\3Y@fOP/@TMAX.2(^cE[KZ]PT3FB=e5>1SG3EN^9<^YZD@8
ZZ,ZYR6/&\N,@fKK&.1^G/;Oe5&A<]fG=W0HMa9R9c+U;)bfa@^27;TI6E3C59_1
bNJ[A;]F1F&[K=g3HI]V8-6C_dFDAC7X@4\(<If?D0&K?/RJBB.OdVc2:2P,^_#V
C>;_;I1fGR(QJ7>Nb=,_STAd.Xa?Y>VH+#[06Y?E^Q62U]Rg:)Ob+?[_24eb7,1G
#\&U1S,AW7FW&<WB6W2Fc/W8K7L#:S?6#217D]FZ0?3ALN?Db_PNJ>]_Y:Y@UQS<
V:M-/Se6M[9WP.:,EV-K)e7F6(Z)=7(8S&X=)RYFT^S#c.[:1==5[fB#aFXV\LNA
C4bC:dQaD\(a=4GT=JgWO9JHEdB34++bNUfdgeNUOcG7Fa50Q0,_OAg@X58QH_.d
R3()Xe^@+7Sa331/G4e041##K@L,0[-N<JV/3SVO1DY.61CT_LG5Bf,]/@N^>C)2
eWRN+;[X0)CS0#L_UU538F3[+OT8Tc<PPU)WB/D-NWO\S>_V-d05E[WR&2F:83_f
HdWEG.d[73:,D6ND+P21341-eaL4Y52^=K3_,O3dTZ6CW@L_BLb>-[^5X0C&+cgX
<[#7cX<Xg1d<eT,7Waf2#c4Ddb/4XOCBg?CHaJJH@NJ;M<CFJ8(Sd[NV-2gA9P;+
Rf,3Y#M#VEZEUdL]N0&fUM3J0@-14]_X1B(PW0G3+DRFggKN4]=<R[]^2=IT2KfC
-aN?gd5B>)))+9R^;63&&W#Qe?BQ?KZ9BJT00@(24^HNPKf0+)>3fa]D(#FSN9eS
V<NH&Q#Fb8DDMS<#24MW-/@(13LZNERD:Sf83.497V+E5&]NOP,=?cQXXJ9UL@E#
F1;9UNP]C/551LdNK51<IW22e:V#UgD/aeC#cK-JMYcC(S:HZVM<Y6DUTcOd@.UO
&M0cJLO].SIY)BZ.aS2>^K-GV2G//1]8UG,,=4><W9Sc@-2K\_TW1e@Bd:BN]f5K
1AADSGPKZKO/FFZ[LZ8-LI\ROSTGS[d5#B])fC@fGf^6G9=N@2C[Z1&_852A,/DW
Ec1M23SRME.ac01.g?I53SELEL,IcEX&6P?K7bMS-,1N?<=2H0P^CfgO^:0YMIQ;
cY]/0B1OeVc#>,LH8&#6]&TZMF&6;b?fdOPI>#S0XGI?]_:GHQXgAgd9FK&ePg(+
<f^Hc,_SXg&=)Nb(/gLaa]&A.PBD=51[Z@HP8+g?ba2#C8P]ZS,TJe+>_OUYMRO/
2]a-(dZa4=c4+GZYQO<3>84\^E=6#2bOZd,,\XQ4YX?]VM_9FaAB1[LcUN?V)U=e
7gcaOU<0.A)WKQd\[;<#@8-[f&CJR&7\=8BXZ8d87.I9=YW#]a/4YGdgXd0436M(
&GHR6;VBMf0Y/W;NPM1g&NN,TFC72=d=ZMFHbNI#&#6I>J+_JRIG+)QW)a;.aJ&Z
ag[22J1OYSGWbM6f7YJS6S(35e/7[;M?g7_\B[@GFZRD=E:?YT(fQ2^J/.MJ3,FS
8HF>6\A0/^.6(OV_L\SWEKa>g]F9AVa^HN/S]dA6\:=1#UF>=IQgR3_Z<AQYT?CJ
7_O40V>&R(;7GOdG[)&<LE);(8E:E_90.TV458#EQXFBSV.N#(,Q,RfM8dPV-6(@
IK@SeAV;W@P8WW\O(<c0b:37;8CDNf(4KW02(,/7WX&F9P6]bL+]aSN22b.NZ#,c
bZ\MT(^JR\<LeKXfV\eE.\1]Xg[?MdI?H+?<d_SEaW;(Z3LX.]QW\\]\g#6gHTW,
gH,T[5IDe(S\DVJCQ_H7Y<K^CF@b7C<J_K7dCc],FVVX/L(\I7@/1B/=Q>>F763L
-<gg3.42VAQ>,ZcS2_GM:V?-ILc?-XL+8QJdB:gbB13A(@^5+F5IXDKDS9ST,Z4.
=.(27K/f8H+4UJ;^4SD[7(eQBNLUHF/e&-gDQMZUJ.B0:-^SBbg?55H1_.Fb,NG?
1Q]C:FCM]Qf,)(1f,>(;4059+PBS:MbH&cE_YL+?LNH,G0_7P.UE&^]C,PR=(RKQ
_e#0QZT,a>0ce_AA>g06QB:+YK+[X@9&2WQ4:a.bg[SFD,S\[Z]:&.L.#M3NB>-,
I?4E<H>NDEV(+;A#/8(NL&;L>5gBAc^TK,b6P3CfA_7HB&^9)Q9LHbRgNBO7c+N_
8BeI7.Cc<O-?aC5K#GDNQ-JW-I,H?L8=:5bf5/W,-C8)MAd.)d;ABdMGB+R54Q>I
^)J:(<Y[8/U&M/<fc?74@bS+B3cSUfO6T^P[Pe#OgAWZ0fV99BbP3Oa],>_(@XEX
gA2-J/CB5QW5@4c[=.@I]2LE+WdLGe9(TT\e(eI)U_Gg(F=5d&;,64f(]OQ@OeYc
0NI^@NV/#UQ[FSI1@&B1;8Q:gf2B&DR-8)B>YX-0>:9MaY5@SW,/C>[a-,N/PHZZ
W_?+BL<_FM7gFSMbQe^P22FQ<+\&M76V49><W@B3fR-RX(,B,K_7#LNY8JISOgQg
3gSS?@\M1XYa;_@(<5c^Ng,6;.2=NF=XDPUOb/#6CF8T_1/ea/^-8.\YVRJTf>Yb
IQI54_WVYK:#_/.55a\BGf,LK1H,dZ/eHWM4.KD9dfOKD_S(Y0.?14SN@?DM]DC(
I>T9:4b1[0/7P_QI(T-UW-Fb3N4<3_>PXBSd91aT\Na<6D06KZYcTCAKCWW\\d@.
X)Y)T>0_.BO(6C0Z^eWRNb>LL[L+Ya(CX:gX+5E^&^9BA0ZDUIC(Z[=TKD3=g/,,
E>R+LFXDRKY79[^26>Jf,cPINc3&MORICZHVNH_X_>;0&E#E6L+1a?dCYg3]1;cL
+A_A=Ncbe2RUPI(=1)Y:P),Fa=2FdR>f7XGJ9CeESIBK_U^Kg:/G@Xd;C[FO7Z,P
C:a&H5?HaW.J2D=/L:BD2&a3IFGF?/.J,XgI,b?W3g<F99Y#:#eQK#,c[16)&HJ/
RDJ(6^7?#@J)V4CSR2;:?X6Y>/D127M\Yd<g5?IATG[K,N+(d8>b<B\EM0&5^V/9
LMK^:/Q+/e]Lg>=c>Z&c9LV(a.fI7[(M&/]G&DI@Pc)I5-c\X>M20[GFcQ\I>_Z6
S284\U\(I^[,O[5+56>7:=PCB]RH7,[S)W(F,B^fNWU_f7U@7GGdBId7U#HPN4M@
SF4W[P+<;G.1Ab+b68BfNG:>>QaEN3AFc>8a\A;?\\Y2<L:eO2eX#.6\O<Cf10b0
FS^I-bND4+KUPe9WcU]HI9[;F\DFHE]X=ReHZ2UG0=LCLLe1?+.]^,&c5gD+Qg<d
cO7VBZKS>A#Ea=HH[JeG;9K;Sd0F^EL=?GZdAJGB0VR4PX#F9&a+M+SMLUHdCO)6
GDVO^4SDQH90:AKeC0/)#C#cI^aX:f0eP:ZD)gTb^X76c@EDC/.MR6eJY::?E)?G
@5gC:1D\f_gdO2S5<4HEROV#aF5MB,Gb(-@VBcU9+1=XV</IX+8_X6W;_AZ>P:<B
fKd1R2BHLH&L@<U\O02Yd1D-)0dIJ.:PC6M=IbK,/>RM[WG+IK]T3Y2D+WR3<cG(
5H??-de^f8BfVf&I.\619(WGH_N,5_Mg&_JF(_:Zf.XRRGPdDgSS].8,&/QQ1D.F
a3/9NLT;ZA#UQ[@^FFY<::X@H&PPXS@X/R7-8Y3Fd#=N3BcgCMF^+Y<U]c588:eM
^4/R5S#9fJ(-BfS2YA(KSTF6e=//_dQ7]&&]DD?Ze^0_]?.gW0&;gage;@URYMN+
3a#I,6a:1ZZ:QY7W(:\RN/S@5[GP9380^\Fd>VBB^8G\Lc^TKZ0\D4O;E7L0]ZA<
354G^5<gYbHK=KGdCX]+??VKg.I/4CUJ/C0WF82C7f+ZSEZJ-?:/W@<TVVV7c?PV
E/R8WHD,UG3#<5Q1DS#d=Z/\BAMA?^?:,:Ga-Fe&X@Z09IUCQQ.1_G.^<1Y^-S->
M4Q+;F@Me6O>W9cHA_eA@+=SQF?]H2SC,OC423ANf&+V&gE[b28Y<b5f7)V5R+D@
G./^X[G&gFg=@&V8TS8Cea?5;K69TOC97:D(RPQDGdg]ReU<9I=Nf..Y5?S>GNB7
dNR/&Hfc>(494CZQJYL=N)b_YYNfC(7d&6gD>OQ;W4a#Nb:1OG8SI[aFB5[(Rf&G
e..UBE(JfCICNa@=6]GFVADcER.M[ERfd(gBaPT;08.eBGGBCE@=a1Ga&>MOYcZF
+XNgB6\6N36O[6U^CRP1aA7(TF:^NY\dLIbEd8C7-Ud[[VP-.GSJ)CPUPb/^2M=6
8J4?R076VZ[SNQTR7W(aOUBC2XbC_ZTJebcbadX>IPBPbZa?/)#IV@=21/;;@H<2
^_&Q(UIC3\/2@b3;-KJ3e[,LJ&T:;c?6A/5Eb-,e;dGaQ2f\+A],Z[-45Z(>150X
KM2R.DU#cHYBZ]/2_6gS>9H8LQ,2>2;e7;CQKX[I(\e0HG=gMQAcC)5P(?V[]FeU
T8Q..7RY.Ve^CaOBX>:cR]c.6@a7AVBTcB]=O>Z+1<#X79RXB3)S;NO/Kd91CZTA
TV4H.a>4LG_XY&7XUX657P9X0B9c<Oc,I<cPeEd?G[XLTF;Qg@[W3aLDXV4HZc:Q
>B0<VB&fECN&0]GACR\Wc16;/6NfPE:9&>BTO34fLgL[?b;5>JBaCQGX/6DR>72/
a=(GTDRO<4QQ^)8PW,_R\WWcb6DO[F9I.]>,b[AW1HdD-g;@eT9DM1U_EKS5&M6;
XgO^.3)\f]\&6X6&#EH#):fBH:)Y(C>(Z<G=f)fUZV0_\efB\4HX0EbPa[DUS6G3
+ReMgI2ZCg8b)8])-U?XBDD2.0(.6SbOTd15Ga[gZY^^edE>UO,TSd1Q@]SLSE:I
/gR(KC98Q#:>C7FI?L]:D.P8/C:aK9MNE+fdM[:CW2F^M4#ff)gX6X@E^SS4#2/[
VAY-fEM@TVW54&PNCG^RK:,+9788XHAO/2b2=0C;D]4<gJ32G,W7U=GHd)6?SO2f
RbPSGbZJE7SWK=9/GY.X<g>/7=KWG,NQK)N)Kg1cFSd#SLe.>Q8OWHdV[gT0SENV
_IX\][W&8DCXDSZ2JYU8c<):)B?9eV,S#@faGfADM)]6GP?I.D\R8FJ3P6FF#M\^
9HE_g=[[._DLMTINDX+7OEW>-DX<;DIaQYK&QAKP58XB)Z@X[-3C1gF1,LXeCWSe
?<^eS>OV&=3AMUF^U7XOXBYb07,f(2:EZH@VLL_N[KeY3[&VR.Y[J4XPI2EPZd>9
YT]:N9Lg@Z6B@_?+)&(d-eJT5/R4)3387B<b4BR/B4+YXX6OZQ)g07JJH.>ASH^f
28K>V-..[=VVc?gcPLe6[JYSJ&9;FBG2&O.0HH[LD32L4)#gVCf4M^J)H^:/Z4Jc
5AU)M41>X[Jf2];:PO18>TJF\.F8aB5T(_3V@@@K)HQ[=_a@T@3_eGB)>>;W9<(-
J;=1:,YK+=CG9aC;,<HT>T;W4TgXQ6CX)cU,a9IGN?<\_J94@HSf[g(ZD9Z4UgY;
[@=@ANgX@VJOd0Dc8#>0O[/:5)/_RNZC9Y:E5b^H@dBDYRfT?.^fW9T&0bd<?Y6c
@PXH,<^/T37+J-_3cV2W7<Y#Z<cQK^5fJU9/1NIe1MDLNJaF\S(7:>MAI39GE^eJ
ag>4@KaRPa1Q51K6<EUAWHL7+BfdQX)7+=X]9?C<#F4I+5c&3eME<K+JT#^8b8a_
f4f15/g395<@.8T>,\#]SXHO\7-a;S]YIM>eFd3OT(2H0.138P;Af7-1)gS4bF72
_.JCA-:X&WX8##bOaEB]f4(bHS)V)e>+KcC^A(UD.PAJ@6U-;5>^3)55^?W(QRVc
C4CRZJ+JU/6^69:IV/>UI@;CKFHDHZ7C89,?-K_cK=I@=PJ.M7-S@#SbMZO,R;-S
=L4J9?STEaA6AfY>7dD@8_IF0TD199<b>)&:Yf8H;3PFEdK;dA;ef]#=TTULcC,]
c/?<UBOPYZG+bJ4-IK^;Mb@Q+/2C\J.<b(WRe6CdIZ(:_#e+Z6Z>2c83bLgMCMb[
FENNd=DE+CSFfN]@N-XP=B74#?(_CB_:?KBBWMfHFDMeVOO2.]D7IV5MA6V_gZNZ
P>DL2\MXZCJ7;LAIX=,T7P[U_(-DC+ZCg>Z-&4SX)=ZNgR@1?SL_b&c:AJ4c#7@c
dZ))A/:(Eb(WQ69I3^)<fU\1>c3M\NX6N9Jf6<1=aaX<A6a/IJd;N?GNKAN3TN]d
;?7,+W&N:<d;X-L2-6D7P0YBU<3I=[(BJ0>11=Q3(c<PF0&B4U9-M-[>Z;Ac^,9D
fN/HVQVgO7EfE/c+.JL:=(KWd]4Q@WRTNg3[3T6/e.Z1[,\DUK-eO1Z3=WA;BeLX
HLTSH2^Cgg5V/#2=eUG>>-QCI.#>D@JeC0;^&MM:FeIKM>AERbD4MW1]8HMb;BbH
4beGHU-MARN&&?McG&^):XMD1=LO=5JL:f6QN)ZPCe:WT@?N;J<6SSe5_^e<0G12
]0,gCBY8IKM[F<R&1d#+?5T-&:+0[T;H#B[TAe(e-Dc-f9Wf@Y<[Zd,TMY__SL]O
a6ML_&G)=^)-83\4/N0^K#Bb20L#+<],O_:cTDHc@X?WT//.&T]YHQ;d3MaBP_DQ
\GH>0Z=\K]S.:D.)aaa41+gY\I;GI7G95/cZ5-U8\QMD+U(KgRe(PRVDJSf5G=UP
?^bg&/?+ONcG)AO#OKJ^Ta6;1<)T+N>Sf4&H;SUF1<_TC9_\07]A:B[.@3f+3A7S
I,cF?77JE#T4)3d[IN>U2HSASZ5b6e-M+Xe2@)7fRVI)/.)<,+^H#&4@J5X(\39-
X/^^@3>#JdTL;ObQF\EeYP^0I-XR(&fC^9aVB\<ZLK4f.2W7#?_208S>XO28\6P&
>DUd@&N>:W.dOa15gWc=A=1BM4GF@Z+JJB-FHRXAb;;f@L(/0]3T5TBdc2763DTX
VH1T.<e?@(F/&bT6?-.gM067==0-Z=DI&EQX<NAT)&PgJ6<ZC)L.0Y6K4&HQB-YR
7;<gE47U0:O@@FMEXZ^gXZIdPe)/8:J=YXNMf)[&;(E2KE5E,dGIAUV,F5YYZ/^@
]3dbYC]b?&UeNR,SL4-(gXQOJ[1a)1H#_gL:]bM^M7=G<_+TVZ^_1b,dT.#OA2Vb
-=Eb._fT:e-J/YB5H??ZA0,We3W4:Qge6BS=E?82/a14aTdF]g#fKNRdTU2DG-6+
J;D\W=ARLJDTKI[\_3S\7SA4T(RIH<HV#K]C2Xa9JP)]8\3((XF7J#619\,g[6g4
V4N+#2VW&[&IBDKI\7)LONTW:0Gf8P>H)#8VfFSV]a7P^6RXc-NfPKJ2.?;&W4VR
cUW.[EaG#4:0E<R@ge;3#\O56aNHaMJOe4V/]K3]gFEG&W.;MQA2#13-U2.I@-gY
0>/d]-&GQ4;XdR@B/-MQ93.L@1cRWG>)Mb;T,PV?X4feO/@,M3S&e9.Vfce>\:-Y
8Zc.<&0>6IQ/A8:UPeQc2-LMU@^P/6IF6YS\d,+H:Y/VA)11<d#5IP&KI,06(CI,
T&LR1b6C6ZFYQ3]cR=dedb3Fb+@ONTM.+?IEb\=P8[OP]PfJX;2S=a29&[&d5Uf.
_Z1W,VKbL]./;Z[-cXKTTR[E^3N]dMeFRB-,0EIV-5NNSK5)10CbGIL:+2#41(BM
CZGEMN=VPZe1O94.1e:-3C07Lcd.^K-Z6#K@Ob:=X8DM>1#6LDDGX[6G[]+d?_LT
Ud-Q5Y8^I3KC.P]#GQA8:c^bYNT=4E<ZcJK/e4JAc]cF)dS,V_>VBO6DIDCS/RF(
YO?F#;-FTf/-]?Bca^:HcT+1AKMI^dL05L=fTJf)JXHF<XI:[9A49K,1:Xe?aX[A
&;;L6LY[,>FV?cP^=]./8W#[B/;5-R4^&)IVE@@fU\CO>>-LgcBe4VG.fK(Ab+X.
&.SBbP>85IH8GTR6IO787\.[:4Y=\+K=U#Z:A\_)/\=^02#QTRM,R)EZ,a\E/>-Y
J+AbEGf[\=Z=ETJa,eYCfgABf4UY2Q/+H\BaecA>&F(d(>:BL:9]^S(bP8/d_##e
[g3/O11QM)1JZc1P\d+A2fN>MBR)O^[T0.AMF?G[[eBW.9FWU+M>9FdgJc2W2&bc
NO3)J(g+f8e-5AU9X-1A7B^dAD--99ZfZA@bCL<.O?_N@1]I-5HETFRV@8](>A)Y
K72]JB@QK/Q1Ud.&LZA-XVWPV?M-UTeXF(A_=c3cT9K8_5;e7L6XD+#d21RR]>/O
(Vb(YAY55T1K9#eYR0JS)RQ9;GUaC1gBY:24eO#[Ef\,J&N/;TTI:5XE^8M[=J)Z
e]5b+W9?-fRW@DCOEEQYCf_&I#OQ5f7&=dL+WL]V+ST&U==eKJ5F7cJ)G[F901Y_
+_JE427DQV1P#C:?ZM[7[.=I8Q=BaUIb:^>I]]0:LeV-BL+_T,YYJ?Z7Y]>72)<5
PNPA:K&F8=0Q;VZ,/8SWe@1:W+L6bX+RVM-_I35;QR\:GD#f[,-8SE,/(XBBeTHK
CBF^Kg2X<QJ8#2XSH)SKQL-H+F/W1^.Z+X-H1)+[6ICgJOVU;:U]L3D1EUa3bbP9
deHM=A\,MF5;0)ZY^cTGE2feM=+W@F<T^1b<C.2gS<=_04V?5EE)B^7+g/BG[HI4
+2]JYc(+9J;^>584:c]H.Ub#?-dNeT4/U+SK3K7()NOb+MHKbE@X:f\O3/LX:<8B
5dJ)\\99L&0;\KARCf)gAON2Y-UCc:(Y+^-A;fA&Qa6Sc-Nb8HMZJH6]d^_+S0fY
HZEeC;BL?/&,C/NOIb^RAg2_1#^^&WP3eI=\^@9ZY8F18W#[GR2^6JK(c&0fSQP3
fHTY2UV77ZD>#Rb>VCX<?6gAUFK.#XaKM#)#([6ARee=C[J4@L@T>T1R;55@ea:/
L>8P;SSMN+aD_fJ;f3OK5ce>^N9-b6[I&6J#cD^4R^g5#4+K?+D6X8(]8_+L+BQ:
d5FLAGN3/,Z\Kf,Y)A5)+F68WD[T0A1W2J0E[6J:.f,(D+;)XTTT>]dDOS>d1RNa
Q+9V6_Zg.C?G-4DP\a>3?=??-B<+#6;Uf8\<dW3;@5WQTTLAAS=7(cD#4bA;BccG
]#2H=FFPC=+XU,/Q#4T9Pc/,fX@AZ)/c)6Z,58(3=CFX)9/+Be:^6,e.7+G@:CT&
/SB>^770KC-Wb#R\GG4;cW)E2YS7V6VJLVc(HNd>FeMe8EYQ1<N)RJYQ12YO0e-L
8/)8)1;D:P)e8JGJQO=Ge2X,^/CTS\^>=^R2RZTU9^#e7C+/N+Jf)GP?TR@PUKg(
S3E+De^7^\7]YaOI?Rb74d)W:gIIQ^P6Cb\]gLW-=\2c/=DSZR_gT,K\Q_cH:IH4
B75XAAI+0YOK,d(f6XH?8KG;V66b8beUWKE&,_Uf8K1=97f0AX(151QQ\JA\Dbc5
dG,a0=56?3fb3MN2+/MOMIDSae9-X_M#R<A0B7UGBCE,.)a(;Xa9CY<c_:JKBEZ3
B0<CXEaB)_&X]&+@dbCBa3N#dYYPAc_=MaD<0U#<Td.F?(A#URM_9eJ-Q_W@)gQ3
ZJL(UM#DJZON2S,=.a:T)D0QYc&4#d]C0eQ7D>gNXd.fa&,3?@IgWd1&&?[Q&RT(
/9cZ1;8BZ&L<TSTIN[VAE+3/cQ-UIg,\\C)XQFHAdW5Y(Hd5CC#Pbd]SFKe8^/-=
;BP),4HC1YU&]Y7-Z;TP(O&<E9-598+)f:)[4Xd^>:DR[FVe)/_OV8;Aa#G;K0=g
\B_ec^.FQ;S[f&,J8:81ff]Jg(9^7L0@=Q:<O(B(0?]@O&EOg#EGE_g-ag3-8+OY
)@ed,A4Kb2>SW@IWD]Y>Qg(If2f]A2<B_Z@N7YO#8MD8>)VO:BO<@SB;LO].HB+W
#Y)V5RDgH?3\Eg.GYK/;WKG_ANN[fbZ_2Df/e/AGQ0<.A_)FV.@e?S&CYgE(<6B-
a)UEUK?c5X2M^N(9Uf.-(\ATWb4I8MR_H9A=X\cLW#b:[;D\1;HKVZ5[OOL)FQ]]
a)N;UN8KMP46LbC8ZA540dbKCCWC>)7Pf>8P3E)6HP?0I?52RF]T<^8[gL7:V:IM
J;ZYWN(6_:68462M61^<DB(:0\VNSgKQ)=P9(;&;XA9Ze8ZO#de]#VL=W;(MO>c\
WU-@eD@-bV7RTDM06:,;>/C;gR-dKf(D(VMI2EGKe82Y#f0WXcbPX[_(CHIB9gY5
@,F3a.S]MB<56ZK/M@@YDRKb:JHUG2IF04-A=(ZIU9QX#4Ea1<c])cCK>eD-GMZJ
ceDYI78>HYT]gbVVE]8)\^gO@-7S55DR,]H1GIfg?)C9IG/]5AD)C3Hb[BX[MPg6
FKQ=[R.@GOBdUW.(>_BTN:GXN;0.R)VaV6RH+^X?(/gG)gKA;W#c+L6^,4eU57c9
+9GQdD\V2/6[EEE6(]J:^6-]CVAPZ<GUHP=&PVB?:&311CN:&7+_AORMU@6DQQ,K
XL\(9ZP#7ALFffDVQTGU7f(S>1QN:,D5/agY-J.2070Q;:J,MdDcG.aADI=KS-a?
b0CT5L<@XZa^QB/5.AM4bMMEVV3H7HT:(4WCVJ1,&,d7d,)9B09A+G8MWb-64YU6
d:>YY#ENUYQYRS4;5BZ-,FQL6CR;CeJ>CTDY/A3EWM-#FE@QPE\KNCTd@L^HV6<T
R0\<UXg\R&S3DZgD7dZCV&d12UXgUUJAN#?J6d./W)V:g>Za5=O_d>;.>/MB\=O,
CcYJW2J,&+A-:36U#cD,0g&\2I_C+.I^/OG)L+4S-5_.J[NaI[(a?IJG^SA>+@aP
I=#)e<BccN7&-+g<RAYbfCa#d>V.O<^H2/B-VU.8D7SM/5C63^?\&9EQXf-CC&RH
/,CV/d=#aI34O\3A^-g,P/UQ^-WW#2\8e))RWX0MVfQ9[Q@:3&43B?]gW<&/&DFK
fYTORH7K-JfE^Y)P[)^/?+:6YG(BYX3,IP:5Vdda4Cc1.SN+2=1\b[7I<WMH\64Y
:)Qb:V:^3J/U/J7GW1;4O?e22U92??Fd4.>).1\98D\Ob@ecQ]LB_0VYAL5LFMXc
:ESJJ(J/[7Q\MJ)g.^#HQYa,GU^C)CA,X:bPaF.&<.J(4BdKWZ4eZZ(RZSYDc8_-
D7R.[SaD/QS(\_DUB;<9bbJab3U_g=c[09Odg#+_FQgWXGIDFK,46]8-f/,b9gGU
>N,^)NM^MIe.6fLY&AS23UICX\<d[f=bO@PY0)0gW#Zac@LK/VVJEH+_+ISf),(>
eIJA5)H<128\PD#aR9<:T_)S^AREF?F.98cAXCUI.efK^(J@Z3AdDW(<SPJ@,(E(
2#[@,S5MFa-<H2[5@(a3TH:8A./gB_Y.b)a.H_72HR4K2dDf?5PGJU8\>facIMY;
I:^cA]4MQ4J?@59+6)XMXa)D=(SW#+M::9EK[Z=:=:GeO;X<7>FLBS<@W(4N<N/f
G\(>;8gJY/V;LMWSg5/26\OVQPgc&LD7Q)-><g\VYP<ZdVb7>f_FAR=8d2:g7I[B
]Ae9CDIO]N0_4=G\f+fd7d)Med9[FZ5:\J2U4cJ2<\gEYROLM8?g7=\#5)4:FMD>
T+3HMg6<dK&L,BFR:9/(HSegN9N5c1ZK^b1[d>G98ScPQB^KbUZH7Z0?gFSFVMOT
<:6BD^fWVPJ41a=,:#4+[-CB^VQ&6(+9:GP5;e89Xf@WK2J-ed1]<G\&-3_K:(6J
T5Y<.SKgS]YGQ9cgFKG<&,KKFa@Ce::JMM(NaXS:ZE9J+1+41cZ7TOIGYF9I-Q+X
f:/?+dbNDZGBQe):<YUKPH^[<6[/#@Zc/<_)Z1)HF&ZYVH>24^#VNR3=B/=aTRSR
c><#dba\,0G9VbbCeS9?\&,@+CF[G+HI20X7X]-Y\+E>3+FRSQ+Yc.]<EFU8MVdE
+EI@]AfS3?b?OPRVU9de,5&2EAV0,.5/H)Q3Q;.PB)\<IIU)TaDf(bDC85DQFK=R
0Y]SG\F-R_B)9@.;F#5BcbE9.KaacZ5O>J)4B++Q9/9THcPNNI2,P1Cg-7</OgR(
TaM@P<#<0E6/D3PO#=9YH[9[/[<^JEZe+228.M[;A]_9A1\@g^J+6g/TJcPB61O<
b8;@(dW&:,LE1^QWQ&Zc=JZd2]\UFVG))72>&A\<ZR:fTJ#Z2OWM_B;]X4/>/FOR
g_bO>ZK=Y.QWOPc)\cT\3B5X(49a):[\fU_&Y/.YZd,U&-=A?b;/8&bA&E0;<^HQ
RGR=CI:0J3#c_S\M5P3/>ccCQfY8c&>[\47<Wa26&MUCeZ>gT_/14bVYL@/,ZOB[
c9E6#Gf5bcK:0[[^dSZ.P3S+aUga#8-aCUT(V\]dbJSD@TNOXa3,V^:Z_\&1Eg8(
Hb==,DKaO8(Eb#LX:45Xe>6daOP.YHRML&-;a;W/WdUDVLB>A59YC#6bDaa3FH(G
O-I/8\HP0\f[f/1g7X:UEUPbK&,_Ug<J3W]N.0.@4V#Oc-BTa4H187&Y?,C.:d)#
IBE](MQ_^5MD,dJW.a(X1,/F1+B;2+.\J/6b.7C0d4)Hg5N.aG?g]dGU7DA-62Xg
XJ0;[S]&1#NQ\N8GZ>PL#T;Y4JTDJGfFYXM[<B][?L_;@cFQ3Oea5R9(W6S_;Ka8
PPAI4IB#C0:bMX59EG6=gE@J:Q:P5^dbfdB[Fg#.UE#K7+0J5-BX+ITd92XF1RGU
2F<ddTL@&bPa<M1::g<C#NJ>#F:+DAe0S,VQ#ec2BP?)Aga9Kb\T0-YMQ3/ObM_K
Y\73\eIg7C7]&():V<Y]?FLU=>9OG;e+fVM_GYcH/b89d;KP.RL4E1OI052+-WRB
KQ?<APd#e?1d7J]c9+DGJDU7M1?3G1H@P]3QZIX7Q//e9&@4e+C(#Q]QV1>G+aYU
fcI(_CLBB7e6CIT?/+g&MC<SfLCCEM<ISFGQ:D/R51XJO5aP9<)6g]N.,c=[T9LT
U?&H6T-;2TGE/VF]N39ZdF[X)>/5#6[T>M+.Wa,-KHPO?:++#WP\dL/-Q:,S(]HF
-KdN).L1VFdMa:9&7ffT)P0;4/>>(SbR/7TXD=fX9H<C77O=N)M9^HZL=a;V7I\c
.R=>Q?I()L,UF#X3PC8gNgc\1=/RbQK<9bT+SJ@_#^eb_^Udb5Y[fF._^[)0Cd(/
QN61+4\g,M1eeT#;BYDFU98_EDLA^9ZSP6SF/5ZC&7Ze#:AW3#gNMW3SOTI0GI>;
\]N3^F<>ECS(Z>[IeQQ:J6F_<\8_a3X3b=Q\JL03b0;HEd3+YLV8@,)-_c[QYS2V
=UIK^N#cMGH):X:PPFBS,KNK:.2&Ra6ZO_IEK/\PO74-XBVP1Y(XEP+=^=7[=T@Y
??@W20e-^6Zg,K7\eDeT7baSaeLb2-RaB-4Y(c3B?deH\@CY^+bI\_X>CaA@<OO^
ed^6[/MDTH-FZ7DDD0K^A^]b7XI[b<<,b^0c-ceF6X2H?-OQSAN60#=11V^0UUQR
SA&,_Q-2:P,R.HK5g/ec0S_1&dYObK;1:cN.Df@Mg)\]2_]>J;#gLcG8ec2UDgTH
/L()dSNYW4Y(;Z0OGc>EW;(&KTV&g=I0I\QC-K?SUQ-d&=KFWe@I]^]50S/-98cO
DA7:4a>QO17g:9BHB-)ag=H-(NYc#:ONb([MXDbD5fSFWA5<:3ZZYM=K2IZ2?<6K
&(5#MPNMG-3Y5,bK#H10=fYEbI<EXSOZBJHN0e(]bTUUOf)a57#;-RG/1YQPG19A
8V_^02XTQ=]Y&LM<535Oc.d:C_R9T5.&Dg&.N#=E-.J(O)aB&<@(UJ5bEJE,5<b[
aBf,]5Qf/@#963/)>HY.ZHSGTQ_A:L)6P;cbRd\9HYET@dG,ISQ6GLO.8LQ+G0\.
4TPP+,=#2V(O=GRL9G@7#/)#@TJ5,,P4YG^Wc&c5J3=TeFGI;a0Kg2O.N$
`endprotected


`endif // GUARD_SVT_APB_MASTER_AGENT_SV

