
`ifndef GUARD_SVT_AXI_SYSTEM_COMMON_SV
`define GUARD_SVT_AXI_SYSTEM_COMMON_SV


`include "svt_axi_defines.svi"

`ifndef SVT_AMBA_MAX_ADDR_WIDTH
  `define SVT_AMBA_MAX_ADDR_WIDTH `SVT_AXI_MAX_ADDR_WIDTH
 `endif

//`define _SVT_AXI_TEMP_DEBUG_MSASSOC
//`define _SVT_AXI_TEMP_DEBUG_MSASSOC_L1
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Jbv5ns5uIqspCnP/c5jJHemKy8+DGrvWod9IMtKGAoUIUvhp1+c2Fj9DyTrbiggT
A1PRPe5KmtSuMpb23VAS1j/SAO54N2ipPwJ9ew5imRjno0Ip6GrL8eojiraT1VjX
q65IlNQVat191D1F9l94iqFqfDfAjYwNzVNUVtknIW0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 10688     )
Y8s/Auy6+5aGWOvC/7dp0KJZTG2SWb0Oel/QxqGSe4gsxMX59TNr0cx2bv5djdm9
B8sBe4QTO49DCfGlyaRh3b7P1sATOeCR7coQnf46p/u+oAxfQ01xuWQgaGwIUpQ4
NINCi2MIkOzoR4RBbsP7NM3GnSM8jypzjCIIpXpXMour/vsgosYSiv1+trC5moN7
C6X8SU5UJ8n1XbgPFuKM291ZNPYwdz4TAK0opnLhAYJI8hqUXMTKXjngxNUGom5j
yGLG387rhtAF/pdL2ZtUProDMjqFkiHRTw7M9QXdFCwFTsBMoft9cIqwWPxb/6UT
QIFgNKmIT7Kq8V78Y+M1chcLlVrEx6ai7rZtdNTVRM6GhmkEBq2Xx+VPhtm/G3p3
FUzNms6pwGGGbx9k2LmTfUjsDtAe4AOki/g8STn2SihoZ4flXXxVZcrZdZz+YqnE
3fK1i2xGQsAKsZIRmksAgGxiDLJjj1Lxs2R8xkkE749GYY11SRDsRdVYSOYRL+p0
AN2sW6dRVALfyfiAV6rVK2X0Ha7La+o+I1/IeVucUxkvwphKb02fczz5fM8QTWne
DeH8hnx9jMp+vH/WTnT8DDBDcUS5htFLZ3xeWyW13HydvFCTfo6bAw8OgUcKnVaM
MvM7DuOV+HKWS2s3G2hHECk57wa2vfS8HH1XXkWketCFG4V0aYqQHmKvrSW8WH5w
nGEx14CFcUOR821K5Wc6SmpHm6ba+3fLntrlBgnMbEI45P4xjDiIYHEJm27VAmIl
ftxP+xoFP/FMugyjk7LiZZARqwakDaziI6ZQWZLGu/96YDj1d8BVmtHGAGV1kPAy
e+Fjays626/X3DkcILxFFj9PMsl97QYwMFbwTolIWFdy6UiNFYkSz9mP+0TeCx+O
JLsIdaKFSrxPqMEzS0HrN/0hFkVdcOVCrK6NOdaqnOKHhFckvfBnVFufI86e8oUT
Nuk9ddoZGxU5Vua9FOABmq5IggtxWFwe+oWMZel0E2XqNaVG77XOuVBI0F937xg5
ZeCTg2u4jHMJE8eWCHQERnJzK+xdFnA3d8+31UmAtlAwZxCdxy01xaFRMpi3J1rG
va7OCpbrFVEnV860Uh1mRkIPED22wx5zbz0Le6vAvURi8oiG4je7YiFGqusl6W/g
1GXYa0mxdgsXhGhUm89cU7eNDcamGpXZnPU0mUYRgB+i7aQqKTv7ZGi9YIV5uHxC
G0Q9EslTB+iwt/8wQogAOxnCdGO7rp9KaF0ISofE6f+fKx5QU43OKRtz7OrNy5Pe
8TMyWFVQ9UjO/cv15AnVmVmEQgdZZQl3Fc8XQ2MozgJWxSa8pko+QebZCLSph3Oc
XoZkNWNlcSNDVlgLwywX5iGyi9fIC1N+qNaT0cOPero5SFgHQzL0zZnmmpsOljKn
oEgfmCyrx30dgUGnxfrdpu2IEyln4GdmMcnABtAEDGI7OgmyruYFhXQpXgJu6Lr7
cbqN9y9W5EdaD6RubQnbj7wJLEZfwLSibEljMfZdbiYNEQhctpAgNF6aXFy+QnaA
zHmFGURXxOjUY8KYedk2UV8dQTNafPK2iBnUqG8Tpwgd7Hy8UlMWcrOHhDvDYtbE
mvk7N7aB/Ok284IHfFzUJa0v88U2IL6RD9jExC41sY3/gFdtrakdZWsbcyM5vS5G
h5yYxMEpjPb+RKb7RAt6lyQV1D5HZZ39j6rWbbDQ33vMXFLz9smw/Qs7JsQ/6PrF
RIHKosATPfDok7pff8TzEnBj2WhOgWJNznIF2V1qOojO6GwOkudbn0DnEjdlcdv5
Z/zU6XOr/bHJElveWLTey4UQAS9i6zoMY93x3ubqaU8FKgVqXX23Vskej0f4m2LO
O00QQouNp6/HAoB1jZ9yaYkjChmtMXKtAR1WDdaPjjdykQrHOgFVC1bHZBjcI+c0
6nxtuMYvPeYkp9LytOLvIqVRFT+AT4s8pJT3F40csGhmL/FE3dhD2TVAhj/qlTVh
+dDV5W4d0vIDCY0pTeTyUIj3YhJnIFB/wths4XQ2Ui9smdwcliqOtzkBWBi6Jnb+
Y04hiXN570Grh/fyzbdQn0NBwVhNDE8zOO4g7oTFoZBR4YsHWsilq/ljU9Qv60H9
XFXqyy5At4F6r3GEigpwfbDZxuz5ZxKL5Mdor8L0zq/7/dRsR6Y/GgH7kUgFJVYS
xqfq4tOkHkPwe1ETjk+G6cbUE6xbvA7V3bwaQvEGb23qYRH3WZTXqkg/H9rvM9le
my9VCPMy/gJgC0sEiyIeXVmIZl8kzayGg6tvUB7A+RYqrflQHFsHZMozbl+mZpUS
qz3D+DMZZ3UjBL/HPR3B2yMcjdlUpnNYa5jHLOrLYCKQMhM7V4mEKXGSOra1qWFf
qsfoRtvaJx4APrFExTEbBjdos8Au62lk2oHCxCU5PhvbV7tf7IsjmDQRvk9jFAg5
IdUSzL9Zc2howitcZcJxQvXT2OVz88ZNJt67KAzT6smViEstgoD+DVqxY49KGtog
JGTJLL3CcZdeAEhKYcghAnq1p4bG3ws/paFzeHU9FgBwjEA+0XaK7we7Jw7VhkRB
XdICckvzK6DM0Wt9VI45wu/T47e+jXcmWPgI+LreS2AlXBMmL9tfY1Ea64mVaRMW
1ojsY+s4vw/xAK/WJ1OUGvJw57EXn91Rlx/7zwF3XI6xZT2K01U5sq8cCVUmBZgb
aYK1Qe8eyEF6SxqXBuwlgZAQVbaEa05F98GGwf9JqfbiCQB/zPLxsDY5zACpMt/q
bv3BpsQB0keVPJH3XQ1Huh3/rHC4Z4h5NcBZOGmoGQ+EkBqyprrtBp5/NWDAUexI
ueWa2gI4mMCDiYwYGcKwI5D0sCDDm1KkPKWkSlIe29C36EeuHySmEeE/Trji7o2U
GFYiQKe/wj4PmpLSd9moP2xf4XIAZsLrTiNM1DR3bcpk5Rl7PnSIJBFXXIVk2d0o
Y1hHjEIfBdR+xyVEwzbfUOSaiNwRN2Co8h0CxtGapw2m7YkCjG8CF2/FvnajQXAm
UFHpdBuTGOVo0hkPq35ugOryQVt09GWpl1L+Nlz0LvU1VfXc4p7YJlIxXqAG5FVe
k9pVXh/IHWcSrIz5LuUxXmSic+gHSfwKqmgtAnpqgKuuPsKlMjToVdvzXr+deONA
nHldTfK/7wqMciZpaU2gRE7VZb2x51Y4EYP4PLVCMTaxIBWHNL3LAhzbBMtr3dvz
wN07xJL77lcHTx4SgIiLWL0dJyBF4ZpKQGGE476bDX51AEwYnTcjQZRL63d0xNC7
Iiex0ULK8ykcofJlgIdldf9Y2lIVaCeN1EoTchgakLArJWwmhpvtow0FjfldVYMi
RxxT+k5iTtSv1cWo4ZJvw0dmvOEGvRpeifWvl5srOOFzlQQqNRDoBYTTqjhT+Bnv
Qc5ENnhGa8f3xLyxQCSUB+KUhFYxXJ6wZkjA3LYaz9xXxPUoIlLPBZ1wJps3uXLl
gQmRTi9KRAqndNHNn1V0jCiJYoQb7Y+4F4n76Ov0BVmhrJ+tQbboR0VZQxEX96OE
IWy5fYXMvOA839jZ+my44pO64OZDAszjDi7KFTQuBM2A2OBq0RNGF1jniPcz0V08
d3b30uSiImJBIZKvAJOUP5ftobEgzalra5Q7IQpvNgefCGCAP10diiQNgnOmQXnu
WhBc89nXnmk36/NQ8eKyGNDQzHFWkyZSFYshYZwuzoYR9Rc6jMLbLBR0bI0v3hcF
nCDEtbtvyxAGpix2jrAxm+LDsOoONhHelpM5DqHNVcod59SdF0cJMP3zs/zNgLKK
GnCiDIVx77mn5ctkFqTpPZ6JEGPmks92Z1wdM7s+pAOiYvIb2/rlOjLKbdHAGwq7
FaaSt49tUOnxhaCU6h57Vw2WbBPo2fOxpgH6ES+C/ee1ZK+eiYOa7JlvFiq+BYHY
Ujh7VNXydZX5s1yU+PNuIAllQ9ut/8zi7+iTbjbyEjVFSTSWNjJS9y1Xa5rSapXY
oKFP4AeidcDh91LFcCMNvi4KM/90gTF8ZffPG4e2yX3XVtZe+b3UFSTIPGz8/RdO
gfINARRH47woHjk9DXpoGK8yFvTp6HWs/kjq/fZzrkCgwTzlBeAmELPQMf+yZ2Ou
8aq55Vht8DjJnp1Vspnuffr0w4rtQPwVYsU9UZn6WQ8RCoRRdg5eTqgxui0wPus0
KlP7bchPNwrqV2kQkCT22b3BtESopmnDHOcQV2pgtbXFk8ofN2q85arTLERwemmN
Cjh7nCmcAuLqhsI15RfX0gllfC+wqtDC/jtxE+Vn6fthVgNamBrIfawoFG0QqGEb
mqhcUd56hmhzIZWe/8u/NAjQ1bq+dz++4qWvLeI0UK46aOIULCSbluFTieIhmreM
3nDuffRKdlrHnGWsRT7agTkTJTUGpklKVZdd6nxazw70UpNymMCCEVP8XTiT0Qu9
a+rUIUxnJb6OVEGK51vFkWvSwrKVtqpJ4awMRa46cI08ZFjeSOCQ5vCnrFR9yeDK
5+TA/4Qr3Ptb/mrCLtUeSabu0UTmUz1PnCIlVZclKwRDT4PFTgi/v54vfoIH6X4P
9iAuEgoMg6WSsdyCpaogRDSichN5DPKkdokUmHKUreXZtLAZF/AXC0ozCZVazpD6
prfb4Km0XnZVoVaih4rkymxHmUY2Ry+c7Ab+UT8ctb/POzirpC9N6ybatq1HTa0v
xdzpObSOr5Ax7GbDm8JoTcH0AWg9+/CNhRo6y8U3ZGWuftBfFgRPZoJkvC/d2wa8
aa24bCTVpratabYH7TQc9V/xSNefA8DSJR1y/CeR5ijamIjpNg8FmBE+tOkJL2sA
TOBEIpm9iX7zCHfjTVB95v4pix/E6vhxDsFuxUFm+S2HOSdhn5u4JiEZmFfd6HJV
NSowZ4qryVcZb+NleNjXFNkLRzaAbVVgZ6ZY9WhVBodbwTScidHxto+84ptIkl9e
if8su6idHAn8OLmylnzPjG2wkfEGDJkZD53BelIgPT8XiZgLxhwoY73nVUdxxgKu
+4w1k/usemNpNM7DbWUliticZsQ4N4X5sJY5aNXtZ0f1iSkSGutIqQP1/UCMmaQH
LMgymRIfgJt+/+WDgXOLsWGDmuZEawImia0yO2mOQOuLsmXOvjRVqNuU71OEyzil
cZpnsqZpo67adJnKk2Uwca7Xyvt2hQP+r1hoaFzwZFT28LdkzsAj3kpnfylPBMC+
JDlNHy9iwacSmI+MQs+8caI6E0NHYu4CRsJE+13U2IbP6JIs41CB+K+9xDB/ZcFM
3rHH6Ss7KPweurOnLW9sdfZTITeacS1hoqABqHvquftQbOxk2KRLrs7QmQW9G2/8
7BR4HKmM1VcDL7HoU7oLtBM1zLMjjClr0A3BkwJQlENmLrAJqFNt1ss3TtaMLmNi
kdeeJ+p1WK4amhkrPn6qHUyaXj3TUCfmJewrgSXqB8LTjrSwhoSs/1ybeoOTJxqh
SXyBUarwj7LO3eXM7KbenKp8cfKciKhs7mMGiZ6Svjn13jyX+GPRFGYYJTqhhb9q
BN7UVX3E30SJRkMECpUJW5rXnxkf7sP6JV4vEF4sNYaYNdGT3ETEGRZmeATaCzOb
oc2J8+NVl3DdxeenwOFBUILXMQXSKzEdmPuBY8WfDdVQkb5jEJ8TgnyJMxALv+xQ
IGSMM5aAxhdV1HP41VHwAvy+cuJ5VYalYcz6bhGj9hGlDifr0NqssA/7HZrqhG5g
iZgY+KUOv7QCgbiBiIvg3qOBNANAgmdlj3iFLM6MvHcoBvLeWnpObSZ/MoVrLxNs
M2j7MuBHmiR3472OdWx1mo+eSD8Kmc3gazt4/RRDCobTBxwmOWo2kae5fW9NbgQy
FKgNeRLDuHrjvknLzNCTqbYtXOc1tsIQKLpXCLFllEQHdcp7Dl+TyEpFt2IVBTHz
CqhnQ+AYIrj7RPRZBz/1qqZrEZE4f8oPcs4w6rzXx4ZxxI/Fa5P5suKP6jMp6bgF
67Bz4a12o1TzBKCqnUz6q4nO04tg5ucnbi/X6r/lnezXfu1FFGew/LjqjudAvG1p
XYd78hQwcitdwNaA/yyBRWidBP9xlH9tf181QUrG8lZtrZclFG35zBa6ucxYuVLK
KywQlLypBmT4MahFaDsisWkcjhfVYzsrGjlMMGHf38RX5QIP0eGkzc4neFy/eDHL
vZIkdSX5zb/Gn7frroPE1pUivvUurW4lQpNsLeq6DBGbIGCV5CJxZtJ+LhpgYS2a
IGPgzIStNQN7Ih5AUL4j8toHqgjtdTdWXsLW8qWccnXU9LOwhry+A/cILpAMlvDh
fVlRgPx6oGJxvkJd5sTqMtH3/uSd8ms/13ZBgLPNqMT5HUASzqIYR/fv0SKpdHUC
7UShF/n8BywlWFODQqAdRGL4GqNjsHuCBaVlvj7KInEiapQAyCxu0tljZOGoqVM0
pIbXKldY+Ifc9V1CaIqICvx1/LYpj4d1nuGDph6czgDSIEgncw8qMTLRoAzdSBTQ
DLfs9YOuNJAh1qGFquc51LQ6r9ApxDT1yhgO9u6yBUXuMqW01kyExll7q+ATBjDQ
u8lzKAp1SalMWbk0/N8wvOJV8JQChwlnYezb6LwG+JdHh0lYsH6o0hjY7tp2btje
F7P03k5otRiIY5tRpGc+Uc2+dSqFwTG9TJ+tFruHNbQRLe4aMqYmbzG+NWFCpSJH
RdIJWjsVDZ6OPi6JePCe9fp4tLWoxMN97i193cGRKozeFH9UOyPov2sw3dR1D3kT
OFfDpBBMmb2TtIauVYgwlDQBC/CvrEkq+2wDmKOFFGUzHGtkgZf0Ov0kqK+iECG5
YVdmP4+8gjhcJXMYxn5LDmcVRv61JOwQxaxREUBYX9Jl1JX/SdnuoNxV8jqzlPOe
Zh0xazGJaZX8n8cxlpoqd53nDiRfX1YeQAB55NCv/zDWsQoQd3acHsGRy7pQ1RzV
qrQsqNxpsaKJ/yKCSmVTmujmRPrULsjKUHbgTuf1YOGHzgvpv/eSg5pAPeR74Cai
MRO+H/nQdaoaqLkErWNvWGVymtrnywGMRCHF0tlY6aWKIqd/GV4qDlpQgo6rqMlI
kG/GL8NyaExLTa16B872OiXJ8AIJrBIm2Cir7rwp6RKATZmjyQDAkoGswbye3rmp
MxiBMfkP//6Y3hnZO/IQrlzpIBIZEz6x9BawyyB8rPJ9aV6mAo/nvxkQ7E6vANC5
6TEQ6XoVVNg4XmfpBalFMSXDinN+ft+NcU6+ikjKPpfkFuOKmibqNJvjPuFND5pv
K06JXKfxy6ZZWVNzlxD4wp2JGSMr95ZPwViSiYHOQ/WRiTTz6huHZs0wnYkzb9OS
SqDnN8nljJ0kQqV/GYNSWts4W9sZ1Ud7cH8Xfn729UDN8/109B3sRe3exl62I+ur
P5r0dk5IXyAmGAEzzwQhCCCGam8pHxRok7h/884FZU1eeu7m0e+RZK5idCc3oCVj
UMhMyGYtgbygxTKMwOWVlEf0xjXMFpBRSUp7BqyNq8p79B88Qu4HDJBLEcU129J4
52A9zw3eGOil20cN7cyv0a6b1RMPd7y8+bxVyxh/9v+ZXix5cucJGVkscFHaSd2L
jscnXf904PUMkuhlfvqfYnfWeF4ddtf6Dtx8qHpq8WlMyBNb3W0tOgJPdr/CvkJR
DszZRlinKy98+pfd9O9ZJLqy6tUIiXpk0M3Pc1HgJAISsLNMQ63XChU4B0cXH8mG
OYq13FSoz7Zph0fdzozTcCg3W/slpY6zjFp/8dKPdv2MU60OzyJjKogQgXpXYm5j
ZBo9Ivpa1mjevTPTbT2cfBICEA6d5iWW6RtRTx200apH+w/aXwP4FT/PeWxBb6tO
51GkhQucrpn7+u0yVDyWEwBVMdug/rq+Zjv9rIQYLhDhqQ2c4QUmH7rtZtTNFIQ4
qYALPwm1YjJL20JHzDjTVZpO+Y+S5QryDNMi0bEdOqwD8pDtXmdtbE5HyZzV1I7v
t6pKju+5ssFzryZXhxTG0B0YBaPwZm9ZGCHAbha6O0nhF50d2o//405EcFku9Wgt
6jygNyG6Kz1t6VUdRWFV9UfavVbOLEXQGCYFFIEI82JW6UBL+45/Iq3XUAT+j3nB
aTgfSuXUdlo5YfSFJsEgX0KPDNmwdSoPUeETCEt1EBpR3j4RgNG5DsQVB6XMNTQg
GnE8voDXYXpaEu05xGklSHU9luuVIrFd7ER5qM0WMG2Ais8VFsuWrSLTOpgXLWkX
B4WUgBGBiPR+XR/LQw3uw8NsNxVWo9cLfz19ZjUbds2hulpRn7+vvqGyr+4m2ALJ
1q8cQbD5BNE+DGPU6UAfiu/TnmvmeKg8YBdTX7eF+nRuShfhEfEWwfJ6242jS46O
HrG2DrswaVoE3YbLv4pa8SWmILIJrG+jahC/0kRV8IOBVFJrq7f37u6UFzZskSah
kftUkqwempvR/rsqcCiRySJmxqEb8ZIfQT8gvae9r9rp6GqXgMTYp7tpUw2/7XWO
Ok5JtKdACPzhxrwIJdPsINOQ3jZFF/19wyA9bQpLSbeMpZfsvxz7A5Q+sQqAsTDT
mcfzlKTSjAOggxj+jyVc360c5hlQfW7FR/f63XlQH4ihdT/Mofzv+1nU4grOPvhJ
aM1Reb5CMAknqmPa+N4ITlchjGeTMT88+50D3WgzekpEoqbUvm5asVe0lxw7rzQW
tr7GLRMSG14GRzcRdK00ypzn+iMI0V1B5+s/7SCgWhlrqkWno0xk76fccLsZmp2L
MDfRb1ssJxG9R5cl560SJCTp1RZz7Em7avGmSQ/iMwMg2CcDtfG0LelYcUNp9r+l
FElqt35dcUPh/Lk524LIrxf5S/PvOaH3eC4N8jwHthgA+iqYJ1QemtEb66EdJDMm
H7yH87PWWS0OhOR/5WsLdVqNmNTnsC532dmJo10NyTKXck0nNwG+xuketnXySY8O
NsMqqwUIU2VUPIW/SzKhcDwThkv2rK+ljXWzEkgQsiQea3RB3TD0zBcGXgxsEGup
/BUKsqJd2U0+RzzW19F3QLjJL3bClo/dRJ7kfAsO9UwqUogQXFhpxAHwsshbGV/h
W0UtAmZ7mD8gMpJufmmUm9xedN2jAOjWjxPA2Ruf7BrCz9jIvpME86v2V3Xemjsa
Y5m/EHyAlrC6e+ytjnyfthRfnuo471W6TvjMBenFy0uYnlIbPUS+MFkLQFbh0PSM
eiIgjD5VFJixOY2FkZw0bzrgCoK6E+IVKmSY1pvC8NwaIQNFjhe6+mHTdfoEjwne
2Kfw4bQHhYFIJB7vnJIVRQtTcGISMm0aLWTMu2SHwPQkPHHY9V2S39qdRFTJbHK5
JVls0uLZrzcoTfjaWVdWAhzbpuvC9DuhxGXs2InE5oP3l75TYuMK0JLZsfDbqk76
NwCCtFf3u5sEc3kr4KZWTfhTbNti3Cp8DWJncuGbc00Zi1W45t+8ANDMJTMOqTGb
M8YPhUD1X3YjeO5RTntuAe9hvy+eGrtpw7y4EwxIVoxGL7/GYBp1vnpHeKRaB47D
eE7ul5EqMKKVp+wANXj7T3u6MnVKdBcrDzYbL0GcfhrOAqY//Zs9kcuNuY+PnwOl
0v9MR6hL3HxuZbRZAIaNlTmvf3ffZrwrGOlFPasIp0/ZX7l6U9vzeAtetwbDF8FX
Pze8Mhael5mzehzKB+LyleJYxq/wA6RJv4vWJOlubIcaF41GY2k9cr6vG+/mdbqG
OKzzUqKk4oMaTU2TG775SdR6R4XGZtJVfP9Tc+PR9utLRgobAVf+NjLcZP6ILEP2
qHpISEP53A8iT7m9dv9BJbjzGLEUAM/hTFfGDbc+KTPEHf/BMuIeOnOXfHkqy8IE
K3Yie5UK/F4qwDtaxsuMZelAmODciomdgh4BsjjA9QMVujTo12iaA0eHXmBLu3SD
uSzZBVVI3lNYn2rqyHsZ2Se1FdSHxwgJdSz3XDDIxgMmFVRaCSPg71F3c1YjeWlm
jshpR1XT7kzFEByGL6Amq9GezphxOh9fjghOcFfGSg5cppocHlz8kYdhxxi5mHc2
CKhNo2EFOOr3njJaV/xVQjq6DNd3rK0UEm4IAyzcvcloUwGpUnpio9o2uhaPCMdW
V/a96j3swb0DAS2eZyq6yXgDhfx0JDMuArpv7rHy3diTBleKWupBoHI0inIxdxiL
g6rJ6H4MkEafDlzQOGPKRY+6QtldzdQKGCSODlqQDjLLTCbbl6G45PrqdnsRfXzQ
2AcbRx7qEHDTtyBmpd4msSL96zONO5cm19H4IGHSF3JcIvJqMbLcLIc7oDGubNZG
QYCI2Ja5nwoff3qoVA2sq5+0fsKCBnFt4NhsUr4NMGB8VUWa5Bsgjoa4uPoivbpG
UXkm08i10BwhZ2iB1Ro4OQo1efJF18dy/Nt8erTaUBJm0pU3YRyVH2RqSZWZa0PP
ptVCWKbb3WJVxzHPrhBCWBry/FdL23LFAr7NMucsSReY/KTDfOvQW21CnWRL6CW7
aXSbPp5WjLuOLr+WMEs7spBoN0oad1Zax8L44yFg83GCSEpF/mhSSP2oAUazs6i5
uEVNVzlqNq0CaH58MV+Ir2Dz9/cos5SlM8QI4N+3FTSPRaVM+DwBjzpv7ujSM9KS
QkQisIuRIlOGLsiIGzKm7mY7HXudkBrq76cMsz16yHbIGZkwVIUCCc5IrOjWNWWJ
/83gVjbL197FTY+yxDAlC1Ts4bx8R6UwQdpsvGv6Gy2jMMNZkK0iKshvSTpWxJeq
eCZFQQDlrxvSp0uKPQr5LUlqVwwAg2sEOgoutppVYm58tAaPigodsdsKJpxdqvFC
nAoIfWQE7h3tBYWlIC15vIFBRdf0niakscHtHcpakoOOWPc+pxjEm5T3LXZF6Xhx
5e1Az6+dF1OO0eXcoCbdsAwnFYgPTa7NoWQBNdOpfJiGB41TmTokZYMk1kIh+jIa
pE2Y9z7u3Qc5A4jwm5Azs39/24X/XQ890BrM8rLx7Qo/NoXBTO7ZLksFbfluYcJR
zvkx6fwUng0CkHl6Lyh9U3X/512jM/OiuMnQwSw/LE4R85KZL5GJ9bRvBJ4hpBnP
7H/yusxsl4DP9dYCy+YNc68tQMZI2YyF/qiiMYZS3sPQioSd2kVu0UurLxkaSEAS
y+6hRkGTTlXBjia2bzBgGTiQFc1kkGYQhi4ZjsnnaiPLXaK7TNS6qttfKh3zGATL
CZIiGYZ+7R5FdSXfQiwQOc0RW/P8MMLz6BnFnm8Kj0l7x61yzCHmBO4rCRFnvalG
hyDtmyRYSoeKHo3L0ZtXvwWmjLWbNUu4t1JtqMfNKe0t0ZhqH8i66pfNEi4s01jn
SejxV+ZayT24C5/is2KKY+Fs/Q5tRznFg5SawAr0YZ2vAQQjYSf7Wwxr+E2TL3da
YGHwk23APQSm8O2upLZ9+z/O2ZcJi7vN+ggFdXTlGnB+LDqRjrRu4ELp/qGvgkch
LZUUJ8lG80RryFGd8LvruHFBzhns47ncRxgHDEAy4aZlWWoJK9kQULwJ5RM+5mRA
uw0vaKtxjSPogmT8ie8oWj3pDNy3VnjV8b1M0y63a4HK1Jvx9zZ/fo0Wlq5aGbMi
dO3tEm+Ukc4ntly9nlQqeQ4UV6IZHnjkaOIN3IBWUEf9pGB30L+IXkm9wIiBfQKS
7zgqUVglCYaQq86nGdJMWcfNbCUKBF5vBR8ZWhY13EjW6X2+vZEJLT7Y4cYmUprl
XOoPbFINp1iH6tT3zL6ReGvEOTZDMwhSW20Zz/q7lUnSMP2DgqACqbo/OuTVHLV+
mpYtByJqLwhywEYb+Nyi5xEphaPmmaG501KgIME/CZJ721vgT//XJUQJOrMMJTsO
pNQTO1euEOfcmOV0xpIY/z7xGeqmxK/bWYZBB4rH+PXTXiUdFAMpYCltnAYBj4sB
w6iP0zr8dIkLlqUy2c6IMTyAp8LbBdel5mKarunG5PraJJoe8M5XxDBp91ghrv7/
yzCNUBD95pSctgs3tKSnFUcCPSgIwI6cVAnq5OsBoSt/P6Wt+3aCS+SLpVYjKvUn
oxUYqjGPS1jVFgONsH1Vo2nx5XmBExdOr2VjK49wqLOCYSB6umoKw3uwRHb+nDMT
25rLR7E12BDfV/FqAuZ466nWdRuymaxIeWOqACOhUkm6KCLpMgXkVzTcHcS9x+0U
DsPuRiYB2zH5STOgMzyxTaJLMfqSIdBb2zwHlXTdlDH6fmi0kIt91qHAJPxVSd3j
rB78VsxStxg7lj4JEPifUJDt/Iwrv2ycc7AAyx1Y9hY+EEDsuKBic0azMeo44FC8
ncYZ9mKsS6OYxkdMJMPkUzIf5QHY/Qx1ixhkLjnq2n4Iv8WAszrDItYET2jj1AVB
wXDZ5dohI3A8+c7mC/dCNpqqYw+EFiQ2CSb+Bexqg0+TmqAl+yqV2C0t41tHoIR9
XNFbU1sfwjFTXOG+FvFymbkcQpubVE8IyqLIz0whE8R08ejaHcstj8buV6L8SYLZ
eX04icrrowrPd7dROponVb75jDoN9zejrvX7gMcebGhQ8eBFYgpJNDiVenGP4DJW
4Y4IHg+65X26KrUH0q8r/c9hVbp9iY3Hz+06uVvsbbwV8n6Fg46QNLuzfVJSsm/9
wHw+SgPRSnFocraSHMZzBTNm10R0lWXZXbB4dDvWB2gP19FPsSO63lCCesgk5LFp
WDRlJ4gUehSjX4lJaquMk6c53XiWP+4hgtDz34nG6Who29vdGFbFPegSa34hfRp9
nxetJNgUkunKC+1OMs+xX95f4cKe+3G9avUxTwQe2cX7zHOe7rWQEmZtW70pVmiY
wx0Jxthc+q13Pqph23uNrQC2TBTUtDor9WR5GjUY5WyiyxBJxvqzESO+FFoNbzdW
Fb9Mxy+Schi651Nk3dVm8x7qcMq4em1kTUL2utV8g1lVBhi+HD6xnsLw43w+esXE
NhWDCrVl3zrW0yaiLln9ib200PMrgu0wHtIrKKJmYmIA7hp1h3nCxBxnfW4hTbNP
T4LZJHldzPvmPi83OvXSoXhV+G65RsZ4BrkDrOxd/vVbJ1qr6afWhyvGqODPyh19
CKurS7Vm0ZbYb4LoLedX7ne1mJtvsqZNgqEHbjqjQNyQ0Muuntnf0Z/8R0Hjmw9O
l4lwbe2o+70CrHmM8Ssezr3q3zaryae1a8ncOqO2WCtYVDvEOKHw50QTW9r1SCVA
+BBX+tRcwPluH8AT8A6Yj5EMMlgXS3ag6B71PXApwIdqFdJXfI+dZQS/MJ72/4dA
EmfmOmOzVwPunN8hBK7J54c/x11W2Rcj7+5oygoGBYFqf4nky4gVBTBegls6tzyf
Wmo5xm8f78enqasjwfdAvgqsVCs9umjKLXmeoMcsEOs1yjjzIg2rnGrKr4nH/Y0l
O3zIPZvWOiyK/4a77BrsRv7zInkK72cDtqrRhs5IpfSOtQ1EPo6vWD66GnbB9zxk
u1/LbL4NObAeQ+2wB5wGnQI98BKGLdRibs2m/7AbNV+5QMDKO9gRezQlbjDxQDYa
oyiCU9lEbuzDAGUkwcKPrWxagrWIW0P7tIcaWAdDNjzRVudXO+R7rPmkEM6K2GAG
pvSStusMY2fjElQ+tGDAcjVOHReYPHptFznNr9dkax/AxW6XSDGm+p7mLji+rp+4
Q6cNKqCc1AE8MQ/E/n/6zJoDyvP5BDEEWqRi/Ndz3nxHiVxLanEGzqSpofs7IiT1
ouftuxOayVXMpP++QknIL2iiUCX59gZmS8bOmoZKYoflnxhQl/TuHJNLeWKI3ciL
QQaUl6Z1VETPDGZ8KncxfPxlzUiUCRZb2hnuD3lHMVN3uKTQSiY0wEJyBQzCmy60
Q+ty+5HpgSU88IIMggI22HQmrPIQzaqTsEdwH/nmAbY0yT93onBWK5nRQGKVcAkp
nv1scLQcjTqn2A3h4p1Z5kFZHVDOK8+0PtE9oSe6YvxkxDvz4TRyTN3YjpUlkaHG
U9ql7Kf+5W2jo1GuXxs/jzHS4vUFaGlHx4ABWf9sgJhgyHsnPQ0AfdlC0YQrhrxs
Z6x3CUZAm5Bh5JnXjLSpCrUJybMJCm2Lep70Bi/3NVaUXHGDnhTVjQhFAP3uKI5i
5egK5yhJQUfoDGHSdHtkywF0ymiS9ekzisdaHvk+1scw+a/spdwH5gppsFhetzld
ktUoPYZRFA+JLC/Ad5aKboIpbuLxBpK+Zn4YVsXT+2tdgE9yAVtfkTbqFFlqallR
FQW9XvlnnF0ZcaZwpR6HEUgy4TDm/iAAYkDVFOgjMaAkG7LI4qIQpMp8WP1IokWc
wbmZ/3CiCiY1w/zXw6YcWfstLtFek8S43/araRkJ+6SQDgIzBwbZur5yv/PkiKeS
`pragma protect end_protected      

/** @cond PRIVATE */
class svt_axi_system_common;

  /** Report/log object */
`ifdef SVT_UVM_TECHNOLOGY
  protected uvm_report_object reporter; 
`elsif SVT_OVM_TECHNOLOGY
  protected ovm_report_object reporter; 
`else
  protected vmm_log log;
`endif

  protected svt_axi_system_configuration axi_sys_common_cfg;

  protected `SVT_AXI_MASTER_TRANSACTION_TYPE active_master_xact_queue[$];

  /** Internal queue where coherent transactions to slaves are stored */
  protected svt_axi_transaction active_slave_xact_queue[$];

  /** Internal queue of slave transactions that got an error response */
  protected svt_axi_transaction slave_xact_err_queue[$];

  protected semaphore sys_xact_assoc_queue_sema;

  protected semaphore slave_xact_queue_sema;

  /** Semaphore to control access to active_xact_queue */
  protected semaphore active_xact_queue_sema;


  /** A list of system transactions used for mapping master transactions to slave transactions */
  svt_axi_system_transaction sys_xact_assoc_queue[$];

   /** Internal queue where snoop transactions are stored */
  svt_axi_snoop_transaction active_snoop_xact_queue[$];

  /** Internal queue of snoop transactions to be deleted */
  svt_axi_snoop_transaction delete_snoop_xact_queue[$];

  /** Queue of transactions that were a result of back-invalidation */
  svt_axi_snoop_transaction back_invalidation_snoop_xacts[$];

  /** Reads which have an overlapping write during its life time */
  svt_axi_transaction reads_with_overlapping_writes_at_slave[$];

  protected int log_base_2_cache_line_sizes[];

  protected int log_base_2_slave_data_widths[];

  protected int log_base_2_snoop_aligned_sizes[];

  protected bit is_amba_system_monitor;

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param axi_sys_common_cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter UVM report object used for messaging
   */
  extern function new (svt_axi_system_configuration axi_sys_common_cfg, uvm_report_object reporter);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param axi_sys_common_cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter OVM report object used for messaging
   */
  extern function new (svt_axi_system_configuration axi_sys_common_cfg, ovm_report_object reporter);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param axi_sys_common_cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param axi_group transactor instance
   */
  extern function new (svt_axi_system_configuration axi_sys_common_cfg, svt_group axi_group, svt_xactor axi_system_monitor = null);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE
    /**
    * Checks if the address of the given transaction overlaps with any previous 
    * transaction. If there is an overlap the transaction is suspended. It is resumed
    * only after all the previous transactions to overlapping address is complete
    */
  extern task check_addr_overlap(`SVT_AXI_MASTER_TRANSACTION_TYPE master_xact, string master_requester_name="");
`endif

  /**
    * Waits for all transctions in overlapping_xacts to complete. Once complete,
    * the suspended transaction is resumed
    */
  extern task track_suspended_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE suspended_xact,
                                   `SVT_AXI_MASTER_TRANSACTION_TYPE overlapping_xacts[$]);

  /** Indicates if there are any full AXI_ACE master ports */
  extern virtual function bit has_ace_ports();

  /** Gets list of system transactions where master xact is not fully mapped to a slave transaction */
  extern function void get_unmapped_system_transactions(output svt_axi_system_transaction unmapped_xacts[$]);

  /** Gets the list of aborted system transactions where master xact is not mapped to a slave transaction */
  extern function void get_unmapped_aborted_system_transactions(output svt_axi_system_transaction unmapped_xacts[$]);

  /** Checks read transaction timing relative to the last posted write transaction */
  extern virtual task check_read_timing_wrt_last_posted_write(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  extern virtual task do_master_slave_xact_association(svt_axi_transaction slave_xact); 

  /** Deletes transactions from sys_xact_assoc_queue */
  extern virtual task delete_from_sys_xact_assoc_queue(svt_axi_system_transaction sys_xact_map_queue[$]);

  /** Checks protocol restrictions for non modifiable transactions */
  extern virtual task check_non_modifiable_transaction_properties(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Checks data consistency between master transaction and slave transaction */
  extern virtual function bit check_master_slave_xact_data_consistency(svt_axi_system_transaction sys_xact, svt_axi_transaction xact, svt_axi_transaction slave_xact, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id, bit check_one_to_one_mapping, output bit is_resp_mismatch, output bit is_dirty_data_match,
                                             ref string master_data_str, ref string slave_data_str, 
                                             ref string master_wstrb_str, ref string slave_wstrb_str);

  /** Checks data consistency between dirty data of snoop and slave transaction */
  extern virtual function bit check_master_slave_xact_dirty_data_consistency(
                                  svt_axi_transaction xact,
                                  svt_axi_transaction slave_xact,
                                  svt_axi_snoop_transaction snoop_xacts[$], 
                                  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] snoop_slave_addr[$],
                                  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_effective_min_addr,
                                  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_effective_max_addr,
                                  bit[7:0] slave_xact_data[],
                                  bit slave_xact_wstrb[]
         );
 
  /** Checks if the given slave transaction could be a duplicate speculative read transaction
    * This behaviour is seen in CCI-400 where two transactions are sent for speculative reads
    * one before the snoop starts and one after the snoop ends (if the snoop does not return data)
    */
  extern function bit is_duplicate_speculative_read(svt_axi_transaction slave_xact);

  /**
    * Checks if a duplicate read is expected 
    */
  extern function bit is_duplicate_read_due_to_overlapping_write_expected(svt_axi_transaction curr_slave_xact);

  /** Gets reads with overlapping writes at slave */
  extern function bit get_reads_with_overlapping_writes_at_slave(svt_axi_transaction slave_xact, output svt_axi_transaction xact_reads_with_overlapping_writes_at_slave[$]);
  
  /** In case of WRITE transaction, gets the number of bytes written into slave memory based on WSTRB */
  extern function int get_effective_write_bytes_using_wstrb (svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact, bit slave_xact_wstrb[]);

  /** Updates the number of expected dirty data bytes for the transaction */
  extern task update_expected_num_dirty_data_bytes(svt_axi_system_transaction sys_xact);

  /** Gets the associated snoop transactions' data as a byte stream */
  extern virtual function void get_associated_snoop_data_as_byte_stream(svt_axi_transaction xact, svt_axi_system_transaction sys_xact, bit use_dirty_data_only, 
                                             output bit[7:0] snoop_data_as_byte_stream[], output bit is_snoop_has_data[]);

  /** Waits for all the conditions before a master-slave xact data integrity check can be done */
  extern virtual task wait_for_pre_master_slave_xact_data_integrity_conditions(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact, output skip_data_integrity);

  /** Waits for slave transactions with overlapping address and which have started earlier to be correlated first */
  extern virtual task wait_for_other_slave_xact_correlation(svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact);

 /** Waits for slave transactions with overlapping address and which have started just after this transaction to be correlated first */
  extern virtual task wait_for_later_slave_xact_correlation(svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact);

  /** Waits for transaction to be accepted */
  extern virtual task wait_for_transaction_accept(`SVT_TRANSACTION_TYPE xact);

  /** Waits for the address related control information of 
    * transactions in the system transaction queue
    * which were started before xact to be received
    */
  extern virtual task wait_for_master_xacts_addr(svt_axi_transaction xact);

  /** Executes the master_slave_xact_data_integrity_check */
  extern virtual task execute_master_slave_xact_data_integrity_check(svt_axi_transaction xact, bit is_pass = 1,string desc);

  /** Executes the interconnect_generated_write_xact_to_update_main_memory_check*/
  extern virtual function void execute_interconnect_generated_write_xact_to_update_main_memory_check(svt_axi_transaction xact, bit is_pass = 1,string desc);

  /** Checks if CMOs were forwarded to the correct slaves */ 
  extern virtual function void check_cmo_forwarding_to_slaves(svt_axi_system_transaction sys_xact);

  /** Executes the interconnect_generated_dirty_data_write_detected callback */
  extern virtual task interconnect_generated_dirty_data_write_detected_cb_exec(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Executes the master_xact_fully_associated_to_slave_xacts callback */
  extern virtual task master_xact_fully_associated_to_slave_xacts_cb_exec(svt_axi_system_transaction sys_xact);

  /** Gets a string with short xact display based on provided transaction 
    * An extended class can append context information (ie, the source
    *  of a particular transaction
    */
  extern virtual function string get_xact_context_str(svt_axi_transaction xact);

  /**
   * Returns the requester name for the supplied master transaction
   * 
   * Note: This method must be implemented by extended classes
   * 
   * @param xact Transaction for which to return the requester ID
   * @return The component name that generated the request
   */
  extern virtual function string get_master_xact_requester_name(svt_axi_transaction xact);

  /** Indicates if a given transaction generates a snoop or not */
  extern virtual function bit has_snoop(svt_axi_transaction xact, svt_axi_system_transaction sys_xact=null);
 
  extern function void print_debug_info(svt_axi_transaction slave_xact, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_xact_id);

  /** Gets split transactions, which are split at cacheline boundary */
  extern function void get_split_xacts(svt_axi_transaction xact, output svt_axi_transaction split_xacts[$]);

  /** Populate resp and data in split transactions after transaction completion */
  extern function bit populate_resp_in_split_xacts(svt_axi_transaction xact, svt_axi_transaction split_xacts[$]);

  /**
   * If complex address mapping is enabled, this method translates the supplied master
   * address in the transaction to a global address, and then uses that global address to
   * determine the slave address and active slave port ids.
   * 
   * If complex address mapping is not enabled then the address is converted to a slave
   * address and then the port ids are obtained using the legacy methods.
   * 
   * @param master_addr Master address to be converted (can be tagged or non-tagged)
   * @param system_id AXI System ID
   * @param is_ic_port Determines if the address originated from a port on the interconnect
   * @param xact_type Transaction type (read or write)
   * @param is_tagged_addr Determines if address tags are present within the address
   * @param is_register_addr_space Returns 1 if this address targets the register address
   *   space of a component
   * @param slave_addr Local slave address
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @return Returns 1 if a matching slave address was found, otherwise returns 0
   */
  extern virtual function bit get_slave_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] master_addr,
                                             int system_id,
                                             bit is_ic_port,
                                             bit master_port_id,
                                             svt_axi_transaction::xact_type_enum xact_type,
                                             bit is_tagged_addr,
                                             output bit is_register_addr_space,
                                             output bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr,
                                             output int slave_port_ids[$],
                                             input svt_axi_transaction xact);

  /** Gets number of snoop transactions that returned passdirty */
  extern function int get_num_snoop_with_data_xacts(svt_axi_system_transaction sys_xact, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr, bit is_pass_dirty, output svt_axi_snoop_transaction snoop_xacts[$], output bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] snoop_slave_addr[$]);

  /** Gets the number of slave transactions associated with a dirty data write by interconnect */
  extern virtual function int get_num_slave_dirty_data_xacts(svt_axi_system_transaction sys_xact, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr);

  /** Sets a variable indicating if id based correlation matched */
  extern function void set_id_based_correlation_match(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id, bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_xact_id);

  /** Sets parameters used for sorting transactions */
  extern function void set_sorting_params(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Sets parameters used for sorting transactions where both master and slave xacts have slverr response*/
  extern function void set_sorting_params_slverr(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  extern virtual function string get_ms_assoc_dbg_str(string dbg_str[string][$]);
  extern virtual function void set_ms_assoc_dbg_str(string key_str, string desc_str);

  /** Utility methods needed for correlations  */ 
  /**
   * Gets the minimum byte address which is addressed by transaction
   * 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Minimum byte address addressed by this transaction
   */
   extern virtual function bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] get_amba_min_byte_address(`SVT_TRANSACTION_TYPE xact,bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = ""); 

  /** Gets the max_byte_address for the given transaction */
   extern virtual function bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] get_amba_max_byte_address(`SVT_TRANSACTION_TYPE xact,bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");  


  /** 
   * Checks if the given address range overlaps with the address range of this transaction
   * 
   * @param min_addr The minimum address of the address range be checked 
   * @param max_addr The maximum address of the address range be checked 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Returns 1 if there is an address overlap, else returns 0.
   */
 extern virtual function bit is_amba_address_overlap(`SVT_TRANSACTION_TYPE xact,bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] min_addr, bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] max_addr, bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

endclass
/** @endcond */
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
XvwrqlquVkdiJ2qqG23QS1rbYxE5oo2pR7MTrajb2G4Y5VLmhzbG/rcU2dzEoFkp
qZCFwbY2a2+9HrfgQWrM+IWNeK0NdrKOb7JUiMxuusYriLovvDhPYi44mQSsDax1
KR3ZlsLPIJMaBV4DRWw5lIT17OC1LawBcJRf2FYNLCQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 11813     )
WwsrhHWVGmGFXxvnIDDiddOrsmiRAc87OPjzU7S0siBdtcI0OTK+Am3g3Gv8OSkx
cibTJsp95tY54qNTbdLDKfzFfJ7afR4N51+ok8SfRBF6RgYSuvedEbXMXei+ETFB
tR5XYtYYvuPWxG+n8iCX3oDNrWxvKqdBe2JuQoM04vNxoHTbEg5f2CnD9bFLE8H2
g3Fhhj3PFmhwIt/boJn/8sAaKv/3IZlob4zDJaN1s2dqrKZfendqg9c/g9joVluV
iYwiadYPonTZ0g8nKoeaT9UBxRv1D1W2LcU7jrABaSxisD5iZC7QJVfZSRI5kz+b
BLr3UxBiiyqqzwIqIWu7QymZKo0UzAF6ERn+d1dqyrkZ5TN8Bz2Hxg/u4WI8MGrf
nqDIc4Y2IT097H9fbP0xuXIbIHMCN7PF7coBExeNZurQJGiqvj+5fcjowCX5jQ97
tJRzEDjmvXBj3BINWRUe7G67C5yguBBrrh7/ht2fWqMWhNzSJMeXDwNYu3zhntC3
6FBepDCvdy8rxHolrWtW9mGsQ9We7rFVCtIy4lZsE197+Ya/3Gy7+ePDppWnpNdR
U90DZQUoBfpWSf8w8MEATa0Kg7UbraejLT2wJxTGYg4KLa1FHGRePUp73CjCCfME
TBnwzfdAnLLGkN6qo9a0qsU8Fulq2Vk27v8X7wndVIaFUgJ7d/EjVfjdWqtB1FM1
dccTz4yjGiE1uBWED58X3JQLKwJcEK9iBatT8C5YNv7eT1m0saUl6ZQYwS6VnE9z
4ZOEHZwP22+yvvqJA9kZfO4JFhV+nMEssIWkQQr1QpPN3a43BmDMu50B/T6Bv6DB
gA2b2bRSdDEmkz9Hp/rZ8kMRbOpcOEQ6VCs9ALXDhRBf9OQw9y7cWs1/LIaZlk3s
ysh8/C6qAiW/C3Dz+ZhSIeS4fpiGt+MEgX49KaUO+ppkpX26IT1hYZbvN+l9NraW
5k2QE5BOOvzAShbSzjX7PhQ9XkJjgdko4mopN0Tlh7LntP6kFzU36tau9DXC+KVL
urHGRUpDDQ8Spg/ZYJBvscHEAsgdIeQPbe4em/YmIqbNRPVRna6CwuNG6gAdFkWb
Z4AVYoGB8VRhIotwbkG2iftHm3B0qTSc50e/PKjf0A2fCQ6KobdBMwKvlxIfrY6B
brEGGJUdssYDSWV3a/ONgd8SIIHUjIimqY9VfDK/Xc1Eu8wnOqRJ4y+LpfBBWeHc
95CyBD6RNYTDbNqRBEdnXIv2nqzj6Y/3zjVn+INtg1F48mv3iEL+P/Jyos3r8jvL
aZe+vwNuIqSf02uie4Vap6MYq64xvdHo7bozlgBl1EwlvhA8ivlS6K06ahBOvVvV
nW3olc8dbtPSEg4ghUjA9tqB+S7NoNZJjZUjtEh5vaar+MItOQgwErHnNqQ/vgwm
XMlij1M4rv5Sz4qDlB1tBToF0TTTs+ThspqC7ZFcPTijUK0MqCc16thH4Ro1dlrK
g8YKSMomFu859DWWN3TsXJA0fqn08Odx9GZOwcQnroo=
`pragma protect end_protected

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OfJrdiR2HLSaiktYWewqXrrPbADwKnabb/nIxtFcCoc6+1PZ9qsZmDyQeYbkooB0
0OXTWMFtxEOVFxBuO5FVLrzjh7iTiszDs1qNAjKm/jQ6robnnlCeSzGMQV9HjYBB
UFFOfASde1X34vZHlEX2K5dj0cga8FHh8sdAIDcb4Mo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 31247     )
fmKvgT/KyyLk6fuu/3VSusMnuiOL/OPPCobZQHnexqxLYRsXVExZ9HZPVvPUSc/7
lOZa7xutJrvo87w457w+hfFp6TGpZTztg2MtR9034ljyjQgxqTNR/JmCSi+Yh8GU
fe+G7OvVVUWg0UwtdgMWdtbsGvuiyUkf51mUOUeehkr0JurNHGZKuGqvwY2+hQPr
VWctM33QKW4q/BrSpwrnrsceeHgw3kDLbPnYJ3FtbgFoz+vueBDa0pb6yy7hNEWn
7EnTAFadKMLyuAnxcOqhnqBZIs2FuSsg5EijxYrEqqVO+/XAOAsuYA/6PkxRQPpN
XhiLqm+ekjhrT5J91XC4BNxZNR3XEMZXeoUA2EJHyMvqVloYlwuIbf61Wii72enR
5RvCCcXCUE2CY1XknoT0PFQ8V1lp8dGyPQWSR02IgSd+xtJMtd8AbuvIvH3TbvNS
KteYRJrT2VRrWH1SFactIvnO4rhLLaeBIoi2jedHuGipgNpU4GvtvmYw9lWYS5W1
Q7m8jOE90T49h18QnT8YQ5JvRTuaWhIgfRFyrU8qhTTKucdvxRXsuf0gjSPKWIII
5AtkySzQ1Ya07pS/tcu/FItnLTmo+EuESs3FPqteWGsNiQPlcmxskYbEbBLRT7XW
tbJZEWMsq8LlO8Du/Nx3sMYdank0ZoFEzcRmLzfkS6RkJL9yH1+mVGAD23Lub8mz
1w2LHRuxAsRVqN5gOqvRFEyhBpBoIzab/caZ4cYiXzPC1BkjhCCCjH+GNgCsNOcT
WtQeiXe55aNN6UVEB6OWl4Tmt9MxBHMtaOYr+npyK9PfT0/xGOeYXeUsQ9hubfqf
Rq5lWzgxKir4Nsb0bpDlnbJDyTA6fniMg2coxwGYvj0kfZu9ulAJiKwB8Uf8D0AL
XLAi59lrAOq1OEsTeppJ3Nad5AmuMdkO1+8CVIVFW+vtQvuuy4wIL/LksPaL+o0s
fagut1Qg8L/AIGPKzsoKYbpZZ1goLlU3RgswJ7BUnkD1ZPpMoGmTPGqFtupCxscX
SaSuWYN9AGSFe1+GecIqo09YBrxyFlK18XmR8m+TOSDi7XfgPbl0No9SiCFIExvy
7FvCMEePcGDAJvnmqpVIUGvgn25kDL7o1psJaeBK9WJfd1ujOsg80nj+UWJpX8c1
dWMBsWzofRwV7niLqVuXW7klZLHsojGEm3IjHJppfK9CIBmoqxU2+d+aWC7pwbPX
k+oniqbt7G9wk/MbxIf16s5nqHI0YeAHRJfQThw8Y5In/eFmnVod8ijNA2MufPwa
NSIkc9bVGt0FtZSpokC7LnHgGRN0y/nHaQCLd7GptketCXoIVY1qzV5I9jBYXyOP
PC8QtukaSj1mX9lGjo8HRLPszwgCSym5q/Bu/mAwusKiB2PRxKkLJ2zAoaip8pUu
USw+ql1+93Q+0OhgUhSOrShTTkdpNvK9yyAobFzmhprYxFCyWWFLH+kN0xJfxg1U
Me2GmlenQq/qVONdcKqXEEvQSHlonwSsi39HVIc7Rb4P962VAlPTB7EqXxxNuSwh
p7oucbVqhpL/KiYYe0zKJTqGihcesuiOKV1S8tjDX3HXNk+hZTjVfSHNlQIFrUHd
wPZHs2JJUv/Snpi8XoV709CtNjGDMVLTymSFtfxu7ymRjUzSbKnbQlO4nLM/kZ9X
Hn1ZwYZ/XrcncxBPhBeVGqiGAQqz4Guzo/uEwdnzUaSF1GATNX7z6GcXotg2R+RD
DTMUvlAs6IVDZEJOidIwp7yuXmlwki/QN8JhD4W9XueQZuzO3+8uA2SahaVmhH2U
yIl7aYYk/OMikJT7WFaU83d7E/z3o42wfgTU5tAkvhbEy4EKx4/SdwftbnKCzd3t
BS8+JmmPHadlW5wxugiTrMQk7Ds5hjvaVqpQ12tWXbYsl0doyL3wLEea+cdJxKFD
iWTO3ZV8poJMIRtMo2qh6YbF8vS5nEhL56r9puec70IiKd5YNDZGAH2ztyB/FL+z
leEMYuLy8TKrcKZewMIQyFqtd+AA2JwV5mslfTa2wUExxI55ujYm3F2H69Qs5iTv
AyV7pdiMz08LsmBWG6hLCM3j4F3qso1GcWpois7EW7A4ijUgh0EMtEa5gzhwKeod
j2Xnw9xq9unwqRwoe8+QpzrnQa0F11Cbsck3P1zFxGitW7cgR2kbaI202lKQSKBV
NhygyrTqITT65HqgBeHOygnPOsLq5Jrw84Mst1P/kgXTesq/gHNpk8B5/MzvYAw+
vE6uEDth9w1zAfySC9RFaCjOt8Bz0hkykPrNcQPly8v8J8y9iNDGIc4lDGUwJQ2n
24xxdRsn82m3vo8dHZy+fCOh4FxQHcy7sVU3hDnY+eRCteHP3QY4m0GNprKU7SsS
Z8ygxC/qArFW97Kl2xfhFnvK2CS3nwXUXFAsLYJyRYiKNAg/xjtsaKNtIn2tZ5UC
qrEubgZ1GSvgwPIHPri53WfYUaGUOwK7CDqJYOgp6BAqp5yjfoblbipAMTdYmWoW
fKnwH3Qis6Ze17hfPWv5SMnz+ODA3lch/WgIeiW/x3d+ZJ9KRM5ajw0uxMhqgTW0
5Y/eCGIM3MPC/ReMK9fDCXoM88PxbMb5FZXMrYu+srVfz72z4ekUKhTaoWu79P8W
sDgAtNoQnO4wDKbaOCOl08QFROjfpXnF+cYYh7M1fdMvfursKAjgTScQsVUOqmRL
x6L83P2SZ+v+RwMB64zhf1lAKmocLARWma5tuGRpQWAQfGWWOyrcbBirNDFjPpR4
Q9Yv0YN9u44ifUdcc6v0BSY9cRVVjlAYz5YR4koWY9uECxp7Lo8Ro8kxan+MHWr5
NUP7fG1pQ31fVOtAhuq53zt20bfZ9HSUYSLAC9bVF7KL4mBnUbouno6aUzisDuBa
CIaCq9jU1EZeLmwUJEVbzDNH5H+efb1ldfqinQD3vK4y5bB+lWb/Ytp44Fjn9ibj
zWLTdlCDHMSdgWn7axI+8RQyeqO9cbfcKGVwnf1+sdCZUFWEFT75zwh7U5/Ja0PA
jOpymNxR9xF4XYCe1fkbSqu3j2iYJDQav5mjHpvGmp54BtwrKC25/94BmGKwhAx4
0GabJ/IQXAlRnDtb1Fj2/zEB9Z8HzxOARW4txgLgquEXucb2CjMm8IMm6h8a8e2Q
5oz71PpO29ZpAxSgWIIwpoG+ncGZ165ePXRGgdBOQXrMSxo/kKw68CXU+6qTf6YA
dDLeBzPBkU1jF8G81tpW1ts7oGk2xuxt51xeXVMRf9p0seQX4la3qfCw4GmjSVxb
KkpXTvNtyJYefIvqiZzk5N6EpSBIjgBIkE/+pQFB+SBzgccrAKI5GGw+RMdOM1FB
e8toTB3/dprR3SMxl/RmS4uI036eY+vh/Wm0uxIcyqJKVucOt/8pvXzdP/ge+c+k
6XB7QUmPFjMq0YcMHB5rkw2R28VMFnfJTlwyTTdhndXtVdn3MudQeIGLStlk/DAl
3FBvRaFUrcqWFO7Y1Dyjxisz01iUNJ/gVaWL/dJlLCcQNutWO9qW3w7Ze5ct/IaJ
2NqNDBSHQRsA9s1FmvvvsAGSgW3EAe+SJ1bJpvMt5G5svv35Os1l049qBusKZ+b9
f849AYQMjeslJDFRdXZ20qO5mYtmPulYf1RBB09XKGnZ68CsOlXgVIK0UK+rw015
6YpS1ERK9+fyxFXs6FjFb4xeZq2D+aXAqzvQFdenbvSL0pVMuM08Mekb+93piVa3
ctjvG6NUbO5VqU5XZ6RtvvoTgoSS0h4iDQmS3sFkOMICEJdBJd/QCdXwfA2Kpyo6
knPxWgDYiTzAiaymSqZ+W1a4ozT91WuVY1a32d1BSOqnmx2JJ7VtGVxMlnvFovX8
xKy/Cwxc7RaCq4gtcq24fa1koNtkY3N0tbMTmfz27f1MJ63HhdAJO+Bf6hiB3vqX
Qbqg6mjK+4Sn5h93d1nLnFJhq9lo9u4ZnjPs1ULDoCJv1snPi3bQU+6XNZnIYyRw
oOs1jyeIZIhwdHAwhCJV+wBRHkWFpcBebP1A2nfbwQ0T8/UB9iKhZ7EU2uLmCy3Q
5rV4NSZUbffO0n9sqswXVV2kRgiFDX3d6ANvmOe0bjCikFAuWnbUBaVY5975+TWZ
Q6ZIiWMnGhVaDI5nnfRbcHaPIeCcs64AjEBzU+rbRuiBDx2mwNTLWdegpx+9937A
07v2wdMeXsuRWZIeiyjSLCEHXLQE2DguCFA34GfciFu53M6GmdiMyvFsOyCLypmx
5w9JVIsdbtBck4znLZ+0BKsRA+Zc4g8YLK7UZNVGBAzHJfhg7tz+753pljgYvqZo
EGJeValwcw9NAJVs0LIV3OX4ApzF3KYTYDJaMjH5YtJHpSrdmelwFEHkQiKBbzMt
CQjC+Q/q6EaqvgUL8Vr59udMT+Jd0GZRyRr0YfXEzkXM/+NGEksztsg+dpZmogrN
/mb7N9/9+ilkk7stzqiacdqkV0YJKmq0I6+C3z7JxSoer+tdi65ednG/s/c4b0T8
wbpGuuHb3DKqVl7AODm7l4zJn/0llCewtPWb0lN7aFWu2TffQf0kpTsHj3LDluP+
wt//XX9oUfY4+6kVV57GaQCEAMMXCrA2sJDwSLjoQ4mhJ9EGsJbL1atoyf45wyBd
krCaE6YlleqxQRxx14u1/gsUCMcsUDsCKRm6yADJ/yU9Tv9n2npuzAH8TyZ9rgo2
j+s2rHx3hUwAKKfjhN1dcD0t6xmXkfDNoUYQ2FkDqD/a3W6kETYOYkjeKRL/pi98
nARjOufqY2scDfQ6oHJQACXAxzYAex3l7LBTBQJQXgnQKWwpKp93xkzx7UQfiCN6
pBzBdx++v9WHSWrqulg/to5xX5c3cfvVsHsqjqaaou4anjQPO1QwBTd9RRdASG2/
deEa2mIaEoqcKxAltfBaghabB8RYhK0x7qsGcdVO7G6SA/NetvfymMMe1TmxB8nB
8t3/tsHyij54jRrolFwQ5iYlHagu1CIPdBgHcMVrmvJ2Iqv5tRzSKDTAgTLVNGce
8pRjYV4AytM7SRQ2I5oqggsJpW5zvv74hAXVgGOzw+kzlmTHu+XpuPX+Cwwpgcl1
bel7bdCY+Y7ddj1l+BWhiLrUbp3RoVTjvfXdVram4oFb4VTBCF5/3C/ubkdgZLe4
xFODnzJPXfJES2XirlENaOQw+Pn9WNKe9xlrajLPvJQI1B5Grv9C5T7/HEtfNIhU
lxm7zR4wUGlrYq70wdLs2XBl0iJHVG/LzbYxRRTIvvJoSaIq2R3ondQv46zaSxpK
j9y4D57xWfdjo+fj+Jn86xZpb8IiWiBXdrRByh9sfVZMm34V9vFzQqvd8167Z6cb
YBY70ZWKOZ4FYluysLm+nZJkUxVfdZi5s9GLa7PIDxdwqtDqhQrTSUlw3exNL2CV
rW4Hzda0sAsBg96TSq9sUgM8egzoiBch6EmUT8S7sNUYo7o0+T0W5lFaSbh7T7uU
BPq2zDrgxbZXahGp2k5ROFMxl+jgQZSQKLy/ujqVETufHMLO9ZOSrc7EDqxIN4vD
q1jahxVTj3jJUwE3bEKODaTXjOqCQIzGly1fxXfIScONwxgrstLxBditYPGh9g+h
nyNQ9bN/pieAKMpkhY8K7Jtl9o48cT0LC2t0BX/A8GEu93uqAbargrf7TTgatv1l
OU26ATPkxBUirQTK5CiQFGJ0HDLh9xoDNw0mKkMyivMzD/J/NDdClLpelr5dOlpy
MqyqQ40hpA0xfqxgCTJJ/CkICESfdk3kuBfF0TdhVYB+ts0S3ppTBECXkQIN5VUx
X0+anVkBtxfJs9DzW1oYNk78zR2HrU9IMQmL7g3HKCD0RVMLrBZd6ArzK/8IeRAk
Zrw8cskEZgP8uvA55bntRwKSEydSJ95ZoQ3bGTN3l65s58EWGY2BulbkbPkkP8Et
7jWDPimyfRti6W+nIwoI81LDcwezOTKT9vENAnvoaV9IJ0TIM64z50k1sMzHkIMR
N5g35L7khPVz7ztcNx1Nv7Qito2IZ/QJwzioW/ENxVMB0khkYRzSks/1QUKvQYTE
//nWgZe+I0fwCUG07twDI5rfG4sJewibjPTpXyOir8eSBWh0h7Fl9KtWLB8ksMBA
3a51Zh0W9KYVH7xlCvIYhNKXLg2l3d7lGdIQFgP4+gNwxiFrDglxF2S2osvlMK8J
O36UTP0Ty7T126eUJetOjYimrUjHuO/FFZRr2EEYtHlISHyCZSPNlsBWr2ZHohaV
ZmSBSrYPbBEkzseCM8NXRT7GteKvkOsXkHVKzxPZvH9SDJbeEIgfndn/WmAM8Y0Q
vZgQAMhCwaTbTIPtVLhSsQOmrXCLNufIRjFROVOdWTsGIrbc2W3mAyQwH5nafxq2
SWcXgIuySkyXBlfZejcnTvmxKU9/D1rb/mkq4Vm4NT+k2VTeGPkV7h106p0aroO0
C/nAklYHT3aCkD782mQER8DPCUc6ECGl9aPRERHnp1/P/hTQIBuHkHBFU7j7gHdh
oJSSTytWh4osEAfMDvtY6OPyOMyrVYxtLVh4kGUs5wQ5SGxNZHEHQ6hCZKle+PlQ
x7eLI3SRxfIJlqbZYkvJrCqBulXiVHiV7/hL9GB0IaKSVBA3LCrtcy9B1Ts4h2Aj
fgbCU1qXKWLUtS+4zKplKrK8V5AqotNdBo0C4FDHhUzF/MWTtPx80RYghR9alv/g
McDc+s0He5Z0uf/JS5UkltNZ/xWL6M2BGr08SM7EL5w2uav30EkL2Gz2s1Kmbkzu
rc7Tpw/KdT+TwbCQpjgbEjE8mCKndlWoh36cSymuNW1gytMeTpflP9+16awEeo6C
k17rfM1kKQKttSWd5Z5EJOklZ3EYWHY9M/nLJpe+n+p577bFj/PjIbJnEbztoDXu
iCrJVai+YobifeWXuoASLEe3RMUDpAA5TUlmaZ1Mj3ixucZy2XFJMcZmcgHyz/eL
PIuyQjRgMivSLcq5Ay9nXAiTEsYPahBKQ7nVFakxWoOQMvHa9oHRXkMxKhnlBjtq
kKEQNVz1R8pNkCxykb15eZcWrNjtto2+pwUl/byHRNJof20n628n3RutwRpyxymm
+uuaV2K7NjDlYDZkRlvhHhMc+EDIQC8rqyC74kY1+84dF/js7rzKrR8QelJKsZmW
XCIonDRNtJXQ/0aPdRVOXCouLpGz3vCDlqkgW9K3U8WkKgIceJVBUK4kdO60HX/+
Q6cwYqZbQ3VLDxoKwmr8uunIzujx6WMQxJ+teZArqAO6AWJaWTRZtQobnfom6v5R
qobI89WURb4ivLqff4ePx95dF4zCXQpVfDw2i1HR9h0uT2bMbSX5KrQrcJ0h9HKU
gyKoisJ4BColgpkgjWRCCO/lSWbOy0t2EzMdsYi1UoqIeh9MpAw7A7PjTk9xyEli
f3V1MWfVfIxI1G75fJfmqV6FZWof3+ctkXdZQNmumD9e2q6vZr86T8to6xoSUPNU
t462PVuvn+/Z4rhXdzmRVkwU6NKhCc5UIy18VFj2yXPocyJgIgNn/xxsjJqTCn+w
j4Jn4HZCmK9o5NPy0xPIm1fOwAzKxs6UQhe0x8oA99WfsS0+e1gL3fH9QNtVZs3T
++m+37EVe24hhWtJ0m7QSTNsRwv73op/hEL+DotK+Flo18ykWmIKGMiJkUVabscE
KRL1G0QlB3Jev1cmZ9P6nzj35JoNXRcPu9LUYhyLodhZhwr5k8+yynbDBH+kOSqx
CSAgqsPgSHjJ97eNhX+oIn1BqapKOj70kNCyQbgfVW7yMir1wBUzB0goYYJ2hFJh
qc0S9k+bzvrbl8c0Vm/t9A5wAxlMnqF2i+2aYaXMHRxVXZRDrov6AgjDW2RwVtqN
VimuhY2xBvG75uz6o4pB2bxiMu8EzTdylZesqFeg0ezTAsXngWaU6ZxqW1GDDiRU
WOfTH38SHtJCMo6sHi4mTtgXnlZt2bmZGmKmcnZwhG0/DfqAVGBYq596aZz0SJ6N
PvmU2ARjrLxtAKxDRjbIMDygloouWtPw6JI7vDIVtVrgB5V5bIQQjVlOjecXoom/
ORCR3iN+40K3Uuyp0IFBW4yk8r32QRDSYVZYdDreWwJCPaepeN6E80zE6Q70BVAm
K++byexPzp6vW4iyx/8ZokdWWgiv9rMKPjBxbpTbhv88hL99PPDwMLbevJpCn7ca
KSN36CiaUz7YCbt7nPKvGhfA+RhRODLNuvCOgpERcWoI/QbWrfE/yBA7HOhIlVUK
ezPYLjMRcEZ5IDHuuooznZ85JCif4dTWr3ow2gPj11lrdnb+suMX7QKvo0U58c9n
USvv1AHla4zh0ik7qocBF4YS4Yl8BkZFwWICtaHPuFFZlMKHfxsd6HYR6/Wumusp
lKJnVHF8Wr5OdRF6ggGSCyzabTR7mO0CL8A5CgSTowz7Ung7r1jHCaGwg5Q5YfOU
yHw03kdtGKZz1Hp5PeKCnPD+WevsKiNkrVU9H9einvw9/Tvm64ZGDNN/8rJ2rkQc
7U9a3sU7mU3/opqjF0/9mIX9LNBcwx0ZXTWYfR1cub6dUyN+WyqZrqb5xp3uqP7m
51Hb1fW091sgf4wbmkF+nkIoeaU+zj+OI5OZ7h0YproBjIAiDvHN90gUsHxbmNAw
59xNfJ6NezAn902z1gh8gfn/uCIE0Yo1GnWDm2uU4tHEuXZiMhTOWrhZ+vfZMMS2
bA7HvG2iEv+aTquM5wQsdpjRMTOw41sDWiH/KE+62jEaai3dj2lwjrSbYghfVt6n
dTFAPZ/dXcv7nDNkNIwCEoWYZYKDiGk61sqKq06pNIQMMRL03mIY2Q9RYzN50ifg
8mL/fPICwMCckPSQ5lU7jMvkrtqvJUc7lw4khFdMzRvq36uzhPSGCYPdnMAMsw3P
e2mPK4F5DMEcPyNZ7hlqcb5aqNnt59vAfo+53cq0XMP9lPsgYy5aNcCZjMtkyEJi
pRHHSKYwW0OEuvBWjGJ3bYQzKdlkp+A0bwWerR9yIeX9qJo3gUr6GHRUe/hnA4bx
Ii5/TnX31v7r4MAuZ5rn2HyyPU6n9ZzQY0CQB8pjLj43ExQKrrRI4J4FYEotr+t4
P1NYw0H+UFEPJ4Oui5uUeTFEgEkhMRoXo3HChIMtOo0+lG7TQbwVgYsA6nXPrd95
0Nwch6Y32SFmbODTa8OkN6jK+Nm8omXpzI8a24UdFzuwTgkkcL/LL5SNOKYhgeTK
deWuWJIT5d+L7MHDl3Cc2UAbkwVjDMi539S+dS8ugPJ218TQU1bH26nziMyiye73
sbrYZ1iXyqY36bY8jJujJsuBKzKjXjvij014SQG2U7Z+bCh61NqbrvJGNH6aqthe
+Y+gP1m0NBqE/dvQ2LwoKK9XOF0f03F6ctMjMFIoYK0qAfAPdgGYe2tHtp3540Bq
lKe+Bq+dHHAbK+Ze2fIvyUyX+KQJTqlHzRnbwkgb8zvRbqvpRnBh32j1wBjT4T/x
ZYsKNtl0bjnUH956rfUvFmBFQQq3zJlWg4lRrEYlVL6MxQJxs6Gni4fP7Crvf8Id
WL/4Iu4O2w33w7ee1K4AdgK6q4IEDVgQ9JJjv62Q4cIypaQ0mWScqJ1VWRYmL3Rf
uyx3lDwxD0bjSugBeUZneiBUZg6/QdPY/99UlRFzRFdXSDkPpsrdy/667nK69BRm
TwWBevoYMF8RTKglWHbq8w+AfJ7nNj3VZ/K7UMUmXdmuWz8+3XHvN0VwJfW0Xzs0
N9c3tjbo3jysnnZ350xexYRgOtd1Kj9Td2YJ9lbOq/WZgVQ5JuZA8fpcLA1tIcf0
xFuT4BuIRy+7aPqoPweMwPxSot4G2/ouy3oN1cjomV7tUYP50nJ6Dd6LxmI8sZx+
axqaB3tteZCBde6/05C2gAleCGbxm9Gl2wTOios4QD7gPq6gSaLcKFOLFzNsh8sS
9MtMIQY13eU5WF/vJmBmCjPlvCtmRv2gXTr9ope4I+SNw0hDmaV4i/y4TKyUcHTL
YC86HAqKCNyfoz7gIikOHVsGked78uroXLbpXLDQLUa/IwPGchK3NciWrpIvxUjH
teyzmf3iYihuVLpjR6smGsjjYAr44806odqQmEBC0IVeYuPRNeyuQJC2tJz4xPYh
a8ZXOELut7k2tdzgggIVbPP1VNysNTSNgt6pQEaufDALzAtiNUBRPFhDyvUpE369
qWm2Piiln62gIc3+4Sd+69z38DFanrPyL5ab2mIR+oxiiNEiMVVKXJ7w+BR5hcdt
USd4QT1Hc7rNKZDjbSpU2lOamySiBvyjzJ+zKbewpbEC1dSRE4vLj+cbxf2YGXej
N0pCtWalNPUH2hmhOmBgjiL++MfjgddkdT31ROdjT/m6QqMu1eMv9F5tgwuGmTmO
9DAWbWmilIC2iELTa8pcCfMJlDY8uoixwhmxNO5v2x8RgfreVbvPH7Mmnp+ThF2p
wfkQiYlpaANEtwSp3wlFY7EECYE3WdYWV2sVI2Utbp7LpIhcDyZ3ap/nnJX6VuxV
14L8eaavam5dGNWAvWfxoqiiqsscr2sAZhfzO7XqueIG8NkIMcUD7JHdjb8WF+f6
48wXZb3kWgi14o8T2SSbwnD5mboCtyH3pjnWaBV4v90zzdTmby3sCTbMZsfaWGAc
48TiIZhIn6h9NeOJg7O98sAE7l8q2s87aOYEQNsXTaEhYLTKio5VPfh6PWZ+zDIh
zSkqKu6Lmt03S2OoZYRiwLgcjz9McJFZjhqIj6JxSvYb4X886lT6qJX8MiQofZYF
jCjYQmHvhz9x0Sbm2rZPSJxps8J5DO/biJBy/0AWm3HC16JN20KyiZD/x6hB4hgS
ok2LgsJckFa9K1ZE2a4rX1woCtsTEkGvI65gV8xwn9WbL5eYk3r0NtwDyT2jgH4m
CDQA6ccl6YkedhvKl3C/c6xKtYAma7v56S13edywgH7CjMYXffWU9lEGQoQIpy31
Fk+lj2hWHBURbGmVsa3DFpGiTrc21Z1MumKaWdISSkISOjo7f8SamXVyhSgF7fKb
eu3gv1ZIAFrzs2KAASirCPPi55gvdIdg7IkCCPpzIwR4lR/S4qM+b1T06VvlUn5h
bi2escKis7o7O8wfWmaf4AFAKAax3C9THFaOiK575tt8mqK6l2vKNIUGLq7H19zP
c8rWKLWmHlEpNcj7/yd32TqjI1d4x91U//oyy13pzi5UG5O+idjKGJ20ekaP7PYH
0t50VbBDMzRGclhgU3vxjf/ehmubGsGDxJzj/Hc7fGRrZZW8ibrySc5vdUQZZ2mq
GPY5lK/pNUIsSz9wno0X1/1UPYMrmQqgP5vzuwmmibUhXbGTWdo39YWWn/joP7X9
2+r0f/n+ZesmY1MwFdiE+RGXYNLib8qVQBEa5LaQ7AUmwCqQsHsWC67CgjdYbiSZ
xP9jQEtzNUouHFU7qMic1fKeNAeX8Uwk9MzXKNPHY9mpson4/aQZPRFDjnsk+44E
MsIBMdTqlzJDWfW74oAsdhxSRUSZj0xM7FvzEQnXewXCchlgl13RydOYNJbvHpok
84cEy/vA83oiR1ioei3RuoyRvMBGw7yLvNtLnm6/abbibEFYFBIvWUn1Jk7qe1Wl
MkLb9bpqeJbUyrMpuaGRYMQQ2DIRKjNn0LuQy58IWHUbDnCRFrb07nSvpbB/ct7u
7tVYbH1SZ8U3l+zkJ9KcOHLoVKrZyrkdLmCl3ez906ZXipVFSSgwTzBzTLrRfZJ9
30mFM/TcFEgnaV4jYaECD8lyxVJGXLgaPEULjN8EWTjlHf8hJSQiD7Pvb5LzY01h
9wnorI6X1ssNYqjGKaSqma96aXtYm5B6VvrhD2Y25UPkJvKCYWT1btYVgOzwiYev
03LyQgZP56qAakQN0SCwnKRsSp66/rUvUQTSMBtbGJroq4mIwpzgdURvsG/v7G2R
VtYlFduZsJzirJAgVvptcneWDm5D0gUOzbL7HvQke5gKmSNxzz+zJLgPRRWaUfcn
f2k01vFO4Uzx5H1VrB6pDbgE1mn52r4UfkYnW28eUE1zq4x0alqMFx6uJj8QO2QK
48A+9f2SgE5OkBhRsuv2//mLGJbnzjbyxRDKQ4SK1j93LdIQc00VM9WKPL8kBA59
uXwi7RSpj9ybRaKfWMCLxIUyY4j/zFAKAXSdq4wbq7FV0bHa94EJ5kk3Tg5YSfWH
D+Igcd6tlsMEN5dHVyge+wjM9XeXCLvw8Gw+7xYZqMud60fYOCb8p2w0Rk8BH++V
AWDC7LReTJCzu8Nmxlw7aq8Ih4LAi3p2WDkH/ghxt8eKH8N9jEzMdvB+l+LhX3Qx
/OLTF/Bu/UIAHjS6JXxLqWU6TjP4I25nYlj4Sr1InA4Tcyhwbb8Vt3+ZzRFt5K0S
mpXG7Jw99S8b3jzyNjKUEi7MFJeIg6wum5icpVa4uoEx1tuFN7DTxuNZjKNF+mN+
q8LQekU7m7DmJ9E8N73MHCli3zgOD+bBfyTkseXfKAcPWn07rCd1ww5zsbNpvhik
O1wGVvkjQP7Go+GFWpLinhebzKK7jJXgU1Vi5bZUGZdlsmW79tFzZafRmc5jqrzt
oo1Ond5lWorzfBzWVDnZAZFd4ICyJOagqrnrujOnmLVyTXuvPyQpHa7wYUQw3JS3
VDc1T8O1GVhwWWrmLEJu96II91qXpQaQiI71etNP9UiCUKsItPIWTQ3dRDD63VgE
sYVaDCKfxTZGDW1Ju8sEIGFdx+IVeLNxtZVjh81bVg2f2pRgCmEf9znjRSm36OQz
oLj5tQISk/3SI4lVVRxJHpGEBkhttqxSj/x5V+waOxvbEpwWxrwGFYl/CabDrrIe
tPx7LYZKdved5ns/qLu2jv+CS/zzkG1U67Op/WGK4yTGIKI9Ly/L3GPnISTr4Drn
hN728D6gy711YABv7HlDP1NsxNkO3f9IFOozuqUnMNMG6MIFbKMmf4KKhOmRJdJW
Y4V5ZSI73snh2L6IHqsVqlC+J4CUiTWZJRccKgvNQvsJU/dVZEEpgvzjANgpj3jO
akeu07lntShwl1nqTiWKDyKJkN/PZsovVWYGC9cC5wJuC0Q4MM+xKL/L1T3kerff
4WgPBOg8NPKtgzxZjwie5h1WCeAHcVyw6WTt8mUYPeFWR1NEBAiTzS3U3RGDJJHw
SH+VR57zkvxVVI/NFxdCYaG6HE1Gk8FVTV0h1wzvyltm2aYnM+5SSjCgr5JyeZcs
GIpjaYEDsZi+p2xsJeqXdmt4oOdsiWYgqUWGhyktPJljNswxF9PjJ91SP7ApOxkT
s5bt5E5MiW1QVKljBZqi5tpCPWDkZ9cL319aHTleYNGpumWm3MTpb/EKFxMd6G0V
kIj4xvIGEFpy5zPl3U3UABryQWMiOZKyqu5L1uE5EEnxwxq+bd8QRRR7ulOqGyQH
q4rz3bVSC2Tw6uBs8aqQM4Q1kXlKlEnSJF4kDPUIkm3zQh9gT2nRDwp+oxpcbuBR
n9O5M5Ya8Ztd1+exhm2sPdiRei6hyuA5ksJYBjeJdBJh5VO4M6rqQjxPVLGoV4aQ
uh346x1nNN9CNZpIP513A0L7bCCRzgqTJljh8dhQfzn+LRV3ZM8D+59Je/iUc8jJ
NZupUayZBQLeaWIxahtRm0ptYc/f3XjITEXrbOnhh50gB1xdz6LIR8KGr344xFeG
BTA+/2bG9Kq/3nDtdGMUvOSj7cDc4r5BnUVJRvypJbidKsV9PrVUxAFaPQipbeUX
8eT/viVGxVHrx85doMfQr3+4EwoFT6gUYZJKFoSUDGO3K/RgCV9UfNw2/KmIE2Fr
ORhO6COYk9LULYxH0ix8g9wads9RjlbwFjSkGu7eooNylVtyHz01yS00w7suUXKc
lSLUe9SNFYGw2uHYaohARXCiEZyzu4UMWZY/mkYM7oHBWgfqf0o392hh68qG3bBv
1FCuodb00xBs/eCHE7ytZf/54rnQvnq9ftIMVRKCXq53AH6G0SxvaW120Vy/7OzM
Pe8ebxt9RAqAYJ47MDH7kHVPQM0RN+8yyEs4cPaEezlLdWAKGR3/ZgQa7UJ7rM0q
1AulSUPCmNJ1EoGRuZwhmCicrnca9pnrFvIwD0ES03S8vhx+WcjeLjCjvTZ2NO5K
wec0LsGUSfkpGvnwKNijKDEVLVw6Z8GhwkigripPqo00QVmln+eLWU1uSSG+ETzS
hSg58J4apRNnPlQ+sktoRWBdXrLL1pwYB+YHh9+cMNsaTQZRCUgI/hMsdoWyIbhQ
jgRky8ZbLykGWaKouKzYPKSLOGwnQxW3Zo5TOolggAOUfUJ8q0qvuZadlWXQLO6z
S14bpkNyggSYJE5gTTtJT6qqO/NcXiANtlv+5V3ktl6Hsa1q7MS0iO6yt04s4phm
oKzoEWnHpmZf1TaHuwEuRUpCTFmWjywJSAsyB5qNz/Qhg+TvrYgyW2F3m3NQMfV5
dMCnFQdzz0fhHPA4LorSraK4dQtGMgAMClH6+fJoKRptrWAXFy1SWBgCWnrqPWN2
kQh7mIVBT66Xu70dhpFWOZOYFz7t2LotvN4y8Ik59TrWsgfh8xIqiI5aJNKLw6et
mUSVa7uyBalCUcF3dDWdp2qjCkQntUcUcKe65RAqxB7dfPvj6cWPbE0DATpo6NhZ
v1olnFcthkWU7qpva/FCRufZIPXyE63FY8h9QmVnhQzMUbPCQHhua44ui9nZzmnq
OtD0MzL14GmEb0e+s/hgUWhSgN7q/4XCoWhdVQNl20XjtHqyjnAYopquQWvrNG1I
8XQPpmTyjaOf9xot9wBmaDw6M+O8FsLr6S/EMnvXjtphWXZaaZdCjDiZ9cVWNZjF
eX7CrsTAPjbo0Kdi3hdaOuBuRN2IOIVoV2lcwePPsTa3nlSD0UZDoU4eB/fVMsE+
2Dkw7TsWkffoZDrxgl5rJBSnVQC/0vOFi9oC3WCnFkH3TXIf9b8t45PaTbuQvU7l
CW2t4ZRPo3wxjof2pN9L4LPXLDjRCeLjFb3Yaz0VG4IlosWnWgcS8G6CCzW55X2a
L/jW1MW69ZjkrQ8+zJoFxTIW00PHL1UfbnzljgTnUYIszCt4z6OrFk54WHlnTw/i
XafpTKVBMQGctJQ+bumkGDQ8HzyAATS6rWW4uryM93x7fxixe9iby2Si0ZmkE7kU
1IiNu4g0Io8ymZH5TgodYssbMEoQAPuC2CEf/EIgixkAKMIj7kGr5Nm7LLflA5sw
oQUY0myr/tcIujHqujRu/jY8UbloC2CcvnxGuP6K74eqHa/9OQHF3vJgmaUv25Ng
P4GHNvSC7mGmRBREz97skVqh5rYp7kWNehVmEhn7evUcdDd6MhvB27P8sfLxeVWe
jilmZ8kkHfvqdiExBC2wULILE5FPtupz3iGJz5PKANzlkw85vL7CnTStI4cDZtL6
JlrmpC6pRgVTaobKQPZGAWfzXHffpz4DiXge7T7Q8ktkm2X3jM0dmzcUyx9i16Ev
qtyFBuGQhYNNpxys2U/WPYSWEho8E6OlJtqw7g5X+V+wVuKWPH0UQXsJvxsnQt+w
nxKcBlN7Tw0mPUi5lteBU11i0iXO7DDBqv/Tp7ipzWU8Fm4wH256dmuEn+tzfwp0
yKgntDqYkAz7Iki3sh1Gq+b8mRL4eFSXFZ9X4IzB8ESQnGXI5nCIYMu/tdZlFPrB
dI3kHqF1DWZwEvAlAxcV3STIcAiHJrhc6J9SsNx4qkLZhrQtn3ATDeZ6Csa90+H2
ajH518i/QQw+QebS9+r1LWuyJi9EUkyCQ83xZhBgk+gnLuf8qg0ee0+b+PE3FePx
XWtlIcR9Y10kxnGFmftgMcGCT8KuMg+BVf38n5n+EOt3nW7DfEjGsty1EZOPpXt1
Yxu4CLaWsW+rWCGSJhhZEVsJ5tZfH1OZRCpVNXFAizvoawv68tBO20z031ZUAewt
xjABnCH1oY8dzd3KXBz/XIilwAeJawgROJaipbAUYkc5ASf1Scnocg97DfJffZqD
GLgH5sYQ09B00NHpGOtVw3wTJXH6XAEtlKpFy9ZOZMhL4z6PJ4SWr1Y4Vwzcq3LO
8cwlt6L30EEapa/KJMSRHUjyYl/dd2iDAuBTZi9gya/3ywIpXF8zswZ+G+ir52AQ
1ndfDQRtQ4zXwZA/AX6WGTVRlRHihlV4zXzHPt6PG25UlGYW16eOHFZDU9alSS2Y
LkK5YdW/qLymC5HezJKh2hhjS6zElbftjSEJ44JHlgZ0Ov8OXg023GWF7ZAC3dwE
4THvT9cn3BKE0DayNfIVK1JlaoXlTMtVPniy99rSVHaRd4dCS4al43XyVCkKYFmO
bZU26izgzhz7B22ojHaMeIgdR4Kz6XT3v1r/RuvOVMQDSsvQrput2W5tCAtkca8o
Fg9SgPSaSmcDwuAT+B0GAVl6KtRT5inw+p2dzhpWgscGNCTeZJSQjW8okdHBocOK
iBxRxgn7Ad3RoAojL4sUDfZ5YHvNt0MfVJEE25HQ7ySjXaI66Vo8F2wd3fvEWR7+
x40cUqh7EKVqLZV0K/rG8iUYXLfOi/WOgHsESppSkWR4+eQQqvLvxftdfdVOeKVh
VDJJnhoypgGRqrGd2onbHcMRvOgzY5adpF2sX/XZ2DCOVpG5KW4n26NNeetWI0Th
64A+TNDtAGfu+J3QKSLMf7eT7gFEeu7oEFNnSqIwPifOYvV231xhCJYxt746uMS7
asHMdgk9C1Iu0jkwqAg96rfbvLsEXc6/nBDWMA39kx8/eSBl2BFYB1Dyvs3drONQ
2+bb2zOaNL/XdsSJQ3zpdSCqPuN1QCCAeXrJrdREl8/tpaufEgvOqPrhMQEQroUV
aunaL3jn6rI6/x0IE6rbBJHBJGgk3Ll9m+RE7dSAr516h3egTCRJC2TOT7xgHP4A
/SxlHiHQ/Yo9O0tuL7nQa8V1OVi+05/c/yKLm6EexLpRFceT4ZONzlFgoSU5JuF4
Lv2Xuf98nIPQwSRg8W1WRAjdveRBiTtRSlDvurv8QTCFKzeZEEWoUoS6kDMf1kQT
dI4iYTUgs5sUl+raRE/o9XDhDSJj3w6agUQvDmSAwW+qYBdS8XKKmjI4+S8btv0s
qo1CO51fvHO3onuSngKueR5/U/GqYOpxhv6q6z7hWWwdikQXjDUkhyDEog6iaI5O
I1FAvEJGl5Ax6WAMqW8rhaT4xP8Z13Z1GgFzVuDOO/pXtbVYU6zjfPMC/ufrSbHe
pyYoCLohkWGUTXK8fIvml2cKU8gK7UhOyhfswfH6L8AkkZMCQOxIczmpvxsGA9iu
FViM9IdM5JLOEhctXtU+3h3MOy62sss6vTa11ybIPy7IVDDCrdIKzw7b71IXRHlU
jQUTKhXdPM9c2Ti+SccOSDOWggqjZ6pvuzlu541kBGAQVn3AhAM2bYdqvC7Gl4O5
T6YSW5+BjS/0tyVYXq3fOvQa1KdZrW5uZTwBlzKzze9Eu6z0kx1XezJxEurso0EQ
ejVubTIJmZbxYUX/PInF9J5YAtQv0+9425RiMsLSI+eGFjmjQkrxHn8By0mXLJLQ
n1DsKLoCiOvX4v5eIhub4beWKcaXTphoBqEO3xSOqcH06/b4Wghyoqf3M3lKZ3Gj
jetr1U1JIQ4R5guhkh00KCGNkLGECMaor7EhJn6RxVk6ItLgRVsdV1oJsofqVQyk
l4NAFDKQXtXMupSL1HqtqSfbEcNbuQbVYNM9IfNX3H47Vq4fIh/rKjBYLHVeeD/t
8HhU8Evuu3VrqImp609nRkSIMWGVEYA2krOL25VMFIMa6dEum4+RaZkg9kzTOQxn
ytccfR4zqQFRcG9aHFLR7yA0RCU4W0j/E8Y9Gxipsy/H1zyZ2SL6i9jNQY+Uk+Jz
rIpgWWwMrQ+Pke/lWB33zml5+QvOtWqvoO3Pxjuuy2zcsw9DxCMDTrQYX9D8HyZD
C6YPcw8QiHfvjGnXkxOrL5OXmjn+gwjqJRSUfuw/mcKmXhS5gwsiuqTYzwtpv1qE
TnQNAnoJuuIFDH99Kb9UozoUsONu73xaY6KoREJLIap2XFYbiRdx8pRoTq7ybUif
JxGmNRSCe9CRKZqsQBIOp5zZ4OB/whLgh7DdgjofvDLpAy121grLnYdcwr/e4BO6
dPQU+Qxvy6H8EfFe7a2VO9RqUiwVOBFwNIYvHBm+tbR+Cjo59zS0l0uSAPVZQBCl
72C7EJPGD9N3lmqwFzj7QeIc6PCD1cRzZFqKbTrealbMd2Uq0X35QB57/V0GLwMV
G1jDCJp1i71JqQbAyuDWXAwVefNYWbRi6mIedwlqesODkOMfYtLCAVPzZO+RWQ2Z
MaAlAhkA1U6GXhIuHqLX/i/uv+hOfQ1u6mSuMuBQR7Gr80MnrXz9b3o6L15nliat
ozfaCFXrO0ED4nsH0f3WJmTCQQkr9afE0YwrCqp2Fm2kX1iRPMD/wp3oOtG8Yqyl
z/1iZV8NKMvXRVZq69XQTpRBJW021YmYvZlWbRrRxRHNU4e2OTIY5hO46ffAitkb
vEHdfTiF6Yvev8YVT9bQLxXtp29KOCF900R2bYNFBkAliBCAbuXAPPRCSv8eJ8bt
2ZKQcwyEaIixFoomvCFXtEyouDq/ggTkd582wckP32ZamfIEtu9zGLf1yTh8QBq4
7WFnR2Yfhyt6tsjkt39okKMI2K6hDiZtHK3gznvlf9RPMzh8XMlARbUzGmFObxIG
2bFon9T8dYk558X9NDSStvfPDVVo015LB7ZOwnOoV8uW5P5iOW/VNyuiKABNUCnt
0z+455VNvZtSfZ8Z17yzAE+hHdmSEaC2n+jbvkE2Vn90MlnMRpBloTa1XsyNGBzE
2QtRV7mTww2iYxnH95Per98gKdCVQEAWiSqJPPUB/YV5NaxdaMHsxtFZ3b+Oulsp
FRYI8DozUMo/FVh/u6t3OqpgHlHYmWUmFePN9rq/DFwQ36GdhAw4jHKnR06aAIov
6mqyzEWw59dS0hRPyyfJjWgzpjHiHyOMqLs6tXOf1BIRA5xhEpFkWyyBRkml1DNR
jGB6H75FqMue1+KV9+SzecIOd8LaYSzaGOZzFGiZZCOdil1e/zYKS4pI4CyL+1QS
ZRYD68/sm+snYAg8PkPmG4KnNj6Gay4NGunQQy7RYmslYkg/9vzo5tY4uAo3GQ5U
dUgn5UR34UH7OREfJt+X6hcXLluRlWa/tPgTIREGljRyzEibnC9REFWLMg9Bdp0L
hEU17GVHpTdyMxt7iI8x0K+d/IDZRZXI09exB8/6AR9TMBBcLdBgaAYwctyFd40J
NOBMFYogLhMlSu0oTRaDu5P260SmarzM8/KfVIpXNNcnJ38TkDMbYpOGoOHJEUdO
I9rX9wTDiwoLnKlenLKdYdzqE80E4VulVrUOv60/AkFSvggNjyXhP2o2fc8AmVVM
Tzy0QB25HGA6qOhPM9CSyseQ0Tms7yB4CDF/76WspMYU2eqa8KQHXUNMgsbIuzFm
yfGqst9U933lmasVkP/2HIROdIGhR0zF+NmcaQhBw1mOkcp1XRDCdDuApmHdBbvt
7ajYtu0t+jC44mMGX8/tLERzivUQW4tFZjPk5mtyW4XMPFEcQNH7Dav4jUf0Uv9t
/UlSaXp7gJAUolqRLT5+P1GNbKjh4GiqntVRG5zTGinSSuFzJjKDOJItDwkkUYyW
WLlIk5ZtGNxSZZPett6lzymkG/osR5fMNT+pXbiXMLVNHtb4uzf4wdgDszGor+49
PjJETdpxk0KZ7BH7PntqrkPBkiJmhj77dRGYLUToJ2ZK9nrvp/LhGe5xjCD7o3Ow
N/GbDO+Fjaax1R/J0v0Xomt+FYWoTyG+xsezIRnUnTWyF6TV7gDPyqACwkKoA/uj
WPtxDVkIg8BVX+2qQ70t1t7eFB1gBaYiq/nJmRm2OrQk0ih6pgUINqcF6kfI46+S
wgij3RjU8ezlY0F1kBYUfvxeyIK6uT5aR4J9DqznA/nPRzvyFIIBwTAUC3gs/4ZC
Pt5QrW+bFV1SpzpRDvbYuyB6w+rYMm+mUDyMJs44bjyJzmzB9SlB2c7UkU+uoJOk
uGT5zajNvsZ9YZhlklYU40nuD0PZsdp0oHotMisLDgLVVH+ydXuWLSEcBI6mVmlQ
RrvICRk1kSTNFomqgapY+il63+YtaIYbjGC1b581X7QJn3xpqjH+Z5kAz+R/sqDr
q7sBEltZjOu26BsYbSli2A7Fz4Y7UF+b/RUDugt2ibr3j9nGVZdgQtDx/czG/bqe
knxw4FCadsUmwxtaX7g/zd4tiecAAcNQr5lxuFwZbvmRKF35llIr5VJFtC5cpdKj
9jl5V34GusTpXXB6iGTqVWlrHjMkTyKi24U5lJG6xbdYtL9YtD/bWp4n/Z/w/Ysz
DneBXMKOvrCk7E9puhnmR3mlqigqWcBQbMYKcUhwA7OnTgliUOXc6BSVPw01KTwN
gGuF9qHUJGC4khDz3+5XFzWeTqrux2jFmOv8R+98EhHFiUJysJmNASClr6gm49sU
1hvIbQbvLuhuHezlSIlUCp/1ZHQ1Vy1d/C3lSme1JCYV9SuIMyZErdo75LXMsMbN
+pGQcnnfN5USoRRIqJSjYUHsnTo1aC9Ycy9xGqo2HcJLDIdlXzKBOVGEF6pIYX2n
wv5822/f9wU8VFz6LRWXRMciDD5/sjVjNg6J+sRqHxh3EZzwCER0TfY0d0igTpu/
AqL2E+gM19vFD6TInnM74Al5pi/plJd0yvRhbkZTG8CuuP4E5uckMOSEihemF6vI
2v0oBbOgTP9n2oppXTFvJBACLF//nCpOjb+t/M9ICMKvJjVaVDQ0yRyaGW2dt33W
r288EwOBmLhq4q5LL37yJ1xzqbL0/9RmqoileELNoy6ogW4ZZ3ZNRCR9aPmhr3Wk
J6/GWVwYOo6Mkc2tbfw3lCePBuhmGVS0NvMRbw962D1UVNGzgbLUbkwvhKUo9ddB
Uzc463dLZ/W9XYugmw8OAEHMI3K600D6jAuA4RaF4hqTF7kmdRbibsKyoHh+MPuw
4fP6HLE0bPI0Sq6ra+/VU856PSbbw9ICEtQInFXV0u448rvxbU6XAugHRq8J59kb
mCi2ezt8alQOLcsmOgbtqXK8Ky5Pn8HjCWM+nFTLYj6E5SQ6YZquD4c2t7At2Nm3
3VwcFSRtcbe/xSkAR4T9RgeGMMjXxnNOFOj+BbNq3e8L0t6Jmndf4vBV5fe6Tgf1
tC4lK4O+Q5g3oU5/HN5YA/AhNGQMYZb+J3K5k77LQCwlteKWJZaxS/x2sejaI30b
TkFN72dE8EaPFFgcugBAAMRZVll37c0KYzFPHdk1/tzMfzeGI0ndcMNhdtbl/KxQ
21LxIlIPFStPqdAyLwgITBnK1gTJUFNF7TAx8CM5jQNjJtOvpyYLN6lNvawUntg5
y4NR0XbaAJClRV69cr4XDvq8Ais35g/cyGGqqkUqh98eiCEK+WvNkqeJwSCHAcGe
dwqyQwpm4EUHnUIhynHXmS8WJjT8L4UQtrkwFr5UCmxKR0mltTcMasjNVrXaBiky
9BKtmDRP4Y1Bgp3XYDxMyD9OdP7mAPk0aFjznmOkuyUiDnF5vjXL9TQGNnUD8qaJ
qlP6F+AnAMkWGfW2fFSJomqeOihz2PkQia51HfV1CIukyy7BEImucb4pczJkljSm
ChaH7dSdzPYhK0bg1UKkKHz0t+W/TR0XujT01KNM2c9WslIsaWeqyJ2DX2GHBKQ6
rfdHVWHL3lzPYBaezQK9Q/Yt2KStNbcLpcKixYP5UB4ueST9O8InhcibBwrUFfPh
38+HzdZm5zFm5qhrpWZ3BzaxXsENX3Hc+jBjgYkxSIp+ruUk8n5dXuBhgdktOgEP
XpG29xvP1sw2IG3c/G6WRtAP3QDhJdMBtsCrqZN7PF09HdJaR0c98LDqsbFRq+v4
E+KGAX5T9mMaFj3Fgmo5jvyJ8K4OBxalh0CeCOGYdagEz5IAtMFjNKkmf0HL+YP8
lw7SDr69PuaJjreCmVMRZJYVphnkf+0Udl7vLWKSXP9QIW1FoPPp76q7AWAXx6jJ
do7uoSPcupqEBMGgHaatXyqkt/AsOWOxuzoPZG89iJjqxGVQfhFANCYSbkL97T4j
niuDBNmTTse4t+LgIkYDudDYAzQmjGQvnCc/ZtEHP5gSSQkFYiKciX09UIgqTHE1
hp6v8Yr6f2DIuclUzkWrDLGgRLCxla7gulLHttH7tyR96ab9ipzLgQzXP1HvltUs
FWJY2iO0oLM0wKTNWYEhY54jnnpw073YZwLSYTl5+d1V+VOYhHQYjS3jrRbmdmi2
+Dw+fBO7DpKcbOePvOwZvwuJdhTnPINTVft+4QRBAAJ2kfjYzgtidcyny0qKsNND
KzIMMxP607R/6VcBkDMo79YyzK5UWbalULXusVLBDrh7+CxnsLfbj7FIjE3aWTeC
8r/k+4xweVDboiS4NolDqnAC1C6wsZ+LeIp72UD1GX/5uPnrl+DIWUtb4FY0MQ4G
geMh1CO2N/rV8vQwXzEgJWRPCgD0O1S/VCaqjxJlXaqxCzdq3E1Pc7sURQNYi1LE
E5Kkms2R/H7dhdHd0XUZbE9AtYkvXHSdQTGkgALyP6RtJaAtHwm0iKlnMBng1b8w
uq3bEKKiS49zMp8ErP0LfcZuhP+gtpFiCmHNf2vVCmGnVyROr5Fg4lR13PFzR5ok
ULvAasmfOSxPO/vK5TAkm+/MWFk8Trz7c4PRUxP5GDLgUeZRdxx8XDHYzqXwQ57T
uuKnZAZceWm+sWamZ7rHrscGK2B9sBeDmMwwzNcYKWz2kXeIMXs2ySDnqRPgNk8+
FaZqifNKOGzG74zqKT7DQNWBDcSaZzTNF42dbIUCT9IcXsa9SuJZZGLB+xdOL5Dd
k030js1kYC0jEc6lheH7NzHWm42EMqiMiN/cdVlxSv6rkfnLOEMrha6bAAamaBVL
3ozsLhkQsyEwb7Y31UTKYcU/EhLyqoqgJ5XiGhqJTNvh+rQulmjnVAokKZ0bwXEi
SC+khjY4uXnSwyEg5EbUvUh04oc4UoQ7doAOtuYUOWJHztOoW8Qr7F7i+WbclPJg
eDI5thqT3XbmPBOrE/ibak5dQxLk33pikFkAHpD3/TmkiMXr07Xp9IIOaHLk6PnL
r0Sszr9CcpgfGLhl9+o8C545hqBtxw6BdBwuypnHKPD1x7ajwG6YbrzvF7wWSD/C
1BDbZkhSwZvLemT/YoPE9kwfmpzRvxemsjJCh1gtSjeXyWZABxYHhi6vVYSdiuzi
OlglYsigsp5T1PoeVSOPjO8itXm3h4Us7vIXxsx4hjl9QQNZ9CQU2jwLHya0lhco
jIWPGCcQD57Oneh9c/Ob1A31OdAkxO7Jp0qylxflpXtNjOVxU/TNxQVpko9oaDTG
qFRb9s0CWedZDCmxkhV2LYlk1ZKFgf45C1WO5XVQyBGdy1uaD78ZQZgYoy+c/kQd
yEzHyfcgPzcx0fD5uhFazkmk9jfL/seCrbu9GQbQob+6RNebo2B54GHKoTJ9ehWU
QhhWM8OjTZavptTMUC5gYrCt6ILA/HR1yKPRjxsDK3qnExeNon9dADTd9jJa76Rp
Sz1Qh4fnT4k6QHnQfCcaT1UEZ4baax0bkctGLHdK6FX4sSFKh2jia0kZLqhI3jQY
ZEMuHZACzSE/rC/XJ5fJH01evsv3voyPuuZFQ9avfsZ4SiNE84ucbDcjoGnsUzxM
VWMBdIm7SSKLzhkhw/he7hPw/Zck2ZuAGgzUbmsXc1q/+0fDjDNCWHveieI3tRF4
9xJg6Wjhb7/9D95lAxGbFujy7l8+Gdz5yqEte/9BV79QRl8OuBn8PfkSRB0nlc9W
qON331m/SsSRNoICoSbAtZVSCJgGv+uhfBOccNweOX1X2+P64Tud7dtYbRgNLIHT
DIIwhewSBATc3WIi+NhU9cUd9VLMsiybJzEL/fEY78u2+aUY0F6u6tvQw01eZFUJ
qzoI8rvKPJc5Bar4+BfXTA0uY0UKKvgSnA5TbEMhf06mGdLxdC1uQf9vdZ+wWCZg
8YHhctMN9OlxkcfDgmAlAU7MkpbQMnLCTtvRAmChxnkKjq3UdS54SI5GEZaO7Au4
11Th76JeGinAwfSjcvFx2OShxaljhMxUcYPuqsoCxFME5IM3oKKF46Gqx31ER5BV
sRa2cStipN/A8uw1RWrmBjA/msbUxmbfw++16/5hrEDJHTrwt7EEyhyWbaclSW6B
d7rbKLVPJjR/y7xqLEsVQnJZXD8shEPl5Jxn0Q0m1I4p8zWikDlutWWXdop2dXP7
EKP6vSKgedjvbqdjwWRrlzHQhNQ2vAbHXhnwZp43Q3PsGCoYdlnaJhi8T7PW+Tcc
RpDB/Cpvt8U4G71kiGao8P6cTkgSYlXxGOs96KG2NjOM4c3P6YxId0u/q5eKZ2qo
CmlBvo1HWq9X0o6xCloBe8NCJ8uveG8vsbdFuAtc2Kij2/MLp/XsQHCcaw6JX1fx
NYPuSzA7HdEvzX+o+F1fRtwjMcUcBf7NrtaBmlC5iDLJ+PVsOjv3K32y6kxP/73I
XdRGvhkaFM8sncoyKybnxr+JIRMF4ces25v8M+UxtDDhChwGNo61jGR3dPFM5fDu
bbysnmM3fTACWQstjlbtUvE0BBlvwAedPUCTwvwJXLef/CgGU3wcl7n5hiF/buHK
1muDuNTPwnEGCweDvBHenkZZoFiWaIAZzMyffOFYKhJh/bXzCHgy4n75vchcKePL
34FgKzamQvv9n8bHJXEgpPW2yJeG0dtTYEBXQbbESZfdVtSSAuccqDg8y382rQCS
YaN6rsnTynDcNj3EZ/DS5aK2AepQMbfrfapKCXp9+SeU4qFQKTYs/+Row5HKYZgt
PEWl4pgVIpDwn0+5OrKeMHFZLT092F4mfLdOMXZQD+rMATbozaMZP4vHCXh9QRlV
3NNvoDAZpYJXSYkzvp9thBVT9YCGvGP2wj/ATZp2duz0Bc1rEltRPeGLnZlpDbYW
mHYnaECDXbBAflFVyxyN6ic5Uy5eF9dgZmqIuYOC4n1RUStS6tBh+3g44PtVFT2D
aa+PZ9+3fK9KNS1X2sTI7Dbz60VgQGv7Zs2MyTVh+6yRTv+i8ikPmCXg5lToTWXU
gI5aAV7jRxbkZeRTnS1+7TrG8b6QowAnXNqOUOilI78sKaPIbX4xE3IUbRMUszz7
auahBaTBsOHr3ER21oJst3xaS7vEU3M0kDkxH2C6JrAZzuAFsUO+eq8u+yN1F+10
YNZXKVB6TNkpaz2YRRjfC+09VE5QtL1H9JK2GYIIjUCs6yjxKyo+XcTCIJrfBqVW
6lFQfGuN/pkCSIU91CKxLTiqNzKRBW8+y6LapWJsaQ5GDpGorxc+2qTNBu4+vSev
CisqsaDuhOGpB/VmIaNtHvX3ZHecZtoeXvelf3BRRnLcVTGot+0nqgX4OgopCS6e
BQE1dvESHGC3k3dU9XoWfUEWPWJRq+6cvrJyASVhGiILu+EK9x1bG3Gnia4AItZD
5DLymxDRJm3SVJ6Tr+/BjAu5WXu8MKrhpXL8/0bOSRHk0Cxirf1SqoHtK9HP7GH/
mwY2kPcrBtAyoUoy7BHWRuij9UWBplNxi7P/8zyTjHbCpSszOiO73kyI1Y8Shufj
rAfblgmf7ZNYNw4GkLePIdm/KGX8PZjUZEdXbxFWodAo61sFjYHbZHB4tg23ty7U
xwLte7eQlOeAN4rC2fNaQxciIZGKqfW4KZhUVZ3gjZj3xRTvWayMaBYq2n3RJrcK
IO4vIkBlOGbKGGdC5mqimdIMoXNxs6yTdlxauhRlS1dSDeFYagrHQwHM7wPoXEk+
DKqcSiPxPEt4iV5TuxQtIZClyR/csmx3VoKza4AZI4UjhUoIzAUWWi1iLWWS5efI
DncZ6n/q9gPwK2OltKWZhZzozZ+q59GASD7t4DVp7YAGKpjQQHQyJPktWWUfV0YH
Wk0IHVLdWltCxBcmTyhTE/i+uogpMGh03RTjzuYRG+zh0wDg8SESL3ZR/msAj7Sg
R3vuFEHIlgAGFN/tDCY5CugN1iUDUS12V7OZioxYD+ArFv2gincffh9IjxLwxdta
`pragma protect end_protected          
`pragma protect begin_protected          
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Ye7+MIzMJd+7jqbSYPV4I6rigWzxgnJswWXnjvKj5M2BwBODC188/fzpUBQ+sVFV
Ns0tt8gjfpzaJIZHOJ1O+IUh5ho7lKmg60cMN6Kt/He+gXLrwuCQG1jmNNHnx+65
g1/AUzzqvAY42iMZKrKtnaKLdNCsSGsAtItdudMye8s=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 32437     )
jYxcQP5sUSqT+vDPcqbhKdtiFElnEjpm0m1zVcctzaRBKlxgKVfioGZJAOKKnE2m
EhIsTSRZgr2cUOn7AMQhXVUQTIrF3sxyxB73k0CI1cZYmBJqXl7CkMx3TgkK7cvp
74X72nMMlWBUYiTWye7L6Pfeda+Ev8gHCJg1NL14JGrAv/y4bXAc2PdoBkvuD5nw
Xta+rR+cTp+JXl2iZr/qlSehjCmUNU/424WSKRXhdsC4KzBZiV9IpPhZWD3eWuRC
9OHjSlQ/UoNM8IatQW2sNVJZdqae38yuBXjzY40p8/Ecokb0nvkA4YygIOWVRlpG
SS0QqxDcWRHiwndwvomTBCxCfO1mqp41zkvqHRKm2MORg29XOl77stoAfFEhrNWA
ezCHmMxHoTmXXbZOPlIQor67hP0w6Zxzu2Mn2qiMtGrqwX1yw1eSc3dkBxDg5DR8
RToUYJcjUrHSzNLWhNXjIMy7T6Gd5XAoiUPKtZwVCCEUQEGGHu9zRABFeas81wla
LbyRUDxI4J06oaAeHslDFTALJnDlQe5cTaxXTvxMma87fEXaKgpBlM80G2ZSvzNH
gb9VIP0CVL3oxIFIq53wWc2oFlIdw5n35Srd3fnU6RHBnhYoBY5WAP0f9cKQoeDj
Ry9wN6+V6/2cYNE+WHmh2GFNnYoehXGGIz7u0/1CZ6/mjZiByV4h1KXzxXNKzbIG
8RHW5wZxsKeRU9IjsTVw1oKF1eNxq94UcJ9OcCzrSgTyFbGBPxHT5VjxldFB3QTU
THVcxJZKwEhpo0BsY+evlNnGzlKAi2AdMIfGdAtS/Yf4ZesnsIn2XKZmeQKKKsvx
6wbI6FsieGr0wAA9BUeIfac1w2QZ5BfEGYSe8cQbhJqRky1rkEl1s/bw+B70wX14
YxL78SVwIDsSTSxW5Fp9D/16f5+d+ogq92hB66lgRSuRtl0sTmjg5smqK2lMtzM9
Rr/iWk8dkitGVUd8uuhrFmw7X/wCAuYB/amMyDZwNoy1WrqyWjhJuuWr+uEm+VNR
xY/r96zuGqoWmq1fLeHOuO7zRqPAkgyJgClZTY4GKSrJgW7tKlxtV9MvdkESsG6C
8wJ13t3+2rePQOQTss9ZwPX1Zveq3KGW/Rykq9tJ6S6mzuLX7xFm4TzVtgvM29I7
WWSo/DmJfvt2JMp11OCXfvXwX3dWJxyVRR9C3wKChq8aUTj3hhS1w0l4FesFYdU+
RtQaA7sshmtnHcWGH9DcCQvVAe97WCw6HmonNoQgqtIs3zHtrZ5Vr/pWZnyxqb7G
U5Qxj3fL3GSQVH+g5dpwQ1DflcJdR3OCBwvbt7EBWwVQ+WACSMQZqFgfCPzQwmIa
NF2qwuZdPdzIs5/aaINPSdNGbp05pJIT4MU49odzRPN2TIN+PY3NqkFbnRDav2mo
jcW4xXyY+CqklVhAzOmYI9sB5MdtIoa2KySFuaSRbdp4X18Uykmb98LT8dJVSgvg
sIacGwEW1BqLAjOPSD9DUFUCZK/iuPGtoIzDWhrFNtyaBwzgxFSvpooTMSol1XXd
xjN9kdDvs+1UYaulvdyn7TI1Gm/OUqMDbIWaLryO6c0LjMO/ZMSXL39PKhZhn8dn
`pragma protect end_protected          
//  vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
daxU5QuIaR57Rh+QD3eKssrSEMI5UTN5xpf+RmoKnX9/TjAP2Ztz4DXHlnKg3G7f
ypvbnGzg9FWPES9ak29W1ne7OePOxfFs2RKWFPmRfqVd1OidCViblfZ3GMx3Rs5l
n8f9suS+HzPnfNzvthIKIaViJW79UfxRqaI0T4BdA6Q=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 212304    )
Hni6DLGbDA5TqwK6742bsQA7Tzblko3WSSzkBhl/K+ODKRJA//mZA7QwFagG30A9
VnDz7CRIkcwN9Iy+8dn6e5h30rZ7AFlhC6VNgdzCEOfs67G2JIZtY3YQ4FX4YMoH
ve7aegqNKk6COO7LproN7naoNhm08Bk7ONWMkMNDyneLhLWS5fuHDhieBM49BuSt
gswcdIMXLbmQgRHSMUBiA+tQ0P2f1fka21OtVUrv4HDAjo3ekbTMJwVJn9dXVp3V
jMuwdm4C3tEH8QCIXOaZ2g73DaZp9hAFW9aa9TqQkUjmkGZwllfO5pxhkSeF6RXb
XPHP3PeIsezJfpFA47/d+DfWXDTTFMp71jqAhgM0vPv+foHLk3cd/V2tiVrisx8X
+2L9ZTwhrES1I2DlTuDdG6fGXyTkc1mp/vfhbBlJRuke8YTkpCDDIafK7GDWLUIw
mJO7S+nmLjVe+h4x454GYLPTlE/olDtQpNRdPHaNt8h8+MoBZiQPqf543mDS3nKD
bMhGcAKhYCOWmm14gl23zT0EJXeZLUjw6Xiq9yqv6Nt9FMwqbbcyboR5ersywmUD
WX/oyaA1Fi1Ms0w0k4kfnDmJWzGapy30DDeRokjT3pYo2EOfN6R5rZBYoZZzNPaM
PN90R5Le92OH7Tp9331+9Xk/eTgH0Oc2uYyQDKEfDIT6qgkcHF6jIy73LtZKgL7p
9bL2h15prhSUhD4dsul3t5eGR+0nwCQQTWQ2CzuGMg6/B7VkA8pEdbUkKsWPHJ+4
1j57lh9Acj2bNTM2JeaglCkqfkhUxpNEO9WuDi2Wy0GAaFiGDUhyvIlQSGMV+WSc
0/aU1RMSMPoDDh6/QVqeS/mUh/BXZF0GFiAo0RUHg7QOIlPIxj0Cg3DjbycGR0FF
C2wag7jbbbk8KXfb0yOxHCIWGKFHUpn+6LyUNG7TgRzCWZaLl+Gi5q7kicF9JW3s
r4+L53XosHqknhEqpoR/KpZzxFDHHDqFMc5A+/cM8K2w7+epNj4FM9kPbO0QJZ58
ubs1Txu5JX8nM6E1r+NoKQ7wFeOwQPu9/zIPOSB/y8UYKCN894UM5dCQvInfC9MT
jDazuu3BFyVbjf+NUFQvX+5geGzzqYI7V/UmOeiWRbkVPaI0izHiUdo/Iegd9isr
Chi3JhabyMIzfTyC64+J0I410QQkfYQIxcrg+jr7tgNQyzC0kkFFd16hichhexaH
fFxXrItmQ10JPUYZJ1C+PP9VWh/qkVK7Cp2XuuKJ5jsaMDiFk9mUaJXdVmop0ImW
rNmYNUCy3gkZZKT03Ie3x9s7oxU0RJt/SzSivP6ZnhA9hN/vSXf2CF84J5kOO+Uh
Dsvp48a4WsQcHxib6pF4YW+CLfXHXXU2YgYtCIiDHUDImF/mleDy7I9F31JWzL4E
iwHvXrH5jYF/ndOABa+pVhPixqjQtC4wdXb+Ugu21RlW321jAzbgLLULClErnz+p
sZzYPMR7udWIZffSO169JNUyoahEc4WVcCVz+zSNqtnr+rqpDwGqvTkbcDKS41jx
bPByQWIXgA7Y0BxWoXwSUKgfO9pVgjO/NInYwGfF5Tgjj8p4Q1LA0k7vnyXf5xQK
oWvMBeY0kphwkYPitsQQlJCrkxCcODn6ixk/pS9opd8uoZ3Yps1elxSAHRwWOi/R
a4v/fuDGgrDD772TGkZ0FsdhVxb0jvj96U9U+82zEsGemJcawBONRK8gbKitGdmt
wMprlcLhHVDI9zrlLR3mN/0gxxccv+rAsTZPBmmqaSJHgge173uMamAGg4qvw6tz
HXiLgiLsq1Up3DNqa9Fxdaol/l52I4KcPfZVB3Q8+v7VariSh8Zy9h80NQmK/p3L
Qe8+SuUMpnWqnKwaGxJvAFKOp9TRSjEFzaWaxgU+9zN80SWllR6WFPQ1tkdUpBl8
v0Y1COds4fkFuKkPBgvH+zgQpteyKyp2tfYKiT/yUoBKQzi5jNrl/y1XVU9lP4Ik
d4iriAQmKSzRLI5y2lfYR8FhAFVM58u1CkuIUxzrSioLe9spvSSgxay03YpPTae1
zipnUbHPk1Qut+bdebRtSQgR2v38hCTfasrXK7Z9Znwo/XoksrZnnJS0oErKdYC/
nIiPTkek23fg2Vf+O0YmWG9hek5eKeAj3hLxmodR8bD/31S0lR27fHTHY3BqzxG/
jva+cOSSj/bsGw8bsijVEOD5M7RZTxG7acfGm12pqf/nyhzdF4oCeIJvQzDJTPBj
tuoAqgJFudq0VSGTD4QT1wMGHfy6l4FKX7VawEIR63j3yOvTPNODjJmZ0GT8DR4H
8cLjTCEVnHRErE3bAyHq5B0ZeZhrpwaINK7kNNDMUsIUAsrTLuUJNFbCoFOa930/
1tXCZmfqMJUR8YCzfArf2witkYDun5vbGaTaq4/8bi07ocshtKw9AOrsJK13FJEU
HXAuzL+zVeYpIgnXa06ePkuKK+pVqLWt7KDkBIjKLc4e58u5CF/gPubxYD4F2EKJ
PqP3ECsVsJWsoVVdf/SdwuK07+QF2eNWB/jpI+pcvWl/LavM4jbTTeytoeQ+v3WV
/1WGhU6x57EPjD9y3UmsZslTPFWfbmdiVUZX2qHMps6C76heH3+gFrjJnuBH2obs
XuW3MxUF+xLdDWoJP7XMVdgEPTWIMEs6TXTKvZ1kjtBLEX/azTDHLG/lNtGPSVkD
l71wI6YJ8vfgBc/tA1rhNsOk3Oc1ylvVe4YqnvbQJgKJq8+DLJrSPj4MqLAIDtbW
NW7ICK+EW/VDOC1MbgXWfFUmaKFlF4EUFrtFBlhq45X+c5vxVdw9JN27ALmPTm5W
o95leKmtL/dHyyuLpRmQr4zLcdn+S4nzBhMZJPyrRICL7eYLzDtffvJnVXhOw/D4
7gZrEu316XuIm4NrWQEyK4Oo5GcGytnTEKpCdBU/rtroDKjs9s53eLFv9luqsFKk
o0zFM2EYN6jnyiPWNvJfdDYC8+ZHUvMEAR/V+vifAfgPgvFIBZKVp80pntTGzz+Q
MT6VSR8DI0trRzOARQc+L4KnuPYp9vEa49K4g140LtNCX7FfE004vEnC7RW2CVq9
UMfbcb73KAMyklU80ByHekWJ5QXFMt6xAxdxBZNgtZr9HMR8MDh2iOLAhGQkBxkN
n/y7pX9pdbYyc8sE1KZQM9czVgGjKlcZN6l6+fjqm1/kFEzbZh9IMIWPZPwRNPQJ
Rx+kbedXp21t/TIZauc+29ez2oCjG3VecycRsN+o453ASDl/h7JTI3VOm4vhg99M
dY84Pj4ZRyWxlwkaKQOP47nICkIBM6SppIFQB38H6iO405yLO897Vq7Kx6uEz9DS
C1+MyLeFPJQSNBHZjp9pc+p39Qm6QxItVJTg2x+OiVanAhkRqw59z8JLrF1pbIZC
etCDFE0t5np4TuHIRc16QzjFzbaAzUTcHfvYjwQ21LB+QZSPl2eCwLIiuFYdIfnk
L4z/0X1OPwkH3TMjBd9/E/h2p3rMADm/N48KYB2dCem/kl6i5edSE3qaJ26GITWF
CjVoj651Ngn39+NFP76GcBml5I4VAFlU/E/fHCaOFkGFYlYo+LD4CU3j0p9bj/IQ
ObsSSOIR8FDx6fiLr1a0j+IKGBEDn5wcV4okj67V4W2Y6o6dlIy5oLphgD92rKlT
IfBLLumndzvrdnZ6MOdejjuO0rxWnTMQCAwn6gwJqNb5ID8MkLGPx20qkBeByWcf
KzzPRZsFJl5OeMrjnKniqeLy4qIFp/XSVbdYChE0a4BUc+stAa6AGIzGesjt0LhF
uvtyYsb/RP/MkIlXRvbqIHawQEoz7U1Z4SIGdvMQzpWC3i7HjpV6tndUq+Lw2smY
befTklmHIR0Olbi+vc+TDrlisBcCv4LpSwNkkUz0tUTitd8uvwUVjEt555g0aHTx
yhc1M2p7vhsdU2ujHITpK4Stk/Aef6pYliS5IxQOSWTmR9qEfH+Gswx0dCw18toO
BCJAoWXK2FcabycJLhyUtUhARYh/DHfkIKTH6u5jgGlVq1FK5XCWbeh/fqYZJv4A
OdwoLyor2dxGDW/0wb+XjcWmILuMszTBBlS6YXJOM99KBt23iWJgdtXl6MrnCT9/
93+Dw/y9xKgCJfda760RiVpHRCbDzc62Bmmk+N5Rau3j8x2FLAqkoIr8FvnKgL+I
UErLN8dcNd4I2CS+TdR1iycsqCpJen/S2bKCj04brGPz5TCWK+bOe4rOPzppsl/H
47Bmrs873rKJ4TRJ9FV15aSoYL6qwDSGPjPZBQKV7ZrFp2LKpSslESB0kbRdwObF
aL3QVFZgJW461jm8Hmr4kzNft98rYKxUnEoDvv1vAr14QQuRcpScHUQOGrNIGKZ2
YLzZonDC/ssgQD6vLfB2vR/MmPwvwB+38az58KoujWoc2TRln7DKrAS3X6hgL90C
hLa35HxRHigNnZkvxfxNq5D3kvJS+I7o847NAu3Aa7sMcEpwePfHUM2macveOSS4
F3utmMAe7QmvzoCMDtn8p2ZnYEYPNWV9j3RcM+fA7q6bXPYmTOXEImeiVA8GV2Zo
Nt7g41o5KiyJlHR8qtgk7QBt1oW3PFwxx1TaJFMCMoMfT5t38WE1YgLS63/hUEkF
XqAjoG7YFq13tW4O/vV0B82CAZzlVyhWc4DINyKQLc9g1L0FAvQwQZsrUFZrvg6p
a4vR/ThJHf55ito+VGS8m09LeA0xUrEOg4eQl5X6dh0yIU1fOl1xc3iOXc21STjQ
/wJJ+M+ePCoaZtfgYCTYiCSl+v1X0lxEFMApRgE57Z4vsI36YnWW7x//o9Axw8m3
7NQPNcpQuePw7bZGjxF38MH2w9EhhojRlsys/xm6HiWtW3aY9QB2wjICP5lkb58j
4jA5yzJMbp6CEHiJUAbbl3hhUv3QQFYudsnDNtRYCvn7e/Lc9G0ZIfECDXIJchZy
2HQ9mWcFMRFcE6vdVVnmGWgfZ/Ya7tpR7xmTKbSuCVGuCD7Pvm8S66Il4MoRkkrR
rCFOPb3gcdUmZtw2fQj4c4jg6QZ3rhhJhycWAfWyJScoBVYHlRfZrTxhbOzonSgR
C0HF1SroH4PHgPXJQV7Rgx72ZDKbbJlMEOXF5V9tLTcSCsECvCvNPk+jVfOXrAj6
rEPLb8UJXxgpFxe2DKQzWQ+6l1INru4RM3s/lQhLX2Yfu8k5lrDzHJvRF86UVcZI
MYHU+ZxJuZ4nNRQE3n4MCSQpDYvnQGOpYKq9o1ZpGRk2bkKurfav4kwofTSIz6QL
f451iZflQ0l2CgKnj9XspWyzorz9C6J+yt5ZBf61Mh1+QGNQiWWtoFIHxeDRXfop
kYEIcQ2FdCF9WEB/Xe7Od/una9PBEGdxMHrdGNf6aACa5mvaiA3saHlFq4QIgRaX
X2353TJGhm/o+ZoV1sDMYEMgC2DlTs9HDXL868KgRpjUEa7P7JYqYAqw0ptqSJ0I
qxkZoOiSGxsJqJz2Lpg3Y3Ci8qSRzvY43OHydWYEkUB3bFlL747676ZVdY3YB1vX
ri1hiE0XuCiwAKwPiXR9Qo2nsFrwFzOF1tCLnXt9fJlbFY4VLPX9fVelEqlVhNU2
DuOnB3rUKx1HUS7dZiMy/JpZEE9q2gGuWIOcbElDByiB26qjSLCRWjb2le2lSfvX
lY4xoqGGZxpeo6JOn/diwZPLGowVRp58BEwrZUfT2QGiydd1FnwJTNOkiSA9kuLt
JwiL/fTY6Fpn8b0z6WPxuUlz8tQLQAAMs0qAhYU+5jwk+MjPHSfqbQXNUcX6MXIu
/hNDpr90fFbqgWytbZg7WaGaucSNoW4C1fOpmnyjnbeg1O27oHa3O7ScVUTYZRvK
S3txCLanWikUH6+Pc4o+51RTAKK9zGiioV2B7mUBuTTLb7AaibAGoKZuGUdMTPS0
fZF9sgUIesaw/cbYOfShqY/kboF+FbmenwywmP4iaHoY9y6Pe/ubcsa0Bw7g8X0+
NXZjg0Ga7emZ8rbs862N1ELkHNqNeFcmylfAIEBuC1wpQRiHgujfz03J0kosiu0v
2pCVF5J3+ca1dSjY+E7BR/G9s8DJiU0WSqz2wDmi8gAcrtVWykoHCc6GGeVzwKgA
+K76Owpi/uQ1p38PtTfd7Pd1aVEvpNejcwyBSINpYnwIJyUucLl7+5wMz931fdn7
b7F5jy1DQCxtVw/RAodSnYmeAs/MS5CVCJ/io/nHKgU0h9ypiQtSjn/r405L/xwh
Aif9XUVXriyHpUBtjXd9r1CCHUA1eWWTUjsR0mCLBHzWzPh8MMe9MAQwDDlnTZcn
hfGI4LMrRF6qhnS8BqBjerDEBdhrr98U7kD+No9cIN3Vi2MiqWccQU+sqHb6lvNJ
8I9xAlVfzIelyL9+gQ9MsKrm1O5XverKLrVTAsHBL/fnHAhJI2ljdDeTKAvqFPAm
NXDQ+1tNeYdQdHGWqP3eIwENax9sWlvcHms0FGLOwLBfrwGCdKFf8Ee+90HXTm6R
X+WSlcmkMax8HyQAHeIrkJuHw/BiSXyIUl3KcOh0p0zQUuuteF33/+jzZtO0h1Ff
ZN0ifLa8Op9LbgMb4i41x7nJN/wQssazLsfZRwOfJgnlktxr/2PfGsRC/L4p/TOS
vZa4Ifv9dWX0z0GXpksFXWwRqgBUz7hmemHk3GVP7vsy3QUHXGNmmZRaRuu31Esg
MlCwiwmaqoWuqzVAJXT/D1yqB+e9TvpLGfVW7cKQFSsXfNQ4hIRtag9IjJn/SsiS
/LTYy7xVRL8gXAZog/OJzhZ7SBa5fNkChQeCaK+asBpW0bVsuDrxWtdNCXVc9808
SgpA0FXXz6FloGO4oWD76WZGt9lTZjFo9HXtbY5EA59nSu/MmtCMuoPqT5N0jSE9
kMmx+JekrMc/uSKFneCLsV864Rd0q5n7gMu97L8I334slUSg+BMwuZKWYPuVj4Dz
OL1ZBjm9qFt2zGeX/7eq8FUASdJUheP/6b61H3E+ftqZ4n63KNmrNxQwtlCyu7Dn
qgJj9ZDOoF4rCDqvrvhUvQqnIBndr9CF7iDIABFFQXSiZJErlycKXpOA2uqw3K1s
EJcW5xhnTASFjGkr4Gi6/gFlZ6xarvZso0Zjf63CFw+Xe4DeHiCx5v1B85G7ohq4
IyreOEBhPu7Vb3RknZJUPHQHbQwEHQIaOmQVpeH9Un3SaKQfYWKVx/IEcUQmdRZi
KM5QlNr7qM+EoL4jFYRQT1gNSDq+gYegCtr+zVTmoOO3uVZalvjddfO1oszBVVtP
qBhxTdU9QaFNpo7TgxFSCGAScmlKWg3rStwa4S874IAs4ZXgX4vHGc7ZzIo3WdIj
HANMvjc2Ol2v5RV1d36zQg4Qcnbj1qS3jgGmjRabUyjCNHKJKAauTr/yLI927L1I
rjVYFz5yA1meKZ9pZ2Z8hUvmUjvzQyjZYt4MN9eMu9SQJagvGsuVNFzRP2Q/OX8C
P9LseF4um78OvFQmXADwEKW9XlblS5j3XcNe7Z2+hUtC2zA0Xtb2mF1qH0PCrxQN
gAvIIJ0NdwJKdeNWaHwIDKywbiw0PELmNTdIrx88m1VKFSUhqO57qtt4fYVi2sS9
0KVPRjsbvX51fx2KpqHibOaH/bqV82rX7rMwImcjtO7VRto9mvzN2rEN2N45HgGk
Gw0G0E6nCbZfOTqoQuCWoEtn+9mhFf4JiVeW1bzy2w1qowoo450wCVS9k+b7l/l4
7kDHL2RLuIe0zQWnsMeL63itHATHuvHmuU6umwzP6KDK3QovwFTExKka32eKzyX0
GtOCt/097dXanYsVI4XWv2e2O4wyS8tLMn8p0DrNSor5KQWTgXChCmhC9YDyDh8D
REzGhq0tJzuuhPlb9vA1ya9AVctYPujM6MIXAKo7CmqtzF/9g7UBqbHn+y/F4V04
9/MwRTCk9YE38+nufYcHSzJ8s+qJH/VwW8AOGUFHiE2VKUm1/i5V7pnFdg9L60yk
RwFX23Epm7By6qkL/5xlUSJV+KNXeK/6L1dsHv9zySRZuUZLwITs81REnwFCjsqg
lZz5zSRrN8jK4KgaZIAHXrrWKF/tgffs1Nb+BQvl+rPUIEQ47gRajnl5zGnxdBSC
EU8eIZR6xg4GjkzAThFIAfZLawYOz1yDRsLN9imUfCxd/a9sTWQzCSF1uF6vrIvp
mSr2EuI7Nwg6WAzJqr+Wo+BUf/B4/TE++/s971BXr+tQIsCmXw46g7acaLT79Yh0
tLW/rxW/J3OHvjaWyDGUgoSu+AZzAvWN+sFYkxWVGXMIWpxayRnuvIk+xGDTxhLh
X/Jw2kTcjTUMeybkVZ+LEMc3yrdqtkYehE6rshdy8+JBggwjNe9V1H8kyLQ4w+81
R7OCJK9vV++QdCREwzzj8SZDMQiFq0fjJD7IDqnhXmBqObXyfwkHqRzhD4E/g6fJ
qcmNDLFHlseNmBbKUrsvIr4AVmJAoL+RgWTxUuJ2/py2unIZZ/kBzPeuvw0PxBpG
weg/Ru263aNkMh4oDlVlsCVUs+cr42BD0uC4GmvCkhquLq2zi/t7UnkXgJcGXN2t
rKVFxdWSHIP091eb6bZBooJ+uxTjNJJ07sJBpCoIWWHfjRXfvWze0SH2+LvN0aEV
Jj/EdIf1plMsDM9w5ytOEfKAKE5o0aSda2D95lH8SP/SfI4C0vC7P+webc8s/ClJ
3NHwx0ARcqTW09R/eXezP66qyYSaSgv4wjC4VtNyEFJFTLY+6F+U6hexGEhiz4RS
0XHZOqVZgjN3TlIWYwXhUv5fRScgjE2lbqHTLApmP8GUDVoSPwFoPH/UKH0fv2Br
9e0JDjObDOINeu5/yooSrYEYSZZOw3dtUqKqniZWABhWrQjmwNKI4g0qpJGo6CDN
bzIfmUaaMslq4ktGE+Dy92YapIP7Pt8xV3/cC4RNykG/aC5hzAfiGRpjVy6+xHdr
IO1bim7+EM4JyQIK3otY032p907V7HHun6z7L83aCA+oLl1duLo59sY0xL+3YgFq
ic4jdV62s8carpdTrQKl1lrWCxBpajIE056xBlvUA+3JTkovZndgQl9/81pNIFdv
3DhXQ6lL8GSDpjG2tOzjtdtFf1LZ81EzIIDpsE9ALOjJVJ5AvxlQCNBpuZFAquq7
sjDCrzpM0en9EBQdEpkWT7andcHYSB90V3vmwYgVOUPvsFpFW2g2EPTbrg/SfQH2
tpF3a+Ap8g5ws3Kz+QJPenzbtUXIQQ/hOXcSmZeVAzBXryu6A8NurReErTcI7DuY
2GT2kxyPsv7YbDcYTWMPWX4HA9qETHg+JIZzDX1ADkFlrcFgiNL14EUZa/0T25S6
Jqmjfr8nIuYNrk9JwjhO9HbExIJhmraRwUn6HtOLEzWbDXxseUMTwBn3PaXVworM
yX0okEMW3UWLkQnNIbbXmtKkFL+d/XCWmVgQiti7l94uvBU3Kgm6Lre5dYZXCjm0
+Td7jNhfur92onjKy9wG6mkHdsBmSAstYUkbSfAThHX3qS7FhtPBSBmwY+CYfVRW
fC/oAYjReZj5hIfumE3t9J1vgTdCbrVFZgPftSqGuSYmS6EDdwKC021zoVg7TmXK
InEP1DoIxCUYQfFu+jsbm5CJR502HiR4nCaEJayABo7ux+LHiFHOxKtwMlSEsirK
4U88SFaByuMl+i4yqcCcbC3eBlRjy9i1jhLoaJK1+Y5Xcq8Al0WY+wrYIH38eZaI
B6xVFQNBJWuzYQRz8q44KQw+N6uTAPrWxmUxlthLFG9IJSTBujJiDzRwXBvRy6GW
RwJ6NabL0DnHjLY3VM1T82E4wAA5UtB7niN9euPJH2lVDXdWbbR4DKXrjsrKB+e5
PluE27WXAy2dNIXhtrr//7AU99PRXIu9/yFP/2GBhLpgGVqRo6840M/QzLMps98z
W8q9fy6QZdRCmXyL9EApTPcJuiegkw9D4eRSJSv5Sp03jHyPKGk1DAfQxZwACIln
4PEDwTMzWOs3R6qalAuo208XdWIZorMPFehl93hjrtiB/kFGbzmgQ80twCTjy2Mm
egs3zXZ8TbxY2YznARQk5D2xIV5tdoTaAwYHkxiNgPaxoXeykzL8yKzp1YEemHvN
KVTUug1jvkKrMMoJkq3RLg9EEOR7BNVP+aTfOEy900wPcIRGetKQCHg67z9MC6rZ
40kAI4fpHdicmBP1Daue0nJMmTdxLu3j3UcjeJM5GmpEBZy7oZLPMhfJDZ7PjKbt
LMuP/BuVO7SvAyy+wDAN+3/RxYfkd2XcteEQU0gcbB7LGqil8pECl3clF5Ov3gfB
JKIKKF6vscNvKz86emVs4GiBZ/lZlMODMlhCqeS2/tD1yWX+/TR/PC+mtki/DDZG
scjfcDYnTCedbFzTfKgMTIyXeZsHaf3BcAeC3bjFEusT2fP4zfoITJKKHafoCufg
rQKi/PnQRggP9u3Nst1IrVTM6LkIQ4VCAyvMwbHKuldgZ9Fs4FAS0OMwYbUzBd+S
Ka6qsffkw9GRYYCr+p4QPFx3QBdeOm5/Qzrq9JswxwZZUM+92XOwkirE15KVSU05
OazvjY1+OgfM8YVng9Do+XTpys6+P7l/jGtQMv31in438Z/w6N3X2+i2Vh+JaB5x
x1O35J6hw989yZLtI5ProegsGOkp8prfZSwmBDkmwYeQkEPjng/QIVQ5IuaZ+bMW
y4XxH/Ex+EUr+53Tzy/o/Z8m01LkAkYbe9io4vhnEedbjr6vntyWh9m0x9tgQ1m3
b+/VO1m6giFTINWx1hMyX4etiqQUZTGNomAR2sx+u+aEsNfSwW2EC74DcpEwpaW7
k/v/8er82Ony7W/s0GhP26CTegn/9AvPD/g7qOIY1uMrgQN4QmCsGnuO/oUWWI86
UyQHA+zL0ZhGqBD1jfHvwjW4mnhdw9esZEyPhFUNnXC3J6y725e0QWu/sQkVw7gJ
xSVJGf8CM9p/kC0mE/9oP9yA5lEHz/FHpMjU3b4bTEFXYL4c7JctA123Rt95wsxi
xkfKOdmnCg2ECghVxjgckollNo9GwEqPUXw0wpcYO4WYpVH/nkStBfHqSkEVsiT6
/027oTe+aMl6olgw2tfhqQA1ZbNRMqQJrFjLboznOofkjnGuTCRmAFVSKD6SeFUn
846pDQHMhLwSJlso/2N+kOLxcExbM+fQ6X3LvjhWNXpw+yUoWXgO/NdmXsoWjHQa
4Zmu6g0NvmiKpZJkWq3LgWC6NuMyJghZjvDi5H9TNAjTucAw7ncq9bEjjvh2ABDU
DWvOhZ7mtFav5lMI4e6WA5LNuqDFrEGUzvHSDeBSE6dGIhAv0wHOdqhMcqY5YWvF
9PQ89BdWY17/DRqW3fwKRpxwQ290SaDp4kueUNcnQAoRe35aUVEEk63Pycgd5o7h
kAcWYQdw0XrmOVdqRwkqAqTduzU0Nlcid4p7iEMMxtebMbuotcfv8zh+p/qLSkBP
u9wrWKuGZpOO29zIYyrrpqC8DnleRfGRY+2lOx6OFqTf3R/X0El5nysvnD6yMaTD
K338zTEQNjXf3jBcrhB1hln7DCyAx/X46nsHlcSp1d7DKKSg1hF1ClwZIQJrhpAR
GPirODMkcB3LHRZt7MBfS3qAi4FUdf09u9Qrhj6UemrFco0QCiWW2cxpj6PId7J2
rkFvAYc5P84xdPgNZgmm+tUKIr0nIYhJtyAO4EdG2YlgNi0eVmN0hbOV4gdevtUG
jk+fR4ALbGwQowqxAEUCPA8BLsT85dpMCtKqNLbYNEOL1nzti0I+xUzwkPE5FLeQ
1RZCbHEDeov5d/GJCI2CXrumF8zhgbp8ihQKMgIOclb0nQ1rhTBNOq6xFKFoRCgz
jC6WK9gdkrD6T0dP2dk0lPDFb5RfIJkBUNQE4uHyOGxNLxJWErnF1C6wS6VoOAT0
nD0k3x+To0VfdWWSkdhf1/VKLDUcrKtjSqeLG6GpjHLhw0N385TaPxvENoYt3HuN
0HT9BaqaBg4fjyJZOTj22fgy7BV10SI0a3HC8ekNDvEp2eb7J3vgl8BqdMma10rU
g4TmEwdVXc+1wrtTcVOcoUqL9mr4VsHc9+trMBonjzGVqLBBrQ3pispAozOtiNcE
+h9QoYg9kJwlCJSCijmkJMKqRV+STaEolDYcsCkudvXEmuItAx8BrSXp5A4q1dCW
hkM1dz58JoWyJU1p2hHuh4CfXJ8tc9SpBY03a67O118NGJ+mD2vYoN5oYu2ePOw7
Z+bmY83o+76h17PjfOUOyF2coPatO4GHm835A9Xm9y4fll13aYWD8oOXL/y2DVgk
7Yxo85EMftPmYjMdDyk18t5ryk4pdJCsHUNr4B2PztGiUafJNBUHEmKr1AM2//it
bYXEmQjJdN2pO2bi+7EnnKbzA3kZYDxBzLebNdYYfzTK5ruT3Bs4SyRWuoJfQTyT
vSNBWw7H8D30RvFJGdJYyrpLshvXsfodNUmNh8JsgYjqCqmRWN2/f7J+HyKr8nsB
PVntbTT52wAnXd82mCyz9QE8NE+WBxrekxQ9/DkDRyUU2KW9V15qnH+DWfpS9bji
NoovzoyIG3wvaQ7+vimxY9XWH9F8uVB+/uiE3e38QtKKtqyQF3E80js5d1bUoMVX
4Dc+7PTtoFO/PlP5xiyRQ0aXOrUKf4H51r1dYQYSTyxBBTYVG/B/XNGCOc/uyfQ6
A+A24jn+/vGQFS7nI9baPnljYIcZuo6lGApMU3VuGe5EmZc/UaGyn7ReUnXQComn
Hn3xbXhK9QoRyJ2NyhUYGbWWjZM3x2KW/Pky5U6G7SDazyV7KCwXATlwYR058YtT
p6XJzRqfgxvIIHm6RF1lqLPlQTINkx3gz6t8UdPUkd8kb81/T+2rKaYqbfKJk0C2
hBQQnT0VMWAYvb95p8qNWs9jcfPcl7zkkaOcStPTHymMrrPg31ZHUUVdVBRsKSx2
zXvc8EkpOhhm7/ClgmUmLRWoFGvxh9bX5N117XD8lHS8GF5sXtzIJru1nqe7wWrr
2cKdHDDI9FHmUJF/1zSoqN1lddnBrSgWlKIkhm9Mo7J+AhAf4/ll0ftQItOdVAOW
K5YY1Z1fLEoP6qK65VfUWEGGRCdprGXPRlgnIOr8tMpY6JLXNjnPXkq4FacItZzJ
9hbU17rt/aAQBOYpS1Vhnw+C55oQNIJKNff7QLd4p3skDf1KJ1cD0Ja0cPK50EQ8
UkUPyxLL601On5sUjuF0/wo5+qDIyoKjOuH2RxxvrTqolUvZpE6xTbAEEZFJR5p2
emg1DJ3wA22L1YMGGEKj1NR4avwWb4svauFLnw2MbXixKUFTqn2oODjBFlxtWVW+
aA0ik8BOztBs3j9NBGY7UlDYeXUiZav5J90Xhwjv5whC6GyNaM3o3uxmslD/+y0R
xxo5z2Wyzm9gKvFRGjIp7LxAm6B1C6luvkemsvWjiq9GbiJGrZqVHoQeOruibf4A
Z1+rBD7V1e+aMMe1/HMRJU3NASVZhJjOU+Z0g9kqtzGg7aYTMTPtdzpoCRbX7K6V
7lmHOWn8JVBwGQmCwQ93krZ5leTdwuDFTGmnEvIoAt4IAshHVRXIDXC71N7DzM/W
1R75jQGkcdT6HbJhBHJO2oAW8eAP3p1zPHygzaj1qi5DNCTXmlwDemMrpC3y6ew4
1b2P6r2t8sC1BmZPf9gLjFt0anv5Ey35B7FdokaJ3Ngk4VdCcz2j5fHUw+hS7vZ5
Qneu3/9100oHi5YKTe44e5n1lqtOKZarengMVx+GJHtoZcG8gznf9jMCzvpprkIy
HS4qsV4zBL2qf1tuce2cgdDEyyeAZgEPq2oqmyHSlQADbTRHojFLq8a7VmR3zq+l
agu9juNCIa0w616fVrGRCu9x830o/liFGKpq7HNioRAJv4wJkNb3xinOQI+UcnXM
45PRLfVl7A7ciYYaVoPxeor0LkAMt7U7d3GSW67Y/TLNCG57XBch5d/UOaoHhAEZ
sTufobT5OA/d1wGxnna6hYBRvGHnrgGvU1NG+GFb3rZUACBoi6DsrIXgsOq/rLWe
oFmdKvhHcyUwK2IkRb5N3AM6VAGCjM6snOef/XAdA5YFjQFK+XG3q12jhMncsIQV
b6i/7xU+zviQEDi02YXOhN2gdjYQpP7YpsMhQrXF4xj9xj51Evg68Xms/ZSnNR9I
pMOweU9t6v6k3v1Lk7MYgaOP7slS4OOUkbR9VvciligfCmzn4aNsFyYM1kYkcgVb
OHPrehqohwnl0fPDIcitginnnc7RiqekrVZHn6sYvGQdV0btK5wnZMLvOxgMtEYI
Egbtiv0P/1/Kq/ZqzOqdMoQSvLxw1k6iLz45ch320ns+VXfgMZn0CUn9Q/pxV3DG
RkIEawZXB/RoWkPos9G+Bq/zKBAwpstXuug95DvWEZ7VaQGssaZPMT1lzPbomUwM
JTEMj1yEwgaYKUMc3reHtaTbH0o9YFObbuSZ1mjL3vPjyFSS40w+2QQT/Zdm6Aln
M5AJek/25vcaNm2RX2u9iNpZvl9Q04ORKiv4XpG7WZcAIsfS/kOY557gx4S/qoVs
Hh6Tv/jnG9HP/NPuwZtkGFrLllgaHPM4melDxk4dCDawISmAODQNJztjxDqlXpuR
70DlpQApTlETsawVDem5at4pmNjfmq4VJqjFn4Lp1BHfz3A1QLqHMdWMDP9svc7P
XZuTgrOOjqZTO7boUsd6pfDEo6PiMrTxWqT49YCUugfyII3Lya5Tp0NbdvN6tDSs
GMobXjWX58s8cglYizwPwGcLTr8s2l7MSbmbieIrm4Vhjx5Fn0srJBiZGx0jbfyE
buw55z4xv8MdAbT+ICci9Bwkp+3ayDlIipVM7ZDrtDBiZskOYxIgOQAdH0Iu2qrc
67PhDyFu9tAD2j5Ez3wnJ+vEOi4Qqsph0RqvrO3U4/QJGgKgh/BQAMoihKxxXFcn
VwunRK1AZ8LgwgMM/TSKTqL0Zt7tF67RQVBpKzt1rOTr6GcN9BdieD0MA3AnXjuj
abDe58BU6kFQ6+T6oPtYerptigMdy7Tw+ry2O91YkTRfHwe6rplS02IzRM81IBUr
Sn5ohZYsBbqAzeSNw1dibCgQVzASVWYzWmvZQsmchk8nItIg9OyApov9WRMRbj4q
Gpkylq/7xF18FGr9j35QAqtpvzxQwNKhbI9JENQlNInwHD/tI/jNmIulvjPFDlTW
sR7G2LxenmtHcFJoNnX1RkZOpY24asyXS4m9IEfTNSyIURKhF06Vope68Dy1Blbs
b4uKwzFGQ/mhBlsKNkAZD/lALq9CN/k7VdcoYXOCJHQLaR1nZ3Dl6cwSejPlQTWV
JObfP/e5ZPZaYa4ngxoHvbsGqJ6nUC/7WFVfl5doVCLERLjEgwgB447+byCJDbba
mhAWEbzWY99g+8peMY9XFPkrpSWYNmGVPHcw3MEsZwtq/oRxpCTTAYnkEfu4etxo
qEV6s2vd/nGmUyi/LbZ628bP0pgRpbfWU7FnKDg3rIqwFKbWVZFFWR34vodm/D8J
4N2w0qKffnWsU7U82DyK2SdX6JxMxHwj673OqF8DiMZBPiKk8r8UyT0lCHdCXl49
0CSAKc3gWHikD0VE31GcNJAizgIwc6hbkABhXdmFbgNALj9O7EE7AwwT6buKxfer
wsKHeT1/hogaRVBMQdVG14Tb7/ch8HBGO9OZLfa5eCd4zAggpthwGMMF7RqhBYO6
29STBSqfz36/Srt4k3KuKHsT6Nhws4uNG/39cYPlGEOelyGQ+4AclEBT+yLevtvP
4p3L8et0MP321RANcd8Z5sZRdpyP4/wHGMMI7LoUutD9t5pIvMecKaaYUYH5foTA
B8uh9I4T9tqVZxsDsSoyJuvgsccpQbzUR6OxAVu6B/g+TzLFi7uliXLf2uYMjDjb
UiAXMgDXC41l7bAr+ADn4qZ32gSF8ZlXCx9ibl6VYM+kVV3jbNAKakYYzKg2SvOl
GsiXUMdySsDoKiWMHLgd5PsUjFd6r8lBNWmedU3h1KhVDRG3DmOMPUIEEC5C9GPw
TNGeY9xL42F19eb+AtxbumMM7bIhZh/gcbL+bqUuGZ0Vgs9qKzjzWUKu3e6Iidr0
VocTYnfSLv83VVxPW8+cKV1LJru9MneXIoXVCvhAM38tXfBXjjRKxfZReetxtV+Z
y1gpzLHIGXbQ4kQ4xYgRqkCvcWjkFflzBZYoVTdmzLG/7txlaJf5R3JNXb5GJ5Ox
lvimu45T8gZuX0nN1IidHqt7kK0taU2eQM6JnT7nOGasocvNvlTuBbqKOx8Aeu/Y
UDLYjyBy9OGrGVj9PZWX10eHB/IgZb3UGJLW6P/vCfhGRG93xhSn9SyJoYuHrMcC
n1k9HFF7RNX6Fd/SPffJXr8uS+qnAFW5XqQMx50OrQ1v1zt54dhss8+PrLMNpoNP
XLqphgp/omZbkUjrpwRprnpnMB9xZhAHQfc8RZ/2rYkqnZsvWnbYf1DjMdz5LLbg
sVfY2W4yk5apZjMakKoGxxGZp+R2M5+piU4OEbCKM/PdupljLX+j8JZJirCaQmSU
bAT8Dlmd76IKTOQCpAL3g0LkURki4s9B6WCyV3b3p3AzHrmhO+LWUxkWnsPmZ4PW
MEeLR3P5/dzSV+xiJLLP6xzCrYIvtOCFQKLVhdhfhNziUNGxQ6ZHOEKIM3A89Ex0
aGmlGx15biHIfFPf4JYEipSwoE1GJqoh1Jbx1Er5F50N2x3mVMEOmme++MZBbZys
+Lix+1FxBxA0CDYc0oQOKzBCjfrdwuS+BOqZMImH0i1QkyUBKU9i8QuPgEBU9NHF
spaMJM1I7uusp8ImZ9ObTAsyVzlq1EVufCbrELSimI+XUbtQt8Db0+ahx2VrGeNd
ydu882lzEP4KyL1rj0on2KdFn3k2NYC2pBmqxCK4y12UREvCSbp9mcYU05XdkuM1
b1k7dizfsvIDlePkNjbqCcDvzf4PC0S2+abcIXHxYS9m/XKK9M/2WdHApu2mE3k7
f6jYig0f0vkSmFqMp1nLcTyaMHNT1is423IyEaq3o7Qv+l0qZDW5IAny5WPCicfi
KDQSJf7N+7qJeXIyFEMNDL08UpPOXF20GW49AqXNpjjlLw6ehkgPmx8Y9jqdDx5U
e2jgaT6PUBmJ8PliKvVFepB1K2KjsIX5x4MNXZ31JQeY303heJqdZ0v6q3t1GoL/
DQCgqI2Z8yti+S9DEIfJ8dC9YPka4YzwT00yWAq4rr//xvhkY7MmQ5zJoAoFc0jq
e2xLJBwH4qw10CCndY+NgfKSIGJ2VLWcaOvSJcMZt9nJZcuBRavlqg+BgNgP25Ew
txtrFENpz9FaY76L4wzvgUyjsTkU4xb14EkrCxEKlle0RipPXkjV0dAzAebEtY2i
HT0c+QwijUjuWshJuIXiOAvezI76RKOVxX3JDTrQ6yjBO8SQkrckIqe7Dqm7QVem
z4i2LTMvPBYtjW4giv5hjF7P44Hzd6MSiVb2Vu0vPT7NUdBFsQBjT5tJ0prj+0/G
SbbVkmtB5st0coBB1U+h1v6et2/1KrQNPnJj6UYGjc7RbJISdMxL6rmx5JIs+gHc
FrPmoQs7HfPHrb62p0Y/jODHnqf7R3hYmwWsgKzOdTAdUeMDSyexHF32VQC995Rd
YQ2q0CaSrfcwfjIyGJkPCEknMpbfhjbJZdkvkcAxvUiC0WowfZXYt3oUPFtFdE4V
1sWt2ur60jsfxM96uAvKIEkx3/uHlco8SfPmQqQ0Pd8bA1hkEGcUuKpqwGDVd9XS
3sGbASpe08S4nOkhsSCuCs1iJR1XfRR1LotOrLAXtQcn4IQn40zLKJfnBH9QdDUg
fu27A/jatSeIgUlR+4BLNTpJrGe5VfB8U/7iro9Lbigua7JR741unMUN3qX4mD80
UN3Xv8Gi4UGRDK+bFrpn7UXD7fzot+XaxNpej8rO/bL9pGsIp7TNi+ub5jCHjRiI
Od0hWId8y1fhM+O3KbKlZNhPfnkFuDiidLJ0CTCrhOz0F6KLM2V3835OEnP8DWUw
dpUV7SPzaddYXEiUL6DIdVkX4+ExZ6GvDTEv0Z0la8xuBo8WzkQtpeyHy6dcPZt3
aLNKS0Fz6LJ3Pi9NdJUtFfpucUYLHN7ajFEbxC0oCxFYIhK2CYhUDG6ZSn3uCvj/
VdmoXqUoKLeCGiSYt7/TWKgQDa8Lcu+GdNoKO1/QC+A3Evj/HslFAY7VhLKbMyzD
BVzLylg/DkRJEvz5Mj68xWgQHPiaJNxtzeF2gu9dy5BykwAzlqo9yeNfE+nChaGk
8FGFowvVDnYzAd96JdSQYsAtdXb0lrJrI+UE2JV1xg+7s8M+/2cW4TaOOVR8XQ93
n6TtMl2Da/u1U6BI8hAo/vNqMPFi0S5O3X6J/nT2+gsgJLnJSiDMzhoZhP+scyZo
wExwukHtKgGQ3kT9cpXdAegdbyK5a4qtDpQtv9z7ONli8851XY2wVeKj6wa549Pr
HNOOKSLdZqjUka0cR22bsCAMaJ1AKk8iy7+CHIDIhawRkIm1KMTt43z9dWWcq8R7
UV243swi6jBQsQZhFloYkutl0wCYAz/17KuiNN0etMZ9epA6kn0UMWaRZg1LCq1u
szp/ISxL8M5kEKcwoIs7nasgMVsr4v6dQN3huWz1Q+h6BREk+Hn/4g6z0hR/hQqJ
phOL7Tx00idDq+Ld2qBdgjz53wLS3fX/nIq2W7Q5oHRUhF3aFrgyg9ZJxkeEynsR
7vIu/drroH0p5O6y1jukKbDNyXKMU/IPYCglzblIPscK+7uQoNKgNygxYBEabjko
3+wjqEOA9FGzg3cjxxcnIkhIam76BTkEOoUvl/avrOU8hWQRzXGqryUx8TsmhfSu
wfPaDoJmcBeoVEk/RjE1wUoudL+MHmohdTJNXBf3yRdt43wYW2z2tysmlTxhVp9K
SQ2ZhmCDffvd1SIm3K2pu4RE8ja4jzlJZ7gpRIXb3MhAGI2Xihd1OMVbBQeSdc+w
tyy3IR5qwCCnsVMUj+JFVM21apsqDx2I/zsqxMP4IAcnEGLhDKXPbcOMpb8gkvKU
qLOardekFFLYb/JDt5cilh3FRztMVi6xXh/fqa7qWSJz96YjXmhG6j9Vd/cssWPx
LUkyb09eYyBNHuclVZ0Kon8cN62fdAwUzweQGGWjTu/kTyKRBnfA+6KRpCS2R+JH
5KUEWqz9/x3oV351f3bbmK9gBN5pN6WBMy7gH3SFW1VoSPa+5JcCJRLZaiofKYs+
bkyItQoFUvZPDLu1vd6cJV78h0HW2RNZgoXpnAaVrU0BeMy2zr/PNRIUCKSGHcZK
Cp5E9JXNOoveXt6519EqejLR1DDX3DrMl1lo/1qbrcvk1aksnsa7ae+yky17mvkL
ClaaaP7JBFRm8rwBfEaxZa+aiSsCHAxe6f+4nRbJCQ1dK2SRrR45UWN5QLgAOp4W
opG2mXVHEc6u6gDC0I9uyTHw87bbB90i1In6EJllQAXn1siiWYEEhWPpRQ201z/8
F5g+gaU8rxZ+5BpKlWbAodfACGOupgCg+TmMr+3ZStnzx2qsRcEy30DJFDYIkzT0
SwScVXAK1Tj+90+l6Y/t/I9t6gYG+G67nyo8GARglczVOVFmpTBZ6mMvq3hlZeuy
Kg/1By8xRz+ADDbpsKWX6SclY3uzVMSchvna7tqARIcBTkgYJxnSLE0Hqhicrhg0
EDld1Y/y0knCeoREQ0g8f4VZ8iXa6anormHeZpn7p/q8augU1R0AOfJ+Xn6muick
SsUEHy3iAqtRchISYoiSfBJaWyNiuwVVR6JVB+Yb6dtLW1GBWraNi8HDaxHSiMa1
AsKHcz8SquBOmhTJ3RweCz4049Rl/KEo9w8NRgfIdYGgpGrQjgTwVesQIu5ZrGGm
O98ClcxbO4HaarKphhxE6IIvTSn/t3Grdj8aoS06I4elnJMHmPNJCxlIw14e8bgi
XyySsNAbN5oHeAg2akeTkF4Hltv8AABK7EaW71VhvHp0v+azl7U16piTzLbIhSfi
BS+fap0lETgBiKKeAN9BNdd8fkNUgHpmUzeL5aMW002dDP56h2msQALYlMQXmgmm
vsFllaCxIYiBtWxOe6raGFvI5TPsh4EY1N4wW6BNUSXtj7AbwSczYVCHkpMxjnVx
W3FSAEBlLKBLi2sL77uEpKsXA+dfRIRixLC+S4p43srw0d4KnuAfnr+IxOPu9NkY
I2hm8cINkVovUL8CnA3HR3Bl4BbptuUqj9CMTZt+dT2/TfRfopyQOn7pGfm0A1yR
H+xxoBFUCnVekODXC9920sueuWKz3kCns87KnW0OUgro4BbTVk+aswci/46GwZA2
K/BbHCSYmG8yKwx6lL6V5CE2+hzSFbFqdTNDGQYVb1u4jHuvg/LTSe+YtQKhx5gG
+Iv/oWEx5WHuRxWf+EDixmviOKzL+r8ZtdDOQi0LbANd+zDCR5jv/gTZjf9mRNbA
kbsJfdUMkjmQD5YvntUx3IXt1LVhOmJWdoEGIbG4RgLERtl3WOoNw5C+jAw67f0a
tXY89j6gtKM6wPv8oNPRrQGutkUO1eElznkl7zDgBtKvXH9GCLyjmDr/HHuzcZXB
cCWIzru+t+AEzPisx+u5YPSnzfDMaBxki+X18iNoPscvN2rDR3kB5Z7bzNsAImc2
ZJ9sKJAUh/i7dSG7va9uNtVZyVGnd4mxLNNUU3JhihfbJkQzzjIT8sFI/jzr+Vzl
wA6q4/gwhh1XfyClVim+aTZttwtu6blOvs3xkySNkDmjYuM9oVDglH0ngNA7OR9x
k7Kil3AUzuFeZGwy/pRQ/Tf6rYKbttcSCRzmxGoueqnoDJm8/o+ecM9H75qQ3ekO
MkmnXDM9cEkPqqaynuVpDXgZgxsA1cLToa5di7+lswe+cBowaor1He4xaL0thebE
cz89IwGrMo3rRQgKD8eGPA/13EGzIssIDae2NTlvPzqLYUYHVf1atHlro7RwMnjE
vvkQJ26nzp+oA3P5dyCjiDn/i9QEdoOhnhl2L4L0W/k4st7mM8MS+0G5CP4BH06V
2MsroWWjZSqZscIIGByXRVccP33WQTvfESA+o5TUt3uyIsFeLYAEwIX+XjL92Onh
FG5jgWRZXKqWiYVWcH5e9cdBrVz9EHw/n/X768ixs9OVrpGhhorAITWG3a39FFEv
xC+AzmNJrJ9kFB0+iorrn7UZa89lb3ugCGgGZaL4gGm4qcwrpIV++BM32EmfPp7d
0kjGO46mtOB2lyaj9VvrUcHwUtZp1+QMBcNScPR1r9BbB3+IoErXfC9ahl97WNCQ
EzPju5SGuqsR+VvrROFox3Chfb0IkBXsvQw0ogs217WGLUuRsTWDTZQGfAC04BG3
oLk3/cErzquXLZFOccdS79phQ+HcUUBt0TmW6L64zRMwuSUOn6EOw+5F65IpLh5X
WTCglPbEcQuO+NZxePvc0oOPD218ufmmO9Y8Yix63DzVNef2kHKAHRZkL6M9abZG
YzMzVZXA8OcYTdFqbVOo/pf+HWApJDIY+UdM7G6PVENepCJRguuwq43Xkx8iYMtS
swrgti5tG8Y8WzbVgQjXLb/rEDnYxABmOgA3UBpxhY+KXUT3PZWnhMfJ4VFT5Mvk
8j3jYaAkw16pBqV3v1C28xEO+aP7FiUiwI7sOaklXpiTLtSsN9rtrwg+hjB5FleV
rwrMPiKiy8P/GjPDeAxHoG4dUCzVPKjRBdgV5QMJJDMVgZrBDMdws+eGRyI5uKAs
+C7BnzhFiaf+z9/3AHp7hp8fRIrLk3sq+3O5n5R1uV/c8FuHiZujAmQBgV5DEjPC
spcpvJyW4AwGMkZuG5sXiiXiy7lqJjBK5MZb6T6GPG60nHHT+doxNhBXeXnIx+1Y
msespJjoB0xTjZ9z5S73POB/uGMrFbpv9PVmdGCvqABNYbnlGHVrLpgwyvUJYkFT
lnhejGPgfrZ3fQWavgClgK1SM8+JhHdxkFwVVxJDlD9mzinCPa2Dg5hB+CXPILxe
i5tfsCdiYWcS/4fxYFGOxJcXMN2R9dX8pS0t82napwWOJsM8a5zPAfWDi+QazZZQ
/PTymjLcltzueLye/ft3bdsq2vZ+2b8GWYVqjdeQsYcox4uIKBtZCp6z02lxMUN+
gZD9cLwvKRdVqxxfzZ5P/lgvtERTTLwHPbDczkmEauuZ9sqbpAnPAJsZsvoeqfH+
Y1UlbgSOYVtKa9kHaKi3pMPBBhBm7UU+wALXdv4IRd7UQ7vYfHpmzoWID6bU0sns
MQuI6RgwzK8ZBsBdhiPHwG55S5h/aB81NNCmQS5lD7uB/r61aj4qBgO8yrY3dxT2
07gXSISiUFhcbJyOkwIfv3/mq2G6mpuKAhvJHMCNH9kbXpf7dIvKGD0/UBF+G7Oq
0MAaCmLaS4RQqnwGk77PL1Xyujm1a1Vtel9Bdd5Ox/ORqIZPqxIEXJNJPQP6zTn/
9eycsQfajhnA5da4xhdUctY8T3l852kRI/ZqdLff/d9oNFvJvPUlbp+c/1tqkpk0
3SuUTK+M8emDpNt03aUD42JTs3jnBOA3/4LhFsirdNCXUGfhXBTHSWYTUDG5OT86
6ueWN7RnlfWh4xC13DniwAOZOZzLgbyL8dC14auJglubStNbpkMg0P21IzC7JI3C
rSQMf9F+WrJKyh7Najz8eqLJFDy+468peWLAAgzZMrYRItD9AsgMDTYpvT9xUnVX
ElluEzIXBySTzhcwRdfwEX3Xb03ZZp81Dbfk5SocN3w4UCktoRmyNp5V5nre9jtC
E82mGnpaDCfvitNvCR0DGsLmP0B35ThIq6U2ih+PynPfmMr1mmyfJWRKxCjdTrdl
HJeuocXXhhXCTzmx2YiL0/SG/YYuyraEOVxxT6PV1TIYj3FzI1lodXNrl8HawTsN
17HHIFLzUu53V9OzuIB5mlZd2QRkp1LVLh/OM299q8LOwRzYN9AuxoDO6dYsIqu6
UdEk3fP62bskBM//LckMHJB69ZMEtkoFYB3bhvTqG+HEG8HJkCU7Y8Dys4Yfo9Gi
LCDEdD5f8bBVJgEEy2L+hLK3emvAh1EULhHlFeSQKUZtxKhOpzfveRwx2hEBOTKS
2u6dMnwFUKlptUjH2GAkByDHW1G5dFHPZhF81HEnPesbtnD2F1ReZIyNc01qXZGq
Nw4NMo0VJEa3yMKELdk4fQHvmZG/R02XY6wZ/ebMOha0BqXcfPw8LKpz2PJe33SB
ANAeMEgZJ6irRfKLnN62IdsUprj1TjPiOH9avfhj+yN+bt0GpEEcHaLTIMjpfD8C
kiAa3XPLk0gxoouVKXG2zKBLQqRL4T8jPL4hBlpo/6yyHwAa1ss/JBPnVlq9m9GV
n1qtadqyQS57y7QVCzbOgxM3yCh2p6V+hdVWfyKs1AzGZ8PXXaKbdZg5f4qIUj+O
Q+hFkVtk7nRVSialLxDg6p/7xKkJxLS7GsGCDyeGK0syneYTAW+X6dvuOLPTNcJg
mntCjgCSMFaS4hw/DPiZRKdAo04SxyjrOI4UkAcBsMTFooiHY986a9UBADIFQY6Y
4qF/k5ufO1UHLYWUdm5QoZIkf9M344i57UIBZ1yH6FrkQs4sRYifFjzVETkefuj6
8Mj580Tcn4yH8O/SnT5kh+//86oNd1hV+UjfooXh/s1yv+Y0vjHOceqqxjXisys2
ed24wV7hwSG2BNrPRjnTkySme1yW6o5fbPD6NAbC/vJlSmTra6/50WuYKX0vxBJL
9ZctssGUyQbkWVrlWXtO6OHEd/mL7vc1DoYM1LrdmpIvSKD1iIfbHF60BlpOGZ6V
BRBAFdED2fZG4t9544+zsORUY9D97JyIi5F676NNnpw2KWsMLZasrtWXbvD/20qZ
+g7WPLzwD6ff5p9X7jBnoKGmb4DRUce7Gjy8SoWdYHD5L/esDC9uODxBUSjyTymG
X7pqOeKNq4kMZd4cMh1k0tpyDEVxpUfHxOm0MVxFM3wJ6OevhKfPGZYzcK/HxqqN
9+GP2g/ObzukaEHIlHALxlXBppjPXZSHGJ7BT8Nq0fddspboXO4sllUBEBRxqNb3
NKwLUpK+YsD2OR4YYGK+mub/gCWbF3oWYchoaRWBKeg9tPEmPcYxVsB9naneieUH
+bly/s8iogQ1qNMO8K01Dqoyi9gcefk6h3535sK4yEXjFYGkX6sdOIfbEavjT092
39xo9RuBskv3lGsb9YXVd1YJBCTOq4WQyjydny2a+kLXFLsTvTjKmUByMfwGFcSN
zSjJKxz+rFSKvEnlvGvlu8cCw2uM1lDy3Okl/mFUvuYdCdUTnGb0ssrrwCF2n3kv
XHNVVAwkmZcY949qGWfxgzpiLqFhxiPJcSjerrpdsSiFTtxM1cQ8SBo9o6R7wZou
PnIBATWwQ9N8MHC8ZXxhyS8IjvmzVOPZt6Yd6V8Ztquu4QiJOqXIZJSJnpZWWutw
zW32x+nfrxfG68xg8WuOB765m30BKZY3Hz+iQvY8fU/CFPqgXspmdhFj5nlajxA9
yluSX9E5DGSaqXiA/P4gdhKOludb0oXfjGVoUkrvicpdOstF5xJU+u1l1cgCmmQp
LMxBadGOYgLMhly1bCRffVMPxP9/OopbCDCei7Tep4VbWk4+kDLKGbncMkAZGQsb
Wb3GNQBw0O7fhXdatCSaCA3KujHwKkuhp5vvfQj7H7cQwUZeb5+zK2Uva+xtBWXS
XIf+wG2OA/PCCmQlr8NtUPgXHU8d6hy2BUbvgwcOh0z+10tcL7aFlNH+tAbuRl4T
MwQbxHFZ8583SGtXRlJ/Xz867dbCp9xw8hE05/wORFIncVHrImSAFAY3ocMM3/7h
9slsHQCjj7ny/HUcTHuLMnGigqrQiib3o0a9J+z/ydA5DOLINULAgud0KQLG9F8S
u3P5cuXoAlZTcVbAVLgujLHAN8JK1jw2vnus6Xby4yUgScVOMG745G6Bcy1NcSnz
AzJGZGDv4TPWoFr4TUNC5Z3ssuTsLk6ysVQlw0LpuVamjL5xyUsDeZoia9+qLUMz
3YtELiSbgWaMiFFgwpG+Q48/vhDfR3eSuoa9zvjcorYl+NQd8ibMoPFpGL1iWEWE
IuqusvsTyeJRIFBJeCVCrYQgcqRjOfFwr9eKBW03IuKycBG/eC0bL2PqJ4pgmKVm
DJyjauiI0aMOhkwoD2E2kABWv+7KzkxH2hn6ux2Bg1p3YL29Il0YJZErBEuoz1GA
DIG0tb9/8YyKox0Fqtf17iNkKRzLGx/ZNqvg2/NuhzrYKtZ0xvpwqgySPW2nTllE
nwsS/9qNip/j2akSMGdzDutScpldL2zs/brbYKZ6yDSVOKRDPUv6tMgoIryyXNtL
XX8m3cuWpKycZGjIsGzmU3I8SGs+/AHsQkYgdKLEovjOGZmzDY3v0cZV//pSnZhb
ghrleSrd2RgALpe+ZxlxZ53dPSEWMszLkQ6OZH3m+8Q+qaup0JRq6KeCdtSz/8Ej
jT5IV6+FbwjQdBPj0+giMrwkWqEdfjOAa2vnUMMaUmaan2kFAq8yTFQMxU1fQDMg
9V41KUdAVnGyKytCOy4gBqYOw35sXy7/YAD1SzfILTS6qJSQRppKegNClZ+QjU2Q
Gi3c/KZMOR4pKgoT2drTlky9NbmIF9/6fa/LS5Orf0A1380EeVSJbgOhD2VMe4nl
yc/HvtvQxwTo2Yk3hp0AseXU3X2Dxj6m2FtpYKt/XR4nTtEDc65H85+dOQGpU9By
En+a0hMChYM1ePMEJqJexyzmdLeL9mN2V0WTH+IwaibygX7oq1nxYHkx3F9kBbF1
Fhea40sywq2zliLW6qUXR/2/vCYj1LrFkywuGjXO5Oc5x+lDnWsNfv3O42V5b51E
ayUZ1i9uVXRkL112NCf0nKddkxdXp4hE7spjL6tgq3odTs6WbxpKNzblo8sBK3zL
7y9lS6SmKvQAO5mQKBgOhfkjRzT4mCK9j4N9mXcwsJQi4+jM7VsGWTawSsZuTM6a
SoOcVz2mGZu9SK2KAx+G8FvmD2q2j0IekTNupQW8QhlGRMpsGUZtVMXpWW33Wn6z
wcYMIjcpLFsCQYlxXT5nGh+Rsax2SZFJ06iU9yAx/Y+LNA2Ow1v+kxOdmoxgW/ig
jNv7SOpNK8QbaeBJ3lDarGBTcIXQWjBmqwFOBnftLO0nzMQdOTDjSa+jtcDoAZwa
E+xbmvvIR06te7jkbJwKbiWzi/eVpPmErSoRrAwUxklEwjMLcJdT5+4/DwtBAwvr
PzYxoj0hMOf7G1CmTX308+Ebr0ylwfdqavdbN/7psv5NEawjLMpqmy86EN05SfcK
s6T3V6PBbLtU/HtIUGUAoebb4D6M1j/5WuzOXzjrVhKG3Zkhl9yvYP3d7AY4DT9U
AeQz+YYotK2/M8hbQBQwXDASeyRRi0ZK0As7Sw7XAmW3WWYrI0klU8CKPB+2ywbK
yu3aRfOhigmZrLlFr2y0SOj7XKaBFgsIsnfwDzEu7O4TVXTBHH/E0ALoKq4m4aNK
QTd5Gozo1Wwx51uzIx712x21Z3ZwTC2SQsHSEIdxtqjygJB0N4z9X3ARwRUat7zq
FMYd/pPJ1Q0OdAngvj33B1TiTIEb0qWfNusQYJfy9ecHsb/dVY4hN6h+QJOTp/1F
GbhmjYRm2zB3Kr1kpET7LLGMnxeSnfBk2Hk4IrC3SbNzG75HSzqiI2QGiqsXcO/A
rsuPxn7NoSeOH8cgARpHBxOYEwDKfclK6DxoftoKajXKDUgxd0TKMvW4LymOffTT
L+zm9RrwM0xTfP1Q3nR6SaII5U1hsiOOkALthFq38iUeMxd0GpgMAxE4/1a9sk+e
orqGoI0ohQy8dPAYQnHxYRSxahQBpScMy2kW5iVMM/bdlXZkyCoimcR224ehDTKa
tdUHEt/KxZPFhHi8dHlUEZcRsKRcFggutVwF9IlzEJ/+SyStGZ6mSe+NJEB6GHLi
KRR2Oum4wcjnzSEd/FlvoE5MOgSDAzQfjNF6CqHlNoRNLAvRkUk8MI4En3YKnfiw
IYMZVHn9fsypMubk2JOqiXSBGUVDbxHwV46kldgNfDQG7jmeNFIA2/771xIPO8uG
amRTzjClNgT9lJgjGHMqm8daREUrYBdPdHtIX35xCSnlLCZhhCFYUgGO/qbSM3fX
VwrD6jBbtOJvADP2aI5mlGnpfcQ3IrNjhdl7Zpu2RO3FJE3ecf4GO4SN73i1D0Z6
kq3CMV5DofMHXE5FW7ib1dnFHmKICDhNYXj3ecsH8y+ySl/iuiE3UzTYaZ7CTEfn
ct+cO+gONlguD2TlBdrGg8wmb6U2nxs9T/C0515BjfT2mo0o3NsncQWgKs8+PwhS
9OO0QX4C68KX8V9Jaw27/P4scNboSuBvZNWVQ8gFFJ1TwhzFq+t2Jo9cDjAZeBsX
DTqPaauRETJJzJ96G7recmrZWN42OwmJ9fhKMG0TDwl3MqyfOy7SAA3cP23ph4Nl
ArzasU+TBEkGp4sfpcpxpyBwVAyl20eNamuv/bi41oDwA4WX6/FEGGbKZtCX1gF3
Ye3MQWHBrKOMdjfgWkQZiCcZv8r2S+Zk5g0W38+O809n6DGFOh7Zv6c37tUlnWn2
nxNxv2rS83a+QitiyCMp7hnyffBpGChaNqt0ZfE1WIXdPMt6vmo4T5L9O9aGpU++
LZx3twctrG/dJm4e5UG6ZQDZ0m8LwU5D1+4hsXHSB3Yld80k6o61Wl3qnMMpd6Iz
2P2TUPU4+/YAg54X94vd+k2E7709c6NioxlYcPYk4sRIMYb8PyJ1nWwj5pqaHCz0
aDWow2b+YCVfWJuPKJL0xSyf/nDBnayIpwduwSoXB3kK8uHvB+6i0BGb2v+yhl+I
dbJ0N9ahtKvmHnUaTPytAAE7d6kl0zDXRM+xrB64EtnE03cBh25kSiH0PhB+uax9
0UhXNqSeiPEW4me4SS98ravirXu2TnA75ZAkFLdsRPmtrp9mo27JtCKyQSplqmuI
vYgJCQvmgQTAqJeuxdvjdHK7cYxL2XXZf4ndX1tR8egYEN0RlABuCY/1jHYU443D
LNHREjfWlS9+1CwjDmhK9Zu+A1K2WaSpeph/JSiFRHKpN/4ynr95qZ7pc99tNX4d
QtQ9BIlPjsHHSSXzARSu/nK/82oxn0jnEGWfN1iZWyWBYfhXjW+MDEZ0JriloxyZ
tWMkGXxRJq/sLvNdNA6KVGXfUZN53XeyjqzSK6cZb7fChvlkmDjQgZa5UiKhkksz
0/QjZQmyauer0/itNX64FpvpiQJ3tL7BUdHi7Ijl/mJcpwW7yhsSyIjUiiQAh428
5r0oFqB2DMgjVupejoHlOAVfSGjAPXGl1GrFAcEZn1Z3/FprqHngZYfgYe3BUIZB
NHT4V3qX39GQKYhIo9M8mOY+x4nlwcn15GC3daLPTWNaPew0xy8NepeGLzbVrcNd
GPLZG7z9aCCOCmzth6Qpzr9rqXeX4b/wOyu1kC1IqaKabgQQCHG9rYsql/bkB+Jr
aw9T2s9aqcjDZTytG8YUamUmEYpdgEcnVIfH3U5BnZENHLO+CihthFouxyartmlc
PgI+YsQeB53AzR+6qxIjdx6kZmd/mvCYgzt5RF27IwIn1jIXpb7lMxoDJwrzZEXe
AjH7ITRXgmHq6T8suBaVvmNQTzhc0JNJGNoSWMqzN/z8URW3nWLpsFfWNEkMgs19
og1voDJafmPbGiF+7+qUr1x+INV3w2qYp0LeWT1cRKXr2x1Syfv0iF9ya/vCe2Cc
AQpNxVN0dCfPUNfQ2RHvYtxCr4CLmDG+UPhLwaD54CSUjTK8n0Yq8knxZLkI66a3
giihSnYO0MiVjBNoie1qe4uGZdOjKjPArR+I/dW5NQT0Cae4g4SCU90ewt38VdDR
3rjlkgrlUFFU7VCA3xENFVNpCGtdEDURxoXtCoRj92ShpCqJLAU7nUSB1BcQ/hFl
B63K4HwNKVUTt8AhG3ln5FVE8DqA4JIssuSJ4t3nBsS2cAfa192vzC//iXlwzIus
+bFVM/sTp4ZAuriZnZm6bX1vSlD0YqZdBb1IF7SzepXDhLt3T11XKhkuOA7LU+Yu
zB5INDb/wJaYoflK1JucjEjZxY2V1A2nzhNgLzcdm5Nq0jPvuaVdCHu6Cwtc77+k
c1NbOFb0b1H97Hyo8fZHD5Pr+YLkeI1PhC44mCtuuYmjaBGyqjH7P66NMWcSPYjJ
hfED7libk3CAXvCC+uqD2+CcrCF3ML5VwoJIXQqTV9kH6iZCxjJ7mMNyLNvifqTJ
2zaXpS4hV63Dujo1l6GJbNkjDSiX1pmNE7ZpcHT9FSCV2ifOtIcs2H6bOClVlqs6
+w7uoRaSC9U548ozMi6EtI/a5GATf+twfhSWx4j9nRK9pjG3dHjFtBrOJI9eW3U6
Wk5nMEslRa7Xj/hkp5Lz6pa75ICqLUwoCtfDxrvmPrW5NfHuVigKd5lJmA0Mc0BM
v6lOLN3t//mE3veEUn7kSGgtfSuifGzW40pupWwCS+QIrUHXQRlF/KAJgODVlS1Q
tuJW3mm497iHjyUhnR6ktpU4iNPcB0jnQCl5pj/GJ+kMV173rGtZPBSGmmnwirRN
R/uaUWTWPyqpIQC35vBa9rWZAMejv94NwYn0d5oJG73s0s0a+ii8i7bYwJReXUhG
3i+fheD7rAi/ERIYwBmOHJJSFK0LbYoNjHlptQlEK7WxclnY5Lp50zG0d5vPvAOk
+efumv+n8HLsLLlIPEp2XmNEJbe1FMATm3b26Om66gRRAWPzQuevtEmpNzEdEN+b
Ls/kzGIelSkS2bm1Pvh9mv9O+Rpu9GnTzDlTik2RqL9Hxgh6CZQEkyONpklEETzl
GmjWKcsTxzr0/5VgZN1DGkm8b27HLPIeubStGuo89DOGT9Tp21HtL9S6MuA/apf9
TvyjftZS7RxHwPE1DpFAWmsymloj9w8jJDDYDxZQ/250rDtzDEyMg/L5LKt4pikm
kfmoINqb3AnwampG4z9CI72UlWl+x7rjCSCNi0Gq1YqBJZ3DSus7eOD251vjgyuf
UGbvb/aPQsWdPkvwqLWzhSgqDT9mzEWL+cAKPCj7mt1XnzXrdafQ9uIaFUvo7617
zTF68f2XCzxZZBtvz4v2vmq8umeh4dXF8VfKKLNPQXOkuCfQTosLapQHRczPPSg6
BsM7E2RJ8sU1wLV3n+qZi+tQOfTtxK6DErgrAic33D/57mi594VMl+GSCkyXiw5N
c8B0EIorl/ssESIklaBIc4q9108YQC5IYkQCNQof0Cdl+6yuJrHBtfAr+Zk2Chx+
GKdy1+Uqid7uVXFsIiH6RFtFxzebce2TFauWiMJB9uwsepN3cGEFHRxc4S0pGJNa
jd/PiTBI5+BnGXbdIRYQY8GbzJmwle1WtukYSiC5di/DtNDLb9Nh3fxdSUU91VKo
0ntqco4Gk35orBpTX5+pOxIixZ+5afoKBCr506m6mfGolmZ3rdfYj7uvQZrr3gGW
ohc+lo2Gjb3Z/+PFCr3PFPniThCALFf5Edb5/fnqwOEdBgnHTi30SulGt9egZYcr
286cgm6sAcYSJ5f3jME9rakGWU/PWN+hy29HIoe4AWqU6WjIZ1zhBx0KqVwiGCw9
PIesbu6t6yBb8U8chwyxxxW0aCeWnYoqIRCUWcZrWmy+0yZMIU1Cs7qNLYDV2bO9
PkFAeL8W/B9medp7yFKKRUpu5zA4xnz/m1ovDhf1q7q63BWHRFYfhj+eku7KN7di
69lvnTxssMeOWcGKRiJd0Fe3BZFNNrfXA+aGrMK7+GbSwrgvsUXJrjgcdbCZynob
wIb/120/TFmu4J91TyNS4dTXDdAvVjFDbtfbr/dGODIf0D3rM68T5UnnzCNJw0kp
eLeYZp8RfAKwPb17pM9OEHWuD2zPgCqOI3lPiLoVKM6KTfn1GBA0gN4IzGZvVrdu
k9wLorHBCah37kvXzRnQ0JFmCC23GfUk3FcX4HSMUKwsoz6QdPFf7O7uHEXSn4xP
K0VdQf8/mJcqrYpTSb8IviTSXi89pDU8nmqp0LOyHRnbRcy4liuFAfBOz/OBlcWe
vzazqRoJK/gzRuZVAAxnT54sYNAXGuFmVmG8M55rQ2QBRYjlh46NulssC3PIwxEX
2BkXq1HgPczVF7BcyR8czPvrIVkeSzx7OvaRB7T833iStus0byY58CQrSIx91Bpi
vTlxkOg9uu5G2VmCWTb98RpcwwJwzfyyUxa4PvvDdD8VxrTdirPL8RkCOeE6ahs/
tAIsLoG1m85nuBBmbr4m+6EEuCB0AZoOm1VLVAq7lXaRYtr6qB2va06Jaqsq7NTp
eztFv5sAGbkYwlnGFIkRWMBxRk65BWnvgw/5Di0DN0Ii645GBh7huL8ZJrae6j8G
CSeaUAzWT9+NT1H5jR7hwuQFYmPU8j6SYQ02Suc3ITIt+1ZE1cFLC/wRgaK3X7CO
EBu6RAABwVCYnkB38caNeqA6pPTUuexTbcSTKhs3jC5RiHu9XWFH9dMQFG54cq1X
B25/Dqj+NXvRUXDniLRkzBDY9lxFBbrrhJLB7KC7YPNTkWYMK16acQYnQPgurkh5
uMyz/ob19amsyED/vTI4PTowrNsVTcvbif9xVZiapXzIXVqNkedyZFebOUzb/jXy
PLGxjuOBx0FH+8c556qV70QW3aUerQp0KKRtWcwTZrZg2H/Amkg7RnSzGQYaR2X6
AgzAFNXL7ycrHgqUbKSkQf9Vns+ew07/vo2YXFkZ7pYWEenrBOrPFJpkVZgZyd4/
BkNI72SG94Eku3EbSEt3ErLfIDcpxdKROdKZDemZDfZbIa/orFTc+Uw9kAEbk9Ke
x02cCG9oxhjC+eWTxF2nIOpv3KPhiAnrC8xkmLztASm9ZOojgvC8drkjAertnszB
jBesMOVoNn7W2zVjItYsGlcdL9DzLdRK8xkK2LHjh0nZUH4ZLzhOKMLNYY4QD7cf
Shx8XV0VyStUDCx4/WCwalrpgN4vbSBAtwT7f5Zmk3uPLFjzeb0QhBFbK1/wCQ7V
pg3pjM+lBMBeCQvOA8chpDi9u7X3XmYBmD2PCXV+hpKTjtxB9f7Fac3NuOOYylMa
V/aiczy8dNd8drOjRF0196W5amiN7pfeXCwkTUD+wayLWoKtd/XUvC9u6ESq4uno
jmrlz1vrOH0FPlhB+VNMT/xFw749AgtYDgw1gqwL7rUob7n3Lw3ZuvYDCZ4yOHen
HWjaS+oUzN+eWeeFdFbZ05HpYZab0U7ipjQQZ+LORUAxFx9jFzLUKHxHAeUgXhCT
XOmA+4b1Wc45uVau008QendKKt2RK+T8KkzwTPHwq/BRNnb6ia/ux7LHQO6kwAfR
L09+vqNHkQOosuMoieyUo2hk/B6YGRN5js/biVUgWzk75NOCj0nJgdrtvUFxbnd2
M64xQdoZvBBasV1xgyPYgNzYPjHtKNJTNHxQXij/F2xzlY2sJGfXaiKFEC7XJhn9
M3vBH9axMLrCnmEi6eYrVLvOsxacGQTC5DyssAoYKOwCUllwO7bku8KjRaTfv99T
DQcSk37r+qL9TszUKDwW0bNum4IALKewaei+5JXuWYZU9AqV2VwgAsarO179Gh9m
GsIj1PW88rv454bwbIo41kFtyrgyL5bndeSzrvbFQ187MH7oErB3/MfV3jE5Bu3e
irKjZupcVnRMLbyX8DFhjB9q8n0BoUhsjUrMYIsZyJaH2t1mjaXg9zo8rwS40etH
nnDrF0YDIRTFdijJ++WNcmd8Ry1ebDhzsik7Q8vmJ+FzfRJ+8OwjERMkHQriu6lK
e3WSgxRn2zfuInX3NSTgrIUDvNBVGq/z+YPIaz/AKbSOCEk3Rw4SfpRbaGSUjVpS
Waz+zO54uHc38ncs9iyVueNs3zD8mgXqEaI7eC5M0BQo6IkeWX9ekwfQaYULZ78b
qtvLsuMGHdSIXkQB/y6RhZoYaOzvHvF2fndPgNQgMyLg2wSdxyyuE+9ZqHEN7qeg
Ymt7pV1hnpfvx5wrdiSJ5GqIrq/sN1evjfRPk55hUxOU+P6a8HtswnCB0PveM1Nj
/O/zRW4QmuElqyPIgsNhXvVDNBUOMHiufiPcibOmAg/N5JqNAvThT5lZiFDEPPAI
EsRxElSmapv2WN7MCGn2f8fyt9fZ6a/Zwvcb5590lvpkIJmZ7ul8j1fKMso37uSd
eTQOYbf2O9A1Z1j4LVaM3a7MiptTIq+aMX7HyQv2bxY0AgwExNph0NaFHMNtIEfL
fdmSf/8VaquisHzMfoeAIKYxWPqvoU0K5Np3p5fehTMgLusR0he4BjJhcClTKxNw
/UCBzBDk38ubnQO+aJmLcoLkJQNJWb+Eys5mlNK9R/IMOrkTQ6MewS/JM4oCTQ+X
P1Pcz99iKMZhpXM4k/ZETOgxR4WB7bEWVkjhFt8qk+Lr5GxK4sDu6kkmRjR07Vof
C0Hcrc6+fuuRhV+zKkHyUyIaj565dILNf0B/oftntbBZV6HlBQkPcu+EZlfMudmf
8bCljNncFU0vp8UjP8IM2DKf5JBidbluAPmUJ6U7S7FuNnwJ8pcI4EK9wFhK1sJD
5JUPmHhutDVPkz9kJJEBasBDXad5GRrhdWZHXVMmDO3zcIr6oY0Hj2pgVJAhHzEu
cSjdMYkXN4hN1y6wGKYvSoMfwN3qgA67t+cWuAsgxDVCCGMMtGSWe19mJ0OJdyfH
Q7EUoLwwzAzIP+UOl+0T8sFmy4IBWVt/6O+f3VT4kueXDqwNKNaOXfeoGdwPgSNZ
9bwNoWJC7zSpo0Qric1vB9knb9kgpR7USF4lnf3T5xa/g6X1J73IysBDx/PJselc
CT9qWEeZUUbu0rRfhogkBCWdnZkGqwS6hF/8pna+X2pBx6BPg0djWAgIg74BlwPm
ONlnD+Qy9rit5vgPuvUNtGBU3URFXMGWkUKb6xq3qtKECl179VgmMyPc4kvpouJc
st8xGpgl+2UnSqpFiAeMXMJ66NJiXCFmJoZERG/4lUHlTPAt4zoF+m+xfFpb5sTs
vP/UhG0bsjGzeLWFlqRn/F47rP7JzQEZoRoZrEVvVB81YreCXKC/6u3M42Y52UFp
xUnkPAYyB/JBfdCRdirUV9A/hUfIF1SoUiFM2qdXCvUV7+daY/1mkge6GTtRT2bf
Crn3kr95YJsiKR52T3ApzN+10u1NqbupFiR8vRn4xgP4mXsDir51l+nzgBvf8oMA
T8LAZpRR6Dm55h0f3AlKg4J6/CYySuGVw1icCehurbm9ebPCVaTz1L8Wwq8MLgEq
4hgY86v5xOtkcyeqzOop1PH9jd3YRHQnqdwAo3X1ThbtMErJg2W7ZJ1hXQR/49gg
KTecfsBGUcL2Cz5gEezhhaTuCPpGSJgjLD/JzljsUfHFudApNRDEYaPGefmgmBsJ
0n07fnlkhJdjAQj4GEMAeXq6XdOQb9upofsMxjAHkJEdSUbOyuc8tM+Iw5kBpCOh
z6C80omFcA5j0vZ7Sqmrb3sWlukq4sMmfF0e0R0wj15LEn5HS9bxD/2Purk5AwFs
uqL/foRTJvEJNSBYvnj6SCaT3OgapMOlPH/xVHUuiaUb3jcJudYsmcbkMwr+dFOp
tIUxSH6gvWOJfRN3p54B9PVezLUF8ePFFnAAUnBeMaHWD1czCZWdABhE4cj7cKU5
Y7zcmuCHWGKg2KeNjmfmkkvthwMnfjTjvs0URFzxgPO/bjkbOgHD/0082DzAqLgR
FI4lhJu8aQdFeJgt0H018ydMjuQ/qzIHlqqYYIucyoU6wVRu356HIuckutichQgK
G7nIQsRf+PPtEi0vgAhYqG4bUANN9/NBMnnqwOVKgqsru1OEva2fADm/ZaZY+bAh
ayAFVKkC1lz+TNXZHejOPbAF9jCFQLGA6wKgqKzPTB4nIvp4IGpbpRfewNxqwa0b
3UmlGP/H61J0PEBj2NxmzKrGtcInLGO/lUQxeaUA/cu9KXvkGZvjbAqKMbUfXCZ6
P7p4xCZ4iNRZHBL2vfVnBmFXSlhG7z+NpBEJAn1sTKUWVqGS5eebIy5NODBk2T6W
I1EvoUPRcu1n7M5GTulyQeP3Hs4h+lzVIEgl05+3KkZ3CMmhyPTLPgjqMLbgB7iB
dDfulwllUPXWDG9roh7IPXJD+0/CkfYVExK7JgnTSKPzPHmAXniX5Qh5KxzPUcPf
jaxSoKmDx81Lj1d07hWWw5SmPScfY2y72AzC8VBKxyePmgClxReMLsUsY245mVj1
EROKzVbmd3wBakxDKaw9XWuHHd0XwzD41U61RbLnqqyFzIVlx7luSxcyaW3nFssS
pms6wM51V4LrTRpJpHPXLigr4VC5PUBkaUEZPBjK8+owbu8hsbOiCK/v7liR9BrR
GEdqeUe+Skr4WY2KaZ8/2J16sPTRTDXO4JPgM/xdhg8KPeY4m8bgHa99YdF5wXYI
Wk4c5cZIQUKn4vdIQprTUey19+dhoUz9/uckTKYxwijh2vsB/VHZF6fk3c6d8GzF
Rv/7JLNnnRv5NPGyWSwStKNVPuGdxP481LXtXEehqjoXNn8Vg8jiDWCrakldInL0
UeDx8Up7rF0uyZ5Qhpu3wT09qgBs8mt90z+mOVy5Btovs1Id4BMkSjrPQaS6nBNp
XJcRJGDXp978UZ6KYEiq/5Wi4XqsoXpDIYjREZV6SUb0bUmS8SQKJz7LWM+phuW/
bbi+XDXTxlAxDmvkv8oj18dSaiHxibCccy+lRUcjlJWhlx2v+Vin8YyxG115aMFV
KVlQt0AVsj5w26G5fl7eFQX451gBajvYiWfCMObqBAXiP0xfx0Un9Q44xydUGf4B
/wRomewn0YDVSmEYjUeIP5kFXh9iM/AZ7raq0Q11QBLLPbuDFJusUa1obRZljOwI
XzFpYr3IYXpVcdVp9duoNeqFQT3eCuGntDZXVIgoCweXMKSDovUn3L1oa/rBiMxL
8uOsK/NSsvprP/x/X+TWis3xRhw2xLFGyw8/WSKvxS8p7Zeyx4Ucdp89GNy8EPp2
jTMzmuQy3JPatKUSNuv6zoPbKYRW8eIgFbamNaHyRoSWdLQnQsWqSZD/pcPHIEuO
1Kr+RA518tJKXBLpJxc9mAfkLlg2luefz09aZx/8APLpx4GsNhWO68e+9DIeaeMb
QBGKUxmaiygprC2O94gXdG6GUSYHfwUMK3rRrw+spNOkTdXaMFUHYVeE2lbAB0Hk
j+AezBQnhcNm0wKF63ZOV9VcLqf/hYBCcSjQifGd73MtgyjOhn8nxSVQucjixZFf
v5uiQTPwOWrdoKdr358Y8YxRNDA2jZw5SZXf3yXIC2rbR37j26sqGQFSdHplmcE3
Cd11HEDJ5/v/wMlgmSh8gsHRpfW8OqsUYcuX1q3GPjhgzIxGflVn4KZ7sMJb/fJU
7gUa609Yy9xd8ATKscjIXrOIfc7eGNvURGU433PNRzm3dMT7ZvC0A2OnuYQuSSzx
dC0LrHB2SCZoJ/2Mj+y0z1wEHntTJGo5puIzUKFg806CYqrzTxzGt+2GTMiJHE0/
D9FFt2cITXjbiXVYjLiKZiwicHQn7kMg/JEz6XZH+Fr37aRRQWkNAnrUntDsW0EV
QDezToQQiA0OVFMJ8PleobRx4iH4Q6hyXQ/X4U897qiRNmBGiQBRRGtw6EaQ7xNN
ahYdh4c77n/AnKKO90dJfqk7I2HigFkE+/vrI6dyx8gxrGeinX9Tp9zg3FOeJ/rI
4JmsTRDX/eirc27GYsYa2b+YIao9VfWSy7nt1+B/I1TT6w1v+WcqX63u9fpsSS8t
IEwvWLDM8blhJxA1Z4OFaR+k4uHDEreBUmzY8dEOPmaJm7ciujPg0HpxxAB1jFqR
0FoCTI17kHWp/4MkJsabGNgMObQ4l4GdtfQM8BEepqukHtQu1QBYyaK+qaU2XB1T
Kw6U8ittX/Lk16f+gFDEd5wpbvqW/RixwrK5TAN/6/WuJQvUcyvwvJoPkvwnF/rt
eMVZ2gK0/NH+qt0TIBb5LIPXoLLcFRaA/x+pA+d2SbQZH7x3UCn+j0nb0NJ6P1ae
S/EGSWPvPEf/P1zluAUlJKe/63PMMOBpyuUt04LefpNVZ+0jSVLIAPLt35GlgeL2
snf27iXCVcrgJNqfBbJiYWwb89Oyl+vz/kAWo672Ok+xOnuHT8wM1aEWSuPz608z
+8TgVv5dcKSFhQF0YfLCN8IZ/4khwHL/RfpoGAtgrk4aeMGiw7UISmbaHUDKbyBu
O7n6mvix1mrBkKGV3vlODQTsDBhCGabKW/4pbLgBtFQ85g3iRErDrHsltrFdsiFP
SJdmtTEGqZ24/LfOpv4EjQ0fLBPcaYNwI9qz4jMjWbUmrODo4bSAKxSNvcEZm+B2
N+nQn9vKvhJIzj5FNite1ju51RCn3p0yoZwi/b14u4dZjhM7EeCQX9M77NFp6A0L
o82P4WPEItkN0pRiVGuNV3BUZgwT5XhC0ublZYNT2QJgqpAA1JcKiRN0IGEFBV8D
8GXe+yhT5RN6OHBAsEhC3izxV9JAuA3jljqcXm0pgUByGQhB673o84xbqgpohDS/
WCz2Fqj5oMbAwb5eWm0xUqq6WBvB1KC6RMET1Wzta+Tdmzt8xUFCDp3y+pM/jw5W
N0geIgx6iA+bpgVYMRXhfloaf2kGaucc4vON7HsTwoj3kQjRdWqjpmoLeDV3GqGR
QmPGWr0gNatmkFDiAf1ghZdZ2xve/FWtS7jkYU3f2GeQZjrZkRNWmf+Yr0A4gLaK
IBlsKbg7qOyXRnT41HrG8soyGSJeZmj/VpQvf0acoG6I5FD4nMg7dWkxuTUY7j8z
D1eRlwF0YhWZHiU/W+yD+9KHIGJLjks5Tgjn089skffN+nPNZvaa29YBI3Zxru6o
ZmaDPcWe8IL/7Jp2ulExp5JQ65co8rUq6pGR2mI6HydEV4jH9Me3HfKkzT327YwL
0ONux3u/Gz+Co/SIrNM9o+VvyDhmXcaMuCK46TK14cDFmFaqPWXzTG7BlreEts+X
NZrmmZdOD21ZmlnfgyFwx0D6UJ47FddpRP6ZExTKQKfpa/J8VOxBnFo9ODRUVH0M
aq/+CSWMxGLIt2s01bJ+lQ7OFDqGOgrRK8llMJYsOOtCnYIVvQ2On+B7Oah83mSK
36+wimJbLqBDh6hbZcqRp5mWF3jbZ1rRpfRqxnwEhBf9r6QxwonF8WhFy8CnnY/M
SVwkPeSY3wilJrEbCfkwP/8ryPVpWSHAlBF97MQ1tYUWUPi5cxhInE3Bb12YdR3T
Gqs7csVuezeJ5sBWB2X43fBF7VJLtBHeSVtoBB8d/ohxxr5NI3xk3p8XlPvxbnLG
9jILWjqptmNRuolrgA4ym02/tMZeIma7bSJP7RNjG5sQpLCLjcUrGTnrgCCBbr9n
sJTEhKUglw/4GEKrAqpAW5Vc84sVGGR1X1uZi2i6Bq5QybcsejWaqSjYsDgrhcx8
FSyAHbduBhYBeT3mdWmSII+prG5zb6AcyM4cptXS3VGD1bkaW+tktQ901I5PMBLP
qQVlWWkI/h7ye1PaV9NIHnT3a6zKMjz+Gg13WVk3U6sGiM+2wuYKe2q9ILlvDCGh
ogthl96doUFyYV3YWDSheCwJAROUFtdLlBTR370SrkHt3jO1qo8O+S2aPU6bv6Te
tEbDHCj/gVBRjQQDqROx5Aa24vKyBOa3fWVS9emTiwyt01kjP7E4cGUKVUln+JmD
C8luU9LkVxUaSK++dR9M5rLC4QNSFeweaWDGAEKfh6HGOJbgaEMCJa1/gIF71cbm
uNQRO77kvVdI2rOa2kbbmbJnFuu8by1PIcHDdsG3Lph/xJlkWxB31GGCcq6DcNWk
tkOkcOLN43vdlhJL3HiHtSzO5GoRK5X9GzQzDo8bfjVIttUfU3RzBaO2N+H0SlJG
GrODqC+N8xN56GflJVGa6CkNrGuzIQqoAxThTiwFXS8aSKruQJFrrvMMSJliX34r
j27i6+FFOk2f3prWQrU+iduWBKAJgKNs1N0+yO9l5TzarPALakyK9uvpare/QQ0p
vboDd5RpyN3fJej+KJf/SgzJmsj5ro9uZ8CvH3FHCBR+xkUH8RvWaMrFKjt/Ffrn
cTxPPIzYLbeDGKvd3dVi1cnkc5LBCuvZoXmiO2plGdL94Wzqcf9jxVYpguyyGSr1
a2ZG4mR2gOdB0DSdoAVv/UEKhdvD9x//nrqnwfH5vVa+PgOtulu+nunzMoGPL743
sN6NOF1I0zOKKi0yYvfIlzgKsKoqVzHToD+5zq4UmnQT/hlhAsY20LFP+jPB+OsU
UdT2NVYube1x60uPHH68S+UHybCa2klEkpD3GN4Qn1Cy5qf1sQ0TdiFaIqCFZsw4
lJ77tYs7aEtW9072wXsMY2Aqp4ZjhepG65TK5aLcqDf1I0/Q8Ph3oZqSTyOzaS0x
ai7SXtJ0x9dj/TBR0J44VFFVF83Ip/VlcpAw24QAYi29x9DCzvKJ4ZjfpF3+WBPm
gEXTIb+uYM6P8olEKSCbT8a/9st6uj5AEtiUg8KPkzH5XEjdm1Y7T2GTN6spEFJ0
XLLu973BJggMZVOGK1VFuV8JpbBY0YT2sNyKFg6gjiUFOlLJRTQEXT6r41NjkiLB
xoMppzKNynN8fdQ2I0gTFCaI4FL1MzHEBbRH2uRSIovIzp4oOzuILGiRW68HD1l6
KSGaNVTdcr73dVcJaM2U/Ob0n+JXGSH6hiREwoJ1j3pu4P74zRDR2I1cbR050u/v
WQJATz5hMMDbghxYRZL1bfpzsYMmTwVBmkQLGqKJAIeIbx8rU3agUauXVb6pGFcp
EyZrzQF/x6dRL5vQRIrZC/MS+cln0CK9eJNgxF2JbPRciyPfuMviuzKv23fxwyCi
htLj4n3VUz+BiYjyOZ+rItnTtm4xzTlYfzersgpC5jPVo86eIuhyCSVnLTk0UjuO
KHjmj+coh/pZEq7oyrMR8nS2uX/kvo9gmRq4BDSOraiR/9vAxpQLUCjcK0N39JRS
PVZ13o6kGzAsFX34NTWYAlkJ7slT/vMPVb9NPOiM+TUZKSH8SzrDVPkSTYEd1hzV
fx7NiYn0gcB2UigLxBFdvwzTS2psAV5JC8TimkWmukDDq6xKHVlK1n2r+UEqNLl7
lSfd3f6fn5YYHmwKNv86jP5qr5I4RMIj8/N0GUA0Z7mwY8ZwCHRUK3Sd8rRp3pu5
5lNTht50+uecbGwfrr1EBs8TUF3w9hfOKkie4+iv7KTLKo8xGZm8Cyg4l4YNlfT6
+yIs9XJdO70meEzSb9ZhzPfpMkSaTYXUB/8NWfLBwoyNwpcU1YlNmNN7MB01V1CJ
cor3Ye9EQedm/raO0gZarjhIlqHWFRrp0AHFtFzrSr5g7WscaSQWgzhSKLQ7nynQ
Dvv6c/OiCMW5erXk/m2/MfsqFJaUM/pN6zBQ3BgluO0pc7RoZdeCyqzc5TYPlGof
vWCMIOFkBOveHCpgYNEDzed/se4wEyF1JNmFm6RYwrYsuZI5mU00/P2SU6GSx6xy
3d8uHdsP6JPehJ3RhlsNnXqS/ScB+GYOfDw8YVS/MC+iR5gBLRlDxk4zIeRDKQNi
b/rpCGlEtpTx2mfQ8pFGX173pHk2VvfNC5jW5xC3vJ27Gbo/DEQFIYCoIepEzSTB
rSB32xx2QEC/u2M5BeoJ0Nfg0+5D/skWhvLUro0AufVXDxnD2XCOfS9sNTI2/8Kz
IQLZmK1shXwHkyMJJ5/wYncsosrZHBta1622nlG/NzUzoCUUTKkveghp8wlfvuWL
3r3KNSn1teo868X+PhA1wehxrdNRxXo3dX+S6nqIrBZ0KrFr0Av474VWWDMhOmj4
IInU4dSGdcgP4m9To5E6Pe2Nm8CdmpzDBOZn7pSqwqZeZC+qbwQg638p75B0004u
vPfmBmchEXEEa1Z4XDVgowo/s8Y6GcbfYjXLEfwP1cMWoND7FG8pRJrcGPgcj7c2
6O9EAgcrGf/cfLc43VNKUQQq+aGrnrUQBiBAj+w9bpnpVIJsx/X9cpf9cxvMTYv+
Zpyth/UY9v6KfEffYmpCFjdoyCGXdi8NpSHc0dcylSaezGRxvjXBM9u+4rDxQ5hm
x6BQzPYHzem7cycSqjp0K+937fHtFTTKkLKz9dUq2ZdEMJkj6SNfrNe+sBDm2ynf
Y0ef854PtMpyRXTBs2sfmTL9X3vnw+X0JyWc2mCNBAGGJjcHWhzMivsle5cjgTlA
V0qoikvIw+/gN7oVBC3id3lDC0XoxUQ2dHDvYaxTo4yMUrXUPovSIYQ1lOprbpH4
Erp65iEoRqW/2H/sRqTaBn5dLwHx2N1iNcFniszarwgKZEGyDDPIgyxxQGJtBLyt
R/ClOY9fbgfmTB0pt94yD2Hk8kftLfPRtBi8xf55a9jTOaMUW4sU3raSasFEb1hO
57bN6M1LsNsSFssW4+HiQmNyYbSko8/UYtKIKf4gWcitTLtUU37me4kwupDIi42t
DrEpQibDbcPrU6hReks2dTy4RfcbMULBcUTolqvdGo1nhYD1gYXjv5IMXoHSxm3x
EDKrfoNWaWuOLum09DPMyeO1OGtjG7sYW/fatdYB8iRTLGqqVqdq/rPrx5FEFsN4
QDwjIvxP3SsDZ6CZUOSL6axafhz7rI2kT1HKPjziDFjQDF/oUWHvmjGBhvEXJ7hl
AFzOJGhVVCQu8KZPt+DpMr6ptbFiU0CVFxjd+Na7tALfdc+4WpGVqNk1VePbQ4yA
rNRz8X93WQGogYEG4Ed7YFU6MuVPFnaKvyMIPltCb7F6dA7C2UzXNWGOVjKV5oYJ
Gh1g+zRjrFX0BRpFhaef4CNznxeIEA/QJXAwKVLhlS47Lz9jomlyfQLe54cGtvlU
Mbjn+XFiscobnMjkqZXpXxuXnpoTER2vjI2AD7K+xjXVK6ScoF+yhrQBgr6URQ4M
vhO7Gg+oIb4UTeg4SwDfdJA/vZluzZnyyzo/vRTkY3JapWKyrViuGj65pCDmCrGU
1r3FrtkfnTesyP2s+oyoFtB5Gl9hMU2y4yLPho+j4iWznU++0I9jvFNDRrvk0+Ck
6mNeEcRey8gEdip2fGlT5udIMQsFoegoh7h5sL/5ZyDD/78JPAxX3cyn14gGGfnW
6Cy8732pgcLjE5nevYbDiuPGxOyS0mtuI+/KLeFBm05WTEq3AzrVMKODtCdC2op0
+7Xn0DcI0+0OnNjSkLt8W1C8xk6IxAq+qd7SffREa9JgAHHUto4Wnped6ZlwgQRC
QZ2ZNSsJDY8uCXxc/owhXPWOx8mUtLWi/UJ6GsjzsRKD50KmfU6xMRHCHwuh2otL
b4RjDHBzWspHt3pEnCnwvmpcOWWMyGBm+weOwpmkkhneCBtf+Y3G/kmR+BHnCmGQ
ke6qr+S5VCsrTVXHHIMSuu4w9n5+WBmFv9RqvzJsnVrtCiEiK66tqOsZJE9UDfqv
OI1EQchlCyObqNNUqi6iXMrA8AJCb8QtyM+cd2hHJjDm5FZJfAKwC/oxfQ7iwFeQ
RngjNeg41EKaUf6zAXN1vMrUAOuLVr/MzCPnFRJcpO0o/sIOgLI1vzcf2Kd5m6m5
R2dKVBqP35to5wA5fil2V/A3rSnqhGm0Ot0E4UVT7UcIMAfWqNWmHO9EkoY32Bnk
ACtTF1iWwWDmwB3GcN8t+RE7j9kBeRTxsMGe6+wLERCXnj4sp5qWkTwGii5Zn7/8
fQ2hcSomhz6bn59XB0n/rPXPAo0qNc4VBak6sAqS1AYQVts+EYIqxEVAmxwjvHhW
FF1vp856/9GFMTS+ZKPQOeFNyTEgn9dZrQEd7mInafYLPvbvQ5YvrTmW12Cj3FER
l32kQk1F8GB5ltfPF+rrvTm/2Bpfc6nAjqNmLCOK9N1tl8MZDLmAfVWFRyNocI5Y
/6mAofwcmT5FRBilw45JYdgcvFVe4SUYD8pzjNZAzAwIufpVm844fnr+SCd7htio
MKpDY+IScSFF5+S0b+joasX/kx8OTY3/0ftu9SoKcrjxYEXJiFSkrVjAyi4KGnr/
qQ8/mhr4bXJ6rSSOYadAEHFAQvSUoQeYn3qiEqiTI/vA1SjM39wcigy3EUIkg30w
azu0AQ+GJeuJOoBK1tJ3o2sC4KA1Pn/RatVSYmfZi+BaPHdma9Tq3rQ3E+B/vpo8
K5vxbqvTXvUvqr9YjtQMSz1SVUtK3fIvibZB/fUyIByxuQ2u2ACgofLTrmLzcozU
kvIfvFAUYlv4xf7VaXUrDMZPw34Ot07MYb8tyU5gsbYePycFTSHNgRxVY4AOwooH
dQBe0XUFVe8UTFHCtrCrPF4WGBo1JloqtHhhrFpOca4m1cHG3fPOwbbcDdoDKWKC
RDB32fXEWuvkVgo3wl4QcsETI4528oVaizbCnyBE266d2jRBHAMUyue5hmnbdeC9
dScabQK2qNXSCUQsRk8BrrZCM0NkOVh4YJunSnho0hDlX0hmve7KhMTAOIufei/q
3FCWrCBZclT1hpS8vAVCUTU12BNxTEC89R9LdY7mfZZEm1dmeh4R6OUMj8LAVhm1
bUXKmB0PEL/ElsS8VC4XNf1gw3denGFtUyFM5t0blITYWpEdgZ6Mu2ZHcUIiB09k
AT9/eOsvSh/IGHy328spaTYfPMhGOjV3R/6K3JJzkhrw3LpeVV5aj3fkl36mKv4C
YgcUH6ChTYajy9NKxLOSbF5AMtP3A37227C2L1TIO6gHJfX6QZ4ZZJRn9u5ZN5Pp
Y8RnE2cUYeapY3F60lrA2q0KLJvfOeQaZvxSPjxQUXMqB9XAGbNeLU7Qsp6a3RAk
EktvNswiIIsBKeE5DhpIK17wKd4KAQz7JNIRdrxQCexKAzEnH4lEtb08ZrcNYzx8
fOXZUUpZVb4l5WVSQ64zyG2CnwHf3GDMzuFKDgIzkUdIeHIgx2CRsivhU6vVXTJl
dI30M8eZ5pvdgLZDxWJ5hmaV+hURKKPqQFSjveyAIcyD/P2r2+ijZV0qyaLkiIIM
bA/KzqBLxPWYJ3772L10FugzfMWLjkcRhLTrQTPq5FrnlsncvN3MieTELkXmn7qp
lu4aHR9xJ/3N83Wvck3fVNxVVrY4MZimGpX53czonTkg2hPvaRLhQYn4haY3fmEA
eqA6uUKxJsy+9TwTbE1KZHqhpZOpN3jlqd3Hl+R3jGAoEA9OU5AKAPcd80uw9LJf
/FXgPDq600Vc5q0bMRqbc4GrEAxsv6EHy9zhsCbO0vQKKpKZFGxjQu4d2Ix6axms
YA+d7bkJUOnR0j0NrHaW3G8XqeZ20SdtntvoE7zHqY0AzSeixBoYXtH2cmBz85IS
PUgLf7ls6gnPWYWlnbxlKnhn5lIfeq8mF8kM1kB+aw7KbmH6QBXd/Z+AdZ60kgaN
iIsHk+uerePElnfLJx22p/Ij37UbLEVfM6FIBlD0sqU31AM3Aawrj2HhYS60mu0a
c4mH4BKkShS9h80UJoYrMwmgMP+plLZlv+micZa4YoIg9+qAsI2PIKEJzPqRPjcc
xcrVX/oIkS7JavIJ9Cn6Ihq1s07vZ+L96+LicmMBKN3SDXdZQ1jgZCLwkU+a4HUZ
sxR+fb9pZsDEV78s9YQBXtbnrc2xg1JMxxdqGQZimmlA1RPKbm/0N2n/W5MDaQq5
xVumiAcGeLrhDdzcYfgV7md20+U2sJX3aavoR9zgpG4T4lHaeolWNZCmy9eREc58
fQlJoWGi8rj4dPEDUNEALol/CI0kLWI+bqtBrkWKmyy/5A32LPNoO4G42Pu/A27v
N2LLcz065JJl3bCUGmMn3hX7Bi9qKtlGMh65uvC9PG5ffaumd7bWz8klF/S3UQQZ
mVCY5bbvM80dUXUK+PenKRPpSJv99CeyNMUb2tGIwbE6MMykt29mSvwdi4NYnHGh
qW76FAxZS97/4v/8g1A0Dts09/VLdV3g2WwRMZLjFwdq9ymviBNP21pErKwNjRTp
coxiWvAxLV4pDodmqTNSCUyeHAI91RyDKnv9zl/TmupLbEtSNe53mBDXx7vmLTOP
uIiehnlraeTUftLoiKCC25mCQD+DIqdMospqyDsShI1i6jBL3wgDxV4r+kQB0kh/
owKpfxC4E/NVNis/z2r3bhnS05jrt+eDiOjUuIVuhMJW8vpqRYj1Xle4kGfAGlVs
cM2c+7NJJMUaFm1Bskw3NlWrSSnAT3yO4e/75q814VQ10VVxu3YN6fIfnNqzGrev
4BzL2cS1NhUzTXewzRNBF+W6DHPlB3MK5mfLELLdRB2Oz6D/VXFlKFSbPa+2jGMp
CaFQe+KIvjtQnanhiaqPUneVO68z98lBh+87n260oEavy6LN1kP20oLKs8wtnZqU
Fn50PDvpseZMBv69eslMJR1gkc1cSYph4m/oYCPddDVIoOO6kcN6bBJRVE4zTGUM
lIEobCde2CmPWj/FVTn0+KcbYgmJY13N7Yv4dLK4nJhK8HDXUc1Joo6p8p13UlLp
KNsBz5q7NUv5bIs7B/2aiEpLsLRqFazHDwwi1r9ffUwbVHF792UuBf37Ks++E/XR
1HkoOklKFWXmWoH7NwksGPmf282aveJagJq3Tb7UWoaEecpylDC8r9pYNM3uhDWl
/5++U0Ky+43zBW0PGxE+m036z7vWgts7SQKmzhTG/wvd1ZIz3tS1DZbIJtf9xQmH
52tj8A8PELP0OqlbV1LmVx/0/BSlDSf+uSS+/KeyHV4ijcKYCjQsY7aHSqv2Mm0b
A+vaQHwVNYNYIxXBoeU1bcJFh7mFPB1DpweE5+ZoKL1MMOgLGadIRxUtYAnXprDe
fQxSxxuviF2Qx3Gp6TUvaaMEohj52xTpTR3VVYMsicO5qeQOwFCFiEczOCcdWJTp
lKNY8iOCcEHZPp40FXRMnAQ80E/N5zmipwhiNS3CnyldHR1SDECGIRipWjpzVmma
MM1JGSu6wKAZKdN5RqG1nY6MAAWn5hOzrJSUrKClmVQ/XZ11PHnMmSWB7QbGJ4bu
xWKVk5zny8n93bKc4fRh/tGvbCX6ObAlFTMIN+co4OV/+kl1cpkt5+TMElqiJiWn
3/jMHk09PH3xFaOQa/v3YGqSK0zEIUXpBrTfFrBlDwERNJa484klIQV6BEpkn95R
k7Y5iaL4cAsc94o5T9ICeZJYkXAqVbYgZpRErMbdwBQG7nBdwNxrnYbZM1k56/a4
MRHNJJULg8X3etO9HB6nQKb0L8GUDI9LTEfH+oz20vySh/JTvz3u3prNuLE1TjYM
OpIRToi99R/0VuvkRHR55kERAHtPlTv80/BR72iipW+KoCQNCEHUOIgFwnPyVJp7
8g0nxhR2IgG3BZfJYl6hJDCGUK91zSqdnZFoN1Ct8RwdIRg+96s6nH5ZBeBZsz5A
yve06HNM5q6huai8mBJEf0n7qyeDl+y7bbwYqV2iVnu+7nF5IW9c0rJd0zuv6xoJ
lSGnOctsonOzugPdi0ICATkKIOlQmx/RegpMuAnPrMz/kJeL09bDqZBnXXDhfxbM
CR7l6SU/O+mB2c+xmN8lQ+b/J7oc4R4M58yEsFSBZmwoaHtDgQyu0kdGGuP45b7h
nmcLsuF5VL4DhFhtaT01PEzq7l/EWYy4F5JGOCAohuMH7Kg1T7ZHsvSTumAQ+RcY
/jXHIby9oW6DI9sDyNkUsWetIKVq2V+84tzWggC4Hq78SpTjlqRlA/kv7g7b+Z4h
A+NO2+6OoppURnIq17D2RYt/uK0zS0sacRP1TQCf+0UdEk5BXQQs/nD2I1fCt85a
Sz8C2/flrIvMVXWz7oi1m4ZeCRmfInrPwxiFgtg2dCRa/ZEVWdyHMHkzhYXv1lQg
FEx1kcUftNiaHuZ7THZLtGeOX1mmX90Ewr4ULFG2yhMkGPQCF72AuMINv9JwnNmp
5Z1TM9dzGWBB5C76DHPQQzCHM4yXQaTVCuGaBeYKTvC/eVqCfKeVCCHFW2UsEVf1
jLtSmaWBqxA14ELTLPbNrfFsMKYkcI2P8u9g5CEhhp+7Hg3DHnEzxK0YrK2ihKWy
hqiwnSt6jN0crYOq75mvcIU3LEtGVTtGI2AYrinJC+zWxXAdQy6qESe702k5H2AO
XG4sbbdL/fAw69Wd4lL8GIENhLkR7lIkpRtCjVNWc9sYOJbVPM5OT+NQertZzuw1
m6fENbIBPtgODURZws9lFVGEtSkN7VqdZVfX5R1zmuTsxmPPlUuJimWcEv7m2t0e
U21zb5Lka9hncCf/KQCoBEyZQan0QYV6lbtfiqmEctoMPD5RIcgMHVXEx6FstI3s
eH6al4eP3Ea198pTaRyHtgSrnbXe9cuWkvjo/oOmgPVK4LsFP6t5JQFsTKcePek1
/lyAGB8FW3FCxW/8ygOvTwDnVhfO/AAbVzMyCmx6aTg5jh50aZoCAy1LuXwyeTWb
cIq7lSye+CJ4EHyziT/L0OadKg+9gXKzJayafW/KnFWKxIytZwSzr9P3sIe1RxlP
nRmuXivOamt1gtOo/GlMDiRb2z98PbG3bqCBNm5LtNxlHTn7WOdgPs7sv5PHQy6W
DXFOe/Tn1Bh6Rx+RZeYtPxzq9ZRc7Q5k32s12RrN9xp1JleTbPpihTkJ8+yYKi4N
kSqc7btVQcNz9CXi+aiaAb3LSgHLC6dMJXycgAzcxCPhRd70NbKg0qpNoyuG9Rc5
ICHYFSY8Elv82lG8OJXqB8MvZPLJztsqNnocj3wL0NRwKyNGWGvg4+5Puc5Eb0tt
IfGjdUwNj8c2sMuny+iryH6hlDs/jo2l2s5F7b2rDiDpiSmptr8rqtIfqVHrq0Ee
51NYcyjhjmwxDPDtbyuelHJi2k3PcTtSSTMFyz9m8wFdQIEJwG4SQuhiEOQjYQBH
LbBR6OOkq6efkQ9epVCJ4ucLP1zcZDa72JyDblXGGnPEsBJPRyQpB+rj6HOXVOW7
btKDv5Hl9fPsFdKRYScXUOqroFhvgMC3P+tDFRsjdcU6fOkaBfATHzZ9JbsH/5GZ
3eqdL8sV99OZCeeDX4j42+pT/RWmRqcFaAug+SUOUdGsgs/u41/R4YBi7bjeEc4V
PP/Cf8WhE/c/iUJsKoFTl8WgTQvgwfcCZUw6EJu1wA0hjkcKzVDq+DijmZhO3GhY
NFPtJJFa5HfdFekwBW4XIjaLP/17znR+x1i2RoSE0BFQ5BdoW9+f5uffBcHFW9x/
5ZMfV4UaCi9kQzY31qvq1eSuSdaxcSlUcrzHycjdLSvw/Y1+TTUWsH8+A7Ro3IL7
2rtH6PIzZ6PVzXKlsNsYjFwClYV5BkXlpSjXIAmSEG9pApSFq+J/0NBHo378RG0s
SzNlw6WGrIG3LCl6uSm8DvowhpuPIpO18xXOSc73bDAbHeJXTsuRzt3B7PqPZ25H
WumxFf0k5wBC/bGAIu4vTHNgyAbwMuZAX8p345Ly4bTHmm6+Q49HbbWO1wzxFiqE
9eV6ZKu/SCf8L8k34yyq5yJdnhW8WLjO2ceN6TqnpJbHx2rmJyfp0KILI2nvSVWj
Mc44aL9XbHn+SeFdxu6YDWpVl3vO+RTY3xuRlaBzTanhxcuXVK4OIvPlg+sS3qax
3q/7pzOpAMzAkby8N8BNurBYWSfQrAoZTBEo8oUWMecCE5ntKofRU7ooY6uguHks
lgTEmBVlouw6NnIu5zI3ygvvet/iWTjRkfMzXunkpiyhRHkc+W9UzAtMyQvrIMkA
1aH19xXgJ9/LdTat4s10RKyJxPkoEVVj+MrP2kWWQniU64t/eSYKpUNYLUB+26qV
LhKdow6mEpLGyncw8v0rtSEE0+blTlXyi6PBgCn/MI18C40hK07Fk2c5ExOiS9ug
ocys9C7OEfZgWDluIPaRWd++K0K2LJ4cW+8v92Bwtiokfo9vz7m7HlrTG5bceNb6
UN6qOaYflhYs162ezO78w9Z4F7id1gySAo1FfiQ16mUJQXw96+jknRaDgyutLc5F
1ZhoKYppxeXkbIOymC7uwh1Ln/wRRrXpiAaiHkq5l8gsL0ws9OhIU/QTx7tYWzat
KJTkRbI1xvRsVxLbZQOCGggYhTk5A7uBHmmXUxE7+NMGfxX4qfAJHTVLHt8JcUl8
td28ekWqGGXISD/zGCEcHgZY8N8IwZIoyhs5wMUoTsjqJNIuTuEUR12N7wkWhKqA
0a3LLUWqWaHJnOc6ChYmpd8J7gV0DzX56uuqLP3Ov6+bROoT8ovyE6zH5pu3Tg88
L0771n3ufxHo4JGL2cAe/1sdSCnqdxyqAUOMWMfqQtjPCiE5KG+DOXVlaTTVpr70
373qp9SC6f76m0L/uKPkipKwFRzhamHjLAZUT6vk5489Bjr8cpm2HNhpT/ndBOHR
8VjL3MKzhJaBgQp8gJdTClXtsC19p1H9LifcY1r14q2AA2M/0Eahxb3faH7fbNEg
8jXyF1Spzvc/EPuJmpy/w2KSbeUP+DaXEHApA3Wq1zzyqOn8rL2lYNTK0lRoJZWy
jMTsff0WusSeJvQlqqvrjJWGX2TRnJCfinFkAvm/aNUcTEBCy/Qx2LQiMWurxal9
24pKOgEZUuhcNnxREbVxQkukLHdPsoynxQJh9AM8hKhIDoCWAPCTtkIC8fP77UyC
3GupGnHqxK4vH6mnqKzAbzor+UGcUnYg+btpgVQsX3C+uJm3mfjt/XXSg4inVq0a
0c48D352y/2hSUfylHwLkyBgv+SaiZSC3N4/5uUtDvYPXWZ92PIobiwptTjr0Vbd
Vf4dYQT6CGqdcvJm0mRye/FQf5U1WZ9hD2G9fNdNDAKWmAjNbMxGBcllsYHpjnh2
fkrz8QRU2c/CNd8777KxhRHSSeN1oV8eRmPgCPsGXCx6tJl+t/Ij5sEIK5aOJADL
S+WKjbG+5yV/QhyF3fF+d4CGj9q4G896gETrzAJH8kKUxfCrct11tRNJEsdu0LpX
4m819QXLdfdQxbtOqtM1PfLcyHOTk/hvjCVVM6pb020O2kCKS5jtezjgIWSWb8Il
uzxXHg1CkZOxlycCkGez0Oo/apksu+4086ZFr/X1tWGH1ImIjUZRKvyDDH3vYc9g
2bnF95xwkJzdtDFR0lTvTfvvYD7DO+FcbKwERnsd2CRalSwdE4H6PpGTZSKhnh81
mXkxd40Xks13YkPcn5ony47SozdLjQaYDgwiwjTJ+rvZLLe4dfVZQjNxH+NgDXf+
Y+h0ABpiWYtMNNdTRDssyveha7rFShTu4aTg3HSTUjTos020vIPwUca0mRAk+g9s
cbPMFTVqrF/wyksFw18r5xI5aMeu6zN9AXOUBr1TbhJqpB2ZVn+AoQajIAtSkkKP
BHqD2iH+5b3w8ilyBubmWVlv305EwGVJ8Gwq3D44ZeC0YkvoNmuoeLcYKfw89dcA
l1XdQMS7AeZ+iyZGED2BzShRUkWKpdDyjeGf5YJ2D0zSOLeJWYA+3RhtY4qhAMYE
4WQ+9ZnGu8oWRoJ2xtJHfEysLQHmP0zqRhQXO2WKogG25QK8UKiSxHZaZvCLrQF+
aWCuvrEpkhEgcAR6PyBAOJISwRS3fbOnb7R1Mc3kBefrudKF+rxA8w7a/ydMYzja
SeqF0sBgYg5Mh0BRQsiZGluSuMSYcrNLedfL7Y748ZwgnMopa8wQcwzEHIVXqsa4
NvQpOYF1ET+KwxbmSfBj+22BxSAtuJRedHueVrAxE8fKlTbdvkA2ZjPUO3TJ/cDX
eC/nHa52UcS4c23ALdwZTgU0Lmhav6wTvU1xK+iT3yu507B0A5AAr63AvO/MmzSe
rNnMb2Iz4tGQSSuWWNF3KZeRVuzRG2pzWa5hoe6rCNLTR7ebgI1NI1mmk5XGGtel
eXx7uSvO1LOZV1YVsgChEJpVghHxe2EWlhafb1gKgc81TmseBO8fDdilB+oLIcrZ
zAcmWDSYw6+Rv5btvTw9KkW2WZdWBs96IQ5I6u11xvbG4DdMa+8OkGe8fEFp7qsj
l5G7EJu1FAG8kyg3pqqdbBEWvSRnJy/FGZj0VwvScYwURENZXQeeHifpSwA2KC/V
x8tA/7qblhngwPpJ7VIPASlcfxS/+hEss4RvrsK03Ihlm7L3oH/FRmmU/hBQ69wf
FabZ4um8o2xc9Sm+cGf+/uBuNOf+MwjEfbDibMeMLVOyNi4CcSUoTjY3m6rDwJRF
1mgILpKJsTAj/WiN4lR71j/QU1x8W6wJrqggr+uQ6sgkzfUtRFCx3iy7G9tTR6/J
imnN9X3p0jIa/DSZt9XTpakLvafqNIvSWZwVgx8flAUEO0gc1GtdC/Jo6pD5Cc6I
T/TfX6np0xIdNP6N8OJG/UEnc1DnzQy4YHeQJuWqE5btAmxjv/+wxHw2ty2rdPBI
6ZAsaAtlZzKxcg+j6NfeeCFu7QEsFpSGaMZs5BQvY5CfMFfxM7Y/woOi8k9dNBta
4BfKHrreXABv67Fa+7OzvGPNUjL/ud0FvxDEJzckivG4hI8oQTaCA90ngJ0wVFFk
SYrO6ruBhGSo5TMnm3jQ46h90c/HigBpDoascjSm3WQbPbxoe450z48ZKkKa5kb/
mbkU1aD02cY+a4Ns3BqQJgOHcPE9p7Sd+GSlm/2nkcnZAdP1qAmNZLjP7/pxzBug
MDa344APwIE5T1Zp0SnydHANeuMwZhwI8z13xkp+o9aQJ1LU8OQfMCWmI9SprJbH
UPjRu5MNJsQXrJGbpngOdrw6tnh8ddOTczCWy+oIQJyYt1YVnTSL1WGwGX7qMp/k
hIhDjbCZMn9wOWfa7ljLsc1MUByNlnroIWkUWRgmVH8qrhDWqv/IyPjfZq5w7Ikd
hYOA1CyauKZacpAYjM/ZLaZj12cBOq1NjQ/zfFvFQwB285lLwGGtgn5fkIGoMHCu
wMmP/nYa/oX8zgwKOYf/qIjfOa/2pxfkrBfE2Xhnvyn3JTSxE1aUW/ydZ3bOCOU4
JZlYldTXugeo3Ky7ts0NyNNVht4VrN0EIUaLLbOuHcjQJOwcwstysUqX59h+fJYK
pLnw1kWO300gSorOZ9/Th5EJcPT2EBahYgag1da6CDP27vq3D2WxP2rVgr7hBIYG
vjpjYXnsTr45RV8JqlpTtZYGS1XRXN3+FrIuoUdu920KMIlxgGZglG11v9p9V8Tp
tXwVVMEqUOofIzh398mrWm6inP2HK4tlk7AmQULyeICCdS1AtPQZb9PB/0u5dMej
2XxVDp+w+VwafCrsC6iKbqTQOj/Gjc1N/WP9w1wstyJXD3l6sbDFaG2d7CvQU5o4
nwBu1mDIsczKCvlpOqcBzFUb/+McFB7WW4134vhBSVu9SZKed9C50xZ6rfjktz5q
jCW1hX0txfNi8zdiyqWVIvtI38fJYIIvNLvl7McaJDmjW6YzO5jCe+7QnU4vkvmd
ibIOzw4bwmCyDRp15+AWNOy3U5E6muzW7Go1+pygCNY5D+uHYaX1lCQaoYM6gN/1
MGqpdhHG6v8mIWXw7Cd3SsVRx2f5EWO8TPCYopr6ck8ckwoEV1bOZg77ncXfyYzF
anfOb62u7P2yrN7WtMXkFlQuKfwFHUv4psvp9f9F+yqRGL6YreDiDZv9Eb1N9yiW
nWRPhyhy8HcV1djeYhIiAhfveEixf8XeDjjbk2+Ej/Y+eejQLl0AzVcKvNdsvrYn
h4X/Ijas3QxBJadk7Whr5reyn1glZsVAIrMQs6NoZO+jiBd9+rPBIBKZWTY0T3by
HadX3ZsEv/PvZK1fps8NL9w6pGNEdPpEW0cIaz2aJeayChz8W5GJFD1HhDDAMzY6
pUpv92sqe/+X4poyaiMxnTeNX3Gdb2+GQHX7KizdM9N27nmtxX+1KF3+DyQNCSbY
Wzv4/XE9KdzuJD4Na5+YboNwz81bRGYaKDTEucf9Kx+f1WW44tRogaHKndMClMtM
2r1Y8e7UueNSPzVsfHudByOPfkeR83JMpmumRFeIt4IbrEhxLjM3tAKNhB7nuGrs
rYzfSmlSYgJD7s9B74PeQwPsMk+FX+f0MJSgnRWOV2G0ALzZPoPsCNl69DuR1tpO
5KPO5i0Rblppo3Xal0eciZF5AdyFW0v8Uq2fLondo5z3jnQSlANWgYEUk0HdTfSs
D+43yV7epsaR7y+PAcYSc3CpFx08iaTxKjw1mz6NdsXPWS6aalwKPfegv+hSl3nC
qvVVLUATXqF90Xvc9Fm1Oee4fjNz0GL5flWpwWzL6lisgf8ry0iKRIKc0kYsZghn
Dgirgw+C3hM7N3GZ/vSp31nF8iKh68nugreIWc1QTRyjhYaTv4BKzqgbVGcuqBxH
9LGnxRQ18SMsDj5WDH5PrHqNCy2MhrztYUmqYTJbqw2GKjTz6kq17IhUJR+yBSaF
zLQNgYhrxJLTjpNeJO32F7F42EaWcBnHFKFkjnsL1LIpv6BQWUu3q1f42Q8Y66Bw
D+8LSZG5Js8QH8EKX0uzpaUIKNZOxpfrq8wRdMkGZMMBjUOwFTtzLaKxLKdzC9gT
36w0HtA9V/dxelHaJE3NcLNBGP5M4o2KFNq7uAkXVkRrEmCmQTC9b7IYCA/SniR2
QL71Qm9cMXO9R0R0HRWgPorKDdkSnIOFI8iXLCs7d8wqCnY47OTBgwlv8g9u+r38
Jz+piD8B5ULaDaRnk4Q28y9IYT8jkmny/tuuVNeCE5UyHrXNJ0Kw9q0hGYBPiNCT
Fx6NByGfqTM5vASWbeq7sL+nbRKzDndeGNrJ1ei7wIQv8Goax0jpUd3P9LXxK2Nm
duq4aGV2jgJAf+U2T1jklIqkTCd305S6Wn04xAvsp1tzgLrda5DWq/Jb2FQoJZ2L
cvshLslwI8NMa8RzkuEW28M/LGxC097rKb5F5pnwi0MI3+SqRu9gGmhnIWsAh/II
A4nMjAoJ0dOKXsmKZXf/LngBOwGO2evUbLwNyuYgFArt+t+vfCduoaK6zkuFRu7z
9N4FoXk2ETLH7fLYN85cvw74Nfe6eRY3XeOejfvvIHrko4PUMwYxgfh8KfpaBUBT
nuYGg0GrCe22B4F++o0NF9g4pANQ1e69KmoNGsmuPE9v6QQZnqTP18XlHpfO2mJa
HrfN46bdUmSs53C/e3L+Xofc7ulgVPoYiG6HCoD3JxCKgREQ2R2oAjbZxouqJRKM
d6ioGbqElVMpds6bkqPY2xQHEdsH/IijC/34FC8pYZsGytrmSIioDdIILWXelaJ/
DR/D/OVmBp4mPriGtr0dLA+2VIl4WoMkiEtliu2UvQBp7cS5ccaU8IQsTlYrTCg6
gDzvDtIfsDgexHPFkVJHS/WWTCvvwbjiNBH4a+Hyr1cGLCr2vkS/SGp69/VRoqEO
CSF5oHSzxbWYLhEDsynSIVYr2by6orckTSi5VxMhtu4GNHN5yAqzt7DQopwwxQLL
EuNkT58w6L5yKECh7YAQkcCuVo38Nw4Yeur1W+RDFRolZS7IRhT/ucbDUHu9WL9V
7m6IP2DhgksNOnTtubJ9ZZ2MgSbvyYHFlbmUEdbozPR4EZEL9GNqyaV+jenK8RWK
4vKY9H+F69jEtCsXHDTinzjwLZr/qnT537Ua0h4wssgjsjGU7g1DXIA23/CmrOH6
p+5+pGYd4P1NrVcLCpBC9vHS1NBrN/y5dUaFA0IRC2O//wGKy4maW66wLCT3kMst
cWGwQo0vHrfPB5nBozOXnR4w27oWAujDxCEXm4LZU3X7Q9pdec5N87u3joM9xSyo
zcyhnow9e7+cW/lL9qXFuUw42x5xINOCXPKn3qZ79i1ZUAnjivOma1JLl07mfX75
d8NP3RQizOmPQnCAHAAczEwUJMGYWEa9CrLb1qXcDRN4rBw5vcrR2a0/Mka4FLKb
ZwTZd+gzft93SZtnWJDPYOFrcptXnaND/WHMIgX6669IfkJCtTHdRw6OwEZk0bJF
sV43y8TKi3zih3MguN3jn8UknSDw76tHKhhVX3EjpQu+Hbm70k7VLAth9bNF3KRA
Fpd2/1DBKoZ5XVCYdqgJI+2RUeoKbiImjah/hSFg06CEhrsQdex3sONL4WhZSH6j
bDnFLcSy8BW5m6Av60O18VtEhPu5H/kdmdjeqJ9FIZNYMUL1tqtTQ3iRjqv8Bw0A
c18H4vV5/WyJyr/2Q1PTe5eMDqn4nnSf6T/0Y7l+qP1gU88QTZHEN8O8mDKYynnF
xNsPkppmWpZ2O6bmJ2ydzKgzd2E+A4nXFgkNwFIaE57jsdgBKHckiqJ+N1wL2PH+
CoFeDyL5VH72iKAIQ2+bDoykkaZWqY5Zm6tvA85vQ9I5DH9J3SE69dUR27qWunmZ
GhnIxCUVXhy1skNcZhgH2x+9reOv7XGkk8tTHntVGqYfBgnawZfkdmxMzjEJMokV
ZKW9zT4DFcQaQQImkaOUh16O6vpraQPTMFN1D3wCOsilGKXfhSIuFQqEU4tp6TMj
QVcE/8NlROPrnX8NfSMolGKtNTsFMtowZ91OQW4xPi2L7uHbZXnKh4E4VcuF9SVI
opxI7tUcq3LX1y3Cv5U1aYfIv+/LaErJO0oj6nMQyyMSgcgiC7kh+BJhYySCgJ7E
Iq2xmz39uycTzw3Sid0juhEeyhIBrGKn6epiraoXyDU+ZowmX71ns2Z9cNhQNwS7
2ohV3zBH0Qp7F3zrhuuGX6iSW2psVtc8PMPV43rRrbwV03YFYfvUBoHn+wkh9F19
T522bfylP5xMNA3SKMhohu+dnoKjD/+H/hHDrQ5vJbzOrU/0RStA5fTxeF/0Blm9
aEl/3oSnnNJYRlJwl8rmrJOs7bY9Je0Q7QkdVHUnbvCOk08Qs5pRD+7iw1rr30cw
MG0DAmkwhDdFeHNyBKVBjvVluVvEJAU0s72HYXpS9a5XQJ5hHM8mWgVVJ8IraKHX
++EuWZUoo82EOiGb0GPSOiT0N7gP8gNuSrwg/xzG3BKxnSnxgup9TnjgLUv2uH7Q
9H8nZHKITpDyUNBAZiL/Did7D/6h00oGIkLK3FSgZNVHJJ+YtpIZUWq1DbXSPmMm
KI5xlSR41XUO6I0NspwOOe90JHFcV0H3MzFJKnWdH6RPkZJK2N5eQLPEUWq/Rgpx
gBi0BO2rLvgqIzugopb6YMu5R8QvNBG79BSOwyKyIgrAlqSiL970UykME17vme6a
BA+TIdz2+e1Tgl4H1wEhikKtzckYGb44G71V9TRvpVhaOkrLz5hpjcQKILEt8APr
hPL/nyWkk3viYTEtt15yjvbgSRiMjpsCroCzepi00KJeJGd4tj4uyGNyZdNMa2Am
LiLynmTx79nY6KU7EfpdNRK3WcAXvEt9aEMpNPH2ZpHiY61lHBgRaUNS5ZI6H2Dh
7oTiFHFX8UR8e3TUgjwv15Yb5QuV+yLbrl2sCI8OgeUJB5sfUli/JwaelLevwBBZ
p9VkPDDzVypksxgCg/TJ5bo0xzEf6YOagU7mmllviERM77ydwMYL/yL0sFBtl9IQ
g2LFl+jzxYrNiSK7k4eFVF5AZwz4HsbQHyCO11fz7qcFCh7HP0xoa8FyKw74DYKM
1Au7443qdltWvmoySdT5BFEMEs6IjUeuX/9NLc6jO970lthus6lwN6Nh6jSx2V5g
eGviWkYzyCFO3kYglUdt7bpZxXGqU3d3+7mVQzDue75ZAQSnJF4Nc4gyuZEbDtW3
ZF01jzd78vFkxk76gaMmwG/7et1SuTwrf/1Blm8FGYYB3ns6D+uo7zJOT3ho1uBZ
+xFWbUbOb4SvET5j14MaeInAU4zlz9RlbhVNwYPSiT1whLLdQhtfjhv2iDAuOPgo
66HwATtpkXH5R6UP8i/OIzqKvnii1NB0rvQ8Teahkwd1bPEz0FEBqoSQJKNF3HH5
TcKSZLDDsMxr00S72x5ALbKOLA4t2x5mwOlo5S/+V09PPCVhGCUxDfPHlfNLa7zk
yPa2WjN0+Q93EADg0lMK6opQkj8yvPPbdC3b5QP3YkWWiEwH23Hp1He4HMZ5k/dy
E7Dlma2aLAEPBxTASc1QV08Bt6cwhWsDW4dzQHY75EMrO9X1yO0ZnmfkCMshycni
sbuSwUbTb1JVaSYFvDLsi7q5Sl6ywcDjId6vgFbdFlojbG1iS71XwDCJQGIsbOme
DJIVGlGIhR/cisgVh5aefeW1oxvoNtSjwSd+5e3wb1q/0dyt1biSI2sTCq7E557w
5kb9NziDE7Krsjj8rmJr5CjppBTH98dAr+8uSaqGFN+hWdSsmkM1ATS5nlCem3xu
794Tv9Hs6maoIptUqP7G8YUYA7dwRUG+IhuMMoEIshe3wNvWbnOhBkwRv6L/qP1q
yhXfWgFM2we+tPP3GbXRqc+8x3Ntzx611QPv0xb6TnHY2cOFIyIk+a975nDegJBn
9JCcZV5ZJoWqzwW4wY3mnFeaDkxdpuMXMo1l2FPbxUiH/AvXHZ4ZGesB8ylavEW9
Eb5Ef1Q+synFgTDfAtPrJmkJYHpEh/a2PRRq4lmwYTTYL2BAOeZObWahqyGwnH7S
r+t73N65ShnLj1gWTusIb/2997y6KGWK3vwpCl/i2IdZvhoWF2oYBbkPJA6rODuQ
p6xEmZdpW7oJ21w2SAvaX4kZHTPobx3qpPVmNJag7nRQYK2TyEtM+h1z7FoCoZ+Z
LTNe5SgJlh6hEuMDchv7yDmHSwJZzWQtNQ3YMRIZ7FwatVFto5KNfczybzsW79tL
NPKlBhneNcZvqu5MxiDuwqRyZep+t87swl72vtOtxcVtJ9nuyr3u0Wb8WaV5JcZU
Fc60GCK+NVHcOpFVr4LCnQ0GMXGPV124jvBiO+TVzMdIg/iC5ikF1N6QFQepa9fm
nPQ3g+2CsPpkPB13IJ4W1/WpuwwygUCaj57u9Z2b92UsZ/tBI4CZlgqO0OCH3nhI
3RWszCj4p6MGE7gXSmASqccl8QbY8/7AGr3TB1HXXzgVZMkH0IBdJKwn9Cwwdeku
WTISJqBTQUF9oRPAYQy5/jC7GcfPHzhHPppTkiNuK1cle+/1BjJxp1y8xqGP3eXl
EBzP0UDMFWvjT2hMWKxfN/jeQPGN9RO72xCMxtiotAGHQRKhaANDnAVOqg4D3r0l
ZfZhBH309ecrTgMTffpBoX/0WJpwfcETtjbXHT/gnoStQFbS41kMZQ06LTSNq8fs
rSl6sYKF5Rz4m5Pqa0HBYTQipt4/j3K/VIOf0BgJAlQwALyFb3f8oGLDnL3d0hw9
f2D6An8p6Jg3gb2yHCu4axDcM1ax7wZsQo1mXySikb+ifRA+MVRKgJxt111a/9HA
cfr4g0lUhqFMCPRi1waR/1BHZ6PdzDVLuTCFwoyda2r/SuruE+jl6PIBI43EqMTI
GhhSkt5gAQ9cE6WHBKlu16D07wV8yCysLgpxPSjPJQIr0X5eIkwMTX4gPoEbqYxI
VMiLOS93grGdtt0oNW7zuHMsnZgJXiXRfPxWc3zJYPEwdkbNXl46WGuokeamjegv
zBNf1UXdddd3LyX85Ny0wIHyGjMcmenxG2J8GWwUH9AZUk5/If0/VnsYhIwj843+
PTc7N6H3KIrP0WMN5pjjsTWzyyJEM5eobXMWZ5sV67AzwcwihX/pL+5x2IUc5RYj
ALpwcdmIchWhZw//g9avTe8KSqbzrVtgAvs9xchafuONtQgp0a+8CKQ07owCCpTO
xgbrHHf8z2oyZYRSmpgtlux5d7ncTQ7dOGx6FXU0D7VNuSCa6Ac0AT03cdbYgs+M
TY4Rl2Ap6y5ZKH/UWMaJd0FqHCNvVAGkF/+mgZCENYXBTjCHaBWCUCovArYkhUv+
2REjdAKVjbUYYz8BihclAKl4nZwGjb5Xotup0L9mHx1rKh+55cWn86uYn+2v+K+g
FKCdxt9Yq7K7p0n8+pj19SBBJNRoeXQRUh8ljUYg//vC3Uf/2WmoAb2BiEGncj4Z
hPtgEjwGHbFte1wJKuhOYMqjyPSE/P3B+zo1qW62/gw71QzdPT7P4MKfN5+D42j1
bm3/QSi3WWnxFxo72i16GtkaQrxwPXCM42acrGi5gstS6iPZoMQKVoUAszZ00ECc
2E7a7gaHy2X9h6dkTTAMMOSsGIpftjkifVdxzuabbmjJIFOvfKMeGEGTYbQtjkeu
qZBrftlwMIm/Lw48XSxdi6FcbTBVPz+a+ngpBJcVBwNezRkPUewDRmpAqFJEjIPy
00g9JGRnlkFIk2zxNT1FkIxHC5onbP26FJNnxWdgE53mxJM+UM+yAyBQKA78gi3J
dMq2BVmuDXoTultA4fe1ZIEK2y9bndqu97MtxPVbp2f8tsXydkei/u7EQMUifDDu
ZeG7rQklo5MIVlmC4QK4woCJWE/ShiTMP8/GABcHGAjgyfCCaM80Yi7rXwmdEFSJ
AkJ5j5gKpKvwJTRjZkylta0C4oRWQKUGZ0n5+Q7jIFAiavaqghYogSqvNbpQ4leI
CCfLWA3pIY2X3I+gLd/oNKe8vYEkktBDFcyhgspXXpaoNTxCNMRLp6AKz0NaQmPv
IIeH3U59cM08mkVZ/QVXpFLXZJtVEzBrQk5MHMNBT4baaDCPTKveICiEJ5OOv/Mh
iqRTZHnJ1OhHrWTmMhOFIlJtOpn0scPRm6gxbbx9EB+OWAmaNqQFT5WtLfPq3DMD
obwbAS4xmxocL0gBNWMrazdB7iEYfTnH042V8MVxA+rld2NUvhm84QmJqUZFtn4y
GKLgxAmZqtQp7UM/GOQHjjNhGJ80lZU1G60IUeUVW7EUTx6uObz0uN6H0vp53nmU
18c3REbwogtGFiRYJnIChmNA+yodgztiQdeNMM0Pmk1QwXP57d+1HPIiWUmO4rls
U9k0rZREOJ/ldXFyWO/YPQ7EZ9VSGD7L+S3z2YYSRYy8WNrHT26eJBA6wZoZ0Vke
UcH3MvXPOU7WSBIjZNMIBieXbwN4q16KhqOF02Qdflv5xy9YvkPHU38j8llBYmjK
2kgy2nitOasEo24HoVZbLfvnyziauSXR3YtCo0ndKIcXKgSRiz2stvtdPELggzQh
bX/33VoHmDbspI4HVSpUs9etmt7sMqaBHPX55JN4PewFXfhGfvx3LNTHMXWwGiVF
WM0RGf8cRu8tHOpvprxBp/43yTUFRnkcjKMBaB/gqbraJItS70C5QI7QIAFbzWq7
K61Eo8Zc2d9TCgPFB7Jm1nkNtsJe/xbzCkZgCgfSrtFACzqrcRBvFIAN+t8KCj+w
HTcL1Na8x7nwR5IvfLjj292MEXt3T1lF0HVdb0pcBifjDaDY9PIOKf7XhvhYzs8F
CKTU3uXtuXm2QoMMOhGbxDwPFcHOLgPbAAxd4KjWE1eIwQGdm18aMwL93h29LIlL
+VTXAvlB49I8ofxyO++7xDKY9QXi+xKK4Z+dvMGRCyEOhczbOg3V9GXK7Z2KUgiA
Dc8qMUiQI1L2DFDElddIGHtZtzD7tn2OpyBugIxAxZmK0Ku0o/2kR7MZ7uxleZKZ
psyDZqtS+0trrHwnV0ZqlkaJeL11ujVKZBvy14QkIUA1TNgleOvzuVKLAqdjs7kL
8NKdnQrNSIaDhY6WMUXD4b/C7Lwa1v5In77CmPrAzE5U2ja2J5Za5W8KqIbHYA3+
TgrxR4zlWRZ5oCgZgf9YBMPvFrJBBBMPySI6MkBnCVXQp6LQ7nNpAJcZJ/t9URCY
UMwkqEBKNhfkyXyZyx0sjoNNc4az6wgYProe15AohKd5Qxxlv7FPD0G0epWAvyER
KbPlIFU/EhfbKBFxsGtO3eAWzMaKHCzoXLE2JR67r2KCZnipYvvOiY06s6A/llVR
qWDBvkSGTpbX+4uhz5/UQRtwnPs2EI1mjuBASlAjrXilTcSXLDeaNNo/80BijqT0
dTl+a03/Sd4FchoAxSHHtZ5732PmaPWLdIluAWdTM5/kaOga8ufUvtfZn8tXCPT5
YcAjcXKFxtx937DJY74JqL74GZ6XUr8LYFxRWlC6DiNd9nXUmIFv//iEz6PYW67X
3BX4irB/xzOIKdenNmSZQ/m/jfYmg5exN2571hQZN3khdTnzfnSqVf8NTgowZ0KN
zugt/9zLcH/NxHBnTO7EsojcUMf3LrOe0hvvfk3Vd9aJ1ssL1SMfgTSKrFh4qwfQ
0JjjsKByJ4YfYATIsghDElABmTplHG+03sN7ZO+7FKbBiguYE01FnlkV6YeEm/Yv
Yf9x/MxHgG8B0eYT+MXgO3Nr/o77UwXscSjTl+EiC6eOuSoqiHK72XSrH2960f2x
sl+KaOziYnw8XGH4713ci5CLoRc1iQwHtcYoFzewmgfk64qVLhA40qvaYi0EP9h3
VerVSlWIRo8pEUNNm5nbx5tdQ75eDgbMnLGt+ORz80yVq7gOog0I/o/oiM4CgsK0
lrPJqQK6f4K2Z1RsOKsGhBymXRwh/Tx4MqWaCjgfMACBtudKWtvwmEHeR5ml2ohA
M+05wn1kd6nJH6XfJRO8ijeIdeAQn6C+3M8QSlznqsmNrTq8OWpHRwZZzrTom0ut
/NOSYjYNXUQDWMG6QI/ATjaa4Y3O61BEC8IuQq/nhy+8eWhkG75kDc1S1AiiSjen
RYwrbQnlfSErNKkkL/5MmdOe3ckQ7XUO3gfVSyyP+FyT9rjLdH2ZDf46i3F/PD3Y
jy72x/xMYEcCC+kxd9QCUfOCk8HaWz0Cs5ae/7xPDkI5cnnrmlLPwmZqY8HKXPc+
l9Dnf2rOeEo1m1DaNf8K0IC058uYkH2aGjU+k7tLoZJk/COiTFPx8dI6jbAzNPeA
x45Uo9lpIeCFmM3Tt+yr0Yougu2bdqRU6WQl3uDdHrXkXthAGKKsDuOhdDmAkNVP
pC/bAvtk8iJLXUrOW1MrI/xcMYVy3rKqS2BJBLzPqDmaiphp7L49ugJSVzCvPcmm
aQSMY542MrroR0zFe0UCmTpa9D+6E8dfpjkT5RP7m7agUV33YDdue9KLx9nagNAi
7/uDLcN/TOSFOMoHveUE8Iumdn/+3Ig1ztxdXUssyjtff9XMgzpXQTEoi7fi/3EW
RmKjApg5RbQkKOpan0o2XO317DF3MNPjbqJx9H57sxLV1icXO0QpU7xFtpfxkPWq
+1EwF/DLN5nLUZK4K8gvWNBB6Sn94m3OIc2NQQDYhfcrZ+cPKUxBC4xqmk7QCi4O
XzpMLQ6QPYWgdL2r1vBFZLglxWboNA6tvRB5AmayYs+I9cBbbDvFQlPa9iNLKMYl
VI7LNYTQtytFE9OBd4InP6CoNurXB5dkn4bJ0YQq0MNX0lZE6y2gUzk/Bvda7xvL
Z9eIJa0PROcPUuN9tN6ijteJ0eO7TkEd0BPDEwfD9k+Yd84UsNzujhueMtPRIe/A
FcyGObzDCxhiUT/ygFjdvtqcQvJg8/BNPEwovV5ibn3sCOqIWIafE26TARtNnyif
LNfmLzm8yHFmOvs0c6+8K6STtsB4iv5FRqUc+tj7ctjBG9VAaQcd/Oo6eaLPez5B
78qUWly+GN2s1vPFUu8RCkKtG1mZd9i7znAk/eCmzcYPcsyichXYuBEUIgM1OH8U
K4EdfTeXxAHPesUsxQWI0pIw9y3ePiNfI0oIg+aZDL/tYzjqRqeQW8gjdNCtIGap
YIiPYZ9Ml+EnNMgPeY4aNLjatkCuQqVl0N6GPuQZ7hvB/fXA9mT8O5V5wpXbCAXm
Fl7NAY9S+EgDD6kO2V27gmc13/ZwsKBa88SXPpnbhKUVB9mTq03Sa1MvAXYQUcJw
nViywVLF3LvjZo7hU2kpLeT6nFGGKYXHGf8JXVxFKwcb9ITIVkGwV5HxLVzwfxIq
nY3aVc60kzjtR9W+lkTEZPa4Pj+LmIuLZPQQzWANIWRfcuyMKr1d+LXX3nTWd59u
34lRDmKHCB43Ns4em1s85wJJt4F4Yxo3ew1SfRjlogREDNYJ8PaOL6h246wMFKPB
L1XACFvHL7cWnvKqby7umCY5nf7kumr+Z9jEZb1pi6dhRVUHGmx6z+AwIHqJVHOI
b2owLCMbpKU1WLm0wsRdQ8ihhpzxU/hPgsvLVtb4zxczFiCdvotLjFnbjX4bfvCE
mRVWCK74czVexZqE7b/6d0V3FGMf4SFj9LwoBWe8YxpbOlA9HNh73t5/FNnugmMp
wOehMPh6RgIkyE3SS1RiOeeA2EqqU3HOlyBIzA0lJoYkqUGbFeaMH4gnn6I5zxwN
6IosJjuXEoefgfjseAScjQ/jPuB8YdCu+HZKcrzE8lHJQrVBRBnpgkuIcrwZUOR1
KUwlESYhYSfI/KIylBnTi6f5qQ9Sr7TkBllT/FFJXsNwtJKp7WOhhguhSpN2iurg
Hvqj6Aelc9S9suyO2d9U7EqRLuko+fOMb+buMy4QnLcEQftrx+qxw7gE9h7XyS09
KhHTv2Hsx1WXvGwPu814LN2XhHZg64Y0jD91S9kAgIhX26EcMqoOSuasAd+or+vc
mBpR75lFBvjlzr3uiz+KJyg0HGJlfOoqJqyWxntrrvnKBWzw2lh2acPg6MHE1DzF
AVuDmMmeB2WzpZUiHLvN8HDON+EEOwJLDwqj8twAnHYAN3MfNxKdLC7e0uekj9W0
DkLWmjUj1W2Q86GqRlr3+svZ6S98zriKJOgI6U0C/4b1xWb72uaq1QyFNS9x9DlF
YxvPy5J7vTVipTOQD0d/zAR5EoRJbVV9F2zMrgqJIv8dzf5s9VXAOAkUeT4VB+fO
2fWO9hcgQAT2tR5H4eHdYyKar5F473IlOb0ITKjFQxxOhPM7xou19XdyykeID/4L
TDdEGxC2JegzMLFMXRq1W4oXAijd/ZAlvs3j1tihZHZEcyZ6pQ+LzLy8HTdDOLe+
tVEEL7J356sUm3qZn49eOMiZpbAdByJLHvBlwx3uGBEz9G94o1M8sFtcPSzd71bD
zAT12W5cpYfxIUgus6xhoEqbz7OKuIGMF6yGXkNkU+oZxy1JZ2bVxUtFJKtfw3ly
nTfEneC+2FKY2LPw9/qA3FHKworRZq6A/jwMh7zpFGe40wAu3DW6NaRIibliSLcO
VipDq55l++6yFEPmAoIG6xlsNHGY0OxtvSIHnNuGB+epiP9L/Yz0X1C0JLQbH+CH
AZ89glnqFGe2xOb8nTvwRTpNIRsn2Zgc66VxpnCUOjQ5QAu2yu+4AGvfDQ500++5
aOjiuMke9PQFty1ViLalRXUXOffgAoYmZg1uqpEs1XVr8nmDJN5/pzRmmtM/e0N7
AAVYdCY4cb1SJL3J+oD2h6H7xTp03YN8BFdbChLN08rkrgax/7ya8/ln5UbQXhkA
d+ajFsF7Pozs9PVKdGT4C0c/bOrbywgLjH3YdnHLpDItpIp8nrk6Fg740ZAk8MsQ
TQO2lcc2WtuznOlkv1+u33u5Xuxz5tkzGBxMoBYe70WSXpM56LyO1lIY9HLPohXQ
g2OSC1KOmLS+wcWrpEg+uBfkWUWCK6r3amBA0al5TxLtWywKG+mRmxGgAHIokPSp
rX1xw1KBiGYEtFD4jzqYPa6gd2CztQlnQ5pu8Z0aE9DvIQhZ73ChOxlKnwLuM2Ts
+0YXM/tJeJlDj2r6d4wUmXBtPs8xukWYeC/1EFCj8xU8BIIHR3I9PLVWLGXzHGll
YwwBjjbORYSfwKwmPulu+kWiJwurOzf0G7biXgdcI1xp8E4GHKlxzE0KvazdKzTN
y04CYR13muHh2mm2qBMQskFS4Osm2JKpNIDTNmwbt12ZAd6qkbZ1ds8RdHjNTO3A
CpgJ2X73enQSXX2dEU63Y5X+NTE1/kjoa4XQ/DbvXd7TZOnHuugnwvC7bULvJdEq
ZLLkDMLK6LJpcSsG/YZwe3ozF8+NwJW3gpbZE1/2/hoCA3XOs/o4FF6wMcqIcqX5
oTERjeAsDzebuDolkTiI4gTZikEX1916NY1O3RdR2AZTPDpBFZWe2H36P/Jsz+na
s4kI8jcNUEZ7QfLt6ulicY38VDOJS4FV9zsuiuA51R3cMOGD9fHaBh9ZWK6pMC3z
5GTQvnLLeqBi4cLlohRU073/BVU6tmjHQytfY3VwVZl6/eIDp5gnKL02A1AGDFWz
K4qPf6bwgVVmp+CB6GeIMhpoJDpv3kaW4DLcQLLsPTTvaBIbfEOaUos+dJouXCJx
ema7UWxOY+1ZwDpxCaqPOO1Jze8p7d2uvt8uMRG6p3n0vsRgNKGngi61UrlZEIpa
YjxaG8EefaRarq7aZat/UQvfFHkm5YeUgeB4XJNObFE5ByzmsTAsW9FRIlmdQclS
qvyxtKM8h7ZYiewxZXcHN73fdKkUrkPil1yjU6V45IO3dJXrfiZGlOIuNQf5l9IM
Hv8ry2sUPhxQI1h0+sc8cYJAWtwuE1xubTYYTPcHZl2704Xd993QGjFnboodlP4b
M0nvi7tklB9UFQ6WTGMkFbjKC429IibrlwsehOVgTS14jP9elN6EPxTv3MFV6WO3
cne65tcyWcIqA/OfmENrL9hGP5PaPgRqFiwxTWrGJy/QRTX/JvLB/7D7Zm8WvjaQ
FKhDKq7rg+H+yNZqhYih3e9rc95+I/mMTvsJAdDZ0ycGlsmpd+Q7QrdlQ/zQu6DP
pVU1wpvXyC/+7TYYF4RDuracFYCY+iBhce8+3D3sE8YJDLpNjHYID8mWOuPfqA2w
z6mytkhSFVTS5aRsSOQ9iL0Kv4VdIDfbVQmAt10p8vGovDxIwQIdzTFxCk7kON2E
Q4Q08/D8UnYOxAj8zZ8BPYdCWRvXVSq/Xvj2SdiMRSjovxq+eOpnC0/AKmLadNUW
urZStLtEn+AHfMzHbmM+G4ae/sfL8E20thtigU2p7C/NUJD5lAZf8jxnbhjvwuAE
j7J5891JDYDoWKpzfkrtj7rRlEO1KUZzbOHc2RLpSJlbn/Ia2wGqKAo8MtFBYB8S
xaIqxd1LI5yI1GAmeghQM8/mi1hy2MfZZxePTO2PXy876mrt9YsoGBPkYgnmtzzZ
Jy/O0WbGp9EJ3Uag30eVosjsLjPyV+/yWND/yi3srn0xPSDGMFgVUR6IVZJ2vXlX
gf+WwfOUXc8pb04vR3gvaVt2CCEbJa3L1YQvKOKCLsIbjpmWCjPip6Gey64EOxf/
DRdiT+JgwKCpn5WA0gEWKTzNnTf9gAj+MDF5fCG+nGtFQxHrjDUzWIU/mfsVpBVv
kl1doqn2bcCcuSuGcx5ckFCOr3tTSN5BX11OujyeoCveRTbwaiFEh3Db4PhMn9+g
WuzuRkrdwm1APCAIgxSoTq/3Y4fK2ECftb+CV0AYwEm35fISBQLC7XQ8zcZNiSV1
OWXbvGmEuPXSs5XT6JH5HdnsrUIXUiPydAuzj43js4OCVdIR9a3+7xDZb404oAlr
RGJIJenSFuKUiE4SC13i4+CH8mpR1VSFMY1hne5dvnr0wwI5Si6k2iopaMDhZeX2
GXpk+VRLc70tqBAHQ89S9McUSNrRjS6OlcUDnL5dlW+KlXTxeLU0sY8x1+9D79+9
+rl1ZfU+Z6njtiNgiT4rbbv1SqSvD9VFNeMUSZFWLoaNE8Knkcw6mOVg6P+Twjxj
hfdzEjNVNt02+JDV2uGmbYn6KuKLnBReaX9Ywbx9GdTWGqTnzDnBrU4AWVVehczH
JBEcg4K5oOETntl8mg1avR/zETnwH871ejrhQ98vEjHe8fGTe9tzJ6DGrhvMBVMy
2ECDuMPQANfdqavkpMvff6NGqlRh0cgu1AJ+/swn7T1w6IQFZZbzKQ8Qmxu9FRsM
jNXLm33X77zHjT+sMal6hpQF2//Ct69ILbaRS/aak0bSIsV+YUkgTIlCZ+T6KryS
A9ljimWp0k7f74AW3PITBmf6xB7vKsHuG3WObC/zlxsapyB8h7KcQVHzpKvxlP+3
jnPGY0hkS+Xxl/cSgpdjH/HPWw535Rg4GABq/UEKpOGJrNieebaKNjq1YvSoC2l7
giUjBdtGri+USubwKKw0UZDN51p+/ZFPHNalAWMOuamORlML9URexAJ5mxoSS9kI
QiFhULDciUYjATvFsgXlU1Vxh99/Gch1nyX2Q606R3ogG1yixYhegmIGHEy0xCwf
XH2G2xZ//MruCcxWKmHSgvm7760NK2SQEG04djJ3dsvx6JXz7YjRRM9dBTiNDW7t
IEfF2/iwor8Ze0etntYKOTYRaqGySL6fRE2vZP7B2RcXiB52WcKDWmF3u9xbjpQo
IDPT+82aEzxWBndAnZFz9N7QtSAqpfRjkJZrsNhtt9tg9TwnMc79IqdyUiUVXzSw
+fmLaf7iVrEYrpHPRUqa1RKu1yhjaTNkjZ+zPy0GX8lko4nmqeqRb/bApB+bRVIL
MQKit0kB6gsQEf43I0rLJOCfugQ13E6zCRmHaXZUwTWUqaHP9EG4K0hCAReqm+K+
EuAUs+ysi6CpceJmMcAyKvTno9J8ixb+K0XvZHE8YUwxrPgiQk+jlNFlJMzVeKiZ
yLZXIdI+zZPcMKDoa5ZTgqnbkkI7hmXp0l9NbB9zi8QiROft+Yd7BWzD6H3/fkCc
IWg6zPGZTOdUsosxb70ANnl5mu9cYsRnWUq74E6/ePGag+5Wf0j75v80YSIqOwla
AtmpKlHTsUjCnUC+YbUMJtE5ZVIVzFAFBYFfvWey9dEqSE6WgvL5IqT0le+d8Gn7
wctpixCK2kSc2LtRVZIPZl+gQfNZ7RXtxzxTNxqpvxSVjjR9cv01nYuFtCQrjOhe
ylks8/zYLV86WMdyyPQqh5UXLLOPZcgR0FjkxseRQvAsTGH0hsP8GgI9jekRHfBD
DIHxSuaZ/RxH2JtxILDnYhv59qOYcZHd9Q1XbtNeboIuWEG5MFInCg7wehveSVeh
UdYKMs+IqOOrsviJF+OdXC9wemEwXdQLCyqKVedc+yMvsgeDLLYGnfxrzMxbc7Rv
RJoLOGt5rCZ+ZA6ZTZqp0AfmWzGpM+HIjE8gc3rj8ZwA5J3yrQEtMIrmi5XkTzKi
e/7Gsk6nBJCGrJkjlN7yaQrYjOFKDoh5Jkgrh1vBQd6YuE2JZJutwavfBmtnEd0u
Tbv96VcCDXO8HfGdYwbZAtCC5KDuyWFNHZTR8GN0aULh1z/vPrhMETsLMDQlfAyT
qoGvRqtcyF6r5GXG183Dsol2oxmzVpF12r0E62S0aQz54LMJy9Rg8vWpxJZ3ScqC
I6jImrBuHApFHdplBalprtVqrVPz9NogPP1Cg6u4d0T0jJFuonGWehC+a/ldMaQI
12VpkmBSvnFiDIKTF5MEk/yEewCzdzVvZZC7H7JD1wY+QUVJmlwmEhEVUBdEeofs
Bm5S8Nk0CsVZzoOoFmj3TlAf2Pkz1Sx67HWaaOgEy3RO6IBhxbO4RYFr0CcHWqTk
SdcqnuzGw25hTN0V947s/GhxunCeOjvYo68KF9/I3MaXjgf2UXu2lhtYycA0LKX0
sm1dalJe4Tz1Fla1hSuRC0iQccC2Y6Y1CBdveWVare2w3qtoJ9GWxAvKiUbOfj53
Jor6dCsJT8KK3b7bKKRU8INKwcAG3MEec8y7DCK+8BMfvyJ1PwrKxA+g0R9+w1De
QsJHy0/V5KOH4IbCdjlnq+i+bZhw+8M/y2meJ5l9jWjYf4XVnm/iC1qKHoAdm5Xz
jKVWJRk1ZIib+2zh8FPyWpmuR63H5sefZfM91Vp4Yd3I1rozu1coPwZA1BDXOtFp
+vWXrja8HZY5eQ62M/G2fdwLuXcCWO52n59yzbBOB+F48z8YLVRzzEg5ZhsM3gRW
rQA+eLM1upeT8h4NNPYXpAd6RL2+gATP3UHzoEUMwjJIdSbyJzufx6qww2s5LFvX
umq7BBbYfom5a6vCP7ug4SSxkvp6Bzc4I545MTDbKil5cuwpusXc+h1Bhh7vcW7j
O346DyFVeYhJCtpn8KjrB7EA9mz0k25Ot8qEvk/DH6niQrV7AkaG3EmrwCHc0K8Z
kQgLKs2ftbnuB5KWnJ5g/2uj9oV3cEEm88En0ily9Hsg/jhLYGULnfSVXJaMspVB
yV5A08lA44xmuzcgXPZjhhPhFr+MJ1QSeFRv+XklJftyJQLh1EAoF94ge2MtQWlo
E3WNLpoYQiS9wWARu/blcAI0X5LStvdK93XAmwaK+7CeplSC+ZyZxGsQfv/LDwwx
FVmz5mX2mFX+aZ0DGF9UX00qwUszwD/xncDb0EN7CWpSg5C4+Yaz93HfMsQBMdKe
iZgTYGmnV//SDz+s+ZKdQNhoPQzSUTqhf40BcG8W+mut+X36lQEDnQGfOZDQ7Zxn
NAQS0FNHu/DjnPcIHNO5cKhUOO3RqcLGiY6dTXuvPUPxxMkP0ioVywFFXwEpOztd
PmtXDfYmBjlGokyCgHNluiUboTocCLLwiHl8bdEKiNGRz4Caw8CgH3/7vgYJ9iKr
3aSAuu64FAOi32fb9hKRreZCF5c2lXncdjR5YPZeCNxjDqjy3hL5PaEzGnafAxHW
owdGpAx1LcOtpnopK8zbHpkXFUJsC2PAvDnhxx+sDCbCGG5Rmp5xmPyZo7QQR7ig
SXg4cmyA7uaPEdCMqRKr/kh0ySssX5g99CQcLObebGpqcNnjjv4fVYQqwNaPFCe5
EUiw8sz2/Z63FX6HDPYMZa6ZqbjuS9le0b897eiF8XN1EEsaj4HkmVOy2DYvmT0U
TzJNblJudVKjWCuL1zkZmyC+EbvtdH+ecsp5TWhmWkebuduEHN+JrtkCmM6jFQcG
3o6lXAh5gKkLDK0wqJVDfAVJC863VcEoFJB9VHq5qgQUTjSBnqYDzgS3xbFbeqxL
BDlJRXh3JsY3VDjMlLVI6j71KKS5ERL5+zXyGGH9Lvsg1WXEz5dAmSZZQZhcAdRS
T1StyMxsvqKGvQw8tU75xgPFuLo1u3D7c3sCr7Bi3t3LTOClPo+q0B6tvv5TGbG3
SajS9sLh3mQ5teGdCSsjxhZMBpARkV44V1SM3szrZXH2xT0t3JGatvyM50haht8F
kq7KP77jOzAzuoZjbriiFhxJqNpHOmnbpzEuUfq/yigfT71NXCJCNnjRqqpJTsxl
ImnLbfmhoFe2AjPW7kD+cuXeUZwWKc8rPm/ZbXR3OQzrDvWRAwQRExVhxvyvqvUO
ZTufbfM04oB3lKUcuXk8VrR036uSzRxBN5UU6b4c4jFopA0/9EBIWWzRylkm7VsS
02AJsHDvZeam5rB8nRnVorR+HCB7ADnq/MOmhNfSRlr2BwVp1fNff+S9bJ2x0sXu
GiX64D1zwB0xgKZi+FFgbTPMilwpwPdcctNwMFI7YA0lPjmeTPGozBbG+IIwODQf
JngMS/2kgyH0k2RF8DML3+MtuW9Pp3TBeTEToRCofH1h525waAU8b/o1LisBM8Dc
BAnkAe4YESwe6CPJKTAY6bkRSzutdXK+TBI3YAVEpOeA40ahDkwFXMbyA5d4BTpK
4+izj49mh8+AtbY0jsxSq4nM/cS7YmUJh5w+MYnKCPaQcMt5lvczJ8lPv59DvNeZ
YHoGNBze0W6psI69TFZdEKBQ8Plz7kQkvA7Rm1badBDX/0QqfTyPfrOeX46llrvS
tzdzLco47BnQbWixfYkbeEqWpuEvFMXdUMJ6c5tyjThmcc9uPJWcL/0ORcH78Ypz
W3XLpBsXiCMm6DZyS6ytxxtp9rnsspBcjk8t1MLylnoUJVOJ9mdlMH9kBZ+edAfu
ClScgKuxXdMWwVVUshgB2JTJAVQFuFKDqjlBgSAWSVcCFftYA/ReTOXz8oN+UUhl
/3lZZ0RWgbVIFHhUGzpzN2l6V7n4deY0MQqz7FUsNEESvTu51LKgBv/vMKJcFgJN
QbhBGjY2OLL8dU+U/xckW13knzM7C94QU56/XE8ntTyxkD4S8srqVRCxNmG4mWWw
DZM49ytpN/rc+J3jLCgTE+hKwP6HUgJ7WBj61aaSsDcCZB56jL4AA5NgBf1b5esm
QhDuiUHFpJ81f6l8kkp59ClC0i7i+4myfcyGRObI+DZ7DSck52gyo6ZYcrVWOk8F
AwF4sBK//lH7xv8xY02YTq2acy0j/38j3WglkwJbAOBC4r5rW3n94sWwT8g55aVl
J5uAvituz5sY6NZe/jEgbIDEpUnRixJXIffsN32+kRNztw1R0uYyVCyXGzQGvrKk
oXyQ6ruNDnmL8/rKyXMOjpfbK80yKGNTSKTf/2fUjvUTmNdgW3KhbObSw4iGPh6x
Clh0nsgGIQa4i+u4aNFCh5EYe+9pDcriQVA77N+eX85f3Raf6ogIcE9nmc4qVPS+
nD4rwJJKrNJHpOmodJZ3kuZXdZg4tcJT/WcFxPhciy0mW8mk5+yicfqlBBe1rn6j
mC75y+R0F9OOAFmlWbHCiSyQT+ID4XdT2m/4fLpsS5CwqRnKd427YgQZyKpgLrAi
eGymnAGHtNH8owb8KTxVzsDbTQ4/G4r5R7C0+ZF2FpJePlBnH0fw6GF2H1Bk6nBl
7Z8++21GJGy9lp6ed44yDcIdK1m91kfmQlwsyaE2lzeyWD0QPdMZAEeCFMSO2w/0
6Ojg6vgT5xaCVN8Tp6e1CQ8QtiPoqtKI9dCq5QIraQirlA/ENSVyebriA8oq3SfC
isVi5gZaa+K1aalREUGcpclqzSxP2NdbqdLDWw4o07ZE4DG5LnYZMga4cdFJXWsU
YDV4uuRDt/c7Up6cH/pihJBQ1FvrgAdQj3lxVJaEarZrScSdbF/ELs/7/nJQHf/e
VqvGE0+FVCohjEv1ghpbdVqz+ZLcLoM3CzSNvBJUorsUSFFSJcF/dlxWDmjj9+I2
NuRa8e7CBYgwVKPe9utJB/DgtqfEb49au+MVURAzh03I/+W6Ilhfd6i/zgnbebZ5
6kxSoUQdc8W1GDWmR98ZblLOZZ+0DB8DiFGEKzsO1u07zNEV9uW72rE1BHVMM/IM
k4yx7JXfTDh88fETHpEZNrA5IxNB8LNFuilAOJwveQfR171MWot9cYMdH1rH1PYb
09e+Gx3vw0goyxoEnmrVu+yGXDSnXUuVfR2pKWThiMiwpRGE3XrT6J/lvSY1JVsy
KtN5EJeobBWQbiwgP/tZ52c4JQGz0RkageAMjsiflaD2cxHmZD51zIs3Ibg7kYAR
2r0GGQNZMGQTp1vY9AVHMj2Eg2uf9iNe2qqC9XjHc65ndOcd3DU0pIm8rC5YpftR
TsdQM5A9xbBgMd4YtVFsnPWlgPsjjXB6Mph2yu4tlJVRIyy+J72orGVgjXKv+Au3
hOTEjvsMW6tSpj++aGIt5cID6tguzRALe4UbzB2G+8+IGujvxvYYuTJ7BJkDlsQ5
TI/3zz2rXyC/1+aYPoznnnsMUdwKEcUUMDOWGxWsZ92i9VQ5+QcFAAUCXPCKU3rS
0EBMTB2HEeddqZWSjwcwS3GrM7+drlD5HHptQaPvfleQGIoJpYiB1USbJp3GULa5
EI2C37CCBSVsTjipBibMNfx/j/z3pjzHhgdO5Krxbxv4nHS/uS1kGA71l7RHVaV4
YQX9PagEHYZjEFgvswDtlDesrwLzxLAiXvHPgoYRTbDCDzapsvfFQrlyGWSGePB3
HK4GyBrpZL1/S1X989AynUwbOrCWBaetIzjERYY70U7KXCg9s/RnGY/32tyaSKYU
/EkdDRyTxPZ5TUb2EVhpQTyW5Nl5jySaEM4ZWxyh3IQkm+KeNslZnL4OlqgpOSZU
HFxxPdjsEPpZaXN4df9chjFmMlkvhhUt53OkG73IkIDhz4vUevBgdnevNoauHerH
PrGVft20s8NQSaIfdTDStvxTGTnKYvJ3ZBazfubLjRSCdCCKfiv6VKrcF2GPpFcn
G2UY0FmGPxmjqC/Z2D2Y59Hx42ae+71qGeuxUorakgxUQsAJRYFVwZCdsVFHPKOD
GudJp7tUnLz4K/5jh50ZIushxHu9+X+XA4n53L4Yvzdrfwz+SgKgZuPhFRf1euqw
5xeef+49DIlKiG1vbUcWeXygiAUChcttwHfQ7qw69/7MUqcSjKkntW6xgJC3QfK1
gfJG4wNtS5J9DbW/OGboN2fkT6d/CTtqbB2aTNJfnmMqsABU7NPxO3xwA/kxtnJO
U/WKItJabL0811R59cEpVUNrsGy/4QD6K/cn4vMu7X6OXBIw4LQignHNDz79PCY2
Uef6ZnGvjzeMUi/rSRYQPscCePGSTNQTci38tkk+ilJTyfbeorYUnxqF/h64OFwv
88yVERf5ItHtWsbaLULMk9gll/J2wAjhwgN4IorE7MVkqT2B/6zhQp3oF7MGBFXj
DHdI+ZsXIBENgo6VKOHZot31XuNSLMGrB4rMtYakCdKfg9l1JP1L4tsVoF2Q/Fdo
15Rz4Us1H00F2oOqqwXrUX5uKJd9SmJW/W9Mo6t1pcGo/2gRnl3TagQ3aaqCa1po
8mTVgVLx6X49C/XWJIbEQAI+uj96rAU8pUwbF98WoIVr6gymwg4rhP9sdPp+x7oz
cOFlvMYsuFguxIZUUbXkJofo/Wh6jWY8lKypV6xjB6cE73QE6/ZA6dupNSIHyu2h
D9oj1iPi4nat2MOenNpJuXmXP3LuBH5IsKDzfERRgk62T6SOD3efAeUafnyzjV/m
JJ2nEZrWYGvh5meHx/E3AS+RM0D5FIsNo9RHRPGH2dliitUPPM+olYcIibzaFQi/
5COpafPHQbHTyrdh3lpBiDg3aaVB77wb81ZOwyb4+o1tXS7DuKgXMn5XncWaZUs+
slJvzE5d1izHW+RUflY5lSJqohceNqYNO5vH75+7TUyUCHJLqb2Ue6mj1wPL5CO0
xiqtlitHR+B1Pl/sNwm16thq/AqjMV0ZxMwdK/SRUb4PJgheLsTtnVNkrvExxMxu
DzFFfJB57H+QSuawydCg4KZxgbHqT7hzBQXDgiI8/sIVme7qQKmE+lQeJ9ArtGe3
bn5ZyDcrv0ZqzASfQonn7kmap8FRb0tEvracgLCf2eJFaUAdfH4GSowDgrGdkBEO
dpsLFmTdEJufaW6MAD/AAMrNipL0jLDOMT/EXf5IuLlhadugcB1c0qqsURKqOKfk
bEorS+IRve4xV+98gUNHtsuLds6DxfBnSfSm9NFj4mZC22fbjSmQWmViqLJtoDP4
S1YVlsuMjEkMS1e425fkBwaGStX8bH2hBAanF7s5EKJy8CgsSGn/iKDVWHII13Bj
aj2B6jVLHJGTf7NwWLlzvdKuXbWfT5oQ+Xm8pjlE3KsO3xHgpwkq3gWyQDteDTqG
3zL9PLdlBBsGSZ+557TEUES7ET1ubCIOUQkVR/tJ75AaKHMl4K+fQ7CGb08uFQ1t
noLopvPsgE61RYThfl4LaiJSHjJVG1Aur7kMvECdrexxYMFzPO8vKaXGn2DAj3f5
Iemrt8ijdrP+eEUsRzvgQ00VL/yri54k5yWiBE+rn9+UlrqPEbgzjCKeFa8u3sw3
89ToLbYB0ygORG0CgYh3W9oKR0ZSHlV1U9vKuriMsQxQAXahfB9HVtZtYyhv5tyk
lxeSDvZZfy9tWLa9/J0Qhsj1LVh0YJIismCqxIiYrw8r5HiWoDYWlkGDr9Yn3ctQ
QGrpNqu/mc//dRezB7qm0MyXF1dhqZixY9lKlnvg1PcNJd4rJxeICN0YYf2psDyM
2VbpemN3Pu7RW9jQcnMOjCuE1WokmKxdM6rq2kRIrxEedGrtz0xmhOXfDgawisBz
PY8QDO+p/kpaCbJYTMWNYPrlm41GVMEd43THZbQIyJrNNEFVCZKpvfw3jVHwyfXt
u4AXuVyuHUPaZ8kJDw9+aSYGmAxAgJO/TTxmHlXzWeiUU8zNLz/aTlaEIjbmawhz
X9pPoxZ8F7j1MIbUu3wQbyWAO13erug6hvHkEZ1vp4JIQGjyxXpuj3kyax/7rQB1
5pczRe1Qfz9GVLla9xaqzmJNoZERGQBMM5SEhMh9CT3tAHt3KnnXCk200T4MhDbL
oiFCEtUnH6AKovZLHqGErsBrDfxcDP8GUazHjzpNIE/kjBKu/v6bho7GR3A1cVee
GhD7U3PF7B9ZtweUARhgophON9aQj6H5DBHXjyCtR/rLKzgaX0thoKXO7g6vo6Ol
PRnssJaK/QV+lBsBXtWyff+sLCoKFxDFHPPfwHvBWG+SVlzKVeEi+ATPzmetm5Bh
pB342deKJrZyKQ31McQEBfKBAiNdp0kpWHAqyoALKp3Ds+Bq55xxOmd+2dOYm/Wf
w39Pt0w1jmFGm2lkaDDxUs3jduB2vOwgHDJsRyr59aTVOE2LKWddzxSD57cSD2dy
0GWqCN3uewEmMVIzHNys9z3zjEz2D8laipSLcADgRnUVoKleZ1smNewpzGSQRSIm
6n6sdHYEG2N0iVKzdr+QC3nsmHo3SdFhfHzgsED7ZPM2PWEnn+UnKOHGXcRBIScV
Pk9ygprYeVXptsxfo6NxY1kc3lZiNlDFVRr5fCPFp53KcoZXgoOorCBc17lz0Lpr
9Vr2O25Mt5AH6EE/9vY4Q1F+xwKEEbT8TKUiyGS3x6kJw2UknLTSDGd6SaMyzAKK
1ESfiW+c4eN7X3o8SxdbabNr1c7Ql9GfpIW6KboAxRLqod2KlD3bed35H8szVJ5s
yZMB2Nd7UicP0q2K3CAGsabpxrJjtcLFohaFKj6sQ4Zn07iC3rI+YaPeiAptHP+4
M7OFZ/+O4e+tVJ7MWRuJ6Lf6YwLCsmRfwIKOCTiEJYMVxMnJzLUbUstFFJQBO2Bc
WWbAIPPhKa7WbzVEu5U5cfht4xaPJvItba6qXr2yBd5fZ0rVRQG7XEGQmlwnW89J
ajhGRShW08RIvk6+qzP5zkrNjTrBWs7ZszWsNrGNPR8LbdjyaUmnap2ovu5RLOea
/YIzx4S2MLG1dgdZALrsY8y7GM5dqGk5ew50yfDdHG/EXwSuW4YQNsmhVn6xL1cx
dGr0gYolXT9CNGET7/13z3Ujl/kCXA0tIGS2mmPdLGWX5bO0e5yS2jPudQk7zMXR
b8/Yx5mQxalmDxiYA5tZ+8aPN2yyOvITMYUPcqDKZBiwL4UgC5bpkB5HGxuTrsyk
B8+p8kGsme917t3WsvFfnpU4VOj3wywmbltLyDUSJcAcVequnKD71MmUbixv7XWu
/4VgwkpRiW2eTTh/VXnL5PxnlBBB4siahKsCTkv825mzPgddC1S+QVqjRVvJ8k8L
fuJESlD+RgXelfjhMrGQej0er0lPaguvJIG0h5Z0RZt0k5sXeJyP3UxeOgUlNOq6
xxOwRscZrepveWcjbqyMvE7T/GdolMzf9uuyJfY/4sQJRmOi4oTFDeySiWLIlEIJ
dqe7CcBIdcV57jrIc9la6GQVx50MDTmjW+UB9NaZ4LImxzGDTE9h085mp6hsMuLc
689OYwhRofN0piAIEPw1FY1oRPZSaa6XOnoE/16/+YoPQGsqB2uM+DfCZZABMIHU
BunNuNKjTq3tlCuUSoVnuKZKzlJraPldHpvDXI9mfk41gtLIAyqUqwZOuibeqXEg
RdtP5/R7DE0GZ374KkyCr54WB1l1El097tX/k5mQDoqK0ZNknOOi9uGiIjH66S+Y
Rc4uEhkp3QSyQl0ChYdiBR28eey0mgrSnXtzlj58eBFscmXjRmb7ur3/oPM2NtfS
Q0dD3yk4mfcm1d7AI4Af4oAm0Fgaum2eqMpvp+t2Vg/oVFULuvMFUU/YZMXyGFX/
9UikyTSjedkHt5Xx6qwnj/5ODJAU9pnaqbvxPqeJZy6hmvIrvGvQ01cLYR1FFIk8
puvbxgLI3u48Rm2A+xlT/69D0CEOAqSjl/kATCsClfTjAZJmR3I3QP4UIDbFpUfP
QH59vxc9xjLwTRkxZjqkXOH4VNOllPYMK8lfp1ftWyGAJZklVOjZX8BPd2ahkonh
jJST77Zsa3H3aC1F/CDLspK6PQODp7Pi6q3r7zeUgvpM+jCiQvDCsctNf+QZ4+CI
WrcyMVJKOu7/RG5OR/MESHqmUraDiRwHI2UBKzc0XDFd7UMkCakD/Zpply51Pe3N
F5hqCrc67bmi1xXsdTNbypc9/lnxIuA1HnrH2/bJpewg2nhxWKdv4i+6Tk/S7o3b
0r4TdeX+rDK7mD4LmHs/VwVt2JVp0rn1rHT+3okdRphE9vYyHcRojRSAjV0Ki+E7
IckINIL4SJIvd+dFGJ1TKbHrv50uKVqcdlKlQDd/Qa9M+bJxmumLaweB2HUaEqk3
cFm1IW/EIX7DBlJ1vmIU6ujM23T32qJNk4OKcvKuGvyaa0Sdobke+6VLh3tfTjJY
pyVwhOGTcLFqmVFndF31pM4oaIFxqPGdJgfQ6JnpKP41SdbLbH2YJsN7NvQiw8rY
qrKU1IyD6e3pYtPH7PIMYMYyARO3//M/0rOVNMg+nTlJjU9r9QJaC4hSsDAScn/D
26RqPRIJt/jydo1+Tc1T413o7WJy3j9OrwUlwuJrIAyj9i1mwBegGE7NMMV2779z
C/bUO33E2ZY0+2KDbgbS18MpbKNom4KBMDHH7rRBdeQvkexFZ3Snkq+/XWUCvWxN
yIW3O/Cmj+FZaLVg3jrECT0ZZuYMXWeN7Mob1/BkkSLZcF3NFi+ryqqDRxRFTI0y
fo0UXtnCCo6oEmw+OdaGnjDpHVururhoWwuT1rro6hYHnk7oSzhH1inCe9rNojoS
XNcD+sCJlIdIh82FHxFYvUwhZsLRxiSM1XdFEqlVK7KRmHapBGVK9Dj5f5AUAxeh
l1IOaYKqAalcHSXg2Z0mwKksBX8Lmvp4caFPWcz6w4uJUHwB0ytm2KeNbDyjUZQi
p2Z65hrUmH8av4AaahdQYu6ShzFEuVczoWm0zW1cy9XiofVvC/8A5tuz8a0KZ6Nq
QSSACvM1tjWXU8J2lDvQEN1b94T8dMf5pEnWdFOHq7hbAQK4ipl8LAfDuzHXJEeM
/kCGyT/Otor37/FwWmTROc9TD4vNdFw5Tx7SvL6TyyIIzutvyhJIm5ePvA3Ofbtk
F5zrfO29vV28CIqNQ+DKZQDz5zSMg+KUNCQSxtdW/jIUe+LZ+l+N3rrVsV5A9EnL
hkBjm3WSPa0TTclYvssp/kn8Sl8cO1E9+UOnlw/317NkpHXudmuItBuF3ioWRpUV
Qh165qU/VXOqgiMXg3ICmFIQHehqcZlbV/36NSrdKcPsGxNYsGS1xervgpTZsE56
/8AYVD8nsBdvcsZ8uSfBmCFE6l5Ws2a4CRhmQwDItZr9UGtKCYCzYQRsy4AWuGzr
id55rhdalv5OVqqDbjIXPfz/9kKowuOhIJ1lAb6BJL3T3mfcAGPvCacmZQ5dvFKV
qbj/KRjw0HVPYioip3/0Fh2z67a1R9earJ+WPc433QJyBahVo5hU0aZmyMvs92Ok
FON1mA+LbdSChrOmLEtxxZrNYqTlKzvdjXVA2RKZbbO3OWEhNs8skMT5F+Id15/I
pZqAJriR3V9x62acNQrUJfuXRXixaQd9utjPAWw7MN9nPAKuNpRyZyMRktIuqy8K
2iW3XRaZxei7y3dbyJB9CVRi9aWFK2ZaEI5/6Av3r0TEmIaOz73p2ehz/78xHg0R
F7dZUPH46DT/dlhEQNLe00bqEuhhmSK2aVMpFvbI1/zcDjwVc5sjoYYnXw/6fdTF
aisOn9+LFMuKruwTlN2PlTa9At9kgzCfQRqyMMMG3Nwy2VA00lLT1shGUsXaksyh
OiMojBsNs7LNbD7QYR3NGQEQXO2iIBGGCLkGeIHXvbodnCfytS9qDXqMjHDZPRBy
+skcw4liOWMgr8SzkyApbpLGdGMUsfHhb7/ByWyjU9PrOdr96VT0J7h+IAopOIG4
r76bHaDlOIAMZ+ar2I0nslihnpz7gVjcWQu/kx/i9jnhhzM4VVr9Et52Xv83l89f
qMrwg3m5lkBvtaW9jaLHzfNvrwtyTfZITiVOg4B00+Gn7k4SjCTJbD5NcOAdXP/3
it/lFmIGasRf9jT35FJJB6fi68EhYdKDGUib2bi6y+nAtdBF0d5hmgDCexGpAOit
iy1n+fMmQmXq9RnuDja5xVja62LasHhdVC5JPrpgJBYrnfNlKdagQPHrvObvFoWK
O2qpFyDJD5sXmSSTa57KUZTvAorK/wwgopT9b+i5HEuS8eOq4XyqdGCC9zZdJkzl
GJL1gt7aLfPPHNqX0BIn6RzY6mXF3psv0e8L4n5gNphcUbT/wf+WMs6w/Ao1ABK8
YJ6dqWnZ/VW1xmFGhOYlA1tVuzeOs6oycVNspbjtDXBjJsudFsw1ST1rs3n86MGk
4MJZ6/IgAKVw1GL1VppkbQN+JhpAJoOc722hgJFLQLJ4wImmbzUkLlUMqetjBxlr
LJErtnsQx2b8dkVmJUEKaxMc+KN3KlFyeaU/N8eUANpMsttEi9GySHZk93o8wW5t
in+PqNssuBd5DEfMhdoJoFHRYF76J61mThtcZ70ZW/1ARv3Xwkf/K8O77ZS5DhH1
bPK/+o8v5WRe1bf8X6/+AQbuqHeo7QYDZaoNvmrLQCF85Lb2+bftDNgoHgwOQ2cl
tKjiULayKS8LB0Q4iRobiNGnjXrqiiCZ6asaO/zvmlSSEDvXQLklEmXyD2C0j/CP
yLiYSMc3EsBIL9Xz2XtOCHIR/oi9d0+eSQYVxX401kRpgR7mTs4IRvxfGBDIOh8z
SzxYNznEjDGi6VEDnTBHAU8CTIdx/XpSO2BRftkJQQlY5ovuk+yoESo0Vcxj9lQY
jHkYYR800ucqkK+vhFwhuVbUn5ZOiWzdYVKlqpauRiFPyOJvXOKECRE9prv6saQ6
KJ74lVw1iw3F1BAwpj/qSE48l7D5QUXwT9tZaD8idSXaOpLx8I/oZbGxgfvcmy6G
1SaUXGlI23Tzjdp6a7mVdWBdCC2fvyEbo2QGs3KVgO128b7LpRpyZJ43Vur2bTOP
TppvCkOrmVd7CjboUNEFnI3tN0ywirUy7e2ANVAa/iffcr4AaF/evNmMmE6mUtJO
8jNyO2gUQwbKS7qgBRyqtsZ4h3qtZgnCvoxUUGDwPB38UYgEDRcNpHliVv3qXhpa
dNr1wkuveEgewGhvlX5VD98ZlFqT3Djb5FfWSosO+K3ISGx46062GxIGBo9vOmLj
CMJJL8Snlr1dBMsjKVsv1tp8Mkn8ueLlXfhbLFzKY+grRDentc9p2rNP1BoUUAB7
BQGoQCsOlFNHmlCJoR9MOf8QQcCvwMyedWSbJM3zhvUF7jyxAscOpkpvA6Gk/1bj
x/UVSdj1vxpZdxlPAszlqsiSed9p9oCQoKXuRfZfeHnxhkLI5skPSbPPfoCBfE34
mE+YNKfRyNw7O9mJUPI9FlVJgpXRP5DyWSCbogPG9sMHUFwe46nW/rnRFw6/nzZZ
WQFRN/ktEkgE7+xrhhhR638W6lBSe8Bx3QFoI9xrOlmdj8xWr9nOMHriQ7cM4P0Z
E7Z2avi4kSph3JgIO75oWdGOlI/qx0TMlob+KaLdrI6J0LADP0867pIRjI/Nm+gS
KSWS+DEB5/7/kTJg/IGlu5WSDfN8tg8GKflJuy5oTJLLvpfdfYRKvWaLxWejO+nS
7+OlMVQIAu/qNYMfdMTSELu9rEDSNGFCNIIF6Do3YtUrc5CeOCfjcHFHysLdrz1r
7b1z9kbeQt5dM5ENp+LggOB2Ky4UHNl+wgw6ahjm4x5EyCBy0pSq7YsWjnYVbiwx
uDU/e57kiTRU0JILzsqTN4GprHKArdozIsidslPMW3LWGS9umNP3VInTQlGwkmsj
bqMbD4RdSIp3ceXwwyWN9004B5ZgYPuzIQxJJKUOfXDKOoF1AfstrYZ9YjKNQXcA
N/Gw8IB1vLFmTgQpMVFW2HwbajJqeG2f79EvrVBb/WU7E/z8c0Hdo8I03eM5qeV5
vSGhLHiz14LZmKidMLDEQVOtlag7MoKiITi19h/lQoWRdWaKg6x9XNgoWBAJJkRv
Q4D6bbeTYWk4pmr2vY4ZSK3AcwIaEmx7NmsS1tjrNm8FTPpZPwLOPco7n677JQ+T
M8rdCaXPmHfs8Gx+41vazdTZecSxwpNGpewMz1QZJSIM3XEeU4J2BNLzTYwDbx7V
SQ0fiefLj8nBDKNY2dC37fT3i2yGJBnjH4oGnYXMpQquHi0Gcs/QikrBywz8XXx/
zWG5als1KavExsFwMx2+XNkJn/1mnKQcKNI/ACF17ezKRvkEFN8IKtebgSIEz/u4
LLN7oBAwAa33O3TkaAozymQWu30urgypNd5sMwwsn+K6eqNEQjpQ0Z36R4HYWusS
GTlwwQ1bK5fcsFOVJenL0CMMUeLzHCGYA5Y//qFPphKw3V6APf8eE9CurhQl2Z9F
o1coLvB/nDz4DuphR5qRq05QyYunPr0vCQBnPgfuuiGCmB8+a4907BiocEkpKIlZ
Oy/eFAxR/9bEmw8YykQ7a9yDHo8dTYunOHGhpoum5YqfAB2rdWQHuka/mncFABgH
M0/0zoQRfywwYRKkTPdMjzjcdXnAuSc+jzVNInDG9fwRopahICSOjVzHsmr79CGU
RCDfk2BomwzqSmscVVyNihv5G5dYG8NsYX+LY7I+6yeRoU5uay9OycUGhYIqFCu7
pWQIbRYMI8Ms6RN8YT1EYSFugCHuYQb+hm4gsLzepnCPKEon7zkVffLJd6mONQtR
RPShwsnnYxshJu7AnikaF3oKPszRv0ClB2jZlcrJ6mlCr3CMDseJtHwTOE/DKqhb
Ia2j4rtnmU86zynKS1s2UstGM2f6N5zq+S9Yp0wRiqSSGf4+xVhFJJN0SEyImzRW
h7JzyHmVXi/tMy9raG5MxslR9COFl2GguZLkwTs7QqTBVWJu94ZHrOWz1vUOGNxy
RyipFWh0xPsO0dc8RXUh885eCXakgt4/jBoS+FC1IzBTQ1q1yPaw14GbfeXrfp4u
gALiBy1OU5/p/xC+YP6bGg0xzhfgLoqYBS9AKhX/kyQpEpnfwFatzozNGg4KAa2A
i3ttzGMnlEmdONL3/ln3wx/7l699FmzGdVDWnRGyH+wk/nADkm/Zbky8qNcJTVXG
W897lCJU6uxBU1rf718Q6HGYInGRLpta51sKPuuJzlhRZAw6YuSiucpGTAPnVvPW
RVnOvfG31vdiOhd268YBmfx3szKyEFfrJg6b+bgI8uItltHjOIKm6k1AUQTntjzF
VyGHZMLYmSLZKBVlaUO2fmeyVX+CIefr4k6+iL9vp5GSymSzU/BVbYQU6E68I+03
OXFTbV8E4bHMu1WOLf8fe3W1B2qisk2JImnnVGtzSgwwLsEkSHoTaG173mSgZ7ia
ckDZ3nGhou2D/oL5qTJT4ktQNzqeQR92z4OEQFteNErAncbwn0uCAZy7twLlq9aw
o0buuHyiBsIAES2ox6Xae8JiJX2/MubJ9tKT3Xy2wQUEGLaD9uJY3T5xXwJcgIpL
VRe5pANqadnODOXihQNEpQgrOOmSbuPxkTT6pk9G2KcnwV4ZMmQlCwUjDXOI9R1h
soKz1e3rNlQ8UQhYvjuNtnjk0acXRC7/kr82giMw/Fzvj3+8zz8c3mnVrUHJavAW
Ruhv2V2v2v23/gqcyBAxk+JUQ4TUNmDHPOeIfwDtANjPB/UjxenV5xuvFdVBFfRC
NCfonZ8gVCcnQYO0M8OqfJn3gR4Pkg1cY9QYNX3LXhkFI8pmTszqgEmtv4khj433
XsJHf79bQCwSEYds3ruySOZtT6jJ2/+8bcmRfS+tVdn+B5pUw82w827L3DfvIomh
y4SWTfE28FWHSI1ei1zO9bH87+E1Eu9+mMrUhX2ZIkSnhz7/UqG5fJJl8M0mEbyy
WaHQcq7kCSmpQjfYdBsK2PjrjEpnHYu3OjkV+stdY4VzLmFLEIAUmJcagVDsL/Gm
JdElwx6FrMIUqsrP5u96sEgAUhs0juMhkauq/wTj89BLN36sa8hpcBpGdOnK8+1g
LJACcS4e7bjj3odp7d8JwWqHn6InhLT0yGLHL5LZ1zpjk2rLwQGyslAnxI+VrzPO
Jx9GWAtuokf/wbTEouTSJADhtvTIZ3e1VzuQBn0ycOh79U3pwAwfxBW8AsXk3/YI
DAUJBCIG6G+xlzxAb4xWHtgVuv0mPE16JP0QR2Dm3XDCgH/2UY5CgtSKOdjQ06IV
4YW9+C+Z9tBMWKrAnbY4HpmU8aEw7Ka5oRGdANFCyY+lJk395y7f1fXwBwI7MmHA
3B764MGUEwgi8tQGFDsIJXoWGSg50OLjhoa6MtbDkUSE2XAKXFc81wMIQFezr7Ao
yj7p/EplHoOBjJ5Tw+cfvN8Vp5NUIYFiHtJZ7pnbLx9Rl4B/GzJFGN5hpdq7cVz5
LbL6PFHcPS/6cXnAeW6fgjPBzFBOf5fqKv5Pf2HPtoOZXSiXMqWQZjU2ZbcDfzGF
tMvLbN+4GsE8SpnuxLejglNstpKSsiK2VaRKiTVV5WS+F6ziruBQS9Mw8VWbJpTS
f4+WgdxYfyexzNsqHiLxxu42UL1zZIunmHsTiwnJOaFXuMTyoB+F4KYLA1MopUqo
G2cwq+bQ0b+DfDZpwLM08FandeiSCp8lIReIyAzfcK/hwBYoCqejAnRhJW3Wn997
HwAnM/9EpKLOmarG0FRRnDaSiJJ13gPVEYy3pO4eESeDhq0H1JNF3QOsjqeNUxdi
AfQ6eFlJlC6/w3mw0sq2VVHPh/cSUwuQ/ucKlsZEvdjzqxLcki1UyKrahXWH6p14
BKDDcSM9ESoGglc8hvm3Fmpv1Wu1DdQhHBL5N5IA76dnfya8CeN4I8j1yqCfO+k6
RZ3V7qJJTvra18KAB05uQB++GAyOpn5bKs2YlSonFq8pZWUhfM5F/n4QZALWL6d3
8LrgnxN3hdYWKnN2o7RrwLWen0RaKK7SN2rhZFzm4qVIXHPqACYXdJETG2Whdc+S
V/QE6LxxSKArwpBadgaTDWiyLPFv1g4FT3frtybdxgcI2YrTZYp6Gxq3yHOsTY0e
ZCqSz9kGv0r7B96UPkYOiSC+aakZBlU3TefglfOzdsVmjX5iOyy00SIDi5CcA/84
JgLr/dsmEtO1xJ5IdeRRqlSAETuTQhS60zc8hdxKv7ENRhQAK1vBfqSM/MzizICQ
Ei688xPDCha5U/G1JeuhA2gMS0bVYSsbip6S9VZ+MHGqLoU0xHgbCUoFl/QOGrMF
lRvTZGsoh+TKNx4vCKLnrxkjg3r5Tn4S6SCdsldrKeeouAJd5cp0biz+nHXsPP1z
tmT+xc/83+YRZHyaFdgtfmiRE6pQXgcvarSWOkxH4E8TZNgo1qWs0vO70o36ZzgV
Z4rf1t/4wEKoY9/XX39FSPFnR+rRof5kCq28cuon8mjCtnt5I5DVjMHxHj7/8YOk
CMcAPAsyIA1OK0Vf7Ffoj8lqmyLth2uV/CbOE3TQfMkIZYyR23UHgfHy06kNZT9a
TbM2AgsKwCxFjrvGTzQh5icb6FK7uwEq47NWZ3trzIENNDQ/jcBaU+b36MpeNJgy
36jymRj65O7kdRexdXm7GsDh/OadWW1Dqw4ldH9fPvkaAYl98DUKvHBlaApPxlU5
3zzVcYJxR0VxqOoBHq8d48C5Jj5Catpq4XhAQHNPUhyuzFmGuAbbJ3F6xZ4ul8Bw
6cbO5fJeBW2UYATXYTf3muLCVO74+2l19CNCYNBpO9Hk3pxt9N+jHHd+qSFVczg7
IH2vp9NYMYyJrYBVKbTT6LhDNN3Idndmk7ptNke3DdRK4RPqyv6xdcbbcD13A0mO
SqeGgEOWLvhn7lqlaw6O3nAskXwWWq/HIt0kDPJdxV3FVCDYdnapAXiRFiS2XOWR
TV2LTcKK01+MjhmbM/NIaBNmTxXUrgo4+DUGr4lmoAHmkA+tZsMPsmiGkRBzH8EV
4wy8EjYgA49FgbsyH1QWpGTUE1Ba/9LSeRr2fbRJ3tc+qdyMw15YQGsU6QWwa3RQ
2doM4TTq1M1+tXz/pBuNE8mhQzZmlqunou7/4CI79C6QVmIo//IxjeigUuz5WGX5
U96AHsFyydgf8RxbHRK9C7oAcPpm5Dt8CfM6qZxhqf/mSlG2J9H1bSF0md+7W+p2
KvDgeFgv1y4twsedznaRhQWTgoQ2x3+EIpEpum0QK2d1BTOWCE42gj5jcNNhi4az
94jVM0HK/dMhsSN+PJmEH8YkZ0yv1BR/Ux6hMHieCOjz4+ds7QLlB+JcOYAoVnBx
oJH18QatQIsvXPSBn3yX1WkvVOQ8JdG24LHrfdWazmB85ptTuMMepyZf/20pcx3c
mu022pUTuUyfXv4K8nt8qjxfRDbwVjA+CafU3pV0hlX1FhiS/P4Qbr2yfqvWuXCu
o5xG/sZYaCDRUtIBZJ5p2OXw9pVHsZ6HHAb4iSHYVpgqyccJn9vDpBYav0rXOQUv
LCcze0oXhZLQnT7uw/13H6PB9msOci3zbvDGxZj5IQSRtSu7+X7/b8S+/WPj4Z7n
uav4ncGqU8TrAvqLo4KioOZvxVLFcTu/cU72hAg1IIwQt5jlFsTjLT5CuvP+9lFm
yEY3kQiVJzwrXS+4TwF63iP7AoQjo6OVkEv9zPtECnOmxshs68nsT46YuAqRTblx
M6oP99Y4va0yop9LFLvPXo6/oTpCptxOhsodk1mD1ZDgP/+cBUZyhvWieq23LrA1
+MhmuLr2CEAPzodrvRi4h/5litlhKUh6JVQ2DKGVUMeyqdzdWG5q03QCFZ/zHJUA
V/l5Or/OnPf+KKDuxC5Lt5a+skug/EtvTsXxDzfsgfK1nSMPSEoTsvU20gUaHn0Q
nSqL28PdgiQOM6k3/pfykp/gbR4iQnH2EoorxBuZazMv7ayB+zfRVtZPTFaHgb84
+4bVfJuRNcOFTmRjLXUwUX6ksFxhs6ZA2UILfciNJYRqkRGJBSu5+UHbEAuTm/VY
Fo+/W/jOpM3nFZa+33TqSei3WJuG6ThxCAJdkNexCsfu4Svq3ROeJubLy3CCKNMR
Z0OfdZ5VjI14zW5ADdC8NvvNskPgUCJw4y9V8+AbGQ7gXul5kkFu9KV1ux440XQv
fgPCyUmKX9C4UKVhU2p3/aBkxHFU5wo+uPqzMpCKrksCREMrafV534GdxspkLWtA
sM5RUAKvkUb3za9TfyTm0WYcmHQaJOnqufxMEJ+noFwwB5r+WHyICw2IGpYarZFb
9rpyvmo8zUruploNIOYA2h3jGNCG9Zm0kolGXhtqJxSaDyTwTjteGMYtLZPldduv
ONvmWscgX7g5NsvfBuGxVJeWzKJvkY2XwT2zF1nLyjidpTn5M9erdx3kyy5NMnFu
LcLmxkcf6Ido+uKp9bIuI8Uqhk1DXt1FtDu96hvjyDXpB0i913ZtCcR21Kh7zWOO
/M6dBGpQlHp7mYKD4H40qZRVqsvnXQ4kpLb+Fb+kmrxKGp28sflZrdzs3t+fVgid
aetKNJ2wBqNul7pvtytGHrFo/aRRdl9pxMOhLRXUYgxDQyPGUyCgwORL4C1JzsT9
afK3hiic8Ip4LL76SXtQek4jUQWdcfK78M/lgzu32yBdQs99nY6eJMWSXG4uxtCz
C/75OriP971Ai97//3dtqfqD38v9muzl0eexbPtd3Lmz0SoZ8hu7QjEaDEHvUPFc
EiPLSKZu1YzepPZNQgNlXXklpeMJkBngImJdgPO6SpeG/XszVwprg4mnc8PLqn/N
uKR9yhAURZXPIz8bUVrCr2VCoPOT4GzXiNvLsgJD6yNu3Ltbl1TTJ8+rTmnfsZ8X
AMe28GIB5dTbs+zFREywqZLOla92s0tJ8n+lBiJRc+AFQAdsB51n39l32zJ5EpEK
N6/oLiu++sy4u956fpHHryyjcTaOYpnDwVPyjTTvKDptVvzOH1LxXRIfyyX1lWCE
cOayF/nPQzeHJHOlwxbom4YV9tZH0hK6U5DQOAUa8Y37mY0W7mUFgfqtOaSDp4k1
SErtEKNgdmwkcK3EMZTQZkSzJjR6XEwvcl0Ez/1LNnNM8hqprJ8MmrzE6GfmZhsJ
5Ar0mmh5Jm/FimyKNNxAcb4qC+PgS3Klzggr7QdgtxaJ8jP2koZQ3m45L9yr+H3k
ymdvjWMlwtxsrJBmBvtGh74OAq5HKywkcESGSxRSJu5YidZCWa1X8MhH1HoVu+dQ
hBu+xUbSMnaDxL64S6oXZcLodS4nyfizA1WzZTU3DbFaNOxfXyKhupiQIpBGHWxk
+VwL6DKo17veoYQvjgtyLC5DEbHXfXZ1OhTrFpsCGYs/rFCg3pUKtquoS3XHWabQ
HrSN8LuAGBjXkRDwwQ55BXMwK0DsnZiQtOEt+4pK2tqqHhty6ZCjk2hqqSY6/mGq
eMyFvFujTc+41H1+ylcdLZFh19GAcan6NsVyEZjA/ASo9UwBGDoEevEbw9Ou4Sbj
+GVsXpwDp7lxqiS2lMeJz6SgxAHpliIrnDS3lRQlo3BqnE7w11ZagkfiM5Qw85Fn
GrhqCjcWPkPYBtl9pOmrdy5gePPTqp/9GGpMXdI0DTYOiIioJNVRw4g3W+UBYlSf
6fnbQzOr8ipbalaWtTthM+4KEw7koJEjfSue9Anu5Os6bm84tl3LBbNLKIusnwkQ
p7E98HSEwt91El4196EeVJnrRfawzdsY3zs/okBZxnwivOcD2ER/1SWrh3DiAKyI
N+8BlFOwfuBNxSx+FVhQd7AHfEsUqnziRnoarzio2Sc0zx9lTmcIrrQBdH8mhlUp
Qo+Ju6iv8GX7b7M3BQ/hFu1R1cMTTyceosehV4oqLwULvaDQgaixJJzcsLASo/57
GTpT+YFjUyvIgvLhH/KZ8kq+nVtq8QT/cXs+CO21ItjPb/BrkDo8QrJcSxuxeX+m
pxjFvGCQtlYLS0uhZFyEioqecilTsuRT+w9J0bkKnGH9tRwqw4xDMALfS3oYo7YP
MyL/oAizgzSH8aBocAzguT1ItzU77JTN+zx1nXzVWdqlJUAs0MStyLuJx9MzwDuT
mpUQ0UszVH8FoFX45pY2EboZFLBxzk6AeKKQlRvQCit880z7KzWPdHRNh8wVsShQ
rMca9PWa4LXU+MLvYkrmj+xKB63vCqJBYU1ZdVxO7qmb70kNhY3i7Pxv6QDEgndV
3TBvxYgOPdz1rvwrlvv60y4eaIyxRho5VN3cfY3nSK9Pz+stbTMjAr74nc6Zn5Pr
iAPLXfPxgob8Wu+u1e/Lf6nkXhCsvAbY3lk9G965xHHmZQuUu219EKdT9uC09s+W
Xv2cCO+POllZ3bAABMmP9O6JIIMLGQaql+VWwgVtVq9Nhwr4nwdaRQUgedm0VrNy
gGjbHDf5+VDWpa0gs6OWVMFjY3fHzFNr7E372SF4Py3WEWy/vSi1hZ3r76t8dWB7
UeFk/Rc4ExTWMhhUnPFBOo4aEy7n/Cq0E+0b/hgZuQkxtJH0zXxTsvDO58reqtNn
9lLZQrQm8FUeD8Wur0Af7wfapSukFrEAeDQPItB9qBRBcxQwQtWSc07ZDw7bycRM
N73kuVUBij3gRt2kZBM88OiilERgB/FNp2g6JY8tc3rtvlGvrve0W4RyJzp57cj9
bXVF8Auox6zC7JTM2Ar+PfSlyYk//OK62oxIJ2gfYdJWtdi/wA04OGpPQy4S+1Mf
2ZLMEAPcnhV0p5yens29bT2Ob7F+VJWwZkZ1A2et9mpALKb/YOnY2gAROrTLJlWf
tzjrEtAgVBjEQRrt3q0RM+bAjkrQ1+ZsATcKCeRQN4IuGHrHxDbG80ja3I6TEmqz
kqbcuevW+ZYqcnWA30nRSicEenHy9hoamVMMHV10N/Dq431fa2hPF6FB2Gr0wH/u
K4XqStLZbU2mfZVo+JFBn+fdIV5axVPHtM+cpep0jOwcn0BHcgJUoeBR/efX9J9d
cYOA1P2at4LAhbIJ2UM8/ttMzBapcfD/dz7rKzQiNl+CoBlUYinswm3d5CwcuAzW
AyeuH0wJwkpACFlPwKqCxfRkTwExIfw4t7hkRzUij/HHHl/iRX16PXrxqxTvIRQq
gUAuEtPZxaM9+03Mazwmzy52/SrC7W42C+rbhMFxadLNSPNbaQNLKWBCOowNup3W
3FS6Pgj9GFWFYGJgbPx8euwc6CDgvodUjMjpJpBDmnJMsvPkzq9/zoxFq1G8xVFc
bUSKZ4oaF1B4jGkebRfRnbv9mKqMJVW/PbsSl7kV85jR2dB6xMHiep2BCYNG/aAw
rYK1MA4WwR515MI3+XfhVtQMd+f3yD6Eur4bZWoJZnJj/WqUrXwP0wqmJLLcIApi
M2HOUsXxjCHuGu74ld9M/7Db92e8B5KrPDtrVIDc91JUQ6TPI99kQnsrS/sO4aSW
wC/KSQxpEng5ewrFarAf2SlXClAYKhaoo2O3IQy22P/+hgzHz5efnA9VYvL+jMpv
RrpLAT9EOAL1zX7YG1MzrWwJq01BXx4pLMs1+imIF00tJJUHMTjHH1fDhQF5eONV
ILp0j8A1fO+Sa2TqcIdqFWmjqJLnQjhIaUSbWLHhwi2dBy5OoyfbpO4zJ3w7GQLE
25b5R32AacdKV9OHpsSqUmGGA6JS9m8b+Zrbcb3KIz7RrTmjszEEdywikM2iNabi
ie/XYQYpv9df3v15MOYmhNn+fnI8E8BLxbI248bv3GB757WgLln9klvRtvR/ZY6B
2Zq3hXg3vsjSRwtk0/disgFbcFWQkRh2fkDsg/SzqVNTRn/dlN9Zgpw+ltlTOo2+
+ErkzcGrgaGEjNKtczHujGwRtPPOFRn0zIeocCOsYiYRRqOkrV7fH6Maikh4k7tE
dSOLYw9hk2Xak0IuLp2XjCEMG9rOv8XmydzChKVqVvejUmKNEa1svZa8kXKCUndG
XSgRR7WzKpnyRkFVa9lo39Ga1Gc4BLe/oHnl9iczCUk7mCAVqhSIxjlG/69QTvzU
pljZR81kcwX5GqHq+31SHM87lji412GVYJ7FZi4NuzMKBpdXCFGKbMrG3MNIMdBL
xaE3KxtOAb8k+OvxSxo4Zk0FkEIVa95u1iico7BwRd1+g89hXcNkQrO3heBoHl+R
sozQhrq/ORiBTIMFEaPh0y5vuP+Lvwz2aBLOZx5TZdcr0tVHccV40HAVtdaLhuGY
8L560osaEQvwaMdd/a/hVbBgl1CTAQF0+rBZ5Zsn4RpN2ZYUmTM0d4papTH7Q8BV
80cZGd/G6TnBF6F9frAn0wuEOLgEReCS1CnRB7e4831Q2uhUIdEVj2dxFsjHtXBh
EAyM8SvMJQUs4Wc/MhN8a9O4m3rCQqhHdM8+fICYAPl40ulGMnQNHCBIRePEbbVH
Wd5ELshu+nrwZqYupKOk9wSAUKS8RPF9cHDniZGGutYVsbKFr7NCnayreQz6fe7l
+y6mb3Em8cGwylZbllZvh0RV4HKkGo++nO3qwaK8X9ToCBxqcCNlM8N2dwv4uHE8
jtygZyoc8sw5PzhCNmJMwIE2b9tDNz1q973i7Dgyz2kUPJAVhb9R5wo1rQoPduP8
qqrYn57W3FAOYE0lkx46BMGOu/+IakVjVOcWNLYlrkK1snEvA5tzLkXC+fode+QF
Hwd3GFnSOvDNkV86+IVidZJ3Vwvm5Dy0m04vSZujVqo4D7KqvvyUk0dSHhtZK49g
6qUzd3/5EH+X3YZhTftnMX66rKGYZz7VasZbjZpNekk4D48WrxZB/2B/3PhW+2DI
Yfrx6TFA8uLWr67QADIEj4OSXSA/jnCdpVM/7z992jv5OEAFd7WilTqht1SPzzmV
Bp29xyY5djOjyTZdXk0Z0cbVytj8CCoouQYSTYg9D9sVZ9ZzKzVVci+OWIVuXlO+
TaH4aKvpQauSNm9+8+bjKIKWQhaDrRAmGAghxTB/zkLoGw/yi0E4PSaNu6hdqen4
LmT3ZT4Vw9BID5InNTxGp2fhWtORjIuTR1ym7YvvnVYUu7gWxLx0dALdjl7pMNPU
cOb7E0G17PoQQnV0kDbctl+cgSsW+NdyfkGVYEQaXNOsg2pKYEXOEtxxkZDCfHPL
/gSQ5aew4S/EqACD1RTJiiHBmLVtE8eTbr10GHb/RWzRvTGkSNlyChR2GboZlhtt
ZE0U0M+c5960kc0cOK1HxcDT9z8+SN8DNerFNkm93EDDI+3b+R+CRwQkeoYLZ/oK
Z5SIDSFY1wKiZa1pHKg+QeNrYAV50/DrwHbXGCQw4EnV66FoiTouokNvBIE+uAVg
XXSYfQZUJlz1g++Bc9U6QNdvrEpTtdBInkuosfhlfFKd7Mv8KcIVa/86wSxe0xuN
C60NwZP5zpqP4LGsx8wNUkflQOXIe5WsK3La8NKrb9Mtq7aqPbXspgEUUlQCQBNg
RGWYMLuFGov2U+uyIIBTjLs/ElnmuFn8+uqV4L9DUPZzTMTzIRwI48LW6Cu3xBHN
TFDCL39nv3KnXLV+3b5RUK3Vca62d2zf8QByUAHbCRYfEf0+t8zYGZa32K9Zz2bF
eWTtvcYgLYTqcHqPpkGZ/TGIhvnVSxw3TkQ1rZcpUnCo7n5uHgJuhcikXp/KOG2+
VD1D83boscBi6drq75jgQpC+4JhUxqwexMDqmLmPDq5sDmynKgqszpe7GHVV1aPx
m7Ri+Ic+xPVxyVNaXaEFlcAJuvY6Wc6y3PFKnB+v6mrTJzDoHuMfU19jl7jSSSvr
bCzZxoxwjNpIy3f+/LWt5YCJrpSG3IF/XpvmvS45glfl7F389GTlSdpeAgXf4vWe
o6KgV5MlhtMHSGgHdh3hits101QX6B+iVhh8+UJ3Lt95Kg22xl37S9J7zNynE/LL
m1YzJ3LQF/HfYbIqMiiNnKkDU4rOqjGbGz07RiX/B8mTWJmBb9bJTCY4uelg+gm/
95cS42UD+y5hNl3dQgyi70Lb4Fi4tlDZnyzx3s6DlT8TEkzwNhBioeU+lKmbR7//
fPqO4K1PdNSQAht+6+sVmStNmQXp6EnzSjH8Qmycz0si3hnkfuzQajsYRAPK3WCc
itmFAAi5WBf+1ixmCZW51XidznAiImquGPhwepfbGlIaVJDAKXql+YJ+OMi2SXvm
U5E+vPER3p8DLM2OuX8Dtig7AM5cAphY018I+/2uLe9hbuSDy8kpHPjoHB5aJyRR
NC8LZL2KrG8CL/mbEvh/1F28ZuC9SUoe50cCvAGHQ0sIEJ/YmRCuIhhBz9u1gUqN
0nmd1dlo+FSG/B26LFfaPCX+lnkzWUcrbV21Ck5DCUDJoTrBhp0M96ieE1qK33oo
jEW5mBuDMHXJhsVidhlJVdPpnye7arzQ9tl15uRFNOCqYBWADnAncz+ZkY8B8q1+
QVbi1qAGUyizCq4HtSSf/QoVYOGQyujfuFHkLQMpB+apkSYS1eJtnO+GZZPdcC0n
lcpRDDMIaYcY7KJXc1to7M0I7KTrQ+OFxyfRwRqP5K8a9+9m79XwAQpbqzZJIjdr
OrDE4m416OblhvMRy3RoCTYRmzW6AiKBbJpLNNK1WCEkKjl6ziWa5Hzkja62rPub
Nvv54xja/T1ifiU/o2f+K9XLnTrYRVS3omEbroRzDZTXZaDj87t/u4I4lop1L4ix
AZgEGxeanldV3I04LiJoDAoOYY2WSMOjlStboUBDlEglIFsxwrR/gRBkN0TD0qsM
91lY3M1+gps9Q/wpJ8VASfquHU8/PGdimsXl7D8wc8I3GoEj7LrrjU9xBCr2caGZ
avFF61IKF34hq70wYglWLmkQb8gngBQhokhwZKojF5FAeW4esLyPVUpuSEvc61+z
y0nIDeoRn/rIJS6d/0GkJwG/npCCQOrCxk+T2OcgV+Ebx8HdnHMbM4lp47Vzzfd9
L7oVa7lVmD3QLIiJeXy0Puy4Uz93QUeaV4atJIbSrx+nBZJFmhvngDcmIc06P5/2
ulDE031vCu+LvZk+ita7ydaOJg1QD30ZX2o0ZKooQp3k1pcphs80WFElD4cLPsIz
L56etibjd/hWMoiPtIMzQLE+34PPjsV0EIItTrdr3G3yfVMnFaOAlaNc2Sz95uVB
Zl6e1SsEZoQuvqLPNWcHl7Y4NRJLr1oR9NC1zS8YFoV3+cM9bsiECTk5epzUBj5l
eo+XyThmM5tN7Rqm2ttm1xGuYbyjmakyWdoPHTnuhcjPK07iCgXMJLRpGPqdNhLb
Okr4cSpbgVe/4qUMfgmik+Ogl0kMAPgbJmjNx1zKdNilzC0AbPAYgJ7PAmIsZwLR
G+sXCwJDQJdQzygWyeK73yzPxItIzfEpjWF7IpdsvPsu5pSHmab0yTl1qrGnBIdL
3pgkec8dmvC9y8e42ZYXIkCNqgFQwfQWkrgI8Gr4gMfL1bE1snVkkMNvMBDQamOY
d5qyzBd8jLWAJsZVukNkYmUGVYOpnbO9Venm84rVs2kKtTw44AqMGqqwG7rqs6hG
Lm07drxzsekDcys1dUds45YkPgxm+sq/OGcAsGvs4zc6n0vRyc4UK8wbsOZiP5bO
NczilbVR/LaHsq7lFqY/hMZY6alSSETmkvsfNj5EE0arVwF2xIegeXNJBP/6vgrx
YQwgXMfa0Nl6/t1YmBvBCtgwvqCqCcV8q2KEp2+TjPbRXp2CHUtvYSx6ZCBv581h
qX2oZeEUrvEH8JkP/j4e/fO9yu1XGROpIxoYFqNNAfdpoGAc9D2usvm3HO9UO2qu
3nl0S5+ZrmXwKzs0JU+Qf4Ra6IdXTB5iDbpD5Ay90PV7REzuChHXuEsPjKDyNocU
SvppSHBoLYk5l6io68xarYJQcuz3v44hWXWYJc6Z9ukhxMDldNAYHbnBmLxy/G8n
jVlU7+Rc6s7b2Y+H5tDh+tP69PIWQ+yDN7fwq9tIKg6XXCcY9RBTTeDQ/S8oXQZR
+ROb5iDEAO3RNLmtiUYJ1Dof+Anzesq37sorJEAB0NmsOl4JKQQMyFp5sk3LZf89
ymNKvut3fiT+VlvnwUXLbyq6zSwLXLoxoLDQeh+/6cybwXnfC7C7dRip2NEBiDtb
ICX8lqS4PV9pvgiiL4FrR335+o55ruZCYibazFfEsma4PViw8oweggvJH/5O8m/5
Ut0/Md0R+uoHoIfwWsJYD8IA3SrRmaaB5V3H2s/4fju+kNHavjKdkE9AxlNF49DX
tGCIVL2GlH+ouGWQYWHi3df5HleoZrLuDIB4DS1VwfbGytVgqQC2m28ntXGmlhqH
2VIym8Q7UrE0SPQnE8izB46YPR4mDESsqq3SJ6pSI14ocZqohqOkBp1TuW1Zl5Or
gz+80YOo9YiTxQspMb+igUalyOu3cfb/y0wwsVY+7+nUMlgFpDbHkTcBAKUvmF2i
VE6Y6ypBMEisMt4TvpTHcDq1wZdi0nSOSOQcy0k1Pj1cjrEeK/aKtUpbezR1MBLu
sViO043xmQK/BYd6B4kGtysIcFcTligytFXOfYwYpJQHllLKmVdE0UU+P7BFNCQo
FL7z7MLS17G/WzKRGNSA94vX4HFmzLPUVESeFfNqldpxoQ3sPwXury6Xa66iTuvF
coV+nsDEYmx9qwGpkSTZxHuyC7MVaA7SbkX2AfHHJuq6NDDO1aMtqk3dUbVEvdi8
oCKsfNXfxUqTImuWHjchHB8xH6dCXGwgeKCzvroQqmrIfaHnpncdSwWoV4nRaRoZ
W+CMa5oidRrUGgr0DsUV47e+uUizd8AzV5Bkv0yzSHRLS9xkGtDKYUYOkEdkslH5
ZYChRP90l2xv2f4Nqz3sxTg7uttnons8DJ2L0YewuxurQjY2S0rXuAuVuRoriQ22
VYxnBGOViADyrGMtqEh9t5u9sMs3ABnG5wf337XCDbNMSl4dFK/x+LWCHRFODyo2
ziN3QleEgETRowSgANfkVYyqJzHpXdD5WbwA/eXR8l+pBHMC7zn95DTy8nCusaSE
vq1nUe/BphJxszZAH4IQ5stM7BL6ePIGuL7oZ6xSaWCF/QM5ixaIXlboKsdscqJL
2pi6j7+pFWqLwgscDTYuHjrieURN1iMxP+418sFI+FMYHPxu/QPSdePSNVPe+fF9
IRG+uAwPLXCv+rUwY+UUVnOFuXwhFcvbOQXYKQLUW9aubhUCmGQ0RpH2orZxoxFP
EqMSB+YGE9BnN1zVaCa3vUBMxCqRXDrk9Fumb6pCy/fusJrhfiC95A2mOHJ5xfRT
trNehNmyWhMCNY2KFpR43GCxL6CAa+XWOuaT+azo9gZYImFNXFRqvvpheYhqEvu7
w7g9ww7hauI2R1QsrcKqUxcnt3bG12de6LdP7vBzxRxakYrDG8ShYA6oi50yb4k8
F6rdFwsdj1/v+WBwWgAHrDm01TKqkJ0mGOqsFb9YU+I1X32IZhIgae0unVeMG8DY
XY4h8iptQAx1r6nTNXlV1PXU7kNokwNqHES4drsBLy95ql9+UdY+z67ED+CddcIn
ME42YN84M4eF5BKBKkI4EuOMtV+S9c9rDTBI6fmEM+XdtlU8iMUSuJnyq/6Bk/Xy
jLd/v+MRo2rDyagi9b52OyDLQoOoAjRd3PL/tV4AUIj0zJFJhdWGDHlhab1bfgDu
jtJnM6iVtj5DbQHWGC9EfWcDyfQqywOBD8aLzqBhZ1yrMsXOArEpomZopyWs6DGy
hBRDSdOjTgmrxh0UJ97CGpRx4EsgyLsmm6T2hicLmGuqe9kK6br7h8qMklwHX2Ew
L7xY5rCLFDuvvNgFvw7kTPBdkL7JH6jy2xFjGP25C01acdAUfAhfwoJLMAxQh6KS
k/72b2YpUqnpnYRRbSGYCna4frNAmeQTVyqmuh493wnwODyq4gFll0WA+1pTCekt
dNl2PXjCVh+1TrETIGxpfOX6hKLL7suR+uUjNVxSH4IUqvuo0nW1i3PkO41h1Lnt
pOM1/+V0/bwpZbAOxczubMqbbknvm167Gg94LuOELmkVPUvENsl5fsqYDHpUt64q
guMhufihPttKAhBmiLMSQ1V126MP22kTh50y81W2OwnfSl4oa54EwLcLwaM6+N1g
6shSKrs84ac5tC4xAYAur8GyLoP+QLQbatyVX17CIUYEvwf22yrH8ZT/79F79NhO
P+MHH2wgDLVr97rYkSBJ99AREXeIKzV8C0GGSXyyPaSxMizYBvve9jkVvt0Zz/xN
1xNv3hJkqPq9dzD9Nc290rELdXAv98ClO33oMcMqwOg+Hq3UMB/FnxZzfCvM6JAJ
+F6jS2RwlG57ZEzzOpZyWnh/gwjf19/eymlluGzs9byVxc815L0DTkRBeuo73s13
R71Ucmi3RFnanq1qlgyMaQxSGnoSFn/kEKmJFHEKqgdsyZIzHa6l4ELRvZn/brBe
fqafW6hqY7lykINobGN8dICXnOPDZX5/VNkmq33AR3MGDzwaqxOEMena3EGijZqt
rVmIgdLOHU/46zoDrHQd7xNUPm3xZ8gNGotMDBdXTH/XIs8Ywqjx0+5Kkczr02Bj
qs9AQjJPN1xc117y2FHkvf1he8TCKQpbhyENKyzbceTHI/q0SO2ukp2UgEAIgxaJ
q0kZCMjOUd5jwp7xeznkXorerWHfyacCAkwNTfcfXIGFIJj6enwEWBEC5A7gm1oP
wczvzB9VRx2Ps3kV/ie/l6r4R6rjHzAe8TXrDHIKJdBGkltXP7wsEvyqRblT4DJV
98QMCwAtqQxBx5OfHfsaBugz0HbTgxyB9J4ruFI+x9fmYjBCSkTxBu724PBcrMKe
Pm7V2+RiOfkjwGKJzkF+aRY6Gd8SdblHv3Jg9vd9v8n3H9OUddLC0oCXTrcMC5dj
zumitsPHEUg733knd5KwN+v4G6zgrnD2UBAI4S8dU+aLznJ2vZs5URGgCxRLFgBL
XWa2orx2iI99FZWKxoRQ6gIjhfU6roASxLvBlmr/rkkTnmWrifQqrTvYjTXqJqnr
1TcEd7X5bHdwd5+T1OQDo+TCabZ8tEFRD4rjGzms19NHPZ7U7zKOnHaXrP4cHHCA
gDBmmyPre1ZWsnUWM/5Xa1eALKapNlJU7uTHvBN/xhu+rrMvQJO441qd5sNwED5a
CPfZAPPsZ1Y3IlpEglG7k8ZJiq8KAV33ruUGKAjjl/Vmq42qwaIM1OHddgkUHdqZ
JfEHGNy512MGlEzGp+QaEHjjQaotQu3Ge/Hfh30HDvB4wglzR0A1awXvYlwV16hS
ejTkRQ0qLV0AMpcvgxjB/w41G6LyvZIcwkWuNz6D+E0LOME8LtGbMlCcYuPnjq6n
ad/XiGmMUN1BmeNU3v71v4UHBhseDjMm2ci2Nfsrg6uEOimKHK1+0Ixo42/hlbye
To7lQZ7VjyWSRgCJkQp9s52rtdLAYINuAYPD8XID6+RyWd2LcAWcxqHy89pF9H76
nbOzliqhaopRjixFjDfMjM+b60gtnlfQI2bR/RJa2JIGpxYMg9f1i1bjKSBmL3oD
Zbb3CO1XDLGSDIL/UG8c80JSiYD8ziFl1eKpjsECPcS+Z05CHBw2S+9S0j3XnPW/
tR00saXYZ406x7O9E7CHHXxcDBKHfii64qa8XdC+hj4TDk8Q3aFNd5w3k7bsEn8a
tnv2RlyGI9fSVLz69MZxf+ZYNYAWig4EKIS+Caq4/v1etwWet9F/tv/rSnkXpt7j
sGW2lutSL7FqfMViEgphBlL8N0gG5fI9qJSowEyPyPx86MzrpH0FoQmBimY4EnKT
KKpDbSLsvJDNPif3J0ld0qxqFanOVCh3mWl07JJBolHuyENWGlu/TdsQe9R3UJ6e
Xg/BFteZQWHO3lLtFYLbhxdFl0V6RcksH520ftl5za+CmfzLJ/UybldRbVKXsqb7
0URasdKicHIaB0uGP1UzI9qRYfvHt/ccqqx6qeI0jHV9EusvLAIl6vHpNrMJprVE
ODOGgvYnGyUdOZleV/BTjwbGHmxK6J2FB1d9fswzoaiSuj+FtoOCl7aO9VR8c6HD
YWnLb7XEbUL77gr7QPojCNEaNo6YJJ1MyKUUm3mUTZCCjTmfYnPTCG9uS9MtWR1p
/JSnrd/wNLPZPx56MgJjlCs0jsv6WndT5Et4ACSQM7GhU5OD0dW3P2AFWgt4U7EF
C63/y7KIUP1OCjO6gv0fpFjj6vCczNWgcEMuBR5t2O0K+eBl/HFTScdp4bxQesYZ
Q03LEE1gSroqQc9id/+jZGprtujFnbKXzz6PMad9zvzMLOk4UL+QPDmcf0sn6jX3
EnYrmeLoHUB+puhqNbyc8HMYZ1MPvjmh7fBfQUk/kmiUDVEaGvjcwKQCh9gxEJgs
lzBFSa4Mh0Gwg46KxjJVveNwllVTOVpwPMIMXHO8Dp9qcyxXfwYBl9aAmZ6sjude
FgZRob+8TT72frkWqygUjqPhPLZJriod4NBqc7l0NiQxqsIdDOEX9YwkzidjEPnb
ZuvBgHabwgRMHbQ6ixE9mxJMDKMGT/0Vnxov6PZSXtnWNvGbxnKHBwMUY0gvqgpp
sgzJuVGOFxXSgKSFWzIOV1qfYLXNGwbKvX7wYxfn/vDkZFJ9j4+lXmoVuqfjzjO4
5v77vekgQ5Y13gMTkqFKojVgPjj3caaGtMz1pTnJHdarIOy+JzeAC4dQzShX3OCg
CwYtTmNzsHfKCAXCyl+XeWXDIvbRtggeuLxOb0SukxBG87bxzFW4zfwy3VdTvxBS
bOMc507Ym3XKbfHM4MlcjipP9r80oDwQG0VfdT6PJzy64QgnkoJ742BfNzugS/7L
zj29CLslZYhFKsm0PSRh8kiqm7bVr6yFJIigaLo+kH3XEbxHhH1GafghyBTazR+a
DvCC919EM0gSJdJSl3Dl33kv7wJFAD0IzMxs3RvQeG+aLKNPwWjmaQeBXjP2z6Ly
AAk9nc+U2cYkob5Fl/PdoCIoLTaphf/sNZJ8qA2uXNc48lIJCUetEO+wTk2oM/7Q
Ub2JmqlpbH9TpwJN7SUsEK9fYvJGkPXrcOo3/LXFUX/JKO2MKQgXJ/3BH1DZKqOM
5txXDF0zs/Rpq+dRGZQ3uIWGL8l0lnVxpgpyw+qeuv+UUHWi9h84mcVoqMxlvPPA
YamUkiEzZGEu/d3HGyRBkBzqL4fyXoFQ1pPETRNwPOcC4tw4wt6V4hS2sWgdhElP
2wXHtfl0+Hh/+TI3YqBkX1pTweskcNCK9JpUGbV5HCkM69go+07gBFXAjZXp+teO
+kBQsyNEn1AxpC/n7CUMiUVfkUYLd5wSbsPLwMcUqUusVpAdF97cWd/FHs3cQ5N/
SSi4exzXVI3QNAXNLPh3IAa5aEpHONZNvsf10YeMwo2S0O1kJsf8h6++X6YZrz8P
4pj3DI0VvQd2IkxpqEWxCPiiGwr17wKyxMJbnAKZOdRixjtfdK6fT2txgJPRXSNm
hnJ9EfSMJlBvjty1ExaYSk5KZk6Kyqmk3lzSR9Z2OErgY9oLu8qIfSkkVk6XpL38
nl/9e5UigAjdyg91ozC5V3XFkQpwbmVHjYtUJhc7ggjaMZWvJxI491aGUYM2+dqM
mlH7m95a9Y2wvdqt5peJdpEK7uMvvi3Y2Ss3ErZjeXdF1afI8PDndnhztjv6WUaB
7+6pnutRRZGZU1BuGooPZBWp1efxKjRYvl9mLF64UltzbhNZ3RuCLOllzO/AWMxj
xTitpfE5HJVg3SaFleFV69hJQe26aOXPu+Mu+zRL4jLVv0xucWzyooe57WQD+xJV
Aa+0jpbG8zj0l5iJJEf/x10RSyc+txHm4NJTwQzizx+UXhwXjxZanFq0Ng4ziFAM
p2XZ9HlfajhNz+4HR119TSorERKBGg7mpFzmRuOTp8WiMaEAeAfMIkeqf0UAmU+3
r2yFvHOu+5ULAucBrVMIsnARVDjZNXGQwyYC3rC8IvbevkfHFVx3WrIiIHWfwdR0
3wPaSWpq0D4QagD9nD91IC04iT+qyqqfXiVvjSTKmthkDKvERthBgGs9ELiMx8aY
wU+qK83BirFHJhlC7VdF8x2vynbCpTR/soMR/8BHoUyy4FuGL0gKG/gAQKGB5fe0
iK1h7Pt/wqe3ifytfLadbohyohcCTI1K7Jir9FiooAscE7h0K07RljO2sl+J/jTx
aGoFLrcHt8ocr5KlFcUjZS66MYbZw4oWmY7NpuKJHHYwzBPh0P3nV31J+jP9i2H6
v2BCqB6IsKDKx0f1YG9Wp+mkiN0fp9GslKSngBXJThuv4/9RYSvFLB83Hk4HXTab
BTIPUZNBPdGFzyvgktG0dFHW96AIVkviShcfVIxrbEncsNGEOnrdzJigJtyekVZq
ACvUaC7AcQ744WbnRMgNlPCKlsjgOy/ewUPWArfXxk3ah9L3LTSkXdxmC3JIqmsS
/dfsX4XKaMgxC1rQr01F82WZYC1PEe/swtqc59mv7EBDiwbLGozG32Xh0Ho6ZWv8
r5euo321mVhHOqR+GIWrHD+jWfH7P1tWwFJ0rPso9bNQiRHt9WeLQh+226im8GCW
wB/Stwi0/HO/VoQFuXujHlxuGTvtAKfKWSkpFD4cAkIFdXAiwm0SkP+YcSrJXyGp
GQH5FPxfmutHt24a3B5WRQ4UAPOjBY1gLnCEQRyiC/rZ7JZyWxTLSdIQD3xqT+k8
6KYTrBUIhzhJ1IVnfqvbRgUolrysdDB5gV0Dkf+lIdUCRar4LgvOc2bGGZC4CXUI
W+stQ2C7tSTDvaTukIybOFmEuurhlA/O9rMhYJSRqUorP8LhEBN6vhF70zhcKWON
NjEYPzGr5q8TrBFSq6Odaq+Tyb1rEQa5tZQN1jK6Xgdy23IImzRT84DjmBbBXaCy
6AUDRaM+g9gUIOT+YFyefWJEXe9Pm1cqMKuxKXfIhDD2bUOY1ie6zKWORsVmBjZO
ssp0VlmekMHNKZRuN/zcJrGdTcr1Yz72T2+CThrfWZ3sRjt1XKTBMV/knh2sf7M0
pehKJA6VijqsUNMJQxrKiHgAM5DJRW0W4L1I44omHZdgDbKx931E3L5wG9MD+Mln
DjxYFl5Vd6jaWvXz+fI8GT1i88a59Tt3fjCj5yPMZU7eRCYK9weyYCBb1d9ZvSLf
F1MJLaFWIpPwXEn7Ueh7clATz4La6RUDZocXOuxu58Ejg6wI4U8lWxabI6CL+/1k
9v4fAROcc9e7J7qg/sWu0uBC2aq78dSchIRJIVu+771r+HefEqVx8pRX412S65nv
t716B0HUVOfGWhfeaSuNAWTEA+G+PIvjlgU5KmrR1ZRlS+f8xuEKFg/bKZq4mSDc
O+ofdgW9pyFeWXikTHEftPF93zj9OEguUXxXOUMRrpUCOIBSPSLQDm244AOzw0ux
hEjtd0c132ZXB14coIdrtRzTleTfgqfm4hmGDQDXz6lRPv7a4BGiXiPHQlhcn08v
3bGzGDj/UTRDewaPYteC+TK2WgUvcFaWk7TY+6tz5bx15064QrvmoNvaXw2Sf4he
gmE9HQeL4wbgpvU4jTp5F0cn005KPAN0FEWHhj4NLC1jzIc7zDOB+rnUp81NW8yB
he2xyzoZwrRdxIhtRZS8L/TNfirqPznzCxsF6z/n9ZUvwiE01jRc9UmR4cdExeHV
gjH0t7ZTrfGmcJnE3jxdrcZXa4YlonaYqsoZyJELpuZqJEzujeVWbfvBa2Jo+Z2O
+aaTM+8jsx0mKR65k4OmJ06Fm2L83LuRUfAFGTGOFYvUbVk+PEq7fLD1K/6Om/uf
g4zrYvPuD4yTpT/cjMFFeq90r5zjjT2mjuYE8CKcUhz84r4iqbUA8DRHR6GKCz4H
8QOHWp1SFXzbiRst9QcZkSjgV1FpQwgXC45gc+Vw3iVPtFisaIaNAIV5uAZprAw/
h5+SocBlEVIOAKjY3AkOQ2P7you89kQOIYFDk2II5bXM4dqupwymRHa4DoJzW8sH
yZMlrFXhbsFHhb1HqhVLbhRZxTIhe5Q44AyvOeFtJjqNNxsQrsyte/Gcq5bsOi+8
k6wIpA2zz87N06mSkmz+fwDK0qS2E8+zrWXAkJT/XFNokI4S+K335tcLmEkT02Pg
wbK7HhaKiIs6uXFvuwRmhhZ/c/XMhAU75VxIgxkNARt6oBieF75TTpx0Ot1l3CWl
QiOHpAthfqyL3kAPdjs8vSUbVHD2I5Q2FXKH3nXl11q4fU7/d0sIKFp3tbXCIN2P
Tsi8M3OTljMetlHeUGgx8nsk2zPK6Sw0QiVMcCz27odI89HPIO+txTM6yEhlhyq9
24TLxW8eIhmHWApge3zgoiZYtQ2ppDoedjxuM8BRFUfb2J7Mlr6nGEGAhkz0rQt3
fVULSMZBLBYSLKouIz0vz+jKpWvQOQ9icP8ntGskdgrPvmzEq5H05+1KASY//slt
3caP0gO+vdMXs4ZrhUgFbYIxL0M6kvL0791HDzJ1ScBUovn6HoXqgRQOEkO4/7h4
OZvIT03SM9Daz5UYHqXixFUvf+sd+hYzK0S76/SLIvmGTLELL77foXjD+rIC8GFB
N42wENQDVMZHnKFu/EbDoXWJ8Rxsogn48BsWWB5AQdv7TGqJtO2LeY7Fh6sSF+2l
MhNUOgJVDlPJmRib86S9AnZjKm5F2IWFp5mRPv06ltS46Qblt/msvq4VB6uGGN3Z
7YtOJX8MzBYbh6R//NM79x5LyBWGBwc8Zkv8RJQ7tETAnNPa5NRR6WHKu8/4xsN8
iT8MD66Rl/w1LdhpDbCQGTOIbw1s9Ge1GtGY9jg547TRqy5KydZdhupSjdc0Z86M
S28OqmreV9Z25McNtlcqZZt0Q6Qyr1hl9JJ1n9QIO4rdS3bEeOQpDbGg6odhF+P8
2QjAIcdCiCYHziWket4cnvFKtkX7YybqfXsSq8YlcqxOPYtay6XdmcdyEDVNaSxV
ypSNA3X6iEnkGVRKBqfm8AwVeFKqxin+OhpmuNR0ySzUBqfNEZkne0Il6nh+kcdm
TgJwi+m6POTSgFuis6axFEBws1/A++x1xNrj5uOuwmucm0BGeUysX1/Cdt8XARQM
1EnkFMJDW1mmP4M7+VJV8OhuXWrn+3UlCn/aEB23nSxfXS2rTw4rvY7sYLCSI3v6
+xz5GuCaF3UWKnOQRsLXzFlaRJ84YzpXXknG7+LJ7B0w0WsjmK/LRJRhrEs6WqNd
99ojWzcSmXI3NzI1xz+JUu0uQ2bnndlKYHjdGqL2Jf6PLAYZER6VHP1ePwPnaccP
5MKMgLQpBAUW4p1TQvcIpdV6rrcAY4POrphg3w2z7tlmhF53Mk7zwncbYMWq8MjL
7jhMRJ4x98M7nXzoFiIn2w9JM1OsNPffkjO8ERC6qLzH55X+QWaUG7m7andYGvSG
6/detMtLIYSmAhIv8EfAeezBPckp/eADiR4THJIvu9PKa+PYgMYoR7lRD6cnWvx4
M5FnX6kIvkSDtmF1LGbb1mKPOTxg+lDwJ5NmPfvGcPa0FP7roDzsr+wYBr1q3m05
0TKlkqE7QfvSDAYej4ZN3k3J87OV34RlPTVM+fxNO0NmRaS6hZZLOoF7YM+W+moR
xGFZacdw7kzIYF7d9CZF7BfGijXlRNpuD6oJ1I+2a08EQ+B14ZYWUZveZTHdrPBP
toDwu7j5jRD1qwKXGohvq/I3aHb7Zs2O/BOHWeGDYdclG9UHHSxxThPH/qSYH7Kl
wysiaKbo9zv7EOhO7JVpQMOC1HchlG7qVkH1X5s9CSgsfYvcIEAK4I5aBYbFHv7M
kTdE+uFBBsGUC+jt7vp7UIMULHia27WGCZlR1Kw81vNAHIsMJ6aJaPaeTg0HhDgq
xBavySS+3QjxHkGpvRwxWVe9TziP1QtF8WNFi+zeza+PEYGCLM4LsFYqPMzR67aV
qMR82bcL/0ygjuNk6mSQuclnqZzuSrg3RbdXfP8wkBujt6Pl0qJaKlNjpW+QjEfB
1HT3pFLBqyPj6AacswyW0uDupW+ddAfRa3cyqnSb4opBrbFTKlxbHb+W61sVU8ww
ke2JB+Iwo7nSj/xaDMM0e6+2ZNv9hQpgkLMK24YcghSYoc3O7PF8zv86fkhoi8el
nYMoqDpClqb5RN1EX/iDFTtcUM3RvpNo7lVS+4aEmSYqTyAzNs/GRMFxRXnpLam8
9uMBNAvt/IYm5/UitIyBF51ssyl2xKRFpj9CQnOohr5Lf52t7aSbHVIZm/u67L8r
XTphwgD1dw0VOTsn8HkruLwbT6h7EaYJYorBVFz/okkMRObaioss+0KAPUF0puaZ
Sv+EvxoHFFwrnPShNbJAfN/4XBo0kGJZmQNjH+rdvzreRafa3SkloNoiGLNPYPE5
fHJH5Sb1HWzac1rAKGYO4IwGUDY7EaIXIyCYaEpXYXVmHTgRo7gBVfSfRHZYEapV
k6Q+lZm3WxwAh/F6QHw0uA1W6bAJWpDCaCDS79LxhWUNei6sGs+72UIjYj016xE7
k+fYZEAa9QKAtRJD6SFZVWFbFnoBeIxbAVaYpA73xSci0mlkDYNuhLG1vK2YGt3+
e3EQ3i6Z8a8VW/uUkjbxMGlsOlCRUFmC78z9SgtePtLTzqK8x8lwYtTtUkoI4/dM
IYd8C4iQU3i6OXYRIL6GL84kS1xG65zgg2oHSIlypxVlcoAe3ShK2/YhBpwpM4gs
SnIaQ41KtP10oUzlpy7fHmhm+Rp3mdHIkLTmBNb6f2Aah8CzQJRHvM/2Smwhwnko
ww2IIhSZzh1GlDldmDrCdPWvCyYyUP9cx5LCngNlmw1ZrhDLdAhAli7X6cIRsMai
TmzFE3hBMZXk6bqrahsj3piL07JS9tvrXC6kNEB7gSxvJkLGjtjmihnbs+mtQuRW
ty52x9R0sMPyQPAuBgI3QMbp8M64AW9RUhyNGPj022WjnbGKLsoYRza0VEGVPWpZ
jSuSLonVdcbTLN05IR96oWLJbDFaqG0wFrrj68ZsC7i3RuRkzqoRCj9DyINamZO6
B6zsqSSAXs1jud7A+tBql6pPgUGb7GCCS/MUPc8Zw4vDnb6ukK5eyMHBouFLF+mr
MNPXYx0wQtB5PrRJqqSVDeJOxWCbYjC4hCmqTwliDUPPHo2QwM2oTrZOAklFhtat
fs49JFQuk3PH3Bsqg0FLQdsU20rpC1za7vuTyvVPpBuQh48D333t+EAIQr/kOJON
14kfrE43E1hzhL7UO+U7Lh1Qt/yLLJgxZYo1+8HbeiGrNpiJDzUGcbmS8lYYoXsb
Cz5UKYFeU0QfJg3Vk6z9BlXjG4S6uMliJuXuGjHMytxvmYZy6KCs/y6mSGsayf+O
EHGUN/gzWWMw4hcz0bpaSx4gE8G6ivd6ABbBa2yAADsC3D6Ofnb+Kv4Q4RqqE7l5
sctrUw3CRQye6Pqaf0MBdKAXsLQqgBmIF/t/DjmviKaLjARyMo9pzelxSAaD+kI9
RIuISOqsmcT0F8UebsdnMsnlYwh5MTtE+8susNYr+k0FOVXegLSpUg8zjfPfTWZs
cYV7VlK/2Sh4vUfeMlBUy/FGyKTI9uYdfG57ZVc2ezjkoPEUIWyEZ7PjCYaLCep3
TKrVZbob1GwDiXeIqX+PVdc5r7er6uynRxOHu/9bI/7q+8+KBbL2JwN1CcS9lzMk
JSXlpDVk2f+kPTZru3qpMzNY7x2ZxiesjOn+++4gGF2eDhizIqHkmSjYtE3ByG+s
Rn3rjvAR6cMnrUe58O6ROjaVCg+Qa1pTFqoD0y5aXHys/B66Hbq+HGHVEA+xls9R
vEOmVccxQJ3+x23uTq6BW0Im7rOG/q8BgFRZV2+vIubFTscr14JEwFLWkm9hs4qJ
j8dcNTC2bW5hLQGU2wxi1eTBUELGBTbDUrFkCuHGBMXlvWmG89B24N7ZfhiWFKFD
PFt4amZqD2Vx9TqY1Cnplrx2jPehTxJRVd2jHh/UQHU5uyC1omDW/0/8rZhhRSx6
68mdfKxQHen8xpwpM3rC+GLC86Cp9AbnuiqXGWdiCBaEsLFfR4hUk2Nhqrzmtgr+
YW1i9JEynKZkshulnZo2AZJUhTeybG/II0mHaO4KKdWgTGTeUzLlLwRi+OvdLJ9r
cPLRte38llUS+wB+2B4OMuZCFBmJvuEG3da/+nfPJRsI+mZovWmnomuU12JmUZ5X
tj4ugrZ+4uO91UUsnxlBrtXaqLAR8pErDhAOP29iR4/wB/wQnZywDCwfKIt3mLyD
VA9C37LSEJqIDFTL5cZKy+SjZQ/DZiigIdalWVrQbeJIEgAmGMQ5khfmOtwt7Roo
7w/FIZuLfSsC6LyfErrIMlgLzXJOkPup70vmCIJK99e+56WdDO9X22H6Cw7HTpxh
LSBt5rRp+5w43eZLnnRhO85HpQSUR+UUE5vQjPym8Jil0QMPPB+19jeGiVOe6Day
FsyvovbOjYNaxcLdTYKQzFnEGRfCgwGTgvluhAPI678RZX0yLUMvkUduB/RuZ9Z1
C/3032grDhUd5b5Pk2fLw5CGdh3TwE58kdgyz/NNUA09Ytu1uKw115BofA6epOP2
5HQNSeuubShUsfHCwXUTcHUgLnIOURAXPLyS6tQ58VJrNlF2EpsmewDHYwDwX7+N
Teo8GASDQzFvCwgOMDUFotuM0RzdFvDF4NdMz9csn7DxoOiyOfz6xUbu8y3t115K
YUZaEeBPhQm/P4g+1MUmyivMSfZEiHifG5iTrI5kEn7rGEGM8XNc0f2lKkPX3z96
PTH4I93w3ZlJsF1dUqx5M+lNOceGmOpBQ+f1wxyl4UZm92pYGqq/xWEjlLv4FbjM
n7ZxKWNTu9YtgFrN7MgAPYQ63uGiQPHNZVd07dl8+jEFRpqitxaDORz0y5R6BIsP
a3swWXj9Suig5xKriTy9FXmciEFffH9W4q6qQ7AQ48f9rfJcEAY7V0K9KwoLFNmH
T39GGp4l3jjM9iLcBXEme8KSRmkv0QYy06HMogDSt487VmYpFyz0fV82BhdX1D25
GkSkeHVfoYaFnV96EDDwYbDBVmGpYEAZFLJ9jQBDCPqmOpW+zWwpF77sjbdcZ52C
/MKwDNbcJccGSgzQhlRJ25f4dblkQxf3sAYNaJAGkLvHPaGefBYxOrjFwlSZ68eM
yeiyViM2hk+Dm36kE9TsD5NERFnGCeUzDsj23hpTUM8sOE9JzpQ4C5sVP1An0Y+P
UdcwKc0Srqk0mVbNUvfrV77ISE9HUX655jwDuIisd6rmVapcYERUESzh2HAYUF/L
3HXYXJEd6t7dp6IOP7jL0sz/oy/E8lwSKmA1PZsJYA5sTpkwTTDRBESGuNo3+9oT
jWfumvuVd8+/PrFP9QMnAfsqHltXgn4sOWUgymw0MyjPYHbhZkAYopjUQDlIj/s0
vvoHjOTQ522ra9iTPcUO2KRNFnpWB5rm30ao354qFXg8L4MK6VGo4AiHZwo6xnzM
IaWzj8TEPH7/N2ECkaTwr/0ut7mP7orbkoEGEs4C6zp3nFFXx6Ayjey6zBqOio3n
PpUHUnHKoUuDi1Kb4XIjoEcYMKToHNkefiKCa5OPAE1tN/yFDdoSNyAlA3dtOgqS
1kFo0nmmvuxVo1bXqSaabcnVHkeM1NLm5GSTXQflV0Sk6eyrag1DGwk+r7nnJxI+
zDpHMkKm0X4k14nhnEw/O8w1P0ESSfz9oXlxakKXVmoPDDL7tX8S8Hoo4n0u9ve7
4RXEJ+B36oaaOppwK58R4gRKxWyWaWvRWYtu2z0tY+x8w2tYuFi0uUUVsmt2LX5U
eQ++4Rp7JG6dVjp42clfR2hfTNB2tGTOzlSjX4QZFWD1OdvETmCrhuIuxsKxTBYb
OrtnlmWFidEG89Tdsdqxjaz6Q1zAwRIV1D4qicCBFSrvyyY00p3pf0kSvdsaG1lE
nYMvsVkmuGTodRjhCWbk81dqISshrRc2pThF8sQuVrsEC7N3izV/4yKhrgsjIHVO
GC39lxTJMM6D1Z991Gla2R7SvVmVpIPHfKTUQ8yAnNTnHXbuCM4KqY1al6ysHPOt
3ufAOw5dnohqm/EM70EwijyeEDOQqUVySlX6hBjXEo4d5Ni9qEFI66ziGMLbU+VW
QP9LiEC+uRlEOP27DazWG29LYd3d9aUDGNNMYzhTA+6QiVpzogRIfMikqZgnbPK3
fm9xh9s5bBpP5xVYEETjeIvhlGXthNpUnX2Rk5cO/nkEU2OfNA8aJNHqTR0PhTfz
0JIlV0TOq66YrrP5qgncL5b6i/4ocFLEHhrMDSGs8LZb1rCkC+lZC3Q2P2cH3dPu
hcBw4WNL9QPyKWUMmZ0KVnqifLE5DvRRmUr3AGaBnywg+SwYGDG38pMkO/r1rHsY
sEh8L62jo9FDf4YeQDv6PExCsRv3BSscjCGC0EhN5o9Rtu6/8q7R1PZMGCwHG0VM
2nvqwN4Buco81QpgAG4fpZKEX78Q1amIcUeWVC5RqyFJM6e/nxwWYLlrSinVU4IY
5Okq4Zw6y3EaZw5TNFdOHEhL6iGeqq3EEsLuLn3hZD+5CcputZtcYLINjK1H/4KO
cN3VT9pGfluXzhYkOFZCz+uNmDEcoHqhUgKQAgrPl665iF1C5QHatiki3KQ65ngj
t/1U9vVSJdwRTiqkXZGQLeWC+gcVtyK68Ua5t1sjbfYY3ioPWlos5+IFVgeVVTsN
WhXCcXthxg2foDESz6z2Q4FO7asp6pwnRVsT+0IXWXRr3H91CL6u4T18bpckJWbs
1tbRphO+UCN7sEBrMkX5z9xpn7FEkqvcLeBTd9XXqn54++Q1jqbfXKnAHhFSfc9Y
0iSgSS+Nq9B/5qWKY3yr4Y2snCFiumqeYNMUam1NbZqE6/AGiM+x2P4K4aYT3vuY
p7HBy76CFwsHKpHUFUJzZPHhDKJl4Hgu8HSs5gMPojLL8x5JnhHfM/jD+itMepf2
F66GNn7HqYz/ggtoy7AbOOH4zLVJFoX6P9xj8e1b60wQd8NKzw89Y8++4b1hORrP
bsC3pQ+XAFtflK7k1mnpBPEQ3/JCCxRLrCAuIg5Xq5cggoCyg3tXtzrQaJHc+UCO
p0ITRPoSLPVDxC/dyqaaege+bOvL18fDVAPecRoOEXmOPbIu5O5FhTv5vMTHSyGr
ZDNRxmmmtPecK55PihcaFFWu8ayI1V8Ly37Ex13ZGi1N9BzQY8sSYbuzayKEcmJW
/y4ZLCuDuqSCGXdHvtSy4LIQ9slZxe62rAfjC2BSCIrrNpSLcNHbH6c5f0Kddb9F
9OQEvYJ5vaP5+kPg8FmJf0DX/ZdmOwcscaUgAQp0iDbtv8P31e8QGzeDHONT9qtI
ZB8G8+5bD8w3tM78QT0VI6df6IhFk/RzA2PYM0fW/bNaxxL87VAEa4WaoaG3s0Rp
OBX6cX+ZjKQ8bi74bZISbEQ58izHT6U8rFnjS8y5U/ja8PirPoq6WAGoVQt1RfMn
ufGzTFXXq+OMoT66UuO8Cs1PTqWagGNFRNzGzus6dJUkRYbCVLc/uresQxJLy8I6
f+PIuPB+SuH258Y5puYPnjk1iD/dvgyryXSfKuq47Qs81jVC9et0EtkoY2v6tiIJ
CT+vXuwmLYtc6vp9itkseGD3aeQPxrYWtlNffzqfJMKM9LQKUkFTSkLsE8h1exL8
hSsjtgdeJI7jnJRXJphEKLsJt98yMEDw7y5aNBs35PyPNXnIsbIdQO/8pv+yuFRe
kaF9wOM2u96RDhuThR1bVvMiocrrijokN4I1W9oR6sm450ZaMZ1f7X4RTOgpmvnX
tCwZHa2+1bNLwGKsv6vh4lVyRbyIcbd2ZJQ6wX02EvSQo96GGGJNTMYip4vNm5CE
th/A1gcr4i2hgwszaQKQBt6eq7OpFS5U5U7Nzu3+S/ZEJrOKOQ94FVSmwz0FNo/P
89Es906YQxr6q6D2rSy+ZhZUNC9F8jLd/ltvs6pIbEm20ZLnc40WOG+IuUu70kls
QUuhIj9qGZj3RHztf8+pvafYXP8meN54lEUJgGkHb5k6AUFh54/lB3F9suPIHIep
E5yd33dvu+NZ0YXqtmZO52AXyV8QR3SAWYQLh6LXTFub5mnYTkyHLMQARyY7uX3P
N4mlxwknXSBN7ffhvyrtHZV5B8AvIldWS5DPy2iKMzaFXpkgpAkoNd4xmOJU/vuK
xjdF7KftFL5Xnl1M+XsRGcLT6907lA5qahT5JwT+7t9QboMQxakH4eb11X/tCQde
vjZPYahMyUUdqfY9kuEB6J6SKT9vXGmosPcR5WMHZEtWtTAA9m4wghIv8nUuSeQM
DUslb4DDPha3YOunjryfb9p9ai55EUfq+2C5BzScpxVi7hFn/HCSLG3yhWOItg9P
EiZ6cARcWQE+jkE3TlP+JM/N9aafEIy5aJe94HFzzW2T0AjdaWmiJlG5lE1UwMNd
sborFJigatFCLrDU1ONfBETcfsR/gHbABMgssaeGxLiJ06vcA0lhj+jpcQ6eUBgJ
TjKolke/QLZPLYjRuKsrKARE6LvimehpCTDmRZdFDv33p0yCO9W2IvtzQ6aWy/Io
N1TCZnU8h/48gXyUu/sBu0D9f0k+7TD4kxSHkpwpqzPNTOfNVuteCO73JBS+/Oth
6Y10aT5NZNPRJxFwkL/huh35ZjFhBajgG1g/qVjPdsmsPIG2PEhrKD+YI7kjER6F
8McQNm2mU2qsCKqdYgGGjph10tA6K6MFbOGFZl3uoxzeBCJeAePBTFdJw/dH2ArO
UkRIk3l8x5AO+ptyN+5HDqY1mKD+U1xmnk0DyfttS9asdLqPWf7jFjq7QubLk9D+
w2kppQvFijLYQdDJ8GW/d7SuwfCgwS4iCrSmNnnRumJeqRzZHqqJp59WwxmrRrly
KRZfE6J5gzaCgEDVLkJy8UfvW/s8CG4myxzTDunLlUGk75fJKw6A7nsnECgvUimy
AN5HnPkwoqw5Q9w52pu68HJx6WD5Jr7luvUHtuATQR6rDpjhKV1XluB5m20rgHHO
otJ0l6tE0jMlbmdzKw/BGyfkX8S5nZr7y2/e340wOgRB5bCF3AaZoBPHMUhD5Lnt
ElMM7FTygCJEbnwlPP0UNFsjaoFGpnI//iCLeISRdHgzYX0Qg4JzSsQ1OlhSH3TU
zP05ui0O87YRNPnAgNTn5z9TInE9dc8TZ2SU5CIB9YbmtDFiPQNwPbJjJJ8HKahC
J51uBWmxUf1V5qUN30llgl/FUpeWyY2syl6Lltomy4Q7pBMfxYLVMaGo5ibASweq
WrD9pi/I1jomkHICY9zgMco+f8VYF5mguIJYscCFa2H6Hqg+GufTZsO1xEVzfsNw
3w9uKA9ZNMxuv+jcHV0eFZwqvV7hPZN0EjSsdFcEK2H8sF+wTHnotLyX1StUopwR
qu1cBRcRDaLVhxGRqCZw/g08ygOtXdZwA5CNriQ2lWHLAXXrg4oB3jSdEG5jhs+y
jUJ3G+MmXdkGCOvpXEh41q/3+mAVYEZ5MOYrAiVZ0OZjpEX25mf5Ap8jy1QJMoRO
/vbCOsGHz2fJ/G5Iz/RkWA85VmIMqsneN+V26ljLuvEzIRx78yZzBUwAbznmz8yc
Qak0xljY1xFswezg5yeXM2Kaqus6S+FG4UZmwStU7KKXT72diGNjVNGbxBO4DmaL
DlClPp6Z8umXCBG6LK3G/xQwrjVibpxWSE7vwzBAX7uJU+bq+1APvAAvlytvpszz
+XGwdVWVP42okYzsV1cGVbEBI6ckJFg4yBLg9qL+b7tUS93JO4FOX9Jyafa3EBsa
QGhn7b0aOvu1riEbWfKpCDG5P2oNqTafkk9CDyCJMC5O4CqnP69F2ovHuaN2aumx
r+QWP3goeOAWZji4fbLXk7wugSfR3C/EklG2SuBH1ENc8Ns7CIxYSe11ZtgpoIBM
mk6VONs+VXrNBEEhTsXbUOBMK4azdlm0ugl9YH61gkVvhdiZSeoF1cU7KOykbA5I
0Njdq2lzgH2K0xo4oVSE5DBun53wxStyOfuU9MMnNICEKldvSFll1HeAEcrvpGEy
Dbu0loDT6sVYMrD467MbyjTH9Xq0JnXtnSchewGQtlymz5BojssJhYhDuw180GRB
9tHGTJFQkLzXw9w3Hdyug04VuvHEQKxc/6o9xUKBoM2gCIdoSnn+mSkk57whXeFl
PnKYO8qAsGMZr0FEOHozY3Twnu2ORisX4axICeW3qvy2zJNWk+aWQ0Il/2DHJfDj
QHxxY9X68NS+rAZHEzi2QIA+9Srrh5urIb+qY79Sy258W8O0WcPUud3+dBoL77gh
t1ZeoATNV3JEnogVvZKFO7qqDQCWMXfIkBGyxV7/DbMVvm28bFARx+WGTvuAKrgQ
5L4F6RfWHsCR/aPy21k01vwfxAjnJF26kiqJJa859zNBpT4SDiL3mRgTtynq0gmt
fErktSiZSmQGIPbfaYwqCb15EERH5SHo3OUVgeYouDb+onlkIyqgOenzVwgCTubL
d/WTfw6OlH6SjOSYkSA+E2DtMAr4Fc1u2KMkNrInsNCQ6rmcB7WeCIuErk7mypxj
vCZsscAX2KgfB7A9bmi8MFZq9ZehtTxR81SKAJoXAdcfYSQmE1MA2JsCIg82U/is
rr1xigP5SIYmVx4FTy9eC8nL65XMDo4zib87jScwepSu4rh/7F5u8KoBhL/pGGvS
sywcTL/qaKMrBYjgrGdg0Bh0nR4dr8zAkJyHa8N8QIwJR/9tT6H3MMVfZXZ0IzD1
Zf+9VotcGQDaXbwvi8UMoacccurXcjvwh3a/vI+oXKM3lkMpYDikiqFmSgadwRXS
cV8MRyHQY6xsTRgdP17bBeis+ln/2iv0R3/TQRsghfEH7tzooP8AjtpkT3S+C1qi
3PbB+e53uhQjXoQNYgr3/VnaYLuy5Kl5YOk3qEgTwpJEeru5W5VSd/gQmJGVr8P9
J98Z3gX+/0IpXIsPsBdAj4o/TGsufribbyJ5Jv25v8Fn/W24B2G+ZDf/2ftStsYq
yO5n9xfTPrNmvAmHg2zhO4Xgi9ClmoLQ9udxu6yqfo1N/f/UcMNaZIORCIEj4jcz
LLja6M/E8zAFMZpO4Yab8FCAefgjOSNM8ulF3LP07cnqxSe+ZxSDtwCHWFHr1196
O50YZck6/jjoAGMluVs6IRe5ILXMzTFlZWug+Xv+2m+iiVUtaen7o0kbzjmUuWTe
WhoZOo8oBkKtjHK2bK3F1b3mrFkIE4r9rZgW79rYQdGAZZ9shPJf2dodvVKEIjgu
mMgNeL9VLYd4gITkSPxj48O36wzPZLS89agHW6FLzCDPG52u7Lj5uBBm3p1irHDN
qhV449Ak+itWoogPnBiQgAcN7U3//0hdwGvfrn2pW6vx1FNluRfS9pJ8RWr9tWBF
9wTMfMKKdX6qH+FGYB+5WCsxgRDXYDzDAhLi01bB30Dk2qZ/I4nkuP/8sg9fI1VZ
6OqOnIFqz5I9GHjR4ImSBlntQs3JQMuVHj0Wffcgh7SWC8nUNFAKlQcdwSsdCf5U
+d5UOBslTO32eRRYpTazrytwozLng2Soy67EiBHBuAPwlZquIiflzlO9SK+t3W6E
UT7nC675ad5VpDMJj66AexP7wgB1vRWfrlnd86PijPGZ5GiJOwBAUuVo2AcPz0WU
DBcGeebjTcMr9Mvmu39PPatCMG3zCoP2BCjfR1+OMHmqAbzT0PiMvz5flYPnBF/r
cqV+aRcbivx83fy2fE/UCLdG6V4ZK2JB7/Y7E2n/Pcs7Ep/aIXygqELWjC1BMGz9
eSnVPFXBkWokDchYRc3nRPw7WWu2k+KfpyER2UxPmecIaSVR/tnlTa+m9mcXvTUw
T+y18aHyEUTBtTnqEGH9cAfhnchAFJY1bkJAfC1Qe31qdAOjmKBiBQmGpXc1X3+g
4vUW/El3w7CtReMmREPCyqJTd0Lzn15Y55VRQTpV6xY2KJQzSOW1z/VQ3+6hHHuC
HHFQlyNdmnM4e2+HaMGZHZXLvPo1hXO2CoEXZ6leY6j9Lt1t52DXeh1yq/Npq2R3
bajoWAsGBbLl9NxIsASrZaNrtZ4+V9jrfs5Rr2s2QKTEAo76Lw3Jmgc2uEHEkXBV
28znwkKHdHg5toCsMxpr7wZdLZsghDFpviDTmyPQU+m4DDUNnD8milqEM3d4dA8+
gzT8KCfQrFjtA0iLCZSPKWjAo16z0tS2SMCkceY7RKvUy/hA3OYQybxzAzQn5EpD
yi9VgabZjQa463pqKuRojG6rnVdSKJ+fBoXl0+/FcmSl7qP8BRCBtWV2CL9sRtLv
0t9S66mBCygBKk32HBpYeGSAOa5FXqqpq1HTm312bmgRtOxXHe7Lqo1Cmg24QYkT
r0knMEjzE655GEw74ronhFkZ7s1z9FXhS+KNynzedN81Y+Ax7HDTZh30n4rG0Spt
57ktTT48CQTsWAy6bpwHyJC/4mm/6r2h7DWG0pbwl9MSJxH8I3lUw+HwfRC9AMGI
JwaHKtvLVB7DRCtepOoTTyrlB8TS5YW6xLMVh2VK1aUdu4bPfVbWDbYZ517h67NK
BTG7VkRcHTFJa3A/L5NJ1Sl+Ppd6vk9mS0RJltyPkp6rdzFKwEmcxPJY+rsWKdZ1
lbwCyrIZ12w7C+sc3kLf9KlHs+0DRNnSFb+Rc2HgNmt2ifCh5dq0JOmf4MXtZNIg
7YkXsKue6KbnrK00xBUqB1yjUlJCSmZFBepGf1myMXs+ol+XwI4CiF1ov2Pzfc22
Sf+yvZdoZOFYds/R0KSXwKeujKvmBycc7Le9n/pZbZcdZBO6CUQgWKn4zKZVuu4H
ErE+y15BUNbPYU1uZnm2UflGICtl/MiFfSiA9+VCnsQlRc2U+5ZcKffyeJyZxSWi
Gu77ge7XFOvJam7g8KeYCKf0VVm3Lo84nJ/TU24GQlUE23i3Qz6umG5EuLDmsRSx
FcwfdBWOuzcj2ecYMxE01HNRvbnQq3UAAbQN0msdmb0hUEQwytwcJFv2cFXrOh+n
lXN6WTpCpuuxaCh6Xb4ZAhFHn/PC0hEO3vZCcvVFaF4Mh6pByy1Z8O+zIj4lkCj+
CjrN3lwO1AT17z9sd0snbnnl2XtTM59AAOa+DP/HSCsbKEUlXWrZ4uwOgioBzaOZ
fWNiin1qLObobWYHQDQqS0nFpeTl+bvY0nmZVp5hUCC5jlFPrrzX8s3AKJUqSqGS
mQZceOlxakivac2ynM+oEI4aICKuR0uF86ck+djCD8wUTKA509t0yd9kFqe2JlPm
Hli0kYTprJ6IBtxrgrqs6GVkwlwfJBLZwEYcie8f2yCabtn/4PZMyGuEJhTsKul7
m0Ds07K93KsCy8VqHPD9eMGKksOXLxl04NzRiqvfyBXc+qGMQGs5gYUgr0ItaU+4
SPMDMHHNuKppbc4LkXis3pYIQMKzH3iVIAR3SSydGPRs++Oetd+RdV4VW/tTbgDZ
/dnLnkV5ANsnQAcwKFmNh2Y2af2BaeJECtU6QhK84JVxzjMlMBy0xWA1fVjuLCpR
CeeNOsI18JnlOUabw+oFFPpN3X+YU790r/WGWqRPVOWF4CK7MMDeUQ4dQt2PZQWA
4KHjoBuUXPlMuNJHgwqQC/dGDLHqcxM5fcK7ts5pqIfmfsZeNXYvEAqM59LR/wCO
g85YWuu4oU8YWnAAqcaMQiDG+0MRuK7I9hQ7HoN1PdRCI5bqlZE7fCqu+U2oHG4J
M+Etb8alHb6yuzcFIVqjo2VJYO4toHHsGC118NP8UMAJcTMzo8ZeSuY7Z/t8a5qh
33lK2n550qVKRn49znH7soK0Clm2YYgkS3D/Yu0iQ2RhDL68K+agVWJBB2oupH8t
eJxoePicsXmymIxW1Fm13vTgHGVC3NxW13T3GtmGHLg/68Hbz6pw5fmIrWq53ahd
yJZ3IXnagivb8ii5N0T5fktqfyt0OJnDujwlTlZ1Mj+0VFbmKhi+18LxYbOfGMlE
DV6gICGyiM1sb2MjvEzqj317EdN/V38wTD9fDyrHCINMynYetJ/VdTIE4/HBaCB8
Kec2ROrjzv+jBTk+qrZe4/Q8JoFV6LNxLnUFPd/jNhmKsWPLjS5+Yn7q37rX0jIz
eRjA5pm68YW40NWCpvrqBtLA8rhh0geGjjPx415rXKnSJBifho1Fsgt46ecwYvmC
nrFNw7AYK4TqLvYhdY+p254KMdED9NkRudjolRhRrW2IsRCFEdQWBFiTAeNXWHaI
XeTqQRnMw0DUQmEgiyA0rB+G6gu2KGhbAjFkSR7Iihyg43ydvrxEwcEfanVU4xwM
l10FSaPlmwbNrYzaQX0qMKwiYqZZMCBRCdVRhuHwLt4AYa+qXIpqlhx5HZrkQ+Ro
Bx+LwGUaHjBsGKxnMfqdLiKoR0pT30hyT4Ys9UD0TzSnPX0NQzjmQVDXILqamp4F
8N3eUT9Kl6w4tEwRbUZ0q52e49zYkgFRab1xjFWsADOOTJOt+EfYfzJXfw9hmqar
3LEJRtNlf5yzsI6iwQlZziwYGW7cTTGayn/TAYPSwGYFZ+NZ2egE6WrNthsEG7hA
prcMUIQCtrF6L7qCFRdxdCp2rfEalXOY1Z2GAAWBIhRTTJd5Zui+DKwrqUr4BYAc
YVSFov47mXeV0udQoxtgTkd2A6c6TxLvNEM8/cPVzWhHe/dldCX8JGohLB/elA9m
TeEDqiIdlVSHAcnR8gvvLUVqOpp8B2LjMJ/Pvbhpg/1edj2D41COjUYbGStHvYw+
80LZ1sz79et+sXXkmk2QQkbg0l5UUqPdFLGh1iz916H8e72EhzHncFBOqBNMr2nM
LfNWKwavkachvV+Gpv/XWmuh9EtoVLxwkx46uF5VtpGS2gwPswZBTVTMsfas/lTI
yB3/AHhCWi6Zs7ytsPXaBxkPVaOUdbC1j6YtfU2u/GYjnXeDxgyuGSI7+F9TL8QY
kbcSouWNxjYhCY+Ag2GdqXH8EmUA6JO75QgRSbgKrPCX5l/is08P62jHySP1IEL8
3c8agD3NbjdSnIeFzvNmx8OpnCziIvt99h8nzuueIPQZTMPdz/Rk5E6HwLEJGmra
dc82OGI4h02sl7ysN83jtot5bsESaLLGAF5txMvraNWQ3QP+0dM4aXyrBqJHZ9mR
3aRNo1Bzivw60K6/e2vS34AIgRhv3m/bHfLJPGjRm0CEozGOsYPsAfj7UGL24txW
pxxPj3v1nUnnGtaNpqpA+LKbqw1mSO6gjeYni3YDf97a3WpWS6CBzT3WiGkKQVa2
1CESKiGsmKFyu+5x30VI3cLdZH2rHqgpAerOZRYkGp9PrV0Wzb0Nu4CE/YS5SHtW
fwtoYueeUTVhZaj9rMPfD8/xUemi+4YOSkOYyhGI2t9l0q9Wtj9YOExIfvoaEq09
RNh9UACcgIThYWmWOZ9b/27XyM2iXJr0iOOS0lYO/vvgjMxTxdi1s4U86FXOX/B3
oWregTR3Nhkfo3/DUXDM9C5I6FKndrmagTxx+hDHUwopoJhnLe0RgPjlSkBc15KD
6TvVYykBKffqUqJLIMqnzSNbGIm3HADtNE1HcmU5WHK72VBoZ+Ppu+QbjrmGLM4o
1HXSNmstXG2xt3tT10XaTnmXzeg7zJ0skN+VD0cLY8wZyyWbD5TwyH4W1ok6pHEG
9mafGTltKi1cQT6IqI3lHS2EGThTjfBCVIvqtjhzl7rVFkLytmnfkEn/cufhCtMm
hFY+oGvMNsm9tOdPnU9hROo5PvfZelDI7/csMNj2hwWTWAkh9cPWSSEKfuZwMfcJ
y5ZNhdnEuFSUcftKcC5odfcqcsW2Qnjcx+B3D6McnwcNpRVcdVz3zVI3nwI2tGHd
T6R+KroQ7aqvWeMGlsgfL8RXTbHa/Vv0BsELjKaG0dwqJCWZDjP07NotHesr9pzy
NtdgarRcJnYSq1W8K/5qQr8ZrdYXCN7JaRZD5Vm6GnBhrChdijJakAzZ31XMw5PX
XOokNuyIvUrrjVbOUKjxbFsYeEKV6ygLeTMgo0I3+MEECNXhnMEdjL3BwAzEcZZ1
tq6xla12bM+D0+B4G1R+QIJTqu/z6uiCFkV7PBwYVjoatewNZj/tNL70oNu7L24u
0LQztUrG6qictlLGMEOnC+cBV1fjkL1f9ebmUd84MM+narg41rXb7z/8dJ6YqpHH
tJgo8PGKcZjAl6fbBtBbivuIzhKmSJ1FGD7ibjVusFEG60wOR8zyf4dbAuS7iKfP
7eLWWlAYmK2OFB3DKIL1C8QuqLRgeWjyFCMZZPYYjBNalMV2aixlB7ouksM1l7Tf
C5kpWdcSERm8Y95N9yyAygCwsdr6WBFZuk7p4/t/3CYCu+Pwr6YhLnk/fwUnM44M
PJf3VU3qftxDwAZvnuX83pOvMFPYOdsZxqAdIcQBAbxMnyXg3Bvw/h4zRPixkJb/
/P6lX8UddX2FDDUEPJlc5Q1CGh8AY0PTK5fm/mH9B/jwgNJ4sL6ZsR8lns2qNL0Z
lrcxEFhZMTWgOlCX7taEM9wBhVMcNFO9jQCo4uu3epML3XwRpmozNmFXyXGA43Sr
3XfjwmWYQCpi/r/sx9kuMX+HX48pRl0A+WYa0bxTIvrCvYcRjbr0XVboTMUDYpVR
VFd2JCAExkO82kAq7jk+jR4nIKiirG/Cqhk45ggi/JH4j+tXkY3JY7jArxaAHs/m
4efpyA1fUyyJ0spdlr4m6Dp8vOla0sbfjwIOOc1LSPjh6dxLvg166OPmNPnUK4gR
38SXOvGb+QyIvmgnmGWKGG8jq10HQ2D4wb1XBeErlWx+H9zYM/YkOmdx0AmTbOe/
y8/lrmcFKUTx2A1Bd9HrMpe9qoyAskYbcsJJtVoRo2/T7178bE+w8HaHACtWzz/B
Tm15Aww2SYDtAwJss1czDZGevSgoVv/8e8d9KsVF1mSvZqMENQmHMJfXm14DkmM+
4WDB5rAW5tzFPEa2/zehuRCnVM9YfjqQjcVKEgTcZQG6VWLAMmdRXIeh6J3ZpArb
zkhjQ6FMEQ8hMCoY6UmHtczvOmVBRpSBRanNmK5u50buzUpytcLtOBroudfjQpUm
7O7xZluDhwAqhwOM168R6lO6Qp8pgyjF5rcq9Qefdrvl3EdqvxeSndAjj4asUw71
Urc7VXi/ILBPuZNYApGWUfMP2YDgfbdDjZG63Z37OTGPQS0bfduB+NSz1sYA7Wh5
uDEfPisdjBFVakw0kz1QafbDXh+G276fkoCTkoexxJj9qUkOcqbXeIZfrkArq5Ob
ee/9e4Gbkx0Am7qp062LTu+RTZePjcKuUzZDHnIAhDAebD3lgnGD6oF2lHsF7xcL
Y+3bxaI9f1oisrTMnFt0x9tAIq4AKe1XMm+uuIHJ5us3XVP1ju+rSOFl57U5abNg
E0AEN961homupwE/mYrvpDRmseB5fvqJEUVt3JctlXw1UC+Sgo8dIkFXxBoULvPp
HqZH+KC/Q3H9fUpvOVg+AOhRo+GlgfJstgs6wDJ7Vh16R06kUdjqZ3qRkYVDda0a
8Op+d2Gy1B4pltpBZDFOPUMdyhaObkZ8glauyUV9PJd7/eMdFwrRTkpVIax28K52
1/2F4HVSxdJ9H5EZLFaI4dDKg2fQ3l+ziza7klQM8W+wRbvB07yKvjcYEc6wdXg2
N3nwwjcP4EUqrLXHT5KEXR+f20PQz9l8WGhfeWO9xwiqdMbq/REKS4h6Bo8jX3JN
WsXSOd8Q98dawnvcIRG0WNVBetW6vrikOKriqhO6axudydxVni1uGAWintCZTqNG
01nmdXN0anUJXZZtRwKXJ5DXVlF00iYIqpoV6vbNxMnHUWPEq/HjDd8MrlSCWtKz
2Jzz7vPQkTSOJX/LTAJdWsOynGYsE5X5c01WwSVSnVpJ7JQ94QrGEDXno0DGiLgo
DADfiaWsyiUoMfHUAPyeIqzNx3b6afcz6q5sRrdQp6zTuCI2S1TDqJFpDG5BCecb
TShdAItKxwALzPDLuXYuaWX26Diu6ZwzIWRerh8+zTbnlNC4uzbH98vImJziua7C
iMyxx6IpthrKVPWMqWTmFD+7JnmbHv8te5nHqx0duFCKRlvVm+E5HVACIEWnb8ZP
+yADnUVHnnybXJeHz5SFvgaPWXb88dlgLezlguQl9hKq3EJcpW+AaTRZGLT7dFKH
s6SZcSi3Dl/fIlz256b7Xju1VrBb9Ya8GxSsB4SCdCO8al3ewvs7psKBu5Fkm8fz
/JgybbXgPyPk38bczHXMFEwzVCmOitpSrK17P3fegDquaByLiJMVhcAiqHDwPl7f
TnYp7WuZP+ot/bmfa5uWG1OCanz0Ws2sWpdPkVhW4KExrIbH7nYt0k+io4VkjGYb
gqezIjB1mfNcB4+rld2yH++jw0KNGBhCIq6z36CvWLmYQmhfcp3WIJK4GK/ymjA1
rY7sEgGuzHvdjglcHyE/MkrvpVN6qr5HV59xfVO57283YVNPXORFjNKKTEFvNAGZ
x7MLwsQFQlw072+oHUBCZdMHPjIAshAHgU0zDAifuP/uOj5CV3hFcMLu2bletUkE
pPy6DSNnjUmB66ehwQr+LnGQ6n7lo4zoU2rOH46DvZAEea5F13f2GcaSR2+1Eir5
Ndzf0vLCE/fSMprxE/jLZywRENGDEwcO/JieeWOlR+jP4rZvaGSU4g8sXVZUEH9J
490VzqplJoin/sJvKhmVivstRH754vv9DyBwgaR1whXx2VW5EvNb65Bp+0fpDqbI
9M53rwzyofI5WSefD6cOmCwbKwPqzsCJpfL63lydNw39YPLS1BsZaEVdIY0WbuIw
YO+p5Q6iqYvKq4+dQxg4cQA4dVq5Yw21f5690JhfyVFapk19ZicvQGrjkiY2KsYo
nY7uultTYU50bFK7m0SXm6QBuYsgoUdD7M4keRjVY0guo3YRG1Ad8116wY3y02kC
BmXoLvK6malGeTChSqL/yVvftqFL6Q9dYxTqn4QiUSwfencSQLFRw0Eb263soCbJ
mhxVJiHuRpJgcw9i43LZyNpxmSUTZQleFQXadNNsaUhMoJIWzKDK8citlmacsi09
7phJZAb2YWEsXW/iiAa1eV9Jp1Xu5MXhbABkx4lMGHbLrhdUBMaefrt2EzllklWG
VUqe6D59ZYFMKNgJJToAck6/+COMP5IlA77yn6/R0YIhMojjButw4gPgwP2AwkH5
RGPCwUoIyXpYSj6AhfL3Pg5JDBy+PMf4asRu60HfD8/uLur9O0FjMvbOoMyiF2CQ
QQwXorpcj5TUQS4Vy3iYlFhGij+PJt/wgYusOhAU6grZd6w1Q0OWeSrZvAg7vCO9
EfpWDHu1Z8ibTS4l66Lw6vcMSstyKW2aUQUIqW5QjN4Izyh8qAS6cX2kYa1q3txJ
08cSoGJlD2+L5H6zP7eUGNM1RDYpHj5VWaTSLin0EupVpqsSbn2GktqOeSyQ/qIM
REmnGiTBsk00jqEoT7uhfAmotPtRmD9iy2ncZrE+PoEpKFbw77fxhN5wEY62oydo
YORG0a0qKP71Vx18jHTWiZMwutrHQEWmAPG5leJNXigJRPQ8XbiKcOH10YZNuxx7
TYVlbRFuOdNv/o8gPlBLDc0C+WihuYZQ9toFfNx9nUqSIjqIeRgQWHxzKHuV4GDp
SfUBiT4jFjDUx3aetdwvy51JMFv7m83ELmroISsnLODGjMb/J1XXRi0PCDv4K0Qt
w7v0xYsnqqlKf7Nnm+OVJgtKsW6l1z6Znc2wA9ykhlcZj2eq98QumKNXw7WXQ4Ma
EwfmUge32iGxkwMtP6HQXvrVvzK9erUVZ+9Lc6wfKP67/rEgNwGl2+wZxVBQdT7d
MpLovXwXcT1/bx29KZwbEiuLKT8AQYR93bsjJzW8BUyJnk+EfkF7sGMG7DTLihhT
TqinE6aA2EtbiYPaRfipb4fpYZBwy2z5pmkpR7viRmONbwmuRecUxCNnGRNrSJog
DtbgWtduVtkTtfzBBNFtiRrE8EMSEAOC4rCzjZAGldMIjrN2Q5KnJi7FzA7M1Jsm
sNBUzbC1Vj7z92eTsw8CBW6OGH+0w1Em5HmGkhe9e82YRdvnd3JttQeeeSVEev6W
QEHFM4sDZknZ7t/JSZBVc9ictrmF9S2i5zrdWEecozfPg3XSl0qnuJ9uO/FMzaSZ
idZ5woue7N6f+eXzx9MWCipwZi2yDu532QN7qfaK/Gyt5w263sdtL1NH1I+TC6Do
7v54JbAgJR1Tg6OgDz9+XxsoZWzipruzFmpm3Y9SwYR1zKEd54x7+6Elhz9Fh0HJ
9d6vAwnp2WSUpDif0Yy/IjFj7E+aqOfI7//8bqgg+QiJE9KuoF76eAxoiHVPGf7J
3am+j8Int553cNG4Jcai/2LIQDuBxjmbNQrIYzFFm6ncUQzNT5j8lXIFb7V3k4A7
lQCNOglfxQ0hN1vgS1JFz5j5+EJBW9JC7/mFTn8CyGxkHwgVPfvsLATHP+SdKQYF
qcTJ2KbFV+96+mZbKLj+PVpNDx9omJvHWSmO5IiFwCz4mIIzLENj89GwWyYfcUDA
tSRJp0dhflUmSbh4+a/NiBlfirUEA0CC+vRMVQXETZRN9ooethhBc05gMkDa58Pi
Agqz+SXC5FZylySF/B6zRjPp99a6EqXJ6S2jTBxcKgBgbkXtaOnTMYk065HJn3DB
XKleHHuxCEIZTtzToNIVbL5SJwm2KI1Cqy53N7k4zqP6O56H58lSPvOY0pEYcx/8
v+srzQsvSl9zxCUfbXrBw3r49sjn1sC08zrtS4GvD4fWZnVO1aNMRrlcCes3ZaET
SXwm2LhnkklSsI2aTcg2Xa6vHz9/hDw4bBBsY7v3TsW1ZnEzhe+7FcCEx6n3SorW
NKdskWi4aZUBSUuPuNg4bYf0MyzGlCkU4STPWX3DA4VCkfxry5i4b0a8Lz5RPs/C
KbQuy3U0qXXOh5EjG41SR1Xqb24jQM2BxQOBGkEjAJgIZ/j91CvV6UBJfwD89Awv
ufw9mcQBvFFB5bFmcO5sU1FrKQAIzf4jplrd5++cq5bpM545zJ3HfMmsw09RAu7k
aq1HdV5lPDijt1pn2fTYY425faOXyxcEfU5T8ObruP8xRacaOvkzPJnam9/XHhL8
CQ1o50tU9s0Zd8ujUSINkSeP3kVJsMbTNLUGUubCEwmjAvPh9morJUmUbQophOS6
AKndA52CZSFL/ClcjxPVUKsPOBQ79xRjIhESDA9CVRpGJdQz9xJuChHQr5Fn3k4J
ndJzH7GL3TW8e0IZFBDhH1eViQpiL/zAxm7fO0RhzuyGU410Dgr6W6Zyx+FxFwSs
LTIQ2OvS6ZZS/CzvEnOeKg7simRG9AxRuFSs6Ncft/Nwbk1KIPO+V6UE3CEQ/Dv7
vwlpXRXsnvRPaLGy6B1bUDZBVpb9UbqfaKf0Rz3zZjhZOv0gXwXZaVehbS07Y4Yf
c4K+BivcLJdiS+X1mYXDQLp4DqyDd33+ILq/bKKmneVyHKJJH8MFRbDmJ/laf0pL
nf4TNGxWBj+lVRnX76Ok4Ndv7MDrMfHnJaivsaACseVsn/Se+33OPbOWTW6nDHCq
YNJvMRPgwl/5HdzYyCM6RaMRNqYMOnwgS62cFYiLSCjWgg600Fs8T++U/ET7OZHy
0aRxPlPy+48Ay+Y6H+/07uAteGE0jpbKg0vvyydFNcvrPB3K6iKxIJNyHmdS+ZBE
aM+C28U+kRFvdXWXEOjpezsA2Ee78n04zBf8HEc8IsK1MKBBoZzTDiqdHKNqYiSL
hEKnQ1uMcv+Cr65gDkwBZViIVa5lyrT7o/B1I4N7mExnC3VXA3oSNvjNTYLomfNU
a82v4H0IiOxAKtE/wssYY3gH0qxZd77ReHRG+TsrqKt8kZNiTv1kMvKBUUPLWynW
mYwpWu7Z/MomttDT8VfMnkssUo8TAGRJT5BNDzlBiQ5Dgyvq0QkeLODfwtOZ3s8k
uW5Cgk+a6dSJgeHeqe0b+o7Y8of1EL2KGYpbWltAsBjPa7BSdzYDADmIkE1uIwst
XSf+cB3mhfP6wQA9oMlsWSsRkz3UT6d8JMZOLuWtORf9AMLRRq1HMxbPQrNLVP+g
z1gTRrEeZo1Q7cylLiYFTiGppVu4UgjvsGeQR8yE0ahC1SLL57FdIrv3BY9FYLP+
qy1hueMCdNMdBbaVVvn9ALzw6oErhMIUThr6yO3v6DAx93bddfIASe+RaZFod4jl
+MK0dB7MjLWhAZ0SxkEVEDMdjJC6Dl4CgmHeTjSDegzNnpTueKTVBmy+RlT/DJNR
dS/Q8kYAITFUrZoJhfaaPHCDnb2bp483tAsKQDJEh+LEhPd81hJiKMO2Al23cz00
DLAgobnBeKbsESol9FJc9+NmI+32X1JYASTDd7jwnAfoHhCB6+wyaW3yjYyJF3aD
2Ti+jDK5w2EVHrnAO32Wraj0JPpw8CER+ocTJVk9s8CuE+Y8vcrV/9rwdNdCeGSZ
ahVRoD+j1i4orcQcWL+dEccIfL24mEglnp/9lL+opvCwemr+6hFVFWMf5/XpuIKs
0THLGo0sRM14ZfOkpP/nFFSWAjIT6atxyTBMQa8GzYEAa07HdZBOv6njKS8sB9WB
ZQNjeiByNZdAHRRX9OvwuvfVrd8GGR2m/5oOa4co4HLJcSuzXa68sy5vtveIyMCX
1rF/UkiGfpAlu6CjJc51izRHzZDRtLmpQiQBUP53LE4ClLusFkiwERjvuAURj2fm
8pRKYFLp7JjMI1XJyJojFERi/+IASQ5ZHWBxcsWI/4HWOijJ3sCPK1558QGPi3/+
i1OtBQFRH/8SYdPA9Ot/SMCrfOIQDrN7SAV4VYtMmwq4FXIw5Mxi5MfBTziV2hT7
4YJHNgmNUa511oFtsCzw5krJCAKHY7fPG0aKYVMXgEmAukfjXAvu/1pcpMEj+Wlm
KqjAYD470BtqYcNnZjZBClidAgElpIo1JAeMm7vnvRMr7f7fuNv+TO5BXYkGaD3T
DbjJ4kRpAWHNALQN/Twdi9i0od2+dWAaSSvzpdpyPa7Fm3ydul7SFEZ7jaaedMkt
VQbdahF4buWOgNkHlf/ax98ZzKN9KW/FmlBQ6jAqDpxR/mSI1yYv7SSFd9tjgTuy
lepllmpkggeoMotTETQobN/P+fkmlunwwKykRxn9Lyu3w9zHQxmSh2hmJs7THBSZ
L/GBnxinzI4BVa1BxDYOaDcmMAFcZFbDqmF7oMLkw9ToHviVJ9nEtpbEXYf7A97T
jjuub8k+pL2L18oaOtbbTcpyqMkGz4ri2rvQweI75HB2GcLux6QuTLX6bOwkCJK4
E9PbBaU3tqvnUTlPdo0+G+t/8hML7wGETPFiKJdPobJ2vca3UH7IjVmATBtlEoib
QMyHc0EmzFua8nips2P89Rh/XA0N+0trvf8+u3UNwE6IT/IeuvfvIyCUDvKTYP9a
XtTAarJ+/JUbpWBCSgu4wJkAmcUq6w0V0oc6tKqI7NOuG4gj9Ve9rCNtHIYq8Loi
kQd3H/SZJayglgZWsouONC+tbmDwbpVE2RwiK8iTXpQ/V4PE2+BPVyJpAfWT0CKw
ibkUZz4CBcOQ18tbgkhZZsHncEQ8vMhJRCu73W1cTZehfcUTUjcoZ+FPwB/MdUbo
YBcd/q+FUjnb3eVo/7ezpSsJf7nmAfDm/l7i3bnqdvX5cQ2ukaEHMlA0M4SuMGSi
vMjgcpdUulza/wDdonMUuxcvb4CQxdtpsvi1o/KQZYTeXfE0D/gDbXiov1jwuvWz
xcFch/oWfpQ+i7JhjLWaqghshlVsiIgmnquI1oetgEtiCdY6ddEUir9fHHTsrL4L
Uvd63VBf/i9g0xsn0D+3a0hXx4vEF8aMU8udw9856iTsLWS2HJ5WeMND1vQ2fxvx
v/io7uDHYnSm4yjno03emjYsDTbWRKxoLU2WHwrj5nUy7vQu6Si530esBL91mOts
svtCeLIjogfDALiynp6mE9B8V5eSyfjPJDvu7qhKtBAsfbDxNk/GxSoyfPadzGDA
vavtFFws+HQtRnSZkZpG1HCRM7mO79DosLGttiGyr41IFPHQNom4cLVRRy78Dsxr
i8v9EEcqcIlBUF39wFaRPXyKYAtUfkkYIPqY5Pd0gNg7sj0K+NQqpEim/R6Mr7Zt
ZJ9p6rLiLLZ7nz8y4uGIrKNOfIj9FoaQzcRrvkVB+NrntUskoOnuVfrTV05AN6+q
weSx7Dk459CL5o+vDARguWlpPTSA6cuoiH2S7UAJzz9NYXHyd6FGGjH4CKKcs/SP
fNff/E5cm5sDarJvP1/flKy9B/T7kEjMW9v66BWklOBwRXwJNpe3rNAZJCGHjR3/
MagMWPLofESEIEqDKUoI8GgPeytxtzwpUuAesvG9mQylT46qJV3mSH3ClMm8ZzMg
OWwySgvfa7bQ6+SdhBdWo4/y4MQi2plNs/m1a/JzphzazNVB89IpMbQ0tyAYdzxC
8tHRtTDTAWCOVIvly1dS5W81pIxQPTbMrPnLDs8MCS/47r/eyx4hLwUNnqqDaYVU
ilD0qsGmAOmE2sotUouPy2oD0Rd59fY/oJhCvB51wtcFfuXelDrKxkl/ZydKXSBL
/w9x3PDL1dQ+2MwzDbOb2EUmRUSeH4g/e27hUDTsvHDxx0XzFtSEWsQcvOrnaiOT
1zDHwmWPPLhetJ5buSFbPT2ePoCiqCSby023H8vd7meAoI8ehTsTgHGXqi53Xbd5
NUpSUwM/rtWKHQtarmJ7uvxrBPTF7mycdjAWquDkaAnXZHOjQ3Ycow+/WQUILBCS
yoH/GO4xCWc2w4hg+IaSZhq8KL60FMFUwaGF/qd38HQSX6km2diWCZGdLRyRCADS
L7zGdj4Mcl/FhcCgoLUHJDh/GUewCb+6KicWmseCHG+uffPETGI9fVybR5AyQG7O
ga13Vj21Dram9dP8JVprZ7++1Y8tVd/pFyOzw8i0jztvT0HlMgXlPT1dztLAwGA3
1OkmsLaZL+aQjkSu7ZRw/LEnYGrWl+DtD04d2yVBrrl1Ejr8H9/jqiu38r5RJ96B
MoWPmJo5UaRKVLzLimHA3T7sppp4OwMuPXsVZOIjxD3uc6C5TJ7GVxLjKHc0YuLG
5voUpcUMWmhpdY6UwRHz8YMQBFLhOpXcCtCyrLMPA8N6vwslI1XP+dwBuk9llCbo
EFpH2VhqFwj74n+MsOFaX4XCNwd/qhV6//kieCwMsehrG+oQJJd6IhwypAcA/y73
CEfV7pyp2DMHR8JaWgjkjDbObiskLpOTvs0bgt+hsY+/LWHa5G+Lb1QxpGMlnSSf
0LZj7qMwi8jqO7tK34IAGeMPqEKczuVhzq1tYc+gm9ct3IHhzTYypDwCgnS+aGgi
SmQ9ClvsQGXVDWZK7nFyM//z1r4zH+nkejUThMXrRkgaDqDMd4QLx/d+hmoa4E4n
3SBo7x2vPhYqO+4privbgfN9oavljmbspXNXPXemkJf6T+wGl9v9F/jZUcrPvscb
KlxW2s1WoHRjKcemv2mYuaYgjb457m6SsInzgikBT/s6QDuUfRr9N7Q1k3umV0xQ
VpHShM4TRe+Qp1BOZWxa7YoqASe1j3G09jhEVrQn7hbsF9WUlEChn3tupAdNwg4L
zSMc3pgbnx2yRxhnfromDN6or/Qa8hA9A1oYvGPfUHuEAcDGrJky1nKK3EIllA9R
AcPTfi6KqDZa3A4KYBSlBrBXMzTq6oneSKr8wDEF9BgKe8BKkL/rkWDNTyP/T2++
OF9kxNyM76lgq8ASSRxC0KKpBhpSeYJo/0W27Uhc83CfpbJBDI6UqTnbZ2zJtQXR
h9comULKS3hIfY7aE2Pgsim8bePo6PkiPj8Usg/S4gOmA1N1pW042swEtQYXxcDy
fspvoOPylZj8peWw6qIUL7aZPsVeAos7wNB8tL/zdhNoNhXhkmsZK6lrdNTa+51d
c/T3nnQIAW71u8wCNoD0Sdte6lDRP47o00NNfuvug3WXcWKJxUWdFD5XddiZQm24
LmBzkt9FKaqXINuecd1J6Yh+gjNICJ35XnwTAQJv7KzWS67gb4ez9mKNL7da2x8x
atZx7i1Ym6DL0GHyFZTFCggnwD7GpofJi54zF03Cz4WalaeLayWqk4I6qI0xAVn3
m/0JpvzXE5kwrVmaZj+h/DJRkdxJw2XtcqDIPwdwtQ/pEtL2UsG8Ra+cRwrsJ+wS
qJEmUBKaO3kt2i0UhZZSz9tQKnpp+Jaz6yQhWumXwLAOo6edSeGMNAFsY82Aqrwn
7POyCT1dldvWrhrV7ub3TKRA/4w12p7Eg5aCFvUwukJBgT7L0hemLkHsCgpgO2Ek
fMIWTgA8Dlq7ou2Mgisjo7GzzRmATX4gYErl3Fd/2b56O7UlVNEyvT5U3Jkguar9
oqZhAd2ID6jeqW0jrDCJmNo2j30XrbB13SvwWlQONofZQm466EpNoieM53WHP5RZ
vG4dodG2rAgHaMNdhzS2szXc3L7VouZdO7nlqIcXbRj6MFdHhsCHJLAQHmxwDQ5Y
6+Wh0fAJJt/+SknLBiFdKLn1nwDr1+YC7+/disJM4LIhPMJhWIYAMXO3hofghhwy
dKo95fD40qhdYICMQkG4w1IEoVRsE3z83JmAAmueAt41rp0of6hC5xEL7mMp08r2
4l7RiFsVgG5fqtuOVljeCJQOqneyCZ/4U90MgttB25WjLUpWvY2fneZBihnN5aRr
35Hygffqn618+a5MqOjyGcfDTJPRa9EJonjHYUGoq6wpGyaI9cVnayhhiMP9DTtm
vtsyA1pQ0m2eQIcnz/LzRfH7iED0/Q2TqfIG90/5zq+6OysrLdFFve3/kesYVWxM
ECYuRPrY3l5rcc3G7oHW3HQ6SGMoRs9isrNMaA9rdXa9SEzsgNVyEI/HYOlpNvZG
JGdH2+non7ph23rqvbZwAv+Wv9i4DLG1XjiGydaL+yZezy71gHTm80H4iLMmKtGk
j15x1vWtQFttlHz99p3ipCkUeMIxAfLRrlINH0TMoBy1sVqM5u+1+eYO01hCEih1
KEa+YUbx9a+O9rPy+ff35MQuYdqLcU6F4v56JsjRORi0j+14GwBQeT332wqYbF8m
DEE5K7qqvmbjvOoW9uzJ3bs23MGjTum0Xk10BMmxpDG8Nz36TXo6dnJqUqpYRJT7
8AirKa/cg4qI1Fu2OGpgwhSzNqbTgQt3EaBdTv6YLTOiO6jI+DnjZRyBQGK2vnAs
Vy76ebjSnV7eMZAkzokgZP2tpXj2NAeZl47uEIMnTpnzvfNL5H/AjWbt+N9TsVp1
LlqaTeCGG2zZQhyYBiZivjgU6RLkVpCIqaN2M06hKekIJoENhfDuxxRcbB4419c6
tptHmIYH14jjbMc3jF1gRBtnjAAclJ0HV12wjUmmoqPCnKN+t++o2XdjgGMtdnMy
cO9MydSuHUGQeUDhEqbW/VXisIIG3rHhu0Aaat5napqaF9Qr7Gj6IcM66fhEr9lG
2HGbNVetFzO/o5X/6MVoii+NtTUvF0Qp3pF3Xmuh1/ibQjbbpUca2H9SAnbjdwG2
AC4w0HpgktFVYeF2iQu3qVwKNyTEKLZqBoh2eskHfeQ65AvOfmiBCztSf3x3Xil2
HVoT3HozI1AA+A+MjiU/dYV8a8Pe4ekvja1kdH+BlYNX82fhnL5/dJePd01mjvkn
MBN8O0cJxOhxlp5ISy7+ea/je6h5h67Ay85UH6EV3QsZvXzvSIaD5aJgKPcXHpv3
Giuo/Z6Ss0L/epAlNzfmvi9Yx67OFML3O3UgM6AXEd43rRGKZ3AiQ8FoFx1QmhLB
Pg7w3gggD+UoEjleELck8P6SzPQ/u6OdalkOhbvWr2TK/1UFXzoh0Xuwd8IHV+JC
v3oomGoxT9LTrRT33U6fjbKpseuBhYg3IciZmCFC0BbNUb2a3OxJ81KHNQBccnZP
nY8IDbPCrG/CNcJixd/cQYInMsDBdCU4cucYGm2uM6Qqkk1dTl6LQ+ZCE012nz52
JN6aAE13JEWMpYs36fVvegXxZ0P/NJ8/bKIxAMvN7s/pMad/lNLUI80PctAeZVld
TFqptDDV6WsYJ2Cn9qiSMQSYVPlzjMsux3OwlplvHdgklyK0wwQmsCno9iSLYUf6
IB0qkH5QUv0fldogPmqq2Tc9ny9znC6k5eCq35eN7h2GI0wm3ktX2DRYWntudG/R
xvlPkj9C60gL0FZ1bsSQQwxnaURn9Mr4nfOJvk+3ADx0hI4neT22KuLC9BxwB3Vb
lyaxIcvwqHhTabeJJAKRP5c9KHXuooXGNBwxGLVt0QnenZUUzawRCQ1z/nvxGq55
qWFV+2L78tkyJ7cuo0wgy2tUTajbzfZrMyuxAtmztf4Vb+/8hArHb+4qMODliTQF
vkU82Hec0SRg9rjJ8vJHp3hkK/kWCg0v/ORU1+2EM87UNFZGxx9nyCJEm0yk5LP/
3A8mA1fdMVqB1fORQZudROOOBrhnKgwe8kp+joPALhZ7VoSSzRHt0ZXXRg+LLksS
LtxVQAVioVf8QOKdHcp0hi8+wThiuBq5J6kRRlD2U/veVNVbFVX7tDKvdUFfK27X
GQX6EiRy7YlEnSBBcDaNGKqZT8zo/x24aqnyhErsOe53Uc9f+Zp9XLGOplTTJ81A
tCUmJpm9D0bLA/ZlYFCDF3m82kBfgTpoUmLRjYhzIK2ncTH26ExsRtM8k7vlCZi2
AyeudQuPdesTZsJlJlEAMP2at5e7vT7bitveyJP2vkFV35QUKuf1juEusb5wt5z7
F9geEg1UW0KKBUKqiB3CWwKckl31aXdufVyce1secQsIp/oPlsyAqooELfAR9TES
JT0mjlY+tKQjrtCyu8PeW5QE05S0yRxWHVW62D0NxLbqjLH8GkidbZuAYZ2LkscB
k5+yCku7NPXW4dLcAlWfwJTLXbsalDtf+bXI4wtNxtpfwGi5GNi3Uw0J0oZTNRf5
c6d9pdXjgXHPjXrb2W3vGe5sSeKvJA1U2aolO9t6sYOJINNFOE/jwIDPVB6BxJaL
WQly0MwgiLzx2+W2ENw7tgIyZTx+6EPV4L0NUl3Jay4G/5cva517/BX19pn0G55a
Wq/Te1Vk7zXKHl1eRr6wheya+AZGQNu1eogSs5f4DyR07iAcnJEjGXT1QTFMTcrL
iq44ScROSoniaqMu5+qbwAxqDni98RZx6GB6Z70yM9ZCB1YK+GY3mZW6gBCvZ7Jc
ZJGM7Cusv3YZ3W1XnMqzE+s+ePdoEUmnp4aLkFJmPu23cXQrf7P9LcR2kp5YiR1X
2IXKLjLlAVppYzAOeoatUAV6x3MhHAUun3Kp0XToS+ytl33K02ox3/bDugSGtAeu
IhpqyvOsk0uaBfTbM30U/ImaqTlc3+JIhXrPxQEQQLFPMiTi9SJ8JOqzv9ugLxWF
R5w0LjtEs8Q/rAWI8AdWJSbB5a73AZ71vj+3PPCtGD9udSsutrupIhRcuke2V2uI
woBfEboaoftVqxBJX5C1aLxanN67hyP0oBNLVqOAAmLESCarR4qDEjYhdUPY4aCG
NQCnn83me15YINKXEFPWJHSKnARcm61BTFT2KoxgYdY21w4914OjzR0Q09XBlvSG
frcItuhjCj6dlHl6CAybDtA8TXqf/u0Vs325CRAaaMVCVBocDE2EUJAy092ljU3d
kKRpvM69tfhGwLZXUps+hFugg1TwBt9ork4YcCaxtDWMZwkzK4/UQJSUBBFsLsee
AZIqVxl0eJnxG39yCkmLyVpkIk89I/hEMiwQng+USiDm2vaQpSV+hVutz0oZXoqT
/aD0xOpJwyjmNv6S13Jo7Eb8IVvHBmlGId3a4WxqSuRXDn4zE4UOE8VGTmAjpxXJ
nyZVcK5oSrfhSJZ8CVKEhGLgoHGSvx8AYINQZ7ZknomZ3N4yI+vHSOoG4QOtZt2+
ZUboU+RAJ3oLux2JdkboO8Yqb+DBQH0QFebYg3Og/+l2Xc8U86b3RMHdkj/QvkWm
YERnMa1ZjTLbvrjy1baPstPk4HgzbdAuq6SGFsed5eD8BWSNV9vpKCr/IfJMxjzr
NARUYWhV8xGXn1EJi74TTYr+R96Qd82P8bk1ns/RdsFO9RNvlZ4fb/+hyC7/7dQp
IRME5yG6gXZZEVJTgtg8SL+PwVEBZVH4yHsEopVlEsjvmKHAxVqrW/J6hXKQyYSb
tWxXY8JJIzGCya5zvBbph/2jLQJYCUi9QkTZs4MCC0ePLuyRBiJoPHr70/DpScbM
3bMK83S/0plj7gPZN8wqSkybc0Na1IJH8JCYy7ZNFykKJArE3aCcVGq+QmSsXGXt
VPheFL1YrXlpqQ5p0Kvrxi3r5kt5XaqIRRgyq0MGH6bI/FyapKQ1ovsZ1WdnB7Kt
IJ9Eok0OJ8BjciAWU/nuPzj/4A3WncVNgWtwRh4a5gW8WW1BYw8sJwJ3/JAE1fnP
504vCOHRc1jn48o4Yl2k4ll+fz95EYupraXAZEbvS0gFm7EnT/LruCEnDGW1tbvV
2/hyo3b/nB4KtT+GW1gquH63IcAph/xTdUcqTLpBTbN1ZnAbbpBSdYAeOSAw7V53
rtkuQgqGl3lZWDza8slGWZ10hMpJMAwen6AnB1LOy3pDmoyC9mNQk/umJ+hU2vJT
mrynU3BpEpGhKx5Rca93/IEDSumiQzO/DFk6vJMmOagGtEv6i6fRtZa5ejvuaUoM
OIPeMwzn7elWYwsgDEDTz9/TAx2hYan48X5CZkjLIHRsjlVuEPZgRVxq9xQiWNRd
9/oRnAjAsYsIBOI6/l4JRjt9ul8co2TZiAzzZhouexB/72shP7Y0/hFs8kEO2BQC
CudsL5UF9RqOLDJr+qOqCNRd4jthjuTaoNxosSH+tN7hyKbjmoWyLtGEj1GVQamW
kVtc1Ph6QgbVyRxDjYlOuoR65/CIYH1hlns4GsKzs/6A7SpcpuiGl+g01cQoIsZk
00V+rZ7M0aSSWb5R07dBM2vasPg6kByskkEfR2z27Zj7SYCML31Bwh5xYrJQb2t4
0lkS19mKfI6Lzu6ZE/Aokg3vyrx1JIPlzls4lNRIYagEkZXcEc6erAvvuNuVV84m
DkOyucLdxuocR5hsAl7jarDQtXmvYeHy3/R4rxyEQpVWTikBrT1CnYEkvqVZswWW
oJQ9FvGLd+QI3m8wd69VQ7OBi/km6BSdt9K5gRF1XYjclcdoshNVvSI7IUgmliWJ
2oIRZ3EYY0p9Tt3kPI/rISkTFHE8LA5wMWb+zktBe+gNUNEYXz+dYI7BEqwEPL6M
0jIpZCgrZ3YKvICDPsgui+F9igYBe0dH0VN15RtCJ4LlPNPjTTPNw4ayLRtsKYB4
YznMlPSyszCx+Vq8tIg/TcW2StKcmh22JSgaLsLFtz45tS9mkFYoMdPcPu4tRYvp
XkHvybGlYVzEV5WcmPX9E7q62Aozoh6vpb37z58XkHJzHvnVR7OoDoWc0OZp1QYM
pz27NAo2XzIDzvar6u92IUK95Gzb3qw69n56f1slEwQDeu78zKBEGYauC25NGsTn
PniGmgNh+jZhsGFehG1MmTnSzwYQMHuldlgNWbhmexM0aA403IyZfhqXxauaB0pP
+33D5W+4qiYiW5uqviJK2ieUAqtCUZMboz9bv5u36f28F2HjSMIrAV5ccBjWV5i3
P9fpLtih7SEvEFz3hYx3brU4ZPLDpUXTyIVCrG5zhMIZ/nMcfcsjji+1e/fKLWyZ
G0qqLxhaNROyyMUX5xmlWyWuIx2NnPk7RZ7tEoM3u1auP/Ia+4veVvYtRZnE8T14
e5I7SSXoITTVyxSxlsc74HQHqmiLKhUbQB3FdEVyreJ45w3+fmepbEt2Fhk96UwL
kD7/hZw26j9lz2R+KrDpcmF7H/eDQmvzz5Z/0QQhjbcqenzPeXsTnsOFnAV/f9FI
1xaC4yyNcls2dWRnM+RR238F1troye3FtpztuUyBHlq+Uwi1VGAAIC0IjC5c0hB4
Ozj3ozoljTFmDPT9yXbiBt30ApPNky6FipKkUXN1Nqv8Xccgy9JNRuD4xpHp/jW0
bguWJfDsFbPpzSbbJt0NMeGz/EuQATlJkYOgrddnapGzVA6kRtJpuPXi3nxqPl6c
wyb9sWhTv7OSgWQ5Vy1UA6bmGVFcLJwSxr4+T6RyPDTFCI8tYEviCQVhL5CYRp9K
veYGvH8fgwltCbXGw1ybS+Svn+ikhFLx+wa1HAwYCYhY1neRYXkj1RbF1vTaEYiL
pvfNB/cDbjAvPGi/zpHgNwqM2Nf6J7MQx5Plz2Gy6NG+1kMMWDvi7ZlebksTaGJU
+jz/XTgaJ0uvkbz6OQGMEGpGpH/PbW4udYGu6oDG8bKvWcEw5QBbXBZ3siSVeMB3
W238UDMWvrtVMvqrQxZyN8bywROv8CqJqqb2uKI8ZoTq+Gws23H0sMLGsQa9ew2h
xCtzDZXl9zhJ9PxKbGl8nF7jcZJgWLewR83mntYYwfIzfh0vGwYSQvFvCuw+ZDfU
5hfcpyKNvVTk5mIBIcs193yo5tGRBh4yzXlMlt0FNzMeM01HML6DPhl9Qmtft7yg
J/Wv2IamKT23uACokbNmhPzzIVUf4ik0Eg1Je8RuYqx1fJWdCOrmIRuq93oyvfpD
ws9J4Ocoo6M30ENo2Uu5qdk+9+kjZSXOIC4kZfZuaFLN5P32QSP04VP7yi9hH8DW
bQmbEYaDxLFur1H+CcGniOhPyu9EDIJ1xh9JyhXR4LNuYhU00V3xASh4qPVGS++t
jbDxk61jN8UlohoIFHkP5X1sLaNckqQJb27cFGUgca9uj7bPnxivIpP8OefWPbbs
gvnVBaz1z4+/XthNd8xXs0zzqTEfs2a34g3zv/xvh8IEyas1Fs2/yJf5qwQoYmLw
yw1kblbLMEiEmKEpDSg6M0La5Mkqo+yRcq2SgRr//cnUfKajyaLnp7Un1paUOkOB
8IlgbhOBS9i7GNxWdjpM6MglVopt2XBWmrRtjAhWTo9h9fN+8u4f51z/zr3cb6qs
1zY8QmbCy1mTlIWFT+P7jjUyIyxIro3DiKQcciuL1Jvbl8dfDvtgD6huUnwHR4dx
KvqJQx3Ucn+QfJvkBuEY0oIdbEQutIQR4OONv6gqoVZm3KkM/y4oKho7SpVJrcnF
dhZhMMvy1GT3mW4iJvuYR3vPgPiUBDgnqkTz+5Y9Rfq/YcP/DjYB1BZrjB7jQHj3
mnj9ZvpqjDBhfbYc5fh9bJ7Jn835EZoNMjXj2hqzzhrh5PSvDvn5JrmrA5RuoV3u
Ohpvd1zef0zXRdtbBKqaUQvj3V2Q16iIpvTIGFvKPfOdAV69B899wm0J/gA+zoUH
E6oFS8N+qDnvesUmOfP1FoD/9VlHLSOPVsTzYey4yQjn7w1McnxU0Qy4Z4ry3R7d
rEaLbs+dRHJ0PGBgn7pBKr1Zre9Rswa/SMiTI4sLAllMCsvhaL5aar59q9KDdH/8
TKFpf8aaTRFnJB3uudmRaBhUwmjsju6d1E/bt0p+qIlTCsf6Il6rapBuAmQ6zzZ0
iOd4hKTh99Totm4OHq+/PIH77dfGj1AZs1Bo6qzwK6pheGWXQWJ6fpwEdOfC2FwR
/OY3KGGJsNVtu2BgYREOhsFS1CYm4rTctZIC8YJnk1cQAtMfBNhfhT0usY1976By
xnHEJQBUjZxhSgYdc/E/6IK+u1+Rg+4AVHzndDq4LGrwEBQ7ugC2vhaed9CF32EF
2G/FwX70fXO54WgKgpPsDLGdbrCc1Qnv/FGlUW+aBdYgQRXts8diKqvaKN0vmJQv
cnpkrsQKeVgdHJi62AKahA2KduQEHuaah/4C70KGX17Zojli+Y1WcgTZwTN/k3o4
jAZQCbMHlqgrQhc7eFIEOYzJ2fadeLdBf4VZ7d3B0pzB1tcb+wWWLlJHYrs8ksPf
hwKpvHSyFDBgYNqfdW4fmuJJnq2alt+kme0xyU+0+RjpNKNMT5zxXYmVam5J14rL
8DG8qo0fp1SkbdFa4hbkwb7J6CuRakD7Jmg0wmKOf6oAFa6Dm0801eWkG2km4UK8
Yyz+QdFcVkyiuuLoLWgHz+iebp0OCqqZrQvF07jD799e5TkAEG2nGX12p32hdkBk
kkg1W9q3RpX/b2DtlRRvsnO8ka9/0q8JM2vv4+SHM+xLwzreXM0+HtYkmuR2kZhG
HHiOzJ5qzC7CfERs1yTXw2a5UeFeKjvRw0ykiA1U6FuGJaCd9oDmEksVXx7e+fka
WxuxXkS5ou6mabLBMyvS1NXd2KjPdhrAwGpf9Kxy2QUkPNLwtJBijdIVu9XXQpIB
+SFaWH+Et+36o2vl/C4FK+EIvLBY/YLpv6Gr1bf2WpSfsfsu78wv9hPx/RCrzuEz
Zt2eFhvbrUF9KAAkOW5rhSzMxiMhl0qnRbEOqnXCeHCg2xG7WlrAuIssL6GTEGwG
Om1sNjCPQVGs2rtLhedC2pMRzrG4o1fMjKmTstIeGj9nUhFs9yA1uEWHo/KFWlGv
k/MwPTvyZCVVY7S0P6NgTmJ0AN2w4bIz5rQhAzt36pCHq2y3YsJdbHXuhdtTiX/E
lV24Yoz8pif1jXRfdU+Uyqiepx966lXncZINpKw2TKq7qMZzxR3p6drBlHI+5A5Z
xmDIW8UpUIlAcpDiXtJXFm6aM6qhNNdB4WpTjD6+gHta7CiUAfyA+aTUWFDqUoEB
WPC8cxrG8iyV+1uBDl45wsTK61FXmA5fChBjtsCtIy6A+Pw1v53r0ixN8tloCQGH
bhGrJC4E6Vbx688T/ctMJ6rhKAxDucsSvL3Z4ZVIuHYuD9qONO51eMXpU0RzpBvb
Pf3kxy6k4MGiNfBbdJYk1MmmSvyk2pAv+NCCOwlG+CSbbSavgAcjq07PvNdkZFMA
9UpzsrSmUSfBAQGlB7I6Zv9iN2SBPaf0PxdrYV/6HOFTrPHCwcNBZpUkcZoFRHA2
UBw+Hyh0aOO9Vv6kezfSgMwJPPVcfTML4xvtU0g9pblmtcIOl4HWjg5KeDwY0Qd0
kmK23kBLgWpWumQ+9fj1sQ7t2Gl+CE+pp0zr9OnUI6zCTZRl3VFhFjIjBu9JEz2r
JtfA+h9QmqGIzaM6UeRX3bwW3pBXaHB2JY57sAh39K5ReIgs70R4rnNPIE7pk7RT
+Hd058yYpkLbRpNlEiBYF02/LNGA/uqTL8FmHJHylQqj6Thm0cyL2kJo+As9twHt
P7EkICwEx8CseiMusgc+fxUEloPH+6bB5k5wv2hHcFdBekHORXQ4Nqs4Vb2SxVV7
GkZ/03yaQpDUEX1zxNVpSdPFvXMYdSkkm1kp1paChue13PIieR3olbVnHHpbQXuh
AJz8F6ivfoiszCli/e/srS1bcS5qST9YJPUiAjrxSDNZidZfY/PWNg5sSK2hOVCe
qgPQmb3mq5YsFx+w0e15h+RlTMtycoCvC/WaJY+Y0NyN5cHbexbCgf90YBJd3Mme
0V8JYhrEjhif5x/1qF9bkRQzH5JdTPoQ4o3qkWhiOzuAk2X0sLQiRlO9aB43Brz6
IkvC+du32AzHmCB4R1EPeWxnWZQsYtj33nGwwblGmfXhrH3Hn5YnU4jQk7wmHLQt
nIQsAZ8FZkg/Xh/98F49hEVT0b+3QuM8QE8uEYg0iTwO6aVL5ayHxYR4YrUEYxxx
yyuKhZUb7Anmt6e7LmZYyWoB/CxQTDIwtJ4LjsA7qfn7EE1ElaGI5ihKQdiprFK1
f1D0ze9sz/VQnE84GAM1l50l2wyt4/g+48Mbcs9yJUHYt6d5BuIZIcK+p/ysOnUY
dkckb/CaTzCRzHlG4M9hIgzzI6O83hBBcrZBkUvI8xADKbLEFb6rG93fyA0ITSHW
VzYo078dpSkUjh5dMlNly/VcJ7Eigv+W9fQmD11eXHphZV/3fPrFeYTGWYXM6F1z
fNgjZ93CcEv9gXCijS+llmTA0uR82w4hveso8pQVh5aEqzyNbLGZMUyppo6BJctP
p8FGaIs1xjYyXDI2kf+XkpJhNB8kZW5Mv+/QIii61SVbpP4fYAaB1fcTTiQkP45d
Ht8HyVPyN5e105ygJdzwNFjpmG4WObdFpPP48ZiHY7pHMfY7nEP0lupk/7g9F8/D
1scMY+FjawNgNwH4hWtRu+TWNn/tixNB67xy8CeJLgco6Skt2vzWkm8D9/IbOPAR
nEwEV1/S2aI3tQxjpnB9BTNa9nRArxAOZBTVlekM1gtFd7uqSodFRoxWF9Kcloi8
tmwnlItxVXspS1tI/PHOPcSzPRFLqhS29syyJfax/Gi42UdQy77GanByrBf9Yy91
g9CZ7eUm4LDANqiSXxXwlLen0JOIRp1prr9HEUehfqWET5fbl843tZ0y6h2+3Ah+
vjVciSejffjahKmzCS2KevU3bPpNKgs06cDNoWITZ8AdrBfwvcVTxzukenVV6lXq
NDWH0kTjbgT7LDCNsYDT1mizfPXNoS8OCaB3qwVMXG6rJIaqejmZIezE53khimoV
udpQxxf5E+mF96iZRBfAeAsSleETYjN6/DgFqv6UPbPU9uMNC7RZztGmm8a1saH5
p7In1QbfqOw03IxJNrZWeL5YDYs+KjLP3o/EBNom2CV0eMfHgKskLMaZk8DvExw9
Oi5rCFPBInfbIsPfWwFIj6ad22NQS+odlIv3+M7LXBzAtD01o8tJOfimmPr/ekKn
rXyqzG2QPRE4PKMlJAjT73H1MSk4PpennRxYRmsHHvqU52pw45RsH/6rQOSGJCXW
Y+FcB0zARf6yDFART1iH6YMhF06r2OYv6ZNNKEC46zeIECasEPAALaUY/rU7zke0
wZqfE29ueiISHXfSFaaTXgGP7bbF5Wfn6DsiXXn+XpuE0LZQw6lRKoBGvSbKvmQk
SdpMdu6jxyQQ54dPsQARZQQ/L8/7RaSIyca/tJ1R5DxyAFI3uFD9JvkI/OyGtN12
DnWy9r91KpO0QH79Yl1bHYXPNistrh4+Tpr5ysSQCItmr+lpwcFLicoOr5skUuRA
e/eu1Z1459Z06bnZ1wU19ayGZuoVFsxFW2EZ9Kd4IUrOhMNbtxs0fgwPtcBzMEnC
pyW/vQ1MEVAkhU7gW54tnImp44Wz1rlb84wW5OeDCyPsAQcG/Rd82sJpnns7HfM3
JjJm9Dar/u87+WYhZf+0GEW3FzFleUUhyi+/V/hyb3g90aL+8Pkc4LNHjr5WlzcR
oHxwERC33apSr0AqFv7ufGIqmVVp+bDkosH3FDvQ0OqcySCsOoU5495XBNAvJgYD
jGF4xOCbyzZzDB8DozFhngVIZQpL6EggSFg27oD+dO+aZ6cj6vVHDMvtcKEF+xZ8
RnV0ujA0El0DqFyN3upeTR/ShaaRrTllN064+YHlan9yo95ORWnIR2VID2k4eO39
A2FMEYoUjVlxF6/WbTi0bACvP+5kJ0iOxGY1IDMbNmISQW0A3dtqHgLhMRof3ZbJ
AQlR6cvzEK1p581K+ZoXY1YF/oTHATidmtV0KPjXk8S/9GOh2Vcg68CkId1+8CoU
2tNkct6qrIgwMMANQMoptmTWM+zNfX2jtF2goF4GViKiOCI5/fJG0LyuSIV/bVYO
bPzZUbWqFji+IM8Ah/X+s/uQGhyexwu8xDm/CbNhWx9JDQcY8OxcU5a5lwyTKp/L
fov6Ls+L9xytfBNPetPbLaeljMfrXqpWV6kGssofCAVYy2Tfv4N5IdVINduFBrjr
w9CHXLY9PIEHU+/3anQcVvZrKt6etA72+TUVSEgyhSw9W67yVjebbO+pge4NFHG6
vzaH/EeClS3xDu0cJ+1INXnAz0wH9K5Or94+dBt8VcidO84xpBpV9y+8YbGXC9k5
/9gGVDZtiF2lEfC/p4Ay7wk1rAl6QxbOIEto2XwNp2UiLXisA0HGEESGxtbILNUO
DGC8oUHEMptl14qS4Iri3Tk8q/hrdln6FQqvVv/3rROosHiz2Zy5sRgrlOupKpLy
Y5urinhMRO0FeS+ySbIMiYWms1BQZQ03pH1kB7bXJN0XtooA4Z9ppfHmzZZDm4uh
MhLmEUkltIdH3qoF51IFyHtCmXHFEXDTLPW4MT9+B3mzZl3zWxT45+Opx/pVGZeR
9z5foCNG1kAjKQs1pCGHIPmM5uSxnrdM5O3hqw6IfS8MSZjaH08NncwCqpSegcKa
9LE6ytBc6p9eDuAUQHhiAX9DcRos1uxQPhWK1eaW7dY219In7RBrdd1Oi5DgEFXH
52cHoLKvdBqeHSuvzJ3U8SAQMeoC2Xh1xn2J9M+Jv5l+xRs1CRFB6SXMnlWMMOdz
f9eqZlXiZeBF7Om/3+2OvlrW3N1whzFZK2KCaj8Ousr8TcRP+uZqBbPU7MoqtztQ
t9ElciazXCU/dwmtN47ujYpWPD8v2scLfn2a9NRRMkYgWjuoXePhfG8S2PPR4HaB
HD0g1/tznxrp5g5l0wYnoEmf83GJuI4whd2LgTdVaQvknCgr2dSrn01sOQTrSgFq
8M2xPp9M+wwXmD9vEyj8Gm458FPKwVHivTOoswGt3hsJzDvVCiedFmohTBcttJ0f
gAbbNRNfD4vIZKlybJqztekxZxaT7pdriMNb8zXl8u/kdh14iHzjS108pDKQmFcn
8ZJC73PJUfwDKLMIm1PVcP9GvsOQYnjHeDCJNdtVf4fZNdhVvoP0Q0j6k4QyHG3C
Mz7Ree9evXeuZM31v2NGgJh9DP1zaYQym7ttS310cHfQkqrAxHO6qJgN4HOFhiUH
enlDaTKmYS0GuWvYaF0MQ5I5iJYX1SMET0A3GabxfR6G1qVDO9sAzJIKnZcdt/f1
BmCG2vYFVJ3ljbzAF9RVRyP0aO8Ug8Wq2oyVjxChOyrzs5piXkfbDAqWrnKmeQtX
xcZ54WDWFRtCdD0rOtsnhDmLWB5IqkofTCcPl77rFlSK5MpT7K00EVgUDQG8fzo7
kTXJjjLuj5eF3fXAp7D/oKDrgA/NEzb8jqMJdRHujNQrCaIUryZHvWW7sNlAOJ7S
EBBt8REsU4DvFh0NMRk61kOOlpkyQtBAF3sutacVJqTKD0sm3Ef3l4udn5c3PSzf
DCo5oLNGHsmRzyto1GzOV865q4gc2Em4y4zVvbJna0hO74/XQu0mdsoFIUj2NHg9
x2pW0XY+SK0Jbsc9XKNiteTQs2MJIfxyzZfJdx4vVyX3pj+AYB0DPmzyFxKLRrYG
VaEjtoPE4xJY33CSkvajWco7/HcatBH3/hXNlTz+lEqV1rCwpup2Ee+a8YYdpguZ
Wg1gs/TIHvCOX/tgYkMKAE1sc49dyLeeH7ApXP2F1mc6Wrx4uTGso02dQ78loSrx
fxZAHghV0foDW6SPBzJp7o0Nj6jbG86ECX3gbk96ZDi4l3GfpBaQihsut+oonfRc
dMhdYkop5GcmLNnP1HL/AmiNq7dQEydinUNN5tCBLCHujyTYLX2SgkPshpBGe7Y3
npOYoxCLelxNyWYNXv1oxbf3nIXgstzxG3nY3s2R+ri6jRSWhByQ7LymzbUoY7Jb
H1rnS94AvIZdU4MoozAcqHpQn3Nv16eWQzklaSuntHrZPbXsKdlwbhFsQ2FhRbx8
r36u0f6H+Q+C5PstbSx1gbyqtLZAproJhe90ovLq+CexsBq9bC9pSpTQ6R2+mcKk
I4CPo4+Xb5rTFwvx/VF2DWZTwek5f/nwW5qXQ1sK70iv8ZPzJ837zdEtCZeuDZLs
RwE1EJORtkbYHcVOX9dfOLq+bjvbr9Dk68d8E5qK/yh/WYGEtv3AUrOTuczp2Jk1
MlioxJFGiWTq8gz8gzcR0sphLtoEdyhrI3vgaEnm8bkTY2mnrCbghU6Z/CarJ89j
oZlef0YzpzNAe4aVi4oiQrgVcEh/Xc0SEw/G1gjVXa2OZNL0+qk82CIq/6PIv6CF
m/06AUxny8B6RfjoMc16ynWOn0NnMiGNe8zxiBq92TaXlWRWm3bx3KFBf+024LOP
+BxUnhCc+jAFqvbih+Dy1ZQ8enpN2S79avU6cHXiVLBoY4Mdu6+qLkFDazZj6lOW
OR4lXc5oUxA1TZamX0SZ2mbRXX6RpMyxwnsExkoVJvkY3VvsGM8k2rpM8/yLh4hH
yB3mG5Kd1dpuFkq7QdoZibxDTgh0BVtNXYuvQ2ZNH4oCtAek1Z3a20DNL9heiZGn
0i4airgjBl45ezBzBML/oqc28kx5WeRNuY8a6/PxYmQeBPJfOiIxfJsyV0gy555h
NitLZot2w9faP1s4VYqiVSBb0tmt7UgEuyuXyyaNBH1tCmlrbPTo4mJtaD9hn3T+
YPpiTooD7LhyabKCw3DrzQvddkk3gWs/weqbAC8BihkTNQwGpeS/j6Cw2Xt0O6GS
VZya6EPQek6CQN4SLt18qZt80ub2xWbuZOi842hO2OIkYWXpMbEH83PtVWsuvMa9
iHb1X0DBAXBhIxrsb3Oul27v5jB86wX3NpxQJDD4QnhCdt4bf40142ofDn1vtLJS
8pVYAyznlCIVBKqL9qHpE/v7Dh4EC0XZOla2h0MKeRjLZO2ugM/Ai5zp+RtjQvIw
T0PqVcQ3KCpD6c3gZ4RJTVDoytuleYMtmQban0v6S50lZC0esqwZkQpi/aN8hd46
CTYCmDhzuBKxr4q+ujX2YzTHBxG/cZHdx8QFyuDF9YbpnuaN7vt0St2IuSU5gzHm
SZHLKlHg4ym5OfQLN0upofvtPwoNwI2va1ObX69aMB2XZl/Q/h95O+J1Z97bokWD
aB6yJc76oGcrXmFykHakh9mZM3YgyQPvuklUX6qoYL8KE1LRzvXPghklnbQTci7f
/BpJ7v8SbqWLGWKi29JwwrM8NTF7QF0E7YxDqJoHWpbqOOxKv4pczrEVM9CkFMBy
Xqmbl3Z+JgxrJVmsq0r9duXLYvNqrGcTlS4D/oiBKQAmReqb7PP53bkWCzXD+iYm
EtnUczQCIiK4UHUGK8TZdqYgpV4ih2SC9Etr61Ll+6+dGEkbYouw/4rf3bILWGRJ
Gq6bbQU5/4sraEhbKHueSi96kveFEYzuRbBcbckuix0GxWN0SZFK3Xi2Tn0sQwgk
krPBmWM0arN7C9HWOm/Pm7nR7Rskd613fipCWIQmE25ZhfGEnvXivmbSIWgK5kB/
Onf3s8fM87ymSzzDdhWak4kTrzBrCZshI57s98c75PGAnFEuPTf6F8Ez1GUFrFzk
pNt6PXPXJ3FvhWr3rGe7jJb8QL5nOnxVxU3E16vIcY+RYb83wkUe7bHc7EtvTtwd
kAEZbrjWBflm7x9Gac/B2W+r3Cm8eJ7Su7p0RY8sI4I6MHKED02A67QVsjq54Gq0
V5MErZ1hHLXdj2JUPgcE9HXvKkkynTOzXEJep+yDtUeD+q/nEV8KvUvRIUgF5b5b
aR0QFDdMvQSHhYbX48Qt3Z0HTFgM0ILX7WE1pGiAW1ELpeY/H0o+i+VF6Y746r9l
cuGXL69hcsOduWdTtO0XDe/Z4uNKtjSaJ1nugCgHZUUK5kgBkHKiSPzMNU2/YQHo
6B7YMvvVMse0U1YHLTiLw9PcTzz6STLs8CNuQZsj2do3Qk4zn1koYnGtEKGOlWGY
oyHrjSHkeUFVMtcMiM8PAmqXjnt36tbrqm+zl+p0HogzVdaSV7VLUAVMGnuvtcyg
qfH5zzk15/UnRfpmoWwZJ9Gdh5v4rCD7ZcFKaWUW3ARCXiUS6TmMwdvjIjFGFsBB
f9DyE3lAUO3f+RiUbuJLma2g15O91ELSCBAhbbwhZX4UoSAM3Oev52it5Wt05NQe
x5Q4RDRLOGbko4o+3VI4X9FGXR5TN0WgfaWsyQP17IHpQ7OtK/UiyD9eRfDQE+Ms
pQOvsQMWm28Z1eOMFjKKAw8DUSP4TEjT34i0HXdZ8ZmI4J59vOge3Qk0OocEGPMh
Tlaof0zsg5dOAy9kGfC/y3YAx3EQ9O4WdyCGIGkBZrlUeH35KmA6DCe0ISsjRIny
5Fl37scfeAnVbYftBJNpq5/J6lRqfx+oo0oIoY2nQ4wIfIRtORzFvrLzEofdz7ac
s++p72LBAFP/8NVHxHIdAUNjaZniPYcgIGJFHr8VAWELt3jgYlJS5zR8adg2siTc
G1P3aEgS2jEjSrYA7H4CJ18a/Mu0ope9u3Bz9vBderE5u3JOecL5giNyXQ5RzvTv
Ea1bFNsx3oWSTzvwMeBESEs3zb3FXzBI5M7kTbMiFSzFjKNmt7cUrWaDRln9vEND
HRZOPpfTVh2997UNKksbuYnvgOfM/puTsj72N4evphI1hUb9zqxtX3Gny0YpnHrE
Pl2+uGSdaZsYQ8cUzZMVj1jEEngd4SS8XHWNKa6+SgCDBM7sBz6BVD7Cqhzt+5+7
iGrTDW0id1nnbAGdmhB6YxsAWyKrRFAd1SChoot9D9BTYeX+Cq2NOsIlUko4z3WJ
ggA3oBOdssmNafIHiwXC4r9R4X7Iyy9qk13rIq4c5iQXY2NmrePehMezc0WSRVon
0XhzIrSXgQK1AsebU/vsxNbQXUYfC6j2DBYJuBpH+a5ocTLjWDUPViKyqTa90W1z
KitDfH/bgxJCe+aQt4XHu8iSEjgmH050LZg2gfZyaNcwOU2YMd7tbkFqLfqd0SFm
ZuPBaOEeAZab9m1EfrVeTjQ/qEi00zz9FROHimGm7zMpzzbQPT2Sg9YE7C2mfRJm
c/fuEzk98diW4jgVtOvIixORPUwn/Ch5o8HdGSb8YaOc3okvSvkhsW62FF632vKy
YXlzR6+Zc3488oH443rlr2f0U1dOS1dsxB0EH0YzqnfL1J+v1AAs0FIOueu+3TiB
uuFsoiPw56WcpocxZYydkJLrgCSK2EtXRcrstxNexCGAdHce3RXYYYb04eZ2oiJk
zms6nisNQB/qe3rgk5Uz6md01jLhEeN3Cp6/HSZf3IwbaRIyiYrcaT/MGvlU+eJI
cDjsRzvyS0krgMxM795o6SoilpIkgEAuKvPdNWKGdOEqwzdc7V016KVjkFf9YnsO
MEDWP00400Qb3kPhe7sGNmB+USEy+O4wIrhoFdpQbROuKUCk3eQ0dA9jUIUf9j0s
kdTV/qf6GFEoUlMNywVM/yFY2PA9tRVQ9SPtJCuW3cEJl8A+HbqHPYxlu0ZNIdPx
NtbnHNOfIH9uGSBS9O/MiWpFMsHGRnb6pDX9Hiuepm0hXKk/yLE2vDuZdAKqmmYb
3229SL8qqNWdJ2yW5pO5B9V0gimGToO8rMiawR94W7huxCQTpWw6v5h6XQRGi3ZL
AvYlSEUWdhYXzYLZqhZum4sgN0rZL0Klqx7zlnJpI/gEdJ4t3lRu1eX0dNhVHlY/
1T3GXk18FsAp4lxCdSveqTCXOmnegWiPt1GNdxiJ0OWkEMfMfFeCYk19e938vD4R
YI+5ovQbFGNMscjADqCpcuIXJIM3WVaeC++ew1sAVH0lPp9MznIanjTRgr07u9OU
0Tkw1QNMRgrWfeEsAOVOL8JxRWtKcuperdEQekuT2NPDd+7+ef5rwqYxLHFVIlFx
+iU6tGoVajCnKvDWbIuOPuOeOPKsANQvFsxMV3JDNhtb+WfxIb53nWSQQJCBiZRb
+87eNmhrJwnRzE7b3Cgp4k204Hm8eglw8Vpem8hpJ9UPL7zNOqUZ/XPBrps2UtSC
HWPhvX7Hgw+1Z0hdcoQe2sqq0keRH9My9j/U6WH+vDwXgONnIdDcNxi7IjPN3eVK
E/RA1zN8QSguPyvvJfJHpdrRyJ5P0YZXj4McMciA6oH0clDhFM6nBxq/HQYURxCM
VqLfLy9FnLTv4nzxCiVO97K3E6hf16TTvQ+nPug/r8JIzlqLKetbzWuShcjvtUpf
9DOPBFhpVbdYJFRoUM3zJDQZApTYIkOD/KUULv/h3HDhv59KL66x0bx49n847JO6
wCc0SC24BJqbBIDiUPNb8zwLkJAYkJa+J1T60ZxZMp0En7nAdypaVo4asEutebLG
CYCTYa7STvgX5e7cNe0UwpIOkx4Ol2jtE76DFVGXiE2y+/K7N4S43Rl3N8xv0GMa
mQlZNoLU+wShi0FSU5tEdOu6gcN7KQNVQKQybO1jrwFoVHWBq43XS8IKTNuc9wXg
8mJXQUcfP2OYnRfYcIswZ1U5nYG9hUDz96iMU7Lln69JP9SAFqt6mF/xNd02hJMl
bV4efIq8Hbax+8UiKH4xuWSTKrvXhF/z2q4R8tJNZpRg0zRMJKf5zYxj01O7Ckd8
QuM6NCR8WnjrVRdGMZVjllYya0hRUXUc2LzLc2sxZm26b+N+l16Iho1OLbG6xcIG
uSC6KB9U2bMj/5JsY+GFpgQj0fKaSz/iJT43sctaOPGkvtJGO+QMbC0ECkGcgmSn
U0UZJau6YvwavH87uZVSSscPKVDXyk7pltCT2tP2ZLsbrNryPJnPbS7PCcRqavCv
LjrdXzN7Jc0lvYzASxcJPWBWiP1FqiqIv8QxsVMEEdrZrAxthrWo7oC1Nyy+gsVO
oEF1Df6TUZqzgrKO3eDYTnarz1foU9e4IfTycGhNJ3zavzatVsR7Tv6J9Jr62vdJ
6iDuUlED5chywK2EohNGfRglVx61+7Y1i71Bpwafy5jSYBd4lsym2eq0RGeGa9rn
Akfd7u7+HsUkuRqBYrqeyP1zzzeHtdSxvkb/JPlKHVP0ZrTsOsEgKUMLSIfm8i1Z
eNluH5KW3s8ZZoPLTfwkPcxbaFxhLG2QzVFxl/TTVHvg534tJ8PuDkotiUzAR0OS
KpdIIv+QDaDy2aZ32rjp4dCbKvKcg8yA+Kle0XPKmTNgFNRufOW50zEnaaAdROzZ
TaKmt5aM931SrL5jaLzPjJLrK/tsn6FD+inrgmn3kRyITp5j+FQT/O8A55qln/ai
rvZ8d9hyboZyXmoUt6b1qJqGtXpw7k9w25mi7ZB/aDP3bBbQg1AYOw4F6HvQ7WSc
IfAnbqHa0GXKgiEhWq0c5xTUEWpimFZZWk/kGLycP7lclyisunux8UBhEeFzOdj2
j6Et3XpZQ9z5FlhGvM0OrNOgZlwWfswrXgZPfoTbahKRaqsTVeyac0cFjfx+S1nf
ZKlEk4aZ/+cuXjFqaOBAnBGh77MON9l/8cSKpVOxKBHBHq9AfKpu2Q7x999dGcE4
dxWYz3OeUinW1PUULj6wIghkyLO2YFsZEs4qt9+BL9cBcV+5G07DM7t2ThQVhq7T
lSBwBVSpHingXBfVyzZz3ZcBz3Qd8jN081g6dhd6NaJuO4wBFu2Wa8r85m/fQX1E
OM/Zj0dE3GkH+1AyV4rVban2uAft4CCOjX73HLx1k4SC4K5LZlDYArnjjEnyAjCb
3G7KvS5JXLFlmfKr4k4OxTtn1NLlbpoiJfkinM+dA5vr+KLPhGu2hc91OwbLIZVN
P0xCDHoWcRpXqkDMvJ5jWa4hQQXxxDIHUheycZaDZPnK2inmBnTw11Ntv1bToY3c
kc/d1xmBvYvM/AH+iR+WoZ/BefQrIhV3gYOflXhcy7A46JTbfZPpp87zN0J+Nhiq
6jwFwg5Qz3R+m/OiX+fUyoumQ2EG2Jc+YtlndUGMM+wt1pTGKwA86KXpwDaMfMOS
B92QCCseyk8qrvOzkJK7vqsPoCKRhCMS6atNCw3rjypbYnHyjdQyCU7rNwTf+RZj
IXDnBrTsjWAHwZQViNCST1FzJUlebo1BtcJHjRowLHpxXC4vFIZ4TebbO9qChfCl
uRA9CaXMyBXK3U9zDQLYblpZzj0ozfeLf9FNdEYwBumCRLkS6tY6NJ/ryBliOzRI
KIL3/zWSTLLBe3+h296JIYF1ti7JLsJL3j3lZKU7NhNiH+vMcLVwKf5Ft+cazsri
EYvwvWEVqUJJsMm6Ek98ZlF+zOfktNvxL3SZcpKwHg3nb37LvSOjcGV8W59nHcEC
2kERwsoe96xp4IkldVKE/gVNBL7nS/IpL5Yk1bpWD0MEiTSs9X5GsakLsmAXcwF1
Ft5rIo8VaueQ0Qn5oPSYw53Pjy6HecApLlIOuqrOQZw+keOzIr3wlyUhmHbasP4e
hfyLBoJ9Q9rQQnBvmPiVedtT5SVp/EQx6tJmyES9kA97/7IpvOqEbE6r7XHoVYAp
F3w07/QHgqF9N3j4QkSR/auZZ4PzBIoHTfFqShuyxJq56vgaR1SQJfsolylU/YxQ
hzQmHmcNR1ueTe+W+DrgUA27EOTIsl/LgfX+/vjhS+NOx8EZ+U6aiEomtjqPvpZ3
5yi2TOWwOADNBzDT+jTegegsfh6ApRfGy8qQYjxLkCMnir8BdoiwDBUBZ30DH+p7
HF3Ol1d+CVy1PphWJIrb4/6dLKI+50E9yFoHAgALyU8IJNRvnbnlXlWAxOeql//l
DivmI5xv8tQKS0n5mA6ORz6RGSON38pP1aofMjiIaB5RKtwHGufFrRYv2QFk0eDa
9RJU688TkDUCQOBGhyd/x2PLe+kivwK1CZKuxLyfAckaTFRSolZ3jP7WIGUdOue5
3GU573EpQTwJIONkZQ0Pvfh2MwUVTkImS5eorFd2gFKgDxhKFfAyUz5aGpJYieam
ikusnwxZzAaOAThCo802YSXWdBkj1ZtJeMk21xSn7Hp/Ge658pokAShonM1TPGaq
X8D3xNdnsgrml8bMJQNJlvnJ/zLS/A7l2ABejFu21Rw7/nKtgeKMtUH0wIDmVKz8
Njs4hl6B6yTFHT87ILZtqQM0tRkVBXH6Uqx2xfISEq7O1lnXfIwmjIVhgaQHxcHh
ax8ab8meCTbvNoWDK7mUMecOdvVT26rJO8v/uX17MunVSWGo2wt8mfL55DstMYUd
Qecq9K47Z9ZCrArvjGT+eMQoHREVLKXFBE+BwgXqY+8NUdwE79A2wFpdVJqfeXMU
cpzW9XrD0h8F0phRjYc5AMOsD+6eEK5rMdjkKPndgTx5/l3RsUPS12yY8FahR+wm
ZCLp4qNKJlxFIokyVBvywflbPYKumFbxwnDtKP9CAye53j6WPj9F54TOHJL8G3sw
wRG8LLX+J08aOiIQG202kIGpNSBbdK8ZqU7yAgj/VuqRt9GqQR3+7u90pw0zRbtf
tnGqkzUotTD7+Jw7iJrXxYlnrhOD+4WWcMsk8cP+f48etL2gWZ8SMgZ0nTDdM2wO
yfU12w2cIFh0zX9lvDCRg0FCjrHr49SFu0URdm4pYY14WkYRwpsS0eXAJ3MNNXYC
FP5hHoEupNgs+4kyImxiig3TyY36NkHT28IAG82nY8usWyOIBecqpASCIF0nxWZQ
lO/F74vX2mpDsCL+cRYaRjfXoaDS4K2Fcs3c1i6WZ+tsx9T5iR1+XXayxuX/FrV+
WoRkXAt3/D4NumGEPVrcwlwGy+fdQPlt0wytP65+t6+ZMwZORHUmYG1shwcWoMsq
STr/bT9E+HNzsYYGVkB1aotkdSriYRx0gRcFIEI70AVw1HtSKn0eAYByLEcyilo/
+v+bw8ulVIAZ0xGF3kw60HdYf+rrYGGaDrG1zFawm337m/TT+oKy871D2Om1mg/T
EkQ8DDl69+CIK6wi9zx8WJvRBmrnNeEHD9W5IzU8Yoon43B/RZQ33+/IxOcoLUjA
+O+ngw3lotGuw/uLXbdHJnbaa/tPhUL+Vzo4ngA7T3tl9SWpihOp3ovYqXEDinHM
yHDPdpVuAfIM+TkghuKnzdbnbE2/0vpvpVpCR0cOXfwtqHKsbAznGsz1WsKYskqX
ZzJImfg/Zq0aCaNBMdqHkQrc1ZgW8UpS8G5XCgWqvqiJ9et6tRzn1QWSbBIA3H83
ck2/DTG60GSz2om6rXs9AjtB6OAuu1SHLRgqeAossPdMf4KVhbYLW75hc/c/HzyW
Fr+tFDX8fHsmnjO2QaCu3aRfCIgKW4UrVN/NVGMI9iNOhqeo+gEyIe+VYa1DxM1o
5dQ7S5iGDvhvQVzS/+8qnRAPdc6WInOfCtZgiQf39kslUxxS0kKtgJLNYs7MMgyP
Zw+wKSgElM/V5EEkJ741PF4sj5QWZGYEyMR6MIOP31nTml7VW6ZTNe7HLqMdoo8B
nRNa2PL28QspDS0LK+a4b21eWD/cQCdWsFJAkQsNbaP1TWVm4Myj/HaMumC+EPI+
xYllHf2BCO8DV6Kjscs9esEwwKYnzslYzlK+0hHodr3CUSwf0N0hYzOwx3XECUji
jSQlyYjVS0bVRz2/QswYzD6SbzPmpc0yWTFzXkoYuCxdjSkcabA9LsMxBoYLMlof
2NFtRV7Abi8fQtl40bwzcBsf8ln7KudPNVjHVZ6YO5kN6mjeanV9exrBmAQpTN4K
MmKvLL7CFce6+bFcL0Q3Gt25AdZwFW1nCr+ifMy5c/NvVqrDNjiPOFrxcj30hIhT
9lnq3DEtVXH/k3d20k2tbAhg7J/IfrbFUVPvk7bWnPTIZF87kv81YJpjd88WG2GJ
gVaRtVOT7j/ZLHmxqfUivPD9ZRzfcZXiGthtyY1DcfzVll22VFbXqpZiWzPcaGib
3iBmjb6G0Ap+vHHEcSZmWgKv0a5+kb5DmhDhVH0bKELo9o5GKG1doey/myLZ7G8L
FgVg42IIc369/MK9zBHSOqspYq1F29kt7EnV8b/UNOQFHfWv09XEBXmL3xyUX2Yc
Z6gfrGtyVc4maBRVoboXmnU0x2wfkCnksBl/o1NlZ7iNmrvqSugPVUEO1cEWeKwC
w607tMcdNsnlP75JEBVLTGI8AcFPwO2tfqKqf/OVLgLSoPXnpsf+fMq4U/XXnEHF
P5Zz0374Xfos7uQwL/gjU/UmJ5ZHhS4bMr2oUoUYQeI2u2V/Vy2BjU1nsQwnfyio
sdK++3tC26z62sl4fN9K+jAmPSOUyILmaRaxEZh7INvKdRfAj1AKYH/8brVTZ2DF
LJ/o45y7u4m/Pb5pS8XZAd91jlvWx0FZWBj8M+cnObVVqmUCwfP4CgCd/ikk221E
Hyn3McEw2auDxK826T3iKxG9rBaWY4+Red261COjnoGbI9B9E5Dsx4u/FSylraAY
cMfWgNwHzyMEtw0XFhQCIfgDmFBFiPLek9C53t9NTOsixtMygR2JtzFjTs5GnoB+
duCQVcHuP279JJIgMoIjGnqN1VrajRqFi9wq7ziJ1WeFphgjMRuRARZXpbEvb14X
c0sY2vDz90UloN8Uezan0xIkWtKBDqvb6tGHiQstb/f0oO426igVG+fnoMHMrS0x
4z8ROdiHMKiq1Z/OwDiaj33sEMPyn7KQY5khN6avGmOhwpzj5qRZXjS5QZLWB747
nuplshEdSHF3HXe5iIPEsTAo8ZeA9Fuq1XbytRYk5/1Lf7TbTTxDZtZJ1NSi089O
CfrXZUjWkZrnOOYxRCeOMaeYAY3bFMd6jicX0fsKFUMya0/gxLcNWnZ65OtmCcSK
5YaabnAabgkyMVpO6OmNFmfxvaZcV2VItDRS+WEOSyZCHmNo+NeWmNkRDcP6kmvf
HvzXPMnOifLjfQsXhB2WSdQNIXEDejKQ91/PZL89LlbGAeUVjTZkkV+Xcj5rxQ8B
M0OmsIzmqPNak8NM2cf0vkBaLTBbvoLpmtBxZo6LPNtdip1l7QpyYJz+F28gEvxL
03zfbMy450Tbz1yePVjkIlLZeInjHCoqxrxOG53s87DaPeqx5ZxRLX0PS4POgBH2
EMwOxIvKdgf7gfmLFZpk7G/jbNxzEGiGvKzPQu6XlIaorSUOefAzgAikCWjolPAJ
b4CQlcl3h6ln3FdddAsjjEELi2VwcfVwSYXGcRSEa0mHhf9n3JL9R0LJFcMkhjQc
t/QknPI71k76AG4yWMcPZ2XwPffCNXPpUAtwKA4ZDZLw9SQs23brlfvCWofJ+Xph
PGSe8GBUI4KyshxuZMAMv62FASyDGxwoaWk0roks9zZdaFOx2QR43AMp0EjhUFaq
7EXEZOEJre144VUL84KDltB5c5kL+59HyDNCkhv2/SDCoid6XfYnY6UJd+mKi3N0
K9wzAa3Af2SjB36ByTcEBZHdmiq/c+2+3trdmqc1OEhGCQP2sBkp7jrwXHf8pl/o
ijOOyY6u2oo+8py5XcQrB5UTKrUmiLtagrai4XFFk5NtjRZmsM/TCxaUotZlf36Y
mHK141VSsY75Fu5y0q33exog10MbKvZ+ROPMeK3jPVeM+OK7P0Tg6nUDZKHd3+J9
BjAB9/BdZrfqjXCUWGgHsXEER5NvTgODbu2Vj4NfGw3OE11EGlV6cc5HBN0vCnmR
FNAqI6JeYZjZP4WJ6n9LjLUxWL8EKyZdspv5pbJNdBTzsXQZR09ue4AYmhSCAHa9
tbM0v/vof6V3eBW7I5z+7ZZTTzpOwrbDi87yu1fElAeWM6nSIsfnaUfW1KyEL2Tk
DA+In87ZLiTdPHI2P4JeigWPKKGNqZF4ZR012sjJ6R3HpGolUVpj3D1OIGD2wrEG
XvDA6kSKE/zVNqSP83qqYwbex0jdEPxV1x6weBtfko3asiQmYGfZ1MbvG7WIa7Hq
7bYgyTpBPgFGhWXZw/CmAgqS56eApuBopob8SS8NloiAcFT+RUxyB/yTL74H9Suk
/ZZN9KyeQZvYqIVpt1qNoTRRYDcA/IR/mOl69lafr/4VYl7NhvOh8dpLyxlWphij
I5IIYqZOdEHzhRq74lgmtKTlb6A63hcT3sXVTagvNV1yj3qECfBLOgxUpVuTAfdQ
HLe6rcouvMdANIN/6R/nbZAajSi1OEvgx47NOSJfp7sXEwQhjbDa95NoXRL5h1hp
B03nYGVpFIkvsjFqo3K286udimr+AglwX0qO4HHC61a1Gxg8s34qZODbxQhAzPIL
UOCDEuIDgS5GaX+SzuPY/jbSTWW/yWLUIA6H0t1KgYezQ6p97WrK0zXScioZ3fVo
yKdQ43Cv2DNgTX/roLGCZWzIs767ECYlADUlbTe4Ujeblu32cTkHQKQBA7fJNTCv
JjaQGuPEa//9dvAUNxQLK45jmLZb6td/sTp9uy5Xw61itwMCMkFnIUynM4Ig7RS6
Jj4Muk5NgydQaRNzaoilTB7caP0TY6hVmktmYhYLkeGSkQKMLbBtHSzxsYgG4aZg
5npHFY774/+C6c36ibaIQIS5bP/fQ/LC3uMvm+J7BObqMxrZX/DIWYUTWu6jrtkM
vFPM3UpwpeSg/PIeRv407Ct7LYluCRoT+yfymuYOYr25ahDTS5cMZBXVSXD3i7lo
JZSnQ8t2nzr5/D9zyVqvGqoC2OKQwnYsLkNHKxsuNk2IMUQwnsI+1TSBdBWSjyZk
H2uUevybspgKBygVqvT+lMZQAz24RjTz3St2s9o0cIZoPj6dwuXvkwF3fFbjn/uJ
jHBVLc5ZxKqmzyjR2qVVhqznajoqB6X4OqjlpWcpRgPPDl1Fj/lzZJi4iQJcsQdN
9SoIdhooPaw9Efx02Ay1By0/fu6fhT1+YcWE5nLxtt2/jVVOSzYSYmVKzzYxzOGy
Sq+2m5J0bNrKYKuoZgi5Ejb1919pnZutlKtbecozMuCTlOuC65u2/GgjW1E7qMGQ
wcsnjB98i+oXGB2kAuL91c3ymkLDZJ2Q8hC0mYqHfgjVsHs86vzzyOpEA3QT4SwS
olb+uJOCPxwpZz3wY9ow/wsNbxB9YL+HqoqaZThnVhR38tQrsGb2cJ+YYBoE+kf+
Aca2xeRHj+voD85Cinl9QxZUFrp+YK/CQ/M97U76w+W3oJaXzRVF0+OCtkVC4sYV
lY3ODTZ15b9GVihhI2tsyq5CavBWKc1LAjRnqwzGwuNVNez7QmRyd1QjnHBQaFjQ
N4CaGeO84Q9ij6Ji7UAk52qS7ey+AHsss+oIOEjppWik8Z+yxD2lL1lLbpT1VfH4
eADw6c5d75FzKOdUxIi5JlUrSbcyoj0m+csrWRVq6AEa50AClSLPFP11ykFLV4pB
iSaBj9FLVfKTDad8RtU3l8z4JM4nKXCfWFbrwVkB0TOXEe1/Sl6TUN3tAPi4CWgq
7+GqHxwdnMDo90/SLgTFTEcVHHZ3BDjndbCwwHDBYAHTlozyh2JWH+D1CslUjiDu
hJwfZfFSbLqMqs0DjEWDiYgwTQTcpMjk1qL9ujteBt25o10LtuOLO1hXXqRz1pv8
Vlc4PyFzyQ+FgwUazJcy3jHwOqCusASyfyT6GJgN+ixRfSHanne9YGDZQsaqQbVc
lvQj2XL22gt9K02yA/VZY791NYRr8nCg36LNF/x0Hs76WP2Hn70fauHLwDDV34su
F2BOMtFr8uGcTDyBFTgvu0rKhx/Yse7IjcNRsSP87gqvY3ps48wQTdQW6M3gEiXx
/+QCJZysBzrKsIpZuzqXyVfe4cRkwsBX3HvwPIjDOAYOevpjeXaX8VGX5soP4vfW
YMqKq0e7EnfRVLoNvkfVtEDxQFL5jaEi056pAs4+ZJAizHwuU7XrMFj3ABAyvQMf
AMey+9PpRuF1S1WV9SBDYiq8JXkhIjlPhnKnYA0JYpRHp/mPoBeMEUMBRFBtH/Ac
TC5NAy05k8G5vcxSoMMBKup1qT+/8JifowidBoGvYwiUPS+91JeenZ4E1FDMj9Ho
zzhrO9OhU/b6cMxU/QWRBsJUEFd2hUV8ZAyY4iQtwBbwQ2zesocu28ttXqbAba7k
LXRnx2dEJI9TKe4sFYmNk5kkVws9cu+dlugr/PJm0R3DjO2ulc2ETefHbtRLRWIU
8ScYbtiEUCR7syvMRSi+FdX3k8NOzJc6LoffZzMzWKQ693nvQYdfz62m4RdzbLw4
jbCkK6NSuOgM6If4dbtKPzvQHtTesrDjCMEg8qK5FygPHCTw/T5rf5Rf8odqVc4L
aGmdedSKqI/+6k2xbbyRnzQLH46LyM8zpDIu0L6uGkY9AKHin2ekaK2iSjUfraBe
oyJTR+3fvsPKXnaZ9MOMCqPZ/XT6f/dq0sgLUnBUDV2wSfixKO3MZRd5uiPq1G2V
tgpSR95yPq2RhSmncEUb3qwvWcxkmzi/oWzr88EcabUnuTP67vgnc+oJGlFpyIeh
BHwV0lZA1Y327rr4VveAeBxKYUSilXpQPGZbvvdj7c4R3AkQ59txkE4TfoXVOVGR
NbkRXdLKaO+9n0By43OWEp35K+/CMryi1X04voQnUTpuTBDoTPWccjutgK+FI+2u
gO9/G8Q7YHjHcbFP2fXPRCxR3gDpN9oapqSzBndZdHSMOvsKceClIEDZoTz3VOAc
J08hfgCtIyJ/3ZXTukE9pRS56//RCSG4BIOPMj09uALNpF/xWWSOxuOt0cITm8dO
ccCzKQef8qvrDSK8UUM19v1IPwBVkynSGn7E5SN7GO+53HuIMCOal76NpfmZXhoK
TYNCfyJpvmTlxxobbogwMii+A1fHhcHSN+S1t4nFv70mwoAcistOFiYozax4GWZp
bqxSBC9DCggnhLgNAecHbBrkaT3qXrQB98AY5BnQXYfPzl6CTKbWAowEdDZPwlvj
r30GkbT/z42E1ZElQpl4HL4efLdtdwhkb0K96pWAWaz1XlmjMUVqPKVgQDrg3CxP
N6IGTbX5Uz0cWUrgCu1WsyNsW9ebtnP4iIklxf2N6UkG1D7iDauttMWzY/XpbnId
Z7NGiGNsxBRpX4Tii+koaQHL3jDAykpLZfgP42b3dVZWPiHk0lr+DujitCd6L1pi
1sGykuvZbQBBf8ZWRZutg6DxLZlgN1+YbVthEVTs/nAYRIKmsYuNbAMJ/oNBMaTR
wH4VhWiV5rQyqquLA84w3DEPYoNZvER45PaZBsKBHSydLJzjD00UO7abVbUxgXrr
ANks4JBv4/zhzuEJHZl9k64B+fEp9Tz85fDwQMVACRTBKFIc6Px2z1IHsMLI0waL
LTNUi3qmPE7nkSJ+UK3HW0GDFvQGiScUnfH6aTNIFV5s7+APnLPLDHzeHmInlRE6
RWqPxJuB504L+ia1cLzyYZ8R6blu88GLjJzw3TNBWv2txkDhlbCY6Cdu6EAO3VW+
1KFQ7+MMAbe6DUs75YikYCBoHlll0dcHLHH+chrVzyipriPOGSTxaDuBFdR4c8Qb
CwSedJLUw6sYimnPxRf9OQGspAZe1Xil51nW8lGhlBy6YozdsZBOoLhA+MpchQni
4M4bWhJjRu5AkD/bGSwjogUOdxg0ZXXCNtLL19jI8e+bzVRnrb7GNAr5soPRNRCl
CyHO2GgcNrQTOE2q/QBeW0vdOPdc3cHI6lPnhp7LGWl83D8xb9MJyjv5wE/QWk5C
1Y00m1I7iHaOEVLt0y2tXHb4NiEpPof8TTMqQSiiaF9j4Hq0VxVLKaBmW6qd8HUZ
HDGTJLp3CgGwR3W7qq7BUijWKCyh/ieB39/Lp4R5XAkaZUybzppuz6tpildCMlit
6Riryrdx0YjnJ+So/BJ+NC/CRtJrE1uaIgIhMpP25cRF/khHZzriS+XssEKsC71P
UOYwWD1snzNB4h7/IzwIQc+9JMbgFd3+ynCjtdP8+KfUMl1tYk1kN9x8zj9AE1vQ
u1X4dSLP64mOMgfDPq3jgmcEBGBCaoRlCkrJVb7d6g13+LZS5pIarhWVaXzhcWeT
IGQ6l3L6FxjcApT84pn5K1zfq+CNHQrTDoQQaRTtHGWUJ9FLl+zIVLlSECFt9V97
vSUoEayAis4fy46VvFJHrPXynjnZg1TtYJptLjwYKA/dPsZtfx/gUo55jl5pra4q
9oQpluYWyUhe769Djly4+SZrqXtIuuKc1+g+h2fFCl+rjZ92+E6Ag1QBF7nwTqhb
J9HWf6TPiIVTk0mVSKLMUHjvhzHeICtlIlBqeLzvdceI2cZhvhEIGe5GIeEqnJyv
D7kLnAjoMjHofGFilQrBI/34fcWSJ2V8BY032ZdC+3exvZiaCbJKfaz3uMbj0dBQ
BqsO+aL4mp6b25gZJXpInFlDqwF6MTymnPTiMX3E/YMmxpPilCGWn3JaPH8A/KVe
HMDeSnweCKanbWSx41sGelQjnGjZO4oIVmnEgwUc7D+0YfhocVkw3uz8CZbKnueX
hLmEGmNJ0hM8NMXdn3wMDpq4MvLYmHx0IEJObaUdnxajOns1DYETrBxf3OO7NXnW
P6L//mktJQqRMFIToYYhYM0pRaYDJTqv3OWsD8yp+P5SncdmNGsMP7+mitDn/yTr
UWGXkLOyB+ihR2nvOyLjIVQ+w7Wk9bEWgS8UkoTGF72KbkXXF98UuqyIAbkiegUa
Gv26/euJFkiCj5JnRVcvMYfvjfRMruqLhlaD1wqbVk++WVvNFsPg5iSzocxMgy+x
W7FUkcXkOukk+ApF1qg9U9la7FR38gJfjWPpzjEM28oknVbkvnIx6LmcRE3V6M8S
zfPlYd4doVeq2mYqmP/rmKp7OlTrRzDvKnjvmUQS1JsDdGd+Hn4dOO9ZocRrRJ+l
i2s3912bDqi6Gc1YAvjB2Q62BhjYvoXlTN+48dwLoLQE2nacwaabh4neH3vzeOa+
jK+0bqjma38WOfphiKoEasitj/ncs5JFstDZPDKMCy61EaG6wAM/zyRng+5qX3/B
mXFVxyAWQ8AMBES0U+OveAq2y7KI6wdE0fTKqRJ2V/zrEWM+K9cQVEuzEIhxT1Xh
gQGSacVSJB8beXplqX2MgpDbq96JnMlDOC698PK81Z2Qexr2gLnXFJ2DGwngz9Ek
0lHaRWh/4qN0RbsXLjdUFNs209u3wzEryyBimylK+ch+ZbggW8hqijAodN+MS8wC
5eYMH8N+EdjurrN9zB37xQWClCSvqI1eojjx03EUncOuu6F23xcuNt1gvRNZnbne
b7QyoKPt6a2d1Cr7b35sz8emCwbeqEHXy29m3dXBAQJLZc6SSklx8Udhbgsxxjie
QpkyC/5izuv5mNK8MuPPqRkHUyCgonzwOhRRR4aCwaKWq/s4FJe2wB6L5ZgkGZib
F5TbYrErW+yuXwifmj7clFBTiI7DSsal7zzeiLAECMFl38KvfSIMKq9qh7wcOuRU
6RfGBSQF7QSdjKOQvz1UNtlixCARqEcrA+MFzztWlcjkVAP92KSamwzNIvzLY41g
4R5ud7yjAR+NNFLZW1n01slc6dBi50ULbELVANKZqnHxZZ1XQqltjFLP2AV2nycJ
8BpnOq3cHdjemE9QHjTniVsytSwvd8ZhSJuJOX+VG96+qgZokjUJjfK065KidSXb
eG2q4ENefvgSZ6yCSS3m6p41sdlKMxnMlAHrJgzo0QXs+CzWfHmFsowTpo/SHY1I
Vfcl6pAn7p6Qoq9h33Ekkvvc2F0oTUrH8/eOut59eD4Qnouox1nd6aKhdw2p5wD8
Bb9eXQMEOuzrOanpfZ17RfqRbJveVn9BVFZ4DG99DPhgjC11Og4z0m/jpDwwGnlb
al45AQEN57H1+bsNoKASL5tqxSMG4SK3dlUOu41dSABN8LbO666gOELcrXLhqbrr
l6efGVl1h+7J3wzve64Q7N4g1TyarzR4lAV3N2ldb2A/ibExS4qgcrNoOBrvolRb
n/hl4au0LF21YVdk4vSQiE+XqcBi3yCn+IJsGp79aUEyHKNERY/f0OJEw4NcKFaK
QWgD6es/3O/y/jjc6zU1MhNCngOP6Uf0D+NC0j869LclLB5P2gXr3sx79X/g3KBd
o3JM6ySLfm/qyQYzSDvYShoZ9aLpRfdiXvjufPzdt/Qxnb+2m68Obkm6XdukpRnq
oQLS1wSLrhuAAD1+nkLveq5ekeHemNqxoSqmGUOQxSvKZ3TpA+eN5b7JGY7/PHru
FlxJIfi5Bu0Rl851gnIMb1rq+6Ksi3b/iJWkgW7CFp0PYDtxsfL1g9ub7mZGpQPR
ebffp2/W+THExzE+GMI/ARL8ime4Zxe+SY9dCmTNA4feh5bZVdhcwkBT+9pYPre/
gYWeWWtxk8gaY/2OHHvxHOblvy5zkn0He7KlnibP6Lm6GprpRnDN9ReuHu9C919c
t82v1RZN6SlQfn9y8MUVzTKmbILCAVa+iNCu4ovrzeMWXx0KpJEn3ZBh8sEBvbqf
qXF7OebQketD9m1gmQDBf+GQZzQzIo89i7HhfCGIxPsQn3kR/fn8pluGnif8KK48
2r54YLOZe0h4AOxAMspTw84cYEBpRdxgtqJIeOiwi8nbjjCQnH14SMyCVkILRnY0
0YKbFPanQojZb2Br8MLcTG+Z5LS8mi9/6PuA0OBZCjfjmY/4s3VHkeJK+Wb3xOjp
ZEEpyvgGkNgUlwCPt6chJ3dsWXA6qA4y3OA6mi5ft4juJfh3Z9S1Vt773l37O4ZM
AYJwFPt8ygobsClwTdq6C2TM6Qcp0Jk3Dp050PXdMm5nPybP0eCMFYlx9iDsIgXE
OUDPPRh3SZhqtLUSt/qcscmeEBnsXtkytt0AGfRNSsJjHcjkS3j2qyoeCIU+84td
r2VpknPg9cw6DHbYFCEukeldXt12gEKvpOfufx5uf/zk0v/ci4XZL7FwBh6puHzH
UHmg7sBdts770nRrF/T7SniI6WODnczeF0FmoyLHa/NPBWINvZsXJtL+Em2/O/Xk
kxGejfjmGYTyCET7VS+jrS6XTTN/kArzMinHLhA3h3LSB8nwlgVEotwASnMo8/RO
I9teRKzYGEmEwoZSiqIbDNp7lg3Gyy/Fb1ZxJbMAIaN0PS9qHAyLSiJdyZxEIl4K
95MeAVOsWlf4Ih8jAtyWrtLJbH0hPzEy6TSVseyA003VWrjdMJOb00EtHKO8+A7w
yeO+woHwUfIo/7DHhYrA7N3PIGsQy7KhL1JAlAi5YSatpXSXdGUspqHMQnjbXpu9
FrGfRtuRpGfQ1oZCANC4/p5fvLfpp3nhcopcj9ZlQHifwOyPXtgO9JyFOFVYRK4p
7w5JNB1pjva/fLnCTVD/cVCeo+PQ7MaaTTPr/QkeZz6+VqJZvWxVGK0VIAdOknoq
xV2ZLYNLFJDrxEohfiwrJIjfylf8KE9F1uyJAH6s65ij95SVl5RehP7jxcnE6cC+
q/Om+G5Fpxh16vxwdp/B+W9Y+OjlX7unExVNhYKtDP7ms6Vb0T0D6HhGmH8QQReQ
WWBlkFyfXAsXCxFVEWvSQpexs+UDen5f85QXn1Rny8pzBRlnrdKvSyw2MqAphXzx
5jaT7A1Gl0m635RBZDsTQGFnh91YWTLaRoKAImlNNf3RLBwf2083TxlEW5zEuQOD
mD9M11hPBoYymLU8MRQ1FGgmXNckMnpuGKgL4QbpTC5fkY70Xnc+aSTLeqOe6R83
GrEcgolcQLSQgXNsYdzPxJ0n17zj4HlvVbJ2j2IFuXDxodwRMa8riZA5tfYELFzL
CifoX/k68Vu+tab5WBGEDLOwAQarhKUAk7zscLAiaUkDFFr4XKSi3ypYz6KYqlYu
PFpoNnBaK5FXW1qFOligdP0l8Yhb6pAz7WhP+F2XdEn0QVWQMUQ8cQyj3yRYZQpb
XgRw66NZcViBIASHcIyoxiiswG+MAvhH/J3H1TXqSywv5YgcdrS6mhIMKRIKDwgI
zK3pwPQB8iRTCUHExh3gjJnjZDsod435NzDeZGJudqk5QxshPN5Ptn2TquuK3Qco
TFuBtmmgIxyGlOh0ZbDGaTAreuP3U+nFigytND61BqYZL0V9/UdwZ9gVvbgezzZr
zj481l/5UaxkSMA/o9EYfDvWrRLJfr880T1eUwnVsxYt/FpZMsyJXguvq/cFdzCT
o9d8xLHtFgFeo3TOMKuvdlE4aSTjKgKfyXdr9w5YkUmJFEffgijNfsZ4vma+v11j
wVQW0gsBLW30S6GQHVJqSutqSV86YBUwSvYxML8DEthb1HWc3JOHuah6UPUHUMz3
3dVAYACvviavASw6kyHNjO0GvkmAuTEJv/nIztBz+h9GiNp7N0zPeOibRViAGG+r
s3gZZ9LLdWCSTYokgLF8gt3vc6oLIsHHQ2MiTxjIezedIpZ3vQjuhHcSqiGs+ytN
WwBn/zN5JSwGii++3/YjsKTy5ArLyg23khIRT4faHowMZErfBjN84ksXcF7ujvAD
z36my0c5rbHeO3qjhYzGAWWW8HtwG1zRYXGwc4aFuF0/l8vuGi+3IQo3KgbXm8bh
J2c4+zX/cYGz6c/9G15Mp5LIAwNu25qMsolmeLODPvT9D+gQeDkvB3ANuJBTEAIL
Yf7CVf5big5cf51Xdjoz/5/QV2j/2/ww5w7MoKB41q8tdyjI73PxozHHPfT0b876
GmiUJWFTKBVvtR/bhuW3yrjmPBYj2KJynecu9FiOqrzlel2+gAHreg0qYe5crjV3
/RS5Y6mB/TTRe0YiKddJAWxLHCvxhwCvRKdgRpsyR0fTmiIce18699MOFB3eA0hg
mrIEj2CUYiphC5llfBoFoXootLoZZ16ziHMgD5EQz0ictpFs+MpkHYUUwdIaysXX
GPJyUZEbNcTnOLya5/Iu2IwQl55B3qKubjAyms0gxHc2FJsCIcjGppSeVzNXewr6
B9KyopXobYBkeeCb0wpcUWMgPzIgzi5LcaD6QpIGN21Z8SIp+GgHvyERsYO/lFOC
cWGQlXt+7XyT1A9+AuLqT8zd4DyVGCwsS50CLrO6/zwP26OKnGDFCnITxjPRAhmw
PkFakmusNuLeIJw6kMRfciQ6LEB1PuuOisPTn+jVSztpGrFcpKbLJ1IaVFjk2e1B
g91WEj2guWcR00vKElkPDahQGg72K6TF8Jued16rRhZuqBAFp977ZBxu1PgaZaXA
yN8bi6V5l7sp8sIASNkhk9B21/hDh5Zs8sVzYAkCl0SRrhjZi8zHG0tvHWkscjiP
qQ26iHjoatG3HBDYuYI+Ptqfs1GnjUNiX0rPG6HH8UqjYEPPO/LkQOy/k4w7JDDp
3NGZOzf4ODV1166phWZqwRgWgrnWqKlZL+xTvSIusJcK/iqcKnhV5gCJyg7uGFEy
Dl1tqCf3BjXH/vdt3gyyGcnbq5hEU6WWuAg3ZVbHOVIuvG8K7hGeVukAwyMv6q7d
smIUevHVGJw0/0imjI2I+izF+dH3AREKL4K8bOTKQ41Aeclwn3bgy7TDWl+I9X4t
1fftJnL3iFZ/KpF4sGZX1+omT5Po6UE+p0hDZiLt7Zxi8TYJ9StKIQjipQ5gp173
ABuO7RmM2VvNdF+pfcvlvmfM5KBxp5Dy03QNPFswZrkycWxg6npuuCqZhiLhSnEM
AX/A9SpJO4F7JjSnTMKc7NbaJPfR73wBhJmGWusWZ0haEvWf7WQ/GJdvBgvMM1TA
oVssfy/X4twq5q/gMT0BC4yz4qayOoBWNKVc5821vPpXkYYf1ZnFobFWHEOHpHoY
fxH8dRfdvVfPaofNZSacZxcqFWA9mYBni3v+M6oSj1kxe2k7FL68xG1k9l5gTGZH
9JeHSlZC4mwuujTqIhipsHOxniSBBSGbmOqSPt2/2G630kHokE936kAXNu+Jma2b
rpZrcEcyPDdLm6CWz9Sl07V+T6DY7yzYQPK/3IYn+i+iEXuBNPjcd7RcReALe1v+
KxDgAu/3jE2Yzlu8izOczfUdHUC+79Egx+gTm6GoLc+0k5UY6BSTr26yHM/L1ewT
KTxpQ1dLdC/C0VC1Vuc/HUsUMXnWwRzKbJV90t449NPrKQP933mf+RpIe8BuEqMj
fsewg5naDqIXX04qd7CrIpwTN/496ANKlsI4P26k0NP2M4hZsRuf3Lt+/ea58MyH
lvf9Fs+bkgNYyIAGy42WYL15SflpB1GOInWickrC0mSgC6kwf59I01eAbZcnnnAV
Sd/LbNQbFpMKb/SlvP5ZX+8ggT221sex32OeY8XzsdaQmpETEqnJ7Il4XW9prQwU
hIO+0/ZntDXV+S5asZR2s9SNlR9lNO5HxDA5bEXFjOi1TecxTkxWKEoCh6vEJkJ0
Hy5gSyjDQbRo4ZzsOigSImMKRPb3CfhqFR79VmppNlr6HHvPIrMdtLfKIlRwq6um
xxYcpjiYa7tzdUqn0UOyBz6o1VG5+b5FhvGKYVmfykCkJ9rx+0RcVztz2uQf6wpQ
DC8mKXD2Vgs90QxF33J+aqIAwryuWpdbKgXPkqDOncEsBzF65U5KaSqLWWhfhA5p
N2ViYsOujduN6OiQPRum4P0carQCU94jMf25DV+EBxhzUscI8c5KTQMoMHkMLKL4
vjSk4o12mJZz/r8BWie5Kp/D0CBtmjWVH/DpSfrqnizQvoNlg4pdVp40go+SF+ZA
IW0+bLr3wE7ByBSJsf99sMUZq7jWwy35BNPafCfz4AYQnF9Kk3PJ+DhghvZGOnoL
3EWLm8IodBfDPp7f/aIyWFBBQer6PGiRp7hHJ/7Pb80yxWpTjWkks8H+krQsnetX
tLyQ2I7gmM+33DQMF8bgNdq2a8RJubEAyT885gHJX9db/B672+Q0i8Snjhd8LTk3
cm3RRch9rgZKu+QIzIZ589LxFhFmUjTtqKQq+0dAgg0/gUJaKpb7ghhJQD1isy4T
n6W/pW8g6FS11Cw/RusV9oKwX+8TiRmMsObeIuD+ac1WRDyB9M5Twi8jatKtN9vQ
KpO8TstHpLjr55sq7DVDcamcDSLQ1GPOP5NdMSgmsh4FQq0etWH3fp9GAO+zTQf5
s1kCiPSGbGTmhg77P/7Su1PGVrzeAanj6cDOKoGvgjFXUatxZohhEwlRNCHKiCWF
kAnSsynIbpsDGVj0x3M3jSFdBOVTrAsZBlKGh3AqjPSVBpowmePSOuB8ZYLuFSgE
EONpUhEAVR9pYy/jrAGmr8D2oNN312VvNgU9LyyT0/s9fvJdsbIl9QTq2kL3r9z0
ApriYCa8p/Mivb163K5YbzfElAfXEvoxEa3dbyIWdTfUAgyZBBpPoTYywK69rpXn
PSO3gLnugigQ41CMATe0t0RC5cujmw6q/DhErXEln+zjPa7ScNBsWj+3uPF/6KYT
aTwzCdVBi0548xfPCIuMTMLnmUxFooAKQq3nrE9+mo9tT7EkRLhaXWcg9OOgHxRj
U/L9jU73a0aADyWQAch9x3z9uzRDtC/livNF05IvDRDrA7XGJxMuF/NRx1Jqw98Z
TKaittlikOx0CY1vp7ihEEHQqDL2lxV+mPKc1+H+5Lvyj0kwcaDVFqFRSRIv2Isg
Lu8PYS5shBQgDpuetl+2OCrcyDYBg05p3+F25Y636Zk5YkVj+nRP+rigYF24wq1k
mSvuKXjE8hGqRfv6gqJMVz2kB44ESBwbGDVlvu+tZ9V3cHkrxhqPSSPM7wnEZ8Xx
/AA3CuKoi7vfK1xxJdOA1hPUWXSW5f6viAkRVayn8J2tcNvQJr4cqXiOKNgxWy41
mEa/7va/O/u2HnDWQjxxB78HUbMoYzxS9eC0eVEp9TTOLgnFHocQvR/qI5EV2sNW
dzwxsd7zaRhd/Gu8fk2Lq1qDIsuNm8jfj5GziFAj59MLf6A184qW/k1qodW2OtXH
4Exp4KYwzFvCospi7L4PpEuaHsjVrmuOULN4f6N1/kyLh/bRTNmtU7dRwPys9rzI
tUwXIErhYs84ZnyQdJF+SsshQ9BbN+I4KyyFoUWQa8dJPCETeZM3gVVsNu/exX+k
7kzea0HEcGkv/Xoqkx79PeZXHmeqY2qe4IPZePm3wL9CejxbApoiTrU/KhLqpLsi
ujPrZPLTYocxJ1fxrOgQy9X3QdZmwTjJJbOBXktbKk0JClcfU14h/kX/XcmyCgdx
oBO7gX9G/Ms5E2w8H94CodkMvptYtfbsy6dYb+my5xfxBSlvPrfFyC6wyi3HbFpd
zeQjPKufAfcWRBR901ygnKylQwmh03N5l+Pt23ZyXiqCESXOuCKy5+UIgSWvH1gN
aM7EzFI0oVHlwOfpR0F0cLv9jZsFUebfJM32P1w5vAqe1wwig8sfLw+Ys6foZzEQ
ZKtAwT63IdxIn7hMN/X/j8YaxpgiIAhzoZ9L9EPcNVpEmFl/Ixw035F0DaRWPrwy
0zVK4TEyS4TOeio2nIi4rD5/slHkXm/u1Na9g7+uT1kEtxw5PcRa0ICbKBx9kaW9
VVg1M6Omnfd1WdGsYRu/LYbplRg+LzIcohsYs1mRTLmqWnh+p2VHKTaPfULXSRO8
xohIURJcxRxYdyu5tFeyXZOLyZmN4ZVnVM8L+znxoSHHjHzlVyDhQLZktX2gSghu
MBP60T1FaKsMpJSoB10leQzFcSZJOmbPXM0SiPRxR3y0fBLN1w1P1p41k4avvBrQ
iTgP4+yfDAbhzz8tcxBMg+FslkHy5Kn9kTlzLlEx14Kh2d2e+LVP3Gw0J5hJjTmf
wsKz30AaqKjdiuYAHmfftXLMY25lByd9mgNL/oz0zz9fi+if9wu9oNxiZ7YA43TM
5F2crakyunJFLQRAjqJXhcN7xSsmvtcWwXgSdRoeP+Ns/ndXy8K4vMr9G3ggq9di
wBgAY2zwUEQURMPmFWgrh1dwD+7cbErTZw6sPkO5g1GILkfn3v7baaAJdhFMCMRu
o0n2LZJ7hmM+mHzur98ust0eoBcYHZJM7szOrhBUOevYSXVOd3yNVvJHJSOA4rgz
rX87hqXID/DE4YCBXXoOCZUHQzr+4zzfAg5owcseTfOyQkNbZXwZv7GIkwEvYnWH
LYuWMICXglWP0d1lSieKiBrmiaYi5w+vkeCvZZMaXFnN9RzlHzqNjZlTF/zlL06N
Q114rniEXufrbRl1YG5LBF6tS5ecsUQ7rcNUlSPutf3/g81M15AYI9IYqbpLdmWE
pm32hE8rjN8PX44QooyfOEg3/langxvtvZ77QGaQZQVpnTNjvKFHHJcRIr88zGRG
/551jd8Pc4BFDPpdX7rT4OvILsnTkAqzn5Cr+v/xgdL8HTPS5WIyFDJZzbP8fGah
ooYYvacjWUrpozXfXl5d0o4lzJlWwoz9AA4SK7NbHFOTHg8pAuTPvyXMOTn1HMuz
jlu9dAYZBe5pAcG71/9TAvCRmTZlqMVl02Hg+s88OZSPs+6alKLl9jY66j2U1Qkz
yeZc7QeWP767krpMpqpBuJ/CbwkapSkdddwKsJNq1VekcoXNNOuHvgcIOq/wo9t8
TyRZlm3v1rdYJF8qcV0jhBxd38f1mXTq2Rh+sC/UhZ4BTrPV1qOUqNqA0Ll094DU
m93fDDXIpT1bBpxfMrv1E6AiEF7WFOcht8eFszaGGqx6riFVYLf1e7jlnOujeqNE
wDhIpzB/9gQ6BcPsJN6Cva8qp9golFhXohhAdPm2jWxwWKKUc1YD7q4jOZQ6k67B
a+28v2quAJYnpDx3Q4OsWpJmxGvB8kMvwjqStld+vNJUeFB6UgvSkS91uNLSGp6o
oFe4aPKrNEcdFLpmabY8VirV8l04RTIQrfrQSjPkxVJ8cPUc6aYtTbQ79+D+VuO/
26yhnD6YCyJMdRpSihCibd7P7Lp/+0FyCcNRHkqvCOVPgMxm/iq2HPEQErBgL71V
a06vGDp2cLx4JanmXywMPgXda/8PqSEc54xROHX962iMV4JLCgzeo46ArzQyVEtI
7++JD3XYmoah+1t0LfBcX9stwDREh5X/2xxY5s9UqT2VEiJ1bmJiKJBVFTc/zYE+
0w9qz8cFMMLGRk3vcdnqM0KTVkLFb1eNo0SMQBQtDGf1/aoIYyCg3R0nsSdQ4j0x
zZ7q/J0HY7t/s1HWsLEO10jQXsxoHhhA7Xtyeg/MNJW/Rbqinx7gw1W2QwoiUyTQ
rkZN4HSK9d1gsZTuWSbyVydGqyLyGL32Tk2lKnw3PcAjJ1C2gWTOY96fgkCQRkmE
GF9bvsoxgU4N6YUtHOZ2NtezqW121G9oGFKTbPe6wgNHB45lW45NMYw8VGQOeFBo
Mkn4QjZqAegEjoLD9+OHx0vG69dqMmPMZvzKrqTN9HSy2EPFxiL30+Kdbw2l/EA4
zbhbnMa63+hS+Dg1WS4EB66eDCv8+o3ua7s/+c6rksMqzs3MOYAR46XkUxHfsvyP
gGHyOt0APM1BN5/7GbRw//oGb4fSaBBYeNbZPHtQLPDczMM8UWQUnHiUR3F0NQzl
LbiDVP7IeqVXJvplqyTJSbc5OzUGCaAbWciXrN9C2dUeV24urJ8NCgZL8pjORohC
Bof4SxXgRGork4YImvyQyeGukDble6Wx6ueWaz5VEhIBIJKCGs+FG04i7ckhjelv
lh035IKrslvChQUBkYuMTQ1iPprQUgnss3q9NpPSfJb2hRlnYxGq+IftMNHW9+/T
1y1VVa7/6nt/YD0fa5gP4jEydpNq4GzepsgF5L7vgHrALAg7VqC8olBEVM4VLxZY
vEqMdoMTUxIU6jew7YbfBwmvge9s/thDkAdHXpsno+HS22PYTDeGz7u0y0vgU0yT
uSAO23RVS4U+7kBHqiC1Qh3F5g8AaZVZ18xtEjXr0306lAY/Ls9wVbQ6PgAq6LSy
5N3CxYXuuYxRo2tb4NdJxXIq6Z3pimA4OboMbWsDJQKfx+1V10XcO58mALTfRiUw
XB2Rw0NoooHz3XDbkzPptVQkFUAPxmbZgR3ouqW36vYw8DY2qH7G7EFQgALQNP8G
tGkmBRDZBoxJb0fCjPPr7Tx+qVLb1t1DwxQgT+GNR4zHZaNQORvFjPJeZYqYcAyj
mrH9mLjvoUOYP52/oKsbdxLftvs/HURaz1CBEoAJDHQNUHo92XPrEoIWmMGYrS86
00Qw5XJ7dbc0iLV6xR6DtEgWnw1027zc0XuYNGuVHMyeIPUgfqmX6y6kZ+gTUeUb
weRkkO1RiSVUmmwIarqF7YMt+ToHoSKgkepFuFbq0xxPFoft7f7SITGYLSp8hpkK
eN+BqIxItvImqxNAYbGYCVUMKOnpwZIJRDB82fNlf1JaJGwGGgldEPtCzZAseX/1
JgX+jz/HCipTWwfS1kNbvQzT6Dh3yKjyu5E/U0yFFv5D1RzMWxkIAf0TdlFRF/Cp
EmBGM58M6emk3bwC06azx2HsiovyeAIWmdR4eiHLAzum92Cdk+Bg1VmxR8dk9aDo
MfN+U0fGE8ZV8J6V1oHMXD++M5AHUYo02VXVcSUN0KIM+pmyLycMb3SJ9rLn3Hml
O+yRjK9hubQU2PBqHzBAovlGxWtsInwaV4VYSWK4gVNeUmFcHP7+tlaJTLu0y8mi
Hl4wnd9cZJMjcKamGHTUPHnbcnvqKoqgjwwcnZlFqWjOUPq+JcZjN1s172zkYHN/
scPHuHt7I2XL+0W6u+USebTOQpZ72lQ02ejKugAeUJsgsvKk0ZQxCIegauGZSFhC
8ZVmWKnoFMtfq2MI0EzRk9D9SJ1nRKlkTBcFuPeImzuh59J1SI2WY3mhNKC4MMor
P8OY27qQr1F9XYn78oL2tPHp68HL18DwOFBt58JmqRVMh3yyGJWosvY3NfkgTqMS
+iQFTLWetysiGR1JfgVupDcRiT07MVd5VyFvlqdnxPd5F5w4unn7tLrfyrM8yzVt
uRb5KVEaimzFVpyGJEoWcyxlTnesdhlOGHsk/klv/n8VF/O6r19RPt2+R/3G/Emr
KB9fncYlNJkfBC72WwsmH7Opn111Py1KNelDi8hkIm2DcRkpwUvYNsVUu0CPRwUL
lvpIJ7kIhU3j+EZc2Vam/GVXpUQSWeFxO0SIhNEIEoyX1cCGF8uVhQ/cIcy+FNkF
qCyOhEYXquaKyvBc1h8xXd3Q9v8bD6N2nwRp/JvyDxeSZROkLCteBaffm5Zb7RM6
jB1DlAHT9mppnirMze0e9onPigo/9xFZCh3qFeme1Ke3i/ACmI74jc4GZ7cu0OwK
kea2gOieXmC2qsCiaHUZkNJMvDtlCTVahzmdlYlXBT0nqieOgYBuIZqm5TdRBi8B
Ju72193qUz8F8Ye965y6X0LaHtXWVJCUeIpgb4FApFnPPTHFMuevlT3PqVCjX7OY
g0dDo7SOMSrCxd+rNBLC80v/67HqCgE+IJSMX0mNKhO8bmHJKMtpkK5xgN+m4GwH
jUoTAM/+CD9UKabYUFPevzCu0+/1cmSTZQFAuzDiQE1LJEZF5qMhiT7Me/lTg45t
PY7ZTG5wk5v3webeWy+9mxxLaqf1gpyD9ngrtUPqteiI39digu6aLNF8tCsnovjr
mt1BlINurErDZIlm1PqYjrliyRVWnLNCCmpekD7QJrVCF2G9wSnDOxrubrmbAjP/
69TH5BJJzV/KIM1LhAn33/znnVNhoQkjLDU0IHyZj81sYH0+pedY2fjylq8MNmwL
N+2c5kHWnnRCtXBkn1qWPKlA3y8SlnlK0l+9Vd9wzXgaZYmvVEKsXPkAr/5yDk5J
lSHC+F0VPDrMcoggUvXWUScoZtUodsBIp5p7FZLYHhhKORZb7SyqjIlsFvP+nTCI
dKLM2FnTh3lJ3vtoBLSozxFoc69bBOyfjwrIo5RYG5v0k/mLOD7EHfW7vxawaUrV
iUe9XEdPI57Ittny+KdHdQOiADvR2a3EwQyTieOlFWicmWPp48WL46NPxaFlbm76
4AUceHIPlbkjDhVsbYQa+47EWrxJeBJ8ASOYz2YOn9he8Qmvww1MfYorECQMWG+W
Y/RB27NpghsXr5g3Ar759N9mQRDD4Wg0WCDNq5dqgATzUH2n3n9L9aI7ZD+ggZV6
tYJyloONXe93PAOThL+ahfvgPZaIRC37mViT5TKfRZkMEZ3gP3eH+3JxgOPbhlSe
dVVSk5+DfcZLsvDtEXNOfknTk4FYSKE42A1OV0UQYr9O+tpRmkSw1Zm65Koy4c1O
sdeE/k8LUcYrkICvu5UWGtvO1Jvy+1jaUgcB5BanZ/K56GxE7unfvBzxHCMz1FEH
OtFMGhqYEFUpR1xFnKAiq4NlRtIsJkS8lLRAroKDXfkEUnQMQcSOJlxRplx4dKYe
OjIt8b8K3G+s/wYa4G5WZasx0qdB5v7Ber701miHPZS02EDOrKB1fwKUzwqTJlow
RGzOUoMBWRGQGNvuq8lbT60FRUuUgFtvUhxEVkO32UJKmTvMHKbBtVY2bXF5blfc
7JfLNt+GSL/J3xt7GSEuQvZrVzoB/IUzp7VGO+NWMggKQly6GXV8Qt/ZAJwEqWQJ
/O0N2O3FHKRXpt2W+9TMXkvj+oKGQKk1rGcR3LUr2vAS9Zp2ZroQG+U4wXB1nD6g
fctvApu47p6OlFJh0whXGF+kBFpYQwaPEg07ivREpE1VXcTWclDsoYnBfOQnuolG
SyqBYrm90bopgm1nPPbAMg676p/DxDWoeJsQ7FzRCANkfECSFpEgwuy5wiYHDRuN
UYEma/ooH9mNb1X90dj+wblk6DmgumE2k4KAznahKrwvJCxhSUhMvTJ5lgI0idH5
rJ39xPcWJNW/E6rYcHY7xhgNmmw/eaMOd+A4SoS8GjHEkgzUcbWI0DBVT9onAw8Z
Un6wuRD/TRF43+mIDTF4hy5vbzw+yOk5A1cL5vmw6URjMp+2HwqQBNbkaFvo14WY
uP2NkvPLOuwucEU0b3S37d6YTYUS8OUjiMbMKh8fY5tW/goUH3pNi5LZWdI/rnly
Dpb3Uf1n9R+v55ZFfovk7b7Zdq3j5f3fZI7gowskV2nlNWmtw9b1MRCs665MU2w1
XXPx6NGC5/ZXcG4AGjwC/wDMYAuKL8u0MJIHsh3JzOn6wuMEsE8o7MuTgE6/X0ix
gZaC44zNmVuxSIRWxBLyEdNxQynn7Qtobidt3fVlAhGxWPs88mXjbUB/aOEpRGdJ
o3zoz34wUGgTvGFT2EyT+6yCYPRaoRq4BTfaHOGbE+o8knHM3NXVJQjrXLshAf+1
XssgN+6hNG5st24cRyfAfgpnGeZssk0NGbTa0sWKpJR2MMtGZQrvaH+vKnZEm8qm
U/PfdwcmNtpzGj/T/1lFhKXedm9bX4729GLTObEnUt/jG/0QzqaTyhAOHfszcT7H
vAxMkbZK6l3pL+BF6dZHuQglZWcl5kTLtiYZrhH1BUsLYALBw5+ZECFFTF9MgSSA
z9fSp/J6ZpU3qXFiPToWAQYRQrx7qovdUc6RmWvu1GQumjEDriUQhp/rhPcCv0pY
q2AcbJqlEXCScenscqvtKJQp4gfMbwwWNqlfLvpsVxqDVImZreX2zpcIDJmqDoHu
6hcZ1gKxd+skd9cZRH1k6DH+z8klHtuKTuk8JqBCw3IdqRnlMbL9z4srSRp2Yl0i
z8Ur6KNgKtLmi/+OTqUCRS4XUdyR3tUJB0Q1t0HGyLFuNT02eY++p0O85ckocOWQ
NBU1OqHeTO6NV/ZC6OZxM6OlPceSXmprMLKAa/5zfHMFABTjA3qs1KNoqf7zM5VZ
paJH5Je45MJakAYhaFI39MyLp02R0RERpyiIrBY85APBKm8TBSGOSeHKYZmF3LiA
9Ap2Ahrgnrg1Qvo7gVYhDQMv0a7nYE3A4HWnLDBvsgPgmXSXCgNGEG7OeXr48PnI
h3Kfo7yxPWB0stw8lEm7nPpbaAMq9w/jsAANH0Kq6EP+KSAQ0YrNfRV+L2BtrX6r
FWW+a3/l93nh7Fi6DuMs6nGE4dSQA231mSDJff3y+njSTSALYP+rZTMeUJLI/EeL
o95qzAJHYY5+kFoNjgWx/lUd1fcNd5BzChvBizDnv0oBUr3vyQCXhfZUpFwoFCdI
WJnVnPElcW6t+N84YDA6C+2tAhk14+1FJKAcZQoeLFWALAdhNvmF+0zUPJWwcNft
6g3UuoaiuFQZdq/aCqffYXHD4CQJuZdId8nOlDYnmw57Swodr1mEYn9woQRctkX9
zUseDECVqBBqhQmMqgq2hRAuxvzDQBu7EPvcEx6rmPnMdioMaX3OX/olzqt556jc
mdU8/OLvNrdVS19nhqYNQMxv9Zeo/jPDZo18YDPgl5k8i0MjLrq72tc52nC4TPA2
Zkrmghu4lNAPU8AJ3xt07yR5cKrfcXJ0Zpcxgfa9F6oLthOAyaUXAGcTjrCX/tIM
TfxlYuG4XnCxK0IG3FCL1dspjqld1lykx2n5wLmQScl/A3/OgZf+Sc5iyeX1G3tz
bYt/rZqXTpO1/4mW9J8Dffdbd6JeuUR8yPQT2PsEGLloB4Zqieu0hYCByInl5aj6
Gs0yJv6tWYeV+DncEHF9WGCY632sTOrBIDYNqwr+j6223z8aIJVsUzhNFeAWYjRu
0d2NjQ037AU5McNlfnQ9lqJU4YLtkqbDUz8CdpJYcvOh/CXpE0/cPiv/4QaysAI8
Gbyrf1oELCkPHyvvHL1KOA0nC3JOpsJtySR/gdV/Jrimio9nXXX4nB/pWDYIWL84
SuQnB4aCsR70bbGn3Y8RRE4h9DT71zsI7BjiSsDs1WLJgp9uZrMxczwlXod4ssrN
/HyNObAGSNGUs5mSE1XhJhQ0KmzypPVYKQodgDaUTm4mlPPrLniJv70woAgUbnuy
hWRV72kHR5u0p3/zLn3C//k4h7TgBnWp5ulZVU1Mi11q+J0BNMPAPH25F+6EBMTT
kkQ27yqC+V3ZRdVlc704g1KhI2agktIwgrvWGkD/A8pFjG5bNM7W2GGVtFukHt6a
VzXfNBTuNNeYwfsvYzf1Fg+UYrP/AYRz5l67mE/qSo9d23tJytRTFtMi0NMxAZL8
jH1S+1k+Re/JlbA2ziaiVa9A+RuQD7Oeu4zDBd0mGPwCVxyz2HhpovpSnrmDS1gk
abywQuM/1ZYKSoOCTchT8vtN9ACtZFb4OOFQnA2KC7QW8iglKKfxXL+Y7v4Y55Ci
nccCtvvo08gC1vXWXND1n3lP4uNqRVwYNN9G0R+fFJ0+jpGHnUtd1PCc2ARLMYVs
m4itR+OHk0x/UeM9YQ8+VLHOdDOdoeVwvdNB3tCQOPuu1sUTF8kLTQbqxbHB+XMB
S4b6njyezWtSEvhW8xD4eumTqxcOhqGa/RJdGFIFiheJMvfwPDqaAhgqSQRUMetp
p82xoaCwLGLSx5J0hHLbbK++AEpXbyFWb0DKfMDRxoJP6g7GXyeLIvgCNdiSBtxV
8t4Vq6JMKDYIyYyxESwQohFyHS5TLyKTMmLSlA0g/ar1DkDKcrqR0bCz+Lyvs8Fv
EIlVB2Rn294vT2/r47bBYXUIHydrS7pLnrCj6eX5VL9v5BIGGoBL2ihgbZFyIHdM
xyddM1hMuNqzXe6j3HsblzjeqPxmzoeDH1JdZu6VejSzG4czuDB1ONktDInWJFml
slFCa4odcAVsFs6YKlzSL1ays2byOcqkZgXeZ2HRplNYX57dT79e/al4cvdIYub8
45fywcya0GqHcDMbPWuutmzlupiybnxg3SI2lTHBVPFL4oFRESIYZVZ9cYNgHi+0
GyUE3qEUmVH3HMfmuTvHz3qJcnVIA4Lap09wfDV7fHA/mUTyMiP47NYECID4DHbB
BjYCG5SQl4fBAHJ4EZNThU3ai21/nkRRQaGNlwR/AZ1usJyRNjuOF4HzFnE8mP4O
hozOun1TKuwhUvJrbB08OLGKkdeU+HqAjQqzLbkSWR6hK9+tSmhK1bQrIWKoOMdI
3PxWqGOVMW0LENWjdvCqHLGpC+sUoI3wy3zUv2EY/a2mwlxaHH77PI/qApcjbDEZ
ZkSL0p8T5uKGk2UIDVxCWZdlG/Bgv8uKg31hJ576rhoQg1cwr887LQ90IGG34VDY
mTg8fJh/Lt7SV46+5DC2SPoDRoBvWji247BScGynkEnsGladeqgvYFixZOF+IwJm
8Lw2PyR51BJzVbjEIUewFFVNcENXauMIbDIR9DzEUPpGF7wqOgm3LWI6rL1RhalW
N1tGwplTL/4y7s0mrvIgi4qYL/3b0dnMZ9IA/YD1Wq9uHslh+P9Yv7XTwoHSq70K
nYDAhIAmoJU3BCx0nlfbkaoZnC6qAHfCe6i4w8NYbWvC+aARst/2nr2Ec3hBfEy9
PdKCN8DZp8U8tC6E1ym60WPpe+fAsRNsWssccDs209BKNVZsRMMdh4ZWSXIpCv4U
lyjtGkXeTzkllEVNEIfbWCdDe7fMez5E08q+WxUJqsbpp/T+KaIru2+bWiu8oYoj
wumyb2vfz485z4R7cS1CGC9OlFPBnk121GUwqk9qdWlQtTQjMGuhtWn7Lc3B1NEn
wi9G1Zn6a2rjTfg6ClpJSV+nMsE+G+ryutpULJ91ceuv3LVYJLS0fWrlqXncTO0K
MMo9HArJoG9Nf0Y6FDdCCHRyJt8FmEfShDghOIESdjQYBBcYYRG7zxcrTLJmcLZh
mEqwb8Q8HIsBkWitxqpnttFWMOFrUK3cDUaxfUaeIySUbSjHqoikVsGcDe2Ekln8
/bMIsJt8jYdwbUqYvkd8WLIOQkXY1CiACwbpG+1RosIn2PjrboGcs8RHKKXy7kR/
kcq9ZAyN/8NLxfcAsLKmoU3R0xPsDQ1WD6P1F4hU/wwfkHcK3fVoLeS2wsG+vvjS
EKqMOJ0/fVvSUK8cEYgNxllCt/tYLZH811h7xO4gBphY8Zf8CxjtjcwfIL2+n+oK
Hn2OlaIE177ScvrUnW1viOr+NyQ7S58Kj6CpDGuJgIlZVyG7n0eArn1dLAUbN7uY
cU7KWXo+lFE0NKdMAwYO+R2kQiN/VF+gjxY+/X89GXsOROO76Fzbc8ccgqF+ocR2
HSCHykojGIteKkK7iGPHuMtwBzJoNbyZHoeXb6oaEsN/TetrT/pV1SEO8GPH3FmC
iVo1yQc0Ln0yel8sawvxt0xRf2jTbRWUjsasC7WyWbYgJeMHBZpt7IMxX9LUBgCN
EILUiact8IGFBdUaHQzyfzkP3ZF7ZWSz+ZllI3yiHXIkqTRFh4F5hxYH2HGdTspx
YS+WaHd+JaJnwWVcx/N8XmYp0xlZm1vLaoWEcVgU6IMHkNx+IY5CihiHcFzWmYca
dK2cOWzvril1qxQXzZyigM7BSXJ+ZGfZS6cq9I/5E5sU0iTd44cSEPA0riiIXZ1a
F7v0HnYK3QLK1RwBy9fUDnqR3cDZi6fC9S7lk2bFsNEb1R5W3d9nLdQS5mZrZsMh
p8Gqy/MCL0OBLmIy3U2VZi29dsm53HeuI8W2xXay653j/DjphbzRUdy8CfwVvL1f
d78/PwIPuoot60YRJUJaq4rpg++s2tKfGP66mRmtacJGsvpeEKvSO9x8aD+DdzxM
TUsFeZMwtloOGeoHU6L+jtMLGcZMhDQYWZudg+NTaZrBnQLY7/Y4wd3ZMN3qXziv
6QSlE8BVJPNeJPeQ6VRFvwKcPpGTHT4ObVmjlFF1ItGE84Tlq6KaBNoTnHkQXBav
19zfOlomiKz+hO7dgrpu518/McWdaCe/CXHQzfuMFV29Dx40zOlmVbpX2LKUYqmS
cu5E8JyEfXVI1xqHzWQUr1fX05IISdflVWc/HD1UTpbZC7ks6TEO6O8mtVZHl8AW
Wml/JNIaihYzxPD0bJVen4KQn+pb0AbCyOp5CyfXykcVPpTjq3a5zP17g5Ntd6VK
uVcvGF5zeOVAoLvbOH6PUc7htHnFQrWZ1DhrN1dCEFOZloNy5eEJhDyPZcQHMKxs
TqEZDEJEAwcGDcEuP8xhGdJ56n+xWSoW9QFBBaQma0o9PJkWsSt2tiK/hsNmNX4W
fNHIV6+uqmGC3gyBz9ctt+IbqucVH+vVpB5qBWG/Ci67tKv3NxbsuCRRBp169b06
Vbg+aCwRaGzAJ9zoXFSWWFr2T0H4O2fqFOMH03AYoN3kP3bhI2JHAmZyVjqDWBqd
heC5KTwfUivgTtlL+5eiEMASZuWEd6u2ubnwxAjIDd9OnlfA3z6QNVqxiSbJkYR2
CdgEyT0AAM8iSTfEfS4UrAyHvE7sfE6jTn5smSkqdxkxRGvy0SCr+nwbZbGSEYbe
myU1Cyf0mNr0G+DhAnyVao2OFAfEm+pRy8dJQNjzEVPNBSaHJQ6+nrPxJxaUd3Hx
Ogi7EtC9XVCpT+eV7XTevM6p7/VQ1PPp8lk8VBf7KtxdfCcSBHaMPeBQ7xGH01gy
KCNe0WJnrFwcFAutbor3ybPQLiks5pufjbLWDHPb70zVnS40rhU0oH47JPSo8GrM
9rv92BI6TrB1ph+u+AZO653+GbkRCm7AOqfTxcdzB3wMQkdUHcicF1iNYi3oh0aC
RBgGMPlKjvNiIWvz1MMQaOikRgP1hL4JrnSuuJ0D4GBAasBfMlHXdfDx0Sx70w8/
mm3kgsmELH/KcRj77z9vane3YXv8o+igHLcDpcsgqimzJJ/tDHs4tQ+F2LYOkbqq
luG137O5cdOyZU0tGYferQX9ULlBD7forVDlJWWr6ipR0p0QKVAZM7f5ZgWdAUX3
0ypnwuAtLLlTq67hTkJsI4meoKQZMe7Lk2Syj1qL020DcOYxxXhK/Zfv/WFz0LaI
eLLjfQ/qnhhkQo6Y+6mVZI5l3kXjpa6+9+dr0jLT4VkctJ/Q6lqEUxQ90hckDbUK
1j4gFq+Pps8MXqoZUt2GQKgcfhIfZdRNuEjiC7DmsVdihKqKh1YZNU8DixzvIVin
8jdyY5u20ETSbqsTK0AT+CZXWCrC9xy0YdvIllm6mBzI0pmBxl8UqzeJSzx5El/z
v3NCUu03ss451+DhWsy2+XK66cAspGBlunqsc+YflStnPIiwVvoKR9MUioxogJS7
8SGcFNWho8U767x5vSeVM5U5L+lq6M6IuMYPUFyWMCjGJ2+J9tgtg1F3CeIE0BOW
YOKz8ghA4NddJdaoeNHANfxKBxUovXYM3LakShUkFRfYge65q55DiJICQPyPwtBl
KKWxswwt2kUeWTzMWTDF2idhQENzlGjdFHa0uU5fcfPf2xvOORwp5Co9elcDTcOq
xThg0xEhtmGoSvmSbksDtdbhBjCKKvK92sNYIpyItXxXhahSDu3ZcStnXDw3U70M
UGEhw3hJuJjmJCAQ/iZ+gbS8UkmZd+tzqaBMl9cjT2BhaTmEfBWEny9yiIyW4Fje
xxaUjG38ocJ8YDPLjpjVj9plN3Iy8z89t4PBQyo1So/CgitazXKtsgOUqGw1n40Z
FQaMKUAJXipbUCsanNHpONgMuOYQZmS4G4adrPkHDAASWjKwezqn7wMq3z+QWd48
XsrDYgUiTSNvSK+q8HQV0p5FqZhm1CJ1Ehmqv3vgQFNSJl8lx6QjpsNF4wSHtJxb
/QrAaoJwH11l81GWf32muHx/4SekeNYuUVG1RzEtDSNEL5/TgNCWuLN8ArOzUAKT
4PABHbi86xc7/RojbQkHcb7ik6YqelzuH8MdHx/MtDgCr3BpFD8y5HWZARTyM7i/
qHHmygcjSlnj5aveDLTmhoubKrN7Ts8mQCKy10ftc/wFgwCxu1evmhmXgQpYtP9Y
cgmHPLOvImUWkYcHvmJLO/oWnoj5Od9i8LD87IwbM61xJWf3mfu0dcXM8uH00w3V
2Cpi+jdhjO8qHN9rlANkedbydY41ToUbg9qrls+lYKlSKf5pFMLQrQJSQhNPt0Gz
lb26HrTPbOLmg23PD5TsG3P8L2bPwf6jSn4jDsMyTIJUBjEClC6c792H9jFwOV72
xiiAu9IFscEnP767LhjHGLiZPIrJF6D3URscNyNao2u5lSk5FfkhSPtw7LEzuJua
zTJ5TZIUGN1E1o5v+PfUMx4owldOnhb/GoI303BiZRozhCJxdEnu2aDm5ymkm4e9
YdlzsRm9Js83nq2kOSe5qTn1CWjKDmb5J8DIA/VmnnaVvAnuATcu+KPw3+TCYBX/
3O7gRMDDlNhBLQprxQUMly+GG7h2VOe06DvnKVQdZu1kgEn8gKmNrT8BM1bquurP
849csM6EdCztJTTZ/5dfUXlazjsjGYRkNvJ7WdJay6XhrRJ6P2yLWrL/Ro9LugAJ
mumz7C0Vk/H3Bf6+ml0tfGbzW4vEGbKuaJoxsBWxNq1cDDtWNkB2EtV3Hb/ix505
WvzHDT84KWv5roCeimGpUXXTBW6HzRYS1bMPBqK0EOc9B22k+94FsIzQabpE0ddj
UKYPTVN3y8Cm9yrVCpZi5X56XMypjY8xOLy9AmcoI9uWr3ybNNeuC1saHkJ2Iy2N
uaVfAoy6g5uY5Ao2Xmb+jzJkbzpgJfrKCJOss0NZLCbDzImHNQf5jlxAa1xDIbcM
D0jgDOUkqfgq8slsUFLp7ZXZ29sgxItcqoXij5vyKQk9fvwiMjpwMUTNSd7RauWR
Fxqae04Iq6n8+Fap1HhGdyXFimK01oe7+kE2CuB6RZBtA1Aw7hwHhRPGggyOECXb
PtehnjFvxDdzgBamYDoGyxFiCbv6AwcmeIzh6Qe7TwD8k8T2rhwMPiktoExUK96u
od0qUXAjV23GDrkoDu8u5V/bSNCjRO3P9C2szAT1QDMS4E9ZXehKfPwiHAT3nvSS
sRO+6H5SGrSpmzSMw/gVxIQ8DfweKBSWuos6yGCbh1mtsvLjKTX8NxUY3hjeU/f8
nVRxLuI8frGFLbyKUtLZYrSaonElmRNJigWf50mb4e2MH4CebKDWcoB6nNc1EcNP
PbUAR/Rr7BU9Nn7kNZdMzsfRBBVwwwFf8gHVCXPM1KWXmQhKtp8HE+tB+Z7K3dtu
sepN6SO88Q2IVKUPIUiI8ZcRNnqw3IRjkXm1hvA0dm8Yk1BectWg7h3oPQj4Vxh4
oBKns4eYs6wzOc1oZAqhj38vn9jK1XsnuH2GubGTDtm3lc2sNgc/BoWv91YhX7Hv
Y9YnignvtBO+pYIxi4ghmsMpdjbFnwCO0O43U1Vb9CmK5cPQOvAyXv4XdBFP4gSN
qbikOa0XNuVp0dxlXQ23WEEyeas62rYxxu/smZ5WHIIhoXPZUtzTxbT7dqkrQ++/
MVm9QJ6BRDAnXiUQVR1DebdhTavgOc6K63lW81AQbcPNEuypVUyJcIrba2z1EB2w
a3WoPfEi/kkU3Hd+/ZUZ1rI6s8ZKs4XfcrT92Zxm5eOe3mIwbnFmxVwEfW80w8W5
AKVUKSGBwzfLJ7jq5J3zWC6dZqlHRpoSlC6eFrpXfU3r0CY6Mk6Y40vpVHoVTRXZ
phgXgyELoc5YMx0+vSRU6/1qr2aiykd0mmr9uvxF2EOXTi60k9mtdcmCaIg8E/sI
9sS/7hW05HaSnWeYTSHtZzpDfgnoRxBQSpoiaovSW1P70TE+i3gJ8K8DoTnxmN72
8zl41YBYFgxgH41ABU8N9meIez2tq1nEb9l+lZNTAmXm91NiLJlwNBc4QKssU/hW
qgEyRnSW8BFbyF5VBFfn+CF5qOpvodrksT0KHc5kLbEQH+pTGJaJKwt3FHccU14w
8Tn/ZNXQdvK+8JHQcGjteIEv3JpG3jJ3KvRHaU7Z+owA8enwJBdF9C4RPtM9CzY7
oe6CxPJyvu+c7m//hu5Cr81ocbPNWtWg/H5q4MhgQ0vNpTYtWET/7mkhI3FDw7qF
+nEEoEqo7uNj2SLhAvlw1XTdUWoPKyGW5MuqiGS2LbNV7jvxlnOIDqoreOVfwzTX
ahkbFcZeq6X7awCp1hRbvs/lXQ960n8Htj40LV5Yi13F/eZyN/iJtrxpNHHLXqOX
NY84uadc2ckTkzzTIztStS+LKJC36nwkKRKdm54tGf4KnuulPJQnNL9xpX7R57WG
Z8CgD+nFs3TlDQvtM/N2ZKeCD95SqH2Y83XapTXiLEuJWrAya9OZ0VLLHDhievnH
cRcpYIWEwZjh0D6yLGrJjOFwkQ4akzYD0hzdcpWd+mPD50kl7//nzowXvfwpTLng
aGk4h2F5hH6GoJ3qgKgxoeLHoZG3KpUgKQoYD1haGsoTMwIi/WGFCtiGA8LqlZAP
TEmjk9ZB8nyMwtz/Yz/Eau/jXx8H7xTBCCIXLjAJLXdb0pc3+Kz057FQoSCpJF5Y
Ubust6FUVcLOTmbObvNfDOqox7o5OVZ3v05gwGwijmolafSnfdVC4zRgXVX3o/wq
OfQLtimKuh6+cmSHlO8aOSG6ToipKCzAT3JcOyQIEr0T/r/deMn322Q9YtPQ0DiJ
N9/RPTNidwXExjY29PmxMJz3bGC8e0jUondcHFmny54SrbBFFSC4ssDeDp6g8LcF
kMSvythwiWJj/L+y2ZdlUixE7DfgJxIdyFgD+2Ef/5Fo6lm7/4MuIQxZKixGOBzI
KY88OUs4Nhh6lt/X1sUr9gj4Dm2UkCLei94QLE2xIsSO4mL5XozvSsfhncvcyCgs
rjJUeA0uS0nqggLnSd01Vj4h3XhrpBVgHqhmGrtI3638eKnlk7dbbAaNj4zKDFu3
WGy/ON20aZ+msGYtdkOe6HteOBXimy0SogPTX2y3iverlwJWfgOf9yPO7FPk7piF
/yJu0lEol10+WsnGXnnfMTxhH7kod4pF9rsLnySeVYdE1gpuYFbU6q0dw9KRv18H
8ZoOcv1TYWA/rEYb3Ucuki9NvIomMhURCTAIqcp0nkFFhOv4AU4ig21HdhUaCcMm
xT/2m8sQJ5lPZzR3ZAYfHxRNSQa4Q5TsszF52JK8QrvRii6t/SX9ZdGbMr/vqCTF
oVJkAT57ZXvLMvMWfmZXXfDqzdaGkB5plV+peIJOeyIfG5ThnvVsmLxsnNR0Zt60
p+tKC04nZhkTkRhnxPxvDoWswdNn1IgXQBpJOLhiCje5HybyeqOCe8A6l024W2dy
1+spPVm0c5ktBwQ9jrWgDwwAmr6hNszDmE4mK/e63jRbjl45E2qiewNHv5Mt6SUR
EPN+GvYuAKQkjCGuXr++gpaqvy41w/+hT+ZXStVgomfFN+LXNtw0PQQsB6KazWzo
zzUjlmFgzPJuJ6wZMo9OQk0Mwomgl8wBgjCmvCY37rCXsAbekQe4KWbvjcN9CpfI
LAC3+XjKyiI8NOOrDeEdIMLZdhk5y7D+exUn0PENE2JPIvJwypn585hOL7+jBr2j
tRK2QFMnbnCWl5hRtcta/eAYhj55yBH498T8YANe+jv5lWhU+Bc3JZeHrqoH8CT5
9/yWnauSTzsdPg+9pjegDt3lBulxE+Febh6XlZzFhvlZscpv07MtHt3UuLYLaaPI
CRKV/jiehGUkuoQepckUBXC/zdaxUcTYPuWjnnB1UoyOv4AI2xU/9xtlnCZkFp2l
VoxXcOuSBhTJZOR3Zfcyq1rt9nqjGp+KR6J9nUr85xnYhk4HOP72emUr9+oKksX8
iV1a3LWgL13TRmryCYY/c45MyxBwUG/rh3QFKLOGvjMGLqLdPwgCcMGaNQYuUz2R
VjYEYxnLwx/RU+h3Ei7S/KKtqlE3yO98S6Ecua2vc/PeKVxAx/Nm6fQr0lTDce4d
FkmzRPQRHwpxn9VmGKasavWzh4NgcoU5JTRxF1mfcBgdPYMavh3hg7wEEXKpO/8/
px37cAufvVbqk//1X4VAQmtDGoeVmweAJLf3fA+0BVyhrHXyEWkKyhisBIbOsEhk
2NiSUJDt87pwxbffaMLNzOaxsXCVGLZM44ytaEyUih6/wxMg/03GLXK2pnQV9e3U
OM7TJcHGfj69/sJ0h/Qu3vVkj7K7Vp7bODlDVqqsKmLuX4J00AtdSpDEAL5OQm0I
Lfg7Uq7Alj+R0ThdH90Dnrs4ef8pXxC8zK9jNUWHL56uXjd6GHO/kUzpL6R9Rbcy
6SYDyox4OHCAJ5WvebuiwZ0zqpGi/iBrP8BT3ICd88z2mtGW4jz7bX0NfxO31kdE
bXzD1Qc1S/ML/EKd1Y6dVssMMZHuFr/O9vt0Ke/KEaB+Ff6IcSu3jg4wGW4FYRBt
Bkr8D8hpY+cjczXkZLY5e7zGSZRxvO9xZP7bpnTD1hiX5PsWVafdEZgUMg6ztlmx
cdzDmdO4ArcW4oFLEMUW7m8JFhtVnYOoNjgDIuERKs9EesfvpJjWrMxNLtbe79ex
awP0g0X4RHm2MKa7pYSHuMX1LN3xAj373B/1VjCE9TpYSg7VkVP1RX+5/IOo4RtY
vOCUz3HRq1IDOwfyaOVVqzYW1zqfY/eqr2tSAtdBzEED+nTXEjnwNWSUoCtjqvrB
PnRJ/7RsRPFWoWBniZQyLxPkrCQIwhp8bqi6l4u47k6HzzgmYUZZ1bs2u8vsJOiv
rFpkI1qH0gf8q2RRwvNiXZy9HivSvkRKtq9kEsFqqB7vu5MpoL1r3L6S5NF48KP2
I8bC+mrPV2EI2iY8butPQ4WCuyMKWig6iTe1vGrJaJqqKIsDxum0g3yJHXHsb1UX
Pgly1w4yKuxsVWU9mqhecSsM++0d1SJ+CKaMY5EFUTO1xCXxug1TA0HdeIrhDIlE
/c84LD7NTsXsKR1c5uB0SzexU4z6AbdY9gQH67lv/n3Q4VCA+E8JE0iInOkXjIa4
FL8eXuszIpbeHHR0VWPI2p7yfhIwY5BTYm8IC3Y2ZBPipYOC9psnae9A8i2yBPTa
gK71M9/PN9LBnpO84KygrGlGgkeI3AG9xfMpj6BtXV/F4QZQxrOMQULa3Or2y6iA
Lbio0JX2Vs+2h8BwC0Z+vjuz4R+tf2wp3MuAI3fEqvauKHhda8+6Az9BTwVf8EMz
4Pt4Hva03VHZTOWjrDf65Nl2P8iTNgAdTKgGvlw2hfOlMg090oSDOx+6wpAUzaUu
5jo66LMzwyKrQyN0WspWQ1rx+89ZyMwf1ZzqJU1qAu/suOxwUs1uOYvfRAx7dNOq
RlDkPuBUqOijMS1veZG3dZmGyo4yWJR1bTHU3P/gMuH4pEZtWluuWf/7rirzDGr1
eaTZ7NrMNPkLxsoVlcEmw25PvPHzebPzCSTloU/MRh1Cx6FEoBQp7QZPv8oKrIDq
QC3e0tuRTHHNW82hLvsqM5UmjwjpFQLsvXzbUjYO7nAytQr5aztmROFiKenOA+1R
fsw1iZNkxUwLsdkHkRLNVxn9+04cbrxLdkTtcsrR57xLopH/Ipqn3qQwuhGmxp9+
nEkC7ZViIFafWjp2sXcYlhXQuE9cj0DSR679rqg9Vh4J6PRc/3bihR4s65Dg9COp
eKlF7G1tKaNWbNhQrLoik6XqPHtYQVRv+5418FQqbLH0qz1jRIlcv/0lxZ/CWq0N
K0UA9bDUxHk+mFiwq4QcyKg3hnXnfg4UzabDQaK04pXgxzfeGCmOPzaDGx8uobZ6
fUR7eV+aeAAKubuyipPHx/n0MvqgwSDFCiZaiTotkgdn8Z2HKB1lnfWfkLy6NVU3
k0gY3GCuVf9beXYUkw86oMxbsB+aI6l5yZFgEiMsAXBopMY4RHvuiDWX20FkOxjZ
MDdeafpoQKryykVXm2VujQpbFIc+hL260tH0FvTGoYlwp8OpcagBMD1vLe0cMpZi
Ke7A3lvfXvxZ5zqXXDKad0G8dEdHWiiFEawKsYVUe1560Y8JcppLO53tocdekfW9
CGtQw63DsTLE5FYMg7z7vKw30p1yHCeSMIwNvj22nlUSwoxG1uyZXVRdqc4Nh783
aFakKCkgQ4HE0w6ek2Ht8ZmkLgdtnHGu6y2O+CpWfN0xWZMEodWozwVMtbniCbYU
PuhYiUo1Q3dbmIcFhnwwSxowlRV+67jYmN+26N5xRymhRzYsaokCKjSnLG37j3vM
cgy5CW/9OfZCNvi4lui6XDQP7EqmpW3Hbj4KEVSeUeS0yHK7p5MR7bwZ3kUtwU5u
9gmz7/aWbOXVjVpgBF8JtPkTNRt9S20QKZ2NqgTknVqbh8Wisw69bn8oGy5bN59U
xauTNKoM8ZwvcMstyYdKVPW+G7c0hjxl84P7fNm3DZFjnenoL9yS7MFleGESzjoH
d1Kh5bRYyOq7Cj7rKnNZFDUbxExU09r/fciuGanDtgfUMC6WpDjmT6Zw3GPbkuBY
1QN98QU2ynoH9I6ULGfltoYzG3A1UVMJ1RIX7WRbt4kVMroyGRFGtkh9979QCXf2
EXxLaXMdlb3MGGttfM7ogRc08rMGkS77gVyB46ZB30QcEUESwmllPk/SxbewYBxH
l7rKWI3dj5AIU/J+ctjCMvM+aWI1mBLiNRYKrnBKg7RV0wN9UG2YLncMS6Zh6qkl
xyyH5VEv4g4iMD0s7XsNhIYKepaVxouVOHUcn9P7udjBVvDq7SrZVw/LF9D93cTQ
lSdukR/CfdXhhEUqfauT1aSSPsupXZ6/5k7/7VgqM71o++U7DDiuKFlbvq97ZkuA
6hjcK1T0i831iR+EpubPY2cKoAZuyg1d5MHWr6nepvvw6S4KAjfrYQjON3fnXjYd
vP66n0VKWWs3OlUi0+creFX0bEMShR8BU+SWrRGZhZqmKG2lTg7ltDkRyMZuXIyR
gElj9xav9SGwZ05AHo5g3rPB2bMubZf3CI5YGcFVzkdhoLHYizLjNRiG9S2eIAtX
ELU1QVeBOlwafcNYoeoDhczTxqf4/U6t9D5qoE9VfVvWddwsW9TOFMOZkglEosp4
UwUsRRnPcBo/xPDg07s0k+e6BX2u1iOA452Cb9QHlKRlMQeRkVFdXUYV5HMH3VeW
mppWfIvlFKAqq4grS8iq4WedkZlFbdhe/L+3hJ46+9m8w42y/GPOXvB20RKNqcpR
jT7TSDp6ERAxm464xrUVAIn40Z81rEHbfTt4eTCyLqMWaIDOtB1CPx0Mw9Mq47IW
ZfvfLm2AX0u+RqvdiO0GJHbaHD4FNhacyFsl+C3V6UQF5tzK1k5LemHOvocQzWXn
4Ew3nEm9RmMwKGZIZ4j2ZtC6KZY3vrHqZ1Sj4C6821jPicn8WUUO/zdQtgLYSVn4
QVdxQC8QQf/An60165dK1ariHhyXCRTmUqWD9+uTNSRIZpoB7kArCiCrQ/PUYY4E
LgvfMar17pmvbRiH6IouPPAC5WIQoerkR6TVXpqPrBoycr36Nll5Eym/4PYHjK1u
RbszLKu7sGCvYJwPA+5k28yDYklyIFwVxlQO+lOThBABF2ve57FtxzaRwHgizWmd
T8QDHGimZfHp9N2S7xYLNCnev7b/3K092AuUs3My1lL2514pe7OrF4YJeHtvo9pL
vl3trTk2a7S0BIyLpVQaPluBKgMoxfIXCkesqj/F0frFMt9IinE0L5ga6XQNvamO
J07POJD9+GNHWcEkZrsDHO2cK6jBMqBkif57Dcg3BWg93OEwo/ylrw5nBa0Zw24L
/7TFhZW9n4DmTsCOX5WrGoDK23mmJIgbrAOAep1O6g32Yo4ccLndUXhA1tRAwUYv
/Bmv6C3slpYMj8WZbAOeFDJWAxddiVjT0XlkIwYH40ON+J4HADY2zRzMm2tyx6yA
VC//VxbfRr9c7ZPWjUuvZyyqeN6ZDxD4s7eaCl4k9I1RoT2BDQmy8gkALNh/uwJ1
HvEYnxiqpTKRGOw1ex9A60PEKuMDfPHfIgjV9KWVD1qw7Ynj7Aip7WwFzelcVYLc
ycCe1yWNe84TP7PwHfp5oBp4mSxuI5dC7ZuEwr1hWmnTdbun1W8xnB49o6F46iIA
AE9GxLUgu0BFr0leC23FYOBjewys4HPLEn5VbHSBzx/d+JJmM6iQdI+FqdiXQzjc
Xh3gEeQ15LM/pSTo5kZtMDQ+agPBG08mm2Sl5eAora3mHIUc+jxbt96nEA97yYSA
kbfuF624D0X1r+tgLrPcRFvrZvACAjHxbFTbMft/loZKkAESOmjCnWz/os4xXMB6
l0vV1hkJwfa3G2st+yg/Fmvt4lE2bwPRw8EJfxK36wvtSvKxet34TXmfc3wFx9e0
ekEINqL1L7lOLO5MFgkH3KbEyNkrzk1oN27QU4Yq5W+IUdueyP78KTRpjCNfat/s
fvDivd5iWiScWL3VQ91zTVDpyOv6OtZdRNqDhlTsEgMbVJpUrk5Pv5w3xPchevVH
32ou35jdF3UHEN9BJSSOW2+hUpYX7mCbli/z4Qw5gQs/d9X7y5mletPMG7dSEZHW
x5lhok6gE+y5IPApDuIvY4rwFl7LP9x2iUzQruy2dG5F3ZiTeJcznU/9EoAkYLow
81b19lO293JMdQbUn7xjPf9MTB/Rl1CExv/ggTEfWvdDzsxYuXH6GZG6ZGvQvTq3
jdnBYn6+8ynRj5LtK3H9Z/ctWLmD9mTneSp28sTd4eiJgXs1otq1oRPExi9C9CRj
KojxcubOZIWa6rWxefRk88yyf41yZw4Pay0U+swo8+5k9jBirBPR0fVjNkJgki5B
U7iWNmjQqexzDUUF+Xln0zyMq+NjwcDWRWkfdOfFAQsGZzPwOMaWHDO1+bN8TMbQ
G5IXgZ0uI1sC+vml4A3hu9V/hqrm+l9nvfCo2Rr8SKeAWI9jWGotF1ikucuy4zBf
o9x7RqfXon6tCYCVBqgfDcxpC2gr6w/2Bb59PkwsctDHh/v+vM9p5Q431+WsmqZG
QGnFByHlxVNxyTg3CgS5qPjBMPQoepNInQs+vgVbC13ilSypT1XM9exVkHB+H2i2
9ziKTBfWiCUp+cL9yTvEz3TOI5ocCabR0OZr3ElwHOSsIcI/aLKlaxDqS+TUmgHd
JTO3ZiyAOJCrG9t4fVts1Dwg5YQ0FPZ4BhoVdQwMly2Xej+LrrwGcX76vOphvPs3
yVIOBXr25/ytQOq7qeljQZ7GjUJ8dUrW8PJcxzUeY6vylK/RjWhTdm3Y2zklkm+t
26QKrvzE56ip3CY1sMvePiKbGHXD4wgBSojZelqourLhdDvglzuQUI34ZslK3Kek
goBEpsky27QsLB7JjPnR7gDHeh28tQKHaew9T9wYvp84MJALi8GjrGokH5GUeD9s
XLEp/xn6nTj/fwFc2S8t9imy3PmDV7h+HkhrhtmnyYIwHT9i0QPVZHXWK7pbiMbG
4B06uO4ztT/G5Npyjk0vVLEphKTVr8O1ZCAs4G0dWzKm1dX6WpieBA8TJwg+KyhY
hs3S7neiZBMlBWwSD3Owo6LD1UmOM30vYGLw0pzC0ovvqWMVO++571RBJRJiQu4b
n0HcFjyiMicqmI/iNDWsNW484d8/MJeIFamK2NlTBMhWj53SaPdKOATqhYrU93Vl
k5xjMSZ7LZyuEZGtbtJncxTfqAhdsqGZEZwp5J3C71HxRp7ZJXkErVuD9YjI1RMD
c0bwnX9UDYfNHd8aud+Xe1qu9qxl7pE/Y4Y/0Kgnkz5pTC1rXcGn0S/nHb5B6oV+
57NoPH69dgrAGV1n8CdcpttrLRSE5BMNnmqsq07VNZ3ZkeqW0slvgul3KcZdyVyA
wD14le8eu8/aoiITpaBGkoTTdKOAHDjju2gV7du8FHFQDOUPiPpmXnJhFzXMUHej
WDn8kg4wPWSGBVNPzW7DWiigJmyHdV9V3C9kjidAq5v4K1MJXqN1VPr1Dlw0F525
URDgpA/GqAt5dq28ySCp5nZnWG8RXBzpOPGxZkvNNcmC4j76a3Ixm8z2AMTUMcbl
v52Atc6+oJHsXVpTZbrMSb1oNj0BmLuoZrgDQCInH0etEhTmaO+urf1IWEWGEiMk
WONa7yRAlraMcAEQlx9oFfoT6x8iQ5GUg9HV19L8JZPmDqtJ7aaTSa3EjlUrKCX6
xDtl0DmJ0K+2Z5VrlXcWeOVuNyzS1LDzjAgTGZencjaLf9DIlhszr4xq0mWpOIxJ
ZZ4VVYclcYQBQypc86W2mHuj4e7LQRhduGCRJHa3JusW4DSKy8Stp1st0TTaE0pn
BaQATbMGTyk6D7zr/V31Uwh4kCqwmfCB77WiuBXNh8WjMbpOSKsLrJDyKIX8+OxC
85yvnsWl6QrzHHruYTb7gPHwRMOTmWjM/gAw7AF9sNzhqYz6xvGfbcXs5bfj9gh2
mZ8iDfsBQSr+5blFpemAn6Mg4mV2x+08M+ATneuzCDMQuYQO32YbEmwk5X8mHhUb
4ua4adlXfLXarZkkiiP7O8di/i24PKmZRrEnwn/el/8QjQ9131/1AnJpLMdB3cxv
8HwtxOBOwCm95eYOFZKHNFGtdgJpvIxZ9W1MP9DklwfCOLMQbQW7nXfrCnFl2xte
avNy+WlN0kheMhTCFJ+4tHoAkjaTD5h/R0Qmr03RpruYiuN95TpFl3YuQvNjSzCB
LuT7r6uWcX21lC0t9X4oa7rL3bIhtOZQzzGVlfi1LqOeUWliJl1LVTyUZZn9RA5I
Q7i8qneDR6ynwoPfrUaWU+d5E3YSPU+oBpMx6zB4g3dHzWD2Cbq9s/SzdIGmi3o+
pPah99zUxpQv++HkuHtzsdYbf/VlXqSmfnhJxFqRxeVPuC8j7Eb2SL5pS5bUiSBS
wNqFwpf1+0Fag73apXZUDmErDBvEPpPQy3eny8Nfa1kHOflEsu7mRZ7ExB83bM/k
IdNatS2Zh2oen4uZy/tQsqU9UibdLFIm1wz7LdoDFnEwYzCMqeGER1KWoXODRDNv
cxAiyzc8aOWNkkJfyL0X7yrKUT0HsMpLMpBQIkDuAWFROBFJ8rbRaq3QcKneb6c9
p0SzMKuW4QhkbjL/WKbPG/2znz2Wm5R9fE8O1qWKIZgIwF56uc7IbpjSbP/vAHPx
6lMvuS+B7OeCJN7dmw50MnYSB1i34xc8E9l1rF+F8MtOee/eRlL79X/LuKKo8pIp
qdW2WPi7JuQDl/ZCUqB6DtfFGqvDK3Wdrw4Q9FAqhygYVWS/7LPDLZ6uyVcbQOZR
8RI0kEKdLmuVUMs1S9bKfrxLf6aV3Rarb0R84a0rcaa34VJdgKC+xvEBi0hgKEhR
4oTw8GqQDYtw75a+Iq/1KQHSqI8zfOIcQKhrDcLSOvj0JZRtgnhDu3etcDf9H67p
WaRkeTHDZqsp+5EeQ7Rv2nKNhzmGayF48gaTWAtB69rwbHVDiAA+zF8SRvHv1MRI
+B2nT+V71sWfl6g5sB53L+/5B9PlvSiXtM6G7uIJuB+PCGZhjyg+4OAfDmdf394+
D+XuPrQhItBseYpC3uWePeWojjcXA6Lb8I/G+8quHWZ21OFHAV8dWsap79IMsDGC
ZjnYrJ23TqURizMaa5ZDNllusdDbeGkMUqlWiHJWTmw8g6g/+ME/7LggNVPgQV2K
NNqRb8IDtnigP0abhMXZtPJtW7wvD3MNWOC1vUHavWI9gS05MP6GWpBovDu8UBhK
1FgzKcoTM+7gIPeDf7Kphp+6UuKH7PV9oq8oPXd3m95aX/gdXoG3ZECQJEKZggSU
tNai5/WU3udswdUTHY3co+BkeryAcxTi6zhisgQ80BU2dzrHT95Frq8jseZtQNb2
hmowyZlYTYTBwyWIORZ2L217N+ekaFRMTjJDDt5h/a1NgA21STqhlNQfqXjF5ErI
jikDfHcWRinuCKD8LWsdA578v6jegSGBl2NwqeD/Czegtww/WFixF9JC+lwnEOf6
GixtY1cqjO2ZFsXutKfLao55Jc9K3tejNuCZNn8GHEk4EaDPGA4VwtM/0/JOXU2m
xLXAmdeU9Dy99f5sFTt2xmjYj760A4ntjRUjpjP3pnxamaavtaRV/0NmBwvln/Vl
Jhxo3P4ePGaH7rxxx3GZhnP+yQ8Hqd4XJE2cZ4JzT1nhjl9saK9JBzMWbidyNB59
kPLEx1uIRafuqbyOVyd3mHfMGalve5+xRcJo7gTYlQ4ITMr8FkZ2nze0/a8fICgR
91yLWqcZGiwARYXP4ldu49DFpDcE4RKwvzQs+3e1rwo2TOzenc03lHl3vZNOMHn8
NijgHjmyHjW33WmZs0qwsBXmHUJBb2S1/0C0px7ITxaO5hCLXQsLpqvGWmdRp6Hc
K7rXIyeQE+kfLN59zgIt3GYKgAC0m8lM5AUO22xWRMjnn6PRMTnFQBlRtCexd5+s
3vtpZ8ExPGGM9vNKyZ0GBaqbWqAbpW2LrlWXfK3cESmGCRbBi2IaippUiWTN9b67
M7rrfxrOki5kPei3TCTUhgYK4+vyrUJ1JeJd0B1JDoY5AA42yB4sErJAIl8gbD5W
GIm/97qujHtUhu0kymqPLpf7H2so+rzt8HCx8Sxb4rK9KZKmVn5H+pprYglXe7NX
P2BTswKdTercI9Ijb7bK/aM8TzN1znpggE8uyeo6n4LzShmK19ugpszpx0XKmfCv
/kHMGaUtOxC7w56s60aUkjzxSz5/4LLynyWmWYJK0JcleZEFn2PGvnoo0UR6uFc5
bcgG1be19+p0XzKSF5JPli7Pnj8q6Z+tn8u92iMJ5nnGGcc238W6cB0YW/idKZ6x
Cgg7Glsz8/sK7F1nAWlREFyO6FDIOLVYzZrevzWpcMIExPP74ib3sHn+5h+Rk9+O
0FhoqRYKTO1VRHqHLQvUX9QfBGzi/I3Eauv7lgmR5KK3uEeQD2zQBGsYRH0Q3M//
l5VAk/HA2iCsDOnbH/0tI0idQDAgnnbCnc1fM3RDZWQUx+RxuS2rl60Ee1sxnYb2
ixPTP7FSvseJ0QJL/UMP5QPHMZoGdFfEBeQdXBglSkgxS8t+MuqfCsQzOXkMCShN
+3T5p/lpcbrZmrBPv8dQsNthX8XDJsj8M4Rw289qYUqwpUEQjfbJnRsytpdTHsM9
J/y3z0fC0LHb7W9aiWDbHMt9FbXTd9p9s0cr5yomPDwU0WRjLh98RzDkd+KM+li3
fsaL7VIKEYmydf6FfngUyAnZtn51yHwUryveOao49YSkmrOBULs+IIxlLoR1Eiu4
oSJI8R0JP1or+aB2pNyQi6wrop9Stb0JwcNmCVwhhtdsgslM1Vvn1j/rL4wkkjBD
5klYiu9ojT7n80p09s7uu5is38VxmjYgFTOXZfU4xtyw+XudPGFDfMP0SbiAwAE1
gtOpyWTEMHdvM9oe4ZRPv5MjRLjohuYPQldYBF3lRKL20EBaxqyPeDhxgP9xZAje
Sg9SbCPdDFdkQdyzi/PEIeENimSZY8S9Z2rNmle6WntArGFvlA/vTtx+Ne2GZE4j
ZdkJzV30zcwXKc6gNaNAu9Wc4pGpO8d3RFYtTAYqpz5tfDzFFcdm6SybvQOTr5Ys
a5EUJOIC1jy3D8rYnmOOutVrP0DKOTrbajOE6WQltd/zH4yhKxGN4U4Qzjefm4Qw
l7izYOf1SGOLEC1dI+46+8NXe9pPCOlocOGBJET3zcXlJ8NRoqIF89zI4CIalp7b
ENghKjwCxYMcRpmkVAC6ykxra+YTWQnpByR4JoicwxOPC7RTaCZjPXT9+oJf+Xyw
e0QLyMUBKj4qwnRYHZiSFsjr6WpdzGVBlcAx6+sAFj2n9BOY1rebwUGrRYIyvkbs
IoRX9GJfBLD+C0RCloY4XcrNI2GT1M1L+o/IMO8Wmq2ARhaelLinLTuM+9leZTrF
6pWWmhE9785dnlVJV5jk4ft0GoTs0U0Tz3nG8iT9vbeJTtCbvlDyAVSf3zKppnj0
Je7CVE4pq+yczWT4j6DxEXkb/XnAaJ48ubM5RWPs/8em+Brs6T/DwVJz3riSQqJW
/Ys6N/FBLKPXfnbcAFMuZ8UwhMDT6oZCihPxy95DpIPGjy6BtJktvsDy1utXsotG
drh3khXIKeKGqN3lb+0WZ2ZM9o7bdspyt+zjedFnNXE4nZwX/TKNG3Dowi6UVWEV
ikIejnChkk9NNEQXWntQsX7CPBsTB8KYy00M8mWfzwZ6jcvBfmreayBxS/wYrmRv
ljOUBQnS5Q71u++NkF3RLhOvJLgE4MhNEede+OJHfFnelmpjd4Le/1KysHXuh2i1
ampaYtgwJyV8vt4YeeeZoAXsh213CHyJSXEjs7FAVUlEbUvMBdzYa3NCv0tCigIV
9lE1O4mksyWvEO37PR5tWjmBETD/i2mg7yY+XQQxBo2dKUbQDk9qjsjDmCDK0ajf
gPgPxn/2nnMsQIcvZSYH5Fil5satdF08XTJz+XiJie86kJFrEKjw1D22vURAqzGP
qsBZsEF9lAJ4Qox0NroI919k8YYbMM1YfroHdw0USJkLtszMDe5eRV52zx2V4gn3
A3+X63qqTJ53Uo54hPwfC1+F69jxRJxlSLrGQqi1JTvdBtQ6iNmlXLHrK3UlPO0X
Rf4gkjXjgL7wADZtEzJShbNMXd2vnZmFtVG7+R2ENZN0ufz9V6pbSNNm+JvkLhB6
eTwnde1zEro7irkw2dIEfW7gkmV242fjlJaEfenRxhwqWFMArTYtaoq6HywV5LMM
bJxxquFy1YdAMkglYtXpskFL6LfTfKTpWP7J9M7fzC66K5SN2nVLuXgPf++usWSu
8uWMUDQOqmU7qlTzJWRmtmhE7wlnpXpkm3zcvDBdHcO3MprQHss9dK11C2rNZ3Yn
CTKzgqB86mP0B477wnsdhUDBSiKy06HcpvUSXj2eiTAlIJ8yllOXUP8wA6fD5s4c
ac5raEwML2pymSfqCc7eWfqkAGl2Q5+P1yJt7muMq0Nz9Zb0w/ly6YLCyF2b93fw
+IP3l8yT2GNaG2XBn5pKEYeWdVb88Bcl9mInnj13cR232wuXuxmXQtbi77tpiJ4e
hnj92of80aLwVCXgKs47PgLKbtroO4zDepV1U7x05CEqLh2fgHXhwVi3KbPT0P1m
Uh5aTFp15gc2lMNM9UAvY2RaAeABp1jpVhxkCacGiS1tLDi+8jaYrZQXD4KPTt11
ijkxjhAqpBbQV/dHn1YofZaHwHA2dZISidOscJcKXd7z5KespnKjDzzg075gMJj5
nYZ3wM6BJ7jNsBEwadzraSm5idNTwpZGlwg5ExO4c1ai5A0xDJdH6gi5EdYglFvJ
LkOh6Su12skkit9yoG1FDrZxMWfJE9T+ABR4ano55iSxDOUJKGOX5zIQu/Q1r59h
ZXCzj/fW3GQcnPc4aiKiS7IhPnjpjtaJ086xJk3HI3cOFs8Pw2KJWM4VKnpUiK+5
PvQPdlOOv/Sy/ofKvQ28FUZaN4ywUeyp6nLwEl3a2njFiUFPpwbjOe/SfI5zCPRY
PavGaZG62CPpYXa6oOywirVjA2eu0/cFxznz+vLrenQV36aauULFo6WC+9jXKq8v
Gc4fKV+t02GegRgUZq+8TNcyLyyahhhnQw5Bg84Le8+LLW9oGDHBbdK+7OPDHaPX
ld0Duws4+YdYtbbdOyyt7wiajFKMqo6it0iogXaFOCQXMFVuyw8hcrVgaLRa+v/a
vKBZ62OQR5O1PGjZ/TCbqYZ2ijIfCK6GjjPYF5C1cO3UNJFTJd2aUne+b9e/oljE
p9ERcUrN0qUCf30FeBWNzPicDvNybDI3827mpbaOz7PjJbBkwiFt2GmW5I/tSeid
escUdyujbR3cni6J6hy9kJ3LLOn40gMqkXto2qZ64LN8y+Q9yKNPsChycPIn6TZS
qzWpehkEtAwDbohpTsaMxDXRl3c7LCCL1dxBkez9kKBnldy6nrkAZDQSTiNaVy7/
Ocv1lC8UoMqiMcir9czdvaZ7UMcBk87bCNt/a44dnG9pMqOVp8oOoas3ceLOkOSj
T9ly1fwCWt/D0MBaCNhWs0FksLlOmMYXP8pLjp2miBelZqZEA/VqWAn2amWVhlAv
mee9ox8gE5vN/TjLqCGjSzd6oug8W+9x+FJw0wjjXdPbv+D7s8/jcSEO5lBQhHQ9
38zWEckQVrYvsrSqTxRzNuSKcqoaYZiaUIyvPsHzSCNv6nxFZgKbOSdnDgtc5FAf
/2BCjOiO4SofTXHu43NOWAvyHoU2xbiZ/yGYA/PHKcaXH3n1etfwChxHSJasbFUl
jdRxlgboCy/3pWLRfKfJfdhOBTSY6Szoq6fbhwI9zjSBZfZ+S3u+edPTdrkQPNn3
mlC6SWjdn9KjL1rKtIrGdlpfidLBFg5P9dC3AuoWhBKz2hS1ZBTh+ZQBIlr8p2SG
gwxlrF3R59tnbtyopJSM1iNJpU1Z2GdBgyoa4HK1HunHWEUgms7wH8ZfSgP+N+1C
gx6UyeplWyAPxy4JsTtDswaBWtKNgeaSeV4KvwIQwkVv8fpSv1msktg4+h3HW9aB
yYeVCpWeOvJ28RtqvEUNVAIB0H4pjWd1VaI5bQgLfAz1nTzKNw/NlbNZS8zW7NxI
ptOrN1cBNHUEfSQld9lWS60viYYL5wW4qWTA5zheAyjlwUBADadLGqxp61AK0xKP
LbEXrXDfIINjpBUyT2uPYP81uXbX+TF6kIn0IPYheH7NWvbO7RxORz6a6ea9y2LM
otlkjuLSTu9rISPYIF8TE2WB6ddyZgc3vfpB6EJ24o/StPaMBGNXZnguJDXGWU7B
87MoevVt6j+erqM1cFWhIn0Dlpk8TPwHewGqpxQSkLBKBek9vHTN3MK+RRFZv9/L
gzRveAoqNO0t8QQXiioUL1cQKBaH4STYigI9WWJhxxMktSmLNgRrYzoyv88tMweS
8dhSDmRhGnrPC0b8r2XNetsc2HyedLCnXiJvp/0vdivPGUiwGQw3TQO08+7McvBC
tDsMxVeg1/+ZW5cXcc6Eh6O0ftH7sVOD6NrgOBPmIenAkjMSdzYEpqcoxJOvxIEr
aKwXm/xpf8jU3Bv9qj9TxqiI06bXGBMPRCoXMARQU0vi5gcbHwPl4Qo0GVWNiSUq
nWu0f7RxxtkaACOZ/92LQke5CkjiuUgQYvHL8lcoSyCDdCOQ7I71uZhirUlsTzql
LjRD8DqDCdvGRIJSlIJTppq7i9d5TQuoFImXwP09PIremMB2nJu+S/zn8ATvjRKj
yLfFPAix4ams4pHk62JQwSLXAO9oiTgT275GFGfJINyjSH3V/i3xk5YmfoGqIY1x
M00UQ7qeORQixgcBKIyxBr13wk8gBGAwCaLCXKA7i8aM6fCMkwk/uSs/eaAeFGk+
pFmfvkL92k7kAa7lB/EERmltgbPIWfRsRaQx1wMaZWsEWS0Jj2+FG0FbuPZIsOAf
3tFhQfNyDVWhxNP1dT+ljt2aL3ly0ZxLGNo0ARVIqPDIFY//VslIK1ldQzGuxrIm
yX5Kh0yiClFBFD17tVQk+NsxPYaB0JxWuo0rIxD1AiZ0MVlRzBqGEV7r9YAdiNvc
PrhUe8K8R4v+58gDK/TCsZE+VqzYytdgYaU3wocXRtkmV2tM1KUzi9JVmfDqNdjr
EwNZk0WG7pkoWpojh2H0rFdvo2m8hqi4hzPOU/HOhHcKhUFWSXdW7rG3LmSzTh6e
wRpJnX1lEevnK1jA2KbR+bh0ujLFzFm4doAq/62QzVuCV1PklJ0yDaCS3cCqgnsp
f43ko2dt1Ph/CyrHvXdEhnXT5imbTTuY0FPySoazLuPJOXvoD+p7a+vE8i1xvDm9
dm7zdoo5FNH34GIeZLXpbhxedNLaLJtXpKhdD5BOvc1ovXUpmHpZYsotBtCEPk2v
Hh1p9wPoyyHvNzfyEVAMvojcznBTECwz0wQFCoe2nbIZTWY5NPXt/PUBCa2E5MDk
tiDNNUAgCM1wyO0QQ6QoAbYANEdcErsTy6mz0KiNzrvR+ImiqknoL3GXBHLWczLA
GeIgDr0xlVZiYH7xBg3kG1pV8zRltTw4TZLZD1lY1+cK131f/9bly4/OkBNEzCdh
Ng4s4FQ7/ORFqIlpV/BvMDEq7IIz+NAstGu8DQ5lyZRiC60gIx8dr8GKZYb9k9ER
xHsAPb0SjsczP9yddj75Eqck4QEo7ZOVWVToasb4W8OSXyRU46HvX3qZ6p+kRFZ/
snoAcVp8vutf8yhJtoYAd6hHOVUoxUNTAkxss53lXy4pzeCyonOzGfWZXuTqofqI
TiWqHgzvKEVdPzUZO8p1Zv1E2TB8YbOD1OsjTgDbzelXpR74wMObl6xXxhWri85A
t9je2jkWHb8Mbsmgq0xUV6Dqx30d+Pl/7kqGmMp4/oKv9aO87XImt2ePlOkb373p
m6tGYcamwX/Lc0ivzK/gEROfkT+lc5D/jwYceCsQ1Jns3jODeUjW0D3f1TEhuUbI
XxJZbSjpautRtfFohlfRsFS81XxWGmDU/K5E8/zRFKJIb5p0oVAImMXqx9pWB8yH
0I5bt+MFgK5Mu8Kv77C3AyjGRXzns00XVzdl4zsYo5GpFH10eCf2omdSotNe4Drb
IrM1Bol2bMhBnQHQ/nk8Wbpv9MJkNzjdbmgdUD+oxn8JRd+G38YDSTd2YZHGGsSZ
AbQObdTFxf+YYCmCFP3z8rlY7ea7lVDLsYPQs9WgC0uguPeso7ik0xE1fu+NknvU
eK2B6RCPjx3g7baMdAHz8QGNnSenzmUazePt2iu2UAes3pExBVk3732F3w61eT52
bCni05c6nOtxrcEH/8DwXO2VoyjMX0d4p+PT0RsIO11CYM7O6nBXQNi9iB1SAlP2
HUu2qauQQxwcG2pMPB69JaJr3z+G0kpDoAL/RiRZ3JCuWI97neP/9Jh1E7gKzSpU
Ua0VeVg+0JEH+CPnsnyvN5HxBC53xeL+kP1lkzDHJN/QGbqm/m0zXoT9tVkbcQOw
esT6DkpFqlzyimkDSVtOI95wUrQBl56kzUL+OWYsuysyuSQYMNLBdsSaxn1qSCsW
706JnDrQA2S2PrQDOCpKRapXoHytDDii6t9ag2SXE1+gXc9+vft2XDDvLrfuQyDd
nGTbcCpdG61Sd5xOgVfldNgzX+NV9hXYygacN4yUnRzSPMHHSVp50A70OfuZeCfr
BoG03+GPFPK4UxAQZjQT8C/scdoVYZPoBQf/WOSp9cyCt4zbHbmuSZW8czuUA1l4
lgwq0bZB6KVweAnMOd5LOsJUH0KF0sYmPrgof1RfY1+fOxJuWs19QQaWN929UJJl
cRlZGSg30EbxkaJGKhqo3+DrINlQqzBcnyuBBHVQpOz5vMpFOEK3zabgponFqZZw
yEt1gZV4CLfbJ6bJC7+Nn3Uk9ANj141P0nNR39IUVHR0XW+aiuyvEVfnSt1qUy5o
JOTTUPsFED4s0hYDFvYI0nHgzCSP2jvb0UXz6nXcnJGLwZLlnrzHhxgmOFRa8Lly
JgyP5mgRFFU1htKcaH+tvV5sVNVmArimQii9OMN0t6v5pHn/zxhIJaygQ/m6DUzT
X643qFjW0RKGtd0bwRsypjANg0Mwz6mCt48osK8lPoBStSZNJSnEfuh1G5Kbk17E
LrPV9cID2sPMjUJRx6plK4rf8L4oS8pIZJFnxg+Y1/orKyoCTJrU6FQSFBUbaSX7
7rdeQHBq+tT6di8ejAeyLSDEC1JymiDBjhJi+UjFTiDzgMum+MkrZPb34SDbWN0N
wTbj1yonrusr6Qu/CZ1POlZa/nw0H8+FAiAsUMHpSoxtXZjCnUAIc54DruQzDs6F
lfNt0sVNagDCBp8ivWDBfKIVdNZNiARwS+bEBUYKyu8fmCw1eT3vCQ7lK97g36WD
Fgd/Q8dtL8NYKBkSResWpU9oM1IDrXu0pyEPT3e7+yoAbnRLIpe2I7phpsnI3UcV
Ym9vasNDvKP4UKgl+rFov9oUwPGeDPVV+3MAFO30IpI7VKjK13FCJq4PADSbcVPm
NuyNgp8+XrE1lGZ/nzp/FmhPEkMn5vSJTp0BYBjM1p5Ar13933ef33ScxrXRjDt2
NrBOp9MSpoWQ4PeRv2WxK0iZ8Pq7i2tj44JEJxTI5k59YwAI+Dy8z2gGLust5ofS
HpO4sjYTFBv4j1HSNraEkvBBkyQkqjLzJnCW4CcaxZhSIVAgNL3GNwKe1bkAF6bg
5k/sDqDk1u+jLKbLMGbsYkOGiUbeIyAJBZDCoOvWB66/RZkmMgEMOCeM4Oq+2kB2
gGfjN9BGrrH9GLi17XBF56P7mMxTfO8fKweJC3eiUE7y6UPfF2BFwQ91XK8ZRI6N
3JvxD34XAtSAihuYOzyrBGO3xLHO+KWPRXIX4/LLwdZl8Qco1Yo03Y95fQ8aoWLC
fTPNZZH9Fwd0ABrEZ5qD5BLboxkyWLbImKoiIupB5p/uJeuWWclSLbX9BH6coX9w
jlSq4+B/va3lYHGekMRaJrATb5DZcDy32zH9hnxd/XFufmNPteR6JHfzlaAmscw1
6TTa8FQDGJZSRY9c6QoQ1aPjOC08QBgdD/xvaGRxXUfQTf+obciNidfPKz1QzKmT
3jZGAR9qPp6K15AHhi9MNNPG4hYI5tjiIkTaxh4qftXhS7Zh6c05WVcLaCSjku4r
nleb5fzC3k4AkP3BhPsqV1FXeWp904zLn/Yvs8ong5FpuJ7l3TAopkWEjFt2AqwT
z//aYy52y68l0+XT+9Aib4yDgDI3skxUURhXh+Ut+i50mZxwjVQn26IbiBPchc+U
IlDt7Cd+AeBYFWQP08EHHEDmHkD+NOhLoTtlIYwcUfdycc96c7jOdm6N1RfOc/qp
X4esrRZfg29RKkzXzEOPVN1jpGZf6iFInbG0Ac+QZ+k/iyzT9Hh62yjImvyKhYs/
FCUVuTJqIf9DJrUKlMYFgtcwOiabnb9kqd5wMbkzp/Sr29UaQigKjSYB0TDi1c2x
hsWUyQNJJaSonw6HR4lt25KQa141YvTcQav9K773UE60t3QGkmuN/Ad7V/HynTVX
Ob0fadCVdoFsooRVnZlW15P4cVLssF4uOxSnsrSEcJcp4bFjGaR6YO17Uy+UB0DW
4yCkLcHdXRW3CpquHEIQP4MSSdL25ttijboDGTixjtCIYkAdQkZXANpr3cc1xxxp
RLWyx8lqfqpB4vimjBg4y4BzLgo7LcJvq02pmaBghV5l4CYF5XlT3RJuIyrN4l3w
e17LEJRMUAOu6Zs8XXzEe+sm49BV19R1i1xsw/njy0hwe29SpleiLfBME/n/yKm+
E3xjM1UdB0oqImlUwCgQbHA+oSocT9wOE2G9FJQ2CQBixccszg91aQxIKEmdSORD
uniLyOCsfjJnLGWh15KtpH+JrQNwLgXVyHOJOXS52BYKYS5VhsANyHEEL/zg3+hD
4nWs+z+hq6UcP+T33SSDWJDZ7NvZgbc0RRapxOCFSXHG79UkEp9Auj9Wa3OJGBLB
J5XZ0E6VZsixekliZm00Uz1CexqoWYB2dKJSHHQMc3NIkdxjrwp4A9TGQuPxnh8Z
m7Ak3a479mNj+swG7JVj9JaZ1mJzDwDuNgIXMxLYpusgqErKPd460z81Hd3R1CS+
t3+89kITOm2X8jqZ3kpmTBEVUPErCe6f6+7NtsB4pXDC02czaf8WReqhc38gCnoa
eHlLJzJ7F/SmgJMU//mnrALdJ9acug6ecgGE41LKRufOpCdGmooQPZh4692lf6gN
fHzXTumbLV3ofjkHxk6MRoN9GGoOW+DSqdJsvxfYll6aAna8CkpUY6YkTeZ03/w8
FVjvgmAD1eiCjXytbn4bNbtuCxikq+CO7+kSysr6HRo39GTedMlIQgp6yemvenGa
cQaWdvwTjuo0ybF+MWfysT6rtGIu1bNw1s1+eh4Vg71/60KcesNspCybqUOIQ9/I
8QK6nbrb2L4V/DvMQ4rVl/m07DC582yHwEnnj59E6psVW/VyzapH7f6s4/udNBXU
ey6gOAIbq2jhbJyQQ7+caOPAcMnIpKQBRhRZRmpcYauNQyOUhQ9zGaYGT6aGO/87
DrY4pSfgipPqfPcoxnGMpLeqC8YdFfdliSti2XkWlhu+PPK6e1FBmEG5Pb1fz5Px
/UU1kHS8xED9iDZo2OX6ayEtRj8CG3/RzFss0Z/NFg5AYsAylzDQwAZeKWMgDrz4
KXV//rIo9JvuBJWi2LdyKrtcR+Xo2PaKmSOm4xGT4uFJMSeLiR9FWgOKlvzpayCJ
RkA6Dcjv7Fb6SjPxC296vHFWvrah0w38AkhOkjiEEJyoAi3dC3ZiGYzV12NL+m0l
vWaVve5UqtRE1CIA6tORxEINl9miX40IpP/MqnoafOkT6TkcbbOp04xkUvY0Hx6v
dpTSAz7VcERT07P6Lg+rVfRS5w5p1uADodje3s684Buq7XK6RQJtcJTPwv1kCtKO
TPd7gWdqgQYLBGLi1as6BKWJ5S5V+ec4+MWLbEPMovQZjlMCi14ZVxdOJ81KHW1F
vhRXL3aTI/3Upjmy1n+8igD3aZoctPtJiMATTAvkSd9DfWEoh78aesniJgonIoQq
m1sr57gU7qXJWQA2xldi88B/gZhlGy6Sy5b7LcSAi3PMlsx6flbGJI/pibk4MgHq
SMp1EsLvbH5ZEPz37JS0KeVnfUs53dUVs/dswLTJXXuWoyJRtJLwjmwssjBIF7Vs
8/I9O+r6HfcIEhFr/WrRUeWBPGzpBL8seD7fwYfilOcZqaYI9t2YtBX2RIm1KUxQ
X37TvE+uYcWEoPi9Zz/wv7Lh9SOSzfgmNdVZl8oi/UTz/7UbDNM6pDXQWCRv6/e1
LtlbglIr/esBNNzq9BlwmZ9TH4wcAutqebDM1BBRGWeTvEOad0VGqsSyF505PBQW
buX+5AtxKvyU0mu9Wflp52pqDE0sLWTQwr1phlcPWVmTnk2CKxR3a1FLxi+nRjyM
9lxmY9HtTmRpvxOHjFjN0NTEtoxMRCUG7VV2Giganj27mhZxJWOjZzVx0M5+XrP/
+kBJ95U0pKZ4WqX0AQLssh06/xFX9FXHkP1NC3N3KqXqnQ3py3bLcQMsIBpdtNHN
cLucfurb4ubUkstjBnn38RTIoTcOJvLu46fXROw0Sk6UnJ57IrWD9Tdm0Uhcl9DJ
GVKthUJN9MTNmu8JgAFOPbY1XB6cjEoSMtGO0LNDceH0dEXrngU4dx1LMuZe573R
edw3l0wixU1KQCMJUKKqnaoxEUwmMwkS3vXtRdDQKNr//d3bVkatlSrUseL9XPg6
f6BKc3wViO5YEj2l16CLydAFBCxksTpGBVqPo6rLJaua7WIonjhHoO+U5BM/xn/t
ge2wPZX00tFiQfCYyFMY9Ggip99/Hz4CIcqjOpyS4y6E1JRudLVz3nLdTF8b9/Gt
fCETFS8s/rBd71OUHV7iikJXAtu0vZq8eDgDLbv5YaHblYEZpqY3eZYv7Cdk18Nu
4Pme8Fm1PWQFjjKqQUu7D/OzhwffjP8iOYfeNsmsps5lFsJYjGfue83AeU0Fsr4U
9Y4VPYzoGXpScrfV/71+lGaJ0fPIwHiOP67U3n2NanXtIxpbZ9XilVmwvAw8vk//
GYLoRmZ6fXX0wKAWn86cbwcA5rXstRnaj/rMVFkik9OD9F4HR5/8Rw34G9OobTpk
eFXgaV5u6rFNc+bWpwniUbeNyyzGIhkYgloSRjiJcMSSIXGmUXHIj9oVg1iej5k6
P7SZYVy9BfCOfbN7KCUuTAUXqVWf6mrj7lGgk6t1yAGt2EREz6A+pwxb96yp9LWw
hYGzGWuhTkCHF6DOj31nGwP25bs9G8sfrkX7LWjBeGjjBXqKC7ySVqzXAO7OwdNr
IyF2Kc08bmaxKM2+drOwYlsWMnDAoGFCl/l1/IUquP9WhffrZq6Rlmc+CuE8Sh+p
GUdX0CzsZJ1y+DJcBs5Ccu9ws1UNbwPDN6IWwYb2ChckUdX+husAzbIdjswqqJh0
YA1b0BOUFmq1fc2X5DSYocltnin91nb+6Ib+waID2rowWeIbdZ4WNjdA4UzVawdG
5WMeLrO83TzXVJJA9BFcrHLR3YDzWfz+3d0cf8RR25msqWtLt5PptcsT8QlTnsDk
r3Rv+icx1UlV7UCEA2k/ZuJhH8Yd7jq+1S5syl+M2l381TjnOR1ZbkqtLe6T6A7u
FeotnNgLD3dhNHhU41yJI/6ISfZVrMucMfA+boTJpn69LEYosL5dWM5OuFxrOqhe
yQEM2PyJh3e3Ge7Nnikh0n2yohXB5xhoVOue2kIcv/a1v8psBMH/kF4TrycqjW6a
kHUGU7/1ysga9QIOysrJAmZTVJk9PT+w3OZZuxbUFVYfMwbWlAx0kfqPpC+9n+Bt
vGNiwls8QknNbkKKsZ+AetJ0sXh87h4+FMYhcC9YmMc9F59WBzFuO/JTXs0NODiq
PwZ+IAUoXUEbuAhl0ytk9mWaYVjWrJlAk9QhPKWdK2LkrFB6gifupKVt4lC6daVN
dUhc41EHZ6tJgg5/rW/maXoQkPJmSyLEdQKZi58OSIHWPLHvhzQW8O5P+uEM7lVX
f2jLg+6RgLkKRdA2xQKVzEKI5ETdN7fJWdGiMcQ8J95yEnQa4w+gIfG93LeYR6d2
fYZGZ4p4yoPjvXWNYSMEtWtHRtppQGTsQl9spdKHqkJ5vLrnNQAH/RxenmFOj/Uo
MOU8GwVXUJtESQRNMOhQU+RG62Wr18VMx1i3Hp2f9v5l4mWUuAPBYAfkkVUd0SbE
PoVvqPXkXvONcNnJX8yYm24+TFEIoEYG3/AJHL3Q2/z/3bGV65FNWszViPCjgIXu
x4EzZx49PUbGL9vecmsvwUnKjKNGTcsjd+puwo7nxe50Ku4Ebxw0RKdy62vM8dNd
jYAZmeSYU0wn17kssIgG3plTfSZE4eqIzbU6CBocVNBrKi74G3dVu/jvggBeu43G
Ec26FE2F65pnyVJab4+VmIfmlMHfRItbFYEIcmGEfBl3N9bsrhkPVmMfXy/PliC4
6nWR1Wueme67ZBElMMcC4XtVYCx0N9DE6u1mw5FVQnWBEeZ1afDBScTJzeqF0EKu
05y52Xb8kMNlLIanX5IDhxPDkISVCXjjh5XQ7h6o2eHcoGikjlxn3Ydl1yUb9xN4
w1/d3xDWHmvmwTMsDCoFwl+p8LKi98q0/irnIdTbx5/X+gp8SpeAk6NnKLqWHjlu
MqXtqKbDlycOVeMyoDmXRAPFyImTxfDUGnMffHjj5GUaZcgqLDh/Slnrz9FTh+BW
PTnnw1DQBMXc76AAoSrBecXbE6SrRW/FS2fv2M/5IOc/y5hw3AunqAhOrNMMEkXV
aveZLES9OJrXtNASk0MB1MX1FVRLb12lM10JrsBGxtuei6BKj3qmD9dh8waQ5HAi
Fpo148gnOKNZAKWv+pbpyjWmq4UlCY0YJHEYGJqleGPC8/IG4cARLDNkNtNkizH7
4NnsoNXemzduirWfCD/hzVymf39KH0DevhacVdLh0Cl7+JRYnlDkARRIZL+K8lX2
wTru4b45gZPrwhBjZxoR/3fywFZEMU9B2ex7dX5JbkQwINtrhwtmqkckYW3+MY/U
H/tiTjKUIKS1pwXeolC8gzIb3wSG4wSEEl6tTxHTpS5vmmWzjvP0ckkecyWYt6Lg
dND9rUeYNJMdRbn4+JyQ9iPRSez+KrQcmSmmZiW78d2ccbQhS66JL3ds4khga1QJ
zGeUZVT9jo79wMBoF2Jrike67JGHic0Sn+dgTcRqgEzF3oaVp603DEI4yspDCyOK
KdTM5vV0FVBO8CgkgBbDqk+cG266xJ3DJErPWXSn3f5SxjbuQVNhIPnABpvv4zz9
3h0LVzlz1F/XTxSUUTQbgC3UvpH0Oy+9J4fd4qkh/usWK91oHXk33p9JJmMjDI++
bPBreLWGDfHi+NFXB6QJMJTCiJH1Dh/5xOl8nTRhQQEXtFUDulUAq/UkLSNWkwY1
WVGYzGpbihbdt5KvspdD+aWNH5k0YZWddN+8qpOQQRe6xRHg5qvEnaISiwxU37Rt
k66f3wxN5wI+PIY4lVGJFhPJCHKK52DrU7BmxstoHgIyvrYDxGigdcejgr0rR6AY
uZ6lQXUtU4Nbn1gXIuw1y2yaECMllwdK3yhVimZQEmGfhyLsTSVbppj+Znn+XLI9
hhw8JZ2L/RjvhdXD0SIqBpf/7pNxTPiPR7iJkSu1TRgadDo0YCUw6HrkX3LdqQiQ
gPhU3EKHOH0hYBJ17tT9nskhL34zpPoELLYtrL10BN5IWkJkrMT04vXwfGNmO4BN
a9TZ2SPy6Mw4y4Rp1vHQWtcy/wa4uF5GSk9yjGcz6PiutqrmclwMryQF9hBSIdC/
XE74DdCvOe2LN6daSjoEoSy1ZS1RE/MKLmlcfXlEwkifGhGyOuNRlm9EAzVpqmRu
g+k0gptPxTRZKhqgsCT7fDFhQaPvKjT+TfpIOf/gyV6Moy9f838zpMyQA6MP6VNG
VlA5IP7nY8yheZMc0rxgphdCRUcdZUh5OCuW3cjESMT2sHYXdGyEGcEc/m27gu4a
USOmzlu9N6C2XKeVQk0BXVe175xWhUH+mKIWemFBzlOeix2/ZCym6Q2mI9RqvVaW
chknilHlecK83+z+4EKz3FGRJ6alz2QlRhwASLk0vKZlrnF6y9C7a8MFYFe8lODL
qFeUE6l7RDFPChAcukS4uDGRh2uqvtD5iNqZTNBM2XaAkYDNWa7feJT7HSvDfmHM
cPidK+6LoBsTBnxHgEOXolOQHe6KoWiHW600BQcy5AfN6pKLdw+/ovzSvifeFwKf
qDYa4WdjwTWJylRAyM26rauPF8pDwBTfDmGhm/LRkbFRtBGQLhCfzfg3mFzD5Gxo
OJ8h+xmimqdi77KkTB6bOgSok88m3E8Z3Rk2V86Gq/nHX1ZrIucKn5D8dXAiGfTC
JomedDmP9Rf99TBdXlDmhxqD194ZfM+rV4A7bcu2sn5+tYx/DFqp6qNsmjB4aYTN
XkBl5JVHwi2l85kR8MXm2SJO9nmq1jVZtT4CxP2Xxg0Exz54N9YsGIMjJFfUybmz
KQODEMMQZsIBmLRNowjKncMtzgQllsi7lhy6DoCxRb1iEDmA7Bcd9YHQWHOyVp8B
uBJEGD+hTAczeSnxCQGN2yNdan8xQd1sz3n1pYlEybgW8jXvnwCcMHAvvX86fm7m
VW5EKk7ET/44Sq59p5U6O022wPVB8/uCrFWx4qnd4TTOGTNQtf0uBXqjcTA5xRk1
dtxipnjK2cUQr5Yy0fBVFlsd0CUNYVjhMg9S251YFwo/ajvawwSiDUzh9pjvuscN
6Epj1hJSa3xbAjubjl73+Qs+JQs49W6sN7YQpCk66hds4KLrpwb/cPrru6bhwX7C
9fq+zEbRkiHSi4134TiYqfqci+r+zOSJMAj1DtxoiJsgjpC+PWB+UMS5BomfXq+M
tIW0EeSvbREHFNnBOupeXIyt4zKqGucO3yUMn1tYuhSMkWovBNIkYPhHYQkmiWdT
gzEHNo8/il6P6TWu04+MWceWbWuFpATLQosATQKGqfSzWB4zdWCtN0+eYJtuRxmA
Gr9aTZvxt/EtoYX0I7UHzA4mCe2nEU5CNtN+zsPeQ/T9mT+XUxUUN4oxQmHJMpBa
s1heJ6shu6KCGkAKCISxOLsz7GO4eKSNjny6zpVoXJ9BBIwQMDqhbr3Tvz25FIYb
5VAtoANd5q47CSc3KbV+PA5/FfPYNxj0Y89RtSGmZyW5msIQmFd1q+foZ7F9FhXL
b1+Vum6/9Q7Fm9kHGqH4870eAQkfxuEEow72xxxsHu+Yn2SFgkRUBYFxF/RYqFFh
tSIJPUEdeqIZqs0ipHLVNifBLuotyW17DeArtLR/Ub48XoYZqBnVdWMRDjISfXPi
iJZrwDUgfO+36lkz1AeDLeE1nV0EKwN5CBZlfrrGVXgxCGbCwO4/Pz53z3qOMrp7
D3U8oUbqGdnQRQK3mrZa4uGfEb1915F5PRxK6sYircF8qk4EcVQCatsQLZEy6lnW
7nPYFWSLRcvCHEXd6fepzGl6WwF9e5f9T2sOX0AKkFspQnLSy6+26zkj33VOMf4+
xfyMYldhf0UrIFYs0IDA0MJHTaFJwUVPvTNnHQbekN48dI3ap+HNt2bFhdWO1zuf
xcVDSMZpr4bPRygDfBKO9/UXAUzBgasDILPZdepjIwgpZulixsPTvg7GQQULMWJx
b1UZ9a/MZ7dku9cQ/AU++9SB1va1rIydIfg8XRFscwcZuOS9ksok6j6g9TKur4o0
Y+EZqHCyFXLkuxa5zlq1s1P2w/v8tXPwf20zL1zYNMWqgafiH0IMMsmWLes/oBAZ
1byrD/DLRVpyM8bwNdtdNJ8R8bFXjIOEiyk6l3TQP20Q19cSf5irHUFnMJ9wZ1jH
wF1pvJOc5/fFrxv6+fdJB4y4PROiF9ewNO4iJm1eKBzLdz4k0a7Goh6qWAmbCEHK
OzWL7J1owWUCg7JoXUbtaJm9x3nXFFx+YGDO17RLf+cNYmY5SAddCh/gVJQr2VcD
40/cREFKbOiyRsh76uHSQ0mGAUufFdiLPeIV2VbjGN0MLoMEhWTasf/b4DjZ5CeH
6c1rpfUHAaeCJ+es/IyTy++/KZioTVxw8rIh6hipPnFPkC2Cqh+gX53Wuw1ZMKWY
DDgm61+fM3dARJsP5s6ZJe3JZAD4+r7xGT9x2mViSg5KmjocG09gK8D382skznSX
+o/5yIlpbVIddAPeNbJd3AKYOfheb6dOMEVy4Ivh9RzW4Dpz/eWEkMK7DCUJxh18
S63X8dkg892W4B0hOnTkvBh8VaeE0p/e/zqAjaJDWEb6Kxyp5/xniPHR1dC6+rwD
0il1Rak5UkiGnxj1unr+mb5khgcgDUE0qAlQI78b4lcfJ0HfrIKCv10YVhKvsx2J
SQHA4AE/eRfye7C9OhQMJFcxuI9K26htFHDQ4XwZZHsPiozKdhgr/25BepgFgQyq
R94tzSMzrx1BP/LJA/qaTeYl0jva+QgKvmbfeQgPnrzPuv5aZgeezcMhO7X9lNNJ
PSjRPjFnxcdio6HedV2Cr0eLJjmNR1VqDUbX35tZ1kMAi6LPwLP2lO5TOSv2gF5t
kqlz4u6s8xO1kxLps/lpcbYPHOjzMYpdgG90js38TES02XnHjDujuq9OMNkZMcHU
NpYApYt2zFzjsF4EU8J3KfPkyrMcWbyGzAsrBR0zbN70Ev3yzZagOWnZpRYQFqHh
eCTGmo8fbCVZRfDx38+sjr64KDZsFDbPYEvDRyDIYJpQJ2swuGTDgvXameGcgdHN
Ki8eLAo27E7hw9dDPAtvj+5ZRoX9K35nHtQyOOn48ivjkZf7ZHON7GLFBPHjSTSz
gNydeci+mx95qkLkzsxnn5Xkgh8XpaRcpUViXDVR2mXhd7qnEgDVmmQ4T/QScWtc
tf4HoHRIT926oMbrRNtOlgGjMBMn1bp7MAYlr6Hi8N5u7qBg+Hq7PPbawlALVzqq
i82KEGThbDdzLngE2YJ1zrI84kI56ooY8EmtfjF/b1ucg9M/e9mrcngegqiOleTg
G14z0vMvDL9Ad1ysnmpJ7A9VDyZeiQKKfFdGr0foioX/v0XPieXdD1a2I8YUdrE5
KgsXCAjnr9pTNtRcwymyoW/MwMeKvpYTZAml88acUYU7YG+BOOPX9JSkjcozqTQ2
A+ZUkBtORhvHJ1kTUGVpF9ja6vijr2kJhA8uldXoP51w2IDHqBN+HX05J6qs74hA
fiteMYjqlQ+f1fBsey+b3dJFUEzfFxg8P4jBmrRbIDzArsKmzdyZlRgSf5Nz7xP1
cFu2BPJeDHgkG7nIcARY7v6J4LS0rbBfj3/gFKeK7MDICSEeDFh80PxF5cg8L+hu
N4CVErXrxvJf3UueCdN3vpEyykRpUzH924uwuKTGtQeq9ZSecowEX0dgdJKOSSpN
uwz58hQCIm8/SZVJjkVx/z0mIzVcGmlpWuk+LIv+PrM6DGRFN+Gk8I0Uy7hn3KUo
XyCbUsTPlsN8Xi7qiFI8fk7wdFybp3fSVKwUwLIItZYpdJJslpq5/FK3/gnYQGZD
MAP7yFhks69D22KkL7jrsuTTdB7aDfg1PTKK0Y7U0ihGazoyDkE81OgeCY6r2KBL
2Xl5FRwBhi/iwvFO8JEBiX769ra5lg3Z5aF5JG5iONpHqivlPUIiyYH1IiEMPnDk
M6iy0AuVaqc/yf8iYBRXUOl9CYm2bRT1h/P9S1SceRAJzKub870dmqMPyle4PSan
YspJs8myjhE1PKcaaGDrPhBm7NqNiKscPNjoMf3sdTMluWUcz+8cg8ojjcUS/V9B
o4MkDVSZzGBhwcg2o3aMiGF1Qn9g4gdT6w6m2RupyINqoxaSgKviETgVCDeOqcLe
49IICTAjGeVgXVqc0lwAKidZdsNk8KlRJcbSWPd6RtO10iKKnordkFRq3lyJ+Xuw
g8xTG1kxhTsdbJ66yo9jWrgSDSycP1IP/nm7iS0GWGd9Edr/BXzjABevCNyWQCC8
Wy0wDjM3NXyY+Og6Her57us3mqx1RH2v+bgMiJDTFylIsEIxNW5a/9Bm4istwKnd
sKJZaentTAcC0NCgx6qmy2JeFOb8z1TX0YIQwO8ya6U3NBoY1IYF+aCbVd/+nNcV
Aufk3C9/CRMi80fSJB56hvQH7bFk7nXIjnCMK65qjbyGfSmv9fWCZ3ZXp+GEBkM6
cZshGkd3PNWuT3oJOF+ZoSeFt01qWBVUMvrIptnnOWj3f30wiOKlKxMdTtcy+Yva
tCTHHrcntAWj2aPeBTjQYpmRmmiGDFETld/VjEHoagwsxMph7Vvt3jCpPo5H06vh
jw1FWobryVKbxDYJx/s50hhyISZFHPmFyTjWMovQjZhOjZKRZ//WMhv4dDXjGLZC
UvQVmPfwF878BNy8iI0k+92wrmQcPvzQ5WDeLXRMtjmDn7tzKle9leWibIRKwomL
u9xtyqTUNtCL8I8N91+zsl98W+SGCQTW+zaaMoud7/TgsTQAI+398aZJPtXIob9h
B7dFcv5ORq3eo9hcYTCeL4WeO50TLpqYB8pgPy5cLf2SuJz7etXSA8YO/FA4yv+2
SIovvhbRw4zj2Awyj+5+NbW5Ayuo/OQErmxmZrVQBfMkKETINZ53blV4E0e2L5dO
wlpnLsBHDicaRyLDJDDfay6lViQ5vXApdOt2cdicyxFQbSyizxtBPA0trG1eS7hr
Ggj1h2eSrAAQYkUY2IEv+tje5xETX3VGUwUPitI2/zfOPwu8Ayb5iS60xJfqh4vw
gdlf/F1NfVIjBwEUeMaVBkp2BsWDFCtVP/XbTsLoSKhPTgwk76VRZNe53fY9+9KQ
c85uTgYF4bh9cMzHMZEKAFwL9OJPMg42OpGss9ta3ElE959TrCGl5jJ1fgNwIcCo
AmucpYaoKTj4MsD7kRsH9gQE1xwqR9bU3cVc0ijHpGdZR6AolFYMv7kN0pUixBj+
tgUfDp5rdX3T9kOKznV1miWxkUAAq3aZ7HKsBik6k9bSeqpym7RXAyIHy1Yu3dkh
TykHAfV/1rEoe7sFVSnuWn+/yYdvhOnqa3hExV1XNyNPHS9NLhsYxt2Hkqpnim0h
G6TCF0qFDgtOaezgUOukUEFyX8kFNDzz89Wm/SrKZV0TZWSuousGslkH15EESSOi
Q78uKtajtBut/L8YreK5HmqkYX6ixmrVoKWj1+eOBP6IvcD3LSsXvWo9n/Ek3xsy
CIApBILz2wuZ4ASVHCXIidYWEx2H8MkD8L3p3ztXjFHmOiEmpjhkNKV9NNalaK9m
LQ3BHtGucn82MBbm/vKzK+ge2qft7l8d33ueRUhWyvBA7komgUra2TqjSBjpeS0C
Rjw69W45lQxrp2PjSfvo0LQ7lfpr0kBBuewBlNMu1JJGShYlbsGkHZZRcgRYUdP+
Alo0SR9YsqPL3kk8Sdo3ef5ntCJ5EWjmp1eO/S5MMhwf78S3Sd2e9CeRuewYJ0ZU
mDfXofkOIlzkDwVuUftcopntqhWCht9K6vw47+ZEwSiCYiwLLmsFcw/2UX9oeUHV
sdegJmRa51TNlFXJlFp6TyE0GSze71PrYpRiEaSjZLEbKZJJQVOdW7TUqJuCc6QK
DNfKcHGyBpgnV3UTEzHfETslRA38nSZzJL63tLIEVWzyZ1FqdOUixngH2/LLlj5Q
BH07InFB55aD8abbxvUefFPcORVvmbIrSfH7E2zgHFJjaGa4rpi7KW1DiJU6WAZg
6WLQa3sdA5UZz6TXFiJWKp0SgSSN1Q1BrpvDAnMvZM7f5v22jbeORcPuszk/rd9C
51NYpISrisBgrLLUO9s7y9j2DEalNh4JUYfNQbxBQ2A/s+1w6p0d9e+K/Ahku6RR
Nao1HaA0IdW81+N1Z7V8FSkft5rnZNCOlkLU+joHZnstJlUbG+YxSQI0XFR2Ni7M
RKGIprBmbhHOv2jgY53TuKImhdqtHpcojLM8lKx8fjZtl2IjpTmS8XDBFUZueqSq
zehc4ixqJFd1U+/dWRcUu35yDaUVA8E2hkdt/QNsKd+vLvsegWfYwzKm8TFAzWJK
a8LsJKBtZb+0Wnh6yZnFHC2k75EMTXmk8d37b4xlYvjAY/Dz9jN1akq8pX71mBvE
3XPzXwc/5NXMJC+b5L/lWdIzdKQTCzICihKXvHR8g6wc5E5GpaoR0D5TqF2R2TFA
oje47vmolZFRilISjBHIjwu1Jcpt0Ij7vAy7vO5jTzIRd9P+OQx1jTN/QJqPjI+Z
dRS4lzSLPBysdGt56QJ/rZUNnRrWVfWiDlgDLWX+nkkcRelbr90q4s4aK23dc+W4
LXDaEIwSbV/u/HpzZ+jp2PTFo+9SSFk99MUTxvUB9hchIgK7HvswioX0xx+UViKA
jnQLDgv1jePh+P+H/g+OykegqMEEOxzhOWbWoKgaw6daBcdDvQnpCPx3jcArvb37
jP/az2v7n6PLDqLYZ+wdZ7r2wGUK5EiFzSLqWffPVubkOxJ3Pi9rWbBocLihN+Pl
rQuxYSz8pok0eOgkpnZklhI4Rci1B29q5AB+VJCUosEgVaFpGQxEC7n8YAGf8Gec
pjU8yT8AsdGf1zdfVr2SNql4tbQx7+iQvl7KnyhGSfB+MJeRgwRInD9rjYpwULnY
R6lX5OkInQbE4kXdqX3lQxLOQ5uXIMpnaoL+ZmVKbnrnWbPJ0/n+dnpdBYActrwm
2nqJ4Imge+MMQbSKJixyuKA5fQnEqHMTb1mPcKqIjjfzPTk9gliRHWS+ctOQuD1Q
7SM/0HdBLPFVzJ+sH+mH6XJmR6WvJ/8haxsaHOYsSAsvXZuIXU/JgyPDlokQYtPR
YVGsZQu9Jv8EmpmxXGIHR7gNNEFXK10ag30ww2a6gd12V7QKC86QGrpn/v4/nH/4
F3Sh3Jj84+UndVubSmjWyvEveTXaVy1pY1EcWi0nFJxv5u/IHiXSPVs2pv2DnkAW
gZA92cWlW3ZP7gzhd2B4Py2VSWlcR3jSiaw2mChNOGidcuhI+y4fnFDHbTc6Hws1
ibv/HQa1X61528z5OPluy5tSsRP7H4KzVGBLmzhXtp7xm9qoml3cMPz/7P1tCF1O
sLNMixmIs3KfRRw4mKTcA1GwshU0M8PerlVh1ZU41XYqCgmFYWXzS200YdNwEDFV
2YnMeWECaud/RYJoN8Ytq9TzKqnZxeFKhIGW63d1tXqQhDRFGlhgZDWxjDZp7mij
Is/w9IBeEXMpJ/yy3cxd8r8DtpN32hvOtxRO8vHhL2N8Eh7TfQxY82BjXNOg8Hek
og1RVQbnHEPFzTKI0bD7qhFGbZ7WbxpJjDLGHpz0wT8QoJPSj4FwXefcHN4gliKX
tR1FNiGNWcJxEp9N26CBqvqnwcyareDYjAwQ9cI/9Qcd7WLIhFS7lh+XLZiHLLQl
otlldELJ4rG42LPVEql8eKw19CMIRoK1Q78tUhKPXS3hrGGnLFi0yF+/6BEcVwYT
Cu+X+3fDvUttvFSBv5Jr/5P3b6e+hz3kZDvBp56feL+Z/N9+frvvSlys7zeCDeQZ
0g96Un1S+s/8YU4P2Grx4/8e2lzQgM3i8IAQx31y2+UM5FguIR+/Rl5002DO8Ewy
mnVPz9SlGpy0RkX/OomVFfyREiYLyl6gIznQk7O5m2obhKoEO/FFPa0263nFx4ru
aPsaSzFxcAM0aZKf+uD/DB+/qUwVFiNMjBMGGJKbVBwUO2N14mmwphCW73lUGmII
tbzF/HoC7qJ/vPx9MjLO9lRKvJFW3ey8oJHvv5RGq8M4n8xw6xZVkOsXxrlGKg64
SR1gDRQN1CEH+HmsjuQZlkaMHO+J6u6t0f7UPn6hDsr0Ae8XHArGQApDE3eJDqXX
c4Hg7ntMCWTGNahiWsZsdQ6mDrGNBauXFWJ6CU4s5HNEvspinP6fZydn8K7U0swo
gq7vLpMS1cpwJhnLJxwBtMdK2q+xtU77hyzpAHS9OXPIXSLbfaqFuh83Ql7VwoQZ
NG1nJg3NMINwhjRpV+k4epYybAfPpOaRxfnIt3C3t0LtnmJasvmho/9b6Gbtb1rR
13VmZCgnLgPQ6H4vMHVyfyujCJ78ce1/xxhcIoeaipOLFWH9+XnrTplB+VQODyUc
alCyY1Of+xc7UFLZZ7aoanTWKsrvWmOluwkp2JfMz+Juim6v+bB/wODHOkPjJc0G
6ZEMrwsWoP6DYYZwgqP36gVEE+JsAvlAf/APznfyzH6H3qQ6p8EG7FrSTbwezaN+
WCWcvMojqNh8l5MqLG8VST5ZroOBdE0Ln5vpWlgYGvzYRd0Z+AZh7troY3EMquIi
dlvRuo0yxzhtrnSJIlJJEBSPNPJbf61FqJByz934O4o4YLCpOkPWgxCGB7Z6SKHU
JCmUDH+/5qoYcfbT6iokjsIxThMmv5h7hEC3sZgx/RJ3U+TJJmAXidowcJtlx3AP
cwLdgyfNs/UVuI6ogkiP5uUojoxefFpZP4URTOgAcTrMv1ZDSmXwwpSkGy6Wspy3
cBHDQglMz8rDVYQxMknNnAM2jmRcmV/LTUNYlDeObShzUHCcjgURYwhyjzo2Ms7w
REJ2MeqazwME5rq5ZWKON11eNqbNUM14KtaD4KZNgcKqmM2r4VJPoMo824/XnHHb
mlUPMXk77wIaOLiGGt6TPFai3SVg+d4m8z5XZD+qlZfJNv8WqdNjovDJkMGVqoGW
TdEgdiglj2Omby9fyRjm2/4MDczZmK/M1tksj5Psx8q7Gpq//jDhtfJjsLMeRyd1
GO7D8kCy3QcyziLGHwyL/mM9rDCAL6Tuni+POc2CWE+tlDNfnqB31ZpX52AMmFgj
cnblU/3hQ416FAVltXou69skGnp0mBHefzycOhLs2Q2RtwN3i2gp90OnIbknHUNY
v7lxbLMtvYvl+Ontjsv8kGjJaI1kPEI6GiDQ4/YkuM39wvIgJ9W3ZcHRnUMjzszu
fmB9aNbQKQpCQCnxHh+lOoDkSe4NdPC1TNgVuYiaIFf3iCOV8dhnF2JJq3Gr3kof
QYbrEiQVvDqqOEIRGQpcknqBZqCQW2CGAe1hw3vAzSOwZo5BR4xBHhEgbDlvv+Qq
hEVV3QteZW/Re5iWydt9TYVhi2YWr8OA3neJdUkkUuOqw2O8oTlkmoVKG70+F35X
bmvF1/EaHDbqnpgR8SE7HhMm3AxFjPUv1L4CPKvANpyWMGgsjFIXBhpWwVlxxQek
M1jy6KdqRlnu4h7KTIGHTzQ1o9e/n2khp6r+IZ8IhFtZKwkx0qsJoxYVk/VpKzXh
6iRdakNdIcMt74CI7PO2nCN23t0RZC9isD1vf18JeRcQ0Eie7sIE8QXqjJNapoPS
VX5/s3vLEWlI51x0l2/dDgpUz1xMee7H7tHaIMPQisigXy7EG7+IMJEt1X6PiNdU
t4KYBQP8QGB1cO2tj7uTTNUE7PkVt/IGMU3is8hpaeYshW1BssjcNgs5VL2ag22Q
h5IN7pR6Lp4eJj3uISkusaw6D+J+eTnHLn1tZfy/QdVCQkhNDFzOl//bcMoMsw0m
L8I2ImG22p00P2V9+VTdLDeSp/qCio6U5l3NSG2WunPoVJiFXn6xZ3d6BZSEtvv6
cjyDoUIQcY0Gc9lxpwKZXmz7OsWaPI6GZXBs+fgp6Ur3MKljsZgkmQnE7XoZZvHz
Bjrv542eW29SK5DZhu0yQlG/BoXvICTXuKCqq3mSVQKHK9BXUMYM+ffMOBJiu+lb
pwYjA8WY23rHKPQsyyb4D4Qhb28bb+dQOKQ/suu+nkrMWFx/OBUC2Mz5y+tCxqwf
kC37NlKPCHF1KtrssI261HSrCB5CM5pBg4QBApFgfk7EjXfYKi/gJ2g4gZR5cK7p
hbRjBpmIoZZcTNXRbG1flgistGeilltXfHEPps6K91my//ceOgG+XAoSLO9eLylx
DG4j4jkdnnsbTPB9s3AD7vKYLVkQoh0JY9BPkTCnX6sYH7mry09MNxag4OrQYbu5
I/2gWUC46sgYRgjOatJKBeW2PP4dC2Qt48jegJu5iCT++i5MMOG6/A92D20WdjiN
M+pZBkzPLkWX2M61H0hat56aZCRf2W9PoPF6Rgd8UhL8WqC/db/CivGAXfjVJwfS
LMJLs0fQYDIvlL5TVG8W837pcGSGqnM6aj7yLlY1UU1RwCnk7NFPEJiHZGde/SEu
gnr7G8cEwlLmIMsx5yQM/3LkPu5cOSPR1NUoFldzGv+okJzNgLHRQj983LhIhTw8
U6kAkik23+vpWJRH/DVGPlCE1XfQUi0ZDFGUniuwVaLX8jdeppFeXcKwJ52YmOjo
4QmclS99WOgqmKlp/ph+wpU/1A92ge88ZhWu+VWSFtrbWi87b+Zwaep47C6zQZ3F
AxciVqwJ9To+y4xOcdKaG8HMg0N+sPIx8Xl+RtURilC1qvoYeoTUkyxGkgsm6Fv/
iBT7xgsW30rnLnNmKa6kJzHxf1Az9Zvdk4yLOozTu7+NBj6SDKDqP7ilh+ZNDDAZ
cHPZFW7QaqYIBC9Q+3uPrxXAkX1JZ5rBH/EKSYzIob5tACJD6NYeWUhQhFQzXxqI
HdNlpyD0pJ2AyNwsSk3grYj2zYQKofynDIfVBHnzFKDSx4OvVUGG8kFWR7yZcXoA
OwS6IOAhtHIWpblqBb9p34CzlHy7f0ZwLtCorjQm9O/7B8Nf+R+zCYXFtGgfvNzk
RrUAkPAKpNhVvsHKFlc846XJmIcTsaMru9tZUor/P1vnRjdKRJLokEERmc31Utiv
aIqoRC9RwBUissKxz5DUwngJcoeG5fFhIQDGmS3psg7Wtj0FHihfq0t0m5Wu54XX
D09r9LbdkRVkA4YKMTDVtdGq5YzM+oJiQ0ombjtE4DxV3xt4XUk86PHXAEC1ZXSf
naBoYWYrq24Xa+Cr/rUgLSUSueDOxNpCmCUj7qgE6FK/klMuw9Y0s6Ucx4Jz48vk
5ck6+SoVQQHsIk4639ITdPnQ5tfj2awUI2hGoJ/VzwCAa2EXSxoDmiHQ/b3u2F3j
/lS9C1ChHBKqRgKXr2zdWdg95wz+eZOvkivO64mW/ZekAlMWydbYNR95w4M4GP2/
xIJt92fGu/Vv7k/XrWUMfuMYtk8rS7YPNAAZ0hL0IpHaOGw33CkgBmZ7iZl+7zZG
GqodKjhv+LYiQop2fEQoqFXpV//HjOMB+H71TFO8f2J4xOELu3AgWtA//LGhNOMB
i0uxdN//fCMrkmI5sViSHISSAETSAavq5/rVdm0mkTowasdsSuhaTdBqxz/Em3SF
sS91hyubObaqZR/KSNQMKoxmIiVVbGZVSf/uUmvWpyPueFhvJkKygdeFrcN1vyKq
gBgB6nrlf+r1Fh7FU0AA0WK5Hchwi/q1dT6JFZ7tOoNCgKB46OAXfLFSZKuBuPO6
K7p9edl5tEjXmE9umQNWEmKGwPXCThMSNVzrLiTDkBaCM/OU/idhpBiTvdkP/zh4
Fk1vqZigYOGe0RdYrUnbrD7p4S630UsK34qtMrVpY+V62yn77T9i5e36u1+biMPB
oDDnpbtklgSWbyiJKQG8IRKIV2PWaZTIpx24iL3Us/uv1rHhZULwJixdiEKnZftU
owSsRzWHLvl/YRwK6G8hf2UMgMtu7xAmBrbnEtH50qzXPRpB5qlDeQRj6V6hYOT1
PulkzHiI55wuRBNh+u2fnQ012Hw9A4dATdjy+KXcgokN3LNvwdlgF7kP8raAJKEz
WwkiIOODfC5nYko1zGYyYftlD66sdgQIS1VeMey+qxgUY42wYjhuUayVLvZ/lxw6
Flm9FkxzeNfmUFMsZZ4++Gx3ZWBom0IQ0h5+8MFe8ryhTVgCGfLt+1Sdas9j4Fvr
Sl3VqWLT0I3Jm4coIcGMOLrlppEd8FsHLNeHkBKBRyQraM3lzbitRMgI6D3swDQI
7YwjrP/rIv1buj6BfTATZUumr4mxi8cP9B5/7MiazZE6Q7mEqNzSBoHdCC22CLaC
lB8nf/uzHhg1Blqnv+/dI48zp3O+wRXOV/n4STyxgth5g+pdqUaS3uHa7bAj8UYk
vnOqK412/pqnmbG3hm5O8nO+1nA4WAPXQ0j7pCT1CrAx7ruARhEa5mZ8PMaRzJsE
4Un5qKRsJRyPWVLPtdW0NX8B7lT+P0Fj2fzpNSTOaku83dnEkgvOxd0wU5SHleNT
kc1TN55K4ouk9c4noIjazBxxjDx5mikem8EkzLEsWOPFwaIErtfQEZ95ZX4xPipJ
IyPNurvtVgTts3a376cAvO5wVrDHDZJOMPB5AV2iJ+RUp389N7gk5aKB9FycuKyx
OpVua7J0nPk+gElmxJlcbaRzy0kiEPEvNp+yj1BxF9oaSBOWZxPzmwlUKRvUMAo+
oVOPrCXZ4bNZu+Sy58XT+0KbQZwwJmwE2DXThglfxandyFwtv6baamlztD5pGuKV
2fv0k+QXODERcAI7BWe1o2JlZGxHsG34ekJmCZeYThmF+UY/K0saEYkyiW8lxYVp
aEFgtqobLbIv2Uj7Vv6ZQ3p5ME+AM5ZnLPAvd4H0wlP29Y0yiVseBd4DwRnoL8uc
0AjTGdwszRCGRmail/jwVzfSO7X67jjqYe031jIsjQUsRAQKvqUjRyCSEbdXDODq
owfmmFluaIoCrVuhJXGC9/F1UHikcgdzxtHkwttXgu5r3WnhtGRFKkc9cJmMBC9L
f30NRk58iaqomqAJd22PXIt7xhyKeW4TkASjluP76MWrGgrwpCjqrA6mgLwKxJtn
e7EkKZ/57b4HEe03faqSSlvU/+HfpFf2noYVHCOKegKWau9OZQtz/TNEJBi4Ln3a
FGfounXz3EwyEjc5BpgLqBwp4fwmVwqONhEJ4Ay+lFJQ/YXtZk+197VJgSQdpemY
vKfS8VXPWUebdxd7qRebqFnaNJaYFuiT137hRf7b2ch2ZzYtwnlGulG7T8fCPnzI
4lEPaFKh35JDNLtc3wyGVK6vFgOhMKsebIsYp2vkMGwTRUW2A/pbgZ7pcWhR+7MX
i5EQ3pqwWaRzqRqN6R+oWJu/snXqg+rSUsk8myLMr7Qz6dWEpMhKnyRjxwHI89HX
nuWcpoVCoxEwnRwKYk+9UOvU1TAccZAUA7KEhb7u3Jma56WKzxsXagT8HQHgO/vg
yzOa1tY0oZrGsMh3mUMFV+NxnaI5mj7dKhBbZk0iNdRgN3pEzuu665t5PeR5s2Xb
9mjHyaZD6OTpLuimhbKPCajBDE9wH1ctgjrXftQcIYeh7dIkSNne+2E8pAd4+Ial
NWa7RuszbnYrmmSltKScxmYaZMRDcsIm01BaYGQLSxMUt8B85fIP1GVWukqlm63M
tdKYPJOAEtJZg4wVIWJRUOjpi1T12X+gW3ZlwXsoArwrFC26l1aadgk5s/V5mZs3
FXcKJmcg+qQRYnm8unFOY8DVb7esH2tCxvufSpArDdyV+BXTMqbftYuSr+pGpxm2
mn/fG7WoTENLek7t4notRUOSLtLSZCeul+OFvvCBnNuU0E+1JzVijTsd/umuRcvZ
/qbv59gDZOoiu6uudiW4kkqqN/ywmmT614Hx79fGE+uDCnGVzI0TLGxWLBG2SRuG
jnZ05i4NnbEtVWZ6PeTth7mivOzC5cvejo5f43n4MZ1uJCJ9Igy8Vit/60JJ2VTP
xhiUEKRr4h6WjhoMARDepIspAa+j+b4TFQAjCjNsCWStGP50GVBAs7hTvKiiT80S
V2Y06fPFXkesDUjry7g1yMc/bEpGBL1T2l1lLlzAVAunB8pNBF9pWN0mx8qEBx+3
7Kfs4yqvMLqolQmGP3K7zcOTyecgb7S5tHBNSf9ogkzEATO6gC4blGU3uO7AR+R5
iMTOT2YjGcwcQHuE0ZRMvm6BztX1WvsTQnlC0T79UHN/nW0+r5UqJ8eay7GDjwNV
+pAsBu9wM4KjCYUy4RTtuyjA/sBLQksruMPHh7zxSH/phusPG6Tczq+m7SN2AKV4
agagQDdNlKk+lXI4th4nz8jTyCN1dMlN9WkaFhn4EdYPF55GR41OBJ8V8rMVNAtJ
+7zitdNrT4K9GepIhvVnB0aB0iFVe/cNb1YdmRzVz/H0B7ctj3CrLwj9sShFnhEh
69r0rEnzAldArGC8vtLgW2Fg2Fc6nXgC6IQqzVtE052OK7WsD8FjgBwFblHQN06c
H7m+WH1h1VHiU8xpNq7kKZ23i0HeE3PZnmJS+GQJJlkf4jZ1cX3G4Cn+BhI07RBl
0RwOfVZSyE/ZaFF/wqwAT2x5hU8tJwcD79RBkLl3Q3t+9ghNwGIRljLk4DGqOZKL
XIba8Eo/223BoHwoMySD9X4SLx/+y7F8BkhiignFfENslOPyhICH18znBST19tJs
JNkGJNDjm3kA5MGuf16rAKApW8DSapbPVIgm4Y/7PpeUKQ8aDHfySCJRFwYsa43L
0MLxRZCLzU6yF0/RvpJwlf1wxuNKoO51cHfeF8gkKNU4cry5gVR032AQGaYGBFyn
6eA1W4dF1CCc+FHqvYqOO2V+ORAnudAefc+BAN0+dmxyCwKMdEppjPD9S5559tc+
+pxgqYsMyIYPaS74TzmD1zA4hKkrLy8agsmSzCOjNFubdLJime5wYIQhi+cyB13O
nrsAFKYJtF/8P/0Z/TNQPHw2ssk0aOTAyT1pNSXMAF0NZuY0IE9NPfowQmKI/fIG
uZwx5WPBPxNaqrBLHvF53iBG+tDhPVBPeXfQgKaZwzhKYFq+UQMfTOLYVbyI3QTM
+vxd1h25hgbFa0D52EkgwstQ2Xn02Osl2sFZAWiRqrA6jUtcWZy0qarJQOBw3wvz
Kr11NmIXgOhW1X7VWSApmFrxnu9G8ToUn1q+jAavYLyKYM7OdVIsioFAU+BBbsPl
SQRqI3L36rj7f4BhHKApvwAWQg5AvWQ2D/OE+WAW95WyWMb92PVoDgyGN34HYzmr
8+grHEunuOTbjTs6Eem3nMoti5Zu8yngPt30QAtXia+5//B6IJonBUojWx897G7W
AzK9TcUWZyjfKgzHpvgV8zbrVgNGR45PG/dJMEUYTmwKtOTWER/pF/x+nDjowryh
1fCtuSuUQjjZS1WW0GuUIf/cIIMvFLC9xlTP1xfcAy4E0nzee9HIXEiHOfoay7kl
q3hiAcHkUkN+PmxqYig0yxnOmGmQMuacpYFcbsGFq6DFoX5Gb3G2SS/yehh4P/8u
dcCVyQxXCC63mgdzSPfU60hkaGLmSZaZbl+ahDADIedmkjeXw3cb+7CBiC8iH+Ev
LVtWb+WPVAFjnYK/7llVzUrXEctfeJI+lRtpi3GkI2IdbwCQ4wAaHiyEh0ug8m2B
4UtGBq9kF8qDhGD65wCi8a1LKaUsdLFSMNAE/QXYANe/iwpI39Jb2uQean5AYHnw
443c8grnT+l7+bt0Y90db6fixy0QmDqxNtveDM5902cfaTMcFqiVkUajLMIrk/M1
S5NQULAMawR4Zz76EItqKhqK+pfQcpN4CLR+/HgZlLRVK9Av7fZRbnb4fzISDFOO
o8Jeet7vzY5UfdIwlQ55dvtvI2IAaiobo58ZeFTxDHAGmUXl3p8AGKKmXey2N5kQ
AkgOat38hhVJ4B8vdUC2DATG6QcGvMkjhaQcmNHYzQ6Zf7MpZNh2i3JFhgPY2JMc
nwhM2PccW/7RNNBolw0autLPxIVsrxOAYSQL0zcLSa1Uoh8w2YGVfXgbgkM2TALS
znHCh/nbS75+L9gHGAgJYEcMSLTeEvo1396zDv86CObwic6dxe44iIpMheAf2qdP
2k4dYPQr+AgNRtLnlLNe+93Y1MW/DzUDIpOO/FlOlLxurZZhj7oGQk0HpmhA2zGS
IwQkK6eKFqTf9SVQd43VL3c4xoqfPWEJRnHH7ZXDRfEDj7Tu530KZgeVqbOCY/tx
53ZEuGZW0Bb2m64IPtcKCw1h6xZjn3F8XHlw4QrkuZs/0NthP04f+4vOrGMJRm0b
w9AgGyswFA6JbfQiRa/QpCUyK0eJcdtQqtsWz7hRFf2/bTdvMtAgtYTT8yN5aQEp
DpvwDprdYpgR7Y12YVipZN+nZWuncUM+1nItnfDis4Z1YGl1N3z2U+b9zjz9Zn63
gEip5NRwPaBvgVbonk/gpS/O6VKkbtjbL4lDxZYtjLwWN4xAXqIRUi+PNdI7MZ16
aqEU+zhzJHb0YpjNKcrPK8y6IdFKanEInBleBX/InxOXsWC9kcYn3DzpoL0NLeHK
G4cJkNziIBQltWIqDRaqiet6zY3OnK00GaXD+8GFWB18obi3Vl2ucbAGcYAwx0kM
wLW9hE4WaDV3ZZV7MNOqM+1Y1h5xO8XPcPTwsh6hDdB35HRpCby1jTKewv61XkRt
CwT/YUs9mD0p0LFo0uGNkbhStk3WJwDXFUsa81JOQD5A05E9iZWjZWoOb18ZS5U+
KM4RbL0l9xwhZ21VfSuePtvBX2pJHK5CYTfooKZq8LAYNUYU6OWZc9W6pECLLpZg
ezMkuhCD7VCSQ6Henfl0OQ2jNQDZ8w+YSDOKnlxrhPztSzS/mXOCDDMxTaFN3qbH
wxC5BVMcl8Kk87UTZdsq5JCcrwbOBjclVntvHRq7QBJjrLtQPLx1SBHaXlpiv7+8
Ua/jeK1swn8bIUoz+oFh4bbGHECEUajSKKDAvfJrzNpNCZZZm0QhyaR9yEemOB4R
2/Wmqyb/m6rNWO18CFIyQXcXMYFDtEVaKseFV4UcWxmfMiu4h4G2L/tZ8cWHl6mh
yvVCX6jXnrz1zWAdpydURWHnrEEnykSeecUPUo6xZrCfd2KWyryzde+76jSvF2Tn
mcjRUJdLQjmqJ92jCyPvG18XxwKWmUUYZsRstN/8O+WiV/4Y2dQDjn837eodiwJF
EN6lT1SgvQHmPsuSoMmXyYHVnuikaSta0Am3qhBB/0xreYXqdVnZSGf74crPzlQI
enhC9fKFVSIvCZg7x5+Xswq0IOaQRnquTdeCEdNPrbk3y3McYzgkcUO/Vl7CaFpj
0zBmjFrYZWfbiweMZU1MR/gGlXMQr6xrq/s6TQx4m+ycGsDaGIhx0NNGE/9ODXnD
6mufmoVR13QPyhz3ibAg5ER2vIiiRpkXES3slhr2ranS4WI3uMa9HWkW2dkP3BaE
xnIul7N6RBBCghYKDHQZppUJZ9X1QQglHAGjmh1hS05lf02AQv30ULxIw4gIF/RP
KwOTot87ObX2uRfXD4mOf+CBnTK0NVcxHO9kgnBIQL31jH5yE1qu6CWI4Pqa5les
4zvMeWb1ZcKCp/bazqpGs97Xu/A00XFQzSRRbn9+0yeO6NodPGgBK/7gQ6uKz/xo
nEOWChAJlHomPFvCvtMJyBzxJpvm2a1E0/S1z80yUsd2WIUyn5njRq6qGgfqYh9t
CZ6cDgmzR1lTmQeQgzq3mYncajE9D3ihcJuDqtaQOeis4APUkamabu6WjyPiXmos
4AKZ0q3/6isc0HY3I8dysqvzK3Ivsff9fFdbLwKBLtc2V202uSjfjh9SG0DrywqR
nOXy7yTeSsLWdPRZgbdvfBRiTqVEtRdDG3EJppm03vDKgHg6PGCNPCpQqty5baBp
bPgbi1kSEYjkC3dtyZIylJ4+PNeucC3bsq3b/SsUy4bCNIcG1zp4c6YNwLmdyxzR
dtWbd0vooWPnkaMW+RXtH+zYBERDvdRrSMzsfGlhRIOiIYayoi/EaHHP2EAuVeb0
ReFCfbz6y5AO3UXd2yztLaWTTSz3lEWk2tDqhaNPEKvovYjkJRN6X5SHBCR37paT
c0VL7jXXtNFAZ+kI0s01Z+PbEzO/ucG/TlNxukmrQ60Zts//UMWoVAeKG4rSwfEP
PfW/nAatc0DpFQBPwvAFee1mzh5VjDgfWzDx+712lOsF3RRjcZwt80L2stP6BlGJ
xqhRInI9CvqbmPXhLTzcEmqmCiZYkPO5/JmB7Bf2G8Ko06CmSZMI+NRXZfLf+mNQ
oDLSU3CUZgvEBAdLziXlW1KvX5Jkurh87n+Uj/i7D+9Gru8d4IsMt5YBK3IMMcdd
ybO4a5drqzIl5/I0jzDxgVogWHKA6Fu7X4xQfvVVLgSxVj9F03aNidQelm2DrYT8
bJAzuNffcI6TXgoapWH/+qoigC8c41jWMcIYIh1V7wWtL399f2u8kTkrZcD3Nsw9
5DAB96J3xiM4taPDn4cVFDTXHOT850KsGjdkZCw5bxkh84gnh/NWc8vYS/OnWmbI
nFi/tUVl4Ym9G8BiErRS4XOVa3VPIwCVKgLngUEGzGeCoB/8Dr5A+nQEOARCDjEs
imnfyiu4k9frJDlnextH6q+GgcixjRUoQQc3uyplNwLfaVg5AlaNHOycX/XZgE36
5SY/J+5Yh9SMjWKJXEPys2JrvKQUZcoERH8UiJaafp1GagzqYWCHIXN2CJkKWKdn
pq2IsNXa6PYIEVySSRX0k4zoYiJ/UYLe1imL8vaK+AZ55B2TfcnLi+0emOsySYfG
us+tlnLfyHsyZxOinYCsQEDBvGRfm/unFMftk4VP6uU+8M67GrhwSxht/nM+iFT/
yKUpcvJtZLpI35nuxQ51mQ7wuEvvdetXLCJgr7ujEN1Y0luQsd4uzQk4uR9qcPT2
j7vcFS6sOB/rYBsFEb2bT8+Upx+TZN3EwN2z/25F2hyc9brXAvfd/PqcWPcpnld0
RuXHGOxe6p/CnzQ9VQJFf01iCXIBxII51FMN47G6sDBFlZGfFj6wdc/Of+d4YP2K
SXowrn+Qt5dNNEGueBFrEQLmp8aiVPUKl20XFjQa3UAD14nBJEarMItfR1oeWk+2
lQbhcB3MlErLC7mAXjBtrPCT4uV4/K0VObttXj29FS5XxwRndxAF0t/yCgthpHxN
1uXjtqR3yWdxuPgWaGvGbsHqLoprdaM9/2UHOpTdbb1aAwzAFTG+jss8NWPXrequ
vGGV6Z+jBuklLa4oLcjLRkINLZUmr2jk/MRWSkK+0cMioVC7bh9SB3xLZyf3/+b/
Rzt7A7wfl1R+af7/eDBugnRTjj0Ui/ZPdwmXhoqsYliy/W9YGtOK1QMV/jXRagqo
XPtYOZlMlli6Y/g3MOSqt9PF5wbPXYZqewRRpRMPUKN5hNATSA/p+0046tpKoSF/
VVEnAD++TMCd2YxpxEs7nq5poDR7rZKU2FKtKYsavsaFXNGSLphwzMBBaZXMEAic
p6YEO+ZFidNh3r+ezZTHYoaXEckakA3ntcirCt/OF29gKZ7zI4CORxwQy7osuOVJ
zek/FJo7/IS3FX1Com6iJVBnuScaeHXwOJuJzqCN2Jj9oE2CkRNhDj3602wRJ3mK
N2HWhCdxHJzE25EUNGjqM2B8YhS5ajO2Bu4S7tFtHDhhR99ADB0SjWXsFpUHLWsG
OkY2TN87dIwBmgMD0yqawBtPFsKu/pr8Aj0FiMpwwht/2olohbebymgkcwMPd7q4
kKzTK3bWZLlObm3RYdIYX+3USHjpT5YGlL4xAqi8u8aRYKKcfOzYEMWrOtcXwWac
F276t+SKcn732NrJ09pJzGfwG0OzW17h+hh/Wr2RqXTEOLm07FSROhauyEn693wa
5iQbOS+KjJPXWAwe9Ei9jUmhIqKJ/KV9f/T/7ETUyy7tYs5gptbQCOQrRZXIoFQW
ssBlk6m1E1N2Mjsw1svkTxTxpwvu+w7hLK8Jtb/qby2FNSUfS05kAikIaKgQUjgS
CTtbKJ/x6rWpSJb69SBLxZ43rtJbOgXYZGPqqH+xjepR1p03k2z3RziWScXWUBGg
ksx/3nufeR26RBqIMFCH7f7+6v/z++RXmJU4LV7nN3Vy5lb57KFZlsQGDkhGYfXu
nYeDYT101BCFyY5D8Spe8bZ/L9us5wzKUeLsK5r7dxOoVoEb/xqHOh/6Q83Liw/6
zWUw9oqetKr6kGIIJxHXf5Q20BIGS5CvNUErHNauhtunzlVHdSwgwvB3WW75+VLd
MdeJ9PLu8HcuerqqsFjdjiZNj3B0nDq/Q00+MkpLPpW1KKV2AxeYFEgD8MX/p50a
icHLhzAoNaxMeYk3T/CFyw/YX9apOc0AseEBcOaxMx90vNppC35PCOf9+RDlf/y5
MoF8Zl5nIGkyK+Rn1JDECBBumv/LipOXdWIetTqFt777gEa//AaC93zMNFp4xjjN
PhGgVmOaH5G2LorpXPi4sp/fyai0VflfvEc4alJ+KWIYkWy6MNjyAb02uqJ1o5qo
UE7jKW1tWn1Kyl0lx2j9sc/XH3KYExvv/iMyFWxdujX8D61rnXKqeGnEd5A4NP7t
K7ecfoaiZHU7ldgngOUpJ5oQkDvUOEwpd8hCe6KY3jEDygRIMbvZBXcyyH9/QP2f
NbsAGnN2z7Veqt4dU6WOjGGcIJWFdqXdy3H1cpRchGSLhzs8qbIfbh1LJTPD4oM4
qYY2Ya6dG5WWSqGFa0SQhoAWPBxhmEs1oxeiuIhU1Xejmy07/no7DaVL+UaDUplN
GkqiDV3i9PonZWOKicnjROLsT57WEPi4/inuyXVshnWGUHZNUk3hC1SYy2dHuFem
cvGv7/SawG3UdSN/GtNJnOPKHwC2kJ8cy/7n8lCEnL9VKUSEVZfG0TPiSZ7z2DRh
93AwC2LhXTqwkWmMdLHA7u9rfJTWtv4AkpOrhnkao2cyiAYUiqMdpj8sKZYo7usY
aLn8nEwRrAOz9gst6qcyRBKcTYjvWty4di+k+1EdAZd5yHt4Ya16C5cjoAv5w2z3
q+4Y2t8YZq+3zAwRjl15+vCB8t4VbDNiWpjqDeuVXQKEm0bVOgg/qTEJoXFutE4e
P2ZWMg1sxLhJKDhbNhhhXOmzhJ8+WKRrXuZNoShEo6ndsXtdgqxXwCMzRnveWK1c
GxaEvMN+RAVWs2Vq+rEFDZLnrHnYmrVZpAHSpfb/zNT1YaOPsz+BvPMeX3QaFwzO
jj8XTCbaCJoQEmUQ3ob/8MiUZpQ8UphJ2jZn12M62dwlpxdjfGK5OQc5kduuQ2m/
vAoAcHU27v/bfnkS2vaDPEWuwrqRHgX3kh7qYNV6CHaPa4CpQvqsXOKSY7ZDx/fJ
E8uI0hF+DxT77y0BdgsD4uWAYB7sNjPpBHFQ0NBUmejNFV3hCMlIgwpd4SIJIEV9
EKmjw9/4vxdzSf74chX8LRrySnrvqqllZUEU0k7uL+fBtedG73q8CvAu5pF1SP5F
5sX92xez3F4yD7WvkYUm/Ksd7M1xdnwBh4iR3AZRAQZcOn7neevfLIP4S/xFaDOv
WJraG5hSiTTdqv4pFPzc7PNSImdlUV7qD9y06pJ6R1qimgfD3aMUYSD4HAfbAdXv
oPVga62fe3DGnPElcKBtMb0ZNi3dO4Bwv9BrTrIutIss889KGTFLgsGlwgd6CMGi
NkCGG58ic07PWOYr/t0dP3Jcp+sy0mYGsAP2sWMEZ3sqdxZ6GVj6k2aFTgz24nao
P8xaZA08l5foDLPgnATGa9vf7KO0cjW2yuaG9JsysCKwkrzXwiQ/0j3ZUD0YsC4u
cI7LKztpSs5LGg+r2Bwv/jT38vumirpVTSXhR3cM+VLXX3TCHCIfZvPdzXNpC3ft
gt7M9UY1v++on3cAJ+YrGf/bfQbtRpVcDbzSReRKxajViEoA3Ab0dVt1QnStLPL1
kqQOs5zB0gJogu1vlHthKbQD3DOPvxjsga8DKd9BIS3x8W+U7QdQTHliobs/YyyT
KrqEZ9nPBO2kQNaQgsGOkTxsH8m8RK75NSZOCf6flJANsZRbKYPdSX3CYeQX7uJ3
UPaZ3XlnkOBoeoSGW0kaJxCYnVvsx+MmCegt3zeyzQGci83yeSYb65rMxEQKlzuF
qGgtQxBRz4KOZ+5aSSD+Swb4b8fwN5oWimzqxOOL8UArYfYeOTxNsrH9cxLICmdW
TVmFCjdCecGxu4yFutBHyjvBQz70bdKiWC9KqAHNPZ7cZSpmyAxgbucdMBCvB5Px
c9ZMOxN0UtKXJVKN2tD6l0OyZQfAvbxSZdcGGOqHHqx7ScYk9Z2KA0kbldTzyO95
aKMjSf6/NOOF6bg+qtb5ddnYdzZjPLiwMjq9NWmGwgApK3iyvNLIyIYreXropkZy
e4rZcchUu8sWNQIXB38xiHbEA2HJQNDYxnQf51LHSj+SCePn5Z6iNZbE2WfFqTNt
u75qsEW8LkA8HHxP8bzINmwOmy0y/329/yBfRLGBhkj3drVOEmFCpRVqUtscQKSQ
W31hyO0B720uOPkW3Ok1KeI//Hy+PU13l+aljyU4eXXA7laN0XeW+F+WJYoLC1xA
3SpIcN0qZq6OlkdQ4vdpamcUz17mQtWyn+lOhIxeroCuuJpaG6ARwjOhyOWGkizw
bxPBJ49H+0q+sFFlAuIwW+qf6Bm6JLEZRthtQcjvsCYhPDGO8Xwka0frAgv0KzeI
koBKNrgvyM6UWdd4l56EXttzsPtgPIHnsIdbw8F/e2gjipitfzMAiizqXUjblQjx
ZYhKKq7IwQPx/HKLwIfDo64X+3mxQ9BkvsrYD6UKoCIL39g5gv07tMCVL68MxGEC
l6Eun0D9kf0+EdS1by7MT/PGxLc+J7+HKQpSAHRVBzdo4/jhwg5BDJW5PmiGpsPu
fz2kDtPqSTQUwQ6cE3565i+ECMTXXIPeRXpZzp08uqeSvNixL87UJI5q/JOtP+IA
1ZcyOmEFTBVnva4/2KQE5VLk1M88uYbtzNn1zw1XwaBaImKtW+xHSETqIfOC2JEE
rnFEs9Nseay0wQBgumpA2eqBR2dauzV5GmcDF09+King5LUdYlXjt3LaFMgPqkt5
Qgv9EMHusKVSVWRwjVJolvqe7oCi5nmk1UDX3+UrnQBhKsv1b6NeypN17BPPRiKf
3/FJ/NEKp7niabH2D0/rKMaOU0YUAKADK65b49dcYo5qBxP5/jrN/HsaflSR/CdV
5aAWsd64NeRVIXeLejwus7CqeXlMJXPNmkpkD0wnumTWSBf6XrBYPVE4Een5COFo
2DK5z3bQar8OV3OPYYYFdMsLZwMtP4pFIGPnVcgEwaV/rHTzdOfvbL0ZEjNHk9Qs
Kx/kaUB2/+bq/06/tK+rTvfTqpc8hK4JuT4T38ogu8bGYqHMrLEPLRcaWSd72nzN
NiuGaQOJyA/nsfM9W1qOlO2/orRQUxDySdd2/Wuh3JrEu76TE1dsgDvAIwIPUgt0
YoUlLpsT16QtQGAJ/dTGAQBB9hlK4coJK24ubcLrykdLZp8cSFMXnlxae/OeqxzL
msCkDjl94mSVisM/PkLJjLZyl4B7kZvekhpeOUW2rYg3xUXDAoKaterrRG9H3t5V
O7cPfY3bnytKcQY2pJ1J8vQarcQ4R/AAgGKv5lM6bzwgZF2ETxTLr/jLd/3dcIVb
gm1/BsKfqKqbubVhOnhcuFiSQTMHXkbd9/EcmJK2vf4FAgy71dnYdF5hKhlOtaQt
FAbXVEL2FR+/cyWjg6z2vPJesXkvYixkbjklDONifrBrwH7OPYY3TcZcm5JAPkrd
M0+KNwOmsn2OVl65KdSee1EsNEKxEniZaIumzfaR8cji8fuuKAQfXa5+6UpdVQ05
Yua6gQwGSSXCSe88o/O/3AHDo+uQUWj7ezemJcqLYFUW+Nldhqn+WoBj/QPAZG48
F2nj93qfgSGbjznH9O8X1jM89ABdVmqrsnMGZ6cQg3Q4+FWH1Asj1QG3IXoxispp
bAg9RLErGaf1U0XfWmww4yj7LaTZgMTdnP55u0IP74wYBg7OucTa3ViOoy3Ghd3+
0rLxJdRjCYWLipawpcIkJatubcN0krOVmhM6J5dts0FZFpSNVHhBI4G/rpxaOE3x
39e917exTMDBP1CHX9FA/tn+NId5Tp6XHpILgb4JMSdUTdGIhSIz+wwHikRh4Q3E
/fDJVC0ebGZpnMVKoWVcwg+ntZZfK0jLrfn0iLWoonk+I6vrFQ4m2DooK1EAD1S1
33PyG9i+YlpOoMrppGv+2G/+q+jOHK2+0IdsO8XjHreHV+97NvpzG+cSUnIyg5kS
ucX3d5dDaVspz/xxqwNSb2vbjqV3xCONbgl9uEk4mn/GyZALPew/39TjbGXRyBD9
uLZg++1pdJ/7UqM0F0VPgaK7J9s7tNxa2e1DMQGyyCkfmA77HDgQgG+KaO7S3zF5
f8hUvgE5V7p2c6Q656I9jIZ4WzXXXmLigbYDNut5xn7+JMPMCHT+I2Oj2GUMuYo6
0oOEAx8BfHQlh72gtnUkEdqgCH9PPJCRz0niKUh9RoBbzx6vaxHI7anB0ZRFA2NY
8eS8Qal7fqqsyh8BXoUO9nVeD91lQla2uVz3BaCM5x9qDGFUoIV9hOc3/jQf0Tbo
5WYEtv95kg7pamqGwNOEJhX99EBIitjpJsQGPt+i2TA7PZS32pXYH5nOZQ1m4I0Q
IaEpSiR7jaDAhB6Q/2jZlQ1MB/Go8gfpqRzAI4VE3BD+DxlWU+KRTZP/i93TioyL
rD8P2KMz38Y2ZHzWWU4uu5DcL0yc0j3uRjaC6yos5UH3Q+u+vOYCC14pDRO+jphb
LLG+ujVDOkppBvPThGK4dq0+vkFZTDYSlkLLwhp+DFwvsXPYNLheIIWV6UizRhAl
+CDVy5+fwAillvtxWZV7oCl5RXTDsay5w/tmUsRIzEYABJaoRloszvAGkilLWYEh
lseIKpVFVx79wMAPiWfrXtatusO9IWX4QiVj5jqjWXGzBcb2YRdDzMukKbMZC8+L
n6G7kRYwTVmFuA6yog/qYNWHWNvKY0FpEhcU0d1yVcDQNgMMtAIXeTRMjgjZqxcV
gpbQokS9W/ugjdorWrwbWp4WLz2Ci52YNOhti1W+tGXP0FF2lLxr9q5Rck40kW7X
2CE7E9Vpwp0DOCCVjagu09OaCc+HRNDzg1zewD7oyB2T8kfiV99yaxJA84Dt97AB
PV4QD9fNRZMJGSONjoRnxiQCyR/FpnZMarbuABSJ1aYub7clMXaRl1vj890feJMq
uXToYALun9peyBDSh4JJnSRdexOxrLLXN1i9vA2pVTdOj0bZPebjyg+BQwlmgANS
r0u1w9sXVghON0o6yYca9OJ7y2bSMIUm8JPu7qs8rU4J0cTpUDgo2Lr1m+TsqwLU
x41WrHo1PFnCobaYrY55pTr0UgqSJFP7ZlmOe2H+lo2LGtl9K7x/8QWMg2Yyi9Oz
CXxtbtXx0lZnu+x6XMCtodRI9xvxqa+HUgM16QbX9wXrjjLfse0iI8CZ1pGBNJfY
wmQi9KUIgGvQsdxr5J2bwmkIql2r7iExHdsZ3I7uZihyLgbFoaeMVL/AAsek3SiB
bse+rnS62mBVE2IyV3pTawi+0KrVyYx8uQesAptcJF+kIp7hCiLUVPFJYVy4SiKk
TraMUuc3Mn/eyT1alGYPIYAlTBGbcelm7W/Mt8TRgihxVorKG5ZeMoPPPRvTYfgU
n5JLsshz4lT+1VrfnZPZlFLXTOG6W0x8AUPRCtD3EMNdyKfpiUM6MPrg8s7l+Dgj
QebtDRNIuqTG0D/XpXDpzXJuKxRm4tYHH1KSg7+SzroU7S1Z8lEzKCjtSBj9Md40
US1TrAw9s1qtEuA4SxpyNGyQ4lNfwZP09B+SSBaEWhShMQ6thFKFSSKtrQgkuO4u
7ic+hzvyD0Ual3LnJoxrgPSUYqhm3oGLyz4HHf9kncK9F7n5Q3Mn4li9RNx4+gMu
J5oNycFiEXHcY+M63XWADtOyBjRAN1itz0C6tkVpEGaII17BKhl/jze5s/zSEUrC
iDYAwX/YMGQO0w5m3DDK/cmXSbXMb52Chu3w+SZCDyAzuNXugUOxIM1OHFqhwpXA
xaoGERTzs7Gds+rQbgCtSnbcUMV3IQ9HhwE1wzlq6LVO+ym69aqrn8WA0FUfJpTY
RhV5dcrGPY5/ZfhvHmTV99Led9KIbWfj/bp8kK9AG8G1CUIV8HCXDZ/fvdRXpZ+2
8HTJyPDChvan6s1atmS3e38Hk40a6foqMJI9d74wFNWB4JiZ6VdjCZoNi5YY8dY6
KP7e001A/gFq6rGLWKpdSxpF81wTD/4OB+e25FAubfNNJQh60uZwFFPBDVuo9tg/
vwW23v1F2RAXcdQ0uxj5/Ofm0DCwBFypSN0/s8Y6G317q6wiCIcId+aYDetoxaYl
q8Csh4h/pFeY3L0whnTT3VhpLuddbLAxjo4jwKSOw1+ptq8pJ2FQSHHgnca4ACx1
ai9+7KIcx/O8pBsRCTJJxXHcfvAPBgCfWY4pRmSIHDpTA6tC7mvgS80nhxfIe+jD
Ch68d9VYkjYQiPfeh4UW0JUe5yqACOF4a56O1tAVJOPSU00ySOeLLIgrYobICFnG
ZhYjVClL/8XKbC93q8O+xIMT3VKh7sve2iy2FqGj/rDwumTa6zle0iHCCDKLp9HQ
diNK1gS9KhqfmP42xsVkv1qi8HLydEtkvUta5USrJ44zEU4yUsPeTZbjYZP0po/h
mk7w0Ugr3IMJzVEqy3Y4+fpErAgb/o7LzuGjiucpor4G9THMWtYzcbWKmc8oKqem
GqaGcPAPHsgA+gXrytOtCLJuVKcsr1kZMrlJ1R7oxlx1VwI0u/j9U4QjCK2Wjfr4
REK7Eyc/y48ADVulmE7BpHRNUoLJwjpSPBS/rBteCXFuYQrF4MMcZFHLmeKR1IIS
IfGLVlQrwi52OFNDIsiHSVj1zDUAlWzNoMiod7A6GC25aAt+UUXRx5W9GK9WcHOi
V+/HZaBLCNFmMIuAeizVbgrBjvZrfMc/t18WvORpFV6A1ZZNOnU+YHish2thE2N7
wSFZmxiBlDpmli4lifLJxbEtQZQmbLUvV25vS8Nd1tOzXU6g++Iir5QcnzvaYZWY
REr21c2o3uVRFHOEwJ5lahbON9iMggpkTrOJdxiVs0NLq6Ytu0J0JfHJwUQI7l5e
PWrx9X9lQbG5cdwXG9sx2rmKb0X7PCphjjmDjng43d/vyVg6bQV5ihJV8/ywehz7
88oSGeqAPmOSm7dSpR4MAjxllJX4QpIUpEu1lLiYnQuAkA1JAxNSjGOC1z4wKdUl
V9i9EqNElQeYDFvoy2NBO7ci7kW3LMU/CiNX4f8N2UX1zNz2YSU/iShTAhnBPr6T
3IO7KLuESDZk2uxJrDktNgpxWTQfbO6gNu61ys2vG9j5zi3p3sy4XVXKHcwyKmo8
QRrMUophc9C0w5PIMJLun+3un39CO7YcxmCQJ9FndG8LJAYc2JhLEDgVi2U+/iWZ
q/qSkVpOSOUnJJAYFfC6m/cRU229u97Y85UPltn1f6F4f6Yau1WCsNIIjvTemFsO
xDqa/uk/hnuHq45effxLmtynP4oWq0a5ZiU7l/KixWVBWi9VUtOlPmN6iQ93flkM
vgRa1Vy0dpGpK5No+60lzbJc+1Zw1npSqR4GH/STIqhNvB/w3QaDaU7JCwCWBEj8
E7bONiSiihnNjrhep0UjhVj4gxjDHw1IdutvC8k3Y4cx/HfmqwJeRa1D7ylPHViO
DfQTojUZ849JLWdB2AO9PlTl6WZ8kjsMbKhKu8Tmf8meS11srW38E62snf74+Gy4
fQLrxDIchLTDKmTLHlPAghu5OMSJDbZFXCm9kCdepdmHCOA0I4VamdKkDePyp/wP
XWiIIPcTgCpFp2Sv13hC09Qxt/R3YA/QGDl+yxeIMQdCNcUUtjr5Q7zA2ptxUFz/
BFfxK/KVCVeVUU+v7iLPL7zoX3w6OGeZq9o2VX1XN9AUTCtkt+QVI/1kad+9kciv
UMkK3068cKPUEi3FvNmvmffQgX7yKAMYYMjJ2rZEo/CYUwsGL3jLkXggt0tMjIvw
IyYHxRp5gd5cMxQ/uPlwoOPaldxK/25DKyUmaIuBOtbrD049gDHmzS95ocw8quXx
qFAOVWW7c2jxoHhbgEK7WBAejZpsSJd2IY6w2b4oTS7XsZ5McAUD40tBfIQsKF4E
ej3ntH4P6ez4BXbT5sKkLeESQG9qBGg6+a2fyrqYdohA6na/YvrUSkQ5M0jAnU65
M6FWSB3cmVI0f3/JJ/bsLgdMMrpNFikr1ErnzcPuNsN9uHll4Flh9Tli+gZN/dDO
3BnYLRjlR3sLv9lMHy3aMdpxYp06xG9mco0TLGjy9V2QPUCVvB7t7dmtNPzwF6hR
IzCDzLmp0q6tnSuYYcZf5eJXNxPwmF50xU5Ur5UaAXqecnqQxFgyogtblMgLKy5u
ngSmkG/L8EFNZI7nfXruZMJzK7XwouKaBlqe959XgYF8foa1iRMU55nrxjesNSeK
88IRqpYUsT/aqFUqlI47jaLx4U4rnhBu8qlOyiB63RHFIRYEdotRZH6z3dJVq2XN
TSg84utOwair9Uy/bYQ1cYErGdENoXRpT+dd7xp/BmrZYhZGihHsnefdoUbJHSYA
N2xLYZC83jED5DLsWBNQgNVJWjxsN4RDGkEqygwk7FDP7UkoNOVPVq8KsTzNU6jA
j6/FtlE4/lG3zRWLpvh58pa0U0WcIyLb1IJDtvyKAx55tS+IGD8KJpL13juIphJ9
8YNvvTnNx4U4gNrJfDuCtgjZxb4fHLi64YEdELIBf+zK1BLUQC9fKxkBvbEUhl6a
qOIvnTTXT/cuo42a2tC73m4C/r3MdIX89FsMdWX9FCfvIcIU2mo7qxYvE1EWvb+B
TL6Ywo4q1ghhdZYaqVQbb7WguzC6IIsjtNKA3A/LteQ0E3yQ73Qb5ezQNY20WbM6
oT5rF0n9Hop/KFpiRw3Z1hU9OT5XynCRcKqSbnSCqBARlTv3/UckPSSbj8FclyNn
JNraDdLlXueG3Cd1WXyRTGHZzlaUIIViVPuk7cPxENR6Bs6bcotR1yOxnb1zebAN
THm/6suC1UWoJCNDNeE4AEMGUz+jscUfe+MwJUf9iI2meCE29P9/j5qK8R8Pbcb6
PbCHGMJwzQZJAnmYbEFuNYrTzYe42oqitMe6UJhmwhtgljx3ziA9oRcQZ+7EM0wk
bUUeVNZd0k1NohIiXyFsIHzigbKMeEIH1cIBSd99WOOixwvBWRiaU2nVgbQfpKx7
yta+kX/sh4Hk+jvbp5KiSptj2HunIp7BZHVIqyYFKPMY1ys8XHXQ1XIUitK5ZQpT
F7kMmtm1pWVV5yos427r5nv2hLRRDqs/eI70qi+KPeL1ZZIMzTqoctPpL/jBDu00
YT95FwOIfA6b0hcLZTqUychtcN0RkCMgqUDnoEdGLsctimyfs5GG3ukTWy0ldmzc
KGk80sMmW6Gg3QDBhLqV89hFIKAMI7tZ7jQPzTkJc3QMov1OfcCV6bpaUoldQvXX
U5pZBqs2bpnKLvwDY03UBqGuYvvB8c0s+CdkmtinH2egg6N7MIXihO6WKWLZBqxl
1U8YxrpL67LgHvMl9btBrP4MUxcTL9Ah1LxuTk04/RhVGxX/yBM19dISbBI5JQZi
f7K4oUQf5icRptwc5UZQXO854Hapj39QJYPabofAwNjx6/V0131S9UqmnVCl/+B8
thFypu3Jn7e1UzKfQC0C6/1qJGHhkoOPA/kEYS3de4N4T8UivPtoXyTHTrR7kFcU
PlkGPQ865SVqcRIqAzYbhrX6qQau4CIZHyf9oCkGhvEZHeiEAdjrIrrzhNP/9JnH
Ue04238XzN0aFSz7q6d7j1DODsnlD0keEujPQiGwAjkH5auJFABIs8SvqnKTd4G6
x1hd+1/teXyULxqMYNjytwzOeypnJvLDI7EJ2LuLqxHh3tMUwP7xOluAmaJ2y7UB
mmWuesAwZ0hiSzgwTQnumXj8QQHDmKAL2oqaid79GxPX+6bUG/huSFLS3LmfI64O
yP4C7+31ma7r7nuT1IQsa1GhlNMNPyj8XMw9SX2ZHTE2W1A8ig2D5cW1YbTM+nc3
H4FliuzBAuWo6gQF32EtI/796V+UuXPPKGn3gOjokJyL2GFSniSDZfJT+1WrYC1E
z3mkhT4+Fx7ZDKbL8qxyJgDax+402P2oOsKHvFnzErDgpEYnzXVa0x3A4iUMBV3r
RFG2P5JagliZ5TDaPWXgA4ot8c3tASyAiGeLZm00EY9bQtxeuk7a+sffcIWv+1UM
3YOg7e3vPuthSXhXX5zeuzmGpfIyz/NXxl85N4pHJeM0P4Fy1Tfxq9ekeiIDkh3O
Lhuj09V4EgFVYslbGNpJHW/P5Nx8gXVrv5UV1dHE3mqh/UugEjRKt1JPcH51Tdsf
c/cGWy8WQJhWC+aJeVduqbsSStlbEXa5h6ho81PtMnHw4ZkS0tNI4ZxZ5OnmD8VP
7cbxtPguwIu4nLIn3xqrSw8XyZXCq1nNHsCdRK5ReUzAvVwSgywVENssOoG2++tw
fizKCvg411apOJL4vwYgosK0cPqMmRlR7w7Pe1+zR9gbPyko1US/ZaXvnWYGFpaS
6WDMdpTLMLrAG+pWwoj7C0YAKJsy9x+zau1f6Lo+Bpj7kspLinKoBoyRGIRtq3FC
5VZ9BnLBLg8q+YnSlI9gzThO65c1fHNEDEy6I2RZqoKhMfVeLgAymqZdH2Yfj5k9
hjYhUv4nbULhuYSFjHygk/1/3KPe1qZYeBgj88q4ibspphgLx0hs/cCAdLkaD9C9
kgGju0AUdDCRR0HlWO2fuJW96Tcsug+9hbu2kfwI6yEExREF/IJp+LxwvjeJfvoD
HcTfZ/+z/pOwLGxhr41pLP+r6uOhR0PakdR/Cs5QRR5VvLZN+/XBFpK2xw4jCUpz
CiqJW5Ee6PLA9IL9AvchkOfNu4njbrpRGZP74dpq+np/E72eLiyabxmsHh70FFM4
i4JhTe+fvSHLbeHo8Hr3PJOwOPHmXi1fd/MyD23i4s9Tgiz1jVtojtx3PM0BEUc+
VSqHSCi5EHQ4OAVfEDzoB6t7lDLlNg6UPsQkSSXWXWivfVOie7EiKJu3lWaY7rvI
uYc8RCyhdxXV73gjhiywP8RnOfL1dp7iiwNcOmcBLq4nylmBYne6eCGEKbb8K1Ye
61QQyHDUYoKPXK5RnKZ0XvIw5t1UwwaWQZyBxaWabtw4TYDb+k3Hgzr7i1KWczut
S6ueCRvoZToqwQIttAPuJcTBPabjS23+1KFTqViLGMCuwxph3n4rJmq+e5jVfsBL
ox3MRa79xw2uFB2jKtEdGNMazkwhY3dSkb6eyziY1T2dkRX6xarjjFhp9GhoXBTi
/Pd5iAu9Kx92evNTbdKVkNvwsLOVlMwLuzDwdo15TgdVg7hlfo+GFkrqzo6QMRfb
fRjz1jTunDf7FR5yGxltW7sc58c8HoCb+18EjF3dlljEXTLcP3h/Le7reIlWE5VC
nO4i+pQ9sd5epSbX9j7KNWpPUZR2J9gBFIfAqk1Q0KO4nqO9tIR/M5knv+V8+I7U
zGi31cFEhYVQCvHG6/fx7VaNAntB/o2MMXmuy0yjuWU2UdXYyv5mORFhPabQhj23
5Eb87mu/qLwFg7xgH9MCodM9uuurg5Lw/ooKxrYVlLQS9sdK01+Y8PxzgnyMieIZ
V64CEnvqPQR6CiW0G2KshYxE7tzgqxlrCzAGXObFt6xit9cHx3V6Cq1xak1shWWV
JxdC1OjnuTpZ5HGtyW8ZEWeFMyfCt7PM2Bn7mslqbDMMVjVv0/Tv2AEcd5Vg4mRy
turq3u36pRa5qNx//A7DaT5BRnKTMUKnb2scdPWl9wHbpgkXjkyOmIkIeIA7PmJX
ZVey5mZysQABTJlQR34+L5ykDQYhbu8jg23UUXbGu1m0jEIAwHI/bIqtdQ2nXo7q
eH7WgPHDdLF4BWSLFfiM5LSuTtLGPXXQJLjEnKORgyjziOmJmsgixA0N0+FYDnSJ
68PXNw3ALyRgKQNZj7haulMN0bDrQ+fkEKQX6K5p+fJtQBuvdEwSaLE9Q7rXQ6J8
LRUDi8SPa62+g4N5a7qG4Q9FhryKPXjGY3Gv4MftJGtsTmcqO6F5Y7yo/JNq4LnA
NI8KkWEeG0YNa/xz9PvKMx4kgWOm1530P3taumLHulyuYKyFQTVhaxeNvwCEKz+3
AqC8N5h9XrtX4Jd9a6S3eGvVFzI43ONLloRWC+zfI/xpvWyroqCXxohxxk14/31p
19jo2CErExR5ZsjDq+LuT08tuFZ3Ml1zYV4hl1JjsaFCPI9gUQ95EXbiB5M1S0ZN
Cjd8AGdMvRlhPfSFmFRX9ZpajOgS+yTmKdUpCdrthvLxwtkRC1qPcxIzN3Pf2ivc
6hjGXzVPfkyELZmqRJIZHCl4b0OirSViar3+Y/ji2Q92ZHoWh/m9CphlxYaS86k7
3dlZnWMx3a1kuT7sLPZqWruPVOz0hfSW+vZ+vRI7gOOZ7RoOdsTmRSEGQqrvq3QJ
erOsGd/BIjkfk5CuCDQd8GGMdliuuLvQEuUiXrf3JjvKF7JSKEHtVtGSymy1SKqS
oukV+EMt6TRlLWf0n8vN0Novb85NjKSYHJVAOQ56BYHmx0C3CwLS9VeLe5nxjDjj
COeJj1GpSsDenfkxa5XK/nKkMwzMOK270cSgn7p7qX4Wpxik2XhhHD91+/b2lx9X
+CtntUaULvUsf5899xbOtI3Rzh/LHqs4aUfhx1YtyFhsbVWM6fsA+zSSsf7KQPDR
YicJqOGWy2WPJm4jGQPeO/xtHWK36+xeYFlqktyS/nGhTJ6aCK8Is0x7bLoN0Z+e
sra36/OtZVcV0M1xidmlm6SFMi0dP/x7rGQlzyVYXN+Z2M6hZnDpRobRqFvs+GZB
+IxmwN8aX6H2Pug4R2zmPLnDQnhsJCXPYrTN/2AnZUKgcGt4nv6W66Jc9DbhKz5j
sMVhvFQSXW8JJ2eMEo25P3+a3L2ERaoT2mry5AVkBOTTHDZmkLUFeBIpp73wR2Ud
DDwlk3S8nF6FknzZ8RALYnngRNI4AmjDeKl60qJaKOx7kMKfuZG/I0FkkeHrV7d7
mD4WG+SaETeqOPCtpYh36F2cN/Cae1Df3FTqnDzBLpeuSm1oNThfmbSOyA81ODHr
V6n1laewNRbZyqe/UP11fbOIq7eOK0XqJf8SKDT10jARFbxJ5mAu9OU6VbQWu89P
ZCaD+jF6Wz7u/IuxcnCiZvZQYRmM2E+E87e+9KnY0m1j4MKJT5ejU7DArbDXuNSX
cOfwClq+aHMPlpHx/RzTwP3Lom+SigHCZg2wxYBckm39imnAHqyYoUjAE1YBFwbY
UiH+6sElYJ+UAC/9NcxXaK8yGcxWC/IlDOYis/wE6+FBouDSsjWDazS2QcKXRr+F
YRH9+PjTfee0jE0r7WfuUL1cegsPE4rdcVRlAFhAdqehdYQ+yJ6B6nOyNist0Msx
vGzyKx998BBdzuHpr5ts10IcgKtK7pcCFx28PxXmpzv550+IJQqNvUMaW9vZ+k1B
H8bxLMjZgTVadArylLExhwMZ3VvIEtDcc+tNWqwkJCKFT/2cCqjjVuROxK6bzV85
iePZRuEFv/FL1d67XEake4I15v7hd9W7f0JvmrtDTa7J45juNhzsj4QFpOtZIGrU
5TUjrrjyw5MzMPMaNbh9iCaOR3bT4Sfcdd01B4KIEESxb+zUB2ZO6lO+pltrI413
XQoz2biSC0/fO2qgMcj5vhefTTvGkZ6z7s8UUQmaZR1c239yg4COS2CbtitKWwP6
flHY+iV7WJsU8D/UE03mNW/VczoA3DEl8lqcnfAQgOasQnZDD6W0UmmroUnfFnrI
1gjLZ9lj+tZBoUK9im1NPFBuPZCunOVVRUgBMkdPLZRXaIWJiAgexc9eQVGdqRJ4
+RCC+cA2ADcm0RohVKmLVIza/SXQZNdO3oy4IOEyTVF16eFGCdCzxGCVGKBl4t4q
EjL1wiA5Ih2ubgWZseVdNe1Rzii6lJQOAckWIudskUo678aX2A6gB8O1u8cxRt8G
S5c8UZFezenZIsjGj4SKZvVhhZlIRb37cWiruH0fBVPFnEb66t6f72avV63lNbqK
R7m5knfJLHT3f7pcF84kLw2vwhaUB8zr+Tl2asstlqu9wVqOT6z43yVIbkHFcyce
Rl2f3MakdVZeQ+d9VVujiKG3Y0Ph8djL2T/JLU3LgbdhINaQbaoRJubssdo9/yls
CnqmUfLrnpaE6SmnbgOwPZndlPkzZCgwnS8xo9z2S9At/R66l/4WULYPDR/zOstj
rqXCsOYouGxHIpDQ7+XvsunXRw96XCTi3VdgoAoUXvdsmF9sLHsaASa6f1qYbc0e
j85rSQKTQmkjWlPELH5tZBRcKy8/Ff+hobxGWTRkii9PIk7RwIG+dt/3eHbJv7wI
gOU8n+S3y05uIA6vcANRVhg/N5v1Fm/Z4dlnTlgN6NNk4q0qfpNsLZt/YwmsCdRc
XDB62lhRIGxmaMNzilrTNfngVHDiOxeDD7wTwj0KGyNFUq8bdwOWllPmMtQOTgPX
XOVlx+dsA5nf6QZgCfEGXAnVU8tjq1sjnGVl0X2BAQCPrTX5DaALrMBibwg3uh9F
fGEBYLtXFvXHnu/ou4giIyeqs0dzwdHJNzH7t9+8Y/uszqgvwrVLBGBFcAs/uIqp
wWP2PIkCOtqEUAr5mPNl2OmMDk4psnEii4h+NrqySgZ4fsV6WBKqjaj6AwjNHbnu
Gcxn+0Ojt83dw1SUXjQRu7NR2e2gvpT+WgWCLFC+ARyqlWX4HVEGyXQCUPddGoMS
txAC2YwGQ1fVVPyyFwki0Rbr/3VrD8J+aaUPdCG722/HSWOOfXtFuvi5Kwuobj2h
7gFsW48zp17dSZ7ejfmVuZjiiND/rQqJNaBucUlCaT0PcKDWK8exLJTE4zAygKB0
wDTA8P8r9SBgx0pBVqgO5JrtZmbnedNfHsK5hYvHuBa4WXXYY5BxWkBagosevjHw
4ErqmKzCz5qJTjWiNpPvNF34B8NO3ccxHVnn3+ca7fqJXV2bxfZPtSDmF5g9CASt
m2fQlqrFWHJ4RqukpPtESKTWLq8/b1gtYJ7muuP+oVzxbW+zzy4FEomgCS4MU5mF
aeTkcP5QfzBiJyrOo0br+ofM+tuZ5RpgrnfN8ghG5O9UucAUtZ2agaSp5OOIkodL
N16WyNhw0IjG0R5qn7c54n37sPOMIp4GLLP4NWjdjBsIuXM7yuhm5/dE5N8RKqpx
h9/AQNgtTIVDhjaHh1oMy9cCm/N8yH0Z2yUtVadq4Nvyp2k4eo/9/JTBLBMajZYk
m4mLPBkS3QeaAsXU8uMZ423Qxw43A8NYfkHUgbci+yweg9FeTiWXYESqVAl2+upe
9TexQSGC246CXyTxCGHa65Mx3YHcdfgUXqqio7ttjLLIoHx2gPALnS1c4bnzQQVq
NlZ6ZTaqrvp+Of99Curys4f6IlEIlL+lld791Pw9sn2G0OD2o/qHTXHn07QRAKcq
IiahQDU4NFAEc/5wKp1e3t8w2b82jqJFEuiSaSLNnqRYkmAatp66w4S5hIQXm0zs
+QK02YowR2tgxAQr1+NVLO+5BjUsDqeX0xvHpp/MnhHf2MIHjoQDZeFZAHJjTb0x
LIkVTGP/g+kxAeMiwQQ8s7LUds9NP5G4SJ0efcNht8XKDERFub55lGvfe7mNchZg
WI+o4x6LDu8CEEpJ5O48WYNa7p1ZSlf3nZK4eklC47zTW8Bax36EWYY0sqNKpBkW
mX+ZYqFe8snBtb4z3Mpe3ZG/d1iMyIORIxQMkwRAzMVsfnO+Pokc7UkBki487UDq
4Cwj7QQGM09r1YmOAG0haaO0/MgzeEieVJlBU9exw9r1oT/MiG4PJNhfntSHgzel
CDfG5gBUbeRoe4gVLFHJUi1hnuViH/tjNGFXBnb0/kEDLtOTUBQpA5h+vODHw/nK
XNNgwp5ayUGmpdIgx8l/O9+T9/TjikgOQjEWWK0aDnglpafAokwBne7WdEpzng/i
GYH3Cs08KKVZOHj3MSsczqsCdA9+COfBcLgBakINE1dpIxnn845zHzwxYb3tvU2C
g60+ur1TTqifLxz1KTVCgCAD5wOjapaoSAYhuNRCrs8VClocQcBSSVU1fUyGtGfN
BWnDG/J4LH9V6s/Jph1CMZC+385ZiPPu4LSmitE6Tsqe6PPXVvx8i77sSoCJhots
wVTexpXXUmSt+xb2zqfKfULnKCIKAYy4NDgDx4YCWBf1svC8LzJVpBpTDLwYx6tL
OuurW0cnmzAN9BLBG0+3mF9/0OnkjkidfxBHhHJ8bykyC8d43TImP64uWBanztOV
wtZU7AlHNCzujgPP/LZrC+Fw+I/0VHwtJ6FtyE1U58UlloPagqtTXp550mnMXpoP
Bh/TG/zRggIkIjtfaPp4KKyKlWXk/bxQUYEr8tLqnQpIVasTu4ZRg6kc5k78++eA
vlMMRpzAdRoCSFIIrvNiapLobQm3VxSE5nRPWgvh5FHF08ioCdD1S7Yiz0uwUw9S
88RJeCIfo0rX12uVBv+r2x2soFxwMic2TO3eD07AJydqwdeFdx0pRc++t2Sc4OYr
mtFlYKb2jcofREmZBrN/jnrlYOJIn2QaoUFMD6AiIQWlPZMMg89w/UTU0VULr9v0
Wg/ZzgfPnluflX1CNPZQsmSI3dSCG9Opow9W0geLSuAqZbqjRjXw3aEJi/W2Q8ZW
uT8AsMIFNZ2WNnXPwChNKyuVu/VEmT8aoA7FJlegxlDNzXxOuUyQuSIfuA4h22cH
oQHuTA6ivbl2s0rtrgy91Y1s81GXwT1PfZIDdlti6V5En4dRMCPA9gr0TWk/NlhE
9RNN5WpX+9aOdJ/T7CYeTtqpjwDNAZpWrlWWeqvHmp6+a27n9/u+znrOPsmcNr0E
EbP3KV/LMX39n88MIxxAm/HYWbTi9+MmSE3fO9PjEEdXpjPIIAiabflvqExEFDvP
s2UXb9IfWFoWJ2VDYZT+L08rMdV0mnOQE5UymeNOAj9R79mlETpr/XXRPgqVxrrn
sHIaDXpperhAlt0WoivY7fGEGWhaF4TRQdrsxHFNkheA7sjb66VsNx3S294JQZ1O
9i6AsdyIXzTmC8hguBSiKZTXBdqjEp4IIUARfxmkgOV0aYDE8vM+uQLIkmKkLODE
ifs1VVP5oF94xtlkSUgiv7AgZyTUb/aPDOsco6SnvHirGYBULy4FXX9Of+mJaVGb
HSb2qnUtPZ4pKQQc9tLjYNOP1WsvZPQskgaDUp2UXLrpzs0qvOF1Hc39n1WXlc9J
8No7l7pI1rdH6ZlZZgpBbyW2Ct9lzcIBnjT17nirajA5lxg68WJtKxP8+KC1aoGy
9t3mZ2G6wzUHjdrPV7Svb0O8H7y6cu7l9w9SSIe6/Tu6N8hcucv1kB9j6tfV/Ce9
Th9R2G//ADXaDjzVTmzNXOLQHwJCt0Bv+Inrf+3VUZKmabkVrn7YzcEDXHF46oiv
r7Y8Y5XPeGSm/oZiMH9yxuYITopsfs/AginR+UfZYEe81vEh0vyRd0RM/Y+ScMCC
SFha44QJ86V2lhMeUnOn/xq5rm+JpIevG1nMf0wJryuJ6y8eqp+MFD2Vt35+Bl09
hxC+/2I1UnSi/4qjw91MxZudJzQok/kw1+f4qOBUJ14n0dvI98vincvoYQmGhe7V
fPGUHhZ4MhUG99IMfvc9tb/SJqRzenHPZWNnV/Ma+8hUNxayRXMa9ja6JWcMiRSO
wJNaKQC9XdSwH3NOuju/pp1ctvDWY9NkPgwtGiz1wWhyfvIhgwcDzp0Ck0gPVDMx
w7n8uwf9yVo5IuDkddItJU+Y8NbuK3IaaUwW0cUyTSUOlHSvbaw9x2iWDLi/vAPC
4LKmpVxb+jkDDk0QWmic6XCE1YZ89OCt2MuaulH4d3xE1GgKx0tzV32RSP6fAK7o
7J351UHvIndFzOzPn9Pf0Q==
`pragma protect end_protected
`endif
       
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
H0/ZRNylEHPhgQJxUZY1peW961PPXHG1ymg+GOdZDdwmo2DtCikaCF3+TA+OHAy/
ajxF1kPX9VQ2uD/DItfTSZj4TZ7AYzTmejhSLva/4PPdivxSo6YwIOygbwW82vLK
b+G91j1MdCrCONDkcXIJigp/cCfXlnYXs8kTTFCOt84=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 212387    )
p/DZTUo7kX9Xdi0L/Ou2syNxZhutxSLzWd/C+DOT5fVBI2FO6s8Eb6mMr9ZfLUeY
2sHZvrsiUfVfMVLucDF35Prk8brM6DKUVQpyJR+gq9q0+UgzaEKyprbo0yyqCJvh
`pragma protect end_protected
