
`ifndef GUARD_SVT_AXI_TRANSACTION_EXCEPTION_LIST_SV
`define GUARD_SVT_AXI_TRANSACTION_EXCEPTION_LIST_SV
`ifndef __SVDOC__
typedef class svt_axi_transaction;
typedef class svt_axi_transaction_exception;

//----------------------------------------------------------------------------
/** Local constants. */
// ---------------------------------------------------------------------------

`ifndef SVT_AXI_TRANSACTION_EXCEPTION_LIST_MAX_NUM_EXCEPTIONS
/**
 * This value is used by the svt_axi_transaction_exception_list constructor
 * to define the initial value for svt_exception_list::max_num_exceptions.
 * This field is used by the exception list to define the maximum number of
 * exceptions which can be generated for a single transaction. The user
 * testbench can override this constant value to define a different maximum
 * value for use by all svt_axi_transaction_exception_list instances or
 * can change the value of the svt_exception_list::max_num_exceptions field
 * directly to define a different maximum value for use by that
 * svt_axi_transaction_exception_list instance.
 */
`define SVT_AXI_TRANSACTION_EXCEPTION_LIST_MAX_NUM_EXCEPTIONS   1
`endif

// =============================================================================
/**
 * This class represents the exception list for a transaction.
 */
class svt_axi_transaction_exception_list extends svt_exception_list;

  // ****************************************************************************
  // Local Data
  // ****************************************************************************

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

  /**
   * Array of exceptions, setup in pre_randomize to match the base class 'exceptions'.
   *
   * THIS FIELD CANNOT BE TRUSTED OUTSIDE OF RANDOMIZATION
   */
  rand svt_axi_transaction_exception typed_exceptions[];

  // ****************************************************************************
  // Constraints
  // ****************************************************************************

`ifndef SVT_HDL_CONTROL

`ifdef __SVDOC__
`define SVT_AXI_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
`endif

`ifdef SVT_AXI_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
  /**
   * External constraint definitions which can be used for test level constraint addition.
   * By default, VMM recommended "test_constraintsX" constraints are not enabled
   * in svt_axi_transaction_exception_list. A test can enable them by defining the following
   * before this file is compiled at compile time:
   *     SVT_AXI_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
   */
  constraint test_constraints1;
  constraint test_constraints2;
  constraint test_constraints3;
`endif
`endif

  // ****************************************************************************
  // Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the instance
   */
  extern function new(string name = "svt_axi_transaction_exception_list_inst", svt_axi_transaction_exception randomized_exception = null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the instance
   */
  extern function new(string name = "svt_axi_transaction_exception_list_inst", svt_axi_transaction_exception randomized_exception = null);
`else
`ifndef __SVDOC__
  `svt_vmm_data_new(svt_axi_transaction_exception_list)
`endif
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate
   *             argument values to the <b>svt_exception_list</b> parent class.
   *
   * @param log                   Sets the log file that is used for status output.
   *
   * @param randomized_exception  Sets the randomized exception used to generate
   *                              exceptions during randomization.
   */
  extern function new( vmm_log log = null, svt_axi_transaction_exception randomized_exception = null );
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
`ifndef __SVDOC__
  `svt_data_member_begin(svt_axi_transaction_exception_list)
  `svt_data_member_end(svt_axi_transaction_exception_list)
`endif

  //----------------------------------------------------------------------------
  /**
   * Populate the exceptions array to allow for the randomization.
   */
  extern function void pre_randomize();

  //----------------------------------------------------------------------------
  /**
   * Cleanup #exceptions by getting rid of no-op exceptions and sizing to match num_exceptions.
   */
  extern function void post_randomize();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to. Differences are placed in diff.  The only
   * supported kind values are -1 and svt_data::COMPLETE.  Both values result
   * in a COMPLETE compare.
   */
  extern virtual function bit do_compare( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );
`endif

  // ---------------------------------------------------------------------------
  /**
   * Performs basic validation of the object contents.  The only supported kind 
   * values are -1 and `SVT_DATA_TYPE::COMPLETE.  Both values result in a COMPLETE 
   * compare.
   */
  extern virtual function bit do_is_valid( bit silent = 1, int kind = -1 );

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Returns the size (in bytes) required by the byte_pack operation.  Only
   * supports a COMPLETE pack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned byte_size( int kind = -1 );

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset.  Only supports
   * aCOMPLETE pack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned do_byte_pack( ref logic [7:0] bytes[],
                                                     input int unsigned offset = 0,
                                                     input int kind = -1 );

  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset.  Only supports
   * a COMPLETE unpack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned do_byte_unpack( const ref logic [7:0] bytes[],
                                                       input int unsigned offset = 0,
                                                       input int len = -1,
                                                       input int kind = -1 );
`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Gets the exception indicated by ix as a strongly typed object.
   */
  extern function svt_axi_transaction_exception get_exception( int ix );

  //----------------------------------------------------------------------------
  /**
   * Gets the randomized exception as a strongly typed object.
   */
  extern function svt_axi_transaction_exception get_randomized_exception();

  //----------------------------------------------------------------------------
  /**
   * Pushes the configuration and transaction into the randomized exception object.
   */
  extern virtual function void setup_randomized_exception( svt_axi_port_configuration cfg, svt_axi_transaction xact );

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object.
   */
  extern virtual function string get_mcd_class_name();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_axi_transaction_exception_list.
   */
  extern virtual function `SVT_DATA_BASE_TYPE do_allocate();
`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: Provides <i>read</i> access to the public data members or other
   *              "derived properties" of this class.
   */
  extern virtual function bit get_prop_val( string prop_name, ref bit [1023:0] prop_val, 
                                            input int array_ix, ref `SVT_DATA_TYPE data_obj );

  // ---------------------------------------------------------------------------
  /**
   * Add a new exception with the specified content to the exception list.
   * 
   * @param xact The svt_axi_transaction that this exception is associated with.
   * @param found_error_kind This is the detected error_kind of the exception.
   */
  extern virtual function void add_new_exception(
    svt_axi_transaction xact, svt_axi_transaction_exception::error_kind_enum found_error_kind
    );

  // ---------------------------------------------------------------------------
  /**
   * Searches the exception list of the transaction (if it has one), and returns
   * a 1 if there are any exceptions of the specified type, or 0, if none were
   * found.
   * 
   * @param error_kind           The kind of exception to look for.
   * 
   * @return                     Returns 1 if the transaction's exception list  
   *                             has at least one exception of the specified type 
   *                             Returns 0 if it  does not, or if the exception list is null.
   */
  extern virtual function bit has_exception( svt_axi_transaction_exception::error_kind_enum error_kind);

  // ---------------------------------------------------------------------------
  /** 
   * Utility function which generates an string describing the currently applicable exceptions.
   *
   * @return String describing the applicable exceptions.
   */ 
  extern virtual function string get_applied_exception_kinds();

  // ---------------------------------------------------------------------------
  /** 
   * The svt_axi_transaction_exception class contains a reference, xact, to the transaction the exception
   * is for. The exception_list copy leaves xact pointing to the 'original' transaction, not the copied
   * into transaction.  This function adjusts the xact reference in any transaction exceptions present. 
   *  
   * @param new_inst The svt_axi_transaction that this exception is associated with.
   */ 
  extern virtual function void adjust_xact_reference(svt_axi_transaction new_inst);
 
  // ---------------------------------------------------------------------------
  /**
   * Searches the exception list of the transaction (if it has one), and removes
   * any exceptions of the specified type.
   * 
   * @param error_kind      The kind of exception to remove.
   * 
   * @return                Provides a handle to the updated exception list. 
   *                        This will be null if all of the exceptions have been
   *                        removed or if the exception list was null when the
   *                        function was called.
   */
  extern virtual function svt_axi_transaction_exception_list remove_exceptions(
    svt_axi_transaction_exception::error_kind_enum error_kind );

  // ---------------------------------------------------------------------------
endclass

// =============================================================================


`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
W2dGzIRVlazmq7m1gOl42aI6SNUR1aWrlVPmEoBEODXW3CDaJN8zZ29sH0e7o3F/
RqobAVJVVUpWmE6Mbj2NL1BKs+FpXZHrlBcVr7vVNdu8dhsPMBbltqHRVNQllVhn
frDZOFA13ibDGkK2LDfPbOU7ZL29MitTm26sdi03KVc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1325      )
+VGjCKmEEqwjVDRMSpWGuu/QjwrEYCgi7Jyj5mUvigQYTcrGe7MkmCI3Wsuq/f9c
AZdhtGPDFHByQUO2rBm3GOyh0xhZbMS7kOttTXxdJTtKcigymhW4Ve/b2vFpQDRm
vWKc2kfNxdMPiogTXMGqnB2VwHyH73XFx3iDntrqqNLO+XD0d+EaqxXRHwgeVjDI
+SGQibVeqUmOHUzC9czbu/aGUSQgwBSA6HYczC6oEv0q/5fMBaooMdBWOIVSFbo5
1NE7EBSGbeE9ik0WNg4OWW6hPHdYEgVUAny46cNYxljl42crgWVTbmHIydnSe7Jn
SDwjUTba3gOg6UKluInmsGQ72LnBNLYTyq8B6T5G8JVbBablKUBgVHnB0atVXqti
GqbKsGysZxXm+AR/bG9emyiZ4od9EPVeWHJg8WGTnUzBiE4GSpjfH1Mf1nU23UlF
t6ZC5I6fNFVabeC2E1ORPaZZZZuhrALNHj9G2wPzR956Tg8x8jwG6SVE8yocW6s0
h69S7oK83ubH8h753KyYtjbc8HpINarkbkJXieVg09ThJ0tuTrtMiQrkSJKDO11U
K6EbXxiT+PEXTeQw4pCg4maOEGOD+KNEq068NNWg2i3Xc4NvFv93DkwkseeDB+0y
fqHgc+J/NsYIDG0XLt45tNsHe9K7fldPuxdZUc4ayWcNJ5C7vMqgj6r6kMKpA6nC
/wN1hHJyFpALHZxuYBFv5P/oF5daufJ8+zOxLvTjsrJ5SwiJ0XdhCO+Dydi0dwol
VfwGePEheMqvqPHn11T3T4XMLjRiceCYB87B/jtMhXx05UUlNsUayo9U+gwXH8le
IeXiZRetkST9KeszOq5xGPIh7j3HgJtQQFyS9BcxeB3eZXM+o9fgdriB8s5J3Gl0
wWUHT45nIERj1DKGTcsRpLMXCPuvnKjypLYQgOMr9yjTB1boS9rC6gZmuBZnLBsJ
E9mYtJBh2YXgJ5qRipsMjqm5komQejQS6YLFhKTiR4RNVwbxrG4ExGbdGWZf3fFm
i95YjTec3VZOhIRuqN8OghS2qrVAegpz8W0oQiSofHsoE5KLEtR9NATCfxr4BeVd
Htk0JAdu5gjEE+T8JLpbZNYukYAlh5ttYAbmsaq3RnR5PjNbldFRVwFT3UTCRQjg
DREmvkhiiemH32Q/kaYRNsClu+Bn7jotAo5W+UtqJcO+9jQeg9sbIZgMNzMzGTOX
9fQ+hYQ+HXGX6qdtXOBUVviCKk9U5SHVGXI1S3U7RUQAj4oa3OkV126tFUNCns3p
hcgEFH/f9KdozZ78IjI93vTXq5Civ739F/+ue07XxA6WRGkeMrX5dWL+gPrJSq6y
EgMIDjW/dlSDD8HwLByjs0E33ka7roo3EfysJChNpJ/hunwTpg0iSmeTQXAmwz73
KTPxG310A4ZFMQlp+8SEW+DTdxs9N8P6tvJRrCR+Jhs80I6T/suQE/tcQwKW2xP3
dUv3l+3EhYGK58EifLrIc5sAAzUJZgjZxyXQZDB68QpOm2heCuuhI+5Vb7G2jN8x
/iacNB3iOP7Nfc3XDpP2QWFJA87LEPsOlOIqI6f4H8fGnoBzEIL1p15MmZ2+CYe1
l3gqt5aehpthkznSjmz1yb6eeFaZw4WK0Lb7tAeMx2sJo2yMs3WkuzyhRAla0Htw
jXz1PSyIONaOly8ZWa0floUqcxVFymAxA9Xc5MWaZmnSEUmT4rkqfrSo99o+1H7B
1pAgCFtRKYthGdLmEu7JcVDc7Yv8PITN6s340BkseT0=
`pragma protect end_protected

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
JRJOj92hZvbHiLT3OIAogz1LOeFF6RJlg5/+tm3pTbCzO+MmfDV9hqVdt+pJVyY7
W06QvhDUC+frHRNoiB3n9rsHb8l05ZgFxIM/VD4KD7FmBoktzQQU9bDxmdmiyk2a
aM95fjFY7NCGRqOU4TEwWokqCAMLe2zlVvokQu5J7gk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 19700     )
2FMe6K4e28lyU1Uf0KoePra10u3d4dQwAy9G5mkD14iJJWibxLDOgx4WaDsjcvUM
+S3u1WSj/B6rP25wGQBU83s/9caScHxn/MqRo+ldIFvReoAuhH4vBW6TfW+sAkwe
I9Uq3sJoiIBkZpOB+QZFmEf+YG90RqgetrXpA44p/eXIJ7qlu7TOBCvQH0bbxNX6
D3a3ashasHPF4l+oGpNgRAhZ8J1oI+g//sPFB9d0ntTZ+vWPx/eeYphVkm4u2qQ7
T/5GC5BbdjhIeWLvNj2x0GdqY3PT/VLQOusVouNMDcm9FIjP50Hb9GK6rlYma9SZ
yPZZ0f2EMW5xCUtLD5pdA2JbE/Euw/duK1D2gVoUUSTshMn3jxv/LJKdTbggId3V
c7UFObNdj+zv2b36Vu/+dOn6/3LrLxsIQ70oCpeQU3p6uP+mc8fhQhPyB4tecUEI
ZQXRY2Mp6q0UVOEVYJzmPvfHvdj6sq5+JqQFhDdxBfldrqL1+ZZgLadhYSsEDt8J
bKl1o4JTI30kGwRis6ZHAzWf47+WPF5//+BMSM906N60PCgJFwlOY31F6UJ9/Gwi
6zLbcj6q14aAgrk1UHr9evKh3KknQ6ke8Br5xqCqqW0xJyQ4OiebryQPyAF/aoS9
qwE0ApPFH2ocfBrMPtftdOXyQBMrMBNNc/Qn3eh50u2RDYTlUQgn7CF7sxPqvCVb
mT85UYgZ8Xuy7EdedHbsLYydRK8CBnYVQLQCAp/xwXa48NT4/aq979utkqbhdCPB
cwyFFu8Pnkuoar/3dnq69sfvijTkHML/yWCOM2kq8L5iNPda9f0qi3lSy5viTCU7
qnKMqWQrEOH1NjJwe25xvviacVp0JtLZWtVB3HIPSQIzdwYGDGjuz38ThLePMUbc
jLyyO2JWvEzc45Dq94TVr1QE49vh0XDGsB57hvFVAOog6mPxC9XJZf8oRTNb+wLB
i1PCuYeF4RRIUO5vWDrkee9Yg6j6QHa/9ATH/JfhEztDjLtVOuTAClqEEFR/kF2w
s8i9UlUPnm9j/Ha93NhY6MeuVyQVCHs3SYkAf0feFhCa/SgJBBKxBXyupFME4KI9
B/+zMxRvicue+bzV49vMPN+qYxFmdYrrhzrVGn36DZH33XUR/N2uKnaVhdDFtSJl
eO/0X6mlHnT68EiiDvRBGVbCUk1M/Dn05odEm4H5I8196hR7ReOYS+eTGcODBnZ+
pDnJE4AGeb2n1Sr+n0YUZ4/jf3ih3KudRRxdWArOp0BujKQNQ6q0e260eNaaKJzK
ZJz/9Az5O/mOof+BRwvWv1/nxjMuxuPcmE8jDfupwZ5NW7dM5k/rG0oFrVRL7TYx
cMJm/xWGb41bWz0FeIbAiFwX323Tg8RsRMjXyJ3c3SWOo1WeEd1J592jXlWVlmRq
xrW2WpwfNDS9WwmBf9XLwNcl2F5Vfiz2Y6qaEi7abWh3LnLdijeyFutjFZMnHjVE
+VbBzUe8E6iclknzOz1hxMTkiL+Kt1WXW0KzZB3+FbtHI5N7wWPB7FnQg+H1yYF3
fKcJCed1se1bUa2TRjcUkYUPP33qfJNT4bevUnS8NgCCY8h6JCaBsDTZ0cg0LZxh
gRXJsBVFhEx8pwHjNB40CCYGzF629HXuIzKTbMLPpjbgmdwqsMbBwty+q5Pnrr3D
0ZLx4ACkUwr20x/KCReaTf4lyixpmzwRZZLcwSXP5hm5Z0c/NQX5tQJtSCwpTyb4
uyXW+0iY43+2SkVw+U9nAh+gwSxU/VQwcQPW1/oJtGBEFA6dRYZcJo2JirUtVdHX
dCGQA2IN4J378WQztrxUKZPGhamu+k5MkFzTpqXg+rVz+fod6d2mLAgqb3Pj+98f
+rhAWuHCQGDuc/c98pIsloU485oEJ1gPxvf3gLg8T4H47PlUnbe9ejCl84TCb05J
6h8ILKkNBmw2/yaiyx2Nug/gQi8as/QXBDZM0waV4uVVOS/xkZYZjsNmjZsG2NSd
+CY5to4Q7qYebjv37Kwfc9S03CJ+PY74a+y6djTp3wspX3LzRbQGMF6yiZiw6T7k
Jt7EDycwfydu7PhGtrR5r3z38oFEHqTgYDu3T48F0QMJsKD0hRw9vY8LsaXbrVuu
nRfVhID1cG4ez6yIJWcJRqeW9FO+azF1ZZw8LJLOauqgr67PeMAepJuj3QT3a4ZJ
5+kufiqplHQ1GihJBqR72CNfUaokWUziExr0nIvlRx3MQcqR8NkIUGwnz/CaTD7F
7s1T8a4s9kiOlo7bl20Zh6wlcN6cIKrCvXwSywFsIwQy4Oo5GIpJPv2kKP4BC4+K
B9Okc+HE3kpgtdMz/jjO19vwC58cfPYQO9eoq85LLA0NIIBXdeVACwoi8NlmDYcj
GpcYPqOrP03lv7thWdFAwOCNrS3PdONWRdX1bSTMlF6gl40HrizFxbnOy+C/Kqow
jEhRudcKp8ptrV65es35f8hhsbebJmYjOQRujuVaEKY2gq9Bgk925lcs7c5+UwV+
XOduxnEKaRKLCQjwu71ngGlAMXGQ1vI5SZfMhpRjK88Kemhf3CHKoU0/BNevFFQF
HM+R1p9AARnZIbrJxHjkiTo7vhAFVDYVQCo9oNO4V+7QzbCBlmh5YW5nGP5/lGNp
Q3vwlWGw87K14LicWsZw/EVXP93gSkqpBQxvazzVAuCxkyA7+J6nL4BgR3zZeF37
0XeA/6gL1TyQi0NIarDrCh7l/6aF3rqV6CzRF5wAxCwnFD6GnfOZQB18l8JrzQCU
IFY0oV6o5YO19VccMplEEyqwh44p3BICkx3zf6W0/rk4lIfEQPMOs+R0sav/W8p7
XlsTcJfk827LRJhfilm6+DCQ2UgIM20vfvmgTzY/FfWTVa2cwlLzR9c1o0Oxurzh
TzqcL1m0bHUnnqDDTSn9bUkwTEvY8qSWeH7bS+kbXY81DSXVETc4Lc9mIJonWs/U
aM/iWtVqa+EC2A1zBf5WfXeKpOi7FAulNt97rbQiTnXGwjaNxwRF1oaOU5N5uG7Q
pwjrx2v/J/LDOC5AWgPmq5Il3wGYa+MRYH8KyJeydmdCrkI9wCjL/UEQLzHN+wwb
q7bDyuVCQgRtN+8lUDucol8OiuJBcCYcTmsoWdMOTTFjXFEL3RIJ1SydNxVFg4j7
gPG/qjEQyzfYj55uNWAxyOpQ5wkXcyG1khl8QcDblBjb1zwba7GVI/tBLmbfwf9D
qUD8kNwpAzbKKxrS1PLWdP4VAxYjj/UihBwLZbwut4xhEdtLfXAfUKHp1Tn5DY/8
xqiNRa6oUVz/ZLp8RCgd2+Mdu7xIHo2PTSzATMseLJu7ddMqsEhmioEbigZ3Jzi/
cmkxfDsk5JIYZObTbuF3x8MTQ/kGPr7xSvzZQF9AGbFUSE+ppf2YM1fKqqfE0/ao
kmSnEQRTkEcSZWVp1e46vJQ8FAWxZ3HhfJAVMNySur0Cfg9duq+T47q2B+yMCquM
itTuksEpgDTUj2HJl6omphK7cf7mSz77gMnfH1+cMyFwVABAJ/+p+29NiuvvI45c
25r1fu0pUR9sjdPRh5OYnEbc7EtryhxzrRMv4wG71eoOCEMS5bIrJGaZ1zKdoogh
4GzCI6LdIEi9K3bAUj8f6H15F33n4lq8E7B0b1jjwwB/WkNbT4mrZpwu3Tcu2+G8
YsPpznSTg/j8d0dWvBUI6lbQNlDYzUb/y92xppXA5NZPvXCYGOruUfnLXh1edC6M
h4eEElst8XYm1ouPEtITpi/5RkOUe34xXpUzSdndE5puGPy8VwH3XlPryxn05RXu
4D1pnq1ZyuV+1PIRMEdrP1FK/IxuoLbUAAcV+sbcEWsadkcODTl2C5dsv6UgFxJh
6KrJEsxx+as7fm2Ra7p7oM4NE/0GB6Hck/+1iy/v8Ta+Y8Zl7ugsZEz3N+pNfPMv
eMsrkD3mR9cv3OWi3k30nETct7DKqJb5us418KA35jNBCRsX7WW9OfbsL4Xvjm16
eZuKiN9CLdvP23246+/U2XQHPTvib9AdEUyvUlMQlcNUR2/BpBKwbpo4PJwsSzN7
pq9qLPMaWeinkYgY/rSoe9GhixKIH1LDruuPBBeWf2a4DUSVzR/bpJTEnOdzT2J7
C1Wlfh/L1Rd3xC0zAmc5ZTBxF1Tskw6TywVJ4uooEFezo/UY7Jmr35g/Q5PplXM9
UFfg7vJhg8l7ZuoiFnida1p8AB3w2k56IDC0jYNSYg+h05ku30K25hlChtdXmgXt
WeVJFSnDMG+krxqTaFXxQgU5Lw9KvIYvzeCJLHIhZOBRc2To4YSLU/SQG8NMvde1
L2M1PNODpJBmmRfDBjbrCV3V3Cg9JuYaH3TF1kSfVih8RkbY+ATZ9W8sTO+rZgrS
yKrzK1jgeLDMPllSGiay7GdW/AwxcI2j5zo8+58QKh3zGQPCuc6spo7a7DbduG0z
cmdNjK4SsnRkCfmTzUmoGgm/7E6XvgibgVDnp6ogsy0zECE/sx2G9FL0xzLBskhU
FVRdKLlPCPO+ojARZaDKCTyOcFjxhrDLIlsIUv9nnA7P9Ml4L1pB3qLpRsN5yliG
lwPAakbfmrgXPkNnNjiiMJcI0Yaa9FIKKiua1VljLz/O48pdI5wikg39CMBcOF85
otL5nTU3P2JcdUtTlcDpf8eMZh0zzBL7idWlSi/J/7pyPByv+BOdXYsb6uF2awug
kMVKGKSneMb9CK2VyKwjlLVeiM8W/MCDc+zjoL2ynDq5YkWJ5Ag2x5w/orvQJ+Oa
GEc96YilpBOlE5tjDKa5edPfYfCttcMAh4aU/eymgrfaaSjP0MZFZZ/F6+IUUT4e
wfOkoZDhe8qblDLj5LADZ/kfmH5AzDsSrw8xxFUrBtDJmhHvr7tbUMrw+kFwrX6T
cKkCh3VkTp6b+jdnDbhZDFPANwYe9Feyo7ZzAeiWRhrO0MMaxDrR/2QDi9K9TNfG
ZQ5fxOQLeIxwAZuluG4YPk23yuFK2TCxAZxsWmtq3phXBcnl7IR+Y8qJEBHAD05T
V//p+bHc5mVc9A0dspL0vthyraKb856ISmBELMqTRQK7MOTU1LWde9fO6k/1hAGM
Z/sZvRDHACibE4IiAUqVgyOEmvTdJaKdkPmiyFU+NEeQWLpP7uPCt9E37CEuKH1d
Sxr+NCo7hyBQOP6V7qFEqVyvP2tYA0LumcOPBDJDZ9DNN3iF+48v/v7SBnzkeaEU
ztWgVklwa0j9hX3iX7FX629FcgT1dbguGn4BTPRH1wQ3x+U9N3bU/VumFnn2ZZcL
lttQadNShZ5Kg+HSdx82l1SyIoXCrdkqFNBKLRr3kI10gLQ21leF8sjG8+uhhV0y
VdOj6BFV/lbT2VrpvPDGuDSUNqykrRcN7zDPRjYYoNTLGj5tFerJ4cGdNkC4xpot
EH++ERFkbpVPLKB8z/A/YxcswLTVMtKWy8LqU+9ZtMDmvFsrEfPEPEzagGZKnvzc
9FYhGdZABy/yNwgbN5TUnpUt2J+8iIK+R+P00vaKTzjYIacpq6ecEaah3UeHpOoS
rxeJAGUgVCQuQPCer8r/kdqzU5tMjIRoqECdYV4LKPSS7OEr2SWG2mkROba70rEG
nUe+wGh8C4Hm6lU27ZZ4bl3n3L26lEj0eKv+lGbTwz2UnfC0vjU+vqzDxv+CzSIZ
u4ct+gwekemV3v9FKoeDUc/S+kYN0AQNv9zonNjfbpsRoGUg5AdJKHpt9NjVDEXU
1fNqu74VezJ7pYuQAwDrwom+aSVcyA8NUlwbEZChHYJf2VQhnbdfihip27h7hnPA
UNrZxNs85xcE/PXvQ/257WaoYc7hAsRbP2JsJi3PdassQ3RIe644EfXXhKh8runE
lUFs53OijX3LZXZ9hXW2jZMTIqhn/IZb/vqcm2bqY9Qg7uxDsgEzc2V7zLUfXtWD
0M/oon+IXszzSXdOOz6LSw9rVohZ+Dtnn4P7cBh03jKqDPhGLT7W0qykDAYTTKVB
TgVdGWVBFLn7d4pg9W00nNs2/Bqw0yx9OpUMR/QgXmtd8euN64UezpBrYgj3KUxP
JLUKjnhGAiHh6nNbYCEVmG8NnaBz517XMDCP/SfE3++MqY0vKY8DeONMGRcifR7A
M+/kybM/oFS+CMa46sYvsrAUaPQ2k+6QFLTaszqM4Rlt7KH3tddNoZwRBKqOKXO8
l8tsHty9fnB6GE5NLV2uDRn+0WZtumWDBC38Y1MlZmHRMUK05Y3xXL4HqAlyf0ws
kZQePk+oEb0O4UWdoZp89fh0u6ErCWb2AAHsBfTMChCEbZ6WbccwDyL+T1P62hiP
TqoZcvuYOv4QrWJrUsUw5UdJS0oD0E5+RIvqT2rOZAuJqWG/ZNLs9AskAGOr4UXA
cqDZurVTl0JXqCp/E9sHhrNLAIdSvkDcaqB0fx7XH5ZAkh0cx6MX3pf7/myomNgw
RfYt8P4lxBNbDqYm2thjWELxGPhO3K88STZq2OuqvL9jgo05p/8RSs3akyQ5iWhS
ye6ODK4NbJx04N1q/KBe1yqzYL7QfMfm+5wzngYc8Fi9INEOj92HjzW4OYhQjrdc
OCnN3tclsodws2+AVo8Zl6wlDs+CzkmdP3ztISBw2/jtBWllQzh8ebQiPKRATzzA
mMiUfwuPqKjzrE49pXbSkf+bbCDGYgYn7xpDuroEn9sx7aFkpFBYfNTOWd+fT2JR
MOss8GdnrYS38V0T55hfQ8YxvDKJXWJt6+hVdN+8tBNa/KhTrV4WMkWWrKEK17dP
uwIQym0/S+gxzCslV6PLrhTzY3Y2+xC30x3MhNWHWTIR4K9pjvl9JWs4SMhLmVxT
aA92cacPpRIiscm3566cZ6aNgQ+DvaQEMJVLWNLVF0VD2GEJuCTW5S40cIZT+PVm
GRXF7D+rVdQuXCxSeJqFt7qaBSdhG6sDxVjGdyPzXCHLxyXde08RY4Vqefaj8Q+V
YL7Ldee1GERhGaWYibv6q007lS/0V+MTbxXd5NeX3JY6OW8ljTCAsXPQKv1h111A
IOYR49SUVd+8jZUCLxpFXvsG6M+gV0hOy0uD6AaJu7vVngX8MyZoHJc7NnaH+Mu6
vWOAglc2fvRh8Ot+Ip/d+aRGyYDNLg4GRSBviQ3+8i+ATA3MdAhILlgVx4hz15a1
YboVBIOvog646HzwQzc+i6Cy1H8UsxTI8LwjLKwGLheAFfnVUxhJTdZKxz/ywnVv
gqFTHPsuruG9BagmlmQz7rvjyKAQLSQ+UiPPFgKuYJeckd6Oqh1ZzJTBhY92+99T
eOoa8oce0rMTYq/EzQtD2YSzlr/FRazpqU/guXqVNWv9YSC+3iNtBy3omJE6vgn/
osMjf5toxa5567PBX/X+dWvgUJApr/qc7gU8ee2wOAh/3iFB9a3/nRohcr7RxkMa
Q6NQOEQ4l/ubVktLI3xa+BzO8tUaT2maw+RURWGFR2NbTjB0rsTMrxai+NqtOxnS
0BBJkpe+/HVT6Qdsw+DGbNCl1AhTfX1l0tbOheoNsF39TDklbpbT3C1UqYX00Szu
usQSGtE05vkjF3sDGgpXMzCE2XO1vjmgUbr0sKb3XVFMDk5opD1SSECpa1iEtI/R
7QJQ8GOyfgMMbYYtFPsbLnDSEaG84PwU4PaKy26iNU5TOjycBVCj5laVa/qH7Qvc
PZ/Cd2s5LTaahNqa8LGiWP/ErVtRgcxs00zHzi13Glvyl+wZfcwUQAN6zqKmAiQd
W5HO4uXecGXu73996BXJY266b7YZQXuuG3YI+kNHWXM/IpiHaltNAJoRGeCir4tU
bFwt7+3hfFAk3uLLb/Ou/3m8FJOgpcDnQNAtRI4igMx3Q3O75GivB2R6Yvb/NuW6
0mUrOWblkQlH+qsGxxYnpo1XvBJMA3aVITRg8KeKz/SFPwAARu1JZPSMwerC3eY2
69IY43mkuWtwuC+tabxdZySqncfv6T4HM/cFNhz97cdyJlultMt6z00ognma1j+r
VnUcTk4RCv2AREwKG03FtVISJzF2wd7Frj692q+NUim4zghzHi9pMGDcxw2FAYy/
AwygCPu2ZChTNX1LQoXjWDw2LnCFL7Wfsnyp2fnzPuB6Wf8ZNq1BnDxnDtKGc6NY
jXAQda5AJYz4LPoZK1jwagcB1FV0MAO3ApSv5x9V4x42fEqDIcyri759vWF3DfZX
J45ZTtRRKWTdSJbcx8na4wBBP7bZN77aEAybZSmEHT8Jd8U51q6IXoGcTXErCLGG
7Z52TyGPqM1mT9XO6HGxQPTRQwDVko60Pe0Cg1QQcVYWw9afzJHUV6aH+iBSUeeD
eUDUcENo6Bni5SZDfhXeqwIBOGHn6VRCr4feRnlv9+PXXbQHszpTvQoNVQKbfMIO
wnvqS1Ti8QQu9fdV9eMZiSf2k4ZJZYxIYGaMOQ0BDAn6Le0xfZs+a4Pjr0PmsOD4
BM0rKU4xFIpUcEhEju3SOXc4C8LtdYwNCBJbNbtHVfV6ELv1pTpFrVeKpoDCb50r
Ct28AvVvUMPF9m8thRelSKE5+fd6HboSsbdVIorhhxiD5cr3gxKIetvzFILrmbzb
WAmZQOv83mAfZG84SdgUygV2ONvhR99hAO9uLZX8+sIvwBPbGkBSJHszFxdJj8rf
g72jVAOdbEcerGn2o8aEiAmun9vwpR2RtFNJyzl22EzVgIdmMzv/z59aWCaX6XzH
YuF9xWafZN3ErQBbv0Zn49JgQvJ7IdyiKm1HSUELB4LsBBZasvoF97iwsN+PGqPR
AHqwnZYPwLk5zFNZCuS7+ArXQ7HqpUV1+Si6giYipGn1o7rqbR+XL5c8v5ujMYjA
R/eCD1/rJeK4O7uSQcCceN/Rdt8lxyyM1IyjSU5fVIBQg3BmEtleFI8PnKoDScij
RToJKdVFNp7NiJUrfR0NJL5CGqiPE9j70r2mC2UukUxwu4xxKqu6ERuMRq5qG2gc
9JXELIJGp6zpZEZFx1xt8c6mEaD7gTnbn3nc1KT+R0dHYJJU1KXhfwxa0+Dsy5uz
STLlPFUOER064POdTOFuVD5ETfGkK/d6WnyDIBRr5vvtBbwCVUQojJ0OY+xUzgaM
BM+OGYvyARIJCFrZa5VgRg5G1hGDU3Pim70nZENb6sv6ngaw/n1xJvGnr+YLQ7U9
ecu5Niz/6rty6NGGIgme2+ESAP98kDPO8RF/rAE0tgj0iQbFIpPMIUS0/nP4/UAy
uSd72rz6NY79j+d5PeSep/BgjLnFvV/BV39sQAraHAYdLnKaLepgYtsdyY0ANtfR
llirw2EU4jWP9ZeFCBDeZPd5xDnPf2BHW0au4NIK7pDlX9yeaUnwF/PWmNRpvFdz
dGIJun0A+iGv6iY7VR1oqM8gu/D8c+AwA6tPcdpU5SB0bKxf4tVN/UrtvsaP80Sv
Li7MYuIAa2/8He9+/J9Q7+FWGrZMZFmuSatCxKo+sdWX1DtAWfNIu/LyvMOe52tJ
S8TeURgPfGEC7v5penylsY4gSZ9cO/x1hT3HsAGy5MEibSa3kFEElRWvfT7OnVDK
1c+nMN2Fk+SIdcIjbocBy9PlpjPG9+ZuqZtd27k+4h3YMOaelNdCWiEXDRMUtrFu
PYiVrdRYyj61FhxC428xW8bai3lqv9s6oTYt3f7mU9XnzwzigwSVh0pAnSf0eCiW
o/3rIR5J0OWU3RqTxkFGZ4EEC7tku4QkyqA1Kqsfsd2AbTaQBtBjZAURfEdQd3M6
yBDuXflQw3ICJllbsP2gm0xPIByIFqCVVbgqv89SLjAM0JK2AhmPKDHfwpi3pHPh
6WuOJovomj6S5/uvyQtKeXSMJQzinEgZG/UNIlZNkYy9av238yfW5hHuhC0vav07
kwnBpz48x/7jf0Btr3bXmUrrCbmQGYBG/vzxCcizyOzf+Y/G/YvCr+h7TaCm1rSA
Q8aCZVe3nvwGDaF1gOsJfiDwHZQzy7qL3gAse5HBpLb4BEBZIfGmxTnyTkhcSEyK
aUtVoxZqqfgPCswASG1Alv0YBHEwJAgbcS6P2cTOG5Nytb6YYEpYxQ+GGCszfgQU
6QQn+TfjNf6B61FgFPtIWxLR+y95pcHDRGMiFO8RP7pI0Z7qxgLo0jYvuXwxDmED
4BGW0ysXBb5BCl/uTG/weEuwWOB81M6CgR3ttMF0AntAyu53p+8Df72jacwm/JFR
InTbjUul/2tEPZU/GJ8h2RqsmbYmn+XPr0fK6pYIuQokSvSjzJhBB7A8Z4Vsjwi9
DvIbH5nYxSyBtA61zz3cHI3ai/geVHNfaeW6QHsSMDl0gtiSww34lS0gGK9Hp4AD
NVYR7HvmpuqqvkWqwEzBvJKvyy4V2cpA4fHSDlhWmKUZAfVuaRsqBu9s5O+Wmgzy
WmGgESuBV4GMdelDvKp257DhPzTW5djxf50HsgGK2rvAacK9sjWCTbMkJ8qZKpOH
0w7pOwVVd46JiHGyIl2mMuk+toqZwPl2jfBtnKR66uBJ4wrkcnpuAQdGVPjWDvOk
lwm0UjDJZsCpAlY8hbC8M/YqrfdZK/ddRH0jl2PMMlJdEbYaJaAe7DzYIiF3/NCL
F2Nr7tPepSC5lk33/hb0YxUIK4iSDjmdepkNieXgWoNaPmQhRBWX3fY15aj+5s21
vUUr7bMcHmtXN9fVTfHMVW6mizYwz5NJYteB8veL+yBSNUrs1StlqycBhXugTRNT
P4qWFfuLVnzR69Y5emmYpzLbvFEbqD0SDChNO8zcqcSFBDX6HEVOQXnQg+2KnFC7
CsgOLI+gTOjrl5oMOj2ziDMaKhI1fDV8PzL6HoOhF6FP/Mg1CjVBPb3thz393qNM
uLkZXnAeMJLlXIBRdox+rszV9Wr7jEVdCuIhvKebo4YXH1To1kRt0KynaTgImoNu
jd17MvwaV0wA89M2ATZ6LMQnqNAQCCPgxhS4J7si6Qw9THGuJNl1wylcRaWQSHY+
NJoiWfEm6Zh/WtGBSSIIjb7zPRTvmM9ST/7cUF28pd3uTdkak1ttBaed84b9ooHQ
Jw8FYhol3Y38WN47X9tfC7+8qP6kE28TNzrOb070YQtSaPl2PpLkcNR1Q0mpkHxy
mBPvzL6924kxtuMc1fryBgNZEBk0gj4D/HA4E1Ym221PDPr8jnHw8/+krvDDEvTI
Q1E2ed7A+6IEL9bvEzGVqe2ZcoTU6cXDF6f5LXxWDfNns14HZxjW83i8dZ61OIHM
l2lDOsI/xUwERvw0RKfLUsINrFNB+Ntsii6n605neHkPLOySRH7FCSrkXea7iigk
mWs8A1ayCJkI012dxcMpP/4E7reRNvSkSbDvDdNFPVVJNdO+B1dqhNbrgwYfRMCQ
89QB1nIDg2WIglHaDaRAo8tdllgrcVSxfXysvqMbKPx2j03im0jU/7okNupRPCRP
7ZaISFg5MvZkM6GcizQT+1FOvckzp5J8TeqQt+nCbv0j5TSzFVKC/FV78Gwn0ec9
9KdJCHzkZ6tFy507aXvXoNhZV2A2iNRKysridN4EGNE2Kp0IQvX3+8MoOY3Fk7la
niKfdE6JiG6mFE7K8k7sWYldkjG2NaPhCIAg5vbs3hjnuHFKek6xwKfDrVSUHu3v
Vc/ocjMcBAx/Y7/W0wsJJ755Ab9mu/BXfo46aF2bpFjvw7jziUaGm0y3bjW91o9d
PMfBfOrpOkGQm6CqO9i4CW+Rxv9uIM1nU5uRjE4bOTwPc1U635e2NYCWd6Mzld0c
hFl/H4xD0DOTlAW+TF+fe+ujWLej7OqaL3Izyts25o1ZwgkeD6+uD0fRXCthdU6n
ESnoDri3TEiVd5lHKzjAFqxOKJZCxrSlrWOb9yx+wyOkx8X8EcKsc0zcAjZ6Z/1n
GerVTCqEUruvOA96U1A5KAkNGILPadVONPLZa1NK18Ol3S90g302MXUO3MhNFPQT
TeuqVugYgMDH+3JZLcy7ou1C6XfBNvfCBYJuPcNvZyVI7QvkXPhcmbH5+ivXIjJB
QtrZgSqW7ntY5003vF7JuRMV3CM34I7SCMESmpw+uIY04aYGRCUGk5BF5W4aJq7A
/SluAfSVdGRGCkJ/vPCyTV7v37Cl9+rUCuvByR8JCl5Wl2t+3bmn6fXqF6VcM7C1
8vcW5Nqwgeca0VxNIrh7cNdk5/db6ljS67l38hC4D9n8MaWLe4XHs/vL3mduiCvE
ezHN9MNUpsVygb8FL+R/CHfHJZ7en9A4FB2EV2aYUebgtE0IIF9MasXqteLPa5PM
szCuYxuRowrcRe0p6vGywAzsq942Q9jH+67AG2nlDzB/Xk6nDJMTNxjld+mKPxCC
6pCkJDexIseNUYq4h/eAOxbeFInFAbWS0BdeU9SXnG+t/wjoBxjDYVjYMWnd1ywy
/MLLxTiqG01JfXMKsOxQ46AXe5ZRrH8khuIZgybRhMn1feQY20Mr9viPoZRW9LWc
ww22LPEsSxALndPKfKGgr6/Q0A8mT5+O5920RDLafFapTi7tT8Q36/lCcTxLApQq
2Qq2Eox5CflkaeeNFtMPwHJvwSZZgGjWiDNyPkao14X4D8Urw7BSOStVx47Uj3Nf
CZr/YdgaTXumEu4hEj6S6UEA37TV6g3brh1EReSjRZ/tDa/3mkZe1n5oTBsA8gjW
4MPDXX+QT+hTHxWGqmuzF+iYHrgXhxGqIuKdt6C6J0SCFdcaIXRk1NxBkDC6Hhfm
G+Eow3OtJL97aGH0bZbm5R0Q2VAcJ9KKO0uBhoJw0S/RsVveh22qyJW7cPr74UAx
UlBWjK4AsHcioJc5+cwo3SwkiLEfGaIw5TFOmOC8yaBx4FYOo/HFi9+CqVBotcid
Qg3gSxowbGhPEFUYrBZsyoNkCgYq12g+NYubsjyfLYtOX/mNemi+bMZ9Ucebh2sM
geLhIxcd67qZ0t8Maj000/iM/FaosL28UkPpdG56KigD1g3epdijHuwvVgN1ad4l
vURtLzUuamMgWKZFGj/WgtfdsJ8dn2OC/6pp7/HK/03c4gmAKKy18D08joxqzhAT
0P3CgbuiCu57ettp8hxWPGN0wdYeG+Z7nlEgyBgCelAT4PtIidAyjm5sf35VNybm
H/BjY/fYVJgBvHRIqXDyFgKBEDUVvJ6lX30U+MU35sx8TvXYEyt6mQmHS38hsiw1
zh0UBhWupdT3AfxW5rWxDRJOVr5H5oufZOVcOCFv8VXssW8VZEB4n0BwI8wnEeui
yDZQ0xRXbtvMevKsrxMAwGBjWjZcM1WD3Fwj+9/W++onYdPYfw1ZF5x2FOPDwSx6
ublbQiVPanKzbJB/fAeaKeDlPnBvhyELK1uIfDp4INN9eS5JiOW4WoYJz53wmYvH
OV6fgHc9Iy2ojislmLuekHVgy5oVO69R83wSbyqZ/nF+drKkw5l6S8sufZ8321as
2mtXQbgCuFmCnV1c+UwDlaQKh/TjgxhBYoRii29Pv4c2KLJdD6VyZ6axfZ9DjmYR
86VzVPeG2MVR/0CDyo/xxlmodeaIlqCFjY88lzSQV0v8BMJbE3uD5nl9lul4xZXQ
yfkR5YTrO5WI4J+gMAmZjG6XYApP5/NIWIxF7sq+bALQXsJqG9YGlMkfmQsqDzVq
23ACYtLXLm/WflO+81+vKBNnUX5kgY9F6LHRyWMInUqY4fnaFJfarncopzPEm9eV
V1BGrGZUEuC/VQK10mn//ltnZIL8OQlQIYNZvg5M++z/W2pdjbyzfpbbehEakplX
FXY9JNiikM6Xd9h27tr7nkqFheKV8x2prbYk5GanTEcopqddph5rwr2p9Z+JwBQm
W4MxBK9oUupGckPOTM2BoLj9fJ/jd7qawmrwY3hyqFHSCpewaog5++kqDStEmhO6
IojDYNjpZ0rwlT4tJlMsZ07ohnYhl8tvIjFoTmiZc8oS6q95X3PxdyQRqJEALAfL
qygUxRlMfYd1/W6fAYB8fTEhyuwTsNxW/VLP/G3LpLHHflu4q4T1RTlr6ETz20zi
xS4Ha/dMB5xA1mmRYtO0BpEQOhFNgiOKTtd/lplBg8DJXVHD7NUwtpIUtIPu7fWI
M1dq+UZ9fWBi3r8wnAa0l7LY/R47UmNzxs9a0gr5UDrwvjNx+srAXjPBYqoWgsXZ
pG3Z+n3chR4OftrsIjKR+3voBsPkJ9Eb4xXQMajry3HaNGsFdBtCfuItnymNGl4Z
noS34rsO3JGOdQU3IxkbQrieiAje09u0JVQvCt/BZmtALMk1BTZMo7hvU7SUe/35
jVHeg9mwJ/7j+/qmXV1Rlqc2NZ9Pxt6Vj0kOoFeXRcwygumC70j96SaDiopG7cVf
20G1tm0m05DxZzyum1+2sXUEQ7gcWkKk4CiopHQHHf4f2tHwmOLDzPt/967rfR7T
2oP0bMvn5ZOYBTasPaves1p7frU2j7rQfvny/Xz8r3UgeDYPJv32ztWJ5hKLDK8l
+WmWobYteIHxsQUtdSAXwUjUFrfNt5Uy+dX4OST/zqQn6qe8uu/nxDG/b5Vl5x2q
mMhFCScyiQW03x89ZYi53oIR13NX4Lr2dZc69AgkR5VEOdl/MYhrwSDcVMThOHW/
wtXdqscEPNvdWPgDMcQW2Vp/fQEVZtUa9oe3DFl9ORelqsrjyyiM/O+m2d9L/rqN
ZRWbvMR77ha/cULu2KIjmbZxsYB1Pqqn6ivd9xq79OhmRtsgPMOTHc22xsK0J/3m
Mj6n1HYokeuhDu41OfiiMd1BZbzg2M/lxc/8HpfyZK6DUy/eyzIU7Iis9chstHzh
v69hA/ZmZ1avcS6I0TeVqnD49VESDUopalGoEVkDKScHMFJLekQnHy9rl6WpBcao
N5jN+nTdyfH6r+trdPkawiaMrxOBQ16TopPfHS6Mv3DdgcIHKO3pLiokj2tgV5xC
fgRzthDjTkD0Wpn8dTGw5CQx15NAPe/fXujOsINbl2Og6KD+p7z6FUtXEi4pp3cK
9i15CL2JFvyq3GUW1Zgd9GV54SMIx8DU0CMitN6zC+JCZjCkCgiHDzx4WHio4aRk
lfdTdf/lx0XNRd9zudF5/YgUTH08NHuoN1D9cPibwYRBoyhY7du/09D5IUzmnVo1
3yUA9rJFKet4Rdmt2335QJYlEeW73rdPNOps2S7zPOMgS5nnuedZZNFzNpyF6KRp
v3qWWPZY7kLEcY9rpdZUmUi93e6KyMHDbuQa6xrW7dS2r0oqywiTFrw/w00xy3n2
sSUNtYJrNhcVLXFwruKe4izxnKtn9Cw4quwOZNDdI2ZgJLfSY8OSt2kDbWHK1X6V
l8krpgdFw92q9nDmKDBX0Y+ZEVeMEqg/iXbRn294K6DPG7k0Ts/uSZZj4mtFGxaU
BGM/0HnX+U+zea9ElGf5qu+r/i8ZcQUedGNCau7QY5GiLFgzEIUhLI2O9EJTuIR1
43h5qOiQz8UBLSmZAPqhocWBvi0pQT8nuEtmHgRytRbDonLusKwL4bYwtBdh3cE7
LdUvmZ7hsB36OoNVojqnpEJOR+CSFJOPqvSXZ+6hCmHqhmVNbwl6GvkBZR5+bH8b
ltkuuVAfYR7ncnWwfDOv/ydldkrOh8J1aZfM5xlJ3DoU3x+30a9uO89jrfyt3rfB
Eqix0lY25MkRbF+4zgX1fbxZNEZMoHCLnYCYkhLahsmvMkEmwFoJ79pKNfiSZbEU
ha+AHjPuOw37yxWQht7UXIfc4zPXfM393YvZL8qj+mwEnrnZrD9O3d/T5lPPdQQV
zq3GXliYaM1gViNECO2wfgc61NeU8J3fAvmXgCb4CaWoItcRVAjUQwcK909ERXVx
HZrRjIskuz5zwqH7sRLvP2Z3QjuHalUPYADl/9x/SeQPKpTY3Os3kbrUFGAxVuy3
DP0lxZYL8mrw9ojUwrstBZon0UBQsWyQH9+9HrZqktHwzh15mdqWXKw9y1UfhMp9
uGmypAwVrLtklsIbdPZhg674gV+5FqltlmNuEfR9B8ld+Cb4/VcGcegHLVjE8yV1
Z1fJmPv16etyDwdpTYqWU79U0PabvZrj+JtHQmQ3T65dSIORr1V3OtY5gT9xXpCS
ZSp4FEpUhnkluyVQ2z6tByc/I6NeHnsOS06Kvn+x1T3GMaYYhq4Pz6it5Ouqh5Xf
gnae3CdPmetPf36bslWS0Tx2Nl4kLTr5nN0HaDuAzgrlnFvKhgXcfFl12/wVbgsl
rbHlBwFqPWcjc0JLh4qa8nCH/WlQ9BxVFgX5uLAV/pwxiPRmDGtC3lkC3PO1gcDd
iD3/2E6qC0yfPU/wssJwftvGK1IOdQBTql3G6mZKDVYeMDG+nWnZ2m2jmdy2Kkiu
9+RJlZ7vVI0LHBHLPhLAvJ1hAgKxN0O3EGpFdIEEi3/waiPwro8vdO1/AE39BvPU
o11qIRAFSvoFRQ5iiGYNcq5xwS/rqxckIqElVb6yxbySjGc6JmsqzTit4nMQjy4r
Y4XUxyXV8wFa7UFocEfMvTQ7zs6aUFpYAgrkeTIkP4KBlMgTlRNxBUBmNAywVwAe
NtrL5ZfXpBBK4FhwtNqvefERWaVJVmgUqCMbSVEX+C3cOuyCnQ2b0ZeLUGw/D+qq
ur3cYXdSm7dpPzYNzo80yO/tPTAiXHTCvrtyXhsYvdd5Xq8fE8y5vxvERddycw0r
X/+rQBHCl3vCIDNM9uUDvUOMnS19sAgnl27fArYnozs8PNkHwqVBdnAloxSB1742
FZwDereqvo/sZsLsTYBZvBHuREsnl31DUN2JGRknWsL2akZVQlHp8kxt/V3CxixB
DyKa4y5sxsEgvJ+kBMIxlJnuNGyR9FkRQhC8BwYy0YRBPphEwXDfpdZ+LZy3p0Lk
7lzLsKy8bmkZDBWXzUgSRQjTZn9yWLjbh6+KiX1OxHyqVzBONb47TbL9SaatJfD1
pCTbCgq2dfVarKk0CfSEUjGO4s727Kl8PwtMFvdtWlvMEUCE59/f4O6ChrgfNetq
gtsCxQe0fr0ZaC2qxj2oQ4po6avAXuJ3YiKcmRqM6EtURtbxSxsCKnbzYnYJ40c1
9Yaj+0MWkrKrPWv6rrFAswtGUjUS2Mm/4hhvQ2vp5TDTuKtfts/RO4U2l1+QhRPJ
1H2hJoa/JsIb0yGyV/jiCIeh7zW0GrGOiAGk5dKoXFlCeBh4B2C17vS6FeTCdORl
gxn44iXq3II4XHIQjETTUM1L3ZmrmZC+FoPNNsYDAnwERTRHyEW3PwQxyS/GiAMz
ypYX7VN3C0jX4yTSUAY+UeLainaLvY+5UTWQ7/0fd9/wltdYd/AR+P9+HIdfxDJY
8K2Q3cVxKoiyqatbHHaxvb1+Qm0wY6AT8djas5/LXYUJ9O98fWjCS3L/QwU/Y2AT
3owKL38RutJENTQPmGZIokfpAhSvkyT7sYA2xvOJghj6NdWhcesPneFyVbZxzOIV
MD/J+273Ftd+8B9wMyqTrxFhJun7Bbgo+9xJoJFy51hCbgAo7aqs2HBaPS7yun7O
rtMuOwJsfHN3JNXb6ijr/XYQzgvwGThBYWczxNi3UbOTMMKA8HvCc3IFZXiKRAAT
NEUMEFytYda4rs5A+iZyTHpo8UQHMHMw+mXLTdgAz6vtnaD1W0B6v//6+5z/YR1b
6YDNx7boYZyRTwSsxmvpTaaBw4b7OqKQ/3YqBVFsB+dzsdAGWzpepRWWdWQxhvWL
kgZdmZa0Txxe1FyD8iuGBDjuLPLaWZSLtb9TUtcN16DyZHbvTiRK33XzRd9Ajpht
wLerYxIBDIjxVNA176hrauRyMtNx0205xeZ12/2DZc6HefeMucFeaq7MwS8fcZW/
1y9N08+nMM0UMc0mNmtcgGALBN4M5d4hBHQInUoZlngFob9E5TQeGzpdW90evsmK
WOAk1slicBswKwA+ZR7yVPGYjJfaI7FyUBvFpP9FOYcgoeTcH2o8ll+d6fUG4EEt
IBdXd9nmmqsccI9N2TUGhIxQF4/julTRsRgbVDF3JHWo0OCAduR3R8wAcgd1MCZW
gY0Cbv/qgDHzNC0cW4YiiHtuswOtYlyPbLJNc0+SYeILbsZm4k/GNsqEgzKi+A2J
zkw9lMjRIgMWZ+yQsQSRczkjEnLmthQRXypAsmuqXwmzgla/kgl41QonggBLPWHj
SH9tr3drBJt9oeTYzVjQrqPigF066Rr8iY43/PrgA3rmgJoW+mDjd257b6gLxpip
M2S7O+oQ4ujq+7rti7rHOHW8CaCU8IzJ8naJgeesqiIAd04pOytKG8CFskyCA+Ay
JOBUqxe2Mxh8DmtRubSniZdam1aOqzmzd3dSVLylNu4BTCDAzKrejUOUXUqtbE5a
2kgQoe3Kk3/tvzwPoX0MW98j07L56hRl/e6wrcNpgAkXmFUxh25zdMzgoauYJLWj
hnEbSGGTi4yLwQp/3aZch/2rFC+sFIbit3G4WLWrUSqu1p0Buv7j5ejh8PTSYTYf
RHDuzE5iF/24pTL1K0v7wjY2z5Xj7BPisoDsvQhjXcBlEfms21HxwE5U+XGz1isB
kVRzhs5GZfdk/k/67txMhDah+ay92f0PH0vzWKuk6qn4sFGl9h0gA7XlQ6yZzAqg
CCYDM1Y7KHS6VBOR+JB98roQg0yAIElS6vw1fyvMJLWV1bwyHZ5tBGG+VKPVO+Ez
C1Q1OxLV4jNqgiGXX1SXIpAuzaqZI3OxS92eMpj0YlHWdmxWsPswWfnIhso7hEs5
f5QZV3TXSKSMqoli3ulhTTMsInmnm+MviviWjSfA5GZ5jevFl93+Av2vIEbOb4A8
z5bJ3z5BhPxzxwTdzu2ddT5AmZGHJ1AL+SBdeKEJzEb7q33fOTAAHq7ftfBP/vDf
HPQU7mfpeUVzdwh9xQRaWbqBypcPnsgPE5pMcYgfE6OGYr+RZEkdxSx6LloYPv9M
/H1NgJdLaIh4avmRjJACW2YeYPIuv+wEhs2Cm1MX7odFkbhmZhgFg+65yAyMh73D
rbeLsjkR9DaSWJDWn8gF6eS9cP7xeYXoB9pr6L/jlLhiXYvgm7O9vorfLjJGMkKU
FlV3Ha3e7rkz2v2XlRF729p8ty/w556CVOfMSgiMz0QxZIsmt1iKhOAu4RVl+R1s
bkRm77irsiiZCnmY988Oa9Hv19Fno1EVKcud+2XXrYpR7vjJ0mQlqNl62AMu171U
yNd1NLA8DNfomcQC+k5uYuu3DEUvGyxSKabxVxLYMHhNg5L51QdUwxaGVk60wEEb
FluZNm/p40GqDzHcElEp99BPmN2+xjA9Aa8Pp5T8Byc3TIhdQJHXpVpUAgRELy9V
ovYEpzmLWApIhH52ldGtv5iPYxkiVlL9RMsfT1FOS1ytjLDNBO+U1OqGltkgxW42
MbSYBj+0rvwt/VY1ogAMYQYra8NVPC6mj9rQGM7sJi0bSCXsayFum6vApxUb0eR+
TE7ML/kkTM5I6efP8BDIXkwm8M3a54EvtcOhBj/joVYeMmpArhi1vVoEhyEq0P2X
H+A+QZOoXxrnfDu3+HmceiFQUfP1nZe4Dd6hhH5VZuqqZgQJ7mBwTQ9BKus3rWvs
lvf2FiSjqwcA3yL+Y/FmjEvaYpap8EhX4Krujcm0Onfv8psa6lLDuYO2kHx9bnuy
+qAk641osmJAXx3EMxXKBbReU3ruBsZ3DtF+u4Y+6EvH3h8diIVCHrEIi9NEDZ1k
Ulp4f7IKYjKByN/hF49u80PhPc4uXh2O8nQ1G3ZRSuR9nOaaR+3tMC7kQxDs4F8c
9fPB0WJFrPMH1C1z8xJwSM4zRzFA/5fhoPDkZDZ0mwNUQ2JjsG3xo/rb4VD2juyn
f+q09iIK51UudURWQs1Y82YgBwHujIz6WcsNvPttTN3LQeACcyGqF/SMs5uowCWq
CTkld5hx3oZTGHRB9vbq7HR7NqnYGOyDR6dT67sXOKyqF6J04enY8S4oHS1Ssc6o
gVLqcPJrYw1oGKQU6nhCNBYXYsGi6IuYYB0iT5VFvrJbdbogGd/8pEDuIduidtOB
ElaFL/jCBmh23i57ztOWVhAbxNF1VaN6dNIIr042EHYkQDzakcNDmxDojFwEGgon
HExYKZJ8wmYL+zDCD7gBGzMU+4T/hv2H/7LdoyC0o4MN175ThGjyLOz/N4u6qTmv
2x+i9O+RWkwdq54JHTx31A7gPtPSoRD3EhhB9bTpEqhFsw1t7FT19PYGMmPyRFEY
EYf8RAjjaRaW41J9rY/oH5gI3tFIR1JphyRYtOhfvJbFm5A27QlVOLfYlTeBso1w
KO9MNirHjd0u3hd3xDfQpnW/JOPgHqRCm8JEoQ6Rmjvvf6DmEypl4TXjbfjDqjca
eLWUHtWw8C5X0ojEbIIrEPFaCeRgsipnd3ZxY7xDWPoplqFKEh5IYeeGCs+/Uqvb
YIqREHhONJ61hCtgRynKvTZA62E6HkwDHqro7YvkgQnkkqF81HDnaaIrpCk9B7Lw
HtZHhw9rWWUgETaqu609uGJc5WDnkJ033Uj5X3ZpvsutYSc1CMWcH1SUUDQJTYJH
l+Ph/990h1M2bOQJ0woUPzez4F6OaVrz+BPmRlsvu1SuUSGyuDie00m4zk6nMkSv
/b2ODrZ365Y68F97J8Kmk24nFT5iI08EQIhyFeBazRqyKuo6ejC4iNe1EA/RcIKr
gtibYOcVzcZn7ZBMzrHP3EuNzdAKaOCMq54Pb3uZb1SMFIqVJZU3YVwaFXGGHyvc
VSzoc8ayT4JcK20S9IM1vNtNDE24VWiqEjTfmDPSX3W7T8yHa1WwteFKL4/1VDB2
OfCxoOWOFZmpr8a4zzSlAJUV8cvK7EtClE/QGyVfjM4xQiKou0EpzTQGNZG8niKV
p5VBAsnmyKb26t9OVWJMk7X4g9GmyDaBnlbNmcqZ7wQsPSdsWU48rhwiJM7VE8Z4
EeYEqf9taSBRakFkcZzWFGtTUnFp4xjOaxDx7UihsZm0mcf9YxJfevmJfQ0ehoad
HQ4EvMiaQzepP0h5Wu7a6Vb4lyN1O+cqBX0mrXrRkG/m5R/a9ShhQLCyT6EKt3dZ
lunJwzup+FD4UJ9H/YIFAyxyFpCCTI0foL2dWVbgUfYMYhuoedpMZAL0h8USIPPB
qI7FBWNqu2MKTJtVkA+gBvizvaeDeXaqmtH9Zeby0/JjQXsyh/31ZaSGg8Pk3Wvu
Y2NoeGs4h0TYpwJ7W8my3DHsffT22eih7eJxzw2AH/NFwZYsyTNY1gx5PaIIWjqf
fjzLasttlJ5mKibEGd+AQuAfOktcQM1ilsLgIta4E34pKem1btTl4qHnzCTJRYAL
Asa5e15dR4TlC3+DO1yUbyNXyTh9olA/JKmMqTwnalM4Tnd8+Oa8+87OfkNALA2+
fmePxK/t30H+1E67bTAbOi3qZbIrpQr4w0f2ehoRFP/cJaNnZKmroc2l7xCS9PQO
XbjJ6Yn7zdcLfuqpjalbOTOuixsgeN+ChMvjrATBPAZ9FYc4Z6MEXZn9z/4ZNyPl
I3m0+xrdfv64iUR99ve5T+gm5d30ZIAaiD2vpfYqiEwEX0C3xXNZ5SnWI9W2EZC9
6vhBPa3PskURszZxohQOZJ3MHxe5ZBGyo4dsZR3uTBWrFroP/6o+B0YgP/ZfEHvx
vBNGG25jAf3WmpHUY1Lg9Kxxv7YTeiU0rAONZlEp8C9WAp671rKXARJdjXmNvluP
aEvn1Y4gimS1q8FklKNJvXFKQBuM8DscLcOzTT9CubLElvRutsTFh+E90uetoBYl
yZeZEv/eMK46DSSQlaBuGyt7rq/rnN1bx/YF0OsTrJC4unGR4nW9N2lSPmNTRBT3
lEe1L635QGDRJG4MBIedPkUjjaJLYo7GEk2aYoRxZXj1BFvI19+WQ3cdun1pkTiz
2FhMs9wndG0YBSaMrIrL9ONcvjv06xJXzKMOJV5R2Ot7U0SXLEwfjoehLBZlm8e8
OCZ8tlqSIvnhA/scH41J6RSSifmMLkiBaotGd404QEpQtP0DEImSabgMIeG8v0VL
Rcyd6+Q1E2AjPFl7OWJSfBovJpHaDYAO+r9/dl6bIXlDHaW0x+S/Re0WurWIcB/0
aaRTaFTiSeXLwJKIFYxRu9zpc5N1VhM/Rs3T3lTfHG2+Ffy0JVb5FNBVHS3+gJUG
1mJWYAWhdzPnkbYIy1fy/3fxVURxKVKEP9yyuA+J57SHmVrp07MLLOX6YdclE9su
iDKwrKq5EaOMdwlCGPQabQ1unnODkJ8zuXVjWmBedUkAVNdChDuGg92XY2ZsDEih
89Pm66HTptD8I+OCjwTzEX9iICw5ywKCIO9MzRUpkk4N2RPbqZDjGTntGI/v+lGJ
62JwwG1fDtAmhpDxH+y9poN66GfbDY1n9m7J1sC86WoWRzJ9cA/EU23YsolDoEHM
oDh17nqfKDC4Fv85E1gha71zDBkXDBPLXRskJAp2yS/MGDvbuE0LmWrw+IAK5qaz
pICaPYQdIXzo9cDfBf4gOo2nlVi9drcZtsNasIze8ko9vBV5xbBMJpZ1QIApsoq0
LGsnLi9VeN8rjmbY3LHPRzQwI4ld0K7Wq7nmqNALkJJmom4r89k1llyKTgHroejB
Q3q9YJiKeBsf43ueMB/U3HZ3eOvSH6xX3SaGVDhk1yR7IiMoHpISxVYw2ZcNODl8
w196+6kxT9J8OUCo/b7iT0kT4id7ROJziumBGenRrk8racZUG//VNtXRGnJRqJXf
KJsKC0V+zYpn+2qnSF0hPCZSkENJ7gE01AmOOvJMCjDJrWiZI79e8SlLp+coPhCW
KTxrEeemc8T5rk83E2Atg5KUcwws883UZOqrDE1t3gEOndgYYaziWOiywN+HeKZx
T1arQtyS8Z5JU+saIhtOhOLoFQZYkNgW6ke6ogE9gv79hU+ugfi3ZTYk5hs4pwly
iG2j9xTPmFt6vVp6VUlmNJBZP/nKzqL+B7jdGY5gBK3CKa8Gr+h+W4g4AaTlrCbD
BIRZgb9dxZ67LRgmC+3dKCiTARaGZjGdFtwUmdfGioRGGgQ6m8PdjPFBJqLq4B4p
7NApEcmqv0S67rw/uR564MGM3LKV3aFjZr1qCvGGGC/QPhG78f8JsU9yGCzK2Usf
bToAf0bYoA0g079s3+74gt89nTYccw2G9TzLaqFR+wk5da8U4EIvqr9pdFRlXxWw
XcN651iGfQmGMcHSO38fbsiTfr+JZ//aU/Z1XquLRsMMX6WBHtANQPOeJgCvwIzR
fk+NZrWvPh4K20qM0AqBXkCPfCltxRdXRxJIu3/rxm7E0PsrfTAeg1nYA81zJTdi
3ZhO+WPdveKtpz+eEjEdZvywxFeJcVNs6Yoa7SUJsswzoLx5GDllUZsQEpwnE7jT
CAI4jZk/5cm1AbZsYlOn/1UW/DDl0SmMqxSSESKCyQOH0JE7iz/bCxAifM6ad4XX
LwOIAi66TAgpIMWUS3LybS6B8hIsgkqRgo/bX9BDTeyMyTOXqpTdsFRGtYCp9OPv
nf4kBlnURJOwuLUiKlkbibRpSIgjKacGb2LHjLuUsCxHCBOq1JLi0rxWy/IbfhoR
5u3wyvkF4scHmk/ieIe3HW9Z9UfT+neP8eiveR9aDb1M/HBuOS57CUZ+gvNaBGRb
JqW+9N8FPEQTgDeQExsYyOTbX7kimlr01AlO8Q62yvf7XyQRz6cSjdAg4LXfhx4j
Q+3QqlBmW5rkIpxn2vcoqgIn84OHe9fbexPQLDq6WN4D3dqOS02bndf2rwutUcSN
7SGJep880uAr186Qaq10xTOgOMUDhQjKPNZFXrDQNz7YpDmiZXoDpv4erpUJc01f
t4nMlpE5ja3VrtnX9SGiSbqc8GF+cjH7XTpCld5z+B/XCr3vA4q9mAXv4SIKwZrL
D7RjYWICVVTaApwgk+yIibDgPo66wVyxiLx7p/+Z6sYmAoGxtvlhADKPE6IRrj25
lz6vmS7Kn6+iGE5a49iOvA2OhaUPJfM8GKn51J36Ld/ECKsM7o6tBoDu/TjxpvHj
FKBXjT0wp6iFQIcNSH2Zk3b6jhk7bYYuK/ljFGZsx3FKCJLcm5OPOrzneCzjWHb8
01W0lRNm0gpBNMwYoKSQuc1trv5e+/g948MQ/4y3f97+nW7nDB39yhomHe4Audyp
ITrqrgMxB/UZBs4hH0m+yHGrFvnMiJQRnfp1CnvHMKmxs/KpBqC9G07gl9iafqvH
Rsy1kxk9aH/GX/d1bcnyLJiefKGnF3ZYCDUI36Wyw8D4qr+IxePM8+tIo43pIuBG
P+E67RJ25O85viFhkJgom8btGj2uXLkeFbpSGUqY1A1wj+R44hTekk6i85Z2lh/U
F78LcV7GHy4zJi2Tg17WS0Di+g1pHqYQa+CPgXrnSGQyK0e6slLCLBx/n8Yuoxkq
Y/9s5ol8xOh33vciwUEOcXJFDupEo59aGE1cQVtm9HB0Sz0p3y4chDxV6mNUWLwR
EgxfIgPrhpuKrgYuzVyCtngKGtdULupT/2Ebmi5t6ZwPOR6Evdcq+uzHpy67RZk2
qLGTV/YmTIB9BMmm+i/aRO5EB3yeysme19cqKYzSyXBign3w52qx+ugrjYL2IpCA
4lq+8a5J1PUU+Z1XYPF3799m1LHfQeS3Lh7PD3rRCJz/siNusBuwLiHfN1gr3ITt
h+IR4/kbNggtdv2ETnj2oI/DdmOoUHvi74cKzuSk879TcrBq3abtijDPaQ62kK8f
`pragma protect end_protected
`endif
`endif // GUARD_SVT_AXI_TRANSACTION_EXCEPTION_LIST_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
cF0/1lXjCFbX93HPr/pPndrdDlgXVHwm95iiqe2LCNhJmU1HAhDfZFloPczxRxKG
JvPZ6c5cj3QZMMF8t6aRjNPMp+nFEO06zzHmEq+VjvLvPdBzcAnMeEkgI47rCF4m
XGZHLKMThIGIBVehMNnnxYji2b922MKZaz94iKC61N8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 19783     )
sJ8P/xwQxY/TjKB33nz8PQPp3rAfeLrDg4kJMg+R+C9X8YaAH6baPRiADO53QT8j
1RhWYmZw9j6vRtCS0qk8EGPXW7m8N+Nnw5jq3kkhIYSiljJCbM60tJy2rsKcWBbh
`pragma protect end_protected
