
`ifndef GUARD_SVT_AHB_MASTER_ACTIVE_COMMON_SV
`define GUARD_SVT_AHB_MASTER_ACTIVE_COMMON_SV


typedef class svt_ahb_master;

/** @cond PRIVATE */
// Note:
// This macro makes sure that hwdata is not driven beyond cfg.data_width.
`define SVT_AHB_MASTER_ACTIVE_COMMON_WIDTH_BASED_HWDATA_ASSIGN(width) \
  width: begin \
    driver_mp.ahb_master_cb.hwdata[`SVT_AHB_COMMON_SHRINK_WIDTH_FOR_MAX(width)-1:0] <= beat_data[`SVT_AHB_COMMON_SHRINK_WIDTH_FOR_MAX(width)-1:0]; \
  end  

/**
 * Defines the AHB master active common code
 */
class svt_ahb_master_active_common#(type DRIVER_MP = virtual svt_ahb_master_if.svt_ahb_master_modport,
                                    type MONITOR_MP = virtual svt_ahb_master_if.svt_ahb_monitor_modport,
                                    type DEBUG_MP = virtual svt_ahb_master_if.svt_ahb_debug_modport)
  extends svt_ahb_master_common#(MONITOR_MP, DEBUG_MP);

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Virtual interface to use */
  typedef virtual svt_ahb_master_if.svt_ahb_master_async_modport AHB_MASTER_IF_ASYNC_MP;
  protected AHB_MASTER_IF_ASYNC_MP ahb_master_async_mp;

  /** Driver VIP modport */
  protected DRIVER_MP driver_mp;

  /** Flag used for handshaking between phases */
  protected bit drive_data_phase_active = 0;
  
`ifdef SVT_UVM_TECHNOLOGY
 /** Handle to the UVM Master driver */
`else
 /** Handle to the VMM Master transactor */
`endif
  protected svt_ahb_master driver;

  /**
   * Flag indicating status of tracking transaction.
   */
  protected bit has_active_data_phase_xact = 0;

  /**
   * Flag indicating if we have a preempted transaction in process.
   */
  protected bit has_preempted_xact = 0;

  /**
   * Flag indicating if IDLE_XACT is becoming preempted_xact due to
   * SPLIT/RETRY received for previous transaction.
   */
  protected bit is_idle_xact_preempted_xact = 0;

  /**
   * Handle to preempted transaction in address phase.
   * This is required as the preempted_xact is local to drive_address_phase
   * method.
   * This is needed to especially invoke start_transaction() for preempted 
   * transaction when the address phase of current single beat transaction starts.
   */
  protected svt_ahb_master_transaction global_preempted_xact;

  /**
   * Handle to preempted transaction in wait_for_bus_ownership() method.
   * This is required as the preempted_xact is local to drive_address_phase
   * method.
   * This is needed to hold the transaction of second INCR which starts at
   * WRAP boundary if the last beat of first INCR receives a Non-OKAY
   * response.
   */
  protected svt_ahb_master_transaction wait_for_grant_preempted_xact;  

  /**
   * Flag indicating if a rebuild is waiting for address phase.
   */
  protected bit has_rebuild = 0;
  
  /**
   * Stores the wrap boundary in case a rebuild is required on a WRAP type
   * transaction.
   */
  protected bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] wrap_boundary = 0;
  
  /**
   * Event signaling when the address phasde of a rebuild transaction completes.
   */
  protected event rebuild_addr_done;
  
  /**
   * Event signaling completion of transaction.
   */
  protected event data_transmission_complete;

  /** Event that indicates that its time to fetch next transaction during locked transfer. */
  event           fetch_next_xact;

  /** Event that unblocks nulling of global_preempted_xact after sampling is done in case 
   * rebuild happens with SINGLE burst type. */
  event           sampled_global_preempted_xact;  

  /** Semaphore to control access to driving hbusreq */
  protected semaphore hbusreq_update_sema;

  /** Assertion time of hbusreq */
  protected realtime hbusreq_assertion_time;

  /** Track if this is first drive to hbusreq */
  protected bit      is_first_drive_to_hbusreq_complete;

  /** Track if first assertion of hbusreq is done */
  protected bit      is_first_assertion_of_hbusreq_complete;

  /** Handle to next_req set from driver. */
  svt_ahb_master_transaction next_xact;

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
   extern function new (svt_ahb_master_configuration cfg, svt_ahb_master xactor);
`else
  /**
   * CONSTRUCTOR: Create a new common class instance
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   *
   * @param reporter UVM report object used for messaging
   */
   extern function new (svt_ahb_master_configuration cfg, `SVT_XVM(report_object) reporter, svt_ahb_master driver);
`endif


  // ****************************************************************************
  // Configuration Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /** Initializes signals to default values */
  extern virtual task async_init_signals();
  
  // ---------------------------------------------------------------------------
  /** Initializes signals to default values */
  extern virtual task initialize_signals();

  //---------------------------------------------------------------------------
  /** Drives hwdata during busy based on the configuration parameter
   * data_busy_value */
  extern virtual task drive_hwdata_during_busy();

  // ---------------------------------------------------------------------------
  /** Update flags and drive initial signal values when reset is detected */
  extern virtual task update_on_reset();

  // ---------------------------------------------------------------------------
  /** Accepts an incoming transaction for processing. */
  extern virtual task drive_xact(svt_ahb_master_transaction xact, bit invoke_start_transaction = `SVT_AHB_MASTER_INVOKE_START_TRANSACTION);

  // ---------------------------------------------------------------------------
  /** Internal method that accepts an incoming transaction for processing. */
  extern virtual task drive_xact_internal(svt_ahb_master_transaction xact, bit rebuild, bit invoke_start_transaction = `SVT_AHB_MASTER_INVOKE_START_TRANSACTION);

  /**
   * The methods asserts bus request and lock if enabled. 
   */
  extern virtual task start_transaction(svt_ahb_master_transaction xact);

  /**
   * The methods blocks until the arbiter grants this master the bus
   * This method is not called in AHB-Lite configuration
   */
  extern virtual task wait_for_bus_ownership(svt_ahb_master_transaction xact);

  //----------------------------------------------------------------------------
  /** 
   * This method is used to check whether transaction will cross the slave address boundary or not.
   * If it crosses the slave address boundary then transaction should be dropped before driving it to on the interface.
   * So this method is called before drive_address_phase method
   */
  extern virtual function void is_slave_boundary_crossed(svt_ahb_master_transaction xact, output bit drop_xact, output bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] min_byte_addr, output bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] max_byte_addr);

  // ---------------------------------------------------------------------------
  /**
   * Drives the address phase for the transaction.  This method will block until
   * the address phase is driven.
   */
  extern virtual task drive_address_phase(svt_ahb_master_transaction xact, bit rebuild, output bit is_aborted);

  // ---------------------------------------------------------------------------
  /**
   * Drives the data phase for the transaction.  This method is executed in a
   * thread and will release the drive_address_phase() method during the penultimate
   * cycle of the data phase.
   */
  extern virtual task drive_data_phase(svt_ahb_master_transaction xact);

`ifndef SVT_VMM_TECHNOLOGY
  /**
   * Transmit response to transaction.
   */
  extern virtual task send_response(svt_ahb_master_transaction xact);
`endif

  /**
   * Executes the steps necessary to complete the transaction:
   *   Completes the driver's seq_item_port handshake
   * 
   * @param xact Transaction which is ended
   * @param xact_rebuild_in_progress 
   */
  extern virtual task complete_transaction(svt_ahb_master_transaction xact, bit xact_rebuild_in_progress = 0);

  /** Drive the default values of the control signals */
  extern task drive_default_control_values();

  /** Drive the default values of the control signals */
  extern task drive_default_data_values();

  /** Drive a beat of data on the hwdata signal */
  extern task drive_write_beat_data(logic [1023:0] beat_data);

  /** Drive the address phase signals */
  extern task drive_address_phase_signals(svt_ahb_master_transaction xact, bit is_drive_along_with_busreq_assertion = 0);

  /** Ensure that the tranaction is valid and that the handle is not already being used */
  extern function void check_transaction_validity(svt_ahb_master_transaction xact);

  /** Drive hbusreq signal */
  extern task drive_hbusreq(logic hbusreq_val, svt_ahb_master_transaction xact = null);

endclass: svt_ahb_master_active_common
/** @endcond */

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
RMRq2E9FWeZCtvSPqVfnVum1IHYk3TycEpAyFnbyPX7+9D0duSaN6YOIKXrNJEG/
/298wxNPcDe7W1sgWjyWR+DziIaxj2IXIcOBJ0+mbNzhsMjigLXIbVnPahLUhTb3
lk5zwBACmIwQoTB9mMDnbYADD20ARcwGT316UZ5wgDgHkIjFFXG60A==
//pragma protect end_key_block
//pragma protect digest_block
5ntEhKUQWnSMRJj4TqTESJ4goZo=
//pragma protect end_digest_block
//pragma protect data_block
+D6WTFTFcvLSLymp0r/iHOlMoRSvmX7PGNleR1iobhfZyg705pT1/vID4OuFkJal
DSmckH1t4mWW34bJizO/WiaKJhus3Mg4OxFeGJvUr8iqk7Dt/vf+1y1BpSnJ7jN2
5haVetWc8UluTg9RCnKGfUaKb9ardhMhOdfJXkk2P83gmsOcdzoAFgFIgjoRO181
Jp3ZSInAGMwbT0XgZcfT1O98J5KszI4Ll6Ay+FcIMvtb6p6q63yPvdgemSCSOpqJ
miAI3vjR0xI6SgOVp+H1QIaqH8Ys5FnVCLatfVoNvvTbG2p25UMWmMH5BCuF80Iz
1S+3Vhiwbi8SNY+io7ScUn1PNhaUla8L0YICjwXx/TfK0Orh212JiFhXUktlRXNN
1zEIJCE14WkjPBK/emkK8iSVhyn7Z1kSke2dXiXXvlhXgyTvYn3GKmrCRN+ANxZt
0puwLn0tcOytIHLC10CwmpkdUnOgXbNf6vWYz48CXLonzjLyXi2n378w6PQ8HyfR
krwBwMTtwoBzM8OXGjIZtER+X+THgNQNGYRh/0Ga+2CM07js2n89tlZtohpPde1d
yt3nQs+m89WD0fmlHWWfHa9WOptpOSNtV+Fd8bwIzXEsSfssABZxglyMekZ0/pJw
OHECuTwY87TfCoXFI1FbVKxP4vkyoVhHODyDCpDKVbgW7bzSvJbOxDbPwlv0wNMI
NyHO4yeDev23GF4C9LE6130dGQRWWkEApT914ja4TNLkkkIR5n0YFGjKJZMOa1xf
wk/3W1zHCXjPDWTStPLGw7RcD+1thVfrN9JnfBUnhpDohoPVbC1Kxfcs7wvTgIzk
X4Hu28BWazR96rr348d2h/AP0I7QbcZGbzvFDgAZJt3b4KPi7o5MyFjlwlH+/PhS
MN3BREBn+TwWieH/7KZCUW9tuVlxmj/uwwWT3+cBTY/OFppBEK907j8fbSzmvUV4
UhMu4XdxHkOSnin4WCiEiShbynjeLUyWtvcTE07Q+jk=
//pragma protect end_data_block
//pragma protect digest_block
In1w6KtZj5v5egw3mn6GdobrJYM=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
f3pJB2Fyr5nfwcex9OJHrFCgPzDjrl9KJmVcPY93L+WIBP9l0nBbybhKackCcWAC
JWXmrLrgPf8u1J/VbtAAkMgjwKaqCg7ySFNCuHRLN4QtegPzfAjdwJxASw9IfrDu
2jdRHD6Hi/WKNsmTaH4ImWQLndGBm+TRgvKTw0kNC9jn3rNChhDhhg==
//pragma protect end_key_block
//pragma protect digest_block
SKk27FM8iSW541P3oiHkR3Nb5MA=
//pragma protect end_digest_block
//pragma protect data_block
fATmmn4CTHxztFH+c14vb4YD6k+T4T7ih5w3uFjGL/NeoN65Qd+Ih3gLhWFCPQh6
n6sJ6zkz2s+Ksfpl6w4ZFvD94CYsvdBp5xvfhJ3/pzPIfRRL22dVvT1Eh++AwhLy
BX0t1hfENTmqeS5vT4jPRqQiIVQoXIA16n8VKAd0fCzoONNaFWqe7syL+Durqd4V
n8rVuUMrsr4IVBQyLhzU6s/rUomT9Qzb8HD/cdbqmkFVlj6UAWZ5zsLUrfLy+tGa
uxx0oeYJAIiYArIk/nlzCNAZ7a+g2ionUEv1Dyl1+mkjTpHk6TNGYGaErMmctl9X
vvmHkJWLdKzxlwfHNy6duxIn7dHOblKgiMm6zJ5IMVB3aULrW5qj2/8FT3G9A9tB
EE25dXqQ3b+dzqUZNeI580KKqNAKs7rCC9HiQtTvU91hHiY6B8cu6KGGKtZRKDUy
350WKdkk20bU+zG2cmsNsKmfHNQGMbe7AT2PgkYCTIEGXHGep1TvY/KyP+d8Sa0o
NrGzpxHmgx+9WbHZM6GLT3+7VhNBQAVJcHjnDxmKOgwioxV5X/roeVvbRuvMt9Ru
iamdwh3ylRwpcFcHutJuC+UVRlG9hQqvQlsPNGAVrpVd5ezCd1ni6N2V97zk25b9
yfyAiEAvxQnD3hssfbXKV9hEoq78/HzV/Hl/lL1VfSfAUffTJgmMM7KaxR9rHbBf
jjPwlJ1kupWUMkzWyXDnEkd7WAwiax0EPE+oeVVkGgPsTonS6W7DG6pmrjuvqDz8
vXB4+XjSlc8F1ZYVhaZ8Kpsa1SOxehmQrLGW7ErOvsFs4trKQnvUvcXCEB1CUjdW
r87lbRlu22GnIycWMkcrCTUGGMDZF9HN/8b7XrVoEhVt3NLk8f0fF4aE4Z/UyWEV
aeMd7DBMnVbEsD62t5IOtBJybmQH7eo3nR/b8HRE1AZwLgo6DPiR4eAwmHIcc5gn
LFXuCXdR/XG4twIzRmoIhDRr7TOhlS8ZyMvRjNCPmdsMzc2anSzogKNxqHzZph4m
xM7B6kLs8KYoX5O1oRt7oas/srP7hSd1i9TpbwA2vTJVr2C4UkxBNCBNes4UAfAO
rWQCJXU9m2yejDD/V9JEogqQpf/tfA4/0/bb2IPT0dMeoOuEorLstt4v+MrnW6JV
pOdUV1y61cHdqgAJ7d7g7kBu6cibQFjPqCBQ/A1rE9wCXVpeKpHrCV6IUBCQEgy5
cmx1C+fIH7T7JH/ileoWoN8qnOGjqYOLzRmZqXTbLDXUY7etVtmCcB3zR+8OX0GS
zPoZK64Jns5EDR1p0Qx3Xr0uXhmHHBpiopNAVABsSEyi4ySvUbbgdFXhuBUn9f7o
U0EkmeKmnifPcBmni/IkD1YspxjaqdifTyJkGN9BPKMkc9C+OXSio9aZ78gE51E6
Ubuct3ZXb6X3sF7RlYMKh7mJnKuuskte4ijSpwdLFpK3P5Zgw6SdhPFrrhcRNhJN
MekGOI58QalKgI83lf4+Z5oDBkMYCp/UVfdYMbo92pTFT7ToMsX//tFRY6UQneya
ziOGKefowpEJaPo4h6AlQPoMLDucKjthBYsfMnjSu4l6i2Vd2qytBS03iSHnL9ke
znVpfRSVwLtA8m3cReJ9utUgX0qyzOvWfT+9q9BSVKg28zarhlOlDm086Qy1kAGx
K31UpCQYUhVILmHtyyrSjcczFPwBXi/sTs2SDKjBwSxMQasbtRnK86VkhO1hK+RY
pDC7cZ9OZrtBY49/rO8l92av/55WHag3l/nBzKaoxVqaK3GcVAUn48Cwk6qOHkj/
fUWrXtEajIkTwMv6Ou10XH2hC89JlrLTUUkJmFxK5693mKkGtIMZKjBZXedotLnJ
0Q0CHeJKG+YREs2qlq30ig8GxM1RXcqL5X1GvGIh12r0FQiLB0SJJSEVZq2yk5Cz
rP8gCyzrEl53YDzdq0Diq+0KQFBlyvdooqgyQUP5Zp+qU67qD4ZikRlHzxPCOG3A
ZQtSYWxERck9ymSqw9+qovrZfO+jlyaNGbu4sBQlF3975+DdE06HbMidT0IaLzhu
xD4P5t+T72y0wERGJ/4fkIuPW34IpB9Y/RbKj3xiTQb2bAu8q6Xy4nyBg5Smioal
U0OndmMPsTAZME3HUaoc2d8rIGq+U563escZd27p4H9HL2bgDYMcDW8rx196N4Br
FNwoWsYxDGL756VF57Ja3Dw5emkwjOFsd0d6lNkPr2jxJzOS1YYRgtZFxdeisczu
bp4Azy2eO4vsXT36YXDgzzqFzYRu4KAMedBSCnNms56IthNgnUT/E9grCSAZmS2W
gRIOdGovXggjaLkFkH8e8IVTTK6Aqv5RVAFnBedrxiBn7T/RWK08tpYSo/p9MqaH
Fq6Xf04MFElOT1Ttu4DU2GcpO62owiS27exn6rwvaDFwp6rWhlkr7Ln6Xoj5aC7E
QRIjAdHwRt0MPVfgt4uQLQnRC/bg0hNE99CI25B9LLErCLzu7wa8r8NxZCxRPp3+
o2BDsWmdbYrzoiLcCtT+0o5nSEVJuGl3ZDi4YNqRpQkSkoMhNOTynW7DNca01Dbx
kkx/fxub+FyR4NwqXbZYn1qQWX+PAHc5Q5B2mjkPbLY6q00qzFj2lzlFct1CleIC
7gcBze1PnTHZHMPhOO/NvBkYbly03oEMvUTs9PU2VR9OPfxYYUPsXbjQdb5rxV2D
Ob4gwD9D/sQ7lDftnunOIXJErDMJdE6IxPUIXY3PgM4O3PYMXgHAPkRPymZZPVd5
gRkKFWGEUDPHBofZEHn/t6vLCZq/VUtwDfULRzeUMbxSVSm3DJUBVUR0HeoC0nKc
p/4KbDMQudGutnyURUIT08/agw0XcyD75VB5d8ItXM+6UdC7Zg/UP29J5oP7tzLQ
Drh5SESWMjxnm0D6F9pEGW56GALdIzvbSFDreRgaiAAaXmT3TBrbNPibfa/IfG6U
CszRb0FlZ7yZkP6SiyoNtq3xEw8CHRf6TvJQ3tpsyL5Z4aoMLk9LfR/qtnx+nxGw
H0eeS7Vw/ZZyNIGNVZeX0pBPaKAomGLbvYan4osv2xvMcv0y5N/TDqz8COA4zx9Z
wx1+fl4t1lYxeyUa+hJtCbGoSnh1BGdUngvcxKpejJ+f/WX9TYG7pi7iaZqGgqIr
Z3r/sj6+KqyXSvGaXZ7MULiolnA73QVnNAPmAkWZauPBqVAdS1MT4oXpozZnRLJB
UOT9kMVx2IZhkl+D/oIKevSZ6DIuSLMzzoPeUwviMketOJLh2AAG9oebkKDXsQW1
FANZtZSVgynUuJ1Icbu2WNs8vHVGh4O4DtxQU4QQiNLO0yINN4T6d93+hiN0R0tH
cuGX0MLgnT2wroUq0SlrvKttq2flmEEcBIys1qg9A4wgNIOpzrNo4x1NWJS4nsmg
vnVKMzb5SYcXlJ/g4DYaNcg9dfHpEvfvHmmAshu0YlUNv8fgD1j2NfqIn95XwRFd
Prhs6GU4gXV8h5yiyefCo9p2dhyZA6BcB4Rytc8IBr7MbYIl13Banw0iKPJ1hkwO
lqZLX14/yjgVtMNAAaAZTsxnculrPB0vrgBO1sVQF9wuwx7QjAHQsL0cKzeq5uqi
TO6NhecNLj5p54qK1EYsm8uOM5l4yNPK0EhL9q7vh8AXdW5APBBL165SFMkpS/eG
6vUWch2jhb2yUa3MWkkCV61fE2xqMi1rTKFN52WAHVZSKYGZ+/mmSfWdGcJXiVKc
QGf/lAte6Z7RIOw1EP7qXKItdM9D2AD8Usf7UIZdMXqbojmlK/v0ZZMaMsSfM5Aq
XHTy05BSO6GQHoSFdtFNyF/t9rPiLJgRy0wCNLDokd0WG5+tT9zkXiukxfmK7YpS
SoBgjjRl6UFUojgUxNC/IeVRYRJWvj4kUopZi+i1Dn7Ty4KabKDdpSq5mz3WmGWP
fAEeVH5KY3HrgGpC678hy15QgYJ20+aP34y3xaHvZUAMV1A4NbkAlPQL+sm8SYIf
0xHVft2XKJzp5LCw0IbPFbf8z2fPvxgpQ5MIlihaxSP3bNzYIVsey0SiEWts1WSE
PNykQuBi1e2vCciEqHuOajfRbrEsfyOS1TqK9MxznpG1dC1gZuiQi+1/gWinDb0d
y40QHbgrfWKKCISPJMHlF13joDn9URFQX//q8ICG8WwIfjQcICjYYp8Hh6dneXOm
QylE9QmV8v2q3oyD9i/i8AoWX80UuHueeJIlN6btQMf5RW8sF9BdVZq8U0W2OkgW
XiH2sfib/8F7NWU3PR186A4o/gi3vuyueddEfTRD/tyObcKzFnQ7f+cA3usozGJ3
wgRLRv+xAifVN1tYrAD+wMlp063rnzzWT+fOCDZ2iwPq50p/qGU8UONjkVXQ1sdc
VWSfIhXAYF7BibbX/kdAZWLiJXtsnZav/+quqU0/L50ThCdeq47TM4DWZGmdl8Zp
7Hn9yoV3Q/wHN0MTHEINobq6jJykXafXuFumFZoH2TOcOyHcHWrhxvQ/xJpjcPc2
t6YXkJlYAW8oUMgCbu5PJ3VPbJrQ8W3tOefB8BsPAtbPnEU516/fm5IQPxQRhESC
JmhqQutNEnuINvXWRkpzomo98QfKfYBR6nIvtK9fnY8NJU6/6LfyY0cNhHGRkQka
DDfcQRfdWq0V2SuY5nwYTPsq9IatjgO/ca1puF9VTRDQ1sI4OQ/ifUWN2pvWSskH
uSCVNWtZAfG5YV60/jmcTN8eheQ4NhYOGnLRDmYC+A9/WxcaBlvaIAw0NGz4IS1Z
YIdtyA3rGmxH6yztURX7f/NQ+BSpEg19pma7YduyUa1mgtopy3lJYUcL7yVnlt+T
dN7buk0ZvZ4xpGrD8W5PyV1nd7MWrt+TY1hgjZdU9ZlFIuQEIV+fSbqcbIX8I4Op
LP+aYGdxr3e0/jTnoB09ofq+8fl++fRz4Sa5bZiDqfpU6vjDaoSpC7UhGARUOLWm
Lil/PHfJtAMOnL0Ky9LSmN8kEqkf1BEamWYtOZP5zsnFJHAxSchvX05+LJKldkZy
+RmeDClykooURUi6dU2Mj+zGJqoKB8xzSylayAAARxshPiUy22CG921lxWWyovvy
d8sITr2f3ZCZbVH1wPO6l5wPZt7vuvKuTLlVyVtW4itdGxwcf+zCmQvJAFXYqaqy
5Kwcf3lLagQEELWKMfhLxpjN7YZgDLPXRvkhgx4ojRH/XKAeS31V8+/Kb8uSDipa
RBouvL9Sed9lmT4Wfi0mgakH5WxRskA2RHlfFM+ubwWUhqE7yHduWAJMDzh6xYp3
pNZj+WwON0EZYMrNSjPvUA9cyeceTel7+dI4E/6CETVh+91Pat9+Vq+l5mmruupf
GK9N9EHrgyUt4YBqDJRzOVLA/+NMV+YX/wZTqfP6kYebUdqbSXXF2NZVk4OMmrDv
os6Oy9jhloQRm6MOsiDYOoYJWDa3nwEeLEQ5QGu4mrHdU/Te2ocZ0JloSro3YYuo
jTPxBneMlmkw9zwC08b2xv6HKFDURxLj7riWtj5Sov8HlCdc/7z0bTDTCt8961bn
EwLsO0gHKuUiHNRkPAFj97AyBwEE14Etz+TCs/jT0GQcLzi5xie7fri8VT+NgBpu
EU7S+dbrQnkYh6c60IpMCc4IRn0bgNNi5IyIlSxrIYebTtbwf+H4bDO/JjIfZnEf
+khV0mW1DS/57PQDUl13VfI0lkDmpeLG37myqagB2DoNrTyxbEFIY/bUrYzVkwtu
Yzl5WCrqJaWesnYOVDZLaNM5v9ObvLLEp0tUGI9PvR69gskpZIqnx4D8vvNqbgy8
q7PhB/6WjY+nITrQg4RsvmncPpg8L8T7lZV8XzB1KxrP4Y77a6eyuA5tCnW8r3fA
feGXnRlnd1VnPvyjy5PGnK8eEk0UjdcU5eDa0daCRhfy0q5L3ZSgBlipccghCJIm
DSEFV3klq86hxxmKwMmYLASXeu0qiuWXRrE9Kjnuc2gSZ2nhcCVjHoCXPyMDoRzG
sQAQFwrunKGww41wPvtg6QTBVRe57rSWuKjeoTa3CP0fyJ5V4sQydcJwzi8WU0Vx
aotn5B/A9IOZVQGV6nyecTEivQk0aQ0jbEYk0ffrtsVPS926w400TjeaG6SlEw1w
5zAnvEJ0cYYT6NOGKaOfogVAFaXKl8oQ8f+qqia96mdzOCcvPWRukvGzHH5Lht84
gzqtrPatRU17/ukkgadSug8YlwGXkahgIETguuLi245ZGlD52UgEkCu4zaToWh2W
qaoJz6Jz/EJQUxawWbMIrhxHLi8Sji0PebjtDBG5uD6QcqVNS+G9ie426mBOoRXR
KvUEdUYjtnj3PMKRW1ZtneHjJlgBZHZjoqEb6ET5fsYl7YLjBf0rVUUm+FhAsDei
/uRk4EAmPsMPY22FBVd1uNiiv1BFPKXOFnfdTp2ZhHdJxbBi7dQWjJ8nhuR2mSgZ
vuhxKGKifu/hVsoBTEotBKl8Vfikg5LwscaQVcUToX2bTVYe1kjgP6i5kIWB/RKZ
kxP5PoJT2stbzPfoqbsapCqYwGe2j7aaJ2ePJtfc8zmufw1JHDNxFJ3Zbpm/hdzr
5tIizP95Q8Cra8wONF4Vy4DiFkj0+1o9cV59XsdnRsK9AwM5SZpJKQLyVrjG9R0b
0pD/l32SIrHtsOGGB6fjbypasM1f/90fAdYvr515AqAcHiED0eOxmlSKmJTK4sas
5iaS/qXDLw4hWT0eZ+Z6+gyH1+r0oU8XWQqbvYJZqnel6c9KMsu2T3AsIc87d6Ku
cGjTMGEww1Ez4acDL+TSWUk88wXcgESgg8Sn/3YdmWJGFy0T8NmWEo9yU4XkdIJL
8zKWqdsiGtQSdUoNsvbO0AN1jkEEw/tDItII2LRJVR2+Z9VT1PvalSqMybr8Ln94
zQpbo1Gf946+x3ewjKBC4egdUbuphAPH8Zns8pj94JJG3snBGKQl+1ubDezHbifg
L3f/jrNtXwjynxIp2I1B0d457RJ0Pki/wyTK8U8S9SqUch4NIKMu78R48HmNeE64
JsdzeGT05SZ29XBtg2hXPoVkXiNSxZKwTZ9D/k85VBU0IBqw9vJmJIGkxBy8aZnf
kXDc3UWSk9cJfM81agSpy2shCrbg9PwzjONS/kus+xZ6XLI9fopgqbdOuEfA3OnX
LIBn9OKw/TDWn67XysUeq/fr123MgaXwWpXEjxOMToOQCxmqtL1rkYfGGpzEIQmx
zYnAGtT+3cYp7PDyAI3qCKdLuIyUTQbKmUsJb8z0aA2oPtdrT+aUNUVVRu889JtL
oQ/yvQBPm4kVcLWkY4TP0/yT8EHDerD19+O0VQ0p/FjsNPbtsDdu321o325AkmZ8
LbwWrBT0r62oS+QuygrgyheZPf7uj0YTo3Vz5QJ89dZcSF2HLEjPS+wC+pn7/48/
oRhEOYtIBUC3fOtnYU4/sCt75Zyy771PYAywv2ACN/n7xsd2CvZERTsop+xUVJAR
0bOdvP309eCnAmntaHjHyUNs4a5rppFlIQHTeWLQKFDt199RlI8hp9yx8eC+P2xT
QfC3y96yFU5ES8W397OaQLPzu2ckRl6yEm2hh4F8KzxgWmDd0wFp3kmTjllDYdNu
8KboeFoKTaL9+vBkD+U+9tZhRAeOhN/W08I4vNFfWaYyy8NdOXxidcjKuivvwXHS
8VZ77zRaQ3nO3+zTnXDwo6f8JYncPJT9NsdOAp31BLp2Z78hmgHOMP/0ZnR+fuU8
2rxbaaw/8bDqRzCGlL54kfu9chzzE24NJtzRQt3qP7gk+jWMAQm9NBmeIggp+rOq
NSHuYsBHnDejPk3fDYK7afnfi/2FSukcoiVOtdf5EwUwxgJNRVTPP8xliGjd6UEJ
Ai2N5o9EFOEXlp5UK/N4kkfrmGZSuhED0pD+5882y5aYeY1Fcb2RXe14MSzxQuxv
x5PTTwVR2svl6pzBsiJTtC+RYH4cqS/ai7nVGZB4NEmkfuyc517+5/feLDkuz6sU
y0c3wqR7ezC0K6M4ZdvJFKLxJszmBJU+1O4v4Nf2ADKCbUDff9gOWKXWchWdfPE3
Hz3pdeixm/WnEGHytcK1Wm/KEFkEqhGoEOME6J3HooYfxgEA0NEv6gQaLqfE0z0Z
+KnWbB0S9aTO7/kUNpx+jJXJBJ19YXBPSi3ETWIWX7k3pgvMn3lmH8kvn27B2oky
uYEfOpIO3yh5NiucAzHuk5qDC+CG5Kro6F/fn9oAWi3YohN8duIeaN4U6Pafvc49
bjHtsGLB3eQTaEkKbVICsmNfnqFGjWmgrhN1kQM1UfMnLM828hhqjMQwVqRoL7Yc
0zF5vRtZLI/y+QlenisYpPuy+/z+Qmwly92UkxiaJ2K6MrlfTQybosdP15yJL00I
SCOGUjZCNxnEl6qA4EZmfGj/V/G3OuVWrAG77GMNd9gsxIXfB2HC6MJhhkkIZo3f
ErVbD6HAq65V02AvidxQGq/6kg7fZgpgTN9yFlGrWL6IQMflnucwv0P1hb8P+hsh
zL641H07Iwz1744CLuXtEpQhp7B6/aysFAfipeqvw61QaUSiBy3e8+2l28W8KOhk
ZGbIQKaUTmrVczDexsdsjSimAz4M//207aOEYWz9ekUweA9E9i5DHHdU4emjyJNL
rhsuo7Mic/1PPF5BuAmMMQix+TRCPR5DlZKKQk6M8oH4YMPW1/ADK6s1ILp0zpMv
i8opKgeHWZ+1VETX5lqr7IZeb2sUQFVQoEjLCXwig9wZTi2peNCMRzqwwvmbM/Bu
lfno+mtVqxXZ5s9uhdtV+Z9M8oWRBcZHXJY1QLblqeApf1+t3aGakw1R0JSn0Wfi
i0aQGd+IYWqbNL5BHbuyDfPgPY3crO5Vk+4KHIN+OQYx3J8j1Dxd4TGuaZ05gYoJ
VxpiZCq9oXHotMygDMVX43BrjsJ9N4Ak/T++zDSuUbTMw401T5/E3mOVIi2A4/FV
uTFQ3uq2RP6uaBCcNpInlre0+G1YKeXlRgh7iQ77rda9/y4pGluNbl1RhfKkUPHH
l6SZattHdV+1qNuwhcRwhyrBT3TCQ0om/UkL8VekxxFTlfsZT5i64gO9v8cNjOaL
Moyx69xGAPPVZJOzH492bujWi5KhyFk5QlJyWyQa/4yu1gQRiwBZXmYBi7jHAwoa
5e8hNhW46UL14i5o5JJ5gP9mV9qL29cDGyv+qKpUgeSFa61Bc69oGpNOHbvBLfvT
WXVsKCfprpRnZ8gRaPBy9LldyQ6PiJ/CXwEPcbcSfcTqBrSO5HDopvCNW4ci0dWc
8KCtflECTLcurp10/GdsIol673WP6Wz0J0Ktt1Jk0wdsrmDpV52k+AIlyXwPbr5/
KR8px7VNupKg6s0aqIOFAeA3yXrD9Jj440MDxMZVQcUd2Buo9sW8ja2mivfOjzGw
aE1XiKdvWt0tNy77BFlXILHpxu2ocvu37yQDsaUL4MbyPZ8PZukyAJ5OXhi1X06r
t3DOBauNH/MHmgzdI7NNVl6e7POYTeVHGdH+KTWYh0HZG74Q73R4KcDYzeYCR7HO
p61sngLLcgqtPNnUL+g5yzBHpsEbHIQRRcTmGl2UjGIW6iyh7zPrnUkjngwGPzZA
lZrGnTW4iztmvYVqE7F7h2bY9zuWx/RPDkImkaZBCPb4aw4X/OuAbmiy8CiMMJiS
AN7Fp18rZXqStkCeOKShZV3lvHFtjDkeSdD3TtRIn39LRA5Cg2HSxvBHq2mLTgmB
JpNRdO2AL+wjHhkZ7kKDSzocuK29p6CBMbizAWEHkvG3egOFd5rreipNYMJWjnPh
oNnydJE8Jg+9Im7vXPvBMCXqeTiIK4xRcsPegih51yao5k6S34WKLIJ2NoDz9xjH
rCD15NIVLp/pPAQ60YHajNAzWkF+z+m6hcMx7y66HWLMcpjuLNsiEYkEFajIJ+Ad
kG+08tzFJ8UntO74kqOK1ecbEP5qELN1JoHdM7d5EY6dxFIDk6INJP8LfPXR+RVE
Ox7xvhfQTKGwvorsPLru3BobU+nM36UASS6YX/NV4EfLL4o661Ga6cQfpZ6ZoM+G
pBRJ3OHcVNJT5A3WcNp8e62P30zSBOkylfIQLUWqMm1TwU2QpjAqA0j5OlwqUi5e
WtW55kgRDHm/WvHUKe4HmmjF3VMl8ER6HDfcIyxQbDdZdh4Rcl4W9ObVQAVQiAzq
j4cLnOQyjRSrhm7S1tSbBIjkjMGxIJjhcrRytNu93jWO7G8kPGnhsz4xGSN4XNpV
GmXfEPn7oQJK+aICNScbH/E3KzfeTM6VkDRFtnkuyVgdkVfEczq8A0PfZubdLhTe
ZdOerunANflSyfK7NsX3Q+Ch2kaW8Gl2jeM/RTzZoNHjEV9NLfN0RS++bOGTsM4i
Sdd8ggxrmAAKGsX76nZ35t4ymW76w0l5N+qYKOywD/KnXiHyZfAn97UY4FtSfenn
kauw5dx/S3f7RuINadGiEEh9brP86JzcFlzaMx6E7BEnCVKtg5O71jWvK2ZXij6f
HQRsROiz7aFTQR+Y47vJel+ySou9cCqseevFDoAwRqdgWOId6oRXB61N5wrsbpA4
L9BEei8tbiv2TlKWA7SHqmUqUgcXx37/ch75MpwuJpC3pg30zDdW4VJNAfCg3eZe
FwbRo4G8hwaJDDifEWKDHRS8Ww3ayvqhCLrxTgiG6q7Qcjd9Hgw2M4SKPrkuyqfm
Y8XhcDBfwcoNjCbuhggfuKV7yd4SDN/IV0Obx/7NqzW63a/cERRI6Ly8a/NXnRLn
ENTMTc/G2sNdxyYq8NTGKH9XjoEUpkycjhEty0A8yQAPwWxqv3wK8Y4pArvNGqB9
3dsO59HKKmE243whcZf0K2y0plwt9RoHgXv77cRZbYz6b69C9pqKQL4FGJuMMRNN
IgGJ04gpaKYLMtOrvWV2VJjD1C47DK3Z9NggxGLU5/XD2XKTrY4CNZIa627fjGvz
Qf9iRWlH0ZN4+DOu2BWddaq2xFGciNgcyjJU5rRNQACh9wzmEgEczrY/67+T6BSx
Or38Yl0+7qyFr7Iz7G0MFRYM+ymzEvi6iaBwidotm6a8lxUvLuFHK0Bwb0RJjdM0
dRRduL0ahCXYHD7NHh/GYRk6kPkvBrplgcjhXaD84omNcLQMl49kSfDqbmwbmN/M
FAJwxqOV0w9YblGgAILFiIA6M9MQhVIsAhf6q4DUpZD3DPBymg1y0W6Dl4WvsTdo
o98KDMgJO0ve+6aszqxlc+036Db+ZMLMIC+ZyJCviMIk1Hhw58uPgOabuxv2U5ji
yaz2HF4VNIUAjx4MaBnu/pHQW0KXK2IeZCs8pJRG94GOCyoqpcmcl/bqhW1O02Yk
eisgdAIzriLwqmcbLaHv5GQ6WhM44ZMECvF50h50yxdgzbCfvcUJP1PSy5EHbYdv
lIDxapr9x1rW27gx2/z6HQsAeYQeJGJc0kao6+dQCdzYyjQW9mmySa+eifcNkyGE
N6KiYehN6bV2wJ4MXnkO1wLkJSxkNwbAu1+tvsg6Iy1bfBJYNSvOCueu+jIQAC/4
yeMi//LWdk5r+f0WTg//KpeU6XyP6SQyfn2iMLrwX/C0MRwfUzP52ksLI9wJohxT
wIBB53thgkUIFoX9de+pPQcPbe2IZavKF8/ZiLF3fJITobHHd8n3gUI2u6GGCBia
CMs0LfkEl7mGmTgWIZjYENLdYRFKD7MIlTBzkA52lvlx8/I4Bj1eWTLqSNHxK2NF
EBnWXxfT8ruqHuFj8vhMo3LH6lca2gPS8PkObP2n+ppnBIzGgyTpGq5Sf0eM8UzV
v+PDpPAjwwf/aYR+E5XxqotXzuQdlIOVM6HTwJfFGIC6jvtMBjDqyt7zhizI/eJr
qQ6k9k3kT/PQIjQqKj8TYfUpjDLKY3X5fVbyQ1hzKCSaZdOWbka/yZxBmkDxlPBR
AgSJUTEi5Zxk6vXZtVWe1X+MiIwvK+wgF0zSGanv9R5Rq8ngbvNBS+4CV7Uyo+4I
NoXaEBELGgJ3iW9WJkJXOjit4WMLWvoOJpksZcjWcFpq4ZDrhtbpSyPTeL5K4633
CpClyZaM1W5tlXnPrtgcT3UrHYzki2XQq7lNBvDGpZZk9LsNKRH+jLHEg5RiScMa
SSo+qCqHfShVlsbzk6pf3kN0mlxfs4p8/3Pm5qDdrqiBpgVnYCRqjyie8zryQhsz
eWuoShG89CCwSdLdHvjbTcleLmdv5gbzBDXDQvEIxJvnj4e71yDcGrjH+5aaLEkZ
k3aEAJL7PuYD0t0LP/UkCWLbb4alGGAU41oadIBsyPJWa7sDP3O1RLyzhfqaVCYq
OhQf/Lcvfo6+I4LLvFrJY0vPoTc53DoDMmr3QpCDi/NbPUlbc2mvZ1hzQrukdvpG
Ibg6W30IypEkEh1k2Qw0FzS+g5p4VWcsf0Tr/RCp5aY7Q/fnSG0dWuEj65UipWtG
bZp8sVPvPjwUcx2PM675ay5pOLg7J9OdFiZlx1/L4kAsC1Cq+q1a1uGT9Loiklhv
e4QL3o3Wby0djCrQ44XhVDq54Tg8ddV6n1On8Cz5W+CojoOmEb/8Cum4uN4Yx8co
6yuuMqrVq3oOeszYUlA9gmFbEwGwLrlIrZ//GLEixo8VBUJjd9ZRUkNgqf1Os7d1
qqf3/CdgB2qHs3sepL4n2tkXsYYhNpM69mPEJaWJiEphr74qd1PiT+A4ehfmydb0
PRG59s/OXjkHKySZu/m991+WX2hTLMN8vni4JXJsl02EWcHxd3fBHkm0BH2q8hb+
Br/0Opk7yAhBBhg75iTLtggyFSIKoiCpPPbOwXHBVuRGmmSILf5DZ1SPY+EiqaSr
x0qPkJX0QnWr8w8doi3dZUueuFDUrgm4LvZ04P+5riTVo5ZPBFfi0tQ8VlKIFfM6
cHzTDNt3HmxOqWZfNoggoixddJvMs6PoFY4D0ArkMCRilTb7kYm0QXIzsRI32Eh/
HBSYGD/xq84I2Mg/0XQTUg95I9sw3udSWYfr0/fx3udglR8aT8OWzjgZyaU6TY52
xNNSVnwSFnqX0QJxtNbUA6CIRnYLm4Ja+jUNBV0q5p9qQGg2mw2bmgmZdIGufZsM
P6wMVeaCDEXXOM9nM7p2DVdLSB9skhPcCThApzTnndI9kLKvlaTdtgWRhr7eX97a
CbcdAPc8aHRo8bCglVNlWZxFEytd4WEED5h7cWl8myiOtyf5At4bXdowK2QJ8dde
VSDgRDkQXTRit42qf7/RDWB6uwYOtcBL+fln9qe9Gf1rY7TOrcv7aLl6jeLjQH5K
n2hhoDEDuPTn9vvxHdOfVPBToM/KUVryT30p99Wih/vHVjBE6WC1SAxFRtDPhGUt
ia3R7rJzLqRLPM96ilT1X8hiPYhgXfuU5GRbO4c3L/6zaEcoKRJUIvBAjuH9KLZB
gR4XzTouefy+jfRpYEILPUvwwUfNziAUwdA89hUZVNcO+3Pw87qsSxPjK34rmEqY
ImDvncw0wMPa4GVKJ2qjPinAUoQcGM36G4Svvtrlc0THkSh7X3Hx3mU420Ow5PTd
gcuajrNj0L3mCj67O16/Ql4ihTbRlpoxWwFioy5Lqr/2qYMyd6kP2Li8xdJ8eofP
4ApFKv5fPOIATSTdRkego5Tc6dBW/fatJvyQo91BvnjrCuO+BJjsGANpSKI0KiJE
CyQ+UAvHP/YPHlBcQUOVeEA+RylmDO/YrVfRHDMViZf24RRQYkYMQTjZov1273k9
lTYPAA+nxOAB+7GlPnv0xHJxUKLlS6x8eeOJyE8tj7LYfhx8ADNoz0BQbQPCRjII
kw5Wn97DQUznrtvWLkuXFcUhTsLZnE9kI9gCZWCAc3rIN26JZhoAa1pla/4dMlpk
Y434nnFuI+Hw2XCE4M64BWr4CZcfQK/sM+kR1Tng/jarDOOY1EJm2Zri2OQz2+aR
64LkgX5s3tbN7/wcEprKX8w1IxMcGGESM5qizip0MeLuFt/kGl3RI7kgFPHOpWP5
1XV1fLNLeHdn05LHppBjAJOWygOXgmrWzcc40/3ICP2JzBWEqlLfU1T4d7huyErc
jKpKWz9IVoP/QzBACI+cgB/TGJ6AwVbXkF33LUL2hDBTYvB6tS6EeNdID5w/P02O
gAGZaE3A93fcDHaS+sn1vqtTB4A1xSe6I8b36qcFZFRMaKCfFLB9fGfiraGt8gPe
SQx6pYmH+HWwFqPhavpEhaKW82OeE28f0if+5LzpwnM/AR9/HUG4SoUpz9utonkr
N8ct8GcRmoE6KtZxe20fXaPnDpJ8xexiCWkVMz657g16KWpeGDz/pW/18HiKusPo
2c1jrISrOL5rYNfpsWBTN2WOsTm/UHo69NasqMQIVatHFcL7k/d8HtHdwm9igbLZ
lwqFbVFqrKWT3gjHHEGByBTrRpIK/fFE3et1HMFQBglG9oTEDjOdU/Xlzm1ek3dN
42jbuTsgkAcN8LilDqDFm35z54dy2fr1wWpvSrAcGps9hBujji1vsU02s9NXSseR
6Pw13xX7XGwx7TG1guWImXgYWjCZJkLcgvZlysDZtoavhqsMs2OEkyh9dauq+qfo
jzXL10CAdBoXSaWMWYlPfxkC2c+fQ/AUxjvUlxKb/Vi6L/yaDiKkGlxYySMQAp2y
Rw1jxwbMrxah8y/jbG4c3DZAH7PuIbenwXyxyU4MzQ3rCnZJPkDjPudRtKfWjAwT
IuTM4H2QQ7yCMwJPBhbipUMqVDC0oqZMMBmiStFZJR6cEeuThi9n80oQZsl9zBW1
e5iFNjsy/cUwm5YfMedYfQSKPbQGdEqDKMpTjezOlPyVjLwBHZFuTQ8FQE1SrR3+
BQKs01P/ohgh7RVVdGNl0yfV4jwfpzR8CJfkMnIibmB/R53uPa+M8EB7nE+TBMuA
7DFcd1d47eO5qgjkMPl/3+jSMJR80+g+gQGGs/NU9njctozp+ZLtWsBW3e+9BUjq
NBN4MnDnXP4zQ+wYkJIzXEjnItvNsZ6ZT227F3Q3fFAueCzK/tpAzXVvfrTQSBH0
BfHq7l3amrjo/fMRUaByrfzTAPhpl98AyeZQt90sJXoy7gZlL/AHbjwFvg4q+Tt4
uc1zytayBmIPTeQ4UxjIjn7NA+hrqG5vNpJ9srOLqXPD0vj+9W9o60BqcI+KjfOh
mA3NE801XNc/BORxHnEukB56qucN4ZYMsHsxnZy9yIa3sIFeGBSXhMsV8oyw3urL
sBMNxJ/v9Dta5pr0QqX1Tv3LCSSsZqRGbia6AjvUBUIW2WPC0XArCX7L4LCFXBF4
NR5hG7ZGrAytuKPY7w28QKmSbn8aKOF3zGyAExrmKG2IFbwULJqZEPjizrzcS8AU
BV/mezcoehKbwK4sfhUbMnefkLgt3v8rdjTlr4iAVe6cxqGXj7Vw6LhSW1ww5cb8
CO4Rs2x+U/t3XbU+IXF8kxHJoDceI9pUVbMJMQ+1SXNorVZPxpyLwWANxipI/0dP
YzgINSZP5BqQswARbyiHS4U2ykPM+IIOuKj6quVcvpfYAjhRRG62gfyXhKrK8WSW
WDbOlwUL/nfSenjvGxYNLDkxCvBVTbXEm/LNJJzwPXNEY1ojofw7JMuE25YHB/J6
ZOB0qaXMzFPoZrcqfaFPw7TSwebnLmm49eyPlJyAtLpIxxe/qXmxzgHKMv6JsYNS
5S4kaI1IHjS7xnPgg16+zg033UHWRSRvteYBXd7XWiqYB9oyBpkwz4mIke2PZQFt
tS20xAWDKrPb+tgtw7w+SOFfutBM7umnk6olSV+THai0rG+x2618cRzY4r3vPevi
lT9qdE1WlOaq8CakNLO7TfVUWUExSkQJUYJtMBRxg2o=
//pragma protect end_data_block
//pragma protect digest_block
1XEvfwko53hCedaRmHgIPG15dPs=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
BWNOq/qINymZnHet9kVAm0NV2l9/Ta5zWYpqFm0vxbpWl2qzSWAx8saJqAB6WRS8
TTF55nWtt3LCM0sqUjNqbJ3SkSbfijzaqPeHKDtkJma6L/J/YYh8+t0cpgvzcQzO
yWVQ1LPlix2lTgvPUlwKhvMThleOWLmvIwfRSRFtj0fGpB5Hox6jzg==
//pragma protect end_key_block
//pragma protect digest_block
QozlpQuiLuTd4lyMhnXSk7loZt4=
//pragma protect end_digest_block
//pragma protect data_block
lyft89/Afsn8+RieB/6CFO3JR/qqkvn4lPLw6SR8IvVcpdsWA08kihC9Su7DoCKw
NuBb3R1wEaLZZNbc1l4imfwhh1LJJWqU7Cu/HQ0p7F6p+r7FnvlmZjc1cvQpm8Cr
BOmEpWPYQ4wQQtneu4NNFibUeWVsKtqAyCGoamuxC8GpUl4svpRrqS5s8JBf2jgN
LDDXaNMnl79WNyGqEqXwqKcfA5lgT1wN7ci9DyueEEQGRTGoAVTuxwlsRijxolWj
rSi/wROiTu/azLx5Wr2pLtAVMOXfXRo7lWMzwoet0PlXCNOTuhMq7uqFPK23I8YT
+ObSqaa54t0SNwSM8BGsExjL3R15BBLSC0YiIKyI9poAPqXm+3DxGBnR4X6+z2Cc
KmxtmXnUe3UMHA73KKjAhMMT7APL1Ae+gqrGD4vW/XkbpC3R61lTb2f5jQfWM3/X
FE6PzCVfN2wb1XDvCoMKMjBEUTUa+GtALiW7yvc5NRxLYUpRHwLbV5WBjrUXMaHM
l69n/GGhN6xtZ6g8/4tODUaNKg5cOJNlgBK85d2zBWLSdvDgEbg80egvGhxDzVGi
5KT0yg15BEv8GG1zWb1ZJ9zzORl5iqj7omkKP9SH+xhdYl/kqe7F1lesrSA4O9wO
O7IKeDP02h0R7czjw7r9pzEpQMHezx+rqu7PoaMj3QFOBCKdWxOLzXOaNoUAsR3w

//pragma protect end_data_block
//pragma protect digest_block
5FKYA95zvJvJwOPKvulIxjWD3uk=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3PYqG7hYjrB3UXDtJ/AKlbUC9TQGCBSfUltTgBkOBgzebWY/+3TnmkB3CproxPGo
5QgYYvG3SPkCRrtxZ3riZ5LFJyIJMojaIB29tp76+vb8xhB5g/J9s9FmE1XZprSq
MwGDnA3VGbzDFCXJhWRR3OD/f5v1z2wrljCmEP49UGLffXikFbJSMg==
//pragma protect end_key_block
//pragma protect digest_block
B4FTm2KomqLDcz9pha61PL3XLKA=
//pragma protect end_digest_block
//pragma protect data_block
KPRNy7f5777UuyPnYyxsELa5VXE6PbqsyJxs6RKmwqF+JBqeOucbXeN54MCLV1eC
NnYivgwFV8bK+sM9Wc1lGsJGpbQOT++zUMsaa5IrGMacqEpdWbz+0Bn176retezm
7Q84WY0JJafYO2AFYtz29SNLeUyQIp6FS3Qs8Lr6/Bu/Xft61o28qZ1UkT4IfwI4
uvRWNJNTIcSFfTPih2R/f0Rzw9b2cHvsZDn4ZQi8lKqTsI6NUTVbxEkRXnGRDmWp
nXvoR/DbAWbuo2ylV9pFZCXOpLQz4nRn+yvXVx4wv+Z/kdeppUidX00x9G4gqZGf
tt4MnO21dQ0sTv4SQOc2x6YD6HRsjhKyy62aGRWmE3cPqvxyjJl2BQ2GaFsg1qVb
Y3+eJ90uxDDrKl3u9zT10vS2ZQiFnsCbtm3wkzi8oYTEdKhbR2RIZhCEdjGhFYHY
SDwxjMAP7esT9JQYAPhw5ero+TyxfwSSfRjvBCa7GVRJNa+UATu59jSrX6EYou5d
+Kxfz+q5YbG+ToDWRBRQHyaprXulOId9rpa8ra8fwRbAvrOG3tLs12hmH1DUBGni
UVr61Ns+IWFUqD8/m2ZRxInQyxOmRFNwZnouxn3Uc4yl55sbYsMCwuoZBk8ylS2l
ahE73N3AYcbT5R5+7e7EyQySfqAWbXOIoqb9M1yF2fCm4Vpb+/zmyNnW8YDAyLHP
3p1kgCgHixQ2173htvVY3LN8tPYGIxpzypa/Z+1G7CCQ/joeQq1q6C9bq0dS2Si1
XSHrkb8v8xK6R4jxA8YAoDladtFJBBNkf4HYl+tgOcbTyytmA9R8VruvFPqalk18
yHkakYTWL43kBFap8HlVHxcHvl15bIPrluCQtOdCVFEuUVbnRtymimabFTKV0/21
iaprtUtEH0NI1uIvK0i26AEtEWM5NX3G9dkPZMBF+MGhOwMofGCBGLdABZMc97H6
MHGqi1UTyOXOdAk62JXH9q4mC99/ErwCtzdmZ82Th3+KLiMIjryFocakdtXL3sS/
69O5PJhnjbUpAgtmcqBKGW8EjlZRjiUSB2cUWmd9JDxy4VjpxtaW/dMQeqdyKZ+d
NvZ7l7mKFWolHpFooGXDYty31O9EQ7qGvqCYx0GLlS7yksjdw76GMmMoepi9B8rF
kqcjbO6GTaMcvXgT+IDHjkBo4OUglSmKWWYQq6rFOTM08632O1cglc5RVBboX4wu
KgaAUN6T5/3O4/fjof4icZimZCqHP6x3AcM6eGStLCnRahSKIE4N7/HPWORVteiJ
T5r2J+GqHJhwSI+I3xKZ7Y4TsDAy7p1cGBUSZqCIlgYJjzv3jrxmvWVGaClWColS
CW1XLH/tL948D34fhW1xSg9F2jlAyyx18v9pfVwcX4XfjxQC71wDJwcisH6wtvQU
YzKdJCDTxqP4sOLEsZrnvwYFX8lSmb6kdiI3XGfBfAV2xjcK6LtUubjNFreWqBYL
JPht09k0qd/ImDpwrmBDiHcg6tDXysyELhMaWKzJyPsoXL/F1nFsNVo71Ur9L3PS
E/PekrPTJbLat3QM02/yIZmbdWxC8eThf9i43C2b3GZUjwcwJHuqBzW16l9ZOlWt
lA1C+yHGAUwcUl07q+IMnryXI07kxmveXGnXto4JXl13bDQQt3F9oJScF4gnL0W1
bsKR6aoE1mSR6k08eX7+MC0ACGiBxOkTjkNZq/AZocaxQLwb6v088bmfJTcN/gIW
W/1LCdEre8tIVhPLFnmmhsrwsroO7PyaC/A8k+Ev3iWUCx/WQ47X+ZR/mMdYBHNA
QuX9vgIsn+cJ2yc3NmhR7RLaxuveB703jzEYIQfnO9+mVfAmxKdwqkeyQYHHsCsh
8xFOQ3AQHiDSmE+qwwIA+zNtpmLS1uFUUGFgTn9Jdbd7IHCqGluxJlAl42z0WrXQ
mL51C2kSuSUCf5AnXUT2vZZHBSVBenRj/WyV4I24JyV6cjC/N9k3Ty0LuprSq714
oyEZAdDvBLJuByRELScib77qSHX58KXo0+L+aKsR1UlNEsmVcRL8g5+YbnYuUjo6
Xkmdvht4HVtegf13kgMfZmxHq1YcF+UUGbVc7q1LSB1GGwq/Yrk4FW5mGaCZU+Uc
jlh85u2Np/Ird2lv3vMO3ghQ6GaMka1xgIHoxaunXTnwLld7sFggYpy6lxx+aRVm
IdegHK5+MzjQFaOElI/ok3nWwBiEoHTGXN87GsaEWZym3LG2DYTjsfS7zslE7/RP
aFLIfUBi6r3V9OnyPJmZONeTU9OQjgA3RIl+5MESI7DKqiTF9bv8v+o6VhTJmkh9
T61TXopm+FEvKBgYWSiBYUS4ReP5kQOmTas6vBaSnZeq7ddse5eXg8KqEEkN1w/v
FI3emEgoe12p9Uw7fpgudEkCF5V/1wpe6YBUsNr7nfEQsIB4xPr16PVTxKHWT0e5
+sDVZUzGjLyCaoY70RyKnqhut2d5HuE09JxG6xc6eZtV+dXUTxYjKkbl8C4yvy4t
1z5kITOpqMl88y+hfXmz7OArhpiw5FSbdeq2Ttfi1XwyNh0nx8E1Ilw+NUmWfmu/
YDNo+EGv6O3T5JQmkMG52D0LaI5kD5Ba2dLAi6srb3f7NJYdkdlpAhLzmsRDEb+i
BsjRl0AOKwLOQLKkpXs5ZbLwaeslrx3XwVYXZdTpr/eBHqD5Oc/Hp1rq7KwOpQS8
X/bZKna+P3TPKQkgXEXi7L5n//zWgrI4Ym9ivi1+KLAVt16AxF6Krg6Pj8JngDRD
xt7r700jwIv35JLWxpBU3oj7C9pHlODy6jn1CiwWB/d1C7o8yw7WzWmeLR8dwDof
7IBobhU3nsA8V3mTh+lZUjDVAX4HI9ojQb1kR/XtklFVbhH7e6umN6sZ/Lrcp3Ll
qwtP94Noo/lTlg4qup4+qLqAvp1LSiIB4LWD0ETsmuv2a2Yz0EqTJKGl4ZtJHWML
11DhBlDmriWoca0H1LYK8j8fI4QJadzE3/e4PX3DGs+xRpOWtMzP2tx64/VTRTMN
WlbtAaiYXyE2/6n33aFQvBVBNKoyxEYP62TDjXKZDZlpU/hrD4RZrrl73QTKQN8p
K/P/Uy5XrcYNVIM91xzqGYOARH6g7Yw6c+bG/Kuf6hy1vFw2PdX6G2sBPbKkmv7X
254pBhOUrYxJNdF//CN1bl6ShV+uxffNXLHkgptuMMNVgO0mW4BKvCrqwMKZnJMt
NAZdU+PtoA07BsKWpDdMNGhD7wFjmK0QqmvmBWoCBS0S6dH9iBNwLk25S9qsVas6
STnXL7fCnhVkqsYR2xbHlzU71tpSt2nI6wgaMhyjSatjpwyWwUEfFCPDjEg9DTNs
e5+89sp2ToDvl2UR9g57PSqpGj4DipAL7slHP8/SaMfZMpxTJI7vs8tbhEuf6tAi
h0Z8AIq9skBfMl6XQ2nShTGkMiQvjXuuNUTTM9TdcHMvM4uJ9OEk+DODBfUoV6vY
WPbQwPYLNlRGVGqqNPSDpAyi0kouc9SDslen5qv/ikSdbtZu1rSW5WUBbRWuVJef
+F9YXKoX0fgJYdtor9b7aPhAdelqw68zVqSQlv0YY3gmBO3CZ/elbfkqvLVYNPgF
YP2lsVxsdWwBmONaLlEn8bY+zHLhyGTUOGqqyCZVQHq0vLYNfLvfkvT2hmhrBNQ8
9lGKndjj6TW6iKXjdOmcBUvbpwnEM8zztXz8rYRt2tKlTN0Mb2CSQ3nCqATUlcHP
zmQlJU01yhODYWxiAVRoMKpVbv0Wj+BObXUqa4YwvYt9jU84qj+ORpBMoEpW10Nf
xixYNUAnjnOd7lkUGVoPgAw+z7HBhov5ar7/U5+fupYjl0YMe5jChKzYwJla/0Ow
ewlzEMcs+KmatMh/U8BEFaOr/sczWrbMksoZleGsbmv3F/Lc2dCnqP/pwfcDwBM+
x6DYU/ocTawgXEVIrU9LgMlmx82bpLSK0mknwGkFeh9cp/VtiDJeyNV6n2qMpJre
XhxD3/R3CN3D23X/nXY5p3uFpNUVYDh/pvSQEq4sJjX+dGyKsoBEu4FlfQX2V7KT
ik47LCHZQzr01p4dTHdrrZFN9PZjYENL0vPvKuexN8OWp4eA9ukQkaidkzTNSknh
kvAB1ymUtOs9cLu2jmckKfp3m91p6B/mx/qT2z4GWrlKjKFQWsMgfLLrfOeY7xI8
WMHZ0EA8lI8cy47P4JvO2gidLKsaESrpca4pRDhte6+V66uKQN5L7Fc45EBzJFcb
xYxdGfhIFTxaUM7/EOf/UYwWZOwOv5QkN2o2pZr+Etp5eAaGnWj/eWvEDNIMFewt
lWAzKhXkg1SooCxj77uGL998Jpoy0KXms81cM+/I9DKUHpkysz0+oAq4cIJgx+LY
0ymPAj3PGDOYFS9FVAolfAxqBmztd+mpVbuIK8nmg84egj2XrdUvCy0Bl6NAaHDQ
0/H1Gaa7XVIAJidzo1R4tCECgopKjrtHVQmKyXOMguMXwGRAyKghFvpv4mLXZlq4
FinZ+UjVGNAjd50Grg6mv1PY2ZtAXuK3uHYrsiVEEk5Jsk9/zTwGaRixVN01fpgn
Yy8qTPb88/xVQSKDqWDoJr/7Jk6/z+ZmFkcRS/3mLOdo1SgG3jD2Jk56Uq1ULH3g
Mlg9UI3O958dyPr0wzFbQ1rTm4aYEwxcBDX40WEJsOuClKKS+vVIiXWsXKJxDqx9
vFgmYUwYeKbogDziVeYXKdDaoWRp5DiQ5gFe2A7+si+rmL0dXVpj1yxUetrbk3MO
NXWR0jS2k53mN9kR0tlh70Q5ZLbgcOtyNR+CBPC+rQ3/dj8KuzvXk7ocY9+wmVT9
m9k2pNw35LaOndXY+EK2SSGlv5UIZ2XlbxbaSP94CxRZzoXA/cVhVukjZYg6mO8/
kTdUDAHWXoJ4TK8zzpnH4pBMDNc30Hikb3OEml30UOnkeoSiXziCI+h0TNsdN30X
RnMGpCYj0LIg2naMaf6R0VGNgTBO7cx//DN1djsvUfPTt/4WbfJVCCCxyWtYJtkL
UEdwD/nS2nrWTdokmBbwn93aNqQIHbeCWkyJa5TFMpMpcA5qkD5xwUAM2vU01j12
BtaqaJ2n/en85oOrmhFRpP3EnF41I6aVtDTfToPTY9XtPyLubS3frYfkBSGfK77b
NnQV00MFGGW5cKeaCtzNnZVlhbplOcRr16DX78nEp2/WpVJ6xZlziP0TdoiFrrWC
9tuf9dBcwdaXOCgTWd0WV/njxK+wo0zSgAOTqhI/24hwAeT7iSWkhLZnyDbkxVXe
S0mVUtHkqreDFLPrvpLAIH1Pe5ZF0Tx1B00fwJsNv5zDF5e1di+aReaxLQNFBfgH
qDRdEXxf6rWMi59M0sywrwnBtMS8QdtH+OQO7fVwgQnhmKW3V8g0ooPgd3k/sSz+
B8Qn7w+ZIO2E0zwp3xe3odM+gTOr37xVQe9kTx8Mm9wSp0otYfgyuD95jegwplau
47gyUv6s5QizeilPNMGZxgi5JV1IaqE/lDzZFLfoB8OjtA4m8oy29bLqUpwmnsfm
HIgI6SqcPOCyRVcBpbdduUR4ZWqfSdprwAdOBdhi30xU48hn6WerWzjnY8SAz+wZ
zrDJranDIgjNpIrXzQG0Ft/ZySRsNLSyzIHbMb9zzfEB9it6ByMT+ZoyIAe5EC9h
ylU+adimoa8FP9YoPMKRoxxqTxgTQgQPJI+fD0fgPI1n6ton6Vea1YtZHkPvbKVl
xz3dqKsgNXkZAMNoMz//ATi/mfhMD96QThpwe1Mf9f9YcT307zuN0l76k73bgxi2
IQUKQ8Xpk1F6qNpUpvuMJQtB2F8FC7LAr0xpsLDcKwJsgn/iu/y4L0uqiQbHgq2S
Km8/aJCgKFct4mjyUZUqJqN09uwnhIdwexnVCcPqJqLp/V3zm+BpjJ01F8Wcg6o/
p9TgZ1djKSUmMknz3E9WfJePImEBuDtBALMAT+o9NsN3aohfkZGdnRGAgszi2xeh
/SrISkt60olzwOCoV+ptaKIB601ICVIfVV7LMT6wYdBKg82Ybrz9mY253mQkzNkB
DqGcCG+ICYP22xLJqKQI5uP0xyy1GXFzGrCInYJIa2J69McUIMa0dD/9FoVLRqrt
xMdvarPC14IIHFVMxQrGPiVIDMLxn0TB92EkeVL4Oa0WNwBAI20P0zN6vc/a6AKe
tgnFJPCazukWjlQ5sGhUD6d/1tszy42e0Ngr7iw5pssiy1MOwh2v362qe78FneUp
6RL5vQ+Acxv9R20IqI3kBXZlazPCQexflho1PNpBEFL6TQUDiHOuXg5gl8qu6sQB
KDIo0XL7CzmYboZCqUa9TELhbXs+zZpGXw7x1T+5GOnxNFzD3d8yeG5c/yLTeRur
HSx2nn2sEEB1mnsELFEz3MH0A7/hLzzZ6bsFAzIgU7RFjokg2NS81mkbZdTJufrO
Mw2dQuDLbKY4Br7QNxydUNyVcezygFo3ADaFELk1/Q7Bw/wfmY7DKjxm6mcuUIFe
7lqutUEyt+KMVw+EBBpiDAwETkvhN6dOa8UTbkZ67E7Bilk5CqXwmHYemO4CUsQ/
6CO3zL9dTC0rOVOVoIcwXw38Pn1fT1iEr1o2bTJB2IUlZPYsgX0tpi+mMwy/z1Ju
aj1JM2RIWbKgkKpKHxHHnoPavCmwYyBQwpglZWdB6I/dQukWC0rcsUxS4Kkm1zvx
F8tacxNnC49catzbO7jeESylo043OfJDR5TakwWwiS5p0jkmvqBgPVBzSqJbviQm
vluRBcZXKEDwAXhauLd4LaQ07Ok99CavHEvKnMvAxt3CIPmPq9HJiDml7omZsxP2
SjwBqKiRr4pX/DLVFHvEadqRDz+2VebQYF4R1F/elA81tIIinbEBDE9kVYc6nqyc
mDtFH2xVm1e4zQa3O2RnbMBNs9YkdhAkk2TfRyTocAk/pYkcQ6yxn+hFZ9UqSiN5
ODHA4ISDms+ykWg94KtWFeWgnj1k/KbSQIYQ6rSoaJOvu95UCu1rAAQ2c+ofpoZc
qyoK9to3t8Sg6ZeHOzhkFC1QFKu9wHqLOFrB3g41CnJ9wWqBuRbmXSxP2GWpp6zc
Fq2hH0Z8n2ZDnE5IZ3BElkoiR0/K3VkMfd/9+X1mf6KZivY2XGD9GSnD7/Yv2aao
RIAcrE67x6bg5ESlYUCqnVrXeE6A29zTN4gUgRy51xywFwLRfdObl9CSGvx7dPQc
tqtnyCPigfO5tvSrYmYIn7IZnWyEU9TJpyQzF0/9x5/FukM5QcVgM10tHT5hsJJa
x9Npkgz6o9F87OCBrfuXvP0Pjg5bADMklhFtn5zoio7NMX+Xsc6k3A5j3cXIEsa1
TBfkCoD1V9/H83LZrxqEOfZMngmZvddHKlKiB4a8+RnzX5TP304dNSCLXnT1R3yZ
wglQS4eJO42LTGq7WjS4DKUi4+7PAJwQGnXN7YO8LHRVqMPiAQ393EHCpUyoQEFW
fi3+sz5Y+dvBHj3QdbuqQLX2/gQa/mETFwnJGyGK7D8OVSRp6bO2dbpUbCxkkRGH
/yY15S2LSUuvgC9peRjTn6pWrEMXmOTsgbR1OQze6klxMvki4DIiMJQcwFZXpBHf
6ZvENmYeYeaIR4NlNLJ+3WErEp1NJrMRaLxJdVStPMPWHkv9smQB3BKNiEXQ/gsy
a+5Gw+fXgebXfYDif2/HGiXWY5Yr6VHNUlNywe9XK1lyO/Ra83sBSIbwncQRXHeo
HYncR5P9C0eQMq3nH+0H3ZsP1Q1W8FHVnvrbQPRMf15k9E/4P4zHe29GE4a0nMHc
c4imFiSnxLcbWmGMqn3qsMDlVTeHJ4dQELdKePTpw22mUaDTjSuZNdGodHME7Db+
2h6ylkZn/FxYo0XxFjsLpw6eZmEvQvizPa1m0O2+prdnBK2vTKT/9jMXgSR6L8nr
uoWY2T/acC2QFh6yjmwXGUkPE9PwMsweelsqEq6+Ajw8TwQ56hYH3jL/ygE0uZkB
+G2JH0lwslVKTidLW9ECs56Wjch5OWEn8dRPkqGvM/jfRUk7Yq057hx51PqHhcnZ
b7Z6p+wDcllDkaeB910FqQPAEjVmPck/YcwLoenhO9fKoee99XfiKAssMA0GEsE7
nfomK8UFWf7Om8VvCRjC0/QkHcR86l3EgY4id0XVjQOkHutHAPHiaCoMcRq4zhnR
i3IJ0ZXKEWynQwBerH2vlZ910y3NnpygP59NbXxvOU75gxsVVc1+Z2Wm2c3Un1BU
aFCJMWIOQ0U8NA/aS/GLO9+xaqEMyiXt8QMOkDCnCc8fbB9wJEUYU3HXI+QqfZsF
L1o3t+ZaPryX/7yoOGozqQFhrYiSF1TX5ghQVrfFpk+p9IETca6Nn15j6uUZV402
XCCgThYBopUJy3EjutHyiSVwmhUgdWtGlJchSUiqk0Wyt3FXep6XDfypPtl/IaUN
TJC39q15KiRdEp+2m3VkEkDT3yK1xP0G0zYdfjZ3/HKXy1CCaGontZwuj6AinS6z
nHBfgx2SnnaovtY1exjQHFYaeGX85jFFOjr6L7Tv5jUSgfpNKucoD1067yajklh3
74aWa1HghiVcgh1geb153jN9t+wKEjGj7Bs95NCdx3Y144fq+HCAXmHu17ZLtCz/
vUGI4NCozdF/KIiyJ4SBXs/QLHHRXkhpF+in75DBDgNAzUOP9OK0H3fB0yOZxTtr
JSyFjTPc0ZIxA1EK7geynck1G0qidIV8AUW3ox5P66xhTJV4sLYxjhn3aDFsDKZ6
dGDQ7iDI0oo98r2WaO5fatxV+5XFb+kMmHp71eU3cNQDQ39DuwAJ690vbVDDQzKq
wquN/G1e762gGVzCQCVSpWIwH+NnCH0Tocznnhjpx9RPtH43CRM6iwsQ6vtYaPmi
vYpTY0wqB26ywQJWEo/60P7LA5izZpAC4MyBjh8hrLbxxvzmBBs1mFJ0Th8dbHpf
CsfmpsUS8Q1dvlTUr7fufOEi5Cxe+VjwrdqYaL4s09TuBP3uVI2mre2KVOAY38fF
JeAQd2uxPewhhY0MXujk7GfrmNgQeJvmXnqo7q2e+PoBfa+5LJAhrwlSwsDMxSSI
i48HbJxbFw1ocFngM7avCHPe7kgEfdZbCOCQeOIg68sdOpcj9EbETV8fvvAlv+e3
gWK4yewEFz5WHuFtWJB0+B+HOgMKXjEIyP7NkFZhkB5u/nKwJ/IQrwdNFV9VF0Kx
G/GRJlWsNuXOfURvzWmYGgtrF77eAe68NjEsAayribcX6p92gMZyteccPeOtJbYk
U0K3uVHhwIvIomulB9HhAeaUIipX+YjtBbMmq2s9JsYe1pIsojfLRWhxYXHTBDUU
lbm3itkAZXfcR8uWF/+zymEdNw2r1fpipZy2uKlthl8LxdbhlsJ2xagxoGT7eKIk
dsdRhWg4sz5fGOb9ktNNLXiOnb9MPGj8/rQ7Dqo45rpxEKCMkE2xxHiWpkPqvVw0
7RQzucmkzq1Akh1lkKoHwUehL3iAF3rYfjV/2uKUMT2O2s7WVzQX516lkhLS8Iqh
ya0098Wo72+ws+erK6DbzkaEu4/r7lFBqoWtri6x+1Jn9ljjA/2poTZLMhPcxWwJ
r11j3YVRn6XWE6FZuELJ2PwcKKWFxBfgQHZBafqBJJ3fiOygiRgsDA1u9fIWaAfi
LwiBEL/M58qvVdMxhXGcaJ7y3b+j0KELH6b7Dsvm1FbYBgAjBGVBmINYfdM500ot
dA6dXUwvPy9Ybz4VlA1b6sZXBQ06BlhTiCd2CvCkxm0XO4+3McXJJ+RDjA5GDRrJ
4zAC9q3M0AKZhOOWIfWwunHjuascqoqARJ8vglaRuSgI9f09njXs+quxzEGjnTOQ
/QGNVD/dD8tfSmcO0Fy/pl1RHFo5JG2KIgyUlPd91LJx8iQOc6XT5ItA3uxWj6bl
g9fSQ2vsiPQBROF4N8DfQ1LSZWK6mHoRs2vbl+sO8Zn1Qo25PU/rTJhldG0uYqpe
Df0tBrMGCg357i+9N6BmJEe3LYUdXwHAhKO9NSKdNB3xMJJMyEnrQ3J9/OCaJlGJ
ndOmDT+opiwJSRRCD/JUkDmOagdPaGhXtRzVto0cxGBziBwwdCSD/SCWA5/BKwFY
rIjRCTbE6hhWq+tIRVhESFVufwvZUwejqGbnaaj5a+D2RDUZh7ZoQxJWQ6m19l/n
R8FVeDjZnYghRdM6y1P/xfJgvZZdJ0WJeuHbjADKSszFCCTLlN4Hfi7jrE6IqGC0
ZXqM3aaH37GzkrHggZBWIzRz++90OsOAEHlhmjZP+s2blBaQHXaiA6AbnFrSRJO9
nd7xdUWynPEt1SmzvxsD/oGtMsGjL9uaSvXFgqQBabh4on1qPseko1qHVVR4f364
tBcxapFnLxp2b4JrN1PdSHq+cnuHK8sOfFBbKsDAr1rOAP4JrtBs65lgjjiLn5a7
cCCNJEYs4PVi/hZ5IcA/y5hGCvCKlegdx2C1mzwmg0+GePib6CEJrJvab28eoxjk
/gWo1z4ltcB9cyyiA3I8BK5q25y+fyAk53P0P8Kzp1Lw86kvQR76O17rUP88zOQz
ojk01Yltq83c5FhTmISBTM2Z/xBvGLFFB66bgXu0b3/HSpSH8tbeTixPwOVA7ZfK
WwSOSHqS7e6DqZbQxULfZAs/CWL24Lc2RblzMbRQoclfavaYaP+IVS90ZsMEgXcV
HRFN5xVPcw7F/GmiCCFGFA1HGPv2TJU11YXEgGC+ieE/dB30Rela0RLsPrP3/pic
bmuBN76d5ZbIWEhpPv0sGFKEnDQBKGZ74/irJgmbhAL7bR6fwcRa5umyReyVqksh
JtmTsY1wty5BVIEJEvvKNl8bXw92dkTZEBJolNLoKX57+hKhIc2PJCCPD/Cf9HiM
NUXErZbwfOxxM290aAMuNR8tcI4Hp9CBm1lYUAhom0/SBUmQDrKBXsRPZkN9Af5k
TfiFBJO9uQLUWa6VB3TfGWiIVqIcU9VY29sLAH8mDAfo9DuRE9WcTSEEikVS8QoI
k3QGQrmuXBp6O9TJ6R5QeAOLDFm2LzGpVFROZQIwovlX7snzN1o2tb62CYRybbM0
RipTI4EXsYhyxwj0n5tS+G7jH1tEFvbxiboMtGW37GW3LaUc/FOLhvUf8Ck95PRx
dOGJnKGWtILzO8tPiDlEVmBM+w3D9VFQsvpeabilbZcK6HzGlEgJdRKCiFOdY2eY
wshvylc+cr/pOwiCf44C1z3Qyoqbi3dJY3cnEVp9jlFHtikIXQsurjZWZjNrqLzu
g0+HNOr3UQ5eYhNjydw8wz7JCoxzITMx6SIaiLQ6KrKg64NP8NTIqSt2f4Unz04z
IiS3vQvPkKotsLpZucFO+YJ8WWH4K9FFq/GwIwYtU0sKTLycbNLXLd8mKaoh6b3u
4Hygvmb3u6gixnCwunL/Ik0BEtCnaM764R7jwnVaxRbTw7GRXKbGXYav69Eqb0bR
IThJ5efUOgz5n6T7PuvECfyuMeFYKC1Oa2koKNlMmTCWYEY7QX+Gdb15nHttRz4T
LuavisT+D39PORPjydv41TtNH+YB+97LWlB4HaJLj+NjqtqFh4rJVC/ytSHdXY2F
4FjZr4nYSFAuLMQSaVAT/fAP2xb2gNdZmiNObdgOPtSU/l4HgA7vGVU2qRoqrk2H
8HkzS+tdXxV8qV7biD21z92rpe9fewpK2Vya2PWvjweZH1gU7SYDCHGdO/J4A1NZ
arQF2D35dsg5UNL+6OX5B7bNKA3RQE9clvcW/JDJKEkiEj/ZOpB1c4SLcbyes9c6
3zbteLSpPg8GCz03yccAJYoMAp3mONc6k+zwokEFccFGXYJuX5j7FNV/dB2ZK+tl
dR4TZb2n9JG/wB8MDTCSXgm6cdYs5fcOVwD3DiPfjw4IltCjZ3XT44a2pMtszsFr
Z8dQ4KP9xlT7LZiDP28YiZ0Ik2JAYeL8nYpZtmemmekc9gmValcK4NkHvFjVNSXP
EDKrFOpeeUYdtRG1CDrRI3qT7P2xVV2QuPcgBqoFlYdMvgEnvNEsZYsGCUTltYzQ
ebMZUE+FZn1G8TiTyu63NW3bxP4MLuSJJ9t9xRWde9jeD1dPUODaTLMYR7dJ19/r
8WKHHUcqjRO8ztHOoE8yYMFqu1hq9uiljRPBr856zdbWzydn4kfYTFaH0BQzRI7r
i5EcXVtWwEkiDmvJptpsL1QN6m77pDmKOD6MvLW3Q1XekIyYIOn6jHRwYkmkC72B
LHqIJ+y1Tw6e8PZ56rdTDjbWdZSAQh9EmH+rS6bR7AK6VIzn3gKCafxVf0shk4HW
jRWrZEfSzCOf5Gd044hwoA4KUMCuOTK4Y8Z2H+UME4EKuKK1mYwn5NcptaW2pICw
eun/KNi4JhGKzVr3BnXpPqJhDMPZN4/PRu+uxE2GSnyVVIoLGITev1E7BSfRWtzR
LLzuV8WpGgBPYi0i14LzHaQfPJfozAwKDWlrDrWg8Tej8KzgQhNjwLctcd8gmZzO
4RXzBtv7FSUsUFUM1hsUbEqRzV48wf9JbiwhFAGDUCmM1MorIsM6TY9Hqh2OQBVI
ERREkv15jZjpwuCXCDUCwuvgq/coI/qFMBgYpMVp9YjM4Fzj5VyKEPfFyplrShqz
47v8+9GInnCYJEm1wvxnzcr/6O0ShQoarNbdkI3w5/R7CK0DNVESIZe0Zq+1lKL4
vHomQ4AcDWZHbG+7kPGCqh6j5CQYzcSh4jkuo8dXaloXqPXZhyBDI+n6Di5t3Lup
tQicmDi8DzMuupvpE98SapnHI5rNaOE5dVSHzoZPyOI+RT2XQgq0DbNusr53l+CX
hS3F94pmM937KVQpnFfTOxq/ADfDZPfMKT3NwRHCu+D1KkmnABxM+6A3yZa3vDXd
PpngVn3ftpF+a7w/ZnF83kYCwMrG7q6HvBsmQMJIrotBfsagsp+Ln3DqBd6GbuEd
6o+XN8hZg7A1Tua369KPFK7Qpb2M2djiqleUXPCO+ULKqnJTxnl241K7MAgaLPAL
Gx16gIkF1bFUM6KQRNcKuXgvTbZkGQYofGQ2XChYwv3IYqrfcYMTf8KUcdm6cnBf
0ivsbdl2Ix1f3Xi58XXdCETdL0qq9y/MBkjNyNsz9NdiMI+vkFbQx0qNJr1F5Gmv
frq+lblAP9vomlQDAoS9mWxB9N1Pfjx945eM0TREuHGnxBAGqhyns2d15sFNnQan
dVXkEZvVa3D/tSh43l4VQavQVgl6NQ60Wn7k+bmnG1Y4rEYydBuIb4+hR4d5/oWS
1yqXXJpXkGPuVOmV+nBOYNkTH90fkuZ+/bCKrnLgnfVsjgsjHQlbUWNd9uinUDmV
VaowmwKZwzuDOL+zK4C2xHi0AkSjgE6PlvGjw8PwsYcYzWRibB+jCr2M3qfISSra
ABObORlRahln45x3ULWoSGu+ywN3ONKCLTpQdNAMLzhlzd6XJac16viWqpy3Wqr8
myn+2CyeLL/oj13oRUfqvlys49+LG/77G7Zq481llCX7hGfCQtX54Xk3m9cBKxvG
ufhhpKGTwv3dgSwsyM0S39595CH7oXgZ3jrrEmNPPxIPCvaVNZYk1W5UbuS1MzvS
b9rup8ScGLGEEFE4fyAshsQE5GRxEcuPB0HWe/2/IBU0k9BppsNKiWXN8AfhcvkU
NN42C27HFPLhqp3lm9Mo6G353x1giR5wYuSs7L55h0nE5b75IKNZu60LhPIWpbPK
4GLr3jPo8Jw9aBVCceC7b9nBs1Xtp1HlzysuPhleD7RP8HxFTR7mkY0So/ca7203
HvX04ZOT+i93KWgxlX+hKSip54B8WYlbgzRX02tPMfnpmLK/FnO72uUc7NOVCgLZ
4xQ38QdfyipeHBfmnUG8ToPq1fbW2wZv0qUVAqyKEmLKr4T87reGccZDfWfpXPLM
ch1tAkr45v2ApJadJ+G4QjwUTgbrcUPqf+Eo0RNch9e2jQvHGfDqHxOnrvhtdL8A
glzf4czpKeGzvkCYvv6JWfMcxEnZXUOXG0upKz5ybQt/q99WIl4zju5VidVlHm6R
2wFtWHustHplkY/f1cLh8TV49N9zRxXqCv4I5cA0DEfVyTXUBktAGCClES3lk00e
N6LMCbhL1ob3Qum3H/mRmwENPhULY4OFP5e9QoWTu0OyRnGSIj3WjLkNnDcEMP46
qmpSkXcfyhE/3/m5g4VG8QnnrVfckaUnp5eXwua5YxmFH2IHPZcLfMouRs7bWbRc
0SdTMP5Mk2VR+fYT3eDTzD61Y3g7bp1/+c7uXTjvSkul++rmT9/75Z0YYRex9d0E
tSHYxzVMLdZPbEmy6tHJPO5LQA53VLnpO//dTWcOTJnazsqykBAshf90gYeiq5dm
tHOoeVOow7dYYWDwkmUTRj3ox6JaLOimd0QrfAFnRNjkV1fYpVw2hor4JE4/hra5
CkuqkwnWQkesyxZh1wXiMtWom9DyDAJdRL1g/N/z2csfMgU4b4fGDbPykUZRkDzh
YCip7i+eIHPjDdw9x1j4FFZp8egBIzCM/qNw0vPKK79Sm6F4yO45gG8cvsXNxBmU
tkdZuVyBoCpmMGT7d4C9T5SX8srCLX9ujHwWMkOaYh/gavlwdPtvxOzLCPyeM6Dv
X8zfMtPisxqvyovBbTRPIZVkrUfCvYbQvPK68ztNLWuI9lwXa2RZMqyQ8QXgDcQW
5x+CwLHNFwhoCD9FlP4m7L+Lljd+cRKyQlT3Lrk/FoVCyOBZztRPQSo26vjv4oC2
c27lN0kpjZroq8SCDEPF/AICCSZLS3WUIx1W6FlJQRqBfZxOb91FgzJxcQ9UhNNF
FaEuRyMAN/ktcrG96C68Crm4MvEgsERzuoYKBEkMWdroPzucmhGuiziD+ufhhmaI
bvDdURutYn4wMMZirx8tYN60qnlgZiW6wEgua52i2REglDz9cl0/SLt39LaTja7n
ipDnvBUtxG280AHdfYpHvBDC/dW9Lqg3PWU7wXygpBxjOdGcuMGhqyfWbmnqpfy+
Bn1X4OHJnVrNGAGNeMBtjoqMFJoe8+IoG+iLq7CoC40u35Y1GdKaVCtnYVv9Ckpy
rFjt7NLP5guv/LlQM9qW908zsQ6pAREUuC+fujNcBB7jplqFcTfkoybUWI3iuTre
Ew8hyIc8KqD5CYl08ethxbEHjvxr6Q3CoAnZBjiuv46djv8d+YKYfEq/RpcRJoeE
azQs7yKegZnAB9BzhlogZP+WS1OVTv4Ht3jcelFHMfxJXwp99vhsy5DvZisTBLeZ
4PTXnzTKsm20nad+2nsrb4k0G6VZw6oaI+2qrenq6nYIrpcKdtRAQpEwktIBhP5P
BMqZfy3IRzk4MeNxDPZGyNqAlRo8cINTapUpCcgW8/EbK5BmgPmdCVKh9dOfGaaM
Iy5qVUluupdeazVXikBeEzsRjirRycSkAq7sufsEzTzxLPNaxCtWlXMm5vEUY5e2
wc9cPoY8vDrQQCD1kojkDZSg4eYB/3jhU18XzDbK9tqy5aO5Vpm7BtZ64M+iTCUn
NN8cMbnSvUkQki2J1jQJFpYTl50X6A/+SP52pPFGNIotKelbdv1nXEEP+HTZ1AQe
uT32cyArUab6wkCfcDoi+Luq41eoCsNjCLAFfN6Nb8WHzPwFjNm4HEAhLPkroIBA
c6NHEngoiJsPXx9X6ncZWdmaf7BqxhD5cJAYXKk99mdIzCxpujBQyo3fSANuIZeE
Uz+RyP72ziZV9CG2GlBcb9cMv7lrsY0iUQTQpAetfaGAURKmEuwmwdw9HR0OQ+OX
tuhUGKrclBNWx55bNxlxlzuR4ZmmQQDnqVLWSr6bGbMXqxqLVKJIWC6M57zcLHNA
MI0qCIIpTTUYK7n45EV+RchW27Tld/8y6gAcqBBYNwvpWFOiWMNDXELW2TSpQikD
Ad5pzcjmYlfsu6LRmeti0pOHTNouFZTNn6m1lDv776Tu8WN+/1wNjhWo6157SwQb
Jd1Y2Lqv54iGkZjA1bvIeeJCAEThsrziTDgvkmodFZToraJu0qoPIr6jJHoqxiEe
M6MLcRC2vbbSpM/G/Gmx7rhOlgAptVUNO5Mgk1/mDEm7vx5M6PPxUbYgLxLi/DYq
a2VbdYebRD/1M2DHPG5J49rUv6ZmdaQZvUja+Jp1TqVwm3EQqNpATa2W2pG4wSh8
VFlPNAaagblGrE2D1RZW1a3jsuxgoZw09slvks2DPMTlTyo1SjopRc+pwleRX9hL
hHXboWqr0TekcAHdXg7vauVFLlqYSetNGRrSGtPOCGQZ4xEFOUxUGTuARI4gZNRW
OzNXoaTsftMt5Bm4u0Vj11NJL8USyhMomW6gQPNQvSxtUaPHP46kMk2PvAkWvihG
pGKxgVMxkTalYWZYXF9XQHA1BUz2Qd3CFKCd0C6MUMSwyq3XaoX4LvfAyjIsJQzo
d5PW6BqdtdkxA5mK+zhIJZ9Lphnv9doga8gO/Kz+ay1DbeoBLfKbRYueAKSbYBQu
VAY+DEgtuL1krN8gIvJQerGr8Bofr8TjJOYDMf9HApuRsE4liBSypAq967620jpD
std0pAf6d0Kkk4RGLGmiSaX7fu2+SVPk+tQQDchawh/QBfUthtmSe60ts21R64nD
/4YfqYNaUudyQxRn5gUfx3BXgNA5CXWQcboW/Y06f3NcrJF2SAud6ojf9f2LG/Dq
spflvMXnzQitWoyHo6Mx+9pRo/z4fOEK53i63/SYgxPbJ7ZwLesoV5VCXmXqwYLB
RxY5YBLob/ciGjwgMxAjMZo75tS6ctBFM2l33M5WgJ9o50yJ/5+GiZtzpT5iQvQ0
XQToMJiWg51TLHtJsP3xXaAMoyh7AsBCWkvsdZdDIQJA9qlcrndsQqHDOn9RQEsZ
0I7l7LZjcuNMdGHRbxULiLG/E4Nf1RvUYmSOszWMX4JIcdTKvhanuNFL7P0fOhGA
l6+954hqwo4yOeCXTzOUTxglqq8jtqa3vBndJ+LJQrubsoadfxFw6eQOAdAyIP9r
u0fH5gVkUDiHcQpIssqjtdRJdiazlDqNwIAypOdNhrzNv3qbdU/8UhlM43uElXwM
BQWQYoWcUzHL+VoguueMDkAxHthObBp8hEB/AqcOzAF0IirMfuSG1I3saDj2Is/W
626dxjufVtT2WxF5SrCtS/QZpUBhez8Y0hNwPx1wmnTqBP2XHmEWUKSzHGuewq5V
MENUfKcnwCikXI4xbw1l9XFbxWz2s48XULCyC2IvRblcLcvlJWM935aDMeOj3+NP
k+6OHalycM3cvfK0uB5egRWVH+Bjk4ZNlZ17Eo+zN7AMkRiyt1vCgvgmj5pLLt5g
7RRpxoSTXcoGRLrJjOHh8QWMOHHdKXc/4zvjfb+Iho+BEC3yloKq6Ge02awAveTI
XZJgZ1g4At2UdNUeAgweYG+X7lyzVV2dDI3L3VxVml1UZfnZvUbklEnNuzIOfIgO
OvuFKwm11u5csHw4vc4tXMyJmtogtGjezEenwIuy9W1WDUfmSerY6KHVMsPlEYvg
ZAciSUKW8WvYeg6yiwqD/hUOb8VmpusFZwuMUlD7fGN502CUfyCIOA54sErb7nFW
OtW35iPPR2Lx/thqFjXGMo+OT2oMK5olKeffBLsbNk/C/6a+4riMtHDKp02NI8XA
ZTj3g6DKfFo7yT2WYprvGN3iBjNmNZaP6R9fSNm7WNR+ymPVehw6upb5I4LFSne0
S1gL11EdgaLBInJRbl6q92vM/H4JCgLc+Ma68qTPg3MqkYnqSz31VeMmqPF8VPfU
1BbN85+Xx5efNGItdAg2F5ZUUQhYnKLje+hXAfk8ubFIKSSN9eStt+3GLPTbBny3
43zFB+XXKf7qjaDxTMvYMrUBC7pu71GJreONjyVpncClQknrrvvqFwSkSuk7WeSB
jXaa2oMQHYiSD4WbiDpcw5dQSxSohS8PikTgylEXBYQjRaJb5smgSINGXU+WCcyW
7GOqoyrIED8MguiGk0FrkvPD/l6brka6t+ykiiwjYQEyPbXIVouCqrugQZ16f6G8
0azvmzL8sQFCmYaxMR/wOG8TyofYF4rODBQBktAF2T6IzX3cUpb4/QYTjnKocXCp
NG14OIScDlASuyOWEyLgTVM6vTdQ8LZKUmJQ/6Rjrw2ZKiKbi/CmpaD4I0M0MzJD
UPJT2lpuCppXMXmrvgGxIFh22PB+ARaj8fjnNhWTDBdPhk9/iwuPLCRzGwBsg5Mj
cZLJy1jxlORyYLvShdi1iDlG+AYBj2vQY9yWmgyKo2vuyyGsUm8XcgcwqqWawVTM
j7NFzWprR+sBRWAe4UZodShTgEkBqfSLcZUYREbHrIfVZc3AFA6UNXfsv1KaC9oc
MxfVt9bIeOwS30aStwqwEEspuYKnhkBClT3VqwLkW3f47B+Oe4rtfOhP7Bbgl12u
TSd1TLF6Y8VcKbNTgb+hhFbqWm7StfTbOy6McLTROPwBMxcSgEt/DidraFD0ZLW9
V/GlpicOGpHKyJMvzj1JzqQm2Y9ySDsMv1DPYxSWmP53qlZxaAeON0gtYnwhqVs6
dnFxb+z0Ny7Nd2WCXrH1jiXq9cjY+NwOXYPP53x3FaBDWpdpY64DnEMTLcclkTFN
5YnPjUQr+qCanROBriXQzD62KHm4mYQsl3Du8YmpmXVJ93CvmLT1oekQDcGwZzrC
YtYVm9ajXAS+nWyPCHpHhe8qkPnvnF9qjbwnpcHj5I09gZJXcABoIqI3NqChfpSH
ChikzLPNmWcwH5sfgYVsce90b9S/VYIQQ/OcmKRwo7Np4DPQb4lXABqtuvhWunSh
8vG5ipU5lp1UqQUEbUzsUChD+Pfr3HWpzDzNzm32CkNRczyAk6qzgkoB+1t8nCQy
7Q5an1Ms2VDMR5gA0hHmoiOcc/bamPoYYS2NTURoGAcQ7ZnlwGdzhKHvg9B1zFg9
xVMexkhP0gbF9RiRIMsEh48P/sryrvZcc762YjG91itEJfTrsSayyRYzJsXivyXC
rzuhHtQxHkbGqFvNOj18GD5xrOCH67XsegO24DY+O339cicAYdBpDifES8TFP2OQ
aS0GHyNpQ0jpZfwbLDAGuzgQ63ZWjCDBWICJaBIaFddixVNpq0Bu0XK4H5urDbIa
mOp7YNXVJdKhTznK8nWrkmojs6VAnhuD+Eu5N77VF2eCRJcwNuWvb3+cD0zv2lSE
SXODjvISM1GiSjNcGYY6e8JO9Z45jvzMApjlppvMuZA3maUPPn10FaxcgZIMth0z
fujBKltV9UjBBwA7VmTOBLwLKk7HjD+c+nLeiB2IZDJyG/QDnd23N0h0EIq+sNFH
c5cYZaDHJulND/PqUQ0Vp7buMLrUq3fwQsOX5uuGm334jKqY6cfPdVP2osEu8N3C
dnhUEAjN/Ywvbd/Uxp1jwB2+UtGgzuLaqk/zBLKX2pHP+xmidCO3uIo9OXZmH5wU
UV12Wf8dEr259kr1BNTsC/hFgA8XZeffN7+Sg3/GExf6pvPm30eHo20EA6PGiNdS
psK1jDZuDkRFobDD91seTe3hplopSa2jEPgrooB2aj+8MisXiu9jPzz/6Ap/wDUK
vwpbrzCZL0xN4ac8fQzoAY0vTS7/8lb1TdzYIxCeDCAYrJVzz/O92dAJ4VeggSI7
YCEb1It1rl72iFTHiFhuPpFU/lufZ5berYI/cdDP7aBu6iv5nsKacjGdCOK210at
GaRpjULMPnMVtKn+uU/4LjSzmAieI4wKrnydScNoAgmsC3aeRGHGlj0lNG+oKVnn
XKK+0ZhYvoE+jD4lyWaOZRky+onUiDhPD0/rP9xTuOkWTjwv0UzhUXMtnRyPuhqm
eAWRSzDpl0BfTgJkjIK0nKd744kWwiVWdMFRmiAFtrkN62t+l1fCTzK9o4NxWufl
w5MWop3eHD7mV1S1TCgCGhxR8+DYl+uWkqKM1TLNfCmPbufUARl0rq5faIzN0Dmx
V0VRI7VQowoFb7aAQDOesrsHrvOS5s7We7XLb0bwtPBlc9dUvK3nBzsX/+Q1be2g
tmzzn6eyxfCxdNl1XCN1K7paHQilq17s+gA1QzaSoGm5I9ibWORBZQunnma18IVB
QXtu+xa7cbwbZ+UB9sYL2NqLOdtREAHmVgi0jfBbHmrSD4KdoP3ae5EZy+FHK7Uk
H/1/DpZMFu3sM2NCdnkC3vllHshMYNiSkD6M3DJRK9dM0tbhAVQXIbDaudmUbOKM
jAJKV8ejauLJZFyL95Y8SLurUJ5kzk7K2BlRARUeocvWYajleI2lRiSOIfiXTs84
hX1D9DR6U3ZEDyNE5O2i7EqulGNJgemmvpvn18U96DzuHUWto1LoEnWfJCgyhq4c
5IvfMMFNIAa97uMNXr9bFq9C8UAvE9k/LRoGFPr+Z6MDrSdmMblJYjT6ksXfF8uX
3Jptk/OaJNwHcNFy+Kqsv/LkcLag1kzj14A6O9N3T3aiz5I0sZVIJmVtYFknk8Z+
l4CbaMxghq+Pnfio+cBUilScPQ85+R4HYEAidzIsmttJCjEaT9iG2H+iwZc2//xL
SG9IBE5rCg0C98WMQ+HTAGID4JfO5uwbnI2FuN3HKjX/ewhl8HSV3Lt+2dffGv9o
ePZ3/bqQnu6x9G3hXrtMqzBTITsD7rP1pq63f1GQTuGgOB9C11iE19ejpFrS8M/a
Pmx0dFMLzBPudwDYdQRNxFI2JHMVt5YH6PygTwiCv57ZHhYqCXcaHl0xGuKoilqX
bGZ2MaAaWpvk21zlFwUBjX7IbejSpvSxY6B2sRNoqcL43PCeliPUjCvjAw5ZTPGn
yeg6Wlm9lq1UhsZ5MiUKAwWXIGgFD8aWo/VfXBgVvSWD4UTUlmA7Z7YqinJc3f/a
B8vORtXO72G0P4x/YMrak2x+a2eGoFTd4SkgyTJWCU5B0VKILbe1trXfy1Hru98s
CH4SVHGH8ghDnaZb/+z7CQfHswYuZwHN6AwoePi7XL5WrInSlVuOmUtOPB/R5PvM
nVmnm836YenuedigbCWADsR+DY3+9oRkoKO+lLgnWoKIS0HxaUpsDsvVjJVGs0sg
SLcj3QBcQf4pOln+2WQdWxuIWBagk9N8dGl8n9MbAJf1NGfgDHjpv8Ahp1nbmguz
iXHRUrTwTCPFM5u4k5+2kvW34Hb3LfG0UOeMVOw6itiOFNPSH6T7GuB72pxmAYuN
AaaVz4aOKYjjjwj+fkSS9Sh7sV2s/C5D0Lo5hSSGuwpVRcX/vMRj3GIQO5UsK1WH
AFR2i3Iaky12Tn1strfr7ttPXzQZSnDYCI5IwrVnUM+2sTrOoBSUbTesrvwckGez
djiylCDaaJ3/3HQdJBHkg9cljZU6kQHeH/cFIKw/q3Yy7FzbVChZeuliwgRVEE7l
Ac+0x4WEkWsz9ZtBsMQGQlT7EJDQkbQnVrU5C2A6ZV9UE48oysSFvomzn7GcNsqz
7veTx/aNlA9+w+1ehb2LFNAhFhJYTUzC1tI7E8gRl4KTxxQbrwjM40w1sVL+SVQv
xKasRKtjfUcFXTb9Q12rnXYfrCltZjIxiNPFTHLdW1WM1tR7Z0Dvp8XA8nuYEVjj
6AIoNBbGyz54K/8hnCeLiip0Z/o62wUpr2LhVWqs+ZhUrDBL9qOh7pry4qdD0zk2
oZkrY/38nAst7Gs7bBSVAp4rWkmuSfzMj/J8tVFtEh1xNdEwT09JUCpcol1G/w0b
pRs9EDn91x4xdr6ZzszncVWZoUi8RGro0GId7tIm/Te3hUXHR2St+BaS1G6nzbCF
uqWFQyuOFgWK5WfAldvF6fgBUEkRaKzv03P+3EwE898HhidZbQqXzLbrOUSTOjTp
Zxa74GmoAcSMkbstwzPkK5dOR3R71hO8MYdcT2ZNSKV2rmdjBCb/vK9p9qJdN/xF
3x3ry/j5eYhO37KlcZGgUusER4TLmTIdi+I4itSNJF096X+HO2wqVL+N5ECl8xJA
Vih86DEpLBRtE2T1TnZTYmXrrwNGH848fVt3h3cAIg0Nm/ivCj9mL+DiV8dachao
TRy4tzKuvVMjRL4GtOQ0gYuYE69dp9Ss0csu5hdhijsXLq4JIHWnTBJYhEj5lAY1
QtzbWRk4xku1DBF/VsN18NaGk6gwKPqf99Apvul1twzLkVnkDtQesmuB/sdx07jj
7fv+mTULbz4Hez8otw2lwI14PtHMGgx6c7jFqcDPvzP7witVYfOxZQNVAcBgoQav
vMMFt5c36XRASm99Iz0iiOupDxINISYPdoKBok0qXknIRWO0GKfFy/d7YQJluUW8
dmiWERQZq9dnVzCA+K11pVu1C8QvmcUEsQGxOt4nkjTmPhaGtRTAbSmj/No4HFnF
GTZimhdhCBJmm9sdqdWJ+8r0oG6fQ70NefRMu1huJJIUNz0zy4U9FTi9PVEMqWHu
0WVVS2fRCqZR3ZAu/HHbXKw/mJX9Ra47EEoIJiS8OGIzki3W73xc/bTy0Fwf6L3n
N+vW0xqkWAlg6Y8XhZBh1CX5T01hhK21wvUPUu6c2riO6CPUrIghmN5qLAqbI/XY
2o6ISYR1b8epEgqFMMTSYd4we89ShfnnR/LxBTCyDgyYwVWhaQlARVftelBOsZVr
at+zplUxq4fC+VfIGPS36San6smLoHBj4+NjzRYXYCgSTNAZHJt+rGrYESCC3h7P
or9Td3ohaFAio8fNJxzd86uV70chIjujxNWoRxWHvgBybd6CW/WMtEF//R9dADID
P55JVuH6E2xsBDIf2q8C+STLl2oORLmAZ1WBgR7v5g5PFjc8MNpLuQvkR/9j45io
wxbLyvXWjv93v8JW6004bP4QN0oFfSzTsqwgVUtfy51Iyxt7ZLnOr+ssz0gpH5DF
qfkrvVPK/I8tLjqU5gp54KR4ygZrabef56L2REI3Rck6/hkYzpss3UmE/FfS4K/S
bVoywRKnfsfF4W6rdpxoEL/KDAtcF4kgsPdsAAacqLxKX1C6daU+voNrFOg+HpVR
e2CVviY3iVjC5kpMEU8nqj1SGcnhiAOHNuUUTyO4UuGYVvaGkEK20q0AzQPDeod6
QAn6NXOPNWdUwyEHrD2NxVpYnR+edoA78h5Zb9NBtoLb4sqB9/xdirVv0lkDvz6/
dhHs7SbVr269XHY1en1dyF8bf5ivRxtfOxsd5rHaNoo+1A6uTGl6GupdmSTMhedu
bADxUyhw5LDFps0dggyn+To/viR77ePjQpIw+VjcfDfgjpnu3fyBkFCFk9eauAGX
SW0cFj51QT8vk47iLJF/JI7+NdjlPjyClw7A20d9S3W5tQEc/4pkaGHvnqmwWAwd
jwsKqZnFktoWagJoEnwVVCT8EIu5/feo2z27omuDEwdPaXW9ETDQ/TxRm+bUdwzb
JwsbS6kkPGyd55RGp/TZjhWRi6XOrvSK3L6kmyNWcBzbgZD2SWsVdh7RiHY9KcZ+
RWtst1CbeWFWb4Ig9kdC63HuTSg8OLAXqNU5NBJt28UTbpVC2k1wAvermRUDGR0w
ObjceB9F4l+G9ayMDk/S6BGiVsw3f3RwVsXTwUj5wpW/t60zgGR27hGTJ8vvF7t7
m5agIbI0m4PctuSt7zlEVLZcGknrSl2HT08Mt4NohdyYa7XdrJoW5BQfHqF3R4rG
uUTTsC8ImEnnFunfHEUPzqwEaJ/zPYE1I0SMZLH1bO8dRN4zjJ2acEvDSGqXoZf4
eoTtHMXDJvOwCUh3y1HDaUFsT11k0GEQeiLDT+Q/Kulk5dVE99E6anFQFAyU+Tfz
Q1wRdPRdbSu7jgTyDIlHaJpp32yPBbxfa2z8HLsZIn28ZeJ+ehTcrTWTXk8k9zxu
A4vFayJhX8t39/rUwKXW8iSWLpSga+EXhK9ULykFVjMQjSPW5sctJsZBi5VmcVog
C+Cy7qtr3l+L4lMzIsVjDIYTkrviugQeo4tvlrH6lAEq5+dgXcG8eJjkYzUXrtzg
i5zBBNYbj/+0ptSRZHbkMqp0NW/sS56iT+BoZhjAUFw9Dt1KkoOikOUoDyI9KE7B
gFVC0C1Eav3V3F8fnMV/YT6gLMKRq0Y7Or0LlKt9uhU1eYhZwvtWbBA7hthjuPFR
NPbpLWP8YJApgxmmpV8NrahateBhvpGzXRML54uErZUks/iU5Mpu+3JlIH+xiHgH
WhUMayoBVjOF5MlUo7xIxSe3suyqkv1CnJPXjsDYQrKzHmwbeWiMbwicbWZqSieL
aEkqH5HDPwoCifutTNc+0r53LtMVPta9z66Y5BB4aLvP6HvDMSt2mqV1icZbf6WC
OFyUQxZfAWkarnyaZkeorhHBq3qf5bcUwaB53BhJT5SDVXDSUO7mbJi0E478QQjf
v02M7h0G6fMkw87O32czfaZqKYY3VLQroQXc9hyEkweCwEDVA1lVMvwwlHUYfgs7
ghiJ3VvrMMr935p8NqCoa8zpN1iYP+zuON/pCPNE3jm/8phl99Q6m4K/eM8/LWN0
dHiI7vvO9ySxxOzNa+fq01F4SkZt44kbMoQC3E+B23SbbLdqeO9J8ss7ETIBYIpL
eG0IJaT8/345pp5PnOE5W9dESj8YfsTAVQKTN862cBCkeazUCrmf2E6D8aa+2VV8
7RI9qHjX9EGPFj00K7tAvx6jW1gTccF58z0XXJPR9Jofhm8qGA/rIwnVo5QoyWnf
5F7Amib+uZN1JElmPsDaWqZbXbkHoY1urjcBEU7FAg3I4m7auWtrD8K0omLTh3kT
obRLJsuKZVjO3ML9JuGusFoYxITdho6G+tq1+p61ZQb8j5wXpkcKovQY2Ag7K9wD
eQ20wyOQHYoEhxxcStekaJM7UfjrTbcWfwc3FKxYYYqwtjjSVv3CZNRC+5rmX0TB
zUWE9vcnXqeJPP9Ynb53B/99/yCu3/MiRDZEdE1bau5eGkkv7r0+jzwLG9Q31P0o
cit7FA30QMD0c/GelKc+hgJmdcQAs+6ZbwTjes89Y3R5fvXMwMrh5W4DpAVcHz61
2fD6vqmibPc77EcQVS0nSTmXEannFnAANUrwOltUyJr0+6CBTGXuYHc1myDcosfE
260+nfN0j5ljVnPll6ouWfw2ycir7iltXt3RjY9qX96roASyNco43C5zh+lvJc3z
hVq8+MFO/TgYdnT3yYppmelNyC0RXwBBfDyNY53vw8iFLvuBiOm8Eif8uyOTtdJp
ArsJn+UlsMxtoxGzxnUgJUc/4OJGvjzhP1XOksooyMbKO8T6KMrbsfWEtn64NfxM
1yJ3z2j9uW+LLq9p4UdsAPMN7aMEIkSiyQJyjZOrFAfxlmOfS/QFDbigyW+iHEnV
8Xwl6L/qT8TQvAla17Lwl+SvQ3X4lRWTDk/Tth3Zkt5c86tZpesSmmFqqyorzf/P
mfnddYaKNmEfOyPI/aWqASjuUa+ArAev62CMG2SAARYSloUj3aqitsecQI1cZWbs
pCopIC+dKU+1f1DGMhVVJ+xi7TQwmvLrX3enFoVJUP+A160fKoq26RPkDiq4pTl1
/54Nh8dulNGUTr+l0vsTqpuk35fvljunHFksjgo++gStdNG/Va9kZVUXOW1eu4Ki
Iu6NspLnu6dzBuoeKWHvnNMpGBZ99FhsA8xxbjE177JQcc2uWGp6RIPH3+s7OZSi
f3rqdDHuYa/oSZOOOaLgW3AjxDn/H0wfppKDX1Q9rOJ63mW/lo5eu/vEj3Rjv9pc
DNgfMOUNj9/hRlRpbT+gYu5oWx/h+o9vkCVeigLr/u2sLkDDX0lzjzQP3/C51kC7
W9s1dmsbih/ZTuo50mdJiUZS9TMxXa/Z5W7gh4zkDcJL4vOhQ89PdBC+iYZ1E4gX
jPtxBid8oX6gEkfZ7nWIzwLaQoSlvCE2R+eyALCafFm5fRO/aJB988XO7ehvlRW9
pe3RY/u3rbMNVMqpRvEC8eLPoo+h3VWN2GDAKI1L09MMu/vC7TndIJWlYqW0JQpq
Kh1rZRMjydStVGelDzo3h2YNJGSmhtBg81tDj7Se+kSmFO5XkcoOtR62BheTZClz
2XgLnK2BfquBV2S2Gmmd3HRRghO6WRBnPRmfANtgQZZw0nUohhvfrb4x4V02e78e
2QKiYhqOt7ryFUzW+eQG/9Wps1nTCACxPWU9N8LSJ67x41CZNIDRYu07YMUp2y4U
YXfz2MZ5Sn6abrgzlIbNP8GHLssw6yl+Cp2sYC+3JxCItwElyUQn7PO8tuAorr8T
jvn+kdN102R9Q25MHcVsH4kv4u7aOLQX6cNVJ00S1BLbLWFRbEkyCGwBr16XLN73
AacLSi05LsDdZuipBWqzC9nRLV6xQ8+7gne98Cy/zpc8v5OT6W2bt/FqlKT3PcZG
jwx9vYHDEbKCTUlQ+LU6YIOWHXA0bzZ/xaARuxi909rn3IUNID6CANen5QHBlJgQ
h/4/u7YChlNbrGiz3x1VMlftfymHr6vqKJH///PnLPPSP0S2l8iQ+GFuCBcdHoIM
9GYvZ9L8pea3inghQorUNQyBylqyMzt5nhV6262HeTlBZvonD8WlxFv25tC4Hwbc
0zvPZonMelvUYrCBpBBYLFl4qZvyFn87aaACx1NCo8JhlWThi0PbpiDMq9UPNiSq
XMvWxhZeAhKyqlKlihgOybvR3/ZP/+jrmKxOIzv8BuoOQebY617kbIxERLer5OBE
1wdIMnSpXV3mc/hGK7XchY5lw4YRGH3MLsWvxlfgi3L2EWqR81CbOwX20j7S3TZG
Vawlvj56GNwNNowxyJBpL0wGMOBvT3ZU3HyAqdh63R1x5Bt7wS298uDOZf/Ypctm
v1LDQT8vm0NpzhYJE8QrjCIxPCOrBIKWW8RM/qJB5DMIwU31W9t/zuJAeqf8tquj
TYdWFo5AzqICvqRUDAte3ryTJyaaM/IIMIzjUaTQqkVp0HCe75L3ZAZq1GUzVNzy
eR2pfF03ETJRNrpmsA8XqATUw0EGEjT1058BFC1yuposIEbScjkymaCP/fMO5T+4
4xdU+fKHhxojLf5ih5BOrU1olGXBlRa59uFkxmHdN8OqC4QdHGNv/doMcNBM7BbE
6dSk77M4vuBepqLcImzNAqMbdgAihWeWYk0MxVYugIqp9WpxbF+C4/MJzFkkTPnV
hKgwSQ2Q7m9P56rVy/3idjJRhkyk1dJlLaPbzyaDxrDf6toH1JNCkHddgqpceG4M
eOMy4gOuBR9jf1QI9KFjP9mdBLA6e3eiQgaJUe1ED8p5tCX26ILybMT6wXY3dHas
Drwbo0VfX4Fp9vGvlgHBaMxPSftgNv3VrZftiw+9Aaul1UIwT3ZVaRyH3iRwEY36
B1oRck/iUXmp1ZxgWvYqcNcbI0Vmmzjts5BHEGaV4QA+1d+brz68FmHDmOV8NCUd
ZC7waDDQCEBe+AKjanm/AZbWQokDRX9z6Yob0GG5dkB98V/jUNt7VUgGZb+RVF2H
IAqlsLhchBqblJTwpLus7D/No6aGMCDt5T972PYTNxAfv0K0cvD9LgK+WjLrb/CG
5UArlRsFBuezZ0RHGOgq0GqvwPnejLDcek5sf0CxJKpfkEPatkKxqwLVXPSRdqhU
6OC43y15PQpV1ZRCGZMLQUb/W1H9W91F9JCuIVTFzUkJVy3XaBYHe0X+0Oz/3YB+
QVt9D7OqgZaYcqkPLp2IqljaGiu5wc6jUPrGTn6dTnRbwtIJqBoPpqT8jNzIt2Mo
mtrdSVG0DjXAHof6m1pMffxTClgQ5m0Udm8rrwBLKCJBL8SS+vSdTBVoI9K5jHoP
3EHIBbLb/VE3BpPn2OZCEMZMJk4UobEf69zBvWJe08L9a3PJT0ED1sROEiCaFrI1
VjKn9eGBWuoE1+JKXGY5eaaG6moTpr8cKfEpLhesoKtaJVjWIT8OoZO5EfQz8Iww
bt1AGzDnwkN7jRyjCOuiuvC02e65tHhB2vaBk+mxXz2w2pz0z3jqwQltVLmUqSY4
bb1WfXC7DrgVd/f5dQaG1Ue4qJYSg0FfHlELSDc/KvXlGEr9kEMZ5gneoTiKf1xy
kYgaSN/kL0/+PHgRTb0tjvvnAIxozqQ+qIxTwDUk9yq7p2Mo8UvL8C82SBo10tGE
fIb1uaz7PEOnvXIgl+18sQmKjX6Uwlb4VxExZnbLpao49RutaGV3ev/2LGyqnJLT
BiBlcp3hOxJEcqBmM3MDEzVvajyD8diIsw+sG+7E7jbwkJsxwtG2jZsdp2Cfefgg
ac2tMwrTJjpTz4sZ5EGu026Urrt3b9ZEGnNpf/JODKBZOTLlIA4BvOw4hJMH2OpE
kh+6Y350UtmAD7LT1MMIZogUltc9b60ZOMil7zHZi+kDp2FFpbVsYR6emyGcSUN/
YTcZFmPLFFBf0IVHr/Ev1nYPMKXHCH/7pyE17l5Qdj6hGY+js/BsYJ4jTYmD1Or7
Yh0lW8ORrPIwutgVtFvLS6DPKsjmgo0+1sHOQOE8Nf4OyCmEgZ8xpVgdgwBx2gYi
NRTKWedEv5vhbgOfhveEYsbloa0XRNXrhmO8FBl00x5Ew9kZNce+KuZ1xqJWbCPM
cFgaopX6iULLu/Lo4KmPxPHEbOgYP4WbMoWhfZ2sanfATJy98BmpgRCuxaEr9Ff7
vt3p2r7FhozU1szvD5GQ/Ucj9aHg1z94LuKOfnKZYMkF9GDWXVD1Dg7y2qvdYNmt
ff3om5W5OUqoyGhciMb1LQoCK8/4pmCcRKJ7snShek5U3IWij0SI0fn6Kfi/1Gdp
dUszjm8GHXcz0jZKo2sS464ZjU1/WYcvhESm1X8i8OqSwqV1ppIO9tqHmlCQk8eG
GhP5eipZZLNQFQdzs5RBNk4027tP7+468/QBVSyvJGtbjwphRVtAiWR15nV/qgeO
af0WR2Cssk94UnWuRcSRm9BmwHDMmkH6kb6rVmb0CUmTB3u/C05dfzpnOj9noVVx
70YnEIt1xrMnx8Xk64uIyGaov50tY3HA5bsBgfgHgqTsHKZQUGfA8aBAdtvBZHB7
WrW8LN1gvNTWb4LD845nttUnxE6Xhaa3U7Po8XDpRUIGbdgj/dPSmJ1yJgpNKmXk
sdZkbkv88ykX9QEY/0IWo/O1P4GznQdPPHplJjJe2+cN82f3RyqSUTIhCoQzd1Dl
HPp66RmutflqFsQCThp+ZnmHBy9WyjE/0xm6EGn5zkbUL+51rJ1w5+OfYRarDPWi
d9OAmRwWUSIEW0HK/qxPcgfktXLsBfbirh2/bySwVKz+XB+uizPkXDlBAB7N/d2P
0a/IN5S288Y3M+0cpGURkm+0aERIjaF12L/iQ6P/S660gxyeRmihxMTZo6AdJKmr
YxkUsQaUq7OF7Ow459BMDN0eu99P7/IXlrLwQQOY4OcAWOiFl0dwwc7mlsTGNUvg
MxvbOqhJn9m9h9UVA13sJlLSsfa1KOgjayVAM2p+mURJS+zzPg+ONS5WtNEH5z50
O594CK0IKMllK2qx4j8hJ2/MQpCNaY6pp08rQDKR5jRaewPBuVPhgtjzMMDsxfgr
/s4z0H0+OC82ikBUA/q2mQ+Pq+nLhGheWD1FQ1SRBUMaiWn5AYzJOaUa74YLgogC
6myTYrikm8tf7cDqkfc/AEx2QLP2bKDmY9fNYR8AzezHzEVVp8R2b7dkjJjA1XwE
LF2RjOCJC78qAhL4HkghNKzdPwB6B7mQBxCxOZQcqHjUGeAGGqHBcmgKBCfyN4WO
3uEUpF362229QtuB7UGbOnZvFc3rOBoM6LAOW71XJwPttw9Zr2y13fjFQqtqItjF
QSt3b7NjtcO5ZvvEfeh4KhFG8IHpz04fiWfietVOWzaNjtWO427BlQlht1iWSso1
hSrj9T9dEATLBC18h0L9gS+YsMUakybZiS3wWNs6TCNwR5Rdux72Rft8UohWu5za
oHWUT7uRWWXrBf6jsF0IHJOwUbMD4bQwgCM9lKTEWkeIRq7zJIJWJ2civiP3yLZD
DjYH2Ozy85IOap4qcApdjba4nH3K82pzMlWD/Yi8ru1HXeAtacI03jSO25BuEGfE
LSNC8OZ357KHwrbDBIfZREJ782oVMZ5jm0JQToSLq32EYTApOmjIAAZSbQHd2dSc
u5x8iVOgtBAep/9sYzR75F8HiJuh9Vd45HwNsoqKCi/lbPgwKl6FHORkb5+LOm6Z
HUN22tZzEgUn61HLtPbHmc4SZ84uRuAFSU7rz+/+cT05wRb9Qrua3bxgZsR7bUW3
AukXAqmgYh07zHTW57eyZpHwIFbJ9oC8lgqDpFIWdCbLu3FVXKgHjRDZH4SvY4RQ
zdt5uKRN8b1Pvrf6KoqSovdAemUWpd5AE+ecsu3Ji7lLaYJ7xhL0D4wnodtfzQ9K
R57QJjNtVrWSae1jW2rY+vE0ufQVrtsT1PNStTKa3iYu88KDZiL+AfFNstK9SKpQ
1qyM5yMNfu26NL893erzu7xaY7tzhN2+Cc7LdnMGCnEJrvgg8ulPFnBL55Q/qJH0
aFV+pulwYp0DK0/QBxcj6wMG5Ep4SYJ8IWhAJN5aXIA4brdTEyWecPQGdS9AHbbU
uJhWDXFw4b8xn7HgwHLx7sKNvJHkXfhyjUudEQzl6hRg5VHN2yKV1xWyI8y/2UsV
Yw4Uuq/whu+jyx/CnrFGpYXucmWM/5XxP3tUmG5Dzz/utj66/rbSzoKRDgN/IP/y
0SZqjLgrb9sli0LFuxaWAxOR5k1i/oLvO8Sqzu5GdIPVhk6g1et0myoRZJNYr9rm
eYPG5h0U4WPkSQtWjMxyFFAW5EmCbHgjwQ3Nlxw0LermM9DFm8aSSEASrJtE2Wcb
LF7BJMLAriF52PvyMclOvJFsnVGDkZHv+EDg8fVLP0FB8ebdL7t0PakV/bK7PdoV
mbC2OfjMu5svJ7li0+x12y/SYhLViPY81X/sNkF39AwySqLfZaLdrnTsJiDXNKeg
6ajfv1k4MkzR2JoeOcryeb+sa5+rh1lcHi/nayjjknwyT0HEmtWLtUI9ceh/geHj
qwLgTf0kP1lu6cPaNxvF4GTtt05XjeLD29U8o0kFcg/2D8xjj7inVt1TFVe+pzP1
zN6sN6i3Euvl6NHvwfqTtGj+3AHBeNlHH66dhZUFffi8yiO0zkqg2ayav3KZZE4J
aF6It560Xes3WJj9Xkwi2dsFA746CnMS8Kng+reZvB+YKC0s7Xtsy4YuziNevoL3
oWhL0naicptFRDSkEQrJssMSDCr4jt7aUaWH//Fokdonl+lhSFiJzdIx0DkdyXOi
0QjxN263XLbv+Y5qtnQiLvvSoRlbjiL0X05+roG1/UCsNX25ogic8EoSUFWL8nJg
VS3vj0F+NaGcVDCVP7owZZ2ss/MNFXTOoFhtwnVk/dz3c9xE/JgU0H3PrrlR7UGj
W8UFguVZKxdE/pxfuKJKhwnUz0Jj3B/5+vkBfE1CNuYHgdfbhJNUSzqPIaLbIe9c
MtutjcTSFd13odQ4x0eDf6XxTVESt2JR7VkNTDXNCKStyxk+KbNorU/71TiaSTK8
9wavrGzldd5j9BVGVRJ69hZptoZcLqO8x/g0+mvZ64VPWVr3gph/OT8L3yRFdyhs
1EPHBBulqbqILxVXjoNF4syvha4wprUNNOrGXyDjXjxER2ijLeFesQ3qCQZU2Zoe
Pvb0sEbZu/jtFDug+4Xl04pGgHkR/N6kaRl0f2a97xlg6sy9uICBpoe39YyNsBGK
foa7wKfxN1OVk4B+37IgDxRP0ucpmrsZ03aFnkH11wVM9f7VUCoMuixdMbk0pjXX
g6rQDqVRJAgerBZeAud5Zy9ieeo95f0LrHDVP8t+qMhjBhHFZ10omOn5/yitcPfr
FmCoKt79uoHFJ3PdjN6k61aaXIRcKJnZT7cvO2XwoiflVnRdMnmTHFVYznCno4B8
hQJWNbDLdJd3aruBALaP3hKR4wswXC3AVKtV9qiHPjE6XwyXEiMBVwEpynE/Qbis
mmhHtYBRb/MjIk2Vk3tgOyTCCj8PLR5MKzIvbjsPhxdA60mHgOYTmFwfS8dTV2uz
/wVr0xintsFfw79zLK1o4sOCsCP4asW+jR2gl2pGjf+QbbrZoSIvMk3vnEl2dfX0
w9p+06axerZSQsXSeQy4jXfnbHO0iTiXnhRSHHxS52ZyPufu/V1CAzoDvokDgED+
8nIdUayWfFCMbQKaLJt+NzGD3newbidnbThjOqCrh4bWWKImbOHBnYBKkDscfbJ7
wTiw7dBe6D5cQIm+ZOQ2W7MuDGafZaQhAQ1dug15SqQEsHcUIPF/7e+X4BzGJveK
MkAcUNKPwV3KOW2cMPZZZ1UqwE+iTDpF3LimbYOD6v5zQZcRLzDBkCWVGF+oU/Af
1ekIugTcMtsKhw70lHO2vX1T2ErT3pJauSjrylwECpVt+XD7/pvZyTZaXLXqvACh
suS7mmOIyeaQr79/UdcHuw/tQtcUMyp2M36tyO5Imd2LiFjcNGZEFSz8X75c5hF8
syzMp/8Ox0wJrK+7yHj5ZGLJNQNwdXQ5UwzN4kA4SWi/E8d8jh3zOUrc3y+ID41S
ACEZZ2Ir61iVYkjlnPFhJ3sxyiM7/IJM+DtCa9/110sfIFkPdZuRLXGx2WHvlQXw
IKFvdau8XeE+L0OcF6/ndW0mtQvWwg1hDi1QExs6sjGGr9Y+rgyR3ZWIGwei+d7W
QR9Wd4TAzBE8yxMRxzmtLjhm0lwqEqy3gvD7Viiij9Nlinq5BzUczN+QMs3ARby1
6p+gG2meOLiyAg6AJwIybO032cBNZV5cR6zYh/yT20sTuJZLKLpORPb14UwVUnNB
qoHMQXCLqbjQMW/qRa7wR3knpZvbUVas0Qd765XkaHqpI+teVTZHHiTO1CVPKAEU
EHNyIkbi09xAINAxFxEdzHW/6IhkpQkQPYDzDIwMXMktGcJDX5+LcHJmEcJknaf1
5gbjUs08/diNMz540EXYt4UcPPAImHc846IHhqzD1zexRu0BAfNrgtsGLImYbaV2
ZQKw7+8OuacrSVYr55/s/VT7T+5StAqBHkaUyS0tvHHo6JdOOv6rRIioRKz9KSWd
oe+CcCZiIWdMAF5Z3MsRvtMcI090TDunIOvuC/ZMz4N3vjjEaxCw2GkEx7zqw/pI
HD4az2WdDV72uUoYZXlTmUBfNo02vPkWoNwpUhEwv39XK8BwMyvTzpvAtsa/zKNQ
aYSFFKxDG4+JpaexTSnOrhIug3+Z0zH0gVNLp5nsWCa1qQtlcw7Hm1fQjb6X8gq4
KSVZTsLTN8c/b4eXD+Ah0h+ug02HRHORvkZtz8wXvrCfTjK+OUxPTdNBT5llr+xd
ktjDXQJhTT0BPDCw3QsSG9dPMHJh/4G+WoiMPqSgYDXOnzsWy6HANOfGf8JeQ8Gd
3X6P9LV8k2hGqGgXO3B35br/4NCzkUrWKe2AQO7N/4AogP8Q50CJSsbTTrZbvirp
yzPanOsCZsTPf/RkM6WjsI8vW2p9pgnM1WJUkcocduDhLOynSY2R1XD492IfEPtX
C1xPIXeoRJzqDVBT2TDUp+zGlnbbzOxOMORTdqdtTi3ndlTdIWI6aCh+W53Ltqmf
ZvnbQPEbmqFEcLRhlInG69QoiMVGaBgz5laRgI4S7muDNtZnOCA4qeTzr236r6pI
Q0vcscYcEv/hioKfvFAeLT1tEymVjd857sOExJmS68zEZUA4s0akEefgMxwBqtY5
Mlt1ecYvCoaoluQxoUItUBZMmkaxd9w07TEwXEWhkDujzn1RxfWEO9+o5EptbEHf
f2Yh0gOWoO86uWZ5pr8f5wnNnkLx5HCG3YHDTqiJrH7lw6YvwOpRjA/OD/0Xm7fS
2JjF3ANnayBz1yQsiMvzS9pl1tfaq9cWVHeGkuAM0PA98kf8ENclO8WN2F1gf+KG
4lPUq0VSj3HlutCeL/GFld8gxo0HJLWe8i4PUtVmHwakvWFUR+F2ZUHQllF3XcUW
l3vlc1N5ICa5955+gb2cS7wt0L5XZ8mY1xUscs4ELRLG+h95uS95PMD5etODnuvZ
z+kiyYyhcNPitO/v/ZFo/tzGWRQHGA/GDdTbOwU9sjgUQZwbbeRDnrhmLuud7tli
efXDLYwdDlqhcT5rVubpWUTywVynBg2XT4xGuht+LhOy8rXAaYItmQtjYd4etrML
BD3nAJ+cr+S6cR1lscC3TBCTS53gSst8gWEcWU7NzUjsfwUrRLRevQ0m4b/ExHvR
URtINidbmK6Wevn4WtsiiF9fg9tZ9rX+gbh0JoFnVbVr+mxxUnV9ssHKIUXNSWdS
TrLmxgdE9nP9LaSWPYmyBSZuBZVq7Zu7arNebJdGXbMjx8Zh3MWjrnlwh8ByFb63
QWEaDZhszykL45zh0uxFO0JeVzSvUcNNVYDH7JXDCeTkoxPgzuXwe9yLj/Nhq2cE
U0J2RvwVRJ6QwkXc7kHjO9/NGMXklC4tO7p5192nmeKmw06SL3qW/LOlS6GeQx+m
fjASZiCNwWoJ4GAycqrkR2rOupihDQi3OyUCqz5qW7NMRbshMEWxzZFCwxrENicm
Av1s3B8+8XlgZ04TneIoaEZ7+VH/5shSSMitlmpbpr/vE6Hi40B3eC2giNVC3sdM
WMQfVxAj9FHCw5s1UZPICHlR30v6lJ/I/LeG+rY8KCXrmDt2nidrUloxZFoZ0arp
nUmk743b3r6YGDVIVUYnletxPI6fkc+slOAJdQzYgcYGfTeaVfrJ4iBVemwRyA6E
naHa5T1BDT+C4XVUX0v3mYpgy4xXBuHPLq3rKLFIKsGz1kEwWNvHQUDBjwfb4S5o
x4wHiuUjlkj4NlCFG6OuVnL7tJQe8yDaEO8T5U+bOiGVg4aBEIPcymE6Og5ggCKb
fncnupSUFWioyE+DpbHcvuBX15DE8M0Nc0VDCiyy09xH71IeG2+/TrrEVdQVVHsP
Zr10sdZODnuotpwv3vZl+x3iwvmiM6ypDUopVMQ7RkGwHTDBwF6iTpB/ZlbeiTam
vYv27LRHlIwDdd7CebN0GVLd2XerCI7nhXYMyFSMo5YztsVI9GxMGEbrz3KRGW22
6pselof+N648WHRGVUNnCNssgT9hu79GOwbe/l54CrfGgzB7DYxBWX2ctL31KFgo
12Qy3K2gnnLW36NpqIfqb7DAcgZtg1l2IdFCe73awO+BgRaTlxrslOipN4KOoRNQ
96SEH2ct3xQH+KLRg5+YPQR0MSeJoG24yHQTJ7GsBanRP/vj5wquaOzVjQTepZsT
/J5lpwXwnYbHizGl16JlljL50phc0b5eickQvIzVEuYQQ6Gfh8oE2dzrAXxmZd6B
x5gcU2poQ7aNRPV787WiF2Mw9q49f8SyLFg/lmDSZmMxW/hGpAz3z/l8G49zdrvB
uxZZSyRH5U06gW8GBpqWzg0TeCNpkD8ydxm5p/O+2R37JO/oaYRMdg8s69O0Afn6
3DVTVcaYvBV+v1FwsFCLsfCvDIfEEQ+ep3pFfa/pCM86OKBKjtTlk4l1o6E1aJ9G
e7wnBbECilMzVGGl5ZrSppt6p5ePqmFJ4sUk70NAmIlac6LtglyDDu6bM+JHfdma
FQKWd+598ryFH3Y3TJ4R4TM2nR8JMjyIt8PoV8ik4VaR/LztvKEWq8rh5Cweih62
JIWIipRd3HqNxSLMrNCssgdKfW3OPvR6SKGJMZ1fkk63Qwds+wQN6ksvCPNS9n0L
fDI0LpOlndnqWPAxl36oqtBi1WOWHfB8dM9/MHjn58pcbZGpKo3AaaBcU36++01v
bdmOUlQMrC0rNUj2Ti7soyPIrdY04DZu5lB3mCTKhBN1ngw6CPU2uX6z8f2WMJWv
C6Bdl4UQH/zbCdph+w3nQdwgzzSJiDdwjWbxGAyAjkl7EZw8XpTi5LVn18g1wSrx
9g7rXCeh4JFNvDkMhLY73YpFqLenXtR7vm6e4tL5hBcVje9zWB/LRfpgCRLXWU+Q
SvQKRvQCF/XC1xU2zMxyml8fyqK7/DgJ022FqDEVk7Zn6l7Yy0nm95S63j4sZZAo
eaed9SUVOOCWQOc5oE8g2lIkQPFl75fcQsfYB824f4Vr2Dpus7b6xfZcdoo2P3RF
wrTXTPU3Vwh4ZrsC7H0VcnXJYyZVSa2KjUUcuMmYRIbwZn2Vi8fGb2c7Hm37yx/i
IvXEMbUbYhRzrf9wpDEBbswB1EAoJEzOqqcsRIdC+JSVYMFTlaHsvElp5hjntNw/
iW147qLeZg7/OooZM4zeyYs1iBd/y7dQiNgkdMR9n6b6mIqZPjaiIjzJ8T6DLFyK
EfpP4AEeh16ngD7iKaDb5qe+OrssM3ZRLh4JajoodKdFotKHcxqyVroLz2YrF216
YlyVCwXNi4XIZPD7v1u/Gxv1LY9y/ODa5VW182DLUvILOrSTMpoeXIS71N265GGv
uIAYwEa/a6I8uT15uYKDCgf/phpfOop3BFgYl+V1vHf5D0r0UoEUctdLy9k+BpIA
4mlTARiShsZo/d2kFPGqAofXbGQ/bQpLPTYwHGYwnX+NSQa/ZuHha26LD7SAcp5d
B8Dja0PbhJc2YIbhAuEmI2onmiD7k1BAp1NPpMUD1B2BTTGNUwOVXF965fLEeTy+
mIOHDz/5xli9bRDWBwKluMkxzBeZA4qRezJ8z/QQESYcI7kj2AJxJI24i4NbWvne
y4H7HuLEasROz/LnirTy/6A0LoeaDih7uSTluQ5WLTWETRc8TUscbqsyA1EZQ16Q
TH85EHDpkYWKXS1sOLWnfQFpT0IEBTbk1I09+ZIx9nD2evlFsSOmsWeriaWZYTWD
okcpJlMBv8V6BAz3SVpqwAj/bVVFmSvtbVn3hJl9OB3ZG4cPaUcRfna8RxToJoKW
s4UO+DVaYBgdFpkYd3hGMyp+e3VJU1PiXnisgoRdYh/nsj/2hW+VGpZoF2+PSV6X
hiCK1qO5846iu4w2/SgukZ85wOZ3K6LXzv04RIYmae0Zp4FLBgRwyBuNUqDFJDFe
aqFyUgT9gf+GZVO9UxPkvQrf/3gM8iqXEecT1imQvf3wgDs+oGmAh8wUKaQiLb53
gacd5GOxq09imlzldDFNjX7LXgM1NNZ3cTRAxrBb6pEIB5jIGk3UOnHD99JFg9hj
4CzOeq2KcJl3jqThBnGAWt5vsSanMidTFkFI7o6211Uppk0TpiYRBuRMDQ91+YG1
qys/MbF8fuuQZ6gcf+aCW3HYV/ilebjPPUlIhqiwtd6dYE7p215YSVzeoQT0tx2S
/jn0OlJzTRtOd3TDRT6ka0a5acQAMBUZUaEkhLlKXgV1o68RE9YAAFJREWcFASJY
1o3vGVihUxcEh2fJeXv39LLQkVFuIyk90pVb5A+/6hcg+uGtF/FLxssLc9hOBGZH
K78MwRCewUVXg1zlsTH7Erl7Vx9jQgHoDVX+juUyLnO9WMw8djGEXWab7mtmIimD
sVz0ZJy2M/7xwANJ1HIhAoiLveHBsS5aFktWxosElQaGXjOWtUUyepCoGh+OQSWD
PNSTCFTZJgBBeCpTPGgcvW+7MebSgrsxeBHYEU3QfsaFuxBl65mJLmXeZl2apxXA
g0XsdULGlVwvZbeDG2C1H+cXWMXEsHBX6rlBOTN6EICOHdyMZEOt/4XWlbCBslQB
Qs58eMOGgK9Z0XAbJZKJFQ8cH1NXKStt6/NWfcixs3VqWECULazORdAN9RF1J0e5
G3SR7kBae0crzCllOXQh+aJUFCIsq9BlJlfer3miEtVg71wlLWvdZCfPoA2ipfYW
OX4Pe4SC0XwaECNzWjkWfC2OWYegn7IJanZ0MjYJpSjx9D7Jh1E4U5PbLxH6hy1a
adgeIUb8m9BkbYk32T0Ic+6/UU5K/D4n/oPXz056FYiQ/Ko+Zmkc2jqZ/GbNcbB4
aDTGPSJXAG34ua0UVkN3P+XBKUSR8CtWZIP9Cz3saEuTcyyT45lpoP02P00AotVI
IYRZA8OXZP37NfuC5KSySZ3kAc7+NWAVOEVsgy1M70M4MCtCUd0afBa7fOQRMNeL
0zRnBTQukPvPBUVOQu+2OEd0xvsjruvtHpRrs0EelIWjAAz7PMTNX1erwQOxcoDl
8rZ42OF3HXa9yvGLE9Gon5VxKb0lUT6oOUJAlh5e+FY5zXL9JT9Nato44ZdZZdoP
qb/W3KX2asolhxChOxKIthynlDo93J52GP340AVNJBFY4l3QrGkd38XBwRufBmfS
LnXda5HpSy0/vn4LSvNjWeAhW44KDC3LdOuwInXuyCB71Wghdnhahtju7S+ckJND
7831mRuu1CAjwHXmF/5aGLe619xEsjeOD7niXYu/cQYpuVYiOyrI3NAp4fxfkX/E
by+LrzZRQg7IraH3pgkMMG9MjCRzbv4YYmLSioasopDOE2bNWtVvhMy0eujxHwoK
1vuPHrjfP7zCzGpFzW9gg0rSHAzPWkZBx3SHljWxb4cUlucdd35RPpb55V6ByshX
YQB7u/ShfLQuiWzMZp7xcrzuKqD5IA6anUaMfZ0ZIqZ+7tpm1vB1UQ7bE/kCKzsL
u/7jHX8wYobxa8sWaOE96liJPFFVL7c7FEk4Am6ZRpEqvR0WNl+UXRVb1M16umQB
tMPwxA2ekpWeuQGrxVnfCcuunv6gjQPgYXsIDhGzju0scQEIgVt1Ul3UK4NUt3dr
//h1NwfClCTAQsM2KnsZrOUgYyZivewLASix9clxtNG8SSDvCsbewSxo8JnFS+bL
ZzeOrWNhDwO1ITVQxhCMwob/wXwOrfcr+0hIZrjEQ117oTJtikwuWppGqaa8CN1P
rJk3ZinIwMD/Xn5nnFtpNxAMx+cO/mas69tHpPfvLJyij+xam7RjgvBlPlhr6QIt
ejb05CfluWe1F4MG7rkSsEBU2gdR3hBqb9A4yGiECAnC78/EB6NgUOKYeg840IK0
wlnkiQho58ppi/hWrQJ8pbQwRrZBAofa5GyqYOGBLzBs1opp05IDX42xQtNECQg2
RdJ0y8I/2RIGDOy8zALt/qoh/NtVdT1PGpS7PwMIVOuZnaJq+K92+aPttlLn46Cx
PlcvFwIM7AdkXnwPEDH/BtobrDaE8F6dEzypgn95oR6P3Mu0IlnWKAOiQGiBOYbI
nD2Jiv++p7X57cMHzwvK9HQzcl43oziWXuiPAnz1ERxLayZFoc3Q0iNDn9v6yyiX
MKmVkwlx26apV48w9TXq1IdFieNjFlSUPYDEyE2lHFfV+A506p/zrrwxXrnioZcv
i2S23Z6r0PzXBr1eDt9xKCyAPhw7Dzno/frgGuSagYmvmYOPPXeTI+2IZbauJ8Vo
sqSdIpBzTg3vuzefTq6cnfuOrdzuY808I++hUKkVa36NLVAzkth2HRchkBspLd+2
p009U2HxnqCGbqdtg23HU3cuGx+pJC8PkOVKo4U/WliFGmGu0sqeESN6feNWISJt
Bfj4g44N0I26QWwFP8yif4eA3Tb1wfNkMT/wZ6LTn3CfTik3SWDv5H9DPcLZKK4/
dubHpGh8ajVACFZqorlEuE4UWuEq3KhCQzQLTVqw8EjhuXt1mZGh6t9xYRqYkrgR
Uzb0o1cKAS+yjsaqjOcqkbbt5G+P1aGRBKaljCHGOtA4QFMPg8YyBbApZK4CfFis
govLt6muZ5nVhgvFIkc4hoRnx2JYbMKvX7ArcKEP9wOVOH3e6eNZsojGudZ+Z836
NKKivoQKgB+vDyEPeN4B6s76oe9xo9Gp4F6z+aUH49XMwmtK1wpuGKZXwXUbzKFL
aYLztfP3fqj5TmAUcMhAsD2OSSwegXmhhi6SY/5XSEvmiSaw/Jz5hAvTC/7e1tch
EonAlczOsBqn1dCupogKlMAJCseu+bkfGG0QdBaRBRz/xF1L0EMELF/cbHq8KD+k
7+SE1BZZd6+b2NdM2STKJ10DHkzbgbDlBxIPHXqGHUv/DPwp24t+fTqqKFFtplKk
Y8wFLboFmJYgWkQwfxc6A2SsUBAsKdRJvxak183WCilEgnjDxq9wcFiMcnoxgyBa
7cDIK7D9gIsE+F34apRF5wEPWaGodYHuRWAtNbY6j0SQ9w8R2xX9lbCoRRTX2TsR
tZJcE/idqOLXG5V4YM+vgsGLVxSaQWD2+BeBajb0i30vCaFDCvxXsPABwJgCb4Ct
sWloMrU1R74G7fQnywRWQoXSXJTR96EyH1HW4F1ioedaIMxRTeZEwZ78u5+ZSYSr
WVggVYlsbhxwpJkjFlRiCpSobWy2kmgd09JTj9YIcOn3Iw8BpaFkuUyxwuC+wD9k
0jEEIh2NnrFdR1moFws8RbMDUWtMOJtirfpyj3xbuZDVD3BhCwxEx3mXlq8RqLdF
+fFcXNgAY3O2AKWC9YZ3HE2LUmHkKwZDuy43736P+6QpzCxQD4GtlOP7n3pq5aYq
wqTW4qxh0Zyym9MNkM36Zj/fHXgRehUQigVZpZIt3HJHUEYbN5SBqLi2Oc8xfYUw
FttoKk0ACMjQid5GUv5JQ+gF4VTN1pqyuZTVb7ei+vbCFqGt67b58hGSIfacNCpY
kW9x/pDUNdyinX9fWaoITsP43gZggNgkebMlDwowNtaVDwhVjkWE5VkGhbB0psuM
Xt/Yb9WLkYnmFBQhnlfC7w==
//pragma protect end_data_block
//pragma protect digest_block
mr63HFtspOO+/wgi4CrzpTYOwLQ=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
imtwEq+W4jDdvprZ+c+hxHTGILiVsxxaVHYPHJDt/l8s1M2G+xDtUJr6EZoddYic
UT+hk61VY9wzFA3x1eYYMCSXmisGljPpiIDXlkC8UfOxb3rEosPeOxmxXS7uQoyD
sE5DbQ12wXlNPWUkQ4QBoxTInCBFfPwH/pUcs7leybZqbCwpKW4u6A==
//pragma protect end_key_block
//pragma protect digest_block
DJD2zw3Q3Rer7NWic4r765KcEYA=
//pragma protect end_digest_block
//pragma protect data_block
FSGgktSf859poIs9iJRBf5hcDeXcd5EZ3MeKg/IM+WlvVeynNl5+bvxa3uwf0MP6
lpcWmQQIxy91lpqkqwhGcqOm4K9aW33NDxL969QQI/mw1Fer2fpQ/ZHyJZIZs5C2
pgGwjwlBnPhsS8GPrMyDAriHLhDziNmg+0XtvEZ7Jut+T5isBMBgJDitc2N+F6C9
S5wJyUW8XIOlT0FlqWIHNKZ3XoOzeqeWoirtH/r25bFJhiobTChIT0WhXFuqYHwE
sb2b5WMPuLNdGNvWpqfTandzbgXN9H+DzzYP3WyJUDTnlgePj6GSBIV9m64klIk7
g7knAicr5tsU053nzS3PJLFjofMmXWp4so+PbWotjs5DtXJXXZ38nCi8E/9qrGB7
BCTnTO5bYbN717y1+y9C3zgCyCuspgVQy5yQrmqnMzz3rw49Gt736V/J9iSRQMlv
tNYAUjHoJeRcVMj3z5Gtwp2e6Ejl2MmkcbMqG3i7sz/WFDVpswy+V9KtMueYy7Qf
OkPA/HgL1m+zIUrm8Py8dlfw5sXkQprvbh+h0dN09yNndVIj7I1revWbrfgbU93j
BMTpPW//58hyBRfC0uwnbLyFQIyV/3rmWq/vMGNbNSRbZPHBfHh5WGpXfxltK7NG
erbcBSTDMOK1j6Cw/AJWXVnNzndtXwPBEVpK0mCRjoQ3y+psseqLLNLT5wI4ecHE
G7PPwXycmONfniMoVqW7Kyw+cP+0fDHnlqpGQRMWrt6J3dzfz17vcDWTS29luqIy
PNxPY9LaBlH5u1m8k8n+lVexW5jw1iBLw5/1nG0GdxkJNtIuZu2T2e7/Kavqblap
HJE71cSvlxvJQvweoMwUbX/AKL/kS6yftfG9WJu5Xz24iCuXox/neCaDPOhXEqOb
xPvhUYTDTswIuaSR3pMxPBC8F+2LILU84xoPxBkuFw3dBYb4OSUpVHBjsrep3r1S
LBMqxNu965n2ciopdrQnfWyuLcSDBwF5jl7OfvpOwCPhGhjlL1aPKpQXD7nNFnyb
ZKoMZrSLyPYIxcakoLljWDSNVWy3olAffsT0SxQbbMcyBP0XcIPKzu4p7Me0pgCj
qATc+exwp9+ffGWKIy5tu8UNaM3RQorIhmZfGPn4LMzG0MB45OXSg3F4OcWnGUQp
JM6R0DEzvhMrER8jzar1DPlND+SNsfU/7uc99DTSUXGWswxeQu2Tv7A7e0navG67
StONy1/oOGYeX46JlQIpYCICVp92qvY8z8UWe1Fwa4Fs2imOW7zPMjutIWjkIK0F
SSouh0jIRNiVr9Xt3sIYHUGBzTeB1lhSzLPJdga08+8bog1ashSFHCzH26nvZlLO
B0JCpqUEMhNuUL8V0Bq6GFd8UWqoM2QgBHgsJSTCZ4FTVWaN2SbtS81txSIPx6i4
h9fPQ1Jz76mMcj85h7zM4uFafRGeUh1uSv7Ft7NMDm3RXlbtvBLsrGKlk6CwkdIq
bDFK/h4MXkCi2aKJd69TYGj1SBSJlKebo2WzsC2KABMgpw5Qteuz36Hp7wyxtADE
qBVjb7s7FNQ4PKSaBRKMKlsfsi7OYqMDZmt0er7G/fWNh9lABDjufgmk03nHgqJ7
c0igIASBl2r0Sxe36Al6DwljQihYTIT95iFPeoOrr7Yf0kc8VoKClD0fBQQcAcVV
9TlMUnV5Oj6Nq4SUVcBCz1ARj9Tv612+3U5hVzqaAecnufQxm5aeGoArwr1Iao5C
D5NSBhWHGgVpH36Moidw+rjN4ipIwCC1yi6V95Rb83evy/jXHSzto//Dr+4FL9+1
xb3KORyRMCp7oWyz4FJ4wf9XuCB8QKs5BdZk8DUFZy/MvEo1Qu51pqApDxKPCZec
WLW8EGfNLvCPrGVzO894rwqttyw9/RcptQHNOUyvB2vWPR5PvjBlF7Cl3f5XpDAf
9KhtLowVQLRfypu0yLsx5bnQqbqpUE/NF530kdjir8NNHS0XTBVu04V24d1XBhTQ
dNlBsPWpJTQTVnG0IG7Rd+yXayYQhpTs2bfqTOxDScrs+WN+THT2Y7/1dbWsTEMA
vZakFuMp2nWct7+/Q3Y0yYY6KTzaNJU9btxEzfc/halZ2I7d5ezQJ/bMu8AYXE3a
LGy2vEse+CVq+2gbeYOF8LotV7DehHm3Kqkav5rcMa4eqEJaGhUaQoCeqJtbNiim
plB3ANLSkjgdngxWCNp6nTMSWKXZeg8uMkszqva5VrOv6+FP5+opfUzdht2+bo93
zP97He0zRSlXGTX5xf2DLOJ8LhN5HEXPa3xXV4eflBzbuHYQ3EgsRHyn5gNjoAx/
R817xmDWHJDZFZDhXW3EMX4ob4rJlxmY/E/lhmdVTobatQw20sJ+Fj6bncsXZF+F
c9JSyIIVpm61ZcUqRX7luWstHd98u29UZPVUkZWpYnI=
//pragma protect end_data_block
//pragma protect digest_block
6O5PkiTjbJQpV7hrHCYviDXI9oo=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
VzNhEKDGff1sDOL7HcMXLcHjOV+6daNFSY0YLrbnXmRdjb17YyAxKB1r/9wL20p2
4tTsEXmeKnbXBJxNAXiwBumOvUBXN29jLRwaZ8jXqoQ1jvcxvGQZtAhpFk7iFS2C
XgDZS/+7FqLlPUSjgzvCJYfHcjMWYH7w1LRi7EGEtOC+DkP+1CU1cA==
//pragma protect end_key_block
//pragma protect digest_block
J+6SaLxM14O9OaamL3pTPbilGww=
//pragma protect end_digest_block
//pragma protect data_block
n91W+nZlJd21KQr4x030AjpC/MkfrCFsW/EZmTBpliX6n4D5WCZ8x2vVfkZ3MdlF
aC/JIMr/OFlid/p+ktqQU4o6JO3NI+y0GmACu/x+KYfkapCJCGdNpoWfaOplJZY7
dEHiSIiK8uFdIobZiqgIo3cwUtoLFmnN7Rkv/mkNGfKSNjkIw2QGnImP07FWvhyI
QXBkpJcmOOkw2zMe+fA1pQWoX8FyOzSqDtKVavnKA8pnPIsHs1EeD95PJoh11vg5
W6LesAJDe+E+tPvxQh71fz+Fpx71njmaHzEYAw/WdtA9aBwLgbS0D1WFC5/AmZ52
nN+65AaPtTMG5khZPETbHa5Kx2VI45pNNn7oXPKdf4mjq6KN/Wjz9npAwmBja5py
s5Xte9VyG/5Cf9sSL9VWQ3fHj5Q9QpHWklSwoSzIVeCx+09gfGM6DPr472/fOPxJ
V5h9K2TloQEnA7en756N56ALxuDnxsQEkkrcDrlXEuSfJlnor18KSTMq++IMaVP2
9OdRSS2MZJKaeXI/fjJ6bu8gIgoTuzatPWdbONUpWoYP8Qx3m3Tvp5vDl79J9cIa
fMq6gUTz4FVxxLo/6/xbT//EwXrZDjXbuoK/wxdHsc5FpSJzsS6jwf9UlWSCQ/jP
I0x1tRMDFPEL5s3HoSL0Dyq6EW06Qn3Qg4Ik6cQpgMMi+8DHNzRX+rZlK4v6mWZp
sq+msKq+NojtzuyMptaPbtFcm227MCqJWwnd455N+grz47N9wnlV2zYrd7D4KFtG
B2K1+0KH34sWbTAYuGaTJou/qIG+jz/IBG9P6Bct7cBXGcGmwl1BSWOtVniObip0
gtbYtibNe263C3NeLfaDffaD9ChQQoip4RikooZnJ2RA9M3ko8goiAn3iaR4+LbI
K/pS+lsrxCZq1SZfkXAMWXLsM9wOe/SoJAIXX7/OC7U=
//pragma protect end_data_block
//pragma protect digest_block
WXunvoGp+6movjHqGhTQ+8mhDYw=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/jgj2HfOPunDlrB2IzfW8elV7OtIsfHwOxzWlbs2PLm0UhDjgOgi47PtisArf3iW
qIko+hxQvCoOWv6qxC6qWXM0GExc6XWPUK5qeUBHmzXaYIeRlR/Fg3pMOtv57cFE
r+xOeJp0SpSIjfG0hD3EnDhMBlfg6m2uggZPKcKYI2lB9uO4J1s8CA==
//pragma protect end_key_block
//pragma protect digest_block
s5Q8k5SWHqKwTRRTB14qBN/4tkU=
//pragma protect end_digest_block
//pragma protect data_block
+CnlgQVx5EyUrO8sVxMsiuOkLCOe0ZPZM49Pc5vFTURmnbWfmhrqeV8xVq8RpYW+
Jp0L26HKfVxCPM/RnvawoWCFcXr3Ahzxrkw68Yvc3asdLYXysD+3NTm6M2abWISa
1aBKHrFQ6tWSlDqgTxkRDK7F4KFXYB3j+yDelleD2jXOmZBbTm5YtJERGqi/qhRu
7zc0t6KMThqQtt0Vme9fzwel2woWFRGLy7xZms3CHuLoJitbH1eQZBVfYmrnSods
xNCqQPGfb9Phvj6aVifA2Km9KpO9KcSoT6U4vR0dhaHjXCCwYLYrF6Oew5/QT80e
GchhT9C+NxDt9+C/cDz/uPEi+MvTOMHuUyn9cA/H0SLaNFNtOONjoSIq/BKSGsxS
Nim7CINRdd50At/JTP2NE0CZ8GLiwCmViEy1Y4QlapiQFAGUZEn05IRp9d5lQGdc
bsLW+drRZQIF9/NzS7PzZGRfpEyFSPlsjUS76LqskaH3Wp6pgDfLFZb6nOhcoWUc
HGTJSBuakAQX/rO2eRJ3vqxg5H5vxOMwU0CylASTUzScS0B84iHxMlvN0hSyVEpD
PUWjjwgsh6gEj+EQvscJwYsZEbFvTm8l9Mlg8H/JseWiWKXrN4QGRZdZ+SSTcEpc
FXfPCUVbSWlAm8BTPEn953Rby8g2q8k8AIXOao2ZQX41t2IdKnHX2JMRybxNee4Q
m20btbHZx4LMs1q3kTFJWeXKJssjFNjLWXHqdPyeVYeeEGGY+MgoldZwKPlwPiA/
X2WUsfkFD1cNVebMv7QOV8kpZeFUctpJjnf7LLkxoUz57rlLPLW1XfxhcyujX2j1
wnXQzN8M8Y2oAgbZfDNmEXhFaQ2gid6tbvchLhAVmUxZvVitO0Xys1QOLfH3ZM3A
BriJt0OgJNtV8v9ub3fpKRITCQ2cIUlN9L5ksPRh+UcoV4OpH6wSLXVFqPusIMkP
qc+LX7pqTxE9u4VOKTaJdGALAuTInpWWcgDtK0v1znjKQIIGtWUSUIlY68SNJNM8
hrI7I7unGY/FwLnJjIJNtAh7nErbocTp/jxe6CzdZ5QwDfG/MEdnDQdILIHA1hkA
xXW4qQL4poEXwTEMi+YWIC/tW27xmy/3n1515OtSvOkI3vB3Qa5tiQjocGFf7B3y
3El8+iawof7HwLmA0oILfM86buKtltmTuGMK856eFGhXiDRDVFlivNxfu+ty5nir
Jw0zbBtQfUqDKM9ugiS62Z4aUzetotHo9AkQWS9jJ65rKjvX1C6G6YMNrVHvEtId
KN3/wX4Em3tlLBeyVhiSajrl1ftw7onQr+ys9/8cL6lccrZ2AFRherhy1yKr47b8
C6WhRxCpl/S1E745YP2AZyl4nWd561RpL4OwrwdD3eA9OcWybQmsuqjxbw2sRgIx
qdWptns8oWOGf0ekiQojxjNwWLb08Q+hDDdEH48zzL8i8FOmOeYRWhynHxvTcW58
pcTVDZrkz6SQCCxYe6b3h8mxMvLh8rNgmJINXkW1YWGeYL9yadrk12Pkcq2NRLAb
vBWIlkjK4phU5yuR3HAA3/lhQUv/LWTxPp6dT6FB5vW3A0I1BeX3Ci7+oBzmaWGm
P9boNUEXqzOJBmT0V9yfYBIjc1/0F+QCoBnKnShqUHtvSPH4mr+VT1I48PNQaqxr
L09jgRLqmTnQnm/eEzgjUZUhruI6KMXlvAU+hdainWSlDahW/LONRvKBc6qpY4Qu
b+YdhP3s43o6ej2M2ZfUCBJKyhaLowGXzfc3rRVzviJcvf80okG08bFuyiretObi
y10UuNIghDNGV0kXskKaIO8dxgJCA5U/smQFKDhm9OM6x8zuPB9VHgbQYtmo0bG6
s/NQOEi/DJ5npuJUoeI9g6QFI0GehY7YgtiF4ZTMgbcUljGgEMNtRrGy6KHOlMUa
8fdVc78OpYAT7LluRaSRBSmKHxvNIirjA211+5WuOfF45Gc0b9ODrZplNR1i8nd/
iPlQ6Gw3EWigWRl0285pw2+xEoFY6nla6iAmCsoJ05B15sfuSPPPsZz2tT8uubaY
sKeBIAo7s2RXetAHqO7/sXgukM7bG0BFZ8o/jr/wQWBkwJtYi0qrooOyto8x8QEY
lufzUhtqzhcwKH2oSiQ9PUFB9mhhMZ28eJdJxdyNPW0eLI01sy1ZLTEO3ymNaYSG
oFJOIx3AIixVajytpRdxcYFZvO+4Tgblj8ECP2fn9F1FahmbkjaU/ruEgat5OfCT
Nv1oBJJSroC7D4CJt3pq5YnEtkcg/r7A1eTCnwLR2hg/xn0liZ4QGwE6sLlwT5LR
N4VWnKQBcu5MAnAg3t6lSESXGcdikoI3VBtoziJJX5W2fAHeKXvuWzlXtC6nHqKv
DRPce4AlCGN9Ekil/i6Lvsw4bbd+Zud9DrYzL9zYDbjF9dq0UGgIeInkyg9cLxUo
SPZWS9T6Iyz5Qjv2gRGdbJgq58cP1Iil0Dcc0RgKHRakOwBWEXE60cb6w1a1ZOuQ
wWL3AcMToyMAFe4rRNbHM0Wuhv4FyW6nGXZwSLrY3aBtigMcNBim9aOaJ09rqtpF
fJaAp28Nis+I7ecKmql0Pd8fhdA2/FlitK2txCW5Rf6zhIwx9SRXb3Hjx9Wp87yN
v1FZhXprphdv/GHlqbraOz8KZdBFmp/KjpfvSyixJtW5+eIDJlHsQQAvgqm8AJw+
r1VfWSOPaUJnptClac+SN/1kGVZTyVUSyBvprDpPDUrWpVD39YW4cI+maVw8Gh4n
BOaDntCQMhokohPad2yLi/CsLoFXsn8VkbG+7JoNrM4pxxMN9sWz12zllLhU2/bL
wtOwVRQ1qM1ZHLEVKKZ2e7S5xlHaRUaY4Ex1QOpzc7tWVT0D2M2bbJekbYNsnc2C
9CRrLJ3tGlxQ15ea+Or3kCOk8sYOs/mPOt8vXhUBGaBJajDaEIS5gBDxBQCflWC4
NPhrc7FRWQmqITJs8rM8qn70iywJyYJ+wTgX/1jiNRz63kft0YSO60ciLE6z8cTO
Zq6WsIVyMpYlZgjkmhmobTrHxrnkgsI1klIQje68WcMb/hJWc5rj83Yeg8fqmnXJ
lATS7Yco1AiO7DpsEZ+qYo9DypSyCuQnCXHJNaQLETnYe8AfoUAxvSra47xkRteV
PZj7eECfSL7pBfcw0ed0tJvTdOQpURjxs2Y3yN2vKbRxdREmtuR9EG4OcuVNER1d
rcpwsUijWSp4Quoqs78NTIXWvQiJsDjheR3zp5AG5E69HN8smWqbUBXINcSht8sT
e+Qh1cTVC1zbCZWODuc4gLlf5VooZISoVq/OY5XgdmSyqGzyapjBh0uZ6vjBRA6N
iAsPyITn2V07WSbugOfsOY7rCUKjSVC0iWQD//3SSSGfn9S9+5FWFbaxOV9NADov
Zm8pD8CngMW31xnEILfBOlkFHqbr3OJRkOA2N3cykxZ5v7tyofeTu6R2IOtz5mo7
3QsFjHsn77mHbpvY37giRM3p6SvHHUodyxgsWjkxHtDlc8lF3hDDvf/dr0C+QIeL
X7jxlIiqLntom5IhnQDF3UKvIAcbOiLYoZvBasaJgYUaGJ7wDSMewkYgTaSuPVKC
z1p5TA/fYYhkoAHmSXR84gomfUxKB0GFMUlUCkJ00zges+HFX19vJCE+XjRe/8Bl
7QuqiS+qtA6DuYAnfk3pHBqvgqZGWwvOqTARvi0KphK7Swgqjvfl+lOx+wgN1q5O
GiuXym8qxUdIU/b1krzGrRGC0omz71le4AfnVnihmUrOjT4mIm3w/teD8GmSvSge
ZQxtbUOo9quQD9VlO6Xn5zWuATN/mFAM6o0I5S8c3Bn1dnB805QjxVMvpvWac7nJ
GzTPUyyJG93n6UaGMQK7IjoKcJoG/7xcrfhL4LIR03ZgmN+4nPS6BGu7pgM7tUcn
ufz3Ulftl6soloC0GLcnhImgwbVvdaOB22lpKXapcL+SFi2r6AoBVgPRdsn73S1h
wvT+fkXmkv95EZH3Wh3mDk2l//gASHhBTAYXnCAHfVOG/5R1Rs3mlp0gdoQZ2bJB
9gcm3DcwFZRGHF839WKmRafuKpDNTwj5Vxd/x9v2Wyd7UCPH6R4CL0Qbp5rxmsnz
uuhWqGnYb65l/6VeNycRdg2Fm10iz/Y1OLwzEM0gT/GiHVNmqSBO7GJZ1FZxoEou
4gzw7RLgu/F4jDHSim1rXRu4kQL272Hwx0xiYt9u0tgUIEBAqzCTLWjLQfR37RL6
2FqZLbA6POxjIMxVDb/Ol2Mn7w0K1N28E92WF2P2isJ5iT+eTmVhOatrwBKYgaCX
dLS6eFeR9a/mGwYkKVmqEeLEWfjZhR2Poba+NTXAZRqboApzVo2nAEA2wXR0zcMg
rw0+HKFLV5l8Le3S2qtEOCDbbXyW3SsvQ/5rOHbzc2L2xDcHx5x5TPY241dXaB0T
LhlAHTJgmA+OWWmxWBrJOjulqaeKfGbTL8ffs85NyXRZk6UjkmBJVUknAXl2G/8Q
t9uc7uayYxNPYq8X1fnF8yvOaVwO/hDziGwfVQ3GjyCPiuyyyXeWyqQpZgcfOaFy
45eBj4QbPgtyaC3khh7VKKBxK74j/He8Du9Y2w+Hw7IVaVY8+Y3Bivf3Tqi/WvBj
PWfRw0IW0qTfulx1E2HeiIRKlPNCL1IeUanlNm2O/JZ3AmnS+DSd3cPBeNQevZbJ
K1mhOLwsbHI/Mj1wOqxym8d4Hz0X4XXFogkrgcmtuXZq56p89KQQ9jJqSSIVqpE8
mG+VwK4bigJFuOOwLphGg1v03WDBQSwnhbbsWyrmSt3bxPvmpVsNo/Ynt7cqGFAU
zthCs3z5hMzbpjyOkDgrf4G4r7luU6PeLR/SNCDRPsiKPtZVfJIb2E4EMQCfbdhC
Wyh9eAyxPskBPOiZShF00JEjoWuFRbPDEDjzD47zKPSGgfAcp9SIs4VlMeaDMo+L
UOIGs2VH5fL3I3mKzmdCDa198FO+6Gc5+vA+MyUugE/PVDORlugCbJb5tU84rS5E
Z2N+ZCoa8VSSP79bv7QkbR/lQZC4I+EmMnZTW4xNnqDyM40FK3fyzOWdrDZPQM3b
kFpkw/I339gmKnJxjdq5Zsy57aTzc1uJq07B3e5P0CvSHc+6KLz8VzK4wVdP6zkF
XAvixK8IkqMUOogJvR9knj2Ltaiad/e2uE1ZcznNQm8WyIcH0kmmLPJVRmJ0k8GJ
s7J8BtYSzlFwOf6TurlwNsipyOFcz2M086Iccnp83kyJfXz5EmfNXzdv6qlLVt+1
jZKejWWBjZtLvD9HYIv0TibNUIGTOUBl3+trTF9r6ZqhiQhVlzhmfu4HrNgipW6f
bddQsZk5XSnE3YDlEdtlyo+34/HIJdUu25838Cp2haywo7go0DE9YiMt92nmxSen
lWploSnBfV9GoKUJKdob8glaTGaLLLfP2NpxffegRBIg7Y9ZME7hosQk8XWQ0WSc
82UyVUZeGK0e4e8IpnrEuoneLNlX5PoVuRJndWD8FAHgl1Q2MJmEpiPX4HXJxXOd
lnYYM2pmTvRETNL8OJDsD95qSQQqkKaFPYzXidswIbUak3GGFTz8rq2peKm+aDzG
R6aJZqQiv+Jqypfb+hA7mXxkGoEQVSV1LOrIJfTIiIc1JPg3BQijAnx8oCDMfnsD
rfgm+ld+5HHJJJmzsRZhcNu/d9U9BNDhcftQb8d0fcGl9zw0ynKT/nFOr/YFrst2
Pva5iu2aNkm2db7wpl4WIUxvgZ8A8T6sE7kfVlbNgIDrVuJF1HBpXuJSMiWL79Gp
FsNedU9/PKJgGNpytkUk/l3QL2zbVxMuOFOo0xGMeVz6ojjNKQ0PTvOudJVitnUh
/bts1KtUkQUwmhBOKZi3L7PI9rvCq/x1w2H9AT9TWceClmxg66Ya0GKOsECslS7q
SsABHn1xKTAXQx1x5fIr1R6M8FHM/SRE4+AkwbFLWfkv3XicrmF5a/zeg2yRGbaG
sNX71cLHHPdVzOUpL/4Lg/8ZLvqrXnoAUknjiQqaRDSA7Fmdvazd9SH1vLD0PR1L
MGQxuwVAtWDYXkLsXRoccpZhMSEFJkBNfDvZAmCLX+KFaLC5ruW5EC0Dd3MQy1Pv
q6pcC73JyxyVE0zxpyEiAjLacHm2NaqC4+D8e8UzfaQFlflisOGV3n5/eBtB2AQZ
kwG6yirSXj3UNTxneur2Vuk9T8BGBGqvhtiISU+AQz4sGXArKHNLbkNXc2Uc5iQ3
I94wwnhsklwaW2sYhjWt7gDXZgN5s6heBC8sHj83TSLohnw2v5Z7kHqDAyojtgM1
PpZceB4gN7coLkrtjPfKbClXbP2Sbau/wYr2B64l/vzHDQqv7IRYm8XxbRzmyy8V
GdlCjLg5ZkqP7HllcYSqTbF5RY8kxnaxAV1FLgNIXwrIcp5thWP3fukCSLzL5Zsl
cVXwG52nhwrpRihoymSeqsOd2UAbRzoBtrXBWvfBmPoiXbL9jmoDgB7jD4eRlHwq
p6nPzu0HZoYTXd03tsKov/6FA3ZrghwGMMIWX0kSZLo6Watq0CqD+DMwtievypRq
hfSsx7bEddtRAUpqp+u/y2aEs9xzZzlDpn6zcjGDTta0qPC1L8HJwkV2a8fKDxm5
7HDZ79MRXCY2zVKScN9Nshyvw6Dj3LsQA3qXtahSVCUv79xy7CAr12Q9IwULCnfl
fLzukkewDh3YeFjOGhTBC2VEpPbD3tfiAA0QN90S3BLHpZER5d2efCtdn7jlhffg
AyF9HUDZhAcFPD7mIOZi7tqVJQtY1gTdFGjqxP5w/9Ljhp+1LK8uOI5ucii9WjY/
k/GzmHBLvz9OppeqcSOjjm0jSDHmNLcq1FqKKGoB6ydEBoWoZ1iIEOPM5OxIkjzf
DPbCgWQorwH2jqStPxRj272WuSI8/Omj81EG5gGMhVsoZsvGyt9rc6xbFtr99x+o
24LFQyDIt636OmcVFSGd5iy2M23lG5WSmhCVWtLBiJFNRY/uzqTta9dHP57ughNH
55OHBZDaoWn2JiBWibjUgKqDiAWVsXGE8PRt5yMZCtXKTXocQ+26rAdagf0j+4Fl
CdlwbIJNw13CjhWAXFYMTSVPnwTivqXYzfdFqyMuZSUEJtT3crrPoknXxgh+jQ4p
WlNOQNpkp/6FG8Kfmqxu5L5KWM81Whh7QqpQeQII/1HPtvVhitIhIZ9FCLuG1GWH
rARlfwoOGcmad1a1OPAvOuHfLjifIipju7eQwq3QXzlyGai7tcP8xrHezy+Y5BsZ
a7XIThzYgSFmrdu9EeujbyaQhCG7HV53pI0piavKwMPzUh39B8uBEw81PYvnmWSJ
3m5gTiWDx+P/XxRP6xgYMMV4onS1iHhcfqfNb/BJ5Jt/yecbOIX+Ke/SYzde7L9D
OcoGNMDWGzyxOqxRC+h3fJ46BckASCop8SlhGd4mZSxvJbOtrtaH69MGHyqfZd56
UnsU+/LgJtH95Q5NRIxMP8DLUPpEHi3fUzmZgh8NbRbfglgUU2GAPTRiTLb6UC/v
A0ABddnkoP5OWpe7dYQrUuTynTf8bShiceEMYITYLgijb8cf9xTQMGa6PZ3LJHu/
A7YC1ssJXR1VVBMO+QZ4tpWuaUeEcBmWdM9Y8LDYheiPDEKyfAdyddjH2M28vhX7
//ZlIdBGJvUAUA0v+LUw7D2aH0SCLtURyzY6y1zwybils+QwCHM96sU/8pnFEs0H
MTr956VmvEWoHPYEuxBctX1eia5uiZ4wirQbzN0G9djfdr7YHy+FkGccxVZ096vv
Xn1mua2mvUmz0Tr4nA1Egssf6Jpp3kyy0vEEHm3931+C+vryIILUGHrOCfEWEsPk
ZTRZTP53tWbVzIKBkyWkSxLG4mK8uwu87k5w3rnICNwous6ci7OG7DolKFg6gdh0
Xm2yaSgPhM8oakGt/xVbUv09jEsYArbm/YeU/NpJvCyUBx9ztZ/nphftIOh+vb+d
fiheoaaSMZyEf8bkUo3u3eCq4VfPYkBj41Quf8hAyajg03qzbjbPQoojKMmvvVty
rjXpFl+fKm+kDUUSRWBWl/KQRz1FhPGpruiFKAu4o/8H+oVUDcrZ9QYdG0Ot46Zb
CSEvuQOBQu59dcxiuU9CnzXGueSDcPnS2HsOoydeoNDD71md7rLwqny7fQm+RfkI
GGTr7xVlYt76LAD98hx2jaTKBtt0FY4lSWK8kc1qtSuYtSMJ/o6g9ibSL+y5rZZl
8vfSaQyLZoUKyVDPEJKo+F5Vxh19BntTdw6W5tTaIC1PryKgwC/2crhmbOJB6Tnq
edPkjq8CY5FOjtQxOPPtVN9FZOQkV/wcuv9B7XwK1AA79NvGU0WNNeaRmGUHCGDh
rgjXTy0gVgOVanSG4oXNC51jxgJBuka8VhOTj8v4Z0EBlyihcSj00a296+DVN6dv
gK4SqUtEpFiLZPOw314ZB7wgrL8lYjV2hbni5QfAzJmY56xzbAKUj1/4h3TBlIBt
+pTmS/a0ykHE+r3Pu0U5TUieVzk/Fk+UCVt8qW52CizY1EYi3wwSd60/oLh4C1Rz
lzTXmV0lNJeJ91/XML9j4vROTTM/VaCfDPzRnbJ3Leq3e7c5vZT5wMn5JwiuCH8o
yplZ++9bbk4QejSaXItlM4XHs7aDzKnQuzayGmXn/uuJfznlcSFJHkO+GX3bKWWC
mIgHEajXpBbxazrun0XSJPBZVH6aTxHY6XOqfSOctPw5cqKeYy4EU0j2CE95xfdP
EPhNchQ1I7XJwcbNECeHcEYOEM4C6PDHxYdj6o+9FpMc6kjFS5EKhw57ZjXm0a6O
m0kFnvqyUSDcr7SORPg5baQpk18AdjJkAZK5Krf3NIExLJqmRcVxYLBPyfS0VhFK
b1dPmtIh8VuVPSzHECV85yufOMiBhdgN8+XuoY6xWjGybgge7UedUxIYZEiTxcdM
kzyVsyVKDDrqY6J02mqmotCcWvbEc7kPIBKajykw0A4y9CtXy4J1oNec2m4Ul0no
31MTy1vf4SQUP/ZYlLJ7pa8GeBZ/H+kENtujROBthYXNwOd4P5mzBVrK/jpuA3u1
T4cZWgFMiuSpXOVvK/89M/FDQN+sY54BvTUgnyH5wD5scvzD4H13geKLUBMvz2u3
H+kyfbgXEt6a/NMg9aPZnl5mQOvXUrAVwaGjcXG82XQqeG//pefrQMoVcQzGXpjS
oGyf8HmC1fLpydo9aVd61Cy7T+JJkOh7PhDw1v5+Cu2+TKDhkCmK9UmM4H2bNDOb
fX+A+56GGzrHRScgIUbck5EFfQXE3Pv5vrFW9BxifTXVwtnlUlkF3LI3En/YeB6G
WvzgmO+iS2+tWVZDKGCIHRQn+6tmIfPjb1hG7jn2eKsz5CyiBXzzPV/OHvfLAFJH
qeZ0esH7jaxDHWqd7E44j3jPajQeKUx32TNuZch+RNN4wrfslw+6WmyjlL6RcXEs
tyqnSG7KusvxbqNk/OJssrViPQ7USIOnDeZ/Zv9VUuj8iq35M+YwEdA9iBP+wI6o
IJxDvTdlr0TN2NqeONRnrxkc7LWk8pmKxMLwDSjHyfDMcjITfr7FF68AMrezcECx
CxBW83HHgJDDdIiufJU+B5ejsoi/C/gpjo2K//IyJ+zQUtTb/+jtO3P7pZ1Fwkwa
LMyDoYbni/A0ecm83FrGa3ZSj5dGxHFoouC01xX344YKUiJyJNZNMp3tI/30L9wz
b6QlA/Il2p1+kMi7vMv6M9QopNvfIxVHKbauOSJqCbpMOPYgbZGOdPNLYxJsqCjb
7oO/5Sde56E3rt9WEZA/L4pTYihztmRIQuRoNgPNCkiuisJpRWphKQ5cHV0MipYl
SDIpnXfwknp14UlNeD5axWZECOzVOpWhgFv/LlupWM1l+q/OvHRqz5w5vLbV9qz9
UNJ5yv7lvez23tYKSPodGxgykQEz1/1PlwPj5zZl1nv/F7ZVEw25CC7h2UpVAlRz
TCMneR49rlG38OFU98t6XRWpZmQpNlJxeq1fz7oysIlsgJpadUOBHwQqnA6MbC7e
QdXv5UIOyk8wfepjpL+XnKgDhaa6S2HZcz2DBzxwxHfoB3PKjc4TIOGXYwX3zE+n
OKCoPH7ZwOOVCTqhBQHkjxFu4KZ49Xvz8QOqXy4oVni61HEyLN8QG4I3Ps3tyty1
Cvw4jsAWlY2/pSm+Dq4jrWFIb8iSfdkgnXpdexpyPTapBwe4LPu6Nix0uPaISmWb
TLUUsCS1F3gmSqrhIwbuBl9xIlwUdrZXSf7IrffQIjkHJ1XWsBMeJP/38NVsQgvY
XHIMDUv9MWPm+CHfG5C/fNDSXLeSHCDAjWbL/xV7MItdKc860YlXE0tiDOIe0SZo
EZmygVGLCipGEAuoDfcXD2xpJoTtO22ANDo4bov7WlpCK38QyeeTVmykOW9MJ15+
We5SvWlQF/FUhNAJ1/4/h1SRq44LIG2D/7hnQZ3+PghAc2gVc4StC/R7kQ8dYNG0
tX2Npj8CbRn6YCeXzpGUSO/5ML5bVng6SU6bXzOvhgjB21PN0no5VRnbNKRtG2MQ
jhUGCI25lJ0ngjrNHGCEw8+wS/hoKeu3vt3yBNXRZgy/K73hixHn2jX3c+ud0BLy
MrSi+tS57nS1i/mMSgPPnNTeFEitj5z0B+38j1bFvPzRyp9NAZ5rr57nak+Q2hgf
omYmhzQljK4wPUKkGpYvth7FEier42HvreKf/wIMzgqHxYU07YIWuvORgOjhOucI
6CYXqOi76JlJEyU2qM/mGZXKphwSnxj7+5uzjzOd+QAtePuKxmr3AQazEXCm+yYy
KFBfATfuxcT76dwCJJFYosJKvm+F0dJmQ0r8sJSkA9Uht8qfZwVTzUoNaL2NhIXX
9sriwT5Pr7+jUEGQ2SoDFh4v4x270RRk0DjRA7e+UYor3EHSzOpeu5mNacSY3FuO
tcHhh0pFkwjHIGJjJCKNkebAi9T8wwE0omjR5JYSUg9xezUaLkDP1M26wMvvvv8g
OnTo+0OVDLWmx5SSaJbpTzuTtBgqHOl3RXjwjz7bxEAb41W+a3c9h6oA/9OboJnR
AV9upOaCvcXomwB9NV956f+HEAiUMiJdCKtpxhiDXxCwzlZ+yAoq4HJVwVKETMaH
24WgTuqQBfzU/NN3Mr8XSyjOuoaB/pb0xo0AmF8Kj9ZLflv5gifExomIR4WABE+t
ZFDnCG3k8mG/IXu0iBPG/zpXw7sun9LKHPNoX9AYei7DKO3Zl9WL/Ohl/cD0yMit
FjBL24REU+aZ1rW3qoigUYlJ/OU/rN+cTBp1GPM7GO/hJCVCUuFDviKlx0z+aswP
sgCET2NtKiIcGL0ApWstrw0F50CQYM/99Vx4oinDPFH/9gWcT8/GmyyFBMORPGw1
bPVYvBri1t/X2UtMMCrvgZXxNhPz+V1WBSGtUIgkhJYyNwbXjN6Nkh/1e5kkUkdP
Z/Cauc1hCpsdKpQaYXxBFANdhy4bF12OlG/1XOgs4sRX3TstUW/ZXqgJtFr7laOp
n5ritKNTbdApziX9lCBchcyu6k8uyOk9eGVceNFrcIN/16GCb3j76857Md6sgrrh
qBz3l01mAWCtlBZtgtp6BF8UgYJsXmexISZ6hSIru2rAqgMZ60IjvB1PPxt5sBcP
q412VNIpN/o2w//W/pFTTRt6Ln2/ILWvPwHGN28KW0t5Q0YLs7QoiyxLokSrctSM
mw27F9VgOu3b/ZUmDPS8kKOzcO9PW/yxvVToZEKP/k1O6c5A+hooT9u5ToHOoQSl
PLFiV84n4Kt2VOKWp1hQHB38z0a0GKLTe9vtHN5xIrZtUJP1/X+l9yEfwb7zQr1j
LylBPNeHllJ2NA5V24cZ2kio6yjkzT2dsH2Gyuq3+gQvHpJChedx8gQU9LZRWJ2h
Th8K4RhoxF0eg5x41KaIDYGMith+bdj6LwnLPrVOpiL1pjvIc78fPJPEh0HlTIZ1
4QLjaN5iPRzWGzSXF70cTqh4VeCFqbQtk51yswupS8Edxkeo2ozTKOXItsCqfQg6
Q1eqehaJp+Yjiw+AdV39WcBLkzfy1DKovEoy9JhvoPdDzssiiu3l7OfMbczRrfwo
0qc+UdCtAtBeMaj0ijlAEqyIiX3M9Oyb2453DVPPdryiLPJIPkvG2aUJ27hBFsVf
h2vZoMBek2yufEJuu3Ng1dfO/rB/iV3lAVLBK3HoL7xkkgjMffr5GffxFuPVB0Gs
CTL58Ks9sS8a5LTSaWfh7ZkEZhCWd7bWgXkJRNQREZ5cJQK/RiIboJYL1yixcZDz
JRA4JT19BHHCYVVlMADXZMRpJ590TMIDDhZjM4Zd6I5jMsRlsHDfBSeCRvBmQOCt
09PTCSKrLtYRIJb1QYJGpdU4XUQh/zJS0/0gFMCMCGLuw67gplo4mcIFkwoW5fXe
VAJ+/4m7c7GHOpjt1haxHLLDg81V4TYlCyPZqVyxryto715g2ZIp+d1VcqViqUfl
1iXbo2ibEKuXnhDAE3EWe/PDxWHfi4qtCL7PZJPMkRf1geNh3jBV2hTCCsj43Vlp
xmYuje3p/ZwzoAYudD4s2CbIYn/SBvfjkQv6qsz+wIsFJ/Oncev80tfUQui6esJr
0Ob3u/3HsBqrGGq8ukPzsncjGDBNs58Jon83MQXDFZmZjNRnZYW/EUW5fm6XXFvj
WBYQlVRI6hSGDT1wBPeuDLl3qqcn5jwh62ATWBPeTGKSafOZGrQAZ95cwssoaAbv
RldDcdxc1RDIhERHNWSMjY4Vf9NlFM9knPcJ51ZxU+ToyelRtm4LF8jp9L7IuAnn
VDPeAA+LSUq7BHwIQCfasTTFtvh6WV/s5PIQYQgG7MUA77kvD5PE0/VfyIo0zIfL
+in2IaCKTvvAiOVfFAMV9vJGhd06Bgu8T+D8vFvm2tMm0RnMb/h82EDKGM+pIjzV
FY0BVyAGTOePa4FcxfdCprPjDkgwCahPTCfjBxqd7JuTfg+VNfowN3AazWmpVq2E
sUqHNYd+07Z9SED9XpBNW7InXkf+mEKqqlv02bovEEsp7FNPbxuapYbQdBJAjC/V
JbsWdlN3ZSAgL+m7V0raa1Mhf+9RQEKVUGP4lINM8S/z5UwEO6mDZDOlyyweb6MM
BiCeJc8/19X/qUDbFhSs6SPkyxUQ9QRcrMxrbEbR4EqP2nil132apJWJW242qWY9
RpUM9Gta1qN/JciNKoB+1JT+SfSDcVT9UK3hfDeD7DOKGbTxnywuvzreKB7bH0gx
gc8Bu/OOL4bLjkMIxTM4bzDMGNFweZRFRNiilNzblTWHemsfcN43FtmlAGNNlrbe
Ck5SmNqlnQ/CGn15J/E4btcyiX7O0rmmqZxPbmeJ2mwtmDMBHYcjtSNcQFHjUtt2
lgooq80d3QGKh50goM6ZYc0ziry3xL4QnI5B9sXGvxLo5f3SFSxWNVcqd/+dwEMB
QdviYKHcPBRRf49DvzPHutfTf7/BUlYZ4Gmu/mC7WCtv1fNAmzdpBnpO+f/WqmXH
CcbqyVxpE++fnIWOltYu/cuocQymVjWTz+zVlFQ3PLEFTqQZuQXXFdGSkp8LzygC
s0edtX8UeN5z7yGg/SVJ1wdsTFqOxdUiKAVlh8AuUJgmk62tGcMXi9kkC32nTXDZ
6iXI1XBVDbCIDAIDyebofrYD3QUR0Gqp67kS5kdGJuZ/EbLUO+6rcpaJAq0BgpLS
HTpRYkY9QDcYPhJ2KjN7c93Bi8olGcD6UkuhK9pyaB1Y9HIlqg0POba+IemQi/7t
MFz73egSf/mpf1JYt6hb8Sb3G7Qe5hadc9ZxLmXsYhVkvxtPYMJso4wJP1scqoLw
07AYJmdv/T1OYXxisPgWUvOpYu1IYGyxK+6aiDl4XNmQxPkad2DJd/zrHrDnjE0k
2wme6m2A7/YA5Eqg5yzOiVbrz/5XQhlIkOZ7F2TWx4k9o0s3GFz64WMSmkaiYKi2
x2w9H2coPVFpFJOLuOC9JQ8CA0bDGJ6uShkDRL2TXKI/8dPHStoCX7zsuRecgrbD
Jx0ZfZgLmHQzX0v5LasEnDpmYuZByG2z8sTGmv1aOBi63Cq0ea15MMemjRZpAAk7
FlSJBlTuYm3KKbBD/OIcqkxk5bDhk+H3h4xLGYGineCcmDqdO6OemgyOqmnKrS/n
TJr/TeWwwunoO42HJDtwJ69adFfZ5+gd/CzBI7/LGR00p7I5YNHAA/2oGY9ay/cc
MD/oQAdLZNqoVAwYUmZdbDqcpYOhwY8GiL+qsEVVMzODXVRIIB9sexI56gOM7Ljy
cKDf1KPAVnLvjIhpXDzTHkUonbrY7Z30/PQys6b7DL0drL0o2JMc5LJ1sKm28LvV
ZF6BjzOlpI7EXGgQ7gKcpi8VIx/Aue2CiVRa3biqSdyKQnho2fDoqGRCbDDq/ROg
kjzeuZZGb/jL6ltWNerkH62BL5D7zexFJu1IeNJ4LSoa6OdoHSSrHXIFhwonop7s
lySAaQ1Yhi72uVRQYSiUzUT3VMCJ336dk2HzVmPcF39TIrHWclIkmFkzYmnH7uxs
wzIEDnAe5I6BPxXWDlp8j0ycnBsaAhwz/UnwPHahVju+6FjXvws1xc2vhHVQbvDL
4jGV/H+EfXT27fIDy1TPSk5nSkUEoZPJgtfdMVr7QF3ew2yWWxKqeOKIhya4+a/4
g4dp7p+llaqA69xw4tJMKLL2c/fYQLfqwslxCgrdlFQaxueOZEp9pDnkkCrdzlQv
yOMiBDZoViZNAStgvG69Zk9/243VwRPZLcQWkdrM2NjoD5+KhCQn2cTzhESHOcB1
XU57d7nWMiC357aR5nZpVfh1nLhNqLv9COi8yoojw12hIun4v0MsypV+tC3/9Rf1
ntLYXDrd5uwxJb9seP0TYREjRgLeNyLizEi5Ppwz5JCNz4sZzt9eCmXi4KuZNvxV
ugkxuy2SDzLcglEoUUuVazahO0z0LNEXHUATMszVdWJmJVhm5ztd3X82JFqIJjWJ
0rTtm5EKTwaoRw2ayrlEYab7wviXQv2vx2ltUQoc9b70pqlBXRZ4isE6A/zAV2CD
yZEHos9BpXQnHfGfFzAy+QbBRutG0yGrAbamy7nNIA8bM3kEvjON87gOBZ/8yXJE
DMOkemVxrjpzU7pC+7enjPby6+lVuhMKOZnJ5KufRvt/n5FVBRxpc2Kv/7XjjAzp
nAoMjGB6GUGu7QYgrELoxS2OJbAzPdc2cYrHQvJd0Uj1m9nPBXhOaiD7Zbh52Ps6
IDpPGJZYKRC+ahtTzVnXHircHOSXOVgk/2ucZSjkgkvnFAA4h/axGcerT5OlRlIT
LGnxytpGJFfGAZitpRfWucZw9SXkseqbb8rk3PIzLu3+6RXzl/h0lg7W0HtRiBCw
A2dFztaMGfEtndtbO4cvTLjPqwooSU+h2+wya+QO1C5OOu+h4nYhMYtjdYUgakRF
AYDaTk80MvdJ0WFAZlMxAjvLrBNY0eP+hjIQ14KWL3XS7VDC6oXRcpN3bzxnlMCb
vMRC+3b+eo1xUNr+22MlvRZ4TBmP9H8ZaBFcivCXbbUbqZnAZJZ+0Lhs4yYvt7yy
L8j4FIrT9Zm12sux6XxV0nM2Fe9GNNv0VNSqP7qFWKT6DVjlpf2BK500rnL05GRh
rEPaF/Y9LTUXW0Fex0Kd9/7rGZO50u4MwvHxeTAhrN9yi68dSr5a3xJthBIWjMHA
W8SigAtFIIWji54lkKNgHW3TYabBogDJQA25lbueQzJEEDu1hK3HpxkPu6epzDrs
vFav2cHtn1qfbUiloGXVONed5scj9mC3h0H5L8BZFAuVIVSD1JiX+XEDfcqMuAvy
gocJASmQlFGAdAcopJYodHQTLRHZxxzu0FPN3eRuPv56XRT1AqBc+Oe32cWTYogG
BGMKFNE8f7vCZA7JIG1d6nv4QQaoQ09YvBiI/w9OQYdz0RbMl/h/j3fcS/+8ka8a
0gX70qWH95GPV3p5Q9/2j+LAXrknhq6Bq2vtt5XTp2XAbX27GqMKdf4820MUWTgs
q4ynvzZ6ml4b87eUDeumTNPNdd54P4ak+CZ9BRwLs+PXkIOUZKSJe3U6ouD6Hfo7
d11HQoCb7jOm6OiaKhIUEp3yhFML4o/B2BPIeiYmjZURfkZu3yIY3NNMJfSVj4hd
N59simLu1hzzqK7TFKmRAM2gCYvPwR3Lsmtbp6GgsX+AD8YYJr3R0zzzlWoDQUt/
AccyzsfPXWHbb3/JMzJFQYAODp6lLwR71dE0wAaEIgbwpkrhFOOiaCu09GH7Czod
kt8yIZd8vQUatM+l1sYfFHN3N4YHtQHIyA7WtUE4O9NW49GiJE1FNJSAX8/qky6m
BCTsQm/1zkUWu3HM5Nav3u9Q7eWuQ4G+vRXBwN9kNALuq4QVLzUdg9CMWKBhsQO7
M5+dL805Lr4hufOpomcEKIyXPEooMb1ElJi5yu8sj+6pLColFysXQh3Dt4Z1k5Zo
s0KGXKrcSGwiZodHzi/DxJZdzdFf6U+RvC8mbH4H+JSq1ESVmGPc58cypGCwjPVs
fspqigyTnQR8lR5TPyPvhKohZ29JaNKYTjK+RHDwUVYHPbcgBfKgx65AP8Z+jv9y
VSG5xJd3Rgb9LolJZvahPjM5q9oGkeuSrfP1x2r2ex57AM9DlRCwfPIhTU/K5GJG
10eEu1srxb19fkIxlc5v4kStlEKMf02Dh+Rrr5d4dSYnPN9tJMbSvt5orogcTXuv
zCHvlt/K46D6aUv4KAEi5HlKU3CKQHKJFhnsy4Q8L6ofycw5kCHlvJ70idvJRt3n
XvCp3US/bJcY1bYYHHzoMIjpBJwW0ltTKH9PJEtfT8mKqLJRwLOEbANEwotj1z3K
8MxUi3BbeRmyl/RLbWDPNjFih67Se1O71BKPQLaugRcsI80q5zR2Gfo2HJmAPZdi
cCzKd38NqBV0Wwx21aPnUuLQB9z8dUiK5BZ/cDQ8GJ+qQn48RYhYqL9pgSYS7+RF
p39BcN9CdzmTllpSszQRu2ifZdJGE3dgfftXzg+kIF+ixR+RvcShQrCdCPwKJtjD
z/Rw8Az7k0jCTkx8ZzDxxPWIslRYCYdOz6Oy//5c59lYvEoDtn2nnXLAFDCwzJSs
yJDGzWfDbTemCCfW2NbTesa6UoFCKXKRTsVN7c1X1PVP5sestMx0F34+IqDh5NXr
dffOUHhf8X8kgqjDEPdtxyVhAbsrCOVZIFzjDcGt3LcxWEf7vq/AIyFM+NtQaGU7
BkK9v66Qwe3BSBSEhG8ngyqmS3tTG6wi1RDvllIiBfZqibBKVGyrR9CDYYsmWzoR
jsbfR49IvODL+4K/wXvv62WUXdOPh+LYkaFTEJDGY/cYjHNUc/yjBRXUSirm9wQQ
73VfevcFiXV/MKaDCq8MifJ31zYYC8L7qiqqKdUpgR1HVjduCPXBsCaeKkVTWhcU
bo5us535X90791oqmcnPYR+2+1HGzNSOr65c5lgP72YW06k83pGck1uupWSI1Zrg
cwFq6yuOn+7MsupM/2qbV8pKI238yCemizYnMvFaS9PWavWujkkKIxGS35Nj9jvF
VCit+Wr1JxZ/8LuZrrMYfVonoWTlnrIRnNiUvbQYbbB0HpC+WtYfnJzTtSwj3Un0
RvHOH70naKCQXdgMdmxjomo9xHgEvIQG0TDSlzk5if89ZyzdGetA+loNKc/uQ7Nj
W07a+nLdlyjPCrv3lGf8PsPHqvFvhYxhzHaAJ27l3Wz+9FTmfTsOUdYTkjD8YhMK
Q8VAJwK6UixYwQTkajmnfz65c2fnQdv0daI89dqijWFX/wBfG980WUfStWfXPcTE
jHfqXFdK2W4YLhHeyBsRIFq4B1nryGDkzPa/bWG/NP+tDYe+JZbBB0kIEKIn2ZS1
1OJamvmrfNYaTf246er7adAF4mCXqlCIY6Qq2rWCP41nt6oHNZvViCtYQ1VjH409
SD5RLrx5iHplbef/czv9TCqIFIj39Vh4sMfMLowutICGhTHu85+WAtytFC9X1A6/
A9wayMKM549dwCqSTMFD4p8DEOohgfQyj2eHWB1YBZZYMFKP6FngSr5+yD65VVC+
7pCDhHk7yqOVtBgDT5WQgSUBHUCe7RKkeHWWwyo9SDYLnouwpw5pP6hAsa7p7AyV
wnKTzghRJ7yK6bp6rzF9KolSfKLoWMNUruOEz9gHyND/Fx7j9CsIeeXjc0/OaI7M
ayAPxSR45EMD3qFMkOLUbGifLv3SLYTSFwdi437355ah0YabXU6L9CaOjIC8nkc7
k3Ub8pMLlfxHi0RzbTe/Sid9Nevx0JLbkmFuDt9sG4Oic+j6HBcAahkoGi2h4gFh
qEfNhQVPT9UFTKj2oWA0L9JU7rSevJJmFJYWKe2lisyYvdZpH7RXIto+KswnzdSj
6LvVX4SMXlJvsRz9N9e7zCB6voUz1FMvhreK3fRdcnYWqKJ+sGpB0E0eDrZIVpw6
R3U8n6YqCKLhmtNDewI7SDseamL3xtijxXy7F1tUmUGDCoiB1pDgT+dx4nBFCIlY
/mKNcpvKQtqAYdtIBohYov3tXciV6Td1ca+wX/kMn+Wvba+qrd6MO7B50gOdkToA
6uXHrvxfzT1+6wqNtyL8iKa0yt4UB2YaE4kLmTCONpiuxpfs1C8uZre9jg93bEnY
3SDWYKbtztfzoENtZDMdZNjUnlmiJXhqCHSrK5hBtjUGeIxlaTpxnzkn/z2aDl5l
mJEGde5wv3ail6eUS4p1X3FXRj+Q07XfaJRfiCyZYxPwyU1ZQaJzfW5diAzElIFw
aWF8KFaPo6pCNvbozo9TL487n+1EkMtWzt30Q+PtHbdZu5c0Tb5Ek3tEWIbVbCqa
fW3X1bhT8lU7lQrLfqThbTxd3lyUOXe9YQS1WF41kRVAKyPjjAGonI4kxm7JCEfI
NX18YZ4HBS5gF3ayVxYPbDRWNNpAlwhMVxU9V2t817FtktG7kzv9kN0706XdGtBz
AvGxOr62s48JqVUaRyM0h2/98Ges1+UYwy4c9vOrQbWnXA+Kk6n9dA0no+JqeAXY
RW0YRXVk9wN5t1Vwz8bFeegSmYYwRuMIpL6mcMt75PAXgq53Q961195T19ah7yUh
gFWUoFf9lKDC7GjP5xuTH9F+o6xmHYJ1IX4Nb0tD5ZzB/myXwSzP1Fzu3tDXEfEb
diPsjttui1tAWNttwUsEjqRtSOuEHNynm1D1T/7UDMxNPM84D+rJELzKre80NbnP
XZ6ZRkntBAurleEj5P2PBmRzzYPtO4vmmok/l21XsFZTTl/U4Dj/KVkkdLuIaFhd
eG/urcvFAreR8IRnxDc4y5M52RPHH2DHPhyx0/M9y/8lo75N6PT+H/GhkG49+IDc
EDJo2qMYtEbIQeHD+dVRjAQeCV4BPeObUQrzRlZ0yAwSk4FwOGZ2ZBVlw6d1DPV0
eJ+mQv/aVavQzLz94cqTAgo38gkyS/8jV/YCDlgxKZxxCOqTETVBad287WUhKzXO
oSXd8uPt2JF0MzzlOLCF8EAAYv/nmeykM+1MzpzmeHrXgAtygo9W7jkUmFi2n8ax
0/F5cKTLJ+OikTwvtRUzcH1JYIZgMSbpVCGGWRw2bXC9n99nrN6+BRD8xoWLevl0
T27PJ8GsGDYdPDjCRbnaNdZc0O99qXvYDVXDs4vLeSVnGREcEVDsOOONgq56QcOm
KXarZZDbX0E9bxtUGY7J+Afvl4vn6lla8fhOMkKiI+XrEAD08kwWWU43yOuSHyxU
OU6x1AQpVns0LgTCUxUL9L3JbSPgW+VRqBARqFvzfm8hOLttiwFkcp5A+cKen5M+
8Z32MGDuGwSSf41QkWbmt/WG0X522eAsyKZlRCfJtMG6pKfHyUY1fALAPl/QlIYz
/FvHoQeV+mYhHbVFX7v25LbJ6/MIG9wgxeJ3vN/CNqZe9aE0c98yQdYCL6dkZHa0
iENawItQQD7Qg5E9FstMDvXY9EsfLndgXu2ibENJ01VTAjCHpPc2Im5R6duYdrjX
pXuZ2PVsA4dXcLW0STvJsMup3ToVrzcvpCvh2mQTKl3FoyEQZX/tO4Gop4P6wuh0
u/m1k+EMKzjM4/WnL7R119cBOHyOkD4RspSfAsDg9Ai6wpX5FrO/A2BtTmAZK7cB
bdztKdY4x9ZG6deOmcHCNjrTjCFWlFeriEUdUzxhrgdeRHglWRZ8agew6w/LG3xX
4x/zhA5hgdHLh1C8BghlWjw4SiNZnJluWq+zdOV+ipZF5nJUMepbxH3UWUv3bTiy
c2Vofvgr7ZXRYoK1Gh+IujGtwBilMUrdfjz7vUcHrVm1NcIvaDLk4iSCARFV5zTg
WxpmYaeFV53fn62Fsp/ojJW+6eXVl+HX53SUXZaEwtiBmUnsC16zgqydFUnxwIkP
NdUd1HhMcICX0AU/vn6CK12Zv19uv9sEoDRyL6lmRjQji+dqaq5NvvD86VfobWMd
Ja7EiOksZ6cOXTbteTkN7kN4ZryB8sKjzvoLqhJP49LXakf4aGDtw747JHu+nG7D
+btz/+LFsqY6NlS+E0yCpeQc0P1iRkykNo8/tdWWPgIAgVSH/HQIKe4XXISWlxO4
WxmgTeOeNUAWrhpmRW9zFT2hbcbsB2VOfzN+ZJtaN0gMFnG5+mo9GAYUYfvb/Av3
bbokB+mTlwRuEpaOYBWaiAfiO7cBovO4VYmxHjxfEjxZofbawMtZurC6PJWDM6zI
gFP8J2/HHNeBhHxRltnh6GfC++oXz9QEBG5HmEBsHHDFaEtRMKawfDRfxnXDpnYb
04n4rk/Uwu1rwdjtrhEvAcFbhC6GnyZZPF8TieBkPFF0i9j5WW9L+muWeAIDwziN
bSTqzoinbkWI1amY2paXeZ1Jz7gL/O5WBiRGoZA8wy+o1foF3ZaS1urCFD9hMGaf
zkucUqBvEzu1tyxow2t2HRxUSFZHMAYCyK5U9J4k96FEwmUHERnGZhYTnti6G6To
ZMe51u+Av1nz+6h6gUmFfFMkyY4bLLndIL7RdZsdSplurAABzhHtNPbkre260882
Yu/NIh4C3DfZhkXKGI4qmJ9m7kfW/6CNKsraOgd+ZJ1VrZjkV65FyF5+RUg3U2V2
+qiK2YrF8mwCrLUjph8lpBGdtBckgEAAVwej0O2FsOpcBK/b6+DUti0OYPQ4BBxR
TkoMxj7mhzDdn0lS9gAux8FPsHZtslu8RBhNq9FUDtek52BOx2yRb8s8bFUg2MWC
MoL+20SxcLeo972PNWmZzcDhBU5U5Eno9/Cj+9lc9+OSGFEquR+CnDYoPLqmktsy
Ps3jtHfbelHurmXV00SitWDuN2t2JRpku7bRUXaLppTdXRm+OHqwMOjwld2Hwe6p
OL7HTPXFV4Rmpgs1+FVAYENEcOw2hX+ezXd2AODfJ9Rhd7GAzttGa0UEHHe0cPde
b/GVqV7W1n8WY977CednuOINAKnoXuCHYRrt7orBE6xvjRqmXsP3vHB6YOXEiRQN
SU2ES3UYW15KdWTK4emNfdhP3xWBwoMgTFqMvZvuetM8JJMLIolywGrJ8WU2EAuC
65bTc+GC3fnf9GLOp6L2FeiQwxWKg/Jaanj234Z0A0EFn51+QqKLF1kreE+2VhVn
T0gaVG7eFsxF+IVcFL2OuJJEoG01zx5PKRMsj/mNjG1VUoF+IJlbhzkLZU8pL84f
wrFTnkdrjFMuup+BShqSB9/kitJCs0KISL58OzcJqDqcMnBHAWFp4WkX9EI/GkIz
adtmQJZfrKa9790eEdtn7iCbOYg5HDQ9xr3X6BJVHskXScpQL5qJ1tuAiPeMYmk/
vKJvRKmo/HAOzBO4F+atmaIl03JpDHbpKTWKRewtBDB1w5yZkih337Er2cqVNhq2
SFqK5eUylRbjPUHlLK2EL5eXM67BWEoFcDSWgJeMJ/aPhTYoRZ6plgofqUxqtM4Y
h/BAmMMnOUYobOZmkx2UVbZgncysAg02R6PoL4BXuX71GUDKUkM18Wn242NQbAMR
ZbxCxDlcVw74xoIOX09bbEKreJnquNeux1nWoAcQ9R0pmp+5fJ1xv+2w22IXqsaW
ikzT0EeQbNWgPbEwHxg6t/3rYkxe9z2StD+rRYBt2ZXr19mbXg+GbWONdqOwCS+9
fVFNWCQSMN8sMFHSvqjqZp02kI87UBofHb9VCHylxeL7X+qg0ngZhLGKHdCujDyF
kKG4MqHUqqKvkh0tjoz6j53wGs54ZJRFks940S4EMjfHcd6ylYVRkpIcE4H2tHWy
KL5TBiQxFqQgRs455a+bg2OIul/k2bnfrz5zvabnX7/xtLKUejIzptIWem8O6T+v
ZqrepjoAp1HdGEKIMx1LEngKtBwqicf0t242hlc08QBlwUXDFEKE24lu3NvM5EZV
Ifj4L7vB37YNUZ1kirFVhDGHmbh3pZg4zcKnC6/eikOSANwBF4TdbzinPBlvzp1/
VSo4Lv6w87uCyg1f5pmdOBVE/sEbXVsfEMGRTWFOBoCIrGEjqiJ/tVd/LaYEufE7
eVU55cUm3TMjW7q6BQCuY6iHip0ef1FYJuDeZUiql5+vqSl2bJnH74xTYhrIddYa
ASZrg+2F9OxfiAktO+uJL2xX5peOVHC+l2hkzoUu3byXIw6gKkQJkPB22pMPNted
XQm2t0MIVjXUMVZ0pFEZ15lka/T9oa79+Y9y9wjf7hjvfdE3UEwNuazBSef39Q0I
itpnRVjr42kU+2XW6ZKa2Y2ITncpjbjbYY0rR77Mr5o5EBuAv9yTWvXaW1PKCjy2
VjV8vIS3OyDpmnAP+XdyHSJsXvSFyo52ogplysjAftAVo1bqq1dKSQCVjF2gNS7k
7cGM4zIRC9kK+3c6Z4Pd2wpQhINvA68dSq91DehF+kQC0S5S10NG2jMt4QOpcWd7
TUBnaocWczgljWQJhGZcJxMe5QyiLm+slqUiA5YiOihniqrReKefxMwBgAC/brCr
D3kjQsqHJZThmMA6qOu/KOwWUrEM01/VZp8h634g0O1bEDfw6h8vWy+fzgYADq3y
rq9yVOyvQ5ELZ1TedYqWKuOVtpPsdWwEnQO9ikGtqQGsiWnwDvS93swzAKjc0OEY
iojQoK1YzQZw/zDyrJI0OUF09YM0wAmyDZjdEq5wE51PA70cM5EKCSLJO70Pd1/M
ES6iVmiFw560p7+ybKU7d2Dw6aIzJzLJPC4jdweJ9fJJO3PhEsWtXITJKPQz3gpB
BxhvybfKeU2y3f+W53E1DJMbbix/t4UFRoKM05LDf52NRVOP8q2vk9gPyyzzq6dl
9QlKktGdwdijss38IrG8yTaab8QURO1i2lXPjw8JzJMnSdX2+Xww+uO1vY4TmqEY
8socMeW/F7REHKW+pty7xwKq3kJ9E08Vj7xjjzEHSIiC5cR09zJF9kzUVbcV5wkG
Tesj1ZTpM8GWxqa2tEBFOW/ArjatMOxQF63p+JYW/a04G6U/eiM/rG3pR4fNi135
b2JQ2cyKuXMANBxHKRL2DBxAj7Sua9tZ66nC+F9oG5qqexKIuWnAQVWWHi84uTck
XxkDDYw+gfyKfi07yUxDjitOWCkf12yuEqq5+NHpUS5DCUwA3CRz6TIy+kdw/DOY
DN7B0t08itPBBG66A2khdcTjkE0i5elgchXxa1QVdKzFkbbesMOamd3fM9hPFpnp
seKBUwfAttSZGLux8AnBgQt760a8rDDqUZ47MBU+QuUQgwXOx/E/3jm1u3rdQ+Z8
DXVZP16DdciOF13opp9vHMM3PdHdFPvmFt0FJeTDcPgm0zpFW9VAip+K7MuYuKDg
OiOcqodaKGoItrA2PjPr5Mfs8Ze5V9Nq++DH7bUOEm9+PR7V34bhsijSyAh1XgTz
179v0nodBgJ6o79pVshWJycZ2NmVybjaCl/hr9jXmArs2ym6X5mm6wnD3kUVJJKO
A1mPwlooho1eVKlbhUn1SPKyUGkT/Gca7lCh484nECyqWLyMznMtPthY9SigialV
GUDAX5qhUJgSgHNl1N9saQ8pXwBeRM0RJatazqhdH5+Umy5UxF3nccG35inLJkCd
ZyFuS5cytHGbeUtUJH2I/WYCtrHB6fJEaYwKVhajEqOfOkSpNUsaoKYXU4qj4fsA
yzy04+LgKx/wMVXIGNLtkIeP2EVyq9JL8v1f7Lr4LYykHQlEFdO9hZpoumWrNMik
mZeTv6v+VWU5k0qdk7TLuJbpjyPYj5wFuHL4ZnudYtur4hvpFkPAf0hd1oXt7fX5
0IFvfbIQ99cjW1cisRbvliC7elIkN0mBZFUaDtdFM1skQ9wXPfv21anaXKLQ5OXS
YdBMlgmSgmqf/DmMBI4AHq0pGqAPLA5bY5S5POm3JTUGITl7NRewn37h/MF5v0Ze
n9aOH80ACuDiw4j4OEezyYKSXbQ/uxwQ+vJ5ezV15ru1v65V68xhj86t1AnGCEQX
LK5qJOHFOq80vHdiLo9gH+vNm5PRGUpSIjmp/XA427Zhe+75mZxgkRTFGuY5tqZ/
9qpu/yEW8LgSJ3qrGN/YByKJXY/aFZlsZcCfQ8YXFYHuqUVkQL909s+hsuTv9xMy
695qtYJ53gKccN33uNGUJ+zk+Z6Hu9VLB/v5BX61dkLhY2a3/TswbcDnJb5yvtrY
yM9YLQXpijipIgGLfiq2K0fuRTxpW6dSOoi8Mr5cq6ZGHajrY6xjhPnlx2ehWydX
g4KlXfcEl1witnhbN+rU1fjWFtR+iJ1jwXqyIjRSYd/giOvE5Ha+By8gur9sDgE0
5wbgYP8iVgAUAdLQYynie9ECNrczQzgKsoybcqVLdfXJ7+4nE9GmOPAdsAFW7awL
IlcDOkDiWcsgcqTSni7m9KwHaEFOFkK/Y5kW0WY9tnssnaIiJKKsUDrCZMkJdQXz
i8TqPLjdmdi68Ic/WSV2tfrE3JnBGZEfzPKeiCc3KFAYGNKkCWa+HRb5HmmTS66M
7YNlUD5r0v9pMJZHSF3GFx+NMcvwj4nUYhju4w0W0ThMNtcG+2nKfAV14LC6jXOe
vTjgS8WBdtOWT6Lv9P4JRFwCY+QtFFVYSqfQZGd4jnBn2t6yhwFv+aEh77bW+MJz
dQTo1UxwMdCp45ALGhC6B4YptMftQtU8J1EboR41UbADMlfX25hb5R2YtF2sVUrN
sKzeol3jbnoqKUKzkTAY5dcRlYRL8ix+thud0wqgdAsdW3vUdKh3YyE1BT/eEomL
o7Bq9bSBUpxarVQoJwNiAjKL/N11UuuhFAdbyCFyHafKi/H4cRVHLIj9jOqIa/1J
SziUGs1jabukZfbRs1npirtPyAr3W0vH65lomKpSGkI2y8wyWJHdEap5byROAlVz
HWtPgLIOXeG6hsCHK7JsICPCuOYEyIpLnRF656HAsdsQFJqIwzTq6VS8S6JaxEFS
ev4ew7F9el5QVEKQB/IXjNFYbTmCAXruBXPuQXaHzIqrpu/bukUalYPKlG8POOoM
zcdul7f/ShtkWqJB96gRtI+hRCBrn0VaXtBRjLE/TcOhNCDAcZwunwcHzJZ9qvtD
fB48ooaaWTippqK2T2YDyXyRVBx9V7UFTu+F27rA8ZH15URV0sT4N5kATKUONTYa
YQqoSpvJ1zQd8s8fOwjPS1vf+WH6aOn2UCmML5J431qKUDXPXKuj6wf/1UqEZZ39
Nb9kTd4doGUtSsUnPtcJ/ofTSSzTdZKluYsT1VfvDE324ymVIj2lOt5WVTdEx0zW
NDgjgOgrmOziY3hJEn0ByxP0y0IHt+3RGKzStNnSqp1vvXGbEJcSCBnnS/XiSsPF
QBLWzGAt/QZj7pXwaJp9MTNIv7zLjTfjVq8mNnqDLIOA1onLItTydT+1yjqa+IIf
TDvgWAqZKhu8XalE7/NTjCdW7JbmNKsAZCuCPKDrznlnaSm+rj62xY36JvggbY9z
866THCfMM6Y3n6OMVMq8RWQzi61RMrTOiCc1wQL60D+DEjbxKZCkODrY0yW2SDzX
FmwskMfi3T5FZo8wHcbAtlw0EB5BeRl6oH4Or+HTTxhzKGMC3TcK8DRz+Taqrk9i
pJltIHgNkn9Rs4RhbSxLyC6EVEs3eHQNmUMNq5FnSZV2Ih1BG5cWO9aCwFLXF3Xq
Z2XSjF8C5q2Ud1XuJZEEb/GzQqcrVWT9dOAKGcCu7xqwT3DHEMjotjrqwFqBHllA
YcaAnyvORqzsOzcWjQTmahajgT/suay2fC9uutU7bjo550eK6lfPvTDK3r7dc4tH
Nc+bD4gA1P4EijhikaXHtDXACF4wc/1HVzoSLtZnhfKfVUHWUy+6hPWQ8LgGshrp
OjdIcKhVGrA3JwFaL3mLpZp831P0+lfg+pg7Wc2X7hVwiPOS2JXtfoGaIM6U5ni3
M31Jj3SAcZUIJIdNeXm55dlO1SPQ8vI3bZ8YPg+ryw5tMRiLa488R5sA1OyoUD0e
SxoOoqHmt6ZaOHGNOMXsMXcnEjmL8GbwDQbg1Gcxh+oBZgmc/m1dPPL4Bxf0gMEv
RPQkreF0rjWFpCoRGEdJLDcC3AHblVhl9QBrnYwU+mlKLwTNe8RwH+vrikUEeltq
G62jjIg2yb9wFtHENnElNOOMsDB6B160xk9Zd/5JGk95wyY7QT0ocHFlDYZ4c8eN
HJXMyHI/I0jbhLWGVSJUCIAEfDpZgv/MgzGOEqqyN4dMFxzjjtVRPqc7KYswyf5R
yIW+M1LC9c4XrxbrdfEOy0+/eMwWTMeDSofx2ZfLiX6uOnKYn60+fkozHcG2yby8
Mk4POzWevLoeRt5eUdl4FY7RJ3OwviZ/mBNkpgtKOD9Vw8G/3f7c6BiOPAuJqEgT
7ZSdSKSHGfY35tv5Hvh2HBY2IbiAoNCzSxRd5RI/Bj4SnAF+FLqAUEkx6vkqdpQC
qH6T1gOXBdnUtrcMNY7KCDH+m9CLKRw2/v1zKBxGIwEmDPmA5ySODY2yRKwOfenA
XuvxacH7LjHVrCwwLRB5BUCZIYHXIAt8ZMFoZPRZNdYwIJqNe12wbRycCi23jJvk
/NzXBM/B1tkO20kFrSc/zLEuYDhA3N7DZOh+yKIRO9sEUES0teS1jgK82xU5tvVw
pE3PddJR4lxLuLKxTplLpMp1YtgAWOefjq/1iePTWFcWY7Bi6VD4sIzp3uESI0fv
Kkb9I2/Z6KUELStm1aNEJFmBrXzpcGBGHsesqokBcP13uSZlT+QC5uIRbJBOPoYf
DbhIBSy+wjB96t8ZVNIC0TJX7dnW3f1YlsqB1BTw4buTyVtdSYWOXH/KmfOFmhdc
oXw2Yo74yaGoMfBE1W2Feunq9MoijjqZ0qwZ5cuAk0zdbuKMpN2nRsP1ofgSSjpX
KIWdn95Muq6UOEGP3OTXNqrGCofZurrehuwFaYFyrIzgDrWRPe4mxdU7JhceSFQF
wkBAtNSpncbGa6IxEzejmACRjw1uXxeg80YaPqhrUJyXIxSyGi6fg26so39qvOri
x57vBbtbPptUWAkPzUnqBXZlD3NDdyWfcrLnaRBg4X6yluxGErseTjfvGc7WkK8v
5Fg+i0Rag6oWOOnN+p56XbI8WzX01cHzSf3it712zDLw7ttGeDUTYL4vjtw8fav+
wZm02mAFXmrbjrI27pZlanMIOUMoUe4Dn5R0+3xwWriJuA4V8OIftH2KF/56vsgg
I3xBb2SF2/cOsFxhjPCGUOTxSgieD7/fnYHoUM780zkXLS+Y5G4Pa1pT9Nkrlrsy
wl3v916p5sT9kmMdyxf3S0Xc/2uM+rNLwG8n8xka1uLv+9y/eUTMLV+WAUisY2u7
EHtXnXxyu7m+OWyFQNNRStOdvWNx7RzAkD7rn74+/uqxMmvD/vR4U6gww4J8OJ/u
W1i7ZUHk6sx8x6NG5xfGgqXR5XcWD8s10znpIfzjSXfaF+VeW3V6fdg1Idu3hicU
ZISqYPNAYpvWm6FSBxnOaFkzaURGrgHULKnReOWtlDJ2N2jJqfdRKjhSzagqG5Uj
R3BrUJ9b1eBFwqmQfdsUxepjA78+Kq/3SDSs0VsGxikUoZI3DYNjmUkyFsJUAgIc
pJiNxp23I57UZgeR+O7MYlGgb7juFwSB71QOE2f9URctUOsRLL7EGyDPG+nwe98d
HYzO3BDiROxqZkfLHfl5Ym961XsX1Qi8imNP23ROd032XY4SKcE2ZQXLmk0ijPaQ
KjaqOpTI+aKgqzjySQI0C6o1adn+o91Nwuh2LevucAR4Jy53Zh9YNF71QxNKt8/i
fzch65MUyf35Quj0ZV12fBWbNlKYMGiIDLcoW1PR9BLBMgnM4UrAA8XcyFsNRFzy
5g3tkeMp176Qeqhgz89Xra9sh1+UoKSCDq2rTOMph+onMVSyYOCjSfPnGPgkIYh8
YdoZGa+E3m569KHYWnQ5bZozz2bYRawoSzKv74cB+nPXhIOrydAx16n5EicdOusU
hpu8y5JlH1318z7W1IxTV2dDddOsh9EI5+hDq7UhgL1Zmjd7aIvnaGnW9S1AKhpv
x+8M3j9/t9dWoinib0nOPbmP3WHBfVJdilbOXSEJH2uwFWB33UTxJjfMCEfH68IL
87a2gyvjvO/TiR7lSA9Kcnhqg8UPcc/Yj8BHGVoaLueKf0peXC+Whlqy4tQ6ulyV
UcUdM5OYn/V5a1bsgz9ARFv9yWgfSQWSHRnmgPuwum6x0GyifzQ0vvA0l257tzGz
iJCwWk99EGJglR5wuwO6pZ04zZ0rvHrvj/yybMoXDMaVFbOyIySkvp+laHknml+l
RDA+iryFBjIA4meSPuDmIw7bs+jQxMhzzAUHLV8rFY2vNRXafml1CP6khKi8tqOP
/pf3iyPm/TO+JauEMGs/u4vl/NGa0TjvuosxbSmxB4NBNCR29ICIU5v0/6y46r97
Bl0lLEWd8jyIceS6EoNL/1mCCmChkXkVfcXcUuY7/TZGkZ67j+TXzYUPDporWJa/
8X5l9w2PxpD8H0dNlTfi1mMgcIPGGml+/dCVVqEqRJwX16eFBNCxyDfw1ZjRx4JE
YdPW28wkCTHJm3gAT69P8/E7417aznxoTvQhSr/03Z4zkQ6LUKSAryMWJUamEu+r
945Ctid/WXUFJQ67W9xQBtKwt5ugF8LXcjzOlVZYlvlX5okePfzL3uzk+sjjzBpu
T2n8WbYbnG68tbug9KO4Y67ii2GvVGoWHWTIL0p9z68VueZIX77KPY4MiY69gg3y
ezWkseIDdx+LrAA0lP7V4JDHGN2YaUo8git/CAPW4cd7ngya1JpuE4sy/IEvQZ3n
mXZXTf02O9usBOpUN7+7XalAocYQCDJWpDBoF/pfwtGWf6wNKWyX0Z0+7ep9Zj9r
OVL1Oj0Aio62gkGJeHGz5IGf9LZ4D2osIevp0GhJZK2L/JzckrkIf2BTTbk+y1Oz
HH/TNMdJmc4sU7Lf34pIPRV2Y6WyHXyhPN7Ct/qgTWwJcWMH9d3L9fQeHXKL+JQ7
JSZkdDc4B1r+9Z4VZ0UE1HjWDVMXnKvcjEASpCormphFy7I5IXJM5YpmI300WDWu
f1MIRq/GlNbC+HjugZ7uTzQCJcSD6Ghu3OU9uIkANNmU3O02Al4cNzxN2b9GT03V
dEeV7DLR0pUoXPY4b9hxnbgwMnGztk4zkUAZvJBhSciqIszAIx/hHG20i62FAHpD
ULMU8nvfet02Y1h9j6Jo532Z+jrOjuzSL37kmD5j9PsSvNKNGxjC4Jsy6lGvZinN
FLmrZcuVvdAgN7s4dlzZBeKWoBsxf/cr8aaAGcxt7/ZCbnKdvc9ld5Q8ygKkOZ6D
JwHWdE3m6MslFS9s5rayg/fgMG5PtWLj/ItRUKiQI1VhTOVytN/MDqPBCnx820IP
X9O1Mw65Qi1JHncmrGsg3Zr0/McHgkAoSmQQmSNRSf/WWso6Oi7w5+cQ5aghZQqA
G66iSdgBaU/PLHFRxuY60cSY/qe1EA0cAnUOI+rB8uvx448uGYV+Q89q34rcDINv
wHh+Gw6GP3PjVSfLc5rhAjy+aNYqs9yKlCOPt2Zk42ZuPxTTZ42wpriZ8R6G/FEd
M+LrYLiizyJ5kw6qmCUFQT6tyejYzPxmKEbN35RoMps9+8fXBAMix5mUjMFEV6dX
iYuxNYOOPc6YdVAwzRwv+ZkP4tMwwrhIZelnpeqY8Yv00QutVQTcds5RRsXeKX++
H6Vr7JZuKTiMhuJBlwcIiBJ2Fh+i7sjDAxfi3sob/l5AdpjMGZi7w/at5ZOyGqoG
kqesQywh+ICKngnBVJoHjpWNi+OUNJ8anIN/gRyFNQt1iVlh5/yzKBJJibKDwIii
sTGfaoYu6SFwc6lyay4LWwgFDCXI4+TeaKGGxLb5tarq8QJbMB6RCWLdsCaUumaU
+6IuxJXCygbvim2QaZHzQpUhvOccU7VXlQ+GHd67JzhLNBtB0jSTyNGp9g+Kw3QW
K9SLbZ3mvxBmsIPCvsyeBO0fi0M/DSI8uSvj46cl8EOzaPgL9MM8bLv0798xbXX3
Fqhg6m4D4zc7P/AgLBzjXyHn4CbVxwAcrD5ycV/VrNqGVZVgdQuiaQhdohqeJION
0ZcZyuUUoZu32o4nHo1Dye9pu58Iudw0LUxUDp2v42mpgPRj0uGrJ2lFLW+rdNvo
dQOsC9sgxrxJj+d+LM3vS4jTj22Min/BvkgSAMAcG5jK906OGL0T3ZdQ/11SOp38
88h9L5jtY2Ck2MTArujdcydA3HxNDThYZ2UEssJdNHcXbM3nJPP1mxvcsslc9hV8
WdhH48wmIUtCZYlN8PE/vWW5vHx97jj71crhExe9Xg6H4EuxZx0ADtpA/h7M37iV
UckAUyoMC7qoIubTJrb9uckcZTaynQP6AGSZw/8++s73LF0ynHyZe5vzxjwXFjVS
Fzk93G5C0D2RTzoi6H53e6kxzXvq9Y0U4/Fqw4J8kexXohTVBPUJh7A22P/hLRxS
7ubM8VuME8ibx//GeWfApSWlp8MDALKaVQdOeZSzOSOXRlbHHsERS7kg521MPAze
cWwO31dbp6sY816U+ozc72h0UttWk//ZbAKh1p8hfBTOzHsA8FHKmuY1SSgnVXU1
q9RQWr3Ln9EvOW1DZh51KE9rawkr5TAl/lmcqxwOvwwRd/YdqZp93PDZwOmcSMeJ
G/Ue1e0QrXssvnLEkBk7aZl5MRvHsmtPJYa92UMKwvhlbEi2jigDol0at6wdajtT
B3BjEWRuM+3Jj01a+10bRmSb/xjlgWmG8D1M/OIcx2XR+e1KH3rNeGTEK+p+4P7p
Zu3V0RiC7FrHRk6MVd/x+aVUR83WeysaVDEmamcIM56sopVNiFfkYuUFaND+1EMQ
cidWCR/spPEQQNvjzvRp/ztVwKWQuAJaCKbcoyjZux7CTkDpjBqZlTQaKrIpW1V4
z+/NhdXyFjh83HL7anEkle15nNpfJMIbhfj6CaoHuUigDCFR4KLam0kXRCBE2ChN
WkBbRvG8MMACKeLybQv9P963YjWDO2fJNxPfZTBxA//V+ZGUkQzMKzXS0OaxqCoS
KtSFdwymdMDiGSc9hBmGHZbQj9JFP87oy5crK9livYr6op06Dkwf5cWTgiFIPrzL
w2qnfvAX6rJjwWUw1vSO/XNit2BhbF+LeWm+L1s5A4y3K5blNnS0AX7sdGUAuZlX
zaILcBucVw+hjey4KsKlOYX5rdlj5Kehha2mmPKv4wi76bA0ZcLSxmhw+jTprRcU
mBJV8FOWw0/yd2gV4kvFxItTAwQ0GboQoKcTT+ClqTWfYyYzUu0NHER0fFUs2//9
XjYZVRM6F54qBj/LpJBLbvMuAptn0fv9Jl8qwIfxeA3kGabtk1K9Wj7b7ryAP67S
prMVnEzZ4IfvEqNyrhK/ZCWMYYhyQBGvpyEOEM8e4rxd+6d80Z2fuK5MwJ5Zjx+R
HDwSSnM+K53mLQM2h/gVe8ye0OYeOqjDgJCO3wObpkuLT/4FDLQOdxlhfmgknkvg
qMaS4sinHc+eHy7A6eANRE0FjXTuTHaeA0IVOhSup4pf6tK2MiBckbe3pzaFFA6/
Tk5wsLel9u3dZvaMFDyTDQNfNy24RGiL5EziVMbLwEMKtCGxVKiRikp9lDR7uJQc
/v+ttcQChRXfTE+bOvW4D1CLM78H0Y6k1/ow/5sZQvdu9WafPSd2/8QfNHmAKh1P
PG7zMgS+6swlkT8a+wd9ABZIp477rjdlKYvv1yYQOmWCT8F+Zwy5XMlSkqBtc8eZ
oLPZeouU1nmbp77imC4mmzKkwMA7XfoHJBjHCSsMfO8ichX9XXU4uMTl/HaD8wj3
z67i9ZPVAIAbqymMGdLElWh9RuwZWcP2yDg6hlW9mUcoo65vfEqba4bP5WtmlFRH
l5YTrCs6sMUwiLj4jruwVJER+3IOaFMyrb5nx9UdhtJIfq95J31BsSxW3RuzZXKv
o3TH5qC2SH9VfP6p083sk5bTXQ6Fk8lPTHS03R2XHxEi2eeT9cue/+j3Ni9nPErW
qOCl7B297/XZNurwBxJxxwhjB5f09omDDVAQXjj4nsCgemcsAc3rD3jnL6NgpmCC
WbGn6F1aMUm6/UxtWxJqcHHyDbHWiq2ULrH+q02jjEfQoeV44gSXEJRuBUic95Qn
x3ijYbHYq4/Iw/KiiNjxkPsVE9HSPxM1Kat9XHKbyXh+Wg6btCXFFsWBnPd3voJd
rPqqh/CPy59uQVCzNyIBWTZxdmJrHxnWavOW9ec9NtUJvQg/MARDYc7SPgstU2O7
0W9DsH3W2iHMkwPsg5V4yExqdBQ0NxJwiKPzrASZ+B+Fq4dFA23LqSPOnoqoc950
XhSFwcm8vDO2F8OGFDYmXyUr81VS+Gxgte+IV6/Jd8TLtQaFECVSdScm9FujEmoB
DVyWyHOOiFb7yUP0BjEwl9lUhaYCnfOBPQJ9acZl7IYAT6YGGj7fa8Km4/Oe2srx
Ftl8kbX8J6W1eW8ahZhKcddsfEufTLYttMDJTPuR20H8MOD7KnL1cL5N+Qp0O+Ol
pbn3EysI4x3psMjNjRxBfNsWKXN0tpfldIoH50HVrgPNi164M5X3jV85VmMFuuuX
nVWwLxsAHn2UiU/yY7jFIG2iYtsUAMaxbagGmqBYS+tqy9O1mvQiSORZJ9ATsjlL
GcIi2wfukiOR6VsBIrvJu1kajwbTJzVtdwrDGrpKBy79PclIw5c8XoDe6i6BTtoI
COCNW8uPok21wxNVEIdo7RjmPlez0USudJTstJ+VWAU7XDP9VTdsGyM6/pqniu39
Pz+CdLhnv2l7gfD9SiFEurxsg6OVFYdUS97JQ3HHNWtp5QYEX6YoRw3OgblhHlmP
90wHJnfiKYnzC8xqBfOMhp1t71NiDU4Gqh6Y4VZNnFmJVRNxnnZCyrA2zBoQKnjd
TUuefAFbWsT2j2CgS/0W0F/HODzLwMLul4YtbP0MwCgkfLcXMoFO6HpCuVM5wz0v
YvImsuKY1k0Vu655Gg5WZ0q0DytDX8LAglwHnrAHVYtg6Y9faONJWzimOAsWoRaI
eJ0n9qt52r69VG9OBEV/wUEE6dTN5RGXToD8m1vXiqjipI42Esv18gcqg0eTWHkG
8F1G7aspAm5gDRXdaKJgb19BO4RjHHZygwAHK8DjfypA1x8W98q24FHvGlenTA6m
N/OZQy+cGf6ZmyfLrIde1AJ80DAP7/6CAxadTlBMhXYLdp7F1Zqy1nTEVb5iSqlK
Ilq4cZAknwAjrv7IcqYMSf7q+UIgA/nESXjaB6S39YgpH6nJS+vus4hWMmw2Pc9m
/LOyqiqdrmYiL8N1wURl7TEQrFKg7v8TeT91frw+0SiYhTwgpPeAVL4Nk0rmEius
z55lEBqvPAXvx+w3sZJ6z1sjIytj+CkUka41rRj5MO6sHynmx+hNpgYbm1lUxN5O
6qCtAyoJY4ZzLO+f3Q+eDuu+d/LI3oCSokgITlJYMOdO/wcNAc0XT6dhBvdZKE6S
ZpA12N+x0Ks/1HX4S4ybB7W3ioez+MKNCZijkREdC6TFGFkLK843bcSUgufjV2oP
0wTqbETnbWuRQSsyOlIFqbYOodmEC/hu7aMMvP9E/pcqL20O8+l3YgIiAGxyG6Wf
0GwgynGCaxDPg7uWblz+5kZcT7nHlzEBGW7Q8Ve96HIYYFDYaKc8T4U7nzaD+IrY
8NvEMfnbY04CYxGsODS97X+4d9dK+BfIjMJjT2pF7n10sCEpw2nWsJ3/5vKA0hbB
yxVYgDMFChTLH3KAtuRR4ule5cTDWtSMa+/GVa+YNt8BRWEIJUtUw6FQwMABJar8
19Mbd3hE56pDnsUNo4HwilfLHoE3QSTLinjrTFLvZlOR6da8J8rgoNHiIB7TZ3U5
8BH5cvxPqDYsMu+WrvESTOngpOIgWk83azo6O7D3GTPmOCI1av94ahcn30fZnerY
c1YKJlM90llsJWNcDyi6THhyPdNVEQDrfI+oF4XS3LS318VPpf5BYIpwD9MMPFZ9
Zu2L/NHdUjP7KC1S4iWXxd6IQlf+dCA0cD6rMYepiKNtDTGkXV1mwePR+KekvE/i
OgVKAtqD1qiVM4Bt3SdL2Cl804UJL+/Bl8rvQAKgGeVF/ZUqtE1th6hjnyrvDdD/
DvoSTFNH0wZFDPN56VjVZ4v1JXqrs+gRb9TbLpjtkjBXu20XrhUfuMAeAfMxbc0g
ec/2tQ9rH2Vo4fVoOSDx3i0cBNPWafwQtO8XUlNHYEo4/ALCkDvxKUUc2j3+3+8Q
eV9/BKjk9Yi9fFaIFBamd4YH9rNyVSGvSN8VbqG01s8JIS0WuWWaj+8XNsK+bSf7
s6TSTCtGEVVH4O84P4aMPeLYtvO09IZ+UguMI5pPg8ul+/Axo3dTwD5gLRAa18Nc
j8kPMsA+YRCoSNCjvxf5R7woVtQnEO7ma/tYjJLd3LUOX9n0MGucbDne4ol5zBpC
z9LxcQh1fWUyimHzL/l3BUmC5pHMoshYsmrwwwqI+j/sY0irfCMyMj5RgZPIKzb/
SoWYzTR1L5Debd0TWyoiaRI9rDnTTwpJPv87Yl3GXEWT5maHwb7A4lT2PJVNk6uz
TXIsqcNfsNWHpiW636b3LAoNoEq0DbL3VJmX2DzIuGkV0kzuRSA6Tha7PItzWCu7
q7sYQxTUYgjMNKZBncauwGNsm84HVfNSFk1M+icur9HgPbZLQbumM3FH6V5MMuQj
dZQB5yObjfW+kCwfxFgw44K5LhSoJ9pS+PcdcdEJyRFWjf0ZQEVkIzwkIGRIqWeo
xrNHifP2lI/EkBrAlB16RZM9uMGYoIpZsE6TLJ0IetDdmKW03QZapa2T0Un/b3a9
SboqjUWRSHvDwICEhkkhwIfpJcTHG2J3sz7P/Xjg/oIWmw/FSf0zkEjwef/6sL2V
hdm4XL8a/++zCWXQjvV5DKib75jZmuEdsnEs5eJkoFkmdDnNjE/KNLaIUGdlsx8T
HIsvd7OhQP53g4l78ww6j5N5oGtBXCt6cxs2Bb+ejS8HqItHOBGRD2g1U0xzMysm
lkDGA4ZAvFlBnlW2iBJ0QXWED8EMt1FHRMeGSW5JVob6T+nKTMSp3FUyAn4G7lcN
HqdM5B2ycR5NBKqEHgLGbXfSjkreVVdSssYzboHQ+ItNBU7TOH8xjD7kOStZy78I
2qXgk7L59H+AxUOLzxV2rYpZgxjApkGJHrEjvREe8pY5VIO1wkfY9Mtsr9QmKLb0
vxVrgAmcxGOs8JoNbssGciULp4Z3WVEaSE1IVeIAXR3kYnKDiPDcFoubtYdPRCw2
xhB4DxUl3sphFnd+wW2TbbGez3Uz/JOOAuOwN5sLeEshj4mV6bQEnJ4LC6VwtCzW
26tfEed2FIlx1xK0bl/LH1R+bVC93HNlH8nM4dhjxmy9NOafAViV252ukwUMvO9N
1xBL+nPD43uLREHoWwZhQ4UXXF78JwU4mx2UXZztf4Woi/56hJb3M0aaEQlX2UsT
ami9DMY04y+gKspl2DpC7+4od3lZCvhs3wQuuWvIgEQ1AtgjyDNAHgRQkY0Oplma
nmE2ikMeOHlJ2RTXmYRIYplt3/8Lku2ZLUQrR/m9UXatJ1NmaMgbW7t8zDwqX3nc
q+TEaxjDLU5I2AUwePinze6fCp923Am8CHdhWB8z1fYEMEZP4scQJTx0t8vXw64y
cX/Z2tRsftVqXe3N8Mzk+6R9m028QAAK8DvAiHi9IYhTto8mosSZkIj7iBKBtqbk
9jz+Zd2fjd58kJG/eso2yMLhOAtfoKtYdyE+Bjo/CGtYEkVKTz3NRyVKs9PYOMEL
po0c/Kw4M+GxQxe9nPo+p7+LguJWFS9O+SRWO4x41rCmRDppEP/gq4EE3S2rGzrE
Xgl9bnOeDCAdSZpqnTK1TV2c9hbX/D77AusHjz/AzwCCohMV2Kck6bcJLQyFvkfH
DL64eKqa8efbsBwe7mS/uubYnSrs+zcbEvrf1twutqXWEEswdDlL6cc8dDdYILru
KVpaH70Rh4d2k7QIG1U8hEXmQ2goYnvd4K0FaC3GC664cCKGEp5CvO5JCVA7nVKb
0LcHqOY9XEsocHFBnEsWrdr/IK4Pcmti7yjAeb0V34zKlAeK3NB5aSQVKPVaX4V8
V//Zjul/RA0y94MdbOSj89AinM8ovR5kdptqmVtiWPraOD2Vyi6TkJBL0DmiqOlM
4inWiFp1Z4rIHtlWTiHA8i2i1BN1M4ZG0SN/S4Bqd3XK+wrAsByzEQcGK9qANgy8
n25SEEzp8XOg65bF0oVfZsgoEM+zecJAubWMbNaF0uo5MK5erg7J7uCoCEHnhgnS
VyzkZ0dx+WIda1aeYE/XPR6x+37GZUFN1kufh4kVKLWjX7+wWMFI2gwRQ5shclco
avtNRWfArfjvavRURfokDweu31cyw+f5Vu4llZTVjnJrjuSgTDTJ6CmNqE6Fjc5C
fXhtVSxWlHuIWG534EK0Cxe18PBmNA5gQCK0Ivl0ZGGaYi/Wo5mecE3GtrEIcwvq
z0nfB+/yWDcXVpKMewBWypXprfnuBQj3OSUJTZQkoRbvwR/+gL+vfG1ACjklcjS0
ZnugCM3UsBvsIYeaXHSp2nZQNLaVxyEH9l0OhElCHG7bUaz3EuyFBcS9IwYn9xLg
QJS+/zvR+LQ8c0d9Qjd+xra15w/HinyNOeEC6ieu/llPciQGSxi65MXcGfdjG3UT
H9xWKpBFH8whkgrMDqu5eJNQrTv5ltvtzW3Gx8uFlhcUDA1/GBC430MQOaH/PNw1
dRBKlJ2F81gxVIsR8SY0idw7jAGTPYsUmFxSyx6J7N4HM+WqcacNvJ2nkrFeG386
Qi+PzKSHpHClo3yFp2zMhPEZsKM78A22BPCQth+jlZq5SsxJWnxAnCUd2Go/hbWS
UGSIzJNogOgnonQM9YktAz/FFv5o7EYdIHW8RMbAhHk18l9eIcPQGZxZctMOEEzR
MQw2GW3Z2VbPaosaAG3ruF0upwxNQVd8ntOGjk/eXi4etvzESCpfy6qTmlqNAU1i
/q+KkSNHCwAojkYD8Fo+878+/KTruHywdG/eQ0pxiqZBB3ra1lfHm0Gb7aoBg8Uf
9jPEzSIWGcgOIgEKKg1DQVvN9gjxYqUx7GLoeFk6FIxNcffhg3pTp05moCLSIwe2
xgNO6IYWGyfkz+Bi8kAdaRIAqoK6sIZtKdjH7F4lJ3yqOHbL8/Rt+5jlgVMNrCJw
Uhu5eT/OCSjiybFOpWAuJtSPO+PafVrUE84I1VMRa4k8+3ctZk4Z2O4PQYwDTs0i
W02YXcnmU5ak7T66NyTW9p/yoYJ2kLg8cC8qqs+o5j/pK9WKaQeQXPj36WrdjIxN
DxUUi7PNBYWcetEIYfeckWyMYwC2mcEIOBn47bpZOt5kvCDQb8Swtj5bZr2mgCRK
eHH9BEPkCsHzQ57h7F0hlybY2FmMl28Uc9K5q+cbXO/3l8AcCZYR3xU3mVlnksgH
moVfa2vSVGrrNeIke/shbKOafAvCqrcb38xtzq2vb0vND+B86nwoZEyLmWz+OXGU
lLCBbl5UNz4Jr5lemS2p1X/g7BGsQI6CAbiTo75G90lJBQOirg9dSgixVjEtqyL1
pyhXlKb9jixJ0fajmvrixXbcJhezyGAr0ivCvuFcTsPMlKrZd/vFpczfWCcPVsN8
ZB+ldpW1/e4HZbO+4EbrX+a/DlhnCbo0eDHnWhAoh1zRJEgYSvpAUnjie8iPI4qp
BZDtQurpZ8vaPdo9EUD/6vEaIhenjQyrpiHHIdM5ZDBT6BWQQmmS3moSWhJLemTG
I8HWpLQ8Ih0xKsoqVd4xR6Ktbht1YbUh07eFV08n3ZjvoqUmSEjv9eJ9xpv5Bxp4
Z4gw3ALwNpLk3KSz43a6wYzqdcYQhVbTnUL37v7MDbgZ3BO+uB1VOqcDGFClEyHX
99NiLDY6+fLrySZhhT1QnmidYTqYegSUSyCWue4a1DY9FXEhwT5Xi4cTFoO6NTmE
bB6N7g2sLf29VSS56rDz+tFTcM2eTTKV7xWttqE6nUlT53RvAzJn9PurkbiAXOpU
Yzx39FNc9lgN/hdK20qew/aIv/6fpRfIJ7PzrKcOSnKjf1jkmuEhyBTI9QU6H+qC
6AS8oKoYz+6nQQ3luuXQgyA7KCtOAWfy86S6cyRJWjexMvAZKU6jhPDtnKx0ZBEQ
Ajbec/iEIMIz+rRy5rd82RFBUfdtQMq1CebhYfspcFbq2jS/VDeAX7H3rSdDMLAU
PXdY6+eXMZfLLQxdAp91oO5gf4tvXSu6AEwYyk8bVwmeuzNzigrN3KnVuYtt9EyM
39MZqfUiiR/Sfr2SDsct8w+b7bWZNwV9APTyvn7ALiQCQ5hVXyr8BnopHZNcWbWU
yKiVeI6E9/GxWTFDZJhJy4Mm6jZcZcg4IkPEeVno2fCJ07Paf3VIeULEnb2uzpfy
B09eV1tFTsoIYx+nrMy6X+PMhE9yXUbabxUZNZ9LP5eoVncq95h+wK1lXBVf1qSJ
TAHGvoOV1iuEJ1dnRmoouelbTxDiZebT77y4OGpH5tnBULER/1zMvcnte3UVgdwV
uIXNnpww392Eqd7wbelfIVyB/RtKGMYjSjZ+/xNd/d9vbBodVdQRGV/V4vllGOPG
Lxdqbgax4RsZT2oN5cw2l2C1BMrlY2LeZwsfsZaNIvDyaM7xKLawm1y6V7bkuC3S
yOaXE82tX1wZ9qYCW/jXPTFY6PUk35IXP0ps+y5ESKoifESaLdnucHSgj+bdOEoy
IqJCjmWcZLokamjSxhRlAZ/ZmCVNCNppeo+j41Fnf+JkJgDOycij3gQ+PtEUOpwb
rdlvCthXh9tU2lhWWSYhHqZmCJnhLAhhfWPUxVVzf4fvnHOIWNopTYH7LxEB47JK
0sWNyfBPqOQeVQKUwFZ7AiVus+F0RqzYjJxvem4w/5+fxej5gB6vre6ZFzI4pVkA
B3cckeCo9/tPbZ5T11cVkg29aWHw1T5GU34IgQdJWmouty2PRN1905+Xlq5rOWfH
cjoGQmnilZ7rXLulCbpcxYhYkaAQa9unfyaRkP4JlHJot28iiZwV7ZgdqcR7ewSP
BlPeVu+FvDN1G+tNqv2ZMUCLJtfV/jW5lO6V4gcOcjrVvLBGrA+OV9fapl56j6fZ
zWUlqKvN2c/0HLhjXGfSSvmz0aYPXiqoGt/NbW+ZqcbOsC9PmPI8eGi59mp2CywS
20G/ElvQF5lgHYrY0SaR4AyTS+n1vM3DoBj4t/W+v1aceDYUWtiywjEea9GHxs9B
nxsTtkFZ+fuF+NiFHcZTH2JcvLs0hAlOrM43/r9wlAJT+SnWB8ssHjXUe/8ISl2J
AB+uqPTWaHJQHhAbx/Z8dAi7jPh3jrRFdd7SEI7nUTlhtNq1I8BtDN9AkhaNo4UD
3oarypl7AI5wjdTNqdSczQlk2Iy6ltiJAzB93ZwHh4dCin/CrME4LQyczWoxLW+V
jCtb6agV/7BftU07b2c4/mhHPdCrvjwN6QhBUhRyQ70ihiYzKXXSuKk5oGCR85kK
ri9cDj7yVYexFugzdlMTtGL7XEs8H5CgbzYy6cnffQ7KGFQvZWTRo4fmPDOOaadd
SidHB6ZdgbFpEscl6Ny9Gi4cNBomJ+epoMZts9f0os/vp0VPKwsdZB4/o4pkMV73
+/k7WU+O33d8SXK4+RVZ8vK0TW6J4dr8Tg8OcrnqtL62u+By5ZHTq02m6AebwNUq
axtJHIy/TW+hm/yA+rgg+p8EW9buBqYycchr4mMn6dHv363vK7JvyxgCGgzqpx+c
veH9+vnehvEbzAnhKtRe4UotGwnn4TujpPU4Sn0wDX801Ef2mIoOFPmjC6d4YA5Y
zLTGyJxb3OzewgLxPN67IGE9E8DiTPQAHECLdo1TybpdUlOUXSyV6rvHzWZL0E8U
mroLu+KYSeY0IXWgws44Odt8nNa/YLKVlUzPTtilsyvSa424NZYcfnUJ0wE1bkKB
AlPFGM7t89WQs+SrHzRn2SANk8m/dUDZ17QE1V0hrL69OAXvu44m+QAqqBmkenQN
3HI9sj2lwelNOXMAQPfeX2SB168KEcDvEIb/7sN/BbtuE+9xC2uUSJIYOW66ShtQ
Hvw/749gXBqKq1FR6bertdbAGNse8eR/jYHXy4LSmU6Xlf8sM1eqTYNLEAPeXJkN
Fq+tPFH34KdOrKS46puPPmx6ynfke8PEMQcj8QOcEJNHmpwJk9BzSlPOzoWt9iho
JwrO6Rrwjb3nPK2RqGT687eVAuatlPswttjFVxdEhAwqlq7nY4kdjph8/JORNDO1
VBBLsqHu+Vu+vKeAVp5suueuUuYAdNr1DM9FWxEncMDVT5MUilh2C3S6YV+Dkav7
8fjB1RvGOajN8ipdG8okIkIPoImVVatOCQnJKYm9oMbFy46D/lbP8OAyGU5lP5Dr
XQiUu4O9VmgGTDPRytafiKYwv5S9Uj/eDRFxtGzbIYtq8HU19Q609VpjwZ5IGLsd
VROJleI7Zyo7yRKEFGthHSKdC9jxNhqV5YhnVERGdc+bSSsSzZkAgleOmKMx4kqK
nu2BTKP1WIsc/d7EtFNfrN6eULAewykICAQUIxTu6vitaqKukvqowoQFObpkZ1ZA
wJyWgntiiyf5jR+lPFdJwZhjAom9UlssvMRKxZhnRKZ0Dfel4cA+JRXm7FbwYZRx
ws2CcUKx6QSRn4fwu1fwwDoL8nhu8qNrE/CvYFNpmLbD/oM0xBVuCJlPiRfBhB9t
/xQTEKEZNq2mk7HWYtK6fDlUx4cTHmOsI+glvAz0Ykofo/bw/wd0JLW6FM9WYI6E
0ucsgi8TY0VHlL6aWthe4r9JIWLGDCaGYzEXgu+IJU8BEvJwRBJZLxj91vXSxaO5
aJQzB04bktrxIfoE7ZCiICq1IpnDlbuDBUvl3701p5XPvYjG5Yw7++l7lvvetvTN
uqh+sClx5u59n+NIM0oVYTIrJOPT5TR9bEj/6TiahgLT6JKtmr37Le0tvqRHn2nC
b5AcX0xVDXk+tOfQOoJunM66J79hbOPCrg336iwmf/ng6ckmeYfoOqrZ1L6yupP1
lEY13fFBpT6fkmM35vomdNS5yc81hK155h+z9Vz9Y66cMdS9dDEWXY9R472Djt3s
W2xXa9n+1aPhoVxvpJa7aTn962X6W18KQqpr0oAo4WgqyYguEyC7pfYrb9QbDup0
M55p8qEYTGGh5eAU6PK6bpug3WPGtzOtZX24K7oHbrEo1azyoDWB3tdG7+MJhjMM
qRotkDx6dtYsl8q4vi58NRdexDJxZT+M5VKV/n0XoPS9HOaCcVxIZj3G0j6m6QK+
R9LyPqU8gmi5dC3/CLzW3KfkgrkdA2bWRKCzOtygBlmdLNm9+6bwOK53zkp3+3YC
rwMcJa1AonIlnZKHAXDaiUi/OXDn9pWw6wOm2a5XnP2u8Ut6n1jBLxsT4vDa5W6D
LjMMfbSDNszSzhxKtG7LN86IQMFof6yRZ6wckQvkIY9YLdvTC8rgIYuiC6bN/Vqg
X190dj9iBDS/RHNuMWAodMmtFtw1BwAZrbvuh+y/NhCDaB6TZPfW5l5WRqPfhGRO
OOp9Wty9cZJcAO7y07MUDLWVdxmhi/XgL+PL5DR3cTX1lkWS8NU39eDpJHjasz4p
4gR025lxz643sbTnoz+mw62r8nIiJPc64OJGw1b2CJtED+F2LV8Y2lxgFt6+tr0t
vwZVqTGyeGFi1BT1XlccLia7ryC4+7N6hqLM3d3LvbI5g7qI4V4snWM0uRjCPR2J
bSi/gRzl1FJyMh2AHMMw8nnjIN/ml4oMw1jRddd1KAEC4PMhahFeAb5rp4Yw4O6A
BlNLU73KVJXvNx2sMhD62GsFnAI8G0wWZqAdoCrXJCSMZ9A910FZTvFoTG1hnEFW
9ukgANepFZAscVqiVabzXp/S3f4iFnMsoznumV5L6dpaqRjB49T+hye+dT6poPW3
Z84nT7u/xk3w9Pi8jjOEgQVcyuxBKB6Geb5cAUqzdBZYqGYxdqPPnjOMTm8T+nXR
BWYu7tfoLGOxPJdQkiDehjFpHx8ojzLD6AtIciiCaIuVDw/iu5tfukn8CHH7AW81
Z1iAc5QpTlpTUOOfx7htPEtRl5Kl2hxNFZIh32AeeYXiEI0oZOS7S4+eTKr4poFE
geor83ith+JszT/l272HpwsrVtLkJ56ypXeJZ9t5xhhAO4Vpc37f6s2Lr4CuPrRC
cibi3xkUhi+XVp1YFl5M4bJoLaIsEG8JV/ocPLFsfWyoP5ddHy+Z+ZlviyLuqms4
vKz+48jtcxxvpdv+wM5C1K3Vx5s60/DqPnn5rNYFFC/mTuwyj8gUfnt2lmQ9gtR2
uiH57NiPhkfMEgXOg1oBjPi3QhjFfvspeNX19xDuQPBI/1XFYDtJHkJtP/8wY6nT
4DsKb19HiB5Z9sPBmO9++pXYSx+3ygFPfWXRe6p5rJXGvuNysWpBXWUfgdSq3Oix
2x3L04C2EaGWz0et8e4C95sZ5tafwaylIIqb6BGVlXfG/RdlneNadgI3BMrkEOk2
Ey/+YsaLtt4z1W3dexJcBLTF2jGP3ue5OlJxVLcLDeL3LHWTIENe3V5rxZEyN5Mg
7V2uVmsn5FQvCcqyLftCyT/F/wtNYiAC3jIJoGDeEu8g5OcR9cmbPEUjD8QGrfjO
JQbh0gULa9kzrkgKDons2LBq5+7Xwex8XbVsKCqWdzEXXxTChqQAtNwqFA1qIZfo
AtYmdijSOLV3T9pJBDfdmRSA7ny3jSPaTeGTSM9NcHtGUidaC62zPLQ6YuYtzBOm
LpYr+YzyOKQUo/GTYRctScC34A57TGwbsGxUZmDIJf7vqUQulVbbKKfP0Ht9X+2p
f1mtKURwWf178b60XPiNXfkHAEuQ37ha+dq3j+uVFUrg4oxNfxDHE3ofBhM5oyNm
j1BtvDqnBHzQbposmQsNEfFRnqbOfRORQUfD7ZMQavlh235a9OUs2t5Q4sIvuuRp
3OFhPCa4cSg9PLzVzYwxfThhE4VnycXJn98uiXrh/duzUWxkCc//Uz+Pi+UsK7nk
JIUKvNEQPzT6AC5RfSzq3XM8vZzOZ3v+gW7/McFBEJA5CiyD1D82x7+F/TVToLsS
9kSvmIbAuRGUVbkUs6qKOX5CCLezxUXKufWzOrFf/bgpavem6ldsmPDOE+Yo16Me
rLY9YL3ENCdkO/G00afBV+7Nzz65eOLY5AzH2exI/1kt7m+4hXErEoGqOsfTEmTK
LqVIN3TYrV/K+3/gp8nRxjqipTrJ+B9/xVVS4wn+3tSuzU50lyiKIy3ia65XDTZQ
jppWhCrYg+ES0dDr3/+PqXOhlPa89f8zSQ8KffCHj+9z9xtzIIVqXwEPzV4rk0X2
eC93cb2IMIMD5/sXCT6ZUAGwLeVp5qkemgd/9eL4Q/lUbckczUulpFaHTrnNsNb0
nY2s+Cyp+f0bWsAc0YyVrWMcdypp5YSmzPAA6z4CiiXBxETp4sUCWvHZF4nhwXvd
fJOEISzhskOFNlOOoFBsDekZ5F6sxArE/JLh7Cwj4hPcFsJwf1gKQ7Xf2+gl0sqY
U/yucflI+GynQx4C7RzYj6hvur/1PXZqcvD+AZjpu6LHwswk5zV2+VHkDhz9cUTT
nAKRjrncPcP4u6rZB4ixx7w5tCl+iXDncKi3FrKfrFMq7Zbln5H7RgZ5tFfogRtv
Fe37khvtJ9JAFH0u5RHI5Qjf+s4gU5SKlh6k5aVP3VR9HvMKf8trY1o3NdyevLMP
7wgaHzizhmvehyXtMyUhJLIlfSmAFC1/zMC5zQsljABIr3uNH5XUaWH9PrBiELoK
kWM/V+6qEQhd+PsidKHhO9VOEPAR8jVsAow71Zn6uDOt7CAtAzMm1zyF+yOtTBP2
r++SPAEm7eTfV2yoPQRv7pi/1ablZ++SJEZIQkxCr4ASwpbp+F/yHKKm4QtsKZGV
IuT9pJg138m0talnJrpQjg5RXWM0hPJiUtbqgVy61KVZn+IfYv2VvIM4xj/Gvihb
Fz7rxw4SuVQLbV9SpLkMmpbeQGNao5Z8muu56orYyLEzGuU4dKf0Q2Uvgx1k+uhi
+HyB5N4dtuKWlEhmAmb0/XP3rtK8IJ2VTeUkp16zru/e7YcPRzPeDHen3VzWWXQ2
ALaTyqZK5gJaJEko+J5uvZHeuhQASRZ/dV7kY32b6d5C22VjJdolmcstS9wYyBUO
d1SrsGItRMukRsXuBsiVgozbJ2owBvFl4uTiBJA/laTe45knjJDRyOmuAxIZ87LM
TlatB+kaoqcAkHeAPjtwuTJHsEwUVat4QNrxoyTY5Ee4TnJ8kiS4uJuNZidk64B3
IvCRwCgC2P45fwuo72XPbSEvQYG9+an1jMWB5CBmVsrDOvRHrvgpqV+Q4m7fSbQi
E+cM2Il10OPSjoyJ0HgPW3KFyGAW91K85PUBl8tvpCXj7v9SdM9LbcdrBocmGPI0
t1lxJD0aYX+RJUbrAO9+CnCaHp02O8O3ZwIGtm3cCLZcKVuv4QY9cqGJfjJfVgir
6FPyQhCjee3b2uKGbAiijXv0TXcrPR4VdUciYeEO74qD0gpEXeD5YJ/CwddMoMiD
9P4uV4GcsFpMdCLJ4Jk3ZZJLukwJAn9CMKcYbvmerkBAkl4Gx6nPMAQ3elWjFwYA
UamheJsAlncmiYUun48fYdxDqFklO4Dfj7FOvqJvZFxZNkNbRksdRF4QVkVIsRzt
DEVTJ4DX2/POR262jZmsvl8fcbmuw35CMnqBzFpMkV0VJQTuSI8etaNQRIFUgyX6
UArYDNOCPvow0TpgMeAunnUZ+Tw42vGaRkP8EMSVx9F4emQ3PeEbJ6EGgrjZ+xET
2Mu5PMFtMlWAJ3ib84DEA5BiVOvyxERxAcLeOPC8nmoXoWCBrbkukUvxMKmDuUKJ
RlkmL66KdxCH8i6M2mjlk4/8k+Npc2kQTXNowUKfSBTfDmUtUFSwoaAqGn2zz6eC
FnvZPOGcUajD+o8g6Bkm5zn57CS1Hae4i8eONguZ8lR0OZ4yuczXQGhod9jHa5sU
XtC4bDpGAt+Edis3sM6Az9elPpeLp/8g0VML5tCdcihY/Z1QCqPM7Oi40t3ueqIW
n0rlMLDCb6fKhzccdcK/ARkacj3fUgLRtaUdufTnLbm1k1gjFgN403kxBdW++JpI
pCN0NV/fsIaoHzidf4GDbffjOXHVf2DAlMkNwNpBIhQyvQXXEIEay54Ytqz7Cesp
iVu34q7t6kHPLMIbZ2yOntZolrEn0smY4433AQgfNcEsNWibzNDIyEYCeAd5rnQt
4rMDWH+FhD7gt9J158G+RBXB/s4wlE19QmizXl7DE+D0XDujYr+MVAoN6rc96y7c
Wt6Zem5YVJ6mc1fABmNjW3JCkzuWAlDZ2L7YuEJc9dJopWb6hIJfOFfS/ut2gyPv
KS8AFh9ATNgavzIg/mFjymkaODlj/wRP4MlvlKMZQfkcoWaBH0IooGCnEx1T5agZ
tYLzw1qwJ1h/0NaWjHO+PjNTX2zDoy3btELPT01YlxdohV9gEZ86GWhlcUPG7pBR
Lsx4S7HhzOnR2CoCVb1gPsaapFzyh8q11xeA0HRqTIpKiXx2TytVKTknVRDEoqUn
winrtjM/9+8/2Xlv8ZOh6jfWMjuhGW3XEHSatg2FfGJ+q6rigPg9hvEJ4bZ0oRq/
MJtV+E1bDZNavSVh+7Irs9Q27d9giuSq7zd1N4sKEWDq3BtS2sqh9mKfjfNblrcg
DuVOUYiWS2r/NwZKibuSyPtt7JgrVa2LlYwCA92lVkF5014MzF9s5WZe/fjjbDr5
RVQjxsMpuwWo5Cop16el91EI/GY6hweedJKctFUtqq/ket6y1AGB6gB6TS7M4k8f
P9XWHTmMeP3wk23fyDeXey57YSuvlagA6QXWmT1iyPTGR9EQ5BufPt7ZphDYaEyU
QOVFpHA2KGd92SzyRrusJOkx+2PB+Cmxieb+rYupu4fQWGT9cQItPwam595EtuXN
zV3X2avHXk5rDR+Y/FaQhJcYEN69eT/J+foV7Egsl9tioe6dQvd5jpVwsan0nIPM
NFz4eh1yUGf6u5gXjo8gukCBIVSU1WfMDj6TtCFryQBKOQUj9QLJhzwUGE9cl/cw
LwAZzzmWS0CM31RmyR3KWIwZKGDv5fwHR0R5o2rUEqBwUVnQIISQNhqxnS2MfMQa
TqvvIT7besi7OacATzIFrWCJ/XFC//LzEwxYDPHnYdLktZTVgayCSyQ2W3P0gzJ5
W46BiLZ2IooK7KhBlbhHxMAPXbD291z9BmlI3CSjYs4CL4wIL8J7tdpa+58OGKUJ
0m31pKNizh5Wyzy/xNf582Wn/bHnKXvWlFiy303bTaXoMiSXm+oQh+/RZghTpjOC
xtKDgSn6RZB7eEWosG4kNhnJfP108ZG1r1jzbx7H8iQIJmHmeMgH/6AZ/HDkV8I+
EnpY213nIGoI6vv4Ms/jmJoMBbb6Ow0OnYoj49UkTFjVZXBE7lUT3/1FYmY65y38
nGy861ldFOBQtQRL+7+BtMpCs6pkdKiDv4G6Mwnu3VmQtZJvkCc/HrHgwnZwliId
q/HzdLAhjTlBE5G+U+feTM8LH2sHC5qBAL6+aZZxYzwSgaOycH0boxToHpfChqPV
hkMhnHhAbraVh2ApUNtsXSLcQzejeKJchfLAWoxjubcOGnzAyVnmbB9ACMHGmLCa
+zKg8ohXx6WBgO0rzw447R3YoVQUbWc0nKVOB4tu/IPLktq2ffIujtWvMJJjT83N
BSWI87RnsEilUAO0suRYyrIzvz2WV+YMtx/y8tWo4zuRAFbLkXDl/0HSsSyU+ZJN
BjU7ssQszrG0nKcI44furg4M608ip6UHLutvruJy+T9yaG6SwVILincwawms/3qq
QBLj1C0/dMlQQ10kDdpyfRZNiPOWAkYhkAkg8ehqL0KkwaTq83IrNmbgy+7YPCls
46wW/MACmD1ys+2cSUaV6wczdZg1cLdxszEvOSZ7GkGmw94/R1pykQwikYGNqYOd
FFtxYLmlhpuGL8PgFvFWPIrXHoNWzUOVdg3xqZzeNDteORbdllPW9bs8W81QwaOz
yT/WamZvhXHCtzNu/pUbEzdPpiNzu+CLyegl4K6MNVmbcIf3h/kUoSkI6jXemqXg
tX2lcsvnsy+EAJhjKdZR+y6rEfYAODb6kv+Ez1cNfjVFKznymaFd/lhuv3w8LmN2
tTeUVw/YxZpomFJ66cC/Ta2bgnLNhCvULkQMn8MsE89FtC9QlUYXwW0/nZZYoJMR
RJjdQu15R5cBnqljrmfAYKCAkmA6EZmG+fCgVW9nAszP3v4Krux1bXWsLtA3JrGD
dX3HHFsef0gd583cE1aVBfrlzL7Z1IprCJV+z+RbFCo7RJbuoFBXR5b+3BYlADT2
laNASxOIhS0WrnhxYHpBQ3gAP485A/pllziXvAHqcQKoG38CGWfDh1ptSAwXqyqt
/PpujLdtRAKSlK+m1sBVPkZ4xGVoOPnyUAekdxWrHcslcE0Srjypm4ndtbyLT4XM
4Ej9adx1zgUx8tpI/L/UJv5pA2z7KnRSmAr//vY60NL+QZiNxdIFjzKP4JrE5lhi
xxjM0uZdEDFE8tc5PmufUfxL5PhyrsHGnr0n5EZuxolFpCgv9LSpu0buuJfxaAXY
ID2l2UtqXWU+WJTWIw+qMm103OTX49GvnY7SQ5ChTS00oJP1aopfAlzI8B5BdeW1
nbjEGpzrUBHaRrBt5ennobPiW+TgANV7p1aPg4yDsHZ1800x0EGfWA+rTBRwmRVc
rW5WmxwofxOsrc5qPw4MuINhU8/fmQx8pbYMXbHUjhOI/mM2J56bNwtHY6DQt3AY
eYnkRD9hS499x3RrtZlQnVhClZveXHeRc/WbuGjxMbR3WSIV7KQGvSG4f+j05AVT
nOxA22Np0tOV2oVzPN36A3QfEXLFVMAqG2Vq5cvNrivgPzHJBF0J7Zij+he8r39x
31dqwnV0vV+yR0OpgmTGioVYye06ObQgERq32Nu57K64HloLIWGK0k2pB4hitUEt
lv9P5xJMQI/h9eeEvTX1I2ICr9YbLQXV98TyzIMuhJrhEz12wpCn41nw46hoHucl
Y1ZbFRdhefZsQ7FttSPeXAYQszGmbX34YQ9MFrrbdRp04Jdg88tnLZffwwglxGZa
i/RVJP6BPvwPmxtDVculwjaeTzjFtj00F9PJ9ILiyPutEUoV6JZLhP/iT1dvAzXl
JkcDN/9HaSmNAjamh+uqIMFurnexuFkjzix9LcJXrAKNwHDaeGx+QbW6PXfvhzyQ
26zxsYIdda9Z2/7E35dAXSwM9L2GwbbIW/Fu9ErwzIEIqysxt8FSHp8NHrh3JuY0
yqbAJhI/mLIuqxcDvRvD3EdtVKVtDCWGaik6hnBQT9RHwiBkLWgZZhyXm5Eq4+ah
j1fHm8SkUPJtv8kMLml6Zy+XYcl/y47FZGmcH6IUzGOWwNCcYusymf6Ram0Y15pB
bf0MRKH068OJsGfvHn/BfiSRGmrvEwHWZACn8+hNAC6n4VcNAXXeTIbUEE0vTPl1
rVUa+4rxVD56/rytZhiysQJdylgNNXGKYj2NmCQBgxgFtYio9YBZ+e9KC2859Qf7
cu2ohs9sqF4Q+YyQbpyfIuWYd8CWg9XkFNUjScJMrXVwea1g6YSjUzeLm0TlQ3AN
mLC4n5ryvRSosyc8byudLoBr98cu3M5etl/+S4cqMkm5S3lB6rcjhD56bSdDTNGw
xT+d0MA6SDoSE61kzXGOvqvJ6+Q3borgz3JXR0tm9EJgP/c1zJYYODp1D/GqZAsn
BUhIUJxhnhcrRIrYmKn7XTCu3QeWtYFxBIczy2uDlvbP5pwg89Wxq0RA2wWn8hCK
Kuu3e7YOmdsItJ9EMpeUn3FOfj/4Os3cgCJTH10fsaWlGfXkPcMhKi2T+skg9X2B
mVT8xhD5FJDucOOMoJgvzbfKwxJ1qEiXP0EOcJcRq0UnaPrPo7ymUMlMzCAtoRS6
Ck1ImKuWmxlTJe5KHPI6C8FnVxSFf2/x7Ya4PyvyiXiZ0FIOair0YT0qME0ePYwu
+M2EcjpfyegVPbpIhdTwiat1HRt6IhyT6PawSUks7kidYHX4fZ57b9OV/xaEiJVm
OglJklWUI7BizNY4+YZaT5R+8ISwil7M+J1FKGKUFMcuBjZQ9lkZv3n2fKpLAynJ
FJEbI+paOuSae1ZhBEQA3oOaY+9IccqhRJuGOpC3z8CqjNvvd8rIxosfXMMyLIAX
metzoDdionutaXFaYJ9uwV5GxGHyKC6U5fg2FATCtyLBHgcuuaQyLtRtwvoof2mj
9XDfs8Syx13EOO4DLpMg7uyAhmvoI/DBwUSxas7rDyupxDadWBVwLtLNvW8IbrzG
VJykMaHxUGLezjW7JF4N+rIORC2u6O/91mZEu1LMHprdGa91douxXl3ceszE14tK
6nhL4D3MzyR6E7KbdHv119Z8vPYaWUeDIKDIGgp1d20gmBwJssPR8kZYagGHc6jb
aeZG9Sy8fbbathiEUzxNd4VrQULKe/H7DhpVL5cyk0vf2vU8UZCkgN7lUcrIcL8G
rgp/sg+UGzOydgM4enTLVsot8r9KQjn22k8Tg3ERJTBJ4A/fte0fY7x3JY5sbCTY
/wZvBUdL0qmjmliZyUy59wdtHH/avr3h8xGIsKSjZNf7KbCV5NYqUp2UID9gYB9g
Pv4lxj2097yvwL8efEMZNhBXzja+OY0TBgkrHSL76WAlVESVTcxHliu+zcctUq5p
AsMJL0BZ2MVbiG4gaYHgQhW1gt6TYhXeBQ+eaDvYcKCZJaKrnV0VfeSXBzwsEFEq
Zi88ZIbW8ywT9zGGDDU7Icqt/5b3je+nhNT1GCctp7YGyMtEO88yuXIGHOJ7Xq6o
WtzcDoWfJSpjV5vbHcsZ34mcyolp49eeXUWV/OLr7HPh47bLG4/dsQhhFyQNHZu1
OF7/jXOSfeBMIJEzm+tDKjvNGVQRRbLYlGpMIWtJhi+h10S/QOm03Mx1oXqQjvgn
DxwP1eRhDPuEevB6BtrIGDtQo90dDCdDZFSuYdrAnxZc/1bfX7q7H1c2IC3qg470
SnUaqeQ3PUX36WNPE0ftV6IvZMSsLqJBePqGiHcxxDsgvzFogyQWmBFDJsaFbIbK
S8EUdmMq6JuCGzZpaYKqYINtpRaAoaVVo3Ol0xTmWLj3T1AKRhKWiuvk6ADBCdBF
cFoXlWl+6/9JAOIUX2Wv9oRFfPCvaEpmOF7FM9J9qx2/evnLjgD+Wywt7dXM9aMS
ofyDH80G5YmDyYrvBGKsC5yzRLsg8jPq03qLTYibbLxoZJA+bK58dm+Y+ZTORKN2
eUw7HH/oKzlPBkU0fcBAC8vMnRBM8aIQBRTamnhggO1o8ryRJz/nOZyFXwRFGTz3
txKcIRzlXE76ps4nUBHZFIOPwhsFklcfihbShXngOb6AJHj8X0sI1c8yC9JOmgJ8
FVLgcXoHbYYXa3KMc6jaoXRG+TXsBc1fXs1d9EpWBdl3qYZRmAO8ZBGiL2zL6ZeV
IRo4TubZm0/F4xM3Xtizl2I3oHM4RRXJvJzZrcWx4uES60N2jh90YPfUAAacl+Dq
dgtK5V39O3Yljr1AqI7huJ+FYzFURuEEVHKmlAkfgrxWI2qHjPdwVWorhtSRVEpF
+6Abb4lbuFff05oXwYg1p3E79bBRo+q2HC9Zmf9Grl+A8jFB7vMnCr70hGOZ7OPn
HraktUQbefUQhdeQBe+l8LctcjZSd6994hvNoGohvf3xOp2JN1Ufc9wGKPTEIlY5
Nrb8KbuBYEUSCFoOyzhrlNMSc1+vLELUaLaagcwzBOQCuTD8oVUGpVTjLVAN0Jjv
1CtmvMCO7r7w7SultPxgoUQokB7MJG+i1iRjeq0y77cDMAzaq6coOsmwEdW1Wac4
aenlwoUDAkDZoZTKjFrb4Rd0Y3/Kq+NpQLzU8y+WLUHDEmODD70uQdXi/JNyVSbZ
HUR+eozkQCvH2VI4jimcjCZPFU1aNBuadduZFNFGzgtya2MJYyEkalhYAe4vzhwL
be4Jpwj5QgVVGebF7xK2TrgOiRPV7yKdCNgFVID1HYVfGEZ5u/cKbdxXVGCF61gB
yEdmle7k8zVvlVvG2Ytq0eXwF48//u6bdejiAZyGcbxEdMiK0j7SGO42d7pyEkDD
s9E30cINvP5qtqS+PiqmvGW6ZD/oNk3FQiL3BatsLLMpVvzkzKGNJJ/qpBT7dZzU
8X4g97/Jk4lp5PIXJMi5wCbYIgPXACUg0NWLczdli76HUYd+RAgvM52dd0ijJ7P2
e62ZKW3gsukbrmuf3iZvKlRsJIpb4hy03/rCbmSMnzWwspF+QtLcDS0aAwO9TAMU
poDgNce94sozU03T7VStRXnpubiJDW3m5mr0Tlev71Z2d0s7hdJe+GJvpYPV2ISV
McbF/AhtqYP+10fhWiH4q9WNe6PVc6U7zI18IJX/7IgKrr6aYZMb6pLkYFk03idx
FgLOX91/451eQ+VypXJazsfJ1O61osyo9rOw5MN9Rf3pN3JQE2XnZHp7xEiw91vQ
43juijweqtFAlRnO/QPX0uDhtu+3AeHlUH/nCxdoSZ1HHtYYIUpOByVnRYPu9TUn
PUm0xjjarP5r2TaA98XJXRsd3w8K/G8UPG0tbhDZG7whWIS8GK7WB8G+pw6NmMgl
WuvqHzfvvA6S0j2M2q5/RYS/T5O2LxunlGYG8z9Si8uS3FlVG8YPATqstB5mu6/X
/EcXcrN3QhD+2GnrJO0jn0CXXwNWqcNlTxmCXph/TAHA9Y4CTRpIvkLn+7SMUO5f
U9jiXYJqwzGfAuhz6izG0wmWEpqItQGlPx7fk0Gj5+7cOp5ogaWcETt2bNnvo7vd
yCnf61k7mWth7A8c4OprSv5/m+VjM6RAf23O1W9Dvvyx/O7nc2ZLihCDmel/E8VD
NNE4eBy8OKfOOmAET+zPbgTE+fcub3AWglSI4L301cElnsYVeO51X3OkaBd5zMtW
BTKuvsmaiaP5u87r3Zzs8LNlG4M974tGlfF89Yllb/IxA8aHKLMYgElW9ulnXzSR
VV/iUp/WjuVKJOW/joqviyvO5UGL4sfHOPPNEE5VkSlZbPMLBfqTTJcbjQczoQx9
19YFkGVTI7REJMKBMxlYEjFTym+nVAqC9NRXCH2Xmx2JeWUyrxEu1kre/2+rZNmI
Co2KpMVmn+b1HdRVYpZqAcWyJJL6QPJT+bIEhV5cpOHCMFKCoaqG2dSQm27ZIOIo
4PN8nwA83ryaskfigoLYzS7LQKsiU2uvIg55L4AzD2Elw0Vq3aZ10+Onf8Df+6XG
WfGhBBL3KZ2nBEO67BfUzzt/vPjF7kykZF16bfhKrICllhDTADJNaOaZT/8u+ESR
CNs62n0Y4F7seu8SVBepPfgYhKfcGLnazlTKj5VNTDGvF0l+5p+3ix1R67aM83sQ
c2gBuAsCILl9mpvywvhnIzrAoOmBcG3YaxJpkrlzMH74QdpHbJSGCfund9yb2wOn
ltMIn7ceMkAlhAdnMvKswCDbQ4v9Y/B7U15R2P5WCFcku/vmuMevuqbztASXAhqB
mLAWskgzZ6yqxctnCDBVTBquP8bAZuYz8NJA1eSpYyBhRWTlKaJzfrGMWZuawcOV
am4SzKPjZCPVgfzGnFXUPYj7hS7yUpPplB7IF12c7Sn3YjSsk1ompv466e6KTZpl
3Z5eJL39Dio1ceDmDIu+0VyZoeV9TDrPAmNE4m6RWeDXxE3blPDx4Tu3OlrHZigg
UN01PAxsOLmbrTrzGPG5wpSqA0FVvyLIViBzDp3C1VOBZdkA9oEqu4md4xxLo4ue
Pa/zkbnsl40rvaZf6RvGfYXCuinGNr9KcqfJxvV7u+47ftrNQOCerkB0dZ2KKozk
jJnFXZW2xV9Hz/kwAgVRleRRGBNfY9nWB9UJTPeYAeex5bZKVEQu8XqdG2wQEhkP
tjDlHdbfEI0wEUSIFxDx7sYp2mWX3sDjSq4LNpKojd4QUO9UqCiKBAw2epjqI67L
7yLZpLqeDg1FeQtiZhtuEZ5FPhUUGnj0W6zvJGi3GynYVUw7YpbUOYT+nARyzfQ9
3ZMlWF4ZNGYZuKNb//8UeZpsVeuhh461bdXKyh0eBK3VHijiLUWi5556OoedfZal
W91XSIJjqG2+gl00FVxXy+wws7n2l1rRk5sSoxBbU6aizK6i64IeYoZfyyFCylaS
axAz/Afk1NKgB7/37QTOiZeex3/ZTw+ukJv9YukvdehDQ0H3vfgwUE/xvoZy9HEH
xGdDqJ4ka8UXu2LzVoyrNZrP+T/MFyopQYfWMtNQKOzh48bQJYdKdFAjGSrXaEKH
lJgakYku0YoiCQC0MF/hV9kuztH3XNJM8iIQqCQmyZATrL3eaoHj9W2TEDu1cnmg
zb23KuGNbKQo1Tl6V8HmL6YemiT5BLp4DTKfsDpt3M67MOWi+2zRp0zGGxPAyj42
FX7SfH6gMv3XTGiM2Dse3jCY8uXvr5djXf5RxrNewp5nibSSUeE4eGQJpUDvY89w
6ZJ8r/r8GgvUyk5QefEpgRjTTMY0UT1WXcidEsU5HfZsL3peQ97NQU9N8bHebcU4
p4mmgZ3rGwTNJwe09GeV43yj1zifXVHph9MlNmhmBwbHUXI4ONkNHQIlOLqa8gCe
kCGz/ACufhYChx4yXZdfx5GOiRtbNdS3/lOzUQkfEJXf/HoHCpLLNdGnXOQfGy4I
8Du354z3QpN1KL4ZBWUba+KtWngH2yxqLItdp1dN7YV+EqiOXGVvXSU0Q9IYwK+z
FgOrNiE1apQI4kcZWHt6qm9pCNUo/bKtxHF9CYAy5MrR+hPdQ8YqpC5bog0h9P72
8rWX/bYaqvUK5SOyIOQ8uwnSvOG5neoYNlZXZzS0MHh7cqq9+XDvXtAsvvq0mWpv
5i8gKAGFo9I4eieYrZ+UeD+6+XTwfthrVz0kB12aOmkDgL95czwH6kc/OWwQ64i6
nCZyqA/4m4d7Qd1DOED+e7+SMHurhA8LsbWz5BbXioq7CqjbYStYy0kVxXFbJJA0
kXFmRBucfVpob8SroBDzDSC/NAFxSW1mjT/GreHGzwkc+d05qgxvb6wpfl3sTDHp
2En5F0JT+jZV4GMj7PwF/p2SIPyQOii2LSzH0X1k+qTpuoJwIRHxzkilXmch4P4x
EX7sNX05sAuS6WfQtUvhIUfl5wUkUkDHZUA4eqNy2i0LPBHcMv+umVVTiS3Zwq+d
yZFWuqaI+kg31l9/0UB25qEkb//DMMC26b/tLblM/iK60XdezZz96xgUlW9kFwoi
oPniweAFcpwMBd53OpFYKdOe3WZfXwR28UPM6H0PrmdYYqsZb0F2GH57HW9eCkb3
0CyI8XxKKTtUQWnVi9CV+WhjZMPwGn/TcdzR9bNX65XsKks8R2L0cuwsGwc0M8EA
NmV2DKbdd45C8Sw+/g1WIWwRzsDSsl5cdDyLrO7MATAjEeq2dADXLwsH0vNlWaC0
+3Mw+0xEqQD0H33untjYeLQqa0t54SMMeDooViAShnX59K+UUeG5n638+DCSbZvG
5TvFjEL2ea3+UUGBoxizg1zF5LjvPVE6FxS2NdqSt7bre1E6CqauAx6QXF/1XBXd
Dsss7g/0fOHEzoUGzRST+k2liBWfbt/EEsh9hDLZt2pkkS0Is914CDgClNGRpurR
Yf8oZAc1op5wUkKVJPAjwDOm7wwOTUc2IMDNhUybG3hFuUTCDUNmFNLv61ackn+/
s3ax5I/dIwlDwF4/AAJ/gUe+Amxq1o0ZpFhjOFWoOD90ryC6IO84j1eUQDBRWHxv
to38QJLY4S9aVMl33dVWSHI153i/DmPMCQBp1dw+o8JaAxxjwtvU34gKBJvUMDXr
9/obFqjhwIV8ZQctOyVhIVaL1q30r/4cI7NDDGLzHOY2SxZIg5ySrNyxefuUHB6K
eEAFRtBmZuoOYy1EiwzNDNUPIgzMzI0wzdz7LVaZwggt/38WwHuq+iM1p5GacP9z
Nhk4Fl0tUbmZh5M1wEViOzshWfBgDZ9KQ3c1ePZLaYM2EUU07Xo5r0dRi3/dp4ZT
gwCm1Wr8/bFABgCIjJKlwR2p836MCfE8XJzgmKaZ9SRgXTYC3HUUtpZU5LGiT7oh
kysFXVoccZDuWQSw5rKNwXiB/7Wp9MCU2vX0Zq2IELMyY2ThLDKbXL8gRimc3Hyb
+DQx/OMCtPc34SUzsUHDA4VKoCt9xncrkGPQh3OmBq6PJX6ATo7RpMlf+UNUfp0c
PF3DNrxPsjrGCb8Exu0c74W97L+G4E9w3M1fvhERzgt8FFX35GLYrNRYIwMqTjec
VTAY3Dpcit9dJiPL8rxBQ5yQ/c/7H4AjF6AqkVTAtjnX2wduB72mXq5jnnBfQ2U0
E8/CXSRpxXyVfkJie9Nrt+wS52UXqCZyGb+yRydmlzeGTD9GbSjqAXEm5LaZ3rYS
QL6I1/+K5CFLRO9cEXqHGPYR8MrRnV8eNM36zGOA2eDvYZhcjgaFbQiUCBuoXE0G
LPB7qwo5ctXVKrtqTwRMgXs4sLjkkG/Q9UlqxXjn/4tmjNftQrICC0D0zgAJGeap
fXWG/rYRGvnUUZ84yEm26zUhjMXbz4vJzUibq/T+hmkRU2BIJgH5+xmxTZ2Q4liN
8uhCh9PjpkWw2n8ibgifi3zO6UfDaNE3jJWq5wNKexmIeyBMJ59n7xZiY1CL+D8m
spgB6jm7nIhy7ssc4tb3Av64ziP9w1/SbpPa44Q8TqTGNym6MWJNh/L0fKpE2I44
/WiNX5RUtKcsBE21k8JYphHVyyNPJ5f4eNrkqM8SqAoVRR8iAAiFSkCkPOy2L4gX
ZsYOvcErdPDqc6Ci00Y5i14ntikhF3HLu+DHkg69uv5oxlxbblp5e6sUo7vT5zWj
6IrPB4nrzhPSvKyK4lKbsbrLUpIkicsVSC2blotiVNs+6MNzyx/75rbvZjtzSbBT
MfaX6Ndr1PPGv7JashiWK8CbKf6I7U0FACb4P7TYwiDnR6NfrScWYoq75gdz4S26
U6MuRJWdClqYF/N/WTzU5toKpr1d2E5lZItGz0F/CnA21zzksTDfauOJzPP08lqj
f3iltF3HF9obJ8ffKDvOnvc2SYL5d1v9e4FDPkcnsrVHURPRMKY088ZZwJTH/e93
w+2jRY9NH9gCM2W+uaDpi5N0w+h/G8jWu9xdJblBaxn8YfHVtGv2GO0lFZLmUJ93
hU8NHWVXu+j6YXGALJkKkEtwWohLUasoPu7X30kKQjZVF2FiugrXCGz5zLp8oUeu
JtVsewvjXyfmmxcdtB1NQp3eGGf2ks4PHcYXjxFjls3dvDwlZ+pAeJu3QsxCFf7t
iX6NEGB8QIKZEOKJfsjvhoUgJ/gPT2tfKdaYJwXtXCjng7E+psx4JpCqtGKpp0UW
jqODa/2LyIXYZrriROcrvqfVbQ6gPhrLbw3ZiOBeYaXZTZxsPhJ8yj3GK1/AeJGo
jN0wxqBjRrh4lqu/OSwNkx2o7Lg4W926bQ8NhLpar+5dvB61TS9t4B8+9RxoX59s
POxMvJdEf5TnlseeNcaskSKK3RmBZrN+BlS8NHRijueQ0BALpIokC+P/C656/RQ+
xl1uCbwWmUV0FkcANotLqvLfWLfC+iknoP3G8hjncHElH/IJwksL0wMcygbWUUQ+
0Eaa45DE7UDE9jrEyw/sGVJHaBR/Jt06kVSV/tIx/0nK6m0uFCMPruk2l/MLTJrc
jbgvFnQFEuUWlgFwhc6ikaZ0zJJtkzHCwkSCrTlsqmSAk16+B4eis0Xn9ARTKotr
P5aI3k0PcC8dGRCVxkZL2uvUhJRkLwMf0vf0o+nDrv+tPfJQgzqXECuACwB+rmSF
WA3SDvFJNB8CY8CMXK6xz3KfhzSdFe46mviXfibICnkUDJbpMjFFuqIa3NgXXx7l
FRy76cjlA+pYXw01qH+RjODQmKEBuCffa8volLMtt0b9JrR6Q06npuv8Xs/lxAZ1
3GfGW/k4iYGznPwO9MS/YpFbczu6gGIZ49XWtAku7ENXuGUNYrJrcGKcOPwW7nHX
uP8/GWkHmpT4zkouMYBczqktekZ1s8CDtPi0xbS5wvEN1APaFFh/1t8AxhD00fAe
Bjg0Ti5ILHqbE0ei53ACPCInbfzPkdVrgeUtyIxPQXlEm4yWSqOMjkoDRjPnabkW
RynIVlbPDQcm85MPoWDH5cA6Dg6aZJpzjrNjI9QTzTyL4Pqw5kjoUzJ3snnUHzvi
gUFZJ5IfnQgXcvXRyJlmbtiZ6vYkJNoWO9QqX2r54RxnHXWMiRE7eJTCz+cc2+YW
qgWZCgOnWuRe7vlWnqfdHG2aGkaQc/f2Hxl9bVfRojdD0SV3fVe++hIsjX/QJABK
lkQhezes5Vck+LhGOWQiKnHSrDhm8527LzJsPVehUECgRB6ay7limf7IIGjnuy9g
m6C+gUAgAoDw47jNwUk8MfP1MK9rzA7vT8oNlz8TBf3N3h5IOt/qHizs6oLPI4jf
AcvYnpmlh8DXkSTJwE3JNsUBcAW2lPK8tX/zzWE7AIOjxiv1jRGY66/aAzqD03bN
lSibxU8cWpx5RiT8xrfziam7EVsonQCYrZLMBigkG2Phfz0131jynAtKZbtZkwQS
fhhcMrPGvfzXlBHAWBsSwHgH1DdLiNqwUdUgT9/2frHtfJU6VMMwUbzqXkyP6959
iB6oBjJG7WBSYnqXoAnBReSv/rQn9WePG95AFBO+rL6/bWC4FN7xPUuqU/P854xj
hkD2QyQMLUzYe3Bfi919AFmf9KURshjJwSFNkLp0B2GNCnt6TfuuYwwx9mOgNI7F
eric7y+XkFng/KmbMqhK2ykB/SYqeAHoBmCrhPsd0KV85YLLowKaucYba25p3Crx
+4fJD0LmCLBaSS4QlVXjeud4DDedtAY9WjWaWcY9UaTN16ctqwzTz3IjzgymEpxz
rgNjBF/mHMTiTnhTpb7eNeZM/inYRtP6RznTk3ihH/+Ds9xpTNrQZAUUS5jpztTf
ZWAO58fYFahXarzuA+09oyRlKLT6hdydMKsGNqs/W61LxQkDzBWJ1iWcbAYZGTx1
rUti45aN8WoHC6min8zrIDp4vnVawmChVJbjqzglucnxnhHPJYhCbI0J3FtcdWXn
aHnjuMQVUogsqx/DzJ3CC6ZqCn275k0zwCtM/8Jr2b3FPSnNY2XpCF1FDtuWd4K4
40JJlhvl1HBEXn+az5FuWWPItwd7kBKzJczMPdzOAtMhvrVZF50FEZhTwiXuwu4a
dv/ycq+GuncGXMwCNApxGN0wC84KbwynCJyeMiT76JKQ+/myzztuMRmD+Fh7VH7c
slmIsT83/zXlMKDw0Iuiw2sYWu+zJSvE81lWiuTgLBJnGRezZugILE/MkomCvtgN
k9hBRusy/6MVNDNuAMvQ09ZsHvnJYg39Wm02bxEIOja3MzEkNcq/8TcVU9DHvhpR
zKgL89EsFtNi/pzkOOLtJ2MeIqWwVv70FHXHArPOzNAgB8wbFHJIFx9+jYfIBgUJ
6WqsFQKN9C+/P1pMOEtqi23jnygrzop/oKrC4979nzbZkPki5QIqPtUepvq3iEGF
YC7SSsSh3VFQjgX6IjvLOw6kGUt34oT/4gY9WQrOTAE2v2WIRPkDVwgNOjYZqLAQ
coZ1ja86msQYiDJMyYbQjS33X81vhkOnKy/cxm2PzbYH3V6oN9dJGScNzEKzLYrw
4aHD9BBSM8QiwNQGkCTmf8+y4Sd4EfYGt9N8VkHzpkZtjt2CCkLCJxv+JHY+P3eo
JbMw8EnhZRS+zo3wsvVAQxOzZUv7+4aZPYfIdBPFFJw6BUze2C2AWdoRp5vkUb/b
cCOKs4TXnxFBryLU2wYk4jb0svCvi0XgI254mr99cRu6nreT+QtTfVFZxNlXik/w
hm02n72PuRbrw6fWUA8t/Zd5DVLdL9YjMOTvdMw46F3eOeBdVucBxNxfWSDNewgZ
Ge2+1sQNKN2ZZ7WjxVYRgk/GvyZ2bvcCvIEh/MGnW6EdshaYTU6d8XVTsgnS0qAy
8ap0+RK3McyvchVUjvcVkkOZPjUhm8BbscMymiE1wqSnyqMdcEcSYndA8VOTbXAH
YRpedJuLaW44X6fVnTe9UJc2c+tcEbBzH4zzsxFWQZboxRtoada9NsFRz6yyck2d
K/o8HcI1jIlf3C+x0g+7zQoZA6cE+f+KHzlKuQSLGeSwJRmokGNL8lbEM969k620
ZpYz8UYq/ZFaOMmUfdD2istZwcJdmk1DOwa/+1vRPP3o+krarZTSttyqZsFlL/Fw
bWJu5AeoS4oJPa7RN8GRGdpeYfGjgEKrGD7IVjmq8bJl/taSh7nNxyDXwyk90KBi
6I/24hHcldPXMR11XCjpmBbwqLfZ7uuS4hD4i9+TzUcSs4U474p79wQSbBWSmUPq
CDiMe84ogplLQg2UvQn+PEV5h00SZE5m+JxWu8G7v9GP2RExuXt+MlBdaYm505gM
JUO707U/9E6QcPJOb6IFFyAM0dEzkoMA1h24wZSrDraArdhDDKYZaKR3O2xH06IB
/OXXsqSulBwvdpf71iWtsv6CTPdykx+bxrZ5GtRxqqVN0jF1ULwH8r/KvkQWHEwh
mXml62YG7gFP5Hib0PrSASMD0gy2hfPS4DYOxy+nPE7Vk0BQhqHaHQI/bl6d+D8s
3vIBZi5QQklS21GWRx/uFXNkOZwRM120M4r9xUf/ZSDwyRxw5p9VwA5dQS+FMKos
MMuCKBEM/ISWLPX2miVpr9mE0XjE6gunyYfisSHaiCSDufF4sNjgWozxyi4famOZ
YT4DZCiOO+N/6EoAm+Lc8YUjqxGqWpk1HZLhnIRPFRXNNy6UxzKDHgY0GG3hCIZ2
z2d3Q28fedvg5mniFox3Og4gn28baKygEg9gojtfrQaUMlYHwonFcU23lbOH2UUz
TVUUmwy7X3CBk9+xyov+pkfummcNVXIy/luecA/utewNjSB+zKYjrj99eRmoFJ6d
zF/5Lrw8G9LR/Sfi+S1XpGa2BJtplD4yjP3e0t/0Pg6edOgNEe0+zfsriMrsQ4fT
MMN6TnhUyy1nMbWF+l1bqSrJChvNqw1CaAzAoksIneAC3GTw5fb+RCrOp9lsyoBn
HYzJSlAs7mvp8jROntj78NHIjO3csFrDBzauAJoeLAv+Im68ZDyWTwYs9m23AvJZ
9Ov0Ck6oE7+AhGApjEKQZfnucmGQRt1kbEStDiSSLy3mX4fF5mPUX9pgPTWtzWQM
7zzuY8vE6ZFwGdzrzu++lcASW3yz7++jAXijCOPobqmklX0pozhXWCBv1nBu0WyZ
cHeZrEzWhZkiQUcdmRkHuSLr0cOcsgzGY6GoFB5IHQEdyGugPGBDgBAIQ3k9Dd+m
jDKDxT/fE7c+6GlSXDmO1Bwq/hbi0v7s9TWkWUVol8yubdEIz/LHb1W++3DwLDzl
yZ8JyC0AZGX7+TIuz7mzVb8LjCn4J7OccijeldZgNULExSZVXvg7NCtrhY7GnIuu
VZuatxcU31gdGHrxtJaRTzYcvipp+jZS4yztPahs6E5CYtK2SazxK6knYNRGR+QO
vmI3diraT3VtD6PoxG0HjGXAYJ8kSg1cdl25nsAdD1frc98wBiUfgD2P72fG1DD2
0pIq0SMzn2zy/7mPFG45049aaiOQ3WGN8Cr+1taf18CGwLA82tSQI36ecbwsZHLG
NkI9+0ZBRTLqgRhw8+WwdP0/I6WpmlzSoaXiFlClt9hzeQ0YlcriSpXwEG1y9dub
0cwdJ5/psVRRBlafmkNyFZiDvAPBJRoi2ysGeL0nGyHNEqHnGniPUchSLcv9nwQF
R0mZ2Ddw8eCl/GaVXXlWuWEffc9bPmizMuTsUbbSSWsyqO9pHPf43nqR/tifKaxv
P4UBr4H0WzG4dB/ufu6iZ2QgZTK2daly05UH3ty5fLf+c/aEQm9Is7H44hEyjN4u
eWkw6Alos9nS71neghYehAZDqhXkkPgeHs5Yy0THSqTqtKOZ4oKy9mP+lgiieMmY
fgKEkDPH9j1xYO1pyQfllq7+IyllPbOFetLMDVxQWW//aAusudRTW82y0D0FCey9
tX2AMD5YSVPQ5VS0wLqRBQT7K6tji5WLjJnPihpNxGue1Ih8rYGNQxFASwZo0/BC
X0/zaaytqcFqe+RapUq8YW+DYtdxy6io6swJ0FzQBtQeBGvH0YTW2vf6meaJqf/y
YVoJuq6RW5OgNcYe35ySd3pRj3WaRYUqug5bRxu30pZiwiF7UmWRcIDaSWZ0IrSX
H/HWhZTbTCK2K6BbRnI7Pu4VXZ1RRY0UDchZLrktCZo2nrKkPJ8CuTfXgZuiSGpf
/5LGW+quR1etzF31R3L3eNvizIg2TGFu1dxJZ+r3sxK7cLM6lkuZ213IixiD4n9D
CfE8Z7CQ6/0a1GNpypXp30mj3CDAvzbA7tIR0RCQb+72JzBhQX2mVs3yeo0vjWEJ
pdYQmi6jinSxsATGBTajtP+dd6L5MCwg8tZlLe8FIL2OFYzkC5ftHQ4iuLJe5F/q
whrH3f4vQKFJ5c7ogTx5p2i/ghV3XM0DIODPHjN/snqY4VueC3d5XxeQZcq8I3xv
+AHOZtaDf6QMlpdGBoH9u8mqDDdNRlcYKulzj8gHqmoDzVWamk0KxWUr9XDiO9RA
p1fpkDQal9G4SFCemt9D4lwtYmZrvYeSeiyvKktSo0UfoBgtnw1maINcVnlKiExt
yxA7oEoeU4zH+0G9AwYeMfMRSLs7wKfZ78BSsIXCfQyrG7uwFN2holEy2nkWVoJz
YEOH7lApqbFKOwmtUF4ipBD4q188d7mmADj5pUux2DhZaVi/H97j2mzKvtXS0GCF
VD48yOldZu8YDpr9swkmovxpwQ2yrnW3IkFkg/Q7CIUz7TvFyZiHQ4Ffbvwn4dpE
N8vDLXUAHO14c3Eh0irK4nZDCzT9vaLejeRwNeSZXOzWC+EQmtMfkuBFHlckqsK6
J76HpkIA8DSytsNmunsqb+/u5OcgPyVhtakDNTl0mzn6nr2QWlaQVN2xgd5ICMo1
gXr1jQLgSCNUYjCCmX1Z7kV8tl6aaEMg/ET+S4vlM8kByuKp68ZYM0s9JObQU7Me
m3VUrC/QnGxfPPA8u/5qvQ50jsX8CaRv37FSkKJzBglcrnc+QdAdJ36JV5TY3gV7
PBHkvgojC/FeJHFbUZoZIduLGoA+SHqcosHTBO8BJXG0fsgGOVj305lfJMv0FC+L
3amZNoDyR5xqwrDsRHp0U4WmLjzc38LB+tnACcCJbntez8VaLaKv8OHhRq4bOz3X
d4l6XN7NDQDwGvYFWtzAtIG+B1p9OygwNlVZQiK0a5f8A2sBw8RojxdmRS3NqoVl
3ZpsxHjreYX0lFOgT7+x9l40ymvXgWCRRBUBRaC15lCA8+9mqhwD4utwC/E08AS0
0ZhiNyQic6nw0jxPR3Um8xt3sJz0FiKZKZuJjlZ7im2TRqDPUmz9lp3hqU3cVMXa
GvCLXCKYpfLjMZHAv6gStUkIkRhoLA94xU9MOZwyAaDz61sHioRTAfV2UcoaZvNe
RPK3os1aUvsjTIX6g+ITza7PMh8poTFd2yU2mg4dyaTsU1V7vJFgh8ABUffMPIYU
pyoY0shPevUIJ9izu5g1IT1PBFzID0Ey+rxQPkyFan8EzYqSseTGdlWUKLQ6Gpjf
6B0NUCKAFY7QAXBKVx+AuMMZ5vyb5yVvDq9gVkCDghVPmtBSBl+g9RfCofDfCQyZ
Q4e2rLo1+CJk7E3m1zBKji3ku3GRGA+mlMdllD2rSjAv3Ya4cOpFBEgrju4MFtou
n9r46qOPkBC5hv51XLiJ8/fS8Yt1KI98BsUczyeB8/rrhGIsJR/95pLkwpBSEiDA
ZPFvLzuvga0DNLzUVXgg+p3SMXdMy3Ed4eN1KP+3cv+m9x3VvVPCLAWbhmXdMeO3
cRSi3ivMswL/lq2pTr1aylWJiUe5rgorNrm+Vf5yCsbn71SFIsmJjCe23dKAcBss
tWCag2A355g3Qs8xSllVIbK43KuHVG3HUd5fmG18+hXcdYJhotB2tmcvm5vyddcd
t/J+ryfPBUBxqI8JCnxgubKz6aoEoM9qBKrm5slSMd1QkjTaSAqMpLd+uGGOlbBc
G6IBJFuClFTZTTvy8aC2nM7Hy7a7aZ1hVftjN5uj6vSiHYR8DedaDxE60AOAVThD
tC1730aNCXr0gsZ6UAJIPmC+Sd/CMD0NQwXW/EYWcvYErem9jsShAXz9uCLdb6yv
TtDrAW5ToGDTET5uv90uOnBo/zjQHf9Blin8t+LO/7/WKnZ92xsWQx8w0r71soDi
qDiClQb+BsnW8szJmpWY02mug+YFrSneGVEhRRM/YR7x/i+gcT6HoPIJ6nQFlm/Z
hiCDlnUcYWG1rTU8RdMDTdJ4yuF0hWKD8RLtrOfM7hXtHLeA1Ftrm7VOMvK5ouLy
UlzoBjz4Bl8HkPXL7gi7yR6GEznoPOKsWoKlPj686Wi/tL5HZYmdAi387Ds8CKqX
sDkfNg71X5+YW9BQA/GPLKN4HA0IrhzbStTUWU0A7wIDgAiECahCtWqqOuLIoyjD
mXyU+m2wH5hPM+6zHUd+xQsjHlO7QnLhpDRQXP6YtjudyP6hVeYNqlb/Xv5+GOUH
d4NV9eLA42IOCzdbHzuil0MFquNUcwofCvc0y1I9uShvr8a8oqZ12ELYAdrcjcbE
p3AXtZgGfFYrlYDNfWdBPkupc9ldmIFsLKNkx+sq60xMNyQeL4aYz6oko6wWCnJT

//pragma protect end_data_block
//pragma protect digest_block
x2txFmx8/lTYRs+Cyh+oN/CB2tg=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
9ZCqgaM2iOzG5iCCQmUMDKgCU06kPm8ZjabXbl3Mg/bWpsd3crQZgijRNKnO1Wh/
OvHf9G4jG1e6Z94mSw9SeWZ1pCA6oeUPOuX61speYBzsm2HuMDfYES7YvzLayCUp
GBNr6hxbstT4Cxm1m0cW4Uv8PSlkcQHR5QcovqcrNbpkwoUlrxLYbg==
//pragma protect end_key_block
//pragma protect digest_block
rnx4cioOUs3lw1rhTLT440VTA8k=
//pragma protect end_digest_block
//pragma protect data_block
YrRapbHSTt54GnfjWnoBRDeQkor7YYgxxiBa4uZyR6upr0LgYfOG3slOemBitKKJ
WYBjgTM9J+WsMjIhCZfo/i3YnwTRuhafQEY4mV4FYrAsOU/6RLrycmqS2gRKJi9z
3bOEzfxrggrJ35mVjTpZ1ES7ejnEzJzFPd1LfGTioDhHAliLhfXlSU2N4FcJsQOg
vEtsfiEsTo8Wo9QDlNLNirijYnznq8SboI3rkZmFKyxELLdmDcBe8wdqQq7Nq1mf
HZFhSeyWS2wPJ0Lntdx4K5fN/EWcIP49EuN7kTwg1kDm/Ifs+f1FBFF92df3jzT2
JLBmwSV6kKlaVP4ullO19CnHRMFVSh8gBc5iRcb8eoRIKwPe/qD4TOEI/BBEuSiA
tVoBSx0WS5BeCEg0fUHJQNEPAa2h7QGoqQkfF2M0BWDbN2lk3dxUWqkbX3oi5Pay
xEcslVZyWdy0mfH30BeiZZtEUE02Key+4EhbXTfuQit+qeAE351qOPqPNltRFfOj
zpRqXjTFtCKNEvcpGlrhm1PwmNGBGNmlrrMgtlshOWEKh2Om9bRL2Hj+qGFzABB2
aIJVs9XeUgddOW8K7LP0mkszPf19vx/jbk7uU0yQsmkoBjiec1iAHKVrRqxYnpjb
l8M1lBRsn4ZtcbELE2YkQQG0yg9DrOfUrrrmD+cNfyzHUQLxaOM6aW23slZUc/mX
lQ68DIRTabLEJHYwYZCVFHRjXdCxuGexlURAhem+dgtzU9WnxtqY+C2Rm2RpP4ke
ImpH5ggNwF5O9tjxrWCBfsp9RjBt7N2repV+FHc4ib1KUvjyOPTFClRC7lWfXxfZ
5HgySNBBhjMgdU5vndnSAdFS1Sie9o+c60p0U4LNMt3vIhvZj+kT8dhT0+EJh6QI
I7Uk4VGBNxTAtErXRP5n3rKie+oihSkqFWM9znQHLaD5nJhpdPE1xf9zpeR+UlXe
n4tyT6bTtdpCAAA/334rvB6tbgtIRcxl88ltY3WW5a5S5Xb/3rAI1VeY2vN+wZyD
U5eYYSLoXQtWr5QKHzBwSUZ3zY3m+o6bn2yLqnJ+y10oz1F4ltm2U4cYrdCUlivc
uGiHWUm5q60CfIVrxRtovjSyaen2Eo1TNbXTfZJ/s+SceCIicPRLWAOFVv73Br4P
0nqV/0XRtwJFSXLwZyamEeWIRDkOw8CNwOuHYRH7Cgsv4SrOTKyX18qVvBaB2EGN
aajDekiOFD3qvDWcksNVeACwYCG+QCiW4NAgImFrRq21u8kZ/QGA78mngVhtunvY
vx9+UxcS4Zf2OhVekDVLii3jcDL/3NhLnD02mmddTgEXOfAtq9l6185FD0asCgsv
/i9IHhE+6dZzg4NN7k8XckOftKtaBnmIjQ2o35TNzkbdWM2k1E9xf//8OuVQSG8G
iioBeUquymvHrJOzcQr9bKrmGMj8nXrelNzj5tT8Jin52dnVsAjILblqqjQqdvT0
terQ6b4lqHy3DUgXYf4fJ+8QllwwAEp2a/tMWiv+i80weukX2uJ0diHhKbK/alwS
+uP8hWR3uREjleHEIuh7VLVrl7s8UEfw0imCQd40ucu76THkipy7Og3FIDxKjcBo
JqvOqj5VWgylDrv2rV9h8xMNhpDqpoXDQ7oGU82/W43drLjSAgtKAR7V7u3+Qd0q
LivaHCkGeKzndmmCxFrgOTUJcSD1fzAUUpF4aViWeehH0+4RwjMSBShDnk0VmFNn
aCBrQkrh3rexm/tsSQALnmJ6qwHMWucunAbVqNjkpjIJvhqJja+EIomzm3sbzVX4
sleVHYrUBj+CrfQGMXPUS0KyjJrxwR+XRPeAXVn340rv0rnYm69hYVEj/pU4pQt6
C6tEO+zYTOF+A21YN6txhpRp8wV1pRNPQQ57+XaAjKL0YghIDlKtAZHm8tcfgUbz
DAiB1jFovE3hEh9KoSZAUx7X/aHDTZm8ZywhAszp3rzVkrdamQL7nRHiGXOKXpDp
ts+DppBF8Ib3LIrgE8EiEJheFXIzN9gM5FB/kIFTjrYsVXw1eP+D1tCY1PISPwwp
pOWbomvgIWb7RmuIfQtHhKfXlE3MnIKUxOhX2I11I8Z/n04lJQwmWb2g0vrKi9PN
6qagOIVydPNujXODKhxBNbIdCPyTgOQQEBgbrURJGXH3XWe6bTt8dIfa3QXV5Fck
jS6kLp/mQAXPnreu+9QcnzYh7SJ/drCi4f0Ojw7jlZm8dAew6lcSqpUihY3JvwoW
0JHfAoOHkZDRDOhfrFt4+ZLGYE9mQla/EgmyIa4uv1iLERiXukpPRqcu7poV05fU
XoZLZdk0V3IUqIFbZJEiRIjtHyFlzb49JJQk23zNICeoNC0486N3UaPf++AOtHh+
0XEU+vqD0Q2E7l7r50ZgQA==
//pragma protect end_data_block
//pragma protect digest_block
zgt9tfCeOv4Jovh/N/WhI/ioPKo=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_  protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ctAX2td9VQZXfHDLDySOCkxOvg4GobCwWE2hbVON+Hpy/n6dgTe3J+62zr20n18u
xyl1USpj9ZLmEy5S6gy4NlhGQ3CBmuE6d9QqmkiySZSphdtPbP2f6L3R5fcpQoLe
Tk8sck5PMSL/6x9L/0YFd1eDKHOyCHz9aVuHT1aABFNnApj8zez28w==
//pragma protect end_key_block
//pragma protect digest_block
yBV5nrGXWEFqHlZxzIJKrR479FM=
//pragma protect end_digest_block
//pragma protect data_block
qyDGrsU02/61fun471yjyGqHNFRBtZS/bgCzesy1ZVTCI9BzCudT/MS7f4NODp7C
/BCGAxIpmakyYiVVVC+vU5FYqCWEuLOMQqquNzAlXQV2qdXPeGPHNKYjWQSppVTR
waxiU6NtZZxW+MuCcQmS9x0zkWk1j0njtsmGVBPQwxzeIb9mI47ULeyllOYkMfoL
qvNmldb93OypVz7HVgqU/WOrqcW6qMWp/hPJH83ur9oq5A3+iCxmuBQY0jAM7eZB
4AIPNlY7gedCokCtI4uhenaN1RvutYuOGYgnX7u8rhHOF+uthw3zWz3bmPQ3DvZc
g15kppLB5BfLmf0pPh0xqctw8fw8iYFPLKe1YtN5BCjxSYXSXW/kHQ17A9iCF5l6
1/MGFwZR27PfwmowBRxsNmrVrOFm7QfXyFTS/rI4UNLPaDoTrgkccDNiS4v4N6KX
aKD/UO0Ti4+tXwUGHEEcQFjkR+Osg2/plPm6FsoB5atymr5fZUjHl8APuHTiFpIp
kDVxURTdB1/NBxxaIp3dBQexXd/TTgz11KiRZDWxXasyZg9uuxsCy+GkXX6G9OLb
RdskxqRz9IWv5te/g2kvdmmkL7VzbtNn8/gF9xrM1a41hCOw9c3dXpQxwDtp3MTQ
apxA1Lc5ORZv3ZRs/nBHxS/68Bx1q3IDjaTkFhbEH5bK5kD1RZh8bNcEMIQylGCP
5lRDAPRjWkUOMxh6+k5K4ZhnoyNuS/Jy4H2fRpCdaSNVGr3tdhbUBNnTOCmVACbf
50UtgL3s5AKprnRkVu3qW8yiLn5EudpcsdHvZVtCrJ1dIKQJ4W3QvGGklrnZK/jV
thxPCSSgAv0RkUlJDHvsVFK4U6n42/T3eLSG2E2IdDH/dLPIREuauR5NCfNKhQfq
tJRFPOx7KMFoEicDUGCG2FjyGiWQmLTYI+GAmUxOBM2qkvsbZFWFALibDEGThqfW
tGKwXYCTbqNMT43ngECrTcCCmKB8lkBlYIqGiE9LL/r1Sn/Q5HFc3To0cI5nnDOK
urNjs0vVdDSkD2L4qf9EHRfYZ+QRnnF8NXkorsPoqzJE5xaOYZyxUEidDRKHvn0V
NO4L0jpPOgfEjF+RP3xTsmKA/O3OwF9eUmkjNT9B0cSR/sGomna3zrBUEg06uuhx
nXNgb2DKxGlNJ7gxUHjcCWmzRqbAWCUBofyHvfP0JlPQpDZMoRmkWVcnkJ2+/C8C
4MI5eOurABwlouWVLLskUJfznW8p8jBVevH1j5LeyPjnXhXfamx/WtIwVjN6qUOB
5BmRJNqReeCoEq7+FhqzsGGa9cpM8ZETGaeqORM73Y71tjauzdfrqYomqPYlHAtm
WztHvjOmFnStz8B9gXLo+FlAP2FIgxP8hGDPvCCwqIcyCaxTmLLXFQjGvnSjBc89
oZoakJ5fuyiCrOCSuBv33a1N125rWIX9KHwrJqFbwR8BQYHgVt6OtouQ8f4iFfEj
AJwwJPOf5ggx2EGAlUW+M/3PY/axIbs96yRGGw4r2y6Rfu8oBRgynBw9XnVm/ZaA
g1R0oXRthQu+WvuBP1uM4OjE0iEDsfnaSKw+WGn/7osPZQB/9y+gn04tZ44Owd65
HkpOkZHIIuyNm/guKzsjwZH7h4FrBG7nuYlblxjVEKEnoPgohBvSSoIFF3fraTpd
3F8bJyuPghVlsLYQH9n5eXSS1YrL0ah3G1LBKugu3dhgAvZG2DGZXWeKnCcSM8HC
SOV3DV+4EhDcryWx6sZDdqagMvUkBk3Tl0i6IjRCIXHDdPSIxiQ/7Q8xEOl5zsRK
Fl8nABORTNL3z2rmjaKnYYPekxCT7dmzVUGRRMi2hJVek4WlZk2b5vsgMfx61JUi
49QwGyQKqlwCSXIJ2oA7C2fnvDwZfh+nnqdVY7RkBrtXK8Pwyzih9mgwAUFaZYLr
8Vu2aCiiyN2yWX4NhURwHbxHmDKz80SMaHfY/d2QFcDlm5FS4q2E3QKVCYp1rL2r
mFzmBUq+Id1KzTtdW/jaRFTWkrXh3Pbyv38KmpBhBnBaE+thAiT/1upx28fQjpPn
TdFD6JuFX61LPcBF38UHaT93uT6cXa4qG9PcvqUE9bTws3tq4u5g26yK7igxDwMy
XIxmr5KS4BZfojEpZgyCxKwPqvhe/jMmTglPG5bYtUS05NDeGFQaQ235WZiMFVVt
cT1PXn9GrJe9PmXsn8qGwUBevTVLgLJ36OsaHGjmVC3z0hpA0fxdOzSIU1f3Qbnw
sMXgRCRUtU1c/COSjpY7GS3xfRTB8pDJCa3qmA8PIf4ZibacUEYsjgwUNR9zA6PW
XsSJT0NetkHwIOrF9jAeEI3eiwSU7LeR+BwoRxlG3C7xsKZQ3aLKngOFjjAWIvQI
eHtDGP7083q5Fpi4Ik5/esC2lw8IXKYJEo0D347+KsBVlHx32XQ+KNmbbuwRMcle
FqWP9XGzX5/mU0fmAkfRwhbT0KOD11XPy3Dc8DmIpY7h52+lmLeyKfiw8KQk+DxK
wNdhQLVGgdZ7XveEcepxUXOeoHtbSkbABSnRNSEadgQrCYpNx+gVMcJtWn8VSvCf
e0l4ll/UBuj7ldah31hp6KXnsh9n+IncAKG2sA7wGcCmDo0lT0iyrl6xl81HBZnl
CVqn+niIy1RGUVzB/wTQCDKxWDLT/6yMyLXpwOa81tYiyEYowYzvv53fxXokhn2I
zGqpN7OGK34R4p2/bh3qRbAh8dO8CZlgktTHXqCBBmsGIOw77m8FXNJkV+JHtpLV
K2bvyht1NPzlfrbscuP9MaUYY0+lf5ndOtFfSrDWsszmWAROjZmO4PtDP9rhEFRW
DtgrkH+MDXbJcVx0X/Jy9jrmlPLlimZGbuOmniES0lurr1oRNj2QudHeqmF8y64H
+fdDNKWkAnJEkHMKr8JZOywf7bOWUcy0FuIZoPdyWTXDC1PbnUcNar7qgQcewG30
G24VhtcJS7E+gtveV7onr2VGcgNIFyL80i0fX7jIa0uzYfqERfQYVX0OCySElXcd
BxVBoiXMbWGKzTdUXHgFsa9+TlHKFrrxZlXC9usqkr4nYlzUl3YPl1Psy7B4u2Y9
QZx8gvD7nfTap/L8w5bEEvpLOjumSfLKBEd/5895IpB6m58AWofh1J27k37UjESa
lllnzWHaSGbLgKxhDHP/aXHIoOZZIHUfr2yNezB9a1PkMadbHE3fzION0YD47Y6j
47la9P6dReo3KQo+RJR9Eux0o4gZSSo0+jK2JhGZSWNRKTubnkMdEmXpFv03fB8z
x1i6hSb/ICgn2rfK6Fuhh3NNcZnLBqOD0np/qWyYg4/L9BqQwB7mKFcywf+Dpa3H
YOul7V8MGOZLRwNixoZyoeRVHsKRTKtqs5WpCVD25h/QPWgvO1s/f/b+5vwEXvFo
w320fXIhENkoNoeO+UDUW3JdaGST/8gvE9ltc+p7R5R4lWqDrfQ/vHOxs2nGfCI9
RKXeRdDl/bJu7gHBsjkcKWSxlltjt8Xuu4gYhjeOMqL50JEa37bbKGfRduL6BYTc
oYXgbZJ6XyHlEQTl9JcqNciIXGapvoKu442El0Yt7qZTUA1G9h2qylaZECWB8Km5
UBQ+2Ijrt5Fn65WJasgibLtJg54gEQdTQ1xNEhlKFL+c9qz2iNOcvOdDexWo9YLl
ASsJM2RcKVDons9wf5kRShU99S8PcrzeW8oxSmQxiMacwOPrJtelqrT29ZuppRwk
29M1TQSg28JIBjKfZov5XxQRB8ITTjIgYIMmyXbc3c9NDa4wizJTFCDrJ0rVOmsK
mjNJp8mh/+Mr2MdAtbHtTgJTdY+TrqOZfALR/ENTfGlpPzamik4AMPje2tZA2f5j
w6SiqGEORroQEnXEHOD6tU+hIUiuo4ondISFxq6nZUf8BcZmpsn6xONnV4fcwvA4
XAduQZj5QcV6o2CnlY/HAXy9WyAqXYsF+uwY8Q7WDOKCZBnMW7kwcF5y9YQLB7Hq
sH/8DJIKpxmNAWuo+4S9o1pXOEWTivjNn+kjjdNGIWODANlO3G9bJn228Lgbp9Zl
x2HLOQ0LJHCiDLc4mv2wqbN2DEjxIoTfuz28BIIkiFe5rFIFFS9ZDHvDHEy6NWwK
xNOZ51oAhkum3bdgU+IdHNtsF+ijiq/sA4pVjPOyIHY3aTW+VO3hZ/2p/rCRVNXa
bnBKARuYuEUt9C7TDGkllz7mDRDAuJ39nhfxOmkR5+qIXfNz6fso2pISIosOusfh
+0K4R/KMy2jx8ucXZ8g3/FUY3jT36ypDKlxaRDJj/yBVH+rIBB/fBhF2lRitibCc
U7zb2CjqKVQQtd8s09WkuK+RpIIsA7ody9n9RAUca4/wFW4FwKSk5w0HtF08tkZA
hakS3VZ5aVRW2rUbFpJd5ZuQs6cIx/aRuzvtHkdVj0/pevb+ESIY6W1QmW7EfUMG
CTUBgcC9NbwQWcgrFu8g7LtxxGewDYhiiIS+9JYX02pwjC4HXt7XrcG56fPtIKnt
9orvW56akkXEJWPMPTDiTbhsvqYUZiF23MPZicwKHPnw5F6oOWo5kGalU1IXPBlW
UGCkBNzk96VPljJgXXgjb2zaWtlkKyimqHsjFViKeKzkI5lrZ7xW/bG8nyAyJIRM
I23LbFq8Zegczpsx9uOlICk7neoF2I0UNsnZL5K7q+P2K87GZ52bpRmKY03r+zLe
HLbpmSHjbNRkTEJv6dPZb2JMtaseVG6MBCWPs3HCD3KN58Wy0k+4vlebJKWyITOd
w+VyNajhnxp5FUL/bdrFGcWN+ROZ0HWvBk0B/xb8GEiiI88LxNWVbZFlZNr3bFkK
4EuhCSKCaKikkPdN8+QUxfESTHVao/cF/hhvEPzimSPQHcWzMWMbxPNPQZxdGTCM
tCnfgb2jfA3un684KnQsSJxSfr58CqLZLr2jpXXYEY5nY55t+W5kSHeR3/GIuPSO
YXPlVqz96nLtzqbipHzt9ueHVv3KGvFPvf2ZDEk9Tc/z6IKO7vfQif+0QEa+7VZs
AoWYAKR9UkgwlSKk0KmGjoqzYAON+4XgIo4rIMTethP8m3benC7ic8r50sNubFKx
tPXMbtGKaGt29pYyTdYqpp3FuYez78jbxH/HihYogplBwvr4DpLQ0B06afR9p0SB
xt8dJoJU9p1VHxTzIXf2d82wtR6NzH2gmIU7rDEswJxseDFwyjhfuGLeQ5pJG6Y/
n8nTmqS8Q13bFpuVCYYgHmwiT2yi8WCkVLLOwMkA0WlLV8GFkxUgBCaT8Vtmw7Rg
aT8aKfYrzr/Bdsxdof3gKrcufHJ+v72RfP3I3vHa+EUSjn4fXixe6cjyrJHCsI7b
BHPkXzD7fq7eyRp3NKyxEZ/BkodUhpDFdp1iMNOlcPSw2vI0EqaOuMkBY2q6bUnR
N3Js1UFsOJfg4g2/hvbXSaP8hbd9jbzv3qR6iMWOn/SDejFCBKS8CBvAzsB5Nlkj
K7cQ1HRmQchZO+jSkh8iuAxuyK5T3Wab6LIz4Grqojui8y5u8wKETEhqDAzF2vS9
uNH3sVnXHloSaxNaYa+vlxB3L9FAm9iUfooBzMkqLCEvHw849b3EjB08WCZDUM5/
9sDo9vqgJBHtLNS/AU+F/kLjMUlWxiF838usI0SdAT5TtVA3q+bro04K6hpsPRQ8
w09v8GDma8buR3C76IjUN/Z1SQi3WOksx08pg4NJIpxo2X05xSpgcgZTXldxCNBA
CkP6UrxU/B96uujSkuUDI0UHqqHNxTDBnEsY5hJt18NmBkZxVoZ6P9vNbkLAwdYK
CApscdgY3NeQXWDmzsyyK4sAO/pDwvme+pKtDkv0dZlNFvfaX8AYlwuhvytbxA2m
ORodyDogqC3JsH6G//tFg2KTZvebaJormAPLFIB2lqfWY5w60Z6lVXZQPovxDHXe
jACvvFnW+hlb64hV8nDPa5aAKf30EoxY7YCWvCjiCPIK5hZFO0it2J6dJdGHXu9l
Yf8hba6cOaf2JsHNmWYTaDNkjaJYvHwWocIDZHua3+Wom0dTCntsGFKNzT2F2fx1
64YlYaMMVWKDps0kJJViRx7qKUrbKjYgPbrvpKS6lyAb+HZ8NVuspuwMX9/jHBew
VpBJxtNmA1IfaSSZ9WaY0aZXoIbGZqtU5T6NtbCDTXRPtvqes7suBvD/XoQvUWxd
T+YKPH2Vg7rIDZ22BW1Nkjt6wqm+zonwwV2CHu4I726eBqKEAw/LgXydIi0dYWTt
NdWOoXLRu7HM8xREUfnuSix8lDOUu67RxG/qNYravkrJwzXFNcoR314SQH7ix04O
cHqXtirBSNTrXhi6rua5xv9ANjnGZXoiZeE3nshoBtXxxpKuMFMNTkv2WGzTvUp3
bTOpw/7ABRN1RelC19EH1FyApQuL+0wRnYeRqEMHGgxpjIRQVWtg7i1UhJiqEWwP
yVEFAAzniAPFlNqPVZCeoH2SfECUyYVb9r5T+wxiXvUu3lOqvdCuZ4GIjTkEoSkx
3RHbO+WFZmnZJ6rNpTuRtFKgHpShi4JMNRlQXU/DWUnpGDJgh830DfmH+xkpRMtH
jjasJw0NMDPN3cM7o5IB5JIOMYQotUNg5dFjeA1g/z7eSyOibrSdRqTabDMMKvGZ
/OqpGrh6GF4ZTSt0lnjqxxC3l2MYZyg8669THNU/l5KYVom4sjaehlFgz6Q/Xmu9
CRe3a5iXvJi2K6SlbEOzlH/SgGgGnVeSDNwePBY6HgcM+NdxfvejOobg5S0P3tja
Ga9hmz7p5+oH9/8VwACxd6La7OoSVYpX/C80s3yCVATaqTxmQse8vttzTJfuZbCP
iDCHzKYQsJA6jwSHX9EJQxNhSc0Jkmu+ZAmyWmh+C7w0Zf9RqT8u2wd3l4qWyqhU
ml707AgAcH3pqdRXpHeYY7ZTBsaQjhmirL3uQNJSZU1ifYKcRh2dFkeKswZSXBAp
lYnlSjhW9FxNkLoPYQtSCjY6LaUJxAbQjt+ivTIkPc/DtTiS53Q3VebCWzhbRU+T
tqcGFeCQ0/Bi1UMHiBez62Fz0OvpQ2lW7CcjAAaN1K9q7UR4wiXQ1MiwWa5lmmwi
cyYxKEh0Tw9GlVJDE1chJROl3jfih0sP+QFNyxUF1Gv0BPwa3dIc5+UBvRyuiQiN
3CUkifxzJkTQlMDVvii6Fm0Ti2CkG5Q+G6iJw+k39zw3SMyV7cg7NLDIgY89g0l5
O3K5rTGElrq0jibpYXzZ3jwUxmANcx0U3EQnMuDhn2OzikZ0LhWEFv5zmn+VJ7MF
5p3KW1RlPlZh3rZVWabJ0gq/PE67PFBIHVncFYUxLRRBmxkM0YoMFdsa6DDwkjp/
Na17rGaxlGzoPB20MdVji/WIj5i+r8L5qGVI9uyvqvhsVo4PH97p2yWkTFZYVTT4
B0eKcoDPX20N+5Fx6nRvL9j2qqD+WVN/mlO9WrnAdEbVYlFkBQwnq51qmBGuwuSH
4yL6fdHxjeidOyRyL7EJkBYBSxQISKlac2/ONC85/R/iDG4arU7hs5/Ph0et99lC
IZYLuyW9OneXP3DVwpWy+xqLYU8KXDzHQQo5w/3P+wNU7tY8KesQPDNlty1pjA90
CAIBGQyLNsq4eLuy1+TNi8pYKAs4kgkltp5QRzStIvjL+4HXnXXxnYhJ98J2rtSO
JGECRC/MQtFOmSWxlCvk/0oLzpaAZEFcXkFTwUNLZQEcXr/HwdhPZAo7uehpO5+M
JmcI3GR4ap+pgIY208eQTUPToQqXhurQb8avtx7pFnrIFN8+W44fCHkYdd/FvkQH
luv8Ua01Cmri/rUQtipoHWqI9J/o/hI8MOFcdsT35tT+Xn4oywdP5yoRTeBDk+h5
NxZPNyzjZiuucOIGVdr9KM7Xz95q9XC5gUQUC3beTzl74ILEKcyqsjX+QCCiWaYu
Gw2J3wpFFjcX0XePdPF4AmCErBJEy6+yRVWtQ4y1ZuRM0HeA0lL1tIPm0Umox4oP
wiRdz0T+ILSxZUDh45eAEW3yqrsCmnD/vr/+nyaADi/hFkCKjhdfVntDlZt/VFGE
FjoKkFrVcmc9ptwnWIWExf5jfkDYWG9wbLIA8jIugVrD/XQqi/sW31owuzi7+51m
VWd6wKzTo2qWT9HpKCSQ24Uh1ZXm3SSqyFIagjYnkJRMyn+4pUxD+w19LnISUVg2
xM7/19YHObqjzwSQZAIhx7+Iog8MD42vqPs/gZ4s4aELBxM5i6TR9Hc2FgYiS5Fr
UvBABcPqxmasimZQ4aS8xZc5i4HIVE1OAz5XhsYntblQmFqoYSR39c2vRwTvU3sg
Ij76s8mRsoxfSXNZtK6pazQtCxHj7tVD2REuGNXT/r4m9A0WvnCwDAy1USBdBpQ2
eNNImQVucBCxuTxysxquVq6oCKtAyPbDyM85S/kZ/kyXDiuzSvvbStOCwJCWuMbk
DcGc+7fQ+OwDSUCxwLhis1cLTT7QpQEKL9gJnOHngFpb8KINe614P7mia9k01Imp
uILe4rXPgkySXtHMh9egW17baDZv9Ybqzhd8xtxipJG5GScXPgiT++wp/Uq5uimW
YKGdywn4jwpBqG3VC4F+bt1nqTwWRW78VEXQO5mwsHl5hkKfdDby+Edpf9Lmz34I
AEknpTrLWo1b3PwizGbybxZwWc/MQQw0rLZCDmbceI8Bja4dHqKqmUcVJSL6zvAX
1OPGkMehO/tQfg+Hd2F8j/NnI67FKom7/opmdljg4t8bsR0theXINhKzIiUOeGGK
iwpKT33ZBh9mokowtJwgHGfA1hZvDYQcVl6RvAT8R0EGZrICSBMKGC9QLS7xlWlw
PLKh//yF7tpoeLxFg+1HNeBtYhiEiTOWmf/j6suOG7vBIR26TH/ReP6keLueF+V1
HN+cRm2TKBccXsIXHTAFe+RHq6JUS55kKJ/pau0GxoxC3D6nBO9PSrZWT8lV04N4
XSpYFkvstxEpttGM2WwjUyGiZHCbQgtDmiT/p+JoKmqQL1wzQyE6JpRsAqgwglr6
p7rQRoEvVijiArCCNRpAAiqux5ON6jByd6duN4vPTyhDmi6TdQIVa5SrlEGHTL8n
TzDwzqU0TUn3hpE0ToETQWE5B2AxuOfAtAwp9cxO/xZCEdVZY1eDFyhMFNxZgZR2
mgp+tnZqEuXJJ5Z1rxcy6Zxia5ltANQRs4E40HzJFrzvypyRwRD9M6JpPC9VuBDH
sLmnHzZXxw7Nvt2WbjtbJr2Vc1dfB4dWTYQA2ojR8VdyOfy1uF4JvXA4YaGtTRDS
NUPl2dFtLLFUvUc78bN564IHiVykKT70MmdcfJ5NSes/FJpUPNAPsyS/SCBqYfsL
g5+Oyz8+QDl+DH8ccHyYQrwmUb63m/TAz+5lPLx1OHLJkF3X6r1zau3SeIuGyL62
eAg4PMf2MS0hzZ+3h9Em2bxOLrb5tNwo0P4TOYziJBIR8IdHgDY5PFo1QF2UbFwC
wzzP/1jUStIRDJ8KdfP1DXmPVSXOmTgRwEKoIeiOt1Hh+1/DPb6YcgrQ1Rd4Gi0b
tM/TSy8SuMBRXzuGO9Xi509sAtj0i9TW/JljCndEOGmuf8Ds+hSwWZ5bwAsGfJVa
TphwqGgEFN2BhYexWmSQhtG2Q0Q0EDDxSe9GgPPEZTVCR2GzOCAXDSlZCxV4lwPm
zWjVr8LVll6vwf8MmEWT8WlLNekFWR76D2WNzkfH5DmPyWrlHT1N2HyNuvdVoeBM
Hq8YSVqjhodvooEnmWfyp2aWDF83rEZfsDEO/0uwUCWfv/FCnGAEpc/avF42Q7ng
eBDCCGQIpD0M71rPACQJ6EfKaxIug6GyoBSs3/FPh9t8DDWQ3SyyrV6G7tGvF2Ys
T+LP978N5TmybmnqCEzG8QBp8ZMKouo43o8e4Twjd8bdypqUI7a6RhejuHr/0dgV
fw6gP7eUf+V7LL5KgsmdfHrPDLhiXUiVOggnHW7/co0iTrUwyQsl1Su1vjIruQEJ
LzSPaNHC5I/0g+yjep5Gw7WJSdAvVXlVL00BrW40HdB5+I5yD7WctEju2AWknLph
Gvfqu78hATMcW6bg5Vp2sVgHmPDElYv86zei24j9JeP7tl42/IOShyLO+X36diG7
Z2CGR4kgSSIlXWpPIA9y/eTxYd31Fk44FIPCa8PLlAOVi6tQWL22+4qrP/wAFPjO
AO6UlMIn8/BGNz6Vt6JICIYYXmcCmUM5QgdxSV5J1bilEgTf28H1bU0+JQQK1Nh7
UnS8mQOlIv77MuSOTcwpjGgva9CyjLaXqq65bt8+8xO2PtM+GA22T0sb7ozUSEoj
qDNBI6t/NBknS9g0VgVTy+2x/AAZGDGjy/EC008zUmJ0MXJOY/WHP3AnBy8uY6Ou
OKEoxDVULgeHqXBOLMR9yUGVf0GMU7cLlQzL5XrR5LDV3ixfmabnVOb3Hp/x6aWB
iyTsxCh1Dj7SYUYE9kfdWHvbIK6mESBAeT/Y+n3jKPB4RKGhtnWNB03sIMUSoUSp
t8WPExTD/QwDu8adlgQIWIZY1KLUrKQkAQo24WFUPtkrF1fh4psluy8XsanP0VFI
Eqknn1/aZYn9TyvR8h5GQrYCTCJFu0PMjH3sbRGQkYxmeM5rDJ2S+30VE+bJGU2c
RCoDTjxRwMQqlyWEWCuHRAti3S7U+k+mei1Fx7IjKTGoTh1oCTN+UtDUbdVdBrKx
fBfhvU/22vSAY4Bw9v1HSjBFFME0aRyM4AY/MajHPDGGq8b3t8JE/hIxduVjyfjY
7eZaaaV/1I8kVg+C/RNKa+8letZFOCpqavVtfOdzfJmhHVpFOelOnMBHgtlpgHS7
unGBfuRRKCju12NGphWnO1gVjIMI65YeWB/iYyGdQyv+FXC7BBrRfXhEWaJML6CP
MigFEiwgX4oNxPbj7koDaldRpJIMbTyTWMWdIccK6JiYzKJkN2ezPIyU/wqLE+e8
UaP7LTlskiZrJseuy2XoWs4L8b/jcLyEESaINRV8c26C45KV9xOyyevNholNZUHt
DPcFxO7y0K535mcQ0OttvguD1QhCdsVrDPVTp5Ro4x9HE0vWU96JOudmhswB+g7r
Z9TkrDGFCcBnt3Xg+iilouvBxXw7ewsA4sUtUKVXFMkab4ouvnmXXigMlnXCzBPC
qApoByZMvsxQFcZR+L1YfiUEhe/dnuvTdWkeYMJ/r5fR12hkUZchQbAlyVFZqvye
F5wTbsFJjq07tT7l5R+uX8sEUZDCTl7KwbdyCteUJdgxMwveSCdMMQop1MpPosZu
QsmyWhs1S1Bf9fnF5niiJIv6oHhPJU49HHywGyaN4pOttXuma9Zk2wVH6aNiKZL5
FouJpK5hUfbgcp45vgsnHpSRtHbhL0Jbp7xW8qGIMGRG9QTGWoXoe6MzQcW0rXuI
ouz9z7ypSJY6HQg3iHLtCqxyFmrKkJq9y0u1pCeQRrODgqkNqG/X5vAea7MFiCxN
Ygb2PnSvatZHOOHa8nzkeBqmfva4LpLHfBC0zKT/t6G6qnhH2CyZUtZ1BMJJYCEA
fcBeE5lHslJZnAucXHUpJhYjPPIsro192BF73JbTGSDKlVuxv+0dzer+e5ZAZIQM
F1lZmhuPiT1IJjm00B8Xb5CiPlhebCo0gS3F0I90THdMw+WTz6vXNV7bXNvbDD+f
5KAzauZCSTvW4PVirJ9D7MbhMXxPsuJoCRsFRgLECnZrvKgZOviafbpliJh9FPxV
hDaIT/kN5m+xSFSwVjh5ae9rbeHXwMylGQ2ErlZCFECGWlwIpECLdy63m8KTBrfj
wMEflzoW2q/+0p8y3gRPRIzP62QhG2SkS9SBgEiSJRP4ivdKa0V4Z388doeFsyT1
fMHyfkPV/okGeNcz7yj69NTJ4vb0V0A+WJ5gGXS0kZqTwRgW3ZF79UPWKsorYaRy
/KMQOi8e/OCpKh3G7x+DfW9H7a7mWjBNbKfmL2+QvV12uMIq442oqxVaSUj1EVQn
2bVr58mZ3chJ8duHdZFluH5N6BXNprA+j54wwidPS2Nh01al8maR3lcCUd+7sFfH
XwlkcO33iBp2fEQTYXGOuX2wV4mdpciPpWP/TwyDiBrf1ol3b+pVb7MPldFaaXQR
eWSUzR9fLgTeR//kzk3OrO0Qmr5X32p0lTh47c67QijYluV5IXUbRxVPFlhrBO8J
FYiSSR/v/UwOvbs1aZjjb7tnjQJJC/TGUI2fZaUOQ4xCXwGmTd7ax6cCyfoiqfxb
w06pvVlpbWU/8ieOCTEelCwN7iENpK41riqyRiMYclHnnxB84gAFk9d74+x9p17s
JpovE0YmZAI+ZgkEm5xeQku1yHE9Se7fvTltVJ2jaBkrgR3GeMygQ5+CWGbOYbxY
63xI4S4bvNLzKMFNeEJKzChgu3GLfN/uTIcG9PK74Rz8lyuYzBqwIaCOKoZI2WT7
PRmvE7hAMgUuH/PQ2scLNqWuwiUSOvmvoV+Sa2Sm6jBPTvNrsuuEjaHIeh2sn1GU
jNxoaxq7HeZR4fbMfTnR/Qhm22DZ4PtqPEcQIH7CEiSmCyY6p8dKI0U21i5H6hqa
ZYXsc4xRCXnJa/H08HtNuSXbLQD37349ClMMNNDaXyXrQA/UNuF71nkju0i4BPxb
wHoWCQQF3DyTD815n2k0pbQDAIwfNNgRzfoZXEnT8aPQwKRh3liFrXvvHMWktLg3
FNw1ssBE3qJ+Ds4SRJY4dqQf8APNtoTTA4x61+x/JsIfPi0BmsIITnRCVwzqa8Bt
NvC1BLQp4sLBCTGmtfZDJl+G7QnniNlh2hw3kTbeJRuZAghr3PtQrS3FP5ahvuWo
EjoCmWVd3KD95rLAxutO86DrPW6B2+JkxAWDWNepMH4jiqS40emKiz2KOqAMWje3
cGRQjx+2q57851PHtvavU9V78YPkohD5wVVwRrVvsi7Gd8R7VGeUVtk0pCBQTd6X
xHqOUmkkPMvYPeT61Rzk+gxdolOTVo1SgEFo0lj+AWzGk/53XWMcNt5Ia+bUo/W+
6aBAlUnTdr2c6oIYwCIMJ4t4oYBhF5LGHJ9n8/jSpzZTXAGAHQRboIkj3Ile5K4Y
jmnP4WsEYuZzHtwN08PbfOHA4DjFtIZCfv7A23lu5aklwsR1Bur8I8Qe1n5LhYCF
YR8hoXILw3K/+NjH66HHj/9kx6fIYN7TMwhtpYIScXBYXcTYy13ePbgJhj/3PfwX
JfDqRmyF5U87CuUIirJ6Lv6Fld6+RBis9c6EjuY1SK4djX2uG5XHBfHsYBt1mnj5
Z88fH/GkbMMaUN8d7eXr3rK6tJ9TP8hu9IA0Eac9BtvSVBhOcA6/cdQR/DYnAU3F
9RY+YGTLQh6V3hKThlEnqoQeY3KkbBXqzuLp3F7JNaTxISaCxgRnvcLUcbe/Zh/+
MCART8nLSF+rF5pg4Dm1AcytYugK2YlQdKQpx+iZvGwxlJ4z74BTNFNi+2r2jYZp
iXG7ygrjJZVYC2YeQSYs9gU7qUdlhxGQiQH9zr1QwQYAul1Y2/0SL212vafYsW9m
7oCIDzwiQsRvP6MG+/vQBmvytNCHW6IrTe3vNJN9K6aPbPsuq+HOBQVmdMR8wOGu
9AcZ0DZFWyHfbD5ECCjDzMPflWOhXeJraxZ5GKoa/Rt6p47yLzue8cZALy845P2T
pH7NrtqPHDB5OvQ6dAUd35mX8Tbk/bEzTKFaq5oS+pzjQ0P0WEUp/nDLGmrJzT+/
1D06fbdHLVojxiInTeTK63ajzJq6fXV5fD7wmCUHC7eljzqqby5JjNdMnCNHR+my
1FQuDeU2xWvbA7NrRuFl0D+6tpcjM7frscmjz3KeRWNi8ZrsHgejXRKLV3rVkUzo
hHSaNuUmxdKhtzkHAco7oCzJFnOmlI2x5vrtELR3RUgqi2CIIoJ42VIuOLYnDZ96
YWZahS2EEqa5XIKrfg4SohS/QwLWmtv+eOG7p+L3Pcg0ZD6ATT5Tr86eAA5Qu8wv
wX2cgvjpnE73G3a+doeUgDGuwuhVbdxYI2uMqv9aulJpdkq4RXNs7K2tLFZ/cbsm
fnUF0GMsRq1VzkYn2DP8FLNwXUqIHwGx5hQ0kyyhvixbU1rt+/y60hrFDHn4TeRT
nSZUCsG6sMsa3ADZEKDgZvAHt/2GVlAKjMUKGDmKHRgCwPGsi5ov7L9MrMdQoQMl
QRLT7VnSeZvLSsEyFs+Vx3KTXANuvmqdl590QKmvK7uKogAO8a7uW/yXybot+DFy
ANrMwR1fb3t6OvtZRE/cLyoZ+l91JwnXNsIEszrsMs0RZ80l1WEsBaWVoFTtpX0y
jnHbswKKnycmV7vVR+6EBGcR5JUARIhF+LzsN3Xbwt4Zrcvw2z3LR0e8KIrArSn6
uGZh3Fs7/M6Uht1m3idPjo9G0+l7UvKMGPjpNhYZ570Tq1hPpXjWL+P+qijQakHy
ZawhecKMJN/nmFSetSYREPyh7lJm/roy7yJ27Itpot8HfqHtY/jywOcNDvH/fkkn
VEp4nHQ3SLgIh9eI5wvPFVToup8OOIHN34niMwXb/yEAached+MpA0u55Gha5T+4
cs0+dqZHSV+Tgi9fAEk3hLJLsz/GT+GryiDTnucWm7w3CLgw/06jqNFXRk3kTw0A
WfjRxAzLSvkmsK9OThfrw2XIzV3yS82ffDxWUAYIuEyL3MkXtL0MbavFuZoDhjqt
0by8nj48OEgSRfALu1ufmLOn9GQFAQ/IXwLI0DYIYkB9TowVmud55BuIkxvE5ujR
q8/SaLEQkjRHDLbJ6NQRZmvzXhSsABKZacokdbpCwBsuIgi31jLS7mbOsQO4W/Ro
2F1iJUuY3lg706qcnKqqrlPfoLz2mrNRnL1ZczwYXUydsltVLhs+ANguQfI7RAfC
oToTPUp7ORpe3ejDElI36B1Z2lqPcgW5reWfFg1CkQ/qM/I/1IBxitKLJExE76F9
U4kRTZO6ipt15/oOznd6Z7ZtFK8bQFjfsipl/KXa7rHzMhmlbhdIM1IdXUmvfpvS
SRUQqmTPlxgfBxiCJ/U5FHpZ+5c60KFLbA7aJZO4tXYhUi23v56PUq/Bn+392aov
/foxAQkzpRyTzwoAXlO3Kj3hUd+GDMlBjNYjKk1+y9IKOPGK2CWnKXIcYc8u0w8L
jTK7xjCVid8zlMz6TVgMNAgtEyulEAnayvqTQabtkjTUCe//fA7ASoMwM3L3Ys+o
YWP2rRq7WnJKqTlIAtJMrbZ58LGeFlpA6p73llLtpZvJA/1z+Rt5pmG1Eph4ios/
b/QJRRyTwLUPopcEYg0xvwNl9jz3ETIiDT+EyXENw512RXiACiRTsMGtXPkClYo/
MK08brvoTvwXnr5ACkjFfyNQj0aXcN0CKJfvCnXJ0mdHFyddEkHZZj71p5k4eDEx
0Maxiuoap9yQLcLAsi2you+GKRsFwIQYBJk8oUvMvIiyrVr2+GLO60MBZD3P01kK
8vVDpxsnr3Igm3vCsFoIidPQFG2zAfzyBMnYZ0eBd8aMbDZKyGbYdDxx0jSs5J9I
kKjdjHC9I2lVvM24cG5crqE+5gh7Ry8EwAfPqDq7brH/7bZt9yzngzMOA28JWlZf
HBLvmfu/nFXLQ+/YD10ckp/2j0O1IbgobwX1EZt/nuoXz+CbTDjxg7H+ZtA1cNui
3WPw1vk6dHtGfdGYuxybJe87Fv5jmYC6vsbrjANcqz4bs1fwd3PbgSrp9ir1bMYr
DH+jzj1phf2WuI948Zkic4Y8Ns8e7rs/O9WNHb/sDg/CpL8Xoqq4MEAeR193nDLa
PhzL3fPOB3GubiNgf5PvsflDJZsfmmlrGQF1PCczGYD7Xrhk/p/fdk3atk0mCiXW
3u71B3HD+p6TG9tduXf7SPuTt2+cI4hqYqCzsgEYIm3AKZBYcJ7IdmzHDME17FDB
AJgNJJf3Hxy7VsW/jWT5UCe0VOR5lBRRxTeUdZKeh6OrQKaTg4Lfi1pY8adBGNxk
nW7QB8BnNDFBb8BRzlDzmPKqimB9u+RxfBgxkNFXOPIT6avIxBxOcJCPW1JZEcUi
82YmvejaB6BggX3hDJwoe1WcKXdxQ3egNE804c/syKIBsvbCFb8HX6vs3iV2cwDA
JFSdN5KuI+OHPQMgNm81t2hJUglMUEmjL8nM5Q//fASUIlofVfOtozEW94AAcynn
bk2rdSzkIgdp7nUr1/dmeYf+NwAWDvGSz+Wn9ofnaZdtqBfsr28XAKgisQn0fgz4
7KAc00v2Z2tfmr+2pwWwD8I5B9PoK6HfsJvA3OLd6mtSTYh0X28JUHfBNlnYmEY6
SwX0QQqJziAzX8/ChLif20aWEz4oO5kOLbSAvsqhJLCMvSJ0ZZh27b0KVS+UCmbX
gCKzbem8lX1EZQu7PLK1axXUDiX4sI034ZcTc3sD2C+2tqG6DoqmK8rq4D5rUuMG
MPysUtN+wRGIG/LQIAPpHx1QskR9jCN42D2uaXj1yTwDIGZLvBclwIcG4ibe/cET
S4EcB8X2WpQHD7SpsQUctxb9Op0QmN1+uo4MU9DgBNn51lCCzJfBmmnjyrCM+QVy
9+q5oU3uYA01f85ry2oGo0Bcr4/uJ/r6TBGoVuMHQ29Eg1E9w/xV+iO7Lq+k3EU1
KV2HDne0D4jw8nyoEE949Y5r90ub7ctcobGhUwSE+LH9EcF8HDWDaqhTcC4NHxfT
PbfdZ680S6vvh6Q+Q2ufmFn1jYwVGK3AU0/uaJIvwCX9dYnJFRrNS8krHh7FgtTA
MlfLvTnNXUrR3sPdb1LYwlT2jBZuodJN5STGRdHSXfDQ9HfDp2rOJ1tp0NcDxfN8
25zpRiQBrbHafDOHy3NRBttqVhfKRTJbqWG7X6RotKGnrNlFRbzhNKRuHCCt8rYK
W8kB0H0fFfIySDrwHQBa1g+xLQfeeXLsD1yWTwp2xi9MrPIS5QB5gGkUMRMyNOFd
S3Pv/9bTxy+4oVANQLKC8p6Bvs7RqaOmWBlWPuBoT0qgPiPZFiaH1xb0vW2Lvct8
ho5+qZYFJ+s9s9KB+i+zovxPlrDqye+yyDZw4HC9ZMLpg7Ubx3EBZthw1J2uNDyq
fBmIeTIRbw3alkcHi7Qk5Ca6OvXqlTlR+lA5eehWmodmfOTcyHhU74AXn6AiZSMc
0RyRy9rwC39JYpnzcdzGOv6oK253VT862mujgL+vaYaUONkfW3EUVvyRhRXAzW4o
QrL24Asznah1JR64zJtk8yKhitOi4TBujnlo9p7uvKnktvzzGF//BUnMHjtkO5AO
6zDivjOyyc6hPaSf5p6qMY0Om3QwpgRmTiZdecIdjiGDu2fsTdkgVV6uy5WJ57PU
EkjOLkdqO9bkRaGUAmyEUkMoECgbD8rPVSJTSplJxV1j25r93GvGRuDboxPPJszv
nipeZW4FC5lhB9pv+WMtD0sHZpQztGs1Y2GMf0i5Z2v/pB6ruA5fP3vvLMVNVvI9
1z/ea5yc9W811pxjLuDFMfGaNOy51x1VYCxsA5Y5SSTK6gPyAbbNtaBsD2y3753Q
hU4XAEkLMPg9rJD894XBCSs8oIU8FykaxyA4GZnr9U8UTcNZEiecxvEagJdLpEI8
kZT1wzl1hyXXZW+AZ344EyBILwGKco0wS9VyJwEWO2GaxVKyJKL3CHdupB+J+KhK
rKSi2Dip8NJJBg+Uc65Csc9sVioLCw95yyvgTyXIka8z2HIOp9qqtV/3xNlV1e+k
ZaGq9Pq3Jlgf9S9J0qAOexd52F8c/JCGMaRJqlCib4dzvmsjc+U4Z3rb4Xocy3Nn
0gP4XtD0yPlFfyWg/DUe3iiCJHf1UQq2nrXT3B8oe31UPCBz7aPKUkVm8TGZrm24
s/e96yf3S9TI/xH8jf1WOwJ2wh1s5je9ra+ryrsSYIwHpXD8hovoB1pBYy5UXHGH
m17hL+aiyNtjHXXw1761Nr2a72C+p98vbf+2p6cf/8+xXthjmmhPTA6wH/1zt52H
ihL0Aouz7PLLVeljKb7ne2DEEtvDqTsFeaNsPUPx13TVp1rIn+sYn82KuiM1k+v6
/YRkGgs8n6Sa/CFNmtAucAmhw+Zac9Fjp2yFO50/ay9V4J7td9E+Sqre1PmkFZCH
Err+8gdCfbajAgFJYjsL0n0hbn5kcCVoKa+vdhL/9foiRTfT2GBExRVqiMCD1Xew
BsOEcakVOuUnzg9EJrmJjFq226lBaVe2l2Tfw9m/f+Hfjzl7L0OG/eu5uv2vuWsv
D8Qkmo5hfhXtHdAJ5AQdS2RGl2ORgZBwQOpVCodrNIanCxhd34aZ6Rl7hsCoo0gV
fLBcuDj114aruMcn49YoM6btLCSTqYJoVoa+NMnnQTj04NBgBrSwrkzzA++nIbE+
w0qPey15p2IIJgF8NpKis2v8Khp/HFChyiMPeZX/9Znnc3kDGYepGpgQPz+N71Zx
650VTPy/bsNcu5geMGcKHdJ35VheuA6FodZ+u5jQrCXCusG2evZxHwauvZ4HtaYG
S8fRilGejNuflbY+U3Gt0nsxa91RF8CogqZNIinWPFtRaDV8XjsNRiKk8K3ev8el
0gcAsHBhaa/eKT6a7BzDNXKFl4sxZ1pj5zLsloUnOA+ROqScCWvpgK78E9laatZG
YvbwuYGLK5DKWsf343kJ7JdwO/chn0ynTsdZ6y5BopStastrR7r1SzAZ0I3wWll9
TUhC1iHnqSbtNt20Jd1tGlq1YIDWnsH+2X3IVJ3hsPd5GzYRnVga01LONFMhzlez
XLjDYocVHld4SzTjU4zLyIfvlhu0IqRkjG9bEPnrUmaWWrVsHq6n0iwlaHtuzlhF
jgFm+44Lng9QVNcNtTsB8E0G8YJCQuhL55Qz8zPppV3M/tjDc9XweWOayS02q0jU
AwOR8kPHlKbPnPJ9IqKE3d08uwAN6LG7zvTWLor4c/HNLCFIgUnHNMKZkgeHwe7r
x8CGi6hKUA/rgUkZP/swtR4CNBUtKPTbT5Ubc5nolyj0nYVosS6Ma/E/DDvdt1S/
vuGqOHbMJGxEXDKHgtmYoYBfGvrlKPW25NhdQ43vZ8QRB77mLrZ7Bqjr3RNbUblv
Kv2wsh+nFTM34jNkPaPsYXMIEGB6rv4tXWrzv66/D/qsjLCgV64a70j/uLQJOms3
vcTCuK3jp28qlVE06r8VUlx1iagTebdlnOwlqK0BBr79ljB2zXv5zwN/FbWSx2ne
EDfhUcgBFQDyoIGkvI9cs1HBH8xgjzrhfuTjqLYxIs/CcS7tYGAcHlR6etdGZbvt
rrNgC3troYEwj4rVDrNZ2VxkE/G2Uli9Len1hfHlVOmWGCeUUrirbMuW89/3GgIT
7PdTkLPnm+Fi8vVLnbbdrlboOF7bRVN4Gq2iv56Cn/q90ivQTQOxJZ9AqGEgwN9W
Y9+6pbsf91/Ke4cJbvQEfCdiUqcI73SJk7hSVIrSAwfc4cpig4TJJeUGyyOvZKPH
7ybGz1B9g22ozn+wnugHViHMbI0kLgvjEKXQt+bSgt/UitYc4Zlc1fSNL6ULkVUw
jFqVQbSzzOpi40b4CclNvi0yTmE+BCbWgIfKc2P24+RqSUxpz3f4A1pwiBwj8LMd
C+720+UP55PgYbZKNZx+QLnZMT6/KigzKioxCIaZuHFEKLJlFuBcMPb8Amg83dJy
nlEzIcFvXJ2StTlOrQ9z7UGwatoz1cqpIT96jj4JbSaZGlHsTXpDorgNB0ko0cmV
F8Upq13z4t4WjNhd4tuOaxSONz0HhpJJEF2owMA4MdO+3uP+Qp0K0cQF/jqy6sNW
H3bLqlMbWG2jCj44Ym3RG43VfPMOB5+OedO7lDpiQzUU0Sfw6rIMg/4xXKweN6FG
+5I0cpNRsWqRBGgl4EXUX1LH/pPb23dS8QE64bq6mJ4jnq8316NQnlq/cn1EieZL
FSTu6GwfAscA0kJAFWnTBjSJDuyhin5dS+Zt1PFIDwHpsHcw8hxmAbKzh8GqEm6C
wvEknEBimM993nmzUinG/ix4OkD+NFnq9M0tP2/Uvn9JosPhfCTfosRMQp5PDRT1
W8zG6fDr3jUqWTIyESAyHq9qNxIpI/OH7E3DXQpnLYCjWJC0RanAPlGMgs7YYkKG
eV/AINrnNC71kFipjvC+zp8NNAI4azJepB+Ekn2v0KITOvTmm/8BgjkFLZwRf3Pa
TuM0R200E2a5grTXfiCrDreMIJw0jjQJWTmuNO998AkToi7xT+Lda0dJQXceBo62
yuBgSz2tLJCITliExxu4L5C+nuvyF1TSS8c7gwqJigEWVAZv03eM5BNVnTlYPW20
/NcfTGBOjs8AG0k7jOa2QkCWHPteRUlw3HrqE7s3Bt593aqRL703B2F209wl4+BZ
Qylty7rJfxvvE80rqSLIENt+fl9vjQ+HZ8EQnjOVloWEg5WS5LfTOiDAiVyleWJx
jrapGoojxR5DrJ6FpNG3Yx4KMV2K6bVXV3X82SAYNWuDABhDAiw+bx/lfYsvrdzb
Js8tROaEN6skLNWePdB0m7GvIsqp7cYRX2kHVTZLKk7IHqby6tX3nobG8lI0P5GK

//pragma protect end_data_block
//pragma protect digest_block
y+Ufe+ZK3eyddFc9n+4k5q/OZKM=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+LmXl9Emmf1KyL6vpfqm34zlJcih5OTJ+gvmGJ1ziUHcUOVQKpcND6tzKTRAc8bv
8vzsFG19WQVA3iCVyo47T9EmGI9E1rey270hc9YLNvE7wXJFmeQnOAcEXryo12RJ
uwUYGoBoTarvwmdfdREfchaHpF2QjeGO8iu3Y57y1l2RfFQWRZiLjg==
//pragma protect end_key_block
//pragma protect digest_block
tXhaZZHvEe4b5U6EquojWYkDkKM=
//pragma protect end_digest_block
//pragma protect data_block
DubXnz42L6UHfB7/yYH11fRop6EiLd5IQkKaAAFoSF1Nv66c9p+MQXnIXtK+13lk
rXx+nSVfVA9boNg1UeSnTkLAa80ZNQZO2MK3sSsjM27mgzPxBc7WpFUs2icBZRm2
rqKBDhyYa1N/tAr+ZoNjw5fsN0jQ82h50zU/Wx5EZdWhTLZXKikfzxqq6LilyYko
rM89qmtPEXRRRcG+ungygxI62CJQzg3dwhHfSxiW2XC0kH+G++pqmOOVu7x3jQ9n
ANaG2J8yWpfwP6TQy9YAO1vvyzGrcI0rdxaCf4qSz0ASLnHhCEskRvlO/125WgiC
JmEUi9RYuqXN1f8vQKNSkss0+mbh9EXXXy1XY78PrXG3uSnoP7G34K4VR5LK3/Rl
9vhvhc0nvphq2d4Jv5s9lJi8H6AvCMgXDCoB9tqFe7zrszy2wGou7yphXnAR9sB0
VC3TaU9TZXzX5hEX4PE8+Rlfa5ztLgwcuQkktZIJbjlBDjygHI3A+FLSdqRajC5J
ZYsO77wmyyUy61EOLbFRJueR5vO2VAFHzCJwtf+MMhkp746J1TGNkXrezSOAx05f
VFfQiuHFpa5rgraRFe/jTUX1A/BGRnK6bzuZ416tyJHD8iuauB0hr4NRlEzubes2
oNbsHtvly1U+4gl3ues0mkL/S6J/SNFvdu6ox9UBbG7czq9XI2UvMdysqvZyQVlm
lqywjhESkmrONORC5u0wpeSM/GV0YmF7L6Unsx96TnKJXp/YF5rq1dFzYJTC+3Br
WLswZJqWk/B3qniEEtX6IPPDGcz5mUYqDOlCBECAgr4V90jhVs4Uqp9dxBfg5UOQ
iANdpzWmesAhXxeGqms6yhTD+NM5n54GA/v/duMZMU66zUA9P06DdNYnv8vLrSnJ
9splePuGw6+oMDZM1B06LjkWIiKNLuD3bh/sXiNVyPiEjTKK3gD6NeEEtn/pOUm5
+78Yfc0FV6EhpNdVRLk1CiBjrOtsepH7a2TU3udA2+gCIqKsTbmkyLBGewpQsPWc

//pragma protect end_data_block
//pragma protect digest_block
ciXUkv/PrcniZtGtVK/i+dbBqDA=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GZInSe4TkAIp09+vNmzNaywi0Ym3tnpl82YbTyoU8zBGlZdA+rtIyQZABo1hSrdl
2GEVp5Eu253NrKsF4zQEm8v2DTJzyYU4MRD1OpTmpNYMUaCXEDHEVws4SHel/lXo
nKdWRTcmVZPkpkV0+J8KPJj6TXc/cCjY05B6cNWKmLnqz6DSBYRPPw==
//pragma protect end_key_block
//pragma protect digest_block
rtFFd/ljo9EOLUkRPm7tNeu8GWA=
//pragma protect end_digest_block
//pragma protect data_block
fLTz5UqJNrLUNuutLYudgp2RQEXd7AWgETljr2SylKplZBF9n53iuAFYccmpRGRO
BZDEq0TNJ3FYTuDX+ykTnSX8XZ2xVVCHkUPlXvodCR34nqsKErx/YVq59N/XCju4
8cEnauepETz7/TkdVHSdRiNPixFYQ4dreiesT9ZrRB4uz2zNaBhyZlXEzgk+A7vh
ragDh0O7DY1KBQsRKOfgXeZGozFdY6xdiXwl2f/JSDWGum8gG6Q5L5hj/Jb1hYTR
GIfkg48VdDV5RMSHctzguKOqp6Nolv75SABs/Z0wY08i8n/owZL83ZXuiR1HkXEe
bAN0hRevXH1Ybco7Wq0v6ba8kLHadgwaa67LHElRIFelOQD3guIpcd+SS1dngURJ
P9lwcLmmGsa//Q2ntY3aNPKIB+4AUQsGJb7X3DwZR6xvYWVqes6Obf3m8NjUb4m2
zYFEwzCELrTkz+ayemY8ciVi2uqpIXK8e4oApin7CsewJyduN/GMkKyyVbNhY4cM
h7EwmQyATQSJRybOK5AnsjBNUy9VYArZc2jZHNt/4bITdkIX8xTrH+6lHo4Z69W+
ixl94ZzdS8DmCNisMlUY+8UnsddDKBYT4VDz3yLTGzU5U16SnvJHwXckihSPipX/
jG3cRLK4HcfkBSKtZr/W8IFMcFDmg4b4NyTknbeY5bPC31OmOR/3C9BgrrcLcL6+
qluiv8tfDqh+LE05C9AJDFlt+Dce7nnLDYmaXlR/ktPvxMlM3+T3wPis29xdbwpQ
RdvtWHRxYLlA5eZcQiJkXmb4ZDzQcQK3H0mnZX/gWcomJvE/W6RzwwdHw0+7Oeok
MLoB/GdT1JtN0hojqF35v98/qC/4X0BvNr7wGc/0pblTvvc+UVCtAev/mNccNO+p
NUR/j5ZCmU9iryF6cRAoxqPFlMXdf2Rny2H2ucp39mHGdw3rf3LvMifJPNCTuO7c
g+dznAwjwbN314KbNCWCCDk8qWf3GAEhGtsBABL/6gwo6xdFO3YLO2+736G6zy9F
GDBwhWZR+VRp1d9eivS9DR97bo5LzLWGwyRNHTxdDv4eF9N7dfroehBE110JgDbn
pFS0lQ8Zq3vBmjknY/ea4DSqe0sJCdoT2zMgz0oJ06T4So3Ugw/qdk61dx2cOUdt
NMkuEd3Wcj4aVbJGUYSmiln7ZtTk1NhWn+R8BkAsQvwDlFrga5Ni2pMEE4PqA8vc
R7cKFZIxayQ6I1A2KMiHfnD4ExW04qAoJ9UwFxjPWWuHc3zMlA75Rrei+bCPjTe3
NO+tm/1HQAhhi+KZQFwcOP/yIkc+MTSEHDeqkZJkXUT6qHe2gLFNfUdxP4EaayMH
NQDCVezvRVqBAmwYr9GPSTM4nV+kjDlH8hlUiyXaOIKNEvnS5EGUCBi/rNGLy5JW
X0zyqQGWNNrt0pRU9lkQruusMFWeoorO3CnhW5jtYEN0HZy6XUXYV28cwyqUiLRg
WzCHcxnkxZ6VN+mpEN5ZuEwDLoaOlkR8+XKknIhetM5ibv0Isl+f0q19Bu+pEzeg
kEQmNsOPOj5qPXSvZJ7kurskr7A4j3t93p+q86sDuauzYW8EWXrg/FfB/xAqzoXh
Ye7a98ieReW1GxAIa9y9Fh1fBMSvw2RfcagQwSy4gsTbhbGAUlxSYw3Yr9GCHE+U
0UViodUblNmQvT/Kbg5+QIh9V9Vw/gV7+qi+P1ZN6qXLZ/Ue47uEt1FVboPmAs01
acw76xJ4HiscDnblSAdg4PgMGuwN1bi6Ml0582VM4nYJzPgDpZwTwthL86vARFB0
ebttoloDRrGk/gxHdSR/kk6qBwGzE1LadUBNvBf16/0xqeywnGEzbv/FcZKLdn3m
55a4xA2L5LHS6DEwyYLFixyjwDX2Z0Rxc8Lt8hSCFFuEsSs8+6SWLsStz82LI71C
UEiAXWcIeexfDePW7lrniaaHvPAPAtnaOURepSOnFydcixLbWe6GYcrXCX/Boygm
NrkJHP6e2BKHq1M7UocjFy+kWESzIAYhm+0+vlMRmk2NAmBtuFJ0KypwouagyrxI
Ely+l7cgz+CgbQp1ubAR1ScDn/UD56hbaDw9DWwbTv35NGw15oQ8TAR33GRrRRxj
f8gLyDU6noECgu+0uRV7hRvunJd0u+yBvYOcSkx0fko8ZW4uKCpZaAG2UZLzBQqK
kWNyO5+PNNHfGFMbey6McjEQblWvss8lbw1dhjC+S9933CzhBvRY9PlEM8bqa9iO
aN3cJdqJeiwhc/jUcyq9Jr1o+4Vx9lzv/Kxm7ZeLxLXGs+YKkaoqAbSIJjdnuss2
esEYX+yDe0yc8HymiLIty/ckFlRh0ZQ1PvTX6Y5z5N9XDzq6MgH+oyI/tmX7zuyi
tIhY6xeaaX39YcxomgNDQvkxspqjvcxKbK2NDrbXylq1euxnbTC2J5uPa/ZgmyeY
WTkgTeRRH950JfIGYPzXuGZ6zuvZZzNme7xYceJejZHKPx40S9Rq8Dx0l8dkETe+
Wy1uEtN/hKbrbwlI+9C7kUDckZ69v70bwuYkooCBrHn05bo7q6Zj6gO3IEbugIHT
GMXDdM2gHEHQ+LwY3wnIFcu5shexNqIzpsLWmqDGr057YbLBdmEZz6UwN5JQ/q8U
RV1kvxnP3eJOAAWz4hpbiq0uM/wGAzFNcX1sz5PCRlKRP3vzd65MBl2p0r/c09YJ
LFowZyOha+mvlo0MKQVnyUY0qXh36VctIaRiyWuR9LJSJ4nbGwgmyYSenaeazJzQ
CVTLbWHB5Qs0MydoHVL9H9CqyHXO6wQlyEh37A/BrFLgs4ga6Y0kS3c2himZQ13m
sV/H34LoeYZ6R/PxyivPbVRhwzpFSc07BaFh3FLD8Xeh3WaXbxZz3wmnt+IrqnfU
j8MIujXL7aa2CmVG2qjXIIt3+eP4s/MqBx0J22dtRP8386Oc1w3CU6LYx5HrvzDd
hhuar4b7F/8QJS/bKUjAvfkCBQ6ogDCHO6OGTqs45C8IHdhjxnrsQkoGswf4JC9+
VtSzJoux0JdG8Thskr/i2HPXvKZ/+sO04bui4NeX3ZEoViDdN6m1GuCyynkZBAoR
C+GQ6Tp4KSkAsgtRiRJX6dTK2C/itwkJ/J+uDaAt0KWLWEskaxEd0h5GonpgZ8Ci
UKjiNRRmdlekH75fbiqhvc3RyQfkHfMdMWWp56vO3/gzPrTwmBU/CQV86WRIe9if
P5PwR6qxTLgrNlKK/cuZI8iXfnC/n3d1GI+nYftjefTCUySiPMed2qvGqSQevVSA
aDJBI+0fVQSXcF3LBgf7ysnmyf6Bcg2pZJy37pph3361lbh0dZd6XpU7Ed7AvWZ/
K63ZOkpbWHmHmwM5Lp1nlt8GWud4UhMKAZKuuRt0sbkrSfztIAydV7EqQ0oXnqN2
ruyWo+uywH263/x68cNffpVJcm5fYykV2LjmXY3fBORw0Q30J6AQ7CSVrHMJ2UTH
hXeGMT49qE48RyxoO380IrkVUJ25i/C9/KqeJJdAmim0bZ0U/JrYOWD0adR5Pc29
3KPm3vXpZJ38kwBT8xlxo+xVBry7oX8HgEOEr2d45dD7ahyAbuOwb+NezF6yQZQl
X82ogcU4JVj4q+jQ607Q1F7KkNMpMO6uGummoqZLPbsqVxyaOWKDZiwH+tHuoyLH
I1DIJcpVW+qk4dVh7LLbfgTzrnnhZb42/o0JkjRZDlcQ3ERPI1qVrVMfzh5qOPqY
FNITmisL+LCRBKP7uaJiQsPTDC83I4DTd378wzGhTYsbX5Ve7LZlfLqfrwAEGT6U
uLyv5r4KNI1J6PKJN+TV8+7QOEUUvmoV8veCLnRc/pdZB+v7TcFGclToYzxhl2UQ
c9Ww/rXntbCl0FABvkTRwTa8mRvL2n6v4mHu3FT9cJQOpXUzLVc100C2moYhv1WR
g4Kh1UguLz0SSVrUhDDGJEhqdgVtAG/jnqFEPVHPqNzYF3hhawxMWmdzFs/SkZ48
wFg6gcB5vNXM4cAs2gEzNHBc1Dg3rz17upzOWcLa9HNszWH5rtrWZGcVbfnn1uzn
6MZQ+CDHmNv0Wu7xVSCXrqP8tHU9B1GpJjA89O8bG1cbpbwUGwgYtFP9tvfPQtAB
H918MG4xm3m2Z5iOdny9ue/qyWMY6liE2Ln8yzLoC8kuEqc5qyjGC3bXSU9TNex7
8TMCpG6X1ah9CS0ndoLrPQudkhTyFvLhvArFrnS2FEh5IopqaSs6LJOxAQlV9toy
xTSm+GFx7BL5MpjKYY+raiE3Np4bjeeXIufy7OXLQEBCTmm3T2Hr9b31W8LddfPT
WcBQ2GoHWVilGQsQ/7H8sYlbtESWHiQIJh/49IabJu54ViGy7aRtI6MasOdwMbCt
PBzLNgBZgNCByUD19RaQqeaGG+ue7wMBlMZeK1LJQFKgxolve5LkqzKmsjoVoyKL
RQrmeSt/7GQ/GFw+nUDVcOEdD1QI/gIAUbTG7ea8oZJDeA5Ijw2XLdC+SMRyVGzv
JaEf0zQyNrXuWbf+Uh4C0/DdFf+G/Sn/uvxJWFrannZVVbrZk84Xi9WOKnzmhSts
8rJqvPvGO4ZbUdmDVOf2LCRsVDE0F7XxsM/zuc5uZ/eyHTjRx4Z0TR3g4kGQbaD8
zYB51jckpd+EjG9MRpIbS/jHtFpAGAQgumOj8As7VSsZDSmtJqfHdb4C/kGFtT55
c1lnJbYmw9ZVKUyUchbs+ij5/Wp7eBVUJ9mtPgtQh26Py+PBH/z5OxhUEBPRA9Ir
YSyg7zIHCx5MSwRe5xLWdfeOP2x1/t6SQDqv+uWght8hdUHf11WtBOjhnUNT+ZZz
/SMB0APNAesV7KC/YPoSRmWx3ZrjTUOF2SiSLDAkDARRl1Tynax8VLOAmT0pr3Ph
cR6NNSag1JwQg3KHzg/ItRmH6kt+pkBxxDQH0YDcBK8J9RZ677jUXQq05B70de4u
M0BCmkVYbzpVvbP2ky0BQvdcXzAoBF6p2zQ/8OcKI072k3h5BsxksTIFQgW6PiHX
tQiGSxAoOO8pTkuI0G+bl6Gzte4xEqawAzTzaEFGIEEp70VGaYbSPQ+FWk93xVhC
LbEOKCsBnEpuejb09REON38bt8Cqcdki0lsS8DEUBfyJul0I+DTRXrjBxkYo16aC
pPQbRplDf/LWHb0ld1KNIF8WzDX0DkiSsVAfZHJHskw+e3G6DquSPwNSFuWmK3po
9RIbSfFAfHkBrPXRWXbRaCUPldZ9I0Nm1SCOQ3pf4KmeYdEku8G8PHMalOlfw6wl
WL57UvgQKPrY8ldAfbqhhGIbPbd82VhMr1yinKHRFcE+3NOUEhSm4qwRoXJSEiX8
DeBk17LnTCYmyyLAtTF9UNs9Lsn0R1rYk1uiF6j3RZgYDNSPG1ZpWWxmOpODzhx+
knXsLvNY1FwvCNf8MLmvcYwNRoOKHR1u/e3/QFoFbbOjITEPzIKMYIFclWwLVl0x
2p/R3JFBHQX/nSQ1N2zcEGakMJdq6tzUGD4fDgDu2ZyrymrcOR10mMM559rxXMJj
jEcJU4f7h3p/rDp3DIG09zbmc+6hK9IM1Ye98Kp+ffg7xABKyWGor+W9Emx1Vt5W
3lhbW4sA7FnUzMID1OtjPY1uM3pIfS665wWbPgRueBHbutw7e/MpCsIBfmBbA4FU
hWPSp1Jne2It5HCTEk7q54XgTtI9OPzLHwnWvqQGz1NfazOb4IshF0YT4tK3mceJ
ljDUqopMcNFnH6ufzbBM04XF634GY2ckpsR50AVfW6urrt65KVgPllIQCHjglSo0
HKKK/vjWO1QQqcd7GfCuZ5waOLyW7NJkueBBKxtdRgruZka1U8sS5x50wSXpQPvx
iUr2KXbF+lJNCx2BhJPqpSelb5tlPjA9fm8qvEOLB/k8a9IEu8WSn67jr/wawzkg
AGjAHGbctEFZyIMchKVVUY8TSx2fT0dSHRvNvkq1zmxDZ3BAwyoblWYiTEkoSkyc
UgsJeCUgZkYhCPim+755EcDEE8/Rx8cIijudXyBfn2+/yTqxVqN6e356ZFNobAH3
khB+4FUne0QeYLVmJS/8y1K8t20oPEvcHUfRi32qHoAtFp7MNjXCrm3OMk0OBSfI
3ybdl0BhZMtLpjyC7FOsvcjfattq/fYJjto6V338VRokYnDPUDrUBxQ/opxNvQ18
8HS/lSeZfmn1q2quZC21OYAUOby4DiNiILyFM872D3J5a78fWr3YxtMi1gQX1K9L
GVAlg4qTgXnJmaUv1cHzNGvETKPTz78pPyOJmbjTwaFuG1KPX4b2roAIi9/gWg3V
kqfcrfS+Ke+dcqKCjPXWWlHAye2lCJ5LMtf4oBdm9iR74N0lLiJ5JkrXxWOblZ3A
vMcc7jjZcYoNV+ikx3kNEN28SUy5qPYVquv+rB1HfEXVYLBut7EhIIeMo7aOX/mf
/gm92ZIS4CKkP5vkvd9h65wPqcxdEswWH52fnt02rFFRX69GxdH4fVvn2pL1egIY
cCQi82wnyfVByHZ+XewjifY6ju7I2wTqJqFQCsbWOYYPKAFE5uR6jTfLjMnTg553
troSX24muLA+vdf7aLlcsTo78LGhG7Hug7qGqezrjdp+/3Y4dGeTFbfokmKBeMIB
yCH8vu43TVnha1nL8HzNxR7OTVidvc7pYypBhPLQfEqVDhqL0tLoEgeWPemCB9C2
c4XxkuUcGpZKPOhVb6dM0A+2QVVo7G5yEco/dUNMPGrXwptBG2B7MAflRZjscyLf
36NrzMSULFGIn1VquDxbSh2NgirWoginhOqBS2VuO0sY+/ZdsaC7MsHXdDBJGgkN
ixeTigR++aY3NceM4AE9Tuy23AspI3hBV0foCHlGF7ChWxlyqvVUmdAT4MZOMY6a
ZTBsreAitiYU+Qj5egfELw7oV8rHZkyROTzuLXl7Z/1Hah3WS92fXlyr7e9UlFVH
/ffBHWPZmG7SFoh7TsCZDJHCsGcTO4+rafvr76IA6rN710pJxMrbBS15FaRzyEdM
8wqI5wsx+F5nEfVUW89pKFnSLqruohVWW/ePeNP6HVbMSGs1GwHRtEdYQsRZdKFz
DeeRoY0pyVWzH9QvwM/uKj9JG6dIAZeghWMqOzALZypo3c4BS6QTnuzbL6VgaTob
GhGmlirjAlAghLLjZoBhcKF/RIX7mPpbbe7T1PmD4Kj/eWuMEVIklx/cbUI/ZeWx
nPHhInMjeK5FfDVq28fDL+cbtLKfzEKewGDe7h9mJkCUF3/D/rLlTmF1SLOqNVsz
X1DOgCo1CZ0RJUAgv85MBmSQRRL1uQS+PD6s/CNOc3o9FgSWxm9HbdFHWndYy2e5
ztXJibEKvSmx4WJtvS9JEHG+e9xB8MYqJQn4hkRHPF9kRLU5BpqcLj+3k6tIRuI5
thLOdAii9PPRTEe0T0Ts09459ereWXopLo4kRB3EJF8u1RsYHtcIKsBQbATWOmz+
+JIaWTasTzTojhYACNEggHvi+d2sCoJIAaVwuvj8v6oOVwevfFbouyGKnD/+u1J9
UUiYF4iZWMS6m12MiQK0nehjGOUGMPuBK1BPY7JyXLUvJeoBopheriAbAjD2dv3p
TXKyounX7dlhQmbQclpg4ZqocATVkO3BlpaQls3z2K5yWN7Zhmrm34bPL/C6/J87
+PH0aURAgFWIqms7JW/iDgEd8aXlr+1XAKZEDJlw3l4xtLrXFR/6V/+gZwNlGieC
T8UUKtpvR59EQ9Z/Kod5Qlx8G0aQlPving10+utEQak42/eUmjoTCqEN6NDKSsSU
CINv8U8fbytBut8e56DvVzC4xEXKdym4SeFS1oUdTZhz02vlRjzoJO8eiEaaTXaG
rB5b5mvg8zY7GcHTtJHEW1KIddkX9LePDSqMgBO/5ZDi2mPVKIEUdTmnuEIfFNbJ
NPgM4C1PBot6Bld69RLwQj9HtdckLroQVazevAMeJWWI4vmxdRKb+vc99FzJ8395
J9jhl6xpO9bpdEj9uGJ0tnlZd44o6oUbb93VKXOxr01D0PX0KnjgLqYgHhnrimQ6
NnnFsvpA/GVtavk6Ixx+QKNjOShPdOwNZQ0s4XadaRgyIsWDCUYjm6O0fLnjiEJt
1cycPgPkiLvoP5cqfcztKqkJsuj6g0QMzIn3VKcrzeLO5mJvAqJIawuONbHIPysl
m7Fcbi/88xJFQrf50NZPTE1r4eKR8jOI0AQUpaSzaySUPwj/aS8RcOnQiRLunqE7
4sbxHl577m0W2QVF98/PKOI1PESRHY4j22WXVA7q0eLCkTpZDe3e1AkSkADb5Vzf
dfUm9wspKrQXiNB7tZ05nDVDVVNko76O3NXc7wjoEYSkowK/ifDv8NCnVtHtScRT
W/xAsQofBSXhAhhMaPFWchHXGj3Q7vM6NAnoUipPO7iYvS0Rpqxz1z8x/9PgE+TZ
WR2Cv9C9EfQWpzamqAJ26p9LnpePIo1qelmwBf2pHqursgHsQ/ObYMaU7ZXDw0/z
tif5jnOtc/j59nS8fhjiWLde3f04PODjFiPC/IS0o7o92Y72QUPNgww7tFcV9F83
76UJsczEFv5jCuOeF8fkeC11m4gIy6t9iQNcM6MjYvPZ3XG7bhYTe+iuaN86V535
fz04NtSMxdi1vMEEZPEBPUV65qW5PkgL9oK4oGPKAIuzHBAty99M1fE+3QFN2N7v
KPjQ7qrZNjQIXcmD4PvWVO1K4RAWIlMasBB2RcjqSDQ/lqemT7rrj0PiNlH6jC5K
mua1PsVZv0caAaONYsrqFid80K5Bk8xi/LxlKIZfvqR1WGFFtKcV7RYDZKl+Wpc+
aeufJGWBrdlu737JsYIV2DUq3rPZai5L3fX9bW0xCxRSvsXaELWWwXkRg+JwRcB/
9sTKaBPNuZ/N15f6q4Hy2CumDMOH9ooxm4EQiWjVr3h9EWd4/sVJxfVsL6YmXCqw
88TsbCRWRymoSRjRUJqYzs34FEOudWaLfOyXgsopYcKRWoq6+PjTBw8dhO2eClLV
H16V2cGRYfFx9lPsOjQA8v5hIhHhe0cWnDRFJbzJjMtz9zu8XIQ1/J5oruOuRTl8
ItFp7q8xZiPJ14bO4RU3YPdlkKimdEufKAr6En5Pq8rlsZAoOONF57p1Fzco+Dvf
JTARehHMk34Mu4UtUIz+cehD8n87Yjt/SpM8X6ey4k7DmwbXMIK9Fmxt+IAuzpBw
SuUfMdOV55EV4vbgNu/B9kUeSM/QR6DRyo4fnqYOhLeFowu2egFiR81hpgrgoeLO
Qb3Y7axKtEiWCuTml6vlekMqN3yzV4OFJLucylzg9bpGOqyIPOdJSpzq/hhZWVwc
VIHbfJ34Zci3rAVhczaia5zzAwZhByvwie85kpizRQvGxylgepRblAzddp41A7wA
L6tg4JD01vNaanPt9L0epyk0pvI2fc8kr5aEuAWNClagGJBZwtHf7FNwfsWvfj5h
WqHp77hBlYFaS8QReUKcKJKaRBFpNBkKqeW+Dz1xaaDhvnXabHj8dLzl+I+jIMLr
iG9s3HQJ1dMTG5/CIFk6biHaN12ZEIhfHazYBh/4lqQf/RQJKN8OzdBvKBfcJQaB
nUydxdHcbwI+BhK/D2Gw5umhuk1zKIjlBgzI+GZnCTWMseD4bvv/tWQbVcIsreVb
wQ1Czb+pOwYQy8CKt8cefG3eF21jILkmhdQaLkmA35IEjU2Uk0mjcy89qxdjcM8N
gpb3fXQhrNAur/aXuJyrAQszRUNppE71/ao6SXGf71Th0TRHoIbbz2sosRTypnd9
h3seDJ69eQfytZiStfdEcuFd+i1/s1GWRv5jzQBeGyODBMEJ6Lml3KQMemZMVmwu
TDlFhYnuYHH2gyG9wXh9jpQZeWaS9PWpnj1n85AgNNi9jhksXiChcGeuyF/gY3Js
Rzqd7nCb2ABF8O2Ytj1gjtDiv+zuZqcwwIJFrrqX8y8fEd1Hihga5MJpC64KH+nQ
Lo1yzRJs74e4WYh9r1Smm66gIKxyOTqdlTE97wpQcve+QVeuc7eAw9BowdWJzNE6
riTrzvCpAjzOrS++3gJ9rCgRqLOW/B4MfwGRjPh4Ho8M2GAoU8MLmZvQXx8b07Cw
8G9o45isxs7yaE6AJAWQrCwTx7M/aHwmb+ZOfKz5Ra4rJlzaBjNF+D9vLnfj4F/Z
8YHKP0qtQw2ue16ZLpkW34oJyd6OtCv5wBv5QF/xIZBPfWLEqK/u98+mWaee8B5X
wk/1RSJi0EsJSjTQEagzUWtsrPNWLtvVhmTx96hmgjZNSCX3uKgYM7pm+WN8lGlT
6E7TIp8nkcs9wzI6Z7AdXJ7uw4YtFfF/tbemhuIy2/faiIpU2Fx4g0ml/tbDPkds
BrU+fM5cX/DcK3c+MjOqDB8c8Bsd662v6S/MQRT9krbPNjADo4ma6NXnYg8RmmPc
8oe33QId5Gi+FQjm/Xb700qlbL0Wq+0ofucjLwkncVw8Njf/3LiMZ/JB/bYr0ez0
TGrVgptuI1tP5yOkVoeQh6NgqdWFoAJF8696u0402Z88gPG1xOlShvIY/n2KwmJo
sVbBlOUtU9vQfwk4VxyGzxuTT0ueiK5c/35UCkDpfdMa4+PFVt6RXLQMpB1dLIUn
WjqcoccTAFbujfDBNiiABFwCkh96FUPbOxg9cWmAWiKKSXiHT4NfvFkExrVMHp3j
Oo+ERmM6w0XlryYAtRKg7cPet7g/ihhUbTiVl1NcCNYudV3E+xSrnqto78H0ckC1
zfyyLNmLv7Id3hIj5aIvs4eAafdMkgmIcyPXHai7tLyvo1g8dM1nCzdRVFaDydTY
xhJ+pF4vCF1LaKBV1ilaBKTqyeuJfZKUOQ7ZoxaBq+lClfpQMd3rW/91+2Qfhgqi
crkayG39lz696N8S1Q9t2DziKzb/V/y1lzNlOQ10zCw73GAUDIHpM5zx3IWs+MGZ
kKduU2bmmzqqoOxhoPlp4Oam47AV3DpGG/Y6svX7+CZmBUoaN6KAJT6YUvmlTrW2
iVoxI17EFXnON6DFh7Y7OoYoeGgkFWSGjlCTOQQRUgZavbuRYYnSMeLaEgflvhBu
nb+g7yVQB4u1XFDAQI70xYtdbh/KeK7GrBn0DXmod76yo601ih41clXCAsd5Qe7G
h9zpb/BDZETeTzM45BNYMJUATLcrV8VMhouscZTjV7guLmfUdbJ2o2T/d7fIhmgg
+kZPiTenszpPRf1bKgb7zOwDYhr5S3mvpSYv8REZWbEg3Im3OQyJInrF5uDCMh0g
01GTnpF+7ICmgwezyeWK0/ftz7xKiqlDGKWhYlbnk72ypnVYsGzsPDEohecmR+OE
j3uY4xAMcJ0O+0t+wn2QVRN0G6/CvgAWRUPCr373AegAlKtfKyxD2WV6EQDF8OcJ
AAEr0pbJ6b5mU591U6PvYJU7K6lh1yXSNV5xRzOnb2z/url/vBHrlNAp6dGadY7e
60f7CqjHB75JLwOlMxJp2LPYIuWfMPWQjimrQmqrNuTMN1EWJnqFWn6h+RcfZxts
MKgWHOguCAMi0S85zJv4K4KE+pMfmoe6eVVBh3vOBSqu/lxRxvIbfwDs+Ve8sfcd
dIwd2qtnuT6g7juYuZ6f0N6AZXf7Pya9XpdDEv/JA6roIkb6UT5TwujAMOMZQs6l
npb75xLXpaYR9NKV8lTb7goWtFgu22TV4kqvZEd6/creDtpR8OpC9bNHvMBqWxY3
AHIscF2yZP3bQOBVerDtkdUsClSnmslI443FHp0LAPzg14UOJ72CQhMVJZs1Ieho
zKZ8rt6u8qWk+BEKf68Ib0Vn5q7CDz+WtmfGYjE3cXugu8rt8bTWF6ACXRUvVLPm
7c/qMATkM/IkdZ/MjENM8MWaprWK+Tdowi+Z+/4RuCcY089UBpwAjmLLXShWhZuO
EP9ynuAUGCUBE5ORsTCY6NVRcql9Bq4aYb0I2MsQYlYiKhmNEcXbz6XCRNEQtk73
KHp7dmsm1QAiiU3SEWwMS7VZHNqbGzMEJavx9BOWPvVOw/fF4nsQO+lX7xIJlnhM
k3lY4lZhOh5aoueeJ68hBhL8C6pXq+tp7flD4w3gQJZJQDNQBbdneWr9dzT/tuMl
ajN2sIVaI+Pm7m6h3Ikk+Ak0dfc3UNGWEzQ6nI2xrckeeEDHaFlbK2wK0x2ePGAn
xaoyDBOB/gI7k66H3DDCKk9siEFXvYAMr9LtSxB/DCDp3hCHR6mQ687qPlRnNbvs
AmClR8wPDYtuU/DnoMAi7ywBfgxrSsn4Q5d54uo/TwFKqgXy5IQEoyxMuO59QBJ5
22p7Pzczel0heAa7BRUF5zTlyS2VHF4nBPzv0Ym63ye0eBNJ5Bl+2ySPqNy05pxY
rsYTzx+QvBkVCqLeq0mW7wy8stAUU0U1CcB78k5MVmd2SzU94CWFj4nFDv7gbY1v
XHZoYcTReqycF5UipWpEhoBu/6bxPa529YwwtwYHep1jzkio1k7zY2w9/F4qd9Op
qlZzW3sZ5m/3SqIk4vVlBVvApUxwkxRBXBAhRm29jxfj1mMN+inwjoW2DrcnL1+9
bnqZFwWEkOVxtaWmwQX6HUSf8f2Y+Ti3c+gaeP+RxlT7sukgJlM2RvoRnYETCGRa
7HWgndQmkctv9QN04YML9Yk8yLsAhaiZvgpNZZ35wJYqoYlfWgx8Q/zvSvaXEaVO
2jl0Slie7Zsnr+VcoEjqjrWkcVNNcQFQ16brkfc+cxwVa/eGB1mgxd3xKdzQtRtY
9Miyf3JbGcWZ+vwyPFVyKdK5pOKGHKTlefuMaViubTUQ+cN+6RFYtuRWgLlKAj5s
OuldyjqzUQQIiZT3x0io3qcX6NGbToxuTM4Aqe9tYjLeD67B9ibAFjMA95QJKXnY
5XMjkXHgWJp9/n9952Mq90kU2kl3/ltCtGUp7JqY/k86eRZs36ntXSWdes/QoXWZ
u9tzSpEFxlqWmWAVAxDRM/57hJMs37hXnSrflDpNT5QlMS2H3ObnuUChyXVfiG8U
AC6pIDSsFlOm9uWKQ7ZQuFTlp5N770bXQvcxoz9ADDH9+ryk6mzL8gfp7/QTKBWO
bmiv1IK1WkmDt1o6bh3KGA4XlR4ahzVu/v1nW0n8nNQI4MPok4bf//fQt2i1a5t8
oLWzWy4G3UnoWP9JDNBNVk87i1t6z7Ctxt5PF8Qxgb6IUZHeQcHzPu8vE6EiBiw+
Nyqo3zJmhU4BqPc3VbGUUiTejckSI5pFddVfiH/nOnfjrM8tstss+pp2b+AtU7/q
S5cAC2ZTO+B5pBukStzs9fVYsQAcFhOq9CFpWLbD5lssbv2G6BVEcIWbMYFJFm+b
SMNi4oLNuusTg3n8xWWnFNaGY3eKyqZISupG0Ge9LYThheEe5MEttopM0EyAgq0o
8hc5v7Lo/E6NpjUPWlF7cUPK5xJfcJhZFAVY0aNxo7lWuSodKwIwe1Hd+Y/GtcSS
BRalXMpQ0gFru0vfJQH8OqLjnCagpuozGbSQxGZY80WKQnYoP/G0SYxNua8ty3rQ
10GQ5VCjaPJ43LSeToJC9pCXEh9xTrrFpzQJC8SGOI8CyBrhXf06ZLXn62xTeFTv
7kf9Dgvqfus379Y3Kk9OL0beSU8gb1hsPCH2ENsW4gN0xVvLRv0sQM0BKuscMts3
VY42pWcVnxOfABXNyMzmhE4ni3w+6farN3CWpekjT6Os0JkqO5O/SqMR2uQeU9ny
qqqMnh61R/0n0eU1iXst8J5RjQy+iqmuDIUUJ/OA05NrLhjjsCOZDwrhrEt9mu0F
ItMwUgXrOD6Ind0WdIJmo6cPqaLmHcVPs3gR2Scakue51fgPM4G4+ON/SgOf0vUU
B7bev0lP4bSaMaizfaJGrImVJJpExQm7Q77hHSDVm7qErcpTrIfebGuIUuhM2aG+
yp21TOgqaEsH77wfBuYR9/cD+84AJdk9vxKA1fObwgwsfScipbnj8qE+0bXH/GXz
suvb/3z3CcI7sYC048ceICdkn35lUbYVcjQF4xyyJpxSpIXgpxMlrizNpa1mOajV
rfXL9QvrWyzjkRaditJxEy70eUwWJKdUBCPC2V56ofgGPbfOt9FpCiltCE3sf1nR
mI1/fWtyy3YeKHTtlGV49oVF3YvLCTuu5PKxsTKceekM4ha2qWtXlEmuz5QWhVOv
Chn+X6I72l997WucWBbUK584VBUpNgawkc9k2nA/sPYd/wIvNz7bOdCdSHOfN5n8
4uk+xcOqscRdc4xx0jjL64LvNJKVGwz/A0QLKz/kdva+tr5g/Um9Kcu43BKAX00C
ui+WVIaP0gw0dHxva/QnkIZxeyECXbNtOmUeB7fyTJuyrDZliCqK9fTMluaN2nGX
Qt0jb7152aWuSpk4R8ePE4smQufEt+gZ2s07i3mkeKn8AOyY4SbjWHgZ37cZdYa3
uVWXAsAdJnlxZfS908me7svNPgtDVbxG9SPuHOk+hqwbVCuYETBlkQfHg6DElFgn
Qqiw+FvGVVTSTQpYz4KBt4qO/sjLspX71J1qus3W/q9oE0/rpgJSVpnWMSEtfWyH
XU6Jc5x+JWLO6rwE/nHHq+0opAlfKNZ0+Obq1S8CFag6FkwgjtsHeJoMr5XYyF39
MpDK2rFswyIeTYE5kRk+zMwD7fpOiXpbzRlpJYFLkA7T9SPcqRc2cqxZ1Lik22lT
mPpWRFZC5V+KOCQGuSjQczX2nMH1SgwqC0O0r7dpC5s4zxJLw3GFVYmsbZbGg6aV
H98lCyTVABZscsfZlIEh52+E0wcA8tBeVkk3mHHsR5xvIMGWRnBg2Okp+XY97fdz
y3Q9Y4CvemsoRmePq4s13KgEsA0vbI91cdhH102a1fFYvdxAA3C3D94ObsDKCXnw
/uCzR/4RUKBgmDSssDpmaWg+/jhhKt8Wn8H9zFjp6dlWv53MwIvkSzjvxHdVGbjo
gQVDH/J6Fk97B1941MpyTlua7tyaVtw27KTqz5QoIpgSleDlQha/JZqlNdFGNrJC
wxhPXUghE8J+JrUvn0lqZ/R0Mk0fPEmjJ3U6CxwgeFv1B9CY1e4xmlNGRWGW092g
bWVKUKH+8YHcCzn45xhGPd25EzWK090RaptqOYs4rz80+4KIynlFUSjr4QozzuoY
PbTeFt+aFrDu6YmtumzVgEjtNyip8CZ4rtJurlCHeefU83Lkz+QJNVEqavVKA3ib
xB7CzAj9Rr7vW1NFmHdrMEFNa56SCH9h5kAnDW4CLLSaGSAZxwRD4HIPs09PMdOn
3ltd1vU28EDH2IddrSDZl69k1QQBdD9TAPRPOSt4xXDK32Ev5/roK5jnX/DJzMw2
R8V4YmeVDK+Pin9L+vdHwdnbNJWHHCYlJOR1UJfsfaRcElRDn5o8ifVPwsrbnueT
SVuf6+/j+9mTXqe4MzhZS8DEQzq21+G3Aygw0/aKRAyVAadYM0FewdfgIOLJ6T7Z
+kbeOCosMfKQgXfqKm8oYJP1CbB8tsntFaoOn57/salT4Yvcy5LkNcwSvlgxiGet
FnW0cSuCqmk66O5pnZIOdRK/bY5q3Hr0XBJi9zBn+wDB5fDEUdnc1OW+octwwfyt
4F54/kAf5P4MDF6CAQqDKPTwtnqkcgYRXxK6CaGUtqr4oTjdiBy5Ox7x8XUcSWIp
Wz7DgZrtMSSoE2zT1/YJn3uWLMr456PFn0nvwJTMTC4GhMRKZq3tHSW8cXRSBAMQ
0dJyKkvbHpkJNFpxCqA/QpkY9ZJI+ttIVvm3GJNZeo1uuMPlRlAOvtYF8RuuqgEL
OuOv3BMerIwQYb4JuxrAqaI8eYL32zEmnxR85+wKB9cxrW4Pmm+E/khyet7fGAvq
vnYOTDLJZWue6GKFwZ7oflXIk2JnZpzx88qgGiaZzbzAHzlJ4w1FfvXxAwCmZx6X
btB+MK1inblVfZ6tlPfoITKhD9bwSQ/lAP0pH1b+OTyJ/VK4ePmhOQSN7r4v4Shj
Cr8vNG+YWvQtnwHhozRjfxXIGdiRk3YKcE1LQG009tE8jbrnUJGHrW/fTl7y82KK
ytkvDhTg+5TiruZqzKvDmi3QKEGMBPYlf/uYamYxUpH4up+CKaGAIjoTxR5p48QL
tafPl4mrEgsqOnD6CX2yl5GeavTTKgIsgSK4LYJu7Qr2r/vDaTLK3zDnlut339ti
2uNPNwhmSlX5F6BmnX5x6aLZ3fw0OK4lBZA5YjX6HEoh5H5FSVvA2ZTFSCL3rxK/
hgDbqKX0a4AcUKP6HwEZhIbYL8LX4bZEVotyG5RQ6BX6+rSHwd1SYA38U7uiv6M4
aPeFlrrgL8bdezhZ6WA7AmANOZurU8l3pqvAxqz2OfBJ69JWX2p2YbcC5HEHU2Vd
6whv4kd+OyXFQt53niuK8H01mSH4BDKo01kw0h25U2MmurMcGolWw/G0Gflqf+4b
jNJaDfytvshzQnoK2ON21b9extpUQXISCZt80gK+2ddK0HIMpAVHP+MdqyhMvvuC
n/QlHdsfuQ69hfV5EIliHW0SaO0EGPf6grd7dIrj3asI26RgVZdfaCB7AAGqRpCN
skaUoiz0gh3QMi1It+0e2HRl4hQZM8CqvptWxYKNnb6mjPbqlOcyjzsP2cvh6Bux
Jbl7uevwnIZQTWec67qcjfa/8Kh7c0VStlzEtKp54FDiTaFXROAm8aQSVC+GMiYU
OEKvdx0bd9xHK0JJqmbuIWjCytJC4OqrLECs4D3tb7mwShSu8l8trl46n17D9ohH
CWeVvnFzKL0NaIMMc7a/ByedBXKUMQ6VxkXAXZaRlZu7NwbhYZE63z4p6zK8WROv
mN+GUORphGmjW4OyPB1QkihHMl6Ov4bk/79BuKi/RkcQf4UVZ38oDTmDoxgAOIjr
QAhHwoP21YOYiyieTmu+h/AGYB6siyzIi4y7kSylJoX74WI83QqI8BOe+g6etNHO
fqFWRpBvHFSYGmI+H7ah6mpbC6sZaIsNkFYXASPvdE/7dlAQH6l9x3uMQuf9hUUS
3omnhoKw63aOG3I8GdnIdKNPBX8PKSwvQqs/VFNwBMvmqB9T38CST906HITNSQoG
YAxzHLVg7QCVnHSdh3mw0oTEWpIWJ3rKlRSEbFhnMr21Bcf6XRVN1R8WpLO/cbu9
CArqCwbUoBa0B9C3Lfxa8Q1nYvrrf69KBPO1Gp39IgnoFypvuxLGqgsH1t/JDE5j
MOfPkM3B8VdOiYGnj93v6TxDkYRZvHulRlfOVpIpKjRljnL3Vx+QmODtbZeJsaKV
8EbQd1tfdTykrLAHg/+pPU/spoycOZcsS/ueQtr6hVnSviCbx/wvjih54Bs3ZO6P
wRk8v/iTzrDcV8AtTEnXQghlD7xIUd0GpllXj9iKx789sak7FAwVIeEGZlb+cYux
WU7CBhOVETLNq4uYbwiPjcp6MP4vk/iH5vb3nigxDUgGiakMjIisqMhWuKm/Wt2P
lJ6jywhuh6Ogd5aCKwIaoYqoAl2UbAuZ0rx3QiUPfeNdN7NjlMAVXlzPC8kG2U95
PJrbwOQFco4eaLfk2cn++al6rl6i5yRjezc4CNFzVxnz/QoncB8GJ07Hl//2lXn3
83G0c1s4RP3r/JiWPArOpGE+oEjWtwPHO3Ue8RbmuzZ4ySBppZtl+qyu5FnnOFJd
Z1o+6e8+D/qlzpwkqyxNYzEYUij+xwKBPWGIz58GahDobl5Uur97dTGaQjDVelDP
72JwS5iIPLiK+g4IzVc2ye2ZhX/C5Q7Kfo9TlCw01BZg2UWYORfOt7U7/+KlgXWp
hG+YWF9HDY+YHTMRKXvWWo4Yl32/PwnuJsrm6Z9TzN5CeZfEqq5C/M9vL9qaL5R4
WM7DmoSdGxRMK0TzmZuGSkun848RlgBGwEtjb/t0xWKOI7tdUd+l5VplDo9s2G5L
0sUTes+Rm+XdXdSpCaIvMinufZwpH529bFaJZcsMJ5j8UzgYYVEf6egqihWqE3/c
D1egG/TCGRt2IR9js9kDo5v5tS/vlPQLhyZtIGPzR/FPbH3ShStGYEPbgUDVPQHl
v7mZceibUFjJG8UZ4XdFwH39lfXZ8xs+arcdtqPl2HF7d9R7FSoIUFBFUAbGojnC
dcCxKacE2qcbazSkhBuFqITYBHo+1HQJ+n3xcc11aJpPXfL/YQNb7uPAlwlMYpF1
ReGnQXZFn90qMHs30kPq0vuZ157ueJkqco4bM8/ltUberCstKvcT8lvnjrd0FmtW
BVBog3fjSwhSKzQw1qub9/imOGVSzpDPKND+3+W6tqipmj0v7LU69EaBK8sHysWX
xPq1O4Yc4kpgLpXAw88cdOF2PdyHsZ0HxIAfR/r++UeqgmgPZt1wqngVm6hYI2HZ
EZ0yixv59BV4V0yzNetmAc7M465RpmdGbUB4feGuxjLr4uDk3mjOO2lqPWpdepmV
f+XJsmRUVXhGmWiE9+Ds/Tmee7HTMJp4Y8fKEMCUWN1W6qPvnMFfRtaxRyIq4UGf
yHZOSy5E51Id6qNwgrCdtQdPYC8fxvOG81ELrkidYp3r7BgU6EromJ/3IMBTPCzf
PGRCb3R2sEaGPHKqsaK2jh84IjzieXp+bBIaYsouTwstSvoadO+0eILKQHXqee6z
kW7BxN50621/DBYzsXGUDYhsAec8X8iwsrX2znOxkGdxoeWptkjf+MQoaX4WwR73
ylvTPTt2+HqAhyZrf9GE7n6N7nIXUv0gd2yk6w6Trg0Pl5MuUSe1CXbG8hBezejA
1bmnJ1d7PCfNrAqKFWoZgIksOvWJoa8+bXErwFwiScpAQf8SsGfLVyiZkn/5E4Pb
Fuv8WZy68TJojr3R0vxAziiLNoaaempXuHXeBVPquYzjnLnmqKKM2HQU03aIBmqU
hLHAboTilpuaaq541ZI0WLBkSXh3xENE06nRxTuS8tJ7s5pdvtAzh+nbI7Q2c54+
MSl9ibYcaLKhI6NnU3gGTw4cD/tu71k4segDhBsej/sn+cKSuJK3x7oRVHyMTY3R
KKodDlLeLb4ByyG6p5SiiCbTHZAILI+l3hLECkhKVwf54MdShMTs2RzIui/bKehR
XZJwYJoqOVoQKQzCMoy+ZTbrVEmJxh+aXjpe1zG7Pdlcl8n+1ozvgn56kTtBdVdB
n83BhI49VV5rGr3Kl2AAlDp7W9lrPjVa67RZ+CKDyKNY7b99dsFJGU2yi8uNSmDn
eWUe7UtjRJNjl37azOJ1gDzlZJ6v9O4Xm0Mr/iTqO9DspVnSrLLLj1eSUxZ/+9Al
i2ly7/dDbYps/nWwvSxUbaPNxA9Appj/IX14bRJasXYYX7217/8rUPEhEqsafCNd
cJ80O42b5TVw5DNFinVJvJDSEZZC8K73fSk2OGyf6zb4rMltzN54rtxc5/ABhg7g
dE4hHCIdnaAAsON4H2TWeqkTQMkO9b6QctAyVg9MlD6k76C/jKA7XaC55OeMdHFq
9pzjQbeRoUWLeZlPyZKrkh2ltXoMty+RUVu5GBZOXtMvvw0/l5nTFh8QRh9IBGvy
ihZU3haiKZoMC2f+5VNFFeTuke1t8zzRUtMHc7dcw8dem93U+rg3dWcnSTUCBcXf
gcMPMXCTe5skV7rloSOuVPldXiYwYtPY9zvR9Zn090s2BdXB8EWOH1K2g4VrcahO
nHHTBF2O1hz24VpIskl5EyY4IzQC00siaPAdAIt1bEIc6XGs6ITAGkil/BrWcs9H
2S6yHdh+jwzoYyVNvwa6GmcckvuGXryYmvWlnXGJSo7yqzMjqTxr+xRUasnjqQFl
9Jatc7Ku+U4bf6FL/6ZdPz9SQvkEOPwGETR5TpQb4vrnaQohp+Vl/aJHi6bHBGHT
syUs7ukAeDNyCEOHeHMNZAV9uQS5Bm5tEjNwH8SASFjbBwDAuu6tJXItgYLEhrZz
LSpoSVnaiP/YXmeHIalWMvLYDZJfrKC/9wFDmtDWsxCBuhgJVIKh7emT2gLLUjF+
gxv59nhAAqVm9Cl7S0SmI/s5tvtj7rYIb4ZCxQk0FT+gsPqwxAwzh08xVJJiMYIQ
mvv0IWGlzEzJJLIP5mI+YY2Xn1yIIgDsDBUayapb21SH2PMDgofHzviq9v6RQ/z7
+k8Av1SpgsMdtvjlsjpbcIHO1X2tr7u/CS7kp7b2nXYOdixoMqbaxLKrIK7E1ewH
y5ACDi4aLiHD5c0sVFv/X4sJ1SA9jLkFjhiRbEDxRcqFn4S+D/6tQCIH72KXHsEr
VzdKsbYiJnI6RD8h4KF4REk4hMkAPA7yT6uBs5rxC4/HpKu46jmqkNwCw1JT6ID5
2QCJLDXaVRFYllaMsXEWqYK6jVe+QpDBFsbkzLcWRVCCltrj7n+GXVPzgDmpC6AJ
wkz1zH3wQZxbv65eZtUAgmD/2V5JyV8zJk1VQxYO+vQvPwzY5jhpSbTHPiVK5QXi
+ylw/ib9IeECp6p6Jk+lS6tgs71Bo+yZgTetNL0fY0l0xnswxiILfu69tmsQRHHz
0O5bxhYyXGHPaPceHrOECTq6kFDJFFZ0HkFP7VgsMUGwaTnSAi1JyS4bS92CBLUy
Kg7qJHxjy0kFayIeDF68+vyaCZXpHRgo5wObLCGsOevsTsjS1VNiQKV/dlsyXSTB
UEuBKb70kPJZlqW/gEEh47ZxrBr190+BlsGPg93p3As+u6zj5OVwWl7YKZkOdPNO
G+KcG3GRxUHg+0qvpelxngUTxqnLf4obPKQxePtXmhEte/x9+3Q/acBampcZJaMA
XxvJwywr/8G7VUaeYgEyaYRV0PtGAWNZwlS70x55B90sNzBbsJearkda70EeC7eR
TKG7GaBgnTCMwsQWJUzq/ZVOAeGso2OPpy6RgCKgvVfZrmUH8Cvxk2STo5eIK8O1
hBnZ42j5Kl1oyoTtoHJebR3Eb+TETaLZpUgGt5IJ+Ppsw9gJg5i9SM4GNhGd771d
vANLyMIQEnrv4ktQ4eYQ/kvVDkC4GJB7kAkBpz0xMdlrgCUyJPh2nLfEZ7fgTzpd
7gc1pWgcPTcDPwhLSRQUdng+khE61f4z2KLTDB8VxEtwutUvZYJeMQSCs4EDqpog
OO9MlWNMaxrYgl+l3qr9WBiIXN2uAkEAEgIoDqxrjdlfiwFCezCLvuNMATG1RH7w
tpu4XX8PSxcjqegTuJ0rRCDCbw5aaxrQX0PrbZYa90GLS5EuksOq1ly4OvRCm2Pg
Fut6wzsJ/5OoZPxVq7yibF9ei0LHuQ5ZiuGGa0pCexIuJuDGK46rkzooBxBU0adq
VsQmryIVectYCJrGbwR+MtUrS2yy90S1QVvtwfFBPjaIpCeu+WntjG981RyCI57O
LpJ9iE1gHsyD9M5xVyhEvakAtaV/fy2TMdw5HGasqkH0ZAo4CbSdiHSTlxE4LYSA
pAwaLz7Hoe+9OnQw4/o7aZS514dpb7PIcWq4yQmL0wIneQ8MXRNGLN4Sbp+ZrLA7
jE+6rEGoCqsPMLkN8AHHpURLwzhq1QtBqOJwXVATNlRGOrzgCFlyzRhxT0n+dtrG
jao/fzY29pgKHtwTX7lrPaAi/X8P2LI22mOAAta/CxRzODi/8M3J+yt526nAbH5+
Q3Tcwf2vuGd26mLLg1Y6aiIFeSvN8ZRXQ7o4r8MeumDviOyMJ0AyrKIkrOW5LtAO
iif5UhaupjDDD9lcyk2lw3B3q2kv8pmoW1mpjLiNHSJsYioYylQDm4esRrY2ap65
BX9t1nXVv6zIz+470F0TYP8UnZ3EIk/6ss84XsGChPhoplFmOKJfaqSzyzqry4fy
CGlpso37MJQ4Y9mEGa4GkQj46RNU99wGyPCT/G+LX1VrbMEXlhXejZytbDWOG5Mg
oJABUaHnrS8RyDkowNW5+9SYFUjIkZthOk8MhRRpzzyLyovCQlDy6Wh/3gn6FcB5
zgpA1Sj9ySYtPkHN7pcf8NKBV09FFTTKxfOA7MuYHMVVFeHbPVLsR8iHcQDU5OW2
06A/6feZ7FtfKlgq81o5BSduJLvV6s1/rv9qU56/CeXjwIivltvmctrqiLM1nZbP
Uhn/D81D7Xzh5ViKEJYbPPZX8XlPil52vTxMNqjkabRMPrhWIEjBEx+tZ1z7lj1S
MjDRDrlZpNVI9MyXYfbinsNvH2l9pFCJp9n/1jQEWmvPWLyVSqVSkBdUb6DEQ+lY
hLHHt7IuAI23zGeB27kjjvW1pLgXIMe5m+jST/pitsx2YzNw7R/kSpixs7zG1gJv
RtzcEjYCi6COur6OMbEVzCSpCd62GUjtnEwTvNBhtQZ8xeIKwOfqwWPaObSiskV5
K/8qzU8zrvLANwgvnzLkNqDa4r1HbI5QE6LOocg7o5tvgrKDC7OGUlGCRk15LTya
dGgluZoyawsQ/GgECbONaGbphd2QHKxmw6DNxikzIWw/pi5WWrpGQvoRZ6G41cew
UwWbyWKxpWBkY5EZ92dive6XTjg/cXB9ZDnCG/gDK3a4DGE4y+uRkf/8gPXnvgxW
THkPrHOCdiuOuHgWKPs/hAYgxBbL+nInGnz1/RZPUAzd2qEXBwsWiDz+MGqY/Bih
W5Op1g9Wf98qPlqO6QLaaA+Ow7OZsYSj5eiC5zTJMb++ZuU6QBqQ6qkYPDscHF1X
ZrWlvK5w/jKuTfscEvD+AHwOMPyf6ZfrWL8JOfuXVjaZVpye1zg3tWM5O9hYOL2h
RZQij+32woCG8b47C2jF+uBjIjI0xWpYmxBK52bxH5XP11N+o7ql65QseEwtrrgU
ZYAygvz6TMDQ+vjHVsDML5GFHJyMRSW6RtuJZhvb1d4kgy6EFNTpwxrZa9zc2bm7
9knA0gg5wMCdO2BeqD5IQ/41CSx8igQDtddOxsFCxCD73WM46wY+v0yPXAc43J/B
TfnjNs5fu7dOlMfNkn30Yv2VkoDQT3x69wDUZdVQRitztTv/D5Famz9j8lCoRiDR
rm94GdKc3oBUCao5FDnIju3+clijmh94Dp8FErZ/MS9AqVCprUdaPm4e3wkiG5U/
Nb5g7eVILJW3m4lWc5IsWmql5srVGjq7vPmszz7DJPvtyVXy364VNNGObBcLrYnA
uOhIGHZafdIY9iUdW9boKFvcMqLbTmZrhnzRAA0YzEIdrbZxmOiCJkxFIbt4njQ3
uMSbCPt0pb4iDEtJkOgdjFoymZWTLL1L3hFLizWiw1lLr637+pYkCPFpiganyDjy
dwd+pNRZ7Wa9eUkZtF6XghwoA0BnTKYgw1stj3vMHKkyMI4db0vCzk7KAmC1m/lI
NcofA0ecRPmvbAvZzDUvUj8VyRg2g1kn+AXhZ7L1m1mT7tzZoeOUn7twzBJiOEnQ
Sjng4jNNG1fuzGPHmdzmlkrjps0lfGvSFhPSb0Q2bKccxe8zWZp5sCjHduAj6eMp
CGq0WzVOJbWdWpCa4x0680Ss/nZ3x3iOMdx5pCaqCg0frFw9+8vMdckT890vFqjh
GQ6lxS0ntto5wRDMF0oPpuy3Zp9930AYaOFCUZQn+rOzvUlPEkF2xgUi3fZKVtz7
AheM71hgrIcQd7uJhnPBwsarAE9T9xfVKGg7+/M3rS+Kkzm6q6KwONxo8F4jXUpt
XtRu7EuGK0+Evfxr/YPx5uf5m9kBuiaApanRPXJ9dPKeUhDxmwu8bmImtunHJ2uw
CTb2ume4ZhSPLDs9S9qUKgPZdVUvdbIfnNUeuWgpxlv/4yppeZ2WkdvnoVshcttb
op8m8uHcXr+xA2c9RTL1wzFeEoN0yhOEJhb5Jkf/HCwIhVD+d4mWLQh8PYjbc+gv
gLudYel3bKpVqVtexVDySa21srpfHrnhG81f/A0JrZhfWnKDoG7IL6BpAH60ABwW
YGSQHFPgkB7hQm88oRKu8J94GiwZhh+ph3Fb4wsZM9wTAmrpRyL401UuZQ5/jzof
uloLgTPeQh7F4al088UNjLI2chopYgFLMAE+jxJoY/Y8pIG8r8Bi6Yhz3hBo7Xno
Y3mRp0gwYzPMCkHVpWjucI5cfV3LcIW/3dP/PlpLnDJFflnQaGwTw3jOsdNXIoJS
YraFC0yI2vrMn0SKa2+UQaACKpluVP9Elpc/a/wE02V+xltlwmcVy/u4YCfsv91z
895T6PWDI40ynuTR8X1Rwx39ZE7cs23HUj8jdIyxqMlw9lP0NaANDLseGyXsnLRT
PPKKrgf1wH53j3itaKTBO7qGOazU8z6QbqkBPMpO11FgeW61SXP0w/LerRehgffm
jureVH40f6EF5uFT/BG5UMK/GnFc9/FeNEer6byEfR/XK/iYCd6U/5Wi1fjRlUc7
nv41obw3w12xf2XXAval/vuDp8gaq8azyv8A2I5nsoKJOr1nnyyg8dEKxClbxpws
odXMGxst3tZ/mCWJzmTkaxlR3S9w1gUlA34sN0e1OvFQKioILykGVaZD3FM8WIa+
QI3cie/KWLtcMa7QGuyl4MNtHyUMFYHzD6pWGXP4Uw0kATL8vv3LURSXjLPcztFS
rn7rBU5gq1rro0mYtxWXX4h8dXnFVUrqpBissg/J39y9QXBRjN8RwTl9BPVPh5NM
S2fsUWjfAQkKViBqQapnLRucYxBDvNZ7cBCyRWUoh6hiYYeQ/JOeAzzOD+g4yEm8
HXY7UjWhKOzNOfYM4Qw6X6Vp0t9sHSGvwwJ309aMUWzSzjJH6w5ofP4JpSNzKg1l
J0IdkDUgarvD4GD0ybzIJ5vuThQcUaWSi/d3zKtlpOfZZblTeufEkPoWEjJGLYbO
LcE/rm8e7bIL8waBsYTeeXXmRecMrYJIt8Rf8aVHbLroS1JLzDscKAmE0vnLb5Np
DzXsBWLr42rt9o/yU6SFSSjClPkpDdaVWUhz0gpBbwm4z5wy4dM+6l4iKmdkSJSb
Uf4vJ04LDCYMqiVSh1JFH2YUBK51MCMXVqVdtplLf98932EREdYa1cAoltzU4A8M
I35bRQuMlEvhb5jkNj3XFQSSivbqDEiTgWkSSiPJBV7u88YSTf1+RWHWXrPRIbH7
azHNWErsck6vBfdFqUiJBGllbCePLDi75BN09/GhSeH5UifmVazVbc8CCIDsRHpu
1q8CrxtA280/FX6tO4NIdrQrhplf7lrjrmKeygbz8rs0WimkkkKWpCb+zd0IlvMe
8cxz54N7N2lCTij+zmPkFNDdbO5vgfzxouvszJifQ4Vsh0y5Hc9sxykH2fA+SXNZ
nghNH6/yJcfEswDd59CG3c7CDfV48lH9fEHbfdikgjsKMxMzwMvnb32Eioe+HFLj
0i8AcOu49BIugoyAIKqRr9nbdCTjXYvvrERDPUo892q0vJpjPyCNO5BPOQxF+W52
vfKk2TYZXBFFTM91h62qNEFsoUiT362mKWYBAxnu9JJhR9X9kF0AHk02fsmIYkOV
yxbqBQLLZ/fS8CICZxSDfAoXcT06a2r1twmZsqts1qDICII9BQ6sGorfUxEDux7T
KRI6IyJKA5v49XfVGXoL92V51VhEEayFYLTKDN4YLoDD6usqiCLZPI3I2jtdmxFa
kRB84apyjSh++h8CSw5hpau2h9ly54fgCgJACg0Vvh1MVYrhUqqUtxCxvtRubMDX
X376xB21So0glmwoKfSIodxnd4nuylD4FFYEvXNHQw5ESKv1lPzgBI2L+Bv+Mcxi
ETksaeZAG+EoUuyrLt1f3pStFvuB+QUGiANY+bMnjP4lt6w1D1tQ5425eeAhB7IJ
HU3u2quwGwA9HErohrmibn1qpSmAxc1Tj8lZl0j4dH31aWTEYN7ALN0QUakZomTt
nGchOf2loWHOGGzx8EpK1XLAm9Tlw2EcBfuW4Y1Bm5XI2GCRZGzJl71UgjzkoHwl
DhMOHSQEzXQGq2ACJjxZPxFYcgv4YZigdoXKl7QUET1GQGZBmCY5pwlBkwohtzoo
SHoM/rr8o/wWJKag/Vivto6CWLLgTKrYE6MDJ/Lf6cIrHEnvyE6BySK+Xl2p3ArY
1ZMosdDJTt3nM4zWl3fdn+lwcDXuhqG3oQVDAKBIzcGC8NnnTqynXzj6rZOmknBu
s4N5ibT9cAEvFLBaRpH17RjA6YPJTYp0M10fAKaKS8hghVq6akRd7KlywBMN6opZ
cGD0HS+v6g3AEnefeMAAf+Ov1OMI4LMVgwswMfZNaZnkLjDUx6nOxqS1O6yG/jYF
/L6dRFNJdRYFhh1VmkzcfCYV66nScvVQLbPQ6FconHM/T59T9+Ah3y3su/qWhSEz
6LEidIUJh6L/9/hInxrd/U9Aw9cJdF7np0VVJIrJetqLfktGyT2ASYTtqTsIdb8h
hZZKRr89b4yoFZ64MJvwuAcj4agwv0yrzWPQPsXIWS+4v2woXZD4JQr+0IuY1k8c
AEMBt0Tk7NnbRRVviUo8lGjgn/iFCPz5RK53H8aCIbC9OvVwqxg03Z+Lhk3gtCyY
sjY986Ukk2uiDf7x5LndBh5ZgezeqNLQSuIifmPpLtwpsXVRRKB7XuE9gLp+peJ2
jpyfrSEuIwzBzgVYhwbok2pB+rPuFJaPjEYyRHXgzg4HOwN1IY/sHuLrq9AtU/8y
iYI2AYWazrlpoGaqg4JaNdYShtxL/CAAFAcZrBEzw2J/81exjGf9pK4cq3DqUzIt
vQBB/SB1AWeYUGDBVC4sIIXu0kureac3bKa1dk4y3OBM//UEM5l5ZKdCIhmH6Gp/
qsL5Gce1WF8sHTYgOEueV2jYtagQTBlQnbUa/A6btetACiY1qvaH7c7anu9pcXjZ
o1rUzx7TES6++xTg0XYezd+5tDPk5+iultuage28oUqWmhJJZTaAyhtmw2/1tcai
VChTdOpq6iZHvf0ykKUuKYJBI8xEkFFMMZJpW36sNBHbAoBImDr4m9cIx05T0HQp
H9/JtnTJV0x2b+UapfGzOFIlpNFV9x+Kt2aSjkawWIjvyMgcF7oPodBni4FsmqQS
L2WLr3hhaLa7u7UK0sB89lHE8R5f/JkHS6nG9GRMVQgB2rX5zKiR3n7yAuNDlo5R
XujS95tLsaAhsPifaUXM82g5Xni2o4EaQ+a+K+OkkZqyOPPyPMKUCfAzc/x2Aze8
X0AFKoPYUe4c+TE6D5jHYh6nGzqHExM0Yky4Ojdk6xgosKpv9o9FMi+ZNCFNhr/h
0s+R4mB1sFaFCeoASSxhINq1XFbZmUG99Xc1RYjWfPA3gIUlOw550PKO3njrKVpZ
YQqLX4oTDmNR/rLClK0zm5Fps/FQBvaMEyWy2SQaTS6ttppolKpU1/DDGayfKWga
PMbfYfTgjPrk8o9DAPhd0OMzbPWSJJ5x+0o7uOhrT9HaOUunpzpYsaNDnDkf0u4k
1iFHMvFflXFUqcuBUyOpuaOaR0enYb9Y8fqRs53xw4x1VYLcqyQ6YLP5GYEjP93R
KggUZkKIRL8OsyFzc9GXVZ2wT5fDD5VxwaF03SqA5gbUtqMmEUM4DDXjm0wYE8AW
GxvoL8xg6BrWygqHjQYQLWQsfk58iyMJ1ll1SCrNmbqG1CaxYeMMgM3VTI9M10ny
2MrqcQPEcbDmVMkPbUvQcTwJDouCMsGj7GAzn3kWQxyXJC14CujvAVPyOffGTMLx
JnT9FiVm4Z9S070gz3BqeBlb2WUybNjmk9F3TH9lAXPkMngE77wQTveaWUoiPZsn
1RyJeQy2crm6spJVRHvu6KNd5VyfXXa2cgC1k35mceqHzR2ewmzBxkDHpWAf0Aix
ba4w2yY3CyzV0h8UdlAHpR60a+JfSo4EJjOs6HwIEAGYZamAhqHzB2SWi/dxAgXR
aprf4ZEXmp+vUyUmXqxmdQ+A+bQjBU/IWSUdPvdxOvSq4gWQb+vFhrxSyAnHSrZa
W32ZLpzAutCBKMx6ykLa4t2VSHuP0Ts8v8T+jB+btont80McIaS4kMhuH9VUCjXW
SqNsbUdd0W6uSJGf9znl4++eY6N502cHT37/CIm2dM8BORTK45YnmaIf1spOSE2O
XegI99bXplJvqGmjlzB5IiLpMcbhSvfvUlebnrBeDXXYuBaUQ9XihN1/V4DiZLcc
gJFldjZy1FNXmv4tSzeibGgyFZ/tlOW+zFD47cL/a/xrAjAEt/HmmLFAXHq7pqfG
tOQWtzr/ZguPN5HcflfV3hx880zIDtB/FKl0etygzyY8QjfL+qkdQ/zsEDugr1uD
UqJjP+EndCzvmWYGnf9rJa1cB4LsoJHM+tKoJ0Kynn1GFiiRfMpkgE15otfkAYU+
OYGY7vXUTpgmx2CsREArjXQFyCxQ37J/4C3gx4ot5QujJDkq5COzgU220+eiT01g
tTufq+sJiN/FVakIao3n+0oNNSMBuLnaLhuULJVw+HucHPlj0CoqZJnPgmRS9PRA
fS+Ge+K5z2Ew2C0M8bwqPhJkO9Ht5MxJR9DiUBIywDEdeiPEUEuNt37r2mr4lrkv
nQa8LwcRAj7RDLW/H3yKoZJwQxOGGTQ/YoSCmo8AA3wTJ6y3/H65GprjoN9SxqZH
4npGr/pV03HlRT3mcEFSRh7KIovZQO8b98ldgtBUhH8nrPynL2CnIZsyW2hPrdHf
O7uzekV3KTFNJyH2y7QeY8/6ZjMM5iU9ZQDv2mu5Sk9KrIok9qpacgCdE+3/9aAC
UiQRoPJtHfGUiZCPaVjaKpFYJA4JO3I6fBZ2ELiaHDjeD9pnL+iLp8+i9fPCg7Wk
vBYKfhNyo32EMBokAYTRfVTit1B3x9QYvAMUmrdiZ8QH8Ti08UVJXWbfxPnzrYCs
8YPLgwNzWPAloIznx67I3LN8MEsRbKdxmpkDWlPvUS3MY1Sk0HrEsHk81gb7zr32
yy9zYKZXP9G/6iIeshFKDDCp0zBQxAiK6wEd0CEFpb1v7m6cRlP83SmjC1iOPWId
pc25sXYMRK2X6RdUbinsKcNzrNiSfaZTsxWBAIwkIFWhdTc19zOQBkdvrGrwkTFw
fkeJThQSCyTbmtz2MJv+J436r3MG2UVgHfhTSmgZi6wkTQrwHkcI6MhK8MmZ99RL
rffc1wxR4RnXdhKY07jqToLFOoyWzfSCoyI5e6V98OjF/ecC4NhK4h62O85TNw0W
vAEB68+sXtS7EGjJLnDoXTIEmHz+I1V3NXv6KUIvXfLFVb1IwMFLTc+sI2gG87Tz
Tdd1Fgi1NWKmZ80IAvOi3OhXrolPareKDOR1VDPeJ5gba1T9dItegm/q2d2gcHQ8
RKoRgQJiasO7bXsEW5gPzLCZoH8GwDB6GJsNfHSnIIDsJmKyXgOYmLKtVqmuP0va
N1WN3InZHnw/cmcgQztlunA3+3tU494NvikH4Fxwh/YAuPDf9yxbHomzA8a+hQnv
ae5PdWxY1FJclRJzCNfJnWL07zXzzyjIjSUuTLd2OV1Z+5rXld9MtYAacPzKar+L
Rgqogu1tfMpVHylMgh/sAdymnodcQFQB7Lazmh1q2RlsVTZM4If6m0clRwxTM0pu
Up+GUbebeEahW3ddLdUboLQv9HmYcRKcatId8ujBiyUXZ488LDrpY7R/ClOlzvHq
RHGlyQsFvGdRHlqq5B+PEJ+BUBBKBzNJZseB7RXw1UtUf0NZK00bZGkb5Zmeseka
kPvaouxG3GN7Bf/BvRLDKUpggpxJ9ncB9p59iaIEWyZFX4QHFj6W67a9YBFKynxy
9WLOjQXKwsrxpZ8ukWGZgu6tE8rHEFa9oQ0plTCAB0YO5n/OghtH3YNy9XyjOb/v
Lh2Yp4i6LFyWoK9TBK+obgkhAUbB2yUDvF3oPxMUE/QWIpsvvTXkMSKgxfJiIgd9
QoSxp3CzQgc7KqIbShPYWHMKYevNatLImqFaUxLwLABpiYf3OOhZkLe62jPZSon0
vk8/I+wdOEfEIs8PpwEfVD7/msanwwxpWnovWQXtCzulGsqVkE/5gFVZEHc2w4D7
OjRjhO0HgbOrTI2yg5j5eU5Xk3Ow39lVJ2EOzfNkzfyEP1BNDy73NGTlaYHtAQGg
QLG6UM+P9JDkvUL0H+pyG7SQ/O8gMT+36PTU1DcIf2fOkgpvRYTdc6wuLNSC+MQM
CF9u9j6ticgUlCEiNUv27jsLOixaFyb8DLER+a39k21SR43Q8R6A4lfhmdQ7taDV
U1Ry9Un2EZK2vzRl8BRvK5rtDzXDkrD/LHh0O76OFa4suSfxVPBKnC9FMvMkq/1y
2wG6OuSvHFraczrwdJcUGyeEOIUU+ZTVVc6NkO9WFbp8hmuWAb36bQkRgXiHJ6po
dwIQBt+SOpfamFtAZbwQ2KC8cvG6rziLRkh+JClSD7cl7t3a6fgFODYEusZ/tg1v
qS27XW7XhTsIQmKr5j0BLpJLQJlQkS2fweEnviNkVVmp0SanHnHi+GFOZbhH5KjQ
VJ3KZKvW3wuPr2NznZfINgNVPbqjCAkTHvZi+4pcGmOSq5HPFzJusrkQulv/KZr9
p1uMpAAgAoaG69z1W4Epsbiz1afevF1T7iPb8cUjbmuwmXlOHGh3l27Ba+a09kRn
sn1e26ch0E00Z1q2CjWqehKZTLAfov/x0TPzZTy5W7Qp41VLwzV4fUhMletsVlRu
Z8Bwd4lfxpJj2YNd7CiPwmy0Q50FhkhTXppjKOljG/E5ykOotlCZM8h4cvDLZHim
EdNX8aiD0PrWgv6fpw1v0zRDeSh1/STbFaug1uAXpx23ekqatyW3ZhHcKItU/eQh
FeEeKdr2EWAKw6pLk8LZazqF9/u0h9E91jkuJ9pG9RotK3bhCQw2XnCpfvwA4Q4m
l9TsP3VOCcBs8s2+Qw+5k8Sv5wVq2mOfaGSDSEmgU+rWhk1jFv8UGnVFtQNkfUN+
ckQhFupc8KjdXQ03B9KUMIcvdDHdcxTD1naIdED2xUvrAV0al1lwe9osozxtrr/V
dNOLtkV7ATOY18GxwCM815za6FrUuTxl0N0m8TjfKCY30eGVwQd40ZFmAZKRQxl8
Igp6Pr2998/OxqmRCrtGWStRk0UM9BCgBPwSANati+GtL/KyfnLOa7Tabg4hA9Xf
uKYUZrI+Q7g+or5HYetz4BntDYBzSGL3axpFGrc1gVZ7AA8Yh2LFbSMUfZFm6+qX
P53wJPS3f7qfxS29Jr5u8Lpi3Nt7g45ptBxHhuNerFWXFrT9OQfJxnHTHC8FaTnO
OEIZRDQO59jkr9mEClRnr/vJaTwPS30IU6qolD+OCB5zLoLTDAGdCT2RWvUtaDUn
orQ24ZZdhF/HQL+eYQ+KAJVteP7WYboKzSLbZbPcXDYgAc2tSZ4Cutfx+baEBmc5
+K7MqLp91DZRdCIaHbb+nERXsSih8LINX/pEJzor+qky6Zf0kQEoMMAzj3vPuJMX
3te6tDJ7l8Wr5ooCh1Ys7nmL+E04guT+UMcJfQ6+Rd7haK0nsRTHr+WOwIsNxZn9
E83KjvqFdIxRgX05Rwuw+xWn+X843jCO4Mv2ZfQ0xZ7Vxd28H0s1z6V2fE/JDrIz
Ruw2hOjWoa61SyZYQWfbfrTdjnALJodpW0bdwEuNl5vOiszWXmJahipSfetU/dfR
5KxWc9i7dZvxU8guyMbwV46BeZkYHyGmT9cKh8W7/a7sdKqOQ3Ew0dtQX8HNnJh8
yatin6fXHf0AJZkpq/jHzry15cjv6Hhl1/NIj+eK0a5QQomsn9Oh6vJnQbFivpyp
/MO4z/xfnApR50JbAi0DZXMXsikH1ivMATtsQlwXLo1rOWxbvivxFRVHYbt1+AHt
pQvjEnvbF3XKK/GHBxi35fV1wJHnJPoXj16IkuIsAGmAkNLVYQyThiG+3i6xEiCP
GglZpD+FGtXjVrc7E8o2ZL8a/fI8Oi32tBTQzvHCozTrPteML+xCSCP4hzY0ez9W
tf3T1diqdX+SBSBXYpgReOLBVoyAwgdGypmHxbA2c4tHlBjXpWmZ73QYE1JtPpfg
HAeKdpY681KmE2vX42Jsv9yQzC1RsetTPyz2ihey0gpiI4AvOTfxVulhNHXmiHRd
SkOzlDoXClm4PL6iZnRUHszxgX9DCNe6gDfNw61/yMbSuMaSrCmCQtOLijm/Ueg9
Y6giJg3Miyi8had2fAuJnfjaBcnhoBvujiWv4pz7c43Z46pDWi7gxjIGOJsEKCh9
IJYYc17uMdTUPCO9rhFherL/JS5C1l8Qff4N+BjWP73Do0cn6lqHLhzxYhvLnejO
nmKxi6CAKsDJaLa9TOM2p4Mt+9pJtfhmPDFp4Xmd6Xvsa8f1vAKOFGfKYhw+kKXB
ExnkUrMcogIxqqJwlt2A5I76fypkkNne9WTYEIpAups/Pj5Yx1dufwbGtuON0Hjt
ZR5jCGeR3hFwaNFb7i3X6q80iGiYbPpfypDRSwJsLJd5N/yT3lGk3L1P4eswIfuC
PAlYt9tSfc99YxTYA0zmvk4HCQnX54ALSqTXNvYCM7Ea26ZYVh41F6as09k6ERoF
TPhgjKEBITDqAjtb2VU0LZPkWNIEdN10lMfoTdURq+h3bkne6sRUuBlSMIOln/nm
IesMBX6MvYOdzYskFVspivooiGTJ1wReN7fm7vUWB6uTVkSyUQ13UiYQRMsplFqy
dB5rQ4JdIqF4k5Mc8AgFnwyMMI0Gf3p4yTseY+GOS9gGcEsYd46UVBJG+pSewCwl
g1/e8RMxHCj02kfuF+k57b8Rm5pe/KNhrDy9cP84/66r69Kke3m1XGJAz39HfFgX
hv/TYOwejYmgt5mswuY4rhxQB9gDgbLh+Jj+nue/uB14dgCIsKE3261tqUe8VzgC
RvUJoBU6j5a4nljskBqKLOYvT3W7usO21EcXZITgxCMnAKZ50WdtAB9ushmzbjSM
yssLS2I6SlnEo40JtW1Q8HjrUnuD7pcKQxffQ+T98uzByRrgqjrysmhAy4bEi1fV
ctki00T99nsTsgTPpvp+guAtakAghpyKbalifl9YfDePMg9ai6LHbbYIljBVneHP
GDD6JR5Xn00gn+uZiR1c1rsZrx0bpGefiS8NjnYs9Qua9tjaGvAW5N306nRv08oP
+nCpWgKjXdSaX0PoZQRbHJiVWowFDBkC4IfUXz4Zq3B+nOnpktV4Xms59fe+NZ7D
yAu7rnMF8FVugwPPCDjnzug+e11wVmItfT80S7PULel0HQxqaN1dtVUBQwymEPuZ
6bvVrly0ERa4B7uxAWWR0Zo2cGyBfeAMmNPg4ca58F9MYLSdLhUKKTQRszSAui7c
yBAWpm96v6+3pvcs0epay84b5SC5iO++rmHVhSsRZJsVRD+oavLGESmqG2BY3dYM
39nw/MQj9f5avbse3HE78y4XT8MwAr58Ei3mbDe8YwbIVBPRLyleTi0hJndozEYe
IbN4csQ+YM6SgKb+BEy4A2U4BF5oznInsA3Ou9UcZVHQbHeVvlLRA1FixRWWs3nO
tJ7xxPehI2fA2q1b1vANzC2KzEiUZnRs1EtE/aycmARFwFaHbhgwOsjK+3T+M3xw
/35DLclKOkO3VpkUIhCp/4pyuRF+8yRwTW1xqgkWBbsTS/bSdwnZjGJn6AyqY/c3
TW1wPg4gbEMld9F7l4zLYD1D2fGJWR3WiMSmhymQRuZjkPaYMV9e9bC8JDl6bAHB
JY27jlWGV+RKP+n9UD1nFbsNCDgCWbqYoFqOP9KgtItaHZjs77YYWvbiFW1dosJ1
RiPSnw3ylKmdv2MrRE3qJV/YqXO/Bvl8yafflGtM41ONtb0SW4e64DD+ZudRtIOp
WR8c7xFKfvGPJNd/adfMjFUunCHOc96CzbJlRD4oAti6vXknQW1ChNLPdMOFJ1UO
rG0Tf1ckl70q/zbTMJBRZE2YsPOxl6pBiWZlf4B/YVj7cbTHakNPBp/Tji0Zd4qj
3T5RrhhglETfhSxuIxPGUDlNf+796yqpjpZdhly3+U+f/AlhHnHgmMJC8drn2FmO
MCvuZQH32Aw37zIrlB+nvUj1ThrKi3mTcI8VH/UD5uAjfc8y4oNqqYmT8HMGdbda
T695MD+5U9WzqB75LIf9qpQoKsmLAwGkKcbPzBXyAcYsVgJLIOnk5wwNA30Tjqu9
62eEk5iiRg2l6UOV39lK1zPOyg+SDn0gNvVvXwpg4qICBMxkm27j0eE8Rsx2dy3O
1Wc1t0pfjDXK2SNTn+p8weDJrUvu0XPFxBqkW/l6ZRBuyyltmnu38CZvXHnuYYSa
kHNjwiaRCoQnhaLCNURFVjARGPzGrnLoU6RWIwPVolNh8NRXuYmm1eaPnY4oeD+P
ribdViMZmPCIwRE11/JxknlTk/YNogPE5PA7amLj14OLZunv/GdbXEItASv7ecPJ
dvcyhvre+ztfa/GaQI95VdUrnj45ih2pwDJ+e6mN9qrfPGAAXxeSPXcCzk/NnJR1
o5KXOsstSYda4yQXJaqImDswCnAtxVc6YOmgqJrKy698iTx3vFP1MtZrkJKoJett
D0lZN0yuNR4+iu05hybvOisR8sOUf6E+RXnDsaSOZYUy0MSnbBkGXLDlAcyCfr8y
/OHOGQrgWj3T6+8/SbCg9DsqOQSDmuUNfCwADV/4Rx4jHEWP7LVKOZqvKCvqbbRs
9twbuhGh9vjGx+z8Tv2Lxqu9kuw2DadvRS0cNqbgd3QbukmML5heEBIxH1PVIUAY
Mz1S3/M+XMbmt0XtrcIwmVC9p9zd/tk7SwA6QLXz4XmYctAXCfn4i+MPgfCta+P5
jFoR72w4ZOyY7xlBDL6cIN7wLAmlySJ8rqdHlcvXpjj97Y8YygbcSbXqu1aKG+//
fl9Jkdm7PtJCc+nbhAC3Gc3rHvnWLJOzQKMATwZ//sycIy6cUbcVisPq2zTpNOvV
3dPOPPvsEM04E4cAxW1NYYc64oeU6nCHOmQzcLQdl+DSA42t3NRuEpW1BZOwRdu4
S8JlRYU5+QWKbdDLb0lbXNYWX/1paXxQFi5YMatfJ4WMQCt/6MSIZYoHM8in+V0f
82Y/WOcqFAEkPd511tiOTKMmnAn5S/rmrFCB2pkX/Ezwy18AuprVCTg8UhZrQjuK
5Rdy31aLQAJwpV9/ZqJ5QwOontYoWObC4X42SgiLJpxmDXb5GO2B0/y6R0Uxsh/o
wXMsU0qYm03fBvIP7sOyorT1wG3G81ITU+Y9eE/jbhoxPTGwU9W5ZrOlnBHPnXjb
WZwJld3M8Ea5WxPNM+xAyHnBhUBkpUR44S3n4k9EewKgXC1d+inhoS4z7e4x79w4
vEuoz504Ib0KE8/ggQAASeggJmPDkV7ZJKHHDq3KVaIGngNa2vKXaRVUjHM9IPfX
QBOmQPvDy9NmXrbGarrpDoEEazdcWAN7YdWbrlINrkRhLF10lUQZAI26kPmcCgBc
nVSatVCIGKE4N4FfvaaCn1MS8u5kQn0xAau1gHPaqBLuu1UQSJ6f1E20r0uth2n8
1B3a8wl1hQ/C0DIrWgpirIWwjmQSYgIfIcUA06YkXtX2Go0oPbv11s8tCyRYezOX
ydWx/OSXHWuaSD/SSnrWulyeWuObJlGGSgr0l66UFQYWYBC1Wk6QDoS4g8n3ekn+
a3JxhLz3a3lzJSWcJ6SmlnkJteZbtqfraXWj67oEM52QwCT9Bd6fD+SsSOul9wIG
HQE6utg37dVHjH3QjiEX5iXGsOHFiUt1WAPkg9bPGRFBGb0FIvpTzfVQzBUbI2N0
Ucoq2kEjghL1NRLtMuiGq2Qdg87XW5Zv3EGWGBumvdiWmrMFIHFd47SQ1Xi/Qi+I
VDbSWpt5LXKhVbwXoJD+jqVUmCAoBJtzoSsGu/2QsDyGG7Lm3WR2UzM7REx9NIdF
AbMHHiZL0lR0Xi+N5KaMG+xYzGNaSmWF7L5A8/v62PSulC5EiuIFGRDALjekXxd/
vNQjdch564xUzR6ldcE7SyeuJcswyIQhYtwD8dHKuWLwop0vSFfAIu8b2X7NSXgi
tw74LoS7ezvoFRLonmt7npIksoHncj8nhVTbIr2N6Gwx8CuqaBpPnUCvXv9yKVhn
bn/4qzLFjWidBQCqIpIbLmdttpus71vY9znbJUbPsUHByDsOIltN1/tbKnfgjjFq
CZwww/0pZRZdPZVNUPhKfalTgOcqq/V/c7MtMCm8da6habOcT4wl8Hpkqsh/T1ot
/bEfAxn+MogL/IyFNFWOLvHgsPwv37/QFryjMGOz+S2NzDDWpsYYXmXcC4JswNpg
4KB/JW52MPINrz46Ks3ms0UD9ljvjiUV0nPrp2PVk6bu/3VFTN39rC+wEFl+baht
MunEdLJe5V7R8gt48yAi8PuT+Ud84UDfvmtcJybYZ5dho88tSwx6RwQOlkecEc4W
sISGG2D7P7E0u1AF8bs4FXdpXlFUhBhJ3g34AsSJ6tyIOe8nqsZWjjxS94gzYXJ1
aCI9xuXnU/UX+vximQ2R6Leu56WN2AlC+s4c6OKPLZN7MT3ELTP+Eu4QMlEtYL0a
ybGPrP45S0X6XGXA4cf+OnAxWAJ6faX65Ad8jpvrQxTaFY2zDg4AOOHeCEcs0/6o
XljAu6wCRT32ZwedrPEoyetkPjAdMLt3dT6W0LPoPYytI7DBueP3LAQziE/xwMBv
j8cTYyZ2Rvu2AjM5zf4s0bHlu59XCUF5PMugFMbGUNmdv0WScrxZSj5HZmTewSwi
IJcZmn2PLez7b7za6I56qH9c988pxJkDt5spTOlhE3iplqQy+AkG7MF0/EmpOkti
UUB8JvWeAjkfhfbXiBbqE2cFDLZI3ofHP2epB7juD5zyy15Zock+dGmSVSh/VS2w
WPP/BSKaAVpY7+gyTCOambKi0gY3UM0/uhgQ9tDZ9zA6ED1oLmqa63HNP3NnKbvA
wEa+uDT6HyG89b5le6wPTFPuxHuVkgcu+3seZYj3b1AmMUUAx4yWqM0Y2Uy+lGKY
bG3o6iQug7warw/UuUXCv1+NMGDmPt5LFdoO51LFA76ITJCjGZxZYOhrSeWC66nE
fnZUkJslcIk9O65EC9A69sUUNuvrO8Pcxj1lb7XkE4Mc5I3iftHbc35BFrSH34x9
u9ZZ+gGHL36gJk6OcRPMe9lQ6TP3dNXcOVD9/MR6C5HLvuD/yC61U458ooo4M5Ui
2zegt549VnXDPgI1xqOJPWgDhKMNVbIUVBmkLR4QDhxp0sZEttAn0aODye6dlFdv
hPk+r7DwgwxyKdA++9hChpqGTyC5wWA01bIqxwcuKAp9A82HzQpLKGfcERZ3x7NU
9YjtzXGa9F6ptoP9+wAuw+7OKtz/ruuN8jcSPMJBrNbepBXzq9Zn8e/HiaVThzBT
Vq2MAHSdS9+JNU3dtja1KjQjmCMxHgaBhWFef8CZW4frI16k0xff25N59vgGa+Y6
zUUc86SC7y398d39ScNgIhEI9Ilp2pT0dBN7bVovRlpkiYsg8QuHN+FNIBkQbDP8
aWRb/Se5ZWdgynijI9E2o/X3si2z074bWsmIkF3VX7oFeXfVfDW3N6b4Npy5QgUc
S78/SQBU74STjmQYbhdQxkQF3U503/zyduADn37Wr7Ex3y3rVZLFZrCBwQeHkn5Z
z4nsdTqqiRBCD+ndpRebguvQAjJHLODreD7aIf2EgZF1anZlnhXMx3YFVM26oBeL
njY8UkLhY3lcdf55zfn6vK09SekOjf5x7Q3LXrc4BjKI0mZIjTnzB65UUAQMQu9w
XpBpSuE8B5gL5tKIUDT1HMeprU+pMGLSIdTwcBfpOqW8j4/0GB7YDO5u7Nah1XhE
c7AK8Pn7mL4gdOw4gjDK3vBeUKubK46dCy1bjP4lwiFefvx3UeEQTjtdORCE/aFA
sfKGamLui7mcp6Jlui71ItYGh1H7dRAz3MAPra0muSNlXhRsN2Up64enrZolVT8x
OEb0IBBnfVelxi/CfhgbPDrkv1NWRF0fVeEGmyUgLRVia9AGcEflBhzeIF0efrOR
4E3dlsZmN6RWhCtu5GUWNUWxIdYWocPuuGaf9sy+u6yfooToGrss6FsWiKswgGOu
aP/E2JBKoTWBBWZjN2slGVjlM3a/PohVllOVCwNerbE/wVshLfbhClDPXShSkMrw
Tt9VAoZEyYK7m63wU/I7XqknXCcvHXJSST8JsLp5IDIZR6S9pnj2lAToHd6WOLKt
wHMGf6gR8jfZGb3KoODwzPuujRoaRCqStDcoNoC3HlxTq+8UwFVbIy4mQ4vnDeCN
yBlLFJ46nSc08KSBKlzrYmW//cRyiDgionHrBVLlI6pwJXo5tuX4jf2HBf3bNZ+W
YftDWzko/ZqMBd2FdLg7SLhJeHVWN/ALbJ7GAI8JJmjqqqJIlyjNYOAJ5K5uFsu0
jVfrvTmwLNmirdyG5cQIiFHxnN4dNEoUsHN14+DohX4EG1ZyN5GfdyXlLKBbaeHD
lfZhA28gIMDMXJw+ylamK1+qTq53kYJxev/m67F/47dFbdH1SGtwkeSKDu8LO8fF
zpo1pxTWN0v7s5lWviXrxT/grzk8bdlzGSrOMZUu1hy0xWrBwzlC/Yc1o1spRvVv
QKCSlYhwWoqo+IslGgF3M7/hi7VZNmnX2nI7kK4ubb2xqXbE1Jc98aQf7wPmxxnA
XUzu/XbpNZ+px6aIIUFjkyRHsrHYoJQOyF7tkVRAcCayI4OJ4iSDbg5qqOzI9lwY
nG+2TC75/0Ll+wZxCtNUKR2Pz1ZyfvSWBLbGd/u61UTdgZK6ywzAq3UBZlt25EeJ
ygJbANKwW3YM8XP/gBf7YVQdYQ0Oh5DcWx4/4aT7w2XLV4lK7+2mTKV9JK3l+wLE
In7IuH37pj/oXvYPJaRRZrSWbhrBe+WhR6UNc3n0taRM4ndiMBGFXOrIt87/BBV3
A24TfqlaU9ltFkQCj8Tvks/sqVQ1gVrX611Dj/5zpm6sWSEfbtSHcqJcABuPE8bh
O4lZA10z5LShGmj9eJRjxPrjqhN5UsQKdTPiVNf5nzTesN9vP04Vrzt9663MIH8x
4dwXOtAqiCJgG5pSlQs4Z8hEtjpAoKkXDZRkXji2troMEYmwUDxKlwll8ZOZtP8S
WxcGyR5wWSkCO6lRgmGE20lRwE8UAgbiw9tJenrcPEVpErAoHlXgXsD7Tw1IR96e
/Xsi3joMMalQO/SRw8jXbAAyPtYOzbHVCWTEOAAOOt2zKVgCl5tnzg7cD2W8rlj5
MoO9/J7YQA+MF5xkiVI7NxFhtyUOr3jqsZoNf9n5TzhqQrmC4eLcKZmXUPhz/HEA
U+jukScUXXIYCCpgpPwBLF49ytFlxZ6uO174UMlFHna7JZg7HOAR2rUqWCtI9c70
zM3MksfnfQje6wOXzS9QLCLE0Q9cDCuLvogb89ZSLsfOB6B9bz82pHYoKwmSRAMT
MVfSRPg/zDKYsgYdkE5UPCYt4Ba5s03VVsRhZqnO01+wd4EaPYJe5jKPkoe9nJXM
v+cp6BeqHYPfOx2HJ3NxC66/OWJInByDBSOQI2DCQBPFeQMRM/f0EsFZ0o95TZUA
KCuCiUawX1YKHzu9GQSFDX/6oG7QkLFj/8rXU/qhZnLgjIy+WHvioZdddfxMmRH+
VcPEcINanuLHcb/o0nSEYg+XMgZ9SCCIBCvt2P01i88NLcl6Tq+4gPa9oR4kpB0z
EUZh+mK/4KVj0/phLAjH0RPceOAA3rhUF2CHUzm3yLzuDO6b85/7aHzOk854Qy/t
uPt5MKp6wBe+wCsgN9UKeHXiWAgJdOBISQN1N30wUdf91og0G4ziQSJMwqgxtPYr
JBCz/23xD2uORWAKLu4epX+1Y79yaEsU8l9Ayb90UOay/x2iAXRUslKgcrvv7F7n
LFXmHnbhGG1fCcU4ci6rheb4OxUWw9duJx1n0ylFOcT8YnzBcNcXL7cd92KmFNaq
irWHlVqYEEcZz083yOKpArlfXiCOYh4Jwe/vLM7gTa4oqhgPzP+FP/xornGUnWVG
xry3LkXMTSn9uc0n7RRydYyPCtuO0TyXpQWEaJ9cJPfx5m4UQ3JdQ99FlOpwCZ+B
yNBkL+gLHAVO8C4KKWQo31s+luLJMukV2aM4c45WAtMCXS7rWADcw10dT+QzL+j7
Gx1H7Gs7h4HKGVduXZ+ORBfpMt2geuhHwymk0n0HxVYivJaAk7HE0m5WUUgrxyNn
Z+af71F5jc+/bNqgrXG29it5k2Uo/sMe9X1BkUa1AyZ8DetvhQytwjifm6SIodF5
9kHiN1cUYTKGzDHwr4HI5nRQdYkCfaxcXBBBDkwzxGUvCUZp3fZUgw0unn+nVI4P
c15oaiTwnj0p3hCRxMhwEC8TvC7UoukSlHdo85zxduVe3S+cOaWfnY6PWB8IY9+X
6XWbSrTOx2UPMAvc35bWWkMseVhx7OIbM4b6BWc0H2kRK+JIyL8qxS6MU5UBjVg3
dr9EGX2s9hASdYEWG9o1pO72mBE+paS+6XiOtIAZ+J4ynK+yc1dZqK13rkRdRbA6
zPhgIFmP5+c9H9NXRJuSahhf9/+2G4QBPss6ZdKmDDkYWwGHx5jbEKeQ0m5xPCMf
ggGwE8Sn6wyRGlAR5cwNauboFKJumdC8UWmhBKEyfiXkECeTe60LtUl/a4i8iiae
lHCxhp8YhgxgcBekVfVHy6/G2X2mwQyzTyjraDP928xM20uXqsNbfc6HHIAZYsXI
vUFLflMOOqqcZm+QPSfXupnHJC1zJb9z2Gg1QYf9AvGSRwf/MxZ3+JYuywvY2sFv
h1k8uL/TVY1YSLIaBhyPFBwLM72ylpgO4PThTRyt/okI5TIgoQMEgaXo3gHizdZI
aUI1+1GwGIc1XAwE3+Vdyidp3WgPtDsi7OhMVIiKTKFVgAwI0+++6HSgW0TemHIW
o9guKHOVbmLBmwiKSSvBfJxNGRLH2lH8K6ILSA7e413UgIn/PmEXEylXhg7y8Sr2
UDNEZgMpF2LHtI/f5svfB5RIqa83yC5YvmyGBcNOwV0/iebKwu2yeOty7Cs/Ojxv
0vlpB5swC/WBIZhjKQHXxuFxMGKz0KLzEiNQ5/uFMd6d9L7pSpJgGYArusPB0H5D
fmuBHLqHPCNOCzB4zo/pcqcC806VqR+d+r02wO8IGoJYPAs7fNL6RQt9/LS9wp2A
RMXnekZBXSfoYIdDKr3ykYpz+PkkoWkO97qlDyKDVUhP453xw6l6asP+cfXKYszD
AzxSzngrlrXCzupf6332yAPkabA3+Amkke2nHJXRh+CNIsSWwui1XkGZr1i77fo1
frtZqYqrxuRRiVKY84MVM+exzq0nCgrt4sTPvD5g0nIe1dWDsDqkiuqy+PKb4SEM
cqOvtCwOcNx+SbFEAMXqa3dJalRTBdCBIffoZT8b9VRUVQ00h1HSOBJnclDkXsRK
SN2bqbr9CUrM4doslFeoQ/dpRT4vX4iHCZN1DEDDpuT5PjnEq9RUl7i7xMhdWjFa
NTGIx8D2XxhK0//JoSmSwwH1vlvAy5zj/MEkLNnKCu9r4Ag4pGxUMAgoeiDw3zkH
hmMExum3hROlg6FElCwx3kY9x8BgzsprrASMsO234lOVAQv4LpFvGK5+KfSIFbLV
VwNY28vgEo57QlRt6fa8ekgVWseBxCjReTmZn2QMeKNmk2P+KwBcXusWULnZYgKf
yc4LTpnTXjxxbaH0/trh9ogoJSRdpYxkRc9SBrstHKQBuezKNnfHJ6pNB++wIem9
aDuDIN+HGkqY25tvscsYFWKQ9bl9yCPouyvjQPuvTU+CkrLIi3tl4YFn3VXw5JpN
1lp5GpoKFJL9+EyLYqQzRmPHNQ+dWYkKoGQAJoU5tMpkNStARduTB3qn10vvbjo0
eliioYBY58LKqSiPjwJ89XPze0qVPVUaHVT2prUJPZdEsOjfoEf9H6ig/WuiDIR7
CX2yAoT2/IznMUukc7ruuA+e1r+jxfK9VyzhSHfS5lQnTwB4IoAQG2ShlRuHWKFC
TUmcXAWl5YHepR/DMU/ypl91Bnde/1EyjyMx3kvJX/FYpLUhIw7/xwE6TGWD1+yB
dMDXP81d6ME9Edn9M2V/mXv+8iXA7Z+f0DXloAUX4M6ssf4uRRRkK+j22O17I4UL
lPRzLWzYj7kPvVT4B1Jz4vBLWTX217xSA/yd4IzSQ69dMC838yTH4VFRjubTLpP8
KR4RNMWY0RPzt6uYzwrnoEIcEGBVY70qObU5VYe26k00yMPJt8vbxNXyk813DeNA
EKmC+D3VP0ffOEyQ8YSPxZft8Dv8xmZYEBa7lFAjEi7WHI3bgDF+/EGP1WJGyXno
KqoswhaWzTVI3i/csGS+XUSXXmsUouB/x8pWYlvMMBV4Nb7aJU+tAjtmR4IHXc1u
GjrdT4w0xGhWlgD45JYfruXgLS8OO73dlKHUCniA7B5Mzm7+XVJGGwJYT3WgSc9a
16SqpJrjUDryx3+8c4V5Y1djhShbtYXk8jRMqpscxK9FYU0/Yckc51M8kZ0jwlDE
hDhuy5LhBePyueAeQ4RBb2eHvGECcF6Er8324z4dllVnBQPdUeeUAFeomH4ZR8Ad
47G4QgBxKlseN1NY0CKQGyxflWpVuJrPWpUtlzNJcDBTMl9pzjN4OM+J51fpg9x/
mTrCVT2XHnExpg6XTukt/BPPYfgzrBpuYy9DhMq7a7/zIsxC4mKh25SNJk3E4ZfB
z2LAWdwyU1C0j3GehLB9+h78eBj9t7Tc4W1fajOynQcCwrhoLfsKnabrIn3LMe91
CzASh5wbuEKO0V19+fJdI9fw6GHDHKZcR0MhS1SLXOUb0RBvMO79ktfLr0kGLTKF
gL/55Py9FKGsLorjUMNYaZDrj8JNVFI1rYNcoSJ0h85cEaa2Pbyo26S3mzYGMHG4
IMDRTHFUgrPlcLnecytIbqJMMy1fcJCJaCBp/w6Wpsgi8jcqOExrj8f5iBqSskKb
EnI22qxUM17+sc27v81l3B3SB8gRSnoXYgFop3Xz3sB30UZZNMMYGGHIkuFLyX1z
2M9qw718q6vjaO6UJwjrA9yyjm2j/w8jgwsVmXm8lI3f3bHJDHYVCg3VEcYoR3zt
RTUstkg50bvzXUCva244KNfFUEdvlzQvLCMLqlT0/C0SXb6O5/pj6MONyXfYY4kx
nHdwbj+0hQICLLCCWu79bffaUHJ+sEZkHUaL3Z5lW/bjWjwDHkl2Cp67FxeNWSWG
ZT/ZkFX8GDr4hrLh5SNmLIoOkrc0IhjzQoQuyilqISld0BFf9iyLiBlEMoEubA4U
4u9zCpHYX3/U6bphsLniU66qwCPqwfCpNLqXaXFqC3qawhyl5WEVsUI3y13h2j09
VXhncLyoq2gManWsubMpTgq4FQKXAroVCYApcBP1G+ZGCKPVrRsHyxO8jtQcKhhQ
oWtrColG/xscXRnhIVbmoDnyJ+y1bEZdEMaauw4NHKSU/IamGF3R/92PcdlIvSze
cTe6ej3bxf4a6AAvP1am4IqTiKyhSeCN6BXdEPOpwd7Njf9nQkJsBoNWmCtzR0gJ
nXgFQdO3Zmv1H8SdfMUUZO0GVGWheE7BV0kICn/hrGOXL12hRHe/zI5rSioK2rBd
RX2YcOLShGI/orFU8P8RGBIFtB7vrGjemyrBSQEDJzHhHHyTFvvp1YeiUOIxDgNf
dWrDI0akrvZclxAc47V6ZGCZBsXt83CiLh2LUjfiRgudDFy54jFio5N/hk1ghNNN
2hCQ6SUPKysM6P1ZISwKJGfgtXjlCIdUssnTWadHz8q2mg7peDEscBgNOvgGbIUy
/R6dOFBcdwYV1upwbGMCQ6r3pYS1oEO8TnmV4RVouPmFSuXBAJbRwtQbiT/oaqct
9vkmIbd5P7iJWNhG+TcdrfQGZS9lUii5HZ4V4NIefntW18UcpeOmnqzj35wWdDlU
SwwJ3EnTbcan0tHofRO79h48lMbK9CiaAUdKdyjNDtcB1NK745qo7MAOC4X8CwsV
XH7s9JuvMQpzPEDaLWSQ+6je6DvCekVJnqAU8zFPX6ts2/UWL7TilXOX0nxViHdj
opjiOYpAiGin02M3ANrzvQ0nR4FruDtHLNSA9XAY7el7wrUi+kr6dbNznBPzy+6f
+pnXH9hUqEUa+gjaBhUVVyanya5LEq2wvY5Ito9xS1TLjsFfX5Jit8jFe96r7ivK
EMupO4b/IZQrN7A1qFOUv48ZeQUT3ju0VIC82aylLAja6hUjaWcYII6yue1HduyB
cr/bewizocKewJbDsf9ljVTX91ve09kHMhvOE2ZmI0FhLUhK/RTwjalxZvPsr6Zx
5UWi4hVQMnduke3Gg2uJ7zVlIXsFu+60gYwdiPjkJWmpSnMcY2FJRp71wwYyI6eG
45x3w8Ydg+/ETruiV6XOjB1mPoEoWnL29EJq5IiCSx4e/5nr+Z5P08OLuogcC0ww
6dTv+nOoShTwCoKf8B1J/0ip6ILQApQHWH4JkkyiC8YFfvXli2dpogLGxS/9LNto
2tSX2+FHXAgzh1lsltCwmjZm48yx2ZIC8S/+YiNNfKZOe1n0lkAVLnCA324V+vl7
GQ2eVANdRfQ3+icCFj5N4evymlaVpTvm0g7oMkXdLRYT8W9rihG51MVIO2DRyTwW
7Gu0JpjIYaRSJnWu1OK/90Qrly8NKDzydkK07fR1UMOfoImLiW/u0/sbSn5iX0sG
Bmg6lS18jssMrzywiXD80jErvUzR7jXYxZykzU9I0Di8weFgIAD5oWJ/782jCuaK
SM13n5ImOZNbt0KGtSQdS9pX7FL4IsIPlWiDIhdA1OxerD+ml860WzfiNxtEb6xE
fGW1DivaSDHqfEen5fOvfa4yV5ZXYSk49x1JEyrwhD9rgf4J6GSkQwjUnXv1yzHw
lSfSF9ChDdg85VmjBtXz8aVpzbOR/m7/vjPyemflIMe4ubYFIMES4xw1PdB+mSMB
QYm364vc/WciPyIg4MARSzktMa183wj8Ncu1Fp4XiskPAxm/gz/4TwKjzaQV5dQs
ZJfC0LnBW5Ujm3XnWhFjYrPQaWkHLAYaSbjVY10jH5uzveDJJUM9+v81BNEQD/4k
iDAE8xy3cfJDWsPOHRNoVVB7UFz5H/QwJr3OWn60mqwviuMEpLEI0y+ruAJmrj6n
OzwMpCKdfWrtaodt29hVBA3xUA3Myh3byp2Ez9liwefomJT7Im9tYLEKrSwm/jV5
feyZnzqs3X5Uz1W7dEKjxzmpug1hIOk0qfK96qMQyuJUvv3xMXe9vvp6F2e9T1ZE
t0wesadPe+Fu7atEjvjUKMAmupHgfMZzeL7DxfMkzEy/LD4d9TRdb1R06LScICpj
rzwJyqHhWDkV8rsPrCfLfLMRQCMPM4q5ntnfCdECsbvUmJ2ZGl66HTmAysJM4kES
hInmq4zTN/Gfjn7qrPd6++nx7JBcK3eaI0xt8VDVmijp+90avAYg9kNTxAIUVs1X
4Q3yBcWKV1f5+PbT0IHLgj3Bz9690SORoT3mhaf/5FiK4nzV+Fad/qw2RTszVCge
t3BPpRpyQa9zHSb8FJbf5UX3xnri+M7VgqjG4PsUATtHrCQ2/uqzScSSTKZ5171B
n5bxcLewr+1TprxF1ljjtbk1a8r4ph9PAD2zSr1jJzllvKWex89r9IG1bOZiIIrL
qOWXb8N9O3/8CEp/VLzuo+wham1i4ob8dCY8JeLyHrtEsJOWLKK2Nv4q1ZIYkweP
MqN4UWF88aQ7ZP2lwRbUrwF8S6zHbWYCDhj849spX7j2ZLYuuhiVu8swPKWbhjFB
invmGoaUmwOCeIlSxTHVtUhffTaPw/WfIwXDFUjvT7UelcW6CCdc8LbfkFz7Shuc
BH+KoDoT2DtQDYFMC9XLCbeWBlLAtyQ/PN8tl80QJffRHKE4XIE1A/avZgwTUUt8
HJ2DesZVNY3aBNc6qgKvbiHlC2kW2O56blvL3MEENlEODWzCeAl7TQ3xeC2yck+/
UQM2Cg+Ayud5J+hVqUD6qRlx5XzpGiegV1Azonxri55aX90dzc2k/IvSHerfWKwO
OvhhY8iTeEV9w/hAsWTY+r8xK0sEgZNvfi2cHieDbG+lhKPjrPvyG+QZpHj+BFSw
dS5S9kVLcgbO9Ix7TIKiSoyvYkO/Qvc/YUzq7Q5RnJv4Q/NlTICl/4zt22jMPjKv
+Jw7vEW1Nf1lLPBrBzl3lm4/iD/37gTwfj4vqKvsN7P9J29cBj0UPZYhPfpblhfi
cB3ktmF0NN5fSG952fyp2pFJ+tn5vYdYeMr1Cnez7hhbuNL8CmAlLhi7XzSR51ux
+JQXqRMOnRolINhWLET0YVoykNGEJxFZD1OJDJUDAg4UtUPDHeCROq3LV3SWwhaE
UwsEYy5WetarAt3tgv9QGI4GfdzfKh+dVUeC70FWTeeesIPjzksDN1H5HVO5yMcW
3Y/GJf22R/CdKf2KMKVS8xe3pDN1GmnNDMqLGyA2F0CWMtEgsPkeF2a/Vunt/AVW
wz64BRuV2H3isjG6gI6vS9i+yRt7qOlV6B/nQBJWNdpHoIU1lUESExcOfqSxd/K7
ChHUqKLKFqSuItCtLKSOMVfMLsG6O+ojldbqc6DD7Fr+e+Z4xvZpqZH2VeoM6wRm
10jvlb1OI1uGoYOqNs6Udsg89NCkFYEE/U6piDgo+AdSGqSobm8/Iop9lgViMyew
H0DIV1ahBhY+XjjwrgsaL9eGPah7WSt1c4JYKGKCYL1kTEyJAlLENCFfE7ewT9B0
2asvXrKSJ8oYXtZR6uxk3sq3+jlxkiVyoVvyo2knC1sA5JlKwKobZGZymEidq3m0
VjjIX9k7jcu39CK8RDT4IgZ5SPN3vPVdxYhp6SRi+cUufrnciSt7v7t2UFzDFrQq
QkPIOdwkwcdkHgPphJZe2j5eJxkcBZ3J0j5BVwLWTB0w1jIku0WKfA2tXEm+LQB0
WeyMprzYxRv5YOtulJFmOFaRTez4lF0KC41Wg3RBbkkZuC2BrL3xqpb6Kg8mb99s
dy5NzoUMyKNtKNPInkqIvuPxJuDO7MN9TmUVYHR2GSD6+GylHDNMBxCMB2v/aIHA
uVJob83OOu8OFP9pwwwwBBembQ69Awbqeuh7JhuEXKDXyXJwBjbOZ6zvPASjk4Xh
/A2zU3gdYFd/+CmL5/Bg5jf06XGENsE1trJn1G1jZdZBP2fdYqv5rLK8jW/NWjRu
Os492TJJGE/Ri6izleYr9wgVNVpCydNBJF0E+sMbAylbhbrtR++fFqZzyyk93B87
bKXcKz9qSPR5gxZVlOZNHVO5m9TwY5u1nVJ9tUlZcreksUHiCi4at9ud/SmySliR
RUPwmgDkEY7RaXIEP4A4IUT2AET82hVIJ1de7XAKTGbdbVcJEYIWFHgLNl9k1gse
pXsX6ZatMHjO8dq++vpahGNjwQBVvoX129qW671abyogJm4uIMoMcMDf/ZZSap0N
La3L84IHCMC93olwwGuDVugnzDZJq9XuP0PEt6NAiWZ2gg/0RNP1433BEBiwWtu/
wHlg0vDFOSR6awYdjplc2cmjhIIdGTr1SSUaT+kjSx3AHmCeRQFwzN0qaTJgCGkl
+d4GRVwmTYVH8faJOK3MGuUx2xUWvjsNh0Pbv3gGv3BKs85Q3vZ/ewpqPZ1CY2zA
Pg2fc2dtN2JVAc7aZhuAV/uS7S/yCNRLfNCEs/XTZLnq81OmhCVm0sam3fWuNfnv
LgdiN+sGJ1zB35Boj0Q6qM6EvLVFUhrXYZmBd6YlYEpwz9GtDR+t9a8mfvJKEp7o
kZ1ioo+h+9EZoV8I0G1wNBKSh1/RS0tNAgGcQBXp+KYKgV7gFLnZKz9aglPGZ2Oo
BMUfYWYpIOUmHIHRkbG08PHo/IqlOc1WessX8WRUOfEfBJj9N34f2Oro38CU9cuT
Q9pme5FzMS3EGI1jkA22fuu0Ju5CYj9ouLW45TAHqfqo0IPE1U6oJpk3NbebQx3c
SQdYoYWF00PBBY6Pp4Ps3Ft/dKDqChkwhdQ5YGvSRpZCDLgjnB14YAoKA2IGUIno
oGtLcqPcbBVP9zccqw7K7yRhLw4/7sdy1iknvTqLB+voF4HwrUPNkp1gvoJ1OZoa
iZvVGJ4s1J7etLEOlxVkUdwshCcOrVRZ9Cs3wgxdnu64xQDE1Y8NHnuzqF2yDGBg
XU2eIux45N1NlrbZ2PIkHAagK3RWtZy65sjXi6bkN28RjkCpgGOqJRxvA9CYTty7
/9aSsliDpgvDZEqKZr/UXUnBxmp3JOMKTUck3gfL4xjYJcbIrhkPsF50g5QKcnlg
bzDI+If2BoCJ8NIVcogsxMl2YLprDz6GCs9OeV698onUJ/aVL3Sx6PAOa1e+apZD
9pq2nLD2c0oI+6TeEA2H+VYNvZyekwnQejds8wZpTR6EpPZduC5p93J9ibR5CS+l
s6CEvfv8xqv7UWm6kFzvjOpTYrFpT0k/ofOrGwqHSWQNkoFSpc/Qv9KfeQiCq1WC
6Qf7h9FX/3hJd3MmweTKwE9mVL2Us3ZtnnBy4hI5r+HB/+1StU3sHmqywqF3tOFF
lq5QkB6e9cjzM3Ptob5TlNPmJzzAy9oidBEPRawjwtMiskUKUwcSHIkg3iLrS87F
oehGAgNtk+iYUJoqYsCwQwmAj0DJ0bZjNz6SfTRENHDrOrula7M5oojE/xC2oHh9
s88Xnutv8xROc6VWfR/+NbpNLbY7d1x79K2182b6Aiwy3IsW9mKB2xSqIeSjEWnc
xBbCyI7TT7/eMfd2Zd3xSh9VrXs8qO0ZB6OVoj+SCbPLVl4jgpo2AV8zH2qEKcKD
a3SavAtGGR3+hhywW20Qg3czyqvNwrGAA6wkgH+dQM3rodyDTcWg4tQN8b7RVpZS
p4Hi2EGDbbrXKrqSkZohdMxCd1wea6YkXLVSEV7mBrabqz1TpyNWFMFESO9EnpBN
SLmi6N+B+v6OdBNgWI3638+RcLsiFMnl3Ay0h68K+mP7mjF2Wvw1Vf+vGA7qUN9H
IxKkGSHUo4zb1AI8aQlhcUsuOcovMn8ZlopL3qaM5SulEJ7fMcuQEPCG82bJv1oN
aLPOtPJC8W2nEsmissPuHAZU1Jck3uG2pjrc8zWHgq5w8qGigi74djB2dKzOMFdI
oOrEPPY9k7oBvvKrtp662BbzqeKEnenomAbkuXkZ0FKCdYliXzjVTdNN0qzTs+Wy
RRpihy6/9l4eKh0WWgCyaHpB3KddzK0qWlE2Iq+wPbwwnpvZaeq5H6JeyaK7AQKY
9LpCNAMSy6VzxDco0TYesLdV79gdRklP5wzXMhi4S1+3spRL3eg24E27KaxWSrJ2
yYAjNHExqE44pN3ln00Sg4YxBUV4tRHRm8isUg447L4rUEu6TLnW1zRVQg26aTdY
lDCDHsnDwr+kMi+Q8fjx8ZYduOxIIozHDpP1A6znEgWzHN8IEDJsv0+WpQSifDVr
6yNlJrNR2XTjEY6DhXEsm3v3hCSHr0An0pwcCSrydzYgXCiNEx1fx1gG18maQrta
TA16hBuP+0FTRK9SQz+Q9mWxLrt/cF1ZaXZqXldMa816XKNMxVhniRZks7WLg3+I
7SYGi2YSvk7Gzm0KrN4xCWAU8Dxf4ZWzodbCjw9aSvArpR84Skg2fqXFCMrjRYQS
7P/F2CSCnZB7gpg2HexfNWxRuJt6Eg8QMZp4rX04ZfTt7tf8Hn9Kw4k7lp0847gd
LoGzR7iSwmmBiV9W/iT9SyrHSOyIELe6SwfsMSb0fQoSdu+WVwdOQTHgsPK9ugQE
hPsp4IFefbnIBBymIXy/Jo7o0kwzMDqBuW+G2PwbKEFH79k+iUVKHKPwiJcL9HmE
oJUrpaUweeAu587NWS4SUrGZVC3HUx7Wywbo03JtlX+G2tckAWhNce3DnoAbByci
KZ9vX+BZ6YgG+w5VKrNFXb3t0x3LBBNYwQvaPQh3byC0ZV3tXA5QjEkBpLC156t2
2QosthMcG6kTxOOvIFI+IQZa4T+hvIsTSNnC4QRuh/qVJ/J1nCN6eh/iraNUxyAG
bDsbcPVjuBciFoI/aPLon1BYBSceyr8I193gjoiyYH2AnStzNCq+YnhpbFcp3CFt
5SQyFahs6vuLJCan3vmnsO7MS5p4rssH43ppG7abZICXNnVCOXGQzCUfFTyITWmJ
LBsmmCnuBqrCrxvFbd91aFFVjpp/wOF+IriTtNfU9qlJBZ6ymeBOX0WMcHmDoZKc
Sk7o4rZPpvSTVf6oZffHL5b30vKiUQoU/bUymFAydVsi7+D8EEDS6D3EXiY7ZiOZ
YrOOX+Fgz6KJ+MwiUAS8ipGEJKc0dFYTVNEDzS9qJ5CZmy697wa0JH+8BOawogm1
AyE+iG6wdxtdDa28d5b2xmzY+1LALgKgWWsjpDNAuoQJXA4Z3eQNgn09Bh35/fzo
CajsSjH+WsN05rdza3jNvDEZpo1f7ssB6RMCCwUilRYrSubGmFg0213W68un5hFZ
p+Jr16YcH4/G/1fU6sUbE7vqVYGtPGhRO44jgSVZwNVMjxyf9x7TnLbeoADRjqPY
fTex9sCfDNqEXsZNi+aidGJAAzM5D+JLwMBYbYpSl39xlUSShmnA2caBebbFsagT
/7wbiovzEQMTN/L9fj/ResBHghcyxNppLlFvvvKnFbklH97N8y8USrxUKq++HXNU
TzB499ucWe+CNS0X9LW/bGou3pDhmo60hIBTaOdxwWZb4AD+6YNDBQUUFdCvw4AX
xZV3aTKugJYSKxZBkmHx2ME74TMaxgM8/FVYvWwoQBg3IU84yl2KnIPEMjXFPIju
aIxE8diH+RsTPoFSaduhdbT+T7Q07UgGSZDyZikuU7syfV+7br7XV+m9UYxkg8NM
TM2KbchmY/D389srkOoGnl+U3q/iVDq7KIADyubktx2ZYIyKQ7R/CwJ0vdHNa14G
FhxQEs3h5tKeYFktaOZeOZBFNM+ZWRnVR4ao/s9DqsAc7y2zK7U9fZZ79wkUfiGD
Cj4iV+8z+a9IOCImxlC+CBpPv21VxsC86E20C+VrAY/iYJDHVyiYNQodvuyBL8ey
AnKx4cF9YfKV9RIkwQPQ4Dd6khh2k6TLYnJPtmGVypY4a1qhTZpx+9IW+Antfsg/
EIEfpOTrVsfKIe8xq+cvrWBjTpBrxvVZwAAd+nlQ7QjH6authrvh2362NCXqknfF
JYbEetEFVeigF0pkKYLZACrqHlumpE+MJpn+yrjE1Cg4U71WG6qGg7SxhUfyLg8s
krOQnn9uLkZxg8uhcxrhWTkXLL/UY5D47J/mNTqp4eKcc5M3G/7rb5byqCUpEzjy
ZfQfqBt5QUopjiQvjVdwUeHOhsmTyx73/XMMHGZx/1ZbBa5CqHrvQfHudor12gMx
lQk0gqkcIWc9/8LLxsqL98V9YbMDocF/xASszT5y6mZVl9MEQq039e64ttj+MJWJ
6oUC8BS+7nGobrN4spIkL7NuChLGgdXeWulFjlCl2dh4crPnHEWjSXYhDxKb7aan
RF8NHF2aLQboYeMfvvwykGCZ63w7JTWBCmalM4DFQKyxavXIfS7E6La54/0bdhkE
JPDciLJsxRXrnkt3Eyd0rINMRQ+lQbe1gK+3r4cvOduUOu4odqO1iLLgJuTANIvD
cvXr5MMM1y7iZq7zZWrZktCIo/9A2oy/OhqQggy3zhA3is88RRApzi4RFhGoSXLc
ebDRPfAeWagM3qXZPKKLU/cQKXD1eDi2kjcIvhC5oSm+/jXX+KYfUOvtZ9xCeFhF
rkE/pSGHjPsJplaQumEx/hcoJU3TAobyZUgVsVW44yck3jbg+HavDbNrEjq1xzEY
rIku1p4Ij03kyGj5N2NikqBrAOiIUQixR8WazV3kwRyzpqmsW29l4RVYRj2/2XOc
jQOPxgcAPRqASo88oUryOGvp3JXZTTo7QBJMh+7W88lnyMzQHRwmXBVK7Gq4fBp2
7GBOMXexu4LCu+3CcaAmeBp3MndtEFuplnNoCVRb3r1OFfSenE914Gm7FdqM1c9j
Vu1KX65UAAZcmTwHgVihLfvdkGQ8SmYHUa8JBydTMYfGjbWUSDur1nGp4C5o6Rf9
dkA0cijKIavPNYHwbrXsyQpfTK1i1M08pOfaVWSLzP5INNne510rZ6ab9E7HjsP6
7efxBG4t5cm8MkcYAE6/56xs2xXOA+4BMPz3sdAL7edEYM66vsEy7PimgIsMFA+Y
BHiwO/oPB5tPr9fYlrrwQf774Lq9Lp/fN56oo7WF0Xx9HQufcQMaDEYFOTiyVPUM
nJu8vK78JrtVU355I+PH6XX3e3imOEnr9v0+YWYyDjri1HIuHU8ZAJ5cey5OFvuC
8EiOoSMCLhNF8APR6NL2DtKvJFOtZz0IMUEeuqgLF7hTR4PRPbT/PXqxPrw1ExU/
4HzK2BVpp9FZNLpBV/MDrAolU2JZ23SIcPVlyiLwB1XkbVLmBSxD4Fsz5hYLT5g/
m8j8eKCNiXZGmGCeDVJ5ONlWebz+gT42oomqkWGnVFKXhFW+/6PC0uKbYUb3SzAd
nqBpLmXsHHoObeSJJSolKtYqQpppeYgpEJFaLILW/obFhmOfYziUrjZojYUV1yLN
6JS84DL6eWBir/WF4dSAE7gvRBAUkhOv4D7pNvmv9WdBvlMLkszMPFkFjmWyfat/
jxppuY52RCE8LKr1UHhIp/2Pbbxw8sMFaH6FwxVc5zsVcE31WzUTd+uhxKTzBZ9I
lM+AJ5QIykpJEvFdaM3B25Q50CASE4QygiGqiwFPmkN3pD4k0JIWByabd9OXNMlc
Z1ns2fem+EsnoiJoraLh5X2bcO6B/r0Zv1BI3Nh8TV5Flv5d8d/WZRCZn7R6D2iU
3dqRMEmDWxW+gsrRja4JFyIyY0+l04008eWjg2O7k3ZoDasfDpjHyTjuiTFEJjcL
RUMMh/w+nm9uL7mO7d6KK2I/RYftgjXkAJNDPVYbtlVBkZd0ms8NbLlZDPT7Gw8v
sK4oc5GDOi2dk6G2cAcl/+m/No720HvpA5YBtum/u2Sx3VD+pp8m0Dk0ANoZz9sN
RpSSRDMyBE5cxp12b1mhdqu/sLGuOtnlm9ONyUY93TFlP/xCkv4P2awTgbxr61vE
nUh/we+/LTnnLHKjB+mu/myVl8qcmgTuRzVt5GD7MAArPfVES2xOex0t5HRq/37T
bHmkMZNf51NAz8iNeGI70XGhqKLeV1DZt1g1rKnJ3H6Qk/rU1BhBsaBewHAuKt46
FFiz268N2DM4DHOY+ncI6spKYmRWYqjdnzs6HJy4YfUeoMeUbcHEfhsdMPGx9wdZ
ufvmmU77mIPeQ8nyzpwHyuYlI7n+nbU5QggXZnlVxtnO746VsoKAsYxfqdEPOQ3B
4q2IvpiavrpYVTpDhrpZaGfbaCaXApeK1qwQ2fgjCKhJQ3+pz5EpCJAQR/B9MnI7
vEIE2cI5GBDkat5Cq3NyXW3HxnKS2ehE5ZnDb3wrNbX/Hz5vHOLX4VFO/pC7MrBT
7kF6v2XUctO3tlFyfJqpryGSFU/k9Jk4Ga9xM7gk1OCcS/78SdXEAecB2e3UNuFj
+PcvG8eGjwE7BF5eMVhJg9ftOYxY/a2uN1YQpmqh3RTFZOXFN6yoK9oqxFoZGbfF
6t2Rd1aMvpCi3VKpxcupvQyEJmE+8kM2Qs0GkPCkCQ2mPPKHsKE08IpG/vmCL6lU
m2zk5C7LlcHTooGkv0nGboCYer1MC+cmiTCge+H+sr2IZw2fcAVIK//LeifAjeve
NFQ7bPNnGvID3V5gNiUf9qfy4L1yTB75k0eVVn7fSKEg+D1oKoTNEpcctUh0sOEV
soOfoiID2OxTXSVUoiSW0U6d6ugLsYCSyd3f50Eh0KdqC5w1NKVSCdmsXCRSZCEv
sk1SpRUFGbRqbF1YPxDEkzzScDN4HlIyimWRHAWoQF17XGUSZaRYylacJOYCWC0V
CG6SNWChjTybQvlj3S/WTIiO3p5kjLrtegYcmHVk4s4Dv0eku4ZirUzbk4fgc2bq
v7ODgZeFR0RhUubEnfLWY6pNMTLjctZ+vAvSIzZbF7Ub2vl3ys+1DSUVQjp88jK2
46DasUBgzyt8qx7t19Q3jJXjFAILFE64CnyPtl/HSe63lNm30zO1h2VEC9K4o8EL
dku8XjgT/R4CzZfkABDLVyYc3XTptmVD/EQ8sZQN/UqOCrrB1RyTJEdHe+xJuPMi
H9ULWD+TUfqfXUeQaak7+JAFZbwm6dcuU2cEEtx/5zARNCxOeXdCKw+nods5R+fw
egIKwkcWiC5BRkIDlftWRnFS7ZUof2MjV/2Zgr4Sjlnj+uY+bLaVTp9M3rH/jPF5
qTtgXoJGCPE6UN6DGws5lxmZ4y0Rbq+fhodJ9U1TKEe5wEnK1bJViZX3rkTbYyR/
ZfjQ21ekYYrvQERumaVaqLxBEqnpwfpCHGc5Z9CtQHhO1AfAmZQZtuMiSCreGe/F
7GwuugSU/a7WPMpaxhuENqJMHhJlqNzqTCtLjgngVPotOt39fB/rJBD4ry7Ioms1
auOAl/AgPJukJKeioB4+mzRTjZwkDtf4ACbpRzG+5k/VEQAcFveK/Clc7QhapNWT
gdge9CSSd7q4pTmt+mLHfiz1076aBB129hFnhSNCQIAV+jflWD3CIJihUFUkMFD2
Nsj/JYfpKA6ebEGRdHyymUBLwvLDWBRUz0L+C6NSfjcORx0Aw9omKCmS8dDNYy2+
674/DU6Bvr3yJdiVYGhGjGr6QxbURKZSkFnYY1QVndWqKKHyGXnjXH9swTzy43LI
07O9tbojancfP2BeJoeJUdOCO/HhP2IRcSihwgapwDUB1BaUIA0xnz5PpAlxJg17
mjOYySNdaWSJKZVsIBPFl8ItmzYjnPoc/kZlnTElVi63xd2JBq5mH5h/tz2l8ibR
CGtfHUa/KnedpP1E83gvklHfwnmpUkTMIGOEwsZPR6GiIqm6C+otdMS+7YfSezNI
980pMNcdoMCww6LlTBqD3FyML7IUOjA204sVDOTopVZU7HAq99tCXf439j5pCsvn
nmxr51qCGk1pKMUJWkyaXKksf3ACnsnaeHDsJn3rHITFiaIWeiE35deTG1YlyHG8
RelN3u5TAhnWjTKu1itK5vnWWhyAxArgZ1IzG5COBmShLwQtK4j8JVnpyPTx5QJ1
jlhv+qP1fMBOZJommqYvG4LRqbk8zBOMut6hoq/npz/opIcXGM3189sIWCs8Y+bx
YJAvRxQ3vdtvu+8kOHlYZKv+y81cAOrWjE32Ke40isbTmbxSj5PPzJ3TC7irmb5Q
HUvJIkGenjPPd0bXEJoNlZ6K2Vcct5q9J31plhGbtqdkNbW2Zr8A9MpBnviIGLXO
TEOJmg3SvzWaRmC4aoEExF8l+w/o/l6wsWIonYGclzA2C52lj/ocUohUoqvV6M0i
gm7lsMj48+7d0V59ul8hvSBSBdGAoU8ur0gdC3qiXL5kRdNMwqVjw8EFBg0xCSn1
uyxTqrdP2yA92zSGP8Xzl/lfUTo8wlLMx0q9Bz4sZd7vY6FeXGw8H86uX604Kv0d
kWx42xsALvdhUtmPwg03tArZ/FasuRnjbP2OUUJ2iEuuXxMrWA01wbgR6nkXKasT
92xfRxKdHvquW4kezLYWCzt02rzrs9vad87cEG+9/Y2Nr/4U26YML4zTels0t6Fd
z17bDui8s8/JFnxSkfp6vMNmoSL9lQjuKrkgz0dIOrfftLouBZ/WscML76jCEmyX
dOUmmHbk/oKNsQ8v2PagOVGaXhQ5YJWbX6BePcfR8+6ZTiKyi9/8l8Ao69sBUoLK
MvepwGv3GYztWxeCUu8I0brZvqr13AaHFak05fRXIX6gqHBajDPh0CvQCw+czhXu
rqJ2ZgHbun/j0KnsV0hGxyyUrFhgHvbEpuaQLcq6LSOK/7shBzVn00rj76ayQoTo
H2anTSC8hwVuBHpnabedTtAnCVPYf6xc5PoDTBHuK4bmpomo4d7tWJrwE70+WNoY
KCzV9A1XtaqNNNtxZ7iImPz4VUGK0DdbAGZmx9RI4GaKn+HaLk97rEoh90orpCoT
Cwa3QskukBp8V+0/ayFtF1xC5R9KMr52Lr5McWlylPSa46eUc4iVZZ3yBMfOeJu/
gj60SWLJjbDIUZ8RuOfJ40j/fSO2F5yQFCgrP/bq9xcs6NBBjkh7HLQvN7oKbUhI
rGhqhJ20dxoTTNLTPczMaocOFYbwAD94XFbjtRFhiQVUHJwIDH6QEz7AK4F7NxNS
UdvNAN15XMDtQWMWDHEp3dCEN+vgV7VB9lJSOAZR6wNZO8jgNgFQlZlQsaAD61Ow
oxUkN6CGuS7y9U/Bs7el1AnhG50ewtBT65bv1YLNivng0VIcmuLxH7lQsMZQrgk2
eUuX4HGHg4gsxDqm0aFS0H1rd/L+d3mKTKKc0atamNHe2HsPPSLnhCncYKRd+F/u
CbvoR/fe/xxysG61LscghILXAhZ309DavsShp7gi9LIOHJtFN/yjHTFyVzBmUcBP
vKg5obZAXRSCtXLM/3yze4kjhgmXoV0HZlMbSHxqVK6hEiNnZcy0lJba7UcJiha9
E3VT47e7Gg8G0i21OFXYCjQK6g54kWM/t/2CwNKdibbP2t5/AYJy49+9rI5PPoYp
4kngcL9+CDO+IebNvWixXCmJVwSrcUyJrdh3vVdD4lv4BkgHfIfow15f9IBUZ//U
V2h01jA+tTaUwgx71DDEHo89v3m+nSmP7Z9jn3lPHk02XCNA3lZ3Lek82w/z7Tsc
izpWW2dE2xYBnkQcLMQsRJeJ5BM+9Ok2jzSJY3xkvtDwTfLnKV3zdiXi8qe8+REA
rQMZAQJ4+vwT2m97iRySEkfJF0l1Gld0eceFTPP583TYJHd8RRxDnZ3RttYQEZ+o
oGIo2Yi21Ue1VjwgMaNqywJ/ZinQTtKfpPowmKs67g6bN+7eHUUmP2XzvDMVdQ2D
fUvNdkWujnhS3ckb6iaMujyqkWKH9Ts1nZVvO9ifJpAGPcjXA/DOM2HR/VOAmI0R
HCnjdlsSS2R76D3bguIADKq3DrKp9YcHCXighWy0X9IyYbt9N/yY9I6zN0BPFOWt
0UnLr53vGsiYyZX1/5w8HxZGo7BnimUQ3o0a9QJsPQ5y3wu3Q3pyuj7jovbtXXZ3
Co1EVNeK46lXYTnN23+K8RRkMn9+RFxvAav3Q+Uo3AEjvJrKJ2NwxzPkUoK2AtSl
prvlrKVjzyrE/k4App6WgbwizZAhyzxC2t9lXyZP3ybZo2ZrUTQ6hE0C4tTiAyQr
vk2bLYFQmR+mbCs5wPHVkMDanE4AuIKb4vuX6Bs3rXkk9v1Hz3/HerqU2QiaBpQw
CCP1xSz5NMaSdhhWvoidc5PCrUEiPjFra8XZ3hbXbXxd0lAUXtAhJodv+u1eigXk
ssT2HgNGd+itmNQsTsmER/mxG418dLN1r5osWUDlnTqzA3DiiOxBvIqjcCPzXQL2
uVIiVjgndtBYF0vgWIH4OBuz3SZrLOe30kvMHRgkrgIE5ytnRR1ovFiGkplPYW3h
rZxT3u805UEh/aTVVg35HLIyin4bF8QkoTQCzHkzQBVVk4Ffxgs8RSvy+BQUcp4N
hS4hR/FBtXGHGEH1yjrM8GhgcImX+Wp9ZSQ6ThtJerPoogQpOGcWzD+5Djc9rZdd
emQy4Gd+DDId7C/gPRr+kBATww2T7qA76sPPnmt9XSzfVkdzx5BYPN0sLk8XIeIE
0fE5eWMwqelwjJ7RSyAg7cUDM7xdA3hLO6KCmCeeaStW7HYm32t3j93FSzyo0I+h
r7nQNvIPWansmGsEjNYe+BSNkh9RGKWRxlGEG6MOBfUJIIv1O0Z/ndk+Bm+SIObT
eu0LiuEn2NiGDMH9Rd4o0bIGKMa/vb2LmwIPAerwM0s55+OGmVgvhUYmtLjIfq3J
e9XKy9XtzEW9hjJbrx/5aJHUTCy3No2jrVQG5ty+mF4nKmvsbe9teBcMt0Jz78G0
bSCpUzwqsWpPs+y12Zf7IS4nWYHL30qnAuYpjVHj7ObTg0MWzoYcfY9DULW25bgU
iHruF0SFTbpH+s2Qfic5Q3IxpM8azybTLsP9dBD41JqTtl0kPeAJ6+774I6Mh5z0
uKnYCvumOSvOU7uKXoSKUJtzDFn0ljk4c5cixpYxDtg6Ve5DqfL6ZIF7Ys0YQf2k
K2JDdi/n9Q6tJbElY4dmANVkEjZ+wkUF2oPgpNCTnhIQBRv7yLi95aNL8UGGqUbw
1I7X/ZHYLffWUcernwN87BRQALqK3GWz24kBiETJAOeFAiiUkBo6MxhIKULqqFUm
ZgPDHUNVhBU/iH2q6yjoG7yJtQnRDS33NoXJRlwrWwnO3f+LLEZpRjhGqtxpIPx2
3kBy15YKxVkRzHH8whVHrEZx2pTHhA7R3hU5uY++sXEucpT9o6VncuGpFp/k+cM1
EdpRNjzjM8h9sATO+Q2gk/rtsdMk+yc7VDboWWEZc2isTGtk9najmnq8ykOaTTBi
7LnK9ye51leuIyZDe94fXe8WytYUG7ZkoGD1YNacQR0/EF1YoHPB34vaqH0Kah2K
Y1vue5H7gCz6Yn42VkOBrq49J+KuW0tn1ZKbaDUWHZT5PKUUuO+rY8VZ6NYbx77/
+sZ6HPk66D//Ce8mEU7Po3T4hTZPwe2OzowEfVf8o1nd+wDnOYB7sDKL9vo5pXmy
YHu9lwq3vqgpnCn7frgaI/KLXvaLzzp1oYrK24NFguRv+F1kzkhjINBsyl6qP8dk
4q9oNNxuTZ5SVVfg6A+MBjiaEDbfBUHJjdMsgW4/Ol+icDxfQa5566RZHJvHt0QP
lyktxz7xVa9Vpq7q4V30H1Kjz4bGcDG7Wbegx9ue73EecbYO9KnZ+dHVmEaYWT3D
S5ZKuU/AyoqTIA2wWBlr5IOhOxELN9BM6EQDhED/uH6/0hqhOSH7GMmjWLw8PCgL
xyGjuDYJYo701kFiMP6N17A1kOazzPauceuRY6cql9y8pKV6DSf3cNVE34vZu9J6
+8KZ3R/7k3rIJFjMnonNlC+HvTbAF4Cw7/hgyuA83WDnTENV5NYOVhnj5DWMj4Yf
cjDLtaa5BAUrmSp8ZSW3NR8SK8b3jjmQ3Lf48gKBQZtuipGr49uNV7e1LKjtLNSQ
Eu/IV5yX2lh9uPXdcLR3PFfmebMLCv9wByRB9gxUPnMH25w0V5ihIYDsZK+2E/Ll
IDHwc/L7JTyKk4dwxAmEVL9BDqTzq1aR/45P+Y8fOKaE7Fol95T22TMO5EaUejwF
5WE0wEDYXMwS03Xa8IY2ZpQZzd4ZtDent726OT9Z8s64QmbXqHVaB/dtj8cRNl1j
zP/iuz3RqyLEOWldjFERBwmug88t+hwSwYMSZ0YRtL5fQTW05x3ry65QfR4iwVRS
AzAvFn1+sg+RHKRlUhemPeouWlcCS2020Aht3ZeX1POEuShiqrAzwsMMJbhKkZ0B
JZ0cykMYT6wrGLzW60Ir69skmWih1U1b/pyZa8Q5Mkb2w/b+rkRP3odGaOlhDo1l
4W7sL1Uk2SZE5zgOt0ZMLspr9LsbH7435PeVaeEj/AzOD9IzU5D2cCD7RFG83w/L
J+B2j/nt5c+eFWyfY4t520GfpeYZZ63N18aU7/wxSiYprWnJb4WprL59Di0+QQDZ
C6p2VBxS4QCrlW1hyjr3FzgE+BortQKoWuEKC0BzRWXx9rXdp7tpltTNYhVSAZKE
WpT7XnGQNDFLWwwgqafKGw0Okj+0U394/tLDoOhqwnPGiIHdTvXFeRywlQ1PpI8a
zbyq8BBpRxjw7AshkehfwtDV+5o4YRgWt2c2F9Fu3FrGhHlmzLq+ao70B7tliocE
g1K2WmPeVAdLR+pfXzu9IAdlVtWI2cGSyaBuwhlx1quw6RH7TaclyEEGjI2Q0FWS
ECTLCY9qZ3RDwEYdzoUnO3+1nWRQmur4L3l7+h264olEtUYdoUuRwr4QKrmkewwt
OjRGIiGLsi+QoxmaHsOG5mVWGBYkwOVVRl3AST9BKqSXk52WFbsn4WNlYy+ShCoi
wrRaUSjaFnWIJHy2qwl4pNhKQ6QaJOdQoWMRMSnvLXD522WLla2ASn80EVUbdsjR
/zEYsLWZGBWQctuYmbPRqQxt47pvo4fc/PZcIKN17IIgUMbJ+D+UYq6x21VZjAne
brNQIWT9Jy8hqH6inBQYnn2g21E4m73bTlg1jehMGO/XItD7Kq3JhlNBpiPStCQ5
YE9OCGah3ogm7i2OI170olFYAIoZKNJw8auJT3RLamhNEpB7MpPzs+qiOnuwk5Zg
1yZjapUTr0yXMlSP5x7bU7ihC3vhEPsV0Py7WNLxaQFjp3j0ToZyU0Ydse7jNy2G
349dA/hRH0mwcSDA9Ct6xcQc1cJkc0v5XU5x7n6Q+TAqYpAENLP2mcbT/3/spvN1
76WM4PodNtjFsrCYnysmv4gPgZQGrrHinYO3qO4jv7uA5HK0eJw9zfecTxDgdTPr
v2Ix79pKF7rfL5kNYTwZvg02l0jCiJDQ9BU0P9cO0f5hKUcxh9RC0BiFybBpYQGs
hve7bU7yu+ZR+7ha1N3BJwNwlbcj59Qut6C7xX9LKy6U70jJrX1j5DU1zWqupOzJ
T3w9UM2vfMcBCLYf4kaGiiSv03qxGm+ottG9h7GghVyc+iFhvqrnwcsu8GScnjO9
xYmYfshvSl/UJkqzri4mdgX7FCRBzuezFfc4hD22hsFpjLy+ZWCNmjcFKQNi6ivA
q9oXKoUBIaun/r62fBZpACDK4L0gr6K0aMcKyjTYB3U/F3mcQbUKZpaNUkfTQg1T
DbleNhcMpVw1tXsBQp15Y+FTP5UjzHSyrt1VQJJJhGijBMHKQeuXKomVmsO+iBED
AbJhO1NZTdmQTDrlA/cyuDK3ZpsMt8/gI5BufWPLnw2Vkp/3DtloA5DSuh048Nlz
64KlPMS76AC2AEgezByEzXjC16yUQLHJW4NGiAjvX3078m4v1655k48WpGzpJ+Kk
Vxkm6G5VKrX4Fx+PfHFpTW+yYlhPWMsN09FdNW+N49xqDlcjZL/BAmDCuxD0mI3P
uVZmBykPshh66VUnqvI36wBlxN88IXMjFM1wloQtI/W9uPc588ShPMnD/9rbTuJp
LWrM7FfgqhOkspTq3StlBEkBmbSLJvCBeNjsHmBKZkShDrv1tiABDV8Lv+yWeMCJ
CalHQtKabQWHEKVTp8t2l1uwzExIjUnKxO2iSOmC/szVlDRvRm7l2DX+Qr+EvsoH
4yhE1GswuWQ+S8Ttk8l63w9LXFQbd8XG0pThmu4iQa67FHTjTGSaF0xFFv1nXXBt
qNR/GG9tA8flUIzhtlTseN0Bhc/EW5vVlydX6MsAZiHofP3jXS6GYAQk0qLAsRBm
JZGIXAyoY0OKIyCCrUeTyReWYqqd4nBLUqXGIOpCfm8PZIbaEfcmd5UWKtzyMTpx
sy38cfJffr6vuAxVwL2/BqOp0NvOhPbTEniYW/xDtD6dc2r3ugazB3k7XrQ2t1sw
KNVHx/BOKN6rXcZVo3GqlK2q5TM9rR/r7rQRneH9ONtijZxZWSX1Jp5gXQdR82Sl
4Yuzjoez0Q09d7b1VRuyldEm6mxA7Cw/q+wZ+HfU+B5gt4GrCkLYTlbMDAKnLcsR
VtdthR0dFbzoQSlHVJExUQnaC7nUTVgqgiW03hPySv3ircdZ98O/DPtP8O+AL1YB
GYlAWkSmZFn75c/t5SpPpeGSOixKRzcyBvSrGgXYhDrUPg/iFQHg1kElA46rplGJ
0s8Pyad3n6jtI0RwSLLkyzu+XN4+Qh3D1OO8i0rT6pZclEZuiBcPlP3N/9mb/a0W
mel9Dw3WTprQMJk4l5G6HLbM5jjD73WnFBPcQkagkGujoDL2SVzdDnm3dp+1IB40
oPlBf1up5ZwwoP5eJtSEj7xAj9Nu3lsCtOQZWKfVLPh+pFV4kNdwVL7OBIq+KhH4
iZeLuKRxYi2IjHz7bg6vQPXkLCAJdS/aXCpLw/qLbg4UbKEpgPAcTirKy25/tKAf
Wa6iREf6ASYsB+65W5bfp63E2KieKluF2PCgohd50Kacohkxl3imywQ5qzFewpQ+
cYqF6KZ+1/HX6/+1gctqPw7wNi8qAmh8ZtrQcGQCc4yL2YbzANl/WknHSZ8y+atc
+5NLfwjgSmYP4r0r166pTB7Djs+OW7zkcaI9qRHnhFqhaE16gO3jyydaZ7iSufaj
VvF0q7ZvODh/ogJ+D1lDxp1Wg7CHo+U1NdcPVj8CZ4qymNY7rHhXkvJ+g6UXNgGS
r+b2qChVaSokFn2vxOngcZLn/Lj9Zq3kyzk3Kp5Iky4OGq/WvWQrV0uXJyj8YdX3
3wBhcXZZ7f0mDLjhyHmEWT8CZSTOd0/goY6l36A/K49Ws0PWdkR0WwFWPhK0qtA3
+3bmvJVQHMB8F1F96pO2tJpojFRGabZFpp50zDO0jArEzjnNViUdAZWoAlrAeGtS
WHmz1R8JYBFvycXCeF6FhwpeKnhhjJr4gTInSMvIci+ZfVv0weHjWF7fiv/tnnNN
vXOycVYd2jiB0beyz/1LxmV6BE7pt4r+7V+qUr8H5SNKrgqF/8DSjks9QPhZbYWM
NIKmC1k5fix8UikI1pA1FexVAVekZGKyIKzXpOWIJBIbpDFFHcvD8GVO9ZUdftNQ
h2O+N+BN/CMFeNW0NqqJENW6AJtrMkVn5Y7yRXT9vh8IQ+FSf9sAcKfy/sA/6LgB
HlQfbK7aHy6WiVoLZNC05AuYVIeHwr4I8/MskqN2+K2SKUdGyHgv0qVvAzQLm/Ns
Q7FOVeEL3YdEygaLb9m+C7ql3f1Z0x+S+3w799+8T0owCrJVwmHL2iiE/rQRYJtI
DaPhvoSMleWUpLe9bxAm7eQWv/iKyTOYBgMwdl8GY+yAZauzxMYzJWWlsDchqMBR
5UgpQbP8+b8EFPvtYF3bLHpu5M7ACwStntyv4W4AR1PiKbKLFMTVICExiGzSzkp5
I7fbJDAPudIsm4QzyVvYU31BW2V5O6ojE1AnQgJQqr26gH/KcA8taVtj8Uvb47hF
1cUrMyOVbfwblAe1Dphjx/mydv0jbEqDDKKij6d932EIMbzj+I1TXMDi8V9tG/Ie
pixuh1ZcrgpS2f/kiwdW5QF8PS/QkMDLIm+pEVZhRvDKu9ZZTBZxt10PXK7n9iAg
JjcPfuldEZ24UcRgi77HjMeMFZGW3x/k1wtjkAg7F/kNOpdNswS8DednwrJ1LXNg
UDBjuNsQajo/a9/XXCahsQbgQgkzTad/VSCSy+YNYvnlVacciCvGCuB+Dy5k+MwO
Y8SLlAVPyFP54Ej6fdXOYWeyrmSspq8Lx8IwoI25xgGRrH01kdM6LhyUtGr7Da/Q
vMSHzPpjMryIADoAIHjDWd+0gZWYb2+NdvbWtRUU9/VRVnvlfSapqAGTmcxMQ+BD
tHbQwOn8ViXnxrVD3+DvgBslUoccJ3NHzpIoUqlcTm+iSB0pgM3OugnhfOoQO9Wb
hrMwVFyARzYgRXgmXhwLGfoD2PMsXkSLNeWjuHQGrZkeGhgDqK9qa2ylW+RGzlQN
KXrVGm2ehId5aZ0uglW39UYahTDgJuTFr0+ljAtbVeIi2h5rdZptwEaIPPKu1M98
YPiXBViGGk5a5duHQPbC5zjEVnHXbybjO/sq7sdJqJfbiq/3DxCNdrHh8pAuOUWo
bzhkl0qldLy2QSdv5h4rfsESLl0fFpMkQhvTONEXp3b/xXX/Xn3LKQOKRqmlEXRo
wyamLNRxFklA0Ae3Wnqz6VCbRae65UhR/S/TL5FzJbxtZeMemPpVIL7XJl8CCxK1
FwV/mfJEZ4zhZJLi8xMD0/LUjyFthdOn62Zyk2SWPTaJnC0BvV5SDpWo8lTJ9w45
AFgJupd/NfpW9yeD6fYXc1TyOVpAt+bfuRAWBmu1tVssIVJDWn1NBwLarYsbkD0d
nMvgZZ/OKHj4p4/uCPc4U+5PZtZ2j4/g+SZGKfvF9+qUbAi7B3mcyjjclYn+xi7p
JyVOmUM6gYqm4gmHmlo26a1QKbGFDJpOYR5KLSIBs77vRHqCTueneSSHtpkxX8SC
X2f8ck7MmLEtKr2pLQMGY+gXuXcgir4e/nQ4/l7158bKR62vZghfU7iGLm56HfWV
DpG19to/fRFwsr7eDJh4RX7+sdN+pu2wbFDRu6sRx/rPUk71hUM50dbbTFJkRpHL
59C7MnEtwycH20uhNlj/+XgqMIlzF2dHMdiuExhsm1UF2q0m5LXef2QbPFuqxQSo
1aeMCfEH5unym8fh4Ae/16D1xdWPsSL+OzoVX4XQbyt+pAs3eO1Gy4LGVdfi3W3I
LelEWHavg7KOCr2ZDaW2WT7ZPC91X9cgyty62Kupm3x7UJ3ypEnMAAYFVqV7d6+B
lR/yixQaGXMglay+Zm27rDEWocQeN/8hm3Tdbtek8P0aCD6v980ZZV944W6J4Jf8
UAtypy6BmyKFsfFDzoBLAeNa0e6z9HrKsSl5UVkUGY5FLAMYvK48fubxeOE/nBT2
ljstaMFGrVCUzNenBCDi4plOLSdekoX7wD2koZAQbPpMTWjWPwoqkXCS6mUSgjVb
AFxKs7Y382wHBwWPvG/b+bDVhEaG0rSjCSxgNL2m5MEGLuSXOFTh1BvW3Y4RsD1N
E+A8mEBonIIX4xEzT5d1aKYfPzoo8klFkSl8Z0MDR9rFZ14eUF8kHFmcfZIU1WoZ
BFyjWoiL5YwDXqH/JU8ULQTR/4D9kLU1bUt7IW4CMwi0yvj8HQJ20AJDSnIWjZiR
XsCW4pElLnsxzFa3P9dittz37pUj7KmYjWJZUdsXK9iWWC5UfcCjd9ctg8ZwBa7r
vwiPkYJACq3CjTQIgPZ+hhjMHgSYegPauGOICKw+2SFVme6Ne/0s56/kw6vRPFaP
qECn2fIv1maBfAHsGM0nCK8ByZz1ntC4g9sfMz0IkP+KdJEveaAI1Sqp0FIVI5W5
ZejbZ66in3wmK4T78nmcjrJet5kC/2Tx1V83aXcp2s1ghNRn4USN+oFrZ5dkZcQZ
2ByhvVprqql20mV4haYP6HciL/T9/pplGketdX+OiH79kge5RPj+Vy2qaV78q9Z/
bYh3AA3E5NrDvs3znkYnJCnCnOwrq5cEZlx/cC9UsNrrX6ZhXE4k7hz/SWegOTjw
hm7GKVSQypcyxVUcjqvyagQWp/8jbfDHYA9mrwkOF5sIWixvmNCZHJd36sVhuFjc
QbOuQA6iRRwzn6NruEZaOO3ikzlj9VaxurvBUhHF+d7qv8YtOi/rji93qyjPn1ef
YLxR9HTMWxXJQ9ez5iBxQNJ7gVsvqvDjlW5F3hvLq7PjC1V/Uy2Ng75L9c7nmOdL
bXFgaSb4W/6MaJXUIDpPt9p//CpxIRNFXyL2zMf25qxGw66FXsutqcJcj+fW9k4u
69g2BJPu0IKypeg3r2F5XUYACpMfJurPPfObLCdVJySkjScit3SsS4Zc9nQeiV1V
KLSjxq7soh/7agW2RdNLhdn+RIlCEGsA1xLyRKNSAtEjCslR+sNlw7alxddhLIpU
J4tnP1jw4dt5xupjXfl7NooMlBMqIfp0Fwu5CR6iy6D6GV2/lGgrsXv2dgXSkIQa
t6DTIl8NiVo89bSpHdz9Gxqbs80skQiv9o5F5FTX3dkt8peXdPOac+rTDkfduD9C
/dKeZyfE0PC3RLock1Fb+OsbbQAkeI5FGUSOnb+123T2jZaJIyKTK0hVxAN684uu
EMNrrzmUC1jyIqXUv/wP9O17gY8rlWDweia813CtMagG8SnP3UufEFDeW4bdHgmP
cWVLuBld8zXA7uT6mISTBv7riTqMoFvy3mYYhSq6Jb50wiyXmjHfuata5vxbibYV
gruso50rgI4hPgvWFwd44cetGbam6LMuG5m2xZqMmp2T9+i+YKmFR+wYF0KOhtDi
JQnvehnkZqrKy593iIYkGPN0grkChVdIDJFkuEDSti3vFAb/1SO1MfqfCHrkTkAV
2rfkg4YwHIoUTstTGT1ITX2Yio3DbaJ7wz/+TU0eSWSOoUGOm8w30qCmX8s9OJvl
RFzZ0Ne+qKI9K0UjF7vXPQD/0kq1VI5xXkLUiNAbxiPhTlWqpQvzSWa5ME5HD8z/
c8oCEOMtnjw53Fw+piHUSZDZlaepnfvhZaiH8MW7ly0as4VPT5J34Uxib6DZzsdd
oS871oZXwBiQxXOvHLF0CyY7btRjdjLDsxp8uUF7PPZsdc8EotyzO5c7eNiMfoBK
2up+Xtz1jFQQkXuVH8pSqI4NunAnXFyaAx3nC0dooJp5jsoi6+cOrKBJibtT05by
E74piPR5XkkfOb/0qTn3Px9WfuH5SXy4Pf5Si8TaZzMtsphiZ40har6JkmpHlvrz
6vQ7MVJj9aHghCK7ZV4PpuxsJvUhJk8pzs3M9gRvWTOqGYgBTcqLj4allHgT69WS
QcMXii7NUGIBEKYFo50z11tRVQF6OwejvEPyvbQl+8GZ6bjC8tLx6NALWfiC20Kv
26QVXfm+iVw6IKqY4VoejcU96lqH69BuA3VEKIynR97K6oV2yQHwCmgLVQJxsFua
LdMBncg+Nl2t/rcmcW+FKIb1XNm5W0UxGuOsDcj3fqRVkA6GRkk1ibch3MFos6OY
8kqK7VECCfRimvt5vJNQKhCBV8WedIHSXWg0Lp0Ja6fVpN0fztEhnU/journEoUI
4d0Udj3BISz5qe+zx7VTViV7AUoXqa92oMoqTte4eGibDiJbUx31hg65JIFUybOG
oJu+Y0u92yDa0cxwkh5RrgTqxGTSGDnOTfS/W9KT880/0DUa3Fye/FWdTGQCQgI4
SksV2eZjG1wIuzRkl449QNhLDE4ZCWT1GYltEbNHFKl8y531mpCbVVOo4tnXaJ9p
RcpCTQDVRt1H/YkvHEgcPiugzTeYlrTibrf+KiPO8UL5tDhapl6tDVgO7FpRFh9D
IIZPa+/8Xqvzp3bg81DnpXAHOB0cHBCyanwM+ydwq3m61m6jID0ZhE2c0thS66iR
036n6m4od8RLidxfXTKVw2jUjA3OoDrqzjKXhbOSxl5zNaHEHybSpK6HWNa4eptQ
Ue4BSthMnP1xXCMFjxOjqtsoxWQu2dALpPlUAP89w0IADtkJYTIK/22V5DikL4il
Cpi6VCCbGpJwkOB3w3luttXf+SXHppZ5GTOwnwt1uZEcWt8Mlx6ZyQ3ktB+c8X8n
VWlqsb81HEZl8pMt7UmZOYZj2wVT7HAw262Y3tEOStk4UjWIjBENldPJv41rAzpE
5uorSoZCR8lSCaO16zm2BxbCCl3TutnOUCLFjUQ3bgrIH1dWUsGZc4+n1dLbhIub
4EN9iCeno6YG0l8X+vnflJN13HUClkPB4ZbV3G5A6UCgVguBixvyqRJlEG679+/i
45PTz8xCbey6ZL+DQV4C415cj2KXD2VRdDdRH6/9X0QgukPFrPAz05ww28mtVLNB
p7UYzmT5o0JgxN8lQenDKYb+vCy8wvbYG/kxkDTrmuawhYqkPIIivVBldfcaSnXs
/9ws5fmPLj0Q/NiE8nT1ej1SL7YJ7I8J249JjT4RkSB7r/Jl+JhLVYWNukT7oQBD
9tyQuKYn+Te1QGykbXbaqRlWquTJb9UHvltPc+GdRN3U/bQQ6csA+vlGQ9Kbp1+r
otCswRA0Pt6MTjAeIN6v/YBi6kDG7ubvHs9g7j4Zz9Woa/x4ZkxG2zHoPAb+c/T2
Ys3j//1YlxbVAl2gAe6kYZtm5Ce60OncpCuGGftmW5+OqOVxH8wE4baTU+6ErFB1
IKKf+Xx8yDmH72flXHjhxz3yCbhW5nqo4l7R3VRlhxj4/qS8EG+gGJn4TqYWbmkW
TkfG7wxRVz9VUDjGPTQytc4hrWj/M53CupPAWHjT2k5rvYXGSpXpd26OEm0DrXev
xhrQ6wW5THQ/13ckrjEtsSY5/v9XbRP7s5TAy2ewZ0l8JAU7t05RPevjKbQSnmxG
ZChZzC5Mkq+2tWb9Bw1+lPyWU+4BRC72OwM+Ospljm2q6V9WrZta3vgdSb+oAz39
zdotOHd47NWtsULs6iyG7BhrM/K9slYOUDgBjWqHmPZD9kmOKMim9OCsujfvkiGw
uVCS7x/M7sOa69dz4Siru8fNZQOy/Z+h0PNe1aoUvOC/Bt4d94fXJNV9jIxhUa7J
j1g2MQLfZn5diCVynIBCfWRu9lkSlmmn4ThPK8YMZWaD4/87Y2JflWPlzyhYRvhV
8qr78L4c7rdq1T2UqumcUBUpKqA0lH1k3FZDi7q+1CdFXjOGebPv9cgP09dBlN0e
FVOUUFBoYD6iYpCh2CqQ2wal8S01X/0Kr16NLA6vctVEWt4RSs6BNNwPs/2O7XJe
AkZaVfF0ovk53S9vnKU6DjcI2Vu4D0x2PBkGbq/HMrnoHuZErLecKj4/tFAQzVTi
fyf09eDTxbVeWDvcYnlm2AF6IuulDeIf7GaRhWwea5ERySLKPYUlO5AdrHgWmZSw
IWXqjd4ztryUSOew86qtlMrvukPPceMbihW7AFnaG1W5wj3GE7s4kvZF1X2ZDdEj
lt5Xi/Ffbb3mnKnOX9eMRLwYYWuPUe9mOppoWaigepsvsv5SCbxv95JTJd3skl3/
VRHjiL1KQyxTf8QhArQw6SbpAaL66rc4LJ6m5rx29SjrIK14hijXdaTyVH2W+CJz
G9ko/YYD5d/5tmJukFyCp/N2ADvEPLgtR4yvz+92LIQ/K850/6F+XkgDk7CDwyGn
wvxnrjBmz+t3DN2pXXHvXwaUTQNaEmUgo/US73PhuUAzj0TEwcBLIxJi/GZeBsge
8bFPfg0OnMXEO0TZeFpr7Z0qLZyld6/5dKu+aPpqAloa1bBsbpDAcuXTauHChlzv
C1dG3QHt+ZLyiJ7NplnREFBeA37muMZPBe3MbGSGLfk0rNjqx00rncczwLZhDvTz
uer/vwpXd+XOlByCfSybrxTjFls3wbwEh/9ySYH9fXTkYrKuJf4iU25ZpE5zSlNN
o8/U1ga3zz+CR7PEv0JgA/+Bw7BogjixSe3+raakYjiADGRApJ+owN3z/ySte4JX
ChCv8vqeD3SWjX/xEMq78rc7/UlXqNcd8AJLkIgqkTWGQzOEtI4zEGaETuolaWje
NTqogZdhjmThxRd7JL1xG6jeBtRlr8MsiVRvOMhm8lo5RHwrhJTo34WdpVBzDOy/
hc4sGroZnb6mO+eJgCQvdGC9XRwvN92FUujhfSWSuiomL+hgYitvREIxA0fN7Z1C
4gkWm+3adTYxmb7rJBTt9QJ6X+tE15lw4a29COiwKPU7OjapNI3EpvdCrQR3yOtS
t/83AFnYmikCJEW+vI8xBOP5ueh8FLOQWPbHQnQBPFvfLgUB8+rqgv7HntPhaAzX
Qr/+ga7BSOjNSB2p6MKOaXQPK3xF2a5NrVQlGEhfqBDyv0ir1Xpd8y/OR7CQdQGE
AZ6rNx93YpqpPDEArLq1dTT+sByCiqme8omy4nxDbGG54/T74phSqL0Sg/TIN9BI
+qAzZjjLSOHg460CD8xcMdtqZKClL941CJXmf6Oi2swgUj+9wCWAM9thhupm3z2Q
r30ML0xxQ1Gu1QFAFYHoDU5tlGWc1tc6xO2EWEsXtg2N21tqMO+7uuOPmmxN2iah
MhgC1kavR8ZUiCVX5skN4qXjIQPnSP1W5C46ofQM1MqPGoVSmLb4NMtng0tMuHk5
45t29kh0XKH+Jz5AAZBcX5rGhhOaDdDbUw4+pIwDnDE8ReBXnL/jPM78ZGU/9csI
ZHjmBL6kq3+qC9Lm/AUv6rvCvqRW4cWIIu4zIlkJPiTEBemiMp7gyqSHw5HKQfJ4
vjYiJDj5RkBoODQl0WvxM/8L2pB7hZLwqvUa20kTIyiqhjs5T4KVUXW2eBG82Czt
zZ/p3wreghMcT58BQ/gQmFhGnLIn78C0h9Ex1VzIWHNM6ObClI1qhZzAN5lKbMam
uQ0ijkWo6FfndyzMywHcQXuK/bLOrajBbg6me78c0XnDNWPieqHRHsoKpI97CVtZ
s0+x3pszYoWd70aOkzrfB0XO3ZTRyKglexhHa/c6styApEE5APHPRpj3hiK2NTHp
47/95nQZXrk7v7fNtGIbhPJnJ5ZVDiro65nzMmnbtec4vME+KR5yIwECgFiUhFCU
vPu86uYbDgFjltXVnPqfTOikiWy8xyBeQT7SIguVCYpiyf5wxgqYQ0D6TrnBbnKN
cnT1gR0BcXnAIp3AjknlEi1WmrwYasntobPIdE0QDztOD4tepwtCNMSUDY93gzeu
ltxQW3ke/8/RWe7tyOhrj7K5irnO6eQVtx7NLf/euwygF6SfHZH5JlZqLh2bvniK
RlIXT6nJ60t2xOVHP/UQApQ8fDBS45BkN6CKTPHIMoYE9gFDK6SLRDfEDcZtz825
DdE8Jg4jImJmp29otU/fI5urMnFsP7zoWIBmt19bVoL94FJ/pybq1jIrkQhgth+Q
tVBZ/lIcAavyNSVSUqkf1veraIDWc9RMPQKa3ZnRayK3DPt18G1hNtDLxWDUdDDB
oQ6v97za/1mooRfaygr7qhlng4dKG1InI+xkZm/Bfdaj30vXE5b+E1UrHcRtHbw9
vRzmQ0hQ90fpfWkkDKF85W9DzrYKr0CF0zK0TM0AYHWT5+37sJIEe579QxUyQNYl
GwdCHvrGlblYEeAHAXgAw61ee2q6AzTpTMVidN73FfuvoLb0uB631FhEWDzEpyzM
0CFV3+vLB+nVC6PKwZJ4mg1aRiJXjuAqRObzyER2PlDrRAQleuYVl+opQPD7VCxx
qa4My6ZwvuKChwMRFnBnEhI+fuKyGj0gLgHbodSftbhfy8iRzYUF3s9u/UUeStNI
kj2AlEsqRHLAIF5FgIB84zrq2iS4rfJvzGx79wnL6SmmgxKnKwOfC4SIImgtlN5j
ti2Hl52YLDC+ZWS+TfxxwoeyKGb/eXC+8zMGF/jaWvigpNWJ88cvOlTI1CUZaxm8
I9MqffVJDCcwBVVQfdptUuYMKy3ll4sPcQA4KLgzQWYd+DAdXMnuqcsvJoncAYnS
i9FVpF7Aanakv3DCytq9LbUmmz51faVyC2+UAwghC4MKDiTLGw/54EawUheidmW9
+gxGle4Ik9fLqS8dH84NWbJ70zxF+fcTVbvvEDSg+Pb8xQu4xSbxkOX0nRki0x4j
JqB3sjSsxkiJv0/FSIp8xKsxSEsGgbid/YJT4zP0jdpWOxIiWFjH8pg6aj5zUdxq
I6K8mC2kPc7+8noN5jYR0QjIdtFbtdVsLwzkFyeptzF5wwdteYMcidvoHPGPNriy
xE1ArCXgHczah8KJp9UfS8SJxnxBQTvbQqztZ1rMEOcsjMRg+v6Vkb7/fHHs0UbM
WyxPI94rnq/INLsBxAC1/HukFWeKgTTlTHl0HjDA46dDe0QwRdRVLAZsuNC4Iftb
wlJn3bEO4SzqWmmdx5U4h/TQ8zgOUoIwfwZfRZvhqq6eVGlzOCBXsjLnPKkUarA/
MduOI1FRUW9Nqyi43yXWK1XecTdM6KZcCMDAfsstQpN3Mmg1oUi7kW1ArWKreWEQ
ytbknaFao+ojzcp/EjtGmyWZ3CNpJ9qpMKTHjIhxWN1cNx16uC2bUAZURA936ApP
1Bbxygv4C1XPS1giAHcK5Q1UGU6VVv6CtpTKUEULFuNKfFRBGR1VGdIEqmocei/4
LSitVhFUlPe7G+nqg8Qa3hrC2zkJdtFWoNQX2TSBEdf60+S8FzBDtyGPVx56IpNT
3UfgtoneZj29P/2hkH0BGVemRqMQIW4UaXYpaQlISrFMHjoKGjFBmh+aPS1GUpXn
v75NM8U98ZXAAQzgFlBJCv6zZav0xI8HG+2YtOxlxKFGLtjveD52suhevE8POHo4
STnuNBFvApkUEf5+6oZ7bdd6qgBJQOgx1NiOrn1iTahG/IkFghSkT9+5wj3IjzUk
U8K7sMZVisyle8UVJO/uzSf8UnVTKVZINtQn7BCfxj6NuEMvDA80LuIKFy5ygTUF
Q+2w33p464+FLCj4kKZ+humyIwrOKKUdrb1Fzt+Ko0eg0NyQOAWlvdx7DzlLBqY0
BvLORtVifCFS5rhEcZHNyiJjySizmUkhb0jNiPYvwP8psv23Xyz9jh6eBLxGkf2O
L+aNqaAT15p1Ar+TGhDn0jwuV6Z1RfOa7MThsKTvXVq4U4ci9LGJt+9IhXvhv4BU
Hf2VDc1sSSM+eUdxRPCutPEd1hVeqwPfd04jR0foY60WQH0JUUvaWw/5zqS9LvFG
8lPOw3pykmp7NZ1nxVsmViknmHJliCWkCRU1YTrehSDPcG0Ac8pNdXRM2ZcTnVr1
wJpC6uXv2SHzluE8yJXKlOzQLhy/M8Ef+shNoqVt/GY7AR1H2qytc0fyvmugAm9W
Ia3E9pYPu0bDePjBgsT9pRToBdK4ATYX9EiWmg4kF+EGrz7giaHozE7EqWGGVafe
0X5JHMbgDe4A4mlvH8I7P2n9SYnw8oCPOdIaqMzzLGAgVKs81kMUw5d2Yc7kNP7f
cikhz7em/C8dTHirkLySbrHUfy7C6VbqMcSvT7uh8XdNSr7qqT8TkTt5XPnL2C+5
5gbjt34wPTbhajCjDrBYloRfjdp8Par/Yfo06dLPQuNlQzj+MUgAHAdSw4byoa1t
xjRSIXTW19MxFArlwiIHwzF8p0fukkrft81K6nJ6dlMTPWgzHr5cSGaZmeSZwZCg
Q2vlkMxHutCzUFTRSGNln2Ivf08Y2r4+Hltkcq47p/oSP5Z1xT11BR0lWNyK3+eR
/SQu5KsBGP9ie8wNHEqeW/CVHNYrXWyRUbxnUuPK6lTr2wm6wPdRSOFoDAInZWG+
QrRnBuX4zkCGB0w9Xa+KA++QoL50mVMf+CRZK42KGWf87LcjuKCHxksmnzmy6UDo
+8ld0ma1MhvI6uuUVQhz2dFobRnOSQRmiVfzwJ3TpAS/L4TgIytEYGmGaZvAWNvW
KpRFAgmF8C0gXmC0W6UWAa1E16atA7hWQpHVtC8TMe2xJ1gJeWSWXnhIlp2d70px
x0MEyvCg+uDSVKaE37VlZ0SyUSJM7FXh/GhfF6CwLuNoa9TGCn9Gc228MQjA+I+F
S9i9czdF9w9mOD2X9dJM9zhlggM20M+PoKKEdl5mGsSqkIWdJ/yHqJpbE36APysw
/0hk1CVdeoXdypBdAxLtJct+AcFR4iw8lhcPu9v0O2+jUUu5E7qoqKPFW6pVlEiv
LR+OgtNiGC/jZJKRB7BPkRtQb75XXUNOWZrtezP4LVkuRgoNZtay4Thrr+yQgG7v
jHWsivmPFNbHc0+OBm9sFJa70kZTm4xP08xX8CELhG/9RnvmA3rg7X4TJAjrX6NW
4bxidIyKjhfXdLBz59aEgTlvAPTzyz7O69A4tDLVCui652lcm9EQuFmU9t0LRIZg
BHdLUmO5O1gMkVT59iXr5dmeFVTtbPvIxHTdM62pkaGX76G2uuAL8ra8XShOsunl
jTBtRuePBYMZdoET6gS5cD4kYMM+Q8QRGJ2kLErfKEo4DtREFRmSGhDQaUpqgNIO
rzX3gNuK07low7bUbyCaCWcossbjykhNn1eCw5bAlNaXjBI0MOeKu2ZHQ7X6C7m1
N/sNHzFvGIGtHIMYnyD8kcKzy2g8o7XnCbjsU9gwTpI2ZrbvjanwV0dh3d5lwcwW
d8Tf3zjV7M+xv9iehaVZzs31oNTcDroQ3LeGQm3Rr6BUYVewfyPdKJ/fMRjOLWCv
zP7wrTK41kvg216SHWSVNv6poMTQz/LBeC56eDNryEq7GdoK2dGiibsOs5hM0iRx
DOUxuaIzpdh5RS2DbmktxGPB8ADocn2qOE46foiHLFKh1j+obANCumnHO9BHBY0f
EjcjVYZY/ApJ6PROAOhuK+6xExm3ZQ2B7LvE7/l3xGUli7/SQmbvTlPUCgW6OR5R
pSJjlm9co0h7KkD/rQEVMu0smwyBJdADZv4ttQz0JsjNY+Tgwn6Ntw6063Z7iatk
JEvM8gBeExXawWiAC85aoWUaN3s3yAeJI9H9AfoUsbG0G+Q/reG7kT22PTH3n0g6
ZI91fmu//iWxeiojPfLpNmjikiLi92S24JemuDf3rmgSmcT7lqfA6GYGuM9vj/H8
zZ12WcUkxADFvPvjVfE9CYu6SkLjbj4Slh8EzR35KBvj4FhZozWB8z65PdxwmuOk
q7M/9Qx4jCTzsH0O7OityjU5znfa9KIdGRiOZmvt1dDUBoZZw9wEPSD9uTwLPB5e
xH1DBugat6jQKmPFkqI0ATzTj+Gg56vCddL83/jxyR6rCJ3EFMgF2ldaCQ6lzC9V
xbBkI3mpDC+wORRveh12y2Gkd5wl2wuV4jzhWiksVB+MXuyZ5ShpH0lYGxAV4aTG
9TEJc1ftVcZOeVszxdyZElp098WW/JkPZkkzqsWLGxOERigyhEHjZ+E/zGi9OZew
OUP0zY/aL6swf5WMFi6TMGBvUNZIMbF5J3Rq3LQkXdrGfBe9ur9dewdNh/4S3BSX
JXLi1qV8FJqFSUxhUMxHE1cCAZq6v7BxGs738J0uwIMoWJhrl2cSuLfyk2pNcnlc
tFu2AEmUHFsTw4rEmOUyH9d9nFBF5rLHDfE9l9CnfKjHGsnmzt0YEBLb6WUarGiS
oiFrHiLxtwjcHEf7EMl45ZC1cbHEhCnyS1LmkAU0TnIkK8ojoOv7HpsI1vaXmtb+
EFA4VTl3hvE6XuLsjq0ztA6ryKpCqcsByOxJ1PiYpBeebZyV5cK6c//9YWcH/BAf
Y4hEHg+UDpSLfbcqLu66dh78Ym53kTLCugAgVzIUxTaZBhGLaKWdqbq7eiqIL9XD
nNCmkLC1L5yphaxeFfgnCnAtErjEN9K8kmtQS9wCdqA5SCsAua8AqbL2bmzhtmAp
/2gsW999cPynoZzDEQGaArO08yyHq+82CYtBPeovkzEqHZ/jFM3SC+rFD7T9haue
H8ShUb/mPsVbMY6tgesXRPMt62BBEzlRqTB/D5ERZGX292YdEuMUWyt5zQ90VsUU
EcX+76ee0NXCyfDfBCrDaCYeKwXB4wwOvfcnVAQQfpHA+psOps0jKl5eP21hxKs1
hWCDIPLCgVW5FXU4LlLSWRgy4k8XDDfPEwSuXfw4zFj/fXxWvAhb/0fUGyHW1er/
najg17K6LSprLNALMLWMVWxxRgn9cBYWFEiG15gxTi6eSbvWjW+Whdikrt+ekiZZ
hK6uYa5BZZGxsWYP9CoKEGdNFSRUzMJsD+VF95pmKN/AQzlLEkBG+pF1uKjC9Xa8
WLuM1gkVRBHYR/9vyCeCAH+85+pMWttrm53rsKTnDGzo0qpIEurvqqsRwWh3eG6y
BYz7nddzQdOJJBHj1x0Rik6DarPgjfhL76JzQNGo/vfqAKg6UsKGMl1LJSuGSyl9
5KK8mq+XExR7RwcDP40VLLVy6Q3oppMeF+uyI9/+VidCu7dNWq05qulCzOmzowsl
kWTPawwHl/yAl//fgQdQYQx4emvcm5L6XpE+MPH1QMOZWV/dEaoxmwKq0I6ibSJy
9YxVlqP4I6nN9uxEWYESOCJURfn+/B6FB2J11s80HxMcb86mfjvex0XoQb/toffB
m5cH6qJ84WEr0/HU9wycYKseTdy2q8+DiWOLofTqVa8Mq97B9h5L1LJAvmrLfdUh
m1e3TsxKq7D9Cqbqi+FHTXEU+fnVQh1IJ3JgJD92sTyzN7vlyyY5hMLaejHhofbe
+ltBY5IRDtI1/i6nxc+yaeu/R1ZVv7vlnVm2RU1QUqohxGx13WbTVisfU1wuS6ZQ
ZpB9BHXU+cIgbH8wkC8MuX4XGHt4bQB6wVumUyzld36ImizOQnf18JFZH5vPwThS
242NkIFoo6bGfEdHsD/NqiY9KnCyHpJz/KBT3WnVQF+iJpxmJ4GGn+p86LlYGOM8
JC4V8P0V7673qJ4Vk9GZVBWKnqH5zKW07ZqQPg2j5O3V4zh7PcKpGIK2831jre39
wfROybnXhrjLEyrEUsEfTir/B2+YOdc8J2IM9uv/67TGfEAaJD0OaZweu/j5oF4V
dsT/FnqYMJE7yybCD/OeOLI8ofrJ1C7tAiibSRb58mGgEjkk8/6h6sUl5XKCwSWl
Yn4rVpIBTAI5032d+RVkYvrm/vdJCtyGj/zRB2EVc9keP34MG6onTsmQJXGKkbCB
ENmTBDY7/lr5Thy5Tx5a6+RnV4/aTPMtWB0MUiEJ6emHwL2saFk0ttiHDHgqvCvw
b1lXdjHxsaq0QfxOh4sw5u4Kss5IGvRWT5IIuHiqjzn6qa+sG233LRfs3+igE6TT
7qvsr3dafbkJJ98K50y1+y51CX1rtLV6lRopSwdmsabRp/gCXq3iMsNQXbS/t4fV
WY6n2ROP8ZPA1iY4H3Nmqmndbgw0rQmZBRQIgUS8CKIuAcbYHxjT+hxfwUalLD9N
1VG4cyaFufc8lvH/+8HJSgQnlk+PprwY5Tqh/cRc0Vv3KJN6xtjy5BGGcsQS848D
0mCmXrlmYEIsE0ne8TUajm/wonuvOEh5bWTJaqZkkxc1hR4VlUzKSlLMjjcg0HpU
oP5SVpRgY6zWme7qpJ4Nx49p1XdglDnY5A9RS17boiyz3YABHR4Ny0gxsZU9WzKC
8Ps3AvOqNyWpI32d6x/t8BCGnV5i97mfwTetsPWBHSE+mi4ql0tttyoi2KKQD2ST
CdvOgNSj0k/nfBaMY7oKs0FcoAvg/S2o4NcI8HhcVjin2KsxNdi07CjgZSxHZW3y
JTQSXilHdhfsc9h7BW3CeYEOF97Q459vjnyYNn7ovIqItr+Qizc4AEO60xPb1I5P
OzNDMAJBFtcNZAkSBF4L+MsXvvPJ6Jf6frVOpHBk3Sjrpln5P+eUFL5ZIyDL/a8B
ldJDzydCB8rBlVEkqYdw3/NoBCiC8XT9d/sE5o1DjTh+MdFlE1Me8FkIXScuUO2D
B3VWS5a6eiU50PtAhJ0UyDQGPWrwhRwK/6v4Nkf4mRL0ZXSrbn87C68+OCxfVsnJ
pwwy0RerAWgL5pPwex9ofm06ofSsFP/afHidrGJD9u3xrnbWO/Cs+qoUdmMo9L3s
rSomwpZeAqlE/LeTksLwHKdVn+aa95fwq2CVwigEHLm7BNNvnKHmE1Nzm25BgF1t
5bqXEv6DdIazb5rejGm7xsjhgd1pBtLnZCPa248ThCgF5mlH9GJUc2ts63+/JDci
v0gbdpfAHWi8EEoaZpdf4iMDDwcmoRJCuENhbxb3tYN08g6x/JIU6omDWURv59eD
81r7uAMPG//wQdQ8Bo+zRWnc8ftWO+GB6sqI/JqNjRXbIUp7fvqgmKQz2z1U6/yb
uBBB4OaLv1gg9pTRwPOaKfAPxuVdzKVevXoNeci04fLrmTMgnxsE8bqnb9lYHxZ6
SeT7szmWqti+qGZINlK5DZI0pNK8u74xq59Kb8otM1Vq0o4LfwdGibHODunCRwtM
W4k/HX6T5D7GjYC7UyIKdXItL1optUe6TvXmwr4OAXGQY/TgRXhJJWDAHUlS7Cwz
Lsd/j5ZfK4MDebNG/S9asvnBbUUMVum5iW1Y2SsO+W2eO1okLjUJPP6dy+GsWzE6
ZGOz36Y5Sf/vmgsMq/qiyx3lK12BDrYYC7DtjwaTGLIPuLm9toK/NkhII9U0clxE
ohoaziHJ2S0oKDHOMD9key3VC6sCqLGMSDtQpL9WUpCBWb5WnJhqs25V0GHSPbzX
CqYRXL4eFZ9V/FG9miRBoqgxS3chZ2U6UH4iU/nLREBne/Xyd88jBt7D7otO23rs
vs69QlJuPhBGKNAH0B9uoMbcKySEHp/fWUVSQLsCIhlxWBhQUbWOOqD90hJUD4xl
+efY5BkZWSCuWT113w1J653lpqDyICrcrXoZbsvnPcKqgR9oXtnMtJpb/kquN7eD
M2yMWBCKmr4zhuKTErD0tVhWTCht86r/J31BDexlQbo3SymUgYXP+OLQkQmaPtfn
noHNEWbbpGBPL7K3jYQR8EFdRZI2OlJIAnKt2PW4N5i5zaaals7eWKOKMFNWd113
PqEzDxHPnuGlDfaIC4budcW88vQOGG+8q+B9RhlKAIyMQADdyPDJVGFfSXZJpD4a
0vZp3g/SySHVWNe+h5kzzK66xt5RwMnlC7RGNtuntWs6DS8DZKK4O5/ZxErAVM/W
BMMN7fx8u0zm4QSsY/pTpDkeo/OZ+d6xT01z/5rNa8iQScGfQ+JY9bvDB/CsbDG/
JHaoLBtYQLNK4/Vk/L+7mG7W0sWET+EKpMNN/6YrwFTiTHGUhyfpz7Ot3RGFk9Sw
uz/1pFNPClyiVyw5kLn8jVf1n2Vp0NDXIW7755MMVoJtxeU9E2dsXA2qg1UUyY9L
83xWQk6GC2j0hL3326A1zg8nv4ZnQBlJgCK+tSImJ0EIMjBGh2CN/hme1ftyzDcI
OIKwSQlr+WJGWil7bRX8lusrpNU4CujUOWzbNzFXkqJCGZqISpTpFekx1T6t7lP5
dbBd6zswRipoGenV/un038cHodh3Q2t4z6AKl5kFCQChtoyKkorH4ds0C0kg6yyV
EU4GYce30S9PoNYhysOr67OtszGnuRUVx6nHiJzH+bKEQbR8CEW0v15iOB514VL4
M266R8X3YAeSwkdZCT1v9yYC4BMxRBWegXaJYjuMb4dE3c6pI5fWCoNp++Ex5wIa
5y7gAi+p9q3ctZkGz3/7L1Xzc4HFYVurG8VgiC3mmOh4XVh7zuH990+Fx92lnKti
CORofwC74u1CywXDYQHARVqFVa8wEorE99LXoPOvh4fpbHB02+Rvn3NKURaRk8mj
abvkC1oIwwH336LRGeFXAoHi98lrTusKOzIM41VMsNJ1552gbolRc+RKSdijR6og
kV4YGd9+hYi/ClA7vk2xinJu1U7STMEyyApy2GhSe2UswT8qWeb6kplaUqTliE/1
Q/iXzwt0iTpw7/kFRsWGkRRajC1arlLsno7FSCePdMU+C2NphvIYX0VcnDcRdW1e
8SPREA5Qrn2QQSePhyKXLARkuu/ul/a03sBk9YCjOVmIIZnZs+VumExKzivCB/L8
kJFoUMIFHn04+lSdFCkZOLauieGN6LssBeODKIdWNKpKSH4dT+1GnQt5q7UtaNWW
/fW6Hicpr56uJYQ2RHi+WIP6xNR/+gl93lC2H6fkDO5sLCgYI//5f6EcZ4hx2jBI
qFo0IP49pxew6thHT/Iimjz0iCj0eepH9td6Hikb/Wwo06UzPzu2leCqTOdgLY/W
YuE0YM52O156LiX6DWDQWqefZkzxUv90Nf+jJaZG4CdGLk4GQ9yMRG1TV0wSgVZ1
zxJaFiX2IMzT/jtBfpWamRDr5FiOo7BaIm8kHBO2qNJRBhxkRrJ5yv5FodCP3x/J
/falIe11fnoP6IOxo0q/yqnQUFz/BVJdPzV1UICHhFutg3ftV65DT3c0phEmqZ7L
mgahW0AQiIUtu/Wl+3+Zm73GRfOaMZQqZI67Cwg/POAyU5tmxhFIuPnI8eB/HXo0
c6d6baGyt64Ad+Z5bXGunp/QcCAN8q/09aV/NUrHUOvRw4fVsf20GEDgndVqq3KW
e0GMtQvc+2Kw3G5GvwH1oRfZvpulYfqDg0nMUiuZ0v+BAQGRrMLtjZcSL68aQSyH
5RMW2wkBXC28W0oxLb3hQ0Wjja/woE7+FsbpvxHpRT3502ZOtEpC5uVKSpuvAGxt
noaxR05F/KAWpt3PzM/BKme/TPrW+8fX6rlYwroe+LU1tjATnde5fH8+ejiCmrSl
oIJRVT1ldYRrQE/GI4OWP3Y2FRaqCwZaiJZvN35kXDxdvprwUUkf1u3ADOuMP62a
bVk47LduwmJcl+pYG/BUExuqHdE9B96im8e0gkZ1jq0IT38nvTLBDjwYwkA3wFIn
2gsyBfcYFCLVIXP674SF/0k7AO+UxG0W3cCxhPRoPtaHTiKkuu0z870Hi61kpZVf
iFE+VY5smESFrNj1WBgIBhUvaS9nz8rSkNVU+Gvq3rRmWXt6mGv46bClEpjfoO9G
FD06UYqfyJFcuYIsYRWITWKqkGEMtB+yk5gcoETxunLAqAzrul6NdVgd5KH78hWd
tCjNTWefl16rarZnqi57JtLgqZ+1tZrczx80F10duZ540DhdS7FJ7+J+Op43J0WB
+kc8YyOqx4dvTS0HuaKIuNSBM7YvgjvJz1ihlbJDR643eO9TKIc6YPPF+cH+Cu/g
n0yf6E3LUz4x/JB0vVE8adP6fZzuNsJJcEcbsMQIMeuh744LcF/TVj579OyOopxb
Xsw8tkI3koGcm8bZ2oULoqba5TM2k+AyS/ra5xu4mHpCLRikxLIDKORpGQzC3Wrf
Wra41mHhe4XnkMgYCzSY/Eb/EGcGZPqKqy3UNmadfz+1RenKmfGbTkd1tSmLiOQL
ZCeILQVcpmirKl9kZij8pNH+xsemxByUleJPcUoFcday8fl3sD60C4TwsW9hTlPQ
wbEjufnZLW4WrsGfIUjO8w3UxDTIPAcH9orezxjrlwvzSTsNN8AQ8LkyWjYbIK4e
Nps5H25Zzrlp9st3ns54qsvX4JoYWiuaVQtlD9WFDnjopcu2+g6H0G+AMw22kVOO
klguakhw5z928dsYwMWEF8hei/Zkl8MLzcKliqcg+ZqxbiVxgbq8rgBfdpcmwb0h
wfGH8EHfRlFxnP8DUKf6ClWx/nyxI/aXVNWm4d0Oc178i/vM40U0A1APGvLl1xJI
P8W0LOqvV7wnZnKCSuPwj1Vf/nw8sORjrqFBtyVqF1v/y5qjMnqUxbdxPrU8Pp19
LmkXDdzolxOjK7hPYPk5hLr7gLXoDr0apGPrq8/mn4H7TzQSABiNHcxgmfbd+cew
20SspYCBZAswffbi69B2viRZuyoOPPkqfgQGAdrGwnygLlcPledX6ndWbhDWtnbh
zLzH/yr40UCrt+H3p39XoeYTsBgncMIRejeKdP6yFvGtmgSCIhBF4q74V2JF9H+t
L8rKlDo4G34yunVgfhE6DV4CiyYgNo8bIP912c+EdSj0U2HYRQdW4oGQSs7inf6z
yHkQ3m90kJjidgFV2rZH/iiDmpv1qJ8C8uRTOunK0F1oe3VjVEhBT7S8meoRusxH
reKnGml9Y11yg6lvZX5MXgjyGrS8gS/3gsJkzWrUm64/NvQjluYnfyYifVKPFJHO
/LRCTO8amKw1bbtrCkTC154T6VngT+d8xexL3CwCEMyIg8fUJgbELVXc9wEptwL/
CXXfyN+X7Rj2FhrDNdKpORPIrd51pdzoZVpTt40Dy5ANoCy6QwYrNK5POsTKe6ay
VD6wQCHh3k+WRzyWMrD0CQAopN0SdFNpfI9JXM8vcLpLncg3xEB0Qg2x2W+13JiD
Iz+9zMtTXedaUBaiuBkKkYaPVjZPm2MTNMhRf+IglOI9i3+5Ssu2AoHbMFgDHDYZ
2kXOT/3OsbgepIVTL1uMDWsl4kyW252O2m257euXkoXvwqSHGk9qTZ6n+8kier7T
tuk+arGb/jRn1GCmDLGs/vts6X0n9yqiJmZZUIdISwIDkpSUe+0LtHcKB6zBxyWW
lbOSorD79q2nYRPvTg2Qc/mOtsjWMwRc73Qd+unE3HG9fPCU5awSfKkZiaVeGPFc
4bFos0folkgIU/Y4yQgBx1m0LOOkb7/JClpWMTdmX/UboIyv04CQLzZ/H7z1kwsE
Qt3J5Kvdhw/fXr78fHKvIqTvWOkn3SNfI5+tqvWu42S/+fbco8uUB2g+lqOgmG49
MN6yXuvsxOaeSffPOB+6gda9LquEEetMxpBh5U6rCKxzxJ6nFuyOp3qvIiDiTjOH
G2h//B9XUpHM/HnX+7IFy1jIWtYvxpJtPMQAltsvYghKWNrR3epxqpyHR34bcIIa
ZI38X15C93XyCOTZP55opsS/f4ofwPKvwcE52R8GDm8Tt167hb633vP0/FwBJLG8
ZflTa5cAYRu0LULBcF9eF1T8JvYFJ/YrGNJeOfIV1r67N5OmK1dTucVwiH8wWQb9
vg8Yjn7wMyuxhsF+L9AhfXzfI5roJwxvBZv+/j88KNvYozBu5oDPO3VtTWReoRiD
UJGOU/4L7/LOxYetJkLkk/l6282cdJeBr9Wdswusk2h6678YTB4+OrEMjINHRASV
8JU3Y9eUOI4IfKHuySSAp+uBZKCoqepqKjRfzOAQlksQZpRAg61K/YeNd2OH+azq
BBZ77Z9yBOITeoY5MVYvH+euNvYvoSTvuDXKSSH3GuABiPVsjNTtGcHhxBvcpdK4
C5CSM/KCBNkjq/o+Wt/W87pMMmZbjpVcn0VUF76iXy3yK7rP51Opki8nZvaxhPqA
eA/c1Pdy8gPpcPEZH0i6pNtND2pa3w7g/E+wv7frs10+dpVJJa/FEOmTGhzsLCL1
b/yq4qbn8dSLH9TWZmu9++uuA/7k+1BTwF9p7nFrwZ47oEvEWF/mR9SUT1IoJwv5
7lTav5WWtTc9PLKsf3Jtxq+yjcAVROuamrmN7QF4W6cJp5I508Mv3JAa0FXMz4tS
zaTkPsDGYTYxEFatXGC+Jz7r5Fwtbk4L4cd+817sOUQJLdmVqUirgg0PEPPq5voJ
clzcW8Ld0u0W527H3/hLK2JkHdfjKnj1XFkf2joNLJ5pSTcONCxGGteXVd1KOnzC
mCILg2zfMB6RiQDjirxrio2h15DtZjNs1BqPT20vJVw=
//pragma protect end_data_block
//pragma protect digest_block
FKtMoMxGcVoxduJrLYZoK2r0zLE=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
gk9wLlaMzhQ+1zNHXyqJMhhzY9++fWwoyUgLfdX4Q+5IOyXCYTDJePq068dpcfrY
/ALSTDytPzNkWP7BmOzr6W1yhoHYdEli5E9yUDlD22p/10x1yY0GtDUOCjVseEUT
Gi/vQZwtEyc0coUjmiFHrWqQLVFU1qLWNv4CovROSs7qb8grjX9/PQ==
//pragma protect end_key_block
//pragma protect digest_block
DwIQwIrztIRqwXPt1n3lZEYspdw=
//pragma protect end_digest_block
//pragma protect data_block
05jlCsmN7uRHOp+T9eFa8dhf0N/nNouIgHhfxEXXTTuvShVCG/5F14/liLxipuvp
ltMPMTiE1AF9OMUiDu+0n710MyPvzWcMdJBFB8xPzjiWh48Xxaioo+xcypE7i1g7
jP9AFIvamUix18kveZKW+mFoJxIdOOPkJyTmMDiysaQuqKFD1ENk5JkR4d9F+R60
GCjGRxTRtimU8p6wmithrtLGOhm6DRPF5ul79FHZHetoXixP1nO1rC1vbnmEuxtJ
IsPF5DpLyxpmBQTxLjbp1bc60Fa5XraP7vM+Kq2cURtikXOfnmT4mXvREHVAxdXh
jU3SUGGsD1mWsMCnsFGbxMzy/ZwqRe4mQw0neBTHZCJiqEiWD0py7tA41CAbSsNI
1lKUs0d3cQyCfu4b6U7ZSxiXJ6gIzzilaGhZPaYj6f6sDfVkBCZBi4NOe7gouJB1
vgXxOvOj9O2l30T1xpDxD4APZRzob8oHsAnFVcuzR8unZvWfJGjQIOAN5dnl2rbF

//pragma protect end_data_block
//pragma protect digest_block
QE7fPOFsWYaBXsPci/BRzcd35xg=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5AYRtR/sUcM/RccqljBN4gPYTbGz8ru2dEs6Xm+DVBVz2GbDv+FIvoszzkBpbMXU
b+/k1WZVfj65SOMQO8bmdiYB8KsDqt9maooqdiFZMn1GnwM1NuhaUtKmpYwdMHPz
BRinEYpgaqVGLbMa13VH3jrdcRLksZGkqPheOj0Ve9jEtZWeNTYaBA==
//pragma protect end_key_block
//pragma protect digest_block
M6A9aGb+fBL+QIwRcPcHSYY0jdg=
//pragma protect end_digest_block
//pragma protect data_block
VlBsratDvmlZzGU+3LUuXaLOE25nd/30xIQwSIPD+Jnox4j7Mj1vC/eTD5gY/A4F
V29qFPbhM+gQkM9cDcNENvrvGWZjPLRC0qQP9uTHsu1Gan/EjfQMsufAxwnYjSQH
uH49EnSSifgHKFDSPBbtbUY7JUspTxwwkkY2gvQvVdz0ifSEmuG1rOixii0jbR3J
/J7J8rqzKqXcie+vYsAPwgLffuYx5XXXPfFFVQKI0YaCY+abiK1Fx7S/x5Sy04+T
jP8pHKKQl8Dc84JlmzS+ixOXMi1TNKpqP2gCsy1StVdmxVTYH0Zs1ps5NAbvwBwZ
G3PvoWZ3HeCwIZTiRvhPtOWgMy1FTkjjR+Qn8mr/nOKN2iPfcg1LdgvwujvpoL+T
WdQzjoqZliB1yHHsuv3YOAVkNaRB06tmcWKT4srWfj3X/dF4NOB661+/hgTv1h7l
neOsaMX0ElYFy/Ey8EQ2JKYDVaT9q4cDR//eMYMSZI4yb52QBBkbbTcY4bZTFUsE
5LFKDE098Pzf2AwXjMWHBzUE9kGUoGZo6FVY+0ad+DN6jwqiHwQyOrHTXHk/L38y
zw9/XaI7ipsMScnrGZOXD6Pvr2hGlzkugK5UMMj2cifBU8B14HOGon6sg75XkcJZ
mYKoSwgStXkR28dV9qAEiMpOpPA4mXqYTModKOymSfB4utbnxFrVqVenQvuoBwVi
WYFdQ/fXg2Bb6L7S0jC6L7sm2V16SNicA+45JZ6e3HVBUb2lbrwncmfDq7L9VXsz
EodGGq4LA/fgeXv6cjsf6PPpCgKlFCisRPjHe+kMg8yPvBFRsx+8/4yvXtvbN+v3
XHclS4f+FWo35ev8gwxW8TQV/mLDo6/F28e95vgLwXVXPTmwNETe0kFyk3y6RSWF
FtqWBFPNe1q5T07hOHCL/6kK5z27mZgvnda4GIgR/8tPLs/mdrqAq8m7pvxdzLwS
4siTy9IdZwHkU8kbND9Tkdr1Cnr2S64bWjtzoYRi+IxTt91Njn4LH2jzQFv4JaZD
HmSng9C7fJyYPu/5xyXilLJnOZMfuyHacG3S/rrO0B3YohzrgXFRuqHdapR7jkRs
he5V1qMSLIrA26+em6BQntYmygZ64buHdpTXqwJnHNds6noAT6mSK0dMjivfDtwZ
gD8YQG45nevLaROldazg8qXJrmGB06KQ+RLtC+FKJLz6e4D75NUR2AopYq5gPGtY
tKJrIJd6nzSthPXHi6FdchRDAj+bN3MZRC4eyW430u5yIs3LCsuDuhhNj88gPxlG
cry8JWk20Pi5IP9KT0TIJeG+Jda7fFmuWgD3Mg3P1u29DEl0oAx8Oh2NhDi8tKIl
KjGZQiAp7ms7Pf18meCZ9x2QELvkdzRyLnCtHirStAMdeJORD3Utac/n3kSMhqgB
ZU3i6liR8Qc/W+wbghQcH00TnxRIi1zAd5mx0oSnaDLDKAnwziJPmqMN03Mtow5y
ewtuUtiv7cFYmQfcfUnjkPa+5hyKwxI43VHCRb8pRyUYj/Kot1i74oLuho43Xpa0
nnueDabMy+OI0EygF964RApeEdY5iB5OVpq1YSccr0KuxyR8VKl54oMrMTnh0JX/
cgldBwHmGRNWQ64pu/28BM3GO9LzaF68Fh09sGxU+y6Uhbphoz9Mf1mWs3ZwXUim
zzBGqChSacUKKb7FFv5kGFu0n8c0hCUAAGbc4PabRHA4zulSlTiMBYUXeFargSvz
rG6qQzjFXFV7LtzL2Cd3dnbIDtU+Jh3Al1Yh8SxyndFOkvHkCw+xH6x1hBtt32lS
WIlbuqPn5+T82Bt2jLZBBKMf06N7Bru4ST4uhTovNcI3h6Ly+CzhNnfdSSdoMsEN
KzB7jnyrvHPs57xxLhqUoamhjdNYAnTUIOVla2FKgi4cuW3F1iQ+w055PsA1/4s0
dP8E1k74C2LBgArCo/nkbogF2Ripb5mVPBZiOuJDPJsWDRHrpv1iAJrZXdel66Ts
ZUz+zpeC8nBYC45U/J9ZMC6aQdv9WY0ZxDSWXs0gR/V28tMGNGk16+p32yzD40Cx
PPt9MG18VHEdX9DwMjW+W7//je5TLMtQDsuIvNVMi5WY9eAXUyDNMZdvWUp5hy4q
+oZfJJnJIgjQL4smk0YlwWzGRjsAUKU3/lN2MCqR+uIf/aLQ1tsi9JsO4I9a9QR5
fzRHL9nfC+UKm4PJlt4CvjYacNyg+t8i1v2nK+BvvKuP4F5ojPdoarqfJuywcP9B
mwxsgcEItPZfenkZ3Lcd1P2DzNW/o8bPPbtMrb/W5R2ZVnwlH0KKu+9r1F/FSWKU
rZk6n0eit3b2lt4lZNbrHPitmN2p2286TjezZEYW5r1g1zffwgehYn3cTXLGLlq1
cHSDE+7GYcbb0lANitED8PX5XCRqo+1zMDF1I/mIfUTpnvLmeYXW4OQUqv6EzcVy
IDGu6GSLWGhZ1pPOb03f2j/t6oQoeYtuwKVDF0Lhr4dSFUe7B1ocIEqIeB1xbC3U
uGLgM3E5k0rBWE2YPLTbQvzt9Pqe8AFOeG8W0vfwIPynN+fbgIY2jND+YvnMrbQu
QAQNUwiH+AT2B41hPji43jaTy5pMds/2oQvKAHL75wiBYKEyUAfmZxP+E+wlDa7p
TDtPuTUZqN3Pz9ondauQ6MTePnlYY+8SjZSYPa6mCrpZeJs6CBdG1L5/hPvWyo9D
gXKOnxovrGQWKORqttQXiR18D4sSJAADiv1BtMNBxYHd0SJau6z14RGbOAtSd+it
0/7F+Gjg41nflO/pmIpU0KHDVnYaGkmJSFMJaYn21lIPk6TcZ0t+wakBe9lfijcD
Tpj9HXoMwURnOWazv80Jne+gODr+fTajojM7ARYuSsU/KTda48pXGiVzT0N3gVnk
p2Dk2Sv81ax6ey4hkBZ8fXFVg8sh58cx6q6Rj7BTaJGHHlxqHaWEvlUq+YxS0rX0
qLLhpBUYfX0D5/EjxgC9hKV5Dsdifamy2stDFzb4M4gVHooAHMqU+lsZ9SmoL797
0hkGHnoRZeiq9woq7ZUl+fIm3vI9v1KyMxB5zPqq/s4xuiVSZChkUdX1mfkbTnIF
b5JT0ynBZfcYnFSBDh4pnloajypFDw6LUn3jF7BymCxJuasCURWUCrbliggSZm6M
rcsOZLoBVU7gOZGEuwO13V2VAj0dWMmfs5pT2CsW711FEqdsv/IPSLFjcJbSzurf
2uTa73wMDwhuEg5ySO3lt/xojT/8tczBQc9rlIi78HWYXHrVDR2aKJK//mSS7I3R
w8n6aQHOpyCBXFqfqN0AtKZ/8eLlcILFsSPJAUWA4qn0GTXSa3n+K3WH1kcRLrxc
Mv0NWl4etht7XDtMpYL4MqCmzPipjD+IHrhB7IyCBFG0Cn9RJaiRlcgLep5mHfwH
pLWp6JW0ZgDBhcwim71T98ZtdQKUfFI3tJuCkTymC0E2IM1j1e5iqG4BppIE7YvX
duBaR12MWZiYt32R1LYRgQacuRU5UBjCKJ70rttYbnBd40PuffFuCcPpKb7wmj7M
RNP+iOR73OGU97V18ZgBBulctzHWpMhfW4IXbtRvWNm+AS4mcaqupQyX0A5sDJoT
O+m27GMeO8vNgVcMDX6OMgPGmwd3ViaL1Ks3FSxlST/Dvqsec79gF2uQ98EsfYW6
llBmk1Whi8q296ZwtFHwbtdYNx9JpmRgkhNPfgKZWw5zwnxRePKDu37RqLZfUy0m
oJFFrHaTTlxGKzun1d1/xAgLCJpI1RSdNfjZbNhAdf/VMyohvhnBBPnQUYXXrwYD
/Tm5zHrhNtEISyb817DGhP57Eix/QH+JcgwLCB8irobJpvWSgwPWiDpU7/WEwgp9
lcGUgrmOzo7IfjVdpwN9EpH04TgEvJjXLkIsta1Vf6kRgrDt+7T324hJMfUYfgsE
sFtz5DPb2FfzmKslxwPOU+aTNKor17MSZKWlsVBuJKPJmYfEemRze34HiutFBjlS
/FMLMhoT5dKPNKGDCUK4Q+aYNDCmEB4YLW+JG/vPrVOp8pOdpUv6vSZeDm16fIFH
C4j0rzg6cmnrjQDPzqtoNLxw0NcYZ3yY6YJFckQnuOSZeWZSyZJbY/4N6HjtAca1
RcWGd2wIous/MmuuPY0tpWrlqHXYKjbBAMWOkvuYqhpkQlxqrJqxWhqzbevDdhyr
7jFujvr2k9322/YR+YNE8tCqwe08kNr5Ug0FbfBd7RXk86Xyjw2Ojf7zocz6Det8
QALpuYUDz5et6WwDU7nxXRcvc1ftTsRjNpWQkpR0DxKhOheedeSuCrNQz6cLUoIY
GKdPAMZk55Zu/i54f9pSfCh3q7hmBSFRa1MIXZ20zQJiCRwnsDDlPWBYRNskT3tr
QGFmkkf3pFQTNo7CRzVa7dokloazNAEgqS0bgg8qVn7kTJwuZEvQD76NfbDueYLk
JA7A4b8B1pandOrykh/JbeFfhyB4l03iCGgYORi/gEvevnB40vYW5mGEicBtGarN
okpFysXj1n/BAKUz03BIGgjGJcVPMFn80jeqZJc7SNUQvl3yHfv6bEEIy6ZBPasM
iXt4LIBaqoQvg/q1vPn/5+piAGmXM82vF8e0RK5+QyFsB5FfkFxKs/JKWERXoO1r
+VL44uBQZUASrHmMXe1QlGwKyLHWFZjTXSJjbIbBxoZ0HfWF8RhVn9llAptIkjlt
lZwU5lWlcCmnf4d52B+BTbwn1SFTCeY8EGngaKyFA/kX4u5QXvmURVV5za6NAt54
KA3zSONvNr19Udo2whWwNkzyk4Lj38WKQVaeTULIPTqIc6WG6r/yEJ/h+hQBg9UM
JbQzUOZJfuLipAWw/Vee4xnl7C0ZDsBlnEAylsSChmCinEdktaaNIE1EzmwdUHif
mUx60wUiez5ZhPu7TW5qjJuXukx4hLv8zOpbI0G8z8vcAfe1UXQ/Fw9ksVjN26h2
n71hJLWhhHOpZxoTebzLEeToA4HwX0inyg5iSaQ9esKt14ksP1+qJuBw02Peoqo2
CBqcjSCZ7qBp0fQ1NmU1KLjl71D2mLl3WWt6V1EaqfMOQ6Gy6y4qyreCLnG9n+91
qVFpRUnRJrSon7diV5Pc0be37GDPlw+sXuu34qldiVegZJp3lWgyuyIjbMxIb+Cz
SUf41mVEjzzyg1jhcH7o7S3wzp2OoCfc23dZGvMGgh2B3e/YAm9ucRybUu7fBOM1
3SRFvIRNQyZwCoS3uvZYYBguOmMizHH6qK6p9JrJA5Y7eyFjoAUI/1utI89Hp0Ui
+IZL/Zt9n5aPNAwSC5A4MZ8PHFXe7sZFLWjMsDDsx3RNCvFca14iluYobHfsLBC7
0C61Wky9mfowHnQUApcYsZP3336q+4IkSqoCQqmSor8kqXq4HBWKXobRe61kl63c
GQ1INxZ8f5ewk6/c5NiDwCUNY8iDZBNjpUMdkqZ52vsqTG1+vel2hkXEJWFrK1We
Yd4rhBUWlGqbI8spb2M3pheL6BEDL8uM5bTsYyZ4GY0Y6/DUR5FSeIKSd9iCCgkt
6gkfEaiE2npS0h8FJouUTKuVdF6rQoMHHYXWkpDecAtLHoR2qx1Pb/OwMCVtxB/4
YO52yKI0vhjpPzvZPSiV127RKX5Tf/LvlBzfSPpo2rlD7XDMWWTswsuylBaMdgKr
8ALnCXQqHhkr+JbVeKvafhPQvQB8bID62od4PzWsKaivU+Xke0k5z7KhwmS0dR5N
NL9txG2YyddDhi8WiShyWm7B7WxkOf8yylYnt9aBbAdDyNmS4WglMq+z+pWQ9hKS
gdilmfAZPPhEEiXN5xUo8WU1Jfwdq6Y8cip6GZ+lPiF1h2s1UeoFxPr58cXEEn+L
+ReUQUWdBv+JxAHLE199KyjlcSThWRKvKnvyFGJxWYCFxmdjukwgW8mqJUSxcHBj
S3AqQFTY75gtKbi+XFbd5YfA0kTSLdHGC7+3RTp3N4LCQGhWQ5FzuBFw9EThsLUP
qCVu9rHSu7NW+ItlWI5XYvGEd5KIDOl6QYA3NRBP6EjN9YOpn4RCKbc7VMwBr3nL
lrEcEEieb33zzmNaopGGeQ6aCdk7yLjv2rUfIjJZHcwAnvBjMJXXwUK4QInQzSdt
rPhJ4Ieg9v/UkMSVWvF+hL7ZSYUYgzaoWtsFc9E80S47jYPx11JLxN5yoq1WeiS0
Iiv1PEOxOlzBP1BXFLqPZRYoNgYnjCOYOeNvJIVFY5yZPmv7LQmsG9tW2dwELcSp
aPsM1iAFh3PiMMLLX1xjmzvtb79qx/Jfbti0dp0dzFDQ3hIrJxKhu+bPjUJWuJCd
y9LLvLb0TH4brvV3vovB9dhhU8qvmXZTQxFQvNopAOj930byLU7rtcqp9EFHmFC7
OiHj4UHB3LBKCbfx20V4Li8jytuMj/pm46yKxpFfE4tPJjVFbDYUi2Od+3aGWapL
BzOJu4lNkn9tO0Ek1oFQfpzX0BANwYLtmkYUBc3b22obLYHqP8L1ams/4hy0b0kY
ujxqKKeYvSVUKEVECBTs0w9IlbWgF8eaOwqiagrxTPURvIHIasWY8K1Fd8a6UJJp
ceijlKSThrEt3tfc7fBrSmrGE5Mb+bRVhNPBVgcnJkwCA0aYjAoRGMlOUlncCtuv
PtahLP7O9QWzflPRAhUPI/8yExtOrI+Bu1u62fEbmNyEZOZenhFMikh4WiiA3Lbe
v3F3H/h+BoTMlFpUj8P47ZcduJ20/Pp++m4hR/VqQMYXyi1oS0u6uhLHmTGVPBNK
PB+PIIdI5wfRYsbXKaaR+fBDkCWwfaRnq6fWytq+rkv1vMW7B2HdFd+3NJpUipR/
9J2/9AA9waJA93oa1UBPWWBchGh838lyvaelTwu2tLDTSupFy4U97o5QkHru325V
4TwnxMq8iIl2KqABat5CTKpdZY9WNR20Pqc4RHYdVVK0HykQlvLFcLM+zOBxnSDz
lz7Y4lAni11Ie1HgTs+Hi4tFvivGyJ1TfegNtaVK0bNsqDj+SYUZSxsFRcxCSIFI
lqIjOEbdbHdKkDb1+qTKuPgoMhxX7bK+HhWxE7Z+cjZPKi17jREq8OEFzC9aawXg
EKNN2Sm6lPTh+u1aSnRG6rWymrQp6829QoNIIhWL8u3rdJsGULtyQfBvjsTAw90m
PZyoPLahHAt2xW/bTrnJKsQbnHgQFRz/J+B30TMFk+gIhNmqFck5Xh2hlNUBR0rs
1liS/ze9YOoz/aXvVV/oBgl0bLEqZMNqURB0mKaS5ZWJ0jPMGpNZJTQJsFpcDuTx
OZC2OfD0bJMthAspDl2xiBeH3boyY4o0UOqtqW8zH69jp28FOpOeV8qy/OOuZRXV
ssT2tsgKQHXQqPjoq2/SoIyShSGjYRn9NcEgaA2hAYTISVRee6caW8u9L860f4TC
jXVpOHJBIlCClV1e4U6hwjflzn+KmSj2GAo1SgMR2d0IiKgJK01R+jrWJNsI4pyi
IXYbPG8SEgeVDREl43xfS6J6sXOf6DVNiDAsA3+XXuyC6TNKoV3NTJID+RHkFnR5
dbF6FGesrNg375PsMe2x3KlzhwzAdBMAjY4lN67o+Z/qmvuZglr8pzL6OuZ73ibm
8Cmn1A30NQG5xMQ1oIKtYj9LJt/LFwW6g7lVBEeIfdt52ZIi0UV/UhAWZdTCYmBx
YjJ63kZyEk7/L+eqtXemRUibXzHN9DPRqJcxZhex4XmcGycsye90bJgVqs5F9NGK
4MAD+OSBndparA6o5+y4Nx8f2RIiZyQ3nbV9lXVUsUW4Xaf7YUJ4kllTH2UQlPgz
S8ydEkgUKyo6euyTiRIKMdW8F+7+gzwY2IfozaIUiX2TqNvQuCHfGcfYyqo9QcXy
wwOajTmHzGZK0oeiQN+7QI/2IIjgeb98Ui0212EcaRXM1VxQOakZo2ZpUxcU1T8f
tv1RuVrS3YetUmnv50VhnMfqnR1XGXz5C5yN0c3kT8rppw5eXcgpfcj+pLWx4J3J
R6Bo0llMYMTnH+CW0KlGO8/uTxe2//NCcm2/nSsW4Ek0QIrLwO8Tj4for8AMffNp
2oX5yeu6BkEkmPt3rJqnhWq9UpVogKtXqdhx0lFffbVbiOtf/3CwcijRUDUULqNJ
aeC7mWkDM+naklnF3ueRjghagq+/BkBncdaO0bEahZZcYgvM/Ju3UPBJsshLrE+h
3cRyL2zgz65kLvLrtCPbvecOb7b2NY0XfIQcmbT50WM0MY//TIWNQtWHe6fyUz8A
gJ+xj42ZvzHEkA5Wk7NISpVGHvsZiEQWF8YPWztq+t0fvmkzqV6F3JXOcFM6kj5c
0ZgeVTVPpRJKo4JxIJDvZPCIQ+fz+uFBFgOcy6lu97AhMkQWtpyJhK81xOoNVxF9
nKQXiclAW8Q+TeJAPxNmq0iE6e6SLAF2lsKPsebPlcokUXDfB7+kloz9BFTWw2Z3
u8rsP/1m3uX+Fan0LY+NVhoC9rpW2+kaRj7VhwUZmkqL+wvlWSh5uDZZ0HlDhUhR
wtHCOJefvOd0WLR/fyYBLOAc6NmfcGcHVB3A4TjR8ElvmnUaTcN3u9NqouXdBuOD
G4YTG9cmQUuU5iJqafSwezGoYGUU5EzrjZMg6NnhQwu+ZCQzEsSKfWMBiwpI9/cR
sglzy4WpBuoarNNY/WVn6fW9K/qQt0IMUD9fhvL3EqXyuKoeDaDfXrXtYRkfrkxL
KXCZ7Yy1OGVJXPJMwvWLaWzAN+3j5YslAbr8D/bVDfbhMINO599oa29imBPVyfkU
ejW/mQLouUhMZuFjyTKCCw0Rvo21BmnQGmBA123lD8lmlV63i6oWP9dl+6vSYrz+
3qy9aOl24dMd2Ppi94a+x75sMvC6/UurK+QnWr6c7aulXxKGVz9DH64QwQqJOP7q
nPodWRQ+89X4HTCqRVv7Jks+pC5ZDsyS8zdFDKJArjeJgoV63J0bA+ND/zqJgTTL
n90cE0drw782f67cGzqg6fQJGktgqTdtIgoMWOOeQByPP6sJ1ZALDhwM8/g5KCZh
dDeEB5el/RW85S+A5eRq23J3XHsoPelFa8y+SyCHpNMNLCsIkmvQf7M9EBfLAINF
WMmLObiS8yuQ+mAwVFmXocUVj5ECq3gnAwolW3ffuLZyoagrgwlTyS54Jk1vfGXB
h++fBH64qrv2f7/kn7ZEegEvEBAv7GJl18wSehEfZ2XVYIa/qaihQZsHsiD5eXGJ
Iw1U5c/uHxZpWBZIdE2uOCTgzknQlzCyi2wAOk3oiEXWlOxRimRQTE5prxWrWakQ
MRbXWOOxI3X3xdMHM1WdkeYYqN/lrWGIQ0s7OceitC+HFZgpMAGrBnB1YBZBVaEh
WjdzGeetrVGy5rIFdjKLLkZt7qc37cJTiNPpp8g/KP1MP0N3T2+Gkf7rpBzQpwjy
GKSZgyTkfwQTAdayapVMWYd6PqXyxSUqkO2x09q5az6SVkK55AdIwP5kenLjLgeq
t0MysxHU13+tG0jOPx4cJA57ezI8/ue2qEpWNkMOoABsi/G0o+e0NXGY9AoR6Xpy
xZO2Co6fQ+6KF+zgn4xlUzkIMQln5FoHSR9c9CEOOen02i5azReBPxxWKJgZ8RZV
INUX1xzLj07J8SQ5FpiVMS4ojj/cT82FHsA1LLS6MboY3caskh5lmVArntXqFiiA
Ajti990lkePMixsMpoIGRn4HqdYhGdKZUQJQFWXXyEUQAvDT5+MF8ztc0TrqqPTN
m94DdIH79JjiN2iTNR8en40wtoXvj/zUaPIaS3bMqzbVnlXwEwXksYY/BcA1+PJa
W6XI2BBosPl5pUT5lITax5ZieyXVeej1XN79H2Z4lhoQMMUikIIeVG7cQKC8Nucj
Rj60ctOoE7hD8QfVcSDf5CW7LnliB1mo3LjBgEczg/86VSbMAXxJODirxMh1qJrK
acpZg4JgYmeAdlQzNLbAp0xus58S1kBz2wUIRxcM4xuNa0lOhKHB0sIpq2zXvUoT
CPo+vsJby46iIJAy+REFsZasm849npYt1Ibcfkl1E3XAEB7KFe4Rv7maGcMZL5my
gtPKsVM6r3Lkz1Fl9ZAVNh/kWsyCU9yMzqtOd/wNeXVkYYMtGie4Ukv3xTtBJloy
dSZYN2ZtSzlKJvkecgdQfRmirZ3P1jTLLbChxq0xUIfHSkHDqk80Y+Fg3i2hIOs+
nROBCWGxrvLeLbKO3ysctAP3RnzEXC+Jghnh6ih+2krqyOtEm6SlwSnP5RqqKGyX
ApycaeXeyq0xOwE3ZVOVGtIqy3j9ROsang3TI1XsexDX0WpaRmVbYE7flEME3HH7
TQoThfbaE+um2gWAjb3MWnZIXNxcNOSoll9WaolRAXcPq9XtrjROja0cIy40FrFP
VFyB7dDqrd4FGo+GdUw6tNepsfNjShOf/w0WWYuIDjO9x8qRqAYDCxcOjaNCbwBI
QttRwGQUVWAywy/Rk/OuFfkOTNEPo3Pq1eoWbaOJWRNUljIbAoZ70tky9N7MfV4E
uEHCIsCUaroejn2TK0cN0VJZ5H/9LSKACH3HAw6xGDD2d4ikR3TJf62wu2hpU+Zb
FbTl6Fnjs/lAIp5NKrmzaq9+/4LqLBcBlnIQy9Y7SaZWAJ9HmvObz/9KvXYHvbww
m/mAsgBgmfDQidktKAj0slqtmFMD2zBicVUF6bqjxE61Gmn3elVUkUdyx+VUvjXN
kJXb0mmUuTqE0DZcPCm0WVutN/B/x0Fz0LT70WSuzc/Rrcr+tVY/VJKKF+3bE7cV
mkKXuVlHnwq1C6YOPSnlsMReqfHPIlkluZZ/3gT7sytkwlDlgqiEnjriEC7WEMbS
mVFCvqpUSh+BgSbN82AWBdMAL2Yva7g6bHKieXUxBFjKQsosmRNm6Y+Hb4zMxEyt
g5DQoNmfWvVnl3gNrzHTZyTJPXR8Ltp7zvHYIJhBZ7lc9v3xTPNFjrccI/gk+VqW
83thIVok1pVlh0tfhR6T5mSXxE5W7hIwzRAR+jHXsq4r+kRX97RCeb5xxK/ERedK
f4Huz2V3XjmVBLaPTPTIbiY0sX5iL/eB4BB5x2KudvafgXQxyWFFArAkcFcb5MyR
0+zuP1v+s8vSZ3m6s3Xzi52CRSJCHNhObiOH9hW7RaXlgE8ELTH99nzMOl3/+uyv
GlPe4IIIy5aa4msOFMzOYOnVSvq3BP9pk++HaAol6wQJIgo9vCgaIPRl6mYZCmFp
VxbVJc8iitSukoAKcU3S4tlilyXO9yZYXhTWUkY0aXIYuXxfl1AOs3rq4z0Znuer
njy6oWCbsoiVWeDNHwq7NKeol2VVieC86p5HdD2Czpvebh9C/pOSa1UoOI7KS+Zx
zMCYURhJyNoU5+xh2qqNW9pWmn6bkZQSSH+cKraEQyvkDC6Ieb7gc+dEOIFxSqno
/XXzC7j8AVL/YyTOtG1UoE8zeKoqv122XUEZ2PdqHlBCDJRGfvR2Isxvdsnjg/18
OKdwxvor6Dq8k2fBLWSqbdKBWYFNTpPfZ3cv9nEh8kEqM64z7W7WnESeeIVjSnTy
v9KVXXbE87Z7nq5+yJHcG7rxAaQbW+9MkyvGJpZ0OmuqinOQYRhXHgVbuyKKKEzC
4+SsSW2yxHD2Y4xUpB9txFaNUx0WGLWEGqPdaO+PPe2o/QG8AYWRR9r+Qzqma/xK
WDGeu9tNV+QOsEcG9hmv947atU3NZcPCqPz5lHHlMptRTQ4CwbieMndSMBAbvDN/
lNssXNWhtfC+r+m7K+MIipWKWvFPdxYE7iewZWJkTWPjMiAiKCQuKj/zx/xFYXwV
eqLa235pl8alWqLmwr+1MA14smszU/R4iQn6YPOksxIHHWEw7BZLZSe67pxi9xWj
UPU2IDB6t7mTAKaamTT9HE/1WEbHx7ZNuuU2LdLnny+Qa2wzZ9hELA6IpLGRIwTk
wH9skHmhYW8ubcOdrU9jfPi+wU5M/vzu0XfvIcT0vW/zYAy9S4jrIJILhKQv8aiu
ajoMck/wezxeqz0Gbhr+atoe5B7c+i1IHFyfHsHBBzQOfGLkz2fMx/bZJF86OtYI
L3S03CR8DlSGqqWCfmvbUq1PG9UIc+dIaJMgorT0etds0UT0zeXLAn3Azpcp27rg
Y/68SeOnYhpDRW5Ftde0c/rgvTaaY5iSt4WwOEhGuh4qWzx2W/g3DlhR4Ij0cpAB
9QcsRdixFbfwHVUIqM7s5KcVRe0lxSqzxlGNRalqd57+kElSKkNP6GBnXoPUgKaJ
ePLc0UPdjbSs84PCgUX55yCG2P4+jgN1vnQNbFYc6c4V11BMdLiTDTsm4ID84s0P
ipYzogQOAF39lAQJFdMQY+DFiO8Lxaps44FJ0d4lkis9YXpigxlMXRFO6Ze74SyE
NiOEq025iW4mGllfYQCTs+MjtKMXIYWEQOimq2ikeY5WjWHL+k2hR1vD1O011ZBW
c5o2nn28bWxg0yiBYv5P3DT5SZqsD1z8i0yMecHyW7+lR/oVYSaFo5n2SRQUQvXJ
HKjWVohuHeYTVIsXM8toRLV0RGGzmChCXH5Gmz0nSIvl3Jy/j9vPk6yqRdNQrI8g
5L/CnpPGqfZRMiZf1XrB/+7gk3Qax/tavQ5gPJKPwNk3/rHwqZ9zA4YWuB8Kn+Q4
vpAtN+ydH93icqiD5q5/zC/vOslMT1R/pwc9oIhg53d+VGNRSNtcPFatYa2GYvsx
K2aVJzbYjIUzqwbWK69Nn4g23JvhhgNlKQ+vSVMVTXHtMv3k9CLFTPs2uMs/7KxZ
fhntbTt4juoSrOQorQToSxCgYdIjRi8JpFzBnOjDMe7aud+WCp1xMzzlLsDrwOMk
1TxpeU8TdzNf/UyxJHKsPtws1l3KhsRDImI17LHIFroWEP5ELoJKO9We6w0uNOaw
xv9V7ZknNdbzKx94PuiEHPZ2hFdi7/69oeiLqInes+vTA2Cpu5DuenEc2qQrQ+5d
xeclauts4qzImDJXdjSJM/eC6wZ7QKdaupHb+gQ17cJKvplUIXOTjL+XImZtHQHK
oSveNu/B7rNHx1CUKkKG22UamOP3ANpYrmsg/8Dp7ZEu376xWq2Tu9yKRAxIP4Jk
EN4hvC7R2705IQwIMjUPWyK817eMQ6KZXifHHJfwWDaDj/4gWOegVwqHbjp9CcUe
vq6asnK3aIU9rnOrFWMzgBfugrHqjkvrlr3V2fiL5BlsFSjSklrihWCmD0F+1t/N
wM2wpLd+n+dbx+VllpJInBhiaY0KgzkTRWi0f/VQJho1//7lMh5i8FOp7t6YnN2L
PgkFXv4X+QIhUXfB7qNyNAeYc7blejI3ewIUe5A/Eef2O85bVdFR0FkmTZHwRt99
17TLK907d3KoBYRpcbbI5zlNHZNqOTkDkL4b6/X0Bg35ej046tZet1m+x86BdYsz
WooeMDZXVlRwLCQ4XPO5VMg0is+fIn8URLiuDOW/AbwGi14zcJEQHZo+7cmCtLwx
D+R47hM1t7KdpDjfAo2oYJNfVguEdmvxOTNJtYij5hTn3JLfbUi4eEHcT0nolHbq
lUdpjXhndV8RGf29Zevz/L+6javpRyUpPxX0oeG8asKLQBq5dM8fYte/CW3aq/Br
stuOZciHWtQF9NtEgx14gEV8NebRFOC6IMsGcXbHDN0umLqdAHghRRK57l2wlqr4
5O2anm0iSDecOn+rutWIYEqjAyiEeYPkuprbsHZeIkdGRfCX9qLdNiQLHdZScH/a
iYQRwpi660PHBHM9cj5YVTg6qarAGNQRoBmj6bHQGd9B+avAOY4gv6n76n6OFS1b
GS8XYDK6E91elV6WO/KU8jVtR0bKAlW+d9ilJqtaN20k5i+iUX9LE3NswTdZnAST
vgULF/nuQGRl7VfVaok+uP/CD13dgLAv+3+WLZ21eEMh//nJYP12U9596fN9ycZD
1+71OnWPOq62Aqm26b1CFksTWcXvDa4KeQ41kngrDDgEMpTMEog6Nun4jnEtoF6F
zW50KPURw4R3w/A0lAIWABFMAGrQNsT/7wOYR+WmdT1GM0MP26lwRfuMrgrBMPn3
ydAow0g1O9Eo4LdQCuoIeg9xCnRMGKM4VR/XbFKUIo5ijYcuqBVPj09aF+W6Yh3m
4x/jsUXuv9tPqxqRLzWleIWmAU8V6oYefHbzmixe3lJzD+DVfbw3HLmU+PoVPe5q
hzg0yrGE5MNI3KFf/K94fqKfaYEZGmaYdePVQ0Xwb27+FzABLXgar70s0AKiYtgc
g8Povl41vBXxOvbLSQejoTzfJpQ/H/VCR2dEnnlA2rPI7oWTHp7FsKFstrp8fjbx
7vp6SGgzdSqjD0mYfr0rfFzM8rS7mhbE7/9PDAHmezBdwCLYcz7EowsVa+HDQnDD
fV+kCML9H+8ZMZYC4nvGIPU+43BJyhPWkrsOk8jI9zTw8L1BgqXpvonzckRWyy1W
h5+8M2b01OTIht4QmgruIFYZn/4dzSqDIdz5L4CrHmtG6Fp8Q7cj3ptfk/w+vgts
YnxOSLCWxhUO/xk/kb6nXLLFaC9zt/+fX7Hdr0ZMdAqMeH4vqn6r4XfZB9WYwmBI
8X7y9t3b/3tsENSfYzvMkUIH0VjsZRCIbfKTworl/RBtI8d4ZxCANlsIyPexb5jS
PE+wE55nsRmleRGsOHCrP1sOOnlpAEnVoILvpFkltG8R3iTp1+RafZW4pC//4CSK
d2cMX1Xr74zsG+ok7CXYyBpm07vTczYRtFp/K0kH6Jvp49DiYxzadko+fqwhV85h
KoFn5tcz7V5WYmgtj8yiLIA+vX1UxlE97ytVETQP2/OUzkWHPbz7g7fdJibC6yqP
CrcgaVTdk2kWdWYKGpCLvORpMO/FDSMclq1HIxfj1kL/l83Eyo+PVx7CxKNmfpQf
rhxDDfJ0zSSvz+SkbylYy1xcrPqI/AwIEyLXQrMI/+dzrLXiayAPCotBIWyWqpgR
ZZGVLSG8EXDOJ3fTByqQaHQSTLgznAC7k8H6BcSBB4ET6kC5jrSWWMZ5PFoCQQn5
miKJAdMVcFK40u7ue2qG3u0GYEvR8+LRx4M93CZvsUklbjM5LpZ2yfOcBG5VjC4/
1ZLdz35DzhzGsTrP6i41U+7nyfatYHFSgEBcQV/7EBK0CG5NXK+6W2xji4q9/nvW
/49JVmC1qxpUue9dxlMChm2sgwnI/UggyTAgQmiVj+BraxforTXwfdo73KrzQMbf
fQMk9wCT9QvePK4lUct6aWEXRCdZhI9A/8iDglKd1bZ+nSDIeCW/V3rqFJEzfg4t
8vns9PY79ccPQEc5OUjCRCKAX+E44/Wfbj5GZwwltyuD883Qa92uHtiJxWqN5D+T
F4U2ebldJG6Yd72mmHAk5w+hV0q3elrV/JV1Xq9i5bzVMCn5u9U14c3sLvv6r1eW
u5lpI0ZgMR4zWmCeRU1E+uX2T4hU0kzwD/3bujDhmJx2UsPXcJLbelWsydgC8GlE
n1H4B3vZsrJpsqZfk0/hB4rtp8ODBsgcaq/Gb//KMUErM0yHoAkfHnuOSu3e6HCF
Knc8w6u3Bi0cuXQWTsn8AR6DjCkky4odEk5oeN3tdswqu8jxYTJ/bXWLfI2JYjc9
ZBs3xGCpdIUl7ehnxfsFB9U9pyF/DbhpoM+eOCZa7MFkyT3daI5LtVO22iGAU9+i
Wy+6kTexGrQrVNXhk57mOZaLsZz9J8n5HpNXLkPCk/LSx5MFZUZh+aVfIUm95BY8
6MsD+u4dHpiHVW7D6ojpN1K3qRqitmDV0M7jvQVEocKhc8vw+0u95HVbMlgG2qnn
q6stnTeGcMl1SJ3ENkJKX0NH8ZzZRUgwru0XDo/XP6zuxYc4sWQ74VaUGMdfhwjr
VhSXy8RFXIJvxrJRjLUkVLprnUBwLpiLj8eBTZpHhTqI1VDYrdSG91lkpO20Bdqd
MkvUqzU75TF3LG8/EEwqhIlL/rmo5ew3wrcRQcx6s971tJzIUJ01u5q8vNeGwxvK
epZf0tpFDzgheFbHzGwEfVTXIRKN5Npz4VMMblI3la3Fn+/1WbaytUsH6THUONgW
36iM9JlryAvoW43lYnbiDHmgggdqSW+n6vcSXcvfFpa4JWH4ORM/dr65Xzknhxnb
zGFONltsZKZz78gd7A82qzUxTZuL23cep5sGoUnZ9ot+SLhXDZRL6QcVUXVuMN/f
AIGtTKTwfsnWO93vvSRXfycVjWZkBUZHEcH+auBG+Payh9I7IcA5lDQs9GHoPnmO
4qSOWBbLWmwrcZIVCgirXUXOsyuP/kHj+5OvCbmVyspuYiquJsjSAWpG6MnP+7Xa
fDyXOM/cWGK2Fskznp9bJ6aBWFLUasLFQCcd0mdR6dHr54UAXwBMABAlZukgw3Vj
cLD2d37fjPC9aB3oreYGgvVR1DTWITF3+2S298x2vMLntUdY7IpOBr6nEoSZzQr0
kWzu0oQvoPIZ2pw/nFf2+aU7Os2ds1FFA5jLMcCA9f+WnE/78alOE+2V6mt2zm4t
Av8Eg645JQLBA7cNIjkQmB6yyFqbgmA9x/y4lzevL/Soo1adtxOpKqpXyEXHCpIv
Llruu5gGi51c9oA15N6p6F7T5OpzvdWmT71igeoVnh6B+QYqESalxBp1+eMJyYE3
pRU8mrwCSZIlKU9f3cu28IOd8w3+4ERFXGMguiOHDm+/Fr55laasii1prRZR8uQl
aIMdYCLuVIcWmoKcpwpqCa963YO6+FfMEjtZC0W4nZbrrDbfEsI6G4A0qg+pwgVD
1owwCPH+o2g3QxrWRIlBnRqFItNQWxpQF8+6ovFD+ODbUcN8K40C04+PjqK6noHg
aNEw33nSDqi2SjWXbEu28BgVxYH5A+YgSUwHWSiJGnAkOtifdHY8/7a4iJTFYWqQ
YqsgooKwdzRtmZk5JS+EDsy/WEULp0x930BfurY9/7+eXAt2hAlznjrd6qTZTXlS
o4Azr1NU3KUxn9wlZIkPX7YY3ozfWNXIpYGSBOBWbcEm6if46wyaGG29Jmg5qqGZ
nrtPEI54Ujdwh5L2CIQEcg8aZBMGxPKCQgCk3VF3E1Xa9H3Cj4Pn7hKNdHCq9lAv
MYIddaIWTUkTZmZtf+I4hRPMPvGqTt/HYn2G84rYyJsl6fZI5vV4DdorFDP5Kzl2
ITRxjYZq8Y38ya+YKDS4OppiJKypWvGES/W31SesQtKu2q3O6oeEml+XSS8wYbZg
qGODAQ7OHuJjWq0w9QZxf76qwQpzy5kympG+VTIZraW06o7MwrwOtxJUTiBkr6VG
FnRlp8gJjSjc0SF/RYZxcv84KjZHNc2HQQC8Bfky6IaRu38Aj/LZRuxnFTAT5ehk
gx5y8mHJgq+Bv1euk71eUesHB9EQilvHkifCRt40KLuh5EKcjzS0Q4VFBSxhYsey
c/yagxXdNxSwpQLetdOGMCOu04+jzwWasAwneOwJQQf+HtUW16JXouzCGYx2U2v4
b6MPet01T7ATQNNmZf3F5OPKmkuV/Ew3rcrLnmPcTe63qHe9aZxZRi5H0MhYUkM3
pvDnELHrS5A7c/5tmpQdysj37N4zWRCHWbUyWrgmzexSEMfLqNrnLUKRWDvMgTpw
bwdKTMeSvbqHrDvAqWubE9TuzFrhYRf+XbR024mirOvxGo50jeaz4Z3sTf+Q7Qz1
eywSgcHuvLlnULDv1fyrOsuVR/LBWY8Fi1ucRGpYdaAfm2jbOsU255xMhlh+v3Gn
WZ8mu6prXtPjV0OcJ+OWq8gXD8Y9934mqUFpdE57QodP6Z4FdogQvzYfKhWSQt2n
ALXa2IMT8NC/Iwk+fZ4WnUV7tpmY8Yj857gXLyGfprJPOLQDFUBa+kIQ9OgV+yhV
+alR4nRVo89iQsmh45MnN6/PMLdBLOuktr0qzquTHJBawOrT1B6x4ot/jmnsTvb5
Ye2FWS4cFL1+Myg3dYUKn6D3O3q4x1PSGjDOXGfnYZpeWs8BL1ufdQQqro4VubST
LAzSIP4CNPhYkFIrcrV6P6KbK6wuY64gE+uDZyMDV2nT7jQ1ZUp4limJSAXRmqhu
qDg7bl55poYEe5cwrYnmoHDn0WrTuHG9bv2ogfsmgl1pxn9um1LQjw8a8uyH2TXo
5AqkYz7rJ/DJGWnjwweYG51OU+ij8T67f+A/FRH9ityubbwci7Z8qsYAig6xBaUD
VNIQxLwy+FTDEafvg+WJBXSJ/xk4hPkv6rlB3xng7FbyIDdf2s5DKaAPTWJCb6w+
e4l28b9qvVq+Hk2cW9ufTh5tJrAzeD477f0vRGI2BZb3KaU1zbznMi9Go5wZ1S20
tiDru9HkJLWyKvcqFojJvzuycVGv1L9giXFPSUGu1jA48ZfJTZCRoXJJ/9wLexxw
A8OXDcwgFu7KkDHjpn5qZFgj2M95cU0bzF2Rj68NFl89BC+B0lyrKahl/nxVmJeN
EVgeKQG1HPrIe76QxPmG+jLBt+BywSCjWnB68/8ahVrNrxDVacuiGe6Mmx1M/whF
GZ7ICd4fJk6tL9iwrM+4cIqhCuvnWddtt48lh/fHU4j64qW7JvTYM8SZirME4aJA
rDs/d/CxRHdsLLEp+EnDvvUVkqtObfTR7LN7V7JPcp1vE2ei+uZdRHuERrSNOhyy
P2vtzLfhrAfMlyDeiYWMskMKHR7+rnb9txPd5rBttkbJQ7iUQS7pxKEn+QqgRXVL
z4b8gyO14CJGrU0t4Kduj6uLdp/1k8yvjyDoKp+0bui1XxhH0TXp+Axix2ds9ROH
SOHYkXSVFDyyPmhWtIhTqgcCzWVspEFN75N1PBc8iF6uAVDXfsSaG8YMQuPNtCPM
krIIbrCcwKw2rq6s7Q0GzcTylGS7SaXaropQiVe6noGbUxd9Q+9oMKibbeEhYBK7
n3Ke2+wh/xIVraJ+89/ozIT2YtyT/w8Co7U1xERzdFwPd9T2rbtUsez1tjaVpxao
rfEGVgL7sga/23CR87Juta5Ock89dOO3B4F0M9pykFoE2lA0vJJV+Gc18WCEOi12
Dh/udpWx2+tWH5lAwtoq4YMYlS2ItKA1r0DZWArjcziX/oTeLuEK7IQ2HW8VaBVR
vR4xRfQppSXOhFdkR8Qwxy23B/4LZnZVIMIhWjKHMI/mBAvYsGLol67R8cl9vusR
Ra7o7u+s32xU76qE3j5yilYbXyn7grvD0+/SWituwexzlHxkweAdA/lUnGhRT2Fi
deDRbWWrjAOLto1RVQe8VhU7Y3l3bFnLLJE3soF0HOfcNk+dLeQECfEonY/HicNq
HeDKUXNXQtmoP9bDQrva9tRpeE09YtXgFsZUa/9t2ESl6t8iF9IXebfTUREHghE3
OOEOydBx4VI0kcvAYzMYzaWtgiC+ajpCOSFsbEx5yv04/wLDW5yjVWzPYXtiAjqI
5aUpSaDEDwJk89FZMRNhsMTJRNd9eR6g41lclkI/6IlOBfze4l0pmn0J0TcONmHw
Fi+1JnZ+vEPe18ele1qlVo15upKLpnh38SFi1BOcLFWcngsUvDlRb8CtJsZrD/G8
0U85qd3xF5e0+7JouOhxJqRRMqDLC7eaJ+OTfG+QFMaYrN07gxs/W4VUHvINpW/A
LGJ8stweQ3wnQhxDu66yT6nR/SsIIv+FcqbrpOYBddiZlyGYiLc0JMhY42QqAt6D
U6SN5j1tB41RlsBDasyCOxCon2gPYLluHUT9UepFpo7Zvyhw4tC3rw168W/8sdhy
o8FmCJGm/aW3mQScknywZyTuKGrtL1xzVWBjydASgypOE4Ds5PubiGeXwcJleBX6
urtH7omTgyUyrbObpLxxNZiv7o5yxRlA+MvepmvEvKMe+1ytU9uI5/DSUc3e3PTN
yScM6OFDgMJFt0Vvr/IdYUWTAozBDXcLoZaxITWYfZ+tFH5ku1HlaB9dI7ScMqvP
oRxCKcLA6G4lg+svOeg11kwEWw/wmncEE5izDgfpAcmTCNk7OtpcpZLIiAdXWTO+
ycgEb75/IDr/jJEbNuKfj6oOFhzRGf8xKcKBgLK9ZPCHkHvwl8Gz57f4WoFhEgsJ
7ljerXXNxzdhUBrEViiyIYY8vdAMV6V8CoHinjAdg/xo+OsdB0bGWjCcXXzGgi2F
wKh7/GA458+jq/H+i9P21ruhMAkITTDONk3GRYKw+O7LmvRLG6E9AzzkB1BVvhbH
HDQafYnz1ukhJlo1xwA7OlZZwRaeZn+9Yir1NhMpKOzQLPstLm06kesfjZqtoFb+
qAWTwKfpZACbjn//Fg0WSbu1yYWYEjfdKEiwP25Q1E5SfmMbnMhrrQCYI/RyqsNw
NR2cPSt27q96vVz39jI8yuzMkpwDS5vSFjA2Xva2kPWwxlqRgn1HkJdEmJbp9D4k
cOQElBeM/dnKu3SnvfEd+aQbOkDICXUWqc5GTLcGQ0t5oHPY+4/AXDPhMKhACgyE
R633fEoLOD4+GbRyS+UUi75ng1Uso6ecJEnWj2eYj+dNEmyjQLENAPz8jfSIIJMe
GlG2OdUI2Zy2pG+B0+Om01zdw5b1wKAnUkf5aqvgz5i3UHwi5tfGc7SCiPh4UkKt
FKqOszfRNH/3bDg0Lt3kjjg0bi2Zbu79xk52CnqP7v7NT4lAIQ5GtO/AoFt8hlTf
LZQlNOQ5ZM1HsQm+Qh+Fd483Ualns5Wt+9xU0fcigayS4vQNGjLIqCmSyfJhspPc
6U/pbPGjHAY8DwCLdI1jhOq7MIeqUAjx2H7ZONAi+YvhSIYtJxNwjAFThFDJMs74
OKRKf7SLOdKY8h8FqWsLwoPEeMjKJzI4gNPDJRbp13t+zeutmcmaVfHkk8HAhSGB
Z6YMCYgo0Qq2RXXuDYYNxJzD//Vkifmv4IXh4SzLfRfhAXcn5/BhZiwo/D3DgnFi
3Yt/yQttJ03CHmcoWpB3573/N81uWDw9Kin4LV7po4Ry1OAr3K9arMTT3BRM8I22
DB3vo3HT0ZDuevNjhdPCG6vybpIKtTXYCf6dzLw9CLXAE+MtrZ5Bc1UOQ3KqBhkf
1QkFd/ZPONHMvCCJ23tHUFxzkSn8/31hsbi+rggOzsZBlGEDAh7F30ok5mm8pm6y
wkRqTXryXGI65a/pQvma0ImkM+Y0UrdQ1eqPiygU8NnSl+fYkXB+M2tqzDT1aCts
zyoRtklT4/Z2pxTFCTxl6vLFXPtnbljmKf7NktmRyLXEEhBqhSbajTEk/cV7k8En
1kQIOrWdSaH1MsqL4BJEcmfz9dhwbo3wjmWPpqBRuTyNmlTfdgpsrYTsUImxQuWq
1rXS4mYfSFzD+1QIbSOPpEeb931WjnFmYlHHI6RthbLORobN234nCYhsYYhNrJo6
W5/XXfPB4fLkJ45Ea13LtDnu+LrZfSGEQHh9bMyLHgIMsQlbhxTCsiPj5lvzYkIA
HTAgerSTKc8TnC8H9G7R36ym1wqgLb5I1Hen3V6/TT7ASz7KCOcNA2z984eDks5i
lmMoEeY8A4kskp0S3wlb6Qg3GrglgTOUmYjhP46At5xMJCsbEDTqaHEgUEG1jIdO
PDh5OmMR/SUA+gr4b5wlYCS9qtZ9EJeMCdLCbpjGLLmq1fy7+TAUl8YkE2u8hcYW
mDqu5H0AbtqQn2x979JpV7AcsZGz34LQVUiyu1A2wV0BunC2obvb/zKiQ1JgKITb
0ubxUgbTePXhfOweakNqeThW+z0xmgAzEF7v2vjaPeJ+ZXhA4KutQkgtxHeChItC
hCXlqJv0C4UbhA2e1lZpsWiL+FZt+vnFJTsnFxIW95yZC+xB2B1sYXjkynm/Z/0r
NmBEi1gOI2UVF9SP6AShlUgePbJ/UWi45FV3XSsR7DTpwaJvbesxpFQ8MjLC8epp
hFvMGDQwlkIXbjXo+QNNxglaIH2X3A0M28eKzmnTuTviAqOGs2NbijoXqWwJ3GrM
1LJ15pJQwQ98om38vdiqgYH8PUvEeOCP6o5u0J0WdM9aRtYx+k9AKPm/sUJCjZok
Hb8YM1egUgTXQfMwuDQqJENnzv3aD497ywIHC7Tj3ho7FEGv+m7uBBvN15aKUcTP
bOJFmPF+60LYfX9Ncg/1oNigitREVQV2ww/QkK4+1sMNLNWWGE73sYppYQ3Pj+KR
UYR0stm5hky1SpMfr4xAXtxQatUCMplvk2mfzgK2/llqYtA9uVie56AG+npZylME
TCvC9jxJbucpBwhfTAiYJVU7p5D4OYIvm1yg+up7ICcNk24tdlyZ97sgNwPDyjek
aHvNdWMqbggiYlgjx1Dqq5xPcMtYGvpYqDQ+BE50QGmiHrm0SsCUGkOsVXas91i2
hD2UL5F9RSYfFU4xAbEYm7VT1Xon5WKDEUpn6N7TiNUYwu4kXxM74jOIuquB0Grz
HkRRdpvP40zpQhy74HfWAPGkidmxIpS68BwVQeK4dW62DrNKSIO+f60FiEXD6wHr
Zq8LzMAK8vwOCmxBrGAwkHVzK8vaJH0OMBwePhdMX8BzbkOz+W+m3a48KJArFRQX
3tDejcxng5+qGZ/Hq93H6IdYtkp1fgkfY46WeZPaczedB8qo5nIrD/KbD3RrKW/6
yN8s7p4qBeOD8nSgoxqz8EnyFY2JPwufpfOCTeJf9/C19NN/G/M4piFyGzScLncC
QiJ/aCHrfeZLIUlAKBDIRLaXPL2ujr5+e2Su419noY5ZvbXrRCCzylcYvJLpwV1O
rdNKG2iO+Yjk0A7I/AuhgMJcORG3E6JXdUq2kExoyvUPcIj984Le6t8eS4tT9jzR
dfbzDY4YLvT+HgAVNtaCiXpOOsUMdrCRUdTsdYcR6x+zo2/dOyqLAAP7V69LDLzO
SgWdV3/Gj8fVASuEDfzt08l2Z+/8SeMfkw18lVfZoK4D391NjDBrMBfv+JMwjF5s
j9u5Nz8MHnK+Mo/XEpNPDPyAwOLOKgZ9zu71q6p7Yv2TiKFNoZJjw4x5TJz4zzLv
yrq7zjkxOzbiZbBvCOoekTrFM5i3LjFsHo3jVs/6JYp+fv2DCxnIMpuQZD4UeRez
ZZiE/uZ6GGSbFY5WeWH9+K4Su6XF2bwn7ZmD7EqMGUmZLf8pAOnldcRmY9SJ6DCj
ZgHydnQA3g3frJcOG2TKL4+XIcGpHx+EdCHM7Ee2p+W1VCLsKRqZLYPNq7UE8AOL
nAVoRBViMQmqCTbIA/I0u/s0zwXhP8MrF743dNmzxGcwc9d9TgcK+J86+O+1dbX2
N4iKvgiM2ZGjMiLmh3pOUIB5K8siWyCV8EHjOG2HcnDGcRNwEetyZ8PjWm4wp8FN
Co79wkjXPXGeGxDofX4nOdA70mPk7wM8p/bUgGsIapqRI6uhkqwNnwtqxMWuc7dH
9FR5UK+9DEu3H6RSHPxcLDoQvA2GG+iQtxucnDMdYzIz8K/JlZmJyeS9OT2LXX1A
tnbX4Cq9tNwUraVbOiJ4HvCfwdGnd/Rx7xU4QBE94/TlwcdBwmeQs/vnr1PpDhjV
fWA6mMCVp2nAWhvmxytWDdnZN0aknYNj6PE64L488s5IJ1MUtxp/MUM+uO3H1ydy
YGXgC2a4JPHnF+mr44hZYlDf72SLywZrVA/Mfx0GvXTRYkDR5fnwVipcX5ohIA8+
cYPnvXVJhyGDJnLF9NxPB90p34LOIRNcmVlXWBVPOODrYv6TQSQ3imsaC0r2lxSN
ampC0WdZqfDMgrcgkmYS0YUSm/ibjnGN2NZ0ZTgBzrZBpcb/RW+r8z7nbhs4g4JM
BIqOMx+i0/W98heOtTWpuzKk7a3vTP2ziu6QlTO9scOlgBREjExov8YOzvroP9sv
zd74g5MdzLO0NSsBzMUWlNdCckyQGk/f9RHt9XUZTcVB2hZAQx+xLNnW8ceh1ui2
WqdhaFhu89gAJRFiZStoQuQrV4lZYJu+9nDYxXvBWP72Cv8X5hRY/BEA0zjM3aVb
SKyVwLyWSH9VHXbbqSSwxYoTQ6571xCzjEMKFe9/1liUpszXaqe08Kxl4dId31I0
NkTVvGdU/HQ7+TDo6knQMp1C2lASgVswIMPY35lAz3RjRiTJYXVKoaN6FnAxCVqN
+O955CWwcAOGJ4dJjgS0Tw5kGnaII0D02w+xFMfJ5qQvaBliNxc3ZYhwEZgmH9aK
LLgcmCiRM3i6OevEsE8VcoS3hvnnEOPqNv3nGkBo3gTzTeS8JimRwcuGpMHwlmOU
6I/+A6sxR3vvgFvdH5diI9TmMzsnjpES//2N9XgNZhXOEhy+UMrSaxa5/A4+MgFs
/QN+Wpwj/uz1viUHEgT7clr9B3wVxV5f/SnSQIXiiNsJwNWqlDtwpuFsNHpc8xBm
k8XZBJ/4kkV+2t2Y5fGzwUM5tPfo5OnWzVavM3d+Pqe98Cbo0XzcSnAGpcwMZ1YM
YGCUPuhFtBwV2+7taQRMUOfS9QtNSGuHlzAaoJ3IHaSEzk0E3u8KDJMN0QlFjT/d
yQU2aGln8W+vYkyzbOkv2t2q0rxPM+kMcwXM/B9OYRIKYtN7aDekCforI2l9ZuVE
V2nDoSKYW4otIEhUWs0SGFqS062Dx9C+5u4Gz8o2wtRv1PeZBsUQOr5jlaOVvZCv
95NqIlK4y0ESVVQd/U9NFYM1FVnpjToAZma0X1NWW/diLqz+APfwDqDr1PD2JO6h
8NTx7D//Bdurvs0r0LZA8VG/a8FGPCp+fnTt1A0yEOFbLh1iy4EZCn7QDi432RAT
+9xpsYb63oc3CEFSdf+d2YbvEtgO5NXy3IJh3rKW0cd7kw8qs+yoCTuX/b2j7hpK
1zMnI7P0wHiBuqzoPKHsPNN0JkYM7NyWMnoj1lMkVdPLP+CdWNYcDOQo3oM4t37L
jlduHpVN4koS87s5Q0q76Co5VAcUppZj1RH2fhtAQ4OANbQ6xGvxl2cB6loFl42Q
Il8hv+Aw+jhDWYBgXhsUx4zWPJaBnpbyq5GmTl1hDrgGKjvHbj3TN2guxIZkmWse
pX+ibmrfKBzBVrwGgG6C5w26Cc9bpig3rOmUpUOl3cLYikHj4hXn5IoF3+iGowBX
/WTX5n1RKbNjDRysdp+bIMJR6IePzkRQGkbITsjdFm+gmTVEQDbDDklWBBh1BE2O
5j0j9aqw1f1rtN1Wd6T3QCjKYPWvjp5zVoSaU/MD6qumVAD+kLpTa7RJQRQ5Ovii
l64FDxHeSt6ho4OTl0MWhepH9qE4NB7E+jfEF7yHAXCUKG5s3Ng2MB4E5wDTJ3D7
f2hQ3jpGWdq/agsJsZKvN/lIigPQjG0eDurq3AlsYvd/lvdRoOYeS79wEm68dMB8
x8lmG4KTmfDWCDOSEeZ9oW6SGD7seHeyIvXzRchO6zjbYB4vgP1/8ogQuusXVVlZ
qJVjwQP7ibmB8N6UxyVlinSMCc1/aseO436sGwOhbMIi+i/szfgIp3k0zLi6gyOD
Qeq1jTP3s3euYIe9lo1liYmQrQGi6bK6zxU362qYi8I2Krq3rpohw7f78bpRplMG
HOWVyBI6rTXkKjTiDlv+8+Oh8tMwJv8Qx5YeTIuNN/PnppXKS4qT66NPck/SVUOZ
DyEgwAkpn0bubH9cMip5M/mSBT43gV4G/lSALiYAIEwiHqgGAYwOOfo5Jeqt5r6g
LsHBflBZUcmzLLzLHT3ZmESuzRv4mJ/KgEZLs6K+TuQTdLEe457v1HR4JpuUtkIP
51vesgTZV3SsfAqZbOfts5sQwB6KnQpPFArXZZAvQaOTanzpzyYYY4Rob6YWey+l
/WDoHOFHN/IExE3ymTY4IaWDeNaBuQNJjMHG5rBLzwU6uVfa5hJkw/ySigNTus00
ZXGfYb1feiKvXCp/ej5KK6RtXGLHM88ik/aaqJT5ImQ20sci9sWmd57cfrkun2YL
w25xnsVUDvTro8e6Em2/A9Wl0zs7+lUCeuuQTIj32i8ITv5KHXg1+ZzzQGwmOQON
18rWw+ydZvMOQO3t+TBYsfZL74NKOU5c169d+7TewbgABp+qQqdEKTMnmSRmemK1
0wMBt2AeMdrm3Io3OiNXnvUp5CJ1KmNq1ri8XAm3TKZKWhA+zoygywTieURxBPw6
vvY7T+AQqU2gowKPlWeZURkKyx6ffXxk15CWM/mcaOP3fuNYeKKapnM1kZWxP9lC
74PvIYDtmcHFRkw6biVNmkHJzRxNdTlNddP7ZQ21wfY6IJC1LdhMZTrS/LjfNFyx
7U+uriTQIplMY+E8VF1M03PvCCrXFtN6OnxZsURpgwYG7S/OjoTVCpo2VfpS0d1g
ey+1fx+UQ0ptF2nT4uMnfZXOOHOvgAX1kw4B2UzocGjA6tho/rrHvezyqBsugWYr
AtiRrmHe7LrXyAJkWYaeYszCys2VPetUuJ7jtBB0BPHeC/WVxJesZpxMaArG/LKO
jhW8WN2uuZePzdSwVRv90k7VVs4ISw/1d6Vd5n+BdRLjT73/HVrHPrQ6vycpeIR1
3RUjDHy2l2t2UoMW/Q8rqb82akf+ly50tONQhcYKUTXdTZ2zZF8QWmLXGbGfQILw
l4hLPJdv1goFAfRW5CV6/OOBa0HePacmtbq/nAt/49W6DhAnfssKpSyU5yJSXsjx
WaVkttBFgEYxQyJ2gAcySZsDI05ms1zLPWolU6BiJNJUdsIlTcEV4bFCQZyVmrmH
GQsVM1EIaPW8ULuDzEjJEHZ3CJ/+1pVLplMf1O71eMVqT7lUfhrIqizGb4QaUSCg
3XoT+tkBonASq6752y40TjHHzWs6JWlNBdTyq5iGTtWESfDy6cNS6lXeRjUwtnLO
T1uhvL4FWzeplXfuA1TM0cijacgiA68sraVaBT1wu018RsTr4Y0iDbWD5WOHDx/P
Ohr3gKkl5UNRIOhvD1IlHeJdv1Lj0sjN3sdkMJ1t2WkA4IIgsoaEZ8QbWnOBzZY0
ilWaLI8+1TaW5sVNANoVkr0xoZcceXpZUPToScNZux9geu95KOBgY28mRw+VgwBF
OpcVe6tFbvrM2P8bts7A1qynvEm7cgQ+1fGMJwL3rizxZPUgb5LnqORuTWD2OAUe
557mRGsf5ImzlPjISR/JWSjme7KfhixoLyl4MPd3rsf2KFY6eMhlQf/0bynDXkYa
GR04tBOvlo2oNvDoTbD8Dgqo714NCbN2vjTxORhkVWGg3Y6htdgMEVgNhOyA8gyJ
UNIPmc/POFsZyriIvU1XqFk99f4LVkPb2E9CTvxhFyTyOvlapA/Lt7lEfWLVYoIE
IQwGnm9vrjFvoyvP86SuuoCNSx0IEqabKX3VIZUTLXzNR/D2YDbvkTojsC02QzHJ
jKs0j/eUlqqWtGj1HuJYRh724W03AUaozZ25bHBlYnR8PMLXw3gSc4N+iDxnO7tz
gNzNXjiYjS+tsLHCz7RyL4C6Yzbj9NHSr0XU2AK8kSnGF+whh9S1UI3gIeNw5jVC
4GBxN9PSnobxt53dsjXCbZ9hOCTFHG/fGm/D/1omaiHQaBS/z41QAlg2a3D2Io8u
jD2usPf3F4Vre7pNoUpavX7QaPb5Vl+P8CfgWjy/6iIeys76XGkEPilF6HLdkIdF
5DbVjNKTMBTfnPLIRP78OKN0XIPNqaI712uUCLDtMt8kmpvUSuXCSGp/JbZm5Pkq
GxI5usEH+F5weOR/atiprn5oRHk4Ml+wRWMlUH5MW+WdsR+eW1M3thCr4SgGcFwq
JMdQpMNyok/8Z96RBK39cn8aXnGIpxKl2IZLnVudlaUKXBKqcTXA3G1We7e2ntG+
FE31BygrvsyoEDR+Trwok+pFMnHhgiYwkl4R44o5rJGMJHPCLYj4BAWmOv0DTFsf
HEOm2JEefrerzBFNK8frSCBg0np3knLRIFOGZ8iH8Dlj3HVbHdB4FhtjnX9zlwXk
hGXEjBaKQdzRTuBIfMazfsbV7ojjEwIocj7z0UxeEpk7pGYWhjWLjFFiQfblPR12
//7vv0yTvwss/rgNcT7XhrWwqouD5fi80iT1jAp5BiMf3PZlzeb20Y2BeLvCsVjW
CmYDtB1itJ2MopfGZ2V8u2MCTwxKh8V5yT/u2IDRvwT/eFzibl5q4tNpPMVfgI+W
uzmd2igr8b6BLpMd/iOJ+dSVaHQI1UHaNlBst/MbKwE7Driz7l1W6crbvQVII0gW
tQG9JUAEWqOgLcK6m8+6rW0KtOpE+aA1qFRJcnJjuTljgO67IZTW4VjkmkEx2fhG
9feCPI6QoCm31jLY1rvz5I6HanYCbL7B+dECh4uBqfkPDxNSU7U2YLsdZy3z4t8k
Q26PlQzSUqzbqjrVB+HLSr8yvE2uYHeEP8rPdzFZcsr7kX8J9bVwtBSFCt9ZYcgc
2cjQCtGaNgMPNvY+xFpc2ElyXSV1gOYPQmtQJRqc0sLpL980EgF+aTsGkGI3Cevp
B9uOizsdTpgE/Oa3//SX+0EfqIato5X2kZsUBehHDnrUPzM8o7Q+yxEc+HPkfX7y
ZhY4LyrhQ75PH8O0/ytg4tVDGRoyVSHqKx44TnbEewIXQpQvCGl6CeClmJBpDfHU
ZRGQmfsqxra9ZWUQeCOpZ/ENk6MHauchwjkx2ietuQirUYdZnxgC4QjVD+zKzEvL
+uery0lXtXAZVO4OX4Bh78n4iDlD2p3J3i+lL2iWYUHaTu45rS+BqGTgvjmnk7Ke
fHS3+UutfUEu3iV6Hf9DMOoUmFBYqM8R5KTKpaQxaT1suW9UmRqJ9pHBCC3Xl9fe
U8mkcQtzHBvQeaSTRT6DdK9UH7DPPJERB9nZa2fM5j5eICrtxS4sIhwwZUp1AeF9
Vnm0jIxtOLt1dV4iFoxviQ9qNIdQMYwoJz2TEJn99uu0CEVXVUWYNOzb/mxooq+W
E7rBoReuPf3izB8TnxI2bNfIZYc/J3z/jeuSxQ9nkBFe2X7fhWMm7nsgMvDx8oAk
my2qUdJLxZo+NPqwBLZmELeocy8QJC4YOZibugn7C5aMUWldZ+cTmmiNe7f5d7Td
0SIsJsUPgoRTHy7Jir4baX7nojBaLwZ0xg1q58zkL42foVtft/LrSgD8bEkiq2Nv
sHnsTNBb/gYb4OzW/qdz7aXSZ/h1AOR9X7ykM6GbQJPz/kcEWufN11WB2vfnApi3
qOJmPCKHw4FhrTbAy6fjuKIqfHGqw/rKLqpFEQL6QgGlk12SgGm6sdofOb1Q1feB
dks5bOS5hwhEVM0D1U/Ud7c8uazg9v0xm/1pFmTkWohJt+kfvyXMwyKX2JdRvuns
7EXXmynCPQ2l9Ce64QPkyzo5ahu6cp1Y2iVQrzZEMUpdzd2AaicnCOw5chvUuul4
e983Ux161HJN7/rhwjVXtptvDAHi61V2/bqEY9IRMtKJaK/DUnbv8ZFbffhylpaQ
1zLVqClO1shq1se5G3+n4LlbIXUjp4h1sb0VYQUW0TEqD7JYnPrS7pzn3ZHJbO2w
gn3EOB3CHyoPzJx+2mUzhqyfVUfRQPBqsHfzOTghrTgocf90h0lkCB32OnZF+R/m
7LhX6I9MmX1ldzm1VVHB+AtxzTgnAOhDAWVOFUpJ+UikGJ6hC0qLYPzt1YPne6/j
taW+dMppvR1K5gSAXPYf8sIT83UYKzC47mfWIlI6b0ZnewtjAU4r4iNtyyBFvnvp
q5St2z++WIJrihKQ7XsuB99xLRIZkuiFnCIjWVcojZPx17sG8PorgkYoXEEDCg47
rHQ23Ss1JPzrCx430JDNBzVd63beXkhQDffNIPgsgQk+a4b/LtlJq+le6ofoawkr
zR4FTflhjX92XjZgJlcw76rIIr0AaaaLi4ZuhoudBX64cR7qtr3WsHbES1autqn3
Bnmv3sk6LR50qHScHFlNWWujDYO4ZcYegt87Ro+R0CZyGqvTpMwb9VP+Sw96e3E4
yuo1CR8btxbFPlcdBPfxyld/MTibzOEm2Y2C3fdNXKkxobEMjx70PRuOfQ4cKVV7
g7nriexXJMhTbZir4zuGpqdRXUbkYTChmDer4oiRfuAS3mS2wal47xZsZfKPLcuc
ctZ2ps0WylXjRBH5PLqfHgg0YzlSlIQu4n3Zi6TfWqxdLhD42FZkkFKOQHiTM/eh
jrOuApXFehWR1QcJQ/d+faDJKKBzRq3Z564Yd8Sm4otvi8aV+QfifiHyBhAUCEJS
5HZvEZqAaftMjMcV6MAIDP5/EQUbYarnAVwb8KDM7Fct0FUqW0Q6Ujk/cY02AUPF
nCqC+GSghrN84i7pMEFGwNrn2kieVLc0VokpUjDVjmHUfNnEwgtEfLDPOGlauRst
VPINysQXvvDJBhTA/44JW9bHeRI1PsTtWCPIFvSy9T9wzdPkhj3fqIESzh6r/LTN
NthimMkgKE3UzCuCWMdgpwoMmVqeO26qtgVMtjW2I3fjJqJYhWY8Ar4KrXAo2y1H
3s55USEIOLbXeJnB2R4JaY4M7qf/s+XxGfswoQLWkUCHOEmqG+I9rMgHb6rBNupY
17jMk6u1LQSqKz3I4WdyHJ3x7UIkeKsbGb2t9aExQEhmsjfokzVdN80lw9BLS+Nc
STstWT8K7xCbIuGV7IQKglEcdC//8MGndaVh4bSCwL+uyb6gp2W/d+GSE3jV+4wE
zY8Y9h/4KppbHFL0C98aRco2T9lLJb8p7uYdt95iKA6we/bsHDzXMREhqsW+LUCb
la3mMy5agm4LrbeZ6Gzt97nySxo8ZJYtj4swkB4e826NZq/ZA4lk0mBMrsVOWOhF
lm4V1IaTbHJszYww77rZ6Zn9W/GSGCZGD9w97AmJ4QXwDl8fd3sSoNGzSzPRK55D
ZAlTbUDu1LvvFcLQKE9BMEXOyYE3VQgnoBIBWQ34Dr0fBjVAN0C4eowq9SFcolBZ
z5e+PlAjD4AA6RW+7cDstrVNAd1m3JuqImailDWWajHNietTJsvt7C8g+MC0LwTD
4P4/ogUt26kGBx/B2dVGogkirMXtPJWdu0gtUfXfJFH6IYrejxM6AziZAQG2yu9v
5RBb//PbxIfK3utqur4lmJqP5GenaRX9oUaQ+Mkf949LMXD6thcjW+dR8AfON07a
RoKctBgBfxn7w71OfRPoejWXY95dFVe8P3ejD1uNxUFaCIUCyZayEQPLeZRqThRv
x0U2p0JPTAhevnhmMCe1PmOavhcfk8s56iDaWtgxizOujSfug/9kuhOshaHeGPui
tUZ/z8ts96Tb4eYPNocyA056YQ8B4+ytOAmObGVWC0uurReRoVETkrx/lb4kv6U+
ZWIKKRL7gEzJ1HXP81jyCApKSscKfhyy9aTxK8lOsq/Mg+ADofgRGKwB+k1KGeRy
M0KemONSY8cKsYs12BpLTPIMaJFrUIA3FKIMR8OwwBNJlMo1CL5RFQjW0TsHkKP/
YJvq5I/xuWpEcOaI4JSeXEGSBjIpggDqY9a5YpLUg6YTMGT1rfKN/A3sEQ0+0iaB
FHldot+K7drxcPQWpDV43dNnuBbsnDP1cLDz3CXguKMYfeLZqtghwedkLWtNu4Te
3tfIXQSb+N9K+M1WvKAH1n48TPXK66zL3mmrecjQGMsLbhV0tG0Ouz+gmZdqsVFh
2DkTV8GlfPNa+mGkhCVqWF7kB6fhGEVLFwAFQh7h/guOaS8xovMZ5k9Lqied6k2Y
B9CddyU5e2zIQYAZSLQxx0JCXZrKU2k57gAwCOBOf8H+K3tSFOV4UdzH+fVRvtQv
BHu1fxJj8pnQfitIOJYIyduJyziN+/1c4iVAEGpTLwfhYjzEuLlSdw7LxhWGd/sT
frLsuB3il0O9/MjJY0/AZTt+kkJ07g5uuTERNf+sQt6NYvoWQCsuVXLGaso07HME
6v4o1GamIKIJmytvwBnJLQhXxfTQZOm6FFNJEF1nbEx2I11H7Fc+//Dy3nd1BCIN
Mq41ExciyG6yUI4WAhnpCfj5ZPyKxMZWrNBed0qQmGfDpyorJ2atjZ4vmJwdCB3U
7J7Tf0s2u5jTvwH6WCOC5LWE2AqGSpuPSBP8CUqG040v9+M+6bqeZs2FLprC2I7l
l1UUl2feiYCPstWfgwRWU+HHm8yqjHg8ZO8s2zhSkANdrz9jesx1WSVye7a9uQ77
NZlOLNzb7kGJz53+RgecTTIqkGCiwmn345IpZgBDJZlZg5MRj0go+X1+eNUN1nL3
7Xn7S+0EQTLUpNjcVdPxe0pGVDAWAxcFx6OIQjYmdOMdEyb7oPFLWXq2ulifZQ5J
I6Z7nTt45QhasESPNci7ld1Mygh/4HsjDZcDJ2vMHiGZR98KON812/rZLugj4vG+
bHyaSKez0rNk1HpQUD9VXIZjQyGBG4ePFTPSqIoFprrE47s+hcWDPJfA8K6QlTJq
1l6dpQo2mmOl1kRiOSuMOljFyY8UW/F+jRd/SIGlwMUvkWI8rC0W80omm1NQg3Lr
9wYpeRi3mmd9ynl33xwPlIYwkihEL3ptoBst7c03pX18tbfOcf6h8lZ7KPMagDp5
EVkjfcJPRB2BGpC5ftbt7zG809q3YLKKWhxQ37D65bVzmHOsTJgIDdet43S3ewUC
WJGp1qqF4Pek3bhMnupfA3fO9mhqUXVjVeQRpQLLGskbkQtlvh8ds3wqGsJnRjbz
q6rM5Gj8huJnNqRGsDz6+x9roF9G/5nvpn4MLhBC5BqB9T36q6j4zOqMrwigs5jT
t9ijz921n6BirkbKcBpz/y/NIo2YaiAhO4/SMT9m6SSbtMzEUGvuoOtP2ELvmAtF
u/guiuL/TNA/X7HOU58BQFJRqoe64o1hJkRl5ZTtn8KTijbXfdrvnGG/iZ4fT4qU
Lb8OTgzvwiswEa5BtvhRHquj5Fdq/XB6K8JgKYv4trjU1noRxVi73LWv6QmIsR92
ReNFEfNkn7zJSJ7cLkgWpfiKuIVNiwkY+GdNqg8JwLEbtlpBK9gkZSiyYgY2gw2h
4IQYNUGKs41B8zLlzyG9IU9OYd3b79tiTN11tk8Bkr3URuzo/jfJ0Yu5SaN8axeg
S4uXconsxgNcLfUuBB2x5fr06hQinXYrSiA8zvvZnhvNxX5mtfX4NTsCcnS2jrb4
jggiSr5mN1NLISh/2m5mcPCE0kz6rhl61yoen8a+xpBkXut6rV6BRWD/qevOnrAf
63EY8JM6zujcS8Hw7MZPAkiLE6p7SNAbHz9stubMlMJK3BNYFlpBI+sbv0ORDp0V
e1TUYV2q6FXz58nYgKV1QMzwGZNczhluSoionfi49VAj6pfxMg+tJs6BgQFgODWr
4lHfuxnTJzPjSXBZsVVMQsGTmnt6bqL5yUXL3T1ppnBRDEqp1E7jZmF6wVps91rb
9/AfvBVVsf8FQBxX3gGsqxh2TmU7mEs9NQfwf124WLIWTzYqImQj1p7GQjkgAtcj
0+LZ0RX7kKfHhU+LNVrD1vmrlQVt5mcxD/1aopRkWPd9uNbogj71bKT/jlJ3YQIQ
1AosOUf/ub6vP4M99cQlSzaaXOIWqFmwXLqK/B0PXXody+I8F6tx5L501mbHlcLR
NV0dWkgim57CfeT1oenBTApK3pgDDVGXo3GmzjngVyWfXDs2qKMceTwJf6ZEniQH
TCXtkQVlHLw+1RvMlAezGixmfmSfdt4327udvLkf9aPm7YbXjuANWkkDo5JMc9n1
DSA8wcsH2D91dO1TXf+z8sNdYGtoAQeUaVv4wjYUEFIPY4ZKOrOLa6qQ54p5PyUz
6KAUvE+Mt2WYpQQdu5fmgIhYuevf0fvE+ah/ltL68SbYWG339rjGV+hRBd9cKc9S
GXuZgD68fCTFbhgl7eGfqkSsXfEriQuDq7C7XZ+8eU4AZYvzMt+ADWnKjSEU4X/s
YLMYFyzNu+0T356KAlVSldxrseIIbEq2B+Q4Bg12D2leZOdQfqrPkAUvdoimewty
Md7fsMFfOfc0mX2mm6AqaZd57/WNiGt6t5t1cLZRQVlJc+2KqCpA+335iYIxKMgz
HVagfi8MOCQUfxnx55ai+AIItII53F/hHAJoHUv90/ob9AJxHmamEdq1uco8ZhMS
dATqKJqSNqhe7H5It5IVOOSFw6UD0himDsJ1eeefWPvD4FY4UXZlIMVtdABjo06T
95BGN+/HjWitncT+3h7okSL62vMOrFXfCYe/4IHW79VJHjwFYbpz5uSjDXk0ThGi
wWUboHShn7+UR0wlG/GzaZ34Rlfq5TxflgJ01aZZqzZZFeO6ysXcpE8GDjk7dzgd
Ns2D0V6GV4pqLfL5TJ823r/BUGYW6AVMBMSEpB2zvkOCL+ZcaOpbS/00OYKxjTXk
Lp7EyREnNvmTweYJ1tJzTxXlfZm6/aVsgStOAAK59R2pmO8xE6TxgT5ENBgvwfxa
4bpmC2cfuKNn/DBUz4TwgKw3AtxqVG+M2JXc4CDvuhflNQDPYPzPSrxAFD57NU4C
TMDjlLaVvrPcxTVPCT3LvF0JTZ8i/kUB3k7ZWR18PeGUEvaC6FUrsNszm85kaVJZ
b1MadpV2qQWuVn79lAjLVownSQffPLrg0i1WzPLbixGcvRR4J38WAIDFzmhXlD0T
vxsXdqlgVsrKV9owIWeJ9XLvuWcBpqMPDSLQnVzW73VOiUW6ml5Mv04qJKHcKMOw
l+f5QbW0eAFCuCBt6wkzf4cWA0i3+rAoCQL+V2Lve9fEt/vavU0arIDbWtj9FRUk
KabWf/Jz3nBE1oJckCx+9OdSDfueDKqcmpXzQJZn4H+uMIhij3JYoQVsLSr/FhkF
lNPmyd0bpHteCyX6VkSWZC3D6TTHoGW92bpYSY+dmeRYTk1YwAmV5+RDZ9bMB5Dn
DleBZtU65KzrrM2lTYsvQ5V34ScZ+1sHvDCtTa0RXIX+JThpyZR4b7YRtcyLeQhH
GasLLBVz8E5fqYiv4DcNFhdh24mDtsA9wnssSU65Y86hEQP9fQZx6wKkZc7mdjBz
3ztl33tcK4xPvFrTNV7Jr6DWolRJZ04r7OnI+YKtfP6g+lD1amE+rzRqocII7o1X
culWDbR1lQ42R+jZVARf0cfs/ewMF1/EzkZm7Z2SJLp/XmhD5VXU3HZ92kGvSokR
E6FodB6DpzD6+Bb+D4wKLxUJBzEFW5ppwKZA1dIr/++gOMbq/2gjDABQHUk9ryU2
J4pIA0A/qlJquMux9H8t50m3p8g/tHEWuZ21VbQytUDjpYGzgTohUDNN0Z7y1gl3
awOUHugeMeU0m2kScCa3cssQwhc+zPIqfo/qLoz29yZRNr997djls5PPMUaToD65
yQ7vJ5fo6f2HSU0ELgCBchkIwQLmUpekgYOXKDPYdrxQ5rsHyFHkCL4r4uSaAlHD
zeZpU3x1sLRI9iQXfBNmx/kfQJawBIniXpCJLW37piLrGxu5NQyVVO3UMZdp4Rf7
I2EpAsu4P75FG6XnvEtVqk9R/sAumn3O+QeWn6Q3TBOW6aKaUwczRwwI6SNtPr7L
yfvsTCwGUY5S6iryfGXTRa3n/YoPl3+k0ko0/uJpGCt8QCMaDAYUWkPHCKxnxV7m
2m5go5VsYsoX+B9Hhjyp2ScZVABMyp+pY/IWhR+0bo+X/Y5bhAbfDvvRfRYZKnhd
17635Uzr0D45cP4Pn/Ivgif3P7+ODMVgs15WWkmlzXsosZVMCaduC0fDykKDYWdD
Qhaq/0RyphSfY7QOhsbiO8uH4WqkzTIVlr9NR7zN4LglPxZ7N7J0iTOfGTsxXAh8
p4y3zPmS+TqJaC9bza3KNLRb7piqsm/Y70FHmkpz3bUCK5VKbdgX5F7Fg4hO5cvp
IaYabvgZuxaezpF7OaSWaS+v+rDJKlABioawKpJ1zbnPKwSqgSkP42OdFRZCIQif
6DTMFEnvgDGfquHqnYY5gCZacE5A2FrINFQRjPaE7hGxVvIyILUeNLZ5a4MezTRp
lfab/JLdk0jNy9EfFiMR2L0LxWPcS1AHS9I4kMiRLkqVrsxlyTdAWSVs1w+m1Me1
bEO/vq2VmWGlu/qP3la6Bot8V1TSZpX0oXGzVYVAvXLotrcQxHKHfnkFifwUXBSW
YAT7doitc/aNuGkkcaELjAa/McszkgzrHhlU+zmc0JSw7HdIEk+lxecLkB/MTk3L
JmROxlr8S6VlTpm2vWNmI3gVIuPHykE0jbL1dQUpGCFfUBtwRBkVGzLZz6EbZrfD
D+tZ92NKR41Aj3YbrU6qqQAzk2fhC0iYlWvXwNvMM+CevCnpDjzpPQLEftNyOapM
4TdM8MABfwihnZ66rk1TpNPJCyTtIN+pVqjY3aMNKztU63LGycEYSWmjaHzxlzAu
ElAEJuAPhAMdosis9sfBA7QSOEZc+EdInq9KWn7yOx7FGIn7JbHsLDX0G/NeeQGl
6wg2OH598/a78qUsCKohXcMcp3JYId+lFHdmu+e383XrgH/vUfSIEZ8iORlndIkI
V6wrjXuiRpauxTNhO3yUvX+h6ArkHQW8zeZiuJiu8BWUT46f0TkS40INcShaCWhM
twUnCVxsCupOJ1Nica7zYe/jrH/Cf7+VbSHj1bcmESe8a2KAOL0YCpw8pyK0tca/
ck3ZNaa1afWc6f3O00RNAzMnievoyK3jsuXqHx1E12P4cHfKEB3OjinyJEFl37N4
p4hgY5/sh7XWAbE9LWdGWYzekt6B39560idqwLGis2y6RmAWLdm1V/SndEMdeMXL
S4RkOBlsLA/OKXY4qflwr1K4FpIoAuoFORAWqyPJnM8y6aymO99EWq6ao+h9JfJ4
yfGhHjIPMSWhViflCCe0OSlUBlUBEbBGnkt/qCh3u4fKbAxDxmwOf/a19oQsEx2B
h6TJmF+S0dAbbvS4SzaT5hqKsXX8ztHjrq4+qz8uMI+Rk9d0qNrJL3kmG9R9Zvl8
m4iOsDlvZ9EI3kGHGl2MGoQm2jRdpuJriT/mCCzDj/iWFEZ4cfDHo+SqmKZlh5ZA
/4izqmtlDJEt6/WIWiGZoB+jyf/IlRezBYMOZwopxyQHuZh5JBz5h2EfBJ3CJYBI
NEuWKkk5g9geJf9W/YRTTp1z+R5tm7zE/MLY2Zzd8KA3AYfBOQZRP3y92HrsGkBw
1RRVhyLaHAQuKDlFbZP7Cu5tuQQ0NUZUOEIRXlZAVgBw7v5qReyRMRs5SPftVbdw
WQN8/2XHwNBgXKGGZnx3pW4kexrHjkS0OqCDgBVzf7Oa2KjUxrEcFILPCnLOebqf
y7PNCG+5pLvZO2JGUNmtwMB2CHE2x58KnPJ8J6ILaRXIGYxIdWbtl1r8v2nuDqPU
Nfd34aI6ANmCDhvTvF1ETRWfDDWFck8pLIdhG0P3dBgNukzGM+c2Aqbw0fWb1qEv
hC94Sj3ovrMPEWxv+mUU/bmUe3hAIyYg35a7BapK7nSg5b5mVSuxLDIAHSIDSRmq
3WeQWojz64qHsOkHuY1YLlVkkkuFyQh7IGJt5yeyhKQ+vgrSz3VZ9RdSdjq8Lv15
3Y6IKDEBGzQR3ASF1zQqD2OrWokoCDjxhOZE2i+A1nLrHyWDjLzKmKw5eeKDLqj6
n2P/z4Tit/KGHmAdMk2n5Xh7S7ukjK6BGVHMVCZHXFc9Vrq7YB+AgnZpdlWPaz3N
ZqGeseMiD0p4tnams6FynbYmDrnzpYOyRMaCy36QBZ6+cLJgrWQ/nTVYlzzFYkjM
S2J/BKtFAguOi3rouLNJLnu1eWODA0Az/gd+kOz3PRuL3ldIRDMbozejnc79oaDD
YGJ1ETlWPjM6v7WWNrE6BZmhgQXkZk0W9/cPw8nyCMzrVNDVSRCmP8TLhtNdKA2B
RwIzsT7QlgoWJE5DYP5XRL756CUb5+/UieDqmP676TuOIbcsSFqiQbXaPp8MsCJ+
V+HiJakUojt34e+FcgDGf16vfQktfgEPc92pSj0DbeAqWqoUcPgxImtic4k8JecJ
wCleTcTihhQf/zjxF+BbFaWqyGQE/Ce99u7cHioYDvHsZYKszof1BHjcrEsc3Q/3
9t49PVYLw+Mhma4RkCsrHrpS6oD82lOrBRMYjA0gDn3arFUppP5YgRxkVnRSClNt
n2JL4WRFIpLIscQuyb1AkT8XQWopeASTD2pK9zwuMmdW7HhtRP3fJCWvAm0MjnYj
34MqfbksYLzqgPbxixjhlieigfP5xXb+RW0wpXjDPTWcDW/lMAPONMCYEygFaeS0
fly58tp7tOqJ+bJngGMdM9zXjyqDNyvSoJWQLxS+WWde7x1Ksak4WVU32Xi1k/vv
fLLG6qb29jkeS+nqhbHnAJYgfNrXs3N1P3z6tlCKmS9B8qBPOTnV80Uua/UbhLzE
6TSnzyN90Rv1b1O8N4ai+0vNgWuFDGvD/T3LCvfGugSfTOk4B4VqRJxSAONhHKmm
UdZYA+GI4nBwZNcqvxk9uQtb4SuJzEKrknA6RJs/jxIGWZM2g4sfnSQm1z1MX4u3
wNBQJ8NMwusB0YDnazgxC2F7o9kvlqELPJ+jPnT9xXaBXLCGMA8FZqAiNo2m7L4S
5CF+xGfkPxNvA5ltpGcmiS9shhNoZO7BFzEtSlI7riYg09cS8l9upNj3Zdd1Go4M
kRimxCtESKw+05slHAEDoUJVR0PNJoPEQjvs+6Pg/VlWlbdRrg/WFpEP/UfFmkWE
/8DF0i/3z9TtSqldHpjwZTdOR/q4Hxo+GP4Lozxa8DHqo7Fgmm0vhcBIoseOyhaj
XP/kOrCKH7dD+nk4WZe4+VF9x6qZMSHSaWy/i015Sq4lvA6mt4hXeuTzkeqJYs7I
DXWRnCAHm39TbxN3yIGHVVnfYo/6A1PaUPOrIOCqMD1Mm3YICyOsxi+EeGcD+S51
rTz0Rf4iNmRPFlu+ZPnRuCXFOTincIP0DamEQkUavqYd7khN8Soi48owll9qW7CD
e4lTjK5a/ypWMnAUkXq/iV6u51NvpnsnG3NKuAaYs/ZwcukXshDuzTBtq/MhNtLG
/SE1tadC0aYZ6JyRrxF3fz6OHGRDV3PaCkmQLiK2Gz7sNw/zB5+ADAZ30V1KfFer
AhWZ9axRv1IUKqHXPrvn2Xpb/drKTIFEWew3IRJTtz8Jram0YDRzMA6PP90XIVET
ACc43l50F2QxGE7BqK/QiLD9Z+I3XT7wepRCNVwbtFGqtNgCRtE59XBfXefPQb9b
4lovAlXj2Y+7ZFsH69ALRQbEY7QMZ0wrz5lNcc6CbvAo4nGXM4RvTBo6YTp/VLP0
kEhFbIW8TdBlcIaYnoLl0bAMVFwHPswPAQnqLiiVycJPRmG8CeXk/cxColjKdL6T
eUG5f7ZXq0GEo56uUxgCJ4m0aLjgD+8c2XGnkOwh9thId/tO73s4hX+GMlUQog/c
Lwd6T5M8rhMUuHNrJqRoYuSICZTMa/mKe6A0SDQ2L8rRZZXk4U3dhK9rw1JLlG3S
Jp3N/ofkBMneEpoG//vvWWI0cW6SBmGhju3ZyOd8EyvuwLBd4rl+ILsvSS9oL0tt
kjyCDRooYAdF9s5E1QkQfOl9IrYV3eEdC0Zx+LbYE5zeDl76LcqWsUkv+FHwiitv
0OHxB+Yji0FyAChZRoLOHU4+TOpcCxsPI5Zau6YRQDLlc2QkLpwme/YZtBDoircf
PjoMdyzuN7pQK8sSo5dQRZWjIIujuAEY9QGl88yDA4mdETO+xvC1xqQ1+qJ8OX6H
gkgEVJInbRPaEOpHZow4E4Ubi45/x75yv7HWmLyIqsAjsT+Ih3Qgt6NTDhsZ4EPz
xs0VfJwfgKVhycZWzVtWxoOrJfwJgJ42MoQhUebgdcwyMWz/spUIgTzp7Uz8gIr1
rTbnyvynRJ22q1VGm/iDRfiA7fbMCkdwYOR21Q5cE9q+Y/AwdsE60YgoO/SbD35m
QBmXK9Eao0tElT5MFcvepAypOWEZweixPVknHLbPqdnUgKys5n0+BOe8gg4W6UV+
18taCuiSle3c49bzI+4yMLmcaiBoh+Ata5ZWPaHV9B+UEMySMKqQlydd4am2qm+b
oxstFJ1abClEqVnWhffOMkTTdf0CCAL+clUegPpg4WQ21nmFuO7Nesq0ZjxVRc/V
NXAT3r82irDrt9yGlT0KhKC4eeqEbGJN9dkAaiGRfMotfA6mIo5TYrdLS10AisZZ
opnKmkWE8epenV69ThjKlAIGrgpJ2Iw+Qyk/GpoAMztNA0k0Glere5HIuqXvkDTk
oB7VPpQD/pVaEHjmnSTcKZarEg3GVTLwVXhWhlPzjKE1qVlk07ojq+2O6lF0eaPS
WOqK8ap1ajTbkIa1dc0l/B9nqq+TH5qkOe/6ZAO33JJz7ZXRthkNCOEbBU47e33f
R3eSnbEZ/56Mqu2twWakHUV4AQ3xm7DF/PNLdxOa7ELVCbchBShGsfOw35u2UXJ0
A0uREmJUn0Nn5pzl/P6+hrjvaCoBcvMpZlXpnLJQzsE2Wjw0adKzyz4+8Qlju/gQ
GZMIklg+n2XFBSNPYd+kQu3bJ3iVP8N4scjCd61BKvyMgdkf7XLvVRdtFLpmEdIo
kv8AtqTCx44cPuU0DhX8BycxueqL4QLAF4y/88Zrhm+1d4WqJJCjYlWXcKsv7Kyd
KJEtwSyIvwePLM592T4DSqXRuSkvhOlnF5Sprjwo9X4rj79ar5scyYI4fnGomNWh
YSHUlzgH60574YCHYoNcnIHahFPYgPv/gfSnVnIEZPDbuMTyDdjewvE7FpoEjgCX
LWzsHlmpEWR8GcJ7bdXsu9GTRHWF1ahJkmmNu9OKQV05c+U+3xN5nEziVGGdOMFn
NztEzM0fTOCCF9n0yMoBmyRgPDB+XbtwXk7izBTQcS9axzlAaAUN2a16bOCqQrc5
WdixxCwSvpbH3+YEaSbBFD7/+cZ0+fuoeYvHiW0SORx1yGZWpESH2GAWnuvVsjH4
+DGR3enfgk+wc40Yax6HXNfcY62HcrzYSFLLPAfpAv93O4mvNeAoJFsvhNzpISxb
5m1xwHu3UHTToDLKy8MrsXqY7Nmv4mx7BabP9LwWsLdvVH/k4vIh5LpDn0uny2kv
RJm+S6P0srA6AnP8eqE8GSSpx6GdHSYSTuCxsp96RLYYH7T07DOsLq6UAseIFvSP
opeIj1p6yRWj1uxuLkVUpS9c/tbbCcyAmA6veYS2SKsZTBaaw3r6zrlzhyzmSrk6
29BYbrKvyJP8keuY80zlb3dF0vsgsOd5ZFbnczKaQ8iIrW6MAWoSodGXnVtWMWF/
EV6ZUOSGP7x7oYKj/KrjHAMgQWaYAG6J24QAvUqcHZZupiwUYRWE1rfaNl2FAlct
KDZPBKK6q5ymJ75QPFGQFDn/R7/H3Ov6XOEQoqvHI7ZZnjMNCZ/0lBoPQB48AtqD
90DjhLCDCaiKa1wYHhLMfwx5ysVXXRBmVHaibl3A1TVMNay/cKfq7nCgQ0D+55Nv
wkBAft7Gv1BpB0PWi9HoDutU4hSeWOA4cjS9BAvKCjsKRYKgkHaX4y6KAHUnVfjb
4pEW+Rq0TZtX0CEhrIU+Fbj7JgDqJ+nrEd6pvw7/x9HRzbC0krDD765yaZaXOxXr
EHIBfLE/w04QdJUjDi5HxyQE0rBJyOSB1gRMMRNRo+CO7ukk+xdW/MCDprca8ghU
f7Kj6dSpzBMnMs08ba1LaOlefONu6UuQwPSRXguy5wpEtIh2UGWm2K93H+iHhVe2
ntMZWA0Y1+C4/n+x00qgcrSj07cFX5UM5CUP38nbrFEcFkxDxXvvyUsyOJzZX+w8
XTBdhVrJHje+vFZMDMUPqzwSSw7oPUOgJnh8QOt86uHnD9pNwAMm8VNlLZa/T/pS
5ztc0fqUBBeXPBWxbMAiFhN0HXGcMjlSe8DzwBFytS8pg9tpJ7uCYZKaThE5wrO4
cKXEvIoT3L4fTjTeg8wDIXsxmVxTOFOCGGXNpk+ktYa4eQ8DHfaeKf5UgAU/yfbR
gIKWWUC0PHLupNmru79qLAJ9RS6yeizj2k0EjfL3loCSky4eanqLg1JLosJGzPZk
y9IQPxieAw2FQsssMXIuO9y4tht7YWJ+Gi4ws+kCp+AB1OskE/AazwFUM0qDi1jF
vYuhX+9zpPo5YnJoh3c4pB11V2lu/aCIa049NesjdCidPLRSOdEVV8eenCwqXjKS
IaCEf3z7FiMGacGPnBF6pV0ja9Im8tsya52WYYTucIfXFyXpy+AltmGcDRejQyxE
Hx+s5opS8lJwkIbJxty/ibFbRMR7tRsmm2AGIRsBGSnNtUmxQvlsU9q+7y7rJbcq
e/VP9XcIERgLufUrMR5Uo9LuNbsG9Afwa/y12Jrv8ralFHXcAdO3lVT9uNs+yN/i
DEgBHchjs5T8QkvoiOQzkuTPMOiWQgp+MXaVe3QnwhJvG4v09Jz+h6rUC3uiCkGj
n0GHPJ9weXg+u0v/zIvYYzLfzSdY1E2FRlHNqphnD1hlkg7RwCbDYUvVliO4A/GU
FPNmxpjgq9v5xX8fGKqspUGAXIIF3A8q4PPjdtWQk1y3GHrNubNslNEDhl7oel22
pMoRX1tu9MyYZr3m1bPSdDsbQHJK6HhA6epN2gXOM9TKpI8G2RVG1sHxxNT/veKk
Absr1GYseI77/TePN2W8Hgz1flHPLUHUC6kQYKo++GGR+KeRtQRxtBAI5lX+WCp6
Ko8QyfTjKWkTPnYOvfwa52L88MQfPSMqF7G/KQIcWddffSNEq+Ck+OrwNYcg7ToJ
aQMPd2oEM4gNy/CzA6ICzfa+PJciOsXdbijjf1JynjbX7FYcELLvlS0GssOxVcDP
qSX5cfSV7oDU78d61tivZ+JNMDBrKo59USpY5Pkjlz53dKI12XazFkCRbUozllIh
yd+25Y3dWhlUt/2Qurv0xZhCDbSshqxQoRtgkVk1HXTtyqMQLgSVkBoTCED9fn8s
DQNlY0pmcq/i91rpmJsZWUPsTFrSv/RUgOMdSJVxKeqQS6eP3M4MnO5dfQwF2ik+
zNLgWaX3oM3Y071qgq4n9ZweJaWZFV2wsl+VyPtj060hcd7KcJXjmMM0JHWCWWgo
1O1iUNR8pbsFsJdYFrb1IBS82QXTXH7ozg7vYbTH9OORGo4w1eWbjj1Y72qs+ZLG
df+v//650WNYpfuRVn+CDl6t2SOWEX1TaUgjqTW/ggl6PJRsr15Bm46uyjxA0yA2
G+29vtaNKuVMlp79D0DWJSHOPoPUjVuM/tWMinKHlcc8qLihVrqBZ3CogRhkB8g+
DGv2c8an3itaak39p5bUSsf8bOrd4aGUjyNvp3sy1lE+douuCm7G96vYbEY4Q9DZ
mK+MjIKD72qUvpmoFkXpd5JQjoabe3hYioACwvNfOQDMK207ImgJ4jE0aWew7Pgd
rT2MvbGd54v4SRJes1MQoDVxQyY1VQbssvKH3irNWE8dmU2OMHWNFHee/eLDoT2J
6Cjy3j2SCmBcO6aiHO+1NtZpAFq/z7HZ+HgBD0DXiN67kZYqCKxN5yeh1EGzwK4F
c/B3tc5S0hta07WT+B9wJqjKH+r0KyqsDAygfT7DbJempKB6crutWJBHyM7dMlFl
RkIko1rnX6FVDKxoJ0K7xwkhZ1SPInoxBYzZinKQDFONXTNnBVvybL92BU+x6g5/
eO3nkofaxiaSMGf4pCW5PV8kmmW13MO3d+IZJr09bfVh7PVKeA6ofeRl85S+qwC3
S0tjyVayjz7CcPOlwbLckczLJ9fZqXjCud5gxiV2NxsTbYnRcaeodU4EiAq6LhuU
URxsR201f3esGMuQ45togLWg/5fkeRMyqeTQC69VLcUAKOI7iV6HB/xJTYPgiS3T
uWOGbzT6s58yK0qGppWp9lvCqXe1UqfWPsk7jQK2emjiRWhJefZHfBQ6ftogDDS0
WwLQJQFY8b4TxC9YNdxNjiAbTtcJyMwjsnt/gMlsQ5MmMZAJd3Bz7hcL7nT4aCwb
NI61XsUlXNoPAw7Fu/PMivNDuKp8lTKVlOL6r0NGYlJI8fDplv+2a4DsdVa6V7uq
VT4mwXKuuGNjQIeejbnBRO2++vC00p41IOwPAFbHvGAweJo9Q1Bf8vN0pR0OGbdC
oYf9bFH1DZJBYX0K/kNsREUPdeu+Kn1DGyLMA+B/tK9mR1y2/XmBo07j4dh8VAds
vRuJdxlCygOFr/JKk830IH60mXPW51NpU2vV2u7ybWv1giyh/P9vwTTt2AQc8rYM
hD0Vgct+tac++xa6VRTu53p/1Ubvs911PLFuGEIFq11aWmNlWTUlY355ln/w3/1i
z2B7H8K/IPsf7WFAYB0C51GEccqbHc0bWYweY5SAkkHCFvP4g5w85IluBohZyKEc
W++wZPX4cK6jZXRByGEkbNo8q6ohgSocUweM8Pf0RmtG1/R1cS1+iVgT8hsqIUTS
d8cfxHCTduLnrdw9wAttfURwFQ28l6/CCj4mIQ9IP6kd0uKEl3cEiLSYR3u0MQ1B
kkSmDH5r6h3MvMPXlTs4m0TlrdxB0JkqUAB2VTARdR0y4Y9J9uY3NZ7gs25SCvy9
TMT6kgxwiZ15h2qqR4mcUlYXyGJAzFMIbb4bTgVkMQmhFeQNoTwXY8UBgNrOoOCz
job4c62D0uefWFzHnUO08swBZm8ExRulkvmz++bKH/bPvS3Dlvy2yLIsPvI0FMMZ
zYS9xwATV9UPHOfuGNaGDzNg55SlwU07nTcD8I2qL9tre0oD1l0ZEX0naCxcvvaX
F39Fj7lq851GA/9rFQW2xNw3bV5TkF9UNDoz9RS94o8AmsW0IIZE7X2Hn4c6Xf+6
KyOt9yQ4x53oIbNpZH2E+3nlxyYP1ySR47kl+JMfmcpzfDvoXEKtYt0w58CLHvLs
8KMyWzulLEBoPJthjk9B2IcN6DU9AqNUF59mp1DxqoGU8ZJwwF4kc7bcCEilN367
S2HZISGnbEUEN2KIQTQUMA==
//pragma protect end_data_block
//pragma protect digest_block
14yq6El2JRpgXiO0YwcZjcDyAbI=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
9Z29vpDsg4KwBUnkQPKnHU1Z+FB2vbEaykA9vo9fNDBYCKHGn2IHaEBiNfSzDTtd
w4ydTQa/Pbw5kcr20KsVj0oWdr4GCNpNGw821zIZiFjuAuF4Zruv3vytJDrkapfu
53HJqaIOVCU7uW0ZBUnk7nJV0/6cFoqo7Qnmr7hfyEiHbAhG4GrpLA==
//pragma protect end_key_block
//pragma protect digest_block
D/UEvR1kNHWa4ce9assOMFmosRk=
//pragma protect end_digest_block
//pragma protect data_block
FE3SLps0fL8kKmBo/nmiD6nGCLG2nncHDbcpqyC4Dio36LAzqqChCLGLxxWR4sV1
b5CEC/qEsIHCILXDhmqA998mtF7D7dqa6iZ9EJ4w2dkNsHjCgSLtG50sSpoN7f7b
oT7L4/DtRaTW3N3Oj3lhdDfx9l9jwTL9NQPbEQNPz0gdy8eHvbPCEVhzOGi48/Aw
bFSQc0fZA8knMlmDhcjS6EJ18qC5d5Cw8UVTa2Wbxt7maB55sIYzl8P6EiVRktfo
ZvpBjBP7efMmCh5RaDX0fqajUo/H8Z5QLO2aSEtFmtPeN32IcqxDekuLnAXxY/5G
S7aaa2/+tQuZJjO0i3VUcyaqLMTKe5mXeGq81Pm7dEL9pRVJbeEHlt2ZJ1VjDlnw
E4sPfsxx3A9EwVe5tCMN13hBmskxt4jcfYKan1iJv18fc63/Ry5tfs6902ee7gcw
RBCcNxDmKSfbVMxass30+H/nFoi56cau+pE7TmdhyR+6GZYWM3dfxZ7DStLxMeJu
2/u4KQfM3dgr8CL8JibIOMMu3hb0oFbr61SetH4d07eGXtXJeWkS2aQPgPoPBE8V
8hQ3sxManKW/FAwxlcRx8IkHWF5icRSzMv9z0HPPv5JmAIa+xt4e28Kut7fjfYte
3yVdLAhEECREMNFC3fKhLGrnXbhPPaZ5OK7tbBeHCHv0OlroIJazA9RVCS2N0QdA
KqkSKEQwjREF7yz0K/398V93cy6/cnpwRWReUU5mW1KmPJuOKmiKjckaq41pru4E
Oy2wm5AEAATVtqD/6I7hR5JEaEVr1FsQ/C/xB55gAk7/86NFeQooF9SWJZwZvBzm
WmAIGzPzgjixxRR3YCK/9sEszx92s7BkSl+iVQtM+/VPCRwm6oXxZH1jR3VZgler
xGjYPIsC4NzlG1JR14arlCYuo/vuj1dQFBlYBAm4uuhh64S0dfbzV0+nn0BxZYbD
rH0nCUFDQpPPL51IQoD35aI3zHAsW4yJMigGXmK/3b5uRu/D/sryxwwqUm85K/FK

//pragma protect end_data_block
//pragma protect digest_block
BxxVTs/nH9RU84JF8u1H2aww3yA=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
F5Sl88yitou8WsX+S66TUckrRY4rvbM5btf8X7EtNonVwgpW7wycHGs9eBhKJ8G/
MfXg3LE3/OvH+KqCpA4ImqsB2SSAeBTyL7l2rTAXTzw1DspbTo5prFIprUrUA2yL
ULJYCCeiBXf6JOMlHZsGQO2SFyofFpAg1BRzNYqZzNiZn4koP7BsQQ==
//pragma protect end_key_block
//pragma protect digest_block
mRMRIJgwzSqSvjKwrOhdp6ukj1U=
//pragma protect end_digest_block
//pragma protect data_block
ZLxwOUKPguZyACZXDHs2K4y6p8mcbw/HFQpMUH8zimu6xCBbw8wn8/t/nQ5mIw4x
FzZjA/35gGkfiTPcFnCfyENGcCmRmkMPSXobRaY5liho7p5RTL0Mj7Uai/TCZclV
8BXwlIqyQRZD4yG0ZeJ+yRA3wkjZONpDvZJEtVU7Gv3SI5WWdzHxe5oiZmXgtW1Y
IaHNnVJ4qOXTSPeRH0BnzOxTftSUWrJ6LwPpD2GUlnMqDqz7Xy3yoeNdhasnlpWE
zo+4drDW+2LtEY+uhbOVrUL4LBq0crEHnHHApgNR/7UboMF1aOMXI5NJuB3a3Emo
edEJcErY8gXjEPLC57Ly/80TEyVBecJhObyAWfaJVQNSoE4jxMveXj+pzBar9SaW
ARHR+hkhOdhPO23a8b/6acklfYq3/uwGkBl0MJprzPW4RJxMuUeF7bsVO0Zxtz6V
b2K4sBEjzESqQ6Hkpzvb8QIr9whTDqSmpdL1zNcjaZORLxnomsYNjWULY/6g7GcL
juztbAh7cBLxZctCBG2LHIXXHgWj/ohzfeRlyo6ETLi+0c4WB2dQUvotG44D3Uau
/nE1yMZNKueF+x0Nn2dBSNb9xnCDAtqEjv9/dm/ViJLcMErSUmTgVgEyhneeOPOb
QVkucs8oMYxn3aVYLg2qWAMD5++YDX76neAW0EcVXA9+Cy3hBl31cZPPf9w0Af5C
FLeQLRohuL1vJdq9vt69pBDsQPl4SOmvsS7MfdMMeDEWPzR+L+CJURj0WpldIlCb
Fsx0xMgabW1kOb2g3XKV4ZFpD4jKOWre0REAL7p35xiY4yf5KnPGzCimI4wmqtJM
w7AOUMNzQLlCxBXEZCbSlsyy7uY508lcpTweu5IxyJPOl+B5QCEe5AVqRn/FW81/
ZMMdHV3tjKKp7uoXAgFwwTgHK+smn8bNHWeGmE/NwUoSyiKd047suZFh3T0Jhy1Z
x5bYsDI9rqp3tniJ4rj7yIs+xPaSVzEbeikDvAMUd7XF+FQ+t3kOjY0Qwtt1ppoA
JFU3JIJ4gh+Q6TxwMNQZ8bn0sZq8AFOZAamv2+WeaJgzjyBdeQ8E78X8WrGLaaFR
MU5SpkmWJuGbbnNQR2VxRIvPH6/QqKUhvpJEyH7Fe6Q0FcM5FLQnk1T9BQt2WWQy
NrwfHaF9afBPbyoH0BskePBx8fTx8fOmFXTqroEJ33s+v+h7xoU5NXnr01v61xWG
yvuupLwv0kIeP473JaenedJSxN8Gf5aje6yQTdG5RK9/24hWvw1ZAOjvylvzhbTm
3ne8hkUNJ9BFKmSeExKZagtGY2PcSxNTgwL0EHbOPsPT6AaPQospuPjNoUk83da9
1EaXdfG39ZRCFOM0KfU7JIcWySQZkwTfcmhHvdAhpOHD4qrlk4UqTgTItd/0ic1D
ZFJwcEIU3kNIzSfcFRHvg6re7y8yaDueHsN4Wk9VN6wHrP3sHfyAMOjiv1Cm3M0X
eUn40JanJdTJcr4hJkIhv1kN0rETKwLtRpoWVD/02zl+Nj3efOquYbmwo+oNcL/y
LeaKP13K9WT2oBslTIU0BFUWAewivlkQP+s1GMskpuDLzWiYcEPK9Xrdt9qYPUVC
KupWyxZE05jxtebzYZzJHC/ARjiDLb3zFhFPreoIlbPLrRUMe71AbQ77dWW3WsKk
AYIKsdLLukn9iyQYb1T/aM3THXepDpeRxFji4mX9VAjANi2VN/5l6uEa2DLsfNpR
fUIIb0zVMc8Na2nfu9CjVpzN7Hl8Iow/ltrG9AAms0+TPOQ502jdtRmfFPiofW3v
LQyt4ddx8QkE/QzELqU+HgX5tH9BFG+UXv5dhzPnu6xerBSttZ1JISCuQmRrL75U
7Y0sCaRi1z8XIm81yTGKNw1bVbKE3C404xjgG7u9x3zcHv+nLccu1wuwj/A1Abvo
VL1kKTaJsjQASY5vfxNoq3hOP7JB7wAtoAYConDb07bmB+XYIMTDo7baxuDe5IRZ
DhVxrx08lHPomDPuuCGUbrSYIPVjiF1+YOEo3Ck1ChDNqOU6DU0X/jyjcsDOFPjs
OKaq4yJxbVxgtmyH37KaE9BXsN3+USDCaE9yGW0vR4R8xs+po0L59pvH1Mn3LYwi
kJSKy7a/DRWwSWuU4tYEHmCWba3v2Jtf/44lWQEA9NWZ3j2fcIGjtja8dqPvaVfT
tW0bUc69+mWAoeEACc8QXy1f8+0d01xetZtc2w7Ji3phftI8AsP1TnzkcUwsvgJo
K0c9mnqh+FrWgxtCoFCWnaElY+68jyOKvknEibgCpYG41aaLc3qpeCHTbIe/sKm9
pj1bBc6WjnK+Ysdg1EXK5xcjunK6RWrnd5lbQ16vv+qzngUn+7hhQX+uPlWHgNTD
BTrbfxgfNcZvP3bRofyvjRZKxk8Ndw97DVFh+82QFiUsjYKW64b54wxJryHUzR4b
zozHWcjj419tgA34iMGeGhJEX7UcPI0iExYik8ekTvFWSDPUJs5AaytFOrytW8oV
r8StXaI+FSKzhy45iFE8BnFkIgz00gj/BLlbwT1cZg565aTLPVAFEDNtTPdLP8Tr
FlXhbWddT0gUa7EwNoTs3SVp2KuZhsEdhvExAI0TCJxROWyN3QZJOiPf3UYaTDjE
Vs634OX4eDCXQ9+v8gI8TwVzyFz9qxmePyIgKK+thiie/mwBS/qIi6oAJfJOnKEZ
fFYZXgcMrce9XCAkfNNXVEVZ/vTtDhjoRMWoUiysKJgb7tyHx0AUUQ5bNW9jSCdO
vgeMkgynpYL9WC2/zn8IZShLjIJD+ggMBUXank2SvEZ384Ug60cPR6FV8VWuGerh
nPuqfHWlDjeqBDz6XuvNM8Sv2rLkKNDf1NBRNr/vK06z+Twptu3FXFVkTbc8LgXj
BwzRDX1uLzD57hTV55A3tAVT6fDu79ByZ6VxCWrmwYDYx9huCSMVck4D6ztk+hZN
JUS9oz9g5C4P8uzJZUa2yid/cv07B/Mu9fKpv6sq+eAG0zbggbN5GzL5YH05Uyq4
CvX/5GkJDy9UNs+OUD7IUaiJ+ZOweQBIysm7cTmcK3EgXENjssf4apfKnYW2uncS
7cjRdgWx1upwgPCN/YMpQZ7aiTGW3J29UlSLTLci5yuRyCGcQwMWQjdWIujJEAly
I8skGVwoZCB0EIyJa8mHCbuu5uBvk1T7GenEvjaMeiD3sgOPlJEJCGTXR0M6re4u
YCTpai9qP7nHXiWVMe8Tjrtg6WzKrGb0aPHEDRHZCChbFO/zAen0nP1muSviXYDb
xSMKSlfWNdMfoUNNdBZ8tIxwx3rrgLrR0IeL0+EmDLc0e1M8tyU2yiZ7NQT3TQsR
HUqfCORQOM3Agm6fbIWeguYCBSJBKjdnkrO3qJ1zuhR6BFJV4FJ6+qGgP7Nuo5Hd
KImMHGr58FmtFetzq0/AEH5XsTDmPenChP+4u3vvwi4AyvvvSSrxa9OSAcrxMiHw
u5QK+M0Q5+WrnX26U9n7PC1yRwfmZcxVDGZ2DJGfKvgHgWZa/HQ1lJpPcJhYquTx
F0qAQsXRm8CM8dSSJ9g9lWoHrOyO0X47DV+Z8hgJ/4Eat+vCssQ57SMJkaVbse3p
K/jS9116Eg5g9vjxXzrBIIQd/HKOccjNqPJ5gBrhz/3S3d3tCkSkt9GR6o8HAUBQ
hkk0MPf28Cfll/J5t34yOLyvAH8etekXf65QeicdUqOE7TTWT8G3xG1TuBaG8gFI
D4ep8nHNb3xSDDXfQiWs1VjYnx5DXFfLmPPTQnDkxmNAVF0n3Gu6lGkDg00m9j2C
IZ7KoM2jWvH8lisovJoVdqLCf96b9pfwlc+yikZlPusBrGAvSpp+9p68iaGD7MFm
I2M91qUy6FKLd9q+bmsEco4fltP3yqMBr3riYCIpPhXJfzbhFKQmySLET9SjRneb
zvbuif+BM5eP59HgV3LCGRTfiAhE51htg+tIxarMUPXuDghnk4dwevCTp3RGzAfm
mWVCHw4jGF0SOg9yAXBfOY0RLdM2hue+Hcz9lTlwnYlIF5SjImAgy3xARgbbBpXh
EvWuNH14Dv4J0HpD6R8r6Rh43f4qIj68uosUxyTigQIxo0xorB+p4GhthD8NUUOq
uY9bO//qF6tZ64bwg5FILCANmkN+OQRfavng22FWJdSnr2++45o5P5U94B2K51TP
s4loNJURudiKOtopHBsXg3QcypDzYMLIa7egrQ9WqzOTtgjVnqN48/gZv7Gi28me
wLobuJD3J+iTH/iyOwiredpkrYKXzkYPpif49ecfhAZZeR1plthfzSmRKhJdUz8N
iP6SDtdDUCmpN2+Ltkk4HpvNHr78ge38Mop2YDUoeArTY/iAZsadRRkgnhdvgqFq
lE3SJpAMVDABECrp53ReiaDjIw+UmRZzfNUigfT9UwhY4mTsL1c2MYeJ/KsT25x9
jgLhwoamV7xscF2uotx2sIYIL8RaQgTL9g2app7TyqBe4QVEEdQ+xKuxcz3BOyHH
GUUJ8A3SpEHUm4Q11HXxZmRtf79vwKZgdK1FfPU6+2YQkIeQJjfBL7ilnSaEl035
yBfWJSEgLC9wupCLHAJwCBcWEH4IclGUamvFSQNPDz0WPGa9jAAH0vfwNW3m9ZPi
NXYk17WrTIByIHD55kwfX4UaFHLGkrDTgdfJb/4/QZYjoD73269lHYWI7LpRAYn6
h+LJDNDufTgzp3rZVao07k947hcFycMw5zeUARWyI/pVCNUvbaf07MBOymty4Re/
YpFmfgcapwoAEZ9owrVybH2vumkjn4ugb6SnCknBBhgjJN3SmZCWKaPo4LdK6S2Q
U9qIHXjP1EcI4cva79Z0MbThWvfGvfS4pWl1ObPhgy7LNCU92RSlyDwPtCK6ssL8
l4cdWn8tghU6THonT1cesC7bakpv6e0WLVrm/Tox12UbYl4TZTtAE+qiGNmV3PG7
Wvn7Z/m7f74TCQvGGEN+k/03hM4or8v2apQR1xQO6cHuuhQPUR5VbvwNY09EkHoY
U5XSe3bxqFtMX2uN8AyuMyGdfxkfidlEQlVPrzOMmya1nxStozhcHov2Ox9GnNtH
/CQ37FKEtLLJ64Tg8QMIdwqLog/7AIjgBWZAS+m8bqCXV2k5FaxaTWLeO08778PX
fqsFPLobM+tLQ6WsddAM8WeEp9PvhgJMp+BSnEbRapTk6kx8w5hE2zfDNT4joUt2
gAv4DyMd8atYN44Be/I21oxI2eF2gVGbea5QQ+moVIDIpqeHtpdu1ZdS4fI7Zf9q
EXXdDD5QkuDIEHSM3wiPTzPnRaA65WxKeDLRkY13RecWV/lzHtJgZrVUoYGPYX1f
z51PbxjmWkvOmPpgeKjzEtZEAam+Vj34r9fLzUpm3RDBWV4BAh6fXR7AsHC2Pa08
SN3UGsTZaz7AtcQ9I6YausF+BSdTNTGaeovImFjwR4CnAZX+x+lNo1GESzkrBbdd
YGQLhJgZYQnrK1MI+LjSdDOTN83nQFZBFbfy6NGCQN1zzUX23qtFLHkizMfIvYE0
kvXFw42udUVugf5jtKI2k5wMcXtkB/KRCreSrA4msVJrMIicZVawsNOsfYS5v/19
chql8UZ44KzIaUgbLZqneiKP/1HP9RbuqxyVfaI2B6YbqW61dKHjQ74Gjmib5CgX
A6PmT/frnpaFskkTsL0xKjh2/YX/pJtavbrqdF1ghib0NgnPs+vI+eV3tWB5dozr
yMSu7gvDfk9trXCbBvY/gVfbak/4sdg/DakeDWOXQ3qmX4jmnHOGbKfbAr7VKO4/
qk8Cv6Rwrscrd/VgP1TmZ/9cygLzx8Xb4T6wo7J88AxwZ7XMkFsfGHEweQaTm4pf
txFQySK5TVMJUsp/KjXJB+K/sui2qr6PGJm4QSZAJ/635Sqtj7VMZXTiY4+KkfNA
4Znxe89/k9M6Yl5DsdtS/0en7QzA0lOWiht535rU0OyFVBPEjthTfmfawIN8k8o9
8NOYMqtuKD94/VqKjVGdAnHEo6dAjRde+20hkqQ1DudQ5+Ven1xpPL75nhwTossg
AqBit4z90VuyFvkzJAZM9ovd3XfxtgqZgEo54GbboOgMRJELWUjh1q3+HeDXr1Sz
vQr/pqlsU/fcBZ/75QxpKS8NM7s/8atIvwW1AatEh0CoCAtNjiO1N2r9fI4aRy56
in3OVNOiLQnRkxy4ryG4rZK6ho7kDqGHNh1ZOjt4wRminkledtr6ZC3cNmuK63Se
qod+Lgqq1p8mtWELn0ZYnhGfrmP/Fn1QmmFWuYSvxwXXil3ScndnvSGN803ySIab
TV3t63F6/tB+WHKo2oaN7OVEhFsjKXSbpPzQxMbHkLBv8NzgobTkERDw+q+h+2FD
W2rxIyElYVAh5iVEsegBw31N7gxzwJ178D2rvkFetrB/On5eyF83ALFpEfpF3Zsa
SHgFk1LfhFgjoosGeqUnD1b1SzYravS8Qq+b3YtNwEohDDCkFaCbz1xnyvBfiPXE
/RWVPtk/+XwgS2eigR1LVw737CbFvd5Y6vMM4HQY5ZrvMNmhBFTDV4eMYdbBudFp
S7IoH2OQpnEVZnUYNQMnIBEgD/ebBQ66Jg4IcuLd7e5njM99AwDHSBz65V/zPzut
IRYzvlzgm7qIBMT5x/kuHRFtpmdDr6b2PuFGlAryv/1lHaNhQfowyildrcg/hoNc
nExfbNSkZLtrCjLAsORgENEvnPdOd2K/Sm25mCq643lGXvFVVop77sxpin87TK32
WvdeLzvwpx0rhRbdKYFZMGRupM6wWQsJMmLpXREjzlNYDgBaFnq+GpdnyXGFmcte
3m4tlxZGFMvihfaeHkZftzCZTqNqVbnH6zhkEfeoDT0enEBxel5rukSTaQI6B58O
bKKyYO4ymVsE/VBQXjyFaS1G5GHIiVXxPIiWsffvSELszE25RveMC9U24h00D3so
N9SM8oRMowtg+QgcqR0hffcdSNGhICf3pQmpoy6xnirh592vT0mu/83EIEDpHqYc
AqhuIABevuMWnhccWH29OS6v9iiMQrnQ+KCufOvw5e9vhx2Z1ozdqMEV/VE7hAzF
yAylYaUcTJEMWUklewiLCHYoPMzwqv9q9FdCFIsUDL7Bgg+6UsFOV8RSuG2reIf7
zL7hUjrAj1ba2O+AQPc/Fj2935csAbmCtzfXxV+tV0fzssxDI3fG+M6EkMpGt4YB
7Chb9LyOXcoqilN51fg5SZi0GXSfVYhnQnnmgdwyMOJ0q7Se78IJ4Abp9bTqKKEO
agv3RUbqxLRROKBlTDng1sfZAOg5EwNaQVaT0mbxJDF0q7FuC5ho0/mWM+WOwzO5
RLRVBT2eW4s+WovihIEzhQ3H2AzISnSnYOVq0ZYGXQ6T6Wa+0FQYorGE+OppCVDU
s7PSxamhcEaJxseY5Z+DZQf6ppQJz3RaJTt2f0eUYF6p23DLr/danA+OxLw8puDf
ma9W2pqcxA9iEllx0WmbmbhWHxvX/CZwn2J5Q9uoRnYAbSrKOpNmzoye9+ML8fr2
vLL1YKVvWSFC/bzxfYcLS1YJyhAWuyZFAa1jvrderzNRsz79iIUo4xQ9avkSijWn
BRB2UqLR/qlqn4+Ly7Ky0XpnTX5WyCGXAUKFZ+snVjNRAGgr5YqQV8qbBKkfO6uX
QCUTf7JkfUj117U3i9NbgEvg3gSEYIYlnGJcF5m3EZjnUyQOw0TPG08Vw/krrUzT
Tmpq2cvPAcNwCFKJT4IjAo1xg71gU9ezZvRtAVBu7wm+ti0EuCjidecjOmJm+/4i
0Igyam9GSq9T+eCmog6SMOSMXhw9MIA4vU0/lBWgGK/EDfSLGHbaEEuS9o5FOr+p
slMZ+A7JrN7K7zY4hjKMjiK3q4tbq6b3s8p/tIlimrb1v+NTRwX6b7enu8iNU5tx
j+0gRNxhuFA8G012S+kBTfuDh7aUg16Wb22BRisl18G+HGidgtbth1hQ3k/NO59d
KHMF4gLFsLtqEwCNd47OPqGhJ/MfiU7GTnbqWYPhGdQpaHvTv3Xq7PGKjoVjWF/s
D9sYDjH3p/TSNudpD5bVVBRvRenreXtlwKUSTRG/Gz+MfxvDK6o9vwRefF7Rcqjj
x9vWmVqj/Msm0vijzxc3dSBzxDGbG3+PlekS9uAyrmFG65+H/MjGWhweB1vyCxHD
mcSNefmOTimMhksYFy0bCwwKUzWa8080fTEsB+8bG4OAOKr11HwEpoV9OFBAcWLV
UkXdjgSoP3BR15yrNGsl2+otD4XMsbfipn3jGZPm48/la87yvwMo242syJwUKAqu
4zDflc7kcQEo3Js+eo0fAP21FkxA1iUMTmjWBfns0SVZZ/Xkwghk39dM60Gva2J+
dB5PPnO47Ln79NKFUG0cJilm2ILvB/xURFDzSz8a3VfjPo0jFxAcgSQLDW46yMuP
QS5h0cUueHmOHmSmP8Fn9JMYpGrPfR9deKrGPuTsQPMFjRa4MMjWnZvanSLd98Qv
YOa1BbH5eu1HELBz7POw/KWmXMbekMOEaJeIvduA+ccLdmRaaPdk8oYZYdBDthh1
Px0wW7AqrQ6r0r2LxrchLY1j2ywU6mFR9Um8T44hdo4/XF/DzKZhWQIEHMZqnog/
Etl3debHYFsOi5VFyeAqe4Ck5nArwbbD/Y3Pww2v7R8uOnHyaO6uOlbrGl+jMSc0
V6tY/oih55O8tlEljUXEy03lSxppvHINvXm4BCdu74DDJrzjleLD8eawo9scWaxj
UU6eq/gl5mmDMc2kuIb0TpxZy+p8jTMfUfAlQd6W2z9b2LDYjJf7DD+IA93NMP73
YTTyGhWLhMUI0ZuBwJ//IFowmE0Srkmfj6Ss6dcTrawmf2vhAs6fsRDSJ9jxfprw
4FA0corYhxxD06jit/0B9eqqN4wzvaVGaT1/Dp4QB78yX9JODJl9NjoZll3EY4jO
Xc1CQa/UjqDuUE2yNErBt+UETFOGGwd4L4WRMwbw6H7VeH/NXZxT2HOFtObk902R
BvV4Z17MSmK25YO9ck+qaBsQqjCr9OzygpzuS+nIDOvNXsQf0FA0kzqLFwSM6Ii9
RjRn9RF6G5KDw64UljMvT83nU3NfdtkZ1opqmyGTjzAsoE8tAOrtEaqcd6tXo4ng
eMALXGvOP+HbzApGtEWMLAvLRENWOXF4pu9s80Gc6TrR1uNgZCGRMXAX1UF+lsd1
OIpTYtgQ4DWN+aK0N7QcbR6Px2J/QBl1HRPdG9DT3crMpUwAxypq6113E/zTUVQu
jB2us3ktgtBimiLW1xS4zAI2BiBXSfa3Oa0H2HEn0OJ3NTHH5atgNqsX+GsMZepq
cwAROV3hUG+kyNkaGtw+KpUiSkeq6rz0YFFa4WN3603rRlonDBtSYCqxIjUMZZf5
vyrVqiCvf8p4q8YEHDfmpa/RRIrMn6sza9GjKPMPVmdpXaQ3ljqUQkG6ejqdfVFj
UI/E47/dBkv3RHDwL0dGI8i+xxfrGzjFvDUpbyymrZUK177i/I6gc9HvPiZIaF3X
RYGoM86fDHalKnE3BqIvem4UQ+7KB+VOcVcNnEj9LpZZ1PeiaMcKvNXy9qFNeQur
JwrYosrcfL1VMg3XAaefdUqemDZ9MkF6BJH9DwixBJA8LzWB3CtzwcwzOQGweXaZ
vJUyF317wMQ5dfgJJ2MjlkyNXjGUAY3q12/a3XhSPN4rGUtmGePcPZ0hZb7AC4m6
kMpjyJ+oIlyMR6ii2ykmnlZOmWFGtm4YzNCUqvFqeOrafABUEuHCgqZFCLCjm4L2
ygsXMj0/u3mu/nEnBXqkp4rMZlK1xzDtnCLXNKFtFNt3u7WFagWOSmr4cgPmSU2i
c611ptD2uCBBLeb7o0jGokTF3xOEt+Ikl8yX+TTZXvHHTiYHrX+8cyMv8CWvRMX1
1EvkHbejxATGPyiH7UX0vElSQJizHM6LryRrUEpXLqpcH1ecFW/8lR7X66b9M5it
TGOdhEroVeX9WIM0MGBapCflhHcA9PV40WIEcKL5ml+V66VqGwqGgvIAwZe2W9bW
teHa5ILUXQfqsVb+mQfwyS9SpObdfiDlsGm4Ed6fbykwpAw5AdXRSazJHHwx4HP1
LTTXJBPtu11MTVjVqtHP3/d8PAT87zJ4HJW1Glj9JkMhRepOGXz1/qX5qvkCf7Et
WonscV/UmlECVuzyA7LV3fMxEIpVg4lgYDtTeUQJfHLVvDr+XAD43M2r3yK5Z+cj
wBrcWDo/VdbkuPB4kwVxkTYKhj1MudeFVABKPmxVIWP3dqLSuuKqnAgnY8ngxcgz
uqEMAvXadnAbm+tUmTSaHvSDysAITc4RTcDQyl6WTmpFHueIpD58/5/yzDGBDWYJ
F/ib7sD4yPjuCibKbvdgElMGH9M7e9IMimmRx0Kbs277hr6oslJuWRlZ0DYzQIWA
21w0CdeUnzA/tvsGub4Uu6EMVyjE/mx6kM3mw4rXfLQX2noGkr4vqhLUkfpUyrFM
NvShE+fcgshgeCF32qkhf8P96ePfOa3wYrmYa4dItxI3phpYVEWxp51lJdeQCYib
MARQfKPdzPj0Or3m3ygyTfbBxuXNL70SVrvsQpvbd6U1jaKjLoSMzV6p+qTO57Ep
piN4kB98DvEqBR1Q0pLgq5I/OXGJ4zNctVb5fzJp2QV9aUvkLn5gJSE+f3CCvrKy
YoQmgUmwMpvAVH8v0hQVDsiW2z4/LTfL/Kw1n7hehAreQphX97Yfi+nyLGtJssrq
LxqZ+DJHE9VifY2VvOFYhBAT6p7loUuz/p5c12uDkCkMFiEwipC+tKteHUlbmJQQ
awUu9wvl17b+yYWivG20RByB1P21e94UZHhSByFNs3piRzFQKyaWKjn3jHfwrnSt
t0hmWqBEYwVVSYRktFgFzoSIbq5fW4dYvJKnMc+RZ6DeBhWBzfaEDJ/9nQj0zRQl
zyM8JZSruc4nxQPQMEQ/JIx2BFkEiVx7UGODPYK4HGS4re2CS5h19Se+h8VzEcXs
PzZm8d19rs3y19nHPzJZIHUBa9JrgL5JyM8VlzMP9L5catn05ocn3pGgstou6tQr
w/PU42m9JIojVfk4SyUPsCbE4wvotTw4o0MefWb26IhtbGpphrwlM6zicdRGHkEN
d9Nh8HpINEDoGa30PnuORf/pmsF51puTkKWw2dAi6K3YquySzda46MGirPDy5SbV
5ixw/RAkEi03AgfLkyGoVel8pMicmRBC4MJImKIdsLE946/F//PLkioKNs9v0DGd
hsgICHrjjvBE5jHf86AG3iaiPc08Yxn/z+q/HhxSej7VIrL20C2XiFItbTAmNmzh
hEF0BmQ+A+RPFeimLyKiUQdtIicPwYYaHfHbWLYHo306JtF4LP8hr5QmRUyULw9e
HugFYr/50Bl14ALqUtfmDloTKcTESFOWWq37WDa3zpfS2kWsZTfHBxn4y0Rvg6z+
dHFjfGsMUa4SqVUnDPJVuo+NFskAgqLifgHVgJJPZ/JVfwj5VjFwC9tTxHQtjQnu
14pf4h4P5hePi1oGOhlzpV3r6nbPyKwSFSFi5amZcL6jBZfZaM0lmLKeYomWeF4S
0FP3mot9UP2Bo72jzLzN59NK6EIOPsipVrflPmnaS7/fFsAZ9GUN4L2MViklTP0b
n7NX0Khx0lNXxctg2on5FvYYvCWba1qkuVwF9AirV18FaPe//UjWtwdEavdkL44N
l88pk6RjPfaGnR7+WizeYO+HFm/PcqLH3gA7yTMldSWCkQYbve7DGhTnGVkJudat
SxoP59ANYVt3dlwp3zXIU5gzko+Hi35zdSNVGFzAIgC7+cA3/U18K7XA732U66Al
+AoYVQCp9APuC9MW9LAZO2EXZ0GOMYMvbuMRBvcoa5tuD0XO67Zhdwn89AA/YP2c
qycGg5eaflxa4qkVVtKMEGIz1bOjRqlpEFeIn2H+6pIjmgPq0jcrkS3bTpInYulP
am0muiGt9il+EpQKnzkC5iDCeQEZP5N3H0F0cqD/pIVqMp6a8e0FlBkcov/XUJtT
91LazooAGJ9Suju/CkgVd+rM+eyNpKMuKqJtavmhwbeLQl8UQf7KMxf5dO6m0bVX
aaAtQi9HeYs4fhSym+UdzzJ3stqds6/GhSNxlPSOEKeXOrJC+z1AUkfacD1qnY6Z
LlhRxKFVXrTNTobGO2lL4JVQZyWEJWqosZHz5GoEvZxG+qV/zjQrJM2bWVtevlIc
r0VHApB2DQKwmpggSNL8KA3S5Q9xUC02lL1LjgZAA/x+VOxPoG56kxhXauVBl9IL
34R2arvOZBggReXGOJ+La2NlfCRmqc4B6zp7QSzkMtxJ6zQjyQsSdd1/EpfViofi
1A4hcKRWbMpv+OjZ8UwbX1WYStZHXO4ffbf+n2zv5tCHt+KtMRYHe5xSEcJuTwjn
eA7CPQ6kKFBX2jq/UaqkysKpotk+hJQKTRQQbCjvPN3DG6VTwxoUtfJTTGTUD/xW
IM3ZEY8BPd/LRuY0vKtKiB0ZadYcW/fGH0kTNpJpUijCeyi8T7h+NpMaaov8D0hX
4Pqb1MHA2FrsLlIU2J5OZIve3rOhfIht7Mz7ZIQq262WrFwkLpP7U4cmWAyUuba/
SrFtWuDtBYH0ogIbYIaWi7TVwVV21lOKSUrvIDHlmOpQJ72KczQXXoVLgMCOgzAJ
ELHsBcmwjLj2AfCeNvyLHLcACYfeX66GcJXIoH2HP8YpmC0FwIs7b3pS2t+BbQps
S2dfrFqnp/CAmbkfrHXm2kWvWjlQUgEesMbbtSIz5716ab0pStXrYax/lrQ266Uc
awrz2FnxS6JL0M5oSlAhkVhs8JtoiKiBS7c3OmUI9gWQUjXJUScelWRNZjzjqdXb
7lt1u/8beFP6Ad8YpAUqj83m0617rwM4dMsq2bSDi+eUMh1Bh1rgYIn7BlpCA580
OMrOtXBBP0HHtyF+m0iBDVVh4DN7TWUU/fHVrmpoOd9E5lO9bWJlVZovgeuvgHIa
ZEKyVqmwaPHtWKFgdizEIlBiWXjcOLYGNjsvxXly8BySUWZ9cTx4ghvKcTn+m9xZ
qQ82NEk2/JnTij5dDCoX6laEAKpC1YYr5FeZHvJuv+7+X74Gvno3ywLtkgKRvDrA
8/QcW8wtQhTQ1GBtXejCxjC0Bux2LRu4jgEjgQuvVknxKoDDPVfRi2hktGe5qKxz
a7EJvZr6GA+jCd2P6x7abnCeFQrsSj4e3Quux9znOsctDaYIKAVB+b8iAaYrgvI0
VspsJJgXBocwUGOxX9ClCJGlSsVQ/iLTdUux3zAsX+XchuyxHYRS76ouJHCYvvyD
9JqEgqcXz//LzBsCBtsYw88Kk2X53qhAbWjLoTKM6yRoslzKGl8WFp+7QimSgxqt
yggjWn6kSB7T6f45jRlVK5ez3DTyAeOpUGmK9exOQUUjrlH4dS6hokAWzJURmFst
hEA2g7/cxExFRnmbJ1Qj4kdY7TeaadiwrssF7cI7Ya6Jsa53KByJc8HgiDvGzKDJ
F47pkhmqvgA15Xe0DTVGj4I5jwgdKWBIRzNlA7JIqPfAeKof6s33zbRynZpePUE7
ZMdtUH7f1lZ5PKjci9VroQKM46p7Ir9Tgd0+i3PGiok1aHijoPSB38mJgA6sL0v/
q67ljoIMAVS4nwQsu/KgEYapCQiBmFvG4/1OQZjzjQHvGW0ZBYi9/MYc129Arl8j
yxMGHQBtKadtM+DIDFMG/RXG3gZUJVL8A5mcqsCEYbHyIU+kE8Yq/xYSnFs6Paik
LIxhbLpPJnzXWyiyouWsLxaBENgU/8LIkJ3RUr1SkTwAvZjl7GCBUbisRpb/dw4G
GNEcArU0hTmYpY89bRUTygEIygcTvdBu7izsQRKO6CDXqMOoJZcA16mx3YHenzWS
X1FAcqrmlAg1vTwjhkk4HqKa2ZbUZqEFaxC2ZjFBk+AP55lZ0XS4Iv3PqkxhthdJ
9MAaggvvESqIhE08ywuXug4ljPNNmmO/7+n0/wnVUnVSH4+LdcM7oLHvVLE1NrW0
I+8LnY/KgS6yH/UjPrltYxQ7p7iBkTE5hE0zMt0myWYnCcyNjn4TKDICgWqWzlrM
J2fnSjBO/hmRSOQWTwm7QpaRul3VVMEo5fKACCP5eiY863Fo95G3lFCJTCxsjNpd
DSaRHz7FQ1P8hXiRWEp4H8qb1OGXKW2FsLA2UQ7bWejQ306B2cz9bHduSBqRpzDs
xWKMigl8vfgctL/QpV1r2d/f+Z0B/4Te66bnvlHlBpm6GKjspMZWkCr96Alg07d9
+5QNto+hJZLcC14Ew9BsTJh72kvnajzgajzaweUaRnKhJuCQRk05e4SnKLMQLcJK
TGgp1asnc6/G73N7OCV8s6aSSySMAQBfguZtcdY/ImuNLD33SEyCRCeZyblYDRQQ
KBjtVr2zGy9PN6GfaRr3+YRjBqOkNy5ZH/GBFZdeurZTqgNiRZDGCUmDLLNcWGrc
YPj5AY8AEs+5mzkQ5eWlOYxdtoGtO/J5ZuAFgBJhvhsl3/5soBu7OTB2t+k9lhZK
a/PhqwI42/jnVvc8vBF9t6MSKu384hjqWbJaX6U8WMti+noHcCVpfYGsbiJizv4X
lQfh45bStVpGduwXpTmoQs0MvgpG+QT32ELuZPDEdhPX4G90DUf5Z1/PtY4n8nl3
5rViZ/GcvQ+h+wW/k6JRuzfr/Ud3ln2/VyhqYZaGKTrpnw+UXwx8vqyC7Iv6EYZD
6zKVdfr9KKG7tK4W3HUItF/sEfov+oxrOhiejuNu6V67tSWsv4/jaKyr54OgMkky
G8ddmdmV80UvXzohszsKOLeQd9vjQXMDVp15tcpt1s1EooW60HHm0JGxVp6ZvMMo
LuB84dqIPEG3qKGnCpxDob3oq9XulODi6ka7l3WZXMLXL7cN9zcgCi+hH1X2ayab
hTdeUbLqQITjzxq2hfuUZTyrMkq3QqKdvGpObhJL1LJKshIy9iW2tAJnXMSQ8VLq
vSihpasi/4a7LQZsTQdLSfQvRmNAnd1kCt5tvTSzRvEQuoPRwAFoVJ/5aZGZ64BY
OWYZyO9wqmK5yuxyIXRM5hVLGzBb7B4SxASzoLwkMJ6vq8hXuPXuBQLKdaV0/l30
dsjF9ztjx+BO4CPqYQ+CUoajw6oTKI8vd1v/rRy8sWNHVuqxyFuH6YsvDvE96LwF
EpYDJaPwyTjoHXq+7TBqiLFSByUyOZeUMUS/A3QXZBlOzTd88HjoVZXEbhVmzz+z
RLzFxt/JQaHdz0feY4ZwWKjnW4nJsAV3O1kEZgrgjVfP1dYb2lLP6LwXyUrNT9NX
qHGvSPu5YPo6Lfxmf3EqhBAFiF+xUYOLQRDsE/5bNtOCAP8lSJ7XbJkF+ck1wCZx
oXxsLHxrrtYdhlVtK7sQpHn+KMEnbUgbLqViwUmxiolFGBO31/5bRx3utndSSfD+
0Uosv/RqKRwiUrxCQo1Pf2EZpC7I4UNtf2PxwS+i2BfGoTW6nqTldsUn0aXhE7gA
B1ZwxmS45+wQazLeTL9eM+PMhZWwjuz1iXnwfqgsFApgltQ/zSN4Nwd98LWeZwnx
wnAHcLIFJiwkxPpfTbM7bXe1g8CtfYH3sIGPiyKDLJe7pm+5G5tByJ54wVkLeCyM
u2OWg1Tu5H2pw6w5Ntb6D1lH70Bf0FlQvjTWHsEv9tHThhr9Ko+ts3rO2fqqkOBu
Kb2L+HxnTtbRlkMml2UlGE5e2McoPsVOdXDpl2EC0ae/PDnW/3KXX2H7ST5DFpYl
AJNPHM2vPMFEFxBq4GYjVW3CAdJdbzerSfJ5Ze9233ulXvKDmkRUqZ9W+ej+Fn/S
qQuzpwa8aWCB/gQExoG3mbsZAFcTHC8PiOAs5BVsBnpj3UwSNx/iqmXLiTdyDO6+
OF6JqMI3ep/iOc4HFHqaUIpvNwKA6dUTHkyomq2tu3sjDMtaoXidOYcv5SzG+RsY
n7z49/Fykv3pluqiqdF0T9Qu7vnvLSP+lb/M9TT7cAXwVJO0kZw6mVaEfatLD+CI
jdwAqYbeg46eDIWUpnkMtoDnAzNZbYG8rlspTu0F5XYtWkk46VFyuPHV4KiLR/nO
r0B8kkLyNkCxh74wllY7xoiHd/vbVaufmggz43oxcCZVNDLXul3LPAPEbQlo4UBa
JP4CNiKol7xpMy6wKXz+PDT17TQyUCzQPKpbGkJN5Z16wNy1g/XSIRHsinZwiBXs
ywxVVAFK6E9pgzBfiBqOxoUF3ZaTm1z16pWfa7aDGlY7AjpPEczUo5/qbQQyFC78
DIM+o5SlmVvoCNzp0wf1aUafLf9fGEuzy2QYZ8/FJEn/EuTxwwxDMRTYq1u8TDaY
SC98BKv5ae7B5tcawtWAHckVHTkYqd+nb7SxtpMBqz8TkZemiovAnp3z64zxx5qD
mZdMadbPR4WAobzIrU3+9wnw4UYNjk2YAtxslOtNo4IIpLmWW+ezPniyJmHwevwe
lCLep74y3E/9fJ8+YaSoZxEkSe08eFjlfwG4/Jq1ORbaNHK1cT4cUdn0KucFQGn4
Oi6C6POp3XCL5HrXhRuVpe+l8GwepfuWNvSfkzLr7sSwjGfU8FjLIpLQDSvMD/7u
Bn5IvsSgrt7ND2CwCzl1hLie5eda3VeFNt9R+zpJcf/KtkZr/iFfdYqqyuFhSUXm
DD43kwr8TTLXIT8VrCrO+VTCZW7m5O76j0mzOgCXV7qIALxyhOo7aliRKe0/aUhD
VdCRBCSdA7XGalXOaI5l/EacslFjxGIQxq+J+nTI5+P87rRZW3W2O8Qd3aHmiFbV
Vh+6OKVv8cMQXA6xrEiGD/viVCQYRPUMQ922liRzFNDDwBJNPzqtaJf6Qsl5SeKw
ADd7c5H2UIGGj8SzQXil7rKTMrmRwAf135I9CJu/CkTc5TW/cg5LNDv/TQSCVNbu
gAsjI7Ll8vvE7hfULmhyp3bWVca1DdBCTaXEKBBi2AuJyA5HrbLCbIJmNAu8Cnpm
76tRp3t/DB2ZC20AHjJONNpRVSzdehBNzGA/ZbUrCl3c3Ylmr3SM1cRaLLvWVoH2
3HRMqJ/hl9MVsgaqDrOL/stk8hSlDiuID2ckVVPF9tuNsWun0yKLscfT5KniuYPF
YrMjvi3c0ULuq78VasKyRD7NNLkc96uDQdutyLBj+iTyyaorTGHOheC+lM2OKNnA
05A+eDCA8USo3Ons2epIeA+akQrFbb25287zKT7OX8r5HaNPACGQmv0hF+u0IHXK
Mb5XPrB9D+WxsTa1Ft2SjN/EdcTHoDMsYZkFW9riPRBU7my39T1q4ctmmwXvfk8d
+v52E7Q1YPGc407outaE63F724N0UBqZRPwKTgfSiNMmq8UvxVSasiGR9M8p51V7
9HEfmSBITQt06C9Luna9kPX8pzzAn/FgeWH5jjPF8Nbd4ZHa6xU50BTEtw+BzTtH
E6dTl6PcrDbh9S4wBF/gYVNRkazdjSdh2XlQ6nARgSWcuEIvkX2V0gxtNL6+RlZX
c3rVOPK4//hs9AdSHyxhKsvdI+K3l13+HJXPMerBvP0i0TKk6N0ogvKxLItsQdvZ
pwgxvE7iU3RH8BNQHCJ++L+Oiu+zFqD9iDojQdDC/sv3NX4OTcVL/pkZnV9mqOFB
TaApEcIsO8QyBen8qHyVDzU0S8KC9YbuCDpmeGHWAQHghNXhgvv/Gjo23zYdjimn
+cEKDJD1Lz5EgFJdbt3Se2t5ex7JuqGD59KPmJcKXk9RPwKksBChYUMdG/Bunay2
aPYo3szrRmgFYzDSso1SaclwXVHUMRhTix4ul9w2Zf0yNVrm/F+GgCPmXIi8vJE+

//pragma protect end_data_block
//pragma protect digest_block
UrbP4TmUN1fPXD3TJxdNCMb24b8=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8EQgkVtnO7JqhUhDgUv9/sKM9qa0M5UH+6Qo9tz5jHHiVwu9juphpaY0CGSfEY/w
Uq7ojxqSicLjoyl90W6VxnbaKX48dXqyjPmsrueUvQZnMvKI9xDs1DXSO2lqzMRz
hQEUkcPcvKWZoUpFhd4ftbp6coSBT1+qy0RBS5Yy4sjU0aBHsu8DVg==
//pragma protect end_key_block
//pragma protect digest_block
qy7DkYRyJutM+dQaKXEYvQwinnw=
//pragma protect end_digest_block
//pragma protect data_block
PSKy47hK1qN7MuwynwbvdN4a3TA7NjyRXp0xPH1T9YPgJYZk/Z/fMYQmpcBrG2+5
gI7cVOVKOBDxcf2l3X9pekvO0a4e7nigFh3CAwhW1wa/tXD45txBfS1VulplV6LP
ZcBQHqicJbrN5uNuvht2dFHFGK9kEnumanqO2UJl4zXKvx5EffD+SIY3HB9zXcz0
vjmqWbWWdVkbuB0t46SPAHAzgTsplzQbrxkXFGEco4jV79vQGTBvFSCmkw8IjvLL
Rw3eJKW9SqRuHe9Bo3gKT6hk6uwW6dC/CgMLXSB/nsuLVn8vMghs81LdRDxmBs3f
m9Vf5WEUnHYJ2rfF6VscAd2hMS8NfeWiV6R2D1Np1+Vm8bxwoE4fyEfRpO0S/m3d
nNZRSHZnJK/sIoBr6qoPP6ifsEWjdIMI35fT5WUA8p5UcLtB945hahW+uabntFlL
+xeAxqM2v7MDZhMAE4OnBjlt/k8ci/MAl6laW68j1hLHWRVucOgzhlUxgJLA0Sc/
UBjFIBYQDC86yiPWjUIBSA==
//pragma protect end_data_block
//pragma protect digest_block
+bx3t7Mzp/NgQfpDn7s3K0gjKEU=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
xqppKb4ywuTw+6n+5jL/iX7UJ4oGVw4EgqLz7IaLSY+oU0vxvqWHCHTo5EikZ9wi
jRmFeK5w6XC33Sc55zTyZO47xR8OXJCKEbh3nLW0CwrvB9FFb5r2mF1uAbboYMuX
TgJhj4HalY46WsBjG21HprZvel4dOE97+Fl9KxkdfYA8uqOCTQ7H3w==
//pragma protect end_key_block
//pragma protect digest_block
c9YMCFIQXGDYbCKELv4MoNt5zps=
//pragma protect end_digest_block
//pragma protect data_block
g36dxjPB5RDpC3ZplYgWfiSEwS0QQ9ocf0z3bVhMonugOdo4qdrMlmHvL9b6MndZ
LGVo0pwy4ud7IUIiqFkQvVUN1H1VNVVuC8PQ3sfiG9OHAgUQz3eStb75HH3yQGHA
JhTOOXW21QBg3QJROR/epRpjSyomKTRtV0y4UDUWZOd9REkVkpi6DzQ323M8NNWN
krSor4OzSnMKg7x/DNxE9QZbsjmH//odpumF/kpiTrG+g3udHord4fj9ujgSoQF8
dFnMp5Raiae6CR+zrPpfgyEeeNgNDd1fxzHS7/uPufcu0HpTwhTT7O0wZnrBnN7i
/BUdC/twBYN10AD77XQyX3OAhziCaBfjl2EouIobBznm1JHTUoiXV2dtmrjLZX/F
xxRKd7JzvosH0DDwVSQfkw==
//pragma protect end_data_block
//pragma protect digest_block
9TjRker1lE8QdyXbLSBVPIKhdx8=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
SMlwqGLXt8m+swc3mPoU8mf48ki1W7ZU8Gne/YDARSjUpCekEsSioq4BH4vJviBo
IcIPvXe2Stafz6SS0yZvXhMn4ZZf8xjcZGRxyI0SlUjRvIyWIuEzsoAc1cPqw2I6
t3iWUP02VINtvFkAtB6gM/3iVgB4drbrvEWiMjTNxdPxfc9jkBUbkQ==
//pragma protect end_key_block
//pragma protect digest_block
MNcjuMKMv2Fp8J3y27qD2l4ezwU=
//pragma protect end_digest_block
//pragma protect data_block
S1www/5qJgV4bviF0D3aVvV8sl7pHln280pU0pkzthOXVKyO4E63ztsHtu2w3sHh
tcqtjBn/v4LscX4BigATZHrpYaiePiiuoQxMixbiZ4+gAnyQz7++m6626m0aRRG+
A8au9aQRag45C6yPjZvyBvGh/Rn3DRrhtBqRWb8Amnb9RXcpOZlQmiD97TaGGGl7
Enxfh0kW/CjOxSDhTGl/84LUvj9wnnw/7K/Y7yoPv7MAZi5ZrkrvFQkzuVSm+rkc
UwK+hdFCfBjRezwdcL42xPNhzC5i8LmbVzv6ZhrS0TO8LiwXQzLFtEUPMIft1hFu
zFHnEynHM/7Xu8dtLYC6XwJkRjitX4STiNpeVg92iUQClyU7WagBEMF/G5dD45mE
p5sq7PkepSZ/zsXoIMkaPUqvTh624seNw/rKyXOZ5jT0N1nGGI1aCw4r34Snse+b

//pragma protect end_data_block
//pragma protect digest_block
GLsWnGv+JWob1Wy7GVZ64miEsEo=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5uOMbGgLSBkrNFaOfbIbB5nlyvWFNYREimY4gwb/SPvysLmdMP/w9uiZgq4hDEhN
v0W451ai6Sn7pPEKW2Us21+MRX7p2K3WSpsomJgWlM2NWEJqV1dN2VpeN8lkL9D5
P4UktLk/jP3nauVtGahfdtdauQBCREeT5yMQdKR0lDiGXD2CRidjtA==
//pragma protect end_key_block
//pragma protect digest_block
I00ZLNjSgkokHkL+UM/On4Tia54=
//pragma protect end_digest_block
//pragma protect data_block
eE9YooIilgZ+MTu0qWEQS0Qb4HuZ0SXIF50qIaflXaHoBufxxXp+489ZxBu/FDou
yiDAQ7npclLLdvCXkJfddSyOuZ+yK6NKeAHnTQXnDe71Xlpe2SKlA+3kEwwxDRru
eacm9eB6P0BSTL+aWT3Ykb5O2Ng6bznRHjgH5fHRih1r4wOHm+VpW8crPZShBMio
6fjJ8C8TJsS/tGQ1dK6YNrYfPRiysyn3DiOrKKH4p9tdl/bt32p1RqeCdz9djhQV
h6DXmE2K/BrPuXiaKSyoMvCbUGlk5jxXDqqhktfN8JWETn2UwfR8iTWPUhNBgoLi
RSbb3eJeUtqkWCX6XG4WNC2OiiamPxBo6QIzcolQthS1Fn1joVRysnn/rWSq5T7M
Z1JRfhE713Ju7zVFR7CC9+LZbECpeazzJJVOxRpCgwhBQm/fXvAprRWfXLRQGdDU
me3J04ZGakW38hqEW+k5eYhEH9z41NBpu9WJnRKhnu9Y47GfC1feryAP5hVpieLa
WrLUxifgvXoqEy/wygNFfcBzB78saDw8JqtG7vm8B2rhp6QLzKs4xb+aUZANXoTO
y8lohw15slF1cvaHZaShoxYywd6KFcLcG/aiEIKWX3qCh/qq2nfiODzrHQf/K18c
M0IKoxjQvZ5c9gpkPwe172UeXl+peD2rTXMeebinZ4jW9OP6XBlIRIbKH6ovFxrb
STjJoYzkWIlSYvbKG2Hbx9RsSRYtXEQbGHo7BUPPNElv0oQXMVLylPwcw9Eowspa
C2O9eLv7tp8MAaqfG2CZ7D64WQmDjEcl6nfm3b0l4rRxNmMECSpeqmoSFGgGLzEY
Ippqu/bteLjc82IkjRUzK2Yp75Eqa64gWedBqs+LV1DpI5YChmb9URx1rm5ZzNla
55L6dIEcAdsKGdp+dD/oZJe+Tja2uEO1CR+rZcOWgoTbsgXzzrZ+IFspqUsUIyfv
n9F5laKrmzRLZ5J6bUhySsV2FsJdSZ4kyy4ObTxkKDcZxPhLBMgDVncEPMAhfdfl
arhqHOCoYsP6G9ATjwM7BUYQok01imfsbj1Z9X0Wv0dbliWhsccBwCxzRX4Xbe5Z
hX0E/4S/TFLWe+kuEIGXDjndwD98DRQo5NBBf0kCE6k0A1gWorHDrU4tAJiZ2Nqs
yKWmKxsRgtt26KTHLJC9OePJyuRfSMwCLFHPepWRnD9x5spx91wBRZH/GNqU+W63
KbMeAFlxUrguqQHUoQGSW0L1XMKK7/4LEw8ZQgKACElRg7yhunfQe5u7H4B2w5x5
KE7QP3mLioG3uhtOx9aNihP7D9WW7qn9QZ+M/gBOvvxPBsNnyRfFvlLZCaEy8dea
mV73QcppOrYKJodt6uRJQEBA6ilKVFM9PYL2LpZwQXcE81OyMHT4mzOo/xKtxUsh
JGZnoNMabeZiPxJZhwqU8BbqdaLZ49idb8PaQRhYDokF4qCyW/RHh6nBQfaJGpAS
/BOlBp6HZQUuPxhPdCG+mRASqWxAx1HIp29HJydfJ4aick0sfmW9AapJzsU7MHJY
3VNnwL0PsJjiXfSESGcuXr+qwAxNo6409lKJSFQiLisETYvO7w2twT/v19hmgLcD
xmImRhCLGLndcHCa6WFiceiY06MhndD8I09SV3OQK5vG0VC/ttS77Hdu4wIIpDEx
pNuV8ld+/IhBfENubORhkz78tjfobmUKAxP5ZWQzs/7ecf2G7IAJa5zIqqEcCoVw
u/PbzqNwbr/5d4xdTcdO/ouNMf03vbw8KYdKlBrYaEBic1B3hEod8fUW49T9Ln3d
r0gufB+uDuNOJTYDenjo56vLnxS9Hk42rPJ4tdgm0N+JZ882Z8uePli7x4utHIZV
c9d/Tno1HDEULB2doodsMe43DqJSeqMFlg+xos1NZ8YMKsaDOCUvBQZOhZyWoNdp
cbhbc4obCGRXt2Ck5+9tXtiOBvQvHZDUPeymQ7aATpigQJ0lIEBB4etTNXVqgggU
ORJNG3gFlJDLI3snycjHjiA+tkl/nvfMt+OZH3o0tolL5KJB5sDfYKiPy8iq4akV
GeglkW3ULXFfDs2gMoE0IQO4uRvJ3zSThdXYPSqTKhxpIAFsztIMzC81rEH2w0JJ
HAO/V3IT87viXDISCRX2UAtRE53P1IRfmyft2er67Nn+nPuJnpYlIjzyx87zBvoA
VeGH5K/vlGUNRQti0CKJolxGaHwmiEmy0ohpZP+bQTAG6pgf3kKMckQqikfwTeJw
GhucJSQRRtSJd3lP60Tim9aX9ghwffHvtXpkvJTF7ehR7FbpRcV8n779e4pyqdth
b1t5hyjTT/UretaXYpwFkRl0UQe6sTs5vPzccRq2qdWlAKC2/XMLpWt9R6/gbk3d
v4UivMRzSVWToLirt+33f7GdN62Z1jFtP6xLEXjR4D+QU3L0eSadJPM6cGRemSCl
t+52W6S7rJZokHG6svKIAPhqcIvidPKhLO9E9javy2s8W/vy/rFUAe2p15MFgReG
rgPthA3ny6/BtzyF3zjs6kukV1Pkib4YrUvzmqPjUViQXmYFAMsdYodJ14W6GZW1
t2i/hWaaEiuU6M8ug9rQBIgYG86GASwHNprl7CZo35SWa3HXwMerLKrl3XA5deby
PJwEt9GuBYsja8IVHtB/r6IL0Z8FJPTq9JrauJjvX1AA6dxyBu93SFSXz9h/eglX
H/IkHG6cfck8IKzj7uZUnRa7vkdY7NvT2wLuEO0E9fTLdu3HXgqKQRnNidPupjIW
16D54GGVUhyYaP0mk5WjIW2JuDIibeevujhDpWwh7MAxdakp68JaB2TtdWhLCQI7
wyzCpeXA18azF7W8LDuGkLab34c6fxmIcL0n5o6q9uzVko88GZC60urqznyxKi24
T8Ewa2wIjqTU0htMcJ84WhLoFe5iVA0lfkPQN8C7i8dTuRARezp1tyn/sW+jfjxq
irI4HKBsnA6BTPYGyUyOrGtFpnBelvw3O8UPVcNom/wRDrJ4DKvRhWCbLFcc35Lo
V38hPu+YFbH6oMwkVVdzHf77GqEfkRKHNOeZ0eZKUE4qE08OYKgyta1T6rNrlxN2
GFlf3eP/rLTEqvdwaOSODWjouM93LQPz46GT56Hppd/fuD2bMwywoB39BjJosvjG
gHhG+ENKkmO0sVdRkHlIVZji7zr3cFfFfnSaVBSADUc27a5E7azuuQ8NmAOu9rJN
qPXkf+B8NutUXuLbN+lSL9qo1U+Xqgj3lnhquYBGU62MIoOORtTfRi5GkTa/rUGj
u3FfTQ2C4YiGe/RjGJjb+X4vMWLo4ixIWAWy+AQAWxh3e4GLNFBWpraiZMC14zAq
AVbmVKZtf1GlQnvBnfw+KiO4pYqpiVC35ztimaMFe9W6q+yJ2JNgoXb6Ai7hOzbc
RYBVMyJi8rT+GbiBLGUwPKjXPXZsZC+/fFLBW3R07qtDaViM4zlZCE0X+fcMM4J3
MW+IICZLZqXBrb+QoZ36NLq/LTLlqv0BUO3u7DoCsepUePkuRx56PlgKiPqHd/d5
fipy66zA56ottP/8N06P9vHl22EwhPa0YASa4v7bzu7DzLcGkBBwl8nzX+xME7Ew
LzPBJiBVYdenAIIZ0aB42HUVdhmgkFJ/hxKITXsAlQRNBxhUH98kKpL/+hxhGo6i
Gig5j6GR7KC060QeaKvx3O8N395rXgBjjdI7KIYTBWbN5+j1Lex1YL3Dbg5gLz7B
bkIokf3aKQDS3nXV0NM5ymD0kMXg7Yl61LwpOSFMQuHlPd6sIikAuM0yYMtpYFVb
rg+pTYWTE9Tt0ynwKickabOzI70byw4LChPEtW+4kDluF6evUP2CEoLHUFFcNKpi
ZOl4FLBQaKl7CVNOH8Ur3EdhYewMull4xfZKbquVb7OnhgsTgppu97w4gQtK22HQ
oEc6SJ0o6Y6st+LiW4NzWB0f725Jey0FsXf1FbZDS+ySGUp41oo8Zxi/hh/fJsyp
YNa+Rw/c7+2pbsYfNICYoow8wKbsFM9FatFPqc3lXkkcO70OqT+t7ZuPVfSR4Xgd
sWfjapWJbiCTQAo082kWOllxKjC2QUiloTDCFTBw3ZNPmvP/X++YOC7wDBvrNjsi
uvMf9aLz4dsMZ7PHfAxjqv5SIy10OUNmnFYS8D4q3lr02JK+u85WGr3d2jiwk/ZW
rWcvonfyzPtApMYdZceju4hqas+OyM1XjJCqI2JfaRYvZkeGo02l04loQPbSeOU/
KmWdoQPfUQY+hdlJldJoOh23rKFSDBoL+fwd5jlUEzKxYZcbpOa+DTqeaMRQLgwg
yUaN2EJLgpXs6CluQGlkq5lVy5FhoB7HMVHIdWvOqCs/i2DxK6Nn8k7hU5W5KitW
N0WFR74y2R0txicebhe80+5mkKADjXFJXOo7kwpMMAyJS4HVzgY8clfwT4mhBUlH
6wcv1snRp3hI1M53cRG6dI6+loaN64pae44kMgyY1LaBXoAjMvAK9pgBdpTrrGTy
lQCPpAXOh+hhnblI7GKleg7fuPc/gidAyyGwuYGbzpouq71Uk0mNlfOGR9IWc0Mu
BRwZvxXgPJ9wipplZyZDUBENCdZmDamyIM8N/ihPQHtXtsW6bw19XubGqagkib3n
OlJeQ9IkzPr4ItRqzvyGmQLMbgMEwC8Q0BPjhXXwdtaGpuJDZ8SxoOxi22NvsOaM
OnjXwuYdoDWxqnRLBLXQaM33mBO8OyJAkkM4+xiz6XG2RFDDE6IrEN7zuxiEjEqQ
0yS3z1S2k6Sr1P0JDayAKuR49bMyG3+IM0zlbWuTst2Br4lymTZ93mWWqEPh1e78
V//PLG88U5GS6BuXzw+0t7TsBapLLOja4tKzuzBi+UcOSh4bbMSWnxAiwlBmqQYY
A8LbaHFM+griKBFyqhj4JVgxjVTQIcNZeqnrP1EMYAGtyJPlcQk/pK/YZTe8bUJy
EnDO8bTmGGmHyryBM7MmZgELi4J+rnViZsvlk4MW5iPTMq6SMa6Cy+hTaPDz1mm0
kFXjBpqpfeDre8AEh+oN7RVGw+dy8xUOi57KG+f8+qFyKqXvASzjzMORAf6N64lw
WqtwRXkOvAYSGX4540zwLOUU92mhAy5uLYRWHCWgq9gllqlHFHlVj0ghb8aIPpTj
CuZshcJGX1WLaxqYwR39PI2sUB5qsBsn4xgKI47p2m2MJlE05/HLgz1wwmHBhdTB
wOkf0z9a/jyPlR0kL4FTmpetaAFeVwprVexbKvzaC/3s52szKrQIByKT5abg280b
EQr/ZJblOuYIFOJ5WUimJWoBj6+JsNvoZq1aUkPVGCfcprxROiTDSxEyxu6T4bo4
Vk1LAUL+2CufcX4w9gzHqdc/pnJFMy7qdVFU32I0Svz1Wo1/pbO38C95U0jo4GCy
Uh5fgBNLe/aSV9imWkdy0IhZCEaMW9NrGetN5OfjM4waHbuyV0HzYm/2g637SotP
+qVG15Dkrw7rz8QV70IR1fOsOoLZ8YBfhA93tv+xlrBVLDBjQiaT4enue8JM9kqW
fq+XADRB1YuoRa+JBfjxHJWtoZ5MvPv0EiMg3YIGeJFEmeHscN9r/n9GOwXM+h2i
c/QMVQ9E0rxleiSsGrfGWk8N+vT6CHLAGcg+k3iKqBuDo8VDCPAsfRjEBgvhXIM2
De8uMZntA3EfT0txSR8pmux1lBl4sO71eYXjFKIi6P//94tm0EPiCjXeTjiKX3qN
53bORH8ceRh35wcS2mOeUm4AI2p7FJjaMXWyF+6yDv/07u4aZSghHdgVqsTHA9to
lO21SbmqURsdvzpcxAbHINiSctrliDLSVmPihEYWmo2MltJXYexH/PzRiyVZbRGg
j8/1xRuMGwfRHaksNWWOGaS8uQNdkKFIhbKbaIWrXbZyoP0HXxlk/lCaiCkyoAHf
gkn9I64qTCVCEAiUphUPXulYY8lyqyJQcj2zLzGkxhK15vY9MKtXGzbwZ1JD+YfL
ABByg6TlyVJxFseRFPATP4VMBqYtr9pw7hjjJiLRZRgWd53fW4gUF21B3r50+ERn
A4y4/2KJ4gBXTaCJCo3eaU/kzzVyMGGYDeT+sBqSF7AWynvIo/CGO8ADSkNRJJLF
EKxbun9KmF/SCK3SsknlA/U+hT4RzQeCUeu0md9rh2fuxmuv5e08diqL7aov1qXc
xk1evlf2K+mAq34mpPKrJoEjDre3e94krOQu1SNn/xmF3pLRuWw5iAbXhgRqLuh3
8p7FxBHYoRgaGFkQ/ZblxGw03OrSnZ3kPu0rSyLRLtgYdITAW7iLwVOoAvPBr4Sm
9UXRlMmbVw0pisSHdpVBArdKT0O8tBvnhXqdoNvX+dSpSeWlO9pT9jbngJYjrHey
fT8XMJKtQ4zDM2wHdLRJu75qRzo0ikV/JPj3HWTSU5EYRd7gDkC4nBZo8MRV6gjO
nZCCH4KKfUmxnb0s/LOVe9Mkettsff06lNpVE2jKmbNK3cr9JKOqFpz5wYWhY89f
i3qC2vOJz7Y1X0TQ3AtzKxAZLDmL9fxw0WSeal5VdjAw1KyTb6wseIVpB2ICvoAu
Rj2zBSbg14LjJXPs/MXEwOMIZce2o21d+8HsOfPQrfYoGELs4pV9UdIKgeYyuMQR
ItB56KLIP5RQjF1Sxs1o7f4f36k1YPAMkz/5m+OIKH7WCl5BJ9NYYEQgKqRISIEK
NaJXOTYVmM6qki7Y8razX23ImhsxPUq5G7Xemg8iIjBWlQysNszj+RC0Fx5bttGL
p80ND7KyShnR2ksXkXdlN5WfOm9J/dGWBWC9vWDjs6SvvzH3wkQKjKYOiE+ZdV3I
RKwZKFCDCkvMYMhe2N82H8mw7/6jH5WMOkMUbAXAUut8DjVawHDvZ3JEjb3GJiVI
WSLMglMMH/GjefvqqQm+2RsuqgBk4Yw+2rdffzAxSzca8lePPs/viojODcG/eeRi
rWQ9oWulrpmD4NkyB6F/3UJM1cQNiIZ1LdovhQP5WqAN01xeOseBB9MAO2kqs71b
AalWmdQDdjy7kFyCFs9fa2NzqGo+WPOa2UPjENdQzCYBYP3QH8i/BAn4+Nf0Ku32
0oAq2K73aXtTB2vk5moZqudVD8FCwdxHb1E08FIct9iqpgGBSqoeey1goz7x2lVx
emzGh//CqdVgiMVOCpWxTfFZtyT8TaOeocTaLxb1RqxewCUqsi5Oe0MMCwGM15wV
+ypgWqWLb50/uZlt3VSbiPe3svfLBxT/xl+qR4j3uuU9L/YlZLRKjmWpZ+dgJpNy
TOCWDqdj/4z3uPXaYfedAedkDXgIv4UOBVRZQappebTIoM8qF2yW5h/Zjh5atVPV
Z9rd5b6WBhGk3AtjtgobMaErPw2c1KMYpYrqrc1H4s0TI8pTdPq645XyHSyyJMGe
CAgPM13Hmm+5Z1IssF/NCa71vgAwf6gm1DcTgwyHHUWxhr6nPDGcjwAKniR8ncW4
4QEGsKswlyX4ivvWC+8S4+QkYNAFlwc+Inb2q4fUCrq86f1EKJWGRtx+m/qRfhYm
0tjx08P0EhPTMALtjH23uviV+71NDOl8udYnZwoSQA6apgdF2Mzc63NpDbSXiXof
C9PtQAEjHuwzLLYgIAjnmgMV5EdjwlkKI5emet5GPt7LSLeZuHctKzwczH8ngQxd
DzFEkMfcu3RcQtEgimZ0Zc2kABaykzn5UB3GE/1l/kyxkLCuKV01R/Kd+9L76VDd
1Y3a1LssfW5I9rvUncaFRKYMqBrOviWZKj9vk6JDXVPC1wrzi8In4lqTbvzEgMc/
oPCJgSGTUXEBPFcKdLkN3rnQcVykePPu6G8hJEnnVx2VmkXRGMClkHk8+rZU2Se5
YO/fgrcAymZW+fUkCMh+sqOuXRKIZZ3Xy7u+ZB8vDSqfLvLv/lg5n6/b1czryQaO
V3/Z7DYOHVYZzz2wNZtP/e09BeA3knMt20jvmdO7Zc9/MNREygR0yl+2ioABwUb7
m4IO4/sBvOAGAFM2lTZ6sKWpQaZ5ZgHIp8mKmZx9w+eWgtOl+BNvhiC0lg9v4cCF
4JFJy54DTqQ94NH1hdbqKEzZ/0mzZvKFljfd1mBA3Uadnc6RcIK3buGsaJyHIzu9
Een7fDltgJ/1ZTg+KtjfmaGh4p+yMhcBoft6XjtoiljoTCL9yDI9PYDxY80MVgur
9f9pct4jxBguWdn+heQXJHSb7mIL3MOxc3zVjh1U/7rklIUo53OmEZuByZ19wJ5h
Dj+8HjOaCAQmgmajawof1i8MoAyVi1Qi27AigtWiDk9GTVkVA6BliPZHDXi1N8W/
n5yjyGglflMXjfJ+P7PQFxyK9LWadNc8AQsLcmgELZf7wy2VLx/b59MOx+di9W4l
MUnttEeE4CaCn6qR/PP2wfFV4KUPc6oYZ1HFxS3bf0A8Su+BxjtQh5dN/LQZpKB2
K2oQw6Eb8qfkvN1monDsMQMBiC1/ZdLLu79fb0QOCQtrW9D3dRzYKZLagIfpyOwV
bFfA8ppk6jVGAMVYtSyLG9CvZ6sVENt7WlMIrtCj9t+hTCO9G72eJ4Nih2jRy2bm
9+iI7ld3jaZEzwgrsbDlEojUqvw2QBENEDyFNVk7Gpfwd7cW8ftZcnG5mJ7JMspr
WsxYl9liZIF07Q4ksqFw5CGyAwICLq7vQ6CwgnJT5K74mw1gOpm7Qy+Al+LlyUOC
cGfaW8Ufc2hOTrjQrjGRf2+uAEx4W3rnfkzxMRPXOMMutCGrLoraFVNGZKOn3NCj
quNkY8RA6FWC2xUqMhEDlP/KYIodo6pDS0KhqltC1sOtyPcljWLo5pfnQg99Xt+l
ctRYT2hvnbrVgGVoS9faPrrFDe8cwP9x1WcNv7/FNCh8y3iG4bzR9h5coSdsl4Et
5o50fvqJXyyr4nvELWMNW5JC83XQ94bqu9Y+Uwi8dA9O8HvNbtwPDQFChPCtQHkl
GeGZeK6K6AG1Qnoo9xig3liDspkABSNlhjjC3m6xEZ++S5zEGrz+/CcQWnsBEdYE
mKMh71Hz8bcgzmaM7h5VtUSDIJm3QFCQGj3iNKK7iXoRQshzcJ9mXL+5wg8jSFmh
yF/Kw5Zrb0v2Txe2RESrbRslZAlZjD9FpReYEngvwr1wjmkrbMk+FdEKkP03jEpf
sVOo8pi21os1R+o5VROE4YUJ9pzivv5J/gXpu6egSIL+GeholWPVzVXQwK60bRUa
pGR+VLePXQEJiOXAe6atlgC0IOyBQufNQ54rH4tkBsrHsG1HJXobQmr4rOPJS0A8
TDtZHPt1GznK9noH782JfK/rrR9yhMrN1ONbtDo2hvpAa3M0qTZM3lb9aCKCzqVW
Fc/BR/M0O9gh1z/5ng/uc96wtasCJSBWrPVkIuAmqfCYzsYRIZneAf6ietWhQ13Z
vJr6d9cDBUii4C23tcJozKvW2mzQ4DYjhkdeoYRdULqXfkkSQV53rY4odQI8zozg
+hPfUCJEPjZ8eV0YP7Se/vre0I1l6tZB6HdPQ0vJWHZw/okBpSU9CRU51/OrJX7+
pGsMdzhA2EJ8IwfaU3OIQYCrz28v5xcMTEsrkBS99hUQwIphP2zfr4V+T5bRWadO
CcbrSvdVaq3c5SGaSZBvAEfFMd4lyuoy5QYjtmGl7ERXHAiGJUuKruUKjUoVcGrI
Nil81QbQ1rJAaobBkE8I5VqyZXWLIgdQt9TbRjGe+DUl1jRvNwBuBXN9NGEoPIZs
n1Z1B9iscxwHZ/JW6aCAnrgKnTm+0RdM8M0QbOIeQx0vQQPvwL4Ful7txa/li+Vo
P68DMpqMOpOhQTui/N+QivsnTPv92+JZXO9h0TEVc/lLAnq7yzLrMSoCtrKVmJ+G
W4NFt2P6QmQo2QN9RLKkvaMvFdWHXjQcSaCE65ESdB+ucdYDi+Dr4uYZ3Cw9ABo+
OvOw7Ouwh3KevLjJVnKlFvOi7hWLJ31k9hzxYcQp8tVaO7WxPpP7aM1DqOG2YKHA
8MMVj9unKH6+HMxapTtlkhD20GlS0xipxKqRzuOqo8dD2HsEoZoseAdsw6yWfJpf
rFZJ/hNE72VCEKqrg5ux80jy+srMNg8Fb2Jm/ONLRJyte6mPE+M0Ls3S/evi09XZ
53J5b7aqB2P5qDerQE0/OqmcAqQGxB84OC0kOD9p/JeLgfDKHX9H3wgdeZvuGnE/
VwC5bAOWAdRiHK1JFQegvzZ/uNgWeqiQesMfo3CRN9wxgAZjclp6oV5BVEVL3b+e
RKFd1x+V+O3TN3UEP3FJJU/m9/wV8hHz113eDTD9WEhm0lkkc3gVJmdEL0JBCAO8
kY0Vk04J+sJYktU5czBvoy6aTxZ5doXR2QEV/Rw6yU5k62ZtD5/UxHDs01GPIPxh
UsJN5h1/ZK+BG9PldL7Q0dpMemPtwpefCkDDCTjaxJkLOHcEL7g7ZQ2KTievKJaw
eqmPPUfSshfg3w2R8g0nEADTQuMgQmO4WSZMwf0FF/PYsLotmAj3s2mpo5Ad7tfc
G8I7CB9h2IP3you53AVs+XWP/zX1gfaOeA/vxyJfjCu6r7Nq4NOE4ACjflOmvBEd
ALby5OwZVHuGzUYz1246GXFop5HcUw5DlwPFWhh2JRY3/unL0gkjvhw3TpxyFPny
WvJ+Yd8x2lZ2mDiTIbpQiCf3N1FbZxfr3Xh3+FlJ3tnU40FUWXHZiDNP3laGNz8+
ro2bPKz7xzTVH7e4ZWKrhAhsJDmypIHNGPkavgVriCnBbEJQLoLoWUDy/NkXklYG
wjSAlrkXzRol+F18dhHlzyP/riwYeLXTI1xBlpxD3TGcWUsctYeUrDZr6uZjfUSB
dXANEmN5KHcl4FQWw30aV5eiDjR3d2pwJEKnHo/MxR+gAfvznfg/2d82Pwkfa0YA
0SrXJMTLQBKSMJr7wNjGl/KghG0YBSU7p8PW96Ag+b8MuAf9dBGWmIKdV3H1SnuZ
ENtHoULErPIM4Jna+WRKOFGSmIhKXXA6zUntJBBatYXB7wjAf7BULcrE/lT0GVhh
8fvw56KTYrA0kxj0w+Akg4ChAbaneJFMsrtZ9bo2Nf41lVHPZtnu4H9U0FtgTxut
my31z6akLFc3I+AHFWA8vXlP2dkBhF7rUDeteQiCupdDeYqTsToig9KPQdv3DRq0
FWCqB/8gQlHXw+4TYUHErjR8DpX2rtUNBbHkKXJ3V3X+Ht5grsEhU2y3pg+5vVbm
yPAEL/T4RYZYzojfa0sTLopUgnogHjxVYbiTtxOMbpNW9dmG8MRon+L6n7ZWUPlU
CxGgKxKS5Qn4y7OsylioD62LliabaVvJtBRGOuxlMrPvxSGI2ozT33tVup01+NEu
dd9alYTyRrRXCbgbPvJ+AcFaSpQXF6za6oUk2RKeph9g/170do6S5gjFTgu9cs9n
ZKqbiAzvgxu7N5WKjG3vdzl41xBiii3mqQZTYThxrbDyx2/ErEq+Ubul0I/ZlqFP
uJLaPJg4umYih79ywKUDQ2To0fOmFp7Cr2T0Ci4PJzfxMS/K9FVGVYMUcWCpZnC4
6M7lqN2RIN18NBUn2jknwU34xj/2E/GHYwuGahbGBYrjcW/4xZg2Im3UuZEbaPRK
IaD764Z0xmSa/geIezPG/4sZM4cobwtDTBwnUOKBI+mdGhYkM75PI9brhPVkGq1B
TU9dPVpg+FWwdLpRPkkOi7iXSp/zlAn/+wnICg/ic75ZvP59aajiaKIkgu8dkhPf
a5gejp4QQmQlihXc0OPdJI4P0DhHJBPVfAtCDCF2ICDXY4GRyZOI2zqzOA8HpWiq
hwwJ6OT4tW7ldHMvDzB5xf+/Hnw4Sr8jP6avRzBtSLwG+781PWrGKUt0/JO5U1iX
wLeZ6YZ5/4ucCOAJ374XsUHq59cCgCNZf4xA1OItj7boI0+ffu/8cEG2aPRb+CCU
4Qvru3LDMlYS/nJII5yvqqy7MBmvLK5BchM/+LrkyJaKLowl5qkBwyF9DtQigtjN
Ui81xG6v/9JW11jbMT18N3NTyGiWSwC73myKG3VReh7FFVddPACKVPvOi8Zo1U06
2aY5AZ1it55kqg3Ie2Ba0DydeGBswOc/6RMLQy4lUrV9tZvIL401cr7vcOqTew8L
GZjJ6b6tdmQg5EqBovHjfhOLBiyF6NRR8fW6feLeH5SPEWdVxhwgN2y7XTJ4zxQs
2w4gn/6O9O7E7uljgAMhFB+T8WY3y5+XgwBhXTj20XwE8iA0KQ1tUp+4wqvBL+Er
XQRloNyKPW09Zn8GpVryrqpOHTr+Ekfx9v/h5gylfs8XtEPTv0WmPNUXbMWz9E7/
a1VoLjtopRrRwRhBQjA2fqUi3wHtoh3o6qWy9lqLlpIZQW6mao3bMwt7WGeVqiY3
gcWJJV+zxrjB0+5Oi4EX/wJPzCe0mGMG2tGZNdHZq6iNrY4CAIPSBgleK1N3Q2TN
NdZ4lD0bKHD4cKVzzcZk4GJJpi70tQPs1Nq4grndK3IB+QXPs4RAFYTLIeYBaEIT
wv7pD/4NusZiOPcsc0lvxByTkrQxFAo5Jt3BTCNNQbqvsBO2zgz5jxYH9vmqsN/x
9l7qJre5WTWZXNp3KAYVG2YW/9+VxiiVwotnyK7SopJlRW3rnp6ShDBfUz8wTBqZ
0g/srVny/0ZfM6li07ROqoyAPLv2Ev2iw1KAD3kud2PCcw9zuXtV/2IfOnon8k2f
j2L61HdFwuzGGQ+7Vvgyc29eHqMxpskdWty0IU8s3MpTq0IoI3uKmZM0Ijy3ysnv
NPwAvDrePglreJG4MTB6uEID+7K3+cOGaJe/3g23e4KnrpkNXL+rfh8cvE1RzT8R
rH9x0VvX3XNq//5YhgfpbGKYb22moRNMik8+hybAwjfdBRfVkiWB82s8+/dDk5cW
Unzx8JOGPdrjvpfoMG24rD4pP7B6CPAg5i4UAFmKZpcDOQdH9DP8CYKR6gkZvN1S
J+CH6omQlWjlpjSVDy7Sq7K5cCTsB6t6j4MPnQcwwjCXePt5d+QN4wDC0FvYvRPk
+C7Gsm/F/nvtyT+RTquxuNVIBNQMpC8uZIABWPJUoe1NuaIZNiJvTttk6ti9hADr
jAa0qyYoZ1unGOcgknasdCBA8Qfcnf+g9Mgw6CMhMkzIp9LastTwz1MgBSMbD6Hn
9MR/aD7An8EJu8XvGXFCY3AXhFvDhE8wKbgfa2O/pFK7LPlNlbzgc2HPQcSxjCK7
7nsuuxqfePo1KL5ZJCOKsO0hVHt3Etajza/rkYAcInBuPs+kDFEAN6kyBklyO44I
mj2C1XNY9K5XMoxIJZ6j/3ut3lNw9lbYRcHBIWQsyHHLTcrtPRLdcfLWWHX1/JVS
6ZY8s7kfZtEUD9HYNU+SPaHAx4dil4Eg73P+JVoahhFodzqTMKl3w6pmpX970WFD
W8/aRkD6r767NUrR8Kf25ChhLc3FfddI1K5pLzccB9r/u+9JHwpJD81KzeQLknXZ
50qsYlQgBVqmP3P1BYLOxeG1FJyarfsivgUmW/B39SO8PvvXaQgNNpYm2T0xK27m
E6jvFdVeeCEAv71uiAOISduObdtPudf+gx/p54Pn+FjPAKS+8PRpK4yuLUE/vYcU
+xb9HvKn2VvTCzcH2d33QaGBvlVRYq7EbfpUzk37V05o7fuc/ngribsbwwcNYKhe
FmaInXYdCKBlD1KwYqkSUupNlIivWQMx4hEQfKDOMJ0CATC2ixy/1LfgXp8bbsqv
NPTL4AS3Il0VrcgNLLaXaKcIuMvEbv14FwIpKahQQzrEBtD9ND0imn9F8OAARcs5
+LB2hXLF0k61vm4i9jKZe2L/U9R/ofhbBfNMe7BzNFa+qI0Ws2+OBkLW8yBnbQhR
2r2evn2baSEQgTtzjFuKY1yTn2Pj1NRSns0xndudJ/ihZ96akAiWGGBbEXvX0YJn
LP/njUDVooAr/aDeqGQVWsWds77UVeoMsiXSin/PU3a35nK98O7fod97t7VpvlV7
XEMEOecw9EPCWT68eTfzrGV9gJivKJ9gzlCkpJ+MgMpGQp66PfXgeOMtstePe/x3
NAlXVhmmq72UeITP5b+BS0N8DFkUeEFYH+37635eqRomt3Tlx/6kaaOD/5FDQ3ER
KKDlbO8bC5IAFJRkIpde0aNSzVbjJzzWfFX2BCRAyZD0+Cc2iYmWERG7Up2uioqj
E4cKKial66LHJMDvVURT9Gcr9uXfBhMOWDrlvcA133wIphyyMY2M96/aoCW7lL57
or5F6jiR8OavUYj8NLZV1eRRxVY3+n2e882/ejeAvAOlq30clhmYh8NOpBWZ6K9M
RMl9j+Sp2knmXUQtA4onWcE8JKDnPikpDJew/EtnBjmFXsALXUjwu9KWvn9DHO7E
NtYw4JeY2cXXuMGfXnI7vaqhlOlM+nRaj9o/P+9ITh9CSUvWbjjRj99ahiO0Ma1k
aad8O1Mzte/jxjKb//8uRzKDQs9vojovF4AyUd1YSyjSGcOTdlLVSpS5wlb35l5j
MJFbIvMQJof9QEP54PxY0Utoj5iYWijEQ1pWDRz6YtX5A964GShjecB4TVBzK3ti
YJNAAL6QC73HBcvL4CtpLBTHLUQ8dSkOGd6yIx/pjuJDV/vutAhgr65wcD+6VG42
NqCtrrl4IlPAEIWQyK1gWBDlaBuc1+ghYsbU9u35q/aO+crLQDj6g3A5DtgbwNHL
NQltdrepruUBD8bJuqWt4mBqc1Y+D27uotPloVL0xIDPyedzSZo4kXEgtFWu/RSQ
c6CmrUSzU2QS1Tv9Keqk5/9tgo11NcjTbPdd6R2faXUNFXW11uh1Ji1fOiBsR2gB
VXZ6C1dr1TJ+GUd2m58BUo2JhV8dggyFJerV6noTAI8s8bFAbyqw5BmrRzIUE9Y3
TLi9a8DGsowegF7rGHRH2QUgQJdtNAkDwiqedzA1eaW2H4qzOUTgDDU6lOn/XDRM
WP+u1fVpV78ugPR5hgoLRXXAJop2PMTOGgyVFZ85+CvBjajiv+HPuBiDeFiOrBSh
mihH/wq/daSLr7kX0emrWx5gv3vXLIBoQAK+jcxxEAEW68HO9v9SKdKs183TySrC
JdqucfyNzJ9EzqDm7d3itaas1S3VCgUCcKKDVOoAKqPUbldMH4xRQWLwiWLk3jiC
m6m/3VqH/d4wqxYFxjgoWtgmrJ3BQ8supvznO9CmY0ifbA+Wyxdz+eyMa9Gc+HUx
rgRDrImwq5D0P6Xug4aJBNeJe/7mm67c0QJg4cC0eIwZmsL0AKHbMT7Jo1LXoiCw
VXg40nAL0esPJwJ2Ou8qSjfd3QWN2d4WiWlN0Sg9XvQNnqkSTV9U31ZtYC8McU+G
NWeJtyuweN2VMw0LJSiGkOcqcf4Ji4+rMgOJR+AtjURjUmdLe5TcB/GVLiH3pBl0
TtKw7K/dMfO7rMVQ4TmKrLdP+GKbEM3INlkOvu/brPKLgfuLLArAYjT2R6/cRDOD
+0sRj7aNRIgD+bb6FHO58qYwrhgryoZZJ317A+yX/t4Y2XjvGwETPjWuHA+HF+nK
biX8COTh/qXt41mc1KVA5qP/JpdCs6qIUNsvGDoUolIAygY835ynt5MvmRVmilMq
JR1JBfgbiwjfmBFBIWmkOigBPB6bejMCvvYX7MeajpLjRDVKC9+cJJo4sJjwWDqa
DNUdjF/Y8ta9e3Q4DST8BQwZuz+4S1kxSoWi/yjEopy0PDYtqOT8fDiRBPr3dOPq
HmQGWbemajPCPbbXsGuoR8cu/aM/7+yL7Z8opS57Vg21Jz8YV09RImE8lLKcFMgX
oYVIAPRToNa0B/1/P+rC3tgpWUuKpNXA2r0YQlXR/FKsGN6UB571pdRAyE1YxSid
/F2oB0rfHGhekfb17tllpi8Gmwhefn0n6NeYkmnhk+0SKV7fDRTXsuwOwZYbrNhA
fm/u1gPKJgZQuzjYz0oJ7jyCmu1CzZNwwWTi+YX8mSYwvXd76gv1vvdGkUwzTfP9
Po4lQbR8cFeeR92p/MVn12uWsXP4AbPcGKr4I5p62BAtvyFB7yx+AIpQsoECZ58m
BsPstu5EY0SKGGp9YDPRXxoY9BHbA+zG0pqJ7yx5aaD5AD5QAJtMj2hGcA2pGPQS
FM+yu5Cnm/XqNgG/fAmYXk1qkX/m/wLb3mdAYVkaLhV/vFOFQvjoVvBxYJUWY4Y1
RKE5ieSMlo3KqWawT4LNmdA/g8a9qpMpuRsn+ybPY6q2hJBxcjfxyu7rM2BeCKW2
i8qkJOiyXCnh+e7/gexnPaYy3WQZS6WJ31O3tTGZHCLla/XhiHytIgiPHYCwAGs1
8d60CWNV0VoYbLzg9txDGJGV6NO8tePJpOSThzGE8kv4HIZdNOGR1/94ifnQOKLl
BZzP+DmSufSb+ztz1JrEqgx12LGAvtk3oUH3dJT2lG5pDR7BUoI5nky/FqWCFNAz
8zRCjAKhung4HidWfR/rFJS11JlWOwe02g5uNbyOz/pgCGBroKc3QketHDGbp2Pe
pn4dx3YMuicZ7dP3pab0SNnlcos46mpRf9AIseb08/BlIKvw0+Z2fuCFzz6BAy/n
yc3FjNUNIiiUjAMTYC1cwOqFXoQN3XoNT0ax6cjkpd8+yGEVFTuEPAin1l3UnCMc
wVM5Ov/vQOcs5dyUHHkoKhU/IqQNsLudMmwi7e3QzSDLzkFKZa8sIwhQZ1+m8Lr2
NQsCEO4FFsVlNHBp1cyQUS2OMgaPBOYdjg824+0Tz+eLxEfHQ5K86Onhm07ToKB6
GJmdDlcJXcUxBZiK7m+fgf8Z3NagSo+kFjsOvWrF0SrhD0MYJPUrKMrXVAG28LR+
ojUdpFQs/6bL8Jv3mEIqga+FOZ3nFfW3Z2PcVwr82E6NgZ6SnEjWYLj4ChRB3Nah
tvcwO2j4182k+CGRfR64kGauqfzrcc/ff8rwtJHijCIzfTkBZOYey9U0dPhUXI29
JDmCbncDnRWUHM6lAQg1490309DL81SJuFQeqGXqaO0z3Jr7D/IdZPnq5jzFT0lt
2BkJPqPd5JMcTPTNIJIEeSAnWun898maes1PKSFZO0umAVr9Z1h9xP2ZNxHvlJ+O
dD1ohoq0zIwN4+Rq74QiF7PGWGLrsJ4cdlV8fELQYZB0OPK3ptkOQip/R87eiUF2
0il/JhvGDZ1FoMmi6E23rpl1YjOT7y1MnwHHoBQVt29SNGLmu4sloZHwDykAA81g
WtypaMbNaSKk/pV+mO+2csbDqlfYohKfYT8+qKYvPvYrXTpLQkMbrcZY1WTE9VB6
wuzbPdB14jUe1GH80n4Mxa+sgzutx1nar0e7SQnJPUBZgBENDec4Hhuvf5lp+6sf
Gnq0jxGZBcF1av2+EdwCKYdzIAK5t+xMxU0Avg0E/MTk6D/d0U123q35w4q8xqdB
3Ku2APrn0SVqtGB7trHLqrLG1oMfGzDFtsLIXnArwKiUh9IAg9I8dMX5X182SCmR
02Iccraw6BlVzr3AxIyVv1EFqCl94/SaOtgEzb4HcYAxAN1fZXFYqM40Ju2UEebT
efNXyOXoxvtZgwHuJn5mDb5AX2jS2AewneKNH7Z2PGor43LQ0M9W2iEx1KsmQjOs
gSuCNd9qWqSeeVc8YdkfkfEjMJvzShkMJ7M8gmKLnGRmwTnxzhjxEGiv2JzUcCN6
icr1eUqUHNzFIdz0G15HXK22XHaVM8+WSQ/fpphJgvpGuGlDkbhRNxGmwheggNf2
38JPii4rRpZM3UiiLkXi995qMy7ljo+WWzJiZ4MX9ntWrIrwG/7/vxli22bxirrC
ZOs9Oi48B4C9WprGjqDZe5ffS/o0ArBrl17ulBV8L+P1hU4KLAGVTXiziUGrD8xZ
t8Og/aRyUs3BzYdUjfKbdCdOVNbJZ+gemUV2iiAOT6b9oznQ53+7ZYmip/y6wLJI
QW0TxfevFpaMHEWxL0b3BKGpyxjNv/051HKABe2Ie3Ssm+UY98iNFX5hz8SXjptL
KjtFoV9yJWyaW89cK9fbdHLuVxu8WJm7XLt+skE/mw2olTaYnO7Ui42+QwUM28ya
xzKolKtqjUtg98liEIMVtjW9QFSYtxw5iru045ppyWshhJXfFgUoSSs2UtwgrJ8e
4SUcNwXt5SLLGTu8GFs79+2WN+aQ5tfa8IRzUUpYbbjjrFgDNeVfICd7oli7rZaX
pPoQS8ft72sl9iYKtctM3ZrvBP6z7p5IV31xMS1dCqF08QE/JkZrWnoXOjVfdUfL
+Er2RTAjquZpHSY72BvHjqtBYqlhxOnhZT2DsLgEhA2s+Gp//Lnsu2mAyLKA9kcV
hlAy6Tyvll7lcMu2Tg/Uex1IbcBNBhmd09bJA9npO2Lq2/Xh1jzci41F+GPC5OM0
4B7rHfO+LtdCALRZBk7mcw==
//pragma protect end_data_block
//pragma protect digest_block
W3qtyrWKh0D2Jtl/d0Mwgj+gwvY=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
tKDlLN15PDeCzyX5kM2eoMxs8UAWB9s6pAp6RHKiDxloz/W28AKDK8D6Cw9kejBz
lNn9Gd6MUK1n2CU5dralyZJYLgpyBjMbF6oy0fVlfZm67KLAPhaofuy5Cl+o9YSD
xLAs6YcEtf+WfMQ/rOav+aqxY8t6WwiW9gqxmXdBCYUrsAJxrZYVoA==
//pragma protect end_key_block
//pragma protect digest_block
kQN0y4lLRJ23IC2rmn2NgnbPz38=
//pragma protect end_digest_block
//pragma protect data_block
IKdxVCnUrImTelMVnWRRB+qNJswt5nDzSmMzjHvZHJPMfJIP4D08gajetInOM/vu
LfUEdkLKZbLbozZ+6KmvY4irfiJryiR8t7bgtvo2O73pb65PQwXb6tWdaiqv/QGt
JfutXrZWC0zTuKyzgluQ9dTmSWoAWUqJH8LA6NeNJqzKns5tzYMKTS/33nzBXAmj
m5VFXWMXF93NZFOPIGZdB5sQIKoT/gJL/OJu+Qr31Gk5E/v8rd0DWEJvsIZj11We
IWjXluyRBB30KNMioPb238yXw06nKxLWi56UQMUkXGxo8KpnsQiRQHcvC8Ds7cGA
PWeYB/uFSpcaa7iF/ijmvOm7DGNitj2Pw9kBgIIDdsdwEvWu0JhOWie8Xzz/JBY8
X7jLqFxSTREy3fG5Ltb8JmwU8iQVHDPVYxeRGqihpDcuH4fJ3gQPpYfH7zDnecop
QwG7xMnXOmmY82t362erXH0lFCQCKPfdtmz2ZmzWW2K2fyGI8rGiXon8vBxBNXhe
21l6O+264s0ImIxEfZlUEA==
//pragma protect end_data_block
//pragma protect digest_block
LI2Fz4++7QB0zC5x3VY2R9mYov0=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
UapcMYLFJtIbTos2eV1Xncfiie/OsC06qWDbtwCHITal08jAQUCjtv1CLrMuCo3G
xycj7tSMWQlPBalj7u+cEMCwvVSvganvvPFfpXlLJx2pcFdiwTl+e8wVcG6SO+dc
m+5QeIVshGu3caJxzl+q2NLBy6aLU0nBnNF6bLbEMfqnI0z6b5/Jdg==
//pragma protect end_key_block
//pragma protect digest_block
dl7RgFMZBHcezYHzOaj8yMylsa8=
//pragma protect end_digest_block
//pragma protect data_block
2hCo1EwVAocLD2WiUqGOiY7Vze7luo1FNMkSgeL0IgruPrh8WVTZywD1Mz93w4VP
DWN39SDsGoASESzhAwBwmNaUX5Xck9pokK2HE5wFX/fB1GpiLDkQuGXz4HdUtzk3
PGOk7z0HOfmHeT8XsrFR4tYEhSDqh3RYIHaPs1qtWtoBe+wiXlGiEZMyLZ/4vkdk
b1WvlG07OaTc9sG6VLKsLidB4eLpj6oB5ypTtym6/ylIOsyYPt53yF7M+1RhTrCv
mefCIqyvz7BTJxvZYddklNQSlwiRd15fP0F8Pg1WUodGyZXYDyuaXZzZaIXDI+m7
P/h7bVHC0mGkF1AIDjeWoWVV+0/aDmuYfgZgpHPsM8+QTp6lZs765lE4ejrGBmmS
VyJSqIkjRXZiY4LaMpRC2FIUcUtfzAyimCip/UfodSCAr2JXaHg98x1baKBF7xbM
DU1oR64sKCIxQaVeEeyUN4RdY41Ys69FxffXBEl25GvabdhLBhulQ3YMwLQGda9F
CuK+X181zI9Gn0P5mIQNAV7jiecMswWVRPX9s3iJaCafXMS6MYeubWQspcTubiN2
U52N6KV3iMZCBxh3PyN8WM5YDvoL8BIV3n1qGPeeAjlgIdIfBTWnq4qP8u60uDRS
aOH26taabCxelKvTj7tscy/MpNEsv2rwiLVIsqUk0TDvNRUR6mHGJvV/cwkSmqVp
I0OeRyViIxr6o/fr4m8uNCdbu4SJA3lXpyD3IDYcxfiLkhwjqa8EjWE37e7EziSj
FJtbV4d12Naw8lqi6WNOQ57w2W8PcPCAuBpY+tsdH+iWE6SnVNADp5VSHoXHg7uc
mwSYz5WLhEhtdA2WfrfV/XtlTlaoII/a0/5XMQNQ1uB4tpEHcI9tqdfqEX20iUhv
WeDS/ip4xe2X2m8wkpkxeywbAGjvbsDCkfRP0Tz2xJTiyQmNULXewao9GMXHOqEH
YG+6eGltQJiSS/6vEQEoY7T2zq0D8qgakB+5i9fqOaa9YfrEH1qC+vz6sKwe+Nmk
sAZYGT4Qg7UfXu6dy97FYN8Joq4w4rNGT9UPAjnsVslvQryLwor7oRDyIyjM0ANr
I4eLeJOtKsD+EYdUpkkabID5KkAjqJEuXfE+LXwtXu9WdYGvEQ/f88ohAuwiZUWk
HJlRHb9qJujjznYaFv0KIweSLH7sbKXSTho+JMDWaM73iDUyiufLsaNUgCIARmfL
0exE9s1zfQUTVCvCDyFSfmqS4i3sP2ske0H+70uFOy7pPOGk5ORzEhyiTouQ2Xpj
LyuGqeH+QJ4h4eBWDDcWBnDc3nu3R584bY9DPgfAL0JNVPOpHolZMqjWDO99/JN5
wREjWCvE7mqnsnBn93QERXsOgaNMoK633P8GfdQwOGJNZZp2YnuwOm6fiv3t9Mgn
q+erp4ou7Qx3oScpT8O0kUpxpbLpvRLzn2T7wakFbZ54X9POY5xbJy5a6R1ju1tL
1chwgMQkqqIf/Bj1b1hLwTUlZrPY88Da4KqPVZv8hqRVMGPwexge+Wgc3UU2xtX7
WMP3+u55Srass8wHvVoE+gPc5jhwfBtfi4qtYgGSFPioRN57ZkyD7SLFjaxHQ/cU
U8ofzDwae5AqGvBNEELNfoBf34nsIwTYU+qS4dMqvt8/D4DNKjHUyar8/XfqNOos
3mHFAIJNLBNQmm+e4ZeS4LykWH20C96OFH14xh/y/CSYJZSQac2UbA3G02D1CdVc
fXt0qiaHNDyGc1dkGQEnyY+QWQqBNF1OXW3q897ky0j+V+OmuaBgQrzoEnLDafD3
c8hYziaoFjFdhMnBSBhgm9zHivjIxX1g5QeKPgoR4re4wkC2fgIcn66yXW5A9JVw
ElRKLs0L/lNlpFF4fVcBNbmQj90xdFlLn35CO28ZEuqpyZB5SrsoL9UO1Bp7MBuy
iXo7RvQiJdnnSc4R99eqlfhJOTz1rWXOxAieNL2SRYkcSS3pJ3QUGWQOM7RV8cjh
1DlYc6agtkdrlAjnZBVA5qBd5CvM6ZLA21hmbNFQmZsb5WEleUVIRC8irt1a6tXq
fpWLk6dYCpuk0njKBIroVoX5X7NT4BzeWyYlHCemRwz0WVMbQOxHA7wxpa4JqYhN
YbLB//FnbJAL/tviXOImGjDeIaV32appn1281sdtrUqndV8rMqnlFNbR17DdnqiP
mVkjS8/n8cmxqy4Ea6ajnQpHg0VHM/cKoHR492tNKM5HvwKT/nzB6OM04TqH3i8M
iHYqMmyFL+zl8gcOZESP/ryhSCq/B6X3prPu1pug1NEsCXjtVEXureOrOFaTq6au
96jV1MI3vnyGzUswZZFlSPtgKOK7xQbmsjJeXxoz22LIgPGj25cDdaHt0tmwvYyg
PoLNoiVzCr0cZBbNpn16VJyR8+hjFGS40sj9Y5LBWAXYCiEulm0Ow7zSkuebP3PP
D49gjAH50vw/yOJi5gYMJMuC7g3e+mCL7pczL9LFarwltUG5kYQW09AhWt4rhXLS
2yJvzhcLLS4/sDCSjj7IIYeAuduzmQOqeIG1+TPoJZDgTW3Vpg8sMj66Np094C6Y
ygXYoK12UYbrUKLRdg1FmkN6ublDRanlLjTgjMQMGnGGYhMmecupR4my5dLPCbeD
7oZuszUDxTR3wNCbBnQPC/xD50QRmR5G/Tapfdd4ltF3/owZ/qBQgg4ikb3+X8ud
rdH9pPoGEAMoY7a0IJj3GMx6Y30lG/VyHOo7IfSFVLJOlHnxVCH+YC4sNGChXebT
9yMASXnAcAaJ5CH3NeuaqZ5aBT34CBSGb6ieswmL0S65wyNu8Wv0Uauz7V5EMbJ8
HSrhh3kAjGiqEeUv48VDug6GjyTLdsZjGefBXMD9nVPFk/xrPzdgTZS7MxGh4Vb6
FCuc5iMzJSeX5biC8l15JPpEqCLrNzUxK/jhnrOqnC8DJWViB1n4e42rNuwoNXIi
dYMOO+OYAjqwWy7PaVg00stjhfV1ZfgkNM14xqz7MnXcbFgrRo0oEKK6hsZ/M1jn
Lj4dJjbjgxLT0XLYjncTIwC4L7yGkG8v5zBgKX8RaoUG3VmKR7uRhVfM8FozQtjv
9okJ00f0mX7Q3KiLwqDmu6Y1LczVsT4R2LUcfUq6rmxzt7Qy46+CWEjJwW9xrI+F
JT/i6bk1ibqN79LgNrXHNmSxw57jBLCbUsuX0th76sHIJvisCElXkGmM4bM4lO70
3QeGtbWL9bHGIZVEb/uZIE6vIwOvodVFnZkSX1L+GczwMnIy0Ct8h5JYhxk1Ti06
19w5GNHuu0BFTp6Q8O6OP1vmZ8/YX/4txYdsO61bNZNbCFBAmNflXjK9U9Z2wKrm
IYr2azknApe3Bx/eUVMPUGDp3Ou93A4mppDvGdwhsWKLHioKpblbsTU+GUaygz6T
mCTSVA6HUvSrMcX8c3LX9/OQpFbh55uXK8/8lze1hNJPhYb7Z+4/fn8vd7oOmbk6
XPnAucKptNK8f/67sYzmTDjd4Bzqx/3m5aIdBdx/+QQ9e6RcUZB956i/wYTXyMhK
v1AtWyh9eFXR5JZ3+lUglPleby2OqgGTSPr2gXYPzm3Fu9R2fuTleM7OJzcNXxoE
J5tzJfcINy/WjrqXCH1FUfUjLjQS3ArO+EDBg+amx8HIpB94/JQmd0YjADbozhlk
h9JwkKtDWGRCjMVsDSoPLdcfSsFRi92da80Hccytm6RozO766aFHswp22gbaIHEs
ewZ+YJ49Zzy3YX7+iX4mrrHSn3Wj+owW53bBoG4feOXFk+LkGa303hcOv+btw3OO
9WTqKjUwIPMWeXQYXEHwdDtPlxwdbnHa1tHa9ZnqlD9+JLa7uH9ScLBsnv9oe+rg
c5BmEhKN0oVt3IHiyeJ21kROUgXmfP3HpKKSx5ggRmRCmitTFmbxKzlp79Wy4DLi
ZE9he6WnTciK5GV5l59KwH6BvEHar9LRjnZ25cupia+S4+iQsV7HkbL/Sy4DMCRA
8+rwOrDDrAJOs55V6BO0a/oE7uZXt7wriPdCMsxzP+w0dE7JGvNwfhIDOOF0UgdU
/eRkx6tLPCexBlE0tn3pddsTB9Eqm9oTmAd0Kh/uPDg3riZnOwsOXRqNrkbHO+i3
qPIoET+5aVsMBs4XiLj+456US5pTMlz52Qs10kkTCaOPiCy86deYUbtgSxnsr2VD
CuqyErwsragLc79vpiakSW3sCzSkQMiHchGYQxeFDv4A/g2lPN9Lz12w3NgU+Yng
zH69ZrMt3qCmOZTJW7Mqp0AgMFqy8oXD7tdxhkTXKxNkD9NZIJytCsyTmKA+Smrf
BaygbyjD5neTmJrEbZjyc5Q87d6NJcrdyMXYJMdttOhg4U6P/Dv0pGCGBxz/3Qqf
v7+l743NWnc3Ub9JEH3sRSpD64uNkuhAM5xKVBl3hippqJBG0vMlrX+zgAy7eo+5
BhRsFdiXHHHQNkiWuekbFyhX740K9iJ7hOVhN9zsEy+bo0WsxA1nCJsyig/nR/vZ
8I7fFjD+ehUGytNLg1+A0fQt4n4ZU2eyLs0AT4wBz0C8G/6ln2Udge7z+DPNxG+Q
+z3Q7zIIcFGjV8Py4Lfi+7YnD3gtNfTHRq+VX3oCGd5AoiRAte8cg5jsVgjyk5hd

//pragma protect end_data_block
//pragma protect digest_block
d2QoA/qZvswcFGJ0a9pGKSxKW4A=
//pragma protect end_digest_block
//pragma protect end_protected

// =============================================================================

`endif // GUARD_SVT_AHB_MASTER_ACTIVE_COMMON_SV

