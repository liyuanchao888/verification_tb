
`ifndef GUARD_SVT_AHB_ARBITER_COMMON_SV
`define GUARD_SVT_AHB_ARBITER_COMMON_SV

`include "svt_ahb_defines.svi"

             
typedef class svt_ahb_arbiter;
typedef class svt_ahb_bus_env;


`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
d9lpraeeXyVqGtk5Ekoocd+eSLciNWKdn4cGm3S9fnJg0n0ydorT9onoP2155yP4
JniRqIufnEYkYFBM49w+wdnF8z/rbnT1Va8F6zqrYzM27syMHxkCEqzONZ9ntZU6
l84YSZwFfko00BhaxR6ykXER4mdRilrhtbPtE+XKuvE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 3362      )
nVLQNJ+PKhlQRHK8Q1XHXU58iltTZxC9ePDSMKFoZBDW1eRGc+/Iml2d/RFTl21q
mzj+SM0pGNi2t7EmBaF9v9apzeWXOWpah42XXNl8IOntfFqTb7qjsaGP9XT+HsEi
fqdwyLRxRO+IAOz0RMSeSpnxa0DfEF+84cVyx7CAwbRIjc6ZB/vzq87nprpvQIor
N4moCDE5bP6c5a26rjxo2XBNdTUYRjDEJ+IBMmJZN4LuY6ECV2TGGHCslByRaycZ
T2tXpkoFyfVFO8tbePInVMj5Lpp5Fj0Q5+vBBFyFb/UPp90KXsoo83pKiaMKKGPR
GDhh3f7lJbmOabcjd83wQ5S1vDVNdxTTYWifI//TUYaOAe2PeW8x/Mj5iHx3b2uU
YXVsK9jnUKjC7x/nkzwMp5zz65j1LRE0KTZ6/uvoLzdeYPD9UYhz21jUlyEkDXPG
nJvya0t7gtynlVFppz4eiF0yrJrl13bpz57sWd8H77eVkCfIL6wIysIVSk2onoUK
hjDBB3QvbGlVf3J9FexogH3l9uTfNhPmpRUTSrdT5K5iinq5hVuM6T8F6zxQLdXI
OdP4LuW5X8h1DOqFB0JzLVsCnPq24LEkQ56phdVOrJ5Bci32WkqMRXXuZLZhrR/d
AID/Ka8aJYJfGhVCEJVGuxMtn+/Wt5RtzyL6PO2j6gYZ4KNmbf8ohIydJFErC5le
xum+n/zOc0shJgAXw9Zu6WIVnlddFCZzOlnK3SDVyf7XVnGg+peM8LdwgEpeU1rG
Hp52fPzSiTTJmPBu1HrL3OBmXZMZ1ZBOUe8pjs5BYF3nmA0CTIgT3i575xvS2qgl
Zb1y6H9hfDqKEvcM8a2dPgOubGZHcFtdesBjhP9G7/V9CEAVZS69nDhxFdNhCK6F
QRBre7BOyeMKq+52nKKpxVgDofMoRTRnEmLbevrSnHUWAgLXPd18b2nULDohqB9b
K6qYzOadOFAO4ZEsGo7lCh2XKnkVZgNJL5LUQFaOkFBjNLf+W1u0HEJDAlMJIzov
7bU+uE8RzDScKaBjqtZzKiXdxOk/x+CMNsiOFjBMdRLCJH7idq6iFxgBPzkhP99h
AuLvYSAh+afyXOoTjwVj/uEc/KmfzXKD8BUln9xniAwlu/xVvTMDPWIW37gURwY7
U6+4sErNg7NYTo/f/4Zfe6AZhKo88XhNo9wzb0cnsW+UD0EkuOpJZq/iRAabboRu
CjgbkelYpCXkbZKC2oLXFMAAOvAe0HHyjMkt9ucIc/ABEAnFHSRqAQqYy9JFXpMr
FtXWjlsxWfZdOi03EWQXsnZ+IenzaVxxueArPjgEkFYvcGjrMLpNbffzmndqutFg
gEhaCqLDv3EtkdFPyPR10i6ha8+ALjgqQDa5w8kfAyTiDAd+kQlgTSAN5vKzf2l6
cKsAAHCt2t1mghT+tkQxkBUgiOpvXsV6V2v6AGBpqIsB1FHXWSml96xehp/xQaHw
7hK7HzpiacvG4feYw23QPi8iGWiADDqqijLsbOQRXzmw5e6zLO2zwnKGwTmtA15V
CGrqJ8PjebfOQ+yJtP78YS58GDL4Y8abwkDWUj6bF1Aw5gnCfX4PENC1QWfgH1Cz
wVa8oUw983PMhevyb45MO/Uqjui1pwNxFkorskSY7Gft0HmN6my27OmRFfcNkJUg
uhgHqUiuJ0zAwjWHSH/eJzXDhVJuVigRDG5QPjQcL2chcP1fS+hJyaBvn6QZ3ZSZ
YKo+pM+FgBcgKIDyAk9PzJXmW6weqhG/Il7X3AJeAuneEv/oRa+BMYrsn/Z8JnA9
zWm0h3IjV1EWJUAN0/DYmIEosXqaSkOQfzRwG1LNAtrTdu+/vYdp3bwG+qGZ2Fx1
pejJfyp4+sq+iQuL1nr5SVI1K82ySwnme20ui4x3jGqNPMC7h0fXTuFcIigvzAyy
MjnhODEDWhUTXiHNlMTKD6ne+CMGyEMv/C8osLvYulj6s3hLJz4Bwsv+7raH49FI
9CFOPEeViZIKFdRJv6nHhVGOSlt0q5BmEQgewRsF39HvIgcTpUvTZoHdu8sHoivW
dMblZtPRaRhgenlhbj4ftd7S5PYrpsrPx4qsfQghUSIXeCgEfgHrSLov+03J7KJM
6Tewyemte1TesaYWsRXvTVF5+y756o5qCBGZhoUrxjyh5AZ8f4nHcip6MttulJoI
+io0j/fRjgFgJz/8y/LbyaDW5e+97DwYDq3bRzYrNV3hVECve18XbjddkaTMUd4T
rRZj+/uE7zK10Uw0+NwKyhNC4rC9IxKHkwAORv1vsHYWSPxN45dq3p924LAPfgCS
d/3PyhJTUCvLheMt9aTeYWMsNIXmDe7VXMn1w6tKYm2aJ1dpaJian56iUeokRNG0
gxjWG6MF/7TfMBeVIPY0V3qHazMcc6fYMYmfNgEjlhtG2egiRjQ1c4dO58/FHF5T
rQwaQaYaYqpP3ZYOpn1Oy8mQ/ltZ79dOER8ElGBt7qVNFNjmt2r22TXngAdY9z3k
Rz0/J6UxG4/8SxI65ifOGhBZ7vA9YbD7c06teZMB2EpvGi10kWwY9lujoGNtJb2C
ooiyg4vCe41pd3fHZ/bg6dFO67MR3IaDYBWJ0JMqrtxakoW1i9qF0ncl/P0R+N3/
cJ0Yjh1s5sDZk0cPffVuTprTgJSuY8a91Ndom9HYE3rApiYrd9XAzSl2iSUGe31M
X2jNr0tjWMfG4KS1r3Ev2N08sgzxBuEm4BCFohrpH6dnRzpcriVIze6PME3itbtY
OsUN8I2k8NZwOjQhKTLMvWxeMJHbvYDZHBFbowMV9Adnq08P0ekQpo6PoLcUyLes
g1xAFrr85Urq4E7Pn9N9OPeCinpmD0w67jcj1KnXc9RJ+X2FO6bQ7rAgTCiI3B/w
GxZhDTJy/uScXa6lo5+Kvf79kP2iWfyqlCBQiqtjMmvHNBRTWLeZevCn6VPE28qa
hb0lJFOnDijl17Yc4NmpOhNz1T79QmPHMqEsVU1bY1UyRLBgxVtB0+2PEGmvdnr6
mMkbDHD7vqUeKq7f+t0LV2Nv+RWaUjcpyEI9Nglk/SZkXroVH9Y1TzeawqXNxVMO
ChQuSE3g9TAaR2bGOyvn/tcAyNBQvo3iwXtkD0zz3kKfvpVvABXrefiTEIC7rw3o
qhKIzKQfMyVE2rjf4X9om6tjRTq02kQKi0ooQA6I8C8mPcmC2S+bDgEKPZ2oyWMY
AqmPmOwetsSundzNvo8sXHQ9zS1r/qE6ArKrPNHm8CGGygfuJjiv83M8kfzAmzy4
VYukhQzmBXHbQNZXlSrvqnnav/dchIr3CCtQ6xIy3/MOrfN+lGuSCQcxdzAypVFr
nNVkI3oRN2HeCWNffzdks9olYdUM93WGhVzbPTvQUJhVumwVKOANmJdRP8Lk+BbJ
9y1O93fp8XIEA6K9MBA24GRI4ZOriJw9dq4MgYA+vLAx82ZCg6g+877k7z2So5eN
n8JOhGvO+zonCW62GGz0FGbPdBsOf2GjnDHUxFdtltFO4zXOwavaz50D/JvxI5L2
JEhVywCsXVMxNTI9YSC2MniQXztgHBLc4cWanZDQMUfLAnQwhmTF7QZKgSErBxMb
AubkYA6JsAO+/tlMrO7SwD62+C+jr5aySjcxQtcN9QxtNNUQzDm4Z3dvLiRA432j
CxI1fSd94N07Sb58XchNxwHkaIsaH95LvN3KvAd2ZBlc5NWKl+AJxAFrFDLP8BKw
wA8UlxNwCGOq9GyR2okPanbfY0v1SDJM1kbJWsFWEoxNE95vwVyFBayxV0U6tZnn
zV5Wkxi90OnFYn3etmCMEEXXS0uMOUGv34d7wqNYi/mIgcaavDCn/ZC5eaVDmcvJ
vctexeaojaISkUibNE5vE7+1wDtGyDUfNU2uP6XX3yd6+GQ2SY5nIwkkQT2ZaLMj
l4C0DRaEJCpTAhuSFzfQz4MIUHw8bW41heRBn1U7ZIe+NybnapenAJKrlCpoVipt
B7Cx9PNM8DjmK4EGY8qsF2bMNYJHxzc4ZfXF6LmGaDfTygL53j5stv2LNx5Syly3
zEkOL4sUrdAr2PR4cAMOwKRoXR2IgEhYilcI/P9OEY1y29hKLrVRx3RL/Hk176zQ
QDRSzUIafsQY+0mGJW5b35XayEncLUIKYGmjIWCl1SpyCvx/rs5vRwhIdsL/7GJk
1Xx0Liz7brlyRMFkbyqFSgloGHaSaszDG4nuKLkIUUsuvyv+P26GfBexgsp/Pjnp
+7l6Lk+XCyMr5K5TQfLIsRSLi/T+zlfjqeI1ZLaJ7WCR0EEW0X3djv0v21c8MoHu
2X+CnFzlTYJjBrjhrVTOUDH3KLaAx2G7Kvk2bNDliyeF1gh5Nqk4MzhfqbYeY1BX
xyXaqq4eu3slSHwz6sSQ4vSAgUhB9fdgwj+WwkcktZ4Jd/BpMAJw6fI/1drZjvf/
0Qbyt+w/3AuUBAfnlmUVwVW3kYhTW9wPtkTyj75EiYR0sWiyWIpjTkO6Mhi7fq2X
i4WVDzFJUb+FWbiR+c7xXQ==
`pragma protect end_protected

//opening this macro for dvt support
`define SVT_AHB_BUS_MON_MP_CB_SIGNAL(signal_name) \
   ahb_if_bus_mon_mp.ahb_monitor_cb.signal_name``_bus
     
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
QVm9BdgfNL8szriyMKCLROnkD0Qm0XTGLNs6/EB/ietU43OmydKHKmEOmZvHQfhI
iMd4pyjYF1vnUCZZpNeQgxk3upsMQ4rMcizFavciHs/5mPDcll+xXcm3s0SoNNDX
fnQmFa+qgcRCUk5MgucpTJi6QeYZB6ElguIuNxM3tss=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6017      )
gTVMij1o6FP6qqkTExq/JWYg6hDpPkLDt5KreH//127/a8rgmjSEobONrd5i2Xw8
jh3APC4whiDBfKnyg4pyWloymOUjOHfO5JZKbJ+UUDdyH9QR0mE07MfB7deYB+Rj
A8wb4rRqYw4kKp6NHUWyOl5rL+7v223WVHk3Q+EDtUGw61DWjufM3I6heVMPB96h
oT+4dPJpgDISTgaLTv7Z5WTmRPpgXb8pvo+iF1s0EFAjLn1l/zdSk+DRMxXek5xp
PsZluTvZZSetLT96RKdBzwCx58UqYiiO4foI7XEg8H26XMEwufOS6Xq+Kga1TBPY
LB6QbXfaMUohptYj6dvWr3heyekZULnZalsyFKG+m4pxVEH7icNzDtAT5sen3P4a
Bgm6yPbht5zILroFjzdraVnFhrHJKoMCQhpBPE3JNrGlLzT8DHuAYfrcNM8Xp4TZ
yhpGww4i+HItsZj6WdUDFF5efdb5fMlHljByw3aJue2FIz6/0hAhNbOis41JPIFO
U1/BYkhLgIOAseKqT6NrhYMVCAvbSOIzlwMg4u2JcQhLJDWP0ky/ZuBU3VR/0ol6
WjCmWmgn0yjRAj2gxt9KfmvAbHmMyGRRv5Chly4vB5jod6GrWK25MImB9LnKCR/4
onozjfw3BodlCvUYFqLkjpV/72WZV1s5VYJBYybmSVUfJuPMDaWYGenKDldZREdH
fTyQsI00QrCUSLYvYBmEien06YgVrnjSwI9RJuZJ5G6LW3eubdxn4SzVDrVnMYN6
JyPEP/hYPtHQO00e6DTzcDkvsQKoKgj8OeN8bMO9QunTxDef6ZkqCawNqRr83vBL
Zi76kwe4oLfPSxRfm0KLIwlO5w0OqSisWsaeMkUscTPyamHuDk+vyz4Cl4yr3QGn
RvLZtdEgGJu0soGw6dAxxl0dnM8IzAa/zxVM68Vs6V2uDgxnB9MMrOiO7fXxMV/i
ct8ek2O59ISfRV7VvTiJKWCJOYW6ZcU0wA2R2Jm4ht9Un9yDylDpsA0GbavDrefR
7bhq8VyTm0nfuoR2OSgv7qa6u+M5qe9KP+rnkgueoFUrTcpvlgesmf6UBfLZ8rIW
AOdhL/tkCW1xg0Y5Yl0GP8CnsET8ZS8gwWDTPWaDagQrIOmTuKRP11InVH0gSq9Z
BTzvZ0Q6ZtwKZQP9/XjVSnbL7fEvRsy5tJwmZvwbMU/sQjUsSgRHva24chgc8vHJ
8X60S0qzBtrK7nMKk5JYzHD9Zq2rixICWRpSFzB0RL4gmseGoJPhcU6QZ9f8Ny5C
8gOaTHgelOCHlVlBYZoTMN+4WmB7mfwMYZagCo3ddat72HAw3BsdDD1I+twusv6D
d0+j+JW0dUrnxCib8kWjYDOSW9DTwMTmdLw7k7vUzil/79JqG11rtyIW1Bu+xNeP
Hhk4yLbTR4UUw6yjtzxeRKQSYqC5L6+3TQomhfmuDf+VRMzjU1PrWUAE/nJVWWgo
LH7RbMY09Nsr/Xugs/5M3ow2tDSQUO0CWz9W5TOctaXBybfb6j5tJHZ+ZOKYjj+f
A3EFzR8fux+KPFrqjr4sJigC+3mHiEnLh985tQSp0sXy6/wgR1NDF2J+1QDXPpRM
PTPzTtduwGdX9+3r7EUCEmZw5FwGAv61c6CAKtWtHOyfydXA3AKkUKgqpM0Vp5EJ
BDLwaFRpWlRt/9+Yq3FPj1LMvgb2g7FUQQ7WMekGWBl8WyYY2hKhvpyO5ifsUP8d
fz2kx/fuFtLeKx/ZSOQG8du4thz3AgHoNowGGlBuDqIeF1G+2Mz6Uf5Y+zwpFpea
0XdhxMMQIQOcwR/c75ZoSgTCplktTievKpjqDlC87ScJXlMErf8qEaFxOzOeYFKY
wwPLqdfTOY1slyj6vmAdjQTlvhqnsj9xQfbe9orvwM5wGHNptXcK2Rx6jRO/dyeU
vCdttiOPXupvckqSRCDCrCz9vEwf/7QV8DbNdJlhcsanUsJkibRETcvupzoxqiqV
yeoEqy42QeTGszPz4md3TdsvPTZ95N8h/wnYUkRN+KdzG0Yvxai0fZoKn+DuEavZ
c/A1PvAvY6ype9gQHbNLs+ak06yle31O8SbootU4OnB31ihZXvoIxqKPXYPoABhs
BqLGiwbbtDa9tqmdNgbzViava1/M/f05op1Q8qVZq27PqD+tuiVH4eLmhOannBY7
P/521DV67s4Tz2Wcq5DfdJT4UjTYpUGqeF2kvUF9p+WphFABwT0WGSJk997OGs37
HznjyF6qmh2Vye2KM+0u1oAmSTZTw3hOTcDdsdEvc8y9jG+aLMza3wOWsL95THHR
yynixxYgNbLVW6NJzuYpNJTn7orMZ7POaTZBs0BGk51PMvA1LK43rY7KVY1xNH8M
7qVxsLHxPMWsBvM4Hj2DARapJtiKigFBE+uS6ndRRyRjSlD4c5syw+9kdFgs544U
aZzDrQ0ds0WhKAXIkosHVNkIl5HJ8AgkJ8qkcZn0KfeMa5dWCE8UZ4p7xJ05/5v9
3ocKl9UHGb8FVtIEfBfTnPlP8d8CJSYr/lUwDKW+PVfOCTwt8y6CVL+TK5TcZEzz
goHRzM51fV5RYMEJRzyacpp4tr93wAWqHommhGCRCK78VmUYeqrOQSAAzSPwvnmW
wtt9mELHyZULhqLtpwkuHAhrB+5vHEwJIpazvu4w9VaEbOWpOGDfdSDSJW4Mlsq8
joBvhxdonq5j+pUVk7EnF8QA8JAh5iVhgOzsF1lI3f0+GGhJ3KhONHgiNzj2oBEU
3tlCChDnnypcOugCmG3DPxgCskdT24xHpduXJ7bGLfMqtTGcLdQPDLtljIlGUXxA
poQBzOwXRdVs/r++QWGXSquhs2va1UjDgekHZN+a7HD2Z2S75Jp0eBzc/xKFKHrn
izX4UN180jSAlWjICcaf7yZsbz7Lu9nPFw8FstkotiKWDeMhsgTZOeT897ucD8ZP
C0dkaJbNi4qssVOvwvMO75fh6XoVkp6RogpR4hdYbYHfqYE+D9Q87XfrlrVgsr7O
GcgLkpyz34Jjywsszl9ysRTTpldxhTekU0nK8Vf7ZZ/ocXHVp9o08LX52ltlJMo9
a3oFl6x0hHW54tJMNtJXosnJdYtIlGkHikIHnxmWizgPkV/eKGejZFkpj2m16yGz
H6pqu883PNXzjTFV3RMUMT/NFM/Pizwe8cjtJpa/hymSY7tUtVkYr+cSdCPwRDTK
evb87W/ROKssCYwqvxTBaeoFSDHLvlO3Ym2mFlTVOqJH2wAS3lnykEOA9XEbWZXC
MiByPrlkb5HvhdlVgjkmEHrkR5lMfb+7HktbnGNc8eAsVA4nQpc12dB/Q2qZiPzt
SQ6M9GAF3t72CkpYf0mwoS0YEwgBysjiaofz7Ny8vg3jrckdhe+L6SSaJSzwMHdz
XUPcGuUca5bTGxB7ePdEZThw8Qm3ClMI5HXAce6IqWEq7qs3IsxLFBiTynG8tGm4
LMO1KimlEHepIIyFcYQhmh9hBxgR4NAvhn4bwohjPtGM5qDHRruNk50fE2o1wWY3
MPLPGkLDawpl/6FKzXQXjg==
`pragma protect end_protected
  
/** @cond PRIVATE */
  
class svt_ahb_arbiter_common;

`ifndef __SVDOC__
  typedef virtual svt_ahb_if.svt_ahb_bus_modport AHB_IF_BUS_MP;
  typedef virtual svt_ahb_if.svt_ahb_debug_modport AHB_IF_BUS_DBG_MP;
  typedef virtual svt_ahb_if.svt_ahb_monitor_modport AHB_IF_BUS_MON_MP;
  typedef virtual svt_ahb_master_if.svt_ahb_bus_modport AHB_MASTER_IF_BUS_MP;
  typedef virtual svt_ahb_slave_if.svt_ahb_bus_modport AHB_SLAVE_IF_BUS_MP;
  protected AHB_IF_BUS_MP ahb_if_bus_mp;
  protected AHB_IF_BUS_DBG_MP ahb_if_bus_dbg_mp;
  protected AHB_IF_BUS_MON_MP ahb_if_bus_mon_mp;
  protected AHB_MASTER_IF_BUS_MP master_if_bus_mp[*];
  protected AHB_SLAVE_IF_BUS_MP slave_if_bus_mp[*];
`endif  
  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  svt_ahb_arbiter arbiter;
  

  /** Report/log object */
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_log log;
`else
  protected `SVT_XVM(report_object) reporter; 
`endif

 /** Handle to the checker class */
//  svt_ahb_checker checks;

 // ****************************************************************************
 // Protected Data Properties
 // ****************************************************************************

 /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /**
   * Flag which indicats that the address phase is active.
   */
  protected bit address_phase_active = 0;

  /**
   * Flag which indicats that the data phase is active.
   */
  protected bit data_phase_active;

  /** Event that is triggered when the reset event is detected */
  protected event reset_asserted;
  
  /** Flag that indicates that a reset condition is currently asserted. */
  protected bit reset_active = 1;

  /** Flag that indicates that at least one reset event has been observed. */
  protected bit first_reset_observed = 0;

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
WHaGEwMpFCQ4ujA2/tqbgTVDBMWg02fYgSrFxWgXr4JVHFY60Rr6+Z2xDt5wI97X
jcFBzv8ernOyn0GR5E4ihLsFVMh/sh7zQ3dUrOGJV0m00GsXCitM1IAcz682hhZi
qJ1GigY4FDhEhE30V7LRYFEoBij9xbgVLS3Q2Bu55Os=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6138      )
000xDCH30grEG1YUReJ9BroLx1hBK71L0BjJj9KWCGbqoYd17/+C6/+/pmq5+UwM
H9AWEpmURF16BY4mOhru3Rnz7hA6UYTS+XjQinALlXaM4aiHwS/xknOtxnjfg0ai
O7mre441QsFA5w2hTWXj6n9yWMz/EW96njORnOf3CBg=
`pragma protect end_protected  
  /** Flag that indicates that the dummy master is granted */
  protected bit dummy_master_granted = 0;

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
b3ufKc2dqBrXYcEUz3CRvSo7sa2qQVGGRoMlyzeWXBXehGJ2EGYu7FMOogRgaNpp
egw0sOyrOxwj0WQHYBUDVmR43x8crw2BDgNAkicsA6PtXAQNBXvuz4rcsxWTAdy8
sKbvP5Elzlcd6nJJFQxE+9z2HsFkay4el5RGkJhy/U8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6259      )
E7IfpaMoWq7t/7ybLEL7oezqEaYxoEGuIHRccRaCNH9eUgXE9kCGP8T4ZhhR97vJ
0ie6BQSIS70cxKA9z5MAv/FIiNBzDTIzY5KuWEhNuLvNOo4WWoSVGHtjap2wrHKu
8YsYWJFiElNGE5KF2v7R+FZuPnghJQgsAaWlsaQWKV4=
`pragma protect end_protected  
  /** Flag that indicates that the default master is granted */
  protected bit default_master_granted = 0;

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
olOu2PIMLUIF/KQjTi6a/7Vc9QYfTClCMK+CfQ2n4PAMX6W7+RQBeI74KZWFlk35
xJku9EuDRqB8QAB4CHgHgEdwW3PS2g15+3rWRTmjiNusBhkHLrBSP2JqQlnAvQT+
jkUG1ZyUA91cJaz9GWrc4/N1VcSLUkI2Ih0x8MeB/KI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6380      )
SEf1Ir1pDglcnD35wAS5P5JzChNSxKzmMg8U2m0z2seRwLKCm6W0QKUirqi338C9
qIG8U27eFuJSsqkiplrM3YyQTeAJ04jsgn/tWVRpymQiL9rHzf3Rvb7JQu/v6IIl
c+ahcGt6KxKndXfBv+jujPv611QV01boUdQQygmReLE=
`pragma protect end_protected  
  /** Holds the sampled values of hbusreq from all masters */
  protected bit hbusreq_sampled_value[`SVT_AHB_MAX_NUM_MASTERS];

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
GpgZF54LGBzJnZJEMlWwSrtLN3ay+gyy8Uhi80GuFo/UPABBGKXaiiuvhZ8mGyWP
4SKbaN+MXDz3GxQEFAtFY16sg2SATjig1BHOiqBh9GYmTexGdcKJ9a0GfVfXx5Jc
nyhj0y20AnQOV7uqt6oonq7uAQ2FypAyEP+VflP58HU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6501      )
eFyLsbxm8m7JN1fFN5v1pIc2NjEjYX+R5ODfqIXWdeY2+XDrxhkQ7TYsfKqydDSZ
OqLYAgmlDZGPGNP3zYAER1PQCsXLN55Ah8n2S4ISRGZLDxQijANFx2QDYWvUO5nc
AWA9gL/XkTbOrUjDVIW0v9g96kaJdN9Eqv5dwtRD8c4=
`pragma protect end_protected  
  /** Holds the sampled values of hsplit from all slaves */
`ifdef SVT_AHB_MAX_NUM_SLAVES_0  
  protected bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsplit_sampled_value[1];
`else  
  protected bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsplit_sampled_value[`SVT_AHB_MAX_NUM_SLAVES];
`endif  

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
O0yzGSEmPfHxuuRu63zceViyZoyoUw1L2HP9doo1//YCV5q8s6kb0EgpWGZq1L3p
+VwWKcZ2wm6kksy/0/pFSX1aFQoPmBUvTYWGrzuXG7AiAflTO6t8874xb3RWlfGl
2MrLP6MdMIHwU4NnDmtM+7bS8Gg/pH8Wv9uIgxEbsvY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6622      )
Ho+qFuJHyCaEMhr78GubcnB6nXHfRQaPPckdqr/TpH9pP70EsrKPkPSh/XoBR+Dn
BlshT9pwEAxIrGz1ME5CKUqmBGxO0YiuWHxm5aRlpFCb+8wmRLJubFyTbTYAa0th
rp9c+JtSwMW+glQX94WZXHrE0YXTFXvby7jUdhImK98=
`pragma protect end_protected  
  /** Holds OR'ed value of hsplit from all slaves */
  protected bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] consolidated_hsplit_sampled_value;
  
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
kMhpPbOHw4bNC8B885oTCtayeXUhznMLfIuFRwTZFsg/9+58EpGGhSXPc8LtLURK
X+1N4ZN1rZ7QwnCODM4gQdjgflBsOvG7AFeOtfbPUESsaUqRBKbL63Pb/bWqQOej
KvQstjE7UYSCgAf6/6wL/i6+KQXhN2TYDxi1tA6uLho=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6743      )
LH6+ipOPtMtQMqC91JQHFS7Wr62P3DvzpNgNqMYTkjAepgrykSCRDt4TWVG72MTI
6AOmZkJN3YFTdvGW8TdNDxO0hcv4eLdnexqYqJO7QUb+4FggsiRp1mojEXIGUX41
skMtOKcCuA1BGljpczHAzUHE1Vn1iaLaCufbAzPYmgk=
`pragma protect end_protected  
  /** Holds if a given master has an active split pending so that the master can be out of arbitration */
  protected bit is_split_active[`SVT_AHB_MAX_NUM_MASTERS];

  /** Holds the expired count of the cycles before EBT event for a given master */
  protected int num_expired_ebt_cycles[`SVT_AHB_MAX_NUM_MASTERS];

  /** Holds if a given master has the grant maksed due to an EBT event so that the master needs to be out of arbitration */
  protected bit is_mask_grant_active[`SVT_AHB_MAX_NUM_MASTERS];

  /** Event that indicates that tracking of hsplit from all slaves is done before the arbitration */
  protected event hsplit_tracking_done;
 
  /** Bit that identifies if the transaction is a locked transaction */
  protected bit identified_lock_transaction =0;

  /** Bit that makes sure that dummy master is granted the bus after
   * SPLIT response to locked transaction is seen
   * locked SPLIT. 
   */
  protected bit give_grant_to_dummy_master =0;

  /** Stores the master number performing locked transfer */ 
  protected int master_pending_lock_transfer;

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
QD8RxbLgD8eO5vOysgI0evbXfd6gVKZ1Ug+sj2tz0ZHarSTeuKfCwEsbUSFzxk6l
ilcxE7sUbhdJa3/WI49g5ymBVJ8qGC/kl5NcqcOlnuHntGbMx7kKlAVLxYPtIQcK
sK9F/3IJ9Xc52UHwWBemwQBQuapoo3u6seV5xcoNx7o=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6864      )
9e1Hok0exHOUJWJ/8cMfSAaxcSXBG6EUNJzfvyzGKBa3WkzMRdeJIyJf4hnX6WHx
T32zZKOx3+bIFmwweDQbgp43kAni2clk5nSS50crvVhWHCX6NtH8N1/Xqmf+EIVL
dD4AtEci4GRtBqcrbsWnu3AGSU6IoA6tQiwpJWMiuco=
`pragma protect end_protected  
   /** Indicates if currently granted master driven addr, ctrl info is valid*/
  protected bit granted_master_addr_ctrl_info_valid = 1;

  /** Flag to control the muxing of addr, ctrl info */
  protected bit continue_addr_ctrl_muxing = 0;

  /** Flag to control the muxing of write data */
  protected bit continue_write_data_muxing = 0;

  /** Flag that indicates that bus master is identified */
  protected bit identified_bus_master = 0;

  /** Event that is triggered when the posedge of hclk is detected */
  protected event clock_edge_detected;

 // ****************************************************************************
 // Local Data Properties
 // ****************************************************************************
  /** Configuration */
  local svt_ahb_bus_configuration bus_cfg;

  /** BUS info */
  svt_ahb_bus_status bus_status;
  
  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_ahb_bus_configuration cfg, svt_ahb_arbiter arbiter, svt_ahb_bus_status bus_status);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter report object used for messaging
   */
  extern function new (svt_ahb_bus_configuration cfg, `SVT_XVM(report_object) reporter, svt_ahb_arbiter arbiter, svt_ahb_bus_status bus_status);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Monitor the reset signal */
  extern virtual task sample_common_phase_signals();

  /**
   * Method that is called when reset is detected to allow components to clean up
   * internal flags.
   */
  extern virtual task update_on_reset();

  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();

  /** Method that implements dummy master functionality */
  extern virtual task grant_dummy_master();
   
  /** Method that resets bus info */
  extern virtual task reset_bus_status();
  
  /** Initializes signals to default values */
  extern virtual task initialize_signals();

  /** Drive default values to control signals */
  extern virtual task drive_default_control_values();

  /** Identify next bus master */
  extern virtual task identify_bus_master();

  /** Track hsplit from the slaves */
  extern virtual task track_hsplit_from_slaves();
  
  /** Check validity of address, control info from granted master */
  extern virtual task check_validity_of_addr_ctrl_info();

  /** Pass on address, control info from granted master to all slaves */
  extern virtual task multiplex_addr_ctrl_info_to_slaves();
    
  /** Pass on write data from previously granted master to all slaves */
  extern virtual task multiplex_write_data_to_slaves();

  /** Drive default values to data signals */
  extern virtual task drive_default_data_values();

  /** Drive write data to all slaves */
  extern virtual task drive_write_data(logic [1023:0] write_data);  
  
  /** Wait to identify next bus master */
  extern virtual task wait_to_identify_next_bus_master(bit wait_for_hclk_before_proceeding = 1);

  /** Returns the burst length, burst type */
  extern virtual task get_burst_info(output int burst_length, output svt_ahb_transaction::burst_type_enum burst_type);

  /** Tracks the num_mask_grant_cycles_after_ebt for the master that received EBT */
  extern virtual task track_mask_grant_cycles(int master_id);
  
endclass


//----------------------------------------------------------------------------

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
UgtKorr/fyVZpr9TF93fcBZk6Mn/KxhufL/DDLpqrzfGITx0szia8bcN2UkCFr0S
hz/zqEkcVbUOMZvG8pmixDyegS9nFaXXjrGehyJezSOO7JETa0EdKB16HNpsl65k
gCqtVSNsQI2IVdqIdA0g6DdPx2O3DPX2OqN0NWGPr8Y=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 7446      )
zOxmrt6x75oC3YAjUDgQMIuSROpepHefY22AiXMnUs9+87YqrQ7iGWC3pOJaQWuF
PhFVk4yPjAkr1Wyixeoi64yHv71RVooaXphP2wJrUNgGaISV5TxbhahiJ3GD+Ltb
i2je4pLsXEcKlPTFAh24Dv17nTbo09rgYeYGLWHj6YHVyInLADpWkhBirF2jGOMv
jxsPslLTXsDId/rifMjFDz5qZVKXbw7/k4Vxebt2HvwLjSlCXj8tOqdzNBJQZrqd
NCs4U5cAdYjKhvs6GmwVLPh5xLNw0/kPc3eW4cnS7fvc4YGPouVbL4Xib1NUuYzm
h1y1xWH8sjGTdN8zCfLiTJUn+5NmPfBZ7ewQtsK4BNg4mz44hmgH13aAxsHjueGW
Zs7ePetoqb4yYtr7PUbEjEt/e4dDoO7THIk4oDS7BR0EpZgy30TFOdK23buzG6Lm
DS1XPqOCh6fia5/MXUreWBP+mEHD/gJtT/hL+itx64Ced4ljE1BrDHt7So0tPMmd
Mevq9xvLWWjnTkArwRFXOpjA/p0yj5RNEYFsxoo64cTcagV86/Nh3DGTTqe8h1Nl
RsH1cTakf972adLakRu2PxkAYHdckPnxp0iDtRlzMOMFV5gFHtugGBNhuVb2w0ck
OxzZpoMHtYa0pBBj1STy2BEg1U+WRbs1w+nTuZi8qsVEXpmOFHedwSnElGwAXSdn
mUgIzhAjvT+V46aqpvQ1T+ZKQX/vB637QllQcVLZXiMRppZYimC3tjgtpzcxdfwH
BJu9a9zlYv6z5/9Hr8fl6A==
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ItnjGAC3R5ITkdloVDF9SA7+n+makvJwn8ZjwJUDQog/4lHgG9VkKFX0Bkrt/f+9
Nxj31JKUw/FmGvzv4nfBTogpZxtGym4ZH76XPE2K5hD0ZzMl7lYk7YG/lDcSkxXb
AR4qzVcIhio6bOCfFxqQGoDwVm1/RBVrdiR2d9IeJOc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 15692     )
djvZDjU1IF7uT3QMaYfI9K5V5LJSym3jModG/x/qrK81vxdKgm8pfEYMRCnZSol3
buz/eO+loEW4RgzI9GKd827K41g6Xi4Umg2cUavldscTUyaJ0KU8i/HYr128FCdr
dSUvL4PLrwCVTApBIDzEMMd6KUwfpNVLRqHQKmFjfxFy1XyVqvSiBg+/x6owIM9Y
3uEksLbPNvq8kT/3MSM70bSj4qbO+1xQtIPpbc3vZOlkWANROef5Km/dGu77rIfL
ABfszO7LJiqfKlcqYYKZwEt0K+uBMWhgeVvjjKv/lBGBMEE7+nDC9h/deRh+Ks2G
9JnQMnV7653SG2Gir6tE7vKVaJKcnP7CI/nlkqh1ZertF0AWBN12KHddm5WHPVud
jhibrnYrp9WWQZyJigqJhYhoEik9hd7yOpb1VaV3K3IFm3g9k+f6xg5Z0AuKiOV0
6d9asAuoMBILDzbouAgUWufP1XzrmDNTN5mguQA3PnKxhfaM1mqhX5RIpr0o1JBH
bhqti+TjYsib+m2CAabSvbclsjv3hmIccQvCGZLkW5t8yPTqj8XMf/jFofUPvKWB
bJVFZx3VNpiVM9i8tWBinuBeO7Vg4Pb/5B8v8AKKWuaVxN8cwKa3YpkdLixlfCkQ
BnlkO3rxiZf941ujUFYytImEdjgmBdnvwrAnGzDZZu0YpXIn8SmZuwC8ArAwNsbb
DEd67xdHvqMUGtUVgxGuzwelE/7XpL0MySN+w7MkpygffBtjYsbOvFFS1nfebwh2
pQS4VsyN4mogQbR+raXSP9LrHYy+Z9eA8jBTwOrTs30Uvzkx/7G2uWEuB/fjUokv
1FiMVu+nYTvjwNZtBXRXUk9AjNWjeePvU5nUXVTJ1q2+AYi4jPAfNOrb6jIYtPMW
fj2fBUYqu1zvKPMI+Z63E3hfZ3PuKqNTa9x2IKBxPhL6kx3siOvfQ08J2mHW9PN6
TGZRGBntIEVu4ihE2GuVp6fMWiaIjVSGpiT3qNEreG3fvubVogRNjfyxEXUfmKgi
efFl3U9ekKu5ViFxmeMpzavan1vGoiNaxWkikIAgJnsIW2RXQZnV7gHAf5TCijDK
tkwg5PMg4ppcXdcVRyGribLGqKRdZ7PDEE4jwPjiiDbgfQzSx5jT10zuvuJTWdfV
MuDmUuu8rHLAsBlO/aBqKd77/7cesJIT0UR5aLabeSL+MRffMa58r0qejFnQlByO
xV3oZ+qpUYBdumgwIEMvIF4sZwGpeF5yC6VHEfVlWIoZ1zTNtf8/Zb1xuVs4Rbwx
BDdmPLGcM4wqzNqaBGMBKidAMDycv877YW+TcP65scE+iGyAVb3ZagliFsZzMTSR
ve++JfES3Q0bStK9xeUDmrH1EdOsBmv0ljNx9Hq8tkowqMI1yFpz12SqBPONdOKS
WxQM9owzyMmnHmup2BY0DWMdc78liSJBidWTQ0EHV62zpDeCzL0LWtqI1s/BL9bU
reilc3ve/aweX945bZ7EiNaiHZffFVp0iLu7nSXlMn2nMwZRWfpLZDRxFo5LKac/
r6l+4rGA5OROUtBZR9ZIAabRGa2MfLE8ueAFrAWb1JLXbL+ISG7gTB9+yd/dU5G9
gfHq1saQhrJnaFmDtieYzC/h+nAuX2+Cu7lfsCpOjVwUc7dMlOQlQPzQ0YMOsE1z
wpN/xUIbESMGC0oRby9wNdE3YxyZidSJzd/CG18SftKIHVqofO1lpiGM7/8R0DLE
HVC7E/aF9EDcVS5vZp/YyVd3mvmpXogUyh/zaCIykV3v2L2dxA674Gy4Mhzmchu6
EFug0hxL5DH6ITfd00/qZmeyyH0EhjY6IzWrYsSqvO0T8hlrBLlWvyThwF+ZJ1wk
uWzlSybUwChLF+TafcyUyXOeebBqQIOhsWLk/D/bPBMepRrZyZh5HRj/JpbDpiUn
tQFOzhnC4W05rJxb2xUEt/KVN1LZYBL5Oj565U0Hd7E2uy/IRrFr1jityXFgAs7t
2i1GhMVTdI33PLqiEZo0cA0fLDAkMAYMTCUwO+/QCrU/p6l6YKwYveGB6k4vQ/SX
xt6whuqsCP2nwLhfe2NR+rXSE1q9VwoB8E1GG+CUDkW6ut0jWzI97XFv1IaLoLy4
xfTGA3BbtwPXWiifZ52Q8mSu8w4HPlor+L3vgTTCqzEBL5pskzZxaC6BHFTvpBS7
pOE3ZNUtHGihWM0LW9aOTE211k8LFBj5i1N6pD1lpH2qvH2DNVcfoN8CTY9sxONI
vIGdyeCfvBvT9OXS+2wTpM6DrwAmXodLVDyDmKufwbKL+G+lJKbI6yKTUd6CTe/A
Q6ORayTNndHAIQ8Nlfc2KFXVlNt45te1rIKbMSzeWd8V6EvhAxW5PSZzbc9cvJVt
oI4n0k0nO7TVPsH1j8/0Thnw9X5FEQIHI/UpPUn0hcD9ceq1ILNvEfZPl7KcUxF6
UKgziHKjtDL0ZohWGt6utKd6afG4XCozbWhph61gIZOpmjBUcB7OYl9SHYimxU2h
+joKN42OT5tYIiuXM0916qQTMgaoNgR4QTEglewkUmO5QWXs+kdkg7pm3ghhRcpS
a1joND3ueLNpNgL6tdJ+1xFTux7kx5LW/c7NX8KmUeBdaNP97r/do7Ku1rAQv2mc
FMJgOeB6ddrnBbRNvcov8awSgpZPAXwLiKsSgdejzFL2Z9E3J1lHiw58G9Zrs4xp
C5qjeygdu/bGjrlPW4PAWlNvqnq9TASCBsB/lGfG8qvJ/bATd9OrEkKNDEOLoQVE
Ph5fYeoaa9CIRX5ecbGnoz1Bw4myTqRLN2eGc1J2Y44kS3rXhe/kTZBrvOfc9Clz
QxJo+a6D3xdlMG6eb91KZr59XszsXv6rPldfLzWacveePiZuUkoSdxmEaKEYbUGg
f8iSna54g8b7HfsRVRxhIPav4RSV2d0O3QaBQXzQyWuQM8/87SKLiWMSh1hE0TQc
TXjvM/VmDbRpB2vh5MZ7skq3S1uiS4jnr54kYKvGZXZhmETT/LRdyAeKp+n27F1o
54+svDBYzOXoNPMMsWeQ5rz+qf8/dr+1SfpF7pR4VRL49iysj1CBpzhRTPYSzBmM
dLFf8wUf0sc5vB9UxSqw+4bU+DCqfzCsddNY8zJvmftSqpfKtcC/fEK7HYJA+mfM
AxGvDTiDz2ccI0FubnNRmO2ae3r2peCffYSRcOd9eKyvk6m4LvoRdco7dcsqECt6
xoQmK+6LsT+ftYcZaDC1/yqmb4lGgzt/9HOmvdZdoqqz3QK+zK16mqKNIYVMWaUa
LJNEZ/ecUIec+plX2QVSOBE1jaDUS5L9/4AHv/5fC0vIrXoYzs7vCCjmtblytzC7
ogbUBUzp0qLqXPEAAFvWrpTcZiVQYeAj3knnziNF3fmI9vbNILfAl/6xyNjzU0Ag
ZtBbEBf8x0CMBQxkOFWg2sYo6M/LojatUVdPvlI0PtkmUS1nLIO51aAOXiyB4wly
ZdgPze08AxTseIi017EHeyZQ8DAQhE0MeVXdQqwGvtx0GmuCnqM2/eAY/jOO7beq
N6xgu9sSKozVsMO3V6dQmWAyZm3kLIa2KDd+P/5Kzoo5dvjijalaOyirytN98znq
barNQYeTnD48M4bbi4BmY5a4WP3DAjxPExy6ngR51CpKNpZLwwko7EQmp89iARSA
mw204Dg4a3ao1Gu62rvnkrmAXtTJ071DIxiPUW1dbi2FQrGT0z4MErlAAnszGZDj
c2LcV4PX3yP5AwuYreUe86yHM5RNgx5bRhMQl3V7GUln8/Sx7I0pTv8oAUESpBwk
pU2DlmU1+jq7HLUblcxvePQFRM07yWBINT9c3OG8WyfI9k1KNw0i1klR3Ty2DGSn
7hFy4PWmCN3Vi/5yYvKNLDs5rJAZKmzLSkZ1Y+mWKV33fLARNv/KkTAfiH1uhCPC
GFTqxuqtsHrgPPgzUU2RnXoHRq+MuDnME9oGVnFQgJRRJ5VcUQCBDjFvweBdzKz9
RjskYbMb+gomglxslMSCFnL6d6VbczMQalDnvkNUxVdRCL6VQ3QMv7Xejrz5JXRv
7ZNLb59IrGaiPCWNm+lJk4BKWEdq2K0YnNGGcCjU/f08qMq/YTJvSNDfOKqREiEp
iVuVKdOYzVStaF3Ry4uABXGcjD69EWGGr9M9rC+TsFlwtKYE9tTM/3ZZAyO76ADf
FzEWtKC+eS+sYG95qs1KiW/2ZsK2S5/6CAIQmyGJNb8I6KV2gZy5GyQI5Lz6Z7d+
EpMHNuMFlpJ5HGcVhNx6VZVaulaR7O5kEUnDBLJ2A3ZzUmrcojkhkZb+808icoBj
V+VI1VFInQCeikrRJG7zxBOjFDgRhPYji0ltzkCbd1Rfv9LDRTezqVE0000QyAbq
hkhIz6H333/zpL8//riW5lThDmT916OXfYsFmmEah0eE1r+xhJ6DUnnbltwetBUk
4zQhwbrSa57NWm2ClnHHkeULCbp5ijR0AyEYAtfXVxvGjyNpENjzG3g5v5hnxtw9
Y4FJZdVAF+/EDHKCJzM2fK1NkNUIkzy86wTJw4tCqVK6Q+PxkgIjKdkpszb4QdHq
tpf/gECAxNTxEaz3w8IG26MBUgA8unWb3BTdbhvIkiVoOhI5h8U/J9n5ldWTpYgV
kLyIvEPMwrYQIitwOhi9m45YDqAPxTMDBYRKYLQ9iZUO2+kAn2j7mD5CnUvW/WKb
qLEqJRnGT2Ftvv+wFD5CqrPm8nPZCagGN7GAChCxs2y+5nRoQCgz4p68zEz6fRHH
d7FT2Icw8FRrSEVmmR3igwCuuH+qoxxE+h7DQCc7uMB/c1cnXMMnbv00yH3ECv1E
mQtQoQDyOBXubnQ0yMnIcaKHDCjWjdjBqV+3lOpAv+w/FR6yg1wd6NzFq1hbPOHv
KlvGwXZjgkdWlaR/OLVLUtHsXozdqz2qCIFYVP3urMMJW2MlS9LxxufJItgkKiS9
pQbOpNqb/+EclpYM8AK6Z681kzXKao3gT+LxIgLVOstxhRXvN5dowD2RQUl38Fwu
Iwt3mM0LnNWu44GKLNLOzy7iHA40MjD0LJzCpEhmLy7x50+P074EFaKDhG6VcmY5
73VH3EQ9Lb+Fj7RxjLHaFmSr4c2ejcLK0pPNvMY2lvF2XFnBRsbJjhdPVynlJqOC
VArQYurwbWe2v4mkUR4OlWLmZv2lmCciUNvJ2NnxxdhMTjPZ4WANf8bjpMCXIcxq
od8qV9+Jgg137GuAGirx5IoyhplJK4bPCKn+IvJW2UzgNfjB2KWr4O88EeRbz+qs
GQEpNkYA5O2oSyJuPdTFNV8tfVrD/5afr3CuYZPLw0BmsWFsVR2UfW4zN0GxMjPp
zr03YpQQmiXioMEEF0LJt4xlChBksJNjbtLi0o9s+DAcn7JnLhfUFpXiq7jblh2x
PcDWkJz0ykeAe4wYW546Ln2oLeLf6lNk3+Z1AXsGhs5cheMAACiW2+88umTr7Per
dnRGmfknYPUER9CDXztLmdCbviO8CJCpKGExXqXNlvmwa3q1VSq/b1Ix2ehX6fiq
xL2SWXRVA1BAMbg3hvGDwd9SyxEDTm4gnWbBMHD5HVseX1O004eAId5/WVXEYWLs
X3Ee9RaEtFwle6IebtvfLMZGh/QNNSa2pHcj68AGpPsjJLp6v6Ssnht9phiqSaok
j+PGK+GheYRcQwVvh6uQM2EMWhKUjVqm0PXo+j8DFWfQHlsx/H6Og/nb0/q8h2LE
anGvXCkCk/kYfPX/1f1g7XNU+aIuXuIEZV2I5mT9VYsaBHhB/nQJ4+4MmzeoSwk5
UtxDW4aiYABrfk4e56uqnzUbpBg6FLxDl/FulfLM0Rvr1x7dVELC6ruzWGftDh4c
2bNHoC7U+Jjc5NMlDbVKz1QAvQ0t+FMhro4meJQLnimIQqA6UDerA0GZF80pq99E
z9uuPGydgyckeWpLxrd6jiG+T0Q4kUKF7I0yVMDYgCoCI93Q2Bd7YnWbrQRWFkVQ
EZLr+guXkRQf/lqtlIuJ1g9vHRHX1R8LLkQYoPRYsxXU/6du01hfPfmmxwF/+PqR
zbxm6rEWntEdqRt2n3ye9h/JWv1VsduwkB5Yn8T4wMHCZbxglouYoM2obvC+SilR
mR8uLMd2G6r41zBsC5ovm98d0l3KDXvmIaPITniW6wKE9E8QaKw51lfGi030OaIH
eDqVsDXQmCCUlzONdDPFc+n5i//D/bZ8tPAE4UOqdvApG/cWirSurl7kvOvAmz3z
FF8/xDoKOI/tb3Y5+FNccwgv5cJw2chwUaE+tmhMWSpkq16f3kmnoQ2Yd1dy3Jtd
H8NGpetsNR7tU3y0O1+5NeGx4nyBRkaYvagfwQV9x2hiYyfGGx5YiWvt7ts2sNzQ
M4DR6kFKbTj6tbmHS56ijdchtOxo6bOZr7PqnWuplk5aBUfeIWIqF2oofnjidTUH
m7zc5ix0HMCdLYg+L6/PGHhj06vcRUHV2qdFQBE8L3BaDBGdCtSIAEzJDrpDQdIG
aa69lq3WUazNpq0U9nyxBv8+5/DJ1Q+s2YkG72gz1IkA/5D8wOPoOBPo9DZeMIeJ
eI/YCrMysUTfR5/iwvXuWr675IL9BRnP224mhZ3ZlG/B/JwC55SjJTtHw9Q6q/Hz
1qGB/CK05w8FJiZqU5xkdmeyUJTBp/1NIpJNayM7Io8tTcvApPYa/dkwIf7f/lch
5kzzsMd9YLrhIVHV/YkHUyoYSBFfMnV/y/2Q5yB8zOkntS4GgAcWHFFFewsYn/Ts
6waAwFVdo86unsF9MJGOcrhp/7KHersZgTJ5R02PqjtbhRGHGZsBhoVk2F3Zl1a5
VKtHhpOxbkr+lA8LAZ73bNk4tE1tcsCbATZF5s838uqA0Vpy1nY9qsHM1dSGhSHI
tW9x+FL7He4WAukStUWzYo5LphvWqrH3jrrA8TEIBap6ddbfj6R6bOBXE+JpkkHh
OGFqMgkNC6sendqwwwm/EUGhaS3Cz3vuBC+6iqRhRG/t9XHUpg3/zBEPTlP8IRPr
O8T2hZlUhBZdfkmv2KY/pC2+3qTDZP/4GRWwbmPKBLr/19WimRcBALX6kr5giS7h
GcX2ifWcB7Zhb5L5z5l7lqn4frBGH0+OaAMBpvmUgLrguDsF+l+xS29TlnwxWAsW
Oo2TJFEjo15shhM3qmuyoV5GCEn0xbZl80BGNsfm9zT6Pb2N1DFFbbTx/7wN82QG
GfUPBJTUIrdDAT+QC5BqpAn1yp7NTVD24Jvh7OTe+KVbJo1174k+rpo/9h8NNXxy
PwRZqoSNWbbk4emayZEhoAfQP9lcStHP9EY79zzvA9ITzOj5jibFgedn69domAgx
BL7dk85gVvSY/Y6vF3mF/teAo5ptO0yU4Ixyn0MYdn/BsO7OMNwAKJ9NPxgY2rY4
fl161S9gUpxcrLQYmp5MhrPipCYSxDAiAGqcIyGb5Y6PnBLDaXBdgUiMJ1PaoTSl
72IKH15L2L/vp5p8L/yueso0MNGzzRQtOOvJTyPNZuEPDpQ6gUyByPFSryHl1PBb
7a3OZ4UYEmjtUMIiss9L6iulVbBSfa3ASYntcZTLgDenEtyfo+/j400mA3BnLEjK
/cKCEy9bOsHXuzokNzfnP7SCXpdpIC0x1k9gFmNBEcRrWtK9gHBlWtjMchs4F4Nf
yxZb1Ydz0holTmXtqy6v/C7c8eShH1v3kr1Y0SyimbJflvyDu/lCakCdMYC0ddmu
N/SFHA9yFPkv7PT5Q9itYhyo8Dgzt4KJD7hxav6zMg+TfBePvM4DU5LaSv+jV7An
yqqr4JEGPYaLkkZ/J8ZKbpNCag3p52PxDyH91tLo/DdVhZAYLpZzwL/0PO/r8bZ7
2ccmE8Pxkh61ZmQ8u+3CdQihdeGxOyr39oKJHXJRn5nu1LLbtk+w2piBcwfNzIvD
NwrrLcD2Uw5SzCprjolMCNpGTNjRDum9P2Nr2btS/If8Lv+uwfSd+Fq1xVnt3aAz
8bTJCLj7GXGZ7HgYW1/DMbjTA+Dmatmm3uy3HWS8QqDjftiLc/gRfqa6ssw6zxAO
F59+XFHHO+t7IWmpqGQ/ilWJHWa1edM8WXGRQnO3U8NWCqDmyoWyMWmqKoNSVTxd
61MHeQqtEuf2uRmM9LCAq0cutGf4y9it28yTOeKWrbDJoawS0vfKoKtJj5ywzmCV
eKVsLelRe05603YC/j59Jr+4QMa8Q2XzQ93m+Hdu1MPDaNA0xILcb40XqD8bLD3w
sIwEA/Fzdd9tImFNgGBWR0eo9qxN9ebYbRq2N1Fc4pburmqlHCzkShsm1DWlDReI
LkfCI+XVTgMrf2mHk30hlukrren/gWhvLiJ6L2VtZDFYv24sIf6Pq8xMbY3NrSRC
a7UUyCKWgWCuZptL1ykkwXZ+pzMQ5ubvuuPbai6LN7zNxvlVCQKStgtrTIOm8r9Z
APmQ4+gwJJ4ms+RKvLvbVb8yVfFt7F1wNw3esGXUMxWSAfW/REjaFZCd9Mdk9iAV
Q4z+YcGJ9dOWMIA9d4zbgIhTpkVy2mDWWoiVjleTTKRqJF4vZZgjh6uGnxo8q4dW
boHO3duKy7VFPUl5lRH58L+zfO9IpeRhbCYGqNlUQiXywzCLJeG909sXPKnHu3RH
ztdde2Ub0y0c7ZLpq8TmNxsBclbNiPaAKArcWAka+JjE7W8MT+RbAeFv3NLesmuZ
0B+9Hve7YDeHLyd3n2EOkzoeUNmsHY1FhKOnFAA8lbBeoWYuGz5+yBUiAaNx2O9l
VYJrlLGC60bx/rRIYMUytn4OaHvrMxq+5XDaZPVG5XTKWe3hYmbXOXesIGgQ8Z1a
jWUYsvvAz8urD/2tgw75tvArYX5W7AflODMr3rPvoSAoamGVlvgxFW5CS/GGWu+2
c5iiqxDQU+hssey8mq37r19r2qwqbC6yLu2mLSLXg91deU9Zm2b1u0yj3AJODmC8
uS169NnF0XLTjfkIv/svZTLuN/OipXqjAjqdVtUwyb6CXU7f1RGdk/OfNTn+MdVR
qAnU00BboggXXe+63V5JGRQEvNreFdFDkrZ464Eorq47YPAmUx46u9PNrHQUKxnz
io9K9JZB4W35SaprEg6aLPgqVb1YDZkzcjhV0Ntqh2E6hjXLeFS+SLxWeTYK+DYP
6YBGicSy5wj15+NCVky6PXqtPqaKTtWQ9LPeNZ8jRmU1jX26O1vT6frjM27UvzdM
+DEQ4H1V/PihANjNLoI0+Bl+QAwnVJVTkkyvFrCF7QAt6994QG9IDC0BKoWTkw7b
flvwn135mTYJftsN/w5ROb/7HN4HuiFu/eSVYgHQ2BTkbwwiwvV7d6DFthPwQRKh
URAzj0dcAkmzRFL2lJEdfC8MBXLcVsOXfZhe4hTxNuaQfT70vABGmzkgZLEWVbpj
cJI9FRiBZmU/1c8bbpFjmfWbGJbWzsGrYGwDN6+295u8czOAApphg9apcbMA2TMv
abUhB7Fr+UUCpPgof8TufhDawbd1uAjoSqERPihlk7aIUzv4ujT3sYbrOmLXxXJv
FECyb2tWYOhZdu6JI0aNge7UEP8GMJvTJT74JGzej1+1aAStm9BmJjZBJdueUmGD
uI71WkMORSL1uMyuRB2yknSzFAGnhNZdyf4u40l4+rL7UNo/15XxlnJVoBztz1pt
QMAbh+pGMmkGtQCw0p21qa4/qDLfGsYzfGCeh1AYMQAk0KloRc6ZLPgX9LfDUYgU
hwiKzJDF8F9DK3xVfKI2TQpFFIVkLJ5xXXP3xJHkpa7DleVd6aJWV5YkVDfcvxCL
57XaRfDLYP3Sw0GTdWdSh5rcaaLPnxbV/FJuKYKqHlArsYEhOUWuit3uz7eNwmM9
jcuaDZvlOgwbGmux7ZnIQdf1FN3Myj9UKH2iCzHizgyZHU+tx0F4MWlSytmCdJGg
gbfaFILKNxSCwh6//sznngvhwwT5tpe2nw0KTzrBHBDisAABUpFJwE0wPpHo0HzG
TDWAc7LcTmABjcVaSN0+DiYMC+6pcrhVCcO+vgJDnHP1Cep2Le04EzmtybAnaIR2
FJEtGtABYChheS0aWEyEuk/9E671Au3WbYOg/8n2G1nz6zq+HcD0Y+P01P0E/Qk9
IlYUBhio5Lmesjmg5bpT2po6oumaLBHWiOEjt2GwuAvJhk5DWcKZ2P/RVYXH+v9z
LzYD65QcViCausiwM0sxydtuz/Yr63sJZR1ovVN0s89f+JBeu5NY/Pn8AmkMc8qo
AR+JQ28gj/gLlpOe+CtjxmwtSSOe3n0EX4GxDemj0rkLbJ2iiESQwJdJ/3sWTe/S
Nm35YM90Swz7CaOonCce1mqSQQN4O5Bv3lnWLe4NTafsPggX9uj9N1xfT7G3fgwh
yF9G5uRGgreoXUA1ssuo/svhnYJPot/DEcnVXQuiPRRUrXooMKI8Jb/MOD7//KiJ
fQJzD+Cba1NqwOcJqfd7M6wptm/0gepKMLHLkj8sG80/fTfo/wj5kOWLJ0NgNjh9
oRXe59I9HKl3z/VB1KjWstNx2fmJV3vk3gWiSELKcy18SfuI6KwsiEZ+R/ScgRmX
hsaJQNcdegfcp6P4Zh53NWTZVchEYlF1x2ZEWyQXIJIF9vZNQPND/YuIO6Z6oPLF
QlECiKsPQITxlPK6tTiuFw2X9xHrV9A/bc7x6koxGHdb5w4l11NUysfJzf/UyUCD
S2WK+6Qm+xiLfLHpT5e5L2VYbziKtZungsB1iW+dbg03efhw4MtPBISh5IeJc7fj
nm3qtoqKyfAcecHDCxkXsiBVawKZHR7fAxUv/X42hYGVVRYzBzwbMxjrC+HVU9/z
o8NdatP8twqmUjR740y451oOoNcpliiZlKM18c2rNIc0O19IlF/XMeTh9unDV//m
FPyKqzLcMNhxnV9l85kd6V4Uu40WfDuuJV43pL1/Y9YKtWKLwGfoshieKb/wr3oy
WI/ddgYzkJ6qD237d3oOWictVAiss5sfj+2c4/Fg2GsiUpuNVQ2aK5ypBfsuie0J
Tfu6NOzwrIW3iGKUOs/ZpQtistXbNoMwKF4gKhJiTWzKcGXRqA3vP4UQiO3cZHCQ
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Ctho9jq/9drUGVO/5/RaghudkX9fLAuoAOiy1oQTXQG2l2R/WQ7zY3sStKOG8t6M
VncY/KpgFhHB/O/kl+10suUge0zX38Hex178XW0sps5IkHB6Sn71fF4ItHZqaWFl
ItpZ9C5fZS9IpVc/RBOO4HXEXOYqKvl54BTj7hqr3yk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 15823     )
G498T8lTzi36/0RO8cAcuHxjsTT7EvAzIM0xTCI1/x+KT5BbB/6rwrDQR9VSjZq6
B32BlpJveJoK/vTDEt6amWGaqgPJFPEZLo0lhNGvi+4Oh1d+4ub7hzqulK3IafvQ
u3N4ORjjUr2RDmfz7mUcXelBtNWXXJdaoc9MsgCHQtvyhwf6ydPlAFioaJ7T/XWq
`pragma protect end_protected       
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OUjrjfcslFuS6daOwx4n3RFOTK49uBYxTFyZ4lrt6k8Kg2KHQAM1fPxZ4hY1wg2G
dXAR89qtCaXPGSglRWmq8qORDGDDYATC4qmB08kvu8OFbgbNwoefZwfI/CAyyN3B
n27q4DBQNZmHHG1U5SaU6R/SCQBasnxihnw4/i0etMs=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 16537     )
fafZreWAMpWzul9+7iHcu0wXqrtWZ4tTTfQnf/7XW6POQy8vJ6yHEc+bIIIdRDI5
0g9sjmvZLAyE3gCAXmd1njqQIZKl/BrRKXLoOjlq8no5yScOxKGdCfqijBKEfaWX
80fdsOnFcYZhNihsHJFh8WdKCdxzhVJmS6kRODxGWBfnDbtSQ51kh8a7BGX7qeFd
U4sUXZ+pLjYJZLLqjYzw69jA9vn6jvaQvugluTKMjnKioycw8r3/YSMUrv68bldi
oV+fdxdFW7t5lz30Lo1WRFUafrSo7WDrC1sTF9cgnZkJDYxZR43hTN34GhHYaXqc
qJRv1P79C/MLruQSXI4s7zpi8sM8QUD/nlmw1nbiAcl3w3qmQA502+JL1Ccb3AOF
s+w8n+RaiYkK9jACisff1hTSfC7QSmJZGVb0fcuOVob7RalbOVruJD2lUx2lHwwv
ZFAmKK5QoRR/NKbDo9ya0CRV586bk9gcOtSlGJr9jDA/puJ3Pvg4GsxgWICznZTQ
MxHB3RWXbRjpqbuVGF31KpcJYxfUJrb/iDQolQx3kbT5NP7bk+KgRyd28Nhs+ueK
zL2cwjYC0JN4SUUeL3otZecAaw3r6d5DneqERtCUHJ8Mibto0nLcP4mUVRH77lZl
clK2tE/J9H/9BnqgnbkXri48BMf647ykIESDvh7q3xO/I0zxPVFNEKmQvNg6zu7F
4tu8OqNW4Hd9h2PEQbPb3W//9MCKTztNNt3/eKz/ZZ33lC+sDwkc+cjORtdlXbkk
QZNPmljY9+K5LiG9Hf5YiPg8DtQwK+airjRYvjjJOP1qHPisf2hDEdePDogE2QjW
f2bROPRcxR8x0G9dUZfNuPwU75RvTdqCMpRPCBKJmVM3vNGydZsvq6cS9D7UQZTa
Qo4Z7Obw0NFO4I8eVKzkgHR+bFK7zTUohKMJ1jTyi0PCtCscJCJJ0Upuo/SojlFW
`pragma protect end_protected        

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RpwUaVf97NlRe5BuDhSLDegDS8MWv47FY01LfblYaBfPzsjNSv/uBDyVs58dL8HU
WGDX5x1VM5bNNcSIOwv4dxoSHG7LgG/jab6fzTbHJi0VcD2r4Fx7SqGRkgLJj51C
XQ60z/UKalA1hkdSqh0tw1ds61XJ8Q+jlZSU2dNxEXc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 16789     )
Yb3odByEz3AeGwJw0QF0C2CIEN06n19rG5XCECqHWniRORLwjlUgeMcBMGNz05fh
AMi2v6w5W6ZS6KhFcD+2v6zO3Ljm5suysu+opcYqLWLU0R6VCHxnKtjee1ZH1uvY
Pc6M3fUs+iaRZPDx6iKfZd76LmrEHDcMpVo6XtFoubRY8ZjXQSP74LflY39A9SBK
wHL1Cm/EESfN80daDt822KyYpiyBfcgXfcfBFcWfp6qvefYax93BisV9t5Edc/Ga
sZG5NsQrM11VtdKVKpU2o5oEfAbXo9JzbZfdtoFUo+o0mieQhyTIO+cXKBqVy/Uf
nkytJhUvKxwubct1+egNGg==
`pragma protect end_protected        
        
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OphS20/7w3KYDP6jpH32czXVUblThfOS3ErT6Hn6KF0Nr9hZ8XvpRvVarlgXmEy+
mXB/4Mm3VkYbdZQrOBZTdM6+lLPaTl1UVsSRzwd8YiCVogi+wXp4wxEQ74KmHJeU
UYKjBViqLn3r8sNhPkywEzdbeaBz7bOqFSvg8VQLHXc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 21526     )
C8CXXZZz+oKJjKNrU+RVsLgv0/zfmNTXinmbjBTl4YXnKGUvOOfURX0edJD0BBjf
JusztYsdiNSloAXLWTDMMnE+FEDEdZ+QNXexgQhvaQ6oa4qXd4Vlr310+h377Lwr
+60xMAN3mhJtd/IyouSao1+9xEQEcB7y45apJvxBUhEPSzabXuopwd6AMYaD104Q
XYY3YG8p+oP7lU4xRcSMrBYGoVcb1H+CX57QZlyVQTwax/diepLx9ReRY/38yrW4
/lqGoB6JdO4Q8W0wi24L2dR04wfk1mDn6Dg9+gpga4Kukf2keczN8sEEvZQuJY22
/NzDIYaWggQCt8s5p4Ex0YVcnBlSTXInZoJODEP0dIJD9RJPq0psR8RVb1yXzroe
z8bxSjNuYoYH8KlWGRLaoZVoK+01aSENNIBVZd8sDaH2SWYRDQY3Z5DRpMXCbGwa
DEvNLCU9pS3+XtQGmcZbQHcDsd7i6s+V1552JflXriQ3rop1Z1Ire4t3sTdypFrb
sh8R0dCvzpy/eO/Q6m5UfzWHhIIFEdNc+AaWjsQ68A3JQPao1YNQ760y5QbslYJE
Pz+z83vWXegqykA59TQoo2DGHRKRGPQYNNlX2P9+GDsCeYOuwQFAs67F7fPus3hP
D3m/Hl0jIPhZFLEJ4Noo7Ktx2lbens5krM3ITQ60hq3fq+pbFWn1X00Ns+fjyXVI
BRb7lUbtRMx0Ai/QslSEkqtkhD10F1YrkG81dYUYLpmRFfBTTiVqqf8hUHQ1sUsJ
3FYhV0pZnuGuycA/0uBZ2Y4f2pZeCM71b25dWU+oUkw4BJHamN/UapU3BVnhycM8
lNVEYt31YSKmiZvbulh8kL7ma6RRpF7WG7kDLreR1lAeCmeXvHwJXRI8CA2uEucr
RHdrZ2VkVNjWVK1qCZlkjl5cnhhuHex6KZ5S3VZ8sUwjfnKJrIhSpD4L0lMEdGmA
OH2QmTFYwYUAKaCB3FoSCGtRGgjfapdWviNg7N/A+HGrTmJAG1ji9e48zrnUK0zP
R6c7wGt2mPvGo34pZAxcQJIANGYDty4KyaMizCliMeixeh+3zIdi/thm1/B9wNr8
omYRQY2z03FXUX0Qex511qbpWiC/qnfQPcinJf7eJazaBqmhgQJukRCSRbrY09lY
muuiRML5ZsA5zyUvgmah3WIBPL9Vi9TuVrmfhOrYogxOIwaVjHwGdrBrvepuudjv
wBrk23vOs4SmsN7q6fSmzLRF3RbgDvPbK7I3+eHOeMWrZuRsrgG/JXoSHMveA6vD
C7cQpmNlVrSZ5RygqkBmdu88qBx9R4xSFhMdUMAoX8yXYZLth32IUVcDVZW4/Uhs
kclfT1mWmFJ2qwmMCcggeXKVoJ44o16Ffmybd14Rew2uw3xXoYzmidUz/B/9i38a
NELlA5Jj4ZgWMKrqzIPReh8P6h2yeDRb486yOSmGqnIkdak6RnjbDCK6YpjgElBK
T5E1OjH9q9g18y27RAN/DxZQKj5S5xIV4OrQZ7AAQMvBn84KNWVO29vY/cJVkWfs
prHvF/HFmx4VlxrxhzTroqQl7Q28WtpZejbDucrKcWiXVZkLKbNLOAg5wlSH/PVQ
PKI/yF8oZlqs0m9CPDRIRMwZxSqTvj3HJPt3EH4mTfXb6ZuznyGzo6bzgKp50scR
aIAqhe6rIdqCnV8zoS6jlja9cFHED/VtYJ5C1cx/WtqZPrRR8cKzTgBRdGC9qCkZ
RquX1qPeCZaVVVrS/DpMPZBPIiKPx+2/cZK0AHLL3nLzPiOF9hsfRNmYBMF6Z71W
SJeZOeIk+Kw1/LIlFILtma/rtoXrchCy1QETa5uGe0NP68xuuHZnSGwXskeZUzn0
Am5A/Mm0MqH5GxZ2rEcTZqKL54QfOUmznYncpeEeUF72dvmMkgP3Sum7Th7tRtya
xiguPzc/vo1mcPqCd60Ca6aQGDD9wZ6K+o16oAI5xlFD4s/eivqRzj9f2ypbFsN8
wh46vDE6ByJlJsnW8n+ttjVperZGidhvRkI0tJZvgSAzlrRcTpxqvoe2ny86HVSZ
XEljri6QovbqUfDZ6Y+X96AqS3w7LNZpcZPmLnXnmZUx/1r1kquWBbyjCLAt1py8
y2Dr5X/20c+ftkLA0X+8MrJzHkroCtaNaZALlQFPIpRruPGa1At47rDnZkvOYTDV
Pvne50i8YpjIqnEBc0xancYAazEbWXiSzvv4LuHYsWkiXfCb4D2AegwY2CU/lv9i
wgxaJ0UMNoE3Jax2FKNV2pOeOaDwfJIFjVh6a/g3ccBcMpVdEw9KGDNZs01LrC25
05x8PT1CeDGN8P15mHMTnCW4xv7+AOQEjRIvXdZ8Hs2+WE3svyc/0tIa4eBhLMxL
MBs33jqS6FeiWXRdGy7kh3UzgiMVZjFblR5d5FRis9hUn2xYkNj2cl4jAYftjd+Z
6C112H79cgQJRRBp5RPZtZciYIQGjeFB3dzM9uzEDDNdHdjW9yVMwF8jsE/1S4Ba
5DV7ngKMWhjkApUFg5assAWvwy5/42Rd6QabWjFYU+XK1DKf9rm2bMKVZl5feFQO
okW6qFxz66aNSY8Kg1UTKt/BW9QRZXnl/2OV1zIQ62urVT+i01M3OyDw4p8wr1MK
PFrZM0OAeVAWgh74e57bRskM1DxRxqHy/yZUftscNf4StOVHFamWu6sOPN0d9t7/
brdFT3UQ0e/RU/JW2/OrnHOeOqtaEFuhTLxjA35c2G7oJUbaGmCoTavuhcJefI6g
APnM1PsdAl/UA8F0MEfCVECzXvKMkyqnDH1F/GaiPMNTq+pix8g/MIbRpg582EmJ
q8z8gyze53L059C06H0n+ogJZMMxQwNfQ2xW8uKp9qDv4XICR3saX47z8S5SiPw1
hJPptEwZzbZkR5Q5roqYURHk+TMQW6I8r3MwO5dfh6kNxjs0emzxb58/3dpsjnyt
wFm5z/SsLu+cBLs+wXzqfstLatZGAer946yqYu/pGbjVzDX5bSx0kP2FmL3bjW8I
t82bMlNTfshTopvfX9RgAeEHYaz1jOm2UvaBnbq7+59QeLL5plZtrIbaEnaVsPQj
J3omfp1aXQnF0uBStXM6fMHNzPfurhq/hqSKaq/vzJeppGPKHv5hQ6GGHEjWc2aF
1GWsQwC0dljvYsBMMQO/LKc8vcb6TlFSh9pGitMkhMl1rxeyxb/XFJM05aubsj/3
6sdyZMSrhrxsh2DdYNirQzb1IAvVMZZZyjpi6uDqb9ON/tORiqXelTAoC7VLju2W
13oc1L/mu60k+ZgF7cC0T5+YOCvqlb9P44bebd8MGFKX3qWHzrZfsPYsqJOY533w
wMdbfCoblOkweJnVXeXlb1kP+VLmRbad1AoJVf6yxHqwMgc2ok4rL1aPnLUTwUbg
yNVp4/zo1Dv4SS/rvU/AHboXwld2fl6Sjf4/38iQgvWAWuRPt7GMUqQ3QeI+FZrU
AEdjUV604UEFU3zDbwxNGZQkiquvrIfOqZWJyV9i8k64mpwKtsfhP6JBQXfzxfHJ
CsIaRgGt8q2E88O0ncoTiJrZrEvWOWDm5DxS7yzW8OgR7aJmJLPivT137Z4vJgW0
GlK4IlHRs5tOrwaMmJj2kKP8fsCJ4iCDbs5+Hip/wwKiRm9KmVNzyyYx8m+D6tZz
0I3svlz9ZYCkikLsupT8Xq7/3dDdTrRlVC/ejFA7bEUb81z0Apknuo7LZBI2AyDi
p1js6B2IDDf1c8/Qmmk5bt1dvxiMNXtYoQZPgJy3DGTeW12yRrlkzGM9O8Z2dqIa
GjbnUuWFMEZ0e6A6tLKYetgbcGSop1hJG5ERC2GlWs5cThX0RdO+dLWcwO2xkWLb
Oe2uTP6rX4AJKG6BVzEQiePk+9YHIpFdQtpP35VUaH5sRWq9Fcjb1dnrsJ4WcwTI
Z/rt7yFcFETW5Wb2nBYuZx25vMgSpeNDbf/ysfJOrae25kfCosWRjZMMhD+bKnLb
FMzXnUZ6cXEOzYhiUmTlNSJGQx/vX4JlQ9+ToFrcZ8EkmttW+qFKgtsa6jRoZbrS
WNt4cfiKgsq+TRTINM7bLc5f6fYhiH/in6qLEhA64+CRpizlEn8W901lpsZL0v3n
m6wUDz+yCa2Su3t3JxxsaaKbaTq8sxfpU68h+i3eI6x4S5SW3P3Q0iBGqbT6cm9G
Urd7UrxOTikZ3m4oMl8CqnvG3VZ1gFjihWLj3dGRSVcVoYtvLbi4T973HNFhtNoO
Cr3YiAAL3qj9vG+gBjweVkNFsZMoBjrmiUcTcH460pPc+lJ4fzbc2wrp2Uae7aRt
hmKDyNXUwQRRfaJnE3ypxnBw05cDa0OA+aq25aCKEtYyZBuPLUvaf3H+Z/KWfnDW
E2LY8PgrOnMkq/BYRt4p+C464oWrHAlDsgwGGzryVJiN/ah+BKx7TerFmPAqKbXW
gGIRiajIlYLGoeJpJ+N+bYqvqpfYXe32qGUnOohzpFffeNwfUsctDTCo0WTtDfsE
FhRSDULp5QeoEnkpPlXmM4MawXbSYTziYgDnL6gZRfUY0cqTOGzO7oYu4YvZMKuR
pcN0qMpRlkj6tUv3NlnFGi5Pui0W9q3QkpT8KJRohi3nVrCStOM2XyS2M/JgMwBz
cwSGI/g/N734UXWUy2kRXHIGQk3ZJfmLUIUoWYaFbk7Clp1qUfE9gwQMpHovRkJ2
OCjQGNxIKGoVKSoUunuOyF7bhBC4wclRReCZOdV2uodPhE7frHZ2VQTfJjMSXgWd
FCnTsFOVST9k3HAlXGqhMbI+Hd8LKdlM0/UBIxYByPg2rqwIaHMYV0IZ/uC+38hr
rGj50LWmqovO46d+aibAc/0DgzczVdItOuoyd72zXPcxnox1/HhMHoWTJNppqv1Z
aNfru2iqXoeTPRrVVsFesr2/lQNts1tHzxmhykD65yoqmwTwowwcWWCw4lHgfFQQ
Jlm9scvRhcLIUnFocneNKMG15z51/uGgaCW6UnE1bFh8Sedj5IfuDgIL90d7hCNo
7Iu3KtqVEELKxfa+PT9TM76PftX5UHohdD4vC3iYgWJ1xEudvkqDpu4k3fYGz4JS
5vE4d7V+wMQnXM2oaCGJdbtXokfQKPJxyExmVxXupRagqd2MU5YHiACQ9LJaIUt3
kF6tz+J5NnUalXDF5HfwaObn4jlcWa4ptZt6UcdBvqMfhTk1gGyWuivRCtQYpz6Y
w2A/aHDnLAODOBxIRACpN/mKpJlfR/Yvg7igj1VePf4j16vF3zu4ta1mgPKsULAa
sUOFVFTaqBSno0k3t+GYzT21zx3kCqdjQvxRiniKvr/AUoQpgr32ZPXwcpGL1In7
cqbYXdQNt4aHLNliIiMeOkYtnHDM8vgnZE47qd7Za3HVby4wZ4Na7QkYSO3dE1nx
A2oZCTVOFwq2P5gA4Rc2AidSUhU+X/oSGqIJqFDZ9dHT5LV8SyHNy8dRrNQWZ0u8
zM3XMMyqR8Gnk2m31O6Fvxr28T72GkN3thpXiZJrZlZjf+JWhPn0DqPt6mqT7H/r
QPeJc7tN1Sz1WMKDyvKCdo/H6ZWRKRnzSXYHcGIEJKZhrWrhNjOp2U6WcibfJEZO
YUYqTHYnaBTl77cB3NfvCeMv26y0ZJ+OV1IXWf3E2yCX0KWHHq/CBnvoh/6P/Gy+
WsgNKu4M+ru2wCukyH4egHlQH7WSv8UAUcB7aIaWDolwo2rxplKwUZY73uDRmT+E
0Hv+lFQaufVRlujDuqNOFdrYMRBzfkSkJaa94+TQuV8DytKoDn2jDlTUKR5egGB0
E8F3eZpUlY2/yFZf5RTLnPBBBn7jLe6E5B7HrX2SkMVs+YvWYHuj48yCg2464GQB
UJ4ulh1X1/0Vo/IsbUGYxxdWWvTyugbSeoT+iMQAU5Eg3ymJ9WJv/7Vj9Skcaddn
+KaGCMZrVducqU7sowAQIeqQ76UQujdkdo4bzezj0uz3nFoSkI/wZZ6gN8a5/9/+
ybTD7Btfjz79RXPSuA+ClRwFb1G3Cup3ynyX0x73IR16ngijN1vq98QyQTKmCpd/
hwI0YDP7zKHKUhuimzJXyunlyDDOtAqmhxqsXcwXjM2OXSBB90hlni7m3WfQKFy6
MqDMK/YD8Wni1KWqkhe2bJnOBvwANY0EKRAtgfZrURC3AruO0P1WUa90EDCLcuPd
ISVIZmQeA9ceBzkA1mClAhDa6NhH6Waxv4+Ki1rSkHWtk4egOU1bDiIcn87YcRpF
GcnoxECx2pP94Yd1qiEgvRvaOnIGtegwGJihrsHtpMCmnbVKi4y+tFM0EsT5SzYe
Xk3g/0ApUUtlS7J5WCP6Wiplj8Z/GDG3+o2PtwFVdmMvutyV5gub8LxEpBx6/yq6
`pragma protect end_protected             
`pragma protect begin_protected      
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
i0Ak8NU/DIbED1KL8NkQEgUwLuxYiqQIP7VVjOkkRO7EL4nDOMjnUcYod7yotbw5
WUz/twihE0ENedze8YoeMkwh/3QWrsphvc7k1pGEOnr1bpesXd040Zx75Tg2NvZv
96m+FIBBzzlz3vtnPUeNxskjeoenosbGrU6parRVH5o=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 21760     )
R2V58srwWzyOVpcYA+X2ogEoElhwsngLHLfNrUgw9Fs2IRMXTEKRqWSN81YYyxSE
u4FQHbrGrJSitDrY+OPXgHMrQM1RnwE7ALV+l3Y/2exVxa3fHg6sw7bxemDOdfZ4
+FlCQrjs9ziw9QZYWlEK6NWnuw19rMcN03OQB7wV79Ok+6HOH18KEcz2a8h5yEkr
rVSN9Nnzf+ONw7djRvp9EyWVbRUiFVbWkzd0wcCLn24Q4zgiFHIvr8J4SUO26T71
EyDXQJe6o2OTRPeszhNLTxEUc1vou/CAbut/vQXPlq2/gSzerOeayzu2U4YXQxGN
`pragma protect end_protected      
      
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
lpAbZBgGTGH8kZ+zUNs5YiymXJeXTKCP9L0fgyW1VtFFmHS755gG1/f8wRupn7q0
qEGZdm7c1KJSDgDg84Ifcs3sscODKO+JJDt6hbBb87es703nrc4YMGV55Jq6rgyW
+UA5CiF8qf1+maDJxDUvRiFj6EPfFQ1/Ou5ZAz4x4v4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 43052     )
6JN1XZnXJBQ4E5D7fK8bx8KFaHAbyJCq4f8RHZTpnQwRAuvwGKLUC2KpZqvId/r2
lA0ZFYGrsDI0x8duWayLHiVQODKdamvP2H9BPweuRGHsLT9usMEbeWOD8mFouPp4
j9PMHPb+dvbrWget0VuLvcl6/LfeU7jSSeNODuYEk2HPBUX46PEjKJSuGtjKctkk
0bBcVJtsW6zuu+3ZkNvnjv1quJoNoZPuygXycPSXfD/qGzi4wS/9qY7sKpt1AFGP
tHZKf7DAVveduOFiyhL5oyadplQaF6VNVh9DW55JKhrLqnTMpDHDThyVg7Yg0ewy
FXKz9tc353gigSfVCMWLo5QVsx0g8PwJF85ov1w/phR8Txv+OeuREYF55GTmu3/n
l177/lVx4T526HNR4JYKCQkq/bGoVNtqr14cmwTQMko0z0c5zsYq3w+hO/bFsVkk
jX2u1e0yLb0R2FgRY3vHnnFKJA2nIFbijCu0eLmpN2NmmoP639lG0aLgMm/T0Vu1
9IuplvEHoVnZhjoyv1+BkH3vpb/Q6r+fQ/AeZOfRQaza21SMjNZWYdSsoOoqCFwG
u4dS7zmB5LZI7hjPfWHgysuu14j2I2zHKbzUFuPjHzfVvgPlcVgdYMfwC9qAiY6E
bPwGKBN3IqNqqALwpIFnAaZADBC6tm/SPMJiH2b5YyQqe02nHZeK72rWsBGMdVTR
/WLWjaz3UNeiSqoxX9LjS9pbUm++8pTTceKqUDUxNnZV6/BGNaPoZ2hSdIyTS6e8
OCLqDNBXIeAXErmK1GS/JEz0iJYUoYEHfMLDAztiDNeFjuk10BqiNqUu7nUS+8vv
uqmJLtc/bl+3ZVFJw+DAq1WT89+IZ6MTmOsBqzI76QdVNyhLRb4lPIbb23Hc1CdF
BiAvJrv194boHoKL99t5l3+ypPW2n0CIRhBd/UyHY5OPViGRBP2p5ll9keI1d6U8
aXIyUhemJ0DE5UISHcLGeRLHhIksvzDTLIbiAMsqWbP/3gj41ZP0XgEqryfJB01/
/lNaNPoPbqJiu/Ha8yBolY8NJsXPia8cweNcv89YUUUzgQPx+moBwWg1k6L5bLDU
MFQ1A2LlT1eb9+djL0WS15BGKbX0f1GxvLphfcj5CO7aMg4GyXRQP5etymBSvTyR
uIemJtv6lL+BHo4dNhIi/jYAdEyYi0p5fX/VvvjNPe2I9jWBbcIPVsJuMMuqVrJW
nTVni4VpR0iuEKPfji3UEDoYP6Che0rzaW1x2t4jBKZmYJY2SdmRAlInXxPqEAHF
AulWHQQvl5eOo6WabRm6M6Yka154oPduw9WpBgI+6/m0WAnyBjgztm+UgW885ZPb
62Cj4Q0+sh/JoeJLqszJhLi7h9MV61iwaeB/G9a/vTbqU95hMJ7UmjjNsulCTctr
w9IHhn9+ONa88UdDVHXgYZxFS4PaJmOXNZnJTFP+htIK5PxZn3EWYb6ritc5YZ5V
o38UZlm3vJKvtINC+KiKEN3nHT331T/RuNFXZl1EFGnJRpQZN3/wGT3mKcrtefYJ
M4hKsRYDCuIOR2XGdH/oUravaNbf52ZkDNBFTdA3uWEI7J1PP46mqC56zROjVjlf
VfSHDsGfskxoqlDEh16+EO4X8anvjxRsPzsQZXPYFBT56Ko73vASLuMMCcOQxH+a
57i/UM8/nVaQ8xOkXQXtJf1qP0nhkQXBXoIInOMSFNlnVC0vlxvvICJH+yGfbT4i
4ApeUDRFaj+koy31sDPj1UOkaB/R8kNkXmEmlb/p1kIVObF+AqsSj14MU8hEnUkj
0vUaXoX0WuS1LUtS0jjCtsC56aaAi8YWeWHbAZNtb8KqADmzL3jHNC9Vk718E2xK
fO5xkI+BumXDP6/gEKhaB37WHfG1vmOrm6xoSad0GYGf9zVbySj+w8xc+JzPkkk7
L00VGslAR1VlcQYUKbXvffXjt3Yz0AmTRJ7s5T4eCpBbOpWwxV16TZeOjLYQI9qC
HhqulAdqJfkp+sxNmShGnMzkIKgxfQNeFg68uZ6Lve3IRPFD7iuULc1T9AJhT9HV
VzQx1I9eGQqxLvrxIRzJz/MCevaklvJT9udUquHzV/jVCSKHurNg6vRRTbvtAqoY
jM/vwFKNmFYdkFsPXn0V0rkNdiRIDKupzD0FSfn7if5K2Dr5cDaO9u1c+lqEOjyK
YJtQpX6PlfqAH7/gLnFYrNtCowMNwb15EtKJd6yqa9SQlv1H+W2V3fRPXiHDYwie
BXepkEpumGwTY1Yy47RQJS9KnbeT1PJgQ8tRmNF92KeebraPTJ3qVQI3fwi3DXiS
/960hCNGLZJfEVBjX851oEglVm5xC5nld/Cm0/BiPp4Kmnc1r0x/V1w5bwFtWxsj
tIQkv27lwIWZeVN/IhDJ1QxoblzR3Qicu+7l2Weo2GyhvkQ+a5zPsedzIz4jpVRO
46ebMInZANZxOw+wH9madhrMJkW7Qk1ezppd9Imw3kLrXfwvoEZIsZiDANNWSKoQ
/i/yKIavv40/W3TfzjP+LqNMudNMXM0ghVeNHJiIOx5doB2EzfojFrKcd8ZUi0xS
wQiDjFfhujhMGqvolHN9fiiRcYNf9URXv69+zKy0fi0e3eS5yPE6q1iuN5aU5yJ/
xpayFq42nEm26ehqEsLk7+Aw+KRVdMZ9QKMQhgDvfkNCuZYvcUiaVw8NNXhi/J8A
4eDUv4ji9LBiZ0pCzeIMYRq0B1Wbzx2gkT53N+CVoZadGFcaq9Kj/aM6vLlaMWBi
q1483p++vBtjo/7cBzyuI0IEXntCEnhv8JbRhw6F+7aO9RnSyJDQz1ulWVS4WuMV
kH5ViP3bmBNBhp287MXp6pp6Xzbr/qrgHr4PzXp4JHpLQm84fDvb3Ei692qwDd3k
03b3NT80DGXmQbSfSfjwiHGbXGRk/EbG/G10DmCrbrDvrD9LxKVTOJr+UFxyGWJ5
he/k0l2JT/Z7g7EgRw+zQ3ojFyLKlgdq/pGFqkUDeDPy7iOchY2w+OM52A6oJ4fB
UZiU/6Odqd+XfNjlKRLCyhP4eCptGVxxZFTrryj72cZCk9188ACvjgJuLzpeR2t6
/bhvpcrGpMtq2bMbWCC2o0rOigJC2YcowBGiCoQiDY71/wuC0/FnwDk7P3R6sA5b
FWYXKhi6St6pQtPfLWBsp/oZxagYemeGDF+puvvqRdJbkmBYzcRrCgA9BvLbkg+R
Y84LUsUl7G/Nea5qUYA8Wm6n6qkNJmgO96aNSjD6nOgcTlpuqbwiQBVCgwcgvij0
HlsYTEpju1gV9nzQz8MNxYLrZWrmlIOGofYpJpN+6TcomgNboZeR/OjeFb9FbHXC
vJHoojJwv/kcFnrAOulTG7w+7kjVwW5zXzjniz1V0N2x/nvNZYLEsAOQcURp83Lb
/6/7aWkjoEqWpCGCgwuqlAnu9mTdalKhUYP/2dgSALxN1TopyMmZmQxFqmcw20ks
t1aQ2Yu21FjlPUJdztOJqFNsRqieTG7CAMS929T0/UsCRTFVpKrSciA8GFLzaSH5
OrtaE2qv4nlLiA8paZzsgP+xuz7rlLsmhJ+cb3CCP8mloYkgAmX/2ZPhOLSQAuYX
tc707hFh8/dy9R4y8XCjVjO+Udj32y+nAf06b0tKoJdIy6blIMf4AMt5A+/mOiEK
wLsX8B9Dx44zuLeTAHGVyhIwxSUlzODFM1OKh7wKIiD4XXyejtMnE/ti44V8ZIOC
hybAzbM8GVaQ7WMKG4ZKgIBJ/JVH+Td+XiDlBdnSH8JuhZZ+KXvFQ8G92YtwxxZJ
KNXdcRJXRjftbasUnLO1OOVgHE6J9/Ehhs9ZWdUxtMnhJ46aDCvFJwfulUq+NRiR
Yfdh+bidtSRqKz8lh3vZGbFQiaoh0wEIC0mEmfuw8BjoeF9j8aiwn6wvEMue7B73
jGh3PBnxHdJBNlFK+tDjtJJX551SrxH+BLjydlHYjs1Fgat6i4YOWjgeFKtXU8Cf
VsyxrG/IBNi4PWb/zlwCzIZHhh6F5mXDh677WO7hqLWsdptQNXuM8NbwPP9D+YHV
LeJMBW0NEuGKMK5W8DB8Tfiwsu8xC/Ko726Lk6fp6C5edS9NVwtE2Lkgl4X4Z+0W
knpHRJ6Dwh0T4w+HjB6kqZTd4LI5PN2ANzeecHmhVx4rmYjdArQ0waYpXNDkvWTp
2AFKAdfoR7MpgYpHEjIA/qWXcRaumknRxQJ19c6wrTJovHusY/+gk825jMF+L5cE
kzZISzJvsyflIXZonuCehLRpfgYSA6sBUbD5UKqmx1fJYV6b78Z24T4GLU77Tpz4
XQotkelrrVsSmPtxqSiCQJ0nv93gumFq9cg7PtyIbvY2+dijVkp1coQhl5BaEhmT
hG5Ra3maC8r/ULEINoiPTz4j7C7BaFxwOoUABNWMgwUyqfj8GxvFDgTOj4ahiDee
EbI58VWXZfs9FIg9btEARKhS+rgw3CdyYiDFL0ZHPPIKRKT3+jPOU+p8g6E7hGGc
EtgBsClyw7YLglmAqKfoDKYTp9ew37rFL4PhCuC9iVGRQIzs0RZYR3n2ny8ORrRG
AbH8SDvsJM7GusPbLQYPCErimM28nC6GIv6KPAFvX7GMIqoF6PVCMLxqHaKr2fut
xE0KJ/4skFLZIr02sHNgstE8Q6jUhVBpsaClM523Tx1Wd/Ehm0ko610QIsulohpc
o+4v1/m3BXZnReCggSrEhkT4ClDbMNil3SoSX1hcmTqjU5mGg4SQAFsns+ltWIcI
4TMp+byDAICpGXf2jO64R1lrbPkogCeXp6k/KqtThI8TTSQjd4kFOF5yIyjByomh
06eSP0wlIjE1yXzdldymSw+THdOvsEhXUCVa5/5yU8yYo/FZonWPJSunV4cBvWF/
qUj27/j51md6lbHBWoBBBDDrgRKDelf8FnRDydRjfQg7j/SbFexLxWB2fhbSqIo4
7BMkU90jDJzHXPZFqKAAHECBn+4g0DNlA93SotWAGMuePgPEJLjH2rwFpnwopFQA
dgm7wglTzb04+3dagOJQ2ceKgq8LzIn36A45F2EmNt/p3J13adz9YKiezT6z4n41
HvbcOU+biHOm/I2cRElccj71O+U05xIIGpWPPZCsaobRYr+RDTkJy4da6Ew6a3v2
c1ttz5DbxpyJZmVmgWc/CLWo+XxXFk7rC83vZGrxTsy3F66qI0CfptYDd9Slj61N
JMQavhpw6aXMrhdeEVI8MfdmRpsaxfpZSriV4rWA6hxSJytDYGX7xv/xwL2GNJ80
UoyScECJ0vc6Rc6kV61Q8cjsedIScktLW5G76hyfOFCT1Tr95LxkvoSbGEYR6D1i
N4rIMrb7LQvFOZQ5MyDDi4ryfOrst+vQuXG1BVm84oj/tMH6zY7hdZaV/vs0HL2Y
xHavSGmS212MaPsKrqmCkEqBgvNYZB3JeYCflaH5ZPplCThPyilQHJaY/2OJck8m
1t71VjDkuFgWYEzKR0MW3n8Af/CAkfpACqGf50k/totx5M5OL4efoV2cZz56Wr+v
7Up5uFTVX5vMZdwGHiDFpLe1oWQhNE6QM9KNipCDk0iVnYeMl4aWOhiVxWjfxI1s
u3vt9okKzSuiuwdNSCWhEQkQj2YfBXnCG1dKxDXT8QwCJGu7DBfrMJq+/DD1b054
5N7KnUw7ZgaTH+vWxJ28Hy9PC5pOaJFDCW6NcHsrkMJC1RT/RVFb8SU5Fm/l8AhI
wi/8F/L/6MKBxZfswigwdCpiZybT02HmltrJL7Frv0pnXheXtWmemQMU/zZHqRsP
s8xKtvHemO5dRMjka1KFcaK8bs3QbFmAKm5lj4UOwJ6SkY3e+bE4IXmuGKsKcAIj
D07/Kk9j6y9ihbsb4yqUaL2BLQ89SlclsOqkcW6zlwEoUEZv++gvMH7/jHqtCrOD
vOZb8PuVvcBoOS72bro5yq94l2QlL1Z+zj9u4gUXvk/cSQFBadmszzcVxez2bBqM
7bj5Yg9XaqCN8HsfxjgjLRbOJCkINYWW0Z//+iyuZZViIW5n7Lrj9rNbLRPUXtBs
bJz8B06fIVa4n5ODdH1fu90q9YCETwBDZoQwXGhtJN1mEWfnAJ9bKRt4SZuAIFJ/
tGOZ0pvc3WpzSsVf5frLwtBJGFReD/MM/4TrLId+XJlnU3TIOWti2wARmHAPQWHd
mBP4TzJXJZAXNapn3F5DZo0r699PhLOYM5TCyx8QMwVCupVaxCMakJ8qX7xKmek6
HJaX//WmAVFORr2jbH/ckQNX+ri0vw44solRq0Yjpj6c0UEm0AGuwzrqMcQnlt0+
Brsi92+rnFjymK9b69eXmCG6SJ/mULYhGsHASkj01SQ7phZ0lCQJYOoO3Sp+LDrW
2XOCOPVRZOVgx6vTG3d+RpELhHraMABpVqisSkA8gh/ElWXriF6p8X7WiKZxq46R
bXDI/MEm8aNhxdQSdWqIsN9ei6i2V4dou4z0dXXEfckA3TJvB+abUCC7edL7RFx2
ImQZIH4aRBmw2uKnz+MF60r8/AzDwMiJkFqRwd5kkXyz2UM/ZPSnJ1MSbMbN2u9V
ggK028C88dQmE2N+L570c2Q3/jLz2Jrk//yc+CeqEGVkPIgoR3ev6oJVZB6NEDkt
QJLxfiuTrcarusfemSglDPRnHF7/LUiuHqYgJ+nLfNfcDQwLyWNVLCRz4oA+Hcij
lDO+NTl67k7Mt+6wHBFkNL6mu7ycPyxMgsgnzLcF/c6u1lcp+tgtCBHMKSfmHYsQ
OxAd4Fey0Y59f3p1X1dY5pgzOSKgsljj+Oq9bdxmS9gfPEGuVMc7gROEx34h2aqN
F1nz7ENu5txfnDBYKIayalZQcOcCFo1Z5SFfA1Mso8poHPlOUbqVeIWdF2yENK/t
ctBBBra5U4Lkp+Mp0T5NSrlNEgMVhZROiNtXFJ1mCiQwtTHK9D7NKOEZMYnNUtQF
dbfPZ4f+v2Fm7CDPVPvemTCXkcrOGpJQoNx6RfUzgs2PZRXFSfPxfMXUcrov5nDf
Em7TTi1Gm1SDiv4midMvOwj68FKRklulpHgp4w0Bt9d3V3PQp14rz6e9Qy/NE3lI
udfLh1D8u8A06w/puTKlJNJkwleDpMAOWeblKfX+yxyOaLt+etaanYddCEGbvfKA
y5Ic8hidgFZl5i66MEluPzV/sTqPUvZ0El8yLn8q3trDg1Z+Bp3Da76TQfSbmYjv
qqNN4cCakjp2+O8/KlmbYj3iqdrj6+cyopv4aUKlGdz23qA7Cn8zgrOkA3gQYut8
lJenUYpsXxO/Z4vbanzc3n6Zge+EjQdPeanvQGUiK33KtH7tCIOld66Df4iN+6xF
mzJpP+oJPZRbsTY7zbkQrjr+171fDybn6yRFfibdE1p1rLLKmvYC1tpXwPhrDbDN
eWvzOkQ46UkHAPH0quPfj7Zo1VroFZWQTZw55XocrglZnldhiqMRSQvYdcd1iDCT
ZJj7EwI4jqK1iag737aLROneHsdk2EEWTlDsLkHLB6/9QlIm2hyyj6BRHWYMd8+H
kVqXkk5Yr8suO1QqZZ9xRr6GyoEbBh04m/hDs91EgUToIuYhaOwV1Qv7JBYVb+Gw
boBhng1DZWtIWDl9are1y9uaUWvwDeDGWP4DdpajateozLzaKKmruhZx+oRj7coS
9Wqy8sOPnLba4zrZFPK6/ntVSzPbcF3LZsSeUfDlpNpayF0p+IgKElVYOKCIgah4
ntlmmEyq/t8sK3C9V1IqRtk+NikLB5yg430ncKOe/K5KN2cE6NMRwb5SCN3xuDnd
nNPUzxUrkck6X97vJeE9WgBfggKulend8CIreBTCRbu27ark7zP7pAfAE2rR0vyq
5DXM4vN086mKlBzUUGPa1gIxLuqz/YvURfIR6SHJjgSai99gLW3rR5l+PahvYT+N
4G3oAjlw839rSjMxrQrzHWeggBCKVaDAS6Qosxss6l1fN9u5Bi2b/0r00qozeEY1
W5xiXWWz874gUwd1Q5tFtO46yGytrkayjFAvU5judq79mEZOaJCOEEigNP9+6GPN
lxG6M6v9IyxS/WJL8dEJF828d5rD5Jfo44a+KrjtzitDeS53JSvg9BcBuriDhhw7
kgtsNANvXmsSoOyZKDxWy4P/4QhEhKxCKz45TDjV9I3LX3I4aoVqRCHiKOdTPY9G
lwwk915tKlPlrbBgLYV9RUh61SHq8T6D1GdszT2T1ygMa/jzlZIn4ljJhgIAb3Tb
qTAVF5JKtW5HWG8W/N0taymvcN3hoOXiHDwsI4qmQjyxkOp2nU2o1s8gzB0abLl8
dmR5kKdxK0sbC9lTofyyFwET3wuuJSvhA9Q94A3IMVKMUi1t8dVEOQuERPoDgLu6
bUOVa0RcLZ6W31PZMfCGhK+PlRQG1jf89QZScUgc8RTQtFXu7DSpIdmoS9wN6I1U
BIn+nXUk5zZjCtGJ9Ya52DGgtKtDvCWqXnVy5ZUCBGxtMv3i04c1CtCq2t69wMFM
cwiPKUoKSEYx9WgM1cuc4tz9XVJwEAqx4N4a2Wuz3YFdm9rq3QlsTfD261aGA+Zk
f3YvCB8BWkk8QSZsr/kz4z/gA/Ub7F9df5NLbXI07xky89MNf6IJMwXbnsPpJIRr
36MQ56XCAk+wHjRvTLxeX5K6z1AZ4pLz/eBvwW56luYAyQmfOmXKBmc3L1ON76LN
WZmdS/QvmGQHh1NMbpslujvWZljxqSmtOxy2cLV7ZEz/B2Ajon3FtykQSgBGl6g6
6y1fcexYdWeG4c/8qV7tfE7bNT8H7eRWZV4SnPRBbnRCaZRT6Qo9S4G2TnjdtrIy
9je+DO2cSK/FDbC4x6YZEwblHL9awSRdJVyROOHzR3GmleKP06NB1yEqksL9WKhL
Pk/m1qyE8f9NOXK/LBvBkbgvorlkz0TRujA3cnHGN4WnoDn7H7U22l9eryrG397D
9PLgXkdMJHtTwTJN+fDTnXI88OEdJ+5dTha+eYz/iuAeRSKzy9/2Bf7Xqc/Oo3DZ
j5r1btKaOw5cy8lWxqL2a79vnIIqQqV40ekc4ZT5whQOZTYyaNQkai2Z3Tp6+Wg5
2Wcr6K5qFGH96jGnXtV8XK1jybrboovOLqGOdsnhBCRZ06+mtqwNTvS9Z5dpjrbB
zGFiZFvNxDrMoBPy/uDLEm5lIn+3zFxB1Kp5k0jjtbxnMLO18InMPgEDaDj2yck8
p6NF3HZEy08hInWuf1kXkBU/26sNIsFYUueb17pHrC86YmT+jqI9io2rT8MyMLCX
89/pFqoH9eiX37Vv8I6dWDKiLZCggNVP9DokFO6nWffux6uc2+BfwNpoV0DQ39GS
SgD4BUp1mzb//tC9hfNKbxY8EEGqla8lv5bH9lF+Sg+W42krSWNO3/7+oy0StEnf
Ec3e6sgvTP7nH6S76h4WfQObKfCCT5XN7IXsgxYZe4zaRma5h+a9P3m/y3NbHRtw
/W9LU1liMJZ1xIZXc1oQrIKXtspg0UiSn2Zyptiz0D2fNlqPWo0gaYR757Vqkz/0
HlzwR02DCEGmmx3aYrb66coZ80tO/bZgtHpUsTbnL7sYICTx1JVrXjvN4FFiWew3
+YmLQFKClj6N1KXktx4Q2Hkje2FC9pr/tRrgYJSgXdnF7glX2j5JnjFZgdgBzUUd
JEBnwxUdyvhEAPIX5Fr/qY0mbfA5XiudmWs6hA433uteQrPoNjINWz775Qstr3Bd
is/P+uTV5i7Vo7sqKXwhcmLlMq0JPIdqTuL85jVwvkb2XSq3RkaV8wG2AxXMmOQD
wnT+yRlGS2zVWJ2rNl4CuLrCy4PKQywHlDXZYpG0YlHkLVtyptbdRO9/czAC5Z4H
py3abkTJY74JfKRd2J8Tq2NqUAaI71Z6t2zK+G9JWxYJJdizV0aFLsMqwBWDsffy
SZPLCuCULWHf3IyKe4H9ZPIVO29DBukJhiRjo8w+L2I7DKTzR1mJQonwzpEBKLcG
tkslsLjJOlFQNT9S/fe9+x3+IMXSoIfyszsYgwe54DHDC0pI8mN7n6ZJbhu2GyWe
vs+HHA8WE817AShmynbPbA1dpry1IU+yezmG2NWIfr9TxwjNHtqYAmYKzzNs625t
cb021uhJiG4FyGdbYPhY0luCm70/SIF+J9dRsBCCBSs3b8QXQkxJrRX1XG8XQJiT
t2NYI1e3ERXNeYZoWGEkt1okgFpIjWRTD9aGAIdLnYLt4/MPEHgZVl1Gc/5g8IfG
yKLVaMWW/p5ya9YMq6yaDgtZpEp3UEdGL8igNPp0PeJpOWEYP7tE0VveB1j6VwBq
/i86bI2APiH+vIHzZJna8BDXfJnsn8hK3x/FyDELPResVaFmwSZH7JcIXG6RgOpy
S6UltFbz5DnV3mUc7uC6U9O8QJWefvn72wQylB+SxpNdJT3GiebQ2vY2IY3DhUdj
bNN5q8q3F+hJpn8M9ALY9UjVwMQDOpArtX0ZjY0mMom7TKw5oKihnB0wg/+gRmYZ
PaBX7TEbq0+2L4qxSw/M3RzV02wPysprBE5AIiso43kX+ZvrrZ63Nz/mBGl2abbK
y6bWPxbHMLTTgk2aKZsgBvBDjMZ4nUbSuzM/yw8IZjQeUF1fFPcvZ88vxaBBZSO3
KaZmzRSJWLk/sBm62tVmOKGA95WswGR6WMO1/KjlhVHPVGMGH8Auuc2iatnUf66B
Rcuf0v86r759xXjnw/L8sniyO0Vy5StqpAOtXBGFp3VKUFts1mAHuQ1vQAHf+Chx
Z3vuwSLEBJMdESGTIk+8j5Nmnzct8eT/Q6J9lBVNgDCSMHAlBzyJcY6JW9shhu9s
/MUHrSn+tN3Qm111XlofS6+JWrREuj4NXUbAXrtE3k+FBWPc2z2Ag14NrWymCisI
H8wcgt+34htQNrTJp895JmS2TBY2YoAtoobzw7ZkcDo1yafjjyiCgV0D4aU1XJ7R
VgRJ6zyMgad+oP54OFvtHfitCi7waCr1YUsPnxEv/dW0vqYTB9viKL4nEIs+LviE
QltEyfURpLxyMT4IYz1w8YGaTXfKJi90d5p+mi4CXqbzA19GIwwxNI7KUl/RRgan
ghy7HFNpdr7pFXnhfGGBjgFltRsFIH+C4Q9BI9taOp49p9RRMbUokYresSOJmmg9
qiTg5/tq6Xft7JnK31n+qzYbq5bwtzDen13OHUnR5z02yhFIN5U2QPlvkvIABWrg
BrDx3LtJyqgi9F0aCMg0CYntYfaYZV44i0wov9YF9uoKA1BDgAqUdLor648RemIp
ATw85/W+64ihdbwUH3bH2NeJNDH21qAdBMTKY0HWrK+0tCYiCO26IcWy7/ay/1oP
kdbA74mRW97BQrenf1YxU9cH+YY2sztkmNa5H9x50Iv5mhWO/KiOAXHnOCeyi5dA
rgvWK3dtBFOBPPobS2KgREJKyU/bj5i44sJpp32X0b0B5YTt9Ln7ga/GC16ZaLhv
GsAHKGlrRFASDTDm7/rqc+Bajm9B0YY4LEOcse4nEOOqdMHqkCpLrrP5eMwZOGdI
KwgfCavxuksQ8FONkMY6qL8+de3vYkdnuSKSb9X9LAioXCfjb1lnUQYhRaB7i6YR
C7OtxYxF3JaHwUVGzxl+mLlHMmRzAU4wmj/jzteGQpW8ZXGRizBHkF991d39H5dU
b1Hxy0gzBN9iDRfvObrFHFQUTh1uaD/oUb/4nryDEp5pcWlNFM0/tWIfN/KzRLVs
Xi9PgvkFzvHYGq5nzWCscW6si3q3rerO7Sz6L5/7HcttAupz3j4MpDYh8AzpG8Qe
8g5WJDf/McXmub323aOskedPku7X7OefM3N9xcIRRp6yAjRlBdQEtpmOCAB0pmEs
On0ytSHoQEtTNWKwEqrK8u7Yf39bBhPfIi9Wpjrg91o9HoQB0zFP8qUk4oFuhbYG
is/ytiv2KC0pUIHWI5pFIFA0Q2baWb9gKR19JDxidkigti5nHKb0MHiPQ7+2Xjok
4RKw1w276GCOfMTtD/MWU1lQ36MtbF3vw2FSYuNZWICvDSg0TK9EnU4x0DGsOuW4
Oejjr7QBX9ExYFYHLKzzhIEfLN+6+p9u7PXKbMWtbQ0cAu5LfEW0OaD6CT0CVrZ0
78fR2G621B2bPD5cI/HtIsFnrJtV41v8VxN0Zit0sgO5tm86DtjnnETjaIC57Xfx
KJ0QzYqCBrA5vurEVFHg5iTGGAnJd8QeZYhVFJCHReOfkvcudGSTV/LkTL9RfjIZ
ft3NZnFws20iTwrcPHDoyulEwzHrhKtzqNcvosPd/9l0bCB5HqpkpkLAFuaOBssd
0CtgjSPNBOCWbSPJC9hmpI+Qr4sgREH2m0fWZ6M8azhiVQr9d0PyFvXRIclNMWko
OHaq6b3DVMER558v9LpUAhgGylii/GrWu/pOs+l1S3UWh8eFIhWLXXs2eBQ0Gv+c
DzSZebgWceWYUDXAyJZTEM1/kSF6VXz/b4kN4O9EKAS1mJ4ZpmGPBTeirahaEJuV
27+V8yBt+yE1LzlyZiGDaT74qodfEIE3I9rRlUy2nCrXb66pqiVO0zFscvvz9eud
6bxmEV1RDxr+gHJQitljsQL98PT2xTXZrEs45nG0ChDjXIwbJLZKYOtG4lQ8ic3n
e1oC0FZsV7lLh4jLpu3qJz/mYxLqZ9rpubHgUYt6FbGedad73G/g/wFIYoMiACMH
Mlaq6qLXppKq6DEG6gL0mwrqNWEEXpW/vNzlo/Kxo+gtPrsCooajIPMLtME/2M42
xe37SxkCCmB8pV8gqZPvHNnM/wCpr2IoEVzWV6ywe6kFMpBKHjlUmaqp+QrExD7x
nj1sFvqHejHGpKD20luNG/B9Ly3uOj0RCQO/n618agUghRl8WiN3OA58xuVsqVU5
9GgFjRDGg0ctDueQyyLPBbBu+sdTHJW7tw3Z8poaNUJ6kDP9cXwXH8Oi9QqTgEoM
ZMj8sQFLvAoEuJ8GdReaa614f+Vb8i4v4qBKj5ui0dUfIfXCRdiNxcqeT/XVRDgV
U1e0xwt9qtDzCtZye1C6oD96s3RhQqA7c0qc4544ImcY/YUl3KOhS7bu2ComfzYA
Aik0BRBxbzuDf5/45yXm+pT2Bz9IMQBnns2m/eC6NtvFiDD0/wNouENlj6GV6yb2
6+30lWASjXaXcWycfxDR5krtdAQJMAGMZCHXLsgFU27Q4vqSFFSQN/6SnP/Zha7h
6oBk2wj/kqNJgl9G8A3go2Go5ozIGzlVWR48qaxbTMg5iSfy//FOLcfMPTwmp/B2
Dc0ePTS9Kf+sPLylXNchRA01p5DinA858UxMtr5Gn/lqL9vijrMH2JvASsU27gc3
dAZCiWuq7H5qAkxRvuVu0DFrE+hTVLKRvbZSsGo74Wg7citJjmjgeJV6U9xB6pgl
VWrtQ7bwxk56pxlPTWosAg+8RvEBRsKbpa7LpxnZWrawZu/tg2ajNaFGAYR/obne
sCJA0Y8hxakRy9VEZ6yrCPv9/E5Zjtjteqk2xhjtI+hXEspzAGFHQZof70AZvBit
yu0Luhgi0jexF91UZLaaoDVs4miI9WgKjRlZHAAMSSr24xGKCJ8pVejQQntd7V6T
Sw5VzyfQ4EJaWVRgx4kOyu8bAscO0x35QFxUgkobtZIK3LfT9CY/tC+Fw9plcBIb
fl7F5KhSDNx1zJHa0TQvuP8QWsPrgj9XVWqiFBW+Cugy+W0pviRucDCjJtXMfs3X
eo7EY4KeKr7Rc7lydAm5NbCIO0S6eoSaoeHl7gAGG+HjsCL/t3/qkyHpZi6UvIat
F4XM9ToY7ULhLOMEjLa3YLKKw+9ACTxOiD6XaKIU/ocnGrlqepAVjEi7LJ2vaEcy
3elqphT126eTXbieeMrg5NxJlDKmCLHpg7bEPKfh8V1E+kRWacPeWSrd4ykQ2zym
6y96oBCUH6ZnjWGcHrd3WnRwl/MPLOFvny+cYRKtMMyp5l0RO8VTNkljyVhoFDOV
1AKd6lu7A8I44poMYbs4pkDf496qmlvKSq2gB4ZrIrRc8d7ijhEuuEBO8MyqjbA9
YtTKXSeH9/V6kKXkFbySnx4aclQyFK0QI4MN50oUTHSzxkUqZIZxAZFkOEPGYIaD
+nLP0JCb0GyVv8f+MHGL/gKNidX5lJw9ZXDd5und6D887bLaTcwbRMrwWzQgzqpd
Fudm3dpZyvZVisZ6wiF7c3RWFWlFRMCKUDeLllhGO7BXM3dOtf/pnOJ2R7YwoW+M
S+VCHgoiwk4A26+ahR8bJMECMlwz0mlKhqV8/dg6yBaBfphflPw4f8QRVcEoqMLV
wnEqXbjLtz/wNo9pa13q2TR5W6Gam/SShttZ7hMS9krytqEMEalMuQMHmr0NZYI/
GTFXQ0zLdxdWmovQaYGq3GirG8lDkKvm8o67szu9mS+c8/9+YNq3iq/a/mIP0Dy/
mkap8ChY3Du1UnhtSKv8nyvPSVLzdD6r23ybx0dlQEGygCsqonfjzn2dVJd7yhza
7lH1rofSU4mU3WWNx3Rp6j9re8dI3YYcu+5okW5T2NaQDWzzOycLu6KxkGH/wlgR
iIYplIa3gIOK8hxrWJ1jzub1BTXHeTPcbjmOkAfrDZbqezq0Lo0wcDQRow+pYVg8
rNSOLxpYVTZQVb0E+Vkf+KUoOTEwaJeSBFQhdV4taS2gPSQramcWLw2GJIfbDXMB
vTdx+672GKl7+Fu5lypCYnrrFwLqWUriD8LwFPZcYFUmAj9GzJ227BZYRQaSwJs+
VLe0o6BzSAbyo69Xbc+YFEBKRZBta8+jQQPoytSrR1TaCQkLu7tA3TtXJXp7DqHN
pI2ov5UbHH3HXWNkY1Zkcdf3EOVPG7X2Rogo7vPBHOYeMCQGhsl2kGSKQN2mM49C
FscPGDF3dsK77v3akzCQJXqyyoVU/qTQsFtUty3oj1cHeUzrnS/WHKGrUIqJPotu
ZBKPJ0tqEekxzvP4CHY7dc5hZQWI3n0As5n+AjkPDqPTBYhdC9CEXSqFUU54zktF
mItqFpQ8XnLMWzitLt/O61kLtrXuazyS3nWAiziJcIinKWC5lQxsjOiHrQpS3FLe
OSKUCBJUwxnuPgi4s1PjRuQRP+BqTpmnVSUXlhhzVvLXmz4hbLTpbPlsOXP/rIkU
qDfB/eR59THPusU/HTFPYdgo/cOvZ1LlaD2Cr9PDFHyI/3hJcYAy15jtWHQKRZCJ
OvKrAMcCub9xOu8Kcijm6VDw0/tnQF+exLws6DmKVjsNgoc35HoaP67R9D+4/Dp+
1+x/tGsre+IXrnQQVa6qDJ+6xoRAcMlJdGtWyRcYynVW0LC04LYwylqFmYEJ1bn+
n6akrMj4hNJ/DDqfKWtRzw70qv631zFK7YXkRFY7saMm3eqPfBjCRn3jyXpLqRgj
QYGLqQBmI7RhheZBOVQ6yZ/QyF9Jnh0GHhGku5EILVdS0Siq/oXmFbtsNER/txlf
vomiLZDWNL24meEdoCv1GPFnA+m1AJx0K7YXJTMqBEv2M+53NrRd9oTp3gIlI5WW
buyxMlSRCA4aOBZ5az7F3z05i9vLHGD1ja+tRV9+a1A1YswgigLhdeUebxJa962Z
TDDSKvmoImb9CLebherVl+65lYgHVQuX64midEnrXjiv0qSgpsslcrzOs13qjJG5
Jvf43C9ReGYV+chg1vKpKww8KD9p6olL+j/Ct5vH9fa6gtabQ7aoDKA4PGA4F0vc
mJWVHDFdTYp64IUxSaj/4/aR5n2J0xN/7m2PHnAjXuV6FhvEE1inmd75959iqlpw
ZHHIbw8RHKSMkSfTkq+koBxYLTbcBu7shM0ctw0cPGCSHsmRFko/2dpOjD2yc97H
iMioZG7WyYM1HRINFBzbCLe1oTw1TLWgM7dX78ojJylnOobT822LvLuDj/F/HKl+
4Xw+cvKsTp1Mw5EVJyn7mfUQIvqDINyccxjqckOSIFt0hIqICdiD6n/4MzxhBpZY
XGNmyDq9dl/gON930VphDftJVx62VxPSt7JpIhk3ljC/pxForLPsuzHeFge5V3/o
zLirZDyywOs0Njuwz5iVVQE30KbAWQhP5GoO/lS6cuj77F0YP6F7Krgllx8HgLfJ
wEsdz3rlnq9DXq2xgblRfQf0QhMaoB3gUMR2GtWXOYdjriPKUNhlcNcBWvQma1Kj
TFOJxeTHyfIHw7dnI3Z2A0NSial0XilDeuecWumu//Sl+KVQ5NLMpfggiIDWwCGo
eJ5XhwkvZKGr/iF1zXgXvdSbhWvY1+uvOD9y/T8Qn/Zx5bZgW/3X6jfTTuqBgsRr
uNdKmLnMUZCclSmf3igKuWs7by+58PCRAb04Ni5/4dTwG9VyTQIfK47OurHBQggU
ZRPg+qs0Aj+WCuy9NBOOd47VCxlXtecMJNygaMcJ3v98aHmbTvRiJTVy+Dqc8OPe
MgRDRzhCPiN9Qc7X+mquqJvIMxO/nJnBSdMCN2MLy+S9E+ZL4C6Yi2IQqYHUDQFF
3CQWEfm7aAGcXdInhdbx30p7G0/0+tPlg0JQkucfOjNkcA6v0n1b5hqHqnGsXs3f
35F1EAd4ooDP6LsNibCBNzFNdsFSVrWS4AAWeAQRV1IrvAXOJ+k5y64cXdGg/DD8
YH6kTT9AjE5onVVgacVIVSuKZvAlI4KQVNNWnWucrPs+us8dRSiIIpplqIKm0QvZ
nnxx8Jgm5OTWuTO2FZ9lgQia5NvA9VqA/bfjLWqMVC25LvMuKUqgQFp6qEVaQB9/
NES/A6MYWN0oT1fa0HflFd8Kdnap3BRAqkwFnbG9LlyqXIPuW07UsGUC0FmZhvCZ
/rEFt/CMLZ7tNGjFjivPmypkwB6txRcIAysvxVmauI21D+xGSPDxVS0/qJF1a9/p
0N7RoeHx6uVQEvk+OGqcW+qDPlX1EmnXtAOtk0soE9xhYdi7Fy7OlW2b2fT7WEos
k1EaoJSpGZU8cO7hyfx3j6yPxHsOifL0gOO0DPqKvYf03Jx84QIHmxRkHiSShSAk
1DC7IFgPcYAwwtcu7LFJBAwMjPEelCC5EleHQB6KA1Lm8DmgMjZMtyRogQbkwf2t
9zPmsodYHmSqcDVo3vFoND33jeEA6Dl/aKSFW4SS9gb/tWhzHQYVrAKfEBtOdZu+
OjHVW/5H33ZxzgRsdH67k+RY8A2D6OTeSU3j7/VFCRbznkU7cqrKxts0NmNTTf72
2w+S8fO6XqRsm7pha7ozRv0Tw2ynLx/AOWDZcDZKIpF5rAHHarDrcYUZzrJkrT5r
y/SExxt5iBX+pJ/yWD5UigwUf5wn8d96fGAkgfa53hh1YZE5drIbsryDbA8wdn21
I1Wjs0m2JJSGGHc2XZDjYLZy5qTcbk5AeHajN2/OAkqGENlv8kdtlV8KvRH2dza8
5TthyKKO+qV/Bhv9Pos6+tBLjudQfiQj8EEg4i6x4qBxk4YnoPtUxu0wQj+DMPDd
M59Ib9QWu6CBnEP8Ftg3O0Jpsbd4QmtmNTS0xUEcPf+aDvEAxdGj+Me66R4OSnRZ
I0L1Kl7zWSK/1ACd1KBKSJLeZ6HupAVH0le7JTJ35M86v21/t+ZEaPGXNC3f4hxa
Uh0Q27ZUgPLWFNsk29p9v5JwAzd5V17usV/DDKYWGAl7zZ5TXMQ6KLo+urvQsyi7
dgftIBmVTF/K3Ssdb6JztpUJCCsnuaLOAVFVRQhNFwQmgYUgiggf1ewVJXCFj082
W/zPLD2x2YtuTPlWS22PBPkeLJCDZSC5UcCetMUlJIazHF4Ti2YUoOv2Qp/hlWai
tXgPlJJBLWj1g7BCBtC5SO3ASu5kO0QlWr1pH/A0YMEIOuaGV/GTWq/fyfcofwXp
JE+OZbwZ826KjenomlQEMEia3wPrb9+Hxr5HlmNOxJc15obhG9PrdjjR9RNKLbwJ
4tg5sZJGBfWSoQBPkZ/3sjfDCcpHUOnAQj0TNZhXBbdEP8z237xrA+yvCl/9dS9/
PsGOhmARkXed6wT05AZ2MB1iPjsUcwE+9a119Klg/IGqDXRQHpcb/aMZekvFZ/sA
yXx9oyRTx7Ou1UsWMXyE0T2SuBZnSWjvHjxgC5RUPx1n7M/N+Qgn/hXQnuAjgorg
UTI8SKQznb5nn2QypLOmradrvcB+Za0NzNBXyZpV8ZHga15uL9r+qJSRb0iSrAzV
tQLcd+08AwqmJ9iaRgx84gqEOUhTJ1Zw/vERJU7DJvRLjZgEY50JKyg4ZoqGCAWx
khWj8XTUsTgvNKjuEJl4E5R8N11FKUOcOULpNoSWcRR2gmi+1d4+1xGHLraILmS5
T1ABjNh3vKsF5Sf9KoT2XyJdLRTsOlkVjmKHHih7tpYX+eteaIbfgoZzkrUn9pO6
9hfJD30hb+3wiUPMUarAfdCPBffJtLn+YFtmNvkbKS369sGbjb8gUvRmeV2dfA9H
fpLpyRuPEb+bBulSz5GD2bv7yyvDnvOHOBImZSbav15Q32ucMz2GQxjzSAm/m4M3
+uGs77NrD7znX5KN/4vz0cY78HMbRaXSgxNSMYwrtms6n/m2C/aGMnFQPzA4Cgvn
PGuHPz7JYVwZ1p5+7akAkuUq1Fk1HCTKls+BYU/wsdA1U1LqrzdOG47wmaurXnsS
GtiysZAi2Ukg3ridCMJi8+hXIbCESI1FJltDN5U8n//oRwT64S4iv2xABgfv6aHg
5B8c3n8Or42UiuU8kZIEoYCxpCRHOTc4DqmC5iZk2mPHbMDv0aJ15geyYFiNbl2l
fp31/aQvUlni7d/d0DHe+6/+a+IQZuhGRHRqtYYijhpx25G2wn36FOCBcvKmixwS
8y1IKiQHE+4Ix6GPj9+6vWzdxuuQXLy/XL6azTQDn8/S5QYQuwF+fWcStYmg/Ali
BuMsUbwGqJNaJgdOUhedRqYC/cBVXkmfnGzm79PGRROwgSt1yhsd0qccKjLyQloG
RfWcU0c/QRzqsnFqPANavQmsULkwFsTfh+i4xQgAp7YA85X37YoeG1OgZxdvNsxg
uJ+t11EjZ8fmoKLwMoBvKQXmhVYinma16doS818pvuJig8cazlLIqEan2ljvy4eg
pzKjZ8Xi64bYUcxBC9lhlKorQ93EixS7b1uhsGpPKzTxLMiirv735QLh6CpmGYsm
6+iWPAgagx36S2Ng8VDIJFq31RyPmbwHTnK7/clT0m37AAVFIvylZurLI+PlNLeL
DBgReRlvjLbm7dL9VpoOuGJnVrH5GU5JVZ8tYvazmJygtL+qgKclDydedjG+GPua
t3x4CinrWlorn+4xdojaftL5g0J5paW2O2IW8f3zwWlAj7gx5Yigc0GdYgQrw8oE
JyP75KzWtEZmuhHGTxsjHrnx2WtGzcl6ezqUGvWzpwcL+0dDLnrbBuQhn0+iPYnS
It6sxaWLmt1HsdxQcYJI8irSqduAxgE+RuCnQKrTWwiTZKQrk3ldattKaRaozng+
vSCRj9XNLXoPD9Sn/k3oTcOnVPoJ4LaOh0wCXGWXYGOIdx6LiwZsyGkiaPKfySlV
u4lg1+uSJxtq+M8y7ZlQeIW4fu28FVQt/W8/8KKfQ4w12fnmkrzO5ry9SVAA+rnI
av8TyLZECapWNqngrVvYFlfHmOvxTP9K28k1NFZSth7kgovd9atO5lgLek4K0Ey4
9EYpmV2LoOa3aANguhCbHbUsroVxKKI/yb+cq9c93Nprd7H2bqnCvFZ7sNg4q8Ke
zvBpHnwlXIUk338F8sXpN02YNHOexOWNP+tSVJQ2A3RIktCSLtG8evc5i2RhfLld
1G6Zh4nQqTYmwaExvaB6Rv4MMMkIrjDOlYqC4TwxtQNFG9/X5FXKf/dk3ysE3l1u
w8guq5rrtDi23+DX1oKYu7kUg4TXgtR4Ld8S0kv+P86nE8WhY50R4txJYoXFOwlU
gg14ImD/YE4waRRynZqKzWHkCXsEUauufAIWmB5bTmollrBv7o4KtvHF6IaisC4a
d1DNQYA88UZysjcTw4/DAk3aCsjRRmFey6/1mcWxPeuIEKhxPQPrFFNgZC/U0W26
xy1imdrV0WrYyUXNeKj/qvxHUYAOkBcaNEk0nZv9XIGSsY88xuhSlY4UFWdvcX0B
BAWTyrRvHwZ7vLPkDzmbcaOi8IMVqzsR3M8EQO7VAel+eRHZ40hGe5Fx5G1F9ahn
eXElXUrWHx53qcSEKuVG67+77ZnX6U+LTT4U3E8NXby2PdGH/ALf9xVkae5OE40e
scd7fj+/ZCI86moOymicmwd7tQHkxNDFm1KZ+gLfnvHQppRlbu7QDEKtGYbXIGwS
PXpHwbzx1G/iGsjJZPZDuSgE+nP+foBP1F1lJV8WdY/wo4kksHSFEgZ3HQ83UBhT
6pCCuLEFr54BNyuYDQqWy0mmRukiqN2ZVHgeS/n4ZyjtsU1DNJQOpUz0jAky4TuR
I7Xb+hw9jRnAEvssK+xDVope+9pccDqYCjJMj6NZ3qSWu3ogMY5cQI7xLUx67fdc
Z1KpZHXlQ8pxzssy6dTop8My4neejVuXpN5LcxJ1vT9TJrv31DNFd8UsvPmGgeh3
TmWPesobzQHEj7bs6GbQN98+aMF54h7Lb4QY2yxBSl/aR5Nvbn7CI50rpzLQA4ly
LUnIjMvcEB/RsPaDRQrJeeNeZh4RpqnjmP1n9oukCsGxJG04RihgBrHXhbwg5+kv
8zDg5bL98xeNwfAiuOpxxTPJmGKRx1OrJZMjY/mSy5VsbA8dXILKYZSNdO93X6Qq
sBQLU/QNNpwUPynx34V5uDXJdrn4wldCwFU31nTiDAbGPnq3yU3TR2D7nejxFBmD
2vNjUC3DmrU8Z2vemePX6+FgVlFzas6aYYLlrI7/kWOKhuCG0LW9MQm57Of0YKiD
Oy9Tit2+iJWiMzQj4ANcovd1twb6L7BhcdNcSwn0XdVQpcWAUOU71Q/ILnHPmjHL
oK+gE7ZQ8Gl+84QTT2y6flc3Vb+x1yRYByiYoyWc0mfK8p/nfp+sGFzzwYI1JfDt
2RFj5ThSkigi2ZtCpjHyPKiIBLciiN7DdUk7zixpL/w3H55ZQQt6Tx2B6yfbGCPF
Yr/W7Tjj6EtEXHh6Lc+eaKa/juVmM0EzyLkwJxyLyoZs59EmA1A83qxrUqMtiwfj
sulrg9tzeMPlAJGhrvQjsHUTfDex1KPeyDd4mhIGFQibm4lYNzFzv1TpHTcECggr
MlvY6p7Nka1o/pmGuFAX8TCFj6k2bXciK9wEg+zRM3YAVp0ZGxm0draPLppR4nIc
vsx9oOQgHOp3vtpArVOhdg+kB4xkyBjgEBg3AQi50oqC+i/ZTbFLoMWE1nrZAh1e
u0+ODp0baZvlomTAQwtMiV9gjr1DKWeSFewW/HzgdHkovjblD7fO6ZmFrU7sf1P4
Irk5wEYV0+R85F4Rvku8Adh+7PnDPSJoCwuQydrT7I29iygKvkfskFrn2ugaUsQA
frlJhLuYf+Qk1wt1itcpI9UpfGBV6FRRVI8yjykksK7BfhKTC8CHPnNZQGJG0Sdb
I9kaToqm+yworjh8BKVKSfdwZ+2qmYCIt9Q9fA+KjgUis3o7JkVoe1fI00S0/OAF
UqX2xjlfxIJgyo9f97QaHVq/CA5ALURLWZoqaEyoGu14PpU2cacpWJ2NwXvl3GUO
DLeAVW91bXRInmSoLedMOdC3QyuAL4+8TsOhVOuS4VQE3PPThNXystNnn6sCEn5k
kCjfzmDuHd3quS+FtdaPmpuu1VwG9N1iJ4Tk/AjXa06USB4ndkHi/mV/rHCZ1JdW
W5nmkdLDWoOeXXtOqnH8wiXbt2uzuURJuxI1qbTxH89Rvch/zAImVelywPgq3ke7
gcaLSqYbATyogD1hJF40YAWKKtrQBoC1ugR3d+MiJNhVJBWkMDMl10dZjbsQs3z/
7HNU1S079MtmFIUhae4qaLD2rGaBRDyO26u+JlSuh6uvJ4atlDFiVRxweZfDJE+y
FekXVw7eAdlpM0l+1AFBl4o3SAM1fKeglpQR717ISOQSnRjZ4hlidtCyoGCAoqKS
4zbP1JKEs2DfIfsS+bc1cLtCiz2LLdwiikHn4TPOrVVuFBPqm6numC4KhELkIhhn
ehqejJpglOjkhTs/KjM8v5lhe0iCeDhDjNkSSo+Jat68zJy+CjBkmTYKVY9AlwiD
lkavzPNziSPvn84TwKI03bE/frok+XbhV+wIwrYEol9csUbmhKI51/BrztPs7aY5
j+RKOwuc4MKdRzzg/j0DW8eNomJ2Vw9KCNs1VohGXsI73WvrOrvrlA+BKwvR9VK5
LfrEzJhD6+d9dmQPeLCUZntUEhtpTMrsiHA8gihwwLjHOMObTITxktbydmn+V4uQ
pphv2qJeZcCzohVnbkuF3O6wZ51BpjPpIeWvT+43dfhp3Y2/uI8lZo7ARS77Ush6
1xDbqfaXHeI84nUl2aHIqMZhVfzwh4RukNVCvHH7ETrHNeLpztSgUN49bYYXF0mq
KlXV9P6ZZUCxGOPPtxBnl9jtcJ/Qm3xS+sJFlo01yPqSxSdPo7PETqAyUMn2U9sd
ZTlJx49osmdfO2KO22DxMcQKqYykyrMxj3NQQ5I/Ai9OLg8a07B0lsq1UtKp4Rrs
sg7Omeka1rKFFmERld3O+ySoCBOdSa/DaaV6UCViDNnloODr94Tszw4yN0KX80Im
TUygjud4ZKEObB4zjDW+/xA1jwq7i+5WWe/0uqTziC8HkaIPHPvHsBnjQvr56rNy
TXvXEfnSbpNKzGWms4JfvzRsDionvK/ZphZwA6sdGG5Epc7ljy4O42573R78duQb
VbYbdxp0nmKCTN4u2CNPhj81NPW8cspNW+pvqK9mAfCGyJy6w47cALFDRHK4Qv4h
KnRMBHCX1JiJKORDWqZsWsRiG52YZgQfXZ5T12SZ7MUu49FynfUdAcqBvUPWE7aN
59+Dv8TOunLmc9BPA0bytDlPsFEU+JnU+84IUjEYx9Nr2WOhrJNMaKaR/qAYZOIK
4ezy8gFz/dizRqxL6fMDgj3+ACJeR+YUcHKRNyTWOlW8ysV380LjqVITKj8EJk+E
zpGg2P4Mr8a8hBJcbfHXh1OTTNU9clseuF+rdRKMm9oUymO61kIEOybd3RbIQCW0
arJTPGQhqKYFfGgkcHwcbQPx6bZbmibKAOcwX3xDEuiVoEXN0zNgoYJB7bq9ma5z
Ikxcws4trbAcLc/jp7le5I3hd0iHVqiQ1V/h2RmwKQAReZ/D/UeJ7Fk+85488GQo
5MctbVhrIdxWZPfAblsHZlmK3od8nf4bnMVJUxcesb4HvWyo27Xtt/2PRl0uqNGQ
ZFTgJQPZxec86oCaUqikUUcNky8OBiuAlccz7FWITd/0n60lP98hT1ZZdWC+yOOf
N1oyNfsLx6N5IlaJkrymUNPFNt+k7XDMapbVHE5K1aJBkiivjQdajCnzRuX626GY
CK/gBQp1OWsbMiow1J0foAU2HxJntEEe3INOY77rP+PnIP/VsTj1JJ9QoWqe4UiX
bPxE8GSndzg+ilgPwJLn2dSzaaWewJJxD3aOxavdGte/FVya4H679dFxJ83/cqUL
/X+XnuLr/LM8eqpiS2dYmZ3vaxYLyb1iSFgXQDXioqNs8UCrO0MXEr44+N9r9eUg
769oxsFHT7dhRDi1vwRsnI7pZFkpCbSJeEJs2zlvRiRGbfhgN9SBtqSrE6nbijcd
Jp+81/ZP11qn2PdivQc/QAiTx/gYaxfIj7FbhQ+5jq8yYA3n5fCfxaPWlN/ewAZi
w3IyEZll+XMx+Bu9CzgOJL2kMp3xvI9+SrfmQZ1BP8NWjqt0mvm5eLaQ5sRmaMEN
Jx2x28bNUciBoAGscNdGugI2rbY7yb/6XdV9V6/5/wP8u0L8TOwMsEs5TnQYt60u
S0iyVoUtoClUwbjT08oNpHV41fxHvhIlALQvN1BBA/xIzuUKpyr1EYZ6we7eVnuT
OLwDdIJu5BckeSwWr7R7NaPOnhf3LGvkTncyQoX7GpKpTJ2UGUCEfNH/x7p+lzaz
fev/0oHMwCdpR9czEOVjXZxIW3J9HkJt+7DAf28MG5/ye2GBCxzMh7twxF97NhpF
IsSbo4EMrh4kmWMdMkvpHA6oSVjkdpq56tvwlu9Ff9J0ArbVQpQnZCtJs/CzH+h0
NfWgYA3DowiSLiFEMRx7m8Hd1qTP48JWrpDsV3uPBwf/gmKMcBa6QTpUdNo5P4pQ
XR/UM9wCcGXaaM+HYA5d1JFH4MZZx1SCmkw6nQeamwnzEFfVVwhErwoVblQLfpBT
+M1vTbyBwQ3Nelt95hu/ik70xcOar+or0GJi06rwJoQreOwMFj6DiiebhEY1g9Bi
Kwc8EMhFncehZKnXSWYjNLK7UPIanIrVYZavAR19ZVi+EFE+PedeG8LpAyculDD9
3j4zgZkRPxsS5o7aCj8CyhL0OTHEAxlPGRDBT8ED0nujBSkiAKWhbxKqEFiTUQVx
lWpgsbtqsNYSq8uSpMY58X20rV8ALGcXIFhxOdgcsdyI2jlOqln1MoGPY+yZwrR1
PLWR/ubz/QSGv8Ba2CHg3/Os8MVwGWMWUkNzRyl6m1cgnkc9ThEt2skYt7AreA7q
WGLdVj2wVllz35LbnlE/LlLP4Krw5f19aP6XwYnlAhQI8DV6Weo6XCLE4TebUAvT
vplWuRLWs+OnPBv/THvclDuwXW5Kfc3m+905uzEr7G6WZXZF9aFYLoBSGrXVd3ly
ENsvVYqCn0lWF/aCOPkFC/KudMp0sDcFsYt3UQSGfxiE6CNpNN3muUjelTL4/XKg
Rf7AFsRoDs0sxXonFBV1mQ4EP3p2WxP5lEGkpMeBYmpEyEup32k/nEiwjgQJp1BC
kXLwo2TyiK8K3/ZQnQN3hexQkEZ4APM2RFNGF4qXsNbTxMTId0RmJdL1HeAjuDYx
cOIsawK5WNaIgF3TIfls+FKfZoXMVXWZyOfgJkg+r34jxTf61YWWndI8+NlJGVxv
m92t1KSiu50vF5Xvqd6bfSlQ55O41fDC8aGOUEdHyEDHu8TAdgRvi9gyxCSvIEYo
mEOnVyOL4PrdX4LFfJ2ds8REUS4btzmioX51wqUzYJEWzqfYtb2QJCC0yfu66Aih
oky0z4tKmqi1SrFzNrwePoj08HVch6X9kyxtQBFo8SyADefoqVGG7lqnksCvQxQp
8QhgfkEQ8vEpJRxg9BLs4isUlDozJr9YiReIeRFhRgYgjhoVGwWY3rfwSGOrhm1I
GBHnLttO+Gd7+0gkWfjd5TCeWx2kk/Lid7+nMzZX1hpvb/sXmV7cXeqJvHLcyX/W
ErOcSE0AdI4OkZN8xgFFf+yi5EZ80IxaxAng1U+9/WIpr7voM5G4pTf6jCSq1nbs
GSylFjGGxNTLZrJdwQkKoWMqnOK8fAE9yDWy9RiWDVfXNpdrs8BQ1OurLUIn8aNJ
cfOZop1o+Fz++JQrJcN4fwlelIQJiR21oJYyKksxZ3+Q3xII3BnQVYlouNjx+RMR
1oFh6puxxUbXXe1rVgE/YxS+4y+cfbU503hXH0SDoAonVdfiSRgVimTm6Z51sA+Z
vxb/dpS2alhiEkGmUOz5t7Rg3PzPiq+6KcWg3mfErtvx7OvSNqu7nHQA4CzxOY6R
b2CvkqrCmMYmtAEHPLW58fuig/MH5Ljzxk8p7A8UrrQeMGzLWPOZqZsx/omcA3El
zKTYPb6CI0RDZ361ocbCSflNNBtpWaht2Wof9J02sypvrJZSOJuJom6S85gCLnj+
psl4KtzyL3axpOZSbmq1Stdo5feLGNlq6N2UbS9t3H7sdDrAVuSYbNQmElHbOi1Q
loxWlN03/uATiDZh879QaLvRWcYH8TyJxOVK3pc9aVfD7Ue+A1GB6R19sgtj6vBJ
zs/g2whTQqrvmKo821mr6YHtbeIclUPuL+wbfqzgM3JjPlZ685HCmanKwgGOJ7VV
LQ1zYqavRQz9VvXxdQt/6yGgvbFwc/x44LQKU3Xvo5Qt6DuMU5GSke1bbkqLhqkf
BHSNMIhGsYqDZQIV2ziQzhF7erLHK4JhYXjRs2TPk9p8pdEOJfZRzO0XpZY+GkEB
Wc1CiX16DZkILIVM+8PYiqDvoSSCci90o7b19yMzCmc//Ul30DEjV5t8m9BvRLM9
0xp67JgKUROQLNRj9e5qwdBeXJSlyBOFbcY72HzAHTEBLQW2AneKqM/NnLnrW+tP
0SqkeDsarblrddeqLnyeIYq+yZ7VZscRUtbHL+KBAotvWtomwjVYv+dhLTPygruk
K40CHPKWURGr8a89dYUnx5v1/iirpmmxK97lKKFq5J7Bif+d80gH0cciktr/xNTH
stS5ebxL5pb1osC0I8hYkSSrJIQEW2gM4Q4fPfkLOPYoUichSXa9uvj1/AlXwxMF
wtN3Od+SKR29o4WocXNKRM5l8C9zjAGbWecjrxBATbqMx7d5XF03IXArNqQzMFQQ
jM7Xq6lEKY6gckgfyJomXznH77HJrrq4IwC5PiaMD2sdj++IlES4dZGg0R+/tb/l
DH0xMcC2qF+vBks+YtQWsgHlNiapjgynPlftUX1ehvtdjtyfIQ0wURy43X6Qgo6y
Ehm6znHmEvWFMFFJ3f4dIgTKy7HrOYVtJ48V6xqvDRD/1GIu2wQXIWLXzwBtKVgs
etHQv/yvq3TeqOV/84xzwwXDvGKP9U4k/DMIKhPcehO0vqtfpxDUBAE5+65bSldv
1iIKzVnLncCvRSDPadWb126JoBvGaPCtvVjXuKSCBb+fgahRqv8cxZsgADvy0cBH
zW+2D3mCMwWkuyHmcp1gWOsu7G/CitFNNOjLCUfrMakYEjs+RyjFvc4rVBGZhztQ
q+bwnAL75QqXdlldRqlUUelR7eSWOWTuRo8H83kTMS9vy8FEAJX+1i/2o9sKQbbT
bLjsFnbl5OGtA95GPw+zwACFOr+5uFDXxg7qpyQ0tcXPe3blHJN5O7qtGaCEiErK
jEXl6Y/afWnVlye/cJ1qoEkdBB58bAoF9s1kObfa66j32whQHntovzdOPFyLtReh
D2Ap6sE4u0EqxU5NTr82dU7lVD1I3rChQVOWXNi84NqT9aCFg6bC3B7oWkEG/UOY
i0hLVDdi3u6KgDhl3aZBlYtj9UyuANYP9QyARej0KihdigJ2tXtolQd8GiaV83xP
KMpUucTpkVedsmMS1y6gl//V1k2+EdU7O6/AVsgKOCkZQm2+uf/WyNQChrz2PUY4
ax4fgxXHgxeTLSCx98zdbe1Y6CoYu634SD6nhXGfjil95T8vE4jWSEvGABnmGFpL
p3kSVOSIBP8ow5nyGbXR7iSvHeXcwZX8wYSNQZgMCLV6OFg332WMZihzIu/E0Lsz
ifiIakxa5Q4mdXib7NnoPWndJCNVfcMZe04GR5C1/3wbv6+QZyP+gaZyklldNJR3
0wXQaRWuDNVgwNdgzLu6tX70+uLOKLb8tZcJ4oF5Seh2XUQ/F+l7UQyxB985a0Mb
v3pk4XBOgI4ZTUkAVmN72M3Ti1jF8I2ENqEiqh8JrxP5dsrb101z3jqjvO4OMx+A
/FpWz5ZDwi1lf+/eU1UnmcB6YWbimLyD4yJrWm6Q31lX4KrLfOGtLDPvF55VR8Mn
F8cWrEyG67Pslsw4fJuZqj26x3fQesP3xPPNHphypNuDE1mPvclATRbY1yz/GjMG
PGR6O2i8SJvhgOHHGtC/+ccB/fhLx8IDX32BTJOby5Rte0T7q70ztfmxve6M/71o
l//j/sLzRdTTNGmOuBadmzdbZjZyTx6G8K9sGbS5CdWCkgYTkW8ER2yN/e/PIjDK
v4o8rDMgTX/aXdEP1xa2YsAbunHwdbme4IxBo9x3wJFHKQ8//b2X+DNy9mga9KkS
9p1yCI8U7+GQ0HRJjjZmKmqaerj/MOyaMPxso/SBMxOkVJiF4rBs6n1ZlEeSm1f/
tGqwQch8NqA/O95aTii2bvSegVMHqxAfdh5CvMhxBmJORGJOvzY0ZP/XcwErRQN7
rqE6eVn/zAlnarIhtt0Q55lpuJHV4+NO8+LW2Ilhe/5fIC4f9sgHDg0z48W83ZM0
YqP1oe16q0QsBVb9F5stw3IyXHMTXNLbZfmUsA8MJajB9487CLwJtj2A5Abjk/Ii
ePpNmmJfPuBz+KXhhRzaoULzqkYJm43B69MnBxqMu213Gavq7fUUgFwxcp/AE373
f8w1foN+wmp0ZhpMnUtJNq+yQVwQMLZ60AnzuTM7HudT6kAwUnVFnf8Sile2e3gP
IcHxkpwsPlG5Qg7DXrecFkgeamDPTDVcqi3ml/uDzw3dtz+xaeaHgx+o/6CKM2Ci
BYqI8+qp/wz78iirFs1vfyhkHSMm2IeyQoMg0Xi7FvWisAQYw1tVJUWYpuTnxyxJ
+hOgYLlxOKMiLK8gKVbZsXTx9XFsgTiwXOodZUbPqYgA3o+B9nI3/56x15EVXoBz
MwhucwsMyClHejUMO0D/l828CB4vhVj/2e4TmEvA+B+YKsVjwNsBHfIeTKqg4J5W
wMYEP4Xhx725gOgy95+upeEl/+X50CZZ3PlUxfurXkk=
`pragma protect end_protected
//----------------------------------------------------------------------------
`pragma protect begin_protected        
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
GEtd0W7zJrhWsU4bM5328PfaBvcDHfpsC5whE+CfEAngaOMQvq1oQgqn22UqTfzh
slB+9ji00T9VHCTVsPMkEQOTSUb7MLi3ikNHc3CMh9dE3VQ9PM5BGwmi4Pwqi6jp
X0d93nOm1TCh91i49vv0Eqmmkt3spctJ4ivqSZhjjGI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 44026     )
7bPHlHlzVm54mYxUuIkH2dB3P/qo0wjYkUH8GfPSo9Mr7ZHuWdxZrjh4XYjcvY16
9T+5wgqIvbABYVt9D++Cb99HgKgJXt7GiNggWpB9EFcGbVSdAR8WRcFyYEkJMnnI
/1kxMZEVd7cNC6KdNR3Y+crpoya9Ysl6ONOfdKDMVWeh1n1bjFltTVeZaaj53zIL
qVfsOP9KFjrqkZrVhEzUIfP/wi9MfmZ9DImlC5NDYJLhYZX3brnjbvlquJ7NlntD
7+XeaEru6WhgIGekJAqjMFstREF1vVHO4IEa0f82PZ7/s9Ks5i6vAkd7JJjK7HOJ
gUp6/e4ZgY18DAEwtvJ7U9LtwDdZrqpZjTSmU6T3B/iD2SCqEqNRTtBVGceonrjd
yEDzX4wQBBgJjdze25jfdkpTVLZppgtuoutMOV08hPSUpm/5+4yOHyJwCFA5BZx6
u9o/asgxSVCq6iE4fGTNwEcoHE9YzAo0CVju6xsP1SAfd2LoGjqYJDpmHC5mcCN6
PuOCFqMQy1SjlZouiKQK/FsZ45IoFcRZ+kYv+gaHhfJWJPNeq8vLfIJqPyrEmnZ6
IajIK57IzisVPzLYQ/XZN4k68qs/5B7313U1TNzEx8Z7fLOFAcnXWFfPKqS4qJdK
C5GaMQ7OEtAZPuaeP06Um6AzOPqpx6Kg5QlD8HiKV06LHYuF/cGwtmnFNJAkQJOY
apwzvfP2zs+IJAIVT6PkAyJM4Z4YPEfDbiOPRE0KOJPSGUddA46ryILH3rs2zTdQ
ak5g3C0ejEx2xhAAj3zyWFlZ0ZUDMfqiaudFE76NWO8Mn5S55cEAjtBlhRSEPqPv
n0wyomvm0vT+tYhv7fO9N6iOUxaRjpBPo3zH8EKMEx86WE4rz73/xuQoRd2ajJaW
WwuguNb7U1lUo/6ClhAVFZ847pDndvlb+MCgBHTIZpAxzYBWVChSbRJCLm3Yhreq
PS6iWGgsv+y5cW2L3eY3Oe+p2nNm4XN1lEj2d7SarGYuLAiDod2uHU3u4CbC7ipo
BRBUT5eQ1Ou8LJvjF4b27nBY7PLiXu8fOa/PB1squBPhp0HwftPGmX1t8dk45aS0
OQP5ESHbemQfxUDF/UOqGcHTB7FSZ+WB6477oh4xYKVW27iM1g5JY+ASnvSHxmym
8i+yUlSHGWX/4FvEmmc5o8GJCKkNOeTmaBrSVBKUUq5WXNtNi6/xYEwcC+cidmrF
kepgp1kbKMTA9i3gkrFaVTlCMoUg91cwtUiZRBrlVZGLEUZSYcSrLW40rKjyIf5b
kFTPdJP8FjwKdM1RAsd8tQ==
`pragma protect end_protected


//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
MdhbkLrG5taL77KoSWmQNKHarfLJ84D7NXCy6a6PUHKByyPmXmcGCRIYO+YQ0lHb
wmJDssRUr3CA3I7AVuUYtvIv802eRhQYopi/We54kB6LfUdwUe6iMgKnuxY0wkyR
BzfkH/nnOJ52xxn81K66c7rZ0yWlvZhbo/2qsA79Gzw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 67729     )
/wD0V6ye7IADsbK17m5nhENk5+J4TPXbaHcn90vsjECw01lqNjxsk7udMYsnvTLI
jsxZLEXne/jhl9N/igbRMWUgnAuSnZf8gUkPwh6AdsfvMxgEGrOSQTyFPXIWM/rW
A0YlXe13+fSfxaqWbCAWeA/eggK51iBTA4t7zPAchKNWCBxmvktaW5Od8Y7+C3DP
Yd2S5o2p3cVY7WZXc6AVRNNKib6FLGM9+Ur4rANbnT8UkzTI1zxoR1hyRdgg9zUi
GQQl509k5sG0JM74mLyZdQQTnt+1xUGmoD8XGrzHy/Yx3yJjbjhtVnuoKy7Y5OfK
NuILIpJWaiK3hTMN5+uynVhUlCoQiFkYGV9dpkkQ5/COsB3Ju+4d3clre5lh8cN1
WseMqvD7EUt+zdr1F560MzXvYKIH58RsNSM1tazC4egMyvPAwMD27G9ui6NUkRyr
PoavsoZyawWb1AgIMSo/HtvgUb+vzUvwZJ+w8EIwQlzDJnSsD1xniDs4YZdwcmgH
AicCBULbDRLKFIjhUFeamwsQjjIm04ioq9xT7gw6bAzeMoFR6l1IUDkoys1RkHFT
TezJ9P+rV5dNnupUE96m11kJ+MZ9rv8BAO+YVJK/IQdHQvsK72PGi7rnNw6Sme/l
yMZ0kkomrs+/b+9lkjohumuwscjot00LptbIMdxLx8m675sk5f1kdVEwdfQTL6Vs
qBmGXOOPNCpnyxCGfcShqKfLjgIBOLP4dM4bW3f6Ue+15/OOOOhB/xtDPA85gduc
ctiLwjsC75wuOMi/y5Cjmoc8JUHOSS+Ae1o5Hj+RSlVJWWiQ84kDL2F7gFLcxBaL
i0qF6XOKCszMX/5K1atbmUPo4Vp7XBnwT1JQxgAh0pG15wP00uWINLw5yNNhQgD/
eHSDiNVoKYF76BtuGvDzNRIcNVaIty9xQmi7d3gbwYdwO71bVfbC9VRfKHLje1Vm
ishXuuyO9AkejiYHvdU1uqpazvog8NzmaVLHMaY6Wo7rQw0UqghJLccnQaiyzQtj
BY7bY2+wiXiXcFYX3P6BGdCsnkxXtz5lyolEkXnXGyjF09DeunEI8PvxZrdI8CDr
KE49QtNdjrnDJ1b6sbXTCVHiuyj9RWU5RK4cAj8vqgAclOqED5ebLdhmX1A8Ggmu
3uXHXToeGEutQO+gej3R5rRV0qtlB8XICLGFueLrPly9LiIGyXUabKC/v/DY6c6D
fprXVpRMs4qrJEGOTDmR5fdm+UyBA4M5u+Nv4thS8iGW1EOe+avS/n+ZYwq2wu6e
U/OuEeaUgoCSZR0TJoYFoudO9ufndSYnzcLNZacAcNr6HhYPGG9sXSd8ov8K7Ig1
gy6PUeHH5c7d+x6bYcLHfUZMNn7sxOSxtAj/boGMO0+ZekWnnebCdINmh+nBNxoe
/79xMIzbmlZkcsIINvY28dhFoZwQBXPwY2rtZh7bufcIBSPpDt9z6F9PzMUN4Ghv
8peRO4G1uzGKtWAeoWzZVJKdihYgtN0MqUqF+xU+RSQM2TnbaJsmmanL0QUt7nst
GxsDX5Cvf+/AS6dnYWyYHro4gaMJ6KCctrUjasXhVZVyyZ4JfE2d8YxyaFr7SzbW
NAXZnvIHO2ituAsg3CmRsWKCnAtqqpUJzckPJ9Tn/PSwESLvfBI5uDZZGEHx4GZh
A17jFoeNKg4bDds6koSfBz7V671qnv+LGyzZpSWUtjOZLBzzsAAUXL/dPVzWKrW6
fVorW8jNSGHzO6BsPxxcPvXjkxSz3T8O3vSoMq3CFxgYYI533igKIfl3BVsqXnkH
HKcSZzoHT43hecj5HYjoth+uVCBIC334CbaWyTGB+Ox5CNtiYIloDPHdT4lHnFcb
exvMTIAyKhP4eJt9ctpGg7Xlf876I6LaD+2i6/U4S32zrRCgYIYCvB8gXisdWRgN
rdUwlH2jHmT+mQW7zKVtbKwfTXQ5IjoaxEN9aX7SXexs9y3oj5ztIjphgPYYpr0p
WZHthYET7Tlh0t6HPuq0LsGXvn/n3uJEBWEsux7PmKDDsR/xiqKIstrGy5/dha5R
nHHiMdJwXmWo0ngtgxGMC2CWkGLM5s2wRdRHFmWLhQ9OBartNZkufYnhZAHg8PwB
KD1Hb1BHK4w783cjDshPxgaksamZ7Wxx7Q1XcU/xPULslcHLiYHlU72kNKhstFf2
KGRfLfOgcf0YkaGSdWdyM2FsIOXqTEltEAwWbnRs01LNsZLlRQZiZJRhKj0ONi+B
HMoh6UzTKhCT4U88vTOY1GnAvRJfgl6+5KXTKn8VgYol7BVCRDrkOTyRbECPVsDF
I1H0UnZaMHQiyk4JdGCryZFqy9IHvXBIOC6otl8DKWtEQfxeHGAKcHTyjWMPiPWr
G0oVmzMwlCwSJhuxg4hMwYZuGllFAmKGBzoJ45zbDk3eXA0YmW7a3tejzJVcnr4I
tIoNa0ULpiX0dyDJCvEmkvSyBiUcKwVBoBiSKU6Lj4WDi7CT6xENkDId1apFzphq
fFOIs9L59eXIGjFVdkRpyoUmpaEj2hdutGXNoULWzyk6cYHXxQjNxGnoepWbN5Eh
HaSD+gWTUiY2WMLmp+tsMgfXeUI+QuJCTgclIZBYm1ykwy24zK+RUpEMF2vVvC+b
7DZTbytTiWHEvJcGWOs2s0/66VMgpD7EBOrVeWDqZITLFXJnStqg3zLL+6vsQomu
Qfc0HVlsaYb1LIHC+j0Pl7oaIF3C+tZc5T1zvQq+evs99LLfupUvXSXquVYkM3LF
OqH6AgY5bphv7ryruchwivb6OHotXmGVzZYCvATtlXtT4XF4Ra7RzkudKUqrfqYC
FMeYdr0jOnXZanIvczMZcClTSHRXNrgFwno0fSpVSVkd53LCiWPo2+nYEYeoYp85
03hZynAiJ8d6uHW6XbueI8CV7Ok8NEQznoiQjoKgC3SWJz/tcCpl9I1hSug2sRxO
fVgoIZjE05qEdScr2RhYgf70xmV4y7Lk/4LcVUdxKdnmtJCxX9a5RvwBSlfiSbFk
sNzFJSBCdXz9OMlhpuvSzYYiLvwDHYTM02LeQ3kcMbi4hjL1pqgejluAwHI3TP1C
n7RiGzS8NxTw/zLgCr8I4EThhnTY5h9okqUT84PgC/vpkDruAQf/xfbPBo4+yHVE
K6mvdVENCUsXWYpLn+GlIubMSOx5uY2NxrHB3+DKznoSekWN1muo6GxHadNnh1ja
8YiYxD0LFghfX5eK/yiUH3ZC/Zy7kshp06dQWdZ8MaHBLj1ky3Yms49gfSBrL9f0
6wBv4Eb/VHQizkNB84B1xHB2LHdpwTvfJsAnrpisT+uLEidqj85L9GSrhlDzyhkk
eKWffLPDxD/wiDrdm/uLciOisvcQVg3ZThHJpMtsFI+vtex/iCH0MfEb/zcpxuAM
hQDVNDzHIZe8wDvlUGRtaaFjYCoN8Eu9p0i50Y12qzHGm5Wru86oy90M/o1A8zE7
0TJRsNHElJ8Gsqv0QZQIJu7Cvdh+5/1JwN1Gmc274HdwkXH6SAUIgXLsrYHI3u0E
TkbEP7watuPCJPcrwiV1zrH2Z/Q+Y2BNeFuu6lFDb3/wtNaXoa2jja3UuBgsCde4
gANrDe176p36Z4U2J800v5DVe8c0WUQrWOvI9+z1QwN6XH+1jg7in6/cNkDDY5Ih
uQjx87NgLixyOEErto8cm/Z3QWFoYIdYKBJQBeQR+aymRX6dbnAKRohLJHdpMe1u
DOIuXGQDXgo2r1IZFmhEpsVo3zCZ5UwfPYogj5IXALJppqXlPm2Msp1QPqYXCp7v
YhJwRjwd71jXngwSW5m/IiL2ZkTd3v+GmukkCyt4a8XYakMni2Vi1CoCu8/yONVg
/64D2hQpgjdx3PkHPSnUdeBmuikRohzcPsbfMIlpedUiu/m+eVi5Rar/A2uX9vxl
GF22+Q8Dru/malP1COJAwKjmKD1eTyyTSx6fIjnGUFduaOc3SPTc5QmGEbqeMmr+
RbWBscfRVctEQ7XtVRbvCkL3laQUMtRuE8UZbnVbEuSV8BF6kSdsa3MEPn6bc109
p0005Ny6nkofetvcIEdw8RKkz9wDVVAe6ByL3+a4BbIamKEC/jezZuDv/fllhK8h
kfSBMYgisdAc38f2UrYWEPV6uA5xqEHdb5W00rROl7M1EEvR0FL0pg662aBV9u0X
+v8qo5Yq1UaXyo5gL2b4NPTU60D8HfkqBpHM/FuuizxbzzW3lEMCEe6SxTiEHbMV
h3pOBg0sCE0UIba5sB5X5s2odNBZSpYxiTDPM7o5yb4oH1z9WWC/9KK0jnXYquTz
YWTRuqYOC545Ux05rmI6S9zMa/07E76PA1Ec7RbiKBopnaVllGEZulZuY2bpJe7n
qku/sprKeVNElN9uWtbZ0J6+rIQbGseFezs/UfOSjSjM00uGq3NqPydhJFLnGNnN
RHOjz7cSThPnEbapX/BLPFpmZ3g9/GfDIM4rbBCXSQhzyN9DQ0yU187PvzC1z9TJ
vqhXuQ7leybBqE4eWGJ2piSeUkUXaX2bkJ+17sdi+xqSVgRTIndZ+OdtlOEsrpCx
/RIe+iJsM5XTq32RfI7CZrzOPwiMH0e2+lrGfaYKdihf0XPphrReQd3QGyHxdDY0
xRwxTESbbkWv5CGh2cUJzEPzEIH7T6czFRrbla/z/ruWblbHg8GipjJXC+PEMek4
PyrmMVJqNsQoByEu4smxY/ooNaq277BtP3ig5w3RCwUvgWfp5qEpeiXpexBMvZYS
Z+R8gTnpoYKiZ3tvtt5rLqaQ/twnfHEXJJg9eyv1mHW/MF1kL60EsfM4t6/1mhQJ
W6p7X79Q6iaeEiCOntRx66Npia45rU5T8ClGUoErw/wWld7csyvBOZ94064TTw5X
SJcYZLrGpLz9EpXs4PjdbC2FjSqxk/tQxy6SennDesIBOwFy8XKcqagUiHqCpvgE
7Wi5VQn82C3BzLMlYGIi5s63X+2QFpL7lV0uG+NOQ2zXXxH/5BwS1Ix8kI3p49yX
jodMlpyiHEY86zlVMhIW+FPfoazHYHrKMjjVvxbdB3wRSY353BU2XQEdLuXrA8Dj
VuU7ddgQO+gGeuU95dsrSmYnQZJA2H3YY1N5V9o+DVvAviWDPLBWcg4/PNq4YQ/T
ZNsNC+L40AAUSOU1mFke/UcsYBc/HHcLIt4PN+5BWJiu2GIQohiUYO3ruipXW87x
Cpt9SZJfOR5Y3Dvf1+xuc6TyBs8PXKGQC5p5zTZwwm2zGmCoNAi489BwSu37Kb/e
Op/egvyRxYNtll0WnJeDfO8RPQ2R92uPN29XlKe8xg9pj8KmOK7Xeq5krSuUKLkq
b0+E5PcYjwKQIh6eNE9eVJVHItk1wwLNNpuas/hHSGJtajE0+hOBfl5T7a4I3WSV
/L5vqvgCjQTVxCbeScukmSjVbVoPgB4UB+TvbMQryQg9hOFh2o25VWUDBpBys3UN
Ev07BMkcuEjwn2FborWuUcevjEn/dRDuGKPoVHkbMUxeOP4nLbcQpWC7QIJwXmV3
FXiitjTGRYCNK3ds5QMsaCzZFtYI3nOOpWoH0grs6F2i9q8AXyzaiG8Y03XKe6+0
6pQ1DRPzN2iaWqErO1rdQyUS3N14s2hRNXd76kRm2DhSbSiaZs585Badm9/K2IzT
5VoD3N95lu+AeZDlu+Z14WaP5oKqG0y3oP6QBsWUfHjSnxKoaEtCfSwPiLC/3amz
aZV6qv2OumcPxUXiDO3xT9Yz5Q1C0Lsr7xwNcaX1C/g4ANpUM2qKL3qwKVnJAiXC
u/UerMDaljA2X0sQEW35cozX/UGF1dKipNgT944H4AkIkhxY4HdeONPXiqQ9G2+g
uHKIrPuuD/il3+AFfNbwFQYUufqJksu+IIXU/ZSzVYp4HiGW/5457PzmmzD3NJ4o
R9JsKNXqcCOqfYuMrcrwtjO9tDiHtiuWb/9gBrRjkdx/xuTUQtYeJCetB4uU073e
sulhCTv2Z2cICJwLV9uFby+D4Hi+HQP7ibkbZwTwUDuvcibejTPQcXb0PNALHs/v
npTOUyiHK1T9Q1mBTHDEWVJNZZ/sbNXX/Ikbf7F98KIc6U4Qdlrf25UorGS/SFuE
FdyyuAaawdXxr0YX1C3gQAltHeTTIvfcvrQKFqzts5szQS9g8/LLUt6cpvHaPZQD
JxM/34sDKZThzwZ2w6KhHktRYPlxPCVWFS3N3X1qeH4qc/TsreQh99SsxvqldmFd
k6GcNeG0S+lcnfLjhxGCgugUPdUzVemTUj004qTRWZC7OTY1o6RswSf8raCdBPFK
PWHl7idhBeGQ01uqUwzXmHIyvLD4oX9q1ueMtskQwKlYqDB3RfWVc4GTCqvvfQKY
kPhAs1bbEd8dEsET/Lj3dNBcBrlWm6nizWOCgKs4t6N3Zi2fF++4EGcVc6yO4p4P
i3iHAck1O1wwwmO8e8jyLg7dU5/id4XaZMnWSXI8EwUU8VRApfYJwi52AQudiqTu
cfQSU/4vvHLOv2m5+DsYql1q12jPlkt4s1mK7sqrQigkO31o1VjMntrkAz60/Lj+
stWZQ+sbwiEAEVNvMsRXBJltGQX+JXR2bW85a0vUzVIlDn21H1hw0sOpflmoCFZP
o87VWr+osaBrCdWqyXrub2Y/eLlGKPGHUBfd2e27K/pZyff0NKUrgiXTji9eZ3Xf
VWTIjRApJQx/lN1C2qLpVWg6CHl49uAogKjYgvAQbK7m1vbLMUgRC4jFQwb96aqI
Myxnj4LSwtz+ZgZKPSaM+QIROTr1PPAhMxhyFbhUAOjwAIAGROC1vM5jxTODmO+r
ORvFL/4OUs4JIUNF8UWCH1Iz6mhO4vN++1a+Fm1STnBXYJmInX6w0cUduzgPVxOu
NFda/V2ZISONQHG3R3EoKTi0DnTdLLMgEKIb71yuzM71VYRq15sqxzfDhOeR/C40
0aY98fDJFYu5hd4AQ+nU1oPTMKSt/8Mqvv/CKD7OBk05IPcwL72h0vWBGJjO8Nzd
HMJGqIcZ3TZZq/tWMDGXoMdeoSup4NoISJVDs3IGlzUtRWuLWHHkcdlg/q0HVvTy
KIvVdJE2IeUEfLNXiTDKDtCNAhB0SsDvmTjP/nQv/2dEB/dzudF5jWDHdgHbdPHg
zq3tcTuMy1T8tENKXUU5jikvee4twcxYunsRw6kqZhTtpdtIaZ5dJiM3bZy+5dgb
efMYELtR+A0Rl8x6exsCJJxyaQzSskDNCr7lj/K9J53bgJRSpvZVpKaUvJJLzoKJ
HQBVhLLmbDnC6qECGhedE2k9c77GCVJpcFTA7yVEnrKjnCblbknWoTiDmAAjBv8I
u2oiHElXRxZOX2fmy/d1dA1fevvK0FdfxIuYTseD0fHFYG18SX70SDiiOtI9hxUx
5pMDyW/5ZaSiiUzWlL0sdlGloN1HCJQXzGLRVuGJGVK1/3eweYXlSAFOlnTzt4x8
Dl066tm1XJOmh9tRaMenxhK+9hO/ky31iwgZaJp9p0woIgige9ERo8bXmXbqC1rP
gaVM4JdYFomyOzzqBfTTtsz62w2Tgt+KKiuLpePJxq5msh7Py/fFC9NcEyIhPD+q
GT+wgIsK6qvwEta9/2d8WVtLRcfgE+8UwSK+7XmCUkUMqBJj4hi2hJvoD7l2P60L
YgBKxssDcz77MnPMGD7VgHr1oNsVjg6+otDyUAGvVcIWzdv3HIAnnqNhv2v9zib+
ZM/uo1exWtRjqpA7yKVMtUzUB2hPT82VvAdQXnlMh26WVS93PYJNTys5A0VZ1CsP
rB6/MAtHmjxGDwGKRFS899XKJict5KnOZfqCuAUC8NzqB3Z0AnVLiY51nqEPE/5G
DD2Xiv3HqECZkHEVKKm1J2Zs4RXljR1lpJ1TuzIlVhx7HmQ6pzympKFwTsLqa9vD
P1Kzq6/qQxirZT1wcxGeUUVX2OrJIPD4aJR67v2YuJ5nEMBFwVVw1gLr4ZVZ3MDz
6F4pnBmOtjZRaufhCgomVXmNt5YEum5MNUs+ULlbgs5JmHE48IrkbEY/0iKscFdA
A/UxtNPLLwORm+lip3a2I+An5AYP0o6aB9TX8pG4HshcTV0NLMu/QsTnRIqZ4Au3
tZjwuMDESvg92XqjwHFM3egwE/vqb2vehVPqFrQopsGEr8AyXVvz1xCg4hrZmWoX
s3ZZ2PhVPOo7QsH+omdZG7N1rcvBbkjPih1SZp2kLv+ekvK4lqXqXMHwHCKgaBrJ
s5qxSIv1YydpH1kH9kIOOfcQMvzRRrzbPhPW5imNVC1mjqJt8Oe06NPmMTtjF3Gu
Uevkr2LM/3Nah3fZshUKUiVPdy8FjbOyOXo5BNb/3QtE6e8PfZULW8bKeUCG9B17
+DmX3gz9XhGClTLIpHVteT0mTlmUn3v/7J6ke7jEj+0IGAahSjRYNHUH4QDalH56
gDt38O9H5n+WJoyT8HXcYgAMNOE4UT3LkjRHdP8E7WcZOup4LahTYCyiMFMTd3bM
dgyACGc5i1sqyDvve4J0ndtHTvJ+AtjrmXSSUmGtgoYYwmmJYJ+o3+GsVdAbpGYp
sC2ge3UmX+4gc795SnB/NDFAnWbK0iDIUyITEW0jJFFLfZxrgdHx2OLwj1UjMykO
pHEYdT0bUlUYnePujlLT/0QbJUJaNEq/i21mI3ZDtDti04XbFuiHpuxIbxraBUKn
AhftSSbyD62nx07gbfI5Vqbgu8uvSo60RWyv11YK3TceTj81Kzx1nMgE0EAUeVGW
27dkHnLon/ITwpXY6ZWsI+/x+OEh4cDL3hIqTvC9qXZNZ+ndJTLDN5ErrN8VOSFA
6tETJl+ii9xviYxKHIfKUsSto3jbKk8ZVB8l0dBO/ADNHl3dS5+pR59CJoxd3Icg
Z1OCVRqDJKhKNBxEImSys2mVJ59fZGbtX1GlJjcVuQmcyFlclvbjFk6XiRU9/kdZ
J7YM64YHw0OygzVFkWSPZopb8xTDmt5x10B2ga2t0jGYxDxsO8hPtqXM12n+WP7C
AosIcS67VrT89Ef6cVXoGkkx8jqwblnrdfTHGSubMLjXz/tb6ow+S2PKh9hWF68x
zLlQl9v2Gn4xyLpFtqrW+RCE0vvWmHbNR4wLFUuzbBMoJ0APg4QsgW21DDmx2ocF
l1rB5hMlNMzPtUqPV5Sk6FqRFjLyDeK1YFDsi5nou3ov1M/cD/4HEyZRbVF1NCd+
quqTx/K1zixqlvi4q0DJ/3OlhBFIGshYWc6B1dApLsrjLFK0LGLukUPmQsVycalH
KCKvppsNrDBix8txHaCUy98O13iiE11eKyYRl4c/lpdXXEhTzGBatAzvT2/MZpZE
QAn99IO4sU5q3ebstqScvEllDorsgfIGAG7cD0ZM5Q/4kAIpslzMK4MprOG7kHiB
b+zE+su07gurki6FU7oZ2FsJlO9ABnF6+4XJzQFGRYDibUod4ROMRMH//l8sYdEv
Eg1HFAzCVzSWpcTw7gS4gwPcHB5okWmfooQ+E3vyMfakdbs2BRLeAMvsJ0HKSZin
KGvtrYwP+rbUIq/xTQJpeeJACeHNiAG2c0lnGNAZcOj5WC1WFURyhOXZFdF3N4Hw
2azwRQ925LQOvm7Hv8DKGscKm9a+wlJawTcbPbqKWN6TD7bKwp7Mfg06y8Awqc3z
/Jw0SzgX0MTjHZGHhkSmqA0URcD4LakRlw9GKfjGeUD0nr7d7T7MYmT3+gRDiHXy
H/9Q78UjNAB5+w8ACQIGmIzp2DL2gmUEcNAbvEZvSWMKjKWezdIL/Z3buJ11oqiD
dG59GFGS90oP+tAhXxB7zMK0xpyavy2G8rw/vSYQoNFCx2CgjPaSZJy/wO//T0bh
DZgYInV5EYZMtoFi7VTP9ZI0DlkV41SMkPx7huTWj7GMl5Q8BwASUEGcc+6rr8Js
Szz72XDA+xxzIajpMKmp1S8KqpwweyukXc4paAmSSIWbyNC6OhF2tY/aVDmpsDaC
SGcCkyHGvkFD6EiI/h1ZzRejQW0ihtFX2aOWLQUXzOK4Kq1ePG+FxM+gLUcWpdQn
mjqJnHIsFkk+NlZPJiT8gJcG3svXFCRsOUreQ+EDiDnJ5y6knUc5lSrUGG9+37S9
Xqo5SD1SgRpfNQRUZ6vRZoSt/iO6AaCIUHcB7Cyrc5zsL8nyCT4ccp6Tfx/PC6o+
44an3nyI8DYsVGghgz36Hus8KlmEmh75hJ3hNpKerUK0en66K7qRlgbNu4+f2uyv
uBHSVVPFVPkZDO2znkbjPJXNxePu0+Cna+kDU1gtYH5Phm+1YHJvYybGKtggM0s8
0yZSj7CZNS3NLjmvBMngvodoh2e1Xb1Gfju6/bFWYR7o4a2CfPDkvZxYIDQz3Z76
jk9RpznmQHdAhMk+7BVtfjfbsz1llKl/q0ZfuZvRIIwC78KbqgIDI501ofkClEbr
lWwHf5kEudmv5ung8T7UeBFGDU7HeFbaOEc3MKg9+IquoORQaIRQlJU8+LUizzAV
gImpk1PKphFhac6GyDEx0CVTCfSKHmaEN0YNysaC8LdJ76GZnYfapTuW/arpY1k5
pewalsh4InyRapTZXGLBLDBBorxDcPGthpiDdACAFaAxKaZNyASLvkg1WiYVMw4e
ys/gWjKiWy6xD+ZPhsoNzfZrigeTAVQ+7TxKkai85aTxePAyo+HEHXbi8oPE//EZ
ZE5LyVOacaK1qkDILU9Z0PQCKk/8LTLbYL1z0Ytb2DVn8szsSP6gD2a1BVqiMyOi
l2rS8iWWIsp0BYjVEJJdSX+dV5gRjq5qcP7QsxkVWqAMUT+cb++5S8GW0WeFoD27
Mbad2rSzdKqZ5M47BHwRuOhCvcmRk+Vl3GntysO8l7uVILSTq+bZqgmIzt6OG22A
ccneCrXXZtI5F0uAA5fWvHliR0FwJq61ge4uDKdbEgnSBrhkVDK8akxQIkcnExAr
i18kHvKQggSpGb7NWZWHOFfM4jUrB+n36EBNNXBASM7qF1totsfwhDixgy367oG3
pCNur1l5s3jE01+UbsIiamUQBQKl6LOylzluq6X8ATpsPh3sjTQN/JoxYUZjX7R4
iO3WIk/HHpQvtm1Wf/tOMcEA2vG9IgAg5Ar3c40n2GesHGjpzi/YNeeDRQIIUat5
Z9o+0+63WsO006VjA4SMK5hcy8jptHLgQUyrXOoOfCahPFtQSdbK1j9cbRnpT8zG
VOvyf71AAH52nowHN5bp74oDD/7IB7oTi1mtlFepRhclB5XlsPppvjqcHUXHvKse
yKQd0UKrNy5x/o/LMx1DE1pzfP0kRDL4ltt8/4uG5rpWGw0veqbOoyRgF0wPVIhd
M6FD7wDpPtY0xMXjUE1x4GT+VnqL3yN2nuQgN8vd5f4vgginUgyLfEbs7FXhOKXy
PTdmokrKWFSIe8EbXnaubLRjyKpqTjWa9TtkXWGQJZ1ZNU5eGTxhj0lYWwTo70xS
iwNRAEsX4H3FpDwsXdRm0zNiqIlsjYuzzQ5UzB5ePUbEo7gQ5WMGlcHLcJLvp3lU
je8xEqx/i/g/m22E9AAJQo1/YpQYsOu2OWdZIugtp7cemDX4YNUZosWIKEbSV5xA
Io8Gp1rKbTK1o/TBG2BLAmVx4GwPIpQVDJS6xCDow3fmdEFGm/VIk1HyxNHx/Bqk
I/lZweLu7dT78A9uBR6LVztAsSgHN/Wh/wgI1uWtZ5IpEE20+DMVLIXYdmLwlQni
xO4riJWty7OH7cb7STIUp4i4xLiznxqoY6z+ZpbyXq+3eqBAORq2e2kyxXiYPwO7
KwA48ry5LDHp5u+yAzuFiHNPUUOq9zo1fs94AiLAHawxJ9058ELSHoT4GNPs78P+
BLP+bcJ2ne/VGi43y5PtV0fbHoRpPWjou517oJ61cfZNpCWi47Cm9xRUDBT6WsZ0
/TZcII5Qpm6hDR+y+Lv/35S3K1YEhaMRdqXMYq9auHRVdIGdktYQwdBz+yQRvqhL
t6h160UCS9K03ufO42E0WvbvfhPccImsPdL3Jk8O1LCxjhJ8PaYmka2+5yI3UFHM
FmkPAEN2GXrF0c2ZBq0UwdRMrdJ8YyRJ5B8WGjoxBWiG4+IPhS+k2x4wGrSmFbdA
YlaRocwoTTCx6i23ZHauVh9/mD25GYym8LnkiqXKNwMsVRbWtG8nsem+TC1jDsE3
gwiG4bjD7Ac9mCbd4IBg01uWC7pMhaCwFoyurhokZPYNJd00NNQyEWhTkL7kSxx2
o8Rhg9nxR8d88tuSfj/gg37+Pw6UfMdH7XUOPr25j/sBzAAMoPY3Ut5KKObH1aVo
i4AVOmdTZi9PkRSausHPCoN6bwRpmWd5sSi5xeP3bWDa2TDBydKDuhBHBF1vrJur
DazSab8rLEUWpvNkwxx1/Rmkprnf1i85O4o+w8CfaZGh4/i32vd/L0+LuZjF8Ye6
K/r509gyGIUEzA226Rp/YL2VP0KiXU9+Suuj0uZaQycDoIuTN2yG4LP4PuS58VlU
YtMZ0OLvXbTDfR/5xTbhOsDdrv8DYR0lV5Gw4N+iCyGJu3i2x8wa02WOSfMRa+Bd
rBzaYx5s1lUbCLYVrsaEBCHp7JMKdyXd807KF9RfOTk2I4rXWwl8oqcrmF3Ziee7
P0gcrqN6IAoFlbZD1nw4BJMCMmq5XKY66HF+n/YlRW3Axtm2hMhyIr1XX1lWrLcN
4Kf3ERZV6kowkANa+vBKhSCxZcftDBOTwXNiKY7prXA43WUAllSflSn3VjvNsXt/
W0+Mm8A+ccsCz6JKIf4BVEK/KVCxdKZtAKPc0OaYJsSKUGwgtc22z77ltAuqKsfl
3JPzO//DHv2JGPgj+h483wNEgiIIGZsWvxivu+0qfrqG9WiY0X/xjQpVODVZC2DQ
GJURAubZu6MF8J7+hibQTjiyBtHTSsJ+tBI4tA/FSMkbTMeVODSqZL+Jqk76vfA1
0LEvrvIxmskTXAaoQau5VmIKCxImMD8Hc7QTncvLWFyBvgiQJ/wgyHFnnF2WLfTM
iaiveBYccHjvfuSZWwO5vZqfmGz8JoV2TzMsi+e5awsVr8bQ6uf2nGaIMmY0TMUt
23ErbqOlXbLPRxiDw4sq7twlRv25NR+WJf4wYZWAL2daRupZo8mFqr94sv1GbdeF
g87cyUnXL33D2oMcwEVjq40/9fa7LUzomcM4eH3gN/GHl99CCM71zrvcqvSVYU4e
HBZDbRQNfZFXVOslMGu3fycEh1yVl9vKcAKMOeQvWg5DieaWbVQl02S4ww7LRtK1
kNFPbg9HK1OBk1Yf9P8rbEHTSMLH/UW7uFTaT74fhO+ff9jOefDrGl+SEA4uEJFC
fUkVVZ9tmwNmBt6bllJU5VBOBEFOOJKt3P815DQBAQsJyAt64TEGXmpRl8q6MmzH
nuzq9+itdzmkCQK+/jtKKBAuuL4Ivzbf7nmkiMo2ZElzRE+CJCMK0+0iK4VVHQ57
Hv30boX8df9cSqEvL3N+wKccNE4QfnRYApxbn4OwBZqhYpghSG+qPy5yO0Cs3WnA
M+o6d+n5eBtBI5g+KDAdXlJUbMYxEWrcA/zG1Zb/D8OOIKTTPqMy3vgHoYr54qQ9
k41Aj/5pI5KLW1le7U3gUvE13UOWLUxZvYBqLeuzUKsORBfMZfTcK7S0APxAzPpX
LHSTbuV0IHBjtcpXKH8hezt+2W51AUjbPYacUv/BEwt5fmjAdV3hxduDGNcIPA+c
hOdJb3lYGr8Qy5VuJXcg+uH1Hu8rlRTPjHjmNP4znv/FH8gr7EV57GNu/KftMEBs
uc/r61WCzHW7ef1o4N/8GJbezp+16YC+YNk+ISFvvBlSKh8/jeeNPW61SMP5Xijw
sCg2GOUHVmdACRw+3wLNV8e8ikrR+Czmsj7LwHjc+WjqncvVO4qn2NQPcvVLau7n
m1umZtLTb+o5Uqt+Rf60FCMSuZD7qbpwhhAEdRdwleu8pedtV2L8m6CKPrZfG+Bq
Mj/OhLkpSIUjs880sGuDGe5PGw6bMSG8fLwpO0EVxBR08I5mq+s6Y+umtiBoPZRk
fVS7ySW2fkUJl9jrWBF3SK07MnHPs+B3gJk4lTlExCQ/lk8pnL5PUelHYHSd0wgC
WVAtuWKs5FlsRNO3DZQOJW9iNH1UwQVZbFmsFzve6li0kyA7HSL6dfClaJ/R16gn
ZuporN1s0GwCPi2rujElXFKh7ec6X9jr85lK4Uo/uKvauJmLbx8wo9B0XyS9JyBz
ABtlq3JKGlasJVqqjYNwp2wkuW8oWztCsna8K9GX6ctULptPFmF1O3s7yEG4mRhg
b4vW7Z+yZhoIRGjDQQtT/38SorQn1EAFnDNn0IiNokON2AMWERXPwN6FZXXm7Ci3
I9Ilq2t8Cx0+CxieuhSkwysejv88wHfwPvLx18YMkA+3ZXC0DQ2Df4C7G3oZHibD
UpcSIDuip6iSyfMhER4gcBeSBHQKvaFJ90Re25UFU6GQXLyiH6kzGr+nbYBn6VUv
BeB7x7S8axNPNh+1dN/oJBCYJf2UY07Ci0iidW1yBRRA6RYTVmNkjgAZtmOMNJQe
6wQYrxSLUguYY86hd/1FojqUIaB5mSzdKIqh3N3cYbBtsWNwY0U/vhj5WsMLXZ1a
iHxiwGdJaUW6+pXrxPOq6G3qPu5nitQvigu2ENj+IrhNJs1wD6OCc0KgVgqZFPLc
98o4jA+E0Ii6FAuCrNsCMbUUFDc0y77YD3P+v8NuyG9fpVbzYcEGVSrtqECASo2F
lbs6RhS2meQHyp4tdCW6izL7tRIha4cCALCU0uh5Oa4mJRbAzoLKLxbt6bhUTNCL
C9aef2GfFJ1rztV2yrBnfgJnwbAe+JZmsnMtWrwuaJKy6VwVPjzl9zG3bUak/+pt
JTQW7o/j4dJHDlkFcVbGag2LSsh/OR4naGtfz3naBTaCxR66S3BkK7DmvsBis/pK
SY64z/zXTeXyd/n2DUk38QgjKC0jIBV4usUXVKgdBrvp0rF2rvx5ZLFAD/HN43Eg
jl4aAznQ7EUxPZJma5OK824uMnNh5W2yr5fjbPxfPx5JT9gFkqcNBk4LF+TZeDbh
2MVTQYojsxcrsig56Yw9cxbVq60g3P0JjD0e3JIkpZKS9paUL2KqAxSXxMVX6Vu4
84FK9dmaE5UGAuvj4xgqdzRC8WqVktsSynZglofU1N1LH5e7sG3Gve86gwwhO2AF
eZGntghdTaE3Vwj/IaJrW7RVDM9f46duaBXrZHJIreu2LhFxFpQ36LBUwdCzBuqs
zNFv2R+xjP3uUn0PusbcbpJ1kLK9xZQ+q8EQX6PINy0Hqan3S9mvTTSVvkagAEoQ
inuvoVZgddLCbs+OsvfZ4nQKLmRcTWG749+h/0f9VwdN1kGpmy4bYHGH7AEXo8Pn
56sJgX4WHAQHiExXE8Q4aYZxm/DCDlFCdj6SRoIqCG62ysH/WNUCaBgL8rWsUGpr
IcjY8icjT0DSi25beWvUaOxF3QIfIYHSAiZ7yR3UTer7paIOZ4ZmjFOVo+lpZGCb
QgrdjwFgIxs/4ULMqYIm3jhaBPEaNbYVFbWcF21fSRvi/rcmTAN4fMe3bW9++Ps8
MALJ8MLrZNuVQbZSgNFFN6LtSE9UYaWyh8Q6iG0PF399J8T/zgukNwJV4MG3knOe
8daaxJArYZ9Jaa4+3m8Qd6d91ENEEXNIImglYKpV38PgtmsfF431M/eA4OQu+YmD
XQrYAQhvdPMEA7qe4h8QPLbNVPdWAsxUORtmZc/wklz221SQ+VGbPIkAuZTU1U9P
bcuM+a0WD03rEAtWGFAi9oRsXKUefNdoQjKq+GiE6P31PoZlYNZ/L7Gkmy6tKDm/
jmPRl2bBV7hCijklxblQ0ukWU4SDNFDdMYP9e6GgiVzqFsm/UCgTgeV0rdm8IKmw
ZTn6odo71zHGARHZlEVNuDhaa0G5K66wKMOjPV/5psomjxPx8PR5QSLCKslpbyZL
yrGgzbOVlpWkLtWYMCUKgmKdInlmpek1Ia+BDcBKi2jVeQLWLanmLV2S4O512KMG
1YFv6FXbXwEN4ZBG93D7K7jO5HOnlsmRGcgzrE48UBAB/gnNPsHj1KoSIHOp60qM
EYf8/G0sEXGPQaggUVheGeru0z9wuFrWFXyODmB5pM0GzxV9NGFLzSooYp/0BYfT
Pb2k7Dan8knX9X6XruJck6re+ld8DBd9sqvF5/PkR5CnRAIpcVjXirvgfpUJ+/UR
xKLhr7OATZCx0MBs5LQZFRPssB1QUwvVs7W/8OdR/dP2O8V9hJgsGAOkG+nsouz5
59Pw+1xdyD72G3CmgI4nwUngXhvpMBmYEehOGNrS2/DYWYHptG+UN2NNHFHfp3fk
lKm/mJps6mCMxvYPtQi5rGUeD7kXhC6Yyup9Klb7vXOnvcpWJr488Qq257A/Cn6D
GLKTUmqPk00R/Iyx7D72MPbEoVPLWBhWdG+cun3g1zbXDvuAuDoj7kd/UyB1dAYt
pNet6bJECB4pjeZuNNXAIQ88BtB+Tg2Tl3KkK+BCNAM6pSJwZZtCg5wqDj6JX70K
8gj/S6epcmEADFLNKv3NoeedC6amru87Hf26EK2Xcxws7DsVaSNe5xMrnuwJXUja
R1xOVlnj5lg6q3qH4YQ8MGCAnF25vWE7CnN2daRGr79C0VyijbnlAtvTf95r8PwW
nepZ1YXgToHM8Rm6UN6tX82VtD6bbCrbkLWofYYWfKIPQTjDJnnDi/ZMSXwGHne/
uJM5M1lJ5oGIV416rgk0GRJg0MbX3J+zP+oJ8OH0ycah7VEsuGTK2z6jtV+80cjW
+OksvywWFdX27VFTw2zhdie11vg1idfVbadMGMf+P+5pkiIa53zSO2AtkFxrepNU
G4Pya39gTXnvJvctHvmA2kOB5QAN+b2Ueis58cMT61dXJcsMb1L/pwUHOxqXgaZh
qGfzZeT1LwGVUYaIpZx/TmVkJcmIPDiVAJIQyFlz05DPDICGDBWfU1xLc0rqlff1
lPYXA64cUKR47os8bBXDvk2jpVqMS+UtMaQPI3EQBNNytMpC2xLL0Znrw8ifNz98
iyuy7gzOjxmo9QhnfzDqPIHzxcJsqQsJEL+cwe4YIzljoPb1soPU7mXys/uKb7D1
Ch/C9CjMNsqa0ylobbvdkbw9eS5WDoP/R3Lft5hWTB3qQL5LPQK47QuCiRdQI+Pw
AhCt5HUVCkFMtpOvECexDEjIQlozQ6SojuigNKH0jyetKZ46gHMeiVlVyW6gGLAo
3fqBng5gGblg6nT09vDl8W36E565wjZ1m2tz2y1rnGVuGB/wLAE8iyQ9nVQNl6ld
5Ka0lPVDlTKHaZY0tEKf/KJ+S657WV0Yz0iu1OHUhs5nZLVJ1e8NKwUnnT0SIm//
gGivZfcpqjzZYNL9bcwCZuQunHsY44h2Qnghn2DxL2QsVLGYyxGtX2JFztwc/TIH
NFV50PaoEPyJiXRBYk1kpUP3jzreiP2Zt0x7rxTHaVcP2ZVoooug9Yk1njZmOfQF
6TZF8EN/zYSnGe8n579Py255ZcFoA3vcoi3PlFtSMQBQJYPvYa7OpS9wTtqxQ++Y
AaAOsdsdzkQmtjCzL5adxsBxymK8ewQulW/D0O+tGGkIn7mMa75If3ZW5c6amUXv
PCZs8jgAic5R+SWphq/1YiQ1yf8rqkQ8Dq7vLMC3V2JWzLzS13F/owIjgu2/iEy2
sO9ChK8SNsR+0HSEQfjY5Ui7gOwH3xM09dXEdpd2EKUAUUo5SNMLzr7yp3Ap4uxG
eWxF4OJxAPVJBQmxSbTHGBk0apTHTQVFh0uc6OCScZVFT8eCtxhXDw4pzcJXjx+q
mx0ob4kFw33Gs5YANQsKCh2pbbNPQ+2IWni0FbYIs0ucuUx+493Np1pekV+pudmv
RdOqoH/VDoa/NGYubvEsWrjYmTnxmt32Pg2gai0BtcvhJ1vFTknFuetknDUG6KZM
FB69p77m+uDMcEdKGyXght5Uvy0OQhoJgGCJvO63wyjxp/jYJuvP9uzYaw9mXIYs
/OIvvE+KfNCpdjKFA+JT0ZNzwc8rVjaGGCYSNHR+LSgfp4PWNa/X7PlllpcTn62W
d2r1jEmRWYtMGHFw9ekf7uV91jJFMvOcVIvkNTSktQb4dpL88zZZeLI2hDceTpYS
i1x65oVdM8J/aKf/edpncNZuC2UZRvjOAlLufQlrxCt985rg736WD0tjJKSKAEyU
UNLUXseHKUjmrwTVsCd+1IpviUPR/e9lSCex05Wu1lnMRudcaIpnnADjmzjWPyEJ
+kb1tMbDsFqhEiVXOb+WUxlhG2ktNdJewFdbR286JwwefMVhy8PVj6tTodP9Q/0x
yKd2m5ZjfradBA4G7m8FPIpbV1rHFDE3OMus5Ci/biMfB+6aYo+id+D2ckiKEtFG
FKaSr2Ij4uOInKxNEssCzvj4k3ORi9PxFUlwTu50sliZvEJD0dYiaDhGgDuz2ve8
YbuQ5pNAkNrIWz7ApVO1nQZe/OrfkrBjC/LJWGiiEtF9/Rgsdc/D/w9c4LoU756M
6ucAX89vW1+iJcpB16b3QpWzsEN+5WKeFNvF2IOKJR5rgHoW8BFSRSP4XdsZOKCF
DsRFXSgbFEy3O6t0O9m8Gsfdain1PvGoD9Baq5BmItvX5fr0o4fbLB69wT+JQzA/
9pS++hTBvBk/JHo7nVpi+0HuPdXHtCpKZ/puIB3IRIC2CJLegj7eHKHrBLULA/ov
F5V+adWmEAwseSpoLsfmLMtvneQ+pQrmLS4XqWaiDnvpOUB8jApopaVKljbyWKUK
ffyNhZb0cLQmIfTBK/sNUdkrCfuWsjodHslUw1Sw9pTswMhJCX/Cx+sft7MRhF0+
xqsNuLZpQAPzaCPh0akg+eidR++k4YYomboVXCR7YzfyAK+0PPzi7tdTlGKW3Yn8
5o47QJUFIgbdBCRbusp5Yb6jGrmWHhm88wwiU8t6VuuRM/85plQ7FUTk7M0PSex+
JuFeiBKOdQAxdGYf9PWuAc2FzvFShsiW6KHjDPKggmGPPjsGVVLnKxWhMxjN4W13
UMwn/r7ItyrWFWF6qdTpOuBRvOEnXLDMCzgXTn1r+rny3i8Xwr0oyPKmsTc8YBu5
DhbrYBaByRbOcR2zHqL5J9D7qupcUNg86kqF+N3PDc2Ck/4ZHaK4AW/Yd9S4kIT3
4PjIQAN368DnwEaAxMU+Zo2KmAFK+HXH3LNdiqk+HG8njqNbVQuSOuBagGQdj1cD
i2elkZ/8dsfVAW/EvuK1pdK25a6IerqcthZyj5/y0RlwUAuv/ZJYn5Pp9ERBl8+X
fE6ES7iI9fkxbDIEuGuFhYM6+7X5CCIxAyBdmkd8a+MtTCGlCPGSrimL+P319/wg
vcjwodf0Mmf8YFriUPxdI2ymF+O8xS//b4edPGKnBa54qYkRi9SIuAZ1FSKZhZAC
VaZgyVoMiiJ7qahFk9U8G1sDFFkLzBhBjWj9C3/myqKSmYLj4YIIzCR9WksYsziY
4IyqHOGW5TYJKg+um5RuFQLkPgBqy6ZCpZFktkmm8XkeNOjfCrr/1LtqntrofoqX
hucKaaRYic3AxbtJhDlnlZIw3qpJLz4cya9w+KVxOGwdMZypiCWT41JBjkw9FJGL
48gxKry0XxUk3CfQMQuTP+ZVJ7vQggoJk0uL8B2m801mwveAdt8OUliNZkC2C4C9
7oGQYDRI1Ac1dxlQaZqOKXs5I2Yjv8lfxNtLb/frN03ST8LME+rP6/2xdlkViIpQ
pWcnLYgRSxi8mqdm8akDTw6NewiI6yUKTGasDJtnKxZElJ9HtyvHfUWYPeGf6U0m
zK71qe0OuZEV2FGmqO39GIyqygqYbFi9w8Cf/FAGvpfZUf1Bso3nKW3JMM2oxn/x
rZGuOcgjIHHYbaqMvXFOZtQnV1uUiqMk/WBmJsomg04TjC7+t0DyEabuuBv8siaG
Ulb8FUWb7CTs6PqZIwCFGk4RtU6Yt6zITIF1xGDlkhOOJAuxKGBL7kYE+YJ5Dd3W
ZHyZsqOMCtGEaB0DCTsIIHTtFYKr36GorgA3YYG5K7uDUKkWTrZ2DBebytwWlXEq
R4DFyewReS4PEkbT7I1oy54ik22QxzpskfwLSCNIjXqSrcrF7cDB68QnB9a4Gsnl
4RQNj8wKLle6TPxvNXvV7Nj3sCRKEy2Sk0YS+jcxz98vxTaDeRI7KnvB3AXU36R6
rITi1uw5bGN26J6po38h7dd+yy6uSQOEYV7pySdVZHsY3zsFQlx4gtM53ap+GZBc
AJ5eIqTJaDGaJjPwIcREnLlPsnQiE061ufqDNB5NcdTaQeqtQQFiW13p+S8tkSOI
uuUwq8unhz/TftbUy/SAUWmQuEHOY20OyX1NNwvA05wBv37IdWYOZQwFuXpgX9YB
Lu4iiOBI4/aS9sM+AkPWtr585DEJm3zXbwS5hNKrwWoXUfI1XDa8JLRbpOibWc1L
ykIX+1TTSiRIkLIKhsrcB2aWMEacAV36DKBfk9RLeQwx0B/HKjavr1Kw4/GEnaMx
YVO/in2ogEiVxUFENwquSJcrKxTKaBAgZRfq2haL48IXFPWq/yhi+CwOfTn5YrP0
z842WvC9VzMaNcfLYNn8++KjwCEpMLU9sbh4gP7kXeQA7GJkQgITgiaSVq8yemiM
kztZcXlZhdTJZMNfM3fDTlOW3V81x5azT6VdhEGWdnOsK7deSxKQNC9j2HuwFSMz
XYNnvhGQaEB/jlCPocTGQ6do3w2crgAgfBgOW5qe/VYuynHpv6plU1DtQgldo0RT
6ifxcVSoH2UH+TqDZ24XvXNZRmZbg2vEciuf0ck1etr3JF5Ac486U9mUJiVkrOYJ
wGGalJczFE5SdSBQiFZuu6kn4uWHhK4G39gpfm99kgRg+QT0VxkNXFpaRMT3pkJL
WjjCsYpHUd2lDi9ShgWnnwLp78xuY69dBHwlnxffgwB05HjKqaZwnSIyBPoDwLLC
EPl4PTaV7iFRKoR/hltTRNO9kAlw73Wq7xJx4O88zmv/iH36q7AfmcV/e21vemfB
9z8lguDmGf7Iob/ixar+jcAf7C8L9DE7SW0Ya4HfWLnk/IZkaGk64e6KO9ytGjyq
eCn5yAycWQ9dIPNkKE8Dim9KkbUceyZSIzoyutNCJfBoBZRAz1s2fzwWwPcByhTB
g+2OTorudecojS1vCs1GI6t+bvLCyTv6q6c7LG50VanVM82iFnwIUi9Rn8mB7tAf
pkZ+WGpVvOv1j2+XBx3kajkPlkh+Hh8+4DuOIkrmXcKJ3mXwxGbPtRy8DyLbVSEg
wNwVJozbRi/gf5a5FLxMMHZoTAB1YoeQM07D/n1jtGXzJcEvdG+XqFPTuu39lk0o
wJvfi0fm77Ti7GcQy0eeAEd6DxSS7qCMXvugbKjLU0+2VaoH/NNfOzlLdbhDMWjp
A61poIx6EWxHo8WrctnwnpcMizA8I3c5SbQUVfdtSP6kcw2Hv6vJwY+4jKuq8jXH
LyXl64P/l3KoeUS0SrP4YtdfUYGwtLE/JN0ld2pDCGQBXQaueUqzoN9EwcVFsnen
kjnnimjlb7au+nREnT2A8gbuP6XARhK5o7O3x2v7U9/Ktds0HeAJEkHjrlxjU1bY
xa72wJqN6HpQDYNACXPWMKjr3p0O4DDqYUUutdAXhbA5UZauwfjv7lg/cFo5Qx3f
NLjYu7erxMfuh0JZmJdS9xm7xB/5f9IttguJuNGlA7VMFHk4uDWqEDaZY0rQGfnQ
uWWPxGlIuzIz3C7rlpoo9TyXYiz66l7LWXcPNtRAXIwflHnar1vZFInfYKajM0tJ
bPLeKNvF/Ugx3ayNPoI1XB0++a7Z6jkUGOQCK3oIsQ7VXrgDfZRJF+m/G9HWvtjA
lNmfp7z6pG6cN1n+Pdt3CKesm5lu2JnzuJpMhM07lU6TeNyd51tOdV3lREYojDlb
HEvdAl/29MqVCJ4bb4GqEAtVxHOD2+n09aDB/ABcs+aGy7BWw352PMg7vxFfeUoj
9iehIjsS4ikHZeWgXnzu3WO/2HFp3OUX5uIAfKwkogbCMqO2yjNNWqK/jPkylaPa
1uIJzYpF8t8idfzLsEIMS0d69IPxpUGEzXrv7sXXnIU/gMp65oJsM6GtH2nE/luj
o81iAQH4DecjWdJktuBDObJoLip4oKiFFrpUDt82NB3otR+8SLZuo2A3r/KHQTTv
Ped6yj65lHrPjEChuqMP0HvgmrnHWA0Te75H2JKiIFlfcq4wtBWbBYeEi2Uq/Uwr
66lSseAVmktIwxp+lOHIDqZ9vxjEAPguubOErZAWYKImi65smRxLC5hjOR5jxxil
he9g7XVuFd+uYjP1/zwc1iXvE7d+Fw3Pm+AgdozKm+9c99HkKw4wbGBriHGveuK2
yZ+4jxbMmFNxuDxrFTuzcWXKPefIIyBK6V+Ad6UL5bMtco6S+gjvDzk1fHXeoEPx
ZviuNrFRe9ZMbgA3W79L2HgrpFoiG6Zg7uCQGC6yt1v+k+KauuPJ9HghK+VARex5
DxQs1G/BoAiV2JaBLRt0GLyW7AjI634+8gaWxJSxaThDeriqNgcve3T5jKFdw719
aF8a5owl/TAV29DBjqgAFV5E6QszryY1LKpZ649bO0E1JFj/VC5ZpMYT3n3HvIEa
l3V8BPV7XazTDjm/s//q9GQBJFng2asVy0hrrWxBmJkiXBFiDSGLAEkMhwFNS7xD
KeOUYELTdZg2zN64gcCMquUf6rQN+lzH/ujja3oOdB5O6e/OfpfG7CqZXPOwFaK9
Sr696C+LNZiV/blELS/j4oQuN/Qt6OwVFzPwmnKP9X/soOLiS/rIyfm7rcennuVv
QbEFefuo3pxlsGX00g8ben1WplRSB36Kh9IE9fZijbyfN15U/luf2pk4Exo9cm3j
eUODFaIh9gaXarfUm7XV2l0d0Sh8tGDd07B1qIzqckueDpMG8W5WI8fvDuhncJgK
hnIHzYSFtHkGUf2N3OB4Uk5mKv3GsJJAEOa6Dc0EaPyaSxt1s5KZZhpIlXba2PBP
6tWjqyvK+5HUSPiwuJyG6kjgLuuhX4jbHnFKoUkL7RMfYopKx0WLw6OJkYTaNI0c
p+Tci5SXVT/DVmWTvAxWk/LTOnBhkWU9oI0XDiAMAv7JzQ11W2rDnXBYafWiiMqT
9GQuVOCO+JEo/wmIN+9CdkLxbIrCMl9u8OP50fLguasDeoQ2kHK8U33Jkuqunvgo
WBkIqFfU3NrUzlZ9cA+ZM62mzZKo3zZ/uNI74Dt+tqH+Z+ARw1q33h2Lniw0x4rj
6AOOZbIRzasm8G0PeQc7rgM/hYogPSpf7O/mPnwZ14IpsOQ/95AST8DmkUrWRERS
MsAQ1Fqt20o0BtqlZV1fN8KEI+PFVqD1BEKYUjDFaGmZqPbBNVrr6v0H5AURtz++
EW80v/MytUE8oGlGwgGs15UNvszoj+blu3szxLltBp9FkzQZ6clQSHMiyVAxd4Uh
l261CvKMeyroERzQNZCbNk7p0zS14J6e+LueG3r+2pPRpDBqot1L+ZSW2js6uWSs
Ns35iZdms/vd+zc46oOlPr/iO0gIWRW6Suvi6EKzQg/LzZlqQmeQGlyZegoAabsi
LwDUw1We96R842brU+U/1nSIWjmCklnnUgoEkqv9MP1aTlLIxYJZb/q9X46/Jyou
rt5IjshZeRj7VJ0pijaMDageWJ39qAYJSAxx7ErCrPu1EGVabfFyahqE5YMK6Vyk
cR8Stxh89qPSpMeWZvoen7tX87jxKGkPSrYw7LPRl+pZP+1UjpJ9/3r7gOItjaFp
5wrNTqukxbqdFD24+Bcp+OlMEjz9m2KiYww7Y/7nZPcGhWJrsuDiRBwSfiIsXWB6
aOPMuj9BIP/3SKVf1V4NzgrUaYZNw8vd/dzDEt22krSgC41Vwasf82Ja8/6zvnnz
qdJlOPx/BL/CHfSAMh4K3S7nDtqrmvFqMvuL/RC9ocmr7a0oB0mLeH9kvE4cYmZ+
O2P+xeYs7ViUEMUd4N6TfDdWOhSM0ymHqBDk2IHOrdgSY+dT1WPcxlXHQsgK0DHd
6Ffi1HbtISRHQYduwrA/mR9L70/I1IA10+kYmW8JFm3+Eo+eCjjh5QBkSFNUhnNS
TBX3P6Fs7FWdnQlPv80/odxCE/TpwuEqqXLFUX1/iVNEFxBTyT/BZSdKSosm1TZv
tdAjUDxGnrEWnaj9XkI+FtCPzo+H4VzvNF+9h7OvMHdKALB7A8TyXzFIf72vdNcd
rLpaQezIW45gAMTL7AL3LW9OUJSi9VjbiGYNQC7ZXSjf34qXR1y4IxiP9nwq3JkI
gmK2uqMwtDmJAtbNV0iTXgnSionPCfP2IdZlqaDlEhcbZhai91L6fg7RqEFlCWLv
GjN1vvV5SaLaz35ukLt3h7pMQzXaFnP27IJkfuPVZAVdLeO5awcgDdVGqE5lOQNI
9L5jwTyht9jDwtejN6F717kmC193P5RBsHjE/uQPCR5rw8PqNLoHqUukWMRug2f8
Oi2ASpDkr/pWRndwfvNU7MsyCOdHiPzZxSDjpzidB28MWkkH9xCE6Ak0lLs37bUp
2j7mPPrWtvtREaOJ3ikvOVLtxyBltfGkcruvNA55vzpv502wqTRedGzIFnUlou7H
V+V+eTElLOT4CI7xSDFyZGSvLVPXbrIR3or3ZVrINinTFuCkaPX+UitUij43mhXM
AcELMDe2MLQlfKI7I0nRdBIW92JgxtYf+1RyqQHgG6ohbSdV4O8Z9/OTyQfitnW5
9L0o/0id5+YoBk214APViTEwownsnoFzHSph2QX1SX7Eg4dIwjHm5lb9fr23t+WW
cuTWFP01QIG/lrrxL6ZGEy3MG3of8e/Vx86uTnQm5Uv8Ypx0kwGLIHmK8RL4271T
eSX5GNrjkXUI9PqixmCU6yNXFavSDcQWNabUiu2KFohfsKNox3ytjwwXFpCk2W01
mOYTw06GYzd5i/e77gbzm5Hl9O60HQE3JxckSrrKChOAvGH4h5D2esM5LfbW08fx
/pDqxknSwI7W98vNdFwdfaC3QL55lIF+pv1mfaboId0CoqTQmXh3asZWHWeVmwP1
254/wg0hOOcVtNeTabBivzXKf22pY+8i75NbyM5zLxc4oAIcfBiAWcTOK3rSL48w
QeMEeSIOFpUe1pjlhZoeuptAQAWi1W3pJEzEXH+fw24HmdDyuC4gNNcsKYaZItyM
rx5/+L02bQmNZx3oCKfYWJX6jiNvOQrbig2C0jmwXwawcyCfAakANVvJD1wSHY6a
UjgFyDqlt76RGeKgHLl7wp7M+JpFUsiB2886pEPGTd3lw66Jdpj+xF4duz1HCh1s
Sncrcza4/xV+O9yzT9h4E5Tei1vAVE6lb1Jyp5nF821ZuNic0Oquiz+P4W2KeL1X
Z6FkL3OWi+DnjQoMvfhTl2m+qLUpT6FC9/SqOVGdAQuslD1S5/hhHmDF/JOlz/Zy
d3Xi4Dh8jnS7y1SlgmbdD0lBipS4pLweQkXqAl4Prk4QZuM30gldyG4+FOagvS/P
G6lLp2ajByc3NQSPKM1ZJqzgk7ZCyPGpWshe6Ijw1Nx+nEmHgqHODu64+tQpvpPE
5dAmUI8h2llB70Z4O/Sv4Z3xo7CiugLiOb2khGn4FxKFTxuYcyttn0fuCbf/mA4e
7YXpUSS8GTsKedlOcu+HpGfm972UWiO7HzsWzMQVJCpSNqpiMp9uuy4/sckOd4Bz
wSgYOTlun5bPBVxh0fhOMIKJuJLAprJZtoeORIa8Wlwa0TG78v4YgayPYa1+q4la
mGgzkQPwRLtm5MuXEZy5RH9hXl4vy5o/kovzWwypMmOrR1V4NXA0FlK85K9vOANZ
wHv6yn3kc6MoqhQhV8faIbbxVsqTN3QZr3hDwwil4d5iwwGgVE9uPfAGFuDIn276
ajHw1T3amI9U6/DxzzrURMHd1wfAp72KNGahi9vefgHqeLyYZyk5qHrP0WQHHc+y
vW8VXdmtjAiYPnsqpGczVPrnM8U18ZUzYnihMJ1dZURzW9lPlt3Q8oOwg6xrf5qs
Zh2oq0f4xWCXGNbi1KuVGy2AzvRylxkfEZke7gQhikD2qnVTBP/p/Q6+kkP2Jx+e
5ClbgYcA6bHwb6/eEBy1TOuqOMvY9XRA4qKoROEs1mmMYzoGp1AGx6DCj1SJnQig
zTW6wBtoNkUGIfTs+5On3PbAdf4MQHT1aFaxqBgForYlnT84D+TJWCwdDm2Py68N
tDPNV6mP+rpwmiuhqTTFXpm9P15PC4n6t5XdfKWzsX5Ic3qEYQh4ua+C56n3/6HM
bKmq7x1T5HmxRra156Vkl040ZkyiDd9iUD6SZkEfW6T7LXnTei7S/pd2IUaA8rbM
7gCK+EsrwrlFSSjD9z5Fjcuv3EmVUrQtUjGyEVAX1Vr9fbLJPz03ts4vJ4/TXAnj
mEQXlhcIyRVlw+WZmtB8B7hinurLN/ni5OAb1qXVbATdwGuZ5zih3mMxEcEP0e3y
hQAsd2+2IkCKKFHcEL+6tCBNhbgSYhpJ8sHVJfz/BCfWOQtEoK9UbA2haWfEF4Rk
mmJygYbt9v3ab+P2fqIS/SSNAlNU1V9/gsXcwYmJaN0SUIOWx7ImFTz19KvGWiLf
x2hjIIJUZ/cBW8mSrYELriEVg98nWbQzxbzZJEBCZh6wmhlV2H/R6StVhEH6JzAj
En7D8naUSG30PiXRUSCv3aG+NnrX5Gp8+RicdteKGsU87PG748HkGdSYtGjOP0xq
ZCSzmOJKchhiW95TXJ58zo98vtIUp7T7HMPwp5m6r/S4Dzdq11IEsXf1ywg9a6Z0
z2rmug7lURqtrhtyS4AgKENA7kofMBBugUIVYKOXuZjbonDISpyjvC01siBPKS5V
adOG50ljHitibGdtWAYM6xOwr9vuIgRAevGsBHw94VO/+Q6FZfit57RjS/3uldrR
EVMs7V8b336doxA0+Cc2W+EJ2L5pYJssuwlnV7hRuQZSrXxHJM75Gfw0aN5Mo+al
NfErC4sCaIEtwboKmgODQ7kbDFqShux8muPozHEcLxaq8jYmbIcqV0fu6Enbv5Jk
V/Izf0zFh9nlSJW7caMQS+/v1R1R8x8LoI00rAPEKvLQ3O3pryKC3IyPKXXAijbC
iyGUJOB0qyejWoWoWOgtfNxwiMPeg8iSoEevffhVMKXb8zAz3jyUx/OGxPQoNh5P
vTrOZU9RiofiX8vPQ6mJCkGGTjJCpiGIE5StLr2bN0yXOCXlS/AewfEqkkHv3R1m
eDlYwdjHES/GtUDGP0WJKbB1eo+qn1sm4R1ltqqk0JMLJ+/hTcNudmh+AAhVZHsM
2culKIWfH04FXDN3f5Y5L+TLPuyUD1Dy3AwkXKcAkefD4J4SkZHf3Xg/dzJ24td6
v7fFYq8n9gVoKFmsclWtInhNk1qwnZVqVFVQOpF7rkKLiRh036jVjOJQjfe8m093
PAcAntkHUEnKHp9yNBHvcLFiGCSsdEkcrA4lbAsDYpNAzC+h9kVbNDjnwLnASLpQ
3NXgOn8uIPFqxeso7OXRRwoReOkYcQnGka5Mgpl6KDMtI03uMdopNv4QnM2/2pEl
Wt9iPUTxNrViZ0FuvOfzYAzwSKmJi5ByTUs+v/9TxWSOjiFRobl2Q2sIY7He5OvF
z1LQiPObsrDEVNeukMawOhbYt23D3nfBrlHKlDuGbwo7aW1qQjjf9OSiCsTseV1U
477O+fzsijaulHqlq8ym/Qui+GDDZXssG2AIbrFyKNR5eCy/f2GJTbIIC5EpcR4L
CWXmFWOcN55NO8/Pztq/y2qOHo8sNpJlFhezsPs7ANMto1L11C8EpDpsZAuMrgtQ
qQ0Ku/Jx0ZHArqMk280VBECIm30qpYQAIlJrKdFm1Q5ocXSCCzP0y3Z5AbI4SyZo
AdaX5KLV2s3YgC75f4TiUYXu1rjCRjRcydkxMs5tLELJ/C+yt6qGtQsgUS63o7N3
KzAj2pJOrlk/bVZ6gs7+M1/ZwVlxPI7zjx7kHqofTtBiDC2BYFaLa3svnsvboMYU
gu0x2X88vnDCkyOY1tV+7Y/zYk7QGLRH42bO0ip9icpb07e2eLH0SnBpwWQZ83SH
ozPSz+TfBWg/8A8vxqAe9I//2MTZsAgJQbMwH/lGAwm7C9I1eWhMfxmI3z98AqI7
hCZ707PRt/1+jXC7Br7iAZDMYTWptRBG/3UFPG/6MZNJvGqWPAzBewJ+x3FwuLdo
hXLz03YFAx5gyIam7X3IDf7w5xmJav+sp/eoQ8g3kRqvM2XUaHTvRTxbJJA5YnGG
DhmOg5iPp+iiW2uXTunHjBXVWVZLhR5ntc4ZMSACxNSGGzyshqWk5KprTr/GJnOX
qZlW0bN+Ti3t8BFlliO2jFvnP8M0OOSkHPYFY8L748lWoqhEDXioVTW2jQdPJx9a
mZMbcLArI5uJfDoS0vE8gEu/fC6e32xIroeT43egH0iYgQGKjMg49O/aCzyfVA1m
XMkXDSmM0/EeS+WyFBdbk9rS8FC4AHQr8WVcd8Rnx5rpK2FDOW6HXbN+2DgSOvfz
7K+Zqx2h18v0nao+h9KrbX80leZ9oxUaxhdUqpEioOjB9XFe+ut9KJKMLMmoFI5d
h42U5I/Ghpu9o0ATqecY+wCWPurdIYntPS4C/dCkXsWVH0CBBFv887ItIay29ss1
590tHaNU8W8/yBw2939Dlk8+CCVaO4aej9kKKZJtID6F8jufZLVNyrCenbx/KmDF
JawnY73PkpTXiTZ6WHIHP0sCjRISzHRc0FhIteys/BI9jZu886fgvTHuumFetgId
nswS4p9MBlFhMbam5FOYu/1SkFq3p3tudmYUpiqj5B4hUYG97QobBldedmkSiYI8
kPCcdsDS7QdzzsG4Oekf0JJlkVUcixlr0bI6KwWxEhGFVGIsasEug/h6iKtbk3jr
AA66NE/6+5aHVq9IyMOT9YaE+zjkFw3AIee66ky2KqUklTyx1dgZtHRfYiaSvZbe
rIwrillT5yvH9nZjWZO4EsCwG54cw8MDjO3oF0mnCQdFePxHBkAkuHuG6l0okB7p
DT27otX6L848/LwiyvZuM+F4J5+NHfhyuUc0F6+Lt9eQmu/CWoLIYTBfmZtY8Nex
vRpZU2fC5nHi+2k7gt4iU74K/2lTkRiRvoD5P0jAEkMJqKEZZQnWhCrrutS+RjhN
gVhRM0zV3NT0CCSzGKoH8u1VQyaw9dNeFgeIxih3AK9hWx6vpiYrceYmpG79XrZo
7zy5IB6diacR4pwUzmSN6REJbCcMs155GfflLKq95tGBNIUSg4nUKI8VHwgNTX+j
urrsZPzz4PQ7I5X6N8N89TlnwCmV5++tsq3r79L/h7RHj08Ic7n05RjAJvXPJ42R
iYkzQdtNXxKzCrtCWO8UKtdoET9enrQjfxvrN9njJx87pp7ZpS55ZV1nKhGpEJ2F
f5y3g7JFMzfYpdNEDYqX1lntuDT3/swLbslXZa7P38zYyohMW4h3UTAE1yRB/9vM
GMakB0k30WqJMniE6X7Dv/neJlRLdhnP128IzxwhnpXEUZGwGPBzqjBbzClB+8eh
9IIlP/tc/sXEgNtzWrab5ceRbejOkDvCDUjo6wm4OS9YrxlPfspOnx9LHsVCQX3z
CS45BRRBMLSmfKEP9UidrcDK8XZao4utU6FenG1CS2ClkaqtYxs/CVzNnqmd8WlU
bmXdyFGxs475KeEbE8CY/+uYYWzwKhIHBDQwTO/zCYpheIgUnmv7m3i2StmTdSqi
Tf2zJpGM8vbMEVCGDj1lDV4vcDr3cOUWKurqIVM8CMYoisTS5lK4yZJ8FjQph0JU
A/ZSb7sH2hJ5lzl1A08m1gRqryYYYoeZXqHgkzNrfLXHkZ5V1G5sGHiVvaFoHVbH
BLrlZZByR3Qjh3rXWr6mch6xJ1D9gFN97j6OH8NkDSprSjFalCmH+GDQyv9mmzs6
OhjTyIka03yABUGTGRMJlHR9Pf/9LRZiSJWq9OzJtGP+DbkHFHpzH2fJ4jgYM4Tm
hjj1S2a9GgxtAz2nT/bqV0aP1HS40yyBaHxjE/qyZSgnw1oVitCBE3FU9D4eYvcY
0UCB6j94b+uqfzTvoGVoxZGlOaJ/Grsnl9Myio+YX65QdTJaFCHZROAEVojduMO2
3JaQvxczj3IZj5X8DqwDjygS8me+E81aIMb7H05qJN6263KZ6QnxR22+8sMAj24Q
Q9QK5CbmMCyM+rDQ8MzpeBbrBVLUXe/wE1zHv9NKzo1BHzOMXZs2hzQMieOS6Nce
vyc6dtY2A+y8oMZH23PLmdszTZYKta+UJhHYFOVtpCvqP2HXmgWT07YtABBob5oC
raIxckPwOuGSWoQhXqc45vrxieFICckiYURRPTkX0v85lsoC7WUGUcfODvfTTwMO
GuzFqLeIa8TibJp6WCLGf0bwVh6bCa2j7XiTWIOKOlRTKj+mI5MucElMadbr31UM
s1cEb2POYnySp+SpefK36hcLvSj7eI583+pgwHJ8DAjhK7fHIXW6Aj19gCyunH3C
TWO7O1ophNriA4/zxNgLGfNy064udRqJHfDCysxP+/f/CSPgs2LeC9hBiLilvYzF
PjDopcyjXLN40RJvE5sSaubDpqGsNgII5c89/pa7vDHchCtuNBc1zJ2IUtGhW6ky
GCf3nDZJNndNc1HlXFiuBJ8qZPTylOl2wxXEqwMKq/qN3NtKWEACIeKSRteiRshg
oElXMADNuqAKk1VtAAfcroYiwoT3qWif61rL7ovxu5zhzQ9e2vSvou2ovVgblv12
UN1fYMAacgtMCbMC1DqUeM89Rat3OBW75uIew8IfS731w4G40KQQQ2my0jci9ym/
a7PNqdX+LYTMNoyv5HkSXJzQLbSkzmqTV9cD28iovzzhTfFB9ih1y/GPvPQae9DM
q/xK1mmHY2FQCzia7LwJ2lQBVuRaRQpeAY5lEzSJV198wN1cK7NtFDKkXCddbVmE
CfI4tsOTLgQkZWbyXe/WzD+uHG963Sgo6emMX9Lkij/3nZ3B55ubmCpaKuz6N4w1
lpayg0i2+lU+rFoZJ9Cn7tjqBmqZiC3vS594oTTpz8WkK5/qkYTIh7SoL5XwFyr5
0ZHPc7R1ngrFm6rSjPz8BcyoFvDxYCS4i4NjnaUA1JOLVbp6o3WP4jEv3SF1T945
++Yqf14ofp+8WTznoA+NpwKiq6wJRSCvvUWXf8KWQnKW/SPtFoMdbrEUKHWFVf04
EKOB+WWcE8Kb6RJROrvjRiFBphWWj6ki/ct+IJnfUDpHBVQTUD9Dcayukf6PpC9Q
cBaWu9b9+EW7cwiJWlu079rM6R+/oFhDtIhbgf9sHgPqlvtTOLIDrIHWpyTonGCC
Pzw5B6jUAA1KX791QI0lth/LYCydDyYVU4zvC/ffTTDa+nLnFPH8nH//NWglGDAG
JM0gzGYcvWJ7ZO7GyDeFP7fal/vtQB0NtiItHOzcIeEUny7xD8KWOoCGMGNy6R1C
kZZIg1DYXz6Akcm0WQKr6HhC6MlcVIe/RKVBdWMI//mX5uixPi9mjEmK+AfmPPsm
Q/q5Ma0m/wSRGT7i72ijrw53R3EnYB2Nq2rJWIcFQfptycdur9tCHqPnbB9B+Ehe
o5dPniz+w2i1eYBn1zqXlILTzETMNN2BQp0WaFIlBrDaAiFrVJaIGMnmkpXsKJ2c
l1IG2ZLVwzIIIHedUv72Hqn1hsVpvH3XeBNnCCF+x+yTQQLQpCJQr32VVRXpdHe5
`pragma protect end_protected

`endif

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
aqWVHvN9u3t6p7WUAi2fsDBl40qBjMWumHqWHWd2ZDV58PSvG5y+tEiX/lnmqZfK
birQPyd+RHpaTAlwseetQhvWnKDlbBahWQljzKBH5mC4rUkracOl1z1ufW+5roob
bBw6saVwjBZptIwfJBc5JsI9TQ310tTeiPNM40pena0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 67812     )
b4ciAZPsQoX+RlrnapkKNrDI0W85hQB7/zRTmZ+sGT9h9S9Kz1NICI5UXTJzPtUB
G21YLDyD0uNNjeUGCiSk9DeL2ZDq3Knc2JsGy3dAnI9bHPghh9clAIsog7kegGwe
`pragma protect end_protected
