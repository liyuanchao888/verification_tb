
`ifndef GUARD_SVT_AHB_SYSTEM_MONITOR_CALLBACK_SV
`define GUARD_SVT_AHB_SYSTEM_MONITOR_CALLBACK_SV
/**
  * AHB System monitor callback class contains the callback methods called by the 
  * AHB system monitor component.
  */
`ifdef SVT_VMM_TECHNOLOGY
class svt_ahb_system_monitor_callback extends svt_xactor_callbacks;
`else
class svt_ahb_system_monitor_callback extends svt_callback;  
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_ahb_system_monitor_callback");
`endif

//vcs_vip_protect
`protected
]N2W4UN)C7E4.5UHg2c,6DG_Q28.5#bZ3M+=1TZ6[+R(CAR>OKH84(78#BA31F\R
TL7KG1=J[(-4EZVW3+0S,N.JU7_)O;:bR9:9MM;&1;IeQ<f=8:EW<_&USFOZ=9?@
cQ93IbV0W8V6G,[7R<M9^@GD^TSe^>^NGZE0\/@2X5fbN-g5LA327d?TM]MJ2E&?
O=SKMR89RI:37L@B2JKdA@Q:UD@1;DQS<R(-]H:1ME=eC&39SYA1E3FRX?,63?&f
c&H.f/JB,Q7H:Yf<R?/)Q.E]-_:;#gc2\5?<3@D&/R<(S.;f,fWa+LdeM[\fG0FL
SALV+#I]@8)>YC<a<e;(CX^<O7Y7IHccc3[D1QY@RCJE6,VXGSWFa+:K.0_Z6fB?
QG+MGF.9<FCZ.=RDG)[+MfPgUbADaA[8A9X35<=5-.\EF238f;XdN#d,VfX:,G6/
c>833Pc^U7M\Z0=UK;UfK43@XE^UI-J:CY391/=UBUYDgX;,96:ZLdJC[HZHeS#D
W\P,ML/ERB,/Uec)T(Ub#;YE=+L:WM4+C(#&(+,fM.D,8V?W\1G;eTVZ,aGNLW=F
+;4K:[C9cSC;J@7BS>e8ZJ+W^)IQCgH0(&cV=&1GU7<.;;^S#HCb0WcD#68SNVSS
=6@RR5[&#g(Hf@K5YP6FJUdgb7&X5f>S>M30;44O6?&^,5:3@I8:CbDfDX/Q6f/]
ICZ?9B5I]U8,:gG4c/1I^GZ.Gef),B@Z&<D.?g#eE(CZF2F(#,QX5BYd^J2E9JFS
HHf&-8\IcDE/4J)&[)X9a@7HRD&L)#5TFLbQM1dO4-e53>,GX5ZZ8fY[BH=301e^
PLI1VaU+2P9[7,T\CDWLf.ZH-+GJc6ZKM6SPG,c.N=CQF)=DFEgI2D]d0K/OP3E>
;K278/=\D&/]Ye><6c247R+8b]feJ2BA9U2SIfJ_V5bc3/L[Cd5M@b84TK>3@X&>
^7YWQ:[6[^M.#O[&PYbYGL_\?+D]3^MALG29_2@&.])08-#a)[@eIA-=f1,.ObIL
_U\J&[-dd@e/./I];M^:FGC33N^VOVG>A?JTg/C3HUfe_FaHU_e/6D32BA.UDe+:
Q;ZZ83QUcUcf+8-<#(^gR0^R?Y.a-@TS<>AC9JLG]1-1F;/=Q1)A^K:<E/,BHe+/
UE_@N_P&02ZBPYL1.^OW7e4ZA_MD\]]8,)Meb(--]\]QJG5RV47WEd_C4:7S-A@P
&F:76U4gC9S+5PYN?/FU1X<6DYX;;/P;;)PA==3VP_RC\T-K,fNa=MG.&DIeP)[)
\E?^LH-ScSe24bd&3[L4Z7CU5T]>O;\S^NQI(T84G:gXLOD507L_TRcb<,77TJ?R
(KD0-:DQ3A./F[&Qe@Z[>V1G9G_S[1W#@c=.X\OcKJ0+/?cSODK/9QDbT]L@WQ\0
^Sf@7cAT/L,.A\CHZ@:g2,:?_cIS2/0Q:fI;Cf<Fe)(0:O2/I=2QT_8d6EG73;(J
MGf+(_@@[CEaNCC(Sg?NAMc6g4)]Hg:<=eQ-8^#U2^Ha4/G+0V4PCV#8KdB_>7bB
B:()eX,.UTWda/R#-G1V^43/N-,0Qa]8g2U00E^S]O,^=5G5D]UbL\+VISMc>;-G
6\A4_BIGYM0F[Xb5U.\(]fMd2EHgSR=I^G=/\H_SX6+LgZ:AS50/(:SIREXG.)CD
IC9AcN5dER>cW0CV1\Z_Y,>Mc.D0YG_IbcI(Xfc,e0=ZJAW_R&-72Z[a30TG/C1C
O#TX^UeE>M9fFbP/M69Q2CAI+G/NZV8&2W?ZP,\^_:H^Lf6Xd5[+J](a5]DQ@-S5
D.:W&PL1>IFMNDB]3D>3(<8YMV(-,a4O,94cP1HK=Z(F;NIAH4-C1F#/GDO=UK.W
Y7YY1gbW.6B&<,BAQYTM8aOg0^50Qg<RbVbKW]K.H1dS^]BPJCD+SY+_cSSKT/cO
V<74RD^(&WEIbZ[0(529\>(20RS>KbYI=]]WDaG1UM?Y=,L+=F<(<4IP5JW1ReA-
EYYN3VP],ULX+>)gAP:V/:GUHdLNbUXM_U\df9Vf>P/ccINAFd(6OB7JA>H1[UU[
)Y^W\D_OB_PB#;8X/Z(8M=YWCbJS8WRPX6?;6A6SL@RIZ53/A=[PKJ])E]HWBa:3
4<dMFL>9<C?LCKg/I^@.]92VLS6\^[-^B.4EfAEG_7I]BZa]RgfF5AQ#QHf,WS^B
/e.ZX4;2^EOBG]EVT.9GJC92^g&?LHCNaUd>0b1fcV<_<^b;8_>0XWE[0JfZ9^Qe
9b)@UI>EMVc&)-3+aHSbEd,=#WC6/I^FUGRLS6P3T;bFXDf(aeHC\J@XC35XdGC-
1:A\a(V1Ed/HT6N5HgRFM-IC8c\+/U1CH6.X)]A-_6+/_BC)#[F69VcO)ISW:Sg#
W5#25@(T-(>OV_LdG^?,#ZF5@X\JH4N-7LE?8<MS1VU(-M32NS58=S3UL)2aH9#G
D=Q7L>gEQRUO+$
`endprotected

endclass

`protected
+&Y5Db]9aLV^DI.QKW1Y#02\_[a^K=[-KL6FJWS:K@\<(eM+R]_=0)-MHK]U.<d_
,<3GA)G=a?dO6/3-SNC0H>8[9I.90aFB7)D4./4gPf:(ETDF[C2+)U:_H8?[g^7.
(#>(@=LPe/>YB[U5:cR@d\fI6RKH0?&#30YWWcS(V@8Q\L>42@g,1UOTLgR1cgbL
=f(.bgU^dC#^-:<P\L3-5Q?\Bg/+Z;NY?@C5-OTK?QLXAff8aHW0RMRe##T9gP6Y
@5F(WC_8G[L;S/Oba6/DMB(:XSf+ZU)_1;7IMDN2@JM\JX4_Z1UHU1H)=+b)R>[(
[e1##C[VWeBC4T>#->VAF8FOSIa9L-#8d.EfCPXP:WcfS++XLBY<#\81G8X]VY=B
gM[_fG&bCX3C*$
`endprotected


`endif // GUARD_SVT_AHB_SYSTEM_MONITOR_CALLBACK_SV
