
`ifndef GUARD_SVT_AMBA_GP_UTILS_SV
`define GUARD_SVT_AMBA_GP_UTILS_SV

 // =============================================================================
/**
 * Utility class with a collection of routines to assist with Generic Protocol
 * transaction conversions.
 */
class svt_axi_gp_utils;

  `SVT_XVM(report_object) reporter;

  svt_axi_port_configuration cfg;

  extern function new (`SVT_XVM(report_object) reporter, svt_axi_port_configuration cfg);

  extern function void expand_gp_streams(bit response_data_valid,
                                         uvm_tlm_generic_payload gp_req,
                                         output uvm_tlm_generic_payload gp_streams[$]);

  extern function void gp_to_axi_master_xacts(bit response_data_valid,
                                              uvm_tlm_generic_payload causal_gp_item,
                                              int sub_tlm_xact_counter,
                                              uvm_tlm_generic_payload tlm_gp_item,
                                              svt_amba_pv_extension pv_ext,
                                              ref bit[`SVT_AXI_MAX_ID_WIDTH-1:0] gp_xact_id,
                                              output `SVT_AXI_MASTER_TRANSACTION_TYPE master_xacts[$]);
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
HF5DeSXOowZ0I0Uzg6mvekRUyZ27b3ogIYZbLuLgWpwN5sIuovRf/IWgh/QV+Mnk
Ph+VL/ovFSmT5hNFuDLgHSqRZYdt+bnRQEA6wxwChR3oKAz0NRLc2CLVlceZsWNl
c1IV9ZXNgJJdNuAQu6tG6J2/0Xt+UFe4gAKEe15TnFC6ady+GynXzA==
//pragma protect end_key_block
//pragma protect digest_block
Uq8erDPdrdWA0a5DakA81ivYOhA=
//pragma protect end_digest_block
//pragma protect data_block
+cWoTgCoAltkLzmxSaFBPAdpw1s4nxmpYRQ4rSmbfEXL6g2RaxWxhPW/wI///P2I
qIBLQJyqYL4lbHIEiMdz69AkOJBHtPEUDG+VQ5U6fyHCLnkmXYtyhnQ0WSkg4LFn
xJRKLG21oPbHeLChVvSaysUIYhRK9MrVhOkI/c//rvg6h2S6Kh/BxOa6A0dAgYts
oJujt9ylyTsSc1kHYC05vBG75ihwzCdMh3eNrir3eq0EzHRuHqLX9ocseUU13ODM
OD7FMDTqTjA9FShIo71k7BjNx0XGdYTl9245XvmQjCRSVyOmiTx9JnLhQNOjiGyP
gbU3oa6m1TypYU7i0lZkwnujW1WzIvZcT54MadN+Lpk445UMu8Q2vtXSiBY+yFFP
rOoEaGv1A0YDz2RxB0o27CIwqAYDD0CyxELV1ZfoQJQKLVIySY96t033UF5UOLmA
zCrLNbyGcE8tVQGx44VMYb8MqdePsNhpfn6/e+oLM6aw4V02yF4+m+7kUTUVJ9k4
S1nSagjXFKMTvqKKAvQ1GwN1qwBcskElNR//cw5S3nUIk1HGegm1235g+r5P5qjT
Oq//c8AYS4axFosxcc41h1Xf+Nq+PVvv+mzWIWd75hjGe8aXUYeCdJNaf4MIrjNj
+Pk0/KaRk++cdt9fFxS5NTrkTZ13oVNOI9ZDm8GBLAI=
//pragma protect end_data_block
//pragma protect digest_block
gl6kS73Ky+6MErC90X2CnC3KZu4=
//pragma protect end_digest_block
//pragma protect end_protected

//--------------------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
VOo+DFOrvXKORPZawVOhz3C4hMxbBD5ME2qcXE5jExibFAQ4rSVHVGdnl+se897Z
M/4OF202TeSXJwad6bSTv4PDcnDDq9Dbph/gUaI6wdX2TJuJxvwsIJJLD2CMknym
XNl5PI8/W4QbdJibXeiuRshpLQDHL+7Pjehp/fDDlah6+r6TK7m1Bg==
//pragma protect end_key_block
//pragma protect digest_block
iAXrJgUD7eMVySDtACc9dTonP8A=
//pragma protect end_digest_block
//pragma protect data_block
UgtuhcZtzdE5gJJAVzMn4Vft/rzWmBVJJv1IaSQUTmaXG15fDOgkT3Ahf6n9lU5B
oKZPnLcseOexU4EODrL0uiJDM/6q7MG9nPMtRfaYX5SpFsvMF2dTBpcMYTA26G4v
BvYN7dz0cmQO9zVGSyCMUnW1KtUrqktunxlaJaJyXLe7Qj1+2/kIwO90tusk8Hmm
WwgOGVweukDtPVGK2swaxxv76jTgfTaC5Kg1eT4gQBagmgJk9VyjRtq76W2MS4hu
HCPhK++Dkb0heJxzyyaZ1qkpGKC0EMRvHD4cd39ITxvXChaNmIpf7jlF4ByW4pem
GnjYx4nxvPnIrJLpeQcnq8AxvjyWWb2e/3LK/QM9wV5L6slDEmTE//g6egsHFwVD
zJHCQNKhSv+8l/usre7cGc+7mkxueWsW9x2unl6TK1EZtDC7hCIuKnP9+pJTmK+9
Wg2/aTJ5xweOiyGWAgmxo36V9lYReO/MvupvLb5R5DZhPAo9976pV2zQA1dK7Few
ynnlXe0WtkfzZ6i0t0XUpx7Knm9QPGchWrilJA8Tfvuu0G18ZS/Q8VDXIoarozuO
EYLaBEo/Q9UgBhiZHv4l/Bc/wevSeAp58sqnMCEtG7U9ybJVZx+pNiFrlfOyZ0V8
SAo8gK1mBWG6hf/ajnj43zYi4PVw0nZN/HbCIr8iaOd3Un+YBp0wHlhRnedUKdji
V1RiqdhP+vsYgLRKhjpSzKDbitMqQ0kGG069GoDqXYmJwqalZgSXTMR+zgd7cTXT
Yg8LLgEfa89HikI9j/giRMc9+M+Dc8iY4nBMq5SdVIvzAE9X7G64Fyg6+WJ63qBk
DcsQWpEsUYufZ87uXf0T91Rm1whAPGwV3isuD28Oxdtr+HjpUaoAHpqLiP5hDApr
MEr2zqKV+zqopuZr/LP8AW5ZqrFAHq6oxlImyhxqU2/zAK5Z2I1wBhzTCQJ3Mc0i
1heVoZsOdDwnk0kNp+UPWK/1Zs4ZX8nVRiyU/5bDEpAQvhB0Z6dI97lE8GQT1ihE
eBICqtQ1WQvzyHU45K+cF/3B4N1Aw2WQ2Xow3YiGCrea8441BMyRJG33mjRIiAdO
0Iy5fR10eKQXjjtI2jJJ5KJ8Qgu69dRToXqw+FxVo7WfpWXSlNutZE3I55XyFDPG
/eD6IEf9Pf3Z6QNL7g0EUrsDXK0AacAOfdEitoR0ESVzThu2OpvXD3AtMJcCq47Q
TDE1+Y2/riXncJjDKCGr9Pr95qICUPJYYt//dY9YTsW7eXPgOu3JXGdkEV80SMpl
gjuh8IlaXBVad9CVBGtHHClQb/Hkyq2vu7yzIN49uK8mN3k7LJWvN+3bJHFb/QCG
FBhTyLevFPFrvdPzDD0FzaoqgleKHMIFDG3gNmCGamfEcSWmdcOfB10qBTjsFfvR
ZeO7u+5li7QCPW7vmJlxkITs5iCzJulY/51qKLlNSjbva/4aZrNeOmWxQ/RSVaEm
arrkuzFjwhwcaeCo52g/70eIwpnYJkfp54muMWV8xqF+5ZXQ8cNjaa2lqvFnTvkf
F+wURE7KjkHJAzVDWWMnAwxLLqkYeC5wVP4dlAnEImqhEY+9+qivMcjKcORsvp4s
DeITavlueqBb4GqI5kX7ylrjCQuTBisUd1cDzhzP7GFG5WwfH8DFB5Mukqs4s49G
R+8bZw0/8egeOKiv/A4wvS88gfSHtKsrfxiErszZmzsQ5KPn1Wukh/5XKQ4VE8HI
SHTL1DVybX8vJ9U8bVNqPLMkk8nPvALs8aUlhgJXxJJzNnBvkyT1blg/jUjc97BZ
vCW0e+Fi7gxSRLatOw1+4n1tH72POOqgiB2bWslaPzZcQlCLYE6mTD1x3iV3x7X2
HmpPWd6P/jjJBSejKV2vmH7O9uXgXJk4RBXH3CmsVAS/PmlcazWocusWEQ2x1Evm
cQEWd9PfKY2k3iot86Q/1Mia7bkiNjLnlIoOO/D+LvxYnhZuSMQ6vZ4Vy8wro38W
riY9d9LThFd3VDGM6+tZxoQXzvVpRcZBbpKRIQX6kDHmAdEzWugaS0t/1j7e2hnI
gmAglUBKmSPUD/7xC3nRuTw+6NT7n09wHd4L2ZOFDRxQc1XdsHEi6fud28w3yYXT
FVxp+sZPUfohz2I7361nnhvLXEweWSli2a7WGgwO1L7iaWvDZShzQJqsq4q+EqCo
F25s5drDg83uQCFj4tivWQOcwJApERYTvJHseo0sVnSNCP6NGJ7SY9w2DBOHB+w1
C/vKiPv+bpls0GNZLwoZaR0pnJf68iP9UflU5c6nhgQo8+glnpnJwOxunhWKc299
5NRB6fExbWG62InGPXflrHKNgjzl6nKVJRlvYHh77j7NGnE740nSKECYhQTkBRkm
yD1vL0e2J0gbV6+nFGO0mgqzAigbaA9Q+MIFZHCXeF+wHbJgw+Oi3PMptzlcC9LZ
lvycHGzpvFmNI8p5IXzJCF9QRXQrriiJVR7c0x8SGgz5DRpaB25RuYXvtgpinGkM
cvpK3tjVJCQvQDUjDVtNzcHC44JRn+hlUs+mRTz0tntQFKcb8mf+sqnJqdj1mNE/
7g1CKCOplMp9dQ0vn1NkMJmq+f4x13a9GQRds7t/P3ImzEfy16GibcJStJ/elda1
aI9x9DUBMKF4Cy4b+qTplhJvFMOODdim0PYYQ4HBYI8/T4leHy8zf4qhE5Vu7Mso
tUW3vMaFq8ChJfWaq9Y+PdVFF/4Wtkl4Gafh0ibuj77WLpFfqh37XywKU0emCu7A
zb7yRXUXjAifDoWhKI8sLNyytPCBWb5v/Da//uuwr4VLASvkbTmNWwui/F7ywq0E
PgeLFME70PWGKGTMXKZ86ppoVJuL18bixaT5QT6ckio2KAhP1f/V+lj+yJfE0DMe
vewdz2ZkMARdF6wSmhwEHBk2wkCBfbMBDg+CQ2HKvgof7Be9SnMQHjUxloIQ3XMz
hvZ5hBZU7N1reVULWsdQ0pYi4JVwt09LKHkRLYGWbdRrZtKecLNprRuT86zf3otH
FG235+/8u0UXQoge1zgUOjYKT/MceucwH+PwcPY2eFYV2/GpwRYzvdmTw3j38wy1
Bw/XT4NsMJffBQhklrG9BBZGJOPzltrWn3tZN/b2Ynbt0a3rYv811eNVsddj8GjT
STvA5L6L2+pijyNv2FPn5KCbOWO38cVat1Qx30YkwUyYDfHYpRnufM27DWrugVzQ
5nf/alWIZ4iA6GICOz2mZ3+13CP5Ge5ZQnjldymrF1KpW6r3ITpysDyfa/2N5c9z
46NPkEpkUUTFMOfFywLkyBXQP6UCicBRO9YmbrbVlEG86Adun0h24lLzTDZu0gO5
2Vi2K3hK+SL+lVlownYNvRdLToJ/hdoBighsJ3Q+yqxuadmM/m2lYatHyxB1Uxtl
H/PELJmxzljRWm5uPvzva+UN1ehmZ7t1YllOxG0sTYjtrMzVEHO/ncIyGDyzX4Zg
rWwJPAZcC2YnXKpU8gNKFb2/T+B7L8oR8Z3vpMLepyqwOY/+K9Kp/aQ3e3ar3o/K
wKtrgADgRM9sxiPIPT7798TTo2si8pf1HbpmhFadN/QpKSfYk9ciQHfyTv7yR5IO
ZTcRcSyyMfycwG4tyOZb5O61cIKsi0RRY5DqpBm6jk7+9uBBx8RDB4jiMi8tfVs2
H8Ot98QkOOBohcpwuCitrM6MgeyA71ACpfHZ/ZvCgito0U+NaQ/EsWRrGfw5ReSc
fz8Li7PRs9454qFiDDaQuV11mL2YiAylcC3HjlcS0AMfXYBPzz6L5/EGs+Y8CJyw
v8BffaBI4LAoqcH8jE/pb72T5ihCCUVswQnAKlP8uk/jGHZFucjSf8DNBK7znX0v
/pPNPj9d3w+a2t1Hre1HwdeqTtRk3EubxXJvFU7f/sUZvULwQ0spTRCbvPq8ZIZ/
EOsQZByRCbBYSagkNDAv+YhfugVQ0OAZaFIKhR/S3KfZ/fDGuBB3o5ZgV95G3CZM
enVO3m4MOmjclIPxNF6JrqkTCC1K4GvXSwi8WnpTgK4MFjgaDuAnqlueaAX8KXzc
dp+rJsRHezaTs8EP7P3VY92hiKYyFSOjPN/wa6ehELJezj8lLclT15rKIIeu4w0o
wrnUh19TQD10void6pVjAe4UQqUCvWE31/+YwuvCZiwZwDWBFSfXGNHOfvsLNqzE
RT6yhXooEFD98Tohyiu4+0PGom3oedgwRd0wATfENaBvtgL9pouSzdZgRCh4dhbN
U1i2mXdaVHCKTja0g+2DsnvK1QqbUEmB1rC2QcvDlkzYHGLCY9eX1OnDwLz1VA44
9KFtvWYZJcF44dKBf4e036di0B6j/VV1g1LiB8wlVlaOGIuo4nhPEiZF4EPxJeZb
wrZ4Ed1raqEYKWEJfq0iqZE/2rSbCQ2CofOVeHGQccWviaIlAUPg8xeWOnwOIBJw
jObBIlF84RkmJzfQfyqXlp27KmG8AMpP0DTY/eemvUYq8xbCZSCAUW2gmqxXOmVe
aqROaoO08oiN9wELY8KzYtlX33OGuycu5Ez1SX4LXvpoMJluXXh3MssK8vFCOWPX
VL50uv1QBqdVBmDBigTY+fo8wiZ9jKjajzpx+b6ea9Jg+iYVZujsBjCsIS8Czhaa
bTmhmRUchgltvQc0r5MzhnsUD3AhNtIuW8FLsRyfLH4c7x2GwzRA0xJj0A2Sm0Yi
0nnaqlQZhPp8MpHly8a8kNq1zxtrCwQ0LKcxktT8ZyE0nH1sKO9Cfy0o5f74VZ4A
PbVm0rUTg+vZPxDfwxT9xo1yzeot2sWaD4vursCiuhLOIT9DFVNHWGE1XawcrqeM
hFJ4/Ri5Vnak9mseHqCAvj6vZg3OjUok2w7qEB+UNhRJSzacKQoizq6b5Hwpetqv
+HoitfvIDb4vRLGWQLFpDMZioDUhl/7+0rjRIEXiV6MXY6tGgHu5sYdOIDXY1phK
X4DvIu++52I5kJ2KzUF7Z4095W/p++fYESSXCqJu05XpRDDG3GQO0xuWmT5gFzIi
Q6qxbF9/pQKYP9919VbdtyO+fVyXXhDOKiPU1GSxFWYJBw32qbaLbZFqdpdrGDr9
cVqKwzihmCyZtNSw+uVA1RY53g0Pzka4US5SiQTquxlHe1vXrL1WyE/UXAipgPVl
TyH17A7wV47ezR8POe+CkIHfV8oF6U4vZF1q1rk0zGPmIuyDWvLKvOaaBg665C/C
y8GC2VLOVA7bBBtRFaKVxOMJKAstfkSPwzNDLQ3IL/tqSjDLFxsYCp5LvjDEJKls
3KnqJdp0K4CobdDK9f84YJKVJlw7FWQgSnFstYD55m+ouijgbKO4wCpypXTTbXj/
ha6Oyi3hVg5lIOS4ePfBaC8T4JSH3U/dJgMPJQpZL3r8G1Sj21QXkpQ7jflugoXz
+744mz0wwMXpBqWWmCmY69F3H+AgWCvKlSQ4cP3SuEkCA9Oior4Q1PqfCKlvvo3e
9qCCdBCYOnd0SAoNZ2qLBw1C0S0zYs9JoUWwtCaDiuPt32lateXYEk9LqpDga5Po
a28T++Hqu444mcz35WJdCq8eUl1/m5x/2820XDTjYBsXUjyekCbvmdeDoqwKmGWi
oZfUw3ez4yvCVqAdLGDgtsWvmaLe7gDf3fByrEFvowMFbKF68Gnss12fwdjJCEem
qVj9HOcpu32LgRuOWGu3ie9ipOnj0X6hDW850JxH7TktpuWAJBsIrBqmoa/LZJrS
4RdBA80sYDFUtTfnrgk7wNCxrTjURUZa3MIzAwrRYL5ysEhcpb7tSoAsNc3yWWQi
DfLNdtnqiuZMZPKiYBPxkqefR9tsKfrZsL88jW2ZcUCoUkRKVYLa/BTklKCDcSEt
tFqrXxLPNqUSeujD5pwntzKD/zJRa4TqxHmoYKcpiTajlQ7a8NdenSWBF5YtLRGE
kKD1FycYZ6NfpjMFSfOZcGV4LDa5w8LsgCapXWltSdOsGGcTY+S4J+QAmaAs2sRv
43rzi6vNDfEd/cKFD7iafpZwCN55DXOtiI3LYVtXisOD5GcsxRqyP/svm8Cpn8+L
2ehzjG9hWutilfhz9+KXlX+7VeU+giFC3vDy+ecaV9Z5Y2mbdD1Y+xvetr4qtfu2
KZ+rnspF+SFnmVgirDPOnLP2/QqzopUW+xOreh3H+JSRaq+HMsgw3lqmwaoQzBv6
QsfDXOz5eIbscP/r9OOCcERHa48ZFNwu9i54RRcKPJcKNVXQCf3F0vEmasf2zIaF
MntC9SvePU2D07fq+fEm3JPqxiOqgPo5tBFVYAvj+5O0/72lSEmB1U/GjOSffnyd
PkId1yAOGnO2UsERD3W0n683qLD/PV2pYjSCMsIVzmd2Ih8JplHhTkYVVRWgmIHE
5+9yBPCy26gjWHUEbGElRmqZj2/57v6jWJhkvO20mn2cKwEbx5fGgd7JY/b3E2ld
zWdGCav9ktX6aPOximtVbXSOqjafuRNMWTlX7RHvvPRPEjeizrQbMoBuSUr7fZdk
0cmxunUr7eV12rW1z3TqHaAONX+WwNWV9GXWbA/MN+ux9C17+DtKGj6wEChKqoay
NLWmoV594Va8637TMD1ASP8uJat9MKAW4p5+yF/T74d70yzk0m0GAUSPhA+60f6y
2wIhfQU3GizXY27B9UUNRJKIRtRADkEuYKMRUB20Yt3nEy6sWhvJJg1xbCnuneRh
VRdfWPyfmwHlesFSHFujim+VDqsvlBk3AjazHsPhNc2JhunRXoMeuBCHT+v88MA1
Jdae1yWoMwZOcXG5NR0z3LFstHCcAk26zBb6vduq5yU74CG4i8wApSIrY8xBix/P
Izf+uAvz6+sU+S388iI7P0mKK9rSUVIfQtVjncV+viVQEnoTHYf1az2M0zcXCyvT
eOr6JmZE7GdG79dh38uPsLToG6if/ivv32VEO2mcw031l9saqcKydeOENPUBMdin
04HXC/UDZabSIzkrpv3tne0IfihtnAjF+0xg6GAAPp21ESsPwCFPRzvuOZifHNRc
zeLGsaqC/OiBNrq6n6f2GOCSxumLyYnwc6ReeG45uPW1tQY8rt87q2OkMwCFk+Vi
BpPH/RK61aj4qgziTU/aFXN8K7FQ+yE2aG988SqDkvK77q8De2FsEeUraJ31RXFw
Dy3ziVJhxOuifDftoAdvlhqQA3TPx+XG8Y16HMKG0nqoDaefiS1bb4mKFbhm9IjJ
wg5UbpPDjiE8nkGS+8ytDo3y9dwkHWEyiI3axMHrZU9Za4L3PJKn8WLQPBFrzGOJ
eXKrQ/tYGmKM1HIf3zh+AIHP6av7jzkTxJWo099mNDIpAo8RjVv4BFDXFo89nbjQ
z1Iw9kTuDQB7lbrU+MVIhrfOr9UXuh1lO05Rvr0+z1yGXugNKHF9zFuGpXlNU6an
rtDwSewvQFJFM94kO70eQGRoSZY7R9QLRYp4E4DqNrECdBWXlWszgGu2RsY5ktjv
OfYw4LpQw8NZFPHcfcQhGdFq8l68iicDfa32BRSpeYpld+eHoHLdkTdTGllwF86M
upyyaCWJs9qGN0KrPNhQfttORZUj23yCopXzWEWa57f0r4cVShcjiwxeh1uYyG6T
HXsd3h9vqNyUeH0PT5hVLNbp2RIcJZ6mqvmk+vHWXttHHpm1AvOUKlrRir+oMeWj
v5aeeB80DRHG4HclJVB92hXNNG/W/cGBvsQ0AlyBq7Fu4EecPJ94TpZdb+cyyFbO
Xq1JzQX7HUKqSdzS8afD0/oUDb8PVGeCbev/hjr1ajhpSPRoL/D15O5WarDTttob
gOpROVjuztFisper9+iyDF/kAQopXNTK7jpfmZqaa5BpP7QhGUEgnub/xKv2BohD
TkDkLBevtEtF6Qted6UUkhkNrMebSk+C9FpswzxW603uZIWOIKLBXLtaxUKN6hjC
XSiX+QKvL46TDtRi1HMLR/UOIR/yVjbGIlxFSBYZ08Mk/BU8YrWe6ujTBPdJ4H1a
gdfIQ6LzeCnxatBH8hsIF9VvGuhEXYhpLp7vjQYZ6DHQZ0A1mKqFXzba2+NY4DE7
68moI9s/ymO60RbzomvA+Lkzkoij2dCDXenWjGMTXrFm+g6CnUJDTjbAgSVZynW+
8O1OwAYayGt8jQcdaDOMxdIkjJWD6gQCW9qm79MfF7yHSqPsjGHJckluW0quJTuW
cZfTtpLRGUgXNkHk2xllzcez1hLdxzJ9BG7+QQNhiuPHz2/4r5sNUCTRFQf3t28J
E0RnxZGsuPwmgoZbmsiH2P7xFoIVhhNaIPuXS9PG6+6bNbneVJjFVbQoIoq4Fi7a
iZ8B4+oGCx63QcgWQrS1ndlGh/Qpifich4taKNKt3M3YO+1/Db0/zXgOpa/UfXge
ys9C5yP+0Gn63s2/i+TJMsQM6IpzlAGuoqEmtVUwvi8xsVNR0vHrjPZ5fFtupOWh
FTpMAWMXxNnI1C3qb+GmiAZSAl8EQq+si7GxvlTca2qVdNqE065SXNTmM5jm2oBP
yV9vLJLnmWCOsWA6/HTBDPRW+JwVQSIKTFbrTRjVZ7CFgiiABj94CvnRPk3pnO98
xVJ1QIk6eOkgZCQNx3XsuKbfPzrIJBryguQfT1U+EXveM6kLQvqDWyV5b8ec/Gu9
mAY+g4OB/zQiJxHQL1sRb+B8y8GW8n3sAIuKKMDKMpU/YXCgArqE/X6nQAlWH4go
nEqpE7Kk7EqZ1MMYSjyb3hmmkWtGogPB1wGgc4T11mdhd5JkFS9gI0PRyihey4Ew
6X6171LQhNF7zJiZ49nLqOS7dQg6eljNGDmrPngbqftiwklsO1G+js+Gk3c3lExp
8NQlsUGvUSko5n2HzvKwKT+by56XkLiP9v4Dte6Ui15jKydVTIelYjjqhJPr2FXx
Qygy7PXpxhmQ+/CslDj/xAsP6SrppBQXnODPsnTURVzoA97zzg0kGwW1Uv9D+Cd9
gcbht07yoUj9LnyBqxE22+2EMmEAMhUQi/Uw5QJX/k/kN5AFZVz8xlD+j7FdYF9t
g6UtoFIUT71BheRVtrbcz2e04sFRyI+aixnt94s/f1QWJlR0cgTSaJsaan0rQIQS
JS+2fMMAcoDyArghVWa5fd3Uxl7HI/gHvCiaxZuBBU7OBZO9GBBuqlX+xkIEM1EZ
vMisyKwS8OMosLhO8c5mOXN4EGyW6POs9SHxM13o8jvJIKxQO8aPkUjM9F6mmKzB
9ScXuUhvK1htuBNio4f5xVpOp4CeOAq6V3iZsiWxUMOqEtt1Q2Ab+merDJHPturh
gbGup9NbnwZe4LjoUbhFC2+ePzbBr/BPQ0B9GDp2ALGLcv32cqwv+WLgYxtGIyCz
X4HNWdMouq4w52bSSObIv9FKWy6nZq4KVPCCjuSD+Y+AYL6L7//j4hPquaGNmrE2
Zv5rnm6rgi7FsHhLxJXeaaspSUVBJbsSWdqJkAR5XJ3oCDf5QM2344Uh4nPr8ybz
UJqvYbEWzAz3vbv/C3mz5swI8Hsv/7yyp+JoD33agopxONHhJoU90BixZ2Um2LYQ
Uqkt30AqdFvwEJ6aghw/FpQ9XjK4u2njf3PHhft0YsPnJ+j1UPRn3UTkCOtgaPl0
PEBELBVl2o6EblXeB00cVOqz9lpY4MMjsUyiSO5SqJPy2Ibe5uleKH1VNvU0Q1dC
eR2uA3RkyKl5YCfC8x0aaM9IcCSxeTK7+g9zF48HoMrUzZ6fML3qriNuVcE/CjUg
a9GnMJnHCMW9Jr2Ywn8nwB1cXZySHbFdgrmOcmDe60Z4lyN9b3rWpjFcDcTQRiM+
IHmygXNi2qZTfC+WldjldIJdcgtykAMO8PxlzZTG35creUpR7AieU6S27H9nIXhn
7XSBent0dlXcuQlOWYu1HfRhVx5tVXl/kAA4xol1RTNPQc4bd1A+NvSwDshTwyog
nAYlcpfIZy6bZefr75+g/qayHMJ266G3YwOI0YzbEP+y2fUE/PQuhDuAbp+vl9I3
ktt0CksVplEYYvfbHcEFqeh+2jA7c9bpa2+MonPlCyz5k9zeGaZhoKdWlCfA77x6
CnlNRodsUp6XLsv4O56xtRopNETGMvosgvjtiP3XqYHF9xODfTlggyrRxhdoB+l3
ipuP3KdrD2Ia58mtTSPm6QHHMPosv7KXodcZVSnkNT6UHFZjhsKuNOC0kxA1aX2Z
zko7oA6yXdnMl2flzdt/RV86tFqzkVYIao6C4MyYuBr7ljBI2LSZOlrTsg4fCU4/
j86IRh2wMjWwwL0SvWAl5SVldpQtrx90Iquc3EtoE9WkpkLdhwxzKNBNeDqkID/+
UhRGtvn6BX0yyhrSEIrCDefjUqDd89kWL+NmHB0CHLoEy3MU6ohfZjYDPb1q7wv5
nhhMwz8AGN86TXNx7Sej2lzMNMLwY1AJEolQ4ggG2yJlkko45gmHtjJgS8mCuZX5
jmW5NDi9tiwQs1l9yL47Ml8Ccfxmnq2BS/V12DZb/EEly8uHPJUKSgjXNno9Fm02
yZysxB7FTc4kf2bSDeq85BoUOezr9nJitpJTPlblh9m9IvcZD2Q9TjF1ITfxRUoD
nlyZF7DKXF3//VGH1fJG5wuLYPE/CbMiNtgUnqdrQmFHnz56G7edRVnS6M+baXPH
xxG2gTRnWO9iBWkXike2ngajOp+yQzVusRV8fvFVnxkFfjb5k8lFYEi1MjxEzgEa
WS3nexV7BVT+ajUr9DytHuHOCyQ7O8WZiIhlE8M97VjhvhQLMpctd+mR880/F2pU
pEV51ElTobETIOUWcCaijPlvSzhqo733JAiX1+8jyVR49TV35tYaywZ+NjIbQg9X
dW9fONMgLFMlRr+1TxNkZ71VMOYRT6M3bANz6tLf7FlMr7ZfOEZLpQyxIWWX6Y/6
ZtS/QhrJDT+DMITgPywZBAY26rA2isL1PrgktITvbVXRQhA6gGVqjK/GMYwtMLg/
kGq2VRgLK2elSMEcYZu0nt0ntowjKYJNYQZ9F95eoZfg9oJEluhgaM7klwb14xYp
b5CnBsjPWEwAi9isMRZZbvs7/lIU/+0JjPpdWYGSlDfEwHd01y3+Lpoq77Xo8LWq
EJ9tgyWH+kiBTyYHXN1+AyP/XTkIo8Huu8MX2KyV9oEcFv285aBxNXWkpiz22pqi
W+H7fYEJ/KwW9JFweXpfmfzMoeb8cVd2eSheoH7C73+zNM/SzDZv0L5WmhR3V2o5
LwmZ6AnQEuASgsf5gRRH96+aCcaYT8DiDZRnq1AWXevTZxGrTlBTcjaAE5WPVdhg
YFGfT6Dv7iF1kvrIyMrvAMPg6JmzpORxAgMU2qVMB8+0lltu1+idWHyGgm5eS4xs
ZmH1z3SYia806+zftlEeoi33AFObFBrpbpuCRh3MVELff7SJFJG2uHPS5Ctbxvt7
rU4XrfvaLDyf33DZu0Wx+eV24eayLOiyGyoe/h1142umS7PE2jb/LcGoEGE7DctK
0oSYUMZdUcQzbYDHOfSJlosJ+i63QqeNw0skUqyYMGX2+ttWp0DW6AA5mQFqjSbx
OF0JY4q0Qu80DnS/8c0sdXrLLXB0KuUsb8jfeASvvArqPv1DAHnHSVzYMS+xxh0y
LVIribY6GTIDoQvqUvXDw79c+Cy0zTYHPqPZpJxl7bTzXOjBKExesmg+1enB9lAn
c3Lpv/1jrPe6mBwaORlRCNEp2klz0yOcWKPhmE4uK2w5YePgY1xuRio9UevIwegl
yXjFU3tQ8tCfzI3fztfTXDWZHRHSBE2OGe9OeJ3XzYyXCAhzyJxc6V/la/CeM+mN
/HRhbImCujXO6xckMLfUebRyA9areuCCrazBh/YS8zjktL4zOIeTbB36zRERF3ZM
be7B0Pqpjdbt7YSNIfcerlVTeiKDTOpLKc9b09fx8fK9PN5N/2H4Sb8HWtBiNtJi
iXXaHrqSa07uFQOHCRk5y2SAtkjqNWzARPkQ/tNMl7VPB3q593IiBBa6qWMlwZqv
wPInHRfa1v+iGZVtGCYBZtCd3qiWCmUREllQtLimqOMSfGyx8Xp50beld27q7gQi
eQ1RyGRWPlI4Dxnz1q7e5mRN6OuyOUdgRM3YoptynhNOKWooR5VkyX+JLps4T9+O
A+jfBAlin5UOFTWZlYrbVde8F50yCmHxWtsMzYc0u2PihdoEHzBLgA5Zm5H/y1V/
OMORkQaxyO1bLZR4KB4L+7t2L9Wsp/uQHwvFD5KRIP7Rd62aGlYpMS8Y8pe/4rVy
hULXzagDY5pe6uzK5jr7WQYg7limw8SJyVEqwI2W4KAbisjpqG5XeTxLu/kG4mGq
aidMTJGcT3Wshmh3kqnG7+xefEwMQLYynOxj6UjpC8O57i8nFXNYpWzmzfzKwDpu
vGWjMFg8FQohTqgzXdLEEXDPx4fyhsT9knW9JkRHOpqSyDmc2uvv9mXoerTvSlcO
w/Oftl42M1cc8AgpcpC7hWEBzaN6Bmw6F3SZmD0Fv4emOD6kIlHf27vdYWnSAftf
8IbqjSk0tLG/LlgVhY8BXXgpsFySDI17fUwao1Pe+la+djX73iGMK4ClHlCqzsLm
JsbwIa2uO4r6achn2aYpPeGJQmSY9d9FE6jfMWaZeFbC5SL1PoCtrZEwDqSKBHyr
EgFSjncO0HVd2eXEMf9BmMZkfl8WNFFwBM3GW8enCnV3UFbTsZ3vRkXVhPfww9Wj
jwTWThxurN8Cn45iiYDxd1RB0uj+TrlA3/NVyTcMycQdLYbhnSuObuluFEyqdYLn
PjxLuOZVqYc5hAdZAeL93cHKug+0oTy4Mr81qfnwUZNRROdvOy60cBf4VEcwu+e8
7LD9lSPbmW97HZqbM1XbQlWablCmbfinP8OpfkToKQMH+AHl7iJEbRCk6oZWwFs9
DnffDPB+F4ijX/Ie7IczGF345OQTYzHc1JfvmN0QY81otxj72R56zzrwoYSXtjdE
nE+4ilfgxDzI6tg6s5OhXypE/aUDrTdyiCvriFKfKl/IQknOEHYH7GG4eg6lh3Ps
UQohQf6RaR0dQimndBTK4k9bxJFZLdLt0ahtRlo0RuSKG7Wg1mtaYg9SnjoTBiBI
qA7flzrfbqFYtaYG2ksvZ36K23TwuHM8b2N2oPhT3SqtamULwvMQKhePLW1DapZ8
OWmB0wOc+SOJVxvSx4YxY4FXCsvr3VBFvuQgy7K9iMQwU6RMTdZvdtZhMuJpay39
RCC8INXAvlBdVM76MRUWOYjH4qFCxPP/AcMi+VQ6rfTdZImu84TM8mih0+xsFh1T
upFTHhrOHqN7whgTGF7K2s+Kl4FD2LVcspdRQl3j3KVK6aV68L967BeQY7NcWFfd
ITl5sezqS1Td5CRBXjh3YyJafW6iiBFzsdXVIz6NmFTXoSd3wFA/S362sQGzRk2f
og4CN/k2FES3W2TtQF4BMSKrnXrZBbWUTGbJok00BnIgSUrDq95RAZ0djIAQsSWc
+6o0JiNvQerrae+2yLTArZosYl/hfjwSCbrHwEnZc/LjLSliP0musARLrCNZQgel
mSOlRawI3h62kxTleySeyayzZeyePn1L5GaJ8TgTezhHPimZcVkrWrqLjYOJB1fg
5RZHJg/WwMJfz1dlEMgRrv9pbYrjsG2fMtF70BbIXXfJdumApQrlLPZ49jtCDp3M
ImLBmS2GaEOXD+a5daRLJzHbKFWumInt58GdH06o1p0S9eOjAESO5cr97+NL0kTe
pw8mhZcwSH+h867m/gMPJewOBh/dDGNNgyZeMYCfO2IX6mrO9S6peh/jH+YhGWEB
vLxxnHMeaEvhfJ5CQqw6dJe/iZp+ubIQhF05ctgFIFFWhVZCLn1ZvevIG8m5vcEP
rtpA8paZS/8/3BPVh7JTH7s2MqwMztiUlhsPVH0FR4Fl2hZZfckkKwGsgO9eTwkf
CA3lyRqtz35Pqe2K/Lu8GmOCpCxo3a0fOpyD1NlyEr1kkEGxOTCw0tMNk93xuWfE
pPqi2AWdQi3NA7iIPTEaCgm6GqX4DpIBMz8va2aFYNAU99HNf3Eck3MpuhtxB3Ei
F6CSHNNV8MFbABilpHg/xl4+KPWdX87dkwYlY5R3Kh7v+dig0Ccayt78u7dOFlEi
7QM88ygD9bFD1Y9jJkyIXK2oZr9vWLaAP0PULW840anHq8MNm02jHe8shwJW/rw4
cNRcYKQdqu/S0koyBqKSSJmArgWLkuR63tyWbEo0a3i1ggc4M3gbh4Z1GjbPlrlQ
OxYEpZoAHVQTU/h/TH9p54WJs6kfQWSSv1djPvtdvRJfECUqs3nxK657COqjSHeJ
eH84EJxnEigs1BHE0TzBFr1jUA0j02/U1I3pYIu7y8RtupFD0j3LdsQJgzxMNpBh
tYYidUdZIYqaCvgEEN0kq57oNKIx/swuLBarX0gfzTIcajw7cVIZXXTlaG7IDT2r
l1NG9P5gj09JhsUSvTm3V1mDJ8FF+1LUulklDXDwRHanH3SNmvBpRfWBl7L98DKJ
a0/79sfaegcKS8JQ2TWwKqqQLK3qo1kFMT9OF1xke9hWiFCVvGTTw1okvFGt4PBi
rjwanoNnVcMp26ehOF8qaRY0htdkhNYV3lY0A1bz5GvF/FjDoOhfyeDIXVEo5KU2
46CreXAQo9BH7KFgrEbCc5D48dON1uFp1qzN8PWOAgnhj06OlzTfwDP1nhTw/TO2
WD5BPGfwHa2LiMTvs6ohVe2h5pmJruHYaQJznbF/50105eF+aAKXFjByXSBKG0Ob
cgmYWZNlXz3i4jmm7sq1LL6CggHyBeG0e3bW0/7DrmyYj1kcEZpIppZaa8QjmU4n
PZHGniw2e4qbQ5kWjZoWZKcdspHHu/Ti86AACyvKOih2bh/LL9LisInNbrMZ0VuM
tLXsfO0RYV9ZjvFCy3qtO+BlTC6vHhCu3g3cCK7sPTUugxvYEp+3w10tbVU4FQCV
c3DyEnBoqxpbwzY0gM5u12V1MDeNMLvFY6xWf7vKsXL47Ws/eIO3exk1A4dGqldF
mq38mZYY0Fh8Nl5ygkt1dXAaZiQT2Q3sHa5RYs01YKVYgjJ7Uwg+Ve7HQhv0zB5o
KGQbXuj294nNiR7Sk+rfnM4VFiqZCOnEQbAvm2UVxZlQ6fyOqp+N8PjxxLjODhHe
CBof3/FvIwSVvfBoZ9Up1edv86PJcRz8XtgAUujH1ZRUSgnwHfEtZSqPRF5eGbxO
PO/1TbJZ8QH6vWD8PMAMTmUaLW1JLAQtUn2so9G6RyCVBnx/gM92inyHI0bkc4Xz
t5RqP6fU7kJ5WPEoM0pAUKzZ3RXCL2AgV2/vXpa71gZSKibxBOEbamH3JNMPrn3+
T63oLfrlToubl8EoyJa17XKFyV/k6Tl9DfZm4QwYSL75rYLtyxUqsx4X+WfO5TXA
Npv0E7SeVkWq+Y2e4t9BafIhmk6cSllzzRmXj7GWRqIuDk9Cv9Wdxp9Hj4TrPlvi
lsz+6QyW5z6s2/TGSJbmPf2IXwG1mHYIQCdzN2Fzj7imAb4knlKvC1o0B4J5C6W/
AauvuGgl5Ox/dSRWokINqjUTqt1KolaxsK6J1as264fCs+NFosF/XuuNoFvNG1X/
UAwX2k4ByYJxGDfZvpRZ8Pt1bAmiEEaxUh6pBFgcAkWxJnqXLxlcla1awTb6cA8E
9eEpPSSwLlRRW1keof66Psaq8GCnzONnEII0rMo+cT6CEeRZVaJmUu1cSNAagety
blZgL5WYVzJQj42iH9XqK/v0yumuxWgiV1Q6MPt+kLyvW2eIKuCGNCImhzZ47UCf
qq8NBaL/2IRQSYTEuO4a5xHyEpjXrQBHq6z/U9AJWARIe9SIxUGJRPF8G0NvjcXD
Sx1955XQ2tZEU2tAZTcR1zONSV2eBdWJYlIeDqvyWT8=
//pragma protect end_data_block
//pragma protect digest_block
IBVGlrk9Usc+5rWVpqHHjYFTvk4=
//pragma protect end_digest_block
//pragma protect end_protected
      
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
LbMk9j1FL0aJtnW0WtFUOMhQuRE3ebYfqvrawqSY0tCI2MYvFoNMiMYV/wIuNCzq
OUa9ySYYPDK+DrDsIuew/uUL6UY1NciSJxBaKZddjK/FMYyjlpk4ZwRz+tLh8TPR
3efyO/Dea1cmOm3NT6fQzo28jmogm5tbd4qkeUmkq+Z6hAUE6Ptytg==
//pragma protect end_key_block
//pragma protect digest_block
AB6kiJS/nO4z0R2FMHcAGY10KK0=
//pragma protect end_digest_block
//pragma protect data_block
dau2EO4dilfNY/2LMaxl8BuwUW3ay7tKRr3ebT+XeUiRosDDZoiIeAZyj5wIGYUb
TRrlQD7KLKEQKQRVoSFou0ZoRH7nzpnQ/MN7AK9inZ5AfYVJBQM7adKIz0QvJA4E
o9q82+ihwTnOCZobSHfs2idp82ubl7Gid65U5cIB+2Zm1qFlioLhkFhRrxV42zaz
Ys/HyavNptCTf05Fas3etgct1QDwTAW2kAXOOmPc0TJgsi8lPNWF++MWyluyZNel
jseC4X0hBlk6AssexRacGBLWsVwtwqS//tiPSnaQkHCsgoKuTQD0U5KJ1jZ1ssHk
mzcz/L1WyO0hLi/qlCSRcagcQB6iveIxPSxEhA27UFIjdA8QVo/wV+tWiqAsYj03
4hzgcw/eWFw4fQtahYfdjXFb9f6pF8OCoXNWyi/D4FoYgQW7ZtmbJWj4fHa3ejkz
NJ0p3yifUW1f+diwth5ohWibx4Cnha3+i5dNeCod3LA=
//pragma protect end_data_block
//pragma protect digest_block
s8Ibe1MpkVQNBjDmtoZssmT4iQo=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
eKd+DJgEYJRnloYpOhw7ThsXG8XYPxxs4y04oDHFZq6FG+6eMfr3oyk0TykPI3bh
YkEfRmZrHVIybZlmKUpOtex4nHMJYJWqbog4/hV5/OG9Yg9h0RkffbLGs1RFkuff
e2Bgk/JsuicalnINjEawiDerjJ1r2gF01RHzpEzYpPOHZYAbnlIb5A==
//pragma protect end_key_block
//pragma protect digest_block
b0nBSHgxVQiijjPd43spkntIfQQ=
//pragma protect end_digest_block
//pragma protect data_block
sE0s5GUfdV9oX+98Wv1Ley4Sh25arShlQL2kO7Rd1b2DHeoWSx/KgHYBVkNWEcf3
aGOc1FRVjth5enkLbAi7r3Z1Nr7yLF7TktoF8te2kGRK7onHmHbPhvENCCqd8vp5
8p9yu/oKtg5MGRDnBcXyrRqbu4kotlWj6Uup2xbYl5Y2DG4jBw5pFnRpsEoDjMpq
FIHEbobz9c1RsHaLlIFrg/kjvkJF74niYxlFr2T3KQuUit5epzwMJN5sCyu4MdKv
ndUsAON5zojiahjKcJA6GzzyIY0/LI0lOAEsUN3S7eBo3ByLO0tUFowaRj9Rb6RE
ugUBVlvENm0KgL9mzaaL1DMnXC9CkTrhjWMe5n5KQdSUYFJApRPDIWaCcEzvsJlB
lVK4XOFfliKZW8Ws2FOEsECHE1X6tx4MxZEO8dbdOoNqM68uSRcmowR16Ccu13+D
DB+NfhhvxSWdswIXWVEQ14yubs0AZB798JDkTJAejaZXxGZseEADB/hi1C9lqDkF
80aqhigNKPSeNKg1tl7BGXaAleGIIqyd+lVzk+wudg/AEU0S1lM/mUwCk8+v4Oso
6d2mxq/waPItGfQ8B7/fv/AC8/9WuDoffn8YGTYEAGPK2wcKjz3ob3Yily52Npco
eKuYnlUirx7EpWkRLam5Qmm5lZI5s1rY/DTOeV15NbAFrx8Oi3ATYJN7Pil8Z4DU
cOEH18r8haEkM8ewzNog6RTT6ScDrtMMd2VRBLejD0fQek0G0xBFiIBCdcSmUsw6
b/w34HQ9tZbo9KrPsXAsaSxDOqMFF8NUvL09uR1pwV2BhEb5PT7AvDxg+F4wHTuQ
ZF57gpzuEEKPMjWW/o5boL8ILAqDm66YNWzXzdjXlANgStHuXsDBKQq2JFJa5y0d
dI+yavmNBjEpStUrwNa3k+8jj3fL4DQ6jOSVbSVbsrxMjFk7zqPg8MRO1QAN/604
kmZFqQJsyhZtDM7OpNL2Y9376FDUHlPuGuasRl+EbXbjdM+OSH+agZDYYaDaNw4W
+xSytyLlPTEfl/e43706jBVoXi2re+2cF2wNPl3lj1B7uPz6UQwk8lne589c+7Vz
HVJLCUeZzkgqBXYvJXCR/fGJLeLCvh43BNM2Sea0BkZBCtcctlpnGEclMiCw6CXr
VkgY8lYRyUrdiaKxrAkMYpilCffrvmwWoDptj2iqxznd3C8iLUiQTjHDoti2tKue
h68s/pQ87eqm1BCaT2ac+6IRZK80Di10p2fXkdCo+/O7Zx9UJobTauYg5OqXPoal
9eLo0u5xCnItcVHqkeOi/b57uV7gBsmRlVG0wT3DEvayosQ1JqFfXQNGVd3bjcDt
shOg05nUUGD0ayFpeb+pdfNOswcDe6QZBTk02yAlu+HRPecYbOjzNztBtHddp4+X
GP8yImMpvyBKZcYBkpwGxuj1+21sl7d100imalnbFR3XjfalE+pJ2fnnlVzeTJXx
SZnZCumGFUPxL5639KFLsrmjw26TcQLHA+tFYdDegtxYeVBDQtXHhWwS8GkxZ0Dw
1fJg9iq6R5VCt9Q/Jook4+PJjGbKKlr5tE0T/kbrhOWxBVClioBcCWAHBS5bj16G
q9KILWECsr1WKZdlKmlnxJFefvt30JOWGrt84tfXNsp22peX0ULXaoKJcB8NllQg
FRenO8CCs00xl6uol/ttzmbXhJ6rXZdo6zbFITXjqzQW14/Sztp4nlnEgyir07Nu
Bl7pBMmDJZU8E2OApzIHzAOlv57pscEvjYlLNGwZrvMHbMcJ3WY6fX/B3QGszrrI
MtkHc+d/OleBTutvojZIUxTWMxRHncDliifp7KRGlyrKT9jXmpDwl8aafNMm2Jec
t/M7c0+p5b/5slMobOc41ExdOVQiqckJaCq4Xuw6C62ykR0LLfBQbrQWFrR47hH7
bXVuoxOx6vOOWlqVLw9fE259/GyfawatVcfVpGA3ij+9yBGh1KpJlAyCbkdbUV2B
xaOniU3+/M6gzSpSqNRBmKkCUIx+0f049QJzJc8kIwMmXn611ijj2+U9e5IoQ51A
9HVVeeP8k6Rhw8skYMoiwosr2ufx+28lV8N+0NktjxMUSJHLcBibO1P3HhWzzmlV
08QnaJgNxluLeo9aIN9g1y7b5lnf/svcHTs/McyTIUcxK14lSopHNaZ3qMa+agEF
Uz0K0SXdT6454j+TbgDeshNAYeHGRb21cCr5FBit0HmXVjqhHdmeJPnINL8DXEyE
459hmyBYfugHLPtms+OQmvbrC5KyDFOGA3S+BhxxUXKjO2+K0IwytgyCNbfdG9FX
Dp/qw0e8KvxrKGS8SIAEmrKybaL3EwlO/fs1VU5u3TuWO2rCLKUHrHsn/+i9CVPU
VL3UbqjJczDxusJ35K6DrILSh/mX+tDVmqBxUIXcTWewWVHQUMEt8ZiLNIuLANYp
uGQSID37gvYhJXaNy7iJ1fvpUb65v+XgUaOZuQcaeNT1Y2kHDb4djHu+tQ+IE9gb
fQ11WiCRropvw2BjnSCvJT/M1ElJnDr4FSzVKBJBaye07Hv3un9vBcncM9Z+j4Jv
Qud9uZ70EhEcEKE0AUKXD4gCDCcDYXzMbQUFv8WWhCT8DGPGCrEJwUuVt49S3Q5r
r1Mq7D41Zd8ryLgMO3e6zaELGiEe15yg7DwICZiiuzAqtVEMex7mjJpJmww3besj
N7FtNr43t5pve6bFYKwGS/ewHDm1ZxP0Gg5ObxIrfqA3hufItwIOyyVG0KqQBWSK
2l08m1utE16B2x/kxi+lsmUmjWvBeYcfmMlUTQB4PRRKiGtAzxk8JFnHRcPxh6kW
3IpGAOz8xyKNz2v6K5WgZYBWq++CLRljb/L3yMN1A5c9zuKGSkp2j4qaGhq1Jyy0
lFQ9mm5h6ppkH+Y4PS024Mfyw1Ke/f+CtA7XKXAgaFowumJNHwJEDAukGcPJZuZM
6jEtaVhzCZnWgwriRq4ionuZqjt5u14bEd2hWTEeh2c0M6xAgCl6m4b3kOaQ8Jx2
OSL41uEdACT81/fSlSVIqggdKJuMbaSjmse2/oDyUwiZgE+q5vE2BhaBhOwiQ2bZ
ZCyqYULExZaz0khjk41++df1jdrJ0St6SD796m0/LNNa9lhXJEM8FKaRnNzbZkej
i0COkyaytXGA3KHAdp6kzGYUd2N8dx7UkXkupfb5+O5ICjPRpw9xds+3YumLxHfW
brktLkf93YfdkJKvfIgawVhTwvXmeQMXbRKL7Z3hWZdPzoXmkbrXLDDVaZCxmiN+
3Yvd9PVN9SF5uRgbGZktWX6sBf9AOCLOmnZJTcdv73+9SWYIIktjtKhJD7FL6e5a
7zJrhzwN59k00agajXYO2hxKux4ucIdZOWtPc4M/ZMuvAyEGRbl9r9hgOhnSbMdl
N0YtS32Vf0eTO8W7++jdv6u2Ybjl7JeNBxXQ3dMqixY4vqFCvF01VNM15CZ/jON7
pKxPKafOfYNvZiBf8Pe4bxcEn98G8Wopn7QBg61sy0VI6qpGx6n03SWUvrk9JPNj
rVxW1tBr8nyMsYo5God9mTtDJUHFxRarLlNx0GDyB7OOPYRAYDX4s/5bkukbr9eb
hFhfLTipXXIwF+3SJyjWgZHWMr3K0+nRdcNhJePtcMmBccEc0PuJom321Guz1Kxq
RjFSl4MEN6+vgjBETY9Hstv4sDPqmCA209VU74fTGP5R2XKmSOnFIbx71ZPOf6+R
JXvmNQC6MX0hAj87pCYNVYqLQHeCnVdYqbNazlx6/sohZdUkqk6pchP/bEOZelqd
E+NnvxNLNhdhWXMfM5S9ZrlcQTjIghWjKHyK+1keH3vHpyiA3rLsLF7jXnI+653D
xpZM3YbUyWsJl5NrUsog5k4sKcPSyRhS6rT4yZCHwnlaKMSuchlKMhv/q5x0BVKj
eNmvDT8iXlYDIiMxB1+XRnVkUWpmQPX7My2MGIk2mZVzNZ9lXnq/nY4Vbw1weo0g
9wPlE7s/z/wSmJ/d9VWglMaiFjhE6zRHFRqBVgTbOUXMvZHr92lq/r0IDok1LfKs
9VKPIpWLstOs5oiorWUSMsJBpzWVHyK4JybZQNk2Ited4B2wNnt/s4TG3JrIywTt
+54aznx1FI+Qpx1fDEljbZ6BZTPuOx0qNlgYwnwBUQWamS/gK7k8PUqVKuLS0q1H
dTjFy/konl7MtX/EofmUN7DB3vdizahQdtzcC7oixjSrOGsQBIv6gmjnPJEn3/fN
LlPsuQOU0K9qlE0wB457zDMiW4QemsqoDw9pftutLEWGo7Hd8yUqaFcgAnc1+KqN
ZjXE4j3lNeh7B7MILTzkPDIGtA/tandjgWjJZz+Q2HtFKxbdks8VlgImtVNrXIoY
pMttJjmUxRMT2lxTNRfleAzmAoFw6W5mXFGpN5FW1nIDjuznmv7pWl+CTa6RCtL5
omfOmBOIH/BAX+BEEX82oYIi5iwVshgju1wbQ8i13Y5vAikbl8072Fp7PhWXzCBG
Xqp9NO2js0+vT/l2LyEvQTCLhkhtXzjM0CL5Kd3W6GXCFmQpgEfHKi5A8jBQPVgW
kAov83yNIYrpB1VH34Wj8fQ8w6VL7qvWCxaD+sayhzp5K1IlLqPBFhikjyY2C3KR
L5qCgWcJFG8jfB9yqrYLYjRYQPVpeLtTq/+QNoMylQQ+R5v0i1eXhGitO+8hMR3Y
zcOqCUdiF71NPVi2Mdq2uNJF5RABXh0SdPH4807H4xPPwNjnAf9Z1COFKpKTDV06
2pVyzCH4+LE7uDnQskC/w/CzNTfNrTHfWqanzBjOO4U+FNF+1BNKorwwrZnpj6oc
OS5/CTAeWRQZuJxzTYR6DA/y2tciIrmae2XEYaPtpukqZQwle1FSXzfTNSAPDkEQ
Y9GRKQKGFKeL+YNw7PZAHuBBJZtcsn/hVo9Xx+qdH2g513OYWN1qK4CemDUeRUJC
L4wPYf1fhMp/Ft/2kSiZjItPoREdkp23rNU/rRq7O2MUmOvexqawUD7hFoblzdgE
Zd3D2bWXYfQqxa8HvtlAkR4QdQNpzb3XOfDonI6ok6+sWTOwmgwcL1ZnSPfnOU8D
jmkt+zIt1w/6uDefvj/v1AqPpcd3ozencXMjNLdn3Z5x/62xGzx4fLL6Ygsazcnp
jY5uTcL1Q0ZZiKH3UCzTu/y8P0I1CwwSb1uK/AwEUWOiNv9SH6aXDWFpkdmgtQDz
Meh8zqNziyIBi7yW99/c76rhnyXPqfaXDslddSN0c0rEBzRVWV9x+Gi/YV+Cw/07
XouH86ZxyH5sC6Sz7fWXRr5e5oY+ly7rqi6h0JUOaDMrfzZyeF2NOkiJQCuBtrhY
IfuI7z0/oTbyrbfSc0gR89EAYBS4zfyLgu8YxgK+X3hvtbVEjR6zxtM0nJeUNuCL
z9AREGvWcKWz1TTRGKeLj6DI3ur7vS/FUWmQEBwuV/lH6WycC/fu18iZnTEvFfPv
cVUHW+yp29/83z1BNykAqdFvQ9NkdFBRRaf5GMYURsy6BwnB0oxYhSYuyCgMgR/2
ypou21o0/d1CUmmQjw2ssnsI63i7SlQll6k3dF/Rf6ZDX7ZC6Rxzb2lTr6X5VRnF
Ri3C8NwolLjSKGWMRPqP2C92EctwKTdpqbjba2cb2abVjGCwLDwBBvvbKBfdQlHF
U4k3cZiByNCfa7hcTFYMk7qWzq5DPBjywnwhR24HHtkifLOPWp4eHFsu3lPx9Mbu
L0AulOHTk5YjFdjftWpWIFATMuJSp2fjtRuPTlo5iKwCghXye/TgzTkcLXXs6KGb
xSmztIz8cz1B4CQFqLkL09KjVMwzmDX7s7pm1vOus4IdT6yLYSt2DAa5HfmJO8fN
xqBuGNjviVNiraYr5VY+SGDG/FuUo+uWHac7PW5r82hVhLOpYA6HO5CWShX7YfF/
L73JCIOPzexNCMqhKCr5SIdtpo8Ijv48dLSC2b8siCZmfPbOWGWMR8uUOS0tuMI2
GZg7lZ1j0TNqBmMSQD7qC4bGmINwHaJBQs/PEQyP458LAdjBq+CsKk6IHpNgkd8h
ioc5weeNvaw9ER/XgfpzZxljscYAznnaodygVvsBhli3he7GAbQEE072dl0eX0MT
EyxjqhMsGtRQTK4oOXmqf8W0hO4dNcAtiF/StjFLbKOuq9YJR4Lrwg+CuJxjFtGt
O0n0rs57qRasH0nCXPukoyctpDnYm0ll1mok6uo1Po8INCiA8qDIGp8dGoV4TrcB
dzIyvs918DOJybIFnjhWQGYUA7cV8WLLA88emshttCIWHNI95S5I04ezonPvzrtt
5dq742ZOLulGnBDO9BpZgM9w71FFlDSd0JS0qvXe2fMWQJQQmWw3f4wHoQezzRDF
zkOkODM25ehquVUFARoTLpp2qja/p3KsZwy5nq5bkxzVFSutQGDCwXfd9Q/MnVBt
cn6/ju9G0ABjnZ0m+2CDN6ThWvhlC5U1H5Vmren9TDtPwAL+465EEKPVgnVNRKYm
kFRJTHg9Du8vc0kNqCv0+tNQ6jz+p1YDxKp1tQSemXfDxGEONScYJYkEw106LOnx
DVsC5ceZkbW66++Jodx3KJI3pH4C/Auv7T/Stlzs4PQbdQ7CCFuOLlOHa1GUDZjn
yqkJGp/fRmWrLHvgSrKXbKMql8u0CVIPrPESD59exJo0TeNVKzZ92M2kiZHegnCT
trLAkJtDYHUFxRw8U1l8PT26THcPgQ3mDNgUEsr5uk/hnAwQQlOHQvXPXulT8xOC
aiNRSclylFwPqO/+TTXy8laLyy3tePzzjxGzOzB3fdO940cmU+rdgG2SpA9PMBTc
4CBi5wmpTarRWuZw2CER/GYrBA9pwGDJtAk2ew4M+GkoNm8W3KOnZLS91+5nexfk
YOlLd73LoptanOwcqFANANQY+fDTD5NLqWD6jQaR/qOziBreAHldBAR3p1vg+laN
cni0El7ZW7xaUq3hfsdgHq+NoPvgl+OkVQrbp7dQ19OckSu42fHCfh26ClK7AEui
KTTSZ3EnTwxqZzNwJMkxhkIL+/m2k3ZNqcXoPYacsQp1wNjnw81/wUXMxDx/N+C9
AQBzYV7wHUNXf7pNhYI7FBgM1zdHV1oMb9m4uc9qr8kOntEDpPYcYDxUquMGkhP6
/gcCigKMY9RX4oWdQNZ8VK1QhAneFvSJeC1U4709f17aLQ05V3YvPZ6Ym/QxvyXB
YPPmKw1wHdgYU0/iMmehsgC9cUkU6U1U47Lrg7tjkqSpHE1tQ06EIa981ca0KpzH
Saepm8KmgmCmd5N/VrA7WPfxaac8KWhCjFCVbjj5nAQ81u1D75+ZhBNHlQ06Aau+
K9OXEE1VUWbw80O2a0Nb3FDfqI2tw0hF1JVo9HGX31y9PztkRGa2Ny6UvRgwKVFU
lFhY0rSwBsMKsRu02a02MQTOapGvhIzw1B4PzmFnxSUnFNvRBT2wcj8PLt+51pFN
uhA8ol3R5pXUo6DHf+R8OalNfXDXm3gRpXZ7IcG6YFMNzQ6dsB/ULbKCE1KsoGeo
aCfwuJJ8CU6f7JT15EUOLDoEcDZYuLGAGJDxnH+3bkNpAIOU5J6j+ZWP6wEUQDzH
g9BSUS3Tx+i1a3ihErgqf/pxVEQpxZ3/BbO1rnrrtLcl5mkUO4oAmaubBlGrD6DK
9i4vbCFTENx6+9SiMId4iWrRJ4ZjXRfKpn7L6l6qyBhwHZpht28+SAwxLdraF2lf
dWzbs8lTc4XRQ61yGtpdR2sePpZvhKgVblnnoQlz5ag3lzpb+cF0OJXUthQ0wtZU
77CXvJ9ybbGwKzVdnxxe2LdgWcc780DbhG5amwz3g1iZjamY6sT4aNvrdXYTizo/
VsFyC9lniGRuegQXKIjhnTvi1D5i5mowrJGHTFaN/5n6SAR2iXJO3QIQfjmwe1Cx
HYPNn3GzaVXPBNqy6QrJaTWBXn/ZOPFy9BhYbNXdYc++ggln49StOedTV+OxNhVQ
2dPygc5s82AXCmJNs46CnYZCLxsK5tdCTY4gkLHz46F3hUmnCMewLHpzdTuCdyqs
PDAVD1wqhrBZj6aOJg5XPcMFLE61LtpRgPnYl2dobbAJMkJMIQGImW4a0mDGVOTM
kuzbBnddGjz8NGtE1Pp0kH/jZhryIg1JC/3e1Z1a0LPG1dwmE4yxNmrZIZ/Ne0HD
m/FxX07u6LP/X2BtsTQ/XyRSV1WRxok0EysYn94ZY/Owk24yd3zaqaye7Uy61Mz4
sthrGujTX+h2FcpxQcwRm8KE1L9MZ8I0xl2DEXkA4/CjSDwoN/DrnSvVohgV1PTy
ChlD4Gm+HVCqqwK9zJnSKaUku12MzdWJ8OhapHxcimP8wB55u4ebkkvkLFO8Yx+0
S4SbEujqESMFN1qcxjVbZh4OBA6VmVRWOkCw8IoQebp4y1qjLqeXWjelxyUmakuT
154+uvB6FSs7yeMTeuJKlX5+nyXmj8uzu/udZPUl4qKtI96u4kktd0p5BJeplUx8
egj3cerIZm+bhtvKS0LFsabbaEG+/ZfM/3TuhKmvzUj2uLBnsh8qOpnzAhttNGgY
MH+6TJa+OD8kut9lrzrjNCRZ45lvtE3Rh+ZvRn57A6tDLPYQrs99pbYtkYCq/BxN
Y4D6FPBwsQysvYRsRY7uU4Lnju5AMKrPhKUoxxbztJr/n20dVI/48H6pSalxKYf6
sL3TM9F6Lkl2WjiBjswrSBUnfh5zgVNMlcAvIUI8AyS+ReWatT0NxtFuZIjn0nVy
wEyDgPJgR1Plg5IZorko7pQeSWUk3xnSEmkKmXdAjoMpd22L/yAT+bkbFCIv1gbm
HzmS7Hu5fh6xBYSMtqGFZFBXWkiGJii6WCYZPA3k82ctE8JImJOQeMaYn2AIqnZs
93zQKJH/g2IeL/cnk6U7Pi8t0i58AyIO048P2is4bSv14LCmJS164HcAtbmO47AU
Ilx/GLbbTFfosctmq+WFTMPEUo+FL1VfiIoozAeGCVzV+SRrJV7KGPbnzrSjnmDh
Vy/NmxtwGNyFZEViagHuCc48E5p7VAR/HFZGm4D0YlH+2sNjMSoV0VeXYiyfsR6z
ahv7Aw88JRnauzahWduRaJjO/PznmekWXPlTrQxX2gY9/25UUGoXUHdMtRUvjP+Q
FS+ZX52MogEIOA6e6HISRaSHEU+FU2wk+QPYKtcDiFRHYN0AMUfOsdKGgw97ic2Q
IUEcgX1/u2cjdqLyxMvpszCgMDSQoD1zAjLg/ZudSs5IXE544dpakEp5EMT7RSC1
MIrXReOmeYDUw7YptuX9sIsboQlmwMt2JdvE5ncNQMbs+DkAviFvdNB1w614qHbc
swyPoioCnt4RlnbzTDA2vltUl1fAIFzkPSUaNd40HnUNBtJ42B+O2oARS9IOcRZV
W2tF4ZkR+85/NuCUy7XdmCE9ajJG5jzrNGGVBoxDGdl9QsOQB7xwsQ9ILrryxRKT
BDZg9OAFoc2U6QOWxXmhCRf96pj8jK0DgMblqCeZm7u7o+IhbwDaWva4l+QXHwfR
VZ44kIZpSkT1j7y8vgJJGy3WgERI7mKP8Nrcdsq6hi1FrQ/rjShVhgAX5aFYosoB
NOpk4lGWRU55Aayt2F897hf3ZHYNc574n+vKdIfzM6XTx3bsAhoXgWShGuBYSdy7
m6b8MlqLHLaAVn3Sg7HkEvRhX7SFNp+6Hnx8FEvDLV8GDeZcQPkvsRovVUa5iLEu
TQwmzeqT0+UUeH/gYItano1bIcN+OLWAgroeYewfkJexdfShUM+lJPUyH0zMwdUf
T/8nk9xBVqieqskc37rGhZglDDc+yppCB1QEbbLNMyCPHnCvB14aaxWi+h1c7oRD
ufBPT2lEvbEdVBSGJCR/tcnk9bXT0XOhceODETQyFpEuhYMV2UmRC9k7tG/nSbwf
H0WzGFVFmECs7OyWWNKjpuAqBSH/Ljy6huBfdeK6MiLeozz4NCxUIg2Jbe8U49oN
TSU/MSSdDF5LyC2vzNPF3RNm2qDRRYBmmWCHeaiDDgjwnvy5sZJConmTee3umwTs
Sd6gvyjAHwxYXpYtYBARbB8z4wQsgvWKrjjsSUQFuhu22mhFzZGkJOxBK46rhu+P
oSfxVWftvfNKE+XTtp5gr+0ZTEwO7J6CSLYEetK0JpXlB8PCeS2zWl+vd5GZ0h8d
xxndCOcXeS+If8vyPUdM+AlGGjDyI8j6JqoveuN1YP+L51YN+eiDhG5IDFs9Mspi
QuvemdOLDgiXFD4OlvBPMpnVempoR1pyPmANohRk09H6ic9qhMrILeS9K6DyHkSr
6J5Wa5vZ+mW1Y4n7e4YSCL0KxguDbsFeuMX34Sb8t/ajyVTOgAiNvcqYa7hRK1rF
fYQ2CcqKjKA6RRJrTeyQfwEq2tU338xvegNEzFmFCKpiO8Ko6P+q0x4zN3LcN1Nf
rUX6adJnZ3eUtz8aRMAErOslwsnc0GVQNNuJ+8uMr9FdZDhm81Q1a3HiLrjNemcc
1asuryINSrUpGLZf4bGoPA==
//pragma protect end_data_block
//pragma protect digest_block
lx5mEjRzLuUEJoiBCWObc3r3v8s=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AXI_GP_UTILS_SV
