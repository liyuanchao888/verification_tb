
`ifndef GUARD_SVT_APB_MASTER_CALLBACK_SV
`define GUARD_SVT_APB_MASTER_CALLBACK_SV

/**
  *  Master callback class contains the callback methods called by the master component.
  */
`ifdef SVT_VMM_TECHNOLOGY
class svt_apb_master_callback extends svt_xactor_callbacks;
`else
class svt_apb_master_callback extends svt_callback;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_apb_master_callback");
`endif

//vcs_vip_protect
`protected
Ef\B2364ZdODb;&b,UDcGSVZ#Nb#U(AEA^3AgdaC.WT.21g_[BG/((OHE+;d;egR
/9FgV82[2Cb4(:fg<Z^JHI5XU-02&Z2J<]>B=M=ADQ6<G#IBCQ4a;f1QFI5([H)0
5ad=+,<4_b7Z;Z&?C,/[E<:)MVWg#=X20)8#?E9a;2-JXU2_Kf.KYPF#1J)Jc/[P
RW^#MMD5F(ONVKY(57^44A&,1K^H),\/I4f/8]A6=.c.EZEV,e3[YdZ?TZ-_3[bU
HcLRYb&ZC;F,LHFKbc7YV@M6Ze&:a#8-?102O.>1[Z=9V0F6dNE[=63NAW(QBd&0
OeIIU2CKKOJ^ecO.C+V<O+E#_Zcca;dK^;=>a3>US<.#\e^LCDQFH0c>##X\>FO?
F\a?E<YYH)BcJ=IM)PH9_I)2(V_;[75XY>GX:f=BW(K.L2:GW:bGWXY\=&V1]SKZ
2A725R4/;V_ZIW\fWC,&C5GMYeZFLI[DZgVKb.2USWb6=WKLDF3EAeH4.c3_N0;F
=#_2ff:BNgD8G(dH^-d<B#f:d_DO<6;QB4775@LYgFbMGV&P^<GH;K2^Pe9^f&EX
]K;]GUZ_/_\FKPX3>DBZH_c1-(b_0H/ScgI&5?,&E;2WW8PM<J&A,0?>N_0M-+21
KE0IU04eT=->#[OQTFgA^D,<c?V.,>7JM_5@E-BY(ME+e>=7_(NXWBMe7Z7Fd@PH
YS?=8U2H\GWf:&/,1;;c<W+L>-=L-O#98=XaE>10(N-8]?5fO+C9<GTI?S?J)GJc
a\f7W@dV]:R@;BHQNMAR.18@5)6Ra>af4@M/BC(@1ca1WRSSD8N48I4U1G=BJV1\
>aX[V[[6;,^>K\_Ha<60KNFK,\OSSaP8<UT0+O_AQ(\^RB8A6U,a+<eIcc)@g^73
(A5&U(/1UK83)_QFV(/I].4Z._10?Q(KCP_fgbb3-B\>^431W-&B/?dP0SKL46?L
@PLJ,KfQ;YM]<O,WSNf?X@D@V[Zg)?CG^[I<?HV80V6;^7T?SA^S#EQUMH+N&X+^
];F(,U3Qf5E^af1JL\NVK9J5&(:0A^b.:F)5TTaIAC1bCAg7(/N]5.9TJ;#Kag7>
2DU,:&7FZ;]-0BG1CW=fQGA3D#6Nbe)=?6a=JA=;)SS1;4Rg:QYO4U+g?NYEba2X
B_9OV<<&1g63e&cPJ\L\;?.Ab7BM-P[=7g6@GdW;gO::1OKGTbO.[Q]#,e]G4IX7
.,W;23F9c(27)Y<G0CO:W=97_DEUHKRLaC8;)6C;^TQ9b:KIcV;c^Tbg)N[FM9=I
_1/NODFb<__LT2XBaP9g:b=f[.Y/X2U/FD(2JCIMg?2O.f-L2_>0,E9CLaEN>(Dg
WX8R6B</ba;YH:U(?Ae3Y80_#GNKN9=d[W>fE.b[@/\KJ]R8?REf[1gQ8BcV[0&M
PM?\K&Wcddd7?@?(b3GG8G(5,O:?F[YP;HSW8_&,6@DK>VY&f3>>JCND2N.]9c:&
B#/.CP9+J-a&)#+]S36>ZE^01]d^18[5+P+acVb9=GW:G,R5X&4MQT]0aHD7)a@)
&?&.JZ<@Gb=;@2L)MQbIga^FI:[PH6.PI]F=MU]2?^6P\6G.bf#V:;IG5DN@B54;
:/P&N)Ie9T]^Af_d,f=b4^<OZA)2<3KE.0XSY=J;,9SN^8-:]IFA3d#[Dd)_4I+I
)UOcB4\XSQaW8(G]8T<JEL38BUadb7?3IER5Z.F^X-CF1&a_\4HH=efC=AK4U)gc
C0OIBBcI25W^E9LDAMdGJ>HN-gdfOP+^X(^SQXgQ=?(8>c[,HQ-^HI7:O_@Lf.dM
1B+EgACZ>T1g2B8\0-)&E8(R>f^HIWKPG3^7X6]+aEZ[31#KQgNBd4&SF3g7PG:7
X8-XEg5d7.B)g<gN7J6M-fb_KI(D(76ZG\PKLV:-6\9&CCR&>K3:V6FYBH11aC:/
Z:G&1)=_NdB+FOONKCIPBaB]\54TIg8FcB^D_DXa?<T3C+K)5LXIPL)NB26G00L<
PgY>gBaE+YcA.UdW.FA[9\4M1Q>GA5_F0O(d&)E0HA8ZGA6+DXWFKg@+:f)?HBXKS$
`endprotected
  

endclass

`protected
NF)A>5JQ,\f0@E>&/#-gRZgIA8T\bV]C/6#U,1]Tg[,^8\EI(_QV4)SMIELQ.D=P
)0A<S#;VfR=W9#^_L@EM3f4C-]De3O=1W^H,YH92ZH,@9aV-JU#WV^=Hg.F142J4
H44gd3Z8J&2(T]=4Cg]Og5G6,1:[XSb_CdN[0fH==?dGSX?&FH3BdW2?TW[/ZM/_
>RZW[L8OHeMfc@/0I0]@)bNA2G[JS)#,S&Y84&:L<\5NZG<+4Yb)CUZ(e+HeZMG;
VF/G3J@+S=;\24C7&NS#?Ld=/E@\BF?=:eY+Y>4b4;>b/F78Ub3+VfNdJdKG^HTH
Y<TLBLE1X>B)efZgC0,6S[g6#]90;2^M@$
`endprotected


`endif // GUARD_SVT_APB_MASTER_CALLBACK_SV
