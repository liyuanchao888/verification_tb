
`ifndef GUARD_SVT_AXI_TRANSACTION_EXCEPTION_LIST_SV
`define GUARD_SVT_AXI_TRANSACTION_EXCEPTION_LIST_SV
`ifndef __SVDOC__
typedef class svt_axi_transaction;
typedef class svt_axi_transaction_exception;

//----------------------------------------------------------------------------
/** Local constants. */
// ---------------------------------------------------------------------------

`ifndef SVT_AXI_TRANSACTION_EXCEPTION_LIST_MAX_NUM_EXCEPTIONS
/**
 * This value is used by the svt_axi_transaction_exception_list constructor
 * to define the initial value for svt_exception_list::max_num_exceptions.
 * This field is used by the exception list to define the maximum number of
 * exceptions which can be generated for a single transaction. The user
 * testbench can override this constant value to define a different maximum
 * value for use by all svt_axi_transaction_exception_list instances or
 * can change the value of the svt_exception_list::max_num_exceptions field
 * directly to define a different maximum value for use by that
 * svt_axi_transaction_exception_list instance.
 */
`define SVT_AXI_TRANSACTION_EXCEPTION_LIST_MAX_NUM_EXCEPTIONS   1
`endif

// =============================================================================
/**
 * This class represents the exception list for a transaction.
 */
class svt_axi_transaction_exception_list extends svt_exception_list;

  // ****************************************************************************
  // Local Data
  // ****************************************************************************

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

  /**
   * Array of exceptions, setup in pre_randomize to match the base class 'exceptions'.
   *
   * THIS FIELD CANNOT BE TRUSTED OUTSIDE OF RANDOMIZATION
   */
  rand svt_axi_transaction_exception typed_exceptions[];

  // ****************************************************************************
  // Constraints
  // ****************************************************************************

`ifndef SVT_HDL_CONTROL

`ifdef __SVDOC__
`define SVT_AXI_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
`endif

`ifdef SVT_AXI_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
  /**
   * External constraint definitions which can be used for test level constraint addition.
   * By default, VMM recommended "test_constraintsX" constraints are not enabled
   * in svt_axi_transaction_exception_list. A test can enable them by defining the following
   * before this file is compiled at compile time:
   *     SVT_AXI_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
   */
  constraint test_constraints1;
  constraint test_constraints2;
  constraint test_constraints3;
`endif
`endif

  // ****************************************************************************
  // Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the instance
   */
  extern function new(string name = "svt_axi_transaction_exception_list_inst", svt_axi_transaction_exception randomized_exception = null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the instance
   */
  extern function new(string name = "svt_axi_transaction_exception_list_inst", svt_axi_transaction_exception randomized_exception = null);
`else
`ifndef __SVDOC__
  `svt_vmm_data_new(svt_axi_transaction_exception_list)
`endif
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate
   *             argument values to the <b>svt_exception_list</b> parent class.
   *
   * @param log                   Sets the log file that is used for status output.
   *
   * @param randomized_exception  Sets the randomized exception used to generate
   *                              exceptions during randomization.
   */
  extern function new( vmm_log log = null, svt_axi_transaction_exception randomized_exception = null );
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
`ifndef __SVDOC__
  `svt_data_member_begin(svt_axi_transaction_exception_list)
  `svt_data_member_end(svt_axi_transaction_exception_list)
`endif

  //----------------------------------------------------------------------------
  /**
   * Populate the exceptions array to allow for the randomization.
   */
  extern function void pre_randomize();

  //----------------------------------------------------------------------------
  /**
   * Cleanup #exceptions by getting rid of no-op exceptions and sizing to match num_exceptions.
   */
  extern function void post_randomize();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to. Differences are placed in diff.  The only
   * supported kind values are -1 and svt_data::COMPLETE.  Both values result
   * in a COMPLETE compare.
   */
  extern virtual function bit do_compare( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );
`endif

  // ---------------------------------------------------------------------------
  /**
   * Performs basic validation of the object contents.  The only supported kind 
   * values are -1 and `SVT_DATA_TYPE::COMPLETE.  Both values result in a COMPLETE 
   * compare.
   */
  extern virtual function bit do_is_valid( bit silent = 1, int kind = -1 );

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Returns the size (in bytes) required by the byte_pack operation.  Only
   * supports a COMPLETE pack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned byte_size( int kind = -1 );

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset.  Only supports
   * aCOMPLETE pack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned do_byte_pack( ref logic [7:0] bytes[],
                                                     input int unsigned offset = 0,
                                                     input int kind = -1 );

  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset.  Only supports
   * a COMPLETE unpack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned do_byte_unpack( const ref logic [7:0] bytes[],
                                                       input int unsigned offset = 0,
                                                       input int len = -1,
                                                       input int kind = -1 );
`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Gets the exception indicated by ix as a strongly typed object.
   */
  extern function svt_axi_transaction_exception get_exception( int ix );

  //----------------------------------------------------------------------------
  /**
   * Gets the randomized exception as a strongly typed object.
   */
  extern function svt_axi_transaction_exception get_randomized_exception();

  //----------------------------------------------------------------------------
  /**
   * Pushes the configuration and transaction into the randomized exception object.
   */
  extern virtual function void setup_randomized_exception( svt_axi_port_configuration cfg, svt_axi_transaction xact );

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object.
   */
  extern virtual function string get_mcd_class_name();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_axi_transaction_exception_list.
   */
  extern virtual function `SVT_DATA_BASE_TYPE do_allocate();
`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: Provides <i>read</i> access to the public data members or other
   *              "derived properties" of this class.
   */
  extern virtual function bit get_prop_val( string prop_name, ref bit [1023:0] prop_val, 
                                            input int array_ix, ref `SVT_DATA_TYPE data_obj );

  // ---------------------------------------------------------------------------
  /**
   * Add a new exception with the specified content to the exception list.
   * 
   * @param xact The svt_axi_transaction that this exception is associated with.
   * @param found_error_kind This is the detected error_kind of the exception.
   */
  extern virtual function void add_new_exception(
    svt_axi_transaction xact, svt_axi_transaction_exception::error_kind_enum found_error_kind
    );

  // ---------------------------------------------------------------------------
  /**
   * Searches the exception list of the transaction (if it has one), and returns
   * a 1 if there are any exceptions of the specified type, or 0, if none were
   * found.
   * 
   * @param error_kind           The kind of exception to look for.
   * 
   * @return                     Returns 1 if the transaction's exception list  
   *                             has at least one exception of the specified type 
   *                             Returns 0 if it  does not, or if the exception list is null.
   */
  extern virtual function bit has_exception( svt_axi_transaction_exception::error_kind_enum error_kind);

  // ---------------------------------------------------------------------------
  /** 
   * Utility function which generates an string describing the currently applicable exceptions.
   *
   * @return String describing the applicable exceptions.
   */ 
  extern virtual function string get_applied_exception_kinds();

  // ---------------------------------------------------------------------------
  /** 
   * The svt_axi_transaction_exception class contains a reference, xact, to the transaction the exception
   * is for. The exception_list copy leaves xact pointing to the 'original' transaction, not the copied
   * into transaction.  This function adjusts the xact reference in any transaction exceptions present. 
   *  
   * @param new_inst The svt_axi_transaction that this exception is associated with.
   */ 
  extern virtual function void adjust_xact_reference(svt_axi_transaction new_inst);
 
  // ---------------------------------------------------------------------------
  /**
   * Searches the exception list of the transaction (if it has one), and removes
   * any exceptions of the specified type.
   * 
   * @param error_kind      The kind of exception to remove.
   * 
   * @return                Provides a handle to the updated exception list. 
   *                        This will be null if all of the exceptions have been
   *                        removed or if the exception list was null when the
   *                        function was called.
   */
  extern virtual function svt_axi_transaction_exception_list remove_exceptions(
    svt_axi_transaction_exception::error_kind_enum error_kind );

  // ---------------------------------------------------------------------------
endclass

// =============================================================================


//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
zd2IxiVcB2bDv3w++wlvS7IkDPHd70tFRcZz/aPpsEYwwuEKm7SDZFKjn9dBwfyR
ke6kwWM+te6uSAeCy6FMZ5VIJPLrQAd1aS+ooS+WP693YNXGX24fE5xWCI18/+Iu
+/HjVBDL/Hp1k+k9cpShA1FgVZGy9+/oLUeDszU98lys/xIrE9Gumg==
//pragma protect end_key_block
//pragma protect digest_block
4PZN5XEqOxnjcuj2u5lVVXsXWzs=
//pragma protect end_digest_block
//pragma protect data_block
8dGS1fWzvoxDaJoVWuG71epfJmfeGwGQkKRdK1P6TKqmaPte4nh7qSShv+M2pTTH
B1ERjj42K42TrS3PW47DZB72gXdTFkpMNd8pQTljoOSpHq90RmNyyfl3zU1ejG3l
aH6+nFWBAxeyb24c0tn+aRrmILN7aq5Xt7jqPNxHuLrw/GuYY0kvvfFM2X6BSuZA
yd/AVUCaSjnzULgrNo3gOdc5GzVZEygQEksxn39RqvB+0NDCx6f422GFtNz9hve5
OyDdYxmjWsB4LpowTb+NbYJMlhw5I9FriS4Siv6HR8en2SrQfsnVVvXiqY2qIoJ3
XJO4NJGt8vd/LL/QTPZc5bB7YZDNdgjVEi8WG+UM35AHGZJwP69lTO+HwG2A2L+G
YmUyg47AZ3x+WuR9HEmMRN02UIpI5qrMiyrk5vb/RTOXUBwWqsJZ5mHR+td7rn4I
ytCC/9uCcGvD6GxUG+D1rUBLpLEI0pF+zEZbu3Ne6L+Ra6bVdaGwjz2bRh9rlQMp
NzWBQFf4T/bk9+tpuUtRNHRowzStdyRa0m+tSwkB7R8lCSEyitH8O7GVMkyp7Nhz
4cX43HZi6o62FsixWgUrAE3nCHhI2EYEhAjMVLV/MHsTkJSdE7sox2Dr7jExX3fd
Kr+SaTYK5OpVe7stIKDOBND3XeaZn5oFqhhXU6YjX05+kFHknvaoKameIo2YSHNj
rWnoPYMQVTEeeG4WGutIsrp8y4iW5+6JMs37mldJrCaorfBHAeYtie1qR9e5f5Yz
jBWRHGQ9V7A/eLqNVVjZBbmbN851CSsOVsObh1xYfFdlIq/dWvRxlWz3wUaS5zA0
lUhIS+hoS9BVwfVDcvrEhelDaOFGBlRHD97PqCWOMC/g8Tz8tfNsP2WzkLKIM+Ur
N3Mb9w1J6O7BLHlZL9OY44+qHoy1NZv3zA/P8MgCmJBjukoPJeKjEJe6wIiuTV/c
3axfeTPW3huKB13Vuu6xJpVhaibW4ekVlGZHH+B5+YuNRxUWUCDNBG6Ttj+0zNBU
T+/JGUEn5VWT2ElyJ0PrP+OAM+Hq6ehWgrWlirv5uU7qVUjLbHm0qqUiK1fDCpmO
NaDoP8OJNPqAH7SCuwvOJOxkn9d0BL2cDzVvw/SOBnFiZMAkBvvaVh9hWtywhls5
75oVtDBxfUqj+tEwH9s2+vCn9jriOXCDs00dB0tg/Disq4A8yRhfoEqTzUimufje
+RL+okBqsehCMZjtJP7mkuO2ENGiLfRxmvFY+hKmcaJPIo+Bxsf6XMhfFcypJRdX
UrB/NiKdK1LLB88va7WYxXN5tBAtwuBQgLSQW6eCB5PQK1V9q1X7KRQ6itG/i4Wo
PWlm9bUjPAr4092KYKSLWU0J0p4lhyQaOjEOik4so2J7YlEX/+rlwYcaR/TA00Iw
Bm0fpf2xdHdRagANdXKi5A7B3Em7ikqZrWeSqR30E5uHj4GNRk79D3TBC0zgN7No
UyciIy6uI7pqqilfH6KMBxvCtv8AJ8vboI/Qha5HOBEuduwvmdw/zmRvhTUZlmOk
0MNo9jrx7zUn2dXQQu2D9jz2/6Mn8ebpe1GQh77ez28yw6WYkeY6HinS+Qihu59W
y7xMYkI1/Ra38P6qyPWpoXhtH+ErEROmuZhXPxFJTJaK02v47E4lRkYGKKaQC2Zc
vDho3zSZ2nD+w7JsaDNJOmmfMPbVPZx4R8sHDxbpIykYjvI4SsHrbP2CgMfW1acO
lyGnDuyjHutrc/pnPFMzaRh27vq6nAIt+vElmSO6jNUZg4A0c/FNrTkowmoKZLvX
249EeBe+rOyFycvn/pQmi8Iy8lYOg2+XnUEvFGiSIyr/8SjpPm/Ter1pHRQZJjcp
yAAVExgapK+ISfAaA+YY7ZcDo3iOp1WFds8easyirwVROlGXgRabHEphnFpTQguf
zAkMfnqXi05HMMGEqpVbvtU1R2smTdEqqFgHo6HpPVRU4pvH8/wESSz88teQDMAf
FkSlzu3xQ25JUn2vyXRcVw==
//pragma protect end_data_block
//pragma protect digest_block
c/oWTWgouMHNdn4N5P3RUstCq0Y=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
LObeb2YClbnfDppCouXkNByR+VEV+Uj12YDHVnDEVj7QCou/+CHFNaGYw2U0pjlu
s5FRNsIYPpGZ+ngtk+cVaQTjbNSfLMok3u+qhzywj1V8xuF85n2yqPjinnlqB+bv
y0vbL8xqahV4YlSRD1/Pd67in3CCLz7p1uGJwYkXaOpp3aDxBXU+eA==
//pragma protect end_key_block
//pragma protect digest_block
6iosEP56zyK84oYLy+MRDUyy3WI=
//pragma protect end_digest_block
//pragma protect data_block
RL8A+8Z8E+cZWAFRBuqEPSOMUvE5Pfdl4RjSAdy443jTdAYYQWHKUCrOkF+BpvEZ
QFSarJKekx+vdQlU8FH5QmAcl5rzdVfTe+N18T6hj1GZ8TaFL3y4mN1OlFQdML49
Kki49r5oRG5cPVHksXtyUJWXbIQ+A5CCxGnFn8qTXCsJ+lQ0TZR1fJeWskhldJx1
DEWEvLRZMvdtln4tbaXAjUU8+OF5qiZk6AjF+MLhnI7TVZXP/3IzpgAbFKeeZIbc
DV/gFuXYDjur2q78xZgOLxh+sM9rsIhtJMkUeTNGLPSgjFNDPVDUmKL2Qfx6LBk0
B9/Vgzm0ElxDNOJ1t5Qu0GVLDac1lOi6LIO9dhLsH9pnpls1Mv5ChucSSWvswZET
XquSNkmNLulTpSGSVrKSV5Yi5U1XZTZTesNPfKwaDV42K+9t3jTwjIQjmtrzAoG7
b0Uz4Yqwd3hSHczt+FXO2yVYPGslQSURWDpYEjMxWyjDSn0YdQ7af/hax3qVNd75
D8JXF6XvNoiwUtH/F4WQDaj9XhunY1gN2/ilf/XbO90BPop214RHSoQP1JJcocV1
N3q/tJHap0Rfn9Oaxpw/Mh50Crhzd/J/u1JvW6hyRS2o3q5bMHHuYZyQS51h9cQ6
237aOJrVDY3j/1Z/OCsxeeUgjclumcz9fWLtVF4BrHpT2SE0q6Ri5+nXJlKjRu/P
pTsTwYphY9r4gHWoRDbzTOsx40Juv5x+TPUM0pAx3eTmFRKRRGPrpvXMQIWyQ+ZC
0ArT7IXrp/jD1JrqURg2/gwXvJ6OFhtbrKghtkLeOHAJmHtS9J2Kbcgzl6Gk4eV9
qC4rPgyzdWJAutzT0kc7B400eNs0DsNsY9ZfjdbjvOeC13CljqY3ga7Oaxt2PuY3
iMg0v4vUrCcqFVerxhcv//W12IJR9cD+LROjgXZ/tYRlP4HGavsBOvB9atD5WYfc
065cAZCrIhob7e5FccDgEHq+KRe4owx0HVOdxgIG7o/fkUuvJaxa7t1FB4yxgrqC
0g3HGoyVro6k/f2L+RSSWyO8+bl2LIeGwndVocVuVnpWZw0z9SGzM+x9yCqHO8ct
x8b7R3UuuMBYkrT4RlqU766jihXQGz9c9Lrg13NQUCRPtNNE+8+JZAv6GsI4crWq
pziGFFWyu/kCvhYCUgwCIHJJ4pQUD7fhoNGPX+8ldAc0vN1FgAKAf4fAjVXiiqWE
8Q4hXYbnKHfLleQjZepGgsF6+hpvBOHm44e4R040YcyjEvFDvzuWFvuZdd5Rv4iP
Ifv6D5wFvDcdug+ZOa0hLU1H09fUJDZKYWQBnQXTNUGFm69tXJyjAIULb8i21vnT
FsaOce10TkuNVBhp8QR5mTNi/Y1zZctE8ok6mw8W08B8+EQEPaAKywnvGpS4FcH8
scl496SEQiepfmCepPaTHRd/lGTzV1TGVLQxKbOg91FKRVWPUbtzkBKSQvkzmsQ+
thekQwXQ10K3P4Jp9T9Yfz5Nm0l0bnq5W7MYpCusa4VWSBwFYpwaL7IPe6dsUZ42
D+kmATHug8E5L0ArUwbTcd5hPnxdLBjOZ7Ne/HmBA9Rx/esI6yT+uREB45a7tOim
xsP5rhmnLXfNA09aogZKGeaHX/WJGy1oOoomOATXtGijp/XKAdBJjXD/OtT9belj
NzgT+uCc0vuZHtjmeb0wrnLs6tBwIGLD5IZ0caZflJ8Rc2j6eTqRmkNU2anWQjRQ
gxnEryQ5DYqr+xq3rdtgwG6DxnoxIlBi8/t/NmDKeOHBz0Ld1qpgthXQjCZUsCur
MgOd/0jnZ+A2UTPhZqIASQxahWoCRTROqXThp2gmU/jsEZP1ySBp+9uw64umy16i
RpVL3v2eMxjsGdcV0m/qCLZgeyKtWt+mExi/fxiKfdcuNyFziHxzg3T022g0N817
xVx/5cJVr/GuGZBkgZQnyIM4DdoZsM/paUtvkh55pHT0wM/mkK336kha1FEh/T/R
fa43v6U6nahocCXGvr4A75OCm3Ly+384/pYnjh5C/PwA92AfJaRMs1dgP7JEydNy
F/xx9sApYTdyr7QxwrjBUx2OKedvzxskmil/uJS9ZkBcKG1KBrK+1GizUXcuxeM+
zUElsPDHA/8G+9ZquDBQlbnb4gWCGBRjZZMCmPA87WFyVk+PsfYfOwIncC226AYS
DvvfZ1ETVaMuO3+PJ16k+iwHnwkLEqPjizGPPt1I8xdevX1fq6xMZve4DqtIM2Gs
AW363Y5dkEnHFZKDYk1v6q2Nph2K43e8YeyHHmM27p1/L0h59eelJSpwLrRWWUf8
UEo+bJ2RsooSIPBlRYCk1ZJOA6XmE/U08F9uoJYRnEJlzsspjOldMjt/MaJN+2n5
bMzZhk3rqD0XkSo2rLX+Cr31reGy0kV+IIchL8Y7qJZ+MM7GwwpFIs5nzGqV7svD
TEUevu5crNQrS8UJOvHjFQ54UUDDQ9IGvHuQj65CLyxPRSeixAlTVnP0Abty321V
3eqBw2ko531Wt30SH6Wl5diRRZXk9758cdhXFoGqP12aTtBr7kN6w2wEB439pI9g
4BxPKENRN6wB4FMIk0bEGdl+42SU3nquKYAT+qMuGiLolwsE4dzk5hgcjkMlk+0u
Erf83uoVKQlEdB2LqRputw5/KTjFf6Hc4bBVd0UNgFnWkiK0vscZFRU4MD7kNYPf
KByerUkRN5g6QVf6E1j8sK2NFwBW31LgZZo7fPWlJqgegwmxayw3GD9kSjh2gjgo
zsUMBmVCDkou25IIompekpMiAqw/3QjKVyBp2ZlL4HCWGqOR38qbTc4WTpIs8oJ3
ulNOabOemeKGlGQpUKyVwk/LVg1L3kvvmsQVUPE+EQo3/tgrKrCpGsbiYE5MK6To
iPJGygH4BlpEYhDqj3agSyCHAB8UIaGs+vqeCxg/PYxzkAOwzunCwLaKeIcQv1qx
f5PR6UJPnVK6ZrZcBGg6qVhTefvnxgPNKplZSuxYDowZHQoRgSII2QSRVUtiVyAR
rtfep3fJyJ8sUW8cBADGwmuUiZwpoPzb2GG3D7eMcxyAalGfFI2Th7x2na2uAjf3
4RF+Ds0afr3hIF5RKyJdiEl8uQTwp3UwG07ry3UkA/W3ryUr/ZRfaUoaV4LwVMip
d27SrehFIJ2c5wCZA4P79V+wo8IUssT381O3RY3jzoKZhyAfTsLcW6JT/d6Bso35
I6NqN5aiW+wPc1mi+iHO6TnkSqLQkT/Z0DBuu3vjUbfxK1z0HvFRt7nXGPiXohMu
DlYJfYw6QEFq4G0s4TEA99g92S+xQbsxa1Hw2UQoLpcZT5XX39sNutdKdYRBcq39
lnxatm9EDQz6kTsUU0hMGG2rbbeK0vYManZPld5CoHvlcporAmj+Xv2wd4udQjT/
mR0MjNb8XnSWz4b62AN4L3r1ZxLM/1e4wuEBKNvlfVT0Z05XHtA/CAgC2RfAh9mN
77qLWc1I2jCvMuEU2KxZM5jIa7L0krltJ113LDHO1IYV8pwx4vnEE8eh9jrVHRdW
paZw/m+OOFZOMeW1skWTWmzf69i05AbdrLAuAmahOEM76Cgt6/h91j8YQP0+P077
4RA/8PYffdzkwFmh3c9WV1wMzEOzT+sm32wlH1Q5lD+WjeifBZLxSeBReotvKki5
eiru8y6vthMu/e9ukzRNjJ4oKloeHV3Ftwymgkpg2L5+3wAyfvSq8P7lAdKc/s5Z
vgV2sHCwCitdcXW3ueFDY5BPdXGqdFABed7ZUF9PTAN3BAlh2OnqLgs1kXCJqUPs
RXTCmX2rFHYuS5Gsqu7nT1vZqEH1Ygm5t8RHIa3Lx3ekj4GJgkoUZLJmf/pEGbUR
YKAbSUcIZOlqSNCQVvLV1LhpOkVm7EUnDm0PC+3edcOgcsVpFwMye+BFKjaejzfx
C7Sbf0jXYmzl9ifRCZ28XZwhNiWxqGkZO4Jy7ryAX6TIRy7RxRNmc8Yisw8Zjq+g
f9rXv3yny1g/Du2jx/9Pqx6YzyqR/zWTj7xll+WUEKI4pFmCjYFDcS1S4b4ANCJP
c0QHzBsx6off7RmuSOf5mMPwyd8mg6+nrTnWsVBltXeTS2gBkoehtQCjxIwIauJl
kXB9cJg+GIpWLPhap8lWK+8eBOnoLXnsszx84QPW5MjPypQRTDTpwV8ctAkP5fXl
Nf7Tnz47FRgntD8mOMJW4sdmSAem4UOruRi2ddzWNIOAqvdiqs/uiwxwj+/u5rJQ
eAq1CgmzJvG4vjrnkemxkJqzLqK2m85mL5WBaZ3f+HxGY1g66MYT5JStzuRovlaN
JTUhC76Ak93zOCf/FpXSXKCpOutNRLAIbd1HoREOk73FBR4f0jOnBc9Gq4t+bK3J
TfUVmOinmHX5FeQn6IiIM5PnZKS4SjSEyDcM4Fb4gvFYwEmuU1hYrcjIJ28mXS5U
VgMlD8E5ScZcRksl7xHzIPCQaaGEIMZyUMLaer2XEJywT69jqJFTwp03M6m1jmGr
NrwhLbMVRvywG7voIwkpCrVjPC+iG205SG7wt8KaHILOSpoCzQLR3IZc4vZhPXMu
eUd5SBAqtOkwaCFikR2hG/HPvLtrXFhRyFzkMtbk/SvApTXdGQHEXUrVqAU/vkfK
PcgtEe90iKGhWax4S1adwv0JmriFLMaxJBbk7JkQEuzGDPB84SJrso1ZZaXxuBti
5pci+UCfYWof8qucijdJq29bsPSc11FrpoxQBwHxxvLi74IUWgO0hot3WnjajA10
3L0dBeqC1Sf99KxzuM1kVFxUWDo5ZjiIDRdGUr5av9HpJ1NtABBREiILyAVNriIh
8MHtusO/DEeg6/3MGkdr1SmLACPly29Mv7Oj2oCYIKIxfTBNihfhC83PwgoGfzdM
IQm8XgPKx2wq4cUIxDU35Tm1aIsf1TeklZ/GfoH2zKDLM5hhRSSI1cDtLM7oyf9D
mOENowvCRAYcOl3WYe1ixqdvXxach31jve8vF738aLveDMblhc7nFZRPGHMLhpOK
xIBPGYTrFvcYNzO098Q6Q6z9uKz1TH4Om2Yfu/HKNAagmpPY4gWtbfMSL82EjFZ9
ZrC3Vc5lc3EKLgkMLVkqRPY4aBmU6k8GrSZTk+2aJ3Mez0UeLHhBpgl3OWOhPefc
9nP9eLmf9+t6LnXvcczaDDreG76mF9M4Og6r4v8Tzh9BVsAB3rZgQYVy5CUxVwNt
X0YeC0ArzvFCZLR5S7h46XQ2m/1Edi+ccN8UYt8SXokiFaM0hiPrm9TkeWE2YGaD
XGu5ZTk9og2m4XR8iAgS9Rvl4x+b5iT6VN7vInkhg5nJvzJ4v1JeyYC3oY1L+R10
RN6z/SDkIHd1Kgoy2df8M47rm1WsiZ9oivTJ3QRRb2eQEnk8kkFhJDMao+nRAIkb
48LUrgv6LSJb/om3GfJKnAq1Xk6u9i8ix2JrRzNGsTNIKJzpO7VpPwOcBIIWJENl
fmcdXUpPq/o7ECTNpYqt0zGIm+qSOLRYopBf4xvMOiiaoBd+BWP09k7DMPJHoX1G
b395NG7Fvfe+F4P9enRbraXCJCU/eOCcn+gCyFx8gMSis4fMKUkU7GnzImmDpdgZ
RyKOGDcpUemXtFuKangr4Zi08AuWYdS5TR9BAxuAMVCboNK77U6YehKd6QwnRzLw
5HSRwX7D3XSNPjWq/9dyPVzSjBenhg1cR3Pin453fhwdqfGrlr4gELUfK44iOoRu
cbOLepU6Grt0ZWhCW1YJ6iCw4oum0elZAqzlaac4CvdSzfrciWcivJZqaVBmRgAd
pIbshhcuotpPs6TLhlXFKYxgIjqMnjZPVnc/YWmnYJbmHDrlg9Gtn3RWa/qG2O5o
qYrph2lja2e2l8iU/7n+1wendQjtITGukJMeJpv4Okjer6P6VBu5sjo/QGckaPHu
Y8CEgu4p+gBk0pri5iLGKHN6xt4A9ZhW7rp0HUY+KsaufPSshGKqR4xocR7oT/EN
Jc4nOHMUa677PJAjGgXW721TbxHGwoaSq3L6rbLpfOLojiA0Dl2cI/WIBN72Koqu
X7CU6Molpa9tZDUy4SdoSgAgClGOEVQbYRoyTNje/jkzAIN/0vX+jnNE2Pp0G06i
ezFdYjW18hgsNW1twMUkCcbhBnCH5MjfcpdT2E3BY6KlFb4iifi7yPcwz0G5HDiz
hCfQx4H32cry5ZOkG1ufIzmudvgTIXG5kZ3J84gFVLbtibTcUOEFUKdvMbx3Z+q1
Qa/t2lwvJ5oljkGGxwPEGsOW0ykf9GvgNa4bobnXandFBKLwtuc0gxF2dcf0xOEb
4dg9uemG723D9K60obNCu2ng+k8H7x7H9kmFG1sRxrUrI9drhDyvtvCKvl8Z65Yb
7yL9OgxydHFaTF45SYtR+DijftEMqxmlq4RHlKu1Fj4V0BnhsnN3SK8rvkMiRARA
78iiXcSVwULWXX3MIaSgKjmoUAVSPSyTyerf8igNv2yKGeWY9cETXp6HKQJjp4IR
sibeuQ7HEAX9nBodXPVYrb45qp/rBF7lmIyJb6zDLUbFeZhXapCvWDnmJjI9aC5L
fA6ZNu2+RyDZ7gKK8ubqHxm5o3SXHt+Ph2gdHYNGl7uhFCETBtuA2Y+AbuAwbADT
oRVEgkM68GjMDZLELjgiOdGaBdiwMJZmuSgbIw5Mq9e0N3O8efehh9O/EfmjC/op
rZXouEqAqfOeRfcwT9contO/xbKZLLnXPTljxJr0+r5i1Noi9KJvUm5G/73XRHPE
6v7vxYeRhjYa0ZGH3Ygs3yDsvQvRgzrFjkVfpQAhBPXSnrxGkJATG3uMGZxv4vuC
ENG0jrgrvtA/e/MW7y7vBX6n13d3ggo+dOSP1xLud9RRxW+Ah28TC/z1UdYzVEh/
TmK6zN8nlXj+EezjkBFcmgWzYkfkhbEqcnlM+EYoyNp4eMwPmz/tU183lo7P1EbU
R8eIPosj8o5V6ZDUpPXi8cuDIbVcZskiBFpJy9/rNxgUxvkDNCEu9T94hpqqvzUX
u+FwtIHshTWKKm4hVJx6/RvHWiSmH46eUYVsviNdTnxmk+SPVRfiQABDEQSxlMBR
Vqq9PeRpQ0HCwmHNvH5st/tNaMN6B6B3mIxvCiTY+UTK0lEpWFiJhmgjmX87i842
R/xu9ly2sQ5M3AYBKGetg0TclzvCJKm2f5hEtcm8ds/7LucKIF3Qs1uiwncitEA8
mFh5ZMqLsMtz2tILV9OPCninCjViAegaYrfovZ+6jCk3jszxXrRwBzqlxGolJVjk
Ef38icG372pQQOVfUVaG478GtSweyNNnRvLrS/FzUIz+LCxiMUUjoOGe9hBnt02f
4T2ZM7bUdC4tgx+fVXdKYGZ5IeI5vLMlSmNYyjAv6fFYDIjNljz6oc5x2lUs81JH
H0fAnL8Ch2S2b4VfWIKtGjSBlLx9QSQec4q91eTgXkOXKAW7gv9K1nLwdJu5/mYU
KSKx12KQ1weIVHUllB8zgSmkTpFPeqa0//XcQYJVgVOHP3glJDaC4GJcMhQQF2+a
vYmmBsZd7QpFyg2st5d+E3lcH7Gt+wm4uIDQufLJ5D5z8K7qJG+K1E4bpZ3xqJ4z
6+Qr+UpHEuGDDVCBCqAxVwpQ4Y3jTTOv5P9mmE5F8K6nK/ICKylliGWeMRgLII+L
GO7kaMRTAFGzTRA9vZr8qLppo9u3WAqf9Bq+H3MXP+H2g8i9nOe8YXD0NfvLe6R1
p4eTa+Y7xu3+BeygELHiy9eS/wuBQ10Cp42jMyklkPC8TcD3q00Jz5N+24ffSwzd
pTg1FU+vxRlj6aaXnT7TfrAPThD3vgYblWgQ9zvVYlEb5MRmbzhmytYHIr+fRsLN
/Yh5FANIPEFkG5gLbvAsPIE19ZF2FaxCc7jgMyTHn35CVhoYcDHp2afgiYhKu/mm
4Zj78UGQQfa45gDQ/zQacMjFoXGBGE8qg7MxlUu7oVcfmaeepQiqKBKa4avyNvt0
11Vtj9fptb2Okg5I1qdzdno9wNmzj1Y+vw+qMgO2JhWV/fZdpTfXD/fvhhJQIYEH
RcI8Jfku8LVgapl5vOa1Zqm3CH/cYJ862f6wbWtRAbh+40ZBUKAFC7xXfv6lyPQw
y2V8wdB86b9yXnlWzpggTg9xW4JkfIVQn1CfvyMkBQ0vnV7c6m/61kpDpxFgxriA
w45TczHf+yfVgabPociVCVgQP5w9Nx9pAyfFXCLO3F1MtWIXfOI+Ph13/HeHsLys
lcG1xl9Vj+gvO2cffO/eJure785TSavd4Nxpq6xDVxyRxIHcUR+7W0Mvp9vaSAxP
Ad01JCWrpkE31J39NOEbY7zf2TIW2LjSaKQBh5cWHpi4Z9ZdwkMu3JovPcyT38d8
0SwMDIW2oL+t6iCnqw0TjcHKm+4NwYMdULzjYq/ruBGq3yTkBfLNFrtEycS0A597
EcokNhnKEeQR9d/mFdzAzXFVxNZpsItijedAfi2dapF7bDcWXBsR3q8W7cQzXGhF
09/1k1xsN+jYMc3CwnGh5ZdSK6Exhsg7y7HypDQI/uJttjCdFGBJfhu4iB21E6Y+
bxPzIvMsKciTchBCPiHjmwGvGM/4cAB/M+mscwiyVshlZNGajEiTsbLC/p3mem2Q
GNyn5xcVlEKdq5JE7oZimmQcxNA6H1Og77F0iz276x479Z4OBJrHp+AarcM17Raw
Tm2qVs69KL5o6APwWveJ07dTSXjbOxGCqLK77riMgB6ZZE7o6JTQH4JQQriNjaEd
RID0JAYWL5aAUi3A49/ZY3qExULn1qLSH3by8Oa21YHmq9W8G9aiadf1zvUVdXih
NhTq6AAl6FJ40HgMNX8RR8A5EWd3UHJ/HqZjTk/OCVFsLYpphhE+nyfvYyvmhTMh
LblVF4RG/bdn+ihFs5evZqERgcZJ4d8wL48YwO2ioIpeyBT2iKgWIRa4257kS5jb
oVhh7VfJEpIClXlpPvvlWwnD+khUZL7TvrSlDJOtZD/ipOEV1BjutLcgrcZlhsch
jz8N8tyrv/iuaBZu22D5ETVHQ/omU/0bm525ECdeNB628a//QgzdCDR6YDf6O4u1
QKvOwE1eN56yLiemQxnb5Le6Px8aqI3bes2EaWUapa5qgQ2Y+YiEF4pe/Dz3+kgn
lH2K7PXcUrJiWkVtRWZvF1p6fQz4FwqzmdsZm8/0E1kXMArtONW/nTfwvIcryCGV
mQkZSn0fIbiple8olBilgRR5I72wf8hqyhOy1OcJnNye8Ya3c+pjuZuwZPzZmJE0
r6Q/ZRvo3r4L4+AvOFr/s8TvizeHFO+PAV/QwGJRigtuZ7M8PA6giSssL+VMnVJn
14jNCX+UHhijT+tRZQnAYZPguXJO2Ll2aHiKvuyS7y8XgijkRGJ2UNrVD9rc8/19
oopwMUS7Q81+hFsyFN7n5EOY4qcHTEhYdOTnbQj+2W44BFpmBhx7dnFNCOln1y0T
FvJrsB0rOJYaYb6fqvfXvEiZWUp9vmHYqcPLPQzPlrWEuloLGc5ccRAFqPc/TGrT
bCgqWcQVyW9plasFAPpBU49baHf6P+7MJ94/rN5fbnP2INsUANbBk1grftPsvTPz
ahPAXw2emUH9Us29vZLLGc1scYE3nCeU+JE6HliN1pq9BXmn82jryFkqiuZEENgk
IT1JpPt/Xnn+ZvRoxOqEg/veFdgc7+aFG1RCGFdkP33BE48D38al4KNCenY7QMPc
RU56jVU3H3RjNEpq7FpXGDB0MFTvrAYCLb9PpJgn2cNWbv6qvl7KTeP/GGOwPK0W
2t/YGxyxDbfpdTjVFvPpzj92hKxR7+PreawdCJ4+LLEgzuNhWpHgSKvgUh2ZGum3
QF9eOctOK2DM+zJqW4spwmm5Iyb5ODgq0IS1tC/pjx5yoMD43/xh6AbFQFjcRVlF
QpdbiPjKLlUoWJoK9p1AYpSQrCJWKDcaisAYajuBwZadeJ79dsruLJbobCk7ao9r
5wtwNl5G2AhW2+3oiXgwp88mla8U3oabYAxoi7XEQC1pPtc/tMr4dU3rNEvponJ+
bqum3St/eV5JQk1dZVtqnJdvbkCRCZg7yOg+1bJOlTeznE0P2NmZ8pcDlY1g25rI
+laHAHJncOlNlBJ4GU8pZBli3PkmY4iKgOiLbbUWg3vYQEG8gC16APmk7ASuJmkm
vs9zIUpohYd7fyS+XqtD2A/wAdnypBvZ3mRYHS02huGBTJT3NMz047f4Yu9dNm8K
qkX+8Hw9xZzvwoITXJiutqQr7nuUHFq+xH6Mcgli1qVM5n5l9JVkQvAzCffOqkt8
i9zJ7bfLTAq78m3Tw5Q7mv9oBxBrxws+x6ou92qFuYk5Cmptt/erh/iorKjmhCA6
uj2q5pugJuVgFwySFvQJd/JRq1UDrsVWONPRmftzfraQNS+bKGFH1BM4r1R1LmHb
+oOzP055GyjKUEpFZGf8iRgPHQvIacYgAgUvWJrHlSpSq6gNJSmHWCO3cLeBnJLL
sVS1LzdA8+JKQmz4QJFXy9MO/LD886Gz+yfl9SNrp4xw8hBaF1icqCmxQ7QbYTB4
COycz2bGptGzbmbSA2x5EDqAaKf7lP4DwJcpHTL/khLV3kGMtgLssXVK9zxNwBpH
IX0fxc1i4Yebs9qe6g4LZyZKkFbwTwVOL6S5spXa18rzoCtSV9UssnzqLB8Ccw5s
xygTNgZk2VLY5rIAwBbcU18sWUPbb9GIkqCHHgcprQsTVVq3t1PuG7g2xSi8sI32
e7zT2eGn41ei2HQ1dNfOJ26F5+esnjxbM8pfu21RAwJoKSQniOQejNp1CWDaEov8
/nDVXEOw5vlIJPHfK1EdufN0nsmq1QPOA3mlY77g6nf25moeTWUD7ELL2Md32+Er
tbx/Mev8pMBZf865YtzkGzu+510ZIxjp6dh/2tVXoP5ZpIX9nLQHWHmfPUqCvKXV
sB6JM5RvxtbWdjuEOA+Byos7XxAcZcsvMaTUV6VfVzwfpqwwIrBDLE/xIK5lGkAU
bqj0wyH87nKR7n4NnD2QkWaFkq1rrPy4TUNBRcQqRrDSnQrNjpaxS4JoS5qNmp/Z
yLR9exiEEfE724r+fs20+0DgN0uJ+ytKuUXKaSldxvET3Mzqd7tvOyTkEf4LDi0F
rwvq8OWxBmJvjUJUcxEflgw85td2zrvlDaUhHNBbg8SYnh5WgDT83Qe5kzWdZEcO
zv4XdVYNV4yfUBopdX6BBX5A30qxac5AzJfaF660d6UTOy4u9qUrAcrmDRe7Ac+Z
HVl6sL2ikZ1KaXACVYa00oYC77zdBRNPjpPmoT98nnCkqpYTF4dM1ZH6QSj8bj/M
dolBBGLdJ4dvkvnXJbY5HFVcUWr5baT6Kzui1zfjl7xzdTghzrI9svBxkPS/sgGO
3EvDcMs7JslXry6pyvxEbnT+Yjt+DFCq3NvEBzkLZAiq6PdyV2Pgo/AvyrYlP7kF
CclhJmZARqtdtmM/JyqUa509kNv92q7ELsgE7fgQZOOGBmbGjNZmGiX+WwUDqbRx
vcvzZhW4pNAPwmgsMrj9OMSPPKmV33o0dS4njerPA2pRJau5H/03z86SCHnxfcN6
qUyBxoCOtE4yN1gtBjDQOXB/zDn2oGx1Ylv1oqkXi0jl8cfwvA7nohh3/tIEIOqG
KvzW3Gcx85NrDleOJfmECPvIU9BDfRuE4rHKN8klKfivO08Ztx1EmhISKWqzrlR2
UUN+ZtVHAQSRDsTTLQ2fxB5nOWHpPkLGZeg12Mk9LMByZwR2hza2FtPGwbm4eOZe
zXwPLx6oP3qfgBl0GAta29LZ+ccfpICrU98OQB3G9CgGEiARWuzJcpkQLOMCZrmg
HpoXtdQQEO2SeKTe87Jxg+0G6DDeXrcXfBGPinV2ctwcpH2j3m+lCeMhZ6NABRej
UtYA2pU4wx+GFkX1d/7Hiosx8kF28RLCFRSUQuD4C4IVy8Nf79Cvjce5VOhlRU6J
RjY2XO8PB1ipPnVoqu9IZXqvos417cm+kkYyMf4RWbeQAfhjwOb3uRUVPDCTY7ZH
CBXFW8d+0eEcuMw71mhGnA6vg3FQMUyjjcHGFMAvUQQceZjbBDbn8ayoPzJY1UtL
y9nxGKl/0tO3PEypreLAMQp67zy3Ooa8Ha+yU81hXjHosud4//kw1jTQbo6eDSGJ
LfqR6M/7dakBiyKiWPLjIja8UGEugk2eEHMwEG4VVv98ZnKGDo4uvk/p7f6Qp+x+
FsTlonruQ7lyoHhCtAzHvzBQ9KHDyHZrsoIT/MnohuumdVZSCyryQl3G2bPOvhc9
ahuJ5GebltnGOaxorHtKbaaAWgkss3cHzRY+y1qUEh7R84Q6ndpimVtArhE3fMYo
flTHuYlDHdDLBp//DDFcta/ifcRlN6R8tVkzwgWfkar5+7omUOCg/5VPJ5gqa2d6
DtIlwMXAYWJAKM88euklpA0eRrsCMx/Yj04tw/odYEneqZYvQzyeoEu0QJlHfwOD
szUzY3+UYX0sHz6TZnmA6Dyl6+oO3v3ov+o046i3bcO97Gzkf4BuOnr6xmhwRKwE
7rhLCYQCRN7UGTbs0Uc+b/icfRjZeCQzEBg6sSEFrf9nwbTI2U8B6QXGIzczIRCx
MBi4W6HSQXXdBrJGwA9IawYBpfZaIM1INuszmnpJrksi2mj1a9EUJp/lBMh6Xfgk
Y+beJbSNPGZ3z1DYKzv+ytKKz1hoOLIMQ+vLifNjB5R2KXatLimAzKD8D7lSb7nG
Fiqa8Eii8+26mFWGEgwn45pepCq/gmjBXQ1itlrauNkf7M0jHFazRaFfm02jXubj
xx0CbnUE6OlbttUKp7BS7hItt7udUr0Ib23e+onipbFg5RnI0tFXHbIETWWESCxz
FTPIpOJvjcMBSs3aojgkKDm9FHNtqwpo48ITDll2YMLByyLFRDjgJdAeQmmzgUGj
UEvz3e453hvt1TI7yyJQLQ2Af3uSh8UAIezQ9uMc+KAgNfQYkmJTeqg8OquAGSaH
yZth18iCUTPo3ppTOq+GlYO7QYjQITkX8gwGyhY5aQXmXOLzE02n0WzkCPc2COuT
7LL6esKYbC0XdXwttJUqeda0TNGAW1+erCRucXAstvGk0QYCXhDbnjIZTvxtLmEs
apMICoi97IyCdPIuaweGApu/2wQP3st70HHnQFyDYSAH69LLQOxOVtVVvepQ58XI
cvrPZECg+9MwiAjJYZR0gj6EeBS1aQyoWAYDOgmnZ+HVw8pICRCWQd75vu4vKQi4
OWd3WoD+XS96WOV6U8ePhbycQgUQUg0bVe7jVjexF0PC5p6KwXc1yVn1CF1Okhbp
Wr6alq4jGy0sMig8S924XIbUPIyU5gENrJLQNMXh/MrtLBydtZoeEqjx39X8CY2d
3sYY8bbBLoq3htUCvTgU0PDeYvQ+yozdHHVKBjUUctJWXMCw2qwCbAQAGcaGe22J
JFmIuGvXAGecVqR+Pbc3l86bNJ6cEb60tg/agC/q7+YgJTRFzY07O5urQk0nc9KC
6ZDjNsOvA/E9PM//tolXd9QpVJBAM4MpQ8k+9ynWHQvaHpe/FVtHifhOm7s2uqGM
L58F7ctiOnF8iTBCXRZQOK2eyw1RFzFTBML/6LhfvBtz7yfw18DH3L1wekohOK97
6SCC5PwGzrxXvPYhe3pbovvx/5X3FQJiGBa3K8YH24gbfbM7XuKpjKoAVCdbKPXr
qfacB4jKKB9w91SfKOcgVlxY2dsw8R1v6gPzcD9W3YeHpA0QH92s7lAdUYGd8dou
E+jJemh7l4FUTE/gvnvd7lcfJzNVkGBSa1aLDDPPzbheawmh4z20B7K8Q3FwCISd
As+efbfMANo1tIuMf6xxcglawtWSbF8B95RcfLHCNnPPgqmtRxRCDRpVic7LSyiN
eIywCrnqtB+IJVnGHcDTYf5OVPSbW6Z8GzPknBpxwOrdedO2DgnJXxWcxi6pGUTr
IlDJl0Dw6PLDbDji/MmEpXSQZ05nETWcmsIbA2cLu8x+YbqpHt2mqUSnkDH5DS7U
ruizJpPbqbpRpA6OwUPSLQIKSjZb4yyioWzD4P2Rsi4CmHPo33HiKe06hibzyNmE
acg5ezbQkngrm09NmU+HvvCRdIyLmbgJcGwD0CTEkS0ZJuI+uwPHPPRIEE4nuU5x
A60NS5zuhbm4nEA3liakNx+Qo73UP3FNQ/WSIi7kdinGfg+3uxLLzF0wISUueUDk
pMTiCSoTgwSZgvNS+Z5efEVMD9qBo7rr5obPfejesJ5kUZDkXq56ySIQVxSdSjhs
8MWIPOIVkfHrnvVP8TxI30LHcX73MEgKkQcwcdHOtyEvAiKn2GPjXt8z8XBK8Dl6
6xt/XPci8d8uTswtI1BHbmktWpp+f7BSQAkCsVI/LytM92bgGFE+BHjXEzUTegdo
rNjpSaBX+AeQhhv24bEcJTMg0CBhWFLiGjgReoGI4VCrycMHMTTolhGjpFL+Phz8
TcwS4mNVZpdSuXV2xodLMBkWi9ofb/+z1nXQemJpAuHyT3ZJGAA+QlVm/9tYX77N
NTkgh0jf0pSgUGKQJkPw9xVQETYKDc0idJq6nAzYO94BEYMCUUd6MJfg3+sBSHti
6ftRsctuRk/S1aQxnFT39MVjYDYbVq5C1i+f5uYitAuPpHjGV9sKhwmCDwRTWMyN
LXvQQCIqiiWHPx2aliIhJ7gZPZyYN78/2QS3Mng7Z5LKasZsl+qAQehi4iFwmV9y
GxidPfYNK0c+aQFhk1AST1ODyJ8bNMa13px1bdeB8zU+zc9+gt0LGExaBvI6BUT6
8SzY+btZ3OeecYwnYZeGcwPedAZl7O5tgc0E8sTg087trqljD9KAXLB30Fgwfc+o
NT3RTuab9d4S2BTfqo1NgXj5h0iciUv+5qxXP6E1tduZwcT6AQxNefbLP5hQFOMZ
RJNrWan61352uQnE0kcSdMX/2SWOfuuNEe67ATMO4f/IyyJsEkW4VjLpSzHWpK2L
NstTygXMQ6ywV5PkdAWztXrAGMpiQiXrcNJyaNQM6VC7pQKqABQRWdrMpRplJkto
8IYlpbNiEES0r3l7jAQ5PKUhiGoG7j554QnZTh3c9ftkcdIQC1fOnc2puthfMZUy
dyooLYc29eJRnWHvMEpH9IojMIhCa4hRzw7UUyxBc0Id92Ninqif2X8NU32JslY+
pXnpxLoJ4kkSzZ65UYyt6UeZexOyV+FtNKB4+o4a/ux8hhdXjpZNsAZD+/bnQ3jP
ZIZ2haZllhBYl7nDgxyY/1y7ivBbAnUcAoxuz1PhF1UH0YoMChZtJzzHuhb4u1/8
RgcBJgyKB9V2U+m0xUCJ9GTU4Q9HQ4OB+2yZh9QkFuGqEZoow6Ohcy3z2Zh87kJN
t5Qqga6TWwJdFZj/ysH9AIcDjN/7VaCC8ls0mlIWQyBt8P3dyFxhiADbSVs0CPT0
G4wZ9lBdpqU0JW8hpid3Rki2qIXkowBey9Zxa3ODMvsmKp1QJGXgDw0Iyq/goLRb
WLbVzgVJkJikUsKGH9QAPiRy0jqSJJ8SfI9c+lG4lEdgqZv4CttlStEvUMcu/RnS
i38q3vSJGceV22r0ARw4qVZB3czPKyWLZEnI3uL6o4nNMdiACiAT0HAFeNZxkJ0a
TCRN/FQtv5N7bXpYTlL3VHvPeQb0vrOJNkzQMNjJq0DoTcFZOVZYALVWwAjxQzUn
pHqSPxDtRYBWQxFJu9P904EA8Yg/uXRZ0QHncf2M/9cE4mslfFiyCwczatJqspWe
QHf+2B4xPOGoNnzskO0WwkZCr9ZssTCQNJFVeuqbnWpOoFRNpl8aup2EsssSitJk
hPDJj4he9Re5udG3w3oQ/e4Tn8moghR26czhC2G8i2iNEobmgz9r/N8INzPUDbUt
r1OVkRDEBW7Cw1k8ugYfc6XETQ8MA2XYK3KG9d7H+qWRY/2H35zVkX99Jt3w2g1J
PDgXLxMPel50SE4fJ9U6WFW7SZ7atdHgF/ViB67hjci2BT4II0tjjIGfAUcS5u6b
cYqyK5BJox3qbcTUUd9BsLwIdZafJ7l/OFekTfgnDBEB4QvWGAQb8XDLjQAMKeCn
Quq5Ni1F/4I5FWsyu9QuWYqVEGu/ci/RMQBHLwYnZDCbJ1ghYx/aF+XgIjkK2CSx
htoJcP5xSEBGcRiDZwY0aeuLg34Oapo66guMDhQuG61VFmWS38x8oWcobyuCgx0k
QZ62aTQkl+xs8hqHvy2RK+i1bhD6PdBFRkkKw8j5xW4RlKAQ2lmepGepZbQNPrXk
oYrgVPWkk2+RAdpI84ull5uJB9RzBE4nPKFlwoTZp0D+iSd3EJ6bjPq4LFhmzK5H
BayFEHML78g0OvIuYtXGSRXdoJsFJpw1PdRsdOxUMD+f7gzvUMAoLEHyFyFVTZow
y6nG12wxjJ0KPy/JH9sshsEnRK9YH00vI2uUuQRNWoDbpGSoTHw/y3zcNP23EXsE
MgLsiCSUHtGMKuCOdqQcmf2C/KnZL5wfLmEkcbOZoDy/pG/r/ZMxljvcOdddCU36
YW7oz4zDbwHU2FDiJJmyQAckiv3mfuL3glo/t7BOMPJW1L0IcHHQNEKoCyc05dXW
lpa6+n2cU/NVr9/q6IOjnnSEodnjEWpFH9axNrIu9XqMjK+lXJfd8lteEk4/q7LD
0YMu1MXZEwtJRQITP3pzCUeDl2ZDSP774xQUAh5UWqNrqkmFdcoXObVHLmXI4etU
eJJhKRKiujFCUMkNz7R4zWUWa/zV1VeF59fzI8RnOPAFbCD0dLq90vLJAUHVl1em
idQmf0blJGWVgB0OPoiA5/wSOIf516xp6t4aokgyb8bSp0H7xchDnPGM9I3mqi2X
z0/UyLhq7H1ICC6jStQ3wGNbe9KAiVqv+HcOrYdRHFMC9nsY6WAbQInrW6bLgLlo
SBQIDi7r6PtI60yF4gn4XXVnCCcpwlnVbUyDYeuyFc6tNOvlcYnsYOAIfgg43rLg
bttmVQY8OJNgHqMsOeCFGmc65lwOzhiYDy8PVJX8MEhYL5U3OHGtlvYhUdl166zp
th33988v4BZYo60uJXFKz0EYhp2ZtDkqw/Sp9DU+EasWs4NnbjvQvv308LYBiStw
o9Bf9SM2PtbYcIt7/J8HZyE1mwwUw35dvieJ8SSN5npNHp6+uDkJGPSX49ZIggQF
t8X4bBtN+HKG0smNZjEWiZ5ohkx7yltEgVe3e/2DGY3Pvowddd/c71YxoY7dVX9o
z2HEADZBxWsnQkWyJAM13xbjlK6hJEVuR/TABhRjI8GNRISYsBOH32AjobgfRLh5
pLKJWPHwR3HPhia1JV+3ZJFJBi2kPNTrbPg1O34cj8hs5o+zu7BI6m9Fj6jPVd8y
fJQC4taiwj7H1lvKNDMgZjw23IVaz8SEJpqPv/Sqnd0mGIWGSStWPOadS0ZXeGtn
NeCC3j0JCqzNfr9UdzT35gVbGYh4PV3CmSlBQR0RWc6kDNsFZIE6dOJiANSyhKu+
xSQYi0XlpAGvOhi4CbaP8NwSf8L/xUmkSBdCvNGVH0VFx+Cczg45gQvQC6Fr5Vun
ZaJonpGo5WgcooE7+2uP2IJp0dFwW7uYE0GAL6PkvGPx/+wqw66ggMPGcTwebtUS
84GT8RFDfGzHqIbv2Gdn6gIXII3mX0r8QQVZqDD7RB+lAQrF/McYuinsUZQoInKY
g05vwZz6s4O9fn6rC+i9llV4D1zZtAdzt1qR/x6qtQK4C+E1Y/7e5cCc9+9M9DqL
aeFPibmZWGZdEs0tWb61TDjQMFWzPzo7e71oGyh6UqXeLaUS/Zy27rf5t7qT9+Ms
/ncpUhOIiOQ/y98E/TZQ+3Wx/ksTrdq7ZCe4+Dav8pYMUfTqu6UAc3jRZARtbci7
U08ZdzhUXkXCvzU4MIlQK3MoiH/ZOelzcJvA4s56HMvqRylQI/DS29/Sr/a4Btgk
a0I0MBKWKx1hmIVAIjTLSR7jtE+iuRDn9G3jFWkRdOc1kZnRXKAM28pCSpGb5/nn
WRKv5PlbIUHbktK8nC1O/fmuMKKFIIjO+9stxdWp9YwXTBuhHvdED1Zu2yucRe4D
rHegWMoDvLsGS5BEqUUcligt22NQ+VLIwUZdLwr0O51DAm+zZKPbd+RBSiciwB9/
hzhWNyP5pSWGTYcjhm0+9j+0Gb/trlGmumEoMIFH/lFdSPs1fWhMliL/VVFlqxKc
aZ20Zd8rRfSF58tIDDIhOdM7mWlBVJVmzagbReI1vcKhnpjA/XZFAHF8KXwQYfa8
C6btaaKyEKAHapj/5tXzv+qzexRdeUDoBon0l5FzsV6/HM9iwPAGTBFOA5xEDBgr
K8XYpydp7ytZjxnNhLEQp1LrMjCNrqzhl5h5xQ/E35/V140BGaxNnWioGawX1MdB
DdVEOyWQ8xT0dKZPj3kHlp9wxEK1bivSsioEMt57tqevpt14LOcZeEC+cP0XJCbU
Q5qTOz2XLIK/oldE2psX9XH4F64a4Ksnzksz5HCWxDDIdz8ozEQkMra03weRsK/K
OK9x1zwrCqKSQ48a+IDj2iG/6NLSmcNaUsqvi04SsW+fsMPIKbm5pOfFrvNElxbp
OGw//55xMwXZqogAMIovPf9lHzrytOKalIx4ERZZ6So0TaVFaSHS6U7Gk5tJUZGT
eYr5VHnhkxqcY4hyP0DaHm5bgparInAujKkKDACgYcGuVRc0n9znCsEvvso5GB4D
FEZGF9ZbyJHCceegqh9C1RdxZlD7JrXpKHAupsGvRSgUZ7FgO1hr0G6PRWa+e/AD
lu1XT1aDJDMDR9BGWd093H0+yWJiL7pYtsEpbEYLCvP5pI0pV/GoOs69BGsnbq1x
qorlIDJLrbY1EHzjp7Dhs9bc8P8sGWv6N7P2gPIcWp7V9dM9XGxQk9XKBXZbKYQf
nViutBF8sJHuRwquET9o1I4Ng3LUkH0fPSF7ZeKAoIswtrfItQhZjN+YcYoYG4wa
pB31JetxbxOm4MOGmyKB07AXsc20EPc1+K02/hHAotBZcA1SBMdUMUJdsO6UW8+n
9cKMkUsYEEfu1pV87+cEZbLIuuVB2QcXWHG+R20xYpRAA92v6YGBuV2FoTeUdx9e
Ev7TLooiwc1YgyxHjvM6nt8KZbGkqvP1QbApwJO4X9zS+mYwWxgQnh/97D2rhAwR
7V/9e479hKmsOc8Cm+Mi7xcoWEXmXTAP2DeUghHIHNhc5nH/SirqMYAWGjV9a7JI
+Rw4qoiGHtX0Cse/lK1qBI0IL2WRgISJeNoQghvYl8yRUJJKN2n/CfwIwkXjV3BP
VRKnOdgQyFAGR+JCgMY1g+TbboiuwK5IJ1Wu8+mZjWfZKUPnPYvKhOY07HK+EdNf
MnfWv2lGYgb6lbTOWa5BHnEg7JXIPKlOS2Ak+S2H+cxG3nmeCnINIFUuL6xGDBzy
0LTAJxsZ9z2o6hwJWUg+4ObQvwJiJ5TaLN+pfCDketu0+z5fnZky4QcfzdE9hs8B
8MFFakHDda8lWJ2wEjNDi64qy2ZQmEfaBvW6fi5n8EMxGUylAaTV9/qUfnZucbgz
FHlr8Oua0UHMo/AY4IPKB2nOkldNha09PNH0L8uOvoRDAT26cYLozv0ktnwD5sQR
066SpTZriUhFyPq3GS30lLR8fVy3Y7FpJ3PVMVHwsLC8LGpJdLKrZZ12aoU7j7ki
0xcQXxrkbwb2LvI9xsw5WNpnBwQbSwxdac/edDhiynUrV10+4HzuZa/mG11t7T25
gtkWKjJxyDCRw+IwVH8RZIIwyWSKdK1LAjACCWSA9PkrWaM87ADNX9PC2nbP7BUc
2gNXd5hfQ+OuvcMUVpxvoGuV5wwzrtMbfCEjhSGdpgCNTKBYmc0lBHksqJWoQOkY
aTYLryIPSbcFtycqOGP/ArSSbFsHDIxGLDP6AwbgViSNR6rN72wRQnn52JilQvyl
hA1S+FAp5OrC6aSp41W70TV72v8R5GyKvR5rQK3EtJGnAhXFfxTZjZoHj7tTf5WH
RuK6vN4Va1yZdLJxDy52JcE6ryAeyrfMv7RqLe5gs/SZe84878R5J5lvSdBW/FSX
G/Lud14NMnAljXtY6nQG0JBsnP6HrbUEFRSy4SzL9ofUQBFhpnexo/lW8xWSJ09E
LX4ncExYCtdCAH3Lv6a4cq9qDmuyfviPl+HJ0DB7q8gYAsaybKYdrkFOLsQLnDdl
su7Yn9nlLqy308BjTxYuc7R3R3tcOF0rIaGOhj8bf0sZ6OwHz5iQ8r5WQWO6G0db
mjZM/WRdoDiPO57ZSvK0RuTPIAUD6eo9CUYqPAfaCvxxdFqxdBBDxNyQXvf/+xAb
AQjpyxClU8WmfyPEv0TPq+Qjkkgh+QHpO2XJEkWIv/+CLVcQ8qVgURvOaT4SWdZN
eKibXkJmT3wjiZ+1RtXGQCjYdPYcSer/hMU9JYxdS3jntTHrjKEClj6v4dBnNvPG
EYmScYPZsiki8w0YHAAwxi6euCPT2fUVOtCQXnAsSXP71my4TD966+JCkQUYjgVX
CSBhRMOwOsi4W1cf9aCUyMYjPe7O0roYRIGTmveU/Xnwkg1qpt77CsSbibXwgtrW
BmsKqo3aGzi9hQ736yLsD+QY8nDMDRVqbNgV64+Yg78XNV+u3Qllq/jGCU9V57eV
HhxVJy9zG5+6SV8HoMDaTlrLqZECaSc4QzlTAhlnz6KLNlyk3layEKa0IGKD1Wgl
FmfUhybXXrca2mhCEDI+0iihqHTP1/N2HlgZs0pKfOB+bRBIZG7wTyf2iEIc5tyC
NVHUdI0kWsjClG04ppclaRi62BuFWQxzpdPx+XoCfwxn2JvnKCJkgNvRI9W/BCXe
mNp5bvX2by8UYcdtWLH1nu3jry639Toejlb5pnZIYYdNKz/tx414Kfpk2Lrzc6nu
xruK6nSx9IbrojJoYs1YFoifzIX4w7857eqKqDOUUJwHYT81B1MGyFNmywu+kJwz
VHmbGphDrrwXJdSUQ9uwUs6s/KCeAF5UPC0/OY657vid6q4dHKQh4GPfXdj2IB3I
6F8ehqDE73IMs44j8QvOqE0Re2vLbMZe4U2AHyolWldB2PLV8rPXyeg/oXrTpaOs
6EobzE+X/2MHt6SJotFCumrqgObq7dNd6cu8Oiszor1vIQQO3vuwTovf+7OuRLgL
mahqkdAzx8hl9JEV5DxrXHhlbWGIbjDko9H1G29q99bpWJ69Ta9DhlJY+jqzVuT5
iYiaP2snO3O2EGTB7i/JtjLIMUrxpDVaiCulTP98WE8KWyMA+1Pj4U31kpuWeGV7
0uMYh6XK6/M/RwHjrjka6Xlb2oiyhC/MOEJbArmDqSm/FpKtdiOyk0c+YN1VtIp7
5vSPTHOV0SbFpCzSj5t+giZfCQ9fZj1jg/sz+mCjeJtcqTO++a/mCIaNTKs/M7/Q
+PQogDfCva3wK5tDa4jkKE8bLKASRfWcoPj4T7Ds0lpaukGxMiYgZEmNfkvEtW85
4uOPCMWU8I9/lLoVjYnGPTH/g1jCu63Ff4UbIJ5yZA9ckc+ZOEyKa9GGEB2Nz6yJ
N0Ydv2FFwJozB09YS7v/5MNywAI57hPje4G6CBuL0I9QaOCKszFbzxWViW3lPcP+
StmFQMZCUgggy2KVtLuLBwHtxCPcMrlkzUV6qRj0oyBU4xTzeYT01Z/luJSlJ2CR
IWXG0P87cX6ewaQX9+065TxTz0zvN+mwYPhELjSPPsItvtD4r2kEGvq0SZIr+5Mn
7Dgg0V1MjoGa/tJ3V5ZV72uf2lCqdp8PJW+ZaXfqLEo/6x5g9lHWsV7ie3ZLMe/N
Iaonha7JNxUG5OgZRcRFo/DEXVQ/5s+xPfQ82EuY7x0zjIrqei4jVEomR5lQgnmY
grXJ1syTtt9I43MizaQV2JPp2s8x7Na0Yes3f6arWkU7BrJUvIGMvE7K68c0pWZm
sRLGB+x0crAtI6f+wD84QIz9UviNafewaVeRK5NyeuO1r99i29ijZdH3qqCe/FFE
65Fl5ccRoHV3bDvv0eVoumEfh3IfjAy9zvkOlLK0AMMgSEgr8Bwyr/qk+MfVZhqz
KhMMrOZq8Jms3DBwuiml6bFIwSmqOgwVAXGmy9IPP6etu39oeoqF93ItyW/JYdy/
QwwdjjDYLN4RvpA9B0NNOl+96T3DOjo/955o2TBc6C4uicfALIQLvrJcB1ZQlEOV
hm6j8sfmy2Gt5VvBKRZePue0UWjYTCnnUEzyp5ynQdT1eUJGmilNQNTvBg0S5Jag
ZXROmY/5wlqc9hgawbIQ8ccHsevcDW5xqTA8B51RD2c3pgoLtol55udQt8i0Z3No
y9pA9UMql6X5LvZ4ZW0pjNuR/omrJCYGi/Mm5HraWS+r1iPKlJ63GT37m+VwtamU
mlsLHnac8Blq8znpzVoBFbMQ1uE2LOMiM2gfOO39K9eVho56nf57jjlTRAasFlH5
pSlhLDIRBPx3q4xfAKACSNR0b/HhlhmM9g+ubPvB+jBixr9pFjL9ivHorgPNoXLY
tsP6KmdWYjlJbLSPrkKyEHH2ar24zMB3Sasxuet7LNyQ2B36MBCOSRo0JHtRh5Nx
h6YysKE+LYLK5Dlj88izk+QZcDZBBDECZ8t/jyAFQnFeUaiiz4evGC3Q2Z2j/pib
ywuq3fzpo6M1L71Ez4Kfr2i4z6RYjW+adWT4+kxOh6AYzB4UrrN82hwMIGwSU6Z9
uIuXsXwvRXSqTrLx/xh/HjaQadAigTAnAE46jCA8IsL5pVSpDsKF9DuWgZyXG09p
VuV8TRX/mm3xufIXtfEkj2E0nVPvpqqQBsjNJsnt16H3jvfim9rRp9NmukYzt/wU
3Uv3wM6Wqeo0O9+eRoyBzJdaXTive6Qv0ZAJRROchlqgq+TRBwHYKXJSCCPQH5Zt
hEOnJKqwliEhTiVJIhWAcSokq+wRekK6JkAc1GF1rTQQ9vAB6BxiOTeNGtIr4i9m
gD6hK6mi1ualU+k7+msvDWHxueW8g2bt2LI8Z0jZ7U6L0dti8hFCXWgGEndXfbrE
3VzmGE+lmmml4pny22CNY5GJcrDBn+MvF6yIba62yxkj6elocpScKF6auKhUn1Oz
IsitvirwtGX8+a+7kXIYqaSjFFuWJM9zCDMFUVojw56jx8DTL+BZ47bawFnRFP3L
GIQnXxsoQX/Ohyc2aCUuF14weTG/NU8JQGxlTCKUjnyAJzavpNyO9IAhXxtz+tg1
4IfoSeq2fjddSVfgTFts8pStzT9Cu3crJv/n2nrp8kwElk0S2bvrm6OJu2JxFU4V
BIOpnLe0drTg0uHt0wPS2EtlNPujvUbdAWYDpPs7/059Oq91Y1STcySHRI+GtSWv
AdU2gaMDPl1+zseesFN3H7D3S1Mn1E6tirfxP5L6rlXulaMh2qNMFYz6RH11N+R6
PxLWZk3+LnaqZgD5RBcaWPbNHjuW9OepmAE8ZlBE6GKVctseOyNVj/BStwnd6m2S
XlWCxzPnVUd+QE8K8COWmSv91byQRqcW3CMrv/MYnvoGry1oAoFPSEzIYwalv3tV
60LH63P1aQdxPf/uYMhpS8n69enC83H3sqVIv28CVqO+mPsv5YAaxcMtZS0NGemK
Ebl/doaqgCSHSXhg1RgBLLRUARawoJvT03fGzb/bcvFKhYWBE+jt2ihbiFceJudR
G7jemj4mnCFLrgft8hEnNVs4m0VIYrzJzd2aCcukKxERsFLLxhN6I7GfbzkOpt6f
qQbzyBx47tdeA0FTYL8Zx6drtCcWM9vx1IRAMS79KeqWHPR5NKmEROlFs5pEfhhL
m8BBXMcvzJGzW5j8Cr4qLxv9HfbJSqI06AWBzhVTnZt+17o2cyB4nisCuIu+AC73
AA6al/45iNHtPDwDsgdO8ba+cd/tAKAEjpEZxtZ6To4J1wxrj8jG7UvCHw9vm77U
jXFa20VVL43O/uprQVUdxwTykChA8/6cZCIqMh/ir0hj5VpDCjineknL4puyjIiv
QgulziGZBJePxzwp2WXP81YlFxML974T8AT475qTomOHfDnfQK23ioUsPVR2dpAM
KfZOTvdz4vaqe0gR8lYsWxwckhCHTgbbZEkmrUeoJImsx+6tY/gDUqkU/0ZOuQOq
Qwf5fslQ434qWE+UXZkq+7x/J8GTr38qS1ap+MtUJNackJC/2LFXCDLSR2ByzR93
IzHttsW+wYnw1vtY2hqsZrTsq52MuMkOOdRFADjkyU4TZXV8MS0Hq5NHlPmwOuA4
QQFPK1N/toMIGuhHM6KbkoC3plgjpXViZfPQVkdbSf9ECRB7vM2ryDzO+5QYenFj
h9UkzFQ02oD44mOZyD272eP6jFRNZatOIn8vXYlOD13Kxoy09k4b+emjBZ/5tYqs
pWyIdUuEuMFqNml6MCq9pdR1nRxVO1MY3HSVxVB05oC/4dWhFYcT08++GIORKXu4
HyW3XypjrHAmHn6/ixNbKtBzlxH6PC4y06QwzWfyeb5uspghE+AN3xqG5Q9fg/3d
iRg9HWxdlCuAhdCyh5qCBfv8OMRGPOSxrHKvOFWfXaQMdqAWFrY/wB2xlxrhLJSb
94r3JUDsiCY4qTj15Gg+QYe/5+cVzSVBUWxyzTsLu5CJVYBe7r8ljonT1RdnHKb+
ylEM5V3q34bAdfY1fwi8Lre5qfmVBuQa6vl6aXmC5Ms0FGp6rjxGeUVg1FqWQkv/
jOaVDJMnMihI7S45hdjMHgGvvdRq5U7pUy6w6gRpnebKYkpHUV4wcjG9xHcLBkhT
wOaytx6o4l/Dyq5ZdKMpBMmrt+hr9ny/9pL44Ss1UcIwtUHrmtJ29Q3x7OHMT5QR
eh4oHARMObnxYnK8xu6ePw==
//pragma protect end_data_block
//pragma protect digest_block
SdAZv0iKSmVXuuVg2dponvgi6fg=
//pragma protect end_digest_block
//pragma protect end_protected
`endif
`endif // GUARD_SVT_AXI_TRANSACTION_EXCEPTION_LIST_SV
