
`ifndef GUARD_SVT_AHB_MASTER_COMMON_SV
`define GUARD_SVT_AHB_MASTER_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_ahb_defines.svi"

/** @cond PRIVATE */
typedef class svt_ahb_master_monitor;
typedef class svt_ahb_master;  

`define SVT_AHB_MASTER_COMMON_SETUP_REBUILD_XACT(curr_xact,resp_type) \
if ((rebuild_tracking_xact == null) && \
    (monitor_mp.ahb_monitor_cb.hresp == resp_type)) begin \
  svt_ahb_master_transaction new_xact = new(); \
  rebuild_tracking_xact = curr_xact; \
`ifdef SVT_VMM_TECHNOLOGY \
  curr_xact.copy(new_xact); \
`else \
  new_xact.copy(curr_xact); \
`endif \
  new_xact.cfg = curr_xact.cfg; \
  rebuild_tracking_xact.is_trace_enabled = 1; \
  curr_xact = new_xact; \
end

class svt_ahb_master_common#(type MONITOR_MP = virtual svt_ahb_master_if.svt_ahb_monitor_modport,
                             type DEBUG_MP = virtual svt_ahb_master_if.svt_ahb_debug_modport)
  extends svt_ahb_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  svt_ahb_master_monitor master_monitor;
  
  /** Analysis port makes observed tranactions available to the user */
  // Shifted this from base common to master common parameterized with master monitor, master transaction.
  // For UVM, it is available in the base class ahb_common.
`ifdef SVT_VMM_TECHNOLOGY
  vmm_tlm_analysis_port#(svt_ahb_master_monitor, svt_ahb_master_transaction) item_observed_port;
`endif

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Monitor VIP modport */
  protected MONITOR_MP monitor_mp;

  /** Debug VIP modport */
  protected DEBUG_MP debug_mp;

  /** Reference to the system configuration */
  protected svt_ahb_master_configuration cfg;

  /** Reference to the address phase active transaction */
  protected svt_ahb_master_transaction active_addr_phase_xact;

  /** Reference to the data phase active transaction */
  protected svt_ahb_master_transaction active_data_phase_xact;

  /** Reference to the current active split/retry/rebuild on error/ebt due to loss of grant transaction */
  protected svt_ahb_master_transaction rebuild_tracking_xact;

  /** Drive data process used for handshaking between phases  */
  protected process sample_common_proc;

  /**
   * Flag that is set during the first cycle of an error response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_error_resp;

   /**
   * Flag that is set during the first cycle of a RETRY response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_retry_resp;

  /**
   * Flag that is set during the first cycle of a SPLIT response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_split_resp;

  /**
   * Flag that is set during the first cycle of a XFAIL response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_xfail_resp;

  /**
   * Used as a flag to initiate the zero cycle OKAY response.  The value of the string
   * represents the cause for the zero cycle OKAY check to be initiated.
   */
  protected string check_zero_cycle_okay = "";
  
  /**
   * Flag indicating if a rebuild using SINGLE is pending.
   */
   bit has_rebuild_single = 0;

  /**
   * Flag indicating not to call the transaction ended callback.
   */
   bit drop_xact;
 
  /**
   * Enum which indicates the location of beat address with respect to WRAP
   * boundary.
   */
  protected svt_ahb_transaction::beat_addr_wrt_wrap_boundary_enum beat_addr_wrt_wrap_boundary = svt_ahb_transaction::ADDRESS_STATUS_INITIAL;

  /**
   * This flag is used to indicate that rebuild is required using wrap boundary
   * as the starting address.
   */
  protected bit rebuild_using_wrap_boundary_as_start_addr = 0;

  /**
   * Internal flag to know wait_state_timeout is in progress to avoid it be called for every clock 
   */
  protected bit wait_state_timeout_in_progress = 0;
  
  /** Indicates if beat_started_cb is called */
  protected bit beat_cb_flag;

  /** Indicates if the HREADY got determined HIGH during BUSY. Means that beat_ended
   *  callback corresponding to previous address beat has been called. So using this we
   *  can aviod the beat_ended callback getting called again for the same beat during 
   *  the BUSY or even during the SEQ trans type of next beat
   */
  protected bit first_busy_cycle; 

  /** This flag is used to control the delay insertion in reset phase and main
   *  method for VMM while processing the initial reset. The value will be 0 in 
   *  reset_ph to bypass a clock cycle delay and in main method it will be 1 allowing 
   *  the delay insertion.
   */
  bit reset_delay_flag =0;

  /** Event triggered when a transaction that needs to be rebuilt starts the last beat. */
  event rebuilt_last_beat;
  
  /** Event triggered when read data is successfully sampled. */
  event sampled_read_data;

  /** Event triggered when response is successfully sampled. */
  event sampled_response;

  /** This variable is used to store the beat data value once it is sampled */
  logic[`SVT_AHB_MAX_DATA_WIDTH-1:0]      sampled_beat_data;

  /** This variable is used to store beat number once it is sampled */
  int sampled_beat_num;

  /** This variable is used to store address value during write once it is
   * sampled */
   logic [(`SVT_AHB_MAX_ADDR_WIDTH - 1):0]    sampled_haddr;


  /** Event indicating that bus ownership flags are updated */
  //event updated_bus_ownership_flags;

  /** Indicates if I am the current hmaster */
  //bit   curr_hmaster_is_me = 0;
  
  /** Indicates if I am the previous hmaster */
  //bit   prev_hmaster_is_me = 0;
  //vcs_lic_vip_protect
    `protected
bB7eD49V;^8:B030R()7\XH7b[BUKbNZb+@V/V+ZHJDg4+_W6b,5&(?IB(>J87.&
fU<U.Q79N,K/d3N]T(OYOAG(dHAF+-\,D4]4H:_.3-X91W=NVZQ(faPO28caKF]#
+&TBO92MC[H@ZT7_8Ab5LFe^T/418bLT?Oa54C1a@,AcJN?cV5BY0I(>D\;PSUH4
)=T<Z0,Q6P3-5O(\INN]?6(W.I,WW>0KN+:U=\#)4Jca,N/dDK24c?60Y:_J]FJ]
_2Q2A<a(I/39S8/QO97=Z:FcEU2ANg^73#W+DQ5FTMXZJMRKSbQ)^7\[2LSg-DH@
aAa_b^MG:7gL>0dU0Ib10OCc>7^D+1E,RfC+^^bUT^>C>+[U1_\_60IB&E26]N9R
EP<IF=5aSEg(RFTE8QdZfe2gMYH-+XFCEI96<)e?SUZ#TU#.L#4S-F]VJ\I>KRDS
9_baRXK=aY-GE+S>C5dbWQaTUBe_T_TD-66NQVafNXZgL15_LJRWGS?>@H,\Q:UG
T<OPd76Z\-TDDZ.L[dQT)VEgKJZ\YB,Eb)@#0?:eP#24K?aD[>[LS>&a(I64d941
Z4C8A/K6@&1D.$
`endprotected

  // ****************************************************************************
  // TIMERS
  // ****************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_ahb_master_configuration cfg, svt_xactor xactor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   *
   * @param reporter UVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_ahb_master_configuration cfg, `SVT_XVM(report_object) reporter);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Issues beat ended callback for active and passive master */
  extern virtual task issue_beat_ended_callback(svt_ahb_master_transaction xact);  

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Update flags when reset is detected */
  extern virtual task update_on_reset();

  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();

  /** Monitor the data phase signals
   *
   * This method only monitors the data phase signals that are common between the driver
   * and the monitor (only the read data bus).  The driver (svt_ahb_master_active_common)
   * maintains the write data if the VIP is in active mode, and the monitor
   * (svt_ahb_master_passive_common) maintains the write data if in passive mode.
   */
  extern virtual task sample_common();

  /** Returns the expected address value for a particular beat based upon address,
   *  datawidth and endianess */
  extern virtual function logic[(`SVT_AHB_MAX_ADDR_WIDTH - 1):0] generate_beat_address(int beat_num, svt_ahb_transaction xact);

  /** Check if a rebuilt transaction is complete */
  extern virtual function bit check_rebuild_complete(svt_ahb_master_transaction xact, int completed_beats);

`ifndef SVT_VMM_TECHNOLOGY
  /**
   * Transmit response to transaction.
   */
  extern virtual task send_response(svt_ahb_master_transaction xact);
`endif

  /**
   * Executes the steps necessary to complete the transaction:
   *   - Triggers the TX_ENDED event
   *   - Updates the data phase status property
   *   - Calls method svt_end_tr to update the transaction events
   *   - Executes callbacks associated with a transaction ending
   *   - Places the transaction in the item_observed analysis port
   *   .
   * 
   * @param xact Transaction which is ended
   * @param xact_rebuild_in_progress Indicates if this method is called during rebuild process
   */
  extern virtual task complete_transaction(svt_ahb_master_transaction xact, bit xact_rebuild_in_progress = 0);

  /** Creates the transaction timer */
  extern virtual function svt_timer create_xact_timer();

  /** Tracks transaction end */
  extern virtual task track_transaction_timeout(svt_ahb_transaction xact);

  /** Creates the wait state timer */
  extern virtual function svt_timer create_wait_state_timer();

  /** Tracks wait state */
  extern virtual task track_wait_state_timeout();

  /**
   * Utility which can be used to determine if the common file is used in a passive
   * context.
   */
  extern virtual function bit is_passive_mode();

  /** Indicates if it is required to abort without rebuilding on retry response 
   *  @param curr_xact current transaction handle under context
   */
  extern virtual function bit is_rebuild_on_retry(svt_ahb_master_transaction curr_xact);

  /** 
   *  Returns number of retry responses received for the given transaction
   *  @param curr_xact current transaction handle under context
   */
  extern virtual function int num_retry_responses_received(svt_ahb_master_transaction curr_xact);
  
`ifdef SVT_UVM_TECHNOLOGY
  /**
   * Map a single AHB transaction to a corresponding PV-annotated TLM GP transaction
   */
  extern virtual function uvm_tlm_generic_payload map_ahb_to_tlm_gp(svt_ahb_master_transaction ahb);
`endif

//***************************************************************

endclass
/** @endcond */

// -----------------------------------------------------------------------------
`protected
B.AOc-7^Y=?@HRLB/E.JWU)OBWO^O-H4+OHJ?0VP91E@aI+#?[(A,)bVQ=>[f_+\
TF(+OR3B=;A9CP,P77RMf/&B=gN@B8N,gB,2;ba@GEVM.\0(R\#>JN/E9IS4S]^D
0@070>^J]U<TE[N_K9f4=FP&RP0a[C^#+WW8.)N4\@..5:GGE-U6)&+0#W.&DE>,
]A?N?0AR<93ZZ7NRV3)O>+ebBc;aHE\:7dHC4Q#,TE3WeIX&R-eA)56V>5Wa1EO:
L.a3:d>Zd)ZIP&SWMgG]G?BLGd__a.Y.3IfWZ\9^M6F9WUWTNLN68J\RC?;SSU(5
N=;T,P7(SJ?bP;e;bgCA+ReR,,\46Y\IFe.a4KX4D?dI[WT6E\>BP[7-[)<#U5DS
;E?-/A:cPc;,KV]HRc@Q,b]C#1;f?e#MN9C#VT#^\fHXS:ffBJLTJBUf#RIP2MB&
W\(,U<^\V-.1cI;@7W466R^MbBH3d0S+e^DY1=aXU<@b1FNG?+?]fA7BQ4&/)BOO
T?N&8-A-.C5N?_;#5bD19OJQX+Hb,@W7Z&T0.W<=_F-8PBB_N1g9D[INP?^(6\c2
RRg?\B1Y7fPWOF\Gg@Y)(<+D3A6^_Z]/>1f#fe+R<Z?),f9MU:<P/+=Nb^,38XfC
M>?.4R7J[:=41LAcXP>+2B8?O6\&SLSA[dHILEeRNH^:^@Q@[\1<d)\)=T(YfDD(
XZ:/[ZQ,16L2F@K>_>cDHZKVZVc8DI0+3Mf;L/VFZ,8KQO&4G2<7#FBTB?13QW#e
6g&HNc&>+fEC2>]6[JUGN3M7J23&PeXaXc/67/X@546PT)?JfG_/Ye-,If73U^X@
#2Y+(=2f086gMF1Z)b?E:ac35^KF3TVO\DSa+D[1Gf#KE?V-/:&3=\9=eU8Y\cH;
XW9RE9fgQI;;O0ISF9WIb?[@TJfO#3aO7G3U)2#<.GPET[E;_FYKBd^T+4+V&X5;
BaB13+Ka+f0PUGg:?3OcOBJ?1^PS.8d0YGd9f7X6GbfIc#\@9(4D^X;ZEfB(3YQN
?,GOfcQ]+UJ.-bd9&ESQXKVQGceEHFV;OB6=NeZN85ZI?L#0=F9A\/FPT-\c<ZFR
F-Z:\K+\9393S1cfWTRP3/YW1:PNV]4OAb-YN^\=07>7,#N(89;M^4G(E.A;4Gdb
LJHH8/-9-SG,8Q]+8OO)V=Z+R=7/C304Qff6(X[dID>[DGQ7/Q-PD(:QF>Z(\TVF
[b=5]II-,V16#G165OG9,VeDGV=4C[[Pa5<g6.GD4>?5I6c>O4_&>f&adT,4L7[W
^B2fFYLHE-4G^5RH,;7FOX7V-6NHSa,EdS<\_X=@18BZTAXaaQ4C;BTaM(&]/cS]
I\Y&#G5?&5E4IfY8ET(8;<eP>c>=f8R-.f(Cb#416GK;9;e6\N/CS5;EW<1IWN=W
He+d?P9S2Ya5Q#??YbND#]\G=M]()Ed6.]bO5<QH.2D>@geS-2VNb2XTGa8:/:JM
#/,496A[@:&g.T=YR1_6/ZR4eCc;:2MC<&AXO0TB<4.UN^7?YOLHgYMAcfO(CTc-
AS&AC5(aUb,gX?()W[XJgM\&)@2L,:UT4CU>,]D2Z7?#960W#-X;f&)S&LTTL.UO
G^@Y.=,&)40O:)dG8#gDJK<_>/>7YMW-d-:L\bS@7G&56fQ)W>b8I@>/(W(>KO-^
SBB-:#8RLbPK=A+B(\/acD8DcJ);<eFXa5JX=R><2Jb?#INITgIQ(Ecc]dGX8#QM
J7N04,,&38]6&]DAeENB.KNI-2fbEMA8aQTZU4NLDg0:^<??OT?aK[I[(&dOCJV8
5;I9ERF,U:8V]:U[Ac7E.BFC7S4\&N@QX53.LQGXBHK-E(Q3HEb7Z(3M6c-Sf=P(
T1dWH)?.VUCBdY7dbQ\NR125>5>2,a6&CO5fS#]d-W6&XP/AKS-Z&Y3MM$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
C6&;/]IR5QUB;)L0TPT;527NTEZ^,PVXA=+.<0b2fcPMg8c8\09I)(4Z3\\EZ-eT
5C6-4WGg/Q>7AKa?4=gb4e.f\5BT4/YGFV&bAV;d.ZW^/G[U(W\,cVZCN<PP.1U4
K2^\--8E)H&[),<a0dCD=^CDXDRfePFCV[L5&X,e@95X_TH4bbbZDOSFY]:U<U[g
GaIagSbQFCH\SD0U\<20>=gf@?86K_5gLZTZ-<ATU6Q3,/LcRR53_#Je:f<CO?0N
XbJ)CJaKDdV.eKAB=]NbLM&+98CMQSBa-J?Egg_)[HE5LTMdaH=V=6,HIIeTZggU
Q=).J@f>2=-Ed)L]3]9;(Za(]Gf,RC/OM(<D+I@?Sea]UGg-4ZHf6,dIUMZ<Jc?\
/7_a8T#@\/8FM]a@[53FV.46BYc)a6fFYCB@7g-;U</ME_/P#61#-;#+0Le^fa:G
R&c=#T&1\[XY1+D1Ib3cHCSa:?EZcDU_/VO;@#&fUTL71[11:;T^D>=dNIWc7^;R
/abG:7G]a\U7dQP6#5RL@X@g/&^+fFPC3OgFKI&[L@OCB68_R=CFKMf-WLb16HG5
b\aXKIgF>>OAReIGMII[D:&22)L17;:Z)G&X^GbYe@085&Z2GF<?@<I^5^TE>K12
;8:Q#U4>L)@\N5g59B,dfD5ND1aAL+\FQ,<a(7N:[cUUPB59c^cA(F&gW-&J:RJ[
TA6RO?e29_cWd=A@6,JGGHR3ZF;UD<43K1-M,LK(V:O8;CF693/cce@RP]?D8c)O
I,G#;#4a)/FI,GV9KW5SVE_^@J/LHJWYgLd3b4W6eU>7X7L#YNJT&PM15F;]4OGZ
X^_JS@GPP>5NM[#B7/A7752(823WD1K62NPB>9HEHA5\8d,)>.KP]cOgEDK\Y[[d
+0E:>&96&2J14YRMKXQG/56:SZ3]EE@EZMcAbG=3M9B:0,,G/R^eb\^WA]=XTbOX
8C6\M<B&&EC9GE(Z/c2S6RRZ4FEe>LYOGe>X8Z=LU[IBTKf\/BVg[3@&8C,:&dUH
H+6,-WO/?.7XR1HSM=^4H(P\f[2S.b-E>@><aLKKRBY@1DER0;]gc<cEef#Y5W8,
aTP8PN.2GD2aT3:EY>W7NPB3.W[1VYITNRE<7-,8ZL[P9[_XBV;.?79g[M)f,C84
#Q^dgU#EOR=2I:bJC42./[,,\J\;@>3T=E_,HE-a43Q7/3(5.1L?a<\UPB-@D/CB
8W@Y+JU\7/M#aL<9;GRc/R];FC1F)R[.dPEd7X&1a,;Y]CLENdeTX#LK31HF6:.F
(\I)?KNNH?B0\5XbFT.,H2?6N7A6;J(PB&;M\N;&PH9IP;ZEUR,\#\RV/C1acN>^
TKEMfG-)DT:)6;g6S(g(O=_C&M6d>)FZ+-W.S1)U]YJFE:-(L=2??T[W&V[&COE=
U(Y?Wb7M,VEK0BW9bSY#/&ORdP+2JCQ_]b(H^PXRLAf>9a:J;BdEJ^Qg&&(c=<IW
edOf>IG-M7&35g7:0=c\@FZ6=[4[]\@+JY[7Y=RJY8DMV]0ZKU4aN3B6+DfU9[^E
A&D[^fA5b2_X+aWI51HE+BSX\b_YE-Q1Vc,T.;+9NA:((5,b(&2,3,RN^&:OH0aR
OKeCYXDf6+DL?P:6_(Tee^4VN>U]:e9I-OF,Pgc>FVJ5QKVCCF[ZS+FLPcCHgdXB
B<;fZ[c.BCe]4-6/E-QQ,1Y5(4VB4Yc><F8Y.Gaa/AeI-5D2./)ga]B5#1U72a4;
Mbf+<;2W/=Y^3agKcY89,XENMfP6XW54^Ud\U0T)1G<Y;>F=,?=>1;[,4gY_F^<W
:Z:5[4S>M@4V3fb.0f.)a3)<JKK&_9]FC^U]-/YdL4g3RQdITUE[21/ceMg5\.Ud
XFB^(F3V#BNcNIJA:56.W0^V[L[_Ng<^_Bb=>YZ7&5_?:0PZP:03TW?\Fe\;[,62
V6S8E5EJ;.PW2QOGc&&KG)?JC0Z2,C-C//UP=[C;Q)?LIWO_I09)+5ge>]MP2PRc
(,@-R5S@gaL&2O5Yd5KGGOd>+[==I5,&a?3JM<L3GJ@2N8_.ZNTNX,-QL4eFSJ78
X2Fa+[<-g6]abe=b[c<[]9A]>LZ92>FT3<He?T+RNCGG:^PX=_S.G,K+YAK[#L+g
[6>5.OL&K\5#<GRP?O;0O<W?^-8DCGC&BLDBRX;E-SZME5)b(Zee;4])X\I#^(X/
S6ZX:X+d^D9A5<R[/MeY_F8QEOZ6ZU?-g[^e(^>f7dDf-?-M_D6c5<E#>\\0_38f
1;L;DV3_Pe(6)XPX4K;)+6@W#aY>@9FN26WR6IZdK3E:O4QU6\&O6D[GL-+56CUK
c9>bVZdQH1+?36XaF3f0S3d=_Gf>?;Kc]GbI4Xg,C[#MJWeH)^THV.@@Pg.I=,IF
AHF9VBW+YaS(@+#4Y.[;Q)1gUPLUUD&Xe?:&PAaT8_6P[4X-)C>ebM0\E@SeZI=X
RR#64_-QFL,A#-O9MB8aZG\2CR2:7/W?cIVM.7)/5gO6.]Y&4:+/9Be&,?#&X?QK
E,(RR42QKI)/TgP.Tb30>ZRDOFgbdN>Cb693FTA>J9LO[f5(D<+4&VPK,I\gVc?-
6T2;JY>cCLSM))KP#ZP,2LQ_#2^7b&5([@/B5H:RYH_1F@8Af7V):(C]/[R&ZEA>
gKG.4JSKa4W8fUJf11EE@7#R6GEN&))#IALQ=1(BC4/Z@2(1d_S(36e)XMS5:X:G
=VK]0WE;\<F,J@6>6W+G+DZ2Z-TMg),0N5D1BG,gL:[I3+fIMS?K]GCSKSfLBW_H
WH3,J[@0?R)]<Dc:XF2@cR5CNcM[S<[@]dM,<47fPZfD.9CKLGefd?WE3I3)E@IA
cOFOAFE0T<;fRV&7(MG?OfK:QIQNAX+N,HGP7&Dc:KcC_BZDfeT\5.Y543:<CD96
?OP.=K&^V.R?Jf0J.gMNbM(g:VVdC8g>K4)CbYJ\0(#2XUY6KF<<3bV75S?H?=08
Of78-fJ)a=Z@/@b];I_<GLW/0#[:>SX)4F1#_bAWb?7/JbYK:9CVC4A+f<<JFG+A
e04/Y.THL4-eQ;7=[#U[0A/MU@._HVV[0\1VA>CQHT23c+V:1?FV[8.,eE/,eNOQ
HJV@4DF7Nb:.c0;VZ.#<@>@QX(65YABL.YR]Ia/UKE(dU(E2._&X;KW2P&Ec?Va1
B<-@A/GW;bg@X7^.IY313A[HeJ1C@0/B);]#LTZb:;JUe)ET14a2JV9d/;+bY?IV
@;ICWA73_N\(:]RVF>f)dKZ,[.,.aAaPe]0-PXa_]5)b8[fG37[f5/ZR+Fbf_,,;
]&\19=KB(64+G6F5XD:_JQN[c5O_MWfP.8)cUX;HWd.+GWOdUF09dHV1M+NUS8ZV
<Vc#>>5IC5Ab/dIOC,CXNT:G+Y\^c;g<@F)0eg\2TX,4.b<H5#?VUYg)@>TD0G)[
(ICd6W[ML3#>9;gFW&Y/7Z8JYYPYLe\IRPXL,5a;CF8O&-FS]H5Wd)CB[WXe)_+I
QPeGdD#QWG8R))HYa_JI>cP.-E>[Ia\[K;9O3eI0aPbO02KbPdbY:.AEcT,)>C6Y
C?JPeY,1Y#NMAE_JdbD6;3@;N#T&]V0]809^22U?BY9,@,W6\[8(S7\U1]HA2\[G
#DC>2E[:7d>8B7?Ef6)Y;@NK<Mg>2d3GUE+#b\-@RK+X>.B-KJ\8b1AUd6SfW#.B
CM:-2=?WW(TZYR=G\,6HW9STK8Kf930?dYRAE:b?c59\0I_7U6(.V?B8dEVC7]TU
IY//ML4RRUEEeP2IAH)\.^<HQ^0ZfNV@L?V(PX6La>f80bXXd]1W]f2^(;]#ag<S
LTD([e-Y=1b^TcFa@;O]\K)08F#B]X-^(Z?\O25@f\e\e8b):gGJC7?<.+M7LM0;
U/G80,eGFEb_X3JKG=(,<&(==IE_9g01G=g\C:4=+_?PgfD-SXWf3=Y[\?T6e101
.8]V_U_R3L()D+;HH-#cZ2YdV2Xg8NG+/Z?bLT3:OcVKKC68R7L5e_3,G-7=aO2I
PH:B00+7BRKG3Y4c4R(6YZ8KIPW<@c#?#;9ZK<T3.7>^cf#)7?P,G#V.=7TI^-0]
>bf.6&\9J=R>RW5BT#=1SAN/4(;EaPR@9.[3QBY4A&G>;0ITU.9;4DJg1.L5MLXW
(JK.);/Z34#J>EB#E@<[g-HRMKZ.g:#KIXU-21d?O)F#c<?)D8<XL?5V<b>c=D)&
Z./?M?P#ObDZ0PR,J?UXOf20/FJ-F]eKW);=5[3=cCcD8#E\MVA9WC:T::?#)=,\
-FAcNDEU_N#DfI.b49Q\I(BA;4H6JFga8NUNN7AB]/09OI)8C(&W6@dNEcdHWa<[
Kd#C@TPDA9B<cMZT@\AS3=>bg;XeWN=F@F#)ePeO.7\@g^cR^gHGHVX/_2>?ZH)+
;a/SHdE\TV6[]J/SVB>N2EM]&2Y_Z)Z7VG3VcACP^M[aXN^4c]?Rd_M4FK7H8=&>
P&8@MeX#=Ccf:TV+=99,8<X:[[F7;0T>5M55-9=#/de=.N?]<2_[M@WdfDQ@/463
QSd?QcNB<W^/)18DJgHN:TNF,I;8PbD]BQS7WPJ&Z@3L;L7]V?+2@b3R9I#O=DHg
>ZV?U,?bD)O.DFV;9=@Xa_F.R_6afODA\W/B@MBM;E@WD>=K3AAdD7^X02Jd:L<S
HD==8eVZOLcNF:1/6^21[cbQGBgfg@:WHN#1K2e,]?4LF-NKZ=I38(dYITH#M_S^
.<_:QTVM=CX&=10d?J]+.-FCQT=FY_agEE#NBMP@E=G6NR)1/^&+U]G,#85Yb,4V
,BP5=bL,:&PN-51(DbbKIc@^g2\=S7H5^M9X@gYQ0?R3.6U+OXb?SF_X#d,2f=OO
d+b^V4Nbd/1=HTQEG?>.K.U@U:KQbTW23c[.6eA_0#L8O<I8dBS)QO.R#EZ<)H1<
@>YQM]YSPg^d78;Sd+edUMM8(B?M=39VZFQUWY:Je]=<PM.MVH<=;5BbGE/HSLC,
-^1&eQW;R2<.H#PR_?]cRQYF@DaT9^+V_/ZQ(Y\&<UZ,5:C?0D<6BV-Qb?<?/PSI
d7UdA2NX_SG?\CC=E<&ED.K-10(SeKT9.W(R^(>(bEV-EaLI\aCB?]4I]6;91Z;4
L&E3068;3,2#B0L<^T)RT[GaU/@;g^KRY8/_d5-_dg;9C\XV-MXAc@dd-7C3^Pc#
0+PAY+VP\13K.W,?ON?d0Ka62MdF2O3F.FRK.Ic)@<E&RAL4.:-28_-Dg1[a=G+N
^/(Oc?;8W:GJW;Re+e[#C?ZUVLSN>MY29aJZFg)-8POTX+DLBOA3gQ49MV,VV1eW
(XK:\?531L98Z@X8f\4UI?T=86WA>(O,K:-9?,0:I.SH4(?K8dQ9M[bd4KNP1/bb
PR3S3J_IFE10(;WEWX6#WG:=>.f-<ff@>C3\G_@g7X,03[LX9gb4(]SN\&P2)T7?
;9JcfO0I<(ENbR\3A;ID.)2fdP?HSMRSAcg##dY,.HeN>(7RAU[F/?HHJ>B9GW,U
gA2FO8.2[7^RLS4IJ.,e&.Fa^TT4WR,3S(;KPIN0b<9Kff7,K1=.,LY_ZCOPKdM]
a73O1M5dAO8^d5\d(MCP8a^)f,eNN[W(Kd6;7R>.5#FRJ)5E:=V#L[bKMAM-9aQa
X6C:R&E]&O,2-A(5dgV0c.P2J4TC]H\6QPBTb1.H?N#0##..Aa4Z0@@]gA1N<[ZE
</)57^W\daK6;-eQH@K92J\Uc(:P2J]a&5VV7_>,+8dQARFI+E_D2+c,dF&JJ+WR
H[6P6;aQTOLd+QWMGPfgHJ=,???Z1OZaMW:4J:J_T8G.d3TN,O8W-49_D=bT99[=
XU\O(8Pf,L/GG_.7UXXN]3QKE2bPCUb:L7YX1AS[S2_8+_dX=J;++?:43^Y.M9]?
WQg&>O=abY_]W/K0]R9VN_=-fT7?A8?1>#Z0N4/eQ)E8;=4:gX_g)D_]CWZC9a+5
9:M,VC:T_CUEP\5LO,^#5.Z(^9]W=TCbA<=W([D;<U6f3SHQ+HA;U\@?&Z)=#7I-
H/XH@C50De-1dUD-HY0(YLaN?XAd4Nc:1T4Lg62eEf\TB68VR/a\W)We<2QZIR4_
GS1\J.8MgR7T_A7#QDec;B2)?Q757NH&B@Kdcb^UWY.F3#M7:9BMMF-Ub\,@FOK^
bea=3;\Q[C[M95BI48]K09cF5#0C?D[85P#<[OJK8N-YYG7WIZZD3cPVe2QK.WJK
Q?_>Y>IG<O^?]JL7U;N,W7K:_D)SU];7)YO><-//:a4>62&OaVS184VCGbKd87GS
YTTZ_GDP+^Z;U5\T--#CH2-?T_KWAfCF1QGAcR&RT(J4)-OcQ:0DBNHKV/N.]N6<
c)LC&f-G84>d_J?DV]X@d,=5W9aD[BgDEPQ:Rf(X\RIB&/RC;B7P]D32#,+6XdFe
c0915XeTF[,;a.P[Fg_3X1bO:OEF-5H4KD?@aCVWOVBQZZ+6-E5I</Q#B[<;)G#e
ZS4=Z.GAe6c)(;MP(0YA4VNc@Ea_-)66_?:D3cW22S?BQIC5]--3XV5D6[<c5)Y,
8#_Gca5U>D#/?=?E#T+-?=C<X1HH+,FZ3W0ab_XE5bGITgG.\((0fgPcL,3M33Jb
Ad6N6e?]1d6&F@B?MIC9W14U)Q+FC=TNM3EdV^aN-L:CORJA29+X[B<#6NLR@10A
#ObW?KH,:Ve2ePL#W0S87QPRc1fSaHMYOMZ+a5MCU_6NRL:f>E:f-&:IGJ^ZBC1M
\W4>2+=+D]Y[ZUV88\-M7[LS7WLa\6;SCMU0gdQa&8,74@\Uf79C_RE^LL=QNe]a
^65RI#J?e2-ZC/?6g^&L:SDCbVVB726E;bV5GE-SU5CC<d,#fK?>M>QWMFM<3YgC
SUN/IHfYYZA-.e::-aJN5KdA;Xf4:9PX[UNWK(SGeU6+X^-:RHEZ?=R0?Y&@ASZ2
>aZ>-Ya3dAEACc\;fL:+X@_32]#_f(/I[1GH=.MPVdG+?@O&5_4g>HgAAI#>37H1
;Cbg<3J&7X2?DQRX=,873CfTTNd<YQPE2G]Vce:a7AYXV;G67IF-]XBT+Y>b2Oc1
?9)/>Z6C-S-(<cZKZIa<;L?/=GQ4=3LI:OD03<9?)<D;A2FYJ6@T#)bgD=]gX+[D
2/YZ,67[@Y#:fNPKW898LCNHNSd;>8#5J\W,&dQ)>E&G1-C<9E2J#SfVe^B&-KHc
10@<+aISCb]/G7;2,5M<EH@3FP]>@cK)+B61;_;JRG45-<ZTb-Z)/eV?dbXI<:^0
&?I+gU>,[O+H\O\1819?3:E1_GBQ366]1QEE@<8ZQU26bed,>BTa\JG9LLO#<G#C
?MNRHbbWEBVSV#bfARFVVZ/bUC#3b6DB&;CEgQa)M9Jb,;)\O5gO?DG4Zg1^K4Z#
Pc^G#&(7I,BK(KA5E5EW^)151M/g6#Mg69(Q),Y;7,Q(I[3G.EV7)O8:?M@c#K6/
\BKe4TEPfQCZ?<8TYca@g\;AX&;A9)bDL38(CZ-;>M[1C&HEV<af#2H,:IKT<;YB
YO>NH#[>57XL+4Q[.f\fIO=#\^MV6RM[d/_\LK,N9U&UV7W\I>LeKK;g2T=g.FHY
-W58bJ0O7D>dRC5^Fd.X9-c.B#7FG,8]U[FL>JP@M?UdM=_04CN\P+\#BeP5.a6a
NJMJA[8;D^:D852_\81dAY@;HKVCE<J6FS5BMb+JPH1b1NHGV)/MMN&[gJ_Y3D30
W0\76KC/VKBORP,92PR9>Qa&gS/H36.4abeKQdTAL)=eOMY(EGDDSBb(ZfMJHI@>
:[1@9OM4CZ-L]f&QWCA&^YNb3>&U[&:Q91]8MNFL4VI5SWT9.HVH,MH\B10>Z;H2
:2=a^\#H(d6YIX8CY[,2MB[#,?g,SLF==$
`endprotected
    
`protected
FOaS@N6=:TE7b>E1YHAHUCW4H4&>fBTI[3I=LQN:_=QH0?(L-T>97)AFS?a^E_;N
Z\0MVTC84;3Dg21b:&]><R9HEBT17;4MY#@_LQ#A5V7;OSVF_;V/-E?5WR0J:d[a
GU+WW&0W;/2F(=E(d/.P@&V=ID1N+R?H1<O\K)59g\-X67=D0aGAeH64UM#6/OAc
5]P4b_Q)GI1F-$
`endprotected
    
//vcs_lic_vip_protect
  `protected
K35Y#dF>=7c[c5V@9G+R?3^C-_^F@_,#A=BXY3:,NX=Ie;RYX_:S6(X76]6:&FA/
&B;.BH#Bg]&9-Fg^=GRGX)02bC/cUZ>VYFM1cS4W\ZO&QU:MR.N&X7E:CQ>;J#2E
c1.9>I0>X<)&R(_FK(VXMOa<;c=UR0=0fH(D<TTMd]I^WHDD@4[8-E4aB:#^ZN;<
>DN4G:)S6)R9M>cZ\S,D,-/,S79ceM704_-E^O,@CO+M[@dW_V.[cX?_DRB)U-CP
G;[ZF6]^8:G1JE@T@3Z7aH=N>HU:4OET+/I/)aLI@?/?gQc0bRSWC:R[0&G-Y+.Y
YO;2^>.RU6\7eCbY8^=Zfc/1]A[,RKCAW<Q;bdaHWa,H0;I\\C)]_R^?f[POWV-J
3)OLe.GSL<JVQ)B7KDf-STGWe1EV4H1W4;T0Nf+X/EHb0_E#J1F\9>X2H&;1cMeV
87GH=_?=H#Se))9\#Tf7<d9TK]W?aHf&=0XSX.,,6SGd8XML.MY&A(7a4#.D5P7#
?X[EYcBFHXFL\48HRYDAF=FT6#\fEfFDc.V#J8)]6eM9X::M7fB:?6DQ-11M0MQC
8=R-#/DOZ1P^Ob06ZQ9U3CgKe3/Z3MHCK_Z<8bOOB.U7)ZJOTaQBa\)OXaN#75@.
.D>0(/HXIL>bG\>GO0W\aMSP=/NFDBG:-BY5LN&GFE@0b=2MK^\Z>M368^&]7CZE
20BWKSU>5XTb/U><XbeY5cA+J=HA(b=WgD4=0E#W&b\7/[+6KW>=\f[P5Hg;a9E8
]/d>e_O/)P4?L-N)S)1N([OZ85BX-JHYC&@L0,T]_80d#aMCEe-]/N.^U):I7CP:
_#fAG^/-DF[.0D#:E3=@,2P9Z#4L/db@<@E69FB9\.:8Y8G]9_@2g-=TFEB9[,>U
^7]E?T&H)GL:GKP@g0?M@-g5EKPB#Oc,_8RWf#?eD.-:cM=FVHP,TU+1&)4aAZ)&
d9(W#1K:7]?a\=[+K/baGCTfM.]@8;,U@FIAHXgbW;LSCD?</Q\1]K-:U_E#]:ID
e#Bd4N[:.HXNgg+83bC_H[b21VTRJ5)W[+_O+)>W?6G@Z5)IIPK.WKN6_B[R+fT5
QUcX9&U7.]>(9S(f\9;U#6XU#8S)-?)1)72QQ\[Z]P(2H8>R_N#E8d=B81>XBeXc
U3+W5(#=8_&&GXdZAN#J@_OZb@cdURYAIO(D.Fe1>N@eEUN-HP.-Pa2R@Xc_PBYd
-W,&+&3B/?=E@^<Ha<[.G_#^T@g:,E0GBaa^Va:2ELZYRLFJ-@de2\R]H8X<TIS[
F2V6V)bcbP)G5UQQ:d7ANU[VN<Adb8<M>WHE:Hb;0/6-SAX)+.&X1+L>D.FB]+RJ
M_bHA+H5EN,HXAVEB@W<c5RXLS@ZTa-Q,0=P<WG;V1BWPUW_Ye.-KbPUU71_.]>1
\9aDBfM(NI-1B\/:\?SZ4EFe-4M#@:;a=]2(K?^F<+L632PWQ/[GaPK4a+R2=W\(
.+WD-[4Dg-Ja71I,04\M_AB8K.&LGGEU(e=d88CI8PU2T1gPF;7+-B.>M>bQ1dGg
,<W(5-X=d\TS^d.a:8aL]f6.0?5EZgZFXU\=[<:46,aMGXS4FDY/>PNcfcY3-TOb
&O]R^7KE]&5Og4;3521.3GCY4^.d,d16A0-(WV4V09Md?Y063Z^F&PED6fUGC.+6
f@V6Y<&M2+&_f;gcVMD;35#0PTWU&>O6Z-NXM9,KMI4\ZeDK3dEUeN+f/4R_[^RZ
A4)-(#T3(f;X2L=-N::XTU79_1-7#,AZb2c6H>KcC@GR.E@6\5>ZP@DI1<Xbf._e
]g.?\D.8SJOA7F+Z6TCe?LV)<^X00Pc,@+F=Ne5IM,92G1=/]7V_FXOFYa8;1&af
e_5-=[<GU<4d\1bHZ>8bE,B+RCBGg@D/7c#(:7@9)4?dJ(8C@Hg?>UP(<8YB@Ra4
c([,e^(3#++SII8-IO41)W0/CS&Nd_79LY4;ZMZ1dCB1_(+_I+f622ZXP0I5P\I>
1#1g]4>HDa&9TRS,(&d]#G;QNKcSE/+T29P>UT+T>,9X,5aH1?M+=TP+1B9TAOH<
DHDHRS,\/L9&IB9XIUb&5P2(-UD7OICYP@dTVgFDT6]ePX:W3+,,KFJ+Hd:)TF>0
4KV(<6AEabdO3DCZE#9/?:?g&BE:c@-DE(YY3:JRCRe;F9dR<&4&[Y;O1g?P+DZd
JE@[eM.F&##XHYU>6^CT00A&Xf5>O)2]FQU=)J@S#IM86Q4b(IAe,Bg\HR?KceMG
K)8C^3C73Z4?FHI-/e7+0XK#6[Kg#[V)<7@GZ,LeM4?JM,Zd?L(d06D#@V,M-BS@
V0R.V<[a]AaI=[\NP16O#+JLU.@YZ4G6\6\C4YA]gLdVRHH+D@/JceC3,NX57NgU
WMB?&F]<7Z+(G6=3g;[VV1;4gHX@aQO69eO_C6c0Z93\96fC5XJALREB+V3T=PPg
F6f8,GPN?/AY&F&8W0&8?DU._;N[\^V^TH];QD1P_fNdVN?UG@.E15ME?M0RF+d:
EK(_2/<(^+\a^N.0]4eeDb([Q=/aYTU>IHW39#G?-Y3XHD-P5_PJVf#,b?IG;FIT
fSZC.gOO]#TLNV3&,;aCYYg&ZUW+<\2H?/8gc5NL@&XfV]DaePV75ALc]QF\PfXC
WG/OVeOf:8W97D7O=RH\<MK6&&^PO8IdXgZHR0dIX-/YEP(LYbTc-CCVAWeYdeLP
YJ<14.-Q8CORM]A&6;SNdNcWGHXbZe5\ZU,ge9[H_FM[2D\cbPR3.?F#C8dS6.,_
6c3F9^4^SIHWAbITg^FO+1@+RL],01@K-C;d]N3(2=<#J5]M6D7Rf?\-G3eG;C]9
[=12<SIRQFCL<C>=\_6>9=M2.NK+DOHY1+-,WO=a7dGX2#\2H2_cN#S0^P,[9CQ3
JaIBCO[8-TOA>?JFQa1Gd99U9&e>f:+;E;R,#OYfLCM?(Ua=.42T]B35d4>C(4Cb
QZN1V>bQ(d.):eJD@a2bVIJBMYSfJ@<>Xb/b35gPNBf@QM>HRD?#QdWXX?RDaTB/
4)VR(+b#Q1fffRg&cIaTCV=+HRDH(c#_9<=.1<JE<EWJ0-Z[?a/;:]J=]DP(:K2Z
@QZQ4N#\P;M;\M_b_?9DQgF4EX_UK4K)0-(XfR\B4#0-QC+GD&C)egD^DBXa#MPD
f3_.(a>[d+_@L@e9G7eY1+V5PX<E1AH<8RBH51O#eg\09GXNA&;(:TN1_T=V/15\
-6[K=1JLW-S-Fg77.1a#\(dEWWOS@ZHUUJE=^)aVL#fD(<g1YY7<.U>D91,OH^PY
C&7W1S6c]Q]OGBN1TXc5YNT>B;68>4>MS.3/5a^HfIS?C^YGDPFT4K\Ra=I#IVg>
E7aN+U6#EY?KGJT:16^Ve7)/G^M+Ug9,FZcP5fV/39KVU>HY3eDVgHSRB6,J,PL>
059=Q\)WJ#\7Q^U(Y:Q5026<:F/Sg8OdPYDI47>>8\\.+:;FR2GB3f(J#GJGC<:)
KWP8)Ob(]bOB[;](^03/@=0/W=g/EQPPS@eF/JbMa\W]FPNcA&-=9T//NTR_TdQB
2.6cS,?^VHeY0T_DWMC7(W\dc/^Qf?9ZG16,EIHT5DfI:L#HI6X]-G&30TR#7gdX
;cX<^O]++HR<RH-JUd,Pa.4/>T54R>\-Kb0<+^V06>2-\M:Y9=DTLNC+e<N&K>H?
d[]G),^+Z[2:f?\gbbBV7Bd#7.TaN]&RXS),()f[^DcXZ(?-8<8[CXM5H6XIX<+E
GdGaFU+B(58W;UK5H#T1e)OCJW\(RCcW?UM=E1AUg;)A.<X)AYbOcbdJWX-+192H
S,TX#UU#ag)G=WG,@KTEI1YCdO-d/DGY;g+;\(GTd;<Lg767)QOB@A3]?C3/B0?2
O[4baV;BJ]3C,Q<L?M>Wc+a-PH=;@H1HN;>Y(9.1&Xa-QJf;@JZ07I;cdK91BI;c
I&1-L)47?I>.K?>Hb>MK<3DHPHcGLeM@>Q[M&99g)IXO<)C3S6]_E5-.C@0C8:W6
E0^20?CTc+VD0.?F]:DQ,.X1MU5;IVQ1)77aX81ESQBQ)D?DF(4FeN?:/5,#+/3\
eOId4I#HI_PaedKT/eVceI7J,MI+[^gf&fDP[L-C?[f55>N]]dc:MD(4;TLC75T)
gRgY)+T7,@@@?gg82b##1/4I[3AR&L#X3cE&)?cMDC3=OG/T6a]W.&G:]XPW(-/5
&I-ISC&.9[eG6&NO=W[=Bg.0Fad<Z/NV7C6I6-?]T51+U71(c+Z.[X?6;GKeUKB@
Y<BCW(YVYWA(=;a)<4-MQUVe#]AJ,8J]YII9Sa(8JZL[6UP9>+B=PT&gXa9,/ESF
BDNM#\3WY-I#XAZ@/XYc;&5>J<E\7HTE;6YVeK=-1<_6CV\F>F2BZ\-6fJ2<\FDW
0LHQRU_[UN).6DWD@S(eP,UgF66]dVV<F>I9>OKFFCZ=1g/#e-U[@DL+bOMDZL:b
4N-D/@W/[N_cZ_^/,B?e9BD=I>3:7]_I@Z<=W/VF.7FBBM0XYc)0bN>1R.E+PG_E
?Ga#T5,1(T7IJ51EF&W[QVfC;83X]S9LPGH;N9A((f;c^D-MU+U;Z;10I-:62g,O
5cDB\XD0B]Q,?Rd@eLSNbP8O@F30>I4WO2\H9T^[X2IGBUL#d\3[XR3&@Q#V_F[G
6Xad2@8+2a^NT1I]2LO:+]FTT;-JA_@]7_<CDEG>DL91<^@#=\aAFU02(8E=S&+E
,KWJ/O?@VCe_+BJ#<=Za21A8DXCDcT_XE9(O^;]@&fJa_Y,^VdMcNTJ989=Qg)FN
<7]9OJ-X5-9PUNYZPPBX[)B.:@-?SID(R5/,7O\JR0]1]-M,F:C<gg@__=<Z\7KJ
Df#0=PVOM9SW#-[@K2BBI-G/[0f0cS\&T;94K,V9@a/2RAWRGb\.W:\M60VT(R5N
/2GAgUOG/+3T:[+YMJ=[,CK=(UUF/b_Q&c:P&YV]/gc5a5G<gM>P\JG/YF]U/\V.
EO:)E=[2DR#DU8;>O[\e7e-&D<dbD))G.=6b,ENYeC5c+[GL)[A0>g<=[-=WEU=X
g@-6\:Pf^C\_(Xee^Z4baGV75C5#Z&#\^<PP2NZRP\SMAeU:)0Df(g_2VJ].5LL8
AXGf7<f05#,4a(V]F_=a1efT:96b3)HPA=Vd5Ge7Jg6Q&.\6SJ]3TOI5_167P\Q6
JHLU6\HT\S_79N?=#Z7.9CCM74dgO3_aOdE\AF[,CR0\Ie:45[@Qe?9)B&f[R4g7
I3MMb@B,F2-MYX#9/L0<c@1HH9Y^-KD:d00fOG,R,4L_?Q6f(X@CD6=[8cZ..)[H
DE7S+eCEd69R#MR&DB^&ACQ6@=->/1cN.1+D:F5Ge61TJ86KfPH3[8Rab:LcgF3P
-73,6^Q9EAK0+d]U,7/_TZQ2,.[X56@a62R;E,H>1#;ABdaI:JQ0[Be=1;5#cI:X
Hg)c7[XMa()3=1#a>YC_+dN.S=NCU[RKM7.+D<gVYS6+b[1aJ7G.<-@U]H_3;9fe
NG2c@,MA;)c1FGUA6K+B>8b<[e<5NOF&/58;b2WN8Y_;^>(\+::9W504&=NP8F(V
J8eRJ/_UHV-Q]+cZ@Ue26DJU7Ba+WN]\^VWWUf6G+V3+-d94[^GETAC=&_@LO+S9
=<O9VaWTWM,OH#PEAbRV]]D--VW<ZH3<DQ&?M)gHg<GE<./.FW?\3NPE,NXFQ)J)
PEX9<[QJb&YRLG[.?ZYMX=+g5=HdJ&LCNGJY<B4)?V.ZP]2H#=K2?-QFK5>+Y,A,
,&;:A(4XXJHeH+K^8+E=bGP\]gOI@Hb23C72@@95a&Y@RV.WBE=[1DBSVC1D0XKI
E7N(VK#+[YQcZ96Q\#5U^^dc^D@8KTAB[_D^].L3d)d;O2F93LR)dBfIHBLP)6f-
c7eLf4U_+LBOgXfK20TddAI:&4PVK[J@bB;:GBN8T[<\&A<gef/1-J]EAV[7fT;e
g(&=I_)@#3?UfRPFKBBQ:dRX6(CV5<1SUJ;Y&H-WNNcIVA/^gf,PM6+D[a>gLcT:
d).#+@]aT#[S?YW9D-[HF[C6H2])&LN9M8Ib)d1-E#Je;(66V3H<4[fHQZ7Y[G?c
MX@[-1CL#^bIT5?^#,M_=K>1;3_SVWM5I1W>1[K0=I(EHYZ@GNcD[6bZeZ+:AMU,
A)KLK#[^W+(6=8UX?bO5I/XC6>+QOV1HEA.Xa&B6U40^dG/XbV1<:46b+aEb5UBb
1e?=g@(.#;O\7/fD8a>ZSBLT/B]=)03\R<&4<E/;TAN3L/^8cB4&YW-B2].Z#J]P
7[97^?(H9_UKC@=:7D.-@#QE+4FC^8+H#2NQ@V.aIZ?ZaeJZHU2gSHF_#[AEUgOG
#/)SYDOG,Re.VPL8ETQ+M-:T:XB#&14^&K.+eTBg+)>J(_SVDf?C4\YG\=aQZ0Q7
DPf/gF8#=DW8M.@33&f;LO1><A._4H9SUX_UR/#4DM>8LgFY4\_@a[Jg]@YJ2/<>
3R8G8PTVU)2W@A7d<BE@XY?+QP;QIdeX=M+\#C#d5]HK1DQV@)9Uf;:Z?K3X6EUZ
E_ARUN07/C2>:4&1df5R1e28&D)TBa:6CB+7MM5AW+a?N86&2+77MX/JTf+]2:2E
gYIc_E[/?a-#M>3^TcaI-T3c)U;e<8Ab&2b?:?+d/E2O06D6+ME/Zbe,;d9Y<_HT
ZZW9\ZS;#TD@(WLcERES-4G8[RJ87fUdG5^>GA8/[>^-Lf6W6A^4YMMFNJKXL7NA
(Te0&3S9Ufd5S.HTd2+\&Z1Y[.MAJK0GV?=,f6A7@bG?&\=&W)Z>gPg\A7IcL,_N
cc<M[SBJgY[XTRfJHc5]<3Df)[3f]7e?4N&1UVLg/H?;V#&/VJb;eY5PBR3DB+<G
@VIJe4CA@M)PDV6YHe&JE+.JP_(Y#8CJ79X-;@@K&TXRL<@9eaR\H)(ZXbMI[@J0
N5822A6_))cX:B)WMKB9.1;S4?LW:SL54f:_9@.,Q/V24C9P+Y6#b->:C)9&[K93
_b/5C,T&)cXOKab>-.IX:3e<D2YG\&gBf@H-=?,-?LDecVJR=@eW[2VSQ6+-+T&7
BZN.H<.OR:0@LVa,Gf@K?G4g&\cEBMN:_c[B/fP>NQV;?87-8]g/Mb;FCI;bAR/-
P-J>4SC55+S>d[(DTDNH+A,[]=+)J6;0AP&9Y=#S-(V#aGd^QB2G-b]H7X0T]:/#
,?&5,/]7[WUZ<e.[E4C+2I7f6gS1[#;GGVe@+;LH/?T5X2L3=2I(W6C=1<^ZN1-\
c4?:L;.2eON\-+.=e:7MCa5Cd/>I]+QY],QJ:#C2aP7SgS/T#dO)PH[6>/LST&ET
]Yb.9aAL.g]>6CMQ5=;Bf];:,daG2V)]9O/8NZ4^VNHU?R3<)@/9.c&U9^();4^3
0(7ab?=M2^g7CD6LO\X[7_(9Be_SA/@(:dLS+ag9.QMReg&4.d?8/=]XX6gR+e+6
4=_g9c_7HANS&X;(NS@RTb:9=MReZ#3IHOC8d?J2[<L&72cRf:^RC79aHE>&QR.?
^00#bT&DM:6HW+R2LSeW7X4(5ITb\77-MYX^fWgHK.A2X&/V,QD#4dH]?;7ARAg-
+KXaY3UY_F:f\9B1-Qf(6eN@?bM<A_6TFZVTM(Hf-DX,XO@W,)EOa<^>58O](;Q\
#8b>CKJG=D]#6Ce,;BG.#3K,8ZCN+e-bgU]Z_,0+\?QW>9W:C(ORY[ZHeAJ..2><
:I1g(TMJL-+VI&3f7K\;Y.?);T^-TQS7P#Cb=,]?;AJ:9M/@;:=-?aYb=6>1e?(8
)&K7C?OXG.>b=+QGZ-e=9=G&C72Gbgb_:O&>V7CcbbP,^G?E@9QgCf6,/54_UK_K
S^QBK4[XR.2TZ(8bECPPB6d]1VV<JX,a[GO3R=ZN1@,Uef9/1WFWGRC@Y2DO=f(;
#.;e#.N[MDUabR<8eV.P)LNM7TZfFS>[^CbdHRQcbU]0g3_Xc-M26+GUBEM,N&C]
Mc<.;+=0:=a-SQWaVSMHbFV\\>T@ELTH8c0c^;[<)UUe[WL,NG31,&IJ3]+L4Y8J
U-V]N/1NF1<cb#O_T==(:?=0MR,ISYH#16KbF5]W@[#bD)a8ZFA:e^;7@>4@3E49
17JSGPCWF=IXA2&(b)f6RZ7-OJ+B1#F>I>MTbfce:A7f\VM@Vcfba[IMZ=b1Q/Ic
U<7LB[]OF+A?>)CFB8Z4TPGUA:S7Te)(>a)]2K0^Hf(#>c\S[Qa8RaKLYEH>_93-
IN.;:&VJ0=W_E,N__]4_5L:<^3Cg;/eY7807e&TDU9Y:MCRQ3VV<=/(0^8/6VF)9
7:Wg8T^;^ZNU.+&OQ]R]<V[]I@K3QDP(L)6V0XG(&+bE7F1898^W@:+M/52(,Q8&
b+Be9X5dDV?TGTWO8a>B,WNPBBDeC\bKMH\0S##-gT9;NQ4NGRA]3eN;ZaQ88?H5
))ae8IEb@c83Qe3COOY96I(;f7Zd1Z0XR4D-DJQC@IdMeV+#TCQ,E,cMK9L<F;B5
7Z-^D>I4FWSe]e7C;,;=a?YEQR7\O/>4gbd5(&g4(;D,1KZ28E\O6W+6:Z/Sa.G+
/.^&D9@09^5C,]dX;GU@d5RO/=@<KE5c;.K)PM(a)L:.874GI:#_^\_-2TN10f1G
G8:WE1#F^Da4W6@J@.S3___d(DX-BC5NLEVZ9cdF3-bDZ=+UP3N?.-4O2.BB=S@b
N.+>4,,(1(cXT/.BZ^SVeA&6C&HJKg>:8N#ML:>;:S<S,T]Sg-H@aNWT)-c1@N?U
.DI^[8Uab?O#Y\f,,C9+<E6aBGYE7Rg:\0c/NHU\ZE/MgW[M\ALbZ^7EHS/GDXFd
RUdXOJ_.EX]HR6G0Q?gGaCLVC9==&(fbKLGL(L[\-/=G?C3P@X5BfceG2[OQ_I5A
Y&OPdMAU.\CGDfNf_SKS&.7S.K.g]4I=+Y[eA&33E.>H.QV_2fV:22@S^3E=9B7,
59>8]M82/&WNHM#YCY/S5U,H4X8XSEc\M+ZZ18MCK#,H_B2D(e30gg@0AVf]c]We
0@6++12cYWSRZ]LI7fgNP^,.7aL,:#GH0U2#QJG--)S\.VFU9=]K0H60;Yd1f[\L
WDN6#TKP],:PRd\Nd[WD)72I,YPD-TD3CO3L,IWcY]]G\&.2aSQY64WW;0?8b\]5
]a6L4GAURDTbbdBX>gB_7fO:Y0a,F^U2#KGB;1)4M\30-&e9MfYF^:Eg\>7&5VEg
1,?^#OcGJX^YPRbCQe27RSL/:a1c#e(5G?HSa+NAC0eU[6IN7VOLOgf0VS1>#)YB
<X#FL29\aG44(a@GbCW@QX1^LLU28+BVZBHZT.=e.-\WZH?;^T52P,P_UXb(5Vc9
>VbQ@)(>8F+d<XS5V/L.^LbK1O4X,\ZcdP7c?>V<66,-E4QK-\g&R5M+F6K2OgQC
89G@RK?2S[3f>8bDV1&;84]M,X_gNPD0(WUYb8Y+3Y1.b]#aKZAI1_Z0OFCK>SZd
@T9Y[WNIPNf^\8<J2GIEEN):3;PNG/S9:>CZG4HW&\IcF9<Q]13\Ee)T@IP.YdQ>
1<c&:#3ST4#Y+(G48)(HC-\Q&<5<XW8^C131B#0DYg9g]AS-@N^H2@98GFM_g:?3
UW.XP\T=[OV<<@:g=&HM:2?L/BA8Z;,,M=L[;,=N0W7RF^]X>>\NT9_Ec]dM#ObS
/\[83)ZO0Q(LYRD=9QFNEe1TECIKg6SJ9V)4CK.DcLQFac;L6XE/92adP\N/=W.B
J#L,3gG@a:4/]KWfE+SX.&J75R(MUP=.S]#S<,&&DH=Y4N4U]K]D/]^]F=@6/-a8
+X:\JD4>VKY]@Z_M2e3\SA,:1a?I&E^_#Z_&BIT3)E53LHL9A-ZJ,88QCKVa9HU)
Fe,=DLeUQX:ef-<&2=U:c[(.]W4/-&a50\]3[-SWWUc(?<?;+=:BOKW>IfHSX^)J
Z^06dY,6_WR,7bUS/931>)&RN^BH79H&a-J/RAH0fCeQZ840#:M12]IDE?;/<W5b
57@d8,QY7a<&0LC#Bc[S@dJHeCdG-,=W&AO[9D)BW(98\+)O@fZ6_Ugb^>DS=IFE
aUVDIQd(Rf4<V03&7H6Z_Ed?dCc:23_c:b3VG?Vf>VOFV+e>=^:Q0Y1>KWc\]21b
d#/fJHfc8Z[<OEa4g&O]TA?8Pgc=1V&_4N&9:O-a8UVa/#\I<FNQC(SZQ/#13_)I
O:dOEUG1]#R6>J023efPH6aI6MV18f3gCDc\9DH:):[^C39<:H5O3);M0-H:+[aW
Fg4dg-IF0:.\^0AKJ[Y)9GTg9=BO?(N<Z&<F5<^AgV-PH]2W8M^bUTB7#bE/a&P8
N;1]?@gWcM7+?=X-a0,7+H&T.gLOH[6VB23X7OO,MM20)L-AW-5ZV2WC+\+.7.NR
)gICae)D[[>0+cT_F+OU,N+Z^^BfgBd3d6W&LbO4002Fd\\A4&AYLSc,RP0I9B8K
RUSeX+CBX_a2fLNA8&]cBQ[<^Q.ZaZKBMY8,G)9E4]T.PD1:S=cB<)(_[HaN+-]G
SCZ8\<XcQ\G)C2>DP?;6_SZ@._AE&QI?WC,/]Z)DKZ,Y7P(\F]VQ],YaU_;MAUO(
CcI,V?HO2M6VMaEK@.B<?LCg.V:<@CISZB]UU/IB&S[@R=Ada5AIM&f:CMLQ,WJ?
Q<[T=A16B4]4ZIR(?^_5g0TUfP)#EKSG-@=/.76Uff65>\dIV2gD^.M.e3CT>5TD
^M]L:d,\)=XO&3ea1;F346X0?\I8)7]Tf4WD;#N0W6P5;f/9H:.f81VI;fZ8J1O\
9WC@US(Z#dB;3EYV.>NLab/UcL(F7cJe2E9.5#D4g2g+;geAageH99^#9>+D4a0M
4I][0F:7BM@)2-@<TIOVZK]HR4-&GRHG/_Xa@c&YKPC,89U3#2ZO=gAJQ?Z</=b1
XZN&e\XXQ,8ZJb]CXAXV1:-YOaG;dEZ+LG[(VcRO0PbQ0&W,O)JS_]cX)C9@1S0]
O:#b0SP4f.);(;4d#@[<LXe#?L47-dUCJe,(5#;g<(EG0TS\N;5-A^,^PVgag?51
-TR?<IA?\c7dFVbT)&1JGIWLc;5/&C#gNb>VUDV]WDW<gUU=EX1T82N5NK?_QZc-
M_]a[C;;8+9\3FOK>Q#:ag??ebJf7Q,?.SFaJXTDGO4fV213@CR+<Hdb&#9b0#a/
,?U(98WK(>=c^<DCQ)U()e2NCO2d]3[(3G/BfYHAIAM>0,FWfQd.ab?JY.g?f>P(
DD/4W1@-EPWI>b5^M]#L?LgUDW61)U=IfSdNNA6)@?3Jg#18Z]CKAde=AcNZ36(\
>Nc-:B+G,c#PZIdI<WUA7ZOT[ZF5>Y@5X])WcA>-+,;ScJO->WIYA31TZ.:b8<DZ
<J]3_.4//ACM=R[7G-6JC_dgKJKD>54GGcQ,=fAV4WPWKNM0Y;?L0M00V]IY5[b(
ES08)6JA.IKCe2(9:5S7b8AW8_[dWQ-]EB^0b(TF5bgIa#W3dH3-_3P--FCGP@da
#GQ@g[IAG/TX5D[X5cRDCU@b/BgY&RCHWcaZ]=\PI/TZG1B9065VI=(Q#3#(=A4>
L&C(=;a[8a#6<#WX5A02E=>)J#]/U@e4KSGF>[&U872(L<^JJY5.gA;M^723G\:/
7R>I>2.NE6M/e_H9N&e@Sg\^]2+A&]#0KB83^cS&)4N9^CG2<?[F+PD/B):T\gQ5
(dQ51N,(1/(<Zd085LH.C2aOMO.bEW(C:cIT8TNG]eK+JDU9G1O@=/AE53XfdRO-
=O<[)1Fab0U-GZ0g9Q\2N<Z)+>S#\MO5QAeP1-<GeY#bFS^P]2B5aM(S5.;fb^cX
UY\ce15[\CK+DF\JC0JZ>=74R?X#J\aVUH#VJTP(NfGTZEVTcG/]A>PC_Z3RG/^,
.+<bLYSd7(P340YD3UG0<70.-7LKB2V?JY)X:B<T(ISa4g_TXb-[D6>=Z6,U?.RY
b87-3U.VEJ8CX:]D@)AT^[<C31N0)59=RM]5AE7f.-C4QFH_MDV(HWJG_0^?U9+C
AUEM)2IESQgMAX^G<0dX\2T-?;&OYLNH0>Sf,W+P<fC\N_+8;PDa::]g3d=[b\AY
)Q)@geK6#;GHJIMA^(6DP]Q\JLM3b=6WgCb=L?R\O1AYgMOALAOEd76@eYX:A+gD
W2>A9@C7=Qe9#9(AS45_\D?<aKLAb,UT>ag;]BD0g4N]Se5:?L>Z:T(KY.D&Na6F
\cV-+W]4R0cf6OJ&M@,5PA;aX6#QWU_;TVY8I)PAPQ5F;_U.ORE7.gPPE61@]5/Z
[(TOe/A_>2AZLANbP-I1bCWJKDQ;1<g)bX)\?9S;VDP;EK6Jg=<27?>8I-e2b1X3
XF4\?,?N.e1+>eP1(]a9K_/Q/c3\.Vb4)(Qb=;3Q2?M=>Zd]W7W-6HLD_GH:B-f1
P1OYX9FDS)U6D<0M87ARAKL&8eaSBbY9BEe_ZL.CT[-SXfXRW8@Q]8VeU<A_L>dB
2+\HWZd.8.JNBea);KeJdSONY7ZWT_VXfd]XLPb>/O)L3dC6&KL&eWbFPQaXZa:.
(N0d#0(VP).1D:[+H8<F&2#WAMdS2F&Nb_4Dd7EK,L]+;0gT@H##;_,OG55eE]3^
\_US-YH0.0:I4dfPPR@)EE)QHBWD^B(P@/6:>U@ZcC2fUe,?6Sd?Z57YH0J#>RP&
[]9:K3J@OLQ>]Mb83dE+]FHa9#bg-F+EQe>+OX^US,_I3TY+>^(.H=@D,3e>YK](
5[PV-bWH\J=b(G-7@U)AB)J2X5EeSJ(L/:Y)NcJ,@..;Q/SS6>.,(.[?D6;D>2e8
((3CD6H4/EgUgC6Q#^3:UI+DC3,aO_2M816@I\5#F-GY(?SA2;CT5D3bgLCe8IU_
5F9=/OdY=8D@aW==@FGJKK:eG+g.OC(-FGdF#U2/?[RdAd;3OH^^SVI?V<U_?[W_
B#AX=f8>1V3CGaW[O10)8PRO.:TGTL,A[O9#5[\^K+R52bEEW/4IFJ6=R&7HT532
S=>^>;=g,0e3^;&f8=0SBJbA<9R\[ZAT89;b^77BbbY27T7GBWG&E@3fcWS3+K1Z
LNVFNWR3&2(.4bJB6]LT;B30^3-TF?.EA:@TaXbW-b]AA2;dD3d2Ug8)(W=X:_R)
EJ?]=W]XWA.&+FTYL><N2L^JW7]dJZ3DR3bEZ/F==T@g>KFM\,[4=A,g&deIIDD?
.>887.FXJV2LYD^_WG<H7b;/DV(4WfE5f\5@_SPFKbfP5ILXQ1Y=H\=A/[&8\V7J
E=6Q5FYaac)5)@CfEE&JL8X&gSF<4[>K7CAK6eB]fFbaW.76N[)8b^0PJ_N1/)Ra
IdSd&TL,+F-eW>:5Q247+2&HdFV\BZXC)Q8#>DcZ,H#H2\b:;)bVe,Z7WDgbM&9C
TH#AVaB,Cb.GEVb&WL>)5RI/FNf[F:->^f6B:I^G7\:4HU:)/U[e4U[b)O5.85LX
NO#H><3X\.[C>1-E]3BH@FANG++@ZU&<##ZWg0^<e#J@I)bQ[.3RN7ea8LX.VL^Y
O6BIgUX=.H.G\Nde;W=C?6\cI[DKVSQe2B]/USE71MBUaQd4;Y6WgeMg&@QdCLZE
1=MNfRK&Jb>LGg.@[##P^UQJUH<;(_Q>2;I/gIJ:DDFb4<M]V4\^f(IR(E2_AMbQ
F&+e6_eP34N:^7FW0BB_W5:(:HT[c>NM/;-]<B,1H]=0W:dA7(K,P\^X+d0_^A),
W3);##CP^>RTfZRBIUR4BHMIX(B6?&<g;YM.:.D91Z?)3GSJ9?4L:X8e4^+cMS?8
.N_UWF9-L:?)BIB6@RH\X4;4,1U:5EXfRO6Y/]\?+F<?fJ9_:I2fTOZ/=VJ=M?Ge
9WO3<@E?1:d#45;4d-?VZMPT_3Gf6SEBS.#6BgDN,<0>04M\/&KOVVSeReLV7L2e
3I<fXZ-;@2_WSV;#ANWGO&;W(P[DKTaf+[G=6<6R?1_VDW@R_:525.[-X8;7O@X3
[e\3A[Y-LP_Wg4T9W-Hb.,\UY17;aXNZWIAD=0_NZTEG87=?7&EB<f=M7/4BP21D
)MXP/d@(/[GY9PXS^.:TdB=A3a0R#OG3Jc.;R.EP3P),[YHI.CXfZM.0KTJ]7B/Y
MM6M4T>d8B==[N7/7PR1>HB^(Z5_gg_F\U5U<E]JB4JU9A1d3e/?CIRfL6-<>6S8
KHaD9>]b;-FaX?X;&4B1PD)/f:#E/7_JDFaAO8C3@/Ac5-)0N+=3&]SI\7-Y><-N
Ac2-WffBeELQd4NJC+L[G8(/TFOY4I?e)N]EOFX^)I\OD<BWP;7Q3[;f1.\Ng(TV
27Z,8[Ta5W(/>1U2Zd@D>7Je]SJaf-9JDORDSC3):^_#RAK8+&_@L.6H>,X_C&3_
0R^SV6;J9TWCY@+)ZMVbJ4&_4W[A2Qeca>=P]a\>8<BdR]2QB0N@VD;;9>7FaN>9
_=cF#_3HL:K?^R?WJc6>c<+.3])(_T3U8^J6A[g<P2_7L[EWg7?)ag-97FD34=1#
&b4@\bSQ09Q6Z@eA@/01a/FM[6C;6T6]EE]4V)I3RDX8CY1>cW-IaOY0<V:J0HLE
P#X:.U..RV)_YMMe6d7d0M_bgV94QHD?cOgGcL<CF#9ZLQ@+0M+6RF^W<\3S]<Q.
8e97-\M\aBc>KG2ab..Y(.B+N5HU^XM_?&5YKQ]?Se-;<R+IYLEfS7?F+LAg<:SF
&0?g.C58Y/RUI,fgeIfd+))Q/6ZF#0M^=_+](E+XI_aI[a#b]fBagJ+]T@HgIgg3
EZ;3V>dY)c4#(PD<8G)8(:2I3@4\9/RPGH@5BDWT:DJ8RHU\IVea0X^X8-bG8R-K
UT5U;[+Y\X7fSC(fB\]Cb7a.3=9P^6Z-/;<Oc=0;NZ.L<.;aG)FE4YUA]_RA<Q][
XP-J?]@&9,WKd=]g#E[fVJ,^ICE\Cd>A[C0(fIM61ZO7aPeWZO465?eg>0bg3cUG
=,H+T[_EEU=24@HXTS8DVe.PTKZ)(MZFdHH-DLWPJ(ITZE/b+FMNGLF)())_@a=)
5?<+0R/Y&<TJHDTWCbOPC[]++_b(68A]R9@N(I9&)]Cd#NY[FEf5B&0bRcK\E[T5
A,5gRL#=g<+PbPQTNd:B<C/(4-V[J3EMF6KE[GfLJFH[:Y1dD;6Z^[2Yf&/,RcM&
+NB,2QM/bA3\d.gJMK1J;>Lc&JXU3db<VeB_.DR^1/A;TY+FB.G\V&4U+4b2V[<J
24bZD25K^VF0SbA+Q5[D^.R;TCC?HR<(Q8QU>BH)FUF]\-/3_GO8/15HB)FF108+
5D:M;.dT,/)Q7)Yd+1CCbRD1\BR6KT5g_5NC]-FgJ=<A-c3g,3IHQ+J7eCLM,XIf
+2dBB\3(=V?AUJbV&JR4\NR2c>^fEHUL92_-If@TS:.a:_CM&cH&7MfGYaS,;9:K
1DF\+S08W73FEI9YVC>1eTd9XXI<0/OY7C.2B(_BYB/Y[1W?PK30(b/UW(XW?cEa
d&d44.7>ZYaVN@YFE7Sf00+&S_2-+MM/H]1T471@W\abTX\7Q8K/U&OVGNE4(QFL
8J?B\;Fe-W8)3LgC8CBGV1H.eTSPa6GAcK&c1^O.DMY7B&7)@_#G+gUH?1cOcCKD
\9].,MDSCRDBBOY.+0Z(=:_-YU:S37T.VcL\\@D\@Qd]L_<fa5L,d1MFGFX)6,L<
9Y9Y+&OBP_dXKXTF@#G>O#eS_,B)1:;4&=0XD]2EbeU/LNKR:I[3NP?2J#IDV^5)
>B(WMS9,Q^MTFY5E\\V^g1O&QceE^KX6K:D3-4ZQS]#?b0L@OF[UH<,fMT]B:MeU
QY.4A8Af\f7^2gI9]@P7L)&@&.Wgf=gd(@>_(EJGV8?=I?.:C,,9?Y?^8(,Jc(1Q
B@9g]gCDDBDG/VVMQSO88PW<-fONK]<L9?AAX21D<3f7f>CWTOMQWa^aDPe=7[D+
gEX>XIV5\A^K.AfPJ(PPg485CW@VEA/6L:a8SZdT[FP(YV1[+04g7JRBF#UV.V.,
9.a76\LA49.&DdZ?BgI<,Q9L&BOA^U+>L2U0e\d[FYcUB,89&,30:GK=[5g>ZX)^
4,BH8)F,<=;fPJ8)<,S#N<;2/5c;DO4<R:R.[^BX+Vbd/XD[(RBVD^Y_;@+J50@a
;cA3M(cBE/4EI6++=]8+/ZUTETbSB,XYU@L[2dBY_TAg#9X1/)L\TUD3:_WPaKGZ
:JZX.XY)cH\PY<H=PaZX9\_;J8724d,;ZeB7QXQQC&gfe=)>>d]^H@BCTe9,CHS.
;]8SMX;NS^f7K=b0PDOJG>9F^@(c_(CabaY>PS>Q0;C/[9O7@M)X&W&.HTTE1;9J
I=e-fO?cRb+&7DaI??<10E-=^ES()Sf>g@_S;4(.B<JY,f0da=6:)9O=Sc05;GE?
D-97TZ>8Yg&&1(eQK;.O;faQTY]BU\b3eCQO:HPGQJc7JEbHEDDQQ]/L22>M9Mgb
2N,K5Q/WGC.8[;g1)Qg&8QSI0,>FWU/?J^_ODTgY=,,WGD8eF(E+Q6d0TN=Ta12b
J3CXOS?VG?c_8EWMM)77.RBbaB7/Z5F1YBBNW81\?<<G?2d\#POc?@@#0#2[ETB>
+.MT,E&J#BeeaV;2WcSIG7.5==A-fe/N2^J_TK(KAC3CP2[dW)V#MSPJP?;/0efR
\8&-RSYgNU)Eg22JWEAX\M,WRc(+E#N7>1d2E(HJZ=U6/Rdg4,GN020CJbIU2(82
V&DcH)de;HC;FNYS1M05F5JQ_P9Sb0H]DfOM>9+bLfG2X+=BX01@-b[8Q/Q#,>1?
#^-Aa,,eWZ;.^TAE[\XB7)&IC/OU?gSFYaPbWDH2@_4@9e/X=?,JR>bM;+PZQFJW
GSf48P0[PNfCJJcK,,-;F/GJW7[)2^,5?28=.d<_YGYXM+PRe\067E7\\Z5a)AfP
XI\>a-DWNH6eV3aeVX59K_S?TH-,B(KV;2KX#eV;9W@;HL[GBfA4P8TJ#0K:Ja[Q
3&f:<3&-PBTdU]9[Dfe<gO;[7P6.[M1HPQZVNAL.32&Jc]6H._LU<2+1[=;])Xd6
??=Ma-[/gJ)+bV,8Y3ETMZE6SC]O8Hc,)KD]9XMT9^A.Z;E0<12+@->g)4^eS4,H
9>=Td@+20&^Q@\6R>A+^VKEVE,b32e3S;_PVe^e[Xb5O.D6&Z][PZ.5M;VbQGY>_
P8A<F\437[Z)S/(8f8K1WbdYW2WP\Q)SebX(Jeb_ecMQ\).V\1.5fg;#<XJ[IA.S
>cbLg++=;3I2b7JGJ;L2A-K/^TK+3&YZY.:5f14I,H9d.HV1H7;L[O@-ODW_FSgU
Z?<]R_9[_7B?:62/7P]a#+8^,.a)D&\@7&@1T]L#Z.AOGMBX05Og5>1:0ObYQ1f-
b:+EG4<N[;4\SG)L6,>EO&1<_Y2.ZJf#ZM775dTdID)P.3P3-6WfA;?4[[D6I#6c
4YG#21Q/a&48S>H=S9]1&VA;41/JZ5JHPb0(A64D.&FWb2E4DQNI\KIHfY\g?;4.
AK1<OPJ[9S^3>UOYKZSW.Xa>6de]-FAg;7MGbc9ICLbgADa3@-B&/?c@RZ^V4M]5
K6&/1MS)DX<(CB&0Pbd4\<b@PI\EQN:UdZK#4eTM53G-))\:<Z:&@Lb65dc-[@BE
Ma:cGcTZUZ@01#NQUS;Zg/ZXB)CE^5=@bJ+CZ4eVM[9^(_]^?,WOJV,D4gXe)Ndg
C2G_FcGTFGP(f9IOZ:]RSTUdVZIO)=I^#I0[5d\(g=+BcB1J2c-20)87JFF9FY:b
4@F:#=OEc-fCWTGb&OU?e.CcXRb/YA0Ve4YD].J@E?]/ZO_B)&61OJ8RICc;BTW]
X\,G5PJ)??4QC^S&80(&SZBd4dbH^8>\dO>&eg6dADJW.9.H-V]Xb:ERTQAY-aD#
EBFaLJDe^b5QBCf5S1Z9]eER]1>D++14/A+1]UH6CZ7^fW4@_UB;<^KLfDbUa#76
?SbH..^^(HIC=N1[?C]MJ;IF[g0,]DTKY<.L;9W>(gO/9HfO&TT>e6Q7=(_fDEeE
#N&ZdH0C,F>T6GQ>e0b0g(?a_ARIEb>e9^B:?JIPf=0>f]aJgKNTE42N4^Q8J+Wg
::d/RLJIE3^^S<G2IJ--CdK78[9+].?cP-S26R-fZM[DY:GDJ.M9GVFeDP;/(90#
.68E7;@E.(R(,]9BN8\+(15eA6O<M5+KfL):G&aY1Y;-c=/Q45XbW/<#LC+/94b:
PC[/eAU0Cbg/JYCLa-5g&BN_4?8A+WH;E4\M.<N9^cYGA)57\,?MKF\-a#AM#ZYQ
QCVf8)LCQ;6RgadUDFN/3PJ-3QKU(5deW9DFX.+bE.RCSVb]c[<?1DCfG:[8JR2a
.1Nd9UHNOG5+O2Rc)7I\Ed>L->+R\c7M?H]PY/A&bf@(d3D;.bS>?KZEA&+;Q^f=
/5g>DRb<=)8MK+?-.Oc^,9Q^]9JQF36W@HOKGWF]<::LP5[aDGO-SCKN&fWE&^G?
aH>C/,[:)#cWJ/WH?&=_6:OW0[H(__C48.NGN6a>.L9^+@VZ=^>H2&I=0A)A2>\Z
L7CNDbDc5BbSC((]<M/4&9&/\QH\UPE.44ZgIP-D2-RR]FL#UKb^WYR?BC<^<>><
4/((@-TK-Q@?2ccXc/+<\W0CXHVK#<-\#4G\e\(WZFUNYCQ2a2V5(C_Uf1GQ&dJa
S269E9SN^M+>[FQdVb&38gFST8fVYWb+VCIC7RO^2Z2GNN\.d+ND_GIJ\g:61B9[
56Z[#;dW:RPMN=ELT,&/FX5J>T==DKC4WJ]?LMP_NVJAf=bJ8CZY97dcZ\;8>M;C
2g+dHU@d?5BGL:D^N8,fg.F<L96G.MACRXb(:@.#3>NXecD19F?@K9M>SAZ,EdGP
5R?\&)15/:&&JINdI2P_C=3[Wcc#-8aKb1L6;;\V8=W_#6-\42T@[.b]&J:5.@Z5
UKWS,dOC>aK__(FB^3ZOc^T5dU\MC+GYb,0+0Gf;E14O\e]SQ(>B1a/6B<fE4&Ld
=f(?.fV&cS2&6,d+XT74UB4<If6Ia,IW_#=]7VG.R(Q//J+U1.+>JA6R(&V-\0e\
G\G@H2(]<:T9f/Hb6bBYdMg\b2c@5;F+L/TF\3XWER)O#Q.K4ZUKOV:,#;=dMaL[
N+MW2[HXg+OJc)9eEPKgD28U@PIGILfaYB4BF)FA()^:d?IRMD8fL:(g?H,FKbOA
-6=I6VN:bcM,O@[5#.+)70>EY,XR^P4O^(CXg.HV<b/D38Va#S5NfD:a6T8a3<<.
6V#I(bJZ<^dAPCeQCK=(46/^IVG3Z0aH2b+BZ/3WSRA\IBQ-5&V67aBS#)V3^cbb
;=-AW>d1bRA6TMK^P0[6G_)(;EG_;UQc+SdeY=S:SNH=2Qaa:?R^->c22#gQ]VL=
[4EF@BUL-,/GgL(_fRgGg&:L7VK=3RA\:E;8D>G4E./-O0<d(fQI</T5DcH.E_Eb
I.G[7T3UV517<GQ0<Y[R?(T_+V,Gg&bTC</f;A9L:6)IY(0.ae2\95a-,4W[D9G?
\8/@:be1b4fD,_8VW,:V__fgP]^+9LRDQ:?gG1@[?]aaR4P=ba5?-,[:ADA\+@4]
cSOX,E5NLZ04)(G9<BMe=a:JF=]18O0(3V_3DgO+c=:2-&69PL#_,>(+>4DS=2Vf
[8N(11S-XUaHBbcQcF6#L;b^](Xfg(<K4bA0bKZ^U3PH7F5&&4UG1(]N0T\d#9N(
Oe6HX(VZb7Yf7VQ(@V9Q<)C;3@&OO6\[O92A,NF#b&PQGCdZ5N]8FGU&]=5B1L#7
V/0L>W?RWT-PZ7A=FPXADOJ8.XS=J(d-]]TK)PQ3Dg7BXXd;(AKE=4\,/BePRdHE
ZG=Bb@AJLCc@Og8\F,&3IRWRC-8YS;RDb07?K\;BdIeT]/6#K2=RK.^dTDaK#CT#
11I^O4Q<;2f>BgGea_;LT5=FN9-Pg4O^:@_317FA^5;N.?;>9W[F68ObcTAC:8I@
YMB>UN,-T\-BP2=T2E28<A>HUA+_K0@S.N7aQ9CV,)e>F+0[\,O&+[L@VM+BR&(^
&:B.08NJZAODSG_?>[ggaD&=>]PS>1\+<ZG=ca2[BXg?4F<TP1>HS?[Qc4DEPL>Q
;,2D:f-E_0(dG9^Ab],^K(O91..NcYdc.dRa\<#/cH1=YE&7+Z9U@>.P+9(KR/LS
b4BF4F:47ZPC03:0^Q;g&-,BNJHF+-<cG4;@9N(^PHD2QdMM&LM^:JRILY6E0Y7b
U:K5Ud+fIR)YTL&]EU4VG(5JX6e<1CDdHa8Sf[[PaD3GbHCL\;fK+,UY/@3[KS3a
>S++g63FDaa,/:/K6C/TO..XG.1P8c[@V31:C&L,+877&W_K\?C7),-9S]-.,B,M
9ANFD0?HNOL021ZOZ9?dfL4P<ZR[DPLL2c;gf:._eY+;W#PF_I)XJ+_KD61@R=P=
VER]Q\B5S&FEBf2ANC-ICVAGYKT[c,ccL(.#ZSM6O6^Z?CeY7VD,>gEcU0MHb5@)
BES7]XXI)VNMVZN17S19DHQ+A),;@JNHd=e26c(ggYR:)R86+Fg52>5,gMg>?b/@
KV]/T^8Uf-#-Z>_&M;?R/6=&aDMMdDce;Ud[YV9+TB+7<MLRVRI-#Je(b&BRP8J3
[Q>d]f<HD?g\6Bf37=_eQL\+A5SO^<gRR+0QR)g?FT.g>Bg<a0WAYR1(&b?BI1H\
S)SSP7G4W9RTV&O9e4)9#@]@.)@?_SHe1GWU&?A3Ea7<NgVLEeP9P?V2OJU2Mb=E
/S,Tcf#U_2S9(-XG(^c_0UZ2N6A@ZMQMI]P3;IYeBb6\?([3+T2:gC-DEEJ=d1QN
gD=W/0e)3KV;#eIEWYVf[EfTD]<fKNU-U;TI+(6&BfgYZPR=BHT5VW]9K\BgCZLY
GO?_Q#O1S)Cae_PC\I6R+BGf1CWbc?+EZ5#0L828R+:McGcP68H_bXae>a^]KHL]
GdP).Q&>AT56A>9XC]JY,N1egC8.<WQIVA2A5=HMb4C=0:d2@3W6L8:T48e)4Ve<
7^bFP8U<S687OL]=KTSFLIR=5c489Z7aV9+,9.5JQNO@=/d[TN+L?S)T\/SXb&>=
X3JJ]-S_T^#DdHb44;?V98XR;#\/gDB8K0PL(AADgRU-:>Wf:I;5AeGD&M\NQ5U.
??KOed>J;\QRd8:;QIR8><_Ubdg<:UBf><,ZWF9>-?M/G+EC5SNIN)2@I@<J426T
gK&,7-6PXCgL)Mb29f>>6d8GFDUId0DPGZ_35RB4>U[@BeJ?CC&[S&3Q1DN2++OX
UU_.S&#20;g-]+YUNJB;0[3]L<D+/#e;O3fC\a&C6bCg_g#/R\Md_(E6[YQ_?Uef
8J_9>G6UgV.aR0eX2OP,.+:^DgWHcZdg-CQ9V?6]K[MW]g)2IZCJT;GFX(-]gJ)f
+b1ECC9(cUd1C#&I>-CZ)9_U_@?L4aS5_7@WD6_2&;+NaV?e.,B,]F]aJ256@N+)
.fI.H-#@>T<?0acIb8]K,<&.8JIT1g+Q>EKL[=AeD;]IcE0^>gHOgV#9=(?,)1LU
YH>5>dfZeVA.ERMF7;:3W;IB;6D=C>^>1PAGe@T>D7:8fC:]I4CG(_7^O\_.UURO
@2L<7[W(]H10^ec(ZOFaA@K(YBF07EINeYe2^VC<D<R^JGEQ0E0Y49eX]9+;/2,C
,SeX4SS]<1-R565B\-DYcP0KVWL.2E2dC/09Y]9#ZG+[3=QeZN0KR8XeG@fI9;Y&
21?9Y3N2CVNOa+2NOZ&.CO(P>:K[O8X=f^;HLbT]RD@6]^JA\1NC:7?PC2R0MeE2
./<73MAS^RJ[ZY-:ER(R1I+Zf?Y6A2aM[33JH6E,cD,V7Ce[d=]4JKV<XJ=GK6M6
5Z&VTeW5OWVHgF,54<,]558^e(/>BfGKEGI&WS<^CQ##HS2,+3Q^F-O3/(_<2LZW
=JeSX(c;B9d7b#Y+bPBMbO;PbGbIDIF,G?-^M5T9Xb(__CEf:3#)4Z+.Ba:KEKTa
:+DfK+]],O#YRC\_LbV?PM;,PSQ;Y/+^M&PD8,gV_2Z>gb6?aE>;b92GBb?C/-=&
<PTY0(d/:KY)b/T<Q8]6BDXaC[X?#d:[+T<L/53>+>8RJ?Ze:TJ=f>F@E6.R^3NY
<.SSH+JRbK2Z2YJ_BH77QV3GEX,/ObDL<AQ6IgB(6I,Z-Fg?/R,.2c:\M_3EC5XH
]DRE[>@TBXK,=bBUN53L^CNP49Kd=cdX>fE1]1#eMUc>+9L>0\e4P5fWdW#Y#P@,
3aS3P0K#UFb5S;9)P[dJ[L=<N&57?3^XVd1V&O5YAbCfU:FPQX64FR;Vdg404<AH
TeBDGNLU(>P^D.WM53D_=/UU\-B9QA??0,.:6)9.;Z7-AU#Q1NHe7f\EQZ91++T.
,)30L4cIJa<6]0UM83:3-1@cGP,HKO0[Jaf\<Z;Q58T>6(3IRZQ4K_LNY\[Y5?ON
X18=-JTT+(D;WF7EL2eZ4<(@KBIWUHdBK>NAc)ZM>;g5/P]6G5dDV]7f_9X1T;WK
TF,D)0;dR2D-)7CTW=,40P@gP;<#K/dN;0:3FZ4UG7I70M:Q:#J)D9I3[+TT[XV&
c:W65A3=?M3TC^_)OV-Y^/W](fP5f@0V1g<@M+UG+E4OW.#0SSFLPOGI3DAc@D4<
aH#NAR7Z6N&-aJ(6Y>cCVD^fQ27,@=9bXAX([f00>K_7N5E530KYTB+>][<0?60Y
Da].^0OR8f<_EgZfOQe,F-Ob5ETA<;URN7FAMK#8M[..(]gZ;BQ82IWeF#USJD8G
7-TXH,AUX>#Q/#]3(WUNEQ7e#8e.O4WM-+3G/J#P/ZOWf@ZG:5.9\3;X95XZ7#7G
Q+a?2+L=:29<3]Q</C=44Wg^g;FH?X2P3\&Z&QDQV/A:VG91#O3^Jb=4II0cYBJR
?/Q1+X>)a^>HW/TV9OQ(,.:NJS#H&:=&?0TMZc?3?aXe^3=XWDfN0?BfBN[d>J&J
U;Y0=8]_?IAA#S<VO@g04.<4TAHGNA5:g,6FG^Q,QE,ZLVPN=9cR2S,&RgSA^OB:
<LK4NfR(B29bW3YSPVa?.R3:aRYU+X?_O[J8TDd_J;>U4.&M;DKdX-@0DU<b2QT:
2.=Yd+c:_##WbacDE2@FV++J_E]IU\=4=<N<+CY:C?^ZU0[WU^4+cLT4c\Qec,EJ
g1.NF+0<:IGdeRSDMa(>DeB99)RG^6<VXg4+b8FM)ZCHC,O?Hf8-MR+B-WC_U)J=
+a-4DfdN)IdIX^@(K(.d.4+fI,?:S;Ub@NQ4b?gL.I9&YUc&)ge]@ZIWT@-<<GQX
YK7>ecE9I+_VJS+<;6EA3/(LgV1+Y&,>I<<_VKG#EWBR_Y8^PgQOK;a-GH_L,(1-
A7;gLL\M>c6/O+5>0K3QBX7DQINND3XY\8Sf?BUX#7A.15#4d00^;Ja3G/R@dO+/
Q(@-00_5YYC[(^XWA[PGD26bQ8OO7IcUTYfc1DF8;T6K[K[X,M]9a<IQ8J<=f1a+
)(.K@.0:\P>a&@GG5_U0W7CJ27gWaLEPY&T&)1E=(6F;P_(NIL2,a0C].FIL)Rg5
c4DfB#EfY<#<O3[TS:DNbc?4>5g5V(-3Ra:.<XNVOf#3H>bK(/gEL4V8-N-KbAc[
dZ^,;DS3>OgV#_)K>b(WH?KL9/Q1,3S)76(:T&IeHZ\-)K=01EKbbS5OWBN/_a_M
D7f:GY_+OCQdR5?JYRc)-7/YGRU_S#E^:VM/bKCS[;T;_5(cZ#,1dHJE61@@</3A
A:U4GMZ&=AZ]D<PA;/J&@V1N3^32a75#[/H6UY_K__<;HBL;EfZL=]?H>GSF#4M\
OeL/+CSI3J(/J7M+X<WbG,KP4Ic@=L.U.0/e,&[Sg/80C@&3TU6PO.:fg=d_]&#A
ab;[fEB&>75a#V[5fQXD9Gg:&YDe,E,.c?P@d[7XR64:I-T/bG1bING-^^A(^(@d
5SR7BE,)JJ0.dTRJ-N[#g7I.O-EDF=__&NecHCS3-R;^^3,f\KJ2LB.AU]&4@<3&
#]d#aMS>MI?9-:?:U-HDLJ6J4WP.&E=DdbP#=B,@\\I>E63Y:X,C=e_]RQ4=@X.0
\XGS;ZdJO-_:>F,CG1-XBL/FZO=WF]QZ5#=J8/G\54IX.IdF@9;.Qf4K#I/TZ[A7
HdWOOgVgN^8VDa6Z^cJUSIHJ)D<f<O(ce/UF7I(Q?F#D@EU0EKI>ffQ\dUFB25XS
<XU@<MQ3][(Z0/M2ag+\F5P=FP0E8-5)?UFR=(L-CEWOg>0CD6[MabYKQQa6<;;K
?P#N[Be9UgPT0:\M9R?-S?UZgE:W.9fY;+BD^[g.Ud3X<e/(e8^;K.52?>TdW/H7
:G_;QHBGIC00B=LdgS325U;0^RC6<,_cR4VG>CNeS,MEW1bJFe(&]8abENL_Mb@9
\a95f=Bb]?Xb9HF\>HIcHD<1?;H@69@bZE(=8g8@N?VZ9db>F]K_JQV+LX(H:(&U
<T42Z1FWB@9B[19Pe=KNR[c-QIg<<]VSa]4W^2,UJgZX/Wf9d\U?^#NGFMYKO=9Q
cPGe@@6IYe=Gc+.TKd7UG04Cf,,5T.<Y0U(A\5L+_>@XBVQFfU+<7JZGFc>e8C;H
73+,B/S1aYKNXgEIK9.U]#QPe+W.O1+8]&A)/eX-;B2+[IB#dPODZG>T^O,-+.=\
gc.eG#WXA+4g02<1/a9[^_0T43&9LXg9Z\=8F#daQUM++20L43_A;FW^e#<R]E7C
7,U5B>OOYODgEFVW></HW?_)@Pb4^Ec9dDYbJfdAQ5WS7+Y.;\aD0DQ.+Ub5M_:a
WNA(f.-aZ#fV-XJf3^6Y?<B,+61\e9O>/P[g]?b)4]+<(DBR>R_&]YO)N9\<C]G>
6aL[.U[K;=,GA31B^=#0\@A-+N/?/)2FF&@^<8QG@[DOQ&[4\?-)(3MaJ(]]f[b1
/IK=T5eBV.;Q04G[9W_EA7?#/K9a4-P@TP/11<@20=6ad;#DA[/\fCAX&_+4R?N;
]D25#.H5E8+QWN_bF#]<Mba?(#RYabV5<>>-?TaaMWX[_ML4>>BQ;MS9+&&F;]<Q
B13]YZPWA.F:=eVU&DFgf]G@P+@C[gc)fOY9YdT8gI=JR^SXGIS:Y^<1C:GNX#d(
1M?B1^1ONW4MPbW.@DeFW0Jf[H6f&fD0#JA2LB.:W6.K0TDA^(@1F1CTA55]HV[Y
\@8/#3K@GSMM.D#c=M,fADWa^X.Q>4N3&L/A4L:DHLC:@:()#HP\#Db-TK11KJK7
D-KgU26aP6<#NfFbDZgEPCR&(=Og,XY=AM8E#d(bVL:864HAG#F9d:eKJ&c]_ge;
M1-LN8MYG&9A_D]KFLb.I=RPRd<HLC/K0L;+eB;5CV5YTWgD/IX]0YKC7<g1^4ME
<GIEb=B_(#:8b9gf]&ES[CNVG:#\8Q\#Cg_MecJ]39OJ)/FcGCYKGR^GMfF#Z=WL
87daA4JEK-[7FZ+\b#gW^=#KVAf+g2V)Q&()@\1=bMM&7N(4)e,,cG\=b]V9:Y.#
\Y,cGcE#R>M)DZMf0,dK203eZ#090Q4_g\Fb+ZP^dKT@bH62-CG4HC#U)>6H2]?G
)GY/0(d^UHIKb95@dLaN<97:;+/L?(^a8[@3C_HM91WcF<XD&^Z/R3?(,6NR]X5=
G94Ka=I(XbNOBBJ4c<+65A6UcX=AZ/)+e2M-\VVf/@?Z4S@M;-.#@PgDO1_8Z=c9
F?ZBa5](E<1#eF79VL,T/M6D.7f-a26O-Z/e5bUY0U+<15cU=W;S)F9:#71ILR/0
_,a1>N]g,&T#HHNC6^dS?F9N&c[@01KfO+DW)4E,^Cg\G-]E,S:D4>TWL2EFbf&:
;?W6]YT1G9-@:B3(HTX)7f=IHTB\1,5MYQP@&(C3:AdDU[&\RdB0=FL3O.TfdN8>
g&&G)6AdIbHNS/GXdZYd1SNQAP2&33T1=d7Z[16S&-@adN<;CFDS[=HO,+D+.#WX
.5G3VLR7^;V<a\_MfaeKTGKLJ?ZfS.:fb)G\G#)]O/4P>fg^fXE?eL3EYEe9[7TM
B]EQ5R2(=).SM+T1[HG02)L4cH_gOGg^a46bT/HSM36Q4f.[JOMWa\,GV^XYK7ZD
G4#,IM=Q/EBJ.UKgZ_3^,g<H&b2B]bT5<X;?-Z;6M>6efK:\D_MZ:=cY4R=^4<,T
2,(d/c5e#-bVQBSI(07K#V(\L5H<ea5gd?=7GEW(L+3LFYDEXe8FW6[PN0;3ff>H
MQQ+(I-[;ZJWLD4=:K,GKA&aQ<^\e]eW&=@\cM_/>Be2-,BKZ)E0]I+:6HaX9^c0
L?ME=\YU@55Y@(#2G?<[=S+QGOFIg8C8WRT+g+=YB3[eaJBEL#)4Y8A4D3UUUOeK
,N9e0B4fTL?e:KcM2JE;13&b9aEEddS23F@S1AODCX&183g7&K2#.<TC3KZI.WOd
3c;BS0_Bg)EI1]CT<g&MHXUfY8Y:ed&,HHBC^,g2d,c)D(M1b7CS/(J0g,H,;_ed
JPN^=YZZL<6e0YS-YITQHKeX)J-c#24Ca>/=A.5@5>1EDW>CHRWD.Pa/@d9DP7T/
gab^_6@.@SJ:B+8+E;#QLP[#X\?5d&9_BXHN2Bg@RC)02UHaFW@TM8e:Z+UO==91
.2^7WAU0QaP\TZ]>2(G+&7f0#+_(BMD&F<S0O\-JU_:0VH:.OFD8RM-R[B5GGGSL
D^.Gc>SM,^\>0/.=94EOb^S^4Bb<HA]U-GTGJ<_YRIaada@D\?.Y8,Fd@UDeOCP_
)8O]Y&S,9c]\De&8^(JU9Ia/5e3+_H_-fNBLP@E85H#7D:X^?0cUD(LB<(K]1&7Y
BOZ#cG?Z@C(<V>[([O04],<?FdX>Q\OFUZ+R:&TB4FB]ET#41<a:&3LY\L-SUc<a
DB:++<-:)K<4>&5\,HT0,GK6]NQf-_(dK>YH9X&&X;8-.GaD/2JYEYRBEYO>O690
I/7GZ8(0gBdP?GO;:L<G?6[[QZHM_CSR#EWML9)/]1RE=_0>P@+C:]P/Gcaa.KN,
6.fNS4DRYANV9\0J4)&A&4d71e+Fg?4=ET<fgOf&3@1O6aOWe_)IaU[XS(WLdVWW
1XU,XadP>^_cP72LC>P)8SCRbLY\U[03Ped;aX5GPC?ACeKg(PX),WW?X@T=a1JS
K4UV:.^ITQc1.MC1ad,NZ33?COQP:71&f\GG<E=BATW\2\X,a?;2<TE4a5#JBSX7
3E&V=0:ET##a+a?-OCGD9NTY;/UGL]=eA@Wda;>Z9@FDKNeA:)Q?3ZQ56Ba\DVF#
9ZfAS]:#Oe1gKXd4=.@VTa8b0J_B=@/\MQVE5KC_\9.?UJSNQC/76N^8=]&]gbVO
/D6?G]EZGZQXZ33fPa:U\DX=T@f@GPcK<G13.\dW?L5_a5VO#<f#K8AT:VffXeUK
dfQ(gTd5]XBJQJaS-dY4d+:6KES<1FaOY<a=a^.ED+BgA5c>Y2-P[G0Ka;(/d64O
A3GL0_d:+\B7R#J]aO/5#)EZfZHM:0=HAR\O1AC4C\b1C7+GM.DP7>6J-HWgcY^W
gdB&9dDX5HNJ+,],R9Rb/aOg^<L\RFUCFTG@ILZ7U.9^W-e699<AGfbPa;#DgD[F
I1]?1ZeGeaD&]FI)GRF8D1?f-4\-/7\2=RYU(F1GN;4,>72Y_9DReSAVL@gP4g31
YXZE6?7+-]-fY4)\dEH1S<c\4V=I_M<YbA5V4\O;Egf(#[I336Sae[gS/S<TFTd.
0&6K+YPFg8TU<6ZDVgcMWXR,T>WW\0HLZ[^L&&N.C&1<g1a1GeQ6?F^4M&2]fNJ9
L9b+86N_HF?2COTdPE#U:N?B:HE=/YTYHPY9@9,XeP#)X+:;fM<,_(#JY6<^WGIY
S1ePBMg#>fKJ??Oc7B(7=70d4Hd)G>]J@D_KA1@XZC1g@XKG9bKN#&A732&C]0(.
GHdJVXca&WA?gM::P-5Uc9g]Q:7Ka(S&5^H58?C2WXFgcPZM)CG@1-aU;K4JQ)E2
?XY,W@66]f\5Yf>8d=(Y5R6R90P-PSW5Xf-XKA=>.SL;UG4f97(84Zb2IWCG-F)4
e8TBGA@,<6Dg;=1&&IF#1XY_Q:X=_D]FC]-J\2YW0D9f[?NXA57;3P+.<7c/06_7
228C)J3PD(?:_A;ebTSANe.[G/ZRA3V4H)^d)@S8cG;Y<GA[K5fFa+?RR;GVE3:_
+dZag44^Y71C.LOMOHEK:g[Ca2_U;Y)93N(f7_PNF;?TT8P2Qb4#PVGg[536a2W^
QSbZV>aF9&G@,V&G(N4.OJ_<K@,E\?Dd?<6H()RK;\#:O2fB_9ObGB(_#N)SMJ9K
aN+b]fIQD+1OZc0O9K3RSZ0F)N</GBOSZ.<O=5HG?:TEPDW?<_W&+95YLU3FA[Ob
YC3Yaa4R);;JS8]E9Z@7WH4()Y+;GK\D,c+3R@Nd=UDJ:/@JQG@ZC#QDg?4KPQ[f
IfC\<ga)WJ[&H?b&AD(cObU-K^?[g0b35T[4g^C<d0111bZL/=<E\C^fS0e^c@B8
Y=B+HJ4:71ae]Mb?HggI>QJeb(<447b_[95S_-UZc,?L]/B7C=a;385]Dg2,<_.^
>bT[MR,/gdK#IaKG?/c6^U1Q,c(Q(eJF(Qe1NKO[<<CTfGaI@+[^dFQdOU(4aBWK
8)93fJ1@fa_U-V-?5:1=Ug+48,a50MK7C&PBggg[)RU.5/?1[EC?2SG6g40;R\T>
UCQGH9JIQ[W<_;CO>8ZCO,OQ=A;f86e8dHR]3&bZ\C^PD0X\aL,Lf-_a#17_e]@_
cfUa9SF5INOG,),N?H7g7fK&(/8@AU-C5^40Q0<R=f@XB+#A27YI;-gX=9QFZELT
Ed7\[+4S^<>T,;:g@L,PP(Z^1=^1]Cd)K/M/=1X(M^e5[a4(13<GfZQ]fN;]C1dR
_L&P.9A#O^GJ]bdAS:/3.6?U>VL\QX\3fgZa)OBZ9f<d#_G2;^7UW4+7X_M-UN[X
HWgUXSJYFR>=U2]JHICA8(L6U3>A1664c99+2=LX3dV;#I8#P4Q1W>8[AXd<8P2A
SS_&<2CN>c1K7aGR;-01KOV?[)W7fS#W&SD^PR76f_7>a/#,A5NFIa6D9,9g5Z>&
PV0-O@.UIVgPFT(FU5)]P.PP7MELM]#;:4cEba(:2_B\4QXKCJ1<^VS-TcMg^7XZ
@d^\>AYf:f(YUQQ^:NaHL<0TRI64>bF+a-)6+SM0>ZV,R9.ZeSQ(FOQ;[0WOR_ee
G0/aDB8WB^^P.>_KI-C@<DJD)_G.0g,X9V8;T;:De/]19,(e7<9//?f9JBPW]U#f
V;5?@3Xb5fVUH6GJ=Ef5Y=AVU+>K\4XYdGBDGf)0S]V&81ZXNaSOKB4C;N7^CEaa
9-WF:Wc&LfaR+RDc;1HY&f@&MBIT#d<a;BHOOY1T>@bB11aZ)b1</&6)J&U&WNdL
3=c)d;;F_>CJ0KY?\[PIIY9.EDAcXLU4-4QOb5:1c;#b]:IQC0=6^K]a@7/KG2#I
14(6&=3&T+]g8RbL()4UH/1TR&CFF;[cNLK3V-g+8Q>Zc9RAdPQ1=N6]=89\DL2\
-MS/U):4B<_@4C(8#BS9-F,3M:bCPN<29[,KO)F:c1^L+-[MDT#VN@++fDBVaIVT
T,>G(2ND=V/6]/M#U>CGa(?f@b2/X^?E[Q?\T12bJYMQ9)ZLT3CJbI@P66P^O)KF
\4A9I7d;]=[KB4bER78f8)E2E9YN@DJEb7>fU-Fg#bD6[Q/8,gMd[K[3.Q<.J#:V
O&6Da(cSYV.YAb:&(&2J:;^FZ>U#[37[gBRL:U#D#PKY=BMEQ&]38V:J8F\1I-a^
0_\6.KWN[UZKAJRXbDd/>PBX0Ee2AZY.af]4M#KF:<>/eD55eV01G=Yf>1PMZ&U,
M-,1a>5_04f51DHN#/DW+)#,YAddTb9EP[Of7RGR9\W[d/eUgI:eUJf:EWPT\7@&
fE<R2a+GD?+6/be8J6d@^Eg]1J19#I>L+Tg-TZ.;>2d-EHH);>)<D(DagUYFK_M-
@1#05DK>,^<EFMLB[AdgBB.]>/A,W?:a=-aNO8)5fG^X91#5cSB/=QLE51a_Y8/d
@-37?Z=4X9Y+c4ZSeB#_M2H&gDd[\^7,1A9..7>(IJ=)9@K\Z/-?AO\c&V0LGPNZ
K57FRQ[Z-2E\/0IgTY;.K&2X,d3SZH+11F,(M^8>A4]Ig7Ca\B(gfBT5QdN:A,,F
R::V.g+8[(][EbJ]7I(CIL2gaD@C0;@DG/,^cN0ffaN]-^?A\F@>)<d(@_dMZTd(
/<MB^V((()H\B:7VVLb0S9dK]VeL)b/?+PXEJN?X03H>&&.F7XV_#LERE9GVBA7g
INDB?ZH/T@=+5]]E^2W?5WGMS.(HaDW7B7@5G)cYW<OAIP6X,3(2?;7B=WE,E@)>
R4,M8(b=60Z]a?)&DWNDD+\VNW/4/\LO8O;[?>]YY.(TK2YZJ,EH#TVY>[+Jc/Y_
O&44]&]G9HI/P_b(7P&T,D8<QdPWOYPg[W0W].Zf>T6WGLcUI.(;2,W+V9/47.fP
1d>f)_=+2/3/>TLC:E[=Xe5#J@6D)&<OJ^ZB=YN3)#F=I)K,d&5U.2C<Y[a#1CCW
>)AG08CFF;d4=?I<WZIMUIVGSd^-dKSZ83C=]+EC^?>P;6XYYS)K5PXRPZ@]1N0:
BN?QGE4A&?G2&c5^&1>8.g?IPWE_UA\.f(&[9E2Wa[CR\+2N[QS<M0P>/ef,AI=(
HBB95Z<ITDgDXeV[>/Z4X?SF]1V/cLeQI2;1BNJ/JCPI+DQWdA:G&D4+?Y7bV^.Y
BG)(KL-B7K\GaJ=]Z<O=fKBQ;?@g#S5#CQ-.<cTMZS4J,Dd\d(&2X(>>R/dHOS\K
&DVYMYBK.:65CX(?I#-X@LUfRWOY>KF2^>.:IM=c3_.L2dL;>(g[K]d8P>AI5gE4
UU+U^1WMY8C5+\,5=N@A-A-4^ORD_N>7@b98N_K]B:g&WgN3XOU]@RXa6e_Z4-)R
R6:XE22+68S^&XCQMfRL;2T0PbE\02I3HOca.Z(WB[6Nc6N#Y&KKO:1beL@L?]Me
_AWQ)ES8HaZ)V;\?8UJCYgI/:TI[1=YAF1YTJ3I3RaJg]-F8ZZ<_J9TS0[SC1]-[
;93,+U[f/XS_FT?>58>@T^1F@B&f3>XF^/Td)?/C,TL_aKRSH2^[SS4[C,7Ee-;/
g?[XDC5g<FdVQAFJ-BU-UKWX<cL&ddKL7/@-63Q6\J?67V9a)gD@:@C]H<D_\c=Y
O58[;R3E\S+@EG)Z6&VP#,bIO9T-C/a=6TX0[#2;a:^ZDSZ^B31Zb?b>6]9Q0^C?
UbY>H_(#-;_/B((2>@c(eW=9?<ePP2^_ZJ&N))ZEE7=\-+U+ED;R7f9[AQ8gJT7K
I/7I[;>(K]4B5,TNW;@M+9^@LOQ/G6:73<7c/0VF;dVK\1[)58GRN=:>,U#ZT)Tf
HGSKE=VfgAZW@#JTO8[?+U1(8<^E08MGaf<IbPOfYdVg)]8),c;:<a5SKM)G&[bC
1?DPJ?YH5#:GP:<8\YH:&.MD&\M;,Ic;B<#M)B^E^&3).WY8G<^]RO7NDLWXD2@Y
Q=,b(2#,]2^UcC](E,<Q[I_28XG.=^c.HRI6N.QfCJ/9d_P:OJ.e>R+b7J+-?E4+
Q/N7=K3_9#UZLT)+V[_H@=&O)ZK&C])O?KRDHEZ2:5&-UW22P=<#^=FX/.?RIDGV
NDQO:ZF+c.Z4a]ZYa)G?dX)&b&KE@U]N8DFD;ZOQ9O1>EOLg46<N/)P_A14\NT\Z
NL[2QBE_U:MbX)Q4QMCU,A@AAVJVf7VR]?5^_5-1<(9)HWQ8TfJWcB;7ef,\b?&S
]>-PI^^@)18K+M-PH(<]g4cgc:d5+JJ9^/D_855LEbSV&d?d1,C)XW5dC>>9JZ<H
Z&fCf](8Ob6;303X(@]SI/D,\N5L4B7AZBGZ4;Pe\GE@?FE>W(.eZSgMD#=a\;E@
cUD[8XXYYDE&BRcbHC0,OZVZ.JRgdN)(7baCHHT^K2&fR(7XRL).>SDBR:JM<FUX
07NZDJCT[+3R,@PYQaa8:;\#F5:IM7c,d6U0@C+M5;P/(10YYbN&IIZ?NH.X&cT@
LF?g)7WaYI\\(K_+P3f;Y5BHcb#0^Pa]-X<_>[4=]TR.cI8OHc=a3ec]f:70-g0?
Od2BEg(YJ,D4GP.dVb[O8Nb40.#B<f1IBG4O6&C7VC&6G@UDZPc99<dJ,)c_^@[b
2A=L,[K-WQ4C8b]H,B<CZ[;0N:Q621&1:\:9\I^)G=4M&><J21DE5T(SD=V^,&Ne
ef/]\PCg4YH6<9XbH14g@I6ON4)Q&S8Qg<fD=S6&-S1#daJ>2T1_:JaD0,f[NWL)
MN@1G-P-ID=AI>3e99>Nfe&?R(5=Z;1O[Kb&VcHF8fH4#cYK;K8][;@f=]2074aT
<RA/@.Q0BJ@&DO6([<RaA4\,Q^G.?Nc(JT9G3XEDU[6#6WON^]1\D<Qa7Y:YD9e+
cR;RQ[RQ#>c?=#?G.IA-Q@9.XW/Q:.2\KA)4E;YS@AS4A[&]<D34-d;?V0ga&S14
/W(E[)a[.9V^,bVf^>XZWR2+65/7TMTHcQ\SB)0[AHN5T64<:_G4;FSII@Uac/?E
7dBRK&VKVFSQ1;K.e09PWM#Cg7,&._^PFEAd?[/&&37-aO:U:X,d3.OTgQ[@V&7L
I<(3_SNIaaQ[?8_]Y,Y0J,]TQC2R\RSKR4&4d7]eA[2^@eAQ#1WT,6bM.;LL<,d+
8_d@cV^SH@?)Xgg,DZBA^G>V7@4CRb]W/f@&G-40W^e91:7gI4/Q//0(+,@G-Sc:
e.#4/\NQG6.+7WKecF[+6Eb@RI4F?\.A0SD^U&Xf(T\)A2I,=dI_JJDH34,VK5Lb
aYEK3M8T]/0.gOP/b77RHV/dcM\bB3eQ9Kf1;[/<+J_TIZa^>=b_18/3)37L2_A2
=]<f<=X07Qf1]RNXW,DP5Ug1[W)8RB>#T_,#\WGd[d14)06[5R;DN./O^2JF6P^A
W.JU[H6:T15IGBL,N#RTY+LNK/MG_(+6D0\,+gVY)=8\@X>E5JVaGVfAfVF=[c#?
KE7V,\KJXVd]dUU]]MC&H+=F<M4TZAPFSP>EVCd=CBD[2U)X2a[a0-E/QML=<V41
7UW63f#V-.Sa)1-Id[Sg(_Y\Z&E;N(B.0)95E5=:_[Z0K7[IAX@1OPbdf=[I0+KO
(N/Y6gfL_345a(89b>6+-A)Td5Z[AY@1;G-E[,H1SOX^(\&dKH=/ecN60C8GfH-A
R>Q01W3?MV1Jf<QT<-cP>,GJMP=aG&Q)3-T+g92]W_g8(EgRP?ccHY4BG\:J3d^>
&5eQ6U;50B^EWa=KD@X]5+[VN5WA<WT:6RI4J.;M.XT&VE0=Z4Zb4;8Ia-+4IH0-
0^YVH33<LZ+8+)DK_5G3X4;IG4VB>7]WOIF8T+e2e>dK5D4@T6CbO<Qg7?&LaQ&,
I4H;eAPN1aU)fD8Pg6KSX?,LJJ/.c&USW-J&X.)GC2feSL@M8Eb=dIDf&1.-)g;4
>LAAJ_HfV-KC+6UaaZQgc2(FX?X^3+U19#:ICcd#O<S+c9>/(=HJ^[N^IF5OJHc9
-XX#4/:b/ZIT1dN>ENGLY\^_1NXBL5,XA&98KUOScIc5(aT=-?(ICD&F?JXPfUEA
WFd9>IGWeX,_2cCC?JDDPT<AR._//659L90OL]-gF8_B5gF<L\fSS:_48f)5HBgZ
D>7F,]AJ-&_]59TMQ.7NLLFQ3J(4L/4C;P03:E339DZb@J<=OQZa_N9O.7-YPcV\
F8TVXPBF#;B(aDR_N?U_^JeJOCc#=HWR/B[R5636Ie8BMUC1F\(aZ(G/ffKZ#19F
;WR<bEOAaYfcS31d[AN5[[\(1HZQNVOMP+dK0367OY8DZHd.b/@NGG2G0S@aN.P0
.eP=)bQ@GO^VTAQQGaW_NaZPdbb+CL&\QQ[b&eR#6EMfV3]?XK=FMbW,#f;4DJWc
>C2e\-2/A7d+Q.:L]YE6+>2>-IMK@#L\4;:5T>[\dFF656,5IKQRI<QeY,WR6Q62
-&-EPW-\#b5>&eYEY1VR29WYC=3>6IA4-5J;Kf-&<NQT[>Xg2dO#V,(GA\NAP5d9
-IW+c@6FD]M^2C12D?OcAg02+YV@QIIa<9;\3P6T0W2G<C,:+^EJ2DXH33RRD^JE
-eVMIV\FNAZ9c/Q1[KeRSZ9/f1YQ8:Y@6KUNH-^E:0/F>L=:GI;LD#-c(&/[YJ0<
V4ZGC&dYM^^g;(3>4aQD^dV(g&c:/6-;0[ND[H\[:S+/^CKHV#MHGg_TG]\M5)_1
eUH<Jeg,gM(--D(?eg\S-AaMW25>0=HRgEN4TFA=IYW+1cFT@VbDVY/,,H6eNA\?
?4Cb01Y&(7Z94M]TcD.AUV6aaW^CZ4FP\f.ARg0G5aP:_:O?+Q:[DQbB,B?W:W.]
SP2/[67IA.eG(P]g8Jc/D[+1fL@-a<C_9W_@T>3=L&b[N2>0?KI+FSeHR_^WeJfQ
MTN5C&,D&TLBa#[\;Z?D4gEK;M]56QIe[b&K?L0]D(02BI<WMF^S7I\ed?F7C:DA
T,B1J2J-E(DWE-1NQAJV1(V66NaF.PdEAg,3Z7c5J]T&Za9G\#Db>NOIMH@4@E.1
a>?Z&c#&)LQSF1T\d<F:][#S8CESYJD3OgF;YK7A[/,<_=P&P4EDDg@e_K2W7:QE
]]L/P@H6(][9E<@\XfMY]_&?^=O3G@,O&\,.L+.]Ga\VFYWXV8_GOQ+(CY\[9g8C
,>ASQcB<?-,THE1d^TOPQ;DJ]DN#YCSS6/3d5>.M@,NT-?N/;6&(4RFF)K+=@;f(
aJA/0C<KWS\ED#4Wg);Kb44\5-H7+)[g9E=KQ8^TYX3;f8<c2G_@MK1T[&:0C5C(
(IZY6,LM^.a\,c>/AAHMJ-4=-&Y7\)7]ALA?_e)fLQ;YSQO2bZ0>ESbV:QJ;CX8H
3E#)5H4de2R1-QF_:5)OHD9fK3\10@3?LTR7QGfFfU8b6#==,6ERg98dT)f<f(?a
bR6bWXI37S4Q/I(:99NRB>I?FILLZ[LQPS/N)V>?DU\-R8M[N2V9_=<1472NIWN(
M-2BgH&,D@e\,0T)38JI^9+\:4/Me7dR\S1K4M&.^PScd56C&^?09,GgR_)8UONV
R[/N:DI2d6Q:)J=@BX6=+&93VH</+A6EW03beP3JXX]+6e5U#EgGb1&Ca=R[X8Pe
G<3<_[<&SNGSR3X)F:EX0H.V5:KTMe((Ic9gFQ4(>eX9U1EX3LUJ]#cIZ_.G3PNZ
3F&2JU?abT.63A46B(&8N:,Z(O576+_f51,b_1gKKCY&<^8VL]>AUBF;)^/L4Y@A
4[-AV=K>ZD#f+E/fMX2PY=bSF[bBC6S:QGgGB=UW;3-[/Jf+R=?TB)K=)GB4dG:Z
5V(AXYKEMG9=aS)R.GEKZW?O_B?,4SY(D3&B=4KM854V;_BO;H-INCXad.HJ?b>&
FVN&NLY6\B-KcAbR2BK8O_EV7U;++6W=P.]&(QaMA+=]^,9a)Fc&RU:f,U1J)P85
WY68<C(-TY+M357LE\S\>/FJSG5F4KT)G=PMYYM,ERRZ^0W)Z;[:I>g0CR.NgE(I
X<ZXWSP;=1SX^?4M7caJJ41]^MR=+JDU+]c.g55-L#2=H;bce?6J6YH&?F4A5AgS
-5M8V6O&Z(f2RZDB[eN]1RK[ZJ>/\+Z,/g)8E<Q1K41@a-1,LKI/;dCa0dI+;-:&
RFMYR1Z1/47Q/#S,cf_7@)/F9F.>cMe&BKFL93_5aXW#)3B.4WTEagI]#NY4EBY;
/86D66fU/])PCLFMfQ#=5A0:2VM>Lg@5Y&bAe,16GMcH@(I3,?2Q\=Uc&)Ra6FV)
0a0<=W;2]0JbX=2Q1UW0U;E11&^6/T[)O6;JT_.\1J0Sg.;&\,>OQOO[>\ZUA.>C
4,d-NQSH.+1@S?eIOO8C:LY,ePB5e_7NUI=XQ23WU(<c7cLGaINZ&&3Q\H<H^<NQ
g</^Ka_&P(KM6XV40IaU(K6BaF[g>[FC&OSZ6P3-L2+W1PVA#6cST,P?c34LKUP\
:=BVRK^bE)</7SR]eT30WE;D2FSg^FU00=SV6RVOMdHFSX0;T<T+OAVb2[D;(f<A
c/@3,+1Q>f<X6X-2A);F^9(UG9O,4@J#JVRcJNK;]8W<@J,IMW^;^.Ua]=bcG/+1
+Y9QNa+HDX\e8#=0).QCRNbU-/ZIW]&6EXFHI7f_b(gCG@R=cA[9EV#W20/C]@0P
@fTTbQ/KS8^bTYDF[[bXIf2.Ga.;bC6UWU<U&.^6(^NT/R=O8RDW+>8=H<:4]P^d
f;W79G+WcXJQ--Ef8V,)T6,e<?>4T\8>0G[b3=g:5P:H>.dY7MG2Lc;?JN(L(T]J
ED,L0bV8/.84d]f5MN+Z<PJQG(?QA&JC+B?bd4EK=Y[ecDK]2A1/cd80DJ:@^</-
F<D:Eg[b1&<?A2N9IXQW2)BBHA#B5VA>^7fUO0ZDd?.e^XB_A2VM@K;V)6U7<^Fe
R9Cce^:]dY-E=Y,ZHd+SK)J+Jb<RReVGG>f#N=.W.[KES]^H<eR3O<>Wd6@E+E9f
fe^+;\9=E-,ESG?eZb^,LTSBT-&]Wf_L2]1Q<?(9Pb[@:G#:=3<6<fc?Z;&Q4B:V
6HJe/KLBX#H]B527]WTU_.L]#M^b,IB<+)\+Q#6_bW]Y&+,,/O)NNKB:O60ON&TE
Ua2\<VQgV1,Q;A?EO,]d+9B],OeV93b3N9_TX?QY@UC,b:T_(5UJ>fe;E,MO-QE4
##AEV&C:(I5T#beN-0H#eTR?Pec>28#C+OM\]UIMF\X,X9^A[&P;MT=OEIe;d,1]
ZNOA)EZWd+F;4S^=g^?dIc6Kg?I>a[EJQf(HP/JMEMB.184C=12SL0<[fMIO[V3?
/-T<4-KPQ@HW9UaR]b5=63cM8dF>W7]_X6DdUOKU8a]3cbWR_g-.^R+(.f_;JG9;
abN<IUacQ2J/Ud#d1ND-AGU)KP2[OPbgEZ\WLHd?^]LR-Y-4EQ_\,f2CX6GKX-WL
9KO9f)9R5WeOGcZJPBDH7Y#4,Vd\_/CX7+;.?6;f1LSa9ER8_OKV0>/<eP6;.UM=
,ZDIW;YI9U9,\3.72\^^bRM&[5T\a9+:7=-QdZ_U&27bD/^d=d63@0>RU;/ed;XC
5(/B=GbZ3f/[7<.3]VI[;0L_+S>1f\ad_([[b?.Lg3/0)C\e2_.\3b3\2[Qb>HU.
V)K1\NHC]#6gJITINg7?g^)[R\UIK;bC,L)QCWOZEa3&g]>f8OU-6I\f4.bg@_[V
B.&YdPCA7Sg2fGALSM07,<R-8_/1.-7=?T+g4V2.gCQ@cB2JUSTB:O77:M4]gXfD
SbMKGI&&IY0<L\&V=UBcRV-35D-Z#R/a8?aX+A1;YJ0_<QTL3#2H(#40f-<4HLFH
cZ^B:WDd0PIEFKOdL\5gE[91b]>KOGVZ=T0(S@FI)VRW5aM@)ebH0GcK7H-6\,f1
N1ZBRWSbDdJK,:#:P+4-^1SK[b).1&>QZFR:4bA@g>6bKOW@NYc:FP2A.YR=06Mb
,J][O#->GX74232-<=IU?Ge8&KUD(XXZ>FCWdS;\_Ydf-[\?\;#48Z/RO\\NeGfK
@LFbIfCM5/WF7]c?Z\H28,QKQfY5HJeVKRW0VdP\Ke86<E;..Qa>3&\1_8cee_M]
]0:^O<LRL<QF_(_8D&LEb9>ebHe]^LH5cg,C,8+Lf8-c]b0:UGV<TI&bGZW18DNJ
a&\KST[+32J6Cbb4FfVC0B+VY,#_BB0).9E+7&?3T-+@EQLTb1M2BV.A)d<5EZ=;
((Sa2O5VgSaD^//HSGD)(CTUSaDT=:<(+VY6_;5QJQa[g^7:6HS\3PeR-#=#<]9)
-Q?2>b9=2,ZRf+9OYINZ,[gRZ:&-(dM3c2=F9_5^J.AF,PRLTQC>^[RS(_=3=6NW
^3gaaXeT>2f/7@GQ+EF&Sf;>LWd1&?aK0WA)bWg-1gS\P5&?Ud,/VXOBZS-,D<?e
PO71f1M5I\QB9BBLVDYG&b,IBF=:C;./([:;ad.3_O1DZAO2eHeSB)N0c6=d_c.5
?0UQ/Db53d/67)M5J>@BJME+5]]g1I568g(b7V?./dD#NYa(KcQ(PZ5Hc2]#08_(
6LHVX7Wgc]0^8a/]^5+WNg67Eda_,AFJ&/FBaG?Z/[BU.-/#YZ2CY<^fb0FMZ?9^
EOSPbX5-3SR7O8HIJ=>S&Y@-[WfGD.(@[DASM^fQ@C@(D9(RgdFB<EF6##<WTUPE
^(;3FJ=^UVKA+N.dDM^c#9U&<:a=A:[.)M(g+(#^WcK;N4L+U[+&=a[]L>40>KXA
FV@FJ:TKF&,>MO8)^>S=3WA.3]X6+IXEABK+^a3G4bFV^@/FDD8G87\/\V[_[=-[
#T4#b53fPEWWR^^K?:eK(daM/bG[/Ug7ORQU+RcOLdB50BCg[V]4OH70YDS(&4/^
G8^VPP]Q/#4e:]dX<?)]=/==6e)SK-c0_T#_GR_A6e7bO=e;1bBSAWGJQ.16/dFP
=AdS_Z/K,RCAICO\^Q3-0(#J:]Hb99)5)+JfVFg^(B_/)49,.G#Y;N0Fa1gdO_eA
(/e>-L<1aAV&<_(IC=7b[e1^HEI]TJE3/a0O?cU7WGKXYa?50/gKR4H6D+a+8J^X
]U-ZG[[-f98;.-@]#/MRZ:2897c8=K=2U:202?=B<(CM[_D]Z.gAR7>d/Y?EKBNJ
:,Q.N&,Q)VJV?TeR4FTOJTDCH0/.NAC:eLG/R>[7;,2=HXG9bM49-_AV[^B:CG/b
H4e,^Z(PSF1AEdF0g)Ne8]AOH@<]&a#)M&JSbL)(Y1Zb-OA/dA+QB]+ET40ZDfO)
>RYBJa-JMKW]eN/<+1F#[<<\QH20=8ZKV-DYR=cGSY)^<\RC-@(.GH.XfTb,J;&.
6_7SP32dQgfZ>&2=Q<M@JTQ]/-BYKWDV<,[N+DZcgXfDW\dRE/DTd02HUeU6IG>e
84SNH3(.7QCY\?fLgeDcJB\gUMNS5(\5Sb0G1/I[(5C^SOI9b=TeY7c5ZbHT7;]D
\O@^#)I)YP(N5FAMRD.BT@&_#J:Y4&fAG6T<\>-70=J](\=2MN6VW[>0::4I>43E
fSF^4c4:6>CBeZgFBZL3cgZ>GV]=57(a_K.e=K76\&bTC7BT+VGF<&-RAQ7(8CM1
N]VQ3&R,(.]/4:R@QaV:eJ]L/OWF8O?F,L5?.L\CTd9cBM3M_@aF#R3:S<?P.a(B
-=<,KGGgHJ6L70T;5e(>6G:#g]7O<E\=SI&21CdTBC&[#_,)T)D:?6R>8FVKNL[f
=PY>S8EL>SW7MBYc<GD3B2bd=caW<3J#>g>CQICB1[6524U(^Ge)^+);e9QMR&;W
>712c63S5,VBA^,81gJEY+LP;9ZD?JL7F@6^FDBg:Z)a.;e.UZ+Od6?Bf-H9&dcL
I\T\?V>):bK5<5RI<XOg,2CZ/eW1H]e)cX@&I-BV..gaLI.G6e,b-=S5C;Y?QA2E
H+7,--R^_N627TP_D/@0LaK\,c6M&0=?I?Ja7560_<4Y]-W0^-:d(F1M5N+K];PN
.7](&2aOb+J:AW,KcV0NK(DZ_\(eAb,3.+FC/3D&.\U:NJfI(0f@7;dK;IbTX[<,
Q+JU.+@H?SO7JLS^+]EOWM/cC;-&K9;H?gP(+A:0Qd1O</R>,FeeG7cDfG^c]P3:
fa7+eaccX8RMbHF>MRGccD5ZgX[3K=d7e^E]fd)I56L5<Pa^g^R>X>@=<5^PbL]5
9.##L]V:bB>];#XJ>eXUM17?3]-DGJ;DB:)]>_gc\+aS[\VS>Q#C4BW&;2FQN^FJ
#B#=&5-9Qa,SO5R[61V.)<_UQRaO_SWSZI8ddYLPJLd5Ta\KN[G@&[f51HEM.<Cd
Uc6\QZWb?>RFQ2KPN<UN=/O:=VR(FAQ#>98aBf(DUS3J0.[UL&b\-MB<X3SZ0G[N
<BZK.3)8Z\U0N>XE?#Vg9bLc7337+9?HN5\HYVOK2DSIAc_9TQ_BNFNI>)ZLZZ<,
9EV^ETc;Fe?9&9;aXEHNSb]]4+\K=gBYg0/9&Z&\B8\agVL908YeFMD;>G4XMcMa
R3,=3<O^E7WX;[J>J4?bZc>cQPEK).e21Q[ReZ1^AD[L.I@Ug&:+.PS_<V1:29L;
AVe9C5>fO(4@Q2FJM.+B0PX9IPAM.9T90eaf6,?0,[2W(E6P6RR2>?&M/.aIa]L/
4&IGBN]FP/+aTVCGb1QV^,d.J02&cWHK^W/SdK03Qg8J14RM.aSaM9G.P2GfW)<6
IA#CKT9F7?GH^L1W0YE=:-4T.R[faa(SLQcG8Ne/U3E&TDCMMA5ZKZ:eO/KcI7<c
-1WXdGY)YC_bAg<+MD)YJL:J06/A3#?&^NR<EE+[\,J5D-g-2_1[8R.LD@P1C@Hf
Wb]7J_(RL^&690H#Z#+FJJTZ3QMIa3ISa#\>.bMb,_/2Bd56FX_0=8EW8=HIM=:W
&Z4YVf:MVOUIf#Q+?6^;WJOce2He#6J:\M\SB5]5]6OSTE/GI(2eRYFeb1^/<7@3
L=GXR7gBb/=Ib3G^?2@ZGDf/,-):L:XHF?OKOBUE23cX-U\S.gLP37\2^6]M9V]f
IL4F7EC-(),FO3I03E_;<J;9:,H+g#gb?8>c/OdUUS50SD7A[W(OTNG)O?:WM+ST
e,4G(U<TU0_=2VWfFWN:E1g<+WFY38P4,Y-Mgb#Z<J30CZ,JgE]SaZUBV2MI0=<K
(>[;&-4VL6316<,>NcbR0H7CY;XK_?P.TV/g0=+NL(6T62&SYegeNR0N@RFRF&>O
EY5KFA/L3O>X2,MR\O/:.(bKJO?\K_aTgFZWZJ0bS&526#:DQX5K)&-OaN)bKcNY
[UJ:<]L5F<22))bT)eUcf2JJeV:bQ3NQ6AA+J.FXSZNb\BH?YI#Z(X2HW.KW+dJ<
8I@H?-.M5D,?\cZDf\-G2Y0>7+HRO1f,:/f,CIZMZLAW?9#P06Z?^;^,0<Y>bXHK
gcX^32W&VXT=Q@8,ZDN8?e27:]GF6,R>#&K\+cQe5J6ID2ZfPL.c34?V((&fVd95
^3?/N4:<BK+E^Y\VJ32/SK)UOMKA4\\6#WM,KR[Q/-<>3-R]f8Jc7\(b<KPURZQU
]_8^7>2^2U;a#cc:(F3220:;e:1=4N8IGFE;MDOJB7@:dOb3X=_Ib_G3L#NM0XFd
)&gYK&]dGFSP1#9]]VH=b5Z52UbW2E=C4GF\f+feYg]SSFQF/GB:Y8bEVHA(cb3E
;(Ce_c:>?(dMW>?gD(B6X,?TW\(cEXf.P9>^_L4TI/e\GaQJVFK&/8K_.>Oc#-,5
1SW(#E].5&7JJfX4Eb,&@bA\6(&X0(]0<?c6OEBag?#0,87CAY(IbK>-I-Z8e<71
2QO6-VB]+LPQE07?HO.LE]-c^>F258:=28?KW5ZD=YPD58_X4?M998&.L^-KP>)b
E0>2]O+@2ASSNGOeL;)PH.5b#:M@?\712+4?5OQN.eIAOZaF<4FH#J4>2/P<1:()
X+7g]^3^C?10e#G@]R<DIa#KKOa+B\I8I9&aV2H4XYX>fD8G#O6+:/Z(RA[L,Zb8
:A]._/KN02,1g<BZH1J5)KdD)Fb8Dcd_b7(EU3BAM2JbH[^Ga\5C(;+KLCZYA=C\
G\0dW9?]VGTXIaKQ7)KAU]GW9-X@T-J-\K81Ha1,\/T.)0JF1MEd^]0FLJCPb\d-
0/+dW??N#bQD[)8VTd#_VKaKOe,NQG#\ZW9U;0N6cZ:>P)2)#STM69BJ,cYEWSb,
Q-^Gf.QcD/XFT/e(WW@V+]5>:ESCQ0V9HGLS<gcg9TFUR43OO\Yf3L?\LC&T8@6<
/P2\,5NJXURQ(^FUT?4SC61S>-AXVCfJ&WC7eJIUcOU&16.OT7]N@HIR@^O3ab_X
0VLRWS[g^LZ5)^ANUZRL/J;7fHN7b?)/Uec8QMY/;C1VKd//@JN=]=)4J:g0@cC.
b@-BC=6MM?&=8fU3ULF@BDA\/-2:;T022WgN1/PA7L7NZ9YZNB48Ge^bXBH9X3B#
D8gE2PR_IH\\T++4EXY6#g0\^>Bd?6+2]NZ4AOVT)\^>B7+6GKT,ZQ&cDL8=9B^T
fVLZ5fe2bG+cT5Bab_@+^8XL5(H.38a.64BVTgF;gcKdJU]>LM:Z^>U1<c./(^OZ
0F;-cFe[^DP39_OGe6?8&GA0gJf3HFJd(D0.88&g]cc6+_>ZMdd-J>9FBFJD#ff1
MVJC=2cNAFLSA>Xf4_-3L5\d9U<AN+1=M..JLVTM7X)^[=fPK]:4EX662P_3N1@J
^7a/F.M5U4a_TL0f[.FYN<=V7PODa=9>af;/+Q+Ng0N,(.=A__1;7FC^ATJ<3F7I
+e:.e/6XcT@GG[>.<O(;T)P[9V43PL#]&,1EA];ZfT?_1=[Y7N?NF-;#8S+;91g(
K5X<U6FHBOdCR4N3ZY#0>[&.Te.8-=3f[c+BL5B&)1I]OQ7U&/c=,]3\Ea3CX3&0
Y/\1Be9f?+D8D_Y_P+I[K63I@LG4GLGO758?H,R;CRRdJIEMA3RG3\MWS_@CR&2-
I+QcJbEC]]I@X(c4D:C[NQ@K4WY.J_7,;_2gK5)5J?ASR;_,)TTUW[X_)N>f.b1A
4]?K;G.XK]I8A(AS>Z,FHHA,6BVTc-2?D9HgSX13@@(H)ed6LQ4HW@J360TW(VCc
[MX4<5J@OIR-X(04+YO_9K-0eaP^dON@,T5eK;3#^/dYZ.\LD6^6JTADeUO#.L40
0+:M3Q[bK&J,.UM+QEBQ63Ib9#+#0IH\3PC_9VSOS8B50QfT(>4SJBC1WX>3_fS>
2SVF-<XcA\)[e^A;902W1YB20=)Qd\^E6ML[Vb@_e_4_?RLY3YD4HIL9g/=V([Z6
.BV+KG25FXLC)(&/<gJA4/DJfL3+>JLc^0Be>d.\VC?K\]#9A3g8MPFSN_W^T5O&
O/DHd?_E,M88AAVA]:9\EcD4Cg.C_J24IVZ:Pa^.6ETC,TYG=42,H\#N_D3+Z;3H
Z6S_,\I-TR7(?a\_S#>8DcN]d-QXb&-C+A[G[bT#NF&J-]7N6Kf>5-RC3B2NZc:F
_N8E_T-B<+^@DKbFRZC:MGJ_+/I2]V[&2E57f]RXg\eVT?#4/JF@^<8P-VGI>DB]
PDYP3N=4ZS#NXO_BeXL#7[IUZ3?d.C9c\E/AKBb6;OL]:g[8A-FcF#&A9a2TM+UN
.>M.eM<VWaC-00Udb>948/]_dI_3AS:.P4=gG7?O_0a-^QUIZddK+ZNMdDE/?V87
FSaOL,9)4B9(ge5ca\1_KS?3;Zf2MA1g:BBQZZPXD)9E5]c]VOaN_5F<H?Wd9JIX
K40/9>V-9edN0SPGE=cK1R1YMP+<\W.MY//f62bWU7UR.6(X(D.2_8FE#bPY#I_d
TKRd21HQ_#>)dRQe_5QO7=P@eS0&B?C;)ZDG-GCUA3:XWBc8\O=-5,eQ^#,0C=)Q
K^SU;BZ8f6bFb&R_BU_g9^M3;.21MBM^PZf8EFAT_1(AV-Z)J/.\9gN6=c.;T1JS
M)J5D/N1KV:=e118\K^+@G4Yd&HKM_(TZ>Y51:L_f]X)\UPM9f-c8^N=-^ZgT;-+
\><c>\,;Fe4>BFeOC2OeL6KXD(I=+\HE6@Hd_U734J8@b:++c8(f8E(9P??PE1c=
@30b__6JHBV_4QV2(.e]D,gT^:),IH,D#X>#WF.#1geD&A(_=f-LIZ58d//50Y;Q
?<.@<R3/JK2;ZYX/4e;YBN3bLS(NFc.EZP/1MCLg00+b^cdBYX,Z9I9_0#N?/,MZ
1F15693aOKR8DP-EA(>,2UWFEDA2F>WZfAU<U2XH^R3f(R<(fc8H&]e_KYMN]?JJ
8P(.[;Hg=RW/Q-IaMD>BX3&6c(B4HT4.Y1\JMK?>YWaKI0@J1Q&8W;0^D24_#<P7
/&88^;>3UIPCR>6VU,[_d-bTX(J>+HMcW&^4,&OXB+T[]?S.<NH?DQdMPW>MJKZ]
DJTH&7]649KIMJ4\(Q&>-c8Q-:I_N:1W]S-^Cc,eMAb/>407UA]fQ)L91MBM;I\)
W=_C.?e2YYI7+\f:cc8/C(LY(:YI1Tc/.L_6.,8B):2G>5/.-H>H0P;-QBHL(76)
_#96)6/<H\/:K:@AH;DK0=91Ng[)ZS_(EQc4,\P9(dO9_/T4(_(O=7(R]C.<MND/
OT9A/[J)ZKMg<#-eU0UOg:BOIMb:\R+\H,LKPCKYHdVSEG(dNUf+0P[=37[YCI3A
+HV1HK2&<RbTV[2_1MP[JU7C5O<5LK&LY:D>4_JK7DM-&J_/#5C0I.Z7.4(g3V(P
EN\e]E(&/4O;YPXLR,Nc<WH9BeCTgPSH[7.W5R#0\+/MADe26A/b]41#CT4L>@gB
@):cd>WDH?XIBNIOE<90WUFR#VLCfUDC5B]A7^,>NS,T6D2bS/;4PJM7a:3:Z>C0
10J=PVP/Yb]XgC^bO60+(G3b^4X3K-[V)e7Ig@:T&LT1d=-.]c0S:B);@^,]5_(<
B^EU3^BdSI=Pd;HTe:,(10U,(8S3ACbQbPCJ4.Z[a:0SPWeG_LC(AdJ:&2V:E5FT
_-GaT,fFe[61#E/Pe.S@T^^b()LfU_#^U1>::_\R)O_TH4dg(K^:WG8F;d0]bcK0
8\R1dd)N?]+O;d^G?\:5A1AMYAcc<YZVSf7ALVD52/:Oe=5PR0NP@)5P-DHU<B6Q
CNY,^&bA(U-)gR?F-9A4Ea^:CCHDCOcfa6He.TUC7-U=-bNJ;9aAWV5IYAU5LO2W
W;.(JKHf\<\9&e7N1XUW-4e_#:G&K?,Z+B3GVVg1>ZAAe@eJV/Eb0C[:[K?XN-=P
ILN0)1>33Ued(U#a#5I-=ZfdY].6BW@K]\UC&4]WF?NgRf-GBgcbFfWN4IB1,V8[
@f.d/BfXbZ-a_]2].JJNWPE-/M7A=LRIE3eBeZM+[PG,4+e?\)INS(]9HQPafA9]
OFWe6J;fS_^&R_e.fM4-H/(2)IHa/bRL4I@[.0#E^[-&@77F-c;f982bS]FQ1fZ=
P&BBD0-375?3\\AL&1;VZ#CW=BG(;FRRXJTOc6YYZSS8P#[3NLV]d^cF0W<51I&-
+52_])O^BRK15,eS+J#4XC.T&D0c:COWgY0(M1[cGW-6-Ha&(G.cUSLC(0YR)POC
,^04[SJP&@?S0WFK9aW&EXCJJ=:^UJKSQM2Y&E-1N+_ADM;M[;ZdBeW>/:5B2DV5
PG+T0QFJV@CIK/:FO^FE8STUa.>M2;cK78gP,QN4HAQ_#73D[IBW>TB-H.46X#Q3
=><D?[RfPB1G,g)-5&=IO-9WC7<#(5:YL7fcUJfLa;:H?g(4B##Le4W@\fGP@ZV[
+JfA)U8U]&EXKcSBB<K3VJ5]:d)IN]fWdTLBLW6;g4X1c9<J6>H<,)g+:^U1YL#f
\,JDPf:T=cX1EZ28<\-;GLT2\6>a1ZNQa(bfC7]WM\?=+ePDaH4dS<g6/Y+Lb6c3
5N7HbEe0FJ),T2C@]V?VK^fTb9+03J3>4U&&@_9A6/17a^^/H?+2==-Z+Y&KO9+5
/caA2Ma0_(gVEa=>+F\91Qd:C6,TU4e;#42g,.O^S+eOJSeF[&X=Fc09Z-&7EF=M
;d^0XO,.<cOXML]DU^?-K&S\ba7M]bRC7dK/2R=]7_^0g>NGYOg]+8[V0d[a;K8[
R]Cg).JR,<Y;b0_KV5]RK3<E]W,IEISU<@;._PD]_8(.V9AZHE(3[B)[99bdNLIQ
S6JP[Zd5,H)I(5(=NCg+FE,;3=+?TS/\JbTYa;OJRfD@4f=K/BCJ=0R;c?PUR>D(
7cc0ZV^FQZ[d1@T;Z<7@7RA=V/E9<;,-\eC8G,[V>@C?@-R]EK;.gA):@O_T4[7F
?HJ11B:T6b6RNN7<FNTZLJKa>+B[/Ne-,5LA,QeYT(XdZ7g7C]6Q;[1bG9K(7PXX
N&fN#X5^8L-[PJ.^BQ9a3Ha/9&G,KU&CI5]5_OOf,XB#cMZ<DI^\X,gFYVW;\3;P
?eabPBM/BSeKC_S_J+C>_N]D[Z\IXeY1E(NPa^>OZgT&-&@DRVAHM7=AKee,(ad]
[/7VG@QF&8LM4FQ\M7I@fZNB+.c9U9WQJ1R1#Y7<H<.J?DUQ.(/#?V819_[W_S;#
V/[5FQ86STM(d)+U@T]&f[7.\W:CK[RX(\N<RBLK<bL=3cQ2&4U?KY;NSb0?)P48
7-,3(EC5;5WgE\;19&:112bSE41TG4S=c#HC&HC/&fc7NVe4)?<@Tf>9b]4&aLcI
Y#V_[);]dVL#FO(3<EeC=]0.YbCDPA2EfCFN>&?dKR/bL][R=]2BUO5?I)V]58M5
<7<I(++ZLfG:TEBTX=O<B+M+c.+(BZ&8Za]&NL?KK\bO:1K\JH((1.L3O:JUE1Yd
bRX_>_c6NP-?4P^cZ?/UZWEGIe#g5E.GfJJ?>D#<f^7dC66OGG_\R7Z3#IW+>NOc
<<\M64)5<534?CFY3d@;[#&WI&?4&0\8Va/@L#]87a;P:_FPbV<&9M.56I>g/43b
-&2E9C0Cb@-0c+/FI+Xg3D:L;ZT<bSdc,.Z_^Y-N@6:A0ZR(Nb7E6.VD<\?G6ce:
9#M?84J-be6^gd6#V2eO3(V4#Sf]Gf+f3;R25^&,Zf,J5cZA__V?EBXH>KH;OdA+
@f7&^?d)@Me1>d#T7.U)CR6(S0=?VdZV0?SNePDG-f\GB015G^XUZ,E_A,C45V-?
Q2G?cS4]H82JLVe62J>[;77^H@?4Wd-a:A0@AaG6)d>aRb]6;K4ad@SY4IXSY6bV
cV1NT10&<J,-LTGNQ=fIV2\?6IMEOe7)Lg5.W\#^2P11F9KNKJX8<\??<6^DA_=:
:6TFSH1.&c?Q_BSP82HWUa))N6R\4[O/MXTJTd@;VbN[DX8.G_[?\\X;(4JX+XRK
^d09L87DLN1ZN7^Z.d40<<;G2dDVPA]Id->6^?g40941=R=Xb\L.PC_D-IBVNPF;
UU.PE8TQ:,/O.=S+F3Oe35KKN</:@aZH_NG4T@Z;A)WSbMeSe,TXYWWUK#Kd(416
B[[^Y+fG^,BCf>\4IVNOD62#6)[3a;Lcf9DO]JMLA3[4II:/3;CXNeS+U&J5[XLU
O.[6GQ9V9@#>_,VcDB)a#d74a8MU;dXWTG9X[LRT7aJLYWN1f<?=b;a+8Z;WU.CF
LQLT#+fVa/PL>QRB?+VQ24\OT6^H-::7Zd.d&@J?(f]WdR)TJNL_KCeaR+[M4.1U
\&eK8S^IOKaK<I6B3bRN]\AW6<3cb;65;<>P_UESRU)Y\BdP2:95C#(-4@G&V.-Q
4/HAA\aF)EfL;+Vc(UYCGIZFaHHQCBf;6\KTD88[)b^Y&#BM;E/1Q1G79D0>3NbX
R]<VPH)G,TSG?\^09;Z(g:L<UY]g@JLXZIF1K0M7ZFc_f;_5C7ef-+?0O=T^QDW/
S,BAL_K&e(XgOM#6:+5PQ-C9b,g7<QM85_aM_1TgG)_WPc.08XC-AeB/(Y<dRfZ4
5Xg7VGF9Y(/T,V>H@R93B./[KIZ/\C]OEDfbX[5F(DgY^CQ3\:J7NO\J?-6G)d=?
ZT>bOcf[[E;PBX4H\-LZ/FG1a>XPF^2\)Z]:]><ZW3CC8?AF,/eTC\IcICX-PQQa
&GM[END/);RY#=^TG\Ic5FA6_7gHaO^a@N1_2HZTMCbB:VP#_^,V/E=EP[C]G-O,
&59_;,&?FF:)c0O+E/_Eacd/0I>TX?B8gMNCdN>+&3Ue/0(VF&&SeFT(CeZ\;)&d
H3R5=3Z[X;gFJ8BPB5BJEaWCHXWS@0_;=aES[7eJ](]\FU8)H+^E&F#_g:7L<RIU
4^.XI#CfS8:;^43E)B:)-Lc8b8AgP-[>;QHV[(MHLMZXadXAX>)__NK_X+,bQ=LY
I-B[B>LMPcSCeHS58dI)AA#.+4C-bVYcVNC47M2,O1?F#2#46LALaDBLFQSB4@)#
D_+K<V]YE81)(\CMb?PdX>XZ-VcJ):cPFIQ/bYT2&dI7NIW@)NYM0OT,6?,@,X6,
a)<F@UA>e<UgULH:A?SW0WO96>a<A11QE:7:f:)b)4BaC>H-f6L,.S-eX?COUAa8
SK[SL?020@/)Q)QUBESaP\Y25@F.C>Q=3U/1/gc+8^Q5\[O]8fEAD_YB&6FK/PFe
b&]V;NSOV3@gfg/<bLO;9F<57:#KS9[1<c;cgNH)&<-I&g2GXd5V.7402@P=JeED
YND17ICDITIVU1@MV0g^H+>(8OK=PK=L/)4H170S>>T/K.9L9,C4-PK8R@D&7T@5
4US3,:-)7;H;B_M8J#/D<W]Ma=A5,72JT8:=2DAS#W+aLf[^LR(H6(?ReVMOK5Xd
YXVg+-;M\DY\+H#e]63YKY[W+7=#ZBNQSYeML+&A;X6gEcQ#&_&dB/C(/4A)V#G?
60YH5,3AGI-@Dc&fa,cV/2/6B+>9(HEA@>#EVNZ0MUAF-?:-dQW0ORZf&;OGg=0\
eR.f\QS-aS8GLH)WTDQGI=.I-eQ&H_@^3P&+I9?INP.]A8.#-7gKJba)=I5<<AL;
GMQ<((GX/FZ/U&JaKSb/QJ5&BO&<Ec,TLAR>e8_@V;DMVB8Q/eP^ReJ/;G]VPF)B
@CW]U4LHX)+eLK@B?6S/>CG&a/H9((S.@YEUXQ,UeC:65A0gTBbR=ARLd](A4Z&g
0I,P#=]6266,&<_cUBg/eQBVeG[VLZ@aWX19YBFYgL,c4)-&\\U_LB4bSKcT1^/X
/<^R5If6(VWDdVA3JS5X_KLB0X>2B?MFS_RC#E6JV&JV&DPJT4bZUXV/#@MXOfZ&
X&D@RU+Z;D[498G8Gg;4(:==RZ.a..(]Q3)UE_(\dZcL?e[+dMMHePHbV=#XQ\=9
#BG)Z(?g&FF<aH32c-/D4b9V3LDCTM(?#b0T.8HZU>4#BPLeVG,U8L=P-g9E6+ZF
K+@U;\I?8&?WfAL2WR4,\Gd4\=@A)S8P:VSTYJ[NNEQ=,-UOG+_eD.;XR>f)6\@\
bG_NbZ3_IFFN_/N+U^;>SYH)ZKe2KR+YSXE(;3<#D4/@;.XVIV+WMA>R&V[bXO@[
OHcAW-bN(GC)T.N]GfHeD3BR3>)W&03De.<(e=IEe]HTb=+YWg;Z05&b2GV\3X2\
?:8CD.S7F&@ED[XJV[cbOFO8RfSe8,-JD0J;JGHQ_6D9]b?)JYFX96/6Z(FLE+aI
Ra4.BDL,WA,7[V#DR+&=\IGReg7CE0e\Z#Sd4P?&T=GBU(0SbZ)@-G1Bb>&7ZVL2
[77^c&7>V-AG_4b<,c]_;\4e9VMY1[eJ]d.:FBX>.-BZ:8Zc:E^.e5b,=dca6YTU
<V5KHc&:)d)dYg@#?WCdT9LbFCTc]LJ;?b,e?=1^_e^/SAOL@WZ3g)(4;^H0Q+Q^
C@Ec\cD8&7CYQ]]e8ELXA0S1#bTO&a23B(K5#X9<1E\<HY1@\#Z,K+2FEY0D]L2Z
@7B>K2Y:.BJ.C5)CV[PYebc#L_FC^4d.SSP^0TIMD44GXM2\:Mb=aRCZTY]DAP/)
1B7gAaG2CNLXG4>N&1D6,C#DD/<06g(+_LFO>5-/7F[XI)OG?.E?UVOgQ9>(2_L#
=FUEH)>\&J5WUL=McG4<RX_TKD_^[gJ>bOK=?K_Y#d.3bN36I=@<X?]dD>QGJX85
98:#HaQ/Led9ELe<@UM.3,)Xb\D5dHb>CFPf<ZGMK[@@<2#gg=B8+Ogf;1Y3=A;?
d(W1g.b>aCSe3@XH7gW?MVG0?9J//;2WOQC)L+[K.7-@#aI5G2UALS)U833:e99f
>KS)XFD0c1N0e705=/^UO#AYJ^6J6RTXeQeUCLB-/X<OXPIL;&#GdKJ0SfH#W1&Y
JBOHW,1=&XHGG2=f(<c96818TY)O(g^.K&AC0L4FdBVB:GQK0,H_d@^<gIb#4fMN
T^6X66A<8>=<<..c0?]1R2B.ZX[?24&D:K>UE<N_N@?5ebb]3\X9XVTF(,UbM#VC
b&AI,OC[JG&VOU=^+T_\a<b372S]>T=UbBgJRT=X]61>[QDJ)J&^5EU=D,UcTVUQ
Z5aeI1J:78Za:\._V:RHPC(ZB7IF#M/A76W8:;:&BB]]FP:YTFHM_6ZVaXM9&XWN
I:gf?4gbXc0LPOA@gF7.\IT17@?P>S_a@LaFM_f;85(Ne;d9A+KOa=0#Wd&^OU_Q
UQ630=PW3OE9V1:6?;>GKBX;\4(Z?:>(D,=5Y+DP[d+,A[LcIHTZ,WLAg\F.B,Y^
2R94dOE12g5.L8Xcd&9>NH8GaWWY>V>KU:;Gd#AVWMT(<eIB_e03BGQJ5_(6F2G)
N04@(VV0_QP.0ea>eBbE^]QdEFU+)7&=3dR9a4acfB1#_VSN5=8&.FZ\]?Ee63XD
/T0]Zfd.1T=/]5T]X=a8:[F9@BaGXKb=:f2]@VeYfcgS-;.,/;cL)ENWF8R1\+12
U9U.</V2B>7)+4cT1UUNMbH/+<T,DIdE)VD.+OF+Y)3-N#G2YY.AZXMKIT^A]+W;
PXX]QH3#FO[OfY+@,M^b^8YB0;___^NQ_TfH6YWe=-)KH1F3\a1D\Y,06+@AAg]_
MK)^4IL^ZYT-TX.Q1fZ4L=eVcaU&[ENHPSX<JeHFGa=OQYYM\U^/1YN?VFY1CUPc
63>eg]eP;/eeA9f(AUfI(NV@\Z>U<O=.242;M)0U6g&F?_M(>H^E&0d1=U6U6c.7
fVfKD^&AY@G2E?ZU&Q#&7KS#BO^Q0Q=.5RMTB,c=YbSD5MPg)670\TWJbQZL-@FS
?-c^HKP[+AJ<6P9Le_ITNGb/^4TV_(OAO[UU^&ObHLe\d[We#AHB6b;\C7)f_D1J
POSGHdSab=I/KKAT/E^AR7,SFaPbXL<T:EUM0PF#M3d1<4(g&eJ3PAW;XR>f7-eM
YfM9#g?T9C8E)Qaa=f)_[OOgUO&c[?49>HZPe7?b.8Z\V23CaE>5DcX78<d7O-M\
^4_G&2\@V71_P^cC^6VM+2eBEWXL^PCF39g,+I?dSJM]cVHWc#,XRCAQ+cZFZS+]
dGcHJ2L+11.<TH0]gaX7BP.9MgS?U_7Ae9(<E^H^T77Q<2WY7RBWE/7U)D2.b[\G
aX7<4eT7D:S)-GW;^A<K#LE;)e3:B,ZH)\?2c\K+QU65XS7?KD3-Y)c+?=I0\AI9
ECP<],aO,<:[dQVUaZ>JE+/DOdNB0O-)DFgOcIO0P(4VQ4gDR@#MfJIZ?E)2026:
9RUHbaYH@,V)[)<gO9SdP4S;33L#AW,Z2ZSF3Tf7;\3aS1@;H]F3&AIKI_E?B9f=
ASW>05gV:>;]aA5N1\dF:LCCLH@49Hc#]dG,6V\d3eULD.A7KQRVQVYf3d7cYBR5
L1];[0M95fG-JDO9PS:U4^U7bW:f[@7gS7Rc5EAMPTX1cBd1>OF_3g1\743J[1>7
O>:c3F9,BJe/9W9=5@LfbOY1EaC5S&JV64,cM5N6IP7^[C3X)V54QfBB<7U/=8Y_
\2\4>6B;N\Q5P9D9A,ALBJN+c1f.?V9HGVP&K8aC\bKbgBE&F48Z4)PT8KW+<I6Z
b#NfSL/J-#/0A[:9PcHCM.NW?[R:P_E1\[I?:^)LP>?YHYN@U5^Rc3LaL2e7b(?T
[?X3:.3.;b<ZO?VCUQ,#a2KF#[;/__DI5f<)G8YfX,PY/1TS?YR]34FW^ddT@8V9
J,];SSd(Gb@aT\TaQ^R?/,XAY-:7W;6R(W&AM03#RE&\WKY+2>37S+G2A4D#d93.
5K+O-[ZU\#b-,.27)<JafGEN[5eDTVUXCJ22=U99,O59F8c6OB3+G3YGM=YXRa?G
)D4c+3^f:Cb[/NDTFMNU3c5#>0gI?UB6MID2,Z@+8O[TU@1Od,CI)FV\HD&;4HON
IGG36>.)1eBN_?H^eWU<MU(I+Bf?:ESH/+#)QGb7[ZQ.gBV37;MLQ4[+b1cS.+V;
94gcF(0.#W;BF@7G\9/9b(O6J_#R-F3],+_XB/b2H30L7S0YH&dJd[U/0F9G@Uf(
:_-5GaI6b/ecg;BY=()\67TdbSM/NC2L5NB8>6;6A_3>J)T=HW,02+#][UWB61J&
HS(<:D]@fN?O+FNI_7RI\1G[XN2A(.]Y_KOYKJR6=78,^BET-WT6Ya#8>7Qeg,(^
Ja\/UY3IRD;NMS8L[bc)Q\edZaRU/S?5]\^CSQTVbJ01IXUDN4IS0;]E2>+HC,6#
/K[B[7<3HOS0T(;c:eHS8G9;0+QS,=LHgWLf_[#SM)YYC51GSeb6Lfa,&_#ND/LR
@P78:FM:D-ZIa>:H0FXU03XC=gFU38>LS\g0+:F5/352PE+48UWIHBA;QQL<=BRN
PO@+]1dga:e6=aYU?Y#-]RF6e?.I_eGNgP7OHdUH_d8Y_,LQ2;B-<3A;d@J(U2\Z
/c=2K\86a6X&_1D]S0=HLeEC1=+2aI5/PH(=&P=S(8,BSX5Gf#gBM)JCQ-)U0bFb
B^(G)=?UZ&:eL>S)WcF+0/a+T6WJI=6eY9_b1-.S=(Q6Z+-GXaQCL,Uc[(aP^CJD
Db.@L-.dSb<QKIN6X94TJH_E^X0cM@_L=_84D(L3MYa1(=d+b(\ae-e,@W^V]9>H
T)3GecK^Y-.@e;?JX?MT[2f\4E8d-K8b&8(Y(eT]D,_6<,>U.U;HIH2-E>):fQKU
7W@L/E_XJ_+2F>;N[d/:/(-/Yb(ZS6&g=;FUfVDX9OC&a3)gbVNFZ.fVM:X_95A,
L:cFC@N=]K5-4c:,&VK\K6ANbMKb3_,76>R]e:):DQ=4&/^?ZOLS\NE1b/PHS4-g
O&g/QTT0C.V>X>C9H8A/+H-<U#CKNQgP?Nb5fPGB76I]CQNLQYHA/JCG+RaZFO+4
.S48=\=/<DHCeM8.)SIHAC)S;LY)aQ/b;CGF\JO7KX7YSg5a)LML#<2,BJ42f5Q-
>U[;W-]S@:Z]A&\fEdX-e(R]RfDDJ6(4PDR3P:_>H6OA)V]2]U@9NW-YSW-@:)@E
^cXA?_,KVc9#0D>^?3(B3g/AD69I7WTV1gWX:-TX\PbF-S^YUS/,:c5PH0_[#f]C
?L^XeVMGP6:53#GGU8@2640JZ91[S1@RD(P]SMFRBT=Ab4fW8#4@dK>^UbFANB2N
JBCd9?Db??aD5JcHV/@@#J?_7KK[5>1V,)4\O<JWZ/f4gS?L@A0M=DVa#5/(Tf1[
+X3[M>^^ceYR)g+DRBUU:?V99@LbZSR=20G2A(#W-9J&5d>VIK(A2TbF1=?/^ggX
_VEEdTVB10^EV)\8LZ>J5=c?Y66\f.;RM,W-MF+SXBB,CC#_22d\4Z[=.>IM;]M?
S@;E)&[:XcbQ&9@=Y@.<WJbNZYJ]/28DV+Ef+T6BRCN#D,F>1L11ND\NNB[IaO39
(IEgD0<ICe78eC?bNM.QS=8.6)2K8[>#P?6R<-=269G2]bX[88@&CZ]PU6K,ZOH=
/[RHeD_H8O82@FKaCVN_QHW](6NE#P[\-T1?[9F_)<(.3OO08B6E781.T?6_M9gg
L89+N6V>6S0c;(_3c_JYKH=:896+,.ED[LT(g;:VU61@8#bB\VW].cW(f<YWbWWA
73a.>R,MC0Q>>F6Zcg;S@1Ke)fUI0S,/,S0]G@.]KUgKS3.R=U;59.+LZ_KA(F@B
,K/[6a=&ZPIBUW/\\7D)6;CW/V/>PXbRaadDKD6I-<?&62Y#XTBV[-fR\1f.]DD0
-c,YeT>f\?<CR1#75AJf-RZLU:)1BQY>HZV6)-cY(YVLH315#.d-0M/aQJJ4O-=V
0^#fV^H^=:b,FCX&3#Nf<XfYZ.3+M@.bZS;GfL1_c3+W,T,\CZOG=?#-650cO+S;
ZB=bN7T^8LH;3&-3<4(;;5ID@KG,/;;;:/>EZT?:Rf2\<c#/KSP_LP5;\PBa-]#c
54R8WaTV#Ga1OX\K-1FfdR-:R3HNLAKS9$
`endprotected
                    
`protected
&K\5^,g^T2RC\fNT[)>ebLTPc)=24KYc(ZN1>+,I[2cEA^f/+@DV()G]W3H2M1-^
O45JX0<=@1/C-$
`endprotected


//vcs_lic_vip_protect
  `protected
b-1X]P-A0bPJKeEL<FOI@5U\-&[<]9;ZW.F:>8O>A.b]50<KRINQ((+c^8IIYYV6
DB_5Ua:(CE36@S.LE]>0AX5-dH.\5BKB;=dMLHK]g]7YK\YaE6L>f>.30)/PO\?.
bTF[-]dg:.JFbT^4CXcNN<SE6B9(I<Z/W(KFD1RUa_TFKHK]\V]R+B88fA/FN>gO
Vdef/Xg=>V>.,O]PK\W]E,c[4-P<1GUF7Me9&;@I>8(0-R84.gJI<0,\,[c89Ued
OB05#Ne;U_[=MYH^O(e@2O:6gMJ8\DXTO&+@ZL4Pd:XAJ0XE)@+#XDG.WX>JXDBV
egD=_ebf:;4D+36PUO.M/da,G1HeBJ;KSOZ:SCSK-\c\_B&Acc:AHM/A-.=eUPFP
MMVN+f_AOCL:5NX5EI9T57GZV<a9.IXJ[6R2/&:P^[g0F4N?<O2(&]]dI=)9KB4a
T]1>=Z([T(Y/4DHLGY>GWc+6RfHJIVUM@^2GMP[AJfQ@KBcVeFFaULI-J<QS@2UU
V#C\YYEO+9XLeJ@UJMRW3C&2(K53XdO0,)F8fP:-;UE^0U)fJ#=dgX@.WZdbEa-8
bV4bEWM]X;W3M:3:2dHPX_Xd#2N_@+]9V+)0L[ZfdcB785LP9Q4cR#U2C?MAd1(/
V]JI)D8?ce#@<-A\LEO6F7=_g:CEc.KSG,5..<K5K@OC0>fB;8-MU5L57fK3L&/F
:W(Bca?9\=/<\I[-OO[XYE#5)..@_6R_VaG6Y=@<_G1H0KUaE?<1Wf(CY4eeTVR^
U.d-J3@QYAX?#HBB/:6HP5O1VBW&+RZP@Gee9UY;L+\36FE5AX+[cR:c1?W;+Q:G
E9:Z00F-;0)=;5;:]G;YCN^V\L^aAc_?D-M>Z\aS1aT-/O8c<1<67fcCBc\?B;Ag
_L@;0S6B.d]aG#=>@9-NdO9)7WGBPG=5+4>4N[O^gQU55B6UPTCWTcAY/aIQ_5O-
X(1;P)M<MG[?.VSB7eH:FZED:NX:3R4/RO(5SLAEM##eWLgZE_TZb/^bPU@K_UYg
]=PAX<C;?L9UTB84X28567BfeUAa#d]M\MH?>C0/,,]C<]086,_I6GdDTQ3[8^9f
D?:\g)-CNWfBb3:-TJQ8fB_[fLKR\^/(XBJ4HD/9FHSHBSUL0T1@]EUODF/[>VA.
8?/\I;\<,UMEEgURBA::aF@C5FRPW>C\ZeWceG?CRWZ;@3KI<;WCL^F941Y0+X7M
_QL/GL=Y)\@8TFQ@@BU>OI1&Lc,PZ?:WU8b+)84GWd)e-,>ZGXZ8TW8F]_JG?W.9
RSRRVIT+D@#PXO3c#@N6ANK>_C58[POaZGO.9CV25@[<\03(6KJc3N8e.UKX,O7.
U?G/aE\MLZ5R6C01A?DWJ5\\DK7,_G3L4EOFD2cdE(]cd20>A948VTTI)e,[aT0T
OM1X=.#+,aa&\^#8,ZO6/X@LFa8>eY3;5dV#7e)&O08Lee422\cN99dO_a.8NS4:
c&8J93(N[465G.(QL_&K>4<,Cd(/@(Y=5(3AH;A,R2ZKVE2+F?GU^Z=AAR#<&[b2
M8B@2YVKMRg>B.2C64cM8Je:?GXbdR7GJUUH0Q[YV/V=&B+\?aIEMP=g0E0M<ZLG
H=S#UOb(F_b7/)(c_\J8^A_>/>H07ReEC)(CF6f9da812^S96/a&)?ZSgH9N9XQg
TU?(OUIK199>V:9H:?AH__OLNOVYUI36g:.-f-:9<-:K2NU(A=@b11->2D//DTMF
BC\3c818]LE]6:B=4:C?_QY[4._FB_63L9-(5(Pa=:eb.]Q\c;5Z_DS8a174+SFA
b(b2LSNQ=(R>aK90G3>PdCa#4VYMWT]I,TXA#D^PW\>>T<)fJaRAC#SP_:9UfBXe
HK;b-],0_M^4RM?d1BU6=gU8&>^>3+]X89)Ra-,,C<V/#53C)^FXIV.Ib/gSaTC2
\8U.,^/HV95S;,[LP.<JV;^34/H^e<]7HE,SV\LQ[5af+N8:#V>M<gGYE]FN1#;M
YMU<DbCKTg<(bT=31[B-M^QcB_.J>[JGV>-0&.95LH.JJ=G;4;N=aAe45P([cNX4
JMMXZ8D?W75L#?.A4_3?bE;]T3d#VIH,A1^2gIEYe..HHZcb7NBgJXVZ?0JW?9&@
&6_da,7HeJ@7/-7-(1fXO-WXDBb/7HM5T2Y-46KU,Of+<-1Q77Oa7e7#R#P?d+TR
Q&,[g@6WA7g+T3AB@3\WRc_^EXQ;J>8_-_,68c/E8BC2FVGND3+Pa^G.daWf,b[d
_ggV],;D.O[X=dP]_a,0X>TcJ3PYL?\_JR3U\:,^GQD>_FALMX^JCWI4)ZLPTH(@
:^Vd198X2?8aada?BZg\=0JIHUdX5P<_&NB+:MfC8@/C1ST=M_(a(;A]CC7Z)60+
e(ZX\dOB=F,.PHRQ84f91+RHS+H/M]eefJ#H+M]B5=X#N#1b/;QS.2:29a,Kfe/a
RF(5VI6U;)_D&fA5MOF<AK@+@O<O>TLETL4E2A3#Vd8d;JO4e897]1R0R]:X)]XW
S8_g]RdTA?U<0P=3cJC0RVf<&77SC/RZ2LS,Y4P/H<A))3GdGD:&9fK>L]2_D4P-
?G)g4,(1\,aEK^GGILQ[3=&XN&T3(58:K(+SG]&9X^.RVfdNe8SeGaA##&:6)Qba
aK3S0fgEANQH,0&EWR7(<J#KI#Bf[AQ_]9-VegdcT)PF8Q01O::.Q)Y&3_:KRKGb
A^HMRe&Y-AH/L13E[N@QS_K,G1M(XT]7XI(aJXZ(@G)9\ZOB0^9cR6H(#RLD4GPV
617F]S<7L>N5-63a4^N63;KJ(7A<7fHaM<]G,6P;WJH59@OIKJ=_:I:GMa>:C<DU
cR)=D_8:054J4Ta_CXbK@H>IW=.T[IH?1CSKPQ;fR>2R=^(]HT(VI<=F;H:FWfG0
W<?(-IKbCK<81;]8LKgT2V=a#Q27<ba2d0/NI93JJ8E&2DM[H6@8,Z6OYGC(C6WJ
^,Z=;?f6?#ea5P(/SO;9YAgQ#a4E^E8-[/Y.OO6.VA16\(Wb;_Je]SD@QLBf]5=N
&[bNI6Q_Mg7F4aI#:cd5M@@9b1?]B0AWRZJV8V6I0BYW;6(CQD=9@<L4?1SE8-(9
L<&8TDdTEG)0_eO[cF>LESZbWQbKHSVa>>10+:X_6J^DVf=P&A=..MR(G99R9K?d
>:,@LD-.c_+O@EK@@WAR2\)DVK5^,VX+Q1#3S]W85AV.H&:RdJ>M/F^I9/1F-2DM
_WT0_[0d<U(^PZe)H@)+f.OJ;F,b,?U1A@/dCSESZ[5YL=121c30OJ=#5Eb\?O->
_ZZ5e,bAb^-bU\8QANNHF5DYCb<^V&7V8L./>Y2=+eP0[>O#+.Ge0KGHT-dBe^PV
0a5\W)(c0].;OE&P^aI&bd[UF.Fg^^ND13PWEa(L_APBGZ<G.5/eJ[W4]?)2.&gd
(B_.X32c\^eXT)CKC^aG[?D<KX33/\KC[PE(JEXR=9[+P(@H+OO\2IEDE@dgOAD(
E]c#][_@fA=YUfSWVdI_RS\9g2(9dL9MdVMP[[FWCGHK<f63;-dYOG&]SM.BL9;g
W;V@N+2Fc#c)Q5IO?ab2:GgF6AF8g3a8,aDPLKc+^=XYX#3/G&26;YCFbQ<0X.I2
FgSRO,RbD)FRRfN_VE5DL-.?#MVQUGI,TKg;=P(ISV9eZ.P>]+=3,Ug;TBPf1BF=
fCH#P@e)T,b4X,bZDcLUEEC/ES4[44<V]V8f7M;_H00U(NA:A?V/@fB[0+aW>Q@/
1+FcA]beF>SM6HN/8JTM5b@/Y2aWH+NCX9(4NcIJEMMMI8/\(B5/QV].JJJPF0Q\
Zc)c^XWFTP@=,;.NIMZ/Q5dW3KKL))69<cX/:DJ-=V25)J(9CcPCI-_+/-&?(,[.
A5Hf6aZ4O1eE<Da,4^(L[+YTeZ#O^V2UMg>I45bF[]@3eKd/Q7TdL3P59&.E_QVe
Y[]#P4M<]Lec26#(#TX]+>_E=_D0ZG,]6X/(#ZZL2G\a5NV08HK^.?^>9UEd5H(N
Z^G_&^1RM57V:Q8b&gK[;Y9/1(7G(fKAg\-=(#59\b>3ZW^?0^HdW#\AaIID+Tf>
7>?G#T+LVX0F>PF@0^3C>2WfO]J:09aN@J=\Q6;OMA_687<J>)a-M.6;FY)E)>JU
4&EQQ6.3=X;H#UH6g\e22ET^cACU6[ZcFQ^d_H]\:9^W)7:]>JgA<T+0ZS6?5I(9
@_a^\(a=7@NL?Q,ePeRe@?;X2UPR],[UFEJW&a4F&K\MfGg4?E773[;B]6a_2da5
_1<4KMBU;PBac_91c6M8[WZ^?SCK3A:Vc5gC?4aX-cXK-[0;D)UL(e=.(E_;FC#_
8/W\1SGNaaAbL2:^B@L]WcQC91ZP=D?IQOOY-@4WSU+LF22E5,QZGE=&QDNXU,]V
Mb/@Y?O5\J?)3\[eaWR-BMTAUR)<0T[S0]S;A@Z4?eO#@XIO:VZOSSU=+UX:?GXb
O9994Z;@ED4XG5)=.T7.,(d[]#G6Tc+fD@D<G,g]cECQK>?\L.UR/G[#L3Z>0f\3
Y[4+Y#3;<L_[1#&>4:5ca=,I;7fTE[WYAOCeDF]87E^[QVWb3b0/ML\_W5>5\:0+
cC@2SF.YGA\&DZ4bUCa]EHH883_V?2,9HP.:PbF[a[dY(H+-D5^3<f]?L.HUBB4E
8.L:+@b^eLL2UHEfKS/,V&OaIS[g[L+>N@9YgN,@IHVf&3Cc-8VaRZ,;]^61^82G
[ecR:_C/)2>HTZ:deAe/65<LHOAJ\JSKBg#0[HgHB@1WWFIZMC=)eC6VZ45&M;W.
>F/\\_H9DVbd;KI_d66L@2F)KKY\-:3b76PQ^UB)RJP6d88YO@GFC&)M:0FF&E0.
:d-?XWY=VU(:^=gCVeX./<dM16[-<cIEW(7:_,<&>1E3[V<5-^<W0YHaEf+a8+H&
cXN;5O.0=XZ.QZ0USf_(b_eKD(&&AKc2+Ic7a-)_c8]8\:Y-5ZfQ&3^QcJ(N820Z
)>W)C?HMWb3]VY]+CX&Ye54C&<?bA\UQ29^W&_TF1B<Q#><2_T7V6EL#Hc.Y=]#Z
D[WQWRGL/#W\#I>2I:2V(J5Uab;9FKd6@E<?.OB0?[P^M8<S\T0T0ZfG.HYO0/^3
U,&gR<8L^36cBG-W^@AY=>@Ld:)B:@+=OS45H^\B+dGMOE^_7ZD?=>?f9(:7C/(N
D^M3=;FKPf5\bVBf#,.\0?Z/AO:L?E^<1C1_Qb+=P9A;]RI0:I#Wd\e630LHE@NY
1PB+OBTcH.G.4BEB<LggNA6R5g>IL_P/PL<Z.N41LHH;ZR:PL@3Ee0U_E+ID#LE[
gaU#6/c,ZUR-_,^6XFQgD56YJ6?4UI+g>J@9d:XBa(MST(HW9R0OTS+P:/f>R82P
W9K1gNaU\SLQFWR1VK)1S+;3JC@OA;C4NgSZb0d@BW;MN03+(d6YFMgAXAdc?S_;
dQ3:(,K<9eL(/,B.a;U2\cCYe06dH&X/Q..>2OSR.EKC8Wf5X^MZPZ6^>IPD??+-
D+;FPcJF6(<(CBb4L@@eG2HE<X_9V4F1-]2PPPYWKJM0=+(:gG:L150/Ub3b7gYT
GbFS)FbSAR?eD7W],Ca#^\RN)d?]?4E[<gc9R8JE/WKH==-?RT-DOUJ^/FOKN0_K
C\NP(PPBA2:\T##J[:USN?9&40ODY@:2=e49:SIe1<L^>Z.UcL65WPTF-@B5R=7/
DVD)TdZEbZ06c8+WcW3=.0c@]A1=G@71H^\0BY<6BUEbIFd7d>.&[GZ;D@D:IHBU
Q2@41JNT@_J=W+43N0?a[E/b\9eCY/X@D+\?@[SZ2I@0e?:-aN>FU)Y=1IO-+TSJ
VQ<SYU^#TgC2SKQ7_78W/>gbB)I>L3c&gOP;_IWGS,7MX^9<XVGGD2UEg.(C[F2H
3f9g@/JeOPM8AeL_>(&DT2>cd8f.4P&C.K:JB<@1=aX50V&94f+@+TgVg3aa\K2X
#\.TUC,\P0.:=AH3=XA9[EO^9M1XQ2C;Kc4P0,7G31Ff7YdPAdCT])B?WDFe6V)Z
D&9L2Y^5.)a6;.HB_A9.=6PJB/JLB]e4Z_c^;?)CQ<g,AFR3fe(+:XVVUL1-IL?.
V9(Xc8QFQb5I>ARPU^[Xd8Cfg7884ZJ#F>;/41-U?#:c8b_(@0?:KZL/0QZ;47PA
.9dH:TT0KNBNZZf5a<7=HSaCUDA\1P:OYcbSKN/:fI>=DB6f7f9Bd#Be9^D=P(bY
U=HQY\\E/QcECH7ONbB^4/A25=>W&g]>V171K.DF[JVK-L(-ZaH]#N&FH;KVSf7S
R0\CK)ee5#9Q^3Kb&5F,bY>d&Y][B\Pcg60WbT[1I.W\U7MQ>5[(10KZR;:f;=PQ
JJMK;[C>HeMDY@)/_8\?/FQ@,18/<GSY--.\RV)f9=O,UgG@=4JT@1#-AQ;8XbXA
gRZL+;P259&\0XFET,R7)(b<XV3;\3VI<e#9SMI;ZeZ+Lc&UHHL0@)_FfVA?Q;:D
E]cEG@ff)S),b)QdbM;TDG?b]]S+a5BV#VJOcg>d:[\@B2d:DB+1Z?O>L7ALO#W&
LYYQLW9Pf+O.L#7g.]VNKQ<K@9Y)8T1PZ,W46.:]a,R.?TXA7gRgVBZSaE.=V67C
<](7XDYA:),\FCHMT8YL[7<,]H.^fQ,V0BL\Q/O/V9G+5##OfQF=D[4/V^U#6fB.
YaA_GM\&<R2U+CEf:/aeN:=/Uc_Id5+4QH&RUfP/K:SOP6AFU2E_/Z8TJZP5QMZT
\(5FAD:INL15a,L&bCRNg^Xef/I[>TJb7WS.9CMC5(YS+2K?+W&PQCYZKWAF8/d/
cX\a@U)/cbUX[f6T4WGe7X9;/9(2McWH:I-?5YJ,Eff<J(4?WeZQ9)2Ia>B<X>DL
KfAI8cJ8?29f4Z:d>f@/D3_HD:W<@9bbT;I]]Z3_W][8AddZc:5.1;feQ:UMLR/G
aVdVCc/S=3&5<9dJ=fQSaUFXY+MfRMJ0.SDVK^L9TdX5A6VV.-@>AH&&+0(eP_35
LV0UHCa306C5RB+33^##ga@R]59^R\T;6U7e3RU.C)Tc^1gSc=7fK2?WG#\T0UPE
]PLONZ@]Z/-[PY-C]LSD[7:1b[eZ3?UE,BcR8.?73A01K>+\)IGe-UUcHT(9QSR_
;#e[C_1Za1U9KPRYX[HaO-?4/MHP16=CYQf>#=/9WF-\@)bH09_b+f)&df<>=G2P
CIK,dGR<NNSTCadBEA,K@<#RTY9eQNgZ]6,I.Ta97&U7>&<G-6RX]VHM[04#bE]a
.R3H65(1b3O2X#8JB(D<JT_9MY#Mg@@-7F,dMd#8JQL[&U5STa@5dI+PKO3gUX7,
E;PKSF-NNdFc<TgP&36O&(X:9_;aEXa00XC?Q<ZPg;G2/Ecd)^=)2MOB4X;F[K]A
L)K<UT70E83S6]2KW#76eHX<]Y5a?G\G91HV#RP,gfPY:N:P1)9:99bGJ.g8<18c
)LEY=>]AEBAN8cU&G/d=2I;Ja[6Q/dZ.SCH@P3.R0I1U0f&X+R3MNeO?\KgU\C/K
)e+[ZP8CG@PNaHVO[]1^=b[e+=De#-AQ_a47NW<EW0e>WG-.<5DRA[=>F.P1RP>#
H:HD3<#dg1^5\R>DH,<V<.+LG+DA@SC,F72Z(B^(CacZ6g<;4_7^P.OXeV;UcN3D
&]S0F+,Fb=UJX89L^OK8^(@-Y82?;TaaG;^L/<4\[[N\.Zg@&GJFMF-.2S#:T24Y
L@G>+WcIU\?2/aEL8d-[0Y<)d\.FMC.2=]8NOg7UW@g26P3.#I[DI81+O/)#FJOg
ecgX8VSW61V:BXa.VbM:KGRNM>17dJ^M2<b?aUA\DS/a5ZATZOdDW-=3gY,FP_V^
?R^gZ//@e+OKUegOG3dY6^#LGI)T,QBd_1bDgGU.Q6P=@Ug3bEK3#>]DD#WcD#,a
H8HJ5G^]aBWT<;6O)+GZ\V.AaY8BGM:/V:fX-bP0<5O5WM_^6?-;e(-OU?7R26(Y
A\:ced85YD/GE-@#;d.c6^.O^1O#]7+?1.-BG:BeRXWL^g12bgV:b.9&FDC4,c9+
FRLP5CEdMeV1GR-.9?9+5^8AQ]R-7J3Z6_9Z/XJ4Y_DHI6eO=A39DT[<ZUTG9\dQ
af<U/BLUR^K1<7=__8e<=Md,=.BdDBdX?=c(0OOb_c(RF893(DU.CBf1&1R:;?[9
HBEH9^[V[(0FG5:=6<N@4XZMMJ=/QG]61f<HbW+\1;[EG&J83dTdd7<KKY?H2(AO
5a?S(d3IU(<U&/e2_R49DVgYYBKDcV(5A6]HeZcW10]UUeO[4SL6;Va6)]N=,3TT
YY0IaEDY?81G\@<L#c=7a1<BI65U,gJ[VT-aSIeB6BX>3c;6c8T8YLQY/eF9Dc^M
CN@GWMAbJK6=G(4gX,_AHMDFI>WSKH>b9[Nf7_4^)9,=.-gdRPZ4BJ=7,>bcUG6<
,2QeGMB=c+FPdAeX3LR8AY#-TKS)8AY43(?d:#PBAgPdb[<M>3<:EF]Gc,?3A_A2
\.JNVGX,aG0\LCF6(b83N5F>C6eWOcCBaJe\IPb30B5AKaaS<R_3Y[IL@#9NYFgc
Y[V-bLJB3]H>41+I?XdODF1@9c[ccTSI)46Q67QE;G(AF<RH:3;Q(O.8YBH_X:Ka
]J7XEN,:(U<>OZNC>I8K8:+gR7/7b?&J>S:R^_0Z0&+.EERLc\_e5-\O,Lc3K</N
Y.QY+2X&L/,@Uc37[5GZN.]E[:>#/2F@fBJQSXC?B_ZT0#DSPO?#Of4D1Ja;b2?H
JE?/Z\aWQ^49N/_Q_(^A/B]D/.;.MdJa;\2D@0?)I^M?&J<^DeD?40K_&&XPS:..
eM(#f&C:/[_-U-1#_Z:(16^PVWR9.AHgUcT+96c?J#cVKOQ9.I5e>(I+4#L[D_7\
UK8Z71eG0DF_f1/()&Zc>J?NX0gL)#1^bYZ64=-CY/<@Db\:F?RZCa,]<QW[<5Q4
85[a68>S-F8(1L],U#=Q73]eO=E>URUHWg5Wf;H8KJ)aOUc&GX^^))EPMa1MBbO(
R<NYb=)XJfYV>H([LU/42.K5Z&F]P=XVG68@_:]K(Tc>O<SZ\Nc=#-KFW#=W2Se;
3d)-.@PP?+X<.O-RB&)2PIKTK_Zb0bKQ43Ud4a?#>\>;FJW\.QS,S/a^RQFQ)&cY
_L1UZOAbAOM\ITRXK^63_.S2?AR=YERG?5MSWaU>fEIG7UF2LA<?dW6.W(agEae,
6X-8@b;)NA?8aa?)>8)LB4W__C(:Q,=1R&&X/,Z4@P-.=a2:g-1JI>]/0SM#.3b5
LU6?GAJ1?O/K\EGD\=a2)\dP3bLFRbMW6HT(bE^XE?LRKW[ESDIAQ=&,LH=8HSSG
OYaIC,OR64LN&K19F+CVCH=[RcWOK=]5H)_@1<7>T1=91WgOEg7cL]\BR=da:[5W
f3BM91,;(,/Q,M>K,TJdX(K5&dH[+8D+)4K]SN<Y2RMeAb+C>Z.G<fI1X)S2_G)F
USL^7FMWALIG,&I@7+<C+68>UCg(65B^(eF-bHM91I,Ge131K3P<;27.QHT=T(,C
&5TVS4b^Pc<Og8@-]XE:J:1TR](T=J]?BL3K@9JYfX918.S=f-[eYKZ1X2#Z:a,F
YATT7eXgM[_(TZOD3:Aa:+]^\+X[[@Cea7#[=H.2\g-c5^\AU4;GEHL(dPE0Y_^-
2aVQM^eA1d\PATJ2LZ3ZcQXC\7PV+6RdIV&@^/bd;Y(^X#1)/Y=UZZ>B7g+8UP,#
Q09aP.-D/X)+cKV]YXd?:-K6:.1)K-/-VL;Cg9:;^,M3g1e)AJ\4)0gBJS2A,Ggg
-AE@S=EJBV.Wa3>WBEWaHJ2e].=c4GDX#1b=]JQ.ba+L-eD@[3HQ/3d<^AR(P.UY
eSRe1&/a=\cKE=,be?S5-0Tg[.Y<Y?_P,3-KP;&.5a>O&A0f>(0\5I<2IR3IaG)F
7H/[38_Z?;d\>Ue/=?F0\Q1TN>5YI^&-NM[4I>L/JS@CbJL[Q6+e80d&gHbT3<(G
ZfNH9AZUaOcU=.RZTe/<3RJ_J,Q<BRPQ^7cb;&S)FO.F8De)=9_\#0AA(]Y6&/UY
eE(I5+UacE(8ZB],ZdSILEUEJBYZ\f<>F.RIM3K)aCaMS4\Y2)aAFL.f3A]=\^-K
S8A5+ETLF@QS(]?5939Nb0dC1VdaH:Xabg2F15V3+O5OUZ8GI3SI4YXW5?GK-gW;
(d)3NC;NSLXf#H)MQ]Jf6\]9#5U)&08B3eS,1H^2;L&(#6PK<JO-\F7A;?;601ab
=TBcf3HEQ[gSOF9Cd\g+G)M&8?./C&1D;c<T0?e8fFB\4+9:V,<#0_J;YZZ,#?AY
9^0VI>Ub_DK3A.\)-Z5FeU4fb[?BSNY:3]^S,e+PZ,Zd_[+=e8M3S\<dL?AV2Z)N
(geMbS#b/\3AH/a7Q&3RF;&23JL251a0U3PIRM<1-1b4ZB4)#48@=AC84PV]c?+<
=<KO(JD,(+S2^]VC4J;N\JaZ#LW7&Y#SZ+VC/f?:b>1)TMS_)VXM@<98^0DSU2cK
LA:1@JRffI70A98U;D6]RCXIKcM[SC^Fa#]+.VYg[>,Pg1G&INT4P3KgXU]2;T,N
(&E_@GHd6NY2d;E@FT7#3,N@F6f7b,^IVUX1A@_PBOUKJF?J65Kc&(ODBXIK<M]#
E;D+5]fLLLN@cNSf_9,_+f/^b;_^fG)a]F9DEZcUcKS46R0b0K<TEJAAA3:@J9K-
d_2]9QK6J.<^YTD<[C[TERRS:F>)FQDcPQaUbU@5#0LZ<YWEdJS\]PQg?M^4>>[K
R#?7GA#XfG[b=GedaeKOM1&>+^((b_C)XS4O2B?:ULR/93aUeBdOSA2g:d5:>#79
cYX:F;@LI^S@eA<NPaO^bR:95^MXA^g0>XV0/I>+(&].\WI2#5CX7]06^OA>cS+=
MQ=b=c2084Y[\(<P-(3^;\1T206UFO//X@?Q5X&E+VT@K=,3\GfcbCB(?02+gAIB
YN0-bYB_0U5[&Gg?Ad;WO9HHd#W>C[/.C7-BVg62E4\+12/.9&UN22H5IIRZ[4+_
e/PM4g4Z^K8UggEX@:D,.1C2,54J46cO,&8A+eZ1+GP1#\Z^>^LRAWg&\GO;TOg<
SHcF9)=?g9gOA+f6QU^A+HY5[]CT-Qe2g2(Z@5#Q=MN8Q(g7.2B#Dg99ZJZHY]Da
b,@ZadL8A<TfcM\N[&PONL>gN&d:D>W-QJdcHMcF&MMcMge&)g+OZ+TWH;5g=,.6
Q5;[Ff417);7))3T>SY./L3#NAZ3V>AK]IcfDUc>bdbLOg5@f\_0F7ZJBLgQDGTA
SdaFcA8b,TD5SYUR0V\\4Y<6W,-S5A=@Xa.EB[Oc5AD335+&&9cW+gdEGD+O0^d\
a<_[QF7;5aQ.&,Bc?_+QJ+;g3I^Ed=,Ee2c8a8Ha#QEdEd?Q24<>J(DGNAfe4:68
g[RH9KUSQecf5fUPdDO=Ub0BJ_\+0OU+RQ2@9SZ]LdUA&\4#E1bfU7M&@C<K2DWG
cU86^a7I?IK&L2UF;)a2#P>3N[Z&AXafWT/2A9BY65K5=JJ1g]HR,aR(8XF56+XD
6;@.Y?6)C<2^RbI&B+3ASZR&MfTC8HVNd1M=^(0?J&IVB/?7UMAPA#C80WX@0(Y]
f=BL?BB,f@KZ>.,9/a<C3?DVX,-TFG?+RJ,937VbX\N7GX]VXBE=U[AfBfX)NL.;
5A\e9H_5=?H+F>49)gf,D>7(@>[^c2UTRUL)Xa3BHE/R);N590ZIg>DSS8]fI>8-
,SKU4d\H^T=K)NH0a,&]#NZ):O;O(AaT]M7P4UHgNO+>@>QK1/./K@WO+9=L.;7(
f^6P(:HA:O<V58B#bER:P&#;J-_+T/_I/F-Uc]UQ3AgX4VS][F^a3b8:-..G_V<S
APdTV.GLS])G8]SK)DNGW^B:&=9>J#F?B7L\:F2@&9(2#B5CR\COJbH:\7-[:5LQ
JA8c5/1S;3INcK1=Q5\?+faYedZ/cG-?MF<4J:8/Y[)U#ZHON4WbQdQ.I3/VG9G2
Fcab<1+8@KS]J/agZ<dG[INBIM</[K2gCN^.c^\d.3^=LQbU?E@5.(5;L(839#\Y
8,,B=0[EJ>aN?30U8+)=H2UdVV>7]B>PI#-<C=3d+PA4L2>d2eXS[5cXBg?[N())
[S9QF87G7;ZUfge2-(7MM@4X+D\EK@FVNF7[:=J&8^^LG;_Z)QD9>IV+-J20GGPC
;L2?/#G,CW.]AN]#L7N&N[OCgKFYH:aKF,3X;J0GKUaJY>BaVMZ9?+]=.&)T5)D/
LOQM>XT(03E(IQAb)ACKE9DV2V\__YbK\U\V=B3H^DO;W:Na]LK&XQ4);TOIMHIR
N(+5Rea,C5CIKG;XQU_SV&3NVV_LeD4\^UU,R>I.Re:S9D&^XJ7AC.SW-<Y?M)S5
V]d_SO#UIeGHUf.9aE>dNFG9A;K#9K1@;FSO68IPR9E(#d;a+1g_I6\JE^Y0E,58
[Gc&aWScZSM;:38VJ:Cb3UH3^C,57:DF2-:LZF)dGRg37:2Le73#YZX_eV;VJ]U8
F35Xeb(SY/D\ZaK)#5?M)2#T<1.B4>H-W.D\H>[GA22?2>ge)LC31T/[eWK#e+HV
QVCRXWG@0Q4bT(J7f@J\dKEW9gaC5R[beSGfBB^gVAJ1Q](#>]b:&RYb:[M70Y)E
FSTMO]3:F[87Z]a1:f+L\D[NKVP2EK1U0;?5&C_b.&a[M,4YDXQ\#cf:D=9[:IP<
?dJ<AcPC?AT-<O29LR-PRMICWRNeF9<>A;_T+)3Q&G)dD_(YB9g7JER<a/\?Mg<U
&cd@/[>g)d\WeFWC8TD>A[/J^MLf<9UC.K(,^;P0V\Z5H;?c9F(dQ@6_bO0R1EGR
8?V?;MM:]YL8?fd-,fHQC>PLNS=ND[-?[;Q<4+be^H_^4U?XMLPISa75R&Q6KM00
)/TI11VfG4)1=WI]DD\UgWN2B)FZd(ZI2cW_+]9&@ID)Oc+7329;<018\ZZY3_\b
6V:0[Y8(N/9[^8I@:==T]O((N3B@)5YZ#@;?-:NB;JU5gfQ/_HQL9;,/@B6W+#+C
]K(HXeI^/M;)3\=SdS(LMM;eJY5)]NPgd#e&(0:Z8?4aOJY@S]GQN2J61B]f09#@
Ud;,bRVSU&JQ;2fHNb^_DX9]0H=8:A>7,0RSY:7TMVL4LH[/?7BFcSKMOaYXOd,V
&g9LP_=FgF9_--+0+1?0GOD=I^\(QDeJ+6G<_\9W:a)00e#BP9QD6\EXVRR2#-3V
(7YO@&3&Z:=SFNU<)4A+8bZ3Q0g74^c[c;Ka/EbM[E4LQ12;72V:8ZX2HPaM&3UB
NA@.aK#3RP?.PJY,ABe1f:]Y-V\B0A?A)QVH]8N>cTWC_)^J\4T)02RKM/-Y>Z88
.9QUP.JIG5X.GBfQJe[-3g9;^TFR\aeG.L\]J/:^913&S>5Q]NTd.X5bJ;OD9X[F
=1eAB8;-23Dg=R&U-O:_e(:bIb9<SU.)JK^J5K_YUL5C_XDMA.KXga^02eTc+;MB
=V((<GJX\J=eK<2WbeNfM,fI3fI2KL7\;9(?@D&MRIL_-=6(V=de6/GZ9;XSb>7G
PY.M;XX#^TdJNDfAMMU?XCc<M44_.3HO;&TT&<bWM.?5,_DGR6ORSMY\4cRFF^Ve
&<Fag38_XPIdR.A^SBGR;IY]S]Mf^3\g<,D>c.)@,Lb_4=IPJ64M+=@/(F;_GIEG
#L,Wd>,?5Vf3-C_CdGI5Ua,K7CT9G1fcTETV2BALIeQ7B::G&?fU@9-686NP:?17
^,(VAd:g&&#C9MD,0U=L[ER6E6,&=9A1O-=KS.C1M>e\E[G]?J3g,N,CQgTd;<M6
6M&&#UbgN>G<XHHF?;59=4:7c>(a6/;?@cU4eXZQ(@b;Yd3=/_P6d7L1>a(cdE7A
gQeH<5O_RGW/=\a]ZI2RSLVGeG4(7M[QQC^G1MXeP/J/8\)#H9W7(S[J:5S[E(g<
M[8\N6/BIe20\4fR\B;fGQ?ZW1W/eU[]?7>M\/81O)28_@a^aV+JD+Z])T>Na#S=
M.SA,G=#cN719/<_WEIJ>U@GGIJ\Aa1(I_BR&c/F&8D@ca]_?8RWH5U;C^g9YP1L
I^KY7NVeg?+7A,4&6B?B@V],&J8T]F__GO]QLT?+Qf&-XB7](_CHFb<:WT:)7E2+
^)>A6[f>^[<]WVHN@b&FX-[G/g?\#E_cBb:9ZR^(8Q08A1J@.K_.[U4gdPS&b[c#
#a-4M?9cZ:cQBTNN>^Y]LP@+H1Xdf1KTXWONS8G\F:2&GObE/]?>(=ba4aTa>SZL
f[A_]Q,O>]c<&:,UT1NHgXRXW]F:3/aF\6?eTXTGJIG_bF5R>U;.F7ZIL)JEeeGP
E1#C;S,Y#0b]J-68D9;&U.^JOD#b;BATg5@;PI^S:\fF@A^(FD,,gT(AC3P/D\A7
T9:E?UgWT7-:Wg:OGcg&fEH6Oa^6MOQNPDa-:g^FPeIC835<B@OS?YR:A9H5e\Ja
2R]Q7&LKH>ZI+N93@^1ZA[_b0a=&:^\_GXU1XJ_VJ8>?C<8&a/gRF<IHV98.^OMd
TGFXI-?Z94R>\#ESFaTaa6aT76;:MGa?MU6CDIf2(3DeK(Qb8Wb;M5(A?e]\3)Db
V)9-PU54NWBcMHaM0O]:c^9UJ<dfUK5B7<KG96##UI2+LY2KU8H;+]ER-_6JV(5_
.HVOSYY6_)6Uf0SQ??bH9X<A-5:;gdg3,##F-g0bJY0W30^eR&/eJUZVcBBK)/)-
&9_VUEHA07NOS5A&K89CHWGQ0D/a.0c90=aO.?5F<4:(dW\E-1(Q/,b<LB7FNU;;
L6U4NO1(\S=97,V>F@IX,P_X;27dOIZ<JT[cD5WBMK&0cI_E:VE-V6.T]6>0[<-b
A;;#DE4ZZ@O1T5G=?f+IR,C3,J5M/M#\7)\BOYAIXDWN(ALZ/ZE:8a<^YUB)>V>H
ZU\;<7-WKI(T;@>DF\#dZ1+aEUAfb2_W=8VfJNDdOW0(2G8A(<&a3e(P>>(Y5Q[H
RS<S[bVF1Q\4O=]P&-f&6/P2RcgCfO]V),>J]M.,B_&T,=R6FNbc:Ce@5L@O6[3^
?U,2dad#)D-d4X7_^42D7IXBf#D=/aVKXRW[c.PX3WGf=9bDf1N,IbC5LK@U7TRG
1<SbggW+(HRR.KIE,gOHJQ5VUGd:1dXYL#1g&Y@eUWYGC>YY_;1.),-DWIY/d1J7
45G.J>>P@[-PEK8Q88ZHXD(7R163Nd\@?CLR+47Q.SB0;C>AeN\eGc-@]a+3H/T#
,1cG,6\6G]d(\=8K+53<+,H^20;bKdB=M8Q_bb&bP1[Lb3)GNdS)edL+7Vc1EJdY
,f\ePG9NXNU0F_BA;BG?bT62ae6#9[+<b5b8+[3gS&.cBHGb=:68M1R:^9a7>6:g
ZYURH=4UW/,8JIOTEd3F#dX?20_Zg&E(HJ;5:f@LCU9gL+)-UE)_;UX#-T,CTdPK
ReK]TIJa[MO=Y^>&D5((,RKUP<S\&PU]1CBbV7I8.==JIU>9JI[[ARSW]?NU-g+T
#T9.-)2();<Tf8,G\_WU7;Y0I.?X@&5PfQY>c;8@bb(BM=FNIGL@Fc(CeLK-U3?F
=_LOLNFP\^AK/+;8D,89#RR9\[FWEG.BGLfJ^//X.3#77^/1+:&9?]C2/B^(Pg@>
V9>.#B4J9C=(H]CG\T^Lf^JO4UC4K[e)0[G63+SY62E#DY3=+.fee27^&-T]RR8R
9eNb;@AG^d)CA[a\QcL]C#.BRc#BMNDb7Pf8@-<-R6F/^(>3c4CbQPdBG.R9S3>1
]cYAR;@8G7:=[-G@3QXKN9=9ecH25U]_JMD<\48YE):593a>NL6d:;+02@CdJJS&
II8+CW?5H[+/cQ7EH/]ANTKW2:[e1G4\#^.,gPRLBBJ;CdA^@H(,1f@V=N\,>@<0
PI0[eIH+7NF1&X,B/P.D&;:A<J:K;/:N6]SW7J9Pe#R)E5SFQg^Xe2HGW.C1>faD
J?_R;RH8BM[YBEHV/F^]]Xg2TBSP8cHd/R2M=#.Z6U=d_?Lf;H8fWQQDA/0+aX9D
;e2Wfd]8Fgc)HB530O8K^6XaO;/?SXC]c>A,d.-I_8FBK8/:F6?@K6?+Y8Rd:fUK
,NcJ+TYLfKS+=f/2AQ_I1g)R\.[^-f78FTbZJ0HC&e^2,T8WdDD&KaG=c9/ce\;&
T4<W3&4Y)fU>,1->892>4-A^dY;TQYdg&Sd(Y&N]RXI-SU4G/=Y)7M.NA#.+DEa.
X3VRQId7E538YLP(E>2UEdMV)OTgM-&F5JL/WO5E_f::&QAD)P;da,[YLRJRdHg+
Q+3-.9Vg>bMfR=733O[P)E]+R6?N38:NY@^A7-[GQIT]>?VA^_>YB4AZA(a\aF#e
A[A<:YS,Eb39&_g)(4WPVTS[WWbQDI2dU@E36\^ESU5\8?WD&gO)X:?H#]V1.\-=
J65dYeZ(Y+Z2@Za:0#=2Y<U?>b:@@+0fDN/+]JH?1??SB7MMP.JT5#I/?cbG2If:
(<f^[e94A@6RM/]L][Q=bZJe1ZNMQ/L^>D:bbL3G>g>.2GMXN;X>-YS]/=g=gN&A
Y?=Y&Y?S#GL>Cf=E0I0^D#??,Ua&1/N#O(L0A]0f1T1PF+;L\0&:+cW4-(Q87F\V
KYgUE36g7EXL.PW7#[V#F_5]O2GX2N=:5UR)C9AW#a\^Q>8_8I?/N@3b,HebEK>X
::6I4YO>(:eK,JPeRBV-JS^>FB>fcdM:cL^\,c.N\<XV]8N.YD//TL+V#EP_VHT<
:_fZ2Cdb8^-a_Me;a+N&0TMHJf^0e)0U,J&UAWafBac;B:V\cF,Y.7+44_X:+L.f
PbT327MA4^a<F72BHE(B(XG&\A2ZaEZ-Ra)g-\/;^</[7=Z=bZcIM^UNe+a7f(c0
@+a9LWQ5UZ(9VI,9FE+7TUP](ZegHE/?_W2_)@gNPTc:[/&+6gNYUSW+MG+E]3S9
E;+D(_C2P8-KIJHQ30V;=^G4U<Y5V1b>XQM[]D9Ka.0^)6=Pd>>;UM<de?C<_X72
:#[L8eNA9R9INdD0,^;YV@:]eQX:.Wa0,.4Y9A>>Tc#CX2E&YV:SV]8.IG\F\M5S
0?>E:f5()VI@/V=d/&7eW7KTAZ4gP#S=b@5<7AD2/O_;@6#V8;&GE@C898D\8#Z,
=.&=cAf@f7^1M:RGGNGaJ9+,B])C@G0:LEU(>P>(2fa?aWB&d,NT2O(XSN(T&I@d
?Q18e5T4BQ7:V(OR3HYHddZ5Y8&W:9\=J]A(f_>#KMUPPCReDc2,<eV/PRBU/X?@
W#f.KdF2Gbb+JWD)81N63T;.eO6d4+-EBS6g\[Y-T^#.3)6b(=<XdVAAEG0O,+OI
QeaZY][IWH,9T.;EDM3f_;)I/SfICYAgUTffF=WXBTSf;9(g(YL_3^MG]9G:#/5c
4&b58\bY/<.:gbM@D+V=K]RI#_f6L#5EI/L?N)a1Gg#RSY_P/C2.0f\^[.Xd;I/a
NK9@d6^\HXG7NT97(_\6?\8_WgIG.g9<[c-Ka3a;Tbf@I?]@UdWD@fG_C7cG-/>T
SP61WBT(,QCGbY7K1NAb1?Cf)TAgFgHB;-eL[b<c;?dTHP>4?b@G-CW@0.+RC>[?
S;^WT7\GI/T?gRW8XJV8H&<b_;SY-gU[MYE+:A>0=IMVW<2O+M9EQT9M60fPS:>g
PKU=QIS&WY4@:#O?QW-I)XSTb369VOS[8G9R?1O]e^QfcS,R5@,FBD<4S+4c;+P@
MC0F6_-8FTe<I_-ZY)c4UR)+QR<B<gN3M/&R6Be&V+=T3WSe<M5@dXbaa90X2,L@
+E5X;]-P3C)]c-UVI0-AR0d6-1G:+STN1&R8gZ=N5I5Z&f8][C,dWW84#G8AR?a1
2&.-U>:>fI,2#AM^fW?74;L2e=A>W_I&a>GK+?@:5L:)8_0bQQeV##SP9O[A)X=W
c?I^9F;_<#V:OW5\ePe=Q&B/YVW1G/EdJH.S:bI?W5g+Rf=3dUYGXR,WggFdOU>_
Cf,e[\EJHf&)d4VT#;^>@>60DJ5)&SfQ,Y9MB,TEXM-I+V:E9W=e:DeAPg?40^5F
2.eW]ZeF8C]D3])M,IX<TQG7ZN#]S(1fS-^R\fa&bgB:863V#]G[[QQ;+(7Z6)Ib
TQgI=C^J9@cI_dA\W>PA.?>e^Q-CQ\?T7JCcF>XKNT;.B+dJ:GR-3c:HD;=\7^f4
Mg?S11DaD_Pd9b3]8Ldd[54;g1G?=^&7K3TZQ[#R2c(W]<(-7D63\3H9K@G05R\[
.B2\PHE5H(NRM&BP1:A7HO=-RXeU#(P]>P08\^g^Q:d<d3YY.?_#/US=-?KJ]:B:
BOJAU\DaK(G2CGL?b2.)d1>04&J-DA:@_9(cVQXSfB^C()<1N8<B-(M<FBHg-3B#
a.D@&<V0H/SIZ,<>6\ZRQW/MDYAM>I?>T-#AKB=Fe<VFa1\UABQCPELLAB[A41YS
7N2fKX(?SP]C\B[a=\:YeJ^dZ\HMgK919HWDMH6aPC]1(K))W>CS[(G9g(3ZI:)^
YKU#W4dS06H)>7J(EQS7:X6KH3PaeJLfD6C3>KWY]cCJ>)\34V/?-6_K:,V3B/)P
XfEF6X</;;UfM/KLRG1gJec\cJ:DR-?=6+;edY#<K.)JcUI5@2+;WB:2\+OC3<>3
cB_8.&Z)4d522#E63YIU2?BH:03PP<A&OI?^H2-+72+-(LN4GbJb2,d7eAQa=X]c
accZ2LE5babgS\c0ORWKFINV4BgW;aeC+b6<771Qa>0eUEK-70(FMJP3UR4K7[MB
I?,U\dWWJKCOAHBREe#)]0?\D4ZDBE\\129?;Hdf)=.Q1]=[BJ8Y8@\831YdQ23_
e3.2CYY#Z/RU8=JN,4HZE0b,/M7IE]@)RZ&W4^E)JF:JE[8,M(WgPD6=VFJcG.2V
V3,g(F+TeW3<LC45JPKN[f0ZHe<,?<)5.)6Z>;-d84JA8;D5d^8(AX43KXYFSf33
/V3]CQ0.<](Ve?&I[5ZOHI(Ee&6T^J..E4.97Od#dbXd^T7Z:6//WBK4XP<CL?B]
V=T4@e^Sc+\XK)1\UaK.;C+]5)/]-g]:NIg3Q&+:GZ1C1@\gfFb/,UD\<PRfERT@
3<DT/<cY5\Pb.K<S[H(Rd0C5+@Q-?G?&2=DQOC5K\.N)(21cQBf+@8&S@bCdP=;5
T:DM,U,XVe]TC+10/MAL]cMc[VU)+&2a]Ha+8FR?83JC.]eEEF]37b9@Z5[Z3\5:
:Y5DSDdg3)][#5CH>+&=-2eKP47C<.g^/_EeUHN.K>XFFP\[0Q0&E;2f^Hb)18X?
W3]&X2F4DZ.L-?.Y@8,JH>2.,8RB:_5.;,Q/8C42JS?,]PFA)YN1Vg3-,]/^AZ,a
45+90W()=ZCB_1g9@R:8L203:/ODN7.=:N[=IbOg#@CFI.^:b;Z4UcX_?2PRcDX=
Lf[N0_7=D39Z@Q(T)Z\E0SB0H)9+M@@_c>_VYU]/V-#QIVIXC@FMD.,6(XPI2W^@
I6W4SNJ8=;X:S[63SMG,c0-K..];f?D-Pdg@2,:T0a&WEY?4-RK><1V=ALg/A(JI
Q27LTf=adHDfD]FXJP2(+(>F5+@gK/6&ZCJ>\A^gVTNMd&7Ug4I#_)I/D>K)\CNO
cfCc@QYE:F1a+g@J\b6E7f6U7P,C=&[J?Dd_-PI=dBY5N(#cND\I::L?Ffd_fB^c
\dP7>,ZF3+Af5K93L<:V_.3+[?3Ug8X=,cc3-T[/I>:B2\8MPKHJ&5HU1(UGWX&5
<Vb6-HLc39ZaU9U+5C?-0)4>M)G+3?8Q774(2+]UGYL8dXPYS^P@:\fEe,T.58W_
XILVN/D20>Q//>(=)Ea+I^KR@1aUUO2(c[0EfGUUd)]=94::733f@&e22BVDb5W7
IffR(,2FFM3.ZBaA#Q/e^CFQ=6HDZg.>),[6Y8L2BEPF,&+0)O+)IOM7LC#@H_a]
#b<.6XC?VD0#a\8U&B;AN_6Ya]7[BIe/IeQ[.EScP9E.O4Zc^0^FFJ218OW>9B[G
g_EefY388MI@0X9Y\Q#5\?<?K9f-?Y0bUPJXL:^91IRB+=FL_Q=40A=-1I4<?<M#
-g5WBSaD;[bW_d8^<9S+SZ^a3[JPISNZ#18]ZIZ;J^+.Q+bN@V)1J2;]4V9;WJ-)
+QVHB_J=B:E(B4#dICgS>3[RF+,Z2816)LdH;X;e::/SMgRJ@;4EF0bMHAXGZ2Nf
aLN97#CN.cO3[A8\LP(eZ?d^:c6)^];&M/P4KHdLc-SQ8,/\_^=WbVG3<\382Q>U
_U2WWB_A(W_Y2,2+;#aCRCK8:J2,5_Z8A:[[Ca^A9;f[+V\:TO>YN.+OE(\1,Hf]
XSO;I^U60?HJ(2=b5a[OH:M;Y=DTP[2;H7Q)_URF>aERE9aSCKD,HP)?L6e4:Qg5
,I>MK(ZOAW62XPHE??NQ(;(A>^a_Ec).aB)(J)\M,_1A#gNJZ+.,36-V3Ma#)IgD
_eIDGObV=UEGS@f^]aHGUR/U^+\2^gUg+K</Mg]#?d.3e[V?dX82.+f+Q3F1&&>1
P(Hd2bVb,Ed3#7>8LXcRG2=[a<[Y94/I<N)?F.4REA>-9Ob=+C>,EPSU5fME&8VJ
1CH;7c3GG<\P5?K,L,g/HYO@=<gbXJ.C;#&gL?VbV3><2TKTK-5KG_VR7N8g]IR1
I==&I0TG3g45Z#8X+-9(8dJ-7S=9S4A4cgL+GFIJ<WCBfSfWa3321]6?Z(@a#Wf(
^Zd@f;&@]_g#?QI3b8^T?D>@<2g5OP/M1GVU6bD(YH8E0/,S:4NOYgC^C2LPPMUU
\.Ub#./KD<1VO7c_K5>@I)6Ya\;YMOfJ<fQR+dbV0L-^E0\0]?>=;d2LHS73.)9L
BS7XcK0CMX9JGFg(HU#>c,eM]21=S4DAB2TM<LMYN7N3/b_\92E2;;/&D5F9P4bb
TFJ\R73ASI(XBOWHM_0[L^YY1[[:a(_HF03NIbZA-Wb856Ya-2RdY&D7?D,,QdH/
?G2fgd^72R:]5NFL<@)\8W4]98\&f@f,[G;4=(,F9[3,06/S0J8_/b]OP1_/cRMR
(Xd&]Y/b44<7)19<2bF[#FL,11DTTF;JZ-16:8ZO50dMTZ@CW02/?5g^96^X>EJP
80K3adCc>024Pg-SW:0SNW-=LgbgR1+349^eIS_X<0,>I0JD5YQd+P@@9I/80EOD
(=+CG)-HMS8DZSNH7MK\VKI,fP-D(P[XUNF#.-\UVJ99@:]+>IB8<c,CaLXKBCD]
,,f6[4PF]L2]cOU6Y.@&QgfS[b#c<#N64QZ9a=OL-Y8)aR6_d:@XLW[8\_^d(DCd
F;/RF[<4J+,:fP&<)bT)NedaU+aZT0<EF,H8)+OLeHE-TR4]X@bHde:2V]5V_XRe
\7?C]6/BKECaJBJQ@Xd-TXb/HKG#>-^9^16/ef[2dg-DAAG(FG9?^^E3dC86aMU-
F?NRC#[Z/:01<ZPH9NE<e@4[(EWaS@>gX-2aZ5/@e9^2_V\^8baaYV<;C@?_NG26
<bcH&[7S1a1,M)a1fA)XY=XUK6S8WRbW_.8JUE.Y0-[;XP[+3A)JQN\4T&8X-e2?
QPR:d+A@>:P31T,.(<>]9;GX^-\2B9Y+\C[,?G_BJX1-.O/.(M[RZbV<XTfeAHBG
aXEK#1c7)dX^RDU-QVb<FSV89[LB/Wc?(cONWN^F;1?K.L9IcCRZ49P^Hed/\.8]
R/ebW-5+4UTYCLY,6T4<fNb5K9MV^J.^>939D_B[PO>7X#GS023--e/^6_)88@6c
&L[/:4BMN,gZ81d<3-]-GRg9QEN5=+gL<3OIf&/&NUI;E=LIXfL@-I:P#Z3;@J]e
XJPGf])]Z;4ID#PL<GW+:&IFMD4^BB5?E9I1fGBJ,(e-Vf+/LY<0@)eNWX(FZ&D&
QJ)dV,@&ac[aQ/6.+XC^V4VfP)fOY&/Kg3QaX1HK1QT88?-bH-T8H4FQNHYF(c3:
FP>,;RP2I^b^b)Ag=)JgcHYAGNB(MH5XEY#JG@W/:cIdZFN2\D-&^^S>Tb5\=)\E
OK=3I@@TgIJ<2WP8;,ZB]d)=UT&.XE?L^:VM7;&P[AA5QJYg/+eJ\HW9Ja11(NA^
fg1DL?2-DR\>W>)@^VT<ge5A<@:#BH?&>Qa+G3.;/_U<KNB4[OW@]X3#<_/f:.b^
-a(I.#VXQJYbAHTdT3LbGURKf9Nc<.SbZd65a-B<BQe)[c_O-#^@ND?JNf.&GL[J
G&/++eN1[8aEaR@QdP_6b+Z+b@MfI=dU[^N011DPW8QUHZ9c4JX6@ReA9,Y,UEOI
L0,VDAdT]?M5:CO<cHK#_9VKY>CX1LM?C3O;T2[O^I)H,(]W69M\Tfd1B5-SZ:\(
XL0Y_\a=4S@=/Z#OVD,7TUJDIKDCUR2(?VW-3(;GI<FXMTbC92BIVZ>^]/\>@YP.
YY<B(4#@cY\._@);+OG#:&ESg@POg.b7E56a,,R>,?1BVd-[c<HFK9AOS[fU6/^B
K#-?P-<RQZ[-.,PR2)?AQVb3@&),cWW#+gUI,SWV8EBMA/HMd<^-FODG\:[]T:G\
=5X1CJg76]]9-=/KQM6b6NW4SfYE3A2dD2(5;/_20,A]#OFLM/)N9JH;J95DFT_b
N>4N05S_]Y(>B09PJ/5@-C-7;_HJ0BDU39(5-17S8#(@GHLe7#.0.S;<-AI:6.0a
VeMKZI>U2Ee<5(DD^g][aXQ,LW[d@:fQ?KG]#,_bLOUXL-/cCT^\8_XXK7I8;MDY
3eSNI]D;YdPIgeA1@E,_=f8gXeK:RL;HZJ6fBL;<e5?MP]CaJI^#WL0CK]Y0-<G5
:A4^L1aJEEd;K4(K-,8SO?^e_#Ec+fc^5B@AXeEJ(Y/_A>#.OBE-#;?E8VM,[6H&
TU._.bdO=;fV?L39cV&Z8COSU0PcU_d@Y&fC;e3M[=QZYI>B]Q],)FW?I]VA2WG;
4#e5GZ9+T?CeV<K,7.5=_#U&S50^8MAZR/eIOB4(:X?gC]B:@BRD#P0>?+4CYKPc
IYC&HI=AWe[)eaQFE9-@b+&TN,)#[C^DOA#X4VA31E3RO=:DIGTC5_JZ?B4YKXVf
5>Ue.U>F0+_X.FOY1<c+Y/+J;,0<^IK5b=#VR)2]U=PS?EDF,FYUdKae)-+[3DOF
>7f[ES0@O0[U#:K,T5./X[cKaca9=[ea,WC&5/&V2U)8=7fP5??Qa8B,<URGFZRN
SY.#eg^a7580I8D&+N&NHfTYVgbVBa4L<WY2+3P4?TW/,U>E_L0-7e&T6FcaaN4-
SdJAW+B@Z,1Abad<?C[_D82B.E0K_\3I6&9&4bWQO,(:_2cHI2)2^\fN,ZaRRd2Q
?V9_N^IFLNN_.?)S,IQGd#)E3S#+cbdLK0K2^[C:BEHXd.R0B6aPNMT/1M<N[VW(
fOM>?AFO7832VTK^&S:35,+GMd,()LBQW[@T2bR@Wg7cWBAHec4aV?JfA@VN-Y+V
9-ON\2R-33A#_,YQ0N@EI5ZeOY,>,;&N##S=c3]..KE@:aNBE]gPNHZ=CDSZgX9S
C]P-U33:aPHK-:><G^1LT4UY4/U;SNI:L[F3V.O&4aID22:aY)U?>L(B0MI<Y1>d
g5PM,N5R#C24K&2J_5L]A:#b4aXR\A&^2:NOc\3=000-N)Vf6cS,b;:T.O;MPCOT
I?2\DLG34=>/V(9=AD3K->S,;8f)=RLRSC6_X50<g_--[:CY?2P+,EBB&YY6?<)K
.OIE+CI6LBG@M7F\b.&PZD&e?M;(KION)0[A4S)g2C]IRYXEW)bd^ECY^__LYb9(
g^NXb[f>X?]MAK^:UB0XU):O\>@7-V3Xa5fd56)MXNZ^Ca_&>>[M3f<9^A[RWg1b
M9;2PU/^]5)1+=;#JCT_LaBe[U@\XYI+D3S6ZS+]Z377gGDIH2]=57J(\K4OW]L6
FgFa:Z6?dTXdJ\8#gLRJ:a6?:bCOfY+0eO0^/QIONZ08:4aC.)H:5)R7:bWCefIX
]QD6+N<:c]0-;=VV7+2ECO=3_gG0(a7gU/DQLEM#8.P7#@3e6.]e@2^fT)U?a,eN
OFBa\LUPR,[0Bg47)F/9O69M3_A,:NfGGMR;9YHC<e^+,Q&8A_TC-K^H5Nd;gYEE
\9FSCCDG?g;JOb#]A6\Veg]WE1;HW8]_\a0528H#21T,SK(.=&GCK_7Ca51dII8a
B1N6(;GUU[O@@=MZPHe?EY+TLE.=PYOF0:dJCg&c#XQ]A.S6G;=6XeRbc/RcL=@#
_)V9fc_=5cNI]&c9D@,H,E:WB>2C0D<@G<A:1:b1;OWYg#==M53V0N17XM_<B]bK
cEa.eOH^QL<2>U^-ASW.@_7-L+G5#KHGDY#1+BPMTE0(g-[\(&)O4E.(a4bbOb+)
#,YZ/L5/D,d^.),\eC09=3AWS/2]J\>+5Y=ABBE1JS70QXC[ZX/4[[4_C98OF)RJ
.gbY(R/U?OJY:d5g^>Dd,),&F>B)(?Z+fWV[gGN>9]UOAW.AZ+YW^DHUHR#9_=1S
N4gDed,f==G_[Ng(],-7UHBe]F6feBM<39R6A?gMJ>V;4I>U/?O.)Y;5J0T:O.D,
.-PdA-GdHAc[,<4ZUa1SW0AU.(TPK)_UG(\7Z71@e2>M8#OE(76&<fG[a>(##e(J
K0](DU5A:=b?K4Z;_DTXG@Eb5a@-F]/MIY)GSYC/JRW0DSI;6^T[C]c8/]#Z1a0G
B,2@BL=ZDN#gWU7&K[7cP7-WJNS5_0([c?4V<J^ZWJDI<N^#2aS1cZ<<XHNb7FCf
Cf\bOSHLC5ORdb;QE?J27g1JeE?bR9LBJ+TZ)2-_\I&PfaE397V7^B3=9;7g9E#R
b3]#DJF+6KZVOET#CR-^BZE4bW=-T2K(CT#W&P;J-dD=TFbgJ(cdegQ?LO;B78;J
VMCgBNQf-T.2ZD8K0K-cO7d\E_[^Eed4>0dHTKgOV77_TSg++8;fZUI\JYQV>PHa
VC6S;Rg.I;X=\0eY36T>]]?#W23Hg+\>gME>D(b(S@a[X9YDYW4P+C?gX&KbGAL3
@;Y+UJVS3;]W7WZAI=>?J3Y(:.UTdFP9gMZ,&BXJ[.,0NOfR3+[5?^HI:4P)+c,U
TA<^1KE1HG7A(\e5Y)LGW&4WeEW75VDU@I8ab7\NRf-GTD[#(:L\<+OJ[9)1HI8U
3JUY.\HgYRfH^AZ#bW9f@[Q#ECR8A])7<4X#2f-VR#cCZW#W=f2aME->><M)C^,L
L[/XH#D;->C.5GM0W]LIXCAKI/2=\E28^+.Ef?;3+U#CK/#QWf1V)d_@Z;P>Lc[]
+Nf,LM48B_T(-a>\])+0Vf]MBMXa^8+]F12CgQM2ORO<A.+41=7-CI>Q_S.1(NLF
?F&M\(X;fKV?c]9@\P=aE_ce=<[ZHQ&#&G4B<JHF>5<<6U-#UIH@/MKS<BUU;6?9
c&\?]4fYdEc0-d?L;5EL<6>X/[ZS<SP?1cE;(W8+AY7]12e9[J3+gF<-eC6(LdNP
gS;D\T:,5]b8T5X[<A+5\:A&WJ@A/50.W&Vg+.[_a^/N#,ZT23C.A>AH;37^HZP=
]I#KSPP1E6SUYM\:6+RA+3HM(I-b_:gW&;37.&WQ9ad8Ga97FY\4CTFY-?gV:EZY
OR4aW5Z,^#<<7SSdJ4J+S5Q>Ob698L>XS_D93,D+2G7dL5T2>TN(V/\FBDV(LNKd
YQCc(;PN04ZH:bHeQ(AFN)1c_eQN95<01J-=2K)(A52T<U\HgO(^NFC6R)I>0dS-
U3NKPaf_CI\/S.UU)8>6:e?JU4I]_^O>L(f[[fBb_.(b];Pa_AA11.3G[C\KM@QN
?((+S:8=6OMW(]W<cRbJN0a.#>1QKO+1>Y&);]1^<f^(=Q>K\>&/E)+C<\d1-a)T
g,f?#6cEGZ0,2/WAOW]Y_G7(I/1DB.4;EO@HR:V4.G^QXL]SF9db4\W9)FLXF0L@
#GR/FS1U87A)JcbXUg1Z??[HF;SObaXIIM/?fX-@a_C65JaD02+IIY9>9;gLfF90
&K2\3WGM90ABS=Occ.-]P(/]ATRGF68PY]VKF4Y)0D@M-.[T0.5KfUBOY9=N1)Z\
a@TGO8KUGP;dYQ)HedQfR.b,U>1XARUWB_UNae-:=/L6dZ5-RVRO/Td>>GgTF_2)
a^6N5)P7>H7\QO>M]W=f^L8[X=)XQP.^3Q#cEf\CR3Q[3ca_U/RM@HTf0.YQ&15a
.LIcd6]F?:,\.[R8gEG620)+YKc]F^Y;Jg]6D+IdSbMA.:_gE]SHe7<f<&8d/I\8
d+@gH.]JS5.7WNSB1]]cb<4P9.^<D@?,bW05@8LK^13AW9YDCJBd)5?S8+0YZ)4V
[KRGIS65b12KB+P]b8#Nf/7SN0cS5-WUT7+15e?@(W&e@P>_T)b]/R+T?LM.9@\5
,L8g<W6CWM;P@@9beU/b(aI7:;8USWXLd#e2?bf][gba9GN<T4IYG84#GE:DFN-8
,BCE8>,3C6^(><VE5U:3#3=L:S4495Z&-F.a[O;;O<8XEcF7UMNff(&\Cf5;^RY?
]QdW3R]@]d&D@I[(#fN@]]X.8G/X+628dEL#37GJbZ3Xe.^.^#NVQQ4/_9?B9YAK
0&VU,b.bdd+.^MT0c;FY5?MbMD^#\00_WDRYC7d.BN2B#1-eedS2GF>)M@6Q.dd>
@ZVX4b[C=(eAQEPFM1<T)<#)QG[#@^beHRMe#T>b]]056F]<)MMa?8K)-fON+T4)
<Bd9:QD@@.E:eMG:TO\K3T5)^^]C=H5QJTJaeEdZA]&4EF3DM@BYMG4:K/a2aag?
U(@dOBU.5F?G]#^D0fJNd0+CT#cGeaeS6M+\a@)H4@[97D)ga4;S#A9,,cG;)/?(
f#D_BXS]98&6,9]F..CV0gV_6+/_I6M&K\45.=E&8N_58]O)/:#bAET8K3XSfFP^
BY>LJPHZJ.@)M^RU]TMY3X?SgITW+B(\95b?:1BebNZ5f-c2Ncb;3cObJ<<^XQf_
,H]P?#VVBVJRX@D=KdGR[a^5]8I8PU>\C?X?G\STNG<bH&4[CP6QEb=66::CJ,)J
1/P&cg2gRB0.6H@\D>ISUb\:X\YNTPTIWETU;XE?KNJ15(g^YZ/VO>13_dBd++YR
GM6)L&1eQ^P&7#4W.GUTY,H\\/\SK^\Lb0=Q+HdRB5YUY4W(C_fGe+T,K\(e__:8
-_RLN3D5eg6DeS@ZJYQZW7C[IPL+;f<PUU9UZGX7b3.BX<SH=JeVN?L2O3U:b;=9
56K_4@6.UQB0c94O2=c,U,RT+^LeBRESYF;.d[#H.5D)fIG]a)T-9INND5\:R+X>
=a+(3J0;@d--@OR+X52KS1f)@S6Q,XcEN-#@9U<NS/5S@MSU-XUb:BQbFT(_+;5e
/)fPI6?.PC?[-[4M0C7-8_Y:12:7H>#L=aZc:)+DZRe4ZQX-_6c4cK>@eSYH2>4Z
R_-4G2W-NLLM\61^1JBdB&6_^370I[;G_WT@4a@<7?MQP.D]@62XT1.WccK486G7
@C\MH4M/c>HaY0J-<46T3d@^2aL/B_VD@d.SIF2\Q--[/KYgJ<?(5TTFG)_W;JT[
4>e)QLBbLNC\-5+WM6/bWS(:aC]S8V#HS9dNZ#cAI(JUAS,H+MWG-H><:OQ?eaZ7
W?LYH-[+O=N9+Z)cA7;S.584AfP&X<Sb.]&>eab,fI^):gZU2XGf_#5U@J&AD0=A
6R6cYU=\PVI)]Z5c+OX07GX]bW^W88#RHf?GG?FC-]_bDX,Je,+.0HW2H3\9MD=@
RDeBeF9K?Tc77CMg@1IfaVBKVB=Rg2DVBg;7Pc?[bF>g6?RZTaVa^<b&1E_C;^^C
9-#K-Af:PS6a]NU][KC#+GBLe+L;cX?E4M#L&=McW(Tf7KFX9FJcZ0AG@;.eM6H/
K1bU77c;[?_/G\((.0)F6C1O8L==7)FK9A/3WZBNQPCB:,f0A4He?7_:\>_PS&9H
1bd3W0EQeT#)TS0?=2QL0<?0_b.A\G@d4A+R1A_NGQ+<TH7bP-g4<]4KCI3IJY[:
P6H2b_G23#&FGSA7PKXcPQIa+(d\c+_IXJ#9L8S3ba);NdE.6gYaFG/)?.dIAd<:
K1E-.]/RZc7AKAaZF/9J5\\(.E(:_>+(E6E(H9,4C.B9aHJUG[S.Be67(\QL))I8
&[[D,.I3E.-TJO8@U6MSS5Z^c_?DH;G/e#IHZf0Q=,f5Ud)BIfdW2N9gVH_ZfgA?
T::U8a]H6eBT=DE/Tfc@U(_XNCX&.b[2WC_PD1JJIc7&P(<,L4:7J#\Ib+.[FQ&,
R?.Y)<WaINIZ^T6^Y\XWd./S?N41^I4f)IAC(JdaD]1_?I/VT\J[-.X/UV2cWJN?
;WdJ\.a=/X5<E&0:=7X[XCZ9U[0D.3Q9V[=K+IJ,6:EW(_SY1FG<;:5^@0UA;bB9
XF:T,.WO:?&JeE(5F<X@TIQO^?#9ff#(RWF\-,7U3J#ZI-@gGSJ03SH(Bc)YfP&B
[_E>gL@]0:4I0,K8Q]1J_G:J@FRIJgaPA@c2X2NJ6;7f(_PII8fNUQ<7)fO9b20?
:[V)+W/)?cXZ=H.&QK8N<c@&e9ZIeD_#@3):)D:@^)47WJ2e.YX01Q#adg66a+/Q
[/HZ;@9bH4M:8LN/ULf_UX&.CHPZY+&N:ZCa/X\/(6M@7E04XX..CcS.>6Q^+BG?
DP-OIZ&H,[bIc:I2Y_>=)M5SL2,3(F7OO8&d316N^OBW(W6=)I<+0UfOP?QUG/CK
(NI+Oab+.6OaK#Hd0Pg]J+2d26M)YbA23W[aCE2UgCS.+9+L^:+@DDY=.^/P3Y2P
-KX6cD05(,X193Ae8K7+GbTgIH/)XCYFV(TZ:<Ud4JO://2eaGXW9PZ#:8b&]Y5O
-83BXE2.@#SWW4F4D/HNMOHE24^1S3f?e<W7+V<9A8VOf0.TeDMPd+)QbR<:9gX+
ITO@M3:Z(WR@N^<e.9C1>7LgAW9ABZ+;A0C5D^QB?Z]LR]5Qa.5XR4:^T=P&fSSL
9WM\@THN(HdJ[FW?XT1W[)P(8X6IRHGBG0W\8cG<0XBVFfg:,BS_Pa6#SN/-76F(
^fecg7TU_,9+<[cg)@U=</.TPU#g:7fP=+W.7E:IQ<f(aPM[d]8gdD>fF>+TBd5G
>Y0;>f-7L,AV+eMaA;&QT>f12_(M>cf)[gS64C3#-fcM?\NIafB,^>0@:L#Yf\HJ
WPAIA0,H[#3=fCVP@&(+/KYg+Yc\=gJHS[>8Y3(S[/0I<KTP3^gX(:BSfN5)c@Q[
c7=P<>HaEVW^L-D;X+_MFPV=.Q8T;0fS&AU][VKIHIS7]^X1.RQVN@=T(b(]#2]O
366BRR.>FRJ,TK13P,@>bTGQ5,06J\f-@8L)9Z0T:e4&cF16OcC9=F,W0X/G)(Q(
QDb?8fY,CF\dRAd(\(fQ^N2;B2.S1I4WYgAI/Kf7@6[@OY11SfYeO@:MMSJT?9]B
YEK._15g,_Y>NeY]=23Q7UQ=7?FCDHL5:_::J>SG5MedZIXU:^BbYF/ZZRg6<#R8
Z,;5M)7ed+L6L(1_;@Y:F&]#g,5:TRWT5#9CD6O4dHJ#>N#NH&USSebF:/D884Jc
AGDfG#3A;_[(B:\_fM[gDPGEg,5XA@@fZR5L?^AX]6;GRHac-))IF^2,d@9+--M0
/4)5[ZW&YNV#EMf]W2RW42K6a?TE,P?HF>0GEZ]4ZEbGK>KF:BJ:H)R>F<(a\?VT
3E>GR#H^XQH7V(@NF/2[3?+cY_3]7cf:5G<ESOAe5?LN?<RbdX_ZeN;LPCKB\RaX
--;/UD3+]=(>75I319d^M1gfMS,#=Ca=GFbEPDP#BIMHU<5+GAE@SZJ1NHOHD8NB
A^<c;9.24e=Ge?fT;bGTYb20O_^(MZ4(@WBU):BF0+\A>+4^0Y9Z2O+KY>4La(CN
W_RXU3(?]UV=Wcd<Y:<)_EMZJA5ccK7I,52RLB)_.2[G4N5G;HKG_K1X5:1=gcTb
5,O3YHY.0Gf>[R_;d(NU)D)F43.a;5E55/3J];[Tb7Q>FX2C3\[(A5)HAW=X.D,g
KKA:TZ/e@8d2]6L,NO&^3N0VKGg>[E7L;O>R\W#&/KU#6XgP2&EWAP2E]ABFLFT>
P=);.&bbAAGPOY:0L+ba)/e&6RHbX7T=4I&75X<DOV>R7,;VG81DK3C+<Y[]2c4D
H\^L4fT^>6/2^W]<1UbIMUT)S6X5RC=fd7@e\PD&5N(GG9JSXPP2IFNHX@XOT579
K>C^\YDS0ba\5];ZHY9F?BEUffd#\G]^R:20TR@R<PB:I<?T2OXTbT\5GWDYX=SX
)FUAa0_/5:<3Q]MP,@612J;I3PSUS/\.)4g]b:6b750FPM=X-R\YI;0T_.cI_Qd=
6-Nf?RL3-PRe<]S=?KNYeXJ-5a5E>PYf=IFcW.RC(A3^^8LBXa^452OfbJfRV4Ka
F(HF@&@;]U0=e<OYRDCLb3A7KH9/[6[1MK[@dZX(_;-fRV,dZacF<fY1-Q.GXc+[
bbD_;<;W@LC3ZZSND=Ic[/[/bCAPcMe9NEa49@d-@K,86_]O1@gd<S@-TJ_bF4gA
+Z+^==539DHQ9KOQ5=(0cD:<BU_@F_),IcbOX6F?OZB7d8QX>Keg5X;XG]\8Z4b<
I9E08)&TXHcT4UTAYd<4E2Af&?8/TP[U[#&.39e<3\/B,,ZR)J]LN1X4.[#+,:f[
U+WTLfb9&Z;fV/Q:ZD>7W]eg&;7Y-FTI?2R91]R<(a;-.6:;N#/.3^(IC&S/ZTY>
3KIY;TF:d]5&0Ke6R+D_DV/SNS+/eFQ7Q<O>dKOdJ@71;M(7dO\4a=H-1J6[T8;&
YX6[B^-8V+:):Gf#YY#P2-E#,eNG:@S=GOEP#6^K<ND5B+(.N([TUSe?Zd(Q?&;X
d1FJ@F6D-UB7dNZXQ_7V;X0Z1ab(^UH61_c_K1I_(N]2V4450Q[TUA2fJMD8_&NX
QOBG&J?&g<d;M\gXe@eGc2T((/D.GcBXK,T91:9+9X&-a,e-=&d/^9.,7\b9+3Vc
N:XH+U@RH>9@,@YdW=W3V.UWMPB[-ZQFd^Hg/=@9Kfe)ee@SUB<T/P:,-VO2c(5d
4X0X7cG.I[1R,=X,7[dX/=8Bcf&e:fIB?RaCED:9+\\5?6;W[11f:C58FCMFQM58
Df@ce9A/+#gUE,+[I>IU<R1:2V,>Z1][^JCJ\>U_R)fN8DGb.G3(QB>(TIQ_Y@6_
c>e8\.MNA,fP(a7GKH\B,+L3+1H8+)Le:/7P)_I_aWAP3_&D<6O)34VJ@Z<MQG[=
#]GN2c?N4Q<94=<E@3+,&;LX/G<A?Ig64:bFH^;cgGQQ?9LFCC_K,2af-fE=ZMNP
JWcX71Fb@/N5H/87MQ;L@3fa2HANf6&E>W[6d7Ie;H9&N9(E5NJ&bdbe7M65G/_W
MbD(KED<N.V[II?cg,7E(YJK.\I-BJI<GLC)M\1V1)_f3(M<T&T075?gP9UW+XNS
63O8KCY#Fbd0:G:QVD>ed6]?:0TNb&W\E9^JFKNc]e/FfY5cFXFT6Be9QI\;(\D#
]<M_e^@U+)D(YA5:0(fM)Ja#YS1213Xd]FH40&<;bOOIcM(#TS^4?)J?QYb&K<V/
&C;#IgU3>PV,<ZPA()Z)WC^CQ#8Ffa38Wb[=7)(4AJ)dbK=(APN2;B?U6N\S/GMT
gdFA&;6Lf/Y[TGLDW.Qgg5K@5^GO,FEcR/M9edPRH0g9-.HPS>KR>5U-4Hdg0[9.
fe]4Vcc624NK^XBgEY4_eCDM\O>aQ()+)&J\R-/BF;BAMDWRBLQZ>8B>]Rd5A<ZK
gdQ8VgI1D(Zd0-[c.KF2eE1VEHU>&&;T7Fc]+K:)M8@E(>IcGJYD7DC7@N+:9d2P
]XQPJ6\>BgXeNV9(S\g\2F25_Q\PQ#,?339O^/FYZ-WQ[N3U(YfPJX9I&:0@QXV,
SXSZ7C84Qc[_fWBT7-I)<61g\]LbGI@L4_VJY;/4aGZA.6M_f.2-NFgMTO^^\+?3
fb^ZD?E8<OS]7/)V(c:Z=_ICZ;?e8(CE2^6I129UJ=a_L;H8J_PQJWIdGY?MQcfA
=[C4)1JYTf,KQ8=bTH[eHD&4#LAB=B3\\JA>D)(J_(WO2<+,>=6#59=F0G\<.:a2
]NUFg-[7HO3->DU;=+gDLDRAEa3/OQGGAG3A&B:#^I4)NW<5LOcTJ.0d1Y:M6=C9
Y:-+\;2dN8XMa+-GOT8]+B,K3ZH,<498HZ585ZR)]P1Z4;?9UX/X^)8+^VK#STY0
AX?P\A-W4T,1L(?GZAZb@FPDL608dA1GP^&c?NVL[)/BR1[&5=11@6.A>+17>(<f
TXCec/7+0PPfU#ZJC>.7fJA#A3T[U_-1.eIXYB_=@33)_^BeE>BA1)O2aa>UcD(e
2^\Rg[,XAFBERHYg@[3U<ESHFE2D.@&G+303P/4VYT72W9Wf7SXUG#H]:O(5./H0
Y&H=a#T/_6BG3EfC1A.fa11A3K-AZ_]A93Hb5L72LBCY(dMHT]^Z;J^#[cQdAVAB
dHg.L4X/R/W^Z0AgS>W7#ZTc&)W2@?TU,W,FE4QZF#dQ,-^.:Z+aYfGE8_4?&N.U
1Q5-IPOGYV]5P(aD1/I0O<;d&:<7&^DGbFE:,S#-(RP^7XDcGFB&>gIS_YW]b=?,
2+9^4WEe?)SRYb]>bG7PCZ&\_F<dNS.?Md?N<[TcS&1J>ZKGe-B3[FWf(U>ZQKI1
M2&&gNb,1=[-X]7EW4OO6.fZf+E0bW_(5,0W8BX&b3TYa_fKGSe17>(XK<X#EEO6
T<KA=CcS?KV\JTCBga02dJ42RFUVJ:#LGXOPf[b_\)6K[PDGT_].:;eb-e3?W7#^
UM#eQ8;4STYRbN-,THG._^g:50?U=J\g@g8Yb@2MXK3a^5dE3e+#I-]RX>J:(b+B
RLNI].DBfR>XS23g8<;Uf2F4F]L43UMYU+[IbXV)9;=\9/2RO50\16F^J^\84&f3
,-M(20DS&3d?V85INSXD)Y^BU5eGU39+INHW7\^58@#H0Og+\EV+4<(@V_Z5VaQ1
b^ET7,(<fH?)C)I;?/)eO9Q.?QCcN1JIGSM33A\#K\:?H+.bfOYMEQFb@a=Z8J+&
SJ4#8H\-^?KSH1Z6,J.GV30T80f7F]_bMG.K<Y>K9QB#5TJXMA9;A.XI?:5Fg7Ue
Q=(dV#f/+]&FbPD4fe8>2X])\1/29a:1)8P]RadRAGNQ+PM<a2]UC>VQOU8&b5U2
[/+3)-1U/XKAHO=060&cP^6dNgB7-X<ZDg3-]1H5/V@:WHbB=2J7,]S\/LTT[VKY
BZ)EB=;_5W,2(;;d&G;AZD(?NCM,_EU0<9?O@JbMSM)eQfXfC7dIK^WZ=gT\ZJ.Q
[,;GEeeT\4>Dd+))I^Cf;K7L;DG&TWf-XSZIC(+YPK_LY_(5=]G4/d[P4ZbFN:Z6
&1P:WKUaRAI/QO=H#^eGbC98WWNfa96CB=#YCOI/.6Z6XH.aZ^Eb<O_REYE<RdV^
KS,\E>C8MF)88>R<(<B7DYMJ3CF6N25eI=^HG_14R[X#Lf)W,/9:e@Q:aJae1WXK
[I)SEKg)JKBb;L8,SaGG;PRdH1S_95D/-;^R/R/[d4VD+L-[Z&P>,A;<da-AeQ+b
:Jg^D4.1PNd1c]._<:L1:3+>(e>g@KAZg-)@Y\MOae,\XH@NU5@O?BZCY(9>D\B<
(A--,W[()EeW?bOb0,fHc=&.FPYC;3DdfJ6\,UI+8;(?=87GEYPT1BWg9_\U2Y1N
SOL0f+#1_U5E>TJO\AL;a6T(_H^[e\dSZ=[BA_fL/N8:ZCZ5;FG.&?>Wa44:Ndea
X#c-Wg18T19S3)\/OeI]V?5[:FNUCJA_,PF\@JLGIRQe4(REPB7fH(SJ+IZA>UY:
4^6/e/+90T/&Q]4:_W<cP@@@[)>TA47?^2)cF^)5P<\[26=;<5C7][16BNd=X^[8
W]OK<KH;NeYfQR=f/IY19-[PNJSHR.(C?N@HOfXC_61+(gaE(PB\99T(>0J+_gR+
/\P[(+_BM/&ZD5eT)+>S8&9Xc/V8#9E5LB=Rae^?d71c(YDL2V8L-[,eG2/Vf_a9
0fd;aN+T)=,RL_I\90G/J8>U[_e\Y2KGc;bU+4930R)f)O5ce-bKe)fT[/Xg]4\0
1S\\20L4I4E<>[:/c5=..eP&_>D/D;NI;=MDN/R&O-34-FaLe1ZfM.6.F(e8L84E
<L+TD@KKTgReE87U3ZDAI]_:H]8OW6-:,Ke3H2?CG\1JGAgaHU/VR<2(@?df<;,Z
BHH<6\B/gc(bE9_>XZ+6#[XG<M<WYD&+bY@&V2#0<JLI-Z?C@T#S[YUKWDGaM23,
W\Ge;16,F5Y#)-HEO<)]T&PU.,7Sd8S=OU#A<VC>&4^F/43C?7&?-b+-2/gWBX.S
8\8Q,\>,FPeYGYR(X>7#QBC>aM]?QYM[^0AIYRY;)]]Z4CRRZ[^]e=D5)#3e92+6
EPP;-,7Y9f;C(#+(:A-M,)@^+e6WSR^S+]b#:J]5G&a#PO>)V@@6N+P1^(TD?DeH
MN<BWLJGU<^PA)3#[(L7<KG4#5g9XQJVU?)3gA.Q#.6cU>eRR)gDa:fMF]_Vg@,W
C60?^[d//RHE>-)[NHYc:DTF_##X^S]AI\<,;gI@IIR^#/6>K0D.,Q@O0DQ&\&fT
Q1+PfEDZNc]7Z4JbK>\AG_5H379&9>Zc6<=(I@9PL/;R^BE)]@7d=f0TZS7-@]3H
(18,4AMAXS[C:ZdXd/MUI(#0UTCOJ5_&D1.fB^ZZGYH+P[B:5f+/A0&Kf@NQ1C:f
bg;=PZQ]25K>L4b67V:G1eOd^MP1aL2EE?95X1^3S5d7cf<0eVUE.>I7MU,4,Z=)
27P?@Y<)efU+,b>,GJ^++)d&8/3#A#^A?#D(88f?((T.BK,OY-FWN#-M#QbI1>O\
=6gZ@1O+cb&c-Y6,/VMcO&82b^f]S;d-fX3P6_G@GOR<4<3WMd\RJKMG,;J91B5C
UAA&+SLdc9.X.ABWIJ@d^LO3&O<.PUVYOVW:<eJF&#:](39&);T(.#^?H4W0]:G@
OeYL;9;44#4+/3S](]A0<?[7_\QKGY_S;/g63C;SU6Le>YH^Z1\1W=^Q-^bNY+-[
E&M<,g\O\[b7V3/_7e]YZ^A9W,0EM+]8FB.4P&E_7YU@=RcLC8=6.9MK;8##8.@N
M@BWOI/_gMYgVG_#H41<1gU/g8K^,aUbB^YDWJE,TU_NW&3A\C6=XGb\;;/bNP+R
#03[cU9(439G4M[;0#=+ca97SaFA>\L<E2b9,HU9?.?3DS6/J@239(B5)06/=[cC
/0ZU4KJDC]U#;4PPF,T&_3;5=RDCH63RN66OIV7cL(Yf51b@LW@)&IRM\>WG]>R)
^[Ja,4MRd@DIMWdc69aa8P8AEK#f1=Z8)bQ8+#YFF_I3RF0?9+d1(Y1TBcNMUD=f
8YW(92U1@06#W62()8+KYV./,(YSC18-SAU6=0FRFP8d,0K4M_WKP845GYg\\fHd
VPe6P2_;5_MK>:#I4+3PSXWN&#YA1=_ODS>HB?MF]^5JLRI&H:GbFf@Ub\^P5?;.
_WY/Y+T_N+RSAHL,APdWgX<O7,-67EMSVBLL@a]bBB6WUV6X\^^@_8<YVP)O_bbE
E1^g\QF.A7Z<H>ID[;A?J[T==1\=PH5I=A/@OLA/-Rc9HUDbAf?ZRbF,dW)N?.SO
CN.5WeW9eP)-_JgUIT3TWX=&;&./XF,fcS8)ALD>5F<YVRH9H8.M]_K)HgTDZR,<
bP:;dP7TF;^EXQ1R)V)Zd7feE>EP0PX#N8&J(/MdN?X,_D8SB4OcU,ZGP9[;Fe5.
]/QDP=c+W>::;+V>gefe9JcKG6.]aO4]9La\Ga2S]@_Ga#<faAAT.C9=M4?L1>P[
dTO<;L-8JX&\^EPN-,E;+&bPC+P8_gPG0^5Y=W4fZ+07AAD1f(H>ZXEV9ZS0MUYc
0GNE_(bd<4MU3aO_YB^LFI/:TKS@4-,[P;fFcLP?149;MRaRSNDV^/?N]#?>Te1I
GG^#MAK[Z]UbOD/d?Gf35,a9d)-W:.P[8g[g@4,3+e&&TYR]bJCE67L^A\K2DLcA
/.LfY;:UPgN98R4X8TVZ?(6T0A=-US79GJ>0I(YZFM,a[Q^[Nc+5e95#E2LY(TF2
YNGd-F?aD^+K0eC\^bT90=KF+3gbRM[[63F2HZV^+\QD,-e?]<&ZcbD0-6QHgC7Z
(7&MD<TO)+\P:-3PI_c/PeOVLaOO)gS(H7;T<N^3;23-B/@;)=(:X&:2#\@(5J\]
LUa+6<F6K;C9F7DO5Mb@S1>)Q,]R:;:M7S_(N?^3YfKASBa6#X4>JYTe0^;-;<L^
>bcb)4f^cC,SF\-&Z9M,2?&E9^4G#//AaVf9_De.DB-W7aZ=E&(A:L5#\]KT,+&N
]c=AI+UAE,II3UXPd#aQ&-CTe?GIC-d5O=I++YGcJcX^,[P=)4KIgbfT:G7^N-Ab
d#26Tg5TQ21).H>N?fR^^PS&&I/W)Z;#PI^A?DEX@X5@,A3G1eV@N+CKE@U1AR[I
6C(:@#&LS;ZF</83]S<<5JGC8JK6,0]3E@6#?:(-@((c;g\-(O-DG2,dg3_H;C+B
^QHb(g5OXeZJ;aMG&UH02Y][UJ[I#?F]/5g3D+B#dSQe^+YN\-U(LYMJbCARMbf:
&VYe)P/f=6VQXc.-C+7<fGACc\Q])-TbWTgK[@=;eR8G+VYBT.c;PW>E,+,<]MXA
2;XSD3@[WCZUL3@DfP88dPa8FE?=M1><HeP43ADE:H=Z[]G:A2XZc;dg)?G.722+
aOG\\F1aQD_1KLL\(G:&;cRf7cK<8X@]B&g0^B)[&GeS9(bOT(>]I9NXcVC>a)<R
:.CI[C&(I=&5,+J]5A9>_,IGUDK(L24gf/Eee&4a.[gA2-A&bG9EM:=N8aV,@Z8(
)4:R-LWL]Q<^gZZDB>XG.)#G+J3QX&^N7=J>,<UTH.K+^,S=c6R_J-2)#cREG+BH
^#eZ0Qa<>T(HT6WcNW0G\bg.,+C@U]/fOA=JdgS5VR:I=ECH.J=bfIf]0Q2GQEgB
1Pa,(/RDDF.SXI(QQ7@681Fd2f,FFXgcCAW:W+\WMR(Ib>48If\QB]SI2:+Zf/3#
A<RFD9-,O>Of1Fd]REHX\PgXH<_dMC?8V.+1:,DFUI[K:KgZ(UQY3JP1.(dWDI;E
M_.\e&WaE1@@/]5Q\@F,Ne>+DWQ&0E:MH7VG@:=BKY;7E4W65ObQB?W6aLWYH(\V
4J^?L<KLZ;@;H1FT/]BNHe@H4UW/P7I2GP9YKea5AW8]b[;_UKN58J3XL.5dXGF@
F)MPR:a6,OD\0dUMTT>g4T0U@YE])E4T2eTU2P>T)CVZ@ZV=ReJTJ8#9QD__Nb8P
H1?L[d<@B<7+:bF,gCg?-:/c,+9aWEYU.^V8FgSD.T1,;+P8XAN3M5]\MO\W.TV2
A;E@X7[b,&;U(P#I3C5EE)-:D:@XWab?5T?KaeQS?+/XZY4CEV:LW[gI[/YHP.bH
A&9-^]Y0ZD<1_V/f5:12RAKBQ,DD))(Q@,P+8/J8We#:0:2g:WK51.]1&6WL7\G=
Y4)4@=-30WK.K4SSPD5EPc8Z?NU5ff-.87G>N(I+T)^,BXQ2\dH01H=X_Z.S.>G=
)CS#9cZ/4/egX5@YL#5aVe?A@/3&#OX5d#0H+D>8N8e]RF6V8[R+Nf)f9[Lbf^MM
0[+&F@M,Ra6/PQX[<_P^D0Q:L1G^+LeT\R12:7[4Z>V4f?6Y8B3#AK-/P):F76cS
5X3Y0^FISQP,ZWP>+E#(LO\(,.-,1=)NWYH_Y<06=AagcOH[CV?3@&<W]=Q#[ED<
gPe??O;962O4#RT,Y<AHDNEUV5:3b8)/=8Ea_PY<P.BbA2+5?Ld@bH/\.SR&LAQ]
,195]GDePDSd-)([1-<[?Y\P4SXT6>W0+eN]K]a@acfGI(VMENee+BfP?=B;BJ+L
#</KGgB]CJ[G&#FF4990H/68L#?cRbFF>CJ3S2]5J.^R3,;0H=:>YCV(=O2bIf/I
Ac_?P.5X:8B+;,_^&LTY?X^FTT7AX5G96aEEd5M,1-dWP^\d]WA@F7&b10?5?294
?&V@0@4-]\eB^M=W)Yb4BQ]OeT(b>d7[^V6Q&(^)PX4L^7E:4>6,?K0M_c#FWGP8
BRgDNCZR2Za(TeP\P;HMC&gOBHdQA0CM38KAJF,8;bYU8VPL)RaafDAZ.Ug(TMY7
G&1)GZ7#=-+WMeb9QP05&gP^PTN<-d_-b?;KDF__RR-H;FW32BN8ORVd6g)Ob3gM
L]Ya:;M2b8+/]NC\GDT94:Ue;-9AT;A>Z[D/SaKKSXULE0;;EK]NB6^?FA(BQ5W_
-S.?G\BG_9g.^DNWEWRgR]6^S8WZ5NB4MA4aZ\U0,[KX+gHC^2P[[?ENK]c+bHZI
=/\5J-<YKfdKSI@);:aKNVKJO[N;2LKAYU2QJ3eGNWK1adU\dd)WXBSDZH5KMV4?
g;-7[;:@HY#>/JG^NWKRH;]X0,TD&N^cX&K@F:MJd&@/d;38Vc+]RUSeGW?7>0A.
)[Zg2fHQVB,?f5<]Y)?C/G#(K7HZCAGfIc,Tf&,V(<EF<RU_7,0YHK&,5@UcDD3Y
7@b6-Yb286<:5O>dNVH.[?G)Z/1:WK^KDS?MV3(UcBa>A2##.AYg?3[=(.X)+GIe
:]W]/=bagRNMD;-c-\)S]5GY4)PZ/B-N-V-b).RM_3\R\;L4M8ERI0Vb.T3#Y94a
8UY3T#EL<FJ70F/?A)U\3]/dC)OO.ZdcK#PWZJe4.EcH0BSD3#R.LL[W#dWIN>+N
J<64+cAUbgCOBV3(ef8\QV7aI>@H#?9E_,W)CTM5PS_J2@BXR^74B;>ge=Q>YT[G
?C0X]@PT(DE_2aMP[/RG60N?4L)DDf_SSAJZH,8Ke7d?/5FNA-D^ALJ)VWI@a-+V
WbQ>)Pd9&J)bd83>cWV3IQ40@EZ(?]/^[AKR\UR..I62XNO#ESQ4Vg9=#3XUD>5X
?:]g]g@;?JXX7^cGA]Z9OI8_AQX9eEeJ5UgY2R5-5>T8R[33LX(:KK\-Kb-BK2c_
>R,O6e^]c#0UO][a<SKcMKJ6S/Dg\bHGbSO;E4W09]9[Lfe+WZ=cDEbLI+5OMSQO
=I^FNS))Y+#Q]JDdg^\D(eH@gTNC(H>K#B>9)WS>@K#LJZdF=QZO;DLMS94BRSFU
8Q3TEYg\C7R[=U\7\_/S^(AcC0(1?VbDDAd9<@;:HaO;]7eP]b)dE&FIP,,U(8g2
;08c-NS6J1VD3NQ2I5W,/[b?/0I=_-a,\#Z)bVG8:[<E9.F2]R1#3fAYR6]DW#OJ
.>OGW6gOGD@U9-8QUD8E<B9;.NN3aQ:R]/53T:L^aA^Af\[)D7XA1IIZ?6JWCAC3
<+T[TaQEGP?A=W=Ab7.a=,MC]NZU3Jc2aU;@fPFS<+GK<4]^<HCZ);bg2;5C.ZL+
\H0NO-8J_@44^WFQ57,GP\[(_#B]dc6,2(9F#DcYHL]0P0XXC-dT3PdQ,M(O)IML
Qd0BPbS[/8c/(@_7;H<Aa8^>6ZXPF[<(/&Hc6#?.I@bb3>JN#?C8+4T04bJM?>GT
Y(0O(dPN,(DZL5LC9e.;G@8>b[4KV#+c&IBQ_R18V/8ZJ+Gc:UP0eH)GB\d81?)@
dOcSXUaDHKFYKJS,,cWC\(a4NM,/+9d5E=?6c\bLe.bAZHA(\ST+00QN@F&S6<7/
9/9MFaa1F+QPdH9IVOCfQ=OQ67Y)KJWNQQKc@GK\g1LGU_HT99@;Z=8726?(\f=.
fTW6P-,#MT][/Y[[V?1O(_YE,DM4;H])T9F\STXZO\VF+UJgg+4ZN9I1S#,YbP\2
K,b9^&(P0g5ZSEU<[T2VPgS->C5c;5[.4JN8KA#bBST&IWM&6MZd6>.4>]7AgL0J
&J3=REEfaOI/&gS81?^6f&b-=La6gGJ9g+WN+J[.K(K^G8J._1A?6)aN[TKFD6a1
4;[Neb#^:RcY[X&1HcIF+ZM2?3;.<0b1#EM\d((SQF0Y+;[X/M7TDUc+J/GL07W2
[cIZUFEd-#I(,10&F6c;UE<NAJ]Q1(8D1M9+_R,SKa\b3]=:cR0R)Ab3\<1eI&Wf
Z5Z9_fUC(YGGF8Q1)RTALQSD);6KV\<;R>_ea_;3^\;TR\RPIcXLB<L?E[d[7CbU
=G&Pgbe<N;3F_;-S]CY&_?/,E&UaO@=MVg,4@<-eQ@c-\W8_>E:M:?\:&(37gTCg
FKIC>O1H4U4_>#Ff24F9d\=RODSMWR)V><<c4^\JB>YQ3a?0W<6&>]L7/H&(/LF&
ES]e,I42\7eE+M@dW)I/7XPT3,B1P2DXJg+,,;S0^e_^N]Mcg=X(N(7eAd,HR6XJ
/dEB)[N#]N-V;>Q2@PDc7NBS+Vf0f<AS,.OZ+c60LXP<IAVV_17/-V2eB#CF)]<A
D#BK2Y5[6X6X-aAPgc4M]7L+^@3P.EHNd^#26/_dF/E\4@R.RbV8^+/eP>I)J[8C
J4PC\?HM=;81(W?bO54^@Q>??(-,<;D-I>>55#_#X48#LdT5)4\ZHd_?BBc_+Z@a
WQ\[g2J4eM:A]5XZceLC2N<.A-WE\]AOXZ98YJZ]UdAM//fO>P/VL+Q13CNd,a46
OEBH3EfDTAc+abV6Y.aI.6c]3CK/^;X(^ZX1C#(R?g.4VX&+409SC5\+/I7-4<3f
f[A.K9S)T:BcBV[b?1+=BKL4W@78_.VTMIf6U20dM\UA9,=M.3&E\OL13g4\dB1<
+aaI69AG5WQZY@^D+#./Lae2BbB2I_XcZC^7>+9aX_VFF2C,UH[-A-2PTTfSWf)b
>8Tf;Sb9\T(a2^J5+,7SX&L7UU_@7(\./T:T9]VZ/e5aF#7UBe/;ETeb+F<LaPec
6\.bVGMI4T92\?&SWR.-@/@P7_L:bUJE^,LPQ)V1/Ib<0=2,fdVf/(?6@07N;7H)
?L\,Z3#5;Y3?#,V=gZH:Q<QCabT1[BND?+>][<7ME:9.X1<R8)QQV(\]3W7B4[TM
T5<JQT)H_>0H/T;M^MAFEOD/8CaKD_MZ=H14]&_e><&#/\9DI,8K<bR\;S4Zc6=H
?8);^TbN]CR_7Zcge.D9L4DLX2ZgW0@DRCNTJAQ\[e00-bFH]HYO?f6^K7+[H[8<
HY78RP28Fb9F>LPI=OH=#3ESbVYF=a>bb;SHeU1PY&f1ID71:LPJIVNI:,VFNZX]
BD4PKD:#3_4Wd9fg;J;5&PCWd;X9+Lc7c[Y)Mc-5JDCT:2VWX/PX5b0A7?^+[JQ,
EP,[PO&KF<LHOJ)X]0UJYA>)YQc8#:NH)W.M[UC<3C7a8Xed3;=1Y)-AL_aTgW6?
GbW#@193T3)<c3b+[YFJ\PO)J(6NJ[fT)T[dO#;H<(cCA^HP?)JVNMX9Y=b4WDO:
O7D;Z+IF(P-.7X0OAB_(+FS8XT(,gg3ZV3D6NfO]3@U;1OAMb;7eBO9#P2Z>fGR^
#<RW^)+-KU\^2I5?;JcUV=[#0C19C2&gVK3KX1^_-\X-P_05SM067^?A27(Q&a>9
0USH/5<S[0^+SE;4LJ;VJ?eeXQZHL_8gb4<<^M1T#[9S3b(&a\WLO-B@&XK1I:76
XX@gD1D@=GeA(W-X12[a=)9076^PgL5LdB1C@6]=KQ-ID-6K1GOaOI6J8I:I<-8U
Mec;X<R_ee(8\0&[S0:;L;^L^.c84DW8T_I[R[bWYPS_S13H&cEb6e,B^Be(4X2D
MZ<@U[JZFQ@]<LVKcFPAB>W<G8C]#(bGf)B4#1K\^(R-LbIT9?ZC1/D09I/4J=d0
?T1+\L(I0WU8_:bBQ\MICNT4d1^X)aYEEa@Y,IDZ;)52/^=TA@P:G<1;MVe:FN]9
E\)6cCa^PRH3Nc3c\+\(.VLgKFF[bC(gV<82A2O1F-P9V=_PJ(<Gf#MY;eUL&>I@
5;FG[g#RCfY[:=TBK#<3;E(LC;WGC:9.+)/H3SL_XY2a;L5e/c0#J?V]#D.gOaWf
9/3)EF(c[3L)NL@1Y#=<Q9;_K)ZR4<M<^dUUagI?b0((JD)JVOeP\JN@K@B=QNRP
MR3D?8MCDY;E?c\c(TIbf?T(d_)#LM+</##(c9-2YKK:E9DS9YZIN[<dAJ6:(g)X
e@:H+eNEg(+KG^W+#I-.J?CWQ]MBFNY;\Z&E9#EQGS\:Q2IOD#>PbADG-ZXBIg-\
2P</e[Mg#_X1RXK[&VZS=OMZFLgV/.EY3KO>1(P&-]JfabMc71@]W&?Y0[6W;G-6
_5LK?(HEOc,d1S>7-T(<8N5U<<NaE+PTGJS>40Mg/+YII6<[2+RNUOOQe3&HG>X5
MNT_S,?Q;Eb@gYga\b;U[7Hd>PW@7UfgZ]2-MZ\S473^KNg24+0?2)T=dH33b@;;
VO29+E,NQ\JL7_^#OX#>N^/;H1Z8V?C]MJGg]Z5F7GP:aCcf>#c\ULCBFN1\Yb>#
_AX[QZ4425@cIKS?,>ZRTKXSTTEBZ[J><VHV3^^EfG9UDME+7./)I3aDT<&GA_ZU
-KHUA_P=FG1<K=WTfI_Zg/;BUPJ4M1_gHU<d(Ya7Pc+WCN2X0MeNE5#O6&:WZbLA
IUKD7P^E)X<VIaLQ<C#8D6)Z/b.9^Og@CDgS<c^R2(dY<HAQ4F#:[bZR418=RVJ2
QRVC?368C5M=YG#b2V,:PEQ?L]@#AYIPB9Y:7O:#b#eNe2ZS/+E_b[R&cAJcD+YJ
eGTMB2)C&M\2DDg51F8g&=CU@WfTZ8ZR-;)-M2Q#;&<3a/4TaR;[<,@G/&T9LN#H
fG)SV8=\AP9G0&&ScQGL6RO,eDCb+N^&)&G.CC=SANbf;2LRX09EC.D.12O(?E.)
[BHOE-cd;89^A>K3B87ZfRf.A/ffe>&?FLT)G#7O6E41a#=_V8FGFCV)</Vb0[XC
EG\Q3=a1N66H<^2=]b6@Z1R-36X)T6-eS(2\3\V0ef2@M(7S[&0(-4)gY_5-_P/B
N)00&]efO=]cdIPSMG]W1BV,GD>aC8JBZd-_\.NVQVTg#gSKK.N]b#beC^A>GF]U
X+LMHcP:^@UL=ZQWN.GIB9Z&fX@RG),W#J)TSZZYdZ(^#]VD8DMD;OZJ^++@T9?/
;dd2:\/\M3)]EEN0bdeJRJB;(2TNH:>Lc;MI).2@2>b\c5:.Y,[Q#71UeFRKe(Jg
#0>e(LMFa,QO+9I97.DU2HeHR10CUX=]BA[)R6Jf985WENfAc)GOJLfDYURSXHPJ
Y.^2(\dCe[O4(#e>?HQ2>B?>RLD[:IFR/KXMF1aA9<a-b2c4A0?bXA\D:C4Y.4[\
K4O?X)DSU0c&43TO@?1F@Y16NUCMB:T/O6fO(AGJ+P_1Z0?317<P->bSU5ARcK/-
+ICCXg#g6.0=5-MQIEIIWVRSA;Y/gZe6AJT(aaL.,4?\H^#G?bT)dd7&c4U_09AD
]@NJGK&>6L1;I1>C6==,IA<2XJQ1:MLbL&47I5+Q-3_)\gbU+D#gaf2O+S47FU[W
B_N(CJ@SP8,-Lagg.0=&gLP)=D#bbf@,b9bL/7V^NN,@Wd^<fb]-CD&X3fYYD:#9
.]Z-F?8?Q_&F<W_aLDG57TIAJ6Y_IG.A4HU,U<:\<g&VDDEEf2QKdT0#6WX0K#??
XJH=cDfH-F77fbVYcE]2VE\>&ADJ3S6VCa,N?g<K5HB.75KD7a)VA1GXOg\M&_2f
CT<LfMgT1;[_e0\J/;R@B9L=YcMV:5Z(,I,3A8>#F9#,_MH3)?XCfR8B<7=7A#)(
R-(A<e^4L(+bL?e+0=IC_,/S;RK=+a\N+f^gd>>NQ_c]Z-E)&__Q7Eg0\Ag0f5G/
7MNH=-H@@Y/L_PT[T/adL>,ac85NZ+Ec/[HBV&;<>HAM<@U3(U;J?8H,Ub@XM?K1
VJG[<:MN,Ie-b6F/.Z)fdE;6??Gb=GZ\2O2C7[B;/If8-\[?D7U3S5PIFHGd1E?N
4bMbIN.,I@EWH..E2A?5>gG1+1Y?)_\.c0U<ET\S.5UR)JWg()I65I7CCd3aEPH4
\#MJXbAKSSE7Ef-Z1AVP4OVW^/2ND?c_/bIGf4(08E^F\1\>2SMLTRI](TFO>_1O
P&d^X<.)?Vg:cdY\1adW^:e[).^^?+THL2dSG\#>,e:HLSK8,?98=LJ8W6+#Ue82
baK/MXa61(8f:#O/&)]&X#-\6[e&^Hf@MLP-YDb^@]M>Y^2>8<\Z_P1?E3(1Y>I;
DM+N4=_(#5Cd,2e#T2L]M\&eXA/F#_5Of9LQ\6FTdU2G+-DK,VZ8]Q[T:Q9&La8]
B4XeT/J8;eeQa5Z\1K8U7.W93G=_SOIS2\,PCbFbG1YE2]YS,agJMG=_c6J_QbW>
:X0f#EKbEM+(Rg>=F@P4&-DS(AI(6S4V&Ng9\_ULd[/F&=GL@cV-.\H[f](BM&^D
?QI0,P&;fFO)YY5C].(U<[VS_WX<+TdTR6F4J7O[:;E<)O+XeCTQC#AJ>X=\G1+]
Z17G6[P\[b7S+cFg6+/D;;UMPMJL@B^g+(9BB<8P/Wg.+X9K8G:_SR@Pd5:XKEY9
X]4:?N[09f0+c6IYMgVI8Ja6TRY_;K,T)>AFDBc/<UcYDWJ\1P@EDK=B+SO<1BO-
af62O@&Dg2Z1_]>aRB8RLZ3#QU]AV(C1A^^cSTY70T^_X4Y664=L<3[&38D+,,U3
K,RVdI#[b;X[ZFb6VYYWbYI]SU0/Q\L.9gOU;bPW.BFQI:SSU(SSON,e#-f36JZ-
fHa\N:L-IV:c7.0HbTKS:AeLd+5-1HRH=_R9X@O/L^M]>QIS9,/PWZPW+P^HK28)
>YT+dBZBXJ31_ZT1DC@4Vda>4ZY.OAd\gG?75?0gVQCaPHRcd@4Cb/S4K,UP#<NC
2dB:AM.OYE[RTQ]@^QH0&(0Dbf:DOFVeE=L@3JT=EV;WXJ@Zb:#1O/]MaX[XR@K4
a;]>Q_A_GI&BT80GX\b[K,NB(a2G5;>29NEM>2).1?]0VGQZbI:.eeS:KD2H9SF7
[]4]S/8fDJA0S;Kd#M>NSgM7QVQ2Q?1:c-K0UYXRX9XB4G7a)&7-JG9#+QTO+aH?
A(?:V7V:D9U.cR9I:IA1@EZUc6:IU_/;,fRSF8aK2:HY)MU1Lg,cQ>#b_+1Y0:b[
-<R0<NZD&F[Lf+#0A-[H_:G#@RN404CJCI+]E-H]CQ<0(.AWJa3YSXV7TcG<F7V2
gJ@/^6JdV.-K]cb)6cPQ22TQU&Gd1CD.0Ud,g_R?F]Ub0(LF>.<AFTe/DP#,[LU\
W0SV5eb;,?fUE^:N1[>H0[R(NZL^4:2D<7(SV/W8:aW_=FLL8.ZH95@+,gQ?KSR.
:Q9F6LYKHPPb13Da4=VYPB1a+(3[HX[NSQC5P1:SI]1_g8gFa32\6EVE0@YW[2G?
Y6WM)OZ4A2K.0J?^.RH#17P&JFYS@Bg:P1J?&#HPg+^+GgQHMR.>b-J&7Ed:Sb,Q
^IIOI_O[?_.MAE3/4.LD9>1H4,fR]F>0>YF_I\XBUJD=X25EHB4?#,E/UKZ3a+/P
0)>FCG47Z\+d/#KIQ\BH&8fAM#SDIM.7QcC7AJ&N/f^9;.Y2B2/R)Z>U+<2M/=QK
OP9_]/?&e39Fc>\[X,f(E#1)Me#V(?a/Q[W?fO^>.bN>I:LX-MQgF\H9T@]-IY5f
,<)FGC&,O?&RQBRCWa\GO5AC1e,b)NIcCNQ1H7UZZ>gJC(^>364[;/BI07?;N@5.
PWTR3.9@\]>N6J(E=QPY]>(<)GL0[VUDO\@TaF&gWTA?&eK73eaQZEcYL[4K[&LD
=,<O(Za?eK,_C;&5),+eYLDZRG_FI#&UGD9c4Gcd-CL]+AE-UI)#0WJg5S:cI72:
7L+ffW\,;;I@ZFWAe3S4XN)5T#=:&CX85DG;X/[752EJ:,RD=2SN&(NdDb\WQMDX
2dCB/5462f@T^97d&:?C9(^O4D;;7>6P5Z]8[4TS:S1S)Q0YXA3>aQbN+e0bDX>7
[Q+AM?QcK^K\OAb5Md&&P;.;B_[c6](XS#bA^E5Y8\\OXX1&^g5L<8=/?AQE&+LL
/=K?Y7-ECWG_X6L^320XMX<A&+^)#eHaTZ&A3gcNMJC&ZZeU3a0]4fdAQK[eED95
J>;@SOA]OQ<Z2.<[<P)6AH;Jb8^O,9g?&JP_A^NZc4M;0#>8ULSC:Q+2OTWR7U>b
6(P0)6.&;gFDV-;a/a30HW^X@dc>.;.L8D?_M-ddZCGO>J7)H9>,1VEUT<6-E[Q/
M/-f\4=@fPA7-\HW[#a6bDOe&X?04QQB].GAc,>5/[U1[OZ01gARE2T=D&WF)9Y-
S]#ES_H>3YD6U(a-f#O[a\a;gY(0R2/8g3DS;R@=(;0BD;9FVX4&+BCB=f4:H0\g
-S+BDB)#.)1-5f4;58_(ZV:f\.V@66[dP\.N_1S2=:QN:Z@1<8g30W,O1A;DT.Be
XVL<I@^eg)W?0N_?5UCI]+C>V261[O\f/?B/C3^9c[BO(V[c&d32ULZG/TL?2&OX
?a6>:[<c5agOSRKDEZ1^GM@?Q0Ve-C-C:.fXA074+I(_bC>a(06>_DJUAcJY.^8M
4&dRH+++PQ^G6?1G>63?EgbI^2b[@_(U2?&1H5T.KH:GVD&</83X/X/)g1PNCMe<
3Q4.JZ&CcR@8D0PeQC/&OP6a8>A\Q9)6YH5>Q9RfBGe^U?\XYS+>YW2N-<W[-.d&
83<J7cI0I07FTN^]<9eP&JX?C<N6+[>9(+@RA;/N?AM)(7Sb#::(e1_TM/PEROQT
P[19_/cc7,W^W4JA6[5+cW0FT)H,IICc,dIgB&;dB@U5a[-U,8gV<O]CCRH9U+U-
2D5X-20cCMXYLe4e&Xd<cRc:T88KGWDYMX8?SYYE1V60[@V2VGe;K:TU9P5J6Fc\
G[cL]Rb>L@@4ID-R13V?UgfIU(FQ]P:>WP/4);bA2(VHY6TfTbb4G:3Y>->5ZDfA
d7M&8>7eGW<7)UVA]/.gJ]G<#GLQc[7[(aVZ:J&;1eK9-HR<K0@bR8UO+6c.;/U_
3I\f9f,]U?U&5K2],d)^T\OCPOf.4)2.AR)GY#gZT[<&Ob3Sa\dN0_C8-6/9]>8_
E]7.)=RcR;8YRG327J0c0KYe]LTE85cB^WSPQO7g(5Gg8.8#_C\US2NX?FAOKe<M
5>[K<^1,XZ:>b;K+d71Ng.aL+eQ9>fCIfNC2LVPSC,GW]Zbe(,G&F&>\<_F1DB)b
WO44b&;SXLN(6[2.EGUWWeJV>e2(-;6)C[#7<fAD\@J^ST.@TLS65I4=?,>9C1d;
)^B#/5TQOQ/Z/P;c.=9c9U_^G<(B&XE-(P>VS:OHTGC.^3&P56[&F2&_JB^aY^-V
T-\.?\W@F@EXRH)&;Gd\O<GLB4Q066BfV+_=]YAVC<0X#I4GCK.CO9b-.((,>,X/
E4:=eNL9(d9TVY^\U/XZLd45=\Kg+8X4b4:8MG[>QJ2HDDZ#GUb0A94^<DK[0>Xb
\796D4P0(H36&(:6TV+TW5<BCQ69HJZ6#;gAdGD9XZ@NNR^aL:YU\7[cI#\G+Z<D
[-H&W8NT]YG@6:,FTHUW+FU8/DCWH0cNF8Q#L7M?\1N\N^K3PWFNSP0_XJ(LG9:^
H:/b&@aFK4;AaB/YCX?Y.X=+>T[HF<E4L9cUE-2J^Z/]CWe)&F8-LU3G-PBKgK0)
0a1]PV5E3IEOFgV813[1^HV;8NbE[7&d^/IabGYJa8_gS6/A?X@bCE\Mb3N>/Q(_
+V=]BdF-RC^QFWMcX4TN_3J_M99M1Q?]#Q7P3P&.H,RNRIE3efZ]LAMZ6?b/Pg)a
2K6f#5=IL;0:R#d7@a3@ZS-A>,c8_E@[3Tb.Pc[OW&8PG0KND;KE[-=)W=7a3V@/
YadL+OcA-AfV>O_Ed8/:XZaC^Tfd1D@P/6#2_;9C#E3BTVPCbBQ:A\M>R-F&/]2g
8\&,=d:D3O3;W4KJF&^T=eI7g5UQ;A>Nf(6[H5+[CJ5aS&LFS]I\[1+S;:YT4WWR
[:3?5\WWN+gUVQN+BeL=>TfXH^)JDfV0_e(ZX(/>_MA56DcI:W.>]3e=bD73I5W3
cS2E<BO4_bB69B)6@NC.=Q6)<VJ=64_UJ;-3JFH?TJ&.dO;QTbT,/bGY-a<eKE].
FM5bbH3FUN\Y:UfbT>_7##H60g\ZJT]1\.O1C5g[_>>\f;E?HY.Ue<O6bDX/N0W8
,F\.95/(PSY+]gD&IQE?Rg3P<b66fa+ZQU)O8D4K0CPg,SgM3cI8g,48Z970QPgJ
][DG<.4W0R]7Z@1OU.+L^3+H3f76d5/98PY\8[,/^e=_:@4GbU5(0\.F10OQaSQR
]&O1R9cRI5OZ4WZ3^^<Cg^M^#GG7<fefeSR4AWHC>703RHeSX_^M11bf,9JY,?4<
Tc-))1c:>?TR6@FF=]I7da5?X,#^Q?G42)PX^cYbP>3;]N9;9Aa0DD3YGJ+&d;W5
TM<8=[ELF(E[@=OReJQLBYIO]J97ZcY@&AB6b2)Z\g(^PeP:H,RBc\AG;K924VT0
b#?:,3dB\ZI3-+C&Y/L.RPBZ@V>KYSD4C-().AL][#_KJ9GMU5T/M.e24TUNY[I1
&NA2\Z_c?e@ad4[VfL+2B-.Q.1;HcabXI(^NNOO22=)#>d_8ZJfBAJZee)-587\G
J//g?(U8;F[@]7Rb)A7]<NJJRbDW4]?;V9O[G17eE[Q\\<@.1<<8;-E=K^YfaUF3
#>370TV;O-.?1(Web7SEPD\I2:K?0=3]B^M-<d/ZdY(@G_BO2+O5>1:+6Va]CeYf
bRO(bG#+VWBBZTgb9+J2PU1,1N#LNNKQI;AMC[BG.gZ4[M@OEKG&b16G)Y8X5CZK
H(H_?4)@RS?8M4D05?W5Y[Ie],VgH2AEd1AC>[:YeE)>WWM6+\Q#7W>W#L=#G&fB
:#9aSN==JadYMH6f0He^X?(bg=Q@1cM4K+ON.g:>F(J;CNM2NT)#LTYRDMS^Ab4c
/>7cU907A\3S?CVG_:<&V]5dCJ<JC>K0\@7-30\X;c(J4M&(8&gXX5@[6:G2GF/N
<MKITI+BY[c#T92A9K]BY</8c7(76P4K9-&^ZQf.P(aDRA<V/ZB&[?d-H@eMaCF9
T/eMWOc.5@=<HX3K7N^2UTB\EB;P.YC>GZSJeRYNY6I<][YV<>fYFHI63=@F0)V?
>XB;E5>BbYAB]-+VMDJKVC8aLe.4UIVJFVEY:+7#9I5bS?W;-K@EHQY-GI0.#bD+
fVY<L/9<6ZY#B;d&\EQ@,O(g7g7#Wb_PDUV0?]=NS\b+932[b-PW]CYW->39d(/G
?[=)JddT/VR+ZG&(JIO<-K.2V]/_#eDc-B_7<SIK82IT;9J0/,<KZUDY2a[XUZOS
?]DM=;,NISM^1]b/b^)X&-WOKAcZ)[J;J[ID23PT&;+LB9,Z<NX^GR7fcB2+1Ab7
2IWUSN7_4IS=9Y?c?(ISCZTgcKSG5_aSb<&c/Fa&GS4_BfVG,#VTV35.cL)+6\[(
QOCbPYCT7TY(_<;/WFP2Gg.?&]_B[00JOBD#)e4F9F04CJ?G&6cMc?_b^O:b7UIL
eJ.+24ZVUa:4&6C:@F[A]K-C)+<)RdWKcN.[[FGgF[=);-#B4M/e_FBO?e#4H?ZS
>>\D;[9]=Be7W:J&>Xa7;<<T7ML=84Nb+NDBFa-b>6=G7gEYXQ]_T4]gLW\;S,GV
dQ;ZfAHbGS/][d4W65ER#2/BT7NHSO>#<0K:6SA0\BIgBK1H.EEZC#C9<TSNZ<3<
/[]W#@6][?PeX1Y0.]1++8)>?bQ(>>:^Z2O(M<bdP<-QSQ4,&JZCc9\VO1AZZVNR
?.#Z_HOY+2JSL>M&+5?f\5_29?V0c_9f38>d5S/0OU&6A+3T=#4dM\<0X,N+2E?#
]#.E=SJF7Q;F5KF9@]g,L(G=\-6(-gI&9?@/H-VK.f,g8W,FRKJ<SdP]FfD/G4A]
G/2MQ_HJWNOSb49DY>]Mab7R@[I5L6G37W@_R2M^gN[,X([M]C0J2&_eR41F3?E5
H,D?4e4O9cW.,9XUAKE_Xc>\SGa(Qe]>;DG-3XANQQ8G&9#RLILPIgQE<&C(]]_.
@IAY=Q:)#8REb5@HT6-)>[(YWd]XS(dg\\O.?KUfe+f;>eR4Lg962RX_b]X9+H7U
^&\MOX])=d1.HJSUE6Q95<e<2-/3&)P4eV\c^Sg)/S]0&,:0ZUQFe5N[-\\-NdG7
M0I4C;GI=QEAYa1<R,cTVbNF1;dK/U_BA5=[=f#RR,9VbZF5VP+c(-J]IafQN9/B
JV(OHe>2dETFMS+3Yf7VV]:..5IfZDJ(K\Vd4,1G#HVKSMO4G>^[HFNIIGE.C?<L
)gYRXNcZ7YfgREQ.eJJX-.J6K(c.(G4TKfC7YU#;YO\ScXD35W3a2)_JS4].YX;U
7)[W3DCKRbT\>VEJA+P1Lc08\]50/3H0@?937Wg>?/60CYM83_=&McGD(YI)H]OJ
P4#M.JFF&eK]E)/]3X,EGQYVb<O;>CVR>67[1O9HHT(@/ZZV&C/7R#P(//16V]EF
[>cCbFSafP6Z8AEP;,fIP?6TEZU=8)H/1<BMAJ_Q>RI(,MgMS0+^8gSEd=U#4<G6
Y<(ZF&@V1R#(7)RP.@?#RD>_:(2NO2O4M,?B7X1DS<WM@=/\N[4VfT?O-5Fd-Ib+
CUO3O3,RU+/Y5CZ(MPUXKd2##09[,U/QX)f#4BAO8,7\Y670J_Ig0>>7EWc?>[&B
V=2#W+482e?5MMRGdd[\Y+T&VDC[C8cXAGOf6;:@TP8#A.TbH_7.VIdf-]74?g@g
=(gW>0++fNdMY0]@[T2#fN2X\8eg<4KJ\J6CWcZ>HS)/:gY&_7,D446PP@H0fa@/
N1EXP>LUO(#66W:+5&=58ba/;#ZYJA[#^MGdeG-,T@c/RG[8E.@#0L<Re7&a2^&U
EW>)GH?F@:/^-U:4]91#bW)(O2bWN4.&S31=M><6NCWe7c1J.A33L_13];>@0RSM
J7;58ZW>FJ-c)H-54[3b;a>YK:^E\6Vdg[/]A?SH-2+])ZUG0aedGa_#M0aNOGSP
J#-gB<.[H[#ML)d\[TETOfQ681a6a@U9LU19_SR:ad.HWRPGS66]]F;ZM#c\N_.\
QSa,#,@d?S\+O1/1cG+H-RP&15Zc[Lfa:((KU>XSOcECdD0:+6=+I^8@ZUW)1fg2
>\F#Z&^N\E(NG>J4]UP.+E@@M<H4C#RT73K1PR=dbRRSED6R;MWKQ+<HOD0+,Xd6
Eg>,I>\Z(DGV)Gc(EH5P_-:O?VNA8)\&TBKNgVc7MQ(/TKVBXd3Yg56[^SXc\1ZG
8Zd<NQ/?fB_0X0F64D-\J#._5B[1T)6+Ec7Y6OLGf&WJEa-^fg8^V#;,P1g6;^-3
9U5(?68TgBg)]K[1ce+9K[=E_TW>TJMVR4UPE(/Ndf)P])(18>42eeJLHY5f_aYO
A4_W[BV6ZW_effW.[/cO5?5Sf\IVV+40@I1YaNQU/J?:;MZQTLXd./2BSa^Nc]10
[b2F]aT+6gg_XHR^.bY&^>^+59K5LM:cOLMKU\X1&/Z-?C(UDOE=1O(G@@+SW&8+
598QB9f^9K,:N:_5X1F\<8&TBW36#\7.+A/U6a;dO2N)(KH@PGQga;VHQ6UASTIP
K?:+W)TQT8(15]:H]0G8KW@A&0J03_^5E/TeR7JZQ[,NZ4K[M;PgQ.>PUZO-,=S6
S)&IfQNU/Va]E)^UZf=^+O]LO;g&E6@JH:2CCHb=H-5YbbdS0,LT7G77,WLc7GfL
I&,H,/4D3.aPeT]\)K;J)RZX0:)OPE;KB&,);91@eM_Y)M#Uf-+a,CcZ-9.G=Y9c
GB@J3;Q92fR2:4VZ6b<?I2F;M<W1VKD?-1.g5&86S@?)N:4\ORXGZ\)7_5^gA^JL
g?),WabJ=AY[N(,)BP;K#X0QJLLS^V(<fRSED[XP34P7I+,F?>&QUX#MN?(U#P5R
>O:-\/V-QV&-bBZG6=E>+[UK3USdJ@<gL_E-5E]\=BVGV)d?V1XMB&C#;2f5-M^A
)P+@B8^<e&VLT<Vc8(SQ09)0H0+CPK:ZM_4.gdECT5N:8g+VdX_BII?6,CLYdP+N
7,:\F9>SLPHdI_+P[H5QQ(Gd3NVbBEP;O&b;J_ZQ<e4_5/[dR4aE&5Pfc9M=eG)7
^bOX/2QH0Q3?D=WIHHJ2:0C06WHMd/P>F/@PV(:#&A1:VE99_+d;5V(Vc[H3FR=H
BBS/dTV_f^Z<=QAJC;:NJcE49aIE0Q.NB<>g;W)Z#faa<MHY^/b>FY/6bRa&M]NF
8MYD;^YKV-L>OgfNICP\\4b6VgHW=SY=[6a<8I\fOR;&@^e=/)a7V,]#A2#H[BCL
_\W.fGNH<fK1H9THCW=038/-Y5/21bGUA&KT[NXNLb0?;IE7c?W:Je.&dKUJ]RFU
gCaRRHY6Qb\ZH3>>4Q,&KE2&D.FZG1<_II742C:(HM]T>?e<]XWQbUBS;Q-EV0AP
H:Kb5BL&I?;?^\W_:HV0BO&7&,dOHRg)II045N0)>@.LfOM_FXG+bg\,XE#P#/.<
5ZKHdMLb?T&;G>^9F@\CBT&=W\G[YIQC#P9aM_P1V=95F/_^b+4e+W9Q(V,3#6+X
\L,fB^4Q->,Ue7He-CE<5TcW5)SYM_K?8U(_B1e1:VX&FP6AM30#X#Y>Sf?F1WTb
TFA4D;^#bd=P?:_C3gH[1(eL84#?D973C4aC,-5^b4ZfRQ.-WAf>>a3^O;P&=.JY
#4Y(&XME8&?:c4MF4a+YH,B&QPD.2?Fc3OIZVG9@Ue,>)SB(JPeGY8-Z5=FO8.<e
dSU<))cP6S-SW(MC2(NdK(ZTM6?[V.#)E]02(=I+,/@?0d^378[<V+BW<Q81?P(;
>&2GGFQDLg#,.Tf12:G6gRe)>S&d;LNd]E,&DSK:;M^+-_,OQ+c)_:Z-_)XS4)Pb
PdgG-c>@:c49BCOGM&3/\cP3CS^dG6:a>(D;_c]fVdERRX;;dR\OTCIF^ZLC\aFC
c-BO2>]-_++DZEFJ]>.I[9L-QEa5eW:B^ZO5<H>V>8D=f)Y4;EB#4Q]S^Yc8eM^c
Q6T289f<?L[A4Yf=^@fBR:TGU#^N_/2HR-GRf=\^5@A#5J__9d>\HfDY/UI;P0SG
N9c783<Sd81/&A?YVTGN.].RH0-/@W#Na8AV=8I1[MEUeQ84AB>ZV&UH?cU5_:D(
.6?+BO_0fLL[5C+VgY91C#W15B[X@?T-XAN<E\99TY.^+ZUOH:>;-g>9b9YY[-D_
d]H=Mf6A#SF.A_IeVg((C7(aQg\f-,b<YBB^8@0>-R,I9=;;d>S_8R+&?2X1^M;W
WCOX<W+Tgc)MMSKGc#DO>b>fSYOIccN+A4C<gGdc-ea=6;Y<0J^^]fd&Ag4&&ddH
M63I.gV6L]M(N:-\?DeC/#cM0^@T(58a>=-MJ-23KVZgA3dG;T&dQ9/AbNV_<eGK
M[&MROX+(UJOgO(:ET=S85974ZARBJJS<0ZH;Eb(5:XY0,A<KV7Q;6(Za[41_-cI
M4>ZTVbM^D^/^5R,]J@ETY0T+CM/(0BJQ.:#BCN0d][;0Pc_CTOBZ>g7gWC38D68
KPAc7+3UQB<.ISJ/O_,:be_G^W^:?78Z]VZIIN]^H#)QLATI;B)O:FNPEC#?,cD1
]Ad+:9Pb^dPNW.98;U>17.=_2<.C>DXZPR@&8UI7:SP-bVI^Ca.J]c4Y4PBSL6Z]
I0b9-0(G;)]OG_O5/D?bQ:KOWF@bX\=T.Z(<1^_0RLA3CDH[QUdcAA5\Z.IG2>C6
AJ_\ARPL_]UU8@]H,f;+&512NM:K+-d\@<1N@ae,QU<)&E/E)3;=E-+SfUf=;2,a
JEb#/+e7_:GM1FA-N9P(.3J].PC3L)H5LR>_BReM(KY.P/(:H.2U;T[?g?0f[+VB
\]^G02e7T-\9[Q3^/9,2R?ZaNZ0>I9=X)c=_/;aA)PZbd21N5;C&.Ec\@e2[,_O-
7-2I4V(3F/,703<S+XVZ3HTFMJ=^RH7M<,A,@<F9=S_),G/B<&D8WBgU2][aU3_P
6OV2Pe\d1:Z0V#-a7:C(=A57?&<eM_J9DT+d6d?:(2S97dI?>W[]6e=QV2>[Lb3A
DbF3LRHe)BOWHSWN(R\aZA=TU/d8=RN>W#Vf[<A1GFE&XQS,^H]YP//H1V(a]T9/
]g)ZV6:(c+DZ^UE4><&-Z.S-O2dgW=J[U>KXU5;)2N6:;ZJ4GUZef1SYKbGdDfHd
Z)GfVSTO=S-7XG_f=O@=8(RXY2+7OMg_AND@,ZO.+B?0ID4+G;ISMTg=V@fEf+P[
5.YE/aAM_3Y,V?8b)@F8A+2Fc(+W>BJR<dPINPA51Tb&b2:.](fAgg6(0B68/&<.
^b;;>;F^Ce)Y4AO&[>U91DP?B07H>R](C)DJf5be39X74bc+24\SOLKG8FTKNG4_
X#Y&;;,T#U\IMdO31]EZBR8d&8d_:])HO^G>TXSG;>+.48c3agGN:KT[6[R<R#[)
<D+W&N@I=KICP^LGa.;Q&@^ICC8E1^#T&BMK.3UPgf\#STV_YCSPS_7E5f^2/@@8
5@Of4O-\53=cSOZ_/AU\fgE\?>C5;LSIG;eID/F>I>S:;/7VB9gI4Ee;9JIg:#fQ
QGVgMS=L^8D>.[AOMR=WOLD357GVB6\efdC:LBJZ@CH6Zg;N+-;3AG3;YB+@,#N5
0S-^8Y[>B+7=T+8fY?NMWeE)M?fU=^\N?)[+CAMb?#N:BRCWDZ1IGJE5>dY/V_7g
^PX_4U[_QFO#c)[G=^e7G66.,AF_E7^JM5KA=_B,CcH,[[g#\=DI^UHFK0NfE_9Y
G(R<GRBbW49.0feLa&SZTY+GJL?OM__->>C,AY]ZRZ4_9.7b1.<c\\0(2eY@T<eM
HT_<^\)]6BBV7WQ?HG0W-DB7a&JAd)D171gD.)HNO:#4@_<5/Q=2W[;b6]7^)Y7:
bF;@eY-E[1FN6W:^ERdB&\J;+W?HAME/VdFPY1QPcF#\5BRd76JVI(+5CZFN&E2Y
;gc+[b0T9_a_.g7FB]BNDdbG)M:7(-5YDT3\-d-,]]OXg]DU]-C3.+3(JOJ]W744
J(-2&:]SD4IL:/cf?W;DGV+7,LX:bdgNPGW/ARFNEbYNJ0:f##S>(cU]BEaNZd^e
-:(KgD-;9^\5G9^L8LGMbA[,S\?_8E133^6Y).UGRA&0[S87L_5[\C24U(Na\SfH
Q)aV_c<gJ88TeF9G@\MFEHU7)1Ea3M/@[N,1BA8T#4J-L;SPcdR)2W.S+5G3<&\B
OMcK]:ZM@Y:DIEEW1J1I=M1_@AN[,2^:dX0=]/(A1df.dZef@K+_+=:^N42OcNda
)N]IHAT:OE-:g0/X#2.>4Xa[bbNg;NB2N6JE9.Kdg=2Q.,85SBD57dXHUS;M6N-?
5bGI64c9f--;UKL\W+34WTBHVMbT7OS&gV9C\(1eC_V<DIA&,AH#8IXK&aJE>PWB
#BLK4YD1^[PVEL)E6=D02d)GHeNJ8:1>+G.c/aX1HA.AaI4g/ge5^8b^<OZ,Z=3?
.6^Ne_HcAZf+O@.&faMV#6gfc8L,0/SE[OK@TX-]OX41(NVA/\6Q/E?TGG56c,R)
0e/NU]&&,<SST.(:.45+].J3+]BSW+:;DYZD&J9d-N=aa8?:])?cLf[VA[4G-BED
EZe@aa/L0/F]L2(Z>AT135]f4SS#Z:/5<O.^Q4,8L2X2)g9J637Q+V]V11_><5]-
7@+IU4LaE0Fg5S]]Y7?YM/6/0SP[\H6QTMJ9IRAMD24,/L0P<@[gF0J=M;-;\;P?
IcYFcU2RAUC)J:&Tg9>OQg09QbTL.SUO_/L\J.dVJ0QQMXLXA4.H0?^7Yfg2CA8Y
K^Y:QG._MU\BVS977_P/(NV=aS>AAGS)LSXA)BgU\-N?^EOB=-Uc.g@MTJ3cgca)
-9GZ4E]<c2Y(?ZYSPR#VMAELf@V#Q^D>[ccS#dW<QW>-a.4,S)Z:RJ(O)W1Q?;AU
[GbeDB#1[Mc6aOcYgN[fXZ(e0B1.B?K,@_#LXbHe3U3V4-d<[XR=SSCODg^g>C<L
f44Eg+2FAgeC/FBYAdF[I@d_+gYfJD)JWdYa/RLQBaU.LRZE?A0E[_@S[f0]MH30
DQNJ&f[RGI4LNEMHG=BK_QA2<\-7QVg/J?Z6=Q\,5UHIe:E-_RFZ5@I3_]KeMOfA
N738]5H@49>C_GY1f5ZR<YPD2g8@b8K)E>fGB5]^._@(2WFOGfc[T&^01O0cFaN\
@JJRRc?U:B]MJH9@^a6@15S4_c4bU:JMJHPF8E,/L>>37@J[_;DU5(_:OSC0>_@6
A;51N]05;V/Y8)L\LD)9RMPNZ@.b)ZAJ]eI906F&C#^fV,^_FA@Y15c/59BX,)#X
9L4WZFg],SH1CD=3[HG[E8gAd+<@0CeANJQB27V.3#:\IGXP.L-G&g_KMHK^97Sc
^5OK?b&QC?RG2ba)c8OYgY>)d?b[[8KL\D5gVbNT(P5U>1&Y,[e4Dd)JB\\FHDY[
Q^V<=8@dEQ6dS+&O+g\T(-O]a4.EUM3c.:<^2=#:C\6gLF,ZD</TIM?F#<&L(Y(a
3?/E.2_U0Bd5N0S:8TdZ>VD;-=<,#H\\6Z;_&D@42_-Wc]_cHL>-1.7^?6g>>O<L
d,/Se^I#0IMaX?/Xc?]6C5e:R<RNf^fdI^CZIIFdH5CRB=V6EY0JTBI9)X[eZ08V
O^CXef+bH^HT7gHKOXX9_@FDe75]G._MQ./_1?Q73QdGc)R2=e?=I6DBC@S7Wa3^
c-5S,U[c;76Z0>HI@W3U76R_L,Q9QO9Q9[1=cAe95cA#e.GMP?8+b@JFF#BXCCIC
58+1Aa8168B^#UXeR\b[3=VcD,H0_[3WRYbN.,9_L>GE//P::g>431PfMgGA1fF3
O7FbFM<)ebb2&df3N<^XBMS4^/BCG9,@75_YUQO@b4A)LQD5SWcP7^-baaa3[JL.
@TP9R==(7?8]3_<FL/HdQTOI5AV[:ab<IA#PEaP:+OV967G;JC_^V=71g-NM6JFA
7#48AY,B_L/Y\B4=,5UOe00;M4EV>E:\^2;,-aOFe)UV19IZB7.42,D5b2dO.-N:
;QQSgN,Id?V?&W=GO__Nb@BRUH8;B[]cEE&XfC4T@g6DN4T=bbY4V,FX=EKC/Sf2
acW9K@VH[L8C5(K?92H6dB9O4/@.UOPQPE2A#0GC\SaUdEcTVMZE6-H#0T+YRU7@
PY@g,#ZHQ3WLDO1.53b&cT0PJ\S+gU0]g<9=HI)8c5(?57.bK+?;4)[FPV+YFWHI
QD#N2;CD>?e_#Cc-?>We\cC-;Ee#-H#GE2<,B41S3/-.V/C:6(YMLH(YM[BAP1Sf
4V@5DLN+#)d_T(O.92QB.JX5TI<@]4Ae9R++KTf46aEL+Z9@-(TCR0\I9)]CTV<_
TUfY1QcS2gE0SR8[Q+_(14c+f7/d-eU,3(G(DQN;VZM9LTOILI_H[_FU\[XVSI7,
XU?#55HW(0;,6LW(B\dTL+\QbQC+J>N7P&Q5O=[(BN_Kd,g,]b4Z&_g@G\Ce^9VN
[-\a:aR5+D<<7;IVYDAb9.<L=d(DK:+9H:06:0CLU<O[\/LK2B+RLQL8f9^V6eMT
PBFC?],J+-6acJXM-=0G)#<NLBM+EM3-\3;LbW1=)?4_XR-=),&4ec_5\N?,O^P-
3;aI[I5TTJ\H.7>.FLd4.:.+RR3TV[Y_DS8,DVfB4&)fbWbU5@Z.4;?/MG7UYTY=
49Y\d2&>L?RDCTO<]M?&c_Ze31<:/O_b,;?I3QPR5g43a6^baO6N@g(JHWSR3.g3
0<,3\=<MA4gA?/BFHbOKIQK[/8A6QZ7DaRcKS4M5TZ4^SdA9#39K]<+J(GdV#<&\
cVI[HE>^^JEgUDF]2b.d&IM?W5c\=4OH9D,_M[8@@K[?f&MJ-BZMLN,CcLK8)\0V
-,cd7GcI_ST>?XJA77KXU,;aH>;];@FD56[M-=Pb+dfaZ&S5KC-D95cE\HFe__+H
DCB=J7U6d,B+ZX5]MV&ca^N2EV[\bCRCL8-8c@fc9P>HFDI(PI2cL1X&>IFdJ/Jc
-WFCV--bI;W)(IbU[@@5JA^0W6IacN9W-c+YG99C6Q,)W]<F>JQ2X2N1T107C1@7
]+NV33A:Mg^HZG99+e5a@B)Ff&ULfYL4S+^<V;L5]5AZKUd>+@g:8#]aa9Pe[EHe
63SAb)O>0Y^=_Y7(;O1/9+MWEC4_^Z:04C3XAb]57?Z+98bW.,YQ8-JP9F)TM8L^
/\E@8c:;LCBJZ)NYa]9(d\AW)/2f->W4,5XEH_\@#83@HbIf@IR,4O_d]7.e/LU4
FDQ@=B]K4WPY?^^VYU6SGS,0PgI0Ye,gf,5+1@JZA5Nc]FX3SGYUSU>)F_HJN(H1
HDD&FgV/1\EZGXe30T:TP1(a?cW[aDfdB\_;,QM;Q(07cG6Q#?2.[e;6AcM,F>JR
PVB1NED?;T1c?:.O85d=eI>D711cZg6e#MQL1c)S-F@KDO<DE/e#X]H<#7Y8@,T3
QacLQHCJ&/C67^HbQ(RP3P2R?EMTa/9>U-[F[/.a,#gN8/L-6R?7ZT3JC=?AeH[g
8HGI2=ID8B/(0KDL)EP2-CEW)Zd8Z(CW]RfF(\+1-;XNf9O.6e2Q98:E:BQS5?RX
ScL<.J^IL,CdIGB-Sfc89F#/B/]>U\X\1Vg)2;Hb(NE(8+Me@F9fT]2,fg8a-XE&
]:I3WB28.4@)9(F0#SbIT^;/D>1-6-CPf+J#H87K^\?ZXQXc]:<+JT+UHYLTeX26
]#aKX>g+BIDN&-V.;WR1@>\SSdRVIGfdA>a+f\(IJM+MOL_XYQ>A:0@bHGC3._HV
&1(c)C<DZY2G</fMRVJ(B^#>[:2>A8O&4cB;S8=fQAcKFKY,6V/.L[(Z@X:3;P<H
3@)?9XOaFg2S_8#.UaEJ5>Ob7JZ0><LEb:&BMNGYP;cT6I/DYc/JYe(KU[[13RJB
+^1dHVeP_J1\[,P^5X+fc1V(]I1XKLb&^:@e#QREM9]]?S+L#LB32:R0.VPCeD9Y
=H>X<CJQ-+>8QeEd^)dee:/C8.[BP?XOL8PS3&_b5@eIZdJ>6UFBTd-dSU.</B=Q
N.XEM^=)<_<&?WHT/:A1YA.,TfGQJT@6IBR);>3:#T1.c3(9/9I9/0)g0<HR7QCd
23SbDL#RRC>8<Z,1a728FRQ^>]8A5#Y=aeJdI)7:)fRCe44I4:/D):>X7E/2RAOa
E4CUO9EQ59dDB?B<5[6+#+B8(&&THLEG0/:OS[N+c=/:UeVVZ[)YI=f=e4EDJ5[R
<6;CM#G2L6K::T,&W@UL1;ESg6J96<N>@]:D2FJ4BeE9;@9-0c;SWZ0==,:XU_D#
,[61f-ZGV5ZKROgJg@YaY#[\V(bH0Vg?e[a0f3e@V[F#^.@5b^BG09Z]+V605+LK
c65&,gQ9+R-+_1a;9LA?)D:B(ESW)&JIP^W.f]-V4d:0L^Kec^aZ^)33;U/;6fDQ
_=H@/.]b\EV?MAYf>;W-)3D)K+Q3+1UI:_1?M2Dd2O3fM;7)SBd<O[^T57T&5P#X
ZZd6X9,e@QbVO]M]S9DSI@EXE17b8OHg>B]CA#-VL6_S;.Y3AIM__DGQWRP<2Y2f
AI-AKQ.H4P>#DccHP3(W#AT_Pd#3)QXHAV@/EDdQB?;[79fF.#&?d3/g81XVZa@A
S):a1WH5I(+S@]\:E:E-d^;M034SO[.LF>a8&ePVgd:CM;O^)aGD>/=>.K/@bUPU
:#^=eUgPb+#\Q\Y^4BEG9&KRD7X-VW8P\I4f@bR-Y-@G:7YI>>8eU:1],;8M=?ST
\EBYa^N8MdIPI8N:a(60RJ>[5QMJcB@9]CR>BF3^@MRJc#3SD3=@b8-f4Q2<Q;-&
Hb63XRLW7cVMaWSR<7(H[,RUG\X\Vb>ecD5^Y2)/X?>FE&N@;CC.#K:VG]=@8WdD
.fGCKI#_+LM_@6B^P),8@K)6OWcK_,_O:1Od&0NNSE49Z)C7,FU^[JS#8#D,A)-M
B@_VAI.7-BfbOIbD.-,O^U3\UC&Yc5@KERAcg]ceO@G(XVQHR?b411XDUMZMe3A.
\^.4J_F.)#<T^B<4)(@N;,V<)=NS(aF5?@@O2M3gP:H:aD]K8MFKLL0GO;@&T]RR
C2Ig&J37B^+dSPg\RQ4&dW]IVO,KJg^6e,;7DS+Gf_;3b<6aEfRCbP37RFA?.g(K
056SZ[[>:-D-B9[#9X.LgVS.3MZ3dg>d^:T.N)A4VJ(#,U_3:=A,SE\g=^AMY0e[
JDHL^+3?)fK9G99.fZK3#=M,d>6JK/g>B?.^f&U>_\?7eAdFQ7;MQN?gDQWUD<(Z
FK7=Dc;8\D.V2+Md@QV>7IQ-ScZBRf-IBd8b&ab6>\(f;D/Gc9?B4C7=:8(fd&+H
SB+c]Z.AP8bK[&5O.cOR[WL-bM:[IGc>gAe-1b6^NZg4&8PP5D&W[.dFAEe_d9R:
:eF?X_@U8P,0-?E1IL,[=d]3g6Og=954Ba(TWB[AB1V3568XJJU5^.K^9af8+QU\
RRH(J33#3179(EP/>9d??@_W:+Ie.FWF>g51a5SSTH_YG?3P]B79Q\C^N?8cW9]P
L47X.OWbeVM1.4+HP_6,JT&X_;8^MRHe=SQK6B8e#P->g__P^]Z[@,O2/6AdC-IH
I6-cbSDA[ZII,H:[_FZE8VU;>/MVe55cALPA[>P6Q>.;=b@=0>4JeG,Pf&[NPTT0
082#Lb/?aV70:@.F^RgJ07+(V+Z]J\D&TVRc:+8:-@Y-KC/4#9J^7AfWVP.Y5O:,
aT#>@(1KZU9H@TONdU;=La@0ZDU66NI@bIN+:DA,<5g.3fB>[3-_]:[VM;gP_G55
RScdU98Z#D>aKM=@.9W0UG&DeO9C:EQ30c)?;&CNA8eO^-A)=DXR\9UKGCAE,D,(
MKac5gW37=U2E4\]R8CH.>G5>>LW0B75>HA^La>@.6L3bT)\N._NE6K]dcUGL(f_
DZeLC,#_LT)65KFPOJg,4F(:6c#dYMDSF[g5Y4&X&:L;Le?90RX64=[DYe.[^BFZ
G<<Q+JC4SWa_YODP0^8c6;O;Ib-fD?0[cL9/G250M5P7e7T^?@>ZWgS5I:@D:gAJ
5D/18))K?8[BA=fSP5ZQEg)S(X+e@()5]2G8/O[3C6KXF5959EB:CO#7f#/)DFZN
@9cRb,LP_G6A_A7_e:R)\,8BKYVS#AfQMM&I<W=\aGN1V(#J]>1JBeJ>SgaD<76X
IOSPA<f8c>^PEcY>5>5U7fOADU8f=J:R6ZaY)8F]3LcDC\3?LdSbL-/:,&Pc)+d_
3c:2+I(IJD;X@6C^ZK1gCNQ\=Z9g^Bc=_ZHXAT[6gSN@5Z6<G7J:).(W6>3_b]B]
=Ug\(aDEe.[I=Sf5@c_1H@C#Z,2QF?O<5A?#6#EEZ7XI^@5;aU,W0EQ;gR8(=83F
Md158bY.B@cL<3T8eM&=AO&Ia;+VH\#b(RD3(+L^B+,aY:c9;&EZ^cYW\5?(bEJZ
Z_NJdZ+^f,^WaR#V=?SG:PJ?M3Q9/;7>,>G3YG.d5WMSD\3-19=^LKGg5J2]#+.V
?+QD..?EQP5PL//(+;S9H(WQOY8:136@>FYYU#:.c,],6V>eGWOP1U0M#Ld(H:I2
Pb1VcOS?E]=HVMH&Nc&M5-I_1-_e8()96NNQZ\3gSD8SR>Z2S/D_G^JDbYW7@RFU
3(g,K.,]2,6=AZYKa@>5,@/9ELODa2:PBbBH_[[.\8;Z?EdQ(D4NL,NZ-#+NKTQ<
SdIg>B9Z^a7VcHAfTZ^62CF+8(MFgA@E4Qb60#2&<NCDTC#2GQ;K.c^>8@P@Sd+]
RN0CT3+.CE)/+-5]\91DDN/KGJHgH7+FYZFMKEI=\c8+g?TECgYGgN<9T27fd@a6
fO:O)\M[^8Gf6E1GCRC,Z?Q66D-=]+eZ^D&,WICOf;E2e1ETLE62)@b+dQB78YQ?
M^AaP#-QL=ENWc@eJ;?F93))EV>3XZ<1Le-R393X[MH#8)UU73.;&ce;BTR)Qf8Y
45PHXBLG,?c2CR/>dX7I6A^2G+>Z)8__0P0A]60=O73,I8@e,HP0PHd00=NQ\^^]
6V26<b9Q;9C=YL[_W^&fF7_;1&3[6Wb.d^JA2^8B0WdNLVTES5TT6D?L)OD2F3]0
2PZ4IA+,0L^/JeXeS#PX.UaVNX9g1Y5\dg;aY<O_BVP+G\^dRg06dNQY>b+ZX.cG
12(Q0YcP1?[J>3,[-.gTg_2NgDTJKV/T5E#U-Sb1^^2G@?WW77+CS5];JN9E7X\B
3KRR:#M0NN/DU:2B_4EM;KbY]?9;W=^BVL8PUPL.W^S11d/_,R&=V?VR_.OdU86\
D\Za,/;8QNSgE\Q6N6FT9^]Xce\P_4GI9/,2=Za\,<<7<W?OK6=\6#DbLVBM[5#>
38?aGd;)BRK^_QD6#VdbWGX>g-<Re4@_?C^6I83]&SL@@gWNO^e\C/.5VF><Q?K4
#Y=(b]3-90g_:B<X&&N>;C^Occ^=PY0]Cf6HCdc)L:AIAU[MKQN3F&EdX89+@ec1
-=1:0A@]LHMPI9\a&E+>+Y>7RE^C,^R8e.G&E,Q]D.Y),\E[@XS\(7aC0Pe;8I8R
B(@^:]Gg(6^BQA4Q_@<)3[b?\2T)8IF.0B1dg(&UIUBD7NHg]FE3NV@BBK?.WfZa
6BF.NHb=6Le^(ZcIfMe9/I;HOcZ6.Z>W1Y=Q_3_5]FYU[14<+4fI+&TFeQD;UB31
QQ+<7>^XNUda/&]L0)#(6QP3RFc\eGJB>$
`endprotected

  
`protected
PHF.,(Df=dgY5d=?a9BVgUQgQY].97I0T1YQWQJ=G_1P+DLUeB5#1)LFW8]#efJI
K(aEL+\3Q?-Y,$
`endprotected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
bHdJZ;CCRe5P0[:3H/19R3g7370_4@)C>^:8_U9Y;7[(7cSL\CH#/(5HG4<Q<EGP
@N.\90f5<G/X.56/8MP:eNQ):\>2d[=&2fD#FN8:K@Y2^(=@?2a9B(=LP4d=c<d.
S&K5FP.=/3[GU75S1C8>C3BaAC30_:3A+6&,5@@^Z.1@AgS&H(e?IZ9@/<=FU,E/
=G0JDTb?U^W6I^O9bVQbN+\D;L+E-3#9RN5CPRND+@ZWY@+5>&)Y1CI.D[#Q.SR=
GH&;-EQ.3?Mc.J1OfTM[^&N)GUJ/62LJ<$
`endprotected
  
`protected
Udf(=EJWA_e,N5N<[f\I3&?YBOY4W\Z@(<gTXeC2,N(2N.I]-(f./)\@,GZ5T([K
\UPDP<65E:O,/$
`endprotected
  
//vcs_lic_vip_protect
  `protected
[Q?9]eQgLD:.H&GIL4,OR&A8ecG_?WRSc/1D[;18]^;54bUR-gMV7(5_6\@cgBB;
==aO6?>4<^);DdM(&9f9H)#?3dNOE&)_W+IG]DcR,Rc6(B5HT;-V_R\Ja/+D+<PQ
+M+MS=AF5/S>9I(GAYcN)KRTfdeg.7I9gYS#da4MU(8EI^W-/&;U@>N8FWeS]#YJ
Q34I?-CaUOfE7:8H3L2[6OF:0Oe,HM/Xe=Q9VIXb^JUT?;>FbZb<S0QO<^NCM3Ng
=D:ASYXW4846B[&1REE+Lf68E^IJbNA3VEY7YX5WGTBH@;d1gBX^(H#;Z#_>C,).
)/VMI3F)TT=V\7b:FaB?<WaWe(5KTQ^)=(U0^;b&>]^(Dc>,#d3fJ/OaIDL#S_D3
=Z-G4Y8E:\>D/Mc7XWZ,L2YKg11R>Vc-Ha3XJ;-:;_WM8c..Y5df\]HG9#7R-A91
:7799XZ)J520a.4CQ6=XWcC](9.HE&R-49B@A?5efBAW0MC?V6&S&:PM[YP^)cK.
/N_ZIdT_3?]\-K2Q9:(JVDBG/1.B<\>:W=\>V;YR]2dN@<LPbdS&O=6RcYYEEM&0
=#3c9KAOLI>([87SI58P4M=X:N7YB(,8X8a0C9QI-1+Ue7CgM8MQe\Tb27d]1,ZK
5.X?#.5Q0ES)fT7#.37XXO4B1E[]@aQJ-/ZMAW#E9g/MR3,f=])c04AeN5_bS8+?
P2>5?&JJea4E=]]&9f;C:F#LI-+FD4XG550&8^,S[BM(OMIFgVc]+b]>IKd2VLS<
fLYc^4>MN11=U>+[(1^H?3:\7.OL\HOddV(2EK2?3aPN;9K(9WSH_P8b\&-6+G]V
Ze.G\+NRQ(+WAFUa@26-H#9W?SN==CX;)-S]&F<)a27](Z8d+9U.5LN[A&_2PKRf
7)gV..;&-=V\H]7[,_N&SJ+07(Y;1bU38-3MGTa,E^#Z])_R>9[Z=H>8;G<1<,<^
P3+];N&SBX+ZIb#).L+c22HfN:(D,QZP)V1T:&SF.:gH7bTY/-Kb@R.?Og5V^T\W
BC>.G/.M;>Q(L0HO\<PQF+HgF1d914bC<TD@O3fEP&MH#/AW3EgKUageC4=RL41E
-cXeS[Q2.UEd+BSE5-T0c(-2EL-bP9d3c>JA]R7]KKJ:>?UONK]3PXS6IQA4(c33
;W6M@1(/>,VKICKFTREC9>^]dcYRJ/;5e)II[RJ9<C&2Ed0EQ6Z>f6B8e2L7=[Fa
+fee_g0.3-]KN;Vac0B-9-:fa/3##TgQNTcTL[T?C//7)_ETGLLd/<9NXP0:19e0
2OQ;gC\B)1AF[=)3CKNREW,ZJH7)<<9XCQ;X[-R+^OI@V?/T]FNDTZ,RX4d40UY7
&RS]&+f_0CEAW0_A.eVQK(FY=[:G,U>,[gV5[9OB4LZMAX-Qe0Y,fBa5L;5A-(2T
_2=T_\g6(\<b<JUNNgd&32aJXDDSE0#)bY;N[,Sd,+EF8V=/7E70cY#6W)YS(<TR
S5Y+>?PG-D.Ae0X1OA1361J3XBbOT#O@K_5A@^A<Gf+aABWMb8/@gF7eHJ_d42MA
ECb=&d>N7.-.dPK?9:abES[E8C+5MK8BZSa-C41#SG&-RQ@cQR&#(036)O8PEf][
BYT>R5M#MCZ0;QCf>QDCVaR+#L#WaH6NZgL1&gbW0T-,4c_+.JdZJJ3fV]7,3IFM
R+L25@-]X)<Z2SK#>.a^U^A[EKG?Kg.D48\1DVR#agTBDaMF=.P^()NcBKM0/cdD
^7)SZMX<#,V^>AMF2<bA]G5c<]6;;A)db\JcX_33g[:IO;M2E/M-e@S&>SKg1bbT
W6ET1DG..OLW<Q@W;0R#5a9X.Z^B_?:7:ag2IMJ3]W_e/K&M/dIB6Q.REg^Y(b]P
O84=34XHI^C7\FK+]\:?d/]XMQ\8S<[D[3bCR).[Kb(cU<Nf0^CE<(8LW(fUX22C
@<TD;-Y5U^+YeQC:(DVACPTQG3dTR?@,\KU0Me>_gIV^>S>\aa[/Z?d:H5C&88B0
bT=?RSL\VO.C#&4FU?.U++a3Ld[D](f<B7\-5>70gZ6_6Ub)-Fa[&L2EF=3I@Z7W
TGFJ+dGf;F^:/f#I6K#GZLSNeaKgD\L-QLEcVJ0Jcf)a\gb:JEf7cNBMV077W&&@
3F_B8f92P;MI[IJ]OPPfPGZ<-S(+Q<,:cgPAbc&b#&9c5P>VH[7BM3&G7NV9(e=7
IT_X>&S&&NT_=378#b)WV#NR?Z@F.K6-Ad)MJ>VC\0XEFG4\bRX7+0#&HI@(HcJC
,6N)43f,<@>YfZ.H.4f@G;AO,N0C_:[#g3,SC&KJ(686]6b0M(<=@52GNgeBSMd0
C64BeDc.R95U/EGdT8VR15Y;,7=UG[3Q\8W/T#E;Z+H(UU+;U/eX35eKR#cB1?RI
J1&/6K[J<-/L33[>g-.&aI)K#RC9XgKaSYIFN^\_BPd0539R8I@A0)3=)1GG+BNg
YTg]Z]7(a<8\H?O3F>8A.4WER_^eWdII-)=5/B9&,8BR@.9b7W6\E68Ic1&RZ2@W
#ARM5a?gZA<P[DN+6-X=Mg4H]2,VC#LX7;#GI&-.1]@d?eBK)8KCLf2VRVR0A-.)
dE?:E9/?5>YQH&O<.U,eE&[MQ\^[3?3C8=?V+<L4B#Jgf3#eF;17PX[1.NGF@L\2
Fd94X>#dbL[NNW;;,.1,3(&=8a/[))?dAeL]3a7S^R[I4>AM=F-;\LK:OG:&;77D
.)L)_S)W+LNT(-_bMI7a#YMG^4S>a@;YI\B#,2O:-WW+31-OTA&K4^GW9fY>U,ID
V)Y1Be]ee]OXJFQI3UCH&I99/_4e#]@10#6S95dHLK]I9NS+2b<b&\dRPD<IM=3Z
R#8Hb?.-a>1^T)(c&TPI_eW<&=Q,#K.@P;b\YBg_GZ,/S^L<2-g,HX.&^6CBH3Xe
7\50#:.[_f+eRB__C#f+YQ#.N\#1&)NT.6cJeY5M,,?a,1=fF^LBCfMCRdE.dN=a
5GWVbe8L@,?4VNP3R6Q>1<U?>Gg71H&3FO/B&-H\XE8fG=[=fc],2XW(PWJIIENc
dRHN1U)0JQ\Sg:BMNf=9Nb5LNK?A.GLT,]:?VI\2NNW2N.:9SG0U(8:D2bU+Z=LB
H)Y941IZI&7-\KZW;3=/ZP]\])^IDFV]d0#.g>CKV8WX<c?W5E.3<&U3Z+,:K3ab
=\=0,AV3LGM_cA/bPg?@A61+HXI3=&6SJS9Z?/+1,^QDY)&NW6\0\U[V,8<TA86I
Zga5>\b6:3A4U/Y0TH4Q,TfU&TGcQ@S#_POBO&C][=e_<19C^RTKc<W>(c65ARR1
VGgGO>B;2N-Z<&GEY1B\.;ag8)2eeYK?T5SW-6UN^N^a=g)HOX/)IJE]UXL_2S)C
,-D/PW<L^A?cZUS5:dd?]d=]=I(V^X.4gG@dUE=BYGgQb))/HF5g]<e2^UT=_6KB
7CS\^?Z2&.6;)FRgS.9/1Cd/29/9P]C40?4(GUc(^\@,CeCd]1;CR&K-:IT5bO2d
C9EBa=7STfVCZ(;&>fXB@(9B^8PU:54FFW@cSeOWXcU#9F_OLf:F?P^KK,<S)^CV
2Y0?#0,^MebaE#K[&a@2K7&d6O+/(fX-V7+MKBH^U/+F)?3.9b+f4<D_E>@#A?Zg
T@0L112)/RR)^PYc](X+Y.(\@]Q-?#a=ZZ8aSI)Y4_dU?MNgL1ddg,1VL1YP05e;
:g;AKP:]\B[51G02:+=C()gfRDa6Y\GKCE@dTZ.4[OCZ5@YO^<PI,c6)Q,>-RV9J
U0@68=/=-=85[#/8JceX]9U=:<8E>1?I\[1F-XdJ)\cK6RTPE()8NKN]4(HTW^O7
#WF?A-SZVSTWXW#RVV0TSOa[>V4NUQI@U.Z/Eb>S(P(V4>.UB^HBc;@7IOA-YZ/W
faX<?6TNF&B<PV9B09cQd8J90-7TV5D7MSNF;,F]OH:>P7(daf&Gb_+,Y]EU).MZ
d3BaSOJQG[UR_&>dZOdP17SOE-N;85+RfWHP,X2345ZPH_VT=I7U>-0:;/#VMNV^
fS];14eZ-+<03+29#b,_Z8IV6^&F9A>d@VY]&geYIG_YSEHS.HB,8M2aA&J_K2]O
HJL2c8=NUg#R-G.Ad]d7AN3@5Of<e;ZRT4dWB@)+8CaBb,A@dWME)HfKd&dMVI^<
E>7,OcGeYg?2fV2X@(84c\/\7Q]5e9aT9P)_OCKQ5J-=PF?4OU:T6(g#J=?-T,Ye
WgU3)eG4RQ>UJaE][YfOO[=]?OR>0P6P<P^_@S?;T],<:<J/6<O6#P9g[4:<9=fN
=[J;\Y\&<5g^M765#fE^@>7/aYA5GW[]cL9ZOS&e\5&8LP6JU-.U/>&e09g75^&V
U/Ub;?1EU21A@R@c^WRRGA6A8(aRB5^7f5N8B<;Q<C3@OD4+4#<2(a<.0[bLB4R@
2[YWO&TbTQ>&:VXJE095_#O-Wc0(LYY35CRA;UaV>D3<U6(0Uf&R:)Z#YW9N:\cD
8ZF>\a:8+6_3gL;b,2)YHVC-QBPRQ<C5NQO[]HWV]/FT1V]Q;(V/\aEM3XE=#XU1
?)?95]QKLZ9QJ#5>-OE]E>>D;77+)B7QQ3aJO&G^(].R4CDcR=HWfTD^O3UcOL--
>ZK@6LPWGALPX;Bdb#8S]5I[:fOY@5/;JT3X9cC1@<LO]6?>D>G9gDS4>=V7S(Ue
A&5J[Lb0CF=UOAR#HE=JD8JBH]1YX(FV)@>bD@:O@DATeBgWN(NGXEAT\JZQ1DH;
A7]<?X\OOJeF[;KXf223/aT.ZJ(2ASKFF_9GO[_W=5_BRM(A8/e4g(U#+ZHG+@SB
2,OJJY/+8JCF3Da6_6f_^],5,(>e7?:RSeA3#8d._;d+G#D<^+KPe;c4d0MWLHVU
39ZcQMD]<+/+,CK[g-IIUK[SQ+GB#>4F\_gW6-0(;5B6OQ[AcU3CF0L:W7eEa#42
fE\O675AJ7G-HN4TNb?,;;f=&V2M.2@E0a<[<b[UR&Q9&gaO>dX&O3dG+=L^3L\U
bOV(WGG/8>CWX1WXX4.\H4d&)SV<Z8&ULTc#VY@dFSJ12P-5@.S6.c(OL:>&8KGR
d=5Rg^K4EC8/\)GG1+Ob][:A^d?gb5d;L<X,A/.3R0V\gKEAYR:[7(4IL[W6J]&F
9/;1<T[<5)+WXIO<_Z=[d+X.)eV+:KIJ.;A0;06WJS_g#g/-CLTEO?Mec=4e2HBC
8-Z0M(,a9XX\#F&0QQ&Q1ZE;4ZX\945c@Y.M&EX:8dA93RHL@S.8EIb]8QcGd2Ye
Q?4L#YHCSFPP_L?dX64A<faOd,S^TBVR]=L[)R43ZS=&OX4;0)NB-^6,+3#S+ge<
fA\HWQZaZ4Q>,fI0P[J<Z?HaX.H5JR4:5-PQ+d-6A[PRIOQFI]<81e:Oc9fT./G@
:QH]65P,cL9c:db(eSa28)b0-FQ(M&7DE,P:8+c=[4IF1O[.Q]VQa=:OP$
`endprotected


`endif
