
`ifndef GUARD_SVT_AHB_SYSTEM_CHECKER_SV
`define GUARD_SVT_AHB_SYSTEM_CHECKER_SV

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
etvM4tY21jpBDFraLoq16WcyGrte7fmp+0FW6cdIc+J9W1DmBoZr5nePhsgtobXW
WfuRhxd4vXkBZRw8c2kpHPgLiNDN86biJVSLO6GONa9GGYWSbdm/fIS7tffe2H/n
CsrwVihWMBfv32suf3vPc6VTT9Gj80RFmtSJLih50iJhhRmAQxxK2Q==
//pragma protect end_key_block
//pragma protect digest_block
qPDEaRkiSPjWLb0R3TY2qapBuYY=
//pragma protect end_digest_block
//pragma protect data_block
DCi+dhseG7DNr5q7P3O4Nx2mNyFvuB7ohZt1X1YJKKLyaiX+uDJf30QgAKyD/9sD
KWcBJeRhA8uhXCNgvKkY+aVSZ/kZbWNeT6lf6Ruk2NkuLak1kD+gDENcWZMHHqai
5G/PYfFYKJQ6luMFpBXmcedzRMSzWJMoC2h0aAIJJfqNgqTcFTAYyfwQAnZOQ2iQ
v2SFAmrET0j0UuBMzPFVbTZXcAdxS2vzEvHT2mv9M2ufkNcKgZBjzllY3sJDZ4Gm
eYP/AdT6SpCESjtD2NMwVnJLGaXlQ1lTwFJwR42tmK/rEx5S/DM4/8hrkkNaUKSH
UHb1q77/IQwH2b/gf+D4go7/OaOm/0WjsRXHgYKhIqmuIYLMo59K6I9ydXGTgjBJ
kb/kVSfypjKs6+otR9pQYGVTHZIXvVQm8tlCD5SXkEl00Qr/OhtnSYWTvD+utOGx
qsRflAj06PG2LavtySI8l5C4Q38Fipp+T0OQPPaWSbyNtFijmDOKQrmcaHxLprFR
RxqmNeSvbjjC9Xj+1aOLTUOwabTI+Q4LS7G6Ek6vbpC3ErCVIQlTEwPfuaVYs31J
5Z6Q1rhYPD2Ea/jqfbUXYWqFCbmg4Z78gJ4yGqr9iRHzhwGQLz7ylY1h4S/bipVo
uBBLJWmlKcyqyGPrcrWQWwjFKl5dSldutwXia/sMBEwOu1axyjLU1xk7LI/B4ZWa
1SL9D+ZOQMdKXc9snXllKvOjBFUUtX3I+TXJ3YnCdOIQGcE3uYBEvlRtoAvzyNcD
Uksl74NCxyRu5JxLn5ij5JxbfyEiz8IJxe6Wa7uWeI18PJFhAUPpYwFg1p7YHKyK
jv+G5+9XEhvaT6UENRIVRpH9VCSG6oy8E76x0JFj2qvMHredhtygMQWjY6oSoeno
0+D09ajbHMxmOp3sxykasv6HyuYnFaFIEzTDTVUhXZrzZZ0QHddjlbQxTz6mUbV2
260uYv53TTmfyYhl59anA+IKleLckfQAUaSbQGS9mCpNi8LiFlGYLs026gZWr3Fw
fVAsN+8JngSnVP58CAFFOsgwpU/g/Wzr55d4438I9ttRAl+dFp+3ui4ZI+GI5T4P
P9ej9mb1k9Lu4wnkML/1xiOB95NRcw8E6kq6NN5FVc9i6bAhIdgJasOCOkP6IBkh
6UfIGBAy3CtHYHt3FKIUMQwnNFLvHMr4XftRDT8R0PXvYMWXjtz8iXbZp5nYwLHc
pypjxiiCVBRc5WOz60pBFo5ieWMH2rUot0aUtz7bIAwBWqr7Lgl8AfbtXkyLvpMA
Qk2eO1cSMLm/gt9//yHePF+gHFRaTgYc6VyS8Ey7zdMNj3uVW8dxezOQSqHBDnpa
vm8sY1bvQg17rxBi7PZ2AMYxle/J+WiHo7u6EMG+08DRaIEiyiMzo+pnrVYp6uxw
zFa63h0KjIQzy0GkTXhFnyqf1LCbtSLLhIeeED11AMAzmFAlBdgblD0SrlZUrNwQ
JzQBjOL/FgGbWDsUfef/QL5biQcJi77gxG1syJtYhuRGYJb1/eeEvp0qxUItjMVT
QyuqYFLuK3caPI9YSX7PgLSkzGP0bF3kqNGcBnl13OubIL7lUsBsvodTjSbX3Bmz
Au4RPBrL+1p8vLW81AxVixa543CLBd4JhZD5iLYnTlHH4S1MPDwuhsPy0IWafeR+
VqVgnsg1hEwkffi69nRwiyCcz+g+mxoGnHODurXWRwxs9JIfroTqqLxkOZSTILp6
FPCcgFPLlynkhSZE+be8aIX8oHj/295/j2aooZpYNjOkUd1aV+C4KRUbQ0EbbbYL
rpj4zK4r2raFQCby8vo94sbjtJpWKojU9xIt9rYKceytFCTETEjkUeEZhgAUSNQp
lVoNt8yGQFmIe8cpYTM6jbCi1aXoDeiq7tBnuKdU9GxNw6c7mugT1L0woeqhdSss

//pragma protect end_data_block
//pragma protect digest_block
5fflzQXB8FI765A5bOQvwlx/Sq4=
//pragma protect end_digest_block
//pragma protect end_protected
class svt_ahb_system_checker extends svt_err_check;

  local svt_ahb_system_configuration cfg;

  local string group_name = "";

  local string sub_group_name = "";

  //--------------------------------------------------------------
  /**
    * Checks that a transaction is routed correctly to a slave port
    * based on address.
    * - This check is not performed on default_slave if the default slave is set to -1
    *   through svt_ahb_system_configuration::default_slave.
    * - If svt_ahb_system_configuration::default_slave is set to a value
    *   in the range 0 to 15, then this check is performed on the default
    *   slave also.
    * - This check is preformed on all the slaves other than the default slave irrespective of the value
    *   of svt_ahb_system_configuration::default_slave.
    * .
    */
  svt_err_check_stats slave_transaction_routing_check;

  /**
    * Checks that data in transaction is consistent with data in memory when the
    * transaction completes. This checks that a WRITE transaction issued by a
    * master is written to memory correctly. Similarly, it checks that a READ
    * transaction fetches the correct data from memory.  The check assumes that
    * a transaction issued by a master completes only after response is received
    * from the slave to which that transaction was routed. It also assumes that
    * there is no other transaction that accesses an overlapping address during
    * the period that the response is issued by the slave and the transaction
    * completes in the master that issued the transaction.<br>
    * Note that this check is not performed on the transactions that are routed
    * to the default slave.
    */
  svt_err_check_stats data_integrity_check;

  /**
   * Checks that the decoder does not assert more than one HSEL signal
   */
  svt_err_check_stats decoder_asserted_multi_hsel;

  /**
   * Checks that the decoder does assert atleast one HSEL signal
   */
  svt_err_check_stats decoder_not_asserted_any_hsel;

  /**
   * Checks that the arbiter does not assert more than one HGRANT signal
   */
  svt_err_check_stats arbiter_asserted_multi_hgrant;

  /**
   * Checks that the arbiter assert HMASTER to reflect the Granted Master
   */
  svt_err_check_stats arbiter_asserted_hmaster_ne_granted_master;

  /**
   * Checks that the arbiter does not change HMASTER during a waited transfer
   */
  svt_err_check_stats arbiter_changed_hmaster_during_wait;
  
  /**
   * Checks that If all masters has received a SPLIT response then
   *  the default master is granted the bus.  
   */
  svt_err_check_stats grant_to_default_master_during_allmaster_split;
  
  /**
   * Checks that if the Master has got split, grant must be not given to that
   * master until slave asserts hsplitx.  
   */
  svt_err_check_stats mask_hgrant_until_hsplit_assert;

  /**
   * Checks that the arbiter does not change HMASTER during a locked transfer
   */
  svt_err_check_stats arbiter_changed_hmaster_during_lock;

  /**
  * Checks that the arbiter keeps the master granted for an additional
  * transfer after a locked sequence
  */
  svt_err_check_stats arbiter_lock_last_grant;

  /**
   * Checks that the arbiter does not assert HMASTLOCK when the master has
   * not requested
   */
  svt_err_check_stats arbiter_asserted_hmastlock_without_hlock;

  /**
   * Checks that the HMASTLOCK signal remains constant during an INCR burst
   */
  svt_err_check_stats hmastlock_changed_during_incr;

  /**
   * Checks that IDLE transactions are driven when the dummy master is active
   */
  svt_err_check_stats xact_not_idle_when_dummy_master_active;


`ifndef SVT_VMM_TECHNOLOGY
  /** report server passed in through the constructor */
  `SVT_XVM(report_object) reporter;
`else
  /** VMM message service passed in through the constructor*/
  vmm_log  log;
`endif

`ifndef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   *
   * @param reporter UVM report object used for messaging
   *
   * @param cfg Required argument used to set (copy data into) cfg.
   *
   */
  extern function new (string name, svt_ahb_system_configuration cfg, `SVT_XVM(report_object) reporter);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   *
   * @param log VMM log instance used for messaging
   *
   * @param cfg Required argument used to set (copy data into) cfg.
   */
  extern function new (string name, svt_ahb_system_configuration cfg, vmm_log log = null);
`endif

endclass

//----------------------------------------------------------------

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
YEw5Vn71OTgBuxZtQDjHdptjBmkUyuqitrFEiaij5jDCe1lErRPkZGwjn1s/5jLr
mIOr1KUZCu3HgygCYsBEMgZPvpUfE7G9BLaU4YNRUAK7u2vvpeD28EtW32cXtlck
WOWgkDRF5Si8pAtXnPPp0qTnFcew3dnIYD7fo+d3Mtgn9cgf5JYhzQ==
//pragma protect end_key_block
//pragma protect digest_block
5xvZPNC+RdircFLicv2B7m2pEgc=
//pragma protect end_digest_block
//pragma protect data_block
BfzhLLhYMTY/ax9acZNFgDWG3o9DPIZw3nG0kIZVEsoymDye+zAljKV8jiNoL9WL
CvdOUGUzkJ53EV22Fx1jo2o1mBsF+Ma2Al0Syhn6AuCRH4Ypq+Mv1PFvZW3F5aOi
W4J4S/FHJsFQpM7uaNaRKbcyvAzJPmdCKgY017P6H7VS4BR9wKznr8LxG/XsmX5+
WzdZiOt4djoc9tGFohluxb8cEbyM7vS0CDXS3epWKlF2N7wEhyjn/u/woETcy696
pKglLhWv54r4nrJm/GbVd7+h2DEi2Ael3Rf6LMCkpGK/sdn9GGylsJSGBB4lpVYq
+boz6xHh7153oJbnMY+VP5bINJQvd2xLnHIIgPZsTrN216JR9lNZr+ZnqQuFwQ4u
xrSjLZAot5OG6IECyFJvrlkEH9y3R7MMsvvFhiRJO8+xqHl9F901gsTM/TW+jZ1u
M8SXRHO1b9nnqkCjwrvq54N7pcGlkA5NZSVFiMjB+qTDyoXXV8yedLLS1901m3fW
pkxU0bXlgpD3PC/g+vX/2ZlBxvIuJ+ZjQ70itIma7rFsYT8vDsn4k8SvBgCw0WxC
pSFs7t9+LFdfu317zgUPgF1aJPARsbCRuWpLw0wyaBGNDaXVQGjTSWMSMSFklx/F
OzKgsk9tUtL1E/1svjP6jwl6sZtJwdIiYJlXtbfNiVm8hYqwHXYLdiQsN0eASp40
Q8PhhnGLOXb61UGW8uacJZz6RqCW2MSMALglr0SO5Nnr8Npqq9+kQU1fWmHdx/ME
/1Eb6b8gka0HtHwPwP2e2ViQRmBY7ejUnxhSJhfvEFmSNql8kKACAYlAVFTtuO02
i7GSeXqw7XUVCYIHcw5qXhPph0fFwoDz5LWAtr7hYjOttqgU7fudjqNK67pxyApR
PGsPUwXl5vn0gfzgD/FIMp+uxmivstCaJjYjC9i68lMji8EIbTzHgkjN5Bfdafxs
qPG1SckOk0BWXcvykcIYbIf3TJRhnEz/+xP85kxnGEszWqNMElSY4p5xboMWeuav
qG7q70Scw0vBM2oQTox0N1ckyJza7cMkWYXLvCojC+Gfpl4dveIfWHtJ8blKNPNf
ntYbbMp/aCQk8OO2g6vR5w2V1d79vVw3Ss7a3LuvDSDMTOpk1Iyu2kfriPGt0Odx
jsbv+poFE+bW2WtyiJDZJP0EwnEybiP6UXe/mBz1jaQ/ZQ/Jd0AhNnR+xphokUN1
GxmTw+GldNQj1smMWiZSYQW730CalGNw8ZpMUinwQm7F35dRkCYqFBj2mi2TkHl7
Ge70novHwZUNUzN4Y6sNRrKu7e2svf/AppUitrS7FU6O/CapYUDxUqVnipt5IKfF
Ws0SIwvcWQ15RlDtxRlt2xApSFm5hIqfW7Fh6T8x010YmozEiMacEakWkMTdI1C4
GfyI6YfT6lFQe6pJdBDOmI4u+mfcx1/0zosUCNGunVA6UjxIwGINr77snMtFJJnZ
aVt02RCpeHiHxPJRzdkSB3RLf1j0NBzzrchBsut8GtUZsnb+YfHbuImdvDG8qdAs
VLPtQocqNPmS73to6HU+DjZtHN1ZHvhR1F7UcC5zsURNVMQGcknaS6CI+DUUkDlN
ixMGJMTdYHNaJxumA6CaVOgXIqv/9SUNMdDOc7v6Fb7Iulc0AGCkc7VoSrA/XZsg
Oa4bb3IxgFFxIRsG1z/nonkkksKrWg7+fyW9nR5zQBfD4yY7gDyBa5h3lRE/20yu
ga+FSXfvlJRcor0fIbk7/a5JXOKaA6Nlx2TroyJnacuOt/B08OO2fEdArBzNnmwq
uNT0gRrf2sszfzJ62fTRdwse955mNBZ7t5sq+NBUeiMeAh7t3u4ayVBpXLLyEAat
NmeGbvDN8qM20JDOaCGY//yTOeh1VOzHoNXGtK+s+Zh8nDl0Y1YPlWANiizegdR5
KEihcMKPnRadzdbR4lo8y05dpfAtYo4gOJe9R83BZUrLVMHC5LitpjdgiEUCc2d2
BnTQhOEqQB574kocVESxtTg+N66Al3IRZEpU4dWj+/mrkRJMlsV5tnWDpSlUzdtM
T8K7KInJ7YRRed+NhZRKmyuKldzd/LYdoHdzYlHb6Tr78Dh0dvrTsSskANuteUQ6
FLAtaw5jHJS3ZQ4asURhZOOk+U3ZACF5qVizA44ZZ5SppbD/C0T8oQ8CIfmgESU2
gkKaob7M+qKdschMFftXudHpx6sO1Pd5ewSR7l/mMt3LiGs+7wqjTKZYI8+YF5cp
fuzG839vFVzyqkDJ/rYd97UZ9hrBzjiT7k3VXxqE8XHAzmJdAx/6V/4yNCBgRcpC
HJXvTVGyyWcgwVPUxc9xMuQ8CnGqQbGiy7gFjBSdTEdd6CABrRoKHPs1RPBtlmQS
oIBi19d36D81Eph5OX4RPT7IeqLV+wlgqHJRy9gXyOIcTnQV0RysXAUDLrjemMLa
roCWtORoTq9BpztcNWzXht97H75gCqzQE6BSKUjPESwa5DY4NZyD+bmsaAtjVtP4
RSL5H3NomBK7XE0+wTtN92qqG7X2xn7fPNZxOpv98DXFV7XBYvMCwKBKWgQnoA0H
QMDr0PVdvlD+4bfI39d2kxN14YqDOHRQjZHcH6yO9mDmCk1INsyoix+DminVL0DX
n+ukscG+BP55nZtLEmHnz2D+Wal+qSDd7k+pFxjejMYhB7LVzZ8HQpTlb9hy7Lh0
use1KRHaxF4cabY75RusqrjeaUmFOwS25YI5z36cIUOMEhziFAZPyBgI/4xpBCD5
TNMoxPmJeMck3CBJCxymleQuh3ILFZk7o3kf7nKSIGkKsacEkPKZaDaL69gKk1Ld
Z9h6TMVMV7nAuTAx0KhDQ0Fh7W+lFE/3q1cLJlkl9YUzdj9qXtYEhyEczu/CrLrr
foNI+6zC7p7uCDmNWv+R12Su9/T7F313/cd/sauIUSPAAmfRsbGybBoAu6Y2+rPm
pKtqaca5ZrSg6oTgxL2jLUD+CSvvjYZmj8MARW8fFpZda6lGCi4o5wVwFk7U8akM
hnbPeyqJicdaUkrbiVb4DWN6Wmjf5/xpNNRT0bJd6z2UMmz8ABmWI+WTybmuGcJY
H2qTj7n80/KXOck2VaOq9cLxeyI4cwz0xNf2c5wrbbSZcl9XsPD+MLPyV269dlwq
VQfIsDLJoHP+xo/Dq5L5NodWa32TUGOqcNC7WLvArpbgCJ0U3uP0YDACcd43HdV9
QLCmD9XY30hmdHT4CFk4VoZriJdXV8eJYRy34I792vt03i8K63vZXZwS0vV5Me06
p+r9FSpnfDmMokIuZ5oT9SW2rMu7XfY3aH3yvvMbbbszZcsM1ayj3sFOx7r1ov2U
NJEvQUBZD9GW3sRmHsiiCRZBHtkdIzOhHPLyRvxfmfZrrOz/KM3MbZGIpC3MDiqH
qG9N85DM5KbHtxe91La7vQVTZb9bxlTY0vEPW+WnCr/ybPNJ/vQbY6DVxnuoUJyA
LmQJzz9vkPhSXGzG/fr/feOS1wGJJGBWw7ZmR3ODvQKY8ENc4zfvY/4nuskHnE5c
FC5N2MEbM2qsX1FOen4H8Dt6YZkedqzkgpCuEP/wTo+O+BUpDw7xUJIO8I29VFgS
xw7OZYkIpJlz0uyA08btEPAv5K9lHZmd5I9jI8K/1gKoUncpWdp1Q9P3ys3QvxC8
g+NzaWlg94A4abEb7tPq7xyjNkUJ2NfhjsSmzTLq1B+w9WemcjX1xhAaJgAlnLTQ
28aHLqPWKfu/JQANY6WWavovAB22kvitNiuyDKrw0LDDHoZ40rsYwBjhWB6H2R/a
CBp65X2liZjxX2WQYo1+Wmt8ygo9WJjZ8Ayk1VwsVRxqCXO2umrMJxZ3YWp+x9dP
vij+eiKvWQUiEkaMmaH+oVkPZA42tzImvCp76MUdbuZQpFH8/oeDtNwGmMx7iuC3
vtOtjoISNeJxKJV+sPlFHqpY80l6C88QDXNhgDV9Vx3RGC0TQyfv/LqBqo1F4LVx
Kj7a2xeTYL5YGpIU7R9b/p5JwEX05mU/MV2qWTYEkQKHJNU9vjuiQkz4s67XLYd5
ryu89wiYopgglfo0drx8zy4z5Er0axESbgE3pSCIad1vQ1T+jszk5GgE6zeAzpfv
RSITnBoZ6JKLWVV5MtTs+bxAUQn6NA9L1bE/iDxZrVTaLbVvYG5xHTpMJGIWdq6b
127U+PEohjMEFf0OulweN+ncLUTnE+7ksO8T2Y4uOccZ3zWJdkT0vBnxDI+rTuL+
IARmjDKVkn9O85QPbkKNIFQZPT8PZpBe/wgTJTeRJgBYNlCK4cPYwXC9Vdh/LIjA
1FA5NWnLji5yaDi2TfscCOoHUVTEYh3IXtsivGobB8B3Lqk6QNAVQSRPWotaKm7U
AC6gi/fGIrt6hN16l/lp0CDiEnXkKKeN9ixq3fvZWaSRt3zx46mOD3Ddo/RWbtyK
IVZxN/19Eklnc0SqDn+hiORgAp1wt+2KStqWnjFhiAfR6J+22Q2u6U1OwtEO7yni
OsePMNCFTVOldW4dG4BtD0N8L84VE0eTaZGrC2/aZC45LVcPUjX/BtTA0T6yyteD
z18uOVF7Uu5KVsZfmHisMMBpM0UN9+dArw4HMzb0eWgk66yY2jX4iNnWgqDCJZrW
E1GxK/u8yDnS6KUCp/wDc8zXRfPUSk7s/r8FEQSs6Y7jUWUqdZj9rwoeRgGo4hvX
Soq1csJwo9J5Gvg+yucliXKAzKhApKrOT+fuBOqREop9sy1advufT2Sc4LmbRTCi
VIbojSZ/79vyIxu2hUlb4LVg7H+PaK9yk1uTKbYximEvpCmbjgJtwW0lyZb/7u7O
VvsueDDAV08YPoIBq0nHcH1m9T7HuJ8gNxHuyicuE21RoQIVYTxoAEJ276gaoU4Q
OpPnHi8RA3y2nd4rW9GytMVsCfKKiBWCUpQ963QT6dvhhdX62YgjdaB2DwJtzxC7
cqGgU1QtDyQexVvHlD9Y274EPeXXKIuShETDOzsYt7WtwTZP0jRX3tMXqdKQ/7dX
BgA1mWInwD9d0PLGPGcU8UBpz3YaLBEMcNqMCSAGr50bCWblGOasFYMCZmxVRUXF
IkCB7NFe47AOZ4iURK6eOsuYRZ9Xj+90oTwrI9nsDBQ+eMTkHtiln4Pmd3K2nnLj
48sH/tOAw7v7er7vFezfhv83EBAcFVXWgUMHnOWcc6HLcWra79PcTla3RA6LRtoN
U3yFi0xA37gBubnZu5yD7H2qfv9T9gy5yh7UcQwPnPoc0Kyaa3wVKpf3GB1G2eva
UD3X+qxhJa5pzgIg1w/7mUYaUJ24kl9iseG84+0WwVypVZhgefjwdtewx8r+OmY4
2Y0YYvdjTGGGlqWGeu/EH9fW03pA6z3jSK8hF6/eW+aDWMcVxDfhEu0qfgIgJMu6
w9M9QU+q4sMqnREghEHLQ52EAg5IYe4J2gX6+nY4uE0h5vTcINXnS/s6vEg0sNfB
lUGIZla3P0DpdOO6j7N/w3b204HIC8Xxl0cNg6r6HtJrKnjJvhj+gnrd+gQUD2HD
pM509dxdHA0zEJ4Hrv/nl2cKEgGZhzmqcP0smObFFr9VmarF+BxaAjjTJW7CmPxm
HspZQX65ds8BzQpsuhp4YrsNY0s1tO07W28JcV6Bksn+ODvWer4jQUP5LUS2lQTa
fwWzXbeZuEuR5GFxQciC4LtDhnFG4aGQvmDvdUPDqNebZ7ToCGjvsB6AdTgJ+EB7
RE8yWtvDGW+TZkTNsydbu94Xu+rrCziva0g32utOL0uwMgTQk1G4iHG8iJ2OZQ53
Vcp2+y5vsrWre8N2Vo6bkI+JPueUr/Pn2I7fZ6pWDpbR6WFUp2dFdV7Y4zi0eVXZ
awG0w/mBsZuWMDAbdCtgEjI0TCGzWEQGVrAQLCUdNRqx9ggT611K6q+vjgz99k1/
YbSwvP5Ag9YuggQeh1C/6Fhvx6Mt+7AV2dEMWoxAVB4xIYDMTGkJqvcqOXPrtTna
eI4cQPFJ//hPCwESU+wj2a9cwko/sYx4Jp0+3jsdEBZx0KvNphR1U38AcWpUKuRz
4LtLqvnXSkeOd5VFXHXYeBEAvXSkq0m+pQyppmbji/PLv51O5qXPtDqvoKS/P9qN
Jp/ab1lxws9bpKF/Zw+J0HxdGxXaJ6EvD870IC95MN+Frrar3tII7sxeI8LOHOPS
1h7+ebscx7De17VJapDId/qGAflNGr8E7eyN79CuiZWGUhcgyy4tLOZW2B+kcMoV
Nx5kKDOWfwt4YGN6Jp652mv47PQjc7OHkiDawYA0FSytnUSkxHs5182Uh/ZxV2+w
IAs5k87EQxA1uuaO7RTtx63+IIb+HljmMOXdAxeIIVAZMbGxKYc6x2hEs9e4ILO3
fSqyMc0aIDgMPLson73Qnx3VnMLJq4ZSUXVcS8drUkyh39ZCYN++zNtD6V/70gxL
8ncS6u1KMVqN/F75OKglZe4vgw00TSJREbESVv1W5YfOhOnie9PUG53C7gA1CNrB
S/doftHZ78XfupvhnaI8O/OnS7TsKVhR7lZQEMgAhfL4UiDMHkaVvxqv0sGt5emh
7RecWJmI5CZHn5+QRc4OPUBbEJNSeiL9Lyu9fUBb+MFUgI2Mb6haAq5xNxTUm7H3
NqgJoeMqbSfbNAYUo13cYMOFST2Nom5OP4zcLbRRYSAjU9z60qMA8rvkZtmpPors
KD/gzwsyPOZVfF8dV596HKxG0UE5hAGjCYFp5s2Njj6KOCCQJ4JP1KErnI6kczdT
VJVyK9B6+DelFlAmLkh/Uo4/AR/30U61lpJhrbIPE+AUwezJ5H438/0vIj5I1ZIF
IrmroMPLdhSnq3tqdbn5jQFd9rCfgiD6aBaWZ6+xhNZ/QNaD8hxsT5RMPF5BKQRq
1g3LlKBBTuyYpBnHFDrXwFsF/P7Z9VvUeFCQg2JP79gmFokEWFIDDMAs/UZu537C
gqW9CVqTTTLNJX129e7OK9doqUvH2U++hL4pUbhm2ObRznPAlA8j64wE3B0RpXEG
nTyyewwGuhyTbBD4Xat0zwjKhaNsStnaUE2QbKYLGoEzWHa9husk7Banxss7BMsg
Ox5Xc6c55tO37aSQSn+eZ753D23NlqX4rn8CtTgiBKU/tg2jTaTLv248Vd8JSGrY
WNcu6WwRud5ZHAMx3g6MdjEwxxEYepk+wa8q8YeinKRy1bWTSV5cXbwSf95ORRCK
k5pjFaPTgfD7cDNj1GWDh4SKWPuTUhf64xyCAHTvfxwD/l0uox7KWK/qFq2JGDXr
C2vjWaoJBc6ugtG6bZA6po+UHRYfME1Tc1YL6L6ZT+kYp98MphOAoSzx6v5Fd3qy
8fC0RNnW1XAffpAquNLIOuptIgIlVKC/tMIMHs/cOIZGtpF+ytc6ZxBNiUQ7t0ef
vLCpeXEiZy4MCfTqxisQ1U9yJ90FOBsvoZUKryfTQhUXF+E3oQMXg60nvRg6BcyT
DquGz76USy8679QDWnTd26lKFeKVNy9ikJ5qMf66kT8FPLhR3J+IdVT2X5mCAedN
RUZ1i0XavPP+Xg48tPf5BQsxXXg6rpZ2oQjj5izlFgpE8kKHHdFyfPxBx7cwxZe7
KiLb3PftULTD/3Dhi8HbrFubM4JMUMXi7EeDrp94kLWclCK8e/xpMf+pJVyEyvQj
XYl3Eqo2PRNmdVx3Y+4aN4eXlDuCXzblNQxcSjWKfUHEZwG8OU5ADvW96LR9h5ak
086q9iFhzN38zt984N/+4PrXDtMDqrb1Y7g1bKL+K0aQ/LHqtrYNGxpbXMPJZyus
wJtGMzBKsc9M1Jo34kVfYERHVxgpMYEiM38wdmacSsySKINk/LBj+QXz7960cbQJ

//pragma protect end_data_block
//pragma protect digest_block
7FWLJXwgsKbJxqhsQtLIbhAeaDc=
//pragma protect end_digest_block
//pragma protect end_protected

`endif

