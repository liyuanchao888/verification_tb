
`ifndef GUARD_SVT_AXI_MASTER_MONITOR_COMMON_SV
`define GUARD_SVT_AXI_MASTER_MONITOR_COMMON_SV

typedef class svt_axi_port_monitor_common;

/** @cond PRIVATE */
`ifndef SVT_AXI_DISABLE_DEBUG_PORTS
class svt_axi_master_monitor_common extends
svt_axi_port_monitor_common#(virtual `SVT_AXI_MASTER_IF.svt_axi_monitor_modport,
                             virtual `SVT_AXI_MASTER_IF.svt_axi_debug_modport);
`else
class svt_axi_master_monitor_common extends
svt_axi_port_monitor_common#(virtual `SVT_AXI_MASTER_IF.svt_axi_monitor_modport);
`endif

  /** The transaction corresponding to the last cdvalid assertion */
  protected svt_axi_snoop_transaction xact_of_curr_snoop_data_beat;

  /** Internal queue of snoop transactions where snoop data is received before response.
    * Items are popped out as and when corresponding response is received 
    */
  protected svt_axi_snoop_transaction outstanding_snoop_data_before_resp_xacts[$];
  
  /** Snoop Transaction */
  svt_axi_snoop_transaction global_parity_xact;

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter);
`else
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_xactor xactor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ACE RELATED METHODS
  /** 
    * Adds the snoop transaction to the internal queue. 
    */
  extern virtual task add_to_snoop_active(svt_axi_snoop_transaction xact);

  /** 
    * Removes snoop transaction xact from the internal queue. 
    */
  extern virtual task remove_from_snoop_active(svt_axi_snoop_transaction xact);

  /** Receives snoop address */
  extern virtual task receive_snoop_addr(svt_axi_snoop_transaction xact);
  static int dvm_sync_count[];

  /** Receives snoop data */
  extern virtual task receive_snoop_data(svt_axi_snoop_transaction xact);

  /** Receives snoop response */
  extern virtual task receive_snoop_resp(svt_axi_snoop_transaction xact);

  extern virtual task process_snoop_addr_channel(ref int acvalid_to_acready_delay,
                                         output svt_axi_snoop_transaction curr_snp_addr_xact);

  extern virtual task process_snoop_resp_channel(ref int crvalid_to_crready_delay,
                                         output svt_axi_snoop_transaction curr_snp_resp_xact);

  extern virtual task process_snoop_data_channel(ref int cdvalid_to_cdready_delay,
                                                                         input svt_axi_snoop_transaction curr_snp_resp_xact,
                                         output svt_axi_snoop_transaction curr_snp_data_xact);

  /** Waits until cdvalid corresponding to snoop xact is received */
  extern virtual task wait_for_cdvalid(svt_axi_snoop_transaction xact);
  
  /** Waits for the crresp of a snoop transaction */ 
  extern virtual task wait_for_crresp(svt_axi_snoop_transaction xact);
  
  /** Waits for the cddata of a snoop transaction */ 
  extern virtual task wait_for_cddata(svt_axi_snoop_transaction xact);
  
  /** Waits until crvalid corresponding to snoop xact is received */
  extern virtual task wait_for_crvalid(svt_axi_snoop_transaction xact);

  /** Waits for rack assertion. Times out based on the rack timeout */
  extern virtual task wait_for_rack(svt_axi_transaction xact);
  
  /** Waits for wack assertion. Times out based on the wack timeout */
  extern virtual task wait_for_wack(svt_axi_transaction xact);

  /** Waits for acready assertion. Times out based on the acvalid-acready timeout */
  extern virtual task wait_for_acready(svt_axi_snoop_transaction xact);
  
  /** Waits for crready assertion. Times out based on the crvalid-crready timeout */
  extern virtual task wait_for_crready(svt_axi_snoop_transaction xact);
  
  /** Waits for cdready assertion. Times out based on the cdvalid-cdready timeout */
  extern virtual task wait_for_cdready(svt_axi_snoop_transaction xact);

  /** Checks if there is a snoop to the same cache line addressed by xact */
  extern virtual function svt_axi_snoop_transaction check_snoop_to_same_cache_line(svt_axi_transaction xact, output bit is_snoop_to_same_cache_line);

  /** Checks if there is a resp to the same cache line addressed by xact */
  extern virtual function svt_axi_transaction check_resp_to_same_cache_line(svt_axi_snoop_transaction xact, output bit is_resp_to_same_cache_line);

  /** When a snoop response is received, checks if a writeevict to same cacheline, or a transaction with AWUNIQUE asserted
    * is in progress
    */
  extern function void check_writeevict_awunique_during_snoop(svt_axi_snoop_transaction xact, output svt_axi_transaction xact_to_same_cache_line, 
                                                     output bit is_writeevict_during_snoop, output bit is_awunique_asserted_during_snoop);
  
  /** Reports end-of-simulation summary report, checks etc */
  extern virtual function void report();

  /** Triggers events for snoop processing based on sampled signals */
  extern virtual task trigger_snoop_events(svt_axi_snoop_transaction curr_snp_addr_xact,
                                           svt_axi_snoop_transaction curr_snp_resp_xact,
                                           svt_axi_snoop_transaction curr_snp_data_xact);

  /** Waits for active threads working on snoop transctions to terminate */
  `ifndef INCA
  extern virtual task wait_for_active_snoop_threads_to_terminate();
  `endif

  /** Processes reset for ACE related transactions */
  extern virtual task process_ace_reset();
  
  /** task to sample parity check signals and calculate respective signal parity values for parity check comparision */
  extern virtual task sample_and_check_parity_check_signal();

  /** Sample ACE read address channel signals */
  extern virtual task sample_ace_read_addr_chan_signals(
                                ref logic [`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                ref logic [`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
                                ref logic [`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain
                      );

  /** Sample ACE write address channel signals */
  extern virtual task sample_ace_write_addr_chan_signals(
                                ref logic [`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop,
                                ref logic [`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar,
                                ref logic [`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_awdomain,
`ifdef SVT_ACE5_ENABLE
                                ref logic[`SVT_AXI_STASH_NID_WIDTH-1:0]observed_stash_nid,
                                ref logic[`SVT_AXI_STASH_LPID_WIDTH-1:0]observed_stash_lpid,
                                ref logic observed_stash_nid_valid,
                                ref logic observed_stash_lpid_valid,
`endif
                                ref logic observed_awunique
                      );

  /** Samples rack */
  extern virtual task sample_rack(ref logic observed_rack);

  /** Samples wack */
  extern virtual task sample_wack(ref logic observed_wack);

  extern task process_cdvalid(svt_axi_snoop_transaction xact, logic[`SVT_AXI_ACE_SNOOP_DATA_WIDTH-1:0] observed_cddata); 

  extern task process_cdready(svt_axi_snoop_transaction xact);
endclass
/** @endcond */

`protected
eXYbId9YDdGb53M/COfK+[A>W>GY4.14d02/-A5<X7bH,,&JK@.=&)eV)GKUV)=-
Jfd@J6]Z1(9?[,[H:-16UNLcfcEOcN(?P@1HU[fAM]6d6c)T53_&<[,>RKfUZ#O8
Ic9d52MH+9Na/5-=(]JEM;=3O=Y/)@Kf>(c(E8(?0gK>2(QQLBU24QN[Y^UHgTDD
]Y20W;2YCc+_.,DaV=@8\V2]QZ<@/83OZ?e.b5TH&8=P<(8J6f48bU9f&/aSH)-I
>>5VebJ]bOP(L+SLM-RK4SE]B^FF&a_dGG,6M>7^Nd6YCA4GP3GWJ/;-;Nbb[PNG
[;L+^.\;C].fV/+Og_WW,d7c@6&IV4G9_ee@T&b_ZY^e?U>,<4>T)X6&ME/,\Z>R
fP(&]/&2DTafU@R,=f_PDGL3F065OPOV2UI>E9MI.#D0^L,YXD1\S9XW:>.-@Z;3
85a_688?]9-8#aVH1434X2_Md1cME^RG[WA(9/-3/C4]<8WXM;g4T-PPgW[9_dbH
DK#AC0:ST4Bg8@\gD?Tg0]S]CaVdUceQ3-U3CZ,GbIc;BWcJc<)f\S[V[[5NL>^6
=AgU.La/B(&bA08I:I[?8Vd-TH10TZ^eK>:+B_2BCDL4IG4IWU.>/&OND(RHEI1M
Og(c,@Va90d3AK>5CP>E^]G=9I_TKe9IR,KHCD[Q(RB2QdUgd@81,NB@W#W>_4Z)
V=ZaY\40^(94#1P/WA+2KR0N3^(LD7cWUIFMLI)_<NN7^cf6FAZ9SRN0F&(NTYc^
N\-=/CAA]B8bNY9O2LMZF,?a1AROV,]2_R>C(0\0QcfZ\T=LV,<Qc&ACL:cM#YgX
VTf8E=N)dSH11-DE^ag[R+UXI<dc@S#,:c-1G?2fY[Ng?_PKFND>Q,FOFKI<8&KP
;.#K0KQFfIV,+ECXAb)73#ccJJc&gPc3(1bMB?W9aYd;N_6OgDe[V2;C7R,H^V9g
_@2U>-6-2)U\2-[b[,:HM<_KW@a.D7/5Xa/8bge)(@CC4MD.)JeBWV>4H0E\@VBF
/G9be/b7Cf,NR+<LM?89K)b.bUb992?<S^.6##deTXR)<,3RGG/b,N^9NSA<5]^0
C;7+XN.ED<7UZJZ_89Ia/7/cJH(Z5EB(UGN,)^5.Zgg5cN3U(0N<5e9:b1(>F00+
ULHUUI=)\3cdDU\2Y/=X<;C+GQ&PFH?&QPIX_b^0M]1,)@VMAaXG>)[DUO3SV611
,FIKPX04YP+R:E[31f,88Hf>LXb<#=F=[3U,bYI7O;CgQ#LKK\?cFf1EUR-Jb(7Q
?POR[c8,Z\6Da9g(:cbEK_OS,><RS@S;AMDTf8&NeCRL0N\NM#7c]c1&ICUSMN/9
3N\&,e99HVbF8bYf^A[[-UXD^#@>I1?#ee8?9&:.Z\GY9-@C>S]2F>=M^J;),_=0
++XF:-1U#SO_FL,RVD]]@Bg843A:afcMPVY?cL/[KPe/3G\ff:L,G^76??B1K?S<
e@cX2:5X@3_2A\KMX-(Pe.dQ3N&T-b195T);LeHb_U90\aLQOKJ^_/AHO6..EJ#&
g87O8NL/c>W#XbUG:4TE0M=CKK[:34@0U=fT/2)83e2EXbI:7^E-QM&Qf&R>9dW7
6+[LPL06UATHbfV_(:ERbIY)dC(JYTG2KMSe;W?(aN]eg7K+BaDK_33;4X4J4BgA
9.B./N)Z:#)1W?E6#/Y+52)9Ie.#6L#B,)_1U=TV#QM>8,J8,/#.;=-73TcEFQgg
WF_e+M=BR#Vd81GZ:1bF&N9-UE(/bYTE\&(BEO[SeAHSH#7[AVYdRN?(\b0V]#?^
Sd<I?@2JY[.40^I87;=)TO6dB+B\c&^N3S-@#1_NL#dcDZMM<LgCMB8#.NG:^LRU
R[A8^2fA?C+84K=Q^SVL4U/+L8Q\@31FH^#7\8]7IQR,LOX051JLKWY#][CgT4QI
V;KE#[\LOfSCANNFg.3X-_=N9F1OOY+=e6da-SKc>,ZAI91&G,XM?5T_4<.[;-50
8-/^)PQIT9GWf_8_dL6Wd9[YAU=d9D8&_RgK:R.2:ZP_aSI1)DUX0L0G=@g@WI=(
^T=a:^1=D)=<=bGbb4&+\EUa5>S[-,X,-KY/I4gCa1HC7fgDMbFXX(HM9FK[<I:Z
>B](^WAfRMIM3Z-c0ObDeX[>MH7CA#EY@Q2KW(F)I;:3CFRJ_&(5C(BZ_QBg+U<_
1fG8@^\I4XK+)QU.b&b6g:YUB.Z(LZRA0c+)f)-e[N08b/T3XdV8M7:H:@Ue/TT&
L#/W\7B_>_8>&b;V4LTW_Jd-3MQSM;C,cG).Tb1>Z,H(=X,V]+GHbXY(0T;-d05)
QYZgS;W1&O/bgY>[ASe>5DgJT,B66aE.IK3aA,G1<H-F?-P27VE=NT?5+Df,(VJS
+f.(;6ZPX9HP0OJ0MW-PJ4H6HQb\Q;>,0QE2:Zbg,fTH_WMCF,9gOS1TMRMP].Y7
EL[b4(3gW4IO0R^Z@Z(7C/(0\9CY=\g7#]<]:?7G@SF52_C&_:Z_@APe>9XdMI[a
8OYY[3]D-[A46Y.(0;IbHFb82LZ,>9W1[PLOZOaC]U<ac_]Vea3&P&(BV=W[XGSQ
\aB)^EE&#Z-BbKA2R=_W1#c]Qe^F@/52fM).6T12V49HX1\40N;,W1,LN8^Z:891
J\IGAa8U(-=,(Z()EN\2;WLM/a5X=9^)V(CJ&1#8/.#V8KKL9gOU+O;.WeM53C+g
W/Uf5-GggPBb:]+Y:T+&>Q7Z>LgBUCHXJL6dROVJ-U@IY7dRN\ASF=/<ZSd8N,)&
&1]MeDVQ8S[4:_HZeA<ECAI1+N^Vf9=ZLR7/#&B4T<#]FJ@0.KDYWe])g5</VQ=U
^FbD&13.D;QO7b2L5^H<PC2H;YB0)+-&Kg5^L\@ZX8C@DC^GNbP3E:#LVVC7W8K@
)=&ZF?>(XF/PI+8\VI#&C>g0B9/VD8eT/XOP#0fX0N3N9P1J56M;d1)P+_\IJ4FW
4S2L>L;W/>XE(eLVS8?0[dY4/S?ZK:)3>Y5LFF<Cg;T5]ZHRa<4#X,bP;;428)bL
4]7YN;B2=+6,VP.0bKJF423;1A+?QXc:BI/R^2CA0C([.?314EebeHb.?cc+42\=
J:FW;PT;J/+AagU3(-Oe-5M2^81JE5LV85@NCEIfb2K#8H96=_#4TX384fQ-(LCU
D98]DBB5XXUYAdd?QI5URKBEE0\Y-?H;(;4KfDT6b^3:JC@JdbL0P&O7A[0=4NOE
+a>\#D)8?]GSW+WPF\N?MeIA>V2^GXQ4eB4e97<?H7b>(NF(7,[5E6:Ac\EY2ZCW
@55D=,&N;(97UZ&Z6dBBcd#a;,G;+J9MUPY/;._>IQ48OJg-Sc_S)US;2eFQFfc4
0U=3Ra_aV3W)DF?;^)1g4/VV;W0dN:D_\R(<HAM@3FB1c(C(Md(?E@NPZR^R?3A0
(gX9JFO[-L][8^Z;@#BUg/P]P=K0)33G\#aMH8.#\>N(2A]UYGY(]_IU^/,9OQ+M
WM&37G0TRC.2@R.)>TRM6FK__\NN5^,UY1VF:RC38gBcQ5L;5.VFL&aNEg>=CPNC
Y:Nf43D38baFdMC9ENfZPX+GDa]b\)-L+MWVQ^=H)2W[K,Hd\>P0T@O@AS(e>_/1
QGbf6Z>[?YF5<5bdFCH&PC6M,2DL\3d-\&W:G<6bc#=D4A&^/GaCOK\X,HWEMaBO
O8D^ETI,^JMHV>W(-dX=2+(^J0e^Z#d#-d42/E)C-A(-^H\6F^(LOQZ325HUc#ZQ
f@R#W2;M(;DDX3C1U1L@GX+-#g,If^._b^c80(B97;5RBG@M=UI[Ob[?OD8dNXDg
;(;3AeW2BUCBfb:E6gVFK_;-fF-NGXT^_A[\VcEU.YXCOU\\>8@WU.Z<L4IFcU3;
/5aX?]6Jab<#UeS5_Q8WF^,#Xb7P@:9M>e8&d40W.aW5P3++)V->44=b]4KDVe76
X]eH;<,#N557F.;]0K_EHLZ7:V<@LN2QS:IB=GCUW,K@E59U.&3,//W)C74JFM.a
1\&MZf)f&>S:>^&4JJ4VX13G7&DS;7856#V.S08__QG8.?)CP^MOJM0B2FRR4-dY
4MP&Q^J4YI459S[4FREGJ,@[c;V<N2,5#_UD#K2d&X>+<&]4eJXR2LK.EIDZ<1Y+
TQ5ZfC,)eVTdXU]V1_MdDFUEL8YG(A](^#LJ5JJHH,35[#gM/a+EQO_ffV^^2<<B
L]D2_.C3R8ab:^)fDWGM)FELBZQ)E#O\\=LCL(c9KL(TMD3.a.]SRa)RPT8^C-/-
K?6ZEQ4X>Y-T?]XC+OQI6NZ__2X<<TdgI7?_5&VK6c2EGEdU<<e(>M4:/Z8DI->_
]dae1Q_;Y)G.dKACODT:K-A8P0_=4&TA>(2LERG=dJC?F<T-^B@ATE&_;\gV8U_g
IMc@2@f14:d\HB4SW?K_/Da1;RN9P>@C?fXL5\=d[:A&e#&672&APG\MPaWNA),-
&^OB/S>1\cEVM4820aDR3(FDS_;bXDCe&2WJeT;\e&CNbF)0Q;S-Y0(9>NY\SQ[3
c-NV?CM7b:ZA8CF/:.ZY4+OM6aIbe<DSDf@d]^+/Oce/.:N[L4RN;[LWR#eT2N)4
g:N=#@J1ZBM3+;7d:[851#BJAeW^CI&4<I>>KA2/HG3c8E\,(R7K\.).H+#SIT&;
K96N@F/&1C=_2_BT?70E<T,H7:M?YZV6SYQ90A.+G8GBC2B_faZLF[/N0<1D-<[[
aaE8e2Y)2DT,TY]FKY2N15@KRJV_OASX9(F\<PHWX:HN-?^O(L2Y;7JCU&J_e);P
SeP-=KcEf.LbI8M8FV)07#XV?OM(Dg7<L\9Sb+L(1U81gfDcNQ1AcLMHUa-9:;)1
CNLOMY&IOE,e>3S^?]CcgS6UD&JZP(J;@?eOcgea>g]Sd;M+@f[F[ZFQQ1MFE_R)
(>]A]8K?c;ecQNaaUE1bX@YR=,FJU^AVd#Y<E3<aRSP^/F++/g?N)NdYF-e]KD&X
YFS5_4;b)JQgNI7076:6)Eef]85W;8OKW/g/V+a,WbQ#N1&/-[IZdc<_RQZB_e;I
>O8Yf;KP13LG<3P]WP=&(J)+U4&H:ZR:+gWDFSGL7T96V5XbH[=0;RI16If5Re^D
_:bP7bYEE,->?;EQ#QOZP=ZE2<\([5gJa=N_):WTEK#A@<KX1/50]B>UA>QO<fV,
ADI1;(G/eBZHJP3@((XPY5RPe<T2ZH0,U#5U(\M1cBE;=I_-Fc-(g)RfUFEBJPL#
aEV-^d<3>)-c=VDd>B5KQJE.+b]d=_I>FU=TRAAVYaT94R._/7Rfc41G;WCdcI=_
I:92-4d3.>4>H0.RJ2T\f1_0E8ZDc.>X5W)YNH=-J.WPQ6V82XJ99\N/VGK3)6G3
c;6NP)TZ[TI\MHDJ@IJ6/1T:)&TZ1eXI;9:29TG2EC&/AS8D?H^/:Q^RP_7&HUU(
?-6)P1IB<1ZgG:GS6TdW>T[(B<=8_>._^KN^TBX(1+OYKLb/F)AF_5M0,#-VIf3I
P>=H[g8U4A7DBF^B1UBcPKM4gVKR/IaaK9KS>BN_KV?B=f=)J,S4]7c4]0J4\B7@
:^DGB2G3XX)[:fFCW)]c:QgWWc0R[AdSV3ZIL4B,O6fW9Y<UOPEKI=MLgRcfUP(2
d#,&H/0VB#D@GQ[S^Mc+_/\O.;1Lg\5/S+UJW0QEM/Cd?EI363,OO.[N)ED8Gf.U
>+1=_(+M6YRRg/<>8]:-U4R[[[NRR7MQQ-Y0RQMM8HA7S)):5bbb1):<E18/@)7b
>W6H-CV7>VBNXE&MAeZfGXLaS-])]0/8^N,AL#f9JQ&-+MV&I-VQ+Wd<_APO+9ZG
?XZND@282X1)93ZK=O__c/3FVU)\O9G]?[E43F=F)-(0\YL9:&#WB:#5SOU+.3:W
N?e1.]:WO6-)_H+91,0:(6ba)MWE1)d+)=X4OB/V>.;?);eX:ALc9D-H2OSM@0d6
4?K\]CCT&HJL1c)K2_+SOdYL5TO2Rg5F:&/689?>f1\CQ-?25<RNa2MAFE\O(YR/
a.:4];Mf3WPb/cG;&F):\1ScJF5H:0:LL?^NJg3T2\A,TZ6\[gSL7g-N>dK\bA5,
)5-^DSW.V6Rd@IIf0;G=8/P.cMGV(^X/K_;6C(B1&F^6XLf^2YY?:>Z:AOa\e[JA
FZ>]IbRJL&3:<V:9Za^B7M9Y:G(RZ1=,A.<V0@46TY/49XF,5B3FIg=.P+1EY#(<
aS7L#2++(03+(]-RC,SE(5(76DAf;0:SQ#>PO_;Z5bVf&SeUf_U3Xef@(bD#;#=C
=I<,fHZ9684@FE+6=f-?.37LO/T00..02R^+2^J?R>SS[35TdD[3WT1FbQL5&:]&
U&EaBI0eZ.1>QdVV+0\4[R8>\fEU;2?A3NP+1E+2PR&+C4EMBe2eX;-FDd7-;B&f
W&^=8@\d/.)9\:P6RFKeA=\628.7RF9Z.5>Z;8GGRb,?.KR8^_^<BFZKVe3R\3Sb
;VM4U[]Q3g]Fa9?d.70P01MfG3GZ^AUb8(UcA;@dW->9@JXL>NVWU6ECG2C)1&>^
0?S0F@AM0]1/d=R>SbHd-ZfL6D8?H)IC,edUXB-9=F,b]E8<@/Q.?MXcR[2C[.M+
1]?A5@MQ/V9X/7gagCL2OR>-H\;E(9<N0+Xe.bg<ZBUb,2K@43EWU[>S0,X:)DCI
8-7Q#?C7<_&]f7Z:2=aCW/0I@>X\Sf((;N;G]5Q&O^3C=&W1BQ8/c5WHPBV]0JO^
7VK?(TR-QbDVI-[7SL;SgP.C_->5D<^E)-7()A(FVYC;==I\JJaB9BJGbX(NfLT[
V_cXWdcC:eAWd+2RFX=HYC7G;bgJ0TLb18TC8A40F>V-B9,:Y.LB>fNgV^UQ3#2K
84O5R@LPBb;S0:LHTOfH_ENW6+Q7J7EDLd5=7(.<99e9cF5<G@?&Ocgd&O\SN59_
^I6W4@&W)&.TWHa?DTP,@?8CJ5eDTZ7A:FG@89R5&6R+0=S>@M?2]3dN5_,4(O=O
B2B83?M?7]M6X/be0dZ#7>3+,)6O2c:4RV@)P?WXK-[P6ceFZ:gMI5X7BO20cgBg
MbX;1]HM4eBGC_;gE0LUYd@)5.8=JN=<,1(RB+ZM:.gb1S4@--RXD6R]Q]\O7,ZC
-;B<[0?\GRY=+U-ALY=^;AC(Q&LEIF@700.<9A[ce.feQ=5e74/:8FfXg-N6Q5S6
T5/?XW_I7.325AWNPFS54FSH5#GV=P(IFY6<WeHA@O/Vg]<=4/X9#U#0GHXDgg9B
P[N@bWAYc<8F(LFL\]76g+bDgK;@SR0E//Z1gOGc^3V4CA^]EZ7BGd9c=cZe6,Z)
&\@4/Rg1MWd[?bLBX=Pd-B7:A^=[[2]4=OF[P(ZY[8?.M]<1=@]4U?\c_D\C7Qb=
OVA#50YHH3\,b&-M1\,<8E,@S@e/OIb4O3I5NUJC&YMHI4;:+I7?B^.25Q)#@7V/
.V/LU79g=]-L6?YU1ggPA,d21J9:fV:Q>RIO02D3P@IaR?U/V6TI6FP70TT#c]NN
;:G(]-SG8\,IS6K,FHR<U?ea6-XHTDXa3V.5I/+[?HgHI)a/ICg/5Fg[FHa,GJ_e
MW9Bf0)2\3Ie2GM(eO&^a)L^G_G#[#HJFg9]1N@ZQc9&/UF:Q<UHUA5cB(NVF5N;
,aL=2-V>V,d(.Va^>>fH<KXC9IXC[VZ;,GK4.b9RWV82&LHK>+JbCQ_=cg47;7V6
<P2V7bGR9)Q6ZP52CA5@W81.6Ib6#fFD(SEc)IN0P^0bA#DFLgXVU>DU9/=Lg3Q^
</8HM,]EF4:BT\31/LE210c[1=I,B<ZW)5fVXc[<A2V9L-71:Y(P/a_cf[1,>:9Z
Bb&f^ABG^#gTZ[@[GAFW7[^a^+YK]BZ=8./^6.Z9),C[TVAP<-a5-Z42VWHPEH>F
./EJJ],8]U28LHQWVJ((3IRd6)1d3H;7_]#.YAQU?d/\cP^Wg9S,8S+66bL3c=3E
f>N9X?NVFJM0-g8B3PW@He&=CN85>,B@KPPWPgAEKQ,dJ8;:<+;C&(Z98bW\b5FO
2]><26bJX#OA9,WXKf)ef?+Lb\[R[aMGL84F(3@bE#+FYU=MFR#P.WW-AS3=Y/Da
9)VUMd53aK1eHR:J[OP9Z>&dSRV)8UI9<12XO\5_\6F)..]/4L8;&Pe\g^4X19#<
.-&>6(]c?T86HC87,48L.LV9G[&-<>1eaN7V(MAG&:Df_821L.8^)e4K^(&5.(W7
W94g<G([IEX#E#U7E34RU[aJ2A)^\7^aUd5YWE-OHeL=6S]aN4CL00I=\7)1,RG1
<7KdV6dK54H/.<e:>=P_dQa7V)W6IPT1NdM3_]>PIMcSHD^8R&,8/Ega;HZ[JI+L
0CB+\DO\L)+,8QaDB;TeV-TPZ9S1UA5X@[LKUFdH+V)&=?)]>Z>2R)>.94.)S(MC
@\2Tc9-P-#/I]&4\4YZ;a85[OXF,5CD,KY:HBT5NIB,gJaNS?_LFW7S,XBV1^A(-
e<R1ZR#VB3T4@V8&gEI^RE?&3CNAJgfE<JX3;IW/J=U[DSOQX0_0Q#UZN\G]1ZZ^
,#XWJ;WV3-^SO-4.N^DI=d&YQRV[F8I=O>^(#M]KB^R6)URH),L+D.<GRIKA0CFI
F4EP<EOdcKF(HX-0e?.e03bggdK(Q3:^VI7.9SGC+B#+FYW9Y/DVJ3+(Sg3/Gg5X
+50ILVNU5a#<ULNe]=NTK>YUU8#5N5:A2)YRN0D0.bd1Ma\/G14R(BdMgELM.gZ<
J>NQBTGKSB6>JT^YM;Q&Y1dK;5+RQ3PeWWcM.E;?gF+I=?VFTOW\QG-aCO:ADfOG
0,B,51XKK4;Oe_,,E6?03;Pd2eC1eaN9(A]9fC&Id9acCL,f[K152GKZ@B6LbI-D
=^98,D4#c,B^91PY9LHK/d,Y+;a,PSN@,?1#29FEecX(O\5.c.B1(K7d=:AV0Be[
W0>NA#Df2FS,-/78,H_c0+EB-BP[\FI::9Re/[EB>&:HNT9:M(<WX;=>WL-)0N7\
7]7bEag5G+A3U_(L&GVX=S2):Fg8^Jf1+_S@;^W<g>?@0&&5V/0RGeeG/>EOEB)6
U)?J?6=?-BXJgE^_IRePPc(N1=3Q.-S9HAF8>^>KE)719V3-a]:XcL#KDdDA0D93
G?^RI-]UX0X6c2G<V<RAYa_N77;\\WZ?.V)N)UVbW<T>I8LTEW7#:RH8T48)<c,B
,QPGVF<>SPX988)GOQ@G&FK<TEbG;X@_\VSS,1JU&6EZOUI2ZB1?gD-S)/BS7M@C
HX[P;9@:^E+)A,L<,;&^7<AeVQX7d<)HQ&9JeEDCN-(J1TOV\V<L?Te);GBW0=.@
_RA;f-P]Xfe7IGDU+JeA3\2Z#ZZX@\IJ6Xe70=T&;Cc.f+,Aef]Q/7M:_KFWKTF0
FI0T:WL@_e/:@M=L(01[[R5<O,;2]A_[MebgHW=a_+=:c2/QKU45Sgb[#V_Zc,CV
-HN0HXJ#M)gbBD\_cRNU_4c<:5C73f)@gP>8LdI]8Nf):e#F7#3<[@A/L#,e9L;I
;)33?]:2=4<(U>JQ?.a..C>XB2:2L=/-BAHD5H01YGP/L_D]<K4B&MfJ\.5#aP6R
WMV0>=\E#+5[AWAT]UUA.8VE-Jf;[bN=UK&@R6J5BK3L]ag@Sf1-[^>cK45B@L,=
Y6c;ZYL2Y^+VR<),4b6a&;>J7AXC)c>gE<7_]J.S]L/aDAJANfeUMgLac#O867IC
ed@3QDMYUA:58GFZJ6KN[Jd7efI_L#8JT6HUTQU4WELC1a4]XG<bJUDD0_;Qa.6L
<EA8(aaVcdF?&b#RM/\P5.Y>JZd-&Y1OeD9P&;[SSU5=?+9><V<1Cb8VPUa147/g
?+b[+6R<0IVU.7Q7PK33OI8#I3WU>eTW0)M[_[?\VUbdYW215+5)^[fG:+Y_B6KN
-Oce(BRD^>WMS2E:E)Y,DU4I[>LgBb#)[IA,_LY-IF(fN11@7,d6+[&=g5cWJHbW
0#0SJ1)[F)ZV+bcdH-0f52ME=3TWL5&MBTd+AH82A/EIYVBfc&WO+^O8I1&XZ;G3
G;;6b=RM^=Z@aAV9P1)gEL=3,D_YB,B/S0EU#b[:aTd]DbT]<G@^#/_0FDW4Mgdg
3E()N__e<]dL=,JRFgL58fOY8JBQ;>.4G(S[YIfH(Ac20-cMNAZZ?H\EZ00c\M8^
Be3NXQ3ET;_Z4])Nf2HOb]K7Ra9B(6J]</+Zcf_W^/S+/:I3I\9^9fG?9S+WQC>J
?9N@L51X+:4>_K0@Va<SQd[J>b2AH2C<1#c6QS##RQE?Yg2d?+4.#Hg[bKNR6)ET
B<@5Ga-.f10bTTR?(SK[TONV\L[IM4.\G_:JO3+IG7[Ba&YYHVG/WU]_B9dGP\@B
V@.221PFX3LIIZ@d[#XbW@@44JWE&C7)[e#bCO?EbHd9GXBQR]eF:[3g1_4>c;\#
,=[gDP@)I:1/JcQOQd]Z^X,;G3Sg^96?f.G<O-g814DO:)g#&S15ZBUR=&O)U>(@
T:/1cE/@=8eY6^I1PMedQeZERS?+J\0Ggc0/.-FC^UH?86R@fG[^B/L+(<X7;_DB
NC1<D[f+@=Z=A]^X]J.9O4Hd4Y,=1491gHD-W@UdAY(Y\;Af\f80-+E2?Jf)e:(&
V_7ESZL[-#fb[#&FT3+G/W^WVQ;H7cK5N&C,[AME[LO,;,3W.0GXK-f,aD3B&fOJ
e&c8D.AUgLLbNW+CBd2P2,>dTIbH]#7<@=;G[A4K2_J2ac&;.R0SYLea/Y=XT7d)
K_PaI=,6E#BB1G6QC2&<OF_+Ea>c<#gc,E+Gf^CY6N=-7<-]>TB/2LADIdEO#?1N
V2IJ6;NU=-UZQdC7\,4f_d6fV1f\PDH)M@ee;LEf9&\F<gE\P40]U4g3=#TCa.9D
Qf(T-R\(>MTMQH7J>U_H0.G#I)BF@[2Ue^DIPH:(^A+,2M;0(DbgYg&+>COLKTE?
ba1A_F)&:MC6FdZACM?WW9&RRa?)P@]dABRX,V]>f+\@,WJ9(YVC?EYggca3G=OT
2[KL8[:-Og..3IcO/8Rg#;#[9+YZ>=NRQB4@[4K>Y2Cc1XN?2251G:)dJF69,3[V
;(?I(U/.0-bAC[75P/@X/df2S6AdfOV(X#:7A-,ZL_]6JdPFJ)XO4f>1G[PWAV])
P/,PL^#XPFS/2=WOdU_)+C&07e7cf87V^J-(Xed@C[Y8)CD>H6bW^)VMfd6+H<PY
1QN?P://KOYN9.#V?,_BaCIg1GUd_0bZ)V1YgA0@G>Z;PQ56;0,Y3;C3#E3BE)K@
R?]3JK>K>RPN&JeP37HZO>gPA.W_JVF.Ce9@FZG&Y,0KE6X/GR;K&&8fbbT@?;b,
CP,L_=UG]6)JI=NMON^G4)WM#Z#G68=,F9@>M4H1]56H0+Z9M>-G<VK3GN&fNd.2
f.)Uc.[<=TWF.cg)49(>eI7E)=_GS=Y2K?#YE0^B?Y85N+5F3RL;\ZU=2S_5/Mcd
^:/A;=IC7@]@&G/8?56aNS?(HZ+Ze:=d/6J,:?(e.1Gg]Q+^2OV)e(P1&8b+?aN>
NVX^3C]&9N&7(]<IO<CBd<8FR_ZLERL9c,If:E.8A=98H6&.ZKO-KDLW?Z3b-1F]
7O.Y_NNZKMN0JA,>MJdW][_&AKP43V^W/0&V:_;7>b2DdRAdA(g\;+bI@[g;M7g,
&3(M-eS),WCgaXg.:+b@S;AMA\aL,V_=aD6HUAg2&2[5Fg_#9N6Y[-3G:&W/K:5Y
g>bad^\Ic/<Q_HS]^?/1D@FJ(M\:FL@18O+#:J-8b6D;9N0&W//^NQ1PTCO;&NeC
?WQOaN=L_.;VY3QD#^JJ8;Ha@)#c;a3W1+6EN?-25X8aI<;\ED6>KZc<L<637+>@
PLVAadB_1@+P5Y?](C2/UUGfcQA:YW/Tb;e=(SU,Z.A;>WPa5Z>Re#DT##O]X#&Y
bg=RSF2Y.7Fa&bJ4<K+AR0UgcMI?5_C;U(W?WLDF4-Bc)cPTKL#SFQJ6bBM7cXF0
,598/]TK_e+R?B/c+T7?:7@0R:AAGWF7)\=<T8MV<.8HJ7;-#89XMWE?+8;9]+fW
<WX.[X+aQW,c,(DM84T[QJ?53#1a\KefQCDc6MOTAX^ACHBUO&=7,SUM3)FMgL?f
MNIDTFB,4bI>GIE9C7+Ab)<NZf:-@d;YG1L,FT<gK9ZV_TbC1D<;M]E1>J,Z1eI[
HFWVLYX\,==WUUbWPO-@Jd)C&#R?UGMf90)(.WA8+10<6;SJ?FYFM83JO.@@@+A(
VH\Z)UJXMEOLQQ2Ff=_B?gdT^0bLb/-PNObDbfKL]&-FCB/d^:1:8_Mg3+[5]^C8
.:Oceb34Xg\cY-8d1D5>)XE8Q]^2#-M]G3EI#LaKDLS8J&TSSMW4P_B<S5UYNaIS
&T-?,:G-MBQSV-E_aQaSX=D22EG4DXaI4YDSJJ_a-5<b-+CgPDD5#+U2gB#].\c\
XD.5#;/8gGNTgYB&cXY@L&e;61^ECJ:89^C.;CcZ77;VF-F-KTd]TeQLJTYHA4/F
IDIWO5_K.g-;ZWD52NBPF]5TD8&.<PI3(Be-F\ABHdeX@KaNNdeA_,a:&@^K6bRJ
LGF-]eZ1VKCbK67>S7:1?_#?>F9;dIH5+Y602JV-J0:Y>WBdJg2NWK_A91P42V?\
Qg&C^-beg->K1_cC,Hg7ec>R0OO/f1A6D/U[>PTS<XDb)X4>RgAR-gd4B/D[(>c^
Eg-@T()Tg8f#@+.>[\?RA6<8Q_&cCK6@\N-=NDNUYA]3>O6\YSC4/eT_#2):.-<-
ZMLEURP&@XYXd.PWd3DF)gO36SW0/Nd?HU[60KHH00UL\=@X5_&PKBfR>?Hf4BD)
]<2/A]\@<#2PSDTd==OE)M;g>Z7,gV)-@-B-X52Xg8N8LQ@,P]DG^O-E&3X,,462
8gB)YI)H+:;H06M]NF?AT4gBCRMHaP7,Y)91[:F/6XKLQ>]E4?WK?>&AYe<H9.B,
\6gcgPBZg-AbS_MRd_O#9ZFY)a6]F3.B^C;_LbBSBZc,E6J30XWRc++NK,T&Ob+2
U/AgVER)ZGf_5NM8R8=7IT:Y=@Q_#1,g7ALPXIAg-7IU)G7TZWGY;)80TO0f9VJZ
PEY^<d4C(OQKd@PI40#E.fOM]FGMU]_.\Eg<A;ee]dTEI;E5L7Z@GK^=cRL^?OBH
_WQ2/d,_gH7IA3(7)Y^-A8F0]QX5e69RLJ,.&OA8e4[^VK3+38C,]95]eFFIB=b&
c>CB9S4e?9?YPCX+EW]WQ)I7PJY6V>BOV:#FXG@Ac6.+K-S_2RC_7;(RP_GYd9JF
e[SA(49U2]&M2Z_YacD@YJO,E=\c9^\ELFIN:T@e=R39.0[QW<Ad(.b#CPWZ1D_U
HfS:H=&E[9Q9^[X21QS^S#N,fSS/Ic;)d40P+fe;8Q_MYN^D:XT9?J=>-gDGb+]?
4fJaXQg3f,=DPJNIPC+=4_=P[:HPbfeM_UT&U,XdP-3;==EX[RQce))3YM<07V&/
1&?9&)^-#69M&]>_R@Hd1Bc2)_:(=BX6^cHOGMJbGHVc(cQY2H979fFUR(ccGX;?
JQJJ?dMf8E#2\HW<VI0c1RF&#()1W]Y2HCE]\/F/C40a?BAER\CUC;GX6^^BH5MI
R;@#UHB<E<3PZcf61D&CdN&V\I95YVf<7??QC>X:7^JUTYGCbfffTN>]fcSb]fAH
[:a>:YLfY^A8L69-4EPJ(S4)UEW/M_0_[:\G#PfCH78?[5#Uc0S[O=_<7P]IITIH
3dKUag0d9T4MQ7AD4RgF#0AL6)(OR^D>R+WDJD6T_^&=TZ5fO&K#N#TQK#LFfBW3
Mebf)<E?QI,AQdg^Z#Z+C?^Z2XIGA4Z9_Q.VAPRYB@C9-:>TNd]YMLT/e(fKGBa>
A.8)]JXIZ.?TV?HC[KQ+[Ec(M+V3FKSE/dX[WB;&?a=bcT8TZ@#H)d)WH5?:QJK_
B1_[#=::a0<H?H07S7U:5K:,Y)g&]bRW]>=#c_Md^)ce4Y?FL1JEebG==EUT8_Dc
+W/M9&EXSg_QfUU5:Q.[I:I+S04MX8[fC:P?>+7L);1@68/4MF\LS<4.N^2.8N4f
Y@B]/XaM?/7.@#HSUT,aU=EO>>[;@MXG6J^,UgTCLA#NS09]D;<KOKQ]7PLcY[M<
?(7?P[ZQf1e(Y#DTQ0K)Xb#F80LK>@&I^B8P#X_56.M\80TYI-HFWdUL:DTW1(?<
L+H65&1ERe4J;B90RU&7TK__28c1)MYRE0C-3DHF[7IASTPJd=VJO[OVKBCM8f.A
A2PZ&Ng2?,&bH-Md]=Y;EEJGWK^+W51b&c?7)I@d)g/ZZ1C7I1+?XgPbHVQEb99e
47AV5JLIPT#L)0OGY<LZ,3>N9eI1>8d:(C3^L=b2^#(I#FKZe^f]7(eg(C#7f7_;
T?;UUKJ]PF34C(X>LF(@HY>^cdLPffRJf@[R9,U(Q11E/4b2gBJ@bZY[Ja8#J^P6
M6eR_S9A.)YcZcXS@/<RU<M3f)QD.b#^P+(?/][-HA:O#)H?ad0\YQ17f,dGXb>]
dKJeC,7@)/#&?&M>^PfC>,[5\-Z6TVg-BK5cV[TS6(6b^Ng=N@EQQ7Cc0aB8Q8V/
+F+D#]K@J],#Bb-@)2:N?K7Q.Q0SN.Y@:=(7NV2c?AG(]gbfTYV<;=J63aG8cd2?
dK2W@?XgeJ:bA0LX=\7/Z(KRO9\EK=-D_<Y3(<He]?[@=DEFbN]fF(gI08BD=7Le
\+CCE7ce+\OD;dC0?Z58[OD;#HM5=7.3aEEMPObf-/81)@8g+g4;-J20=<B<.FHg
39c5D3#/&-_K,5eK]V]^.EQDGMI8dQOW4,fDT7<ML9:YS2K276HSC8[@/8[Q6aW=
?e@cKC>&4@g=(Q+Z_ETYXeG>RP+S<K/W,&@E(9YDEeC,S7fbI28C-^#B?cZbGBCK
g(R]Fc+=a?a4KP8KTNeCJPYd,e(NH.7((5+e..WcD+^VH>K547ZTM0=aeUO\@>BS
YLI#CLBV1;,8+D.(]dERXeTQU1QEE4=cJ0_<C?CT(XX;NZ4/249:9N^P^UQ8Y<@N
<&a/RbXgX,9Q#bO>Y0-OGdc([L#,\6KEePX&VE8Y:J-N4OO?V:a2:Z1V._BY;dPA
e<A3.L05M;R^\ZU-eVbFAMJCUE\&V2I7c_:K>dbLQ2Gd/@GQWJJ3\a>#9\U4&a_^
YYJX/&ZTJP9>;+U83Q1(JF^2&]&fAPUd5g?\\=?SO:1+@7]CNW=gL)Z)KJ\&gO<M
g]GL-H?Y(4b55N@6+a;edK<0US]PB845H=Og4L>]5[ZJ@A8S8MeD2OT0,MBJFR07
fcZAg7==BN7VgX:-gLWcS(06+?Dd0AI]LGW3Z(_Q:.b([66bVK-8:<aJdT48VUe)
1HS-B>0B2?eA2B]Y7)>__01dacYE9c/bBeDXTJ2K3)^e8<TCGK6XO>)AEVDF_;T(
M.P3.-:fYYYB3RfZVd-FQH^g1)S;:Z/a,gV+PdbfO#H5AZI^V>E6TERMa&\3=:3P
E(d)L?T.QS9@MH;5>1U4<UC\KcT.QF0CV[FR>OJ:\GKc2D-5VC(PL-+JV@GP>d;f
COG09e>3U4V(N:#T,AX:LX^,1_e+7()]#OG@cPZ_C(c^X5>=&LX&YW0PA2\M>IK4
>3?0AVgTLeV3>W^5HI1G]\=N9Hf0_=-e3,D32gW=(bF]7:KJWECTRL0O3=>XX>=g
ABQGH#<26G=B(0.P=d]9:TQBRY^J;ZO.:C/(,;gURTg:?.]UDB:@SG:[PfP6GPNF
H8&I7Oe\M^0K^@J+6_de#RP>2:3N1.5YYG8GHJacD7&+aP1N?40MR#H]VA6U(e[I
\NGT<YXD52;S:GRS#0]g[Q_/UJ:[4UQV[WYOFKbP8OM@CBQ7\PFg=d+-&M\XRIS-
eBdZLc^a]cLg/LR&KEc<PQ^=5C@#+XH8:K:dY>H[a5@]3<Q=KSb+))=5EIPI3A9W
S2VW,_VKZ]&86\?8TFE4ac?JW[@[8[/a&aDfZHUO(@eHebY6^;TZ>27K4b8Yd4VW
Lf6IMSAGX9G;J=fCJ#@/DMHa0dANT4XFV/+;,355Q9R1I<3)ESJ0ELAAFd4@7Ec&
93N2[0_)OA@Q=EB]X5bJOT1V8LHOD(?]AN:7^GOfS06>J/AF20@Od99-I3_dHU=T
PIc]&fLV1IGK^D5O[<58]X=EYU,]d;9NVJX#>V[67A2,=C<(FUYH4XOAbGY(dA?U
RSbBQBQ7CNNE4K&3W2_W_LJ[8GV0\fL?:#=3[-c=RdL6&WB2gWNJQBW0+3P93L]X
#04-460QT967@MKCFC&f,U+6><S2=]IY,YGOZCAB)P+40-THJ_;25eTC,VX6TA1F
#K-&&+)STVWWMK>g7aF,++-g4FdgIMO)OB&gE^<e.b#GPS_[EUM.FBR-_#4:8(b#
?+]?4.I.^P.V.R(95:0e^gTP7&Zc<=1EJ?[IEB1D23=9G>,9e..b0H2,NG+MTS8d
4AYe1?Q:E+c05d/YZXc9X@R&Q=\de-,MK8P^U,9AZ8O]6<2PaNRBS[g#e&5X.@])
cg#QNX8d]Qc2c91H1#WI:MX,EM19K)9X(P#1a[F&K<Q=M=#eeX1L_.X?\IUDWM=J
YZ7SRSG9355HgUFA8J\CT_01-gcV/E>4B\@b4gRMVU<]g7L_5c0AH6?5H0a-R2SJ
,BRL&6/e2&gJN+=VeI:H)f;W(88A[=MT^ESPQc+)a#[g-6R+\:VE+G,f>B=A(SKT
XKK\]=[C3KbU24#LTM)9>LS34>1[_Q2XB=BD<8=_c)Mf9=\1A3+2c-1c8&:G;2(<
EHOG&2PN5MIbd).8)F,O(KgAcQ@5-<]=9K<L)QHc1_?351:_XBB?(=JGV9-05<Da
_d=[BU,(F.?DZ0Y5Gag?W;6LN(0WVI+,?g0S6+)ZeGO7_1JR&7b-#Fg4&ZZE+YD(
I:GU5,g].Q68ZX_@5cL,VD+2dJ<->95T5#\+V0b3?B;AT/H1QfP94EVEYDY@CHIV
.^>eOCN^++C7JP8(\P)ME[[[#5VD/;AKgGM\/6X@f/JL#^WaW2,;FI:GBS/JF;-<
e:/(SE/?IRXR>&Ia9dLbK&;-2C46[;]I<,aTR/MV4>Wd1e/f)1;=(<-+IYF.GZ)G
OfXLJYJ4@D3#f+<SO2BEX-W;OT#e>FIBRZE,QT)+IFcKIBL67LGC34N?@0,d5S,]
&]J+4)9,:_-<a\dHP:A+T+9F8PHLE.]@[Y;>cd.F/8_L3^;O<&#:A[+(YS:g3T[O
<HZ@&Z2CSbT3X[5N)XNJWFKL9R(<(&Y0G;_SUO0\]cVVNL,-JBX6O@.@[#2-&D4O
dG;.S3d=RVgRPbF:3V]\\[R9KX6SSOZQO=7EH+Z>][c+YK>38fX1L3A<F;gNVUS3
R&bYFM<Ka(^P5B;D.,Q-,\C2/EJJKBYZZ9\0\0_C_GC4A980cHdcRX4)1.K5Ogc-
+UWR_^.;.Q_Z#[]6#K^Z5HH3:68N-A08F-&E\2?,fK6UA9\64H]>&Y,+Y\XJN=,f
D8<.bg:D_O^BZLOdfV==B9_5,T3U-+.f:=_9FRER:DdLB:LXbVP^6cO5AQP[\C]4
Zeg[ge0Lee)3ID4e,?INHG8\T16b\<]2d/,:bfBYT>G2#0Q^a.P>LY&&:/+IIf4d
H81R^U99^MQ1@4aLE_[]4<[T/W.H[Jd@L&WCRT#4>O-dT9N:5g>>4L67#@K@QD_(
V&27^B6J(c7@BVGg1UY8.]aWTZ1E32e]+/Oa5.8)b;L]M(]S3=KA3A.L+#:egIG#
4_UV]H0.1&LX7XUEA/PGP+L3>-J?1_:)<;->=a+aC.W:<C?2<W28gV8LCH@UU++3
@XC)=PUQVW(6.Q9e+W?Q@H:BT7PGSfJJaSQDU]+A3=R@DN.\<g/(:.#CFKZ&F)_0
bMTdL8.M]#7d-GCSVWZL3<PSL833?KgB/C;dF5(FZ1Tc4CW_JE?1O#QB8>Q>=c3]
J\=8;:.R]D;Z;TffSKU0[-BF1d#B@#)GLNDHgf,19V_2K0\(=IDW@S]geWVWS\FQ
2R])1Cf0fWceY]LX,H(&GYT>McT-JU,5CV6=_BI5^^PM?X1JO=],5/[_M#.Z:5_L
<81RNdG[bWG9>9GDeGO?W<+DZ:X4RSC>^VZD^]KZ8#\DEQ2N30+^e5]ZWO(U;X(Y
1MK#7&OV&;c=&S1JOTZC+FVTe,0I++2]G:_Z9/5]W<L[57A-J#L2Rg7]8R51c/>B
22OfN///5fLAY1D]Z(Z.3Hb^Ze#b?41+<3?MKdQ6,.J5570.W[UVIC[R-=@U)KK?
/EB=1L-0<JZ)ZZ+U;K]MO8&9C:T/RK-OeBP48#gX\g,O[V0@J2(2TN_^a:;T^4c2
E3,:D4XV:)ODOCIE-M#C#;.@KR+&Bf)dM_NSTd<KD;#;6II(E.H5=6Z-Y#3)bD0[
a:>MT_+E<-4UF32J+V<e-6G8/fA9aSM/]FB#1\/bKU1FOKeA3XXEUAP.@gS_c;-^
=G]DA+BQCNU2R6Y:I<@(bT,EMDY#3CS.7S,1HT,DX&-2D5b)eB,I3//;ZdN\TbaX
JB^M-5FRJFOb[UCWbYg1.K:KRGEL7\/6,f?CdgVJLG7\efGT(ISeXH1XSc/P#]M3
]<f.QbNSBX_T5Y#QJBAW<10HKBK;<fB[FeAUB+U=N2<\H[PD?,\b2#]J[_PaK8AW
c54BaH&DY;(E?Za^,E4?WO>SHV&E(7#d:Q;PRA><\TN[/CYg:D^Pfd[dg?IRF@J:
(GHRHaW2<QBgd/,Xf[HNc\F]13<K#7KCKM3WUTN@>GRSL_>N/^X3(K97=?/Z16#H
P3DN[,8[7VPL52Y6_6_M&?/Af,NG;@;D528I09Kd@\[Rd&0]f_@@#WW_HIVB0CS-
VQZ;[SXA^>@5?;]0],V?dC<&e]>9]G;_a\VC,_Fb4M)e2&(>,a@N?-I4Q<FR^.E^
.)DP]NPT@<c\>.VT9.7KH[<[dG)_L1c#dF>U4XNbOc:Q&:B1#XXbbTIPb932:C,0
R@A1,(9#TTK:Z6e9M(Ad<d.8BRT7eU9V[^KA60+2O7Xg\+FRKbYH=,6\UH<UgO4A
PNcG>9dTG/1,c=\S?6(B^\M(3Z33]:R6Ua#8(D60W#Y^)^UWcUC+NKdLC\=K<IA8
NeA0U2/]LOAb#^Wf\H&:GH0.d5:LB/2=PLKO>(]@V@6Q?K,NO]3DN.4K3fQUe2-#
[&L4W)I0@DA;f<5@AH\-AGcTf45LDO3W[LaR::S8YgI6c,QT=E>RIPF)EG_.6f<H
5IKGCB(QDS/bXH=-^GRgS^UNf\Hg?]-Wgg3F]geV]@]?7cD1)M47\Q5&/M2>3_6+
=@NDY+;b(YKCT2QFGEKKB<J?4?eX7QNf=eGCBfB1SE9#eQ29A>R?G\BSgUeQ@1Z5
FacNHV=cK.^-,A;^HIH?ZGRLBO,Kg6U6B[_Q+Z+Y[;NP,F(JDa-RDd]N2gONI)FZ
X)A\BdJQOa4>Iga\e_[7T^AM11J2J]K-8X=Q?V:)gS2?D\\3P2XX_QY?a0+P@07(
O1f6;Uf4CCH^6@F;@aXRb.1d?dQVbcT4gZXFYP;._=6?e[HD8?_E[4Jd7MM(Y#^M
;ZQ6YM>2J@N44cBWbc((&]=--5;S9H++@?cfWTcWMRc+YC.fe0Z=\3MY0>@/&2P[
JE_gG8DZ)6D3>7(R()8fDL75a13;)EWDc#&?a-PRDQ@FKLTOVe976@N4U9\6SHQ,
\.D_0\XQ6bXE,MYG>LdD/YJAZ@6R8+LOb1B=&N]@XbZ,R/R<fGUHV,MaU0DDAI;1
f[2(5:46d8f:X6<UE3OD[<@ZZZ[6-:aJIP\\(=[4MPI81^GKIX.WMCU6?(+L\J9b
J0EQ[3S>1HIXd<^=X<LVLd,TPY+:gc;2,[]9e8(EDcA2b<9)HUW8&#,f4c3JCCeV
3ZC5,W:_[\33T<(R4@-20=2K\c=gJ/FaaeCGRLM+THEO4)HTcdH4F[S:8C-I;d43
Ba)+HREM9ME/340KFWR6>E>2,5-+cMVNFNES]&#8,U8MKRX6a3g@OF-W:C46D@ZX
.M_^Q#+;4LeD=K)MMf0863N2O7&I_N/fV&bFRRZc@=YRLD9Ld]=,H@]OU]]<Z+^3
73bW5&W8A+2#PEO_ZH2\<EABY.bDSd^X]Y=^e6OH,54,Y>MCTe7QdQQ#B(ge:OXO
?=HQ?I.?]<g9M-U5G20YA?&)0.^d+5LA\c=J9&UF>=GMS^HI(Pa5<Y:81=1\>aWW
OSPWTF,.B@,cPS4aQT)YQ@3,2PB,C^]85]\#Vf4W<)X/d@&BQ438J2NY>CQD(/1J
IR&e5D3a7B>[:3YJX:>F\_B(Z:Ge.)a:[N+bb=Y\/9^><b5Ca;6Z(<BfWC4B7,T-
Q?2INFH+S(5^GOb3/S+F-L(dd8eJbBPd4Hde=MIO<](0FMcZ0_Y#ZIWBCLQI>fD3
@.Fe=eU^?)@WS=:-GgJ]-NJY0?#d7?Je_R/_g<>cUGM_MDO^4eC.@3cE>/;gO^E;
2))T1eCKdT+bdEZ7E;[#M10DR1e)3?_R,[V#/PEA3W<AdfIT+-RZ(7H9G^e:M4P3
A@WNPeQK9^Q<@DSc67&Sc=R_5.+(82<D8\K2_BI07DE2^RB04K]f(MA+AS&/a-D=
gS3P4E^dI^D=(&G?S@dN6>0NgAM:Ja?-J<E>PdFI_TM2cGR,V=bRCc]?;BUeQE4a
1f<REF6AA9KH7dA6/5LX?U/004U=Q1@V?c5ALHU+LM,IK0YJ=,I)C[=@^T7/-P:O
#B_O2)[\d]I9W4\9[fV[>KC@PRFQ5XZ?+dIP^,f)1G8\X<U05:bH/F<b0S/HcDf_
FM>ZJVI^C\5Z+A55E^/0Na3(<H)6PeMEc#B(.1XM)W00UYeSc72I9@Mc1(61GM.E
HH(ML+bG3U4):->N&IESU&&#4TV6dJ1H/bH4Yg#Fd];]8JTFVO9>VX:V\>)E?<@=
GgRdNC,f<cU[;eC-Y#.L[9-KfbEKNH?-7@8=67[DJF.^A,\Zc)@e6,&-Rb2X;1VQ
e_]1H5CeU)b&?//eY;S,E<F&E^_N@0DNN/JAM&&ZZF9(A8?32Vd1)5#[SQXLHL,?
Wg.YJE@b?d:[C&L&,5AcUQ,:.#RE:0KR2LgaFEMP3R;&:=?3cPR#ITC\[eM8B7OP
4dcf9(/K2TK,8^FX6.DM0C.VWT:bSA#8,,d--6K9TL]5&]U;[:4\fJQe/_-GG^)/
K\b-^_53QO#CJJN@&e;T-L-7-)MeRFcPED-UaH]=D.dG7Oa<^M82Hg>WgCJ-W1PZ
G:2VX0X//fBQ?\V#EI,8\[O.?-9SK)6=c:D4HJULJ+[,)YMO]U+a^QLS2_gPT[IJ
-V@04247Ked-D].dM#46aK_?c_=9O@N>L^gJV6XAJ:1bW/Ie(4.R1H:W>A#f4NFO
[W_TKZ^(Q8J&1&F/gR2ceO\U_+?DQQ0?D302,/XID+N4/0TR5L1-\)>4Ta&7IEO(
/6YP1LgfZc3Ca>X=162NT^T6N:(=#11RH2g-.B:[>/BWa(3B,R^(:AYd-/JeM^9V
O0#3BMT8.?f5JUB6J82,47\,E&0I3<TT^^afc^BB_,]E7,:(fJYGB.WT69QV&T2D
=5eFY=--))4a1e:HLC+ULD=/F6SH;@Q>A+3^3ecH_fV2ZEH9JPV?GA[[TGV@UP__
[)9)R]EB-2E^aDZMfT]1_U=#\.aPFG=&S/3R]+Rc]gTV5?3N]]#;A5B-2a#LR2))
,9b6?;5>&HQA/,b1K9?KbQG4O5>g6QG-=(U.T&bJc.8G@)WW&]N8(,Y&=SF-4e^:
c4Jg-a)&#<JZ;=f;TQ&-]:-]L9A2YOe.J(D(.XCYQ7C9JU[O5P5F_FQICJeH>:P/
Q9Z5(g=MWP[YR3LN]BD37;@eU^#G4L6QBQeUb)/>7S0FfU:0LK4YUPXHHUc6\T8@
^T0WHY1;[?feO]VG#JQ9SWcC_OLeHF8&C\4FQ9V2[U=\+TQG(I_D,B@DeQFc([J2
Ndb[;C,M/3=J2,^QGgJNgZ<Gcf-EJ&_1F79>229#>&<;^,P?9CWa:9IS1AGA:6[+
B+&B@#G8]HU=/8FS]]OI2beCZcBS&dg.6\f,<5VZMCB&/cAX,O1a>[XHBW;d).]1
W]#B8Ec^YC@Q.=\O?eIMOAMYDAS5+?@F#;7]TQRWaQb5TY0IZHAKVD0+OI7#O6U;
a:A#GLJ/7CA^QJHF^_=Fd1R1?MJAbR.<^LR\f<A7_C.<G9Z#0.VbF=#c2[N>DQM_
<gE[OE9S\/,3gF<>GW28R8M+)eYe#P7,HU[CVMg6XdMECgGG9Ccba<^I9&CP+Y]J
_@9_=>1-e8KCIOa#dC,KK<NOe&9?6]7X__BIB6e&R7e<80H718]+=/LFRAIH6A3d
LKOc+g[#&+Zb?A?a^8V#JEcHL:KgTd#bO\9KbT=AN6N-O32NWY&9EPL^8#J5_Hg)
2+SD_LBYR(9MV\9_+\5>CC;2,D8bA#SUYCU=4+N6:0KWb)=9AG2IOd586=T(e.-E
0fgQYQYP5)\JT0Jf\Z@e^1J]5gLI5D;7HDg&7>:?]>H]+JZO8O5<0EL-KV+Yac-K
,XA6EV6W=a:7YWX^;6BM+S_?@JA>3RYJaYZ;;JNE3I(=<3,V:]Da01X:dG=6[>32
Mc;((a[ANZC3@I?f0\(YY8aPMc@I9LIRUeae=[;(Y^JK+HH34(;/^_g)J4BA<9/5
Wd&D3-[1D_E.K]e3LQdJD)MN>Hg]T.^B2V8>DU@8EVT6H6:/37VL2_Te@4eELeg@
B^HdbE5FF:;FbIc_ba\6e-4VCGRN8g)HIRUeZK1^^L)I2IKIJ7M@c[G-DfTO9?G.
LV4B<Vg:b:J1_C_61g&6,T:1<(;gg9_8UA//MGU@<D0=gSRf6GE?(FE6NXE.U[2,
@R?PSa#A)-@GDY_V,8ENCbI3)P/=?U1eDQ?<^8(#gZF15gcS^,I,ZXWITOHDF/4O
#H1SX3XUVDT4BC6e^\dDc#\aAB:<AEP_R6-#df_67f/+WE\-^Ge:;BHWbC:eTZ[g
NVfK,QRPZFd(^5/C[ODE?be^Uc5_WP-LQF>QL)H,Y-QD<&V@/79[=QRaEFSM)dK@
)UM\F6aKKK=?8Df=.GEe-;XZL_Ya4CffM38O9Z&eQGU#G3;JE&WRN3fXQ:631<48
@RDL2KNEH4A+JDe:>8&g&(0_?(E14,AE;)^T/62R9+g9/b-B70;>>DA&@dVN\Ref
[5EMdRROdP+cM]f&45e[LK/#/IU35.\P]Qe8T)U9O2fE7YD:aZ+OCWKBC9(RaP=d
/54cB]]/W.Pf;50gS=OB1&(QMa^5D&-1a9NC2-G<T;_HS\F1VDQ@4WH<6dL<7@Lc
N4/)&5X&b4X.YI?eXd?&I]-=9FS+#ITL+O:b52Y^fKP=4:c1+>[P]F)PgO;9HU)A
88LOCW^PKWS5S&&7NDP_L.V&e72.;=D\e)TL?U9+>c=(e1b9MBAB:3IAEdLY/6)a
@g;5)Rd@8W;TP7bPE;E>]<?,GMSgN1]1?9#,F,P=dX^JCK9?aHKgPAT.VY6eB2L;
E&2XPDNNe1\<A;QQ1RX._CDN^(fX;U1)=F>T1&59a@IG0#/6N\_J=IeKg&^+H:-1
H.+)UZMFQ;>N#OLS=H,XF:aVc<VT\8MB=S37V_.57O8U:HLU-CTJ>UNKbLXe-7J,
fDCF6<YDI8]YCI0a&>2E5;HKgc?4/,ZeK,a@&g#,b4.\)H8P(bD#.28C^bXN#3#I
5eAA8>JV(@S,K&#+14R_^)4,8[Xf7@8^2J?\-:3SNLS=^Gc<eVF)]C7J&/>VMddN
1AcP49S4P3-M7[2:fF&1.gL&gNU40D#fTQ;A[TY_-R^efMHGYW2a_PeZ:>gZIde5
eEJcbS,8>5TUG8FK^QW4Q?E+I.NH@)\d^LHJQ?GI)D&S,LN0952.H96[1VE3H.G8
Q@W@ZXZ8@7]9<O^^[@@6F>\&;dATR6\9^?O,IFZcdgIY<(D0DJU;_0&R0C+5B49D
bAJ-.V&F54;YO8NYGF;U0>&WJGB@C@O0J^S_.F\<Z25^+@IF-6(WB.9B;CZ),F4>
ReY&1.]a38N&23\0+-J.e+FCfR:2_^,ag/01+B5JRPJ0KE7-2WeL+eP[Jf_?&NCK
O2-DSFc7,a&1HQ?1a7SR_3O7\#IA^\#>BC#^HfgF5c-T#K\V(+LL6VPd.-R3:K.M
L,VFSSB?+BPA+BX(Tb5^NgSBaFX\0-9[9;1YU8A>GO^.bTX-@<XLgf&-Rb4TZ-#H
7NWY.@30@S=bTf()5[(K4V5<+7b/(MK6L4/=<;CP+9VbcYdg1#fAO:14H=edYYLD
I/\B<>XRd=e&bR4&[P\ec97NX?c@4ISJgV[[.VY7Q<.\)]2KHAd=@V]BQ[W3Hb5<
_>+]XCZQc)_LH0NDPCS2FX1Y().0G\J3.O4+5I\S-1R8,-dBe]1_-N@FBaS)]:LG
]21/A?cN]]?Qc+.aN0fHgcGO:-JY8,JU>N?dJC.NB?.1HZK&a3P[M=6.E&BQCD-4
2SbL=TUZg\]F-H+K8<Z)LbE34DH-1R+bK99e3C\8Ge)1efIH>-YA_JVR0eWYCPHN
Z>9GSW,0T_9.LdfDC10H(:FGJE6BdfQfHWMDC83T9[&=)?C45SM(f2cc?=1VHS4A
PM0KH48R]FUCIF?CfHc^+V#?5.AZ&,/Ia5(5=8>G\:;cCB?[KH5NGP)GB[(UR9K)
3WUZ4BGS66+XIMM0C(+_b=P2K0Y2a(G3-Z)beUB&8(^=:;8H_:c(P+D^Q21e.XR;
G@NLUY-Ec6IVMB1X1P]F>7.aO?PWJ<:AUf7@3#4-LI4a7V0M)XTF#TF&+d^9P1Ee
()#0YGW;I)JPZ#73AJZb0dN-\U7#WT__e_d/2&975INX+=2D6>91dca;>+0K55F\
LHBO(aE^YDZOL4=_5-X&GW9W#WP,)@XXH#&,-8)1]Y^?,5VA(fgP<Q&B+;W_8d8N
52F#a2]=#=:-@67B#D0[Q7N:-)4A<VIDY3>74T4\XNcG2KbL]+Z#Y8S9YM#.:9]O
-@H+L=0bLF:4[H4HaV7c]LMg0f[EYM9K2BHB(AHeIP0Z?Tc6U.\Q=Ode<_T:)T:&
>5b1L#=;PM>;6TI(53\UWgAW[I5):G1RC.=Y/1Q]7X^Fb,T^A7P:<M9[4XWAC(8)
D_(O)WE6H(ed]Cf]AAQ^VM3Z2V=N>81OY_F#b@B@(8G>cI5cYPQ?O>c(g&/KQdPK
(KW>3<2FFaaI80<NUH,?K??&R81D7);Z[aDV96E?QOPKZKg[I#U>R2^f56D-+@0I
=,65,MH]K6AS;13@(=_=c79d<ff1P>9\=PW@B?Z:_)GK.Q:XQ>1CdEfffbLZP[.W
3:Qb+c(:J35KU3cYOG9ROIaS6C\D?@,ZHTGG90f)@)eP\-(-G3&V2ZF>ZbCFURTG
5=Dff:SW,\&KGKedE7;9;+5LX,9M[)3=cIZ;ON?5(YVH,:c[69-UH6=;U;UKK45/
g^XPPQ32H]MIgaXB=+-McO-4MOZM1G+RZd1S,3/A6.ECX28adBaa/0>/1=PF0N9d
#XXAU.8/2bcFSSe_W6/K?<OfaCF+#I#\=+WJ9dbf>[.^+300(W7:2#8UBWL9(@Qe
Q(TPI9BX@C9_8G/>9EDJF>FNT[MHX[62,M.P_11gUX,\[K>JN<50M&+-[=EcIRXN
WQcUNI;)ebN?N\E7eJ>B<XKPLG3.4.B=e@.=dA+[,93[)E-_07fKJ71Z,UEbAJ8T
1A^0b_M;<:@SL6/d:PZdFA22;?U;^@4&XW?-S_Y.XE<JXgV^LKC,0NaR8?1_,8Z\
M&>I_7SH-J\cJ[4I5.E#G#BefXYI8Q,/]4<\97C#EE4BP(]=B,\4EY;/>@dMJ7)=
73ZWMH+4P-H5,Ia&&HBcX&=WBcHg+>YHF1g#cCJY[#fbfE<O349O6V-);ZUN;DW3
,f_@1.W9C-d<cB8dGG&W,)09Z9E_+X&ENKaHbWaS[W2S:4VGBR8bTO+28MC_IgZE
M0;\V8^C>H(bF[&;9;3W6>O6;&Aa<c=8=(^)L\;fg>f/FHC,808gU4QaP,Y-ZZL:
#dQd.D?aX?;RC[bW8?&=3-0^2,ME2.[&HFD^WT=SIV>fbaKNb)+4_;SLa7WE7e#4
:\5&)=4F+)Hbg]9X_cA@[=]bJI.<;IQIX4&[LaaA>R2>A_X;HGJTUI)>NIOMg+H@
?>7?)aW2,DdBb7L7B=NJS7B,[S?BJ+;^70RAWd,0ILJ2&>aBLH_RV0?f8YTFYH]T
B1;T:=909/Y9[+R<>NPLO(EP9<2BYe7b,TeK)90?G#4Y(\G+F92RIQf1GHWXM]LC
J>E=/gT=-e@HUHTEY<>IPE,T61dJ.BT2V709JU.eUC.IHT^(KGPd](?7K327/+aO
_3LF()V8:XG)J&FcVH4_+@=D738:BDTc1LPT<:E8bSQ<-S(QG;NHT)5UXV_K^XBU
A23ZIJ+0OA5)CN5Ze_J\H[:1#Z0V^U,9aBLD42[+&LdWAZ6gLf&[Q+Ka0&6R&<HL
XW8=SJSe7YU:2&0GEg9QR+-/=G=eP9K#Q7_P)H9aZJG5@6Te8(75GBCJ-]a)PWdP
D2+W6S7M[_037>+[UXR(<]&]KHB-RX&-;FAXL/e,\4F1]_6#N5ATb#M[P2C&KVBG
2^6eIH1@+FU]Hc+#d7X&YKHeTLaFP;Eb&KG4H(dOOEU,];61G]Nf6g.IO.G\&AOY
\]Q[]S8>_R=K81bTJV??IS?dAP8+8eR-RSQ.=+[,R>A#C,1bP,9<ME19-1IdWeCO
D]0dc[(>Y2\3)&)8OYdPTQ,>Q>b:4>)&WNQWUJg9H6\-HOO^=+FD2)U8HPV6681U
:^cP6_O(N\We>6H^c@,Vd]A]1_/BJ<0JR#0:1EN5bKDAA/UQ]JCa>eFE.dM+KU4V
2(D:?VHJ]UZBHUE\c]]L66FRW(S@#aOB>-Mf8S_>;ARf6-&X#b2@7&1U;0;e75cJ
FIb][O\4.b\K?F1;bSZd#U=,Gf6:eSE;>#GY^;gL\L0#E__da<C/eZ]-#C^c5&C&
@=9Ia93Va@.)d65,(0T#@PD=^Z@>?Oa-fTD/Hc]ST&H_1F/JXJa8GAL_ML8V:Ccb
96?[;+=0E06]0b,P7^H)IMDa<]Y[<QJba=XOP3f,DMFQU7T^;ePe:-#1>-32#&UU
D;.@)S:>KY5a]UX^RE\N1[Y:X@I9;YWD]VF(K<\QfVBfE0R3;c/JS>f]f)X9HJ=,
fEB8+FQS65&<WWZ8>gY:N3BMJAMKUIH3[A8@+,2R.\=QR@aNT[;[;ED07AEb?&(H
8OO#4)DRT]6gg930E:44&7\EEW=F+:f(U\&f_)NZg6^CPH\5_95TVecZEITCg09:
P9NEA#f81SRW>V4ad\B;Vb/9BZH/7SXBM8U)[c)^L,_7/X;74D8Yf9-_6R^2I20_
#DSBP7=GeA)2]gWWM/,(M\\3V1\#?,IOaV1I1)De.CR6#F?DJ60dB:E@6NL2Z>-f
:]RZ)>_976]23Ug1^3\.aE+e4Z/[Z8CQR_a^SLKY0McSN2A#?T(]&bLXD&f&=>\X
O:4MXV<\J8>_G2eQGdU93ZUPX0&YN>9+-c1<XD4#D?X,MN\#aW9C+5A^7XG@FOTe
HgeVRK7J;LO^WSL6:E-XSaJCUc/E8)@GG\^6(OD0?1fJ?14<<2dQ72FNG#+=Q2?4
.V-_HY)Sd0aL4./UCDX15L&?.::3)L7]3\,IP1M.G#Ye]GC>ICVWH1NR/Vg9OIND
W17#R+#c>6:KM^GW),1-A.AcQ#FaZ^]3FJP.CTRd9\5M1_3Cc_;OL_c,9ca3CbE\
W-]17-.5I3QWaRESWEb\eU;=.G@>B\<bZ6OADU1SPg9d@IR+=8OL#X=fW1WJRE2Q
L9+?L\baS.b_=L=GZFYf^]V>Uc.E7TOAA(CA4^ced9+=cG.;C_gQ=F=-Vd;KXM.e
fH5e.YAT?b(C-+W\e:L&1HM@_X\eOY#P3>NOJHQ:/N?3\.J@+>W7:>2#EZUKW=],
+Q6.NBG]f?O,&MbI]g</45.6LAMY8>Zb[@-;;0d6R+;(U6>:&5=5&87PDJebQ6]^
FR>?d#,M_7G3<FM.+TREB)8:6B1[]HgCbS0JT-#G135=O]5ObVEX9M=?CXGNeQ4+
DS^DGT_>,T_5]9eHFH8WgQ#XBV&+3@g>CH]ZU=T_F?3;@VVN,g0I^NNbB,E<)Z3I
.TecAUAC&279T;Y-EKaT@:8MebLBM[2?&@8\V/NAPA+3YE?S,-+T8B2V+)P;]O4[
ZL)3IS2Za1@,GRXL#8#Z?U7;JPgYdJc08J0bbJdODgBPVcL5:5&4=78fI:07;B[O
<bBE7CD:c6L1g/YWK&90+5X8>eJ)a\KdfEZ3ID#NT8FSe,TO5WPf<]K<<BL&d>fO
Z@N0a]_BND8SI@DHd7JA]^e.^^-TPW3CJN)XMd@0U3>FBb1Y7c8N\D;g;-OI];P=
9K9gFX-^YQa0@&LG[6&VPU9PMO9X.JBe@G39A_SRECgH&QfJV7VE#]-?f7b8[[X_
EeRfH:;=;^^3:F9N=eF-@4N&8B0F4X,MSMFVA/6QaPddebQ=O82dQUU?;9MP#:GS
-<a^&J3-XY20bL3;^3MgZT9XcX5/B/47gG,9:5@;-=DG8gbAc-UbUOVMDD37AXGM
U8^+V7RaN2IGUGE=:QGF<?ZTYA-\\D\<b>3460g>(&?_4.R;P66G=I:TGfW1KE/\
]6;;(&e>[A<(bP-FcCSg0F::fIWUR]@1,:V\.f-6G4ae_2Z1PA/0J5_[72a_aYGC
F1AGOQC:L]S+JP5XZ)9814.G5X7VE=Od?2:RF9.ZQ#E6^;c:IK)Qcg44TK;TNWf+
/F,Y=;SU#;9BK.PG,#6M5g97<X++UV5g56Y[ZGQRHeg(3g4.I,YZP7gg7]A+(Wa;
KGH-9Z_O\S@T:/=+(:PHdMON7d(NXeI6GeAQY-;YTP>M\.+edc-?CEQ#-&W@0QeS
90>c]bV\cLE,R,8U/EeEF6Pd1>M4-AdaW;S8<_A7NP_N,IS8gb-Y>^Mc^QK<F?QG
Va5MeNPOa7YHAb78(^8f2/];QYLQb7:\PCcH_Kc(C@X^]cd@NY54>.2L+3MIU]-W
\e?g3),Kfb-\;NCIKdVEXQN9[6N#4=O(;1>RDbBNJ<E09a<5&SYJ.MJ[&-=I&I/Q
QLaM>c@JNOQLLgAN\b:.J&I8#+10^I^D#O2PR:V9CZ;d^[+\:a4H;^6<J]\<8IB:
P,^[U;2V]6DT,96/MV7S_(5]>@W0P4Y&f)7N>3c4GF)T+N-]MFbR]YR^/Ua.=:P8
-FeW6Hb;ZH-K\DFDOY;6g^<K=NbT4,CKfd?ge[H8G=(ALA@U\]gbEd-=Q@T>Gb@c
J?6P?bc)KgF7;SG6\^N_L=bI;;>?6^C5XT;3(,9&R#3R)^31cYC(Q)+FC\4B2#_W
NLNa<;]?E+bId>^(e8MWYC7.K3>;6-VQ=;L/F[>QX5[@8.;fd_/;).QPC\cP:aOb
NY=<>KQcY,Rg\R[Vf^-U36:J.K3R9cIfd;^a90+9a/2<X?7]O8Dd40B)V[3_FJ_9
.PNDDNE/8,8HVf+Y,MU=I#ITKF]N+TYcL;JXBOegAO?A#T7SQ\QCN(UJ0V,R&ZAW
O]I=CcPM.LG/8US<+-BERQ]@=dT;\<68eG[<<LDUK6,4R^)TfKFCZ>DN4447+W&L
J-OFSPHZ?bKP99S1>+g2L23B6.T?HD(<&K#ce[0.]f5US;YDLHfK+[]gBG7?)P+_
KI&M.d&#JK2Pdb]V\4HD0d.HP0C#OG:+]L9V5ZRZ#?02M;RT-Z2d/<[c1_&4--:?
3\c:E=]EW3:#F;Y4c^I+.AO<?EMOdS^@5e.b>71CF?f+UDTTX>e+]_bIaT/#(WcL
ZV,0eC&2-0#IVZ::a5=FgR=07:gW-6^D&VMJZ\_ULH>2c_S;H[9OE6_CKXTbT/8X
Bb[Ud>YE>VXR6=DQ4:I<ce?-ITQ^DcSBYB8^XWSZbZ-b5C#3\;;PZd:.5K(\JP+V
]d5TT[OKSPcNf#.YL.T+Jg.M[QB9AQ:A70AcLKeJ&=\#VI1,_)c?U#_0PD8S)Ha>
DFXK,#a63W2XA9<_EY[J<G<8_<MeEL#Kg901AHg9/N6^g4:3)H.4OZ-Y>-.ELIX2
->R[UWF0O[ZDfTP8J:5\5R-/^UI-N6\\Y:[]<BObMV&3cD/^QGgBNAHREZ/?U,07
>BK_M@-OTZ:aURD.c#3D]8a^MNPXdX\OU\g_0:W@(.=G+B_-gJ?NKH?cKX8?E4TC
bLdOCRT]G6TT9\K4PDQ(/R4_=g>cMZSb57M6A8f@]H3^<_JGN+/TXe]HP34g0\D/
O/@1+M9f/Cd<#2I16W=GRaf[b.Ub:AB+)FJ#EeBFfM0?6d/6MOa/Dc/N;NX6&]_?
/[<OG5>5Ed(RO(3XYY)POBb^Z[^W8YQMT()JHD6_Tb)ZXef,DfdK3ee&?R.JU7U,
]>-4eE0>_6T;Ydg<A\OP#CV\f#7&:IUE#@1<eE:@3HeM([7PTLG5.5-Y0O?Y4_Y[
,#\A3)eCHJTPE3;G\B:[c?)3f.>3Fe76gEOSRV0&4HZ9f0BV,;UY]84WJI7g^WN(
L..)Q0:\:=MT)Dc8d6dW-58]ABA)3S9dNBUNYMXB[NI>KU]M2F>Zd+MX:3@Rc7P(
A>4I1f30_d)DYg3J0LGd[Dc\)G5?M03-bQ;U#)E6b^bH)4dKAP+544F3E:YH#9=N
Jg&P?U@?YLD3c,KU7KSC+U10>S0W(70M]1dcd6F.Z[8T)PMg67^\W7LVM3LQX&/C
:e50dD[O/Ad^S?IQ:ME7?,^=OA2UVJ?W=?I>8TR,U__+;F4]BU0WD/Z_JGH#e&9P
d2DbVfT_b\JWcVQ-S^5]==ME\HNX4bCSK#G+0S8WBR;=+T_d3>>A0C#:6_;_+dG)
A/HR>O#)ER0c-)0XKUcG<e-L]LS<:6F8/5_HV+8BNI;ZCP7^2b@DP#PbA]\#J6\3
.Jc;OV>A:V_a;A0-9=W.KAQ[BgXdJ#c<3P\U1bcB;9Z3@P8O&DF:b]Yc=M>&Y6GS
O^_:WeG]N&TS86YA3b^.^E9C0/V?0e1HY3>1K@;0YgM>4IIDYb<Id3M1=B7I@0-_
3J+2Te9JZL@gE;b/(c],,R(V>54:A>6Q;.c:Y_a4^X,_[4SY2EdB>A&U3+fc[6#Z
G./?>G\R&gA@V^CJcJX[dN:&M;^f?V@5DO#aF;]<[Ub]gR&V/X;24LLK8.c^DFdJ
IEg)6_C@/cHfc@M\S:KZ#7HZTGZf+A^0T66:EYA_QaM^(8;P#;1Q>>G0+#RLS)<W
4^RVC#P\[N,>XLQ\:>S@W-071(ERcQQS<g=.QH^H@Y-#=Z7LI0[]e./OW(-.C81[
II+Q1XDVYR/=WF6[N&a_.S[KK4[-AXB=g\<3\b3/=:3J36I8Zeeb(9<GEe:f5H=<
a3?gF0]c+H46[J:3\>Y\GK=PQ[4<>R]+aW^aX7Nb-V:)9WAOENL,#N956gYL)JR-
^Ze?>E]IY>^E=dXLa8Ka=AV12aMMX(;Z\MH)<)7S)UI&XLD2bfZ3#&>a+X5a#13Z
18aF[5eS>0MPR]]S#U;aBSSBW0CdI.TT\<2N7-&/M+-6d1./UAQgO5S.?J9P5Z.K
aA6ECZ3EfU#I)T)]TJ.69QFF3A,d1HA172RN)7BOFg-,WLWeZ,aWdB;[K;d<;eIT
W<g.M@bJ8J)TW(^<.E29J]>eOIMX>5DJL9Bg@H1D(?;.+^:50>>]a,W1P>FZe[f;
eNU6ec(<c(#2c/4]c]BgC&ReS3Pf/4(OP<629DWQDI(+\FA+TH./G-+TZRN[?][;
&d@#5Za-K7):4Lb,eKJ3@-Q?S#Zfge5eS/;e9?Oac,a_B->(W-)VcFY_UD<&NT,=
2^<>]W@HU2ETTc5_6HfF)R<:[b@-g17)4Y=H-/R4<).MV.-W4\@Gg26.TfRP7&R-
=Q9)f;<_;4-HJWRAJY<5=?@>IH&P9YAH=1<SG#(DdM_#BBEU_fcNc=,UABfXg8da
EgP5fSf5TW9.ZU2R<A[[AV]B#T)T8Pe<9Y[]:ZC+=DV1<OW47HQ]507L=<K37P_W
<,aPX9aZfTf&KO?R[1/gTCfg8IORKaYgW>KAJG[.3RN:\gNZ:LU9R=aC1>VW4Kd(
4#X>,1UeZO#7=U(PUWY\W:K7\195,RWaL^(E;Y4]QV6X03EMFCE@<(Q4;KRc-WKR
[fEHbTM,_OfFc][g,:I:V+]<KX<E=/P>@VRQZdJ?gO)G005P-G=1)#4g:RI+8^)Q
HC<Aa4NQ_0&[J8FCY+Mf(UC/?Wa>(+b+SYY6F>ZK2D3]#B6@0f7NdDIBCLMLI@]4
=E#W&cI2DR;]Fa7IZ3MLa/D)8)-N,d?AM\64JXTWM821JZ>4H_(bM=HG,;1I-EOb
.<LR08OZ+^Ja;[?O=d<LWFe>Hg-T0]cLF=H-AWHS_/F\X1g:M@&9>QD\8]e7P+44
L)\@;;(cO/B2O3]c?EV+;_9(^9I\I5b<Q5Z=fYM--S)6P)R9gKN:QH3D?ZY2;HUa
++.Nd#M3YgA9_.c:@;9]5?d\0g_S@6;KT/J:5eg5U>2JOY<MEYUDS[b9PPFY1>ce
<7],fFf0FH@QZ#U=24;R-[,WDAWa5D+ZbO^1[;Y,.L0gHVT_HVcaA.T\W.MMA=3G
4.Qeg\/<(;RDF=6NTA5)F[<TDZX@P/K0ZR_M-5Y/Q8a^7@JS&M9FJ-E6LNEYRF(X
c[K3E>MU>+ES,E>V>\e,#)f#HU>ebQeLBJUW>SS5(N#g/YaOcbX.e&TWF-;Z-E>U
2c.1)R5/O5@:CCVKV@8f0[/(#7JYZ=YJOE?;X-U,ESBe<QMP781H;J7Lg+D?C)[a
RH7L_c9>GJC4de(46AHaZadb@QUGRg&.OaB<RF[#Bd_6e7/,bH.D.L\>L>:0&d?b
E&OT:<<GXa<SK<7d:VBb;O-DQ]UaS?1;BOeT_>+WA29c6[dC233_A;<6EA_QbH:C
6:Ia?-6RYI2.+,EDb#f<]79H5]a3V+4TQNH1M(VG-Se9>(LWNTd4T004=0[I(F+T
9@8:PK[M4&(CMPTUa;7;<T@LdP\2PUa@)aAIG4E6H\Y;4-JNO:3^.<K[4#(E@XX3
Q)0:_]P8PUVc&f]S1AaI/[3L3RdKF==><I5eFUC4K;T?2Ie&ETb\1Mc^7&Y0#6]6
-QLGGVQ\Afb_(d(@7>L4.g.K\@3A?dV#/M>8ZJ9>3UT8YMU_/:55?^#cM;_cd#a9
/HNc\dPUGYRFY>B0=6=N2/(F9)_6]>#EVc:B+,7BG\1Q-Uf1LH\Sdf=GR75U@b>(
XEA));WYdPB-CX43[6B#E:I?cHg<9FM&W:H(>DC2b2FH+WCALd::gA_0ZD919X?G
9RH81)OfH@)DSebaA:;_UZZX)Q(3GI9:_1-[cbG?TJef?3P[:2g_.Xd3AACZ31G0
\YU,+ZC)ONJGDgXg?X.Q:Y,YDeQ6,<@Je]b9,XN1BbX3J#PY3?C9RJR5P)>@0Q;#
6<HZW=OK/H[-@0H-X:F<P0-AF)E&\4(]Z),HI9SdCbbdCY3VTVBD0eRQa9gHaH1d
]&Jc1L@Na?LIK_dP6/>?;G;.E5?&Z@b.7(g\:13K/HB6@NBTX_8aW:GJQWMM]UA_
@O^^B\)&e.],fKbfWZI18.H1;G(cLTGQBB@E#KY;f&XO)2BOFBd9PI#6]I>MYE\=
5DdP&YF?SY&[DA\Z7V-@L#PbTJ^aM^3+6E?4@WBDNBLe=#IY>/8Z2-KA+R/&fQ^U
6OGW(5XLG9:=A96<4]<AT+3HJc/.b_b^gWWOAW_AUI0^.BEKVL);F_Y-9Z994ScC
d,4GK+dFE@P9(7-9N+G],OM=ZQa7T8K73ScH(XKDSBF9;U=(A1AA,aC>@2<Ca(#G
^#Pc-8L)XG^J50bd#ag;Y7(-<MGf(,/XI\&6=M8#J+(F&1T,P?dFA.5<fg+f?:9S
B.W4ScP&HUL2B;/+^4>;??+>5CP,CVgUG^e1KQ@6\b^a,@#X(B7CaJS)GAfS<PEN
.U19&U:W9SQ+B#L&b=UcR[\U_(NfC/SF+(HTMO9+:b(_3/dPAS&G0-HZ=;IOaUTb
>3&g98-b1<feJSPeLKR;GO^)J&ZP?I[ZIA@C>_61dcQ=M4/MH:IcZLfIM.ZL:cI7
6(b,&b@eRNWA,^AOUR2[B_V\Z-RLD=8[1S<G+dC4-,HC@K/d\TJDPJUEgR<N6&cb
SfW&@Fb?0B-9LB=07X508O<,X.<a0>f_1AaEE^.S9^G);VVbK@;[T_Z.X?KGP,:T
LDP+LYd1-K[B55/BT=MJ++;)?]K>f[NY+TGZ9OKCZ@,[D:>JYBK]HKTN.dBIO(=H
gELNJ9-:W/e]RF.XIXSI7O.35B=#<->-P;Q^b&MZ<6O:_?IM_DE,IX(CPD\;UPZ@
IS:8b<IYKS4&IH)WYOBFVVcH?b#M)KM&eI5]D[[Z&KULNg;aEWbO)9:E-\\0a65S
IG4LGFJaOa71F=PFCCY7D6/[A5./#0Bd7b,0KcOW=M)0^7O9g(B)<fYU,D@7YAPe
Ic_=\bV@cW7VI5</R+AA0[EZE(D@dT\73beNP+XAIHfZYJeM2#AOJ94ACF1=f(5,
Z,&H;DHWYQ?56Q4:MagUFFC1OR2>(SSH.@Ga#YcdNcb3e6FdI^=)81@LOgN#QJ-?
RbaZf9&YE3.<:&3RJ==-@^GQH&1N=URK<RB?=b64,^&+F[Xb73.B18N0M_)8d)02
P^N@2NfRLNg1KE9@g6M1P=_Y-B.\V@a2cbMK93@NRaL^A&RI-XG,J#FBNZVYCSA4
>VG8BE#T[,TX68bWWc+;K4g@#_9X>4\[FF1<8CN,?CD+2g\,+,bIgNCTF=d?+:YU
1EFF#<Zf;GE(H4=6g/^DW:(3AIgIC@e[E_?BN<:@bSR;-+E(J8N&UB/,1R02S#Q?
@c.a)Ce=>f4\(+>;9HX>b0KAKW(O((;Ec?DAN:1PFP38E_Y0#&CQ9G<[bIgC6>#\
_dfJJI8R5.X5-V)=I9-2E(FZ]UB3(US<U^OU+VDR&@JTF=Z3b&LA4L=PN&-bJ1\C
SP9UZG;gF4W^NJ9)E&d2)X-OYG;1?U8+PT3S3HZ^O2CIQX/)QZVZ_5BO]&/[#AFT
Y[JW#>P0ZJ41dL3]6L0MF)80J184,;B&^H@_De/DWXWfY1=^Ff=OZfI/9UT&O/ZF
=_HQ7:2&^\gATD0H2_.g)fK:;T<)/P_:f1BB@03WG\a@8-R(CXZ7KHSQHa,Q8/c.
0_F<?9S_S:3X=Rf9Fe@S+6/GQ#T,;5.O08\Z?JCEZZA2,N:JH:5V]94CAVUbF\Nb
+<aX5T]]H-8LR)2/^?/e]_dY]ZZ]WX;[eMX.]L4KEI&\,1G?L]JQI=T2O&<YO-GK
VFBOAJg04FEABK#g??3bRR7&9T^SI7L><HXB&?HK1K??OGdLR<BFE-Q;&)O<UIG8
(7QQMK)<E>..TE;0,(+aW3IEO&:[Q@bBgDT0W0F..C>bIE^?;S0EEc75?JGS<EC@
M7M)JSNZdR[a;ACb)ab/7.Ke[;NQIG>V)F;g@dBNE4JDTA]]4BUN3F_EMY\gKf4>
LD_?fa2)-VGBJ&#O2)I-55BfU5FgEWcLeZ;(cS0;:@#=(]8RJG]Se?4NWON(4H\<
O(-><CSE\IW1VP7/,gf<Y/0BUbMRBEYc1abaYf)?5Qg@AV+(a5<U-/?;cS.\#2aF
9:N6-cOe?8\FaFfRGF2)6Q]+bfXee0fAWDe-g2V)[Q&3.OHZEPN7b7_H4bZ9W-,V
d+_+1-FH]5>ON(5(FHXETOGd@8?MRaRRZV;fS?U2HLM]I_2ECNF[FDc0G:7cgF2R
P?:)RC^+cM&,eD])7LQR??GN&?CUM5,dab]J]e,@IOC-0;DT>)Q4H4HUX&e@Y4d3
aY)/Ua:RP1c2&14fPa3@a[=[,RcRd7?O&.AUCTHdD4M?V=/9T]P:X6(MPaKXC1NH
fba@IC\cd[M)I5A[@0aYg-b/9<&4N1CQ=b31NQ+EVZ_d1\]T+@<_CNZAMLP,=28>
Q15S7Zd8gF(A2ENc&+2S0,\ZF>Y<=8V)D@(:YKIMg.J^LZUI?T_<(g[FL+;J,O>H
]5_@X)A0Z[3WUHN(O=I<1,;PWBbDa80,:=+;4^NA,cd?-#T^+#89gT)EC/.D[C5P
1AY@BO;?PH\&,WEE<OKH60TX9CM1UP+W?4NNF9Z8f)4+^3+(ObIPBH04SCe0cQK&
ID,cfNDbV(fEJa(G055_53D3X:^A7UY?MQIaT]AM^;I0&E&K4Z7b7-@C(#(W8e<7
4)W2CVD=,GTS+?F#&X(PJ3@-5V[^&NJJP4KU567G2RE3.7RVL8S.T15[X4XP\O_W
TV#5?@I+b/^U2QVWB^JdV81B6R59b\#&Ybg1AdZ4ZW-8IMdBb(G[IcJcUQ>?,=5c
O<g8_:.c;JQ3A-[f@0KW_^)KKV/Hc5(e+9X&1RHWdPYdT0,g=HI>PH00=0K4S0ZP
K<:WP19b:U2ZC9E)=U;N^GUd]\G5e[Q?F9gAa[7KaU+ggG/fJSUPISf?M.#ffINH
JV38/LQ97JZL)GB=G8LgO^/ZTW8E^1O9WLA68e4g]DaAc<Ea4M\#e:3c^1f6:7H,
@>U]cDO]b.RO)9WV&FTW1E#b8ORcZ8S:^CVQ5P=P2RAaFDD=5>BKTAX16[_O0f(1
eZQ0TT9+]b=f@E7<8CLBE,LaO5QH9,4<4BK&J3<WfMFe/_K8dSf2U5E]3B57IWHK
DWc1)BILEF>BTNBQ+FK4D4RZ<-AefN^Xe;W.?-D@>WcYeRaPTDZ2GD.Z@a:3UgWc
.d)/,RdgcD0MUP3J;B2_<:E.S[;[H=CR&K9b:,b&AV#\OU&.g2?=;QPCP@5ZL2(&
d<6I84@YC/Q\V_EP.g]5@a7-1dF7Q>.N(N#^Z_7U^69UUNgObgO,U<fc\^A098=D
07bY#N_[=4^6?>DHe:+?U.f#Z1Df>fDM9X?/aEC3cd0T+_-5;5gR^PeX+;?::O\=
A9=K>Hd@Y-K?F[HZQc?MS\OGAE,RB05^@,,;G(M(<b<>dRU-XJA-@cN9Ge#/LB/E
^&8PWDMbf-3E#YHV192+:]DdDaB7dNOHBQW47M.-5UR6CDe//=J1(6F,TG4Y?QE8
/ORWX48TN=L,_?KLADA<KO)PHKceP8b4cP(XU?\8=:8OQ.^fE&)]BJHG3@TISQWB
]g.10;e+,-#P.7+OYO+P1;T?gI<I62(PA?Uc=g3\FD->G1/3>6J2-c,[E?a5Pb:J
Y[?2.@=I#U+SQRf5c=ME_N.)OYETcd5<QU.GUI]\BL_-6WT7K4a4I0a0-GSR?THg
TUQMVP=(b-VP5^5#97[OgJJ6@IIR0g\ddH^U6PXGK(A=?fddc.CE^gCBd#6GVaP6
T?30eOY0e8G[5<gdXA52I\YAWB(5\+7-IWH(MT^#BKA_.N+:-gV>^J9E6L_DEM@G
+A_5(,/:<]WcS>I04+eGJgM=EATSD=/bH^G,,b,-IMAE(O.b?@^<YQe1a<VB5.aA
)cA014bda9IAe2FR#0GK_Y^Pf5LBL[H7^#b-C=B6PKAW+4d-ef]:98<,Q2EVdU,0
3PEU124MbI[/VQFB&JFN/A3^cUVT0&HUQ5cTG?@a<0)^]c][/?P52B^aOE6TEFR.
^WNT?GC+(5cYU&>6cZ6AHZ^5]^PE953c3/\?ES8HDF>H?\UY;,EX46>5b?1TaJKG
B.6[S=8RG:2WV5.9Zd/+deSD<154N@c5,EB#\b&G#XVEWM<1\K,Uf@1>6^fRNS5_
XbAHd>3gK&PW:cY9QP<Zb@7Z23HXe7d.7CHfV#F9C4<Gc2:,@Q<g(CE/LB#\Z.c]
B-L>)E3AJ<>BeEEPTG)fF])Ca/d3YK]d:]TZG&&LQ7N.76@fGSQf>T4T&a>#,X-b
.8L,aP5[GaGb[X7\bc[CHaP.6;QHdC4RYS(Q4;2EZX_/Y@]VfKP5e_-LX>_G/Lfd
SgZJO6d<EaDRNF)da_@\7T3XJXbY8UPR=0a^+?d?f.[F2])4X#\Y/2-6DQ1-G(;,
gVPg44=-43VJD5be&YW7M+:7S-Y1+;02&K/)f)e:9R;d^_IcJIMaVVL_[aG>.;P>
+JQAH<YEJdN\B^]3IX[=XM<_V=O>bA(INF:)LJ5@gHf=(JGdEWe9-ZQ@6Ze>2(U8
LK<PZXK084W7#e\@L2dFa&&<:\]].RIgAg.O2c,fOV5>H.g+@-0Jg<K/_I1=g@Bd
UK0NQ^LS;eVDdW/VZW3SgUC]U#3MD\6W99H837&077-\KY_0)W8c3b2<^77+KN/d
MVO#;9F22_6Y7C91]MOM?fI-dILR<@=FKIRS+C&9IGEIHbY_XV0g+?A\(&7)HgIY
,^XQRd0a&+URT_Y69NXfHL&:<5[:OV,]eO0c.c]YFNFZaUKN/T/LJ&,0O(>X[-,O
GbJf4>Z7-R-_aeW0+(6(aR2,Rb[Zb/NQ/K6JcAdZ-cUZ7RU>fR,LOYAe7eeK.<Z&
S=#2#+;\CD0EW(7D71^0Yf,^DgfHSR2^GS^Z:FZGBUS_;7V?EM(eBQ3_<^d&ZBWJ
W2M)V]N@=)[&HB]CQH@9&XV8DZ>WP_Z4E^;0:\KXG=6\DLZ.G7E\X(be]bA\2]P2
dE]N47X)R@#g2Md7)0Hdd1GOGf467CY0^6K6<^V=ED#_EAX#f71]L1?HEeGA2BPQ
MP53\];Ae3fOI\W5YY]-;&Ga&GVI6RbaT3R3eabA[+--3b7I64DXLX-?e)<O];D+
eD9b4,ZZ2;?b/Wf[B[b[;cDG?-W^,UU,78?UKQT9dZ]fQ@&P:B7/4\SR0<SBOWb:
T&7/.O&IWK3-^._6U70E^,W;:9PT@<G:c9_Qf;-4CLP:fd\DGNa_&5-F^fgNM^N3
#@d0?\fcaBI6BI=XYdF?SEARD#AN+OcYAU+_9YAgf?B9b-?1d3,]1H/_V7fTX2:g
_&Q(8IS/8W9e_)@K1^>NCZO+B&,=:a\DG.I#6&EL.#+PF(>F)61BP+5+5HR971S#
NB3J<JW(c[0UVgPG04_+_9S93W2WWHW8;fXG2:?JQPA.UO2dJ&gZ:&ONFH](?>Xf
B(#.I[]VRGR;+UXGDQ6,dO59b/e\Q(,EfQgJ+g6Z@Z3-FUF=LNZ/+::EBBYNF(PS
;/bYZ-Y)fcU>]7N(&2ZWZDYRK+e)_&+)UE.\VdY&RbV8CFM94Z^b3-VXCH;:B6&1
L0R7Lf:?W^b;/515NcODIO^O-5ZUS.S4>f@>G9ENeAbUYeU7@Xe[/@VDG_T&20H\
>9d5#2P&(6=4T=:\SNS23=dS+.[=35HFJbQY2=2;dX4_Z2NO5f>:10U2M>D(1T;A
#K,@B/,<WDg>e&:Wc<T/?[c^:YAUIW0?SA56=I4T3cbWFBRW+d.J\VKN-2IJJACd
1&GUL15L]AI5/cM-IO[]N63WW8])=7(a9G3eC]T958CK?c:3A]=.;&#;=/JWFf5F
7?&?F/aCdY\Xa@QWSCJ\5K&?MF^D1;39O7D7/REA?:S1:-gH\16IG-,E\]e+-Y8V
D&&R&1[E.A&>eg=F5,O+2OaP+YJU-S(^>LWF:)CF70)7C,YPGC+g78aGQZ_#VN^b
DQ;Q\AcJ77X0ONCA;[^FK03<.FQUQ>XLEO5NV,Od&<)78]EMPQTW[HOF#GDMTP7T
:>Q,5NM&0b-K<-X>O?6J1Z1[3EW^T(IJI4(#E/K(7>TeFT>1e5RfT3.8eAQ.UL3C
+(K-H89O>-RTQ#VVI\#&A;:?:;O0>?>6&HHVKTR49f-dBZdO\#78Q.:MOV[ga1,J
(4/e\-X(.(_cY=2OR85XI5],9-A^<2&HXG)g)C@=W&c=8dE;N3\H7_OIK0>=gSZY
F5ZS8Y-?X/bV.e5)YZbF\&E+M4+C_8(:RP8eN(IX:b:(U?WI61762dB:]6MARKd5
@e,64XIO5])@D,^_G5-]#^\<2^6D4>eUc[b@/_DL:4b.@:-&K5,9&Qf+J9PK9EHD
EA875WfWQSVMZPQa/f#3?)<IYCaK6Q^/_OSQM\ML;1G:-J#CV,FL<OR;[COJ&DA>
XO/<6HEI5A1.6e:RNd./I6Gb<WQ<5U4dERML1BH01g22)RdPF)TB3g6\<Sg,O/(W
G[aYN0d/f<PRFK@@^:\XG3+[\4RPZd51O\1??F5Z&YT\1O^D.D]a.W<25M?K3=L-
6S>c7)2/XE,e_/0##TK2,5G5Ac=Uge<]_1+2aM0Z(ZI,g_dZ#D&:c#^HcRZ<cKCc
gb_IUV=e.EUA6)40;R8-dI2]J^H^&gZD7OMZ.E8DgDY3+:g_.ATZ(23HIJ_GB6M>
^/TAE-GGU;H;?<^QV.d33[)#-KR-Vf>EJaE;6ZV(EE4,OY6V^.3QfAZc0NUbfS;;
;QJ@g=UNf8=(VJbPSO2bVDOW,#J+eI]AH8Z=6TCLI.T:+SB5\GZ+7M(WC:J\ZJeE
dVGQ-9c80IZ@Z+OGQL4^A?g>bd+;^_>NG;Oc5Q;Uea:/4VDg-MBQ8E?0Me\9^M_c
,-7^3:U5KO/F2^3A0D&Q>Yb:6:MZR+?Y6=JG]Gb6(N/AMa#ZAR4YCEdCcECKN-+W
cf>B?V;f7VScGf0T39c1,d(QGe=MeaYK:9,deP5Mb])>c@+gaZS<Ua=@Z?^b)g3A
(PW:B._53a2fe?-R+1VO6.U7&ZKOIN_FCK;5A_[&_4>0c4@M^]>./a/OgROPg>\L
bge9-]JT7d+0+U=fX&@Tc1_M;c7KSBMPY7JTZ_6K)?YQJH+#RM\.SVHB-CdJZ-=9
<D4H?d6P+>WcD4g#-EMU/>Q/;aa=F,LYReDMBbC6e:LJ_AU-#POJUX(XL7@2IYed
a#(A]HXd4/aIA;<V=JKSaV(WJYW8d?B^G4Sb0I66?NID\TRfGCB_+O]40Pe<JfGb
<>ZR4#,[Oe[K2N@S;PF2FcUX;NM/Z+5RKGLaeV>UAH2_PON6OG[\dZP&/^OFBP4-
N[7@;Y-:.V9DB6=WSY]B)?3.8A[+#TL;I_]C@HHGJ+QUg3W>5</)1=7[<CDZ-SSN
X-]Y6Hd.(45c2,Rd\JV3Rc(cEQ/fODW-CJ0[MNX=_XBgQa^NQN1C0YP>>F1FLb>;
OL5@:UX4T\.1BYE:>Md82=R<)0O]YBT]&S?\=MQ7/A00ZK6(N=2,b@+K5dcRX&FJ
1]+UYVSWY<LcIX<D?f8;<+U.2KD+EYbeOdb&2.6c9YbZ)aST>=(V@\UaR(TVL8[6
TL;)7KY.aFfYVV^dH[_Fa\C(I/Rg?_)]G:+QOG/HJL^/FA5X70G\G2604B7K5[fg
1_)74ETSZg4f2?EfeEZ)LS/>C72)2NA9DQe6=?36:6(4dEf5?<5=/eSbe5dF&gHI
C=)?)YZ_Z,;,d/Z^5H:d;P(<I&cQU5&fN<;EAd/gE_1@VHC2YA[LfT)bG^:..BCN
X;7R=f:A72(FV,>?eacKW\L/Pf2\g]1E-Z^L\H9dMJ7[5WW0BCO8DQ6[_^T.5Zf5
Qg7[B:fZ<3-3DN)4^_,d)gO.&]AUad8=BH(18DWC00HTX<=<HIYee?]_SQ4D8UZ5
NQOOL>)aP1Z?5](=8a+53>->6Bcb/#+0g-5cXL<JLR,\.b]GSD@5L#X2TOXKSeW9
Ad]O[HMI4Q8W[2J<9#^dB-NGX,J4A2FRK:MR[Pac>9cK^BII@fc=]@0Ne//11V>+
V,fVJ9-36Y/YZ>U)\MJT:_c3#baF)5JNJBMFMI\/c-=&FcBbc?FGQGIQOXCSDcI<
_<e,\)]]JNY]3M@G,84R;gM3CS.X.eU4X<5@,feX\1QcAd//I@I^5,NBd:c?+-_I
fNDXbPU.@F]2^<GQS\?K(@TVAHM?K<T#V<VM)b5JJQCeU&W&7U:?dZQ?RZ>-K&bG
DZNJF9;T=eAf#)22Vd(HgL>NcGAU4<_+A)37R@+R8PeU,-1/=9,^5KOKPAN>QL4G
?;-02Ve#)>4:8R>_6@D[&)T8+a1cA&O/WB>1^1,OU2g_DM@<Q7Q)<5e5R>\=)c-L
2J=3.0MK4Uc6]>#eJ;LCg5a=)76()9+PE=ZSeI>^#=</YgM.ASJUH#-J_XUY8K[1
OWX&55_gZ\E0N,X@[5#B\931EEGZc^^@1X;PF;KP<OK4G3d]d0VL_AG)(.:26P?a
&C0A?DL-XUGQL@(R<D(a5OI8>ZM(V5[C.T]+:[FAL\8/9N?MX[>S::dWXcQ)0ZZ&
&&7_\[1Pe+P]^VdfgQ0gY\MbT+KeR0RW>VO;2V^PY^.LNMX4D.6aDTeY2X.5S+aP
Yc09=04-QV>^_#aAaAS)C<7YdFM=W,8_AK.(=3<f+^^UA[4&,6,(]C]e\\AN4Z\b
M.)6TaU5?DZ4/-QHTA(S\1a8LD]+E4=&8GaMN1ORTBSObH_<6a/MB,FV-+NETNNN
V);PIVBAE5bZMc=+FL.EZLDAJ4fH==I1VG/bXH?a>TUIJ)YQ,DOSc#I28>WR<25>
T54N#DA9UU5EQ&:&PYGI3Q^&:W5<IUT3J\aaNf..W(&?B\:_E:YJ4e.X3RY1X^MC
EgS#0TX#D/SNY_SOTV&^c0/(a,Ya]\OX8_Y>3^M\4fB/2G:.>R:K+,])bfB_3cb&
>3H@c\VU11PGf/DB#fSW7PQL2JAdA+.<SS[4A)W3TTYUHVNO]&M\]\(3a=XOOEY@
C-B2g2DLR2H?6+R\W3aES^8I)K8Na#1@<AO/+JNYG<NQ3/9:gK_O-,EbKKa9b0<[
g]9YIGbHH[4&cg6;=B=,;YY3DQ]L/5agE.\D#J;B[Y,&)IBR9BgeTCOGRO#/RIcP
]N),7EN]#H457GNZR9,bA98b5bM&DaM7eQ))T/C>I&)+7-BaVNNc8cccFgLFHIX&
W:XUDVad<XGV6@C&8G5^YXGA<RH2T^TOQ99UTbc4ONb=1C59_:M@T=;bfQ4+6DHT
I.6^YS9+,KVD8b;7QeHMV563\N9^d8b:a08JO_#/KHQ83;D2(1?7(>Xa;UfX,Gfa
,N3:L615:b(c-gcJcbb^L.ESBBYVe@[>b_5JOFfA;YbcR-;-\02+8^[O_\&7D,O3
B?(Ng?&U(T)1XTaC:O/,2b9c;TBP@ELX)Tg5BEOZ[J]OMI^WbEEP>EM.6KdVUR4]
R<^9F,BUb+f5V(C^.);fY^<YAQL>>N+W3+T?)5+eeM,O0I40\SDR&bRPVC)C@g5:
_.^fPL[9)<HcZ(,IHOg@8aI>3C<MG_A[;3;7F1B68F<>?3//H9]^;+\GeMKeP-(B
7@@-UIAVE#8f([4/]5Z.=A65ST(Cc1RN\]@W)/c5QO2-f6]O:PJO6RZKK0@7O^fa
1cF]1d:\f7V&g(&)+#GH?&&[;8BTbd(OE&dLF8Y>_6KL>YDJ?Y+ES2EC>7AN5Ag]
4c41KfZG3P>^R&PFZ3fZ67[eHO^I6@_(TI+GIaTQAg^^_c-a5GB#KAC_WeWM>)8@
DT+JS5_7JE7NJAMZBPP;CKAGK/2D:<;M3cJAI.;46bL6TBZD]#/+;3,5NU;UXAR]
L\=8g?3/XTK#G1UdVZS92Oa\TMdEaT(F;f;[<AWI?ccCLN.76G2]SJ&[@d</AF_2
?2gT<KD=TE9Z0/;7FMQ.G^)KLd-)I/3S;TUIge8.f[-5dE0KZ2MH)8.E-HS^8GZK
#5>RU3HOR,]:/A@^g):(.COgR9:Q/a+KEaY]gB<M#1XR?f#e/^U&g>&QaZIJ.\C-
\.#b:_OW8_8@P#OA<@.?4Hg?,3#d)b,PU-B;JO^W.NDVNdA?0cB7RU2eEN[BgWHO
HJA\=5I8.cV;2;HB0H5+7W@8:6UM:OMSbfC3;35\.&4@ISRNgM[E=1F#J&:Z7(+Y
4R4b&ZC>N/O?c;LQ4Q7[2+MPTPUc7^^\Z9RF?>U06)#+G_E7:ab/F:5QW+7(TXON
_TAJOSPX;0T7WC:HV8#Nb/>IB29Q]PI8&BLU\=B,VEcT=8X:4d]Ya^LV_RQZ3CM,
N0\b0(TD^,Y_D3S35.Nd])e6TcIeXbf0,W;17[II67?7PYCe.HR+GO:EJHaQ:Q1A
M^@EFAd/6.KQa@_DB@N<9/3IE/ACYOcMU[XcT]+aLN93Y=f=54Be9<<>)U]-/I=^
(P?c;;D\,M1W3bQa-2DaC8)H9DMaZ_[7^)7^6T9BZ<)^HA.BMaE0V2-BHZ0,O6WC
I@I4=e7g..\H/>IK?;T+JaV1gG8J:f.P44.^3H^Ib^@,QD.T\:#E^-93+HU+(YKM
EaTWd#.[N4N<,CR)bQ>DT27.S3]E7498UG5b>P&IDY4>Aa+;9Fc(O<\R_AgD\c5d
5>>?94BBE.=-#IL4/U>1?CeOLQd2=JKJe?Fbf4S[0e0Mg?N]E.CT:LBMHNeE)CH]
.2CQd2A@+JRf+^.H[+QV>[W^>^PL;YKAP0<feF8:11VDA;P/<E:C^EV0PF\cYb]+
G=_(B372cede4RVMI,gOe6GWRVgPHG4_Ie&M\,CN)K2=F;.WUge#IWbSb6\GfJ\V
9V6E/5OO3=1R]68ZX).,V>]A<9:O]Y4Md&gKWR=.>15[HD#S)&.NgP<)64;0G2fC
=5<],b6USZ<S5.,a#]:^5.J1?J>=)1,,5[&Y=:Nf>&6#e5DLa3PHT);=]8X[T;We
dWB]O,1O,9^2aB,@7L[KYM2)bVZ3bgD)1]gbBNNQf=QZ3</(1ENJT:Z?QV?49)MI
<TVa+>;K@U<VeCgE0Z0@K@2WJQ(5MdccYZN-)2PS/O(8AJG;d><@a/]DK&#@HPW/
LL4dbQ5L#,BB+Oa\d^SRc+4?]H?Z-@,TTT]#2@5M:RX5=QePcJA<2^a1F18]Ld99
O2,9AV5Ke0D?L?(ZE3#W\@EbI#F(9YQY):ZT(EHeFY0WG^9R)A@MeOC,<:b#KGP:
7:gN2e?GfgD-b+:1V?fY7@UR0-5a9BD&GMe=NddPIY#JJ8+@B:#2Zd/1P<9K)6N:
/eC>8>bf5+<:J;XQ#VOZHT+[#AUN?a_N)UF0A6X^LL7B>=ZV+a&f[:fAOA/R(#VS
3aEI-f;DN]LE4]_-[XM@\7NX@^A[NGaSBSB8D1O.-.;Lc;HXNLDQP9O/.GQX)PSL
2F@7g5_ZIGA2IM<C9JZ=cF>EcLAZP4U:3N6^]04P(a9BT?71@[(FXe(:c>AGJU6O
RfbNc]?)(B[&[@KKa]@5VIaV@B[M<.?DZH=[-8B/VF.b@#HVMMRA0QK)^^6,U<Of
.3d4RYBbTcV4,>JbN?-&F@424M&#(>TTK-L9#X^LQ++VfD6,CfJK^[c&QV[.&6RK
.N@/?BNe[R:1:TBWE6cZG0WSB-:ecYd,DD^+.a]fbaB?13)@SK@&KaQgG@0;MJNa
>ITb[b0,7G8=NMM?c^dDFGf.c>:XRH\O(]0&eZM>KL_IgR6/>)IH)+[77?cTV,_^
7#\=e,24BO&E0<&)23IHbL2D2L5:#;GbF.Ebca>_A[dHW0+ZG^X#SZB2>WT=77:-
b:>>\I,BbBCT)LMZ[HW^?\Fc.;UEd<c5MCBB59.d[a23YHU]U<0]J22J_#.?:(;W
95?X5-J4d-7RgAINC@^#CeET79gRd_]OgKP12)_+Qf:,+UKT<bR87=3g#B9QE)-4
.:5>[;-)7KZKL)TK#7M(^.@PN7+A,(6a9;)6NZd+=/2HV#fUfT),^.F.^CG</L8P
?\@aH9g;:LYL/YdJ#Z\@A+1G=:8EeRffMQ.++LcGB9E49B#&EYE[5U@2^/BZG5ZV
dZL@VK.6QcU6K9[O&N7P#PbQV1Da?LOb:#9?af<O-bFUDQUd2e.7+.AXbeg5NCQN
eMbBX0Ie-RHB5K.=?>R+1EUXR+-IaWS1/Df_bQ+?S8g9CUERNPBAg6M.#2#2Q4<6
HGS0>QH-Y2T-6]KDVdZ@HeYX<-F4DEWRH:2GWE0.<-daR1>8d?1+b.^>,LODRD8P
V?dZ8dd?I[[Vb>_+a@(64;H?4M/_3fK\ICOc1YNJDJ2cW=_5THBQEOK2fYFR]/(b
JRRP:U(>LA0ULV2.aQI_:aDQQ+EF)aL@<bA5DBI>>27Z-TB;:^ZW^(&130ce<eYe
/GYFE9KD&2F@c(M[cEE[4033f<(Id&3X,HBAZX;P(I^&(OH4?FXOS)N),Od?dA55
YKR23TU)8JYVH[N\X=(QGMQdZ9)S8\7;7/==L7AT-\V_Z5UgDgZOF/-++g3OSZ+V
BZ1J[5TDQS8>L9E;KUNX;OZ()X^W3Y25ZF;J-R2M37+A.S@12[DW>K4C8R46.GaN
DTR^W[W_,SW&c9U9@eE1=6E#KOM89Z=Z(ea?YXc?C6MN.O+)&,?HZQ2ZK&EZ2KH.
41D1cNRD.=8&_ORN9e.fM+:WDO1a1K/OSIJKYZRD6#U#Gc><Nd7g?J=16.0L2c?H
#.U-:&)MU15)K4XT.fG9>BST[&C&]cP3R95J)JO45c;=(;F\C6#U5>HEV:T^MYW1
a@^]=:X??0OL97c(V2[^NK#L&M-)FZ?S(H=+PL6@#e6#F:TX6ZJce@6G9=67&35W
1@2&53T[C8b8\g-Hd_SZ1PV/^(=(XI./P#-c+AOL/79XbF^6dF_NVUN7BQ=&3;#J
V3BT3JH9/.,0;Vc[10B0GF&1UP,\U6UR;XTDfR1+GU2RR;+_GM<M2e>/9aMEE7C2
b4=/_H\6X:LY(BN8_[A2EPUc@R>c/0:+5O?4\R^aL6RBA][cQ;=(NP:A>cRQ.1H)
\Hb#1f2a.+I^+79d9FBIV#VC:F3_[;/Eb]XO^#=.W)C?9-?+2FaM;<?X.&fCPZUT
O(R#24H[cAL4-PN,FFBF>;3e8B5[CJLOGOR2P,cdK3JOM\bd,bFg3[74,@a@XI\@
D+a6<aS>^#N0M#C1(?^^VWVCaSB8)9gQ(_(0_fYB=GYV4+9S,[A3gbB@fL>Z^GFf
Z2QWM,S8=IFTM-bU;R61T6G.KdCXAaV,N_=;(?B\1[aV;#JFO_)W\Z-TU,M9@F]=
3H/UIB<8_BZK8dUK2V#/E8#-a>gT0K,<M)YC]+9FQgU+@?_PXMR-(0Zf]L6B<55L
6WO=I8@^TCcHR^g[f9bTKC4&HT?9&WZB=6B:b[F>D09SP/)>A<0^#Se4gLIgBK#7
e/4&0(:MFWY3E75I/PU>\&8.=?MHQYR7H78X&a\J:TWb+NZ,?RV96PK>.QGDNZb)
:??SA()g>1@WKHg^QGM2OR5Naac5TI(2@V?gVO+(/F=D:QKbc22#3cb/YB@45MVJ
b7b&U)gE)G8\JR:PQP\9G?#4[c1VaKgU[1c.]Q#.0I<D#Y66YK8HNSCdZS]b#E:6
/YM_5X6a:Vf6R_49]693Kc6cJ-?>:6VKZSeF3a=4\]7e?6FM&c>D:[)>&GVNW+:W
)<#,O6<W2cHLI]S^_8aMc_f1PFMH\KVUJR+G^+E:RDYU#FVa:9:.B/b9ZAE:=:#X
_IH8P6:Eb1EZ@+_dKC?5)FI_M]X.,[^03\ebgeNWYN3LKQ,9D:_bF6).N0Bb6:Df
A(R5gSSO7CLDc,X/9.eU;c^\UKIa^f+PcfTFX)).QX#>XQE(\_6BEcJVB2Sbf+H>
\NVZY@A@PT<C-=120CKI6=[F:UTFX]2^>Z26&:KJ^;#-F=692P^OII(\cUL.]:,?
3Yf^2(6OZfDeF#@\:R]H-6gE=#?QFR#)Yf5><IR(:1C2:X9&?EJ._@G;.:fIM#AD
Nd4:890C^;RSABI-C33^/NKXR=0/CP5Zc:]dJ6IUg4++(gR#,]I)7ZO4C0e?fW+4
4HZOGgI#>[>Z)\T<Q;9:f.M:2AN>;7@3,H;>?1#U&e#>WX^C/cS[+-7XYD#g0-[Y
XQYRLS?.;G6][Z0?N&&GZa(J+)F]1GcK7egPLE6XG+3[4J]c>DJ0SNdb#fZ_a[MM
YXTcd8HC=:IWD/87B^WeZc:fI&9H6c-W7C,PTdTfY;\0d)0,LeO7_H<#2gKR4XF;
)[.N5_8[4F7ba4O#,R<U^P32cG_T7SAdSV@FD[L&\<D.gTZDfYKH0A-\49U8gH\I
ZQT)c^W63CA5N7JL)Z4XYLRV@[S>2f<#bb/3;9(TQ3?AAN\<Cb77:7RDVCaF^f],
.+EPeC+Uf5Y5=4&.D=BH&:9XE5R97gFb?_QI6O3O?E.a?<gN4^E4SaM)8C-4+6NT
Ce[+0E4e&OK0V:.X)U7GKeW0C(@E53&R22((XU:VgJCH9VJJa&33b\,4FKHW0@YO
[ET.?-N=BcdI+)0OE.#R5P>BK/39H&;,R<#CISGV(:&3NAM3_K)B8MWef,SWCCa=
_IV&Je8T-MEY_L#>S?F_Z/^C<2?MY^^RM3BFVd3X\2M?:QGN_,dA&PI4\LSGH,)+
[OWTG1VC2T#f,L5A0<+O]^)N][UA&5A]AGbD?J(]H#KA=P/)CbV6<#TWFRIg[)aM
XVDO:]IV87IR3(2FBCg9?=<GI/e;&=2.c3A4G:2T9?S>6@)fN1^EC[,2\OIGI6bJ
/ZW6]GZKYCeY/X/(f(2_7C@d5/8eNfLSSg]K:F_.]KdU>[?0)C_<,A,SDSTSEZQT
cUF@^Pg7)Ac=.5_<Gb^#gCB+>UgH:<3<3XSRZ0-M\:5Nb_E[F4194Mf2N.?:;JP=
E?R^7JCWNS[0_<?]JVg)(_IT9EP4RDAKcW;VE;OUI+Ec2)MJJb?X?a#;VJ+#>G?:
6+AcB^gaQ[OLV595H90P4<N;IO+b1U4#Me\/_U[8LDgM_X+9]#_+Lc/CK04<VM[e
B8HE6e^1d=+>A5>YQC9Q@dJ#X.0V>6RQX^;JF;^LeC@4V_;2e0F<8I16>:RaQE+V
\L<^AI5QHBYd>HH;LFe.9:DOgK8=__D:UeY1@/TCYMa]MQB8MQN:<@+PFeD,9b?5
GFT?\W-L:V?\C<V_K]^V&\OcUY\[e+=\#<P(#519/^8#_,)QV<+EJ7QZL@+.N,E2
;f0HTg^4_5>)4\D8:c+K6KWf,g4SU65>3agW@=.&g6dN;+_D24[HHH82dcI5&5/S
dRB<XN,&g=4F9NLOeM#>]-IWNW6_@g(\9?JL&ZN/K]<AgNV[KW#N#+fW+KYZbESf
^Q4:+@M2K[698Q+Jd/I)P)?2ZbSP82]ZVT#9>06A-+2Bd9^YNGZJ4H>C;P^g(X[O
4dHB&N_Ia5(bYMJ8,[W.CaFE.OaV:.;Tc9-Ic2Q;gM&?PC?LALc1UdJZ9g6f@a#I
_6K<@a&3^^S15f-DUTD>]9EN6g>ZI+EN#&[5KA>fbd;<;5M7#50SCQK)FL?b&@R,
O..REK3XeL50D@:?8?T?[f<V3;3@>HLXQcMLg]OO<^9SHfGF&2-edb1NR9E#VLB0
O4U2--DN4CY3)Z)=E?^=dcLSf;(^_/f(AX^I=:J7gTZPK<aCcIH@O[U905>?d)M\
>6^T3RZ9aHYJ.YG933A/#1?I)[-@)Y+=f&EA_MEQ@X)E/Se,aGQ.e^&]NMS,eB)c
(:3X3<93TDYcFF13L+GT6YQ8K^R,45.35([++L6)8)SYQI;#Q9A]+/Ag0_-]3.H1
FDSUV9C[X9L6,EP7=bLX]T38/?/T^3U3GQ_]]K3U>b<7,(bM6+fH20_<d^UG0O6e
edD?cKW.\7C,E#[D#FUT^^LaO\_NS-)_S+8UM\(#THDDKWFbO6Z6O\4GCSVFM32]
ON--=[]I<0@<\-1>O.X9:ef.,cgVEL,W?W_76=//e,C>._.KH6Q[_\6IWV?</ZF^
)5Wbf-82;<6FG)NFZ:g:K6aOZU0AENf,.\@DNXA2[,f7(QO-LUVK;U\_F2RL?XVD
Ke8D2QJ>Z19P[5]+fg&(\a=SN&8XTF=[cY<gW;D@gU.IRJ#BR/YG1\Wb.<QM1+DD
O[3ee+L_Pd.1OC6E;1M7#/S<?SK>II50MAGCJI72[[[^^LK&:9O^>eLKAHT_Aa@T
^9\AR4HIJE3Y]?U/G-BFgGbZ5_fg4_bd-GfgASQ2DCN[@CG/JcURS/eUb+=PIXbW
MA?+SW3IIJY@7QCP,bX&c70RXgcg\@P:9=L;^#D4;Y__<G3(2J69=aV@XJM>D_T4
g.Wf4CQ5QFK1.FX77WI5QOJ6f+B_DD3]MQ[^73&be#JM=KdRXUB]CB+5Lf1S(S5A
\>][O0c81^A5;KDJ_#dg]+e>PSKV0,GAB7_^5CaEQM.E5_=Q-?;RN<=;K5KPa,;K
[39-gZ>a(;e@)Y2eD,0LND1Z55H.3<Z1&cLB,,+G7(NVJ^HEff1_^[#A4GY0.U;O
UQ?8?:E\2\L6.3+UNU^)1Y/9&EdK0aK\+H_<90NP<::O^MDb-?1\3C?F12)gX=O]
[HAD/b)f#Ib=T4.c4[8TT_HFHL;HD1<R;,HRHJ^E2)_5T,J<@S\C>M0AUM=b;-e(
=&PQ>DHfH>;:&5052b/9>[fbcY71PQTdP+ZPGS/c[)7I_6@(A_&\_^&S_DGXAP\R
WHO;][SH?O1-_WK@WIW7L>W<>&F6[2X.b9&J:&FA_@W/<55>@1_SD@NZ+Ie1+MUT
M\,X-3G4-\>+?TLcO?RG&68?,).1C1d)MZ\Oe:2Y=/Y=L@3e6PLJUF#=Z\PWfUPf
]]VM@,>gcB<ED2N475=WWKTe1fZJ^R+D;VOW3g>HPB8&dJMJ;=8H[2BD\dY,,U^K
OUM>E<f@F\J],P(R=.&>b2aD)L1<B2I>S6,D9>[TIOK5ffLZ<b2KL25=,3JeG;/3
@GgPe)^0)g)5U]PJ.U154,[<)6Jf<TS/F:6FE;4;K,_L9,DGH#DQ)XWQHCGY#H.d
]1]38Y-JEV?JWfK\+)NM-dS=2JE2.W<4L4/gL2=Kb4cfdcRVH?D++\RGEGO,MZ@O
]&+(BM(N09cJH3//YX@R9ZU.;G:B6]7,X/_,[<=fJ@W0/\LRJ7#+?:,U#^EL493:
_],H\HaeH_:LM<(b?eR)L16:OO<WDIcZ8)[A<_Gc@9NO559K?,)d_6F[I_6]@(+g
eE.49\AF=)9W&B](O8JK>_OLaD=IMA[3+04@/J<7AQe@Z2@TeYAUYeY,-=[f,.NM
@0/I/LG297RRO2=KgXJU:gFJ)DB^3f].=P0,(@TbPH84A+DdEIH81W<WE8+-X_aD
Ib+MYY-5f^#.U=Ba+V2-Jd5?J(6VD_<-&9:4c-CJH[gZDFO>5fdc@.Y#W<SM..+c
&\S8DS-785>3GA>53D)JZa.LSd<Da2K=C6M8D054g-dR^@1T^[eUfHe@L/3BR</0
8Y+Ue<]>AQDDeXK<gd6dT[;:Zd=U=N_ea.1&_DBUWOT\>HU<K0/8;=\4C^@U,15I
4N.[S2)PA\1bQfdZbDLIL=f\C?DRI_<O:/T;A;c6=ZWQ=H:8934X3H0(5d^CB1U?
)7\8PFb_8#NL,^D/IS_NX/Q5:#H^,@1gc4R6/G:bb6V_aS9+6M1Ff?P]KXS3a-9Q
/R?G;aE:PeA.U&EdT1ZI#=\WJfeJP5Zd^>MWOTERcQ1LC_M[V,0J)5/bDFZ,)^^\
^Pb^Va[;5/CBKA:\I8>24HB(Q,]Q8>3SVg]_9S#dEUIZ3P-KY-2)AgN,PMB>c63S
3B4KVRM>H[e=D/(?cZ/d_52=Uc,XY/RMA&cDEF2(=K^<f,[^YJ1F-(MdS8GH08[N
2T+a7?&H.9+OTOIIREPRNY:+(D.BXa9ZK-GVTJY#:V]dU9:1ZO8E/7=97+0B:#b[
0GH59Y.4b>RGO?68A(A=KP&MgRd8^H>?88K&=55&,P?S7b+Q;??0WZJ_M/=g_=[F
XSdGG3XBfQ4THM^,#HOV(G3ccSCQAbO0^aN[GbaCDL&J//8EYLDY0c(3-PSB(E,&
?OHa@;.T67\0J.#+CQ,bOP++:=]0HTA<#XDS;FF/L8(40/73C^S]E^RF@eMC@BG>
-8_D/WA()./IA-8CS(ELPT^CO/:U-7PG#G-5UZ1GG\6:@FgE6abceSgXFd><T@B(
RL+10M6<3#M4;(TdS;5S>/59+Q5Q40d^DUAfe+GaYFH39K=[ca_b],D/5CH5<1d3
fWBF6^FfX@80)Z5G&;=ES2M,VcT3NdcM0P5L2JX^I,;BeF&QQ#9MXGH:EB<^Ha#+
)>;bGZ(HS=WY=Q^(8_]K97SeX2;P8CPG\CSLD1,;=e_;,B7[EF#5,TdFg]_0PVQZ
EU88DS#bSCfg961C7/X7+BJ-g/,YH61:V/UW#1ZMX)7fY8#8GE\5BR/:=4,Z_B/^
H\94;ER>Z9?/VY;R^&WVRS8#:)B&\b\83<.B,ADF90G1(7,AeLH5SV./Ie2?eMR9
f9^]VT5RgVZ;54=Z#MF+a,]&1E;>X2RIW8Fb-47??X4O0Y)U&PAPI_>8Ha<+/4L/
3/]E)7GN#;>?]YAL<K/cBMgVVFg8McTb]e\I]IB?8)E1A_RNMf;VSQd4b_cedP@@
5L^YNbC(NN(_E&K4cUU36WF/BR9;R_ab+0\Nd9L4.]UR4#5J(SCO5=[/()AU1]&g
AB>&4,4X/@DE6U2@:e_/O[FCbS?(5^\U<X^eB</BR7O.4PZOVXQ-4XIcc>>8@G2g
#V.&a]G1Uc@cI[AUb2Z/@WY=C0J#0ge(a2@M1[1+DdV)]P6gC[7_8H/fUNES>3?5
TEbTX0UA:d_aS<>9T<;R;-(HQTWOSQg#bWC5W0G?DaT1>8Y[FX7?2]/bW\E3LK?I
I.NNX;UJ6ZA7gVCXA-5PI^K9Y4D0@I^E&f^VMVe0QP\:?.aZ,W=P/88^:W]G[4HI
7S-:YZIR8Vg)dca^^J8O@L3Z-/cLG@Pg,1?C.J_RZC9\.76Y5@Q^YU4.dC-W3N?B
fb&IWIe+P8N.-[14RPF>0VX)4#>G59@(IQBMa#>+Z)8cA\Q=Q_IPO0V8\KJFK-W:
>SI>Y1#/8.?EP@GXW0Oa(e[<T^2(acQIT<a\OgL/,L-WcbLJ;?>PF+N0XJN[&:W?
ES_EeEYRBG\KC)0MbJd?W/SAW;cD]#ba+\HR][ZMZ@b+O_HH73XJdUT+\bB/3&eM
6\5]Qa8GdPe4R0J4O8?3F+:PMV<:edcDUfZ6T5X@d>&PcJ[]Hf8APR7</L#bY0GZ
BANW>c#Y[^,DX,g?W,IP+^dfVZ8AKZeN)N36[35+XfT#4W3.8,&b6&J?;G>e)cU4
3B-5BXMQ>9\O^6-4=GS1-=aXPTED&Ge41/4]\7^PH3RY1HbDa1>d&&74J8>YU+K7
GU^fEYB6WUMB7H-S^Pf35>55?ORYY+>M=\X;U74;:JV:A-/(#1X/LF3a5fESJeW&
3cgb.V@=5OGD>bKS02LIN0Z+SP;\.^_=,>_O;c2fG>c.R31V\Q],&DEebPgDDL.7
Wb[MS:[K;eI/@:g6K6/LUIV^LZ?Q/Y.KR3-a1;BB&#MQfUC&eM2eB/H^?.CO@+G]
PX(NOc;U&-0XCdW#XWA6/67F/VAKNLLc)Y4_6U?;/YcIZ]=4.J@1:WPb;<-/Y^X\
7IUFf.3GT<c38U_^dRQN9^)\_a-ZR,SY/@P-3bACZ1-&2<Bg/6)XB09=]KEg3H1X
^ON/ZMH1/7CQPS87ge^g6VA^^_6D1D41BH2C:Q)3SG-f9]Q#>(0Q9Hf(JVM;ROga
=f>B^UYFXZ]M(&6RG\9X\70N,&B@-HU-_]=.S-0&=SJMWb\<R25AJI^@P)JHP<A]
_8V47(B5Z+QJ(FfAaC;aJAEFNAXM]F=:>KV()?GSG^XA8VXfHgd_6ZS9[1W<fKeZ
HIM>@\Y.eHV[]VW14V)BE<8IRM083HdJC[<cgR/>=1c,,EFT_E2/7A&N?d4gZ9?E
D_.^<dHFYL/KPNM^#741Q^1<Zb96G[H^P])V3\Z/fZa0MF+BETZN;-DS??55RLXd
[\GQO5aOP[fK7LCf6</][VdQ8EZe-bDaJ>FEMPWDMb>Jf183ePWG4[#47XKDe3^6
SM>F,<09Z77W6W.+VeCeOQVWMTDT]=SA4]aBYMQ]CV+F9]E791d;Y:+41?=-V0d\
eX9#Ff-UB16AT.)KeIWdg@B=A&5JG8^Idfd88/Y.=0Z9_TTO#DN;4cBC5),X\WQL
9R)b3Iee,cD[9eYBd-e._a0DJ/(FOLE,1&JfY06:#.DVBGKH.)YNX8;9f7+Y1c#:
2P2FHFO_BYSN@(E0D8B].5Xc88=L/X.5gb<^SM:eP6F9V6a-R36_Q89+3G&5Y6GI
X#?E#-D7DeVQMPQE3@Og+H2EAEI@F?67EfA7M>ATWg[?B+Y9W-H5OU&5OSA3g>Q.
@348<X5D7KU:c+Bg(OTBKQV6O1\c#U#Q\H-)&KaR;Z0\gCg&G>4PO7eY:+ZaWM#S
1#D0A&6;TVZO#[5HPI_/9fe]09EPWKS3\H2gcR^:IBeHI<<\@^[T3]4g[d,gXZD^
XgC4XBS3_-@VSMaa.F]B&+GNgM>,5V_&LB>/?<:O^RLNBMCUD[-8a2_2(#9TI@6E
R=D1bH:9,Uf+^D6SU=bPD#=JT9M];XbSSTZaTCI^J?E0DKLY;<F>VX,,<8345VKP
AF?c4I/>L]GW/;Q1b@PPSHVGg(U<:?;:RV:GaKM,+c-#LLN\g=W3<Ef<=[R]2;-S
aN3^0M_W]\cgTYDGGSZZVeGU@cLPdU9:U0f#G?,OccM\.L3.?6EOK36IY.7WL;5K
?VV>L&,&ZUCHD>RdTdRK;2@+.)./XILB0A(Ob1VF<11O&K_YYQS.W>^WJ3G+.cG@
CD#(D,N4&([_G+V[8.E=2b#]Kd4d37>OURG+/=Z6NA9gBTS?E2#HN@HC(^Ge<U6G
WScHTa1Ma/aNRdU31KC[24B.1W:?H+gVeOD4+U7-,8>Y0=:.:e--A;55=]P75:15
]fDfD]00L<K3Q#M?T8(4\[AD-8^f(CUK[U?RCS]ZdN)CbP^9I7LT>f\A;O.0,E]1
#g<g)A?B&4IgWFM5(g8?>V/6?OF;H/,,O^;,TW#:JW+OFS?2]5K??M0dYJK/_.QL
fGP\9[0(>Gf;N#H>ZFB?4]bM[Zd-?TWI>C^^=26Za#GV19Z-Qb2Z6<D/L6e0Td,4
(5.LJ#.,dFgYSeK722c0:^b2_e.F]4Z:g[;((dEN)[]X?eAcU5>+NPc,LU3IK8)<
EK,FU;8WTdP1S=+1KLT\9I-d)9:QD[I)4]K#=?LM7dGCLL=bY.WSb#U\GAf/[90I
TUB3.2;)@;aGbdc)^:),(TG:JGbT&V<]Dg2WR5)UNSgZNeJ]KERF<A)U.(2@8,#-
#dQaKBE/bKC3J@R#>XOUH>fRIQI1@/BGcA&I_YL(fPP8[HY4;93Z_5?P]0221A1R
?.\<>DYL+g3T_([_7<EU;;\S;G-eT=]LM>?X-gM1NIVfA\ca8?e11a>?.O3FK0bL
<7EE15f/eeSV;Jc+ec[&0KPYaJ#3TL6MCA-[+AI2C&Z7PW6T7B>&H&G&F?7LSH//
UJ]XFF<1;a;]+cY<^#^;W;HW76Rb]Hf5I,eHQRV[@&#RV<d:7a8DI12],Cb.4bV9
dWc_>FM=V(g(2[,UMbd9X\VaK.^AD:72,e3+Y.5fPV-CKXGCR6X@0-(T4de\-QW[
VETGg9aDad-ZTTF7P.eL)7e]MI=D?JOegJC?VgXd<+Yd7F33(+MXP=42+\g&c1II
9DL_<DMTJe\Y@_RP?=.FOd;O2FY5AQU8EIBL,ABB^4fbIR(WLQ]_X6TBEeC2C=(?
U8L9aCUMUKHI\1B<@1C\JYc5GgD>9ZJbO5[Q+7::3RQfRYY]@;b-?>\]ZFb6CI)/
Cf@ZEJ--@/H#MWATE;?@IRd2;;eeQb@c(Fc47dfS28X[>7)_KY5cZ=c?&3B&IWQR
)g4IK1fCNDS)7,CYCWU2_Eb[8e.4F;0_2^W3S:L.V=W+I;Q5J\KB8;GB+2MUF^42
DccRaJ.MF<_Dg>[N(\,+/0P2[^_Q=HABZa0dV[#7g-137_M.;O@gG4+=09UKHa&?
U:?1X_EIUF\IV8b@)MNX+Y&4W2@EWX&/e#L_0H,9?EXV@2B=d,e(X.L7XQG_>L;b
MCDQ&Se@KP_Z9&Ua]dGHANP:GRU.bb3;]\30=f4T/_HTS.HJQ5;RO;Ge4Z^&VK)1
EKZDDJT:K5&UJbR8P+(26KWN(TI-@(b@Ra04-<2efNAdS^^[@3bJ>._6Q;EJg)I\
-8T3@JDCfQgCR3@AeL/Vf&\_H@0RM=.G;W?7_3eGYa)4<6Rbe48Z\:RJ88;e(Y/=
.S1?:HL6..6@MK.PG[G/^OFcLG7SHRVe&8:]2>08Y\eXCPH^.S.7NUKFDV3dJeOM
FS4eeT5Tc8URJCMdVE(+77a3#FERAT,Of7\_:/b7W#ZeUC](Xc2C:7,[\cD2CcZY
-^?U>=f#eZc\-eNKT;LZNL\-]C9?U2eJ^^bUI@[b1J(O^)SV[&THcCd,027;X<K]
gQ^&0JCWb.;7CJ0Pf7AN=dU,UdB,\Ig9,]2F0?2^Q\5/2aJSUZTFa1]5^SdI/4f+
^C#V&B8H./QE)@0[OH0BT+7EYbF-EE5[7H(4#2&IZ328@O5&9:D9)>2\E9UQAR&U
RKJL(<7Y6>6Z&g+&@W2X@,/];d6KJ#^>T-Pf[>NXc@7W&:_\0<R@G4K\Ld/H:PK^
)(BJOW@E2-6KWRX^Gb-G::@I3Pc@b]JJI#9N5^CN>5DUW[>3M[]7E3]]8JZ1c;(/
IZg_SZWf>.?U2Z@3:X9b8]+R.?KUcU.(f?>W^RDF1Y;6&;FbaC>L;8f&g9#Ha+M+
]YBC9UbXYN;_T@addSQac<gF&XJ/]/8S^A=bB;>5O/,QA(IVC2OV^)X&V&1E1ZH8
CR]=[UWU4+T;GRC4_]=1Sd#-]X98I)f@?B>QQaWB3DFX39.B?,eDZO#U7/Rc9d,U
@^W,W#-PTOTX=S;),^+[4#\I:E/PCS5XXc+D33W/+]GV8_PFRM;A<G(;_(0_a^T;
J;YaM=7IEBW:)]YEd1+&_8XJGd=R<F;B#],[6_Ff&?d,O)0Y;.D[^EP]ERR@3X&4
F^KP<FXa]:5#LIg:RY&+5>e/6d]/)1Og.6Z;aOQ90[/f,EY7X2-8#R8A#RG\M^V<
B-)bKEeCTJ0JD67,WIRSdK1BS3\]e4]2?EH-N4[^4Tb[IcIPCeWD\#&eQad#G,2L
VPe^4^#1g9[]<@][eD56/8,L,WB4+&f-)gC4d1F<K9X^b<LObIf/_?A)#;R=2#TV
L-P&aCA:b4.;(1eI@OJWO\W:?H^M2>LMb)7L9/5SFC]W\9&)_gD/K4\g8O>&O4#Q
aHXO+S4&F\F3dcHIS2F.^<:&1+Ld@&X/P<E::f>HPOIf2NESV8c+YCID@C^16+EJ
9Cc#89a+gUWY#EA_e,&VW#>N-<<6JX^1DeU10J/[K@-HV72[48L9;>_GKFRAFF.R
HX3P0W;:[:<?,<?IM6KVH(I@:;;L;6e:#:M<I/_QNPYR:(A9e)KG^LTU-AI?)eDa
FX\LW^G,@5UV)]X#\GSfcW.^g-8G[:F?URZ?F<>?F.[#\Z+V58Xba&S=,-(cS5bP
@g#W)Vf?T0P?V24AZSZY=Nc#O<VWC/&e?d\J,_Ta/HU<Rg[>bL=?Y=OXRW9TW\;)
A_(-gMLSdc5&Z;.L4LITDb\-;[CH6)YKQ/#d@I^:\SWO[23;0?c,W#+FP\<1b6ZG
T5&9TO)B&X/EQJBE(&R[6?\+FKUbReXZfN(;3#\@5g[FJ_I^CgM0]V<U,?GaUZ3^
.J&,H_=8a)F)d/1Qb(6QFN7R25LPUZA5ZJ]B=fJELXFfd7g[RU@_LXRV+MV;d?RQ
@>Y9fQU]/W.@Y?(K[HV/f;9.N7+:Z[dZ#0S,AZaCD>+Q>Z66N-La505:ZJ7bR\C6
c4C2)2FYB16&I[DH9a=#/LTff(<fTX11WPE9+V#9)^PZT],D435P.BN<G&:?^;Uc
R#9)SW3B2g:=,Y2a[&b@fP]NA1g.b<J9cT>F38P1AdRH)&3+YIV63-?Z:-0K>RD]
UOJgI:a.7<^6<Zb_5<9,/]C#@S0LEWT:SMU>9-Q].SBg.bI_Cg&g>?;B.-gLF3b^
AeKH-);[e^7M5I2UZ2XGYK+7H@7a/N(f>Ia58(@SU.b3EYR&Z:M6OR:(@AJMK>CA
D#R/_35A,+K(efG&gV&(VAb2BSU?^a1RDD^A<FFMBU^WLU@:gQD]HMF:[27D0XN7
<0HKf0CX7\5DYb]3K2ES4Lbe8AA(9=eK6:_L<cSIOE/;C;f<92a-Gf2FFQ,^Q:Pf
8#[R(&SWJU,b[7YQ3B^Z#QAa0R^VXX:RQB_NQV<X]B/M=N@Sd^5I\=(d>Wc[f_(9
gYRXO2AAb_W3[e;cW][9]JdJF0VG#Z.?.=+bPYTE\NT>Pg^g]M9,PgIV,HUBH19>
A.L>DZD-?Y\,&/4:dFUZ20:OWG&>f8\M2O,..g1dU,VYGK-B&XN@B0J\N#9dCPDX
E#WI99D\aT+H=/>B?+2K968^_M7)?OJ10O[JUPbU?,W[G>)M>6Re2U^=HL)NI5]f
J^HPZc1H?I@E\OPM<?>bQN&;3a1BYMAc0DILRX(HVP1OLNOLScN[G6)ZX#D3JfDa
#[6d0=QLM(PRDVS5#9KPU8)Bb<-dLHY46Zg>]a3HSD/(G],/bMW5;PN:E-H^.I=0
6f4G8e<OI;I+&.W]EYJMGNc4I[.c:[=05Z&f+-b4<\>O<(Xd5/V5J/7VgJAbF[VU
_d78NZeC/N--\IX:G0=#B^M\Fd/eI7<P2Y_)QTOLTX6_.S//&\eF\gU91,VWD.9.
RUB7aPM++O]c]/2-.HEHSW+L8AUM#5SeIIRGYI.F430Y2TW3TC]7X:B[bHXD^5e\
>8T+_9<S[S@TC^]7:]EIV2<,0TXLM.Z(B<+-RK^?)N-2/H-DI:/YF,M>>5;(7AeI
PbRG_4&/IM9VP+54gbQ)=RI@I^II7_5)bb2)e^e,G(7eP:2>8e58]2IA@,/gB.T.
<)1<61H[?.&<C-J/W)DaEYZR\J@8K=M,\#+(9,M1c^a,R3<,<Ydcd0/eURWWXg6c
7Xe_5/QAeX,Y7,-HEG)>?G<+G<.64OT9/20C7AR>_Q@\#NJ=/\7@I00SJ]-)d[Pb
)\9W&VZZJH0_/H6G6fW6PW[BB&[c,2YMd?J#^ZOZY0,V@QeMeTFcA;M;gP6QEV3U
SN;364#VVcHaNWgTaNPHAef._S0Z+PR&RGL000e/^aN=QBL(0g7AVRFS&@\dS#7J
R99]0RK/,^;8#gbSb9HYEA;H>b@FU)g2^&T2Z+TddQd,AIBfPJGZgc:D:AP3g^&&
/WBbYZO>7BeV[^2)bY0:VH+=9.&1gR8g(dC5-H==S?-NIYU;NR0J(5WbdMGP2WNE
-RS/I]SZ&a<@g-SJJ>D@OP>YOO^PI^[&MY\bGI1C61#dUdVDL>+@3WaQMO5N3(9G
O^_,I,1W?#UF/I-_bHAFQT?Rc?20+-./e@.8/b(g_-@IQM;48f4)&ZO<2#4M:aMf
JTe._HIE;+TDAb)&,C9PeDC(^D>fW<C740[\7&&7Af9W\cGD0\^=?T^_,E6XY(cO
2BUVERg>b,a,?+^ZLaQ4#];HG^L5.R2g4cb3@K2fRT&A0W5c3..L#fDD7?/BLdc)
^A=?X3TNQ^daV\AUKQKVR+ae@7S-R+]3cTNgVO7^S#[Ye/H_ZBAD\1UaFEN]Qc12
>&\c@QIA=dWO<L6E=4CZ9ZIRHZ7A7U3?L\8^_We=U;=VYSga5^>B^1g=-Xb9(cg6
23^NJIaY3Z\@[U\#@,)#IEDR4Vcb\-NMb8R4CHD/d\6)?WgI:E5g3Y)@,1<9XcL;
0G(E?KL>N.NMDLe=a^C7HLRI62cRTfa^G,M73gMM<Gb-F;DPSHT2?e_->8S(4X?b
O+#TN;Bb_a92=40<A):CSHFR63R;8L@S@,?#75((0^d1)XJ_9RRcSP[_MBC5cE);
59P<?^g7B2>:ACSCJGf/IAg5b@?CDRQV>4SV(N-+N:g(0<[7Y<d@ZgS@+0_0)G3Z
+<<GT]QO4]]bK+?d>F7eDDaPCFR+Cbb>0+G;Od[aK(5]WHZX/0TSEU<cV6J9LBV^
&LOWN9bYHe>U2Cbb2)gDG8GgXc/:ZAKHcZc:\DY3Y?aR[1NX0J5X+02e7g6.fMA[
9gWZA477]RYKKYD@VS90=?NQc/WeU&,_Y]6cC\RBg.GODN9\E[?^0=IgYd71/&Tg
(IEWS:6>;R+P#(KLH26O5<f5?c,eB;B:gQB&Ka79N?Z)aLW=FO<ZL^J;BS2\PU>#
<5XASU);dO@52J)2ca]-2]7H:@WbY1b=TOK?HC-O#[8b]P\.W^WAEDONB0d<<4//
+S:D+AZ59TG5#_gO:K6VL8+(JL.[YQI1<^22N,3VWdU<:A7X>D;bAf4,CaU&1105
4Ge-1_5aeG-LPD&552>=-])\RX70#9/4+gOMM;KfBS?^ITcOZZ6aG]]IEVU:]61H
-B&.]19;&8SOE:3&0Z:,KXcZSdg2KBN3Y>W0_5S.aY9#.#,ZB/AUEfZ\&Xf@U\RS
.P?=Oc6_S8#>dT=[\C>f[S,1d#H9<09;,eg[5\4.[fN,fALSUQSSH_S>fDM=<Q<Q
65SSNgg(6#:6L2aC;A@I\\0[Hg648AU-VER/?/f.C4QF&g9\N#P^<MX8V47L]gK\
8g[,,3E=&,A=RVP5beJg/&G)=GZ;QH,UcWZ_LNM24[cEX7\9B\7<A8^aXH9BOT9@
?B#XU1.WG]ODJC5H-XR)<I914K)(WEBAJ3E(Y.#=P]Y:[]ZWc7JL](>3Z[WQBWB@
-N87GIJ?.I[U,GPGFS1+RMZ8[+bg_7=8:Z+U]We#8MGD9AC\#.]-K0-1.][GXCc/
.LK:)0f[_[4ILFdFe5GF-=:JX(Cc.++9:[T(1(ECX>T?=ZK22^N<d)6U\;,^DcP7
=\KReQ6)SUBde-6F;SV53_)6;/W4>Q0VZERLD_RJM^c<H(H5cdGXc^JZXG6;@>]2
fXXGFV=_#]R9:KePa]_gK)EKdFHeG;(>D1,Z(f;YKEa^@H7f05Ree6[3VJGW8Z(Y
PGLf6Z7[8R<a+?H>(4@^6#QD#eXX2(2PXEe/V=:I2>9;#\0,HB5_6[2e0c(S?:62
8I\3+G=JZ6)Z4.+55M2G.]3B&069TGW,EE0.1]FSZ1DYWKN_7#6>IcA+:QKIHQ]^
a18Q).B5Lb4@X/<+.a,+=>.2/bJId#N;EPZ,0-J/O?Yea41#5K+:fR&9c\NZ+O#T
[F/@fbPe\3EWNHO@3X,?/(0fT#BARM;B>\]ZPEd94=1-=D4RTCFJ@cE8F<,\HE#A
e75N;ZH+EbFQVJg\7:#@:bYOQ<ZQB4-EB9[V@R1Q^=WW?=5CPO=0NQ9[E(^Z:H5E
OKL1e3J(>B62V/,cT1OI-(>a&4eW<P[,,24NT\/I8G0CI3A]R42S48MBbY)cb+d.
QcU<:D7-&ZUL.S1bG3-3R()PJKS.5L1BGAa/G48AV8/R]HY^)?Uc5RFOD]5df&L\
:M1UeEPA=cc,>S3B2Fa+c/gO_Eb\9C#_0WNgE/f9:b_c5\Y6_;@C(g8ABKK[c=-I
D?P30/,(MHG^eI0WB[LP2JRQ(F&?Z3=PAOFJQ+9&9#.)ZB)57G&ALMI\K++gV>Pa
W-(LNWP\7,bSNK\5-F1T_R0B9QSN/6K)FKH0L72FDZ>6I61I2]ZU)_FU\2)O80W#
20XG^(/?E7BBY:gS:.[E[UR36JZbUQL,a;DJa9YCI3L-PDYCN]c]OK(NR#65HNdK
7_SY.#fKC>c#ZHLPg>SW+11_DZMGLC9NgO\)b,LEe/F7)JR;/]YICcDA+ISWN,I?
[2Wf^+R;#AY;1b.8]@DGPX/.<U_(S2[0,dYIU>Z78?E@@A9-WJ,4.A#Q]H\5NMa/
I+61(a]dX5[]TgK:M,UHZT/=0?S25923bd:-f(HW];]MXRg;D>b=]=(E<<#N]GR;
P;Te654&?R_->dbQM,_aESV&BeI0Q3MZD::?=+WH73&T9AA:P<3C?JK8K[+PNXFa
Z]=J1d?SYXZ;/U()T&7[,M/f]:D^:OB@[fE75g^a(?3V+QMVZ?^aCQNXAYRH9.NH
a&Y.BRa&X([WFaH@>S]&4-_.U<OTI=QG\1FT2\DS4//E-fD/Q1eJK3)fR?0B-4^I
@Hf5L(J1FaC3W0K;I55e^Fc6LL70N6T;XBc)ZgOO/+19RA8G4H:X1887+M6G8S9@
2:&BIUGVcC9W<7NGPUDf,fM6_5U<8SX\T6[63V-\A#^=&CDHQfB/d-NX@E_<DG>\
MU]4]2Tg\?PD[+&>e6@D,#dCLa+0)4IReHF+\1LXCK8]8ed;\K+7,L3QfDg?FUWQ
\He7)cJOCcc@#JQ@:8+V?N9Q@ZQEHfR;1Q;3c.J\V&@I,TbH7?#A4>:BLZa21_F_
Gfb\&c4&)9Ja#@]>bX8Ng:1T[dF]b;:IPXeOEW?bV^ZA#Zf=Aec4Jd-6IHXf?U;Z
?\\.Fa1JXLg#SAB-B(]PICTD;77\B)FZXD<=V(DQ2=XNU/UeR_LU(gW3<fN^O)/T
e&DO6D=.HPS<=d._&FC@GL;NS8\QTSFNR-.S(fV<C+:SO)2P9?DK(X&7&(D;A:74
CB>#5cB85JZe:<KH/Z5@GNX;)3ZJ8XYV_\-d3L#AC#0V=[EB23dZV&4;#A;2UF^:
N,Pf4;H(D=bgPQOM1,5XcI>,HH-D+Ra@C=L-N=f+6L]B@gY=-3WdVWc=-/15=e0)
CNQ;2Y)\S[Q)GPd6/VNO[([Y^+06?Q(2a5]QOGW[c8&PfH=?:T<,Z4K;N\>EP=:;
G,-:;RMfL^57H6aEW?KfM+-QS=ORV&]cg6^Q<)KgU?2_5#Qg7FbX_0cD#;#MaI;g
Z++8dH:-R(.e&EA.#.5>d\F@5NSI2>(fW1?>2^882NHe]S312.(\>^Q5F2@^^<EE
HXM#X_P;IS(;^M;4:5D4O6Y9F5XZ+906-@b])(#(4L<35Z3<6P3]DZ<C+^1EBJCF
IFG7JdbbDc&5<7\eeH<P\I<SG>DO^0[MQQcXQ7OEXS-#\>.C+fBVY1/N_<##X8Y(
G-G0Z-2X@dV:WEe:L,QLUC?85QPEUQc[N?U/?_cQ>].DJHVVQa5=a\WGX<Y&>R-C
Z7IJFNgg+.a<OV]2,A<R\JaGgeI9BVRbMe)QC)dGAMJU8,a_\^+(RVJ3f(g:,AGM
\RbYL@7Rg3/EB]64cH7@RX3BDg[I(J<RKA_W0^ZU#I-#d8?;g>6U>QT&)bY)QX+&
,F^(>23&.XTD2A01300_L0QQe;S.-aVF6P@0<R=BJB,>5e5^bB.-UNH^(-\dHgD;
:^S=,TD.[&[4WR1dSg^AfU-c=D<+OD5PEUR<CY<dOcNU(\O_OUMKF1+Ab3T4gA4C
#HG;(AgBIS?O@Q8a?Q8.CRM&H6@2C#c?N>&f]4dV,Jf>R]96@2IcMKZ2RZ=;Ja]P
R;GS]e2UIY_gU6\8cRM#T)f#X6IW\:c:?2(M4L)?e&eI2XN=E>(eGKcCZEJWRKIB
Vb8^9:.?AN[A]7D+0I@80<]+2Od^XDSIF2Y5NI/]@?U<U.GH8YL9bMU=?<O16fD=
aWWDM+fAG<V:@/7FZVKL19);X+=0115WXR26W8gSH#,IIdTe8V-T?O7R+P?6?3;\
3E9,[a8R:[=NE6c.GQ9J=#Qgd>-\(e5)@/e_cXGT4KG04ZZ0AYSbZ1G8AM5(_aP4
Pe1B;[FQ53HR>X>bXGaMFBaI8=:N+;N&QD:N@@\1DN9H=SL(;_IONY(Q7<2P)GO_
_B^8F>=;10VSMXKUHB^P<EEc#_^LDJN0W5F-OTDL_?B9@[d;A-(0V[fCY(cgggJM
SAU@I4b>C;0@2F(QWMb+^ZBCf77?)1NE&=WZV0Y2:NJP)C[D?N@7\BJ/\@a@<#-(
Z@3949MF<_F@;&3T#b=(V;S9ed5S&/c6H,EXAJ=ZHYW;/OZ&a<<#\((9I\-/BAg6
+4/8<;TgZZ7b@9/d<W[+)Wg8AE<ME^^GUQF]cWA\1FQ-CT3MK)R=9\B6;EFd,J0I
<M00g;YRAc4+9JYV8aCc&dA@)Hd&e?e.S-QZ]gVFe2W,G2>A>/XRF>-@<)gNeZTL
#:3<R-JS\=II&b=3NK,T?P4Lf7Q>L,V7>[@QBOWD67NeJTKVTa0X0dVT+JJI)06/
C>dfCa(=fJ^3X:U1NRY(@OU#_\[W<5MfQ(6<fU:?BR/Z-Y_9QA1A\=BMT?d1+Q2O
:EFHgeI37\O&3FUC#&1?4?^Ee)72be(8VGN1G8fUR9N5X^_[0JTAd7DA;SfZ+=-E
KWSB&TA3CHT7W:gQ9E),D51b/&:6WC5^Sb(T6>=Bf.+M1IPb(EYIaNT\R6g^@/)6
B;>7&=QPG^XB?0LILg@]X6O@(DI9ZUf075^8JeDVR@bK1CW1;J]],I>:GZQ/dgI[
H0OUR&LE38a_?eQ\S-If9dXV[MXZa-+WFF-X?.[,SV:ZEP)b<L6[ZGg9J^_AUOCg
cT#DYH:E>J-9+c>?=1,f#@O:.ONXY\H5JO:33+C)B<gT[UQ3X8@736T-+\O;bfY2
#1fG;1MP7#7FS(L=3\A[^?3HJ)QE6+f\^<3<V#gc:5e;2#cAOR=M@+N:^,I/L0)]
L54)fYUYS:8@Q@aN-SeHC<O3IO^]85.NS.7gQUEUb>IH212Ka<8FTZ@[Q)SUSe_c
bTK_7<,<RV[R),82?UYWI_YgK=6AC_ge])^b^BdKV2fNdBBaA;0RT+2&4DAd1eB>
_3a+(@Y/Af>[\,@d;7#UJbPTbH7G,8[d5FSEC4;>4?RJgM\@c<;/O.2<(@Q@3?b:
X>^;&8TVY]AGGZK1E4+U78G:X190,/cV[=X8d2[ZBT&KQEDE/LLR2B>6)GLI-(Q0
NGdAB9cWbfI@+3HVZ+0Bd>&:9[9WPP]#E#XF<aC2_8EaO?@[BC#=:gDWRNbb@HRL
[.:O#A2W/7+4V6#R/dgDD0Gg7>=Y#E=8CUN(>I#X,NN80Fg07,LE-YHe>2aA;MN]
F7&R5<@Oe0GO?_S>Q@8=[;,9,6FVU#(Z#E\Vb82[WHG\;<ECCE)GBBfaD&+4J5^^
eM<8M4N9TAPQ,+A^//A<YeL^3>9?(,M3BA4[J]HaM4edA(g5d3HX;S#YO6f4)B;V
)WC8P[9)TJV#Df&(6#?R+=1Q)NJL)\gAWPBML&P?^2W?O=UQ0.@KTA&T;NU@1A8&
5=A.9S-eCfXCU2BdAW5<2EMD4>bJ1?E4]YB08F(SW]A2f/K#T]_:BL?d=L8c9?-3
5,)O^K&:#6b-Neg0Gb5:Zg=TB-G_LeRaJ0(4_)&9&++OeV)]NY#^DI9Q?39QH-F3
^;/;:VfQ\]#M/09aeDS3@54ONSA_RIe4G/1I\+eET4Wf9UR>HRUYbe]^W[^_EMd6
1N_U#U9Y^.H2/N]Hd8INJ;+\W]J0<R+7FS.c4-[7b]5@NI@-X6PC4D6P>#2?F)ZT
,@ZX2UXDV]8F(,?.TUF[_J_^]#4K,L@V.f#K,S#64\]M]7<&0V2Yf>UM@/O0b6G[
P)c:(B:NdQZYPf,]/6:_R-VN#NZ48OTc^D^)2&I>=f00N[Xd3ZKfb3,Ue5KM;[54
g9E#La-X-cI:W_g?H6;(e_1D\FT[GDJ)))TSgO)<B>&,P.\?#TA:G&;9A,ZBJN[M
=La6(0EE+.Me25[(TF9,U7eTPgY6&e&J<>9[b<6[FC8<^3MZE9WWO2:+4O(a##BF
?GHSR9QL,HZVX^PfSAc@+&;:?ZHBDaEUTd]6.4J:,G+LA01+#HeELVJ5C98bYB#Y
4J35:.LQ(a&[59.M#S3d_/Ofe/GTVb_)BL2eH+QAg3a30TUf5]A_W>1aR-H+PeB]
S+0EI?6fXfK4&2WeAg\LIXb0:>H_70&QGZ^@c5JDSc3PB@=/=V>c:0eebAVA.]2K
S.eC#M&)U_b:NQDd(_[J5YbSOV?LV5b)f_9Z:dS35GG\=AVe0&U9\OG/e(\55+E>
65AOI&(Fd9#a7WR7=#1fJ54#Y]<1ANTd&@X/IJUgc-7(9+@eXFWP]^R2IMXe3[=X
)<5;-CL;HZ(ZG+1LRfN#5/)^>DDb@_8IDS1GZ#&.3/6<[1L#7(Ce\]ScdDJS4aE>
G:FBFg\abQRagF;;1e]WJ@12.=AH7Y8:SUeKU=D.(E4;\G9CeZ[K.dID3B(DDHN9
gIcEO?PQSNA.OO,#JKV(B&J<(KDgW=HA:=16@-+>ZgMVgV7.9C<7MU(TGX:;-2MF
@\293,?_P=CD>>,\-=AS^Ed/Y;f;N8TDOc-H\N/)gUQYIH2?=X/P++15)Z?I<T(g
&7B8[FI@[N9F20EX\.2[.3b4LVBb]D5D]=W[+&AdQKL?@OHTc3,8&\F._#NS/DO^
8&MB0TFX7bE&cN.g6\.\TW.]W>R8A99GFG3^<3Z15c&=dL(Z\AN,(092d0U]<E#V
\=^f4OfPC9M8S)^ZH6/@S):Y/+@g7OP.83/dN:7I?+:/NLad5RWV2I:U.4PKg(#D
#<DTRW1Ie6[ZGHQ,RUML,.f1SPTV=fEcdU8Q.?=O1YAb0/G6)7FF@WPI6MEB_OX+
)T\@:,ON/-0NY\f.0>]\;Ga8E+JN70?+#^>fM@B0Z<(;=\<#4f/S\HYDaW<0._3N
aAJP;3@Y[d3?f;f=.?ZZ<;N6PH#7(H\ZfYM8L2a@8?RPA0BFE&UfD)JFOK5(4ZB_
JbV-U3OMIA7b5R8(E4QD0S2Sa;0cKLEIg5H&.DWBR2]:(Pd:O1Z2a;0ed\0K+<g(
-EO96M[LY=_85(K#UM4W+Z,G^Ta,I<Sd,7Y:&+I@@K<BKgNL<YA,GQT=@ZK73])f
Z7IV]=)(?dHF>_a#.ZN]SC6B=[JDUG4eL+809HT/0M77P:C,N-ASd5I[VM2PJ^A<
0.._K-,T,_0GU8C3A]=26N0b6B]A\gYfHDFfY3_5AFM,B;]4XS<PSKXM]60]K?;_
V6YK9M\gf8APV>]32DYA<+ZG0RPe4UEPQB^,BSI)I><4_TYId](EGKOJW;+2IWb;
=1>O_FJ8>YPF+A9EK2=Lf^gQ@e:?L31,F=;09gd(gN(,GZb<Ud//.C49)L0736e7
4MV]>0?QXGcD2PGK?_457/0SZS\3L&Be/.Z-DMF^+MZ@[YXTW->OceV#;]\Q>N[S
2-?=V23BRTQ:C?2WY,PS\ed4dMeTTR]KLYY&-afWC=##?fZGK=Td<_,_V/eI@1J-
\+7RbX/4^bGEf5bEO,?L[7PgEb/BM_BZP6&bL4cE3EE0D)1=V&H9>EXe@?f=<__R
5]2<P69[6/A^((7E?9N8f&LV3X\4UbUNG9_R3ACSHFR61bKHFZg4>Lde-7MPAD0-
0E0-a]?1AM\+]<T]Cd/BV#ce[cV<N>I8>\\aE8\G,D7Q[[0c8CI^[bSY=^SQfP;G
>9cR6=-I]Fg8-G?:+eZMU\0Z.g?2_d3H=69bfa&M->HO-c]d<PB7H=(9W[J,gVcH
QN,SHTaCU1e?T5OW;f7gb\05>Zd9d\5JSXTV9/b]I#T0XKL(a,NC5ZAGH@CP=X<D
dAGU,QdHW7D4_A+:9@I5eZ0S0(U^CX?Xg,._3M[2XL91ec0SU53,&=bc)&0VA9gD
DLMU[L:<X,OP7P/ET92&]N_\d&)Z<CQX08,C6?TB/LI=>6[dV(GPf=6+;Va92))2
D7COaN-5&bg]XITgG.WNAUTN@K:Y7WJRGXHYY@DN7G0\C>4C.:KI->aS4egY8/P,
Y;45<=d>93047I<JVHB(dR(RT?[-BO)+-XbWD)O7cRFM<+AM[^Ea]5_T&HZbRFeX
NccHDJD@efPAYVgbBQ]3=f#/,2d(=X78@(<+H)03L0cEQFQU8CR=2fXg\TN,@58g
OTIV[2LCYJaNRRAfY3U&?;U4C(ZM1e-Kg,#99,YXS+QR=IQT;GYN;A>,9>S[:M^D
/_;527gIPV21P3Tf1P2YSJIPP7PU&F0;24?3/W_;bZD[(HTH]=DQG]P=6d14,#Lc
PMeWeC3P\8]P5,/2C(If__XFg&]]\GROeIGTBOMH1aV,ON@\d]0S:=6,:5A;_IJW
J/Od/W03_Y#1=M/1DTgUFM)M-]B9]gR/Q=AYc<cf0-g7(?gHPT68gGWBJZIOLGc+
H#Y+SaD-J_/e5OJaLa>(>&TCL1PMg+S[dUUL>G/]KS-])+GQ)N2.>9:0\BG>S<F/
9L+aC04S\?+4\DF&[fEcD1N2CTY_8P62KG.[M^fZf3Y#DY;e,1[;SE>X&5Y3Gb]K
<:AK\1_WfS]CfYUgT[1[U&c/E,B/923_0S?KSe\T<LE<=\g7X]H/&/VRfR@XZaA9
_fdFM&a;>Z&AdKc_E/W\_cYA^&]NTg,EAgP?K2HTRIeGT_H=P75eeIbZ0=&X=a4M
fJ&=?TNL;P&QfP?g48B:(V23)ZeOb.KAA,dHUJe+e>Z,R;\_cO^C,e+aR<,Affeg
5bcU829V)0V^+aKC@aGP0-3fZ0&cTO6A2N)gW5ad0[EIC6?^dIE_BTOSg,dHTG_Y
f1JG&Y2)f?LP(OL#2T\6W]3V(\Fg,7W.g^,F_3C6M4L]O4R@2]S5R+?5f?]=DZd[
,cd]O_A@:IE-IMQG7cB,g&72PUc-863F#&.gBG\cZOAJ&BdGT^7VNL]([_1QYXZc
I>X(V3[5<7OY7;L/WVe)N8S_b.<VDe9d_YE-geBE\,&]9Zd+&VE\[GgfHVKK+Z07
A,a3:H>()=:F-.<7Y)=EdDLO0ONccH39PQJANTUI1<(B<C<g3(:Dec93c/LUF@ZC
>YTf5gIV-/U/U<?0@Z7GQF2ZL9g3,a>NbE<6b-LcI1:.fJAV_E[f\-Z=O0FX?Uc-
6CC0:ce\?IU^/6W,\2gHbK.GHeAOaPNX)@GA(RSLX#O1bBD.TRF1]Pb@(6QFD.;(
V=ID\(_aRHCA?gDMC+S.)AKY>g5RaD19TNMYM8gY)bR5C7(4U5#3UeB.)cL4B;b(
b[U-We;]<5.,_Y3D<BU1K7S_I0@:1K4D5ZXZ0D3F\E8EI7D+]Wc8>:/S+HdTMCOP
(8FNO]IID553^bc@cX^g\[a:f]T^NJNI+6,_1\Jg_]H/#?cIC0^I#[K89;g&SDAS
_P.#LK#2(,4G1T6TMa5B3<_3dBd(N)Z1BL/(915VHF#EXL[3WDF0^Y+RLRL>E49d
]?H+[GCWO9KQ&>SK;6AV&25P2?f59MA[NU6G(REQ_8ZEUSPKdd1_Q>>cR7@d)T3G
[Ec]dL3E0/?+<#/a+2J0)a6e#[=I.\E^</?,R#13M^5X6>;?[b<K.;/bAD;Sd,70
X=4-AZYS38F+Wd(,B0f]c9\6M6VPK2@KK7R4^OK2PNU#d0)6BWW3a7>Y-:;QK9).
=/X^.SA=ODIg9RF^Eg>OWg(eN.dgaB9Y=AP6db2UZaE/0W#=_M]-dOR1HEc^QGRO
6?P.?8RTdDQ_;;M16VgDRI?@?[)DMT)2a\MUV4_KE0&J7]Q>Q4V;/S^^546PXbH/
F+aDObAc>D\?EVNK8[e,D3I9f@/B7VaJ7F@GZ?&86XN1g34cO<QK78\UaGbG0=?@
,a]#XRB?=Sf6>cKe[@-R;_.::QSg<:T#-KNS]]eI060_SO)US;S]Rf2JY(-NF9+c
8Ng-57gU2a.gGW4^Y,e&Y_,M+gCTL\:(5RJGS.NTNZ5O[UXF\)?//W-afd+Q7\f0
E.bT2?NX=0WI@HDA]X>MSR,E1,D/>)Z&711GcN3H0?;4b2^AHE=:?]0>@BG6d3Q)
Ae.9TZ&J]5,F-?:YFdG\f.ZabLY.W;L_?UIW2,R@c?gX=3:g5\YNafd,TR.C;]+6
e(b;A.aB,O:KJ>L<Ja#RIbRL^)^KL#dIV/)YNXA8e:e,XDMME-OB&(;NOF?Q.E_>
OaaAYVTD+bK:JU7\@N>^_Z[OXR1d6+:2Q\;D=6Jg)/V9J([=?Rg4]b5&f^^0PC=3
S#1=H\S.3URDT,>B&eBK9c_UZKE;I^)@cS@V56W:KJgBS]0WX+eY6USO+6K<^?Q_
<>Cc^JF/N.eb^^([S:Q4\V[EQGC<+T;AT]<Kc&ODH8&[JX9<#YFDTCM?RUU=@bJb
4@.922Y_-9b_R=?)Y7[fDOUaWa?e]T11Z33=CWg7SV)V;aN:NB^T+973M==2+]f)
L]40bU#+4J:df0d(aSP(>P8B@T3CVL8f,(@;/E5aXe<ff4OVG2)LLBfT\N)G>e:A
Z75OO5d^g?HbYb;0_;-MONT@\If^=c??QDb&TaZPOIDefP/0OHP&<O:;N+FVcXHQ
4PeQ^>X#f10T^g36bT^D:VGW]^Ja:=)G&R7/O]fXbRVL[,<g<?=MbC2HXI-a7ZYQ
4e#U#NT[4#7b#\T.&7.K@B>2;Ud<fTY&N#ZKDfO@8KK11^Q2[b:BC)V#7g.Q8@D&
PX6EaP[Kge@X=1>>,X&_CP:TJ^ae2V7Q(fegR)aG:EM^<[)eZ#^BZI\3R:@V]R_7
=Q^SN>6c]MA#M/bT:S-T#^8\LDF/:>1>M&=1IC2+O;P<U--YBGC)M,VfEPdY\:[F
<\6-O\6FQY8_fPg4:[@\OdVIE1XY6XKPF.]R0RV2A9_gfaV)WeDYLSe<J&76);8=
]RF64Gc],g,\c]RJ#Wf>bDVFdR<DFIKFQa8a2AUA&7gS\(ABSNB8JR5J\b?^LX/e
>cTe[aOGF=/F9^(J[,+KG3F5fIcNVW\a1VaGY6;^#(J]W-V@[R#cGR]Y60eCD7S7
1a<C5_YL\MCb>DJ3LQP^M0WMLe+M.5XFB26AR=4aW,.,g)HZb\4T:-U0.XedTa3>
a>[426U5?]>dd[aG[4B]&G^\4YTFZIMe\:ZL[9S#WU+9a&ZW0Nb/If+ODL^#?)U_
AC&IS(YS[\9VI0XLd6OP<ZCD7X>TXg@IRQ>>D7d1.SMba(#.AP6LZ+c:[=0CI0YW
[>O3M.bB0UT^1X:F;WHfDT,-)(H/fZ)#?UXe&PS#U;6<_W83:f?BAV3eHNSY(6AU
:TRcd&6UFM.^6Lc2+88,]gd80@f=4e[AH&HN(4TR1S\@NUI\SQPX_>?N_IAR\-]U
(UWPdeU1\?HU)XE\@WX6:(?abZ-L=27-V#(7)8BC]^)IPV7bM30Z0KKLX[K613/,
e+\1TQ&IC(5@B68UB]TSY(E9^TKSbFMIAXUfXadUND4I6^Ha6,DUR28Nf?DSc^NO
\)B=RPgXPGP05&?f(&_VCNcDK#90B=&?SVQ<@H=U1#UOOSI7K+U#5]>b7;Mb_NaO
+T[QE]N5Eg^M../c?VgI<8BZYbc]T7SBG=:ZYM,b^7TbEW1(NPfL8+84c)(A#_+Y
Ue47LPQ@7HSIH6P,2T^6?[W&V))5KP+@K<dO//>><-I9]T64Vd5[V/1Z#d2/\Y9)
bFMVc63I=X;6a&KE\FUP/9FSPIXTW5P4(UggL.JXT-U6[.#@6+BS-^/fGFbS1GCK
PE34MH#9DQ^:Cf#S5-1H(_d\d8NgBD@Z2Q16U?)S;]_6@XeeN=Qea6D3_N;88<85
3,-+5F4#^^C_E[0K3A/O96@dQ820Q/N2;LdLE\Y#GU[4U:&aEb[d,>JI\AMMUeQ1
.:TdebJ^W<D])J]OI&&cPD<4^f[f=f+95M)6A/PDHd4I2Sc^IEJ6Z_WS1N_XbM0@
;,^gD0YdeXZLNO[OYM@L^YWG[]=+AcRdDR06Y+=3S3BLBP-,\Z=.ae)<?Z:5^cHC
UM>a<O]/8fU.7LAg[YXTgDCTE<SUPC)TO>4JE(926PH(:fH?Na]\GA3D:g+X]>./
4aed:_fe#g^IbO0.T@QI:7MANAIL(1N.;DA)]d2(>M\^EbCg/PLgP6bLG>.7a#-&
TF=AY(e2M@2f>aLdgB]#Sb#Z\_<L-F#A5gVX_eH(CZECbO>[@U08F\YWNfDCgI\&
a)+I\9)DR:&SOAe2[XEg7HC=f4MXHZ=Mb<V2d<2HC).@Lf0>B#b@OMNf+dBU4&Oc
ZD19Pb2BBXZQ&YV=3NIH(JUVXN>LH+-1@(UG_UZWW#1V/2[4^]3XR&c5]4\E9R4)
<2S^#Qb)GS>>D<U<)70\-gB,f,Dd#JEe;-]=[;Vf>PI4d#KPB;P8>02K_>=8S1]#
9BT6:e.R]JVU22bWfTg;c&VJ6_2#Y,cU_&)W2SPQgJ>NUFRMNB=XX/C)-P:]Q>?g
3+?Ae4R2T4)^/&POa(3O>^C#NGEW:+F-a=4f7A:\acTI>8^\5?(C-eZgV@XU^M2c
G82Q^4_=/:>9b;ZYd12W\bZ#EWSS5=;X6U3A39V+J6)cB9D+a,VJ)K#[=-5J1I<W
C/OD7:OR\,AS,N5(9=gUA?B7TZMEB]HWOd?FHFQ-=V3F39KAWI\XeY+1Fgb.AM4>
C19Sb)7[ZB2)E9,8G+8YQH230M(;De^NEG=g0()]YC\[4)<S-#)-QEf>K8dH;@DS
BPK1Z46:,:L[8YJ.M&gH29XG.F:Rg#c6I#OEfaaTB&&@-PXbT5#(DgG6B=@\Y5V8
?TEE==U.Rfb/+^e61f->;M6>C3=?NQ@:NE7aQZX((.+JNGER1S#XFL4c)<+4Sc7E
cSFce9ECB0>&1HDUN7V=5HBeOM.)/.DXDX#f/f]]?Z<NO+g+LQ471Z3@e1?G>1+#
854V8<V6].[(:F4ZO.b9G50NNcY:TB_9,d>8QJ\F+\>f6K/3F4f1c1MG:JGT@L4[
X]:&XCY07NOD_(DZ[:T:>(>;45;:caP)M<Y[-^WEYWB?FH5RO#ebK=>QF.,(,TO)
O]&5@DR7S7[B:Ag4fbN#H&?gGUT.4IS.IYT5TB_g/>]SV>f?3H#J23(TZS\_2FK1
HZ^,1IPN(_C?6T0=5<HV&^^=13VGYg-YF^aTCT7c-@(d<J#9.DO_2H^#:Y95&=@[
-O>UABX,4FKR9)+^T^1K(V;/KNMD)(#,.DRe>.EGV>BdbJ<RXF;a>W<GeMD^?,\G
]130@be]dMeE8:g1e4g>0QLO>b:XFYWR4M<@/ZFUCcT)d\+Ba^ZJ1W4-B+Y&H&XD
DOO+0@L@WJ^@/AEQ#Q&LYGU,7#d818F8LYO9;5DFCNd+86#3=HcNfa2Y,Wd#:)gJ
CSg0e[3NE@SOQ0VC&20I?6[]b6>X\VAHBgc#S>T:Y@c2#-ET4-]=5GX:^<BM:NIC
aD&NLPd?ADb>VD\Y@2NJT@.?a=bG9K9PbFIIB(Z.>&HUf_+?=T3deFA#b2-+#aXa
9P2Bd@WUT;,L/#d+_Bc_,cc\<R99>VOCUDQOLV4eF9d?b40(GE&MW;I/1I?FW+8S
)24Q94(>\aMd\EV2,=PQYb:I18CZOgW1_a#+TfBgJ5b/V+B9gM)DEYMaVGSS^ZX;
)Uc+d0OO(PX>Mb/@0=BXB0V5JC_960I.eU7IdM5I]Y+dTJJN][]M)67,=[b(f2\T
dRaZ9NV\F.=F1P5<V?[-=@;+/0U@,^W#W=RV/1_L&WCF-dSL>^?Jf44;(-#(T^X_
^@aag090V..W[(9GaOA-Uf^4&-8ZS>6=U?BS;Q#<+gKFX\T,a+UQ.=VWc)-fGfW_
/^SGFQN;KY).BV/fb>EO)SV?)d3)2ET@c6Pc<b<e^e9@>[X;B-EKEeZR^:J3JT-Z
=C>KB,J:[Q8DVG+aDUKBQ,HTT\)ROJUI\S2E_AM5S21SN/J0[J;OFZgAN,JV5]EV
[/EOWNB:ICF(]dTGY+4-c=D]6b6LLVR[#9e.T\CK=PM@-<IXVV&WJ_AQ4G3V^7DO
@A^\3WN]f#3IL@]<.:EVGg&,-cNVG[#PP>^D8bcO@QO-Hc^b3HL)B7S-I@0fA8=g
D@Z5Wcf4U<ZA6c5)+?BFaV0OC&DOKC8gb8]_JOdc0A:\^?RD@=e7f]_=8Of:dR0^
Y+UGAMSd33Yb#Ad&YO2S(95EV6@DCUUK>X@dZN@2;T:8R.L5?VXe&FTTb8<Pd^(H
P#<#GaT.0,>V^.IDWSL+2]:R2L3f1W?+;)HLIfCVE#JFXMXc\6+(;SX+<fL-6bMY
6V/B,.X4B]Z:>Y>P>W]B@&.c<ZRPNSWC1<GQaK.Q<QO6U-2M&[50?HA8\3:[;M@)
1g>=-Q/DP\J@XQ&)ZID+O&XVL\Y=W6Q]@]NKYAdAS9C8bRFCYFL_NcM4M>W@U>>J
<eN>YG?X-,Uc66)-;8-(]UU[W&191#5-DWb4F#I50:TVReBd:6967X?b1HNUXJ-7
7-O.].Cg0\D8B^bW\f#U)NJ0RN,@g#b;,B^B5dT^,MZeORd@c_<HZ/EZXVF7;@6#
W1_H];_)^-fS?W>>#&bHM3MLQPL<M-?Q:]>W_L),B.5HWE\[9gAHU\F01NaK+cNK
5DFBVa&DU5:^>YE=)793)HJa]^WN2,OQ_=?-ffD.4,5ePM@[GOH9:>LMJ:E4F:)L
FGE[<D-b-<G5AI)M]\AaEPRXKW;W-RIQ;H3+V^9+B&K7QFdV:]Z#[<6(^5f2[E>C
ZCbC,Be6Ga6&\2:NJR29FAQ]+,8(K;\\T.J_,L-@&-O-&QX8BB<X/AcYIOG4V)N0
D0BDS=.4;b600V2NCQgPc]Q>@ca@UYNK@#E[dV(@TeJNL@R;ZC4FUGO9G/FHa_DA
?eX:g8#e[^(V[Hb[JOWZHeJ3FO@>O?c-SQ;Qg7>g;gAK_SQ&)V-d]e[.K1,fIU/A
1^?F2:&+UO[A:.X.HZGG&PfK>P<]_beG/edST.JB2^LV:A6f;H6;KC2HK:6b]Z+8
)F,J<DDg.AL>\Qf9\JUGDFc\85@SY_OR/)S4#aQeR.^ge/W,)NKN>[A;BYgRZ(?1
Z=3Wa/I+-G]?-<2B4-5,WY6/=.L;R9ACb\,8VO3I9_\V<(cf&?=8+F4YA+,:cHAa
,Nb_)6,OcF#G1G=VS+9d-]YCYV[g[<;RN5<gG8H_>?@O=9Ff,E14N(.2G=]K;#W<
fLaQcDJeMa()I?eTc2]IQ^Neb#fR4+?&fAYXS)BVfM=\YCIWeP[L)&TA8O,#&ALZ
#U.EX]ZW>S;Ee-CHG^2I.5>VHUHJ)MXG5=MGN@7Z;Q6S,J^dUK^Y.2W4PJJQ=YHc
^=,1HJY)U,RS9^LcO/<>0OL5]9PVGdE]LPA<[@P4?Q,T-^^O_Pb<d-Z;>>b;dgc2
EbSD;CAI808[IdUZe69=9O(J-1#;9/F\??0a@:e9Y4Bg9/+d&+KZO,8RH)dWH)f\
BO8\P+.,//^dO#6_RKLZ__7<19gX)(]aAgb)-Y_?O_X4/7:T:b#^:(d@FH8X#.5^
6a:+@PXW0G4b3D/99<=]H+b_/?XGAIPGME5>gJAe/0>;J#_8HJCP8#]KgD@I+g,(
IM]g.aeL8Kg<RQISA^Xd666Q@K319+O3/_7#R8d5LcN0)Rdf_4CLNdCT6&F;;Y_7
8.)dIO[/N62H&I+OER)Z>VWKTfM.TY<4?9@bf9L-UG:9#8Z[CNZba\W8.&QPC\KI
-XKME]&Ra_7<&<1.6I7VPOA,SPLJO,O1@+CY0V>AQf=Z15]2)7\>M\.GG]PJ+)/)
2V-MWQZ#ab#c/dDR;dNT1)<0K9fT^YUN+Q@aR,f>Tdf@&=NP\MHBYR1K-:b[(;3d
A7XgT-VIWd\[7T6SI\29Z?.K9V#,^W[C2D1TUKB@L^N)ENQTM#B]9e,_6W;HG7-E
51TR8NCDK;;8ZT\]P^)>[_/^Q-=(&A.2WbBI^T5OWX@B681f/ag6(Rca_U+cgE,]
#V^g3+<Z(,-\45#9:5a(Qe<-]2)+9Bg.S6@BK3CSS?6/+SD&P6S.0JI>D_1g@TKS
,?Red@9^Z389g(BOVIZ+1NaNRE\;]bSS(&aV<8Bf+]N:AY8T]>gG;HEfC/U.+YgG
4]G6ceAfMXOZ=EaZ/;A^JabTZB=/^(KV7Vd3:CC-0Na[bZ>9Xc,7)<Af\V-K38Yd
9T,?BE<VSYEUK-VTW-KFY2I1LIIdIQKT\>G,V0a37G?;D:^@Q8(/5eH8J=ZVEFN)
c84?W[O,RK@0Z5V7Ed,AXF[N_1W2c;I5MZb+D:^H6/UX17X4M/c)Wa4J1[fSLF#4
:QY55I#[&GZ.9]&]b8L0YTZS8R#7Q3FXRcT?+J@][)G(U9SN8LP?\^.;KH0UGdXV
YD<B_[EfYS0I]\/94U)7dcVeWgN27\3(<S@O94,XeV=K_4,WJX/+)&D,#VF[6+/#
?)NVc&=?/7^6_S/a>Sb=#3[[cb/?MC/Aa2NIS]_K<F.7ERJgQ3H/0QMM3LD2A37e
W&^-Y@\?9&6ZHD/3g8Y5VJe50Ec/=O]5dF;Q1,?46?INRHdG,6VM5+AW0R_[=IMN
(LC5E--N19RF^ZN48O@=,FEDDHN(;-3[@O^36F?c_Z[e;^N^.X2Q)U[Q[cSR#?6(
C1;1bH=cN_HW3A(54R=IWeS&6C2F+bR79LD^-#6[NY_cCQ9fIAN)J:=/Wb,N[EWd
e>c)W8HH^bS^P):MJ+/Bf,;b]Q0K]?C.B-V3>Z:G^V^E4BMLdecVURPN=GaPQ+b1
,QU2R6];#@,H(c@_75_5SEF@d>XCTc##>OfTL?RU/Kd;(7J@-4Y:LJZ?CA62@VbB
d3S.FBLH4VYX@):9?Nc/c/S3B^0:)4M]M3OGZ;b+VFMJSJ9]0^5dHY]__,e-TW[K
FJ[eM?@R_3CHaB+::Y+AYKK)5=YO-C@AYM&44ecK5<#)YVCU,gQFA:3_7E)[X8e8
1/A#G<W\fKWHRP>RK2H\008OQVHHJ\Ie:])U)VO=)fb17\gb.-+>Q)VDVYDJPIVQ
P&N-?QN-5\W:([HU0<,W[6S,.e-e_R1=D^0e^ES5[J;R8^/J^C(eX:0NGe4QCAd[
FeI#GJ\CK]+E?6[;80RJce)W4>N80L?ZLQ=ca.(<<=Dg(;5Tg<c.OgfK<d=)S.X:
I.@5@]8#V6,H:Y=9&J:5B:Z60WB-S]<([gfB4[J@9Da/-QWfcHI]?<08FRQ3S;>Y
0I<R^b23UaC3?T6KdYM4QG2J^>+SDSN5g9,JD^=@LLa/EKCafL@<Xa;PQ:&A3E#7
A5.5SY4D@BGOI]8WSHS2SeLP1<CD?E9e\AW,W[G3D?;a-5]+Mf]2[3Zd:C=;:DM\
Q8g?Ic9Jg=W547^c]f95@IcM&K;G7=F:I[8.<dJcH.fS46ZP5#4Z@[7\7)7b>=03
KSK;\2NE=J(^]]F2REDBQFBN=S[W2Z,2L(13(CbOc=T8YDaSGHRIVc;f7I4X>\,B
Pc\PX5YJgX,,_]BcEOYW_5[L/4-S&@+UD)d&\\@Z#Z796QIg\3X\?.e^[a6W;=d&
&>LcHf6\fdO#^dW+QYJGIg-4TIb.YQJIZ#9C#g5Kg2XSeE<Ee)0,d3LME#(C]VLV
KD+&-\Z2Wb/8YH/6QYJ;OUUga#\)374gc&.ga[&YKI+@.dWa4]1aBYS>=AO@BL#e
Ma,DKQ2<;24Y11<=?d/cTRJ.:_SbZ_ZPY3-A/bW8Hb:?0.=AE/.,ca?#QUFU7GLd
C5Q/R4ZO7,ME6.DT8(^\F=Z?-FbH(]43R+O(TS?&CIba=D14e4&W&d<3fRcG8JgE
6E8SC8b_gCQ/JQb.cHf^@KW;L.:CU_:\LLDV?L9RGY6)>eUD#1D-Y3eg3>,:_4H7
_B7E#(T5(W4SWS_/-;eNbdH+X=(MEeHBb<=d&[_daX_;?H/a)/L;M?T/-^XV\?<0
C33Ie8#I]Fe8E+c6@,@EP6.bA=5E8P@g:fXQRfF=E-4U6AXeA99[?M&^GL9^gC@#
=9[>MG5aIF+<3F[BL&GD^b7F7=>K8.^\WfH=5gW3C2@UA1efJT#JLgMXVf0Jb6c:
AH>X5aFA96C=T:-YI-@Dc21_0f/7(:Ad3=0g^B#B\3]9N-[BO0g-D\+d\49;Ka+U
83_],-;Z.T>6CX1(?eDBTM27YL6Gb3XeOM7Z<_M&(Wc7@>&1,E#781M46GLJb<>+
2DZR3UCNG01>L]]@_6<\g3,g9+1NZ=\=3bK(HO6@KF86[II_>)UdFa<&?,]NVSUb
d@=3Jcgd5YOFE&J/4W??Y;bD,3XYSXY2LbB\;?K>UgW@/D.849WRXRce0Ef^(GWP
cfNSE+-WJ7Uc88g0W,+a@H5#FAR:^fMZB)ZG,dEBGKDR:G.6N7?S#/_>(0\J<O_P
VSM)DHIYSa-Ke]LWQI++.d2Q&&2D-aYd3EI?b-FD580<=((PCBVHgbTJ<8d?892+
GcK.&gT3W+]&)NTNERObE;RT<D2-YCU:Z&>Z8R.dLJK^eag7Q.L&4U]P)R:DZCLf
S(01K:PG]WBB=EM=-Z,H0,TD3gW9+?@CgF?PgHO00c8c\#5TEg_WY#gDH]-A90BF
S9XDRg>V>]/N//&^&g8Q)+FR5Ec5.9&J[/3LI^MZ1H/PM&cPU1\.K?XES^#=AB(c
6XG6]LC>[N&e_cBI:)R;7;d2(f7f)eg2N=9]^E=TBd+1<Z;S-.gf<?cG&9#dg]2L
3N7;C9L5-UI_=XeW;bAMJV745N72#1Z/6#Q^-/BF[]TZHJ1Vg-T>R2,HW7\>T[C/
b.H4\O90Y?/DRcAA7IS]1Y+KVV[aVJ:F^BW2NX;FZ]c\5--@c&C8WRVb@RAKKO,G
/1P:&<=@+MIBELDR9,7\+(BWIPB7f[-Ga(c^Mg[\7CJ/-FIb/FQg07AP5R7S(d,X
[##U&>3BRM<g@S8@^g6<YES]6g6;UR8JTQ_+XVYIM,]29[J])M+[E?Mc5URbVFE3
6cE=:>T/M)22/\=2b>\^<(=Y(M/L6<?6e4#\LMFAdLWC8b=afVD-Z=\:eJO=gc\f
&(F>44\:95P/:fX1M0LT#gCa19M3[c-CG]MgK]F-[7af;M0W6)a_(6.^GBg]C+W@
2F=_V.012LO1\b5+?Ug-/?(M6@3_[b5->2@K)E(C/F;H;E>Bdd=g+58]7LH9bR3a
NH5BJd2FfK>/bS\c(/FD.e.1SN<:3SC)e4,bGb](@g:=8X<gRdUaBJ.WPRI\bE7E
G;_M+ZA4<<0ZG_B]^R3P+aSSSSS:T9EFTWNaC@G0>>S[PY16cQGH<b0VZZ\G_@JX
^\f;W?:XZJ+=dA,:[=DGENE#/[BF(e=^&KAa#E<TC7bb(-f7O4FD]BYYUJ90#+Tb
?HUfg<]WQ1.;MFb;[+)ZdUWab\<^c@F>b4W=^MF-,1A^ca^0gbJ+_^7Z,6.(4D&&
(D8MC6<?[LHICX_T_gEG[I3(GQB=U,>EZU5]SgC<FR7ZeZ=FgU37WK#Z@bg[1@\[
QfXa<RM7GC@T@cZ)T8?[Ee@Z:ffFfK&-8@];;DgO9>Aa4#J0RO/F7Ff:4AHJV+C8
)E+N@^N]>[L>6)O<7g781Y5,]7ScMcdHgMVT<6TJQaQ6GKfb\cVE;V=FM\/IC&bB
<S_U-=N?]B^>6Q,>OWVX(9;(#^<]GS9<gDbe-\Y-7RCS99:4S7PW<\Tc+7^8\9:0
].fSOX1e,K,_:Y&e.22N)A^I)2X220P4NFC/>_8#3F@eQSORbaBITZc.N32cFV\#
YVN4Q:3f(<_B;(bZ;b5-)S861ETJZGQI3XFQ4EGMNTY.PIg)U>+@IH9P]17a+F//
(Q<T#AFNR/=:XDZaYA:8IQI,50GEKU7DgbPDFe;/C(]5#SW800D<K8@G5<03Y)2e
&#D,Y;QKcEeC[TAKQ;2E5R(Z@27)@QXae^[RbOS3<8W^f(J,NDb<9e.]PS6C;G\D
gTBVL05VQO^Kf4=Fg]&<AT7>M>Q5#.=2?/=.#+9H,UaGQ8UNL:<g;@3HXb88X5C?
_G9a#DDW7P=cNQG-Cd<ECJaT)>7gKJ/DJ0c:[#D9\W4@S(SNSaR-7b?#;.XED7C2
/6AQ5N/8K(.<Ua=A3MK:3R7+,Lc0]+#1Bg9T#;H9XFJM6.g&?^WHQ3P+aK<N@)X?
@3??FW+Fa4\A[a2,N<9J5FAQ8E8H8_a=9R1_\IB7)Q[DVCZW#3K@Q&/.YO&D+IOb
P?c2W??^2U<RFAS&6cMacG?&><aY).V0E)Y6<NZ_1V:bXBbWW?^2c>::_ESB(FB)
aIf6(_=?8,F,V=AW3TL5/Q6HdefK/#GQcL:U;4-:[:OVQ^1c0D;XS8_fGPA#&X[&
TLQE?>P8T]+#K^6?I\><V_e)63f\FL.SPd[S35c<=f>7JJF(\@G97Q>B6@cg,N1V
OK.&JcB>(7^WMW.U6;+]S[a,-gc[F+2IgY99dK6Rf6TcBAAF8N9CcdaeN@0;@APH
-41.4>\b8bW]1#..XGIUB;>?2Dc;RO31&ZcC-::HQ9#F;b=WO0#PF0aN>I?dJc(-
\Q2OV2PSQSQ&BKc#YZ6ZD_PV^c\-BB1S&c2@g:D]?cCUEeO[f-KWdX+T57U+I=EB
]R;O:7&DaXbdb<_[A)TYV.DY#L:.)[bE;F3@HKCE2_)AI@EHTW995N3#Ng#83-QR
<9ad;SFMP^M(PLDFe+.6FZ)#T>LZe:?XbT[0MY&eB&YAX0ACBd;.<a1\<G)@](FJ
)V5R(3#_I_ZZNYMaaXCY>JU7TQ__48]C^4C-gV:4e(3+f;R8LN9J<5f5W;CJ0EZE
MA73^3Y;Y(&S4\c=H2\Ia73#=?_?MDgC87g\,F(HQ=Z]<Nc=bJY]+;M&1Q3^BXV,
22?=e&RfF#6U8+Ja(JFcZUQ42-1N\6.dLO:5=DI<L\O44SZ2;KW@a]TQNgPa(0J)
3027gBUGAae](9M349#ZQR5^Ne\JL\?eZ+=?X;,eH8@)C/K8ba\P>=BR)C@[GC2,
W(E+Ke+a<#OVP#,?SGVd?=U7\20<:XcG[]]e91cZ=DU(,[MRE7]f6/B>8<MHV-]>
@0XKJ#L-dSa?7CASf1R(>^;&(L,19X^)b<8T(3fP&C.<^?J5aMFX>?8cP:BO)7F1
R?W3&Y,f&05E&C0?1:K?3PJOAT^@8A&H>?,Lg_=:CM[Lg],)3_&S5\WSA@+K#0GL
b.I7C8ZS1<3#YIZU).YL^I>.XQaAS1<D2A>W&T7XMP\;-V_[cD3YLC1H5>Y849#6
2d2]7(Q>gX7OM[U\.TZ.=+=CGdPHQf&c.&Cac7bHdGMTB<>Kd>>214_HC8c-#e[G
WB5\+QURbP5daPAF&_S9@f=[BE&OR03HBW48W=7CgRN0YEAV\=ca:LW:KIdK&1Y\
/3\Nd_[EZ,gcXSU+Gg:_-AgZ06L.&MVZfG3F\1&JYI3/-K>YXCHN\2@MaL#76[F7
)5\V&YGZ5>G^R-&TG^#/CM>KX=4d^R-X+\\4,6K++K/bgffdKFbV6;I\HUYGVHDX
_^M8E^N3PJ4<P+C4ZN/5/FLHWCKR[d?aV573:@A?J>3K)][(8f#G.TZ]=]/&<O1J
&MWHO+IXMe@0;^d?OS^DS=K,TLdc#Od([A,YD/bJ;VY7@GI<_4N294@HSAHcH^Ae
:)83/J-Yc/M8]T1G4ea_IE__EHHU7/CYGG6-XFHW4S#T.(dVI#-bdVI10\bN0,&,
P[O&gZ65fH<;aAgWZ2X11L&Y4Sf>8Q^NdZU.Yg51<ERZb<_W\)@7B&^LOa+;KH&<
L\VJWaRJ>C+LN^40GaWCHZR;[87CcaY@5#\U\QC,+@9=c@<>fR=5WC8R8\g^9BD5
M]+)FVbUJF=::bRD6>-Lf;P+OH3@Y[SQca&^S/Rf&X)LWb6J]W]B?QN+U>^QM>N0
->ZO5[YE#7<38L(>4UZNdZO[U:NDOX6);G40^7#O#/^#//M,LbNL_e0H4&FH3XX8
L9+[b_GQ;0F,N+=9GEMGFQ_J+WYK;UcCW9#)A:J#=Y0T^GW#WZ6=1Z@bT(A,CN1c
3E6?^?1#4#@f<\d-=JDHOD^#_2<cSZ;(TNfZT7=&2(;YRQ0_UFg6F(Y,_8ZZ6^1Y
2^Ub-DY[<d].DH]a3=4CH7O^T?WP:eWHP<eMcTDA5eJ#V?Ea@5.9WNR\^c^[?R&e
=S<Y]/>P-aQ6)NL(/c#RFM@GF(F-@_7BJTSOS#\ZLS)g-;9B[Nc)JIfR)^L3FGZf
Va+HgfG+K?<_1B?)M.Y/9(\&Y\XcVbPNDd<;aS)U/G04&a[+;3K.ILfZIGDPX1^Q
[3_U(RUYQ?^\70:@g+e)Kf:Z\6CN><OYe/c\:M3;^WG:UZ3_3&_0Q3V;E.&N)Wb,
\-H^-X@3_<:\,>8>:HIT\G<:6M<KV?fO:?ZE^YL-dV^W:0LFDY9_ID)9b_cG<8H=
P4DRH.[EL[X,/1K#fX^U43DTD:aW>@:aFZ1bFdNTFW+]X.T,fEfOIOF,\S/JNEO2
,5JS+OV93\_P0cNT3S7M96MbRceF,\a3Ng.Z(cZ09C^F_7fUFPX(&Z2ZDa<>J<P1
0TM-:=^^]+>CTd?O2=DM8ga@6R@[G&6#_,3OfG<K/49EW;S>MC9S/ZE\+./L=adB
H__G9+U7>>W[WRGNA51?&)R#bLaS2XW&F&3<RLN:I/.GPZ)>207dL?2cVZ/]NEc2
<IcXaK@(LG:F9PXO.)M>.ABNe19AUN99bFK@-5\T:3KPeG=3MHX:1aV1=Y\@?cJI
:QFPW:AZ8>V1F#P>d(1R\]P_P[N(e74Yg#Q.Jg=#UDbT02:PCf.29IIE;F;?^+).
\XNFEaNC+cc;F-13,OJF(V?ag_V;[0J5_?DgMdH..,?<XF.beMK4@cBcdC/cOf0D
+(]c)VYaK@.9[-fHWcg\JLaQ/eO>MGI6H)3+(fR/Mc>=/_\N4FN>UMM]c=.URO?]
\6I_Sf)fL7:PQ/)^D></G-A>+V_O<)Z&-7JGHH1\R5;8P(\V]?S8BV&E5f45&\,V
IGRG2.4KeT&C(]ZW#3;?WLPb03ZSPO(IN-2(UL-d60,N(HFe<8>Q&4JU1WA2X)D1
e=#2\0/YbNa/4UQJM>_K1\LL5.2+?FLeF)=^S4)C-D4ce9[);MJU<QJW5aDfF#ZH
0R[E;5(<_d1D02&53(NNI/Y,SCX8U^8M>_-^+S42HA(:8\\F<V<#0.T(\f\3K@Sb
I:XUP72?:[M6UP]<XFggB5g2R+[FXME;S8bS=49)R4JC&//^1EcE&/O<EH(<^:_6
_B+UZJ&5Vf>3MP\c?AaBN^OeW<eIeWWDg&:O)H)ca]XQY]1#ffg;W#(]cNc7[0=7
B5>NKBa:9g+Ag22@\gg1AcOF]eBS3\SB\IgD941E1V_dFcEV5^[1V+I7aM[15\AW
e2P#V>\I.736><1Pf0gb^PN#R3F<7YM^abD1WG8:1\Tc&=ICdS,O,Q?##1YLS<d7
5:P@KH2-U<S5;[V>a<=V./c1RfU:B8;,=d(8:37E-,X4,_PBN9CMf@4_AC44++WU
PQK?#NZB<B.cea50X1OG>;QIdLK;;+cXcL86,9?Wd^33f;J-OZI@.6F&?=J=N&@H
4YKOf^D@Z(O<bIE9Zb3M=P/+E1/LL9D50[#F)e[g(#DfZc#A9C_b9XQc>Y#K537_
TMQg5<YWI52I7V<#F0T+Gf6\<)N)8[a/Ae(b/0@.]W11?M?d+K];[EC6ZcNLC_57
<10].7#dC5VK7J;-0I)Ud[#B-f_@X/U:_Jg9FO/G+IB^a1f[eL+=2QK0?QGW8ATS
5/3A/.C91O^\UQ:N/V.7;+?#+4>E@R07XLID0;:0>PNKO09WCbU92JW@G.7Ya;IZ
QYF1JSAE-RX<6H\0G@&c/bGd:XDGNUS23A11@LS/03JXB(NW(IO1IaLMP<IcT5RR
#IQ=TPI?JN,G;g#LPP88#<UNeK-D<65W^O,#gL@QKF)]BX,=aV/5ZN,D2L=0UCG7
BL&PKET>RgLTUL^g5.5[M0_/fH[7Z&S0G3ZFZ[;P,&7_>#+2ZM0ggFdK=L,9S3UU
Jc#--.?-2N^cX9&Wa:^.8N&d0^0bO\Y3NL;HYI<3L3/YJ^M)Tfge&Qc3I?AQPWad
_HO)A#26PBH2.fA3:=@=:ZH&XD5F^#_4?M)+[8++I@6c8.E5W]1(6Y[#9)PbcDV,
C3&BWcF^6K6(6EZ=+c_CZ.UJ\];Z0OKCBEZ_;6BU++X.H7A>.9M>NZ&CFg2b@Q3b
=8>RM<G@\9=6^.V?Z\SH>P2&Ugb\F25A_f9_/,);)a,J^a@)T.60B&Z4/A;+R)7T
[:??Z^5#J-)@)BUGXb#?Fc^3F#^9I7#DOT1bRX<./-)0N[>Q3:LNdGG2KEPJ>6QV
4<4f?1AQ6F?b+0O4JCRb)9^:YFeN>Of]-.F0O,6((a@[dH\+XKY).PRL]W4,]+3L
D)VI63N5=b:\1fEFd#:P8d6D9NHF@;3W@<2<?E4[/Da:aIZ)V(N)</NR-GW=RN_^
#ZO\W?XHR\Y-TYYPNa77P)KWJ;RgT(#:/;WZ27D/(GeJHG5Xc>c?BGCbCP+J6YSS
;@WgHG,I&<J0QDd=<P/d,0N,cdR::g1G;K_=XE_R0VTZ2+7@66T_ggRe3cbU06\H
]EIeT94I/R;c:2V5Q=(0(<2D6;KDF23PB87>]\f1#FT(eg;JB3XV78M<AVf7<;)=
TI]@A-(80PUdHT-J::/8V1]4#Z&1Z=MRP?OP/+L9PA.UZD#6SM^>O0Nd2b@52S-.
BLCJBD9MG#IEa?2XJ)/YLX<+gDR&gW.;47ZDc3./10?gJG@UP]MBZ:KAY^I1B;JZ
Q>36EaYSLESOJ8Uf#3)J4DdHUY3_P6b-9WMbG#^\e4&G^>=AZXc3T4eX27UPXG)T
9VR.UfVB]eC7>fG=\f;S<:01gE+CZFfc9U]ZbR]@[LgV-gV=W<Q)#2#b?6RJ4WE0
;B9,ce0@YESIWIQ;\8BE[]SP=(RBKQPP5,9_W\dV\&>;S2)g#5^,7/f>:6TgMUU5
:3Wac^04&=gI[53?&O5RS,S+L73CN(,WA?O0#E+N,WdTREE#?45BP.X3(T2D4+DO
@E&17;&gZ;,QZY]c&_<(_3G9S1T-7S4Y)_HW82EP_9RQ/5N;WLCJ(AV)a;6@5O<_
H0YB?#CJS(Odd.<DYXI<GH7-d?8;-B[ES8I^U=Oa;]EDfTW\(EKWDe)HQC54Ra\.
^_,/I[eO.,[gKc;D3ff<9FYI>F#d73PaTD[/b#DJ.F2UeL9ZX\(]I2N@>Ee;MJP=
<-/C?YBX>fHTeEF:TG-NOMedHeF:X?.GQ#ed0HPM@R7dXG<C.1aG1bMVBPECY@LD
-_AR@ZXc7QW2R(fDNJfR?-2[90@V&T4bdE^E2b^1P0fI0QagC&9OYbMZf;aWJM5?
Qc#IIXU1e2<?(U4\b@^6F/YFfUd1DS-e#NQ.I?-[U9X^5QcQd<LGaWg\LZQ12P)e
5T=1Z_EfQ0Y;\dTSHb]8TD7M5=8Y@de3J3^Z&TQbKAS-QT8dWUC.<;-S?NQ3\(FC
.<X3#ca(-fD)@C,g&5?.JPObDHLaJ>Z1OY>0JT1#04N1g7dD-bN&)<G3MKGQ57(e
ID+^II18->RYXHENc&Y<:c#.&UYX>XO_RDBE(80\d^YLC0+YT9;Z6QM1Yf_=:\gP
QQbAM>Ng9_YYTfLCF)]+G)4HWTCV59EG(K<P&ZYc8OX;)5/8:_b:GXIJGF>BMY-:
B18&\UTYBe[)DTMI<R^MdFRX@MPeS(:&#=@^\//NKCR0dA6Y>\]L/a4&[VON#K9:
6c.TaXM3Z[L^]Me+gR5HeUeUWROTZ=RQ46NP1B>_8[,JaLBTL(gKY3(<J<2CMBgD
UJ)g5E7>]+039;^MOZ&?6S2K?(YXXCD6IYgaXX(1MeVWE0P]P\^RO^-R#AO<=T@]
87@TZ]E)B&cW[>f6PYBPVUgB/>/58Q4^EK&&1,b_V.[Ve>@A+R4a6N?S#.#O[gWZ
9,WNQJ9PaE2,K.(O.+V3ZY:=ggV_S[I9P\3E?.DX,9T3UdBUWS-T&2K\2F;:OC67
R=5CcdK5IX+2c>^,EI;WfUFdd_(J<P>N1WPU8W29b^eY@C)CMOM;(]^,UdDX.-A2
9/(+fHYYdWb>WKHBJ&NXMAW1AB?fZeIHJMF:YY?[A5f,NPb>)_>Z4BFKZP(3fUXJ
HS=H@TG>dMHa.,(b\gCQZ;9g;:Y2]-<:+RJ]I&T->M5cM45OCZDX(B+.V>I.FP88
0bRTgQMNOK\<-Dgf?5<0.C:g9ZM6S4a>0HgbZ&4Y=_ZKbW-BJ&#^RD_8=H(ZOX.F
XRBM<OG(_dAXH.(UAPg+1g=)>D-\IWC1@Sdgf)Lb_@E)&XZW\e[#TdV>YY1]K(0B
MB/gA;[Q:3Z.bAe@^gQb(T-G0UWe@]6\^1/b3?b,1P#AY.\WEI44\0J9C#)1OY-?
g?8I-8Lg/WG+P(J__gLg&^7,e;K\T]<Q2Q]/FZ-TcF8N&=<DW0faG:/NLW)^ccbf
B\TAYU_b4E]?UV<KS>/)X09+4GYR0R?)X69A8\/;A@[706BVQGe5XPY+/6C\-GY-
V&b6-0-V,4&..BQ+6^?eRC]4gbIW19ILT<QK@FTYTCf<D32g#ETVdFf]9PY9?Z;U
<5eU<\^<#K9Qf/gB8?g=dC[/RL))M#?O=5fWaR8KBWQ:,M0>3,>b.=@,#2d@OQU-
,#Y,5I@\BTb[O01P7]@aJ/RQ_^<+1#=gB##9\3#T@9cBQeVQG^a[ITeO):(0XF[c
;Ka>NU,()ZB(1QFJYM.E@QGUQ];YG4-4bdg6+S\MDOG=/ZPFg1bX);X7Q\_NU4b[
A+g5S>94M2?b;9Sc5UCQ;(X5-MQ6YH,HK+:X33]d4S8bb)D/U)-)R[58UFWV-69/
=Bg82Ie/gW#FDf6B(_()Y=U6G2K4NA<H1.,2(I&K28US.=&/45=#dJ7O2,3250(H
2gPIG9W:ISW@3&ZHYfY:DA??66IX.;F&+Q26BNF.?DSEObC0f3,cb3T<a(U^GbD:
B8=O76+D#WCAg9]0\LZ:&8^0#K>&WCeI?;\Fb>F4J.A@>aDX/UaI?f9SCF\Q/F<.
XG?;J6Ie_,^ZU:VYMA.K^+e,g>d#YU_bb<Y.^>?6bL_<MRHX:,Zg,_9S9aCLFFJ.
.S(Pe0=>;T.T7,VK^2V8^aPUP36K[\T;CES#1;DH+99g7[aW_1cd&4#XZNA86<@_
:4DQ>Q6ZC7RP#JADG4_CU4^S4WEdT._ec#e=;fQPMg0-A2c01eA/B=ZO?/g_1WL5
9[Jc-KGD7E^Y4[Bc7NeQ#FfPER&AF[T6M0eO\:PAQ<0Bg29X.bd0X_9ZQ]R>&5QZ
Sb.f(N6Y[/c)fdTf]9)Cg1G3feH/cMU6G,._7A]f_2):\7WAbW7_3If]LYNNA^c^
A&.B9CRI1]eU<C:bNKZW&@-#5,P-NK)-PMa/W\L^B.SBgaQR]75E]:fSV@8)/U()
^f6/.bg^)^9&^-HSK&5B])D5DW0UG4;f1=JE&bY<aFf++/+29bWJ-Mf0P2+c>@VR
aYdPE5de]FW-gfG#d(-T^]SHPC.cF;6@#6A6B?=1C6d>We\71AgB@_)]A\>:VKP_
=ee+VM^92VK@H;0e4R2H.[g&+UC7(LH/S]#,<\)IT_<=26\6\>@N6BgF;S,a^9]g
Q:16_Nb7:A\Zg[<:Og>9=;-F\,eK;HS&&=;QC/T1:?fWdR&+RfUBPF+E:XLE,LeA
HGJa,&+^A#8RRT2S:J^FC#3O_6[XPO(-:-)G09X>ADg87?J:<d2=PU8/9<eRD)d\
C0(5S/c1U7[.@J_RN906)>]b\E4gK\6AF:,GU@E>H[_66W2b:YfY8YRUKfM@_)>&
cE.U=Rf_aZR#)cQG23:^X;-2<C+=72W),89QK]@Sc>N1P0-WHM+@J71<9XH.3I_Y
QL,9CLQ<FF:S812Q+FcN>?]-^,HF9:^]&K#)+0,U2BX883+K)Mcb8X[H\IKUd+KB
6IEdMfOSE6gYVG(L)/@+ebNYNM4WCb3)S>,,B+@@ET::Q(.<Z3gM3XYI9gXF5,BQ
<14_:X.-8PBBB>Fb#Y.(9Lg#O5<:H^0Wf5ETU0&SXG8GE]\Q::O3BONW/^KVFWQ@
W.P6a6KQ^\G.,O^4<ICJ:5-e9dSQL9;1KY>&W7MJD/HU<ZZbQ/^_EbO4Ic7YUGB4
(g&86#SD(D+Ha@?8+?PYY4+?Ub25NE:=:G_OM,S47(WST<\Lg[Ec&_L^fZV9BDbT
ZZ#bS2bb2+c.Sa(da4M85bJKK=1YDgZ8F2S>@=Y-05]G0M2&+;:GV2S]#W<O/COL
aZXa&>[JV:9)G\#IXHOEX^;2XKX0IJN)&7@HR;QIZ71F1=3?^bYA[MTR+NHZ2WK_
6V_@.0fgNEe2^9cX/B5Ia:T.45UdM11[)^O\K8]ZFD;Y=2FXbe<a,SUeK.84b?H5
;@\B-:.AXZUBRCc(K?(g(]XQ=)?09_c7X<Bf,QB+^BPLaH[]@;7@0TJ(FPa9/>^N
R_f53J?]48M>ZR?S4>c2EaSEd?V&OST>/?Y9c?&2]\LF;aeS@[=^2YeJKZfAMU8U
d9^,fN0V<#OPN?<(8dYA6ZAE1=75F(P/NK3(5,3^\@AFH8H?:M#R,HJ[SX>:?>LJ
b(V3ZCcc>E]U1_L9AA]9W^D::1J5AFFAI<Z?P:HA:<YSG8RM74#cf>9PR&CBg;a?
V8V0)a?4.=UJJMR-^_&[LKYXCMPdg/a-2(.4B^@a-BL:@OO<ZJ:CNd((gUXXA@<U
E^KP?0([4&L5_X(GbYX?\15+e0P)8GU,(3J/Q@V&6UIc0\Hd?O=OD7S)O]NS1@bV
-KBGc,ZSS5D2eE#_5EUgK+F]@KW_TUG,,d[Qg\7X4Z;A.;[PF#A[L3-<MeFN2:2f
:GV,L^GPFGHE4cObZbF_g_<aa4])(Q3-<.)4>f_5eF3)D<Y\Q^[Y?L,fPT4U^e,@
:3IOd_aRbf@ba;UE\T;X)+)G<_O(?.(OGMX(=O94]I##4N^#Af/g9TD+=4D[=3HT
+LL[eZd\Va\KF+P[PC==TO1Z/;L#E7\]9BgV5aPU>/;V@d77</@9AOJ?SZE(]V@.
L6aRVab,CU#3g>1THJ;[[^?&c8#IPA&<E^,=.62,B2B]VGJ2]gN]WER./Z422:<+
KW<]]2B:Mc\9F+POA;_,\_K?_=)cIP(SXG9+YSD@\G9WZJA,ec(>K<+L0._e4RX9
TEf=Q2FK+S;]D3JXOaa]6>]Og.OWVV]=,AU1cK]a=R7H(XgaBf3-bd#aFdJP8K_a
,OM&5<&#9<WM3]X+0&M+RN?aW65FJ879@MP=/+6<bR..>)489WO66BLLc&[\XD]T
4JK+9^5_)IT&9MHDMeOc#5[M(+]d:eDB[DBV\CR3]2cgET8HWWRD4CYI-WHf.fNX
^ANZH40T9G3Y^)-e/I.Bf^WQc2TK^X>4YF=T:V=-Aeb9)94)_WD6&@7-A(ML_VdI
Q]<2X\.;_?H4b)LHMZ513<?6LOc=8P61]7:)?JHDFV895S9fOV/#U\4?K/06TZ3A
9ZeTDc89C@S42WV6W?DYKb/MAO.Q<K8,7EJA?BKe&QA@:S(Y:^_O9^E+PZOP4&#:
P-,RFNKLf?<+JTM[5^:C#:?3@6)FX&<Ug7SP\DY)P,):CCSVcWZcIedV(1C^LUe+
=3EQ(\3a2DHK=31A?9^K(#Q=<LPR&#00/,Gb[:Vd(4/GAODN&C8R/cZ0FW+^2&=M
YZc#P3gQCH\gMJ51C&Y+MPG(K,.&<FeDF/FZd+:)_FQ8aT#7GT:da]d3bHJb67Lg
L>]@G/]^8R)<Dfdg(-Y7bd&UfEX-@6;UO1AK>QA/.14cf?Ve:_:@+dH000WZBQ_E
J6[&NS@2]/b@N</SEe-cQ^OL(e5>3fJ[,>GZEJaJENQ56^5Nf+MT2AbQK?eKI1?\
^AV;Q9BM]DXW+8d=AdH(Tad5NN80OdR#\X#a@GMKK>^<[&92QRAL7/=><25HC)C@
PL?Aa(,#5-ccP4.eeN<G,G,O@0:SEI(TV0ZTDWK8&W;JOI)0QP66IH0+_M9=#\OE
8B0eSN/BOU\1^D(B.^?);KV7/;^2#fCd^&?JW5B2D0G;44=&DW2=@]:R(GWg:,V-
(]e/Q><V(eK_SO&,E<F?6^:JQM?_C6WE8:F/UI.ZaCX:-F?Z>TQU5_:Qc#W?fQZ1
WC,Z@328QFG;3\aA54BaTI=/4I>f>@Q:Z(#:51bZD3cH<39NX)AO:+#fZPXE4O,C
8CSWA10Ve7<@@FBBEEMF,297X#bG3US3J)B9P1\^-142<VYeMD=\UB=63bRR<g6O
TNC(/.\.efeeQ?2NT^<<VUX&_BG1aGTg@SK4-T?)cXZGad+E?T^AL?H4;B,&^F7^
-DfX]VbR+3OI.<J^?]d]0X43UcdEMS11d=]g6JAXXNI.PM#OK=f[FSKGTA+@aY(E
0#:8U1(d6<M05-dFD-@Jb&+O.+9agaWdR=^;Y)D(eSD\A3@-(V8A/K+bMXPgW,EL
1P9.=J>D=_N=FL_;S=/#H?DB=A)K&NY-W-:Xba:;1#N<Ga;91?8gX:_8E6(aO^YT
V.5DK+DZ+-:aA<(J49VGd7\6cE]GU;#P3YI]V8Yg-/4,3QN[.Qdf,707M9)e9OE@
B(:S+S5KJ4eL(V?D^OAK\gZbODFJa[>P&A+(0;E(6HZ;0\J7VG6,KMgY^(K]aQbW
fD.YGb-7RgUa?M7<XNKd?4GUT5(]7GG]T214BQZTe\2/GA_&aGTE=HGaJSHcDRK#
(3M(b07>-D-Cd3@U)F[SJTEK8fX,TH+VNX#9S(aP<.:^HcLD5;Vc:J?e^e:=WH>B
&N,,):+Y&U+PdH4;4-]GcN?,f0R(:HP&MA81^-K>N;OMX2-E3VV?c,1GENgN#4.(
K9;G+&-FS178XK:838)7ScX([a57CeTVR<)C6F7I#FCV]-2W4c?P-@23^Ic;f:@W
00bNJY67aJ3OUK0M?R[3e73H(KQ]M19UQVL8Y344GMQ[^T4gdG?NVN-NN.WS^+95
]VG-WO3\ITYL89-Zbe;(O@36A@_)GfQ.&+#0TaK),aO\7]-f9RC-;&aIV4BV:fPN
f(79Mg>E=MT1+)QX/3fKZ\J)Rc.D:g[:f6c]<BLH7K1ZQPZ-^>Y^V[;HANX_TF<>
:#22.[@6eH&\,TXXGEYEaB0Y#=\6FB&HX@9SNROc@\J+a<C_:?1Ua@f;^3A&.XS4
caQ^@-##;fO@X40MEUV48=g+Qe4C.VM1B)>B<Xa8<gW(N<XJKH_IHB8=ZcbFNXP_
@ReQ+;F).?^.RGg27gBBM]G#[OO??PYF15?.A]P\8-.FAF+U-JTM2/X4:3J3NI1Y
>=[@4WR,J;Y3[7;4-#PLD_+;DeAOc0)^H>,?gb)[f&TJUAO;NR_[P;(I.g;HK2C2
PY5bOWGZ5<3cA\4a&[264?A4DHKf/NT#SZ+15>8NUg:R-1>;)L6=]JfLf[(OaH5\
?U,2a,2AC5:Ofb/RJ>)Z8VeIK#Uae\cNddgKURMSW7Q(OgJF/N8G0Y?;Vg<UA;IY
@F)0>:B7c2-dU8OV5&F,a(177J7PT29V0:Y&Q6S\70Xa;DcHK:;Q=M7S,AYX#2cR
:1L@4IVU@4-0&-6;RS(@Z(@2ZW->W=dN,C]BJ15E;<;Z>9R9fOQgZA.9>P.?WbI2
._?@cg/Y5^S4gD@Yg189BUaLUQB90,[OG@>)OS@Z)9@U#FR6-7.Y.cXVG\#R^aBd
PTY]7Y5+#?[\We._EGOB+a)6G0CUD.KP#f10,AXc]0Q2.e6+LEO9c(He6YbER+77
42g/FN?gb=_\&Y;[Z+BL_:XE@G.e=TWKKacVHfC-7H;/>UQT3R8=1fG@,:Cd<#ZE
UI#5-.g,D]gc6W06PcbF]42#De)UbB6EUYR-34+C;;2f/O/UYM=H8U00M@RYO#a)
<B?6?<GYMG2ATN&:-B?(+Sa,_]84S27e264bTFSg)JAVHZf8:Ec)9.[@..E+EaM]
HHHE7L>QXS@Saa3#68@6OPDWcNDMD\=#DXWd:2)?E@=;,<Z]N7&3V(5RN&>ILH,R
\B#^JNCgJ;J;ZO_)A+U-9H=eg7LdR=T56C(39Z]^J9C3C=SNP,_QN^\AS8FfM-Of
/]9^eCTdPa;-Q6QE8UTS8F4Tg(&C-)gA6,Y.MO>0CH-#>Va[Nc^a+Z65)U^6(f5#
BVVKBeM#F)5.-GfF[+Mb8[7A,3EU#HB@=-KS>H<,;+5GB&&;FN2S=BCUaSKH<<NX
Q=XdY),4JAA95DLgfY<:^Q9[>#G:W?O1:1(MK:(dAZDHbTg_AO]KL>&W&VU>cE?+
#?_/3bT5acbcA.fQ+H8L[2cb#4f75RKCfHE5L=T#CVE[X(1XM?JYA1,bC^bPX,X&
)9_QN2--7<fOR(#RKKYMR#U7a+6-a5-JA:)f_FF_SdYTFa;?@UQ.f50E-@A&#?eK
.&GS\C@EaVb\M.5NF#5g-&N0.WM(FDM\2eVW^G+,7f\&>f^eabBDDQ3H46P5X_?B
9/1)7cG#O8HTRWY&+R]KGVaJ?1DIQJc#BcB</.FHRN]\A2&U@^A?FDK?U@,68,FJ
VU:.W5X,C[B4;]+:<2?P&4=;DJ0I.NH_Xa;M+6[4S(QR8ZB;F=fE]^A_7UJ/9+SA
eTFd6()-2YQ5;bM4FR^@a@^&JegVDed:37B##-Sf475TY]&>,TD,F\gB=,F/ZJL_
H=Z2>3CS:5OgEWSKU^aKg\IR]_I;V]d]34B--07Pa+]#Sa0gIe7JFSV_4LZg3gS]
aF2L<TE)KXN2.L.b]K.g1FG?Pc4JC#Q#=@:Xa<5X<RBII&#,X2-A=&I](]8D++^+
\V&C#P(]TN;He,Z,]VLab8E.R)58dU5RbNg,TW.MdW,daA;=VFS8(&V4-YeKR3Nc
,MCdI4H^8N,G]CD;M#cL[cI&OVY&.44IIgS9)WC8,f;:,\a1C)X8N^_#>eRVHe0V
JS8SQJ-gX?21SBV_,QWg+=?;-Q-f8ONaPb;J9]KRV4YcFWNDJbCb7#R\P.0E4LFE
HdPNgg9K5B/TCVO780KVS_ab@IaH0>I;GBZY<?&4S+&=V[;WJG2b214D+7;UIf;f
F]Q-HQ7A/_C<XbcV?XI/[P][Bd7gV(0;WZ.>T6JH4K>;\6?L+g0V7Tf3_M;)P53-
G1641@NGF&O,SD);VO]]]L>:C\<V-IZIYN:/FN)>1_#W:XHQd8>38Q;?][@4J5FJ
W(?_W7=26OW8J(cZX^72E\CK)@7(PKA[Ub[_DJX^K3&A2(J+I-==>);NG;4QK\84
6g66A;O3F_dCS5D7T(OQeZ->DI,A##WU:P0J(0R@/>[VPZe\@aTEDI<e^R:X)Hd8
JK/&a1)F[\RfH_E8>1DK=,WN0/O0BM_UQ&29:=BY:#Qd>.VUYF5-cR4A&3eOg6#g
(D>=(d0<A7bB_:eM3CMU/-I_5Pc8<#dW<?fM9PPXZ86B>[H;T>A]BA&-&2F-4(FQ
S?J>075DcH+&1&gX7\_VN]AgN(X9C=8DJ[+Q\PM3]I4fL&@(_P;[<A-WeN(g(3Xa
f82=1Saag:B#S\5(&.:6VQ_IC2b_F_JdJIR.G=\-,/0T?E>J?Y1X1+PTbB8=#6f@
)V#+(7>1L38(I\VOF^#9fg&+8/KS&-?2=,VNE3X#J#SLP,OS<F^4@IV_>eC?cZ=T
]\fd\6LNg.\^MbDR1TR.IV_\P[KIY\(2L\&X-?[UcCEBG781YgJF/O^8]HQTZD2Q
\.Z.&g>T,NY(67G>&ZeHY4\/,9D;774fS3DTO)aLYA,\^Z.3/gI>4BdBc/f7Z#M0
-g[ZCVDPd.Q/]LWaK/E63UfD,S+S@<F296R8,IVB<,P/2],ULEeBBCUJGPO([?3<
&7)\+[Y&W@/aGH<]DZK-POKdWdE34^ABCP@)FcI^EFF<-BdYP^^I2?cL^/-^S##Y
K&g5a9>;8)cCN\^CJ=HZ0<=_B[V9N60-S4QPAf)W?f,CS&VD#W1TF&7aI&^)3_bG
(9Sa@e-dVZR6R.[Tg>C>QK^0+f(H;TC=AV8;?gWD1K9QBc,V>3.]Gd]J-8RA_Ud\
<:d=]=/,BN\bJJ<^;Z+,UXNfN_1\a>>O^V.<^^<3Ob[6eJfJ3MLEZdN_4\KcNRN+
SYJCc12G&bDa.S)G;D)dF,:>F4D/agX<2\VdfPWP;Z3+]/UZ47HH31F^,;AJC@@7
-3^dW5/3&cd:PP_R>/GA-J:G>78ND+dGZLT1+^AK@d4eB((TETI^(TUccG3b<_RS
Rg@K4-5S8OLZX?K;9^B5;Ng29@fc-8D)bKDa,@+N1=^5D4&>gUMZSE_.(ECF4_N2
)d\d@/=[&K@HKaG4:cD\1:3gfX-1>UBE7+Wff_VRDCQ73JIEdd#_PX:2+,gH#bQG
[c3f81#>;?&X&+V+2\9IU[3Bb7D\F\Sa4(E3&Y75S?\)-;<+P55U-gfE,G539(:c
Zda-4@;+gN3e=Xb22<^.Qd>W8eXPg6FSg4EA_U4\PURBAGefEMYHJ=Igefbf8NfK
-(?]Le:8:[,E?1bNd0:d58LTX#>f@3@0Y@E--f@#/A5CZ-P9f4eT4I\-=^R:^Lfa
TQ?e(5cKFQ2:(RU.c&bAG@?.^agcNNecXLD5V;\1#SX3M3?c^MI0(9dU@U<@.+7R
_RYWAa5XLS;DE7GJ,&P^QW;;=J+GLc8#baQ?G?Lb:OE/+4P72]dGQ,-&A@<Bd]&O
0I]5f92#UP@;b>B-IAMSJ\KUE;#1ge6#b,EbVKA+4bdET6/H#gAL;5V#;R=:TY(:
9^ZW3b[DBSD_T-8R-gMcN<13^-3]P9UUXgLe>0C^OOe;IFFJU,>69LQ2ZCY35RHD
gK+U#aJ,b8[NGR.YG-AV2cM^c<1Z.=FH2TZ81T\G,ZU9^XfA-b+gJE@3#29>d]fO
/&EHX#3HPT+K9J;bL>/W5SKXO?<#:U[06#DG496bDc+I[De5MCQ?7?H48;TYQX_U
ES>A_<@[/L-_Q:U(81(OFP&6P\#SACe2/;LQDQO[C0a=96GZDNU#HZKD1<g+UP(>
g1H:/<7G5@99^09A]eRD6,01T./SSG:ZK@_T1+V\C74+#/WV1e/EU@f[J9f2dOX;
eG7M;1Jg=]e(EUCc+[FON=BcT)Mg&c=5IE:CN6,,(>MB#SB&3]2=Bff:.MR;=N2b
.NW,O2A4^E0./=FJG@c6=G,?>+a7O/K^^;7,O>R^4P>2M8;)LGc.964(EP.;&dZ.
eGY&NWJQ-H/GfE2KC4dd&Y93Y4-?=H6;9MDVICT]^EP/9Va164gWd5gV;NZ,9O2V
\0<b./)3B&(CG8Y#F/324\A;I>^RUAM=I-OOT.YHcP;]gB]0)a+gKd&(BRYZJ,77
-32&6:8K28<>OQ:.\^FEAH23O<5D^<_YcFdfHRRR\,:?#Q1bXT]-?T]Z5V78f8e-
gE3gUeF;_YQEI_6@)C^a>MJM:\=ZcfZN8-SgG,OB<Ad-4XI-&Z?83Mga[bJC3][T
G6,_FC0@PSTI>+HV[&-g/I8_X9A2>ObS4;bKOcIc0X_C8X#\G]P(BOV#D)=>8:1f
-A<Y;(IE?5f.gIa<.bF9#bgJ-<FV80R/c9;-6C=V5GAN;F\H8a1cKTfK_#?YJ]LR
^\BP]0:RbafOf5,I=:[&=R4<=8^B\6NNJFV48L&&e\W<^/U1K2=)N@H63@)8,<<6
,PL<,=K6_(Zc38VZ-ZYJ5\Z4-SKY):28IL](Q-M_gf+K@9JD+S_\\SJ&M\XRIO>P
JB.N(B_70/>@@UC?(8b[X:Zf->NLg5JAH,+bL=+7bY<c2\0XP-W<2A?bTASe2LE[
VMb_?986L+?@=_>0Ne>UA,E^YZDZ,E+^fVVc6L?68_4QRMR((.5TZZ17/]8OC:^7
<ZVA1FG8,7>KLa=?4IVI.(\L,#]JJ3;faY/WZQKZOL[F7M[YD4D)+S=Bb<,Y/#fX
XLQQOffV>NXdB5F12_F=:BYTQ#E.4,J1XA_I[bF79MATD3[Z5HL&M)P#@1WL0X>X
/?BP4aU73W75:><-X50E:,5@G)XFC1J)Hf6;)EI/YcE:(&TeEA,03EbAS@I:c542
cQec0HX/-J^ecH#\Q7U=/.5R4Of_-?&TS:USB5dLDMK[?/FY8,7(AgY5G[^)6N^A
gFcEZ:VFO-M?DB.O]Pc9d(9&aFFU#;M;H#R=G4U-M71TeN32(K&<7G<OOCb?]^/Z
_8DCNQdUFY6C+S(g1EG+E?EWA_^^7_&<21]D&CD-LbTC-ANc08P1cT(]YW]QP&(g
-NEC?d?XYBE8@gR.QW31Q+,GbK_9QVDZ<2>b#)9Ygd(1JBW2IQ)PBI<^U#6R:XeB
df5>1,#G8&&=5XRIbGQG75[[X\c?+M/.H8FTA4G1ZS7dT1-df@?FQX\0^eX02^DU
ZM1]=f+SKFQdV9CP#XTfKXO@,HL8?L,VcO(A7a7&UBT=(2KY00\5F,Wd33L:8#_9
A-b0/8H.@D[6Cd7P#;;cPbTFJ7gTcAIW]:7;Z\U/U(bPWc6IF^8M[MM(5)ZL-HC4
YgXDO#^df=T48QXYO:[E_SSNNgHI/W>#Y>_>EVP#^2-_)Q-H)Y__5M&c3J1@I^dT
>d]=;3YU]:D+fK&Tb?OQZ#6&>56U8AC?_W>JS5J0T^_P5(AF,^_W50#N3SOL^&,;
[/cL]U-48-@2H@6b6P5W165EW(90aLAVSbdFO/UT_/8GVI;::A;<ZWG\QY\B^;U[
TC\AB8J=bKLf0>1Z+8J0=,B<RKaEb.d0]W]:,\;\,225V;aA(9d@,(8@G[3G1gO^
9^AG?/ecO.[C(C?>IBY,fKgU(MNEMS/@+e8Ze0g-3<&\J=/]2ED163UU7,4c:bV1
]SYaK(f/Ae\Ma7Q5<2\#d]d=W3ff4b^I@.bBBb=]7J&0O8XW<&&K&TdYNE>WS3>a
C@<6BYP\QM[>^QCg8g;\@1;;I_c3E@6e@WbVGBV7/R\IXPJf8/?#@^WI_#GC]L/2
A^dC6=>;@QZ_QPR;dTO0_\G21b&QUe#NV^U8K^P:5_SRd\G\;WCgPE&52ZA^^088
Q.Na7TgZ71_,4\Ab.Y@8TTSb8f5^>7MES28OAKCNd)WM:5.3[aG0;W\K<N4@Qb9&
/+9QTM9E7G.SV:&fX;WbU6D^OS@LG?TOeG.&O89g-:TdEQb45aXC^T;53VKc.,J<
?dJQM>MWJPMWG@?\I,A/M0-[;02XR-PKQW4DA(K)B/T67@:67g7]G?ac<d-X7>RR
ZXIU=5Z]CVMWG^A]V<M(0_>:86C\9Z[S+JU#LON;NIdZH2Y0(K)F>(V7RDeXKDCL
MGJ+D;f8c^P]\0:dd&&[UX-3/6_Q;;;,^W_6d:0XSAc1\KfN?:a=\>1)5;X;5>f>
MAB23#([@W[gVJ.7YIBBNc0ER.LCad+R49@eP6g2[-JK6BP#^XE;(9\BB:,21HM8
0@EJ[_\Nb78@CQd1A1e;MF^+C>C=++:\3?A9@LQ#BS[2]0@I<bR5<<eT#cT+d[8E
PSVM]#J=bf&(=@X0GTGB)<&:O\#eISC1ZV:P@8UV0R@,_KM5^>3:F7E]K:N#.]fO
&Z&JO.e5-H+9CaPU6/=]JK<-:_X^M/1+]3JC^.gDICWJ[:gARY?2LN,(-bY3/2bY
C]IYH9\FN\6D[C=)7-KLXN;aYS79)#Ab(aB&#=e13Qd/K+e5&M=_CM+0NJ:VYf@:
1/Ab>GLHC[BeWRON2ZdRDg1S7(0.LSYBKf7@9V);Z>Ac-@UZTWU.OPOYIG?L,BOL
.c2Xa][>CQRH9=6Oc&cYSIa5)R,TVg-:6TZ&cL422^.eb?gP.29g;2]3]MV1N\G7
WSW?a[)H=&If]3K)A7gKD#Hgc:H5JaB+8F;ga6(_V1H_<^KM+a32:2Hg\d9[?7W.
/=-DA9LN22@H^QfL<[:6K^>OKFB2;9&X[0B+N+1.&].YNLgaP8HH3Z/:@E]KU#+T
8^\(QM3UL^Z4MBA\XCRRDPRB4MD[3,1gSBGCbA,NW5O?HC@g_D<aWL#e8^?=gP5d
EF1WGg]WM-8AF52;_XZ2_=0@c8DQ5+f.;:2b;NLL1c92<UP0X[1W#<a1C^=]J6Z2
Te/g_\V,-]S82Tc(gb6(F+OgN87c/_dL0gP2.Z-+/O7-T;D>W3BVS\VICRM.HGA:
8YNfWO9_C-<IBK(YMA)V-7b;0(.<THP/1O?C-T\SNLcJ075EO-<ca2>5&M>bgCW&
ac]d.U29<L[dIOY+S)bfV]>N+#HZ4B[,U;#80H9ZfE_GQ^eDY-fW._BFT&c?X3?/
62OIWbcN4c1F\IQK;&e>FI=E(Q6af1e.J3^_a+,K7]H,:K#+FE)D1d[1[#UOHP\\
Kg#\L4S5<ALCdf@F=H>4.3)(U3d@c8DQ5B)4R:cRY[8G:E?/UF&fM0UT46KNfZRE
3,.#dFJ9F[8-P@:8a+^8;#=R1E.\\3TW):R?@J;UICCS6>/6V^B?ETNIVYUZ^S\N
D=-2C?H+FBI<U21TQI/FY2ST_FX:<G8(8QEJY[[WLZ]/f&:LK@0\5#&dJ07.Y>U1
Ye-2Ud5RUSOB7Y6\8:L?TDUA)W[]e\H,/K6EgTZ_7Q^@NO4:\R.Pg^1^.:5+Qf>8
3KN6>^;6V0&D@-)3SQJAdBM.N6eLg,<XR4=B&ec4@=-H7eK5W[WO.()K+^eFFX,Y
S\3WNg]eZJ1DHe4QZV,(XO);BbYE.Af+@=II4C;V>&/g>7[eAKV8QY)MaB<8R(KR
;WY?D@<eb5a;^CI82fAE::G;3g.[F/T34=#Y3GX[8/:FGFEN9<?&&Oge)dTI0L]/
XC)D3@4RR?12^CCI0e?RRbL0O708V0ZT_BGPH9^S\3SgHLB-F+2XA@Qc>)C#<eQA
X=>@85&?._^DTH1c<PG+3^3[gg)6(&KbZaAJ^8-X(Qeb:RG6DW,BF[/_[+b8-&S1
QNGX<#dP\EH_31_a6.d<JVZe@0cBb][PQ<P+4J4-eIB0J+3[:e<X(SGL.(E#=)3c
YKV)OL6)9ERT.aSf_^_Nee^8e]LF[OX(ZC:9-HBf<)V(>OE2;WN?7G1b;dZ8A@Y1
^dJPL)fBK9[Ta?K+Q=FgKNW._Y_=LBZ^=_MEc\R)@@;-cW<,I\U0YVBMc8Y:2SGZ
N6&5=0?<f2IR_gT@bC[g37a\=b^/>:YMPBgZWaH?2B;5JC_:9FAVA[YOVG2>Q+eT
3]aJ#TVG95VN,:TFJg_11GH-e)Aa-<V_fAcW5L#/J[VZPLF=QS4YfBfGdWHKd>ga
OZ;=d1gA#gLF&9<0DJ[B0=d:47KB?Q)bB;WDIe.PCU@9dVQQ)Q]0,>+@W)b=>[6P
53W2F)[aYN2ba:47?E]&6]./LI-[4O6&1<b[O1;PMIK#a[gcbPQOX3Y2\aJRf#Rg
@fXE./WJPV3.:(W9_=&1MQZKMRb&9^@,O+D^JP+?4W[KP+T1+.;0#a<dI;/+a495
DVL26SY?R+[GLX2R(00TA36K70#PK[XTB[U.EV@fgHT+I?@V?^L:U(-c;K>:Z<6S
dR9J[T7.5?9\ZAGI_F-F?)[.C:PMWY]\2R/E@JN\8;5WIbWC:W4J/4(9)>=H_QZf
bT<VSa:28<TJ1ZHS#QDa]_[2=A4538e<M]>F8BK@gX([\)WT^\@L7(Z]:IC^\Y3K
1=FMeZSP)6Z1)0CQHg+,<g/^X;aO:2Lb?5QOSfgDAZ57/+E]>O,ZFKEDZG1ELV)V
?;8C=Z-1X4fJ6@0]C2NA:/g.;YZZL0DbGgBfN)_8?BgLEZ8Y;eON,X0bOLYTA,0/
=J6dQc>X)a5]3,NN_bfY;g@fb@Md<V,0Of1ZQ]RQ.IL8;&@/E-+\],@Z,VW=A)UT
9_U1UDfP=1HcPf#YNE@L>DT<6PJbWIZg<DSI\W=DYMH+JYZ=ZZ6:0E12#A(3aY-[
WBO_?WUH)L&cF8T1[eHVe,#Nc^19YgNfcdQAgeW(.+NDSb7/d#^0?3[d]+Tf:_[d
,B+ZA_CGf;6#Pa/D^b.gR3CF9?4@]9-J=YQ.MLP\+:+-);MGVJP229F8Xf#V4(C&
MHa4BJB(4E>7S-A6D;e9LY29bTgCU/3S=ED1OJ1SZ-Ldgbg91<eG0W5Mb/I])fKb
6c#3EKLQ0@JHB_T[&K3>c:>-gOG(,H.#DHKC[7.\g0eTQ<^efN0a:\K\TE-ZOG,L
B(cR<LA?7b]Z[:@S4a(;GO++S(3^VKBBS<6K11cgI_PM26=6LP4JL1A)7ST0QB[S
>&FL9-\]W1+;^J32ZK:_&U-=.<a:BMLPQ8AeSL0[RJC4gMT:G\E<\T/O1DY4HG/Q
PH/Me\DP1OZ/)@E9RU1XZN]:,9dZUCE:f6JYNX?e\Lf[R@1B#HVcIe:]2_;COP[<
;050Bf::JJ^S.HQ&1[&ZSL_B#_5WGEK0W00HNEID[?/U@c;HS=<BIVb0QJXS^&0C
..79W9TH4S<^[0b,SC#P04Fb]4,@\HU?0(^gHNA[C#BEM\@+VP>W00f@13UF1B8T
fYT>S5:+11+fU6Ab6Leb3QC\OMGU]N^6,eTAXd<[)^AaCFJ?N5;.g(_94>V)#K=A
0:\LQ9_ZLKGAHJ@QIR&)+De?/W(ZC?,._;8;X2\-LNULDUKALF5K.CSC/H<#N2:)
U&F@Q,N8G=5ZJfK7W7d[^?LHX57)5?VXFRVO2_?E.YB1<YOAHa?BEc#BQ0R-B=88
?(H]2XCeb^F&6,f6PaI6=U1?KgL#WDF\IP_bTSK7(gG;V_JHI/aRge[SG>E/F-6O
4>R,<?@@c8RV2H=J84AS8#DLQ,<N7FI_78b-4I342S6W];U]&,CQIU5WD&9POed@
6Ng=_,gSdU&S9SPD,eOL>G.G-7Ne@(^dN;\=_??[NP4+S>e?=3e.EFG@/LM;8_7g
89+.Kf87\\3TPFTR;N=V9>(C<K8QE/d#Y#2:D)Ff9SNeUKA<4:VSX,03^\PTLQ07
PK+Q0bT6QK=>A6d40XUF.4<:ZPFY3?/^3g85?.ed_>HNTLZeHI8+]4A0G(M-)_aR
PKag62NZBE9Q,##g#2;@B^^1)c+6c3JLH-NbT[ZfRg/@CQ=+MOW/J-Bb4Zg#/1-G
gB9f@LHMRN1dT\c4fc#d]B\>35X@<FQ?3E/9[?ODE5Z<f@:(.R@e3(1OgePe(eQF
?1D.V+WU#/PSZ39gCF[:[,8T4YY:^X8_;e3Y?BP5(E-O+Ta4Eb+(OfEL3gefCFg,
5F?Ze69><]SYX:6>/\(g[G?2b39?ATGV^3J^)7F1c.6;)Q=W@1^?Ra1WP.(YRA:L
(X^f:KM)[a#)FHFegJXWETWLN;2IIKG=8H-^KKB@6Ld4,L;W/aJIDb=64M8\7;X5
,L/LLIe86#]KgfZDf<a@Q]Kb5QEg:G/c#9^CcZbWXB+F#CN#T/]WYM&L/eZb,dcd
IPce,2BGb5&M;(?2IQc)cB_A,_>Y[P5((,@F+#2S:d#d61,aKN.+A^f]V;bLX)/G
U-7#/93/TQ3@S3[J.?<QN;U6;Q[MG-M]SKc-(]eC<HOa;AYMF##MZ5KT/5EP5de(
#,I-T\_E8,<^MbAY0)UTHD_fP+[8?D)^N_))RRM6d&/?\ZE?aUZF[BbUQ0XRIGRb
@f-;<3<dFTc(2Lc@2F\,B5VM)HY)\QAc_I]NT>bEIL)^a0@&Z8e0F#fBJWR=7.AS
XEBZT.:\MES2O,7<?G=Ma(-R);-T/)H&#0#5-PP67dO<SJgG^gd(D@SOI\d6.K.)
:8eE0K\@4SN@Cb9->AHUCfHEPf?HZ5ZHX/-M_eY]ODI?Scg>eWf[C;+83LV:C\Re
egI9NAM#4>(@[Gbcd.):Z?eXUVO-,UT:/18]8<<>HDK:bI90;]B]IU0CB1L2[G&S
\>DCIg,(I1&)1G_5:UFP:7eC>(R6UT1)Kd8aRgd.DR;C>KHT>ZCO&NQ;EHEFT<BU
9eC.?>XE&X@G/HDR]N6]^<C8d\+BG7Z9AgB^_H:-POT4UZ^=\SK]PW4HA]Q[W,P=
;;QB>GC=We5L(IC,ae[V]XcD:SDI.=BIBMgZg#OeEg<OP@B#Z^M9?5bFMXUPDWB#
-c/Q.ACL\;b<5E9[RD);fWT7<eegB/0WZ_c)1b&TZG,APRFbGF]-\=TM].@:UUFV
#+>@LRS,ef<Q=)Ef&E_NLe+bKY<FQa=S(8d5<Q+TB1,GGY4a2>5X#fQge^C;<6W;
Bf#FP.9I72?SJ9/JaP@2H<1^BJ8L?XSCIf\UB5WG8=G-:,YKTCIa-<L+ZL#/_G^V
b/86EUA^Yggg5MXY[I=c_1:TWFZa#Q),[e5;gT4LAF@.CZ<dHOL3aGEABWC:=P20
01f/bKX3DW6T(bdPN2O](-A5#VM&Bf[9=91?V\L?U+&@M(N\d<TSc)/4)DJAfS-A
2,UgBT4DW#,0Z])83a27IdOd5IO6XKaF08LCS=XSPb.P>(W9Y?V9:^#=\1^4H57>
W>O5I):VMVBD/>1#Q+]g?+A@EYQXFWcB#N5GO4]]\6A@Qa8YfgH/TE66J(+UCO=1
+STSIR]W;J.HKHG/=W[&XRT?e^4DL.edVTHgaI3:CL0V#-Q)?EeN7IdCSW(9TMc7
V8RG+.<8R;ZaM5/9XR#GGTaLJG78b,8@]PJI,N+LWDFf23H#L4J:UUGJ:Z3;JTP6
?J\g.Lc;[:Z\><fTA6N[NgfW(?#=@2e^c\0@]e++<?>G,0Y,aVM.c]Cb<65YYE/Z
2D?ZH?Vgd2\UQ&EXU]57@/-CJL;>\^>&/e@_P=/YXZ:1;6\RJYK.H;_)>17;U4E[
c:DA\:LK0e-9IU.]-)1CA@2B.ecJ=/a<Q/:e\->&,7B[3T8MSfFc:4N>9<c\Q,e5
U575DX[?77WT5cMeG\CZ6#]:/4ZE2De]<9Z:TNH+eYD9)F7<ZP:Z?-N]M,Z9_g9J
QJ@;?SH3)PaPL>4f4[^g?Bfb&)b;RV^)#.XK0-HL[Ng^]2Q]Wf>K-QDU_ed0]7L3
\YATX^f88._Q#Y6b?UW(5Y]8=^=&2^1N2GF^=S-S?0R-&@_[.A15XPRaYE30TOd-
Jd>;#H7SP>bbGZZS?/fLO>M=ScKMTbXBe7Q.LO5bc_3^gb7TU#I4.D&C[9.9.SBa
Wf8Ag+>4M&C53fZ/FaYQ;Bc,]]\<d=+3&Z1#&WcPf=.?Y)=+^O?\SV<3,/(#,.fS
C;f-56U]M&#eN@5d=ZVM3IE,,4Vf0D\bAPO/IeA9&)a/8[R7X94(?,]@H2^#7K2N
X<U]3>4LVI-/.;_3JI+,dX^/:M,D5SR(c/[Pa[eK_IU1LL(FI)/Z[V/)85Ff6:HO
PME^a191LbId9KQIPI(Q5XXB98XE:;H45][#]5Z<]<M5_G=M>ID)@KfE:)#S?R-9
NR@b8P;MIbPQ^F7--cRFFTQO[U#L>G7dcB3fXL&-Y#05U(_?_RFFJ<=\WB@f(MAQ
XJ27P9d:/dFL+^6.B.1AMD4+ZbQe+PG(+SV6&Xc?8@X/&:5KbU9RIQ]R;5FBg9b<
7S2E+<e;>HB\W(C+#0b-5dOIQ,W#Y-;ID44cW<?(8dYFa5<;Q@,,HeY9=2SH/JS#
O+^@[RF-0,W:_K;f&DR8K]-9K6JCTZ8^GePd_L?/;b6H#V6[d:9LO?VEfOYC4e.W
W(GK.D3&=B^U7TO\,./,fNZN0d7]DZg/b5ANY1^g3b<;C,T@L4)35K:URgR:TVQQ
XLZ,R+XN65KEae?9:+f&V]T9(0&)63bQV+BA4HL+1]2@SKd?261E+cKL<HOHQU_[
L1ba[4@N9?.#I_ZH9+E?MZJ+J,P+9+^@+g0DP):#Zcb2LCc>UR(0_&<&9Z:[O4].
/I:>/Q)4J^.J;F>M@-B,5XYDX6N\#FO5WUL/>:[#IcR=KGO5Q9>[Jb^Kb2ZIWD8&
GJ,@ZbMB4QDcdB#WdI[=]XA52:G5aDR];^Fa9WOgF[408>20>eeS;aB8^9?VX(Vc
TF@HW#U0aNIX?#Z6gPD/8f@JZGeF3M1URAS_NYcE&.a+,G#2.N[C,/Y@R-0>((_-
Y//2Z54#7@BP=TOU5G3F+6dOCL(gFT9OUK)5(G@d#WHBGYSIRYSI#c1,W@?dg=M\
[MWH[PH8/c2:.SL]g3++QJ,6Tca?_/;83?W_[4Af7T8/,&[<U9cML#EbfBUeKXTV
/S/M9ag\@4bY[&+aXUE]GgXe(/.QF7:F6:F-;DUV\=#cY1);a42G->W9VBb\T#PW
#\H1>C1@[0A:7CSa]YUaKG=25]XLa)@O)?6ZUP&Z-2FOFb.VQ9J&5VK\d>W,b<@W
bIS_C8fE;Ec]&D9#M@K7Z1b?AC&S&b;@TD?&a+g4GG]Z=>I,ROFYJ>\&JPGNI[_)
Y^#=G<0_0/+cQ(d/N+Q1QT7]eUGJGZ6D<DCLJ7:^.d9)?e^&^Q?Fe(67U,INU[53
?X]@,#C0bUCg_E5M:cI/Ud86#RB)G25(A6[LdOdJ:?Y9HR>M]5+Qc?^1[:P]5]PD
XE5TP#[^IFbKU<P:bD]cDHP^+Z\5:@2[:Y?.K8+HV9O)9PSe#>6C138KdLA199bA
N3/LaY2P_;eW,#L06)WOD_8&)?UWa7[B]#CRKX9:-I9:6B03I2WS,M>Uc38_E?/=
3cbfO:&&D7WISaV/8J(2_JC6N=5KFBE)><2X&>7+U&GA.P<A>RZ9AALR0SO);Tf7
+ff6@QdbeOW/fWE-A,ebeA):@d[)O^)/9?QGXU/W,LEF,GJ-<gf7M\7LQOD:\S:&
NG(UA)3A/_7&S4&2CL]KPP:9OJdWR5Q0&L^.,HFWADC47^GbR\eIPH6^:?G+G\f_
E1OR^d+d?H<EWH&7[4C[cK(:YBRcW-gOQH]Ya^WR<E]SBTNFd:5e3e:,SWZ5.V>.
Ra@9?>3.-aPO9\]FeM+2b+2d9+GeP]&fHT>>JdVF0A#3CaA.2ND8V3@/fS1B01gI
&2OX:0I7?+X=;4]f46DZa[@2;^.?=bYI?)\=C0NW2R=@\f]2&.<O2);7a,7B_8^]
+;E+aRSXT4fKZ)V^b(#N@;6PO:A6IC(Z-)HWB(7AL:/c<B#bSR_Oe6Z#BMMYP&/e
L6aEg?ZbR>W]G[be79T]EM)X(OMbVH>KA57F2ZbK94adQS)V&F???dR8PB-S6ObG
B6[3,R6cD2\L_RQCeP3=b14]S@V7,S4&D8d[1:MP.WN57B(WCaD\#YQC43ac.,fQ
GW)_Q,Vf9,M,0Te6[c+]L]Se47K,A<_Pg(L;CWV\eHa[=></E[^.XV.(\XdaEY]5
DDeD,VHS90G)A(7:RHX/RM9c]\LS?3VbFcN6BK8;:):Ra&&/c>Zd<#S?JM?:=fIL
O^VYIDCVB>3XS/C4&HZMcYO1+HH??(Q-6e-0Re^]:+;(?B3VGc(6])<HDGSdJ]4B
_I2/]>/g@JJ5#f8L^=O4YTUVQdX&.O;VHa9.E4@adZ,&.QLZ8VdgBYUC1aSDIB6Z
F6\f<C;:BLP?+f)b:bY93R.3>BDNIF8:@X&WKS>WI]41CNQ8WT.?QQ2#>&.&OB-b
E_KJ/7\M)cc9cKM)B.(XBbc//Jdg09A.H.V@QNYT[baHHW/HGfaF/:W,-YgO+891
I7UW12-KMec<NbDb]C]I:d;d6B=:BeB,gAO(SeUE/>.b8,E:62<P1\2N8C_\0+WY
M&SDfRX>@=/,=f92A=;Q2e<77;U-O1[B:3=GL=6&<;^a#3CAZ.3L0FG1\<:/2,a6
RI1#N/]C5)R-CP4ZBLQ6=&&3eY=9BF4FB1aAZ2MaI46;YE?&A^E6;AND=a5:8cM.
3#dN,9:ZRIf0:PNWQNVE&8b3RAHbUD<V[bZ\aW4(F6d+]Nc]e40IK/,&P:[VF4/U
X6[ZJ#6aC#,J8K?@[GHE0#[,K/&RQ]9,S@78=_8VV^Y27>HV]bC,EU-^gLM>A99?
5>SQ/U)L2SZb2YJP,N+=SYZZZff0L5F9]T88J]+[d@B,GLEe4WE..0D9A1E8:93f
.-Bc;88R3;?+X5GETBSbPBg6JCY5;=#DdPRZ0OYR3MgJ^aW5JJUSG/E3a;.G,GNR
+UNGJBgR0Ff@D+B&DFB=ZVe>F4W5M79b]H^(^fHH6WE;W4VUJfF0/5JJdXa>2\+T
-FVTXAb,^7E5C4,BMKI<^85U/F_86QD<E;d@H?7<3[H/I0]/#?,X-8SE27;0=/,2
Y-012g-DPBKC[9KgSZVbN6LIQd\[[B6f@.aIDNZ,A<L+(6-YR1I]]7]>K4WQ+>Uc
KU?K_IK:<d/dfE)^4cP/>09]N&0.:K(;&7VKMSXTeS5H1#eCM,4faf^T29fFW.5;
N-9;Z5/OAF1:N\:ISe30?;3cd\NI3)D.8RUcV/K8U1f_J)agPJ<(KAC@I(I-5J3W
BFEHgQ5YC9O73NTBP(>QGIe#1fXcOb;;.DTDO=cZ=J<.)\-.><O#:85aaJeS8aJ/
.#W@-VFMD[GQcG?&B@0/f>9,\?N43:@aHGf5+I8G?:(6]H>N^S1;2IA>7DbDa:M\
NVF0JeU3/Pb]TcJ@RYMAPG2-7_KAZOOT1GWFKfC?e&e4QZRCM+J>0Ya]8ZAd9Ze.
BddY+g+655W4>ddJH:/F53LVD6Z-JKJ13#_K-MfA]9>/MbZW&F5WSf,L)#]TaHOe
\-VI;9IV.GcZ@2#eOF\g21[2VBRF3\Z1<d175#Da5G;a<cX(H+)e&[,(G]T;TGYe
_@-fKeS8CU\R[Q=S9_.SgE7UCF;?IaX7=Z&.BZRW2C)g72Nc];<B8WQE]]-L7AXc
aH>\Ia&\ANb:7WaXL;T8M?T^TH3T3(G5acQS1/H8Y+UF:.)0,R;O;,3Y#C/S(@PE
:c)>?SdaRV5<GcKOgaPH_7#P)DFLZGY#<BdO^8Pg0bdQ52g(^\M2HcO9WO&IcGSJ
?8gR/bPeS[<8fJ^1Z8Udb1@(;Cc+dg=JSE(ZUdeJ))BY(>@;>]:0-\I;+cYV?@@,
K1ecc+]@_^RLYSVW3SSf[=;GFgAR[OQOYQ.KaWW34Kg?V3E-W18O[DB&?>_DDO\3
2)g]#9cg)7SS2^[-PFRSUTSD3#Y0^QV55VWBX<KT)Qbf]5(O0b2f?I.4KR1.dI0Z
PNP&(2B#D9A;GR0C_89gNafKM4P4?H].Vg@,QQ5CJW9K3.6I]KNagYXdO[U7EUK<
QTQbLB6eZdH];gaf5I=5W?QAW@?PN]-b1+D>eE:/XYW&5#b2FXe32@b1OcRWM6^J
ZRO.&O0[?@>,/WgC(B\?66TYD56O</RSZ8fBf:-^SaBB7dV_,YAJ@]]Q5=ff:<-<
g]FV=;S<aNYE2&\J?c6:2aYQ5;SW8c,^9,WMZPYg?ge)1ARabM&P2DO>G,Z.21/>
ZO5bZSb(BLQVJ^1/JNOUVa@+2@=G3,7[,(+d[R,/c)N0+K14E5)+58=fQ\XQ9WJ:
EUAd:PLdcXJ1H9L(B]F&dKS1=^f+cEgc+UNgUT5\K-d\X-a&2-.LOA2d7FVfbCGd
>d^Z>.MZ+QfC>TbE80]e(WA,H0CQGKAV/fc.4?^X3S1L?G/P>eX<Y(]PGBP1NO3.
<2W88;SVI1S[(6(_c/A=PYVE?BCTM(DQ#CRMS0/#dJ:KSE#b\CV2I7HgeA=QK=+U
Q<\c]56DQ<S,8BTD)0GUaM;0faY]RZB/Y?6bI,:=[bM:Jb1&e@gMVM1Fe:c+GUXG
-EJ)?)U3UbPEQc042dTZCEW\H3Y1.R@\,O&D?WY;_<39@)2\K<b-B4>IK:6>gWQE
\/D/bXRYI@<W7RdPHC_^?(e[H[I3L:@:16>-K(ZE^<aFc>Y(JgU+2[ZEHD3(.,Nc
c-E+J:Q9Z1N@L-L]B0BY&aC\>-?YFUJ_b+N;PI@\WG+Q76a#D&?0,e6gN+\Tg1e-
=KY37+CaV84>R+&(3/,SX9:&9Y#<O_O-Z;B0I[\\\;-&A+U(2-KS)>C^8>#C4\K<
d\LJ(7]S.\W[Rd]OTbNNc4;Rc=13]=_LH_EZd&S#I)a>,T.16b<c2CS\417@8E@T
GBR4gG5^KM>YQ.?0b@.&EFHF:BQ8Q+)caeR//WODU8X<V>a=X9HX3ES=01#G.61D
bW77]=ZK]I0PJBO,F=O\)K64\;JTW,a:&Z[BJb,LXXD,OJ&:8?N.?81;S+>T+#D7
>KX3Je95OK76#,.HBH5I9&K(D\-0a\]5@DWWPa@@_X>=H(:f;YHeYDV0e<&Qc,DD
FVaGP2UGO86Z6J->\=<_D#(,&73O?3+0YW&O-XT41aV8e5:T+6DJ\,ECQ3KfgFAa
K93-7aC5SR\:?Sc5MY80cP3E5:aOF&5BbbNeU<YC3c?S/KQI4VHHQJDBZe_4cWY7
XW[&+e-5e[>1d#JQ8b98=[3<RH2=K?&5C/HJ&YSHW^efED#3S7T66,^D+X]7,dXI
)LbF\QI4^SRa6=SG0#<YO,[AE7Y3;)<SNM3e#T1;[bad8OgagFJDZX/Wce(WL/\^
B6TC>a]G5/3X&N/aRDe6K[b:WJ\.M;\_?#4B2SHLGB1.-RT:]?PEVMDAAW7b[17]
^Qc[#b[C5EY?4<]D)^-PU#NA+c)_>Fa=XU-dSYX3/K^-H-;CO:</b3<)AW0GZgCK
gaPHV605CE5#])HR]IcP?fTLZY4f(1DEfC#f4GZe+T@cWf4Ca[>/V?YX7&Re[_(#
P43cFR(NYSHBS>dKf^B>RY\?X@>:Kb0H\_+P9JP9UK5W;[FBaa8.K.[-6F38cISd
YXfXec\89Od,-)bGY<e\2g8.4,2WG.LOcN6P.B_VOILSKNLf=RJc76R/B#:-V)U#
7U)eH1JbgH?)e\IP0HTSU\N\6Le_aU:)/Gff)cJX8_49Z<F:7PI_C(RUS6aY3X@]
_1<^7UDOJGR>>W8\R4CDH>#C3-=@=IDW-GG:O-=NP^@5gO\;00G&cgQ,+[O1=R>2
X8?1=B&+fadN73KHeaS.Y?Bf8aX^G?/)K#/\1XUK)86^Fa;;SWD;S+&34I>B1@ZH
?,-=PG,4RUG8/16W@9-LUVQQSN@_8(ERG+][6Q7A@>4UX?W3RLK2#@c,2b):2]gH
&DHG@5,C;IY2OQ^Q^&&Bd05KFg4Y\;2XB?[+/D>^bdU91b:FLQb(=OFHFa+Va2I6
2QQ:^f/WcW1<-E,&D5,SPX=H=_0gK[,LLG>\D(1-OeUB=cGB:RZbWST\(DQfN4VZ
JG#+_;bQP?):GMPd_R>E.-:_@SV?c8(X8-&/DV,)&.]=4@)fTRg&4:Mb6gGGACc4
LGD/V^F?Q)DGb;;1ZSQf4cU-=L(_\2S>XS_0/-DDE=\Od=+G<ZS\/g/7OYdI#_4/
S2Y+O]5JK]<-_AHX/>aQeM3e2a/]LRO+S5>FR_RV]Q^IMA0,.gdF(/9gK&ULa?T_
PC49P<3^>(8:)]_<G/R-:RGK0Z,=-I5[Ce=;7]AETaNB3>FPc:3H_3@C.U+=SY=D
6(@b_#_W(?5-d1&H[2URED8IfZIa,#8]fFXD])T?ePZg0_WA&eGA413KcC3ZF=^,
,#e,E4WFG]#QSPA<2?KgTMDAZC7M;TJ@O^3d(JcH[\&aZd9XZMaX+V@^^6cNFeJW
cdIaGJ]:JVX4J,8PN#4dPOI^3NWAcc5Jcab^KP[eJ66<;@&gad+WWCP&57&E:GPH
TZJa=d4XNJY^8cJVTUb@)C@2(GVSB[5e)L^agc\c(5KY^),bLP32U\2&2/R:ANO+
MBBZ;44._^fKIf2VMXZ27a0(#96?I+3cWR)Kf6cBaB<&IAcfc?V6R->1YRY,+b4]
@?[+cE@6,XHT^Y(-4P]>I_.OEAd8;R2_>A]IQ1RIH-I@;a)(/0c=MW0?:]#30_]b
8</3dF^Zbd8[]SEQg:Q=;M_OE)>LHF4?.8[Z#FCR_DD=T@4=b_:5J,35JL;?Z1#@
7UZ;K\R?I?;AQ9;+?f7b;_I.#)D6Hg><QV9Z5P>ZOL3D16#6Xf3G#B4AbFUD2He>
RAG36E>RgR_/<1ZYD[GN_JDR?7e[d;V)_@-K]Uab-04-Z/GIPK(OcS^LA(RPGW78
CUHDg:8@=LZNC251:e_2566T5g_&I#-D@N[VbNL>8(NWOI]=XXH002[O6E)PLfB(
S4U4]M+C#Y[f_g<7&[@@7^6<B0B8ACfQ99a_#bA.UD<V2:;gAN;/G/B\T2eNDGA#
_UQV<2Zbed:Rd.._J;V]c9EWd8I6^+XV&W;QIQQ:[94CFW-@I36PHD.(XK5F2T4M
deM-DX^?A0800J.46/35_]T08F+@7f/ZNY1Y,I_5:-5R3LE^]=\_=EaC[.KXc<L3
M)Vb(]Vf\OKA1IMU.P8B\Ae[[G00J)/2c[VGBbdE&)FR]6fgQ5UMD_ES#U:^E_.b
O]Z@Q5V49KgEHa1bBV[_-UcJ.^7I99aZJ_H[\WJ0ecgf<Q\GW8ODW^Q\&YS?g@3A
H8^##WB3<M8E[K&UYMPNR?5&,2\>+d:J1]Kf72X[dTJ;#TSLB2/=Y(_fKAJD?6H_
U7?U+?LDX^_I<YEA\Z7P7BL0IbS@/cP@Y-K^8>=HU9D84TL5XBFe:ce.IL@2[EZd
c5/GECGL=<f7J_c0[QE.>92X^BFbCAN_PNL32DSc,]E4WK9NdYd4aVY-RC#0IHg&
Dd8>F@PHIZL@ND5cGH3Ve<N?.<Fc2=973[01()MPTP.>-ab.6^:V:VDQ2;KU;de/
d7&9\)_d:g3Xg[[QETI3\1IFYc=KN/RB&0)M,-T^EV>]))D.1/>XHEC9Pb^94?).
BgD04<N_f&_>=MB&?,]NQ?,./.+V/M<aPQ:f>ZS/aM[a#]?DDSY-:WK_8T[XKcRY
a<WQ^WJEMH<a\3XX&VXMMU3<,]O_R#;<3)N@2?FZM-NeV+LYDG]D+^>XHO]b2Q3[
E=3UR>dba3ONK]a8H-\ZJIdbOH.T@?(0#IYdY<=0;-M=Q/CB;_V9<]/N:(>F\J>:
);@3MB(].;a4f#Q]cCIP.PT1J:-,D+V.8c]J?0b-#)NWS,\),R)01H(_d.8dV0=]
,]\_Jg1McfTbT=EUe7)\_1ITYM:7b=DZ(R@+T)MF;+#e&3b&E,agf_e.\#M,cEQ\
A.I]8V]b[LSJde2\-N/5@_H(gZ\8O?OY<GUgg^+WVSK7IgY6:<-]RQH&)B<C]I?G
Q8?,B2WW,6]>g3?NE,b2W.3gNBgbFa/\(-KEZ5K&VM?9;-<-FB0[S:b9I2AUQLKI
,DaDGdT2c9?eJRE?agXF)J6-CK=2R,U7ZIeZ+AG>K_\,abcb\.:+A>DX^F<:^F:Z
@a6JG\WU=R/5.-\GZCE-:HW3a.gAGf[Cf\(8A;?#),;2_>]@g([+bC2;V[g@HCLb
_,1GZ)Hbg[6:S5E&TcJ]^Peg@D@I-.#SL/T,>,0:-GF,c?_FZe4+^?&7@6;e&9/.
cHaf?T)=?cOU&1LC7:)7bgQBK1X=9F?V<H?e06eV_gb,V69G)SA#_?&IF@,bMT5K
2Q#OEW(?H,GRL.QL@FAW5Y__\&_:Uc(=gdKaRQY0/a&/&Y;M2,6C:D_.NU&=@45J
TGO(egL&1dTL8fO6VM-Z@,WY_YHPg?(:e=O&?P7GNGf/K?]AK;6,W<]+S5bNLHM:
b<g#0G1L<IV@V2aG@03O@41JRDA4:6C#T-R(+C]fCAJ5D/G&<,]Ug2EWLJD/-X0V
B.gOD17bGG02([Ka1^FSFAbRR+[UIgVL_)Z(U@RWeH.^>EWV+]-W9-ZcH2f1\<8F
TGgW2XG77:6/[A0_8^&-=0F]&,(-f_[=2TN#DTdIODXCY4FV7#d;(QNPgK2D7;2J
a^;+fC+VA@TKA5c^KN_\,YGf\JFb98V@_\S8a7#P(T(D-U^28P/gg51)31>IDD\Q
GWQ<3;Q21+D89I2@5<5G.R69>7Vg7c/]:#Q>@R@<ePc2TP0GAeV(_KWU]:/+^e_[
>]<#O0.:,X]9N:1,T=[aH5;:E_[A?=5/JI([BA;DQ<^P\geAecdH.@NTZega+=NK
a9ZG@g1RKgb;7R;2b>1O0:ccUSDVe5D429bAOSEcOdFVY1&1]eIb8>:-D\OHVSf5
S8LR[,K6+58;UE4#M05EY1B8^IB;+?D<,.>(UAJ)FDC-Z&&-aA6,=>)8)[E6)[(3
QZDGXI9E@+V&B?FGDc3JL^4g6J9>XX&eHTZ_c8?JPG2b-6_)7G2+WdYKFO[\/GdC
3?<<--0-(\Q6)MK</J5L:^_#M4U;D]E)YS5IUJ3#Z=GUBADZE[UU0NX#d(3\Ld/4
QSe^/?LGF:=+14_E.D+5MQTF;ac70_D5GS3IT09([6:7CL;D=8ZN/_Mb1?WD+[J6
7^O0aNVgX@b]:b<91LD)>H??,H(T_8]R9CO8Cca9d07L\&[<5P_;a?SW@-2,N4HM
=B_#)c_XbFDEQ5:RPBe7CDS@HRD;QY6gQ>++:]aCN&,1V(c_G+6+O[<L;C&4W?\?
]Y2,0e^0;XcWLQSV[WOAXZ9:74_S\D0Zb7U#cHdU\1J/;f@0e]abT1W=\I.;6J]<
a6&[A;/?0\J@-Q5H6-A5Y6aga=GR(5T9DUB8??YdXO#M.Z,c9D#>C:fJedHB9LJU
1WR03RKc^/(;#RTf)4_K;89W#8PG^^:0EF8c0ca./Ed6JT;IU]5>,U<2&?0__>\9
bF-/]=f\IMQ/V,[P4HD48+I=H)>J^[:IdT(Y1-L:41:VP?P3E^X9P7V/:A23PP#e
=>d+CA<8?&3+g(9XeD+6??^PVM/(@CcF@IN\&]A8-3QZF4S[6@/4M(g):KMZ]DQ2
F?KHMQ>I5Z0EYA>C?_U5VZ+]=,M<L@Xf[=57[4dg9W5TYW]B^T&<(<O&a^9IBJSf
bC,NICR>5UCY9UD?XZI8^DLNbN]5U]T2[a9eG3^\RD(8SBXecS(>OFL[-MJY\UVT
THMLV/VGI<LM@e::XUZ#d;Y+W@;Z6fG9CJ_S/+\MNZZ/+)#4:O^7DG8DK]<@[#BU
X9F;QA@W1YGHd+LK2#443(7T+Vg8<IZ23YcWFP5\+g96YZ?))>.40IK4M5)TXf&f
+27CZ8=;?DAE8IH&aXP6X9P]B9)BYU>=31_gA9,YY9Q/BR/[<=C6:F-<K5>g=.dX
ZYb_Jg=C+Lc-V7.86+)KAG2MN0C>,b?D2D39AZK8O,H?ZfXe^1&NFa+I)\>XE#]#
CSIc4cEFWLM5.T3&/BNH_eNF0-Z\d57UQ<2+-JE-]GP8#Sf<)\XS##J8aM,[_R_I
fIWg&AO.(79d5&+e@(&XXcfLd6#_J9a7OQB1(0-;W_B@9eG)ZU>[>/FdA]/M(Q)Z
aS96(Qc][C\?ggE7KA(PO)d+N46@eH-RG8.?=-&9TBKbES^=9R5:V^Z)9AQ4F(Ob
c0]TSGSM#(e]RP]@EYN][T3(?7@DD5eY<?a2g3ce2]\3,4+.<fC.,-U/)&cWH.J8
HOFE9Wg?NM9c&D6LAKbcTLa1A,LE365F?PKcSSC#Vb1-TTF?c?g1e+&gUKS5B\M\
R[>#bf<J:BRA7@D?>Wc7K,b4-fWE1X\P+NQ^f,5\8TV13;fQ<Hd[aT0&bReZ=QeO
?8,DRRd#>DGT]30/ac&B;XRR_SS_I58=[1,?>8.J&7ZDdLG)>&IOf[I44\]A?5TY
)YC-,,aF:4T+OV@6W;F]Q5b9@AJ.Z#@O.G?TWB]TDHXTW.ZB]HK6\Kf5+ffYHdgK
^MNFHRF1I<AK:Yb_KU_W_S@aY?F)cAL[@LF-^)6VbF[1D.]]D<5HQ#[P(8RVJ:S6
@](G[a@B-U&P#\GQ?(b<Ief1AR@L0,dC5PAbfB@JeN;,T5NF/)Hg?:V5:M?Na8Y1
C2;,]34K#<I1->B4SC2?(#b2.>@SR=:KN^:,.=8W_RfO(AgFe4<P3G4\6HgB-9E#
<:+6AXeKUAPFS7N-->3T)R2E;]=e.7Y9\KNT@NR]IVC[P<JG3KIg.THbab(UB,PE
>(Ye3Zb<3LCf.EXODN02=GV(YJA>g]&6IJVUG5?Pg=Uc\a\;2;JX8.#2.<fO@3U3
JC,Y5CeHPJJI>B8c&)6KO23<^9dL)AAJ<M))2>XNIX9fM6,df23GH9H9DHb7<SIG
6<TGK(\;A[5BAM0c@R3_WSJX_<.H:A2=A0I5dbaZ/#bCH7&?6C5eJZI:K@?_;]X)
aN<X^\V[:4ABF+/X??^KN,)P.8SI#:/G/TV6b:gNM)eWL9N7b_4Z=L<]_<;RaH<4
UAfQcS.Z(\A5-Xg>(2>K7M]d2CIPLNe/\0&UE\9d(FQ0g2A6:H7P5EH2dG23BdbV
dbOX;\DEI[PXTWBX,d.]?5.DYTPDM;_4??)ZCf,&aYQC\-+X<Y45\R?D))IW=eMJ
Idcd;N5g6FT=&bJaZ3BE(17]5-@C&)@#@M84B3[8NA@-[X-SXR(#-2f3EgYP9/aR
>A#YS#(&Y7>ONfFD4@fN2OXdCT@G0U^X=\7+(5@DT>6RQeOT7XBB<6<#BTS.A5HS
RHWGa9[cSPY\8<+XM5X4JC=,/Q,21QT1c+eF^=e:=_)J^>6YFO0(O7L8(1FR:>dR
SVU]W2bdL;e4eQO,J0.AV4J&=IL?3d;R,6[#3/:=P7NRD-e83;ZW;2R[))ZPeagS
U9)a+KD\JZbLC?df::^HDL<\FEfN4F5Da5--:fH\\Q_R?A=]\Ka5E;EMF/)bU8gP
L:195.QSEbBXD-SXFc/)^Zc1]9gJ#D_HA=70I90T<=T5UBA57BGX27Ca;KWSFU]c
;K8CDNPF[R:R4[(##H/ZFFY<.c2@YV(N>W]De:VLP74W?eaQ72>)+,]QW@X>KO5(
LEF<CG<T0OUB#+U#3Q,#O,<[8A\A(CG&CPE@Y&8GQ]O?Ke9e=FJN_DXJ1J+MXAH/
<b,43aJe_X.D]eafIbCMD@?8=7R:eG@_QI5??eQaPeDc7[]c5-ZP##gIS<a2&<>B
cJQNVHKa+C]GYMH0O7W^eB-YX(?>QRcO^PX>OHeC;2P.K>\IEfGUY/3fOReeCcLe
7;I.K]T_./A./3JH-/cV&1<@bO;Fe3D,HLOg5Z)5V-EGL4)^=#IBI0C6,Uc?CKG\
Kgb\&IH[:@IO]T?fZ@88N6+-TR,2F\?]YD)aJ1X9d0^.B,6/XE0BAF9gIV0PO&.<
;/834DPOT3I(.TG&HVUf6;Y==(5\IU=cBg8/Z^QGb/cM^Y.]U(SIJ=Nd>]&-6c2f
::3.-AQW9>72a,V)V_3T3e(D0BQb.6@((-EIMU:2Ue/@.J6.EGRfLTgJWbNKX8:8
O5(RKd@BQ:d5Qd245Ee2I^08cLJM>2)_^DZ#61,KQQN^]PEcN4D^O[:H;dS#@MZH
_64<8IBZfG=1a8BT.7I6f/]L-WE-R.VW:?XU1<M@L_M/A;_M,3cLI.U=;PHddbPT
.3Ue_(\)+VZ\Eaaa[R&5ISb/Y)3UC.(V(9V.MQV8=dTTg4)Ee3KBU?U/U)^+KcK(
RJfIG&MLLF,\]/2ZS7YCM>G49dX91,\LY48-c38N2UM4e4XGcgS,A[dPaK-HK:71
9NLEd1DXaTgJDAc<CI(5=#4D^aJ6UJC8>R^4d@TeMOS\L:,bMa__CSWQV.=.KH+3
>:\[1K<9\8U^cM.7#b82<?4cB6EYYD>O8C)AVOWV[&eF\f2+<U@,Wd[VY6f_7:K[
UNR(eFd^\a/NA9QZR]^[=B-Q[1\ZG><8PW^ZF^)^aU^aLN.-\,LMeM642-HPbX/I
QE\AZUC(4^8LLXcUS]OCCBP4_=,T9bd[R#K2:D8eYb&a@@=;TRaTJCZ@1#N3K?1;
S9CWf=K-dfZW14G.OZ)T\)f,)L\aO_#B7W6C+Tbg)/E+bH-BRS+NBZ^e7dSK-?8S
:2V1?Ia=6>ZgTY1U=ZDW.2c-WXS#d]M(e4?_YIJf.S:6-#>W>2J;,8X/X7U==C)c
P8H7WG[[VFUY<#DF;e)f@/&YFS>g)\+f)U[?8B(41#(3#-];?>;\?I2W0W>+/<TK
,B5MBAY@2])L2K_TG>fRN9F:5SV/Q+4e9VgY#Z55<07#>AaPaSM_KO(gb7.1CaY@
a^FVePOMYc1g8/\T30AHI9MHf1e_XYSTBGTaFVP?=?W/F&/U9M4g&8T@2^11Pf:E
TL:)PdF4d-,<DQAH>/:K,9/C07G6#VEZ126e3JOe-RSVbg5P)a++e0>BBfN_N^ZT
EdVLeg?Q>9D-DQK1/ZXSe@-1eg/8@>F],JSR0O_#L+Z+DO.F98+\f:13F(UZY),-
)LVdHNIO)a:LTB#;SgNG>Zc((?;3b1H7ZW7R+1QRC7MG>]#IQ+cg@D^6dgEW)D?V
_;,fU\?,V&.&(Ag3<R>VZ@V2SIN;^gV]E./]>RRGQJ,-\3T[-X2B;-,A0L1Y=,T7
1(f&RRA=HcfV&.HAM]G1b6JTLSM&cWb97_MZKYd[6^=F5fISE:E]CO+0gbgTW>Y_
YQ9DQRAK]gQYgR9WQ][H#0P2Mc=8g)2?PSQ\05+,-d4F<1[a-39W7&2_[Y@aTE^Y
WED1F9L]EYf:HUZ4E.0K82^SW9V\I_<8411<RE>8JT]8Ze,A+W0?e9,>MCY??OY9
MC#(c1MD[ZM#-TLf_S(_6B[;..(_9_ER=[/g>a=;QWEEa;)=f-GZKe8W_45:U@K2
9];:e1QV=:[M9?&?QR\+Ld5Q=#1Jg(bTG;>S=T>L8:04eYARK&:^&UG.-\@6U&ag
cQeAXX;7aX;Ra?dU^O0G_.E.dcbW]GD\G@[VO.8YMN9;\Pf5fYBYWSbB[;^DZ[,M
9X#_aRaVE)Wce;@5(@JR=MIcP(L4ScL;>-Hg-^d]<Z]?VB;);f@J[a_+23eYE90g
Y(RGPXT8CbXHV&K4YAVVQ.Qe23]B0/YP=H\Z3aEFM+TUI_,b&a3G9:R<Na-V6+GW
TJ[?c@K],e_2JQV63^BR+RUQN5F)I(ZWS4<Qa7g&fZZbU)QS4&6Fac9EC)7^::#>
P\4UAZ=(f7g.F?B;[/[LAU.NDK?F:><1S_:#KZa.SUEZeYacY#P\E16B.gB+7:R<
^WAd_E.B^F_XId5HJ<D,<c84T0&<JZVe[MT5<4&>7)=G[^J5,R<C&8AUDJ#EGJKX
\T3;C_<X)bHP5P#?IB?BacCF#,N-RgR\:f@6TQ&NUe0P&15(OHDA:cW4OeA^3(dP
De72EBDV6T6XFX-_M>O5c_N\<MUeH-=L&b5bC@EWZ#2^XEfM#]@6EYX0(,U6-50b
D2TT\_>4N=EZRQeMTPJ4U=Cd=>>_S#U\<@(9U/>]/eS?b7Bbg4LM+Bg2g)X)V0gD
JJI&LYWLO;:=aE]]/:SL6&+Hd)2.3)OG:5c\(P_F51G<)GYW7(/Mg4/W5#&1-&4W
JY9gJEcf;O.a<)\2.\&\<NJQ&GX3;0dc&[3,gbQd=cL/8eT9b3+&6gSI,4G^7DU,
YQWgc,TI//1IW5HagH^PDQ_.<LU8cbN6JV\CX29.Z-;8BJLe#?>Be>#fX-::-cZ1
AB^Z#9[)?]MR<D/H5\JYgH[I&5Oe.[;A#U1<63SW;?^8Q/<LcCPCDSCX^A:J)MG-
;J6T)9S9,M-\]/G9ODY5LYGVLRN;Lc?c.99I[21+X)PB#1FOAHBeZQV5+a;+g<)D
\X4Pe4\OJBI<]2C2356,d5?NF1S/RW]CDU269@PQI<.KF=c?C0M:3RFJ@F_fAKF,
9LRL?2a\&?[.&AEDdgZ>g3JQ.8#d]4gF(]baOR,AR[+)=,#.CXYe1bJ3,U+eEFK-
\1\SKS49GGR<c+[[Mf5TA0Y0]\>O)>_5eY.^EFX4U8e?LSNS=c#LXMQ),^A70@H4
1K&>,\.3F4-LB]Q5IUZ#dCL9(9#g&3:GKOTORaOd=Y5g;9(F;NP\PcbR<0@2/AK0
DQ2:B8AE9COBS7<9FZ60:8G?5>[.)WDZ0J\#8eAb),L[F+.=2;Jg;C>&HY7cTEI6
Q0/5dAGLf]WTe<c-.55aCgB0MBPSZHZLa^bTd27Ja)GcTY-LN5[BM0=gYaFR537;
SF90adI]HgQDJ&DYgf-=1d?V(Qg@^T[ZcCXF6LN]MeX@O?;J>Pc9@92F8]NcgON=
D.Cg&H/#I.T)-(agV,E2#Hd\;^)f#6fgc#=;O+(^G+.7Uc<7f<[[UZgJB_EZO=WN
RWdFH<<EM[bY+.<bNZ76UI.NIaAgcd,L1f<75XPNNb:Z7J]C<X+##D-1Z52g6JMT
=@-&PbSSCLD5EAgWDQA2@c-WNVMUWZ[[2@H02?K8?cZ&;(AWM991fIPEb4f,b<De
<^dIY9eQ77E^96eQ5L&U,_\-><dUK=DUJB/-HR.bXS31OZ<>SGJ;GEG7=FSKgZb_
XQJC#>XE]cfH]C.[^fA#bcbf>+ZJIB3;E0O(<^Ab//d/c,Pg5C)#^IE33eB6N^,F
03OX-EDH^_]Tf^O56ZA1,>--a::^JK:\Y/<H9VIK[YADH.,OeQ##]g6P?>U5U8.H
gaHgMcKTV3.</I0/L]O])F#agEU]1JN@RCW0GKbKYS3\>SD8]>M[e2+9#[B))6Q>
ePb,ZGfK>MW0^/A[#<bgW/X=;4&>34[V3EV^J?PN\<.9V8B9X-_<@0Pc5W?McD44
c@X,&U,Jf\^9M0,M>g@gMZ=D3^:VZ\7M-O2b(X8;I@NSO+OQL9QI,]V0UA;@A&.^
dJLgH+?J7QF/>=;;-X,=F1G:H]OJ5MZ\E4?#:ZaUM/e;49e:Z\7^D\-[d:T;ae3c
/0-dD;6ME3HL)9Y95<K1Y.WG8(39[[BUE@,CP#ecHF?eaA/LK[.:88/AabS?OA==
eQCfgKNeA@f+\KV225BINL:ZWJKMH__AD+f&?ee,WJ4F3_Z1[C^eA+CLB.PT-3JS
TCA[G@:S+IGR0fMYW9^;/PCYRbSY2HBF/d+#S1[[RGC=fG>e8ZB..Cd1fE3#IBe5
+?HG&)W0H?ZG(@S?Qfe8=.?O<INXFaCH=[(>WL__VGbA8\HFR0PAcVH)8X?WbK;.
E:(4NFET^L;;LIf1-L.S:#)\d\0I=+S)[W.Cb/FDX7c.8_XP9+CAH44A#<PCFDSW
MHIX)LBJ]]&\bJ,cZ;(5,2S/E>--.FR/-M\6E8HA/,.2]UAH\-3X&G]UPGS8F^.b
?8].(b5VB;<RTK_NGSIK[?2G>ATND.G.>[S(0HM8R?Y<g,Sf<dN&UXfO:6ZQP5f#
.J\;&Z#ZMEWb\U;N8f5(EFT;F-,&,AM0P3b=>B+dCMe4gP3-_ZdG-L<gO,Y;N2YJ
#JT1KK=7Wd9LZIFA#AZ=g_Le+;Y8#.R@8bAaY^9(_.CR,_7)R8NW8PY93L5B>NCM
WV:9fZXF./5GNRWO:KLf_bT,@<e4U_R?MP?g4N(Mc,1PIWM6A\^d.Fd\5XHbcKUb
8M&N79eYS0ZMPLg??V38=fPdC^SbX=@TVOSS.]W(IA?L,,9T@PeX[A5D6A1C,PD?
3D_I8&J..F=F@0S)aGBRUC<D076Y1&:&.RfE8MA?ANS>4CRC9M4BI:MAb]NNG_H#
bCGMBV5.:B?6LA.a1GYG47A3U3VS/_LWAQgT:M08M@MRXKVY3ZYNJ:&]+\(R[Q24
.\c<,8UYH@5Y8.CHFT=gIQY6/GINLBe\1aaGUW1Y/7Z<Q65,Eab5)@N5UdRG59=)
(:#\dW#c7:(DfOD=(@<V5PNQU_SP:eZ7LEG0DI7=OL-W:D2]E^OMKbd+XR_FQMB0
-\a+Q)N(bY+\fYI=8-HHQ=BJdZ#@IQaZX3\:2<(@<AB49O9deZ@8@H[7^]QA^UBM
EAFb.=S?Q[V/AN,VM:BH8e^SEPS)0ZdfLcAgZ#&g]042[F5_\cF>4NV-VgNPJC2S
<\S=XU-G)&OdY?<GSI8JcK>.^JeU@ZH[CFYD+Q9#@)TTD4RR.b:_<3+LI8_)Y],[
MGaV-1Q&B^F@K0Vf.fVA,a6XfLTRQ6Pb6MFTR7(f]d\#ALQL@-KeAYA8Mb)cLaP<
Q>aO9^A&LfZ@a-LdW4X0NI=7dB]??UPNGC4&QS)dMSN0<>?g8(N-DAEfbg(/^?WL
JQDQ:&^1;dMeN^]T?.OfF@N/<W@TAXIXe=23U@I4E7,A4P>4ALZR&gWREQH=\dF?
(f+5gHIR0-bK(c\>7Q[LO&BEXNTb]a4dE=YOaUDNL-dVaN6#O.K?95SGE<#WO\NH
@7-?)JXX?MZ=?3_\J\/CK(fa0VP3&GOE]\):CPR]BTeBQ&QS6J5aE3Sb&),-K&bN
T0AOE:1Ne-KaOf8,,N:0CJN(JbQKS)-X+,CBP,QXQcH2+eU#Z8D-eDBb7bb.c_J)
gd]X:?LD:_<aHD:>(JFKQF#E.JfQ0IYF]-=Q/=ME9+FC?N3/#MV3HF<#&FV>WYBW
U:/P4&G?G=-9SBN\3EHK[XCVMgOV./dKcce@_S-Q2O1=P-L=A,UG0NSDFgE>cBYY
R18P0O3TB5>B#@5#CRNcR\+UEWbQb8XL8+#R,-9G-:]&e,Lf#C,J=R84FO3KYb)H
&OGE+)g:Ua\#Y-fURB40.8f0HCI0/+2Tg/(dZ^,;db?KBT@2M;M03-6W5:bg2+39
c8X=68@f0g[S2c;^XYbbaG03:agGIe@e@ISD)R5\LU\;;-XCN)3d3RPNTN3O#AWH
[c;D&)\Q>cGC+@P=NWXLZM2&OA#+=g>1&MRX&b]N]L+1E>[.Y/UfA;V=1)R7_;g#
=87Td)/2dIB(Dg;[39d,.@I].J#dbBRS>9TS74A,4a/ATAH^]LM5IE^Ha-I8Q#M?
MGcf2F+CJ>A^FGRZ4cCf9[Q-UER4(A&=@JBXSHWMdB>Z1?F16gC23YaGS[)C>4ZZ
cXTRJd1cG-S/O.MI=P#@7=B8?)?.,RL)<;P/O5@LCU@>EQId1e1N3g06DWP/O^.U
84POIg+DU,-PP-1B>:Y^24#V/=CZQ:DaSF6I//ZZFPTRb9ZJ_PdbeaQ16OPEZ)6R
N#=c)K]DNbOTN.bY1UA>OQ?X6aHO2L[=ECc7OX,,I#eBX62:/RC0Z@-,OK>#(7ME
N]^R4WQ_U+VI[RCQ&)Y2W;RX17_UU[E9?cK<JdZ:bZ+WFgb\XV)fYL\8KS7c+CGa
>c:GE/bR5KcQ1<99VU2ZC,[G[F<?e4#S&Z#Q>9PMS^BPG(5@3D0E52=BNeXBRcUK
_&b86ALS743e6+FG-C<#IO[[9@ST?3@\:V46^MWX(:#M+WZf,)H1Bg_a]OMBA7Y+
/JO-^#IdgSf9KJ^<5P812OPVV@W?8.IP]@6.gSO,]V^LWHW>2WSO>da?c#EFCaZ;
[FS[KW^5b>>(X&=^BR_e&.4\J[(/X+)4+LJY-[d=XE(f2b6L.[bO2)eT5KV@HD7<
aPJ[1WO(K&4VQ>UaV))D?A>34L@cZJRWP8=?H\8)VM11C@HN&U6=GfA.#+X&4(c&
MIf>.(bUAX7GfNC9P^OX6LeF9/gCNIQYd[O=,-/+aPF[HFUgWgg7(;dbLY-Bd2@>
\<B[PG+A]4MKR3K_XT:W=2AB3C?)Z\KBIf>2GW;[0N=7R(Y[-0AL\KYKP(2dM,KJ
.A&ZZVBYG2CD3<TO7PCMUX\1.)4A=>O&.1QbA:;BBL8@9]3.Ae)/:a_3Q9>:FKQ.
TfW-]:Zg[K(NH94F;CD=D>9&C.ecJ;=SOH;:U7V<3H3T>)WK\e]-LANBf>c<d0]-
3>AYCIe\aD.SB0F5\UN2FN.&=d5.=1-;8@(;[7+5]=3:C(_:@6[e4^-UYKVC/I4D
I;dK.#()P[X],(9UfMX3,)1&e0PPFCL>(^>M#X7_@Y_RGJ5W:bUW=.B[8CKOL-\.
72F4Y1.#.R7RV0)<_geOLDPa0NVOXD#MOcV6=YX@.I2,)b6L[J1YV,?G/(;RI@]7
SW&Gf8X1:>6-Cb1TXVLOJH\4C5C>cQY+-M(DUSX_JMEEZ2I3MZ2GbW-82M^#;b>R
H&A\F-T/?_[Bg=dS=H@,2c#V1HCNBbP5)>B5SIg[PdG>TM75(4M6\gJ.cega#S,e
3;@Df^P&gZLgMP<19DD:8NCOcGQZN\PdP?<+bYFN.J3Y[\#U7&685@Q/^\LM)Ga\
;F#a?4WcIG5KV?92[\1D),,cZ5&7eLA5?HZ>FQ.^Q+HHB2NOPY<@EYdL?FUa4d3/
X)P8eeSaCBCKST./,8_Mc:d6PAP4/[31=48XM9RS<,b#T:^U1ANZ0E=_G/&6K2MR
_/>(AAX#3D[SOV9c1d]cV2<W9D1?/VH&dTBSfIg6.^f6=eAIZ+O,Z+@-UD_YM3=#
OB+gJZeb\M@Xaf.JbPT8[^dZXO64RZ(9:LX_U3-.9BIKb>gZICJ;#2XfAcHX4,UR
:@YVA;2N#LBNG6&H18LIS57gDN<]=4>PL+\XdI9f&4:TIW8SQIZ^:4CT(U/CCOQM
XQS1c+f&PO?_2BM>3a^7(W\,H0]^GKW:eSAQ?.SO.+]cC(>H)EZLHY>-\aJ?cXcY
.;fgR#8[fL55LF8J0X/FAIYTFE19b]04/a.^I/6=FK1HV&EQdZ-.X^7cWB4PO780
V+(a?&G)SI@-]=]SO/SPcS_DE[+?[Y[g#:_DJTEgV+1O1(W]@I7.1\/WeD\V]U0O
aB_GR)M7>-BR\N^Q_]VB.<Xc^,S1]FE<=MXD=&K0Rc(L3ERNPCbXS::4W\1BeX\(
W:D.-bd5c4e/aK=@-9S_IPV=>71CIA(VL-R\@S1a\@PM5HOA&Jd8DMZ#<4C+1.9-
,N6WT7S,9+<IR(N+-H=H2:;L3B936;&VPJfDe5@(409:8eHCN<GG7cK>D)<DX:JV
]\E-^N2EA;HRL5PI<bFfXaQaI/]=:dMEIYePH0+>RK@X=P<A1+4Gd_4S[1EHOKVg
WAc>(eKT-C1g&N)^5cS@^gW7\F56PRENeUe,#0RM-W/B._^20VfMgYD5KbSXQGIS
Y1]/QZ5X_0bW;)M8F#1EQP6;+#KP+<:^H>A;+7eJX_(J3LS5#NRE[1,^3@.EV2DS
Mc?fTF/=K49H9P9>eJ)5fJ,3O1Zb#AQE;^#.-WDV\(1#UT]gV]_&/=RH/F9?L7a-
D[KaZL&6b?J3gZZ55#fQf\_7&6P5aF@-YB)3I--@Rf&TeA9-.;):YC0N>D)+<6gJ
^Q1QRU=T^0=eV)f6KGaD,MS&?55;VAOS=4a5.Q+cCa]bU,F\dQ;9Da,Y<e0@CE46
8@>TF57--dH9aEQ^O#)YK6A^,V6X3<78PU^T5^aO,8O_#K,G=J::Y+dg-RTYYQKf
=GbJ_CIZ+?\[NBVV5gIW^^/:S:T1+,eQJ@c.;Ucb_AJP/@\Nab<?#AVYHX2Ie(94
/2Q49;C0U6]f;F[ZNUP6F+_U9+f(Y<WSQ7C0?_]2g&.]K]FNS\O;F,U#?;H(9T3L
HIY?:,WQ@6RfTQNG]M3>NQ6F#bRCLDE0JI3d645HO-&8N5HJOF#E9OW=LXZQ#TCg
LR&>./O]f0T)PMa#1D#6IIY7MT>95]G/-R10Tf7.Fc:1&-G.#cKF430>Bba0K67)
6Z>/5QXY,BSOV2-R^:W1EJ6NRfeZ(V#3RDS#@@1&3e=4TI]?ZE,d3Mb=EL<:VZ?&
TL.#gN7L5df?#TOY,L4P+M?fbQ9eRH?KA=#VD47/dYGPRgLA4.X0LK:K7#Q,]Y5>
\Z2bT&bE6)^@=>QULH?#@Z:QG)0JScR[\&Qfa.)_RFeVW0BQ;:,.&Q@#fJJ6O1e2
fR6WXJT-bUZ>cG?Q#SI9=84;;#7Y:L991d(BVM?8+N8T_EbV?L1T1R-:&bGTE:IZ
[)Oc2\KF9:e)9.V4LgR4,@D2^H;08<(YJNL^+5dIZ&8/=(^aT5_L239b3K2:e(MA
[VKfWSdaARQ.1K9-K]YFDX#f5/S?+>6H2E\Wf4U<D;;C?:[Z@PRdV23.Ke]]7E..
_THg-OEI=/MBTN^XEGdGK_7\-A:Q)>)G8_?ES\9>dF0D]gaJ]<JPC+EE4d)XQ8GT
./TQ(1RT4Mg(34)S<HA6,JP@0b8@P<(eT&UHSI9dOFD9<>>TAcKU_/3FcM+#d+2G
DKfG:TEBV.EJ;NAOQTSGbM]O&:,BJ6Ta&-;a;M)Y.Q4HZ?PW:R:::U.Gf:>/&dLR
3D1Y5aPN[M[=[^d7M^3I4]M#+bU2,,.3JDUKd\fS]/ZM<6dUZQHF9)bL55?4/>&5
C,N/WGQ49)G.?G94+eP?1PP.8.e,#@@MDfZMOV8N-IcT>R4;M&[:Ka8<NW0L6_2e
_2,b134X[]:\dP/(fIKUG&@VRd23\,L=a61HDgLP?@,I/-b>70&0I56&<=)d7>NO
\D^[7UE(=fJF[[MG&T2dNCZLe6DZ_I0eZ_?X,)N@NOTGLc)5bO1K,;>00:8f=0[:
gC7e:#]9Yb,H(/,3.:]+:BaM>=R+I@[;&6BM[E-5VTL0BT,8N8^]D::KB0&1F4?M
;)-C]<3cd6#(DNaV=-,4_FgJY-(3[<g7WY<UI50(OUTVe.e_G<?N@>b6b2bN?@L0
SC:5e5Fa],5.TR[b/+[49dKI8BL7NQQ..(PO^QZ\_c4ZI6(P9SJO6b8fF=J=D2V]
6T90,XS&0]LF3gT)?S1:PP\JYf;06EfDR/-OD)BC4XW7KC+d]W,Md+Z,BG1YXf)b
<<LBVPLDM:\1-B2]LDA#W@[JeTgd.\=V(XWKTAM\bJAI982(_g0:T7e=UA?_N)8.
W:K+SW#1#J)CgTC[(:IFE_.-@aMc9)>@g?aP_U@cQ#P=AW729/d<b40Sc(GAI)/G
AU1J;T]N[McCM2Zg?MTB,M@fdM7V<:#c,A7[b+7dCad8#9CN3H(CIDZFPAZ^,7R\
b[E_T25?_<L__^;AZ;G5g,A&#T=XQ7>Y7(9N^>GR(IGZ)O5fN=W#eRJM/V<XdaAI
1S.].^;EH+aP).AXZ<d_bMP\#BG1Paa<D9X@>;AQD+6Z(NF1HK]O;C6C)5_VV4UF
W8g(_a6G5I8\:X>\Y7bK?XRcB[87]fZ9:P.B@KN,<5OU/gPK;Of3(e8]<M(\48(Q
MFA_CPA3,W30fQR,>BQO]f8777SGO/F\I:GWXQD3^eO.@_<A.ScB64T,Q0P?Y6;C
f#G?CP-@U7b05NT]F5@<b\-A[1J6?42U:J(D#>IIa>8-M&RbbY)]6L,I>X:XK-VP
AQgV2ECXVeIQP2b0VVBK2S6TJ9T+U/OON/Y7E;FgU?gQ1Z)3JYNQ.aFZ:).T2Q9V
7<].,7c7SDA1.8/@@#^7L&X?fLU)O0.cVa=^_ZQVHBg)-\6Z48aTU3X.SC)J02bO
?LSWdG93_A,8\T2a>DT^V.V.X;TY)KF.>N;8ee?HNAL3]4Q^])1G1;YK,6ga]1D;
<DJ]5R0MFTIc)gb3NC6__FI.DABf@(Y\KT2F^>CAIK&+>^4Mc6\P,K#d58b>)c?I
D2d6,9&@+PLN9QA777<c5d^8(HXZ;5#+?=[IFd<98?=,dP+NSSfO#ASaNSeEY(4-
8D7=>Q^N^R02)VV)]3Zc;QP1[6]NA/X)KT3Q:e8(dEWIQM[&g2]+B)J\.1bgPI<7
4aAe6.2,AP/-\B+7-Bg5^fBN5J<)d<XX=SJ5]H8f,d+\?2W)8#HgLT&W)/P2RGZL
Z?>@g^.-(IBd\56Da84EAL&SDK=QcI[@#^1=FXgJG=GQVE14BL/Ec_OV4gd(82[\
,52BE?FOeXZ/W=?(90/c.:7a&IdUMf#,SKR<cB+F6@6L2,6MS8?5594S#J:#^,>9
eGUE6-I=AQJ8@cVg:\_X7(PFNGa70]CfPT=&U>2:?10X-cf+IOb2UVIA^R0&Vf1H
b&GY&K1E1:>N9Dab9)JMeUE>6(V6YCEHeR52]I;Z:Z@MPd),WB3g2)d+1[Y+WTU>
N;05V#/Me+Gd;HgE9LZ/)V\adXX.@.<3@=&RG&AHDaC9KDXO^>\Y:&#:J2;)\5>L
CKSgH?RE]+A2X0gJO]g6c=Y^)LXe^F_;<CCb@LJ\E;Mb>;I:#=;eIQ8N1,Eg7L1;
)B>=@M=7cD7Q)<&HMTc+PNKgC+K2&6f/(94O^?gE]9Z[WN#EUZJ)1A@;X</ZU)-5
GMYg5AaG,T)bQ6.b\GRZ22_S[BOAL6gP/7gZEgedf7<#II<6]cJHZ7U41N&@XG1Q
.(-aA>ZBDU&)9b+M&/QK7a75:ZVBI&P#Q?A.BRSC@:Qe@BSUBX;c,QQA.V<gHVG8
GD^TTWd@H742]71NgJ&E+7M.9[A1\;(f<RFLQ[B#Z@U@Q[7<]N<1>@8(H>]ONHKb
:C3L8Pa5T/)][=Y?O_+D\],09abD:>=>LML?/6Q_P+LSW^Z2#H:&a?0^:JQVFFH.
W\b0#M:=OM.GM.65DDU13L>@R<\5&-?+0\^MHO8L;3Z/[4M^+QZO;+A7Y73M5S)O
f/E]Af/^-3U7S[4@82bL@-Rfe.?@-@HH09D3DH4PWNO@_8(7IZUP=Of.FXCGJ9(4
9Y,=8]8:L(27F@#[UbeV=CXg[9E<<VN9K=O)X.Qb9DO,YV_;g=EJ#Q5S<H;=d2a+
LKJB>=4)b:T&B0eRCO.C(R7L+1)RU@,c@3C<16&91e;cB9Pg;L1+O_J)g4)+SIbC
,PR]^A9fD-Gb;D,;8#5;(TX(S<(Sg=[E[/PIe\KV1TN.eVKOO)GAa_>IGg:d)V;e
JT>P0_-E9?J4631-@=4X.1;^29_\@fZAHU0gHW\ZaeMY,FW-<;Z6N89,W1?Z[9T]
KCe+6\\g,gfCR-FO,ATcRZ5Z#AC6(O6EB,4QIHcKGV,\2VCb_:]M]55;U&B3=RHX
ZK;_#+4;=ZVa7b]TH](\X+OWJC+&[<+Qb#?QG?Wg3UYP[).4=4;E?-\+#1#OfHMD
2&6BOOZ_.6BMf)fV&ZD<(457ZUHEc<3b1+QgE+dG:KC=#3_,MA@g2)&-8aa-<XY>
,(Z23<Ae-[PgN),?:9R_-ZG9G8(>fS0A]AJEHcK1:+865g-G54VSOCbEZ=IP[-bG
_&<K;;@d^&]dZMJN/&BMAcHg(T#I]Z@TAfW&>eWZ=CP/57O0(^R-UY<3><6d)Cge
f.0^[O;[bGB[HUQG&O.^TW_Q,W?_3?ZA3Q&9#\?6]MI\)@>(T[,4A)-TZ7KMgH/Q
/LAdF2[N&:dR=<O/Q.M4gR+32+[H+?R4TR?[72<KOE,?W:)RT\b.].7Va?1[=4+c
K[BEQ<]-7524HRVP=OZ1V2]Z>P=@6/2,>C=/:e#^.V;Wgb^)TW<CL)=>Y?YJ^S8a
]XSBW)5I2@PE(Xf9\V:1/Bb:g>-YKVW=YV35JaSJQb?;3QIA??X0.CE:7\H0_)cP
N/[_.N@Y754Z7JE2b(Ff,[OaDAgQR]d3\]B4VWe8L:3A&J0Xb/,8=+dD4e9;f<W+
1)ZaR?#1CULFJCL+VVgcf_OC&:\C3<<Y5Z&fD0_d<NX#G=&AbVBc)5dT7(\&<UY-
ffMXA)L;;Sa^X/RXTb5EO]92g?5;^RGV9L#X)0.\T/_3CW#M+<+Gc9GV@>TW=XQ>
8[.LfDa19LL<7E,KXQg:Z8W<4G(,SfXG[Xd:7Z1NPWUFW:fY8+[2<_4^a=WJ<O-(
[O&P(bD)F3J?ACR1,.\F?Hc#VINCge><K3\CG?,aH>@18C&>EP^G/ee2;F&K;@gC
9MTVWaZKJJ<(^e;2<0GI1f)^IA]K]O7e^J=8#:NKZ^^5RgKA0,g(A[b8P_^B:3b;
GHd2=N-&YF?[I_13]\b?;]<cP;Y_\S1123:,-NVK\44WQ+Z-&[P,3M3_\<?5.43W
GA=3HVAN4Pe53gDXS-P2d.LW;>W-?]C<@)7HHUde6JNDR7SCAc6/F>5c@45LE,QO
4S&K1Y//QL][7U:AggH@]9e9@,0[5N.#Te[.DP#CK,1_MM_IKdWaQ(c<Y^#IdVAW
CA8&W&1CIY]-DF=Y8+/>H3FNN=,DQPP4gUe7\3&J^?dJ@+D?A8<Gc67YBMgVB)]<
gV@95I(-YVST/M7U?76NE8257_3M6-13P#VB<17:D8eTOLDX=AVG84>38^KUJ^]X
b5V.R[#V1T.ffD8bL[IaJcM/eMH_bMeg?Q#7D_2X9_G[_Q-?ANadEED3,1#]=aM)
X@dMCPYU6S;(UCNB=]K]?_6YVfLMJ)B6?(f3V-<)B,(4&580e-N.F7LB7)D/LO\B
3BK1F6FAf/FJ5@5V2\UXR5+FW\]U2OEQF-#8G:\e^08-_8e^dNWFI3Ud]XXb\;PC
FXKQ53.-I(I]KQD)T?BMTX-DM#T>7504ZJfWc(faW\5^VbT)eHB7531&P<36TP4-
F[,83LS]FZ\Sf^#Y]QJ80Q+],7ZIQ7MW\=L1g2UdP;@\-EGE:/_f]Ze2ZFZ/DJ,d
3^G4NTNe)+SP>cO>V8C?b#98SF4:U@.TD6WV7F]7@@a7>dVH/a.8RN2gSSQX-BN?
N?Db\I\^ecf@EW?3&K-ca8)5SCc)K7N<.612f>CC+c8#U6.f6&e1&HDM6W?9+I(H
Y,^IHP1=eJ#7c4(;EW:d#<V08ZR)I0>c=e;9_@2>T0ea3b+JCQ7#F0P+=H-d.fRA
(Eb<Rc61.R>2#U;FdTUUIDMQMJB((#LL^W/f\e9ALd>S[?N[K+CbET7]R:QIbAbc
H&O\0L<8(GK556CC[]/81e&f.R(1+>a4>H.Z-0_XQK(_OT(g,#YLJNRO<CSPMEJ8
f#</+?dP5ZC+G7D)3T,RM072CB7[TY>;Uef]IeHb\+,C][=c6C)&g&ESCH.7?I(4
/60Ng)c^^fJ[A>f.1#-I5GI3:7eBT&<GMf;S8YAD)VV3N:K;2&OCG8BOX;b[5/[\
9-_3caJ3RbZcO:03_J9#YE>\g.?7b?4e0G8GNC0e@?1#K7JEg2?:6.DM9>KX>_)6
=EZDS1\M,7VFATHXMJfgBf@W_?7ZC7;NL.T3IePd(G,]F82RCC7VKedGF=0<WNS\
Q+39U6YL6A#eTS/3T41XB[UgW8)bGDD9Sd2.RP502]5USQ3b>Ld?1IZMST?H/_;f
A/Q>8=EEgO/_eabJ]/\_N:&9f:6?PHALVV\++3,,))0S9Qe@=)GKUJ2N)\XZ(-RZ
f6W?Be30):ZWc_0W9K0a(J@Tec(Q\g-H5cNa/SgETTAR&^@_PRE\a?LDX#<US0E5
=eA>f5,6<8-=[#9#ZD,ICZN;2.YRQN?DRIb8)T<c-0Cd3ORF\d-[b8Z.^T&;PF@R
S,Z[U<&H[TV1++KM0;/\K6O5/2XB[=T1bO(,)=g(MG&.8L[c/,_=\VJ<NXWJ(GDJ
+)#3)U4V]7:&4/bM_dYPVCQd7[[SPJ-E)I?7M&(SR:44ZI0^;@[g9)XEGDD.492g
[)5c6RE5[2?XR^7FGW:H(_>1dDEc5bDA190[H5AX(<,\\d?TTJAV\E2Q;2OG=-^\
>b>Y+W(CKGHP.2M;I/EQL,X::F2ECUg3#,7Ig<A&Ya)RC@ZG3E]He38UVcL3f,T@
:cEU#4R^>f8\5OeU)-I]0,T^MC^A)FCFQ)[:@c,36Z?&TY_Ca^:G^?IPD>F\=@5X
f6AHf3Y,VDAf^WGG^=S<c9O]14^N?;R0@#XM/MNX#OT:):(\c]W-,YM8Ke:T7fN,
)g[<;CN78PcP0-#XM1,^g5E,FaD7F4(^5AOYe7cA]SO\TYD=Q8AO.#T4_B/F7+Ac
^8]be<Ra;K0fB;5[&6U63_,EW];W5([9M8f<7E(Hg\CN4RKM<IRL6EJe+^B(EFOe
d8Ja^]9T,;]0]I^3#RF3O5TN\1O2OW4+^QW,>0bC3[-Q@O(10.2)L&-Z\._8)bdg
UC->U=GA9[5a3>e&bA+I:11(=+2_P9/I2UTPG1I?D#.2#KS<\J;^5gCg1WYOW5+T
g3H[26c02K94Kbf4gSa@(:&TF?P3N@[^]B=+dJJf4CS2fOgI0BI/27A^(KfbUC+Z
664DgIX1P[9\J[/OL/PVF13:B<4\;U\>K6+U5HF<UZLBJ@I2:N.Y9:L.ZKI0PL7N
Y>;@;?A=dN>5\.)gH&CcFEdDV?3DPZ&NK=cAZ3L,NSb:b:E<X)?;BZ-V<b-bMSGO
U.6\>8;M37d&GR__3]gb4C+6MLT/[4,]9JaQ5f.>MT#QNgFZB/@4KP\R[V]JVCaO
.S-,A)POKeZNQ\g7YLW\HRf;1>M9_SKZLUFO5SG@)UdW.c:NVgQO;RU8BPT+2M#:
]H#^+,\EcDQT-B,X_;de&,C<Z_2aY3@g7AV.^9O>336(M4ST>>f3c.RECXf/;QaC
HA6W08=IS<@TTPX0cC0/N49Sg6Y02ZNggAE<,()YY0^UL+2SQ394Ud9X;:O>SReK
10B,XB@/@BX8E2V[\fU0NSJ<ED^I#W6;&;XK2G?Pb^S>,ZY3/TL+]?(:RTL#U5X0
W<R#f2BbFA8@/A6g_VKHcT7GIJ^S6RdV)LJ]KR:S?UZ6Z_:J3)BZg2S]09QPPU,[
D&/g=&Z37LR7XOegE<DY::31UG(Q>)aRUe4\?5_]];3NHZMTQV9(MFeB+M&,URTQ
Xc2,<3ZN[^)G]DaCD-GWZe915Xc@NK[5)-X+-bb.d<+bG1L,?1PdB6Oc,1[&170Q
H>F&,Q(J(cI/f.+;)GV<3&=8S+YQ_;LO?DRfN;N872Ma]Q5Q[cW-)JC3@JNZL7:@
ce@cE(:[Z3=2+BEdU6_5S36A7_1H@6T05H(L/8bHL/g/P_UaCTD1e#8Y<6)4>2Ka
]63]5,NbL[&^TVM<(GS;2\/dJY=OCIH+/V),8fc:],CaCd,JZ-713c:68^8#\)Cc
>dZ-4,1,QDcIKDb<NNN7b3Ye?)?Ab>bM)gP&9+:Hdc60&0-[&#.#5/EIEAZfDORf
VHKNT@0K/]-9(9EMX^;,R<25gV2gG1(B8.HLF4IT0ANXI1/4^..J?J(J09XS(.:W
45TBNH,[M6HQ_,34N+-.HT6\37Ha6ZAg(OI]_9^:F/.>AVL8Xd+(e5K]c)\UeRD&
-6.[IZG#Q)@O(JO>Pa>WR#_OB3?<6@:I).WA-Gc&T5GXLLV-+UVPP1[6cG:<H^LZ
J]7#>[C3K]:eSU/F7APO_(#YU?)N(<OES/If85+X.W8_R-5SQ]Q_&54T\VXI2K&,
J4ERdbO=4b<;+FeM;_#\RF7a5.55,-I_AC?J?fMC-C5C<+SLbV_MSF3GMY482ZHN
KDC6M0AWX--2_,7WCTL<O8CGfP;93IW>LceBB;1Z<U401E;2WI>G4JN&R=_H?H7@
C;1FbI_1VYETL=V6=<Ac^HR\^eI).7beR-WTY-LZ6^TT?@b.;+=:D+,U:_2L@]84
<8+b-d]WWTI/DV_-g[,B/8\H\8J-;:@BIdBLg(Jc;NRCg<e+&0&Ca]F)WDTB+fVS
RK(3^?T,;7b8XN^5WPQ#S33>B=5KX25c>YO_E9eX4BQ)(W#Q_R@a5P_aOb[J6/C/
;&?<E7Q\WCO&357&023]I8b(8dHP4W/IC-Uc7+cZ>\[BIQ((d):WRfcF;W)8R.[g
=a\,9?;#0Y??#OBDSFdV]4K4LKN(X4bM:AKf20<&Z9#Q@#W2;8(TLa<XfIH740I#
[;(=gE=6cVY^UF[OQ2+O@;?T[MUC^>a5&#f&[KA)=B7SW2a3-\cGHS&2D+89/G+L
QL>ZQ/>cE^WfM/PB_OATeZCRD<NCZXM<2-(<G<+WEgM482f>3\LJQI8X8[/TK0]e
ZMa9<9dOQ\H#OONO:F_W1Q@)<2?6T/)d2J2NP?g#J>N<BF](&LPP&:8JYFZf<;^g
Q-_LQ]V)^bfAI2>EV_I?G[4(2-GFNV=Sg6\gZ;fd?Fb@9X->W6=(H5JOgCTOc7J-
N)eYQ/(DM),AY5/CAH>9A3T6gS&Qd#2&N[ab5=)6+D]UUSE&O+CWBB],K?JIZ4?7
UFL=b(PO>&UL4&S:#gB(ML-47S\aYHGge1)WX5H/^[IV>TGeR1<MDE5IN?US9P=f
XGcJ^A+MB8Z&UF/J6ac)G_@):bU+;REe2:9+TNIOZc_+RMAX:cCQ/R27[eC^aI_G
D-BC36=<#8Y8A:LK73Dd33H+#[M>A98BFCFD9EbDc\e0eM/\-KQ(-cV8fIb_&g])
17.-WDSJ:@[37B<EXXc)3;/Z_f8/-DKa&>N<^aB6/A0(aJ,]/.9Y\4d:,N:;45;H
G:;,8VHAN,EWfK3I5J&I6bKX/+V9A.Z=^M8XZK_Y2L.K.J1NY>8X@_,_f+;TdIH<
D:P[GU:>H6I40@=a/Q(ZDXc]5;@W(J:L3Y]a;@LV+D_@66J/C\V&8R:2f8Tg1AeJ
3]KAbf5.80G9#1PgI5IM?ZGDQOGW)T<1-A>^P4N_Gc\PaddGP(Z;c=IK=K\c#3>R
.+6?66LP+0C[73P4(PK^:+&S1_J,f&Z+#1@b+@<?NQ#D]^#.OE7\U(R)KQ>]LC<-
U;c;E;O4#8S+2GH-ANHV0R0Qg.G0I&D-NUZDdUFR3#NVREa6:CM+fCAH\]XPO5V=
FeI9GO&>ec]>HT&37bP[a+BbbCFc[/8b2=;LYg_/WN(-U=cD0eaU>CWGQRC^/=&&
KOM(;^aXL;)[=#Je)P9QI7=#Z4+f;6LN82\>Vc7CDb1D[6[:VG4KC47XBXA4fKR#
\]V@92?G^WR,J<-\/2eL9EEK@;4AbUGMTN]a)-RV]-J<^C:GJ4gdaQ7fLLb5.N3(
01JK;)6_\]eS8:9XcN(RH]1(OJ:E/c]=/OAK46VeEUB&[0WdK/9/9;e.HV7VO7NM
1GEIf811GY^45]CJJ+2S^FIO>,FgF:WAJg02McF-HQeCQ7VNY_K0OeV>-4dNT;,[
>-fX@KecQ@_YP(H\JZ?XZ3gKX2=:7g?e[Z1.cDAF3Y&PIR5gDT>dUP8)16a\>g5O
OTD(@^WaI^WWEU4>H9@d?Y#QZD;G2EV7>L:)Y7TKfaES_1-Cf[M>@N,fYBH:P/[O
H\ZX=E:7UMV9.MPPVD)>dSg[aF)PaC1(D:8cFAVR^NT>eF9X5U4&<GANOJGL4ZD@
BJ&]e@(&R^JK-e/CSSAa-3G+J^bc&#=2@20RWG6^fcBRRE<FP#G7NNW;e5V=M/K/
X<&\b[_dM^\/[;1H1ZH_JS3+@@(1dBHEFRad_\L\PI]2-dQ(0>\+GA+\[V&^46#I
CNY,TfW78XT-[Z43IMU10K^+AVWRHgN_29d(\G02AQ5\)0c3da=e(6<=E4G>.2=5
g8P,J,(-He;a:M<G#e3ELgZg\)OG>/,b_SJ7K&M34W1^J1NF3OSPQ;P;6N\?\@7a
3^bD>TcLY[/;(+f>@XIZ5eWgHWS^9b[3be);3See6bfMYgbHG.VWAJIWf@cWE\=D
[_UW8BE?ODY#<YP]/IAV3TXPg4VVLBZKFW7#60],VbB[4M9RJEZT8^V=)R]X#=E&
_35LYVX])^YPI+]&P>[C_9@O+g8=_P5RbfAVP1A3eF[Kgd_JVMaUPWH/U7fC@X1d
De.]\QOY#/+f^Z2=-fJ/1GgGV(eY_X5.Q=U+H-&3?Z\JV7M@[NF.[+^#,_8]N1.Q
6PI4Z[WQZ?O]LPQ5de=#]990cSJ@]d7MNB3,CWM=?YBJ<E+_HgaL1Yb.cG4A_EHF
L-#SbL[GN6?gPIN0WT:G[=0F5II0R&CU0g<IS-Q92-N,5=C<=]MLRZC&(?K_2COg
8?1?abA0E?Y6,>P:AY+RUfgE96R3[AeVf@Vg2&(^cQAUX^+eBM(LYWf<I#93IS:A
7:Q/Yd&dBUB=S?_,<VVe=?Fc06?7UZf-TB-^3XWHJ:&/_/Q<3UJJfg1CH\G1c^=X
RDWTCCR?1gX5If>a^L,FYK0?^=LIYT+WG-?a4?daH?TIa1;G2[XQ+@XI)BFc1EBW
=;]IfWN?[99C:>f8&@P?bS#T7fc/IJe,dWgU^A;H;;Y(CLD@YBW<L3^)=NVOeS,,
d=0?(_<CS=>_eOF2&fTZDYaQCE2=H3NWUYYKCc::S\PWQ12QS,]2bN,.<]2C]O5d
@85LJI_SAI^Q\9CeeD=AJYe)R8+NFX3B9>D)8B^2aP(:=&A]-K:.Y/A[Ld3fK8.[
?G(bH:PG)6>3]J_81(aVCS:bfdM9d+&A;Qe37U2fS<1cVE:ONg86BC-4L#d[D:dd
.V==-UQ\;20M=#NGaI_+KcWOXQNQ8PIQAC5fEMG-C?TZ)L1R_;)QT^AM6(O0RId;
W9K^5,3NQ2O<K5[.f7H\796Y@LG7]gD7_9+a]Wc1]W(IUJMAHVK+ACTR-W;817a+
X0,IbO2X(8eGQW(8BRWgb#?@^3>:A.\HGX9e[DeE[:5(a:=B8d(aVLcGYG:>f;0R
Q>KK].YH@;f7&/-AeA3J+GW@_DH.W)FY@(&:=.WJVTLe0ZQO?BZQODAE+;]YEHS2
C,^OL7J_#+fD458#_GBGIEXe:YRQJ#^89B/OL<#<>cZTRUX+Y::-F&UQ5C4__6cf
M6/@,>.e>^J+1>_G_6gTe6.E0D,:\#4(5b:a)N40WJ).0g/GaN/4.@R3B..O_MWV
Ud0.\[S-HOfMaGR+[UK/MY:0PRb+g3O3G3gJZ)@5N)LPN@0,O)FL_aA)+&A]&bP9
_AHKI-U3NELagdA^V=I_XK9Y39>cc9;4-;6]W=)8-1/C?@b?c+>OfB-]<)PJGZFU
dAH;XM6T_a4f(<5TAfT,<CbeO>7MA6-,f&+-D8E?Q^&;WM982)Z4bS^),)>CFA#(
aERVOP@=R+7HD=FIL8U+[6=Y-Se1=(=FTR.E\J;85#.O[RR0gPNVf]@_JY_NIINR
FGaG?I:?5?AdJ=d?JTg6JGFH[&;>Tb&3=[[C&ATWYZ:WPOFg-FWGJVXK]gd];AJ4
_&?2ZSHH3A19.?I.@cP+(13=ZZ(S66Q7<F.;9[,C=<TE#C.N\f/g,I9Q^53/b#.T
O/.BFS4TN#\0PN&3ccYeU9Z72H(AL_:>FG7BD7[=c3PgV>JCR&RCVQB9J[HHA<)_
Q)R3e9=a<>6C(-Y:<W8Xa?0EHEPJY\]3I/5.2C5N1Q+]Z]9^5+;:I+A,(<2BEIA@
CXb#3Zb<.<#SDc@&3K0KPgeH?IU&FET&CaD@gUC6HBeUY#9:e/\bVR^G6#4XQJZ0
-bLWSK1DX2JVA)0]AP?MQ7@Nad5?1Mc5/8D(<F6-4Y9\[](-HQ2gQNQ&bZd[=/fY
G,--47faZ?@@b.-_eaSCaN<B)0>8ZAO0E4G>OWLZFe[g&];dU2?Y/R:b7\D^JDg1
]fS6ZJU-&Q<A]aRJ\+.eZ#d3:_[O?eY/HZ[)ZUMLMe;IK2J?3bD1/)BB_Bb2dYeG
39e>@J1<GM)J:-8O^CBA/fQTP4M8O;&FdMdJSGSA=LY9P8[(^JNNPDfI-7feVa0;
MaBJU_fD-VA#,aXJ0^F7I8]XIJaNA=)D:FIXEPI@^9\SSLTNeTJYR:N\RfKG3gd=
cGM0]/fX(E7JOSa2V.\MOA-43f(>N<.QH0#2e,R?K<=D]&Vag+Y_@7=&B.IG)aZZ
31fU.(43U=0].XRBW[S&.EM2Z&7Me-:MU>H8=U[0-dG57(LYQE]STc_7[Sc?Rg(?
N@Z;df34]9[-BDOe7Q3LDM)Z_V78@PUS8:Z,94E<E^dd0gINU]T3EHVO5=2<,eCG
<5-@HZBgA=H60(O=;Dd.YZ;d9d[6L?A+e)f_DWEXYDIHN\9L&BD19b:&:[M.BcF4
gB?YcCJ]XWd6.c4L(Vd+W5ANb;d.bS(6CQbU:ae-LRZW[f(^TIN_g@7QOgEG[g>0
JI1LV/0b<1]fM[7MK<2A=/TB(^-6;_DSTc++fF,fb3>bZ4SLAS<-:>._:Wb..a[)
3RK^1feD+QGQK>b@ATI?3fBL][:L7W@)P<-_d3fG(WAKbXf_L:GaC)5[^5c<Fb6I
0+>WfJ_BDNHG7QKa3Z(/J@Rc=?eD:JJLRJO]L,5dJPG(05+6+SC1Z^ORbB5^VNNC
FM2HN)f8M?7IP203IE<3TL954@52D7g:ZM79GZKYf[AZ<Zg=e3CLC1[aB4+^#4,5
^Z;FPca@<@&@d&G\e1a=\;[fYSRSLP<f4:^8=Dd[)OQ7>-\bJdLbY<86DWH_P-96
]1)+CY(1H8//RPAA.V?X\&+Af3&;&W>HFMEDI+UIGd,<#fM6]]JE^3dK\?A-S0d/
^73=1UfRJ_=0ERD-7daS.G8_]KG.8;6C[LRLQT#)A;OM=8THd4DT8TUR+=8\f#9:
?4:5MQ0>Zc/2+d62(e&^<T714-52Z>)H,[N)W5a+-HA79WAXSM/_d_+.B+^J,P7d
F+f>7DFKTd^e\=M5\S5(:Pa7Z(?20OE.HCd>VR/Y??@#++P=;A5O#UCcNKFPc9:,
cR[#0-\(\L97=QgRBKdG:02IDDNZD=NOGR]gcX3ZN2Y>RTPf#=BX;D./+5L62X_R
^)H=>_N]-a=8?ZO(,e>HCZ019_L>]TeMT\[DW6CK,K16#>?(C)R+D,9R.6]gCSRR
BH,L4:EZFPRe4c4d.P;U;=bVc;P?8W\5DXB&__:SWBRbUe,E9b)4OY@B]&5B496;
Z(JY(R43DHXRD\I]W),)P^^E;/RaY+:O>W].RM8>(@[XM>LWVXOZf7X4SD_P>)Q/
:&OeK^DUJAIR8>cD]bJO5]6)\?b3\W7c(#.Rc^faU;YZd026FRb^34WI#9?^KV\E
IEU5?G&Zf(3]JbKHY_A(7-8<IE8Z6Q?4Z0A/+4gQFBENJ(WM1DAXJ-+10Zf/B]K3
f+91KIT#W[DAXO18T-?fKCT/6H7CG<5_4^a]KV/=SRCKKbK[VYDcZ+Xed.;._GKP
6@QCR51FJP141E:gOLeJA2/RAG;Adb[ID(&#9[f7#G,-3AH9]\X:C9(2N)^1_-)Z
6gD;A5_DdAPT6I3\@C1Ga^&,_B0<N-F5M.BP8dG1,e4I&GQ(9,+JXHY@@_DdRWGC
=>3GV0CR)04)U)\.(3e9CTPZ,#]XeC)\KZM5IbbMDWL<eWF1bBT@I:\7IRIS;C:Z
D6ZeAS-I7D?(.5I8bP8fWWJGI8SOJ;/EKJ-B492LfNU&R\fCZEMS5,8:AAOd,IgB
G:<^.@?_9NZI0ET@/gdZ4_M?PR5EJc>:QFT5)^K+<=0?7>QHe)K4=\f1JYWX;ac?
NK^LH71WSIfH_]Lfg-_>g[>OI]>SK&-I,@BNZX([YDI&,,:WJ/.O98XTg<-6W\8c
&#?b6&f0.?5Q;YBI@_1V\/O4Uc_HIT;Y+U[R3K2M2<W@^SIcR70\U5B[EdZZDFH<
@4XMSO/@4;-D/dIL3,AJ9R\WU)[\MR>1N@Y&:@)LWCe1Z_Wd[]aa^>&I--L_a2K3
+TL<05(ATKW()A)Ma@^dK/O]FJ61Z4>0bf;;)0M6APa3Q;46g=Of[9,DCac7Fc2.
eS0I&Q2W5S2&?-0.7=1,S>Y)\d>TBgWRa?,cS#bM2/d06T&G4#+@:aBD\3XDX]GS
Jff3WPQ#XU^8?Y7QPX=)1&O8bA=Y:WK&g<49fN@.Y/^W:aALZHaJ&b<,_.8Xgf,.
e\2\5GDEG]8Q-J&c&3;IYd(1TDA?U\=b84ZbS4E^=Z-M9H1\.R@aUUdUDMBYR&S,
Y.+V8ZWQ\C^=e9ADaK#,K:X@fRK70W5-0N@),]Jd.GS14@4dXOOg5Q.#I^dOKHW6
?@;^-@V;aeQ7&/K5ALHGU5;1<RE88f;@7XLJ?^<)Zb[bc1ZMR6T7+4?3;/SXGgd6
CA6^D/].@.JN=b?,_9\Na3]OT&VbXR\eP>adbL,D&JNa2<X+1A1<R5M;&b]3D/dC
O1eWL^-BbF/_#YeMIcB4H8XVeO(:0=.2](cOK7J&>U[P6DRX,a7::5X2PO\A2WXU
IO3HKHOT+1J,acUGG(Pa6O_HT0QKX<B,YH]^#I.BKFFX_O,XWdO]YaXZ6a??4\52
:C6gK)]e:XI]fGd[R[<3XK8ON5caBAI=6DBd=N2.7U+V]#KFdR=a_JPLW^KPJ.LV
U:^M?0&,aAM?:N870f04Tc>MI0H/.]KR>Nd3QeW\M9cS^XAfBKAd61-;15OUN-[Q
9F;]UMF1fY)cS22RX-#7cP+1(E0;Dg2@6N:SO-R=RC+6>1=3@TQK?0gZYG<gTWYD
H/E6&[5X7T3H;FOPE##a2ZM;Te[=:SPdKXL^OZE.gU7e#1Z2X+NBBI)b8ST>NdY#
-FfXSPV]GeaO<]OIUFX1CX2dfE[UE&ZU_3YD9e.HNKQG2P#U2/5V..c7>)7]MM3F
@7UZ&BPCHJ/_]<).=/Y0IIHOZdN62T/f#6\;g027X.TW4-XI.W,95/E0La]=Y:f3
G)3]DT\+4Jfee[8B>0dW=VGO/YbOQN0e^L1?(V5:e18E7;1^<#H3Q2Z+,^/Y/8,)
Z.</Y^0)1XYaU,+;J#NEa2Z\dC-G3+Z1V<NP9gfFaKYJKN-e#Y.R?R?N2[7B(=47
FK=UC],C^4O\?W=@_6;ZR0K\P).]T-@U,O]X\C6Y84@>S<]F;2@[S-F6&L8_b=^?
(B,77^b=eUMJdDGDZIPCQ\,4.^>Jc,2SbYVb,Y+JSF2f&F[?1PT<O&#<=ec3<g7=
E.gVASCRR9_EA+O\]=R0\5d-efaf<>A7X,51-D5VJ:2f)>JL,,3)ENL&[?^1BV>R
4<3\LPY[ET/LSN#RP#:B1_/:;@d0TcBK:X5aS),V)gJe>5-.DfM6#,G:BZQ1.Nbg
M<?D_NF5#-7_:\GXDYQ#@B.PW#&3Af;3DK/?FP>ECU4>.ID<dN9\gWD(+6a>gJ>5
V5=SB@4c.:UT_4<eH6(.CX#&]>O@V:&.PWJ+UNUGC)NFS7\:WE\6Sc)_BLV+Z61C
bVdO8[?W+.5:O;Ca6dR5O(\>-#++Z,Ud\)9;BFd#^2>5^J2U_a&;4URLKO:PIeba
_@)9Lf::5J:\+([F7,X0_:T]ERd9_&f13TPbT^(FC.@]>C>#fWEN:@1aHbbWXRQUT$
`endprotected


`endif
