
`ifndef GUARD_SVT_AXI_PORT_MONITOR_CMD_ASSISTANT_UVM_SV
`define GUARD_SVT_AXI_PORT_MONITOR_CMD_ASSISTANT_UVM_SV

// =============================================================================
/**
 * Extends the base UVM command assistant to customize it for the AXI Master
 * Driver.
 */
class svt_axi_port_monitor_cmd_assistant extends svt_uvm_cmd_assistant;

`protected
Z1,Z9dfgYWT[\Ff:T>L;?10/#K9LZ8JN^fcOaC/e[GB/3.2==B^C3)EW3Z[;f+cC
+?<EKf1@[#efA#DZQ2&ER_A\f>Ld#&Z>CUVO4PY,7[BGPGL2fR4UQC1EA\5@W9]7
A(L>A\9:0(R9F\(B@)_Z@>AE92?.G<@<?SQ\9cY>;L@_Q/VDDSX>I.):YCU:A53W
KX=YIg=M9I+00Tf_a^9->9ZZL5TNJc5E@XG,TUNI&VG(4(:(]U[0WFcga07UY3/P
Q=\XfCGEWQSB8L(A9#d:A]aeV2&>Cd[@g-dOG+VaLa#IdV29bMD:RL3@eLJ=)\UE
XTAD#PafQ.V42:1Ja6M>8S0N\Sa?+B&2=1^ba0&gU0?-_+YG)799UD;X#+4Q-1@a
31^PYd?.KR>\8IcGf6_/O:5F5XH\Pe\4+RQOc@fMO>1C>UJG0@1g7f?d9+JdXD7\
H/fgK)MIYRT,Y&GBYYL_K/>[85+[1bWHPPW\XVVDXUg&U8[&GWd6GI?eHP<)=&0#
6XYNAVE[YQ8YTJDV5cVB6IAAb3,Rb9LaY6+IRN,+C>M#fR+M2:]\dA#AH6@EK^CC
?0ff8UXdV,ES,b+^0#9<.V[AT[VDW+.367(V\da^U9)\IG4GQf&(d?\5BO<\e8&S
\B<YX8QTK_PSRKR)6X8E+08\ULSeG?2R\..YgF6:QI6?+F;e.+b6C@>e<>(97]IP
BWH].f/K:L?,WDRb>K/7+;T1>/J:3]-N[O#RRF(<0fR2^^_7#47R]HJdN[^;RZJZ
^#1:&)9:]TMgAKeGDZJ.E#L.^RHd?7ad>#gA.V3Vd=,B@LMZ:09>2]W@+^A2YP=#
X&:2GfKTb)Ve,W-UBIe3g&Vf.?Ib-R,cg6:QQ(BADa7BH$
`endprotected


endclass

`protected
eX_V@@42U4(0ac07=#OERY/MQ0ZMda9+bP&]Td-X?@_QV&WG?,5T-)5[GO-AG+]H
c],7&cB2aF#^OT^<#:?]9CgL@NfPQSa3?f?F)K._7e/4C@MN-L[Oc2([KDRR5ZXT
72^Jacc5:39R.(P3fYJ-5K.5XBM]L53-H1VRX1ebGYS>b6(Z++_b1DIeUA]CCJXZ
?\38>3+8P</0Y:QW,SU+0F\1DXK=e63P44-@&LU[Q;Pe?K/Q4gM:S/RU9@E:\+GQ
+6#:9]Ha,S,+cY-)&^c9CY7.5]5)Pc0A]MDW2d)P:a@QS7H#)DLFPd+DaNV46]0K
0XAJ7?\G137PCg:?TWVXe@eL@Y;8B;&7_,HS3OOG=RO]W[DN8_7cZZ@P\,YZ\B\P
M=f5EP_5ZQ;g]fEP8/ME9+0MNXY@AGA#f)>PAT88e\?A+AFF5Cd&YE@6,5_Z02QF
JcW&^ATMC7G]F9GX,WaLI>)0A5bbE,N3X,c30K(4D5NX+>M>)UY[AKL@4HQ;.2G)
edP:_T[IfIeX+M-(T7SbX@RI\4SUAY7dM46665A^.X&,GI.+1:]dG??Y9Z:2[ZaK
_@2;/3/W:X2)9a3f4J-RIa3R;dSSG^ZH)c@PA[[NFZb-J[W<I-M+C_]=6SU3.HCa
8]@[J0\A5JfS<\b&,F/4)=SUe+Wa&WV[CTJ(Y0Df)dfcgYC[P?#B/M4TT)a:XYHB
8O]8:,LQJBSNV#KeJ+4Mc1IW.(.Ff7J0(LPd?;_e.^gbBFUYJ3Q1&2?NM08C9d66
.6a8]>YV<DA>CQ(DA5]b8#AJ.&&/cBP,.HL4?RB4J5]A,,0=0#DdFY3_1C5TWTV8
-<a9b23GO(CaaC1=>>gWBRAXW_:eMC7,FGaZ_X6O@,O.3(_<Z<&(PI01Ff:)9GCP
<;T^-ZS/U7,WHJGC4X5/1dc75\Ca;OM=CRaPLQE8(?,]g6DL9&dSfE>GX(T]KKY8
Z<A]#=#,6Y8[^&Ca>e8-L8TV\.A+_]S]dXcY8)03a.E<L<V4:)<[QUVD34-A99Q5
Z>0=>PIScIc,JZ4[0(38MVYVO#7J/4[1.T]af^\J[W1/9KJ>#(W56-OUX977J8<\
L9AA?.9+@XUfaWa/)G>UK]4b-6I]=2W@ZYRS5<Xf)0V(N,0eW.-LL3F2#S;\MY^e
+-bW+8>S@A=^d?Q]UJ:\V[RTGOd.X+daU.Z=e^0Z3X6T)34NL@-d+/P83,5X/33,
MATb8^\@DOTF3CGZAAYGd\OUI/eK6f8AcLH^4S/YWOU1W_SK2O3bV#Y)I,N1F7/N
R^O;0?<5[K/PE17CVB4.IYFQ-_G^)U+\=7)<]36^OPBUF]FYM4R-)1e(.7NP+Z#7
0:R#G[V6?[]]d,_&?YVEP7>^K?W#8K&U80,48UIFO8MCM[-FHg=T>2eUaSd/09J/
-=##-[+Q#S;eZ&O9<^dQQQ-5R8#::5e<EQHI.W&/MA8C:Z:_BX1A;3^KC4eCO5-L
IFK&GM]087:?3::cJ#aG//:\>+>PV8XZ6>QZTDQ^NdZK:Pg5</MYGM_;US/LE8F6
/-<37I;)029^[&Bgd8=ZOQbP\?BR3\NgG(cdTGe)VPX^2ZD]?Q4N0Xd(#LX;e;;8
>LAA_6/S@XaaePFL8(T^[XHL3J]6I)=;.bdb2(4IB-2E8dBMTIaJB0gDH))6(W1.
3+(K?A7@,/(+.(c[M7C9N-/SOLQ[[Q<Q86_FaC,.(Kb-8JH&E17R++G.T3Z53?+Z
&_^02b\Q.3>T)P]A\Y:^CcV93d]W@):-(FOeOL+A=CN)]2VMceDa[Q<,<R2+dg]g
A\FYW4S(8OBB+N=G_WYQP5/^H&a4T5+M2DIaRY.EOS:==H9Se>,CKZ<,K$
`endprotected


`endif // GUARD_SVT_AXI_PORT_MONITOR_CMD_ASSISTANT_UVM_SV
