
`ifndef GUARD_SVT_AXI_SYSTEM_MONITOR_CALLBACK_UVM_SV
`define GUARD_SVT_AXI_SYSTEM_MONITOR_CALLBACK_UVM_SV

/**
  * System monitor callback class contains the callback methods called by the system
  * monitor component.
  */

`ifdef SVT_UVM_TECHNOLOGY
class svt_axi_system_monitor_callback extends svt_uvm_callback;
`elsif SVT_OVM_TECHNOLOGY
class svt_axi_system_monitor_callback extends svt_ovm_callback;
`else
class svt_axi_system_monitor_callback extends svt_xactor_callbacks;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new(string name = "svt_axi_system_monitor_callback");
`elsif SVT_OVM_TECHNOLOGY
  extern function new(string name = "svt_axi_system_monitor_callback");
`else
  extern function new();
`endif

//vcs_vip_protect
`protected
?Qfc8_XM<+MSNRTcABd+W<5E\31I\2]E&S2/I/F>IAD;JTLZQM_S0(XLaD1GPFEU
XGZKEELRA5>T7DVY1FWZ&FDOJ42L,3J(I9@-ULE;L5;K]ca=Q.FgL3#FcB;.#JBP
^UX74H+a&T)fgN.:#B=]fMZ[3EGfNJ@B)4=/0=M>W_)gV?Z>=6:H8^_JfUN6<QNS
W?X5^GHc8042@^IGJ\CCUPAPZW(M3W5=W<L4QW.NFL0<LS#E==GY\&a/:&(9-L,/
U4CRW4)HaN(6@+#;/3[d5.dC)6D9M3@EP^5LfT8V2Jdc<UV5V4OVHUeUW)Sa1b^_
](W5GC.4bVSC[]:L\/&642eC((fE80+#<5A\DY6/W_QDSSF)&Y6UOA6&&I]_<XZ:
3X-MGC(:@DO80(g4<Ae;<W8P\A8,XXa-aU3K?HcYEO<:?1OR>>aUIedP-1K-ae@3
QFI6#MKdIUZZS6b4M)E_EeVI>Yed(\A?7D)NW#C(IB]4d1(6eM]GB&Y^)(O&FM5\
UGONFYCV\8ED7Fa@:HL+GeaKfC-:K&>S@S7WNDgSH]^:OS]Ia;CMPefDcQEEU^Ib
)X\2^QAce+C3:2KZ)QMB4b4ZPD(bU17(WDIHgQ[43e=9I]2fLcdfa=TKFf<ce:]2
ae3W<H=^a89BDLb.4G:>Ra/X;Z_&S(0-b\XZHW5PgR816#8S=YEY-IHd3f<IbAV#
ZgP@<XU6e^&e+:JW=:>;LI?EZS)MWQd7^a=([2,KcFHHb\FSB5MLS::^R=W4M>2T
BBK/GUEMY7X;\9/]L:LW[:UL-I0_1c:Bc.0Z&S-,#MM>T.=S)C1@)TIK9B+<ZPX3
+UJ,D(,\[,/5_6WBZLGF31DT0RP751VPg[:T<IVd@G?>3N;A#=2U.UZSLY3YPC-P
QU9.O1D[BT3<,A&7d7@_7GM]I[+>/75NQM-SY=>Rde[E\[_c/\Z6Y:PY)f?gK;?Z
UG+a\.]WA7FNNK(6#OC4IDT(ZBA6>bWW@V_b@U(YD#b2\U?d-ILH:7TfgAF6JIX<
)M/.,2D5-efGT4CT2-\2C6dE@fIL=>ZAT7BPI6@Pe#(LC7S#L)BO(T48#\Aea]#[
#:/9\DVQgN]<YH15MY(0HfAfVIC2^PSBYWNcAeKC.)</6H7DJ>fc/dQYES.>g2&7
AXCfG5L7D2UTUNg.=gE4P-TbXB,,=_HS(GZI?.XfB2<T0C>#L9^W5cGLR_8^YC:\
.:AXON1Z9K@IcD)KUCQW#DMBU1?\O9.HU:cac_9aKAWI>2RLH,#M_7P5W(ZfEYd7
EfgIW-#7<@XZGGaDTeFT;5eVA&^RWaZ0?4EcE=;Ha\(A1W1b2d#\WG1S?;EI(\_g
/P952-Z-D3R8Rf?@XLF<QW?+_UPCT;LMg2(Q,D9DL7N(f/X&aTM)XBJgO=bL;P0A
VaF5fGg&LDFMR4N&R3KW-<(<]-#23[XV7F<4Yb7&EdX^7LHI]ZIA?I:eY3N3K#H.
fg1a\MGJ9faTFF_A1YJ1Y@KY[B#cD<[:D;=e#Q2Re[FX?98?3W[4\SL?3\0:1+RX
C8Bc5Y6F<)U(-TI:>417CK<[0a_VcPU+I4P5U=/+(bHJX>=Y@<g35@:JW1L@YT58
KJ?-42ZF:]QAHQ6J=[]4SSc&IS/BWQ7X>5(ZI1R6N/_7\+PX,U+S9LWG(WTTCdBG
,1-L.SHI;^B2(4+]gaK8NTX,c<Ff\A<D5R2[-TUTGXEVRJ2[aD]X1JWYZW0-CP99
eUY__TIU+2UO&dM6a(CE]6e4RA8?024IYaYgS?9:]RKIRMgK\F&AM;5JWN?N[FJQ
@T2cEM2[])f9A;><HS@Q@g?6]D62-+&)b4#ZN/C&e]_3N?RP.S/)8H0I4&P7/;B6
e6D.[WC6)0-VWOe:f-ef@<E;8(,F<ZODCfg7QJED[VfFLTB4NGG&IV_@71;)<AM(
V0PR+bfd]\V2G5C@,AP6FM]b=8@^fHS1#+^Q1c<^a,JLARJN^@M0b61b^W\^YdVS
:?=5J<4LN80Q=:dGNDAZ(e<FE^ES[Q-eF3N(I51A_^K/VE8PFF^/[R\6CXcWHT)G
DRKT,B-H@\ZRNDA1Z(-(0JWKS:gWI?REH.?Z&,W6;XS\,>9,/8]c6;.<6#1dHY7\
HeUaAR6ebR:Y<9[873U2<B^:@ET<b7]N068DF+BX2eO-EN=G:0bCfL5\)@DH^M4W
gc_L4G/gKd16DEBZ3U6=]+:,ZI_gITE=b/^_7:d+U5(-aZ1O4J)c4A&1?PHaQ_6,
O.^5EL554#;_TRNDTOa[6)NSW>E8943XOA-1P3c1V;T:@P?O[.-H=,Og?]ZS-c[>
TN4(CU223X<cE0\8b/&SJ+Q/LWV4+(GeE,b]7U2@aac5VZH.d6SfP@V>d6]4eggO
cXNe-^)D<CL:M#N6\WVHWGAV;I&3GQHAY/S2><DfF&P-1Q<]NBP\PI,WdGF(/+=f
G^gfA_8-P4,DZ>9_+D7::9]@>/1U.]HJcOG[BXa4[3QYa(R:Md/f48Od<FAfcV^:
Of\7]d7[+WD&5fY/@>Q)>>9+HYTPDLS<5-0Z->aXe6bUAf.ZRK2.dJYIT^VS+ZUD
&9&T@\K3;aSB#)&HR.A9SJU&?JK:>+:53L@g@+80+7N5?6?)Y\0H5)#2B7GAD=MN
?eY=>7HTHR0TRL9dNNA;1>;L->cS\T->8,J\PMc/YA^-3f.LG;d.5\G/1D1=/KCZ
9=:)e+GPD+8cIRU1]<W<X3LRCLESda4F,8DZ/eC-C8N[-W4<34@1/JVcA1LSGWYg
7.+7Nb0[LXV20\dAHQbe5fFC#G5eI&AL+5CN8#0W0T,7[710fbFB[X+WG@;HM?;&
E1P,HSAeB[_JYfFMGFG[OU);6Y+Y.=4R[R(c]b^=T<8D;f9Tcb>F&H(?-AA;>.bP
Q908XTH-P_+O[gD;Q3/CI]5K&@N6f:?=2/.Td4:RQ4\J;(6/BO5,\VBW^:\N+_;8
Gc)XQQW]:SM(a:,>FYf5d0B8=6I2X,)b#?faF1aC_0gP<LZcO,7Lf6gHD]BC<7aV
gD]529O[Qa64H(^V=5[\5D5Y>E[dK8_#GBAaZ(6KP/\1:1.9)FZI-&_-_W^<XcR#
Y]L/SVZ7\HCHPggAOBO,.FZ>XNV&S[MWV2:862;\42AI\7,a37aT4<1bN@g0&VGE
T8;aD[-K8J2)dfC5:1U;/DI#CRO6(6B^&b?&YfIL4#5eSaJ#N>b:ZV&98(e)16AR
3F?:c#\aFGP?:+TBcd8b0J2B/15V,C>9C?3W)ffdP@^LQ6eaDfKNTHVUJ5FeGK[/
M8DYM-5L,8.UG/<.&,F6,6F7Wf3PE9+>La@=g;&N:C\XB0EM#KWHO9/Q]1]T3T?Z
+YE/J,4V>9eWeZG)aTO@YfU9=.J1=>P2^ZS#_,S9DIE_(_DFgX0?,P8CR,HcDTO+
2SP\ZRF.>KPNW6SWMXDJW771fb4?:IYG,:\eK;QTIIO<V52f74)6UR\2Z1UW23/<
X7I2(bP?cNS/BDMC=,<:gUR&-H5d^(\=9E7>M27:XH_>HKL]:/0A61F02eDF?PS;
_:^3-^P(c5T8JfS3,[;Z4F(WBBP1)NBCF5K#;MCZXEC;^acN^(?TF?J@fCN]_G5e
&<^9_?@Jg::-,C>eA-7:dab:YYP=GcO-2)2c.JV/KRIC/C1#Q+#1BX[R>cgZ>H1U
B65#6+7RB?[:J]5;NJ-b2,eA(?-MM_Z-dR/#9E8GU+:<P#M@#=3P[P/,3<dU_CPZ
&#N]K1:M[\5,g/d8Ab+N\Y]S[)UKT+f+Q:#B1FM_<Hf,3BS#G\>_ea,2d@<ceA#Y
DcTQA2,cB>BaT#>4cW#_SEH/=55^4LHZ58FNP;1\]:4#VF4Q:WR@LQMA+UE57OV/
J7MV/V:\beW]^6]Zf.SDY-3D?Q>W8<JS^d:e=PEMN+fQS9X0G>CR?Je>-R8T^Pc/
@R8/?FLS/;^E2TabLg&b=Ffg?ab?eD9TEVYDMQQ.WRf8T3F@71[a;e#JO#96:Je+
+A]O#N-,U_)QD7ObgCJfc,]e#ZPLE)49YEB)1gZ-SWR&e5B/QRdfZVef^/S+V0N&
:SOL7Dg0IaGE7bN,FQT4a(&8HIfLE.B3-)1=CfU+^dT:cf29FB-2@.O?<)Z8bg\(
0IKX7-L\=gO:[Y(gOTE9<D,ADcPN>e<#9=aEXPS1[E]8HKN.JDD[S9#=1MQYCVVX
HMV.HD2DK8T.e/EI0598EELT_^J\)S@(gJ#FM<XZS6dN&VR\NJ;?Ug#W<0Na5,GW
RY:4b?.?\1VC7>V.:OB\47\ZC:Cb3DeeVCRgI\LGK3MaS8SC)9CA2b\4]DY3U[:F
M&N5L)dDKF:a@K=#V_ENbE0&63ebba1f3H9P7<?H&G;T9<+P]FZ&LAS-87:ICR+7
]Z\>W<Z9/GDHDX7TbB9),ZZSMYG\.ISCMOTg27:8/ff]82.)@W&;Q2@?//cNNT@;
RQcPdN19c\L3;TDF1C/Qb.d_\@;]K64SB/\9L:f28J^-<S@J#WLUYAY^&71]=2;)
6Ic_68ZF]]-8=8TV1P?Va2#eHMEXK?PC8V8]IaOQS+3WFXP^;bddE2//=ED]-8?C
Bg>8HKb?GUg2(\<e-7FO\GYEOe6NSCMgY6;F@C,Ad>A)MNOC3&OH?76d8A40-J)R
V^94U)aY/534D3V,-T\;1FFS]8P_6(;-.=7I>&f9ZbK)<96V#6/+:XMCIK^]A0bG
<]Ec#[S8:d]H/?YEC3AHP>FNH.T]/F&A-FBb)#6]5L0X[]Q,@DVSL>X>U3KLQ@CB
bga.Mf@P@R?Q(E4LFJSR:?=Q,G:.\8+Q;<RcBcdXVQ^48VeB)\(NNX)aRFEfOPfF
8K->P;W3PIf3=AVM4<]9&JZ30g&Y^PKRZDL7bU4EP_E#P76^4^@&GA6EJOLOZEa-
8RGB2b[8L<//S+0g-P6)-V>((L9WFBbR;5=SK=>?fOANW+,>JI7NGKHVEVXJXg>\
)_[VN>Mb]^I/2ZOTN+WLNa<+Le13c?)c+B4b9.MQ8D((D]<U7HS_#CAc^##EB<DQ
:aJWY_^PaHbf/PFTUA&gKYa1ZXM0c0PQO#Vc=U/W5I#&:f;.T^8<?\f]\[-=MH)^
0e>B#fVXg@@OV5c+/Q)WF)2EY;S9RMOb:7YcG.__Y9cLLEab:GNIVF=:Of+^4c-:
N0N+\gRR4?5ZYPR@GJLV0MYCQ7S,65d9C=4:0L/RJ1T.E7H2>,6MPDe[\/^gJ[H7
0GLH571XN&KN7;WF,(&.[H6fYFA,e7PU9HdN2^N7MWgb9)X>R04:Abc<M2)#LLT[
>&.MAA6d:aWOa&G#/)RTCR6&9;>+O)U(+]V#4;Oc6cW&KTTdb0]1a(&[+LSB,<dc
f+?Ab2e=:/IYdJI,/e+MK-:fa@;6/>)U;2&<de<#22G)-A&NbKS0bD><K/>=AA>Z
&8Yb[2,6#74&#F>4&>A.C<Hf27ES1WdQE]?/PM?FLE,SU_W4VW/F,e[.#MbMgXMG
^\Qd+:5/H<2+;EX4QNE-SgI?JBRe)^1#g3^9cVXD(O507L6/0D?eAZ]bUe60W-XS
B3\T7,QJLV]C75)#<1OGDf]8#XE5]e)Maa^Qe5<MY/g)cAD;^E,F.IW3900<.Y)g
WP9Q9B8>)7T06Rg:_=&ZIL0&[MNaf]W_6U=e]NfE&LXdg8LA.8:XV.b4a<)0KD^&
@0_CL91F[-4FJSe0IR7J.0DS^D.Re4D2EG]2Y4R4L0LG8:CW6XG(&LG5XC&EL^5+
<S@()@;M&WD^-:@8.SCH&e;\0CR&b]\@U24E:dAcN3/84(V?GG3)3Z8#aM8gUa0f
(SCH7QM4\aKI\g0BP#C#LKL8SWTHF2L5Q^9IT^e1?dT6WfIeZ]4)1X;7Ygf95)33
EXM@OB:D9A\6a?EAbR_M;--bfZ3d83:JaKIX,TTPef@.>60I[WgcL()\O8cTVGg-
04Ka?1:PWYDXQZbT^^,#&ML6+/Zc(64XNf\a::5a.J7NP)^V@4OSICcLO^WEJJ1-
A47g)#.55A]5)P>-[>-gWB/_)>Z;HSOE390^(AcK:9[Qc[/aHT3O2D3L#][BY6-d
/E6_LG9;9@?LKC+P.?8eZ=<1W(4]5X7EMZN[&>Z?^JafO5+@)5G(Hg2.(D0[eKL/
J<9.B\&KX;M036<\V]LO/=\WV,@E^GP@A1(Z[=GHP,D;E^QW5(,6OV:LLJPZV_J8
A>(C4X9>&[46#gY/1cd?M^C=>0c4b&_QQQOQ=_6GO5CR^1WF#FePdF2#4MVJC8N3
O)Y0?5,JI63VGT_X)TG1XS00J_9Dd5dM\_[T6B;_4(@<0Xb?_X45ec8HVOSKOD-=
>0A1SLZD;P96R]@WOg7L\Vd.3LHg/&JX[F5K<N<CI,2L@cg(^^.84;_2.^LI@_U,
,\aXVQ]#_5ZQPIf=FOV8FP&#HGU86Q>e)(IT:\1;?TX,MS2^;0&^PC)/2T(I,IH\
^fa=IcE3>)75KVKJ4D3TcY5VWdFP)eZU]CSW0KPcJDRHI>E&XH-QN+CZ+&UQ)?g-
CJ@@_)@a=2TJCgR09VAERa_(AA=Z<@,1BVQ9(dQ8\0>PaTT;O4+[,K#X(/28(8<S
H(J1&:LRa5CU-&a<0+JSNeN_3;>gJ7aZXA1VQeH8O?)1XY(2g6I_)R)H0/3LVF?V
AC5Z@W18.dA_H2R[/F@Y?Q9O>c.I<Q>F)7HL6/4VH:,?#bfb6bO24KF?QD6[C6D[
X9P@QYP[TdEgXSL)@@6;IYCgaTaX@7^N5Q5H8TdN[&,08,,KZPWE(-9>a3HNcGBR
C1:TLS[0N6P8XE[39Y8R513HKIJVHc(-BN@47TTM1758YB(;DH7fK?OQN0U((AfH
Vbgc\07&S?bJ.OYUS5XWKVL,-X)f?2E7B+1<9BM_JY3fXY75#H7XC0B]KVK#_Z-_
.X;B(dFD-9A.-73VMMTG7&,426d:,5=O.5C73B;bICMQDRON:EHba2+EaO-D8e8T
CJ#O>TS9A\5(Xa.4C)5]17HAD&@@-\HadAg3\,,HP<Z9;34H4Y,-/M&<9b8SFOe:
O]FT2]dF?cf@M(.Y6^C0FA>-XaX_O[+^Gea4UK-,aS3HT)7A+VYH@6TR9KfgD]UW
Xc2SG,HgEVLBM?\^_F:6Df@&(UIV>:>gA_\.6QM@-+.cO3BM[6.T\;3I39>NF5Lg
fg9IA1cW93O5)R0[5R>RG?:<>ZM>JA25:\K0O4Oc?Sd@,FSc8\c@H#/1DN+ACGL&
IRNF59L^,755=Sb-Z,bZ6dA[4]d@dB&;W,;,f;c0Od_-<IdW.XJ(GgT&2M)PRL<F
>5CGB@[:TC,\&fA7c^g&TbcB^#BU9_4L^-#X;/UaFRb80]^LA8RJBHL7M?#<ZCB)
-0_-I1<VL=5-YQ/88,2b(>Q:f3c#1F__@^Q#:=T9T>-AReL5aC?B\HfM.?Gf&I/L
6&\@VE?8OR6Rg2+aIeJ[6f_cVD+&A&M_4J.6&E[KGS237_AYFA1#TL#b@agG+=W5
SWb3GgC7+\)^L#=NUC=ePASJM7/Fc]HHEGa9g]aF[MD(=4;TCJ@6HSS[XbU8W/.L
SKGf?a;L^e9?0FI?Cd1>I]K;G@A_PX7UePT\U8GLbXZ-P:Q6K\_BYW,NLLOUENP#
[L(&UJ6#2K&/-;[#,:#(NN8^\N_I(f[X\@06PMB&#V1Z7A.LbeX&,&;V/e#^#a^@
W1Jf;_(f-ZH=0d8F&3]Z88(>d-7NT_WCPCI2fCMefMWC;d0M\eXIQWae4b[We+A0
S@+(T2a&c>6)1fVe,g3[@X\JaI=KK,82F\5JHDf0W1K?FUJ+L.O4@[6(@7+E<N>?
=9WN^XRbW+EV21<]39H;:];M^Y7[6JNM^^,XX5;]gU<0;?\GXee^4Zd2gPCB[4;P
=LSZ>OFb:L:ZHb#4Gf#e]^Jc]P,HHPbN4P#C9gT>5,/+[gDEE(&>+YD)M.J+8R;V
J<SDD752#\V=V4/VQ.6=9-V8=DTN8@-V.[e&^fUHa5;-?(T@A-T#7,J^4\S<WD>V
b0P>^Q@1d_SS@I>bfD2ZPQE?\@edK?BA@@IC>UJRedd_bVT6@>9BRB^d<FYU-^&4
5=)5CFgHS1R7(Cd<C&.>Nc[KF[+#=0W?/YMgLYY3#.A4g#CW88GcP95b).g<T[O&
BNC_R75/(L+dFY?FSA6deP,dH(1]LD6,:Q5UJP?9Fa<:bZ1MENE^FTD87T-4/WcS
H>b.^\0).3_J?&3E]/R3F<P^7DK2bW]G,-gH-+@@Xf9\Ja;.AN(_XKJ^8_.d+M4<
-_^5UH18K,:6(SIN)-DR[469f8:GRcS-<U^>QVW#^<E5b0]ZaYRa?DPUbOX9OGLF
HZ8/?cgK)>TJ@?T9^L?O\?DY[@[\=_O&-;DI1FKX>X9C-WbQ\c0W:Q#[N^\<:])5
>.;JVJS+[=S<N=b&cV:K94Fc2&>OaY;SOG>6N5EJMg<e>,E62/SJ=YU&VD3P.bV2
d+0R1g)Y#QdQ_EdW<4)+L1a7)#Y<A+/f?)-<^>WGDWM,K&;YW0;P3#70@=^9fT5/
;3N)R>X=JD9P=W:#M-B&fZR/[D/aag[Y7W+faQPc23-<cHWTOS;:]V?3.?EV76F:
\bG8#1<=aU8@PXf]:@#P@GWD3N)99-;-_;2Td/A^RHGaIXW[@>+II^(T4/OCV+5U
b0^RB5cW=(037&UM/0FD[LPT3M+3[NL3BJF:P,,6XIEC@9>V1#9]H+,;Gdf5)MBS
#>68N[gWYaa>X/]RJ1^\-].;6&G4TV,g>EPTA4B+gSD86&Y^_AHXNI/Y?LIZZY,c
@d#6LEU[3I^NYY(OORf&3W272^1>g5(f5-2LVc+cM649fdX.d9+8@NWN_[08EWaW
Qa_^@H)IfY&P=Z&NQ#GU/?:?](W=bb&fQCEFMSKX^+MP6D[<D.^;&Q7#gU&;;;Xg
La8ZVT7:JG9O56>9,R9_7Z.4<5SL(6BTV@e#&EA:FU^,N6_d8<aIWC&Fc&c_1[Ob
RI>V6.&^OH):D>+RNW^]]@HUR\5@F=B3F)?A)M@b:LY&.c\;\>37<1-[O(:AFOeT
4:HC2fRf&WWc2P4fF(&H1c)cdR0a-.aOGR6=(E5=1&J<N;WRJO?F5cC_RYKU.Q&F
gZ&):<4..0&1@G-.4A\GJY+IXT;:?A<;Ka1Q>;[T7JTf:.3_UG:9@a9JMBd\8V7^
VR[GbfaW9U[54-O:cRE3#Ze=+g?#5C5QC5a:)RWC0Ef8.@<_cge7=f5TY>]AJQT9
=U1P[PKTf&=Aac=g?&-1A@WZ@gP8>HN_P1V6)^<>=]T<PD:;C]^&[U/J^JfV0CZX
M\TbQJe8aAfLB81gPJ)/4L@JYJ6&Xa<0-535fU=fIBY\aN=++bPBdYMU&XFYe<MS
EZfA1]@?YLQ7CN9\HP,VT:?#gPOY6@^6cMGH),]EV^J]7RWdW:FVEVf,@LB-CY-g
#88XPP(ZC3F2\[:,7a^a5&5DF]D\,G@V@GeO&c)MTZ:LC5XSD3TW=\Z(E)\FB+R7
?0a>;2AXM_&6W.^EFW8H=>:YP.7KQ?^-YLL#=\15VIe7N=<:R5RFMS\#YBaNEc(e
6N(dZ\6@DXZ.>1A=<aO+G(YbAFXSFE_HC1(bVcW3.Xb9)R1RFHf#gIXEEZPHKYSM
aU7Q8N@a[cHVL9W7OaD0,3]A5[_-N7Y=_7DfRTMH.8?38dcKL.f]fCR6:O\(2f.T
H((T0Ze+O3C:=bQ-fNN5[^TK34aZNQE.FE5.4f\JHbTGRQP.J;4A(Tf;&&XLMJW_
#/7(HDQ;[@O8C/6X+56RGOBQIW(e+V#bQL5EV(5HF,c;NMB=VO/a9a]^ZU_XZHO5
(Fb.aMV@PQN7(G;Fa73MbCVVLL8P?JC^=;U_dE2,USLLe,B&([Kf,]\:K5DLSdea
-??CSBMAXHcfR=16^\&XS0)ZP9AV>;6^IWb(^VI\01>SK(PG6T9a?ZE0Kg7)]OYF
#FIDJ3C>9SUB=+0S?Q)5EHDRX\fA,g;0NWKCO#+1EM.XYWa\._[b#3bXV8)HJ&HM
0SX0AbA8D]TEHEGe/GS5RVH9;Z2T:E#:QHOda4^eB2O168C-8PZN<P6e+LZ<Y;LP
C7/(X+8X,aB&9T/C4D=.Cb</S3&Q)FYUGEgJ3dA_>fLR=84LH<3d?Z>HgIa?515=
ga3f;&J[MU7B\c,&ZF6Jd#f-Y_.=;Z4<^&S:49I]-01ON-+)64<A:[be,f?Z17(<
bIC1,IE.S3LGIDa48=SJ]g)g,:U0S#E#-+BC,]WPOM]2683.<M0H]JT)a)8?fMU_
?+#JQbV,1^Bbf.XI:ge3IKD>#>68<d:PTf8:QD)+50Ud]R:b2H08?P+_LJO<N(47
BcbYYe]V7GR^aIN9C5@I/CaeYIgZX5PfQE^:2e.cVaZ\27C_.TfRXaYe)cC#:I&3
N_4[e@#af7.DXJ&/U[XIDg,N)8/>V[@.c3d42_,R8BJFbM02?Q)OOaMBY6T+\3O#
B=0_Jg,aVQdL7H^5N)5CcN5[I,T1..;gb[H[T;M5aQ3<^;/[,W_-QI<XJ[+/W@]Z
NB)\?YQYS(&J&-O(.3\7HPQEHPSOOO=[I(@YW[#>9=WIg>00C,74bW#RIWf-8LZ6
CU1bY<@,Fc@V#.15=ST)d@\(&2P>LG#V895>86TS;A@NS5<)cJQd37+.\W/&X#58
2R:+^V2-=E1O9+fJ/5BPC;+R^KN::cI^6>1aAX.A:Bf=Ic8WX/UFaA&9_HHQTJSg
IT?9T2OgBdKa+EcTb2J<d#XS5KXP_&ME>\7g42dbb3)([>BU.1X_TReS4=(0KN6_
4=Nc/J3R52^J/.)+6QHB&YC2-#:S66]K]MPPPg;TV#I5^V:^C8OQT/;(Ba,c;@Q-
^<4@,d:c@Y/?/2E/(cE6D^E]Q>R4ZT5@CD/B^L\+/LFd:@dIK3-#?dZ>bb;4_8IO
L&^+K?G:FVd#JXRB9)S,<6HdE98O5]X^4,;AL:#I0Pb99-bCN)g@<9ZR83T+Z6.<
:J/DJMGQd<eDbX.R1Lad4EJDUZD17&XZ4Wf^]cDOX9QADRY\H][UgX_9R-_WVTH0
2:D3#gULSXb2eVT),)VNUUS=05GJgfg4U2T/<=_dI=SUBPFASc3)RfDaRXaW./G(
NP[ZNYR7]);[8XeJ_aKNdF9NX]\C:,g\+X_FC(T@5;7M<1LdFC^@C18#F-;+DDXF
GPV+7G:RH<,\I/Y,]DKLL,?eDY\RdRU3,A74.R2K&ac\&N:FbY@VW(?_/>Q/97Ue
6ECPXW7+3bg>&+2/H7Q=F^O:OLd>Ba-.@)XW99/<JY];-B(PH-H8?YTdRSSNPO\O
0b+F/.^G(ZO&TK2dH@A]&OGJR.?c^C:ad&f&S(-YV;N[1<cP1eIgS@V+YZNaT@>[
JZMJ=ee&2T;bb[W>Bc5AT=UFI\d+gMIH.<.&MTDJK?,X06W_DfAYYILg_09?Xe(c
H.a@cWOVW_5bQBKP0;)PW&D7g@XLVLIKO&9GYD>#).14#62#H:ZaBUaUAL<JP(_R
LM=e72fRMMJN7>DeY^Pf>ZZB#,YJ6J5TL,?cf][aJF5V^S9AUWL,<dWL_.7dL\<c
Ke>M4?=GB.;ZY&;235Vc::V0g(U)JFd4aIKg,edN?<gN^^5^I;:&^-L[[P,Jb_#D
(NH6J8/[e]<#ZRLJ^4X0PF+2#TL@6Z&a2),BReFR(:G_+K23/JT[4cIPYUaeC6VY
PZT8WHU5bTI/6]KgSI#GJ3bF0WFP\YA01L?/3(^<LF:VD]AO6f-]3#8?d>10Qc<&
G_T(?J&/MQcXGR.@.5_M(2Y0Ba4f>ec\V@?].;XKaeN/G)KR6<C/#/d-RRQQ12Jd
E#NaPdV+3KHXJ?BV.)>MJge4HaPOSF.YMNbMR+\23:[d[51,EgR&T)#ZE=#_gW:S
.XVGPX9<E-@8F,P-V8=ZWM2=gEMD6-:7)BWO,PG\@+S=f,AT&..:DbE9>+CH0PK:
faV-(V<3VCa_/0)IPI(#\EI3L1d5P;86XS<\7L3E9XS,?,g+:V2OLc>[PIP5KC/C
@Z(\:g^D5)^>LJZO0NIT8c;W8HOf\NGTI;a?OdbW>:<UaSf]YM7H=2]DLGO+]dI3
cMO:QBPGRQSCG3/+^M?-E6TX::[,g=gOPd4^PGJP92##<X#J),JQ[K/<ggRYYa]C
#B&?2CJ@IH4B3N(R2b,U<)4)&RIPc<O#;=:3P2I;BX.g@^U3PQ+cSfT7AWCC^-^H
aJP1+f9?9BSH>_6gY^g(7OcDOEH8R>BV=eT6d9;gGB78N4CBQ)KGYG<g>41\9CbC
G2\>0d<)?<&4#;LA(YO2KH4Y2=RfQ8IRJD9YH/GEO],)J=SWPg5R@8YeTfJX0.79
T=?3S\U_B+@f&cW23(?R,4W)b7g/Ya5X<]_<QOIRdW3WfQ\JE25EH@E#Y2#Q)/e6
g.;)#&H(4@>e4B<DdT@#0W2>1)Ab:L_aPA8Ie4ZWL+0C#\6XLU?:)LTS48_+J/]<
Lf0(^5YRa[aQ2[ZI5NEfS(40V<AeH,8;7-M^DT?d3cOX&_)&?E=ZC<bM@9,A-P-?
\FX(_;A&=cPRcQ?LLD_]5b#3c1eJ3\NbOCUd+>:MMDJaUK_@Q975[V>^?bNIS6SA
e:<+ZMYW:Y&,N(87_@URU<A>>(Ye6K5Q]VI>SLcM<Q@T,3Y.W7]P)I#aB2.GgXWI
#3JQ#=8aX]?g#ZaTdD6F&bPSdUYF)WQ;gK2\PB^[&DUG8Dg#)RbWZBU4e8bZ()^g
XC2,E;7^647_VXe&/bBY<G>90XYEI,(gM,61<O^b>Jg),KQ@+-RB)ed#fZ<YB_P_
[I)cX]a.J7R)Xe?gOCA@KY9+b767UG)XF.dLPg]fOGKK_4SR(8?bIDQYb(&e-c)=
EdNRK]e\Jbb\d7L]AXC^NK/0B;]cO0,9JHAEf7@E,^4U8_C]>>+K4-5cD0MK?fG&
d]D0H5U)9VcIdG38M=_ZBJO^6QR2\EWF@6:Q-MC-/6]VUA#;V7&/O03g_QZ0;2A3
@ed2\f@aN4Db[5ACQV8F8D2I3+OQbf9?=5KR\1<X0;6O>C3[OMFa(^^S7B-NHg2c
-9JKf[+_APLS4R[:PMY+&B[FM^9e#PC9(Q]:#DKE&R.(Y0&CeJL81+A;;6K[1Z^?
RLIIZ<[UJL(O#HA)&+2ebbRAf#TF<9Aa.c>f7O/bKU22-U5;)6G&C,LaG3SHc^U(
2G+61&?M<3R^N9=V,RGDM50ZCK[g;.IRV]Q6R9<,ED0696E)3U156R_9-;#=>R.-
a=?6;Y;3\<#S#A3N5CMfI<BX<_RWQQe=3QJCdJ>K88<U7_6WGO[(-SN^bG+D-/[_
<65f9L^Mb6YJc:-R?LM[^UTCJNeYT(.O\f52YL)3I;GN:2(^<(MGZa+dRJV-[J.E
D<;K[5#d6)fIP(>H+_@N+M7QCgZ]+Q)V,]S+<OPTdRV:(B5#M\D,M35]G5LQFT?>
F--03@UPWSOF34+1CI60TRGcC0P=QFOd307eZVX9I3BI254JaQ.cY(4,eMV/9UAd
7A6.,gA5;H6\\GK)YT9:_)IeDbS^S3:GG@H6=c_MV)K0#F<FG498-Ob#^VI&TB#9
OSL<PK1/e)XXK<;F<?.I)eC_1fX:UAULBcBFJ>C.cY3WPIe8;T-CGM.9K?5b8^F5
1][,g>f/aZW0B8R#::0:,FZ&>+YW0[TP=dT[V,_f@3,9fB)_cS>ZL;WCS&THgb5-
,J><BA<)2XBV\gVUUVLb>VT68F;#d[>eVX@d/98ZbYQbAF&9dLP3\?)?SMF:Q<6R
/(ZF:dcH41[?.+CASHGT]U>QVAJNG->]NXA&K5eT:c_XU2gEfGRV?8Y@>)-P-G/>
VOR:?ZOeS;(V#FHARV4Zg;dL@1d7RW;H\e>3EL,cbA:H<5C__36Y=:5eGLYCZV\U
PA2##M?9Wd?Z;6e>2D18;U)WR1Q6RgA5U&=@gIgZ5.(2^FM=,K4\Ng2:bK1X:a^:
VFcJXLN]#+MZ\U;V:aG2WS^9ffFC<D5^-a;dNHP&Q=8a<M<LdBF1&/I_MbKKEWSB
>1IF\7I/U-:+029NE7[(:Se?6SU]=/)#19I)<=6?dA2c><MCQ\3c2480P17<E#g<
,>/Ce(cWCIUXKTP\(D2:)D>4/.KZ2+((,GI-g)UHP<fac]\-J>>7S6W))_KF&W^.
<]Ba[##UO=@K2,;HJ^SQHC3;PT7UI<@DdNEWR(&Y>[(XI=CP.5#VEW--ffgDVKS+
G?&F2E[b.d5+39>8Vf-WV8gfZfS>?f/2)?741g0(IS-8-9[?<4a:N9XfH64Z1L5W
23D[^aT1X\?EM-+QNa&E=6Q+N6M/X7=QHE>Z[8+EM\F1M/-T#aYPc2La_W_VB[2E
F@aAeZgR24E]8I@5_geO,</=J<(F4Ed\KKZ4TR]\ZO3<1d2_#XHLFfA5=Md<a3FJ
7O[4MMV3BF].3/4agFLLcTa7(??=NCY[@]J+RQe(&^HN(a89,=fe^&f-bAdc[ZDJ
K7(A60=Y?Ae0+K_H:_MCG27d4F1,P9MSdLUY@HR[-&cZIK?C@D=O(d30Uc.P=Kf4
F6/eOEODT(=c)AN:Tg@EKG7[_d#a6YFS8P^5Q#5:5)>3.HC@XNF^7a>2ZX)T3W/)
:=3W.CaZ5MQ?C_LCWOc=WM.d8?4X=B)5_()PI+D75^S&YTG]#Wc^DB,5EZ^R+PX)
YDeaceKgS1]ANYCVUGJL#=AO/M@OW)/KC4K14c@(_[;bV?bWeBE2U(#,G,/NZ0W=
<Cea0XKUF,FX/ac/>OAQ&P,14.R==MK1;8Q1W3<3g#aHY9]:eH<\83(eDY)148d>
LPTf],I1(fda@R8RcFd&XUg9=&1&(Y_/>EC\D\O&B=4X83YNFPRM>N6F\e=_2,RT
:I<c\E86L?fXBReNC=NS1]OSgF<.:5eNGV;e&I6D?>&f>4YVXP@(74I+?[Hb@7E3
K-2X^c.&(SYX5(>/GO\O?],2[Mb1(;OW7/1?E1B#dTJ0cX^@5Q_L7KJMA^beK^TQ
:B8OIO0)+J-CM/7fXJ7O#eMMM_@2)11/5(-T5U]G9L.Ia?_Wa2-c\TeJ6H2KN1.C
#=S0FF.Z658Q.I^J@,1SFXKU(0.b<K<+C,^HWTd@;-[+dCdET#9.F(C(L8=>7W1a
<9)J43Z)ML)JAF;,O;&1F6R>D=0WE1-g)B4bYXQS9(@PbT^W^+E3PXDNK-3X\>A2
0^YTb=VD)AZ5EJUSP>=+T>B:gBLW.b#[L1dc4U#_A8R.VEQ?L/Y[d](:(Hg=^O-8
#EV76G^KW0?d#D<e_:)F\2I7WS+M:C&PXSRAZ5)W9:MVXAd^W+,@OF)I#_/L-Q8R
:?]PJZ-DLY/+<HETE,[X#8\8N_>&TbY?IJ7[>>_.2BQFY8aA+aBN>6YN5\Q:d([,
6]a4^[SNU970(/8@0)[T9SfL>(1Y4/P:E=TU/DCc,X&JNge_XQ_UWSc6(>e]A7RQ
EQ1Wa?(@PQO=9M)KLBAW2H7=^8B[WL)U^UKgUA[S.VS+-N&C<V8_MNF/XYR7e:-X
ZAaG/dS8Je>,@[/bG+3N3=_FCA9_;=G=)(B99J2TWK6dS?NcBYL;d04]MKXI-:[Y
f#3/#M9)_cTAFf1L:I_M?c6_7#<DN+P\AX<&R4/8\TR;[1):E;<]&@&],:=W..dg
#CO1QJ2&J4EF;-Y4;P/TLH-H,:0#P&Y0g&4fA[QfB\f/4)bB#P:NO@+&6D4PPT,G
7<.1X<03DT@g4M=dNJH[d#Uea)-C0AfWBU4FF[[(e+?M:S?W[CNdBdQ9Q8(8[.XL
E(]81bRX1aDZ-M3>cLTD9A@YDK>64P[4D=,L?E^-UC@Te:L:-<F>)^GE8GK=-2]/
#FW)M8Q@X^T3g([9b?ea\O4-6eObC\acK>@S.K#+]H+]c09C7fZN-VP]DMUd\-2:
UI9baPIfC7C8O>-._gaOFM.4,C/B,OE(c1G1b4cg>Igf2g/X.0O#>=T1-9,3>YFZ
Ma=SObcb;:f\&d(2)e6;FcD0.AX=A+G0JPKN)#J:8]<]UVCAUS/C@fe:R@b)]U-M
#?:]1<FQBe<6]W6Ka/G98O_=OWd/L7^\YN]cN_(P-B[^4#JX:G_;I3,XR>BI()MB
g3@ag=8L?R&95F/7=4E.,LF>RRD9:+]H;d#MgWNN]S2DDGa7\L.4ZZ)QeCSEW\<R
)<;DNZ@e#9H4KO_Z_#E37YPPG[FO#88]&]TC<f=YWC&Q@W4<88SY3.?#]J^@A06D
,B)D#;3)&=2gPcbB44.Z8,:JA2-U3G-[)KeK?_V3X.C\>L_M9)Z[HMK>9^C@/;;Z
KI?eLJC,e_7(?#HZBfDL/CX.5/SRADD4XKD0BI(PGPcUW(4RVQ:P?eO:,+c)?JM7
aY(X9dI1DN2</VQM:UPY\K?;3cD32NE_(K]:/_COZW(77;;DNcWS#[5de(]&QdaR
?df6FCXRZcG3\gP]/:K3YA)9f5T&V/&&+:ebM9f?DV=@M)Z=OA?\:NC^a\+3:61/
eVN.MYC_342P_VFDK0a#&.G);b<5CFZ3.8;\CQHUPL,e?^;I_Ob7T^KG=9KE0ALD
F6I)D3ac4QLH\>1DQ;&XKD,(2aPeI)3edRL+-?0E(cMD>=48IA\JW<K&/\:H:K+L
eFLI:3H,_T9SCF#\CEIH;dfc&U?-1A\^?ePAP7IZPRJH,cC=4(_\U62G(;PO=A#f
E4BJ<cDO&a4@4KXe+UNGIU/HRHcd^?e..Gc-Vg>-QCB)ZdYEE\dHDGOB+C4/8XP2
E7@DQ]X6970OY=1S5S5&J#I4V/f=2Af)>\JPG]3MVQIA)1</WUT1]7UWJN)8HdBL
KTaKb_V=/9==?V<6J:\E8Za_92F.4ee83Q4Q0@c\P5^f4XaYWN@+Y4;=7XKcb>_1
[CX&15T-=9G5;J&X8^4Yc>6K[3a=^Z0T)#0>>IRZPcC4Nf]JBg1[L]d5PGTT(,f=
U0PgJB-AG;X@VN1<W;<,\/IMP0H)=Y;ZS5]PbcT(#S-aWN.VPW^H,]d5I$
`endprotected

endclass

`protected
Q8XDfd>.1+8Z\)L7L>e?41T\DTKa1L-PG/HYNNg6C:CbOAZ#?CgE+)9OSVOKa-X8
CdJ+[JEK#aWWW-]]V<4/FDTf,>&a44EMMAWRT-_<[+e@K0H;<T(gW>Ha+.WI]:a^
O7d4>cHEU7;^^fSaUKZ(+YG(JB[Q413EB((FN0f.?3K^d/#\;DH(d]3V>baK?8>A
8]E9bP+:IV]X^+XVU^VIUE]B;MD,X#YVa^OTPRM<QLRY2Ye^XNgG,7<F]^bX-g6g
).MFSL?JeLF8?g^6?dZV_:9=eY@Q?BcQPE_cI[<U6FLVQf4e]W?8a09LcT<f-8ec
2D2bVCTJ==Z9bWV8=e<UC/&R^)Lg^?TZ]JgRU_OE_9beROaDb=JE(#VTAN,Q&4]H
2I>ADgUBaU\cEWBEE1WL4E-^\7gc6+1#0N:(SSU4X65(K4>7Aga<^/B:L0)E:T>(
#\-)ZN26dLGX4[HL7>Y>ZTW^;-b3gT6>)6fO4DGRbXCe=[P)d5W&:5PT/H9gZ8KK
4B,]Q/8Pg0)IO(BDOUVEIKN5eU]f.G_:S>agQA[=F?4?#b]U(eIR)Td<fQfW3@cKV$
`endprotected


`endif // GUARD_SVT_AXI_SYSTEM_MONITOR_CALLBACK_UVM_SV
