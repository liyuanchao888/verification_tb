
`ifndef GUARD_SVT_AHB_MASTER_ACTIVE_COMMON_SV
`define GUARD_SVT_AHB_MASTER_ACTIVE_COMMON_SV


typedef class svt_ahb_master;

/** @cond PRIVATE */
// Note:
// This macro makes sure that hwdata is not driven beyond cfg.data_width.
`define SVT_AHB_MASTER_ACTIVE_COMMON_WIDTH_BASED_HWDATA_ASSIGN(width) \
  width: begin \
    driver_mp.ahb_master_cb.hwdata[`SVT_AHB_COMMON_SHRINK_WIDTH_FOR_MAX(width)-1:0] <= beat_data[`SVT_AHB_COMMON_SHRINK_WIDTH_FOR_MAX(width)-1:0]; \
  end  

/**
 * Defines the AHB master active common code
 */
class svt_ahb_master_active_common#(type DRIVER_MP = virtual svt_ahb_master_if.svt_ahb_master_modport,
                                    type MONITOR_MP = virtual svt_ahb_master_if.svt_ahb_monitor_modport,
                                    type DEBUG_MP = virtual svt_ahb_master_if.svt_ahb_debug_modport)
  extends svt_ahb_master_common#(MONITOR_MP, DEBUG_MP);

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Virtual interface to use */
  typedef virtual svt_ahb_master_if.svt_ahb_master_async_modport AHB_MASTER_IF_ASYNC_MP;
  protected AHB_MASTER_IF_ASYNC_MP ahb_master_async_mp;

  /** Driver VIP modport */
  protected DRIVER_MP driver_mp;

  /** Flag used for handshaking between phases */
  protected bit drive_data_phase_active = 0;
  
`ifdef SVT_UVM_TECHNOLOGY
 /** Handle to the UVM Master driver */
`else
 /** Handle to the VMM Master transactor */
`endif
  protected svt_ahb_master driver;

  /**
   * Flag indicating status of tracking transaction.
   */
  protected bit has_active_data_phase_xact = 0;

  /**
   * Flag indicating if we have a preempted transaction in process.
   */
  protected bit has_preempted_xact = 0;

  /**
   * Flag indicating if IDLE_XACT is becoming preempted_xact due to
   * SPLIT/RETRY received for previous transaction.
   */
  protected bit is_idle_xact_preempted_xact = 0;

  /**
   * Handle to preempted transaction in address phase.
   * This is required as the preempted_xact is local to drive_address_phase
   * method.
   * This is needed to especially invoke start_transaction() for preempted 
   * transaction when the address phase of current single beat transaction starts.
   */
  protected svt_ahb_master_transaction global_preempted_xact;

  /**
   * Handle to preempted transaction in wait_for_bus_ownership() method.
   * This is required as the preempted_xact is local to drive_address_phase
   * method.
   * This is needed to hold the transaction of second INCR which starts at
   * WRAP boundary if the last beat of first INCR receives a Non-OKAY
   * response.
   */
  protected svt_ahb_master_transaction wait_for_grant_preempted_xact;  

  /**
   * Flag indicating if a rebuild is waiting for address phase.
   */
  protected bit has_rebuild = 0;
  
  /**
   * Stores the wrap boundary in case a rebuild is required on a WRAP type
   * transaction.
   */
  protected bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] wrap_boundary = 0;
  
  /**
   * Event signaling when the address phasde of a rebuild transaction completes.
   */
  protected event rebuild_addr_done;
  
  /**
   * Event signaling completion of transaction.
   */
  protected event data_transmission_complete;

  /** Event that indicates that its time to fetch next transaction during locked transfer. */
  event           fetch_next_xact;

  /** Event that unblocks nulling of global_preempted_xact after sampling is done in case 
   * rebuild happens with SINGLE burst type. */
  event           sampled_global_preempted_xact;  

  /** Semaphore to control access to driving hbusreq */
  protected semaphore hbusreq_update_sema;

  /** Assertion time of hbusreq */
  protected realtime hbusreq_assertion_time;

  /** Track if this is first drive to hbusreq */
  protected bit      is_first_drive_to_hbusreq_complete;

  /** Track if first assertion of hbusreq is done */
  protected bit      is_first_assertion_of_hbusreq_complete;

  /** Handle to next_req set from driver. */
  svt_ahb_master_transaction next_xact;

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
   extern function new (svt_ahb_master_configuration cfg, svt_ahb_master xactor);
`else
  /**
   * CONSTRUCTOR: Create a new common class instance
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   *
   * @param reporter UVM report object used for messaging
   */
   extern function new (svt_ahb_master_configuration cfg, `SVT_XVM(report_object) reporter, svt_ahb_master driver);
`endif


  // ****************************************************************************
  // Configuration Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /** Initializes signals to default values */
  extern virtual task async_init_signals();
  
  // ---------------------------------------------------------------------------
  /** Initializes signals to default values */
  extern virtual task initialize_signals();

  //---------------------------------------------------------------------------
  /** Drives hwdata during busy based on the configuration parameter
   * data_busy_value */
  extern virtual task drive_hwdata_during_busy();

  // ---------------------------------------------------------------------------
  /** Update flags and drive initial signal values when reset is detected */
  extern virtual task update_on_reset();

  // ---------------------------------------------------------------------------
  /** Accepts an incoming transaction for processing. */
  extern virtual task drive_xact(svt_ahb_master_transaction xact, bit invoke_start_transaction = `SVT_AHB_MASTER_INVOKE_START_TRANSACTION);

  // ---------------------------------------------------------------------------
  /** Internal method that accepts an incoming transaction for processing. */
  extern virtual task drive_xact_internal(svt_ahb_master_transaction xact, bit rebuild, bit invoke_start_transaction = `SVT_AHB_MASTER_INVOKE_START_TRANSACTION);

  /**
   * The methods asserts bus request and lock if enabled. 
   */
  extern virtual task start_transaction(svt_ahb_master_transaction xact);

  /**
   * The methods blocks until the arbiter grants this master the bus
   * This method is not called in AHB-Lite configuration
   */
  extern virtual task wait_for_bus_ownership(svt_ahb_master_transaction xact);

  //----------------------------------------------------------------------------
  /** 
   * This method is used to check whether transaction will cross the slave address boundary or not.
   * If it crosses the slave address boundary then transaction should be dropped before driving it to on the interface.
   * So this method is called before drive_address_phase method
   */
  extern virtual function void is_slave_boundary_crossed(svt_ahb_master_transaction xact, output bit drop_xact, output bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] min_byte_addr, output bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] max_byte_addr);

  // ---------------------------------------------------------------------------
  /**
   * Drives the address phase for the transaction.  This method will block until
   * the address phase is driven.
   */
  extern virtual task drive_address_phase(svt_ahb_master_transaction xact, bit rebuild, output bit is_aborted);

  // ---------------------------------------------------------------------------
  /**
   * Drives the data phase for the transaction.  This method is executed in a
   * thread and will release the drive_address_phase() method during the penultimate
   * cycle of the data phase.
   */
  extern virtual task drive_data_phase(svt_ahb_master_transaction xact);

`ifndef SVT_VMM_TECHNOLOGY
  /**
   * Transmit response to transaction.
   */
  extern virtual task send_response(svt_ahb_master_transaction xact);
`endif

  /**
   * Executes the steps necessary to complete the transaction:
   *   Completes the driver's seq_item_port handshake
   * 
   * @param xact Transaction which is ended
   * @param xact_rebuild_in_progress 
   */
  extern virtual task complete_transaction(svt_ahb_master_transaction xact, bit xact_rebuild_in_progress = 0);

  /** Drive the default values of the control signals */
  extern task drive_default_control_values();

  /** Drive the default values of the control signals */
  extern task drive_default_data_values();

  /** Drive a beat of data on the hwdata signal */
  extern task drive_write_beat_data(logic [1023:0] beat_data);

  /** Drive the address phase signals */
  extern task drive_address_phase_signals(svt_ahb_master_transaction xact, bit is_drive_along_with_busreq_assertion = 0);

  /** Ensure that the tranaction is valid and that the handle is not already being used */
  extern function void check_transaction_validity(svt_ahb_master_transaction xact);

  /** Drive hbusreq signal */
  extern task drive_hbusreq(logic hbusreq_val, svt_ahb_master_transaction xact = null);

endclass: svt_ahb_master_active_common
/** @endcond */

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ptnSvzNMsCZaKLsiKZXA4bTr3yYN0lT1wxQmkLGd4Iop0Q6mNWCG+ev/K943RNyl
WF9OKPPKH+myicIHksC5CdfSU9cu9IfKpaqw/cZtH/zpUA4P7hA8wfrm0Fl7xEPw
JsVYAvviNmjNLQAZ1b8xIjvn2IcI4MXfRcea/1LWdFQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 586       )
g5OObxO+dwzdFMH+Q7JyFzJ0HwZO51y/a7kqNG8oBnAAWofL0/DL3/bIlD2A2Bdy
90hRi/oTCv/qhxNt8mTX/rJD036kcdu7nFeFKm9o/m9l3sirUaV+natQdg+svQYY
rlCDWV8yGD1dsSaV+btJ+96LnzO4bdO0AGRqVVPzV94XaGxUbSFviSuesMz+mlY2
XOowO034LmO4on+P18N8IPAja0Z435UBPXu30NlHQgn0V0cdj4c4ce08LY9tdceg
BnBwOWupHtC/o6e3K6K6JTOnSjk5BQGLSzzftvIFkv/sNFkEXTSE5uv1GydR2NVU
D7jkRm6rNCreoSsFMMBATiw0fFH5sLKbB+HTkhRFfxjWQMm1UKLD67X155lGjapd
oHX6VTOj4l0YoevR7F6FnwtYrJ36yN8kmBuM+eiWP7kkC2sOk6aEDwSHRGuXU6gb
/lPqVLELPX2Ci+HUZnP6gXI05Bs8nJ8+1dhMsQxvRFWBDN0WiSLwMGqA2ZwV32z7
CRObTxcIyuLjL8vreiYwc9qPBRhEmkQkJX8qLCsS7LvVKHjCwMCuDfBxAAgKRb3x
J+2d0omyhBcc74fy8waJTh8j6ymgko+Hw40GUPsUV8HqbJlBjmbTajj6LlG0WnrU
TsDIeDMbXrTysaFSFRxiiQ430ArrwarsEggdxmDMTVpthtpZK6JwBgl1+QCpObXd
Wjt1TU6Y2O0mcP9TtjXktnTz8BWX190T8cTDt2svpo0puUWZ8zi7Ch6AVEIbY7v0
/vQ/Y5WwqPrNm+dfhfahUg==
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
fPaUOHWy7ajvJjsAIAksLjKO5Dj9yCUmUggPi3MBqlLaZznNFko+8NXcvjUUphkf
PBJja6qPHmgvX3nqFC/ymt7Vp+cYPFvBn/zss2ncA/kopi5L6bAJOe+5Rr4sPf3g
qOU+EU1IAdBf6+DiicU9aMm4+3Lt/IfCstM29NGkurk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 12208     )
sq3CtsHPFj5Z0IepYwHauaAHrKel4nnqt/ZVGRaxI/i5/wn4cixR1oYNx1kA41NI
005dYE9cTyOcr5RIfFcy7tbWZk7jgCT046v306e4tRFVwtZw9fte8vEKLQOjesf5
9oUXcOQBX39F/oKeFDl9RZWcRGoj5iHLVgfgsn90lt9XzhV+vzYB5yw8F1F/kzLT
XQC1Y5vjniaNvUspZi6K3igHCqBpCYMqioV+tk1GFi7cZ4P6j/DCfg4MwBlEJqRp
BAscddjFIV+oB4uPyfErbU2HuCNnUhTs05FaWya/QMKaFOiFzJ0VgpSVs0O5CLh+
VoJtUcDUDNrdE9U/UwhW8t4Oic7Zz+0YeToiu2Lf0ixJgLc2X4d/NPFBtlR6vVxw
qB44jRnduz+jefbmDlZdRNHPj2FaNrj0jvrgVlpFCNKALHrb8tNNb+S3mTG9vksY
eormi54Pqhl3faduMBvUCxiIIsbQXTnRpJ07F67hhOWU5UgUbrdnxsY2LhwC+cgN
UvIubxOgB4Pj9P/2dfjprlvFYPvhwmW34Y0r3Hig1Dn3xUAZgDd9v4gJERRVK0KE
lROVuaqDDCroTwLNaWQDIKf00wFnSpE2xTo/AqT5g37p1NXlmRfhjhYSm2SAepmW
5IKvrZiluzi6D0qvaNA25MyJQk75AOicp/PRmdg4cYUq6mRFI+3sTFcSP21PWDpW
IsC6fncicsZPzJtSkEUy5pe4qa8q9iDdIXu3SNBeTOzIcxZq4j+wKt993SsaPryN
K39pEMkr9r824EUqFiVPRxurDH96VkSj1MAFkC34pLBTeXeYK+xjy0wUnI4yp9xP
3QxnUYB4GNvnksPhmuwxxzD8mXt6JBneJwawx+pdmXhva0mYvqFcaUlWRP77AGE6
9yGyH33qcwhvsGg6Smqz6xKvRoGr2AFKasJQaHMA2gly4sF1rCQhmoGN67Iqw34V
v2X/JFkLgKE8I+Up3X4rDJmJ9VVqGIuChton+ew4WqqqDq52EzWxyH2iOEqguNCE
/iVAIwUa3Mc8ZRwhV+bHSGzQGoPROz4J521hvyF2RTWsKGdVNR2qXQ4HFdnOI6Eg
DlyPENTP0/hvDLbtMNDPue7RoGklTMntzgRh2J3BjW2qpQg0AJQu2uAHJXNtbehX
pGXHKbI7wy7375OSOn7mWK5l0GOqw4chg+V6BX/Aee1DwAvBHGsc5acBzzvQqpaZ
F9SU0vQD/PQ629nkaJaqiO3jpDcAVWyPlWbnatQGTidEKLyWW4nHlST/ZOY69AwT
DjYZgM4fUXgBpePcjk8tZ5bAlRB8JK9umbgwRiFPkyey/NGrl7cM5+8SJnBGWltU
HtrCT6S3KcPjRMrbtB4MNEUBtaZE120yGKLo9TCy6GtOwee4GZBMz1umYMSinP5W
Q3rA9Q4ZgopClRMFoLmowgqyuYXr8aiVm3B0iukkF1QSAIEVisD11RS1CDBID4OR
il7heAl9+XAiCHfXGuNejZCCfmJthHbjp3KvR4F1Va45t+TYI1GIJHhGkREATcOU
4g7FcxukGbTWbHgqCCTuCyBvstua9xZnGQo5ZZ47p/QoWnzvTlClMZNQpd6/n9U4
CkflPAOAEj50Fd73WYRe+Xs6WkhretkG27d/hAGl66C0WM47wA+m7i+p7Y7l0CeB
/ixTeoOychg5Tyr777dv4lDHbUL7nvvrgaoi9KtBo1q1y+1yv84rJ1uAH3ksA7pw
ig6tF45GW8O8FW9NC1c8EarnaaO2MyuZSqEJpyh4bL576HwuiILaOjIOEJNFj7r/
gKz6Rpx75bYMeu09AEu//xUc/2EOpV+EqdCaZ4uFrq7/vfmgpKJwuKOM/unj41+K
TLPVT7kfiDc/PLqRnVwapFOYv9GPZqW8riiPSM7vWMDg69sFsl1t1CXSyAOH5yTp
z+oi/q9SEzyjgNNZbBGI8yWchzC89aOADV5uHDukRj3szFX2iUBcCJDJNVfLAU9J
teLrnqCECS2o0ra7Sm3CuJ9HF6xiBxtG9XtcWvDKprB8uBt1BkRecijfw10jjt9m
6fozUIAwgz8HAaXFBYN7Eb9LRyax3S8zmSqvcC//qHB+sKBnOWYS03mwwioma+Yh
AwDv5OekhLUrLDjlRDyxsGPr1SalgaEdE8bIQqXBU9nNC0qSM6ny6M8IpfNM/Ht9
o4N1semsVrFdwXXsAyifbyeq+txwwFp/Gjx/qaLZZz5ArQQT+SSvdCzliimadjG3
ESEo/JHymubIqBlrneC+pBFXAE9NHn49mv8y0be0tD2sgHYz73ct4sCWu1PMSeiQ
wZLfIuuaLq28Xt6XP0Mc2poZX7H2M9i+1dN23sqBfnPfCPGKQFc40FEAn3dFrojN
Q5npcqK+IF6DGbSVa+5d1GjXMZ+GMgdmaOExW5tNQ9kZuWYFy/qD652WLKTqOnwb
dxzFwkfJ/93r1CWNvbm/Nj8kBxTqj/vyX6JsEKeE69IR3iWA5JsPWMZoC2wTktfb
ajTXCW5YWSfPMI6QMk+U0y6JM0kCanJb9gmfPpuc0x6kR8J65E00ldQW6BSKduSC
1o+wv6IXr7iVX94Y9LWb6YNJ8cb2eMhOs3sM7EWCIOJAnvHWsdtYhL5OZ5+ewGqr
8XPzDvvDYU1SFsAEJU6trqDcJDplsZZrfzhj5Mp0oL0b7kJaERij1LdrWvOjZVzV
jZCIxEB6JwXGJqB9qWqfFeGJgfSmXF7Qvx0LVibdixczIMcu7W9kpIJ1HKUvXNsr
cCD2luiNwnMBBy7p+SwSWrU8VVx+6ouTr50R0jU4mjMHDY8AmBQEtFF2NbTIF2bQ
IaEfFX0h8x95KcDPDV4uYwoHMndSCSf0OlnzBnmMF4aaFjoU+5wB2h1QgPJp+P7D
bN3CqMq1/118DQCc2XFB5rPHEljyb39hIeeux3OkcXp5Ia6P8MrJTLhoT/l5U0AA
zyFQeWkJEXvHJK/jtb61eKo6cglaPwGXAoFSieURV1gyuotjxgawijZAZJqmLnm+
2AgLwctdJPnxcydGoWdmYaH2mRIIk9ne5K1kMgt0ASg6g2Au97+yLeVVVRIp59CA
+Oid8UR4QzuLrRR9+L2p4pXwA1Drh9JkjYpGXJGapF48e6qB+LZxsm64L1hp5y6t
uSr/x7rTXfTPSkkocyMCGYeMJyRmNKcb3wN8MaTqTIs0qnA7Ow2eNqVfqt6RVJin
sJIIc1/yEbvFbZsEQkvroojKzn8FFM0uLFZfWqWzuv7EntIFHfPbGn45paLNmaTi
MdRnVIhzqXdlpTUb0SmMhT4xddrWDd96fR6mY3rzxT2204rZDz6ppNFsBenlqZVQ
6FJXMWkG945Ow7/QeqFwuwUMkHQjjP6bK3JES6FUOSDI+5Gs+/7urVg6TduWFzDr
PXHvZQwvxcLxAxE7BZ316htwcICwB7/rc/J6MQquyLR7tQeFTt5ZKGSIx3wlmSIZ
Dg10c2ayTxerWTTYOgld6R1Gk3DLJAAxj0KSPqPbY0t+gE4vZx9/+B1HsW0ttlE8
0Iy8OoTmRh/G6lh8K28ijfjGoh7YFSr+OSOkQciZ+0QsPMAAY3sdR116qYKa61G+
AFi0QdxuaA0D8rw4CD5vXe9b75oMuo93+2daUtLhHGGwDIC28/6tOp8KUfwnTc5w
ir07PCauS0G3f03MGsPe/EWBqGxdJzqizAgaj1XHYsKp/oPS1LD6d3OfUAbax2KZ
hQwdrEvDV3iz3+Pvneu70IZQb1BqyJ9bZTlI5YN4og04X2iT8gwro2MYzmOdITm/
C0+ugjOD51NOt5b/CoV5xBd5nEAIk/ICKjGxDnRnMd5ceeLZ7SQl/f0n+UOQE7NY
/nBVWxAynyNN74x5KM+xXqEmfXrkwClgdrYrofAADH2FczvqFaGDLlZrXP0QI44q
AZa1QfC2XCXD1dfj/InvLpH2Nc9j1Hyy6yjD37jfbu2YZVSFvvFVinzuc4iZVfOk
yhTBE6RRhcGWJ9RGXH4RHW/wzTwhldxXep+jV1F6bOa13eBknPeiWCtQJaT9dmq9
vIAYyYOkCzCXKydPWSgSEiz+uQ4Azo8DfMadqur5wyEml6Wps6JI9TAa32OONNhI
IMa87Uup0CDJayPdpegnMIuwZ4oG/osRCdheGxKxu7IXoh30CeNcBjLh5k3BVPts
FpvtNrjlzujKV/rbxtIWpCP1rCouEm1Gig+zSSllPyaH1rbReonV8Ph6ZFBD5DMz
qRA68zCHxpr5+wTqnxkQMqM2cgLw26KZqdfQyhwM0t6LlEPx2GQ9/vZa+zz9CBBW
f7pkf/lQmK79Azp58TDEE9vs2PVAII9LgZZFrFUCuLlR2j/b4Kx6QAYpfFja9xZC
6j/kg5LnaMaP+N0YVb0fIpz0NwsQBZdhQo2KyvvFB9XyskHq4OhmebQpa21f6Zm4
79NPihhYSdlIOlxhfe5QeLNWsuuKVJq1QIIAVfbg285yA2Q9rfEEXj2lhR+FGgEC
7UBFTBxz5OdkMtUrvzdrRax1WEpXMziJ3BqsMvQpCB01ucKCVQI6iPNFHauHFwom
DR3O6IM+iPoIzZbTTN4tcOCCCiqeVqwrJg9oi5z7CQQXy+tusqv8c52K+AiqMtBH
w/ExpKDYPNjhp0qgVulWOTJfxiEjzTDtpeFjp5eGLDEuxb72f2U0RhrbR9HKw57x
JOmmMPEfw+G8f/EktFDbardSADP18HhKaaJuj3ZAQyxIBBvRYzUp0f9Q9aHJhAvL
We/ZXQ+AfXZmGm7UeQi45iMl/dzDyOcn7F/lRjFlyS78WaJHyp0B/F2zRYM15MQb
XHE+0Q+YHBE56Q0QwW8YDzewb8fJ+kZWeAutGT+/B48WvHTedqEsY+Ac+Xapg4eB
X92ypb5eN+OSZCZw/cwHsIlOx0lVK+W0jjFsErIOGvfxgz0Br8jt7JUq2SBFhc5S
KqD3kkf0Xa7CpBqBNWE242M8V7DMb+CYvwXvQmiSfoXrnSKeUcbKOqVB9fp+JE1I
N5ExwKTVccU4THFjbR0XiT+bYNkgxaVp3SG012UmAh5m98crJrYk/EmyVARxa8oW
9vIOyDHN3UGX1LQBoFOMnzef2WG8U1mPP5vt3WXtsKdfgaE17aAP8at5kQBqWOAP
YYNvaA2sVJMUaNQZ/7M/BUHw/6XS0w8+Cm94AThKS2Gnm8CT4YPE8hNag5+TKg1Q
JrtfsLGS+83X+D09IbvucJWsBnOeyv6HWoBoStBjA4+mHzWi25HsLpZoyTGEY4m2
s29E7j3w7KNdIffN91g8BCpxHnV+ZaQfbTpFHxB1v7tR+lJGJm8D/sWT9f16msZ1
tFr5pfLfsq5EbLtlgDYohhl7/PXkU4iyMj/W56lP6ITVwnWOgdhr0mz00CgbyZy9
F7LNzyMZVib9WorSsohRNE6dcwTUGRXHqZWQQzOlQiOvBVMzqgf2pqpAmTOq3eqx
2tQpERiuxESM0NzqAKkvfgdk5wpkFbWQA9tSF4gsM8fbRP52hpcaoJn5bWOv5nC7
vzvFS28ZCO/M6ngG/iU6ExmD0+/9DpGldGC7NIBqv13aw9nUiL/x4o8srUM+cB4G
tSJs/3BkdvGfNEJQpMlVVqCtpirhrt6AB5LLjnOpRWPSqJ311WD6RhYgrkUEtSYa
1ofKs81hS54VOF+eH9jrnzMLXTUGT9nkkEvekX10j9AKxW6FHVxHJGOpgm1A2l5k
xwAbiNwOUI07GrbS7uwoNvwnGOtTOywr5lAvt3qrEAiaGnjO9e9oqKJxNS+yM0t3
mt0vl3mv7IwItuTWz+SvE/EqDXBs2/m+bAIcP1lSWIG7LsOWeFMum/hyoAGZuznE
GXNY0lk1tSH6tX4zq1Hh1ltFlcf18sozU/K4h6LofACoAqqzXRIY/kdNSr18ioiG
sK0BQfae6JD+6lIeRsgf+HGznJOl3mgXtmStFk8Cv0sndbrSgGUiAdiKJcvX9B5t
0j4St6w2emlZe4lI07WjB9Q/2Cytk9GlzLgJnocxu9Bo90DlOTV7YPByGkdUnMab
ZvbBprMxWBeX+2b6MwSOfLS48zkHgqGiovemXVv1VCf9QTYqubsvx4clUC66VAup
38HEPsXMYPKBtX1oHV8swnOKLWIxsaBP3Lqr/P7CdazKT5E2kBHd68nCNKawW0F1
dlRvHSRy+QWWkVsOLOspzfuBxlqCnoX2J+xAw2eHIRlUtvhJmLpIx5vIHr8x4JR8
WC+lupYVPnPwfzC4AhOkD4GbQ+CgqwG0TK54H0NDgG2ywFnHmtTghfUl7S4SDBFv
7YBjCnrhzwNIaRVW29eL7J9cLvlm96fT1FQbQVv86tnwcWoDS/VK955Tq+KtfmN4
8YHdu8/EE23Aah7YWPsDrsv9+Iz9kk0rBE5dV36PNJVxOu1xzMzWZ8zy1E7WJmt8
1x6c3LZ9wW4m/fYdkGNi71d3ajOa50t/PfrlWEvPdSfDBc6m9UQM4KCF3kuIElIp
AUW97JL4xXq8+P4Ydz32zfruw8mNCi0wbLjc6Jw8CCST104e2foLokLMZACs1112
VHGifF/BcwkFmcTI9RKeXLegVvbCfRSf2LhHz8gsr9ToBIIqndliGNC0YeQoghZU
7cRcA4XY8G+J7omVmLtuN51BkNlnY5Hvwlcg7wccE1ZlB7ke6wYjjm8JcEAoVFew
sqvB9VquwwXgu8voGYO08/DXlWvwVDHgEM2E6KBANHshDan+Wm0Map81dBHOmjR0
Va80oZJyOeLJadtSocB/C9rtnR6jEdjfPmvMBPgFQ2sdw3mKJoSXL3/wCoprzWvM
blnGmlV3vZ0CEn6uXhmURetSUB5bKEnr3LlXJpnn+L/LmErQd2Xp9ixr2SWs/VeO
y52Ris/1WTGn4xwSOH3PAiLOdJCpJcf7oDQxZaBGxzYFIZqDo6HE94WLgAXT02w9
rp3uxc4oa/TbOhsgeEKLfy0Nxpa10k235AtbHSyT2mgrJgnuTJVkulJ2P8XrZ8Ap
RyIVoxVwyOdPqcgZ7i2JU1tGMdMBOFLeCVKk1TVezggEM5dy/eTStSS+5pgwaBPi
V02ijpgQhN6OJzQKOGnEaJdWl2qFEgH5jUbcrtodc/QixITkxKgXL7rYR/NeHsIJ
bcoD2FPDdi1XM+FGzEF7W1Y+rlh14Zy7vuwXHgKGS4Nma2uddxuHnm/55+oLWLXm
/e4y+KdQQgcqgYXrrJOxd0sknhG+TAgybCIQ6T3CdS8bwUkXM9TEkHnuPmmJE1UR
IzhxPRFpYLrB8xC526eyCYJoElYRNJD0IL8FXY5MzLLtd0arZ+Xmx27+EO/fQthI
scBINrtjuo0YW77OGP0V6SRZLToCanXj9ILzjaJwuxITbWZEqrrEFYwPSvVeeYWT
IrzFuADoIRSIKSVVjzndGv8q8aWsuflUVFbl3q+8IegYE+aYvJVkyt65D316mYak
1nWLZjJ3HPR2LSI9a/RggJm+NcpGY4faE/bZOPS99ESRK0MzrtIqflzvbvhnWQTC
gCaiIw4qEQizq2sGnF4QEUubi087M9wlyVKqX3D4bYPod6mbA7r1yZXiTx3mhCHn
4xPpHEl9RX2NGUtKI2hhSp7nVnoyVo1c9A27kUxRR/Zml1TrFWabADSFG/q5hMFu
ycjw2/DzHc32gYP8tt9kaBKNtFc0iTybee/h3GSrMAMxAPYxb8izTr8ZwbDVDFba
razguHk0iri5NOZls0ID1FBMHFEs2jMOgRfGZUD02VAXv0/G3mY7uTAhDVs8um+O
jxsP2Arc3JsLeZwfVj8NqxqjFXmalACgX/fbD+F1ncJCbLmFRfSLtewiSHPJ6TAb
3qJEBG+xNBTipm066MyPquepvd7rXWKnaqOwqSGAZWfa/5MgdpPcMT8qDA0toDe6
85Qqnr6yUdGAsudlV3XXA6SdNkgODqAXDGbLBknrglqmG5iyyEHue0TZj7ADjULD
TwSMQ6p6jzFwaWbDv+JEOPyd8n+MaYvmi1iuhSlc4dsGxZFHpQs8hRWdVU/nLKH7
//kciXdZJkuxEKmemD0cBCwTwcq0EzVcy7MADg2Dj58Rt2ET1HXvTivT9g0q7xxv
Cn6sAchPpjvXG77vQg39PDpRI+x9BfYT0ebufvU2+HjYkUX6JCkHvMgtnf5YNb4g
7geOqZnZpBb6hYwdYAHPd++/yBw7tMUrlIaZF+k6LqalTFxo9uVJCKbh6MasAQ0V
e64PoA+ItR6F/hb8JcZ3ho1rVpA7dbFyVpqs++How+oCcO9LL60yEGI0LTVTWtgV
qBPh1cKwNbwaTLAHF1TdtxaSWuqV1k+bBgjZdAgksKdEEHemgvpJ9hKoY0ZpMIpe
PDpnNDzkOzRC87R0KCMoXdV42NTYH35FDdTt99xjzXAgeBjx1iJq0MyKspW9x97d
pA/XkBWRETdQacRRDQQQKvEcHk48NBMYdMXIheA7boFGrghsM/j153ctB4/0IIIz
SmxK20QKxiVQiw1nB4MSEo8D+NCBaFFsFS1fA1+UFXQJT7l6fPUrOoVIpfM7meuv
x1YskKMGKqgdvKKIxVmBTivxC5iR0/eFRsRsYE4H5gQX33jGr0GXLfcDIiXxyVFg
tYu1cfkonA3cndnGKCtGmIagKARjPqbKrD4KuyTCFGlVzDJOps+eUcjD0K1TU8Px
2tlHFUb956XJTFx41G3fMg690RHeShgNy4XJw/9Y4PBXbpcKzRJNkeBjSzYqoors
ZZR3sR6jBiOkvRemdrVphfslPj9BUOL9W+isogGgsZX4SNebXJpi1qUBiES6Np5e
O1whi4B5qPwKwXfRKaFlTPUHB32w7x4EH8SngDUIDp105VLiYvq7KouFy59PH76C
2Kp7BidSWQB1fK6mCNTFZYI3pHDs0+JR11BuuVhRppvi/OimMtUfcLHpyJhqo3/r
lO0RdVE+HHUHxHNRNAk9OoB9ecZnuX6Rv9Uy2ADYIt28LIFUulwBjPo19kLK+SxZ
nOBHpfLfnq1aMv1Su7NnpsLardP8Hz+IFqnHPJrDJuqgAw6JxTKGnyoZctFkKAkm
uIZBhfc589PaQcra+tUHgih1rzh4vQ8Yo4+TrOc/dR1e9cbQUTaKJPFIM+7FsO2+
d8GCtPKA4Hok0l9lCjYOIrVw9VttdoKvmnzOkg81VUVDu/luVxSdZc+08qLfmImJ
R0UhkjkhykYl79mI3P1P3biny5IsiWShdjtb7fmgXNJB0NLSQn8UqnPh8bQb0Sqw
Csty2iAjoy9I49Ev94GlUkakkJ/dc7TqUt5T/XzZynGfvTeMboGZd0DLCyITObpU
7NYyVqgWlC2WBUkgMtO/T+DqVbrGBRSNjlceXWnD1GFzvGPoFQlUJYcUQop4U+H6
04/nOKK/7p+m7Iievdv+8mdu9aC6XXq1LM1yjLSjaZ5r9xgle0JAf/sF3d7cHqo/
dOIuT6luEJIjmeVY7JLDryfCHdCnjPCiORcQpjTg358ScTDTZ0MJIGMGMTWvSUHr
TRAySx/jqu0xcdppu7LYsOOTeUc9OjrpHN9dwSZQH/iYjSWPu7GrrDWD/ajcWqO0
vUOONYeFufFYM6Vwat+gbpOPualqzlNVRDvwXMPeOGFIU4Mcj7k8gPpoCH2HdyqP
YoKAcv/2HddYxII0c+sup4iITZBoEAt1fNR8L9te+r3FT1IsvYlLdJwoph8qDm6Z
m8EFWfAe7ZZsJAG93eivojyAAcenUaB2M+5DaQsmAhsG1qw0LeKoRyrRMLER906e
AeL3DE/tGGE00/sXIT05ZeCnnuJ1dzk51kX5digF4/FqehjWdZhUs8TVhkS4dQu9
7tycxrMxFeRwdkhBzR1Konjug9l7bmQFzWsck3fkiWpegfqxLZhKWZIE9yvwquK7
ffd8EHFMv/yon9QJDH51zyPTESlwcjy6wL3zTXpaE1hrm6euyjxydFMtVNg1mg+1
gSaeuxhw8wxtHnbFqLchh6/m5ki7br4uT4TezPVUdtFAkFmVNGQXJSbRKFJuvcYg
PP/jxwR0LeF3qgej1DkR/CJ9G2mXskqLCgt5ArhZldovEIxUNlHLerhmN8F9AS/n
mmzt5X7aCNpxOWkPDD0h1NRBe3jtuC5tH/UZH1k0k2VRfi3DptPCUspNjh4uFqxT
F+Y6rRIp7XN/3n5g40wLp6vDIKncVpUJoe9U98vnjCID1ZsPwUztH6PiVjTJsI9v
T03sYjH5h8NqD43yJMWSlZb8mjzL5+A1u/HsQxioHJBhHyRvivQNFmJ3GA4pYnPo
M4jdA+Pa96/6dfxqZWrTFIUN2D4JIedVPXByGfX8yiARh2036/ArLSooEe2YW5RU
Kj1SIJIYNa+5pVKbzUpaFTCcX/U4WwWF7axTSJD0rhqiWob5l4+mB4tse5yUMviW
dp17JG5l0gtt5pEW47Y+uMv3fiYl2fJSF9AWewNGewa4oDQyNp2bdzlgEp7xpM7S
MPKe5fyERgmwKZyWbOTHsY6TeoAerxiB3cJrdkW1ycyedHKMjMKRTLENbafAYjbQ
od1FAlP43pFg8tXD8Fse0YkzVzpCZBFlCrIZIwJ9AUObQTh2NB5YAGQkzzMwhoZ6
z4n2CB7b8GuRYUKfmxbwIqbgp6G53pBY9s3kQyHnKH87PdxoImY6KY9ggF7apVnY
n8+zEgAcYMK8xZwb1vUYdPxGP068tRWldjOLNlMiFld/aO4LwDvdGNOies/nripP
nyxWn2ph0O9VwWGDklHHMYek8TgE2qKXi2Z1GXz7cX3o7ors/orxNCgcxkx6DAnh
JyULUmm/4KWTQqUMWBo4NICe1nx8CWpJlfIshlnlHma+flo9eV6mHC7Z2ql6jpbh
Y4/M7KLawLA9JHkrmeku7PrbbZTTdSfz58RAPbuLr+1A0G8srUZ3/y7fxoPkAGT/
3WKbyh622+YsCvErGEKNZ7L9wnhGZc+zkiL4xBJroG9bEQCC2mjQrGMS1G24XuL7
2FGJoe4OUhNf/jVF8UYm/Ik5O8VakFrjp/DdxQW1/bvp2VOFbxABTy4fZikZF38m
NwrY7S5KfR8y0opvZDB8wa5K9Tc0tRx3dn7HUfg8NQYfc4VBEpZE0BIKfSJ0zU+7
xJ1HvSvLXh4G7usA4eQUPgVyI54wieMaRGFckDDVgkmsaPl8jpTbktdZuXraRzWE
Ofx1EwXsp/KvNPOF1ATZMmqJvDLBs5tJj0jWYLaa+VvL/mrCiUcQ78tfz6gXH06b
pBHRUolIw35huBiYttagVOfQaIyCaGKjHO+6m/vu6IHJYcpZ6vSnVDe6tycVG5VD
+g35PnThR+8YpJi3eMjPRpVmbFNwxvrChBOzBJ/QJZ//Hc8cRtvFvXKwb2QmdXwN
iGJeftyVM6RhrhyhKEGJoKko+y+IJWXuDGPjkonLuzne+bHpOmu8AVoj0hJ1PAdN
X1vx9Khf4hDUCsmqN5Kl4jjYByuF/LS9QEDPR9Lhhn6E+qM2demjz4z9kBUIQvnK
9X79h90F5vrcTFcLp70pHUL6V4MwNzgPjPVt7tfVjDwSfiXVa4vmVS4Xl0pRIG6v
94v0fcos7jGrWyLs1FJ6ROWOYDYwpglZx7nuVmrRkreLWIWUAZYXsuVel1rvvKk9
HizRO93twkDC/ZGu4b0VC89uWhUvmbnDbNnjBi0kWC1BBsrKpKrNiItkNKLxv0BC
4dLN9c///fu6YlSMB1kT4AAvEk3Pp7UVBKw32ZxTG+w3WYUZPqvYNU+bGsVZVnA2
xB5iQkhHcOSB8ivqppVKv8zPxfRKLRMox6f5NGLIevvK/QjfR3NaszDU1lDdZsCY
rZ/Ssm67pJSsCTahUjydxkjACl/0EoE+KbnWK7R66tPMa4rr735hmKbphG5M9Sxk
uc7nBMBmxkzJbrB4IV+kCxeZrnfMFLmbV79NsoDIjYaKzdSmLczDYZxlnJuaDSnS
0XAvDUeRpK8m01EhXRw7wq++vYSfBACINBzH41HChusDFvPzgtYn9z4RhKqrace4
rzc8N2ZWDaB6fk2iDk4Pu3h7gH5ZDz+Tb7eOEWLt+Si7WrmdIOVXcq/YmDVt41u+
MLsy1COkSeRefgjNknheVfVJK5LIDmGhRe62ZhkcqvJmdg0RZUSm03yazAvPxllK
N3f2/io9+aN4uN08ML7/m5hQAsQl71qwYyXCSm7ssMfQ+lJq58XoBdmmbUdyATrr
fdHWn1YECICN3unzCJv1x2e5BYmKMgshvswVvrmPRZdQIOvUhe6TbAGFitqmSm++
+6K6H7uzVK2gnKddUBIbexL4AyhAftJb3Dwk0iNBZmmP3K0RVsL1/wjrigeJkaBu
EOVtsGCIMElkq6THpZI0wuPTK9OLjh/y+POfqM0VSqvlAO40sbnLqsCBAJNF4tb3
SY+dNOHlAyL/cv00tTy3PIwGuwGkDse3SrfBIuSF3SEUVOkxq2IMRu65Ne3bcOOc
7m7tlVo0pFCFHTL7jwa9zEZQH46bZxn7yTiU/D0RPSGm6x6TDnfWFTff2IHz+0y9
Vk5iNEEy8xDDzeghwGQRsPZbu1QfNS2X6Nl0KkAQKRHIIbUhlQjktzwahcO3KxK5
Vn36Y5RyIMalRyZdU4OSlkrcUmRQrV1by1RPsvg2ddxrObUdr1ylHa4H4MVS/3v9
cY1A9mP5oWI/NbobLew+ZGy0zacEpFbJ/N4/fin5JwDRaX70nF2311TqByj6Wz2w
ZVJlaxSYxbKjLt1VTPT+bRYoLhWZzBGXRDeCPDk3yPx2N7MN52/1enSuWmDqDbuM
KYhBzfPYjCeuLzbkGZ/ihbJbPwx8GHK8T8PljvhJcUwWirr9xqGxHIXBfKSjXLhs
0LWL2g13vzQ+cdImlvDOgvECykP6JroHZiDbBagLC/e7qzVaaU9/ThT4ZHW3Abqo
kbcC9bb/mUnwWQ3UQkwa113yAl534nKLLXUYJxdRQ1OgbPXP/VSYUdQ+y2iOTIZi
RW/FJmnbSHTpjcaGN/i6IHqv+grdoB2D77CIH2UheN3jbxj+0H/a6dFhYnJKjTGd
hWPzcGcVGwGRkkvCcJdnaWkxysx5P3YKwrvtop/CrkJJ9YAMNfXJXvJ/XJ7r9CAh
GrizidIWoIOoOXjslxlT8JQcHEeHCb3HNc5uHekIViCtjT8da8bJJplIHBMhPNos
ZDF7WMdWHO6WJbwX4/QZJCeGtQQhV3rhpdp0Uk/+6dTb5IrUjdFIRRkghUwk87sZ
vh7v3/grcztvED8Vp9RfM8PfXJBGx+JcXSLjWbV5Mwhb1EKLVfJYu/N5opvFOccs
ERZdG6RQn3qJof6V1FrLOyBW9d7VbMNriAGeLDSvQBIDzBmPNCvIaoUutmej5M+j
s+vzHvLR+HmLcB1qyjNx60jzf0hcUVFI0YjrEKSwmojHtrxM+D1KU/GIEedOnul5
qKhI0PgaJHyq67ws/DwqJ5bKP3Nzrq52FsmduiG6xNPZyL5q5tFQcGJy+6b1iAdd
39aUrrn5Vz4n5Z0cXXuVjErlQFAoabms0iQjDhdayW5VQlzujvBu3la9YoYUYC7r
G7F97+VUE8Gl/sZUJBOEWsNZEwEM+uZYfrwgJsb6UB0bNrq3AJJ3Z6gmSOxLYN2n
ghuGb+A0hH9HzJm6ZoZAPltgcC1jpaxiYqfVrXfxspqV3iw4Xq2z/K3MIb/HFZIy
BCZTEkhMjxbdnL06vVuCTGwDFazHfO6SaXBztpP46bushDTWEildVjgmz8sgukgc
GXsVjrCEfhH5UvuiVeyADd2YpZl46bUQ1GMAET16Q0Dne7CLq+zS4RSxBVKCc9mk
oWp5zjZgF04DUKIKPZFphkNeRKiazfJoqCWbE7pQGdoO5vgOxONdXLQbgOWYGpIN
hokvmGWigEv/2kaUGQY5WqWzRqYOxexAYUzIUVPbkBAYA29G3Ns52EPPSFLMNHEA
0G3D1C21pSSEkizGWktb2IBg49jh1wUtAb/JVg33k5EeXlhYgjppcF4HNd9yCBZs
h+oYrfnTNBAjG1rEKLmjuGM80xGxBiT7BdtnckdgyN4HnFk0/yjFthHHZlsQos1B
BS6nAWEMkdRz+RyOc+A7THMe2HyxKSSke5fOeIsFcbfiXIyHYoFOgnjhhRwP6DPG
uPIJgccx9g8u8LISDYumuiHUisNBvD5sCQl0WCbVOk+g8XULjhCD4Ot/q7RQ+dj1
P6dOLF/3irhNNAJWNp5kO3bCnyDHd2Q4qH19TcRuGVhxg750uvWNYLlBWjwPszQC
id0WC7NuNYmxmGrUoImroLs1skawWD5NbnS6rAja9bTvB93VRVmYBnf2fwe0nYQX
FvHTXpg2BMOCgts41CuPaMnrN7s9NDjDeGRUX6XYS/IFjLWx//vlXIfWRjduRHdy
F5A6rHg667YInn1IjXCpqo/PwPPc8AVByKkIe3lvyQ+fzRCHYDDFakB9VbutwNcm
3RUZAZMCXfKrMFUzdLdmDfqVWBlN2gcnuUNceRrDeJMj+B1QUDW0EkRz2paAN8ux
LZRPWOC+QsW5AW/XjfpB/tWooGxiSGCbe9YXO1JDPR2E6Nim7UqDxhkeLNdSKM7N
3vDxGx0ej1zQ9HDwU4uREmQkrQ83QaPytmpzf68eU8q6gD7aWauesUKGLc22qNmn
a4h38wpiMWRmyHXiyomgEgXIqxxrPtwTN5Jo3Ftl6beWj1l8tuCXkK18az30yRGX
wX3P4QrOuxueIlVZ7pBk6lB8BtqTCcLc18rNkR2353r2/xuMETdPSsQe3kH7yJc3
G7xG1QxOKCYSCzF3gSVXopjxE3YDXb4FXn5jV/ZBYtarVQTwxXjeWKwGJzyoT/3q
oh1YzgHKyK3hvR+ZHzvAgwJ/6DaZoh3X7EGjSE4Iq7iFOcbwO/iExseEU7Eq3ZVm
GFp+oDgwlvywOgE16B/z2jT1IrAg+HVqYvzu6BcPasZVkK2zkkWHcoWBt/tc47Ks
4khxkuoSnqkbBKPGUeVVng5a0JBg49ppu3dm3TcBt6q0aJFSrXJWEJzC+FJ49Wi2
GDwkccObGWWiSQcq7kkMD6bjR55buvHLvn/SbbeSBwYFcAri5di0QC8BbFFoKC4s
1tqZ1mTYrQT6bvVUhBSgsp08nyJHnk/I3LgpSsLGRmQdCWJhCdRQ3uisYKbYyi/l
US6mln8rAoZx0Hy9C+FnnfFswv7VQj5WUxMZGma5+2TL98qTzgEyTcmePG5Ra4LT
fLOdn+/hvonoHrtTQkt09m3t0m7mBj4Pa5Ar46b7U/Fcc/hGafpcSPGgfsOVBHOz
EZJDRpSqYekemmhqNI8S6yCdvWMP+kQnIEjKACLArD160wlkj5qX6rl7/cKwa4Fa
QZS6iE8L0yjPqNweTJD+6LEdhh0oQkyCqwbCl7ZtJ4zuKj/x3r3KXYQ52k/e4qRp
M/ktWZsbvtV16hjjUevCNAoJm4REN4WHieneYENDLkVwe7+wd7vLh3ok1J7rRN7G
FzJMr5T4q+lKqwz9sEP+8Av7dqNfvI04ye2pJGIelOi28gXhHMAwBODoT1pvsTwb
eL9GOjiGChfFjEUMdJrLKw==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
poCfiKbQ51FcLyALKqXm/pzzhiKTxZPo+UHA+zFi4LW+HNbLj19dnRvTZA9yyq+F
vuB5hD34u2BgdjdJ0700GqbsayNUyKrNmp7PPwDR0t4BltzcJ9NFOWUDJj7rqpN5
mRELTiL2LdjDQrFhe+Rp5MJDyRe8NHAQhdO18bbg3Bk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 12558     )
3qYIFBvDmHnqVO/5PzJn8HNRQuKcnfgi0WPc1RGZ26h9HeLJmzBYK7n5ICK7sB3s
tbKW/+R1tloqGUjavuRGa/gMViM6d/ZNoFAefIb8+HD1+Dlkur8FSNPygpfwA3qa
SAcDbYObKu4L9EQL6AkWI8m9AUde6oq/bivbiWKO4s8OJm/tI/KRJilENkpPkOPN
QuHZCcocpbmgx/Sd/ApDoC61BlbAKF0bbVTsqUUvCZDgtjWDfRCJXbaqsLF+gxAh
4k+h2v4eyAYSOd4x+qst+hrtDutqZ32QPPt/0k1Rdlm3oIcDAPuxEbUk5Lg7rwjh
uk6gT+8d4md4f/FVGCeR2yVCA9B9r5LbhmLLBoOSUAwwCItD+WtGA4PCMSoRbfdV
ljHZ8SJqDTk/9GMvtPYvuv4gUHuv9gqX5D0KLjct9H4EDt7ygGsOYnaHDtZeqh8n
tkFg2UVBkTNy953xT+BI8A==
`pragma protect end_protected      
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OTBuJZ5RdpR3l639cDWEa/iwPCPaPOmf6lCywGP5RwElzgWKNTRvA96NrSqBxjYP
Lp7HjxLVJO990oEq00ZhQxE6VaSchXZNKTtjSMFSvM+li9Nvl4kmS2zZ4SFEDMHf
uvn0WMy0sSttiv9ZpZUNjwSzSoiW70SSpMmenGynU34=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 42647     )
OuZ1lEeWg3YxcsOR07LZaEcEcwAtyKxIftwnq0wovcPwh4hbgg7DBouVxeRSrk1w
yZRWXwU2LNRvEc6QFxQMaiE1cMzfIK+avf9lEr/Wm8whmF6RELea50kskqoopA4E
X61CMfrzXz40pbaIjUoEuAfCPuHcTvLTpmCp4hJcxwjhsKjvRRPQjUl+T5cwYpJn
lGDUz4K9vlaXg38SEpUu1u+HiUoyoay5IvkBzubYLosXSF8rrXEPYNoum+ggMmYW
XR086OXVTh/I/mK68UW+gKV9Kt8pUUGBg2R/5cv/Zuw5uWYCPioMb+oqOwWSSiij
r3N7y51tLUq3MpGux3C30mHbsnuXZgctclWzrY7O1h35nriYCaC5Wp6lyvVXEkqU
z/3PaHpJ4qmmxfOzGdUsXEAe6xpmUnclaVTPFwcnTB8TH+/MOSCJp1zYI5n0gyZU
5QjQGFJCbZEZGgS/2GPC66/2s7lG/3soxEuxE3BU+aKRm1LD2hz3/2Gmx0BEZYxn
ljwKn+pD3rIuXg9Dc7WAPST0d5bTK/ALcdqJhoB1M7Fr5PoF85n8XQl8R7WS6hnE
z3m22GyVckAJ6Mkx5aHkIkurkDqszpjWSH4QyNJ3Wg8EFPxDPqbfvbrX7eWklebf
zD+3/EFK+9HvpyLK7AzFRudZvIxsOHvz4/yXB0Sl3In7k4ShBQ4Rz2zauKvcLsWU
4vVO6PBS3AXQYu4nabVB+SWud+gtLL39E0ca0ncsGcPdGOGDle/Oyc2bomdlB5mn
ucCvyKF4DMAAC4FLkwRdi+zHA51dr9ePGtBHpe9enfuGQZx9j8XLqaKy1uX2Hn4T
gntKpMxEm2sLbwCcIGmhl1bAqDAB2ebYVZViizDYsUUrM62U5CKXii0ygLbGk03s
x+e03w/v8ISB0MPV51Ue8FxcgY8KioYOiCjszI5cDPIwcIyOM+ce8l887KlDmONq
hNYf+y1gqy1fuZHQ7xHyKt1cmVcdeHvy0WSik1F8pesmpbXQVdT1BWQFoy1CkVFG
Bym+OgHj4dHxhLTpi//tE4UW3jvhAeXfi1koBX+Ht2CGQYbp/EPMakMB0FXSkSZe
rxkoCpbc3TD9dlJhHMHRhlaB+eXUGhkgh53w1G4Ui1+z/q/gcdZlfr0yIMolXXOU
olwMLfISHS8uh7Dp5OEJG44zhsKMzJFpGYUQL+Qh073rEYDS366oUrlXWYBV/fLV
VLBLvCIPCPM1Ux94itbHU+IlhfLaqEcexKiXCfVle6tL6TTNK0XCadgoz2cwILXr
c6cgx6dFBM+UlHC5qHm6cKxYJmJ+DAnlO+eGoq9e3HpithN1xcNqYBNE0iyk4TL5
zYtEoQEleyrionpx5YvTZ1MXuR2qPdVmlAQ1xUVxe0SEKz9as/egped9pPCpJjxW
TnhVX4ZAosFCm6Trj9Xb2zflWUwV41MGNjY9tyeOzZVhE0RDTz+4O0yZD98tMeU8
ugJdsFztIy6/AslXRFFCzmKvGxxNEVGfpEqSOhQwf+RpagMOQs/RkB7r/pmr78B7
S2HsfodeoNnPvZnvdvyvMzEUqKP0Jy9v1LgOZoNzYAOBHWhld32rK1vmQGLkRTYg
YHUkEHaJ7rggW8D8leC0b1d/F5OtAJX/lT5DCip192xGwS+/UvfuTGZdcCZj7FUR
G9S/g2tUNzBnwfSYGRpyJv03iwpIAidulmlqQ7JsYobhRwuepY+yAiphnW/PkKtz
qW7qrHzGC2HqG1QRT9XwTmSsikb+7J2cWubZjFYi06dSisGNFTdEyuYEfc155F4A
dniQKgmVRuvJo/V78wfi1RyaydxkOQ4n3KvBtq9mTb9u5mx926jPIKgYO3Xw8E6n
+V+wAvamZEtK8KiozdojoWL5sIfU7GziK+hpTUrXS3s6v2peWK99xV+YcMF4FUQK
wJlrDfw60cUzvdwYwL1VYPVQ+Umtc+upOZdn+4+rqofN+K3q2+8fjlsEqSgtBiYX
hv1a3R+6mu/kESZspVOl5R/8zhOL/8ud5mVXsC3yZjPE1UQ7FCB9KnrTVxr3sqtT
bxH0VxsnhDBgQTHsqPAp/aOIGSYbpL9/ZYXRMwimznkcz17zI8gqzQhRbfFBturM
QtNJ9PMlMqjnxGwzZ2dBUoQZarlQazG1mvfg8fYyZ/Tmy1/TUebk1Tqr8IxIqoPX
KL+7+YqncZg6XtgCYrTcVRpEzkz2MiESWfPhKOzTpnUEd3A/yPGokVE1yeaup8Wz
bVju+ret5dkXmsI20CSC0sRgx0iCKpqYwMfr/KGCDPZOiEk4z3MbwNl2DzmFfPCZ
JCS9JxXp4Xsya7YZsbN2Ly6o6KFwcD6rqwbBNq/9eHvrQ6BkicVW2uYAwGUnpoT+
IGAmwQBo6jMaox5kVkZCkv5BCuvUEuH+4uGgxpgkr857xlJSU/WeHtuRKIfxbjfw
rvYG/W8T2b+DbYfWCtwvRALhKcBF/xAmOPK4AtUSbkRgjKvd3Xw9N5aRSocdoZW9
xG4wtDLNNJFn9WbmM9m9O5NH3fWitGnTIluEYHmbdsNbEVjrIohKVtZghm9TeRs+
gcfk1sL60G3Jz0CV/xWCTPY0OZIffKb40IG29hU83kc/DZ+wHBMP3G86mz50Xfuf
240DXADPleBNGfYEF5793HoHJkFXjHt2l5LGYEDJpAPKHywfMEOjc4kYuTPX7Vly
GqT3IXJ7GVkTZsvf4p4nqByt4+TmZJCDdB8X3N89N+24pPaQzoT4S5q/6L3qyF7x
tJ8Gl3kTmP7v2cHE5Y3lRaFzk7ERB/CGmhuMnXTRoGGpHdO3J0M67OAt6j1Klbk4
x1v776OP4Fejatsf1IS7gd4V3G+WcrqsE/hhQhnYKWNf9wIN/laZ3ZmrxInsF9vy
s9V+h9jjcuJX3R0S6PENAAuXrka8V1atvMOg9Szpm6pfcPOxWP6V/bz+fQOXoz/I
IgEpUwOwnzq7v7meN3vRovWUsv2PlbGC2V6f0GjshJd2MGwAbENnNxZkpN9n+uHT
AHIc4ZJNVic8HN4YC1bD+yXE7j4EquxPiue2840bVP9RwhPMFl7nRMnURb81PWrd
QdX2B4eUSI8NPQta8q1xh8oMU66BBggU/mMmm3aTTyUoMM+UQhId3HOoAlz0mQHq
rHuiaPRoM7HfP353EJMfJBmvVM/Pxk1Id7Fxl3KoeD3fjYPnB8KSv0AkdKeEkX6z
cjaKkpOZH/fibS6Uix3I36uq9nEgLi+J2D/jXJxsI81I/VzWDtGKFF2sdynVR1an
zos+vdQ4CLuOD6wLHBB4hFnd1wUwgeRzA/ijofXoRbsd06hkaqZ1BlN4n4Q7668j
i+CjBiwFVPtBlDMdBzXpt1KG45Cq0WMibzK+3wogDRePkbnOcTnYTcNkWQ+m01k0
9WUmLAgsWhkZt7jHVQDBpez8PvQsSTK0jcBkoiDY4YsFSyqwAiQZ/j4PLsFkSOL9
SMk53LtnHsziLLFV3FShWyN1VoOGU6RqYIphz+ZwpvDT358UfL/agBNuMjlxoP16
E0dhxG6S3YLGuEr57DbTnEQm0OZGRXgIab1L2wQASZ9NPsUfbwZ+4bsnioLaSSEK
EQ4cp4C3/26iNQiBEnmB/jSgGy+FDodQ49DyJTPDDuunUk2JKF/xhLe+5Jq/GH2E
82MWqvLKh0ngGHmhHEjXEhz3uCz4gPKJHqfi1PKlUTmIEIAZed7c1P45H5/dxPMI
5dAlZaxZh8ZmZh0XPtCf7heN/4HD8GtBa/5qvFKJ4OzmNq2Ym2WUQLHix7SlYuPF
rWmbGpp+V9l+xQXwGHryMV3yrBlW8GtEHBLDNIQlSy7IXc4+89/+cbqjMj/i4pmb
ps1wEOTJBOG8w2GBE8j+qZ1hahwKD0O8SKkmoorSFvn085fzXPweZIrYmhyQ8D3S
rIrm4E+aowbfixe9J/OKsfy2p+cuuE+ORlTVHXGP3QM+0RgCVDTy/2tAsVVa/d1M
LMZhxVxz/OQs+68NDoupOJoTNo1UuqjrJuQRqvHpcXLBRUlpO1Zkaykuh0VNiPtj
+oYJfjokcoVa3YpCEDK1cUVpt94KxkbrBGHgs7MRVroR70dIHes5Ig3O11zswGsL
gssu2SUmrKiP9oQeouXZaQs0dmlNoiUp4HjtWSyxkgzGqsg0Fy0HzMqtqPfQ9qNO
fCo963zmIQ+2mzS0TD7+uu93a5z18AKiZ8aYLxPmCLlmJemivLys42fL8pxlBGmb
lV78IDjR2KTnIA9wjDY88nRrc9GXJiUngPrjKxXTYPs8tH7T5YJQnBcI9rso4tWr
eYyLoHhCH029wKc45M5f+mw+zJwfhlBP/szumU1hXRBIQknUbQ6GesFhxN2wgLHe
DtejRwxU7Yx9oqkMCG/Y1SRQ55F77AghsjOrOJXRazJWtvoZi7CVYFuWVY7g58pR
bg2irVXcv9JnEIT61QLwK9xUV6D7vvxc2yzYx7kKJproYTqc/vYlAjIZyortJG9q
L+Ug8R1RJiC97VqFcF4JSZ5+2ADiskGVsGW/jfAEx1Oab1NM6S95nVX4sG28VvER
Jm9gH4CaiSYj6GW/RJbYvVgZgtUY9XXsVJwwMsL/xuYZaxfi67e0ucuWM4TA9M5E
HD+Iau7R2EXFHafN2pegRaDzmib2msO6l8kR4XNoICQ3l6OxnTLCD0nDVnqfnT8i
gNxYzsGTwmjuuNOXQk29jIsCXApwjx3qjkjBJ7y9mKxOUsgelzGQKpCTXgvLp2yx
nfk9DXL4GztM6CXSsWhB9anHTZEkBmZEUpqRC5F3e25XQmtEUG6zf81f4CE4WOpD
4FQABUEmnuxkEKeiDODKqAPJN9K204Xkbhwk+sB35CkCdRUiNP/1W9zj3DQiAPNe
X1MKiD0v4dKAWs7KHJqooibivX8l4Y7bb59UZ61nX+dGChJYEJs4lnS3LHytKWtC
TFKSOXiLPi1guAnWMUXtM/JwreFnlvGzw66OAsijeJV9lkhHPoPPg/Vp7aelw0mG
fO9cwod/BCd9ZlQfsd6yIIdjNnBo5HVzzvPjq1ev0v6YKwnhYvegIQssrxP4m2oQ
bEWMCnjF4R5pyEU+kxEuME/MLTDuAK1hiPeKup2MYAxjXuq82WdgU7QFQZ1keOrM
+YfV4eP2iNbBy904PShNReA4M8G2/NLZVxPQJ+ZpVUgaVXVXgxS0Ym3Ohddr3xd4
umkLzvfycvBgL4eeilIH6oMF+dEQggY8hfypvvFEdYH3U1wL05VqJEOWITi2BrCr
F5xLpbSfORWxuvHqxptFswwgbfEpxsYUUaEHBmrfpF41uT7Oj774byEDJJHySi5O
L9AIGo/cQh0wfOHhaTgJLoLrubsJOrXYRJ1BkW9RsVbhqh9wMU1tpomxQw/DHy/r
kwLRIWJwQRboWxO+x4LfvKBEWBtCFp2DTW6JFGS/j3QNPTvZBsFW4Rer0Xpkvmhb
3Uf9VMMVaQm5wqyPUqQHYz6Jw1cZDIyLe65QaEXQBzLHWZHgyaygDNPezgpSkBRz
pJ7ES0b1HCpoki4iMOS8w90uIfqb26N/VcYAsSo3MiHk4Gnj4MZpU+RbepKDXM40
9xoBdv5vOuObkylSGisZOG1eB30+WBfgfJPAtOEdGTwwI2bOzH1UOTa0OsZ3jnIN
+nRXy+0SwMmp5oeRNggOVuStasRJF9q9Ywck1ZkPaLFAmr82zlirPJZd7a2lUwES
6eymfhQ3yVT/W/nIc8MVKj59MgRkMav7wimGnsYPOdt/7YIOCNUHtdLbxv4Ngtjs
ZMOYXfqKvuYvBYbqvSumJkS2v7Pdrh/WGnnK6DUGBYYnRcmNCfm7x2A5yoepqDzN
H0+CRej7LYWmFYCsevu3h9HytYh/rKqxxUDQ6tmCnjB98lvCmgQQLmiG0BXtL/y7
TB++eh3K9bkthmUMfxqEFWYDl0nLDuuYhEkJm/KlN0DMtGwRD1Ox+ZmGTQqDRGOy
UUFEGy1jd2D2ZVqANzIPV6Sjpt0Vh47U4aRxlunSLA0ceRuq6nizty2puAm5cBwP
TCwQK4UroEmBSCXzHHJSNBwn2b66eN/1AvGoeDPP/LJ8rxuz6thi81vmhs0Wq4JE
e909duUzuJ/0B/Rb0qZNll9QUi0XUHi5U/K8WvVuTrlNMOvXvXKIgWcvo/uhqu9/
zrUC3BpiAQ0SXcdaan4C7am6AjVEJFP5y/ITWfn+qWqVf0Q0EqsE4Pi81yXTba7A
CMKpI2CU1iUxugXF0JjXHStd/odzpoZ1YvMfjLWq/vIYFu14XZ1DDxwQA5bW33uN
mHUMVRTaotikFo2Uf7o1gWOY8YFGoIXTOcTumbrGUhgTehtkCgPygA1akKR7FUBB
WFb+QRGAIJbVyw0A+EIpAfaMVlhf4B/G4jkBu+R3jnJ488kR2lLGCbHOewtWQBtn
jzqcyEzG5su12aBWz5x0VX/FKsaibzFzK34Rj9AaCALIbHxF6QUypWLHsPXhoUld
n2BqCfVUS+BbJEi7ZzbehCf3n1fPvZ9L/m1R+psinr45fDTd5nSUJh7HcLGGx5XN
xW6ahpSdZj3t3PBdtWI9U/86ZIBc/6GsvGJu4WuV5s+MYgXMgRqKNIgjRUZ4L3nI
YK+GJkPNh+tk3HihgD4ikU9VAqpNRBI5JD8yTH0ORM0FJeVnr1t1Klmo9nID0M8a
b1QGXbMIGb1mh4wRXvQXH2jL83SFZLgL2Gz/Y9OX3UeyVn2MgrhRdQ2xhaaqKMN1
1Mr+wtii2MAJfwsOZ6xV+K1I0LrUDnjE6IDmnrlVAmzEJbmucHaK6DPUxKhi5XNe
5BzYHs0B9BnWexC65zPEGMXpezR8h4Ujd3wbJWFHYR12LcGLXDxV1ZtWkxKZixMf
oTW60eIKI/tBa7tu3rml6m6XmvJjq/YxjvtY0fFG26xPoY5ZIWNQ52cN36TAOTsy
1q3VZ/XI8cVS4eKUjfZX8weRyLHM7dVYYFY4pKQfjNERjIsi0vIgXyL3VdI4UQwA
VyZnGN3EEfCk6IN2NqNy6F/gyMWHWvcwOLvkE/QwOETBFScPeVdrGM0FJ9D1FCs3
piYg6FUeGSm8Oah2M0iet/BPjyKLnEZD3KX4kQtwkHSlGOgYkemOMNI6N7tRH2Ax
IoNOYKfACWB9Ky5KBta7Qov48ZsKbrGYBWYFSQ66efsThqoJDXSlXwR/ca5cqkCa
27ezkBbKzr1V1Di88IAdncg/OLguXF4yWqWOEHezYT769hupLAKsqCQRIRQ3cS1+
GA1PxT6kAMu45h25PLnN33vPsXGAmmjPKE5R2jg2xLnWGekmzJVROS6R35UJbP9s
T/3zLWuGgwAkiV1SyGZOpdV84XDIBCIHjg3EiibFt6fLpCw/oCkiqEy8dYidN/Hp
ODzU+eB4+ONPoBBbxP26cEjsdXHwCpxTfd2gOkL5+uVVzaX9T2XDgu12BOJzpliA
8zwxh/pudsSXlWcomiBh+6Dm2q7YID6O1/KS5oHryhm5aw2lW4nTNjDHsDlcES91
qV4IfvyH4gb2D1LW0zHiZB82grMzxIP9u1TcObQLG1vD7wA6s0De5sNdBr9TEaHl
FIF6S4FxB2YOtn/daEQ877w8+o9rFgXG3xG6EkvuEwdH0btJUbs87+dh4oNvzpQk
7xGQvg4pxk/OGtE3TYPa4+WEwLWZYKNs5fkpN5/2IRNULXIeC79w7My4OL2cs42A
lyBdX8W+0YxEbwLoICHuKrxp5/xSXh9Esq0K+VUaLmzHj/+/tSLVVxjxMmHp+Nqy
o4cPXZagjYWMhEjIlE/G/ly2rorhqx5ZVE0mdEMrec6IKU3nzgRoGiZbnJN4/hYB
riYbKUl1z8IpfxpnhbBj/hL5W2E+H/OijoR4IS1Z3nxqnjFWV3f8B7CbVjY6s+3c
T6OfBFbBLsfOzZKjQ6z3lgQEnSMKfBsWeXtarwU0MoTKRqEGGCA0I6Cy7T8Pg+ld
IPalexy15C9sz7qKUVukSc8k3HICq6+hK68F3EwKJG1o8z7oY6pQAU2za6+fKK8Y
wi/LRPQtyUwd81aOqVL4OAL8GKSPPaxfmknaevO5QsYBssTYCxmE81wsayWHFQnz
iJTSDyWrEPnLWFPCcpJSmwLuhx2XztZCKIb7UW51Gb1QWToC4RuuHcDCi3n52ueo
FlrY26m39J2eTJyKiHUlv2CVCQzdHiCTBqQyjlrY/0bi7sgMkG4Upr3XMzEZeUdS
dnYmnynHVtK6IiGyALs7Lz0vIw/KaY5Ws5+FowrjOFrUFaIsK2WPfRSgEsu7CUZE
R+3Gej/n5kbfJecnRnKWUYMr+97/U6csv0dOBoULfn3qNsuGfMrL0eumKMlNQscK
G2JKRekgBd/Q4T6RqbhsCOSd8I53Gx37yZIepT3mJ4Hy1bJgGTWyD/3EpJSUNrSw
Nz+rb7MQPFSgK0kueUs/RVyEXZ8uKu7xS2Dro3WijcCXLoVphiPlSmaNSNo64ZFh
3F23s9/M0qTmk3d+Gix3FLUn2BkgOZtwJ+tuLGw2m1odjWQhtDhie9s1X6FUXlDc
WkDaGsVzc6J/kcHj4pbKL4ZjYnnIssWvdolGMZzv4l0Gztz0T47AhKFqS2Dv1ClW
C6eqAFz0Nw8CJa3/SpKUsfwfoHal9ny1PMOqojgAeOKPGXQ2R7FCbk5MFcIvR80k
6iupzBHncq+l20lMe0SlVj1xYDJfce5Nj2Asc7DMn5aBAPcpfmt4VdQddPMu+4XG
JKUsnSMRsKPtKnoujryhM4k9ENacqZL3cO89rf36zLgCVrZOL0aGfJqu96un1tTS
GcW2RALWzj9g1TkMUjCBAzey+FKPHdN3D3X7XkUAzebJhDgvr5AjJrgghEgASIRK
RX06vbQ6hOo+2zWfuqwkCmJEv7xaZgdBAMpWvoO+hhvEd8XtWVaWOM5Ioit084DI
mGlhwTHzkD2nxvJn/iBxPNyZEIVPs7w5p7q1Z/woyb6TdQDUORSmoWrcii4vVpso
np77h3QeM7vlqtYSzadJH6prx45AvYfSYa0vrY+ujslSGgquGf+DTjk9P/BTCjXd
1dYG/9SBi8Oz7izt8R4Uj2AMVj0uKNK3zxQ95BYJErdFi+xagDORc0dPJ6sFcxNb
OGnstsyQJia+ff+kRGfIed1zR0ugEHeN+4j9EGurmgbcOPyUk6aBaC82sB45BvJ7
hD6ngPCNi8Fp8woc8Lxu5oHwads8boEUVh40mVgHCe+A5Dr1gwFbOgGnDzU4eczD
eMXtUNUOmG1p0cjOwJpoVCJonG20iqlkLyygb+YEscQO0wo4BoXlKa3MIOF63ABk
4wh/7V6Ko6AtuROgljhc5BX2LScf6l/7GRhG1qUT9c57RsUm8DwnhFsY3UIf5du1
U1cIB0vPj23C5oQwRi5pDttjEM5QX2Q5eJNMmg72z6aoh5kbzbBLRKXnUbbSAlGt
wMwutX7aMI541dLwsm6OVzkT2/c73ZUkGEIyMVho2fwNhnDu0NuW/NNzdiq9OpID
xb2EW4a0CirtyF5vWhYV/ngwivU6Dpvd6/ly+EXqTBEUIjwgxLVHdAlFWYAsNIWn
fm+Tzjyus2jXdQzYxbw1wsKaqJ4n1xDtA9/26Q1RjYhD5Rbw0S7O/TlimTsAp+5Q
+GhiK+6/MTWJ3dEhFNPREKCYPZX8Ysu0qXy5l8jikeUB9ZKM+iMd2KkZcc6oSktr
tkNgRXRi4y95CxLo2ABmKEar2X7oZAEZIg4U6ooXJSxs7oOgY3icErgTR4uEqKTu
bsissoJ5ErkkyXFIKm8GNGVHr4ZPUnKFtZsjvc4IuOjdKn41bqY3cVb6pM5iWR9O
VYLW2HIf3j/svfoq9dur84ajxjcMfSNzZfsoHYwWj68PkzHfwLx3qOK6arPsZqpz
9zZGHC5wHR5vTZg73cSEpUAiAlwD9h72le1vBQWcstyQtow+wQ7vZnwTnEptpmek
VnFMblzw5lj36B+KhZCmxFBnCAXRB4y7ZP4ZRhizoSLmCMa9K3HtkczjWPdbrvwp
KBw0HXV76u706mlXT7xaLf34LP+NCR4PaublFf9UwKhA6ifv6fFXQYP3C9ZhjYPo
0ggPxuXMit2LnvZNFeRGj8/b2vUEJ+2GDHPsQ0fzZ6q6wjRgtIz0lfThUqVU82MV
Ob5yC2CfsI1nnCJWpRXanbXYpaR6euVeFW7FZhve+tBtpMc7DBgxv3kXMFNNQI9+
ZaealzIQlhvmtGVcbM/KF3M+X+QCcaHAxxTDqTHpY2+6yEtWCeuszYFvg4qolgqC
9WoOD0OrNV+VLjxvRANp751u78fDU2TfI8W23lDUyaZkSpUT0lQ6krYE4KoxLPG8
wY6ffFac6IxLeLw/1KopTiAfjxbEEtHnYL1/cXQ6UigaEzhtXNiuR5bHy7bjjxVf
HaV5TSMb7kmCqvC7zDX6FYmUjrv3iTxh9S8MJl2HvxmRyUHVNVvbIqc7JorA/P8b
ENTpy2mrQIJIBti0gzdtZSuheiiA5njoDc5aSUfB6kNSqzN0SJOTqAI7so4c0G+A
Hpr7mWb+UqSppcV+QOZwTMxYVdDecF4392le42fnvNySTMSd835q5WuF49t/apna
AeHa4WptIddYdAcNZe8F9pywcqqnc+6oVZhr92v8k2z7IFZmRcXl1j/2KFrUHW/o
tPB97EkWdyfAhkhz8CXkPyeP/l+YORTJ3qgwIRedbVoTVdVQX0jVSBAxLo25ZGUz
OCl8MCRulhVq2TfSy+z3akLhMmHt1xvSyDUNNIek7nKAUiLpRbv88oiILPeCo7yy
N3zgtvuZ9ACeM0ldevTxROn7Cr2wk/YsLl9Hxyd/OotoH9brI9HvHmIJeWl1urfm
lnrpVyU5yGdUaoKf10fqikPEID+2agXQH83rnAZaTVrQZ8sw7OdleuFVP5Hcu3nf
wBMa0j+QGSuYEIsOmp0uwGmx5bc4fIJ/fI6bt7C3iSvcOwt6xTQF/mJEkCv760lc
ee3LzyyQiWVwzYtIQHLtyMpv8NI1b0nV3cwFbVDBZNHs5JLDgH4QPTbgiDuxsJoL
r3ogZ4Vum2o7t+f+1s4s29E3CGTF7CROpyxxG4aVDUlmQsHunncllB0ePFRdKjx/
Ri94BSlvgCwe/Up4wigx2ePW0uIvUpcCbPzU+yfYZo333+GsSp8i9CMd33/DSzXF
xVOEwneBj32CxAW1mW2RJVxL52kNDq2eJUdUSC1Aip/1UYyHsfNuDw3XgULE2r17
UUM3LBIBI6Sd15Iy0msCulfp6mTz+JciVGTnpz+7iTHeXr/jpxdo7baoeGDLMU2T
mKDegTmu4sApd0CtA1ZN18IpHP1jy3SpkeN6j8VEMCxc53CnM0Oiz8RDrpbcOw35
aXQ9FqLp1E8EYXk3oO40T05seviendnOSQF47I7gDIMyDvMuAb7hCxyvdPE1Lnmw
aEaDMNTLNXeXxDkBHLSlOcp8XaCtQnPf98hTG1N69zmLK3oy6nFoDxxcHMUW2Okf
BxfMQzG5UWj016N0MnF28j+UM645ZwDHwsna5dchhdSnwtfRrfbtvwpZuP3YYQ5w
usFjtrVsvf6/wWq/hZGAh/fjFm0GbaHB7D/BsIeq0OEBMNtucNess94PTR+aMBw/
YaMW3yyv0ivnFiooi6ZGwfAF1r7o6Eki4mM/KvhrGpA3JJF+ori5bp+2B8zkf0dg
5UHlVMFLwVrcPcesSWcDwnP4pxJ72KYRX08n3zL3gPNkD2ZkRBK37JOF5hskXFSm
/Yhv+M90HEX/zoCO0Ofua3vKJLE4rXsF3Al+KnkOujaJrOn1BCn4zsa4tNRm9Yru
jmxZCLPZG8ioOHhTLpeQkaBtJxCapCJm+sAX8i7LV11MmyTEbE32RGR1rxwd3ac6
Nu+TbHGDbAMj3gufSOhCrkoZstAWpNWjGzFJtE5vxfZ4NrtiWKeLCnSDeBhkD+QK
XrRKRWX6QHH+knJZ42SH2d3er8OL+OXvGAg8pqRG02hQhbQAd6Iz6Q0ht/wpDtQu
VdAzbUHpVcIC3QyYQZp5SxxB+Gn0NYGhJebm3fGQ65Dfh2Kz4H6gU/xe8H87zt7H
XurwsOXXw87+WP6wpqNpDuW6ijEsQFRGvp3rIUJFF2+6z/dGaN/mxWhneNvhlRBK
9efqQHo9Ek6B4kxHvcz/XbM+juL62ge68GhoOjm8UGFDbCs40DE5gHzbCmCgkFUk
9JYtQqfVRRoJAeYjbaW/vCp7gJQii8GX9WEXEaZ/0OszMzfDzK0pxa+K4pkECkAi
1tUew3OSyMh0aKC6gzL2OQWpwxHcnCvygSyJbAGO++wdcEeKJVumCpSVwTd8mo2Y
cM3mwz2eisYdBY/cpRYyJN7CiToAc+IQ/J1qmh7Nn6hvKpl/p4a1lpqVzuBG3nnU
h7drnkMwqgbAuMSUKCqIP/39TybhBut1fYnhcUWfx5nihY1I5MTyZwd/vSq93wms
katA6Y0uCy8V1lOlNpMT5Fll5YD9gCbv0oZdH+vscl0ePc2SozJmLdIfz4E/q3fQ
apetirThI8y0Hwe+16TWtLLhwQns0VZ0/YJ7Mg9BA27ItUNN/e1SfKNt74ldsH8q
wKUtYBw1T93z8fJraO/VK5tV3LpfrLf21Zr5ivZ5wnO4/fRM26vpb6XPWEk0fTZE
pDMLuhFp/t+Mslt4oz9enrj5L1g57kl4Ybn4vrPU1GfMQ5+SGaumgiDyeChUE6SU
+7Ur4AJdbaLF890QnO//50DtW1xq4WvQrgsScVMpAIPzyGhXElxprUAwIljchmlf
FCie57gXpFHscjnsQp2OLihnz+a5MKSuJp1ebbZW21bzBmx5AxL+AhvagGgC6ent
ltHAsqcYAhKapPZwaAUmgVByssKsKxIlnPppOUh93PpkwpJB8W3W4ahx/qUqFDxj
rQJH+UtrtLgpWlNPkMH5Qe8hNSwOE2iahB3HnkTrl52R/9F5WxXZ5qcuVmK7Tl18
4+UIr/zkgc6KmFVKFRXfzubteuo6lDVJH/9zaIGkC2RPO2OlegSLuoI3WengZf4K
7UUH/9LpV7uMmSzQtcBjKfB1phmX55QZ0nEtXUSs9J1RS1lMymr2O17pk+WJUgHQ
bLzAcfgWurEtkQqlz/dZVjL2vn/OhXpKZXgsuGZNmvXzro/roRT1wLU8yxn3OZ8+
ytT2DIJ4dxDmsaIqRlikDQvnGJIO5BtIAptcLgkl6PEOcGREs6lAf+SdXnpdvfFy
lXcySf62xPCIQuhcQdfj7B5lksvEvfONrVtLTEX1gQH88VNQQ2TUljQksrwK0nZJ
QOK8optLjhD7uLJ/bKzscW0ddFkSNdACXD8V+h+hPYoPGRwSm4WFVgKL3Rl9IizZ
eYBp2DAlHcofB/Nh3uj6uHHDbK3lWzfM5/MlNHvKYaigZ7HuII/g0sP31pJ37nkO
Crh9TqAFr4fVoneHFfWHhfXwLlIAzH1rUg5EPPM+khibxsgbgfT4Cs9txwZb6Pen
hGgTWzvlWxXg/iP8QwrFPco4BpqmjLWsAOlf7AFEbXf0oolNzwhqPv/36JgU8EfF
UHhWxlyGTxNm0skvDKgSvwlVxDLV3DuBaPN35mRZ6zi319+Z1fRMySiBROTRQ2b2
h9pK4+CmpNBG81Rh4gRTfoj0b79Nxm1AodtL7post/7k8pog4CKVPP7gLWjRF7Ss
RuYtQ+CoYpAzGTjKHV6bSda68GjS8tInEpl3llyfdcFXqH05bpaN1Ix7xRA+iwGj
zRhBYcuxW/7xshQ3Hi2kgpZlpyL8R8kTtyy0YfRZ3hzr2kk76A9JbNJnaHT1942Q
2RfH5XHwDeBukzwiDFce48NF0XDnxY/KChInkGJdiuhkc4edzN4mu562cQyrQFCM
OqLTqvpvH1puP+VP2Jb24oIdOBrJbPeUiGiK+YxKONevKsU5c663adYFTGZdYnnq
AbT7fDslbd6RDe3ebp9HFEu3K3dPQPdYIHAZizDusy3yXsXwhdkjHS4fOSvAS3jx
6rjzvwetMJhBxHDxGLO7JbNan2Rwm45kV/tbb9He8Y+A+l8S8kOHgVxz2ik9CORe
Om30KLwNZuwqbQ4dStp3AbM9Ev1J24qkvySMo0QERbGZd/peFLS8T7TZwEppmIJf
j8BHCFo2cbGImtIkdAbkk70MdruhC+3sQpH4FpZcyGcxfZqYsmla0Q/fP/QacIR/
qCTg4OXh+t76HPIplo9t/GI9Mc0sje4BCjI8/L2mnzpyqOis1E719tI+48k7Vr7m
Z1VQUARiRSn7WHwCpVO42us82yGoDWEyXaRyFwDnZ1BsgNTtYjanF16QxDBCczLq
d0w2YLf62u0rMrzr3WjAE4oK+sfNCCgeaNSaWkQ0FGC70ARp/Dy/wooZ01WA6TcI
DGqLKn2ibgUL++mOg1Y10rhBBORBSPp9JFbxQmMZjmp9m/sEnM+Z2K19Ba0y5a2R
n4sdn9XxsPpQs4e+675k6MoR8o59UGACrvrW81RUhw0bf0B3fXym6saer3gCkK8t
xIHo9eBArO38XtsnRl7dnF64zDpNasISRg627kVt7YfkSBG1M9ex3vzOiMIFIMZJ
ZPNNTShBJTfEyPED9jrsBGoIfcjw54SHRuZzcIsGNjS8QxGUDQkDZ19oZE+v2uvj
YvknhWFtDfi6P4Tu09ONDgNmucaPVZL0U+vZGIfSZ3Vw42nKGH6Au4kfQvlsH9V+
64gIM9Txw0sZwOvxTdoUiAxwWg2ECKrTsVtyMGP93wLJPAgV+6WJh+Qv49qJ5j3t
5caFCXS1UK95eLTyWdt82cIk4hwlqdrptGGgcV4/nx67cIgrsDbFThpzOhX1irE8
PPOl1PW2siQ8Z0Qy0RcLBYyQSI0d3vPYvqi6HAnYaBy1yohBG/CvB+EXxj/viMPF
oHDZEF3E7c6/ymnm754ckx3lFplg/6SwkffEPaLVrq1dTKwXuEDSRT5mo7B7OcDi
Uh1sxeaNpK1V+4Ot+ZDXiuqjOTRYBLakSl/oy3rYIR5l6f8WfpoGzv0kM2cIr3Zp
I0xEfJAQdFFOB2EzgP9OWJ7spP2t7tWW4j8BSFmR88+9tmbLroe80mJ4CqLN/tCA
I0PwPt8l9MAZzrLKRavNbt0VB+7x590vBBTpCzZTzM8bjoNAdcTKbz7TDd+St9ES
epP1J8bA/G/qa0imPOVEO6+UbwrHiW3dxn4XA4QPQVOlPpU7FVVaDANDt8PvaVzN
ZXn6IsXM0S2svRx1QIrLTXxM/M3x/AjezAuhGp71ynobdeVddilvyrm5dowYRvrT
Z/aZOvMXSkIa4Paw20VisAWvW2iAL6tMb6UW7WlCUeUE40lWjenGNCTqZGTZRmur
8gPqD9o/ijcuk1A8HIEgj9cOaqUHB77XKNqNc7tuKA/6cVlkr5V15Ian9ZOv0zgx
R7DNotwAnfBglngbpprNpzC6GGejKhgmWzeUAGtrHJr4sOzR/xL92YTEIY/pZrhp
QzMfX6RSjUH0S1pWa/jAOUMhRaf3BdUrbALkNKqmU6arHUUduhXkJ3gjSSJfZoL9
wiGjyfzHTAn1aqSs6C2EFPqXEHNG9w2c+utBiv2LW7JKBumrg8WT1IVxc0P6i2e4
0lZkGlKZS2jdFVKSEkffFLLniBbwuiTVRrj3x6UiT8HW+qBMHA/wt2h5XjZ3zeTR
Nj99Xa/h4+cfeI5MC95Kw0YM4hiwB26WKY2xbvXVo9VN7gKIfJJjRRmBgnnrA8B9
28jrafO4OVeXdvMMs2eFYD17sJ5NLxTuARy8xK6g9KQtM611XVjEbNwSnmDx1iVX
z2/rVQEZ1EzOlD0Uj/D2b3IU3taQ95Kl+0gW7Y4FdFtRqOlWGGRc7nofCxYB2Vhm
wwyRL8OYVKlU89bGXfrleKlShkvcgr4Qmh5gLYxVYpw7QgIHNWRRHJbCuhmF23Lp
vHnLMnLBurBy/I2n7PkxvRA2npDQSN6H08VYeCtzR1Immw9t3KkT/iGuGpeUiICy
zNqL92yqN8yI0gFuT9h7xUX2WOjZZwtZerNjAjjOcW39Ysh8l3GbjelOmnmsM1Xt
nFJeishv05eR3BOziPBsqhJ9X0jnBsB9ccecN28wWCtLS6xeqMGytbts4/CUERPS
YNWZk9+oR7TcanN01hZW5sA5llypF+t2ASY4g1xFq8hYG2Lb2xm6GbA7IlpsGYk6
VhqKJNnxzsgNGNOvEKNBPJHOK/L06cJkx8dYMknHUR6THHxvE0ierfLyoLpoP2r9
2KNaeunE12vbDeUZvk1P5kri1DEkgKWxPqtsyvoRm02a5Mg4Ru3iciGhH4yEsCVP
hcYpp/2TBZPL+LrGjxYguO+0ga2pnBW0vT/xYiLReQaOAHHc8Uhhr6ThQCbLTywh
T3Iq3tqdL4Rr1T0OCPeDUzhNXnEBP+7lLvBqsLGpRQX6+yY+wt+0AFOt9OtOstbE
8p1+rHJR4SdvcPCzHQni7KiLciyMf0c4dp3M02cK6vGdYCyTSwY9Tt+zFHI/x4Zx
Jz/q8FS/LHTEQz+ItrbGoA/QRLA2trvzcSsD4yFrRynvRfuDWGLNI/JhwaRSWlKK
tHZMg5kJrRBdxYlRmXeQVx+37iP6bBXEBY7Mem7/axjGtoQdnhJeHsVqJDvuM3V5
xaeRCUYLdIjetZkRRk50o6+i8jX6pAHUrzXeXGaJM9hFDYiGusOZDwGrMzIVCbSA
Fi1jLeUcdqi1AJwlcLwCMkm0ech9ZQhZfsoL6ltGboGABH9x//YHpnA9J0+FHN7f
xievSlSX9wbWgujnINSVvq2TgrGEM+YXnaC8eU4yD0+BONjHKXc/SR8FYcn4uAmt
ueLtPbZbrs6WvVpmyqqAGWZ5b9znJkAYHb/ZwN46rhuPtiU6WOCbFMCSdk+pPVEJ
tGrTp8V/qIzYNkOGZY+Syik4dS5QlWnOAUu3cstJ64oN/jx7gVZCaaGL2jB6yM9Q
bNwz9GEbFRTwAc3/MQ3srgE/aEU0YbAzb7qTNiRaOse7z9tVZA5fjMaUHAEUOj6O
MEElkh8WcdhrbRyEK268HrcdrKH3CyoRohJqzbyF9E2FX7brX7E0UQYev0N4khLG
N9AAkxb4MlTbsWFOvjsoigkX7HOt6tEMjI6zxPCNExO21PBmqAy5pflla9APJhkr
pJ/Qy9ZWnXLZBfj1nzJ00SLUqMiEAd3ihyWQwfAVaGUbgbMSdnsBbDOTGgnHPqq3
w8FScv8mlXLldWhhWAXya9aUSCJVM4DHuTpubUrzhvWh6uV6qy7oinCAh+6sXIum
1uL1XGGeh+7JC3BpABFgTz7X5aBNlAAkP79uWMkadyXhbwyLh96MaNEYJeeLVavq
WHPSZS43iDapCyAH7Yo9g/7eruBLwctVjLIncdvk+9s5Jw/oUng7gmeHIN2TMJog
aCUdtr6W6t91INqmhYZwWTbs0BXbYDHa2K7WDwn+DDCm3ZpW4Cc3fyT+L7GKZ7r8
HsBQKT8KQ7z/sr21RI9iQBOm2N2/qGxvZxR2yo2gDLq5WMnm3fvq9QrqXViRSDe6
rymOaBd3WmlaOOLREXuvzoslW0B61JtBHeWODNOIJkvIsemQ7THyNkYNAIN2RHCx
bMLha3U2hGeRwEiKlNHGkQuelRhHAqeDLAUHFftawqysJvKM0W/G7PWMHgZY85RC
kSU9lz7d5TmvXtgXtaPPfazGQb+8B+VpQfA4WF5CP9lry3tzLswMKANUmfcAWS3G
uv2UQl4JdC3EI67joNa8MpOgLqxM5Fcvj6KmsoIUltVA4r5CmbERjeuCLc4WxSZH
n9o8wi3h1C+ZNS+8vEjCvRayLB9vn/NJhL5i+R4zpgysU+anLFco3yhgqQb6tCBx
Dnu5HFVBvpUuyietNCdSAky2MyR1JONUB9TmnTT+Ph3mK+I+/v+be79EvcmeDGn2
0SgUgFbX1hq+v1J939yxsMn0YAp9nF/B1d//1orSJC7TLZvSW4U/HNldWSEW6xd0
hqRryq41cNDG59kN2FQ0EORDBCtwFBNTDjujvB4F9ctPd4FfY94Adx6QY+BeP5/y
+ZjPIrs+Z97nzGn4DxRaQIHMkaqAL0LNN6zNEJYpAMFfDIqVbwj3P+4YEEVSPcZP
JHf4cNmg/y51AsJpCivUlyHqkAE0TOC966T7JdIsKwFSL0pH/GqtXE+UI5P+jQZ8
nWotlr/nPrTfpMdVaIJFEuWuYC64wlz5L/9i+eDsXcjnTuXR5PBGXYUQOcwIfGIt
yByP9GVWqV6tiTuAlApV4I8sL2VcV7/SWklBkcCfjwZVPNtHF/h+OYPbeVgLsig6
u/aOTsuJpfudoAXnHRViNfhjuTI9l8VvKASMhyFPZsH5AWV4H+M64xCFv/6SvB7v
/1dV9SX45qgW0cevlSoghqJkbqI7Gg6S3ZyVcZ+wqj/9tq/oCv6BmbZ98FJzNgxZ
qdxKToa4UQ1QEUmjPJcrzqcaJpd+4KHyTunZzRGjVRoqsBFCuG1ntXEpMeQUsGQ0
rJfmc5RNIJOku2zgWlhK8vdtpxlJmEPkQZNyzDT1Nix2kIt7m9RN9BAiWtE8+u5h
M7FSYM3YElYBUUI4lxg3gOw4RTh1PbjeVGWSE67NBNRmCGWf6TwjEbd89lGkw2QM
3cpSqYmAz8+5G3zxJ2qUgX1W7iVSVLCYM48Mf6deFRJfyki81zEYtlIy0+Z5rXEW
JhBX98UQNCue01P2ec8pyEMp43DjPo0y7dqOmvBHuXGzH23J+EUJANpKWRD0IbBF
G/Z4zB9RW3Uosz7czzY8ScyXGIjp4C6FsjNLSWn/7u/0xgvJ6Mom7YwJBVSImWJ6
/WRchlkq4rA8Tj3KoeGZoKC7cetwIM/xWzugW2qZPQBJDj5sC42mwhGMSaZ3V08Q
c5mYHnQidEGMdd2/0xPzJX9H6IujvrHMbim9GSUjOsYfNOayX3Cyl/ijtFhY9q21
VNIOhW0/BhxmYzLpSNpnTE3S3rHswRoskmLkShML+xqgDreFSDLiB/bYJKsYDkZQ
kEkz12lciqbvZBO1MyhYl+S+VKgijeeK5VcAfUoUMy5hj35Rviy41u98aquo5m6a
Pzk3eKmsrhZpob8c+bBxl6F99YXgExDkeaerisNqkn4WuV/u7ZBnlf9+b2E6hybg
eYXyIhqIpS1s2wjE+XAOI4ju+bIho2SxNEYNQ4/ygBZcrhn0HRtq/d+WUT1a7w1E
bgdYjSMoccNIEVcETRXr6/c7iZWNWHFIDDMjpgogNj9Gc8zJLK1okivPTjSfzVgj
o1zRkYWmbDRPvFXwtI3M2DpzuyDBydXT1zQu6pgSHA8YPzRkpztuMHMKepgX+NsG
R4ey7YqxlmH/wmz2W5v4TZUelJ71xgPR1NeUOpJOTU2pNUgZ1VqxV5alQnU6UWdc
9WxyxG44lsNcTTJammu7UvbLTzULCRxLVU2OCcgdu34LDDNcQKmi2XEvoeH1AAAS
Ixx9zaoQ+0A1kH4GkFryVvpywu0HVZgpHe8Nek2d/O798F81KS5g6TZ+qNA7nQ6K
L+F4iUYDR/rXToUkVfRiUeL1X1L5PDPEIHmQhQNz0dGR026ygcW54fiP87+o20Wt
XAWUheVPc3tbZutHYWUm4Kr+E0dNws46pvw21C7Fu3EkIlEH/KDeX8VTGTPbkiYk
qA09QWt/r2glVxE2miYtJZnjqWAyNcbng0SAiuOcpQ1J5hgV1G6cIABmM1+wZefi
+4lBLkXxVqyax5DRM6ZIxU7qS1F8G/pnl87wpQYjn57DPIn5GBsqU9YXzvxcWn+h
Zyqi+aplAzGwXJ6pyf4QohEgVPJuA/iwb3eY435QWFlZfEE50cTbP4WcB++3uSHH
7uGZZRk4V40BulYusiy7Rr9JQM/babKvSK6sNS9+fUQweSevpfmFp9XjlewNr9s7
fDOZAJ3XkGUnIVvwTFMvAvtjxYeWaMBZtjmKnlRFsTsK+IjUX+EcxaQsDILemfQ0
ZM60p/7YLRC2GOJfUfgDXIkmVnq+wT3hXcXLvRXyne6wtTJn5qd3b42zcgl9NKhT
jQQ+L3YaGGMyHVU+IlKwMO6jrv/bhg8k3jHz1kLgRfCSIdxxeJ2RClrboEJcxf96
P7Vqm+4nl2zD47gQjby25LRAW0P769AexPNMmdX0LUffECkqKLb8auU5SJAlVD4r
JZcQmkEdmAgif+vfARBO/XR8akxfQTuhRq5BgVOchZS2Qz1RUvLvSKRhqPHBoyVk
gGP/0dX71PAM7jWJVAp8q4e4oUCR3hQMyhGQhBSTiiNd1pqqvjQ8E57JjP1CoObt
AVl0BLnl8lq9XtpbbFZP4TtRxYBckg16KpQ/jcLqoOjk5NYo1DHYRDqoA61w4xPW
d26yPgzcBk2YRChfHlsRiGYfyDb30tYCJc3iGSxYQ161Q28Fww78F7IoTi1B8f2Q
e47i+HkxQwQhqTNlahrmxXWmrgzlx6c2iVdLYVO85rucqdOlDYFCMgvsDZg6rrDc
l22Y+n1QzL+T0bwKo8qpSdA6AE9GECTjZmP8zH8rlhd3T9GeVH4ijuCz6DHlfSVm
/ScrKmynFf+fmmZ4go2tbC1ofaXt3czp74zO3pXo5Q5zIq5VjTCcbwE7bCCTUE1+
PYIZG8GMk9bdUq+8N3lYK61AQvFVdeB1/5Xt1SiWhwc5EWXGtdiuS8/JJ7VeH/ka
ujs8LidgU7QarMWr8zadSiDDe9a0NKMwXDiEEiH3cvfZzZEX565HV2E4Gko4AMpZ
SBLRQyXiJZI6CEjSsk3fIZ24th97qERuhDO3Ttc9nhIxYJZce5/jnSS0D04K9owJ
+04quNgVHDvXCh6TaK0oksVzB93uDR9f4LNlPDFtzrMY+Hosj8ncmS6M5BGJojHN
YuLK39xwrq8+z3LK2pEj9ZS4oKBIuq5/gojSFitz3EjYIt/kj0RH8QsfXpa1iNLX
HrvgfP1ICAJ5tX85lj7gaKaYUp7zcIFaafR/ln0CQYfo8HcPFGSIebTRslnBbUs3
AOW2Ser5j+NEkH0/RVvE0gbDGPqsCIb8/P814x1KFXWXeBBZ14Aj7vy5qTreZdcE
mtDt44Mc+L5OaFVWVG2aJrjL2tZK2dqkPp0PCkK23CE65tI2tCuHJq6mjw6rWnMf
R+3nVUablwucF44d2Y8rKc8p9FNeo1sdm+m7UaNUTOJVn1/GjeAIc9U+H6PKkPta
Wx0basupx2hjzAjvIN6/5DMIC44nkNCrRcrpcYk/ewjG69Cd3oCm1it7VAafmipS
tvLnMzzS9hXBOi+wThJoX6oyWHiV0XN0GSMzYbNwTSG6cDLbO2V9LI1wsrLKlNAW
zvddUMsPONOUzJIlMxDaa8o4WMvF9JLyL4XtukAFBnEWlUYDlG2fYQbXtC1rA0oE
MiG84YEAQREsmHanX2L7Bfkb+VDhH9hv3dUTaG1NCfHK17nfsdYl+6l3w9oFOG24
Ei0zQulTSOeUHbZUgXaDpWr3prEvsDWXMeGMUEjjxGbTL8DOHq1R23nK+fPgKvGG
33ztBR7Jzz46S24Gd9Fr3uOOT0rsWrZ8jrE85ZJEn8h7ggJFrdLWuITgsxkbiHHt
m4bNHVKpuhsw6ZOnD7V/ALkgRNvk02xBez4/ehwlnS0lQhmQAEhDrp631QEgEcn5
6qfP/4/3vIOhQ7/MGLaTMHCaJcutkWIcGbiSEgiSwJtnutzNIj3nIvsGjDhlVKza
RYkDR6QZksWLLYNyFxRzfKPeK1nBpI59rkMiXwF4MGSSDjxjzuPpyJzezK5hf2nH
cdmHtXSjdum5QwXKo3/FE2sSks77j2OgdKrw7ypE8Pz59WZiXvl+mxJamZVfFk03
kGTrsWYLAbp8L989uRTgdKWmmeG/RVk0FK24jXeaa8L6jVDoJEbsAbUauCiugiWu
dezRarw5hHcyCSfboyIT25CevyZ0I8vOtD1e2rsdHrgpPpFVNuYtB23fuwPjN/7n
709LjHEP60MpKCIOz/61t7PHfIT1nng7xMxa90h0RTPtxbTQ87SV+P+4ca6nQ8DP
qykbKQ17rMBbY9c5GnPeuYufsR2KeKoaDSubCoRRlPTnEdS3dC/pGv7bloZcAZl0
ofqs1ho+GQV//QSTGRLBncTORobQE8mXApfoeTMc6YzgOrWzrckvdpPxaRBC1TXY
i4c/+U/olHtywjzcSIt3ACOKJ8wOoevC7vEZNJAsm+m7uwG4JPfPqZn2zqAVAYBb
5BNMCtxSOUg0oZaEZ2EBQpwgeCGQAtEfrnDUvfAnQOWuJofrpQdQA2eZxfUXfQ0c
uUXzgc5oezjG7RKBWrpXLiu3cb8dg8xqm5QiXEPHSTThRTEGYCVAGGxY0ec3/Jip
33v/x236eWIZVABtNHgSW3S3quq7jOpMokF+sKQieQaSKG8TiWFslkOw1Q/j5sl1
b0PzTQYAvN+YOXsgVR4LhiHPC6EbChCQyp+1ztFUUlNBWJYQVUUQwgmQjUHAD1F8
CGEZ+faWj0kLlQ+M0Z1e3Nb76GKb/Jc73/6vzSVYUJiNtglB/TNm1EkZj3JEbAyq
bj7IUAUdyxj+inSy805tifun5YTgLOm+J5W0A9i32OOVdwL8AL/h0R3/4WDtC0pD
mN160Zn781aI3daKVEjc2Rr03fX0RIS/0uvxbuWXTd5NwMYaqEDelw/LtSnrcXiQ
ECnSl84fU/tGTw0B7HwTE4EF/Ky6wz9yzHcbnsmSz31B/Ede2kzrP08JjGTQGjkv
1ot+zr8Fw94KxAsNBKoaNWh6ruIeADg3wNJs8Bjkgl5qcMsqGWE5rzRskE1TjuS9
vNTWV02BCvaj9MzrXe+ZIMAsRB9QehriaJzErsrtKiHkid40IJQltcE5tDtoyvN4
Q0dAESSnZ5gtk8JvU2UICr7ME7sIVER53aF226t83t6/s/qhVzVMshgoOhgQASXV
kJ94rkrGshNqgVuXs9ixnVSpk0BX/11DO02ytJi0sxkTb4YMGv8JBV2j1v1rX0jZ
utL7fOAfvSr3gL8wtd3ViQIeky0nM+dRvrvO2ncrWeq+NPvCWKFoSIyauPKlp324
4ZZcn6dryPgF+TKiaZhOg+rlssogWKrTIocSdgPgNNLUuVMypUQ05BNNRJ5Ex2+x
Zf3Lrn57Rgmp4JGjMbCmHThNxzpwCLG1JOmS6hNnOw0ImWtQ55KezxoyXMnKUNFX
jHQt+m+G2x0yXWBhw6IWOndEeYFnsTnaWM2OCQTHK0tMCzze5/v2tFnf5pmt4dee
Aq5KW0vowwaLbRTig3UHrJ1fTYh/yTIC6UiqalJld1jQi7Z4nZAxSETVRXhAJi/p
8F3axNW9gSyO27YJme+qDRwfqeq9WiRjLj5zKqBSp+g4kH1DfICimfWBL4YnnOwT
2C5+9r1kBeumsqQMBpvZEVKio82Tz6BZr0w7ej1sPWUvIrtiwxCKVB2e3AOC9daZ
byQW18koojvhFT8KPQbGZhbXct6M8DjQgJ15kDqZ6vS8T1dclW9+AKHADV8ITw3q
tHNPmRynqBDIU+n8gQDtPQY9LaodV8fnq30uwnQxHXl1pvbl5SfKFtOv1CdkXZjC
UZ/mBiyrTwMtZM/ho68jBPfhrLtzf8525byJaBQ89O+A5SLx/4gIGqT5uEARXaW8
TUo4Meb43kC6PrdAVaZJatWw+0d2xApxqRkxwFvS3GxAowXJkTBKYSkJok/YwaDB
FAknsxjewRMtRaUzUJOPLzx57dykcGyz0JxEeQ0rQUtoNiYBOgOc51fbKVPISGSH
EILizgxqOql7Tra9CaWpTaO5mr4+d67P4kmmppUak3CXEw1n0hss01F2l9b9xRlO
sG1/Ge9BWE6WtVI2ihSxQXtRIu/iN+l5z+JgVENrNFj1CZJ2YgtyiQh4Inp1fVdS
FO1y+jzqK5Lhv5dYeWCiF+aq5ILag1FCGfRexMdPhTHWemojXmU01q9Hh6fWKo1q
sE48wnbFXZej0WSCsFIOeOLY/r7lVQR1ug5VO4mzulbe5WOCZZvxjKM9FHzrFC88
/HNc8WFYlW2iWr6EFe+Qs7fqyGfdWnn+hTaGCrPeT7jFG2/2vVNh7TMJ76BnKv5v
y2wJVbnaOK80RTTh0Q1mavwyeJnp4Ql2yU/ieSypXN3KR5f6fynPK+zcuwkw70I1
ssBDFppXKyhaDRv/EgpFaUYfXbNuJKKqL6cnkIHJ8g1Rc2Gb/AgXv6XZWAtwKOI6
alyNSfDMSrL3zRtPRuJoNwBoQlDzd84VHgZlsyl6L6VvIz2vtK6q7aN4VsUeFcP8
nGHXl+tsRWCI4hR6bYSQnC+VKZK8B1MjdgtA7ysCALJgZj4lezy7Fs3U5eLwPE/4
lyR3S9rBaNSlBLPeMTHTwmewz2TfCc8ETH7swSGgVflXfIsN0yRfLpNOLJosVYmQ
7fwb09VowNTIRuVSECPlqiSWvMLCG8Edq+f2/elit/qWGUdB4dJrXIqIZDitI3d5
SPqGv/t8Evcu/VSC6XqeMKbJ64/Jr/SYGown9XWb8ue/xO6S0skWvjrqI72LqaAu
wKua+LaxE1kN66fDnNgJi9CMLdssaBjzd6aCErRkmD/OswxWUmOwhVUU0b5c8HlZ
f3RPJvGJ4aw2SWyR98CFDR1AItWB2kTmR0lEYQngjo66AUO70So+j58MX2eU7guB
THsGpyC26zM0vgxycHolJkybUZvxV+ayRYJfODIfTQj9cwV/nJMFpZiBU4TOPFgQ
vJyV1szKYM99vOjVUjVyT3LCDMo6Nhg33NPqOmXLQp/k0Kyjrk3ughKdeF9P6jOa
Ai27PZtIy7gbgG8sPDtuiUFqR+kgLs+64E+ZS4Jo9r4s/ia7rGF1goYG/Zg+Ejia
bv0WKP2PzcjEwolF17+hpz85Xe7X7EwenOYnJl4QVdHvmatuQpBn6ngXRWSQ2+sg
0b/Q8OE7jMrNHsvBiszf/k5VysJ08Akne+YlAid00oEkSYnTUiRDf9UpdAq5INYG
MMv250TlntfDmiD2OHWAVwQ4Zs5n6ggxr6EZQutiuO/40rTjfN5aLA3RBjo6jvZN
fF5a0rBN1iaqnfnU1IhxONtGiEw2UUaDBHOOFVUs/QhLWRgYlwvPiDkRoWMqjYBk
vOkV5HBQbK2cWodYX74HjQb63xQoBRdnSuDun0pTXtsPKGFwwNsm+8lryU1zWMo8
/JzKZNtKX+3ML2YkC9lxyKVeRX87FFPZSmJGCCaQ5KDkOUb6mBxPZwnoFwfQVSzJ
+Ls4PJJr1awDvmhtZf1nnIjelrvDPT1kXGQnqMIjZ6kBwiZgXrnV3Rxk9/fbG9Yy
27c77nQlLLOGpW4w3uf1GSSa4AHYV4BKSnOF8zz0r0zlcj/UkarVfSq52INXz8jR
VcQ+MCWyWq2x6uGDPJYp+d7Y8N0o71IsJCgG+5b66591vJa9DUAO0GQHYdsFwwl5
VxG/jDdS6d+n12rkIDBnjxpErJGWf3nIiAkNM49katWbr4CTAg9/7yIOGNUc+U9D
24R9pYLd1Kc1/BMQp3K0j6WMwlHnrVvDqJTsK/KUdNm3u6Wubxf6au/qm9+giLTd
F19CCuudbXUhnRVuW8kmGcIIOpMRkrnsS+N4SE1nQqXi+jmPnNauscIF4IgcXs3h
YG2cDEuz2qM+/o4LdrEb7l3Bb676itAQ6FZT8/QFMPCRKYXS6p9SVLo0J88j1C7f
Tn4XfSRhPHs8LlBsdysFi1cKjo0mmMsOmJ5ilmpiSIAcKmGFX7dE7NzeQlyumFvN
n2NPPbZZBbwxs0FrD1vo+K5DdidJSjdTvudYa7021LHcpH4gISOD3HsB7X6CFuE1
A6nYCSWCnzk/Coy21I0TB5muDrkVu4krwipVG3rbMncSGE95WNkNIrFOzWbuGEd6
fdSf4Po71UdRA8ibP3RAGxKjo4TVMvGGOpfmaGC1s1X7crSdGZeIOB44SUNAK8j8
TGO+bgzchrseWc9RExTuK17dQi2lbfSBbF5zB1r7btVu9DkSmEKe4JXsep0JZgU3
ncwewUGuiurJdwFEfdKzKoKPJ7Um+br6OjxBF6xUxfNMCqJjrTNIsHvYrHXhBOSL
wdD5/ANEvNDn6an+Ie2v683vvt/AyRZKD0jRPDqlBMP2XtUkZ1hwVtyVjw9fn1zc
XwaYaXU/qlxUdIV0hFgwRE/hYMy4VEOVwCKJt4ZhoowaF0x0hxQssXqvxPjLuad8
b54/z+BiU75VP0RLuLjC6pnSLEOEkAslOhtrMrQR21xeJ3USNeyZcL+dLG7176vs
4VIbicy4X0Pid1VmPxCHCjW8ZyXfKkYc97BAPGqjFGhuw/c3j+MLMqSdUWBimqEr
bVz7hw0FUvYsNsqgcs4xW0HWUjinREhMTY4WC0VfLRGigqV0LfZXU4Xcevt8OqCH
LvjFPA6AKt/iZXVikE0YQjrjwozvmjPQaMHyTIaeDnq+fobs5H7kq+H+xQ3DDxq9
aXRo8VtpgsRQ8BrgqhwAnIN6obWQxVuOgFcxpQFEvtGcehwFkgfbuNdrZLBX4hOD
iZtBThzzy/YEblsWjrjczHzYM1RhaAFQrwQK2JmL0XJ/NVXojeQP7/BS+fzZFLNP
mReR/pMYdyv12WaperKPpzFry9W0sMbPAkDsUqasFHygEdm6/g/Fz+TqnuQM52WD
pr4yq5IANapjjLQg72GMfUX8oo+M134Qh+U7My1ja4vSZh2hWKmWFczwl5ijFKvI
BNoFdS37eagNl3d99Jquwq1FjQci19rc/MGjJsckifu4pTWKvaOUy3TC2AwJlY7h
dvrXEWKVQsx1Jqvu3L7kAnYpWqoCmU4EyST0j6yqAMmeHXLxWJ/ianB5ck8PzSK0
3GTqqr1dllIgfXUK+Trc36TE4gZjY5q0rTCd9TBNyZ6aVwZCqgz3JKy8UN4FKgAW
UfMOfprRRGBDsl01oqG5OF2uxXWVCsJEdo9EiM/LWL7jZPjxoGZPxcomiHdGZ/VN
J0p41SxHN8mRxj7kipgaIm76XNI3sQ/3FoGN/aLiJLG2se82Sobke9gcPdX75UaE
594F5FEzXslBy56C6oRDAgVspLF1PjhR8i6J7Esw55ynIaG86XxVSarb35dUGzq0
+oHORtKG59TjG4N4qUT5DtNCqZ71MN3a9u2BF4F8/vbRehxo6dqH5gTwNWEizkN9
WKl/UdZuNpOK1LjF5B4oV9QX7Z/vEQuFqIYqd6WZxISfSxQ2ETG6h9bEF4PZLzGG
CRbh3+6JUQEcQtIV/KkcBWq36EI67PSHSuPFwlc9o1KvMcN/hVT4OIcSoIVvhnNL
RHYPvVtUrhaOWhMZQdT8Ypqx5Xx8acMkC0lhblNsRCodbme1j8YAlu1eRqkERCnA
35joIQE+pJsHcC18miQqdjiO8yXwukCJZTrUO9P7NgdxBe7+1ySHyKqpX5klyufG
RX/2booyt2J9vNXR5lT74PbMq3bRzbxh9rVEZhMop6aAG7OZMq6+EWEjGIszXcPd
YcekiYz33qEou8//ZU+2GYMKsjB3gN0riymekn5ny+9Nlx7K7wS2tOQXyaZIUTO7
UTjqy5zAPQmbJ7H88xGmsafMJuL4xS7TYUZCSwIxAQc8A3NmHqxdne7JUjp5AxcA
MaiaqGOVWmKT/DwbdJ7qfXDpgeMRtOduLg8EGzO/YUx5ANaFxQXF1LKhHCryXPAF
Dizg60XxtS3gXrY3rawnLPS46dYbFyCXWVuoscWYUtdGme4H+xCi/jmTyLeDFA5j
qi92XbE//2/YD0t4/7YijMJ3Wvf594bQgdHLWw1/aaoPS7u6XECcUyClUcfNsGvL
2EhjsqArBO6PTvo1vOO23CcqQgzAj4+cjTNceM4HW8GZxS0sVM3HQ1ciUG5ZRjnG
Kdjz1u/ZOR1kGbNYr71xj7hFZZgg6vMjIk0ueshevxEYsIkCPqold/7029Gb9gNN
YA96+6wbbVNtrZ4t5S+j3yfFXilxuz9gdDcb26w2rGUeyuXdLUNvMUksDU715YA5
723v7/fDiH7A8NiAMZY+BqUDWQ0dKLVTVVl9hJUyA9VxTVqpsZKAb+Lm9SLnqhNb
dqA0YocCzo7won0d7rESqJimCyWc3zOUzzs8Lw+tdMsrWBBvk7+CjUHgLHcI82vB
WoWhEH3dkj+DD3ccyb/y0MO02IAF4H9twwjQuNIZx+DRpGw1cB+pqFW+wu6Ni61I
zWITTSYqSgZ5Y1GhWOUL34os8IC9dBL6Sr9TyqjaIJQ4514ZpSnl4t0NP47cpgDJ
jluFrIt0qtL8zgKMGdlbAPxQ94UkTrydQu6qMRBfbrFJA3/YP2NGvKPgymTmSlJQ
Ukq+14s5XNuJHshPHyr4jmBegPoQ0IBMTDnTrRtBHu5wE3OSO0la9/VHvsiZHwP8
hesARirA7xYUPS5yMTc9AnCDQpHIhV4wQDIn3rkuoOGbpDD9nuVd2PjB7IpOeeWa
jjhMqv4b1lmZym5nUsrA4rVOhdBQsqSfdNys1onuXQIz7EKrmRPyzVTzmWskumEx
K6pm9zxA2uEmvvv9xkZ6kRfTSaVbnvDTJFWQMY/yz+ReSpGFg+dHzbSntEDB6666
n0E/GNgXCGzOdO78GrcF6AxB6VEnI6CUq67rCLc+uzoZTEbOHPVKGyEqLXurlW1s
glxUKXzLiY5C9SESGoDXLXpR8T5tak4Yt/4xfnop8XlGori4h1bWbz/2PrWGFWTM
gidf3LeGY7vb20Mj9O9MaQg6p2kfnEdXGxS44UOAF+bp3lVxi90ISdto68tJfa2C
ekuLJ7TiQ37K+d8sZuedTTJiohHImnf9xGqZNc9nC/VPMLCY+21ikuuwQZTAx7aZ
4h4833/iPBTl4KtP+MWUb6sz6jH63bclrKr09Ly7MucEBKLOg2smjp6vIy2Hv755
9AgZJ3KkqVffMsg5PJlCfr2Klj8fLAIxdo5AYOmgS8sZ2LsGklleu+smXWGctnT5
37afDOyjF6Rg7SzzY11lG7sZFUnfXKxnYX5d82msEqTlllUdbRkYMXfcd5ZZQ6JT
YirujnpFSW3qYjX+tOZTHehHxlKZzv0j9pFhKuCKQcMmQJoWYzhsbHTUT5JeBAsk
pWsscqH4a+uuKPz9e66pTNWFxJ+m4Ujl6D18qSWVCWXWXhNPR+OraaaudCEa59zQ
Id8u8Ux7Z39hDJV3pgCm1ss5nBlyCtHhWONm2oXT6yjuvjZQVgnIhTg10fLyHZWe
ZbAtOgUUX8ES2oBMAi/eXENTPSfMqybGGqoZ/vtMaoXSvXF+mODD8ZaiuXqGs0Id
QyHrmptYy1BYQAd78EVhI8SGmvIZubQgthAa3VaMzKC8PW3ed6s/CYTaapw/ScAD
m/BUiaZCSUnIRJTvXqep2Wl21LOncJz4gIRnLJiwPqzCf7OD7Yad9J/1hI+o7CMH
NKhZ9bB0ElKLPRrPygm/BDmr8qWthZegGybAb/pIhLs2upQRdpxQGt55kXXaf8PA
BZP6ImyZblcPa+9SDbmZKq/yZoRDzNjr5KxZi/3G0SOUfQJjWwbjmzLWA5KRC/5A
2e845mgqSn8I9paf/PdHFKPB1qUXZb3dX5cdK6jVtUQ6MwlkLElvz/PN6vk4gUtZ
XclljEWIfM4W7QTqeMbie52X0chSmxYffVCiZgXK0gSL4h15Pm8qbPV2xZ04g6/z
wvfXSe1yPUYeOqa5l48jaieVam2RV2uRdluTc4aF3zv4BTpneJyaB84+YB8ibTzZ
8ftw7dh52vKlWB+wvBtOj/k2ZO/LKezOt1PgM497dkKKMnVfReOVrROi3vOPlYQz
XefK8eyJ6ytPNW1lXTvzbkFG+FTu4DlwNuUfi0xEqrRr9nR/1xs9V3DknLZVqeJs
4bEmR8FyFD4X/gy/+1WVAKjn/0bdZajIcwPu8MWvl5QxwGdfZkHQFJ3vaBkxovia
NSlp+buvIiyOFmj4Vco6kJeON7OZHNBvwWr8x8uOB4vhCWgrnceUcYekTFOWDJ7t
6NmZDxEPtoRVdfcVei0BMaZf/hgCPVikIDvxYthftRy/waeH+5bwt9E2HL75+qyC
p3XP6IRA29gwONbVLMWXrQUZRRxL9ojROmGsYZNmacbZ+U8LHpfR1Wk+dUBbn65m
gebx+xpe1Rg9XYotwnPosUE2L3IJClHPFwlDAH+AlI2xTrbs75/C+mKBP7r6rtEC
HWnxqSnBHjysw9w29Q/NiTUBWrRnDD+e0yX6y9h0rf/zBa1RPoYVzpZWMEaQ+D28
OzWPxC0Jt1ibU+imXDi94DntuNI9ZMb1rtNA+JIQnzjmW6+0I9jZPHkdJCHJAh9S
b7PbG6lTfCOB6nvimSM+HlGGDBOXzBWJGkwxse3OsCovoOdn7arc8aC1vEcDmSmK
64vAoPm0Jp9rpGcz9IMvdMApGsBgF6U7B83E9zouTtG0P3NoUICWj3eVIgqMGAEH
OnTBI9lW0DrqhEP8vu02tQX1CZSvFzDDT6s86qNBiR4wE+xqJN8IN0mw4Etbxm3e
uolWzoRy9aBXvKkAabOZHVnL2+4a6paCZYPO4P5SSJuadhVdgbRdagTIliVfBMx6
tEsH47RUrH6snzIxhwUQq0Tw5W3hCTgsXZZJq3Eu+7ZQB6ExgcQ1Bwiwt5W1PBH6
XroKkZWFRrgj+IIahVhyevz8gdKtBPfpthHIr2lgz493r6QkP5HSV+0bYJFuZeT5
SihvKxEf5g+qkBQpBfJcqnZupDB0x7UIpB/nage2QRzBu2yLAxwXYcxvH7F9cnPl
F1M0R9EZtwcxSqODaOXAdW8BOC4TjDpswY+jQGNDOPlOH8DiXYIcAmIDGqDdkPy/
1eibOhahl0eDt5WbCnz0Vxs4ckO3n3vS1huYC9LwEhxOOWDcC1tmILx61u9WANd5
7rWFNAXH4dQCjK9T+0bqo0ZZBi2VWkzaDsilc0DkOl/na2QSKqWi9jBZjQ5UD4pL
8NBC0WibnNeA/i42wTqwewLtLq8eym/FaAsrtwKAndLvQyl7jnVaHVksjj2ESKtA
oM6j25Wjg0mrFjeTEx3jJ33p2vdsE878N7MzfMecfJmifSANg0QkXa5WUVBPgsGp
k3TjO4vKbfx+oOvQ34QP13TEznDq3nqojOY4CDKnIkf0z21o2gqVUuUIcYfhKwUu
SaffECDJ2Oab9c9yoABw8O+Q8xpn8VoLLUTtKITGzJfNZvblwXUxyLIC3bht31I3
GRdx3JGNoiDMsgjgHuxwFJuo9CyIKg7jL6F9IhqrtSzhU8vijnfLLKn53QnqOsdC
7MPURlBhOMFm9EHH1/Jjaq1F1LNeVxfVxeMKqRjwrM6zW7U2jfFTxqBiDoDf1R8V
QrfE9TR/ibJnnkpjsc7DNtGQZj5v5Uw/OSfS1w6Dv6+uqguu9k9o1WoRQ/pbTL2U
2CaQYNE7bmBIiI1JYUcFgMuCC5cH5siQI+8tzt6ggeys85/hvsVxQ7gCI3K5HPkp
63eXPEwK09oQV0mgk2WDHi5q8A6OcCZaMQk6AVrc8ycvQ/dqCGMlxmk2/apHesks
QhG567yr4esilyQcr0RvyO1ygC7TjugvVGM42iCxUwROThOgF468l9LMrFcN7cpn
PlNZl+eLg/bNhXAlboAwKH6HWbR9VyxDMFo31TdMnxYqN9+5gyASRQ1KoYC65W6C
XJj7A8eCH5OfhqsBoe0hhJ/qC4JNJdIV3aCWYChQ01fSAUh+uvmm8p70rqzhYmFz
str4bEinhFw4ijdajwM7bEIDo0EW5oHuLZAT5yeiP90z7ov0SwdpduTLyp+rfsbA
pAp3LbaHfZhYMIiaOFlTw6+OZarCR9dmQP4s3/KhTxsm1/fvxAlArJKw7NV22yxr
suEQVDmiJ75FcgJE6fhNpgLnLF59nvqdxfVXKHTpQqtA/RzSd4eiTx1OdFvxXXOz
uDXM8asRAWk3iTWufD7hRn3AHmBdBRCBS9vbbKd9jsLUQAcUlWPJCMijssku6ER1
xUnomxlE8RVFqgShKoQKoVyzokXenkGRm/D+4sGnqQ/i6lwyAKLmMdkc8diQjwg6
SCI68/G9TtWKy/ZuMoakOY7VpNKsXUI2PdSno+MSnl3PtDYvVm/qXxUN8IRwMTUw
x/BkPcOcZGlv1rGZK8qnpRYo5quc9VwVNKfL+bNr7H+pQ9dKr6KYTO/kskv9Zg8W
n6Ozv8h4FA+Gi+YUANi8w3zb7v5iIoEASRfF0PXF1kiQ9CqHAe/WVnge8T/DaGHN
+JUBtvSj7gnIIXrLPutHX94JQfJS6apju65GcoEqEuJ0Y+LZRn2dUbo8qZvoB1Oh
0X9d4JdIMRfHdCTqThfZb5lFkmxEtpxs0FGv9EukUzmCFm9Cg9P31DXORP8HyhPk
gTZYyrR6cWlHUqfDypGT9yk5rPvdsyZlq+cfuIisgzRxPtGdwfP0WZZBOerIYAci
RM5W/d3OJmylV15I1mIwAJBtIbqCWmcxjlMNcjoc0va6d10XxTkTHxpFVscfVXBe
zRgjruFNx/QH1nQY8hA3+oL64iqIVhtq4g9AsWvX6u/FS4UhWvWnfn1T/LDNJ8tH
2SKcNIFJA7qvdscZ9N1b+YeWpJc4JgrAig39NeeboO9g2uqlY/dAwEe11II2op27
xf6iMNABI3/xO4jxfcgT9S4CHTEdydX7Vk9UNmXr2URPj166u7WYvL2NzJ0u/ews
jkFULYN5/NHsc8q6Ij5A+Fk+fpeW5O9DYOzIABBHCh++7mtMI7yIr8WLMIs9l48A
bmT6sYHWU7rbovAktJJUbSgS95eh5DewS1EPp8Nf8Pq8TkK3MxDtJTG557uRpZJa
4azCxxRv4Tt/WTAeo0phJ6aGraRJzfPhANmg0TQERRIdgxsrsVS7zOVIsfk26BNT
/R+Z+ebcOG4tz54StdbClOhPZuD3MMDd/T2boIzQPdowYZRaE1DUl6BtvrH5QSdB
t8RKVzde7rmW/4SsEM2kuItNueQzcpb0tLMNU4EoD8QoAmhGL3lcxiRqp6itOdEw
YVdnNgHVawS9zycm62Nvm0PMKvoZ5Wbq6eqM5tJYIIQJvVNjMqeA7h2fmpsPaLf3
O93bEat1iNyaNqYeQwRnjU34JAGjVfqYUc/J4/jgi+YD7hlUQzYudqmQ4JbbQs8l
Sdf6Cw4rW7lre0SB8fzLT1/YTqkDBWtG3mXHMD8QG2hVxMXyYx74EqOR7EoBUi79
e7BigkxEKSIw08j76dAlanL3TS+z9oBGbjRm85S5wxwASf/dqujlXK3IOKcG1D9g
LlRsB6RLIpXUxwtLwBhl5WaH2fnTFQ7yvN3PdRb5MD9MrRXQ3iIkS/RqEybQX268
2sYOovp31MXxyHGrZ8tWB7ltsc5au3RTZ20bb6jZMW10hZA0sqME8geDriZ7fQuU
UEJcJ4P7kTJJ2oJ7l35yVa+/IDKOzYynkKSVPf/7fdL/fA/rze7GJUsOkuUvRQgZ
F8ct7PtEchiQxXac65GlTjbQWN+Js3xzJWHn0j+B11vSRmXBMVYiJJNsrRf5+fR2
nQhIoZ72nLFA3RuttYnXKvJGWMriUiL8Fn5BWRxdQhqywg/wwqCCKtGNGnQYOjgK
nlnVujgDgfB73xe3IAM92TumdsNl2oobo8QtHcpGdoL8OlTo+COWedM7aUNWd8zQ
eYwdB00yHZNK/nkDxHz8UZwbhHI4B0Gz6ALlVSEjZ8W7J+poqAFn6lkUa0z8kBCW
b0lg7gfzG4NICTaWCepFkfB5Y+cc5bOZ5gi0To0dUtGYhEDMWQoG8QdC5ZqMDSFN
ynHtlOHikdttXY04HJC1wPXriQsZs7CbrNKaBDlmVYewhcUKwBH2muiTcVCj+xEu
dY3yzz3X+f0Nnch95NmSaOgy9Xi76RCl8huQz/NyHzmNOun9u8onoh5nr3pmJiJy
nacnXNL8ynA0D0Kk6SE+VxvjtweSzEMYnWHQRu9AvSeaiQ2w/nO8y1x5gGd5R558
4aKeIXsq5mH8A61VBsXvG0Zz2+DZQV9p+2AgTfZQ9PQKPBuMcTcPWTte6cjD9FNG
fZ292XIt1U5aetfe2H5SCBYJgpOdXiRSZoutsCqPkmwbaWshAlklpl6PfHR385IA
SRKtMRaiii6L04PhD5B8+1XdzGN/mejjfy4kqsZFk8pbZ2RJgpkfko647mcjWdfr
rlgvjoOrjpOn1e6OPkbW+lzplhxFfToEJq6UEU1dWlX9FQ5Nm5PDn2GsHLJvaHDj
AyG+19iVE4KCd3eEdW9WwVeA27Y0JJ5eEnBDvvlLqU/3xkZZ1don2ooApX7JR9mw
3P4VM7HRi5Qra5j8mksFGbo51MHLrb7IVV8GJvl0JIe5jLu1Jeh6sutxqKgbwjnA
iv4eUiDsr/AkjjWvfi4QztsuVMLb19O8y5Wgs3W1/RQaCJcFNupY+QnQyusYoWDc
FJ/7eiK7NWbZkMTVjM90nUVTiKKHpUmKOjxG2eC/jEcha/IklbGw+b5RIL9kfRGF
xrAgX9i2tPg0pD4yHmeNkoxBrMYyT/2QJqBLeB8C2cv7vZU3/x9+Mtk96G4U81MJ
/tHbdoVTQDHiaHOE/j8QJWJGNq+F+Ahp01k8Pf8rUojb07HOpCKHuNOy/LX8T02c
KDSWubb5Rd5d9zJlVNpjAUCS7DWsiH+izukBSEu0Yv0p+G47Ze1s+NquF6oK4NbO
vPb0veTpXI2wlL95FHSNo0LCmw4uGXP8jv5pyS9OMe3lgCmD6d5kDl+dVhu0CO2f
snOggn8osq6NNwASWgCVbc531BgnTyCkm7FUlX7xc/cAEZhPr1zna5w3wbDVddw8
PkpYWm7kmRHDEUq7zcgR7RSMNQNJHTxYvko8SvgVpy703GKxQEkxRL25rYhcUUZO
31kJ63HAcZPOkhctpP0ii50K/n8onvba9PRgCeRK49JYfQ4AESkRCVEQULNl0KSj
M93427Qb6sAddcdiTkklUywPzzoOcLGXGeeHWwd/j40HhvrD7ZiaiKXnpJXFUjvC
6SEVYwcMpOXmMN+C63VwBGfHsDYIyiAq57bY0gTY4TSgKPtdXOI6fY77mtTDoxED
+5DDiiHDlwBT6yatihUIRe7Egc+MhkmmamfejLWdkpuV40TeF1QfuKyVnfYSbDri
2hHajZtqWoQ9LQL7q4eLG9Ks8GuaxoWGPg+JCJmXogXSvWjk3xn8QvBMdTxcaDit
FbNuDFXWhsfRU2+iywHXEWtLJxhlH+ciqsQ2zx7oYL4GdEpxHans7X7yNaz1JkNF
F6pp14k1MYvTThZeLPv+Qe6F1dWB93TlZiZvP13ggMMxQ41SV7b3mh74j6A+n/zh
YJrF6aksoJqre5WjMgziJgb+yT+8b7WmcfVBbdk3fm+mLmOa7tERpVhPyMOJATbw
x6ItZPpg/VUgGbXwTe95qvgxZ7RO0pX3PvmmUAg9a4WceNQ8hNyEdx42FSbbricc
yDl6CHDDzWzKPxciZDRMgGi9oCIK9vBGftOYv06KLd/N7qwmYD3wSZ8kPMyUzlBO
SL7xEXoBI1MiRujqcZIGStVujAnKkYOeCBzD7HjK5DrfNN2BfIDqBlfu/R/o3cZw
3Zj8pHU7ytehFKjccp8zZagYPhBnm/JEhJ3luepp4btoqf8MSE/2yZTcOSkHwGPZ
WIGDplk+cBG8XtYvO6et7HiCAJZjAzVZnrSpVimPdUk7L3MK6F2WJHRMcFtdIbue
QVugQD8E7VSsJUonxbuemQW0ggrZLYytPRc4B460hBkxFarQVXWNKEJCGIY4fP6X
hKUFSTunqzZqMrqrXW3VkZqxJKqw8H1Bp0UfGP7WQnLl4LHpLvQ+0AF+2t09gDr7
krdbEStSzz1ht6oXzqgVSEHdrJ0WI1TdfP/nOZWyQAzLnhYxMmGZc19PAA8GN7S9
6dbuwKsi5U/GyOyfw3lP9pPc5kVQLDTnsptI1wfBGvjXtHjrz/T2V91HwrckajwN
UTNGaNlshXf5+1jEEuWADLo9n2cMbDGW8fhtY01KJVzoCCYzcaCHtuipoJqSDyNy
8cRIm+ebkjkXfSWDmH25Azbf7m7tA9pcPcKCDdLQE4XXvu9Bwu89hyddLttQePmw
wBSVWioqZkWTqFMzmwyR+I6g+hE/ZJVZ3RyrrAO8oR66KWa+oM6J4EboYRFmcZoa
vlefBNzrDD7BQYZfw+9k/U4jPlcnoVNGQ5nnu3hVOZG/kDq/VO3FmwS+8utGa1TR
fpw950YCjRn6YOC7iLxvVVycG47gG3x58dTgPRXbFWn2AWrjimIwq3YezAz081C6
1DUYh1/LTpbHRa+iWryJcsyMxIrDKFg8zsJG9Egu3dTVQ63s/4vfwJm6wgMPlFJH
qZTtoUn5D6YjPiMS3zn091QkD56HkXSU1uLcwW0N+RkimDlhiM5YimAX4LaT9Qub
r0UjZTTQjbt0AbcmpmVFtMXhP/EiZ2dBmfPOIkDQkBesGAAjxpDs5VRDio5FBIZ6
vP86RuFk+kY9lh9cIlSy8Yx8Yb/sPJs2UW4xIRfcR1/qyAF9SuLrz27at846IN+m
WkqNX5pC32RHBYb/VEtZo2o8D5ve6krLHnIUXIzs49kyUuW6/PKbIWPFoLxOaKGe
2HKxQAk9L97lsM8JrMLuyz0Oz+y1zeRRDWm52ngozG0k0/2gDgHw3/IhxOMN9IKo
rVeixLsEz2MspoewS8Md+L7Vegr3Sb8XGNocVkYbjXgZUcB+QZK1UsJUbAYFb8Df
15TX2AgaGjEOvxURYqh2b/lxj3d9Clk7m5H5KydM7KzUJBK3CLsApGgtIQfZl9ZJ
5Fvtpy1dlLirbsRDNOCncGx3b2GBojNvZrAuthUHgbh3J/P3gMax4KOICwr1vFtd
d4W0ViuP5mfFkd1Rn2ObUCGeTNWhNXRxMU/a2Rt/O6UkiQKwz/jWRm/rVYHVgz0D
J+XzXUWm3dy4P+0VhF/s8XLjOl5fbMwGVbJC+3q/BvUTQz89KHW/g4wjX63tfVlk
q/hq5nupSyBVM/8waybX5KI0deMoKeREau2VH0q+BFH/dqq6dj4yuhmI9ZJYIiUb
CTtkEoqNXa28hziwJYf95zTnJDCIY1frmEQuNGP9nR7aPNYULgqCFXjJqiyD/Mc2
B/AQw1RQYFrJ2t2fW/MFzh17Ux+jzY2szMAF7wpjGY9Vaj3d/FEqR6mSk790yyAH
wuIq5mxLyyrC7VIQ7J4eB1svsf28EC8WlyBQE0cuehjbIs3kmSYr4ksLpjGN0U13
zWm7WgLIFPM+ESfxpawwZkunQAPE2k7RpA6c1n3h4mOusEg1bV3lTEpDnz5E1qU7
xq+NiUyknSK5muq1ZGcG4KeK7N/Kekcv8GYfn0F77WxXlTIllzFLaBnRAJJq18QD
gaw9eIOYCBDp+eKKAwBHEMN0lI95Izq38k+hGg9CLT48Rae188gw/Fb3zy/U7h/x
VunzNYW5xiLJUNa7lw+C+hGNQLRUotpAQS84XNqrZN+SBimCkPwBfdIaZhbHiSAM
YN1nfV5uuFh7LqxiGO65RaVZIWJFhi3VM2Z8jsGYPX47X4XMsVc/nCCBDfYFa9uO
FteHhggqWCHM8gFFSJS00hu2uKP0wnzqoK68RXtlVPUr30o68G3PxDjd0dFO0By/
IchBZINvqYKyhSY0QiUvXFApye1vwfKYzDgd5fg190ISYvfTnw03iErzist5bnkt
lUcbx0B6wccrKInFQ59alL/LZHPyZZUfIOnvFRGh2h764eJDBNjN8Wc8V4kEiXmq
VrIrYtwcnpLn7Nge24ilSveU5Gzzp/jO0RV+Pqu2pZblrkJsNDs8/l7O89brMD/R
w/hwqN63I70v5ug2VWRHiuicJFWgKFNC/XExBmD/Duj79fH8bKq9ho9AHt6WAQHg
+DoePS0+ws8TCkN6dlxKYjftJ5yuKQxWSrcCTmTs2lNoBrdyCFQvDBxytArohg1Z
JDlb9IVBpVy10YdZwtu6Jv5P97UaE+f8hmFZuZvKBTmumeiIHrcxaJ5wRmZEM0bp
F5vnbKkmCo4u5ZKxdzsC+UJ9WNTBP+l7/u6f9G34DOak4AztTaPm/klG1EH3vV6Y
DX8mNC2Aoh12wAkTuoO3urObKOMhDiMmE3PA+9T2yVuLhwhrDFeipyqFu9A/W0Wv
7avkpl0eqb1QoMQv0qk8yAdEbAlU8oSptGLJQVrv9ypYy9pc02LgLA4L6NoVtPWH
H7TssN3F8ILTGuLbp5K9spiNwgH/T1TRjrC6FReVOxTWrag3qEMM0/ryt8QSPciz
NV+nmwOCTBU+XH8wPl1r8m1h2/TZVuPu3rlqRYLfYrPqppWrgXNdoqh+aOSRljop
WKORIhZbfxOvnSvwhp1nt5Luq+FgBiwi6xx1oTLYffeVZff2eRh5PBNggc3SMSCo
+32xGnWLi5j82T7UJNyX6XJjctbSNqxGQFvnqIozBji8T3git7tV4G0mWvCCkkwY
6bYDTINdeEJzrZx4Ng+FTVizD0wKhpFaoPU6MJq3c80eXjZkjA/xpHNmdPZIpBur
Ld6j5a+ojV78PMDx6rR4BlKmZM+lRDw+8A3F5O0S15rmaTSmMe78j1mC0/5Xvpzf
auOhn9k39BVe2T5PBa8vvDu/XubnVn7vjyFau7wuz2U7cOFpyBrObQaFjY4MSOrX
TnK/Vj3x5XAbLWRb/7e6OomP2JKWhtED9hZJiEZ04uiZouEovYk4vdCQnMM9HS4f
zKEmcxt6VPSfbi6TB0HDJy+hF8C0ixJVgIt1Bg9lXtxjNsUU+NPKfCqxRXkuMT9z
0HUBum6oR76x0NmnhmAwlkpa85/Sqv5wtN7X0S2MVOXpzpSIVzSieLumIUTw0dPc
SrxLJxr8ymtwrHCHDaLKIsHiB3Kcul+ahXR1hNXnMdL95jV0XVc57p1Ng7ElYY+n
cglnIbMZfGdN+E/43VH/H5l99FIlYX5Uyg8kE4WcJLyl+Z0zAVQwYplFfJBdMHAu
+uA3TyhfS/PYKolr/ninNJtMbv0KSdiMLiFHn4DsQkKpqQCc6al531g9hAOXiOZY
2fioTmNhViDSM1PzHJLWgLOeglTJXee/V/j0vlTXl8BkoqbZRq1bs4G8WWdq6rB3
8pRD5tgATvo7KXSai1xByfzPKlFnnkIUxbuZ2tI83tjB6DF8Pq/3YnB6yUPQcTkv
OAZ9bBdMIPj09xSaQ2ly4U7/PP9ttGTUeZpE0Ke2Xk+Z+4JtISEqQ6QlmDuSNvBJ
z1EstanvN8Lg1ppm9zmubv9hW0BImIktiPqWAZdpgFEbi9n2jZIgzi5rN0VsAsmx
RAperNRPSH6j9ysFzXGwe5+pR+oniRPH4hCFZYOI8mZuOxKQ9BxYyBCTFucUbn98
1hVGtXyAYZ6xZArSFkdWJjiUGoa7VT/57TQo9OmbVPixHkrgVrx0IZLWntgd0eta
UT/me2XRw+HozkQRiPC+Ena8CvShf5kRFiG8jpEsxuwsFtbOb1qH9iDcDY3qZ3HB
ycZMxc97G4tl/cdwVH2f5c+oma3DqHgfhuvK9u4jFjIawFc1R1fXTcyzggzcc6sA
z5UaUCAH1lF80SPYoJB4s6st3mOPrwf7kBQ1hH3uIw3xAh6NsZEHUOA0nzklzJxA
WyFUMJvmZMl5CZBtP5jwig54SW+QqEO/7ES9veQOswSbMIuQ2cLiiKVGJEe2Ahal
No2TQEF8wDypC31OWmht+HifSxf0XczPbL6RuZgvZIu1VPdtXHDjT/r0pgJ4JRrU
WElFudjLh9gNceFqIxTDb76D9f3isSKDaJtSlSekOxKmJ8CJvTlOMNFAc8DVbqtn
VYDKP4j5fi4Hk3p/UoFvWfxY6eGMwKUzq2GArjJEhbQYTmkZEloyry+6/BgzfCzE
QuH8MqJU0DN92468lF/xetZVfTY38C0Cty+1CUQphJmxS7XWaDk8CORd1rAtrpat
lMvLMoFl2PGyTc8acJoAyPAA0TGw/V+LmKqbSdWKTu/bpMY9De8WHpjqNElNuW27
FZon6dbIOzR6cFYNu+VuKqLy+QwW9yOsNaDQI5z1lBTd8arL96AronsnjqiQv40B
vgCG2av4hHoEYXd59+R/61ByOUDMD0RMr0EcDQL638ORV7djnVDt5h4t0solTqZT
5MmG8+yBlhCBbyng8h3NsAh92haTdhhzcw6+m+/3wUjq3OEpwbHS78bQhPjLtubs
G3VDxIUC+Lw4/hNdzmBW4YmVVvudMYBufBO/aUE+ii9+sGX4+QNudMfNPcy0TeKx
`pragma protect end_protected

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
jOHqTFFC9TFke9v/yrz1SpKhUaMIYDmRBhF+kzYwtmeU6dgVPzhHgASNJk/uafsv
N9XJGNjFzbztxTyYz403jknaQaiqtLg+EXhEDe24CfYtPevTTaIdBCYYncwQSKO4
fUxa/MMWMDD6smxLCnRNSL7MiApwkPpuKVvvu0A9WS0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 44290     )
KT9UcG0fdZr90kId+RFtylfeBw3e5rEEZR1oEm7DFeiYDm12lBA8iJURPjSVoaqn
FzH898cUu2UIkIrWBSwdtCKVG92XQAXbZpylWecyyQMIyclCQ3IOl1RpPZL9wIT5
g3pJ7YUlFbYExbgO08Hr+wiiungsU4cBG6j40km/kgFAzsmDK24xlWsrAzeSia7e
IkgGYjmKlyIlKTXHPlwirYS48BRNkZsNZrJ1+QnI46bX2M01d2bBjxdDJOZpGJ3q
RCtYOmKvre/XMCp9de7JakmDehZLW70+CN21ziDR5/DXGhUfHBqgYe4ugVXhZjew
cTKmbggrGwZy16XBQV2c/na57DAa/NKJcjGBphr/YPgyff7MuO4bqR4yNa9OXhr9
HU8vgp2dtGXFj1aukr1c8DFO1V4wYnuK4f+C7J8AvBksaQZgIBg4g8IdAjGaZWGi
DTw8FJEQc6UtSAHHxhET8zuQiuiJsO2e4PFUVpz4YhuPCQQOAnq+d/aTlz/JPgIE
aisse8iJdlZV7oWxg9hECi5Wpj1fD9XK0JeCPB26ybk8uwDeALsn2p5Bx4r0WrkF
gKwxDMo9mhm0Mnduai5UxcSjGYCO9pQxXCNs52KyvB+oQrJ5wtQ3ajggGWsvyvNN
MeuIcM7w+wR3EVAg3IwL529++NvqISoJyWMrPnBC4T773jOvKbxzzQkJX+T77gBc
cMe1tfqVv+6HEtoo9kjbIXiBs1+o8QyE+AcQrLVZoyLJRyRe3VMnl1FojnQni06m
qY2aJGjkIsuCAYAJOHhysVlgFTekT23sq/o+0KyoJY4qTtsmqOlhMSuU+CV0ULmy
I07fMeApfjoJBw42kU4PMOX1gAaGYHs9xLiFOLN7vKPegsfLzs4T26hVz9iwBNjc
g4B0hm+NZ9+UelQdwX0otGGcQLrsRj8undf2qUZcXPVB3wS38zDxVPFuUWlGe50I
xvguwTbCCHGN+ewhIKBmehODZWIFZ9bgLsXGDR65TE8URLsA0w/TgJC5bif27AEU
G0RZyklfu6dh8eEXiVjPHy3RT6/0tfiL9BtS1jVWT43hKdhGu2MoW5qz0HC3U5zU
9GM0fk6GQUD+LH/SpbZdYhDXZyFV37URaRPmwoPaUzPWFcNAJGk5LHJKzr5kf0lh
957ZS4dzCoNmFiGcM7D04KP5iJFtCX1qU/U9t7sEvGqtDcWwSlDzN8WocTx+/v94
KnlprMAMi8kBbIDbX40/nHUPrqmeVgZitwZsOat7Glid+5BRdZ2BXocriynprTJJ
5rUkvtab7Am3utqY30PGAVaeoFnZljWHmeowzI15MQ63NvpFjz0vbltT8q4vB0KF
y5JLz+IE74Ke2TC+bOXaBa+1/z+bxpjceF7YOBzxGIAKFg8/9XWQk5LTPk55z0wc
Ys8ncBDjbewn37QU3tsWc/iKGds/82ZUupCXSuK7ytIM6E7gebrkSVbz0X+IWxzn
siG1wkgtu0V8AN6IrvGl5ZCQrVLrua85u4ZCbTw5/NIydqd/XlHUCepst22Boe7Z
aT1hlM1brJ7leyA/VKQr2bE3xKCbRtycfeMjuppN5goI/Ft+Dw7F0jeasj0JL5DV
f0SQmUkOdJH6BofvAHUXkB6VoqTsEJEux4eerLKekwuKTN9gk/IkFakpvKttPgtR
a84ZFQJ37+GQT1wUVQRCYZUxOb81o/B5j7vZzqHcGtT5OdoVjUhEArgTYipGZtmw
e7Ou91ccGvO+8gjgSyAHZRyZmmJs2sZ8SZx+7QK7MySERx2YEpBEaL2gqzebyqNr
Y6hD3WJQlPOf29fLKKMly9h2p2SeiX9haWwDNHKfUQIYXj4zQpVdn2u9OTwxrZ6s
RcLZlH3aq36pas1WmMZRQQMYGHyD00CHIRgV17G2WOcmnqK7wHGhpRS/TyWrBi+4
IlKZTFqLq8zfULIHrZpOG4ItrwfuO2kyYOfXSZzeKxuJlnnrU38XWyhYWzKvsN7A
I1v/3zrUq/d3y8hI4Hb4OJKiV0aZqRnnYR4J6sOW1jpjqXnWag3jGKfllFVLHzMz
Z6ZbOtpLq1ZpF/665wT939Ircd2yKz4PQxTiTq5eKHpXo3oOZXa8PonI44lTewCb
1c8YluAtzCZ2+z9TctL4G2DsRGyFgiKtfc/uqA7MRI2Z0CFa6qTzHUrwtPgLzJrO
FAfd5oDkXWf7iBl+gsvi2Q==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
QTge14LMPwc4otqmfNBNxK60mlWzzlWYw4jiL6r0vPZB4Ws+59Z0RB8DW/k6KApr
zDM4BxvMUciMnXL9KWChFgYvvucwNDQdrMHK5llfvZkL0qcEyS2PMr1w7avf0XP+
e7J9u0Y+yJ38AgFgfP5wJZ2dl1mUSrkAaQdCftkNesY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 44818     )
Ih9dRQTqOpOK7uZSR+fcVK8XAP2M7oq5ZE+WUvBk0WMS1is5gAC3/7OLReEPHxva
qHpxeEdyWq4u1iW8jF7ve44ibdFe+n+HNLHjL0ZAkzs/JYQPW1Z86K/Vbn13ilcu
kefLjBgCcZMtympv51j3gIbFgj94q/kyYcp9oSvuMR1N+tMkM7gJhHMet4jf6FpL
vEYLoOUrmQkgXFIKdoQRpG4yk05R3V6c1kje5T5wPOHyX11g5a9LyqSw/3XR8Jt3
zsqhAN/ShMr315RIEfqi0OM58BbyJYonNjQu9Kgj50q+GLebvzaFFUlrE4XfSPlZ
IflgXBH6BFWIGcvbJcBjDY04dcQTLktet/w/wSI1qbLkXzPCC76njb7AMcA/0lj6
fc6aez0a0jFuucvhyupU4PxaaCtLjRcgpOo+cZUTYgHD/TaYd9LrXkqLtUH6Ev9r
J4/X918ZbyyUal81yAG8qVGWXXaYUDkMYy2qREqf2Itx+10cxx6mIySQjaP3kNCn
q4EgN7mAJ/1fVGiRXrlXn309qikKxKC565N9VrLg8j3P/Xrv2rU4RiRpPCj0F97w
ZlGNvCgdjjTj/d58hxWpvP+Qeke+r6TbByybZhPPY7VsVVxH76X+x7kzqxwxSLQb
0QdRQcLZrHSl9nEJOr0tY2kJxDEVZA1BKvGKU9XKYEZE0MKPCuZx6IrwQ6qgeuyE
5GLujw+TUaggfKtsSTsBfg==
`pragma protect end_protected                  
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
DBKI8cdoW/Qrv2rvrKmnixihfVLsrhme1y8gmV0drrDa/UU6U0VXKnG0p+hLq/2N
vgtaqf90C9Aph/5y0EnuEtmvoXR12C9IPVAROteb5sxX6ZhQcryeQ1tN5WFJlynS
95YF0RpLR5Lkw7uBV2bqXZ38iJ6ywZXvOQdesfzxtZQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 92689     )
Zb8WEEufq/fbzqno+KTGpngAfjmydnLzYj2JSa8heEqYAnXdwKf6AhqsC1FoGpH6
u2gVaHQ7kJvfxFyL6G/xYBhs+Qur8UARZIpM6klsOWU7wqKEmKtw3p2/HBUHEAGn
qDc3dmBD3FjjfGBLKB4Eg+pfMPxgjN63pb0wmWHgdNMZ7OpT6qZvyErG84WDEHXJ
GfELSgpb8A0JhBojs5rBjR7iGIvs4raXb3o3vOG7LkKwNKTA5FG/tBD46eSNDmdb
UqsBxQ9m4A1egPn/2SJMIrRldW1dEfZBZfxKlk7Zlb2ifz2Si9XhBPriOmFYhWGs
zlRlCtoALKzhoOYSODVypvEqujGYtDwc5NpNOa/1HcwxXqgt0fxNc+jdlicncGgl
glW4sNunk3kwka08pwp7RNBc9dPXqSasdUVBnL4JdrLKV5YRiOS2pVHCx8qZeRW1
EvW0N0hUAEP2WvL3u9FinIOA/LpTboUiI4EALDyLHJTRjCJuMhWNUEL0WlMEyvv/
opvVMymycAUaOagQ2rjuxHjP66lxo5CxAA+L4GYIicKD1mKHdeTpNesYtNiZWWkR
068dSTCFWtfsNPzwjHHZs3UUkBxG5s9ZkBRIk//5ToiQvLuYN1WtJhn2eqe/MGSK
EI0yFvIS3TWrsgax/yEbzhk8EcVog/84eljwyERHuCFQeAWEEibI+odmGNwyNpOG
yEsoMsMIjiWpLWGVK2z+wq7QfrU51GLWYdGV2edwY5SJ5HUk7jsWNaOT8baX+/CL
E5wJ36i2FhCIj09QUESyMaFfFC6RilUb12/kZYXOZryvMxRMmzSpVM3Fe+BWTDIt
87DcFliDGf7ZQEekZ0EytAg0x4Sqk8bY66uDBpLqcyfGQb0wZ2ik7zY3Bhv2qbVS
xO6qAJDoL6plJ765LT3JHp8vmJstsvhnHepnAFee23tDB6uHnp/5q4zRrRa41sB3
a5ASo551gVl4DzlP0DzaATC5uBMVDXob42DwQgj2inf/Lgr8BGFWWI0LdKAHwYnr
e+tKnHS2pKEVfXeWy+Gx3HLt/QnImBfvC+qWgHmoiKX2xpas/wYq1DTbq1P1RDJv
9HqX0nSRKugrDsy73rSxSRioUkmxGQiS0YEwWbalBE8SKKvpfN2yoVybDJ51aZ3S
8L1pwTh7sKgnQKT/MOx0bBLMep7cQG//q7gbnqZAA0OSFuETBL4NQAxty3RhmmlA
GEtZLD73D91BgwT9K3fk5I9V9Xcj0O7BzpWi2iOT4yEHuRJiZbId5FhEF/mrm5Wv
UQgsBabtBrhaNYaqiSc+baW6KJFtpmFdD2YD1i3FOxDt9z2gksLzMk9fSkbq9qg0
u4drWRagSDu8nSyPOCh+LS42MFdX/2IrtrBGAroKU7qr88Za+GQhUPs1G4EJ/obj
qnZU23y/PRoziiwx1/uqtzae6iIjH9/oI4S7in3aE0MWxcr8kAT1Hsi1zFjHwFB2
CeO4FDIRsfFtkRsKsjkhZ8MjICoE2LcNF8Vwr5znxUrccaiQXzvpKuLcO9BFLFFy
0YpuyDF4hVX6cHidbn4ayT6Hn0PUBa+scoXicd8kP+zeP6Mp8vOeuPbjGquaz4v9
+MqehkhFI9CrNG4BvOKrHKiiYlVy2CFWSaxvBMAfbY60uavjXWyxUlBNkT6JjTu6
SyVPEViPDbCBGXFDmd62eJn0N3sI65bKBnj44Cwuu9+E0Cjt/61ALrzjA/RD5zgD
91W83CWOlm9uB/KXLIsk6v6V6GHONxKvQpVegljbM1Drse/2IVKtvmXg1wffLjNV
u0iGXs+wMOpA5V5Asm3ccSVMYBORSFqWlrzt+l6+eD5gKttrXMwoT+5NRlZo0tL0
KgPiOa1STkZ/Rfvo+xwCDMHtZ4nMhL2M8Ao83ZIekeo11+WHH1ojybDnAuL80ZBU
PjO/24WAuceE+lI16yIwQ58HKCUTkDD4ZxcmCPHzoyaeXsY7V6O/2cT3lh+BA0yd
/wwGUF+0KsScrRwVDzlqKsHMayIYVIG+21tfHvivv4oI446eW4Zmke8+TwkS1Q3w
dWfNCk5zW1txHbU6l0MxQFRfEXQ66AbFdDHdz9A6eoHd2Gh8EntLAdifiyL2mAnX
DshAd/ksAfzuCSuXd+XT+tdeJC770ZInZ+/QXZ5g5rHHOrDRPnIJfy5XTHs6aWF2
aQAyMstf8kddG24F0FZmQhDm3DcYI6tMdU2fdlvMGX80up2UwC2PD0I33kp6SMt/
vGkWygO6PcvHFr9e96zcjpy/Yo6NAkyqJtwrDhXqIIOBl1kLWu3WxB4535CoFI2s
DxSuKgI6uvLLuwOG+zEmlZkFeSkLhE4YV4JDpYe1Exv7uCOmtTnLjIpMZoc4S4Ih
cm2pTgz4FXv2b5ig87kAuXGhX4TJcZ5ENDuQKpQhw2fqRjzePe+55bwscW5PXyxj
+XtdCRJIuzC4aNmp8E7Lq63bqwb99Tweb4ZcOWGLOk8ti51Q0pztF6EdPCHDaOfP
RAzu/Nw47muIDT/QyIbR9jH/yzRAJR2KZko7rc012kMTzHxodrD4sHcWicXg9JGy
+VBCeOYaDwUh0lFMgWu6YLrSZjzGYalCTaVemTA86x0/1ZQ3qJevg2HwVXfmMxZM
tEjNSPkHABjnYWiaK5w0owWq2KnJQCSDdMz88Ajwnq2qj4sF6ysXPkRm8ICmdWCC
Y74/92nsEmgJ/ZYDCd0cLfYKytNJrwqeHJTad3RBTWe0X/tbbfAnHIobEAElb0zB
RFZ7PL8lVNIJ1IJksI4iNF7WlNdUewrCSLDSKVbf4ndeS3ysLb45V2s+1kwvcAVM
S0LnOS2oEJAfSP2zs4+I/J/Tkrhl9iW/wH5heT/f2O+BkjaBDhFaReQFKi6n6IXy
k7CTvJlnXZoocHSBXfUTu846vPvGH7GnyRZ2dui+tN7LZJFxHNw2lUIU7ntCTO7r
mtuPBKv4jE/bbvPPROM7OTNRZFntXor7Loix+o/7KimmbSJhbaXELoIwnPjZo7kP
MO94+U+RoavCsdMQpwNTz9nql+E7Jc4FBVjQ/5hQZY6yytR1c49YqtSvFWBA65r1
l2xX1plVOGtSmonBxgid9aCsqeOm+C6kBMimQRgbVQTA+QHkSCHfd1fJjbhieBOh
dVN7Zb4tBSkxIQX5i/TKW9DkQpJpVzAufjtTZ4Ghwt0yoDgdrfwoSPGQRYs3Kpwa
QTSbWJpvcfqcDWfrE8laKTFcP8dF/lR8OzBXI/QLCtfV8JiBvd3QEcHBBEEy1Dz8
gHn19y66rRgqrlSjTGprpo0MHGurKoPYU48KOQgdcL4DJcyXdVdWE+dakmhRLwdY
MDhEHC2B2+XTUYPCHO3nQqKO1maDmzuE3dfOmhCrJ4L+wGpuDT9uM21wwcQqmk57
Jat/9VYYgwD4tu0EKooiYcPeBTs7X5Pjf64QyTEC2Sg51AGbJBzjqBCpR7lQnLAb
IjDLWxWE+1DfpNIHml5ehQW4+Gc+J9rwHrcuqb6dblikcpDGI6Toet2a3UXTrqO1
/85OzbK5aVgMG15IyUYJ7JSDMzYpHy9YSqnxc3+k28hB4reJiwyp+S1nR42a0WBS
+ztWA3vbcFQP47cAan5GaHFZmVAteCA/+9tx9bidLUOpO/q7xB4xm0eBKmgXvKnL
TKL6bqfp1tr7kNt4M6bEGZSHz8sJeLkRDrdbwplmGs7gDuxlZXMx0FZobcXPGxpL
/mf/9IZMvLHbO0h3NcdG5s5BrH+7LqRsSK4tOWbXE8BmTzsLKynbCzBd0dfQb1yY
qFfBz2xKBtLRokv6DxNblgxUwr+SNfvjqt7HwAmg8kzCbc/RnIqCYmeVeQcUXbf7
TZl65IdLaHwsaCV63Udg54F2I1ZQEJ446JWARqOsBRC2xqbLK0pJ/qS4UyL0Ia0l
irF8TkxhFW0aZv1flXFJL80xJVp0ueVUdsVHRJXyvo57HQZw4KJ7o1WjgBZb9Q01
SRZKvWVJ45W69AR9rGi0UvSKjRXyFYaGjOjSdDo4shv1e5UnbKQYe/2JcsP2FI87
vD6pVGRaSxbsSfTkqvzOMOgqzkifVlMX8uxMoIPoS5Bfw9UnkTZsoGXRIdH1Mp6Q
RWadcdWJVsJ9RRs0V09x0w9BbpVfp6CBz2nM32lmaWhgmvm5HazpYg194ooVr3J1
O2O2YQMiid3HtVhW8Yg0mluRrEqN1bPUhxpgXr9aIpgc2BzF40gTvCHGJqcIBgHZ
f/7zwzfLuLwb79ucDACzsThyKUrjK8m2vPK5CMFkRWc8V/7FSFp0TmXNztRuFD2f
l7e2moMK5eb8xkluKpjARRHRFbjnJXhkEvZS+5gcnWAXcg9qjB3ykCBF3YTCyY4U
md98SlZyDlkI+oxQfndrLMWtiBu1/XCQE2eNhbdndKKIQEc5yFNeo/0VanX6bg2J
YtVooyOY/dxlyjCR9ifHOtjn5ClgtukZEs9AwE2LkB0jL78KuY9r1JWfnSb+zWRI
H7b6nmx7tO8s0CKExypJSeziVLYGfALbv6EDCGnqxyQkEeK/wWMZgq6RtFsxkMjG
KAIxR4Igv99iJgs7lmLyGWVlwH9raoXsV4gyjqiHWJwQ6d1xNfp7BhQPnBEs4LLC
xtG/Kp9E4ZItA1K2yeA0Xh2CVi3kNOBdOiiE8/uAglEG1TonjlxeYveL+Skhxb87
s9U+UoZCadyFOUprCwi2QkIAV5myIK2wC/RyPZpr96FnGQ+alJeTjEfD/6Jcg9JT
T3ycfoCPWbvXmT+nb35MfdHH3pzBcqaxUOig9O6Hy2wMLnyp+thtse1DwYB98E9E
yUUBEQrfrSFimrMLqEPVe3g6A81IqmOv8aldy0YgIBLU3u6C24QneDZu5I3txRF8
QuAGatGD+jZYjdZneZnmK6deHxRf26R+Ovp6IjF4OnLU50ShwSojPedig55y5Krg
KRD1ciW2MiJALMesIwW1Nh3uLh0wOmVCaEu2Mif8Z2GiolUPV/CpygFtPYnD9lau
JrZCIDN0y5EQywfIqh66pnacxw/bns2c5ZlWfyfPqQmakSGRM4YiDUvDlU6wsXvc
p1XGu1XkT82q5UaghlUuBrzs7Nu2ZuYvS6cDrTLlat26yAg5f7fcxYRn68iAoVhE
UTqdpjUlvOjH+VuX92J9XAFrrXaIG6zUppA8NZBeILq1qJkujBGiT+ZZC8xQgxip
QNpSfESNn5cFObstrY6m67VB3UBGijF32p6nR/9ucfCJt27L+GEHrSg0E3MuOnaH
BrNdK+3Un+uYXIXwObOkAuw8CwEl9hxJgGB3A7XTnZV0o+DSaI5oyAK5x5rxlGPi
yMkqueVrJJbJEet6KaZ5y6E1r3bAPTp+4J3o+Pi8p/mjxjF3hdaskGHVv3HbpqxA
WiWZ2r8D5eVWl6VYdzt+WYf7DWhiwlvRCh2dmMkupBj5g/jtZHF4nPGW8SJtRoMs
tfIKp93uJ0D9ST8MXUv+x6lVcmog9gk0UIkZ5UkTNT24kNEoDFwjlCG4f+RPcbne
fVaMsa+34dYrq2Wtm+MP6b+VpXyLJYR+9dYrk8mB+MjLH/Ds0/MGmns+6oXw7uiu
QCAkIV0b6gonmWOJL5Q+L9wiQvq320aDtAhFWmzUablN4EZpgxbTQNhghF5zTMst
P/VIVXj+XK2OIzVozLcSiRYkVK84p3J7wBDGtUMVOOQwssNeCqDhuEIN3Ahvw3QT
8jPu3OIXcuSqRKbseI4WPulSiz9n0j4AesrgTQwXF0c73Ix/lNv1SXlH90GWZoXd
lTHqPQfu2I+zAOMcojIHRsKOqhZOU3SmGaFstD99+A5a9se14ctRVk25tPcwzyHX
5ZoV0zUiQ0vSjyC6tHVKAkQJv8ZX98VSEmRmAxJEyR7AzBIG3Lq+3rpGFcs5OuVE
LbjnO2xJ7JMyjmC8rHZPms32rSQ8MfMJZkHnZbw5C6GkPYvTYzca35L/ykozNEMg
mvUjg9ypWyRMcLhMoTJ03iqoYnuuWtdYGK8fv2uLmko9g3vEZ9ibZW+/49XIIMRr
fAWkFPn/oEhIXaj3LMomEqjpQhpv0xu/uqvyil/Szq0RFamkziCNX4fgpRmXJThl
PymyRClZYiygiISEfe/Br0FYC8jmYSS5Um4pzc5MCJ7X5PKeUzuUq2sQeyThNYx/
j0W3lYhdu8O4cMA2B29OgG2yN/CAHoUP4CooPc6+xH5pFoV1m9RowVEVNrp0rgLW
TUgtUak2yblseZQkvvIZmvJ+CeIIAoYZWxDbQvZxuDXfTNcc392zINPYcJtuZ+Nt
PuJ4H10rtB+ejBQiw2B8vIjoKcK/f/cVNgs1BbWMNONRsPipqKkGWkPkt4PwhJKn
tiPKf2+FoM3mHXWQtojL9yBX1BT4dcVmu6wuHzJljFZWGKfuY1YnRjsfperew6fY
GsRLP/KvP3IyAiPNHZPsTqKiDZZhcBskqT7tvIWZHdiXerj0Xa7BmDIlmVZtP7br
Wy9xTrfDRtGJEFpM7s4CsBZvOwtXb/NdB8pIAAx5IaCNbbhBKXauFLed9ZI9Ux8Z
lQll7MQZSgNmxD8+FHGPazPTaclFnrQLKtC9ISNY2eiK5R5eV2LX/g0ByDmWlpTu
yTRdubGto9u2uiSCbtFi388p5QnQuBRCc3+CmS62CI9HHSLEMHkRb0QMQNroGfXa
QN5ZcRtWX+px1wdkY91hYTanqeEIqxOHLvliEU9Yr5u3dv9YIQSrX0nk6aau469X
jmRE5G7gszUEw9LxwPHPhtDVpg/q6lOdnsyhS5RR4r2bPKFVubbyMURz9YhxULyZ
N3iCZG3jUvYwbhudh8EHc0hnYZFiVB4k2t+Gb0J7x5kfqUlLvDL/RP/J4fEp9gKd
qccEzRGu0I+/DUYcqAdOFIq/yZS+qKqhUZUVTiVfEXpRUAnn57wt7hr4yiTISyvL
pI2GsLuWMD5e6ykU5+LwUhwLmSgLHMqjqiE7AVnfSm8SKogNdBaaIjrcgQsWwWuq
uVNkIC+ewbJGznLo5csrEaxetCtzw9hQ0bhztC7ngSe5cDro4BMlL/YPkzD6dq3o
c14Ru3TPgMVA8/pZHHJGZAHbOHYtzrmzrb+enrWt1myslXiOEtXHlXE4SZ0+IqV9
qToMQ1w6amHdS5uRdOClIRByXogwDCTW/T/VP2SucNxRr4QKAD8Uc1v4087zGrUC
AelWdI4Ls+tLpwsQnNdyNbUxLV7IYUkHt5H5Jg7DCclCo7chCwNGkCmRFgBh7nnY
8kDVWfdE/DM3uTg+R0AFoXhZbW4EtUgdQgSKGPnToyWkK1k72q4xH4p5bWKt2MOB
RaAVKV9Lbfm6Ced1ENneGWJhydZCFKfBJv5GzSB61Mr3pLBUT20cUMB1xD1BGloT
xBmliyNkmrNgqONeEBW8YvjBkFvAnAOpAohzOBtVOIckftj6Uq2SYBP9mjIN4VxW
+keJVjyZcXUggFcMe3DSgAZumm8miYdcB4BIsQCOo5eQSDZQJZpbPlAhvLahZsjY
CGBdBYdA9ci0wrz5mEI3C88Serl2BE5+gkuwHUBySNCrPp3ha/xlW/GSSpY9ZLAU
BbX0CFAjV7mPaDJOpJXxsufjULQUsqUX9Eubvn5agpChujwFkeeYdWu/9VysEP+g
mbDQfLJlfHVqmOhdN+Y12xQuJsBPIzaWTe/XpZPBnvs1UBnajRmiInqebF7O/DuU
bklIc5uIuRRF6+2b8OGYJ63F/8Ivaq9sV+lvi3MOCJaBbkZGcdVvkgluP2Y5/TJj
20L0Mr/hFoGL6wFutg43V9lYeWdJQn7aPd+6CFjATSAGHsh6e9rPCttpDM7VgTXa
bEcyY8UEcTvzIdwHaOPrUcD1dL1ueHYJvLE6+JuVYS6Pjkm22HWvtUNosnqITXH7
Y5Em6RbrGSe+34Z3OEXGaZrWNDUMgN4oTKQBy1w3XKGIuNQL4rhbq1cwG2Fr5k1a
BNunrQnC5TMHIS2x9b4oxdod2U0kzKxcOOpDg5fp073ZGAhVg/W5+/nCGXOkNo3j
DKWqdHcYVWxqx2svTo0A655DzjIpfwzeFzzY+Vv3Lac4RfNVIzW6nKRnmk9fgqFA
8/Yec/v/UiFagmvGhGCgh7RqQ1H8vlJ0YR0wchum13OF+KeSmgxlAo8dD/kixmtG
d4JGNjmZEhlO4gI2e+P0BH4TDdpOqOUxDNDmJ3XOolFt5RFO+5PWk2ySPusy1yHg
fKPRv0BxBdulT1Nzlmb9dibfsv2l2M1A9VAhmPJB7IFYbsOMBhpoRMWyZ/LjqZYR
d6naprIoBCD10I+csJFIbEx4KPJP6vJ0JC2C32v1mX8XWtl14cX77mCu/ql9wXGL
TdK+IsMbJf/IKQhlynN7fIGwIf5VmR97vqLYcupFc+MHQPK/uKRw8Y+26Wtt2cHV
4IZzZSXO+wggvE5uJ7HCNavNRHYHlR/GyfOMofoiB/TPwBtBd9Q4arr5nnRfEmjb
4StPXOzQB9mhZPwLFcN1Txxc8dFosDj8wOMEsPnZTcnSYxXEv49myVPZhQllnTXH
qqvYzySyYBtZB/jmt+csP0k2L6eOboYEO20xXUA8zS3Ru6DYMZAUPGoKUJ3LJrzU
tghWOA9ZNKb0f+Sum46TokfwFy6TvLZ81eq+pvFc7c3hoyxBZck5+xsWCPh3gQ8a
ARkJ25i3P8u1T4M6ozFb72HGTjomgl+tYcb8GjLiO/JjGE5Maas6mhajO7Nh5Tme
sXFIDLf59+b9TOPWKtjXMwZS5HIcdyRUQWFz8qP+Bik1aC/a6ajBHH7MPWmK++4F
SwNppN1iazNivcoVMtxAv5wWT6mTQwd/e1hr0ffG2iHp5HfaCNdnhRoMbdCl+82z
SYlSyz/0shy9KeTZrnWVugKjztc+d6NQV+RJJqKS+Y4vnxSd7Hi0k+547rQIKnZr
4Akb+5PlQOfsZFm9OJ7YEU22yAWmCIdVroi8myGuc7R0UJHbLWtlg16KajMV18EB
M+9qgvy1zaeWL/t+tyYaoM3zAdrkl5P4JG9Q/6FeeI00dwJzp6FO0QXyKc+ePifm
p0xXRd46xYg5xadF8rnxUWaXxuxux/JeFBylUr+6meOB3G7KKKya14QlIYPVOtt1
tvReXF38kbtJoj9wW0Sfv4QvkhxW8XOIEzlXzyb8Yr/5F/RGW6MebYjMrSlwKO02
LOF/eDH82GDpUSO8rmU8Tnpg2kwAfF1BozbMx7IbK7wBIyfzYGQi4mty3zLfVy1D
zFo3VgyCoF29nj/P3y8ef+PAXSLdJj25YqbUWSR6Csm/ATyOG+mUmIKB4ee+oDir
vaVCAmCylUjBqcAoUhfhANhEft+v/W8pBqdSCDPr9rfh2fpfyb13sXgcXkFWJ3y0
EJ/57MMkKDAbdtT0AI+I80CDe8iarErcEMDQnH1q7p4pEOwp6FVwTiEOAPolu+r9
Ku4rLzWOareTv+3ZtskWlHnFPDUjvrSTcKiOzOinvrJkUzWGkeVKDj2zDe/dyHMq
FBOEdTeAbeVGhWaHVUNNhe+JUSjpk3ZOG6hy6AIiF9Jl+hCbYo2r/+Twgk3tsczj
lSoS4sOEjvv3MYrvkZG+oKJO9T67iy1+HiGQbZOJkR+7Ye6l1xzZ6Dy2VTU6G6n7
VmhQyFSAqrEexWl50Whhsex+npvH3hDjM179f7BM/xOhxMsGjIQKZvJ5xQqxxPns
Kx0gaTVWqO3gDHetiQTc9kio91ske42ldWTXVwr+IECe7Ii62HcEiFgSGeUp/0BF
vrmwmEptknnWJIP10CpWhqQ7/lvc0kISFryuryqMmVBHmRzjdSUK5jcb93VDBJFJ
hJ/dQIVYIyjB1z3LuD692LCs2cJYnuDpnLij1FV1cpcn5Rkbq+9j4WLRAX6P0CCH
Q+FWunIW+YV/xT1528baIUvGceXOhW93bXScNn4E6986ZgofHmof5xzR7S34n8cr
g1RZKnkdSoCqAVK9bYKk/lPH+3/96NSPgSO1KrzIriEJQvKWY4y+cN+8zTScfUOt
7tbOsADJM3/bn0/oYRje0f4NP6kVblbbLs98u6c94YZoCVEtOhuNeLDTYTaSRout
Y8mW/nYdTXWbq6V0TAQQZtxs4C8k7rvbuwU5CV3kLROPq2USovz7NYee5DuF0IAe
VUfb1rHt77Yfl8zx4MSRd+Bp09giMqsKFnlA10rnFq/JeFnGxJ4y4KoC2o5Bct1Q
vMYLy5x9eAt+JNBx22DOXIqG/gE95XDo8e+ambguWBiB4IhKoIaslDzGok75cURV
xaE5u0UrtbDq/akc+s6lo9TBuBLag82lQZVLH+fYgO2frawg7Uko075tgspBFZ6Q
FH8ThjYXbtL6BrBBr6OZKN+8p8qTs5xGU2PjKSOuxtrEdOPxEZvxcFtzNxoPk+jq
/nc+rJtk5JEeKKLIA/F/G3j5iZsUnP3msvYw1wM6EqgSkrsQtU2uCGzbB10vRSFd
JAWkq7Y55+nEksz9HYzFuHI+y8EMbm6NU/Fx8LJ0hmp1YuVtdo1BBp9t9mFhCzu6
HLlP+5gWb/HNc4ZX4zxnpo1vdYU4QP4muEMUDWotTSxi+RGSm/purGfA/x/KvPJW
/S/oXz3DlpYKr1OGpFun8s9NBoczAaqUMsTzDwhx5bskxK02BYjWqrtdenSoSQCV
N0kpMtnj6MTdfhjt7lkwSNy61ooW09DmydS4G3oFQEP9UtctxuUjUyT9E6zK0gFC
SHcsdgIfIFJ9U9XLDj1eJHzQKVIkNmXERnkCMKpQN3ZTlzdluxmROHAcbac7fIUy
AyeTv1O71EcCsq4JHMpMXDza85wUqsbmomnBAyHWbQVMwT9y+yxdsiK2IJ+5XuoR
0rvQLiKW47wlPP5YBgHRjjYPjtNt77I0c3CN/VXvIDNI1vH2RWndUWTqGBi/DTDD
B6bN8QavZg2vaJTIUS5fj9SQZ0gAlWuyokE2XYt2R4GDVjgYB0h0shLr4jrT67nl
sk63cjGuaC/2OiQRgfDbajcwfdBh97v7/+j6sSCirT2cGvey4FESaLx+dPyBZSc3
DKfVTa+2vy+mUFfZRhFKkh+g4yAAUYFY/34GwZBMynvwlboLYg2WzZrNG9/7fWvs
OuD1bAn8L35gky2i6p6Vdh0nNHn0/6OikdBjYuejLTpsw1xYqEesFH91r7f8vm6u
hJJMy0eUO+k5vfKRJG7l2imeStLs53CuFz2bgFyuGBejz0jTTeW1reZTAoQxf4F4
hiJ4p479f0T/39CfIMkxjuGpPeAodsKcmmiMRwTWbzsmYMs70YQ/2NtgzENXG0JJ
033GuT778zJ9eoWxHwzCvf1n1sz9iyqI37KXzuTbeJEFU925EGCThVYRMeNBGNNK
BxFF6Fzk7EHTu83fTDbndlcr0R0XMLWGDN0VCpmT3GkEfHErGth+l3tC68gAJvSa
/hP9Uj7BEmMQSBGWtbNJcZ/2TkNFv0rPGpYFpxcEBSnUzIYRl/s+7DdoRwa/qQyN
zt+Xg6k7i+Myv540v1AmpomRncb8CazivGtqpA7UUqcJ2Poa8jtpIOWMiNB+KT0Y
9JEqQu6Tjq8POJ4cjVaSxipJyRXJ+0dRUwB3VaXVbOqqPWQoH3/t4beMd8BAB6SQ
zfaEF9IfmPSLwPvbJyyjRF3Ogx7lzHkR5UDYzLjBM7zCH1CjkVXEq3NWp2dWJ9fx
NvxjJw5L9UDL7F3n0W3LO0dHqy3q9yQXd4OP7UJtOmDhBmxbrs49BBjVXMEm7/4H
Ml+uLY4ehKCloAbptjfjpmjcsZqbuiV5yT7jrrH7MpOSBEj5aMPlGFmdxMFCCQJ4
eHeqtVv/vNcDGKq7TveN9tWWLyNSzg3ho29QF+wr2V4AvBvVV5lNSNBw2e8xd3di
JVOI0FIINH1V/2hZfEGnl+N3KFULMjg+H4Rh+XRtnFkdrselspPOmq+ZmB9/uMRh
mQaoFlYHocaZwxlm81vuHfh+W2kmnBorZB9C5u4bcIygieVgirKiNuo8BlyI3Xc6
/7OifsQzA9vkRYOVU8SxwyOwHGa9yMkf1TrNsV5GFW6DVpiuNZ7v5nAS2SFPx+w9
nu/r0gSIhsZQBTdWmWmyu7FzevKnrf7SSIyxVEb0X60zFZkqU1KnL5Z1jxL68mPx
zUUKUJ8g5RVw2dSlyQpX3L3lw9IPqRDxmzzknrjb50z7JbpLlnn5oQ/jA/+BYmtc
LClI2Rl7aaiNzQE3qp2U/PNHqwhmRH489rr7cXgdg5xczH9u3KWkURvQgAFtjCRT
KQs+ZbaTe+VfSfxuibI8SuJuOucD3JHgB/qxljE8b/PBRYtaVfDNpVsJK5F7W+5c
ZW1Gj7phlqaSly5A2JzBk6tqisDkjjokWCZMEokdkWNw6BdwLMg61NYkh9sKibJI
AVzUNpr4YGcrEhdWD/cgUBvsuWuIlTyh+siEJ9UeASk1C/efbw6VtOV7ygNMMwa/
d+DaFvYe3F1Wksi0RrAqq5eRaD0ssKOeZhL5EBLe+0qKYw9gSCgN/fE/lUa+o3Sg
LHSRnaL/AgFoZzWJYqjB0nNfofLK4SEWqiphlHeCRfi/qp/s55fg0LoGWKDs7gkI
k0ByqlEWX3dnx0V1ojkRp3TayITscs4QxK5YjBkMv36C3xctWTx2DSXBlKGbNaTQ
9cJJ0azwLrntNH60R30hw+Vw3vuoV9HE+J75OSNX1ZW24BeL5f/4EgqmEnN6saVu
4bOXUtnboM+nCDhlvqp79dBVrgwS8wsC6JtFX19yQ2QTj0xafCsX83e+2NBOPa8e
inlo7Vs62DNU6cuNNaWXDT6FdzLQCPAKjvvD4D4Gve5Ner8VQ3fYi1QJyoQOPF6Z
K7fOJB+brZLK3Pa3dmERJiJ8p3i4BhgJ/JsJOIDDrzZTUspM0NSFY2Z7KoXK1KqX
P9K6B2X3yPuzssY+wIKbZL9pglFWnEqfAAaCNtYiN4ZgWAsAQV8qrirvQ9oyCewR
MdbLL9NFHB/sX9yYmikhH5nS/gVFwN6nyy//a4lK3HFQtNzeuY2r/bjKYfGyGPGY
CU9gMMev7/RyFM3TWT9USuV6RxZGQx1618GXfEFHe4cHUSrAcRj4mfaL1oGDRopS
Snh5qHd5W3KXn+uuVbVOlU6maiUNe5rHwbh6fjQ44Nsd1Wp93alfNXcUuSWIW7Mm
9+a3AO4ktz13CkWndWeSYFSg1xcP8XpOAS5SV9HUv+o6/sLaHwnQm1xGz+QvMlM4
d/FsgormDbt/42nu234bEXAYTY+zjNikYXLVAKi+FP7P5oizFy7hW5BmWPXK2fHR
55r0BMEIhvfAqmDl9nAVSRSzQKdV7MNgNKtT3xBRegh+ZYwmMXJ/rCRCSVkO36dH
KbQXtw5HQuBHt0LILdRF3o4SGUPmaia2etIBhfeAn3V2SStdLue7bSmHtQrJfFqe
aSYzz9QO0nDS+HoSyLSitomsbVUrUwnLLxDHhxNrRI5h6iie+MxXj8d8gDmS41He
tn4TiRPxMsx/FECawc9PADU8N+A6phvfZmZ6zu5k0C/4/Zcal0SHXVA/gXBYJoYa
uH837szqRe0CzsRxmD24f82PDPsoHLP3zBHJFOVzlD4VOqe8cdN7xIeOD/RLqPpM
Q3yXKptK2cXFCV0Qr8BeQJ/6UJwyUzkFQEKgiEufcj1XaZ5hVc6kLZOhLyTk5tqT
Z41r999/oYY7tS/rXV9VYmBHFyQJTpnv3pMISCMNROn2iUk01j9Z0BobAi68Q6km
SXheG7eOWuzPjXqopD0GpeR0qmpClWh753Q80bu0ITLeT4HCRsEImRPdmAII5b9R
+uzFD9rBTKvw6VoxH2fDE7VamWtqRbUkAOYbyKX1ScGF1QnhqS7i5+I64ZKu3Gds
dB36FgKRPzlMaGYNW6TACtH9ybscT35x+qbeRwwL4wr1hhXcT2UFZwIRxrFatc7K
Ss9SGRYxEi/78usjuvfGXd5LnXnl+9H/r7wDcss3v4Aw+1LSL+gdGT1yFhwsx9ro
aPyeAl7yyLbjcj18pbQa06Fy1ajoEdYctEXU3HfvumYLPqei4vHHnSNrL7GYfzDd
T2DnNs8GCtjZhMQCZRlXyGOOYEjqo9iGjTu3vWT4iyC/gKkFNldjBkZj92LFSIaz
oxzsOeFGyG5UiPUoinFRo6APxZNwOxLwrDJjX/2SGy2PNSTAVXIe7ttaOQifVozM
OyKI/svdJhNY3oOnyJgdoqfTqmJzv/Ap2hDAcCVn6aFjO8iStyo7uARaZRpwLF6j
bnUNsjv1V5ocdXLQbQLzxeXMSYfpxCWla8RD7ZSMFdVizfirTzPoD8DQMB3AMOYX
sd1sWxA6wlNWow1DKBnzfNw+9rJQnVettvJWwgwdEfmb56Sdf54eWEhpMj/lrAwS
XkZ0Wz3cfflbWNSRvA1YTDBx3RKFcPXHl/qCihr0QbzlNP+LoKNv8oTbPNvXZbPo
LLnF65ZkIOErkkZBvzDFKb+zP0SmZ/lLf7U5ZFQk0Eij64nxGlgvxqN6r57Rqh/Y
l7OZueWiUSVdK7NFeNrz3HPo8Tpb+9T82JRqbbVJ+YfuhqG1NlhO7vxK9vKU6jda
jbaKYCM79CVn+XgaP8o5LAon8CwkwHXpu6hKDVPmW+0ahDqWTgYKmo9bn3ZPFe6V
QLve/Mxf4Yyv3fFAU6pcfpaZMmzbchQdz5n0g/mT7jR+lVKAjqzfU3nL5S4P0kod
epxreuz8yKmJYrGOAIyBA1vByK6pyQVV0TX2TaFnubFvAEvj4DHC73I7Iv8heXf0
4VNhY5ZKiYQwtJvc3tHg/oiHDmlL4WKIMG9wgAOb/+EFTv2f/UvG1aMmT4xPHYcx
so0aJaz7EyVr+qerDuGqBP3LxWwwSIgBrH0fviGR2VZPtK7mHT70z7KM59Ov0m7D
D0xRS4/QS7eJc5Aw+0diw4x4f1oFbzM6SDfavqQ9wXltJP6gdgeCbYh97P0Zd9Ro
xZS6RohIa93F6Yfldg4aUYIHZqLo8uPBvlIgT4x8aNjG7PGkvNTcUiFoLauBqtek
/s9PfAQp7JZY2hFH31NHZ9YC3pFQQ3li7KRGW+N3may37iR6BrETT5O+5vQga68b
nFBTAverN0ulvZGKwyxZFz80QIX4/uUQioopkvRnTVGfqFAfJZiar9RjzPiJNQgj
t4nZ5Wc4qMfG/inuw/lfNtWK1/i1Z1YKp4mAVNG/MPe0JXm6du1EMZpTsZEHOOzT
mDtCCAF4WQw/uVV2EEhX1I/7kTxOlwGsCj057p3PwuKH1/mxFhtw5TyutTEIAG2x
6Z5jHIj/7BOBVcWmULgPhVIFr9wfCqd53DLjMO7Hmfuvy/87LeEYAloOQcWY0ih8
WBHyhLSLQA+HzYmdvXXT87Noi3VqXVHpT6L0c7P2zkb/mDZGnBF8kJyyqFEteUFm
QvUhRXhnQ2rDw+LygUPPlJGt81i1jowRhBPWudY+kjOtlmNFCSTjFP2a78/hD78E
DfdiPzwPL/hZ2XHjQ9XlaLC+TX4AK7fIFal+7Z09y6ylxNE1omotfD6Qt3GOEfk1
65OloRyca/NSzP6cUeJIKneB+BOg4SyZH++/LLO7fxy1iMeXI948AByTY4COcYEj
GhxxATf7WCyQ333EnhP5fA2Cxvxz5D9KJ6xH2NBKrax923G2F8m7ajjtiOlJAUJu
GJ1RJV2cplXiUchR1cBcJu901jMRouXEIMj30iOJjQqbFi+D8YTosvGJ+UiLmIGE
ggon/BZe+Q9uBRv8Que4NQ+JLtXL8nNtHfPc7OHjIrV3LGKtokqIBIkoEKNIUquo
aRAgF7r5JRSBatE64cQ0CGud/yGUbYXE61vSdoIY6gJGnYtwzb6nMAS40CxoPRgK
YghvoOIsC9/4HrgC+yTCVphjTAWKFymFJZBy6wWoLYn7oANV5iC8G9HoUFPbA5cC
im88bBp4jkha1kyqJ781uGPjLOp/BZ3um44pDnQxianaAZl+MWO/QUmNzaVtVq7B
csnDP11vvRZQ1G2XZ6gVk6F9ShpiDeNAYAL4peaTx1FLo/Q26gilxQyYUcKrUQ5s
I8hNnvlFjj8+CIPp8S483/XnhES3RifM6HiTnE0IBawU9mZ7wGbzIz+ojjrv6884
GRo+z+0T1bfCnLMMc5LvlV6WheUjX74RpTFwwTy1aZbnyQAtuUB8zlF46kMhYtNH
6T5EwWXYYMpR28ZFXK84iuRm6/wavxWVxw5NRF4tpcYP4EIfxZHaYrkWVaL+ZwWA
nh0aNbMTidNneWrTzeJoRasoG36rkyev+Uk2iZwZ/56iR/A4acPnUc/QR8e4kO+G
q48HZ3PmU3ML2GVMa7UlSnf3ry9HjD3giEnqPR33rPq/P8xdFP2KXhVWVXHp/sAR
VgnDdv0O1m+eiq0RhNWh/NRkaLccxWnGzEOanJmFTThe0dLxkPk9pcunpi/Xo+/M
we04CNI/mwVZ4yIv11JHanx41oaPmgxQUMHPPSSFWf5BWJ+ZBWQhuTbgJ0jIo5m3
3dZgVLZ0246TgshC3pFsuVTHyopFFzjZ0byKSm7uYizEVkbR1H8IDYj5apd3oKAt
pm9RECN5BnKnGmK4B3dXFNVc+sDs5SN+AXj9+3IPx/O7NQ7yM2NTRWManiSUogtQ
L249oMNKc+crUctKVN/ey16yWiOEXgu1EPe28lF0tXAIUDVus1v6llDffyFIaggw
AzzKk4Bkpkexebv9jawYMXWKsvf3xSQxW2hJeOUGHy2QvryFJW0URHgQxBpy6tz1
lN0JzULzE5aVx8L2H9tfF/+myOz+qeauTP35UVPv7ICCQOxHrUb+/OGM9FKeyGZ4
Yb1dIX62Yumuz3biBhbftlSeFE+9moBsX/gyP7UyULMKvriGhNGaYW5B4I9P2hpo
mLH15yJ+qJSrYJUyQl1F9RwazTdDrZkq510uHo9PLRyAftNagnNp23kAi0gH76Tr
l0iMgQ2AnSiTRLj/GdwvfqoJWWFuaHfAzIa30/dsVIUSVzLPW9UlqHlJj5GstRTy
ZYFirvYmidEWRU6Fa8UxsoMts5UbyiroudKHLYOwhz7gRwrB6gR53QztiVdHNRDC
Z0PYiNIV0iQEmMl0y6hPmqWlkujg8suytFwx/BqhMfbxlA7TDXEmurDTgaFenh6w
/gGEKgdg+q3d6OJEzmqrkNSjtHudD4RRMqxuCmRN2AXxJImcRE7dJpKeUOCwqZDM
4CaH636CzzfVw/2kxS0Dq8FeyTe+qQdCfAjVpoSXIxv8YHRYInK+zvRhZ4eEHCS+
Gp4JO++NiNF5jNF9F3l4urdS0SJrwT+CrH8jTgeCAsFTk6hn8+fUerLQZA4vpPWj
9qnyC3lbe2IQjfz1F/XG08Lcs+yW7jHhlHZjzCugb81nyeCM/QctjOksWBTpwFHY
ElabDmPi63uH1GAb9hD2DW6RihqZXCWeHy/RevWcRV5kwjrrtQQ/0rFmPEqhO4ni
EhNtZokLMCnsZGyhgTBB3kTIFoXjUUfXG3gzY+VUzHmH3gyIbfj/Ye8D6nhOyUPi
zbcTjrHrISJDdII0GiOIOlAvWUyc/aNGpPhE7hTh+/06GSxBtVYYRLtisLwqLMuF
noiICk/B31HkIrP6DubKn7g0JesVAbZ2WMMGrTQG2pSN9m8vw88/cvv1ZC3yaduW
K8d6QzBmy4gMpa97qGNpPRCMzkcvhgJmYr+XHfkTK6T0dR0qtOLUXjukbDu69CNI
ZcN6cwXtKAe1HxiBf77D+WwDKgzBvSzkmsLE0kTiqXf+BwGjU5/74jrOtBIV56ct
qqzI5lL274oQvjW45zJLqQeKKdy7aR+fb3t9el4qJVeHoK6E+oMUjJWDf5KpGIpC
gYF1yFxAnyh9IPFfKCzjuGhw5dLXhjimslxetmrdyhnIot0y8cTrOsqwhujJBFNb
jUM7tkeKm/+bHLEJkK+omIjrmKwx8VR6Hnb0ugS+g6uFFk1oNbWDMPY37Q8eCGqY
tQ4nKCN2pjzrS4ENGIc1pF4Si4iNGWd6ihzVBpRU04+uSI5MaK1zAWAPFNyd1Oa3
OlIquiFdp8tMqLcVqHx/8exSZnwUNFocmqfyZhY60MBTuAFforOZUtDaSsBVh+EQ
C6tHlcbtjoaHIdZhOL/QVc0jYw3+pvOf5M9fnj3184UBj9VGlhfC/gtsvBE8EwyB
kd37qPM1hfITnYZcWHe79zLQZCHVUabIkOv864UZBVBkM6Y1WGe51Y5RSIQ86xLk
E0LZAednX6d2+Iz0GQj/QtTHPm9HylIEKI2tUgAciExCbEDqZ2pELDBgvow/qays
3b9kvQOdnmmom9wPQ3ryvUCYIRWR4vJGbpvUZXPBFM5xVbkYaFQjf56C0c0qZVQd
P7DvnWRPhqjK9KekaRoFL4LbW+78n10WQKBZyLgjUAq+ZAUNE6kzEqPSzapHEXGX
X78DG/Znx6w4LaDV9enPgapNpt0j5b/u+bXkPmuyo8P9irwInB36kgUNPk9MkbLy
MGIG1e2PuM1vaiYKCiFPvWwLXd2EhYPLasSKY1s6EuHTa4XYjniYq3+u19RkCqod
pA5wSluuhZX2KFPIfi6+1SQOTnlwU2YQkmYqHINA/K1t23JIiMJDM1/SBDNDbwtf
dfjeaVLe7ggFKdKNILaAAk9kZCUykeV4MTONp6iVkVAjP3Iuh7mXjjl/A+7FjhwG
OqOnFkdQDH3UzDQiPXri/gBa603Wtd/Ngw79c6TFPE4G4qgMC0JpaHUw/QJFIjNF
DPB5Js86t8ZQgmjtuDIrGSqJ91sLLk1xG1lBKl7Pq7zZ/ikq4L6Kd0AUVmZSCP4B
KPqn1ppHQzQfPB9IIY8fcqfjA9Umc9l/YodgA1inxRLAFyd/x79SC2bDkT11FQLf
N5nJ3fay6gRarJHpALy6IeJ0CGKCrJ9EA8a3lJmDO6hqSEGfmzDf899WYdd9hRXU
d1HU3g5sHgg9K6O4BIv+OQg8fa52c3FOhIalGeamVEMnQ220sux0gbeJ1kTsm8Wx
PanHqXulavRNr72+JJRVtYqyVh0ciwteR5dfcaaEAPLAwaJDSUL6bAolC9tokY0p
siPjQxmi0ZinNx5JeDGsWgP2KR4gI7wyJJ+y+M53kBzcs9v6RW27ssu1EXjaDwhs
6j+RUsase4OgGAWUXO2wCdx4h6DgimDRdq+tgn9ZqPexcGLz4vzd3iArx9bagHY4
Mum2/HkXSqJBMAh5QgSZJZZ0InGWbr9lVYKU0wUKMtVNMk4Dmvh8QNiwSKgaD5m4
iXsDgZ5EhjSZZ61Ju2cLpXQGDUWaJ3bTuwu/VNQg1TRWWppRAib/hJSwe06CdZcf
AP8Vv+ZvDvj/g7ry+OrpJHwL9FKv3PO4RPU3FvlHi9bPQvVfG5o/6H6/tnWaS0Gs
q/MgPMH+237ZBUPijO4K9da1OuQ0alSTyUi4d70lFGK6OfwZzv2kBHuxNUTkZGNn
14siuNbjjpkH/Km5g8jpa2miQm3RziQC8pAwE48pj8mrnI9NNhoWjKGKoAvdjLo9
G+z0n3Es7WO+8DKBpPuDOKgwuJDZGRklosAiBoL3zLuAyupnX2z+f3/tP3j9gq8l
2uA7GlHd0NvZtk/pqpuaqg+MN0jSeIoxpcwLTjD4UgEfouj5Qugs+SFPuNw1jb3r
CGDQjB6e3IoZ2tzU23N0BbyxdHZ41eqUYq5URvqcSDkmqoU1hhif8/09yxSeyQ7B
alhd1Q0Nti94clTcsj+S4kgU8H3dPtX3POPUl5GULhlAU7b3sTi5kUpWPhg4ZhQ/
QDd8qfiERgd5tcFxkPXV72JS0nNU8EUz8OZ9UqCccJ3fbHnAVVVAcokPXzfa7IJ1
C1td+IWzw8rk8d5JOnJwjpbdjPWaau6/AGJeila13OdPv5svQQHgvQGuteQgxSO1
3sJGb92s3ThzKHROFavH73OfGzZ5IhXhUSe4uGSHqFk5f/PLBikOIqLpYi+QlgLJ
cER0DHL2lNcmH+D0j7nL9/fd5c5qPah9oNUoBPpUV3tYtzfO3UqtcjMqHnJEW9Kg
3s2AFSnwdNsm99YKGQSHOzB9UfTBaYM8gjD3BalsaW0PJFRFd5/y0WKb4iZM4vEw
iKB6W/msvK26SZHV5IFxsJfRF+BM4O287iIKXK2sbf8mJO6JGAPpG+MGS3gPx+Ph
uBsMlFp0JdKMBCGYi7bUZdAHptdcQBObSUG0XFlzRnkeofx8xbKydQcIhp/u5bof
UEHSaZw2lxjMFdg3HUNWfyAzaiYwqL205LYkZ4BjJBfufbefcMeL0bwx+EUI89Ak
3vKJoftF+LZi7aFuJsviCDrrVJxVMMGIEkDco6AHpvwpsmUydhkwNwwGqofDp4N7
ab4ekk8LBXTiid93i1jCvYVZaxjl/CQwC4+A9Y3TUXKMhYHzA6hBlqh3MOTRckv4
42A2OK9RstzWaJJCVeNL0wncQpTSJWaqEyq/tkgeocYE78zYpIKcedckgbEPUAOw
1aiWdr0a9xJxAYwxdkdZMbgY9XE4Udud4IYeICSvtiWP9/cpqEa9FAZ/RaTXGb2J
4SVhlW5n/7K1UJm0Z80ZX3T35MjZWS1xtOirTc0SOy1A/aeqe4r1xJo6ZVN6/g9k
Y8ozjpua1IERIClzMjbgsdaM0BNMn4z5F9Pzn1hBTDEILi1MXewusQpnYlnj+5zN
fAqj7vY646AFb3UV5/i1Xu2/NCWQY1HU2cXmPqZr6G87ed3lkYgTLvriZuziKXu9
gFkl9yW9SBOsU1z4q+R84S6ntkIAPodmHLGfLtwYLB13QlgplNQ3tnJ42k714EtN
8KMG32K8EpNlEtK5Hwb+w6q34JFBmby3rN0DIKdU+i+xX+xF6/CUePm/q7coTuwj
Xzq9/J6A5KFR7Bqubi7jtQEocbDcZaf2DaRRNIIa7SVja3JhtsYJq/Y9i7+pyznk
OP7B8fl7B/TkK7ctoqcano7fpjmfDxCNN8FVJECiakjfJQKQa4tfg8v9yaLmZig5
5tKsMf4+S+k7cK+xHWQGYiQR9V7uvkSzORgn1vudUkaMw+N0kumg0ju5+fMIwTOH
jB1/0xGXkzr7iUsvBc2ioxojpwo9fYgpoYH5OpA+gKvUR5jhfYA8uPkymhOFTdy1
EKN6agOQETZWkT10NygeVqHMnTqYrL+IBVWZdtCzm2UG6kF87oPweN8CR9nY9JzP
yYcAydg75kKvxUxOdb7uYT7G78183XzJvXxvCGdd0oPl8xdp3MpAopmuD1KAMXRF
91kDhlbqSYneZpqDH3QM7OIoy5V135wRrmBvd2GEH8rEiZSnVZx3ToFkVGtj0RSX
o6XZgqaBvko3smPbb0d49bteK0IadPHDBoy+9bfbDkRrJ36WuTwQ/x2MlLIy1riE
Dz65GraihHAE+xdECXXfucBCKjLXh5Ugvc4y5VkoZ/idQslAjx98ex8Wy9w4BvCb
3mOQkS9wpEf/fmO7Xqdxj5SE/FTrJrqrc1AQvMUV916oWG/papbPclBJ0xUl9dGQ
M+ffGkZ3CmGCtG9Filfrys1T0HGIYJoa7tBbOflDKLy+iCrIk7FxY9KYQxdVTETr
T2eJDuxEPWhL5cgZ5faDIlx28MJQNMfrm/bbEgX4jQLmq5F3UyCZyvSj6lHIa0og
6Oxj85BAycnDxlmueYSFhaBBPYIAegmqpdio9as/YRiW8rpZacMLG6Do+fVbuU/X
/WVyZ/dRKasSKuZZSUUmSBUHwPxB2dN7uZyOJs9SMZNfaHeRRVfQy8ptz6VE4/ZI
4jzz/yOj6kueeWtVFvKbWkoK+vR1ecZZmSKWXTkEviD7hXizSU1h8TWfisz98+zz
MJJIOXpY1Z/aQPy1KIm5jrYnt2rJDPPzttaPhcVX6F3W2uYMwadBEEh+m6sW2KjX
yNB0Uxg5bpwr0W0RY5bEWbSKAUFSe7GTSrIiD9fScAmF/v8CPGPR/D4IMTL7HbKQ
K2Ud4W62Qb1fC4ICAvXaqJxjX3o3cIaaNUKKNwozmF1+zpvXkhGqoZF/AOe7kZad
PC/UypltQMb7J1dzGCEoDdGpywpAAxUysVZctesDjjq1/3gbB3My+gQcoUh3F2lL
ALkA0Yrsz4N4HQiy5KmIUvIqRhbD46w1uwA1x3A5okyP8aU0ku979LlsYhi599AX
uxyoSHxlZ41QQRXbIxeBP5Y4B0/tLZKg0BjhZ4/EECVOs5xn9dLkS72U4GvdxCjn
n6O5kakRyL3cvu46VfQsMl098IJ0pU7bIWvBWQlTZwQUD/RyD5DNTEsKs7PI3LQg
vTsC3CUO+M87ZcQIk78X9fIcs+s4UDqkveNBNo+v4V4azeTQg5Lrx4dbyLiFe9oI
G2HlbDPKaRp15DrXQ7yVVoZUETeze7BnQDjZKntma6B59k1wGqyBA6kbTT+jqvSG
RDekaiK5xteFDEnH+rwFDTS5TccBGTv7+FNmnBdR/RxxaOvQ4pmZCzvw2wznK++9
dCYkc0Z6DZks2cfLd0ZqcCA9+7lat80vKmTKjS7XDLD1jwG0uRnHBj6sLIfhACgf
i/C8iYi7OLir853cpjyw/Qb6ZIbnEt7bOTI8lBAQJkIUyw2webJ4DAtO7E2FhIs3
f9/b0XdRyGwvclk4L3E867h3oeKflSy3bJDCneVzjWY2FnJ+vxdTAImAvxG5PApT
uhbFH1/+wgI1MdPz7Vy4qU3S2gURuZfQnamew+4ebG6AzSclnF0fBzThWeSIBASX
Z5S2S6ix7CzRPTVu405Z3HpIVxV8ISywsU8LPwm905VQytsU9bisQiePEhLJ4Liy
RmzTsD6WQqkjetJhgcQgxvAvsc0kkcJrAXT5tCwalwvHyTudfeibAIpnZjmh/XEo
i9NMPWcAjDo3YPn0b8Gl+E1mc+TJXWHEznbHtrevqCoFRBmmWHxSPYhUjN9+1/WI
nLbSFaBuE0wq/BaY+6p/gnyOpMndS8pn9eNPZq4oyWaDH6r1vwDKvJ5aLVCAbl2z
uVm0qMr/SBf4UxfofIk2EW2CW0cFyRjtVsReNu8rWkBD7hGxcICU30dEPinCEYEN
Syv7V6hP5i5f2iMAQiYwlTinqx1v88dccUntWQEe1OJ9zfjUXbqsmZzXF36GoKz8
R09+E4mlpJfbCsBiAJbmNM5SxY3DlpjJzXBYs8iD2DUIzgZ0XnhUmIO7rjHGfGKf
oN1lHec0T8YOK/Wi8+iXtN+lYP9sMuOikFzfGxzxy0Io264qhsu3MBnQnBVVeAxE
5v/wvtKhlT1IAVSsbJBvQdkJ7ckOPYA159ZrEwMmYUMu1m++InQYJOrYnif2vpq0
xXVTrhYC49f1/7gTSFCuYGmu205+LGryCk1/mXiOeL+VfDlHxlr6RgdtyyRV0O6H
w0rJ+HCOlP3oM71lEcUsQhTpbOgMdq+4sp6MfXLd6TpgaxXkTtwK/hGbZ+NrfmOd
iybfYFj9p+j37kK9ruABW5FvYt6VsJkyHW00DkqOJj26V1d81g2qWhJs11Pe8YdY
+SjDCl9gMXuAv4OUJUEeDCXwiXJPwdeiYBOhePRpBIVsdaTs0T0xLdFh1NPYuybn
QaOyg4V4eKcB2ZLOWE8GygdVhSaqgd2KNZ6TAsuELwNSBhrq5TDkL26VlPinhKhe
hvmduA0+Yug7TfQctwL8v6iBikFSrLIXFY8O76deIx0cAgWb+nHZKkt8l4P4Om35
ZwoTdNuyM6Npc0wNytv5DciRO+G5P7gUNreaok051xdfaKQ522o8UvMVq9tLfVfk
D8iUJRH7J6HmrDhdUE6idBzDsYlQalvGEYK3D3VH7Xn7bto7wpWPC2vc81Ietk8C
cIhJwGogAfK2BwqjHsNHRXEMlJC7/5lRZitcZ+fZYjuWqheWTZOmBYt/X6HMRELK
+fphav16RS82Z4DDnnf0Pg6KyyP2sGSct5Dk6mtIRYzef3PDHbrxBYGx1fOMunPj
4BJnET+Pn6gYharjVfGpfHOaTsk0G01q7DYoDT8bPTdPihwOAM9/wJ9FJ6d6XljC
JmwlynQGMKjzT5a/K9/najxoOOXXPFaTEYyy801eSn8cDZfqpHzGd92EZgx3exUl
66uoxKIxUtLoar7L67pvt66MqAxDtVg6mV/z1S9bYoRKSPfCt/ixEFIsmuv1lxZh
nNCYlRUb5tyQlgn2h0ZuZ/KWIn0xQCAWhB4ega+XAM6PM+cV+xi7AsWCg0tPISGP
sYvDbjbrLBdUBD7gPTcPgbiNo3bakdE7sgyw/Lp492YU9WgVQniyEli4e/I69K/X
WjFrG42BVFxNIC+GoPKZpf5EAcZHauEboyrYIiuQhTETtS7u0CHoHklJKtoN2KYQ
7VEwgUZRi0rr1JsTuSrptH6pkUAFpZp6Ml+IpooToWXeodfYEfBStfoZ3ZaSwLpm
IHIlK17rK027VEfQnJRku1QHDeETaXCTyp4C7qA6LfKXFZvGVQCyp5z+gjcyQsnR
8skFNFnTqoU555miJm7xD//CDB6vfrNy96Tya1lDrmfaHe3TCXmMd/yp6ezYeBTZ
4MuzSBYYTKzP6qeX/U0xkQtlVxkGOgSr7PQJVhX1zAqO78px86NqhQPOLLts4LLK
3atvnjBzSVZ03E/lvPiLGcZjC5p6KGx9NjUJBwGch6sMCn3UY45bbrQbf19mWRgW
Xt/fYo7cZvpyz9RqhPxwVbPCqKgFtfU0gvek54qNKhI+tODTzD2b/yRws0sroVme
tq0vw7YxT8RmOupygO+oGBH8d+JN1o70IdepYdfRDrwLbri8yjV6657licr35Exe
PbxVNOCElyWWxvSYIL2H11B93EY4GC57rxSduBugMObUR36dmwJi3JT1C8AQqNlD
EvttgTHWTRJoI90ecwuzkTXiclfliBbFgclVUOz+t3OlwsUqePluvPp+o4sxupUl
H08a8CVJvAToJfHTJ9KK+Hr782Sc94o3iOcOiPr3rC9yx7qpDKZKWUAPn2cecrcO
iz/+x/wKWco6RKwWpfYHbb+nxi/CdUWA54uvH/JGNIbBEc1CvAXrOyexVbiVoOro
CDlIoA9QnwMDRXT66LqGBml2RrHlIYO+hCDAi30WV9kWe8C2l3MciRpPr2mzjVcg
hMS3fbERS3LkJQ8SNCT8/iq5ywdmk58OKFVI/WE9PaTXp/XGB5LpTTFf8GkmU2Kr
EqaZuBhG+R7sioTDPqotbuylQhtU8BwCnrSmARzpxBoNy5XU4vvx4yUeevgSm67P
pyJ6gZtLEEGIiFi2oDeBYehg+xKPbcLkE0c4Xx2MaCk5Psscy5vLft9S109z6frR
+C99+AuuWubTa9m6HcAuot+kfff13ZXSOwpMe0+n6vLUSKGMn+X1qOWHjDmG/I2v
Hnw1COn/2+elCwaIW38GbnTr20e6A9U5IF1ZE0yYGnnFS1zalbMY5F1eg7JpoBBQ
F90tMWfkiHX845HBKhlwhVHVUlckiMdN4e9Xvz5+DXfy065vsJwzFFdOKWlSUJ4H
alGPtlvRVpad04hcx/nR1ezzK01vyfkpgkDZ8gvSzipldYFRuoIni2zDqFYwYDOS
OPAz+cbM3g4hralt9JvgyvNQeHVNPQT2cnyKM17MrAO76Dl4yKL43gZj7H9AGiKJ
bOtToqADWhPRFlrDmwHPbDxZVsm4FKVDgHkE+Yg+7J812jbuJHvUooGibFLeRGKY
69aBMjBtd9zTJmJf8IxljO1rrqbRdMtxeoPUlRawcn0+PBWLQJLFxS31VuQFWhbi
9fzgXT38dTRzyy4DJvDG/wTGHxQ04/OkrbwBy1jHPifnD1ChFa01NXIktv5qi+C0
Whc1Zm4Q6CBxhg5HGA8fh2cx/le+7NfWTgnoDS90eXTi7V1OGCQdJPSP7/KQ9pY0
yC2YyJhhfWas7iyuyNBw7xEH/bqr9l5wXOH+Yxci5eRyibnic5/vKAjbmoPYhfCT
InZeOeszBqJaSpquiri7R3mphPEv1gvhwVYdL5c0+ESaoboSSDQabNYtcMLnQxw/
fbCykwBu+wr1zdfghazWjdXkseez9QN7VR5BlNCFB8mSCWmXcJwy6lwJ3U6QPENS
EQnTyrH304HHUDu3+cFydQn5UFhMTat2FLiMDbVQHGX/Fgriect8aZz0KNDSDSj9
6f0ACKKt0TLtQcti7J/LEawoGUlIi5typgfRXW5OMv1cz/AstN8UFltq00TtBivH
s/XZOGEymOWR6tLbuSGbw61FHCQLSAWdInMAmsIzqJVhIaiOouJK7oCJuOluG2Yw
urvcGctVJPu5I3QQzv/M1xOqqnbT5152Pf7CW5S1ZjBbYfcYtwDYW4O1f2xSoyjr
c6cwtf2Y8o4fF0AaYwDcvJiNRQiIjbKB1pwVzAuijMuXeMds4/wZbtUO4wQdqoIV
NDVnq58kCRFOsEXYoBoXpSZSZlIlP4x0bHHNtRjVKJKw0NEBejSWOpeDzrJfGEPi
dCYZp1Zk9ILSjBaM3g3x12xfJy6RyOCX1Z39YNx0OTxFV4HplNbhASxnsVLcK132
cxqbJVMvCcFij4F+4Nno+HiaUraCgimbJzAfv+hq3V/dqiWEalX/m0JJ36qM4Xvj
5aLELB7BO69Bfka1D0GbI4jGAyvelPg/tTBkfhyeQ5E/HrBqyaQgykgSBQL9lzN8
Y/s9MHXWcq0M4tx9jUT4O5xfB/iWf9W8sM6H7jkHXoa6vEfU30O2mJbbG+tymSG3
2gNsIXNNlLYu8hFB32mYU6bsbzgFhxCsDb4VhN72w1wRZX1hKeFSufPQelXF75WZ
DKNt28LunIb3fgHsHH/0UjSZ1sz00Uxl/sQ2nW58u2Rtn6SSLVTAHYps3A+XRWxZ
YP9qxfsss8kzmNd/D+mNkFIBe0VxJWyHVm1NyTsd+6UuyQ5goKWUu0QSr5UjZAYa
wsz9nXKPjgT0lkmUOcA0b1AG9vvhjnth14D0rgTWVAALhXbUJ1ZyP9z7j75EInuD
2KhuZ8OV2pFTV+xIQe1lCXKVlK6BzhYkiGbgWz5x2fkTVAbW5CCoYG7HDRwU8RuT
kzLtYTYmnQpA1Owig2I6mhYWlT1rDthIbMgnJsZPyQ9AydGGKG9a7n4bNYGgyVID
rLnxScizLFTZ7/AJGvemIIUmj6vhNmVTirhzQYoU9lwmE+vX+VvhmieYqTuuG3b+
NyIKl3ZrFRiYFNoY2Nosr/o5BGJNr7s0WzMCOYFD9WXyRUR0GgAWLEXqrLMDe+I8
HrxR6HH4CCBxNeAyJw9utciFdRSCGQS7okUTOr3ch+aEmJx681NYIZ5j40dmqGq0
DglfAGPaPnmdfrQGniRPvIKmm1JxMhJNupaAaD0QvqKLMUxz94pCJOrAkQ2FjSup
cxY6meAcB0/E0nKGr0YhwFjGxdzEbmMOaIJgk73/55/0pNSN1K541rtbGcHKnp/b
0MdkKarvOB8aubf1xvIlzVU6ABVX9kiKAtlE0c3kOqp1mESIo7y0i/47v8EuoFRB
6ubAOOk4Fg3nzZXJptclqCWKIlacWYb0rF3M9mLqgGVcVMPEfAPpqu285Ok5e7mx
aRE4PKl+0W1iEMWni7kKWZFLXouNxjM7bc768QYNAS6dMBDywbxrSYeKTg43BKJD
VfQiX4NcTik9zcySnqm7KI4sNrcww95YAzkdMHIRHwHBNxD5omantMAf0Eh4pV5e
6XdkgBbowiS68k7+991kBlxH/JuA6FBsrviwtSRNqGM3XWx1dT+PZy1TQLaGxvZe
JNxGovBoHxAymdP1o/LK4oEOjjFwc46icwpc2eWEC2cqzAmdDyP0YSgRc9kVC/e/
0iVvrUYkTGEdPNJONzb0gcbiuhn3ruPEWwn9MFQugBZDThVfnSLuLIFLMuFmERSi
71xrT3qkHM/H9Nl+ciHvr1NSfepyOzyOz+IgX1ungjGywk4YCqaBZ/S8UNvRhNS7
emlqNF/ZuzvfLYV3980NNtsmJi3WfvhEJOs+tNEIJu0khJj+P7opqjaUiLWCEoCR
q5IyN/rja8Uq36a7yKeYnC4IeQqqdsXguUl/pi5iIbNbWYUMQbCFH6llj2LcHaTL
Wm68apNdHAwtqlsUOdE3sqQnF/NbwEGD6A1uz1xADK/wPSvdImuemWzok3kNg/j+
cdDiSZXu92vOwfJ80C5mNU2sgfHjuWGyIpuM81VZOyBqd2q/dNuu7G0bJcBzGbPs
P7X9wMuLpD/G1BDYMM4ZmH4C8dCd9EixHMYAdIS+Lc4t/tRkDDM5dKFTUrPWbFsw
r2HXRhJIcw+I0Y5ETIN9k/ut6LKQulgNn8N7nKpgIX7tYDaaomqgxdiELPofgkbs
HEIv5cPUTigswQqG+QCZ9aaHDUeaXpkP1+Jgdpaa7DTAVH7lV2XL3uxQ6VG3m2we
QpVU5sAjtzSs2s1aUI7FS0a1cXzFpY09HZAudQneXOBFmrQxg9EU2lTCKvjc0M/8
rFr4etQKGCbr/366DXZq9X65JS5ajWJTHmh4jBt2LZsDVvuLXlUzkz4xfqbsMTLn
laVSNEJFksCgpllf04HHMm9ziqFr+dIIn4B253XP58FLvLTccsYOEC1enaWsJpYK
hIFc3G5AIUDyy1g7v65O7s5eqbA+xYoop3eC3+8rYw+BlmBRkF1Swoo9LSwttP9e
fs6GjKU0o+F/ZxBtuN0Y2Ho+OlajKiP3t5VPUcUnFfa8R2eSwMcqNdnksmC7QZMd
yH8C+K46Y53y2UUbBpNor2wtNbrPJ2G5dC4B4xPSmyN8gba9o5fAOV8OCMEIyeyq
vTWuBhR5s/xgqI5O3DjlY4LCERxnBpDZYB+sw9McS2vOBixwHOomezYTjX6jSUXN
oYgtBW4Bgp+Qu1eS/PpG/WQLdwAp6cUj83EoO/5yLsO8qZjbXfyKi0vs7s2VwMcA
tlSjMb0QikpNB409AawaUg3wm/QJhVHrv1NAO9PWLPD8Lc0atIElWKHngaJ1oNj0
d8RmOwiTSZyyXBwTaOvPt3nk9wJIFhkcND6ELwNXP6+S1Nuha8Be/Exj98cQfU6R
o51K5LdT6UitZzZXVrg8aaN54x/MenYKDxX6o1OjoQQpARzsNvQmsdibfTbOIuec
2ZDQvm6zrJ6W/8RcgKsy7dLwywQ7tzv5EzX5m0GMxUQIKM+B+iBKJ/UiprvENAdu
HucewQZakg9IVCDGm5Wwf+woaAPAD4cNT9KhqKTHz+G33Rtb3C8lYuN7Xw5hOQ41
HCx30CyJYEkg98+3Y+SGwv2teH3/Hs4wWAh5zr6lP7YvDhnHZFHlxXgvndBZiZJJ
G60BngJY/WDWSRDNOEFy1FuYt0xFX13c1CXEARBaMZ74Yo3xQHj34WgTnolmLDrC
Qn4gLKb6MKAPtZWXzvT1QpIRlzV7ns//xAcCQnPVntv+aWlkvLyUROgPX8QpMkrh
L1ZUGUnEPuSzfe05QfpL9WvlDJaQckuFVel5/WqujQsYm0EX3oWkevDP8zDe8tfN
J8Necr82ltQjtKAtYeQFiyIuC7ktNSILUT/SgRTA4enEfI5M/N0UblTCwOxWFQZR
Bc/o28Mrz4oQNHJ6KKelI70zxr4z3tlmravbgUusZ9fOgRqNTiOT2IRXN79nxNQs
aRT14X6W9NDumdNkREoUHv3hoe6qKmivf6dC9g5tGmm1133yWlGGBZPgsSk7Spew
VILPWiTVG5TFwWkImks9ruFNTpJOa4O7ZGtmB3QU5Py6/U+pyL8J60I3ueLtV4aw
Zk/HaI2+lkf3yIon17Kffh9TRs8B7ssrElSjOeFM4P5mHaMQBWM+uFS1NFXtW9Pk
x7enGvpcbIAfsroVeycOVe8zxJecwwJ9GTrbkGz87lXG3aWtOBT+2BeNtJuOxXzI
KGdjcAudSXR3Q5DX8HXz8hEBus/qINBE6aCGVXISoaf7yOkEr4/AA8uC7b1FRZ+d
bTTRIQTpYzTBzeY45oubBQ6p7j+mIjtxtG0cmN8m8VRE+0itySV065Q4QUwTuKhS
Za2r1Rnd3EcY1EqM4RbCpZxutf5mDhq07AR5qhegnDCTV3Xon07vRE3zX/2pxKe0
HAX8kerUK+uTd4RhkVQWo8Ito7NPLa1rXJ3rk+mCp8lR/RAs0vbS3t1Ej+LIlEEB
l94XotS0+SUiuAjAg8jyHrQ7uxo5zDy8CcsdzE1Vglc/OoVMU86WSU+BK2VwPa5x
vzuG+AeSXIg5bH1OB2ElMGWNadnB2M77H+tIVZ6ajnESGbPwPpicjaAuPcwOdNin
fHsQ2Dgv3rzLpw9lkpkJUFIdbxoO44Qy8XcFK7GhdsK/eUDgtMbSZR/IiLvtE2wN
p/stF9VznBsL9WQoPD7kJGIefZMCcSJ9HrJy2J0wbWTaQggt0coOMbXQnPIYbMwM
4iGKxSPg/0LzsZODDGD++lupstKu/QgoSOm/j14di62NHoXCi2gh6s3sM5CiZNTD
KPhDo2dKcJPDWa9qvJttRq+9eDEZYaxYS6HwADfqUsv+AVVtDGBaIpUrK2QM+jol
ZJev44H/i1E51sR1yp+BnmEgItIgzZw9IJasOiSTj3APVkoA9zw92Jo9kC9wD9es
lV3mj9WQVJKjp2xsNlCaUW+xIeX2xbEQJALCsCY7Sfx7giOAzgdGn5CskbFFK/WT
31FAZqrb9sVYotvLjxTtDB/jBkVcLk/9uF6M2ZuFyyjJw87rZAxIdY78DMGEjTO4
KU2SIfAelI8XS2cQchEJRdErXzYJLAva6CzJGhsADYmFf4ueIeg1oIONdLTQeLkM
COJK9PvxB5noxrzzed8K3Khfb+yKf5jzMJRpNOf/nD4+xF6OluAAPUCM2URu+E6G
FT4U7fNb7JSNp/U4ZzAfVoTEqH47AOhC0VogFsQADOPlrGTbCVORLH36qAecZw2B
gBEpfdBSnil7kUDd6iKyS2WVBkHrxiSuwoCmyctKMH7Mtfyq4U4r2eIuSqY1Wd4y
wkg5RLF8BuHFKRVf3eNf70httrCwhPGhIxfcamPGdvXxKU5fbE3mpiHIOTfQAvSB
I172urhaS1Cz/tK5SqEpCqhGxiX5Q7Kiua1KjMlNeyoy+Gqh86+cZJAHngUrDy8x
nPTWjgGPpHefQIHfP0L3E0Us2VjnTj6UbQaeSaPhe4LPajG/atXKj83ngrtLLr5L
94iDk0SH+Si4ktBJz3qEOXcR9U0qEA5eBph4SJ0g0pmE+NUdCm15cy/OJTsfrNj0
GGrlY4Njg1WKmj4IiJhmyh9BKpgRQaRXcMhQQc69vrmoko/CvpFnu9O61eeSm4NL
y5sKbEnn2zin3C4tESyfHN9qna60E7RBDQdrt8l7v7a57Y+IL7Bvfl3+OnWpR9Yl
TibBsDoo0XUIwhNm0RNhC+q8tIxmMqqE1cdA/b49rWng7I4UyhF0IGPcpovjgo1c
9bFqYc2Gp4EItJ2lP/WSAgZLQqcvjAz91lKqypoHo02eUz1pdCwZKWXFM5cd/9IP
fczDC8e1uxMGH0PG8kpLeVikmIO0+7YXYV9AKh+lrKu2yIX5AjXNbMbOuGkeOOB3
XvEagTCjZoq2ivSb8dulFqJCPZikdFv2IX20Rv7xEsWcs0mE69AX28HvhHACe0o4
ZdmAOApQF6yuWe3v6wRFGcb+MjpxsJBSqF0GnTtfeinPbQYNsDLIkN/ZqP+7Apaj
iTAVW+uBC3bdlla6rijvzsaSppj5RIf5yo9suJOivheasZLpmO2LsCl11Umr5pEg
tpi8iyyiDhYAVJHlElEPm9/IVCg8p8fH03m74VYL2zL9em2a4O9JMlr+PMxBqLuY
djpjWOUObMPYXk+vVTQBJDQAOD92NxT6o+aSqVOcuMh67FRfTbDPoUFI22wbgYgX
DAT5KVAJ7xCyf8k7/xRVouXLmTOg4ITS8BIe5T8VNnugW7BL4Asb4+I3ZEnZ8R4i
L3Pj4S6VYSWl/jyTUEZCtrYCXlt9eSkaoXoKhPxbhcMl64j4EQMFuSMpt8LTE/qK
FKP7h92DkcDCj8fBMLFEGE3gfLoPGOzPUmKvt9/tx4K3Zx1guyopl7aBtkcEcdiN
bBuDQw0VKZZMMi6AmUwhS5xGuhtmoF3SR4UOlWu7fGYdE4mjkTT5kHvAz5cK/qOD
Pc2O5CS7sbM+wDdAqeD0Fwlsdq8hVV34J+5BxaNz1aIlqFEb+B3Bb0KXeZY+jUKw
AaizunoFidPOImEsF6ebjyfhqfCGchKMlV1pwPogRMihAnhhGleF/rS0ByCcv0m3
V95UeLnutq7bVI9yQQq6l9g25Ai74tBbXlv6at2ZhQ2zxt7xE3FFjrB3Lf8VuRvT
vJ5H9LDrlWMZTQo4GeernxIg2CoF4oiz8qM7P8YKVqC6e54usCCzSoPNmyVbYwmg
AIH2+LSB1qQ6nE6TLIIxcP81ja5KlMNFt+cfcJKU0GGdvbcMvFq5rTQhMoRorgoR
Y3EOC/LnBnxXVlgpngL/gSX6b79xxvBHUzZbQGPUjhvSBuuG5Psj1x2UiFR3Su2w
59kGMjIOdWVNOaz45vtgj7PxOuxkdGNU+Jxq7tb+rP3vF3s3h+BAXmvvZ6+9CZId
TryLO1z2Gnj3fKWlgg1cBbKsKeO4IRK5jqqSEFwWVaZhMrAsUqDB4NsdOgv5h6c3
BZqLtvHOLEfLjLQALSDdnVgRgSu8wGkFtgtQtHCgiKmZ0KXxnswk6CMWv6itwu6J
r4jjyEQJw0Z+SR93zRxGfF/lOeLVVwlFlRMbFW6+NBioR4M4ueDiVJWxed8GK3qN
3MMV1vN592hB8YnwKZ0Ncp7xHJ/C4q3y8qlbuqRzMo1Qv0v3w2o1pm3UcSBAoJc/
cDf43o6w3+rWPs+LFFVnGVhSfAA043hurf5DDMxWMSMcJks+80kctYDQdwSknGYi
u1FUbnA3BHnZlBw1xbBkMBgOFG6p11wwCPKBfLLAGWDU/3T8iOlEzgtPsEwVqJSW
nNAygeSuzTloyoUYMMi1D3DfxL4FVSVF/2SoqECoL9BdyJ7H2YjHQTsHkIpdzxtY
sgY1aj/rwuYFO/bYHBOZmftzqlrDTbcWOmrTI1BAyhO/qHr864EGAVCLi81cKFot
wlexz4OlBC0WATmfulPO4oJtrqdBzmoh678Drseh+urI7EJoJuyzLlnjRSa/u9jd
No5Ir4/VRZH/EogTHwUPfA3QF3VyGZAoSgiAeZuz0Oi2XLxFTO0cpED/LmnkU9wO
gA2QIUMkPnv2qLNyu4ZvgFSj+3zPzigHzTwVPyS+o+vozWu+lRBI6O3ZjLej4o/E
NoZJW45VBJ8zVIhmmEHSus18a0U83oRpi5f1wWICcxEzRGadX9OuKrcpx/w3ZgxN
/56Vq9JCBVKn9GPt6ipVaDLcc/VxX5XMUw2JRD9BAIlJ+QRSCuXJfKKIWTDX/cBc
GhwMGMwFhqur8P1cfoEACz0GoMNh6I10/wHRv+4TSoP1lLetT0fCTN6RXqAAS0ko
xMqVgSIoGX+u7y0tEMWqIC9j1HUZ49oBqP0AS5GSEUDLDXfkRNqUndroMIG0gEJa
MKOq3uZ4ndSweS0BkoVMyGqPtUp1tVtltSSupK4xPkj/r5ZX7dW8w8GSWISaS4T5
Oe9/MNvRvPkRsrVptsPn/yltmcXBFjQofmJOWQZYR+d0w3h9SL3kYAeBB3ovpRTv
Cqmcj5rtdOIQiBw1Ugg8qi9wjqb1pCJWz7qlVcd4gGsjjy8D/r3VbF8cMuEEdJLS
FL4gFQelgjc09X1ITmUmOZR4y9Yns4JOofNx0fklg6niVp7iMp4oBETDSs+p8xLX
U6yAXcG3KuivE08OOh8jum9pCMe/gNTU4EzqEOFwhzurnCqr7Rp6tTXRIrfk1THV
sWszv8703a1AN2lMXsgvu1q2g49ZRxnA5Fq5F1BBl9kuW+rRvjIbFMxJKd+CdlZt
P7EpM3ooHBk8mNJ33lqs82fbbbhTMuCszK4FJuHFbNoTzzFrnt+cQGPCqVCsWdDr
D7HfwS3Zt2I5iCNH1zoDZMBFqzz/1OFjbA+9Gv4Ie7VSAuRwBM++XkRx4HEJGFBa
ZWosP5kTWS/T/B+FvMQOITlD1dVXlm9IMyAw1NbBVaPelrh9TSSQoA6Gjf9qNvkn
mVikixeCJ9hxX3KGo3x2MJQYrVh0WZ5Sb1x4kb8GwIip6PM8/awtIoHC5rjmmYtb
JSKwPBP50+C/xaC2IELD576kELXw8Mhb43xKKb2RzDMc1koiYOpHvgkKoCTJbyfm
3nTV7ZoSFgOpv/XqQmM+N4jnGKK1RVLzvbjWo9wadANcw/UDWKdK2VWq7w1kCxU7
EUSUDlklT+LWfvQug0EIwge8G4QBCOEhWUvqoPebnyOo93WQ0C/xEDkR0bzU4Cma
jWfYtQPaWGv1XyIyzLWRSFce8fvRQLg9Ch6PjVsA86LyGXixVrHcQleUjPrjog2C
ppwKLtvcDJ81SFkfOfihrTc/jkPoTz1dH1U/DP/lEELwMiylD1Y6iIMCUlFt84kO
289C3TMhYsjNO5Ebe7OmyEvVO97DDErYO4paHJ3BnORVUxWLY4sgf3fkfk7h++/n
RzQ3lfKw3I8pj78dMsgDYyM1nH8dhXeLdYnQfL4NmidDvV9ugaxWeua/TnOWsIbs
7UvxZey6LCr76gZdudnIv+t15SVaqfwFLAN1PeAs/UzuX0FVL8HR9uqsuLV0AEcQ
19zj/AwIWAWkXE6VWu58t+I8E6NapQdUOE/9YlEbd4ZO3CPOeYgIbOlbbw7/LnpF
D52XfCP9u/shvLMp3RdQ/2wOc1noX5I4SXG4LcMmE3Ie1BYInkKxdjYlVgTRfK7A
AGKr5AXrgSA2eX2n9gDwl6roiadn/guN6yxy7cFOu64NXl34worLdBSExlrov5eP
QEXwu2heN/wyhqwmeK5HQ7c+zhgwLuln+0TCROfNhgndpYtVIQ84QSbFftf1LvqZ
VKWgP74Kx3xf6dR37ukRCoWTfY7hYbbYzWH++h9lXHDRcCr9+Cv5qvNy2RGlAMdq
c+/a58gdABSVP4pm2lUPVq+lvLxeN+4oZdOV66W6Oo/ybTJIa3QeamU3JTTsBPu7
2RNe9X18NY7sBK95Ea8lAUw8LY8ZEJu06EqiiWlA8sb9wrC5wPH1RmnhFnq8UbLd
QB4BSecLEKz63tEMgn9wTFlMJAx3898ht0e2TeT/2zZIZ0rEcQsvC/C72KhJ3TaK
tim40PYh2uJWpdsiQV/Lz8oMVXrCnxfRVdE+jkYC5ZfJ6WwVno+CUX9Zqr1lcWbS
HPuwWANzzbLlqZtVCXQfeJ6KCltE2OjqCZgjmUyDJNoElrufJCGGVvmo8oBxI3Rx
BtnUk4m3zA9MKdzpmC7pGoYjQgK6LorNmteQiQlmS/WLUbr0WbtFogfAKwCincQ4
kShnRoJMx7VuwjV0ov6iJs91ec6F/PKiKRqJIghuvYCnHJidFBCbrC2526piB9mB
5rFM8M7elUEWCFWdaQ2xnPRQxyU6vIWDiykFq4CuwdRrDxIZRjgJ8I2OtikH0C5e
xpvLnUjVh/q/+hOijNSYJoXz7WoExCfjdW0IGSiaLX3IbPLlC9/d8R77ro/C/2Ts
7sf3QJMaIBnoKGoAWaMjeYC7E7TBo0z2GcjffWJZLqNDeQpC1f5hry9+6+khOi9/
RlqIZRd0iDJuCPE62Hv78aJy2zLSFeV8BtJh/WyGlAjMjnJhFnqXv87J95c5oh1u
JjdEFQnNnt1p9ihY8GO3dTqW5sXz4LzqEBBWvCxcjtiP+Mqcypk8M8JeLUsGy1fH
HGV+gNNsrE0EVVqxu2aOgN1YHbLIX3aZw4nr9hNxv64r+ZJqM2JAPZN+uoR165Tz
UByESywWKW/ddaUCWWe84gjWsvLGPLcTaaH7kNUvNCncBwHkB1qnuKeMQ+Dj9rWV
A9VqIi83pKcF7jt5JDmA14R0MRBtVwnJTRKTOBWJ3ayBqs9PQ4jRuveZy8SCzlH7
AmwDzBcNI7xXxJ10Vjh9QS5HTRC+REp1GK5c34luy59HFiR0BjgQrO5/znwxRxWY
8KdZChpbFcCS+pL9ot7B1RnLfH7Pi6ILINLJDIwJ9Pl0EEQoLREDetG72t2+OGzY
5JG5Osm1S371a3pyB+O/R0UNKI6Dd9yB1KPpFzKFsN5XY95n+DZNCtZLZCwQ7vU8
/xjADOfNDvU4cxDw8jvYQBhGvF+WJe1ONjkaA553jfWKaElDB5bM6BXzfeBjLBLu
ETvA1aAblrU7p/13+R7iFbjUrDX0/2QhjUnf0UhB+v9Qs+xTw20NVkM04OojFQDD
u+iJQxfxwuqL/cFJmXNBTWM1XYaYLIBEKy9mgJbjwSqI+WFvzL5vn/V6ZeYdxNrk
uHTiS2Mf8ORDLIrsIFMpGQ0MWeSKxfWYCeQZUlhKi2tP9SyTw8OAS2T7d78lj/jQ
XelEkLFudWorF6vpyKjnp9yN2Ekx9NTJ4bVH6GUUw3L71IpA98mBAbHfqdpBLX1b
x03krVmw1CATc9ojFTQhCrj+psCsFU7e89VYX4283rxihMZSUcOs8+7Mf2ldsUJ9
gSqLTBH8A76hMSmB2yrBP6zmVGwOXZ9mmpsL4+v4gjr67Z52fMXVJ5eXtAt1OXdt
4yF7PPtFl6Isgs6+5zmEpmOGviEJI/wS1LRZpUw5tHNU0clMClt5A5snA5Fz/lSY
TvUV0xjXcZRPnC14Ob6tY1oYGlsYZkQgHbNn2iR6CjYte0qoX+GSAa+DeFBOdq2c
5ScJE2sKSrZmjj8NHHYUGdZRUNZC59hRCmFlhvu0q7CJ8XUo/Yrn41nI3cz9Vsc2
gi4z3WpVb3KVewaATHuPd4dOqQJUYtChLQTHcPGUjY3m1A5N7QHsM8an/Or5FbGm
tpU8OLqYapXaf848U9bkIZthwFQ3up+04sE705VbK+JV6bPP8IAnbNOpjL/XDBq9
dCmyQFHcL1XxST/qiGti2pse5xfFFUIHykJy1OwKLwo8HUTiHy7JuFN/isZD/0Cn
V3UKk4pGQioUj7D7CX7XZYBskftwsoEIb8uVigETrUrZZmXz49AS4c5UClYV4SyX
srzLP9tNFebPPvnBCbhcdsXvTIuAL9NMM9xvjUto+Ja25Tx3Y7Nk1+BMX4Nw5H0o
qqdWSs0X0LH0LGPH7b1zA3SESrUFcv9BU76T5S/nH9/r1ksLb6A77Q7QZLLiwr3A
XxpMj8Dc/HBayMO4b+fwS5QIT1dXmDR2/cqOVKtKeyZPUqwY2xtNUKUJeN4uoJYX
bKnKZoV54OMO0OY7iYx6tu33C9xDgtL13o12RRxjkHCX/pnCi9ibgPPgSS7tDyST
yswkqKR7c+jfjXTl7N+v9d65xsZPHekukev0V6CmdNb27eGGMbizQpGwt7E7Neg3
d8HfAFiHshzMMci4i99qbfYV0Lmnu82LziMhN29Hp8Q7Z3KVeGHXGt9z6u4bACV8
i5Xt1pcBZJoHSbSpFXPu1Ye5kKpwIMepuD1dCZJBoK1PgNR9yk4WcP8i5gRR4Ma6
wNQWDUyZiqvTf/YphUh/5iR9lxBNdNz+AL+GuAEIs8lbZjgLDX1Ld5N6qZoguMJo
79cw4hDQYqjIxndwcj9sg77qzihyXbGFjRcFiTD7mP1Ni8+uUaVZvB+zyK2ESfif
wo6WYR6yCi4Ulto57vv4V0Lsj1kqSq1tR1LWXiP9q0YTbmoZFZTk/+wwESPJ71N/
f/LVEKXQkO2JGv+zA9UfE3dCMSyqGWhViLhPsfUWP3z7vFzwKkEKzcr2qGGL2BKt
GOH60qtYMIfONSvQbnyGaF7JUmCC9cnEUjrXqe8dt2RrZfsYKVmIy9EuMB6gRqH7
yuHd8KUnq5H7HisAbAhakuMoU4PiQez9I9kgkTNpAX4fX67dc5cGDLHF00N38zFT
qkhgSF8HGJZv4P+GBBsOK9OzGlLSI7jsxZ3WoCAwIeAlYtRmVmJF91uBiHR1op2o
3TVWls/Sw3iAEmrCKHUXNQ2dYLfXC6oDKUL8qabvzpJ/nVIKXW6kyrJv9SYdVBMb
1vuNlektZWpN0zPDCyq6lBrCUO1vOlZVHx9Koevfmkr4XE2iA6cwy9BF8KSvdxC/
p26HCFoUQpPBzQhSR9DHoW56JziCuv7GgFaFhoF8FA/s8ZX21H6GENRsTddVACkG
UIurScEyocar8FcpV07EidqHCHMpggLFnTJo9IoGn7NNLVsRzfZzFZ440BpbDtR2
Vz0Yl9a2VOIsNHppGtUEoDRCzQmEnNb/D4FtTARubmz45zumoDc7qlOzVwVP5Nq0
jB1V99SwLgIs4ZKFWVQ59pzjBogZBfDQ2Cz+oUIgklM3KMJD5i3OqtoIjH6uIhva
mckkE/WnXA8ml3eWM+Uc1wd9iOSVx+IoQf5WLtYx3FdaLvxgFd33q4Z/+gexR1Yq
rvwo8nT/uAZYLrzTeC57wwxFvNP3lkghcz9tVvVINRaUNygLuN6THdQnAcbaKoLj
0rrZlAEWwQNkFjJScV8PDsdVYGe1h1znAhHVIP2XnQxOhQ7ppLuW1mcvqE8PPcpY
1RZBzvCFjQnQB9UHbsN1qd5s6PoTGo3EDfGkJ7+ToYxzmZ/qZJQe2TQndlVCUuAO
soR9XYb0UaNVX80YUILcFHWQAU5OouZ1oy+RhOHtdRUwSFr/8wGHbmzy45V0sqwo
IO9k0q+yHgDzseokYKpwsfDUA0pZE2RO11kfxdnKE4x+r25s8wuaXM6p4PP/F5fi
C7Rd9+PbGWV7lKdqPBS8ut48/AvZjmQdeB/FYrpZVAoHwnAUqZFqL5nFkxW8apEZ
VZPs6AO+S6cmLlbTlH1d+BlqZKuKXe6JXeY5ltCmzNNXeq8k96A/2CLVcu3xbwkm
s1LgpJOb9LVGAnRKlPQ3kbKWktj89DrgJGqdiIzuDxtaVlMtTVOz1y9UBcC9JGBn
Eibn754brDk1akglCsFp09S57tDoKzgwLkQyF7VDkMY5v0josOL9ROQZn189gRNJ
y8xymMeRmD+yhELhNzsXlHO8MTSmocf6NuyzerR0sxkShjMexy53YmLpgntthqvd
ZnL++vH6UHIlCHNf4c06XGc9PQABJLJl624oeqqQyu85i/QRWQ0ZRUQXdRQb24Tg
QG9CX6G423/SpIraUigFUR9iG5CqbkuarpealZQpu7cuk1+5MzYrnteYzR/3OJbt
y0LFryTQTmQVe7pKVYE3EPBpsixtq5wOE3EXBVFz4KQ3+mlUo3l/jl6EgP5E1ixp
loBh4Oe/5tEMoCS1kKGrwJYVMhvNu4QiRrsGCn/DdLXTv1K4MTQ+NApbBx9uekAu
9rjK/dqNHcJGaDDgSkk5nLwR4dh4CpLjgox4U4mKPxbBhwkAjfGRjzS8COBL4MnN
XppmQY0CEje7yviTe/+oRAhkZrJe1m98MoD2KTsc5OhnhycCpGY4cjFTO38n8Ve1
Pe1OwMWIrz58cyFHQ51uXk2BeDNyNcx0sYLZiHzzyMWX1O4g+cYy6lSMccbWViuk
KxT2sR59JZndk8faO7fV2lyGii6b1/w53wkNGwLEzrjFwLC7KM2F+ng9LOLHmkjb
RNwzqfxEAFp8F3U09fIu3t3poCjaINN2eIuSV4Lib5uDIEbBH8jBUePXA3QJlRLw
W3/fVaLSUZK7oKDDwbZPTFMGVtCgIoyuII28cwiFr6espA6Bd+tgkUJV6hMh01YH
45AYDpPnURoCtxZf1WZYAEJK4fnJwCPXXSG90tdfg19Ih0SfntRA1QdJe13t6wdU
jyDIEzbOPekR4uHy1ei5V+oI2PAZanypowAwxgECvwVrz4keV2JecToSdWyMBtcI
+Ku5frkjX7gytivQHSjOPUNua4V/d6qiBmxaMkxAAWUboT02Viy9SOgAXeMM7wTx
SAoHCBzogcu7I7MDjJh1KmB0nJ06jwMFAxkm3PyuwaZhrv0WDQN0Lim/ykYAYh1q
JjJwS6mSvgqTgBrfiJKVtKvWxTbhubO5YHAlLQLZFEKI5rXuK7LMY3p2TqisvDBF
KkTkNcvzwSul2nDA2o7GdSpyU5irfMzz2pe9WbVn6sKUtMHK4l030ahpNuMcaqJs
Gz/5PJfqZZuD5DTP0vfcTlSgBZ1TPl2+35tnBOhdw44dW3zo2qspp1iRom4zlOrV
Y2fTU0STcLmR7/HRR+xK+NFjURgINjBtPZlu15Zg3yHziRGH7qNV6GP51BY3AIbj
karOe/I3KwBO6T9uiUKkplnca2cmjqkMYiSfu70vksamIWjSy3s/yJpx9AXGHG7S
q4aRviKmVWAjzIW5SrZ0dVhblsCDG/qVeID4itAThNoBtlvrXKWNaIKj3uJg2tHk
C06GCSZe/8LVEZPHZA/1IVZsiETSER3jLhCd1/KsEuW1gqy1k2FZWWkC+Znio9lA
9bRkWousk2spyQmgf/mw8/e5P/zTtGY0sUr37RConG1tUqRKoGemz7Fbuqz827FU
WcmgzJoPZcPhe4UzVJ4WdNozMqFMzuKhqeidpxUan8fmrBmjnVVk40m/FTQq6I8H
j2cxTAypZbfCukb2xRON3mz7gbCyBjSHG0i5S0N4eHUxkPAtjfEh5EIYGUmxYHO+
T/hRQTJ/W/JCj+jD/ofDOvmzFEkWv7OiyDtW7O6t29QI2v+/gClT8yQ5Aa80x657
K0C2e/pyFzopRA892RHdJdNcPhOqyBkHqrpokB0PlpVgb8zdQPzEHirMWEgAdqJ2
ZT3/WF2XEkkKDADZdqmfqvvUrCwaikpdxtSQj1etNmAi36yEC27KwTSBUz/tG/ZK
CLCb5fDWpHYrEtC3a/r1xNvfB4fDa+0rx4akgqFU8a144ngihJBJxLMou9sHaMY4
E1/1gKJVR7i/XzceJiX1fgZwxGYInzJ//qmqf5KG/rIc06l07NTkNU/p4L0sOh/7
M13fP59WB9YcVcZpy8uj6zf38e0S8G91Msygrk1S1vmSEYR3iPYj+Zni+jMl+8oF
8hDZsX6u8P8ClGgoK2R3EypAa5EiD6qoNrSerKGGBRN4vM5cTYOXlawz0cSUZ3MK
OoQySNrVL9D/RESXWT4n/ZefpkQJPkann8AncH+lni/tJBbu26nUoWiG3B2wM2We
XUHAL4D3bH/tGFYNe7aRmfdyWc65ueDZCTV8p2m19oDiCd0FrihLC3NFPHGKJnmM
AtVBqEfiPJKPC/exC20aF9U3ynS7CJiD1tJV54GfBtS2Ky0u1Jzmk0cfd0uiCXKr
qhcbtuI+mA7n0fHIH2xHucRo5Z4K0vcXGdUC5vxiG57ZjcoMg2bDGF6gzArIOjgg
H3QMW5XCyQ9zrlA+QCGSl14oMbloZWG4BL8K0RweGeTzZcDSl/5YgW7zQFxr96Ks
KBX+i58rTrBC6UDfTxv+CjEW2ablfa8MJZrkiieoOxViGD4Snx/fWHXtjjv0RQTY
jByddqH6lemH+T1OS5E9JcsBr3L5CRiOkAJOOhqAOzofUg4qiVawx+bU9/HFeVRE
Eh3bvM7yq2W4S7/CdzYdaDKmpN9IZsp9UYhOw5BxmhvyR1IwrlQnp4PDVRDOyrvG
D/EPXcybvBtwYoLfW4u+90UolgEVngg0SOdWRdaZud5OfCGspw/tbzgmgMiX8xQT
v6jbkI1pjJ9RdggtAqm6AULE3TvZTXU73rUAv2XmcyG0enGk4aKVy8QNW0e6n8NP
n17DOEsgUENjKJjyz5sb9lBrt2gOPECCa96NW41mfTHdieoVbOBX88cmd1AAPvUG
CAUDP/pI/NOX31EG5d3mTIZR4KP8o3mFdYnqIO/HmX9N4cEYbvkgwM5l1RrP1TpU
9BgL2JKnuoPCzAlKgc4ckB2+PWrZZzu1R89whqX9hIeay5MeDouhl/dgTyeEnBVw
9TJOOJBY+dy4fS1pfG0yEaPrTkdEqm3cZ0UT3HGbGta0cIQBGiglKwXhjf9BOt6J
Tz5gRgRckxXA2mtnh5MXZ78kp0qYL/5slsZivs5pDzdVa+0wmoRASKdYNL6dZ+C6
rE8OGTULDow1WRHN0i8PIUXmZ2Ph1A9wTu2vJB/fU4l2qmtglBnGJ7uPXfFgq1Up
RCwrlckTDhIH10D+vEMXK8CLukleHyg/Pcpfkwakk9WFfGWQrhDEifLD1OrLq2by
odcqlvTU8i3lY1tMyOgInfieHGApxEYP7Wf+9op8yTx2c/k2wwBnbnlUmR/0NlWT
gggp773wAvPhihX368FYNqiY0cE4ciEUhJxTggvL8av+sDUEGkYewB82tNNUI7dp
S+ewv0fMOzgHHG7HD3SZ7Vy/yKmJoXNVWT0wdtkTU4WXeSltLacDZ1kjhXEsbSic
6K7yKm1yng4f5/iZdk1u2TWrZ5ssRExm+ZytHidMg6fUMnbcBL8duXghwFWWBUE0
OLEdyQf1ZztfLLCO8puuM3c4Mdds11oVV/2gaKH1CkW98TVBpPG3ZOVpKtBISLLU
DqdhXTWTzwF1jqhKviERy3PvdIf65XhFLCfBSaOn6Sq9dKpwhJwEIpHg2f595Nt7
ppzhgo+awq+bYaJMVsnppvoaOs7j4w1scua6prmZAGHOLlCiU+qTgZmLI1cG1OAD
eleHco24TT9a0bnVKt6DSCFymqQOVpbitco9ZlJ+yjvWc3feKd24uysCeaeY+qIj
hwRxiQXpfp/tc6n6OdPHW7SJil/c9YskQy3n4qguqJaus6J0kiiMQeb4U8Corc4o
4SOkiZy87MckGPoYPEmbgTsT93iLmcS2vvRj5y8BEcxOiML4uyQQhAd+gRHnTdfK
xXSnx6ExEarj8jKbRsrzbPMZc+u/R3zzgBpHP6DJZgeIjqGOQ29lJaVwy2Q5S7eV
Nw3fUDC1Bs8aYoA0LebNtOd8wSfa03yBUVdHs01OhsWndyIvkcmmg5CJdVsF7cmq
MPF9OVZdSGZZQsucMU46Md1AIvu/3EJUI/3+xOzHjIFKET+wRaQN9cWFTdPNEuqu
zlu8CoY+BJbA/515RQkeUADpbBwAQC2ZRVb+6Dt6/6NcuBjdPh90OAEsxiOGPgrR
nqQVSGHPbRhQo/UO3YBtVu7gALt9I4L87ofXwN9wNlH+1jXsvDtsapUjBelXUl25
S9eBJHz191WJIBNgoqX8aR4vEm5QOyfAgUOlb5Dk5CIukP+mS+0+LCNSCwv0MiUO
KCJuQmN2wyE+m7OG5nCldfQa3OUqrdER8DiCqho1IlAwMVZ+UV6Aggx8SamhWl5k
6nXujH0vFwFvpXbOO3+0zC5UDudwneLFCTGjMS/AERnfeIBdIJYnzn0ZB7ZgFkE5
+H8lIKz9AE+azUtQxvZwNi8vg0lGZYqJPXHqcJdNSccqWXY1YMyuQN4xCp8gcOF3
W5rXZPvr49qDE9C7i2+lCW0XrCDo/xu7QDMlU+gX7cxF9ICYV77njjRv30qddstx
lt6gZ36dq4av8Tvp0eRVSnJqRUfcoEcMmS+OQMgi/pE2V7CHFjlCwiV94BTTQ9WM
UV4WJ9V1hpRLMH5bHJVhRPRCjFs+GNdINctSWEthHwD4+I6J4ft2+C+gOk0xeLrz
iVSwt4MWg0gB/QbFL8E5aQ5ty0Ud9UvLv/LSm3J77PbGT7y2XWonzzc6W/49qied
+CKg6FOz7r3L+fHud7s8rC9plLkNJ9au8OrXMRFOd0++cncqAVB7teJFUQTLWE/k
a7qbi4Lf+ETtPYS+/mFZeHEMYRUtWk6bVfVwRVwllGutS7yhh55+ytyi5ykceQ8L
TpUEcW8zNCJumR8Sb1AphjoJVCr/MRtXTUZkXMxEkDBN2e0bgFK+6PI6n+vLvLpP
giZNoMzOuoWEN7MjImG7C6D8HCxWsdzJu5Oxs2cVvEJgrSNdeIoqS220TrYhQ6h/
1nBE20g4JTb9EYLMxx5PlIZ6C5flnh3cfUlWQPpC9pM+iUGtTVexOvpgcPRDLLen
iiWSg1YkJNN8itg2LanrqBf39E5iqQglp2mP9e8NGqKmljCPf66muZpRxizsIclX
Q6PXhhRviY50yAYCGR4FMihOuk5Od0JBZiCs73OYU1XE4ZQFYsKk2O85YeoqpbUZ
BsB4CDCLEdtfC1BEUotILzhPDPYMrJStcSCvs9TmqkbKssgiER1WxGDfgl+m/vff
AWXSGq3Lef4TpeFdY3Nv9V8RUSUeD/r3yKYZykzOV9kwqqqgJPs51Cirg8Yuk4UJ
EKUE64FSs0sex2nR5fdRkZ0i5ld+3Yi00Gp1U77rCTVb37qP5Qcs0wkR/APAKEmg
XNhZuQsLFBezaDXc2h67zNYI4j7t5svhhiVamms5R891W2a+WL1CIrvFkr8MIgwp
pxJpGnTmtC++8NhYfai97ImpVN6/EIhzMuZ2LLCnz0y1DDFqzr1Y6Wb+v9auAWHk
zyuZXR1r/S/kLFVD7tUllrbY38li7nvx0z7P/9xN4Za7CJaoS2/l/LknbuaSs2FP
LEeXjuoPINroyvMhJrQ3cslvstwFIJBBGqdtV9s+pMeG/2I98QTCOEaRfUCFSIrw
mDFW5K0Zpjf9zLHBFBQnMk1eMftvGooOZvMp38oDDJtWQjJnlBuOp6ZecpY3O9Nz
A/SLYWCwNGwabEx+9xmmjIf54OQYvLgGxxX0fV4hiZ/A6DWVUa2k7MU6C87LU//O
mY1buFMkOZ7RYSE7ueGngtgG3LuKKZwQB58uXpki1/UGWv8Qo2wKn3QHy8vZVZe4
jTvfnIytqmNKvHmI0LEy2Qzp1T0SHQaHKxbx4vx6A6fY7oyS9JoLF76RdFJR1cTx
rBMoLgoEd8Fdcigz2GQW5SYTERWe7kbT+Mj7Ai9kmwLM6go7E03o6xDRGGCJiaWS
ug61XGT2ybILrcCMnw4eDPlj05yAWl+BFLcd696WjoxKABYXOP7rgPKYD+lOYbOU
C5uPMU2lWCjHsdfxg7E7Hn2szO4aF1ws3lpZ+PEhMQTYTqUSZJ1Sgb9PYJXo0yxt
aJ8RvFs+h3oRNFaQOB8818jVY4c1o46SuWXzv0Fik8PB6fmPAMCg+bC8cxiXwWA9
dibiG3khhM6cjWQ03mH0ptiF0NQi11w06VotKpuWuhXjZbPlrTNVOeybcADf6tNT
jfhgIEij/UJJQgTZh7zoiRTBVcSE+z+vJ7NGlHEmhnhPGZYPew9LrY29livwItuV
LCQFh0zl8/osKWfi5FpSKJUblYomrEHTYyxnDjCoRF3SsuzKyjL6hwv2+HHXUdQM
BGrpAOgt+EcYIKHrdQ/2byyM+y45TVsfFoU8+tzAlijTmVp4X/PVnCQTmMc01xnu
1tKQR0nGdWgEcIvbvzBn1W1kqU5mdP9P3/Bwtc2zDl7WubwajslEArEgIrOVSFuV
lqh4CDs/AS9l5hWojQehigTjGJTteqxN1TO6PHUBl7tU19lw9RtYyHQNC6X+5a7Y
HUFNzqBZf2dl//uel1MM351UESdkREFoTC64Sj5NmCsLR7d+wvL3HQ3L0VGVhQxD
VDE5cpQUeNjJd/WLNz55cGfooYAZmtcVSDAcXc/EDZWHoDd+fBDolueVbfjw8EWf
z8An/V7ssxPTBRK1UGmuCrDOE2oj2JRDU4/uCBQoNZ7CM3C55yrLuOxqLBR5cymq
uWyRHup/36o4dNkMFIoqT/PJI6G7fiySnhqyV8Nd93J38zakKsU7XvE90mnkwVhN
yLx2IH74a0U1UFsdrHc8Ve+v04RmXWG+LvDB051T45KmrQB4C+fbL68P+n3i7yl9
YfwtI4iFhoupFQI7h2BKaUtf5KAkzLttWeY+ySUYxMFO7xSDUd3o8eSt+Eoy0XrW
IOc/N+WhbtZ/F/utvFQOmElvsfz1A0GBjwMqovsaMOzMjmUQRYxGUvcTltTZqv37
XrOXtf2iJfH84DvBKGKuO2E5C/FJYX/oD0CuIBifzZy6dWin6H18rM0TI/0qdnjr
OiciIFi8kYCLKJO8+SAPWnceWmzoI1kyWUWPjMtzfcZXV5/18uange7gKno93Xxz
bY6JJ4H7GtjNw3c9IIUfWn6a+vYNxBaWn9uj26UczFXMbHIlDCMgdi5cga6ybo+4
onr8fRxrtwNvxBEqsCdtoEPkNMtiQu614KMohvJ9Z6fMX1jnvoipFsYj0bkiOZDe
xddOK0vNVSo6Jc5vg1HtY4GX/qnVR3W+cMcmckhUqLV9Wv6NXBDgsgw9aGCRA6uz
Kz5l44sEYKqL3Zqta/95Up/9nb+SU2vUnjzVtIhVjhBgIj3qWImPwzQsn2XRqPrb
j0YompI1o+xfQhksgz/WkV39gq3ZIHbImesTCqyBAZz5pbo0zZG0jwkTuR7bJRdK
xEEWDhIN+69dEblEWbeoUvvlGIX5DZJK61NyBsiG+O8DVx3tnF9S9hVbuufghG0t
b0BiJ9cWCYnb7yg8KW/JHged3CiS1Zsxi0DxQO8G4XuVPHgH1GkgRYJH9jrstmqd
BmpyczxpRAlcCFLktajYN1TWmZMlBkraORMs0GkinCbuewmH/vij7nTLQ3FK/Bg6
MJC3oipyhP5UAZgTqhq3aPdSK1CYGrjXZOdFeMcLkSCQ6j5HreRrd1npW0cXyg/a
U3BAHXxrHEtU2HAf9H1xiV4dIRAdE7IlHrXvSUiuBRputpETZ3IC1swdzdhNEReJ
Imvhrz2bAAp67U6zxVVWhVwIIw0gtS5wSqOJ4p9y2NZr4LFCnv1M6V7cmmN9Kdsc
ENcVyleaieDPnGwA1cB2d8t6lixfxBNZEITW0gFQT1qlD5Ad/jtj7/301ktUl2Mx
GwevWlqX6ChkngojzuewSJ8Xb0xN5cJNCzddxwy+rdh/OPXECu1+K1sKMHQYQ9+n
F+4Ggif8/RLLwjTB7wlPFepUuBYNWAVM3rE8WrshziS3fEDxx4fvrjXZ1cS6/8ek
deMCW7FLtkyr6SaW2ESzsOkovqzsgsF4e4ghpUTgp4u6vLEqp2pJGfHstFoih0Ls
NRtVH02wZTjAHm3Mv7S9L3/r7VXC4jMkQiJDec1Lr3tF/2TXFZQcA66O/Cr216bn
kLSScP0QlC2qYZJnzFDVHoQuEeAKnPuxPOr44zYWKqJqnB32tleNsCNPqpLtvwTA
XAHzyv7tgucBIZ0G00I1nqJ5YCQrkCQwQwp9YQvXtqr8XY/gGWYTrvOvcsOqQ94+
K9/jpfRk15g1bzkR/Hp1syHQT67yZaiPDY/XBzcJkL9c1Km3gIcalWIbzjHleEMO
kgyhHzzC7O6shJhBhdMwKlswB/BK23f95+U5UggpkMSrioUvNi6Kzs6Jfw50aS+g
D3kTfGSKoKu3RZUUyPppRn717p5+rgxcC0kMhi0n+E2wEHUkH5gChxUdghMqwiyA
04tKKUyqWD8iwwB/etQkjkkt6p/UPxaLkcTLIE7ggI2oFgGxM5sK++XKlD0twHxx
7nzGL1eI5YWH9PRJyIkN5MxYFp9mdaKB2Qw0qbUO5FtnmsjWm3xDwrBnns1kRqmc
qTyi6/OeNTr64eQKdscTWA9VvHq6yqu8Q9uPKqKNtaHUN0SK30HqH4WhuHnKkg5l
AwDIZNgsxpC17VnuAtvMU/GbIraIGlJHbZ3eQkVg6jevbjDoqDJfO66EW8rGlXho
mUfUEFjlQKRtF6UFy/Zxoa/c/S3NB5HCFUY2q+754CGQpR4BdvBTIMIKIK/2h6Xm
MFgEdZPmZVAeJCZHhtTxDi8C9LQ5htg82HF4kO3FThiTPsH9n9YCGuD1tOSEDUwY
DhlLFXJ6MdqdS5CtcW28v4bRyZ9FcT7OApVf6HnoRUX25OEi6Ki2SpJbC9HcIDt+
5kzo2fzd2Sibqs/ST16KRordIPPLmNKI0ORVMowoWyvp109NYLH8oJPZFHYEoQ1c
OypyErBDQgfFIcODFy+Bx6tVBp9uOrIe3IZOmcFG/PfUUbblCPKfyI+9dWSc4NgY
PfCNwav2am0Po2xAbpZDNc02qyGDuu9OvOvFdRZwdJgM40meL74cQlV0Ym9BXPTU
vQCCmUlRbUBIGm+f/L7hQjW/go9vZgp/6vvIBQAUgfQmlxjee+jT+Pol8GH3AEpj
PVjrKHUSVHbEqaeYVc1X0R0R7yC3/0NOMMZSQRG95g6rdx0PYySg9o3OSh4N7DSS
5X4XNsMrGK5qOyw4QAaVOBxLny/uGdutVG6u3em8KT/Qr1MowJyPpzOAMEsVRKVm
UbsJvx/5aZwvJfqHYmLJKx987gKKQfRJRtovpm52xpIFC+3Mh2i71KTZgpjAUDk/
SSK/USjfxeTHNMH37nQ0jP5o0S75UwQpj5QqQ1ftjDqr5y4b/Y/ES6WpHeBrjf/x
2SWVPs43X0qVG36JvuocmQYivuwnWCOrdI63oleQu9BzI2aYUbrtyIufhv/xnimn
45JOsNo9+mQtp6x/9ofIZ5H7u5I9BDiwlY5AM3WzgLvm7yfX+SB7NKuy1nCRDigP
72TvdGuoEDo8iEnV1CkAE2LUGwYyfYH15+OP9IkL9HFWHKg9qmU52JkK84U/kxkb
EZ9o9irGcwlwYkk34rxrR3VrRpqQrJpD1er54S3C1r+kvQP+byny1tbgVyYQe1Qq
IvSFSg9xOq8NuPQGRFIrnPFWZw5fwOhLr2aKV1DpUkpJSx9nChOuYzLlmAZnKvQx
S5UTjZvE45isKXS6AyEc+vP4xdq3M2IkeGBJrUfcW2pZh+JHHj4Aa+67o8tkQ08R
FR/B0rijSqvF13kbh5yj/12cB0IMnU7p2llGEVxWpwCouQtMvSFLzgawhrio+gks
f07Am4sMx4Jx6f8XzfFZKpd9f2shL0SJkqefnpls3a6cdamfOVLnrvNkGP3KiTab
4HVhW1BC2evIToODO98KlZzarvHbgsTSL5UlVyoe3FNCcl/89i4M88eYhGVTblh9
pAuT2TTSKgz3lg+OwoOtf+S7X1MZXuZtU5Jz1pFhWwSi3Acbw8yN0YpUytHHVyTu
NMxm9b1xVIzSvMP6/XmG1ZpNgTkCiMlLLLL6tZ82P2svN/MxLl5qC4IjpQHsajuF
119QUIrCNHCNdSyBrhLfD/J57zUu3pjnnWQc1qsEFPWZP4iLnQohfJiorpySefi0
fK2nxvKfOxWu48hzlg+eJM+seIWJZEOn9DFKAi6Lp0vGs5DtuJygubVd9ahQjmXq
hmaX+GQY6gX77kITefNyY5801M9q3quT72DY32+EVymBYWTlhUn11iLLrM2SkudZ
48R33TLs57c7Zgf425fhq+f8uaIZe9sSAxPEXHeuHoOteXIRVyuROKOalY3zoDFO
85uxuWmgXaTHCV6pB/M4We8l2SHy6ZsnM0gYG+tPPRiB+K7XRBTipp4QpdduniPg
Vs1EYrH5JtoeRig40fsHyc4ylOHtxIj1wYdaOtRvFojDxprhFA9V30hOCjbWa757
rtB+smkrQter+2SXERbAqCkbLxa7uobhAv6rZo3sgXmRKcCC3sVnxqNye02OZeGl
CzbrfLDezgV7a8Atx5jmMHvkUvu0TAEEuDRWB+AjD3cEuKTUGz3hcKb4MJhQ9xXO
jaIU3s+YMK10MhwpO6Qat3FlS1qGO9CfHGwq6StVYYb9gB1+tWZuGMb8RI4vxAM+
xaNj/Kno9iaauNnTVn8tOX47rZkKKQt7BwzvgYy0z62a3I3dSSFviYA1T2gLGrp6
ffyhYKz8yx/oo8XZV9ULmT81ULCZKr/Xr01uyVl3LD47XQnBS89gKWJfptVrW/E9
0Zh9z1/nUriAa+Aqpzts7IA1UDjM9ifQWb0yBxtLDVPwcmEB1WSKwkNxPV7j3ZYL
ecIKLrO5zsrsmplL5GU/7ECHqzSZfcMigKcagxbMfut/TPzUTD/rqdoaE++dRy8d
Ypu77+zYaukOXrqxuGMhNBvVkKn1+7Gc+SNdxSRUw5rU3SZ4aMhTwh0gMlumvrWa
1NtSVWyaL5zkV3FHO6GsZVacmSV3rd+VzoW1rb+8oPTRB4yAt0NHv7WBACDD0oE7
uZF/o47YcXrpALqZgArPUzsP8iSDz74Y+C65NXLdQKJdbJ8u24weZL/IZNiAJXd4
o4GIozl11fWko0tYl4zV4kJuP6EGZZnsWMOK19j9/Ayi0QimL0Jd7gQSLR4mUx70
Hx6RRtBpVr/keopgDfTzzUIl8NOoqcGPHN0dDp5bGpSCqWisPX9z6SnWyA1f/LzR
HAcxdDMKEMq950LOKCr+WEO6ucOVL7w3A/vLr2Jg0HTubNbZHURcjB2mbrRE71E2
xAVuDNboIUZ7FcTXBRMc6/YOg8M0l9NG2kkwTfGRGkaghKdaVLDeHgdLageFKHUt
Y2i541oj8PdqBe9AjObyrybQYbnWIYi9p1t927KJ6P4xD0bI4RqLYeZmkFVTFM/9
RfoqUvEUOTf+CyM3u+1mUdq/FD7rhq48eGYa0BTelyCE1TzrGsqYUgHz+eYypiov
5CXPwxMhPCXxsecOauohQECGEbQIy45x3DCSubAqIiV3Y4OU4RqF3QTeVB8bdew+
FxGy4yuDcfI1vdNMvQlUWe3bS8ybl5co2Ejr4muGVE4VTHQ0LHqo+kSd7b7h359B
LPK/CDvbu5QBoWR633WLOdwWeOEVS72pt2gLxp0npoj73wEpUFYC19+FwujauhiB
D+Z1hiboSNNiu3q81Rlq/ywHJbB8D/KaJIRsfWAatbo34AtSHJX37xkpSCUAH5wK
PXd5OttZNsad4Sq/poO+TVYCnzXZrR0Rz4A0FipmGpDBmVuEJKWWBpTPmfBvaU4S
cHQ3HWD9Svo4EFPzsE1e5kh+c/ujB26Eaq+WWaJwI21Bzrdz7fQ22dtp9DBMnxCQ
t3PtAr4K3+ebEPhaTMGCC728JH0goUC8NJCTW0gCEbyQA15xcwPrrUhDxpHAmr9M
1bbOGPd5UUugLf1EakjuP4Vg2IGg8YzjbBrzrnDCbb4HkdsWWFjSQ+tJ6J5W/wNX
USmL3cFaLhCmubRmg6JL2b7tIH3Cwd/DEcOvH66WEH9sFNuBg9/g8d/f/CMPbLFH
YZSVTOL5d57dsi/6md33XTfXIelBB5XRfc6xc5kHRXd0me8ocAsc3YWzeL0PYnP7
XhYcBQhcBcBt65Syj5YFF5XCG3E8RNowYL58W6kfvfnP5tcFm1l3oKrctb5dF7aV
I5Uoyrl1v/wtLdpy+2RlE4Kgp0fgyYTN7znE3kx+acZWVdDeX2wrcPkYUg6Ecw2g
FpqlMWdR0XrOYFj9T9fkaE7TVBRfdoYqvOUO6LL/OVR2JWMjN8eIKcCTDmptGHjK
5BNYehk2Nv1nJOYGDflx5rsKExQT3Ws2q3cAyj8oHiTcUdzlgTDFBOR+fyyUEp4C
WG0gfM0XTLOQ9x3bLLqBxJYfZOjCJM3NBbIKedjtj9fVKmYiqEeCDrox28dThlUS
sJwMEw69wc9QKH7p6SE4O07OyRdvIPGMp1znh9DRRllR5yxILb7IapxwY2gpxA+2
e1ptBqbYrx2ZAwbQc78scfrMYld7Xmp/pypmjbzLwtMYSOsx3Q7QXfVa4rtt77Vt
cwEVqxZxEt1eQUQqcuu2bNt6vVWBaXUm9eou7l2AqBuWRg8Ypo+i5+r+yjVyJjEO
KR8SYHwF+zdNAcYgbbMUEA4NLZVGXAJoKBt7x/PE0qCjIHGmZFB/Zoz06Ki1xip+
2H2t4kLXZlKbKmrvs16jiFNtfhS1sQpkHunA7p9/6ihs7MQQJWE7uwSdFueckj43
JcIs9kysRzeezxCAwySfinnJ606bC+FNYb7zVjzfj6W2T6RzajtedxtklLABSYKz
4RUYlgoTjHtSzDo4YU8K5ZcF0bH3RelzpWw3my7+lx0GB0v6UoIUA8a8XtS4A5Vf
TUsXLpGGOjtz2Zc5kVoTTKEGKdVq8thSk8ERP3s2bjlXsV0dAKh+gwuUKhTEVbfp
ESAMGuqeKIodwGu5JR7FkYFnSnsTnBDlE90NEQhaoLJwIBDaAbQyNwiBfSqDn/Rv
TqBQ0HVZILjB1qShS0OOeCTOcnVWRrUNu+Btg0fLF/K/PGlSP+L7KJfjRHqwIWkt
FPToFH36IV+x4SbwYpiTKMA3HQghhs4NxvhlD4UWEANnJ9qw63Vipli6mJtcf4wh
sDmxXiTdOy/ktLM0R4bsN77a32vJLZorRavukjd2uFclu0hDfERYmYhN/QzgjAcZ
03mHXCG+N6rLN4lQo/hDu2/wD7fGTYXMKLB7Ma35Dk0RhPFCwV397SltQ5U2iwHY
enGp5xyvitOp9rN6c/onusXmxkuu5So//Ag2pM4Iw5UxgZ7a+8ZccIt7JTvj7yKl
h8q5OV1ZGqNzhW+84IaOAJD4lF5LzoYRfqE1a4y1zrMeeSauc1cPKDhePFGdzEzj
epkgKHYXUg/H2hBeufpOr0uarqOBMi0RAMBkDZxn+opoalWOw6VIc+IECLMBKPLJ
qUCma73/mwpQDreR3NyfCeiVg+3GYDMlexscTuLY8gmq8/ZTK32b8kH+F4OuVXvn
Y2uIdjsoIL2sv7Z8Oq5PAz7MuPbRfJIlaXWWTqHBE01htnOb4FA42jn6N8ZylGlj
CYWQyiYWxHae/+dhmJLGtGyBXNBhnt5HoApa81qzk1Swt+fUBFxbPksz4vcO4jY8
hvEnvWF0iN13GHC7Wdv4IWUJqXSuRIkdI5YrfbpyizQrAMvMJRNzE87zuQbSZaPv
Obd6qV0OA+X1ha81x4JoHmK4HIB0Y3T1157Ng+OIaVraxVP/8lUn56y1MxgO94dA
CzOj9th4TBLyy9mPUtp2W38H8JkgNj2hNv398ZGM8zUhKbSHD/hfaJWdiaO7RfOA
uxyDFu/MDkfnpzEJj8LQ28Css8uRvIViRZ8Pl7wgE8Roip37MmJ+XfnlYkXEWOtX
kXswx4SubGEhAB09w++hLyWGPuVVDjt25qxiQ0kWbY6wlTCgHfuOb4UVqeGjZhz9
UrF71I6q/CvpTh0DuiUAbtJ5Maa8+YMSjKhNg84/mhL1p2aPbKTH61V/n7aRzPfT
fsl0k36ZMP+NM1WgqCzAsh40hBmqTnLZOVy/56yYke731qTyo3uwO7z1Mbb3ilY7
1KbZOk5k3S9XAAaTTvG1vCeU2kcfPw/TklXzZ+KNxclrk7QCMc4ENLkiztHZ0h+R
+d1suIonYHpNbSazBW85gQE6kgkDBQihn3K+xeGfVVpOPd2qdaBxNLsek4BpYi0N
69mlSuoHAEaW5WCZbHqhSX1+41BD689jqjquneiXkHskaa6bcKn/kcQi8+J6AYF5
mGtAnNg3UJvHtUflJy8BVPlj6rDKh12Xn8hzkNHey2G2qZ/aqu5ypjGsfW766Dkx
/b5t88a3IjwuR7JI1EUbZ/mrDfQz7tVgL8snarIu5dnYXgJqtjUkTnZ/Lqgwcq4p
l/YQ0Sciyv1G5nnpamrM4a/XWDY5VWPwlfuYjahm9YjC2JPrsW6aYZqiEPaxRECW
MmG2EDSYUTYDOVK+P9FvQkUryBYoxvNGZ8z+HsW+0Zf6dyuLpwzNHH9WOOPl2d0V
FbRwkAuuM01GLZstVGgDancYflnQ1tWb0frXkdKTzwgfid+vtynkwDzcAVLd2bew
j4FQMN8ffXYtlg5O4i/gNWAaUQNpHJ/Omvyku3IXk9qKFcJwrZN0DfXfH+Cz0WoN
o7J0TSKBTeJTZYeFeFU/SQiX5G7y9XCwaXUxTeDqKdvCEk33fi/3jMSqJ8uNe7gi
itYrCfCIZrDiMCveWm+xpxyeAQRMbB8c3aJEsy9mUi3HJNNQnNDjZKlcDaRFn3Bu
3MSY999PDTJk6VSN/jNcDR95ZNP8KvEtRXfH98AkMLK5/aEWLOiAtch3VuXWxBot
j5GJp06j3aFqioV7vDXJUkPQ2qsmB9xUlPyUHEMNCPgqlZpcfSQIlTQa6ri/BYQF
nv3/vAaDEQFvuW9vePVzvcPiT+9RpDY0gv4uXQnqdC+ETNFJ2/mQ7irrxRIOIQ4Q
tQV65U8trj8ff42GNwpKUtniDkKFpA69PZ+X01N2s05G33a8IRRR//ALHBLhjQ85
o63QTTcktfZJarWwCMy2egZSFTDGgUpO1CI53sz0VVCsqzh62qqnuDDJ3tVqBcPP
7mdX3xZ9v0oDQXMx6ORvw4Id6tRHOZVrD6224HpjoK9cParvSkKifbkJAHpwunb8
gZycC8+fPHd+AY236mfMcf8FSX4CFt6v1ZMnvvNEn6uYGByzW+MXFS81LQsF9RT0
5cDRQiZZLPbyiMP+cpxIg2fblp+YltBudySrTGe4tH7b3vZOw716jPGXUbjehVE1
I9KBd8ftkMoMtxiQi2JGt30hxip4fD332I3UABuIkiudrc7ahq96V1yQuD9dVvrJ
VEpiI3O5JBOI+c5Z19sh+tAImBu+Sjqx1PojQ39KyD7SXeIiqUP3Aj3uvZja/QH5
AQ8MxDabnzsLX+bMH/8Bqdp/xuU9M2IWSi7YFktlWmrhPEzB/1iW0hiCoLZOX+Pt
loe8PcAyJJ57mOCH5PlwtkzRYsv/R9BHxp2ldlR8vN02saqv9gwlIaMqFHe3+3c/
8WEw87aGVCcyiFQUjxbc2zGD9fwvvdMaBIzlFeroFdQHGtADib0Ndrzd8acInspR
OYq8A2BZUa/cFO97HeErK+a1zNQsz9W3w/NsPbECYAkg7AQJVCC13xUYbWHyjd0l
RJD4D7zndv+jFT7kSl1yeGqg07rPgg9awnGDckikOIqhLrQXj0E/xJiP0Vy2iKYD
o03O+xU3ap68uneSpJsb/fs4vMqhChov4VTHJtMpIAGq0Tc7lQS9155WbS12T/vv
bMxTcQBK0W5SDXrslWywdW9pw2bk5qklQtA8o8N/hhHz1+Fs4e6xk1UVehqDg9pM
WYP+knPA1aVVMr4R8n0E7gG3UPb8rLn9SwHq5oJeUJeS+sQLsnouJazwcBwHW9m6
W5WI3ir7QtnllVVlacFNV1uHuWrkDmqSwBkqBt+QrhZpQxswpdI6Ky6voD0K6fGE
P5HcWB6bAA96jEogLyASWNkFYW63jc4vZNlvDHDSXlDvaLJRiYB0u/0xDaQVUYeC
rHeSdIOD/JpFEtbSgrauGpc8QJcJ3rLVgq+ctgND7uSncLB7RtZjsL4/G7X527dq
bblpQP77NzctSeQTkbJa5deWaros4GsGW51k9GhYp2C6ncTqTlIoRNIv5mUR5cH/
Yf4k/5nsto0chF91NiGgzFV1Ow55w/yb9Lz9OBpMdqdnFgwhG4dBR2z8gGAeAmzn
kiZtYve88x5xLmfM0g5TMxlTn/HrT0RqeXWBK4Qy7Hh6I9AOzWad8y3mj0lovuBM
GvxxzLLyqsFGfAECDv4sobBmsYeN4iRLz8gk+pDUqjLGr7DBPhhkHAVgN7bIQCvM
PzWdIhiHkx6QrlSQLX5bQU+xX+2xCE4I+6mW35vCaknDcLFaAoTeNeIPu5RWVc46
4YTY2Cr312HYnKIriY/ulmVoCAgkdgKFDT+VEoDRUsTfyfJxNNrIXfldQMR4OgvQ
2LrJ81e8LB6twQJ78but4zwvVi2StRpfkpijZx23+SHqKcunW+zlJi5nFpKkOwq4
eMSdMb5bFDJ5dkiPZauUd+ruT5GCjtAztIsMfkrWi4+Izjwzh7Tw0IY3DLw90pOL
y/Nb2r8H0kSiterUDbWIffIYt7ABprHJNE4g+UpkIzmn+k5F/2+rB9Tw7oFQxxxO
NUeFQWDKnHMF2RGacHjYeoYFl+JntpBCGTtPOxIOvFxrYZ64T2/dTWA68xHAlMsO
Obaa0eCc+OpKKWFXR1Q4xoNyHPXasxLDAkOWdCAeSboJyha8MmmpUqy/VsTDav7N
2GQrf2mPa91GyxlUF9bMIFFNm62GyPuJinSJbe0QCLVPk+3fG6YUghiP1K+zVCeg
3o8uDyBwtIio1pnfZlzp0D7BSR2mrJNk8ULLjy8T4gIbQJdXQfW+eNL+WH/hJeni
8FGJsb+tQNgVhrj/XXOcwIbh2othtVuCB3mzt9ZP5cE6zt18cfA3M5WAjGCJm0m3
6t952QoMLnqiruXDixDPLUuWguteK64Mxj8HctjB1rn8dY76m1vIijStkz6cM7NY
EULyxj4DKA3otWC3TL8Emg2Guh60AnN7jx1NrQnh/+TAJKOfLctOscyZnnmX55cW
ImuoR6FjTLxQV4ld09kQZRS8XKUjthg4KFDjmMcOOA7CgNxjBZ4bT012iRZg+BJN
2+kaJgASczjpi1+yb1SgH80ujG1y0+3t6znujoDAdW7Eywp+yuJpf9dtEjgYgPih
4PQ+a8yrQdYwbxKC7gMza+vNYFK0/V0I0knt0qLtp5RHgSlZ27s5i0FRVM7rjqtl
mo5zMnEvrtCRiJ9wsg/MEtdIZDAlA8E3NRGhDXDAVRnE/bY4Q16rLemPx+xgr8IQ
GIREWfFiAazVgEeTMRIWtlHLZ7zQYEWOUrKjzMZMw2SEdUsIW1BBELJdlTPFe4Y/
yXjSDiB+h0ESdVCFJJ4y5YkPbOSqyBLtQCYxoAkFDqTrcK8YiY6B+OctEgHD7eeL
3y8p/vgjAhICeILBwYvmH84tEJnOL/UxNfHRF7c3Hae9T7KQ9xKVhReKyyfIbZTD
MF3RRAn5L6UUXk4O8g+t7J++tdxeapimHQR04c2vQMpRr6toKi9Uukzi1I7wTtei
eJzDVCquFrbsFycqQEN7jm5ZE5ycdcdjqOren3CbEArjRloebmqzt0RmhnJrvL2X
VuZRtf7a9fa1VTLgSxvET6vgeYN314rRmKF4QDYA4bqzx0+dpTE7dxWg5mlKKjqz
6LYJzkc3OakkIEqQTFLHtN0WzrM9PNtaM48VeQ94V+rDlrrR1dnT2po/zY8VPhMl
i/xghuRV7Hcv+Fr6symaCGNEF4jSKL97uXSHqEiBiHJtod6TfVjnt8nvXCN9CT5Q
xJwwrEbMlniMijzfTC3fJPSbXN8xOi1FGoprVwmJwJQwkwkuy03tOMVfn383K7vj
v6RnNAmE11XXZDAu5EPQWZKlgkv+KDoNv4F8aqZfLPMVelkmbeuJhGdcGRXEacOu
n1kCNy8cpueeGkyF0h/FZ8bKC3pr9BUjgCFsTNoOACjDhjXLZhBq2vooYg7rPnYi
1sf+heZLWgr4gpOYYR3rbpZomXBW+Rg3x8wIBvtDz4KgirYLgsyQ7cIQrNWsY8fi
0We0KIHGBeH94+OGzTNtcqqYzanQOBBZFrJrFDM6ocdRbTllrdiB4cGLum/wTDC8
FH/ggl0qCid+Ioj/Us1RO4pW0LPGOLVz8dFTpD0cNa2Qnr38z5wGoZwxgt71eo3X
aFhYoPHp06aVdNps4oVT2+rNm1jAN+RNCnFvxKtk4czy5GDphcoq0SxHTlKogafK
H7zxDff1qplVdnCTmAb/D5Xg/KSMn9UKOr/wq3/spw28QPyZe4dohDJQOFWpm0fQ
34wkXwOiKZlrJP54g2tzxgMfxXw3CT8NMf+qineAiyIFEmvI4dWbQgBcuUYyDk2A
z6dw6WzPF1EKr7u96mSb7ensvvAw7nwZCKwTlH7YpL9jgOFjx0HpdbkcRgPJKahf
LVbZYyg9c0XBMyVkeaEUfSgkj04EsutbkZw1PP6dLGDIF9jY4v5WJTS1HD5j1LlV
asTKBdbL0Da2pYJq5BZt+I7S7U1H4K72AJ1mXoQ+9fAl6UT4+t2cpp5tPPZ0ASk5
/cPMMCtmymBcFmJAev0j7UMuXarGgsolf8JIdjADaWhO+L0nB0pLQ8EW0M4kYKs7
4qrE9vgykOVHWQZ2eST4/AEQINHhlRDwF2glr8NwYIYm4Y9i81Zu8diSlYsJ+em4
+MyIPgvfA0ZCz11UgT5Ytlr0zv9S/WOuDMs94kU9qov3r3f+KnM3vFLOdA2UI0Ld
+2dRQTEf5LRC/F3bIM6TaNz9+T61uzM8w+lKP7DgRKGgycpVZ67mYc+iuJQQ/PWq
xiFOcEpfVPkuADlfH2XEIfE4zm2oL4ymHZU4lLazP7hDrYqPPqjtKtCDaNTg2AT9
uvrl4IZ41+q9g7rCEVF4eMoNex2KJ+gE+vZaRVQEepiGM6M+eDTLW3Bn1Q8GOe9D
cYIju+QMpFDL62sSGUsKOcNOlj4n6W44P9B5V3y07j07uS5XhzdXTWM4EGE7xzeQ
J/T2IduHX+bt7Jffrvnl2Rt37AZU8NhnhWpnsIks9VBxO/HgTeBbHmiPESov1nVz
H7ITmSgJxYOq3Iwx1uj5N9VtKQXCLwN4rXRvve0YlLgZB/PyJtMvfUhVDfpAdvCt
PMkCI12vL7qB3HyAJtCt1Fqlm36jvxPgxn24/8TbAIdgvDiKfHd3gpwqgL+QmAFz
VXNkdKW+expFZcuCpz5kSQ2yG9HFCyVGLEqQyfVPEwdt3cy/IdoeC/dWPMV5vHsc
d70s/QlaRJ1uZaTjuFhrWfh7TObdEm3GnAInrL1iUB8AWGjhb8AEb5ah7SXYgNbK
JbQadjtRNI1a/mTIS9oQSZCdmxfKDJWq+b1yBVIcnva4neddGBMUAG80jmD94OSk
vJM7TSN6uHW79tdRKaNmcBRj40+XrG6VIvv5LuxNrGj73+Up30+rcTWrjZ97WGyX
sRqmX7PXZzVMTnGHxW5/OOfLpmaEbM3fZPv7h+Nb1Q/PE59BDPy/Gz8YxZcFi6CS
Nku/Eub9tny59db8L3EXmexgjbEGrrHTGa1OkxNTDI0ATgVM8hW9DM9ICEY7abiE
ro4Nq/Z48hgYBAv0UtAyuyYv8ybBZdN8+dU6ouX1Ddn1/sUUY0uaIhA6ze/HagE8
NriC0i/cgOF6q4UbO0jwI0ZFV0HAjDnlOfP9HeaKYAUi+Yhoa3iAqfwsLsgR+Bku
95KgIG6gQbgH/WiATZrmviEhxDF5IuzZ7UFdjLHP46g4TOT3GYFXZRK4ZDzlceGV
tzV7Z1XvDJLxtp6cZ2BWrPXEMiMO5DL9V0qvetimKJmOcu7bsm5xT6ha7j4ZiVVw
wvel0K1FBO9SK5tli+Pl7AGvF1oMxpVDGQpbx5MpkiMgCGVBu3lsF0tGY1tm4Tzu
yTOAzZ14C4kS0YE2m/9YL/xZa5Y/byyvN/FyhDmSHaEDeC79z1GaMJncanFZsVBu
v7/W082AyGBXWZMIpcDU+A1NuIIwous6A0hdTYPV9znsBJGfbOcOMRCPdW2MGfII
mSYRA5nm/w1o2vfDYWqTguzlP9SdN1nb09+BfX2KQrUtKbZl3KwQXq/k9PzcLMkV
B/U0TUVlheC0DFU+oz8g86f5QHRHHx5M5+lzwOskbIzNiHsQy4y8Bg39jnsFFAiS
JHw0R1Mw5mtKALjYjIXKuq29/Z+dK9j6FinNF2Z2FHLPnSUr/beGVVMhmvqFUn10
xXt9k1YcCQESlQ1Vu7JQAex5KjYe2LQNp4H7deo0U/Xn/YoCQOc6OG2xWlc/L4Y9
3gvq5hoS1Ld7XM4K3U5XE74wcLXjnA5NjHVW+i+NamPMjdRtDDKz9Qk4PWVgM3HL
r/cJwyvrICfGWcer6EQUS2jO9G3ZRC6b1XHMKrgcCwJ+lt0P+Zom6wL0Cik6S4Dm
rWn/TkTmn9CRg1sT7XZIQdqJ1NLzw+fil98ukC0vmlSvQMkXViCbiZJFZoO3MxOT
OJoru5vNyR81mUNqeORa9z4/oXKTdRkCBH7TY2F7MXRtPpI7CXSgxMpJv+0adYDy
FwKgsgadXUVpXW7011WhLggDpzUF5Ohr0wuGl2HISdAUkD+J1/nvnV6/vsgr1opW
B5W89NhWIcMeltErjlfbVEcRt+0HN1RcQsLlCA5w7pnBNzUz3/9hopjlP232BJr6
6Atm9m9Wr8JCvM+YCfT7f0b5/YhgIu5f4Jy1HVqcDSHdT2zAaG7EbAsSn7gLYgOc
ZTDG1paqhBGtDlcSe2kI04BpI3AvsQA90gbDOVFqkPYGQJS35zGHLNuVF4wCrmpU
+fx9x5Uwv/oFmycWQihicU+zDQkn1Q0RtupzIzPaBwTxmnvzMJcgupmHnB9I/3+h
x4jVHVbdb14ITM/YPMIhujMMjVOXvXYoL8H8dkMU2OQjYXsq2sJXf/jfs+OjPeR6
fU2GdxH3Rx7RNIzgaSDccbvj1og5STSTioPDvk77VctuMBOz30q3zQmUMGlK+4mU
Q32ttUjoSP1o2oZi6nB4G4bN8Fzq4E6KeFGnjpQ34LoKNW1U9gU3FNzAe6sIXUpG
BL2980X8hfTXVh/nqqeerv2HXRqs6PMPQlkeyQrcEAn47HDrpltyOv5A94ryIAF6
K5oEKC71kU/JkHLS4M3RU+6/GTKWDun8/cBncrWGpOSVNk8G4wMPKJ6jWFwYg9/7
RcmkC2JFMra/HD504vhGuG6sL1DTTmcKeLSZncTVl9xFElS2Al8y7rULg2fBZsog
iqdVPR2J5voDcGCfrPy0r56WiT74RGCeuUwmm5XgJ13EeT8Zexf9+ysLqm3aqH3d
zwWvk4DiOBDRFCP+I727z2mvUWiDLhDwpSRcpjkCrOErsHBnPkUbTZK4txYvS3vY
zlwcUTR5VWy6rkrnlPs7HQvVHCnItE5nhFhlm+kHY8bk3SUgJwm7CbWsHwA6X6Cz
gCbsJ7+5OYfXOUSv2Bn1/Qepw6OCokKLUV4noAEbuI+fFCNjJtiFFVPcPGCnsIF/
MjBUSL43co5dmKIWeI4OUFXpYUu8dKRwquuwG9dUPam+yboqyYZxs/tDeZTxJydy
S52ZhFWp+o+E1/xCoQgR0P1gwmc56jj+OD+SX4gbDv6Y7YQaivy1nyrqAGDhkHVa
8qi3ytFqmSojUN67zViCuh+lcNP/Nj7bsGZxLmISb1Rfewut0VfJfah6nyQt8fsK
drGfn/bQ0U0tRhyYE2mrYHkbCSbG0SYdqb1vdpJkocfDTXvcFMp5xq+0SoCJ7kZg
AKrozKKi4ICfTk97x0w2IfymmcmW22y4hrClK8TZoJMUo7vifaVvxMgLAfPBlAZo
I0QsOyf4HF2VN1S72/lBgYTcR/nSlNhkWVwOwCp+RZm2zPfn4/gXZinmpJNtbPx/
+Ei46BiDP4rRhRuXpZPbm1AaVnPoRkThCgRq3YcMEFttx7mmrjvbz5iBT8JLsucK
0XwUQnst7ThBDrbOTdoZSlNcpHeobkOcx3+La09HoMRDTKQr6K/alJ98Vi5gnEV/
FwjMkLaCNWMLdnr/6RYAxs5hX3nrlcvvv4bTUkz6h8+MWQV+Zyg3bxc2iqnSD2LX
FR3nX7/NzgFYIYE/oLdmjVYCH9VvNpPduwy2Ah3y/Pj2keXsXSuWaiL4Y8gkhvR2
lZG+imoSHKUqOt88qa6y64dfQm8uOdxYxa6TBq9Kgc4GOBsJrCuNHLOWb8/+CWZX
KZSsFNJavpD4tTDCQEESvMVfRDqjWX0zJbhHtwbahJJTdmGas1rNQG2T4qjV2mgH
nFxpO39459wSYgIHpj2D9mgplePQS+e4d/1vFamX+iaX2k1/1AiCoFt47jQQGAIL
eXpdQYqW9MlBaMLahJhaItGFQZmqJMGay8lB8v56l9UQDLF6tdlaialr28IPyajl
Z0EPy6huoWXBA9TkPHA2Ch3GoDbjuo1xKyiL9hHXRtoc25uu0fxNFz6Ur5X6Qe6x
JfY4950GRLAaeURh24dilEwoNH+xI8+gN06Xyg1kpdb+P+CzxN8uQenhhq7EoUHW
AFeA5eRhTja+JK5P4L7CrtjtxWPaS0GNslmg7l24x9RPyZClSPobLY/Q5SiAQ9eA
x0qa0ToEDJWhiETQiltZIuUzir9egK8IIzR0LwS6r+EuDttalNlGxJSzal5tFm7k
nIhYdpPuDb/9/vEI7CxnmppO5WsvW4wsPl2H3ubdBz2y6Ja0VlmGOv23tnXN6qH4
snAPhSuHByAlyXXFQiNINsfLq0VKsvLvojKVrfV34npbEx3vg8wATGRgQJfPgh0I
7DOYapOTXJO+UNSeY4nw417vwPEvBHILgPX/5jz0mJDA01Q+nndtZ8e84pgDigYv
TIADoPTt86Ope2U77OrngpdJYJGSfTVDBKhxU5QjoI568pZo61HuL2xLhE2W4h7S
NwWumomBqrfCD4vOfSJ0cvDTnn/8sk5otfY1yiRUmdPYfjiAoU886L6XpGJ7hkr9
o6zHhbVajx2pvkAFcVmGaK8OYrVfc8J+D1rELGZPgO+aiCmVBiFOqfsuSgq7bG87
Y0u5sz5j+mWEVDpLtXzP1IgBoEMIj7SCq0GbAVibSNFy69tKvv6bCYdyi5ybse+w
Vl8OGccO8Ig7ND9bHs4HrbOc6sorrTvBjGjzqcAJv5SlzBYOAmuRzJB7DV8aHITf
NiBF55n4uAcKGdRiQOUZ+GJF0sto/4TxLOG1gWpOP4aWBIjqYQcP4b+x5dpqmIgV
+JyH3xp2e2HDF3bJ1bq51KBC/6Aim6K/6eB3vBtNOGUguoQiO1IiUZl/F4r/r7ek
9+5FoiMdYLSxqznyIPifknc3s6842+BNKdfjrJak/HOX8JyMMoq7L4irQ/1ODKLs
HOtvk3fM+Q+NThzqd87oRe9ryCTVO0bxa3ood1IT/rZky55xnY436w9gEZgWb5x9
/pZEXHziyN3AOwXDdoYttk0gcRFnVkZzLNllEdltJYJOw8xJt6Ekyx2ySda+2vgt
lZIZR0x++cu6e3X6ewafbhHBgPQkR3zo4NC9PTyuZiNEH2EnjOdR6DbaP3zaEcJa
3Fgov6CHuOEG8ziFUNg2NlsTjtHGnbF3S1ybyJOm1FxESx8egp17EsVnyboDaNHA
QCvi7pW6x20EtJ1XvhxzTqqTsPoQvCWaJgNMwp8T62WQ2Kqqr1CsIbJ2dsbwV66+
H6O4E8XYCeokBRH2UvDA8RPU6HttG8GnrU32K/OkwK6oH6xcCWayR0aAyaZec0pO
VI621D23B877ySJEa0dWt2wcAe/HUEj0M6PjQfhDAYfjrjnygK56dhdvmfvdGjOn
1POQ7COCWMD5PJCJOLM4WJeLOzIs6+W9GNCe22nk7/kYrtnex2zuggTTpDqS74g4
uleoZnRNzZajlPaLVrOsIcF95czGBQcRk0aY0X3/uDMDyuVQxXEKESV/NkDLi2nz
eTV9sJ5gk29vZcvgYBTpixLr9cYlQs12n62bI3Tl1W5+bB4Ye4CIREiRX2ExxjB2
ljtnGTDs/PeY/J1ClzB2RHeveez1tbrzqOqXileFgf2az6ChrNQG4cnmdvTaKOGr
IaTRVzlHahZyLVocy6ZFjAN6L80EGw2UoBnKRgZ7Mkg5j4NUyerf7i28iE6/FIG8
E9ZG4D93VlSAo513TGfAWw9Qzv0Me6Eoes/TRl0W/80ZXo3tbw+i9pbbq4OOIF8O
LiK2VI4xFgMFb8x8aRaBiVR5cWwYtgTTnGyJOwx9KDFKyyiiL9LpALWpcaOLJNsk
Kr15BztsIib1Dl8nlTBCOJGeQxo9SvhybKt1rhhjx6+bpN2fLqvrkMjHcSssLVDj
x8RNQ0PeMWyvDI2F4mi+jrD1ixxddN8MUI66XDm+QwWC7JqX8XprO0162XQ+Aunl
uJnx56bZjqLVjyFmzUFc0DgrDLYXd2EDK3eJ3z6cvsuB/qK092UgML815SegKYVG
y4GZ7PyKv7qhkiDdxFy4arFp763KQeosOfaTBIuPD8eJoJ1dVTP1P0sQyfTPuq2L
lBiDS8Wi/xFhdD6M8Qzwqp97UFfsVqCYIMBSPWaTeO3lOztBZCz7f5tjNzqdRdWP
jHYytZuBOsyDE3IQsl3YbTTQ4HAm1Z6obySB3qQcUwc63CaE3jtGDpqMG7EKHZHi
D7TQEM292G7I/G1ZCOBJMDH9NcHvo6vljWhfPBn5w1lTipT39+fQbsdqdFUR5odA
59b3gEdFmT5jHz9pOzG4kxM4dR7hUSsycjH5dp65DPJJ5fFb8JHZagJbwGuG2y8g
onL54Ccpi1dY3HjfJSCm5FeyNRwV5NWc+wScRKM0dRy/nwXZqEzqnDjn4Oxwaq1E
Z1Il2vQZQDhfFOs5jAtqKpkahgKG0ykOwf6/LkJkrKtrcozaUJpFABEdWkK15e0G
F6LOddvCG2Mon9gXyEbzVA==
`pragma protect end_protected 
`pragma protect begin_protected  
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OCy0TKOikztW6GwJiO192Ogkqjr9DZDKrT3UayYlDeZFnkjkyxiUFxgwi5sHPuLw
IcgwRbaC4/r+H3oIMi3ICy2c22WS0eTEnzYYkPk3WCjJ+gb3rC77g1MLSG9F1L7z
lVcRVBJcGIBwzjqFzKpbI9TEP7/2ACN9lJgSgZAHVVg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 94311     )
cIbQAcrxzjhvqM4iBN4SHufCTvpz7nh6O07EnGL0NI2maUBTV4zj+KeYEtKuKn62
YiqusLr+Kc7dTK1DWHPHS3P8IhG57JeYhhPsC3sGah1lOG0M+S8nOqqEnepuD7Q2
I6EdjoRQC2+g6n35yaF4wxmipjEftV/d/MbtdMKY//A1s8uZPs7Lld76tIFd9Hb8
W2yCKJFjMEDKOVBuO9L5wvQSL8lzm3t+Jz3fSd3qdeIbamhcnjvnVAcx4X+ZVFQ/
WiKyx+bylTP3elaAxEw3Nc0nMGNFaoIM99DJV216+8tKKNT4kwcAGq8J7nTxbW6w
YmUAnuaHwkpMJe/e/dJmBYms/qkkANQnnb/Tny0TY6lOji5u+tr1OXPGcO3ZeuUl
BQ53BB0kvHWjgqwDHtMlyJRYVp43uL3HebFaNzzGhmR6/GMM21W72C+KlF9LwfpC
dAp8CnspRvuqGIj15tzgSbnVM4HsIxuD1OfO3DliQCUIWpZEizUHIw6JGuQFBQ/O
Yfe5OTwS0usCohWhBKAJIVtz6g7SzkWP8v+n8k6L7HY8HVKGs22sf3+/TlhPTbgQ
6lW311V7E0HVdbgu+kcXuDHkuoeBAPQA+7qMrpdCjT89Oa5XS7VGbd96K5unLe6s
RwIrteNJYiBSR1mpIPgp14DFk585ZWdECEIv14wQcnFBpAT4gE6UbL/ZT+US0bpF
sqX3NjseR8VSnG9M/T1oB1f7xVH8yLyBbVefMTTjSoRr/lJnGyyXoRCNCurNaahl
/PylVP+9TTVPtRcD9pjC6fPWFMSpgplyZKF+V2nJQGQ95JE1SwLQ9tnIPZGPYqD4
bYsKCdHbJklJZngbzatFKIhU7mF7d8HV2U1k4IXUOoIde+aKPsNXt3kUfDPvUfNI
J7ru08r8Trcaz8LJgapVt5FHxH/loceVEc2xnuWQKI5HjOCr0bKbzhRNo2CE3nBj
hYy95ITh/zSa1SDfrT7WGj9gK6dzvkqQI3/wG7o1h4LWOXWu2gK+lyhN+dwIva1I
OlsExCiuj/bOHIGYku6SvtMtS9dJ3r1zbwyuAfXzkunnp+D663oGBPIVi5DbPMWH
Ev1xa14QJOXU63y01DisI3zjTONEQjJvUX6PyDDgjfKDTQh5CERORnAosFS/28vV
o9pqtrLsgplxbVd7bxZ5ZpVZzytQ1ikBunYQbCiu5fYAa9CcAhCQDMjN1GixO0Cl
4BPbunbZjxAA8Fd9w+4JYIq/sZ2g7ofCDplSvYh4EmP8PP/hXO1dbxlyra5jtZ8e
FCXKTWnw6/Q0FahO+uf4HTyCiqvyvAX1ZtqThusspOu5MsTUjcqDah/4fcc3Nkcb
tzLhr0Ig8PvyGIZEYFYd8xOTZ+MYTDPcLJTl7X+Y+/GcEHW34ufEuCRS9MXqFqiw
WTgWrfv6YSo+n8i1G4R6HITcg/HTBxsU/G0Tl1SVchP+y53NaQ44635ijd+VFBVm
K8uzEvaKELAx5XCvc/qqBFIlAxABT3jgONA/dN1LktVyxA3lHTY2dMpGPcdNIOkp
KNwyfiKIL93BnLvl1ha+ddbT3X+ml6+WQb34WHFxiUcxrPmCARL/Q4lj0kgFlWFf
WYHoy2t7Gzhpk491GT4tJdZGP351vuhMXGGC7ZcdwbQr7DPMloP5FlTQYl86TKsA
vEptWVo8pFKcWeJSfYviqoc0JVvEjRhMdIDCO3jLp4OLEhdUUc4edfx0Mz2324Cm
ekbe5EPgI1X/S55BaH/9sA9OQ+Wls3LvskVO+PeuMp3FF+RRFRoMWgDvxGuWvbTX
F4w4B2E/c6sgJ7HGO7Rt+QWYfrR6sQ4cMaxS/Q+8ZSiW9SSC970ak6I09UAQnmtU
FQhYDHiBwzNN3y5rtVmc1P9Cvm/0Hmc7WNY+SnVOw3uw8wnenkuXaILByz0/h1Yr
SJsl1e7eHfFfft0mcuLM6FQuYPBl62zmFWne/wdLOU84t+5ujw4u6ZVCEvXE2Jn9
uK/ttIgEBkZi2PMNu/5wqEgvl0D9bd2tsKuAya1OWHpvNbyb4zRRYPM+8LC0zbd3
+QD2u7xu/UygrlVZHvX5zzCYlyFGH4PbpgnMfdK58il5YzFg7v+MIlxVHNy3pVi8
SrExgUaCeUvellXAb2SX/AQhRtmy2k6JNKlb+4t8BPTRR3HLpxkv0WSABp9mpk7E
`pragma protect end_protected      
//vcs_lic_vip_  protect
`pragma protect begin_protected  
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
SGnnee2vi74vb5/LgfmQJOcncz7NAcpvt4ZX2kOkJ9s/VFELkdGg3xXUielQbQ7L
7B7UP4LSfT/+cpy8ekCHvV+gKmE1yQvzd8kB1/5qzmCkeAVdmk8U5XsaazrTGpra
NhpK+GMQl+PGclunATroXU90KLf1SQize6y5NFUWXuY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 109450    )
qct9alMCdpJJFEubhQv5Rbx4ecMKy0fTVXEDNddCdT6JQ9i0fidvH82AiTUlhJG3
w8sTuqNWWvXOP7/QdWG3oPJ4OYMdbt9gDWE3T7qsZX1zHHgpsXN3f7xcipKDIq9n
LSWHnnZeWcV9ZnU0IVV4JASiOqyvWSLUgD25qvGRZTBB0QrK3VTLg1aouAVnUnMq
cF5w19USGhobbyiy6nsql+s5xWFJDQIi08ydP6Q0JpWNbzuUDfb9OdpBvf3bzioB
Y9zbLBbmiJpgy1KMb5pA8cjBD0sO/bVX+o6WUN6sqtnZ87uoAacobKUuanOM6Yc2
+urN1E++/9E9FSm0dTwapTOa4mOcrFsJjCZsYs1JwubPBRNiBcC5vyjRyU9WHZwV
nqJ5NDo2YJFtl8aIXICN954/2gDjD0uARFeQABv1u8OzGg6Mc0nPUebmyD4mv0ed
G1K5yo+7VCHsrP/Gb3WgyYK4qK3sXU/1IwRzTb5YGocfs5CKvINQd78GUVBX7wg2
lLK5D4dRnvaE9ZI6+qCcKtH3GqoZ8mwbFrLSVtkO+EKEGG/QxzrgZpmtvj7Q+AN4
4iZVdAryvnOG/G2Ivm78GovxawfpAlfIgPxWxf9ND1HDKSMqQcJ6BxvsxcK5OWtK
lnzCY+NuFSVx9HZWbtJ4Tg9W5VSP2uA1c2j4GTBub+NxQA7x9X5I4FIUhOk5HNBW
Oz/cY78DfJb5oXAvrgM75JqltXIaLfmjhgZ8HVOAtXRypAT5wuNPXXY+ChkqUdeX
51G6lN/a1HapoOSfj6Ix1sEmdV24zFwcVXLsEMeXRQNPnveDa6EK84ynWYaFkzxR
z8kgUlqO7vM+WkefFJVEEfUfQNjjmZDuGmkNX2sKrE8gKbyVcOHmot3A4VZ6bZL7
uqPfpwtMNqd2tExq2rOL7zsbL2mnJRb/PQl+4BOAklhH0Jy8X/oknObySS0CKhkm
WNmU5G+4Mb9gttCT1bxA3RlfB2jMmzuhzMIUVzuBokAfSxeeVUDcORAzmwbTrPq2
cSmjq1HK/5y9/UcN9j09izuLAt3XKQmYqxrzVllZ4bFt0DwIbFPxPVz/gIdGjNwo
MyjfMuvRCZphWshnUolFrLowvPqoezJrzLqKe7On2kvUVZY/YgtVzVbkJAU5JYKZ
fRmmKEN70tWr0p4H67SUjfbLOfwXacl/JdkI/iRDPgZM4jySvmT8uU6c2kXN4w/D
1KnQjEMF4qhTOueHWmWJ7+h8DIXHs7SnDu0WoYCl5LI19+zTrOX+xC9bfubnVBEH
Lb+I5dYEfiulSvNsRmEZNWJjVgvFB6f2MuP3xynSaQSQYnFzNrtRFP81i1vTSYTz
Wd6KlYTkCft5A75L2a7zHPZucp7pSTVWEzbceRHqtfSDtdyY4CE8qQ7LAOPMrzWS
/48tNqz/1v1raz8RBajwqiC9rjWEXbU/cyuGdgcRKT2pAv8HNVVvXCwq5qUMlrcr
8rszJ3xxHQDO7DUaEqZJnEIjeV5sk4w6zl11ztFGi4+9TshdzHRWhjEEsy3e38Tz
5NB4uTMMdaISzbmBw94kwhpHUPlfd37Y9cv5DTc2+rtOYtkgOTuMMN2rdiiQ1Niv
99fXlPEWi7faUvpwAmI3SHAg4FijviAAx7HWmWmx2NV1MRBrO91vnPbPt78EklIM
pVFkMbNzvKpwIvQ5cJS+yiU2Z76zePz+gbJP1tdEbD5JEM4bh9Ngs6hSucl25QHY
o/KgdoG41ruKI274vprZwT1h5x42Ls7gvV2frPpllSw5FT+h1iYX8Wy6eIlsHi2/
y/XBToyIzpFd3J1cQ6qfEgIPA/81UsPifklmtu8HBhAMAO2Pp/JAOrjYDcmQAbDM
M+7tumtcdHGr0NyAdU6JJIXeowU9wbYsThhkQqvNsB44XudjBXVj5vNDe6MGKcsW
szn946vRYVXpRqn+Zb0tRWzeabSCPB7K5mAngA0Y6IPzMekjAtiq1ohVlgQy1IZ3
PMGIKCRVKe6/KhDWPR+iZMJdWSYPy1OTS/mC9fROQ55d2S3qc5YtExQcSsrGBSAd
H6fxiKwFgU0REw7swUBGUleSXWVtq6YFcGpPoZ749gwcUqcqNvPUch33Qhmbh9v1
phmou2EhDaUxQBfggiZDfAf1sJtOJQLlhfUF6kGC9no71i1jKkA2EA01ogTTmux/
6VzoGWbOd1caX4SITXUmIt3/LkSAbYFEZEgMBT7Es9xw1Uule/JQYTIM/RTm9x9r
ruj3NadHmA+X1GmS/SZzkK0fb8NMY0ealB9d+Lm3yULr6onIYotGadGBXWu6K4n3
CA830HnjWqWZo3nCjNxAcecdABIKZwqHs+jngSVm93noAAMywSiJuTJa7u1ukV6q
lWVkRWEDy88kZmDmp45xMx0tHrE9ipjzHLtTTcjSn2Y5fswCBad1JbaZoYVmkKkl
Y5NU4fLDgz6O+q84IAw2fYxPNPEc4wj3BzAWWSFjSv9z9ObCBzQW5SXXPIj7GRpn
vfS0qIQ3xTWIG61wml60XEzvPAIuXhuOzf8dIUeG0eBpwBDR8Vla5Tjre8GrVdqf
8Tm9CwT3ub5VX+3pfDbu4y99l8KERK/c+AhnTXYkL1ip2MHZhG6/oJO9V65qtIXV
wEOYRcVW2WPnBbCaF7gjt7WNG9BPNEWIOI4sr2qzSOOnCF8uBDHKt6U7k2Ww7iHQ
Pvu4yf+c5TvD+CxtYbA83JCBHAH/w6GWfzf+sXxncw3tUo3qTAlwwcOyyLgLZ6zS
QpkYCLfUnWSSzoCum31/BbkRpQgFTxn6tORsSvVOYlguaznaOpNX8t8S3AvlJp1O
sx5YHgQ2gx0aKhQjKzup4dUQgccUeRLN3c+IRTkA7n8VSuRgTyStt8YyjoahvEcw
rwberZXf+9AmMq1qrBtPZd/PP1ZXOZwOXTJCCe8bDSWcNtgmMM9U6116hoh5YM3K
5aWenlWOYkCFQgsEmJVA90YELW4G2GirkEE3nicpA8MKJhbGqADMOpouynMSu2LV
4iBo9QC13pK+0mdMBwDpAiGvKkBL+iuoNo8unE3mz2ykyhKdSK5fx4KkMi199EPs
6XzW3jPG00RJ+iPAz5IkDg/+EtE3RP8dgulVnQBS3QCjApyAJOZhprLoKVT18pF4
X9qDhaUUK51afMEIozM+Qwg/ctpu3efrHUjXv2Mmxy5R6fmjioyqVoA4/BJNVMye
w5ifPhUwacLzpPw9ubeeDvD2sDBTmoc7meFIOVcP94y9uEFsEt9vTTj6PnKW6SzT
DN9iN3rYD9tk/uqzy6drqK6CgYo7LKut4TC88SeYdW8EBAzyS9jmDrev86T6wk7O
/SZybD/nGl9n2CKZC56udEdO79NgFfGUHh8i0tzpSZi63I4H6YLJzitAdMYcA8VQ
e1lV127Dfkvle3nxvnPlS4B/ckiIlS7AnmOuIWn+vBKZQxFC5NHKmhhElrEc3bCy
NTC4M05FJsZJiGIyaZwIsY9v/aucDd7GsVTsnxZahFsMYikRrk/pRSdzRJ4Up9Aa
K/BRNxd/AA5ZYoYunLXs0W56RocMfHo+Y0Iswf/FsUlOF0JGSCPkQ8RvMI3spfMK
FPZVeU54oFsDw+bhcjSY05dgvoplvzIV9+jISL4OsIv/9aVr9jn9xRhWt5SvftjY
k2ob7DFdc627aSKrJOy23F5CzsBEUOMvUq2mnJ1mT+CmHTMLeDNfs/Z6yGq2JaXe
UKoZRxfU0b9cnSRiU49E6XWIsJYCWz9bOKI0Uc1RyxNO1CoN+7TvUVCd/06bg9VU
GkLvRM9mysl3hIBp5VZDBcVgC5zM+KkUH/SweEb/Dq1AkF0uxgnD5fyAXVcj3b+B
T8qNB3oNZ9v3i73sJ3Bv+XnEEl3If0HQ3SyRCbBSLaF/iE4NNHOFVkAhmDU1sBBn
vgz6Re32qPHdxv1xKH7rWiNse52D7c8YeiYGEHwSA9dqn0sLRPiXFjMKwNylSnVV
R4AjPbrGoPcGenxZx14DKGurJhNsmeQhjSi+k8Gv12kPS71DKATE7/GsXdyCeL76
2iiT2EMXZFG7AQ19GZg2lvpl7XLZ5BRsuARAUqJg1lYxHZhSGg6JOW0KmLV53SWC
1vBvf2GdL9SyqVE9/+mPcqdv3WVKJE2ZrI+WqnBW2bft3XzwGwPBAqkVUwKMfqUh
7G0hEnMQaquIgS1jAgHyj/eoTF4IV1oXmu9uRjybYxt37dxEnlFlHOFU9JZUc9He
DlfgDbNAJycKbr1aqUkuQW+2PlIwpDR5YLnv6z0Vrmjql+FbwLVfoWy8biAyzFyu
Uxw5JGtuIckKgD8l3081VJ7pihxyj9UKbkdbJU/NLIKJPDt+EPUYyzWPQ726QB2j
bya4xp0ObDBP5Htj9Uo3ARQyvnze7mZ9IkwEayLfKW29rti4pcozaTLw69NA5gbg
WtqPUbm+g0kAxrZsSvHzhlU5YztuR3TPQmDjEw934iSjsCEM8YIjJKKV1InzvoEs
bJpWaPo76OmVjY0N/ObRNwn1yK8yJQWWt0xOX29gVSmgmCYcdMjJHfLCaZ2aE7XR
/YMtFKOSy0txyMyuH+uLdcHvkQCJZvcntZ+k82JcUCFhNS+cdJtTGC+ULziWgUU8
bUW5CkfdEm0JT+luUQByj9gY1nlaS6zEhcWSxQXt6IxkTaGAt9iyriL9eP57W1fn
TonniVby5vIsB196MQe86hJlS4swoZV97aG2Cwmb0mUYYm8Zka/W/brV/0MJgQqr
SMJ28W04A97Ye+9kqjZxuW/ajF8vrQ8ewVaGVAkmv1dIUmFSJ3cuGr8GXhrQ4TOD
yDFxeIgz1iSxdiv2LnL7mNhRfQj1VfclJ3sWaLybOWfvtpUAbZzzaXZSvtlMsdR/
s39xRi5lnT2hk6+Aiqfzdq5pW0NxnvI7zTTm1C5usNzxL2w+JHPfB1aMsbzfjuGA
mNXIB9j64cQBCcj6J2rHLpCN7/bV2Ww+N1jR5126hPgq4CLlMRT2qI7uJ++4OETj
3mTAkchRgECKYtb9gAVO2XZIluMwS9C7h+7OAn4u2zVcEgntASAL42fcAH5tsu7p
oMFplJOGhUXS3brKjPU6ZM210NnCR7wrikWXGKbnQo7uMt6HAR3YihLGESzfN3Vi
sPF/izEgA/3yxVNqRlOq6SS48aQD3VP55wpZQmwveGN28VJrrIzFuEI2QLgBr5Ml
fZclENHDH7MUC+b+0xxDdU9KtRc7v6Ma9gNds8l1YShqv1iAp36niT6Fdmv2zz2L
loilcrl3Hr5hUuqo2/U9jQ+myNIcDRb3yxuU9YeCGNvZtubX8957hFrbqmD8xD8N
I9aL7Y2D7tpTG9VZJwQd6saDeWBptRC3sEObK0KI66cEpuLFp7ZEPFFR6Be430jE
6oepfT+c4gmt4OC9dq2QyTjjiYgcCw86wftr/0oFtHiqaNWmz5w3ZDniB10UZ1oR
ZbquA2CYDqR1ZuKnEZAunzxzlheZBzJ01fHf3Oj1ahx5DYZdBbRh9dJF9/UP1yuO
iFdhpSnl93xQ1ct0qrU+23pYWRdT9OBtLPqhZojGk5rlW88+ZFi95EaPUzxTF+WT
YBiir5Qol1Rrh4qJD59rUK/GGOQRL6VzN8LNnDh8Q8YS+BA09H1jvTJytSvPqLR7
9UdZ9ppok0s03YACnm1vZNDzTqCos8DM22Xb4Ucan4C0/dUa5v69uJLdlqJjIEsl
J32OHkAkWWQhwl3+sPoIDZNxsV2ZVon9aQQn0d+AVdsPXypCsxne6N9adNtLIf9r
AM7tNuZ56OE9Sm0rtQF50K2tkQ1auSRi07ckAGrm1wZ+X130xGPqT2hb4yGkQpzx
sLPsWIQQdLA4o8cbk9Ikj2r2JW84ZNYEF3h5CHyOwow1cBfAHXnSBaCC8rI0jEQx
yts0/Uuwt8TeCy94GS7fbpP8XJZ81rw/4xY0TWvd2iAfJZWfXizhz0ynR9uosR6/
NF15co4+0eMti98IhRO1nTfcejjCNexqu+xDBfvC/uoScSUaMOut6Qgadp+2kt5e
j74D8tNvo6Oct8gfJRODb2v4AUiIOzd89HLim5LwYnoGoWH+gC/4en4ihqE//3mV
wXw1lfm+3yYuafJ6AOtD8bSeC6LHKTNUWwAHQlHiT4XGOZBn7JefvQnohKdbsmZQ
mbFclwLIT6IEPNMfXVLs9px5iV3pKw5Plp/37dglBIjLr/hE58YWybQymmQD26mE
wxyQBwGjDVXbvfUOMgJqpCV7lgYaCs+rcoarnRXRtFLfDJTs/ELmxojyN+8CRJG+
ilB6cAskw2MyUN0yg2txm8eLRuDq3nbMvQB5GTMpupgwlkkRy2P2k2Q0b394GalX
+FzN4d/jP61pqLO7tk9dzprlJMa3GXJVdo/C+yET7/7MMHB+K1SiwGooTtglhH+n
4usMKV692hcpUt5oSXsULGU9O75Tkuae2I55G4rUn4fD78dLJ9N8VAdbWLi6Idel
DPUQCi25xovfYLFsZNOUkLnBIvpEZtSU8TjKj8D5k9TVr8d9sOZMmy2QYwvcQ3Yr
RQ/ns8co0y/VIsyhVp67R8mgqvrDVEUSeCbcJr9v0yJUSWBT1jS1y+haYkn/MeiA
O5fQDYkjNXDrZ0QAMpep/SWSEp5w23Q2ejxD8lZbuhd8SEmzIo3GxNewU+fXz0IR
01HcrjsN16KhGetgvQ7BH09e/HRIBmuCSF3ub4JFnEEYgh9qYlSljCi06UlJadI/
ZySt0pkZMuvmaUG2xxjfu3sXbiald+xBoxqwWAIsgxk07dy2efa12KZJk6hy+IHZ
w1XgaQwjxojl5CG9Vk/fw4CddX2zFgS5cT2Y5FoiZEAdw+Ak2p9MNnNqD7Fx8rsF
gBcdKUIfc58/8BUYCUzkrhRggaJtNvU6AhQgk7KHaVJccelNg96BIL0D36XMft0v
Q6NhgMiZDEPZPBrCMC2O2+xSOHDKLP5ITnbw10ReCcDbHfLT/iX/3ZS1NITjE4Yo
13VjC2UZ6dqPh05HeOyz5VHM3cNKWLorAN7iWD2FBnOdyluC3xDdjlLyqeRqnLGg
ipLEwXGlpccz5iMCcajYvdYvMwhXUaCg0jEI5sZgXoruXy/PJlxeGiMZOD84QH10
iRvstOknHzwedz3ffOT/gwf0KICVMn+xIcQ2vUmWcs9fWC+QG5RqtIHrIa+dQ4ap
ptEOxpc86o/1MyuuDku3zICOUEHkydm0WazjTyJR/xNnfRubWa8VdnzBJWgqUNBv
DZHBNGt5DBZY2sqbiyxVi8stC906RlyVsrcUKAQC0WYgdIu9bfct/PSSlxbJEQ9i
SxUAhFVfx9ZjwCaJi24OK4nL9urGFAI/JknqoFprea4lIZKpZ+5H17RkfcDsdU8g
a7EM1bukym4p70fBLAfQ8ocOtDj+WJE3aLvRJ6xptJE/osOoL/33d2+TVqgMXXNK
NAviIMdDwZoVvdoJGvXeaMjQm26SeAUeNtlyfxG1c1o1u4P2EoVvNjxwl/vDh2Tf
ry9uKX1wz01XwIFLWs2ochyC/eeZ3JcmS3c13WDFm5WxZU+PWkU5sPIeXzxTr2sV
p8qyrNMC22WU9KKDt6s5rOoTZTiRHGSWdxGuhucb2APpmDOCbO6m6deH2wpb/5Qi
ABGxoONPyJzliD1hnVP9B+cRe6tCjx+j23NNnV0C5WQvn9sr6mB6fFGILc729k1Y
/hqFbdDSdOtbI079IW/vESwOg0b8eQyHXFVY0uRkVgL74UYxEcCUcIAgTTZEvCWN
j2KiMaa6c1Vqk4Bjt9XhBChP9FJVFpILxdcVxRwG738gJZ4My0XxuCVq0DyU9QHZ
zUQKNTXQvIS3ulf5fVXUMnxwh1Op/6zSEItEE4rIAqd4foVVM5+3QHx25bow24yg
HrOEFODBQLnWymEkuFXhf9ThFSqJfA9ZvKa6SHonz8lxQYDV0vbnNRIyeeW39HqB
p8fjwQtAzcULKUzU4J9aZAoGf5dMRO39lHe7pZ86+Q23mSVMj5h8Mv3t7V95NiAn
04dwc+zG4RO5pMCb1KBb3JN3Agth2TFYNQxGcYTvl1bHV9KIEZI90+VxoPWx9NB5
5Lu7HAfLYg/PGA/Wvw17gP10yyN32TcWX3+fgsGJPx9Q5SgirNM4LrRU2Bxdth7k
5dbeM0G7Ek6/0wELifPs4H1emk5bvLSA5bsj8EEs9suBuJI2m9aKAQ8bcIpMseos
BWozKFEwTQjUHS5S9SiZf28amu6ie47UAkXJQyP6+BhBx3WXpagNlj6Qe3POwwDh
EOuWQzYdcVjMRt/21U+SIbS24OzGNE5giSzhIPMcHD6GuolkDL0HiIjw7nHg5qUr
wEnU2rcYvW/hUkHg9+oEKT9LuMDHbYd4LNLB4Jq0Mm6GsykKiA6rujPqoOjr7r7a
+DmAo1HiywvqNk1stpvyXUQwnvUlICqLTAw/49+CqeU8Hz8ADeHXOr7kGY+O3012
k/Li99l3RCAI+aXnJ2OBWYyfiIqcRPAtzvw7YtS/42t0bWVaqQFfRjLyLLfU8ZFQ
2Kn2z5c6o/l16DhFDslj0QmY066Muq75sp6BSmxlRYruTo775Gc/hDyf0QQwXZYX
Y3EajiimNYgKzHXZMvIkfZawdNH1pV9fXeRnmYTMwCULTrSAPG5kmVMPV7JtiXu8
TFXa/p1VKEhTPeBNXaVTBGPU2Chh7dtj3uGySMQmqk8PqgmkOfLLHidx5d2p6Esq
oNGZrh+KGLS3unGFmLBHQwrtR7pR/uNKV5UBGEjiaBwhp1GVQrGfQSUwfEy6J0ev
dLwsqrHMjRjgz+vt8Fz9TjRITNthg7bZWOicIc6LgHgh9fIeOt3t216UaaESohzh
Ze5NAERCy53Wr6hpUVFBDpKYxN1jAWDwxPWI2kBBfvOjQgX8XrnlPcTjKR2lG+xk
Ur1ZhxJExYXl7xK6yPGLTRboGf9yjjxQYuoH1cY/QYXiA2HqmvVhKoGGgX2TmHgz
o4qLO8w8vZ0UDuMUZ9HnLgBH9Z0Uue5C/X6YvJrXXdvlqBova/sjSVfOECem1mtU
VhRqKbRF4KwyyKu1kIyT3qlm/qx/EmPCdO2TTR5oWbF067BZ5fsKCXdA0zyIfP34
2M75FbIKVf3+PqsTjEUu7j65UNcyO9hSbyJMKGDLNXMlFjfUjb4HqS9DBiqcP8OV
uo9Jn+Ra81tYKaOEwz6Q6lCW6ZSYomBiTt9CDaMM6CA0yKhmDc+IWhTsdQBIZPgc
Zyb0hgQDo+peyI1ktYTyhzcXgp/M8gmCJQg99YiJOtE34fFekVcJS0QfEiBu6eze
Qx5cgWyZjR2zz3eGnKz5tFrk6weEEjenpqgF64NaKWRteL4SFGQNFu9V9jdBVEw+
mtDeglvxO8fZqdbmj2dDqtlr/ei6IAj/odlB12VlbWMmqAIYEimoXXV845D2wNHd
2G3NG3UI940ymBeMTyauWIyeYh1Jcyk0e7MipWBWjbNOi6BFZ9YQ1eUZkgaWaV2U
YgC6Dkgv8D0jsa8xXk+b9i/DwU1AHr6Q+kffpGX/8CFhlKjBwCYVBgs04gbhMvGs
Kjq8oKAB2+Eml+3I/wimYAieXce/5cOuCWpmwpsnN/SWlURbMZR2NyWpdw53QgaP
Qs6tv9C8puIZBYYLBLVyZ5ym6Te1qV9C65RJJP7la8jx6oI0UilW69rOjXozSpAc
vPUK9ac7oEGI/nfJZJ51ATF0TS+xNVekrQU4uLICrHPinFsL64WtOZgiP28oW7BY
IkS1fmcmJtylOwn2MTUHvJdKgXbKQEsBz6Z2n+m14OZyTWdW1UdShlr7YwUzdM53
WADqyxV5a/BnJUDxgA+jQId3UH3j44IZE2qDNClgsuyR23e8L3h7U3cWQuzinO1L
lyJkSX1rLOOm3jM3//Oqk7lrbFmJGq7fgYN+vC38gzx7hbyjwYBg89alPquAXTnU
DnTglaqmYnaxnw+HdSaJXov9OLd2m2PgEi1oQ5N1PeIsgjvHKf3I67BNjaq+yHq+
+pVKvdfhVc4XlXx7CvUXI1qrpfQdgpe+ZXzrDxlpGabqluMkTgRRCdvtXU40+1L0
mTO527TeAGQIXxyiIJtEINEUtQgX2ZQATHHxNa7Hz1pPtWBDuQkP8u5ccrX1bt+2
HSMpI7yEsY0ocmuCgvzvZ1ZiAhgHG12t6I/ghaYMyOYYvQABBYg0M/lmJjwqzMGj
Q+EXOplh1nYi4PmLOTe00y4mW2HzXO4iUjiDPbq4BGAM8hy7tT+ItNVuADSpSD6l
WklA+9Dz6pypMLKxVjUZVNRIzTPSSQJgliQKBynl9P73a+BO9AgXjSZq6CNZXdPH
l2EKqEoU36AS9ommFJjMlyGmL01eHEo71kzLENU3ZsA8Qj5LVr0c1XYtOaJ753Vp
+4/gC66M38w5cZZCw9KR82vvskZNuGzfg/6aAV2t+gPHNek8WF80A137lRglSBpU
e5zuCBxXe6hw2NPCdqeWyitgPVKP4+LdZLLOypBhmLSwGfUsy0IU+CF5x34MfeB+
fbJSZXvuvFodh/JgquAfoWNp7l10gznzHMfiQ6v7eSMWp+fdmUvXxaQiCNAAgGfw
qCMsPrnV6PVF+ZxVuzvXJMqiZGPbu6BRXCQBNo7GFcMSXSRVmWnBgVgdDr0vVeaO
BmWKoAPXBjtG7gW6b2W0KbAtzxYqWxUaptIqLho8oKZ+viyUgi9Laq03F5rM2QdW
SwgYzSjHPlohjpEUPava5khbJgWmetNs1qTZ3CY8r39hPaQ0fnTiHXocxlyhr1ej
u0qtErw+i5st3oQkVffNluVi/90+9uIoc5jMz0LJokDIBNYp6lS4BhgHODbbl0/H
sUtr61d7m4oGeDD6P0Q70klWAenJ2Byol4rUZn/QBJ2SGrcX9Eb8dwKsz4PlyK8k
+QhDQw0bHq1rsFf6V1bmc24hbQyt0dc9wnnLxim50KQG57aDo7NzxNqBDdPpG0S/
7OdyOs/8aQTfzcO+ZPaoDqCB6esJobomIt0wY1Zp0VC4zJz+O45V6KQhzu5RnkKT
de3Gs4o6oFEk7VqhWPp+dX9/zHQsVh4DvCO6iipO6az2facFF3pkpdjAHZv0Pxui
4cNhfySAX+poEFX5DKcoss+ljYMxM77rJ/JN3ntmauAXnl3xgYjxDgQc9jA/5vkL
GhiJC9G01YbLbbHDvV85TzdMFDmHfwTy5tW1w9KbD9I9AenftpzQGuR+QbZyBnl5
eNLPaPcMCptf5fdN6ysNKQl9LbDYfe7sTna1O8HaV/AWNWxsmKoaUdwAdSi5jjp3
sA1/Sbk1OXRynNhs5Z22/jUVzjpQyO/olmpfmU5eOmZF6OhpEOLlOkXVVglAByRt
YqgDlf6q/ITph1L07hXmzQsEVs9h8JfvAx2/grOcyFaYjg5UEfE0Ohr3joWFv7TC
WfNk+Watffpf7wuVRS52ErvSnZD7HuUecfWA2VkUHC4gSSLGVk0HdW2X0colNDOs
KG8p/KdyJMpzpF95ji95iuKnzQFHWKU2VE9bo7L5fh/awEksnjJTvkTsWI4RwrVK
Woz2HvMnEUquGKRkrBNltIS/nooki/2s7gojpFDAPJXy4LJXAbnxwv4PZwZ3brr8
5+82cf1Bp373B0KjfT1w2ENXUPVJqlQx1sGDTe/SBigIoKGzN//iGcRL3K5Ne08/
2XzCowulZqcE9ypGb5JdHYIZ9YmHe3AgrXqg+q4F8dmkSfAkjceS7Ihro3nc+Ij+
pX6p9g4kasJZCou5Xhk3Zzv7dOibwCmhf5/MBRCxwjDRWRhAP+m/G4hBGfbhzOdg
AxFQ8RXAOdgIa9WwUcZ2/0AYS8NmxQm/rZYnrq3E3BbSKasD2CfLL79VX8LCBESe
HYVWyuB5y1shWlgyKbkTR++PuXSJwnFARnpJNT7RCaaPuWAbaNQ5OLFfoo41gnxn
bzCIvtsQqpRUDCzToxceL/Kd78OfleUYLhy+OXiHCstVOb2jJwFy62ST+NTYxB22
pMvNPy7ZPvu1l06fehHuqzaX8jH/9l6r90Ttu9a0fPB8UB8hYx5tku6BMa+BgKRY
QlkMpkWwumQ1ycg5p2Fda2MGIO2YhGBbBlAfgWBdcpSe1goE1Xui26KYyfI6DT5l
a56SDFtz/9MG6CHF6T1U3MNtKUxWp8zqtS/Oys+uiOfhRNidV3IETXKfaE7Pss3c
6r5tPKJfcwt7tmkR25xkKYgFoIHsVsLfsPivWQ7zfL8MzA6arjYE6adYYTj9/JJJ
z+Pl6C3+vxUltfFXXUIpaT6xuYQZjbwPYDFmQNY0QajEp9wtR+FM/uUZrRFS9imU
ML+22NoJu19VuArsE2bI8H41Dyz+Ybd8vVFa4ecrxSvwLILLyVJG7N/SasvhOYP2
jkb8C3Kiuj7gT3hp5PIYqThWx3t2UEobZRq6RBtlYaT0LGIBFg7Iqgam/QXfDQaM
yd2f5nynyhEzj5hxxs1bjsE6lOdOimEZnAY6BwKXZJgGIhB9drdZiIaScnRfbOqw
SsndeL+5cJhPrmcS33HRH31yLBh5fRT9AlzYiCcuzZPiTX2TUWb9cUudz8a9Mqm8
8bc71ENC6Ckh2mqFQCcxll+oEWaamRXwrzvwXmROm++wDojFSxlBKrh0myHasbis
87RRN5OPY0by7uUyWqSGk2OhPVBPoxNvMB5ZZzDlmclz/vE5baFnHR0Ocwq44NI6
87wIHj3c6nzx4BC9+SXo9a+lXk8Vid/xglbi6gxwOkkM9cYF2MmVPsY/KhcbKtZ1
d92KaRWsvprhIFFhmc94d3T6aM0lwlohQIyQF6QUUOogwyANlGmYBYR7K8quRPlK
RoBooVLyEw+GA+YCPcL7WpbXe59ecD1jAQsFQXqQwJg9yp57kjy0y3JPUhPxGv9u
g679QlhFmdUDknTbOe2IJyHJtrp1QBwUr60ft6Olc0aLV3q/i2ev7f5vhhdscSBZ
NLUZ62NH8dzYjixhrml8rD7yLjitPjjETRpvGLdwCmPI1bxJqqRdcztXtmB8U4gc
uEx8rI0BL9zKNAdHSiJyBRglbiEx+qUfTn49AXIHxhnI9IpNPvgX6bG/Yba/8MgR
wV1Ir4h2ihOdhs2+q5wlMdDH7qBhldj1uVLHlSMhsYMIycrdaBfePMGdWuTa+gsl
dgtBBGsyLUadSMkTIynMGMeXWTs07Gcw5XKwMgcQdMjwtIzCNfqERr54AIYwQTox
e9um9bK/OCIU+UVy9GkmPP7znzDXWz77RN1E7oD1lhKMMvuFSlGKA1RL15dDdSH4
NPJ9A5wp2PpLYdkcQXkItnk9lUWs71+4HUY6WFv0HYWHjHGcfdhSg8NvOWz7ujmw
qobjB63qc45LUUrMxJUGYDlgkuM56L/j200Wn2IyclBFMoGzANaVQBvTQZdO9HUc
s0pKrZoPi/3czDvq5ypx+Hj13vIMRWVMsvGBh+iSkEI3cp4VMWUw2YdStv+arrKJ
aSs8UtsDbPooHklWb0hHNzLyp8MIatdTAfssYRlyBv5ahkFrNB2iUxKuKlXOW7G6
P9zLMr4vqLyVzw8iYSZ1wQQRlWxN5u2PtDy8GRFt8O5OLzE3/qyT5EaagxKHI7m7
fb8mHwRw+jls3kZY54REKLxzzxN1n6m5K360Kc7OQVx98Qqb4OktGXMMVDDHfKfx
3jtlxDgSOfTD5dPr8xunhro5i0fOzXbQeF2zVYEW4EWYOL5w8SG28yRkvyqIZSDd
AMApnZ4ScroBOw6/tv2j67pNweRd77yiYxfzzxJeI0YgZKTu7WQB5NSF64T+vIng
DStC7MO4xMboJma364We5msUCIoT+A2c5bAxnvM1v2nRah+iGW3fhPTLGwmJ/sSO
UogWkQG/1tR3Mf2YgcpR4Gjzs26gqSYCM3fGGCJafOlMCTw9vQroYVdaf73nyPNQ
fZ7SE71x/xhqtJrejGRGoRUYhs/w+kibMMD8hLOammm2IXsDPZWOu32mA3bVCgSZ
UGTPiaYQCujD9jPGtB8B1av5+t+qefWtuHS21hNIXjJaWXWkkt/GJQneREVB8ogS
QtAH9bjusQOfxuNfxoo095gGyut8P+YFoIssQmjnPnyJVp6j57QNPjYjsYpGqexn
2boHXmttKm3wD/GpIylQCga8WVKRQyQYN084zwdZOMOygt0s03Ewz4MMDNpyJ+O9
XEWuLEsyc9xSwjqkKuzOqpNcnuN2bDP3InHP+o7Zu8j6xds4zh9BTs+VfH0Tf4ju
imH2zt5G0CEHU8q9ya9wrKQbcSAZNbTedgMFDUTAylRwIzLpLW8jCVjjJpuLNbUq
2/D6yIznfcA4HfU5VRc0yTvYGjBI/SjYfZ7H6ntQY3rfKWrbdzl4nztvAhOKyW7D
7rHQkQZmt0afHKqhinQabXKDDsh0YEcXX0/FUCU/KKdXTqA1QWkS9uUpJSww+HSz
KbRjyGr0PTtn9U94p0ukQaSwk5tVQo3VxHKn4/jpgKMR8jwOgrPNMPmbxyA7+iXv
4SPGcdjPar1QKO+ge06RNNhl7NuSfWLyZlOuiTMexGmxNLHLaKt+7uO4B8R/BvPu
aXKZc6oV3qeCyYvWsWImeE6LR0/DDAnrPhA+E+Ffd59RUKUQyZeg9yypqk+sbvka
n12vZWd/TZMr2oL08Cp7S9xW1zetkEYFfMLVR0RipdiWz41ptlGrNOLQG1TDlQ6/
tuJhkxxE0HFvha1hYxdoLwNKs8IzYAKzaW4VOUQsFMVLapF57Htr7ybWuK3WCVLI
XrLlXiAVcVPrwl8FIF/geKef0pNkoR/BFMttstPVuaI0g5CM2tyfUkKKN5wHR4rE
WeDJeP7PNgGXuvEab5mnNqQwH7N8Ds1CTegy5b6xVEOd3cz9NvjxXVGnTc/+9AMm
35VFZDGRsmWf0CWeeruGzsk+icoPRk0YfQZxNxd1gx2/jXdJzhaDMPf6pFfLVl2n
3apPZETgKS1IaK2FVqAWgOY3GjhLPklGl4GdeWGFgUNXTfwi9yjlkQBCqe1jlrCS
ZsGkl4rUoQR50/T4JWMv5RgCg9Gtva6LOSjw/WKP4Yju5/80L9YE8KN2vxh3KSrR
6uu8RLgg11+XUW0LLxDYHC8oTGFl0Pry3Jz6Boa31w742PhlV9BJ8iUw1GKpnorC
6e1R+0M0EcU4MBneuVDsN72kw4nSoDiFrHx7emdNLo7oUp0ZglPcrcTaU3Tp7iuO
ODxXkLVPG/lfqwNcQr2fsx9NNg0nlwzn1Bo+iY4a+FngwdV/gZfD03e2mve4dNqU
gFpdjO77hC0cY6iJJohTjlJbmaFoO+W8zgWhgrujcsD2+4E2mrSKkL+2tnjIjZtS
X+iTURBjMUBcY64BpJkiqAZZu9Af0gGh7myon8WFZ5VjqvjpA3PT8oQyw6XxEgIg
3Q1cz1IFejBhxTYCbxpEplQ0xl68tvaMosToffmS4NlsHUYkH02Y6t9adlYueSFi
fN3apuUJKSMHseTaGw6dyZnMMRsqjFnChnSztxeunjikVShpDPNdhnmj7cWbcCX+
TVX2x0uVi3YoR6eXyAIj2W730lYMPiC/4/9BhGRmunptiOqAipmQfT9UCPh2IQ2l
sUqtw5S20HtIpb7k2Vk/Qv2R/VGc0jx16OaZttlVRaLuMXo7/x906w6p01URoMzn
RRgmMpxBUWuvQibQhPQ639beDV4G7Cu0Rz1ydnLXyZmW+rrTzhcUDfutKbKjB4/X
QVXr0D2ipUWq2U5v5Q0lG2xxWB+eay+Eo+cHm1eMtWtWjTbwRHdKFhjEkRTeAklw
YgVm4dGHkA5Bg4a3bVK2SpxDRuF2PAT9eY34kCWj/0nUvgZnV/hjK6GXuOZ4ZQh8
cd49PoiVpRThMGuP7oSqy9bwtGfOo1ZlMNwdgwiO7ebdTo+fIy3cfSfibrN++D40
N+2MKlbu2A4CWDl82BNEa0Dd42+7+9VDZUk2Cjspv0XxKwBBwUTxEjASx+f8X3q6
N5al9RwQk2LEwsQ056TKK1auUHRmws38GR4HaI78U3MffqmZYoHuOdngbKpxT7SB
AHOXOCIwoiKIaWsXKbimNkWnxT/QksEtPZkE32blceklTi4O5Ud4vtuODkcL7u8l
rKfO3Q/qgA0h/hqhINJdifiZMYaml1FubTT/OwPy8uxIOTGVPGSp8JT5JEFOxwKT
cSd4HkwgT9qILsvvYSflVtIzES3HtcNltQPWQslcDTQ4hBXlbNZiKOhMrNMLefpO
noAuPTzFORpH6yHFde/oZ5VQuHja5TSeVESuQYyv/3Ync3AiXxpwIJdQJzrdrAie
C/Qm/fPY3LlZtKR0mTJ7HR+9V8GLMgCVXFyTjX5Jn0dvOsYI7XbRI/i9BHI4utGH
uOqM+gVBXmGv3ITBTdMQ+fbb8OcQP/daa6R/Yb/Hcls6xNw9I4B1qVMRi617yRDB
CewiqOprooTrrbZIAnTHtkaErODaRZGOBB/41ZehTKkmvxq9kpJOXpCnfiEHySRe
6twiHYZsmXOI8YQCk4+sjN+GPe8v9RwBfm+s3AKB4a7W5FPKDFGlQKP4d8RMLdu3
YAjLMUTqPgaJY5EVmf+g83oIC8WJIGOKJa6gxBbgskBKjb+AKsqcYdgHhLwONRqp
wEf1WgyvAkyWuSBkm48d6cfwAtmQFFbA/r35IqpbTuNDokPFxy+EAChEPUvPpnlp
Z0lXG7QIRmFGqeJNMGl44HeOxVUPVFKZxVmNcN826paygiaTTlrogp6SWfM1yj6m
D0HFjxuLrr8yNnZPNAAowgpkJdRlam2esY3aJ292B0dvtFtq7YH8qbkknuZr/1O2
sDtzDayxoGRZBzQXXjcbYi74rnLRQkhRgNSv86jpZa2yA0Ige/HcfGsanplRzzzs
ksEy2NsJF3/2gcn8PsrQC1iwRAxLDRua6JUPaVrVcLWKKolYW3tgh4aKt6jdNK/P
4tt7MTctUfQ90uH4cxYs9ogYMn5MGbja3EGVXxkVAfnw9TT5tt3JY6cjOkNb3b06
EXqn6pF/yBY5Xy2HWmg8Tk59TFBFG3c0/tmmPin8zFrfaYaS6vDj+Nv2Cxk4hwnF
e4Ar5iQt+tj+c7LmaeSlk4ItbxO5fD/Uss8aNfFOThXFxSImaIxf8Ek6Z9cADVB1
YRhnBeThAKFps47G7N1DF8Y75CvZvxKmfBkHw5j3MczgtY18bJ2Dtjq2cnIGQ0JA
8pIXIbTmKDmrS+febyHdXssokZkhJ11dK5JB0AH1l14ZOTl82pq6pJjmhNDxYILg
8iHZQ7F0w9iHgUy1pfBauKu9sR0mCRuuo68r8twGbjwtrnQ6nXJ7mInPwrGuVJBD
EBwqdkubWbtmiqzmrPSmgAs3Cgo1G8mqeczFJYyQ9hnVluoEidbfDt1z3hutqQaO
GJ8nhOSDSU0yz9MLUGRhq+LILHqn0ymW9D39R6LIFIySeqbfnqyF/xr4CVJ7GEAz
piF2h/az/PKgnwZLK87/MuINY/nap5bceiyvVdt9gz1WANhNVjmQrueNHvEhK15x
JHRswZWyWDesEs/9rzD0fuWNXgOMMk1440WPrcRHpOcB5estaf5jIz3xl7nNv5u2
Y/wHYOJ2VRUTuwwl3ze8ikXH/heXsRMzPxRY1WE10PLSfHmArMXgkwV66kiTQki/
xSPLMG+8sv/7L4XayrNr+vIp/KxvftUCTtsGqGr+zduoMuF6eyg6zGfm2AdfxbD4
WoZuvqAqXGXoPLKoyCUU3DXxl5xHrDxzqITei39ZjefBP/Ksb5t6XprrYYTavAj3
pdXd+a9sjv7v8EOqzFdqY01BGC/Io1EBR+h4wRGp9/xwN2Wb6oCmuC3rW4o4ru1r
ZJ+z+qSZ33CJh3rwrLRq2WhRdwLT038sY8YoH9ral5YEAVXnWvk06+uCtMyysEXj
dnAUQs3KNNLxpHbiOo2Y3BsTinYvkIku9D1ZW9Pl4GzfQVni+XVC9OAjAVIuP41G
oY/qE7blXZveNQgClPox3kea57Qaz+X9vP1x0lxF5Ps//OSRNGkAD4GFz3txywpO
HF1oH9tF/HHDy0hC0R0wJ7EhkpivG6Xl0xH71wFiPfqFUzz384yLGp5HnwrZ0K9t
22YH/cANcN+pavO7t8uuVkrU5FhnOYpWPJ/G1/iBNKTtL7HPIdJbLPB/1qVcdcVc
F+bswA+HqgFtCFtE7WADbt01veJshOgV4iVW/GQvpqO5Gy45wO+qSkB6kyvI6s2Y
Tx4f/z+BzVtl3lxXMET9j+Cpo1n2iOUa4M1uoUAPZHJDeyccqPYVMt2/ufoJ46hB
uG60WhP/FE6GE2PZYmi9nK32Sei5sM81QRT99wh+BdtaLjpcj6CzX7Hn/DSDru/e
OSZpzxpDhA/spDR6Q49UsvpOEXKW8iXradwcx14DO4JYQ2jpQt9W3Rc0CmooDzqh
LiT5fx5Hdyipzjz4vYYV+o5a84gSub/oNvpyWNb2WJFVGP1lLxcB+2q/XOoecxxe
lII3GnfrQbyakfcmKkZ6FtakyJq6FeYJ3wm13ayptB3DGqcX+gxbsDzO3yx9RqrG
FvD4nzzimMDY5QMv9H1MIx+2IelqKIJDJhyokdWhrFyNZa61OOD1TVjamnNEKW1v
zGgzKMLHqEHiRP6VMMpnV2HW0C4qpre0jq5jdaOuOJrTyXBoKb4ddns47yEkMD2B
SkFQoFPhukEvf1ranOSQDZR1UtXvKKx29X+LCBuTFHXxyiN86VZvU5qbC+IrNpVN
ajU1wfnXF5IhDGbijoVff4A2ObUR+gBtWFauwYgOBOEJ2s7+2KxkDck/PMW7rMs4
qr4RYljZJTf8aoouwIxnN8cDYhsWUCWivr9Y7L317MPcuQlij2u2yUsSQJ62UedL
vih3fMqpAecnwQ602HtFrnva1fpmbbPuR0vGrN0x+ZyEeDp5UYnQvmE7pcmx3A6Z
4Ilp4ZC/OGSTksk3I8nI8xQLc/ZB47AsRrrp+tGnZBRvr3S9war4AYu/vd2jlIeM
Crtr0KYWKgOP3NAG/YN8CPXPb1nq3P0UlcIyuN2E2uP/+qYb2bJWDn26U/MHTJJ2
0qbkn+dqHGnXp5YgUwTJ4GqQzYVAI7oRDD7e6xRe+aSKX4BNH18dd8nM3WfwKpTl
k3Eaa7gLh+1B91QagNO2LyAMugVDp/WL0/1wrKhQvmxG669BDfwOwyfOg3RGQlWx
n1IGBxgmaH83ZrPP26ZSRAWG5f9HJz45tbc4Ln68WpsRvwp+GLJgEV9TYF9InMXH
MGdX3w0E5iJnbrD8Ao1psdzzH/nWDe0kn1MiILuQq650zAVfbRV/8Uq18aAD1vrb
Io7z6t5nxjJ2nGzik9khrS1BZsWT+sL5/jloaPuAfIegjnZPIIdkEv1P8ovWZlDP
kxbAPtY8nZhTKn0pCgJnNOEDgZVHfOwxtLUfc7CW9qLwVcaHszSJyKHhORAFaapQ
YpNI/8OPYd+X9JRiTme/ovq2/LXBPJJ+3/xczzBfeyMwPgUgpKsPixO86S2mJp5T
4jVO42SZbTOENTM/6xFtLJJ0yUgK/Pem6fijzmsPquLm+ttp2KzeatmJs/mEVTMB
ZqLq153BIT4EO84G9+QjVvKXPMPH4kIDPwi2NeYSkwDImQ3r9ovgDrwevEvs/zTf
UddDVeVFISmYhK3T2eqf7G7d+brZqLxsJl1GHSzEu8IvcNdhol6mdjg3jXu6ZYt/
FLmSC8cnSFG0zkU/IUn6jXiSh5cnRYoIC1dEYE/wsMg9hVDRuUF79nf/ESqYTK1K
NgzbYnXVK61EUz+5rmbISnRdaEQKuEcRr1cCc9tP0X8qviUfvB3wS22h/nvO/L1L
bfknJvGH/ZT+j7UfIjodXmciqUlQakX+yWobctyk2LapyFNj/yAvWP2hfdzIdl1Y
0MgEqRqf9ZkdaFn6DanZFPvbDV0rBeXj2qY1acr8z6wjhgjbjHgvJxv4pTJjRRAM
HHWF823xAEBgzRpcPndlv/jdtPZym37Iuw0xI5LzcMmKldBfYbI4lfP+3zqsVIld
RPPj09ruPABY4c0oHa6c0SCzz7m1OjR1h2+3hcQWhRL3jlpAfNfByn+/zCk6VN8g
pLE6I75Sf5stWHBuWXLScg4sLrVAvQpFSL2TBLdFulQEp6TP2NiZRenH85io5y4c
EyeosuEwUIW+6cAbQl5e/LVk1nEJTj+8fHQ+omIocgig/JapnXJz/XmHgqF11A2L
ZZkRgn5tqF6g+f1qlPwwhOwakrPGBjj880reND5yPSM=
`pragma protect end_protected                  
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Su3eQyt11tMVkGYzLhzmHTcfr7CMCF8uq5iEt+KIgF00ZHp0YJe7X2XFgmygPq1f
cdyOi6wohjTmurmJyhodgAjYHl8tev86EX9K/D84kNOAhIdUjICEy8seQSzqGoPW
Bw/KoAkEiZ7XKHJJYlMJUZFAEeYZ3hs/FwbJxXaQ8oQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 110040    )
6G+jpLAN6yt2LVfZ/bcBMNmgf6+BNzNzgodkidQlGKJk0telEYoJM6t1IoDflKJz
6KM2QbrS4Iw4Yo9IlpexQxXsqwIy3YHnGE4Nju8wXxb5FC5xgmeplv8Dj9BFTFt5
hmczJRlDrKy/6iPDxo37YXVtEDTAusg9mXQIJv81at+FzHCiKLuXz5+49t+CSgSu
0nUbdkUfSv1sXFQoIlxhbz9EERe/HIq5FGt+tqpcaRahnOKx5tStZkl0pLBFmpqk
zIMFOddUT29nUxDRzk0ldTO1zDCiFEuYgIZNQ4Wq2sgJKcao71hw6cSbW72vYRRS
2WOLQIB6OC0BrxdmWlC64Rgjh+qPFY+VLKsXrUUbWy/1AwMxUb33hzFSdQHIVV0/
uGKwKfaxLgR0P0j297xY+A+5dJfjtw3Sk6r9I/ymQKES8XkezFRlDBj+uV1gd+BW
oeZNrhtoLLE1Y28VDuWB2/35eE9LvkEyZdcX76r7UFpke66fJCangkMpAjz1RBBE
omfpV0yUS1I3fJPgpvnCUsuIUUVw3frnjlzmsjVFTIT8tR6ZzxNZ1rR+YYhDPMq0
KSygiYjbhohlwidGaX2sCGzTqfsv4T1GHa1zXRpxd3r72OG5L6CDyGkbAKf48Pew
njdlXNIrO9MgXL3r9GRwApKd1zWZv0E8QcHIzQVsq9Yo2NR1jX0AMn2adm56GXM7
JGFo5wyBd6SVTFM5R5RN679s3B9LUPQ/flS72CEGkwGyt1DRj6i71E7TcSfGkLze
BXsE7Z3b7YFfE4JhwaWEKg==
`pragma protect end_protected                  
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
dLo7FTPJsW/sTRZPUmBNCN5cRxZikSBscwJ9zl7ii85GQ16Hq3Zvg5pqQ+II2sYW
rloD8bYGVfET5K9llBakV3FSzlXefBSig5oYaOtCXN3dQr/TD5rAaIlQLaIYaq24
UssLTKp7vaV/seO6QyV7GXHQEu/LYf8FMcSoZe2u+0s=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 171534    )
egVD14x9hB93/P1+7qhSTA4YWihHhL2azUX/WUQjtHhYC5lTXX7dqDfD7wki9MDa
Qm+WMAaZ+9sM1Ci98S++fAYy41AtEkHQAvleQqD7UtwthHav42TXRIAZ+xHApL2v
WU4zNy/V42T9fn/2+khYH7EqVMNxaqQOYrEhZsuZDWn9K4/jkQKCoUY31b0OkIax
re+rQMwO2GHtiQptrpE7R50+Jw83x2WBzTl72z5w5jLMw6uenFJUlQX16o5D7+Mz
x8NBFdhJmlScQDcutQRkRPkl6fvf3QXPYawepl/d5HYIK/r6Mc8X1baX6Ai2bfpl
BAoc2Fq1Jt6cjGDi1gWidPg+6Oz1irMKhIfP6q/C9k+E0KLBJ0FFszxhQIGZkcL3
ms2d3tDwCi/R5tc4p4FawAYQQVrSEXGXjhlQZSqp7snUg/fXP7C8H+1JPPLt0wZr
189jh63BwN4P+wXkM4tjbskAtMdHlfj5M4UdChfupnXJ86hYu9cFqymI0r603yAF
YX+UOGoAOYTw58T1YE/jtKnqcSJ2VbDSDFRLcqPvwXv6LhCWr0jDnMuVZDkB0EcS
ZrBXPumonCdjnBe32Q4IMKH4nD++Dm0fUddBSWHxbco/4pHGb8ks+IL6R+PGaRPf
MA2/7mY4+ql8IvXW/IYWblIGxj4UdofBBOpgyVUgca+TU52+HZ5SJEFgEq6+j1Q4
dW6RKP/xOlanwzFiQbj29Pa14BW7wnVXM1XlEbjEnNfZPpR5GBnv8sVRec/REL8G
fEjie87x834JMaukCRP7GsM73LtadwrJ9GX17IxQ7DYULxT785XIBUK1jQZSQkSn
P6/Ft4o+Wysk3xDLm7hAtCdJSoi6bIrybyVdG01bU77DAG3XxcHhoVznR4h1uTwo
nI9EWLH33r3rI/0KLMpEGQ1sXRf1l3Zz/iJuex7wh6kysJPvv4XqMmIVISJPMihx
Mz5mcm1A3atB7yeoX0e5E7uIUvQvCYTnQQSNSLE9jAWThe5pEy7NM9thh2hTN8eb
zy50GIeDucMwuw7zrw98Q4K6Rl40DHmrfWUrzbA6PehzpabUmx29c7sqd/CJl5Lr
LAY6wrIq64ASKISXaeYSLztA6e2UvF3O/3hH+OcOc1tQ0HPFN+Zfy4gILPpj/azm
hT0LvFhewLiGERXHztuSAwWwqklY1ERoXCNyJAZ6sbzVkTrEPOR87Tnyodki30bj
d1e1eCp2njIGGIUDjW65FshQO6kpUy3vXPdTxesHkLbExJeFWSX0qibzJkN4Rl5a
z0J8ZvUXmaeld3/29OxC4HxnWYjoqX+6w4BpbUCc8h+Rpt3B+C718XWnA+GWLxBt
aec7CP2GVIe9URtwdWFwUaH5N9h8+df5xojbbs3Lu+rpAAYnkxQWnDbsEPuCAjbd
FZML+wiFS6z+WEtU60uNc9DuwjZvagPWbrasLTBaAmgoM77uMaHmH5Cs/2DtaXPM
4K0uJ4b89dJ78DA2F+Ub3Zaq5Iy6DQSnkA4AZCMiLUQZCOfM1plVemhCXYK7jwF+
2yQI8g2Qp5kziG4cODkqhTkOlIF7T52ty6kL4ZDbkQ1LkR9kbTq4gskxhYuao7Uo
hPITs23oCskmzogT2HcT9a+CmVJqF+P9p8cjXxtOT32TAFqLC8qpfvbJ9N2Bi8Fh
hV8v8nJ/EvYO1a7JyJf7CldfQVv7Np395+47TwietCKd58gan6wI4pLf2nCBVAtz
uxOxzSvUAhFQSVWvTJ8w1o7xVKdYtfjClAt+UU/w79UkhcNSjqoNauNEXsT2nLRH
PNydWoE/vOPARwbZdyq96das8zLw6Cgr5MqFLBIfEorXxN9Z5PKX7S5XdL9BNGMM
JwJFd1Kg1wmXcgX626caPgRhGQZ+2ipwxxV2jawBXwa9DP2Fh/09Tc8xhT+OCvJM
qRXDyMEaOljm4DOSCV2z4yaKghZi7OcVn+tA6cPB7YcN2vUKC1vXb5MoNwKLfTny
c74M9lzUQx9KubBP/kScvw8olmKbWkRvKjSND0r3BtYcv4n+KhLr9E5gge2jDxPZ
bMioFjZ1hqd7FR/2iV+b15EJYjoxAr4rBCQCFktwMep4zXDuTnwWYq7bslaAW0Dq
cjWzHUrGbZR852vF4rF++th1JbqobzDuxN4Qpno1NQNeY1q7HeoTKd6Uh8GvYqsz
FutuOp8hNpsZTdXWMMBEdbi+F7+ITE3kHRjVnf98k4SoE0ci0uuRECGQEzeIPPqe
AJRPxxWcuiBtZmmP4CTkQ3NGQhL/sFPHIEqqWrDRhqZwpKTThkZaIE3VMvNxKmCN
eqoa1BAh/5+JPHfoRlaNAMPgJ9HcipnliRZ5xNVGbSNNWra4XCjKsgfPs/x6JCKg
H+6L78uoTuXFA7rvQzqPpsNU29cxgM6PeyHTSHdjz/KmuOp37ZJQA+h9anlm0Ff+
b3TQxbIOChQIGcYiAPAotLloZqf0/JYD/e8k9g/luMRq2qAZ9oG+r04CeG8T7B69
j9tcoG6dqBsw6+xm2bmTDvpLELRBqXjiNcEIUKPHolsMBwQg7Jkf4RH1NZWfHcHV
0+8MGIYQcWAk7f+TKLeSBQytoPSz9jFFpfe/GDC4fMfzSM+tgBNJmXxMpR7ZLFAj
IbYl+vWj1XnhB6HVswLSTdhaUgfed0qu2uwyKBNYro8/m/2q61wxAD/CTJzJ/L5W
Kw+dV3H2NLZLfNNBhrdFO83yuyoiaaq9OoKZSMq/T9hnxYMCWaTnITQTSgUeuDKE
+/fuPPT3eQZEj/zT23jKUZvlRxjA75A07wT2aaQoTJQd1gtHnci4bueOkBuocsm7
VlxjsJ4m88cnS65d+w7TdVbQ8VGMTaSuFjCxjkyZgsVF25WPx6JGOOsGCWyoncU5
tsnYPA9PEsa+jmjsrIEHJwHAaJ5p3t+0FM+hj1vcNrSC6WdnqXaYVI+GkRc/Aoa2
Um3X3XIVjs24C7KZmhxJujZI5WXAp2CalQtFxg9vq6msHh5gv8LiukCrK6gz4TfW
VghXriX9rlrJ0c+5VGDqwsv5T8PN2r2GDCN2jDeYkRVAKFIQAIBLDjkQqGx1LCve
AlR21jW93uTDN4H0UdXavNFPxLD3Jh+IuNBDCVRrz2AFpmhemogVtarMWzQaNc1p
e1f3rZPPr7ng69VP9Nq63Z2Sv6O9csM0498qEcPZ/rXgGY822f6sUZ5IvV0tg91b
4YZvdnKMDG6wIVU2EAlpx3XxKyz0teXMUeSdCXHvFhKLyvaU9Wx3gp2cdDdPjrHv
4SesMTLA2liAR0wGRn0Nqiv9hPJRydxdk8IEjm5R61zQGgq10YiUb4MuDbneZx4c
d8iiPPGrd8SGm50BERml30+GTQT1OWaQcjMgzwqieJqM0/PJ0m4KbFKBNyNXUTZC
SMmcS+5lgy4mT6SkuUcyBDnI8z7tskPsd3S0Xbg0EbnjtpsWu33G3gIP1dKPHdUb
mD3Sj+FxNHHwoACRxMUKIYeKMiDQVQom7iO5FZQkl7iiYSVYMiMXPWwJY1RcfND8
I1nOCW+NjvF2XJkx2+5oY/YIGVTyLJumZGvp2GerBnfldUI66XcPxwKcuc1uxDzg
VpFIaGOZ0CVwSVglQHIJULc6J5XtJRSYOT1gUzODrixU3NBEFK5n0dF0GdGNqe6s
+Uz1tIVCwv4wvx1h+B+xe9gGYhTSJ6nXUZVPbwsK8qcHmfNKBjRiElZ60o97gQnr
Zr+Mr7OPEixbwgOmkezNTKntqLopXLoCPO6hXm004j7Jr7JUtnIRtTTvdzjBXg/V
Ny59zeB9RCPEB0ndKIfiqc9Ze02CWO8sOxTOyXD9DqwCAhXuIo6yq/JCuriipr25
GH7NA6kqIRiRD2j9dFHQ3gnsPtONz++xHVkbYFlHmmNHvKGxKXtsAKDgDNufWSBz
0lT80OU7T2hyngDkxMpg2Ao/ZTe+Xbc8KQk5+PG2FdXI8XrI+EJlxCKFI16Cs5cq
dY/0H7pxlTJBUo6d7GYQqBk2ymj8LjlZZSbj518rbm1j+Ix75QaN7vViORxwe0J8
OwFBSTrrHWmB8WcjqGp/Hs8+WmWJzX3BOGUQxd14SvFzgjBvIlfLbYuvm1TGrxn/
0DV1V4Q2XbiBfDi4sjhzpqRegQsVNiDXk9q1dmg083ptR01SVXsVPqVJNWrVuTm8
ThCf+33ALMv9hpwG/tWHA/ZJamxPvpRJn56Iv9aZY7BRxo9dLqXM0hZXyCXFm3u/
uYBovktb1DR5Aztks4BP8V16Xtxukm8UihtfTIYUCrUhcRZOwWzjSaNa99QPqzFa
Na1Hw8wHpMY03aumq/TNj9aMXPAy+20ZHjNdlNlrXlWSni3UfB3GmMe+XNEtmU4M
1L3h15Sk/OIXf4B2OLRyksLFsaC/2ubxPShuEjTWaemLHW0tlvcYFKuXMeuaklPX
ihlQ0FldQ9q9X0QbYRkjhVvLUAw+rBP3SqBTbC89CfxAARfstTVnuu/3QKfm7lDr
6/i8P//4urX+UJGqOOo+B89TktMBL9aMPWuUlEYoAwbJeRiVP3jUqG4QLv5lBh8X
vIb2pRIUv3qsHltg8zxGFGVs/7fTTSdqlbI6XZja60YDsF3XakBabvrvriZkw9NJ
3ib+FX0n8rWeeV61iRxHVyLy2kmyoAq8vqWaw/8W14445/bWegw2/WRj20PSLJDV
kiUtX02DWJppv9/XkC7Oc1ot3FG1r01UlP+TnKNgQUPGYqwfktEGMXHHKziu0nG8
bi9cElwbAQ2/vycr9DpovFvHIe/r8FJpyPHfDO8IcJxmCeT+XOQVuClZ6bS98A25
hZwBOn4iIn5RfmISYv9XF+MMpQluM0kAs/otej/C65mQObn39L6X8zZZjojfREVb
xelZYBnDLdiAv/dfFbxvX0273Ux0geMz4o/F4XyAZKUhahusECO+sem2k7YpBJ1f
dHkkcvr/MCurirb7HKWryDS/kQmi423AzMZJ2tcHsIrXGlbKkNcnDFfJXuMH9nyz
q+8ct/+TMXXJrGSKc8an7afNzugOFIMwUB+B7vkJddQ5M8IDssegsXluvcgIbpgb
H1pEq4V6NpsopbnPj0ApbGXo2FVlgWYyFR7A7aPfBFyPzeY4Wbp3c+Wu73scrxUN
iCQEWhGov+6+JAQhExDX6hRyXwl0VousOhhncTxnDo2r/K2FtqueYbJKG6AdqZEB
i4kwLs4QYSQPlr4+hYOyqr7l3OyISsbPTKwoUxU+G0+UZfix9zkxMtZL4GM7ZQD3
rCAbwLCt7gFs6ASA5SDa+BKHtx2CveXvtRlbCXf2ELYPqcgGJOISR2yQU+InodQY
ruG9X0rw2wSvdqZmsaXO4l8gYDaX8yL6mr4EJzudyaA6LNnJouJeXZiKpYHTGj0Y
ISDAPI9BR3kKLitQ70XtNGpVqKN2nwNDgg7JpHT/8tdEL6p+ZW4scj4Xg+U9BXv0
/Qz78WDukI5yKmJqiHnO1Z+pk6opkOcYVrUH2UD9nlI539DDTc2Y9iZcgMZQj7Ko
mwz0TN5Y00+hf1lzuQCb89Yz5ifSqqSGLThAGvG2QWmg5asX/zZVOP3h5uC2WdN7
p5sJlNR2fUKTzaYhVILjb9BjWZo08TYBmi2DcYo/zeDAP9TRcQAqF5CXpMfvtl+C
rMZMTk38FMuVEMN79DfzedKB2J6Nb5rdsKHzrZZdms48BenM2+dUpjaZm2fG7BVu
+Fl0mcZ8riZXPrIS8txpWz26ybeB98PGdB0anauenoDnUzaessTdEPjZYdfRoa19
i0sCBpcVIfoKvUnlWbQbonDMFieuWgzOHZBG0JRzcVvTgLvt39Y8OmmgKMklnnH5
wo4OWQFJex3BZbWEXRLDQ8Yx05phHwdyMGcdWDiquOZQfe1wsAQWdmDYyfbk8BqE
00zTLk1j+vOarXWcSgVNsm5W6flHYfoSs/eiPFr+hKdWjomiK8SYdUXI65Vd+ieV
PVXeENqDX3MZR65APmGyOT/20QJF8TSF6eqTIzn2zV0//KznHFaAIe4LL2O6bHXp
PHDD9Oz1XX8i69U+dkXRdqUiDZtHApOayKDRpFkAM80NE/1C4j/y6cvyBljlebu6
g63utO89HR60x030XvThdS+9Mc709nfgXvBnSzBV5gk/MdLdVbJsIWtsQQqx5IZY
inC8LS+TQE8HT9TuLJlR088L231Wc/Vrh9kmhdrL6WHLdPuOJYvOUpE1T+oSLQ+K
fcnMzsIEDZJhIQ5/9NqtaEqZEAh/b2fO3vHmLhuIuYunI5k/Pb+T4TrTj2ZN1tqp
AaFyDWRVGg7peSXnzQsTwk7P15XVWgqWroaoJ8VwPt2d33mpwCDosWOFONbXjDYG
OUAbkWZeO/o0bxymMtFaXh938YcYvEHnhAYLjR/ckeeuEL57SI4r8EhjAopdhoYz
92FDVYRhb9KJYIcbojQFYhjweDO7sptpELiD34dLhsa28EonE5VQIXCwwXxvkW1x
KGn8aDMQzmzYgl92vcf/aNHnlnoRWwBsKyxyItN22qomFqDVNYoG7f8HDO9g0Df5
FO+pUP9a+YB+kHiTahIn5r5+fkX1WrWBr8Q/a5wy+oB3V0bQTO2YB8yAPwvzMUXJ
1UoLmWmXwumCC2roIQjUOO9z7VpBYnuto4fcY7D1wxy0KwJHdRjm3zq7lwsEtwMI
xWtj3NA0+qeq5iASiYQK6lCe/mZh5BiIxPbZNJVTtO/3j3A3O/W5TtHIbno3yS2t
THl61UzQTD42Y+7aSXpVNgnD7cUTkRhEwpEJ4AWZkfDzNqUAS/kwG969JRSYNNxY
sYm2lMkUYBa0NsiHgEis4YE72se2YBqDw7ByN2EZra2eebkHoGy6a7j+n+uGdGQN
Vno8Fb4vwzczPVAvSN6kXTCSJks+l68tTEqP3L3aXyOz9QGGNM/wopO0VOg7r1g3
cQCQHnJJthPKhWfL9RI4hyAp2lMtyW8m8o3af9U+RSgsnoZ6IAPM0WZG8zkq/2Fj
9j5z4MWZqdBkZ4JATKryHE9uP0z+JXSCsKxpG9enM2ae2TsgxJhrXutZHpcA5xn/
tZOMXHNvYvkge5TDHREGoYYUW/S50gYnXCyOJfyj5GsvT6fV5y2PQub7JoZDkn6D
vpAfJlutYrI9u9rF8VZX9VA/Zznl98kj63luUUbVMl13mPOB4C40pol50Ym7tUXe
0KwyIOLCHOd07TDmix5dMxTbVDp0QjlnBjh0qUZye868JZojEqAiQEkj3aW3sxQw
bfS4+ey/sIBPqrGqqOGuXZXPtjnj5uBinen7FYHes7bj9KBJFnPcXz8pAUWHXf0o
SlMuxm6raS3kxxUFwqtNRVUPpccKXoojWUDrqn8cCrzQSSjKIvt+SLcyWyDj2nq+
LT6ggCUTcmmp2M2S5Q/nLPj746mpUw+bqiHTsF6osn3SpxprOVIrsh9PbiCOoM04
gyVOVtTG2XUP0mesHVM3jJaDJnHlbdB4WUbG+2kvP94lmC4nhXI67qZpX6IHXN6h
7kwFdUHcekYFgbkhwxhANY8dfexmaOXLxbrz9puh7dyZaCxutUpBKbu9LWvP7t8z
1KEkL+Pz0c9E5bcVOdCwEGTjNllb7sc1J1YQW73J/U0iwlD6M7vBubLbQEo1gJ8L
tEtkrI28gjFZZEEC92dRskAYVAIv9PWzaSz+oyheWS5qtA5hhMm5l7WckT/6vjoN
oJeIMcAtW0PPZKKhCkbs5ucDoEl3dMLpzeP2s/LEGNCKXGLHwm3t83u2uY3SBEmY
j546tNzfswTz8QDRD6y07bQZ5aicPfHJCS884e2dvr3sHtm3gnuKZ32a5CTc1ntD
U9IvPUB6fmQ8NwEwvfIp6AT1cfWyJ4viUAxnebLJr5lhfQ5Ja4ARHTGBxNWMaXyP
dJON07TfZkHqqhHkv6F8hwCavQll5nS2GPsDfrVS+cM2fj/dKezqxubFJycsHKLo
9tCFE5Xhvk0dbKSw5VLuu+xLCP0oGnV3ktkr3Jr4G9FYWeRnO7Fe6gbjeB3JdrZG
5wknaZpAnlOZ8KIiAuV2V7haOrsl1PSJ8A+FD6zUCXtNtVtIJG0OBFmv5z+SGf8j
pm+5tqAw5fXIxgwh9BK+T95+uHCIROW0oJVVmdsrDQY8sfAuIGKGRCi5r4/nlXnj
iUoP7Q4pCupfpIqz0O00EncnL6rXWMh1rhPAscwSjvDMqyn11R77kOiIzAjW73ES
ruYdFWghg1HHNn0cPWldYOdAzAp5174F61jQUW0QxDMWlh+xw/s4FGTB6Rn2Llkv
Swwa0+d2mNYeiM2AW1i5mer6BcPBJNBQspxTeHZxqu3zySyEiIG/snanjBSpEmLK
IzdleLxIYdvoM+H36lN1bOpGNeY6rN9zq4h816cY9TtVTVtK4bwtRTifpdatnDGg
bV3/jJ5SMQ4TK3IZ65/hbCzoWCgr488t1S2eW3so6ZwO+NxDa58QLKeLMb54o11N
imXeBwMQ5gNfWA0BUqpKsO89lDiF8snmnIwublQO388HotBACj9bH0mCjm8gT4hz
ouPo0enSLV9FRJeYGW4vMgmCCKroFXRGKPGMIDIu5rkg7OywbUl9YtFkRRM1NCMh
rYeqeECyLUfzKA3Irz3eiPDNr4hqtGaItAheu07Xkg/L//F6LDJHaz4pMoObn1oy
egYwbvtjfQIf5zN0LFyVUp/3bKiB+xpKA5D9TfKtJ5sADzgY2ZYqXWFl8wJFnSwQ
dar36a0moJFemGsrcUvoWFqkU+rHD3GtrcK6WzIovxTpYJ6j16/l7RcOVpCPhams
u5JG3C7aXBi17Nzcyea3JOhag6u9T83j4MmXcOxxcdqhzk5XdL4xTaisOarSKdvg
eP9xv2ZsNdh6KFAM/cvjfToADyM3T635lO2kQDd3s7Nx8WmKp4UDh4kAvHhCfZ/V
Y4mvn0UmsaS32aUHWjctovoX8tULiBq8rICPIyUs5mN+gRmL72ZQhonmTHZAdqNe
aehO2F2IV0N8WNy3CHziJzlJhpOAwoMj/BNNOW2JgLk7VOWZtdIywyas6QaVJnFt
yHSuJvyIE6MEaOfRjGRGqW/Tli5G8iH9gdnP1OAi4ZF1S8cE3TImAUEXnJOsF/4P
nswvcvjOHO2fjyWzrJr2XMz4941AW8miuiNUMeCDDf1Hxibkr3SUtXSTA6kfNXZn
QQY+8l1NGWKb8KGP9LyqUNkY7vb/+T4rrXCthipax+ke3efmdDvYnot9/nN2t09r
rBCgVAW/AfVlhRnknxmyJVENZt3L61Sz6EyPH31rM2k1jI+rm0hJqFDxlwrHLmHl
Vh54bIN8oANqOerZrWpcvCxa1hfV5vDoU5d3HbxsPkeEQCu6VaNW024+Ms1otIyl
m3p+dXLQuE1PLb1Xw8KRJbJ94B5dYQwcJVkYQDFXFXtnXozpVi5o25IZi34N5qlq
T8GVGvcAAYa0eo4IIyIrfiI9Bkhxfv+LQSlPA4cgnYL72ZhU9uzAFpN9lGQcEDoJ
8CNDFn0hR53H3mSN+fo2E8ZeLvIuQ5Eie9GhDP58v8Sx0WUqMjeca/PsXi8IiaHn
lOmT2byFwq7NnoRVWQtZwUo0DrkDRlto79PXkrEwoX32i346lozECHzK81I0CtqL
61HquE4uMFUJcEEAZ8RRdxU7PG6F/s3/YL1EwwA5sdNv5nv/cmeEc2/qaG8PaQng
hgI4+dXwhcVyskhqmHfWCZVdD86pE/ydsguT4HOUX1oAJ+mZG15U6W49v4Gd7mSs
EnULAdOxP+AdL1rf+0IvwB9bb9PIz8uHODqjPfan80E9i2jMHMERgdF96kOrH7Aw
akHYIhZVaRwG5eauaFNoPcnN3JphH2w4wAji/h+rVIJi6nw3GJxdS28s2gAdFp11
sL+Nk744icTVQkNhKyTL/Lw5vLCMez1jwR3+gYyxyIw1WBFefeaY70UeggevGJZt
2a21QAzmoJERAQy17jKW2kXwY9lQZV35fZ0BR9i377VkePXAB5NqldeBwcxiy0jW
Xm8WWvlpbfFT/Hb7AWA4GiLFWdvJB/kbn+R6kW2xKP56Uv4VS0PWjQ13W0RVLIqp
XFAgh2+B6IVkeK3z1urUHvN1B1aDhXcI7orIWglDwapgXS9b5WO/6XokLaUq0pTF
eUlueqJGQCARAm6oxrkSTWpg4OASaCvsd78WN99CJHb1xIlTTdTZe7uTCNBNbi+v
mPHXqi2bOaRpM+iK+Qhh+FzeNsn1s3rynGYowHbInbHM4uhXcXcCzyL8rB5HQvvU
xzswTk0xPTiZWkGGOs1Hsv/CM2yBXfjuHzEk5kbIZPSlt5mssga9Qeb63qWInAa/
tuSnUiA317Oa4ZDZh/Bdf79R1sexnBSvNOqhXU66Wick7tbHKoWjzmUNINnDb4+Z
xABqMCemMFKRIjNljyuO88KgW24Hg4d5vE3uXJ9RVXgcNdz8G3yjPOYf/WQXqjOO
SGNjE1qtHZAvABTV97sLHY4AeRs2PIfEy4oYv/Xp7plsrcbuIEkYHKkphA9gbrea
+eFZngfVhks8OYPrINiO/+0RP5YnO8IsenBblNWYT31hV4Lb3qXQzbEJSf8eCrev
mP9qtLwY3xHd0FTDU0U7UKrWMSUOAEhKX8xgvgrsAXSJ82fcm70sopA23szUe3Jx
w4fG7CCcSLJHCkgskitHzzhcTkRLiAUbyhSAjBfYwejq9vlNXgYgoxWwZmY7S88Y
UZZco22VyQk37Xm6jarc7ZvRAT2DyEC5i/s+MGXLgBR+s7UIK5TQgvFtDLX5XDsU
ajiHh+qD2idau0czSz1b+Dij0Z+hF2FkAnqHelrxcDzQWKB8MsSYvjLgmQNiokgj
2vC7z7EzL+YvN39Dz4I9WgX2/fKaF1+WI4R6s5dT19ALrMHKTf8FhIj1GfkGNQZo
p4s2E3GqZ6ZD30/Pb+CX33Hsl90b0Kb8CKbWUOjLM/Z48FCwxvp8vikZBOiy/UCC
TqmTkkulZ/eD8REaJpnpOuuJqQOcCIikAATuQRKF0GHg37kVRm65pNov/yo8A6jV
nVF04IPFbkfAB4HkpLn0EHf85EHHREbfbIL5DrSKX/IiXVYmUWx+I/l6kqA/rjKE
fB1kQZdNIsQHDCt3898WPChwBPgourUaLhHLmH+Z3alcFIJ+7y4j6XWVIYvm66kR
FUuMbzB97/dF5T5dTzHYPMEheQ3GEykQMpFlQPiJbTNc4ZpxSDKSYEj5WDSUvED5
XMM9XPEn3DREbUM9Fb/AmQXYQINQQnNtuHbKySMZ5qxy4uUnFtdzmcBwuasrKPhM
S6vZJsRO4PIwKhqFmjcIpL5oSfl2p1ksgMgteBsWoxyhQWR+zjJYhX6JzJdwS00H
S8MnKEiIYKp43piYtosUsIAcosX7B0neS1Ms0XkwblcVJAwayJhBDbQ89Apv4az2
H2owifFMkndLcIZ1E1GkFKUXUyVg1lQ1cBHgJw4kUoL7wDJcdzkklJRSfJLLeoPT
3J+jfv9xHrPFuPGkq/2qmfhq5wOTbkMpJqYgLDsU92ybBODm3dtQagnsV88DazPG
AIdA5r7hMu8cybd5EsykNh3qZ3tFA5ud6PQmcccsmWJvYux8hn/UdJocN+DqpwAi
B8leiozivaMG1xFk60/f58xZFsTXAVYI2/GB+LDR4krGsK5liDdb6V3hoSx3YEwv
b5y/7yUsqvn6otTtklRzUhA7yXrYNMajBOsie+LsUQ8/jiX016looMKLmYGHN12j
cvZomjtyNcUMNPDGfnIkChBekRrGaV0SShYY5ihDatC0kgoWWl4EMldhjsh5yN06
zkDO17CW53TWENk1BuM0UMZTH1MQUuoLKyjPx235ZPSh9DOrWojQMiIypLAm4FeD
HRw4f/rsAIrpDvP4eIgXq84ibcLvQ1RZXjBjbBen97jx2aePa1Z0EIgmdjWdRYNG
xr3Wum4AMQuH7CjYvlYLN/WZWpC3k6fHNvp36ug50pMEwWROVQVH5fZraRntpTmt
CPH8yJTks/YoZqHUdajz15QXULmJDMK9OnIrmTX23Q1vruOf+SIjJuDwXrkjAC6h
RS0R2Q2r2Otb9a8CB2BlgH/bVdrtyktdyy793wfyLRhmhQ8+NoarwPJPPCDPBZvm
hn0HNv8IvUR3xJpqXBj02QxUz0dcjCYvz6kq7VlmPEKgA5bRbrFAobiW1+V+/9lu
+PS8RnOAMWD1zL8kz6emL8O/rj3ncsSjzBwEOQbEOkTskj2VmOCH9QgxvAarizam
QAQjGXLUxtWUpjCInlctB+dpvxl02BF77MD2EU/DVQJW1U2huOxBaWScJETuL0/X
2xZiz0+aqssGggTy+YeySRZcFjrRq6ha6WYlmUVZMJy/sJNGUfR90Af+FQ/7PE08
xgRHwFnpsW4iZJ0sZtrpqgTjNfuJIiQUdqRWOjfC6jTGqPhLhivYGHiYsVkcvUcR
sTMlvWIAzhMYCIQ4UV/kfVT8pUKtmmK8fouuyOQLRtBl9gseaHRxDoaMQj5IxSUo
F4EB27Pmnkk3Tm6i5IsTFG9whK9y+c3sWAiwslwvdlD8uNKfEFDyJfZqKwBokSUw
V+LOGNptfLIJPMNUKzUYuwzpUPSTyYXCvK8hkMXGQkQzUZMR5sshE1pePaKhbs7n
/omWzZV8cRVbsIRPuAqavqf4q+9ih2BGNHpEqDCSGOqwvq99761zaysBAbRjagFX
8r9Nn22RmrLgBfxur8rMME134/m+0lYwbz1YDRxSxzdwmk7xcftUq6wdO+rMeHKD
dGRVTWin732LPFn3Oe7dDFfo+nsFv1fPRUQ19Qf/vm0GuWL5YfFXPcDpxzxWP3Vx
6OGWAC8bimCw5MsqRphHkSmhFJPbYJ9jzwDcteyOSMRX5sWP8y4elRCrWoTKrKa/
C855TMPFgA6wULRkYaxZYEDImJOApR0n1/eeQGOXKgadi4FPgRMFRlG0U5Ps3Dts
nAtKR1vZUnbEb+C2b8MtJuQBNdpLVhjAjvnVtEBpWxevKl+50ksl8ZGPRdXUv97L
qkmF68qseQ7l6y1RQwQ1tULdWtpaD9HsyW3AEz7ZCwum/oTy+H6FE9sakRw3crhT
43j273fVbHJsgvNSyFIGjRzBnl4/LVW5D3JQi9iaDBo3toVeac4ojm8svL8E6Bp1
5Ttqnn8JT7Wg9/MUT3KnBE6LO/9xjGi37POuSpdS/+ijcipUs3P8DhC6hGlZt0gP
8a8c97gRUyVFCnJazta0fRXQzKyTlLrygG8tFvPZ/g8IhhPh2TOJJEFd2uDRzHb+
q9UMpLFyCB6tQr5qE38iR3+Aq4NWItHhOK9coSQNHvrxFxvhWEHmcG7DxLKi1EbG
yfQZwDiTEjSZbYRZe+Kv1hm8AlYPECBGxGPc0U8N7O+ywP5F6pLlZmHwaazfKvbp
RsFqhMpJX5h0l13lwLEIMBrGt69uAreGV1EwtF5zNWm2IHzemyjaTAKB+nHI4N+0
fG+YiuxW+YeWZrXRk8HF4MtZ4RI1I38hZIAGoEz3lqLDkYYTz5Ir/0r3D8zLrLva
yNwQM/PoO22LXZsPVtMge8XMtRF612MlD6Zo1La7p5Snv96CJ/nTmIPkFGqaFhGi
vXL7yzVqSEMb5lCtFsvTvrsgRY0MeiaFaa739fS+iM35O6jKgwrQsXWpd/ddbidZ
5kpM8L8NZjZkBDv5XfO/+aLbae2KqCgD7idaqXI38TeY6a7C6WXQFryBHl5wX8EZ
ANq6bDNfdpO7GPOvBU1NAW1m9/Gb4+3nJT/gTbesCrAKoFmzUb1EJTRDK4C57alZ
4XcjFrTqmOKIHCEfFJsHwiKmA8fnC/2sjZiTPLoZKrUQTc/2/Cira9ev5HFPWm86
srFUZHrUmOXBZCkcV4wJ0PuBCPOzRczViKnqKhfXwe1Y1w9fCyFvRXyScqipVb4s
V5iAioSCBIXEcAS7/LuqLL6EnNSsqc782/g+LDZrJOjZLN16cEoD7eyPqXBUl783
+X67sQ1XQgdr5NESmWAl89qiAiKZCVHqk37c2tSRsTVu0CvcHdjPTBXejzcnbDdZ
DIO3W205SxzavdwCSty0Nb7CEHEDpRf4gyLmfcl3ahyG9ixWtc2QJD/rx09UC7tl
CXy0xZ3tN2ewHhkQNMqLTWosnhQBp/I/MMLUHXRzK6pWMuEPm8LDHIFWSU5za37m
6FLlpZ4lEnaLKFgJhfJkXDqE1D6QB7ogHjQYkekGgJRzpngLSqM9qZV1Z4vxi+ov
nb5K2+frJOoqKU6k2vb3rieU4Vg02oPFm3vUgetI86QVxmLiDbNbWZ9tt1JnsAF8
sUV4LleojD/tHmhWoDI8qWlINiYuGqR35Dn8W79/72IRa0Zk1bi1gedzqcdIrGgD
IJ5HUESgJHJNYNQn0V1f7tPTqIh+mTMn49MgR01hERk+VGTwmv975x7nHCM3fnYa
9ADSCFKPqOKLksAHQzuKiHDoGVh6yjkwqnSB4QdojXK1iEUyHs7dFp5nwWqYSIin
//zMycm0Z8EISV1LaMCt+48vz/oYLzOviWSbBCw8y6EU7XGLvxtCIsM02d4adITm
HjoNKCvmVhKBXpSdO9uNKXBcib/4oj7uhPxctcqM0LnfwWx2BByxGxH1qZ83jl7b
LUzJAPQ93hqZGj9K1S3y6cFv4ZKM3OU7biNEPN+IyuATGDGYmuhBLAaXlwwAjLkD
bRCFW2MuKV7l0z+Gde2e7D2BmPKkyZGSULPIA4IChZrF0G53HZcga27F7YAFKNXI
tXr7/jG+BoDuHpwUY4EqL6QuI+0awpgYeFwFwUV9z00/+9gN+XjDGVJ2JIFxw4Eu
D5n2D/FD8Sgx2SJG4SE+p9/zbytNPnVgMcx+NUyfb/+HWcNR/PbpZj1S08MqC5DD
X8NeDaHMXWIANfNX4edoF2W4wDJqyIwdwTQAq9crbjGjd/4GKoCbfpN3T6hJHdUz
0ffA9AKLlIt2VhUIIRB+qEWbIoRNZlH5wuwasPjwyqYVLTuAL0g6tSEJxMzddpss
Oz5SKZy1iJ2/nXCJZeFRrrCkJ0CcWdmAVwL1aFVB8oR37KbNZuhWzZVE9+KA0rAr
HlHy6FkhUuDzrH+dX4BntsZ9eCOTs7Lo86OOANLwIYaBN/AAVR8d5ToUMdgVflGK
mv/fAU5Ggw+fcpC8UtFs5IydREIgJ+lAeJCvOf7IeSxMDatXLWMRCu5+IJRSIZPf
iHiFOh8/zxsn7Ebp9NujmdJtkCO8TC5RHMZNNAf2Egmou0cCm89nhVQ3YOy+/cYd
1hCHsfsFViioEHdmUejmClO1t4lN9AY/T2tifBjkYtKweBjipsj7XeTUeO+k2sj9
EhlqpgMle2BkcmMZ0JuoeL1mbIg7EtSCXf6Dcf3+jHwZpqNQrITXkBUA4lB+xWMy
fYC6oMM6s1/tMrvzh8a4HQRSXkgzJqBMHu3Xvvwam9qY87LcErSgigREe1hFRW6h
aYCsZOkiJVxD9HrZ4B4LhsdGYBlQJfcMS0niTfRIFE9ex1xlhfb5/Wp8XErORlN8
cS4fEOb17t29TE95UfwaM4bPRY9bPkpZ/PbKBKBSZGqr/Y5LVBbhQ7aGf0C/ResH
dtbym7CxhEwEtWaz50fAdFagcpDNkZ5JVV52Xi0RBIF5sTQUJVA1XrS9imzDeWnW
am+O8P2O4qB0k6EVAxkxgVlp+McgvtyS/uEJD9OVBG9kVytm9r0v8A9lIQenE8Ho
uLBbg/PKyd7JNvMaS4Aps9iKvuw3g0tRiNz9Ke2Kr36xngj+DPnHIWr0Jcjyxayb
c690pc696C3PsS+PfT4rEoR7LynXr6x5lIyO83SIYEpE/l4C88UFVVn2cLAI4Daw
nSlQIyfINbGgtOGylgbhxeea6OZ3RHHCzA6orLOJRw4C/f1zC8hd7/QeRqZw7lbE
/cFn8/K8vHm4HxCeIpn5DNmq85RXEI+oKTdWYfDk5m9OKzwiHLK5pKA6IStvVb/w
hxRAbGX0boHGCilTtmF6VMnD8NqV6tQz2nDghIXB6WpCR3PdGT1bhTlu8ZDf7oAo
AkY9EFGcDHvkY+ticTJ2NwnHQhDqC4v6K1avFeyA9qdhWlukbE3pXjqoR3jCmqrv
86ygGFGhw2vwoeBp8/jfuyfosLer3QKSY0PEatgXxKP16m38iU9LLZ56L84uvxu9
adyyuPp5zePj8kIMDUGrJcN9V0+jfZXSvbKwSRFdLJTOVV4Lki543QcLrngJasdl
tKs1BQR4anzfkaT2qrKB13AnM9gZ4j9fFqEIk2LbxCxI1FEo4cHKB7HvYwdEJkOw
ghq1+Lk/XNv43J3YOHn/7iugx6GocjlRIzLma3DdDJF5ey2uFY1yQnGDMLQQHRVr
pgVzz+zRS5n+KyR9F2Ig2hlYT4eAghOHeLQNPI+ADUcq02QNBlsVHUYpBT9Pyqpa
1U1CG1iMiXV+AEIrElo7jpuYr7d48zSEpc2xdM+l7Z8PMTisVOneAdFWK05xxVrU
Xp7UFKYLhWsVI10DW7e5lz1J6zlvwgNdHehninQvF28fqTVurdkgubY+n8PJg4Rv
YDlNQwzP1AU1ioQsrZla9VEz7ArJku6vpiKIv7LFcdENSAF5dqq5AbI0YyZbt8Y6
9aFUKPvJK01MlhmZ+jP5D92S694kGWpNrjlHB0ggZQJd6ojNDKB0mglgl3uVsEsg
vz76CiJ9W4fGzZSRhZfsvgwrPP36pgm6wEgfe8oMwmTrr37D44/Jl1HJgWnxfS+9
T+TqsCrD6To609wtfGmu/TfvdwZeh0/2/SDiAfxuoC/ss/lwrzKRshoR0IDurQIX
hUD4FQEvLE2BVlXpvO7or5OKkKzx1He17YS2DA5oKO13rhaOLoUw2x6o2R2iSbxw
pdwuJKnF6otTi0t9UY6jjL/EZ4ccdcDBATqiZZoTBAvFs6DtQKAi0Ym8Ga/GtQtq
BkzmcHJGrU7yzAm85A9JbndUk2GhwI2v27VUdlrir5hPd2k55G/6j8JYyz53ObL4
W2KNnSrrUs/Jyu4JP2uGE83MDB98pMTFlN8GwaUyXmGBVp3klwI8iBQE78UIumPV
HjVCxbnf2Sj0joofSYfaIpXQOwaWBNQCS93cqlQqwrgBngTF//C5RaNnAouGmrh1
0HCXGQ1/kiP5jSeOibNYY01yGnNjgWrIyIJNuVDKkPUTCz2yI2ou0kfinUwm+xtB
jgq+yweKW/PQCb77VSXjXkaImiplEzZQirGcCWDq7olBjp2X1vqQQh7PkPQOfOrU
2kmq4Eu6R+ZMGb/TmIuoPcnoHIaghHZjFr7bY6zapJfz6Q6pfjgypEz9CmR5EiB9
rLioFbQ8Z94eX/CO+Xz9GbJCmnYaNKDSTiSJA1gWze1Lt4m7cQ3b+vfhLeVFhYIb
9f+9kqdFipzUeNGy/l7rux/uUXjshLY70LXwATehQ89Y4gnXDr4kBIQOViIEHXkc
f6r4PwXqlDYh0tFe0dX0D08TJw9+lEme4RCFmOCxWfu4hx3rzLhqQGlX/9/fk2GI
7t7ht/oB85HcEwffV1eNct8lFkXXMCx5Zhg5scTr2d1jlaMdL54GK4fmu5U/GsVC
9I+RHNNHvmOzzLo8KscnTJ1mSwzMLIV06Pch3slY7nQVpXYrdM2jMKXfJDNnpecq
9wnmdX/Ky2XB/aV+YOazOy9SCOliwOOmXdd3PNq6dvDdcAx3o5BXcNqBdbS0M8j2
+DEjJPFM7vpkP8k26YZE+NFSBGmnOrtKI1UBW6Xsm7tyQV+gaRZ1gjPyEgLK+WQN
peT1fUQ5MZxA3OObNV+P/ruQdHSrLeI5tnVEaGs4tRl7B+RuKdazJ6R1mn3goI1x
ZUWIoIrWH5xqnOw78WI8n27wGZOfYLIXcYkGStLXm4mN6CMkvkgbpaelCmXM4vDd
NsHfNtkJ2kX2bCCRxdhimOC5IFA4V5Gah9awLtVrNzHT5zCivje1kA+1r+CiKgO+
c1gM/7uB192EDz6BPDOvKmcGpV6Fz8guG+7J9+K6SPNzi8IGZWr0auQjUgbNp45y
o9lYFpgReM/qr8LPzBWBCGyD7rxBnIP0wH57+MNCisnDjGN8sCfdLc9GkjMQhGo9
MIMHkfdY8TThyMbtkHaVs09Jt76O6BOmn4RueFhwZ+9YEW7S+Z3zponjBUSYpvXq
BbAdMAPD82TWGaZG07GemXqMhH7sJkqz2+0m0rrIQ6RZvzMnEl0wEsKXrJls7N/d
DsmO3Fdu1ndXPgVutRjI9cHO4pwPEALt/FxQ6k2ZjsyMuiaCMdZLdz1LNYfSfQ6v
2buChv/ae+9XJWG4pIDwS8cP6FVYO2Kw6K/9v6xdLGyT4VhCst8+2187ok/COVnn
BnG56ZVhPC48ppE4OkvA3tMjq2j/nDU/wg2wp8pNgdvTuiExUqoqB9Robp5RU7Hg
M05fJRWkukRLuloF43eP9ETgnVETs3n95vxCwWt5A5WYwXNCYhCT/Mm0PJGXhtL7
Pf3o1ncgKNP+A2KgTekwy3y0JHmpgezmMtBbKYfAYnUaS9LhvNRVFQ0bdg4sMCq0
qdirn0ATW+WCy/AFqSD0fQnQVukXNp4R5rR2h3TWP05+4lvCW3Ye/vvffQF4fUNY
EfBFWuybuyjmnn6j4FlquEozDuYRCKYBGJcUMhh2jE/OV+ZUcWllEbE8i31Wp5dK
2htyeCJ6YKVbwZqpjeUQA64z0kRNGwwOqS5lfocrbFnk7PxM7uBOhhI2KkEDIFem
BeiGUYO46fv6lodRg7VdHRIw3zVBqoNL1Rt/KZWk1VanexDViJQtdrtnRPNBJ7BD
Zj+JqjATEQkxnAvHExn+qo3XXJAC7ltjvZdtY9sRGwVtBW5h5GStDi+Cv06e0jkR
Lb+ggheW8fMYyAb3t+OEnm+v58Z2fHprlGRTxLMMotIBqb8DSCt0GDdAMLbv+0KJ
xWrnXljTLcXXTlX7O+Y1V0MHBKPxKpMnA1rODrZ9hudbC7OMAuF7HQWWrfxUZlQ6
nF+Jfd3E14SEc9RZUeug63zp9Lcr7pOhTZUuYBVnJ9DEmfiqqHR/RTTTOSwjmV++
QbfogTTNxDhRtQoNTnzxR1dus1JvVjD7E1L38dKJd68RsRqC/ncbZI3SYs5YND20
PVhFbT3uTFi6aQrWPULScXBKGH8SJWWddpIizeYdkOIFsXm3WpaEqtV3duppIlYa
jecjuDYbi5Ig3wrfLH8wPNJl6VTMSiFUrj/A0kNCkla72STz7Ewgx1TCqsaoz55Q
e82JzXsi3vaMJQy8GnUqywvvm6XdpqHsXZc4HZkFkYIJtHipMgQIGSy549xZQ9SF
vSngzwWt5TIfS14e+1wCjKNzP+PT5UXjrclcMsb6o4T16ngmopb58L7dYyOFRdWP
1/9kAyKNhogobdCDSUnM8hCdqYkvOWCxdrHxv4sODSvOGSmRDzhdgKicBo/1zhVb
hEBiK15nAdq+yapftQOsp8ZJR/GK56RjCtcUKhmeeERkyEHE7t9TRTOUKv3wUZtu
P0Fe4S9iNz6KRC0yMSpkK2YyFtm15nJu9taOkS0d6OoRFaEsg/Dpu+e7lqH2ENJ7
T1mpoJRsTOsjp6/gpCpMGz99h7YhnkBzy4Ejjlf517pNwtskCj4lKz8k/2tQ6JFe
KRCfy0WyTT8K4DlUK8SFDjRqRHBumRFbFBe0IhASSqW1x56CjMUOtF5sIU4e8iCY
LxoIgqgtazXxDPd8nTTlYLa0qsIEq7Kw4OemsCL8qIjNAM1zcZvnaM/rpq77l9w8
0/LeyKQ1BduII1gfISvUKQWIsw0XDcSkPVzioQkO81a0s2/6y+eioqjIMjFjEnCJ
ZkYk86Ka5RCyBh+/I0LGMkR905N8pTjhGs6jCnpGUHTJxVDAyqqoSV61O9QWNYxH
94LrGGI24lgXKOt06holi84JEghj7ZeVU0yL+gQXLzbXK9T24SwMtSAwaPV2EPRR
121hQ83O2JRTvJhE65y9rVEcD67tIGz9OeUYt2+a90gW0BD5bkl4QXZDbYwMe5MT
L/ZnNJS23KXn6EF/N0QPC/eIoUySjOVxrj5pJIk8Y+eee46qK9ITpA0n5KGYHHRZ
sTNXktosqgn/kDuHP0G5USiHQn79xMg+BjS02X6ESCA6c8cFpckhPSD9X9r+Wo0g
5xaaeITOX6uFTEnq2Nw0RUOXP9OmKOtvsnUaSzm2FJPL42PhkIUbJ0jd2+jkiVDm
ixpgNT2WJ5ZWn75JuWpHEGCexB0CuFt/Dpz+XdY+k6oIneY/UpuL38eDct6Z/6y0
8/601RzmyHui09kDzLb0A2e6vimuwBU3yxDgVEsmgxwD7jpm1DN1zXf4SElisEiy
NzL4GKJQ07xhPBmErsUaCpn0WoTt8EBdcO5Za0tCgccnK5ZXzJaag6H9yPtY+sSr
AKi3U9il6Oc/h6NxqUsKeGknSxoSs15s+CuGzYMGLoa5FRen5NhSGjhnwyvmI6RC
7f9w20keIF8/peiEPawtz295j2GW7yUfOATb9Pu+GPFu7Jmg3IZjds2Y8hE3grrw
o5+M5V4IG9RuZqS0OdOYK7Io2lCN8JDiBRLdd535b87uAr1lMXID7tlRvstgFFcU
XO+RS7HkX7+2S1HH33WJd3dsKr5ShxmgliDxqg+6pW0Zmo9O59G4q73S8MRHs1jn
G1//VWf3SBAgQ60ILWikXIHtyN1wLNp2tmHnGedbCHOYkB0AA41CibUAwxdmWN+Z
SWo9idhpT/M+r3cy5j0IP+8tnIUkR1A7af0I3aYyHnfgKUT2fPXT3bdT/kF4Skd7
BatkFFo+/imREOWjUTmhl1zXCoPK8wreJBLU5azE1xoyX5nJl85ptwIDy+sB3ulL
06bMpw0K+eGQZ07I8zeX1/s2mLQtIjCDMgP1BoCWUNCoQ+V5ORJ/gJ1BiF261RNZ
BLCiUG/Bu8feUEwmKX74kvkZLZyE71BxH1Bx8w5i8Fjlb6RVezcvpd/2gPviOUIk
aHKJlWAn8Rs+FElEAgyCBgXyeki09N0jIdKEahQTZJZE0cidhlzEWYnYL/mzCukq
m+5ACtx5hnElgZXYcIG0YJZvmeBRWasEZam3u+/fejoitvQ+NuKO/OnTXu2hBxTl
jgR/2x41iJUVG1Zwj9CCuysl7LxL5FNZqFGCnHRhtLI/zmYN4INQHqI4CZhql6oB
z9wOgnf9Dk/5AZPRw4APcYmYtg4kSdNQ1b3PPIwo5ewqJ5SeDTDxDgs3lg02c6OH
gKSRZdGk9qKbYRZW9OX7flnUrbldbRKwuqoM57+ofah1iOylQEek/oyqv9jUjItY
d0XRYXGuPk275rB/nSC7QWbXUSEHak3g7o1Dob1PVvkN1S8KuduoNC+A+oKE1gau
FqmqM36ndPEsIyKvk7HgmgFuvLxCaGf2Kl8OlosBFwK+Qq+wuxpzmsbmGyz8YiYM
ifQiQbuUJfpSP0aIYUgn4MtSfzt+/v+B48TsHTuLCpTKpcJyXtRIE57vtU5K/5Uj
Vw02p7blB+7sda1GnyWO/PGGvaBu/7CSwUCn3UYYlwoIAKM7w0Px5TDYr+eMCLDc
bJPFmSgJiGcGvaDWkyMxcqgYY/5lb83tBxgq66SB269a/TKy70OfvS4sthG7PX1o
awTY1AzjFSCM4EAMm8z53iKWbtb5nUqYOiY0zMcqGfNqkTz9tlOrOQHjjs919B3Y
k9b7niBJrg8TBywdjYLyUooOAHoy+Rh0Dru+G2zdgRiPKmYNihfLRZpnC98Yrlmd
LR93XWZ3fGZ64C8E2s8D28MLSo+EwVq0Ove+Ow3KKNfcrdBbizpeJlPIWn5fJ/DZ
ho2thEf9gmsyqzNKDBkFISHhYx2xduUt5ecLuyB5GJtoCQ3B44a6xYWtt5c1cpeC
g/rmp2EcZP08MrffHw4EYFdVO0eXyfZ5tQ9oKEFi0Ssco1JytqsTU+nvuggWJrTV
dsV56XWcxkNqzzvNc0i98t3gX0RFw/jG5uY8Q6vDPs+8BEBx1Hwvs/KXlfRTrfC3
WTV5zOdoEPwKfNQO24NhF5kcgS/NDHwZO8Y7Ug7GA9GHUZTzoB6BbBNPIvPihJ25
Gu0Yd+m3UYGTkZYIQKunGzLLFYBZzIRHw4UcSYsQdJq+D/0tYiRRdvkudVzbGh2n
0ovmxre5X2ar+A4o1rf4pvzhZk2ng5SuTpl1Ki5QKKOEQpG1T0q9SAabvsupmWt6
7+IdX/wzhYx5iIAmnuS2w7G7636/ObaxBDbjwtb13Lja3l+kcSb2fqZ/r03HYdlr
xDqOPMdlEPiFdJhHewLGRvHZbIcKN3UQe0ewN3WPOSUmCaiD5VZQI87L6AJj08/7
UkG44CFKLVd4wtRz+6RNp6gW1Ro9vHDR8+LVdATO+j4bOUHMTWy8XwpwuD48a+or
S21oRpQOdUUBEUYFFi+K1dtu80yabmzKSyEvoFWBW8XT4+RuomuSJj6R3qIgmmCs
fiHvdYwq8mvlAJI+BlUGhqVLD7L2EeylCZdTB8SF3/7hYg56Zn6iZcmRijTenCZw
3L5eOE/z8/GOzUpp8JcccaQJQfm0CHL8tuBuaxlgTQuVs4n7jC7OXkKuu1Zet42F
Jj06FOUOUSA4mg3fqdjxIjB6lX5M88KJmtGZ+x4fvY4yjVw2wphj5gVZoX1mCRwi
hv00Oillsxc5VZocVlFzu54H5KDwFkArEw4Qo5Zk5rh4/T1k9fgsDR9GnFKRp78k
ZqzfVJ7iHwIAHs7CiGNa07qOuZYgO+69Rl6qhyM2c+/qGe/9v83Z9kiHU7C/yidt
IEphDhuM71S9I2a9IZlFfViIjU9UUq1ZxpzmwN1TkoTjJbmRX/ZvvE4oasE9h5Q1
licQ3SCzQ1RVaf4Db1dcv1lNLKhynhMjMxy/7bJaPFjPHrjrv4WoAIrhHLaKRlhk
zsM/CGF8ogvJUb8wOOtdJZLzgzgYex7NuF4x1nL/Eo0IBOMoDJd1PqaGLcTSTWDP
5YgmIWf7WvjJMSv1LIo2PJYJbfkTxlFmQ64DB9f1rrBPPyvP+F4/K6GmIluBiiV6
NXOpsBnDPlaXABvMtiKNhRqJu3wpK8ccsWexY1dXsuiz6apwf2vaCHUESvQYzj96
hMNfJ67TCaGaHDjfQX3yKDcsvRTmzxU7/IVU5d1AugbOkqOL2nlPkubgd6hd5dBu
8LIrIlCZXDxT74udGCz3aJMSv73sFxPUqXk4ZBaXphhX1WFDkVX4xdQYc61J7O7M
apVg61DysZ0H1y0mj9DVOWsxOX2v4Mhsyk/kL3C6qqdu6V8COwbFjHxgZndF9n/J
nDxhauq2plXKXO1LjEW2W4APIABylVix9/6RlMq1FBv+cYszsf3t+qRoFf8FRXPj
j9+YD+vqkx1q91FPbv/jun8NeHeyca0SOQjc9KDkVkxQ+b6bPQ8SmhVpnLDd/V4g
aCrjYoszaUh51s1P8LC4QrCrGfIERodaWXhM69j5Yl5F2vN9613PoR0+5CYjMCe7
rY8YOhYx297sPIcBWpZzpa0+WT90Id/QgMcxdvOL5e0yAJQzfUIMfz6lY0iLgBKY
CW64tRkyQNivGofvQDAmkSINKjj9JSI3I90fUf1mWLlcdCq9m3haPmS95zrtQaOL
71EaIjTOX0HeQgrmfGRlmnb5RZPnTOTalha9WWeCj0/EqcupOq6D23cssjT4csKo
A5gFufvP/L42HAmSS2JrxfxR38nqMgRFJ0ZmaNyun+Qb22xfgjujYZwOsRnqCVfx
wwiA9ZH7Pmdrzlzm/GchNPM0uJDJ85blF00h0YfdgIdQpacixfO5WU93lNWLZndj
H5SQOMQVcLmTdnwSue8OhOL+Wug1JrmSErwNSeE1aArPbhXW7c3G6GZNo1g0HwBg
MzxRvTprVFGS8Qjlen0yGwIHM6rgS3FdCpWrydJMij5nwkLO497KW06vnVKpDwrN
quyNRpSvzRVpOkunj/LS7s8AIA5Pngut8/mq4HYL7lXbfausO0uI3xA88lOty6Gl
K+k2dLV88IUGRAzKY4vIlAMj8D9PqiES6vLk4vp+gbzPG4F25ka2By4vX9CM2QDH
UFcqT4uDFIqAXOwg9OolY3Q4RuXLPWst6UzXsTWkYEMvX63Eg3Ahh3sYmlLLSul6
HwmvyLk8SW6gBj+k140s0Adhkl0qWxSbwToXJhhije/6adr1k/KAyqL31ln2FN7Q
MuO2nAAIGGkPj4sKzkwzwJP9hpyh9xliCiDumtXrP4pxqwneXwteDnhZlkVIYycs
zFxypUCarTs/OAib0rs1N2pkH20tVOgrLx2/xkRGByxTitYOLB1hBQOYOrpN/Ars
n7f/HkMRqn8uwVxFAQNqz0zbszh/TKBCwv33KzXL31uKeWBwT2aXzfzG85hT9/KC
zgPUiWbtp2vC7p3xDNfKI1qIJhY3DH96gy900/Vxhlsk60uWfK3rbuCNp0jCpUpx
map2/mlNmDeh/SMBcHfL7BgkAZRZ2Bw4QL6FSQzkHgQBqRyV9X7UtFJokidin0x+
RamFXAXDqjrnVQYULd/Yv2U0JXsbZxd7fMj+PEMOpIs4BBLw0i35sQQ5MyARY8mj
48IvZXAOdfMXz0tx06GmzphRrCoZz4KFP+Tvf/nXABW6019kfjBCWPVGSmP6L/dm
uSSiZw1wYDYZ+HmIMDz6SXbIJRWi1Olpk/Ujvmcqy+NBLYtY3JbERufHsVFD/0Gu
8J5Bc/nm4azSqrltcbblFs+wvSeCsiCmFOd90rQIvAA4t1GCRn3klzz9Aq9u91tl
hGDQikHMGrjQdQI2cNU4b7qZaaAOSku+2r7neTaehdAPUv9rvJr7AKflboBsJ0Nk
xNlim+jJif1eVS6Nja9jIVru5BBA9wq5noK2vzTULJD1pdjQz0sdf0dyMXCvne3Q
Cq1jWjcEpL+hzJOnJ7nPWI8lTJpUK0kk9wfklBjvMCF0bkijM3QazhJ5Q0FdT/cy
J1HPeS4BS/5nONwLxog6Ej/lYmPKh5dMIGR1y0V7LMzaD7g14X5sSzcNuBsfQvIe
4dCsoGR6QgBtm1apZMW0lJZvo7BxcOC7v8f7kuU+DrE15JWB0M1MVYIddycK65G8
ljb/m7YLXJ0Fjy52Xa1HfbELH0uw3X/q5IF7YYBy2VA8+8bsoPlQB4Qj2coMZib6
33yt2WSQEd1rTZIzC2+i9K3MsdD0tgRiNwJK4aHb+0ra+YU/7vGVyLrfDxu4FK1u
IF/Awo5q3zgdYgsKQGpRVEfNkrucgkwRq4Gd2UF6npyma7JElMSu8fVZG+RyDMat
1p0NWdcU/67Wf1OcB6HabKrIQYSoMK6OZbhI1+HruXlgF/GB/sbUBa1mK+hwpMcW
l9zcszfhc7+DJAJuaQAlImfQ6W+GV2O1ZqHo89+Jm4zE2235pGLBKcN+c+VrwHBj
RPUllTNWnv+ddFAlvy3zAc4xNe4eQgwfwJzW8wn35f/TW3wPo+QQVdti1s5Oddes
w2QZvtMq/80K3vYsRU7WtIrqCZQMjfwpuDEePDQWnqWLT9MjYV/X8dBToKILBlWX
O4AOIz0+LF5yz7S3Zxnb35hqDu6ceFMT3gpXkxt0XekBNiLLdOHwcE7fng8xktX2
t7hoOtZocb8Rz0Yf5WLcNKPtsRCjNShlkus/Fvw1EcHS+8tPdEdmbQPr8ap1ygUV
7vyZQV+mK/6TAlXdyvDJ24/hAt3TqB+YjsRrt13Vw+KyUMeZ7I//+yjJ+Fnaz8TY
p5egfQlNH59m0PVjblCzNJiXXv9S1/mUER2zguYdE/9+ssqiQFn6PirhGUgiPazB
2Mi63xkiS8ZLqZ0eTIiBXbJLzbUMx2ZQ3qsPi6i99LcskTCZIiPpcSt/bhLETBmD
6vqnTvNzZsYbStM+vO0y1qiQ8AtpWiCJsCtS0SQSBygKbB9HwT3JQrbTRG7XmobC
lDfc/ynTQekP2hGPsU+MagpVNt4KaPFLdSUOVXtNx/Eh5qNfQrl74OuJUjlww9gD
fPxCJ/u5vuj/nfkJryu6mepWJXDQfXs7pxwLx9RxI0OuA8RMNSoXUjqdJJ2PNS3B
WYO4zhrUFGPbWYfsrT5xy/U/cBjsH4bPRoa1UPaPdKssXfYY6RF2FwJlrg9OFuiU
U6GlPHi5Fq8ss1ZgmcQFTZWg2CoyewV+983KAj2mdFBO3z91ej7g2ROtnB6VzGKd
0Wwkvwc5V/JoR2UtfgL2uwqiJ4FEaJ1eeVcqRg3JWOhFDIESySseu/SoqZFY/Tjf
s1JhAKOA25iloNZpO2aX2kEA27ADPJYpaO+q+qVsmJNDdSUuJYeGQRcX6sy7D7Pf
qFeGaH9LMqpmzaTlWH9A+RW6ghUis93NSsG8oxog31Kew3TpyTVei/PVvWUkpuaQ
w0HfJwKKQV4XjI+yUgn1aCnYFh/5lBN0ksAoM1y7nxNHByyt0hN1+PpJGj1/h0I7
GMBBkZEnPtIc8McJxhNsbHpESezuARTCiIQIxLEQskPQJAXb/NBI20Rs5C0R1weL
w6FWyinTOeeG19psPOv1265yx/1VzO6BCpg1c18Lo218d9dgaI4cRnk5frY3nscm
HCIkDxoqc4nC9H6KrA9tGQh6mqaI0+ojW35E4ZV/HlkrCHn7+M9iLrkQayBBQD+S
aCl5KwXeNDOxXB7sb8Hyy8d65gK4KQOlGn2ESjAqtX15ziZQnCR3UhMh4tv+KHaI
uuFHPr1hVTPR03X9I9sY2BfJsjhdyC+bd3kEAWZhWFZ524sezEEgxbU9zgRFuh3j
6CYGX+2OWmQcY3gNvfYOBZ2gamQlBUkLWKxfu5vtubXuusxWWJ3Z+KseNNdj3T25
q824xiz+2HAN5zAC4vFYYfucc7xRYvXgn++oj4tUOlTbbaMNQg9ZoFyWCssuOtf3
YctGb92cWMID51eRjzOjZrN2fWmOvFIJ2sb3IyfQV0Q4aPJW9UzxcL/esnRL1mQF
bd2RzL+RirItBbhP7duoK+6hocZKDVnZh4cjhcrSmHxpqSaulfMBOaOgPArmafIU
2cagfTU+wb4cOy/MuuKRcn1z/X4OXsKGK+JtMT4Es5Fd+tQiaKhD5dYfFsRXDKZR
rHB4/Upko2Pvf/S3NOvwpwxBQ8VZQqB+WzRyT6mKJRvXS67ar5Fi5ZCGL+LXwaEs
OMXF1TRDch6utGFn8ef3Tp8gKxb+Z204Kecmmm5+OClyo++W1nQ9RSyYpfbUF5fA
TL+ImWQ5lSM2qORvCPdra3PK5apgl42pSrZX/N/SsUMOppgBZh1tTxQLzBGFYmhU
VocK07asu3FAcL0K+S2SsKu/J5BNLoZDWLHJbeA52JENdpv3JFOJ73kZiGEbd3S0
m8S6V5dnoI0a64FeYKiqovZWuwiCsUNA3XHHIZYjtG5YzM4BEjURtSFL37X9yhJL
AGSJTI4UUWAf+5XpPhH9wRg0jmIocfjwPYE4VAnBUUKh0YTwEHnveLDKZJQn3YwL
VUj2McU4ne/Kij4GT+Q7fxejMMXDY83Htw0D0W+YxEObqTdb3xdqejuqJBfq13bn
WCKFMPD7tuhekNA5SO7ex92rA/KNvqFxOyDdBEZL0dVHaOZXooX4PJ6z3+WN8UZn
NmBuP54i6Sw3bkL5bworg1xnj+mF6bNJpylml1fLJzuO6273H4Mn/NzrVw7Xmmty
YS/Z1pFL3IZum5i86zAWGzwY7rUalPD+Ywh2lWWH01M8oY86bIsGxJKostRE8opQ
/BpAKqzowJ9TaKJXBtnY6/MPvcq8kenmqzREpk38SzIiQg4Y3XliBV0tODWydf9Y
A8dKy1rRao17ygmFyXc5qdNPfbwWRFFwuycw9XhAePvw4tjWBPmZu1OcYMQFgdVn
TN0DiBxmYbofNqp0oRGj7LNQcN0zqee8qbsGhJk9SP7faHmzB0nA1JHZjeT3VyMK
GUiINr7yYSPo5g8MuBaeUjotr5dcPuQnojOvXm8cxw2PtQnxVVpkaZ7WIuH9Miu3
mm4bnxg7nWi79rpPxG7xcLLmkxvrJ+8cywIKQTt08IfLJiZRf1Nrn4ckh143CNHS
/OGwl7gVU+nSAXQhhi0ehUInieHxPTQga8dkdsoab7Ynnyms1O/HZ4NPlMapMbMU
4xKw9+Hx3v6qh7yux9RYGcb1JMEgYFu+0Bc1dGt4JyzcjAEvAGDAkq4fnikBGGj1
mnfSAPXYZfmq+O4aki/YneyoZfYrePvbzoQ+958Rqv9vlK8VgOTtZTSS3GlSsVfb
2hYUCj1OKhdxHSqPEJ+YWbseRX9qWEeoxH7AvhtwcZ5G7XG1b69wej6lZYiKsO5M
wY98uU9a6q7Reo34stpGb85it0lsKZ8PorkSpWHaTLId068g0RJWQLYH9jNYiFmm
mGDjk4dybD0u+ovdN6ai04AlaSbPIDoL8iUZ++WmQAnj0lJwiEGnNLV/CIbFKnXp
HdCFTPA8Jj4mLrTud8kJGTTbkPflrpxY0pKe4XpqggOaAKwiHag9FxSa8RA/y4CR
mkICCR4ZGJ0RiQh9Pnq0TPox1cg6tL0mpvLScX7/97CFoRfh1EXSlkMQT4YoWSpG
UoFWE5obp/bCSmZ5Un9d3hEH4bo7s3MpGKcY/+ED6PI9qfP9CLVDUtJ5vibZZPIn
5J/SZnTdizHNlG8C2xqjD5CYdlPQGUtJjNYI0vltJquClE6k8XJtQLQw8lR/NQPG
lA2dps2bxaGoQW06L/fVFXSVcKu9kgdMGzHrZYKGIsnASobuJs4Q7lFfWR5gzQM8
XCqh9zw3CSqKrk53N4aMqGNcn0zU3oMLcZjUDohF5VGa0Xd0KTLf/f7LN3ZN5hKt
x1NHrJNpeSUjhRvnKwyheQ0zOxkZNNbmHVDywAjN7EXQmbj/7VKfyKi4c9otu1mc
ixKWTmsCNnA0Pzp6Aw8hLYEHRnltWncE3vaBIo1m4xkEziRvmPNLKmEn3f+5YEjT
hjXDMtLUkdGbT4HUrHkHvzBtHRQUyx524gkCtsQBtE4/xCTSS5A/7f3Dmu8Ck0AY
ifK7WJTcCX1438uZYsYSISgEKKxA02Gpa4IRV7Pl3WsPKqoe/kh384aml7MEgRi3
Pw5PUPBz5glYa4PCxEPE3X9AaXoRE8NsgeafUNIxJYikYY5PI/Sfm4snH3i+bWhw
JC3kc+n9DaMfvYsqWchrVRaEs+UA5ZkdSFOI1vAdIdplpVyTHnVGNyp8EX2n3oEW
H64jq7S0LqoYUOuOURDUyebNs5Ek+mTYjMjYHLuT65fvYyZGqhU45pstpn+e8TXC
07FF3aQG4WGhGx9m5XfRJ0gWhAtysLrsnTC/nBxXp/IAY5XFpKCDn/xyp1zJ0UzD
NvhKKvhdf3KrafJvfsOdtwnEeLUJ/jc8cvnTUua3GVObz9+g3fU0cnpeJBkDLGbW
og2PnIF5Zu+I2lBl46cgddhUdIGakCfy7pCXZGmMJxb++ewFNA+lW9JKZl/vZpe2
baDa+9sAk86G1N+wsydXx3tSJbvIVD9as/YA/uUczimf2TscujLa25D74i5xXp9G
suutGOSRVhweE7mq9ccXTRTXECNXKdpKLfACTrnBHzIFJoUEP++U6Bb5LRZmGEIh
gHniEk6/H+7f37YTa55r9TiKzJzYPXDHMgjIuKa0+I2sP1tLKJQplqXUKDqZOV0H
Z2R8xdk6LHnc0p0ODUMJEUy/inu7ILAXvbkv8H8HpHfD+GdiFrFVbOw5DbCjKRQa
5bkqc3fttKhgXPHjMpc0VQVKxB5XIJfqqB9JIOIi4snK3dnI3wlWMgd7SFupyjCy
DHkPBdRjaNFdvB2iCt84yZv+hN5NczvpE+YOeX2FV8Fd0aaoDGOau4+B1XZ8s87s
TO4cATUgHxXL3s+vqIzTn0G8mvuZZOBRZcGzYvf9NIKpG5+nu8ikpxthl7/zNM/M
CjS8asitol9t6FDof2nhdjA5PwnTT3j5Ni5pAYkIO2YqnqA3TlPjtbBmK72Wht9V
iFAsItpPckEJT+JhQ2eXfRmj2IPpUH05gDiAMpEIAyIHoZYlsvUTzA1pjC/0vFvl
+0ME5k9Ny0pb7FL6xJ8hVGD5EiTrX8LflZb+sQoKNH1KxUWRcuwwr9qmOO6b7Ry6
0caLTuy7zyamGM9QCnWIoWfEKk39wFiF0XvqzaFVpyWFmN9d0yeEO+iCaXho2539
WVqspKx8gwBJgsR6EcJMGkTrT1+8xGfIyv3OYLH/PzeCdJU+BNAKY2H//pQ7x3ca
xbSzwSSQIfn8lV/O9CJ3ZW0wXkqjNZt/FAh17y/XJgxzJUYeQY1X6ijqOu9XA2Ba
PT2NE3NYU3P45HJ2ygqsBmnLNRAocKMwlIa3PzDjrS6y1gnGGPdNNZo5Q5QI85ig
OpWJ1XIOoPqRjtwqlvfEBQE1acTPcXZJhCMJGaXHCAkVv3WkQYqY+iqnaEbKaGwz
M53zbNz2bd6IhwD6lBrSGWeHLLz+g0Miw0kIMsfNw99bR7Db29nTyC1GvbrZuka0
OZ1z18ENazyZKHDfp4vKNCDvUA3G6l7NvGcyNkjYpZMIlmG04xIsdIPAIg0ouZbx
du7lZz8iBu5wnd1YEu+Wj577HAmvc5x9TBGz6uNxfz44g1nh1IDVzLOQ6egF+YVw
Ng2KipWISl/+ZBuljuWeqNyzKX4LV66NlX7GD/LsE3nvX42UXWj5mqGDxPuihutH
+peGnOERqTqqs9gKxzAU/SwXjNBEVSmlTRpe5RG6V7exqRy0mPgGjDK3/Vzf0T3T
0EnDyN/CWgg59BMB1p0qV4Wo8fF5xmztY7q0Ycvlsq4uyggC1Od5ZnK7TIxetToP
0OYIr/Xhjbu1AqnuJ/b6Sk1VjxZloeY+sULYtA2nXW1dXrp9cKKk2RsvnAEd5Wtr
dKEHNknC56/BuOLmHY61V0cUdyJNg8ayNHGJLG4gZn41Q+ji0DFNKR2VKIB3b8Vp
JZ6Lwrvd/Ev+BHOXEdl6XVs7nfJ4xtUMJhEXtfp5rlHbXeEXNESAbqE63SrZpV8R
p9jtqELsPAdVIz3WNHdVMt6SarlXWMpzi56VWGAQHcT/Asm4cJOctusq7F5sFfYW
oARfp/0e0Y2mevoIBZP+hn7QvDDrjt/PKV9ekeXYqQN2ydLEY+NH3evhWpeLlwtt
m3ajIwKRACtR3jdztkxTJQC/4iurQ/2cc0aotpRPK40XLvIsOL6/5p0MTSZJQ5M3
SAQL7Ahyc93UtX+dgzNnHjMKeSHD2cqfvv794s0uuVvs4KZu303dLM7R9zZ2T2Lz
eUewN8p1bIflYH3kVkzJEfyX5HXVtiEH5oMJJ0QtO4U90WY/u/EJB7eyhNjacIB3
8num6JaxOzaTqYjyVYLueSMuuZijYP5XI3Ck00MVBZfLlseTHa/YMCtE8Wa48Cfk
oIcuOyGYdQoFjAp47jZeSORX6B/3leCYA1W+kmLGSbzhZMLJzwJo7twF73IjGhx+
8g+ZRZF/KwmyVPhOOiiCrHhvBVLxJ5I4HHM+lBJjfbtWPtxp/xY7dxtaCd3VioT+
ZWfaCOtTlJ/7J1o1YKwTJRmnLVf+VwJOQVbQfNbbiP/6MiCLijU6C7VO/fUfOU0o
9DxsRZucV5+LxrV/+JHxHmxbwDcKAakdmDZiqinC8i0uDCpE24PgolzDUDGQF7c3
5PM7HPJq5AfX2wZLA+njrzXFk4A4veULqmaXuwp/GD7H9v71HGPkkqjME6zXsj4h
p8ug16OLeH0VA4C6miKwQYml3ea+ZDKC+61f8lIs8bNjQN8QiInZGtmsfkpFNHIs
+izRpMrIGZPEUhYlTxM/19W5dPY7QSFnuxDWNs5nTG+Hf/AS9Cx2nQyo4HFtpsg5
CqDYbLmKw77ZyNkEd4cVUdVf2N+ZpQmK1DQnYnZshao+ftLuNsCu7+woyAgQe1LU
FOEYq3N7ZyiK/8Dy6KaCL3z4/WjOBKVAPmAO6eDE63E8dp3RDzYv1iItK9DADBUp
V7wcAe8uLmkAFYfd5rpI9dhFqXnsPHgCd2+3D+d0EMuEVkM85V8RJ1pvBDTC+Ve+
GvZiNgZo7OWEk5hCawIhn4e+sJ2dthBl9XMXS2l8e9QmspuNu2oKr7UzsuBpbgC/
kSUdmh8mq4JyXFyOgcEVpoTPWxluy40H2mBY0+LcYMsaqzeU1ZLmirosnqXBdik2
prsL1IgRP5YxBQ0kiazq2WLI/qSIIAOFja6pTK/vLo0IiUgqTxFHy8ySXGXd28Cx
6vWh6ChefSLICOR75f5AXCAAr822aNv5MzNWfAWa40+CzyyYtCHs6pQnkmKbwLxv
07uJoCAhnAcEeT4e6Zfb9STBZdYmFZHCxjipepADWDflqEb4KPR06zQDjgkcSk4E
TKtGTYaJhc5/1nxDWCybiAYPsxAzxjoJJl6GFN2XNsApXN5FbEai/K2Wra0nnkkt
U9pgubmuLwlNmqQg2k0N6MELghusv4/GI01NjvJt50pk5B0M95zM473RHsiWR84r
cDAFdEvnzGABVgW+LytOhnMSLDEjO7S2ZCdBiuUpqr91K7c9MoGNr7zOuAqMSIyV
0dAmxnjGHRVd4755fPG2AuTYYxwYNqCkFB9ci0Gj3iZq+R4r5FVtNAsfsGSiHloA
X5jbyBtz2GcDtijDQMlGO9aOS2hGj/YKqhkK/olnvLrNxA8NEpDRvrzNijr38h0L
E1CjMhOX+frUhkjbymF8i/PS8HY+RDssg+eD/jWFjA6jB6ehYSsr2IeiMUEZfR8O
W1jCnK08lgPe5esDxpwRqkoPblJG7xS/YA7H+MfFUD8nzsghB9r7XCIcNB3QNP1S
Tsc1RU1ursdmuqNRATsqZDOkkFjil3ua7LWPUGSlvhXSAonA9vWuXGwkAJDQy88q
mi6B8uppLpKqmH8gQz5gp2koLQwSLXi48EIWkZvnF8AJ3DHZCGsmK1ZF4u62EWWd
PXxgKFNei9Zbhvb8fiLSBJdSl4YzST99oh1GP2JriYteZI9OQ68CO/X6nxjvRa4r
eHr6sUheDdQ1H9qYbs3s9qvK2OqNy+XGDpOoGypx3BexNgvCZpFGtcG5uMZRtWdO
8d47Px1aT+/R8sQIL/90CnXpxTFUgME67HuHEECWqIq1bVOtuORkJJ6gze/3CuYU
91DD8ZHvAYvFSE4asz6vvma5oh3WFnjwxH7qrJC4Hqit9zupB7dbrs7NE3vlG0xZ
9QUjcS5BtJxYQRGmHCIPBmojkvrz83I+7z7as2U6VAwBZ9AGL5qgwEgCCViGpnJu
EjMEXRf0Ckct1eCM8+zjF5HXtfiBQ0f04GEXIz0LL1VCp7S25TShSvCv70sdtdoT
ynzWXXdtOtEkQzj12Olqwq/B7Szgj2v3HEFZMm06qPnQFKUxH8mTOa1EGpctCcPZ
yocmQz7GVKSqtYMOJcXa9kUU31PIzXRdxxB26WDbDXItkyUnrBCgbX+HG4Mvn6Dc
sEn8XcYZvWThN2u2nodU8zlFKnObHw+JO+MDz7VQzQpK7MxV8p5ERYxLEHYXrTAR
6TuyPEXU8HK6Ivc/eNiDBhsa2Ywi9jsUPpDk3NfcK4Dr8wwLRQjanyy92tasGkWL
M0zglNSw82p6ndVkiGwER17qu5GbW5p/6I3vrBNekf32Xa7o8/w2IT6KHxHY6Ft+
LbLeLJyxaW2oL/gUi9nOR8enGZYo++5zraX6NKsl/wPt/EKWGmb8TKEKFDgb05h9
ntd2oP/G+UmKhEd/CRps4i8+uJM34xJ3V6sbhcGZXf9IYdQLp9cWqNaKU9hBScfv
Xo+jTXQCl4tRUb0J/1kr/aIfALSxub9WC1Dbjw9n627l1RFLNFIQdVfapghP2crh
4CYoYFGaJbMIbuKDiV8r9IpSiF05cjQGS1XZqJcPlR2XkN8cc8stqlsHWvXe96Za
sk0LbheEb2TcvmSF7oqJ4SqSRcGN3hI57aJHnIqyU8jCpeNnNoGX5lVoFz9xv8sn
oC272leU6DY5lsYgMhAfloBPAOBNJtCLO5LydqrLrYf1mXrpnfnGuk2DHQ23xJel
vzMJx2/8FZvbdCJsUZ/lB7fxWIHjzIyQZugNhol8dohfbmrVHk/2E4Uo3xR6BlVm
9NMRLRYXNVZ6Nd/0T4wgMtM0+9A/36kz4JVPkqSbE7cPnIKx8gtz57lz8/qWrlrA
6QbMxgSi4KLeS4cctKzl07uHJ8IT1gH2Hj9AwLQ0wGkJhWM2sgvqGyAH8rV3OgOy
+KOP6JFLX7F6ak1lD4vyiU8V/8ZlxfgKqp3skGiQ9SViQxr4djduiyHtCXlZH6j/
70T31nQ3t8IRNpbNU5JcftcPtrfHyJ6m0W15LshVT9tl12mI8xFEawsk+d1L3D6J
+IhKQTJv5enSTZzXFtML5Bl+a4egED5F4hIH8nnWs1LBrcgGyG6XGYDpOF95c30x
fXHDtQQbD+Wm1gY3uuq7uGWpSo8QneyKTqDOiwTsM49EO7l5/ms5u9sJJvCiIAFi
Lhb5GGghg4wOTXv13/yWp871FsqDi1Ft/KwSUd8ant180ot5lOYoRM/kugh9LDRw
y4Cs/v7b/EBSCyCApDwLdl0J+cpzBMmgsT2aUUjzNHXS5swkGvkPAqsOzXslEhNL
oU/bx8SEmPE3rIZH1zU9RlHfaONs0v2BX5Ry+re2fdSH58WtGm2/YJv4o3q/+Kno
IY7l5431o7M/Lo6kzOOTOZwDe1wu47bPAe44VlLh7VGQ+hP5w9StladCfsmV7Jq1
6GPHSE6rflKHCbzNWkWI+Y9PJqs8W1ppxRpIejqkPRWSeMpIQ+ZR5sOtsAQDEPs9
9uz/yBB70D1i8awTikrFsB0BFk/nrL36kxXJTkMxEE9jM3kbHQdS/DcDtOgtJNE5
ZZZZnfzKvYaDEgIFLtTGZdyo9RExPej5Vl8wsyCd2RWsDXt7Ro5f57UmjKLE90oG
aMmeCCsGDrkYWbhUgf0vD++UntHidbG8TYj5GgzCh4WBO3ihiBpQKLiHmmumYopy
cBI5IeqNzvkB89CHbPQv2rysfI7IKGEA+UKSU2ggJMnWHXtgn9T2m8c0BaNWa4Ox
gr3X2vKQXxTIlxyAsxCRIoYSwcqhWU4sxo/+WCJr5DIeDfcoGsSn5AD6F5YmG32j
CJPlZ3K94qgr0/8V7mb8Ntz7I5mlVLSgvh68OqfOYBp+clT4TktWEkfA+ENJq/GC
Wrzge9817wyJ8ByhryJ6F9OzJXb0+7h+x0bnkRiXIT6Fpz5Ujsg63DPqxYDi+bm0
8zHIx8KgMn+C2/7A4II19YpoCZdPc9W/xNotIrhqezARBfh+odmf6+ff9bp0Xrem
UWWeYvV90RM47ALnlLstKlHl8xtH8+IQIQy9wSBOzVfIEaVUIoCYCABS/2Dfe9jB
0JmBZP6G4ZXJ+p56MUXpqW/gjEumW2fViNquI47ndrosy0GovZaBshsi7BdbFBJ2
imoAP3Iw56T+QiE6hymzjTevx4FU+LEvvkl7kvEcJD63PchhUcCNEPxOvgNjqV0d
Fz+o4y/jwoQrW18WtfK2MWMCKp/QCAa9iDH+eD8zh2uP39Ps0NpYuBQVmxBSR7eq
UoHrq3m3Y43u34shq5Qb1MUnZtYY1X9HJJN8l4eaDgWPM0qSkRSHOHl7LZqL0IQS
XEnJS8k68BxL4eO9tte00+zGJpyDU1Pc0IjBW0EQEWjRc/lgEyQOyGTRHb8T3MB1
72O1N03gunzqNmvueTvGCMnTg1H8Pk68leot0lnjG3mIMeU6D4sXqhW1mWcJQ60H
8vy36ySNOY75cDcw0dWTTa5EJEdNpU2tDC+qnC0CKllAiS0aST3D8TvRLlJx8SE4
901cekkfS/g/VC8Db3m0R30tMLIurKeLtjffm4PGrgyRxoCZaWGtDBubpBM4UrQU
EZCiPgz2fmTumcZ3WfQpw/J0SH7XkdIO5tG2MTiMpo6dvAITzBfSMFNltMqxNlPD
nUxsKLusRsLqjfk1tYgzGqelob9/wzpbkwKP82r7viyNxMdJ3w7lN+jJkef6Ayc+
1ryX2+1Xwky74IRar4OelDyQrrsWo26GWk/9UOgmBVN6LhwySbPDXAXJK4QivSxi
RycKysG9znCGGJa2z6TBLof7ybAVHNHlxKuvhCv/nS0iW/1xqLuFGvmwuj5AtHhx
Xe7p+n8Ak8sw4CYEsuFf6aRfQf963kN0zvtSDyBB4gYkIBP+s4fVQcatCpaqQvbk
U3IdRaM47w2QctMkx6qjx10Af2ntmxJAVqRKKrTXgHZDGYRRD2zeurUoMfNAArPb
6GvF0LfWGnl2UrfWyLjAgIVTrkbFUzoxTTIv2303oIrg/IrlByKYwZa7DnMeD9Il
2Rf1mWNkLJ6qSu0617lv075qUomyjHzJ64w5x9FIQB7uwusqanWqqYnzGjl4upP5
GYWgkwMUC7JufJAvEo2L0/kfEyjD6C+6mpalurx3LzZ1kVmt3j4zStX+LTFYEH7k
TwLc5Uj4QII0OLi0NvhX3jOvJUZbI3hZRbtc6ZYWRIYqE+BSw3n6GBRTzJHf7F5V
l50VhZ4GaPHzIPdh8pRZt3nMvquiV+pFsC1pyOk5imYrlyjkneBLAPoswkWH4tsr
QOPxQhS1iNlczK/+MY+LNXVsiPukfYOLnE0SaAWJGGYwxXrz5Bn0GZNMIMSNmiWu
naKQLHig8wFf+v1gtlNzDZgVGUnpOtQ+jWgwQxjqIxX/hH9j3jFhS3ZGCRfQ43+t
RBUzBxJZjpusetLPeL/OWJwAXOq1ajjPmc1g+Vv23CIS+yi9zN19vpl75b3UMMDQ
YbX3tZzHGDwvkgMv/hDlzF6wBQBm4KDMooiCTSCMcp7kwocdaJcz8xC2ivxx1fFW
izq3FVrbHvo1Wfli0DK9frx8HuCO99TWl2G/TDaV+P/z3obfnSeSr4+w44Dxc2hv
eiQj3qDlkxmrXV4vzHv/+2wIEsIvjXzdjMFtTQBc5jXTcbfbonvmOe+5lSj6+X2j
1I7LK65t4EdnV+yWrhTyKtO21Pvkv6htaYVSdz6Is7oYVsHUcPyrQ2UbJXao7HG8
+SwxntYHHFKqC+oRNmXRDcPQdCsCd+6n3Fdc2MMnTrRo/h+NFlhFxUYPHE37J7R7
wvfP6XzRTzjFyqvDNp3iciYZm990PoE22OTmQ05jkZw+M66i5G4URSX9/zkoYmh7
7rqnl1gZDv1VwpG/ND1M9+DPlzmW6LhI796WuCnYgqED27+0EsnjU0scrQGinQBN
rx02JN8sOJVgpfo18Mamrqi/kf1T47fmPmp2Bx30gnibD+E9w6Wy02bOW6W733WY
+KnsyufcG2Qbfis91FjAsOgmr82Q9epFKJE1h9XisRMXg2qg8o5YAgpOLK080hNf
zNYywPu1D23/m2XYa8Vmra7CP8nCWR7uv5zfppysYQzYIRjzsQ6MUcWncTtS6g7l
qIZtiKVw3YqlopI14v6b0JDOWnyv3Vy00MfKCO8h+kH12YzSTo8xKSJ01N+AC7XO
ygt+pEMSvZRibKvWwoTnWk86OBYnBx1rNZQpRqMWDF/WXwc5tkuaeoYzNk73/HA8
vuI6jJ9C05RjO8eMfpH0kwmezZt/OKspx/1Mmf6k7Ba+ZuyBMO2AKmVuwc0KOC2q
d3bCMGyMcDciecBlA2vEZGBvCAHQ72UoVZ0uFs87Hr/pLPDcH64h8EBg/eD80ZoP
tdQNQ4slBxrRNvfyWdjeCdbFW3YLwIHsxtaL3i/CvBKP7K5ERxfGQlEs9Warv0y4
lUmZS0BaJmb865Vpzr3ZNkSBUlRPR4x0bGyRxcorPyuUll3aAlSGWgz/fttmmFej
83DbAS6v0yqL+VhCNJfysdyfzRze3U+CsOpzgpIqXMC8yyPLM72NqVhTMEjxNp6p
BEj2hUp00+jNSNEnu+1t1AAMqzgg18Awv5ccFKoqQyCa0TgBFuM0bQLZMT5zHkcS
nRaiNP9Y4gMmwZj48H69aARjccfFzVtwZrMV3kAXWwlTDsJSSwEyF8eSw3D2PM3Y
893wScqzDvaS/hv95h1vGmlI9FYkpyiDnczoRTr+lJORRBykJEwaZNUmNhMdnTjV
7FkKksomLCdC0r4kpK7ATIuLawqIR2DOMVfHD5igrIF3VJhOpPtyT6LjkzX1e+NC
LPR5KL/gcXZo3qWhrVsG1UpVxVsLk0RTUd47OyZChmbrVn5k0dIkbbqkLquyybVx
nbdyssAN9qZykOasdRthMET9R1VatpxGvJaqxJQwqwnNDWa7yykN9Dd931l5Kn/X
sk/ZJ+0UErppIvQOi/ynd4fCTpjNHFNyEG96yZPg58/InkXS5N8Y29b+HC+xb/Yt
sI0/QsaTKvu0mU4IRXY7iDmh96HB13VBu70uq8pU0p1jjjBB7JNzrmwPDkXKLSwV
FFEM17N4jTcGscYH00MrPhbJE8Z3ZEJuphAu3uqLaqzLssDy3KLGHQ2ho//7ZBA4
G83OHgHNo5zYE5Pk2i5uKLLySkRdZYUiOFdQndlEfbbWCRON3ZiP0o8Mj5ZlxP2b
qLASaRJD4wRci3TyfE2JzSeMiLlQcc37+T7TP8BbZKM7vRFbUWthegMIeg6Bel54
/8yPIEUCCX8AFqvtAIRfj+1MsQEbcClETewL3KCqdied8gcu+1l9mPnkS55jgcFe
UyZxbUyZxOx367eidgu0lPMTYsnF/EWbyNjEI5o/obea23XfVIbPWoUubHfxA5dR
urnoJecetLiiBgcU+jj9YIeULsUdhJu7GK6cW1pW0aKdtwpcGIFDvKSNuZ3b2FmA
0H/QWi42Pan3SOJVHgUKoKjdh9MZdbybUtvOHIa4d60RYSqM1W1mSQnY0ASRo+Pb
WDx6O04i3xupnp/4UkoiBnlUQxiSPhqy0ImvNmGJOHScV6NiI65HtrzDA4MDzrHT
PTbEbrWH5vBF95tEMTXxvCWqgFZVhXbWZESMQElot0WqFuDzFzhEc6uY+FxNdcq7
bbAICzpCiYX7XAr1jkilbkM+QjZzNhGr+GoDG0RnLFNiehZpv3ngU6VR6/ENqVuu
qwhUrgL92RuTH+QAGJA3HPmc03eC1OTODcHgX+dIigttYWbzFAuGkFu1hvdOA9Cj
1rI0PmToUN6sisJHSKga/e9K4HgQ8nzH5f+CRHoe45TqeQL3bOiLnTIv101uG45m
MR4T+8/B4RvgT4gG4j/H0mLHA5G2PSWhH1MTsfthwhnwhqYGpSQ+UIJ5hnvD5CIF
XoWWEzsFnwRi2OnmB5WUyS6SHuPa0zrNe4B7Bw+OK/dCfjVS0A0VAgoofoRQ9Jiy
BOfFT5Zyd34VhxA8dU9F8BMqy3HaMc2O54ivAhJgB5I0BvbdFyG2Luo0oEZS+gH3
uIe9sZ2awM7gkiNZfabJQD8PNZvs9q9GMxqh2zoe/oXF78VZibkvL6mWtQ3Ivv3I
BVb8iEbuQov9qOS9bjv4Gm8p1r0DkfBho6rmpxMeGbMyTGBTDFjcfAK3Ycn/lE12
0CdF5hyHie25F/FsfKFqrvVqhPxBUQ1ieIBlXd/2TJGtuOOmzFUJVwqhnvhIgmS0
1maZrkI04iS7HmLitmNS4eGrCGFU775PVGlX9V4ssZJPksvV2HwRnxRAl+/W1eso
b19QSNO3rfaTwfrHhTDwZR/LBG+BfEBBUN+DMEf8slxDTkHMLeTVZa5PKgFmQv68
NUE6NFsd/nVG4yekNdmVhSxGD0kqUNzs2OGOKVlmCr4lqD5azpHoEgvAEWEsywJj
gGcUhe3U/xrDQ+Y9zn7pwaMsIa0FuY71Lb19piVIkUTYm+YZ/6OU30T0wSX8sA6w
Lzuak9qbCmWtb6n+17eqWwn7k2sP2mYz5Jood6gu4P0MZOYbptjwQirrP6DrCyFG
12ZvoVMlJgZNY+j+MbWhTb9pe3g+IXLRd7AvheeObTvj7FATd4ZvxZWAer47B2R2
LcQECRWIxd2UDvI1h0Gv9TJOaFDtwACU9cNsdQphdMOjb4rUdMdyJp5w5+1WnfTs
kHT0T0OAV2/fiEhIcqwUHql9CwnSop8OM5fKqSZ5Bw/rwdOSCPh6y5fDMP/XWrm5
b7FrZqgL7tsEfbkZQaaaq6G1RlG26hvLFnN29+JQusFgjwVLzfPnTe7j5EQYTEr3
JfFEh19UUv94XmRU3ITlUp1CWqBnXp30w/p1GohT+YgwV1cijMmyQRmtTfJWCNvs
kuML2Gz/nXEwh2TBJeoysqxPj8un9SYZLS63f4+PTsvFjjfrAL717H6o1P8CIe8S
fYuyjOFiyENuwT+HgADe55lnUVKqT8Dtn86Gigkr2TZPXmLElYyhFbGqWYLbwOvk
IXtPBWIsoNfv81f5sfsXO5m5vR9j5INOlfTrcI4u5L1w+F9+JiiNir7iHs2u+Trb
/1IgUlvMS3tLqPA2o/qvbEEDlgQrcHJGv1i50t3FJnmhrUJMIu9pvvjmWPOp5CfB
vdW6Mhc73LMrccsySqYwirsmm3/4wViqWNNiDHwdYC6EFZPwHmdPIrDn46lMro1+
k+xqAR75K5rFp6/o6KWvxpb8MK6Xa2Zo8lFVqRC14SyWlTUJ7ZTqgTmJOkMikKS4
Om+M502ts9jcS3E4pY8dzk1bN5p9qMZGQzqrS+wh8YQgddLz6VbnDSIcUkTKH8r7
6G1MIEG+VfE4ZWoql2ZyNTgFSbcrkkWRn0DCQN0CiKLew4+07+fgsaSToCMTb8LZ
bKA+YgAUJfkbtXbEVkEeTQrjes5jtwDzEZe3XVmX+djmv7jhBZq5IoIMu2HKYf/k
7ktn9nbGtou07U5KsYzyXIAaK9aHcfmSjxtLjAALp0S0vaTzeBPRABvtsgeSMTk7
8Cz2I4sw6qILg7xGkNMH6AAd2SwU8gytJ7C1QN/t01PYJ79hMcoGNSS7WN8xpPTw
6Co+af2HfTRpm8qZ7O9qIT0r1TvZQTVKxFhPbLW/uG/oBzvdlonXdUDQ37EDyY+F
TyVdkrEIikHBq+H3m579v0BWfiS1pE3cBUS2rGEpPIxRmsSiUnodfKuepgM9NT84
0pJYr1MPwBtJJyE2R794AD9/YHh+AuZ29Zk0NoY7ttuw3V23tK/qRc9FblS4wyXQ
kUuE1XSzsEoB2J5NujOMytU5j5vDGi93PsA5PKHw8frAhxwmKcpFRR0UqARvDzOQ
L48Txaj1nSzCgiZdzxdCafWKK1E1DyUiYT8EsomTXKhqpel1Wi6Xw5t6Dv+WRE/d
fUf3r03cVJTE+s5m7Dw9Lp5Nx6Y2lBqBMcCcLlf6yEyQUxl6cMT3/tMKZ84fASYP
DyMJ+0+skYQHoRqoERWVvK2wiypJTx5OPp31iFUB6iBgXoX9d+5/SoJ8m8gdcunc
g1NeFT3NGhjHAdsU8fhTRQds87kZ1BvhFkfOwzgRMtKHwPW0M6s1FdiXztorXIaj
PJspwTV+H20hk0pzdx2NeOhiDdiFnyB/gYZDLxPlKo9454x1byWp93Ures1mw/2N
zbCvqiGBsP1Ye1LPkmPmn9V/063FXTNWo0+bcYqiMacHXDXf/+tEJItyxu7uEbwD
l7FVbJFF34/sQ5OudywZ/h60+NMZK65ZLZoT2diG2MCulhOpBVh/JzpwJf2DNcyw
cT+1OtHPAvTwLNUIs41q+hebx2RWaeHiJkiSMXu+DxG3u9G2l/hKCReqEoLn+M6c
u/1MtdgpGQTdoUaR5ec0lOv+Mn61wMBsgyTC40UdQusKHJC/Qp3FwWuQVkMAkNpE
2M6H5cH0kFv3bjGxikiBZ2zIbJN8WUh/r0JapVKG9hDw9One9Pd4fHbDvV9JjDPy
bftJKm2o6HXlLozqEUSk7lECkEEcekHL3Nj+FYGCPwiFI7UP0TYn9h8RfI3xRv6D
HxmEl7JbvCH9h1q3xku+rfK6NdMx9b4OLICekbWzdsebN05srNewnjCd50IzV+2I
wuNdrwDeKel21B6bRlsAdo/MC8M1+K07x/6kdAjtTyL3N1QhvyjdBp++nDgiQf7s
4R/3+U7RtZK0f17XfOn0PFzB8mOthP8A/9mWfhwB8x7EWV4f8TK6J3WkcP6RzGti
Nj4AB0SWXEEpCi5S495HXxp+yCICDETFlgPd9lYabJE2H8sr9+iN6+zvUtMkoYV1
mJCXg0PjIBrCjSOxXgxul3JGFeZBJVlxC2eToUgUjcA+BLdyDt8vYcDxjvPP72iS
I4n2qLtVWfr/4nUXAAQPdmuJbBOK+Cgvj19SD64vpCq2MuZDewvf1vsrDYdFa97f
J+p6VrvyzvorYqhewYJ21rSJREBVKe6eNU0BYxKjPKPFpNsiyJf/poqILtP+bmhJ
CRjJ/970h/RwtMfMlf/MAAJ2ldh6+uVgB5e/7zmBy0eKFliHWZCL1nZmeQiz2xNl
yGXTIRKNSswOnxya21K8DEkE61YoCo5gmbH/TZiwGhOl/PFicNg+7W/UJTOYTVBJ
w54A1nuHAwACZ2vke3cZILtB4Hm4JAO6l4uOYu0yqPgmJjRTUrHoqGYvSk37wiiI
Xm6nr1Ciwxqtbu3SStZ8C9/FuGRxkwEjcPFgrVqrx3AAtOWIwaT48lPT9VCBLF6b
YC/96xZgfiEhDGo9z1fuhjZ2pXtYEU8RVZvjlRwW88XTjowehEJvKJbSCsacexTq
W69ptH4F7n7lXJmE5BZXXygEAgT17ySyHi4z/4d8GWjFhJkitW8i3/3XnClDyaPg
PCZtF/F/j6aq5dvIxZoDoziynWMeiGABTE872Psv4PAM+j95vy4RXj4bjms/UuVc
VMdJpq5s9ErCr39ZZ2uWaoueUJKa51dAT+sEa0nl/LZz8K9AaTOwTN1lfCENYSKL
HmFHJnS8ZhGTSj13a87k0kTkh6kTCbvzilQh1Imd9UlyzaGJsQn02ub2t6J9qR06
uX9r6Hl+fIQdqs80Jzcw1usBgiskk59WPKBuZqY5bm0heo2JWDEMymLMbC19qIZ1
TTRG6v2EvPBWGsXltbMnaQNuIuzU1iMWB6dlfNO24gSASUPjXdawxJz8bywmMD4A
vLzg/vGn/Sq7tRy+YwbqsrR2EhJlf9W5fRUvpcAmzOToEblcJvM7gDarwEDUAtz5
VQTH4fBXiHUyrW9JEVEkg4QWUigecSUf4NpfUOjv9Blmp4Co8k/DwJbx3x7/swsR
zXWIEqkSYKTyu/hZpUogNgVAxE5e4mlKIMOI/sfk1J3HowG5sVFASijT58jir2Um
4kPfP2GjHkctU7GchbOwbhOoWQG/rc+dU8E0Jh7U/OzYFSIJc/PeHW5+lxkedWcG
JDvz+HU3xP05vbr/qWdY4M9v0o8gRSH0ZYy2wwZqiYwdxDOBpsBqlt9Sj/qLSY1n
CDAaNR8OYlgoLrGZ8FPp5Iuj7eK+6CQi7P11g/14HG7LvxKlSkgxwcsw65hUQVBE
k/nEaVaxshb7VZLCj550GE+LhmUkulow/Tt2V+rqs88F0hEsxWlceDBg3rmsVIsD
yx/l8xx7Ii7HK1w0BYIJ9GMadA67WsG3yJNGi8b03qvMWNiEIiw7kyTtf6En5ORJ
TNhc1FTcL4BtvEgXDSao4LhDDrD+JoNjn0epJY2dIO3E2P8scWoSH8kQ19ePA27Q
NMaVH8lRA3dPPVhwjLVzi3oJNpXVOoHSLoTGNZyM3u7mCc8bG09A8LHjxyBPcxa6
GxNlYPkua8aXme5DgpSibxnPMQXXhYJYohx6QrPKrJILIM63p1xcyvKjcUb3zDIO
vIJ6gFf3djzi78AhVMvG2zghZCEtlc+Bl5EZ4OsmckHu2qekT3kSI3MtfTtdn/Bc
XWo7nNyP1QDi+25YtfY1wNutD88dVFnCwZsMz+WTy7lvRIHDgEo7gCwP/cRPWv7+
TGkcL339Fet2YYlQpawAOX/tJ2hgcqWDiIHjNaEin+171cWv1S4EzDs6HreOaBfN
1zt49Xg6gE2rxTuqFc1iqqij0uYuWZUBk10lBEcImzQ8ZQQLuCSxq/5XJeHOb/NZ
0HgxVn/lm25qG8UHTi/x6+C+vMXSE7eC61YwA8mfinlfBlunkiJRWqwGW8FmvtIa
dfyZyWuX/4QJsYh4EYjqftnrp/zgAXy3uc4KYdzx3lrMg+TkcJFHLZ+uGzeHQQzY
ZzfkQTGddgDXkY0P6QocB5NKKLQ8CKP4kLX1jsGrA1ASpj9a/qRF1ux3dfuqm0Ij
9RaAA7WqQ5kg0lMlmWXtISPFMyalXjQpXHKFQ36XVcTZeZaSsMvnZQKyKDqN2u40
lU4X4AsDekiE8Qq2fz0uZZ+QJuAvFVaLjvoReULh2vxyUwc6O16bDarVaPzbDRJW
XXvbgPCOo1F+Qww8MSqX/r5FtJf77mYpe0PqqN1QDToYxHNXEka3jdVOiseZ2jpR
kXdKGwS3xvUmmARQOrlYBXky6xQtX3BMfeKHIs9T5xXHQLkvWTA3/HVbFH8XAuuI
lxvMn7W9Z9g9aD128yv9aknDmas31ss7dR94NUA/uDihO3Gf/3otOYf3WJquF7Pn
5LsjjKCziAJtBhmOtrzx7iu0WS8v9ZJczI4bmWOZ3s9F2IBoh4glRVW6h5f4QrdF
YTJO7L/J7+rw2loLql3/UDQ2n4jMREBnFEUYlt1uHp3atYaX/hs3S62/GO/F1WPp
4D66NxNBxj5+x82apG3zdRFv8F04tucF8eivm7FLowy+f7XeOW7MaVKxS0PoFTjn
H3t49M8SF8gdPM6nZT5UbMzkQ34eyVkJWAlSJUt+MOaNoH9qn3tEDohcN2m4KICV
3g6br/qYcV96Rtyqo1a8yg0gmFqQiX303uHs9o85QVsiMBn9n43ad99oIuoq1QfZ
dvYWCa33anBxs3r+ZyizaV2t6ofBrFQ549R+/l9eeE9hkIB/rrYTIOMcTB4qNW9w
0pcN+y8h3Y1HHqg564eY9GLsy6KW7s2yjCQXC66/Zr95BpcwBYpQ1+bXGtVchJUQ
iOBiFxETGpxOSOVCDITqHloe2VxEtF8MlqkBZ8qGUx6hTgO6aObmxmH0K9Sg+ENR
8WyTmMMXPIdlBaax+01oJqR2TMH5iKND5+h0a+fM6eVqDK0FR76VSY0NUfd7glqN
aMtcTwO/C01jeNPUZPBTh24CZ+atJSHG8cRQmqJMjPsWgwobVsUhJ//yxsuEtUa8
xKOKE6Y7cqopn/tKmTZWFftT9YcML98E3LxwQJFoJ6XscG5NsmSKKs5kQqJ8w7AQ
a9CU/IASnGI5heb+s8cqF2l5pyQ8xRlyK/yoaeROBpZXx/vvAHBV1ergf3n5puYO
tvy213GxkT4LXZFUute5ZDrlv+vLIpGTw9p0h+P5c5hQnnOpAuX9HNGv5mKX8739
K+wb7N8PFkbB8/9YARXfZAwDXills4Tkd2HDtgyIK66j0UzrzVSNa+GZDZlQBOTY
NN8eamCS1XmExYAsPGDKJJPmPWMuqPP+vRKhvgasd7WNQQAzfY0WjH+Cf3KUg396
cs9ccNWzBMqH7I5jHhkY1y8KSIVdmu15J7fU74c87lRDhkoPfzcfiZwpKkXZovMa
3UbOCGpOzVbrF0PJr4VcbtIQDkBl1fHY+rn1zofEAtWUTZ0gDaGwvi5EMD/MjgJQ
tvO2uzD3x4ANCaLTn5Sknm9VLFZ1HR18ILm/KNsuRBCz+SZ28vXCSPrWxr+WOAyU
Sfu3RPUK1p9/ZvdCUyP9bqCGUxr+Wi+OssX3kpnpO0NMDCULRyoPpN5dEp181lJB
YB0V4GgDTCEMchdlf5A0F3udKGMp9I2PseSpotm0oW5yVldC5OPDl/vUivwLeWjF
QrLPsteiw4eVEo5ADjI3i5yb+plfeu2WKCUMOplvvKrl27qcj+0tuE6SEYWmiyop
OdQsl6Zb/nj1xpjkADoLad0ywgxi6piK0CBnM8q9HZtjtmVYkv3j7gaSpanjxAI5
DQHXTL8PTiDScLS0ykUFRZzwS4LqH5voeHCiRI7x7cZT+bRNXXsPtZJVZQfyygxU
ex+TDGDNBGuZ4L7WXzOz8SlRBTQTKWpAUTDzpN7QjrLGnc94rQWcHeyb0XF1DOSx
YMcDzGQAI8cAneRlDOn3B/Y3NW6gh0qHXUXZbVgCdS4itdC5zQuicUyTG9GXtu6J
9IvRWK2he36af8taKTBh5BqRvNONCLYUOnrrjnKFSAzEkX0R72jtsuQIURR3TBAN
Nr+oGQ2OoE/W08FF7kyIzTmnx5w2tIfG2u2g1BZMDEw9M8HmCBoIfFL8O0/CLha3
42ECZn0htwoeJPMx07SsQ548LBrUkLp4WCu4d+KYNueMn168yxV5yEtZBJdWWJUS
gd1m42rHCpIqo4orHxZeYsEfLhtPMlE7kxZtO8zIebNdi3mbdcUk1hc9H/m/hcjK
np2cQkoK9bZauY700ko7goy3pqSyNza3KSueIcIO7u9Cs3qbQBoggD9V0IZB7b8O
B+fGcCm1vQPUkksagMnmlyRcb/upb3JgH4BAtW89DV7Y67e6h6O7JFYlUehj0/r9
Vv/0F23OYRC9R5+1y2bAbmQPVExJ8DPqf6SAC15PMobrJd+RQhAJc0jW9Sj5ASPx
ijPy+PbOuTuHFvlp0E2uPulxrqy3T7mMnvUZorZW3+LzzP3UahTMqxVxZZ8ejKoT
bxJPTQgFd5qz+YvwOPXGe6AUAb+MQ2r5b1TA4rg3FM1LyUML1frlIvAhvEsJYhuo
sZAvVfDWlQWM51eW5c96uEcRuQlpnZnqvDQtcc5xhU2UEDCVdPorIvB+LCuOl6Ag
xGd6tYQ7TSzxuRvmDLGBUpDK8Ufm7n5Yt5sl7ft/qXh2PMh6kVDJK21r/+NsuSYk
/o1FKryma/QbidPYgnCrRmFG8/AAcRbuOO2Yve2KrxNVrDBM88yMq6ocbBgiJkdI
tEcybzuq3IVrQeepfVP0DrnKf5ie2KlpcTcbxNIIxBZcwoVSh6BymfpCzr/kVKtF
oVJZB+V7Uo9VvQKJd0NRu+wBzGsRUGgJstKmb/+B+7YoTJDAh+r5TO/wBuJkelbW
50JjVU5Z9DkNQzGMZRZtfZS5s8mYnWhz0BsTAGgLiEQGRwp/gkUgUXz8QQqgKGi0
Svibq0uGvZ3ZGScdin2whegX9FoRJGasEJpraTJjqqGW86Oi8/UTkLPXpQTuAuoD
x2IG+Uop+7Fjv4VoVYf1hDYt39TYZidS28FOOVbYEKTCagBUqb5ShxmOnABG2XR5
wTYSBsvC1U56q1L3IyA7pl6SaaFl8sCF1eYEJ2fQjwI7v75d0/6bOtgj+nf2aFot
bQQ+b+WJaJ0wn/3Gl8Br0/WsIFm9EzWrsbgVlYnVMwclnXKKYooQZA4dE/Rl4ELV
B6WKQIUgZTS0fQqjxRQaZrBa6I/48SGnHAZHUtV7mGqm6WF9j0xDd89WA5cRLDWk
i9HrQ/B8nfaYCC3F8WAspOHyzA5NQzkEECRFnSYh5+ln9ko2j4nO4aFnB9WGRw+E
F2IrUlyBRItHR3Z03tpilA+i++pU7eL9SowKveMY1YK0GGvG5cSrqwARfU6pZA6i
/dDIxsgiTWOwzBHTt86n2cvDWDwG/oD752f4Xrib48CqFAUotd/6E8glg7puVLM6
fR/9RgoM4UPBN1jXaWazdCr7gT1l/Etuu/BOcK+J7ezbSZX6RkkpnC0G9lx0BwtL
jF4ls59JESbdZ6IqUIkQ8FmI23t0oLjGCs6OdzgXE1fYQZ/DRrtYtjjM3yLQ4wOl
yC8XAjPDPwURz/xi/SjL5hf0cZ0rbd7xHAhuv/OGBfrExnncGXPnx2BCA+ITFFbK
58XYxdVCyTVzerGr0XQeUxgiMGKNYenPX9KGdkNlkvn8y5dcfJ6XNySY0nodc4oc
6X6eWIp/lqu1Qv/JQU3EoZDCZPK+Vs0jzEM8OwTWUm5eAoSCSr9yNzUOqNencJcp
u9kMJMZSZuJeMlf7NYb6W1f8fFg69K094SVyPTbYaBM/8Tlv82z0VrJ/R+Hq9uUq
mss9ITt2fJKcB0y7wNHrR90GE4eAIMs+1sbGpqKoeUQSteIAS6rWn1lC+Ifla0zs
higtcmOjLAYuwYN2WYerzsKZxGvvx8OuXQkxSaAOatbptTGYA8vNVvFJaZxn0Xfx
2KFo5rzmSH3Qcc7CnX2QasZidFXUsf/G2Uei5l/bu9+1SPGiIGPBf0xnRC3T1ql0
/gmOXW8P8NbR9azq81MuWAfKTjSjAEqS6H1Thyc9VTTWw4cAWa957G8Btc8rtGqy
9L6W0bbRlRBh2BOyWxEbaXhcEJZkbdxBkzgrFdY2dfaG2fgg0D0YM5Rz542C03S5
ezYH5rw0Vh8+nfRmtdlW2JUSALsiffR1/bUkOGe4sR5v2xhOzS+x/xH+EMN/AnF7
y9obhSQE7aF8SKwQMsSOP+/jxBPM7V/heAPLmVejHUSH5ruSdKE5RiKx6vTw+BMs
iChJR/iwFAfAzy+nOr/wNqcHCKAyeiwiGFamfPBHtQpLpYfQkTdqbCQ5ZdwRxOyN
CxpkhGwrN2wzZZ0n6GsHqEER/u10wMqjhsK3CpcsBUz7sjFewi1IOlIrOdeL+OSF
2mjjeBqyhvS6v5TUHtTdArdk8i/NMXWOYELiy+MWCKyqGPsi/pYtBe4B+bPPtZEf
xdnDQ1IzWJP4ZhVYHzQlnr0loxiNYYZ6np+VS462qI9mcTxdiKxtJVoq2e/z+rKt
wb736yelMHyTMFRFnHzXkLJb0f2bpt6ATFIFB8TC3e653p89F4YP1M6Q14OWo5bU
lkrwsN1nAi6RnzHtKS2o9EVuJstOZ9Mdfh0j4lNyMn9fBeYEtn8Vk9bP8i3V5RqN
qQ/c7mAeFYygdQ6YYm4d0Nc9jaQGCRe7gbgh3d+s8oivdHmt3PA+fvyMKw9XgDuY
8vAa1Pa+iC9IMSA15KwzEuGMyCVNFSJ8hV4KRJhJtcr6ENkzBb57fDx2+/X4bB1u
dsN4/A1CKfPYdmre1aEe+iYsUNgpdlKivtcAKy/UBpGIlLH7CkkbJDz+HN16X7Zd
efI4PBArbiSA0Dl4kE/NJZVIQJqbQOZDnSsveNlTXWFaG0ttjR8ULcBHvJbB52ED
feqEHKwC2kfnOo8+Fu3wfJafoSfovUrDQCtxGP7xG8E6L7km/0MnYcRmSEAvKKWz
OxgfPNrD1CvaAtjhru6mCoDf75akjuc/uAiALLT25XITHOH7L5YMtZI8RpuyZGRL
EHeUnnafyB50E/9YLXyuAMYs6E90mbha/Bz/Xht756fgk6Y/yyczPaPBNqiAc8Qo
6Niis6scxVPo+KnMUntgqH6OiH2dg3o2pAYYf4alDJQSQotkyWEYyejxRjydhGHz
Q3ZstML/zVztUFf9TgDYJQv7TN943VCSWyXEG8C/ooS10MKHlJbFks6LSHaeBmP3
nqJRQsF/iHdTFshWjHbTWEear/vzaYDBPSkTta+x6YHqcgCjjzMEuJpIEFibUthO
Gc0kTl/PZ18/c61tIUHSf7iKi63krEpjw2DgybJp0q05v4lvXWNw67dbL7D47gZf
9EF2IRDlrGhe9mOzOY63s4NC6dYkygmG/zlB2wuWVI0cJtijYv22Gb1rfCnDi7u6
v1qa3gGr4Z3cCGK/upebAo/tnA3H/cg/VkkfNCONs9xLuoNeGJtJfSWItzSkZpP+
g3NaIzTu9MXbN15pxeP+Yr/sUzffRSlRupiOhC0FBTzeBg+ergoaVuoHDKw2xTt3
WTGifEV3nr6BfbQmE7VsaDlXoQMDfftrNm/O6RIEm3p0Mqys8Xyv/Jslz9HnBVSt
h6lEqDZ7ybOYnsEQ77xRxtcRp2aR34qtC8k/xqvW/9KXYiA4A5bfWJGaHSRFn3yp
nTYWUERE65/75DcFZfEREJDbq+BPllrJkLjJeXOs0YlgRqhHPBvm5VQ4BRTVEI/E
U1jYf+jHWgJokY0Oyn/9HueCdQfcNzW8e9YsKK2XSehilYS/cZ2np0zSIi0v0MuJ
c8lUKOf8ltDHqao5TvTkd69PZUVEta+cIN3hTU8G/J1s2fViC3DnHSlx6pcI1lDB
tMquJO1qSV4WLAbwTkUUusZnRdBcDuRLyuanO0NJEV/DaEMBVOanOPbA6sSNHMM4
1oJ2Zu278ptcLA/2YqXsbg3NmJoN6my5tNoO7pWn/rdx0gPPgQZO3GPxcjwvcy2y
eIr0Yxys2Z19SdbCR1Sm1WXV2Y88GbJR6aa8d7gyHhBNTxDsMBqTbjABnKRTX0NC
mrUkvm9NIv2f6w/Z8GnMALYWfFl57A8LYFdGiWB4C+N54r8Fn/6jWgGza8WHGHOQ
SdI+j33Jvc5/W7G+M8QcoI3XMHKtFMeRnSZvzcKUyhL43r1SfM8igQRvhUqQY4dJ
hTlBjIEd2NYMrC1C+a5hXAq0Vl8/OxO0XVrYIoGwkI7okFbBg6kzueUlkb5op27g
iroS51Hdo956bPHB1E1nkjmmTIVUcc7lwhcH+/TPN4SmoLoh+//LNXVbiQAbw46y
lpR2ApcvdyX/qccH/4VqZ32bKKoK4e1HZas1EE7AsC4QuDcQ3oVeqZDQ1Tdkatc0
S611/xuLPnnhKf/2GXJylMf6o5pdXkzhjYWqzfSOBy9CF5I7Ek+cGPry7GFD0p84
0YuDG+L5rUKaxZxfVno/XZG782kL+5tq4DReMQHYTjeveSb4iJ+CYMLi5f+TBs7E
4kDsWZzQ16dxVx7Alvu+Jy3CWABM08v8CuREhWqtKbjX1drkmOHHH3RtXg3cjJEN
knHuSpahMBs3EVA00DSqdeJ0btAPz1LbIB374Pfgr4FE68ghsxX1pUaSWZrn/TMn
hvXK6RK48EpbAjYqkr8MbrrxB472zUx/WvDk52VpISEzcYwn4GgwdLXOVcDTTbpN
Rvha2OzOfQ1ug5Rk+jad2hRqWhid/9Xq4EZRlSMA9I0fgWM4FJTCMaebegZtTOMh
kEAd+1NMPc83wjgylx1rfhbRWKeS+0D3rlzUk2DUVrqv8ZsTm0Lx+rjEkIXU3j6V
3fpvkWsxX+z+Aa8jsDiQyarvENR2Qm1SOZfijeIWVfjQNsEzvoLjcuxWqzLkqBZB
7+bTZU4i7fej/kwu4M9ho63LGFPxrsychvjaOBESLDo1W8U1CPColiSkOGOn/DE8
AzxwaE1HHjzZvc8l1r4JQbalFfVtKTRYr7IyxUARXBlENuOnyemdi3VF8ysoKejj
l4XYzmsS2KDNCDLy9ROEUtBMdHbN23zloShfI63xBtDvjYL3a8VfAYv5jbkCwpkC
Y041WNU44QEboMrdU1/BDB1z/C3GvjaQy1wN2SPH8Uap0XcacLgLgLzE9lvLiexf
cyESpwWLtQZAC8ZHqzohTv7qk+oTGoAzhWHH7BqpCpudwJgSOMgkbxK48KkQVk9f
zQlym7bS1szS3251Pm4iLMJx7zrr5195GUhesUO3R+xtQ/NkblzuuhMMHlj4e8Xb
GWqsF7JccqYKOE5C/17zHUqVqdAk5d2Y/9MNGvjDrGwFy96r9N1SALddVVpVFv/b
D0CGzmOVeKtDvUutvdRK/06gHHDdxJrx2Mz4cVPhxmYl4BZCm1T/OBqWGG1KiFpu
MtVR/eLwwmrIJ85rKAiSjNI6aN9xzoI/QWW6wj0ebmPdQklaMNDCMwYJ7v3o6qqn
FpU6LBmMY/8ZCA2TFEoeP2c0VsJ5v3p2Mbl2yeXpOQk352TfSn6TvfVR0o+JS46L
KZN9RNS145r1qEoIeGxJwDKocAPOHC0T7P9ehuJnSi6gFKGZB2ocv1ETRScECjh7
+MiwFCrPAbxHcvw2J56VYNu147MKu036b5O5r/JD3N5oVfBcz45lIUEHh7Sl3pQ0
gBCH60U/uCWh+yEyYJ3B8DYgrsYCIiKjDiZzuDHaAJ0SnvdCB08aH2aQY4NZRB3f
JVyvSVQzQODQl5FcyvG9yBI5nLGbkYf4/+HSPhOpak8E9DWw1GJMQ5tim1yNYx0E
Ys8gm/1fdK+x/sUO88OGNGGFJ1Dp3rS+FbxvXjOSe80yiPzpA4CqJ097s6bqQfud
FeFMY8NRLYlxVhVD8b0qnnQXMdN/AyMYBw2tkpKa87hZdM+r5DBMUw3nmxqB50g6
neJt5/uLGk1X4k/D2ghdUYwK/q83nL97QMp6Yl1lKhThFt8xoa+XRdREjsUk9B+W
LcyEU8nedqNsP+CRwJvUo0sbs9FwogHdZJ92s7+9pS5kMtt9ZrYxpmFZHKvFhtq4
fJzkT595LSUZVXjxfPf81dGwAi1azWJPcJVaLVIhcMBai3tKbwyX4sRO+Ia6wYr+
QzALgQ/y9KGqvKjDbRWyxDLbytkEJcCvMwKrENdku83GpSXbAkGb/FMOS86tJpBO
AIuRkcgVidvWQBmTKXzr5VtBDXM2iaj4z96xhXm5aACbW12MPSVfsLtvmuP7IkIw
tjGYHJVPMcv2U0fsbkh4aIgEyzipoi5vGww14ZFqc+tdgKjVqzbYUY0OS6nq9vp5
gRZd7Dx3qC2YUEw+fr53RFgYO7LSizyMiULDifnjsrhEEx3wsXD4js8pDRpGv4S+
dgA8nM0YNPrc8guL44LSJ1XJYe1nxSljzrID0CEjqHlV+6BLcN/oIWnF06OqXFlP
CKZi07P3kWwhKV6cHWApYOp17NwSGLe6lpLPmCUBxzhR++SIjknxXj729pAB4t2s
1wmKs58ZYf5DPAvmUPiKelQbVhhco7J+tjUqIhFYUONwxJxnnYPQyS0Cu8F+7hhk
y1RLxk0Ag3xPoExgtn0107xh0IB2YzNpADVaOkPd82VLxBqnsNerefa+14rPO5Me
ID8GxYqgn7bAjUMdpNmstLqqj34fZmg+eqoe+477l8C5auUeDgBEbImdYnsYHFhu
53U4coxNkBltKofaRjiAsZq7pM/6ot90sk2t3Oo6iRcYake052TEGooA7kWySSiq
XiQxIj1n5jdlL9WRDipPiXiF2Q2Pp6Vk24T8M1kBx+FEt71t727bP8Cnrk/j75Bd
GH5SS/bDxY5ZsQMPkHMvjT3VBoCVXsUsB+5q6n4HrTKywx9hOg9kJAMcFyOuKS2l
J30XpvHXszwHv8VmTdRQO86QWoCBUKi4FWGy6n61E6E1rJQRxDiYHxTupLei85bP
BFOy+vjmOfCu8HrVat7NwmzcQw2RBLIl8BH1Jq6UplLomZrbLU8/J1dJ2gv+sQ8U
zNinVbVMxwKoK4jCfU6j1PyJPiJGXDVm6jfszchMeREEnys7u7YwHjQwNEhZB/4z
Vpa8Vrnfrf/lrM8ONORqADYsKHJuozDGn1ByxBhssu5IjSM/1inKj11s9L5EKmsv
ZOCco32LnIDNwOhxL49X0lbnufErqT4YDDcWVktWkVgfNaS4ci6HUrBWrBAjfVS8
m2KfpKWYNsvYTQ8suNenQ1rbIdHQhV5/3+9bKgOxOUyN9LEp3WDIvUrmDG6WYPwv
wo3CQAd1b4VEcoTWTvQKpksty23AaUPX7X94F8yfP9rGA9+6JCToHXD4ZD+D+G6m
vIYGpegGRftYG3UNazG4NefKN8FQAUMuKGmy1czxBcWvgfeAOaLbchC/mGfVQhA2
MxSLYNQpQR9XsDsCxD1Ne7NBnwvCr+1ZikpWX+dXU5X90IJ2xtlw5OcQ61Si5gaP
gDAk5C1LFYOVR0VmrXfi5OCEkcS/iDh2gtWTkuJlpNNjKDhOvCjkiU0skrz5NxNR
4D4coe8a4Ed3mJiwR4hyiIlxxPdKsF7UM/wFqTP1pohwS8wIWL4U0X0IbnuBWiuV
mN9GBictDnRkNipEXfYEtRV8D3Kh5N4h3vRIMzgBphIv3FJrgHqSIwY9x9RJHhm6
J7cVDJ+b6f0TpiA9vlbMz87ue5OxCRcmkNl1/krAt0TyD0c4UUMttkjwgq4HBZSQ
zjgFJQ717eob+sTTNcPMrlmCpMu8/sxfCAX0rlqChuvvlRtG/5obXguBLYdZNrRk
iltmL7sLEsqoWxhJnlprReNDG+NHMvL3Rq549QDWSID6tKpruckM8wW0rvn5dI0l
g/Eoo/Aeu7sZ2FiehbWfZ28QjCttWkO8E4JyOXJSHeAMrbBMYoXCGzGpSp9PRJ+g
IkglOC9Ae0UOxTIAIdjca5oxO5FsEjAnwMgqch4kK3bpvk9Ej4+uomeDqgvRNqcH
Btu7VjuHUQPigSqoKJ/3CAGu93NLvyg453e8k4tIoM7EtSpO1j3ktTVyTnqZrjtP
9Ln23N1pE9KsiwNkN1EubCCiDdFQsfEfX+CS1MKLyHb7rjLsPM3UsslOfF+zyAhn
KpzTkFNiSIHPXp2L9e+rd2FiS5DmmUXrsXypIckoEXvi9rHq8vzwFleOAdtVQ49j
Ggtn0C2b9WI95lqdegv1zAzQOS1MI5HQCHN2b2EYD7gVwllz9TLbZqCjFeJ5grP+
PA8AFF82Zt7Tmi3M6l6wW7AGRap7HsZN/+S8CXAnHjCmDMfkR2hK4oSJzUkl/24j
8gXOn37npfWr1nmy6cGjXmHS8RAintFuSGWE2fr82JchBu6nJiUbA42SrN4Tb/oI
2w+a2PMH1LQlcwbxo1tb+YoymBluaoTPI32Ir+6Afli7+Xwy3+4R374algyn0H6y
QuJXRTP/6vjWioRXuEksxpzo9R7vrjYqnRYgEfIQfkffTucjfFc+UjBhl8h2RIl7
cZBgeJRo4zD/7SRfshoJfg5ESKIoCqJbaHxA6RbDmTOPIS3BDU5YsvGjYvsBcRGp
S68c44Ptnr7Anu2E4MixVEb8jIdt/Up37O/PWqcN/gjDrJ2w6oc06dGqFhG4joMj
W3btUcZdcevX/mR62fVL5VK3vGK7dyjKfE8sAlseZgH3rDzbswjlHNq0xH6/l16D
snu1rs4aFF+t9O4ANSeCaHlg/zxFZNAshwul7kUvQ/+EE51tyZzh6skPt3XkBGgj
tKV9dmiQjvo2d7qYhrAQFqU2kMfV/tWHtABu2weP+V+BKdfr56nCTBYTk9gf5Ksi
aFCPAc7K6wpsfTJK0hY+R7CnUFOzX0TBVa6fy6t3Bb50+8keKUnXATw+I8gI1Cbx
X5rqUg39yUSZyHnBSn4pBOzZk+fKlpCT1ucOtA6yNIPcwJmEawme+B9r86tg1UJ1
0nJOgdLc+JOlmdnpiwdhJ23dQs8rI7GdmmZzJFRbwp+6MriSeW3DsMAMxyYcR5F2
90cuadSyc5/xnZJ6tu4GFXXsNUzTDzvjzEvdp2KzM8zaATmS8gydPiuNPSF81dvC
RvqcS4CI7VBOpPYpndplFz0ZRL52b746Kylz6W4QCcs1N4iWbluMZ0j4dFXo3fEd
W4GFpQc0LAoIVe/HPuZYm6InpIvbk/XXXFqsu3idDlotyAe1aFHAcVZou2aQWmIf
k91hIjA2KDxo1opDagRLRJRzXvVGwR3CmO4hP8aqfaFSk6U8Rucpf1YumcARlLy0
A6DKSxyABg+bs/0tubM1Sb6W8q13Ih8oThu25ROK94QXrevw+l0D/vx0fdRmTMlz
jGODundnjAwLRCyw3OpZEqee4FHt0F+G9Khu6Oq8bPfTWW0L2i8g4kOlinYY6yTp
ndIbHGZojqEDOI9eLz/DGn49gMP5OX6acPS8q1Am61Izvn1thkltlA/WWOEWzCrY
saKp9ZI3/+gl0/xqAW4hM4WDI7yGWn4DpA6yOzSlRrahoYU7S76v2C/06zKAYgS/
wLY8OSXVFAN+0avzfWQLj3w2kPQJxOSlKWwgDAlLi0fVepsWCw1VnfsfqKfXhxoA
3U9APOstKtR7LHxAb7al826mAUAsRbgYRiOAGVvX+GZuEh4DJnQ7rjuJcHHwESZv
6QdKZBe9ps6+mE+1HmnL+7rcEgoXgSk2HXpCVRtSUgutjL8hyJIPMXCKTq2Nc0Po
CgSntf2trrx76HM7uOmAhiS3R9wC3tRitpCVzIJuYo8oNNdF7InXBN83wnraebLx
OrbheIzJsWpdRLAOcufd/gj21AMXqv4va8O/8Kr9bvH9dFB6FH8axSt7LlMKe3CW
/6ytNpLKk+mg2zuK0H2Z6prN4Bb5SlNY8+f5rgXZTLGVQfu676Sxv/HK89UoRGdw
k/vuoz56M273rFg7pcE2RZxL5nO2gwTWtC1riBEY7c69xj+wUghKhPFH2/HERgBz
8Le0Mqh0sHZQZR+rUnt8M/iWWE8omobexgURuT4YIZCj2O13VkRkqmnV1cop/W1V
NhTeFXmoaXlVa/f7XNZqWTRVH/INN9JiZQYGplbg7U9txk0U+QdsnIIKYGHF02kt
atqzIFAHDmIkS99ZPqQmuvZOHu4qt2H1AkrPNxbbUOJcyZ4g8hdTZhf74ucjh2fl
vuX4YrRZCPiWx1McZSzcT6icdq4qbRyxuVziyK3bMAzpZxZH5szHXnpyazKX/mIx
LbZMHNU4mmN9AwYh7Y8YePiLE9s0aJoErA2WdlJ0KBSXypVN1VatMGd6+Ukecz/h
BIINlM0FA00pvYv2phKYYHyVdgn0/LIU12yf1PGcq3VorfqQkAjX07/Rfh/yY3S0
qEWBP/tUS3pFGmr1U8fMd1scpOd7pfcoWDufK3zsd0KEucFFNAgNNB+t15tv5PJh
MmTy0XXb9QJo4+/5SkYgXuXRPGYwXZY3BC9Qv0EqMotrNRGJ8bnmDIp1srrT0KRb
7xw5IAhKXUmTPY5rFW/CZpaP1ZPjOGOxrWNZFUcU54cvjr9HIe0x0NBCrMDAFH3P
qR2ST9sHBkgc9Vl5Q+zBS6x9VVLfIEScIvZMHz9u6y83lvdst/3F09Mx8giz93sG
FtKStrnWGcIyx11tWps+sgbOkueKmLft8QAK/w4k9HoqY0p1emobptSreSKr8TaQ
Dd2BKO8iaW8K6RS0n1m41kfqNavZlsghjadEzkpGPaaVM2ePRgm64bx8/ZEOMCTU
2JNxmqhDWD+s1Q63pjL/8RrRRCdnXqybLHS+XPmPEAfNlLtOn4O7ll1htvEnXEuR
ExYZgiONUnbjyRzxj04C8R7X2EAg1R4oYTstau3DqMfjZVuH6AvRbAXTe8BACj0Y
YL0v7Bst1pnMaLzDdjCgB2J0VNIbw41D4AQrRm0DvSet7fXuRwBe8uMVjsRe7TBK
uT3TFxYOe2/kO50661OWxBaDWoJIHsPApBpwp01bU9gM2R/H3Livnowf8njbGi5X
BHNHz5KAcoEdLkj4Rdu3aaTU1KgFoiKp40X4hJaIW6MxUeZ72TR9xCcYBx8EhA+5
+VpzegsIz3KZCJ4EPjhl4pIbCKlVP/g/BaMW3BMCuMcQgj2hsSTe6bVARj9ctVSw
7z2Tfty5cUeOhIoN5hLwtFOQ7DkfQ4ymArlkAhv+h2juF709Sm7usLMfJLnJTjXW
/DPwqcCDANXsb2A4R0X8sXxBspf9gjhbOAufR9AG1mjhS2Z8wHeA7nLoSJLjXoIV
McPfYpFRkXOB3eNhuPDMg7FJlkhSSIjmHHPdJNe390mTrkpvA6BR2342xU5sW7zp
CO/t9qw4RVAMLXChDVanaOqaPEUNs3zBWXHJWX/bXFirc+O/m7Szxw4mC6nFSd2v
Fifq6jbHCvtlSpaPUrIzzVuT7LZaVZ4DdULSD7O8hG20aRXuGKHjsNKvqEFHkFO0
rn/8dGBk/RefjXdX27msxoPX31O2odetXlec1/Ey7FphkYBEF/24h1hNVAfzHSVb
akxwAGSsZW6s+MoBjD/oj3FJmQpfgYK0MGFTs7VLsq3z/IacO2ELHDdP7aucWOhD
45ilRkNU6hoK4u4/CiKAEVSepNv6CzNHjYtW6aW8Zw/8q5zi9QXVc6n57eM21WL6
8KPE1OTusIAseFX0xQ2aNZufPJp6PtDc03vSWizNeIop4laV6qZ6gbHZbsRGk9Ig
a7TkXlSsOIy7ABIR3F1O3f164WOFwIa7VsMQ4vUg73eWjhQksWndjoF9YquNdhG2
dULyyp5zl9SuKZXpomKTItNNyOEz48qUG6cfoVxFM3asTcn7M44zNStTXE6RrW3o
PP0gSz9eybKTWbOCRsXtFZiy1ajWraLvoKiXf8Ecr8pTf4xGUIvP3KZ3sC8cuYNR
SWslS6+9OmlhMpmA+dwo5229Df4FiBVb4NiZ8FZv5i/F31Hx2NEn2TlUjYvcuvxU
D5NsFThVvHl51EniBqKUxXX4OUp6vKP2Antc0e5NGzoCj3H3DyBkjyk7PAXktsq8
9SX9w75O4GuCrBoHLDllFxt+ZZK6pNo5iBp4VBQROtinHdS824WqC9ckc9GruVEm
tJr/COKGe08trIt594xoCQErLP83BCmacFrhsM0PhPEy82KE/8WS3okcKiBMTZMj
HdZbO+jqAlqqvQ0PFX2q2Pko9v3wSDD1xFtlnQt0/HM0hhXRwOdRHPbjrD7UZD9W
cGfxEni1ap5VVSMnm/UK01GwVKiGN46xr6ULGVLwkx3pYFEYKKuQi3PEmQmXgSLO
IsOMCEjpjhaU6M2pGZPEPnlSVF4bvbywlZ5fcsjmZvlMZki8MHkGRyoqheAPDF7K
+9CnFyb0RNB2zTew5KAgAGU19aeTSSUkIALv5ShORN1vmcUW+wfRM1Il40s0TzUM
iZkdFeKkySfAjWY6tNj1k1N7nXq0pjn8A2WTacXI8aU+W76Vz8X3ugPZJ2MwWl7j
OMQfuRvvy1iSwQyMZYuWP2sZMpEfr53Aflh23dWJNuDGVxW8o3ky1yXgneAqlsbQ
DW5PvoCabcDJnd2nUDfiVv5yFWK9rfeZDf68BnjGtPvL5YuNXv9Yq73yhyTI38sl
wIcFeSm0NJUdtTdCgw+ylKNUAQ4hU2QUrzO4BK2uu8zGUMCxzMlD5pRjYF/CVIQG
XjMsQiwqySzRJgj5AawJj/eAklVX+U9IjnqZhkt8RweVwZVFMfqNfoFfFRwNNSwd
N3vGk8pDO7/rhx690cSJfPess4P1Dfuaj14DgE+bsvUif+bmBbkP0NdaCCgTCHvF
SwUSrDWp064GH6MSXuhmY/uGNzZHt1FzjeSe5GbN7SUMqdNKw1k7z3bmyS4RzkZ6
0wVZU1SnaJ0aVBGS1oK3nbn1wPIuJwj8fNtAQ3Iqjqc3gNN/ngeksNvsTMBjfYu2
YsEfN5LAxOvl8QIYsjjBokW3IE9zXyQ9NMvFPn7gsR5SO0xeJg7gWjBcR71LMBY/
wIxHB/3SBHczsH1AjprJohKzZXVvFkBud3chrbkpUPJF3u7S47Z/3ZW2wbUaBTdP
HwCyi/w/4DOrneQKI6ypqwiH1RIU/sfMk5AVfu7N0hGKtBVzMXXoRRDydWvNTJaj
EYEkc3o0C02vzvsWeBDlbRsxurzCnNXIsiClfz53uH/sebsuYJ6x+oE2RRVsRXv4
4C8ey6u8f3KNRUWuqBPhp2praxCG4oJDXYv5tOhCNKMj4N3F9kJVio/wJQ3I2oO2
K5uc6XRjVhKZEGiO9SattxGykvPsNJF73hmV5VSPR5X6hwNUGyOHYldnKjnLNfBr
G7lp1Xj6d8PyHPjxSTRtzoX3lXQjUgJfH6p55wC1gISRyhBG/c4/+l0qMQ/Dt+A2
FtRKmHIKzGO2WLMuKQ8b2veTIMTZRQ2g9qlSz3T9ATCXIUpCCtCCvo5dl2sMwg/X
NKX65x/z1ipgX+ZX9NN76oQGnoCjJ/3+ibX9J7pUg75H3NOXtMF0EhXcWcww9v8Z
7kthq6DfwYqujiPw/0cu76Yphtkm6y7ZRI5ABSmxE7YwHjGRZYsp7neKXZguF4xn
TAZ3NdXMd79u2eqgEy+9s6cHh66qGC+jQqF4LFq8L6L5XhEf+dRflPbgelnXDhMr
HF/d89qh9gZOXI9/EUKdOrr6NAiTdpHggCb6SMfTSnbwdIzWT+rWhkWVN7cWXnuR
pRODWlWnS8WnQqDN03+j6S2uxMcHZKV5nyRsGZJ8m6XZJxMWiKyffKLRBwhUTDcU
XlCjCKIN+gyX6fbLEETaBJv52To3pEBZFKNV4kjsPU1tufVOJW68vspZRRPpni7w
Jpn9Pel2O/VrklhjGsIc2BJbag0PAh30A+cSDnz6/NpHB+J2w0ImPMmyiOma77tn
uPxQI3JfoIqr0crjvMwpQUoVtrJOuc+OzdUzwg5gyBD8axi6Spa+mLne8qyx2Jnb
6jQE8CjhbN9f+wtEFGdS4RLd9JQ4Z0qj6MeCK5ymga0LSnKTb6njDzR4UB1QHiKW
865MDTXBdot9aXhq/W6WkZOqQ+3I7CnC/Zii77jNKKT78SsKFtKgd7yFOYLCxc0A
q9Bw1RBc6y0MbzHjU4kROjuEvEj+FBB3LP1mnh+9gyiIo6JAMZ0v5wQgup9HDUzg
ofdVE+vjUgkAC80/WQdCN55LdQAUvjntforZZxubOD1D8pWtbaBP7mWF8NuAIB/2
nVY3rQDhCpBxlCJDQ5LkQObCEkg2G575B0QWwShiQzkM1RjmLAlei6Albfkj1j6J
PfnkbRLx5GVHt8BPqQvrTXKsrBF9pJfb0sp7671SJ2IeVEIr3dPAuvhgqaDe7a3W
bWU4GXgT8e/4JLQUGxI0FnPV9KrZq9m5JcE0YKEIWWDi6cl66HMSRJKq5WG1lK4k
4aHM7XpmD8WsktculKk3pcO5uaked6lZcYTJ3jqARKeCwIFo7tiiIR8i+dvIwU76
oduVCe1jdIls3LcSMESEplB5V14aFFmPHhbKerHLmz5OjKnIigY0lP3glbwvrkFn
7fsshzEw3lieAEo6UTkMNKovsjGDwN7HL7gd2Pd92WirHVOWss+CF5iuqZmL9L7G
hsXKMsusUWFgTWQVLxftZObGOZ68fpDIm8TfhHuh6Eg1tP2vKGtxuNw598BfrVdA
uzcT3ginwPDMOV1BsMilguVK+HWPCnI5hDeV2lwlQQJyY4U5KIb2unPi6P75e80g
370tyh6gW8IniSNH6GEiJ8T265Ew1vTuyj8GmawZQq3Skn0pj9Iy0TDvLtH3tIsR
UHkeI+Tu22iEZQNUCi57WE23QraX2SAOwUZB4ufVL5DpD2euHdiYZqsSb5ItoeNr
/n9K2kUaz4VwQ0Qq/dU6PLtgoe/upSyfg7Ty4OIAb+pn7JMTL2zmlTM3vIhOqjib
d1jOJmbFu32H+W8y5J5G9pTIEDyZiLwRu6EKfGrspZV7jr0K1mJWiZ/2xEZETzub
mCvC/4PFNDmcJzkIna9hk+GcnyjondeWWB2nME0Du17QmFxDlJf1fSDxFBMYeSbc
rOOm0ea4BiKxy0wlyYJSTgHutJwEWGZw4kJzRlHXaL7+9EeoraOOTrQQ5ezRXWL6
0GChcE5d90mE8zELagZDdlBcT2ERH6XogKZ+Uh9TkvQA0+eK9TS+F86BykGYCGBD
hg2tA8nRk0jFK+XS5qlX4sp5hErgBBFGfheaEzeigmwuTw5Fh9PylxisnQoCY/AO
NM27UqOWw8+2uWbjsBVrlkhqXGydm3Y0cSiFeo0W63DkzoOZg9SZ98s3zh3VXxzP
iIAeE1EHzatCSYxWdlhpv6wa9trD1giPcvBOM+H+k3cIcLkOiNIVKnY1wuWYJXbl
5WJZ3zAlCBI70UXjBaPrVvfyHB5ANHDf1XM3Nl2YzeJbVI9UpHw4esBCaVknFbip
6MBHf2pR0JuPD2iuubFiLYRB8G5cZ0qlxmy2RPIhUXGBzsqoQcAQmap3JV0u0PG/
Tgrd+q1idYxP3VbarVzlMzDQC1I9lS6ZB38phHVlf5fihho05Ls9qi3ZA6jpke9L
roUHr/enXhEfGABV6b9x8t741NJG0ONLN0gk0pW1HY5L3bKbIdKUXm0VDtkru26p
28UBSFSyZDpajlXpENo8VPUtALHYuqCEkXWRC7buQlec1ejRkvz8PPXTYBNXc301
oK8ZSjzOhbKLJwL3/eZYd5ur6xOCRCreQozfxB4oix0blzn9IcSdYpc5AoaaBEW8
ftiNEG8ZYwUK8iCvB4vVTraHJ/6DKDCEtZxe9Qld27zcO/v5/7aVPQJoH/Q9IOjM
nuVSRdwdFnWofX6s5ITwYCVY64F4W7Aa81+cvnIxKXWyu7FAAYRl1GdhN6j8AmvU
AM4apW5HswvmTGE1WZ3zsjGRr3gEfjfofxzPFqaGUAzHox1DC4IFjIrzki0QfNID
Njrs7vrDiBGt+hfVpWgQ6s6TV9ejJq1NMm89XvI1mBa8w2z43fmkzDj/OBOEdb8U
X/YlmUhUsS/qZINbuh2XPo5tnHlDjpOu5j+nn9mghmrnRtFP2LASN6z0WNtg/o6V
inwrDUMLdZDUhDj6V8bfiWpIL6l4Gxp0pc0xe5slELKnzBvlnMfTmiYcweK1i4Z3
6cbRd5tZjcEDLgYSgFaI5wM7xIgbpGqvpZ3Ft+2SiC/x83mq/n3nNEZ3MT7NIBJ3
eQGIKpj3RCDvU/1F2PxX9NmNK6j+ICHw0kqzmXvNlhDpJECM1N4yFHnWeowTLJpK
ARJvMeP2Ddn58roWnC0RtqiOWUoGqATEhXUk7CrkhMQD+inWn+vWr4sM7+CEG5Qd
4IFYKLjis9FveIlcoWXOG8osQYAzfp/U8yRJMlnupaCTqn2bxcJZ3idpny6XsyG+
1i9ZxwzaAVhuJkHigPvjthWiSfbY3ykgRur5CkkGrkNWX2htgrp67q5CmFpa4rVA
twgC6kbV8GdxhZuBPh/Psp5BxfXrWkwD5zUQ7L00+I4N1MeOuRfZfG3fJZ07U4wL
bh21/G9NvbO1LC1pswzNi6Iw2dwbL+51ABbkwdCNoTe2wCeIz++04PsmqGyVyGIE
46NddiDBhgGnyNPM899BLIkPeD2/sPRAIf/sAG6bylD9k9nHfl4wW9WNienKvt99
2WRbvaUZ8+Cg+iys4WjzgnTsNUFS5nXsvgiQ29SvQAJGzBS/uRF0HQmXZTrwyzJv
4N8k5ND+qnmzX6lQtayjUTvYOEvqiRmy5HjOWdpi7LTbW0g9I4qWtZMD1m2+JYv3
3p7sQ9Hmk0FGC1Z+V+Sl/3s6vv8pYn/aJIPgbdsbdJ07W1FuGNdN841G04d+dDVH
XkyzelAgRDzZdLqCHyovsit8lQdpBhuhtSU8BlWpoH2ysRJ3afokWBUg6aH4vilk
PajZICHPR+2VhlFo8iqB7bgm7q9JAiDNBPfxsuRR2+XicYLOx4JQ2KHPFP+/jPGU
gaxvL1cQkplsBQogSx7QXbtVh+ZKe/b+on/ntysHzch0lw4suWF40kLLhCIsGcqz
pR61MO862+pIrM8amx+cR61lqv4dp6VNhYTsUA7FEsUq0Z2/kfiPdhmnTaQeD5BV
I1GvRF7ReywYlmVzFW4KulYSlsQeXXC9E/Nhnt482HUQSti+ZTl7Z9csepePDORc
OkbCKf4bSK1Nk2N+RfGY049djXt8mt+kvwP+0uoUod2SVwc+G8SKcOKnbYrJe+oU
xrG2pSJnPQWJFRX01EnPNGZhtTnqyk6O0TAaWs9ydMegRDgmfITErSHBPgUQLGIQ
MxZgjXeQaYXQ9yLRd7ZfBwQ25BdVTyBqcd+YgRVaA18h0uiLRV1ECIv/Jl5kbrow
3jRtIqW9NbdPzN3l9JaDFqvf/sUj484V6N45Foc68z4dqB93DEENMXe7s9apRtAm
LcoWJEIKrbFMtrMCsmi/qtBvjx0oXWtNGL/DWYkjEkivtw09f81BpTT7unWWhaoE
EGTyF0Y632M9NDAMcrTaMLQK2tCs0zgyNq48XhVZhCd+FNGYKvX0mcUWzo55tQb1
i2jzH7vRLNjcA5L+eWMrYpMwXovhMQhMN2IPoLBu2Aqi7gzfRC2w7GDRIPY9eqFg
gF5HQw8achctQ5TacJ+bWJ9YRtj2gaDwoqm58DxuARGm4Us6I88+jgBvF0jPuDz+
PJVB+XR/443EnRY9wwkE9+/YllnsiGCgFYwxCRuY+bIt7KgzLcIutOLeVb3Ye9Y4
y/NlTt+XHi+p5zavUzOdKfMvlWCIrtkdEnfUkIgItrkgIFr909rVy12tj69x6uaX
3+1Qpnz/KNI4yDCPiqUS6caJsSUPu0Hfd6vecYQ1PozmE9lzI9dldClKEiQFK9lD
8WFBxzeW+R1wh3TN+EmIZTRFuObNOLuXJciDaQnkaP1/lUh2NI9jfwubMylpaexn
JxpWVVRbTBSOsuiEJ4wGsA4Jln2DpvOaqFazMgjjzQ7tzkfSwwnR9SqMmw8fje1I
RDdWPg+XdyzNQm3B9hoA8EquypAtHI49pSh5y0f+JkPEu6XFKxnaX2ZVnQBcZUXl
9IL1EXlB7pdFetjY9qyp6nbUIFIVnmp6Nf/q4hJZSFqL01czq2mlGL9RWtL9/K+J
u0DCudkcC2Xl3V8yjLRA/1yJaUepy+FLNCLA8nXwldA2PDKkbnCfWC3ladURr6Iw
4Eg2MwyY5GJqa6JvkOi5DY5QqXeVpFO4buAdMI82sQ0NWDTzlk8x4ZMtT08C8JGX
dRPr0Pq6aNM4xGHMnCGbw8YGGVUddyEtaqMTs/aX0EeuYESK2EGVEI3jgaXtYNLj
CfRpaJEsWuoN5nCF2/z37lbsxAPyMvwZqCW4yxr/gVlBjgVAf7XhNRF7DX2M+pMv
y9vIRd7jkkPI+NJAEGNkrlTLuYmGsjxyK+TuydwEvukh2pIPqFgnpAFIQElCDRSu
/7F5cvYmoiJLJQpdyKfH3hS/tFQje5QTb7LL4+LMxavOUzfCHyD6U8iwSHBJFbPn
T66+iBmcqPWOSZgw8Ex5dlNtxXjjzrzt7c94m+/aL3Ch5JM74fRvx22pXnIu4RtH
DsRb/XdBrHRQ4xesg4WR3Zw4X7CAxare+tHJQ1vkmnJJXMOkO215/WS/6mVYPdg+
VR7AD/mJIxgKSU1F0ZL+WNVcZcs9f5hpLR8DVEW7PBm7WqsQDeK6msMyVYeAQ1n+
v1fRHpRqUXdCbtz589hvYMrjE49zrJD10G3mHBs/6F/PgT/oTbLVoVC2f7OqQdfM
5Ut4biIkG0tDJ9ZKe3g/TgR+zQVo/s2vz0Zl9z93QAUkyaF3BDKGOQQuKUcnQ3eE
NlzKXmMxh/pVWrBCC0Hv4XHNRdDgYZ5n5qafr1CtuWmRGnbmdHNA68mfQRySslKS
iUnm9nqIPZBVFFeayoUjNfQHCKILKXHnnj81Xv0LILnbW1zA/cNQyYpGlzsKQ3HP
oVh4AfEACwulrE8BBXiMwRKYZ8aXXhCcxYRDgNu106ZmGmtdXG2glxkXSAFMOiQI
+gIS1ry/usEvzSO4GRs2l0J8r6T6onuKczOFbDlcBE6gN8HRWStPJEZmL6DnfbA5
8NsPaphEUdtSmi+yeARGScl7/g2/IcMmL7yRm7lzTxmIQgvc+/k2bVxjMCVMpdjN
BWtnmiRHVeQJCYZPt9zXPBZNi3IA3p73oz9HgiGygF3ixzsjEOP2KdIbpa9qWsN/
UXspOuYvixR6b34iYDWvxTTGlXHctRbZ1rdxkLkt+qklinWQU8NBQ0Nkmyl7vLTu
kuCsXhsqbm4spnVkFyvwIqNhOToIzWdH4AkTxsRfiSS0O9iNPy9rvxJEqnGqVMv3
7RxC2IJbpMdPBqGxumCNTlQfskrDRDRtINOmQ7/TTTz2Ty3rMScy+rdiaVXHSKBr
HqdtMiC9j2hFx++BW8q3WUHQ+vK2LydXZ4xnkXm9wc1/oAd1WGyl3gJ437PRCjSJ
VkSaE6gmDL198Uw3D83EaiYKmGA7tu9O5zSCxtG3Us9Z7kWJsT4uS5A/Gn1YNsAt
xfedSZ9nQiJRKiA7uad1d9bmw46UrYXN5fvcCkUbw/DrL3PlVtrCOTInzn5NvtNI
oGqYmYTU0IoRH5SmeWwOBMx/uBrA9pyTQ9rzVvCiAuBtwn8A497HBm3fyepLFhON
fEWofABK4fXoSD9cPh1JGh6zowXvY7wweDHiYwSsztr1WP1ILT8h2h+K47C6qMOl
eohT7JLM13EXFVcRUqVUoRXiAH1D7wcrM5RxI4O8FuHJX/2x31xQpFucUVKIouER
IAEUh/UpE/VTK3IgkU0oFdkhWFZlOPGh+ra/KSGcMiLwFwGOHTdSOlOtxcFEkoQ9
Nj4ABSFbT9J1vepIa5H/VHj7LC8Lj26f0WYy9zGKhPOSRTEJnKfe3H+sMJ56qMr9
1tGOgrwvAmmFI0mfWckpWkkKm64e29hn1Aso8bi4D/YsW+Ze9BqmMXCsnMW2UKWY
TRMQfepYiqYLxs3KnSI7lei5aq28IR4DA1+8/YMIYWQ0C0iPNXniTyk8+KPPtGeN
gvWzUC+ScHToZJ4BDeF4/Ls5DrPoczi5RELRtQufo+Je4knKUfcJJGi1QYuqT2aN
PeOwwNMyR54yWFLKG7skXd3swzf/NyuKMFFYzVuuUoogToUcE2AtDEZ2Tyl5ttuD
PTelhygCOMXaaB5TB+2vNAsFD9OFm+/WLq8juQif/+aOfPMlK9SQQjXpqaPLzqvn
a0TLcDNExlgG2C6Lk0IjNwocRdYjmKZ7kd9U0LFM+HT6VqxrYvTmIYVbfP0LZjJy
0BNaikwrawzwiWeswhpIAmBd0cHD7UXcd1LOHdRsrAj1U9gCA40X81aEOuS0Dbhm
B3mQYolasDg8ZTND66VhgoaT45d3igwCu4VXIJG5yUoaOlMvQfX0EnbtL/OTdoEp
xLuwFRFZYlAIl1QR6Ey4scbGTsX95hGw0OKu5eUZ3GNfiP3ISQnbJb6eMuXIZY07
+F7xRaNfDRVdLKhG+fT9FossTsMa5XIgnTMCFvnO+8t9JLFGw1j51eKoSHI+h5XH
kUV4APXnJ9zYQYLIzPqvhfGXlwUJeCzDZ/+AdmuzTIqWSl30zG7vlNS846b9TxDb
6G0u9kkJ47nhQarsQIvY4a3LxcS7wxzj76jRd7mK6ubxgiZrsfyEr+DA9GyLbFub
ZUz/Gh91cw+ZmBb6wp/DPsonXrqSLO+eK2F12UjVE/xEqWiAI6t95ehC0C0MMZhQ
9rW4Y97KZyDN3uklEs/z/bHADkNjfDxeSVG0s8QUAPOuynhsLh6l0i7MGsWaZIBJ
lM5wrN1yxmedB8RERz0M5GsR4pLBKab+yU9A3P+kgcPYaD/PQlGnXnBaTjARMJYq
owI5iTtW+tWfqLZEbdChRCmf1DxevCXv1Wyr2xUOCRQJadzpb0M1xHV1gmrjjWab
zWpAxZFKDC2MZ0jvcBg8LDL9m7ohnv9JWNRgLvGQX+9HL1HZGhyd0PfZ3jDdC31R
AIQ4dl0pqQqeMc4KcHuRqn2bVumsZ5fEl+7OklEi+Bm7h0G6JxClSEjBI5gHu7kb
1D8AvkyNHdiHBSg0IsPe0MyaWuVSg1qQPVx3LB5UjpPiIJ7fd/WaCPPsFLKmVz+2
8H9r8UJ2OHKiAh2nYNWc2f6q2026THsSu0Lh9avIPVIltwJNauEQlA8b3B8rdOTD
+grLEre1XP+NKo5zexejXEr9RMYdyHgQJXHOIrFZAczlRkRRpk83I+utdPNxQDGQ
Q3EU7PWN2GUOqzSDCgAIqolrasaTcN8hZS2JRjVah9di76mGTi8vsA/65FfO0GHe
NjebdIsMo3UdftU8F8QCILAK7lVWtJ5bm321s13/DDxw+9vN9xayhvwL/XcXSmfm
jUAI3l++q6zTNx5x3l4/1STeciiq44dQz29QWVkMSG/9jyb6ui2bm5qpXLzRBvmp
Kp/CzzmeMVytIPNiRiKAy37yPgfWylC02RpdRk/5i0tAj7CFabnB6Q+Jpg33YFDL
lkFrSXuATOPehVWNR89F+sHsGcsbDCfyO0Y7pmMgiANTVIpiFelu+xLJF02zq9qL
NnkYib9tOwrzcsrjtezjXh6X0UhtUDKC9v2ko7FkFP9GFCI6viOb8JnSTDtkRs0x
yTThzR88u1eD1dr/u19NOmYiYiEaKqLzkOOsHDcp5Vhc36ocsI1NIDBCbmufyuMa
V5fh1T/+1OpRCvtcVp1VEuFrFooMcgu+k317ymsHXj/6+Qcbh8pqB4HAP44kuKRC
nFqHZ9srFoFA0dRm8HKuIidBSMTp6AUJ/HCd+0h/ah44JCKUHW2LFniQQ7JvCtoQ
ieYs7sOoy3r62gH+Ns4sbjiU5Cgppzs7ncejRJw51ptF9MXLsz3EWAyls0DkuZui
z4Gcdve6sQUmc+WG2/jMkmYoOhM/OgVnI5SFvcBbgGtvfUJgzalNGFxHjHxEoE8D
BwTM9sh4vdn9xd7jN7iNyajwq31g6fCsYT4wIcXRtty1T3q9exiQa+d2zDTQk5Xw
LYvo4ncfsAplqgLiJoVddjJoB/KRd1Y+EEfvJejGN44VFM4VOuA5uI7h5iGAbgOf
i8LWn2YtIfY2ldGO1vmSG4GvSjZpIv6IyhJsXBKG+p889HtMk92xvrmw9neizkV/
FVKHQ27G6t085dP5cFh/OwlbMnMVkV5H3VAY+GjCH6XIl0QNoc3IHeOIq9e8EAIi
jmBvQtZAfoqRyJapDCumCnDrubOO9NZEjWMg45W/HR6iYUFzMtAcklf/EnCtNR7X
Cc5DinjK+sWXjawjDltTMDMI4LsVvqtEp4xBXjRI4UeGqTvPrxSfHvFCbTrg0BMX
kzdtJ8eHeiMVOhSneePzERY8kMaz7tYcypyohBtcaY9ZvGu7HI4tPOLTScMunxcO
UfDWymglvqi80/IZ4xFLRZ0jeS6Ln3pCp/iQlM+arm9YOazEPpkRcxh0QjMOcB2Y
Kg6uoF6IaBsOZ+XUhNve3cRWG/5I6JyRAYRXaafYeuz5WRMYuFkZbtxOBvTgNxp+
ftCree1UyNrBXGmVjT1YcxYz5/XMRDkWQmBOnkR+8EXgywaLHvCV1l7YWFxFHTk9
Up084RTPRFzWqpwJ4Wedl/wYATVTsBliaD3liURrmw2aLxFtknTk6/cciZa7pNzM
XDxxnzsICNF1EafRH4SxTMWwjAv9J6ZmyDTc7yUR/T8iVL/VBTn1gnv2ems8UuIO
S54tWZ7ZBLHHrXm2teRV+elX+6JO40i0pXZoWgve0Fe8nG+L7gf272n7AVmim15e
Wq7AODVVm7DUi5bZXHZBFPpW1ViXg4ey2Uyi+dWha21Y4nY1+SmWA9guYYBkf9Xx
+nvx6uQEz8Dp6mhV+IPd5CD7J/UdhS6Lx2hQ8cGC4TOI2UKlDkaBAvs1Vfb2o/8K
iN+xoAM4zv5PZyQTuAIQn3EyFqNa8xjYCPaR/9hlR17cS96+NeGNB5GpG1kI74qN
yoHWYxJkrUx4vrvC+n6wSCIwBZvZk11nh2zll7IMfrreBqAyEOgxyaU4Pyc3xaWq
X27ITIVEzf+jb473msgEn6igsn3eIVXGngacRpvLTm30JOn2BxQVIiQygkq12IE2
GAVyDGhTMmBqIGpIAl4xDeqP/KdyWJI3qIOw5uLKJIJalj6jBbN2MapHpIIKLvJZ
VENrxBkDYQB5vLQCH5Fdq/FzfUEx+aDzKTA0VSkakiFeC1Mc/JklkiO3QLDqrBXw
K4k8dsuMHMfEtcU68EyGEs8YR1bL5h/9DgEnUSWtSKhS3OtN1OPKBE/j0S52f5QT
gG9ysREiPAEFYwUuvN6U1t2lahfxj5DL3E9+gqFznqV3oxEn1/AXK1yXdgjXMY/q
RxPtLm90UN0LFAvA82IbaWAjwJHYczoO8gmqzpqJ2qMf2rEud3vXdZw5DIpKvsBe
GqSgUDbiG1J+E2dqP3oD8Levx4RXPDlf1WrBv7waSQDatys1tvhmMc8T2wG0AXuT
NSYqVWFnfAH8gPIk2a1bTXe1HgmXdov0bHZUpmBnirpmR3qBBksUcgtb2omb4XA7
U230vCAAzjhJMBqlyYSGqHUcsLKIKsyvAScyel89D2BnZnufmkfS8LQ2R0aZhSsB
qfB+0v6hBOT5rsbifvzsj02W+6lNgVPPuhNIpjZSvSYYs0F+KuT6IZKitvpC1wxA
TCQn7gVic0QDH9/DhbzndC+GkBBJyhRNu2emSx3UVYpw3g8YPKHYnWqNaRjEhHNz
NnjM+N8MEkJk/DoJyRnidfYgzkZwSqGPNzDhDWBkimse1vy2TCna8f85AF0n7rbI
4qXPzg45Q2eX4NvkHLRU6GQREuK1PaG8KMiDH7n7x2Z/xbLESntWoe2GAQwCkFXv
ZTcNo7G01TzR7jiF2Z8S2gV4kpGs93CtQL9zT68cSLiiTATqKpqdxUC/AAVaW3KN
n6bRUHTmNBla1OAPPFjn21AHaWdTTMb3w/COYO6mW7kF5ioIiW3nCN5pVCCIeoDD
xAOkqqhObGI8ZqUaKD602P7S2zBjYDPwH8gQxbmge5lsgVMOkLyVvBOldGKLCMA/
NyAlVSNgxWIkE0faK6MwmtXrccuxM1Mzws/yWBUiwOu0raKLUfGzcfb+OQlbU6ae
oyNaSSmz5gwU/VpWNKseRkGLt3AI37GJ5aDzAkyHa78reXmyEAswfu16dakNvepY
ALp9Eufwed7897x0CADwlKTuO4c29fLf8e1KGj4AZsFlJ0gEhb1aCDkCkAkZfucR
AZuvnnnQhb7eHnRDWrIlGFWArupjANwmEPvW7sekVQYeyoQaBeqv4sRoFpjyGz+B
eGxXiCbJqCo10Ez8FP9x/dreHELcGejKfifSjE9Eszq0E9oyY0cIx6qaO7NAD3G0
eyXcWB6ycUYoL+TdiodL2GQvUIpaLS7m7XRK2bap1FWIEwBnzbfWMDqrvmKDOBxB
OiWtL5FmSir2tYN657wd0TZ/e+EJQ95jzat217LpqO2Nhz2MbRqTI/Yl5s8dZuzU
fEJqAWYd8l1d6GB79gwzY+kgJDeyaIExncVSyuwvkAM0WVb3bOs3FP6fLvw4bMMO
6+B2IhN/pVaAed4xJOpEdBoTo+LZUNXdH6fxyntAWEQ8MDuR4ebm1haBdWIP4uP2
5W/tK07y1iPgYrlnfYaroqT+9BRolU7fbs15hWKv17aSXMby0EX1NodrAsq//fS+
z3EILmCy2Q6P/livqX5bSavfuhQ+LzZTv3WG/wGLFQq4zX+zBGZaLdvwAZutjb7d
hdjMlINCJ4NcUgeRPmUCpDVSxhfg6EbsUEUYQuQErTp/wcvbap/05de/RWSSMU7/
o3IQ7EsBPPQSSWSThkPztgjqpnDSU7/ljiiszIWgr6MBj4l5Uzu0EelkZt7MNiVM
fqUZovlftJTx4o7GMH3J4nrjAS9/QyMDdi51BPFgl3XsVF/7uwZsXl330VkRWbaN
QR30pNraCbn93yHSass8IR8u0rogNi8Lyf/FkzQpEc0TJ8c8zwBppPMGXWCCkgDy
ONlmECWomFWFZWdyFJz+MklpqRUNTmjXnWOhcGjOXtqaFJqAwyYHlhgX8q29b+aB
n9ZVFefdEcctzCd8M9lZyEmevarH04xRiikLnd53ZYEIpHbB9O9zrZ57InwRL1/Y
93dcb8pI/jY5RkzIyb1u6Bc+wAlDib13de3rk6JjVsU+3dzm5ugznx+V9J+Ezp+Y
wh3FWMbFRm0mZrlSLoYm2CYc/kNhBcOfLUWXp4YOC9EEWOBwhGYX4Ao+eJ/7ISLX
ZztjE6fJb79tWBNH4W175hNTZ0Kg4jADj2GUxdNB5BvF9uMWSoeWzKMiN6NjmHi8
GE29I9Enshxa9EqvvQrv3z8JM28qSa20EL5+QY/m6vLj0iM8L8U2B8PbVzCk4nEp
qaP/EKcB4sNns5WdwjfmxRngaCGbJkX/liZxwdlWnjQZ4iatV5iew/g6Tw+KG+H5
+LTqELsbLEmOg9o5m98KmD3Laakuo/0PUKx9D6nC7x/a8ScvBPXNuUak+elngcsb
YvxmjV6ZfuZJdNpYWHdEESdW1WPpLWP5bve+RrxhBkALBiUmDCkPfRkiqH61e2mA
KF2FnizHhudhdTQeAN2Y+QNP5aBh2/J5cs5rikvDqWleafevj2EAIcfmI3+JHq8a
oDTpNO1dXBrPzand9TVj1unU2zALH97i3g8KHbupFpYy6QrfykDFuWKQn08l31yt
Gi9uYwqiAzrJRikrJWSYY6Qj67Pviyn82J3wq8t2yhyG60VpjmiwS9wMBlpruyv1
iIACpq1/M9u3fpozOaF3tQjYtTG096tpHwSxqEd0cSnBsita0OQgeiamz3HrlD9E
3QOkVmtj800YA0se2BKwSGwdZH5hPVooFYX+kdhS0DZ2Mypnktd2zYFAWn3vkAfI
27I/6pXXQ1P+CmKqhzbAHJ4l8buAtH+ufordgLWJwApsfpbfoqB9fVBLLEDBHTCP
Ti21p9OROrMpR1bOlE9lsuA9vZZekl9gCf7hdJH89LjHj7nSimfOtTVN65jmAp3G
ZbTjPkfLyLuz+X2QOfUASNM88kIVkVtxjW7kBSdMFTYMun2+z3MMU3LoAM+Ork6v
6iJfv08WP1OeaMjoBx64o8eKYH5ebX/pv0OP6JQDxmJgib0W+RmbYT+nl1Xh3yo1
N7RikMlbfJx/TiaCMq0k89SGTp92uBvfRWNO4hgcUi7RZIEnjSf7QZkKmRLzVQbD
tbVqJ83L3dnrndmKaW3XqA7iQXubVPFT+4a/B+NCd2ZAhqffJ5P324woFtaj46K+
xFw55+isW/M9uXvt26E2bu5E2MmKLaAjWcZ7JefP3gl5MOjmcjNfx0rkneJN00AO
v3P95OKuKiF3liDKXJ0AbxorYPzdlge2Jeg0YyGqO5+aYZepATeq92vxAWajTEst
znTO0u1xUwH19Bf/PNTyYc7vsFRsmxsVwwo9fsYSragLRICyh9U/R0exf/7mIyx+
E+qnuj701wKfjQ4pUuck5ETRUeKzI1/tFkTTOlktNSWUJo2VSP9CoJyzA3ONshRT
sX0o8Z9VV9uNNNICin6vu2lNC6r4Sdr3HvrURLI/IcJbgBhGAE0Szwf4xE9L0Oj7
twEMMsgmM0+8qGDiKD5fQD8eG30z4XDrYJmBlx2MorICtDmQjjwOUTC0iFD5edF5
20DcLPCsrRm/5yaU626D1fXWlyXuEMrSsr6sV5y6GbtkbihA1WyILGFJxwc8+yhO
I964CFN7LNtz3+ngjZIg7gwWBEzoOUcJcqHSLOY8BWaZHjtpaW9counxf1gwkhkw
Wm/CkRsvXbSwPw+7orcG5wHEedxHRE3oSiNynA8UYj2A4kni0lGhUa1tlyCiGBsq
E/Z//OmQgRRdcFTcW/uZpoaHTZgBygz+fs0RlR9CxX+2abzdLNDjjpIJmsuWA19W
+zlPD0EeY2YD4pYZZOjwdzIYJB9lQxBRuJI8DSldkwoauZ2jDZQQVfMsx3crADFN
5kmeOfP5E7MZ8N8yh94+S5iCeEXVohIm6c1hgbDrkRRSYysZ+ocmIiXuUplrWX13
S/aHJpfkV1TSfD/eNebXiFj5kRXxltf59DJ5Cd7lxTHWEcyjVObInnZXOd8OvlhT
D1Q5LJrdeUbItyEO0/l+ZBT6f8mr9oCYz3To0k9eKw9rRc6toqg8xNde3imISfwK
aNZ6GWlNTe3ywOUWo8K4o0Lgf2kIF5BhuJvuxdKuIGkfzQB3Eb+xwNsk6CTJ6arB
FDMhNnaO4ttu/t58nUjovhzJjuSp1jeyvxwzGkYKCEisqR5MPlWIrsgNQ4A3tpzC
fIY3Pop5uVRxxeBgugNnlaJbS/PlwMhEvRapvwfEqPt7bjiTenDFjmFQQ1O7tjza
tJmju5SosgmLJfaYJTlxLuM6sF9Oqv0tGCEhlm3vVMTJra5tM+WesZEyDCq+CJc5
TkMK9MFV1/PU4wEU+GwoGWpEoKMRXHYH4mIhE05Z+9TfJEfwEUBvKJEW3oViGYEa
W6Kp+99NO6CAhEbM19gpVIz66mNMXhpjSy6bOfE5RR/Bbc90YeXubuS7e8WGQq6A
BTk1Hyit7EAKj9Qx7aegB2iqEs7HI7OTBft2COImHEGGAanmZ/Y5YlBSjZAxCOoV
gjTZfqmNiFeXNDurgY4+COA8lY4IC3woVR/WyJeCYqc3DJtcXdAljjirb6I18qJd
QIn7VlBhawa/v6US/4nL5NK5wHcDyDu0dt4W5X9n4G7l9jxk582ObWVvZ+V6f8+t
wfDEwYciq08eJC7SD7nQfHhc61ZjXpHbBGbAw4+48uyQG1rz4XAasJVg165ot395
D7EYlGDYXOgnNI/uMj1FtaSXP/WwT8yjigOLJBJvCP56lR5Jb8pKT7bI4/Jqd1BP
qv4WA7dhTCkmBYlwvtt3HPLuzNjzHHjXnvevoHFZebx0JC3fAKKzMg2ZWnWwfNt/
75Xo3qVCzd0ONXvKyATdIYHgItRKZAT7OuMewLYhm56a+7E2vYfnTA5F3ZMpXqyS
M/fQrdMkIibtF0apPOPxiNhIQYsg7pr18Ig0dpGiHoxveMTcaPHD/wYYWESClmy1
LbwMbj0MRhJsISA8iGIq+WBG2jKxcnVY76v3tN706ozzWHhdWHgf0eW10P9Y/np+
cyWemf1GnjCzzsGdhX91kPg6VMQpSdS/eeaCuQYPsJpV7VdHR/PXDtdyMnTtcjwk
p9rosiA/D4b7cExRsAYQ18c09djgYP9LHm+qPgo5W/kfbRkRsCjwcLoPBnb7IkvF
KC+L7+pzq7OJ6HTRD8chVNOoiCEY1ya20Et2JR6z9KFtIDgHTpKIINbT7mPMRTQy
tZboKfxIyuzZON8rAFs7k/F2kCwc9Iqu7/Oquq6Ecpz4UDjOLIp9wm8NMVdw3nCC
6myxhv4HH0kmTugXi2uzsXmTjRT0UbmYbDS7DgptwRGJV6pBweuHeXJ3zQj+OVIA
tcD8h2IzTqYSkKiyHF2rQRT0WBjIKSCxq3PiUpHkDTkYzdO/CTX9SbDAC774i988
gXrz90C7h01ZC3FIYr5/V79DYm3v5wUlVV80ItdVI0c06uZncWHxRlkO/3rf/2VU
StjM4fr4rdrGQlNApMDQEmUkB+90Ken0c/mXV7InxSmEUnNUL5uzlBVE8OxjDtlg
iKYJk/aLa3Hdtz+GU2/xi+9rn6tYhn+cokI4dBP8qnZt4ZIRJPqzQuZGBQpa+N5P
4avQ4N/qJqk1pCCKewQNFRY8gSI/jGGvZCXDeq+1oCJeKP/XkIgRkvSpfcq+d+PC
kBX7nD/0XnGBCtUvkJLQ/gdg52N1XqBi7vynkdhR6svYJHcTWSa/Z05o/xc/Fh97
0GXXSFJgDl5vuDDN8z5oIvc4z0V+e0RWy0ocjcPH0Gmu9yQn5uUXtvBTri5uWFF4
QpV/hzGTxQ6a1MU9EM83WXIaKvFN+9bri3Y6ZCN4JxlBZ1MNwomlg8Ip0nMQiAjN
EC8U8Xs7nOvzKdHJsKzlHlhNjlx6TkZagYClwVZ88AsS+BBCsBAEswQultJW/Kab
Gos4DkGj8rY+Mwnq/gsbgK9JOE3ZDG8YCuPFSyIKebtazkJxBcJSRRkHu7t71ntg
NuvRkowK5WNymP2Qn9+Z3XWmCB7FKAN2Qs2Ao8gGMNO7PIsz5PavEOBTv5iH6ko8
wO41QPCz44rhDcdzVe776lhAoCQxvPLpUdXLwtBUpwTHjrs0sgpqlGtY1ANLicqj
cOtmFiBc3+9bnFkYuPMTfSY0gm3ATA6Ah3UwEJEf++Vy/MQBOyGA3b1FRgVWew/J
1S6gH1QYnFxXbgU0aKSEnTOtRAIqZ3eztIxRAD9V1GjSK4Ptg2lEgJCrqSRVfVKZ
1cTG8OKobE1JY5PshOWnyMpGTg2vHVFNuXzCWSQauBUvusYCUubMypUuwuIPiVgk
j7QuKOauGvJdL+nB7K19p8kKtCHmZikIs/c5wnK3l0ibQEKpgE0HTuYzUbSBvd41
c/FFxFp9t9L3XggeaprhD3tSO3gAvMmfFQ8kZ1vmi3N7oy+dBrdVn8qChrPMceRp
9FMGkBJuXvg05VDQ9Sklq6TCrHFyiaD4WgjspWZWWbPCUoHCUyhV53Xg1nKp5gYA
LnHOyqashdDk44fF+dqI4OGdQi007flWIAGLeC/lqKcX6BRUbotHzTm/cbkR+pox
DCrgjFxdC6VOMzK5kJaedxVdkHMsyFOqPuXUf1TIOL9Hsn1pfOVy1luM+PZirJgE
ozqz3Zy/HQRol1AFAGgq4cZEyQI5RHA85pKOh3Jpk2QSeUl6tDnr0YNcT5Bkdfbr
mi0TujqalV3VrRELKhytttCc858BAjBxz1nT77b9txWq5be2s1gfDqWuiEsO5CdL
5WzOEj/ffudLAo4V/nUgV08+nn7ND3ejUDlv2uSKTTqKk81tn+ZeclMH6Eg0imPI
HqNeZCpz/Xw1foI6AhZgrhOIWIdhbrdFy4DEBGrQus5RdyThYxEB/mq4WujFxSaw
t7JYzcO/4dN5UcHDQEeyeslIPgGCMu8bOl43uvFuOAkKI9EO9vTLPGL48RyhLKQ9
CrjGPpyEWinohoQfl7rv0QxuvG446bpD81oOEld85wJnhY5ImRb6nLUCL/u74Wyk
xIs4TVubN9OKZmBFARqg1+MwxAUVWwoLiU4F3LJykLq8DCbHWjuCqVaQUUZ/PCVN
Ib+IvGHUavfezS3PP1/p71VnOjy3D/wu8Fb5WhdpgQWWnIkvv6fIh34j543uKEIR
GBcJTFVT7uSehzpm1cLT/S/BPL7J991PkvRsFvgW3C4d1YaeojfBH02WeMx+uG89
KV5CNy9R/Root6UPucFxcKjpXDucEe8bSK8CTvJEa3lcl76QfrNq6k+3J0JmVcMc
YZK6XQ6UDCW6RYg6EXz35MfKaqSp88OKwEdIMiXQn1DITDD/QNVhvxN2A4XoyEmn
+toJnhLFoqPsBHWIlYkarFHrUGC0Y3mDQtsZTvz1AcRJtuUD7YP6kYSyOMsasqc3
HEPFY2tNITb69e5MrATWTdW/uEWo5xXxuqvyE5h0TpC/TCwxs/QCTPZ6WH8r71Ry
MlK+B25wyk8mzZ8Qc71jAQDqw+H5+VRhANcUH4YynUgkR8x1pd5lR8IgO/ZVF4PW
kz0xyqgMPl40WtGSntddAkpFlWEkfLyIlz8pkovG3mGK6cxZLchKUjTYRjZCeh9N
j2Jw/19FfV24Sbnve7kKrlHafrDHptf4BHbOF4rKudWvHUrJQWs5O/qdq9ojk2VX
9qsLW+JfJcRjVNXFVEng9IWr+jf58t1lBsVAIDn+FraGBw4O0SBB8Tn4C/xHUm5B
QUNILDbCetZmckJq6fPKR/c4d7QR/wgwEaP4uLsbsOE88dzuYJPpXGTk09YQRhBM
H7vxpk85QIzCN+HuqA/25HhooO/wqeyM8CLP9IvHVNZfLWDxp+yiS0Q5qBLnk0N9
kmaWrftLOiVMVu97TEkesTxcOSB6CiwA1eZaGV2Shyj/YZuSd457Oicmm0z3lET+
U0FoAp9CeJz5QwsggdAGDYynojTjWPF55KyIHT3TzPrNlyZfLaevBKVGhbrXCknQ
u6mZwrzRNFkKyqbXoyvZKPEq5lMLEcARaB/KtwIo4dAde+tzNPZZEBIt7EU/4whm
LprJAVcG6jsFPiEQmD0S9kg6owUPd2On1k9GtQpu1H3Mvqnpey4X52UzFn9ZkdF1
Lv//aS4Vn4LPiY44PkCIm8+yjlc4qc/6w5BoZqFqi5RKNq69mwWaoy1MaODK3pN8
3UW1SA/ArZCmnz0X/rZigwqIcT3LD9IFLnvRo6P85o2M53sgT8PTabe4QC0X1Mmm
9Ooj4h/RCsykxpqMnLfJ97BBP4O/VifJMfzidKQUCbBvncCNmYBzgJcvMFuCAhHF
p14G2qBGAwUNvrwAUqr1jUyK+UXfFSydp9EaWLP3Nd9W9Ume3Kc1mQ5C5uSbPCjt
8Uqiw9E5pdjv63zKyez3WTxP8mpGOpYyAuPhBtuU6LhjZusTxm4ZOCt3B1DSHM0A
t9M1KA2fAn0DlVpDWiRod94W0OHBkIxSt72hMzKGa8+gPK9tTX8npyamwCJLSNC6
YtoXH4U5kM2vNV4HelWdXQR3W3NE6hYpokjO/o/v35Pzchh2iED3MMLbZT3nM3E8
RuxGwSCXQG2UC/J0Z9S93NDndVbvbLk9a/sr5rwZN5NqgTGhS7T6B8OglwjiSEwr
VzMPoQDvP9Jh19wR/LaxcaGS8Q3Vlz+QCgCQ15QsQqXy3GKBGddjF+FpEKVIj5Ow
wX3Am7Jxbk6HQ38Q8HseHRZRhP8GQkmxpIzZYSwwDLFXYA7c32Bx091GAIKJb0GG
6UxpanokwXDkogNX7Kl27H7TO005IufbFHqAIxjSkk3TLPinjhRcx/su0M1muQHM
ZAEkJbLyJ8/PxF2oyfWkhX8v1VEG8+LyGIzo4wJoV8SRYqWoKMl/GYDkfDt0hQgq
QfQk/cscpT4U8mPVST/RVeOjsvf9i0/QmKCxRpMl+oDTK5OSgGgKD1Pc+SxDN6z2
X21C9Qdfw0P5OjqkHYLhGSt7V30fNULsapMgdjJyY7OMO94ianxYV43x145ntLHe
lP6BxoW6PudnO2HhprezM0KEPWKEYt4Yd+rB/mKDXTvciJUOEQhw8bWRdOHKkSlF
CLpCr10kyczbehNgani8fVYWEsxHOKW/YGmTMa/6bzzMCab6/cM6nYDyHuX4+ZaP
zZGlYTuxeYaQi0D/H57LyHvy1VBGDAX1cXV4nu0E/yQvIFb/GnvoRu5Ugnc/gJhu
J93Glu4PFM75pnreNRviTtxEivi1XbsDcwBND52qyn6r+gVLsM9hhx+xY5YhQwkn
Vku53GV1/SQZh4mNKdy8pb/suIXa3I6eBg8cnKSgkAblVxeCP/8w0oViNyGw8v7C
F8LPectMOX0Kx+tcZpBcvX4gusZAMbQu8sFxNHvX7+Bwz78iOZ+1zcP/IwKfMVUr
VJffFHU3OtXvTopSDDv3n/MjYFO9D2xNjzFiZOSBaEzem5zmdeDUwLa/64er6uIU
rlUrSYchKGZctvqZrh1pG1pGCaaUeavQd5UjcCD0NV0upjDwAEXSEfV+otojVbbA
8Lxnf1LojJAHlpGQmAMuF9rchRCe15mCVzDflzQMNPQnHZKIwFTrgTinpStT5a9x
36mrREWShI1LRjem5hW/yfucYMDWWrPjsTXheDyHSvs23l9ZO8EGusSrLAvAdpWc
cFyPKeWgiS/CmKQjZ+P9lZ3tTQw2GgCQZMJEL71SPmd3hdDOEqipJDF8R40jawYB
JHM+zvos7pHaNmF/vIIjpIz3cNuTMaTyfeFCCQaFmqvAf1uqzSEJ1Y20txyWgASD
D0H1Alu6xbmJAUCelbOjcjrv8s3Env51UU51MVzXIf+kfwvRWXMnwPvGhMp6v4mv
w4aERta2aYQCOgmcce3W0fTDLQgKvwjS/w9LNRXD6Lvlu9dvkNjTRegOr3ZFroRH
Mb31YrzMYwNkSjfWCVg1YEELnA14dPRnyUR9Iqd3eUbh7xTOu+YNg3q3VZelI8rL
+yiHtvrYMDdToJ+aikJ053RtBisectk3yhSDgr2y7+ZxDdUsHk7WG7GK4dL3jX+/
Lo1Y/eD1p5Wfh6RVEzVcScvIc1UpXXgOY+swDSW4rfKr+92XZCeEIMysj/N8bIie
Cf+DcEJ2QxZ91yVeMSFaAHY03UomUuKe4/22g37BfSDpktNjpeS5BtigqIK/jruN
AzOCpRMJtNIf2+xF1uhVRaU45hAcaDFcAeIahYdoAusgJ4iDOUvin4tm9cwmXDJB
mS8fstwpyx27AuEJW+2vG2hiBczPIYIs2aW0lTGsbh9kvTrE+qsG6i4ACLeLnhI+
G67+45AzxD9LrmniM+NyAWoNfwHqLMlczhERbfuG2m2+LJJ2/yC3mkkHP6/0VBDq
tWbZBQ1WvBVLZb2VIBBwCLCd8TuGl8y0j9cT2Tkw/A4YZfteEkjhS6uXR9Y1a/xS
ayC0mT2rLNofDHs4CzxsvoUQ0GbV3B8b3+l06ZY2JJIOGpupnUKLxRY3qE3JO/cP
ze/wgSlp/2mEt6zpdpj0E4JeMxevKrve93wK9Ch5wI/HjP44saZGdJee8WgEfzO1
/Etv0FEQMVRqcYXOhIp4Zxrdv9cqLI3JgwQJ4iUoE9hNiVyVhcz4IJktAfZ8oOSw
13eb1oca4JTkyBEcOe3+EnkHyJ8LE+/lndK+PoEmKjasDjQS8lTgGBUtHVkBFw4U
QgmG0H/C8FhBI54dsegcKGM+6ov05KMWcdgwjscdPG9/ZN16kqyu17NjI2wAdBpQ
2AUaOPrI/DS927MOj/RVIYSdM5Ub1edt/xsmWsprG0fgdZI8waYv29hT8aBEFS6F
/cVL8XIxOJuowE8SlMvRBIVPbkLTiSdqhmXguAcT1yvdbCWyPGI9t4mi+kBH6hBh
IcO6aBByprZTiHP95uaiuqcJUBEVso0JvoohpG2iMQSGQ/XClLET0NHCe9nyJBgm
uVP4l6RIgT/09HjsYs/Nop1nHbhC44RCAgoFkcWbDi1QG3RRymy2z1jEkRQMqfpW
2+Eb3i2ZZ/LlgsG0hQA4CtwHP9qGO7iUlKV8cfshzPeGH7WiJi8anjqWB5+X3c9G
9R77iGI8v7fsOj25jnz1jHwV5872uUgRUBzwUAy1YgOJiBFaV0cULp26L0e+j9Tq
tWFiXlHqj0A4JV3iw7PFNU56jD88hlntuPSrGf7ALykkvSZ+fZP2xFtWqJTZBAqQ
CnXmosSn4h4jLKXsn4OiPxhXePXJQLyIOa0mfx+n7G6Y02P90tc++rD5ob3UdUob
/Jyx2Ldr3O6X66zsBSVbNt/lAv/JomQvc2CS984w41J/xM6r1Yz0KbfriwGjSORM
czxa2Gmuru298CMj2CHFysTQwVKM38c846NEudv1CyqmAF3qU4DzVp8tgeKWoc28
mly/zV+vYiKdBUMy+Z5A3+LaM28Xy/JLMBEC0tIQkRkG6+oq18UG/ub0Kh/W84AH
4HuHbKrPApjAHCCUTKLanWeAGOkQfBUzOklqLhsoJh2k1rkF5sZCrKZMJUZmeVlB
bKCKDdXzbmEEN17MGefBwTxSd6U+BOEMrxcdEI1y1umk+gBIS3oA6OAW8DJcNP38
CRRLGtnFH4By6Gktq38FMQU87mALMyLTV5qYrXoto+uXSDLZHnK4zzXEdHQwPfHf
00X9j4Ks00vKaqNBWMkcCs/+z9QQYk3tp6nUpHXq1JQvOlDXxiouoRa+b+0vX4jU
O4AbhOUxD+wf5BgHHWFGJ8dG95U2Lz0NBIIZUq8B14e5CkwEMCtsZzzdJ7HyvcZc
seur5emclXybglKELs18OHowI9j+LsWL1YstN8T5X11l+Ts6+sgnME7lzwyxHwgO
cyQjxPO1tYzp3XfXhshCWVgG+we4sU3J76uMWmFcubLCH0uIu9gddBTtpvaiDHCL
ffMsDGVZ2H72p4j+hAc/CXXl9mvQLxAfCYsr8kzgOMDdy2e4frHEK4GOX66zDUBq
G2aKLis3HrbixEwJJrpsmvTeoCbuLJAqbveGtTAED8Fs6WZnOXy5ZMMVALWme4MQ
mENcshBJqogQd8GFnMdmjEcx7C6BVYujwK/hd/urNrJbpJbZg2sONKuGC5rwKXj5
NPJy7jQEfAr5G6bWi7uFzgwm2G0pxwvmWY0OsO1n5J/G9cwnTmf/NQOn866f9ILJ
EWmFrFJ1OpwxICaLHz1pBsZnHh0odIkKXldLoolXTwqyvDTR8ZZ/AYH8dcQxixtn
cyfGz2liJPJUqdX/xjIc24foZFP/zbchcrU7VUTSSWkSwYR2ML/8bxyxPmYi0T4z
eSDukO6W76/weKZixr+0Y/QgYrDVFCavCax6DuggCEIMsZ/gifOWzdM4+Awr+fut
qCdw/r7dJK3B80QepxIpZdlqDIjVvIC4rzq0rQHC0KMEOaCotu6fqMeLdSNOBH8x
z+oJpuXrNsoPu2Z/r69zs22SPZl4jm+VAPHN0i5LDx5MryfJeYTz5A6+zL+Y+e5C
OBSRUJMs5tVBMQziSgU1R5f3fzGGkeRu1z6PFbvQ5ue3fat+eSVZvmeI2lT7fbDf
Bh2tweIi9wPN+1TnpNJCHjpnOycEW/o5B0A02V+yJSmzfRpV33G67aHFJEuokcSY
N9D8RWWWZozJJwNBGwU4jY7MYl7sBp2cw6hP7mLtjNFeRucNf6HycRX9/GDhJ6zq
7x9L2zsmph43fhJISmVee1eIwP0O/vrGT9UM424yNd+7f96yJLu07VSK1CJbP/XH
O5bPu++tpU2JGFyNmSJMDgQux1ac2gd49PRONYt+qH3bBoY9fLd26Y3PoXuUfYo1
m9q9tlG9BhdlA6kURcdVBenlR1/+FWrCRlDf61xEhs6Ai9b2tF+IzcrQUQn9XYP1
WrR+10m7hHPn6pChz1NWtnDoaIylQ9D5sTo9d4lWdT9vL9cbYaUBqUDjHouA+NY7
RpgP0f6yUc3nRMf3RbxAjw==
`pragma protect end_protected              
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
MuacxTrQ7W6gIQOlqfcrxR8ovOZIxiTSrezzKDsW9em7Mtq/K8dJSw/u2d2nTD1/
fYxysOEhK/RpBUtLF7dHpBDhsjkNsV5MSr/gESbVa87QtPqJ+XpNMX6PYfdWd6on
C35u+Oi9FFjOa36doAPxXLUYz/d3KLMLzuZC7HdPrMY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 171739    )
yDBLVsvePOz8Mjx9ssZaiRLBRDYCE4NWF//jVqG5/7LlCkY4HC/IAjwW8UFefUS4
AeK94UZ/8t/cTSPChD5eJROFg8D1D1v9jgHDekK9yqDux7za+Ugw5pxLshAu76OJ
aPpytyCCdVRGhrqJ1Sdrhe0KHP7ro28ctT/IijI62bgwo/fqtctvjztMTyaxgu4M
niX8yHz3sP3Iv3owC0Zj0gXICBzpjtr07UFlVUdgHG0f4L7TDU7hV2ysX4O+sOFL
KGEF1ogb0v3o5IFAWHpZLw==
`pragma protect end_protected              
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
XZLurifK6pQPne7QdfkrkdqBjzaHv6D0MLhOdErnQHv3RT2+5cqrXcsxypsCrJVW
AxMwF6mwFWIisqY63kcHLAEtZz3H4QeSL2dtSdBG2Fxgn0HK5C+QE4YmUZDjyg5X
n8Yoq76XQHR3KXsh/0AbzTtnZLZnFaSeSkbmSht3Dmg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 204946    )
MTIUDwTQDL/NJB5ycybOrivA8p95qM8WWOH7Oxe0PxNNvYBXuJcMMx2KDVZ+/WPP
Y066Ac2iMLFq/tFIJDqrKKGKkX6Txay0XyUQmRCVR6TNwiWE/tPEqBS7H1fCE+Ts
TVvAzyK3F1MO7XMs5euTgQO8hI1MOEFPB9gWSKGvzwpp3qyTtnzF6byahnmLFoU+
NUbGb5v4Waa/NMn5sAKrzgE2c3TCG/9125NCq8A8UTfg6iKVWYJtY1OZ2qYEaGUE
TDUEzDudKVaEZxiwqjrYTu9O6/Zsy3EGTSHMop9N/O7+fJ7QPXjxUU6jil64ZvJs
YJuAVpS3ZBaOQDzvE6s8fy0vWp/nbd+PcMd/mQZzbZBfwLaBUosi84o5UVoq3E8t
VW5VM4L2y6Wv0mCDUHbEcZU1UQSnStEPmzZYjo3idQpnXlt2GtRt0/8jQ5uB91WZ
NKL2wflX0wl4Rnb4kB9jwN5qDzq3cey19ybaRfaDWwoKDE60rSDOw7FpdprQoqqq
rvflqse/V8cNVe0PPbB7UXF3kkYT2GmF/rixb17ecHmi/ujza+dW1qSDgA3gQh4S
zW2c0/o8RcUrSBxpxsyCIe1LZMiQxA1hsRiCCs4MvOA8IrwHeukeLd/yN2VsUvpm
l1YcOiYNhSB8HxS0/iYt3LHZtKE06uoMFey+Kg2JgeEIR+UpeOGQXvWWY06APWdY
hFkWi/Z+/zZID6+haeydQ85LyrZ2Yap/Soj7fQHWlUnOVMq7X4i7uduPRPjQtHi3
n96xPZzjzBtlua8WrZRPvkv891H3T3s8+Nh2b73oJgMNiInlDTFZmGDKu1AxUS3D
/j/9ki/LdI2KyyX8Mau/uN4yI25/Ja1bZxQfdO+zsKBw9/yVaPZGP1+Taoc0zpF1
ZBcQtu4thCPFFhDnkTUhmnEf/dQGuStrUBHqFs1HW4uXOmZE//x1ca3ExfQXE9Z4
oCyd8V471D+RY8V7fSlm2lrflq9QeYSbA4/Pl/MrR0J2vi5GEquT3lwBtuKwGcAp
ohSvmrrYG54GP1/KIL9uFlC/8UrmhauEMFtui/Jij5gqZK3gzIExCdopC49fB3yT
eHgS7YSRuI20+lmT+yk3qQ7bxUJc2R2E/Czb0z5Amy/XwECyurihloD8fu4bq4PE
TC0hVoOaxyeMA/bEh/i9+3wz7mTpdJcIR/a0jfm23Khsti9p2/8sZIgE3/7EX1QZ
OTOTL6QJcP5kPsnBZBlLDEjGIyISZCTkE0oK41s2n0csa3oGULbftUTkH+rSlSkr
Np6VanvjIfe/WVloj6hJy7vCTXrDdkyGB1XWJwHnKx8Vdq/CpjgeSCBGwqzqzHRQ
Zy4u+8M7LhrAr3cmC7qySZHXmdi6g9uZzKjxRzADfuZ7GOoUUKI2Ehud7tE5zECF
JL6zjTJFJfdTnDRsDRZG+2HgAxOYMrneOhxT9kElMtFfMASbAxCXSjwKyMt0m9tV
3Kt24Wwc2OoNAMR1pdKMIVtB8yVzfZB5CyS7y4WQHMvmHqr765AqNFQtD9ohhazy
8HoTj/ljbbuTwXJMe+SFQ7350HJ9WFvgYDVUq2l6iaGUeXSyJgZJBIvNFKS0i87L
NirrTjC+EeYv6Li1Ric8cSsYr1CW+t6lwaOaabm/ZLmzulUScPYCWTCP2Pj6D0Fm
FlUFmduHUsDBs1fAVIEG4QSQrPI3aUEaKtDYftNun0ixIDi1sMavHg+E71PyWePO
t90UND1bmBX2EmMddd3XXJc8RB0x6zkzTC1Kx9ZrI2uN59bGaCtTLvWIkTjnVKKs
2ydXoY+HN0794H5CIBhYu9YG0HvNWRlSFv/tlkz1GQBopS9/+V8+99p+7jhmarmP
9KmnVSaTHakAxKNMDxDPf2BZwTLSZlreaQJ3TL3nsHmWRr1hmv01eGchlK/6bYGN
UCa0WbhU/hCNadZP+h11jt67SOOgFTNuzFebeChN34BHAkOBUjnivxWP7bWoM1P2
fKfaZy84RodWUqrSRkJ2W5mM4GW3vlnJUTaO4q6/AgOxa8wHzugzK6CCHNLuhYiM
FY1G/mNhxEYzm9LNlWr5/8xK/DZbTqe1vgHs3S+CMu5XNBkzGBHX+enRCLUbMEUa
OCHMHjj01uoh6oFzl/02cwHG0QLQdZ3WiFkfzG5LOZ1iRcLN512DJrT85bC8X1iN
Nmy2eonJmikGXFmrfRNV84gipn8+4K1PxUP3IZxVwwnMq5Vfh8y7wEuSz4nwK4fk
H/A5NnhSdQxteWl4UakcOTAu2RcV0hSEWOW83NWzXBuE7njiHtoEy8Pu+D+da9/M
IVKTln/UYcFsENQvEU4mUOryMMHHAR/QdWDVDDLWv0+cfeH74vKMF+OhHZYWsHOi
gARdUScfoiYNCuzYziFwXFShwtzvkCQiRB+6wJwbrzwSGikK3TPK//1IQBl3IN9a
7ZUAuoxViIWq5Yadgz9nj8c8fSPCp8YhxC5mT7ud477sZxoaXtzPZvAFbprIJeGV
N7hX3pQq/8m4NBE1+9HpXsBej1VNvYJyH6oY2CbAHCVlqGRtGrcBkc0wqR0bmjH/
eOBbs0AdWwzNbL3uP0mjwhZ8P6a6xX1hybFaXjXFQhb2ZxmGqWyhL3rv8JyeLnBd
3E0zusSSzUKUa5QxTv7EwfGVgKpjeD8G4kaPy4k2fkydeQcQ74JNgEV3pCcHq3FI
namnoRN/2DmYUw7WIQO8LGMnbJGQka9mdU2hmkwTKlFNQPWRoZPIzTiiiSID8SBt
4jjQEA2jntJNwq4F5PRpXDFiKC1Kxo89h7k+gUyMv+rkG7OwY0estQ2qxK5YF2Ul
yDZLzLzCbyf0BjwpJCb2OcHhowlKGjb56A8lwvOHlQJd79iypkkUb33pGFAYGyL5
NKNOjWLLuqfgI1/k/lO1ZKZOOcUj62nIa9sj5D0K9yM0f03yz/rgp1scg91LEKkK
1PpF/oE3sAO0KdsZukPiMs7waObu1G+7spaF+YYOoTYj2MZMqQWYVOmLkHunfM58
p2ja/3bcyra2dYCqA2Eb+s+Ru5gye1EePZAmXnWNih1fc6SZU9wHV6XLfD1HCCyU
wFV75KU3cvNsOWwUFbHt6UcBZVSB0v64KBAkXB4MZWVwPkzAWkBATNE7NanLkSQw
YMi3loQ+IMM7EdqHgcdg68NjO/7hUhnpRlDCP0cLXUJ/Z3ipP7TADFTKZuzldW6y
6gmlggicDZ2uj06oWQBs49ww7dnqlHyxsRQJMTZwH1G1G/XngCVGXf2Oz4vEpE+c
0lb28PVuZggVTY5RRsZOBGcjxTY/OOjlyF4LM444aYwgH+hoXyMAK/GPE+kQT3gw
ddlGSiEhQEucibS8YXPuvuKUhhToFRCdxljHoAssmGCqImTDuNlTo/NDwwtz4R54
Y5ZSMp8DpGAUmc70TszorIoth4h683Gdgss+b9HKcDElBIc2xHZz71aHJTkf2uqV
q3KOzxhqM9ZurpIqhXV3mBOsy2ghsej2ufF+KD9yKGGCZ6dixaLz/fz6HDdoAF0M
KXRCha5GCiJ0/3+mmtNvNtqy3A5eqNBOcHDVD1QvVi1A5szDCbKvUBn4V76B4Xs9
UWLC+bf9z4kjDpZ8s7gMwfV1CczsL706O2Ti12vdGMtl5YrOFPBMsNCvZ7T/Y6Iw
pax8JZq9ltAwAhqvSQ4KPiIq/DZ4eMZUNTVxOQExl4QP70wZkz+DBAdV//wgLSOC
lZnK0fyxuTzNl5ZXuTCsIPC2DV/wI73Bj2erULbfB4xS7EF6bf9KLEBtQ0k6rdI+
X68XyBSHWYjW59/cXZiooMT7c7TyPOHJOcPr994rQqfJ/a7hNsG09gJrhdKNccrr
KtiFSPpoxu2gIUQnUha1hVoq6z14xAa5EQXOq5R42kX7RnkxuRbeLOhsgvLEqJAK
iv10wTriLw+mEo5yuLFK81mp0S7yycNvshfVCB/4607qT1eTTbm/GgljKw4Go3ZT
F+ZcxJnzo/OZmhrkoy2uMMZ4MtdjVzMoOEQ2OdFU9nrqvopkNnAdPRzAboGIr+fl
n8qzQqFKuQ3AcQQAYowJ+hhgDuBSHCQ4JFXS4CpKwG/00ymMs7TUhk60eY1Z8m9I
CTxgYeoNZCDXUdLbYpMRadSeBWQ7hm5w+h9KKfw2CNZ4Vu+ECmRai014KQ14lijp
WPl+6ruc/XqURO8LTSlNwgQKsOIfrJhkpuwFrSxxUsYKHuhZIPNT9Rn12pY+KKlH
f1oJaXmvICvIQmEovpikPtXzX5IBYl0tuByecLMuRO+RgQCGW+gH2Xf7/ilOb89G
rHpu/q4NuNZN12yFuIXAwps1NAPkruigGtS5XwZjWcqPgRdWg/uCbCX+dR1LfErK
R/Yb9itYQwUHcO7U8Y8rdglDtClrIOwbTH3DZZZSNou1vtZZHrYVvQfySGSkLGHe
pzlqQZ8r6BqkCQ62LOF3cdnVFWQNsK/h/PVMyRjgud9ySSxMbT/7mquC1aYP3bhH
i1zOCcxvantJjCjoOPqJDgpZpUndEaQ7tXCs8zDiAaMgoA0N4r9jAP8cieQBcxEs
cXn1N3ipQdhsW2QJ+OL03r7FsXwtCWwTOtwlhhvGk75Kwj25idO0ZWofpQdXHCqv
c0JM2cVKAie004fWmvBWPEZkFYsCqDsO04EkpQ3mGgIuL9z/jYCpDTsKp29SD/MK
OK8w4dAiNlZfYyqPeQqQbiCgZAiLp9BXGDi9NTbXxJxy8kMzal/8/9XROCf4nVOT
tEgdeUbJroK4UaTxkd3m0uCwOlxxol8LB2H7sgxMio+jqcOc1Y/D7pPvj0n9o6SD
nhn+lCA0x5lOpduUTl66Np7P2Is9VpbJxIym1qdlhbgUyZKgwg+bjdgtiUg8eGIW
Wh/z9HHeWSsKH2kJlhQ0D7vZSzs6h0FGFOi8zzWZTile5g/lUVaRVBr7Pg9BKXNd
VKKdAXu62X2HrEYx+m1ir1WRfgu01gyQ043HRuyMJPefDFG83zxZi/tLBq+4emt4
yl3wBBoRYUSnkWo0UFrVnKtf0vCOIAMAQCL+g8Tdjaub/Z7J+AQ8SDNgl15RY59V
gUpwnfeisRbg9Ztq7IXvyuFd+RD1OXtLn0KOWzteKbT+w7eUAhs8fhke4v+Zt2G3
g7aFZwNIgCwwqE50S3F8Qq7o0IBT1qWMez8eZH/RmpuKGRtO04rl0qGAGuLxyS/7
RJSDYBi8TB1Vk4Pshu5RQ3BQT5PJNqWSCe4KUXNdvFekkWRsp3REc6wEBCi1KmLC
Mnhmv/gsmnjhABHXgu+USxjs8FomBXEW38w6d/i50DQINeg0HpGimScBGLP3BGST
gRxrPJBUBCJG7F5yA91QHb0WkReEJKfdaqzoBjsqgHIpDFojZ8MQvh6AeOZVdgbd
/6ZSV9MpWgzZnVVPmJhNUDFqJKK0iaIkpeNwdDzY7E7BIS3vRLIsegefIhl6jE9c
+druV1borpqUOv/inKGneS3b1ve1K/Nrlm7iN+MjFUgIRz+bR7lJiLJdtR0emuAX
FBaxvNFNcYCPuNuMFHh64IfYk+DAeL6zefq4nrjQYjv/Hr3zRqKOXph5AViumM1q
vBqQ/i4JTn3cSwa6WWkzzS9KgPP/qdK0QU4qgWudAt23wQQsuYGXjXZaUlm+IxUr
IfdKo8qfdI4dTRf6KvmGC+VaoDwpqhV+lnpmouTOfCA91YiLbI26ZLIn/cNr9fU0
Rdx2FpVMYTnlBcowm/c/g/sRvmWvW1CxYK7ST+o34cgW6R0KhDUkVmDUtaXODWoT
GvurwE/4VJSNFhxGxLaXs6tA4aOalkF/5fHUSlHefgtU8mONkhrs0evXf4F+MYsY
jBjB3rS/dKgJCv8P8Qp15271E0i7ryU9oQi/pETPmwSEmCL+0jB85Tg9EHMUc6IQ
VQCfKGW/L+cjCQV9TqAOH8byzEEW/X+pWE/Uc+GTYnpz+enrudnXgFxnBqViS2XX
ATAutN+NiikcxQXK8zSFlvIibmHO6oQc1x8e+xUQ4xaVour8lvptTI0gk6tqA7yT
PbldszOTDQxLZ5HCmFBO6ifDyqSBRtTkHVtIcGN8d0omTJSbTWI49yWQlwC0z6CS
USoxSL6ElCVr6DqjJt5hsgFja7VQJ5lpQxQjH63b6B8WqtCWPFqn2EInzJ5A6485
nsuTV7jw5ud4hWjSkrpc5eUjaZQKzV93dJFwTob51MLwj/FyRb6mfbnVnp9wl2Z9
78K1zOiMstyXVex8mZfoINm/HqEDQ4XW7GfONAHu3BENGqvjcDTrC5FBZrHbsjXq
heBRtv+qCY+DvOSRtduZET3mO71jhAv6hDjQXVFtOyhCYB/dTILlhPiqxPZvUoKp
BwG5l0igTOHfQrgPUTgKXct1vVGpICXfM8k/9apr53yLjBSsLvlxzZUOF7eqr3+v
mG9+XXU4NIh9SyuDL1T32OD9lP+KTiPgdDqloJb9vw0HlMk0o/ay/MGVUiTp1kcc
h2hmJTZTPPb7vO7Lvt6DpaRNNesT48As9MzjzQvUexHXvSPJD9QP+kcdsB4DOkoD
qkd3q70Dq37hi9dX/SX0xp8AGCsQ5yl1U337c/ENowErWlRaPKAKwh4t15PekxFh
zwuexzUDic3tsQe47K3F+m7jpxa3nx9IW+u520yoJtcViSmAqpZLp3ZPkOkJ3Zri
2ZHrNl1tEBjAnWQ5/ErBNahk4NrIT6CsrdkAVpic2gsDSKeM//2CSoBqHWEAC2hn
uc0F4Vw0Ix/fOGkEofhUwYgW5EO+z0/v082I48YalME5BP85RWTOEGp/hH5yEedB
myhRAalRm8WIyPi48xOLZujNLYaxPe1D4rK/CMXMSUuugSYsMcQCOnPrRHg/fHRu
v1VzgW6P7L/AWtnHTfHoMTZLGpvVlwlc5lKg68Kw7Qumsk9bAJW2fyQx0qbkAT13
MKxIk7g5c2tjl6a7OUb0Wb64cyZR2KnPOqhRlwR0RZGcoIxlZdJsTCBu8F8jzLuw
xI+fKj24iz+maujpUjyAC2cVCRcu/ZA84ifS0iB0mznxRiUNZPncAwZtFJcMdgG+
EDu0ZvrnnHpl2UtkgQbyeUK6RJP2dgimCj1X7b8t9hOG+4M90+EPtiOUWE74XdCX
xlUVkdQWLF1U4XiMJtFoa4BRICQu59VQ5dgi4flgvXnLPSf8RWI3Wqhz5YNPBc21
UX4GJC9SAvRndnyVrnvKAJqYFwXzB6NW3i56P2hLpUcf69f5ZWmz+ldtGTQti5to
+JRYSlwsGvoai0v8qDi11qHLWRmNnRVsPTFckCmi4jU0f+hmkTKn3cl0Z+l/6vDg
5TOlE6OT2fyyHzWYuE7yr0FkcraX9hyLX2rB3RZLeI58zy5I0X09fcqu+Y1h8I5M
499+EOgGA9XLZxcpKDFEcbJNzXHMQadN2fkhlE0TfaGVwL78p6iGGTuG1Xf/+/gU
s52DWXMbEo7BCzebGuOpbyisUZm701PvZN0UUO8KgHh7nPKorznBQ+X3fH16inDl
hCLDq2M6OJxODdLK85D26KSK2ykhdPmbRVxKFGCXgfrU7PmABtWKaAvFEyYQGruO
ZjYTSqHtus40u00qTGjdap8yNd0vDnh2EOh6Y5hQElo1MbFzH+N3xiH6jirjqrCN
3cUNLGxlUAYe6BItnnKUf/yWHZD+UfZ9WoOd1u3dqpy3H4npPdHEg/alCcIjZ/x1
xi3fq3mFRpEbrlB2HqJmBobc5ru9PjXivun7O+Zx/vW2qy31qEoN8aMmJcuCTLfr
OTtb/efg+OV3mH/C6kPCF500eUvQzvy+66mFkVOGgAnguM3mS75K2VtOUPYh0trk
ZjMnb+VjJbxxjVVMjRug6efCQRwVfmw+mEe3RvkiuDwXm2OzlPWMkC95i22TurPz
ZcJUhGvAXEr0uPuXVy2Gdmu2a6EmP7GS/LrA2cCU7+GZiwPxTNlKyn0QhPkJloIO
P+yzsGlzEra3NyGC7I45RuNbe9VYUNgkxas95YBsxDGHTyeu9OfoP/mvdlTVRSFL
Mg+NYugA+ib635pHykKEv6TeVORBv2BxpRuq5Wc2SoTQGZJueEhUqvKCQ1z+5bAs
y8dRL25yr9EE5Kwle84IiqXK8/9DEVdIUNJsXCJEgaV16m+WcwikZ3nIeZInc0lS
znsXzpiwKKqUgTFNRU+SaKn95z5xE+4kNqimAVbL2dbWWLR9WifrdOm5rvoN8SZu
L8sZQwlfkxshsXbSGHg3J3uXmDOazIl7HGEmWpmZq9TR877Kman06C1WkdWxwKiU
jubJpLC3nO+XpqZOMryvYNz8/+uIAHWHby2Fv1ZjkTR0ogsDrX6HWTjAiVnK+EfR
gSjdUE+DtYQenMxE2z84ufaBAvAGESRD1k0kKOTlM4bc03dtDW8VbYuNb0JzSP0T
WH3QpzTkPRr1+IL17qawMN8en4kROpbszH1YVHRn2hc9kQTcCJorxNHbP0OUiliR
t/7J/FCR/Uv4rjhaS0VwU9BC2907sM3FHPmHAbl+oT2iIH+biC9QqrlBkq+YpvDY
QdlynV3HRy9mqado/TmhghoPHBdSLluRZxrKw5MT3f8ZYZoVkP5yi4DToM12cImj
xffbubHw8N5/uQrfdI/yR4cW7SuDKkg3MAn/WddAqP23xBaCUhZAmWvhcWbGex6L
WenvFPK9hmhlBhkUjVge06XXUnO2nY4Po8kK11/zpy3dl7ewyHZ9jhl1qWI22HEc
2yxuU2UcP8Y6VcbBmu1I5TMDgo/6JiC2C4Sva+tAlxRBo7Fb5V0YwhluwsOMLDBg
MuuvC+uILYXDZ+I6EATb/0D8wPYcYwsrgtltuPuw+pr9TU93WzSET3o/Lu7D1kmn
oKn5KQaDkFw262Okg788AKJewLHDCfWKlK7bwfvQgVw81f1oWEOqzI+LhNNJpSU1
U0Jr/z4O/8sMTMC3CYzz1P80O8ktFC2IGN06Qac49BU66hiM6XnvDMXtQBknsJ1u
JXzdcAosTWkyd9Yp4aslYvTINXnaS2xhvsyDqvl7pZLia7QkqD475R/VkMVJRNbJ
JONtdjv/3dzEW4qFvOzoybyAd3Mt+33fckUy4yjjo7Cre57fQiZolKw3yCpu1fm6
e1F8jfQUsYseRKZwbaIf00NCWZtXDJtoJ1IyJetI/C1QgFVGMVRQs0V5D02/gQWV
PVfG1kKZNsdqEaupHY2iCsOZmt8JRG0kY9gnqnqnHdl/d5KWc9SeOhsbcrsl2z4M
Da2UDikOx+Afk4UL/UYGBDVwJKpuYj467IC1xeoiYEgrLvcTu8Le6Adpi3pZPvi4
QOaXDcXwWUFwOt4+UqrWOUeqCL+NYVQqyaspQrzBISKY0etHclaKJwWFwGWwInpB
oKUG3LCIWr0KY+gTNOa41EmTyQWK7fhShcrmR6b9Q+tIemG8y3ywlXwBjtES+J0B
U+aNqq0gZgzZr8zeFdbx6P9u4S4ZTh74WAo4d6F85x1EbgpHF67rwhZKIF45YnC+
C/NV157kf+VNKNCbpwWe+wS8bd7H8kzEuDlqRPA6NPWgmML8SnrsV8ufpWDXy3pw
x5ehU0Y5MoPF8wpYN3SKVctS7Bs+jGxlo2hX+0o7p5Jyw2fHQdsHp7P5pZcnk5IB
H5yukaz/OrpungTuGcRV1BhV9G68WL2HwzT7H9/EWAzglVz5G6oWIsixCztIUx//
IVQ08EScXZzHz7nRbdCx+59RYd6zauAvvANBcWQAnaF6lYERd8wt7/v04tCRtmbk
bkugl0/QFutSctsPxuch2d8qeO6AL2BzJKQxkDPHYf5gpRZIY2AGQp+tWUzr7Yg1
r/JhECDAvp4w5qGTRK/PCnEzyPhT+o84jXOfo7uzrgPJWofINGjwjfEZIZh6rJxa
mg77zeou8VVUyWmQYmiEjefHjkmTjOwlgfLub4ZQJiQt1e9kaFZMATLovVynbCnL
xLZJ6J85rIOD123nH5BN9uOLZicg1b3grT+HzzFfZ6iwWebOy8TdAUMzn8MjTlii
JGyg/EtDi+mNoA7CDb3jWj1FwPWaaZkMWqs8H2J0K38o8ezuE3op8c12Ls+epjfi
3BRLM3Phq8SVnbmuAxm0KzlW8NyJ4LzzJVBFT4dO//TZFDmifKtC+aV1OnJKfO1g
YQ/KnKQnVZg/Otp6r61ccOEbkFz3K4Prl2rVnMynNfNK9evlmivmmYrOVquBZHqV
M9jTo+oNFjOWQyWHU6yl9kqKSo+vm5FIDHOYtKN2iBstJJllCho1XWWoF4VcER4h
QKDMCLM/KSdhch4hvvNcBEFG5omICErcerGwh13qEzJTX1dbAgynUCkpK9OmdHbo
vmXKXlLwrAf4KZ0AwmCO420UdhE6EjBZbPZARHVxyvT5/oYoDR0rCUOMlDuDKcSj
fgtW9mvRHApTvsQ97rjiXEQsNe7RjUK6FFE0dc2FUOs+dZchbTe6SejjwkOW4yFS
O6+qxcy+jjH78rtRXz+izx2N8VCdSxME5VCMLOzZQ+Nfm8aSkUZkTouu0vBTvg0d
CvbsU7/0UxjPPH5+9dufL3l1Q72aA/RDk0q1s72JSJhH2J3n0oRxVyEClX3DoH+D
AlXVnjpkGGG2HSrMNXr7Uta/9nDPOfUftespOuWyejXov/2sQq+HQB2NlXi/S40M
RPl0up70aPj6/CG9w7JwyFLqFJ2kMXesEt9HlOdvFcV6aKNyE4FivxpdtNzuOA5/
pQ3KrIEaGPWRFfTNm2m7pdhGB+KnRJE01Md4qACYBSxW7ZDbTV+ReMmB08sEqC2a
LRO1KTrURc7F4AQiMaLCvSVNNYnIM8B6gZXqzElFn+3Ljx/yqt4i83cfbnwRPZkw
vlbWAZF6VVI46XuBFwTg9Q7zEofZxDSLOTXKdNAfeAzQAFjnxFhTwUFi37Njz26o
VG7Hk1fN578LK4EQsks71paY5/g9LqkX2S6W0bV0AE2HcW1S541mSEO1W4ljLpKZ
NY7f2m152Qh13+oY26MJRVLr7/4lgyZO84NVwLYBcQDQM/rWu34jWbSeVeb7XqBd
myr05MYqkJgaWUKS0Cihe8N0LV87HZUBfPfvg2Krf82NL0CyYN1MdKRfwNPjwFBB
kaDaqlB0g9Ho1ZrvY/KnNV0vwcw/6F7CUjcj2GTCzdb7dmK6CQe7VOZpZypMH/mG
tnLOWhKfe+SsfTroO5qQxDUBOsCWUqbB+pi/QJayI/bF6F8djbo972VFZ1GgT66u
x3go4v5P05MPlNUe3uYAsO0ZCdKVPG7IC7ltvAyC15OMggbgvxKKJEaPlbVCY4hw
gmr5NLFM+beQXIzd6x9+iwIS0f4JZ1eymdD0IZe5FKglGEhA6LdVPRu1AlZKxiws
vSLeDA97+kqSxYkTDaXagvcbPIgADNsOy8nSRfXszV7vuDDacZn0hjHtGoGPVXbZ
sof9coopcSMWrnRqduq4+S7Xpz606ex/Zp/Xn21QcoeHSOcy8i9d4+rzoFiyjrp7
LUU3lksQhr4Ff/RW7A+3SWt04xwujhSplqcJCyBkoulMGpJchggQOn9Xyn6/YbmZ
LvYZvd1meK0bB9/KqeWNRsdRJWAiIw+6GoTxPSUddvWfzRRDGkdiRXnproJsrHaN
mNuuhC8h6j12pInTn0jEmBcCSsg9kT4PVEeb78pucRLQo2lw+cPT435m+/9OXsTQ
E/XQJ4h8pTHmXx/Zg8M3Mxb8+CStR2owg98Dk4kvJ/xQZra9jAMfui5EgHpb6zho
cAGB850raoCz7jL7Cn0OuMK/k2aBn2kRfCYhe84ZBEZhcCzRV78KwP0/n9UP821r
6dd4GbCfvzjca2RRDnm0mkGlXeoYT5IpgEGeviogIrayZifChd+3POPuGab9tAzS
ZbqPfo17zM9v3elSfHFJdAdc9rBx1nAKVgeUnCEbxoimyjxRlf1bYHJLqPZTMI8Q
RCevIddGkZbh4ePlf6kiEuIYPxUR7qC+LuwmbTbZfPnXVKhLk93uhU7G70/RFoW9
gisl2eV1s6vxgmCiUT4/+IyGlZMi8UAQiGeq+fQiBZ868cOh4juV8iCbuHfHhZ8W
iOfjUzGrimHGXtjyCNlGLKpYcCYbU2CodXFo1MxQ1WAUHgH/axnOfIBLRx3uWyQu
VHbd4xYaBYR1XIJsD1yWMWDbukoaXmqE0PjR3Dkbt06K1LACHaFwqji2r4sQP105
FdXJfuQspCFP0gWNL0yxbshfeq18kpvLdwGWx4cHxc6fy31vsI4OpCKKvylRJGpC
LXnatXOq1mZNYtL7Nc0wVWXQVmDK208+/BpXhZjvvFXQ7mBvheC2RWmZZHUSdbP2
pNmrcPOft2CPxcNM66qGL7fnpfwkdoA8Fd7pFSBJauRFWbjcfQ42tMHOLrr3PZj1
pyg01jOWvaPP2mOsQ3SFPINflTQoAUvIqCLORBKYJe3fsfSnen4yrlc6aP2Pn59w
QRXInLBDrF/tkXeg4scE7fH1ByhkgJYW89Ic3UNwyTKys/uqVWj4+pBPy4Ww10zP
gomcSwcD1WoH3E9uxRBrEV2ZJv2G9g7+TuubUqis7QQ4B+TyOOXbo4ag9zvT9Uyh
AYUtdS7cQeETNlJjs4h11UsnKyREBEAo2yzgyMhoB11HU4XfCCA1DdukF0Lxf8hP
GD2u2sMvPrakhXcflO/AcRlNtAui9WuI57zdUYXbfscthaBFNAyxHcgKHLbSqSvM
yHI+woJhj11emytc6o3NLBUbQzo9I1nQ6S98LspFIkEaQGLaeuHULwkxtp75g1Pk
PuWNm3vtPeudU2Dk96tKp/R+lDQkOc6NLGAJKymyEU73IDhIksYKzg3AA0zJvGQq
Ck8/3pDtYt8goTZPG/P/1i0M62MPaqdI37Aq321ye40YLAeew258XOtrk2kc2CvQ
p3/dpq8v9mPk7iiKKHYnRGqW0+SeX0fWV+xmbPT1hdj3+8OIHOQzpAb+WrFWRN+/
IWPH+nCuQm3KYBCmOiw6okZ2P1n3bu9OJNqn9HVSErnBxL30uWw0kzryuHnISVCg
JxFirGN0dK3mnA8hnk65FbS0nvOaoqG5Up3EAvopPjV2ZVgJ6NUY9OpxADwoBA0e
N/khEEZQ9YZj6RVo866rdNdfubVTslDan+EUzPuMv07fOHj6JG6tUFVDzaRZlkWa
rzVjh7a0u+aYwEl0xV+6Gu6ZJ+4NOSUAUSQ5I55IUIZ6g7DpsiZf0/6/mLp4Ry0V
KKHkJScE/n7flMXCWvEyK0f/aOcnzbKe92KriDuuuRJWkQNwc8SqNfS1c6QijjLo
JFB3nP+5f/DJXSrm6qTIqMJ0gXXFT16ZUr16mpAZNKEGp6R75EF43NJTMH7ZYZI3
q5XKWJSb6MdZMzfV553hmIvjc9zrjRX7/Ah0ZZiYXiO8tF93WDWmfH64bSuinlhM
8kRhYUAPpRr/bUukMfmPHqiPHTjcSppNAhk1pGqurbYj7ZhyYEDssvpDEMw+Yjb2
EnzXEJKCLDE9P/FNNYXXarGSX8wPAcbeeJ4EQMdxS77cLMpJqEZxQ+Qx5zEjcXiX
weruc+3UfsQFFSnkKLvGjNmddEsUmawTP3ruC/HhVk2LLKAyBQ4huNbkCrj9aJ3s
TCIeQCzvqOSe+mdZn+spKVLFJz7yIAJWIwTn9Ye2aGic0fw49+lyY6GMMnLBRpZP
8DO2+CP30ekcFBJ44Y/o0OeU0G2xsVCkq1tbJK7G9sBCyLkM2tbQfaqjH2w7D/iy
qGYMAOXuh/WnPAZ2oR1vZpze4KgKRRsAR5ZSUnc3AF+RajJwb+atAgcxPaz9FfZ0
RNMDzZ3w+RCg2IEBOCevPLdDB0zgq2C3h/e//If2OVgc6KLvsQ4yMIrF3/hWjh34
g4/KU2QOkGk6KfJ2tXrierOlPbcANK5uF6vJTycux/wetBbv5ew425yUBEr9uJsp
Auhf/p2+L2qdm98DeKUhfJE1xsB+U2TrGg63B/9H+wHVzWBgrmXSlw0cp9Ep4Nqm
9gSpUflePF64Ndd6ca185Wc0Z9DGNjr76YUAphQsSAz5rxUB6rWWY+VrFh278Aro
J7vklpWgzPFn5DNus4LP2FJRgBCT4U0A/InLiKhWiWUwp/SFTY0KsK3zOEPE/H/t
hyrzz0wDwKaIHGtg/ZeC5anpjRNXTVHcnrtvXmPqepnpi8ywLw3i201kSQei6Ezp
gQy0SozVqNCvS+S60UfewbxV3PhFH71RCJyPlMl6yusqyX/iGRIz27n9pwuM8Sj0
xFWgYm1L3qn/Tfa1tmzcjkm6U1B4XW3HJUrgMJOenv0SQZ6RL1jxfxs4477O1P3H
MNwqjFFC3MsLgXGz1WJquLJrmxbl8TDPKc+PasErI6qTSMo2hBdPTvHD3LaSFdSc
EefmA4q3rADzVchF6PxhAtBXxp6Izc0q0nPO2Jm39mhjM0ucWv8NFVR+ZElNBPtl
bG5i0IPCLOGKBxk6DrxNoQymdqb85Q0TYXmDlBI4wTOsipFeM/HcMlbbfFtmixq+
AZs8/MxBpgqjHb2BL1OAPcOkecEx29+3Q/zKX2nFLZgkAT146imlHNLdlrB+PAzl
3/n5DfrbDUlBFIsucjFi/MdBy3XejSGV/KMNilGcguBP0welgOj80A+5NyrB791H
HqPEGEhqRWyUx0clG+s2p6UllV+PnEUu1Ry5EEPVSkAmrqHgcxp3dC0A8WjyfIaU
zsCLRRxmxGGwClFxBuAOjEXnLjDl4DHb8T1AsDJ0wgu3C/FNX88RTjCbd3SCA29Y
nkBUw8WCE1siZyJKmoW9yyFM9OQ2jbUsEd2mRfQvUL13WzPbYN1iDOPIhQIC8Bo2
FyzpqGym5VySxgXBX7IJIHOg9IGo1hqIpwRo+K4XrUr8/AxYIOxT+IPm2Jl51enI
SU0XH2Wn/iNzdD8F61pa6fBomjlAm2Bi3Oe3lr7zjokm4et1OKk9PzYq5hRpgrz4
ezIR870lau9aPlLb8aV1gd7+Ic6XH2uxI+pKCHuZdzphtu/KK3ia7gEjPXyccOuQ
IV4mkEEfaQ5xV9tlce1FpJySwQPLxEUFNXacfdkdNaLPQO8ZA4pMf0xYfgbhnPUW
68dvhjnYRltRf0lMzv1k9JQobmjQhaJykSPkTq/w+kaJCXGLgIqr+Sniu6apy47/
3ntaAdZGNu9rD7g4GJFVIYVPbZ/RkFuXzocilmdkCtXq2c/eplREUOf5jFFwNNtv
5NBCGHIIobAmisltNklvHglqXCTERVGzoEfiwHA0qoGkf5ZAwIp+6hnsyT4vd7Gk
0w1h++fnLa10VnprYN7TY9SvVJHmU7gY4qAR1QwbQ2BfjX9pRSAawJU16d3Z/B/s
YypmLply1QjykmGaNzJu9OayMXlzz217/SmQycc2dpUU1MONRllHUnVYBREt0QGh
1hf+ZZDv9i+mhb7PyoirfsEl/yP24w3R8eS0T326dr4G/hIyKVEmg3JAvwluoZhp
Xt4u+nUfSzsN9k3JjMukqUKmN6raXFxU0AEZeJCG4ur0MHJ3o/oot94fFIjms2gc
WDvAbVBxSAWvn4O3UO40f+7+LurU3r6eatdXAaZurBIuoA0O9qsRY6GdaVQJ8whL
++k8izLtTVIFLCVYH+B4ZZSY4k9Q2mlA3+thhIQhRWMVOP+eyx6ZLmKHcPG9rI83
RF1wjkElc/8fJBTLsZjY0pQnJ00XwA3GW9FnbMAFX76r8GC4U++bwX4ej+zueOZ5
8jsd0kUW8S4YDyecJn5ndilE56zQl9xrUzDqesnpod1FPdx9HqGC42nGES+Gtq+1
rsQ4Q6MpbvxkhDciSM47dEIXJBwvhrzyQ2AqmomABPqN/ppA2YZj+vC+9EOqrnJA
2oNHqvAKgrmlwJ4xsibBdiEaHph/bjBB/lvGUSRndFBK+3qmDI6+Y4i5FZe24nVR
kKMrAy939aGQvUwm2c8brxPUdqKlbVW+9Ptmvb4B14ZDMoSIAb3nlHYfqdIWJlnk
DTe1iwHKvyXaEEtxNxB9Vi+m8hKpUB5b2Vz1UN0mzcvQHtYVwH2O4M0wh2ew+Nts
1smekcBxuQYbtdZKoSq2tUoFmLs/PjLSiXDBVD+tft/p3JBG/5DAtglksyYdrNYe
AG9vm3N2sz9ewn89Ckmjvr7sgLC/6Ual47/9/3+fF9yO8WniPKP9VZhGLzTCuS/M
lLsp+aiVH+OfCTVFnZRejoWXVAosKq5hrI05/Mv1cOL8Y11ta4TN7IwEuotxL4Rb
WIgPjKGJ8ZyQ3sSSorcB5uv6ynjHOyBeA4n5RV87Lw53b//AB3EAQ0OynJqmdY0+
KjFszGLYhFNTufB8Pr5Q/rXA20ZS0oythyA5eRbq9jz/opla4RgshB+JsyWrjK3H
xOLTjEcxKcTKGaDVpvWuXcUX+2Z51zuXSX5M2Vd29oLVqHQJa6AGpxVDHln5zcTA
i108xWcNQtOvLB368oViCbBPfWcd36RVVlHLNwsgQqo2bYnJGbAIHObQKgGSBBti
jpYeDs5N6sN4ZV4gcp1FCNdNMzHUsTA7S/hq2hOj3JZhDqZ8xlWCcDHTFtQWdWLZ
GzUcGBg41h8iM+udeo6ejBg58u0AbeSoJD7MwGfqug+hTk/trqFN1rIxIxX6NQog
EMzKuPcBavUDMtCpXMJI7LIiMweNobkgW7d59mnNm1Kakae7DTS+scCEVHagPCb1
td7146K1WrpZCXleahI7hQoy2LywH/URPClXeM2/QVWaSxOaQkGsSeVB5GAmaPJC
SXLLdDy4PeBmXRqu5sdZ1QzVEc7E0+5iQTegiNlvLhG++wz3ApQPhkPcjpmOT7Fk
XUw5/4deK0wok65lwf48diXE124YEez1OmnvsSak6UN2yDgo9ze7pgeb1NRLbLYw
b2Jy14D1YYanCXnAOIvRlcbIaAIyAA1gkc43kg44sbcx8ty3tl94hmpq6HkcMRPb
tvU0cGx3BxetmfUCr5fudiWehIA3at9kMcvsrckPdSwWqOWZ/uC6aki1cRIiKEJa
+kXtaEI3d+mvQs1oGI6rLxlH7rLIpeFzcZ3hK4qI+irj81hx3wtHVORpwGTmKoc0
k/NWRSgnvDNs90hvcf861oHXt2Zddaq9wT/JNCjg2XMzKlVYXE1iLYghMYqIMUbe
mB7U0IyfntvTzryZxy6O2aWrYwApvpDvm+nCcfAcYU5+SHdKMae/0G90LFC2JvyJ
TW2caKd1Bt/W6mVWktCWAvJ8Mk/xacTPhDpbzM89SZ401QVc4/QFJq7Z//2iPIfi
+S7jyNo3Xa/ov4SXNpPoTsSDvSLOnNP77vbzE87J1PQpv4Dv0zNH563Koa/aS0bm
YmnYWrhaOZKZu6gPZreJL67kDXNLj8pTNUP9AqBaosQX41DPmakBDgruDbDjyYcj
ZD+GtTd5XQFip0w0V7u6zxJymRoSX0V+FwkvreeiVGjzwsqE8lLHh0JKaaE1xed9
/ifKOg6sY3MC+DNlb5ukLES80MBQEflbrAUrmzJAhYzZWbquCs2tCwIgGyxhpQa/
6OL+2w5O4TNxD1LCTAYY3lxMgQUhGF289eajganE1MstpxpYREa4BQ5gPGBnVA2y
w6Y2Diy/xqpVM8ZugKPYUv8n5jqfc3RIonMyG+NLPYY7oAdlXhdJq6oM0NWgRHoQ
tXBKp0zEdtiZ4dC7BYs+v3i2mi/sV4qnO37e+WzOn7Q7dz9EWXrCNBCBp2YVk1mb
z8S+LjXzDMxLcfdW/J1uw07oEBWWacEp15qKtv1oD5sMlyf45SEZawhkQZmlX3mX
Sa+0ecS0xr4ZaX8wD3Fjsc2ZD5WfNykSCu+XTe/QhbFmN9ETRaDjDPg8XX2i8k0+
fpaWFsk2Gn/49yr5CoBXtvIGf5mO9u/6SyaRP2aK095RETWlp4LQeLwMEsqP85yA
deyjPUECzusk4hOZ5ncXIWsjt1lx0ITlDUvdBO3iNE0XJ4jvWZOxxbntV2zkO7hw
AQyI06o1a+cFnaOZFPZXYfRguQ5T8DFU7uNt6eElQ43tkLUhveCxxGUrHtBZlL82
9sRdiSSvtxoD5aCL7DBBXfJ9uI47MOWgjt529fUcrDvud1GJR8xMbmiWjoAICRsM
fMq6vow1U84jQQR1au+I/R1vxhG2Jn+/56+fkCTPs02V63Ez0wv3FRY7K/9sj7gO
avo7WI5kLJHReKhqMoznrwwD89bWnyNBWBZ3T4tnYiuYlJGP9TYtS/TFqdsWnJzc
0qLVcH6ldR2JWMmofl78JxXRUWufmgtEdcS1CmqpcS6w6gO8VD1dLHM2f9NJbBiT
iZGlTU19SYA3RFIVSb0fHULNKqYJpbpdeTe+rX6MsBaW4pAaBftXpv9dtCHu1HMH
O1bxoyCzz39mj4Gl6tZFsZ0npcDgsDelM7zfhAh7B7QBvQfCQ5HlNizI7eNMxQdm
/jN+I4DpeRbBWajd8voVBvbDiTsUeVBVofXKTS3k05zDzhAtNGM59P643ht0M4C7
3W3ThwDHZE1JWFIvxK3C4B6siNL3sFLGZQR3/0hmDRHPn4sCPr/UVfkk18UhM0W4
2m0eLU9JfXi44b6zwJjrBoUsFLdYnZQ8yf0DZo5ZO+7xmH7KCWjqN59IoyZhGep1
m2BLflpesdOuK4oZqzUYehYN6gpmgxpTmBkDKJabKPyMFBugEGz6pDBGSeap02ci
78zpPkH5DKY+aGrPZcldmio8mmU7EguSM6g+Ym0qlv4WzkUy6D1QbHe9gi/0SkFH
+PM/5cZ2wcRNS1JF1M/ijCyak7QtLN+/MRW2g6P3e7XSbu4ZdTdZTFmer8REUCEc
TVkfjDxyDSa67IDcuoR7GtwpGHjPBMtvM20GR11fjAiZs28hxZUjy1ZAwvnMR0y5
NfmfUzuild41PX22QpDGZFfoGM90FNN3V7Q32lSDc8Abep118WbMmhrh59YkL/ji
xkeL5NjDt/9aZCS/2EJud9ym4trb51pgpEE/YVDyr+ybB7AAtDhgsfIYsAqL1L6J
9GQ0UZPTEVNq4oAT9hrwARvEYmoZx/7AgH99zHIrqaVIkWN/V7yowUU+K/L82E2a
z44CuhFW0peNo9AV4apGhGzq5aYDwR46ZLlq0jUweT5n7kwomB+HgYWq2sndpfVr
B1JPRH0H1Y1olnrdYMGzrd1ligsUtjSLJj8S9Ua+dLaaXck1IazICjgkZR50qeg5
+H4ZfKXvDLx1omYg+jcEqQ4VcmMS9o67vqTnOhKHllC8TYa4UU+lpKj0iQhQ3ef2
4ypWnfW5sVnZOzQbjvCWNKrh6WXUImLFw/H7/w5TLYD3874FCAfRkfPzakNSXuZJ
y6VoycqKySVr7iUDMEbvgeBx5oLiAjqBTv1Y4AheVS5Y2H3yMkgMQcSnBDZULzbA
4pEwusq6/9kWNywgIUDCUTYrUiwteD9Opg/0Eoc1E6fkXvKCFjuAwrpQJ8rHvbCE
NEEhVdwqym6IAGOejud/Ela347cTndk8YDAmNe/Vvla+bjw/N1EK4ubOQ1DoFKQW
BxaHqKE1//xqwht9StZmMwPmRT7O9E5ZuPhVzVIYFIitLd0TW1bB8LyorunD/JuX
pEgAjzR0afygrbe78oRJzYmZ8dcQqmPZ57v4/fngvmxjvX54D03mkENv/OE51JFr
fmUXVbk06QkEtwM6j3xyliD61nVbKFNAbgKxKmUYE0Y0YE4Yx2tg0rIoGaq1nRd2
uSmQg18xbSd5TECkn72OXmix9Bj1QaNrvy5UdD8Um/r7NKRcXR9gTobqAROyhvCk
sM+mE8C6vKCKZVGbN20udEwNqxpwDQEoxr2qoI6NuYo+DDZyB/sRdRkn5Iigbk8R
SdsGL7BUobhsFmAZF96t+Zlda2QnE07KUD0GqeGoEt7EWpeJ8DF7p8GFnBTbxug7
lP/W3K4OKmOgDIPxsOQJbaWGaCaluP7wU9EX/2zCJgf/QyM1poIITLMlzszKkWNH
YKerGEFc/RbOu/SRj93tpVaSAb2XB2kQ6ehWVw06BYh8O0K8qssOBdPSbIRzhdH9
RV/KPgGRGTCxWarzYUDi1xkt832ROg8mS5qbGuKdt1Nl+gPbEqtWwXQJhHTSS1Jy
LXzQJgVdpzrUtAAaOLRtf6gYra+/GsD6EJrVRoLRilnXysbRE+6kdvihyoSoBNQj
wmPoOQg2qvzG49bOJ10GLdyW5dBLDMSHOr/M25BiX1XsORZyYluPVEPX3YjWb+z7
S1h/s+16D+nLhl7vvZ0Bs/sXSzznMiExlnSYThbz+qw2vFFWrayHforPgw7x6yEF
pzZriq3RNYfxUpe6qOYyhkTMBCL2S1E+MYE7RBdPDcuQuOBpX8r6wdqrvpZ1bAAV
0wTF03aKBsHD3Q3mo4SVQbhMZBeAO0aVv/t9brpVYok33QCw331PqXpLXH/gyKza
PDEyqTYFW8p/CE0WUfAdKsPrxDTPXuQMMG8uLvBEqi4SiTp687ibzEG8Kx7aeJ45
mKkUZjV3zUIdiWOUnj4i7UTBwRF95DBrwjJ/l3n0kIcx5kd6hn5rkXZy3/4UvKob
bpSLRZtPAq4fkp3xejfH0+OLm5l/hie4Lnj9kxmNXA+61yYUJtsSlGmXGCK3gF+V
F7GMAp2dAZiO0mmOb4C8dY9sYOiOIoLfXlaamhHBs6HHAW1Zi8RUiUmpJ1l2BNC9
glnx/klWrAU6TH6pc4FelhlYgB7dT0BYc4r+Yht46z8ulxnzjYC2MvfFwvbW1h/P
7f76I5F9hrw03VUlinoXJt1VWAEmeeUfUAGB3oTBDOAVasbdhlD3GTHak0QEHHM3
BpnoReJkm8v8mJnEvBoF8lgP6baBBfGPpMtPVRkp1ry5R16gmgBnlJHS+m5qPlJk
JTq0dLQ/Y1kj4fmev9WufKEHJ0hx6zVQkg28lKTNtpjdoFhl3HSE9GQLB2N2xFo0
zZZC0YHyfhf+zF0rHT2JjBlkCCQes7il42gFm+qwMuCrN0MdCkv+oLoU4IuDxMy4
cVmSqisiXzfb0JEawGxAd7Iib4ez+fuF0SrnQas/EtIPf3FN89eOtlY0EXThy8nX
sFJBucSPG2iLjp6Y4a5tzhogpF5tBgqXNoykrcXYE77HoGVWSTT4TvVPyvW0XH+g
fZVkW8owM6Kyzrd8osG6VzR9irpgvmfLO7z5hw2MlzK1ckC3SoutcokN0mT5n0+I
rdHTE80gew1PW/D/gbvkF8LjDp1Id5nPUSNFJndpPCLCRiBQpM8eroFFEoVf1VDu
i9zPYF3/ssC1kCziYNkChD3dxMYlsObqf76ObUjrEdeez0CJU3LIdR732K1GgKiV
RGtKZGAPkfbrPOKoEx6cP+kyiTNfqmVrez4ZOZE4t0KOwe84kBmH/AdSeGbC65dc
4CfSoCAGP6ipz933bYYGaEgkZnpWwjq1W4zvnqiS7HSPeOuwMYrtdoB/RaHIlYwm
PhwkwvuqQUKF6Ko5A3nuuP8lhGKLx1XVPTswpcCxWvBJsOB7q2i+zDP+fBeUylKk
votkhNqInoEyLWkCNWUpDeIpGG+/pHWmisBBtDp9CGAJ1pIQQskNfWOmN0fUcVz9
jRa5S9oIWd+5BQLCLttIGzLUT0ML/I9zVeDnlwWio4jKrjVgywcOIehzsumqPeJq
3zAVhylIDeCdFQUMgXFQNQV7/WlBfaKRwmoyvBRXFbpHIMtpt848X/TIA5GArm8H
tyA1aRAv9Ze+o6oJn5XjrdoXgZtalyE2IMDUinhiOM22d5+6Grx7GqTb7tqLhC3t
9M4T7jkIMhmys6sop11zBzKinwcOW0ypU+QKB4rg7GJhyybIwsa6ZYSVZhcyLv+y
y0hKExIH57cQAZy7yFTmnhDJIqr3jG8t+grzMLCcNd09whM8AsvE0Bkvbfn7nvfR
eBUwQDSkjmLR8Y8hk7OTFPROl0gJuZM0waQfNXoEYnYeVqLUj12uv2yi9qA1Ebjf
Nk8H/VbdF1Zg+X/mYZ7rtcyOSIbHDZlIfrMCRu9I0gJeWMUfG/AqXxMSnSCveegc
vd02yomyQvC2Nz5UhiuNniNqQkI/etg/RL1Sx3Lcgm7JUEYsed24dANlD6KHQLyj
DZFYcIykhLlDog5L97FkSKkunVAi9S4YnDabPkt8dUKF/dI8b2fK0aZueQ/psVJk
CbrXhrTmTadDSM4Vw4NZqXLzJTOPELoEdbkJlg7GeP4vPBrFQsEOVQWxdenEJkQ3
m+XzqP9CUrulYCxJYTrQRYI+oDvsO/XxGrUcmYeD2Q4aQPAKkXQ7fVeAzxDWFwtr
Y+rYpImnB58WeT0TZR38gSrXJHzLoEwJWNcLdOL4aKU3VhVsyNQuAxCStPnBoyaw
rDqkMMdA7cRgJL/vC8TJDYJOZfiY4KjB/bRZzPfs1TR6E8WT1SuUJuuS6uW8gdZ2
T8ZG7ivzbTmzheHhwQ/9SJbfboA8ZTClYT+U7d3Fy31rnN8X76fZXQayFC5uePI8
MIibdHom/BdgAgxA7pM1PiMGkbGCEJGOop3J5qb06Gj99vum54zdhLkqQtoGacwj
skYH7u2o/bOxx8g/IXwJL4/TAp4h4reXHVazCC1x8ne5KvKO0Wflkz72xLwLwG5c
r/0YZx1A8ia4pnc66cvfI13duTt8EqrlTxwWgLcHoVAB/hk+JYDIwKDfLEWVbXjo
ichHRsMHzIWgttK7iQyQrLoGiOiNGRYoVfU2wV6e9NL6CFow/0s0bGvsO1Zrit3A
bOyXmVamPUlLH1YWmB8Xu7aj8nRjK+NbGb80+diehEMfsm2+jAXSjysvMKK2Unyk
CCxngx9x2sJzRWp2DqsWuw1ILKCtxeMcOrT5OGi9wMzE+TyJ624BSV6+3u34j4Zp
tPsbWRknJcmMqAgUHb9cRU4iv5AEVdI/2q3C6DQL1P/YVQX7Sg3wDCqrGqyX/q9L
EvXIb1OId1YoMpPapfAv0Jb9VBmd7LzUyknJN4ZLDlzU/43QXKOI50byECje11mt
+eTxV6A5JbmbCzcXEGZzWSHZZJdD3bXcUqionCzlAUoCcZJp9DjgJENIXbKJQZA5
f8FOIgKQQo8hyW5sGCo5XORe7ToekVjvUQ9BUiCaq5QQzefdD2fzr7HFpkBUGfJo
RgOBBGFp5ReCKF3t9fsuGen05KSSimkeoTANypcjQH4sdG2ebJ20akEEnSAVmSz6
m706EeHVz6KIuEbk2KLCArZFxiM0g3vZqSF5uF/YKAqWMtjJr3AX3uJvJ1HigV5a
vIrGQuRvW+Qg+Y9CA0MNRflhuVx3M3BI8ySfPU9TQCBtBfGfQEM5wfS8ksFwpy+K
nsNEGzpfQv1yxltBGwSr0GajSJ9PgYRWtGkCaFjeEHvbcJWMEaEsxqujehMw/0x4
SBNFJaa5dnevzibNEqXdgDnjRvrhXnYm0WNNS7cnAuhNpc6VAMe5q+SPeqKgxf9m
CBxr0jukvB+WRHDKtxDaBxkiPGiGhr+6qHrLqQewEqfPwKttluhePEPaBCLCkdNi
FJFsnKYwPGuruajz1AqKNLcFIjQozqSd587tpj5K5XUngPosYGd750wbfIEBES33
YemyEMZayFZeM6viGO/ZnHTJ0idCyhhN8LhhYgz3NMPiaRzVH/YEypHL5ARzI5rq
5Nu67SXx7dAwNj4byix8alYF7X1wUPCfbZaKTtmLC/YgWGk9KZI7bgZLonycyJHx
gdkvjpBLHNG4tswYFyMr0onk84Meeqppha8yCVkuYIUwVBhnnT5I8ejHXK46zGvf
EmWfWDi++G1An8m5WUT3t4DicdwdSB450gBUbvfIrM5xAfWpqYhmCmELb74/FFPR
HhgrukpJhRiBWxjPMXm+KgANgwYxSZKFtHMSubkc64zhEEX1aUO3HH107qd+jOBN
0nPdtPA3cNfKOuLFheU6ddFJwgeLkHab006Fi8hH6vVkBMCRTZN7LV24yt/UmVxl
fmFPSY1Z2o+O7PvnYEAVQh43MKGsPsv/VG8z0tWfL0oGHbH9mloJFqZC3JAvkTNe
OsUayGySYzO9plPeAKH+S2SHKrad0r1x08S8TgPn5EMT6gFNn2rsQPNa+ErGQNvP
sDMI3zT8GGmLp2UrWkEQYC0uIhLzOdCOHE7sLz+Ib8VvkNoEGUpaSh90ta5Jtd5h
WvcuoMwVa+cLHPb4U4hZcDOqHl+qAD/UsZjAJYc/gOb+h1HPTvlkl1DrLDZxM1Re
mfnSuXGGYKiWrDipWoXrnR0bUUYOXC4nBQF8oS5t1WfY94ddjlh9OqQq2/5qgA6s
n4/jPBHjshrDzqJ3NiB1IQ+hocqKcLdurSCZ9oikE933wW/BXPcnl2R99n7/FECs
dJRhj5m2zb8ZRNs77FGZ5NCbSMtQxrYH5VTFA7mvq6Zp16FqvqLkplsDZrNUGOyU
Z0cGkmKk8TQPX80owX2P3Pf9uuNaYTnUL2+esqgyRz0TepVfr4SbClFpDvWY+JNp
qOs2emy0zhQRXa66QZ+GQ8rscTg+guU1JCuUdgpNwIoxhraoFfW3xwBvlvTmOqvj
YxdA2gtIR/fSKaRvbTV6Iig5hd29C+rHWSacjd4656silyxNtriJOaw/OC2ToOlX
o2hOMAD2XpGPVbJntrKGsjMykzRfj2bXEx7TvkrmvDPLW6h2zPZuuwPFNvS1Ygk9
UTDS2NO4hovueATNovqHG0lQtm99dkD0vLjSEbjNRGixUCzwgx1gji+0s/1RDnh9
jckWu75xitVfk2Y32ikGPwsmoX9bYD3ppdOQ1/YTEInfvY7KSiiKRf8/HwKjAnxp
Yanm1h+G/BAvym0AI84GBK7tf3J2f5mqWIz1EVhQo8U4QQrOnoiXbeSPSotWmXZc
ROWlCKTqAdqMdCcHfFx08UIsYqUau/bidY3FlDsquKe2Vkg0cvV3ECTGNLXycX2S
H4Uw1Fg8/K6uXGsv+vQfG9tccbee/viFHewcPWp2J0dSSvl0PC9is+baF4vP2W/Q
7sGFsQrXgUi4vGoCduApfk5wkZzLb5n5VlXZ+H3jPsXYuZiRVUFQlPnViE24yp5k
ewgtvMeVb2mu22DRd0EYkSCGi8bd5lBpsNCZ5dRITx3eRnYTxss4tpqdlGn+8PSR
sskX8DOw+aFVWiZoJ6dwO9GH9E2mm6TKZTDckkfOaWA8xLY94CY6+m1a/NUfRmVM
7Cd5xsnamoey7T8iuVN2HR2RORw/ZVHyH1u3PEdU8+Ez0O56ZM7XL0o1kHduEX4i
Bif9A5Z6rOdqoTuS6oNSxbFfcQY6ROlQg9Sx8Ss9K58p24hHGReFTEB+ZsPOEdO8
1B5FJ46YmRxK9fvm75IY7bFAAgAWXDmfdiWPYWUdn0QDLF4H4Eg6mZcpXPZ6etfe
In3GtNkc/IwJY52yXIc+x0SgSbTo0v7zSXIN3Ze91u/4XxWO/hnJZZQtiC4HDzyL
5arVUs2BHsU6n1Bps5dWYLt/sTaEakU7dpoerqeK5zknc4R/lf4eykxmCXMgWnTy
kZMX1lremTNYC+gc4fN1lIxqFt1jZumrERt2grsMy9sPVw9itY7DmTAI2RQAgu/E
I/CgQPLlv297P3kPywJ85cCh4qWG/NM5ZHxCmf31IdiURQMw1K2hx6uh0nobgSAN
6Fzd5jK1+Kmg5bAPp+FYAAOALh1S2QhwZRFHFc4zG3ysOJl51AhjUz6C9AualRLg
kdC3nAeaYCGgSvPOVyUpNz2A/KAT+h7gC37cYyxK6TVW1HYx3/ybMliNKJxyfhgW
s4Dd8BqdosuhF5FkT5LRK9JORjGIsjuS1q5NtHfLlWkbBrhD3QirAGpT05IN54oL
uirLBSRNJKucAas283AKnGImd6uK7BLQb3QSs584pBGhTFI6KyfnLFIAm/aZ8FxY
5ghojTLusGOAfW++WuHBTiIPI7U7DJ7pSRYZLQXnVlw44lZoXbDM89YcpI/BmDQi
eNy1AghnVs5mwroWFqnrN1chfk4Jlhhoub3EQC8uhnt7HYojhvmmOFskapfuLZiT
GmsoXOnL76cYbj7jPuLz6R3h8XrQiBlitMSJkjRVtaYJDqD/WpRWaMixIQnmR4zE
Zk3oWgL2G1z9O3AAUA6FyQ+Lb+/P9v646UPtFUiS6yYdb3/zOEDm/+WxYckL9o63
k4PaGHIBPh74yT5IXfmOfGqYLGat4nOBEDIfrLOURp88DsZ+8ce4HpjGacamMF1/
6+UE9WA/kaZB01+yYVsoo8oWHreQkL4DbyDGJcCeIpeWfzxBPTUOhBh015Q/zmxr
3qz2l/XHgw6oNp+JwKmsH2V8l9wJy31DrqdkxGJQPc0opNywJ7byPanL7SbKX0sd
AzMvP7IB3lN85Jdbzf/6Ylng3Nub0iTkbCMmanC65At8mxOEiDqpj8hYFK3rhiVk
7ib816Tv9fDWMLwQWGnk1PkXeEx+VkmqrVMv/F45PKp0Q/H5SrCEN1RxMi/UEx36
F4I0jA/osY34CLgAFPUqRG0lhcn/Lk+2LUqVCE2rLvhXeIwYSycAbDPsf+nRtoxM
9nk6Ao+xCWfa92hXhMS6R/DHDiPJHr42p8W7+W6XpqWrWILmf5cSNk+10OQxnhjn
xjifOBfS2hX/FNXfUgYIW1IxvwBzthIXqfgCbLnWJQ1uLC37GkSRzzHBvzMRLDG8
ZGc44HQzE3hug7w84k/IBT5UlrCIe6aDijBqM3v/823kK2U+4Fa2SOVJ6HPBYVLu
7pPld/8yUCoToeMAov8JE3zBzatlPVlQ4FhOetQnz4djXt0x8ZYzb3lK/tbbZW68
cIzYpj0587Cbkd0edqsvY49LEMCzc5ln+xe47z9ufpkxhavhHi8fYY4FvAyi/j22
mrwvIzy+EW+qPmYpr8fo73x4WtEcq/ygVAN7wv4bWcdwqRnrgtctssgfJxcXeTzg
heClRahwljxjRXL54PiqP7gltcNjhkRepxlp03S4/SadDvGB99rpqIbJph+HIFyO
ohB72MSEU9QRndLnGcDHtOuLK01Yl8UgVPCjjnKaC2YEsqfyuzPLUcSZZaZAER3c
88NtzxLONMmPrgP7XgEJrTzHpqOp4O5c/OBSvZugqNFuwtQWoO6OL0YaB35JY+M2
DXzBCD1kZfwdGwM/te9V5Em0+3FS0v/6AtPNdHd3Rw1gWP+Pu9AKgNS11yyS9eHe
AnEDLa53Pk4RbkVm/4+StSaIn0x4+h+xXJvwH57iuq3g/0Rv2Ua5OO1sejVoH5qZ
UWTQCjBrvrJHLPBFewXahFhOY77xCBj4mJJopy7o926nvFcSYnWmeLaXQcRNw2UP
TAi1TPLIPUf1WoQDI2fZDieTe8zrqXXD7homH5XKcE660aZP3V4q3NPOBbCMchr1
fDPEjWqHpW63TBiOdMm3QrGm9aqHTVUCRhYV1saLM7FrOrTMP/7Kh6jc6N6kxVHT
TWFpmFsY1IP0SwRczA9bjOamDq/Wglc+HuAsVXEMYx+3yBAO+TMP3MQ0PbBafnLU
i/ZU1ORYACLb9LVtrKdvN98G1Pdt0sHpZdpSKkMuXbKE5DIHigaOX75QVWcJsT/2
J3I+Ag2vN7FVhBeET6nz8v/o21ubHS/OEdmOpQf76OL2cAlyFh0w02CyAxnUDCaZ
BpcDTbigsr9Yz5P3wdAhkPtGVDkuQFWbrin+ClLHCpNg1KlOchnaKzteXGgAQTpm
trIzu9rPgPc2nNYtTJcfzTcveVuODLtoinNB90x1ltfj0mzL3QvlWDUK08L+ssUC
Ux9Zt8KHu6t5EOv3wOsY7BCpFH5qAD4gpC433kdqlD7OcVVwbqVXvomVxYfqOFMt
el46He9CaPHv1m2916A2RFMal5KKfzVinujf0vgYg03Te00SPTW91o6yFQALrMYl
RmZ5LIwHZwQ+vCK3g0mZO1bRVKKdIusC2JLT02OroFy1NUMD5q7do+IfQJCcEZ4T
0Y6caA/GOyUdFFKzDccqNa7Ie8j+EDE4m+lmBRmuVVzXE+hKtMNWGltiQGyIlSlp
W4pnfHr+Lkv1C5E+7oWZXd82FXDb8Ne6fdcAYST/dhn4A4f2Uh49nM54uVJd8DYA
1lN6JKOg4gWJyQNR++j3bPVKzZmvD+Ls9az/0VjDlWKHro8EyCaHUuMefZyEItJY
wEybvyTDymFZer2n7KVUwheXvAq0TH50T5BvhH8u+2/MGvyIiNsw/YY1QXkbildl
JiiHzSsIf3i9lp+jqYVICbtQbm4p0PWamZW3c8UhOcjyuqQ1k89tRFGePbcNTmjG
AhmVLM424S9A90Pm3Ij4szj2mII04Fl58KTxZc8Y5khl3J1mQqgp1pGY0P02kI9d
qpp2sscLQ41P/NlZQ7GTFDj0+DhFjekuXLaNosaas32Lh6U5pOjl47Wsv7oE5Vms
AefnYL+fI4rabQo1Zd/6XKe9+Zgj5eeZ9pZOMmSXNvUTyVQqdnGGJKdzwGjm8yl/
vHMBa4UJcxV4gB+wdZb+wFFbLIkGEBYEaCSVO5AR1pXwCSdHy8hePF9suFII/rjh
ftfX/btCnckxxApqBfgQ9XDFpgG4obwmsfUhVOh3ZgTZ2lLOxZBMqme3GKFLmkqV
ARpdN6vmXaAKjVDEBAUGjdyVI/xaqGhzKQIPT81OkS6Z23j+HnEq4GYL8l1x14rG
T8WVe227CqpCFqpBAOIWjwsx7I5yds1YIKsFMgwtv5Zy8e/bpuNtUBNJmDFSQd4A
v1t6+sRg7V3rbh2oUut8KkiX3zfjbPc2nCfa7NvBz5sMMrcUoo4v3srCZ9eY5N58
1IoiVP/I4L5jj7AhbY1dPhqP23PJpYQdIAD7exol/pqOTD7voCpnWQOzJlIJBzr9
uETZcwhG45gDJUJiox3CgWfDLMB0inr9SsVVPz5TrwXjDoDBl+0ezWQML7IGCy60
zY64MgdnWofp6NggUnAJRhggUoSRU/6kGPJMYqW3hieTcsdMdCJ7itVyULG0TxDY
hoV5sn6/7cXMLYhZyVD2NK5+godsYNH//GJzt/upXK55VNyrN7YA2A113IqArOYp
wQq7XjnjXcmc/7nch+1/MOeD0fgTO691DFxh9hc5YC8W+0hT4tzmkTe70ySle7f8
ufOM5S9DysivFziJxBDogBSRCkyBRjkwFEBcrWPtngJxd0cxi11jnDFtYuDteopC
hdw+vhlayRZ7ZmUrxDH11cTWB7VCLqAzgCiyDYCR7XHD3D+sFbZsaTiFu9AvdPjo
dlJDwVhgXJ3icRhgFKjLqyZ9hQC71X6EMm2CAFuSjqRmbahjk9b6cSDdQgcrWVRP
rAWLrxw4spEjAxVQeJubmvkql644S67xcVdkBJ2iqTHN1AwC5CgEGox/3BnBkp61
z8h6Ap+m1Gj3SCjB84bpqjIL6Xom3MtNMF8uFVf6lvHRIjFAyCME4BpBdFc5/0Qn
KR3I79hRzNEimTUI0LnEkpEipKzg16xNtGwQs2BTghBMX7+9KGVV4A0E6/mRf/b2
Grd3iysO3VBLn7ESJb9v+1BnLcD9WiimTk/k8R691DfBy8U2Vviye/rVrq4yDx/s
4LVJZK6D0HH3DS35SMMBHtJjZGuZgpzGaGVL6y7C+zfR7eVSzI5WXuZdRdQkQ0Sj
s+mAdtF4CZiP/E1ZyOz8GMifnMxPESbM0YBbhr6PMcVSP3zSFQ5SChQBDhFuzI8F
UOQJLo4H9gem/3QU5yYwFUpqzBQPPJtCIdLuP7GgBDLZptbwH+x/H+RqF2kOjxFy
JhZpDa+T0rvtqaRfO0ccGwLCyshdOE+m/Vuzkpyq7ATU/nuqnxRS0YK29qBRfl+f
L7SDq9Rx+CLezu5PVjk6L8ojX+nnjuEhCSJ1qpjRB7+twpZSFhfEqGXBlXfRk6pL
eY4Ik42kIj9igRWbhcTkJnLcOKuSwoLXFCz/oZZRJzc9SOpo/TyrgNmn+JnZaGow
17lncmWKcFPcWRvkRNJckKNOAMfgc2rZ7/OkDgpQyAldB2Oie2eVL1Xc0xgrIOJg
DxCWNldHOL4HQpyZqg/RrFGo8nocV0wptBvTtaYB9s/rZhwOPX/uaw8WeuwVH4F8
SmcWRm8wqj6oc5lLnBRukSSGLPc4WBeu8M410gINdloJGJdiaO+o9aYd5xyqD4QF
/fIWif3TQ/Wz8inXzJYjuFPxttcME/vvwLn/zW6WoolrBTXFFlmGn/r+zinIUH2U
248FkMaw0QeeKQZ6NQH5GgqdSWuK9gp20jFo6LdhzNRWjcryiX8RwJxVZMqfNfam
Xfgz6PGr3JchNySQ2TJ3rJbiO2de5t8hF1rsHumuSTgfcDpDEXKKavSb7n667iAh
M1RDVumsxseE3tN4TsYFqVPsxC0vJjKsqG/uwsvGDFoo4wQpHG9SacnpWrc3hhYK
1xadPc8BoeonoTMPy5nixAZxqHjUnJhmETx31t/r0dPSYYPEI9UKUvPz2LzCEvhb
VIcGyuFCpw/e7tyCHhuh9EGLOzA+kpoewSOZ4vsIgM3Qb7Cj5aDmJ7vCHful1Jq2
unA6S1NIsrUcOLKgwc0q4ZJZzwJsDlngmRdTeIJPz/KgfHcbiFtvcWtYPh6FQXeJ
wdyfukKeSuke0fx6I1pDHtDokQ+twgDM2v8oLSrlZIz25OCx/R1b2hNT/YUzs/BS
4V6vvvUVBS2am3Ya+UXi9dZ2jIVTIucuxqQSdm456uLbTZXbsAfjzrqHS7td0/vw
XjToS3yXoSb78vF4ZFwnQmRC0OhdnG0uCoC2xa9ftjtjOgd/cmH7FBfNKdyFFKAZ
4QBZ95EDLYgsjq3Q21mm/C6B3CK6j6ue66V9NiqdfXpxoa7OlSBT+4m2hHmmlmUL
+Tsj7MI22P5UKjTcf7HkIStQq8mNsMi0Pl22nmA5wi8de9moTXRzYipPra5chTA2
iY7LTu/GM0JJZIoJpUZpA837kTyh7251Iv05eZUCVIohbTGYAxq9ifbn6uqIaAm3
TYUPR6FZppfiETwk6BhDSn0X/M3ZOXNjvmkoS2mDTJ6sqpflZM3IFOr+u1J7t+22
C9tFFlH2HdYA+jQmtUnwXWtraBCwLybPygPxVvirt4c438FgEnx6BjPgzzxPIwj7
cTrJ372wKovttSarZw9WiUpUJ0nnUKSCbaKbYGZmhQPDun5iT/K1NB1PDM5Z3r7N
utLXioP/HtP8seWYrwyMrBC6qhjcdZZwaO5RITQaEsJs034/iNaetPZEcfJfpdcH
+w4FsrEB5yJGj+lga/15vsK8s5WCcGTHScwCEImmsTxOCpmZP/4Bsm96uA+pF+nM
oQ3SaS7qU8kdl7E3/aFHDNvS3ObXMg6BJLy5LxuaEyGIPBDzelWjxyOO9yoQq/40
YQkLksFNk2dbuardC58JVP5x6msegVvEkLKiq3oIyMvM0blqhDGfHVexlipIIFf1
H4ydb2XMogVTTi6ORxA3psKfCrxZlurnhiF6aWxXz5SAi8SAS7jif1iZE1nLnTGg
0HoSLIYkE9zqI+Jjrxsvs9QbxzfABCejcdB14aGUJqbYsfi57KsWNWSHnPNhKbZ/
GmWGp8Z7BCd+OwiUZxk+6jt/guwf90lKh6Sx7dCf8fliiNoPwQflqh8IhVVADNVF
0GDuJ5vJMcdjd2cuNt3Z90lZ5go2SQKQh62NRalJcBOYUZrkv8hxR1mTwd6FR2XO
7YNzxaxxzuo4do0TsePowBWhBThCLIzTgWd52Jgc+gQIePG14w7n1nlpp0DBbFXF
76qwS+VWZ+Z2zY1J4pE9R8Zbon73JtDr2nQp4tZYguGi2Z7kRUdgYIagq822fpHd
ZHYiTBaQBZP+V2QqwnCf5zy/vDgpxgfEvdI3KV/OF5aeGPNIUsqvIJz+qcAl4GqZ
LAyPh1buoyBqvVM6DLLGreJT6ErWwinQaC4zIOi54/GgwZDZJno4R+JQWJ8f5IVp
L5SeVKNijNEerzg21THwzoVcmSXqu4DYtgQdv72iW2/y2wefpDa2zmvXIyePKFlA
KxQSlDnf8QPOzqyoD6YHYNSw43/O/eIqC60vn2e3OI6iAlifSkD4jbI2EGnyjAqt
n5VOHo73v1tdPPjm1kCShG02krsvjYsj/094eY6md89IOTFuNZPONX45hMAWpC4h
X3fqZnnnsyEYF5aQ9K0nIQk7Pp0Tsc6/GOCI7dve2oO5xfXiS1zLIAO4XPYZVp20
/BNK3OtJaK1kbD2XP3uY/tAxLvoF6duFkcWAycCwqdAmwu3pJ3KUBZWMMvuWwVNr
ljzug7g+YAeoHmfxDyEkQK1PcrTRZpaSaTSiB3gggRohFzOrIWYeAl7MU+5kb+LD
yPc7rKNm49evMrd2qewsQSkKAZY5S7lXcTk+WbbExqk9P7ceSsNrZzXZnGxSH71H
sG2C0ytl9JZUszPoF5q/RUtsZeLC2UaQSC+rvXV9MAv9uDpxn5kFQCd0osV7icud
0yrGaZ86H4Vx0rG1O2tf5lW/DR1WMS2kcTCsIGMZ+acJYlcWO8KYZdk0f1oTS22S
yJ0V33Pk5TpOpE5umTHH+0t5Gysn6V9EiJfE9QvVVo/jcglfVmiY5Ilb7Tjte2B9
tzl9LMt37TMVBb4+fovYC548CBIMBUr9G/+r8HdcByYxKgl5SMWjvTP8Os3YRFqq
23CWwS11YxfHpg0Wekh4FelHiUozAfWi+CoBJw8Pmz9n/XZd2mnN5sdENkLaI24J
RBS1cVWbsOoj9me+kKzC57RB3njtfHLLYFWckHh0HkkLpavIgaZpjXm+s2oXlHmi
h+qAipC386lJ5m/K9R8YT+4qmAZfFYt21fQsy9eXc4ynLNQgufqPm0muzF0Y1+9g
rsydEvdtQB1CAOmfYIGyjiQVgeSGmOLTIZaNTZyE5g0P04YoPZXh95Bo0rMjiKU9
6J2/OObDqJk08rzt0A6f3TB9RAlvy5CTHkW4N/QlteGJoTczUOcG82ckqsKvpIzG
QopskuLS9ipfgVXfWbySlGBXy8/h+8bF+18I9RxCHoyASyMxLvYJ35n1n/O6eMR/
rAoNuR+rxtgSYha6U5zJmHTaPLTJvFAJE8f33HguzCWjHbTJkr8aKMlGSD4Fte8t
Wvva4YaL1WgFSZNBTGTd+VQvPBofGFtosrN4mhNBLs6p4YWM+7UbGpJHwWlPSDlN
DM8IkkuCGOVXVAhqhucSPoU/97og+baKU30S+kvyUYgcP1q1rqptA185466Txbsr
wVBZAJw13vHRpadlMOdEU6Hm4Q4xa0Mv/3/abzZoJudE51YYnHJU7wqyh9hmpRCE
KIH9BQtS5zn1w1sYX0HlCAkNO/Vf5m5OYqnOY/QnjMJHdTojOVJysviyMlb4noC3
GdreYrm4FJjXwMRG9i6UbemFPQjOshjC3ld5RW8QsFGhUfjBSANMW7WgQQJKaUGG
we7XlkLg5VClgG8y6ZUFE6MJp0pIXXsEz6fNQ42Kpx4YOngNusX9hTnzEOJ5is5G
210a6RxJUVrk81cJku7FRC+kEQ035VdxwAVybUhQ8ORKZ9GC8OryCjJrZPt+Hchy
3MTYDe8JHJvFJ/PrTykv9pw2Jukdvqvp3XveTx8xRQKllGNsuFHvUOIkSSCVb7jw
qOKZEaZR9JwiCFOx/1ls5MsRrADE5/GqUaaemzF3wM5u0ejsh3yPW9SWiS0IH1i4
GT5FGbz0fcSOFuZyTkB1rOVP0NUhOumXho92zhrJs/J66/NR7a/ef+7bWIJbTXOf
2qOZiLmdBAgicOD5Ml/SNSqH++riGnPWKMQ57VWTBnx/jHvqsTzN+CCStluewOKZ
YQDPX7cZiWCbVJ8S/7W8VuN1jAKH/0gKEM3cqy3GEo0g8KVDChmUNS1A+X1OQlNn
7OLV/l09Do+rjPtw3sPtE+Th5KDHFnfZqtB2ooXNsfqyrHpiebrFGRlEZf4xJxXp
qh73PSWPLTbdT7mZ2ACu5BRJooWlORJGvJsbqqDiotdVBgPq15xzbb6fZKeZENB9
q9pYBiVnrvtD8FC2D2gDL41EPH23L/CJNajCvkxNVS/F1+urx6DIom1GrMutl7Bh
SLT2r0XJYPSP0GsbXJQMMRxQX7E/6ZX4PrHRmyqJKsYa3PTEgSz1hrNQmLrNfJpM
xjN6za21qFQTdNZi8p9SmHf9A379FIrpGsLEi0sPL7PK7XV6XYi+mptajgjFvRX7
tqk7pjYFQq5QrUICkMo7mLoov+AnmBFmZzzmqqlfq2BEor8dxOwPV/QT+WpMRQAa
+5hEFadZ0mTyAVacgTMk8IDK8/c83a+tMXx9FlLjyH/DDWOueqaBajiqtz7JWOMO
oR/thVejwVmwnZ/FGao5bunVjt+yAvXiqq8XAvXAW3/AapGxx0ot8bxdAxcGP2di
nguPXypzQIbfx6CcGp2V3gfOvoqIWZvsMRDwnRHXxbVtWPUC4AxdWYzPE81qg/1R
F9B0WqAWQWS8IYVdMiGLqRdt+Ly3Jn7jdzJQwsa7bNloC06z9P1Xppyq2cnerc/C
M0gB3sAUIdprlJXp3SkV5kkM2hmWMsGquJdHnTtdPW5fkBPvNCoJVd1l5Adr5mo4
rgoGiLB6iUBc/lepeE/sxv+npK+8nK5tnJTvyL0tg2PNT1uUbKsWZTdko7LrXRh9
GTreHKYnDWRstLD35ZfF+L8pN1XanuodbO1hn0ly2Ev6LULXQZJHIbhDf6muR7/s
H/JU8TRGKQgkI/gycvs71xmDErw//A9vSoN0YdrHKiIRLCa8o/T8/3hhglxZteDi
IsIPWDRVVBKwdk8mcFQFtgpEVJx/mZsQrsBO6ANmEYxZEQ3YIsX+DyaA4EmzoKer
1asp5dYlAuwIVXpcA/CakItdvEp0kezSUXjOYFyQ/wh04TArQI+wz4XUoKAMo2et
PHar/vdMQNXL4QXjtC1cYngxols63ejG6tnGxYqm3qgnyQhAPn6M6biIzCwXIoiZ
BrQh6DbQ02BgeGz/w8ovb3PjXatmpLm5ljSmpBBtGfnUVzTuw5VupOa7fJUJZq68
fzShrnD2PIdhUSZ7k1vnrtFCs6G6GHJYn5hW7ya6V8Ci9y+4XYM+J25/OEhpYnkF
u9Ye+kVrqaJPsti+rbZpgN6JLncj4Ur1kVnrnukgaLCaZ3rjPqMVWfwdu7dQyJXk
gJPggexP++3jEwmyoFNGqWlwDkevYwA05+xvWMLzByWpyVlou8jzyu+aBMYmuEV9
TqxQuLEMwZ04vWV7EOQwwt6ohJUPJRV0ACeOdyodBz5MTrgPbR4iEtxO45cjcehc
Db+ieKplBl8JXYoawOqTvahqZgS0LLpMRKs0UFAibk6YyEghhup7eztKc7maNHpx
+ouE6JgVU/FAYN5PHu1dZgsHmv00LHg+APBP9d4kv1u5d7t8yNfqTBe3xLr35f5f
xNoayGMFgfmReXm1AmtwtfDwac49/7XrYD256bQRyWO9htGaSYQsiR2fPaGsDqfi
zS7Hnk3voi7VDIwsjBkIVgO+wrJipDogse2+vzsfWB+QXeD33WJCf5oxvJ8htKfy
yNiOwf3cCJlfPnQPW3fnV7bOR6PGJ2VcVh/PetMzR57FqYBwOWKP4oMwSFgGoSma
x5sexSebz4gXzxRZ5RV5Si6UO6o4rVS1Al/1/Ph7c7mmI3VwLM6FRQtMdbc9nUzV
FyMuKKE1BV/NKemfrrrl1QmqwqCAAqQbJuA1JIqdTsOrmHRUD786+E/KAlJsSTKX
49ryDJgw32uRVZh9kB64dUU1gXYMCcOCXV4fWx9uCtg0h2TmCegjoXRWHAh9m3Rh
CWZrtIjx08GYUB1yqNbmn3DurpJzQp08SPbHCw44Tf6gXh9e7FQvdoCs12h9PbfA
1VGmItCWVVEqTcGMgjxaWi5rO0Y0V4Tl6RiS+FmIXcU9EqxJkIZvJEy00XeQpZ1U
0eaGjHeGOAY5yYIOBfsklxyXqoMMuehFQ9/IxUjE0YGYEwtiCJD8QoDZ3T4rCufy
CXb12zVADszpghnHipAiblk76Qv6wRdPeHU1mB4vxBObnjQ3smHjBwGqlOJ5SDah
VdgIoadqiq4UT40v02PZOOk71iNCr4lgBA5eZUzyTALLbgFPbyJSZp+Qfg4DdZiG
MeHA9X5g7SoRgrH+vFFUK6IKRTVok5RwwPbsIKUoP4aQmyv6utv+Ln+HUuE7ORtw
7aknjN7ehvi3XPXDb4NHQ8MbKVqhW1BgW3j4A3/tndXWq0Z2SrIRnZu9YxRsytGP
31PDOno3lUPGjhJbuazRR2PRXXDkLgwusdTqjQko5g51mg363Ybmjhbmf9oYCW8D
Tu2kntFwIEyFrM3+tOKGuaU6rVetgNpU2HCiCLh4kbjzsAFFKijtEXsuJvmHSe5h
hdw3ZUrlA4+6h3TLo4yGvdZVX6HxAEPOJ7xequ4PGbUJUNtM9HvuIcvXvdZa4+kH
BlcK+8tCnenwR3G6yhrE5+Buhu105jpZ7tSjPeODmBD2aVvXCt+OIQxlqwb5KF6P
7N6/ieiQI0SpGxesC6S38jf+xDxJVtwgX9qJ0iBuMDr+mmGtYw84TZnjVsWl5s39
Ay10XsFvlv6lbQYvzwPz1HVZOgRKvwzP6zzCB+rMpCK+w9+DmoqXQ4JDVRxUGzH2
DEHfSlmVy4sUblxOxE/3F0hpmrO4/c0l+gJyzetaQgJ/3d7rzWBSPWJe4KhzsHdG
nXEIpE3OL8Y4jwQ+0YSv9kQ/NlokovWL4fwgB9sCIflSZewen5gekAOxubyWcqQB
Mx8wY7VZpowWa97dFRGTBNFaW3K02Fw0pyj+uxY/Phu9Keavx8z/JLe3LijZ+FF2
j7DrQKUX/FARnYNchoaEJG2a3e+wX09d9TWAMbqdCtWgb1DafDtjzXJyV8dqATuR
vLGFuXficb2LWFjStQLX3gqY/sSW1QNJO5ciiRnRW/PIIRt8gnfbnH1wjg9kpT0e
LfignzEjEgJQcceAApcir/rpnDQJW1TvhAVYFfrNk6lubqA3SOEwNrjI7/8AAnwa
4cfAUXUGqP+d1zfXDrP6rnO/WwxuoNZXGFPEU51CY/uxEhsC46lVuMdbMO4/Jp/b
YBZQ404yiiR0ubrCU4813M6QiCXA+qrE84oQjiZYN1KwJ/ovbAL2712iMWJLJW3B
UTeeM1oKlf+5m5DIYlu61x8cH0cyg4gmXLNX53qLhGdgu1+eAPikd2d//d0Vmypa
xmprLVcsSp1YkupW98aEZ0vVuVemsR09B2sKWVw7RyIF+hT6RL+vOPMXgmLG80wF
YhpOxAbrdv8tgypj/TK2Etud/+jS+hmJyvksZToVpnLccLakEsy3CXevMP24O82z
Cz8lgIYCi0WGNgr/bfjAtjd7wM66B0uDwwJO+8M26VPE6uB+rxFFaZPfl2W42mCh
qSWT56v1xEf0iQ6B5Gt4YhdTfI5x8eb6Zq+2z3IziQcWpUXcfctJIypfSruR/Y6g
U4LEUvh5COoXFRSlBtQYhvqANSF6WdzO5DzN0NyxiSLaERn8ravVEkY6OEBVOzoi
SOOth7J2J+rLJHEnAXQZ5Nh6It03PJOH8e/5h8BGqCKOZhedaPBiGwtstwlqEQM2
dPC9PSLZXnQbvUnRnksqCWCaK42783JKYCKEnmsYm6Sg/J2L0bPND4XZ6gKcFQjb
yDUKd8upCQvYfGlF6mrFvpdYOFolopDkJhXicuIIoy/2OFARKdSJFdJYvgLAPuwP
xXIWxfXJ1O2FZSqMsrrxKpqz/18FiOxqyHEFh1RQrvrsaTJgnyu5rprqXH7Z1eI6
0/bOkv7XyPquotIYvg0cCTl+UqTpr0lhbMJvQqHW/mr0JWVDgwQBTj5T1Owct4Zl
MSRkLyC6cicMcNl8HXS0zBBKT4Omhx0nWKnqk8CGgDtN82a9LQgOm+FEWMD7qmbx
h1CvsJViotepUUUtR+T1A2vSqZKFuTJUGXoWFwcitPFXKGAuU0RAjgkotouxqKjV
L1kDlitflIgqbkhEf6sDQY9ORDQMRYXd5XuuYDy8+IpdD0/3ZnZwkSujTCOvQspl
+u6MYK8qZmC4aB477QcPGRQn/QU7qfB6geQsKFptNBcDYtey9J22DFax65B9H5PU
kQ8Amqi8iUUFZegUgBRAqftwBKOyJvoHJfYiX6/SA5AYYs0+cd5NKCBYZqRoXhDP
yo3JD4wTFd43VCUX22S53+ZGNPuInBKKd1qDVWH+HiS1Kqf+IXzKsbdKV3hwi3xg
dyAu63DfLphobzHhPHfamUaWQj2hmiUB05WE51GVTIcXtRInzTi+bJPtVrfLtHV9
RDpeD841umob1HgbsXwGrn3lTQ5FznbLUCYXTEtMVjLk1+7z71lbtI28Y89M/BUN
uPb7KbRdmaAvCtzaJ1FjPlOCXhNr2rOw5C95xx0yHXcuoHFTHtL2oWltqohjsw+N
NVq19kugkhI/ZIBtaQuYVGfMNG5yyAbI382yVE3q4Lmo5vFdy4tqyu3VuI7PEm8y
WpYvXJrfU7iChV3Jg4D9IccgwNA8d0R6EwL++97EltTos5dj+w6hkeR5ThuYed/U
KyPQtNg3dzi+Kj/LhkUbo0o1jXnzYgwtMI9EGFftdCYlWu0hqXcbOnAnAM8AVOT/
1x5kJ5qeWNY5vYlqCRSogPc5Dt7e2BOvorZI52pnHqi04evmmh85TNoxwOXe/b3k
SNqdGrYbJVl/gbNgpWw0lUviiFI+qwSiJEjxoViA/ytII2xNV9X9cs4MxJ+FUM8Z
MXqPZUqeZw2rYreWzDhcxGiRMpTkUyUqagSlSF/BjyWiQOjfEvTnNp39QeJll6mF
PvdVlNxCndT0kXJQvh0krC0TvXp5h8IZmiT9+5x6Xxwsb1lUN4nxZLePcE5k63er
JzC6uD5fw+Y8zTkc30u+d5TwL1FX7bqs0aQ6OeEq6+tJ65O1tj3kwfrAu0bB/T+t
kzP5QM8dF4HqwI8tBZ6gFB54fX23eLgfiyY4oIIJhoqA85cGCHmH1J8nsOoJAZTv
I2My5MJcXKeK9B7BGeTksbWljJ5I2JOchJaxc3XzMJPwtcuU7FzWIQeCGIlXItQF
iKiCbdG5rZnzbgonVA+7c1ie8iwGp29/RMwMDRDzdY9aVPUh7z91oPkKIGp1S9NI
DFoiLrzf1isY6iK55v+QDWwWgs14rvrtKysXJxq9hAZukzsNn9hp2WplDt/XBpVc
Ig+ED3HSlH1e8HEzwKR3jzEatyHM+tswhtndSIXVXvBroZFjU/czkk92PfDCQ319
oktZ4YI94S2Jg6DujWdj2S9HIKWqDJ3N0MUONm3T2k61wKOCSEPy0Zgym2JATsdz
etn5pEmfoFdHx/hla0aAoUGMg2tFOo0IT3c+3kAK82kKRzfICDnZCclUXzjNaqAR
M0d7XGLZod0TFQxpSjJMNLLqeToqlruTfNnkDbHmhIPcXNi/5XPpPuAtvVrIvbBa
wt9W3p5k33ObkgWGag02Sj3sJn3YMmmmKMEEWHvdinExaH6K4xaONj/yrZO9AC6g
6SQMa/nv0cHIHPwsjF9riMAphwXL0uPH7aJrTN6qEnQBo5b+F/FT5ABU+SjTjeTL
vODljrMKJI6G+d7L+GDcJwpZ/XgoMVGTSOsCM+76731jzWMUQvPiJmYcVPtVdgaQ
Lom4/6Hj4NAm8S95v1mo7MAV+VK/qBq56fW9v6Tdny/lu2X1VzW95gCZOwgY6AnC
aHmVJzCUpFfDTamZHxNO4Fa+p/DaIPPlHs1/QdwdgkFGBz6gpIz0GMQyVwwd8VQo
q+68XJ1GJQWH/wGSShoczXorF7tvOegEmQudvFxgr45PrHxAKqY0X0QzroLe4V5f
BlJBc2NQKCjqBddXpWtdLoUNFA1g3oYlqnGW5o3ZJ6XSfHMB8PhRuYAoxuoInTcJ
ioPnjLXnpDeow9Xal6nVgGVEIwFOVnq6lmLwhSOFMCyDW34wiuR0DHsK1LJzTaED
EB0Bxt8TAWdj6uT2rj/kW7EAK5DvP3+M0Z39fXl4I5WeEWjL1uNTsYkzX3njnwzL
t8tw7nfsYnsKiQmu8OJIQOBAJtSOenhnei0P+INJGRZx1SEhP1qbOYA4YUD1tL/y
po1h23lIlqgzWxsrC4sxshregbp2i91WAvB1+l2OzAJ1Hz+mLzzJoDPT9fL2Cxae
PnW+GCHDpbeyVl02F8rcQmIo9td+4rzgTZLiWEyL9B5O4o6vE8dhOOgufppXBBq9
S06OOn27gFJF/PVpfADTj+9z0uleYYBda5Iq6ImDYlqofuaTIWAqfengEMgUP44B
twcSTPYLjv+neqpLNk+Mrtl/5Q5kjyiaSVBJuCuVzTtm7nhxSUsKYYhM9Ao8Sjgz
btfG9zBoeebZZthOy5Hd5UxmMjpMvWrLC71N2sQ25DIxjpQCwcuMTsmmuuyBlexS
3V+CY0RA+IjCQZwDIi9qljppGHL7eCGUDo/BdeHuQr4efax/JiHKsBOOVAlCoUTE
Vwlg4jPA2l+Nrd7WSIfspIig/iQxXdSQBJzOelCZP8dCAMYDy8LpCGRZ0vnma3Ji
U7k4SVUKO8uUK8IBU2FJ7fjRBvJyE9SwtnTDOw701bTtGGLDVsDH3tDUSpISpo59
wVHEbXpfsY3OXmsE7o1Tjkk4rn+FtyVsQJ6pHFAJkojFqBpMiNIswca2JOM5dBqo
sdZ+uCI6no8JlZh13iC9eKpTnJRwUDTO7HBMd5bAHX+74CHd7orN1T7lKgy/C7DN
rb2CDYDjWZiYsOjXvPQF0VMgai/nv+J+JHJ1XmEnU/2bcy6SJG9E1HvchcbPIXX7
9uPyt7H81y4N+qlm6xYGnyQr/9FINFkjZExaB3YCm5RwXvSl4Hxohpa2mILsksdz
tLsQVKk/jeLASr0JlxFDZcepkjvW2FvtO03Tfq/f54kJwEzux1nhTNhOLHVoVY57
BN+46J7741WINQeiXdK49u1I9j2R1efjLJN7kFW+AbKSGLrMe8vRKkQ30PJLR94c
w3OvRH1Qm3JuyMiGrIlxYaMpz7/PZ9ZoGK3pIFiTu9rb61jH9zX8WFNW0uPGwqnS
y3lHeixWTtDr7Se7qgZwajY/YGjJr1Q7K8A+zFFLZPL5h9X7q2t9tZX1CHCc4k9V
VVLAO6/oGoZLDKmWU3CWeOfY/8CB3Ep1FuXHP4eOc9qNqjlstglnymn53mkv07eB
z0kAPUsrQPsmXgw8RZrtzGA4tVttUIGV0EWB5PxwoAztcuvq8xKpD3jYNUxfl2zW
yAT+xWASmX6UBG4zsLNzNVYcXW8RYQnyTNnNSy2SYWzACGZWyXXZSXeqJCXVr/dB
FRpnn2FYWvng2AmTmkvxuozY9EuD17NXS1s8RfeJ6A6keTzmVHBKBEFwkGfEspbM
gP3EvUcgh7PQ6dtb2PVMhzpBAVLabJF8+qfYlsrZ67cJ86R10XZdCi5aZfo8C/aI
Kamtn6oHvLTK63ZgaOPlDJtMhiqdsLDWzzJYI+5GcO//MKNFfG64QTX34SmMF/jj
uOMI+DhibHEddQTZPHVshAlq0f6VOq0gjeRYOJiwxa0w80+EjD3mzluX+cja7JWr
tfzMlWi78LfmanJoIjgFKYfQjWDfi/OK5rgvN4Ta41Kj7XB50f4yflXJbzZvp1qv
1oI999066S06SBMTIFB/ZAdKtsGO38ePSNjfsp+NKLaqvgmYgv5oNqZD8BQ+OSwe
kLLZeut/H/EF1JG8wN3wP1HR6/+Qx1Dfbboyw/IdxYecT9/vgJZG6U7Gu2e/ThIK
Yc96iK8ydmbiMUrh8PKGmzNB5SYvAIon+U+P6sWFUStzwOOgD9CA7kIgMVQoxro7
EEZMgpeiCy4N1ZGREhTgjRRTUhhEjHgvtGtfKjMredlUZ8NQVPjYoGxw7OA99Vjj
NdezEy9tfWbuNxAQDO7fTwrB3P4p/xjbSzEAd5Pq29XoZbj/Z9kRsOCriKQWtV8u
mocSVHr8allDuv4Fo5Z9NLU6NYx6k3kpjws2IBK8KQDq0cRV62a+TvHu4eoUNRQh
0fuLf46Aurq904lwERRXW9QRdwUpzB6Gwttga+bSRQVr/1v4Ih7B3TnnqNhfjMzW
NQcUF1ia2zNxtQj25Akq5Lb2Z7TopFhQQHHROM4MFlnGnuw2gxmKuhK+iMeEDOm0
wolo0J2ZZ85VLmyoDLu+YPcduDTzxeHCed4sA+RQqpOvg1io9aaIJxfJaYLbMEdr
S2cf9Sc00QroVHogPuXVX11SkZrhKU+Y6228NlVczqx3qA9t1LwdDnhkGmUoZ7ac
3Z7llUDkqKBlFW85rVsA/SF1uwNQJFqOBIXt0u+GiV440vD+1UEJnu5mqLkUTgmx
AEOoaq9+mUkWG5C93Ir6AQL57BgrebvZRhf+n7QDPmPpTiORP+sLEibUzd7opakm
v5fYy8pP1S58Zf4tgmLxlWWN7pozYlQ00aswdefxyKnpxfNCVc0V1CQesvRSqKSe
c/wnitk3HuL9MnPeeSPhnersfWA4X47lf2b+vKMiPEjLdaDy5iswT8HD+BLsg+nl
uZyI6rp+pa8SBS3twzz4N60HpsSi0GftolWA6+yFttegzT1ex9JaIakP9wx5h3XS
l3xBJKAS2TKij0MvaQx5f8kHaPWkjM2f/Z9zYbrHzxSxQ0K1+VGOeLWz2RuF6HRU
Kb0fPu3qifBEf6ZXShISppy76x23tknHp39Ztm1IfR9PPP/M6aZ52tQD/AIHa8cY
Y+R5Tij2/vgujbEH0EgivzcsHrIldE2kUp20pyQs+lt4KDl9y9lTAb0Fc4vgh7JY
Gv0krpM10M62GRkHPBZhwp77QtcupdF30VuPV4/l/P/DlE57YdC95RelZppw7cgf
lDBzn/VcoTl8nA8T/ZSatqqWR/fQCk1S273RGsmnhjhj3bM7+S0IZlzwEmTn+usu
nHxDl/dNKzt2h30lxkZGzZc8f/I7mQ6D7zsJFUK0nYfjfmRsbBktlOe3UJwtKK4D
0SqA9zq0W4u39+pJosifnpror+ZhVQSZ4Q+UA1OgnUxWoFTM3nPx7Wz+A2dttAcJ
Tdpg++m7nqkC4kB5gMQJjeq9OywBldiI/I1eq7f/NBjOuGVMmNPMQnuBfsmLexzw
+8ntqmGLuENYBd3gipn5sZJPo/o/FLAVbJGCUyLeabJFsHsk+325NfzTKFbA7lLz
sygCLOWES20ivLnmosay5K6CmX5LyXriEF55XDNycHyEI7vb9xf+HwAYLiUWRU1m
ZGqqN1mJE4F9jEFYJ8proqbpWLDl5Y01NbZnkOdOUKgPA8hhGG4Fc3YPdeCCDwFn
PGedrvgh3HzTEZvbPIAMKM2FTAS6DgNvleVTR3Wp0kC46rUC5ytZAe7DRIG1hShP
hoXVqe+kmXctYuZresIaHFLpBeXk5HBqOCqCl9Wj8sTqOBwjKlyBghKrkPuX21dK
tEsaX7WTszKb5KLDKx/HCNwrzCnDgSh0ZCxenn/DKF0+QSkKbLdbnd7Jt0R+uELh
NXg6ZgeRiDUZQzhPCCj22W3TwxRz2QH1i9AjY6xi3+Oza1x2XU3o3AWhoim6Kd8e
YKs/yB8UnL1ceH/shi3bCArNlhThjz32h5NCrKmJL4WU7pIb4Fg+QCnXfP1HMNUn
DmOYWUUA+QYko+cjTeEqJJ7UMFam89Fl3XqMjfc2NxoFMYpECfIEr3+zUiWFFqy1
YU99LyKfHpLazeRKkMo03sA8irNuBMCbolHHOCNYxsB2JPewmOvadF1ohNVvw6Qx
qTsX8ONU6/D4LCb7lcZ5fVv5D3IIutdp/f56vZWSK5FdQk6+0BvgUkd4LViiMi0H
uhFAVyoRZ5nBJF1N1O2hDjTU6j5Bm0myG7wxMvF+OYY8n761cjy0RTD5SulmBCRc
hX8ICc/Q3GG/xpxt0A9AM8wm36JaRhppbyMDLWS+TZDIwgLjqBaYswZfUo+ZtQKN
U0pD2x/sJhvfWS4TRS3rq/eVfvpVCfSeeo8izpK5PJ9AwXtVaQMLleWERzSv79aE
JFqkPqJRHlrB3AmXUjqHgJKX7BncPJOPC5oipECKb0aUrAwJgMYmAKvZf4eE0cYL
1V3Y/0VwjQbFIEL6v1EH9PaWW6emgGarBX9AwqUUHfcdzK92Fl7//91mqCUtV+yF
Ws5v7SOP0zIPZT9FOgo4y0JBP0QXBTCp/SMVdnoP3amzW/iGUxmDz6siNSmfB4nX
/2rx4zYgLFZYN4d9NZ8ao78er3vvPvYsTrMLhHXBnKv/5Irt99MgTxhepN9y+Nwf
5NA5eHddyVbm5JPnKKSbz6cDsnNZX6WG+cSDMT5YQGKzD5dWkpT/TI5XhF7a6dzj
6YkZs7p549PwV21SFJT+TmyUke8XFzy6TgjxNE9i0ZXpsIMSlbw9xdtB+9gQc8hd
Uj+5XrNPMvIfZZHus5EO5RAHcvdl4BV6uQyxz+8NE7ULJ1Koy+C6H7fNZ9HwAcE8
`pragma protect end_protected              

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
MQC4+FBbvfeeB6Q4w8tEJVRv2kfxnLdq4gKH/R30Tv/BIfTbfoTQCnSY2KF+YeGO
OIe+vWkCVKT3doca5oAYU5SeN1i2LStvg0OYt1QY37W2XAOkIzVT+QNdO/Izutw7
Wvd2t99QPbjUNQxYo0y8gXSx1Z8UTOLYTe5iTeBby18=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 205540    )
lWmwi8dp2UTePRvABmpoj1Zsgd1O1goW7p+DJ6BDRkPO5dvIGZasn14VYaDxrqAi
Xsiipr5lrhnmlv16UiirA97BXOf288Re0spTii3aiY4C0bjL9ggkgNq2gudwBOIs
rzKBdpsXeX6FsLzh6JIcShgoF0fq957fhn9NwuDU+q5nvJZzNrNAaJdGYF1sItz8
UbFnhzw1t+kuqW3jfEq0fnRsvlk9955IgT9wO8r41rMxLwIN1eGeO2rNIzrcAg+j
x36pI8k9nfIhLMqcC+AtGpq0U6KlGKBjVPmBmUABXm0UPBL8v2e4kAZr02ZDQtXK
JhS/09gta5eqE/WASf8sKlwI0jsiKvRklC2sDr7jQl3pM/Rpika+N/QjheF4zgdj
fETXeVYAZq2vsyhtj48iq0bTvhYK1Eeykp0PhHL/jHHW3akTZYPpqAf+38Hw71hI
0ecniyEYCNZbxLQB2AI2tM4GYAngaEDPyzxUoo/lixh9BMTiUPEiif0qFPwQCrpo
KXtwZkRlbaHMTjdfyJ8jNZwwCrQuxHlFdmx/Pianke0sa33QUNbXPVRYtII5qPtB
lkbMCS3uoxRD9sY6V1lQ3ZqcXf9DgrMwjxEkj9S8e4mqbYvrBD2sAp9ta772wKAf
XBwCxwghKmWYcDOkS7Z9msL7UtFhvGCZ4RyiCtd517FfpYiveINIXxOxGQ4Z4pi+
XhYSah3VDTmL6Wx9TwUHo6r8IGe9SuaMY+sncLRspdnav0K1eRNkvH0Q0QrJ+XE5
nM0KQYj7X9NppSYJWceH2OWZbNGdbWlFOL15AFYpClw=
`pragma protect end_protected                
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
hzGhMipjtG07lKOi0d3F/2IsJRYxO/I9NIYWrVjPVV8Tqzv/nL2JVkfeFTjhDyYL
/6mA4+vEglueen4ebbhoRSW498K0YW2NT7txZQwa2bQSYwltyNRxOM68mHFBM8XY
YStcLct1BWJF/d6c7ffg2JfHKBwX/d0JV7EDWyF66CM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 218658    )
jwiToeZgAbYWOlg/I8/0AFM2mzlmMlnC5Unox60ivd1k3XxyxdSLDJ3g3u3uxOoF
NPwsRGrucLvN7vEq7con+8A/LfWu7JVeWyDK9Ma/H9q2bEtaTqSJW7Bpbhf4zQZ/
Ve28cpxyw1Mm/TWlz8ncOsa37v5W7U1AwWolA+lZpmfVOoOob9QwcCDVxEpbkvFB
MpXCK82Jrxo72LNQDHOvch4rThj6ABmUu9JJEp+I6OSqmyu7H4axPM8BBzAg0Ou9
Tu/MB/ac0uJ9NUxll6HqI65IoKuoTZcyWdYjNZo7ZtWII7Xlq8DRev4g9eoPuNvR
Q79H7EuTC+WUeYalLJ/MX+KcS/Kb5Sn4Mai1QODiGR/7n5adoa4K5syToE4dViBZ
dWok1wrfBhkmUE8HCc912eHDcFo/gBlG7/WsviJe/t+jF7DXAoX+Wh7g2fLNPHU3
MemnZsyct5EzBHGUIInwJKjjWuz/Q+XOQHhmD8c9xCSKAtXog6gr4zgtqyAUJsza
4BVNzlT8IpAnoTXO+h+GugYDSM+YNnxjtZgoFLSTc7MJzBpVxaasgaG62WoNZfhc
QaGQQMnuSNH8/iPYv7jpf7QNQ/ioyfDtzx6IeGyMDTrMKPXo1+2KI17edXBZwDQx
uGZacLxokDcXNZjLzYfG4xGTseR2ya9hgWRsW6gtQPQUoQvTU0P8b//2U7vsgstN
DP1ql1i9oeot0H4L4cwHE6KZWRME4GzhEQCIoMyy2413zValmz2KzFSgOE85+7SX
ylN5J5TMlgPOwKsyRHfZdNd8Rjg6nLR9g+FCTOLRjFSg8AK5JRGzDW6behG2MiPF
KL05JhRHMDyia6JCaP7RXNdNkbrHApjzJt4suCIsapulkVodGfh3ImXoCOXnHSDd
PS8WB46hGpPPAlhEw4JKAuzLT7yIgzJGeKsuZ4gUZKTeNu0qorVBQVbb2lVrs9tN
/5mGVkGIC8dfga5WMcQyEbYNf/RiTVzlilb5X1oJBCp4j6aIP7OUbRDtCpLIiIZg
+Tm1rWNoURjQZXUIisVW57tHDQFoxtm2UMr/rMGgQDd8HGMKbDtdOpMZshYrqrGF
5sZJJL3C7JY198CfxPppg4t0sj6BQiMP3MXvqXXLzmp6b3mTj77QOuRud/4hgBBN
ZoCydqtxNq5ylTTBCXbFe91vrKQuru4iQLOAdVyqwSevicEe6+6fbiEdfNEoxCqY
p4EOTXntAueqzZXtw/YR/PTBauLUtEjCw0wTUzod704Pz482G/Ni89nnKPXfNHl0
eK7W3Jhw9exH6UueO2zEIZU1pHJAEhxetSUYDFSCF3oPLfYqIhqltGVCbT5NvRYr
s603utCzecTn7W9/4ehOQZb3IckpkPgIwyUeDzeZ8YHU43IxChsfDNt3kX6MElAb
B5pmHYKsKMyWJf0CT70rJY5HZxpj8bDFueGgws2DSyiTqF3olaui9JkYBcSlFEMG
xokFfzgkKZtBVXodONc2EgTLBcvdkZPeFk9jxEu2zcjfNlNTYydxkTjiYOrNrw37
T6dORJekgsEb2ZYCGdXTLErzTtok00zR7wIlkXCtKd8vBo07fbzAPVIHojTLIfiK
K0o7Se0yGd6zDTCE+UotSLyQjjhO+0AMnXj7yizCTP1F4/WF7GWTvP2YCwVqsAHV
dMIpGqq8XxXurljNescYL/DSBd+mjBjT+5Ka7r1TGlmKbTf9stgrBzORKlYxw9xC
0KYzFvB7fzflBsLMMWpHfZs96IRPZ5pE+YDuqph7pXYLQjpHefqbfLLeNMUfubRB
LsP5Zu0bry4ZgtciAmkYyJFmS0vA83CRPE0pYFPfV1kfj8FHQiOyyAYiEXZVXA7G
d4b2du9N6/zEnMmZjD1zExmBmNPXrss5tRza5s9CsdiAHZ92yVdNnuyCOeDx7Dl6
FKvwMUIIYID4BRRfC29+Okr+8vlNnsi2uIjC5llfQH7LCjEFYV5Luec/XiRXbvhC
389nYbcUPnXy3G1JX/DM0ype7YI9GB64I9D0Z389KqhCterCkXJeR6L674fejGkc
wQRnGv+04QN3ZszgJn5SBJZkVqdQmqBkJCkBkLRYEd52yOtsGsowKsNFz+mYtI4k
6ls16JfOJcs7OTeWkTrq4e8gWViV5mMLFxbxR8XFb7kzvzVPxwVpehtzT70b4wfS
2oVc2v/trdGLAh/Clh2hQfT6pplqEgz6A4tsjuEp4H4/sn+nd79Xtphn2TChpxfF
UCYWuwphQp1q+YuIFZEFWw3pCbYVA2ZYNAv5nF5/miZR50WPSRNlxMiI4viVCJp0
A7m7/a/NB4M1aiqDTeI2FrDU8VcG1Se2PZ+VXBkbxXKR59gmIzaxvNDnCX39EDiK
U1UFJBY7K5YGCeQYzocoD24zq/b3aaKMUxW/kCenvU1D2WW+44YRSU8gq4N8FDmi
4gk+LBYclOFQnO8ZXxPtEQd+QSgypuw/+Iyrd5lwadj2jFKKUVxTh535XtyCaUIU
WapjopyUzmrXQ4Irajd7TZP1AVDVThI5MWtf0qBYLHt61ujjo2uGi416/EHJKsXY
xrMdoTYswl8It25LoTLEgu5Ccb+EV+7NTN0rH0q3DsiNHt6Jys39SGaYC8N8/zHG
I2+qRsOefYKKOm5SUUe54bY08rmjUslysoZE0CK8fzMxV/DaFHTZgHeVkj9Es67v
eZZfWUl3qaKtvNQp6bDMHg1eW/S+lpGAcAsOr+b4nfkxA9soZw5U1C1yUlI0DVuv
AZiNeP//FsN9LRutMH/WqjB6/00BONL/B5YgtQEskk1JoENIOB72uOlt0yVduUDZ
GGu+KcwdBNT9QpcuErFeFjeMZYRiPcuT37jES3H89NlTGoIiTRUeAlyEoI5Pzut9
GxBDv4P3xO39yf3xSGWHYkEj6LtsNpvZIXCIQB2hexYLcFr8Hvw96ZEv+VhEdVEs
xJadASWPhkCi0sq3xRcHNiG8z9+1ecxAw8LeRDyDBIpOGqr5enhn/DQ2yKKPOxJm
kx1u6O5LNK0r6hgjNuYQrDX6NOyjsm2XZS4j7Q+XfsWQL5p47jBGdr1XQjZp6WAI
z+LIGZX61fpxiUDqG43Sxh99+Fr8e97KPF58t7I/E+zqIYauzMrIKVYuR2UO2vFs
SgdmXcqHaAh2hpSUYua3hKqIFXwktVFKdDN8tc6CiOidcAM/CR7LIwu2UdgnMReP
LKAKODLsn0XFtThdyjIUP6f8S79PHommGQRYwogEqisWZQkKCLGKbBVWMNogmL4i
zgj1jxLYNG/VekFUYDfiEsIJNQxFj9iZze6jQUJot4f76aShGbopztFPtTAsG3Ro
Eklerq3YmYacUmgQMwW1CChJgi7ng7rHw10ZCVk1Yj2bhcT79QmicPCEmv4VNLhe
L8Af38EoKh/lhoTwCPLt7YSXffXyTQa8oinnW+WgZAdVHWR/ZCujQc9OLK2L7cwH
h9aM47aTW4DcpQHgsmZDpI3Z0grkhxKXvIvtWvaqNR3SxOa+5rEA9Y/xzfVQkVW0
gQyQ/v/j6qrG0n8lPdOwZV6JRG9u3Krz5BKs3RAhw2yURY02aJA2+8INvYHdzuDa
WfRiFQ5itqnaW99EEYC50korxQeiEGMKmuNU0c4AQRk5MJl8IvOPdWMYSCspC5Gi
JSwq9KRkc0LmX5+bpAl+B2DfOaXtWbqocatn7PvG3McPWd3yMNnnwHIYGAwZMKOC
EyNn0w7HG1FipR5NBM6zlA5Pj3CJXiBx4bDLSEotAOMEoBSMARD76VGEs9QkNvi+
ixTt15qKFrDluBGIP1tL+4TU1vaVKFQEpyeYpDGzPP95FqrJ28ue9IpJ60x2tyAn
IexRBuqAyycZor+RAx5la93VW4rSgZiOi3l9Uxy8Kw9u18RfURKNVaz3X2JYSI5y
DRoKX8BaoxsfbmnOmxDSWxh27/kzlTJ3dfE4ZSNEtg2x80xVBKQv1iDrsbfEfMKM
p/6Qq/o6xVUjXn+cD+M2kUlgB1qq4KtKLk/16ui44RmWqtl/e4QaDnjdw6FoIp5o
KfOAA2WXITAuxMVdSYsNaWIahLydV5ZoVrzIIxA4vZmcwXN+ge/8jT8XYSI7SPml
DDd2dXXbqSdvKcr9h1LKsZ0gWZ016MF17ArCqb/DkYhlABGULGIaEjjMhIhDXadV
upSXvR3MLw9zmmzkzmjDuZnAhbLU0Y+zP0Zc7YYJEld08c9nAbrDfDsPOlhHdnZ2
WHUg6uB2YdIjm000m81LnhBH40z1uaIjJ0a2rmQgWZ5NOmUT3pqJC3PR1LN4Odd3
bbMv0nivy46yi78wkcfMoNLDQqjdMNphrPvjw0NcnOgm2iZ3vB50nuULgMG/n3bB
2itvX+zcktWJMByQPMZCqBKjVTPB9TW5OkZmX3GLbFD2de9Ex8WuU2vT/Gi8i0rr
Jit6Ts07XY29QyVMQKUoVAGx/3YIHgkdjtow7Y13xVIWulfyY7S0OFd+b8+BAMDG
HJKziCnzJA4oQ/2tkcCTWG2Jl8dYMk+aGs8rmo+gTR/XoWPDEBonZpg4C45/VwNg
JiGBNZPFbX5wvGZ9okckOflL1m+F+Ib2BrWQ3gatKW8iio+FSryT5DsrpoASHFna
hY3dp2QkgAKPOax4eQDMEKLbpCEv0lOQyFw/D1hZSjTncsqKhsIs5LtDJQvP94pI
GGGw4Rq2/tec7ZRlS5IkZx4u0qKaVhKEoQA13XewqGxB2Zr5PshoDvZ0KFKUcHfJ
ccpAw8ZsacnuAaLmdlYSzb3Klfp0krcdcZdtELQaOn3jNNeraouZmmAVzyCVpjDn
2UIF14OEpcbATfTPEVbz1mQX4dw72BVeIQx51OibpDdGrvVaEw44y/EOLHdYVajK
Phz9V7dloL4IIh2x+HfDNdJadqltyGwus5fGLG3EtINZnOK/ZHX8xmncRjtixSoG
u5ZDYztWHsBrbbchj+rASiJmk2er0hcilspglWCf5wOGaK7KJENVLw+7enrqUT3n
Re5oeyeV/OADF0/4rwzqTzN0Tiiq3Z2gclCBykjm8IdVjjUT7SC3vNpv5ee/xHVC
p054GLtmr6qMyofVYSSQhR0ndYnpXfXyl6DgXKRp0ZJx8knmcAp+w0vfU+RgZedu
MTyXdS+48bbcVZGe1uWrFLqkSW5NMreegToVlDR2QYgP7GwmOAJowkUzzbtGf06y
lNjxNKHEJTLsyVKD3IIi3D6uhcolS/WomVE59RwkWTD1n7iqOWkqZzpNtLDzvf93
DD5yaLYdk4KBPBMRzZmZWY9Bu/EzHmq/I6ewZGTRpqnz7zKAfjG2xRI7SCbdlHtE
c+z0DLdqkpABmtm0B+xFSa0rcYxVOBo6kXZFZZgKybEaMjky+7mh2ovzm2U9Egns
8TNbgweuA5iIq1np+oJHEJFk0ixyTrVoD5x/BOsjVpNxskzrfRaEsZ4gPFiSWO9A
54fSTHRgRqCwQU7l553dATOZYLA03hl3Pc0ZKOqbDe7nIogMxeQ9z0cIeFqV1rOI
EPO5i9KD6/Q8sA7DC6HUWJWUiPCZ1dE21Yi9c1vsTHzHRHspjN9jR8sEoZXO/vau
M7LDJjj+OzNfBQsaA09xVFS2ZpV/l5i9IwD4Tkbc3Vf+6kB/PCNP5Wga22tbRDn4
wwkFIfApVGUXUfhoUrYBiyoTiyys7NDKAQzVEGGeF7bbLXD8WPvxeX1AjDGW7Eqv
eXxawo/FCAbVs3cSpRqX8NIbF5nyowNL89Lj9BODI8k0S/zpnapsk5eqjqB4mlZ9
LayD1MPB9PFO7HxTNtSyCnxsGAyGjSkUY2DAiYbYRXNqUEsnqkq4FPFFPp/VptoD
euUoaFVtxHCQhpgbpGCqzWn1k/pZ8N3GIWoHfZn/CsxyvEx/wVcoMOC8yH95jwOg
GAkPTu7s5Ss+NSGu26RQ862TjPFBFP77yCIszeLBiZxP5NWmeKDCoslqUWotQsQ1
MEpzOR9tHdiXoaanXDEuDnEFMFhdz/nz++UXY5oIxzbOCCRpgs9d4NzeL2CA0tEE
R9QiOaTZzZbeFXkkboqI58VZ0GRGjIRWwxUD74veZ/5CTJr/k3jr7wtKyPL4BpZN
ikxfHF1g1ZhzLE8o15tlpPM8GGLrKZip/PfAowoO+4CR7BZrMNW9IFd9vRifJKFZ
ck+c/rXGFRvrtpMwO+Gm+8JpjAP6H6pSUqcmhu8h0SYuVzrlE221URmIrlkGGR9H
8ujoXciqqKnBQWty1SgPIvdnr4ZgDTZZz6IlLtyrCMeogICqkmCul1sfHac1VVHo
TYzWoEEuKfRSVzESwAn6OghAukfQwFtQ9OpvAWcuOtNe+4ExFkz9HuMI8HIK1FgG
bFtWirlBUmjqJsWP3qa1WP7Ory2I+bZ5i00X8n0OAE8ZK0NQ/pVgf5XaXq4geR9I
Azwlh89Ko+sz3zDuxy6QlB/FuqVQ4ssPk9FSN05sygfTH54+RETVv3ojoWr8f5LI
oz5h0ASLfRaSXqFAgeUVR0YE2kPXf5XS/DC68Nk0nV9yKicoq5ph0OuMw86w0yat
SBic4H679CngPft1hP+K5NKDXnbcSWkT9fxMaoOJIG0FUxZ3JNX/jzE2mYcvXwSY
Ow8RZzZvh5MS2ApBS3N/fUwkTNoaxOqh6rhBtxX42bMHt+epR8Og3f0qZguxkm3H
Ws6XMwhHq6ut8F/vL27z0jz7XjYjQQ+C1nrcQFUm0t3HxnA9l4A8sJoBU85TgI0o
+hFSMWBNH6CXrkK6d1VR44KLZ7eWDUxSG5fVALgrSsEZ6KBLghBqoGFzohY7CWIS
px7uGOPv808LelUWwUT6kqM/+p7oM4B48i8QIYhZr6kvDxGqF1iLSCzibWcgeU0v
ti8WvV1UmmWw/tuWP//AL+FUgMgAbe/jx49rcvOHosLpGNiPXPP1a+THqArFeK7C
TPuLyEKqgb0UJPtfnqaisU+epWA9sWE2YV96bzPT0xO+U4bHtaSiS6s1hw3h69ox
Liu1jE5EHN1eeXUDKe1v5+yfgwV60zMWvF6Roy1SGPbDtDFwS5R9zoegyb4IMwbs
CkU572nSF3Yrg3SGd8VzFYhJjZxhPxMrWw7norYowfalA3IrOtppOseM7fAqRwOJ
T6TANew8bQyRzhT6DBtPJx/k2xJ9YXVe7Z2griNhVCuN+lX4qmqrkX7N3fKozbfU
cEo5ZOD7SCx7u7C9I5OtzREdHM172/sk3JUnjr9MrB8zGaojmxg/e3gkhaTFf2jg
/XW9N6VmjKHS7hLVtyjvMrgPfW0KR5y3o97NnEdgEklka1XhAJx7gJZtF/oftKeR
w606v46hcFrtRRhEthtraYU+ki6TMAWJ55EYe9RVTS1+SXLHJBMoKiSyzkOnNfKn
zczJp7VIKRwvcb6dUAs3pRNPKVuGkjToEtprlkESbSrfnBZCe8PMfSUgmVaKyJir
cxBzsvJ8JmYlpbpUuQpJ/t8r8KTcAn1+XMEPEUtLotAy2Jar8djtrahYunF9Vt+T
9wr+gVyYcu/3AxV+NeDiJh5//1mKWASj7JURaToKm0cE2BSrEfjI/Sg1DSLqtaVZ
TFuYeA+WUDDj0dulQB35lnwIFW55LkOzjlwj60U0uCo+gwWrxm8fNnU9l9qL0yMG
WJe7XUHd53yzCq8ToriO5n1NGx402rLSX6eeuCd45z1pPe1Xo6wv4ml1Sc01FP8J
StRHNf/ZSgOw4UNvt2pITMjbAA2JF+bhL5S0/09LRHdF8XDJk4bdpAzUpCigXfws
fb/fhtOw3/PEizyDk/D2Wjk6sp/Jm1PiN/c6tFnNfd4h6e5VYMluTkoZ3mpVcYSP
vQqsQzeo9Zt4bJk61UsiLrS0OLUaCxfQEo7fWTtEFqwXeH7P1Z//p/hglbqj/6RH
eHlNN+ncItKpwdrN8+gFFP3QMBBO0Bqp9otunnpp9wRj6Dd9xoJ7A74gLfjkvcov
xcfNuaKysJl8XkkG3eW3MqB9YSVrdbfwrzhvi1+Syh3uS3hMups7TRQNPDtfbkIZ
eZh5VLG1qafwSqdL4Ry2zrFXlUD625oG0PSrqkEEAY+EGi+ugDM/oif9vJb8EG3p
sjiL8qh4JGEUCQdoiKjqcsdRnMVJ3ZPQz3NGnj9423g6gqzCx6/kO98zBAGcwd76
iI+i/JWyZE3tycu/aDHtS+xXtLxDGbnqlhnRz1leabzM2XOn8xITmIIy59j5iZeB
dzsT7VTh4Jskb2T7KRKrlbsUAUOhW7K0LTDR9NnpQrM7f91fL7my9ohjpd8IruYZ
+XryCv7jL3r1u+ae5gfJnnhTIZIM4MoM6OrH6eexsY05yXllE45MGVbgv1/uVQ9a
5wugX6kJFuiruLl6MSV8vOFr6ivSGZt0g20N+L4LuYUS6jN+AXysDmaWCvLBWLnI
n5aB7V4iIom0hMZ0+5KDDjPEWfli+2dJLQzZqBNE9P7GposKcM4ONlWK7KZ6VAwt
HDo8FL0rudwtxc6unjVNKGoujTglcaE57DZk4wZ4ABU0/1QEtNqamk0x2icI5Qsh
LEJu7m9paN6iAYGU9b0NY2ZLql5FYU6m7p4lPY10toyFZGqTr2Sud5A57ttgZtHQ
aw59ImOx4Uy5HjUBEV1B2YOmeEHAe4bOqH+jUXoTdpykJ2HeaorxiZHkIO6aXu40
YWczBX9Ns7qMlQaw3Pyu0bJjxoKcUJEd5N5WtZZFqlC7rsj7eIcyKSxu5WMt+xfg
px8f04u+W6m8cmbVn+0eJ0o2qPkwV1xfOps+O7TAlFLYN5uI2fPL5Nvh7vrtCjfd
1QIwS96m+eiH/Tb01+nU6JNbIJQ1Wu9ITMnpCByTQLVkiD3IojqvjjDIqf8kBgrN
h7c1JjYDqUEMCt2W0MamajMLlQeJOgFCIFD0E1GTalFFyl3ndZavzcivEhKUWQHY
l7UkrF1nG/xl7BhU9BOsaZ12M+OmmEUfWUiEgfkfKt+AnVKompaUkPMjYG5dUvaZ
mVdL8HQ6alG40uA82zyTonSocrFpqYmUGvJ7XW+/ORQzVCkxyNhesH4QBIwd91+L
94Pxjqhm4J8A3w3jujLF8w+UrnRZzRHQRwjI77X56kx8blr+JFglzpnDfFnAKkaf
Y3a16UBdtMLw2fpIb61PCaYX/eEC0a3aY79gbyPGs8cZuGHI9/3M5ZtMRYH5vQgU
oNrCS1VBr3h2CicORxNZ+DqguUaFEKFXwwK5bwWDXewFKdMOGVzVy+YyyDlErsJk
YFrfzVV5CRxZ3RK/q3pl8u+jdY2/kniX47wgjLg+aKGV0AafPpLUiocYvGbMwdpI
vbA8JJHV+hAsEcxvKdNgpvYcHLGp5Lz5cWOkhd30iogohucqcUwBmOXNDoyzWnR+
kWONPuNEv3Y/MUi7horzvDFYxH+TP0p8GxU/cfVZZ0hkA/We2wogAzISKGHgpe4W
6b4ExGtKbIJSN/VrqQy+RtJ/rXrIM7MIwkZXplKI5ZzBodbxenxRdHVvOSClBAti
Ba61UIlhnRBPqRn3leq96UC0WJqojQCln08dlJVrtc4EinB6LTDorN/V4raep5pw
8BouhaHqe9DhTFzcGee+tSTZWiU1p9gT2RuS4zz5MoHzoocFRfBy7wpPn86MGGi+
+AjM2an7U+Un9UTIyLSTlgJoWdvo7rutnRc0/YYLrs0egooMccCKzczvEksWho4q
k2g7S6LczGvXYWQANVl99MC940dktqZUjm8+mIeAKtXSSVrnlMDNCS70BFzbVFfp
yDo78ZmY4Cx+8+xB+kWn3rUGWjX+Dj9eaWPARQkKsu8gH2E4WgUNhyBeinsie5PS
Ec6xc2NLKQDzuc22/wm3Gg6DgiaTTHMrhoC6E6UlrscZkVCd2I4u2iCT/JfWKG/w
QUE5Iab6+Xit47xhgcygOxciTRPUwyzULzfUB4mq14RJIubFqmT8M2Ro+v3C58b+
JQLpp+cPE4jO0y1fdDQWyOuYswtPGaQ4wJGlIqLHJX52GnmMUy+r4EgjcLLywElb
XAS/a1NOx4VcicEwUEMMCCtVH4Vypr5+NDGtz5vUjQhKx+P0v6P8QVu0huQs791B
g8zTjDxLLhTl9yVDZR6zjjWQ5bWXQMu0clwOO0/b1BTDexgNT+JpQ8LEE2Loi2Xt
xQbMwDPqEHuNmn8Br7zdXpjmPJWJUyx6skDoP5BdGr6ImbSqlBWyraF3U69cwffr
Qi/Hg+Hz+IoAcUihLunjiOaAXeMBVal+s3zXCXOEUjCDCuGInMXSVkRXh74Zl7Bb
gdXHDKI8DerZOODv6W/52O5KZzRyQnmw6D5EBvWIyymk4k+sn6WjT9P+47z/1i8f
zRg2UKZSvknHifAtuKfTy2I+cntLq+J8/kw2/54QaP++p5C3PGTqEpV459IYQ688
uT7JKydm4PLRGpoTePquMXEYZJ6xZjTDSxhlLcc6OQTOTzIuk44+FbTxuk5U54v8
Kfcr/i6tOzMCObSF7GkbLTH+mfk4Grc3hTiLghSsLiTlOrG+HhlrRVfD1N1FAUCy
fUg5jSo8PmbcKrgnc5R4qpmbr5pRelE83J7wmZd0H6mOpoPrpkEsngkUblGIRazG
NjSh7HznkU8zYjhoZb0Kkkuh+szoZb8Ah2fs7JlMx76XY/HEP6nQu5kWKYra4IZh
m235abbdhl5eKe8V5833hT35YDVHU2aY6pw423yTPDijszgwC/BNoZhOStxXfigs
3m0S82XpFOuCmo1UpFKAltEYUdPmjaObacJ/NA33Ul6BhyYv7fa1tXF4Xiyvyolj
KBbJIR05LZEySfcmq/Jqd4vkYrt9IgTYotdptNZnIRXi0Ske5zmlECc2kLMDt76d
JsgeKPc+IzwkOUCdt/EIuw7aFqHLtQHWfIiDvqhK2oL6fhrldsn2n21Z+TBzxMvc
TzNmsP2rz7sYOYE/r09/cOwutTsGGcS7/5lk4bj4wbixm7iGvL0wgpnh/FMYLuzt
ZQ73CT5H+ANcfkoI2o2ApR/ZUCeAxl3SG3rWMq89dmjDUGATsWmBUHia4u014XUe
b3IJxr7iImg9PWfj9JsG1OxDXAC4myEtzWSVC0lziPJSCMskJEE4us0BtB5Pct/d
5DJ7JDV5Hzhgiz5k0Rd8n5kY+oVo1BS5YNb2kn6e9PRnNvKMcNq0q6aQgt0D9QWS
wmChuafxXgjYssVepNH52y6IJOYmaTUn47CnLisl8tP+l82LOjNVtFnaG/7Aqgm9
h6c362G3jJLfNrvHwxXOXhXbpvjiQ2Ot8WNVfSzFVp0hUxScETBTJktKRgG3whf6
oRv0Hx99Bt0rL5RhgbUSK/vVZbbG0Vyj020srFtvt2+EACt8Ky4qpAw9H7LvTupq
xWc6zPDDVfAw+DXk8znIAPTFQ7APXzyQwoZxtRDr1TDgYjmorSHyodYD/fM7C1Kg
ctvIqfSWmJ6XmjKLxSKi7sQJooia+ImC0kLJVO91aaTfJRzSKhU8tOaOsKI2rDT6
AbrgzugfsHsmD9K7e5/ZnwxPcCQfWqMuzTGZIxR/eJ3zUcKRHGFt5GW9qM5XXQ4z
HyA2qGdOYCP4CyMNVPunm+KNXeKAxqhCaskYMrJ4pdjsXpa7KGkxOqyANAtbYPEv
6eKKaIlBbqbae9FZ+oMCrR4+H5QlrPudetb3/Gjx5QYWSmOvBriN4hNu5tZxN9c2
8ofXT2IgsiQsChAPEkj5w6pyMWVu9KKYVYcZBVuG8jVSj2essdt47pJhS2eU1NIr
85JR/xBxEf7adlQneb+addZASuJ6+GXfubsv1NUmGiYlIAuzUpwEAloOX86qjqsE
O36kPcKiFWuNKgcJJgaY2K1ljbuL9PDFCwiWpfrAl0Sps20e7vnhLk0O6ji9Jsrl
6Ib+QhxWn+mC5v7dsl9H3H08FfSM4GIKsJTBn2/Z00YlJtnIm92UizKOq+CSmruB
1dU1wwDPRGN4vJDh0lFussDcHC3E1V6vt25fsJhcakuLx5Twya5Ttt0L+ipvtrE1
VL2ZjPZRSzWOuZobn6Rgf2GlhcsE3LFpIMG4cm4ZX6oe9JE8ZhlutTCWGR16zB0F
kCBxe2m9aqo6ISpHSbDRVMZea4+xCXaBkEyE6NHE1xOEwP0UqiGYbgSSJYXjJPE1
g51XsoDiMXRqJN1bR6AYLnt2GXE9bhMN5oUZBCYMUXy/ryDm64f13ROqFmOaXns+
vXdOI3eGgRH7rckn7wWJfolmYW8hRRIStiIxeqqsxGO/9TrHT9DWXP6bQBuP9dNO
xzFA5W5T+oBuQhGjZJj35e4/vs3JUWQZ4maRbhmjJ9ls7RvM3ljM4rSXJDRL86Sd
8P1Sn/GLpj1EbjzJBAWdYwZGKHlTn/pG/tq60foJ1x6GmO/VwkGloPYSNB9373Xz
oel7UXyTYKgIm/iFJ1RfGFOHWDO/827ZsWXOY5W4TF7iTVX9iX/wC4xHID1NQyTH
4MQGSvXdbSAwthfQJ5tuEfwhRbjnwDBcTG/N7bA1+etI7ZFyh+eVSVXCtvfAKHbg
OaXoPL1FuvtatHJ47Sqneq2Zg2AclE5hAXzBZStFknS9fbVezL0DcDW3PhdPsJpA
4DwFLNBG/JwyNBBxDgtdTkoxojJq9PB4jYi+5OW7xlTq8ODlUWHbx4dkomBv2Vbr
cUzZ+acQ8VexWHzAUin8V/0elRZL+fD+rry9vNXzjAR0PLDuHQwOMyjPKIJ4GMhh
yg7LnOEWOf7upyUU91Ldj1p3ZcbJzz6IZY03i5hOIeflt/0QxmVbZ52Bl4cHH8pM
8N6HJkxe5DCCbpyfEiQuudAvNTQ493HOYpbwwIQk46S/E8vOOafbx9dB02tx4oZA
qbQyieRamFkAMO+VD91k0Ua8l+vpbV8wmFQnd3tP8g8m67gh466ZHwh4VlCOXQkk
f/Fuytsh6863gcsnGd7X4KEJtY8pdbp4E+cyqtVdKlghl1oUISoTcv6PJVyaEo5c
95WrqxkZQJF/E8zvAIY7XGeGAkZWsLZYlmCUY7F/WKs17lQAgyPTVcBzpEvkZw9k
yXSH+NJbYWM22fw3VOdMDpDZ60dClT3eGEwb8cDAA2r+1Zc3kgdNHSKy11wi9L7z
HuQ/PM4hie66pVZpctAhJhM3sqjrCA4LO2xmdi9tDV8x1u/dqxYbZXtOy4srzvvu
QNdOteGyHf7VePMjzVP7G+NP0m7Ko2q49YqutIKG1FOroJ9aG3Sqvko8fpjQjn1I
Q2Mlt8a5IEpDucjz/aWBE/ao4mlCrVf3nW99/pW4X6WfV0IIE1LhDb/VeqRLiDGh
FvZnt7c9V0RI+yo6BYGJjS2rdoZO4GU2sT9w9OAmG6bYWv5yHAAyCrHw/pFnQ/dp
51+ulXrTzPxWonAyJlcT3AivO/A6969LWtOwVyG+en0GS8R1x3oi23uByJG30E09
BeHccdE7rX+baFt+StSaxUeg20b59YAydzesGRmJt3Py2vGj17Yef+7QhiKEuock
hO0q6mS+csSfytSDpsUo17z+AqifGq9iY3tSrZEiD/p8XS9M3aNmumY2huumsAji
9zQ/u9l5imLTNXmB7wMQC6n3Z1wPd9QGRS/3pr8foHDglSjIl2ZRlra3q5Ylnuw4
hDqLxzMp0L8omLSWvUesX7DFQeXRCz/q0vgdR9Ciz6f7k4yzZun7kgKaGFQmn9tx
zB2y0J/rZq4extJkQvCysgmkLU2HRUGiqxECgtFbFSr1moa46PRXkJSGoiRi7XF6
hQ9QoY94fq2obFh7kVRRVoBPE0k6O7MpGU3TVTnM1ObOmnE1KvtOWmHxzawm6NBZ
pAl/zCnQxbRh32rvoEz1HWWKl/W55Qr1JVHiWLUqFAr+h8UXM/UtAcqFSgFsOWRL
DNyT9uqAPVRy0/l6vC7HJXhIFisAPE73l1arcYFi2sfEa8+JoPNw1hG5BXZEsGBR
aeztYw5iV2cHnJGc1oV2U8groZ+IKEvGxCadeUEnhkdbwbPIG/AwxsUI7f3NPdjg
ZH9f6qi165x207d+cvVSimPzl75D19TrzXzS/Sjn6x9u7Deeae+z6+lqOjxarwpG
g9Tps5Wxh2Ss/3SqNAjhZfG4W/BH8uQ5NkYCCVcp+P8WcxxM67o5Omt+ufFOyC/i
H9rihSxzd4GR5K7WhTuH3Wr2K0trvMstv0NqjSgAwSUYglOhsRmDgVaZmm9FDPTa
lQ+k5r1e1uWhuCLtGt2Rbc58n9SQITJnj6uODVMSehtxIaD5cXP7vU0XC/7QySI+
Jcaj18PCOeblp60OiHnKcrC59CgbrteF8VooBFgVEMW7579apPerUeBXFrxOm5QA
1DPtzL36XfwWDs96Ejl/HyZz3S9cwzldXRxFhqjjZHE13ZZt1cd0MYAoChngmGUc
XkKw87+6gb3xRtvIJqTpnNWk5tbxPfSY5FgwQq6xdwj2+TarNEkDTOgOhUHvbcWk
wzTim55fVc/djrQt/DQtEpOZUN05NT10Uhx5nE3CG/+StX+jsGE7aXo+nmEpb/SV
M+6OHqIk0YzpXQo9qUdBlolDU4FG/5j9H3ALlW+a/wDpxs4caAphQZ3VU1NXiqN7
zeCSFuwoxZaTGZa8DGQvkJCbO0y/k1p2NcDPBlfGmV4anSJAhmtbFvtdteaHzFOb
99bBvSKp2DWZJZJgEk20VvN1r2YPxjLH+db8cAuwfH2tIN66YV1Vb9hoYemEsZv/
YC+XuI5j46mU1JJpsyTREMcQlJpYUNro1QVxzyXhxpaHeJ0w81Sez7QuVk93EcHH
DZj3011ojWyYck1hkQ+CAR9vYW7zngTpuV/LnFGmAA1DAIKmrVHwxENFfZG31uU4
zkSA9oVrCLSweRumGM4bNgWas+v/tYj0CGS01Lo43k0zqcEUNy+29D4eIhf92Zka
6hy8uukc3ryVClN8PUPvH7dDSxPLmNDX0F3qUpy6xw/GsVBu0D+sqbLlNKdUa6ha
CHvjdIQen4n8KPuJwlvRHZ9R1k5O7Pq2L1b6JdvfWgkouhe1WyXY4e1imWcopXpc
eLAf+qV0EElj6MIXJZzxT/XgN2f9ci+PoUb3g8mH4/rhPxx8UxLSZtKDNuWpk3S0
bSqyIeZagF0FfsWTJgszvKww/YfwgXehHuAYHoak5E0pUCxCmkk+HvPCdlqdJ2cq
Zk36ZxWD1cwQGvX/g/JCYw3NdBNJYRxquyMSJIYpIRdzkyeAaWCZo0C1L2ZKfrDv
Zp3pljyzY1gio3zQWn9z5lwLBAVWvX2d93VwdrHcXXXA2dX0Z4D29eo8RqQrUZLq
nKZ4+oYTPZc7VBh+nCjJsUaN6EWNYj9BjXVyNypsgn8S07kCDC1SP9yfHAVCoROt
ubEDFWu9xIGGP8+/9vLORhoN9cQUfN28Vnpvz3dRWKAA8kkji39xHIdHLtYliVuU
wwStEH3o+Y8QTs3NRrm12IQcj+l4XrBCox++Kp6Fjjmg9xZt8dqkYduW+/9TFgum
rSbYTkUYT7LUMJ6K6mI8fAsq1tz/zIUyzWMv/rtpyGWTb6nTeBWQmb4dhxOelIDr
C42bnZD4w8cGJQf8h1Gke0S6IAUspTqen7+DO/yNOsigQorv46isWCYsHE0KoIGg
tzBGaDUlY8Y3vu+u0hbgiBx3qaK/b3iRDVHBiVx++bGJk2H/zhLm8+3MWOj4T8A5
PDGyuXy5BeiXlDLkvLttTYC/Y6sEsTm9fLCoTyyKWevR4KugyKXn8jvgfFGaHzOa
wWNqC7mDlnUBAhcho1jHC/7gmlvZNW7Ppc7liS31uxwgrbNSG3Yh3Q8bunZDk2es
wmrXh0Ek/MWEQCfHKtHxP5sxjMOFze5JkRHHsKXGNl+t7YDbNCP8O/bwV+X1iuFD
bqaO4yky+FVxDesYSCRAwF6NZmPHxLnaOvzSh+0OiTIw5BLQbC0+kLAFGA4YbZCv
u9zMYl0Ip2sj2WBlK1xXaBdre+yngPwxdnWj/gBmHh9xZBmuDvm78tmf4OJ/uh7u
niNSyZO+FUme5qUsc3+RmccBhjfWkLUtItE9mmRJkoLsc1kSnUXpTEQ8klI1cyrq
4QGdmVOZ0Mmr2N1FUvZ98mIQtGiBeGqPD9qGfOVwL/q/SZfwFLmG+ivJSE4hTU2g
P8PZyVvGRK384HDvwFHZD1ESu8EofatvYZ9+V8rirhexiGuyGQUkmK5s/iAHtl1t
qnFjKFF0JWKiOdy/pdNFWD00Edq2w1LSPfjFgMY5iKh3iXfShslxj4JhDNOMpsnV
6vyFQwFZLAcd81EHkBF60NeHvyvtUmxiuE0aqEvK/DAgyfzgBu/og0ISckLXGvNq
htmXRjC24KpV5OqzlnrXTjVXGNUpdXCe3afOsftaMIIuuxXPMQFCtm+HzVP9O2YS
lE1HKX7ATepQhBQUoWcMmPBl+rEVGmAwxx6FHkv2x8JMpNz5hCSjEW2+upHCVXIO
CLxCFAC+60RNSA3hFX15k9lTf0QGks9e62d/WI90tKkyzzLu8l87KIvUWW+otQRu
/dXnY9L7IJ39YebgiukN8Bpdb6TehGroy6gFisXw5Us2wCKqOESLU0lIJThc4zbX
WPHrPrdMfWhmKPqw4yg9MBXcMlV2g34KY+Yn8yyuEf+JATlvQO4N20NAI+YbyRuo
D2GnWNBBobtaBsAxH3vQVGHWrmJcSVAFwe6md3YTFXTc7jKAxvDhQ0U3urIgzMwc
D4PX6LkcvamprNJnwsQcnwdr04+ucB4CQ6oGlyioOIuljJY17hZNfMtL61NYYPCm
sCsAqDn74O6AlMGr5K0eOZsX1xhe8/MXMKyOHfUO0REhNo1p/bb6sNtvESY9FkoW
XlgNjxbou7MBLsVg3q8U9EUCCRGpaA88W3M/VfT8UnL567qkZiX7TwGu1YIQa2PJ
3Vki6AXN+dqFe9rzT/ecksFYpcs9kfthUNPZYrpu7JpVhyP0kbmCRfjnkSoRRBiH
N3Fptz0mudSNor3tRorUsdbpsw/T6uvSZ1RScX/Z3SmAkoXx6rQ5FOz8Qhm/oH1L
ptYL4ICJEQy6ARYwTQ7DALgBVPAd9dPEni6h4vtV0KntuKG34HH2NQwQGUBOYOwS
1VAkA7e5o2LCzEt8DsCPhUPJQFtEy+hl/yEMCfn0zSChWRkDP0uyw3mX1FSTkffz
g47X3H67ReyCkHeQtN7P8v5iofcGtM7iGr1vwukbM3YEp1fviuvZrVRzjfRghfFo
O0PlDIENR28EPYLcFju26mizU3WHMh6w7xXHVAL3BCoQTmfoNepWOsfMVgUqI0ka
fJq0wfp5H+KUH8gUdcKZjd/g2PhMI6RYKEpmII/WBaNuInIQXh/YwPzrM73r3mHQ
4TivqEhrfZ0ZFeOXY6PvuLQ/HZio7dxmOO/kKbChgQNgzDOngy2GBeWuBvA6ei6a
VE3ITmov083754XMrw99wKPplRGGN3DdVtUSbIrPUkoKV4sLBj7dMytOdMwz9EgM
an0SA6/3QIVja3rVPr9BuK6Mxij2rSNgh2Le2fquksfUcgsd9/HEN2FWKSMAsyUF
tZp3vcXGAaD4p4iLTu3ggA==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
QMzTMbBnKk6gOfDGmEu3ifR5e0zRlDUobuTmz/4IyzhVJGtJrbjoXwhmh39dFOJ1
30oCsPDKrrPmAl1YHMa6HHMQKM8nxJR/qoC5yIgGc6hdYqhpjmWfGLrh6jgkDNgI
7JrZbgRZnoFGuQvoH8sgBvT4gAxYuzSuyVe16cq/xck=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 218890    )
UYBXO8dWKRBx7T/rpInqzothV2BntvzcgR5gpFw4NsokyOSUnxX9m4X1Ii1/ANP9
A1ogSjKY9WTun/5pz4KQ8ud7qbOnRa6N94VMgLzJsY5UEoQbVxrEZIBymSJpaOxK
TzO+b4QfvUZegR7mSHTZoyEOEDmSgp4P+llVxyZoqh1G4/fmh5gfZhAbXE8QTDLI
UMwmLIkAza2QAOfCWYPyUIg6XWIYkKWExlsaZZRpyKePfobYl//q/XSgtDBJIOBo
jleGD6aW3JP+X3SVoqbyUw6gvjE9ELhy5CxDM89XN2kiR1xiKB/ek5xvlJx+46AH
`pragma protect end_protected  
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Key8IbU/BE0sacfBP9huE7W+W8jDhdyKXlC7Ln7dlrobH3eSNXOKFsKaqGGsdctA
JarVTnOIbd6wCL6eU9lfnE8mEpFiwyVQFmAUXV4I8fcmt2iuoyabgM4ZrS0zSFmq
fPBconICzhir02GAd4FJ2jZpOHZ2vkpawvfnAWDEqcI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 219023    )
O+3CkqB8i9NSiOOcPs3DJJZBh3yizNkGNfrnR+QaycSVy/6V1f3s8rfO2DfqLyJr
0LciuepFE1b+fgHzGSV/tiYJTCCd86vvKNc70dXwUtDnNDkdHCjJjdAeTBPBRTuF
OSXYLDaCqOk3141/RSpCVyZww9GlCrkQJYOzv8wgU96h1jaKaW7NfRnWEosBB0nB
`pragma protect end_protected

// -----------------------------------------------------------------------------
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
grJNVubIleprPDxQYCkRqIJfzH2f2IGybPRitH59jszgfr6v/M1Ad+jKyBwc5f6Z
tmUFWK7PZypB+D/og1jrqna30NeYr5TnBUqXfxpXdSa8ivospNzXTJGZzEpMVNkX
5e5tKIUCh9NsdMiKDXr8pVE1tPLvQR8VJysFGYv2P2M=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 219189    )
imoFTyZYNbX0HGJDKB4DX5b0MLRPLiI9TXvAe/SVZaZogZzWJ1MkECFiQme0sl3H
v8XSc9524EJElIbfSQoh3FLZToh/PqO/EHy5b2S7EeisvOIN+yyzmi+rbZUBQ5Nv
C6NuoQmcoCelApawa9zWhXTgAqutlGeHt0W0uO9HG7BXPipfjBIxg+PzEL9xHHZl
WnVmZZghVFm+XzXlwi3SGfKcy+V5ih+2G9ApciW1Atg=
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
bNkKeVXf//DIHQ+ELAWbX/1cL4G3Ux0FORo2schtF8qtijAzJoBsKqkPsByYcS5d
vV1m9kknt5QUyl0YAaypT5S+7lsJSZm479r+4C8m+NCoE/6Lr1JDzwOAd9RIUVsu
A49iHkPlnyHN7Gjv60EBjlFdJd8LXSV/+YfQS9Ii+Ak=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 232711    )
HzdsraLGll/8wZ8la9xo0+qh72dedfrAilxl9id5eCmBBhSeZR/9mYBofhuO15Rq
Jm3G8oGP485znRtrTZvIXeF84orm27wpJtqfqqiqjZiT0bO8DIDWOqA8b86EwdLb
+61CsY8j9eN7GV4+Fyf5pMB7JuXrrvNgLQfT9e7+h/bnzk2NX+6ui+UQcnvb7r1q
79F+l5nJcMm+qCKsY8KdgKIWJQBPlyluFEWT4WPSJS/819G6tLIMfmd8uGPeYgm8
kyEavVD//973iYnLgymmNxWI4editisplckWlC+Ecg8Uz44g65LBuK7DH9/OfZ8D
nADmtbkf+91Z9r/j9oBz0k5bgmm69P03ur5aRlsJTjArfSOHeMpW3bMk/W1pFK0L
i1wfX4cQg6iFtxqmKc9JE9H5KNQQA+RIUiMWvB8z9ZINs8h/52dKwGsglcRZAl0t
ZOpLWccEeGvu591hp/sSNPv2qWUaONP7ek8oBZzYmkZXxG0r5Ps2ciiRB7CqZ4Ud
Kb7s2GBTf8bCK06NTHHeiIStA6qh4YlSKblxpUBW1g0H3tzHz4Wj95F891jVGfu3
2n+CLsydNkfhD0pYFVMGcVCsJjmRa8BC2HOv8GEN0OFTQcgSr17Sp1c2LaDqFY5z
HnEYPGPUBOPbdsRHToQmejCO3roz1tgX6C3xxXjxyBnIFOe/qKAdPYE+6r50EZAw
1aVP6/MHgsnxa2powIaQ84vJ6bGFGuyxqCb3AyGAYFUd+SujsFjLSoiSC4is6WTe
OHA+6mGC5QbXmZ1iUcbtR3GoDeug9pbpNFV7Azsk/ToohdSUyS5s5C0l7kTaUrVv
pU/pj0fTRp5XO9Cu7sY1LzlCyllRTQaM3YEs1SrmtWZaz5BB7Q1nre/JY1sM9wlC
3dg72PsXtGrzfsYbGLkwM231F5cswP14Jh8viM/qsKLAzSeI78PrT8uCE5vTt14l
SILChDDyJsv/8Z54f3y24freH6NbSwdnNXJnGQBAmjOGUQQSAZQN+uOt0156eME7
56trsR0sxswonD1FJ3EBb6UbICXmvMGt5NJfZfjf6/SLqZuvaNqmdxjR0w262fMT
nX9yniMgICrsI/2D65CriU3yKOwuSNzR2z8QlG+ExldTg0BwCdH/C+Eb1wKzeedO
fUvLSYhfGl2EMSRzWcee8ktvShsZETluj2k9zFfHxNphXcYEkhVjddb6l2W8hbB0
YBwQ6nA30cnmHkDrVYqfxQRtm+irVROo6kCeNvriiYqlqDvLyEtWGh8K4IDU0u4j
LtAozQft0P5MQYCY1HWvyntuo9gx7AnR2gnM7zRFwRnBxWN1erkRodgdurTLBg7s
bFhfj8GzH5iU1e6Qk525uhfwltkcmjefahbBSNn5lOjo7zCM0SMp2ojthfHKzrw+
lWtq4LecxUnrP+p86tPGgMm7DdyHpVznOMgfnqsDHW+iNI8mUul5BnmGYzK0bzzM
+tPzMMSbMYwJ0BnVDITd9xNXmFyh8yDl1/iND3uTGl6iNruipQCacogk42G2KZRi
WsOL/Jrl2ld5RmznXuJRtHVNmxfifCuVvYaTPRyGHTaqlma8VSl3gFW4edeZXGmP
isKAiOi2iT265z/seMk+Wzhvj8fvwtazeiUdApliy3w7itI2C7jbV4SLn0BEE178
RqFC3RWHE0yzXp9QebbKkBbAm5XlfmSaPRBPbUdLpyKIXpXlsVFsrAHoCDnktEff
k+IzsgXwW+yXDl8Pw+ATgbVsus+3BD3mTIPSMNBwNblUw9aNFym84GgJEK939X5E
vzoVIgZ/V/PiRqFsD/OH6r9XbUun2u7jtuEhdzxiwUTy6+mMKwOt0D/wk2ra7/Is
byL7AofE/wa1/W0UGIwXUGQAvdp38nNMbgXkcSc1Z0JBrf0j12mVMFAEy3LEQk4I
tif1YJ7fzJy6WOqvvdZpYKABgGUs4KUoYq5iAKNVeuAjx4MkDqP4Ski5MpLq1zeN
nh7s5ft28tXBJ2j+XMYwiAA+57VMoTZTAfJWuwJz4Wto5o8vCDHM3Pf0hBHGggem
U1Cl2hafxp2Py4mrMos/wAKJyeAMvV4mzE8AaeXT80y+03dMG89Q7CLNhdW7Rdpk
kfsu+lSRmQXfFWctzKHmZCqcriOpPKSYym9tHqQa9uYWlyIVHUFkrxk7APwU5O3B
sSoeetQ78aHgA+1jp0T4VeS4r64/Z0q/hc2F1uVIPeQnpyKxNxHNYY2ZCvhc6BTZ
1AWrp6FfA1PYyA7ackkcwycTBu+AWNNoX+1LsY+kU+APVwDU0Yg0IYUgNhiN1zjk
yyc42lm95yITfEZYTKfMEABR4ET+rhuBc2Ioz9JLLrdQ4Bm08B35wOU/DHKuWBCc
JU+B1vmLxCUOkgiu3YLKyVTKstf3qZTMDPFQg1QhH25VQIqcaMMUiXJoOoFDRap8
pi9GKp6n2z/h3P1iYcg6oHikZc+Vh5AGIh/AOtDp6E0dMDx4xEMVQiU5iL5G/CYK
e8/TCO4cAhqK17qlPaSnXCiYbERwFsH0OHMQho3DG7sxCZT2MKFBXf6yHZLLgIat
sRdfFdVDh7cBb6DFI0cdoHQKHu6WCTIyuaAbS0VMeQr4pX91Wi4Oqe6yHk9rYqgQ
yUa4xCBje8irw4zfRWHZE+iDg28h9xvtcTCs08pzDM+Oz+Entn1fMsBOB47Xa0cS
+nUODirfZAWy1opjUZba7WfiR5Qm6uzjyAasKEFKdOub1WHxhhEmqh9i0EvbKwO2
FC1KtU6tdwGKZgYM28gz9MpmJLdY8PLN7GDBd7mr3KsH9IGMJFHOjuZDE2pS5zXW
f7pLIsQ0I+g06kXZDnoNd7swWcwJTBOFniOt9LJ/Lszzc/9OdnV5OPu4rVTS5EtZ
Wyu182ETu53dMABsbEC9ZZGB3BVKPFbzMxjuipOhRXWW1iJN9O6ZNcegP/1FwtD2
VE7mdGM4udXPSgyEjdOFj3yf40nNQPxbG4kWZ8m/mXebGRFqdDtLc9/jjJ7al1zX
DiUZaFf/+DboFPVh3aNKm8nhqJdXcAVnfy6OYtv1gUa7nuEgrHvoVnMuJruHS1f7
xcEQM+mKU5So8QCjvzeFb+omiSib9M8uICID9/zx7up4I7P9oGlSg7JnM9HRGJQ/
FO18WZhZ6GwhU/w5zZVIXouh8R8ZZ0WYmu8ae/li9uzDYo7AlxpG5MLg5a69Qq93
CxOguI+4yvPVf+F9bmu1c+9ov568Q4+2dNNDKtHoesAlWBFP1zi87ZeKdoJ5kcyt
ou5udFyApdeg56MP3TnOAy4369PiQWpMZVY8Pzcs/G+xsXfbTyQDmn6VsL1fLq/y
WvOnQJSy6l+Uh9gP3rlekPcYW3YssYYER0OghwQoDIOsYYX+k1pDyWG2DfIMwEwz
xMI41sY//9nOV9j7yXnd1N/0XtwaCOpYT6a1X0Do4rnuPhz1IPid1FeE2q5/5C2e
Fia+B88w6WxdR9UB/P9YumxdzVGJjotiiGbCIBXEqtgmpxMaQqjJYB2G8bsmS3c4
1QN0AH5D6dp6jHt8NzHIYywZ14jLhdOIi0a4UbxUbqc1NiZn9vydbc1B1Hu0JBci
bW7sywJAvFNiiYkesmrdLJSe9cQPIumKZCfnAWDxgSebaC9Ks0p+aCB3fs7sHvWa
PttrBrjgEFIdMeqvKIF7X9iQCwaj5af7yXz6DKNYCUxaQN2/C4ZOs5X/Qhxj9Scu
VsFG0HtFFsVgrmiVlU0Y1aDMM98p+pPdU9n2pLuxDI5upukd3Eww4seg+HV9CnUl
kU3RZs2F4A0iD7l1sGv9+I7VmLcQjTZDS6lHMKj4XHSj39Ew9I2VD3QUxUGBft/2
lH6tMHYZaWF/kK0jaVVkI+ueLpO3ldv4IhEHKE9xe3CFjAoQ0ts+aiXyKUV6QEAU
16cfaK/VgkviU0gcefOjVB385w4+GfAr+p/hF/q5DJqtnhtRf18T05HDmmnHLab7
hBsGicnj/QBHX0or1XVAD3vTB1GDwGoCIkPVYMdDG0FP9b3FmS40cnbFExisGmPm
aTFXZ2rFEurygP9JWSPe5xpcDfpqWleODQePtcwQgyvcZHywrcK/Xxx4jSyjt617
AP1So9Jub8RwsJ5Wh1mqXQCoyADC+EfiU7TocYjOfsqLLXh5MuSDp/U5ja7oVijj
Gg/DgSvSxpoHuvJ3MB5wsCe/KJ8JNJ1U6J+DzwOSiLasCCsUutHt0HySDaDscwm8
DEAYRfb2GUQhbmf9II2UHfm0P2sfWzj2f4OBdVhUAoSoK+sea8vYRIkVTIJQL9ZW
fqyW9BnxiooPG9fwCYh2tN6p7ABWMQmqp4Gq8CTBFXoWDoo1zQX2ozvimlj7m3N9
7RcMdu2UQCi9dMjM+uzM/+5Sas/VJWm9+hM5krbIsCMc8le5+IxShaiZ38Pkf16C
EWFrjUH2Bq3vScfMV2QYLEIPw+PJ46fsHyliANGoENF74leb6MyY/MfibMFTbj5y
+tI1J0lhDEKj+67puo/HY9o2Cu4xKvk1g2UPgGyR37hWglhMHq7xJ4+Frure+6Zc
2uGd/bDedNVZgrTQqDoUxnIuHhewjU6xPCWRgWcfNzKlgiBYfjz8HgqzsBPq2NXj
JpdCL/dLKJKDSP/1RM0c75fi+Q55ti5rpb6VGBjvH6WDLwm5iX+hHpYa67dYz53i
wT7bh/806otX31G4ZKQBvOZ7bSpQiCPXe60PR3lmjj+XeYN3h4mnvMmFwNWVmsw4
a3mDG14AZzGB7wcWUg5ZZKRm3E0R925eCR5wAoUiJ23CxFfhpFhWAQnLqzlWN+kY
9pAVTTsWm598AQFhx1dWI4JNwg1Cy5gh+KEHeEJ/khDxWHvBoiFXwdtQwp23v6mc
8E1bccMfr/tuHUVGnP+7Epm8rVqIB+RNCX3f+UpU5qKzfhiP/bYddLm+mRpom4sI
vseXTUqFL8tbNd5jN4F1sgtfF2pdHnxU29iYBmrLNAjHF6I4hrRg6uTFwys5VDG9
9ruThuWncAgzcQhtVGC/3oC8lJzWECfn//oOqOg4qAuDPf55eITwYO8oSMag7OGM
A3I/MWn2n4FMhgmvpcvRhDuhQ2HYYT8L8KmL4bGVm4YVmWWY8KFGAUtcITBbOGyA
ynMxVqX8Bchju6NnqFb8Rf1jwdfNFy14L1pBSlfFRBO/KtpTWnd32zPH1KiN8bmO
CTx3MHymcE/OVauzqkyJH9v/+SuD2tMegmRWb0tCumitGCwT1sOrHRh6anrIXdz6
PxpS22Q6EStSIHScsDs3g8PYLEfBs9KxEYXCJCjk0lu4oqU2qs3MOQAnj2YRFM6f
CQfg1U2vkzEIe2FyoICnxvhKVlS++eoBZstcQw/7p1TJMpyPcqTQ2KshIadp9h9v
GACb36+buzGP+iJ4Y67NRqtMHJX8dLOKOiYUYYiVXxwC3KHVhvpt+aLHg9FZg7Xj
fZYfB9b9NZQyTnzrTWUA4RTaFcZJBVi2051j+kRVQ6l9cO+TTOXjGutabCX67hiU
QX6J6vfR7jiZOcWEBHfFEuD/BOpyBg8w6yZp/C/D0mZn1jySsXNXJUEfLMRpDqdK
vl23v3k42eSMbD/zJd79CS4xjkDBvfjyTQrP8tWX4MuQ3M7xtnWeBurfAI0HwXmq
NEmVQAjRcGAuU84n9rWhwcGwuxoSeJSyOspGsF3q0/4F/Z+CX0jV0oSPSTpkR0N/
asvaEFyVXMpxmCkj6mE9qOxTnrMBZC+7TQQjMJiUnoBsGHoXFWG3cnLrLUIrsGQC
xDsiHZB6k/pWT+75lWBSFmmGZauqqd5AI+OtDb7f2FDxjJl1AgSe0KT+jiyHDwW3
mftC3EL3CaRWUtB42pQrSYLr9bXWAHMxx3OYRy/M52xiGg0X6Qsn4lQoSST/9zyc
grJA2YuSuQkTs5LN81OhdDA3//RcRvJWpETmRX3/+8yoCaNO2nKMVYSad6HIOpE1
Yt1QeZbGV5dHO6FUDh+SgVytQcw0R0Fqrr+bO6Kqq+8pCerR52ng5sMCvPWJTZBy
fsUjh0Uefr8yXUsyCDkmWV7NsG3KMbJLBcQa0v7mbhEi5cuHuydeOU/f15OZpcVX
Qw1IvGJ88FeSaSfI1zJvJ7Mi/QrsF3uL4Uy9u8vNcmxBkIJU5SdzA8i5TfiqzSLj
nAqkc2NSve273Dndi3LcECLMsSOJm4RGC/A+UdGyWbWcMHqgPlzcNMjFhlIOamRD
5SPRPR+kSJvBOk3Pk1mn2A7GhZE/jOvlKAFsPDWH7c4D0k9VVr0iSnndSE5vgw1I
ibcW4kXS8yG2uVa4yqs/tmYuX85po5qXnICPtdosrZk7YXC29c/Pg4laFW4Ron+a
n2wYtLNv6KtmbWD4JBsaYV+8oM2QNHWpP3JOVixnq7gbx40SiyVsyx59MAjnT7kQ
9pAGWLjQVxnH2zLXBP2FVb/VsLU44u3n01H0ZcUcCz1qic1CJDkoEvgLjr+zsp6w
cbYEUd29kkME/C5EC5DvA75tJUyV3LGaXHljs9fCb0vtUnGNxwxeQtIAl+sihpOr
JI24JVubAgVlfStcYx2P+svDa0eQuEGD8iCrvYQohjIO0fYZi8e1CjqhkNcHvCU5
USN7YFy77+aenN2r3iCxVYS7ssyldDffOVURdlF7SpYSsZ6hbfgMbcSZNFVWU+Tf
2IrxFW09DXt3ig7P6jkg/sDFKhOGkwKe6IbP3Rkk3KCie5r5sJeYl0EW7bPDb8j/
GyW28wOFJOdJVug28QZnqrY+71EC/Nj1oiTcsSnlvQ0+qiRT3WAsZoA7zGwBy6Mi
errfnX805NcZMwsLgaz+qCXlsMufNKyoB55/VK7XfuYBoHIrhaNAEugt+lhBYfsD
qXhR7QkNiBJeU+mvdZcDj6JA8eExD3BmsfQC61iGxDmQ56VWZ6PrHDWS9wnDCWFn
UF89uD3l5t9eWrKWhRSIZ7kDrhZoS94a29/4LEF4k9DIEoxejFSmTMto1mAQAlOw
XupVHSnBnoJLKtowWOsg+8HyZrjSxMLDCaYdhFg1l3PbwubClZ7T+8i7MTF4bFE6
MxKxPB4sKTlVo5nUo62gOGopUfOd1DNa3H7joAl50r8uNkgVZA7BO5Z25sFG7/Ag
ou4lAC/8Tn9KohcS3/kiT83xhfQ0WasxZ3S9i8OlZkT/DeIV9FT2BPrXt1nh+tSQ
9MxcD9mCo/K8mpwuxdU0DZCcI9taZLSUW3alxQkltgiwoyzrmozFXGOXkourtEJA
EWrdE31Ggbcml2DQ1MC0FQsvWP5ggxtAn+2hP5QM2S/MgJPv5++/m2lf6cF594cZ
9YmkanlB9oZ8Iidkog2ThEtkw0YzWGHc+0b1RfclG6JpMTEZ3E60Ymv5YQjRVLlE
d6sfalXQ87s2/oEqGo0HpZhSEMRLmlJlLMXHour2P470KIwvhrR2qzx70biAke0y
U0qy+YU47nygOapLR0iP64egrzcA/DjOzDetnmzpBp1kZTj8Zv/0zuPKo6rVslQD
98eIhqGWrnIQg8kWRixY75iXtHHmfIUuFYJdH1ub5ufHmktzC67e24E66X0lnIdB
SU/TiYo2ytxgL4wxliratgSHjxDVJkjGsfcWljM8bmKtWeIgL+C12QSNQBfO8ArB
uqS7qtkAIcg+UtYBiS1M1pKcq9tmMDbPgypvseVJTf3PDs0OYeAqVE4dmJdUHRoA
lhcNDcZm8dAhIKS8c46BzgxUeTQKYrXQzy21PlfzvgYdW/+CIyhowNlHjgD+cgHP
vhpSEI4YaVj5SQ5QxZQfaZy5VFhhy35onb/eljexOF/yhdvEavWpLDzyo9uI5ORp
M1mNYo2T3/k/LdNNgTE5qPqVeGvozyIzziU8kUN0ukLzuqaTgw1Yd2ewUd0tKpCV
tw6bFJrNoZEYwCwbKSMQDZrb/COyuSgKyMffz/3HLUrKNLQzmgx+AFMrqN/cmt7l
RY2KDeAjJVNnbdln91ZS5qX7mbmxmvclgyWgZXGjBiQXeb8Trj6IeF5NnvdNKlCG
I6k/8aISo8PR7aK19VK19E/2VTevz5puc/l+JGDXlXLcEdi+Bml6j2C9z55TWbNO
ShWLe3tOxrqSOSt2KjCjiqPJxpjvfpkTy6asOc/RwSayCgxHxADR2bF5UrW7IbLe
p2oq2ND782tf8s+phmLjcvlq9QqfYRhjpQxRcC0L++OMJu9oOVnI8VFI94e8vYwJ
gO7K1Cc2o6esYIE65nKXWht3EruW2AqBELmjLV1E4OuAxqDWzLCC0F1jmnFxl4+2
j7lF7fxpNrFWztWgE0HYhZifXfjd67h0a87s7SzgEzWiMN77BleO61D0KuTlZe8X
rnB8GVRX3MQ/eOo/ywfd7JxKHvoziRhUnKXurPA5GJp+X0WbVRM6qCRyVEZ9qE2I
Vzvg7l3c06ICtZX8aBcf/AIKJPJE4TscAjN3S4QfMPX8sHIvMGs0LpAf4N5kWcyk
DwtQ2jMCKva41BLgfo4/LxQDD60l2Qwvaz9FLgmab/bvBWVsoJ4Jx8fcxz8A4bn0
olUVEfhay5VDBmRxXKvMmM+XxuLTGCl7gaMr2B8OlceKyoZhUTWaypfSRgNALXQy
ktEJxOgXATlYdlKja0BhJSLL0/0billCELabwrB78fao5X2P/IR4ztjVw9n+yM3L
Ui5NviR81qPkdymEjl2Ag7JwtScHlrxJBE0BpSEHG4f5EMUVJszxUaWgl6b9M3AW
9GVeGZ0bdqcoFmWUICiZruAns0pGCkcZhABOu0dfo63ZuBYH7Q1FwQs4I8y9LXYb
M1P/y1haB710avGGDJCkWUCZO+mrvYwvTDsuFaeCSUUBOwzA7MmWjTmtV7epp30u
BhL3Uv8ZtkxHkTjzPP1C3XD8RxaBJYa4ECeIZTDAskib1Nt1QCno51Iyei7yQOMn
nzP30Fr3bdKnugW91YyIye/HxZcXc0Jb2991xVNkcuG0s76XKjDXGLBBSlb9/ya3
nchBAqPpSmkG6igiR+c/DPvqhE1vaG6Hvzo3EGagWqu0LBuXmo6mKKX+2S2La5T2
6zU8f38l/PRfsyHGniHLKkrdNblJxPoNQJ8AkInz2av01sUbpuJyGZ2MBQKvkkTg
mZGyOAhwaD+tMQMaCJTJ5SQb/dz5jPhDXeDCO5ayaBSsxRhSSouUUh66C6gt48dh
TgoabT4Kc5m/MAvOij8g2s+ZE6ugOpTQIneraf+m1fdtRzOYqStyKe8YI7zrih/g
zrSH2j4sPLNcKaKmtEGPWpMb7nTv06pJmHzVWIy1NMYPR8+HAbPOL6qhmpWvYHU1
NVUWtKF3LRkPV3qKuyIeGF4JWeppU2Qkn/5z0AAAA5bw4m5csmD9Lr9AY8PTxclH
IMHeYjjYeDLhBHWiIxknCOHkPCVKpeZJ74Fcb7ld17HZUuBQ1k5HRX+6bZ9hdsGR
pjVDwwAICeoi+oM1uFCiz8ph7tPgcSsYvM0nosrpxqpgCvhPvYrprB4PTxavf9MQ
h7j7GfHyfXvMXwBGsptt29BkiwbFt3j59y3ZYxh/YM2IeqWlhUmuvhQW5JeMBYcX
dcRPJMi+/TfQnKynhSnHnj4Ymlj5RViR2KwF/5XeVSnTej59fo5AlP/aztlXbZ1+
X/E7clmGLUp6OA5LcXNjyHDRYiIL+oi15qVuAJptC4RwtETZqdsE2fpsR6GKzSdE
+asqkIvySPzK/1y4dyjqqZGrj3ZuektMHq7zEZvgtWvbdlnCf4p03/DQdkuduhtQ
MX8nxUSdRZ+hFMwnHnbTr5GzRQMlIsGvlyWRmncE2ZjgxJ/LN5+AcmCpGmvo5Onl
4dtM+4eDaDHLiifUk3gmA3Uh05v+0/NAwaElQznhDiDwz/NyXBzSzzdFZqKhYnwA
/hpsHnFZsp17vNV4hA8CDJbIgCA90g0QDcGkMSc/nBnA+yYDq17OAW3qI3qMqSEx
qFcmwbyeZjmL1NNQ8ubJ4RmmyBr9i5ZQjQv9H7dkDucLpd4LJT4XWHSLzxcWjXZa
N28J7X0gjvZie0qNxcrFbuVESZo6Svc7XEO/tXPXdQbJ/rNaxrI5SWE8esYAoqnC
C+tFOXNDs9WGbWOQ8xDgN+ewjEYAT9sSC8lOJ7H47Cti1z/cqq8iVZk+O5RhSwHt
nHelMQ7k6Zu3OojWpSNy9y3ADSmiBbauN/uYO8DsNmTHQiUm9S+zWdP5DKwQo3Qi
4CV0ndSx3kxw7Q6Ut4RzbGG7xRWZxLcsC2bOMS/Od3bJvt5wR/DEYyEvATjDvZMB
w2SVriHK8J4kQa+5GTu0TkfXwbEOAW/jI5rkGm8jWeATMewSrQiuwkh2EdHtYxem
GYTRTNDcdkU9CbyElfeRtFgtElg3t9j0ZuFsrTB4zl8idqdDT7FRERSD0PFhZmu/
cc/G5sbx/82mKoaN3ImzyRoOza39eaaK7pgBMh8BdgyocftsYDKPodIzJHv1kBMD
YDAI2y+vjjTIOjJOk69BRq5YCSjN2tkxi3IRcf/qeLgOJRK6a13I6v9WoiDTBnIl
JMewKXm+MCXaduUDNGZ9JqC9937lT/xtzyr16UaiAuvC5cracCZsH9InYCwTCycD
mvmooA8yFjvjGNpT3k0+L8cQ8TSzcjSCA3/gGsRaeNFzQQOwe7JMeCGRh1CPC/X1
XxzlHZqEOVM4GGHlJ7LOFT8c1cLuPv7+dfwxa1ZIhlkMlzI6w63wAo/UJaGizV7O
zF0X0La0kKEKenxAwpKGx4oMgWwAz0kukcOGeH/octCSaQ9lrELbK9RlFmnvcFfU
Q0i90Z42Clq8tK6Xjje40P8Ebd59c6U+KRLAcqE/iPbnafywfCkb5IckeI9sd8wF
KKwjAR0q2IhMTgPKdX4wGNMsGM/YEyb/pFqtUXhoUPVBo9sgQYGQcO29ml2T/IW+
hlR7FR4uDNMTfVbCcToSg3fSkl/p+LCdceTFGBGX5xajCixd7N1+iKuAgg+aeB1a
L74YgskTMTvU0aK8oIwKhcEjiPusk7xsigGiEnIY1uUEzeNc9tdQBmm6KsrJCdqd
jdWrsuGwdsilOZsDWSfT5848XbUGBs4tIvq0Zxruewr4tBK0AFBLcq2vXdSk2s+x
NsTyEqLnm1lMrANZzE3A/kRTbCCTWslsTch711kjw09twVMnaog1iAoZJeQJ3SHP
3uS97QP6m/IyDcLykapS9/K2BYUsxaRn806Pwqta+9P8miQfAhafXF6jpvItsp5Q
g9YlPa1hg9zuQSbaW/khwEOesJicz+hSnVwwcWbKhcsBvVZ6GUd4DMDOfFl0e/y9
OnZ9Y3Lk+7WXPkoYAozhAFqEPu+FJrKYdM7pn8kMZKZh8dTvcoZ+VYIYI3lUUr1I
hW4h/f+A9qhGHwkOln4PS/1L8PZmcEL3yDtZSlOqWZgAy3QuMUvtSwos3q0WKAxR
UvoKsYHLZj+/gJcy3fJMPm2ZQvrHGGbbh6YAAvp9Tt2ZOUJOWhNV3ABGv2schvpp
sHKJ8jS4GtXIKrpvHvBWR2Nxydw1HoangCm03D1x5ejMBArmQ1hHvrkOP7edAH6q
a6Q8gKK2fIoA8bTzqqGoP7CxV7O5rAF3T5qNSKkffSOZFQOVE7MwrkthFBusRIj9
WAXizfwco0aCJjBDcgtMEDj2StrposQ2NaKLKfjj6ZCRIxXrAuaSmtnn65uYHR9R
0lLs5thboWireXXR5S6tZ07UL378RNYT1q/bwxe5As5NQ5mXpz9Z8+fYp9O9+03l
MCwI9GopG22Kwga+R46borzZ1VmAl8cpkjvVuhk0KZvoYoWrXb7hOwvEGMQEIR0R
rEqbJzjXWPlgl7h+hvNu4JgbYIEX5M4wrGdxQN/+1GqtjxZgzfuDPKiTWOtd0+Q8
ncxyKXMJmCHfwwTObCBjzt0Px0w24ujgbbyre+zaplVKHQT9ct9J1qlUuo1Rinnu
Aa1xFERv5Ce0p973dHSMTdyMegKcUdBRXxA2QFv6mQUA3ZjRolqdP2XcL76M0E5e
aDhSEchxRT5cRiKqCU+NeAhS2WUFs3uS6uGsEBTeM79B+fHYY63JdqnHHPaq9Upt
2F4nR/wnxOKDnyIiqZpsTcTnJs4Y8PGvVaROSaQnIJtQRlUAzQP1zLsOoYGtjU9q
lh4MrltpKfDjhv8x0UOJZlMdxdFdBQo4oXnXwhPgJAo5NqHSrTp83ZODLNrY+L6f
S6Y+78ix9udd2hDIhE0n2HO/QMuVUQiu0bv7pd5cKW7o9OEghzBUkL1ZdNV15Ogu
/g+v5BhSpVLoavxqldgr/VF4Bt2+lmsaWGTnKVZPM+WgjW1cXnKD/YKK0LSxqFea
6ZC+3mVXfuon3GQSPqYkPnPr/AVc4yE69UoYc27WDAwgNi8zxMxbteK3XE34ytyZ
/S7uTIpWJrg6ICnqSCegJkxX2ADPzE+moXXL0ozKXfvT18EuCpTc9RxCVIXXL0R+
t9epooF9jPkMSZ3iixer7OO4txDQYGYdJySu5jHPboyO2OQaTGqR/3QYboQZbP+v
jt3eH4SBycvz7XZSFtQ2y5UnXO9ol+5DlGlaJmnnCZtH9PVVTHYWmYE+p4aHvvnD
eGmj4MRoaTvw8sh1Ex7als1PPhfJ82YWm91V/TQX6Z2HVWat7TGhYrb/fPFr7o4e
aSu1MA39APn3y48LfVVDEeJiVANVagxpyO096mfuteBVHigflP2vHadAMWyQF3nu
noSEYaDwW8uEp99NrckgdP8lpptomq9FDw0iqJ8xpn95dKtgBSmdLDcba4Y9ozO5
edZzGdQe9wwkj95R5Vyu+bxklsLHzknE/WvydlwtfjBAg5XodONep5glFXP7Nh/5
hQ6d4c0EhrGNGQK3C+RGnjLyUSbxpnITM/B5YOlEF+7VuAuHpB6Bv/GR5TShwzp0
KEetnQmNq7FTXsWaj5zAoQF37hhqDWKKvbiv0d7d8+a6o8VGr9B1QF6WWMBjsGXr
ZiDnHImSzJBmLaAEYjjN6uFQ3WJeHWYs3kZq5bf6O4MpjpbbRUMqPVJhtDyFppcX
OcVxOwQDsAShOO0guSPwCzisFydu5F5luYiUBn5L5ZZqQAA4ScU7M3fC2EpQQNFx
l/ZWrQq1AYNoc6DHMTlTEOGWlF+AufQR9gTfcFNIuX+5Fz+76JG5GH74XSWHWrz7
aUVa4A/cDG0sNnQgkk/wchtBbsEUaO5WXptJvVIx/RZgu3nzE881OtXFgCPGbhFk
HT/6HNhPqZ+eN92v3OhWzTA2jqUcC+X/hJwiffnEUAYAayhpHiUYME2/r1jvfLXX
Ufxgk00HeVcxFz6BMkuiaaDVGUuGIPwXbBOI3fy9INbl150K+mhqJNqNsk1dhL8s
kKzfaq1RlY/00SRMoNdfYu+HQ096niDiTTEYhcjKqYaN59VuowIpQoA9wIemMRSU
uZ6WGNHIPikOrYAlhOZZl4yXFnes8R27KmA+HGn+PHU2o0a9vs/YVgHQtViRhYcn
Lzu5RnQHa349NjhklBJr80S+GDBnwwYQCinIEG4AVGLppbBhFm32zViE47RUTxDt
99zvGt2JmGq+OAYmhXTeyaKCqDnDfeHPX96Z30mM6pAHLztJpG2K3ekLbhHQNOm8
RonBMiLuk9/6LOw1lzD35/PnjOYiM2fOceA0Tr4pCDzNJGfFY/fQTenJazKxYkcO
NJy4XFbfNbhTrCDDiShFikS1DwCRfxmoGcFtYNr/787Ke5/UydUUOHScSYzTjhMK
mc0CJvCEGOOUA18GyZ4svEPfhzZBKoGmy/QOPyCsGo6bosLGL6Rnkq58Cy1NHsVF
sGZBg77LLjp/nwedMiKgfDZ+ez0Exe5oFcdz8CpdIgZWHGt4HSn3QvYxziT2Rf+P
1wBMB7XLoOdBy6iNIEQIVI7X15b2vEgVab89mtrpf4WvFqtKAKZ39cbV0pkwkbNB
0oyFJCpzdRdU0/rtFfDiU2esO5sqBISgmlft6/5txBk+oa0NMxg3DZMXYJEail4a
MyFvXBysV+Ce3P+/A3cODU1NfbcrP3oSeLD9V3Cpn1Zo6S+mwr2cKOvtMSbLPKAL
O3Lm0T2k7T6Qjt9cDfzU0Oach6eFJjWNgprcqBSmR/oa0LjbirEhG2B6l3ywZOOm
/u7sOBvaaQBuCU2/QvXZeYA0ojyzwyLkktjzBJ6w1AzzNuj2PxI1uy6jF3aHTnvA
dfFiiJ4m74RiK/+9h9qLRRm7yzBh728Y3NvNzO2384W5VqUzjhaZ7tvI4n5Ic2St
EDhjK3S3pcZsWLzUk3UemfkAPMUMPDuCN5sZ7xyXglni2YgreFjGWXCpu+R9y4wt
SFWyW/ZBzWtFVHFtVnWNZokNlFBS7gmVRf4SURYei/A7RcGvbzaYsC3JlGo3b21f
1Q2/pxTqOWxekGuXBOcstxbSLcGmkFUPwBiLQPZ0y0iYP/yEPtLl5XHxKXY6q0/7
esMGLcsBa6FhHbGKbOWWMXCS4U4InZteSayxaetxwsMUZpYUpOXM/0X2k4b86Nxn
tNXM0CrlE+KaSlvM/yXcGOm85JDPmxbA+e/36hkYncF/JXTEzhEN9UIs/9i5nbC+
LeKl/z/ikKAm9YKRLS9AvOPXNx23KQkInP9WSIr+AS/1sdB/HqsnCYrxQFuL5M7L
ypPYVWy+rU+gQiDYGIXOfNSxzMyIcohZwTHX2uvVrip28OwxBBNrBLy6JZu+xmEN
oZtn/0LW9W7v0DjfyJ3HlvIYp3w26QvSqQcWsDOmZWGNjjcUlDSxMHBCqMDUXi0J
Peavx1wsFTXa4yLt9J2m03czvFojcrFEWsMSfHh3XH/xJHouhQke/4Mvl9aK6MOu
s6zSFGVHpAgkBy/rWBKTyquQc8OP3SiHGubF24i9Ut120vuzvTaiZGoqo3GNXxR5
z4Zio5/Cjw3EBR92k/BT3qCveClvZUxwHQoNt861WMs2YMqb/ERUyY+PI4Ben3lR
6GIHbxtaF08SXhmtN3WSeDIQ9fIDgskI9JwiGxkvdI2jRpnJ1Lmk+5qNx36U8ERB
5YD734p5IIk1TYvrZyCvCbrkBAuWdot54ic0Wz++1vPG03/FWo9Js3WF9fB4Pf0i
Z9Hw/P772TTfKHG8eTU+B8wJhZSwzsLntzKPQEYLZg8/jsXPdv4RLPjGtoEKsIX3
Z+NBvIVuyBlqh8O0DqODf1mQpOT0SAwoVOoYQS0r4yJ2fiS75mXSfFySmCBpNOzY
rdG8uayY5Gy1yft2Pb6CTT97dn7pEbWeGtESukgRM6fbh4Seb3mAtyaVgq5BLoHN
AoW8L9FHCPNiqRHKAXOMUtmPyzx1TIjURmN760xz9U1KB0gR3A4fiykdHF5DQQ0W
Itbg22twWU0qp4nzFM/AQDvV9xF57IUTF6bsWDdQyGHildk3Pf3zv46MWgNVX33H
6bMMf041qGH9DQVdccLXJY3Pf1N255HpPACsRTyxNHkGgf3BQ5Z1fwkWdb7lYWil
x3XuMmnMkPsdKgfiU3imz4qjivceuIv508NbbCCatfjp33f4OzIr/W4tKcjbNVq0
DWQ9oPWsPts3gzZA+VbbPEglCHfkd6VUmI5Ksd+uCOdgx99A4islqrYV4oEHgODL
3zx1arUcBnRaRumuGQGJ3M0MX9ApQusf+JPb5Ri6jhfkjA3HVAFVVa5a55bCS27a
Yeu1otw9zP0N7OAt7SjxHfsGOjzob3ai6O0yL1FPBfe2TWfsKE+s05RztT8jgnrc
+fbNO8VqmjnZ6oUfyT/C2KY/57xv02cqpcYLwXSbIZR1f6RClgPVQhiWIK3k9lgp
Z4HyJf//rQlo5yiWfeOegsKS+T9bNQx3kaXu2zmH92ydBS8jihwHs6yengnn7Lo3
+Ogi1ZxbBbuMi3OtSf5ZJj4gnGtnM5TCewmwjpRYs/iMYG+y1ha4oS4rrxwQaY3o
jks10Xz1RBgW1wnwxdLA4kzkstXW9QId5zXbRjBwymc7U3iaBHsyoz11Ynq2Iszz
3LWdEBhfdXZfZTfmWvd06+h6WhQ5srJwUp/pxqmsHjHDwD/k+Hw5ljiymdrfYyXq
Lrrr2XDpoYB7Cve7t3vaDgnxVjeIuEB7a7zxRDBMKSDEMWr+8N/FczXRWL2bYSpq
KYJOcrrCuAHNiYoIxgdrgNuE2jmfxFzG76l5IoFy/R8MDNpfk3cJssgcm5STQ28f
5fYyZxQAoxwvimS9Zqf2rDtANhzxxKwL94l+Se72esYxu33fAsSH+sAT3q6LxHkt
7IkiLd/VJI4ydI+tnFc9JXYy2z7EOSVgvXzFvPF9yB/S735vGQRyY36ObipjEUOK
z7Q2S9+hhZXwU1nbGk3oFtip0lX9PBKugyshthaKq4/vBDQ7fOAK0olQ7bYQP75+
jNIew6JtSo0u+Hxi/UlGPxR8VxKc+D/Fe5X1a8Ou8X6hMX+2V+LqoOxaVAwMNcym
YpLHjxEGDkWg0HE+nUO1/OY+Ouy7Wk3L+6i6kKFtqhI8RY5XMqBucpljw08fCNzl
QsXaSjJ5/e5HyVrW1JCvMJSiUgRnOCgHz1BX15CNzC/H59ElWpnMr0VCxNpdFQMe
v0aNBUitrPpjtA/Gi9wa6kodb1JQ/PjyOB3601KdPIErPSkllaGlq5Zziz4el6W9
242H2jjH9cCRie5Kc0LbNCOixmH63fH2fQjGmAOGvW4kKOOd9uqlW4PIPsVn6fDd
hLwUgJCNU0AuwXhuiXn9HLitVa3x+Q4YeiZXuj2Q/+qx4rxBJJKvdkVG6gV630+S
r/H30E4wxu8NTQVNgnDbpapZfbSfbKDjIZ7WCSDnfHw64ytEIZZ2VC44boBPL8go
dQNlEjHREMtF+mJhrxX5fs6Jzz8xGI535uqePm/WucbltOSrhWyG3ymAu0ihSlFM
LppjuDd7/MZCdND3lwwPStc3gbkDZkTl2kqDx+KbNTac8QaJ58fD8j37O0tUnWoQ
opkp5JA4cQWMxYXaRcqqW0kdWVMPpTpNjBMLkXkaZxF9mwrUmHVvmmb/kZHN1nJs
uJ0qqoApNeSQ+l01fpGuK8WK0JGlnpHcWZeRm8/IknIKpisScfnBG2c5u9WFeG/n
vF0RI7Hile6hiXr+dQDErCzjagQLpu3U4IaE4rQQe+VJu8V2pTPg6hVUhdFVAkCw
0cJhqPHDnjHEkAsjrPgPAQXNVG9dx1vORn3g3pTj7V+6uxEpOaPMPT2IlkxhQKMR
bYx3MgKPFR5eD5gVtTIIoVHLq02+MdciNIllS7R63iviDeiBvJpDjbDbtJsNtVOE
hNQS9ydF6jTrjzadPOcQAXMZezEawMn9C4N4+H+M+8pY7aDwHjjsQvXUf4rKN8q+
3KgHNoExRSpV5+xqH99EJ1RoHPcbTt5PqYByePQm6qt8pD6HpS/ge7So9k9paD4U
RUe5rSbTMbOdyYtk2nLHr0fzTM5Qum0ZiBPCA1/L646f3lfNng0d25RNFxgdLcvR
sBZCbDywhYohqxMDj4ZvzasjdjffkvTZ1vQpa2UyywII01flIDEYNGT+j4vVW2ET
NtKOeFkSZsB+jwCMa4vHGgcdVnfAnhpThlRTNSGnHoVQDjW0GMkm5r6W8Z78bh0j
1B5k9cBVRmFcNP5OHyjbc9roBxcMBF+emgRRHb7gd3xJamQP4DM8QEBnUeDZZLu0
Cuk0/OWCfFTLFoVM/vI71mW5iCgubnMUb8uK81xxQTR9M57iYsh0Ccvj44sUrG9H
HxAtwZSWmBfv99lWlNy3Uv5PxvvvKcO1bXNR0rg0qgZK2D2xlZoL1RbX2rhLvh7S
bjroqIFE1xFbCi9hLweEEVvXVLZ8c2njlvKzYoZfOzv6g8sI7AM5WQqzopzPIhTH
xkWN+t/48DqZCr9hzxofwVa7I4fG9PydDZvPCdPwH5GMRyptXr9H0aVxFUCvmc1k
zES76vwYkl7DWT/9yRvJ2en/yXo3Q39Kuw5gnklw0F2+MClHGVmPvwQoASkH8PTw
pIgjYKWS/3lIMlzh2pSV/SUTrPL3eFkckAsiK6tpsXvzI5gmvxDi+9Hm8kmNkX5F
PTTqvDcSfXi03A1ycvETY7DlRwyqds6V7M1lO5yn7fMcCqkX2qKw8JTKzmx+JQ3s
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
C5TSdE0RFlbasCxbTiBueiCLiMseR/yGhZ6aMlqqm5SnlLfBbQHP//n3z1pMcK0T
LVFV58NcPoeCec5eKjZ2plvcYBu48ph8bkNuvcJ+5AlSZPdfRq5bWZheDeruJcIB
qVL1yvHKs5TrTL88Yb7PWzzEpP4IxBj5iZqENmfcPfk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 232935    )
AHSY50gtrlyNRQFIBQh6e1F+mj3wS7Dwcbt/7hOZ7dDFlFGN5LBT0pcJ+xVmZuY6
v1LqkfpMqHre4M5jtgRz/o/Bl5bSXYMPmigy/lgHKdCGUqlqYfjvc9nY9Ibmr6yV
eNd130IK1wms4ITdv07aSPVEPksstJnoXI4TN2RyJskTsHanWaFt7HCW9fl5Ut53
eq9ixLgThTZK+c6luiETglbzjrhXgBcGeTrqWJo/KX7n5CkL00M0e0TKFg6SBcVe
GhYAZ+uD8p2BVkZCVWZsURhbC96dQPI7VHqRSzhDq8MZ4pTveUn7U6LvGzkwBugE
`pragma protect end_protected          
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
c1bu596v73xLF+v1CBc8G4EPPIqW9+h1tykFoHY0CF8+yDdKAquUzqbrkQ3/bMh6
jzaqHmDtauqopMztSMRwSQyWS4a+d+YeWK4zhI6kvzrfvbcM4Q75hjPnUpqR45yx
4QRt1ruM12LhsA5RLnut8t8wLXGoH03ySKtbE1/XP8c=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 236213    )
WL1d4Sl0OmVjx33x/DyYyCmOu7E/AEFR7WFnkMYVpC45ASDVxZc7Orz+tAQfeQpN
bgADo0VKx1a4fDxDnX/UB99DUxczTDKYwFSIbFPA+Q2qGqJ1wGMn6Y3tzPM3SXSp
JC/3SCghdh9HsP1N8267HCHzsrzTS2F5CKw8bA7rFBZdOnfvhSwAf410C5YHhUaK
MxuirZdNHPHZjAmSP4/v5yvLEjwXDwh8ZzQ9gbuTGLKwEDahf7rCjIhSmhxprmd0
UOeBjAU9K+Ps0to8qrDRg4/Hr8vvCG8qIlrk+YfBYAQJG6gcJGStRJ1S4l+Fyii7
quwgJxRZwoG4QJnrzfXUX8ozuE/4G2yhOUKkdTB1u8kx8mFmE51j9NUzJn0kDAbl
KWFl3Ifwdj/QsbgJabrURXLShdvs6j9RVVkkFX4ELAQe1gCzh+so9UAhRwSjI3P0
Qwcr9Fw5BR1glzTnOK/cvxuCE8HDh/CweZZHFol/U0ET1pNTUNVdvvm79ficK5Z0
LrzX3TvJjtB1Qt1ut83mfZ/tokBmzIYYWRY8j9soMUJAPlepBjUg0167+IG6jhPD
nYK7Xkl6xKaFv+IC3+ZgrAG+61sUCTtpKxEA/YPjtlayhvAf6xTJCmS/vmW46Vz2
20Nof+fCZoLXMDG1obl49oq2oVgHICJS8PBFvipCeUXoMxKRlK4//VR6bjm97RPf
MqDdEGttp45dvF+hSi/UNTZWVx6uWHr5IFKDyiCzTaivXizZmJF+zBqPlNa2l6A4
4wfsHAkbOpt+ETzVmRJ0zab5OTWUjMcG2ivtpj/yjNTwAkxlPai0UYwxDBe9n/4f
Y/1kIvr7zLPocTvSdnJo51yV+/JoHd7JlEMk4ETfEwS+JNhaim4J9HeDWwl5uqya
Nm9sLGaJ0N0HIvk39zeGoxJGl1KstDBmUY7Awk9gl4uI4meDKflgy/bHQUuQrvAm
vGJ9pV2/35oE7BRiNqkixyGP3Oq4clngaTS+GcbUm6zWRTxFT3qrbc7CFhnk3fpw
TEubJ1imjj9dKXvoKmLJWRg9tf5+6ZmaGt28TeeFVVbHyZ08Xq8C8epMYI8g/5lT
EbgwE0/7J5FaNQ8ds+oJ24tePw4Vnvf/Dq37EmhTBYvbDm5080un5evS6qORh4jx
+mZLmvMy0n5uRAccBbqdP2vWZju2SCLK1esSVYMrzPbL1ejbz0SKpMuEwYEgK4Wu
04+DFXSeGDjDb0CYQgph3h/Byk1SS2tDhQdd+FJ4/K9vFqoSUCD6VA/6boK+NMdL
+Dzpnu0E1hlpMs05OrUie3DUO5EEZFnxkayWMyA5sqoQI8B/aP6tsOjybbqAqeqZ
3s6UrhGhnvl/zGcC3rV7ZHYDeN+WdgzvHzqS7+FVjmDmY7EIyd4PT8nZhbYkiEFC
veVQD9SdBFoVQvQyVXaTRWIyRq5EJt3NEGp/TDTrW1P4Q7rHEPzEVngwtohgxVhz
DgRmlDmPSa0iodF8m49TAzeDe7Nai3Omar9/dOuzMsv7OVjDrvZIGBqXf4gDUryF
UPAag9+1+81x/5QFZSVStFgfPjykpWfZNypBFdUr8s0uTozo1PVLeW9+linHeFBd
ridPAZlq6h4UuII0RsqXZhi3qUnV4uaVJrkCMbWwpZwVET/Rrw/C/uUjlYxZ0zYZ
eA77g20BlS2gA82D+XhBNGuzy/qtvFdPZwUcvC9ao8PAEDJzaz7qhG1jIH28+CuC
uSSvSsDUS8bDzk8XoiajoW06+IVRBfYWoQD9L4AKqGHC9jJjCTW7NWwOVLkdb9R1
2AEvR3VB/8gfcerKzOFrcuU2toUf6JVHdCEDHydI1avxR22NCMY9nYEiagjKqlTa
Z6LzrZ+RM8VbKOdmqH/WmqlFpK/rIrVYuD2ehGjNX1Uc9jdtYCP1HbYOx9sZZJNg
oFUoozTm2bsR4C87WoF/O07utJCZwkSOINsIDSvEhboh8EDv587oXBZXLTFo/9Io
CsGBCCzdxlAgiYAlCvtojmBp3TKRNESQ1NbsvSDX4b3ohkT+l6JxPQ5nw88VRVCw
8rZaJChAJB6Lgk8DDl0LA4oDb40onU1XzpJviptsvpY32YFLq0+1HSR/gHvpSYQk
01mFHRwX92dBcYhqp4/7xDy2l4OLN1wYCOP5lYvzZnGXz0Ue+REpwLUUoI331OxZ
XCD2fPVdc53u1hMCBMw+sv/Nf/eiTx7woPadoPXOW6bQNZr8+Zk9pEcSaIWQLqBs
GE1MBE1Xpld6FUx2ywGfdpMOaKgxjxR4eyD7n+/F58ero+j49P5oFWPg8bkigyLZ
30O1SgTDZmlhzeua2TgWQuMLJGL03BMhBLgGwXE25t347Bg/D6kgUVDSyb1I4Y1A
+ba89j/GjLbKSPquDFaMwKQ9MArrK/Dcs17nFQQl9U6Rt5hMWRl531HPhFrCI4FF
TNk4olL6yljUFBvlsj+AnsxeTTJEL+QkEWBwcfpzxpDAzu2Q6kf2lSsO6XsvlUz/
fWJrDiCPpzVxerqb5C5jzNL3JEFHgiflTl+4k6NLJ04Jk940jH+wa4Vde4DJL/bS
GhKnpmhhJgvm0aG/Ng7oFJZO2KstFKXBVGXtBqKI9wqsJDZj/o63PArSPKxrpMgu
l2SgjYzxrW8Bji6c8jIGXKsh5fFlu8OLeP3EP1niKuEqyjDhTRXTfvDrGqa2IyzV
VLXEPmZDGrhGLwbeRl5X1970v5zirsvUwiJr74iMyPC/aD4RuJ43A9m4m21X2CWn
iWOjaRzeRyAdtwU5LS0wnV00Qf0RSvpZsf9v3Zn08zRhNx070DOT0cGZzAzmpebQ
TtfVsqbVKlTSo08Ql35+SvOkfbWJSUtoDRQ4XRWd89wg6z0Ba4q+00XiTeKZgHsY
m9UHsvxNPqdT2mM+QuHjupimNMXWJHyThO/CBpZuzwdXVDjF3DMKhyC9Jp3mGuuH
EC6P8kPrIZUgURUaITqJmLPLjhRIo2tn6HsH2X53DPW3m1es6rbGXuDwGojlGwFP
ww/NBIFPOI9wlK4+km05gi12m50hlnWCqlSEhJkBbXB7PiNQGlZ+a4RgJ2QS2xqs
RJF9UliXcwRO72hF/SOgG66gJayQz/j2h8nFWSOhxfTfCGBPXTg6lmEL9SK1lhYf
GwGzj7BNtAlvMZjGiVwfPsUakpiGvqR7vry/E1+bk37hqpyHH2fvgLUniR/XllKu
MMM54xpCo9wIxBa3BR3/P63SEx0eqEB4tlZN/1kFHv4utVu3HotZHmGvaR9Lm7S5
B8tv1Yp+/27sxvQwA8/Em8Jzu7gIts9fLNuE3AqkP5yoJGOK1gnt0lYxdhBCKj35
SmEzj3IivHExACXegNU5oRg4yUR5gD6KhPLZgxajBokIiefY6qyPhkpNReQQJHAe
0z9fXDjdY+lTflNJx8D/Tiwp4YBb/ZK96aOu9n56TsyMhKEQdcJNnrM+S/z8tPB8
0ouCbfHMXdOdkxpbA8vwidbzeH3i8OwS5qWddEG3i0B3KoPm97mzgYKplCAIffS3
6xPc9e4UOhKYXoLBeccN0b3OYvYrjl1H4dUuyLLc9vp3QAFkLUwCaMGlGXsUoEDQ
wIK7qvpad/ermZizvTe00X+BaCJYkD0wWm++59oozvzUY8e7431qsL2ZdQY7cZMv
O5EmZNVRjL9PGXfcJKVQwjuVuN6f76d+FYXFzV6MQG/hRZwX77ocrCuf/2Jo2DMc
jWACqvqStUBDvct1zK3H1ahAOXqhWB8JOpscsZZrX3PDYKaZAIjt3p/PeMcu6doP
lwW7IHgUpUwjBQACxgjq4hc0vg1ejQaG845vjtHDDEmxytsJsVnHMHjf4i/4wN1q
NBElvg6G+m+VaGEaEW7E7YZDTWo75Xz10Ai4/17YFhPK4Tn7kU+8NftZpkqK5lX2
uZQrDAQ3+MuG+7fM4bqZ+gMQQGqND9sd/bIjKVuzh8pFGyQW4Hg/YSFa++bfMaID
/ZpJG5Qcg6SrusLyq7E6icfHXlNXRrvlvA68EkxzMIFgdVPQu04MBHT3elWqxdb9
fNLSb0k7iHuzYN7xju2j9i9tdfF/JVtHVoAJ4NE2aIvHTl1N767h5+GRSqRDHP5b
B8dizy/HBqTq/SD9A7PaQAHCnX3I1tM4mpcHhbR7M7N+JEp1+tZxpyXEnaGM9loq
TwPewY3IVgG8/sv+C4jro6aY0dYzsvBluE17bu+E0bTJAyejiiUEnkyFzBF2CC6N
CAi/qJLhHkpiLsmscZ2WwwS4/BbnlOlt4SpWjCeOAdX99wd4HNYNFiiGRrJgKG7M
DCUG1MYWeWmvW09aS2FI3ohNYKkDOCsYxcypfM4Z8EC+dGsfDfySamo2aLSkWhEE
pT7egJNzFgNFeZP4K31rdg==
`pragma protect end_protected

// =============================================================================

`endif // GUARD_SVT_AHB_MASTER_ACTIVE_COMMON_SV

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Z6vHT+o2mzW/j6TYTwv6bOCmAyyDhy83esUM+RYUQrgE5v5aXrcXOzA4vyhzv85R
pfqw7zHxKeEwxYw+joVcvYxnyduRMq2suL8eUJcwC1W9kEYGD1dJC27o6UiPcuYT
RwKZ7m41ecJTCHjH6QldN/q8RO+nOxIY/TXFJ9Tot8U=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 236296    )
sA2iVhb6SX38GGz+LtD9daB1WvU7xlPgakp3E7raspnlHWfn3+ahOTPURgC/LHtN
fdQ7SlWCXujG9pa2I3N6rhgi7xPiKMduhQzG8mv/TVsXjz+Mupz+hNMOYHGhyhjt
`pragma protect end_protected
