
`ifndef GUARD_SVT_AXI_SYSTEM_MONITOR_VMM_SV
`define GUARD_SVT_AXI_SYSTEM_MONITOR_VMM_SV

typedef class svt_axi_system_monitor;
typedef class svt_axi_system_monitor_callback;
typedef class svt_axi_system_monitor_transaction_xml_callback;
// =============================================================================
/**
 * This class is a VMM Monitor that implements an AXI system_checker component.
 * The system monitor observes transactions across the ports of a 
 * single interconnect and performs checks between the transactions of 
 * these ports. It does not perform port level checks which are done by the 
 * checkers of each master/slave agent connected to a port. In ACE, the 
 * system monitor correlates coherent transactions and the corresponding 
 * snoop transactions to perform checks. The checks in the system monitor 
 * are geared towards checking the proper working of an interconnect DUT. 
 * The current version of the system monitor requires that cache line sizes 
 * (svt_axi_port_configuration::cache_line_size) of the various master ports are the same.
 */

class svt_axi_system_monitor extends svt_xactor;

  //`uvm_register_cb(svt_axi_system_monitor, svt_axi_system_monitor_callback)
  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  /**
   * Channel through which checker gets transactions initiated from master to IC
   */
  svt_axi_transaction_channel mstr_to_ic_xact_chan;

  /**
   * Channel through which checker gets transactions initiated from master to IC
   * These transactions are sampled from the scheduler's output of the interconnect.
   */
  svt_axi_transaction_channel mstr_to_ic_xact_scheduler_chan;

  /**
   * Channel through which checker gets transactions initiated from IC to slave 
   */
  svt_axi_transaction_channel ic_to_slave_xact_chan;

  /**
   * Channel through which checker gets snoop transactions initiated by interconnect 
   */
  svt_axi_snoop_transaction_channel snoop_xact_chan;


  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  /** Common features of AXI system_checker components */
  protected svt_axi_system_monitor_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_axi_system_configuration cfg_snapshot;


  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_axi_system_configuration cfg;

  /** A semaphore that helps to determine if add_to_active is currently blocked */ 
  local semaphore add_to_active_sema = new(1);
  
  /** Writer used to generate XML output for PA support. */
  local svt_xml_writer xml_writer = null;

  /** Callback that implements transaction XML generation. */
  local svt_axi_system_monitor_transaction_xml_callback system_xml_gen_cb;

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new(svt_axi_system_configuration cfg,
                      svt_axi_transaction_channel mstr_to_ic_xact_chan,
                      svt_axi_transaction_channel ic_to_slave_xact_chan,
                      svt_axi_snoop_transaction_channel snoop_xact_chan,
                      vmm_object parent = null);


  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /**
   * VMM Run Flow: obtain a handle to the configuration through VMM Opts and
   *               build sub-component.
   */
  extern function void build_ph();

  
  // ---------------------------------------------------------------------------
  /**
   * VMM Run Flow: Connect the channels
   */
  extern function void connect_ph();

  extern virtual protected task main();
  
  extern virtual task shutdown_ph();

  /** Reports transactions monitored */
  extern virtual function void report_ph();

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

/** @cond PRIVATE */
  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** 
   * Method that manages transactions initiated by master.
   */
  extern protected task consume_xact_from_master_to_ic();

  // ---------------------------------------------------------------------------
  /** 
   * Method that manages transactions initiated by master.
   * These are sampled from the interconnect's scheduler output
   */
  extern protected task consume_xact_from_master_to_ic_from_ic_scheduler();

  // ---------------------------------------------------------------------------
  /** 
   * Method that manages transactions initiated by interconnect to slave.
   */
  extern protected task consume_xact_from_ic_to_slave();

  // ---------------------------------------------------------------------------
  /** 
   * Method that manages snoop transactions initiated by interconnect.
   */
  extern protected task consume_snoop_xact();

  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void pre_process_xact(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>pre_process_xact</i> callback using the
   * `vmm_callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task pre_process_xact_cb_exec(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void pre_process_slave_xact(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>pre_process_slave_xact</i> callback using the
   * `vmm_callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task pre_process_slave_xact_cb_exec(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void pre_process_snoop_xact(svt_axi_snoop_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>pre_process_snoop_xact</i> callback using the
   * `vmm_callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task pre_process_snoop_xact_cb_exec(svt_axi_snoop_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_axi_system_monitor_common common);
  // ---------------------------------------------------------------------------
  /** Sets up exclusive access monitors */
  extern virtual function void set_exclusive_access_monitors();


/** @endcond */
    //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------
  /** @cond PRIVATE */
  /** 
    * Called when a new transaction initiated by a master is observed on the port 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_master_transaction_received(svt_axi_transaction xact);

  /** 
    * Called when a new snoop transaction initiated by an interconnect is observed on the port 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_snoop_transaction_received(svt_axi_snoop_transaction xact);

  /** 
    * Called when a new transaction initiated by an interconnect to a slave is observed on the port 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_slave_transaction_received(svt_axi_transaction xact);

 /** 
    * Called to override the expected snoop addresses in system transaction.
    * @param sys_xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void snoop_transaction_user_addr(svt_axi_system_transaction sys_xact);
  
  /** 
    * Called when a new transaction initiated by a master is observed on the system 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_system_transaction_started(svt_axi_system_transaction sys_xact, svt_axi_transaction xact);

  /** 
    * Called whenever system monitor tries to associate a master and slave transaction.
    * @param slave_xact A reference to the data descriptor object of interest.
    * @param drop_association Indicates whether the xact should participate in transaction association or not.
    */
  extern virtual protected function void pre_master_slave_association(svt_axi_transaction slave_xact, output bit drop_association );
  
  /** 
    * Called before system monitor prints all system transactions,
    * using this callback user can remove the unmatched slave transactions present in
    * the sys_xact_assoc_queue.
    * @param sys_xact A reference to the data descriptor object of interest.
    * @param print_xact Indicates whether sys_xact can be printed are not.
    */
  extern virtual protected function void pre_unmapped_xact_summary_report(svt_axi_system_transaction sys_xact,output bit print_xact);

  /** 
    * Called before the system monitor associates snoop transactions to
    * a coherent transaction 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
  extern virtual protected function void pre_coherent_and_snoop_transaction_association(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact);

    /**
    * Called whenever system monitor needs to match the type of snoop transaction to coherent transaction. 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    * @param snoop_xact A reference to the snoop transaction which is being evaluated to associate with coherent_xact.
    * @param is_coherent_to_snoop_type_match Indicates if the type of the snoop transaction corresponds to that of the coherent transaction. This variable has a default value based on the following:
    * If set_snoop_type_for_coherent_transaction has been called on sys_xact, then the default value is sys_xact.dynamic_snoop_type
    * If set_snoop_type_for_coherent_transaction has not been called on
    * sys_xact, then the default value is based on the static mapping provided
    * through SVT_AXI_RECOMMENDED_SNOOP_XACT (if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * set) or SVT_AXI_LEGAL_SNOOP_MAPPING(if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * not set)
    */
  extern virtual function void get_dynamic_coherent_to_snoop_xact_type_match(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact,svt_axi_snoop_transaction snoop_xact,ref bit is_coherent_to_snoop_type_match);

  /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param snoop_xacts  A queue of all associated snoop transactions
    */
  extern virtual protected function void post_coherent_and_snoop_transaction_association(svt_axi_transaction coherent_xact,svt_axi_snoop_transaction snoop_xacts[$]);

  /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
  extern virtual protected function void post_system_xact_association_with_snoop(svt_axi_system_transaction sys_xact);

  /** 
    * Called to override the value of is_register_addr_space in system transaction before it is being used in
    * system monitor 
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
   extern virtual protected function void override_slave_routing_info(svt_axi_system_transaction sys_xact);

 /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check
   * 
   * @param check A reference to the check that will be executed
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual protected function void pre_check_execute(svt_err_check_stats check,svt_axi_transaction xact,ref bit execute_check);

 /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check.
   * 
   * @param check A reference to the check that will be executed
   *
   * @param sys_xact A reference to the system transaction object of interest.
   * 
   * @param slave_xact A reference to the slave transaction object of interest, if applicable
   *
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual protected function void pre_system_check_execute(svt_err_check_stats check,svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact,ref bit execute_check);


   /**
   * Called after the system monitor detects that a write transaction
   * initiated by the interconnect corresponds to a write of dirty data returned
   * by a snoop transaction
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param sys_xact A reference to the system transaction descriptor object of interest.
   * @param slave_xact A reference to the slave transaction descriptor object which was detected as a dirty data write.
   */
  extern virtual protected function void interconnect_generated_dirty_data_write_detected(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

 /**
   * Called after the system monitor correlates all the bytes of a master
   * transaction to corresponding slave transactions
   * @param sys_xact A reference to the system transaction descriptor object of intereset
   */
  extern virtual protected function void master_xact_fully_associated_to_slave_xacts(svt_axi_system_transaction sys_xact);

 /**
   * Called before the system monitor calculates the slave address using svt_axi_system_configuration::get_dest_global_addr_from_master_addr()
   * and svt_axi_system_configuration::get_dest_slave_addr_from_global_addr() methods of system configuration class where master transaction address
   * is needed. <br>
   * In some cases the attributes of master transaction are required to calculate the slave address. 
   * So this callback can be used to assign this xact to xact present in the system configuaration. <br>
   * @param xact A reference to the axi transaction descriptor object of intereset.
   */
  extern virtual function void pre_routing_calculations(svt_axi_transaction xact);

 /**
   * Called before the system monitor adds a transaction to the queue.  The
   * user has the option to indicate that the original transaction must be
   * dropped and split into multiple transactions by setting
   * split_original_xact. Transactions are split at the boundary specified in
   * svt_axi_port_configuration::byte_boundary_for_master_xact_split
   * @param xact A reference to the axi transaction descriptor object of intereset.
   * @param split_original_xact Indicates if the original transaction must be split into multiple transactions before adding to queue
   */
  extern virtual function void pre_add_to_input_xact_queue(svt_axi_transaction xact, ref bit split_original_xact);

  /**
   * Called after the system monitor splits a master transaction. The transaction
   * is split based on the input received through pre_add_to_input_xact_queue_cb_exec callback. 
   * Once split, the user can modify the split transactions through this callback
   * @param xact A reference to the axi transaction descriptor object of intereset.
   * @param split_xacts Queue of split transactions 
   */
  extern virtual function void post_xact_split(svt_axi_transaction xact, svt_axi_transaction split_xacts[$]);
  
  /**
    * Called after a transaction initiated by a master is received by
    * the system monitor 
    * This method issues the <i>new_master_transaction_received</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_master_transaction_received_cb_exec(svt_axi_transaction xact);

  /**
    * Called after a snoop transaction initiated by an interconnect is received by
    * the system monitor 
    * This method issues the <i>new_snoop_transaction_received</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_snoop_transaction_received_cb_exec(svt_axi_snoop_transaction xact);

  /**
    * Called to override the expected snoop addresses in system transaction.
    * This method issues the <i>snoop_transaction_user_addr</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    * @param sys_xact A reference to the data descriptor object of interest.
    *
    */
    extern virtual task snoop_transaction_user_addr_cb_exec(svt_axi_system_transaction sys_xact);

  /**
    * Called after a transaction initiated by an interconnect to slave is received by
    * the system monitor 
    * This method issues the <i>new_slave_transaction_received</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_slave_transaction_received_cb_exec(svt_axi_transaction xact);
  
  /**
    * Called after a transaction initiated by an master is received by
    * the system monitor 
    * This method issues the <i>new_system_transaction_started</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_system_transaction_started_cb_exec(svt_axi_system_transaction sys_xact, svt_axi_transaction xact);

  /**
    * Called before a transaction is associated to the master transaction by the system monitor
    * This method issues the <i>pre_master_slave_association</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param slave_xact A reference to the data descriptor object of interest.
    * @param drop_association If 0, the transaction can be associated to master transaction. If 1 transaction should not participate in association.
    */  
  extern virtual task pre_master_slave_association_cb_exec(svt_axi_transaction slave_xact, output bit drop_association );
 
  /**
    * Called before method print_unmapped_xact_summary in system monitor
    * This method issues the <i>pre_unmapped_xact_summary_report</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param sys_xact A reference to the data descriptor object of interest.
    * @param print_xact if 1, sys_xact will be printed. If 0, sys_xact will not be printed considering that transaction is not matched
    */  
  extern virtual function void pre_unmapped_xact_summary_report_cb_exec(svt_axi_system_transaction sys_xact,output bit print_xact); 
  
  /** 
    * Called before the system monitor associates snoop transactions to
    * a coherent transaction 
    * This method issues the <i>pre_coherent_and_snoop_transaction_association</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */

  extern virtual task pre_coherent_and_snoop_transaction_association_cb_exec(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact);

    /**
    * Called whenever system monitor needs to match the type of snoop transaction to coherent transaction. 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    * @param snoop_xact A reference to the snoop transaction which is being evaluated to associate with coherent_xact.
    * @param is_coherent_to_snoop_type_match Indicates if the type of the snoop transaction corresponds to that of the coherent transaction. This variable has a default value based on the following:
    * If set_snoop_type_for_coherent_transaction has been called on sys_xact, then the default value is sys_xact.dynamic_snoop_type
    * If set_snoop_type_for_coherent_transaction has not been called on
    * sys_xact, then the default value is based on the static mapping provided
    * through SVT_AXI_RECOMMENDED_SNOOP_XACT (if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * set) or SVT_AXI_LEGAL_SNOOP_MAPPING(if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * not set)
    */
  extern virtual task get_dynamic_coherent_to_snoop_xact_type_match_cb_exec(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact,svt_axi_snoop_transaction snoop_xact,ref bit is_coherent_to_snoop_type_match);
  /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * This method issues the <i>post_coherent_and_snoop_transaction_association</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param snoop_xacts   A queue of snoop transactions associated with this coherent xact.
    */
  extern virtual task post_coherent_and_snoop_transaction_association_cb_exec(svt_axi_transaction coherent_xact,svt_axi_snoop_transaction snoop_xacts[$]);

  /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * This method issues the <i>post_system_xact_association_with_snoop</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
  
  extern virtual task post_system_xact_association_with_snoop_cb_exec(svt_axi_system_transaction sys_xact);

  /** 
    * Called to override the value of is_register_addr_space in system transaction before it is being used in
    * system monitor 
    * This method issues the <i>override_slave_routing_info</i> callback using the
    * `vmm_callback macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
  extern virtual function void override_slave_routing_info_cb_exec(svt_axi_system_transaction sys_xact);

  /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check
   * 
   * This method issues the <i>pre_check_execute</i> callback using the
   * `vmm_callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param check A reference to the check that will be executed
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual task pre_check_execute_cb_exec(svt_err_check_stats check,svt_axi_transaction xact,ref bit execute_check);

  /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check.
   * 
   * This method issues the <i>pre_system_check_execute</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param check A reference to the check that will be executed
   *
   * @param sys_xact A reference to the system transaction object of interest.
   * 
   * @param slave_xact A reference to the slave transaction object of interest, if applicable
   *
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual task pre_system_check_execute_cb_exec(svt_err_check_stats check,svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact,ref bit execute_check);


  /**
   * Called after the system monitor detects that a write transaction
   * initiated by the interconnect corresponds to a write of dirty data returned
   * by a snoop transaction
   * This method issues the
   * <i>interconnect_generated_dirty_data_write_detected</i> callback using the
   * `vmm_callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param sys_xact A reference to the system transaction descriptor object of interest.
   * @param slave_xact A reference to the slave transaction descriptor object which was detected as a dirty data write.
   */
  extern virtual task interconnect_generated_dirty_data_write_detected_cb_exec(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

 /**
   * Called after the system monitor correlates all the bytes of a master
   * transaction to corresponding slave transactions
   * This method issues the <i>master_xact_fully_associated_to_slave_xacts</i>
   * callback using the `vmm_callback macro
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   * @param sys_xact A reference to the system transaction descriptor object of intereset
   */
  extern virtual task master_xact_fully_associated_to_slave_xacts_cb_exec(svt_axi_system_transaction sys_xact);

 /**
   * Called before the system monitor calculates the slave address using svt_axi_system_configuration::get_dest_global_addr_from_master_addr()
   * and svt_axi_system_configuration::get_dest_slave_addr_from_global_addr() methods of system configuration class where master transaction address
   * is needed. <br>
   * This method issues the <i>pre_routing_calculations</i>
   * callback using the `vmm_callback macro
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   * @param xact A reference to the axi transaction descriptor object of intereset.
   */
  extern virtual function void pre_routing_calculations_cb_exec(svt_axi_transaction xact);

  /**
   * Called before the system monitor adds a transaction to the queue.  The
   * user has the option to indicate that the original transaction must be
   * dropped and split into multiple transactions by setting
   * split_original_xact. Transactions are split at the boundary specified in
   * svt_axi_port_configuration::byte_boundary_for_master_xact_split
   * @param xact A reference to the axi transaction descriptor object of intereset.
   * @param split_original_xact Indicates if the original transaction must be split into multiple transactions before adding to queue
   */
  extern virtual function void pre_add_to_input_xact_queue_cb_exec(svt_axi_transaction xact, ref bit split_original_xact);

  /**
   * Called after the system monitor splits a master transaction. The transaction
   * is split based on the input received through pre_add_to_input_xact_queue_cb_exec callback. 
   * Once split, the user can modify the split transactions through this callback
   * @param xact A reference to the axi transaction descriptor object of intereset.
   * @param split_xacts Queue of split transactions 
   */
  extern virtual function void post_xact_split_cb_exec(svt_axi_transaction xact, svt_axi_transaction split_xacts[$]);


/** @endcond */
  

endclass

`protected
KdHMW.d,/\g1)QSY_-a(C6fN4d[=,O^g>W.X/X^+==K#,cV(CP.)2)DT6#HL9#VK
7L>I^1^NZ.ECH+(,F?[P@:3^B>?2M6P0LA=280?)5#>^fA>^Q0_]Q/>EA+HfERb0
?E3]=Gb-]J2GggTY1TQ=6P-5AZ.N<J.:IA)##/g7&P@gNbF:Y_2<QOdB8W)#+bOA
c=/[E.Ye;7<3:1+\UXX_,L?YW&c8/Pg5,&Q&S5<T:TCQ_YE,G(Z#Z3UA?D]VU,C7
8^7@(G08:_[\E7fP,3U2V]1.WGQbX&bNFDT[1=25)+=JK,2Z;[-SbF/P4aE1K.Rb
>+#GUQQCe8DMfU6-:e1YA_&0Fe&7P8;Dga1=b]F:(..2f?>_[egUOEHJR5L=G3>b
4cWZD;A55]DL[3LWbO3_<9eY/9TBY.a6>[00&(g_SP--aJH.3P71e3g/<?D(gZ#P
<SPbRVKEQY^\MP55B8e4ENM]Bf,UT+?Mg#\2W^RD6]+-=YP0G07?N(B&N82eS#<+
5U?YO6e)f\)TJN:8Sa#BI4UL<O[>-D#GA2Of^PaaO-\J=0eI[N2]+JVB78b&]CWa
Z?AcM]/6:_>Y0>;H&<1((RTS+0:C3;>V_e]B<:.bcHQUDTe3]Q^(GR#<MSTVNZD2
,@.6g3W6PS9BT?^GBD<+g9J3:-EC,JR^ZE7>/>KZJ2JR.E+GBN6.aM2^aLY)WIWT
eBTOcU?;3)L/85YY]YMQB;WT&]SPNBH8RdAM?dX2055HZ6Q53XI2,41@QRY:SYAV
B^c2cdRZ,4TMI:afT].Td<gA,04&c>37+gX)D&,:II<VUE&5X^I200&O)B;+55F]
40HM26CKI1]T(-/]f&,[cDL/JNBR+B1M<\Y[6@?X9eda3Q1;4Ga-<9SX0P.#?NF^
L:93;VLB)]Cf;CS;KXWG\-][D^+/S,>GPQ,)(JW4Z:CI+GQ_f^1bPXF_[.:V]+1)
T[PCM4Y.;>(T]G7aa,B(J[fe_Y<.4VUIJY52;WGO5-9#->.=1A)Hd8>NBa\/@HG5
g55SLYH6K1+QXB^PFcK0+AC&Q\#IXWaR+0KMIFVZ#S9-WL9B=LM6@&._PF)A7P7V
CfMJB[+6UefNaD9cd.RVY#/Z.F>IVeR\QGSOdf^\Z(U/feA,K^KYQ=8]PM&SL,C@
IQCF43HQ+;0XO17W5-f1a>7[)KY/+gP@Wc@V7J?J\C@&2bVcEP65.J5(8cJ\<#d6
&\JIZW+>@If:T&EdCLYA6R&ZPW@aD63TPEeON.3YJT:9Z,3.V.dF##BPV>OW)YD^
I[UO)\L)>g)-/a@6bW-<bZ@()HC\RKL=.9.MW59:E92>#;:D,=3+T+PO83SQa]0E
_H\46Be0(EDZNR+b+>&3:]-fdCP(PQ:gD01QV_:YSI?e2?gVf\WD.Re&e)Y@(ggM
HWP]_H.J.:NT>IOb44@:QBFL_ZM,CV3PP.8gB3(G>.,=f7TF\:aT?7AUg1#8_\&I
UP::eW_&dIbXZ-C6V2M2QCE<APPW]LgM=^,U+?HI6@1;9Kc9JMEdUVe3+OVE+N\1
^QDI]T^Be3XU6G_;GT7SHMC2=.X^/Y=aBW1K1KI;V/E#-E1^>gGgeE;YPS-21RNG
D<>6YFD\8FFJ@?NFT2/GNN]F(4F)dBc?^+gYaVHGQIEc0D5N<Gf,ORDX[2[0@DW>
[;e1F<.@b\BS^^,F=I#[DWV.9?D?3d0@K1VQ>89JUN@@R@]_Pd7Q4M-1V]_(_/NE
@aL#1ZbPd.Ag]I8(RJgET,\JT2\FaE.3<=_+cLUXDX\G=S2RG>)Z-+W)8=g9I=Eg
3GbU4UU&@Qeg)$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
7G/FTHQ_DE.9:IV/(M&?#EGOJ@FB6BM]:.F>CQ=,@3/GeD7\50=Y7(^OK+CP,B#0
/UD2]afUB_.X@=O_UA0K0:d5aY2H(3N9BPU(QcN<<a>I9OIa/:@(U8Z:4?LK0bOZ
MJQQ]]dKfG#6d:ef6#XUbYgN,&cg[(V9UGg5ANYUJ@b#C\BYGDB7T:bNeBD=QF\b
Q>2[gME6Z[TeVWIb9?[_R(+dS[,S]IbFL1B(G\7g\FJCEW0f0Bd@23e+JSR39XO2
[MR@b,&ZBg.DdeO:ZUNM\fX8B(d3Y\;T,21NKP7;#=PZW7;@2ZO#:/7;9/QG>)&Q
/4G^Af(BK-0/R.@9K1M2M6V83VM@FPC>d2:6WUgVOQeOY)T\PIYR2ZZe[g:1DJ/[
+#\N1;]>^8K((QJ@QME_\[)e#,T@G.RcI.&5+RRa]MWPFBNW-^0,O:]>6(&Y>g/G
@E[:.W.,PZ9T)]6Og/:)12b^QDdVN_CBXN;](O:1TCfF0bM.1(D_+J0F<.OKb7DB
76I-1]eHIY<D^>85H0F:K]V@1]QGF=03;P5IWY97;[E/\MO;gH-d\FFb?J)I+BKc
\,T[@#L0W3=RU];aU:Fa9BF;H6GVSK7BGCb(#UAX7VJ=5:B822H-8>3R&FB^=N?E
/1N\Sb#S/Wc9]ANGKac,-d;XG7J5ZS^Hd-:RP4].3]B(EVX^33(a#Ff\NdR)\MYR
0)IW^-+(=SMJ\&cc=Cd_Y9cfXfZ#S01aY.-;JF7.VX(S@793a,AYaJ+97HZ.83AA
7U-C6OG482]?H.?L@&PJOg+M&&]-7E+D>_7NJ/R(LFZ_AI^[8/eW[K#O.59^b3-]
MR2LIZ3CK.J..7Y1Qd<44(I0Ogb>D:WE95:\@fAL6BT,[fTaC>,9YV5C-Y5ASOIK
IMg@7]1HNe])3]#TIEWE;M4C>P9Y.L39?L#I)W_BbFAI3B#;dP4=V3N2:5;S\<C]
&/I)M.8?=(2Z>K8)=9).8B&(\G<.)6aY:KdUOI><&T:.OD87cXAA[&J=89.YF2BS
f\L\:e79-CAHU:f-GGU6NQYI]4bf#A4G0>PNRaPA.44QIYd^P:Z=@O8X1Y4>1#:U
5?<<ZX@EK67JS#;(Aa2b<L>9I^..E?5Fg,5QN:[HF/D,Ja?.])NT(7JYB39cWCFP
S8VN@aK2\AA+CK^4C:U>OgAbf44[>6G@5GZf8#]\D5PE4RLf(YCBTO(,a)=B+V85
1?:N0Y3b7cD5)\,,3a7cR:L<VLX@@a[=D6&V0@ab\+@DDB-+PTOYMbeI4/RE@ZKI
LF&F+(8QH4e(953V-N?_I?AY<?dC>Z[#CS2J#:GR1HFNK^QRL:\eN)#>f;[?Ve#a
Z?6G0+dP,SFFd5>V(>^WZ[[@+g4&-d-6-PC5>ZQJBaDT(Y[0RZ9Bc[<S3>H^(eK\
PDR)/e(62P><KBHgU.,/ecP)7XS2MaB<M#d8RG<BENAA[fTYML60_=PD>U(JH:\X
7:WU-YR/D?_&gJ[L,D)BdNJ,CE7]a6X:+VICb[H6<NTfE<YCAZfLEUW:^Ge]dSX)
]IJb>,04Z[0.EO>)H=@#,KbGgJ.<A_/f_3bUFb4Dd0HBg]TZ92L2WMH.\X4<L;AT
UL_LYZ@UgC-_;CNN.BZO+(b^]f(D)S-I(Y51^WA>U<,L&&^D6P1Z9JZ4->ULP22@
\][CIe2WL/.G^EA86AS7DLBW]0&5ONb>0Nd@+?^./^-+;G\A42=M4Xcef.6E.7B[
90?5&dA2A5S\ITb:Q4[;,7A+^.3,a]GCQ8USLL.QS;H@MSb_<.MO7)+<G3;cfGfO
17b&I-64IT9&2(1RQJ)UXR4W224/fI#IO<Y^,V3\H\a<[5MU<7TOX;c-.[1QOPOd
<Sg_2+#T3YTPN:[>/K(6Ya;[@W-M1@F&.CD#YET1U__ePAL0da0/?Zb;TP9DC0YD
2)c>N7BS\#P1#P4.3OI[f,63ZaL)\FT<H=JQ0PV7DdAWY>;dYCD);cGS;#+HC/>:
4)1D5J;GONDPXG\Oc==;0+AGLHLRGg=G@OA2^#^Ofg2-7ZW[G#[LdbfdJTCSb@_X
0QZ0ST/a_XOV^<b5[=G,L(ee_^S)E6.aY,OFYf1TT-<aOC\/Q;UVY,]IO:b,WN/G
E=2Q7bYaQ>a95\cdH(O(XEF0c95(451(G55(QW\UA,TEB/eEefVgG9TZHYOSgOD;
R7BSR#a^\4K[:V#e@.<@II+]Cge)-9#>YLGWU?+[7B=4.g0AP4?]RVFWS/(GZV1,
g^7N^>2<<./^<)<XO2>g0O(EL7@:/+;]=W]2_IXQ-Rc__EW?Q^&^6WY/_]?H3e--
@+-A@A?3VY-2(\L0J\01>9[fd-V523&[X4/.7D\7^?+-;43IQ9HT4<UK-^+VIIag
;/RR#XO5OGIU1YNg]>WcgSVb<]^6OZ2MXH#.TZ6,.CaK=.Z,O2(/&OF88A_.2C/_
.J6TAWacV#.\H=e:(^6b919M;_G#FU/.2fW1\XGKBWU.2@/5\QLKM<ZPN_UBG^e[
L2)bg^Cb1\K>2MK2GTa8+,^&Y:1GCP;L1Gb:RIe7Q2.A-[@<gb)_H_DQ7,L/<[54
V@WI_(9-K(E<WH_\77Y7:#e0O6(Q/F#fF\gDD,)N\_Xa9-1=<TFc@F[WeJMH7?7g
Tf?B\_+5&YL6).Xfa=68U+0^#>-9#T0B/\@IZH_(a>G5CgGeJ[AE=1#f4M&Q,),-
>PMBZR1R]LOEbD_4dGJT<G8LBWDeXe/J#c?/TTRDRH@C&U_^KSbEA[UG6BIWO1F8
<Q2K]F4KF;XC]SK7PU.??RHc_Z_.^QPZH(U7MeHCT+]Ug4LXA#51X5fbU?==AXUD
=/eV@9YIU0A=8\2@;ZIJPIUaCH3-A2ed9_&KNQCa>JMa2G^-MEEa@+&JHNN7cJe)
Y5H([W=R9T[:29>G_HNc,RaHMJ=9H0KFc9,1cfHPS:=DFe9=Z9a_aSMZ&D79[VG:
g2_K=cK&K>A&1/,cG9ZM&RQ\[163:2@G=,;?SZAA?)2)X<I99+>O78_]HH])(34:
A7A(f??dNRF.NA^QY?G(8WA@Q@C(EUWO\E6C_gfH#_-+Q-SZ4XB6QJSX\&(8Me#f
+XN4deQc4,_V5JNG7a>EFYJ&PfSE<T.fA,(g]40+(3&;Q\/3]aA]O\DO38K[USC\
3-:,ZE6)OHN+dOb9GNYM4T;3/9Q-72>2^S\OKEQIKMgWa=+MCVZA.^MNH=]7.5((
LgTe0^0c=]ISTLMg&?95e2b4_Q4OW<,dK5Rb8L7,SLd1/2:H/-:TIZSEO_Q]<6Be
Ha3cgQCgf)c_=G93\G/KKUCW)H-Q06?7?\^)-@geLL-@V_/\9IR]:-LGT4S/_;e>
@O7)ReD.5b=PXX=ZBX<94PWBedg(N,g8Ta2.=c)>45g0NLW;C>R5b=^368/,Vf#J
:HdH[_HM4?VQ31bG@)fAG\UYP[IF<1a?4_2DA>,<EJR]\S@KEV-?6T/EVBggA/QS
I(<E,@;CAdX4?O3^PS:gW:^&=_3KX;EIX(g[B)Z]3[0.OM;AaL4:f)9>c.)]cbb7
Oa_NR^HDK^ebe?5)RX0>9VDJ68,/3P:7UaG4N5=BZJC<(38.<XD7&ZSgIQ6=>9bd
PSETaUJ19UT\.KK<DV.156OPCRbGecU9[3K+)FbZPG025+5G0Y24BZe+GXRK=9SJ
89U.Z1M/PP(3[^(AF=P86[2?IHD-QGdJMPF5U9ZX1?I;5/bKOQ+#4Y36X;YNL?JW
;<;LHN:CO&=Ya]+:>VPSB8T&=&fGLGP-B6V1CV#6=eI&@a2AY^@K.UO(-b@3_ge/
(.ICM(-SDX593NffMXL&[TZQUR,b0aL.6B7@D[cF;)S>10&R.QDTe\2WdHDg)]CW
F6GU00(\b;IgO^AVEUXBQ<4U)ZPB/EcXe<)FKFSE<+bLY\DOZf)#aT\CN8[)]dGJ
BV+Y69bb3G);6T7#UV9FdD=[69aD=NV>?c]KOSJ#R_:;15#6b8GJ-Q=ZVX8\RT5K
ZdKRgf7PeVbBf0EF45dXRS)_dD:,@B&MD>.AFSK-+B#USgc]eB;ZNa(8>D99<S&O
Aga2^0Y6_N(BdY;cFH]dI,&4FW]5BYDbJ.G-_T\([B0<Wa6Q_O0H@/eH&T0B4ce@
2Zb[5\bGWYaQcHe8dKUHO.c:?Na+aW\+BMa&97\6?9B^:YgT9TgYA?DaKIQS,f3_
^L/J@7X99f0+b=>D3DeO>gd]?]If)TdcJ]^4Y7TZ5>==>&b,Se8cD,?1=AB&JU1c
ZD0#EBZROK]cYVcGB-)P=VAIZ3:YCAL#a6[@HWCLMA2BeA1M:;bad8;OB-CV6aE0
7_2WDV,V,&[<3,/_@73K6F?CM>2S8YE&B4CV:AXf3>N)Z;])863L4Ec2^1c3Ed5.
Q68;>B3LfZ#A.Se.a);?^1)KM#7WA+ZVONA,9fX,&>Y.a#J2TJ-Y(3^&)CT8?41H
V.367e(;_dBLAT^cdWQ\1O+bgQ_cT[UOa<-+.[L=dJM)C[3#BY_X#)H?_cO-[(IK
0beGR;)/R,78[a+(/QF-.Jfc\1X_+T7SG9[0_b.5P/]T7N_CgH(NM)S?B5aMQaYI
M^EDZ?=M:<^^aZR-:NgSPHb3EXFV(;Hcb1U#<N&V8F^1]EcLPBKX@V8Ecg7TA/Sf
(F,=;OOFLd(T0D_T1;E1\;cf_#&PZ(&\K@@#VF.?OO;@RD^_S-F51#9KBAH3JJFU
=9<MH-H0U7F_,E21,6?X>24UJe9F-gWfLVZ:Ke8+/bHd6YWC@IOB1N?B(C:^<adR
NV_cdYOW>9_+,;/CZ&2X\6#AR<YgWX-X^T#3@PM-H)@Z.YT,A#,U-02b9@c@\9EB
Z[IQagccT_P)[&DS562(GfDgOQafXQ[(<0Q-fg0(+X7FHJ2U5OL.1]_4C#Z]Laa?
MUe3PZ+XO6=U[#RN:TJ>XbQK?Fb^f>b4N(b],0-.f1\\R9C8D,b9L^GT]0a/R3_]
CPQ@:Kb&-f]Uf,7KBdJ/YX\Q8#8.)GZ5<J@=J98,9G4d3XB=4gPF.?AO0R@25LD&
M[BeL93S]+O+f&A#XVSHeCfc^E=.0H-fY>1<Sb:3Z:,^b1EWFH_c<]X2WE.Vg8(g
?H]WJT;#.J(TU;-:PA7cVW@2XE[K-14@RX2)aUC).c@Z\be_a1RU4P+XeFeZF2Ud
Q5O@aTZc>Q<<L-#g:UM=]SPN.C/8D5<[J<?SV)-J\Od1b1[=fg-E1<K.W=/.c]IV
A,:@YT;Ld&+@gURTaae&Cc7;/cU;Y9,YESbIQ\>fR+IAaFM8=6,d(/DE8A<@d(J0
>T7:.]6J&N:ggaPFZYZT=bX@JK]D,J]\UG9(:?@+;L>3(MM>ZYD_<RFgW<e.1f8T
8c<[Gb1SLG/C3:O13]Y[^K1O\3T<MgKYG(?a.]2ZN<ZOA0^93Ib(OOBD@??\2T+[
gWE1T=4TA1+1Y,U5@]BFf0S[gIbe@:K2Vd[9&3GCYc.CWIa-Ef>XYR1M?A^:0,9P
>#GL=cV=5AT?V8gT.JU31db>^#V;B2ZBd4<T#Kbd?5&18-4&_^H,N9&6&bgRS/6]
Z#/^0c<OdGD.U6@3TDSO:g>ZW[M4d:-g93#b62MTJ6-?(7YF2OBXC&F?<UaBDJfU
KB4Lc:\.]dAU#c86>ED.C,[H)VaH.KNcd,)CKQ0MA&P>W@0&XX3L#][f;=_G77_J
e[5_)de1(X]=d>Y[&],KAHC10O<d-EAC0?D@dTeB,7XBB6_NaG^I^e8&9=T/GKVZ
PW4CYVQ76^OaRVGN0/bS?7N)QXME++4G6@VJ=c]bDF?VRdaO,^XZVc5K70\B;Ca+
/0O?f49\4>CW4(g3B8LeUOddKK(UO4#FdSS\e.f:[L.VMLT/5,b]@U1X=5ca2#4=
_/XUcB;Pc;c.#U7:KJ?)RM5+CeJ#RH-HWXP[MJ\I;@2Q5(-G:Ve76QZ?=0JcEWP_
^WdM<(K2[8=RY=EHU7UP_ZB[+M)<Nd+K&::10Ag2VR/<?ST^?g]]EA#L>NU@dX??
[M3LK#E,58f[c/:/^-/>QTE1KIcfRCC-)c0daC(2XD@KXc_2a5+BQ#>VACbV<)c_
V:B((]4A&(MN]\AaQG+U47FR1,?@CHX_W/NVG;98_d>g?N/?)?Q9BQZgS#<eYW5:
T;]]F;.9&b=A:>@e,d+&38:N-RJE?HbC.g5<VTFU:0IIV1MC_[CKCDNNdgVg:[FM
&]G<BgdaaA65_RB1fb,6XQ_30J+Q@^L^b@/eHZY]I6<3P+W3)Z#F0Fc1.5@@_>AS
b?ZD<ca&=>I2OJIOg@QNJ<QeP-5_Z8b/+R>&6TX-I[Q9Q-G0fGWE56U?M5NY5\CR
ZaMXb3ff\-^[0^@CRIaY>^S?2-Sa.R\Y#P9J\2]7J,@4LF;GMPYYETb>BaR6a]JR
W?8.2.&W?aa:]NDgOXNG4OP)5BN[X^J(ZP\Eb7_)]71.VLFdFKOZgGZWE[0QEL.N
]Zd8&@R^+;+OI#DL1aD9BD#K1[&8DYB:#\>5(J\WQ<1+JcO0I=:0,fQa6IX)<I2b
#]R=^/E7SZAbf0LVb<UK\5KfRLabP;F?g8([SOY\SA75WHH-QTF2UN,]?edbKF6H
fB5QUgKLeE:aQe\3^Y@(PHTO+EeZFII>TWB2Y:>TW@5A&UOSHKXKd(.<\\a=<b\/
CB/SKc[VJKGCZDVHWTI=P6@7+UXXKV4M2Xaf5KOB79KDKH5eHgCE^de,a#1S2Y\5
_KYIYQRQK,gcKJVODY3M6XZJOF<b/L@YAK74UT2;G9acECfJB/G4-Yad;B5:[S5.
X2-Qfa+JSS\FHVKP.SNU^-KMaG5DgO78@:6eJ_We#FOXZY<B.022BD]XS>N2b-S=
R:d++d42;b8,XaPCg?^&?:I8<41T-NeE3=02g,GKX(ZJb5+?^]SB:WVIe&NL4>S(
\S;7Q;P,VgM^ZFCKG))6W3TbdePW@S5Z=dFNW;LU/1>Y0;D3OQ[T3:?2G/(fRgcR
[_(^:3GE];>I+5Y2M47\/PW<>\3<TMJR?P>WeaB@CFD0UU,&((;?(R(C)MM]UW/M
\Y@?Z1:VRQP-FC\QHK,^S+JEfLbR[>>a/c]-4&@0.c94dTLMMZBS_BP=DW71FCNO
OEGEC@&AB7.L0G[cL51\5WHW3CEMH=abV_1U=.a-Q.TB6GAB(NLGTME\3Ec[:/;c
Rc)>5_LR0>YNd4I;N4^d0Z=?Ga[C5cb-2^EA3LP->D.CA2fHX3P:a+#F5.<RU3CM
R]cB9?4?5TcE2IV>@E676S&ATf=bWUN0b<]W8<b<;@[+MKK6V]c.[)O[]V4\Q8T?
)L;A]_)Gd@(7+0&]&/#;U9R1.R@(<a/QK^HM-_\/[X+7+MJYH<bY<(K05F+PF3L;
AEV4S&NJXL1.Of]2T&;>b&Fb7RKd52QZJS#;GC\\[f>@@D42e7LdFG\B(,0@^)P?
ON./-PKQC_R/O,[O#MbS@[f32+##8\DJ/WgMR8(-X&COeM:H:D5Pe;2WdR?4BFUY
fN(WKGR\)fdaM9R_eJG[_9EbJ>G^PL4e</-EW12Z0b5+9G(agUK5VDW5;L4EP8gc
C,KBX-3(SM/UUE4;@X;?<1?DP5Mc?M3[:0cTK/P?(A]H-.UUA61dUQ5N:U0_(CA.
1C2EEP)IPD?N2VdP/^JaD;8-aNW.XNUcHLRa250ENfe(I++L2G)<:VB([bRY05[#
-g6e=&/#Fa<Mf);YW,C9&bS>]&GC>DHg4[H45#Z55DH@:J/O5&dSN.TH2Ia,JZ4/
--C53M1G]DL.,0Vb25UGD.dBJdFa&G+HANR.7VS)>CV&db2@:3QJ_dWS=c[/1\Q@
#CO:<Ga6GIV(C+^]fKX&gWLWIDRa.\<2)eXB&b])3+:(bTfOP)Ld?_#aU>@R8@9d
]&NS@<(-b0PMeX9T/=dYH;6X3)TTPHQ#4&[H>UWA(Eeg1>:[78-daASS0GN3d7+L
X]+a3[_+BH?ZI2faVL:NRZ>6cPDEGW_6d?8Z1eSV,QGad0S<KMWbPXCf_@AH\I/N
b+P9_Mg1dPKJ<L:_J#HY9Q[)0Q_^V?VR[7gMQ66_ebUFO;NVZ[C#89;c,-VDTK^_
R6U51NHJ_]J#(3@WK^Z<e.#+bIH473NTFfI.RNM/Q8e&54,5/gURE5GETe@>=?3b
:EO-95ff[YS/f\L/DE]8c9REbI5)a7^a3ICLU\>@@GGIF8d0Ze-IK;8@BRQCc:M)
)9D+C,>Q6NUS\V<LIWLF=4T@5>R=)b^8R0(>>]QYc+Y.5KRD)PCbS#W9A>Dd5=U]
N:,;GSL5&?Y772(dZZ>V;=U3S&(&3CQ3M?\JDGX]c@I=ReM+O)U4D:#VR].Dg7GE
]dMKf[7MWd?-4^[WYU:JL3ZCB6g3.f<0O7Gd8DB\9K,AIHKNA,GDF?O0O(12;O@(
Q^JSP^3aIA=9@&-&V)a@#[9T,N)&]3_f.<A7@Agc@b;YZ;3DVZHV+>[MV,g.:K.e
bQ.XELR7C1O+[HcIaD;4)^Y&bf\2S[U5GA62U5Y;U^#H>Z1QITKS[f#9WeU6)F<I
VQPcVeY4VF6YRTG(gT<[<c)\H3g3V5TACL>:_/<#G5V-?\3b-;;77RR:+JX-I;]-
F9&WBPU2R&7.X8CE)bF][Zg6f-Q7W^0dK&S]Gfb2#P8,[B+)=#Yf?,P;DG6.VNAc
b8;0aa_DXN.]VEA3]RBW7L+>:Ld]2T840^40-U572KCO5ATSa#R6dK\.RB?S^1N6
.-A:C,Ae61W[Rgc30aPY8MSJD]H,GLbG6E.fcT6W[RH&E)\NLY47fR62]U2.1<AB
<;C,Y_QAC5C)GW(O<>_/NDN[T3)BH3M\LT)9G5L+^II4+NPT0Ma+>S:V8BEMeS6T
(HINL0PNV,#RZT]e^e]]QQf,PEO9;?&OZXYag)UJScV28=\bCg^KYbNOa&X3?C95
(U=^MTO4VYY^G9B_1MC+5&8&Zc<]MNETA&45JE^Y&\.0B98B3?Uc/EcZY]9S<#\I
MFII&L[W7]Ub=TaQTR^NI@^#[4MQ:VbI:3^B1+aR/4?;3YEA?.DU/BR/+3@OX\&U
#]Y^=VPED:EL5E]4)N^@<\W4TcBGPR6)4ea8R2U)PSf[af^=?8f3\fdO82#&M78_
&U&>E1E4W0Q/4-[d\])]7[7O^f2/>g3U;b3GF<TCZ6VDc[KC0T)c:3Wg2S^9g89W
:D6#S43I)Jd2_aE:08._)2\\>4?I_D_VJ^@DE#fURVMdQ9=Y6N4GXH/Y_cUFgMgM
K8+<fL\K92P6G8IAH(L6)Ec+gLIZA#JW-P&(.J;B(RXcZQ;e.HDK6)egNVI:CF#_
f.XLA9_WG,&?JP@,/f;YMN2?]++1IIa(YQOCZ[BV[M6JWY[MVYfSVE1#(A413#M8
H[IP]eT#<TBg5W8-^YBP8UH;7NXDX__5eCZBLgb5(9f?M4GHHPZD<R@GLgH13=4G
79:)=CeV_gD)RY9V1g3U/QgP8)J((VIX(3GBaKCcRO=BJ/9@d.c[c7I.RS6VH5d)
:<YDaBM&)CN6X&9^Hg,NI#]a0:gLJ@]WVMMVa6H2LIVZO\cCb>TKTLPS^11UD3#Q
g+\.;-f.HI5_Z9.OeQBGVJHXYJQTGKE@1.TR<-=#>S,UQbS8>Ldg=+MO//PL?&F6
)O<>O0(E5<><2[gQMTH6f:cO&4EO/F=1g08g,R8LCN-0JJQegYWbNO,H\J:-:TJC
(R\4@FGR<C2V+8X-:2QHfc)S>ZK38A_Hg1gMfZRKF1PXAF\1]I-@TQ.Y)&),B/#S
J+V>;Td>_#[gd@V2#9TgEO<CSLVH5c4^_H2MSV5UHYbU1JM3(g:1G0f6EB(&a5K0
,3=TOCL]Pa^&:[KXFXBWVDgD2\0PDB12ee)8VPZg)2:&8.K2bH&1N3>J-4Sga_W,
d?MbF0@0Q<0d.=?21_M\<;G(C1(#R:6b@=@M]ecROM_gM^ZALe4&LB]NeTMTT+TQ
;&aK6bccB/0I0LKg9?:SM+28=3aaX,7@+]G[66&BKD]?,M1V=4Jf1aR&M(O8eWE&
))DBL-7V73IbD9S,P(_++3RDMYcAB-.OTJGK7DTZL>6:.2(HK>,3H=QfI0WfW66>
-9D[=/\=<BSbN;)]R?eR?fE^K.MJeT1G/M@I4P3DL?]E;R?\/]\U836)^ENTdD77
DT<;=[3OGQ=OB9Nf[AXX_JC5FYP@W++#L9gL^c#:J[4H(eV&2(S9P,A2J\D[=,(f
d<2dS(4-.KgZIaNPT@,/#gS);3c?0GUe0-BLI29d)=9@g\>6VX);0CSVW8d=&bMe
EZTAIeM[ZV#X<]5F7CHf9e;@SfUc>>^K@PF/[^W,YLM]K,U3T(01T0f1)^^VgXY@
6Mec#Nd6N3L]W+O44HbA=U:<P?_;MVUb7\E^96L9[f.db[eDf=_dI4;@HI936?T;
V-b7#?PK]3Y=cE\>QH/>JG2]A<bO?+X^N648W9\Fcb5.D/7DbQQ>)7>&2@N]#M9=
;Y)H,A(D_-T[,/3X#TQSIgQMXA_F2E<1?Zf4O+Y_Y,N]^&4fVNG1^RH4bD<E#O3&
_=ABK&_d2II6I7#f)0N8HeL)=EMJ:0,F;6I;;-GC/ccQeEf\PA5[B+WOURPD-J3S
21DffO/@I,P4[</=F[T2Fe)W9FI=G6/fPZIJ\82-Y(H^E8g;Y0cRe,BLf>WgK1,/
56>^-_(DV<]95d,]E/,B+]#N7dEMZ3C,gZI-GS7DM19_gUEVLX>9G/0+Y=BU&&]^
#C_E[a3dE=&E9;DLK:8PD;^YIX]-EY10W\)01eaIN2^J]M5C9S?O>W2JS021/2AT
U9Z3-gUV?1@;#053#)?J(2dVI:(Rb9KL:J&;&2[H5eY=;\ULGO7=LLb>HVL=@5[=
T8Q>@B=cCX>FY:T)?L<8IgH,1(Nc^Y.5YWYN+@:0(K]YcaW0=N]A@7bY7(E69MCc
_9N6eWA.NR>@@>c/@S^C]4F&[g2B1>AA/<0<a><8g9VWCX^35J\=b:N+\Y/+4TIH
^^-?1@:4O>/FDb@a^1+0&9>a1:dUFSf:?4@ZYMK[,CIRE[Ib/6LKY6IWM>U#d>b7
30B6\YRB?-]Mf(V&NDCLS@S38Y(dIBG)eSb)]3_WROa4WJMcO/KO^(I_72^e>^K.
?IK^\fF]^ZQXbbYa-Y^L4[3RO07(Z:-AGD@0V\8O70eCFU/#_HXKK>R1,g=_dc2[
)\=O#=b\O\[Da85_aFX7PKP#<G@eCK1I;,e<]JD3Td+G1>+WeBDFbeF85V2_&cTa
Ld#E)23CP5B0adWSAcEc<#,5AX.^9bF8bJ8J7S].ODY@2)_Gb;7]<9?LCK??3R=Z
05TG5S54Ca_MJ:HecZ>.gAQRX74L-SBJC2BV=QO?H6L?ZG7b_bYXa,cR25dB@+@;
JP+24530(8aMMP:dUX_5176V^[5+]6TAbD_P+bB3@NY,g8:8L/bDZ;^g;Zd>K[RQ
F?_aSQc;UM-e(_+[>bVX(N:dX[8LOGXE>(e@9IZ34H0cBL@)\68(Q+SJ@ccbcYdg
TF>^4(G9NQ;:4M_A//BEEEFZ5,b.B,&#08+MU>EcG6N4\-d7F57Ja.BAf[Ve.O:=
NNeWUZb;AB)6[-AC8Kf)9e09c\D_@:OJGWP>4Qc4]U4(V:5(QO<g+AE5H3\)]bPc
EL#++@VB5_G5=WL#.T1C]Y:WG@8XVcX1;S;eIN0SIKB>C8-DR:JKKb77+BHEKDNS
8f:S5ZF>=bS/9DSgJ=VG^][f8+f>Y?A-56?Xga=DJdEU7W.A;>WSLZ9KSaffBYR1
_Z/B?Z2\;B>2,]RL>/eZ>QQDGedK6@1ROJ+TP#K0C4@D9&HG_aL4-7cICJ^ENF.T
-DT9V@DVNM1b]RF6200)K.T.)ZA;BYd#BC)&G-PDY2616Rf?NYP4A)/K89Taa1fS
J(\]&4]:5#X8K,@T09.Y>LMV>K0FV>YdO<KFdJB>6[/U2gaMVXOG8ALD7WBf&+/W
eg=5S5:DZKD_3_NHO70CKA.-+51_C;LC+_<-\SQKAZU+#?60L=RR]_8^Xd]4a122
(/AV_a@AHN7O]O=9?-P?<6:+LPe=c>.D-@@dG;aRa_T;a96T:7UE<TbESQOIAPSd
,NfQ5E+(6F2&K=9IB,)9f-7,M+#-16CM?3/+AG7d0VSU5e)S4E-Qa4S+5F463IFG
JfF0G^GC=5.5Z.;:XBaLdH&RKMNa4cH8:gK-=MI_aEFT,PK/XH01CHS;]S>OENM]
^dCWH^Z20;H<GBWSQYF3\eMgd]_3g^-F;)VfW1P98C47/-4639P>-_@\^GZ>\0UV
2Z:CHO3)bEM;S#/N.4e6Y_eA6PLF,NLQSQ)^H[5F517MMUg+CH)7\36IY5G>QWaG
[)QYFCSV/6a0\L/.I7K5[;U&^Ef=]+eP0F9Y,gRGd?f,0-K<32/-(.P.6X.3Uf\f
DB/8D39F.M1a3_a17>S<NZHW5)(JK9.\[=<X@?=2Ag_<G=aF:fCJ6W>4Y;))RI.X
UYL?b0Ce;3+M^F_\>28PHgF3WAMGA/DZ?FVd@HDG)OgZ&D/0JF5HU,\XIa<dQZ8^
cL23E5WdI,/;._F[/7ELG#9P=5K.&,.LV_>aJ&55OBW.)R1>8]Sa6>BJIQ&c&JbX
XE78XNH=S]B-f;OI(14OWM9<9]#Z.NVa<dc4)L=@G>H75EQ&HfG::.;d@M-]efMG
TQ+Q>f>EM,?2,#JMbMG?[-M0(VBg-aBWCCG@7(/P6UZQbU0TgALHMKL)C>USbLXV
G.A3_2I?(208Kb@d_GOL/[;Z>ABA](1_IR?O89JM7d2_R38ISQ0M_;Q4R+LP/7><
\N7Me\[4;,d#1[UX-,TD63:#U.PgDS1g)B:O(dXHA#/ESaP)E3;DM0G63E[^e0GZ
),7V]GIaS\L4F]@JTZ7c.E=ORAW3^&Z=,7WaVX:-BV2BMV,ICTT+<)LNfJ9HVVaX
NB.\V2_T>7T_V]G&Z<R;UNbLH474]2#8V/^6[:.X1]9Mg\>fHaDgU7/\_.TGEJLe
1VD7H<ST4W/QNZG=EPW+N8Jd\RW]^6>R=g+MD&0BF;-L/:T>9VR#1#WdF(Lb(Z<P
XL>GF@4_(83[c_DF2IXceVJ#QH2>8S&X)Y-U,f-&a1HEF-2fK6Q@E#c02MA,;1#&
YgG,,5H#.8W[T2UeTe6NR#ZL2UC6&/[,0T\-7G:QUdP>6JGXN0(>6AVNVd5[C#La
-QB6QT@+VVMH&5LO0;539T:TN&1gH&bYDFKZ8&<1D5/G&L6M-QG/?6\P[U?1R2YP
Z&eb6:K6?KDES8b+&7VFAZ;c_O+dKbP+VBDS5eV4/G3DO^[+&R_X@cGb99E::K)G
9f7MRV45WEdedAM]3WOGdP(2/e4@]##@5(GO0=W#LXeSUMUeeFK75#>(G>\45ZHK
C6/VH/E_#,7f8XH<YaT(Y932Y,0>+NG[KMO<:UGC7eeJ6))0C7&fT[M(DTC3(9-E
;LJAEU@7P_P-gf=B)_c.LH-N]+W<eaQ-)/R(CP9&+5Ed3QKfYG[E;ZF3HRO0e1[^
]=[gYFRW+3+]IcMRQTLDdW>KRgUH:R0VX8.X=B9@@\<90YSIH:PEXgC(&O^NLBJL
.BEPY9R,;MS;6]JZBA(b)BO<Q:WL^TNJ@Eg5L)Z.KX/K;)?/g]W6>a;=+Tf<J@OL
\+aINY?Y+O+3@VDP[eA1dP8/2UZ#R^7Z_C#?D]DY\VNO3]<O;gZb=B5;;R6U?Ufa
bEEU,TgV5aY&@]QH20C=)ZSH879&gQD7LOR=aY&^]e<S=@PJA89GA)CF#KB0WS78
H0/[a#?2a/-38O6T&)8M8aKfA8(+6gR287Y_a_8:<aVZWI1MZ;-f,Ag,N^&##&?@
>Y+C^)R#+=f;^T0VX3?+@P)4Y]FAR&g&P@(#0a+B1:LYEL8Td=QIR(3g8C,P7b=I
f&O;>9N^F.-[<fWaDAaK.\DFY_5O\(9N9<L)+[#B0J;NP9&Kd_C+J@G1EY9&39.K
U-@HX1(<XbVFe(&57[F9B4N[)M^8N0#H=69;ceU(beHA_OLKId0<.MSYJRND9Ee)
_[gL=389J\>S^6^G;/LQJUBL\9R\B]Q/8(EFHE6P4\\(cU.:_54L\,VI_5C.@:]+
YN\.9;L4IQaFE3:,ACK)45e/H-Fc@9E\W/?^T.M4gMI2De7/YJ>>O+<)/cC>8V\P
#dP_[<_J8+VE71TXeJ-NAAF)YReDD85S@ZE,cWD=A@<bb@G<5E9S,?@gEJ8)<]J3
PPI=Of^&):04VPD2\.6/VHR(+=8+W&]M2L\8QXF43eG(bNKJb0.DFbRLT1Y)KN](
7#.6Ude,X=UIJ6O(;JV;N[II1ZQ6+8VcPZdNgHg/L>9^RG&b2+ZQBe[:F(YLOa29
[D/K1.;>M_<)+[:,0f-_7c(,68&fbL6@WU.QbMH\#B9\&S&ADRDe_fM^IJ0I+]4W
0A/c]OPaC^<1gf22/C688MWJG?B19WGCQ\;[3;XV3K[2PO_;(E.E=MAe[DRZbH#P
L0H\KAIHRGB05B3REFMa=dM&d[<dAaL^ZX@?Rc?L_=#3Z_B/gA2(QGQ8dbD6Pe5B
(-GXIP,JK0)G58COKLI&IXf.OUU5GA2L&/K(=c]/7)07LR_(Z^;8(Ba&(cgDGOWE
/E])+F_MFO@L2TBDH-HXPP:X(KS=C>fBcBIX9&@@Y#C(Y)Q\N4bHeRPC^SeF9,:D
<+bCbJ/FK+L^L)&?g]OaDg:IG853>:@^@dbdRZ.FTOe7DT)^dd>O4)C-@Oa1N2e:
-WfNd[</g_A#5;F?,P(K3I[J.4eM2d16BaOEW^@,8Ug6=C@gU+(N<dMT.I[<3\O^
7.).1KY.;^?+8Q8.<..QT=.UgF[eAXb])]QP6Pf/b#E5+\=Mg0OcH,;@K2U\W_H>
>W_#FAW;OVQeTb+M]Y-Rd#\,PFg^FVZ0H19BDD)_E^>S<CJ5VG&C1U,WT3470LUV
LGU?:\(fU@<B;D6f1S:a1YYR:7)T_.W&MT=CadaaWeZf&K(M?BS;/FF_9afS1&<?
^d-;^EBeLB9JLXXIQW1--a5W_9E?/ER2V-TRZG)P_E6-LYY\U913/RR>I8^]1E)1
aX0cI&D,Rf.H9.:60#YC>YNeVSf+CIT&S8XV\B7G>QG\-)W6D(PS;Q/P5.XRX8.U
6Je/:V)8\]Ba>V?GLJI748B+b]TED?3\\9d0=S]RJd=D^DY\/];bK_@^)fUS3E5]
/T\Y,@KMf?G2YN:bd^JQ[6PeS]VA(,_7gJ:de6UKf;G4cC>GX5fe)_W3b+=ZB>0)
(=Za3b8?V_384KTdBb<YSB;MT4Ob6#?IQN1NecE99a=+7VQ-(/WXC<B:NN2.gTK8
a2M7Y_HHV#3<AQNT&<XS6>>ZU]ZQ+SB4#Q;;a>fWBYg+g1X<AWE3=WV0RE(EFPH)
-;::S7UPfdM22.MM.6RP4NI[^ZUH+-#WL9:)<TFK3-WfUK8<W2:I)IOW99Bg^C&9
&0^+5<5S(2SNMb.b^K_;L5UO9_NS74SZ<I/YX;E6QNg8#2H]CHJ+dSbM#7-[45_a
4E;Y4YD#f&@3Y5EU/51NLLI/8Odd4C99.7_R6C)V]6F&I>;\BFZ@F+Q^UHO0X1IH
\8+3@3BKA&[DH)a+@+V79,U#cNB<K0(E[FTWLB:LIRb<5FF4O=(DT3JTe>(?RE#+
fG(R_b6CdV3=UgL5YC(O,.3e7AO;KE><&;(CO5DP&aA4+0ZN4Kg&_V_TTJ3-S4;K
II?IANGdH#0UL=[3g-@F#]1)b67]1beBLc=c;Yad+&=afX)D90/;:<TAFX^2fGJf
d7:VcDA&X;+=AMGAECI24b8WacF/P^O>_Y<<1_XL-\ZR^^PdI4@?T2Nc=NgK+GKF
KS&Bb_JD.<+O>FY];+@Ma5E:S0.LBab50FNH1F@/W:HFcfK@79[]21K]4g&V2>\:
c&9;2AY.fBAL3?cC8N;#T6?Uc(H]0d\0NJR/;=J#EKZDMZUHU]_?+8[RZ.;WP4[C
>X[6+W54G^YO^9f>>CcL;c_M7#e_H\ga8KgRcG148#Qf&C;_W]BB/:a.L^?03IMU
<OK]/JQ[RB<Db7=]f/f#GT\]fUf_#.@;G<_AZYfd_+O#Y3,@P?f&L48X[-LK+2\+
d-gA\CbE4WYHN&Y1UYXW2Ua.33af?H]H2LG_<>509ZUT6^K91Td7Y7F-.a#c5+D3
EUaEFaLFL5YQ8<g2BdMCWLSF:S^UBF_DZ0^VSf;O@BT1JBO:_4#NFM@O<ODFYD/f
5I,,X[;Zc2C2A\6PZf]1JVS6gL3)c6g6g_g8)G&+#Y9HA,6G..K8HLe&F2VJW.,-
@1FgceW5Q6SY;LR6.REf2]QSB5CbNJYfO_D^=&UCec?5=;QNRVV<?./^[TIOfC=-
FHR&/gY.9?I0RQ[1FJ95,-b#CY;IJ?cDIX)aZ<O-ALT&Xa<B]]5UH71<]Ge-_&#5
;E18@YC9NbB:(a[)aCR-];G0<[_]-2Cf?fU;WC(LTRQJc=U[U7R1B6?P6R4b8ZCC
#K7f^E3R(MJ(<WZ<]ZHQcN#)]g.bc;A[1c6.-7XVGXd?_\S&5]9-JMZ<FSS?U4],
T)WN+7N_JH3EH&066&Y\VPC6].7Z=DN\L;=,HAD3187I1,.W/H1aFC^3L\,bT-#9
:/FXF&B9Z91M?>T;@;8YXM&.[]^T18?W13MO-O>cP=E/TKNd#[]6T4(&)OTf+.,4
7IPgf\b@PF]2\/<Ief+_JLR3bXW0E^B<]^bCIK#[?b;/N#AC2>3+FHGOK@Kf20^7
OFP\90Q^78Q/HJP_??O72Z+UR3dIabZ1#<a:/I/>K.XUCQfI)7g/3Gc9g<N:2+eU
?/^K&P?<44/XJ.ZFXGI_=N-_A?@Mc5^<7SVS1R/f^6T+^HD#IXF<a.5P\5V@EJGS
AQ<U6\bgaaTD]LSD^_<62ZTEX?_Y^B1P(c4O8JF6X@@PM^U:LTQG>BZ7D;SS5C5E
:OB=Ge,Q2MMG2YEdD9d3NV/]Y-0YgP]dBc=#W:YJGD7I>>fB90UJGZ@1_J1HQKF9
3E_PcgEPJF5cE\X&OAKC]^QHF5GUIDF_TMNU7_):^daE+16LOG,/2#7K:7IS6(JH
eZZY(C(Rd39)[TRR_U]&;RF4[aVF(6gXG&E4Rgg3L:IV\/PS[,bUGDgXYQTf-4IH
W:SAYNT,92MBY<^#Z0eD22[a5b?REU]ddC<eR[1-V+PfP+,6Qf:d4KJL=UbRZ#C\
#T3MX#OW7,E1:aHfOf3UQQ-]Z@&=AQd:?>[ZQ4/C_]3LG1KV/BC1b1(4dgG26++A
^1EZ,T_)+LRF1E3eY(F9(.g(M))E4]DQeWB=M&XX-Y/\O&FD2c1VTSU8;>1HYIbZ
e7UP\2TUd3+&D8QC7bNK1([/dd#5.PD3BCbQ9P-M,9GWQ(-PZRQYUNfU_@=]MS#X
;a,],M:?a0MQ\_0L4cDcVZ2#^V=Cg=\E@=X??NJXP8Vf<GANc#L<(Z78IC?DB\SC
=MP2B;)/I.BWF>[@T&?6-_1#DAQ&3CZ?d9VN7M\ZcIR+L9PUE?[2N\M_B/UO#DFV
.PB31?QC,C[F:O\#a:WER2;VHZXG>;5=<8KEGHF=CFgAM@XUD=,63g0eGS<\=2YS
CVZOI7<G@N:C6;A1;0R?[\)F\g036SSfb8Ud7O?f1?eC.Id@7O@LQ8.9.b9WE<6:
)gK-O.@_2@DP(#9a552S26G,Dfa5RG)b0/WFYC&HOb:]80XB@E6^,OUE0WXD2c(L
3g<]5e_577DN1()6a:c\:94IMMT-]>9IM&dR\VTX2S(dAKXQG.6HS9BTW#\5ddVM
325NEW7GWV0K2V-C-9JS[0Kd@?c[5E;OgGWGb3T2AbPB-_AJFOG=)S1NI)be)gJ>
)7FN,5:M4KYX45LIT_B0W06@\:\D@KZKQ=\M;R417\I5R@0.cb[O9BY@B_5(DSZH
d)F.2e5(5O_K+1/D;^MGBc\V#NAP93EFGa.[U#N0F<H<Jcd@5)7>381)CfO#410&
.X21fD-P;8]J78.cdE?=8eC0I[[1@bg^:#LAX0;Z=#(a?_.)@JH=+]4@gW^/OL=P
Ca&/9-5b.SQW&)PM8/H8L\5;T97J/K))@3ZWdYG.@<I>S8bCQBQA4QFWg9MbS-OI
^R>I-\U)dGOWLY&:N#LLM<<MB[[U:<][NQ0[JXK3(aW45#,EU3P(aR8JXZ+1GB]/
b0:D:-b.6OS<G3Qc>d-L23NXS3B&G)[O6N>ec:cU7VP0GePRG6][fO_dKcF=_Gg+
\?=<f)8.8#ZMT(D<)KO[P#CJ^DBCNIF;,deSDDKH&Wb??KEAQ@P=1ES:?F2caJ>b
;L\<UVS0I<2BXWU4SEQ2UXL,bLYW#D/#TW_X(\60+e>c2N6KE;\JQ2b(&W3ZO[+,
;WGY.(65Q^dY9U2AYY4&\cGQKE]dC;gDf^0I<I?D(U^348Q=1NfQ6?>cb9^X[PLJ
b@(OLT8P077U+Pd,T)BZA?TC>RR2ZZV)g3Qf^=FD8F3QM9L->2K)f,aQ-;Vc#G12
OS/B:7gG&=:C-Q,IO;D]#\:C@T@4XbI^U.K?G4VEBW0<VU@bVG=I6E<302P+>QS>
AYTZ=UW):-#BRVVCCOB=Y<gT4F_,@e+(33GY7><,dC\9(Q9L)KED0dBEfW5b(U6[
&PdeP#TA6&L3=.UIU>ff.E1_OUYW[7)(YJLA.D7d.C[6a<A@b/_)Q(aBS4b),L?<
?&Wb]cTKNE31U@@EPOKGfECUJ,gKDOPE[0K,M4<.^VS;J)#1+8[)BUR)8HE4gD&a
L1-M)<5fc5d[>-Eg=[ee[^F[7AWV7(#9B,:3dF.ZcUSHL-<]>M@I5^4BTdW3J>I@
g]WDYgATI[A8UUBb5&X)]1AVUN3@73=C-ZLB]\J@-(M@c>^--H[cSeA]](SX8OCB
RZ?TS\14.bgR;DF4YEV+^S<gX2T.g2VW,6A_\A#UI#Z4F)SZ6_XRI3&5H/<F,&\)
.<PNTYSWJ<6ab_F8W+7JQECGQY[X^eFM#b)]=3NLNM6RX6V7@5+4>8],(OHI?4]M
WKb036C@510FD#LRX2/:M39&Q>/#[1&c740/J;G(Vg5UaZUE<dJI?OZI]=O&T,8,
e=9BX8V0JY+<^\2I)I^>->G97ULVgRAE)G9^^T2Kc:\2b9TLa(;7_V;SUX(K^\BG
C8HUJWB10a5_\TKF<FF>)VYGcUPP<-:8SC&bdG.32\7gf)RZ/8]:F0-ZKM(\;dBf
:V?\M4?=55b]>U1de9M4D+CFFe<S(3]&CcT36+5f2[.\3f@>=(\ZH)P]IJY>Nbca
.^bG<^W\2SU&QSF=1]JC&TT(39c6IAF^S07bgL4=;YG&>^_@W?5/12O60Zg5N]d<
M-GY.<CGN1K_W0]>g1dPc5^5^V9J(Y])a.bRO+]IIVXHe]74cN._Vg;3.;_,U/7H
CU\=gbA:57?/EfeV.OeYEf.gTVRe,7\5LFX?Ib)W0b/dEGON^<&HPSdN@.@O=ea]
\.d//\CSKKFY;SBcEK1&6bZPdJf:[1c:K);KM)0JQ.X1@I]3CD;,<S<:T/WLdI.Y
J-0B]#UMNZHKgV1USR0Xe7bddg.#Q^ZGf@G6D;aKQ+7=WVDVP4WS1AXc3Ie0=N9T
5f8?(S[fQN(2/IcY)5K>DAg(KH587/+]f+5PeLf2cUfdZ[6\VF&GU]dB[=4eF[GP
86(@6C;\_BcN64;EF-eb:9DE#1Id<3^ef,4Z2Z(-1=FL5YD2;(,?<Q\6[.He[Z_d
B\Q7^YbNJ7^bB\VFK+20CNFV\+g?ST5RLg@ZKQ&#6)3_S861J,DE3K+[Zg>_Y40?
CBFMD<@4G\2HFKZMG4-PX:L+SHcK/=N;)O4;5;e?deUCLN=SZ8&1LQU&8+15H9^e
UK8P)_Lc=/W@e1QP=gW<+\?]1>B8eA74IZF9c>(7J(PU78,]dSJNd9Qb?46P<AQ;
ER0(ITU+4:gR+/@E]4cE[QHUC]TA&1SB.L]dXU;HC8g;GG+2g5UJ6N=D50#5]f>M
R3_2g59E3((ZPd;e82-Oc]>(e+/YH>-NDK54aDeUPZYNQ1GE-gc;KfM1PPGY:dCT
><9MSf+P3E8\Wf:5]aU8KBWJTGL:?+:c[g-=DK>)NCB.c_LR1DY^H[NeYfYUOaG>
&,Q@+(31\M.>]OdB;<6Xa](<ZFZ2P>39bgH]#&gf)84(UcO/V[,]c^5FP[ca1HS1
\aWd>6#Ne/W)^PROF^N^#U?>D]Nc2,#,?e[?2RP?TPJS[G?a[?C3L:4+0>\=,Q3E
cgBGJR(Ce-F225/1/R^J\6M&/C#Z5)e2JA[GYbFT]ZN-IOI;#b;c9.,U7a/ONAEG
ZMIHDMDUM>4U8=#)H#fQLJ^J<<^X;_MRQ0ST^DU]:gbc&Kf).TQ6W\6PSY9GG3B_
AY:cNLJ6/B/dRU</#FGMNC]UF;8U;3g7KQ;Z1<fN<^@f,d.I2@-c4@aKY7LA4=g:
G9[YdI+1-CRc<E(GH_M7H-5YNP:Qf6a03+D6-LdW<04::)6dJ>+/;AAbABFL)GMf
VW+VYT=N^;2ST/Ub2\e/;Y>3[LDMcX0UHVIgE7#X=M48?-gG@E#a;E[L8UN:\eNc
3.Z)M3NZa0_\3LH@V=Wa^21G29-V;R=<Af5I4,c9f_G61MA<O4d,-M=)C&@TR=&B
^)K,FY;D)-&\I-F_Z&.DU4d9dLH@JZbHRRF?1IRP1WgK?CH\P[L@e(JKW.(7=]WH
#0MT\NgE^9[X]<,FR#4fgeB0gU<-g@_?X4EGc]\OK[(2/g.N;-.I.HHOa^0MIL>_
A(9\0TT8bK&fd[L[A&#(<+/C1f1G>M(:1D39+==cG<YKd75#C,UZKJa3^.XN(7&U
(3\>]dgf8PD?Y#Cf.(Cg43J=<RS.>#C:21\K\.6=@+V:-X\R3b/HD4#^TS,/I,)Z
=3QRQcXJe9XYZ_d_H:@EGBgL:A+<7?/+U?I>^[gJ/f-XT]ZJMa>FfDTb8K>gb/TV
BLf#UN9HJ,XH-T1,E82DN.Y:KTBK,DZRZQX_,Q1;XFfW#Ke5S.Q@9bM4D4WQ.L/]
JI009R4c)5UaU6).f>6d37\@N5ObY1aaf&FHgOd9-^gB2VJ?Ff&ce,^)OB_LSb.2
D7;3A]H@2O^7.WWcIZE/AU(D>UVb(&Tbcd+OOSVP;gR]4(Y+fHU&Mg;2#D\L,G9J
E:4DERdJU,?CB:Q9b\B-GRJA#8gc<(93X#U?)J(P+BNaY1AYe.IBCIL7Ld/Y9MO_
JX1#]TP;07gLO(=(;UO?MAGWe)A^RZ=QXV2+V7VB-387b6E1FU\8MIB[\X?L7[@U
B]\SOO?YQKU6,e&[?P>5_G3K=c)ZN5RZ4>(;\=R3WH/,b26e+=6<@VY>-D#&@ddR
HUAR1=O/R=B^JaYM_a61G-L/8>X=2/5D-eaQ_@@N+cX&@+(F4(_)50JIM.b4@H4,
A(_WSF0T:J[/bg@QFQFgF>BOD^Ne282aXUPEF[P;U@D->7)PeK/<NWXRMIML0<37
.?+O>^?#eHUdQYZ4>?e\6UABMI3;;3.f/IeGI.&>;1bCC?a<\RcGfS\;P6aCE>XW
>P?TM;=]?9ZL.6WB]R:.Db(:TU=_0,d;.WM<)MC+C[S>G3@2\&NeJ2\^@K_dS_be
c&L;&Tce2W4fA+cAEea[UMH?HMW2D]\Q/H0g=>bd[.Q]f/?e)M#E0ddH\^B=JP..
@MNW])AYEF;1,Y02K^ZTB#A>_)8CIY5&>>eT=GfSf\PN=7C8^<8+:#124#U[YZZ2
_XBNIe9>K]95dYI91F(O4VRc9&]]g4baP9fPI9.[:gI0@?&SBCET(@MGHHYYY7U;
0>P.NY\448=A/48LBZ=8\XDAE,?Lg6HHUAU?)UT#6#&(VXec=19<33:^]XQCPcW(
bcJK^;@?\Y+ET3OEBM+C?G4H:fUQc=,ef2.&O;A)I1>K6e82]fa9(Qa.>VdM9Y#G
><Rg\(;4>U;9;b4TFT3@[UO/dK7[(MJ5BR+9c1N-.2YQYE1]PFI2G7dT8eR3[&&B
Y50.FI7KQ5@@d&4cN..G>DC5QBK/-8&;DAEATbFN.JgZHE&cgL+^2=86I\Zf.&UQ
b?<B3Gb&++[PJ<9LI6JSV>(T-/E9/85UAM#4?L;Z^eD.a5Y-NH)\.Ve(FMBJ9A:g
Ae?R#ac\D#VO0<+LA:9@G.36cb19/KU.,O^;?CO?^)Q,0OV4fYb(+c#EZ[7Y3.HE
)YfF0-PDW4#I_]LMI4cPV3Xb.@_:TK4<WE6L9Nf\N[:X<Xc5)+&E@DX9#<1569[Y
81E<gR6YR1eR7:0-K_2.48cBgG2O9>=7>,fLJUK1U:gfKGc#3\D->JZ?I:ZNQIUb
I_6E+;8bMIT[85FM53HR?/FAMc?M+M@1.TfC;-+-N:8g]\WeU/#G;Nb=I]LWc[F^
M#1=>6<HZ9D,0+4GY,d+0]6/]I0+J8b++YYST?-O+G#4+)a&4QR,CG\^aQT]8)ZT
&_Y5Q6@GR7>[I)IbJ\dZ>\SLRV)OTZ<Z#H(2[=cb#2[Z2/4(aK:DeV&TZ4DJ2MNK
<_IIBQe5\\_#/F_Fc_97fC^LW?Z01YL.V:JP(#5aV)+25E84<4J9EQ_18a7fJ(P&
\J]ef;4ege:,41JPW=A<9dER[E,+)S++J2VL_dY@?9<cO&,H^C@#M&UY?,Z1<SXg
_EJC02)e337=989+?7@MO28[9TEPc_ZJ/6&bLE^Xa-WQeQN3V9@(eb6/=RG;3LM1
P?]/4_\/\4.S\83ee)<\UaY55M1>_8W[#CB,]#;?HEYY_:MBMe.:V8X5_;WK0/0\
Y9bfO;L2B^U&fZ[2VO#;H4L:Y&/\RM)X<233ebG^02ZFLdS[g+JQ&^Z/>(:.3,)Y
5HFOR3+F#H&-g,;\91JDC4dCb09GD9XTB8)&UNg^4SVD0S(a21T:IB-f7.6MP=RD
DLMNI(g+G34L^IT@>6_V<)B3af/7C\ZTC<LA-T0RRV?/2WaQ?^SI)\dSZ2bY@3dR
9SHEGPeXfSfCVA^31a5Q;^7.LL7AQ0N)#Q^gA)ACU5/4TWGL2A#=I)M.Y8\GQB(R
W-Kc7F)B/#DQX\e0#Y:8c3.V@5O\._IOXQO?BD^,++3<EWK#PGT#^O)>ac<7gc<J
3+FIdC+7NPG(J<V&;/&]M[E<O<.fE^S->4PgZ&aS4F82TTF-+;+BB_U&e^DeSJef
b/ZWU-WgD/+S&DKBB;FULGC(\A\W8?)HJFRMFOUMd:=J6Y@>L]#F^3)2D](^O#=B
1Ze1<CRGZ#7.QZ#dZ>F(2IPM=VQdO)0a@?YA[UbdV6O<>@[2f]?;HDg0S#c(8B9a
F9DM_D)98:GJ(FY6,NZ/>Q+&^_Y(Q]LWRG]7+G(GT#K&31[K+^LYN\SN0[f[]FG-
;=c/^<e3SO,YC8;-3B2SeR,H0A8@e\CJ;I;dXXF-SCX>OD1W9^<0f>eM(74cgd5.
(aOLMQEM]FX6_SH]6+.<a=Y?9:KdJ)KAGbD/cPS=5?Z^#[3Ud^OG9HV)<&(10<YF
@a3O6afKTa6]]XQXe&A(7?/C&.;?9F9bT-4ZUI:L;L/3HgdI;F9_Gf4.e,[;O1NS
)H-<P=T#.W;[GYM8a=4KQAc3B3)/:H9TUT?e1T.X;Z^\E:#@_368>#b(\J9<8NeY
bc@MKf5fEgM27&E]+G?WH\84J]_S7YgK:R=19UDbdJA^.QaHIc^W?bd6c-YM(0FL
f2.2WQ@YY+;6SCFSDAD7O,J)2TU7^fG38FbcK(3XMW07_BRddQ#ff#cL0bBN;cY#
DELTg,/5<AUCP]Z\/GgAU<,LfPd6RH^34K&BT4?9#IW@@7P@_YCKU8L#CO7Za4A?
490Ab@]9QAbGQ4JN461a5;Fb7W:_B0(#C&d6.A7@eC9KKP5g/8TMHC7dJ@TaJE1W
J2FR5GRODO(:d/1O[E61_aDg:V2RSOR+ceA9DJ-A;=9G-d/_B>69Ha+0Z9M62T<D
W_8X?4c;aO-^M#^0Z+,>BM813f)Q5Q#W)7aXB\E?V:_97S/._7XM&DX>FEZQTWVL
():2(:5[Y[\^,gL,<,PNbMJg:()E24:_d],]][F4-)HKM=^BGX9MZ1^D^,;BdUeF
>2SG8#eI.UPeVENLL-SJ+P)8-CX.(EO>H)\Y(\K+2I9=WAT7GL6]IGIE=</CLb;&
>Wb#-7CLQc&P=9+B]<ABcY+JG=Z_C@\9#YS8KM8[2=aOHA1D_@:6WB?,9@MT;J?D
V(W#:,R?UB1SD?PcIAW1)CBHbB0<G7VX[[1^@6WgX#g5XE]._GXS9SU5\KCO0fC[
4/R,BTJD@Ub<.>HDY7-d]K/JK@BH^_DbS^Jb8CC2-?6[&Y\8Z4UWM]dYG(P@,d88
LEUK&\>/,OY<b:b\1;A[b:YJ:IK4FPXA;Vf;YUC&D(:1AEN88:g&]^Y)-<S[VbcU
=faB]BRW6PcV(aMd=)M3._CKU5N(^df-6L@>>9[5O[TVeL=<FZU:WS,e<(ROP[Q1
Mc^NY<ESZVSg2b<#[0@=W76+](),HJAAG/@:9@K\1WF^GP#L1c1,3O>\T@V9aO;#
=^X(Y/R;@94,&8U6,?QcN4I>B7])eOcT=FPVC8<#/&\RbY2P.N&3@ZW(\-gI.H4P
\:fAZ/>JB_LZcPa,F\ZbP_5KGOJ4_9bAd_ffYGH?#d96WRR;Z@;bSRL<J].YV)?F
0;?-G9X(-O>;(_b3MgU3A>5#L]PMfdF5=<MEFK(/IaNX+GFf&LTWIGK:L2)@1_53
>[WeDO2FH]QTb.A&]D#X[D&0YTM8]L4Q@<4f?TQ1X;5\dTPQ+J[Hc8-L0P:X]_7G
IMLf4d>d(e8ZE<CTN_G>UYe.3FMaETJ3(:B4;@.dO-6]g9>30UEO7X1T^?=DaA\?
F#=bfB+[8?=\cP\;,KF,5BH?OXW2.8cX477#bLd3E&-HAG>2#N:CNa4Me/N[f>]L
-NO#>I-N1(/3264bg5J#GY[(7\\Q0cZ)f6I?;e#9T42a4d0OH@<WZN+[af(/J,1d
6a<IQ06D6.1^DALY?0;<?2,.THE=^7>:MON.NP13E-5=c0OP[3M),V@-#<]IJL#\
;IWa+<3cPMI-,CFO\T#9UE\b37#EV-c50=B#8@,bge6^E6W#0@(:HeGQ/P2<3M94
/3HB?g4O8c(@XgW^e;=(_M2d:@gX&JD1.S/f&5eXD4Y]2Yg9_Y[>R5P8JGVDVe1)
ZdKa@H+)(._24M83,#e8.Rca1>);,:AdJ4]:.#GcIQ)#8gPSfTcM9&e)Q#5+^=55
=R3TBV#0-RB_/Ne>0X))=M;85YfCS=GL>g\.>N;3UOXC@2RV?:V)PD:G?=++@9&N
?XA@O?X[4F?([f.&4EC0GM=IMNMZ>G/0+J<#_QQZCOSXZSY#ZF@2.F,G>\V1(LQ9
a:U<ge6?/6HN-GT9Haa[;\36>R;-QL0.VE?QNZ,aaeRS-433V9YB,#ePd>F,-5HH
,)HW&Eg2YO@LPXMSPFZJ/e4MB/e3afL8U(O-:.B79G7)F9L+ee+Q8\98@TMW.--<
P[KQ?WZZH/NBY++>b4;XO007(L?YDF_b#X>Te#c(-XTfBbEg1715Rg1.AZ7V4:MM
PGHWGVb^g,FQ+Q/5KBg-KMb[-_K+c79(@/ULEY+[:fA20\]-I#04K<fS1Ifa@3:d
0e5T3=)\S.1AZ2\Q6Q^]=Xa28]5[)WI>>AY0CS0P3bVN3]XaEWOd#QC.GL0c6HP-
(M?=6OJ:+2REC7>P5dRQcfgdU<DB>RM[:QBYACW77-[9@7NaVFDNI#+g][LLZ-+O
]>;/LRLb4/)MI-Gb;cX7<g-(>CB1O=13I6Z81H4aH2I+O)S90=-3Y=T<(7[W9BSW
B7HI5>018+3,=eO5^@U55YTH?de6D84#4efXT.dO>dfDFe]QLbWSVa3QSK<U2<;#
b@K]1R_8^E4f#]P_,KS[W\@ZXU59R4KPJB2FJ&S5M(6b.?]@AB@1[GF+;?U3KX3G
4OG1DL&1;JWP&M_fEDK@LI#9-NJW8N?P]4Jbe2P+Oa<\TXZe&DgO]A]H?=.80(=F
X/IFJX_O(Y(=J:[(==UF4_(+PCVge48AdGGK7AXI+U2PC>HO,da+M_Gg\d49)dVO
LXRHA-79KR+OH\PEK_Q;e^>?W>(J;R3+VO-.gQC&Q6=IO0J44W0+f6;F87QFIBQR
\XR8M-aIB)d_X4(-@:1W5UBQ0TIbR_/dR3d3c\Yf8^PL&/O;IND(_-5JH20Y1F0c
LV+dC5bBEK9?&L]01B3?@2bK320_OOaee@VF[TO9bYY(+W9IY_43&bR?\(:>[03Q
(CB,P9gYb5Hf<H-O>0eR7_1d7,Obc2.2,BbQSUF)cUFQbS;?WJFL<1I1NH?CcbP@
1VIN5=Ye:YJ_-+F1RCW4B#WH/WI@4CH@;CbAC50,(1f2@GeZbQ3X87I7I]XaE&?c
G?C9BMQQeb(\/Z<WDE(Z9H52.LJ=-TZN(MUP=4[?a97F^,X#0P=B3eWa??e::]J)
[NMN,>TZT,Yfg31G@UWJJ\?LXJC5/PM:T\S2,7M9RWB],^)^6#081]5dCdV[PW6f
0#<(FP;[[RCDAPZ5H?<I]I^^(ab)<U6&fDF0F8T?KTa@R1WG(7^^[ZPG,-bS@H2<
X_QEdb3e?e0=2^?#DA[R9RN>b@8Q6@915U#\3ZFHMaPU<VIX7E1]G>:(4?d[]IPT
^@.Z>+gCK)+K:@C1I6:6=OCLE7/SG-:aC3J,Tf>5Rd<W/&HX.VM;#;V9@?=8+9Rc
f7Xd>/WH6cV<J,EQd]\JLV<ZT??220GB-\_.9Gd)8M\B[OfL?Ub&GW..GG+1Vd+6
7@g)9;(_3VJ#/;:T_2_#S]..GcVQ)e;MZ&21R?J?-E73B4AQ#L/9I9O\Z;C8Y^[J
6&/_f\K.9:7[49)VC)(_4X<b<-gcOH>>Z9(YJQYW&bN7TR(V(2?Mgd>BX?H:Y-ZT
2aBVES2=fY53A+AEQUCC(\f>K>Z=--28\TTaO.2>:>AYbK<Y7QKHTgU=?7Xf5dbU
TH^+Q^UTI,>#f/7C/SA@Q9]AQRY0UP)FZ,05.#eDD(P[0VaLPF\c?-=c]QX=D.O;
<STP4=BC<14Z.@A\LY?a-8Y:2XD2,([MYWY.(H(Gg>414Ae<G]9J@<g<9B_5\BTD
0=SBeH7faP+W3QR4L&+8UZN2BA=#?OMD:<-/bFQ6N7MKPO>f:Y13ASOd@VXOeb<_
)?>YPB?e&UOW,)C\fD;d0O_<L,QN((R:7BaP4I_8^CG@c1/PJ0<;Q\D>-F=.FI:8
O]=IX\XQP:1AB>c+HD(9?=/g,_3SdR<c3:.c2QTg:I0YQ1N:FMCc]5JG_c51;4_S
R:>7ZQ?HSIS>+8b#[PJRJFCM;VAScA@aH^V.)eRJXTL/AZ?KN3eQ]FYK0a:-1:MN
_.S4+X^)O1A<KQ0ME61_,M65G:P\:SA^cAKNHEB0L\CST.GZAD]Y&dRDHZ?Sff:[
NcU07IP@0/eb/;WZ+NZX60NZ-AR,P4f9dY4;;-4/G8>9cHcV_bA0#b70D5^?VB7Q
JR_#Z[^R1M0VeRNFT.,ZB,?.B63[7+W(KLN;.c]bQ6.a?O2-eNAB>>WgG?FeUXdb
d2H<<E3PWA03e;FUf(H2:3?F3ZK8:L@deF9VEL2FXI7#-Lf>&8IK&\.Z\M?S2BOR
V>D5<a:Z?<);&KXPE<aE<SN,F(60HWU))N^1BX)GC[K3UGgKAf6A\/;F;Q4>FZRV
YMTe^)ZWAAH0QYZ:-c(R^KK[V_6G9:_Za>YPUMWHc<OCWLI<D^M78/3(U<3,TQX6
K19E^6e1f\V<QRWU6#N_#+[NgA?)X\(@G7VRV,(7++#e\b9HB=93ME[Ba(EAW9;7
IXWQADO-][W>CfCV(>ER__40W&,#MO3JR:&aa#_5LQIfGHDQ@;/3C)CC7)bXQ6Rb
QFd;=2]e^#;H@Xa0S+:MRUWMc:5UJAP9C^3+K?XA;-.UHeD<;M=0)>c5NYd.WPOH
N(bQ4>;N4;e^8S<]X?a-Z)80_,KcJ<=MUFc^(,-<aJ5<IaT1_SYS(QM?)U4Y._4c
.L1ST6QZ.b<2J(SbE8I9Y5R>\cKEE-W-#Vg\FSWMJGf1AEdR##cK3Eaf\_6>1)ZY
#+UI^>:CBcgcV-0(P:)0N0O26@PT+R9Y4.K8&J#M2]6E_]6R)AfR#47__E+3PeHX
7.?EbYW>ZVK##C+gP8T//HCA[HD)AI58DG[B^\U,d6@J=4+ET6I&^&>B961a<?&d
0F?cbaED0dV?1XF,b:UJ1&_&^9R-_1;a[,.1:LMcbO4S5)@,Cf&WTTaQ2##6^=N7
N>@A7bS1=0=99/;gN;ZZFMB>NV=MZMG^<9L3NVD^ON\X)DffSJ8EC06-#\OX=Z[6
A<TV]N@,J79ZWASMUB(7.5)MJCBVa>#d309&/_VcLSOS@;/-Ice:E.4_dBQB;CG1
XAU,H+[)e\:14=a?8I\ZV7LWJ=T=(ecGSDMCK<gQL;eb_>,#3[O6KS3T=Q[,b/4]
MJ1A-[aO3bL^:#73C?3#f/BUJES=JP/_)gdC63Y[(UZ9N3cM35&]S0.W;+Bgc1+E
dPVb+04cE(9ZJd7958Y=Y\J\^?R&+(geMa-_DfU6O?::;?Q8=0D<f5O;=2>b2#TI
c=(&c8TGY<U2XX,.;(_LVe^[#ATNR?U]c<35U6Y.bK7#gU<;TW2+AG;EM&N)-4F^
\gS,ESC-7\Pdg@4;1Q3_ESF&dEQP\TZKP<GE1)IP<I]M.GX=B?@\Q6gX:++JfB3O
\N>d9FWI-.Jg&),^&>W7==5WZ,bRB<LM<,TZ0FH)KP]Z69J(OEa1MRLJ__:C_1_(
.(FOI:-&GL=&6(a+V.1/]WUT50Z]XGP3a6cfHXOfA9=\7S9GDMHgL[/9cN.6Z(7)
6?&+R:.XP@1@^S:d^11P^ZENDW7^GeRb&).=M\?[54>-QIW1YU24^8OF\7N-,E^:
6Mb\<J6ATV.;)]6:dbW<Mc)L/SR8GA2B)S>T\(47<:dW=JNQABRfJDTSIZ5d)]Z3
)PU>WX-EUfeaT.cH4]cNXd/>8FT8@.W2??c#4f/GI2:FaEP>ND60D5+)LQZ>7a]W
XV-D)\>OLNXVMbL2(X9,35?Y>?[P>F\5LcPSQcI=MOFA48A,:7DWB,VP#b4d\b(X
Yc##B6Y[0Q#;Q.P/[L^YY@D#WMaTH?J=b\2\86GcBCR;YX0d8-NSfDf3I+-_c<>A
>b:V&1M1<7?/?)0G9AVA3ZU->-.5-_0=3/SePMYXe(Y1UeD]48(1OFc51fNA8V_,
U4Y3D^8+A-\;4_KbJTdV>G3C<X2a6/T[21Rc]5L)ZXbHaHU^:7=SeZ;d@,7)5-AK
9(]ML@IS<b_f9:U^VQ\dDdQMP#J_6V<E5b8RgH[Zbge0:?JCa67@-+X-/X<GOR9b
IKYf>8.N9.a?C[/g2?_Y<,-a0<NL_JGWHeeQU6]b;afV<bIH48JN.e1\CMe.McZb
P[[L/cee\+W(2NO/[5]N(-[cYOIbVK1f<$
`endprotected


`endif // GUARD_SVT_AXI_SYSTEM_MONITOR_VMM_SV


