
`ifndef GUARD_SVT_AXI_SLAVE_CMD_ASSISTANT_UVM_SV
`define GUARD_SVT_AXI_SLAVE_CMD_ASSISTANT_UVM_SV

// =============================================================================
/**
 * Extends the base UVM command assistant to customize it for the AXI Slave
 * Driver.
 */
class svt_axi_slave_cmd_assistant extends svt_uvm_cmd_assistant;

`protected
Mg1Y50;&.BKVe3Z&fZ0e,.15</4Z,IWP4_#I2VT6f>;(5PF2?<C>/)d=FIVE5G[N
AF1V8J<H#RKCX#;XB2<??ZZ;K#6JDOH4YVK0E^GK\>g./)Y-LEQA1DZQYKNc.H\U
#)3J_8.ce0FcGU=5[5f81RbQ@HJgDWK;L[H(SQXfg<(X;>EbLdKa@6]QH\[:V?^+
Zd4&N&MY5=A[5XLR8C;YA@O;IYK+<N0N3N7g5=/\eZH&H-KWOD@:YWbgB\N[W_UZ
O)\Kb_R+=0=#cTZMEFSYEVXSOe?VLE0]D7:2A\E4feIfA+WZX(6aTA#)XAZbP9WO
RY\<,TX81:SPW8YF(BgH?#9[GK1+-d#V1G@32)c58<58_@3983N+M_2Y8<C3?P<_
,;1K5FVT;1&;6?(O1bH-8,;UAPA@LIE:0ESFLYL?DFNGd_OM3f]IVRZXfCgbL@TE
Wa<<61KP\57/c@:IEE0]IY]-LXb)/c7+YZ828PD:8f/O6V7Uab>-B96F^_[?&XWe
\6fcH5+&-KB\.0/KXKWZKLMQ.S.BP=3]gNO&B38aUG#TD_G7UcYWJ9X3=WEH)5\>
1ZQOgP3dRF=FUJV<7-FH,RRXF/<V6HGD;WXG7b069Y@Q(Z;__JQJaA)2ff9QfNa=
E5BX(A:_YG&5I#]/XD>e^a[I,&@@^UCDV]WM_/H04GASQ2d60LZ(915d(-6#SDUW
:GE.RGN<:C/OI:A@/WXaBb<.QCH9SWJ.=QZgV+>G77Y/(LS)MT]DaFL-4KY7Bg58
d_X=260/04c#gT,.V]NAA8Q0PJ7?;)3]Q7XO2RQ8&;a8[?G1(.HcVbNg5FaeD\0P
b&X))c?cNNc:R/@//IbH1CQ08$
`endprotected


endclass

`protected
IF;8M;^O&<MAKMf-1[;-N,TH=&E:7Ld6^aFd,>eW?dN<K,[fd,Ka0)V:6THMFYL8
QePB4079A:S@.8[E&9UPBg:I)1bJ/>BRJJ+BX2>=#V+())BX/U=a9c@-G=-dKRZX
3Z1Ra9e].)Yf(U3I:I03QL^@4I8W>8:03U3=?Hg3=?/aag,I^DB=]INY;\b/LNJC
XVWT,fge4:I[;+1TZ_bgDG^V[^]_D>L[Mb)#D#4:FFOgd:2-(c_>7_\LFBJe5V7?
Bf7+B]0IgB\-4ZEMPR(M@P@H?P9J@8LZBF\LD;1dSDcFDA&BIA]5V1&b[D,=F/bR
>BKXQQ6Q>bZ(HHN@5VUaE_0f<X.C=:&I7bO:QSgKW3bO8((/-GG=W,=<EIKAQ@03
Y&JfHM=#A7BCMCaN0/cPVW(eac1d7[-c+Q]cH13K==d4@eI&E+@,cNAID5NRGb:=
g+^A;UO:I#cJbWF6J,05Le,d&FWG+cb\&gdMb-6BLW7F^;IGX/IPS?;[6>DZVZ]?
3@:D41\I[O&V#TI?aEO5\/^SJYN0WIRf.)76=LI@QX\eYVH3Y3dWM>Ya#>Nf5]9_
C0KTQCBNEeCTU\70]O[a=+EOH3J?)(/&]R8Z]#a/0e+C^SDJYRJd=(ZIAbW.55?^
\EX&3]/3c(,=T&BTZ;SMT2Y2)#SOEOSJ)W.^:9ZFKTcR,<IC9.R^=WDXJ0&T+1S:
HMGJ\D__M1[KM#EGS[P82@:V=,]E56H4G=.>M0=EVb,VJcHPABcZ5FFVd&Dd7(8Z
c>O<?>8fM+Fd4^/,9LF2O:d[KAA/>X5LS[(cc5N[UfS0dRbU)@]Q/Kc32H6bBH.b
6GZ__b/V2&?Qe7DaFMAX)QFf09d2[6K-G^H]XANd_2DG7?O&,Vc/+?2C<4DBTW&[
FJ^0_/[a8),39D:37eC]ZeS6aHJRW8W<bb[LRN6:d,[FfS?LSEIC-F_2BgcY1b/,
IWX_7#+_XD?<,J;92NgTLgP@MAfT.2O-YCgXb<c;YEJd()]e8Dc(DB^d4T<d[\O+
2Pe_1^E#1]Z(TU&T[W@0\K(#e5C2;(E&2g#d3G/=#0W1(TbRKGJ59/@C,c=e41YX
<5@d1Q@8cbB<Z>V-NU=Rc?Kb6Va;#G[42@[QeeGKV@g9FA6VTb>@.)@Y,DSN]Ug6
X1K1bDJY.2R^X.(QbNPWcQV0cZ?&YZYGZaVR(^8DD@JY0CNLR/:F#V;N1D,DT29S
DcOXa17(O8CG8;\,PZBTa,3c.c3c@;>X[<P>=FLXb;?SMR?J-N.#-YN(AZcVDWR/
9RRFUa4P?1T[:4FWO-3(>7\6T22A)_#\_gEcS/<Ec?9MVX[UTH18=DK]W<((6,aL
E9P248_54e:V?J]BB@&D\PL8f),H@,A/XZb53cNe=GHbT(G=.dYH0g@/N@4e&J^Q
WUEI#9]]J_E[2^g<ZT^3<Lc75DNUB)\#BC;=a,R=C3G?_<cU/N2Wd7K<VC8[;R2J
=G#.3g_4ND&g8OE:R5#UVggNH]N[@;TT5=3Bc=b[XO5,d1_Q=Ig/X,R4cML9Y_CQ
S@_#6KO0@3?T(\eFT8QO#?<+]^@VQ6HKgR7HZGK1K5W,@fUH34(d0_#H8Q4YJ\#C
/Yg-820JXEYa[JMW[<T/M<V^f]cT;Df&-+W^7g>M5R+>RZN+8^&.VR4C,NM/\,;R
,]R:9&>J,)Z.:EHK+(FDU4W\I#XF=A:\FQXYQLa-8N;+]])++@36,CeN[/6?cBJY
?<;B\JSYHNTH8aX[JUbW_KCS=gAN<Fb)QGLU/+R<V6(-(39eZ6Wf<E4+6S^(a9+^Q$
`endprotected


`endif // GUARD_SVT_AXI_SLAVE_CMD_ASSISTANT_UVM_SV
