
`ifndef GUARD_SVT_APB_SLAVE_MONITOR_CALLBACK_SV
`define GUARD_SVT_APB_SLAVE_MONITOR_CALLBACK_SV

/**
 *  System monitor callback class contains the callback methods called by the
 *  system monitor component.
 */
`ifdef SVT_VMM_TECHNOLOGY
class svt_apb_slave_monitor_callback extends svt_xactor_callbacks;
`else
class svt_apb_slave_monitor_callback extends svt_callback;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_apb_slave_monitor_callback");
`endif

//vcs_vip_protect
`protected
H;_JZ)/Z-fA;:2+\=UYOOEc)N^@F:8C9KdQ#I^GD[I=73E/CX9Y8.(M-W_:^-FWY
JMa?&AD080aUf/a0N8gG_WfVYS<:JX.UZfH[Na>O_\B@ITXS&2Xe4:I,\TdA^KB=
X-,]F6)]W]N>S6bIO^9(TI&OcI,TMQUL</PJA(_(9EJ?B1JHdDG_UHWe_<YQK&6S
&4\&V=E=Yc@Le>QA#SW^YK20<I=(<H&J5>HGE2a]3FXW2gHBeQ?2E9E1<2#e_QV[
H=3LLf6PUcF.?>bE&-d#dQQ</1HT+1,WOgBICYd@9aTDG(MS9[S<9dJ(JgC,[=RO
ERTY0YC_Q^KEF=KQbZA]Z(J]].2D#&N3M6Gc\?d,:CDLSKIYO[>^CM[V@M:_4A3O
/-GW\=K[#_DRVV9FQ>f)M(LKKS.FJ>[V_U6dYUc<SIGE:a[-gX<5)U3IaQ=(aF;@
65>&DOIP@_Z,G,+Bbdg43(.JZ\Ca^fJU8&;)E#JVHRZAS_)Tc/Z?E>MUJ7HVGVZ?
RM77@68Z()aAP&;?(FAF69Y0R59dcI<O>c=cCQdX5?ZG2d?G1:G+XUP-=Q1Lg7TD
A&)VE@2^^)X5UW2QD[7DG,IK></&L1YI;9gCN0\A9X/5@25K>#/Y_:5O88W4ZXJ#
<G2bf0eK5;H2HIN,9Te?+2;^QN.A[a&)N@9GG2F@O?:/;d33dYT5C/4UFVLP]D<+
4,6NSBc<8;OWVKB(OEGDLMT/+/L2W&[g_G.03N[Tb;K-+C0O=c@F438_A4OZO7BG
F2V#22;O1P4O>dZ3Af6B=\0SA9S4(:<U/LM(KI@U8X^+]+LKdD9]90KLROX?_X-d
g/=[+)GH>@YEJA2]SGbCeQJZ[.^YKC2(QQ,c?O8J]g\dXR07ZJb]#]81^J_]-W,c
Cd\G),MKQ06SX7T[O(,Ce_4>\-=L_Qe&f(HLNKCb,EHH3:C//T/]-c?5:2+@Jf-N
/;?eCb9;NRX;]F)OVJ#T^L-2O8[cW8&T8T<,],aO[,8T<K26X;E^1(9I,)U8=9YW
J=P+R?OF-T?7a02:a]_@_144f@/=(.Q)=26_f1&\^IT4?SgIC;,bc@[,/#[F_d_d
7XPHULcC\.NWd8VcRe.MBWSOd;SPBMAEdWg#E(JY\1JT;?^2VROgY8O5QYb.BJ^R
X\NH?dc(_(X)>;.-+<0?[<FI>BV:?7:N/K8CVK14-T2If\e^J9cYOg?-_.4H6cE5
EJL?S:bG5J;+^U2LXcdIZOUgWZ+(8DR2.9E,9S66N3VPK421YKg]S\S>=\QCK?(X
3T=@8L<DN]>eI;AO]d8;U2C76;6X:N2d:D8D7?fA_B44b<I)5;&e-1;5.?+__/,Q
6]3<b.&V(@#ROG_<H?@D<Q5EF>P(bV;J^Q=_N_>VE,@U>8FS:Ha<NX0?RUR4I50C
0R5Z;_Q2=8/D.0E??[P[O&4a@E_a;S[3gSN+(380]JPMR?BTKGF\AYIG6=I0GA#C
?1+(__7TX-G9IS;VeQ0c)G@U;;(P<481Y+c>e^[A+[<RR(,@HGbSgY6HWa8EPTb5
.-T3g97VGT2[(H=-O<RT,2b^]V_IM)3LU5Kcf>DM:)VFV3QC9@26gT./@-1c4Dc(
BR8(X3BEQX1L,F[_8QB>O^7:_>XI<F-dbY6397(XX-W<WU<1UYVAJUR@]-D-d^TK
Za__=6^g5;G2[5@@UBd1R:aMVYH5C^:R@W_eV4_AaX9)XK5gBP?3[E1eXD([CMZ2
6\8.I4]4]PQ-edL:C[JHYWR[bCc1/,;21Y1(V)PNQ7<\b?NS#HI5R:I_Wcd9d-#_
95..ZBE#ZT)A7.g>=0G5fFV(OTXSJ9^&H#]6F#O(;LAcCe)D=6BUa:\)f+J_5f@X
8H.B[@fDIKMHH:KJSCag=L:f<G3Kf7.9_,=U:D,cfCb:>X#c;J1N&^Tb8X<@N6ML
+UfdM9W#_6HFO?NY>S[f;F:E\#g<S;K6d/D?Ja8T,@-Q2NQAQ+Cb1@-94?JaT?::
&/QA)^d/-.]T=&B0F_)d]_H8:L8MC=@?^14B0EbTPS5cJ?W:a>2)]8.OXe_G^QN@
/O7<,Z>2-aa2/4eD>2f8AbAS^FS2cWP&/+LYObN#S1cTDO/7-\d(05:=RNX\g/J4
JB1SZ6=VMM?:>EG3@^Of<La/O.(K9?G-A3gPL\&6NQW]a\LL=T5:IBB<2ISg7cD:
AFIbT78KB/^/bU0E]#4<VZL4a)0H-G-OR5A:SRcReU?P?UDX,5^XDOTJRMOU]#<Y
),><F43T-fdCQfVJK9SITRg7e6+]acTbM>M96TYJ^=,f>G)3gOdDgRT#be8WP8Zd
1g9e4Pg01d/NSaSa[@7^.5W2<F@_5gJW@5\,ESAM.E/eKDAF2<W6,+3L\IUG?BX_
95],H3,eOaYN/>MH8:1ROV=W0?P_/TP:YNLdC76>fN6IfE&MUO\>SA@eXcLI:Z=F
6-<I2;PB_NG@3P?cgd87CSH+@:TIDW-JY9D1&3,4#I+CZ,dP8ba@4-H?+dA@5?W?
F2fVF>/+L<CMEB,E\<Xa1ZGJ3MZGUZ3NcCWNYRCABF,_@OQRa:LTCIXb8.?#I9eT
&#=P22Le.\eCRAA<^+@U/70SX?_L:67H?ABZ2aXR@LK_;:fHWE&64@bL/_VZDRP_
e-TFITTT<ARE@9K-693^897XTG@g61c&;BSIMW+<JEaY2/(8;f/gMVE(<H7b3T>@
;V]0AUPCc;aC\6>G=OA\>:f3A]?<)HK(#/?Y3\RL=(5dDMNdU&\5DLQ),<e<.KPS
,MJB@-fQ]:^P,,]9(^@;8L?0#D24J\VM@LFacec8a_HGK,dJRMa^JZb@7]MXME4_
@N\VFQ18_a@>G?)cMe+9Fb-WA^^J,MP?RXbHabUN,/^a2TB[c0B-P09EXG_MRUU8
DcgJ#;eCZc^Zg)6Z&(0;E_&2K,g-_./#8UgIS4E/HcK(&C[I;RgRZJ&g^aY2,\SW
H&4-CE>:]Z69d[U@(,YU.3:Xd6YS4]a\J2@3/(W.6M&EK\(9aH&(P:8BBK)&<N11
Fb</-B:EFBXD5S>DE]+g0bO,7G0e.V]f)bPO)W:0Q9#bV2^BgAF\:\J@0HM&T37F
RGW[U]FP/a-f3K,#1&<FNgJ].(69KbJD)Q(7.1C^GS,QbT;ZgaFLC9>8YL#R]Z[X
+G,7Z7fP(MDK#U6E?.:LIJ-TQ52c//1,:5J:=2WA3\QO#VeJ?P,/H;NXQ[-RP5Sa
8NAP[2..-_/22I35<?eF87A0?83-+4Y<(G8OLS6K;Aa7DT07f95_32N?dB\:62KW
Wc]c0(4EW;YRDU+f,<^-O>JfDgN=JR8gMK5:5#F1X<2[#2.(9\>#LD.053&Ic&OO
Z+YBE0^;7^_A(MWZP\H=[^:/.fFTHBYZ,)--?PD9KN3L7If&>4OR#G9\G0]H#,)?
M(FEaE>+PV=;[Z5-Dc[06GF1cE;IBJ>V#BFZ5A@<ZPWf4A7&NVV9LOaQ18[SAL\&
/X,/P+P8GJYc+#-,1cFZSbSdIV15CMJ0MU\V8QZZ.IX/;Gf8XW@ESf&fc9[Q#M@)
:FPV#CVQ?CZZ.KI60=0B-J\#^42^&0c;8;DSg,[;M;(59A(1ZcVI?72GLa2SM2Q(
#QJBC]?(IWQ06,2+>+1HWS(Rg&RTcH0]9+@U2DFCf;2:GG]S5L@7\:EYG(B?+ERU
BDQ:O[HM):V+D;)B9>MVXLb6SF&)\2<3Y(OJ[)/YNegM(6@R;.f\(JZ[1aaP#RE8
2LaUFZ8UVO1L08X6.Kb>S-.aC):L96P\?baEOR27G=NS#VQW5A?VL;52WWUdN&M6
O-,_XI:WQ&gdYP-WI0a45dV?XLT9YB)(.F\467]PeY(I.cWM_gI_D<86T?Mc=O^B
^IPGO3EH.4H+/VW2/X[DTB&H3)5eW@g=(DHE\,T9R+Z9/TOLSaW)72;UCf8@:W4@
E^;<#1F6e4?Db>)gQ&Q^\gg9CJ49La5P7WK8P-fF7X[b[PPXP(@.KG]fXbM5^d(-
Z4[9\c^9(AY@P?&:II,8,L?_L<IB/gb9g)=9,b,bb(A3deQQE9,F_.(L_C>ARfT2
13E-ae\TJVc/ID(4[a[SaP\N4.L3M[1.QF\^Y]fA,(JO9HaZbWV=\/;EU(RE_NQ2
S&f.(&eZeKA>2CJT/CVSLM8EJ-4CUFZR/@WD287^bB8URZ[,R8J,&6c4A4[Sg;[P
P31#L6:bUgIU>YXAA1M6+8C(_7gZ;bCV<-&^-0ST\&TDP,8ET?5.@UdGfYWI\U7/
^WOMYI9VT)#&II+,(L4RIJJ0cgA34Z>SeXU08;cQXT)(.TMYD8]b3ff48J,,DQ/;
GdI#,H]/OBcAc5e^N&BfNT^]c)<0]6CLGcg[#>.H)LFVE^T=ScKgUUWO:LSf-4#e
c3/YQX:L?[)X;4-gEMC::&f:P>FNHP8d];[=UQg9Y^<?7-&4?]DDY<d0QXT<eQ^.
UU)Q89b<a^EO=.C7gG2H?&0A]agK.Ga^/^ee7J7f:]R\7YbH],<2PY#[X9G1b-RN
=HRfAeZTV-b+\(--^DPdFgfW>F+OCfH\G6U+\.ZGM@KQ7(O.(L)g/K^72#5-eZG)
=@1P+>Q\>]-PM;aC\N+X(]0NP^CHa)PZ5GB0_<8_Of;V7,C@LP[L-/g41CFYd/C^
.#@ED_FUOK8LPVSd7QeA3UF.;b,Y1(AM_-F4EZ)11If[@DXKF+__V5DRF>18&Q7f
d+=e<Wf[X86#IMW(&QO)7>)\,PLUdCBT2OB_GV&0_T[=_#L?)JQ<WQ)_LZg+?<]2
I-b_\YA?#OU@LY(H/OgM(>85b&^@6&Yg>8_7dN#[\X)7e>>@)[&)\7P<aQV[,OWJ
ZC<X5/S<+4V\+(@=YFW9f.bg&;ZT69B>bLe=QY7?5D:B>M9Z^D3Y\JgRQMT990H=
N\\7gD,JC80\Q\H10dU>_d[4cgEYf.RQI-7<2Y9;0aP#S&a.9f(8[#0CE6NYDBd6
YW5?2^D4S6cOOcV/0M[YF0G\#<g5()K]B_.GJd7OSHfTGgM8[4SM-08Q6cG1a7/8
bE,BGaBSEcY,,S4_8\N)\)V^FN\cV7LN9,FI7I60a9OR^?.WdNI5?1-X6A?_OYK?
NMQQG-EIIB(?\RY>@&dAI=RY98TNb.)&D8NLKa],DOXKg=]M;Q;B=IE+^@PgO<PK
d>g)1,1XX1-5]Qf9)gP+b0J9S_Oc9c/#7eTXCdPW[6MMR9(TH4^8O_I/XdB4V^g\
0YT;GY7B7cR1DDB<fYRaGTSIK=C&JP3?;=&70b=fFf0RF3gMe&KSG&IQX;<LSS3G
W0DeOc>:?<#>>+;?6[;\EA647H15RBJI?JBCXQKXLK8c1M8/ERK,[SH?LL_:CF)W
<>P:9d846F@CM^3K:HP^SAA3gH?2J\D@I&4EGI55LV+2@OFNc6U7B],Z/2Q#)YeN
EK9>gYd6L?=R]Fc]E&0E]JaebY_Cd)-FcW90[:(GPH,).7J)),U3../gB2JR>T6U
Y_;2LZ-8<R7<6KU+613D;A&&OAbF@AcXMg@SJG?.^>cZY1&R3D)[SM=?FHM&G2#L
/,.(fHZBU7a0f/3+1J+4RcaY088_@_<S13C6U0d:@ZW9Y6&X]bRM7[V]RUdZ&C<R
I34(,@-T)CM<>^[?)Ed-Y8;FQ2<:9->6)BFG;2/9N@e7NL(4?T7]VF_74EO_1A2&
aJPK3;K^M#&=Zc9EEA\:gL3R<??<F20U6:NN70=<M;:eYX>2N<\+XU&&?IET@0UU
5V[-9BRMd@e1D;^(_.F-_.82\dL2K&ReEbEPe385e9XVD&D[T/EdK9<[\I6E8;)T
3SK@.7=44P3F7.2/H9440^J<FP:)B,DKe=#\8?ZdX#P21K2NILa^7#CX-b8P/V5D
?:TCUa1AV424RKb:LAUN3Nad\Ug0G_V:cH&-9<aR-T1gI\AZ9]LKbC@5@HF(>9b:
Zb)PC8KB[^_LYB8fDU32S#L^_ETd?>)/8?fQe[<Q4Sd8FELEROI61XdSLS=:/G#_
5.G#:Ud0AB:(A+BTKJ0cdg7LI#W]Y=N)/ODURFGB=UWJ:.;CW\U_^?3d4/]&.5DL
2Oa&Y9Xc.a:[^H&IEP96_>(K,K^1,R_f_]BSK&B;&Q9H^RA?0A8BAK7P./3@?,GP
/c<Uf.PR8M32Hc)?Yc)(GB_Z=5Y)4d9FCUFU\0@fJ=HK-W(U18Q(1Q\+MKe0LBXU
GJgdDIf<Q.dg(A)M#LF6c?fKXE#11G5Z@Z-#O<->E4.H&^B=db[E5LYC(-ZO62CB
B0WJ&L=)6>WU15(L/VPA=DBK=2X[(MWR/d;?:]Q4-AA#[WD?MC1#7g?H#E;:QHJe
40Z(9Y\Ma(Lb=V(dZ)9WgH001RHMX>\d.4?F^4UUAbLMCWe+KE/S1<K6^8X3AU+f
c:XGPF^@=/<[I#/5-9>@/T:/=^3+&ObQTOPbWR70b0GQ3UGTKCdMY)N\RB-Z34d]
(:Pf2E;OF&&POPEVD?HF.JW_U(H@3X41D5fWU=\76@X]U&>RW@<IN68Xg&B)(5WF
.R\;KQQ(VUUZPA[&^L\X1VM\KcM,<d95.\N-748^@RX(fW6\SRG3J=3O]L(4VX2N
<EH2P.[+c4.VTT[&/P<4?QQ)K#T=aN]W4ZH3a/>_/b@b43T]daDK5[Cg]Za:29#V
G7aGGU&GJMF1<[KI9/>PZBF[&+8YBP1L&2CacO[\Oaf?R.[GSK?-K(,f9&Q2RVYb
,1W]]BN_/Z1B&(R8/d0>N:>EWX4+6@<1)DSQbPK5L2KH<G^K\^5.+(D[_)Ta2QI7
V9O+JT.T=#?g&ba062L]2COK_@3;Z,6SPW73[B?L9G1c6f\,J_;3[f1X\A<@((S7W$
`endprotected
  

endclass

`protected
+gM[A)9,d5036.NPFJ0cdJKV;C<08F?UeJ5f=ARUg14AJWL70N?^,)@EKOaMCJC1
<UgNg;]&7d>WAGNaP^c.4&MGcg/D&G0If.c;A)MPC895OLKNDQVYAATMcdQb,,68
+Eb19WK+YFP<KPA=^QbF_KaC2Mge=;36<7]OZX9K,f\eF4gSE[R6FgJJ/5cLS]?T
Q.f,7BefdVSc/Y62&9]_bS[eIN[=5TIX_Q^M\,-0&,B;gY/&24(KLPaRKb5IHCZb
e>9G_UBg[OU^ZBg_>E+]P;,B0BUEfZS(e>C4g8C+HWH+M/eV_@YNR-3bdP@&W7N1
Z52[I)gAJM(=M+c@bf(X,VGBc5+FFJ,_6c9fM/NB_Q(Gg9M<SaG:0]1Sd^N5HH,QV$
`endprotected


`endif // GUARD_SVT_APB_SLAVE_MONITOR_CALLBACK_SV
