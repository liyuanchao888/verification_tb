
`ifndef GUARD_SVT_AXI_PORT_MONITOR_DEF_COV_DATA_CALLBACK_SV
`define GUARD_SVT_AXI_PORT_MONITOR_DEF_COV_DATA_CALLBACK_SV

`include "svt_axi_defines.svi"
 
`define SVT_AXI_IS_XACT_COHERENT_READ(xact) \
(xact.xact_type == svt_axi_transaction::COHERENT) && \
( \
  (xact.coherent_xact_type == svt_axi_transaction::READNOSNOOP) || \
  (xact.coherent_xact_type == svt_axi_transaction::READONCE) || \
  (xact.coherent_xact_type == svt_axi_transaction::READSHARED) || \
  (xact.coherent_xact_type == svt_axi_transaction::READCLEAN) || \
  (xact.coherent_xact_type == svt_axi_transaction::READNOTSHAREDDIRTY) || \
  (xact.coherent_xact_type == svt_axi_transaction::READUNIQUE) || \
  (xact.coherent_xact_type == svt_axi_transaction::CLEANUNIQUE) || \
  (xact.coherent_xact_type == svt_axi_transaction::MAKEUNIQUE) || \
  (xact.coherent_xact_type == svt_axi_transaction::CLEANSHARED) || \
`ifdef SVT_ACE5_ENABLE \
  (xact.coherent_xact_type == svt_axi_transaction::CLEANSHAREDPERSIST) || \
`endif \
  (xact.coherent_xact_type == svt_axi_transaction::CLEANINVALID) || \
  (xact.coherent_xact_type == svt_axi_transaction::MAKEINVALID) || \
  (xact.coherent_xact_type == svt_axi_transaction::DVMCOMPLETE) || \
  (xact.coherent_xact_type == svt_axi_transaction::DVMMESSAGE) || \
  (xact.coherent_xact_type == svt_axi_transaction::READBARRIER) \
)

`define SVT_AXI_IS_XACT_COHERENT_WRITE(xact) \
(xact.xact_type == svt_axi_transaction::COHERENT) && \
( \
  (xact.coherent_xact_type == svt_axi_transaction::WRITENOSNOOP) || \
  (xact.coherent_xact_type == svt_axi_transaction::WRITELINEUNIQUE) || \
  (xact.coherent_xact_type == svt_axi_transaction::WRITEBARRIER) || \
  (xact.coherent_xact_type == svt_axi_transaction::WRITECLEAN) || \
  (xact.coherent_xact_type == svt_axi_transaction::WRITEBACK) || \
  (xact.coherent_xact_type == svt_axi_transaction::EVICT) || \
  (xact.coherent_xact_type == svt_axi_transaction::WRITEUNIQUE) || \
  (xact.coherent_xact_type == svt_axi_transaction::WRITEEVICT) \
)

typedef class svt_axi_port_monitor_callback;
typedef class svt_axi_cov;
`ifdef SVT_VMM_TECHNOLOGY
typedef class svt_axi_master_group;
`else
typedef class svt_axi_master_agent;
`endif
// =============================================================================
/**
 * The coverage data callback class defines default data and event information
 * that are used to implement the coverage groups. The coverage data callback
 * class is extended from callback class #svt_axi_port_monitor_callback. This
 * class itself does not contain any cover groups.  The constructor of this
 * class gets #svt_axi_port_configuration handle as an argument, which is used
 * for shaping the coverage.
 */
class svt_axi_port_monitor_def_cov_data_callback extends svt_axi_port_monitor_callback;

`ifndef SVT_AXI_EXCLUDE_AXI_PORT_COVERAGE
  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** Configuration object for shaping the coverage. */
  svt_axi_port_configuration cfg;

  /** Event used to trigger the read transaction covergroups for sampling. */
  event cov_read_sample_event;

  /** Event used to trigger the write/read transaction covergroups for sampling. */
  event cov_awakeup_sample_event;

  /** Event used to trigger the snoop transaction per burst covergroups for sampling. */
  event cov_snoop_sample_event;

  /** Event used to trigger the idle period of snoop channel toggles acwakeup signal for sampling. */
  event cov_snoop_sample_event_for_idle_snoop_chan;

  /** Event used to trigger the idle period of snoop channel toggles awakeup signal for sampling. */
  event cov_snoop_sample_event_for_awakeup_idle_snoop_chan;
 
  /** Event used to trigger the signal_master_valid_ready_dependency covergroup for sampling. */
  event cov_signal_dependency_event;

  /** Event used to trigger the signal_slave_valid_ready_dependency covergroup for sampling. */
  event cov_signal_slave_dependency_event;
  
  /** Event used to trigger the signal_master_slave_valid_ready_dependency covergroup for sampling. */
  event cov_signal_master_slave_dependency_event;

  /** Event used to trigger the signal_slave_master_valid_ready_dependency covergroup for sampling. */
  event cov_signal_slave_master_dependency_event;

  /** Event used to trigger the snoop transaction per beat within a burst covergroups for sampling. */
  event cov_snoop_per_beat_sample_event;

  /** Event used to trigger the write transaction covergroups for sampling. */
  event cov_write_sample_event;

  /** Event used to trigger the read and write outstanding transaction covergroups for sampling. */
  event cov_outstanding_event;
  /** Event used to trigger the read and write interleaving transaction covergroups for sampling. */
  event cov_interleave_depth_event;  
  
  /** Event used to trigger stream data interleaving transaction covergroups for sampling. */
  event cov_stream_interleave_depth_event;  

  /** Event used to trigger the write out-of-order response covergroups for sampling. */
  event cov_out_of_order_write_response_depth_event;

  /** Event used to trigger the read out-of-order response covergroups for sampling. */
  event cov_out_of_order_read_response_depth_event;

  /** Event used to trigger the stream covergroups for sampling. */
  event cov_stream_sample_event;
  /** Event used to trigger write completed out of order covergroups */
  event cover_arid_awid_diff_out_of_order_event;
  /** Event used to trigger read completed out of order covergroups */
  event cover_arid_awid_equal_out_of_order_event;
  /** Event used to trigger READs completed back to back */
   event back_to_back_read_burst_event;
 /** Event used to trigger WRITEs completed back to back */
  event back_to_back_write_burst_event;
 /** Event used to trigger Four WRITEs/READs address handshake completed */
  event four_state_rd_wr_event;
 /** Event used to trigger sequence of four Exclusive/Normal transactions */
  event four_excl_normal_seq_event; 
 /** Event used to trigger wstrb signalling unaligned start address */
  event wstrb_to_signal_unaligned_start_address_event;

  /** Event used to trigger the read and write barrier transaction covergroups for sampling. */
  event cov_barrier_outstanding_event;
  /** Event used to trigger the read and write barrier transaction covergroups for sampling. */
  event cov_barrier_outstanding_event_ace;
  /** Event used to trigger the read and write barrier transaction covergroups for sampling. */
  event cov_barrier_outstanding_event_acelite;

  /** Event used to trigger xacts followed the lanuch of 256 outstanding barrier covergroup for sampling. */
  event cov_non_barrier_after_256_outstanding_barrier_sample_event;

  /**  Event used to trigger trans_master_snoop_to_same_address_as_read_xact */
  event cov_snoop_to_same_addr_as_read_xact_event;

  /** Event used to trigger trans_master_snoop_to_same_addr_as_memory_update_exclude_writeevict */
  event cov_snoop_to_same_addr_as_memory_update_event;

  /** Event used to trigger trans_master_snoop_to_same_addr_as_writeevict */
  event cov_snoop_to_same_addr_as_writeevict_event;

  /** Event used to trigger trans_master_snoop_resp_during_wu_wlu_to_same_addr */
  event cov_snoop_to_same_addr_as_wu_wlu_event;

  /** Event used to trigger trans_master_snoop_data_transfer_during_wu_wlu_to_same_addr */
  event cov_snoop_with_datatransfer_to_same_addr_as_wu_wlu_event;

  /** Event used to trigger trans_master_readunique_snoop_resp_datatransfer_with_clean_cacheline */
  event cov_readunique_snoop_resp_datatransfer_with_clean_cacheline_event;

  /** Event used to trigger trans_cross_master_to_slave_path_access */ 
  event cov_master_to_slave_access_event;
 
 /** Events to trigger DVM overlap case related covergroup*/
  event dvm_overlap_scenarios_snoop_addr_event;
  event dvm_overlap_scenarios_snoop_resp_event;

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Coverpoint variable used to hold the received transaction through pre_output_port_put callback method. */
  protected svt_axi_transaction cov_item;
  
  /** Snoop transaction Coverpoint variable used to hold the received transaction through pre_snoop_output_port_put callback method. */
  protected svt_axi_snoop_transaction cov_snoop_item;

  /** Snoop transaction handle when sampled at the point that snoop transaction just started */
  protected svt_axi_snoop_transaction cov_snoop_addr_item;

  /** Coverpoint variable use to hold the value of coherent_xact_type for covergroup trans_ace_concurrent_overlapping_arsnoop_acsnoop */
  protected svt_axi_transaction::coherent_xact_type_enum master_coherent_xact_type ;
  
  /** Coverpoint variable use to hold the value of snoop_xact_type for covergroup trans_ace_concurrent_overlapping_arsnoop_acsnoop */
  protected svt_axi_snoop_transaction::snoop_xact_type_enum master_snoop_xact_type;

 /** Coverpoint variable use to hold the value of coherent_write_xact_type for trans_ace_concurrent_overlapping_awsnoop_acsnoop covergroup  */
  protected svt_axi_transaction::coherent_xact_type_enum coherent_write_xact_type_generate_snoop;  

  /** Coverpoint variable used to hold the ACVALID to ACREADY delay. */
  protected int cov_ACVALID_to_ACREADY_Delay;
  
  /** Coverpoint variable used to hold the ACVALID to ACWAKEUP delay. */
  protected int cov_ACWAKEUP_before_ACVALID_Delay;

  /** Coverpoint variable used to hold the ACWAKEUP to ACVALID delay. */
  protected int cov_ACWAKEUP_after_ACVALID_Delay;
 
  /** Coverpoint variable used to hold the ACWAKEUP and ACVALID same time assertion delay. */
  protected int cov_ACWAKEUP_ACVALID_same_time;
  
  /** Coverpoint variable used to hold the ACWAKEUP toggle delay during idle period of snoop channel delay. */
  protected int cov_ACWAKEUP_toggle_Delay_idle_snoop_chan;

 /** Coverpoint variable used to hold the ACWAKEUP toggle assertion delay during idle period of snoop channel. */
  protected int idle_snoop_chan_wakeup_toggle_assertion_cycle;

  /** Coverpoint variable used to hold the ACWAKEUP to previous ACWAKEUP dealy. */
  protected int cov_ACWAKEUP_to_prev_ACWAKEUP_Delay;
///////////
    /** Coverpoint variable used to hold the ARVALID to AWAKEUP delay. */
  protected int cov_AWAKEUP_before_ARVALID_Delay;

  /** Coverpoint variable used to hold the AWAKEUP to ARVALID delay. */
  protected int cov_AWAKEUP_after_ARVALID_Delay;
 
  /** Coverpoint variable used to hold the AWAKEUP and ARVALID same time assertion delay. */
  protected int cov_AWAKEUP_ARVALID_same_time;
  
  /** Coverpoint variable used to hold the AWAKEUP toggle delay during idle period of snoop channel delay. */
  protected int cov_AWAKEUP_toggle_Delay_idle_chan;

 /** Coverpoint variable used to hold the AWAKEUP toggle assertion delay during idle period of snoop channel. */
  protected int idle_chan_wakeup_toggle_assertion_cycle;

  /** Coverpoint variable used to hold the AWAKEUP to previous AWAKEUP dealy. */
  protected int cov_AWAKEUP_to_prev_AWAKEUP_Delay;

  /** Coverpoint variable used to hold the AWAKEUP toggle delay during idle period of snoop channel delay. */
  protected int cov_AWAKEUP_toggle_Delay_idle_snoop_chan;

  /** Coverpoint variable used to hold the AWAKEUP toggle assertion delay during idle period of snoop channel. */
  protected int idle_snoop_chan_awakeup_toggle_assertion_cycle;

  /** Coverpoint variable used to hold the ACVALID to CRVALID delay. */
  protected int cov_ACVALID_to_CRVALID_Delay;

  /** Coverpoint variable used to hold the CRVALID to last_RVALID_RREADY_handshake_to_next_RVALID_DelayRREADY delay. */
  protected int cov_CRVALID_to_CRREADY_Delay;

  /** Coverpoint variable used to hold the WVALID to WREADY delay. */
  protected int cov_CDVALID_to_CDREADY_Delay;

  /** Coverpoint variable used to hold the AWVALID to AWREADY delay. */
  protected int cov_AWVALID_to_AWREADY_Delay;

  /** Coverpoint variable used to hold the ARVALID to ARREADY delay. */
  protected int cov_ARVALID_to_ARREADY_Delay;

  /** Coverpoint variable used to hold the WVALID to WREADY delay. */
  protected int cov_WVALID_to_WREADY_Delay;

  /** Coverpoint variable used to hold the TVALID to TREADY delay. */
  protected int cov_TVALID_to_TREADY_Delay;

  /** Coverpoint variable used to hold the TVALID delay. */
  protected int cov_TVALID_Delay;

  /** Coverpoint variable used to hold the TREADY delay. */
  protected int cov_TREADY_Delay;

  /** Coverpoint variable used to hold the RVALID to RREADY delay. */
  protected int cov_RVALID_to_RREADY_Delay;

  /** Coverpoint variable used to hold the BVALID to next BVALID delay. */
  protected int cov_BVALID_to_next_BVALID_Delay;

  /** Coverpoint variable used to hold the BVALID to BREADY delay. */
  protected int cov_BVALID_to_BREADY_Delay;

  /** Coverpoint variable used to hold the AWVALID to previous AWVALID dealy. */
  protected int cov_AWVALID_to_prev_AWVALID_Delay;

  /** Coverpoint variable used to hold the AWVALID to previous handshake dealy. */
  protected int cov_prev_handshake_AWVALID_Delay;

  /** Coverpoint variable used to hold the previous handshake to AWREADY dealy. */
  protected int cov_prev_handshake_AWREADY_Delay;

  /** Coverpoint variable used to hold the write address handshake to previous AWREADY dealy. */
  protected int cov_prev_AWREADY_to_handshake_Delay;

  /** Coverpoint variable used to hold the WVALID to previous WVALID dealy. */
  protected int cov_WVALID_to_prev_WVALID_Delay;

  /** Coverpoint variable used to hold the TVALID to previous TVALID dealy. */
  protected int cov_TVALID_to_prev_TVALID_Delay;

  /** Coverpoint variable used to hold the AWVALID to first WVALID dealy. */
  protected int cov_AWVALID_to_first_WVALID_Delay;

  /** Coverpoint variable used to hold the last write data handshake to BVALID dealy. */
  protected int cov_last_wdata_handshake_to_BVALID_Delay;

  /** Coverpoint variable used to hold the ARVALID to previous ARVALID dealy. */
  protected int cov_ARVALID_to_prev_ARVALID_Delay;

  /** Coverpoint variable used to hold the RVALID to previous RVALID dealy. */
  protected int cov_RVALID_to_prev_RVALID_Delay;

  /** Coverpoint variable used to hold the ARVALID to first RVALID dealy. */
  protected int cov_ARVALID_to_first_RVALID_Delay;
  
  /** Coverpoint variable used to hold the last AWVALID_AWREADY handshake to next AWVALID AWREADY handshake delay. */
  protected int cov_last_AWVALID_AWREADY_handshake_to_next_AWVALID_AWREADY_handshake_Delay;
  /** Coverpoint variable used to hold the last AWVALID_AWREADY handshake to next AWVALID delay. */
  protected int cov_last_AWVALID_AWREADY_handshake_to_next_AWVALID_Delay;
  /** Coverpoint variable used to hold the last AWVALID_AWREADY handshake to next AWREADY delay. */
  protected int cov_last_AWVALID_AWREADY_handshake_to_next_AWREADY_Delay;

  /** Coverpoint variable used to hold the last WVALID_WREADY handshake to next WVALID_WREADY handshake delay. */
  protected int cov_last_WVALID_WREADY_handshake_to_next_WVALID_WREADY_handshake_Delay;
  /** Coverpoint variable used to hold the last WVALID_WREADY handshake to next WVALID_WREADY handshake delay. */
  protected int cov_last_WVALID_WREADY_data_beat_handshake_to_next_WVALID_WREADY_first_data_beat_handshake_Delay;
  /** Coverpoint variable used to hold the last WVALID_WREADY handshake to next WVALID delay. */
  protected int cov_last_WVALID_WREADY_handshake_to_next_WVALID_Delay;
  /** Coverpoint variable used to hold the last WVALID_WREADY handshake to next WREADY delay. */
  protected int cov_last_WVALID_WREADY_handshake_to_next_WREADY_Delay;
  /** Coverpoint variable used to hold the last WREADY to next WVALID_WREADY handshake delay. */
  protected int cov_last_WREADY_to_next_WVALID_WREADY_handshake_Delay;

  /** Coverpoint variable used to hold the last BVALID_BREADY handshake to next BVALID_BREADY handshake delay. */
  protected int cov_last_BVALID_BREADY_handshake_to_next_BVALID_BREADY_handshake_Delay;
  /** Coverpoint variable used to hold the last BVALID_BREADY handshake to next BVALID delay. */
  protected int cov_last_BVALID_BREADY_handshake_to_next_BVALID_Delay;
  /** Coverpoint variable used to hold the last BVALID_BREADY handshake to next BREADY delay. */
  protected int cov_last_BVALID_BREADY_handshake_to_next_BREADY_Delay;

  /** Coverpoint variable used to hold the last ARVALID_ARREADY handshake to next ARVALID ARREADY handshake delay. */
  protected int cov_last_ARVALID_ARREADY_handshake_to_next_ARVALID_ARREADY_handshake_Delay;
  /** Coverpoint variable used to hold the previous handshake to ARREADY dealy. */
  protected int cov_prev_handshake_ARREADY_Delay;
  /** Coverpoint variable used to hold the last ARVALID_ARREADY handshake to next ARVALID delay. */
  protected int cov_prev_handshake_ARVALID_Delay;
  /** Coverpoint variable used to hold the last ARVALID_ARREADY handshake to next ARREADY delay. */
  protected int cov_last_ARVALID_ARREADY_handshake_to_next_ARREADY_Delay;

  /** Coverpoint variable used to hold the last RVALID_RREADY handshake to next RVALID RREADY handshake delay. */
  protected int cov_last_RVALID_RREADY_handshake_to_next_RVALID_RREADY_handshake_Delay;
  /** Coverpoint variable used to hold the last RVALID_RREADY handshake to next RVALID delay. */
  protected int cov_last_RVALID_RREADY_handshake_to_next_RVALID_Delay ;
  /** Coverpoint variable used to hold the last RVALID_RREADY handshake to next RREADY delay. */
  protected int cov_last_RVALID_RREADY_handshake_to_next_RREADY_Delay;

  /** Coverpoint variable used to hold the last RVALID_RREADY handshake to next RVALID_RREADY handshake delay. */
  protected int cov_last_RVALID_RREADY_data_beat_handshake_to_next_RVALID_RREADY_first_data_beat_handshake_Delay;
  /** Coverpoint variable used to hold the last RREADY to next RVALID_RREADY handshake delay. */
  protected int cov_last_RREADY_to_next_RVALID_RREADY_handshake_Delay;
  /** Coverpoint variable used to hold the arite address handshake to previous ARREADY dealy. */
  protected int cov_prev_ARREADY_to_handshake_Delay;
  /** Coverpoint variable used to hold the last BREADY to next BREADY delay. */
  protected int cov_last_BREADY_to_next_BREADY_Delay;
  /** Coverpoint variable used to hold the last BREADY to next BVALID_BREADY handshake delay. */
  protected int cov_last_BREADY_to_next_BVALID_BREADY_handshake_Delay;

  /** Coverpoint variable used to hold the WSTRB. */
  protected reg [256:0] cov_wstrb;

  /** Coverpoint variable used to hold the RCHUNKSTRB. */
  protected reg [7:0] cov_rchunkstrb;

  /** Coverpoint variable used to hold the RCHUNKNUM. */
  protected reg [7:0] cov_rchunknum;

  /** Coverpoint variable used to hold the RRESP. */
  protected svt_axi_transaction::resp_type_enum cov_rresp;

  /** Coverpoint variable used to hold the response type */
  protected svt_axi_transaction::resp_type_enum m_response_type;

  /** Coverpoint variable used to hold the aligned address */
  protected bit [5:0]   m_address_aligned;  

/** Coverpoint variable used to hold OOO write transactions. */
  protected int write_completed_out_of_order = -1;
  protected int write_completed_out_of_order_same_id_as_read = -1;
/** Coverpoint variable used to hold OOO write transactions. */
  protected int read_completed_out_of_order = -1;
  protected int read_completed_out_of_order_same_id_as_write = -1;
  protected int num_read_outstanding_xact_arid = -1;
/** Coverpoint variable used to hold Back To Back READ/WRITE transactions. */
  protected int back_to_back_read_burst_sequence = -1;
  protected int back_to_back_write_burst_sequence = -1;
/** Coverpoint variable used to hold Four State Write/Read xacts. */
  protected int four_state_rd_wr_burst_sequence=-1;
/** Coverpoint variable used to hold four Exclusive/Normal xacts. */
  protected int four_excl_normal_sequence = -1;
/** Coverpoint variable used to hold wstrb signalling unaligned transfer xacts. */
  protected int wstrb_to_signal_unaligned_start_address=-1;
  /**AXI COV DATA */
  protected svt_axi_cov cov_data;
  
  /** Coverpoint variable used to hold the CRRESP[4:0]. */
  protected reg [4:0] cov_crresp;
 
  /** Coverpoint variable used to hold the number of slaves in the system. */
  protected int num_slaves;
  
  /** Coverpoint variable used to hold the slave id in transaction. */
  protected int slave_id;

  /** Coverpoint variable used to hold the coherent_xact_type initiated by 
   * ACE-Lite Master.Used in trans_master_ace_lite_coherent_and_ace_snoop_response_association
   * covergroup 
   */  
  protected svt_axi_transaction::coherent_xact_type_enum ace_lite_coh_xact_type = svt_axi_transaction::READNOSNOOP;

 /** Coverpoint variable used to hold the coherent_xact_type initiated by 
   * ACE Master.Used in trans_master_ace_coherent_and_ace_snoop_response_association
   * covergroup 
   */  
  protected svt_axi_transaction::coherent_xact_type_enum ace_coh_xact_type;

 /** Coverpoint variable used to hold the snoop_xact_type on ACE Master
   * Used in trans_master_ace_lite_coherent_and_ace_snoop_response_association
   * covergroup 
   */  
  protected svt_axi_snoop_transaction::snoop_xact_type_enum ace_lite_master_snoop_xact_type ;

 /** Coverpoint variable used to hold the snoop_xact_type on ACE Master
   * Used in trans_master_ace_coherent_and_ace_snoop_response_association
   * covergroup 
   */  
  protected svt_axi_snoop_transaction::snoop_xact_type_enum ace_master_snoop_xact_type ;

  /** Coverpoint variables used to hold the back to back coherent_xact_type initiated by 
   * ACE-Lite Master.Used in trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id
   * covergroup 
   */
  protected svt_axi_transaction::coherent_xact_type_enum ace_lite_coh_xact_t1_type = svt_axi_transaction::READNOSNOOP;
  protected svt_axi_transaction::coherent_xact_type_enum ace_lite_coh_xact_t2_type = svt_axi_transaction::READNOSNOOP;
  
  /** Coverpoint variable used to hold the CRRESP[4:0]. Used in
   * trans_master_ace_lite_coherent_and_ace_snoop_response_association
   * covergroup 
   */
  protected reg [4:0] snoop_resp_from_ace_master;

  /** Coverpoint variables used to hold the CRRESP[4:0]. Used in
   * trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id
   * covergroup.
   */
  protected reg [4:0] snoop_resp_t1_from_ace_master;
  protected reg [4:0] snoop_resp_t2_from_ace_master;
 
  /** Coverpoint variable used to hold the specific id. Used in
   * trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id
   * covergroup.
   */
  protected int ace_lite_coh_xact_id;

  /** Coverpoint variable used to hold the CRRESP[4:0]. Used in
   * trans_ace_concurrent_overlapping_awsnoop_acsnoop
   * covergroup 
   */
  protected reg [4:0] snoop_resp_ace_master;

  /** Coverpoint variable used to hold the initial cache state of Snooped 
   * ACE-master corresponding to a coherent transaction initiated from ACE
   * Master. Used in trans_master_ace_lite_coherent_and_ace_snoop_response_association
   * covergroup. The possible states correspond to the 5 states of a cache line, namely, 
   * INVALID, UNIQUECLEAN, SHAREDCLEAN, UNIQUEDIRTY and SHAREDDIRTY. 
   */  
  protected svt_axi_snoop_transaction::cache_line_state_enum ace_master_init_cache_state = svt_axi_snoop_transaction::INVALID;

  /** Coverpoint variable used to hold the final cache state of Snooped 
   * ACE-master corresponding to a coherent transaction initiated from ACE
   * Master. Used in trans_master_ace_lite_coherent_and_ace_snoop_response_association
   * covergroup. The possible states correspond to the 5 states of a cache line, namely, 
   * INVALID, UNIQUECLEAN, SHAREDCLEAN, UNIQUEDIRTY and SHAREDDIRTY. 
   */  
  protected svt_axi_snoop_transaction::cache_line_state_enum ace_master_final_cache_state = svt_axi_snoop_transaction::INVALID;  

  /** Coverpoint variable used to hold the total number of outstanding transactions. */ 
  protected int num_outstanding_xact = 0;
 
  /** Coverpoint variable used to hold the number of read outstanding transactions. */
  protected int num_read_outstanding_xact = 0;
  
  /** Coverpoint variable used to hold the number of outstanding snoop transactions. */
  protected int num_outstanding_snoop_xacts = 0;
  
  /** Coverpoint variable used to hold the number of write outstanding transactions. */
  protected int num_write_outstanding_xact = 0;
  /** Coverpoint variable used to hold the number of barrier outstanding transactions. */
  protected int num_barrier_outstanding_xact = 0;
  /** Coverpoint variable used to hold the number of write outstanding transactions. */
  protected int read_outstanding_xact_same_arid_cache_modifiable_bit = -1;
  /** Coverpoint variable used to hold the number of write outstanding transactions. */
  protected int read_outstanding_xact_diff_arid_cache_modifiable_bit = -1;
  /** Coverpoint variable used to hold the memory type of read outstanding transactions. */
  protected int read_outstanding_xact_diff_arid_device_cacheable_bit = -1;
  /** Coverpoint variable used to hold the number of write outstanding transactions. */
  protected int write_outstanding_xact_same_awid_cache_modifiable_bit = -1;
  /** Coverpoint variable used to hold the number of write outstanding transactions. */
  protected int write_outstanding_xact_diff_awid_cache_modifiable_bit = -1;
  /** Coverpoint variable used to hold the memory type of write outstanding transactions. */
  protected int write_outstanding_xact_diff_awid_device_cacheable_bit = -1;
  /** Coverpoint variable used to hold the number of read outstanding transactions with an ARID
   * value matching to the ID value which is configured in 
   * svt_axi_port_configuration::cov_same_id_in_outstanding_xacts. 
   **/
  protected int read_outstanding_xacts_with_same_arid = 0;
  /** Coverpoint variable used to hold the number of read outstanding transactions with an ARID
   * value matching to the ID value which is configured in 
   * svt_axi_port_configuration::cov_multi_same_ids. 
   **/
  protected int cov_num_read_outstanding_same_arid = 0;
  /** Coverpoint variable used to hold an ARID
   * value matching to the ID value which is configured in 
   * svt_axi_port_configuration::cov_multi_same_ids. 
   **/
  protected int cov_read_same_id = 0;
  /** Coverpoint variable used to hold the number of write outstanding transactions with an AWID
   * value matching to the ID value which is configured in 
   * svt_axi_port_configuration::cov_multi_same_ids. 
   **/
  protected int cov_num_write_outstanding_same_awid = 0;
  /** Coverpoint variable used to hold an AWID
   * value matching to the ID value which is configured in 
   * svt_axi_port_configuration::cov_multi_same_ids. 
   **/
  protected int cov_write_same_id = 0;
  /** Coverpoint variable used to hold the number of outstanding transactions with DVM TLBI requests with same ARID */ 
  protected int num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid = 0;
  /** Coverpoint variable used to hold the number of outstanding transactions with DVM TLBI requests with different ARID */ 
  protected int num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid = 0;
  /** Internal Queue to hold the IDs of outstanding DVM TLBI transactions.This queue is used to find the number of outstanding DVM TLBI transactions with uunique IDs */ 
  protected int dvm_tlbi_outstanding_xacts_arid[$];
  /** Coverpoint variable used to hold the number of read outstanding transactions with diff ARID. */
  protected int read_outstanding_xacts_with_diff_arid = 0;
  /** Coverpoint variable used to hold the number of write outstanding transactions with an AWID
   * value matching to the ID value which is configured in 
   * svt_axi_port_configuration::cov_same_id_in_outstanding_xacts. 
   **/
  protected int write_outstanding_xacts_with_same_awid = 0;  
  /** Coverpoint variable used to hold the number of write outstanding transactions with diff AWID. */
  protected int write_outstanding_xacts_with_diff_awid = 0;
  /** Coverpoint variable used to hold the depth of out-of-order write response. */
  protected int out_of_order_write_response_depth = 0;

  /** Coverpoint variable used to hold number of out-of-order write response count. */ 
  protected bit axi_write_resp_OOO_count = 0;
  /** Coverpoint variable used to hold the depth of out-of-order write response. */
  protected int out_of_order_read_response_depth = 0;

 /** Coverpoint variable used to hold number of out-of-order read_response count. */ 
  protected bit axi_read_resp_OOO_count = 0;

  /* variable used to hold the outstanding write transaction. */
  protected svt_axi_transaction write_outstanding_xact_queue[$];

  /* variable used to hold the outstanding read transaction. */
  protected svt_axi_transaction read_outstanding_xact_queue[$];
  
  /* variable used to hold the outstanding snoop transaction. */
  protected svt_axi_snoop_transaction snoop_outstanding_xact_queue[$];
  
  /* variable used to hold the completed read transaction. */
  protected svt_axi_transaction read_xactQ[$];

  /* variable used to hold the arready of the previous xact */
  protected int prev_addr_arready_assertion_cycle = 0;

  /** Coverpoint variable to store the previous AWVALID assertion cycle. */
  protected int prev_addr_awvalid_assertion_cycle = 0;

  /* variable used to hold the awready of the previous xact */
  protected int prev_addr_awready_assertion_cycle = 0;
  /* variable used to hold the completed write transaction. */
  protected svt_axi_transaction write_xactQ[$];
  /* variable used to hold the address phase completed RD/WR xacts. */
  protected bit four_state_rd_wr_queue[$];
  /* variable used to hold completed Excl/Normal xacts. */
  protected bit four_excl_normal_seq_queue[$];
  
  /* variable used to hold the slave indexes */
  protected	int slv_num [];

  /* variable used to hold the slave indexes from configuration */
  protected	int slv_num_cfg []; 

  /* variable used to hold the ignored slaves from the slaves list*/
  svt_amba_addr_mapper::path_cov_dest_names_enum ignore_slaves_list[];

  /* variable used to hold the ignored slaves in the queue */
  svt_amba_addr_mapper::path_cov_dest_names_enum ignore_slaves_list_q[$];

  /* variable used to hold the ignored slaves from the slaves list by configuration */
  svt_amba_addr_mapper::path_cov_dest_names_enum ignore_cfg_slaves_list[];

  /* variable used to hold the ignored slaves in the queue by configuration */
  svt_amba_addr_mapper::path_cov_dest_names_enum ignore_cfg_slaves_list_q[$];

  /* variable used to hold the slave names */
  svt_amba_addr_mapper::path_cov_dest_names_enum path_cov_dest_names,slv_m,slv_t,slv_hit, t_slave;

  /* variable used to hold the number of slave configuration */
  int num_of_slave_configs;
  
  /** Coverpoint variable used to hold the number of read transactions that were interleaved. */
  protected int read_data_interleaving_depth = 1;
  
  /** Coverpoint variable used to hold the number of write transactions that were interleaved.. */
  protected int write_data_interleaving_depth = 1; 
  
  /** Coverpoint variable used to hold the number of stream transactions that were interleaved. */
  protected int axi4_stream_data_interleaving_depth = 1;

  /** Variable used to count the number of read transactions. */
  protected int count_read = 0;
 
  /** Variable used to count the number of stream transactions. */
  protected int count_stream = 0;

 /** Variable used to count the number of ACE_LITE masters present in the system */
  protected int count_ace_lite = 0;

 /** Variable used to count the number of ACE masters present in the system */
  protected int count_ace = 0;
 
 /** Variable used to hold outstanding transactions. */
  protected int out_standing_xacts = 0;

  /** Variable used to count the number of write transactions. */
  protected int count_write = 0;    
  
  /** Coverpoint variable used to hold the previous rid value. */
  protected int previous_rid = 0;
  
  /** Coverpoint variable used to hold the previous wid value. */
  protected int previous_wid = 0;

  /** Coverpoint variable used to hold the previous tid value. */
  protected int previous_tid = 0;
  protected int previous_burst_length = 0;

  /** Coverpoint variable used to hold the RRESP[3:0] for DVM messages. */
  protected reg [3:0] cov_dvm_rresp;
  
  /** Coverpoint variable used to hold the COH_RRESP. */
  protected svt_axi_transaction::coherent_resp_type_enum cov_coherent_rresp;

  /** 
   * Coverpoint variable used to hold the Read or Write transaction type.  If
   * #svt_axi_port_configuration::axi_interface_type is AXI_ACE then
   * #svt_axi_transaction::coherent_xact_type READNOSNOOP is considered as READ
   * transactions and #svt_axi_transaction::coherent_xact_type WRITENOSNOOP is
   * considered as WRITE transactions for AXI3/AXI4/AXI4_LITE related covergroups.
   */
  protected svt_axi_transaction::xact_type_enum cov_xact_rd_wr_type;
  
  /** Coverpoint variable to store last AWVALID_AWREADY handshaking assertion cycle. */
  protected int  last_write_addr_ready_assertion_cycle;

  /** Coverpoint variable to store last WVALID_WREADY handshaking assertion cycle. */
  protected int  last_write_data_ready_assertion_cycle;

  /** Coverpoint variable to store last BVALID_BREADY handshaking assertion cycle. */
  protected int last_write_resp_ready_assertion_cycle;

  /** Coverpoint variable to store last ARVALID_ARREADY handshaking assertion cycle. */
  protected int last_read_addr_ready_assertion_cycle;

  /** Coverpoint variable to store last RVALID_RREADY handshaking assertion cycle. */
  protected int last_read_data_ready_assertion_cycle;

  /** Coverpoint variable to store the previous WVALID assertion cycle. */
  protected int prev_write_data_valid_assertion_cycle;

  /** Coverpoint variable to store the previous BVALID assertion cycle. */
  protected int prev_write_resp_valid_assertion_cycle;

  /** Coverpoint variable to store the previous ARVALID assertion cycle. */
  protected int prev_read_arvalid_assertion_cycle;

  /** Coverpoint variable to store the previous RVALID assertion cycle. */
  protected int prev_read_data_valid_assertion_cycle;

  /** Coverpoint variable used to hold the ACVALID to previous ACVALID dealy. */
  protected int cov_ACVALID_to_prev_ACVALID_Delay;
  
  /** Coverpoint variable used to hold the CRVALID to previous CRVALID dealy. */
  //protected int cov_CRVALID_to_prev_CRVALID_Delay;
  
  /** Coverpoint variable used to hold the CDVALID to previous CDVALID dealy. */
  protected int cov_CDVALID_to_prev_CDVALID_Delay;
  
  /** Coverpoint variable to store the previous ACVALID assertion cycle. */
  protected int prev_snoop_addr_valid_assertion_cycle;

  /** Coverpoint variable to store the previous ACVALID assertion cycle. */
  protected int prev_snoop_addr_acwakeup_assertion_cycle;

  /** Coverpoint variable to store the previous ARVALID assertion cycle. */
  protected int prev_addr_acwakeup_assertion_cycle;

  /** Coverpoint variable to store the previous CRVALID assertion cycle. */
  protected int prev_snoop_resp_valid_assertion_cycle;

  /** Coverpoint variable to store the previous CDVALID assertion cycle. */
  protected int prev_snoop_data_valid_assertion_cycle;
   
  /** Coverpoint variable to store the kind of STREAM */
  protected svt_axi_transaction::stream_xact_type_enum cov_stream_xact_type;

  /** Coverpoint variable to store the status if acvalid is asserted before acready. */
  bit cov_ACVALID_before_ACREADY;
  /** Coverpoint variable to store the status if acready is asserted before acvalid. */
  bit cov_ACREADY_before_ACVALID;
  /** Coverpoint variable to store the status if crvalid is asserted before crready. */
  bit cov_CRVALID_before_CRREADY;
  /** Coverpoint variable to store the status if crready is asserted before crvalid. */
  bit cov_CRREADY_before_CRVALID;
  /** Coverpoint variable to store the status if cdvalid is asserted before cdready. */
  bit cov_CDVALID_before_CDREADY;
  /** Coverpoint variable to store the status if cdready is asserted before cdvalid. */
  bit cov_CDREADY_before_CDVALID;

  /** Coverpoint variable to store the status if arvalid is asserted before arready. */
  bit cov_ARVALID_before_ARREADY;
  /** Coverpoint variable to store the status if arready is asserted before arvalid. */
  bit cov_ARREADY_before_ARVALID;
  /** Coverpoint variable to store the status if rvalid is asserted before rready. */
  bit cov_RVALID_before_RREADY;
  /** Coverpoint variable to store the status if rready is asserted before rvalid. */
  bit cov_RREADY_before_RVALID;
  
  /** Coverpoint variable to store the status if awvalid is asserted before awready. */
  bit cov_AWVALID_before_AWREADY;
  /** Coverpoint variable to store the status if awready is asserted before awvalid. */
  bit cov_AWREADY_before_AWVALID;
  /** Coverpoint variable to store the status if awvalid is asserted before wready. */
  bit cov_AWVALID_before_WREADY;
  /** Coverpoint variable to store the status if wready is asserted before awvalid. */
  bit cov_WREADY_before_AWVALID; 
  /** Coverpoint variable to store the status if wvalid is asserted before awready. */
  bit cov_WVALID_before_AWREADY;
  /** Coverpoint variable to store the status if awready is asserted before wvalid. */
  bit cov_AWREADY_before_WVALID;
  /** Coverpoint variable to store the status if wvalid is asserted before wready. */
  bit cov_WVALID_before_WREADY;
  /** Coverpoint variable to store the status if tvalid is asserted before tready. */
  bit cov_TVALID_before_TREADY;
  /** Coverpoint variable to store the status if wready is asserted before wvalid. */
  bit cov_WREADY_before_WVALID;
    /** Coverpoint variable to store the status if tready is asserted before tvalid. */
  bit cov_TREADY_before_TVALID;
  /** Coverpoint variable to store the status if awvalid is asserted before wvalid. */
  bit cov_AWVALID_before_WVALID;
  /** Coverpoint variable to store the status if wvalid is asserted before awvalid. */
  bit cov_WVALID_before_AWVALID;
  /** Coverpoint variable to store the status if bvalid is asserted before bready. */
  bit cov_BVALID_before_BREADY;
  /** Coverpoint variable to store the status if bready is asserted before bvalid. */
  bit cov_BREADY_before_BVALID; 
  /** Coverpoint variable to store the status if awvalid is deasserted after wvalid. */
  bit cov_awvalid_wvalid = 0; 
  /** Coverpoint variable to store the status if awvalid is deasserted after rready. */
  bit cov_awvalid_rready = 0;
  /** Coverpoint variable to store the status if awvalid is deasserted after bready. */
  bit cov_awvalid_bready = 0;
  /** Coverpoint variable to store the status if wvalid is deasserted after awvalid. */
  bit cov_wvalid_awvalid = 0;
  /** Coverpoint variable to store the status if wvalid is deasserted after rready. */
  bit cov_wvalid_rready = 0;
  /** Coverpoint variable to store the status if wvalid is deasserted after bready. */
  bit cov_wvalid_bready = 0;
  /** Coverpoint variable to store the status if rready is deasserted after wvalid. */
  bit cov_rready_awvalid = 0;
  /** Coverpoint variable to store the status if rready is deasserted after wvalid. */
  bit cov_rready_wvalid = 0;
  /** Coverpoint variable to store the status if rready is deasserted after bready. */
  bit cov_rready_bready = 0;
  /** Coverpoint variable to store the status if bready is deasserted after awvalid. */
  bit cov_bready_awvalid = 0;
  /** Coverpoint variable to store the status if bready is deasserted after wvalid. */
  bit cov_bready_wvalid = 0;
  /** Coverpoint variable to store the status if bready is deasserted after rready. */
  bit cov_bready_rready = 0;
  
  /** Coverpoint variable to store the status if wready is deasserted after arready. */
  bit cov_wready_arready = 0;
  /** Coverpoint variable to store the status if wready is deasserted after rvalid. */
  bit cov_wready_rvalid = 0;
  /** Coverpoint variable to store the status if wready is deasserted after bvalid. */
  bit cov_wready_bvalid = 0;
  /** Coverpoint variable to store the status if arready is deasserted after wready. */
  bit cov_arready_wready = 0;
  /** Coverpoint variable to store the status if arready is deasserted after rvalid. */
  bit cov_arready_rvalid = 0;
  /** Coverpoint variable to store the status if arready is deasserted after bvalid. */
  bit cov_arready_bvalid = 0;  
  /** Coverpoint variable to store the status if rvalid is deasserted after arready. */
  bit cov_rvalid_arready = 0;
  /** Coverpoint variable to store the status if rvalid is deasserted after wready. */
  bit cov_rvalid_wready = 0;
  /** Coverpoint variable to store the status if rvalid is deasserted after bvalid. */
  bit cov_rvalid_bvalid = 0;
  /** Coverpoint variable to store the status if bvalid is deasserted after arready. */
  bit cov_bvalid_arready = 0;
  /** Coverpoint variable to store the status if bvalid is deasserted after wready. */
  bit cov_bvalid_wready = 0;
  /** Coverpoint variable to store the status if bvalid is deasserted after rvalid. */
  bit cov_bvalid_rvalid = 0;

  /** Coverpoint variable to store the status if awvalid is deasserted after awready. */
  bit cov_awvalid_awready = 0;
  /** Coverpoint variable to store the status if awvalid is deasserted after wready. */
  bit cov_awvalid_wready = 0;
  /** Coverpoint variable to store the status if awvalid is deasserted after rvalid. */
  bit cov_awvalid_rvalid = 0;
  /** Coverpoint variable to store the status if awvalid is deasserted after bvalid. */
  bit cov_awvalid_bvalid = 0;
  /** Coverpoint variable to store the status if wvalid is deasserted after awready. */
  bit cov_wvalid_awready = 0;
  /** Coverpoint variable to store the status if wvalid is deasserted after wready. */
  bit cov_wvalid_wready = 0;
  /** Coverpoint variable to store the status if wvalid is deasserted after rvalid. */
  bit cov_wvalid_rvalid = 0;
  /** Coverpoint variable to store the status if wvalid is deasserted after bvalid. */
  bit cov_wvalid_bvalid = 0;
  /** Coverpoint variable to store the status if rready is deasserted after awready. */
  bit cov_rready_awready = 0;
  /** Coverpoint variable to store the status if rready is deasserted after wready. */
  bit cov_rready_wready = 0;
  /** Coverpoint variable to store the status if rready is deasserted after rvalid. */
  bit cov_rready_rvalid = 0;
  /** Coverpoint variable to store the status if rready is deasserted after bvalid. */
  bit cov_rready_bvalid = 0;
  /** Coverpoint variable to store the status if bready is deasserted after awready. */
  bit cov_bready_awready = 0;
  /** Coverpoint variable to store the status if bready is deasserted after wready. */
  bit cov_bready_wready = 0;
  /** Coverpoint variable to store the status if bready is deasserted after rvalid. */
  bit cov_bready_rvalid = 0;
  /** Coverpoint variable to store the status if bready is deasserted after bvalid. */
  bit cov_bready_bvalid = 0;

  /** Coverpoint variable to store the status if awready is deasserted after awvalid. */
  bit cov_awready_and_awvalid = 0;                                              
  /** Coverpoint variable to store the status if awready is deasserted after wvalid. */
  bit cov_awready_and_wvalid = 0;                                               
  /** Coverpoint variable to store the status if awready is deasserted after rvalid. */
  bit cov_awready_and_rvalid = 0;                                               
  /** Coverpoint variable to store the status if awready is deasserted after bvalid. */
  bit cov_awready_and_bvalid = 0;                                               
  /** Coverpoint variable to store the status if wready is deasserted after awvalid. */
  bit cov_wready_and_awvalid = 0;                                               
  /** Coverpoint variable to store the status if wready is deasserted after wvalid. */
  bit cov_wready_and_wvalid = 0;                                                
  /** Coverpoint variable to store the status if wready is deasserted after rready. */
  bit cov_wready_and_rready = 0;                                                
  /** Coverpoint variable to store the status if wready is deasserted after bready. */
  bit cov_wready_and_bready = 0;                                                
  /** Coverpoint variable to store the status if rvalid is deasserted after awready. */
  bit cov_rvalid_and_awready = 0;                                               
  /** Coverpoint variable to store the status if rvalid is deasserted after wready. */
  bit cov_rvalid_and_wready = 0;                                                
  /** Coverpoint variable to store the status if rvalid is deasserted after rready. */
  bit cov_rvalid_and_rready = 0;                                                
  /** Coverpoint variable to store the status if rvalid is deasserted after bready. */
  bit cov_rvalid_and_bready = 0;                                                
  /** Coverpoint variable to store the status if bvalid is deasserted after awready. */
  bit cov_bvalid_and_awready = 0;                                               
  /** Coverpoint variable to store the status if bvalid is deasserted after wready. */
  bit cov_bvalid_and_wready = 0;                                                
  /** Coverpoint variable to store the status if bvalid is deasserted after rready. */
  bit cov_bvalid_and_rready = 0;                                                
  /** Coverpoint variable to store the status if bvalid is deasserted after bready. */
  bit cov_bvalid_and_bready = 0;

  /** Flags used to ensure cover bins hit for required number of times */
  protected bit cov_AWVALID_to_AWREADY_Delay_flag = 1'b0;
  protected bit cov_ARVALID_to_ARREADY_Delay_flag = 1'b0;
  protected bit cov_ACVALID_to_ACREADY_Delay_flag = 1'b0;
  protected bit cov_ACVALID_to_CRVALID_Delay_flag = 1'b0;
  protected bit cov_CDVALID_to_CDREADY_Delay_flag = 1'b0;
  protected bit cov_CRVALID_to_CRREADY_Delay_flag = 1'b0;
  protected bit cov_WVALID_to_WREADY_Delay_flag = 1'b0;
  protected bit cov_TVALID_to_TREADY_Delay_flag = 1'b0;
  protected bit cov_TVALID_Delay_flag = 1'b0;
  protected bit cov_TREADY_Delay_flag = 1'b0;
  protected bit cov_RVALID_to_RREADY_Delay_flag = 1'b0;
  protected bit cov_BVALID_to_BREADY_Delay_flag = 1'b0;
  protected bit cov_AWVALID_to_prev_AWVALID_Delay_flag = 1'b0;
  protected bit cov_WVALID_to_prev_WVALID_Delay_flag = 1'b0;
  protected bit cov_TVALID_to_prev_TVALID_Delay_flag = 1'b0;  
  protected bit cov_AWVALID_to_first_WVALID_Delay_flag = 1'b0;
  protected bit cov_last_wdata_handshake_to_BVALID_Delay_flag = 1'b0;
  protected bit cov_ARVALID_to_prev_ARVALID_Delay_flag = 1'b0;
  protected bit cov_RVALID_to_prev_RVALID_Delay_flag = 1'b0;
  protected bit cov_ARVALID_to_first_RVALID_Delay_flag = 1'b0;
  protected bit cov_xact_type_flag = 1'b0;
  protected bit cov_burst_type_flag = 1'b0;
`ifdef SVT_ACE5_ENABLE
  protected bit cov_stream_id_flag = 1'b0;
  protected bit cov_sub_stream_id_flag = 1'b0;
  protected bit cov_secure_or_non_secure_stream_flag = 1'b0;
  protected bit cov_sub_stream_id_valid_flag = 1'b0;
  protected bit cov_stash_nid_flag = 1'b0;
  protected bit cov_stash_lpid_flag = 1'b0;
  protected bit cov_stash_nid_valid_flag = 1'b0;
  protected bit cov_stash_lpid_valid_flag = 1'b0;
  protected bit cov_atomic_comp_xact_type_flag = 1'b0;
  protected bit cov_atomic_comp_op_type_flag = 1'b0;
  protected bit cov_atomic_noncomp_xact_type_flag = 1'b0;
  protected bit cov_atomic_noncomp_op_type_flag = 1'b0;
  protected bit cov_coherent_stash_xact_type_flag = 1'b0;
  protected bit cov_endian_flag = 1'b0;
  protected bit cov_atomic_burst_type_flag = 1'b0;
  protected bit cov_atomic_comp_burst_size_flag = 1'b0;
  protected bit cov_atomic_non_comp_burst_size_flag = 1'b0;
  protected bit cov_chunk_burst_type_flag = 1'b0;
  protected bit cov_chunk_burst_size_flag = 1'b0;
  protected bit cov_chunk_length_flag = 1'b0;
  protected bit cov_chunkstrb_flag = 1'b0;
  protected bit cov_chunknum_flag = 1'b0;
`endif  
  protected bit cov_burst_length_flag = 1'b0;
  protected bit cov_qos_type_flag = 1'b0;
  protected bit cov_addr_flag = 1'b0;
  protected bit cov_bresp_flag = 1'b0;
  protected bit cov_rresp_flag = 1'b0;
  protected bit cov_wstrb_flag = 1'b0;
  protected bit cov_burst_size_flag = 1'b0;
  protected bit cov_atomic_type_flag = 1'b0;
  protected bit cov_cache_type_flag = 1'b0;
  protected bit cov_prot_type_flag = 1'b0;
  protected bit cov_exceptions_flag = 1'b0;
  protected bit cov_region_type_flag = 1'b0;
  protected bit cov_data_user_flag = 1'b0;
  protected bit cov_addr_user_flag = 1'b0;
  protected bit cov_resp_user_flag = 1'b0;
  protected bit is_addr_4kb_boundary_cross_flag = 1'b0;
  protected bit barrier_outstanding_xact_flag = 1'b0;
  protected bit total_outstanding_xact_flag = 1'b0;
  protected bit outstanding_write_xact_flag = 1'b0;
  protected bit outstanding_read_xact_flag = 1'b0;
  protected bit read_data_interleave_flag = 1'b0;
  protected bit write_data_interleave_flag = 1'b0;
  protected bit stream_data_interleave_flag = 1'b0;
  protected bit cov_coherent_xact_type_flag = 1'b0;
  protected bit cov_barrier_type_flag = 1'b0;
  protected bit cov_domain_type_flag = 1'b0;
  protected bit cov_coherent_resp_type_flag = 1'b0;
  protected bit cov_snoop_xact_type_flag = 1'b0;
  protected bit cov_snoop_burst_length_flag = 1'b0;
  protected bit cov_coherent_rresp_flag = 1'b0;
  protected bit cov_snoop_resp_flag = 1'b0;
  protected bit cov_snoop_prot_type_flag = 1'b0;
  protected bit cov_snoop_addr_flag = 1'b0;
  protected bit cov_ardvm_message_flag = 1'b0;
  protected bit cov_acdvm_message_flag = 1'b0;
  protected reg [6:0] addr_offset_coverpoint;
  protected reg [63:0] dvm_araddr_firstpart_msbto32_coverpoint;
  protected reg [63:0] snoop_dvm_araddr_firstpart_msbto32_coverpoint;
  protected reg [63:0] dvm_araddr_secondpart_coverpoint;
  protected reg [63:0] snoop_dvm_araddr_secondpart_coverpoint;
  protected reg [7:0] dvm_araddr_firstpart_va_asid_coverpoint;
  protected reg [7:0] snoop_dvm_araddr_firstpart_va_asid_coverpoint;
  protected reg [5:0] dvm_addr_mode_bits_coverpoint;
  protected reg [5:0] snoop_dvm_addr_mode_bits_coverpoint;
  protected reg [7:0] dvm_message_virt_inst_cache_invl_bits_coverpoint;
  protected reg [7:0] snoop_dvm_message_virt_inst_cache_invl_bits_coverpoint;
  protected reg [5:0] dvm_message_phy_inst_cache_invl_bits_coverpoint;
  protected reg [5:0] snoop_dvm_message_phy_inst_cache_invl_bits_coverpoint;
  protected reg [7:0] dvm_araddr_firstpart_va_vmid_coverpoint;
  protected reg [7:0] snoop_dvm_araddr_firstpart_va_vmid_coverpoint;
  protected svt_axi_transaction dvm_multipart_xact_q[$];
  protected svt_axi_snoop_transaction snoop_dvm_multipart_xact_q[$];
  protected bit cov_initial_cache_line_state_flag = 1'b0;
  protected bit cov_final_cache_line_state_flag = 1'b0;
  protected bit cov_snoop_initial_cache_line_state_flag = 1'b0;
  protected bit cov_snoop_final_cache_line_state_flag = 1'b0;
  protected bit cov_dvm_araddr_firstpart_width32_flag = 1'b0;
  protected bit cov_dvm_araddr_firstpart_width24_flag = 1'b0;
  protected bit cov_dvm_araddr_firstpart_width16_flag = 1'b0;
  protected bit cov_snoop_dvm_araddr_firstpart_width16_flag = 1'b0;
  protected bit cov_snoop_dvm_araddr_firstpart_width32_flag = 1'b0;
  protected bit cov_snoop_dvm_araddr_firstpart_width24_flag = 1'b0;
  protected bit cov_snoop_dvm_araddr_firstpart_width12_flag = 1'b0;
  protected bit cov_snoop_dvm_araddr_firstpart_width8_flag = 1'b0;
  protected bit cov_dvm_araddr_firstpart_width12_flag = 1'b0;
  protected bit cov_dvm_araddr_firstpart_width8_flag = 1'b0;
  protected bit cov_dvm_araddr_secondpart_width64_flag =1'b0;
  protected bit cov_dvm_araddr_secondpart_width56_flag =1'b0;
  protected bit cov_dvm_araddr_secondpart_width48_flag =1'b0;
  protected bit cov_dvm_araddr_secondpart_width44_flag =1'b0;
  protected bit cov_dvm_araddr_secondpart_width40_flag =1'b0;
  protected bit cov_dvm_araddr_secondpart_width32_flag =1'b0;
  protected bit cov_snoop_dvm_araddr_secondpart_width64_flag =1'b0;
  protected bit cov_snoop_dvm_araddr_secondpart_width56_flag =1'b0;
  protected bit cov_snoop_dvm_araddr_secondpart_width48_flag =1'b0;
  protected bit cov_snoop_dvm_araddr_secondpart_width44_flag =1'b0;
  protected bit cov_snoop_dvm_araddr_secondpart_width40_flag =1'b0;
  protected bit cov_snoop_dvm_araddr_secondpart_width32_flag =1'b0;
  protected bit cov_dvm_araddr_viraddr_or_vmid_flag = 1'b0;
  protected bit cov_addr_6_bit_flag = 1'b1;
  protected bit cov_snoop_dvm_araddr_viraddr_or_vmid_flag = 1'b0;
  protected bit cov_dvm_araddr_viraddr_or_asid_flag = 1'b0;
  protected bit cov_snoop_dvm_araddr_viraddr_or_asid_flag = 1'b0;
  protected bit cov_snoop_addr_6_bit_flag = 1'b1;
  protected bit cov_ACVALID_to_prev_ACVALID_Delay_flag = 1'b0;
  //protected bit cov_CRVALID_to_prev_CRVALID_Delay_flag = 1'b0;
  protected bit cov_CDVALID_to_prev_CDVALID_Delay_flag = 1'b0;

  protected bit out_of_order_read_response_depth_flag = 1'b0;
  protected bit out_of_order_write_response_depth_flag = 1'b0;

  protected bit cov_stream_xact_type_flag = 1'b0;
  protected bit cov_stream_tid_flag = 1'b0;
  protected bit cov_stream_tdest_flag = 1'b0;

  `ifdef SVT_VMM_TECHNOLOGY
  static vmm_log log = new( "svt_axi_port_monitor_def_cov_data_callback", "CLASS" );
  `endif

 
 /** Event used to trigger read xacts with same ID that are targeted to different slaves covergroup for sampling. */
  event cov_outstanding_read_with_same_id_to_different_slaves_sample_event;

 /** Event used to trigger write xacts with same ID that are targeted to different slaves covergroup for sampling. */
  event cov_outstanding_write_with_same_id_to_different_slaves_sample_event;

 /** Event used to trigger xacts on AR or AW channel can be stalled for snoop xacts on AC channel covergroup for sampling. */
  event cov_ar_aw_stalled_for_ac_channel_sample_event;

 /** Event used to trigger xacts followed the lanuch of nonshareable barrier can be any domain covergroup for sampling. */
  event cov_xact_domain_after_nonshareable_barrier_sample_event;

 /** Event used to trigger xacts followed the lanuch of innershareable barrier can be any domain covergroup for sampling. */
  event cov_xact_domain_after_innershareable_barrier_sample_event;

 /** Event used to trigger xacts followed the lanuch of outershareable barrier can be any domain covergroup for sampling. */
  event cov_xact_domain_after_outershareable_barrier_sample_event;

 /** Event used to trigger xacts followed the lanuch of systemshareable barrier can be any domain covergroup for sampling. */
  event cov_xact_domain_after_systemshareable_barrier_sample_event;

 /** Event used to trigger xacts followed the lanuch of barrier can get response in any order covergroup for sampling. */
  event cov_xact_ordering_after_barrier_sample_event;

  /** Event used to trigger trans_master_back_to_back_write_ordering coverage */
  event cov_master_back_to_back_write_ordering_event;

  /** Event used to trigger trans_master_write_after_read_ordering */
  event cov_master_write_after_read_ordering_event;

  /** Event used to trigger trans_master_concurrent_coherent_exclusive_access */
  event cov_coherent_exclusive_read_access_event;

  /** Event used to trigger trans_master_coherent_unmatched_excl_access */
  event cov_coherent_unmatched_excl_access_event;
        
  /** Event used to trigger trans_master_num_outstanding_dvm_syncs */
  event cov_snoop_dvm_sync_event;
          
  /** Event to trigger trans_master_barrier_id_reuse_for_non_barrier */
  event cov_barrier_id_reuse_for_non_barrier_event;
 
 /** flag to indicate if there is write transactions accpted by Slave after 256 outstanding barrier transaction occur. */
  protected int non_barrier_after_256_outstanding_barrier= 0;

/** variable to store if there are active read transactions with same ID that are targeted to different slaves.
 * - if value == 1; yes, there are active read outstanding transactions with same ID that are targeted to different slaves
 * - if value ==0; no, there are no active read outstanding transactions with same ID that are targeted to different slaves
 * .
 */
  protected int outstanding_read_with_same_id_to_different_slaves =0;

/** variable to store if there are active write transactions with same ID that are targeted to different slaves.
 * - if value == 1; yes, there are active write outstanding transactions with same ID that are targeted to different slaves
 * - if value ==0; no, there are no active write outstanding transactions with same ID that are targeted to different slaves
 * .
 */
  protected int outstanding_write_with_same_id_to_different_slaves =0; 
 
/** variable to store if there are AR/AW xacts stalled for AC operation. 
 *  - if value=='hff, there is no AW/AR xcat stalled for snoop,
 *  - otherwise, there is AR/AW xact stalled for snoop, the value definition is as below:
 *  .
 */
  protected int ar_aw_stalled_for_ac_channel =16'hff;


/** flag to indicate the domain type of current read barrier. 
 * - if value == 0,1,2,3,there is active barriers(not complete yet)
 * - if value ==4'hf, it indicates the barrier completes
 * .
 */
  protected int current_read_barrier_domain=4'hf; 

/** flag to indicate the domain type of current write barrier. */
  protected int current_write_barrier_domain=4'hf;

/** variable to store the domain type of xcats followed by the launch of nonshareable barrier.
 * - if value == 0,1,2,3, it means non/inner/outer/system repectively on read channel
 * - if value == 4,5,6,7, it means non/inner/outer/system repectively on write channel
 * - if value==4'hf, it indicates there is no transactions followed
 * .
 */
  protected int xact_domain_after_nonshareable_barrier=4'hf;

/** variable to store the domain type of xcats followed by the launch of innershareable barrier.*/
  protected int xact_domain_after_innershareable_barrier=4'hf;

/** variable to store the domain type of xcats followed by the launch of outershareable barrier.*/
  protected int xact_domain_after_outershareable_barrier=4'hf;

/** variable to store the domain type of xcats followed by the launch of systemshareable barrier.*/
  protected int xact_domain_after_systemshareable_barrier=4'hf;

/** flag to indicate if the current read barrier is active. */
  protected int current_read_barrier_is_active=0;

/** flag to indicate if the current write barrier is active. */
  protected int current_write_barrier_is_active=0;

/** flag to indicate if there is read barrier. */
  protected int there_is_read_barrier=0;

/** flag to indicate if there is write barrier. */
  protected int there_is_write_barrier=0;

/** varaible to store the addr valid assertion cycle of read barrier. */
  protected int current_read_barrier_addr_valid_assertion_cycle=0;

/** varaible to store the addr valid assertion cycle of write barrier. */
  protected int current_write_barrier_addr_valid_assertion_cycle=0;

/** variable to store the response ordering of transactions followed by the launch of barrier.
  * - if value==1, it indicates the transaction is completed after the barrier response(in-order)on read channel
  * - if value==0, it indicates the transaction is completed before the barrier response(out-of-order)on read channel
  * - if value==3, it indicates the transaction is completed after the barrier response(in-order)on write channel
  * - if value==2, it indicates the transaction is completed before the barrier response(out-of-order)on write channel
  * - if value=='hf, there is no transaction followed after the launch of barrier and before the barrier response
  * .
 */ 
  protected int xact_ordering_after_barrier=4'hf;

  /** variable to store the ordering information of back-to-back write transactions
    * 0: Back to back write with same id
    */
  protected int back_to_back_write_ordering = 0;

  /** variable to store the ordering information of write and read transactions
    * 0: Write after read with the write completing first
    * 1: Write after read with the read completing first
    */
  protected int write_after_read_ordering = 0;

  /** variable to store the read transaction type information 
    * when there is snoop to same address
    */
  protected int read_xact_to_same_address_as_snoop = 0;

  /** variable to store the write transaction type information 
    * when there is snoop to same address
    */
  protected int write_xact_type_to_same_addr_as_snoop = 0;

  /** variable to store the number of outstanding coherent exclusive accesses on different IDs */
  protected int num_coherent_excl_access_threads = 0;

  /** variable identifying the type of unmatched exlcusive access:
    * 0: unmatched exlcusive write
    * 1: unmatched exclusive read
    */
  protected int coherent_unmatched_excl_access_type = 0;

  /** Identifies number of outstanding dvm syncs */
  protected int num_outstanding_dvm_syncs = 0;

  /** Number of non-barrier transactions that reuse IDs used in barrier */
  protected int num_barrier_id_reuse = 0;

  /** Identifies whether snoop data transfer was initiated with readunique in clean cache state */
  protected bit readunique_snoop_resp_datatransfer_with_clean_cacheline = 0;

  /** Outstanding coherent exlcusive read accesses */
  protected svt_axi_transaction outstanding_coherent_exclusive_read_access_q[$];

  /** Queue of ids used in barrier */
  protected bit[`SVT_AXI_MAX_ID_WIDTH-1:0] barrier_ids[$];

  /** Handle to write transaction to same address as snoop */
  protected svt_axi_transaction write_xact_to_same_addr_as_snoop;

  /** Number of dvm enabled masters */
  protected int num_dvm_enabled_masters = 1;

  /** Mapping of coherent to snoop transactions */
  int coh_and_snp_association;//MSB--coherent,LSB--snoop
  
  /** Coverpoint variable used to store the concurrent readunique/cleanunique access */
  int concurrent_readunique_cleanunique;
  
  /** Coverpoint variable use to hold the value of coherent_xact_type for covergroup trans_master_ace_concurrent_overlapping_coherent_xacts  */
  svt_axi_transaction::coherent_xact_type_enum coherent_xact_on_port1;

  /** Coverpoint variable use to hold the value of coherent_xact_type for covergroup trans_master_ace_concurrent_overlapping_coherent_xacts */
  svt_axi_transaction::coherent_xact_type_enum coherent_xact_on_port2;
  
  /** Coverpoint variable used to store the master transaction received in
   * interconnect_generated_dirty_data_write_detected callback */ 
  svt_axi_transaction master_xact_of_ic_dirty_data_write;
  
  /** Coverpoint and Enum used to store snoop and memory read timing for
    * covergroup trans_master_ace_snoop_and_memory_returns_data.
    */
  typedef enum bit[2:0] {
    SNOOP_WITHOUT_MEMORY_READ = 3'b000,
    SNOOP_BEFORE_MEMORY_READ = 3'b001,
    SNOOP_ALONG_WITH_MEMORY_READ = 3'b010,
    SNOOP_AFTER_MEMORY_READ = 3'b011,
    SNOOP_RETURNS_DATA_AND_MEMORY_NOT_RETURNS_DATA = 3'b100
  } snoop_and_memory_read_timing_enum;

  snoop_and_memory_read_timing_enum snoop_and_memory_read_timing = SNOOP_WITHOUT_MEMORY_READ;

  /** Coverpoint variable used to store the master transaction received in
    * master_xact_fully_associated_to_slave_xacts callback
    */
  svt_axi_transaction fully_correlated_master_xact;
  
  /** Indicates if an xact from other master when barrier is in progress is detected */
  bit is_xacts_from_other_master_during_barrier_covered = 0;
  
  /** Property used by system_ace_barrier_response_with_outstanding_xacts */
  svt_axi_transaction completed_barrier_xact;
  
  /** Coverpoint variable used to store the overlapping coherent transaction */
  int store_overlap_coh_xact;
  
  /** Coverpoint variable used to store the overlapping coherent transaction */
  int no_cached_copy_overlap_coh_xact;  

  /** Name of the agent/group that this port is instantiated in */
  string requester_name;



//----------------------------------------------------------------------------
 /**
   * Calls buil-in sample function for each corresponding covergroups
   * in order to collect coverage for read transaction parameters.
   */
  extern virtual function void cov_sample_read_xact_parameters();
//----------------------------------------------------------------------------
 /**
   * Calls buil-in sample function for each corresponding covergroups
   * in order to collect coverage for write transaction parameters.
   */
  extern virtual function void cov_sample_write_xact_parameters();
//----------------------------------------------------------------------------
 /**
   * Calls buil-in sample function for each corresponding covergroups
   * in order to collect coverage for axi4 stream transaction parameters.
   */
  extern virtual function void cov_sample_axi4_stream_xact_parameters();
//----------------------------------------------------------------------------
 /**
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoup read_outstanding_xact_same_arid_cache_modifiable_bit
   * and read_outstanding_xact_diff_arid_cache_modifiable_bit
   */
  extern virtual function void cov_sample_read_outstanding_xact_cache_modifiable_bit();
//----------------------------------------------------------------------------
 /**
   * Calls built-in sample function for corresponding covergroup
   * in order to collect coverage for covergoup read_outstanding_xact_diff_arid_device_cacheable_bit
   */  
  extern virtual function void cov_sample_read_outstanding_xact_device_cacheable_bit();
//----------------------------------------------------------------------------
 /**
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for dvm_firstpart_secondpart_covergroups 
   */
  extern virtual function void cov_sample_dvm_multipart_xact_covergroups();

//----------------------------------------------------------------------------
 /**
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for snoop dvm_firstpart_secondpart_covergroups 
   */
  extern virtual function void cov_sample_snoop_dvm_multipart_xact_covergroups();

//----------------------------------------------------------------------------
 /**
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoup write_outstanding_xact_same_arid_cache_modifiable_bit
   * and write_outstanding_xact_diff_arid_cache_modifiable_bit
   */
  extern virtual function void cov_sample_write_outstanding_xact_cache_modifiable_bit();

//----------------------------------------------------------------------------
 /**
   * Calls built-in sample function for corresponding covergroup
   * in order to collect coverage for covergoup write_outstanding_xact_diff_awid_device_cacheable_bit
   */  
  extern virtual function void cov_sample_write_outstanding_xact_device_cacheable_bit();

//----------------------------------------------------------------------------
 /**
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoup trans_axi_num_outstanding_xacts_with_same_arid 
   * and trans_axi_num_outstanding_xacts_with_diff_arid 
   */
  extern virtual function void cov_sample_read_outstanding_xact();
 /**
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoups trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid
   * and trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid
   */
  extern virtual function void cov_sample_dvm_tlb_invalidate_outstanding_xact();  
 /**
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoup trans_ace_num_outstanding_snoop_xacts
   */
  extern virtual function void cov_sample_snoop_outstanding_xact(); 

//----------------------------------------------------------------------------
 /**
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for snoop dvm covergroups 
   */
  extern virtual function void cov_sample_snoop_dvm_xact_covergroups(); 
  
//----------------------------------------------------------------------------
  /**
   * Coverage sample event functions.
   *
   * Following functions triggers sample event in order to collect coverage for covergroup signal_master_valid_ready_dependency.
   */  
  extern virtual function void cov_sample_awvalid_wvalid_dependency();  
  extern virtual function void cov_sample_awvalid_rready_dependency();  
  extern virtual function void cov_sample_awvalid_bready_dependency();  
  extern virtual function void cov_sample_wvalid_awvalid_dependency();  
  extern virtual function void cov_sample_wvalid_rready_dependency();  
  extern virtual function void cov_sample_wvalid_bready_dependency();  
  extern virtual function void cov_sample_rready_awvalid_dependency();
  extern virtual function void cov_sample_rready_wvalid_dependency();  
  extern virtual function void cov_sample_rready_bready_dependency();  
  extern virtual function void cov_sample_bready_awvalid_dependency();  
  extern virtual function void cov_sample_bready_wvalid_dependency();  
  extern virtual function void cov_sample_bready_rready_dependency(); 
//----------------------------------------------------------------------------
  /**
   * Coverage sample event functions.
   *
   * Following functions triggers sample event in order to collect coverage for covergroup signal_slave_valid_ready_dependency.
   */  
  extern virtual function void cov_sample_wready_arready_dependency(); 
  extern virtual function void cov_sample_wready_rvalid_dependency(); 
  extern virtual function void cov_sample_wready_bvalid_dependency(); 
  extern virtual function void cov_sample_arready_wready_dependency(); 
  extern virtual function void cov_sample_arready_rvalid_dependency(); 
  extern virtual function void cov_sample_arready_bvalid_dependency(); 
  extern virtual function void cov_sample_rvalid_arready_dependency(); 
  extern virtual function void cov_sample_rvalid_wready_dependency(); 
  extern virtual function void cov_sample_rvalid_bvalid_dependency(); 
  extern virtual function void cov_sample_bvalid_arready_dependency(); 
  extern virtual function void cov_sample_bvalid_wready_dependency(); 
  extern virtual function void cov_sample_bvalid_rvalid_dependency();
//----------------------------------------------------------------------------
  /**
   * Coverage sample event functions.
   *
   * Following functions triggers sample event in order to collect coverage for covergroup signal_master_slave_valid_ready_dependency.
   */
  extern virtual function void cov_sample_awvalid_awready_dependency(); 
  extern virtual function void cov_sample_awvalid_wready_dependency(); 
  extern virtual function void cov_sample_awvalid_rvalid_dependency(); 
  extern virtual function void cov_sample_awvalid_bvalid_dependency(); 
  extern virtual function void cov_sample_wvalid_awready_dependency(); 
  extern virtual function void cov_sample_wvalid_wready_dependency(); 
  extern virtual function void cov_sample_wvalid_rvalid_dependency(); 
  extern virtual function void cov_sample_wvalid_bvalid_dependency(); 
  extern virtual function void cov_sample_rready_awready_dependency(); 
  extern virtual function void cov_sample_rready_wready_dependency(); 
  extern virtual function void cov_sample_rready_rvalid_dependency(); 
  extern virtual function void cov_sample_rready_bvalid_dependency(); 
  extern virtual function void cov_sample_bready_awready_dependency(); 
  extern virtual function void cov_sample_bready_wready_dependency(); 
  extern virtual function void cov_sample_bready_rvalid_dependency(); 
  extern virtual function void cov_sample_bready_bvalid_dependency();
//----------------------------------------------------------------------------
  /**
   * Coverage sample event functions.
   *
   * Following functions triggers sample event in order to collect coverage for covergroup signal_slave_master_valid_ready_dependency.
   */
  extern virtual function void cov_sample_awready_and_awvalid_dependency(); 
  extern virtual function void cov_sample_awready_and_wvalid_dependency(); 
  extern virtual function void cov_sample_awready_and_rvalid_dependency(); 
  extern virtual function void cov_sample_awready_and_bvalid_dependency(); 
  extern virtual function void cov_sample_wready_and_awvalid_dependency(); 
  extern virtual function void cov_sample_wready_and_wvalid_dependency(); 
  extern virtual function void cov_sample_wready_and_rready_dependency(); 
  extern virtual function void cov_sample_wready_and_bready_dependency(); 
  extern virtual function void cov_sample_rvalid_and_awready_dependency(); 
  extern virtual function void cov_sample_rvalid_and_wready_dependency(); 
  extern virtual function void cov_sample_rvalid_and_rready_dependency(); 
  extern virtual function void cov_sample_rvalid_and_bready_dependency(); 
  extern virtual function void cov_sample_bvalid_and_awready_dependency(); 
  extern virtual function void cov_sample_bvalid_and_wready_dependency(); 
  extern virtual function void cov_sample_bvalid_and_rready_dependency(); 
  extern virtual function void cov_sample_bvalid_and_bready_dependency(); 
//----------------------------------------------------------------------------
 /**
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoup trans_axi_num_outstanding_xacts_with_same_awid 
   * and trans_axi_num_outstanding_xacts_with_diff_awid 
   */
  extern virtual function void cov_sample_write_outstanding_xact();  
  //----------------------------------------------------------------------------
  /**
   * Callback issued when a Port Activity Transaction is ready at the monitor.
   * The coverage needs to extend this method as we want to get the details of
   * the transaction, at the end of the transaction.
   *
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_transaction.
   */
  //----------------------------------------------------------------------------  
  extern virtual function void pre_output_port_put(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);
   
  extern virtual function void new_snoop_transaction_started(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);
  
  /** Called when a new idle snoop channel toggles acwakeup assertion is observed on the port */
  extern virtual function void new_snoop_channel_acwakeup_toggle_started(svt_axi_port_monitor axi_monitor, int assert_delay);
  
  /** Called when a new idle snoop channel toggles acwakeup deassertion is observed on the port */
  extern virtual function void new_snoop_channel_acwakeup_toggle_ended(svt_axi_port_monitor axi_monitor, int deassert_delay);

  /** Called when a new idle snoop channel toggles awakeup assertion is observed on the port */
  extern virtual function void new_snoop_channel_awakeup_toggle_started(svt_axi_port_monitor axi_monitor, int assert_delay);
  
  /** Called when a new idle snoop channel toggles awakeup deassertion is observed on the port */
  extern virtual function void new_snoop_channel_awakeup_toggle_ended(svt_axi_port_monitor axi_monitor, int deassert_delay);

  //----------------------------------------------------------------------------

  /** 
  * Called when a new transaction is observed on the port 
   * 
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_transaction.
   */
 //----------------------------------------------------------------------------  
  extern virtual function void new_transaction_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);
 
 /** 
   * Called whenever an ace dvm snoop_valid coherent_valid overlap realated case need to cover 
   * 
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_transaction.
   */
 //----------------------------------------------------------------------------  
  extern virtual function void snoop_address_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);

 /** 
   * Called whenever an ace dvm overlap snoop_resp coherent_valid overlap realated case need to cover 
   * 
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_transaction.
   */
  //----------------------------------------------------------------------------
  extern virtual function void snoop_resp_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);

 //----------------------------------------------------------------------------
  /** 
  * Called when a transaction ends
   * 
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_transaction.
  */
 //----------------------------------------------------------------------------  
  extern virtual function void transaction_ended(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);

  `ifndef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Callback issued by component to allow callbacks to initiate activities.
   * This callback is issued during the run phase.
   *
   * @param component A reference to the component object issuing this callback.
   */
  extern virtual function void startup(`SVT_XVM(component) component);
`else
  extern virtual function void start(svt_xactor xactor);
  
`endif


//----------------------------------------------------------------------------
  /** 
   * Called when RVALID is asserted
   * 
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_transaction.
  */
 //----------------------------------------------------------------------------  
  extern virtual function void read_data_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);

  //----------------------------------------------------------------------------
  /** 
   * Called when TVALID is asserted
   * 
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_transaction.
  */
 //----------------------------------------------------------------------------  
  extern virtual function void stream_transfer_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);

  //----------------------------------------------------------------------------
  /** 
   * Called when WVALID is asserted
   * 
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_transaction.
  */
 //----------------------------------------------------------------------------
  extern virtual function void write_data_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);
  extern virtual function void write_resp_phase_started(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);

  //----------------------------------------------------------------------------
  /**
   * Callback issued when a Snoop Activity Transaction is ready at the monitor.
   * The coverage needs to extend this method as we want to get the details of
   * the transaction, at the end of the transaction.
   *
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_snoop_transaction.
   */
  //----------------------------------------------------------------------------
  extern virtual function void pre_snoop_output_port_put(svt_axi_port_monitor axi_monitor, svt_axi_snoop_transaction item);

  //----------------------------------------------------------------------------
  /**
   * Called when read address handshake is complete, that is, when ARVALID and ARREADY are asserted.
   * Extension of this method in the default coverage callback class is used for signal coverage of read address channel signals. 
   *
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_transaction.
   */
  //----------------------------------------------------------------------------  
  extern virtual function void read_address_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);


  //----------------------------------------------------------------------------
  /**
   * Called when write address handshake is complete, that is, when AWVALID and AWREADY are asserted.
   * Extension of this method in the default coverage callback class is used for signal coverage of write address channel signals. 
   *
   * @param axi_monitor A reference to the AXI Monitor transactor instance that
   * issued this callback.
   *
   * @param item A reference to the svt_axi_transaction.
   */
  //----------------------------------------------------------------------------  
  extern virtual function void write_address_phase_ended(svt_axi_port_monitor axi_monitor, svt_axi_transaction item);

  /** @cond PRIVATE */
  /**
   * Called when a read/write transaction is added to outstanding xact queue to trigger
   * corresponding covergrop events:
   * - if there are multiple outstanding read transactions that has same ID, but 
   *   targeted to different slaves
   * - if there are multiple outstanding write transactions that has same ID, but 
   *   targeted to different slaves
   * .
   * @param xact Current transaction under the context
   */
  extern virtual function void evaluate_outstanding_with_same_id_to_different_slaves(svt_axi_transaction xact);
  //----------------------------------------------------------------------------  
  /**
   * Indicates:
   * - if there are multiple outstanding read transactions that has same ID, but 
   *   targeted to different slaves
   * - if there are multiple outstanding write transactions that has same ID, but 
   *   targeted to different slaves
   * .
   * @param xact Current transaction under the context
   * @param input_queue Transaction queue under the context
   */
  extern virtual function bit is_outstanding_with_same_id_to_different_slaves(svt_axi_transaction xact, svt_axi_transaction input_queue[$]);
  //----------------------------------------------------------------------------
  /**
   * Called when four_state_rd_wr_queue is filled with four RD/WR transactions,to trigger
   * corresponding covergrop events
   */
  extern virtual function void trigger_four_state_rd_wr_event();
  //----------------------------------------------------------------------------
  /**
   * Called when four_excl_normal_seq_queue is filled with four Exclusive/Normal transactions,to trigger
   * corresponding covergrop events
   */
  extern virtual function void trigger_four_excl_normal_seq_event();
  
  //------------------------------------------------------------------------------
  /**
    * Called to evaluate if there are back to back writes from the same port with same ID
    */
  extern function void evaluate_back_to_back_write_with_same_id(svt_axi_transaction xact);
  //------------------------------------------------------------------------------
  /**
    * Called to evaluate if there are reads completing first in a situation where there is a read transacton followed by a write transaction
    */
  extern function void evaluate_read_completing_first_in_write_after_read(svt_axi_transaction read_xact);
  //------------------------------------------------------------------------------
  /**
    * Called to evaluate if there are writese completing first in a situation where there is a read transacton followed by a write transaction
    */
  extern function void evaluate_write_completing_first_in_write_after_read(svt_axi_transaction write_xact);

  /**
    * Called to evaluate if there is a snoop transaction to the same address as a read transaction
    */
  extern virtual function void evaluate_snoop_to_same_address_as_read_xact(svt_axi_snoop_transaction snoop_xact);

  /**
    * Called to evaluate if there is a snoop transaction to the same address as a write transaction
    * @param snoop_xact Handle to the snoop transaction
    * @param is_at_snoop_addr_phase Indicates if this is called in the snoop_addr_phase_started or ended callback
    */
  extern virtual function void evaluate_snoop_to_same_address_as_write_xact(svt_axi_snoop_transaction snoop_xact, bit is_at_snoop_addr_phase = 0);

  /**
    * Called to evaluate if there is a snoop datatransfer for READUNIQUE from clean state
    */
  extern function void evaluate_datatransfer_for_readunique_snoop(svt_axi_snoop_transaction snoop_xact);

  /** Samples the trans_ace_concurrent_overlapping_arsnoop_acsnoop covergroups */
  extern virtual function void trans_ace_concurrent_overlapping_arsnoop_acsnoop_cov_sample();
 
  /** Samples the trans_ace_concurrent_overlapping_arsnoop_acsnoop_one_ace_acelite covergroups */
  extern virtual function void trans_ace_concurrent_overlapping_arsnoop_acsnoop_one_ace_acelite_cov_sample();

  /** Samples the trans_ace_concurrent_overlapping_awsnoop_acsnoop covergroups */
  extern virtual function void trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_cov_sample();
 
  /** Samples the trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite covergroups */
  extern virtual function void trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_cov_sample();

  /** Samples the trans_ace_concurrent_non_overlapping_awsnoop_acsnoop covergroups */
  extern virtual function void trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_cov_sample();

  /** Samples the trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite covergroups */
  extern virtual function void trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_cov_sample();

  /** Samples the trans_cross_master_to_slave_path_access covergroups */
  extern virtual function void sample_master_slave_cross();

 
 /** @endcond */
`endif // SVT_AXI_EXCLUDE_AXI_PORT_COVERAGE

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new svt_axi_port_monitor_def_cov_data_callback instance.
   *
   * @param cfg A refernce to the AXI Port Configuration instance.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new(svt_axi_port_configuration cfg, string name = "svt_axi_port_monitor_def_cov_data_callback");
`elsif SVT_OVM_TECHNOLOGY
  extern function new(svt_axi_port_configuration cfg, string name = "svt_axi_port_monitor_def_cov_data_callback");
`else
  extern function new(svt_axi_port_configuration cfg);
`endif

endclass

`protected
+21eI88YH,R;X#3ZYceVVY@Yg&R)HUg;Wd)1X(@@C>OYS=NY#@WV5)3:fX.6eE^O
cT-b3JP?XMXC9;0IR^\7=Z-NK7=F_C3&3]S&_;LN0cO^#8=I71a9O3&dg+2N6Cf[
B/E1@e1F@7E^&:GW-VSE78+F(CNU,P_0;cH4S[RRU=4d-W.PJ-8NE?4fRB-,#PUG
;@#f532NX5f5OJM6;@4IZ6+/cY,C[=-^\M,C?O\//dJRTB@U7b\:aO+\\fSSL4=M
CO:,0<C[CUH8ge\V?LPYG4@+[CdD68bAg9KfSW:2H?Y0B#U7a[4=8_MY^;Y,]\48
AC/#AZ5CTf]F+b&VJa;&P9e.B_,_Z;N.\_\Q5(&=+dT(d=)M/Zc?g.DOK-GaB2g5
M67AY>D\@HeXRY;:fD07MUKc0VE^RA[U:WabJ4\)_d82@Wb1b?M,SM\WYZOKc_-R
EATW]DFMAX1E(@V:3MbTDSaKW[K;ACS+T^>8AgN?H,2Bc73fY,6\<EeQZeUE>YW6
5-8YU09bXc4+:>TaAD2&+2)Xa/R5C_c/P2?YM8WAb0a4^d(4,E56.Y=LZ9207/FB
<0Z_L^;P;0G4)GL_ENI0UQ>_PPC-D5Qd(_e[P\VW+b=;(G]QfVE_V45]&Ve5-;XB
ed0?-E50H/UE]TZ/DEgHQM&U2-F.1,6&R)ga]6L=@.?<YUAZWVbA3gT)-^_B1\ac
4_2/Q:\PBC#VaID\4WG4H&3NPfHHGU@WCJV=2&dgG#BXPWN1]POS,gRJT02X\V3H
0)50(0(X3FNPT7g^Eg+P@NcJ#OJTPQ>fP3>@bd2JcCUE<:1QD4,(SD\[W1A_Z1La
bTQ,_R5DMNe@4N#S+8g.[.AZY8,3(L3HHR:>.a8&GB(UaIX0MSJ]^Hb)Ff/T0ST]
aGZ#CW8OgH6&U9LbeM^4/1+?S\gX\(M-Z\3;+VA[>be5GR9MZA0JOSL523:R)1_T
IfcK_bU9MB0(053L/D3BQ?)ZB\E<U<K@dX@I@\+>#eLQ@&3ARdOdO1-OCJSG\MO]
KS;9#P27W0BT-47.Z\2S6bdbTGWIMf\,Y<GK=TSY-KWW2CbUBd/fL85&,DF^/eI6
><O\(R\16H+=A7d-P;GUPO;FY:90e<WXODI58:NL6^S)3NT2Q?e<BR3c+a?GF157
ZDUM2X9M_e/gg1S]-F#62_Ve;.0?FZW,M:)0LGLJD&D4RRBd(a:5dK_IeaMP\a@?
Z6:I+BfJYS2_L0.bB>+:/7cIR(0b]QfR?4fF64PL5V]+9<Z=F:<KV(ZB(;a0U,2M
)eY<Y8T9XcH-.BB/Y\8:L3.O7H@81GT<LRG34\@WQ0M:^5>.=CIU/JRQ1RL9UU/A
b&EZ5b+4_&RXfcV5F^@2bLf=56<P&/Z#@=P6&Yd15Q2<8BBeK,:^Fd\44BRJ+2^C
bOG&I;@d;QQD?[D@XCeC?<]=_4a=IDLg_6eMbE>c)]1@6^/]9D3Seb@;I7R\<4=/
^S#TbH@g_N)cGd+]N\YfWV9J@V(T;:(NK;07=LNSFI./KGI/A,e)YU8\EN(d2UKX
]@NC_8146GO->9T/PeGSF])f-:Rb3YU,?F]+K/>8][F4WJ)Jf>bF(KGR..Zd/cS[
0C]b;L:4GRU]OUL0H^cK8Y32bbeC,^cSSAG-KN0eI\eZPC-AWT_3V;.+g\ET?JaU
5L6DPSN]YU)@[WXIQ,-_4/aGVc0;:W.b],=?#;W4]=67H+5EG^cMXdeM.Pe:bWDI
Q4_NM.A9MDRQWDTV37[R_F&L0\&IRMU?1[5eC-GV0KXQO6N>YX\Z<Gg&4?>F5VX=
8@Kb9@aN;\\bR&9#D[Cd.<b.<^01(675&E&+N6IPR1H,#^5RCcMcX-FV7I_0_2T4
+LZE8GSb/<dX?JeN:KY_UfT8K@4abd=1>fE#MEENTa7S?_AFZ?F_4MPLfP#&0@&^
.^gfdQ++/^DG6)JFN3I9?d^8FW^d+,6=KA1c[5@IDE\2LLM<^C96CB&4)&ebGR(/
b:J;V:91EU:Q&e9df9(^5IfCL.a\d2W?=E/1(Wf2J/PX=L6;#/DX4JA/7GJ/OKLL
adE\(:TaGMB=#+a>M,P:25[OfbaW7KdbNLf-Ca[HeA3QI>Ec+N;/(dT?5C297<?;
QN1B[N6::LL6G@)DDTf]fHDD(PUB:P:]023C;DMCU=]_29M_?,C?.0L-)PQ9PW2f
ZU[RTd9Sa7)/XP7f7B=A,-YdBVV<-.JALMTISGLM7ZGV6?W#NSb,@N43\0F][Y_L
TaEPX90P+DY?5Xf\IIaUeGfeAbg2B?)F^>NN-=NY_MaTOd\;?eK)9#4c56HGIRUc
9WgX/B5TA&(;NJ(X+-6fWBT<HcELRfde:BQ#OP=V\M>(-93CZPc9^A5WE(X#3.XS
FZZ0J/16K2>958F6Gd.QGEO/,6:-Sb>]?e^e&d=S9eAZ]0DQXMO(^P?>bFP?TNCB
C/)QPL/\]LJYTCUA]1A/I2H]/0[.#I=R>IO^TIa(Z,KTe.5ac?ABWO[fb4I[&3#B
SF=+]VEcN3EGKF-JQ_>7LTSM@VCK>#TNKGG;NZCLO]JScYK;.S08N<XR_95T\T6b
O>-1F@#V15G,:W<6:a(Hc(-1JE+M_a-gBZb;UYHOWK0_eZKY47=DHf+1M:P::FgK
,\#]BFaM[#dY#D#;?&d:7>PgVJZWNWSW+ffc8PT=F16]ZX/@SE7X+]SQM]?Gb;SN
V\5N:_,JDVGID.WYacN)G0d\_:Y8]NHaX2-/M+/,7KFQ5fd/_aR,17Z^&QfF-))O
P@NS6(#DF7gN8a(P9YL]:<=N,[FVFe)\SBbM57bIJcYTUK@,GF_F^9;KSY4XUD7S
VNgP;)DPSJDF)e<=W.[^F@;T;J):dOBcPY&:EU+6I?.YSc\R..T41]@d0HH&#.)G
<)d?gPPHZK\>eYV/H0QR.,6gO0;>GUYN4TP+4a2[QF+>cG?Xd..]J(Q>S=O8_g:W
;VC/N(@-,?]LWHLW1E>O3HR7COLJ6cA^[?XG_&&Ua#Xb@4_M2&<)g],6La>AY27b
WG_QXb\GFX(#YBG3R^[AH#,J[@^bCR4:J<Odfddd5GL)K.GV@L:7M:ZQRD#A6-XE
TWVZ7U_6/J?HUG2GV(2+Z;T<dTe<g8R:EZ:EJQ2UP9;#(+&F5(T/bI6T#4Q6c/df
D.L,R\Q;RW>#Z+Nc/B00VV=XVb7&A/>(,D3P)549^4S-ZU+_BEBI8;=g<X)]A5?;
A<O[&=:>/MHggEQ]RDTM@c3b#H^NV7g;CVdEEaY&fM(MZ#V:;S0V^N;_I)FR1+/B
LSQ5JZ844Y0V[a[(><;f<+Wg98a/:EHOgAX;[F.J7SAQB&R,LR@9[UZW2=TNH?CV
JH7;Jg).Y#fac-c.P:(.9O].U4a9FPA9.&>VNHTf:S?f>ZVO:@@A>db^_dT=(/CV
5),YD0#R(HVKA.+=PHf+8MOS;8fdfJT1G:=d3f),U.CKN1-e<BXT?A-;:g#f)0(W
#OVfg;E93<8a3gXH&YF)79;CG3DLE2c^e2:#_1Z#?N&XAWS65UK2gD3B37gNWQA&
BIa>+WP[eN^C8T]2KEK&SHC\7W)L@F#,K1D[&S<?,A4,F63cZT1)#R_Y#g(&eP+L
9N]fU(fQVgCP\^K@.7cc4,4X-F/dE@P7gQHW&.DBX8?d0&cN62>,g2,.6IP]-=De
HP9b<cc2Ff6a.D>1-B_[,/AI;+7R,P;[69.8g54=_>C6a(EL2<,@,X-b>b;BC,\T
COG+-@&_[fF-G?_>&FgN?(X]e\+6L<cF+3LOH&TYG.4=HH7aS.H+F1A\CZDBYZe[
1Z1@2e?SOaF<[S;gWQ[T6JF5:8\PeR]K>Y4-<_5?9&=A56C_Hd-D/dOC1=0PQH27
Y;Q;VTWC:XXQ;.,/Ec^_;YEOU_P::,&&L2D]^0#NM](A>b++HKT,<F#c@g,;+2QB
5VZ>;G,,;0D6eEOBC2AK4Fd\2D_g6E,^c-)bT-4.Y_M8B<<.cLIZ:57SM8DV5HZ4
]>?Je)CaUOOO=U8>I1NdVbJb;5b@VO:;JgME2E(&C?&GG&#[MbJL1<PNG)Z2ZO;F
fd&:FgUM5)T+RHU]@=<f2EgP^CW;9Y5H3Ya_&]@R#d+b.HS3M4S+ETJW2LcIDgPM
DD[&9I34#B59F4<+-:AQa)2,d]Q1:,-@5-V&U63QHY:7@CR60dESf+R;R<FX]>A\
J)T8<b(K>ZNGfPH)OE:\1O,EXM];g=^(]W?;6]?fE#=X;R54640IR(?98T88J3:9
XVg@V\7G2Xc0f35L=;?E58;97bKYB8bN1>?A^&2U.L9Q&Hb.E=a,aTB:]@[AU]Q6
+FdVaf-Ac7LU^IPg;97dK3W&&0+J42@3,Yd]=AT&WLM@?[T]ae>>6aI83XMT=UF(
6Z)b)IW7W7YE^eKXF3]bWHZTad,Y)5ERaJX[LBA=_=/a+I+.KO<??D\+<YRc>7YE
I8;^W5Yb+MSH963g_N3.(8NHXSLaTTQWC)fO//I\61G=g^G&QKbYb0BV4QSFIGN_
+,Z&TVK(15QRQ]?\YAS,WJ8=dVPG;P5<OAH/,>_J58[X()V41(01EI0_Zd]5aPQA
8SRJE_X=J2XQAT?Y[6?PEKY?<Z5Q>UI^88eLWF[\]R:<a-RES>J1daL6-8.PYBBA
B.:_T[M/W^J[>cRJ<;c<>Q:\BP1aHPSb?/#E70YX&\LLg/(^ATeDK>[>/OJT]4/[
B9XSMd96W9BPIL)^24QXQX\fPYI5Fa^<(]/[A(8<C5]73XME&3:-dJG#dB[M.<VG
6O5S]Vb.\CPU<ef/LPX(SLb\+b0((T3_b/:FW@JDUN3Qf0VH]=+F(85AF0MIF[M@
MAN12F8De>]^<9CDZABMRNL?<Pd&.15Q^([L3._C?.X34.]U\CCRZa8YU)1a6KQ\
])L=A\=4/(f#NTa+,9J8B9_X(0cDPC]#Y5I]<TPDLRS@;_4e[E-E26cfKQ+2T,OV
X(E\Y6YGb[UI?X0H<XYa6VPJ.X0UQRCM@#)U74C5DKUe:ggTfg5aCSX\CSf\,3A2
XS^N],\WV+_W5OAVYX_FV,&gY5MV,+<c=1]O:H)cT,aFU66(@I?_H;#Qb>48\=f:
J^(&2WU>/B(UW5ZWeVIB5EP?.3D+_Y[Tb^0>1aE.M>C9:A((c^UBB.0J?6/g>d4d
TK93/A?Qe_edgNA1a@9;0\(MM)\SNRYePMK[X+V@HZ\dAB99E=fT2Eb>P4#=VR2Q
]4890>Z0,SYQ2?S4a/[D@8-P+:RV(HQ6+#_LN9?7]8E:/J5AO-45a\Jd7KLO,=W0
#9^W6>^A-W,#7SP@LG#RN,[gKZ-DZ0VS9J#(a.@FJf_NR^6V\a)MKEO)=,@#AO;R
GVD7B+LMQE&HC5aD)SIYT01#BD>:WE8]]eC26[Q&8-HRGU)1(K8.JW;P\IGRee?U
Wf:b//=g&X-9PIF9:.DKS<J\20&3e>XD<CUI,@+)Y_#<9YYO#>VG2/JSQ+a/W(Je
FJJW8.+I0G&U(SVV(I@HDA:cPI^TYF35X7L-9\T1-)]LeeNH.g7JQQB_7T<W)gSV
?.DM3SBH0g-5):(9e_@\#U96=3H8T[M(2I&0R/@VQ_IANK,CTV_;MY\:Jc>3A#0;
-=G6AUJ;V(:Yg&DD>,&ZQJfA.NYXaK&>KfTU.ED-#dE#Nf^X8cRJBW8Sa_Xd,J>1
-,dNgCQEBZ2f)ed(^I1PMF@V4W>+CTSK.5&?4?gUCYe>=)O[M/>?R35,,X^&TAIb
<(-S(eN=F?+>.M8DAVa)PGEd6W+@+LC#G+796AT<:(XeR(6,c\,&6cNF.gb4N2:B
,[FI37]e],_WK3MQJ.-@KBcMbVSGD3/e6I=a>QR=[4bNW]ZcDc>/B)MMZ:&.]S@7
L+T[f)MTIKW5H:^_fD7,,Md86a\_]7?J/g:C,gQ:HVHaUaVf._;&-C:UF:V+Y:?]
D/TNe/M.?_W]1GJR7f>8CZ.d@;:0[9G)&Z.-;G1A3g<]&0Z[#_1:#NWOd4M>>7E1
I)^;HUQ8/]W-5Cdaa9fbH#0NGC5_R_,ND),T7^#+#XM\Ha@N_7<X/SQa<T<2CCab
))D9)>fN8XS>X=gSXKA<<L#YQ\9?&?EY,=JbcA>EN2>dQH2c:8Y=:[5YZ?Db1/CY
UR8CL#S#)SUZVfe\DfC_CfU#Z7?175-9_G;==(X;cNacG-E)XW]-^@4D->\<X77f
IU9>#M?N^Y7[4R8\?3&4#]aW?Y3\Ca.,Udb,U\8^V_;]Q&AQW5X2]97+FH5IeB9&
FM=(5&QEe+-8C(K62eV.J\b;OVRD.3&_M&?CKF@JeX9C0QaNF(CSLEA3;3Q?C?9R
f.CbOBb?,/C_a-8##-PLQ_aY&7K&e&a^+:;GKGMROc^WCADI-9\H=K?[^c/,.NYF
64fgZE];52\V]N58-BN:3ZA)__,)c7[JARX_g#Sg./+14_g4[POE=0LV-,R1M2)Y
0=N(3#@.T70MXC93Y]8[bK9B>ZWHa6ccC#-]Gb?H-4+0AXIV5-c[Y4I)g?KTVIAg
EC^Z:a>c1QIY@NM;B+,KDH&^G\)d14.[_VYgM2bS=5UI,eZb1<_8T-]:4)LaJ^#O
K3,Y(#\cX[Q)GFECgH\<e82.c(8G8Nd5V37L1EAOa7O[RB.@YV>PaF?MfO#c;&(4
CH_+GO/.:6;E^+W36PN?#GO-J0-/<+/\JXDS(c^XHW[1A29;Y;NAF=g8B9.SGV:W
fJ0c^&[@9XZYG+a/,C4SM-3Y8P,=&0@72.Fef.59IcSJ;RE,S;I/1Se)1Ob:HWW^
_c+P)U=/3LIPZ(<^O,fa3?OLH1VQ-1KN;9Q_]:dJAEN+g,#g#U#5^X]NKKfBYZaG
8[J,:V51[IR=.ZH>[ONA,F>TH,:&2Q-;W6eKGB)DQ3_P<S.YC@ORVIC2IE.;;LAR
-[;e35c]d.VQM,P/UI4J&bF=8?VB]#Y1(.&,65c?c@P^\?Yd4SQZ^33X>DGeFFD:
OOYgBf\.aT:/39MD>@URB-2,_+@:8WJU39d5[-MDG-YCfBJ(IO]eD50R9#ESLeO.
]O+T3E,<K6F=fOe]5(A,9QF1d0UgcY)Cb-HI;CVH>3.(G+24)51H\M:Fa-&GMM&4
0eHJ]S^OT20c+aG)\d\NO>S0)X[S/;N&<[Nb/O=XBTCg@Bb(\,;V>M;HRD8V2>[V
QG7C]V25TMTaADb#eL_4ZDa\MTaU1MZ)A<[^:5QDL4+Xg[U4B,ZdGO3d4c\-<Z(6
07[&SQ>Bc_S=#==/83/Qf/7H+FAQ1Ng@EgK:IZ8XGg4(VD0,N2b2f\Gbc5Y+(XGF
,AT9c?0CK8A+)eEKCa&)D^?gI-]MCX91-A/HS8NK=9/R45X\V,)TT8(X,Q&B?(8&
IA3IZ:3;NBV-/O6\[g8f@8Z9fD&>OO#:<L-).H(PWK&aRaG;J[;#FcN9PGUdWA&D
^5LGZ)5MS<-F[VF_fGFV5e8&&4<:;LCC):bFIFT<4&)0WVbR_=X=]ScX#\:GKDJT
.bAJ0U=&P<=ZML?aED._c7c2>4#bI_X[&O1@7H09906\QZ@HJOV89C\U+aGY2P+.
\)4bH92(5RCZ\da2HReLS7P0aA>4A)MAdVK^6GKI#W<I]gC6g+]a:=B)?M-#:GfZ
TCUg^d[IUDN+81H-:;eHBJIMT_;A\Q?:5bN+,K1O<2-DXC/0ef9<^gbQPC+4D&Cg
P^[:5c2:T>B\(LfF>P4L&P]c=]/#=\EBKAW#WC/N_UF9-a<EFI5>g#g/\L>I\OO7
[[:e@1FT&)?#EO.UAde)fKQG.:A]<+GEg#LeQHd(;_C#Ea_bWQ^+NgLD&Nc\8W?:
Q.4cI47Y<eHK>&H5&=U-J&^c1@7Z6@S\2@G2\cb(M#Ydf=XcIW_17fZ>b^(H#VPM
9ZX7TD2_;J;D3P5G95Y\]K]1b(V#.;31+Y]U35H8KEf=0^9aR8J?O5TX-]<aP>G4
>\K^ODb62>@XI//TVD^@U=(P4)9QD7+L05XTbFgV0W&H#Ed5NX(5d<@0H5D.<b1#
U36^<I5YKM3[(\MeRQ=XQUd[O-\V,K11_JO@R,Z73=N31@dHMAUI]@Dd(4W<\+/C
D=cC6gc[I?QZRTc[S^PTTM?=TZE52@LXEZ\6bgU+VLHR\.EDCZa7Ac5c@ZLSZ?7b
X]A3(5=TgPJ(.A<D4L4-5X:I0)Y]6-0]#gWW@aV8]#7ZRbNNcGDCf+:NOgV<L/3=
V,V7RO^T?3>8baZUYJecK8c=ZF[P]EOE:#)AeC+fO9aT#aM<+ae,RCda^KFOO&g[
+9ZMG7A;_J.=QKO4N\.dL#FPPAA[\b;CH.G.J?]Kb0a,0@^KUFWcO1X/W-bg#@#8
_JLSKae?.Y(>^)9Hd\eQW8(SY1^#?f,C+USX@,;Y6NYU>IL?YEIACSY0R^fY3XTS
4W)0JD81J5#QIaV7g02W+c@VX44]A@Ge(G0Y=M]\=-7#XW)96&U?OLg#J(eD@@2E
<-9T/66MH.Uge^KIcbA;=aC@EUC31E9X#;b@;)@7H3\O2WMQ:[K,^?_8&9JT.ZP:
:TX_0O0DbSRF#H/6CQ/ZAYOG@,5H\GL2ZYCO3&1d1Z;#?2dd)2aU,fMg.=</V]5+
]6IS=GX@TZDU5&_:^g</H7P-DDJVT5MSGbE-#MSO0LW;R5N>Y.+KbWX?QJRT\1.H
I&_RIBJJ,4QB(BJgO[RGb/9_Q3U:.-3.]FEI<8NL3Z[);cYQ2W[-EbeYJA+8MMbY
8G0H7c[@@/,J;eNB)JESd0#<[UYe4PZV[@:H>Y/1X)ME#9,<V6C9Z#=Y+\NXa2SU
MT5&:>+J=.NPC.&#OXCQF4e_0]4+E@@fJ@H0^Q0U?94c36ZTPN+>VFVYQV\WL?2d
F(f:.EV^Ncg4-H#JKBHg>D+Wd2ebQL\Y/]SW^Q[C?>BHU3R2W/9Q\Q\g.I_V(Jd>
9:G0_9@dMFTBKaW6H,0Z@O[?a8<#<aRW/39Y?,K3+X2DE2RH@&OR6&XHW]EJJ-/R
Zg:\++g1L-.=C;#g0f+NLFd>&\<+gB/72UJIQ)agJNERf#)A#Y?NKHU\))+=;aF[
#]#,]:G9eU2[):CYJ4c;./^<EE&67K#BRK6.K09]3<X^/L)+Vd?OV#Z_VA-?:gD?
e@6(.IT^U<__?-YGaVGBM+LZ#3@,1P])eH/\H._afXFZY\g+S6U(1XV0Q/fKFN65
\M)LT6:[IFI616I+K#H5G@_ee;L9/4b=bg63M3Sf);)&(8)B<^[@TFOKTZ[Oe:aV
QB-STO:B?LCbHZdC[/TXT&dF0ZF?[g;W@cDO@^XY](ZRVO#OPL;P+b+HXC9.\7#\
H=FNOb^,Z>\C<DUNVAg@#S;;P#?I-/B93GN_0A,V7S]EW)KAZJX8]B:fYJ])&be&
7<G8/9/H_fcIIaNAO:DIWPdVR9/X._T]_g0LYIdMeR_b0LR@ZP7OG)A1PV3f[??B
AR@:_f_[g\9dFMC:M>7]+4/ZX?(P)J_GFR3@G9Fg<7))OdYE/>eAB&JK\6J_8a,d
F3;:5FOUJLW]<eE(6G9,U<[eZS12;Gg,4I,=VT(]VG_=9OJ9)+4X?CK_Z&1L:[9B
\Sb_T1\7Vgbg/)U087=7CKd/[0(dRg;N-OF-1;37bXKW-2Pg;10#GAF/M-/FfN9^
NSQ?..?09JYH,5M[cEJ.d@6AU8Y/K^T=SLdJN1bH&2&\.XG:I,VY8P_JSF1M5f:M
DF\?^0@OOL?CdZ?2HW8UgTA._QDP+dXII4^/&eH-QPE8]GcJUX>,B(\;SbbWMQ\1
B<=GgY^Q@g)f]R03cQ4]0#4YMX5d1B0gK_;@\,]K(b2,:C[YL\YCZ,CQ5T&7C;OT
60G9GUcgL9bHb7<dfHOZ\/5fNF+eFKQc1,[C@LRX@WK+(Q+6(W+X/.G5f9;-_D8;
YKMGG^Y.4VPJR5;,S^b#>^F3WC]IS&eRC)5\5c)#?JT^MPGFM<\^bU;^SKB<DaP6
I/gOI,3Bd&cFNO?;V2AFJ-4?Ge-gA/O<e,9Hfe\V&eR+YX,3+P&[<?U0cAPc^]H=
>DeA=(5:(b8:&5?6S7cZZRa)=K_f(>U]VE<-@D/&aSHR3g#?@_VaKUN/5g0O9_[J
Yd45bA=69I3e8+1P;Y(OeBSbV?3E&)I/Db6,UV4CK)RP_6AgAH)(&(DYDG8M1]A+
)M8,\XbKd=/O_\145<B0D-678V?:7AMbZDSL=g:8#R?A@dL#fO-@=6d:8QM&Q(WY
^K-N6PALWBD;/K8M=?6ed>W4UbIVS?OYJg=:L\.fd;)BH]\W;C4b\^W=7E>g,H&S
MKH^<@BRdMJJX7d)@e._g.M44^.(LM53>D=[Y,a5HJV#5>DJ30cW:M8C#?VRAOQ?
+fa6bQdU^:=bXD09JPRBG_.a;9H#CU?XLXDE_f:02N;2EcMXJ43OPUe@]]=V)PVD
_4BN+4dA\>P?A89P4:8574Z2X84@IBH]N73U]?OB+FZU8G;BC71MYC9W8bPgU:1#
_/&7]dHWNM6aD^QY=[TCJN-4?RI8KHI?#d,7eZ2c+QI#Z>c?HULD#W\W_=&3G([N
\S=(HKAXV^]<_#A@Z[4W,adg\^7S2]6aI]Cc.eY\aZ,H,^O=X^EDC@0cNUW>Z[6=
Y60T9+dB/>:)&VOa/48)Ga6<G.T?(a3X/HJ9\.YG<[NT^?Sc]);H9>Y>(]7Q^^a0
S64_II9Taf^A5(UX)QZa#@ga2;GQ^6FP^W+#U2:FIO)KK),[55XM?5Y?.)_-MW-:
VN94Y7ODGT[4CZ>V@0V^(_L9_V^_bN]_Y<HC(?Y.PaR)&NYCYGVA5=CD.._UVV;V
Z7EF[H:O//F#<Zd2aT_c>2NeXc<ZW33/;+3_L69eb:X(/:D;a<75D+BPeefP]W(9
V/Fa<QXS1-94gEK^OHQ0RMG\,QP5XEXYg\aMTg+O9BZ-J=e@H,R@-K&JLVbC;0Y#
PMSCLZUL+8K]7OGLB\NZgWTYX==\>HS<eEQ2[8LMQWd0(9HMD^b:7?&=/#a))1K=
:2f_QGcEbCZC));FC6V2:20_EL<@WX5)GbI]-TKVH.1G1_HTZ>XX@Ee3?Fb)S?<V
_E2I3D0U4L-U6fS-2Ef@.Oc=-=9ga3C5NA-C2RM2ME>RbL):0EKFNI,g+#J^#3c(
P;^C7d+(.GR=TH4\PAE&&S;bIKQ:]9WN+/([O_9X6GR8,E@V;E0a;^CE]3)aW[SM
J00D=-R4\#b2[E4N08>&3P_OX3.,(SL9fRb2]M9))\e90Ag#2abcT<HVf_:;e=a<
\SEeO?>?2X_=4<+22KL(3gLG:EIW0GGD7I&8()M2[aB=L/9\fcWg\bY;8+6a]2KX
P?).R2K01b4VJ(?5JMS(-5ET-N4.NIX)A(U[QXWbJ1TFf[ZPBSX+D\W>O4+A>)=B
-(JZIFNa2a&)ICB5_7Q#e#d8>L3>[SBI4@cMfFRJ^<)51J?]RKb[:HV0.DA&EN<M
?R.Z/[DNY8aMG>PMSKgB2UAU^-.\RJ2Fe,31W1-NS3d\JT(]R/3SEP7HWVO^:P>9
T7GbG3b9QGCSSGOY6</<2P_6FT5;:4EIG?RZ)gNg1RI?fRMPD+;,YWKJ3=13@DN,
54MEBR0cRMYT/(V\I=a61P)I6YLEL^\5[:)+3;+9P4(W(<+<2XLXG@1Q)QS<TTb6
993RM4d;NbO>3FW/VX04F^_#cVX6;afCZ:=,#cEa;X>TE0-BJN7R03I@LN7:OGZ0
;+bT0]9D.0(MK/46S9GP7g\NSTQO^C87U8.@cNXcQ?N2PR[g&+6S@d[SH_DSVaZg
)W-SGM;6-0/>_,JTO^d_+]cfQK7XEF.]M2+bC_5U&9+EBD:W8JQIe&dLLXLge[E7
2Q-^+Ee1,8I@BY358BLa7BYdY/W?<48IceXfW06aaR\5+1TACHJQ6R]?/TS#c,P5
4_+ABRY48??JK;7.6=&>\WE6R1Q.bXG9I)(:fPE@YDJCg[VTI+,Wf/Ed0U5J#0@;
#^KF6F?3?14g0+?XcOHT2gP7_C;DVS=92gX7O^BCP)AR<A)3@29/cVCC[H=VZ<6?
AH:C(XcGLOCNY-A/FLb.T];@<CLd\-bVC((D,I97gf<4\GO+&^:fO.+SdRN,@W^K
>1L;P6#M[JOX8A/_QR-^L,\4\&\a:7f(H>-0R/3(-ZXF)35PU#f^dKY+3:bYaFNd
.IYV2H&4Zc:MKNg^ZF<dZ#.?:\JR(.5f&+Pa3E4&-H032@eGa_^b;RF4?]G\eA@,
PDY]Hb08c,ZCH<BKDYAZ^=5A?LQ#_+2VZ;246?JYg+GcCSKd-I@ED,I[Dc,74)W0
TbRRHCeVc&FHc1JA:QF8M4[A9LgAS9C/^P5F].MY+?aH5RY^J7+d-1>ASC6(&E,_
a;-^3c8-[1HX<XcZ;\RJZ=8T1?Te:=H91W3_:090KN(M.]7F1:OD#G[YYWJ1/1e@
9---cN#3>,?3_<W+fO8fS16\??b..Z7,_0\3]Ngf3c,R8^PaTQV+f>b,2#g>4>PK
Re0O7GZJ1,Rfe8Se[fRTe]fN8\g)bQHHOV(SYYL@TE,aHN]\)36#.9UP:)X#df^F
@:E<]3#7,7)-XOeWN7M@OBfBU^1F1\/^SV:Tc4Z+O-3DPbM_\6cT79?bG_52\FP[
dK=YcR]@cd8@_GI-aW+TVbba\#,4N[82&.^,-_-b<HYCNT8<B>]2a../]1d8fgN]
=+gKBW8gK,O+MB5=d)#972DLLScfPKX[_2:>]]f\1DU(6N(0QGFa>84?N.]5PVSM
-=ba9]gI&>@13NQ69]M]=,8E_W@Kg,;/aOd=UJP.TX]WKOT3TZ1&BL:O<U0P_3L;
6HRIET-6_P]g:E_#(]Wc<YgeJY7VWY#<87A,L4+@P<3328UVR@5)KTfFR&H:DK3]
:,AC_<HE@ASIdB@)P45?V4/L^SUP76EDM;F<8>3V@/fO]W@F\.-C?R+6JNA-a;RB
)7<^/T@L7B\FEQ3g<g_K&gZ:^K.+G-#L63L^.UZURg_DZEE-/9WSM#^,Ve^2d7+,
NaB1YWB0dg\3(0],GWED.N8_5S#?KY/0R6J(-&7E[7X=eV^#LO&QDI.D>+1Qaf_5
\^DQY;g=&GLR&5R)eZA&RYgdMW[MEUK8AAHNU#E4?WCS\Wg[8M4Z?Da&2PA4aBdD
]g]QX:=QaP?LTDP<.^-eLc/[&BNc;e5#&,2a&D#H@A/(bRQL07La9P=(UZ4V;&?V
>.ZNN##_)-)D:aJ)HCd;d9-Re0DJO=DR#^?NNU+g0DL+PO7[BOAOR_6;RGTXM<=6
+b\[/N^F;E_2F2D=?UPQO;J(#&6VDRX<[@9E]c>-?:.WSE(-[X@&E]QbMM\L_Q[-
U)=FT6dId8V#M&9N9,R>D16adZ(-I<7N^=1/fZ=B;g514^g-FH&]FI=G7/<-:?>>
KgXYb7Y3[N10B?/PBXMA\?V7c_].dK3a^0.4Q5ffQcBCL)gOcbD2@U8D6,0^E/:#
:U4?<ag5a<P0X[M))\?8?1@^[GI1XG7[RWR>A2bIRB2(UIU_7RJ:VF,aN#fF_?69
VI(+&IW>GWU</@Wd=\5Ua-[]1?C(@94<&UGC(6]RV;4@L<;_fGEcQ@QLWP)]IXH+
[Z9-O@ZaL.1GSU;Jd^=/SE:7Qg>8/.SF&-B+Y+JVc14DXFXaMK&#4TM1\8>dgDZD
Y]-G?5RLT/@9H:<SL9WH_1=QU>e25HEX2-.UX,fb:d(g2dIV1Ug7FFE=42MPY:fg
TR6&QGK8cX#UKK(ZVF3H>.RGAB?8I8;W0ZE.V9KSYbWHB=06Z5_V7(<..(;eV1OU
IKZDAERGF;ge]>+aUf_fL/AZ:N1DQR[&20PZR0,dVIZ=UL+3V._A@b\?,BN_\QbO
QAIa\(c3&^TF,I9G#11fgW2KX47cQ:M<K:W7NcTSF))6(LP@5W7<OB_&,4_=KC5B
(E?;a&^KZ2WVTGb#&QE#(JM1dMGIYN1+\C<GWF.HB;/#TSTeb6d8HQ2@A13S#:@K
?1,P]\<#2<LA/K]EMJI98)?cU<4<,\Zd<d[fWJ.:^I]U4A,U.]]/ZTJ(O;K.:;.>
WK/Gb.^YEG7N4J.10W(PVAUC40bE<&3?:,_cCDTeKSf1YW:W4PW@_c4V)DN;JWg;
8L&PD[1PF[G-49^^&X2FKgRH?Y-/-UdS>))ag.c[;EOV#DVD+(3KQcFJX+9EBa,a
eX>8=QMf]J0e)_NC>fYDX5U1^8JQbH[R#+fadHRE?36e#XG>Ub4]ZZH9<]U-@F;B
7:.G#.4dJ_XPV4Z6#g?WAPB.,+C/>AL-aOaH^LQc&5HVJ=4DLZaG4P.4RJ)^@SKE
-V;;TX#HAEG8?]/SeR4>dYeFUT;aY@gb@&4W^/)]_?GEQW8UT:+EA8_\J8IU/#da
6QS]&^6IPF=FZFfUA8eD_C^:@eL<I[PA&[/Z3gQ3^Q^K(I,f-131+5ZR,a2689ZP
R&^@]6KV>d1/e49N\&X,fYD9ef?f8@+CR2T<<)d53<L1/EH1VK,GB9>bCcdVJ?T+
ZFfZFP2YQ/HaBIX)G:NJ7=W47ZN]+:XJ,d3@e=E?GS^?5D:RJWTQP0U+5?-3BOd)
[f=Pd>G_@BI4WW=&H]c2I&T2/ZR7#K3R:f@^:M5QVE2,_O[FG0add/de+,0?)10f
]0C+[GNB31dD\Z+J@(M7Hb++7G&K43>]08T3]]W0N/APSI)PGNcV;4B3&H.07+Fa
W:^YebJ<\4MMWbc3e@WEB7,08Z\G4_.aOKM_W=94W#@-^bQNV4I&?DDHB)7Y4@UN
NQA3TcZHG#^0#d<60Cc7.X6(]aGTOd8@d3M:fZ>JOb:c-7^eGa:_QXL+Y@Z_7LUJ
SCN+(^V?VT:2+ZDWbU?Z+5>AJ,B=e3+F.V]?9#FLNJN;dX]:BEO]]92[&gB1&/O7
>#F\KMe3C?;R/D_-SIA:8,3-4,[-_4c;,0YT&9?N?gXX;+0cN2[?3:.+&::e06@;
Hf;Z>I##&T3RUS2HGM&Z#@J,aF?M7.DSQ(B&X>NYAMJUXHYcS6:OX9f\BV1M)1dF
+#7S+R\6A0\O#BSF>@VTCX;8RO:,IfXXNCHC7b?R_UFVZEUE7)R.SF..?)2F(P93
QbfC=1,4RPC+I(7)-UfK37a[be9M1G8V3UMW#d#:[34Te>YY5&T6c4JNNW5bM[@d
H:NLUf[NCQ)VV+b6+?XVY=&^)2)I#G<-=SY-&K>=^:ga55X\E.-R64AEY6SDdA.N
-]8#-.(LTd0V=eL1O<.G:H+7HY9FBP:IUg15Q2ZgBYG.7:dW,\JRGc\E_eL^L/,:
LMU-(TELRDfCXCT<.d8234YWM.T4#?,2_^P+7A/Y:RVeERLb?O]Rb@>P82T@9>N<
_\fF=_ge\b6YU_:GQ/>FNcNb#YXG6-E;/gY4MAOTGH[,=5>[ISJa3g1Z(L+R3]+R
_./b7D2<TK8@Q<If=V8&EB(FZD(T_I5]DV^937W1H1+F-9MJ<@01#1?aBfO[L)CG
cdBC?dP3cA&-SKVB9b^UX](+DC)gSW44Vg_8V?]P_7+dF),VQBIbDK.H4/I[4L=N
Y>4[_093VXHJ[3KH[;M7EYP^[2GH>[cJdO.WQ8];H@EHgOL0[^11M=R-a5TW46,5
=a&#/4X6LL^CRZ?DJ9H5bg8R;N\42YSD&3X7BR#+_.E?<OSCD2:\[:^34^M;UV@K
Z&RM>d_ZZIA4KV,J@)gW\OEV0IZg=H@g<F>g,C>J1EWY9=H>#6SQXg0[,6A]_4Ce
;7deBAIS:B=IAcP(7[G)b-KbB,H-fX\9(5b,LW+/L5]0KKRO,ACSIaANg9J/;L22
4V(3SSJ]bU03Q&,8&VBXYWT2_L1V46NSe@<V=UK(T160ER?1c?;AP(;aN2Z]c8gM
?:Z-J7/.D5@.JP#4)X&-<#QN82<YJ.E43;\a?S,;KZY41K.eQ(QgO(4R;EZGMI_,
&PA>TDeg/MBO,+S&FaOG7SOg7XL>B51[T7a#IM0X.R1D2&,:>6@:?LI_QXMfLgd)
TFL==T>[+NK3<JMbc>((T2WX[XZg<FC@WQJ2#RI\8Z9L-+SGGc0dfY&C?+>0T([N
YGL>Yb3C.]>e</</eZB5.OI/WQ2I2fZ[IJ?7[VGa?DZ:O(c4NQ;.3(bG8?.CgOZ.
97P0cXIa.JL3&MJ5[dH--Z,+K(?X;Bg_03PMSGdZ+Y_JZ4N8TN>e2Fa>_^dBNS+E
#=6Ud_aGfH/.+;Y:-4LSG[TbB6TWg]_Ne1+JQ+I(#BONd30#d/)+\(-UcP+E6<(^
f@KBE6cK>ZB3L]-NQ56V9HAPYQ+KZ77(c??V;CHF.&/O<])FFebVUb#H4P1KM6Q9
gSCE-[RWPI;f@T^-QF803\_VN&N0d2eIH7H6^:_11E<d4+^N4],VXC8b8GLIOcJ:
)8ZP:g\8UbHHb)0;<S8SB0XHP:U8K1+N>YGE6=&]T\].TXBD,eM:4>5IL9DbF?F.
d9FZB8N56Cdg#0M4;>@RF+OQdIHEIT,L7F(_Sd=2a_CP,TXa2NKZbVaS-J;Jf]EX
+683.WO@YccC[:b3/GGK0JGTE/KX>,H8K-QN^3eD9J5=JD=6?YUC4[gc8)Le44LQ
+B3DB&H.T4;#<R;#@JK[LE;I#(KC63&-.3@fA#=2D?bTM,\]a;._URZ66V8b7N<f
51N_8,a,:LUB#L),&GNO\-7OY.K&[@JT9Z^R&5.+MXLT-.S:F-?S;W[@ZU,?;^=T
NDL^KZ6f24:6QZOK9e&:1=9RXMd,d4ffP<.KSGIHYL6W/<]PZ[4/AG-VG7PcP0.,
CMI1,7G(2f1Ff_eWR)ggQG[4P<dY,CYN3N#31Ze:.QD9I;\6:;3=cY)[bA1N,<KW
#I<d4PGC-F[9d&:IQ6DI^ePU4,TBFfce3_=UWIS(=MFQ]YY:BgaLS>YIQfT9I?I\
U,8SVBeA4T#Z=OBDQ<MeRe4#6Z],]fc-HMg>URbA5-9d5TRD@Z?ObdU_V\#(GdP1
\)ADbc@?N#?1GYHSH&F2cDR3BN(A=F@+-YBIOZE,LKVN#)SQNae57<?U+<\U>JE]
-ZGU)MN5FOT4g.@+2)6+C+HRSKT)[1TQ7UMYC0C.NAE_LNHJ3Q4C)G?DZJW+X4U<
WUg1:AM3Z[Wf@E4_ZNgVa.NfQ;4KCdf;,8=bGfK9<DNbDV]NQfW;].YY##UK-:JP
7=0.GMTJJC::SC>]PDb1CYf<gFMZ0a;ac&.g@?&P/(f>3eT\WH.._M,Z)dS3H@,1
I+fO?@f/+&<&^R9dAW:\:g_S/=d-)b1LX+S]/=B;c.,VP,;8#>RL5PY(;c]--_D2
]eTW+WaD7g:MZ8S=DV:cZ.4D:Q_YIYCX<)335b8F<+V,L;()A#6bNZ+58F=0PT_d
#.6YYOB]DdQ<T;C>URa+D&VAV>_N[dA<c9==LUCF(M.8Qf-RD<ENTL@DN?6)@/I^
TU_)\@I@c,7I;Q0CDc.eWbOKW@-Q.e83/f;?e89K5Mfb_SCBUUN6ZeI,WXK0/LW?
GUF^P@HH4fI>MK+TY8eaJ-P_cS/C-BJZ>KaDaN;-LJF0FEF[7KVE9^HO(_.[,d-=
I#AgL26g@aV^XXBM8[/Z/>b[&[(>dgcYZ]61S,OOBeFa:QMB^6ONH,eEb)\_dL\<
@f[=#B2G9S1g^N)W[IEfGdD2;76#;V;D[4e+V-8KGX#PgF(>fI<4TJ^1)J.:4bTK
W#2VI,4]fZ,9M)W#\9)I.P<[M:IQ1cS[\?FY;KN7+0LK\2:C:4X8g]VB[AF,1MEA
E?HS?8R6A^;1&I((]X0g\NZ.@02S?-@TOAN-I(2\0ZAZ6a17WeZWQAAbJ_EED+3X
(f+Wgc4<MZ8]OJd:LbE,YD)@S4-9<-N=#TZ>E.M)gXPVV)(W);g/F\;/6DVGJ2,4
\J^/0L6f)^9DQ:b-E2>PX<cHA3-1U?Z/K4G0G[,bF^E?aVG&Ma,+BCd-SDMMedJ?
d^<ATfG3E-)YPCK(D?6cd+\YNTRXTOgLHPX2F-GQ3Of,gJF\Q:6-e,Q.,B01R,R?
W7KfJZ8FOJ9g^S5U2I9TQa@G4Ga,YcC,4LRC,DY-K\F\MYOCbXSTW7Ie6Y^24HNM
,XJc=W+>VT<7Z+ZQE;YJ2NL\0[4\^,/f_M9Y8YWFSb]^=6c+T/AXH;_0#gG]^gY?
_]Mc&Y3DM16H1.>O0QJ\8<?Yf(g4Y&N)B+@1^H\.LV=/C+N8K.H6^H6/7(_+WTOX
\HEF,.afI<WXY_>1.4#<COfCfcH7BHQEWcCN2^4\PB1A9\:;M3GW90WFTB#EK9-S
:7SZZ)WF#=B5;.:PMf3#G;H+43)/Q:I)VLc);D[+\1F09O\NF;8+D/ED#].3@KKP
4gJKP.PfL+N1DW/@D(c6MJeV9#D7N#?R-@eP6_CcMeg?D3)f<4.Z4)4fB>M\8=C:
N?=/3[/>.C>&3-9KM<U]^-8>&O>3bOU.>:g_V/C((,U[(ea[gM32OV.7]OC-AdY)
83BeSd5_6gA2D^,SG>X=.>P+DQ(La)g6VI7^6(#Nb)7II,YSdQ/gfUVZ#IWXUa\X
9>/78e1O=4J]B.BQ1QZ_e?5?b5LX+T(EMHaU9;&eb@:5DdPOGQSD38#-OF(a3-2>
4)eI4:>S:H,:A2IR,F,^\95;46OR8cQ38D5OTL25FSI<L670D(b^f+7F3cVOcGb&
I_,PWL7ga7/G:S2BEaZfHf,X56&<3bPVBCO6HVb--<@Q3^7d597:<[E?KMc=/#ZZ
1[F\+DE(&?6IA>^#:X0H?9<(FS7-5:4<K+?_MLY0FReF9==^g;2Q5C:)]=VWB?9)
DHJFE&.-AX95MSU?9()NWG^HJCCL;@0ED/J=Sb@,YL.:fPWK&MY/Q,+\X;OfYI&V
J2##c<U^BNWDaH#QGP.>J+\(>BEHO@3)<0YT7R3H:\/@AK_R(T/^JGFfa_9Q0G?+
L;TF(dWC]#F\AL.O+.I6R8\RGFUfTf)P>@PE@K^)d.eUEZ,(6<fa],A2J4SKJL@c
@J2M.6-ZYf)2KQ];U6>6X#F1>,IUaV&b@-3HBJM7BZZ&D(VZ1JddH]UU485gX0H[
6X)aecK64MLVe17K3O_V=a8Q&J9E(;4@92=RV4PHd^>K)\K(3,HE)<D1O;@SAR=L
8W1LZ@/NYY,IQ&8X>&6?9MEeLMD6_U::;,V/JQ[a7?D]EHBO0CZKaIc62JMd6+G\
f+911d.8D-;U_ccGLCYMK9K4gL;08dSgDG4D&;(eNe^,3/1AGB,XMOZ?I-@-LQX?
KKFPIE.GOZ&eYPBcZI=^]>2@LTA85Y..Z_0,FPJGYR05\70KDF6fLE1/)^fERUgT
,(@ddYS6Z7bAB]B92EF1K\N?:)MXI0^9]^/c>)RZ59f,g\5H6UQK1LT35D5gCEJC
M8aWFJ?accfHIFWg;L[@gc=(XSTJ0QV9QaJN,TX,TU2]O#bLJcXK4RgHE5Oe33@4
fZJ??S8#E?,0c:H[Sb<GOL7-H7F)I8f&I1&0M).&CZ3[;BJ5M.3\ag[@W(P&R3XH
fcEU(F1,C_L\fILP,D_)9)c4KJ&>^_Y\F29+90,EFUdXAK8,b&;LX.EIU68Vb89Q
,.&,SPQMX6RW,g,.#U40FdOA=BSCWag.5E;@N+^c9MAa)9OPU(WAQL6ABDG7XT3S
@[;W<^^)H4T;^I[8R7G5O_GSF?:8LCCAHBQYeg9fUPc4DfT=B53MbH+cg1)]Y-bX
XQ/SIY?IB23/(UF;BYbI5BL=ULT)3eVfAKLLT81@25:A0b&S<TR-WcF>I6@XGeRW
F(@73[MGg/GY.,G=-+g[KVAb+,#R\PP\FU2BV=C/&L\+/J34d1)9@^>Ya/KWa-<D
@#D_UT.0AU2c6b\WUM1B^D)HD/+e[BT7f(3dX>F8O5H&WM,VZ,Z#-\HeW@@Le<2g
R?^7G,1N\[)cV6:.YTR^C2N/?G3f&,e.gGGP#Z_.dJ8gXQ3@-5>CV0gC;#97Cd;[
UYSE.?8S2,:a[92/6aA9aT@Kfa>c,,[CR9EQ3@6;GQR6F8Q?U.7)1g<c/+dWO1TV
KD9SR66J+cLUFBB<1R/K=g=^+<CWVa\OWc088eX5WZQF)Ag^aaRI-/>=(6[cTM]I
b1.+cJ9b=_-3EHLQWCQ))?[J1FYC3]S;NQJ>)-UBMY/4^-CXEPF65ef^9+&ScZfd
+T0=X@1/cC@_#&I/CHc:_?Z997#-e<G0.7_YD0\1UP<eTg]KBfNJQdY9^6e<eC+_
MV]DUQ&3UdF3#5/6g8C>6\ACL0E9d(:eHGa:Be1#2d9.&g+H&9E5RbZ0?H46W,E;
1^-<(L#EeAd8[,+..WX;Ig)C&?)B6J]9dPa#ee_9MISaRJ0PdCaP2Ke5.g:..Z)3
7Sd2Q]6J.6V?9Og&J[WA6?+Y[1X\F#PI;2/,.I7(bEggOa.V6V-4:F/WT>(gC>44
VedadDNINC6OIfE:WV_gK=5,_M\)&/:U0:b?\3.IdC&D9QgG/eG9Da./R1RK@4A7
dT^2K6OMGDH4Y8#DUcE\79b^6d?E_3BXSKa#-IOaeDa?]cR/bcM)fc#.2[3FPd;[
]YSQ>=J4?9#,g65>[6C4>-7SIMcY<T17MU4fPg=[:<7>[&8X3MV7,+AScG.84#@:
\g007S7D::&W+R7YK0JPBc(T:ZZXfeEA3=?+PMZK#MKOIJ7OOb8PQNB61E(QWb>V
5HdbZ1M:_0^ZcIac5+PB^20@?XP@&YSWEg9ES#CPJ;]V3E4998O5-&,f;WP1Rf2f
?)]8N.GcD#S/QSb24AINSHHL\;-dN5KP9N4P#+NBSRN-JdQCCOO]U-3ZK1?R34eR
J<P-]FK7dZ88,X)\VWNQ0VL9VGS,+]^1eG1?=M]^E8\<<QT#@,WZG-bT^EZg#3I0
>#\K3;+e/Pa2L(5DcTMMIGNIaN\K59]HZfH)bGI49?F=:#+B/30NXMH>7;EW=>^T
.0b00e6GFF?HSFJ_,cX3G]geScYdQPd\1gEBRU_0d<[-Z-C0=RN4NG9F02+SCDLN
X_8JM[Y1\2;Mf]fOG319LB+8fRR05S#N]bY374fU(gY3D=WH.b(=2@SJNeSa8B6P
gBHLDU3@Sg1/EaB:#0f9gR(7AP^C_;G2gRT9)G]bGF?&RW.7:UC2:4gPC(53Je(V
XM?CXaO<b0WF^RH,[5Q\TVE&DS?EYQ.L^dL;1\g2:?D&,E7C[dIY]e6_4@2>fB6<
+OIZacXX^?-9d-D3V#fcXe^b<=UIK44E^1WW6c,R#UgZ.WR_UJId-d@X#T3fda(B
W[:+LX(8c/A)?db)KeH1;7aLa6#2eI(,+9X[DO1J?CdW)6VYR7N_D23C&#1c5cQ\
NC+C+,Q<<,AF-+<7F\,=9O;CIMU,.1YP<WQ\AEKe4bNK&5=MJMYEb?K)UJeW\[;[
XK4/^;6G.Re&c7[D>C/M4YY5FX?;LgA&\LaL]L,+7(4Z:2@Ac5T:_.Ye>G:bANHQ
KA^Z8UBDOUT>bZc#);F^URXTLX\;M-c4=Z1F-g22B-7UMOY&G7C,(bXBN1898I;&
D@9HJ)S4_dCAN>5-eGDEL-(RMa>R+EDHe0&BK3QNBJAN_JRbN_?Q<P##F@bOL??-
Z)3]#D98d3\[(d4KH6GX^X^#;YJ<PU)-@4Zg<H-UE;QJ41]^cZQa?/OdAP\bgK&(
BaGe8(d##5TK7,9afJ7XDOE6J@2fBU.:>cZJf,0YIR2aV+12+GfT,11R/\,(-R,L
0Nb]O_]1M&)eAaC_#JRN\d(Ta^L<g/D&G]CQG6+[PeGeCe3@39>cW:A<5VZEZY0>
([;\&-71Fb^MQ6^<g.PJR&+M(6X+8<F;1e(=LVdL>bKI(G-^/FS,e^2)fBC]2Nc(
9L4NY##Id&::fdFdd6U4W3O>_:1OUccM_S01QW4e7JBB3)3Rg79f=Y\<-egWS\PM
9S0^Ra,,F+N9\P^1L8?55WFE4PdDNBI=ZJUX49#,>Hc3Bf@7):>e<CO:^eUHf?M+
3-82@66B5_^GUa;G1L8+>cW-F79)9]_ZBDHTd=.T4POJ]MO4CN:1.1J,)Z3_(gJS
8+I41Ea?f6WO7M=O\75_XQWI]\F48B+J57G0/P807R9d],7,LWbeEJWMG0F5H2e1
4ZbP<BX2G=@:3XPMP(?Hc[D<La6?:Z^DP[f.WR>Z(T/;@4^EW3Z&[a+#Df&T>>6C
9F[K\A=(d3\OB\[I+3C<2d4UYb]9g4M<W2AT-VdOHGaE>(d4&>=VVf9,X45gX<A.
b(70:@8b4g>T60d=K\7F^fXWb\7[NC:#Y#:I2--Q-+C<REQWa1&]aC[1?UG2b&N9
M=.d7,GI0UVI4XF1O/9@8QM?PO9LYR&aS2,A(MUU.KZBL?:T+<>:PV02UV1g8RW3
ESIf6\I>@?gPKTI#K=2?a<cO;50G1PHC\IM0OH2WaZ#V?,I#&#FP0Ha<&HO^E<5&
CaVC>74g=bH]CP22RZA98MKHR.\X?6GQ/6J03V8]0@eAP3XS?Je=_ITJ]d172F-d
/6()58WX.I/e8I3HP4A;K8/b?3(;WBU4>N2=9TGceW_\1/Y[9?X_1@Y(Z3/_V5[/
-6DCBHPNeG7&1_=;>QXC2d14)c^=TLJc#;C&W6WB&,=CYa,ZF,C;<\^\PG9Y+/T2
UDa>6-;JCT&74_^K?@5UC]X8fa/A>^\\,\KfB;Ie)0QdGJIY?5>R>01WPI/>#=QE
S\FY9[9U-ZI9>gb\>=76b7]HabP_P&UPd:J9]_C-LZKPI+A6FgCWM?T?a]?@R541
X&JQD.9==P4=90b:L;A]eHMR2M4f_@S1\<1g;(C]:LASbX]Ob\g_EL:_&E1^3&Od
PN^HA2AK31>W/5JOb=;55V<Ree>^\K,a;bA?9#aK[E-F2,J@+eWO:Z?MSZG3+R3>
ZdZX-:D<[F\9/L6a09S,gJGL<7>S7?dL3J?JBSE_MR]eMNaeBbcWDO[^#)0PB^RH
TZd2/E>B]4P(3X>8eZEQbKC/)#KH4&F.cO9:NeaQaO9/WK/YEfR39Pgd5K^/bW66
)M+4CPE6K-3B;?QF8eM3&U?Mf^9F.eFdeVCW:(F@1+(M8M#beC1-)b42/:&[M4M2
XUg<CL/<^4_g5dMSaCBF4-,-266OA3b/?g73JR4Ga@3UU\<<bPQ(K_]P+P>B6^.J
][gU-5O2UJ1WBcQ,UNCT;I[(><6HbGD/+Qg5AeY1Z,/H/B_A+R_BMV9McGR@QL0I
_dDL04:K6GC5C2_#8WM,NIe_5Ob;C,1>G,,M4/(a/e^@-/W8GU1,QEgWUC+\=0X/
<UO9g)H_0).XD)X\U+9HF98M#@&O=-f8AgEOV?A^]--IXT:_\UDU(K1gUHOHg.a]
XU_ITM8AW@Kg?O8Jf2BIU_2eC94b5NP\g_e._<8HA]_16<);>P4.<UfT).+TK9.<
<M65_\DXEB0g?@fN/d.VZXgbNdJggG<EJVFT+DR&+R6b.Yd.X&=EZ73Cf\-+aZT(
_,O;+2M?V;C(H+O?>7QF0B[,?;M@TTN/M_\XOSKa1_-KY0AEMM?DSc]9L6=aS\OU
&JE3]#LaRL,FT4E2UF^+A(^\T-([7[,\W/FdHVE2EDPT-WgTb(T6JHK7bO35DW)0
)L^ATaHgcQJ+61O,N:TJ<R3?<?PJ/7:=9R]G0.2Y.eaFYOG/ZRMD,dXYBHN4&eCb
K1AS-4CI0M<=^/Db1^f&O>M2D)#?aeM,&aYbA[=fD:AW8cJ6H\PC#^S6cX0aFBA^
T0bB4.0&Z+7+:1T&5W@-3_,OA7\KI=A-HOT><.<Pg(Vd??/4B&2OIG]4bb.?2.a&
Kg=V/A7?JN;]UETcF[GJ;HLgVMc417C-Q/^53GdX_2W4D(UX0feWf.bfH5\fe>C<
./D7=\<9(P5OV,cRJO?3=3f1f,.(.GUKY>[8S(&=cf-1>I#-R;ID2M@[a6+&B4?_
7)JJ#J-7VH,T9.f3W?c(e8\D-\7Ob6dLI\BS&?;ONQ8)F&6(-98.P1@9>X#Ga2(4
#,cc8:8.gZf:X2#c\;+[c(>^GKe@b6G^AYZMI>D-F9ED0+&2Z4[6CbeaQXK+KOQN
B7(-fS\;0]][/6M@96aNQF09D,G8gYND_eFOZ=eP-D?bTAeMM&2Q\^IP\GR^U[39
>F8\aVFB1c;3Bee9JaAC(>P;#[LU69J?.D5[,QFH=NC@.AA)La+//Q5&;-+4ccDF
bJ1MIOQBe-2>I>:;(;F,J;7NfOK4(Y^3P80>1dR9?,#IWJ]+SY/+BGA4W(]-X;85
+9ZW=ISEBVVbJH\SC^\\:NC,Se].96VB(-<C-@]PK^+9BYH4^1R<>)ebaHW8J9;V
d32W7#00/>B)[U@2c-#DJ,S).Z]g>[;eMJb0IC[DW\MA4SEYf\F_+Se@Df&-,UN^
gL^:>c7DBQd4:]T36JP3Xg0L-US>WF;?VgD>)^;_@=SGQH][Q9#,f@YJ9W,6Ab5,
cG\Xf2;9D1I&F\_aO]_T>.a)L3dC5XUO=W4(bB^Y7+.,Na5D3d@.XP]U3VH([6(-
NKFJATb?A0S21#4g+?V60f8aGIG.+M2ZOL^-]L1>;##,J7SIHI)28-acP+bV[X4W
VEM7.6R+;@g.5P&gOQ.JLe(\U^H/&WY2X[f(1\P\K2(UQK7A1FHM)#gSc:#[L)Lg
E0UWg>N][AS7UDZ)VOI/=b3Of0>\.C-E4#WUO\3MGGc1#bPHP<gZ,79@ACO4Z)?#
T^&&+K]Ff8a/DV9BKb[ePY(:FFJc=ZMW2SF-3B<Ke;Z=4&IO)721@5Wge8(EUaJ1
)FDTI7N(NcE)9[K;>J\O+^fSO8JaV\b4Z^^-gefDKdJ@J#--BH3Q_K7B3ZIQe;ZH
//eG#3+]>DCBS^<(\ROCLKg:W)1fS2A=Dda#Sf(4;4IU8+5\Z4-8I95N+7[IH&<2
8HPA97PM8?2@&dX,;KJW3;A[@;_5<RGA77VfJC/:9Ca3##WY6J:+>33.\;1>^@XX
d(&b=L/:ZV3cg_)<N,.4^/>aH21YD3]Z6:I]:f,N,Fb+\0A^XMEN@XC1@-gU;IB[
],_M&B6/^b9TY3@e:7C<I0I:ZN<d3GbGAXM2+aJ;<IOM7;+=_U.:a8G86]dAJ2J]
?7Aag8JV+b)OG(HLR0B7,>;RK;5X#[Ub,JbYN[\ccd?_RN2R/4&A]3a;IWc9J?Ac
TSK0f9;T<I1+]6PD^S&7:8b]#fRcHgV(>9X3+J80&Y)2.QaB>4SUO7[1I2</dD?U
KJK7XW;Q(#+KWBS&?@/KfS9FF]A-2&IOO/>81G[6LTURM.>BJZHdSC71A2O)c)fW
7#)HbYGHBQ@/,&RVG)+.LZ10<I?a/>GUT42AgE[<E@T0QJQ42O?:cB1L\94-AeR#
MaQ(MR]9]+G#5;_LZ3O=1BF1T(R4PP<Vd>A)1cC29;#0@H)AWQ7IXaT\GYc<_c3M
T9>R-.fC=#:Q;N&Q<.;C<NHcdP.#YWU.JaPI7W3:c:gK@6_Z5G2,S7FT+02E:,Y:
PCXOXIYCO9^B@DHA7eXFP#;>EN>eC,U>3VE(Gc8EJ?Rd\&O)RJa+-aS&dG4a(V4+
ZcMPGgDZ[X[D7[1Fcf+PHKTd1LQd?;b98CUX]EM&2=FY_ge_B,/2=\+F^><X&91#
MOZDZ9DeV6F\)AA5eO#]Va4#+7>\D<A(@T/[J(92LV98M/1/2cP/4O6B79bW=;74
+Hc@AO:QBR;WUEbY,L_NC8-50EQaTgGHERX^\W+g_?@AM+,F8.3Z(2>SKHV:g&;>
Z7FXFJ[O&bSaC]>0(.9#MfdMe..D_K9ZQ,,DQKY?agAFW/MKJ+Z/OT^;[;8@8:=:
_:#1:_M,HJde<GW,S)c&aA4@>43XC?,/Z5]2MN<H\SQ&U7A+.b?NRG]@V3-Le)3g
gQH4HdgY?UG:DTXd/T(W_P/,f?2cUTKCODIHWL5,4HGa>F+?BU0TNCSD,@5B<&@@
8VQ?^5LfUPE.71]6G[Y2Z>C6WX_5DC@-\GR[B+RUP\913\f96,0fT/eS7IS>,=YD
cZOIg7dM_9F4fES#a)Re,QD]I9g8+eG7YO&_.ZM=MdO..]Qg[]=MY1&A(1=VJ8;<
TL1Zc136P0NS>[/?ZJF]4D-+O)W\ZFOND<:e#:JID/-O5R35<<8.d8I.Z>Ne4+GN
eCWC2@fa(VM?SJ9S&Z9ZfONdG<RQCCRdLVb.AU6>/Ecbd?fJe@XS91+]_1I4->V4
UF>6PCa0\+@_PJL0OG5:<a68,:Z;L_&AHN)DfQ86[,_c/-5]?;g(>WH;MM9P1ba:
2&GGCY2;H560-4<=D.e3(;H^K1ZDc&Ed:Cf19FE.F^dU3@S>+gOV6AU0(g>G&+[J
d\[S5F&Z,2J.(6+W2<PLP/g\I:X,FR&3f&DXg>,:BJG@FL&a1#L:.d@)[38Q;QJT
=]AAC/d_))eaD.VI>ZPZPK7d(F,MI>9JW2&PS2M_;Jf?MCg_+L9PVY,8bKPg(,8;
aT8DTS3T+T[b@5UfME4/J+\><<<C<9_Mg[T,MT:KP)2RVX>28=NI?]IAO+]Y?0\M
-R49VA0d1380@604IYJKL5X17bN(N&SC[W&G^#ZE09fKRFQ))4aJCHSL5bfb\e&S
3SeCI)b0B,eTM24KD_eJeL2ec,SBd1LP2C9CdEIX#:D8e;D\E,T:&6MV7J4bd,DB
R)F.+C7H[K25P>Y[K+=C),dRW5=6<39U@=YIc@fV)dL\c.(+5@NW<&IN1O\L]\Bb
^OJ1LUYTY>@/P&)_DGJ1ZS?7?EYdT/&D9K2_#6[M)5L/C9/bHC=D?8MdYJ#^C?,f
KOK]3Q?Hf(YG>X5REN>5TJ:PMA-a]T23CdNXH[A5UW/C=.1/P)QG3BF;RG);:6D9
F=;af/:>GEKc9==XI\9PTGL8GeLQZ;TWfSE[&+=(NR@0X;W?bZ1ZG:WD=>Yf/_<+
OZIedQ9^LUd(PZ2eRFUO9b\Q]=G#;F]C;fWT/c-@;Jg[3J+_;]3-g)W.P(HZRH;/
VMU@=,+1)-)3E5FPWcE(O5+MI].BV?OL<<1^(IaEE2c-/YD1+I/3S;&=N_#:@@0>
\Q=YS1X]DJCL#+6H=eH(,N<,UM4CPJJ=SU(P=2JTN^7\C.-cZ)cTHX(,)4I_dZ/T
V3g3TJ1d3J[Q#DAMD\H\e<A+/>),&6D5XB;Af5d_@;FdSNdTEf&<S9.A_<\N9W>I
eWA[VH@?@#/HcHJ[)aGE^ePf04GH9LD0TTP^61fJ0Lg+AQ&@I8^dMYBA4@@Q<FE^
OXSXT1P0Mc;3SV1<,_C#;8e^5AS+fDI\W0BY-+8=&P1;[-APZF3\[9B)ZR13]NII
2g#Y_8@^DVM5g\6<[ZDPIP-8VgW/ZeUe@UUe^OE<)eB[#5VZ0.?dC1a]2C(M8b-_
VZ+aAWdF-(&#Mf<KgU=g[g8SYGTc&+]^CO_;c+^34GE?\gf,:)Q9F0/GD:a9+T,^
2PIB5Y3KMSCE;\\,GHGE_X=6JWIX9Q(+0^AeE:L?X:dX^V(TYNd(^,e-:O_R)@K^
Z=#_-9\g3V:1Z1SYK#.67_c+TaOd+H?<5-+<MY+I:cF?_)f6[>Z\@(]eJ;g,NH=3
KZ8=UF4QO^I(KD^d6C\E#]+XA+^W(EZZD(-\6V7Y:2;90=ORQULR#<QcM1;g.6Nb
;SBQdP>Y[.b=bL=Y#IE[70_I3QNYaZ#7AZ:Q^=,g^W-71K+=,XVMNNMP^V2.42C>
T,(TI.TaG2U-;PaA^QQX>H^,^5fX>HOMM7aJD3KgMgV#PMYc<6ag(<IZMW><HFY=
84\M7\>=X\dHXdLLOeK176#Le]_ZG+4?Jb.ZSFEBf7gR&9@2EC8@:\YVSO77M42d
C-.a[A@,1eJ3TP0M^^eVGI#Q@O><W=8VbKCbL(P1:<8g^:d3CUdT.5aaf[[d+e;N
CB[+#CdFd).R,N+VaBU\@[,fID7?SRg+>(81JD\OKUEGK6c)#WUW83P^H3MAX8NW
Q.gM1bPYTYa<)EY;0+_S97a+Lc(GCN,bYeP;5L+]-=.22)fbZCMEF7X^?289f6Q@
N[\N-6S+N@YK7,JOHB/0EC+P6<e=5_)Ac2OcEAAb:]DX0XNO-dTD;AEQM7(B9T<&
gADPVU9gP+N>(>36-4U8Z-&@=.W,+[12\Q9RI7KV>.41@TbS+1X[OS]aG944SLF<
XQg?:I@WB2,DLA[:IA)Sg,2\U.CbI6QJ2N4D4Q&V7K4#d^HOCUEU6,B+1-68g#-;
(e6S?^e0>b7I#C@@X;TGJRFg/+f?C^2CMaF(56D5[(:(5Bd;(>W4K&</=27cdc1T
[gXN0?I:+#D+H)3;P+R]d&SOV&W30H&\;U]Z+LN[b^2ac.D(9E>A=RS9Ga)JP(4U
Z/0HF_-V&c_dKX2P]KFSKF5N[a#eLFDU/=?3BAKK8b+K_1cfIYGEbEF1C4P.[Cc8
e(+KDcWgL[#NRdFZ\T?c,+X4Jd.I@QId(A;G2@1NLM;,^8+?@Y))UB&F0YbF,/FD
V99&A?W;&W/;OPH,^@A]e\DUaE,_8CUIDE]dU)8>Kb;L@7IC)C=-)(Q?dJ].9MC#
MS4,a.O4F>=P;BI/Fd;:eLc^Ng\,S)W2&P7R@;QQ+QG9R_TW5Z7^G/]N=L#\G4:;
eE&FMQF1YKI^0S-OVVP>S,8Y8_MZY]:aNK>4:c\a-<1NbTI3:@8(/K8RV4MC3YNN
R-822ZOS1>@61NX6d9EK3N]_NW?:[g0a5SDU494?08,6?RM8X544[^CL2^eY4+1:
S8#@#KU?[E_7fcI/)G9H>D+7=6DaXK4)8;?CTEJ#+CWT(JLUd9D2[=0@c@.Y.F/^
=<MAF,P;1X3+H)7b4(QG+<_,X\C^8#LLdG]3,T\Y0-e<S^5^W#M6Sb@,E<[&KfJ@
[)YgTFV.+E)I#HbI:-PfE.+>I)YQY.L\26#&TdM<F?e@#.)cJ2PX[XRS=Z/0CA?b
X/\L4ND]-[H[8HK8,C(eB=eQ+aW(,Z<&,dB03;>bX)2?NZRWc/)^fdAN>e?IWQ&7
/W]VE@>e?\+EY,<K-7L/46dV]2HHOd]5\DQ,J/b+22La>\KP2@DC>UfC)OJDX_6A
c@WDWcAe(;;6/Da:<CZ#gJeRSL)OT);+ICF&fS#?N)BEffa7&[.KEAe>KG3A0J+Q
N#-,QIJ:g>WDbb;CSBK(Q4dJb1F:ZFd.#)I7I/)\@^2<6O:H7cTQc50SgbSBD#1Z
(aT4981X5M7&?WFSH:676^Cg6PVGPP,LXD/cT.N]>#W?DZ^EUGFB6_XU(<HCa:aF
0]S<N7YM=N@AX(Y+,HW24[+S/?I;1JVMf<d6a\)5Gg,#&CGXGQ4NMc.#cCag9EH(
DTHeI<Ze3M3(YZ[:PWZD:<Q+C<Y<+[#L@5g,G5/CWQX^@CbE)&CbOfW&UW:F@RY6
6[YL#UHPAI(WTQ2<2/aQW@>4TaHAB(F.8L(8L,5Ca7cfYUeCBTNOM+^R@X6Tg:OV
:\gd9A+.gS&@TN0&B8NcL5S[_DG,dd6+VM5PF+\A(AV399dW:fWKO-(U@@3LC>a0
)Q56FWa4UF@U;5I->PP,C\2aV;^e4a<PIY\5PH,+1-U70U,7<8TPe5R,DKBH,376
+]P[BDT3KaR;N@UN)\#cM&U1Y_d93J>\g4];J0O]I6>Y3&RE7[<0INXZP\V;2LGC
CENOE,2BZ^[(Q9@BVVZP,+F-c],Id;,a@XYIa/gNeK6YOafgZZ3<-M=a;QgFFE5D
5eP#(bB+gVF=[&#>OWDd#ec<,eW)cKI+9<FJea#DT-]7,J.&bP=Zg0;)dAO])3KD
NJeSX)8La=dCE;<K(,@5CNd;>cgc-CVPcS=eG5fRO<d_5;g[C;VP0JO=B3G_4E^S
S5c8MVMb2)#\#:L/];-@?H7/M_:R;GWK?FTgd(\/3JE.A7LTF49_SLCOWZXPU6g5
+BSY:RAg]<bK+;YESAZD>3/^@I-c<B/V+RA+)NgOcROF4?:S,(g<RHRM-\>g&VXP
9(K^>d>UAUGQ.gE/CC0DMHXE37HJMD.)(KA&RK7Dc]I#/7f9/(<V:3f)N@PF<5VO
@L7OFU6OfeWA68>>a<4QZ0:;gf9)]H(E@P?\;05FY:VdG#GNNdM/H6[?Hf;c#==N
afIC/YJe.ZN:SKK3N9If;C06<VDN4ME5<7813M8X^?MU:+4Rd[MC2L@+V>;W5W6f
8##:YRD9D?YE>3+SZ+/g45QVSY7A[=PIQX^g<,e[G\7CbPV>D>:?4X[0.>).@d\\
Q5a<[AG5a8^(,[@>)6a&D:J#G0F,A[I9T^b/\I=Q&fG+dcaH.>Z1GZQG5(:=-7K7
^2K^+N1M\#ZGNU<Z=&Y]?3b\:YV+E(TPcG0@-Z1Ze&g8;AK(eBWZ9c_NP(Nd+K=2
>=2D3TMGCf4C6,6?GVF5H<,X<?MBVG[HHFeX/6+J\IIGgR+Q\Ab,.YcKHPf@6eKb
fXWJ<0b4DR=(?8G/#69-Z29e^c^\P<Q?[JR&g7KGC/I[HMT8<FBN6GRP?J,]K@a2
/NT@THFZA)AP@#fG]g)=O3)HJU?_40D^d^@1O>0g8U0_24]F#Q,CESRg;3egLcc5
A[gaU:<>U3b,U\-bQcX<-YV^e,cFI3:#]/FX?5Kc9AU6D>LcFO?Ygf027I0?GAd/
TbFG/0RX&?-+^KO?8A.OU,NddMILZNb]^7Kd^7O@D&PX?[HY[VBdE7?T9/Xgfc8>
;IM.32bg4LfEDcKg.\f,[D?f4ENW((M2bW7C4P07)XN-4TKUcP,R]]4307-+2FXa
4YeGYY@a^;/G#_]RZSX>82/A(f[BN&12;8W--YBa+dSS50/5b/[2R78:,P?S4<gW
-CT;4UNUDN19AYCJ,-X-?#.HdN51IR7/O<:-U4+b?)MSC@TD?[,\4dd;=81)8Q(>
/e#-B?<#EU:P-SGgOR:^[QLDT/MP]+Td[e)e6Xa<:?8^LMdY;IUYT6.TXZd0+;;O
<<a6JHR5ZECFHOPL&#GUbYc1]>^B?VTEeO&KY<S?]LW6:SE8M:gRM4f_,J8W.AX8
.XdNNXY\f.g>:N&_6X9NG_MNLUd[B]OSV\:#5KS#bb/9Pc1W?\@Z#-:ZdAC.\fCW
7]gYN2dNKc)&HD6.>CJWE6FJB12=c\N;PWFX;dX(\ZP]NDcQ&TCO27(:6L;LC==c
;_A1-^L3geM+RW2JIO;PF(OOL^92_6<Y+HIg^C#+Q@TJ=c^e[aX_aLJDH(3Z67AH
1.HKa45(L&))^PX0,I-M7?)0C24/@0FbXdFF=@(Q:V6a]#V&Q(X._\054ZYAWK;U
=1[.&L,#3Q5\)Ug]T45U^Y\^ZJUG<WKfeMUZQ<:7R70WeR/G_cIE6D:(>5B[I93F
#S[_K&dE6BAP6@J6/RJaUX<QW503APWA[QG6>GdC_&1,#ORIL.gc2@0:N[Ga>.Vb
CIF/;T>Z<c)d2b:R.QUMS@BA4DGE\46[PKH-DV7[<TR<2I@AF/\:SeM?4VTBE-e)
\gdd_EU6#PU4_&QKa;7]GR)RGJc0]93D@[&#[AO#:P^X6;TQ]_/:N4?Oa/_7<&=3
Hd=8_=,A?7KDDFKAgB,_7>6gG/\^T.#HS9WS8SDEFUR;=eR?Ff6RT:D\HQFdbX^E
1&3A=HDK2d.,Uc@VL8]7ELbg]7(fN01^6#RSa=Zc86UV#)gVJRY3c.9@85^_c6A[
(-4#./YV>O:Z]RAS5^M<#VH:bE<3K;00c\#1F(aJCe):W^T^)0\CB1cD?.\TG>QR
&LFV^FM+:2H01>.fI@^-0R1E]IU-c34,\)]^2Xb]a_^U2Q.3L5?J\?aVeR>9f4RR
gWdPM\Y3^]63<bO3#=MS>#,)\Z/<O1EJ8D_4NDeKOZ#U<0CQO+6N-7/E99XT9FIK
LGWY+?<+T8>6IfQ1^L-ETRI(GB9@T]0=/))e41(4MGMELRH)1+3Z4:H6&-g)<M]Q
WK+L.5&#I70d;FK^SGZ;MP9+01]2CM2+bFZa^U-7S=N(L,VcK-N?L6Y.Ff=D#^Ld
0M(ba#O@Q(dBCI-a@c#I1d&HN1?#CBPQ@Z@6ZDGcd3C30WPH,d;4,(XLZ,bZ^RUa
R42:2LQXVT>Te8U7N4?B/(8Y6RW[8\?AL8Pa,.0DWQ)1D#Ne)2Fe#6]26DO2)IC(
LI#X=.UQSGRM=GPAQHCC;CDEa0@M^0SAf>-E^QC^CGS?@\YL;J)F&T-L,,/XfS2R
WDBRP)40;/]-\>\ZOS,;/4I7#]D))d?8D\L]TT@S@1+[P(K2+DB;ULL3\-4]g)\#
]>#^deJ<BAV40BG;)=CU]@P7IBJ2959X9I8IC\1.W0B4OC6:/JGF<g2GU=VMAdWB
9#dXcED/FSF\;XE(1bU.]3&U0?<D4c#>1cV[gS^:>^.MLAE;b?OLTRVV36.C0+RX
2Y5O^/;1<BbE;^[8cN91[4c1V93_L5\-[)O:/a35^L@P(5TNag0-Le[A^V_#]RSN
./3@\bWg3]9dD9?.Y:2)014E-2VU(LTZ&d4eP0?<9GJE3-++-5>GA)?@eZ;[QPDO
S3DS#6,QBM5)K37MEL8<^:0Z:g+3VEZ+Q[N0#YGYFd3Qbf4>^?LZcc@I-F5))Y?I
ZD.Nf7K_^DCMb]3bDL?_@XeBTJ9@:VGO65eY,9JG,e9@c2LRHPIg?a20Y\IMVE0Q
L-WZg?_87ETIP0SV(f^7AX7H>M83=]KcF9c(1Dc#4AU=JIN+4&;+F[f(HTZ&V\AU
#&a\B#[U<Q-,_5bT_OfBT<d1AFMBPJ-<-:J=9^OIB((0QM\\O-YC]dQ#=_IZYTO5
ZJU)^a.,TI2Y+PZ(_/^COESMG5MO,(B1,#)We.[C]e&e:<\E93Z6<-,:2NcG1DG=
(S?IIBXKOG<(_;)FccWFB(4+N7eGHdU:XM@QfG9HZ]dD)]e;2PKgDZ3H526d<8WL
D\?V&:59b8B/(0=T&P>;LVCE)b,->^CYM(3VUbfT92-S+7+Y_1[#I>>_86Fe8H(5
&bI>UCEDM:7W@Jf0@6K#&U2/HF]\(:4bCF-eG=+L]/+<EQ(X&D1Pa>N\&L4I10SA
/=&A#S>Tb_#?D>)\c&Sf2;WQK9IOT+LY-AEB@J6N2aI+#.K,/D5e^&66HE=eeV=T
CgS&AP7Id#6556^:>.IGYX>7X0#9&,Ng)<NHOaE82I@F/9+#BAg#9_:6<W[a@W+M
\-1b(Sc8GLgRG1&Y&cf]H)/bbH>-XFTS4?8>U0#AdV043-;9]QMIW(MU&M.TL7g.
GWg]-U(W2PS#,A\M4@V6/fZDcacP<)/<<OC(<aEB/T^OYc+3C\7Q<L#1Q?ID\f&D
0=4^S=]?8XY\5<L>:BL(0Y9IQ<,.EN8eWBZ)T^<,JQ/B[EEREZ9b@IB)?@><V?^6
IWJ/=8Hc#N/FIL3_&C\ZQTT\H7dfE)_f1[WV8_Q?bJ3_6<S^gDBQbVK#BMg64e&g
Eg)\3PJ69WAUbD9IX)ZQBYM0/;N<\b50RCB9A0M^>Q90e4,??(#fU5H+8)A??K_2
fa:MPdB+@Z/.T:0X@(MUSgA:4aXVdV69X^AK_OA9_(]DZ<7a-UTZY8NBM,9P@O?0
fc\<I6[&5B_/\M:KgXFE<)F-PF/D?N(-C:J_faWY0QgJe/<(\VT>@.D:bB=Z7V81
7/[82L8a+^PK-W[OJ_5H/d\9YS,]4[RHgaGZ;Y&0UP-M[.VA2&eTegX=#FD62cX_
D2O&^EQAU:3&&1+#Te,+1c8VJ<R3/4Wc0bggfMN.>0]@CR7WedRW3cUJ18aS,(JX
(>Q3FO6C\:@,FgK_6AbSB@Z?04UN23LXR17:WG[R///BX7\]B\.2<GWAY?@U<P@>
(;]XbgGRRMQU&R73T3#NKP40I-aB4c6d?D7I\#[[35Ub0.^#\BI-KEG@9H8)a86W
7M@5<C3AJIO:?4_Yb;04B.[11C@+^:bH85NgFQ\YE]&XQ\^-]GS&FFU\NW#\TFId
GHN2\XeJ[7P2W/2YHH(PeV?WR;)]Vd70JfLDfK#=aD:-I.cRGVWLfHN#&6#BOY-1
-6@UZ)NF0(1GK>_>-3B&96EGN.<@.V6Vgb@0WWD]C+1U9Q<dLLa>73->OCU2/Q(E
E;^8Qd#&W(/GbA][/DJAW)f-B4B\CCKfDM3d)\K@e\VJ>UcPX:3AKS0S.BEaLK-d
cg1GVEE#:2S(XCE^2.KV.5-:QQJ;b7/=NA#E^<+V_EHSEbe>gA:\V1=gO2L3<N7W
gZD9JKOb.JB3HLF>2#NE(R)&gfeQZRBKS94Kd]HR+(\0,X6(-AB>?CddP06;fda^
cbge9<-4;?)Xg@U;/<bQFCMI:Q[0RH3M/J_-4:L(9^V_/@c1I-&4THN5L12@3Z/B
GLd-AO5b/=4Pc;8B_J6A:L(QPR(+/ISd9:)G-f./V?FT8Y+Wa9PXDf(2#FSe/K=A
4cgG(Z>-/4+C21NYFZRb+VYW(UMLK8Ab9;6.#]<_<(9(TS5?dYFYV=H2&,1_\-\I
7[AX;0I]06,,:@<<BR@1BL<\CHc8S=CJRQ,0^^DO2FI4af0@5_]60B])N4IKY\AF
-O8C;g)DITc?<.0Q]-H\eJSU#];XA7TR8.X3MZ6B6^X\0UQ8d(V+2dD]BR<fIGG>
/H,=CRZ>CQ&+8Rg)cC.0a,RDAOddS0>?dOBW9G7]WgK-\Ng]&AdUG&==HI/HG06#
+G/G-SIAZ/7CQ,f3DEVU;Eg1\]e8TKg^>;F5EBcf_?@YdRbTK(R\2OPG7&4R;N&&
5S=&&aIcS8H(,8:FV8]S##_eN]:K5[\]]Z43SBRT/1Y,A)1_f9MMCG9ICf]<Gf\Q
LY,1,GQcKfCRgUA?SRgK^P8.f#V&+_BQKD:(?>SaYe)RA-\&/,4I_N-cBUC=PC;@
XSMbVD(\6)JJ1F\&ZXbL[Cd#WL8.T10N/QZJ7Zf+:>#@FdV/495]C^b1N<\;-4Vf
VGO@dUI[S(dNb>CfbHNS)OG5NP-/M?V9ORHDVV;>Q@<)?XX+@]SQU5RQ?6a.#;ZR
dA@g)S,:@b1<,[^I1;OXL0\CRQ-@EO\2+[<e+YSKR>Z,O/2^NQ6&0.fQXI;?ER]D
)fAO8#FS]+8G4R<7^IU8ZS>XAE60@g3SeYe)/BbUg:@X=f?ecEZ;X=(We^-5Bb1^
1WXLFE2?@6D9+:gHa&5),5.#N#6^DDXaTXW#L-6Lg]Zg+9:U>d[,OQ0-05,+L,0D
A3+-P/+g89cXE0[?F6Z#5)&#+cB?T=&R/Q9FeaGWPYKA43NS4YWd&4aMC?6J7JKT
[Y0NPS;&KAEO0Xe+>]P_V<,=V[V0AXRNM6]O/M[UA,@_69U\?&\?,4VWDIX7/S\_
ed7:P6DeMMA]^LVEb,Ud^>4Z>a/JB^,de)#&-Z&c1<#;L[d5c57bT4Y.IQM:B3F>
^FG1QG?YI7cR1?;Gd\O,g]AYKB8gLd,=#bS=R-Y)1,/c4b7O+Z>&XCD_[<JV[9SS
/8/#8.OCK.Hd/g]RZ-A@ELbS#7(5D(,-])BUN4U/FA-.9]?UgO0<&Id:L4-UNIDP
90E9([B3Z2\89^Y9B;E[@)E]H3>F[Nf+4bW6<9:@Se.aJG7I>&4Dd.0[?RFOGOW&
5Q<\?R5EQaJ[)96OX-.aRReVR(1,&PMea-J)@:c?#=g=/14AXPW0#1X1VM=6B:_7
WK#Mg#aSM<4GWY_(JcGKQ&1c>&1X,+04[.c#_X[=4?T=X[??][9+SGE<2fVNG8B(
bW/dJW^<8/OVDRLX.YcM]9b7N(+H1U]9a:.NZXX]P&3GG1&LQ3WCD/7SPd0Yf8EN
4P7K7[McCY]3WC&G,_NDILbC+O69<Q9LN7_\M&1K\N8&,=[d&V=E+\Z4NNVg7&43
+fW.ecfH.+Z,^[Y_]#LJWFGb5PcA:E1@S&e;7Eg2;ae2\P;3>Y=3b@eYD/PFW>:9
ab4OVNa)M?\X+TMRa#8<D2ZW)(@(-<M5@DJ#^6fW4-]H.=OT,OGBU5KGMG7[G2TZ
OGEC\7QeaYaWR+/BJdOfM9UaT?&)<CHS]R02CD\OPaNE?8C92(94>f(IO9I\Zg.<
;+71J5+M\d>>O(T[_7U2?\e4_9M7T@[5XJ=0G,J/CCIWd]3a7cH@E5&11GM;\=K^
O@:eA0+0]1O^RPI#(A4BBC=N,L^RP<<41&3V3)-cPYfNLD^^3O;DZ+_/&Wbd@-DK
QJ-NR:2fAYd>F@4f:;U&0_IJ?(dS68[_b-R1NJET8?:bM[e@4_.dfR7Zg-6-Q-[B
_XA^@6<I5f_B/b\X--0dUL\2262(IDJ]3^N(D?\QQ:<bFS&]B2Jb.B-fKaP5FA-O
FB?;TRL36,f9WOO@e)@.,/MA)LDL2#,^IJgNMFNO;;-R__f_Z^J@)YL16H^SC#;W
UUbe&7X7?Y]7#gKM=^(e4PR@@\aU]-cNB>bR7=>;,e=[c,eP2<42\b_7&97_;&E+
;W6ffY3;;@R1=RY:g^DeP41K@M<2g;JR);:3&S-I.C3DPdI5>UQ@L2JO]6\@42D_
FaMdg3HaWVcOB#RMTFS^&^,Y3UX=,C&_A7:6M:IFe8Q^;3;?HJ^]5:OI=b,#A:FR
XU<=2fOW03==>NEFaE\S>\BUN4M9+8\07)VY)_)aJ>OX65)1\A&)R9?VS8X5?AU/
#M-Fg/7^CBHV?feXE-VNTS])@B>ZOSHL@1f/5B/5Pccf&85;(5-G1\EE0>V6AJ\N
cCT=WRaNIP.T8\OQ8W?VWc^e;MIKV/^+]cDZW?SHG&)3O=SN;gZ51&8]]W\VS?1_
1(gGVRAF5HAJH7A<g.B.e;d-\ITA^\8(gcR[:D[,/.61@W4\/HMVP[QQXMN>-D>O
Tf]Gg9O;64IXBf6(g.?8\E@[:TC/I@.BX)L2YD+Vcf@+^XBT2_GVWCCM9\QXA_CG
gEP@88<0#N.#R2]^?;R=c:T@[GaH_XMPOCV#CJd65)dKG^M9]).6UB;facZXIBV(
P&J@VK[36G5BI_EXU\N@-RUe@WW3TKL2^,e15WfHP),(O;S_X#9fKQU@:a:/aTd1
d;:2&)(+e&,G?#:+\]b=5SBI)0DU2]]a43-T2_NPB?SMYe);e>9](_cUF9-(M9\A
G_/(45N,>9\W[7T5GT^DOV7LJE=U[[U8.9[G,AGJ2X95^/R#-NZ_Ff\cE_28\@.#
+;)WX3O1L0>g8)Z,J\a@WZX;M&5C-Ua8,R_Y2RUNcB(]A(&K]WWY<Ig8UEKLe[JA
:ZEf1]J<(D\95ZSJcTU4U_/R9OQVafY;D25f@-g0b]eB0Z;KB[//@,<)M&U@9/Y+
1A,7IK6VEO(#+5A3NRFW2ND9JbEf3Q)</QE^DYAL4@Rg<g6=b,J+g3e37M>X<=W,
ML.:(59<PYGf#0>:PEO(W=Z7?(_&=cBc3QOA\=SXCgfOd@;^c#/Yc9QK)8E^&dFe
N];W6]HYCa)4OSZE84g^V9/,1IXG@L_)d/PWQ&bR\BDBMPG4;>J,=QV=,ZCG+XRR
,eE@;#-0ec[E&VNfK=NU4TD@<_X?gL_-T+OP#.#&G>9a)4U-YQS52RFCS5d2_AQJ
LG&IQRJ0SI;T:N73g;U_XCR>LHN)A9.7IYZ?a;cUZBHMTH[DK7@XVI(;A>:U\Gdb
5J2,&SB(J6A<1XV?Y+D.>6#G,)1F::^RH[aXO8O4X;H-]\#X?XBTXaX2WYPOSO3g
Pcg&JLFa+4@#(dQT]RL(<6(AL,ZRPNXHc2NMR([F0a95-8.f\e,LJ(5Xg18^ADMM
1X9J)_J61D3>3^,/g7D)Q-Qg\.GZaJ8PUC,7-?P9-M:ZBGSIAD_g?]ec[SFLEd9.
8c]<IOWV[1Z0&A5eI+afM;bP=74]N,I0b>)E<9Kb<?QRd7#+I>+C#DF1d#?>G\FS
@2<Hc^K/I##,NE(0FZV>]OI4IcQ9U.(8=P5dWHHH7G,Q+gbDHN-/gEK;CA_[UbTP
98ZUK&EI/=]<#)(4R(K)K7,7]5gL0eNbbd?e^58JXMA+VGIMAFIUbS+?7P^ZBOMf
NPI6YPTS587D;d>)Q(#?KYg.I,1.M3=K3D3M\)dM^QaV.@U5fSK9:;LE3Z1T=6#f
<=b26VH.MPf2(]G-[SWTbBb<Rb-(83Q_A]WD7?X\KH#O@TT.J+7A=SANN?O>]:?I
YO+_O<b^R<IDGS[AaVJD+&VYPfGU>SSA&;gWCV]ME;g,\4C#^:[K8@JVHDC@BV:1
f_V_4>>RFe0#.7-Z#M>[XA;YXMZ7DePc@)Y0VF(2)V&#GODG\?F1O:eT4\d(bFcT
M-Le9#I<Q&F)ND>f6),D&Y8THa2[feUKH8[\5QJUU9Nc:J01[QgR&.NUUPQKdJWA
J^0B)4@>aY1X49969c-YX8Qb(N3O6.]GVX=Q:TXYYd;M1\fEXXAJL9fR58:(aKf>
TX;]OcJ6Z&CED09:H+JP39b3SA^W(<\gR(a17_a_U>#INcJFPNgB)afgQ76>PgKY
>P0FP)TZUbOSNI1>XXcY_c>T&a-NT;\Za^#eY85KdR/A,Z?+5\_UK^7#eA+fb@36
0E0RFW@VJ?e@,2H.bD71DBSDAKZ6OJ.9JQ9.Y[,FU78,C?;:_HT:GXg:b#ReSHP9
#^b:d\ZgJ(6G33g,ULS;+@W69aHJ@8RabP-gN\>?/695>f[--)PW.O_-T_FTB372
+3Y\DK&W/=DP@g/7a:6G)6>a;H<SC^_LFGCJ./03cNTQEJL&S_Sc[Ec-9:^2XYVN
aAN\a/6/fM3X:b:Va2+XFbOJ^XQM-/&D.3L6Yd;(XKS1JS+L?;M(6OIH;@)->9g/
Y1:Jd#6RDfSU\[aI77CVQ3dDX0JN0PS>8<d&]H<:?1?a92,MTEJ&#1NVF003-=g?
KaJ43VBB0HP)BI=@5C.PTI2aeLA=E)MZ[VU#9@B/D@CE&T+0cCO^(.0+U[?NZMX.
H_=,NP5XBU.Aa\P-f8^g^c(YE(G[)6BJ;g5G4.1g\L^W)ePN76>;MaKRS)f0IKZU
>AOB2T@K>AC2f6[1R/VW/<W<2f,26_07N5d,.0dT-D#&eA4gePb=XRg)H22?\[P9
?_#?g_YTSS521LNHK.P6X[^Wb]9f5)_8Q7gN[d#bdb,P7<+ecW&_B1cRP@<+44/7
Tc+?W\>9V]:f86DD4P[?+c6G4)YObNBgE@cgLe1..XXV0KaZN#2\QE[g[Y=_&,Y#
R8RCBM\>LT-EL@I_7G0=g3PUaQ.gKP\_=,d6WH^27)4g@GM0R?;1<<WZV0Y8Z4D0
JcZQFZ1=0Ab:TaK)N/I8cAgTYAXB5^8Y:A2XAd,(G0H[IIRGHPee.>J>IVJH;=,V
K8KKd&-+8eX#0GK_#EdcXeM;,B<WXf5&>&S-8P_ST^93e=DGfR[L(_#PF,H&(XLb
[]Y)5GY.-NP5IU-_U;)f62.1db)ZeL7Gc_1J5(VXYOVggTO)#IaC7a.CF;4TT0_E
JJYXPARPddIMY,P?D11G-eHR6_LD_DK0aW&#QFU]F5PLa))E8&1Be9W(F&;f<NZ:
20[_@[b^<4U9O)V,BXeDM<8R/gJ@Dg<7DK@7EC?TI\I]CLNWG8LgMa=fI98->5QZ
_Z/,7QRX@^B,^Wc4[AE>IJSg<bg1ED:\>@SI7gcH+K;^W4HM0]#4CaLV0BA>8G(g
eNX0L<0B1-U[D1SL7+U<;HFY:c>W9[g87Cbc6;M9M/VRQ2.Xg366)^bU=f5GL.<@
S7.fDQ3:=(Y=dW/HIQ>?=G3_[(T]?H9.]gKD&<2K?S?(cMHBI=SCSK8gP^]]:CaK
2N(c2&_V-0TKg3]C5X>/,.#7NQ2,f)P<;E&aLW]<+K9,VeL)SG6PLQT<F2D\_=OL
@A?ESUVE[8>VPKMT@CG(^&7LIDMf[MNR@ZRO,=A.AEX(S<fH3YN:,b7V639U5??0
O+6[J;P/G+FB^9(8Q;1^cX@WIC.e_CeaRPPXX@M/<M-,@S:+V]NQJ[NN.-8?2K92
_7L<.D+^Y@[1?4DI4ZgDQXZ[fX_N_-GP7TX[fc(>]M0PZXN1\AAKZ<4Tf/\HO@(6
F.@Q^CFXS@&ZFfVb=PVc:=].HI8,Ge?71>[/6MLc5CXGSM7Ig/]<L8+e1CA_,WJ-
CdTeF0eT:=VRKZ]YZ9AO/a00b8Wc4F6:9WWQd019?53P..N<&5G#YKZ3?4^/]:SE
)c4EMM]7[d;U\R+I8L)TVX/GB0FJ+3<\_R&21Wc/F@R;Z@+UQ]GV6N>8_HOE]bG/
MKESPVgDB+V94)b+\V@6:\88Uee6^;f5MRg_2]5Z8M9<O<Y9Z5d1\ZHH-,C=JZ7+
VJ.=T[c7+:d;[L_&OP-DBfW[>@f8c9AG]gD=8^S03RRe_:\8<d&=3Za\EAKdBN<1
^1UFcDDQS+==6\\=I)V27;I+O8)WO+aI(&<R6deKMUS\NAH?/,:ANT?;g=9\:QF6
31aFTg;CJdB3Ye,I)[K.&C]2b&TX#Q&S/fKcTSf:@8&WGe-S4M51,E5.VE:>L6/U
Yd99fHLZQ6^\?W[Z#DIe#?+6[BF4M[505<P8Z[f3c:>6TDW^Y_BUB?3?J)5/GHZF
Y-#I3N@@,HPcQN7X#1.Ld9bQHg/4,ge9]4?2R,M_eMOa-&[T7F0LQ<//b)W0<?P,
CA-&M^4D)=(XDKZFI+]1NMU14D^C(f1X,:B#CFZfa+[L5V5662D6aSYLJ0f;/;;g
8NfL.QX)-d.(-bH\#IX.=0/<\DZ.b#fN5MMUEfP@96:Qa&2KJ;C1=aF[^a&K\\:X
,R)@MGM7J9S?c\9@,26:7TaE57V;SX<(DZA,dO;98JY@=\A]0NE_X)RNN_RV<^RV
^CTUea>bLP10^6GM:HA?aGF3TQD[V?DYYA#=>JTLJHNKMM?P-J4Z@;FT+7CN#-@[
U=1/(_3T-3DJQ1GJf#Eb#99:=M:;T&N+^L(ALdLV^e/NHI]?e2MM/g\c@,E8f+O#
OKJ0<8)#@bM?U:KV2^7GV0HV2@.-2KfQP8ZP7GFZ,-W[>ScT=84VCHf-])SEfYL^
1^X2K=\V.GC6MgJ3^6)H2^X1e.]#;_E_-MK9/\7(T)E,K9#/gS>98:GY=FOBV)>F
=3?7(>gQH1c;XaTWC^,N7gb_d@YYSV2g9b^9[C6Z>=8+#Q8RO&5SJ6[<ITc<(eHJ
Jb[V_<Ee:H1B5/\#O._TW<c+XWKY7)T2<_,7EURc\:7DV5S[cQ>;4;?2\X[Rc#RP
e[_(UX=+N<V5UQ0U.M+A-DCRG/;9(18L332T^.?I@&VRAQINYRQX1f4L=,P\]<1W
^[<\)&_8L+]eX.g>=-:ecfJD\Q@^\OD?e_6eDPZ]BWGf?W,;D.[+M)#(g<HVTD4:
&:GA(M/K_b/504JCRBZ253^SH8;b>-O6bY4-\(SAOH7+/e=-b4RcU<:3bPS]R7.C
PSS<AF3+>ZQ2N,])].XT+>e6?QDALRANeX]fFA+YU0-Q7.\=e2F7deGH.N1b,)91
>H#)WN?HO/dQ^MX#<MDSPD)#]A7[L3]_I/=55\FUEJT_4,&<[H:1,00VLb^F3MC;
?79).WFFX\7UHDL9EANXcPLfU4A#&]=Z9YN6I=LI+M;K10TC6TXe^5OQ[g@<ODgM
8SH-_0P>AWZc.3)gE7]E]1@&<PX_-,WA)5Tg\L<YgV?ZI&/P^YdOBKV8^AJYU8VL
8dG:V#e<<RX6KP,YY,^1fd:(g8fRgaZ\C5@YQ/F+[>XP.;6>12V6[,HeW+Y\Z;[C
a_6Pf=6]NGZ.1,T7+aB8.c)-_3;6a__Uf_Pe[;3@)F&2(X03;];fO87+[cG;eQ+^
VR2GId-c.Df:)ZN:I8;,8U^V=6]^YRO^d<a.[QfC^:@0G-IJH9e]9eSDHNRMS#Wd
.LM0b\YaTM,bY]Y3:8a:&3?eC(23#^7DT+NP&a/J>;c.0@a1FR;[Q??Q?&]S)[EP
A7M5H]?(LU,CN,J/Ld0@fGZ8eA,PKXaP&XSfDE,@>AFf<3Oc#R7/CN9W28IeOZ^3
X>I^(X(+K+K5]eD@F6=cf^WJ)CJJL8SP4@W_^[C4>?Z,b&[Y&XL1(K@SJZDKAR[e
;(+G:g(ag/8[O/De&YP&^TD2cg6cW:XM&W.dZA3OG.N?cAYH0-QKdGI.Ga/K/2T@
/a;PbbOM\8Y&EB)?P\1f;_(V.>F,WUH,37[TbU_J,LY/=90,<+H=?SPLcZO2^#UP
V\Z>gT]V0fC+.L<S;E)-Nd.@71\D>ddN(Z5U1HDbbC_V;eJ5IGQS[4Sf3,\XYB3)
TacAL)F:<IGc)Z7=-W,86UI]U,M7D8:#_KDbBaU,_59^WG6Jg3Bf(B^7XHUG5H[6
c2,=XICeWMc2[=cL#H[Mg37YEZ&2/F@ZB3gc_ES0DGT]BEa5>FT9PBdYM:4e)DV9
NA6(>>SVaZGYCE]<bA[#/ZTF^bC#L)&3HCYVP2V4>7&DHd@c55F6\_142Z>.W:^?
EKB:8@+RbCK4=&<5IT8V_,]AADaOZ;R4<dI_bI7Y;9O#?@];Y/Lg)+6W10)Wd8TE
5@C^S5d=cYY&fYXM(OX#ANRd1/@GUNO\0Mg@cg-4[_fcU\b&FMHeNaGMVF4RSeW_
H_aKJGDO-\9&3f:#L.geQ8^/&ccVB>2JCAT^ae#&=.gcB]=4T0Y?6@O[XS;/1VNV
#7-^@]a&[[.C>2.c._FgDNM9VLHFOXQg(7eK[eZ^YPP<8]DADFV;?_CV+B19f<18
,Z@JSQ7Wbgbc=+AF_MGRY&NNRYHAZcED3[>TZd9N@:]>R+L>YCG5[EgMZC.Q,2F?
Rc?(f@V0;c0,>W-P4Z9]O2KX>;c/W&<C/S/EG>C;W#/@c38>FcN/4f5@37M0TCH<
9_^cPa.6@]f<.+QS9Lab+dE4;2eJSN_O;ER74N]aW+1MGV#DZ@K(HcKYQ)@Zc\FW
2@dXCW72B^a1J+b2+<\Q[dC^2(R-+EbS(A9F(L_GZR/BHBa149NQH8V#.#B@[GD>
SQgYK0:FSeMd6]/XS)5#_fdZ@KOf7J&Af.FB?^HeHJFQQ+GV;6Z1Te4Wg(?PBe-f
ZEMCf3&A=,/06][/e:[Kd;?cEO2Q,6QAPJ.SNTSZ2L]@,]d@1=<AD;NUH=BY^.eU
J85_X1d>]de)d-&.-OQ:&.2X\_)0R9FJGX]F+N\g^B>&-Jf:P>/4bT]I9J/,&V;=
^9XO,8^[f4G;dgG3Y@a_RK2U#C>V/6HMK_3aH0dB(.HTT7Q_63c)Hc9EG#KaUf82
2^<4fT91>_<,V<cV_U)\NaU;0X5IIdQL40(67C3#Ddb?P+ZKACWbdQgfXX5cY2.5
LK8@-#AHNWdZ1RaO,ULDW4YA^0eCR\AA?_M\<TAE2RgNf85S)N6UW:.:S-IT7Y5b
(?FdKN?7dRU8L,?A>\cJ6#;A7)8J;VZJ;R1)1_,0@EHJG,4QLabG3N5.8,&+4G5B
=B4+]gbH5+_4.ceCU=0Id1f1@\-eXb@SN/^)I?UO)PY@7MQ8,.?3W(CN2\#T8bNK
B[;@;=Q@MYRa],5)T7@cG=6FTe^ZUU(.6\&ZO8fO,3,(T3G4C,+fadB[CR\=96W/
J\=RJCTX[?0HUeY^POeH:;4+4>:?]74Q0SP#3ce.SSBe/Rc)c&I8fFSAYCe.<bVQ
-eC=WHS(af/f/N)gHG-&VMMUD7MGC7,8IJ=NKL\=_Od6H0G[L:;93Ne59MDR0W,[
(D@LWTJE1.1Z&MAe&0[]aYA9J9g&e#+,#=bMf.RUdS7/G?(ObIQTg<42DdSB6)Ic
JOcV9,?K.2M3CQUOJC><,)9H;8Y..aHF__IXGZ8@\&_,T>Ce/NK#K\@DVLVERPRJ
fYO[)<bc@=FY:G(/7eNYL/aLL6T9YHZA1AP7,]=I_Qb47?-OSZdCX9:Hb?U,\Tc-
.M6^deZf-9CS4KS#N<GS6B^_=UTcYG3B3Zadc?Vb&8?U3(<&C4XME=E&BN1^&-[5
1bg>GVcPRgKV=K)QNESdTB,#(2WOP=(=--+aR0A#DR0Y._/T(YUfgWNE\OF,X[67
EdQ;UOZ/C@/APdC#fdG[YA(IBKDQ/5S0H-L\KBTPR\4,\,V@8YKUC-XaL7g@V9f_
KW6)5;<E)[Lg:36>YZbTe/>X:AdP;A;5;N^C5]W2Rc2RRKX:84g3#^/GSPI+XF7^
6P#&T+M&4eCS/5MaBNICXX-_?_FTUQ20P+1-#>##D[2Q@WGdKd:<D^T>UT6<[OL_
]J_-bLg#Rfa8YPg<b>\X\C7O7WN6D1MGF00E[ZbMZaY2AIPEVLVKDYXP68c[S/_,
[V4b.2R123Lc,#^K+U;ZJ0]1\</,]NI.CKe)HS(JR1PBG1+cdef+EB(]NNeA&UXE
[S2MW<]OH,AJ-X25).Gddf95K/V4?.H.E<<::4(1P/,[CV._=0#XB]<?AIPgK/5\
C.C(:T/OM\bgeb0cd)&,fac&#b6.R1Y>;Wf.VC@=W2_AWXQQF-:#c#)&VSOTaK2D
RX5><Nb2FA;E:YA[Gf:)c2F#V#G.CEQJK<(E8SJQ398Z._/-G]+&W)c(65VG^Ne&
dLYQ<K#,ELA4B>X5[6S2\6.dL2R1c8@\Df^H,.7Se#[d4;BMO,NdXQ27ETbX;\PT
3VQU6B]#0>PT/4/eF.2U(&&[&\d-^Z@JN\>@eYTXVg(I9HfBV1NU>2SOEE6e,b=L
TX/(:GE7F[KK4=0T@0adAgVdLAc6BM3>H7-]K+dY66D46>O>,OPM,XXP/[H(9&7a
MQ_L]:FU\DMPLPbHT-CJbP[ge^RF>L+UQ0(0b4G@?1ZX=J>XGM+aSe@7[\BPD5<-
R4H4^df1-cQO73ccJQ6;H3WJ+47N#6Ya;U<2V#^R1V41cXVUE&QWEcU?M/5:/I4=
?&[eEgbL(B8563&#UNA]HdgRK&f5Re+#ecVTSM+PAX4H2fOHV7,UQ8<.WgY1Q6BP
)::C\?7(FOK6RJ@1ea7L+c4PSNKAS?B:P(]/WRRdV=TA;FCX<V^L-7V(NLe+1\<\
WQgT/_deUL8O<;;081Y+5Kf;Mg^B4#-ESf:O92Y<Z8e[P,LQQ8]75DS&?S_8DDS@
O#^gf^J7C(M[8[AV9#?SN5]0HBXG-Bg</Y6a:P10BbY7]]e>7I&]=cRG;W+<<>9)
XbIRPNcc8T0dL,MMFM9JHF2G=62>OMX3T:?M1OT4bSR+>]Q:@_9d1CP3a93:(:PH
8f^#1]DbKeGBWed;N)eJbOVJG(_/AO;_#ID,ZTZ4a-WA;L)AHTe3d>T4DC8_UUGO
Hg;J?SM/Oeb2S<GTIN_F;ZH)18Q]<:29)PC^IK)b=eeTDT2f1;=W)NdT1?YUH1b>
S2NZfEg3_(WBT,X0/S^QZ[FX<>bI8&?_7bfP\D:,S<N&Xf#@1@fD504WQVK(/.=>
3Z2+8:=]W#KQ(=^?[9?):7W&B6LfgePN,ELU\LaG>d#&E80a:6cCTR@b>&?0N)?&
b6WCLJCXI9L.B\c_E26Y)&;YS+Ae^A8U^;5K9=M4APgbc5CC?H)3B_U.A?aBF547
0bMY)dfQC&OcRKTEd/dHSG=_c7)92ed=_-0L)R0>\eI[/29(516;07:\./(D=-Ec
M4[(]YOP]b[[1_TICD,SIE1fVa6aTO(O+eQPW\dX4e6O0<E]_M_@6d4RQ7a7=,0.
0NY9.Q0?aB[V1&D@>eLdMO9dNNb#,JPP(,]I4>.@7O33\Zc@g4W0<<3Q3GZ0)_->
,9F?Gd.F&e0b+cO^SD,ZC_>+X\ZC#Sc8Y>6>L5;^Rc/YS(+YH2FD=&9;?)c,W<>7
IY\.a)EA&0^>N)3:W34g:#P0?;a(ffecI1-YR4AIXEI@4>,]2ZJ.RJ[T@(,[\Ng8
2f-ULBL<@ScFO3>]9<&><B/KHGPf;+X^3-=@RAU^RSc1_]bcR3eGaf1N.L4^e87T
J<,VM^-5@]gX&.M[OF6GLA>^P?eaV9WKE3Z0J1P2[;gIZ,<7<-.<#dH#Mf(#@4OF
d^1,ZG9c;Y7<W+)gZ-FR6EX<3CJ<0cbf]?B=5))S3H0QSWV<0@U/^U+/NJ^<T\_5
[dHULd&WC&7g?aW7MC;e4OYgYQNAd>[IA8T6+>L^@M&YQd#6H.&cN1XIP<e.W8bD
M6IO5IH+_1NIZe[63D_VXgXPH@H<Y?:5Z?>W0L9TP#2c)4ZJYE\A;=Y/b\K(\9C<
BRC1&6fg3ZD4W[7GBB?HGU2BUWcA-_KaDaSP_<Ad;.LK9GSG8IP)[W\U_JY)0Y>8
[7+B0JZ)=GWFOZ_DOZ]#P#O5>M79^QDFCb-e]8OfRIRN:H?J-dUE#A4a+]4\4B)@
&).PDUA?2R94GZ16:INb_M=S_PD\;Q832#JF7PZB<M]ASDgW-_REGM8>[GW::L>/
]0Vd-L#&?SAM:I/gdGS,aC@61CB3P1=bF&Q<,)57O1_Z_dRQ;):\WQNGY.2:FP.b
BJ).T,\YE^[&T16_9Y+K/[9\caU@C[YFH^g?<<f7C)HITNZ-?X3KM-cfg6.5I_RW
cGW.BW/A[G^U(fM##.I-+>Q&)+:6^IO_6e&W#I\a?,+Z4>>^VK<3LC7X8BV?3\L=
VbV-JDD&4G[7^[RK3B446WD4CK8b3[\7fD;]ZVI2PQGC=e=D3N?\T#A)##EgIf&A
).ZfgM5-5.VRH52Z</d;\YV)C)3J3=MFW84<C\I7WTV+Rc5FOXSKf(>-/A0,8dVA
7+=8DBNH_Q[JZJc#g+H\cRT6=WZG,[7=+=JP,Q=24Z<5(W?aJ6BWN+X2c&ab#fcZ
GS/H,/XH/V-C).eb#EJRd77_&LL<1=Jc(3E[RfV4]]Lc1-E0gMAZ\I52@.>^28G8
[:W822&2]OXYLBB:N\WJ0JF,2Y5V:28RYQ>_Y<YCU=@;4H?\+;90ROXWC+6UHEIb
;I-_H7VLN[9g^#6HCXH9.c0._c,9,LYC/.I+/HJ[N++X2b4f(LKD5NGVV^[]C\V9
cEF_^N2BM6,DX4GbgI7WC]GT&W6PKI3L-HUG8]L45/eE))DY>LX[@^G2=EKLO2\A
H]7CMJ0ef^039]4@.KSgSSP?M7]EZ:dN6-g^S8?&7A1g[MDT:.R2<3UY.O>T.AaB
+V<?K-17TX#M5)?EY[\B:DVNP0=G\O4EE.3IA.8Y0N=/=[e2QI,;\cb&@_FDYaUE
:4fXeRJc/7/-aKH7X4])US<gL06GJY0;-ceT550<?VO_VHMN8.):2M>7?DG<eC61
fET6TJ>,=3_@YN<48?.F7TgUW[ZX7J[FQaI3E8C@B+fYLYR+LaN-ZgO[edJVG+ZB
OC9KP4c@fKA&P(@Uc.@YVd-]2gTf9G]_L80])5A5\HZ[OgA=W/@0D(+D<,F^PBdZ
E5XJJ7CQZTF/+c&C?FI9\:0&H//OO6L\,.0W)Bd0)c:Q/+0;<Z]VG(fbaG(><aBC
0BCB;2OD0E)Z<9Kf.4^INb4+\R=IdbFA.R>HLO_V^TI&(@QL<Z5A2[#QSSIVY9Ca
58QK=1#(JDMEbHgN=(-HE2dIDb^./_#VEZK8Pc>;abV=44]A6X@eX>O3J+2UfM-H
3HJ;\[>SfbFAVJF)2#JGH:]37PETe-GZ\a1K3MH;KY16A2Q:@[>f7P[?ZU#aa0MB
6YSY?,F,W>a\]YJ=??KH@QEK0)ce85W7I._UL97]Q?WL1d=C/_cVHR<GbM_KOR1=
BHeQ1;?<:,FEYRFdXeU89:R3>gebE=C[PHe)@)RdUB[6K0[f,,c?U7U9<:c@,bT@
XI]dBG52e/,:c+]WEP0U)MXB-Ld9d-[RI5\7J0#DX:IO\PGDaI&,.<2\g;FfX8\;
#fc;&+SRTN+f]6\DVJPc\]-B?;,]@,Y;__=,GXAeWBb]4HRS2M:WP)IXD-(&MV/d
aLWVO+DPL0H3=7K[)eOTa5RV]S;1_PSH1W2H37J6,Le^&?99?;\W@M:U,;N&+V:E
#E,N^dRZX++#THXN:TB/9RV>]a=]UM?;+MHV0bO7O^daFOMNXAUYE824.UTWN6P7
6#BF<K=e,fWNb:II0OIYN4UVFbWJc89<V6H)3OL.gN1@=#]]C-:N^TcZ))UHKHeR
#FdCGD\KXGga?MDW-ZO:95QLK)IZOFZ);;#906,K(/E62U.JI.:9\2@)AVd(.Y@?
D:/Y?8[cJMa(CAPTU;/)F/=W3c;<5fg7D25K>\BJ3fE)9G57?aI:[7JGXWW77_=V
YY2ZJSM[=C7=Ke^D(,N.6G4LDE(?9CG^S2;@V7RH@_]>5?G.b3H@MX7<U_8SQ6-X
/IPXe4LP:QZ<U2T\-0;_.C-XU(2:L(LY<[gP\9,0[#,+2C(G=e\c?IN<)(9,S\]]
?S47X/P#J-g+7(-7@,2N:ON.[B6W<.cUNX[Z\<eU=d-(?8D=?R+gcH]YN@,:L@?6
RXM:d)MY-DM-HAN6RWZKC@353IA#Q[KUKaPWI>_aC^789)NPVRB;X;5]dXXE+;XE
/JDIF=((agW;[?6SMCPYM&^=5UE0a+0Bf-.N[,Z/M/D@KF+5eC16Ib.)K6V2]1AL
^T0fUWaHNE1:^4:VGAH>).UZDdDSeNFMK1H+3EgY8=L_a9/2__6e728UeEQT=A@_
cRa<D_]MCBULC&25&?C,E8V40<)O69@UA^eUO&V?\+23/Z:,Bc:fC]@WI(ACGe7C
\?#VUH=Df4@a-d[U6)VI<0#;dfDZ5d==N^bKM-QS9e03fZd9-8W#-0d[OY7@I=8F
Hc^^#[ce+1?O0K(88a;]@MBQ_TR=e:+VO67K/4Dc>:>B:::9.Y8TcD_^NK<aZ=fY
3O;4N#8cL/J]G]Le?c431K)Jg4@2W;3Wb&VY^,KD^5HZcYL-f9K0CR,U+09ZN/Y:
OTe>^,0E;<)S3>(G8I2OeM40Ka^BR9^V;+9]C]+2>W?O8OJSW@+7a5>Ag&<C,f.M
D&(71S-OD&CHcWXR?;dR:7B6@U>ca3-]DBQ86GEAJ7?5J9g09U[EDP-:T:KPg_\N
MC;PK0;H##:[T6R@4M4e76,@KK>N4Sb\R]VgQe;7XMHQ^(8I_PI&NV@POPLR8:ed
@-:68J5ME9.W66GPM-5MC(QTNS0eB)dgT/Y=E<3V_<LSg.1AM69GD1bEOe_S?RVS
FX]9_BZEPGA8JZ^GU]?7D94L2-6=PU&^UDG,Re7Y9EfV19I?Z:R-9RY2]T)9.W&E
9[bVF)0gacQYDI^ZT]\#FF/7>UcP?F&\HW_84f&G3#^07/bX;?&H&>.FFQCV+UH5
^gV@A[CT57I+&^F+Q;8gK0V5)@3fT5E)Vf\WVgMA)Xcff-/Z5-c(FV+WGVTRDAWe
VMYIGKI<DJ3/Y3BWaaL=Df)<2,cG777LWGFRE6dGY8P,02]WMK;b?DBU\8U2?A()
2cLA@7R(/gY)XRB7MIJHT)efcF18EGM#<)#IN+BO0c(3)aIPHf2LMQ-3UD-DB\I9
I5fUL,[f5V.P@B71E/O0dg:K48(RFU/>LZ6[\UOc/U;8[3.Y?2)]dH16X-:3RUZd
+>@=Y0:8()S?\f-#gL]IZSXTS#f:g)U[I1IB=7fDHF&?QHMDWe-cWX;ZbJ2#?M70
(F4E38a<?:;aQI)([9@>XFW3OSPY[,6(7;,-VH^^VH#A=c+5K#3\c]D0eG#A?+eg
\FP2(9=6<MGK0g=ZV<IMMd48L)c,fUW)aRbaFJGQ\GL-OfP8D-Q2Ec+.6NRFQfIM
E8PYS;0c]+0XSC7Tb8cHE=QAT,a<c+XQ^4c=:HQYTIM3:+f2c_GCQ91DON<fIbCZ
:C#gYUCYQfM+5FGYG+WP73D#63T6H);Q/;d>>L)\e?@dWMU4b4\2e)HYUg1NS2Ya
Q2M:aRC3C<8f2&fTY4(c?g0dSRYJK,ff6]RA+R^5Z;M]).K933>L/\L=)]J:fCO2
EUQ@\,FZM@Y(>TJf\C:#-d7EVB:)R?[HL/QG3SQaLY.>fM0NAcWB6<DU[D:?]/-F
=4?SO=CAY_5b&:Rg9S0VXH)C;U/FB5VgAeS+WI7P6B6K#3UY_76BZf7K4MAPdU:1
](-a-gUfYAW;Q;/-U=3#H1Y^ZF>1L@O>J8Vg8R7_D\Wg2.8-?^MCEeT?D\+1;AX(
+^??J>#7<KU&@I[a\K5(7KRf7M)5Y^?A[->UN2:V+=1K5F/R4E/:ZLN(4cgJ;_U.
.5\,X/0ON,=_)2[L/GC,2gR3aV&3\7<E^.&b;-9G&ffYTJZ#&]GQ)=\B>e:G]/P-
+TY:d54N\PQOQRfE[CG,W_(^,cXC_a;^U2))QST/HQcBMZ#Z&P80QQ(^.2=<.\)c
/&dHSaO7e8G\L:N8A&][cI75\S])c^=d2/H>5L:B0\R8T@b)/LBW@7cZ9a(5#8[\
g+4]S^b;>DRMP4JMf_NgTJB/ZBF/YM:&T[@2.AUD^^;C<_#7dR:_;<S#e^)M;9F[
=a8QHb2=M(A:;ga<N:Ic5TI+:(1A(I4+gF-H8P8E/5AZ.8T#9dGI/LNCgO4+AaKL
_d;NdWcSb;Gg^/+N>QXbdVUA9(I&0#42f8YKRFPeJIWO\@YB)8:/b^6)TIP-C7aI
0B)R/;.f-SE_gO#,fVbB@ERHG,Fg^?#,&9[fPgQGES0LY7^TM/;\a[/5ZH_=,XOD
;V_#8/<FTE,N#;5E.\.b[P:;+f=XaIA;BJKBTMdQ=RN\CUD1^6T-I2T:^AURW4BW
M@eK9=P35D>R&1KFfOHZ[f:QR0dD1E-XVa_PFJDK6M)W?#M7aV\CP@6]XA(N/UDZ
^PZ1d/f^EV;2+DN)-;>J8D>;=S14-<+)0V1N2-L<?_SgU+LbS73a<_d?JIMXQeUJ
7;>WIZd;=FZ(HYgcb-RW9?E=.T?c=e74KB<?\G8B;gY_K8U\LGRNPNQ@b)/K<dZ.
:3GMZg)bQ2-aA9U-G4F@),VI57UBW11QE?K25O9,>.M@5?D]_\8Sf>^+LY0eG/O,
LRQGE6.06N2gP0O>Q9L[GY?<ZWI47L@,+]P:J1,/3aGC6+H32ABE3?+367#Z_VgJ
@&I>VLgS[Q,O\3R>JLLfg8,>E;W0[FK.[GYQ,9LP&+FU2?BP\+<G+#Adbc@&+M.]
e[=GJ3g=@=BgDG[@6cQ=b;K2]XC0P21>.JQST]AI[1cTTdT?=5[IbOZ)eFSL.If]
8E1QG;<N@+C217d8[XJ9MHeZ87;KDHIg:b[X0K2g[^2(/FfV^:#_ABY&OZ^>c1#J
+N#Y0NA7V]WEB;:=UZVC#G1d6=ANfe#/&8g&A8-V.),U4O74X.DS(B1Y)-XU=E_,
+\JCQGBVOf\\WUW;_M/<T=JIU66XA-)Kf+M6b3+IEZ9T&#;>H_,e<L:aSNQYU,gS
#VgU\=SXN]&0Bc,Bg2EC]/@-O@=+MSU\MNIf;.H9IVe\QM07Ya,]^c]b>gF,fLN&
QQE-7+:[NWeI4A2?Kc^&+(G1Lg4EKL;Y87)RAV_f#\_5?9(&(4Y.U70Z4;WX(4I<
TI<F7O05+RIKK5fT^4WVTM147@^KfUHf^DWEBAICLIAd.dP8_<b7XWf\B]Y.SA1f
H)4U)/0U4e[S^U<L0L-3FY\L?c\0/9:?AC3>&c,&_D.DCdES]S3QFHMed6NMG#3T
X.6VIP&^\XeP0WfGaLY#N7,a/;<@]R11QN#7#-1H)DKK3VXWYdVbH9&O4ZMf+S#B
5Q#1=I:7@=DS(3[fBGc3gee)\;)0IFA[,ge,?XS&c(f?K[J+cf+Ya7D&XJEJ^@a5
)()YdU_[XWQM5P8,=Z9.S80/.^cUf;I-HC+E<I9#DP^<R)AP;&^9LQ_B3[JY@\.)
WgCKPIIaf>;G;(FZd[U8^R:<Dc1BM7aDTaX.Ua7UUCDf@:\FGK:+O3+_Uc#C(IWW
)\;L^GfN1&6=<PU9K>X9+3=DE6_KH_Na43=09IVZ=GO36;E?G,2fSYBKPG90LN_X
&YfUF8b-TGGS[@(C[V7&g2)C)C<R<>ZegN#TKaR[Qa2N[]EX9V;aG[=N5C7A&Gb/
1QKH<gW@,@X/=01??0,&/Bgdb4B:&@;-C@=SKVG>#@eP,H#MJWAgRDF_]HVJFZ&@
.HegAP++V1Ha+:&QI[2C2Q)-BTOLZ]L2A,XG7YVX[^[2f>\b4Qg+aU;c4EAeXM_Q
@c,39)ERb\XSDNEN5aHILYV1013[4#,\7YHOdDfL3^^-B1I#,XKI07Y[BVZ0Q3/e
dL+#W:=,d=&M07@Md_deK80B:)9cR>]>0IM.(H>/=/?>Y,,7VE.1CSKV:_KH#/>g
gFWCJ7A>3f9.:1W6Q0/:gG:EYV1Oa)UQQV:FIE#JU0NW\(KI,aF\KENT(]:R&1,R
:=ETI&VI-(g(4D3Z+-fEJeH(TBL-\;Yb_&12C<_Nc__@15W\VT/KLP;@Ve@RI6,.
GKR58G2[Qg?#f;L^df(faKH9Y&/A9)1HS9c[Y1B67-_((YJED1YacAbRXH\N\)U(
ZZMJ?Q:f)6c#KSHUG<9d=809P9X,\[=QSLG&-7J6C++CPSfI,CBVT1KEb\f1a-QB
Q1>@@U>RT(M<be^H)fQZIY0(+_>7:6W@6Z8BGV+A&5FQN?Ag/#J5SY>51Gf:_](N
C&-HG&d:-UY?QK0DeKB2-0GJa3)(L:SGb1A@02#.X856-8#PNPGeBOVAe\(VZJX^
,=C\0dG^G?4L6#,1?ZX#S#C>)C^<5f1^+bA=?1eK=GU&_\YM;,AYNS/J:QdHE#;[
?;Zf9->Q/3CeLUbdCa#TFV9JA(9ZX,ddgXN[;\d(F9\fL\^4Y98ED;1(^8@(:>d;
cfW-=Nf?e?U0PL4P6<@_.UK?>S2]EV]MSND]5(]KGgJQN.:d-4EXDJ)8CBVa690b
CL-8.-G3KYEIg[A_.K[+dSTW(g39IW5aYED5HBA]?,6O1gMK15]52ELHYb7@E)D1
K:<8ZO4Y@c0].B:K4>LR>e5TD^Z?e]eVZXFMD#O2ZfL]V+PR@Ua-(_4\_L_=MH?&
OW0,X;<0bHE]XC0F9TR(d)WSIKZUQWU_JE_HZ3^5d0Uf8E[YB3M1L8P+ZgdLBdc,
e#dH(EgLX27bS6II54DD=f,,GD2NBK]]3,RH1)WW_BF1.OA=7N&e_;IJ1Q.9]OGa
:IH7(7fJ=BN6>NBQV/T94]59KE0LQL[LHe<2)D)@IU^Wa-A.O_?9H\6PL#QI.9CB
GX^]F#f97b)eIWG_aHX_9F9dS@VZZ@T1#Sb(;g2M-@0#CWJ+-Vb^V5f01#=5/]NC
PXBS)J&,N-^Z)I)^#W(.FJ>#9E][+P)YGYX:X^AfMA)BYST;GE\U/PYINcKT+7Z;
B9Tg\60>;G)JIHGJBA[\>/VB@Wf22E+1OSEHVX0CUL0QK,9=#^@5A],Kf3@(OXN/
)6@4ELfJBeMMV.c/9DO.XL#),Wa9[c5J+.R^9@?K6&^+U(<^gEd3-.Y&/O/A0d4W
3;TfCY3]NT\Ha]M)Q.H18POWGS;dg&G&+9?V8,,0&C<IXI(?V+1:^d-bNJDCHW<8
CUM,H;D5-<?M)^\Ob1)d.[C<LLY,--g)74&&E7DFH<daUS5H@XMcaUS3cE,b8b@7
LH_3-D_(8BT\L/9If555=^FC4=#B9LRcL;X&1UX6CJ&J6?d+S&BMHUWZ=RK^fA^2
S];E#AO6T;KQ+[58cF.VZBTU,&+TLgS\F-:735KQ1GXH+P-20[<V2U3B+UE#;#NP
aB-a>YO61d[&9b4KHeg^gKgKGH\-63C2;+J<70OR?1S2Yf07[Mb,@(BCKMFD_BLd
282cHN<V4S@F;8Y\R1:UC[7W-UZ00gR79R?^O1W=d]\13XW^^b:94e3A4+SHK(+7
:[Mc<.11eA(#a_aA&\<>]4ZU^0)Y7T\7>8NSJX8;dTH8)E(gO7Y:V-?Y:LYMUQ+4
B4SGBLcSK7G2E63T8SI82@V=3.fT,+GN4b]DNe+BSW4@ZKIb\VD\ae8GDIG:NKYb
X]a_^+><3O;H(6\0X.R@JO5;>(:5VF2[-XS=R>=I,^c(QSTL4,U@I6gFL8:FY:@f
LL&J54YI=5:7BHGV7:N.#+KA9(Kee5ZHOJMd7=YKP5g?gdeLF5eT3,C<U&=\K7[H
-,1eCV,P;#.R@2_R->_AP.,02dZF>+(=(<KKGF.K)c#M(?b_b.Vc\>KG,;WbDR&U
1_@32N:c5JMf0YH\^^M(J>.N48G)SJOD<35\(87I0]Qe3=Q#:HP2f&VNK=(LDP7G
Z7gISW.F@LCA5J\1UKa<+]30@^-7ZXJT+DI=E=D+KBIMC/C/JA\VS=GaU=/&/7+#
OX@&ARQYB9^-:-F6bL5gT.C_fMI;2,[O628,0Z@fYc_agP7@eCgb9D&YX:UfN\9-
,>9^+OBHR3a33C=:@aXH;H_<.VS)HNJ]&OFU_/U&)TRg3#@eKBNATg1;;>CIc507
2]QN</#NMOBDfcXT[Y0_d(fGXPe@gS/a8E6IUQ&IPQ>A=C0-E\1XJS_T]YG&W>e:
N0H=gH1N:#?F:+Ng0VW\9U+74=#F;+40&32AW:)D3a;W5+Uf=.TN]:BP.\SG1M@;
&IEW#LcGZ<]&KHSY\<P+dL0J#RNdAaHWUP5Yaa(E^RVH/8?3-1b/I^2CW@DfK.QF
K6d3HC&M@G:B8#ZYR(CBL3?=8EKYa5@:Y9])VB=4C3/@:S9[^D1N<S\?1bM6/@.Y
7G7].#A#ZeZaXCgD06/1EbFFLcQJGgL,G^@EB2d<Y>VfG#>b1-6X/&B(PLUFOOD:
&4[_c]1)Q633DVf+A20GIf=>U,[#]K<C;^K/Y_Kg-]9TgDO6<->S3fYfO[D,.?4a
WFf#FUAWENE4N_2V,-ZHMU\M-,UCB+8A]b1:I<Eg,e3&(542-<M.KS^cF3bC9f#^
Wb)EAUbdW7DXZ:P:?(SP6O9LagPT2N[gSG7PO3<0_.F96RJe;+Oc]DP4fYZ8LO.V
CTH>RK,ZGdDA#N#Fe^g#\J&6+JZ2JXLJCE8c\0I\U\e_][R3TZ9WcZG6?PH<_,O1
W7[Q>gf4P.>f(:.W>F=.g6AJQO8d4ddI)BFDaVR)<Vd_<+V(V,4(VY\H^NXbPGL/
?R[#cEZ52_GAXgFaBS0^K\FE;L>90PaW+)+A2C5=S6?N)OH-4eU@&LdN[Lg0Of.8
K-WN1(SLd;;:dT:\KFe@QO]7A0DRC24<\.13QC(=3DJW0\2D?J+\FHa9O6>ZM,fI
T\cM3/+VFC.d(=+b.^OIcT#FMK,7TI4dcFN.RL(WGR6_T)L5KPdA@#L&8=[OPg2>
V9YDA_Od>c^QgV.CabA\,,J+8BB:\1c?\7).JM@<1eaL\b\ZP5Y:GZT4)_F+UIP>
OT1I+dU6KT9bTcK+_I>+_)1DEEI9EDeNAB+)K@X]bB8:^\?.?A\9:]9\02C=4M9I
19R8AIM+Ca-@1932L,A6WYSA?B,.J59M/&X8@9AU&OSXX;^4,8fPN?B1,&?&f&(W
HeGPg>ZL[IS38+WMG^C?;VC6@9facgcK^.fDNC(2P68NVECSMSfR52@T#;K&TDXT
:F,YO<\V&A[SQWQ4.GOHeK70@GK+/1VQTO/K.HA^;7?a(,X8g0M,/M^Z5G6g>#1Y
C^MUHTP;JBgJGc3^XN+bXX<E9:>3P988&#C>0I1L?\NTB8M0(B[fg-TQ0II]NGdZ
D^2<Cd\15ZfM4A6J)V[gYU.GE_T+PJ4Cag,OXOIaZ[D4c-NN9L:ORE9/#&S(QeE0
I3P)0RR+8d>)-Re?J+(7gE6NJe(0WY1JXf3>:9GMAGR-H?1J2;3?&@E8Z998e#K[
7IBE[QKH^XbAVNTK_Y2S78^AC)&#Me+gfDTaBI7b<9WWZ8.G=T(3Fd1I80;\:^5#
<I4C3EPe62eG#QY2Qc<.01=1;BfBgFd(LKg5@X4ROSL[SXgBWb;.JS9FW&;8>=d>
XZ:9<0.T#-+<b(9]CK4dRJH0a1=N#+N-M^ZCgPg8K;RL;_K1;+\Ta=aa9,FUTCF2
gR6-@YP7D);VC4O1ZaK.Ye^#VX.(\)d17]Ga)^U]MQZ03]+D\-^VW1W6/cJ&[XCf
BeLH6?H@e#Ug581_W/3KCS:=;K<4b=9:/61W2+N8L/.fO4eA\7BgcT\I\1.<WcD,
HFNFZC5A.X9JdHe..8?0_I&X/-JH&^)Df3KX1c>gc)g;c:W,;O1SGBS0fb7AFGd1
8P>,=VHd(gc&Qc,B((=QRG?V.DK(.JG73:885eFVgaHQJHa#]C@A+fbZgac06IT;
G0Lcb)+]OZ;#e3c&H]V\b2O9KY56A4J[cH9,(ZcC4YJL]1DbQ6c4>7#Y_I@Dg[PH
X)=e3ZAeGW?JPGV2,g37HI+aY<+R)N\fTN1(YPU(Adc#+6UW>GKa&17^+ab-@T?9
?84YdPQ^[RN&,R8PCD,dSHZD)Sb]=WZ:5U0I6J/c9O]_eTc=F);a@.b/OR)M7NSE
DODD?WeGVO_7CDNNSC3@7gRY2>_?0N4e2[W,INH\+DE@)\TLVU@8DC7(K:X8\GL&
]L9=fXV+WP([986Y)PK)2[KdQ8T8,)^dL?ZY]H)W3WJ@?-cbD[HgGbV?/@PU&eQa
WTV5(.+bWWQG\:B6^ZeRWG=&>RKDJMf2W/JPU\;HO_D3Q)5P_7c=6W2GU\>eXb&Z
f>Y>TJLH;74?g>.=/(AdcW(N^HYXC2;(R6>.SL8(9KN#-0(KecVbI[-2+81.#GV@
OA@gO(I0P.6Fb<QIeD&C;7/]C&Vd[MMa4,01ab)/W31f5Ic)JKO3FDQR@81YUQ0H
6^(V1KV?)\GYX,A-e@;MFHIYEg6W@,0&<LC4],PG)3]Z=5a<E]^>fHgE9fLU8PC9
+=;(D&FC<R;C.7M,C+=CZ>0NdTB=./VO:U,H0IP,(A>K:CDCED4(IJ089U/]4N(1
0R_]C)LOG9X:dGbL[K?DML(Y&>9;K9>K1O&IX11Z<5-HbbD_J#c<M^<&+R/dc91S
L9R3PS:B&L>W;VF&98ES0aQb+JZX-<g/+2\7/5<f)E36Y52^3_W+WK[YX5-0BR#b
P>EX6)?R>H:,ENb7g&@W87?374;4YBFE#7D14g=4SJ72,Ke\eNG=OK3I>([E,E9a
EG32XM[TG4&3+d2J@F0K0Lf4@JP\-JEM>0J+A4E>(8KUUWZ8F8f35_:AE79,aYgM
\?XZ5AUSCINXF4[6d8ML\W/+=\b#4d5BG+1?.EF@b(?VbE58U8>dc.(Z(V<bQ^.R
?g_?96,BKM4eLYPTaA7X1LS5[LW-4FB[aQ_2\CTNRT>H;RW?a0d&dZ<c>#YY@GDf
=)^e>:2e64T,\USQM:Fa7#4SPCgIXLL\H2@MS7#M,XSQ8K&01<_&=&Nc&>d.V@ST
+Q2]>I,XMK,W>]K&\0?1b,WH>#S7?O2FQ3SL_:-\,&P]D4PO[8R<=-4M20]I6[@2
[-&\/1LMW^UI>fNTD_QDg&fF]C_gc^g/6ZKR;2EUSR0e7PN-V2R45-eCQd.Q>:YM
d]O;LF.O-08IJe<TM@ge\/A9;6;^L/f,aN>O[/\Dg3]Ne;aUb[(_eE@(S]C]I\2[
VB.FN=_g:42J+GZ\H#e_B3WH<&eF]JYC_(0BH^8a3_7M2=&]>J=B.(c8P<1G25RA
cKQ01ce+J2/\^-U)7O\XFC]?:R\B-,QT>-[Q:;W,(WVW0dfdA[FY4NI<HK3RCL)M
C1Ed-9C=UZL],I2QdQ6dHR2eRf:X(1+aA[3e+O0+TRUK7c6>.B.WJe7:#6?b\?6?
9VA8\Wg4_3I.dUdYR[245:+.66[6FRID1-b+R(576SED_g+5#Z0&=<W[gP+D6)Ad
#=f+=AW&RUB<&>.O>C:IY&FaLF?b;AX#C?I=7Z++E7JU0>]B4NR_31ZEHVO=9@1)
9;0&]e_[e?>Y-FSQ3S4g>-,:=D9?b10X23d,)c\-Z+6aWTPf_-g/Bg/ab+MaO)FD
dRYI\?(ASd9@g<-a8cOX4AWUGC\6,[3KSH,;6G8e0_V5V9O9WPXI/_]EP\:_5M1g
1LL_QQO(@-J&KT]>\C_b&<[PW=>KMC)aB[Tf8TeP7NI?Be3_eX5C>\PUJ:d#cFF?
;RP@IgW7MN]J>+G?@UI&[[5K)]S-U6faRaJSQ=Y+T(-6VJHf+P)JB:]C).^=DCDb
R=F=AG:ODPbPKVK1_^N@aB6K1gc>9/N);4b9SB+8b8/]SZX4PDA;@^+2cdIZ/,GP
-,G/I\.W.GW63XOF/T)II_CC/A4HC,1O^;B(0MS-X<T06^b32V9[G.+cU\V6-b3/
Ye[cP0NA5;8H7_[_=/K@Q?DJRM8250#EBU);e&84+a]@(@d4<I?fAK7;PJ:f5V6>
-F_&2DG[>;WIFHaC=TI4Q/VC=BXBfI=]+f4#=FE;&R8_:=,M;4L-MQ,7WLG<dH5@
AUVeNeMM3ELZ6ed^B)cfW:fCN0T9aPRUGD9eB1b3cLV-MJ4fbRf+,85V)34.D)aG
@-N?Ic)RHI@fM]<A)bW@>KT/,/[&6;Z95IJa64bI]?/cg16Y_/>=>0/>G]3DH0U6
2QLP8f4T\T8P3+857G@HPK[M-VKO81?/T[-[GEB1SJXEDI)R>QCcQ>c-6[CXGHf[
<:)[<\-Y2XD_VKEWH5Lc8)?dB7ce79;DeJ^\W9c/(PN8X=GZOY?RJ.17]:,(XRC:
6J,OB:_WLbQ5bDT6d#XAQ1@&T#RZ73J+9TB(gD<>^<_g8g3;]8>C-0]BJLPYH1_5
-KSIb2(c,4g\4ORU0,U5JS-df42U[E#2HW0dBZ4)@L7QXP_4X,.AJN^O5MI6GL8+
>CbXM/D1IHZH]MZ[23c>A-=FP5TaD/2]U13ge8DbXASVDaL^fZ[eB>d>aTH[VWF?
aa1B<R3T).H&(;7V+BR1UJ6H0RU.gF#O,ZJ)dNfWeaT#U#\K_TSODFDJaeX#WWe6
2(MNMbM#.TPe\()B)16?;^.4B/S_:E5Ygff&V&1#?7?Kabf)Q@bCe8S;17:K6C<[
Y+>LdN[9GOMYP]^,SCAP;WE[9fLJ4Vd8W1_f4Ye:>]#\+KKcD#EJbK?;H2g0Jfe-
1gCNJ-f\_GCUEOM=6c,RHRbWR4E3?>(IcAU+IE#R\9>05Z8[GeVd7<17UaK,?4@#
DbBA>\Q@FXEE^DV>&<T<=O/)-9](PISS3C)Z.M8@dHc#b/L#B?]3.JSKbRfb1]:K
/a#>=Z<bIfbd];>;L-.\GMa(gG(C[J^;E3SG6#-//<,5P_&.K<CB)))+(>XG1DEg
X+G#,FIaF1&HF:=UH]P,P\.Nf_^B80-//@\8QJ:B\ZOKb\JO^gVJ+L)V]<S-SA./
M2L1_=SY6XVbQLEL\&KS.HT2&@:-e2;J@eT3W0/FfV-:1JbC6Mb>^80#0L]=V.cH
DK,@(_B+UN@Z?GAG-QVfb-XPD<6F6[CP[Y+KOLg;POUB(X#_>418][#:0dDfde91
-]9W0RH=3E4X<KKF<I2LKRbN#e;<cM5N<5@LYfK)T-Ygd@a//JB3Y-OeH/=K4@<@
)YVEMJLN0SSZMLMI4EB2O6=POZ21a]T\dE&=@=.UDG;G<E0f2X>;H>;#5.LNc\P@
Z7e4#V_e?B6LK9dd)V2cF3DHe)8>>cU6<dAK8EZeHKXPfN/?CYfEPT,8;@@B+29R
d-K;&6eK//H;K6@5L];J,ge[VP\ZJ3;NMUL:[B2XZ+df[SP[&FC/bFM-#-)EY30E
16WAb(gTBOGdU:(>YcQU0-g&YLC]Ie#T:#eH-fV>.M]/AXBE0A7dOa+G1c_J4L&6
P]-:4f#O[-^Kg();WgJ6@)Q.H[YKQ-0EJfUNaOVI@2=d(MMcO1XW&G13\=KF7QPF
Pa?0YPC5;8.,,_Z.10gLATg@ND8e5JdQYZHf+X;cPWXFdK_2YaQDCOMJX8<=-Q6:
a70C[S4?Z@e&TD;-?#4;Nf(\+-U?;W)T^DCg:6&K96TJb>5HZ8:1cB0(,DC4Q=LN
Jb>F/J5J8ccegE@P(2N6EH8+VE.U-+#9I;XZXSRBE]5bKDCNU2QE(9US21@#?OX-
_KX4Y]K=RNDA@fCc(4c-T]J5>0,dENHEY5PeRNKJ_QS8NDM2:1:QXU),9F,9BD++
82QMGd0>PC.e4,6aeTbC8IcTWVgE:8CN3NL_OJ=9/g^Q+,QRR@ZQ-M=ENU^0P2DZ
ae,Mgg\#U.fZL2AK?:;BY@Hf+FRg._/f9A36MS=QOYFTP378<PQXQ5f0TI8<0\bH
a<Z):/4SGK(FCLg2-&_)QG=d,>F+Na<P+[eK^7BP6>[:_)]J)96LS^1AK0.gO[OS
CA)>R/_Aa3(##T8=f9Je8P2TU:Q;[8;;^@H)@FRKLIc9@C6R/2[_ZbbWbH@YG2S4
7@[W<XOcJbcOMbfd6IKb(X/g@>efV2YTOf-c5W=<,Be=F]&C7XK-#((E.Df,7C<d
[W96O?LL+:I-NNE-DQe0^O/1Z#MF_?[&fgR+<A#4EDbb6gS8LGHL96UG#)0Z9cY?
fFUG4L9P@HeV)@dY6R5U+Hd5e9f/f,\>AdVMgI;Q[697HW?ZZfS?3^26_\-05?8T
?e7>1W^XaGG-1gMc0\TIV1I&4g(=5<<#?^AcQ[:,e==YY5@abWXZS.J5CR;5+DGe
+9+=F),_@FMT,419;:2T<bNP^JMDf22\R2d17<eJFJK[GA2O;b2A?_&<)O4N#YHO
?<,S0T\=T5O>M(>d6SY9NEIO\1^CFdI#&7:S/>5e:c-X,Y>SIPI>J>Q004^2(f;P
Tc>\+G0E<JL=e[f-47=-G703\<QE,BGFE/ST:OJ><0DREE,GA)8=^6LJ<aRg-/S8
Sg+K_<_XU&I@[U4RIV9^?V,[[68VQ7S[P<Od?HYX@4MWa.#P0+IJBcI7HPc272^X
<UJ8^\,aU3M\QFgW9Na9D<La7,[(()2ZC]3YS>aOR.CU_[+[WHR101N0Y+68b1\\
C](YAQVE(d;#gF9F;L-=.7AG?Y>CY)5]3>F2&T^H>;aT:BBB:8@bU,b)G664D>GL
cDeURZc&^0WZ7WR=>^:G6#@WfNF0\fNeXMXX;/<=LYK(fH-)VgW?aTbcRcdd-(0F
U/;]X2;?Z#-U<HFS)0_G/NRX3BI[84UGa\1/YM4=-)3P=).T\Z:&PGJYbD7g]b2[
:Y51Gg/EeA6W+-_M3OcbLgK]=e,NN12Me&S.;Kd9QYDE1bQ9<;WDgC/UHB8[N5PK
a,)d+g0:L2WGT]:f,].-a[(;bEBB:6gJ)<7gb7F44GfO6I,A?Mcd-RT@]c>_PC?M
;ZM<SefR&7RfW]BR_DA]1\B1,8e_DK\c2A:O2SXI,\#XcA6-g?TD/J&B95D#9a=]
G&ORK3C6\P5K3<XXdRdLV6P3<a?J6V-/SU07@6@9W0b<D?/c]POdgARIA:c1T=;b
V>S.=bU_8J_-9TLe33F.(HS9LeC:BL@CYET66a\83FD@_cOPBKONDH\.0c8@SY.Z
fK<#P;X(Z@67UTBg9(dO+Q)/VJ0F]R^)DSZ7&<CVgA8,0X8)c]0>ffYFL3-R8J?0
AJAKdV;1e=P^SN.)&NSG30a^[9Y.Z64M;Tgb;cggc9>0I0Q468.,fO0fNW<FNAg<
cTY2IfW/E]Z+:/.@8\845:D>V0+;+)3ON4[X?2aE4B;0Z6_C27@0<J=<>?&e\^QC
(G#T,AAg=0_cC/3ed&7)QKg6dYL/.Jg1;WUN0B@Mb=IKIKMJ5#,)WgDY-#g4U7M<
+2L&]a=A0XV@8_^3=]B0-e\Y5;(>Cb]MbEc?RRRM+FKeHDNSPZ/F#Xada<Ce\-Z1
(KEYY2O/AQP_7?e4I?_Md-:g4+UU],1Se)bc)&g[]5L>VGa??g.U]K-HO?aVAM+V
g6U_K+1J^KJ\_eVU.[D28D/#Dc@:@^IQYGNNM=1cD(5PX>-<W3P:-C(TRFA>E-C@
<(7<IN?eQ=LH.e2]PQSDE82P^@Z;:&U8UADgd(a1\=(@A)7#\?4\250c)[K6JY/I
W=BDQ=Id-J0W6Ef@a^=Xf8C_@@IPPb/cNAA3gO9fFbFVS81-b8698HMI9(37ceQe
JN2(3E8.-a,N[Y+S3>5CJ?d,](:\V7)<5N30ZQFK2#:NIN&L[_SP2_GOYR0\f_ga
3b&f9JIJCLPM=,MQZIY#EQ2VaKQCFc1#ec(;M0ZeVSA0HL_>IHSP_M])T,3;gQ5a
A36#M+BG3@NN27^O:T[\.&0Jf-I0/-^g[9@7U/4V,H;UUTgMP;U_RHDd?+>[LHZg
//BdL,EJ1K^2T8)I3PMa]_fXSN0O42fN9-=UN<(+AVf7K,g6cCFNQR/=-R/9fC=d
:1RD;=(;-+AOab<ddMYS:,OT0,a-RZCLf[M.+PWE0_29Z.G)3^;Xe9#ge(PXRAGf
1b\+<W-,_G#bI,2_WQ&fMCMML@JCVX7QBWXg75])K6PEHE1N/EAC)HG?FRg+V\1P
-60DH[e:&#^ZD2]HKa?ERX/3;219(W1J4H]3ZOb:FPD2FOH@5PVPgODJ)JE]D;,R
4;c#8MGP1EU9bf:-2]T^0ebA:Rc535.P18@Y?TBSZS:N=^1Ne:<F\F81J>=Gcd)C
K6SYf/eU9S;U^VfPc:^dA>LeO@4ER,FZW&<Y7R?>B.CMgbHY?Nf6W-A7M4#6.f2-
Vf;,/W;ceb?2V6Nc5[+=3W.^=N,0FS)>^OWNDC]XC,X:2I;[/#&Z/LR+1I7WM6ZY
;IH+Hd)MabXf.Q[1\-IUHTfgaSb8_:G6TaB&Z8O=)#L02cg\/;+X&+IGA8RZ[/@Q
__BD,+3e?YJS_<Ie-e&JPJLU&abZSX@:Wf/0e[_6#Y#>C_VM,F-HO,]X-\f:,_NK
.ZSG@S,J8MP,M[cSbPY=Q7]eD>/c(gV[9FO&Z@Z7c302HZ9R&>CfI\#5Q.fE0TaT
dJ(6]P<H03>-D7F]/?S=W/67?&G(5\S;#1RUOIY8TR0F.=?@dXFFOa5HHJQ+=^.L
bCOK8-4=2^-6G1c68&ZB:_9Fe[CY^^9O=8gORYJ8FM[3bVH?.RMN=YH7HHSF@O29
Y([IDfIL8Z83W0&0+&d5T]cQ_-Q]M#Ja<NeD#_[XQ[NY+Ec,NM24Q[Wf5C3gbSa=
RFP,0.G>X_a/EgRGPR;TOM]6/=(1PH)E):c8G-ag_?VTLL9PG3](fV4@-g<[[;.H
.GEMZ)Ub((N5XSd[-)_F?2\P+NXZ\.#4>534?e4J=7Z1>c/9#CffPC]XeJ]fa0[@
LHI3QI,)=_=;d5Md-CdA#=5CU.fVG-SF.KD[LL@<0e+]&d&cPS1]aZO6D7PeURTY
7O2&+_YYB4.>[QUV0Q\R[e?gaKJ_^>1,E969<^&:V2>Zf)5MUY1)]LfY^I4J^1;O
FXKBSbT86T1LU0#Q5/,=GZ^U,Fa8-A7XL7[2K^F7]2ME?2]:8JF2;;_#Rb5J(Q,J
[U)41;^._<44NZOSV\HN\;G)gF.@Df[1[4NM<>0O;/QF6G74K6+L_X=A)E:Kb&2a
WYeV8f5IR:^:6_>/?HQ0\UUM[c\AY^EBIZPSEMEOeZ3._PRMZ5:.]RUV_[P0W2cQ
79>EQB,-/;/81e,],M0#HT,GUf9.#YC1ZX@/B=^5G\1^=4+^C,.cG-&WU9IV;SVc
U/HS/+.eIJ16.CM(EgFc\WY(K(O[ER6gAG,c,>II<[.(\Q\P+YAET[Nb\_^](,L9
9Jf>>2,L)-P)27F;G\:9<6f5V7K,KK/=<2Ba;GKOL>Xb):,62LGN4/<(<L2?c?:>
,;NK(J_L:WKH_WaTGD^J[4.[&W)I58^HN?UHeF0/cK=CWKU=<S8MM=T\L-dRFf#S
HABC3#KWC;#GA20<]W7+CIa#/1-]3[?8>gfCP1H@JKcA\J8#\EGb>@4Sb)M@;=E+
1ELH_cb3C@0@:2\<;?g=?0+XWGJ-59D-[.7DNF_GZV3e]@5VUG=3UbDV>E8X/R<g
5_DDX[P-LP>\,))W2aR.+@QGHX_O3[a)+G,d?IYG>-Oa1C5C6_]>KREdPcC[Q/VC
O0;4J&f)_4A);D]c3B.eJAQHfg6b#EVa++6e=7f/H/3_\.>2/F/Xac43<K-8)X@_
R5-X^L1L9PMaOESF3D:NAbF#D=X+3/9M[-=WI@4(K+W:,,8&3IBTe^R#[PIe#W>D
;OcB,fNU3+XMIQ2XK<GE/#II[P_Nc-d(K,@QVQMKSR6=5:5+4^7(DDE7WF:WGI3M
MHGa#/[VEK)MC:KU>L;6e<0GgBY[O?.BUHV]5O-]B;CQ[ENIZQE80D+eMAeS7S6T
1V6>?NOV-@9J7_-/?b@A84GCGW8ZSIaM&0.#[-0b(=eN7]JXZ[[[2\>Oe80;(&,/
WACX#Y;SJ\3b3H_3Yc5^^\a5dT7T,[K@>cVK_;((/4&X)MORR@E?1ECU)11EGc_[
Q@?S-7WbK.c9gS)XG9-4/G5F-/XN35\_B7Y-a5DE-13]4N)[08QJ636[dH7,1L>+
CU_QVOG6-_DV+555CTR^6]2e;a@@A6Jb@F=.aI=NW5P8A97(^\NBa77]&0:S?.aZ
&O5D\N>(?L_1Z=,18#?T7d86e:;JM-J#4GE;=]CAWgJ45EWI3:NQCdL;(Qf1eS=^
0-]8dQ61M[BI-_NQZ(H.N/f&S>2X]7/\@<GIRdPBGB]6>a#@e]dOge&g,GaSTN:G
WKD.\FVX68DR>aMgA#[e=1X^GGU^@C;?2OKRX6FOIV60,@J6E>b]QI&\5Na\:<EX
g(P<7RHLcQAE<2LbUHaa#&,]fE8XP&2?a.WX0-\XID]3ZI/f>+99I&?02/cQKP&S
X9](1F3:&c1SM#0+Vd+M5<X,(2>:DQS)c8FDF5YCDLIESZO+=:)B<VK_&(Z)TZg1
0<Z9)R(O?+5EP&HV;32SM>\T>R-=3OE3dG_f[f<V[^a8.dRaZE:gLV1T1a=dT<Z(
LJ7a(@;-EXXLHOE>I?1IJ=(0aAeg1T(bQa36/4IX9>>NNfC0e:M<F<I9=GBT5?H.
.=8P-)&ITdQdHObLKCG#O;.:UKGOX+DG-@Tf7P8d2C,6B(+)6/4TZ<0fBOQ4.9EK
BK#c#)6IW1OL_BJE4G/=4V]&aPW\8>V9S0^.5bVc+6CU;A_S5BIaI@MS3P\LL9?M
09M50=@JQb4IU5Iec:bYTP;#0_)56\P0bS)(8=ML4/.2/93F2Gce@;HC)23<YcM]
(Y)C(,.BM4QT##04&;>4OBE39A@^5N=,IR9A;ac;f^523c]5gB0>a1O64-]CF)0J
gYK)POEH_I/JG?8Q:07;3U:2L<WK0^YXG-RFOTUA/;JFea4:=cRU&5\4b\U?^Y_Y
UW49<Q+773[JEXFSJ7U,&Ug?J)[/c07,T7/cce6.#1IAKb+JNQ8=bDAH.TV^=-WH
^)QWT]9KQ>U<FA+E[\6,U.GcFT(\RP__K.P^38<&FBQ/N]db/Ob:4MOLG[bL3JTc
L@Ze:0=Z>Y\]GG4Cf?]UK66KQO1MRf1ZUAF01J=(aQPP>SfZ5d5W+\/Q6d^X)=#B
_95U9g1b>2R[OZ(fP),?)Ab-V#SP(Z?\LZDb<2X+M&-J)@U^;HGc5[#]\GJ1@SYT
2WG_gIS7-c^M:d:)O?-WQUD<S:8/FcH;(,f/4.W7UYBg;,QG9C3BZY]a5&MOd4cR
;X_a9a\E>Ygb&bf+]GN+1Q.F2Q_28[9g8P)8aZ([3=X^OZ0ea]O&P?<:])ZP-PS(
3,96EQ>b+2J(ba(3W@,M-Y(FYO,4B+5d=3ZL6G7A]0PKOXRZ0W<#YJ6Ed^LYHN#@
QaA999f2ZA[.G-_+@>GH9IKbPbBXbABN4Af2Z;#L?,F]V3eUZdN;\dOE>3Y(Z1&>
M@;a7EM@XU#C8)EV06.[F.&7T/4Y)1^W;]c(WZ7O>9/I[2+11;@D:@G/7>S7D&6c
^8[M_M-fTYeEZ]L_GeB<Oe6g3T5/PXTE3ZQZH:K3cHH_;N+E^L.(]ST,&3F^>Vf;
6@ac:Ne\J]EYH)=2W[UHeYN48A8ITTZ5aCddc>d3J79EI.<)Y?bRHJKR;T,AO[5X
)7C=[<Na;8Dd,Ad1NIFU@UT5P[N73.KH0DAEQcV&b&<NF-Y4AH+g)55DVNXNaQQ<
Y=8R4GcO@^N[-V1CVVH?-5d>#,XJd3f.I#KXJ:-O0D]&6OF_&L+ZS(3CO:85[>^I
[G09=.._O4(acbQ;72Q_gb,A_>bRVX:H6)aM5D;AdZ6TRA<g-WS1P@/XQ\(?TdTX
)KeYKa(Q+FG;ZCg9I]7+/:Z\=23&\7UeLbVXT(Z\9:-=D-aU19Y0T/NTIQLaYecg
9@-0CFeW>]>7=Uab1=I_:AZFVKCH6X^ZFD-_37HAIg.Z<Yb.0X0#@KKKe1SV)g#F
37W4O#TB48N_fDBSB9?JI[2J,0H,f.5]5@aY[LNDGPO0_+3E0)750XPIY(&O82+2
O0IZ)<+<eW</>SV:3T46/gND(cDa80S_d/>K1]Z/QFE91=;+GK<eLOXeU7N9<Dd5
,UKN7;)0&S]\Jdb0B<&8aGgD8FT?CX,NYA-4@V:Qf7&&[VOU8IPeUW1.L>M2B#QP
OG7]#=U3^0^cBV0fED,)47_5C?DJ?C+VRRJ1NE.?-I0:24H\AG1:A>9/:cH-3gJL
0:7YZ0XSE#Q)Pc[]-bDJM8TY@(:E6GS7K^0KL?HV[CEQZ>38BY(=7IQR;YEXP9J#
,#aF0PPRM9&>J,cJGY0(&VZD9(C@C/M(H.6d1e0C^fU:Zc^9[5CO7fc+@KdMM\C^
NTBa@D2ALBOH-B,3MUCKWf<3bdDAZ1=7U/Y@P8)@&&?4D1>_b]M.aVA.)N_I;6[a
d@/dG]O7XTIDPIB1TN6H.<Wd\+J8>&\@+XST^AC5NCISB/aV=OY#PT^5_A]cP7fB
;A?;SQJN2@,1VGFG64]W9,=SQLeS]\B+F1@HQN3<>8P3;b^ce+4V5_&c27\PSTdK
++QD>)BCfI_9Y90,=SeKEMa:6CXH(gfPb;C8_eb2(XMBP)EM1&([RLg5^U@VGE()
MN[IP&2=+P_=aC0?BM^U)3\K1RI8T[PMZLWS9T?BUe?TN-JMW@36fbQ>Cd-:(FM5
D:E@/+Vb(@5/W+6MG8.](J/a8+0<ID?FF(FWDVMEOHJBL#41b2L/Z&7PJKg6Q;?:
_HW30CYccVKdS:5Y.CS^LdWOaa6T5N^<CZFP^ROf+bH>d2(=Fa=0gXWA8dO=gQIc
S#X9;M6=Q+MSMgV7\O)ZD-6.H)T+4\MO(5+T@&VZ:@eTP9@5F.:Z.ZTB6:f5[+#P
V(K)MH4.N)G?[fKbLaCbVSR^^&deSUN[eGgN-ZX7[bZTaZ]/>#BfFEg[6>Q]G^C/
<))^XQC^A-91fG:C,AV1KY>.Aebg<e-A_C^ZG]G6;BWVGc+4WJebg^fDS1NG&6-G
IR1?-7(&_Q6MfX3FT+)6SHd6YY<4&=Se+HEWX[.+[LM@5<7XYIWBCSQ0e/^KBg[O
\O8dXOgeFBg4X7S0@5BJgJ9S_<V+TK6)1@?(SA_4@&.-MY]&[0/>H&=#PXeEcb:1
9SfU-+KFdOYG&1TUCP]ZC+UYL#=5:TCcD&<b<]5SaY&]KgL74.-CY/NY8R3#Y=J-
N4>5JeIAN@M-?IB106YQNAAUQYHU:#S_+P_L2@MWb1J1K0Bf@e<-a2]XeG9K\YH.
AF1)Q<(EMObdC#M[6JK8UH.2fc(eUGXO&_&dX4L:OZJV2>gT)C_4NNMOJF5R<>eG
)BaaVXE3>9fa&;df1IEQX(RNETC7X]-CAB5CBKTKUD>-:(J^N6@b]:LP<VDP^gEc
gS)&;ZFH4EDFMBQ:#eNIb@C6^YZNFfd\<V+GB&f48::M)N??LDb\+)\JI(>AeODV
_.=#EJW\+0SK/-Cf-Td]IMPAJ1<][97D<B(bbTbDM2AAcF420(84-H@LGW4#S_Ge
7,12<FN8W.>8ZQ>2ca>YMJ[c>3c/Rc=OF3O5Zd@<ZP?T/&/,<SU3a)6MJAQ(BK^4
e^+9(&f<c4baYZKZD4821GD3e46ffT0NOLNC57PLgI8SXFXX1;=)S9B27,=A0,F.
^D9W@ge&XAGV_0AEZDEHKOB<3L8b5SGgAf5TQS&^ab14K[3d3-c#^^4Edd\IeLIb
2V26EQN@#X23X3=DJ<QU(2bb7[#QR0b[O_JP^H^f(^]HHK7dCPB--TTb9VDAO6MZ
5RVX_SNAIBa)R=Y=\-KM_&.44889X3[5L;C5DJYea>RZ?(8dQa=CONE_]\a^g_Ha
1(AM/<X1]f?0Ae.Jd=&.FQ\&G[IMJR<T^#T/GI_B8MVL.F=F4aF]D+=If[/9HR[D
eT>SD(99GD6_X;c=1C?<M_<E2,d[V58bRZ-N?8-&AM21E9J)TccMC+(NCDYMG&bf
+]dZc?MfJ^BEdXD]OBRH:>;??KN);H.EL?TR+BeNC4\?<Zb;^.P)65>/[H+J/+IO
gbSea9IKJ+8\D30[f8PET4Q>Xa7=OfW.S;H0]^MDIY_N<Z__P].)c?L^W-b4-U;=
Q:S\Z)NY]d8_;7XAaUQdJC;\J05<f:4I75a/_M3]XWLgN4;OJ<:W#H8J:39Tg=V2
UfdR#&C[SKYgX8^aFPQ,5ZR)V?RBED,XFY.^#A4EVB;35_La_EX1_[5+I=<JV4LQ
@e01FD=VfUD#3:AQe)NOC<.4B?c+[Z[eLdH\DAIE2e,&OL>\\-UM#9-Q_S3?L<#f
Yf(/aPJPPC+WS81TQ].#_gWNGU@#aI;OW&NQaZQg_+Z_K04:O>L?_H0FVW/\PRc+
F,#REQ3SC8&AQO6WH21_U0S<=JeKA2W5a4=5-AdQ;(U:ED>(Xd_3U0d#f5X9M@)V
3>9Z]I@0.R4Da8P4F=^SKKIe[.S4P8[>(VY)UbeXc#=E2BO\d_ec\A56:Ygfg3Zg
KccR6GTKO2V0]6SYVeMB==dF0&O_C8&W@&5W=D-KS-/+/F+f2[>a1L_5WQ[eX_#I
1)\e47K:1R]>4/ZPg9@0FF_(0+O.)QKF-6E\K&J6:YXYCN&)e:AG9\/1]T2V&g+e
0Fa:W/;7<,&&\eB9.[V:(.9SdX,4L3Y[]@]/E#UM\+.0X]S#<#cVEL:5&C;#@4d#
5U2Sf=/9/b#V37\L\ATHXM5(Te6gN+/D[eW\OWR/TXLS;b0/EBXJLY71R&Yf6?E]
UHV2].M?/CZ\(@_b;DIX9fd;5[dC]5Ge>#HE>c-6/)J(b9LgQQWY;TN,EbPE47\W
T:U&1[\8PE<]1W,Y89(9O6.>G/>Y&KNCV/?X++a7f@BU5HH3dTUR&I85&;d]&&[=
L++00M0FO\\OW?9a)aKG4L]1g=a?GK@+96OPS#f8/3,R9QI@cc.CVUSDa2Tf7Y4V
&+K.BeCcCJ83Fc08N6TUEJ5:7B=T50T7;a@^:G>000+Q&Ae9D\(^LQO2Z5(Y3J0Y
g<XE&03XSWg<.Q)43b;FABcTZO45XX/GU7),)@R4FX]+MeTb8P957_8Xf-Q.b:KE
U?g)TRK6:RfWf7S(_Cff)V<+.YAE8aJI90C)2RFg_##eQ]6F2U6_#O&-\1;gL8>Q
]MP;(/@g]@fDQK2I?9P7VBI=L283/[F28e4)0J4Mc-9=9F1];U?U[ZW+(&/O75B(
+IO4g[@UABVJM0VRYCV\,[>c>BL1&UG+1#+>/:V3IgT,4.(>(X6T6,0Z3UB=>&0(
;U8ZP9/LNH+RPX<SW6@EDX).D63(S;Ng+Z)>/?e)DR5=4fg6XccdF=?S?FJU&FR8
L5YB?R^=J6^9E/;OAea:WN@M;]a#9bX<Me=Ye>1>AW6B8&I6b-HI<RBZW19b)gU4
f:A\L,BQ.K_=8-7&K94ADFS2L&FVOA/56E<+#I8PV\S<YdDN&)/O3_)3CQM^+1\?
NCdK3U2_F)_O0WQV\2d_^6RC(O.)dG<f?I=[<XgcL]A)0CY@8Va/5&e#(ZA.;f>]
8A_5_?(EZ5ZU(J,_UEVOXB0H<P3eZ9X#:[B2:)DK\DPO8@bY3HRTT2#aI@IUX<#E
M/T(\<J(ZEcTUcW1=^ED,<PM3=7d]f\&CId#RY0?fE_Fg@+1VY8O3R1=-](K#4XI
&&#9NU+L_<Z.Db:G;&JJ86=]X4&bdBU(?K?0:1e=@3\+fX6@8&QPGOZDaAO+WI;]
.-V4B0Zc7R[D6L4H]I#CN8bgCBO88G2?Yb81.LQW1db4==QMLB()HSUH;Z5]^UO8
?/[1gJBY_b[=0gT/Df=2&)#9#aQ;-ZdJ2=I(Cc@HA(=W;#-Z?Bbg,Q\C2aCLaUI7
BQ^OgF\+LOVEW@R#S6RWNe;c/XR0_CV54\C[E6?e=:/J&@7dFbOWN>&A>)FO0YHa
U9fGX6P>=C.-/D.E_Fc02-ZJ6.M&Sd3F&&WTLfbF?(3VMbcgEEWZ,g#BS>Q2aLaK
53(.<B.RG_6XBNCdA.:Fa4KI97OGY#QHOdAVD5D^If;Xe&d=_^5A-7ENf?[FA:0J
\>ZE926YeJ&SdUFWcIL_a@)S:7+:<-g?1LEeG-U6XOdHQ?&^RN2>HQ]?80<CV1BA
)8Q].KM;f?7/I\D@XU&U=C+O0Y/08=74Z;7c0MD\\.VH8a\E2T..4a)1XfD)B2N#
[f;.Q7WE4&R@M^T)afNM+8-EFGQ)XV,MHG?)5W,K-1eW\/>IWgGS(X3eMFdVE\)7
IFS:(4dP[15Ze;H8SVAJ)\EV0?FORLg>Bc/-JPV,dRCe\UI:-I0>Ad-dYEA^XD(G
@C(B#&:(Va;&>AeM7].C@L[Y?0KL5;GHGg)+71\H:_aRE?8@57_,fU[&3\EVPA.K
(08DIPUT.T/NA=6KA;Y4U+#b+S..1&_;\84&7]M>QSJFW\;,++L9W)dTUXP3SW\S
ZF6.e^9W-^daI,/g(?6\\D^eT^_/)A<H&VKPZ8fEBd/P5ZRN<GYefG_IQEX1),73
R4K@ZAU>Xf/ZTP[OYP)RNGc?3M]<-<&H9L_T4Y?HgSAU?H+9JGE9Q^NJRD:bb2fZ
3RVb=ce3=PX9YCH[.<?3E<DCFEZ1&9d^92G]U=b4N[6F)SR9+0E]RGcHg&FE7ef(
bQJP)fS.9)[b;#4CQcffY7?5XeD/RD0=69-HgC-7Z=A1Z0&J&WE:?J9(.)?-GaHX
#XEf/c7c;f-+TC(B<BD.]QM^@00I:3cY_QZH@-V,e]NTU_:^JGY=cLK+.@2+,QA?
<UD90H3;gMff>25(@LF.R+a[)YH8B1/Q+>#=S6Ye&]?UMRHbHXK5RCRUI<-MZC8_
@K_@X(B7]^\5Veg4JabUSTEZ:gGdI<TdEK]6V\&Oe21KWK.[4B[>[_A-Q3E52)gQ
f&Y7()I)_K,dG,HKHO@KdAP00.UT_4[1-BfQ)>#Y=,V4ISAWMS0<>0F4PW(VEc^N
C?b9[LI4,YR.eG46Pf[4-HZ>9gWg1.&1Hf04WFREXYGT+/]X/EN]F[U&+Fd87;f(
@I30Bd(fAGc:QMR.>]RFGe#Lgd/_e=J_9d/9+K23AHT[fO@IUHEN[f5#>&EPE6Pf
[);5#GM@TPZ1QM<4N(VXR2WC2+bUHT]>H]:6;2JPV?0Z\051UZ=H\DSXRDL^418+
KZeM/e1H<B(Of#9MHVU8J9()LHZV[M\RPGNR_-1<>_C1MLTaafg(&K6U-7##C>V8
46g4#0#76#aYGR+/V,FG,+P;ecZ\a5M-\S>f.LO2:e-P<H(BDMB:=Xd.Wg03LLL\
UEK<62@JZ48).Y>X[:@eeRPW1VY2Z6=f.9@=OJDf):)KP4#YA6Wd<B0X#g]SVIP1
;S)X8:+?a)_(J;f29(+QW_@TQ;?Hc7BLMU<TIG\JObTFA-56(TIJ=B>4;7c;VACZ
1RUOFR<(aN^FJfZ,,)(c98<aDBW4ZM9_H?bG(R.C@FG<V&<O3((-MWSYK2WGJdV)
2((1-gB_-LILPd)_0X0]B^?U3V)OXEg1KSL8b=,J;_J#XE]S7=L]A>bA[-7R;4QW
,S7O4cQP,0C97S\Ge7)b8g,AC>d6YVL2-C@G(BV-[fH\/-T:S0bWPLTb/D8R0&XQ
M_<1M;ba/0+353QQ?8:.]G<TQZ<NTUG@P\B)NL1/])G\GU^fQ/;42ZA):(\f#IMg
NZIM4-0;0Lg23E#?AYU5GU=5Q4a<>.QMZN(cdCSVMfcYEIF5-K[T>e4ObAb2LJ(2
STZ8H/P[RUUd-6WE?A0LK\,>+CT0&K&K21;G3TN=EGVeWWeadFR>]],?N&e#T?cW
9I#D(AM=(:+L15^L:af&JKD4-X@_O<ad<]?;N@T2/3D5W-5;GT(F3-Vcb+d097(J
^+EW2YDPD3)e-g,Q@O&FEXBN#E6+,;EU;]1#,+/0XV_9e[H[ag:W7]/P:;D-d=/;
b#J#15DScKe+OIVYN)>gbK\MED;?6@8SK.(3UZ^eI9gGANJ-1HH8BBK2^Gg-?Q6;
/_QIG6b=Bc+S/X)\J0O.N;MI?aFIB28HV7:-I9Z4;R0^=M7#aZO2XgL7IYY:\gZ_
F@>:()B:;G8DJPSg+0d5=g?,\UJ9MaI.IS5(0YKeKCF8N>P3+Xc)3TgY4RF>7gcg
FL<@f[cOVV5YH)H)T-L/:::c;ECG(8c77d^C]Qg)X\>MOOW#K8&.1:;_g5#c-H,Z
/gb<2@c5VJ4(+FWL;+MCJ,8caa(bILN71L^E7LKIgD^@2+2-V?8bb74LCcKAL/^P
C^<IcM@W&C&HQFAAJeCVG\a.I]:424/?<JeGSCE+D6^X(Y:W_J.N>W>9+cc-(f?<
VM2K-aaIJa\fY-7Y\BbZ:g-57PT36,=-FLH+00#B-ADHGVZQ07B1NL)e#UG8cdA6
V?\Hb6bcf\?B=?8GO2>0#RO&CPceW:?6W1ZF6H3?P#<M5TR/gNBE0fHZ4[](R@5=
#]:,e=LCV(7TSdH1E[^?dUO2b#T2;RMP/e7Qb[;5ZbN;-V\RX\SVKG_I_<M;-I5#
48(GaRP7]RJ2RL:TSW^cdgPF5;d0e()9<;;=GgXIAZeNbc-2GP1CV3X98gK(bRN6
e;\9DfCU7e5UO#R:/XB<QTX+-CSdYL6Q:Fa>6UJSc93HY[<LZ2YDY1O0T/[f#IP>
;:Wc@EZLR?8-DI<cH3K&<__?EIcM>Z+)T[c/#>CKbF3OU8XB8dLdUSD#(<M\gWb^
6VK=V1\a#7-cG2a.Z/gOJ/b8<B\e6;JLNZ2@X0R(d;?A#6O46N,=LW?(5UWTb)+4
/2QZIN2V94FEIWefP0b>:I:aV[6I,M,3,Seg^6]_0^(>DVc6]T<YH2^Y[2=&Y4ZI
B5,H;8fTIVJ,QGO5<_[#&NWfeQY>GZe[/UWNRD,0TT^HE-4EOLf[aKZU[21TMR&^
O4]\PKbZW:/ET6gC1I#)-KN5/3]2dfHQ#CWTFJ474R3UQFWPD/D4PB9@H_=8M)Z-
HQ:gSNf.;SbDBKU5QGBC/53bcK3I0TU624Ie1=#CQgQ,eUX:776b)b[Y_:E2,e2\
5Z2aLLe454;XWT#VEf/OeU]FISWR&FZgLb0_E/P4H1K]Z(5B\WAI0C(#:]GKWQ4e
K?4Df3E<C.:[VICI;:44GAZa74g5JK4BM6]B>_E[?2a9g+1+(255VLD8AT[Q1TM:
e6aRcS+E=-d)\.4I0F^DQc61Re+BH/-PE:TY#BfVVC-,H0[@/2.F=390M2Q\TM1I
BJa,8#QdVPEMR,[]XEgZb/P@W]5e-eQ;<42ZcIM-Mb&M997590.0V:RR@ZJFBA3P
EDXT1=L:JJW98gJX/dX^-;DFG#c,9.Y:DK>FM54J?19b).Tb8C(L,8W/<EE4J.Uc
1F2c1SDD[J^ZDUYDO)N_&Pf<Qf6;?8:\<5NLgaFHOX9QRXMU2A9@eMZ=AZZDV8+P
Aa_Q[2R8agIeZ0N:LOQQR(]VLE.#D:]G>-70XG4F,73X)QBI8U-1<@N[T.>M#XWA
-]=6PX:?(J9#4^3#Mb7ZS1QBB87R=XB3=ggPHEDXdQ&JL3].fC?;FVY^Z71E;WV=
a1X/Y(PQ@>.]Z-,T#)D30daRBfOO,,T8.dE?K>Sg]@TAM&./3a^ACY)^NECFC.?]
D^A@@5>.XEGHbLU_K[CC\JN:3X\P81P4Tb8CTW>g3>/W2,]DBPG\L_Jb[+/<;GY^
<Z:78Z>>3#7B.>JMU<RF>XXfV,74K+f4N81:4Aa-ZL0KQ&M2Nd(=,c_)Ma:4T.+<
,OG.,2:2X_HVS.#7Jd2#]bIS1+g)&78/8W6X>.D2\DgU8d_[QC-ZG)SO;0#MAF(K
G8A]\T2XAbCag_IAZ^S7T[Q^YYB8;g0Jb;5NP>X;]WLLb^L^MH.,SKe2K>^2LS/G
^4f]Ue;^-DT]>^R9=3,X(B9<23gRTW.HG@d@^1QgbecGGaHXdMW+L2M(;TcD\d,6
1D+(DQ)=FRPAOg+DfRgENJD2aG9YdJE8Uf4X,5D+1B?Kf5_:.\A4MXM=+3,78YU&
Z8Z@ZfYM7OSL:>b2K?aa.+OU8dVGINd9:KN89RY<#ZaTb1#::4\^2c<?f81/3>0=
D5RP7@XYGYQefUT;Y9O+KY-\IW\G@_O8X022IabU-Cc>dR@ED?@;9W2;a7C+OXM4
ANVH?d8LH-I0=3-=+[UBJ?U(@=NV(ER[N2#=C&>7<^>HfZFIA)De7JaH5QOa(>;9
g-Q:2(:bP722IDbH;J[N0P[5>0.#VBC^HgB+?eR>1/D2P4]2Z1OaR;UQ&?g7Z7Y:
ZDe6aeG+8(_STC&B]O_2b1T:(UL0B]]>&VaOG8>,AT#/W>:34/SU53@?^g,3H=-R
C-);=<J^F?E9)#HIJbg#U\Ub0#4[gWG0ZAABd&BB07\RX\IJdKHZWLT<]9;d7g9a
PLU,e4a7E-Z2UC_ATA/XU)F_2\2BKC.EZDM#/f>a,4U5&KX4C.7]b5c4C+C(M8HC
+5M6+eN85-[acO4]9;&/7K].L)MAJWI6#D&/+_.aI^#3\DC,[,g6EbV(.AZRD4>2
6N;a_<(2=3_?d_[MbVF.C?;AC3N4CN6.#f7/SA[M0?)#B^ZaSW3cbUMee83H\E\&
J1=(0&^/6dS]T&b?T753HfCX+9_]b8B2/8b3F;VV3a631d)dY68#XBMU)f0+,[;K
7V/Z@#6]V#?(6PZRZG-#H4aJNROQ2cab[Lb==:X2d@\a-fZ#TARLSPNHZcS[R?V,
>fM6C54E=GYA.MCULG5c476_g?5SXO>f^[2Mc/6XJ7+MdFcVDCX4N,A#A&G<#\QX
2#HRS7M:AT5SO(#Da2>@HgJ.YBW.^D4JdWF53N(/KU\Q8gF&I9gdZNU7dT[eGDce
Y?[SEU9>Z8c\M_AT2>P(eS_)..g>\.78L-6G^@(@5>Mc5b34[_9V(V2e6Y7A4Dg1
_]5T6V2C\I>-KgC=[D]QS[SW;7I2dU.K+0N(&#IcD@?O4Na[6+L]@O.C[X:OG+Jc
-\9^?L/PQW9.b=&LDD4BSE4FV&D].daK;>>[JJeb^5/b&];(D02Kg]S-g?WW53:S
MaF3=T>WAHY(2S?[.#UJ@ES(-b_WTe2EEDBBFT(Qe)BBB;;c6O:8J:aVH6].K.NB
5T+D=L@DcT<ASM&/N3883]RE4;\+#2O0aR79ZeMPeJBR3P+DER32LGXU6R)9dMG5
D#GR^P;:<RaKNa^[XY.UUD/RY^UZD,6#V=dJG>6_\?<J)(,[7U(&[aZE35?_6I78
#eE:BA([78GREBCg,FK+BE,4b)O54PV_M6P^RG.9TAYI1V_ZSAb?35g&N46?-_e.
[X><afR2bUTCAP.,LFIcDY\\(fd;J3HYP,.EM=1;H#5UQDe&7<N+;\a#@979]4GE
c2U-HNKES-a^feIN=324F<d>F(24#X/S_<QZ;B,,0NTG;DKcIG0B9+c5F<@2B_G]
/2/)e:(;EJe2Kf#9J9fN78aML#@[6P_O3AN#S0/W=S.H<W39T@.b.dfI,M_2X]O]
8L^7J_:#&#2QAC=-b,1S>>5GON/HI(R)W.AZa-EG(F]RR_SH:KBSPI]f.6ZSHS+(
cDF_CQLXFR5>Dc?:>GRfC>:Td</8V3cNNCcK)ZbL0Ec)QO=_8V/-MW_=]I\Oa7MB
+PG3SH^EC@#MEHC&>&[N7g4_4X.g^Z5PfO?RLIGJ+/gg\-.N]B(.6JG<H;2I,IL8
2VYa>;+(-]YTX<;<>TY2,65U0<8TUO\578O/]=.V/?)EC9ACO;:3#L@;1;gKAMKO
].]0=Y1I[If)J-.,cL,,;9HSW??(MC0eY6;b^Y>;).)c&KQMZ5c#J)A/5#>Ee&N[
)>-GJ;8R<9JQ6D:gD)FgIR?ML3IE0;AHJc2-CKI>,Q?.=>CQGPI)>AJ+B9RH@4K7
eQO]7TQ7XHGXP7I4LA]UZ_@IF\9Sa;5N,EY[1J1YTdF3V?P7E58/>/VQ1;-U.]>+
TXR[#@?)1(\&V<7Wf/BR0L^95aZ^#a,-B^2YR(0H?&PO)EV@bbGC_,_8[gSWK5<0
?9UfM-M+QBCcZMBG/CfE9c23f65K3<T0,WT]Ta50)L;&9<=A4@Q@B0d0</,,+;=B
>NZ3G3O\bTU,)UGGRbSJM;/S:/4DaS6Q?R)Ee]LKB7G-ILVd-&W>>_IU&\7IcN+:
C;F?2)[H:-c8@()9>\YC?3:eMQ,[=b;AARBUKP(&^Xa6D0\@PLe/;0&6Wd(-8(IF
5Q6b45TaF+-O?W4S2ZT88<QSTJ?1XM-^MYAUUBQEI=<I<KG-&)_AYX8=aGD7JI]P
L@1f44<5Se;?A(If68,Xf_UDa1-->L=<eAaF1;a[./_IS1-GDI0F<Tc,ZEO/+B>9
CG8DQ]FeU(\YI[BVSf9^eFgMdH<;OF:EQ&14Q;TM:(8M11<@PX_1/AG+../#<#_9
),JdZX7JY0X/AHF5Tf3Vb2_YB&CYf3<TI5UQ9Pcf@8HWKD\ZH3:JPU,)WZ4bZS5d
(9>E)eXZ7\]LgD/#:I#+L:c&OG+?aO;LON+^NS;DOd60TXN#1Z)d]CF2SR-,>fG^
Ta.Zg@T99NBF<S40=-SdTJ/ETe8Q9?#@+=[P,cfMRE[6fcI,_4gC<#V+e57_X;&S
cHTX>)K&XYg16MY)-PFGD3PIGYPA7B7J;fc?d1RZ75?bYHKMZ3&0;7a/.WNCDVA.
HU<OKHECOT/35RdLIIbD7BT-(BP;RY_5^B-Y+=/>Z94(_;I4B-P@9eNXM=R\a_A]
E+5T3;+,]E\RXS>LSGVYF>R_D^E,@64+K66:KS0#aMI>b)FbZM&L.dT7,ORXabaF
V2Q>?#Df[[7Z8::L9JG?N](bHH7fQ5X_)6MTG3=GUXXS5#(\2194^]0bTR]3>&#7
7.E8>YFJ>6+TG]NNUgUJ\]W(]GMFZU?RZ6&5F^-Z2;5&&FZM]f3GN3#5YS+006_1
ZQ6I9(]GN<eFNgb_O+QaEAZTcW3(-6CNX@+Z7&7<g-7XQDHOC=T#TGSR0.END>Q>
D@I<A[aZEc<H3)-aBGJQG.49R+4&5NM?<EJN))ca.Z6T]G6FF.KN14\GR7NTVbgY
,P)NXHd\VU:T9&2D:R85BG1V;=E])]_]X20^^_4+_2(U/WN#U?QDSQ9#66UVXJe)
Uf8KF#dEOPWOH(6#]PEMZJ-?)&K@ICfRH39e[9d,&6;24[\.ZO5]/&;a4O]YZDAV
7O]@6)b,\LG&4MY/L.FcZE]P,@COBNgY>L8L#?S9GMd9aH65,bg^+]WX6;EX7VZg
O<45,<)7fDQD[8+F;ID1/8#HMTB>,aGcaW0..OIFXX,Ea-SBC>82W]fJ/)KYYc6#
:&c5Cb>=:e8fO0S1XS\7IV4:8Z[U>&IPOL?W>@X?cXQHKBW51,3333)Y_9;0Z;YO
CJJ(?P2fJ7O>OL.RHI1#9,0\+>Q2^O1g3SDJ_6PQ7e(S\I4TfKPDK,C?XQH/?^cV
(F83SR0G^1.;CWaD7PeZg?UNcB5YRYAIJ&(EI1d:d^MCX:(b-dLc-#)2QA@0N&1d
?>Y\NE<9TfS4=?Z0T3EY-+T&K5_,]OY7HU>;aD9)K0KdJe,YX&Y6@\AMF@-VOT^J
6SRaD/Ig6DA0TJ@K3N0?-QG.Xc)&G\&-MNYdPeOBJc8GB_W[#e7=aa<MT\B^ZJRZ
2A:-;HC51A&\Y^<bWd-=BcaKa_G^2eCd<L;F>-K3[KZI/b=RJW+(>Le5_>026(WY
8^2EVLT=V,WAJaSG_B-VNNg^UO2XH-0(-Wd@8=C<5M6-C>HAV;Q4C;c?ZdNR&eNT
f)M2,Z\I]KYFWMCT[AO&+gDe8d4:dHP#I#SVGQ0#UO-CZ/QA/8UdQIBJNQ=)D+CV
c=N7^HOSK;4S6N0JEKfJA5FU?&M8WM)Bd<.4:Bf+f#/Gg/8eYOJ5E98=Z24&?GN#
>^CVLD/b@97A-a\,;.U?)+2?QgZU9;#JMN8.8eEbMdE=5&23;d+84XL2O:^]1B20
gA-FKM@/)YFFR?aT<g,_K=JT5^1,S?C8e4?)<<>F1Z8;S@\5L.82ESB6D6R>09Pc
PQL[DLT4==aAI@:A:VY&Gc651IRdJN6cV\CRHcYOXeQ,SE1]Kg_D.M<0[M?5B)#)
6-P@AL@.FdVZP.aL@R3;2<>f8;WFaDJ2)DL.CO=ERJC\PbB]-ZWEPU7b^dXg_X&A
/Paa?TO?e&g&V[Rd(/C&R45+#95c[1S<&_R+4Ga/R)aPY3)+WG?[1#B7HG^[(D.6
I0-8+.c+Hf3b;Zd5+4P>)A7,OI;6^c=Hg)5O,<-[-R5OHEQAfVNR3U=;3\fNLZ)A
g;DW[Z>._=P[(^0&0H3B^J2NBUe4EA:H9.?\PY]d.@S6LgFg]HE2(f\8AC(_Z^J0
)K&Y3<-RU9f>bE]\-SU5cEb?>L5.e?[Z#55K=7<7BVK^R1S4K8Y+@U^/-Y55:;d2
-@cf<H&X3Y#D7e&IGJO[E)PQ@;E+2NO]K\H0:MUX7e?[R&]Jbcc;^8-E4^Y,ZM58
6,3B,TY\\fXa/;?6c[/d+#:_BWg_HUee[,Y48d@GD[QI=#8bQYgRb4=MWF5U=Tf+
BU>C5;JITXT4[QLcgO;B26c:H9P+^/H?&]PVL5Y=E@KZ5U=UM/@-L&)c,P.@7WYP
cDAO51M>5?_0(XGC.?a)4&g1?_c&bU_92Pc8]@TL_9.^-KFLNN#3W3O(O&+CX,4K
a<V?d:F9JHc-@(eRFMA2L(?eLC=KdU<MLfM<[3e2XJ96WCP1(GFa)#K8;W3WH-<a
>c1]WM_E^.TTVM@]>A7g?G64Kd?4M:b.U+4?T[0RD@dd1a2Bf<(,FWDC:_aSY49G
PDZ&/bNF7;a<0aS^?N[A5MWaKI77/d+LLYX119EK1D2+/a(@<Nf6UQ>=cZN,S3J8
KR=K2BG5G.EYJb\1&6>(EZeFcd-5](PfeVPYNBPP.C5UL6#b4W3/eIe-:]bC[;Za
G:d^/[1\;,U#KUeP\5&dJZ-g-3Hg8]LeaV0(EAcH(+)EfZ&P/4RHfbd)[e>_g&f8
O:be64KGgY2faB:<,?XEg)eQ+(e(,)^-X)(\WW[T-@Wdf5^#)f/LM8SP[X\d+]:X
&HF6=/@;GET0;gVd#-M;dBLN2_1Z>d49/F#N)]ed<Q@PaO7-c]Q)N3=0f:VMNb/g
SSe)Of;^5:_AA^9c_,cH9bR\Y1-&b:,+5U2XZ/WDB=KG;8V=9JQb>XV&cBHSdZQS
b,/RPBA]90?8TNAX\(:>()93ST1FQB7EPf_>.T+TOa26Ne@^BL^HWCVQf1b8b&Y7
J]@PU?,+bRMLO?cWJbaDaC&]UbE@UG:?>.d9aZ<:DZ6Y-Ebb-,.9c6PE68JX\]TU
N1;bWafJ\[)G3a<H)T?7XL>K2<(FDQGP,Q0:HO_,K0D12-H\3AacO<C^^_2+PL6a
RB3f_J-^<5V(3;X<1fGXHM70^U9:QHYTOIW5J3<]R3+<V0&Re]Ea&UN#@5&2Y4+:
b=HD5c9OZ]MLZV83M&+IU-Jf2RQ6A>a7.gTKfDL?0S?A4R9]IK]40+)]B9:)=bZD
^c/\[]IEFS3M\#HFGG:F5>W^RfQUGXDe[Z=V@UGU83W<;c;PC\Y2X8=YNALY/ZaI
?65;^\&XFVg9b;=(HMK^eT]_2Tc6;DBE7Q71Q)f3LEb4g4LXUf,WVH.UObSbXQC#
26+<IaEQS=2FfGeBQ92V1_^+XF5@d<IN#>V2J5/=6B6OS.C&=c+X1HE)3E(I^gB2
6f2@RY7Y^[>:U#@>a89D[>)E61&U.W#-G.G(9#?Od+2.c?V1ONA#DH+I@[<6/BK>
??G:@EMSKcT_YY@#EX),;1HZQcJS=CDT7OCc_).[]X_K2PgR;20gIM3?8RZ8,3CO
AG[X&7RA.A&4@=E4T6H6f5d/HR(0<Xd-6YDNbU)a7)81VO5:32X+J:d.).SY<baD
:1b?@</g,A09I<J_8?XO+AJN1+fT/[L2:RKS].aQ2gg/]@H:SBL[&8^g4JZaY]/;
J?B,O1RI7c(5-R6@:TNG#-4@I1,);>JN.b8_8)H><cS?6g5_2c0WVZ1CQHgdE((E
U4.96XN7(R)8:UcEW#Z_E.P&&##bJ2WN/?bWY/@C+OaN7T@\#e(1gD5XeZ#K.]I=
eAPQ0JL73c4b)LS2GWDAAH=QI/KM+a0A-DP6ISEX7M&@N&F8Sg#\)/K(eA65+QFA
L4^?J</0W?@WeXH3ZZ(:Y6RaV5-6/G-7CK^de]VX7\98g><WR+2XLWQ-Z7<G@[\V
J/N?K:5[]cWLa&9?P]G;c4ED-<B;>c2?bF7g9a_&-&9I&(Pde6UeQFM2?acIM.BP
>R(F+1?PU@/+5>7D)4SP>F<f3.:AVF&53.\NK[7^f4/a_CV7MHS?d@Rc;aV56OU5
<UCc20B\?6=V>TVGZ2W[P-<&TPP:4B>5L:,FUG.DH4Ve=g,:QS0D.[Od:85-VVYX
OD?W3.c8bZ&BL8[#XWIQ-[+WV8X44^TSY[;;URSS0[\S_?f2N5AAQ:cUG<U0<9PD
4f,5IK5OE&J\82Wge0Xe>5;-9FW+X+PVQI4XAV<fIZ:;SG])R:GSZc8.<LcP.L)D
_a[f2fY,OQPDOZ@ZV(NCWA2TTM)5PLP[c_?T23/-3bJY(.cTJ3^T6UHUAO(#IWD1
H1=^X)TAF)C:HF]P_K&1ORH1OCeHYB3#PC0,SBd&/_eO7[+W#N]I\MF(^)2#:<bJ
Q9Hcf1eML.UBWf[AG+8PDGFC)IBE#HIPQ5/f<SR7>_2SY9I;AYIM:Y:@cWVJ[:B=
dCN>]_PcLPR5P6M>2?g]g6DB>gQbX2I;aKRb&=Ra5;>5Q(aGRZT_X0HE+7EH2KfP
g_80(1fWd<K(>@<OQXE4bB4BE@^,OQV^GTX&20N0-E4EC[WG#3^TA^#@^Q9>HLV1
<L]0W:=YAJC>B.E;.D=dbY0E+gGe8c_+>d>SX;71-:XNED.QDU4U><[LZGVgadYG
JBM1E#7.+#e-?^Ja&2EGO8NAa?BTU?_c7.PA2b/60=ZA?\YYH;(d6a[b5+0]IKA>
a<A&6d1S0;Og1S01[#JMXH@FYA#HE2(6>LLUF+B>+:EW^P[C81V.MaVN=W1daTd)
&P6aP2BdTOF(EQI902.74]Q(9&7[.QR,72K+J\-[Y9Z:fK#9/J]5b&NAOLQLG09:
5K1\SPN#+KS[:Ve.S5X213[E>?TB:\+:?bR#[AK3f:>:7;URM,H#?-)@WJZ#RU5B
]\T/7D5A0N3a,]7^ZFE/,GS<OcS/DKV&@&DQ2VUO-;,PJ@KP:[Qg]gF.W>g6g5+D
\?:c:JOC6BgG=O&;VJPb(1M9V/5L8S)./JbJe[FFR5JNLPQ9e7F[ID/dHL>NSWJ]
.4Qe+O^&Ng-W:_,eW?&;8^US3_1:(,7T=Wg?8aD^&:I;8A=D@K2OH3G6e+6)FV(:
?W7K@8gV?S#Q91:c2=KBCQQ9&^[3W-+&9)[e_+Y;,Yd#2](f9X0RbCGIBS2YA91H
XKd;TK:R29g1]ULb4:QV3BA0B99QdbS^Lg];^a6PT.:31W0>XKLYaJ_-L;S<;HH,
U-8MH6)V?9D6/?P9085];8ZGdFTY\KVTAT@cTfCN=N+FHJ,78S<9+YH+[=\TL@?@
-7VE7Qa7ZfZa,@@:GC\eDGe5\JDZ_G^IgAG0OG66QL;#5I;\PVPfQe&9(G^Q?&6g
^<H)=&E_gd=^>d<f?NASDQcS,,1]#16W(B2gPP/]]HA?e=R]U4>GDVZc^gaVY,G.
\G?/QW8//<B\+fER2+Md^bOE+ITL=ab<27WRN(0+T.W2H#V=;4)A8<WF1c8gO&UP
^.\8cKYAXOZ^>L^@O3H=dDgGWN8VXP@Lfd4M\@9[I>@=[,3TOOcZWI)?@7)GPP0<
^,<T5]E6BP.Y3>KbOX\)4OfKF(I2BQ_A@#D30-07=>:&L:A\HT&\84QN\TCU9-K_
Hga@T?#(AS2ZYVD4P4@F8ZSM^c-Y1A2Q?N\K1^b3L#?NPcH.+9A<IY&+6dPOg\Ba
=S)S46D7O2QcAeHI5OFJ:53,I-YP?OAARZ.8:e5,f).]5#HUMGUG/>f=SB;fE+d6
Mg:X(MdU_fd-<Y+Y[Y\0KF#)QC>@XTPC2&.3[8@Q1gW96/W[RGF?;07]>R.MU?>M
a]#XM]^4ZWD\0&(9KIVUFfPe8,>9f+[C0bLW&Sc,e5POQ+-TWSMVSTZ6GCcI\GU9
d&5BMSH57+U#-::->^.fVT\FCVNa=T4Zg^]U]GS1+-9>1PA;^a4XfQW=f)CF)GWZ
58#S##X^DZD?HO@+YRDc,K8UZXf?G^W=/JR_JO4O,(OHWF7YYBAGNRQ;Nd_=@JRM
IFX^-;CcS/gC_PB7<-N7.#A\a5^,d8DEX+W0BT:3WdaEYSS\]/,R0[>f-5&M&5BX
:6N2d9ARS>=XCN1_b[U=A^<?)faPW2FWIK4AGefUMgOYDO5:MGggRE2cgQ\8>Yee
<X3\YW9UbQ>(;-];#R0fZ\e<1AR;?7_FXF+_M:^@TBSY5X+AB-T:B:KX.eba96H2
O,-\<WRO^7bfF[c[XA8[+K>,K[_X)N_U,e(I7)M472:&:T;bC[T70Ia-G1&KT.)C
>_ZWAJ>=>C.HDNC7efa9??_HK?^SA.5#1a839ME]1V1ZUS@4P9\9V6N3=/DObY=9
Z:J)1WLFE?O/3b4_]PXN#^_fJN:e/K3EGOR\gdL9RHJe(cgY6bEWL8dS[)R<U_[O
4]1)=F3b2^[><5b6IQY5eXb)O6ZP:cB1EL84=]C:JQdaY26-\A^dcM0^;)4/CTR&
;4_#R&(O_.)N;g[TBf514DRePI^[B?S?.C5OQ0+54Z-ebH<Md78c5^Y)[+B_=)7+
C#(3-aR,??W;3.GU(W+CE_,6-5c(9#@+R0=FM,1;)]c#KJO8?\KSCJON:Ia5=;LV
SG>R/6d\4JX<.-GR,cU)V?d^\PARDeFfJ0N]ZbDD+9[_<,8eO9;5FQb7(dfGMM=5
@3@/=-DQSJIc0bG\fD#OH]c.DCI1+/2GDJGc.[,-I6MD^6^d&67H)7XT/D^<3&-+
Ab5Q?I(gK9X?78c9Y)TdWOWL9NA]NPFaJ]P3+^P-L070P-+Rc+a2NcCOH.4A\^?E
7PQY\U?<Z77WC_;)74IRS<1/]4S:^E?VaE&?VG[\c4U9^9gK)H<_M<.NXY\IdMKD
7=0#=VA4H\0bMM]##VR,W#_E5JE,L[XF]7bW^A.&0ARM+Vf+BbUL;#R?-VG]>O30
BWCBgCD2&BPZH0+OQO)2gUWK\BG;^d8;TH.&+J,E+D=BV)#/O+&SCOJQ_ZKJIZSV
?OcKZ7\WNc6KQf9YKMg)B4T&5QT2[H:\36aD[7U:XJB/\+M+6d8^B<.U=Pd9Mg;S
4Na6=K9-.E]QS?d)[1T?Nd]J.E):#7SPU]B0fQFHKDOYKKKIe5Z&5<9N\-L9#4(e
#HXYT4/&H<PNA9:E?YeL\:89ZW,:=Q?DAHV@#1S?b7[d2Ze?MFVK--?US=JYE+98
BB<eC-VeA1fELP\7QbA2=8(B^O+[+UQ17CB>^e2=Y3aF)f[\Pf&/a0@d.d)eb,W@
[^7M=<2AMd3(LOKEfGGY(@5f.aU_AWW##B2#.LIEH&fT<,XDb<>&1^+K867H?<;E
N9Gbab@2P1FR=8C&b-.=6HGaY,BP)ga^XI]D(c-B/a=^D<-CFS-BM?8#f<(H)>CX
P,S[E+5)BOR(1P,G,1.RO9(MADRI=CU.=&RI3;Ad3GY-2V<C^S.[<=\d(HMG3V-A
@2#_9;:#.W7)0UMZ(L4D>VR8GLVd3IWd6IQP7K@0FUXEKUN1UEDZ=EH..W3;bP:<
R9a.V>fZ#T?3>U85#Z+_C-+ZR;FV4\d:3<G50U4<SGK^M0,YJV[==#OTAK7V-P^b
;1>/?G>I4[^XSgS60\90NVEZ<5f[L:_b^S6/24f6RE/<I;/6SC?-2CK/&IY-W-=6
BK)_,_;:cS.D-1902=M4;7+EG2;AfAUF&4/]OJL41YLL_7&fN_NDf?^COMZ0e.D+
6,(fR.aA9HKgMa<U;6=.3]WU4^V:8E/JSPL_b0NOU#,O28ZRCI[a5<[#[5f13\Ca
IbDZ3^RC=X.1@&<c>HVd?QC]OHeL36f5/DOU5]]c:PaI3d-(=-KGW9U,I8])2AC3
5=&e1FRN&7:U=(:B0\542\0MR\IUI0>c.?B<\X7R.]aC/ORXC]GM:\Da8c@WP.M=
L?53?OE1SafBB)d@DG>7QE1MH>PO3DK=1I?b;MU6c<#&(0-NHBJ=X_+W&.5N\F(d
4UN3a&bN1-0@.;&4/SVV]4_?]e2HFdb69V/R<E^0]->Z?^P=7@/DN62=:c3(T)>6
YU2N3&HR&ZcB+=1QSLT)M\+\#_Q&Pc1.a9S4]Z#I(g,0=Q#g0?U:c:QKL9e1<&d[
,^=^-Z-BX5^fg;MF,ZTfDPYeSY&9O:<Q@\9gXaeO6DKaZfA9#Z3:cHJgLTS_9(32
&K]Nd?3)d=,1TYC^FZ=7I[H\^Heg#NZ&^Pb7g:GV^4fK1>RR4]GR-3C.+?N0:.dV
6Of/@H-Z[DU8Y=e#N@E-)@I50I1=][BDAY^JQ3eP\Q?bf?7HIHHR]bM\__SgYY5Q
R6E&J.D.Q^,G>]W@R:gO>;I^QAML-N87E23PE)6>S8Zb.T,bP6NbR4<A=O0DL#eM
,7(>HZ]BIKN[&K4(+T0^1bc^Xeg=;57MX]K.cS-[+H]a5Z]J2RB).O1@YN3L@7f?
MJ=TWS]eYgJPFJ94?,\;=<c^bZH\EW)-7H0aNA:W/E(SFf,,[Xf42=9#?Qf>W^7A
JX0WgT?^bFM^YP=BH\;Rb30S:V\g\;)5Pg<Q7#^ce#a;5.#]]Uc]<^8,,aPU_/JY
0S,1)6;WM?:>A[d>U8KP/c2UgC^Oef)<b31c0fQ_11C\F-dMS98Y):-3GbFTEE]-
0:OBJFdLGK2S/U+5K4^U2Eg]A\b=9L#(b,MEEY53]O(W\a=)&f1JZL85.1?M0KBS
#QUC=\4P+/V?d;/[gCZ[=?+TBT6\EZ/C4SO18ZY8\^Tg-BR2W0cGVURH/4+ZC]c<
#4(=5][^/:BGgU1^gXL])AROT>?]/]XG.&W[D;^G?BOd3&]R-HZ@f<L@E18)7X_T
&4Q.DI/]&)PCVED-)Jc3a[YQ8,5]ZM=9,)UeUeg=LKH)A)&ERU/6;aAQ:&T94?MC
3K30=WJ=E1=a1+?/AN.040P2b>0a[1YR=4<G2aG(.PO>4AfR0Wg(^Q/PH[#;]]BU
7)cM^)3/##B3b=G]+Y?C8VJ2/JMZ?8A&ELDL7\<WK0<[<8X^a]gEVNQGDYK,+/2@
.I-S3#CYKPR=2a4R8ad-9G^+;GA@?(FE2@(S10XdP9>MfDFN&:/K0E=0g&^X,H(I
TLE,CHE+\M26-UfcW9DRQ9ISIg>39=,a3N(T)B-NbaZSWN+ZD(#MFa&AFSe:f=(B
RC2H7cMd5_V^;64N[dBT_JZ;fN#V0Ba.MYL51S)[J\X2Z5=P/(#>35TeESLXHXKC
_e@c4T1X768gUcY8g_QHDQ+11\M)K,RDP_K^QF/?^7L^[SW^&LX9a5;??VC;#+BZ
e+bcDda=89N0OM<U87@1ILd0#(F2O>=S/+[(46G:6B(eJAPC\;(VcM2e\CC.bHLO
XL:XN==IEL&#(S\984);797KB#JYec\1IP0=AMUW?L<FQ&YIM0.IZf\AV9?Z=JMe
N[Gd]@VRSIY\NW^/K22.2[gg-POG31^,>fZ@E--[fHH0PLZd4E=SMgS2GeVZd](B
cT(_B8Y2-,/VT=YACOe6@fPZ)40)S4XaF[@ETcP/CW5b:-A=EM)5TLPDF7D<Cb;C
(I[_c\0^GZ7))<Tbd)JMV;F.Y;6GeBf,)bHI2TUR:(KH7/1UL5-5AMCcNFO=Dag7
YaO0^E+YRAAE3Jf;BO7UVVEZL&Zcg.D(D7<07A17g(^?T;g:Tb:_=.+_VP(AG+-a
GB5T6g2::bUaEWO^[J27^2)eTfSWgX&G;MF5J4=TT?OY#9e)g>E#c#05?a,g,9(F
J)N-_KOT.5T.E,;GeS-<L+I2cVM)V\?QZMQ\_>1Lc2d+gD+=-g_Z<>;78>^:5c(H
&N:_Q0P(A]7C8K])35IUd5_?TUIP_?)NY[dNO1JKAM_CC)R^#\CFO2@5:/UJKIOV
F(+:9R/bT:(D^V80:<Z<=U#);&])SA)>FVT)H6T:,&VbWO=E5ZY5JPTe+HM\D=F+
V.3f4W?Kfa+B/I:AY#;f^,L:OT@H(AGg2X:.DZUO8IX.OcXIf(dRU)DIECUX>&a3
VALVGT4+=&K=ONbUeCa^NV+1>Z0NFU]=c^gGX]U.J)>E:(eGC+1X@f2KIDfN43FU
JJfI@OW9CaVE@;#F^/L_NeYPG#PO=aPOFU2G2M&.gMM,)V6?RBPY9PB=L5M?VAg;
>>=?dC\?0\PHEAFJfBS#:-75LX1PMK[aUS8W2&]</,1Y#]-,6:VMg]HX\RB2;dK)
CPg6V/5bN:FcTL#Te5a>L@dWK;)M7RQP5.IFf=N9HeaIN=R@Zed4EFIcQF/Va91e
QeB(A82&@SgQ;E(R((T@ecZQ,]Y^-4LTZ48J_PSa3&F0T&D.:+c^:FP&Q4<bEN=^
e;=/KVAWWO(IZD[ZGI5f7-0-K/I,,[Jc_;@OfTbUPd2+A.F>:5Z^B57^@/+&JGA>
T&^,/gR^L6FYEO]/<eLX/O0I;B(WA;NW<CHQ8:;=V&&A;&=XE?\,/M?B4\[10:ee
JRcW01RC3gd#^7(0)?0&A&ZLAZJB;M0bN[eA/Ae0J[Jb>[F#cGZ[7)b\OAU4-QDA
H[/]/g]\]=XUMH^>@IWLW1)F_a-<IeH,\=b8V67b4FS51JYF8e&a:d5.dAO^5ZG4
7DM]g9g_@@&<1]_CbeFH>FG?UF/Y\#7.QK?NF[ZUB,7f3.#<f7^UPgcA;&X9d=CZ
_g#@Hg,LKd]G1g,g4?4ZV9>EW47\_5VDM:#3#T4@Z8TV],H=T)3_;[PX?@.BMKJ(
CNU-^-V5\U8G:22K^W&eDJP9CDMgJcO4<,LDL+6T/JS9:\3U0B/3Y?=Y4f[L?ZCZ
U[L/MV,>KM.D@A:2W;0K39BD<3/PFS11N@1ACJ>4(H(LGE+E_d^[@Mac1H4:N;1#
FF3-HSB96<ee6Q&E.,4bQEUX2;A,08bGSOg^.E9EDI31ZYSabfUDW6A:NOO7IT]4
g8MIAX+]1F@LL7XJN;UH.UdEg6D;5MKU\(9SMA(>[[OeYfb0,[CXg-f3GN3XUXOV
,ONPJ:eQ[S)(/N@J:;[8g:-dVI4(PF+R6a=.H@U-7MI\DQQP;VbUY+)Se2W+J)BY
&:\DGe,F\Da@)=GG/Bg+8JT.3Y9NOJN.]/NM=\^V5HgG+POW68cXWUIbZER;4)CX
F?BW/&2-]P[V_BX;8TK99IEeg[2g_4X#REd,YY@7BTCJZ]J>g^XM5K62]64_&gSg
Sg7(SI#U^7,?ce=_f.b3-B9#=gA9BY@B4OT&V>.IOQ_Za/.OU6UE9,^0AabV61:V
2DY4HbRNR.@L>;b6&<&NG<0.+#__?>-;=44^;C&@4M48LRL_P+d.]A\F+KMd_C@]
SPf_Y-T;6FEK3=:PU&X[721+8UW8-_MfeW6SYV0W&FQ0]#&WA&.Uf:0A2VNc_)6F
PLH.#9J(fJXN]3W@V?H)e45;7;#PM.=78X)TK^4OcN>=E(L7Q#:LU_(N>ZN9Q97T
C<]UH84MJ/7#b2Xc_e5c+T>S1VS0.g2\GX1@K1f@YD3Q@R];T&:Q#(CP2d^BUU]E
4;^ag,4bA?PYR1aZ&UcET=6?3C,B02B-F65,=4M&WVHCKL;#8#Q)F3Bb.I/QVRf:
Z:_XZMK_XY@5+?(,J3eHLP@RLD<-?]34>]V:]1JfUf1cg7)9/Y2\]5d)U9D1Z^eS
#=DCY.Pg-fPT6dUZJW;#=F9+8PgC<W4D8K.GbORU<;:QE(9C=ZEN>53aATIKRdK5
,b.0A><O<+\=W[G9(.MdfKCS55]-@Lg8We[d&+XLY&L,TIQNfRdKDD#QVFfV=2T=
)93C5-V(UTQVX..WMf<^K2Lce^_;5&MMd<(ZKQ:VZ/PI7YYI&.>?ZE>RF;=9V]5Q
_/RLe\gRZKUC&RA,0)W9W_ZI9d^G&Q_=G2B;+^^BC]M:COLP2g,?^.;4=?c9<^;e
VEYc16DN=7A;F6>P^@PC\PTNLP-3.PSUOCHE9fLT:.J&b#JYP=B\=X&(N8L8>E>@
#5/L5:bP#&7bf+WcXDF9S\][/CB_3XGV,\aOfgR70089V>1^M-N7J7B)_/O[H8)=
AcA[Gf;AQDJVeMM-,9S1P8L]ESfaWgJ9Q9<QBNW[0B(/2>ZK:;)U#LS7[1d3V.Ad
d-J,_Ie/6H?BL\+5_;X:32FC.SJ?Y)d96Hcd>PH.03?\B]e2\8b.UCGP@Y-6/S2L
(OC04e-F_a4[G&f>cQ9&6Z8D)+cW:d&2,fL\?6N_N5aTNdV6OF,;^OfMV.>,F.[5
2#&UGA(B67[IKLdUOb+1OBc<[5TB^MO8P3J<Q:)eLWEV,4Ke/&b#G&(CS<eN\H8_
NgP:+&+8?S0)NbH^@JIMS1FH(2MDW3FEG2cZa4=[T-g#fT\SbOM_3g32R.KIMOKA
:RWgNR;3S^Q;0>K0Z314Z21ZbIQZW1SAKfC/GN)IR&\ZG2V[e8,9BT=L9OK4/g55
TI>;GBR<ILIaA;V]<)JZ9Z8JNH0QZ-Z8IY-59fU;]>/VQLGTTa?ceI2TVEI?C,[#
=(YJCIC(#_T.U/[LS4_IP<WSNg=Id17:#g/5f2<EFA]SV5NZeXZG?:a&B])?J/c#
A(\4&G=\@Q<B--ZLaT-D)@Z_:fM,JCT@8+6PA)GgK]+[&,A>Tab0.OUGO7-4JM</
[J\H.(5VaTFgEKI0P++D.A]KNUO<23g(J&f).GGO4QQB:.ddM6D-0X4f&DM>.EA[
0+.If2JI&NePJO,,I1QH40QY[20V&9gN6<a0[dAKSBV3bNJ.IC9dIBUb0?-c(]O[
Z;(KePc;c3IBZCDOZ#SE8=V/4WM6U1P=0RJVVPGM;a,)/4c)d<+#NUc0BK=6_^^@
a?Z405:ce<CLR-Q[&Ka@D4XJNN;a^V2O);MPIJfEJ-1G?d7S=3@@R<^H>.R\U_X>
DcWc#cDLTY/6K\OE@S8fT3+J)5J;]/.3<WLW75aJb-.75>?R>Q)1/bT(\;H]HMU#
@8J0ff>80b##M3EFMf9aa7ZH/;25G6K^12]0HaLMa).Ea81@U=P343WY^R7f5#RK
3OD7Zc]Q<C]Z..OG:X7E(B;SJ@9IGOJ:SQ\4#&K:g58Lg:?2)2R<UPQ7^7gI#).8
Ac5XK:b\:I&(DcNXQ@U/[55aP<(L_4@-)84dCKAH;FU.-HGEM_Kb8D.NXCdg^[&6
_81J]KI7dXLg6MK/P+C3d5&QEFA:G+G,Z:<\DR.5P0;C/A]78W>^_4EQ&)gN5AY8
QP5Q\-D+@\V(c_5cPcU6<:UW0?:D\2HIJ./<79Pg#a\D&/OO@39-\#0RSMHeXQg7
F;UgfYH/U3g/H:^&)OG]3UWG]e0#cF\BLeK@1JW+L7-#?2NE^ZEZHR@PIM-&]<eA
G&P?=S6K8:W+Lf369,XcRLX#<FG2S;bJGDN3<f:7L:G)[RYPdd(EQMC>U;Z8f-]T
Ke5(K-_FHXR-c\);+4?_f21<Ec;7;GRFI@eRLXIFK_Q.bSH<8I,]#^>a>Pgc71RJ
T6RbHVd:3+?,#8DCA9Sa9gQEaH#-.I5M)/:<Vg]I<Eg1\FP2W6X/_;-6-C.?:6)g
(9ZKPHL.A:<eR;9@G=S>g^#&&7+2.<8Ed64XY]:R+=[bbOWD4IeQQUURY3fd=8Mg
cTScCHEdJT]G66E23]RML&[>NFd^;XG8V?/.LX-</S6?+NSN1FDMR>Y^EeX@F0NM
YR[.[2NaAPOHVPHC1.dg_6X6_+R>\;g/X&eH:MTMTE&GXd9=Z<)CfM=F@?1#-3GR
#P@gUWS1+1W\]>OSaZPWORc\4##@?#N04WADb1?Nc42MMWT22fSR<Fcb]WDH3W1B
_NB\)+Sc<93SWTc0V@OTHcNZW(R]T)[#K(]bXY^&UW<0O<&G<,Y-T]HM3W8K.W,0
,b2ONBD[FaVZUMd87VC#,39AX?O?0XbbLA[4&>U6+0Q#D]TV1e4PE9g7]<O>[Y)#
&O;^N7]TXa8AB58_:^1GA0Fe:2^1JFL>C,?BLW4O]QT<F5aBTI(,M@CfZTP8KHc2
dIYTX-5B+6@Qd@M@=S0F64L6<85N3:/J9MK-cV9AG/)d8X/L^QZHaW3H;0^([X]8
Z+.Wd3V6F7T/W3RCNI4fPO?A,+6)GX<,DWK7)L)@(\0?R@P\fJ:[NA[<].8+6)2b
B2?@,d1N3ONdI<D6ST.T\bRX=>2PPK\8<N3L+G7W68.F1TaFXS0S8)R&\Q])]OA9
GL8T9UIJ?5-<9Q^E9\bNe^NfO-gcfT#52F.@DAL93<;+4AcZT2aR@=@3OE3L\<9Q
KSaS7O9df+B[ZD;aGfT9?D5\8SP1KO9YGL8e:BEGB\(a@4G^KZB5W:2Y\&MWb.A1
72TIX;=eaRcNV6EF=I7</>bU[<)W@>1aB7.]DcB9BBZ]/]4?P6GXU6\E37/?#P[)
IFM>gNT49a,DIGSMa<3LR@A89fNKaADXFDMM[4OcR&/R+FI^LM.1H0D2X;NU=4([
W_=S_U>->ONZ86MHR=)7MDW1(ESJ#fF;G@XWdUF&YeE_Id2PI_0F\[=a_.dP7A^[
67Z?]6E9^WWgEF@K<R2-_gg13)+I,M8QHE#+X6VZC;W1NeeP.-U]XTR>K2_:+=\R
I.fb<@HLO#G5]C>,[GR[SM9XQ?)XJJ;P0_CG.D9_VE;VH>8W013M)&a,faSIZ3M]
4;./XQBLS4-3YU#1<8V)T-0UD/26B+Se5Db?\\c<S#V=N\&Z5R42[7T<G7->?DE_
(gYdQ>eg5DcMOW>HO45AR.5)/dJKUeX#?I)XZPM0DXT(98^eYRJTBW;0\Bg+@S].
/J?W@]S[)[Yf@#@Q/+9g#7LI_RI,EZRD87fE:BD8L(HFL2dW+G(eH]T37GCIFE>A
;ZN/?DBb\.bS&_@TQ3^[UPJ]07V4?XG7cN3>?E>@>(\?9D6>&DRB=+9NC?G22T55
;(O&0,dA3O8e[P?,WN6e5(2;1MBIJ6KI7c=J_N[<^TIg&MJ3U[0J2MQA<S5GR4Yc
:dK)cb6P9/JQ+;I\3YX(BNE8(97_K#1FV7KT5SNIY+4\8Y+AZQQ6<f2)8(#?-=BE
.39XK?]):^JQ@:5gX>_99Ygc?H^:\E.]:cL82/X?+CLAK@MZ26AQ-K1cV+<638P7
-S99;6(B-Ac;_V-OO\[SL5I:<R?9-cQF7T&M-_WB:+#VYfR#S^44aFYUW^?M18ZK
?>57E&gMV[&/XE7cZY033C(7SLE\>H@e5&2U1fPA13SJUHBF]BG9Md^_H)2U#]&Q
]YO9SDX4^5S(:0+REIFHR@-([I]#B5CFPAb<BNJ;1cK=LFM;aUa]O(\B59d(,37K
HEY8cR(:_b5ZB^_UB.1<Q@&79>aQN,>EgIT0W#d17a[&1+^@.-FM]C6@6+:1,PK#
92H-4bJH7gbPa1a2LTIGE(e&NKQX&NJX[0#E@B<I6Lg^LgS[g6+-E6/^+1XRUYY>
;[FL35V2IE8c\]d(-c#O8D]18b+YF4VdDdDd-K@Ma2:IKFA^]If9)WDYL1Q#VdDP
J9V^/ZT/(RR]SH7cN?1&>92BKb))B.)\?&4[&FLb6Vf0[/925<AA?C^dE/?^CJ[L
b@fL<fZKZPRE4/WJIY]R#&68-U5?Ed=F=6dJ.NWBE6K=_Z13[??U]M(8,IW_80I=
Cfe957/-6J?e(;g@c0TDc4/2S,MYQ[P(P_MR:Z[;Y7_[[IWLS2II@8fQJ&(/E,GQ
d?X16AW=X^]2Tf\JJ?3K0\W]\+E=4)FIWW()NNMdd^TGNS-8#bR.M\6N;-D1JNS)
#19-dN-D8/M>(AZUO5I;fILRAO;TZHXVGNM+Q+RS@OaB.(A3d?bB/2F;]G[PD8JE
JR>PeX;4.bU2G2,7b.U.9f><3U\,6,O(RPJVZ7?-8?>O]MK;YS\G#_\R_d18HNQ#
S](:V<DL)E@-^bLf/E/Pg6D>#AcC8S0MQHQGe-f7=+.T=BLBXS]Fd+QMH/;@,Ig-
2JHCb9=&3^MfG6HH=)?4:CaB_/F;BJP7SLO\L>G@]TbgTBSUTf\RBZF28WI0XDS3
#3ba3B&=b[+6M@0EJQG24Zg+;#Z0g^O:&Q]W>\;LXS9R1RD8=S6ggY&3VNT.9NQ2
GR#NeHGYdX>gIf&IT7Ha7IQ#_(3CMB3b;OKg>[R@a8@)PWLe6a7XZ;bX9;KC2\-V
&Y05([\L@BVP3.GAbPgVc.V(@F9C<.L?8^C,)]dG1J0UfG3HgK=ZO-@g5#J:#AB>
eRD(&KF(^O\80&#&P^0#9YP,Y_VJ=6DCcCIN/)LDJY^GWAG]LfO0bN]755E4-QJ5
?[)>](6@<d/G[OAA1W(K^d10fb^D..f@-d@\IN89VaXQ9.baQR/;7Eg++QJ8)Ha7
2X&<MS,1WDf_#(W1?_3S8-H(=B5+58VAPSL-b]bT\;b\/1]34(KaG@80M<[=7ZQe
d]NG<V4,3U0LBbW06gC\<>2K^<+^.TIC,(UR1Xa5)MV1>)K1@YC+=:X\8PcS&f?J
2;>#6@DLS_0E>R34<,&AO+,4(NAdAOD\;[>H^e)_.8[]V\@2>0FUTL@NAbAdD3@2
N,e6R_bHdg\(;_BY^.T=<#\HI#7U^#,OKE<YN3MfDAO(><K#3RL;-1a&cdU+N7##
6.]O-;]^8/DO5V;=/<[.BG@JE?XBOU1>\(N=<8XRa08Z#,6L<2>e+46S(-VQX,^#
9^C^ZR,\@2PcR?IL#IH?SNJ\1CgB@X:>7bH8\N3\NVY@M(.A1BW8#1/ZFO44Z49U
gI,C+UW6aScJBKXDLEUY@Cad7_?H=1bgZ--?\c_9LcT\->;e:T6,.V&>8g)O<<BT
C8#9W)/T]=HJN^##M_71M2a:Wf9eU&)+[AZ[/W75U>A?FD1(L>;,&=O(7Q=6(DBR
2d&>NO__(RI<V.g#HT3D(.?:).]6S6;3>.P2^4(\a4JT\[HB3E2T,QR)N&7g+d.6
gVBHQD36@],9Z-U=b.D84cQ#&N1C4E31]R5(UC7UbL2a;2Pg;UL574Mf\9_.TIP\
QKcU^RY#9gR:HVbMF+dFN/AH^M.Tb5R#7AagD[.b=66V#?5.(63(W3b;=VVWR(Q:
F5NC1^d1N5eF(]AJF5=X_(b>5?)EbVC+@.2L1AHdggD-8dKL&PM)+L4/9cKDW?<D
&9NbQ[GT1_-3U[XWcge3NT=A_(W&E<CWG88@e<29dC2c.BJ=#Z6eXC?a99Ze,7QK
V;&.^5YdUCDeK9.XJ-TK-O#__5[1LJ\[HbUS>C(S86fb).AG,:HJ<;MDWKgUUcc5
U=)RY^e1T@TX-MA;/=(H]EXYIV,))NP\3CK#\.3X=N5g-JB+aZ^G0X=648,&d+DT
[9104WN(NM@CRDCC];A8@80?)H08:?B5TQLE7;T7WbXM[TUQ<:fYK?(gb1?6GVB>
](aLLFM\-I<+RbZ<gVC3QQa9^RTO+^9=acUP[06,(ULWgSV>\/B,(EA1EbQL)I[?
3>=RFC6a+Ja5V2Y0]&69=&RZB?U(+(P,I&@P(G=f[XM;38ac]XZ_&9+#RE&&]G0N
;A;.#/bSNN<)#[P,=U+_8=-JKcc&@EE9e6cT46HOZa:PSgX=O)FY#NUcWda\4=3R
AX-[B_CBC.+0TW;\Z]ITaKTBBf76=81<aY]NWB9WUeQd-^BMN+TBSGA+c5J)>LMf
,W9E\2O[1H&3GCf&:[&a#dJ?>44:cP1]QOA:Fa:K5:g3gGMf0T/8RHD99(.Ze-1Y
0FUY;,aa#R21-7N0B]I1XJW3Q]+[A6FLL_DKZY4>ME^MUF:b\3^Z,U4WM(D?Q2PW
7PZ=41B4G2]O&U+]I)C#Z3XSb7\X1(YbT+D&+?SRBDAH3\5dPCJ8KgTd3BHE2Ud?
+S&Z0>+C+]G7[Y^^0\+f2Lef\ESCH4KUF:B1AR_@9_:7^VC(gSR&+_2H-2_E&,@L
e0-G:@Hg/+B#^@49#+a6/?I]:76P4]:L:c?TSUbX]4N.0/0B03=^0L1=X:=<Eg-7
QV(IfV^-A3gDZ)&L.FQ.[D=Y<W3e0Aa5SWX#.Y<\U9\@&EfJ44-9dC?&Tb,VYX94
T_6(>PC,JVYaaPKN<#D.@C+g\bM2gE)SE8,4C+&SF\DX#<&#Z^>#QO^cCf5:BXQE
b1=YESO)T^UEF,_\.1PVH@eLL2RRYKV+5,DX99f=Fc29H,d\7A\PMNQ^UT9Vg3Nd
</@YB8.DV2Q9e@PQ[gO&96(VV(4?#&B[)YP_,^#:Hc>/^51=e;4Bf-K,QaPgQ27,
8d,<R>:g@IQ?RD?S>2Gee9a3Y-J3,b><&>+@JS3Q0gE(]H+JfJ@N5L[P5gWQTI^X
&e7<I9LQ?>LY6LYXRMJQPETR\4QJ-SMg)>0g,MSf]d\>X<LL.Cc<Ba==dd<,K28O
VcSfI(\Y&B,_9#T&UC5_Q&8e600EfAQO0<1IXfCZcE1DBI@[J)e=.2@)bY>09\D#
T63T16cS3JZQ<:P#L00U_Y^2N9;]fLR\7WOS^0VU_-,:TR9F-Z91:S=2YfJa1/>3
QI-1f/U^W92LPRQA8,0SN9XJX;NK.CSdbS.9G4QHFM:MTc#0DOW:1-B6037II&@X
;g6&V5N#bEc:-b?g8a2-E8YY1K\R@EI1+MRS-A1<Qg/=6(^/(Se_(0g0Bd@DAQS>
5e8f:R\?-VT^0d=I=5(XR=/X)cP(b>;I0dE/E.2PQ#3=Z#5b_G^U#aGgXES-&(=-
.X5KY+15:fWG&c_NHE_02g5-J(S:6CW@(,XUUdFKfR9,SU5O\AKQ[Qcg9BT[@M.1
3?S<T;:fH4I;1]KY#9#.EE&5<&-@#OF_4/_e5O]bH9K]:J9YVaRL3a&07L+Wc>R(
,&(O8e@KCU>:bUf/Z8L,)^#_^N)?[4)dKT4[(KAIUC=YW@TLP2MRN?c+8a[WDHQP
\YK(W)J^G1ffa>dIA^K>28EF,8D[2gI,E/dG^.KF/Ma?6K0/3#GfaZD06S-eW8f?
bS4<()XXIF.;_H79)-UY.,;3a/_da@36bS?QbP7Z(S#eWaB7bD-Q?K_?R+#[IH-,
<LV</246?B&OH-XGXf#U&OM?cP&<bP2:HC]IOP?7Wgb,?3,)ITKF/b6\;HW&_f92
RL<&QR:VSF_KUSNR8]_aT0Y/B4QZ?WMT-4SJQYbPC&XA7<V@6#QL:Daa=HZRB0=W
7IGaU6I7beXYB_#b4._YUGG.PVSJSFecLHFg-O+@L:@<\\9,V:ZZ-KY?Q\]Q5Ha,
F,OJ2[3&g?::eC)3Q7KZQDB,&d_J/C[;b.1<ALX0OAS0>NYD]@c=Z2-,I=e(X\QI
,TJ-c.2DS^fZ]Jd1dO=?\CedZG15+:/V4B4Gb,&6Ra_[_)MP)HX0cF6:X(]BfHU\
\VJ^gd>Z+AP29#]f@QLYd8XL.@T=7J1Vf8,DXb8;8NXEF131Z:\c,?(LS,ObN9Bf
1,/0\V9JW8I8fL=/@JV213[-W(+B.9A,<(>#Vd4=,a(/SPTNeD]f8>M8>@g=g&/1
BI18QAf,J:T1R)ZNe[7:>B^;;/J./59E54RFGWR\AR06N286H]BL_/b)=WNHWR>)
_>;V7X]NF0UdLWITRNGTB]91\A4<A>L7a=g_HPV7EXXI4J1MU6)?O,)bMf0W1V,g
MB<@1TTF]a:7C5_4L/-;X+)7P&)Sa>a:B0>+AKaL3\,Nb-R]6ec.L,-EDN<]@@8Y
_dK,<2>J,B-Ib40aY75IgVN-?7DW46U2cO(&]&B;8K<,A953b>XQHIZOIe\-YSUL
cV-]>1XIFXRRK]_,dE^e?FIHA23c##&bbf4dYM#MEB)M/C\5J36JNH/(Y:WOR]5I
d3Pg5\8&?I_@^=cHB\R/TXK.e8R:<8Ca68UVCaf7A@:4J_RgC@3fDZS@T83[7J#_
M&^9g6IX#+GD+dcP;W1g5SY]UBEB.EYUXGNR(BKQHd4eMdFPb\LC,@H6B(I/CWA2
._&90#a?38c]:b7..9CcR7>,6&DZQGa(0_Bg9bY_GbRD]J/>A)AYRD1c,S:1aY9C
NR_MW2U/66:41Pe0:?50UO8T6,:N=906=\DI24YKH9(fH+1A6?1\(eO0?3(#0NA7
7H3]d@7EAQF]:9D:1IX&)M&^<NP1]XN+eYR=8Q]@Ba<CGO:<8/3#5G)[C:F:Vf,1
2R4B<e[JQ.+@R<:\O[bF9X(TIP>??2Jd-AJ^KJ6GA>b55O&e)B+JZDS:=ZV)K#B&
;^[/BN.a3ACb#fe+;FB.]R(a>.C.M?f/fD37E1P/-ecdXDBTY2L8T882S#&4FYcg
ALgSX6VB;QDO&YPgc[1^TZ/(IA55WBV<df/)#9V,BSUH8DdMR17fO6:CK:W@I6QH
HUS[6KGJ,bT2Gc+^&EaSN(6,Q.g@.d/I?Z<,XL7+1?d^Te#_0::YUGfaJLT7?S&f
<MEdOL=O4D]#Zc<K+c99WV+5-\][^D^?JaeJgS?KHdKQ_:6F9.6G9Ef,dQ^4X^NY
5d7TCL-;-C^dZPNCH8]J6\;88)E8ZE8:+@;gNNX@db-&?L5C8K<3-H]@STaTD>VV
Q6IP7>GI(#39abO\@J?_<)]UN6N8f&2dE<Y4WGOXd:F&cPVeFX;5DG_+HF\L04DW
Ve1fP2CZ+OP<@C@-_K74E9W59cb?T<XVg)E02[Dba#-\;gSK@bbJbGgE\U(&,.Q9
7gP=f1;8-MR61E.(L<8K>Vd6<K32=Kg>(;(2e@&V-AEe[e\SBL:^DV4^9WZ)\204
0?Z?7MdSWEV\(2)]5\R?T1-@HN>]fWA1G<BAMU_VZ8P0VTIX.2R/.1WNM[V6OF)0
?C/Qe/[eac.A/?=cY_7@HdOS+c-Ra_(eZ=,d8Rf4-HI,6HKeE0;^.H9\VF3f.#5+
.844#FE+7[N4K,=UaF).)?/#POXBD(7,AO-A&(3;,;9AefGg3_5b\DfRIGa)O0Pf
>^0FT4P+=(-XDN:QP8FCVA>U:ZbcI<\K/bR>I=XGHe#bfFD\-(@021UE:;@=E-OB
P1D6R3TD0MG1J0N;>#\:-G>]1gCL4d5-X^e2F^3V@G0]V?Ye,IJcPR#-9JGEK&GT
<&e)V))/LWA2Y&ISP<eJadD^CJQg5LT(JBC]GDS8J7-e@DZ-[SXIZ[-J9=#LU+0/
,._QBK<7JC^A<Q^04+fF^;b16DBeA_0Y4B&O^cR^B&6Td::R?1BMcV2S]\B.4&D7
7#D6:A9Q&B.^IeSf94PFCb[=]QN\43A<HU#cFWW)@>)33C&cSGA6,;b:<,F,TA()
\-=+EZ3C/^B&E&B3Z@NQf/abL,3-R8FM+RLaYX?35U6>@APJ5&^\AH+E6:/Q(U3^
[PSRA3+XPAAbXFgbA2/WK]e@<>Ug@=<=>8J(dF3G194BJR,54;a4L4AVY89#c-1]
Sg;9ET&#I=)BgNOHM0B6)g,4,F-ZQPfRLQb,),gC;RJN(8R(UI#c8\ZI&57>H<8R
I3eI-FS4V+T@G0f(HOVXEYfCf<.&6MZe[XIB2[VW:,b6Z(4;\>Pb\)8C;>g/ARUW
O(+]E6Z75<N8)#976fYRF(eWH6<8cJBL>7Dg>]717[X^3@DI:B0VE)<>/81&U6@V
FS1bTQC+SG=\:_d:-F109S(0](LIY-VO;DO0F@0J>5OI7GXA3DW6VIdIZ&X??DPg
\@-ZZ01IBV)f&3<6\SdOaHOg^,NEHOB>eNR)MgI0](>gWcgc0F:Y-3ALeA[EIYK-
NT)I&:,Zg(Ld\NQ29NWbOgMY\EHbRJO3DU0=(ScD.a8dD8P2c3#F-IP=(MS5YfN&
X>\cXa0OTFX>PZ5R6WH@,13eE)_W#)A4J:;U1YBI6##bU(8CdFH.<9bC-W;e3(&G
dXM?F75;=.=<cI27AG+B+QgIV;T991C\K;.WNYMc1=1+ePS5-gb-FMRM9.]5WT8g
B9fTY:Z:,b22]>Pf7:3:T8WBJHZ)WI,WEDNYNKYb+05TTNKe(=[I&<Xb1f-X2+9b
#b6YE5f=_baMH2:VEY3H>7OS0f/&,O2B]g^HN,P?R98D)O>^V]4^E.E98V1Z=?3c
=LZ+Ic#eI_2S@V?/+5+O0JJKJd#:W1S&O(S&bA[/.=?_a)R<MGf:__-gX-.+/H7:
SdG0(>P8LOeE+,ZERFTH70Y-8a2CY;Aa^I9P-eB30?eJ.UK-MfHf6LdZ4;O3+\+&
E:+]5LO,]c16IO4>1E0>d8.cT59(_L>K]5Z4\//U@JBM,?4]X\NHc(4U4#1_La=Z
@G8fRO/-.;1RB9M&CNd7(R.f&4X5JY+@GK=/c9bVFZ.4Y8VFf(-V.5#9P@+SdB/#
2XAPCQ18LcEL@Q\bZ);:/3PPGXf54R1)C39d3]9)#(G1N)JUGN4S)=:HUa2P1A[E
eEHb?V8<>YgQ4I[W]F)?SB]Ef&e3UTA7D[>LVJ.W+I0dOWLDa5@SH_Pd.PJG^1@3
(YZ(<+&BECg[1,S+J<Cb[YD.BCYDZf;bIOB#1.H_U)R)_NA_f9#aC;&4X<RRI1_/
LLWLQC<HI0&,b;C)=7g0AS_07Y:&<G9ZO7f4KS5K#B-01:a<fC;0Uf=<D?<9P&OH
,YJ^2EMQ(?IHLT28&^<H1@FB@K<#<#X]=aOfA7g))MC2-;:Wfe6=VFG(+YHB_&K]
2e6bH&DXY7L0K&/M=bg=^;/0Y<84bBL]QL0-g6eF1bV6dE&N;M_XYH_FgSO-7-]c
#c8N\66gPQ>d6IBHHUP?1QT0=6U<MRA)CgGR3#D2)912[CfHYE8<##O#1J?GdJVS
8FHGDJdQG3QI>:@K=S]_Te4fH4H7c?QCX2SaJ-LM+#OB>_1\ZeZgaL9BE?_6^>ZV
JDJ]c+P(eZOB1V:a0GB;XMZaFT,9<aLDafY2)S[5EYH\<:_ccRC+_7R(<W_eY9d=
CQ#JN\LHB1fT+Oa)5<LY9\We.;cXSH(P#6f,GUbZ=@LI7bTV?9Z<X[,2&3W8;&18
&Q01>cW8PRa3T+Q<dG6WcQ3KZZ@RKATYU26]773VIY/TC)]]UUAYLM[0;Y+eC\E=
aP@274Y0O3W[20V8V+Z9T&IS3b:g79,7I:CcdB7DgbE\Mc9^R=HI[8=#RYV5LKD;
g\Y1](-G@(([B.9]AP@cL]Z_6dXM_(65:Hf3dd;EaR,#e3^>)Z5;7KMbRfced6DN
bT2#.Y8XB7^Z1geC;:Q.D#8YZTI+0,f;PRJUZV0Ae[SND06J,=g2R[/AD@4T9+]Q
(INa]EE0)KALJRCA8+\=F,1NJ-YY9(D;X-4>-=-^_YHF;-@L4T<f7XY7<LbMf_J;
J_])140R6OV8H_-d6XN&9^K]W89B2YB]fL[\QT:F@3]<.?Z_W6dF,PcK0)+48\LZ
HgACc2X]GX#_8[OVVXD1V=L\^&J,].D65]G3ZZ/c;g[S9A@V5OYZfE^Q2-,O3A+S
IDQHO#&[P4?BQV&=CRXO2R3CES?TY6^R#;.DVXVEUYT?Vc&EbWJE12e5A2Q@T/Z?
8A5@9e/]fB2?B#1/4BTc_AETWO^>/60Cf,(.4+V>?V#VJY<aCAF;0HV^+Sd9N3gZ
>aZNA.SE&SJ[-=c/?;HYS;GS5\FCS8d?U]X#RCK?YWIfQ/TKK(XY?^CSB(T>L?Gf
Z-AdE=f.Q_A^eKIJEX?L<T62b?^:4S3/G<c?GN)g9Z&MA]:@@B,XZO<,/0E?0=;5
[,RGBa,-XT>OF)@efB^E?,FO)D-BGd6agIJ;FI+391c2B^<[00ReFD3]@XBY^Q35
,H7Df5aIE(;6/;#U+b9?a_S[L]E_76P,-g03HGA>(0;/;_N8L+MeYEH;MT>H/+NP
RdP4?e.#MJYM.f>VgC00>g6,<U8&.eL1b>YFY^8IP2P=V7,?^A,HFJc(QU>4P.,,
JL,1bJ/RF;D-g05+T\@]9--M5LcRDMc)@YDWJ4NV-BE7G89Q)0RX5PQK_R&LCb7c
BWMKYX)DU;5c1d<0_ZAU-1QQQ>W6=Y+7IX29TDB:OOGP?F=Id:bg@FR)Hc_eRZR7
PffW)<>I.f;NW),&KPJ&VJ]STI3(F1WB5+S.FMBBbGS)6#K?XZE1fc,<MaY:G=^[
g]6X);E7M^_QI4=@-JVN5E=\3P5V-TY5L#;a6KB^B:Q+,ICcGUJ;aPWgJKHMB1V1
C)cST3W&g&^B;E9)FOK0+?6SR3c>880)&^;&W/HJTN,.:_=7;[<N#JeN@42DC34T
];^E4PI@aYXgKGSU]1.CA:8RRMTW[Ca;BW^7-0-AOfDGBMWcU.6#G.ED5c98STSI
18CE/M#5Oa64STG5(bRc:AAAF?,fTV8>5@1V@IH=3QON;[(00EDad3UadF]5<X^;
IN4W?(HSR#0YIHH6L8Z=-6[SZ#EWScbF]4.F<1cUD<<\.=EL^&Q3b:EF39H@Z\K0
OHLQ/IW/1,=E_-\1LH5LI([Q&RbVY@P>Q=M,aFJ60)=8.?M,@<-UHW:BKQ^NB:,/
;M_:]U48;>[L7/?B0_C<Fga96T;f@\[3@?\\>Y<g7JbA1ZQ(2b\[&a0,@4-F\4@E
.dKA)E.XA_d)E)>d<gfW8MCN3G,.I66#(=S)U@W@DTXGY,BS_Y+7]K&:^V9GV];3
085f=_.0B)F,7<7c=L]K38;TW^[S[FAY5X\VYcASQH\70a5Y9:.?c8_Bb.X=e\.<
AgDFDMKg&CV.P)+C-@_[0SLK=>U61OG70CX-1\VGb\R()CN5Lb#LaHN]EcT?YO\,
d>;?]#NI<gfAIN6I/C)eUKZ3\BYaR6g^6R1bf9_>>;?820Ce&<)4)E2(K8SDNN7Y
\UaV[+I@+?V:b2^N(:MHeJ[Od]>U;TC)c7#?N\<8_)aXG_[F:7ITA);ODbE-_MOM
=I@T]cS59J_7;GD)Eb&-74LVZ@7E:4O<_fb#4,Y9#^G+CZ/1J4[CgAN\V(;>K=/6
EGa4d3V+:177A:_T-W>W;gY_IXLK]/Ce-?P?[)F>W3V:N2CJ.+97S&Q1Q^98RcEf
5M\g/,U+Q4K(9QG3^fNY9YV0+dC4A9gd/dKMPb/F.#T1(3-\]X_D]C\IT9XS<:/)
e8VbR7^9bM2]c:/?FCfSZ=La<Od8DHB4^-VDEU266AJ_H&+U&H=9NK283g=60FL_
H4DR8FZX@;0#<MVM/+71A)L(1:NT6\3g@7QH&,2?^:C]:3SXcc>MPD&\;+_BdURD
@[O,F[+VM9(SYN-8[aHQe[eX7\b@X#YGZOT82-X.\faU&a1IE)[>_<:6B:G7+-GI
/U:D6f\G1Wg)5I.2YX@:#IY0MHdOIUHSe;D/8+[Tecc-A.M.19CcT3.c@-5@QPLW
,,9-NP]V/=+?PI9_7RU]OYgY+-POb/1W?g3fYX]O80Y?:JK?M5(;U1HG=(E0K/<7
>=NB8PEQW0SN,U.&Xd[H[9FC@b+0KFR(b,/H6J6CL.W7\20([^O^f:+dC[97YO;_
=bdJ=FfD1g0,5[aaFWNf>f]0De\e0LF^g:aFH^=U8c=>N1I<RU?dTYO&QZGK>CII
F^HM;6[U)f\/bd]7_ga2==;4[D)HARd\e(7RKLAaXX3M5>,9LK7cQ[O6?&B@BVHB
PX\.BcS^J,5EO=KHL1@UYA<^cR;R(29R.LK_;3H=)0-R+;NKP,;GB8C9I#RgBMH<
NfaPV./XDECV=UZ[HZPgSDb8]K+YN5>LP;Td=NBFf@1LV=Y?(.Og759U5[Q=HOB(
@V/G,0LTSV1NZG?5f3YX>>I6U>3PYJ;)Bc5bXGYFa/e6+PZ/2W1GYgN;B.R)FGTQ
c1G&,_=X+G+cPSgB7&,=+__[QBS+0<g[adcdbRH.(F,KD/:O/GcAEb=b\XG+:d#F
@]V&If4gFXX+BA(gUT9NVDNLBTST\VBOL/2[f;R;D?R&[@2)YedJC(SSONLMZfFd
FY(c?]3BB73;[1\E.8@0=eZaAMb+(;4ZW>@LI9<,#>L5CS?\V,;D1VT^F@eZMFV6
(NE&27>^6I??D].JBEfU,.fc0OQV:)1#RG([0DK22#\FJQ.ZF>TbOC\G@aFda4aN
U76^HJS9PZdX:gA:ZAPRT9>;+QZ1YE5^KYaJZ8;bLIJB9Z:,?_^UQ.Nc?N\\@Vc[
6Ma>/)HI-GCY0V5QR/95cI&@6]J.f=C9#=^P/6f/6Oc7D80b,7^19ZL]P6:.2U.+
eFg8HSPQeTO(ALTSA9D::6&[>O2GY0;[&Y)dX#M(D54SO(b#S&>2W8MZ<:IM_GRJ
TJ[H:PFRX/\E:-(BUCKTa=fL)I>AKdaUU-3-3ULOP.QOGU0:O4aOgG4dU]8L)E\8
?Q+De_D&g\.IMW+>.dK2+?e-0(N4[<;2&R+FL/;<\Qb#0;^K??.>R815AC6?42@:
I+HVfR/NC;:5Ua<+G+2c=_NfF.Scg;b>bU^^2+CZ)D:(QZ>46DA4&;D]A8[K>))/
6^D-B52gREQ1O8gA.;#ISfe/b0,OP(a9)5]FHI5J@V[7IH?-GOSC\AN]e&b8(^]5
--,#6fXbX:0JaW&<@a-[MYFaD[.99AF^6c[Q59^NF8N3JVOAP1eab+?9a+aB^bH.
DLUGP9d7a))7INBEg<,RZ(eb@EZfXJ\XdKZ#.Yd_UKAadZVH2CW;Sb#e&\L&.N9R
IX[f[)CMFR8SUKFFL35WS#Q9;Q04K.=dbSccMV+TB8S2,2eG.P,8gTTg\>gaQ(d6
#:UcIT^^7gKW>NMSQ8L&d+Q<IHc:W01>REO&GK20@<G@>/gE&_8dUT,8T+D&-L&T
960VJF9#C1b\gQ&PJ?I),__NS02V=VHZWQU<R:dSb)/:?4+T7P#8X&D..XBI1:\M
fb#V1#>W;O(HIaCAVG.AOO7VW1ec\7c;NH#HW8]B)(^M6Of78(^3CK8G)_I@aJ6a
SF]D3R4(\SNOC^b9fN9HQDA==,(14L+WEMaZ@^fQ;@Zc5f:]E#WIC-c(+PHQ0P[@
Y]_)[6+TKB>&HV#;H7-;Q)?YQd,.M>@Ae;S?ZB])OQ8,Q21^K:Y#PeR76:FW_GM1
O@:M.fXUV<W7S0)\K6-\Q2YQGD#T1LRWSQd1f+fEWMI^JE.=33N2#BE--X0W&R8Q
4RO<+39Q>W8c=XI>2[0JKK9](Md\C6cPQc:5RDa)(^NDVD5MHBMKY4\)OcHd>JDQ
Ud?(6LIHBRR@I85WO][M33FV6Cd>(6RdSMV_\YA+<0VCFY./2;C??DA>^:YZaQT^
@E5G7ZTJDHYba1E.386dFNE77/FU?UH[(>[IEHS[D?N7I]f2B+Jc&8YYI\JTK7+M
PC4(G6CgVbH?5Me842CcDd>1]2_SZ]H]>:.HN(GVZR&AZ<e^?=3<-9AA/@c]F?J<
ME-c4P37aD_Q^R:F>[@O(\WKN>d)C1F,],WFf6Y0(Z,dZGYJL<Fc1>?7X-OBc^AI
[Ed<\eZLJ\48G/-HNe=.(4],Z2/,XP1T1^3\O#7@C1);/-2@81(;;g884MAK@-#+
7/2fEHRG+<7]A>FSE)WZTKYZe_)?DDSI?:ZV,VQ#+P#[9GYGFYANZ\\VR[4Z2Z6=
a6XY\;J4-PfY8gJf_a\C;/+<4F#Z3&U24U>a+:7#SOKDN+Z3N[]4KMLM-dL8?g7/
WW\JV>V124?,C75dZ1PE@>MF]f)6U^4b@c40EW>9;1T\g80_Ue:7JO\b5.9/Dg1K
(D2aeBUfXa>\FMcd.ZKYa:Z3RQD<9B.-g;BgUCD>S+&+6=Mb#FZVE1&CERbRfcJR
:f_(4bH2Z0FcJb>2/T/Rb51<H3]/(=Lg_H:5XTfJ6_M@NQZ.H4#?dP7=J1)e/b4Y
cB4B6.^Q[VG3+-:,c965:AKIg+Q/;c6>0cd[&/RH]&Q]_dQP\BBV_6f\/fIK&[D[
STC:JH=MQ&16gc=,#2Ic]gVYBCX#g0c?[=_67\7gW)0W?=1KE]:<-SGd:QUBa;@H
g[;g:?/,G#+GW[b4B]ON@^_gO>WHCH5H@F1Ge_aR_3fLe;VQ2fNAMLW\NAEX@b3c
4b)7TKUbMgKL)c5KT>_41^5[T/]?;:H:VAC9+4_1]U_d^8\+6)0P7R#f5=c=WYE4
20fcUY#\M.K2KATX<@ND)+,/CbDR@2#/W9Q7TA\NR&5dB_(R(;:W)KFK@Q9?gE#I
gf9===@1,4ec00[59d[Fc)Y4BB11GMIcdaRS5C7c=V\TKFKDSGX]b:+,BD#FWaP-
)VY5F>J)F@<]MM^7GKEd;Tg)]2<31DT_7DZN>:LUKUTS]:H5f5:\L(0J>NeK1M(P
<&ZM6:)O-3#,1MA-#YA#&9I1;ee<dBK;,L[[AZaAH/.YS&0H>eURYbEdL1UMZIDM
P-7,\9Y@6>cQ4-J]+N5[0M:J<)T7MWN(6eD<Q,=X=0?)L5A+/ERIFb<14a>_)WL&
M)H/R?;e=e/Ue6+]Q=9_/TW@==fD/JO??0QCAd\_N?,KI-)9>>Z<R(C3_+=a\Sf)
e+UWJd5(RI(eI<@)V<T[Y1-65@:BCUJUHb/);dHI9L;>:gA1LEZ,3)X,W0WZ[<.?
L_-&0-IW+14GL8V4(?/,g7UQF(e85MJ]?bA_)_4PbCcYHbWUNb_H8YQK80XaHR7N
M,)Pg10@CK:K_RK?eEb;R6Re1:dgd:AGFO_7N84<e4ZAWIgS+6A&KE/0bGAF>?/<
S&BE>Xg37F#A?+4#6Lg,2)5ZU3YAAa8A),A_XF;,:?9V-YQAY5ET4(5Q4.7V3/B&
)\WgG(Va6X7E#T.\6@LWSTGQW9:T4HAW7>a:K::@VBIaZ=Sa\\TC0=3VE,(=/:YP
gfX]BX8WRG/Scc@-<-f93KK^<9NLD&a35>Q_+>^eFJdON.BA5]-Aa\U1VPTHKf3e
,Y)g6Pc63A=PL+IBEb>#VDF2df41aK,Oc0(J@c8^3=b2U.Qd<@fSfa0OAR94B;I+
@77J-R;7#_NV_7/59O)gF.<R6Q):e&QJ/G]+BA<A@8:JSb2Z1T(/1XUK.c,JZ8@?
)P<EdI[\=;+N6>?LV,][:H?9WdYOR:7C-IdSI@2+#_fFF2G-OT@3>XTTO0&5cVUH
B[1a5HPaN#1fV/0^V4GWD+>\6?OK5D1;]J=2A))9D3ObLLK_TKQGE9GVf<:]_3Ra
+9(E&Y#KAU1H15gQ&CI7gdW6_S?=-24QA.1#V&1PBS7(@-fTOX.JUSP^T\_C(&/O
L(B;_80+MPIV8:eFBL?GeaH_3+IMZ:QBP7]3TEGYaDM7@Y8S7AAbKV-SVe)WE4Ge
gZ,1bd4JKLYCd?/\S4TI#AU;;gQ6&.->c\e:\^b1,CT>G4TO=\DY<a[@82VaHV01
<V6ZKVCbDM2P3/_]]6,\[Tb(J7N8R6QNOKHX3COQQRZN3WQQg<D]LdTc^/8U@SYK
3AU50;(R+9V.B8NCS^^RP0X1CM#WC9BJc=Zc/C]Fd2gFAPC+U;68Q/2c>PI&a0XN
S@+1/GPPc,E@ZA>Z-/)a_74LK9a:#c3Ja^9<3R\.CFa3D&gHeWT7;^#CbZbc#@3<
#(X?YI/deAXB0VDCd+@5K5N_J=>bZ<NZEX.0NS-H_D)b_:?6TP_EbPbK\0,7a#WF
#Sa1f,>:a-YbS&0H#.G[3H7E8MS.Sc2#]48C=,X?db3?Nf9S^^NJ73FEgK]@W]H-
4\D1g([8.=\K,f&IBN_5+6.71Jac^0^8c1LLJZ#K&=T.Y1TfD)11f0#VRY4FFCH9
;?K;;QAQfAY.A]]HWNKe/2?-M[HdC,4e?@JM/]K5]-T6.9U)FdU@W4Y/Y#[:[P8W
\:+f\)^[<]aV87J6N)FQ6G;#0DGZc8>-Z3fIAJ)4_WP9f+W8eB<J+Q8#0([S&GbU
,1A^+H^Xf8_:fAW(7[]be->;4065#=<8Rd/\d<dCX/2BX2#MH2N2>SXF\aE2f.:8
?/FeE4731X)Pe0_0M=Ze\EH&7#RHY_C:0QIO&32f&4@H)B(3:d+-_A@:<TL0YZP:
5-VX.@MUU?QH_=f.B1O_gYa960SH&@-M#-0IPQdS9G/#:b+NaK^##A(0AeP+95Cc
88..,1B8cS?W<>-6e=Ob6(3_21<cbW=5U]]N;e1)/>.-gcFGbe=8b,7N3:;KLZX9
b@:\-HC#Nfg@[dbU@+_,?_GWDLM];^#NCYGJ/4&d/LL5^=f==38Y:RcGa3X&DCH3
B#:R+;2[#YL7:N-K1.75>4<@aY8/.GFY<H)DQ=H_BFQ3a\ZZGYT+A7,/^8,[TG_M
Fb-A&2XF<QC]=gX.)S\I.e=?&(,M>U9^b3;]<CN>];G:I_/e]R>XT,0^IN^B5VWT
7?0C;+8DFL:PGO]AAcI5BBE@=RZ@KfDWA?COK0D)6XH/)TIS(F9_HY3G0[L23Q]K
8+C:?_^Z,7PU0<9X\UY0CT&92D//Ta]A)\ZA:&H)(TecbM?01ILJSSd1IbbZ?#Eb
WQ7\ZBTXdG47_T?()V)&XK-GCG/5/7VYbYM6-+f3E&9C7MM?1-c9A3=TN6QcI(cT
4;>&_KI-dBfdRQM>UgAFB#FPdZ8M2eRK3L>U>TMGf<I=O?>:aNdE@@]B^M8DR8^]
NIK8U7LY+(Fg3#)2C4eQdMPX-&EGW],>JM&.5ef+@O\IdS),V^MX4EaYU#QPf;<#
_#RH/=<.=d:aI?5H=/?G-a[KFQb4=9Ja4]?<E^C&&X/d1\V7K16c?<M@WXJ)g2;M
@LD9Z_A2M]c&N_;N);((c[/Ce.O;4.@,[\PJegE3[>NDPCODPTdg:fAJ(VM;bA^8
ZXEb1O4LO;-CZEL#G8>T?^G2\+\3/)PSe^01B)91fE8gBQ_fRFL9(G]<?,ETHT)K
KOL^a[Q?gZTSA^VOUGH7P9,cC^BB:eeJVH8]&OgL1_S2V,3U7Y;fE9?H/(5<]A;S
FM65=B(>g/XMAOfWN[dFTCeNV)F#JM1E;.ff#K>Ad0g1X+<Od4^?7#Hd-5,#\#EG
_J>]Q]I-bY6QSS<HbeA7K3ZFb4G2L^(GV8Je&IfH0G[?<6QTED(914Y,]/fgN#2@
X(IGCP;<[Y=L4\c#>?W7c4)HL-?0_W6^0[eCeG]X;F(;H[Fd-&7DA+8:1XH&IZ01
)[5/9I;beZY\baON[BK[&D1^3eKAbAYV?5X:K&):5c6+KG9OQ<0EB1R2KN83/02d
4).@6@FQUf>-]:ba,eKA4@gLFP?].]^[+eZfG/0M)3C&(SNB@6K)5#2]@:^+bC@E
<WS)?/Rf_HS_:7VXfRBHK9DdNB1e)F6;-RGQC<=[F0&&5@f0U&c0]=2SPBG-ZPUG
D8X?<&Eg7N?PK02D_-9fMQVDOfTJ:@5:b_BUS^W1J.,]11M-0&N:R/,2:6;:VO9X
CYX/eP[b1-YS.E<YU\4#O<c-T8g-g5&/9?-0QNM(B(5P5CQ;_A3QX&fa1<(F_J#0
64-AX);TZAMgA2R&0RKgRM+Z.CcP,ZHg(I^UV;B8RS6R?Q]_<9c1&PJ(O1MZ@RMI
0I]F9X@c#[_6;[:2+1X7)DA^N51a]IQ?OEK(/)8Ee8(d89[((eI8LaC]3+S-S^gJ
/&(G9G)?fDFJ+.Xb&2,R5b6[,8gSHSg-UgDb,.<TI8MH,U2a_TXBL&1S@&fA7WbV
fH@0Aaf3^dNSfQV@fOF<g]B&^[FBS([cgQ>M[82)SMV5Z4aUS[/;4TW]&DHG:;-S
(bMIEL?\cWZVLGMMHLUQ\V<-EN7S;fNH+8(+fJ>L(5V#;_?W(_7(Hf&e0I&&0RU7
UZS5C7O)D]R1(8BdZ0eTfRU?YZ&+>VXIg)gTTUSK&GDN&<3b^/eG.CW1)[F,E],O
L_.Q)Qd7PKPTdIND9#0JGSDXbFM1e)::_?FKd+QM4OT]Y+-BC/YDCRI2P;.1KF#P
KfHQR@+e[_9;(C?J(HbSSLc6W=Iea9e17c+XG_LI>2K<3>D-O0gODa?:7IHM..R6
e-:gZ@a+0BfPK,]cKQZII)8M&0O20g#De>:ZMH8f(FZAB9/P@5Z0<S-QZ0C.<>&8
7@^WJ3c.SG^R^H)&[f1?P@HJB-59WR8#4RM;3f3]VI:T.R0E34V\VWc=eK>CTa?#
_>?LTc<QBRHG#Z<A/?U]EOXXJ:](>B6GV\6?\9]d5>5D)F@JgM4Y6fJ(aK.g@KTe
Q2E</[FD5CYF>8^2JT+(X5G<RA.Ya8/7H0,VPB5W\g#Rf?6T)OcFC/K+?+)?,(a=
U#7)Y=\0-\fKG[<PH_L\5f.J)+D(MO8Nfg9RZF:MXFN-(M4d?\NY>2ZOTS?#N:S/
8EaNZG,FLdQ.&D-L_/+G6d(8<dC7FFZTHgAU4W;8Z/,9e<PVVZa7,>gD2gOJ1YNf
F2=BH,WBB9U63fa#_5V,Pf^ca>Z;0I3,&,C?8)_SZS4gH4A>7@/XY=5_LCAdGO41
Y,M_8976eDe8+I(e?JGAg[G)T-HH^G0G.G1IH@S[1cDa\3HL<W.Pf:48JfTbcXaW
^IaH<O95<S<1IQ0\S[9X)YTcJL&1G&;f=.8#]:4X+XKGfd7/IFW8>F/g-]8QA6(<
ONUfR<dI8583071,fZ5K+\K8I;V.1F_-NYOQa1e8N5X_,<+Fa(UeQ:#&R=WNK+SV
#R.:[QXaa[Qg8YE\bf+-W.Q1g]-B(7WB\M_B>.WR&fI.R.UEBN3YYI\HBD;=@gQ3
9)d@C6._;35#DP=8E:A[gHN60B+ad8/V#VeJV;IX>,&&d1,U;CP]-CZ[NUM807,P
:@&#KCD]6^eZGaT?;LE1eZ^P#\Ff,^[Q6Ec/;PO:Z>:NN56,(N\:4,G45Y?5c;Q,
6]CbXB)B>_K]=UU<@?-DC>)_\B_-R4X<Gd//68V?e4LY2KVOV]I-_@J.QZ/f[gGL
N)bM=@]?;@?cL(F#FEU++=.eK(8KCKJKWX)GL0P33CNI1=B/4:ZZ1UQ42_cOBMIg
Ca/Rgb=&31.0ffKPbS/ANP)K(E5.2a\=5QaP?^cZeVb+X_dH+2S6>MX,.Q3>4(0Z
[.S,J<1L\b:RL^MUFB_g=aKg<VAXcS>S4A;P\.CQ#UL62<W>39IWS0eNB:PMd>AR
DFCcbP5(2-dbMPTTGWFcY#</?U2B^KZFa_f+d5/8FN2[L(FKP-IK9\(+J7e)9A0C
f]J=@S=21P?<&Q/b_.\[;1W&b)[CZf-GU7UXNXHP:Z9WP1d/ZdBc]3:OPY7L2Jg;
YLY/bLG59XD08FSC2e.ILC^0c]&AFL5b5X\gT]^))&fUBN)NMNUFON=2()[9K:7A
]SeXFD.D,YQcNT9D#L#O[>+)\Zc3)JY#.NJ^WVQW:O0=\b12-.[:C5gVCA:SS=OJ
\D6D:0TA;=64MJ3,LZ0?^E)A]=/+MF[\RC^DR2_Z-XG23M.DEE#?VL+af=1bfXaW
UGEc.UB=&&4g:(8gfKbXedJXRIJ0c:e:e@gU4,XHPOaUgDB]R[(<67b?H5U,ZJf=
G85_6SceaL/7bcKCg>(O<5P7ZW=Y-gLN#F#3^8UAV5JAL4LBO_g)e/6(7F2dLUAF
1Y^.Mg?e\4?f33M]Qa2?AMD)@=S#-Ed,b#&EY@Y.,5GB)Z9-IDJ(KcJUH@7NV,f@
^dH/#dN9B+Bc-MBMTL+CL?X1+SY,2#+-KH_2@=)[@2&UN4->.HIOE2Y?;O<0^1(6
\-4@7]Hc>.6T4+^:&2MK0[baAf<Cf0_IIceS:^(ce>ec@4;WW241b,5[,<X],:gb
c^eELY/L?Gg[a8FIERAd+)Da[Y]O.]_-\QN^^&(7JIZ-;L:4bd#^bTZGG,GM1D=-
(ODK@-C;F(R4M0_.7HG.+,CQ2;,ALOFQG9A5UP<[f7VUb]K4S>WSVG0U=87XR@8;
aE-LQcbR(f,FS?^E1;\]RT5<[A?QJ@W;c.-LID@PeeWTA8fQBP?YPEDTZ(:KRLNG
Raeed-+?BNRZ=61.3&/TB75=:BSPH6?K&Dd37LP>)31BG/T.OUf@>aL)_9Z2-&4A
D2(L=LQ&BMfJZd39G5\[Q7^8BB]1-G361a>-7CP]H;.Td)VEU+1O3Dc0DJ;0OAb>
GZ+K2)#aLGE1_/F^&8MR[P2#b3,)3K4Ld8(T066bKJ]fB)F#A][]a<J5/_/V)2-R
@9/^fVb6V+Qc?W@1ASZ0OED=gR.6<3:&712=S.bWGa\,[==1?=#bL7eI>ec);9[c
6Bb1B\]d4>5_D9IW_R<9A-LFa+f3EN>fX)DO,<6HKC2,.S0<a4W&WX><.,BN&;W7
.:@EgPcE&PQa:0<1G4+[[]U+R@:MWC=[d5)DCJP(4DG/@BI0/FIHSR@g6/f-MZ,.
GP]N=F,&AY5<DS^27^U2Z[bDL?Q)@6-7V@fcgT5ObM>-(;?6)S]G-Q#(,(XW[9e>
__ce?(W^4Kc#?ZEM9;MODH]MfcR[Ld\+=+]U&?A#1RY8M1/@Z15g?X5_c<J>4e:=
RLLG5\43GU<7@PTc8PG;956QH+[T.B[F1C](#EZ:ID6,T/>TM@,c0VG5B]g782E;
\M;b[=d6d4#2JO[9b72,AT0O:2cA&&aQFD(_I8e4A.Ub_K+1L)F7K5V84Rf-<.X+
PA&d<f]&eN02V9HU2LU=#61@9]=ZNg#CK\MJQ7ZSQ[IRP7JAe&N(5fTJ0bU^YO[F
\R9UU24>,O0;5RI3(JXENU]5H[Ff;/QKIf;/<g&Z^JgRX,INfZ?TJU.X;)),QVDN
TRIW]cMg5a\bbTFZ>24c:7?73;I&4Tg0K9@FU67Z>V]Hf/16&@[U+CdVgDG/3[A[
<-+>K-@,[D[=e)F72U:+4e\,5H@AaD=V)g,]9YMd1E,5=IGLe_.II9KW8>VD0>H;
,PSLS:?]L+P?(2>EK)(Da8S2Z<,@_d\1PI50g]C&6fLLIAf]3]WLc<4)J#U0]Ac>
WE7/N=23Sd&NEZCF^Cf[)Y60KOf+F4:@aDFM-[^HD^]K,ZFLF-6NOA/^?^PAHfb(
-@(,<@e:,W/aDYC\]JB\;8[1LW1H]=KA\d\ZXR\YYS<D^BBcD4#<SB/B#X\-e-K?
;I)1S96INJGG-_D)1N=RJV^/,5=F=U[_9699bU/T#&W6/A#+^>T/YeD8R\>IKB6S
O+CH@9f1?Kce=Kg\X=BPL81ADU4&R##\:>++:N,:GXcfMP[A4N>Xg4=-K29:89\B
FAX[LY0L&QQFWQ?PFb#OWEEV.NM]R.:Q9;JBB8EX+1/TSgJ2,.3N7EUg<ZcS?3(]
TZIAcIA9986c.0H_8BT>,8Dc098)aP_7)O?(K<,O&6U?7Gd6U5UD&M7AZ56.0-2&
b?&V9\RU;(A1W\+-F@bZU+5IRQJ&.I5UF+a^RC(bM.ED#]AdL3dVMQ?#P/]H3.D9
@Z191,)G]dT(.=S,,RUgdY3T3Hg5EQ7b[YXb9dRf@)T;Y,N6:/S:/#^L^6<Bg=eC
U:\(-/-F4?9MK-H3Z<fLg#/V;-JVLcM3KC.OJA?RcPMe,TbfW7Ka?CdKL[T3ER;[
4#DaH)^OBLYGdFD-:9?B[,G.W>63[b[WORH2D28)4W\@I<Pe3eQ+)B7_Sb6<HTI&
,fU&-/-OSd#<U3aC8_a6Ge++(PQ/EC1&37a^d\eL1HH/[_YXE65R?0[SF7g/W]I3
=,fHAe[XI0LF=IX(RZN]#e+,eI4_WY&&EX_LTRC0[>0HJLJb15/b1+=V\BXaT.Z6
AIRI(fS+->(/>52?]&3Z[B)&ce[,b.4)4Y,9gJJ+?9H?T@NY\)gD^=,a?aOb&ScG
/c+VGaaNB#7ZJND[;7V/aE#^C+58QcON,V-SH4F.Sa^b\9,RU&I1P5&0B/c2^_(4
H)gSSV811_CfQ>#(IeYB+-fY_OLB.\X;EcF.T<F17B@cCN;9116bb#c,YNdYUXAU
X]]G9^5cVLU@4\W=:[C2TJAOI;?SP3/GCGQ;Gdae:=LW0D#9)1?7>EU_L04Z9RaV
2bPXLWcO3a.J3Mg0.@e07WIaRP\d\:A<3IUKd<?aX>]e?N,5MG7<,4&e[bbV(<M>
C-;LM)fZ0d@CCN&02bSB<9Y:8&AGA0_INNR<(/3&Sa2g&/(^543_;(H_1[@:MLP5
\KITgO<P(RTIcE,9L@R40Z.>U.B[Fa1)Ce@a]6Y4T;IG7;;Y9SJ:9C3f6=4L2RF_
2L-C4.;9fJ/DeaF4R>CT9F^7L=I>#B;&J2.Ze,7MZ4QG-c3Z@QTOKVYM,?GJ?)S^
P:cFMTG.fg/^Xg;:5AMQJZ1&aFCN#8eTIeRV)AQ>IGeA&OQW(Q/]+dKUU:?:O2B1
#\e=.ZIX<(F<FG>6;F8fBO5/OHcZ3U>5d,^_WWb+McY#KVS_,VIL?[GVFgVZ6=DU
57SG).MFbcWZGT?@aYY8JMZ;+C)DF42GPE4V]VRa:=Xag23\R@&HGdB_AZJ&fUS?
eT4f]daA4ONK,HM2gP^&,\Qf<2-Z^O:abUMI1eW1;Q5=_3AcE2UHE4>;U5DFd1_)
-]-I1M)3.#Z7I13@3LZ^QW5479Z8A0,eVg0(\()#)O01U)8PNQL;b]_>\\A)&]7<
.Y7HV]BD+.\bOgU#7-^MN8(4.b&J5322WI<=U=D^>a[8NZ#N.a0-:^_=OS.37Deb
I^-ZGVgRS9_+18+PV76):a>DFOYdWa:459d3.QU4FAE80+#Q1T646)g/9IT>YWV2
&7Xf8))1C8UHX.@NMe.LbZ.eI7-EPD+5Y&f&EZJ2J2(BAUP_@0U83RS.3_4[51AK
^8OG\Ge]+VUD]:;VI:+=]P_QPX1^d]/5ST5IJ(]QXCYOD@^KcGL.44HR,54-cLY[
dQ&8J\?GR-aYL](MgFYV&e6/@E:-+gN2D^HJ-BcZA#?J+PJ11[\-g,T7G8D,d5MM
98(_bcC18S.P]Ha&FOa0>(LBV]&<@,2G8&JAP2NY?SLO[G@.f?,@1VJDTWP0Z-PD
.TcG+e\TTTFFZQ1D32V+<+4dZMM<ZYXL>EUFC_Wd:@bJ2A1K(7?__XK1a-da,HBg
0KS5@acDHePNZX>Qf.EHR1IaL[F3O19B?eHB:0aM]8RM4>#VD<Z6J/R?Uf,O>V=)
@Q5f&(d<_FLP[F83V>=F0g5Q^7:P0IO1EDCa/=0_H87Q+)Bf65CQW85RB\)UaTQ.
)]=PT;:FT,=7>B0b/_&U?A_1JS;+]6SJ581VHDd\=cNK;Z[[,3D=0b,QNQgE<I&4
SE3f.AD:M;V9)/^77c/S@[Ee@PG)f;Ea6RS4aZ=EQgAQP21&BGW\>_9534<f>>_9
G;_SbHHK78Le]J:0gKB\_T76#H-GQ..eY_CZ.c]SVY8\2=JL#081eAVVf[?:XY6_
QO49aVHKV^K<461?WK.CFTG5SZEg=:UZ[8e7O@6TG;Y9Z7]A-MC>(]AJ2B41Kg(X
JegVX?bbFeI9Q(PLcBWRVf;QZMN>MIJ8)<EJP4O.@1^J39Cgd#L4LEB_X,_6NMW+
aB[535cNF_Z5UAdO,/0QU&H8X_E-AcRRSeU[\EB[^0JKM6I6M6SQGGH69W/YCbZ0
#P+HAYQH9H1\=J7<,X@FXa/L8Y6:DgQBY[RB@[&L6@5PUG3UYKYI.?>LTZK?=I\/
P(JZd75]5OJI-2AE:FdV&F<LLJ<P/&QLU\:7MLNV2P0T/&#+>((D7Ng;d_4[7??9
f;IC]]\J(QZYMQOfHgN.?HN3SA<<O,R8;NcBS[?\O/<f:)9J.E=,cF<0[.,YCH-/
X:dI@ZJ,8bSNS^)59OX6N8/=Fd<_EKT5->7?9QI;0;V6[ee884I1N)RcE973(A;R
EAe5K0+5\#M,7?_[)MF&UJ@/fGZ43?Y[_)NF&(:3(=SI<Z60-5Y7YYZ<(5e(@=fI
MC-/9NOa@:8J?#Q@]gC>LCXEV6-a3O<R9EHW7^20X\=d2YRfW1IU7,DU(Ye8R03[
(2GZ;)+DZM):9ZHV5GH-6KI7AH(:2+c[X5beC6FD(7:VXEIR^\[]6MZJgS8GATG]
\^SWbLR(-XE\L<Z<(4a#da))KF@RC6IJ66HL=ZbF),H5,SR3/PbM+@_Y8#<Na3_L
)\1)Z;PCDc0Dc\eAI@d?3_MUC;.;9/(W<dW+G<AM-&/X/VYL1\\AR38dA1X\2RL@
/gH_\QSScVS)S>=(T7J,JTdaDVK.44JD45(@,\BQZ/8MdLO;Y@0?6&^?[E/gQP&F
_D1K;@F[@3<d+47=SUBQD;8AMO-P,/ZPBB:WW6D5>G:;UB@)8-4ab?_(.PD83P^Y
=LDD8;K;=RY9fSAQ,QBP9#-/:^N8b+C;-)1XQOH)R-<C71W_3@SA01-7O,.)P,bd
8.NYYa\T<JRf.XSM[C]d:eZ<+9Igc8c)e&5>X5bfCN2bY.Zf)^=<CS-81e@;0#Q8
E^4C=VO)Y0(<_^JcUMGe5e95P9,b:ZefcHe;aQ4]UW_Y^JF>;aeTeYb#6042<8_Y
GPd<-UTIfa8B6FB;9#LDOHcR)OdgcW8VNW_dOMAJ7BeKEf&6\;23X7^H_B,>EH4@
(4BaO651BT)4DVGB9E>;Q0.@:&/XKF28ELIJ):f3XII=UBDD7A(E(T-2(+><Ad@]
+H.R(fO/)LR8YHU902YPbfd:X45\:cVKFd:NBMK/=&X??+.:UHYe\+A4^^S/76fT
BJ;;#]&-H1Vd>-5N(KSJYKZ<^KT^bTZO.gW+>egdX7:,^DKTYCb^K3HZ+9M[dReD
G,R.M,,N(B1eY[(gP#/M.KC^?Z(YPD#3+,,:N_V8)M,<eR;E>23S76]7UeB9P,NW
M5;:+##0D;7WQCb@6^?#U@);<W;:@<A_3JA#RIRJXCeE>)0VVKYCVVTS:d@@<NId
)&gNA8.a8_A81>^2HOY)<2gH]:N?gRg>#GSLIeIA^X5feILB75-5Y/cf?CKAWAdN
=L1<@5Y\HFAJ8RA>UWDQQ3WB&+<dY\2W&S;@e>3-.D8-7g@F(a./FYM3X^:HABIB
+.Pb@ROFGQN&,ebE8=[K[/;66GeSVb6=3M[U3PZ47#.V9VZ6YCS0^0B,OOR93)E7
-A>/21;V-7#5.MCKY@G_MK,:GQX:fB_NK7&<.R052Z[/A&>G(.0U^C<SX47?N8)0
<UU3Ld654b-IX:/?4-DR_?11-+F>/M?g(/K\?.dK[+R<,.]10C2^</^#3#<A)RdF
FE77NR^+HY5&3QJTW6]MeD^Q/F8-XJMO5&,8HJ[0b0L07H(+g<#63aM-=[;U5d:e
W)U5SZ/7<+E3XLRd-O=^fEBAE>^1#E3XO.5Y48INW>\9Ra7XM98\;3U0a0^M+X4-
K6-@U]_1^.^Yed>^aFLc\2G17,=80\f4P4[<=_U8KgOQ,S#CLa)_E@+QW3MW-QER
S55LPX4[Z;aZ)eN1>^d<@+7(8SffT+\A;<TKMb+24OLbR<&P_=P@Q+NA1c<(H=[b
U,&?Sd)88TE^B0P@S>1.-Q?Y<\3H&].SG@_8K(dVKBgTa7+@R#:0JZ,5P)\c_0/a
X.4[+<4.[b;-X05a,VRcJ?<5=]Pf8B3R(J)C0=PEPVCARcH@+AQN>&9M@&-SCX7B
d:NFN;Q20b.gHZ_g4_FBf6b<H::Z)2+CU5_XTJbCNe78P?+:._6Kf2JB&.e6NK=5
#fVYN1L=7MTX(UZSS96;TA2C(J98@Ub9P5a9<NCGA[c-b;g#VFP&Q7?Q7c<JL=ae
Ga[Z7M.(BM&Jf>1W5cID/BEA5THQ]I0ASgSS,YbV9;WMN3+4/(1:.2L.<S&M7MG@
N8IY+(dg3CZ@W&UY.QSFQdM\FKfA0/IR^a9H#\E.HY0;^&;Y//U;3_&9^Y5^4^]K
]cCD-;P..;T4]X^fZS\e=/<9G0T9[1F^bMH7-a^,M(IB2:+&HBUgP@<&X8@VY:R=
c2>3](Y?@cE_Bb^1\0?<3P(FMK?SOJCe&)=KN-U9Q;[23J(RbQG+ET6]R-V@3c#T
J<B-0PMQ<5U=<UJ2</e2dG=O[U_81GbE=1e>&/,RLEG]D920dg_4L+ZZ[432,A:D
Ca81g+D<8H\3N\38)E[:61AR]:8:L7MJd@0f<N25)AA\7^WVN/b5,4dNO:3cWFG=
Qb]J[^A>EM2e7Q3O2\Se4&Q\=J\C@#HS>,X@&.8ffO/60HR(UKDCUX^&DQ#&R+X7
[>7_eV.BBf(G2)Z[>.7QB/)S.\fL]Kf,XMFgdg;6I75.^B[;dJ?+^(A^XaD@4I-/
7fD&Qd7[L\:LZ;?M,dH&-T[HDE+G]O]U)H+f((#BY6C4IMM^_8[?6I:WPKYQ3Yce
fcM=3L>\[3XLURK?_62>JR[TA)^7dO2PU-+G@I53H818:TDPX@D#46La6NCZSC)@
Q#V9BIPb<+4,-;ESE[=JRED#gdSG.DdD:\5_0Y=AR..N\#aI[</N<AcTW.,cIJ:6
fGXZB02Yd6+PU7+7EgKV7W^\U/e51XU+g22/9H.R#)),>M3g<+#Xg(NeL+g-+W\G
GVS)&,LSOA04AGN)546++Q_bb/I/c.0X_Dc:^X;/R]eY#^Og&K4Z<?W=80KS/GQ.
b2N,6YR6Hgg<CRc4Dc46-bJ/(AON:^F,Q#/T[FU_VM<FRab86MUPdXJYfGG@1-K#
,SAW];fTEASF\J=MTa2f_H7&Ra>;A5\WLE[6GbR<GU?MQ&;0>4f09a4,5QB9#7J^
)90/L/7+PQb#.[]b+?R5QR)-ZR@5G6XC[4=a-1-e=;\L=AAf&+J;TBQOaJZ:CSdC
(gUB=@:AZ0-?=3^&a@VA[GTO@/#;7]b/RQ+)Fb>W9J9F4AEMH6b7K3PVG=7P1U#M
_Y]ZI)OE[YZ2&c>dG?:STJ&,ZL2VS;f2P0fcS;\7ELg)O[8NdaLFa\\HX9B5YcD7
O/BJEPg_?#cNM&ca-cd.LJ@DRSe9g>[KQe@?2Y\NO@@-,>D1AQ1/g.H/.g:^POAP
-7+G208bC=A[dNW&Hc^\gH9OdC[?-O8f?KPS=?JHa4U49&=/X7ZIf9/-V3,7d49)
g@-\?g+.A\4#Ub.REK_[.2G0_?Jd5Y)\C^1a3=;PUMRI;IfDT=I:4b-)K)#FfX,5
F07>)d[[-A,S<F-7.F8.1<C0LGHB>e(BITbf[51FM&<QEN,c;1WRTX/P.U:7d3b?
fRZ4OCaA2V8W8Ue69],E&0>74JCY:IQ(LF>e>4SVSS9>&g?(0R9<8LQJB/+b=c-I
]_D(4,3ZI;]JP-->80SKa<N7Sc&cb=/?Jd>7a3T#KGD@99SWL(Te]aXfgfYf:QWD
J;[0.L2E#UAJfLZMNRR-e5.f=45e<C\RUFXBR^UC.WV79;:UGS_/LJ0-(U3fd^65
2NUW0b.JM2bO?0XPd_DQCW3T=94@#E00QW^fO1d5(]#GW5BP877=)]8W21.7RX_K
_\V2AAP^aL9:f3AC7.?&O^LA;:/ES]]L0<WN=D9\V?b62DVG0@88:;_^?D8Y]PI&
2=Z7gdc:/^7^KBd,QAQ3?=6\G\3eUH&=Y_/Yg)eFWZUQIU-R2W<QVTDG]IA?XXF1
F74:CBRY^]AP\3R:0#LV;S2P6^)+U(?PfTBc@1F,\W1)&IV9Q[6#AAFgg:^ed7Yf
Q),A/9cJbLX->@Tf_\+J=DMU?g8Z8-_)Yb8aY/Mf(3P<,Ugg9.>QO/JM,=E[4EO1
d1\;BMWF-+BZZ6D@A70TF9Q?>g(AE,gPM2\ceeb3eOeIN<N6PH5_.OWVC0CNeeVg
AM151RAg,#B_T(/VWOZ0EUA8Z(NW]EHKaXV_<KN20.B-J[f:/EVW&D\Z?X[[E805
NQ-G8);K8TgP]X8&[JD0cGX32Y_E&R\I&9)4fV]COIL17KBWK]&Cb+[;-N/I=DAW
U_I8\5N5(/W)d#UD<FGW^@073_&N5N]WAAJgW=G1C4N73b@GK2Y@RJ+5dd(G)1IS
O)+Q4GcJOR@L<b#e:0OS8FZ7S</C=CPPZ[NH=L>Z9WYZ\#2\E=/6/P;e@9Fg(E-4
_bKRfg6E0Q(#3)5;@2aXL8\Y=(T./WJDR;=a&.Z^fE==@I?([2Ng7Y.fI^#==1NG
V-F7M(HV-/#8J]5:S&0>QaaE(->N.<FDA8?.8?bMef.,&U,Q40W##F.?M)>9\)K+
?@,AWI6d&TY6;1A3R)705_MLdXT@C#OdIMNB9Ea[SRG<6]2c=&NCXRUO8^)):^&S
\CYOUDSFfT].HaegO@eW/)TCJ&;B-Va_BJ&[/-1C.VaXgHb,^gc:;Qb8d9KCDSd8
S+:].=bP.<@&HbCF]g9A?RFM@4/:#@=G.M+O];GD5C?<:bV)HGc9?WVZEaea9d(O
0a,7&@@E9V91S75\+@)\ZBB<f\2AeeZc2L8^WgXD0GX02FQX_:=5M.?1Y&)=PF:B
ID6(OaG23N2FL:MW08OBCecF96Wd=-_W(;.;CUXe)4MKVLS4P439(>PGJM+YD-TL
JdZKdL4G8<)[XANN^>9fWA5;Tb#)]C(:FSV[IgDYS:HPZOOPSd4O4>)Q6)>A[R74
BO>ePN?EUN>.?c^(K)R-&^VWZYN6c?[><1J:gJ&;bVJ;;f.3\S&A08g#EMR7IJ81
RPB-e5V:FER1)#3.M3]R1G\D?6Z&+^+aNKZH^J#X<JUMWE[W,\?AL;Of>J_;O;#V
MYFY:dE/U3PKf\O9PPQ6aDUeSTb1T<YHC^FTYZa-I,)Qc9d?PbPZH65gQ9:bN855
gV=,QG\=M_=C#1BA#SK8RS_gGG4B=f_PD)<):5]XHb=/J@McF:PT?+Mfb0E-/GBJ
T;\),U]d2XUX?B3A:X?eE^g.WEL^U4VL+@R&PDf/3VVS^R:K)>TS\7aZdd>?FRND
7[PN,H]1E7+JV/U#>@N@<g-9X4f1fT)R)W+NAUPcQ)6)G7NHTe:AFfYf(/SRZMDA
I36Ve.9:MM]O0NYB(]S4D&fZf2MM\&>HE9_S/;K)dZ0YHY-^eU:AELBd8A<Cd<^M
_UB^EIL/>N\5D/d-0_3\3M_2ecMY-NN@_aEdTARMGU8&W&1^WK8&#K1;a3-:>MXI
;X9_YO4&J?[TH5]GPQF/:&FG3[T[ZE=K]8+)9WeU@I<2a43<)8I#-MS-AQ8>K:[/
7,c9D:_V7PUF;]TP^Ea6LN9DMGcMa^6KUa?-[PF:_7R^BA?H^M1==9NRMD52QMQN
d;DNJ_OD;O^WfVYY+3].bTWHR.<UOdfASD05O#gbUA#2LPXBPZ_+Lb+5JGY9&7I?
cg5W</.S1DE8_T#gS&DTA<eO_T\ae45F)RT,B\3.b2<Vb,NO>NM.,>=NE9_DBE65
FJKbf:KZMG+d0VMdggJ?6A>&E;5?/GN1QFKcV8dN]-d&D>:,9YAb0]-T0G3YE>^0
D)gLaY),8aG;@>[&):aYgc/]5&(/Za9>a;42=E:OR>eQc2^DLVWGM-+^JC3.E4WV
H6Z09F+?<O)]H29BI8]TeS;B[V1MC1E@@]21MeCU]f^RF<Y[:.OM]?5(ESZ6SNL?
S.5LN]+5@RA=fBN(/6_UFVT,2O3J&?I-&]L1;O2gdXaVR)X4S@>W=J=WJJb4Q5S,
5Z@F[WB(1+O:KP,U<V[Y.PSOf4F_B1JdfX/NT<0OEd)S.2SGd7]8?(WF2VC1&ZP[
D?0=(-::(cZAQ&,NddXKY:V7Q_]T\HW5dM4O[&bU6:8f85G(D:+NY#)C#()f/#W&
2).LX3IRaIY[2FHFUbT4T_3gDP0I#FGGO,>>T@:g[<FHZOWE9IPe8@J:M:GNAbDa
[6CRLR\7F=_0;<bM2;2#3)^=Qe=(Y7KL)&L;P8YJ2A+a[,2=CaPAC\QGfO2.=<+T
UZQ:?/,70:gC)Tb&YaH__>>G<;b[gFfSS2c5cQ?T&#EQdMD;6+1P\)S;XZGMcE&G
8Y+S7gL.L,-P2>PGESeATM=0^U.(BT0eIXNMW2?:?Fa>K(B==da3aUB.D;,OdZ(S
KcLf-2HA6(aaC?6I:3T-(49dJL)<QEd)S@d26_f-_eZXHV,4.+NOf;:6U[R?:_=A
&Z\)6/42,[BGDb:fa;Ze7@;K<U&=_f@19O5VBeFHZAVaH;HE-+[16]+5&=a(bX+K
e@SeK^(CQGTRR]/7^+Q(=9.=Oa=PX8VW7XT/UB@1CLD\R=^=]2?#UF6>6FZffZH:
:5#X+=+=O[g3_:A/)g2.aTYB9If7S-0(c_KN3_<QgaGPZ[IX:J&E8ECNQ2_VFK;7
HY_e+M2KT8-gUH)_7dPL=LRS^:[TG+.&@]6M,TfG\/X#EMc1_+\;407d0SEa_54,
;=SC0A1c/8W(NY_ZX>MSXeZc-R5gP\J?&&AD(+OM02G1D@N;V[CDfbgWVIb32D]P
eYDa&b64V]GUEVE4,6OV<C;E3WgHXGSN4LgQM/[f0\ZZVf30GDCESZ,)PPIXfDW\
DJSOY^7G+C](7D>M&-.aa^[^eGd8=6;c]UR08NGOPK8WSHc1f6ET3]LPVKAWNbcY
8OGbQ_O[A2UOE4:Sa/e/V-b8gDF8OL\6X=3RaN.(2F/BZFV3gLZ@X)H2[N((/e-T
I+;/\R55#94.F3RY,4Z22>97(CF^]U7aeGBXAbZd8,_-C9=VD3RE=\=AD^2bI<^=
0>41O1T7?E>Zg;LcG(HAU(?DR+=?fQ[+,3#;^E.+eNR_;f\eW>4XU:(N;FLb:>5-
9WBa/S^6aJ\]GBX/CRb_O5?37D,AUZ9,M.0TTNIdMHE3b+X6EBN-#XL?OJDBD]/E
Z.+AQ4b46M0UW<^6IV]R_\ME</TJLC+_b/fCFPVKW?Z.MZ]45ab6B+XDI.P->?:2
b2TY01c@6JXP7:XT8TFA-YRXY?#eWV6^Ub)(6;0ND5b,>F?.YX\@aP85_#_MDCHN
1X-T+E82g7gEgQZO70O7:JF+1U&/Z_[[ZX_LfB5J0P))#^<V6aW+=Eg:5cP<g?00
Y@UE3d)BFF[<QR>WOP6PNYUKQf?66>(AHN70XHM<574.1<G>X>.>M<9DF++6LKU,
N34cU>@=4&9S)AH:Q<>0B^]C+Eg\(M+9KP976_EgG:R1HS0#cg(\;@#I>O#Q+aF]
FLCHA?R[]EQ&]KHOYa_+Ub&[KR_R=JMZT&KEY(e;?P:>;Sc/Q4b2IXOR&,EKd?_+
KaU#[\>J9e8c+H-8?RG?@031M&G;&RF/1L-a#9g1>GSBV8P2VGWRQ82AFe1g&)2U
F+LQJODQcW,8#,856NZNV#2(HLg;]4d&P1cK88aGAA.GgP-IV.X_:QeR-&c>9gQ=
5gSCb\0agVO?DCN8&+aLWc<9[XLeDL34_<_WAPQAC?00c=S5#e?Zc^1V/DcR4^NI
VTT?T?0HYLJHLNd_C7PS.g]9Q(W,].9EZg3;0Z_M@YKAP,(e8<F6e&K+;#?F7faX
^>B5@6ScKV4ZO_\U08/^_56+:/&YH-I+eg8DV9E.Z]0>6g7/UC@BXOW]:7AMBDD8
Z7WZAT#\X>1W,d,P_a1D=94[RTOPPWUOHf:M?W8Z3^<\#=>0/^T3ZU39]^_8@?dc
UPg4TbeT=N2<0SRE^PA[T[KYATeE;1)E^-<+P8^J@2-5YQ:CT<K4fZQd]A:AEW+(
E0GMI\0MX33.]6=EDM8>(Zb,70X]LbSJ4),^1g@U82[9,B=\MO-9/HLgEW)FSBAD
\O50e.gPa<A;6DL#QG#ZE&<IdFd_X)[+C+@/7c1S;147Y7Qf<,#G\#eQI\ebQZ@H
8EJ7/-]\.U?C.@eBO0C]0Pe\#(BJN+fN.^MDP#B[=@&MSV,_JNgC:ADU)9BgIIZN
<L#A,1abS=V/UZ:XJ:B&D9U04F(;#:\D\/>EaaX:1fTJ&Z/9PAb,QHDV?8VD6eaa
/E;@_gFE2,Z77TXEV8_<^TH-:&AAb[U/[1DXG#EMB/&E1.4B&\6eZ0]>#XDf=/f1
fX1O?9[O5b)g(G16NScE]O&Z,3ETG^V)TWaP>fPISL-@?O:Q07?6=)3J51]c(WYC
&\J^3^TG-?7X)XPRUg/-^2>C:J>O19U-bO]1aX&bFc14>BbK5FX<12I\AN4&f=78
fB],+JfOZ<6\@1]:)TE_C]\e-?HF]fBWBJTLFS1D.faK@4U4^Tc@[[IGF&_9(AFD
QGJ#:1g1Q>WQ1?LY&?11JA<95,b><2bS5ZE=JNQfP]&MGaVU_31VY-]FbZ1+A=,U
3T;_=TVfDU\UYK4JI7]@,bgY4A_P&]ReTJO,S5fK&<>-B-.1TLOI.;&ZJa]R.)\P
:-BcYYD3R73<:[@e;eY(MB]LHIJ7Ye+-g+,Ga590)[-Ab4,U7CNJY[03a=>0BM3>
#.a3f1;C]&)GY>g]48_U>E)/4YgE#,[J^R-+GbE<U<].aJ=H3<2N_>#=^I+]LM-b
CB&TBbfNEGBd\WI3TFg4Z0_G1DL?PS-fR2b^&HX?fMX=F.aY5XY:CfS^Ba9e](85
ge-4gOg/_0FfGd,GBO);fNUT<.;XCOS+8+=?YQ.G^@F-2<L]R5R,CT:<5_X)/gQR
4J0)g@?SRgAEZ5gKRJd+/BA=P.fO(C4a==g3I>.7-P:aDHWL9c37Z#S@f/LP)C@4
Jc?8bE9IH^2/a/:EIWe,9gDF7D/fXcF6RL+1G/@\LfR0d3[S^,3P3-81c^-=ZHHC
DI_eU7#gbO=R17CKY^RF3TPaZQ:Ed.JZ<6XUN=;_9eR8^P&01.6a4fJ+ZL6]/6TE
a<MHWBMTH;^O:E_4;R4;UPB&XYAA[FQ2F+5E4F#JSI7g;f?aE5SF\-7+=4GV5Wf_
YbM&-^4_1-?=G9G.#]:aIRMV/D88:Y+R-PeD=_/V,c+,U&2D(<G0GA?+A[6ST<)\
a6&A6Ua3HfNf)gaQ8b2A\C_5]^fBZA=+[(7>GHNVRCg.]c<OgM=&Yg@G=@_+=cTN
DVUHfLM3U?SE8J-#A.[2O>,:3;#Fg3FgRd9ceLQ-M)EVLR4dgVA)R&6A)0HOKWAF
A1@.ZWY8/MI^RgI=VVE,)ccb-DGI2a#G&9UH7MT:)c+LT^f)O9)]IM?FTNC7(PTS
eRB9F_TTX28&H/WE430S_]7QZPbB(Q7ef><T(@84F,EQ;aUf;[C5+,VL4_g84(M>
NP#46;2A70Jb=c@P_^TZ;W[-F=W]0U^-d0Le++Y&\gdAS,+,fF78a?aK1W:0_)I9
-0P,P7=AH?Eg3_eX@[G6N;H08G4A;ZDE#;S>XN]C8IU[BN>MJ;KO.-ba;0\-RS8b
eL#:^)_;gH:I:#@#2P]]:W&N-&V<<95&fd\;;LcZ1DWb-Bd:dfKDd<XIL>^P55\+
P/9aK@+35X])]=#^@P(KdYAT\##I]ZF0)YbV?a&\5+^O6X5/c9M?cZ+TQVS64?]-
MYbD@5EL<M;XN:gIV=/^M:QI[#&0L<;=R5;331.YD?_g4Tf09ZIWS>N=GgfPRY^;
XcA6TV:d-&Qg8bIS>7Q/b,SbU.AFcXbX&fWGX-BI&eK^R^+FeKJK4/1<OXB#DNgC
ENF>)^Z>8?WTMbN6WeX6-XBKfL?DN(cb<]GLT+IcS)8(2,(==F8bgJ5::+,71MRG
(0_T6I<Z=D\aM;CB\P&0^(>-EOIb6H[NFK.WC/5\KMFJO8(Se^4Y]QG[Oc8W12a1
T\IN\5+P(P>21TLA=bJGY2B:46RV:a7+X,f]6bL=+?cZ&A7SN^a=_0F^f1+VI4NZ
8(&9C\a[6\)5Q^@S>.eWF\8ZIATW?EZVCA:ANP\=gON8f-EL;Q.5DD7H6?(cLgUf
+=-A3(X]=a]:0,JF,6[)KPb&]+==_X/VZPQ(-O4BIN/cAHM^\K+NTR8WP^A[?#dL
_b:5.A53R=O(\Z@?HH<d#+@F4UP)#:WA\54R=1TG?=_:g=7XQDYf4G#O;ZX]\bBS
N-]T>&46[c+-0:EBERA-.a4AS_ab@G)E;D(.?_RMbDQM=@A-@cP3[7W^G0S.f1eg
_;1SI7)Vc?#[0&:_@JeVO8HT^#+[.JJD(FY[8A9^353WK6?MP#:0>e5-[_H<eVM8
],SPVU=LV)0>8\gSWM1SXFId6+D:(OWP_TQW[TDT6U=703Z/\Y/)#H]gg=:,5JLS
C@&(=JZBQVUHMEQIQA0d(<N]bP#cRUHK\SJM5\0,ePdE.SU@<<F_15^P&[#><Xa[
bbc96WgHVCTYZ)AJ>A\.g]1eV9dTGM35/B^&DQQ+RcA5#5,A&FT&M+5cWc((MU;:
<4U8IB8W9KWcR:#39[7B+CBH-GA<@1O3<K64LGVF)PeX47HD[_:?e^e,IW:#:?#F
fJ]S7/P]4>?0KTNJdSAW=(C>V:+<<&J12Kb+\//Nb)EWHU805R&DP&aa;Jb\K=#V
)TB;QZ?Fd+B>&d:#R9IP14CcT>):LN4EA1@2Y,Y-I-.<?Z+cN;#gV#13:g6T?d6S
Pacf)XTd7Ee5FL7>6N08?AO)525a2;Q3YI;@LHVGPafFKaD]G5[;AN,,^AX\JX6e
NQ@:010,c=6[aL6X_[OEW-f^LP3F-Fc?@gK8E?MH6V9QP[6:&6O(-@D:Q?=O3?>=
M8/a\P0_L570?UV(CZ04J47IPfPVL^6KRM(O.X/5K/XK3.].297BX6CSBUaGEEW=
\8TKdb?A2SIO.85T#dBSgRV2c&f]@E6>B0O74EGO8M/Dg70FH>T:e2b68Q?L-7QW
YTWSGZAJI+H2cIAFE1HOF-A7NMW5H;[LUBE_]DK8;PYTW[V._JTZ8eC8A_=3a\8:
@WD3,#cZb^-3.4\8Zg4LDb2_8M_3,MRS]RW+]Fe-La07N/[+]g2WA;;4>S24gedR
9ggdL,ba9F^<L4<Hd^OcV@:=a\UP0dJ)-FCTbBbYM=DB6,AAL;]7)]56M\>)aZVU
)M7^ZQ0:VM1WOVR=S6((I:MIJePX0C7^\6,+1:;C@b3E]@:Id<R=/#JRD/SY.02R
]QFB#UaW:R>N^^-T017.=#[[]RNBX)WX2A,B^R+B&Td4DEQ.#>bG)V:aU]/P5(?X
E@4VRd22KS>&305]LP4<]Oa@Z[IMM7U5b_c+YCL1,-_FIM+,LSZ8M:5cQ\Ff=^a?
00f2H#d(((A[O>#ZQf?ZRYR.eBbZR5/P(9&UQ&W,WGR&9ZdSN9?+]UY^O^eOO/+=
@+JQ.)R51eNaDI\BARYS@)B-M954DU>bS(RCd:BEg4Pd-FXefPUKL6CH\aM>\I4T
<(_>7+6L_WHFC+,WWg:Kc@>#,>WSQc?#LI\N,JDAZF;U1GKDR^Pe?f3U3-+G:D\K
Kc?5(c:MUJ3cD0HcZPg_J6d<YBAe,=CG7ea^CL[5P/I/+P=XOdQ\/EUYdWLc<fF(
.Y5.)bW9OM3g;S<Q9GId-O=&9Vf^aa2VBccEe,e]SIC4.I4cd6RA<8@U8<TH#?4c
H;VH_Q)16YJgFQB28&_G.aTH79U:\O-,7M=^1cc,JeXC\QN/,f:GP/D0C(.#b6O.
?:;@FA;7;,dS&+C,gNZJPQ>_)>M\9J)2/e9<M@#/]_PXTQcF<9Ua)+X4M@d/6?X]
__7e9&(\TTbf>+KQBBZeWb/2Wf>TE[7+dZ/cJ7Xf4>X9:<AO@bB8(.WX/gaOUP2J
<bYL>N.2S98@D.@Qb&;S.g<3D90_9T<M[b/)E\:F@:5+TTScZg90,daV7+deCb>a
]b:-?<-1?R_9:?KR-bG9-PTGOK8;>cAN>X?:RRZ(ag6E[;2AJ)C#F&BY_K_@^Rd9
1(WXZ;02#8ZW<)9H9d_VXWC\7.d.PN)IXec,]&03T]B6U3B^Q<,-G3J+P[OBJGR+
Q3aaUZUe2/?FT8XH#b:g@<.e+IcIcQ/B?dXMgd0bYd()1A&S@Je#FEHB1=X1Y-H7
fS>ZT)ecbX)WH_I^NQe_Ybb+bYL4TU+4?+Ne3#,dU7O7Y;@)O/MHXfYbT^J(FFCc
WB@Ug39WXL)P=e;d/UFPH=ObNHBR[g&7+].aaRH#[9>2QB<TTHNf2;[-WUeLfc1V
4@2a3[N^T).\Q.Eb-L=0AaIeYGdW[[?BGAXS/C^J3J4GSdM2,J-Z,.;P.9^<1Z.Z
)f/SeX]R#/7E4IJ/2?O#XAM:6P#,.b+#b(1^FOG.DXGIX=Y7C6DY9T5)YUdIR?&9
EPgU\?Ld>S=Z#BLS1Vg&\,L#R-W_5a^(-c9WT-O_;6^Ka@6bML__9a/=a=SOdbBO
WH(5:@P+DaUE1#_F7=LX(b(._F0F<I3eP>b@<H4Ve;U@WWK.#Z;=YZR)M16-AZ-Z
/>EU=A>4+)ZHF#ND?HI>?>NV()V:\18/=ec#T>_1K9d>C/gM(16ULS7?Ffb.YgEG
-1f_Z-RXfBE?K59f^+V:J<aK10cUIa/9L=^&>/PB34ZL\KTK^c=/;/X<Z;<4?IM/
IUUb+#XD;H:U@bfCIQ+&c,,ABcD_cJ=,.YWA3<155MN/:/7<H@d5+A<Z3HH)LgZ:
2fF::8A^Y9c^X?VcNQ?5Q^fCf.?DPKW4)3R.SYS52SO\V.5V=Y10B.K+WW(@(CgS
H:(M,M0&SJ_N<NdV74SM+#W2LQ&,_Q#gN(KeK6H7?J8g]8U#&M<_[N@FV2KD9K8W
#;bXC/-28[B#>EM#UV>BLK#ag<GB5^4Oa:L=0)^=YCGbZ)JDD_[1a7#I2;fD)=#L
W24aXaTa><AYE\_1_#gdc1<Y12O;2=J3be70d&P=(73-c&NNa#[#Q&fB?=[KBIPN
>GZJ1A_6UR^G5C+C;HLT<4f?)=>Y>6]94RW[.geaEX7LGb=?-]AZ;[KHg9958cV2
fXUa8Y>,5b#g>,.UMF?)NIb0WdL;ALE&O&_CO4Z5._gTFdS4IU+_;bP/[7?\HK,+
+?)6NR\2<.M=G2MeC,>6^d&X4[:F>W^Be[)>T1e<]d&S\Lbb1U(HA#&T)N>MU(9F
dY0_.^0f./L?-5KcBB#eL[M)cY5Sg=1NR].?-V6Tg_e9?g>H_JaGH[Z+20GU;=:9
8eZEI8W=@N3X0\eOTF;47]/#[D>9[-41=P\e[a1AZJ5]]VY<<MeB&^+63d2GXE78
Z2>2VM_FcGbFec(VeNLW:EIB3KY05_KU?M>6(8-SD(9Og1cPe:?a:f)<gK@@D8B0
PZM_:H;E7c=CMZ4MX=DRT]OOa0QOEWFV59V07Vg4^0EU[fgf?O,gBLR:T)JGfbc5
676V+91Y[4YE0S06G>09-7^W<W9gV<aJFIERe+VMC=.,<2W/D8,U>YLc(e9UeO>Z
REF#a&#9RM,I[[LEBH;bQG8>ANFA>&XL9/^eZG)_M#K#dWb8;0[e52/TVY>/-:]e
cE,OY#eA+Ic=->[>T)XU;FXg#6g[9(1CeJ:M>b;JEfM?a>9aSY03aL<0<.FI9dDM
H084a2S,;R#+=c3MZ:M8.1,R,W3VZ_/]Q=@5S(E4B@W9BHWaF[85_/4<HJY)HZ)@
.R<@XW9>TM55aF4;:&S-FT,X..ZY7_c3f82=;/0W0RU=@WVHV+<D>LD#5[T0?7eS
<-]SMHecfQ9=3He4Y@b\K?L]/VYM2B?5&b.Oe(KTC7GDS9a?RO@\KV0HKBTcI:BE
\g)^b]@gb5>D:Me&IPU3[[Ld=T2U>KXE_L6fSFX3gA(<S)Y?Wb9ZE)DMQG?\.8aZ
PD5bTF8>:B9JN._N3Y?E_IdRAZ](=LPcISWb7SH_0Sd=@0_e4::9PcW,\1+_A0eT
4XUbb12EE40R]D;.5PS&fNbA8W6MYcC<>H)H<O?A2:L,26?b[=5Y<[^_<SI^@+T:
A#.-RGFLgV:5LbS,8Lag/AWOff5.A1E.-3<BJ0E^P@@=(M7HCE=fb8=5g\(8f7K=
f)aMLW#3X3ZYGWJgYWE#+DWe:bQd-dNNW]J-:>AEEaRILI_C>>:[++,[D0>O1,OA
U]]?/FNaZ-MZ+Va<42?Ve&86/Nf^<)NcA7[eSg>),#G&2642@N0ENPINKL63N@P_
CEVC&\@:+M,fCd?OK=F/>>J>G,,J-1d&4+Z4TFU]IXaJZJb8^LGGJPGW:B2\-ZZC
HQI<AEg<GT6:&[SdZALUU5C;XH[FQK?,)ML;,eTHHHEV@]/MR#)fE-<>7L:)^E8Y
6+IF/44#/5O(Pc[2XS0He@D-)7\ZIb/9eag4J5-/+JJ&@=M9TL7M?QcHc&M>=)^^
)O/<HFTFE865?L1E)8HPMg_Y)+#TF3LP_V3#KC0GEG?+-G\3g?K\(@QAH7N3M&(H
-YI&W+NY;UFQ2CcR[S@C)ObVaG03Ma2#VTa=B6:\U)=Y6&LQ-5\8F.a&<(LZ@W6Z
eDE[B?SD>cL>TOBORMUB\fHEPb/TQ2PZAEO]YZ\@V^RU\B]ZG)22Tc#OB[V;@Qe<
(-=R].RTG8-7bU?38K3.8<-,B@?TK0U8CJMY<2B1H.X39L+cUTXC^ZYCGFdGCeT2
RW4X57M^69JW_\S=H_DF@,[a7.E([O<&NA@Ub,R-VOPY:YQ8e^G=RF3BfETc.[>9
c=,L-R8F,^3Q=W0]>&GJNU2AW6P7O,.:FOQ_/(1D08I)V4UM.GU]Ug:W&5fbda7-
[+M+.CHa[@TGKRGI8dd6_AQd5>JCBCHBWY]4VJ3DEQ3<KQ]+H#[,VBFJA)MJa,S2
XO\NX/<INce;+-QIbS;PT&C<QPTA6:,,RNM-W<:YKWT=HFOM4;D@PIaH]0bR++&.
6>W-O]()W?BB=c_P[Og;(_R+R1A@8fP^=^B]gf9X/?aLJ_^OS8V;;9.aV,^?6\.&
L;dK#J@N<9;.G[OJIX8?72\baMB/?.Ddg[Z/.Z)5Y#4;[78QLWcWDe1WC/O,BB\Q
52A6OFMKNH7]O??WJ#DD_fe2cQ3[\PS8;Bca(H6fF_[39[>aJ=7+J?\ZJ3Ce#/AC
QfHb3X8Gca+TgDS\gd4A?ZH4L(Ic7c(UJ-XAJ+&[a5@g\F^_;d4:M.fd64[:CNM4
Mg_3JN;0(@.OX?dBJD?2XD5SH;]Vc]b3RLe4Ag])[ED>WKeb7DUHSHZM.KXU[07L
?0];)Q,QgKfa41.)dBLFKXRFB>HM]gA;8g<X0,(0DZ28LE7+7[<^?J_IE,=:H]@#
[(g&Odbb:N;NK8LCYN1E:ELA-Rc&HdPc-5Z0_#e6+6EHO^\9.N)#bgRZD1&6YL1W
0H^8>g5NTM;2_@S(&CTZ;5))>6QQQ/c]+UgNbQ<McfH)<2:WL+^?BdQc]BR>#+><
0^2Q))B@F;VeIdO9MO#/]BHYMCf1_O,,7f9(IeCcTAIOd(2Dc+,[f8fQ?8JEKX?c
\WQZG4=@dBO+CEd+)&4Rb:U)>K.e]7\.W_NB5@e\O?^AIZ&&fRe(Y]G-),B9GHIS
H5QZNJOL@<<GT0Y]P3]dP6Z?5BSBS=(J#.e2R1-<47dAd-:>DLYI727RZGC>BadD
DVIOgR8d\U13_0]K8>Y=V6=UDF?JN02d1:;D7DJQXN?N2\f9g+9fEH?JdbEb[R-T
SQf28.N@[:JX6?.1N:B@cAS;K3&<CEGKB;?6&&0SQ,5FGC,GIdLORL3(K]MSW5=I
[]]>8T#Sd;FT3B#@QFQ35>=T.eH>.8F\RA^REDA1#-S;5KADZ2Q4??K]@OV8N2Tb
M8WF)GH<T7]7eR@H-/PSBLgZcAJM8+ZJ;Y&W0N#W:J8cW:4g=[@aR97b1V]\0Be]
;.8CG)2/RY2OF-5RBUDJN6.0I.GZWB[).-X:QA8IW-B9(H&?2WA_797008FcIV5;
NB9_1JP[8;fW\V6N\a9^+N5IE/:MNWdJ0H,+3IT&1J8\[9(320PN>YJ5AT]A7C#1
PPG_A&G6^dQ64H#T0=N/@JXZEX8\<PR?@[VJ0>b=H^W_eHM?L^Y:ReOcVB5323Wg
.a?88A+e:N0^;+H4gc1cRG+HW(VPB:#LKLPY8)_K):&GZHO2U75(&^N]VVDUGBET
;,_6>Kg0<eJ6/#9FQ5?U;]-3E^[V892Q/^6ggfX2ST5M)YCD&EXM4(RO6+F7\WB?
Q0]N._5T#OS:K(cLE8TZHQPY,S4QcQG[^KV--#W=9dE>FL-TASH+2TAIbgZHQ7ZW
5c0F.;73@OUSb_)V=LH6c;@,JR/O];/7?U6+c.B;]79#&2TAHW:c,LW+D^F<cW#d
FTU0EWYR<G@&G4#4YQ)HdUVNUYLG<IHI;?7eG&gG:80]IFS099QR^7LS2H/K3Wg-
0+.gC\QW+HM<J,[4BG#?2[\0W-KHUTX?T7/-:/dKAXME5MOW=gK[RJ8-?g)842HC
e,2RL;=BHJ<QfEd[a@E1Y5f_OX\UL+X?W+c0:a?g&7AYIb/dKC4aW[JP..ML\IP&
BV9R]M9NRUcfaM:^R))_QU59cc<HUe<aQ[XGO??XJSe\2AG^>4BLB5@AH_a(2PaG
cDFM7dZ,YCGY_Q]5OQ:)If4^>Q&I-#RNUb)CM_aP=R<0?)3+6J/&6B;d07@H9G./
+5>000BY6/>\39dT2Z2;XI7S;CJ;9cGR<GI_g#_<#cESWUPU[/?U197T.TOQ9<X_
ac#]JN(dJ.\I<R=Oaga]W9Ze^KbD@88UUSAU2dKG[U61URH86ZTLVC>S?>Y]WSMQ
;+]1BMOf=N-.300d\9f/f+g+>9bfM<<XKX1KcXIQR#?YWTdQ-I&&3MU3.4PIO68]
aJB9WVgc>,4Lf?;E(Q^DJ>1N;\8<D-,M#He>=/8X+[A7WTZVIFfPAe[^UK+[A>>L
G(5K@NgJ2J4[2e(C+DB/,8AL#TELBBNbGfIaL(^?IdC&U:(P8GRDJC/5S=aA.,.(
H:c.ZOdR#JSXJQZg(PH^9.@PB_C\&Yd>QaG4W-bYH^3H<I7WA-GcEJJZ8b=PT3K1
G<7A4(fJdGJ:7DP@>@L-ETb-&dffW9WKA9Z6LT4(A:LM<YQH_5Q_:I9PBL\0bBf4
gG#g#NH5eA0TN(&O8Z<g6RH#9:Jg_8a0@bOE\DN[3#VA\g)_]AXH.IS;.52_[H[G
1K9(?-cg5VGEgR0D+7OVNF4Ja:^)-0^N)6QPXDb6OL=MIT(U3:4O0ggADGDTY&[V
.;X?]Y&gd+c[P5<E^RA2g<90I/J/8]C+S05^^0:#@#]MdJKH.[13>#^1TA#N3ZZb
EfV0EEUd5.1SG_>J5-+N4U8afC0/S-f3UR2X=/X2,?;]G[-FXL;^>A=-+,V)H,g#
?P]WG-2XG<4[0&\;cP><ED9(;>?G=^a3dF(7H,?I[gbfLE777Q]LS^^2/\5ED#4e
+#(IZENU,&IG?FR(&@\Q:F&Ee5X?IEB42Q4U(HKP8ZbMZ(^N]?8Ba[Ugf4U<[)ND
##cUA(RRATY[4U\QANX6@YScCHJ@,MA9\A0d>D0?8fRXd64=8=cH>5BDNJE:XR[8
8[C;ec4PFf.P;gX<^,0>\J8YQ5AQDVfO6Wf0-<)CISHA_QXL<H/cLK+6Ree[)bbO
ZGAQ46>N1&7BVT8W2cBDR)KVK[HKGf(@9e6,Mf-3If;;d8,T[,USZ@5ZeL;F>L;&
K^4?bTZF^NYO4b(Q-?7+-J10LK4.#QQW=L2R1g:\1FMH5/Q=K]4M\@Ue4()Z9Z0a
dJ^-[7T.TS0OU\aKTZ0A^Qf:d#baU<-13M1-Ze?7__<6f;dF>A#-KU.F\[C06]>&
NRV-7<U+KJ&8[,J:[I;GN0[OO)dF+..,D]A0X-;OS](L]@IH.1N]=>K;@2RT=E^6
,K##-2Z1Z+;,6VG^dNOJ#G937MN)g0-0W_.>0_/4=^[fCX+A=OE<>XB\\ZHLdR<7
1J0,ZVLS9H<SOgWKIR82G59UeJ^cLPRFJSZ;36+7AS/;_(9[/R+EB+1-_QgGN_@.
8[X)YB:)aSDgL#7\698_5C6b>P;8+?W#08Z6\&&PQ8)XU[d?WCg9cPUE1[/F?]Rd
G^agS8+@090P)222#AMQQ./LbC7#Y6-PeND#F9D4[TO,_N#^>9^HVJf7d:Rf6YQe
WLNR)P-P&]Lg/B\\-6)b9a[Ia:)U;>)9/Z5/+(&K[gWIL,+TD@=I&QH=[X>>e0S)
F=c1Y:H1F95/I0F:@0V#E1X#\d?N.GR_FUX1NXFAg&ZZ#6FREZ7Pc^d+6^).7.;3
7Y<&^Za4G6T;-3>bc(-#+O\GdMTMQ9+Z;DK2e-K0a4A9ET_@gZ0H(3,X#\++MNPH
5T9_<IW5HIZ;;3BV[1P>PJ#7;a0[dZ]PH:C#U/,7[][)L#5BE^fQDP@V-UJGb9>+
5S5MX.2/aZ6&8=D\7J,g]IJ88WKAc7.\XKZHVDD\OU(=8IV.OE);K=aH;20/a9[(
0^-4S32(7JQI3B2S#\^AH2aC\3C0/C;7:43UTe,=WG<IM[)2)e4>29_a.T0XI\Ze
?\Le&1b(S?029<6JJObZCRc.gJSc]:C[=D/1e3?f/Q5R821__GY,S_8.T(g8;\We
?PO[407FfFg8V3_:1]2A010U&fR2[YK>D)gX#I)e\F)#_b+5a96REH2[.12H>d=d
5=\YSX?&FL&.21YJN;.;QA[@/Q.c2I&0SP^V/2Jc3f\[1(+_g5L^QP\WIU1gC.Pd
ZeaGE8g&:M@GQeQT0WDTE++[Q+1ESMIdU4S_,<=@RLH,L5/]OIDG\c5HQI2IYK<b
]R>>FC>KUU)g\OG7Ng_Y1J]=XFXMY+.VBDVB#&DVF2Ce^Ae[[^g8>FZb+F/],Q52
Mb6W1+:BZDOOU@?+D8WS=gB[/Q)JaF\/RaRaDLA;&VEOPY&9R<MQ:JHSA45ODX2P
J\f6JO1eg(9,Nd)C(VMA@]B;&2Xgg/#a(Hc033I[6JYY&QF:-cXG-KL018XJBV#d
a:^b):0K,(-J-?FY>2[eYO2-I5eXUCW1A,(VQA=?f_U&gVZ?42.^BUc^EQ?BK=O\
;.Dg?OdE7Bf+8DBWP01?f@L(MJNKH[(VRA+4]NCP1B=O^E)NTGS(bWYOMP;C;L4A
OE.H3N6A:<A_2(1<SU_0GSRM#B^8#ISg[/[,B?dKg4RC.T7NYOAe8E9P3/^3dX06
d)+c/M[GXL4)gM,52QEOM#RdW/RX:S,ecFeWN9?Z\4]?\A8)V(VBCT&M>bBcN]RV
#[W_,V(8Cg,gB+\D84BSMS78N;UBOF,O>I#--?[Se>6,NV2-RHQXPH2NDdJFF-(g
,T3(bH<86egb6_J9@UaD1Q,V@.8M+1)b.[9MH87?G0M6_VQEW;&7<:JY;#Q_L,MZ
757V--1eQ\KXJ9dYdaSKL)14#[e5I^Lf-+Ia3e4];)>Bd+FR=2XgM:^F70Y>03=5
)1c;<&b[cB7P:+OV#)<,T1]fVC&gc(7]bcZEb=2VA,GgQ&+&RJ8PPW2?>_D?H?RG
N)[:LQ;W:.)N(ETZ#0Y9Hf-,:JFJ?Ofc^.0F4/GDe+ZU=9D]\6)1?OG?=0<ac9f2
SgWE@_WHY3gP?#@?,/?[Q5_6OP[g+bNAf/X4IQ.?dV?IK7gW]U21&FD@cOVdJ_W)
BI,J#FbLA0;L^W#XO>FbV1_1E]JJW)cY52]Pg;]4)WNcN8-?\Z;eRRS>F((++VUM
RF=CcF.b[08^ZHOf,@1(adH??a,WHECW=cc/74N7KL0;#T2?5@-#J8#S1Tb=gULJ
/YK>a&6VYbT@)gg+I&/JZf^-^A&>#PN9T8VJfDT,[9M>]e7?Q\f&9#YZ\XM-XO[]
]cJ.W/LP,+Wa/ggKU&WV)],\#7OIeUQcNAK5MfO66-,BX?#R4O/f-:=NU>XcN5[=
@KTLY(aE(WM?9Y5C_T;.60SIZbg9XBNg<C/BX#[<4g@#FH:XDQF73+81b9#9AJ\O
U/4WGAS[.Y]?S@E0POc9>6e>:aE#gF/-5b/>.]@&@ZF1(DX(YQ(T#3#eXVY(f8fd
Xd<d7,;M^83&3^Y@3\3Na0>e,;0V]bEQHK&RWOa,FGAd>S)dSMe1Y1_1LgCfH=O[
#-..TS/(A^6D5T,@/0PZ-,[8B@L6F#I/34TQfZ][dG2E]Fc>O@O=QR093<9IKc]B
W#0(HQ8R);1.H/?(d[==MHIb,NXL,:I5c(-E6.DHfbTY<>.+0;/YU1bKE>^.:7aD
dWcXN3>4f+VNVFY0]_L(S(SPHGb/^/TW0eXe:MYQfQ\J.#F]_U>QJ6/4>I+Yf8K7
@(#M^ba<S>QH:6GR&4OP[+[,b]3=3#[&>X5#9E:B[M67=FHR?W-TT2\MA6HI<[cJ
N,XYU4O-CNB-=XFb)G_RS-;0a5(67#a+ZP2VKb,KW4T;9963^^E[Y2C^QWZ_,&5W
MXLCTbL\,JaGc)2+cK9:gUe-&4>7)MgLWIS;._U7(<HdfE;Q3D[RY=B5WQSITb?E
X,@T8fVDJfa4g#IWPK[Y@C?:g+D]?4G=M+W.M^(4>ZV&ZS#YJg<A=g/BV5+]>I3g
WC<LJ@-ZAHS.++Td?CDE[FPVc;3[IbK27(_-R;+5WJW,Ud.,c:R28M0dL:T4^AHK
1CJ(&TR10(PO+(O]FUV>Xa[bQ9>KY<]\8DfP796SZM;&N(\c_BF+_X@?Fa\.;eP-
+,;]V\_Wg7PVTVC&M3M_FeGB/^MO>04N;;->b:I=EDa1&gALaDT3)[1WEWRc3EZQ
2>;J,&0C(:.]9cb2@-5E-[@&THD]Q3E-#=Xae3U7e5TAG/I3bfF,]E))-Wcc4^dJ
M9Z^2YW^+3W=MDb5IP[OBaV0c5KKO3M>BZb]1H5#IfKf:G_AV-e+VOgU17[ARV&<
H\QUJ&-)eT\+@-6^S=581-6\)X[@UM=BA]77e:6:4Q[YD9A3R@dT1H?QEgTBG.U3
Y6IU1\=#\3;-R/<[16CKGIfI+0:8V\/9(_0g,ZQ@]/fBL.CgWPI6(H(W<]a<gTP<
ZS).#[PPRO)4-S14Z3QEZc]+a;T:TN59EF;J#TYB.d;[7-D[d4XBS:9I8C2K^L[@
bG[(OK4c8.TJ([=Y[X@0GaX]S+PX3D-Fa^)?RJ8D-EddP_-[7+A-g5P5GMW45V#,
cDXSB90C3KQK;?NKEcPWM?1KI(+:a@&CA->LYWJa4Z=6KdgW@RQATII_B3.1;R)7
DT3E4@IHU0c+1+gVJNeIMU2-0@AM.;1Ze&.Afa=e,Z6a.C0cISUWX?(6-S9=EU8?
f\[7P=)cVJ@f);@bb^5BI#W/-PW:dQMD:W3GT/aSX)d5.&:#AO09Q^MDQ/5\;.g=
0?>V7>RgF9B466@FR>Xa6c(9LNJc:0<\b-2ROK9)?PV-PXV?#>LdP+8d>9H3D-WI
U13JV5XIRgWc388:Ogg,G&&dLDD82#NOU07\3CCE?)<0^8gb^ZYXBGb0P?B&[C;X
>Q3b9KUWJ7e3IRSZ&F/6:KT?TJ/g8V]7FGId/N;g3fffBJZ801_C3bVA2ERJUF6[
^#V1=IH-.>,M.f7>6=B_TUO(K6YG=)6=Kg\L[5JND)2(VKPTKJ1K_<_d6Ma[R2G#
L;e2I0Jd&XV)#<AGAADJ=TWR\R:;QHS0dfM=@2IfG6M.]bYOVULK=8Q?KdTJJ,13
b#V-a<H^\5<8&FZf9^)I<30>I;DeERaV2C3O:R31Wf)HH&1+=QM(9(cbYI0;)OSY
AH-QO+OUO8WOdOUZE#SCQXPSSW/Q-U51;W.JIK<;P\_^TRKPQ_.,eCeCfNUZN4],
WbA_^/\PF?D_5R>[UAN2DB4-COM>]^0f^/^VX03]?)3N1[#G[eN4FLKIeY(Ybf0T
;DPN&HVR[B1MBJFK^?>HAIX8\_SG(@E&e:b7Zd44)0ed0_g@N7a+LBM8:cfa;4F[
a=ITFJH.PBX]@fY#U^6QLC5g?[NfaNdWD6T/2U+FP+W=#?E1Z0)889?7:Q./]9=f
g7T.(UA]XUM;8?Ufa+)MHW3C>>&;PWb(,5I,-<gRDZPU^^-N^J<b;5cAf_,.2a1+
((bcAGSa2M\f7O2c)(dB<W81H=GX3g1aF(B?2aFH7C^a,GW:0aDJ80>G4\V:/FPg
6MRY\C3GAK-8B1F#F5(>4LE:B1\.::/UeG>C@4;_>)1G(L&9HSZF&]-#)9CWO3Ve
Q3#CIP,LZf\I=HNE6,5Ec/XY(d2Ud@5VLVdbf8W/Va<<e2EF9&&),);JPS^L;@[;
cg;:IN6_O]M6dgAM[,gS:R4BGJD>OY2G9)71],@#R3-I:1M.NN^dfI2R@9<Fb6,?
]PfTR;:^?3(6]Y]fC9OP4>VYJ>Q99\IfYNB0/@I45_G)R[2AA_/?DI/UFD1^?>&K
?_P^DfaT6=NL=&Fa9_>:#VJZPHNM_F0;@0G65_2#NaKe]Y3-):?PgVQ7F2gM1VQK
P>U2#3ZV2U<I[YQR-_WW]PGYVee=+^=+@&@Je@YQ-VQNG+W<<P4<8c@JgA0K/L0W
09(^[6c4M&PS:2O:0H+(<&f&9WP;4WJX]QN)VaD_4M9VcfM445[Y_1>\8.S26Z(O
&0eD,T.[5a93>BC<DUDY/g/#EJU_(WM0(48KFeE#c;7/E,=.R7)(&Z-8bSTJI[]^
&@LT@MRQ6M998f3(JLM=+,PP7^O.LOI8>B-XQ@ROd@Cb7U;4d]Rd<S@)bY4ac9Mc
,VJK#1,GA?.LYcR]5[CB[8Y+_O--5d;@D[+3CRZ+;)WE8X,a]@<BG<SQ=QFU\NQP
V=XRI=/fYBKG;34bdgGId31bW\W]0?>0_T>WDK43(5fb[d]U.c[<_WCMYNfK9P=H
X#6;SGb/&RR;MX#M(U(/S:O;=1MMTc_\X(B_+Z#17I^7N8X:XA0TDSP)6ZLVK<_^
Y3ad9[3ELET(fS^6_>]2RT7MV;//-(?NP78gPD_J5IWIXS):eM3RHH?0N(9+)c_f
?=fXc/ga-I,,J)P=b2G4G-&UJ1f#ETSJ_b<]Z))g<TXgd0X[V8.J_MXFN.75G4OG
H^8gR>g+.eD#S\#31D?-NV;1P:]FLPYL/AQANQ8.6aF2c\H&]A@\N7EDGKRR1PId
@S(I6W,R/)gd2cD6&aWfIL((BI4P;+-e0f7YgaIc^#V3>N@.915PC6eY)DMI>C_E
<)c][+,QSUOU+Q2WK)_;INg30=S@9HW+/LI2?EUE:D?/b^RaI0JT,J/>^YQ1CS\g
/UIP=QPMGc7#E(aXXS&9S_HMC+d>>O0SCMFUAZ#E9U6[[GJG(/V7OdITW164C<Tf
b@HgMS8CP6L2>b4;c[fAXH@-T[6JZ1/J@V9V2c[[?:1U:Ga(fb#3RM/,\Z)C7PS?
[RJE(;F]046cc9G8-M5e)O\(Q41F752:YDgIf-\(LGd]e7[,f;,PU.c=P58GaKbC
8EI?ZS>3O(;AF8AUc42S>8L5Jf;E2/:XY11YIBN(@ff3J=19L(EK/F_Od3(7N:)3
@011G/Ia12/AYUHK\@W[KZ+3g@9+PE083-aUgXY&U+D>.MJK+R8@A:G(ee@+U/W>
Y40:dDDW]_?;ZGK@F2[3X1I_S:.[_9>RE2C6<5dFI.EC:_FHWI1#S)4(4;UKG/,&
KM&3\D+4L]gcL@O,-\e\g#+L/H26Z_F7<W+&;>NbX\@FOL.1,YT-71+:<WL8RfZU
,Q=A7<bFG[V-f7Gc@7=ge^cD?2D3g.IT6YF_.KPJIC98U:0.>VY08JS<Z6[8F[3V
8:8B)]PAD9;RCeC6Z\Y-2ME)eN&^7dB\E(GA.[]0\X=]:@4)HJ?Yg:W8R@\/MXBO
8c[@V)HEcgc/#gQ:3-<9_2=Zf@7E&;?Ya=+73B\dYT^LK]5KU^6>(?1R3=/2>/H:
L^TBJO<fUdP\?^4UONM^PXIDAN=aTc5VVdTT0IW8RCSd-#V,10XaPM9GJYOI9aLP
>H+BgT:V51bUc_FVO2_[dG^_[gA91_9VT#ULaJ_G?U:gT+I.RC+XH6]TNcSV?C,P
7_gRQ8;-_;<)Eg]>4WGYONa0IHB=KJX1)7\4@>@E[dC-]WGg3-O.+C:FV?gLSG)N
G+6SF.TC,;^+aZ^2<.b#M6fQJMCWZD^Z7MdM;/M86E5H(XELV_&]aQ6)NDN=+II^
,g:7ZL8(I_e8@7BgQc6g\H66@cgEb9.HVH?+c87<VEO0-_?W#@A1/4b5)4?d)4)M
4])g+VMG2eY<a1\6PAXZ=NbaVRADBGf]g/9cZ1HM)-PGNc(//+V3+25;(<(Zg0ed
YdP)K@C:G+d;UNIe,PdQC@OF>_^#;TX7DD@1EJU91Af5JV;.XeD#d._4G#+9YB8N
8&[BV+V2,[E-IWMZ4aCYUCSUEA=)/TdgJb_+6GP-e1VEd_U9):Hd(]g>40N-KKW-
V1USc86([JO9&MFSFAXL13=6@?_e.K[KdDE0[0)#IYLH<+D-+)VR(#S6F,=d=3\O
>)Q^Y)M8KFH]<b\0F74TIVLN>a6K_8gC+BM3WbFBKgJQ?I&S2./>?16(O+I2A4+\
O,I?^@H<(>fL0]2GUGM9ZWAEPR1/eKCT.T?Qf8C,3[:X1E4JJ-Y6aLC.NcMIdP0S
CA2S0c);f\K6GDd0UF^O.9T@0V9HB>I,g=c>2).f8\7]7FBG;b);,c-NKJ;Xd3N<
_:e_/1H>aKgH[61\c-5^Ca@=BCbGF0QG+G>\)4/(M03RESF)R(Z3FC5Uc+:TNNgK
;L2C+gQYOaM]?20LJcb(_gcf31eHAc2Y2Y?A^()YTZGB];KY[cOFgNVW.FQUW.MO
4@;;47C6)PG1d&Nf+O=XR>9C-5JR[2dA5V3>X(C59VeIdQ@Q51eM[FWg)?UfQ8/5
[0VeFJgYb].03@5Y7L?AQSI;ZefX7NQ;2)14Y#aIg4\-7efG109JSRD)Z5I^:J=&
:M=TB2Z_).EZ[)3?;-)^2c/J01W0V_aP@36FVBT<NF0eHb+^/.@NER/QG9-]Oc(H
O(TO+PUBeY1RR,75Gce2+O&Wcb(3H/>THI7RO>3&772VD3L<L]4?5UN+NKXa2I5&
LC2Gfe,dL50&SZR\8#?8LZE-TWOQ9eDJ:?eKZd\GL5]6N<DWbeQ4@=:,^U6U4S/2
WKA3U]<&L/#>Y+SK=7O54=HZg4YY+SU1]=&<>L;:/KBaO?BSYV]=f^AKY/bALZ<R
\X2=U+fa=Z03?,8dZeDDR=EWD-(T1GE3Y78A<SHIBE..X=X[0+\\K4=-,DQ^cTBc
EV:=?(:;U;-]2b+5.],-f,A)fM<1&1.02@B>,HULee^WUa8(7435UMFCF\C@Aa7e
7PSdaL4&Jd>P<;gLD&Had4?QfJ?&cGaU3LXgJ]K^^IGIZVd4a\d)R2>+EDE)64PN
?94/3bgBOIgaW(Y^MWF\]f)L]I00c@?>MU3<K2;9<f[Y=^79\8C+>B[;C=T8bX4f
gCM@8<P=Z<Z9=aVXT4689EBXA4e@FVfTYTAVQB@WQ:eSA)H@:KJ10A4@)8caB1?6
OQ^F]G4+LgWH[dQDRB=6-3FC4?TSCaNKKDMaT\aHgSDfZ3gI=agaed^9LgGWF^]H
QVJ3RTV)7W[+8X]Q<fUd+7X9HVPcTF?F_fbgbdGTME;0M2T];J4)P>M39XQS&\e:
0JgfZ@<);=aEcN]dEY[]&E]CeDAYFa\([4IE2NCR?2b8JQ\C=DSO<fY=bZQ@4KML
CKd\][L-_:HPGf.P(F[E8^E))5K(+G)QDgHM&+P2^+#I\7>g?V]LT=(E?1R>]f/&
YeRZPS5J=6V_K+7HUFTbSf#LX#VW9<+.XMA)=FD\Rg=ND/37KgTPa5\C6cM&9^W<
=)=.WDJfW\-=_;a=&\Y:.VE:dK_S\5JNPYTPO^KIK#-&&?a7Q\:ce=:fXNGc6DL#
PVU#OFdKbZ(Cd2&2a.Y)0;&.:\P.B/)0PM^,_H(f&H7D]_&.K7N0EGHUQa(N_5;X
E:U2]FHLZ5D_?bT;C?VdUP4K6B(JFEd3A/1_[8Ja=2KI_U,U5bXVTXA(cU(2QTFA
ga#a4VF#@O&gO&(c7FZ?+3^90R0VQ_#(?&ZBe85_X#cH-f:W]6YK5f-C?:;Dc&cA
VWceWM0&41:X9;MV7R1P9\K&#0K4^dZ26.+7f_?5g3/?_6WP3\-MQU/;DZIdE.@R
/FR#TOYcfKM?K)<<^>^)KHaH1I]G2Z[(_-4\A2TeI/4ZaD_WfL=0/HX3QW/<&Ba#
@Ib>KZbd.7D#a62#<+1K80_NSKHX;Kb@R.(,?L0/QAe74=3Z[3^g)M\8>M#dR?+7
UU[C;&+TJe5^W_<U=a):=:^,@+S/+b9EEY1B(/01SH?(#)VCG2JdBJTU[Kf)HG&O
.+B?7)<.EGbM6Y#IfF.C-Q)JG\3L(,^.:2J;L?_7<g?&J5fVJU<1H6a6_@_;9@#X
RFKIbN>&-Q^KC],1IOV?&3+M:&S@=4Pb[f<B<gX^MWfX)Y-[STA(@&YSUZFI?JOg
Ld):KWEMF..WP]_\#<V0WZggM>(/YUZTTb?GB@>.I2/?DUbRXUee;-P(@d[2UaPd
IAJMPBEXC6ag3)Fe:-[cZ03F-2[b,0>fIY<XR68=fb?b=^[5bcC\Q2/[KX+01;96
KEK/Y>F=WHa+<I=R3<Ve[)FWL?4M9?:3Y-RCWNI-)?KD:?H6:0be-]30O=/L#GEG
g>I1^aa-)e652FY_2N[^d)&7CD11]0bQMU<6&8ATO(]#86gYLbG-LGEVYMH+feZU
HM;(^])C?_O(/+LU2TG3T6/\E]WWZ-.7ZCcC.^]>HOJRMC;&Q6BbZ((=eY@0Def(
^F28>4OZK0D15:>?d::),D3)M76,g]U,P]STW6S>MEGZMGH6H8/?BR?/QG-UOY]8
U+8MF]b6(0DF#HI[Z@805]eaH(@F^(BB+5LNR>EBE_c;,fIEL3aHB1KIV]UYSXCb
eX+/R_?DW+UEY^7L4gG-ZP/D1YeTP._-^dQ?K;_TH\UFSQ5Q:NA50Q&N=2-DR+44
J8f\;GECZ^1&/(F>)0S:8WaVW>M;([=QS=A:MF>X/C4XbTU?^VfTf:5aN-P)_=F?
d8OBN77d+WH)M<b06\=?KP]0:#P@c48NC1\<Wc9YIcP(8\=V6VDSYe\@STP<X4;[
?5M]3RS5+fNI_dGUI3B6Jg9\AbGcN?7fYQR6M.GcV^0X5]S8N;GSS#M8Z8fER=IR
;g[N5_WPUUcG&X4>[bRa+[PH?I0)/V.(3._SNY8&C343KLH-9KB0K=5M:9b(a,eV
ZPZQ>(H>9UGb&C[/Z9f9F1aS^#YZK\K>DI9#<ga;?:BbNa[TeLb].?[Eb;a(FS98
>+ZC5:BM<CY4#VM4)L(;OHUg+Pf.gbH&)BHR+I-3;L=ffE_&;&W3;S&80-9_.P2U
2S49d,SYAZL;Xa.,FUDA,9Fc=bM52I.=g4Z\Z<J2+Sg\9E><;bIUSXEg-+L72GSL
=5M&.fBZ\]&UO^TRY>X0;9[a3-R:[A,0<3G,fP,&?4]WHHX-1D,G.:X./OY\Vf.N
<dC+S:fN436QTfLSFRb90Q(Ac,1d7NcAMbN)cPO.^Y>c\2f6Fe28e\Fc-S)4VI0T
BXQcV0e20AB^;77B>Q([b^Kf;>MNB^+5F:0MNLgP2\)PIPRW3I<U(BbB1Kf[\N,\
#WBQZ=d\:B<-[8Pc#6F./_BRA#>d98d/=_GXNF+1(6_aM,C2[^^.-aIHDN5RH]#.
5>,TEIKI^9e60C:WAeC(FO(=g6-UK0bEA]?:=<Y;3e@1L#S#QP,4#-+F]4HOJ?GO
Z3Y@W)G4AGZZPC3/K13G^N9S_CO>eGQYMc0_4B7N/IZ]:bJKN;a8_XeOD(PA?I#[
_3#,5<BHCSc7P,)CDI2P[DWS5gB_,FCWePN;d(I?0)Y:^C:S\3K0bHH(GaN9/BgA
;TBH]G0eU1,@f1B[-4dX?eW/N;5=CXA&G2bIc?g>[2382d1bRb^E/SPK=]#QTJ4b
DL8_P]bVBe.&feIY)I3&B^LS>(_2P2K5D(D]]dCAI6J>ZGRGXN-X8=92K3S7H-HR
6H,J/09CX:dW\6=>I@=L;;ZRJe.ZNMBaVID@N3aR#J<QcM2B;?.0^M<8LfAW\L=9
Z=K,0LM9X&])/6<MYNA-=@<Q2^H@NZ3.I6O?;2:[L(U@E(U7<PA,G9g=:XcLOg:]
5D\c5&(5dGG,6EDS+4TO.A(QBTb#HC/=6[@>3M,PLUfOHK3OR;?-75MJa1I9YLQL
Z2B984F=VC3WZ8G8AZfM0_W391S.G=HX7(g+UAQ,bJ_\16f0TeH>S5:AQL3=OOH\
DK;Ge<#GW,T33@:@2[YK(XHT@4NXBWU&A?f54;C41&/ZBa<3BUMFJ.^1aBW#b82P
JWO\+R7_/R#a&1G2Aa3HZ@QG;_N,E>R:Q3/<-aS?=95W:&)?D+3HC.Z&gBA>6\+I
HPQDM^bSYDKLD/D6J-KQf3)Z]CC1IX2-QJI@LV5XO\9Wd9Z._Idg(>2P9:M4#6[J
bN6]85[GXS6G?b7c1JG<,W0EMeV@7O4I?@2ffgB;28eY;[.cL(:3@e8S2?K-Q25^
)V&/J9T/5G)R;<MgK./<Q_/PH-\IR1#cZ?(<?=.IZHVTKRICC]b;4g_^f1Gg)^RP
56<Ae_-Y1U07);<9Lb-dW-2G<g,=V?B1SSN[.A\W25N@V)AJ.^Q2GD-JVM_d@H7E
[,C86)=aQU;U86&?gA+b+C-KFE_O?NC7TW:0]3492(gM5J:U)M[YcT?)S?g)4d]?
.dEG(9I<ZAT0BTdISUgYVe)))S46NEgIe5:e/Qg@3RW>@=SDUO6fTc?FDSPX]JY-
K+6/X.S(SeQ3:3:\3Tg\\_gB3bIFDQGNACL:C.f-T\3UGV#65R-=?FKKK^,:-fb[
9R@U[?36abX=(TRdIUU=#V4C_W;91#g(K&KJdV5aPBf2I5c,CB/9+Je]X2&BDc/:
&E59RO9g[YQ.[A+Rf;X4(5e09K5=PHMKP?@JW;L05.>J@Q9UW<UL-Q3(J?>^fLW<
R-&KL_Nfd1)CZ@;&g@FB1SFWUedC2&a#;@A/9<3BDC&XZM)ATb6d1O9Y;7-M5JCZ
+QCdFdX0]481QL\\87aLS9f&RCa:QLZ8=@F+8/&cN3g;AAX+(>V0<@>FUN6/c_EH
SQGB[NL[MW<)4VeF.WSaI.=R.1gS/4KaDCJbgM&8JWQGC2+cWWf]Wa&=4/FZd<dO
>,2QHeQT]8b224Lg;I[WHVMCREA,\+ab;CJd(UN3L?KM_dIbV2Kb.JB<ERPFXE/>
A=5OENLa?ZE]G?<DUfcP_&MQ>Ec^>+UK7\?+UE1Z@Z_&<T;eHHHgZFPO.YRCRa+?
\PGIC(G:ARLM8-GI#)+],CW98:)861]=359LIUAS[10:[#7VP:gBK)fHXV;5:NP.
0PI;(N95R\F;Y<Q\\5&cb?0,5LETLLb0bJ,][<dWNdQ;X^d5cE1OQ)<W<=bYdOAR
EG/8[JXRC85TUP<2bf8#\2WbSc?ZWg@@O],b@-4RfEY_]gV>dZ>(;DUN]@f5+/^1
\^-:_)G:5^J)>(@:.eD3ef/VQFg?eg@aBeSS[));/4IM2B\2WcOaMdG->Z]C\1_f
TM[d/=(F([f_MOW8AVO[GE<bf.)??SM:I4D#8@C2(TUC4<[(dY(@K7A5=3T(66U:
/YGRgdbDJCYR(b^FZAcdP&g45;[@>QR?FQ@3.P_g>Q.JF1J7/Q/8MUHCBU<;7C=_
\Q9(VP<LQ7&HBY3?W;-.EBXE/#?6OFe,b0[&WeL6L;OcGC2,/#E?Jd@9IaG#eeNT
S&\<8WD9P#33@/g)E:#\d?IA8E87P&R1Z-DBH;65b,_+fSQ1eF+Lb^91V#8ZA:,D
W-NHHB7(Z7>@C-.GL:b6W3LReL72<16d53db&=/9BB+@)4X#<77401\#P6,#/:CV
L++@VLCc4D,&LV1(1E-HSKWDa^=-W8<.SY9#ZP-G81b=R)=c,7\J[&bXPgS]a7b=
85XQG2V=I00;LeR8@5#-=9J4/?ZD4P++f+MJ<WH?^Ze.VBZ,SG44E9RT.]f)>F\T
O2Wb/_1c<Y?\4aFOZaGW0;g#2Y[)[+Z_8ZeRU.M-:[Z9d/+gJ+YgPJZ==OF8Qg,+
CbYO416MgbZ0I_88A#76P=C&RV@#/3bQPP(bB@;=;8bdR5HegUJ1ZE^IKbN5g0dN
<,ITfX#AS]aQ;D<O6NKf.BPHDD(=/-H702=K,ZKdS&/EUf])--DC4N+VKaO,2NY<
@bKA415/a#b9BJTK7?7#Z/<_3EL3HB,@Sb=]BUWMbb6#Kg@ZfVMJgSF-J44XbZU/
/;ZD[9E\Q=2G)>\=H,_4SJ2K)L00@>aOdCB1-UYMg4@2U)^[OcffCEDWbQKH_9eJ
-.E,9&&FLR1K[@#KRMDHB)]&ZD.O/FY9WC&aA9[NbgB:bcEga9KBV0&9+I-<IKa&
C]cFYIPM+CYO??>5[aPf3)gL4@/8#f\HV^7MW(B3^[Q966TILM/-NT6,I&T0\:RB
9.(UI#f=O;Q28MG_=/\LD1HF:J+QJJT4JZ&3GVBXE>F]\@MMV+1SfT]_JXMKBBdb
Y@4\2V2YPDb=O-D\()#B.Mg]Z84LR\Y/VSK?9&[GLD10BCRcReb_J-e9fI9F;1gY
;>:::;e]8c&JUQ:8TV0KOJ>#+B25^[]gRJ1g/>f#+T8a8.D9/PB_+C5+:S/K_#]+
8a#8V2&X<7]@ROX(ER^/1-P3&KbCBeS<&T(=N^JW6C#_f7=Me2]PcYKJ2>T7G\MP
SFF6.g,R6:.L97.Z\d&@&bF+;CXV;_:HFOO=>ZGY^>V40U?eK]2fKI7Nab3QQd@<
4#[A?,5)E^IPQ[?+Z9e1WR6WbW1g2OO?SDCb=.<O[II8JNQP8[][,)/Vb]1B<cIO
[PefXbGF@R)<LIJ#?O6I@))+=b-Z8_YS9Q.L?/0Q^SFX@JL4.DC=O<e(^=YX00T.
FJ?1(eB31TZf=MAU)]X\Jb<8O#L?]c#d.2\5?_,0g4M)&LLV=\NNJK3OK3GbNN,6
]>NI,;D-0P6&==V:I553ISf)>AI5[LF71M):dfU(E#^P#E?Z-.^@+R,,fV^1-LHY
=32VB)bL6>H&_XdGB<aZ0W>OXGZN12+[c)A.(Q1GUH9^Bg:Q,#P3NUe/d=L\4aCe
\,?(N]9:d(F3<IHZ1eY-&0eMM,\:5HYNX8TAc3C@Ea_DG/]WBF<E(dICXgX9VPRP
7.Q_LJaKVT]ZbQ6@<N.L@I;03Y[Y)WFa#K&J:ONEf[]0S+][?VSG8;WC,8Tf3_/+
1;4YQ@80;?>=XDEa-a[77-\(:P7G#R#RS<^d3>^H;6JAHDT222JEKT#R(0GYU;@;
5?2A[L53HF;KB=AgV>d72H:N[+H)W/V5\FOQ[VT#&B5A05]]SI,2/aZSN8\U]&7c
2Ce^VXO1^/D_[GHM/5fD__.EG9F7dXX_K>1?BfAdE9RP>B2GSQ,:5a&&M/0^fcD4
JC2#(O^abIa<X-L\&<O7+;C?3Y?.c6DV1W1#.#F.+U>8HeEJC[fZT,B;<><>_)_Y
(1eT8C=^_D0\5B.3JCg)=8.>YXa)J=L&NWfA>P6fFH-OAO##8\FO8fR9?\CXAL=b
79^?6eXIC8ad8+Y0F,/OeUCV7HV[D(EY1/\WKPg]YRZBZL0-I@<I36UNdDOXE))3
W5;<#F7E,HObR,-T\RF:]3Q[<bZ@5,A1gL:f=\608YPVaDV=^#]QT;.6)O;,);W\
TPNYcR6_+F:A_XKA#SWHG_7N;W@H9N\cN#T^#MS.@aPI+793dVE^2Z=?L_f:=IEg
C>H+GKO&fLES\ZcTB-:_#KG<cW>2,^.X_]dEWLf@_;FC/SbQ/gQJ=/3.+&2/:7#.
2C.WOU\/cB.gHg/\b,GRXF6WL.<&U1eR^Z<<I49X7b1.d?bK]ZIf<8^(XPD_EZM_
^G0T16-@2]OIbdQgPee4>fW&F]RY:RP;B)d\E/,W1KKSMfbOZ(@5QeZcEa1/WdF4
)(Mc.2:.[TPQ\5dFWQA\L7+//B&Q5ZJfN3;K+LV7D8c<(4LU@]U3/KK]>8d2FHB:
_:Q#RT2F2YAJbCaT<9V&:1KLS]/S&Ca=W/YUT\RC^g]]CMYYUeS;#&bZ&X&1BZMY
DaP,O_#8A7X2V,DQ+VCVeW9I&02;//7gWHf;NcdTc0=eI]7KZ1HC7d1:=(7K@f7R
FG8_Y(O#GD&Bf=;<BXKDP7J7dL.7^AMC21A0WYB>>&NG;?MOA&N=S8YPcZ\ET_]\
MWE>;=U/1RZHf&\LMaDDHDec;4Y,+&D0O@^8P#CO==g,T?-bI:#D6>8a[_d9dAZU
IM1<CJ7:5TY>LO=cT0,fcD=+ILgMbB;&Z+;L/4#U.K(\@dGEQRM5V8L1E@D-XBS9
/??\;K/K,>a4g;M[1Mc22<?^BJ#W,(&TcY^?\X1DcYX.0YH,Mef.F_F6.X>L+VK)
CXW:Y/\=,F/E#IFaU-KSK0B.\=TP>>dS&4A(4(-]ffLR<8&:O=OR\=F_W7)@<b#,
8Rbf5&HY4WWBT+/YgJ<_V@8&0DL8Z?@:I_eR\d8WfaY/810L;FKKC7?K1-JHXC\]
^T#C4_J/M\C8IS4G^+<XX[VJUTW8;O8-g^eT8J5fV3U(U7XU/_-?gf>TTA>G^S3(
CC10>7#/\AeD6d.]9B8P/dOOV06X26Vb63fYVF4QFCF0,dW/dI@L6]>^NE(2].17
eD\FOA/8b4^K\EcfXdB5RE=2GU\CdJ=#(8Af<5:FM;T1A/M++B+0Jec,CQXFWH6F
ae+eM]@6R#b:-6VD<B-[@SP8M#MJ)C<])dAa@f.)W88?PAGRQDa6e9U,G@<SD0_b
?NN#&eC/6<BXHU&KP1R]b8,#EJ\@S7Q6C7=,7A.Sd?#Q-a>)5GL=2#_R+J26UF/;
BP@\gUK][PbJRBK=e7b?\c-c@;bQH;&[=Bf6O-_(;d]2-GM#gW48fgYcD)17BFdQ
c;7OPBg,a&.5Oegb#B8XbFb7Z[GR_QaaI24=.14R:?3B5c7KT<+gWYI>TE9&,(ce
4/+)EE#dS9K6:36:MN[V6EVA>;Ge7bK-FdSa\QQ34g?NRE)/)_6)e7_UKCeE3ML5
;C2d4&>EL<;[B5HX/3<@-73g+F@9<^)VO1SdgSCPKBcX,05@<594RgRE_?cJ)=^,
.)beMVB4ZB,Q7G\&-ee^F:(K_\VJE2P>):XO.VI,b;^N>gaD,_EB,#_^8X8.O&]^
\->E+G?WgA<1UCE9J^E)f#FS-38)gWZZN,1?c)9Cc1<NNFbV-TWe&UL9X^a1d.3e
C7\X?c^#DD.UC[4H9&&F=QP7?U8RKAWO0V<F.VX:H0=P1N)7M38+.#gIcP/g49(0
DF]52Y&g=7F.20L310G4<I,PXW,UZ/=M.T5ST.g7J#,Lf32eLcO\L@.JU5DN?>(>
9^(MS:gK-6F=7,g<=21ZHKFWbC#)P(PRdeNL0I+b]HF66IF_+8g1/N?M=\BY6;YV
1SKV8.b8NT26b\(=USV8V&BE7C&>[a<)365B1];:.2e12\#]]df;XWH.a[4W?_&<
8A:_+A3#.VG>+ECN&d)-KXUb4=?FC416(8QY)SX^O[I.-.=7(N]2FC3.P?GYI&[/
Y_\>a>9N]=aX9ZT>eV\EU@098DAgOOf[Lc?12XP3OT/,&HCTB6[ZcZ,:_U.4V)9L
b>2;A5:[,T4(96XL-3fCcPO/=N/]H+GV8H/[dVJZ@a#KJX\[K:(Z[KF)1YZHP,;0
])cVN1#VRcGJ&P@b+SHAe6W6J/(@0WIGV;L[)X[Yc2#3<QK/^P5N9IcKJcB2,L5&
=A8/Y(0Oc-G>.(]F],(D@_&6&cL;V1c0:LJRIQ#S+YUY,]fXCPX]RXQ6/P37T2>H
E.bFWb<e=\(cf&70\e(43\5;2:(T6YdH8EfJeN^(b4gb;,;1F;S\0RKH]3a+2Q/C
<D.#>aU)\gEM_aD=_HC?c\WP=-C\JARd<f9;fFB#6H^9gKIAOMNN_HN3,R[geU@W
.Q:4+@,1R/?Uff>K-9FB-:AGgGGPd==HA-Z68f2@Xe)Wc[0^DI8Lc<Y&dNLJGZ00
_Q4RV50DIXFC/-K6KDYJ=>]f&0([,>=PTe)INSX[H<FPbBHLUA-W3/M3FX[EM)5+
4aL\Z;QMCJ+,6OB++I/,f_>aPQVM\e0fPT@.]TKT7QL6H3\7Q1e#PSXe#SZB2ggQ
5cH[d9KFWF1ODL.34aAH(L6;&/EZTK2K@>,D_\<U<\B5&#A)Z9.Xf;-D]f#V9B>9
FO@b]g(?>7C_M0\&;T2dDc)_)(>4AZ8PXLf3eL6XKb;E50\fP9KEZaB2:?F7T#+0
Ba3I>2N8=GG-Mc+cO[B<KU<I5C8FAI^GE>(/>2A=a8QE>&(WG#A.[b_8a0H5L>;=
A25d8/<FPg/cQ)6M^#bg@BK&B6@]U]^^<9V>FYBBcKf&V9c-dH^-;8D_EKH4;&I:
_WZ3E6=(SN8B2]7C)83gPc9-3XP#9UR=29f367IK<1T--[^4Vab2)Q\U>b]TE]f2
_1^L@>Ug;SY5C,d_67G?]Db[GS+.+D(cW..E8)GR/^M:?KV1IAe9#[)OBd9/ADB2
EJ3@ag>1D[?I_T<gZX=48T]2Z436O^?_);)G+NFXVZdPQZGe4RSRY?K<.86LffG,
gDSH<-]eG1+QR/;M.._gH21Pd(,=88=eGgF>+\IVRB;?^b/aPdO,<g3YYAb70LWG
O<S:SgK_2A#PeR4aVf=8;(U,e<5QC>fQb5+83UC8,@^<.DZFdd25;FePL\?6EE]4
?0)(Fd,>RF4X67\R5U+K4a_LfXGcCP3KHUXL<O-Af);(4f]BVTNO&5M[4\6?AESf
D3<BMZ:Q?T0Z/OY1?eVM>0&GS\6ZEP1,)df2c):_[^]<HJH[#PQbHZ&SOSP<]=@V
@374=4+)PYH)F9S8TdDg:V8LbQ@AK2UT-??PfW0OLYC3aH_NM0\P,Xf1J+H,_:W;
Q&3ZI]&.S7^]\fA<b4B.5;,AfQK_\I^H:V,7=7VNTDWN.J-NR-dS+LT.STX#9<Y>
9082b.d6d;DPKVRU]]?aI7^g&WQV5ebMKV_246Y,Je+B&WP;64CUHE&GB/Vb2Na7
Y;XMcR(F9JBS+&4c))0I7Dc6.S_@/-5?Fb+0-]BcRe(_4#),8T.8.,D,FH,C.+Ze
_5I^5VT6d9_4eD?0:Z#JZSKOccRcg7Y@7^&TXLY2NCQ^BNWA;PRc_XN+;4c61aa,
HHHFfK^P>I.JLB//_+&1<dNP1-=DK_MeT#Y^D_eG)[3R.8&QRFS\YHA02-eY[.S<
R_W;d77_\LK7MJT][BK7^eTV<P(H^<?I.K:-;_,-e<X[VD#)XP1V8O]^?U)d)71,
THC2B=g-LbaCAU1>TT5T&05)6:Wg8-PXWf67BRF_<)^0GI+Mbf&(PJ=@70Ye,[8Z
\ZR#^N@-\<Q20PN0A4AL6/0YM<SBJ=LX)Ne>X@;B6R3ZWB.#&cRee]TT4C5M+@AG
:>HEcbW.Qa/?JNKc-E^L/Qe:?;UG[g(?&\GXFZ;GbUWYXcL5_T3,_J\=Y+EQP-aQ
-4)O.AN5=ZdZ;(A75<G:0W7Y_Y6S@Y@=4\eQ:;R:8(&A(5,fc-,N;YIbJ6ObQ:NW
KC)ZNMVLVYJ]/ZT2PTN-+\6eN?fG9,ZKNREC]#N-_2Sg-8(N&X;IXe:\M>PU18>Q
4SJ3fII<B5RO226F.MA#G-VFW@UAG50J^1F1.;I=5BF2fFMHP2;Z-VU^7:52#I65
LM9d>FZ9JEN.;<L4VF5S&-M.d/2;<;WC<TcEA7AIWTM1R\WV,N=d^20]3<)T8TU1
dU\1GZDaC_G_A>6aJQ:MPJ7(-=:RA9W\1\P+DF\WW,2;899DXf./AXV<9A3QA5fY
91H/70:JUK/HKT4B0NLA=a&LfEIHfDbDGcHaOCPbI^^N?Y;CaPIUK?E_W1AQ;O)T
;)Y681WdDKEO6.JcQK=4\MSFWQ:)QEYZ+,,\3R5D59=\=S55-,feE__U0N+Vc,=a
4/-N&=A4X+e5>Ag)14MOFQFW331YAbZTC)-6_59R=94.RZ,Z?<UdERC5(BJ(KW1L
#XT0R1dTbeB<=Y;X,:IbbZVJI0dfZUCH?G4V^c00L98ZB735O50?OP\2NPeIG\9Y
5(S;40NATUPdaEQF8+C5(QH:eACg4aB#BBb#UZO>&BMC_4e[.>fH3dS\J=W\-d:E
bC+DWeB[FB6[)Aa/FA^_;-b]J8(B&Z\#FU4F6MdgN4egLKLDO)A-FGY_LCP;3[/b
6H+IM68D_V:_B(\X09O-J7Q#?b@,Wa@,JL\NKJfRHFXZE1DT;6IC203b_N:GX.LK
?@PV+a.9K.2d_;eM2\.F^>+0Ng;13[)#ZJ^GP,98:1fDT/+W3>XSE=##E.Z_e,V#
WLL4-X,3LX&HHX/LGY=fBR/8?PDZ/M0#bK.]HE;dK+L?-C?@LWX1\HbV8bX^@dPP
_=(FX?cGdYI^P)S4GU+N^Wa]\:T^,0H,.[?I,04<)M&)G)B#>0ZV;I8NMb9&f>KF
U7EOIbVV3CC7F;0H./\I<,QGGLe?I#=_-O>:-GgGYZ&eMbe3==WRIO=?B3GSTcL,
\60M\O9\/U^#]76NJRa&KW6:dOBY#6gYZMX0WJ3+6&C&A.XK-&;N5USF1D9VN2IX
=bGJ82PY+ZXb]ab#TM-)AFKHS@=.&K7KJ:N=?J5-4+K8DGLNL^F&MKG]dY7WD667
Y5-cQ#I@N2J67ZRL>(&Kb5)(@)UE1;1.83N0UHZg/(ZfK:T4PS6X>J1XcZf]bfZ2
U:\RNXYZHQ6Y[(4RG9/KdW&K&UC00a.>19>3_E&D;;P[ELTbAUY8Fe/dNJ^0B5I3
9U+A;4ZQB8aYOBQS;V[/54<A3cDZ)_WZ?)A+\=C2G[E;<0T@^#P)Le;&4Y1R+c4O
0U\A=]B72X@&-TWWPONKTB9)2P3A)Nb^6Q(D,81WNG[I_#)B?B7RY93VIQb.]@]Q
;#G)6JI^&[IQg0+EXe(C+Kg#;>Z+10)]PbL&7GeOHa6^7^U,EG(8ePaL30bRdH<8
&<2Sd#UJA39F_R)SW^_c];<D<I&7.Z#B@&RA@SX>F-\aTgV(2V,CF]012]B<I4a0
0eXJJL&7W\geC6X.Xc@<&e)L1YC7_14M?[cgCPS[?VG?0KFD;IC-,\&2#T5M#HX4
e41<^HQ;=:A3a>@AN)60M1>&3\U.CeEe--].]6-(@C7>eIJ4MHg8;>EE3_WdE_Tg
/f+[?eB&#:3WD^AJ1UM[g?Y-eBH<;/,;DDG^/CCW23BT2X30F9Q<MH\Ce6OX^@41
RgU+C=MNfKECbX#?^,F(N@(<V48L5GVIO@:T^81/C34+[C3-/S/:BIO;Kd9MXO[K
H#AOPe>&dNJV=A&L@Ua8XQ&[@9YP0TU])eT-5=#H<ELaDa>;4>fRV86ea:LcNQDD
d^1&,CQ/L79QCOEXUXP<77a5d2AR_DQ+/MHK5(Gb//1=^dS:dRZ0G)c,@d4-?QO/
G7_[,)Kd@(^LI^ZJ8:cfQ,0:aKPDK^BJU;I0H>RX:J.JCW@9</N4Q9B>eLH^5UKZ
1/JAGXIdVfJH?L8?<^Y[/\Y5WF6/IQ)\g4FD;g(AU:=T2?5@?Ee([D&B0NW?WQ)Q
_\[RA+VC0D,2P0Tg&1EL6@#[J_bL<E/4RYIUYBa\3Y.#1LX?#WZR)<23&_I<U7X\
Eg(^O82:2RI-8ATDgZGMK9XW^S<[&aR.<X;a1b=F\?bbK^5OIVXBUK02,V7OYBI1
)K:Q+MP+;=KC#H@OcR&S=G5d0A)(>??JebE7OTab5)D)GY3[=K9MGK=_&JVWNMK3
KKS<e?3bFg<F^.IKJO6R^QJIE_6+_cK#.-=PQVHM7812e=b4&fT,P0PJDUCYgBaP
6/?7?Y-07_WDPgfULQ1LWdJ1,W^;:XU5?e339bb9S]/HRe),b+@?UE?GOdR)_ILf
=AgAH+cf(XP)bU2+;\HYK1A];[+F&0XX(,8(\c=S#g&ULe\KBUK2#c^]UD0K?(XJ
ZXK??+S_4&B0(9,((=]6CZ&71\;A8U=d)^?BdN-TWMWe<VM)\cG2ORHO@B:d/a3a
KN-BQ(E^bILU,PNREP;E>EQEDCN;Q3Eg)P+[=A.)3<<+4V2-8=[Y];UH6B8MI[9K
GK/CO^B>[GM8b\:^D,8#Idc-<):_2W-d@XAJL4B>4.AOD8);HdW@\4KBWPXae;&U
d6eV7),4[7\+HR^J-.S+g7a)PVJf[:>0ROHYU\<cg4BK5ffg@49);-bS3ZK)O<R4
2;VH2P#1;g(<G4c-11YcT7U6H)Z8T?ZDbF\^5UFI0.:3TafO;(=(O1T_NbFI@bd(
L8GPf=I5]BZ5;K>fS/EGFG\bdQ?T[0D[P^U>08d7HTGgQ^?>5/0_NZd\KA-Q4]e0
23aC#b1-A7?OI<agASN68D2@?V8ZUF]fIg^)5IO6)U&EDN[Y,ZH/ALJf+H9=e1eM
Kg_YX?J+-c-6>cVH4<afKbR&fW4(>)HeI.VS5,EO+]dD)8b)N1L8N:P#3^0/H:C-
.NL8LaHP^.0)Ka[bM:df?AY5/eN94]4TE8.QUJ)[N1S=dJ4?U.4E;ReOJ&b]Q38;
I5XX6;N)SQVEE>VH=[fU:533I\OESJGI#,90+[_g6ATV9QRJY1H]VH)gBDU4K4@:
571;EX5SU[U[()[@KJL,(\RKV_0bTcX,IKTE1LNV(Gc;a-aQ]KW1Tgf=g@27b\DD
bRd#]cS.)JFG>&9AYG(ZJaR4].AB_WQC78Z-92NR?/,G2S<-48gAOOZGVLIG)C<0
L<+HI_0QC>@3H@O-T3EC47MFRSZF?F]RP[B08+;=,dG\GIS@0=d.M0\=1c7(VZS:
Z[Ng+d?O_Uf@V:(3D\&a>ScdO8\)I.)f[=UL=+GLIMf,G0gV^T97aK.&4(PI6dd;
g^;L#<a4<cebTZ7<##F(-Mb-ZLEN._b&7_.E#J0Cg<D],#d&S9YgK7E-f6(FTL<0
\e\/<;NWAX3E>I3eM;WEV3K.0&#;_Bd_H65,:&WZ)6>=P1F-Z\1O//2ZNaf9\I84
^>Hd]e&fC)HD4-#b.aN_T4VN37J7]H5PX4&fR,6P:R>dS>dV\SE:=6bY2VF24(d+
-PS)P83JVFMN(52.GQVDLMeYd8D#^LUUb49..4aJWbbANK^2TYX[SgR#<<PN#5[Z
,Sc_&UHJIRW;1T+0KfE/&;0/7#9@QZI-b];-K3/\M]TVK3>F+:]TXe#7E@/1fM-F
IKUY(EEM.@PZK>aZZ>9+e4M&A);fT]9]?41eYLQ4M;[[W/agOV4/@gB]0[05AZCJ
OVJ80,V_DSUc\,^4Gf3BRa2a?J)ac?CbIC#3CfB9(Z#8EEFA1Q8W0F5T7Q0J6[M;
803>&3aM\cV\@JeQ>.)W;G/?)^IND42A<a>ecdcS=JE76=P,/G=Y(JP0Le7eJUd,
aX6HeB5]M+<K6f26#A<V5+-I^T(8[\V6X6a+,@DWdKQ>TR=E@@SK2RM#RU19E7OY
./7Kb_:Eb7R+=MN=TOJW6BOD,_T12^/+Sc1>?aQ-N8+f/M\@QeJ,Ib?\@4Ue&S+&
+GD?]Na0Adc<9_L+)+H^C_+Q&+]+J:+MdHM@[#Hd=O3-2BNJD.U=L/DPJG&+(GO?
)N_c69MWQESL</Fdcd2\X)&C[<)]G=C9EE\:,N-Q6=&IS;L=)H7e?,O<fSE-](SE
Jc\-9ZS#TfZVJ\V9.9/F#_82+@CLO0U87+8T/(R>;:0-T\3K@F3EO0..+LC=P>(;
:[=L1@HfD><<5O/:]bWE=/Mf]W=\Z#;06TGMee)c\\+K9VA8CKc5=5;/GbE3&bJ4
Z@TeV;W9V2BX6g[.\8Xe-VS]/>TB3L@aH79S9McPJD:5[?95b24)1\9._CM_1-M9
d^Kb,L&KWF_5Y4]&VL]NQ&,1CDIS&5-FY;Cf0)1Db030U6KdRV#Y4;-.E]-UdKJ\
Q(?J5@WQ+LPWf3gTgK^O9^#T9>[NMa]-Zb[@S0c>U1\GBQ&gU.aDT6C9,]P9F41?
OF+_bKM@XUO:;9ZfGHUVO-:^C.6gW7UVO-(@B^b8L:;N\8&gYJEcY1WR?5Ae&HY2
H@RQUM82A^:4da>XX08&EG).^g?OS]c7IR\#)EQU;VE3RIV;-;L0=DD8aJ<#Y.E_
Wb?K]=<-&2N:We/;b.9/)W[Xg\/aZ(>,Va7[8&3B\4Q\f]?eX(>8:_0C@QS]SJ4J
0\T&\#O.^3=D1L^]eg:Ff+)_GEaf_V/b\L[b=R596JDZ\C11L1&AgS.11RKG52a8
a+V<TTW3?eb3;U<VI=7=C.(B9JK8?+=,X13/8PE;X8CL.+Vf=dR0H[]XVIU4Y3b^
TT68Y/f3^a^/<PH^=<(R+PN)HKWAAV.+^?YbA3IL0b.2.Z:X=^8gNB0E8EH_ZY-5
DVAX[K.@7K]#C8XKNSMLHF&-EdeFaF0YV^ccE++NPQDZ^Pce[ZN#fcC;12<=7]S7
@5^]63Q.VgG[P[,bOTKgN_7W;?+(cGM,]FQa;c)L#L8/?&G.RP_V.W:^80RVg.[1
@KANTR48eEaP7;LLaaAgc?GCWAcH)S9X8^6W_c_#NAfA&76J_QK)Jg8(K+20eF,:
[bIPN:N6BeR#adV0;[(E(/5fV=S#=IF;<O>WbHc7-3F5f<JNE6N8:U]QZa15U@<>
Y.[[Y#?CJVJDA78eI93B,)TRR_2B\cN,^:+7-Q6/ZA1>3/>DIBO+-HB2egH4Of0W
8BD<5:;4?10_+@&dX0C(/3Ja=.,OF)_1X1.4Y([O>1Ha,N6MfF8O[FJ#A6]]+,+(
X=/e.M&]NDJ8DNNFL=QAgUKENP8(--C_+P=]=@OTXUN2FR>.DOM9c)NA[#Q6JV5P
6&Z-XN50EF@PcI/VcBfU?/R:BFSO>0=4_[)EbF6G3DI0_=T,&[^1bJgdQf=?H8A=
3e#eE^eN05M.OL;d-c;VIM#T1d3Bg(Sd:8]XQ+[<>V9La+95\);PST+f[04Jb0F;
9a5b5VXdQJLQ8(YD99D#=)V;+1:5BSW0c.\0<d0c,SL^)CPP49O@L11=VE?)#+8G
D#^_ecgMa9,)QR^H635@</Q9OgNf2\3Sda=K7\H2DT,D8LLY<fIJ/.cc>C3Lg;(2
,_cgJ5CTW>:.[b69+WCDNH\3T]D)2KKH5&UaO;P4QK@K15GFE16L<KCC7aHNYKS@
9BJgW8#&f0-A3,O:fA@_eT&]dVK33-QRJ.Y4[DC27SKFJ4K9N^<6C^E8T)2b;ZW]
G2+M)0659IH]G#UXR@??ed4Z(+S]AMT6F?aSHC#cR;&He(Ab3^3WWgf^TUX(:NVT
6BK8fgbbZ-F=<-#/f@=6?K?GFEXYW00+4,/L]D7UR0;@.OeX@T\cPMTFMEdHS4N,
Z#A\G+7PQZe3\\6gO1;@)\:AGaVW8Y6acTJF[41^[R@f/L58GTY=U>=A560-LJaQ
aN6&?;D2P2+Z_R(gRdNH(S4e]5Lb_,EPgCE<dXTg)P2^W#9Bf2/\<_F>_1Y/6;LF
6N50P/TfG1Cd36HGX3>f^H9cagJQPL=5Z0g=,\c]J-W&H@BY:WH[0V[dLT:@#5^f
8-VLEB[L/P(YYOH\/2UF.XA3Z5I12Se<)^8<CN4^^3X-JHO)3I1Na+g?H[)#2+G^
O5Y2,IM^a;,J:d?Fe3P..ILOB2+(?<07Mg4X5VT+Q1_^#H3>D5#2MXMb#d,e5?LL
Q.cL+&>7JQ^C[TE:b4S8P0TW3Z+\^3_d^JI4JDYdIAE[T.N6_F.[Hb5?WSU@-7ad
B(RJ,<R=[0\4G7.R2F8)5P4-<-VAOOR4A7P4_]5+T/SBa/cZX(d;<G-H?D8edS#.
JJDBUO2c3-SRea:@DY@-ee\T.APCK4&gdgaUDTcTLJL@D3X4C&6QA^AW)]@aZ&YD
Aa?-KaZJ3(45g+]7XNe7TE>S2Y^HIN^&D0)Qd(R]81B0RNVL8ZID?2OWBJ,Y1>-3
L5DJ5@P#5b6ddS9&<@W\TX6CFNR]HIS9,@=^6@,XG?+=>B>aMQK1FLTN>FS.Mgeg
0bF^40L;N-1DG7#H-[(@XYW/YgR#1_UJX5GV8aSE5[8;</4edNH\G9AeS?L..F(#
ZP)3/@AZ+P/WH9--E8cSfSUG#0Fc&b_KRd-L)\dDVZKIEK9]-LJ6\GUU\,@eE=O:
OAXCIeZO.bU3c]Ug\DI1>_Y=F_&)W1429;2<(QH_YgODPdT-eM^C:c]c2>2+X<c)
SQEUBB&@g?>e;#W[^5?WP5]a-DSf,,\H63gN\=PQPS;+._RP):&L:bJ/)Aa7OPGZ
/,@7)g7H9[BWa==X\^_^40Q)9A?g-(;#BF>aG(Eb&Mad:dPO44LaJ]0&W5E4=^>/
:D^eO7<.CK+.+35Zff]76cARYL6,MG<DTD^HN&Y>6C2YBe\9QZ(c;3QXH4eXK=a_
,K1,LKce4COV/U_YY(KR8\@Id.WXDg9M&=Ua4OV^H0dOE.]MS0Y#IK9/8,K7P6=X
(^fE/I20PTAL89II8UV:CHE^O2<0MdG<\63@X.-cA;VeB?+cLa(:g:&2?FPR#)Za
e#<BJ8^\NXb^E?PHJgHR\2M_@>f5ZO5I_8X#JD]gd3gD(Z0M_K_&A?4V8^CXS;?#
_71e\b9<K,OIDZHH.].)<7>?@O-UBS=#27,[_a1^57J=g^JY8UEg+28FVQ<1Y(cd
b\]VA/6XaJ:LRP5d\&QC/(D3&T6IG)#SYFE]NYC31db.YV-JN\b&J2f+N)X@,IW=
HIbN1KIL5(dM])SWe@cA#c9L<gM;b=V9&:/4eP9]OBIYda&a>MYTNccWZH,.VJOL
[0&CBAW<b5F273BMAI/>EAQH@NGP[:WgMYLea?NJNQ0SYNW/aS_NYX<4/B):^XCB
?##L\>AF[-6ZdcD0V5G(^bIbfW<I;E3XTbD&NL^/GC/Wf)4J>?>P@dV:EbfX9-79
^XE#7JEf_RRAMO\K65#NAgTe]N(&cV2PbKK+9:C&.1b;Wcac<6,U87c&YL>&3R,[
WdeL<-bKfV<^a&WC?R;aeIZKdC-SGCA&2J17Z^)CXXfN6&TRWf#E+034Z[=+H8aW
67O(3-=MO<7>dVCVIZ-WTI>:_)[S.^gdG:Y^7aUFEIZdafX6SWZAT26]^L<YRN_]
LO?c.X(>g3MN2ER]Va)e3C7R0\G0#EP_R<E3TJWS32M+HUWLL7)b]f/I4LGPDXTA
9dOX9P?]e@A06(E]^X]7=A:1MN?=KQbAO3@a#dgNR&HWGZ@3O4CaT;@6X4#:?.,^
VD40AI//FCX21(W6#=bH)fF27HAc?C8,YY74U<GZ4e@K?4[W_?AL+Z8S6AY\<eAK
;VYd+ED6E/HZd)BG<O37F:IKD_2)#Yd5;XG((&+J4J/:?MIaE^8/.N>Q8.2U7DS8
afOMJ0O#)VQeKeYI?IJB..^5C?4f8Oc7bFaXUQ]-CGR=G1T:e[9BF@F4?bN-0?&C
T4K/.7.9&+b_dNB@AITV^C/eH+e0B0T=H1^@)JRa1Z[L9c=1aa<OU[)a<5ON(MeW
2/)c+A7JD#L-gQfb1c</B3OT^F<<H\[(B2)9Lb#gg8e&#Q-JMOY\+6D&dVe^1-X=
UNJ+.\eG+KVNZFDN9Ic713UIO[EL_;R24bCEQ0W+>,5B:\-7_>@.BP^R;./6I(1,
Q6-FbG.>TM=S0OF5E1H?Ng\J/]2G2A^M-,)?]I5=:,5&ON[KK+@@A)FQ1Y-CTc]F
RdQdOO4[HI-N#?0D;<a#X@DV2NO=48CIgN0<<4;J]NHY.dA3fZ>+eY[Y;2-QaHI3
-O-Z,+072P_06S)A[B/+WB3c0OA5YOT+-;R;SX&7KN+A_;,J^Q/XMIaT44I1K@fT
1)bd5(M[^:47-IO#:U]X=SHbCWab3O(;f<fI348.9GbUR8Z8P(aPZN?e,[3.)#b=
Ra7@R,1B>NM7O[C83WRDC?V)K7#E+)0:+&4U>X<D#f(bOZI:<0PDO<ICO<IbJbAY
AJbW9bT7)LH,7?L=c/1Cg7<KM<-&)=4dU/-AbEY8/SLF44CJ20/[c];YV5XAA_5J
Ca&ffF-CN]e0GdXc;g(E1#OD?NU=7]78>&dR0)Z5\aXAPZCEOW8-]eLCcZgb\<.X
^(L)aNPTU1#I;9eZAN(dH7X:RdPG3_)#WB&_EP]D#<b>2(J0@6JTR5@LS7M+Y<TS
302=H;F[=9ecW#1J/H8.XC=341eAM<a_Ac2C]5dbAHX59CfU4?Megf#N?Qgb,M6<
9e.:Z-TaILUYJL\gF8_;P=bM]BBIRY1?/a/1Pb2W=.CJVdDE8cWA&:OfT5K6?1XE
eJ3Q4K=dJe<3bO95&PdD1@bW1>Yf(&;HBK^HbCRO(H3X2:+[=3]<,g(R,98Da>9P
:Q-bUg<>&Yc3gIR9fM>JM+2@AR5;+K[2aE1+,ZIBQ66+U[A^&g55D5[A9eEg@A)#
D_1@E-eAd/5PGD?M5G&SUN=\JCc]UPY\Tf8.FL#5EbL>AIS+,Z2dc-G<2XYg38U_
cbC=Z;9b9])#BFV&^0NZ9O+A.4,RbEEN.2@5f8G[S&#9#^.P-=#,d67N](6]?J;Z
#(Z(29,U0C.eV4gA<cK_&TVcL5WA@5X8Id9<?J9;Q2[FW+(NWTQOT,ZFP;V0J5Ug
#gAeL&9F5X^\cT/:PWBS8gTEL92-H7YPO3GXCI7-V>S7cZS19X_?ac?dE:Y\Ye0#
cd]F4[egAG.7O3[K@aY>R6_TO(Q7=O_bU:Q)(_OOK48A,>V:B?C85QM(f5@A9(_)
1KSd^-JN1)^<#01KH6&P7egeCeA[<@XQf=HDT1OV@02Q]PV7=;>.26\]#B=+ARQf
/Fa6gJ7B6[<3,N#I#1NQN2NY?d>CAN\SW8OG<(7dTaQ77Ig[09\VM6U)d4bWNIN=
2/>TXO#C0K:H0a-=e&/J6ET8CHKC?2N9=<QQ8+eM\b9:_<#EHZ:@R/eGBR3GA/AG
e?Ud-QDG9:We=EC.NM0-a;a1/>/OaWIce+XdRYIA6B&E[F\FL590B-A8==93gIH+
];9Z]a2<YS6+\CASRb+5,,@UB5M_g^GAZH81/>GVW><WROJ75-;ea6[SW3d1]3f)
L,84Ucd4U;TgCM@bH(a=8<<<a0&F:Q5dC[+VNC)I+5ZS2-GG.5b48fI(g3c_:Oc0
)9B3/:#TI8edeP8FfJdT0G[C[S4Ug3I99dO>ZP\09IG2bB-HbZ<Ddc49R5#+d>OZ
]e[FK_7Ld97F;ZM;AEA:P-D)EYfOEbJ]Z5W9L61g.YQZ0RENGH>M,O<JSF[#8AA)
A+4^<N=7./KJ7#D>\MbLTG>^(^^g.@.64JW[M8N##A,bUISY-/e)3#0I\-VSWG?)
&e0&WfaNfeH]9N(U&ed6GbAaS436abQ:8cd>c<G8[K;CMI;MLfT57N1?[gZg\F\Z
489Af#,L26K;Tc=6;DD]9BQDdM;\0T_4Hc)]HW31fIaDGO>U/W+QG@YbK0@@ff(/
dPYgd4/g9)?/T&^SW2;VZ3X#c]VJU]T=19[fAJVKIX>DCEKfV?7X[OY35g],@IK+
#JTHc\Q-A0>(c/b\c/c+&5_57()XM=]4/?=QD1OER,^=a-YfX#1I7OMdVOb-?&f>
<M^W--5A94KaYD4=U6:\eMH:7WIC6&XEK-4FDQMSQ/G+HaZ,Y\P<GT7GV;EgfRE4
2/?\=-A)1JW[T4\\?e2\0_e3/0,4:XX;UX6XEUBA\P]W1<T^GH](?-K2TZ)CSf8f
R?\97+/Kc;G)4;OL;12WCNDeEML/#]ETB#A[G?Ed71,[@_3>V>F>E7;2b?MSPfU2
U_O4ZO>,:1g)0b<H2G6X1)BEWT3U:5K1?#:[IUEGC(0P,T82YVQc,V_6Kg(@X37g
\PAOVPQC>T9]^Kg&+G&c+O>BVR)8H+/2a7P4AHE^K9L1.b/Zc@MQ\>1.&RFT8=:^
fIba]b5+^R+BGe<3H.C.2OA0cX6;fD8VP[6Y\K5@<L>2CQ<4EKH>+d?@02G17H<]
2YG71_bCdZOVJ0N<V-N3+VVA+CN_O#ENEW/#WMPAa-UBM@PF0f+NI>]2S8Z<I&GK
9f<2&3RJ-b@74PT8LC1c]bD@?SZZ/bO(AZfF&GIU_R0CXgIFLc(1S:K@U@@GYYZ,
B.N9OW\[;MO8)bLKM=97H:/YVId^23HJ0fP>/bBPNeJ&L7B)#[TK]5F?P)#49B[O
W:a5aO4>Jc-GWT-)eZaF(<d0V=J[K#]XbAOC]QBU9NaJ07dQb#CM>W]>bDL]3WUY
D)#EOZ6L>6&,fBaY4DHWLT0Q1QI8eU;4#-84Y&:Z&4P4#P];Q<@?Y?88eR9Pf2V7
[V,(@X7A^ZK6:(-&^BQ[^6eKC0=Nd+//aeG8dU[<B(D6g_3MDJRO#YJcK260;VA+
N?8RV@f]QW&]&9KRbJd\(C_JE#aM_Xg##?\B_FH^9A>/HYb+S6Y&_]#a1;.CfR;K
M^cXD51:P/3,[0\(Ca>0WJ;_W((-d]UKd4GI[MLRIFJC&?YL168_0cU\_N,cG27W
66WJ0b)O^3R6R0S0S/K>.<,9<S.DPcPc39J6.R\S;^B@X/fCaY@F,)M5JZQ)EgT,
O71J&cD.C3>K#-TfX6eJ<-UD^3J(#&)#<;-[^WK\^[>3SY^bVbc(@f;X>&:&WgI)
>9G9OIVQbbBO0=U4ROI;0F27@]0DT785R)?GK?K/(O=-;e3,>(IZ8U6.V9ABg@MU
gD#PMM9P=&Y.cB_,9VME.7TS_4L56HcN_[6#3^M&O9EOW5?<T#M?TKXJ3N+E-gcN
Y12^67P-@//&fH;JKOA[:KgLKA:c/XP-=,/KZWg073[)R0AE(RPWcZ8(NTREKS\N
77\BHaa&7-5Ze8VEg__EcQK>,60,N;CPfK_I,C3+LGREBUYT87#Q0^dEV:)X2b4N
PAVP;]:D8PcYO8AX3NTMVKMKU.HAI?(^&Tf1a@HK;Xg;eWADT0FXgKIFG&TEV-:6
LG&F>I@K#86ISLM\_2.I1Oc\6@U)eUM3=dEc^_LH@bbESAQ^[B:_[(X?@,0_,&S0
KLJa_MM;\,CBWYJ0C_eWN.dD_eOKbbBD7?9)]:Q-f+0Z&U:H45)7gaL#P(9@4JE.
GNe[BZ#dJK2=DgLdO82F:?69Kg48S0RVW>3,)-X@><=_H(YWE+dE8R-OP#89g;=>
d/:5TCJG?3BE?]S;E7VUDE4\S7=O:OJJN>Gc&Q+bT#520Ng;#GKW2L^K_.VOG?[V
-(9cXXFb_NE64f6)b:&>?O\48fFTXeN[DGg:Sd3GQI-2)W0&?_O7BH1?ED4^Ca)I
/<8#XGMU6<Oc7QCYJ7:>;<5AT51Q@:73?SFR5?Ra3NE80EY;g/H(a>_T:FI+;:.:
1>d><f6:#0#)6WP,-_(&VX])D.P?e)D=g[9Q?8ZE_94+9bOT:0_[Y_8_56KF92T=
4.0U)]X&)#SLaO>RM>NV2A#WaHE)WVVaO]<c7)5AX?WD?14_6J,ZXc-CUb=H\.=Z
X6cD4RS56_?9]T)@\3)<5?EV@=2C2LPN0?XT_Y,7=UH#&RAd9YFUNY<N2ZeA=;&2
IAN)Ud0&Q+]7T..QSdDNfB]83@S0=++<f(b7gX2ZYc0J<EA=86JD4MP@b&Cb59Df
7JM.)MB/K6+X(M3<#]^5.DLP;aDb.=-c_/fU5]dY4?GRY)H/DTN1AR[_fNdg71)5
@.aWC5ANZ)1B-=J7dFSaWVE_V<-.)M_0((,RFR2.b)^97_L5B9fI<U6G(O9UJ9-R
/(Z63I7Fb=SC<P]-d97S&31HAbKg#8[\/MV(cC&F+Y9V-N+cdO8I&VBKD0)[D4.f
MS01LRbQAL5-O1-1Y@Z<,b3F(dL)15R1DaM+Q?<U(=8a&&AYRMS\JE/>K=EC:H&P
SMeK\H^ZE.a[dNWD8RL69]:d_-4-I48ZK.+@2;WQ&f:H6(MYfF4C;7JA4XRAff,N
fC7G<E,3R\\b=MO@G&0RC3=SDbT@-Wf)K4+Yd0VI&1Z_HD;Ug4b47__923^W;]NB
^&L69^^dWJ9K[c9&X;cE2>T3ZT&9U4?GPRW^&?&KaFFD?Ug(80@0B/F:\8P1Obd5
4+F#+;ES1Se7+<>0f]^-=W,,6YTE9]&K.U?Z)#OW5gP0U[@VK<LUfC1HVQd\CF,G
ge8.5=Z)HJX8B\A;SX/]YO-M1^EVaMK61015b7E-c?@L(,XX2.YA8X17-Y)LAF:>
F_dHId0XK(M1S6ISW0:#Na6bfIQARdaE&&\a>AcMG>Z^UK.RN](T?A2:JKH>@/?d
S&WUX9e58V7JK_/dZ^6(7&9WF\=7ZG<2Z;@-6[C&./J.VHbMLG25;23d^S?CJT;]
I.;ZTG@UIN<d4g79:[[T?>N<8H=H1bX?2&?]B+AO+;FNE9,B#:+J:V<.P9Id34cM
+35PJ>WQb2UII#SKIGf9>[O8N44:cT#e<[)0KM#Zg)dS&UbDZ:S1D0f-.?&FEERH
BU]PcMQIH@#J87K@Y&ZU-_&=S9N>9@\91@#VWWA02B0a?P62\=dH,XSfFS#)>A8P
gO@V:OQY11]Z=5SAC_OX:[6AJU--7ASOR^VBMW&eb/QQ^cD&^AGSGTKe[L:/)YG^
S?:66ZV[\(75.R5:[I1T[cbE;<8Y@RV[HbdLgJ&O3-XBX9MIS<09#UM[#A&g/Y_H
Bc_9EEU,7B6FP1>L>G./FBW<^a9Qe5WYM)>/a.UYIdA=G.C.gc@(D[&@N-[(T=H[
8HQ/ES]QdVX^CY-fbS.CWBC(^2UC1O7>[5^U3T>ge;<NT<gB493WHH]Vc2;aL>&f
]bC(UK(BeSA4(&H?J7C;LC1Vf=ZZL;TI^4(EDR287\bG+?<0JIXR\aQBAWRBECJG
<313:0_41#f4(f^^\.[:3JD]3)=a;U<ZIFNaZMIJSd7;(>FcH7<e/D8Xe_I#[fYP
_AB(2Ke2DB1-W-K)Gd,]UIP^bRKM[+24a1:/XB2>O)M:H+aa?a.NF4N^:OW#3=N=
GIT:44cX.W)0?WQc./;+/B2)=If?.OS;aUK)&Q8B3YS]I,]+E-_35@g<(<Cb3];0
PSNQU((\Q7gS)#=@JEdLD0@@S45,H^B^W8.TKYWE=YPbZZCN><6?;WQYR2=_-<PK
ABdb,6PKK,#@@9P/VAW@Y+K3]-Cedf44XgQP#1G,Y\LWJ9@\G8N\3BX/)]+C^)JH
2KA)WD3e4c[6P)-dJ/4U>M76@f<6Q:GV1bBRW@:g;2YbfEQZSc:@EJ<U^YWG22(=
,^F:f^(ZZ_.YVC2OLR?^5B=M^2A(eJa02b>^7\cIbIFW(3/:<A80U,_c29IN/I0M
9EH^#4FfaF<EL4^^\A<H0Peg;1W6O^c#9RI1;8a]_\[Z</#^7X^dB/QZ+\Qc2^,\
1M6KVC(9YM9Z77:X3BB4f?-cP&XVI7:IKEcfD62U]L5&?FUbL7dA?7RMIK#0ec9#
_IH-&Y57?e]H?G3,[<X^7PVW;@b.T]B3[BY6eI#3ZE>8[5M6YS\([WaBDf\.A;;>
1aM5-WN4L[>ZA?M\@I&W9fV<Y0ZP5#Sf)gR:L7]0/\U:3U1]LfeC5V),VYK#_O?1
G&9NRMc,;XR7L:/7Y^[5,AA,67Z=9Q9@>Y&3;4-[VQTW87Fb7XOMH@Z0CaH7gU=Q
7B58:Qb_6;?E]R2D>02S:<;K.O5)E61,;,Y\gN5c4K9+60<aY-NL:NFVc+&>AbSP
)]=\+T7_,d7GeWV2Q>9\>2ddNT<Y..8/Y1K8SQ0=RQW:;Ag@.-0NH[T3JFQV,JQK
,H_E-^?DX^g9=V466@aZ#3?._fW_]g(HT#@?9X.QLS.5^RYAZ1QOFQ(:/+7C-GXH
e&?C2^FNB:/M5,,_D=(+,ZTAW)QEE:)_1b3+NTbDZC^0N\)MH:E(SG0\H9XFCCT2
??52QQ4,=JcXBCT7/OH&[MUK24A8HeU=2?XT<8-,#N\bL8-.)e?EO,#-=FPNNNga
T5R05NNbSbXK)NG1ef8JV(3O^da7d4^A412e\N\+<L\X\NPN;-]FG/c,F?)#:/_>
K+Y4\Q--Q0=(GN/.UH;4d._KMMP90L2DB;)Ke1?.@AIS<837e&;=c9/REE(Y399/
NHZcaH&SBRJR[8\_Jg;eDGG[&;(8_W\_7+c++.VF@Jf-&LZ6fgM0_XLZ-9O2aD/#
PfY.7@EVeZ,23UbBDb_<.:#SSHTcR1\Da=^a(TWPa6H5A2+O8;6=Y#AXc_b[Y_-=
@3ffMU&DYH=_(EbNAd)>K@\73RCM]2RRF:^g]LX/Jg1M0a-cZ_LN04@H=EGTUQ@P
#Y2^;3>ACSNK3Fa?T_5YBZI=VGb4bEZIR3@Db7e@.@M+ZO]#c0:fM0eIU1[V015-
HOWHAF9:eT?>926d,O7ERDH2LIBO;ME8AYXH;VfJ7?\ECfe:O0e47#[.D,L.9VPe
R?L(O;f-e??4>J/c^NBK@J26.\4+BL>KZa-D^e1GF]b?&W]\3;a_:(H5A0e^P+e<
BD(AB94OZ+8g83NB,6M(^M)&Cd7#aNN,gN;fT9_#Z>M/EK[7)0BM)2T=CCJ?5_/N
584V:(1YHDH>?--AP:T\bB49fGgJ<4_5VEgfVWM/#@f2HfOIBQc9eGUF1X-V.#g&
JV2V-5,:41R+]<9RZ7Od)Q+?7RL4=caGCK4PBH^3K0Nf#OLCT/CH+Ydf):QASg/^
>QSZJ)J36VU@)8/+DVfP3XIZaCKIXRF:K/66K?aJ.ReR^b0c#@E8;9_0C/G+\R_)
HTOJOKXZ<E041]ZN2F-UW23])c)cf]95S\]N=9SIY1(g-6PIP8]A:?7RHX8c(,XC
3bX7IA[\IAVLT:L9ZXW6YefNP0&]_(@V0Fc3F:+-Z#S-HOF);WW#&:6_\J5\\:A4
O#b2;X^aM(I?4/<bZO->_>=VSU:5Z&E0QE+]-\SOVb.H&;CeA.,8Z:bZRg[=6E(>
YKQMU\eT?UAV<fG3eUF3W_a4-^S<Y?B48Z^2#[(8SLBK/f3U?[QIYe8^;MA45K-^
]KLe5.2#5#8)9;LaJ[ST/#VHHXa<@_6>B.LVMHOAa-cD:&PHdK]-gPTG1(MMA^[X
&@gb)(NY0AVRB=DF@QLYAVdYCIg/9^F:g#P,4A2gT]>2PBV]F;AFK#][1>QIe+_e
+bA&&KEf1G<=OCG9+Zc6<\0a;U-3=XgIDbG9gMF_^IM1Dc0_S8BK+#._V&Z/+3CK
E2]1>;5SS7C3EQRI,03.c.G.HC.6P=7/R5?3U#,egY^cVG?#Wea<ce<e0d4aH3U=
_IQ22Q_0FAc2ZX_V&GN#H96I_LY9g\,c#a_/1<Je7gXKR/(WSO^>HQP#e).Ma;Id
Q<TZf@0Da1X9,XFN[E>GZ\&EDTaYY&>@gU(@84eDf-PZBg<VO3YaAAd05)LJ+QS3
fQ>f^5LXW_V(@C[:\)0<9b,[387-IK2c:/#aF;?C(1N),O./+F_:Of<3#M)UBRPV
G4]LOP2@D13NQIRD<W(eP-LeFC+?f4][@L>MR-W.<:X9;.2-QLB>]#Ea]eUSReY=
&^_6J6#)7=(0d,7C4+f/7REDU=H5))a/2MQD^>O\9gY)9#>@e3aZT0N1G&1PA7bK
(CEUHVR/Jf1;B&gYU(V][cC5_cL5VIOg^5VD^TdF;f1BT,GTDN(=YeQOL+b/EY@1
ge:Ed&Jf/g?9^a&&O5/W<ZQ)\X/89;()+GZN?M;Ka@2C3S1PgJ^R;g>1L\>Z?bNH
JA-L/DO1GOVO[=FPGWB<?>0Q5ERB+LH<2<FCJQZ#G^]124TVZ;5+KOGJVIZQO778
Tg[2+26ARA?MC?8X8^N2Q2JS\]fWR3^bFQBe0C05aH[.8Ng]&;@_[H_;K1f.ER1;
b^-EbQI^efgP52Jgg[\DJO^fBK]@B<;I1Ec]:ggAb)7,gcF0S]f]9E3X:UP7GX#>
&_PCT3RIJbA]1JUG4OfD[3O^O-8XYY(2\-Q_+HCY]gY:W:S+EC/2aA_ZgL\gTO39
eL-)[C..]N<f::<O\B(87_W5M)@ZI&012:,bCL<afQf[\]#72J<GC020<bK]489f
D1IM.-7(2aAc10@O]T(G_H,Qc0>?:49A/]89M+f/SBdM4Y4VE(O09\2:3cH_T,S=
=N=W;P.ZYP/+,:+SX[I_#1LP#.;SD0P?7c<eO4Pa3g+c4@V5:=.JY6>1PCIU@cX6
(/_^(5>^E[M]KY.Yg&AWcU-8eE-+IaD#VASV,g)d@A_/I_HMD[bC2PL5Wb6+)<Ra
TA076EY5+U(K\^[e<[SDOA-56=@SeG2RKb0>T[.U[f>9Yb2QJ7VQJ,SQ(QX2]@8L
/2_P>KCV]&:gD=5^YXH5H/#eYJK.TXV;gVT&ZB-aA,);?1Ic&d4:],FL][Q2ZAg;
P;Y\GS]\^=BP:P&;;8&LO^Gd?HHK+#/;#RG,L(cK1]\][2a;Q-Lb)dL2gUdgB/W@
7A<6@b4E6;;.a[L24Y]ZV+Q:KZ4RJ7;fE;TOa4W\eX/HK7XP^c?+,T9PZfaD#d\)
0OALAJMFJ4\-fK\9^2TS>KLTd0XF;c(^8YE=KUWG\FM4W7.D@f1C]Oc4^@<\RI_5
6=XU?80,VLEa[7_.3?ZF#N?#9N6PRP-H_G79-KC]U2CIWP=EWR+dXFB_WOK1U-=R
JNNUN6UK^U:XVT+^WA<F(CZ<RU6CG4UK0G>TL][@OQ]2U3eK#<b+<K[,3-ZLC0L,
BZdF@Q\@I9]KCA0?JZ3HNHLFe+@be-O?@Nb_P_AF9ZMNa^:;@)DGbF3CKLRX)#R2
V+-f:J[(=\=V>E>H30H^)R4=E>&BP6J12>^@UZH#0;:\>AbR7.Qb=6-2\9Wf1LNR
_LN&_0@42EVREAW/I6^[\dOY:8Kf<3OLMF92]Q>6E,PD\VEV8QFL?dd_[A;H@K+I
;2^4WB/5=SEBOeb&Q#f3<g0MO77W-</6S<g^#7^XM(>-W(I_[&TVP]TG8A.D\UaJ
AQb7-[_;d0V+Y>T\)K7PA[Q\4Rbd\FU_gKgU^-:;WOGU#-L&U8eM.-Gg\BP]@#D<
H4NR?7\<_gP[bZYf<&N72<F;eGZO>c?B#4KQR>>S37NEPb/PX\[7;CY7aAeX\K9;
W\c+-3-?I#GQf2Ma_H]V99G.2+/W^O1\ML7fZY#KM&HC]4404e[dS9,EMW5\+)2b
gPD)gH7@L7I)6eWP=L\PD[KB_VLBNF8/P1>b-aFQV)g8@DG-OWMf]5HWe_S#6@g2
?,e5U@MY,4SS[6d=HU#bC(a7:5+?C_-.YRAd+8=8;6ZI4,PfPRI]5QM=Ma&cXc&L
QTJ1+:b@WSVdIG,_O4.WDVTM#[/H+Te\_Tb=3J^#)Z&?^aIcA7\0<;G71WA<eeT>
Vd3b=#>7U>T90KHN2&=/b@-VFWe^NWX083_Mee-8<;NQ,WA3B/2g46[dC>G2<RN^
g<#gcZeW97?6A:N4a]N:-T(XG0dY0/A3#RKTEIA\a,,Y@/DOD;4X-?_f/32@<:P:
S4^R=NLI]&X.4B5,&eZ@BH?=U2C#^J<b7A@,V5Y-J?eOb/XbE(5J:e[gNS.,X^O0
G8@?</D_GY9]R[EB\VMKVca^&=&<BW:Q:f>Y3:N47&Y1>O<9fJ_/B@]SZ<BGMe_7
^8fPR1fc4F6+aDd2dKNKHIAd38JV7_Vc[_BNC[>14g0dZbQ(<b.C/eY08IU6,g2-
HK(BJJL9&O7b>JY5C=:.U8_\[4U=5,OTAb4T@I+6/ZdO8]29a.eeM>#+_J+IQUD<
3FG:>))&J]b+1\1X.eRRWX[,D#,d.9ff9&(^[NW-8#SFQRN5_UELI_gS4>].MYUg
=>SF)LEUZ[TLf7BIX;^J).efg8&&;fMd,Q-O0Idd-A^G-cF5RFec=_0TIJ,S3SVI
4>F_.D))4LbgW4F(M>(VJ=S7K+G6<>f.bf<3K.TAV)bZd:L+_Z8TOcXGc)+e@HT4
?CFDFO=FDdB1_N44#C4UM^_@-d\@1K2+QSG)M,BHgLK=K]3FWVA&(M)A+UD)aUZd
1)a[F\]D47J;2Eg2/7()<=C.FJ6aG6SY#g#^7Y=KJ90/C_9Z\XT.R-FV/L]_cI,0
<@)1@d4P9OF<;aBX9[/TX>1UV4,SR:L7&Od&S^cS14f??6.1H\OYGX#JHU<f8L+L
/LFCVUG2_::#T>a:<>@0C:Q0ab<UeNUO86bZO[/G4?&:U1]/ICAM)@Y,ZYF@ESdd
:MXcC2]\Ce-CL9>EX+6SXX[2DPIU?WQ57=,P(a\[,^4F/]BIe#05cN_;[Gbf0623
.9EYF_b@a.@XMa\/71QcEc4N8SAHaF^\W/\fZ71[B@<@KI.cO;?.c44R+]L7?:8)
>f6gDb)C;L4L0M)eBCB>cZN=+U7M_=.Z05<TgC6?DaO(+TP/YcVWB[@MPdN&A\^#
TQbS[4;)HEG.^+M69XV03D[A3A;;HXP8W[Mc=J^?bBAc&2SK;@R2_E=RJ.\R9TFR
M?LaZL>bRTDVPgS,R^\F4-G_e@1U/;Y>).>G@7FK/HHVCIbCX23.K3ec/IQKH9De
K&2/=>)CG8[-bD-FK8a9baf+]DT(,#G0^2_d3E7J^W&CZ#_a[JgXNPU@d>,I)acP
[KZLL9X+F?fOH(V8I)44M4b_OZWVcBPUWXb+IfJ3,U-//Z)#S3#5:Qa.VW9YU\/3
2BTfQ1PJ59&(^c+-4SCJCO-H4.K9)WCaKTN40H#57De3?:SUO:42ec0=K00g0,L1
dc_)V^@=5GcXE3ECdEJ,-5AfD/K#4[\<+V<0f3?KKbgP)Wd?HYdYS7SQ^fV,AU9)
3\Tb:/I9]8-VN7PB_g<.>O9c6(ZVKUb2V>XX8fW?8AB;L+YEDU/G5RVcEXU&gM@b
6P822B&=<N]\)Ha^3K6d23c)eQ_aOX7g##H:QGBG1c4)\@A,LT&80IQ2W<@;+fCP
^W]02:M.bA5-\9JL8H-^V6Q4CbK09:-TJYRXLR1EG2K#YA;)DWIAR1[+QY4fW/7@
VL1<>0Z+Dc3=66NGc-&U?3HC#C4bfJP>+<PIN-080KJ6ae0VWTPa;6=<Ab\b-F8;
+\7RX5(.OR=9EYB+R@d.L,95]N]d\fC&3#BO\Z<)8+.[;NTAUHCTVPD2LX=fN(&.
25C)>2fK,=F=+.=]1O_HCc@gX&YH]5,I+1:&ce-6LU;:WNF_A4_PJC7.14(2SE)g
_:=aJO1YbGD/Bb02M^d=a\cbL;=GG,dRI>A)>:5_VW-BHbTfK5QMMF6KDc3U\g4c
^BQ]YPAN-f1eM?<P<?4CHX_cV;K6L&-J-CA+^Y8U:#HF&.8(XH1O^VV(MW_E31Y+
&6JC[C3L-?[LCb5)&?9?)?;#IMHY[&CB7M2HgbE<B.#MXKT^;10&14)0N,,>P[C\
UL752R6eM@1<HREAK#^>(e>SaEfb732#X8)CM@]dEK8,&,TYf43.BabRT8a.F_KX
J@;.JAH\K-#A0H3f_6Jf>V8WIUCT@@dL.2[KBTA^]F64R6[]:b=,:=226F\X0?_K
LGDC2acd&W]0\ZPR;21CRT9UG&^F/08F-FC-S+.Be?__cc:2@HUTUa/^M\_M^a>e
e6]U&<8_#EQU\>TAgLe\DGR:D7_X(WBMa<=;G,3#ZQDA&6#O#F3\d5)L1H]^11,J
T77BMA<[\4QeAZg2]=9WY(4,VIWKA19b.@=.TeR+dO7#<XbDUIaOP^B9DCZ3R+)<
+SN.0J4H[\d7AWHeED-IM6F+?[#I9BS?0;<EADM<b1A<6V/WO]M0M<C7M<PARd6g
94g;fGE_#6:SMJZ[de[;4B/c^DLTIQ<b]?DT5VP2J8G:?C/EZ1IY5.UC?VZ3_>PT
;D[;NG<T;<T+@/:AE@+GAWW:.1NLO=(QDWebIB/gG2Y]BfG,-.IK-AU,EY[0H)E.
04/gAd9R^.3\JMR00^F>.EeF1:fY?@@#-0A:\/[Gd]gY5C.Ib>;1V0^&IV9D3&_M
gc/E8Hdba1?2Z?a.60OU#ObKPZN:_B\HD4df.U8\2)cQB#N^<H:;D9;-W\/VBP/K
EQ&/6e<#+UGF75VV86VMVEE.;.0,F?Q;b8B5P14PI+YH#SKE2[Da_>8RcW]_0]-P
XU2C6Y<\Q)PZeOUa5N8OA^5;ZM<98d]=K.b5G>aN^L5Rc(ZUJQYM?7J-SfD,UMd(
fFKA&TKC;M]BH;\_IPgdgF?YcZ_\+=>(/d&^C:\)X)9WSd5PKWH:gaR:eC1P+Jf4
QR&T_8S>>:DUa]b;aII=P?&T0TTKG8@09<AA&G(\J+F,LVB#8ALZ_(2,3/&)Oa;e
bC&L[^A>KLU]Kg:d^+3I-W\62&]IX74<F8XMa]dX\c,1/c]TY/T:#>RHZbUJ/X?(
((:U(W<I6Y9fVQHB,XR2W4B8>bdI/GBc2LFMf/J<<GL02(b4Q97,,IRQ@EGMMcM#
<#R=T^ce81A[=W]EHY(L0S=;B1/:HFH#DU5Ja?7X21=<6C.BJaL?/^S]3=B3<JY=
dDb6dSDPXL];-d[.YXMSg<TF>0dXCJ5a\gA-Yd&ffR-a/8e+.,6AE)],MFK_03Y-
R,Cb]F[D_>;GWTBN^&DI+603=2J;F,8gNEK8EJ/(YWF^G:((D)+^[SIC0R&.fgeW
^#V3<dV0@c/[[H+L7@I:bNPFZbP61b_-fD\?bY]f#QL9a6.C2,BceKI#S0Q.NB95
)UfPd)&.0NA=\fHG5[5(L_c?.+aY_MWfS4:ZT?/PJLHaI9\U;X4^],IDS?M8<<>4
0aOU^^RN1E5e7NM1\\Nd2.X]+FB1RHQ/+=S0A@,@67:W+ZS3.7eAH0dW)D02H)&+
=7Cb.QOEeVJ9C#ZT?<+.Q#L,HJFYNP69g\M:FG]A1\UY5Kf3?EB3U@Z98GDVa/W,
W@-,)@C0Y(JWZ^\0-SV_(HKCHP0SY[JT[AT&&Bf9LH(C;cd[6SdY2;4(342fARaQ
1^OMNRLH]IOI[1M1J(JP.OZUZ,RI-(dMAeN6BJTd@RIaJJR<+D,_M6We?f.CXX./
84D^;Q,4&R9S;F]f,50S[0F_#EULHFHf\)b\>=M\V(_40]_DcFCS66WDX+F?Pf#X
RF^94OPc&DbY5XD5],@G2CM,a4O);GS>UaGOEX4cKWQT,^;F,CM]3L/#@G@9Jc);
3MRW.d+SJb,[N[6HBO[g]W)(/JI\8B4A=P;eO)@6Bb5(PeRXg./WL\PBZMEIb+d+
FR=-d[UCe/7+0IE>36U+>;^:aLXJUW.3?b@8bEZd<+(H)AJ@^0gFe6AG>H^b&?b:
_?;dUOZT@df(ac2C:PZ/7PY)J..HI4VH/a<3FaL87\N\3/@b<fT()NR/&4IWTH)#
We-8BeT#-5UA5=1W:A.PIWcf=E27WX9JgKY436QB_X(26L?ZP:\L].ITOcaaVRE0
2]9=W)@SN;:-W(>Cf?OEFRgaPV#(L>@NYcTL]U@YHeFg:.4&RZc7.5#Qc4-eB-3?
g=/(1AP_>Ad0BdQU9f.<.;#d1T1C+c?MEKW8?fb@6OdQ.#F3LZA#OV)RWDScB\H1
<4cR(#DR@K]g=:[9INV2(;XKBF8^3beD(I=U>-HOOWN&1fU#ON?eG0J/5-NZVJQT
eOIg:N9U[L3&^#A5ZW-YbO6]8:OOcUL_Z.S/602fB_#Mg@g^LAcgNDNQf=_1:ZDe
CU^0eCOO]aHQ^P?M()PJ_g_]Zf9DQFHLW;K4+#(.@=ARC4N1HNT5M(YJLDd_H&1;
_.TgVUT;AXU(d]CQ./G]@V((8TLX=OXTPbR3=NTd<P@]B/PgbXSK/d(OW9\Pc-EO
:dAfce\d]^]ZKf?LC;0TQLD^c,#g+E7I[B9),ZZ]Mbc.0]3Z,:S??H^G=DQ;+,DH
dRJLACFVeKUTM)C?X)0=-)b[PQ2NF(<aJ_5-g#(/D/V]C(T\++LFb&]<[8>gV=CE
beIC,6P##UgIAO<+_(<e<VfFS./[52\G#gL[\b34LH\9:E<<-9NZ>RF;#2a3SY>W
9HP>O=1)VGBcdGdXb(KK0:Q0B/a(af_B^=X=c6NWJK,M3Z0;#CT&XGVYC1daK#=^
FU#L.((<98L-5W,^]+ZUg4KY;WPU58WF@IgEZ>J,:e5ZS)X+P@b-4=KQJ&bTQd@_
JOK=[9Ba3Ff;_M]-3Kf8:E,Va0Z:7e0&M?J/@G(JV(2O<6;E&USG;deY^ONLADaP
X.@NJ^QU^YVdW^22J\:Q>8CX3B((<;BBb+K3NBDSX.82DX<B#WYHQ3b)^WE&?:Z.
F]g_7JQe3URQe-GI,Sdb\A,^3WPMBd(C](8=>4K)Md2V?;HcYP2d(ffJ/4D90:)R
N;eLK6Z;[7\3M).2L_5?;T?d?SC+8^_:bGc:)1IR+?C?,Mc?@Zc7K\HN,^0CCUW^
\PX4MFT#Y_/b\+JOF++=+7I6+W(9Oga-Mb)9KB7JQ]KDg7\KIM:<G85:)@X&gHX=
?</Ac=<dU.HW3;TH;2F23)PWg?ZT2@]]]+\D@+a:d7A-?\bL77I1-SJ3IW;JR;;d
3R694@8WUZRfLcTLeTXIXLKF/]#&/L&-[1V:ea+C3R62(JfK3GQA<YEY@<#9/MG<
MS(H>?[N#E?fPL513C4@6cZ^fCW?QA0K4(9;)+:,dC:G-_]9,d[+QDc#HUOD2J8@
7)560e=@NZ#;K.@RVBa-/;c;fT8<?)e>Db0338eA+:HF3K)VbPS#/+#\X0_YOKSA
]VBJ&37R8\4MH8QE0&K2/Ga,\[;KT[:c^[UR1K)G?C&&<9E(V_C?<@ZW<;U_YOeg
9e^HI=JF&9QA=Q(TM6<?/9VdMQ_HZQ4/Z\PQ6WO[B<b5]HX=Q-WRHXf8;[d2O9.a
NVJB8eYEbCM/79PaL2XZRZ\6,+T6cA;d/F(eN6YK;g)D#??4]^68RICS-880Z2H7
Xg)g10]Cb&3d6^0ZQ-?/R0]>WYX87I;H,K6>F4>=eaf11g=EWM17@T3PMCd?Q>AL
HRV;+&\VR=/6OYT64?A2R[W@[NR@9M,9RANTMY-1a3KVA?;LQ2b]c9b4N,^SJLR@
aAJgEO2g,Q+BJ<4]31=D6/H+0H#+PE7/@1.Q(GaY9@+<_2aIT3H2MONT7MMaJXHS
IU7YR+:92UI&gI2;E)J>_<;[?8eY,5-X=WPfFB-3Af+d(?VP@1PQ_@(52<^70>WB
7EPe_[+)WHTOMG9=KLL3K]HIEWD[@X#KK.]SD[OYO)\17X+3e0AF2DVb#?44O))9
=MWA</MIGE,A4XJ<))17H&WcNS>QOV>-0=B1Gf\-/R#(V?c?G0BO_UZRXVL>)P<a
;X09)UbY:.2_4QIbZ2,=F,3>&#_=OT5.d7K=XTeO5U=X>CKd_)3&34X42/,FDRZ/
(Q+TUTb@=-+G6RfS:YW#UT_cHH/2W/-F>V][@d2RHb4ZI^JC9((508:2L<A,gf)C
@aWN[O+[fMS2>Z]d#eeAaJ4cc6O_L:7HN,FT^FEXXK=@RaA@&7(053X0UXJG4/]Y
7PHB.9A=46U4]:2XF8Q+=d:Z65^<Of;fR<OYfDU.C+_V3Z),=)QBc#.a_?cbcHd_
[(SAK\Y1-g18IWeIB>YGJ[RM0-\dg9AS0M9K2@I6<8^]0N-VgWGS7)B7ELH9<HAS
(4#X>I:2F.e:I?B&/D2QC1)WTA?0^KR:PdP.VK339<ULS8OY;<BY47+IP0:)X,4&
c_H[SOEfgbJ<Z8@^YNTAc1:P<SZMI0ZL3EB+&5MN+N^\T(Cf_O?@af6G@B].BQRA
D(de6;V0/deV\aG&M,@I\&NFI,-6EOe]aY(7d17_;bJH@7.Z5<ZH#Xa7^9Fa470<
IBM_L6#O>4)X:J/agZ/2(S(/YF@2C:OVP>EQV]U4-WU99Q+-UTUKDA2\#d\AE2eB
JaT+V;_,8f4Yb@3+@@HSX9QI0QN(K]Xc\3@(I\^.XQ;2b4XOGT6G-gLF@RZF\=\M
4?/\L(B,J0&1:Zf^O1&<R0MG(:aH)3ATFZ;gH(/Ca?/PFAYGR6:&;(_CeU3D<c-E
4)ZPZJH3fH?A)a3YR0=f3S@9[.;d>f\3].;7QKMK9=K/#@Mb2:S=^H?^V[EEZU/Z
#HA?PTd4INZNM3/YD0,Q#;<(FHIaWXLbDIA)BGM36\9R8^X\dX[5T^+AS&8(R;T0
U/E+-@3^YYH<I12CaO>BL?[L3<c/PbFR<D<)Z#:e9I+VaX?<AM4)dP(P-4g=)SdM
2f2()cF25b=I+])5#T#P402\D:E?F:cSA[_7]O[TW1LT3X&++AU24\LTDB5A0A3+
^1c.)eS[0fG^2IAcC+e\(8eFCJIFCG4d(?T3\B9FR/_b-2^K\cS=?OYCNGdC3JKH
GL^2,[PSd>\9FS^Z=DcH_#EOEbbQ4ZWBa:-X7F7a\J?D#F^B9CA)>BJ2YH=,4-U.
<1f?(TM8c42O4KIA#Le;]9DHT-(SIb,O\=dKK\E^=Da?\ZPO,)bL1H96[0G46?3;
?Q\YHK>HLI102+EG3)PH0W)/ffN-WSSMc^2GF[WdCEeLR>6?;fg>_(T0]K.VOU6T
J[LaE&Vb;(]G:8>\L:7YVN1+aV@g\\NfPRX;-\+,P76+1Ndg6.L.9BP-@ZP/=P\L
<?;GM6B\I4C-c0gK/#570^=G369-A/eW,#=PRbd(b)N:1^[Cbg<8C2W/9HN)]EX2
UeU?REKXHfg[T0I\0cY8_Ka2R4cY)NQ74>-]d5JY(f9;b<;V2V^fVNR9b4TI:dBP
+Z]YXT[[eJf.-:.&EL0>E\EOQ:K[LV92:42W)FeC.Ve?0L,5@2.PX9UX;9Xb3DK-
F^b.EA:e55L:217<F2D@;P,_/c5=N,@E(b:-+>^9D9:Z.9&MYF-e#A\fIAHG0D>(
0?7,_JM56XM,begT7,gaD?S.d(YC<]a#AT&0R_07#f2B6Q/FE#6F)(]OQ4#9Z:/b
-:WgL8_W8>=A-,5YVcB([/4J@Mb]#HF-?BZE-9>4?53B1RU14gPaRG=UDOM7GNab
Gc00=ZM>Bad>94^;1->RZ76SN(TZ#)T9=Ef+_S2/=DH.(b[0Bd3#/;8CTG_CM_>^
,gK\^=HPFQ&\PG1Fg^f,U?de[M=0Y=8Hd+M\JZ:R6@cE:#/\#K(T@cHKa_Sbg/Od
+fFROg2YgW=[C=8D=7.cEa>\&B7Kb3(f><SMMV.S##UJ?=Q4+(?[K_<0bHH+OWHH
1/5)&FK<YX.&90b2+,LJXN#C;K]+&f:=Z+QcTHR66WK9S+[Xc?4@61V3eNfTdb\b
=f)=9;4_S#3S.JB,-5Z-YE^<2[XI[[BPT\e6P3DL0B\1DI6O434[?,7R#fg63VG:
BMW[dP6LCH=)?Eg\=M]dHXHc[_(5.Sad06^5+13+cgfW]D:MSL0IY@T=NY6EXGf:
HV>1_MI/3RWVVR7-V458)a7)9VL[V+[Xc1YUK;#P-2;;N43^ZF\<03I_LZ^TdP#Q
10VV;D7a9?/Z26fKf8ZdSLC-FD:RbPHLVc8ECg4PVV6;]9(N+PL+DD;SO(FG[^1#
QC(X6cg.=3YCCgQBc:_EP^eJ--03A5=QfCgCB+LZLR8,&GNg?PPc#fS&5D]=<XM5
==H/3<M?I_?VK:_&I7MQ./GPQ9OaJ]^S<aWJ31LE8X62^fD;(N<4.O9/SLFd#55e
4P821e8AO2E;^/Y&LF3Y7QbQc]6+G0I_NWUEXZLe-,5HZP@@6\<A1;&7PLG]KQaV
CR^_Ib0L@-b7XRQ[-R9DdR^^&EEB2.JUJZ:?eL/-.[OR6PE>MC?9,N)5I;W?GS._
>L2+ITAQa;,LaS@A,Z#WXHf7[f=Q8IgP20FaXaQ.>^3af40;23_2KBNF7P@&P3=e
ZCJc>bHfPS.MT4COgCV:[PDVT-R9;LeX^5Cf;I;0Z#U5OFH#b9RQe6?C[((WLKB@
?0[MR1#T-6c=)W@.#M7QWX..7;f-OXRd=RH2VY?6fL:/)HLGRN4F^]8@1SWGMPKM
67g)EF6O=^A>f\fTIS7G23G9[IN]GT?T(&SCR8.\NaeJBVELPV8;ZKT>^EYI&Y]Z
Ec@:?1R#bIGA)J+?.FE@@9f;&;2=))2cPVXK#;dCJH)P-4gYZC:fUI9JbE:9B5@Q
@K@L>5OL1;(^ZY+dKJb;gbHM/FD8geHY#d&e[1=9WIQ=6U,2f^[]31A1Z\>N5D]J
US.)3Z3TO\MC=U#RVJ7@I^]Z(8CSOeVF;ECbW73bg9(DPXW+IIGd0\TLQH/6BN7V
@C+@1Fe.S/MJLY30+7>;gB8@.DgBZL?LDb^?eaaI:THML2J7cQ&BOFJ-<3<d7dg,
V1S7cPIHe[:fcfd;<.+G^OB4bgE7,^NFX)V&R,H76Ge1[&)&[ZJHSM5@a^_d]aG0
7;^e+dTO3D4CKM<E8I>J&\C/6X,FU;T=gb)BbJAd6BIgTZB4S\dBMUGA=V]G+\A-
T2?@6XCH<.3X+C3]&3&(2_Kd6L:?2O<5CaA^.ZU1#VeffSDOF];<^#YL^H#Uc63T
X+U:.D_NEFa>;=4a_D(I([(H<NTf_.RR+KC/TcD<]5[0L0W>A=3>N_Y0Y.9\d2.5
IK.:V2/Ca@_MJLK_Z^&S;gN6T(+5LbPT,J3gX:,M-]d[H6W[/bDC-#8ACW6NX/8/
)-g[gEC4OTf)V[]b?3L8:DT7#7fZBMJ2<ZP9eaB]d0,e4;1B5?)&Q_+7AMY)X<GT
I<.X?eG=M4C:@e&g#/I3[7E)-?fZ-?[),e-fA(;+aLc9?>4.(OD.;Ma==b-S=KGc
9Ve-OQ6U\3\eDeH=)8352FKb;N.Z+:>VdQW/&O702BPPUAY/dCM)=J795V2SfKYF
^N8@:fOQ=-1_76OE_+-U&0P]+/aG5eZN:&(>_55U6)RN/:YMIL.J8])M<2VeQ@K0
5/\_LT-A<LfXA8@)5^S5^,249YO\W[X&gTdNdCNeJ.e;AF1[Y@b=JRZY9N8O#=]T
<.4M],5E:@;6KD)R_FE.DdfaU^DT4<1gVW_57(Ua^7))_DK_4A1FB=f#I\X\Ib((
g2/CV3WTMCaVYW-cY_.MH6d<)07SW#W_<Jc?RB64F_F@U/:X1>RPdM0,8#FFM[TG
@RaFJ6Pe],c<D_O0E#cSF/:U<L=@_Qe/Q_4+?)JYAT@]605E_=\0D?I^Q[P63VfJ
(@9L^^#YVS8CHe/,G]4^^be&8UOK-JS;P>MS<U]^7L>J<\<;(^a4L6D#6YL-/H8M
7J8FJ;a?YIU7_Y>3<3I];2_?50)=]Z5(SCFf@DY&9##9/8+g8IFJ@@Z)>4/,^P[]
U^E]Idd(;Z_9@W[Y?BBU4#gEeL,/O[GaD\76fK/cW6V0a3U_^.7H0)F\[G+G;bcS
Hg2-##Wc7RC0D#3MI)5EEKXH-MKMeb2fD8fJ^Z=@03Te[R(9&2I)+[GPE[;L@#):
:cX7cH9OTCC-^GZBLH?]R7B4,Y/BIVX3<</7X=D+K&QW8+=D_46eKT0?0RJK)Wdc
>U_):A^_<9I(aNMLPg(PX_R&d^([Oc]DGfD:?Q2>;(,ZZM4P(XZbF.gWdNT?]&ae
4g</1[96dTFL39^R(W#P=WaAfYH59-<eF,+4cg&e<J4=.EdYc1L:7I/>PP:2=B:A
A7gW7YU82U[b;?77VTYALV_c7K2&;D]<MZ,=B.,T@-AD0]KV^f>Gd>;A7MW>Yd;[
F>+2E#;FL_=>aMH68Yed=6=T.9B[93<gV[(.(]N.N(^UBbM1Vbd1C,G5b@XJ;.?:
M^R&BbR_]d3C#5&T&\TUZN:Vc@JO0P4FBX3;9T6-@=OF<+dM/.C0gS(KaGeC?aX:
fFIR]R)Q>c2SP.C/TIZ<)^^f;<X)QW]P6Sc[8cU.I,)(2-2bIO\V+F>_L5YFM-U[
H=?X,fKGUcGb@PbOA<KH)>A[]aA87B9QH5.14C0),&E)R_XgSN(-VE)O7.,6DFCM
e&a(:^Q/g/6Z7DF15\:aF\Z2O4,U2-3T7KBRaXW]<1L<\SfW<3><H3W1Ua0c8gSV
]3=c,W=fAZL46ZL#Z(Q@1GE^5Q>X0:KUKU::DI;b5BNHS;W87<W#^C1C71/.T9aE
GfBcXgJegegagBB=cbP)8[SL7@FHLY,,fK388+ed<[/>B6TU?(NS?)EIM:RL/O4b
@#T;G2,=G3LI8?dMf@U@G5X;8FK2B5PD[PQL^La=2e<]O<bf=9I\2MX3J0GFSKg<
A#IRCV6YH^2N^1C[30[M<J>1INJPd[](F7G::?=XF8_b<ZE?2c4YSMf=U1/aTVMH
.Fff5#H+70Gbd/DNFHKTe/.2[^=+B.2M.J7/NA0OF&RId_<S#BJ2)Pb[PdCJR-9d
<K]D.b_e+_81^17IE3[0U0[d?#4--eSd^VB)O#<61>E=>c,SAR54POG#_/JW:UGc
F7JB0]2=.Nd<31129[;.B(I(M_YZ00G<VDZ/H8S>[HBaX3THOEaDE9CEADA-95#U
P/W&Pdcg#B8.XT+F,,ZZ59QP^a+7T4.4QdZ#>J]4SOVgeEZB)A)66,a?ULebcRId
)Cd^]Fg\a[FKV55HK<6N5M=E:BU.B3=QVW(TF0\)[M6Eg@83,(@8O_^5G)Q2KWaf
7L</M)<ALeG&W5ER)51G03-)_O\Xe@R>M5BB)1N0H)SJbBaI_D]?,;d6Ff2K2^VG
(?96()#EOG7VVT+S,f4NH=S#A]Ce04;,XI01Q+2&A;+FLEE#F(_8eaYHdd-8gC/W
Z/b\HNZCeA+K^Pb50L<#V+S[SA3&ZbV;2c^B;0#[IKb((a<AND;4\(2bUXd\8XI?
CSE.(0F3[M2g.<T:+K^TESX3VF#L(f?KCH(^EOEXNb4J]U^;b6Xc:/PA@/=I93KX
_Z;QM[7[VLHaa5&X=]cCc/X=?@C97K:;^W97=Lac#BJ0=Y=C:&VCH1g8WZRIK._g
&98IS3NI4fFIWHK41]_7YSb?ZRC=>SZ#?@OQ4&M[-EdJ&J_QMJ]UD,Md)-I/#a#5
D:A1.PKF>2;8H8_U@NcAB9A]74CNOQH\]HO7eKIF=X8Df0?6VDU?2/E+(.RCU7DV
bZc[9=d^OQ]&/>CKA2=&Ib>(M<D?A^G14AQ,53VbgDV@E(+JEZ93#T^>8.D7f,JV
AVeL-JG2<0CYJMEb;TQ33Sb)G0XS,SA.<1\X?/8)?N9&+C]A>U5ASKDFK<PeOYTa
MG.(13-Y&G#T^dTU6P/FJA1]2WVDE)PU>XVeZ@J38J/A.7O1>@+#2<UB,HZ@91eU
3Q_@\cbIA0<XbXTYSJ_H^^.DJX^>4d8I2Y8MS=&)BdaOAMTZD(4IMdD@dNc=d0K/
M+(/3fM,VOe&(OFS.>N_L[+YZK4?@gb)JT@XH9GZ<-^,X<;CF6Q->I112LB?b0\f
Kc/dK/AV8LD:P2V/[f^&<d3&/Q&N/&@g4_?VZ0Q=bBD(P])acS/N&J?Vf.f(ELK#
&LN-^?/=]1]eIW,V3&#&Y/\XI6B)BfRFeVCED)8(dPfS5).OST&J8-,H/(BMgNJ0
B2<6S:H^DSQXYS)\(US#^RcZB2ZJ5.S7]6?2E4@(IWFV_2c/0K[dQ[N5,1#C(Na?
5XH6[KaLQX9,Kb4AO()ORFV@6gJ#RfB3)4#FECbWcO/+;I2NI2VB0?H>L2g>-U4+
V7G+2RHO:-WA]<6ZB[dGQ,9Td\2aJQ/W]/>?#<Y6VH.Y1D;DK/2bATF(PdYA#LS:
:8<I2TADFT5AfZPE1K1b5f74NE;A-/@)Y]/;WMXg2,^&EJDfgCSRE)d+PY&3^eTT
bKHJQ_0.DLVcC1PXP#B/M[PVDMM>(CRE4.Da+=;O876WJ=PM&:9Q0<V=[aA&3Z8)
YBZ=M?&g[78=#+_E@ZU6F0(ObLS\4d6(7?2S<9E,5J;SJc4QdB598>47_AdSN#ZQ
557.A6K_bc[]K[P1#8MEZZ+]B8[Y_8e#^T4Pb,\05G4#bPR4-fGH6X;aB0R;.3D,
5/K+]^ZNg7Q6ZCI5g#9^R]?b,R1MEd2T4Q.A78OG9f?7aCN4(0Ab,6H:UbT[:OFT
-fH3,FCZ@#0(61,c)CSBYL118_?DF-#GIH@CeI#8eH=)L?bg=gG(?M+P)=cA&b+(
].<\RN55@5:82S1_A1fc:I_4TZ@:52/_F5C0ePgL6S,QWg[g6^R61N&.SNZ;TKaM
?8Nc0^DDU53LU8(c(C.5GNLf6+G)I>V.;[f7DBNYRP^V.5BIPPBDY?KEHR[HfNFV
OUWFM/\Qf6C@#^POPR:@S_613#MZBW1eLSZdMUOR\@4/QRT;&?[+)&3N)>9O@NdX
7:b2WSB9aSP>+W]J+a/eQFeH5c#-=+=1H&HfXL(HGK/=(Q3.0(NDPaNMIN<FGWNL
T#U3/+Sdg2;(?MT#]@LR)g1H<XKH:CSBQ5[W.I3Z3N.ZBB#gRg6TSc2QA7a.HAWU
C7).\(?:C7&N9K2E+-R^Z^=N\5.E2f;dO,).25)C.;V\Q257BgRb.L[?#V2TeUC?
YFQ6MA@\+HSK?]4R08F@;FU:fMeLZVJ\VPU_38[b5S.B.5E^I2\dXL3?\CA@/+9O
N7NULeNUW335A8MJ/40/86([a8<2F/3&\F9,H_eDJ5UbbZY&a,FJKK&L3bbC\S67
OS)-P>CUGI(@;J^411bD^cMC1SC#97H2L9E,dK.)H0e<?UAMIM2E.1F:8fa#6<\\
UcZW3::g?Ac6@(e_gUI<O:<K/)06[@-ELaQPC&:<ZB9AR,0C/)D1[+LFZ+DUK)6I
2EFG+Xb(_?5PC)X</Wf-#F=b08H0B,e0:X8:E(L_I;)d:EGZD7YT/](XG&SA\N/\
XC<?QEGM5UII<QDd7TARM0V1=EK:P59)3c\;,)VV@4B5\9<FgIDVT,8RC&TJ,Je6
?\06Ve8)-V6X5AOJJT68AV2(MCR=+I_ddJ9J6FX@7LN]WJATM(XTW&^:7,<)E;:g
H[?=^[O&&fW)OgYWG[cTGaG9+)7N2W\bZ=ZCTgYGM1/KbVE=:0?2J&(Xfb0W]aTD
11ebGC]2)B^B8f1VCUX.O/0RN5,0Qb+c4]HgR-Va&QR[fCdP6KbfM)e(+1SURW?e
=0>5/A&NUEU+@O](1(-+@KD+ebe7cKJIf5?L\/1/U>X-1IE9/]]3JHN(1-d<d=Ug
<c-L2?(KYJD,NQ>@cF\dfZ.AHbGaTR8N:3V7;??[O?S_C5IVQP38USaa#fISYBQ=
a)7fUZ1G;E=ED2P&XI7N?V.JAYgCA<;aQ0;@K=c@Gbe/SU]8ABRA[UVgb/&b]-/V
>b^X-JdSVFd[Qd07&;6#DfB-&(c70:@eAZ>NC3>6OIL.(J8<Hb^aQNeONb0U7?1D
K.H3aXaR0b.)\,;,g?f(Ke+8&Q]Tba;O5<>KcE]N\.E(f;X(D\VP1T(<K3#\R)\L
K(?EWSgCWf1[;gLa_A>.?a,:Lb>dP=Pe<BU?YL:.e>QW_e/N5fETQ3XI?LCD\5T[
ZGIVYVTB5fdO7eTMN-cQ01c:\)VfTC/<CUOe,N;YeD#PP/-SE(2+=B5MN99[,>&:
;A-WUJ/=0d,I7+ge9Yc425?M]A#Ve;MY=TCJSg&YGZSYR>-d@^c1LZgIc+dSA3PT
H:fMWg3LF78C.3?f7HM/ZHEDdCAKF34NdPe\IB@=IA9E^UA6O@5+TaQSO)4)08=:
G#8+04SOPN^)]U[/Y(-7[2^@YYQ7S_OaTQ8d@(VVc_5T:7[33Wc]4F?=0]MMHEQ3
=Y_/9(HHf]VWZ-2R@F-b=[bRAE.(\V#=SaDR9V]A^<AeR+2RRE&ZdK-SVfYIS7U-
\A\4^Ef(6F2SIc[)^HT2B@VO(gg7G:Z?TR;TI:Q+#A1bfX=K9#a1gUc[b.]1(?Kc
X=#K#>#dR@d^=<H4Z7gDeJ.aBd<5c1Tb6-U8d>SB>(+TK^TB],#MfK:8fSNS6MVX
[BEAVd7(HSEA5c:^/CCJ5c\PJ\4L8MK8bV-_4Q(Zf=1,cF\S?HO<6X._3;b0d;.B
(_0(e>/.)&[?G1&DG[:XQ64)b4[,)B5^^<5f3Z#CbVBcV5)Q@4U#NR1c3Y,f;GX(
XW@[P5:I7-M6gC:W5d#V4D]S?[S.4KB,3D?N[/f]M(W3:>+;,2g=J1&eJV9Y4X^O
->L)eZCN2>\OdM5DA^[(4^YQ;4CE5Tg4#K.SGe5Zc8c0QRHcGc9HcABPFK4d70fR
V0)ba/.EH4aCOT^PM?F-]<ZULb2(HY9HV=IPdNg4EJ9WA_82\EK/)eVYL46RWDdU
T_e4RS6fY8dL&&I9EBgBRI0\Qa0eZaJ&P-E]^c&&3RP;VPXO0I@=d+2MD\g3Y]QH
b82@V]PUK+W,VGTPX-WJ>aA:#Z(O).JFg8\cMde.IVg^?40W[U0J63+@d^c69<E>
)X.\(#YM)255dII/RT@Ge58\9/-,&9\Ya8@MIaBD^0VN8/ZQ55@V6C((91X<aMg/
cM:#EZ:8YU8<P89HObMU.#XU3>_/aB5-a11@VZcXZ-LI4IgZ0^/3D>3;<@DEVTR7
=>NPPf3_&g)N,Z41e-XfQ[GJSYVaL]AeE1OV[[9[>Qe2K)V;29)Ya>5afa_WVgG=
<U,eA5#d9W+1+,Y^>DXWg:2N_:7V66B2@aY5@4/C42&.5::(UP\e/P?KX)c@g1&(
XQS_AE\g_PJB<G/-/B-XWC9@YN#)XW;GB;VHAO\XT9S?EF0^5DY>/78AZ81aL^Vg
3N1-fZC,#c)-WH+9HO:GU6Laf?AVH-/NcS&&a>HfReaO;<K[(+cd<dO:Kc(V@_a6
Mf>JCc7AE(8f@C?<HgT&2QC7SW-0R\3^6\c.@,:+fQ)&RE:O:4)Z2?XagE_KX@A;
(D@+5K/cIGf&d95H\4C/_EK,;B0a<874QOK5gbJAEd?=Z.L]H,YQE=fS8Og#&=N<
M2/>@WVefRV657,33g:]NMG(S1&+/f:gE.Jaa4-0>BdG9/M&05f:?7VL5@6@+1C#
&bRgAL1/^FbQI16Gc[4ILMbW>bLeXbf6YcRX_0?T?^JLUY4L7PE]MDQI0b8YHQ.J
?J=KO.?eVaX?O<Y(PBfYOGTS(@19E4IX]Ua[?.:WX#Wc[&>BE9\b+;I&P[6;)Pc(
:0&(GfbM_4HGV3H:C]YZU:@<a3XI0NO11Q80R#S?-:T<IF?SXc#EL;52QF#7FV&Q
\g(>dDOb&?H-dIBAW:3aV]OHC?MDaacdf5N]K6KfPe>LaI#:bTJg3QUf?Yb[&D&O
G]_>GGT=<?HM)2:\gF3MId1=D-EI67+<cZ:G6WB;U_LGP2?83RK)37YdVF1[WgNI
4;,d>8b1>,dKH5BA;OI(\0T0=5Yg-45R)SQ2bLYe+NL8S)5B(7dUT:PP/-dKf@S.
F\,=<0:H1].F#fCO+T\@UC8#LCP_O2R4^)2QaUgJV\KR.SQdFZ0IS]?;^6WCL])[
Lg5-K\X]CU#WXY<UOf:g9&6QZH-M;^:CA(>5Y:_R95\KI^\c=6g8BF?;8_(+Xa&?
aOa\[@#75IPE2I/#2Q0_fI?_XcL/[-675\c39#N.0T]3/A95VBVS6C^70#L]>(G.
aM3>^<gRII^9,eOS1R5+d1Y?fCPI\LNLbWVg-HWe6007/IN^HKNFZHN_Z/9:MF.\
&P6JS2MZ1Q-8-.FN>F&F]GG\_aNR=_;/SRRCcR:2YDLFZ:KaS6_QFF7;K>FWb]CZ
/ZO.1M1H3=]Y-;28cI;0NeOAM9CD&+R6,=7eIMUf\^df7Z8HUgaV_DQE_SCEcH&O
;-C3Vf0A4Y5RPZ;NNCMB]VP/:C:B@D5d=)^R7L+?[1AeT#8-C3INcWY#CD+EXI?S
Ef,KT5OQcAbPV4#FMfcL=FF8]a;CSR\K9&f2>Bd:_d3XPJbA(dHd))<+3SJ+RERI
9C\O8)98c[?^N].=c1X6K=R.bB8#EaO_X2PVG@L99/9R;>Ic1WD[FVMPF@U04NWa
70<:)X1Hg)6a6/XA&fQB&/cX;4CJMTEAX<bADGH4^7.Z64C@E=BWM3>WA)d9;&],
a5XV]]75gFG]>3F-_-aWZ=,@6]9:356EX8AE-fJ<(f<b(RX4ZbF)f=+&,3]#_NUM
WD3cZII^cBZP>1Fe9\<R/6)YQ+=&dBQL_W]Y1;d)(TF9V5=YH.FU6bC)X=GZ1)@>
02]9b3=b#BNaSe:8GCM_:Be<LV]@@X;<fR:(\S&XDNWS3gcQN1KYD]V,WQNM<6)O
P4c]T4?V2SS-&WN>Le110>aOB/)]:L1;7\4U1HdBb8:JA])\5bW^HEKbJ]1?0(TH
9/ODA^@ZeXZ>SaG<aN.+b-=I@K+/9IN4>QF=7;>0g(WL:;XM9-&KD?]K..#W5</J
F)^QOT7TIUP_9)QZJ?L.MSDIQ,Z:?O5X-F?S-dT=TH2PRE]eP^CAV5@J+@=d]0Z5
YK8(3YOdZ=:FV(HRK-LM/TMVRTbGb\;CH;a1H#fD^_[:=Qf)CKaNMVK,e/LfbSNX
TEQ(1\eebG_VD1I/9OEc3?UYAM[IES&I#QTNL8J68a7PM/4\4(^ZcR:e_E#/cQb@
0:.9>G-@>c_A4gART+2[J6^\&@bU+G7DgJ4-(&+JHWg]LW&5],2g90&#7G6P]]_V
bX6.R\4]NOO:P)WTa;fN&8I62UZW[Q@+BX2H\5dPbSfZC4(;[7.YUH1S_d+g2H0Y
Y9fHB.^S_E1G/BUb+SC8>,A>9dEa8SN0-;bQ884HGR6==&[H@]V-ALO?gb<MV_;3
X])a-L&HPZ]<8,f)@>C>L;\?[R44)dJMQ-CY:7Gg(42+U3b^@GQVCTP?;g+EUbF8
]L.Za#+:33DQE_FDgP(2g7M;W^>^)O.Jbg,\gJ?5ED185N9KW+TOM,PC1595MTe_
bc[S9>?OfIH]_F8J\e3;#_]43)[_9cI8VbGD_NeURUIU2I96V.X95VO3Z[9/0YfL
FK;WB/;TNffT/30Je,+7,PfdXF)G6=V.=H;5g]84B3;<7,58&HYJ]7)@K[6A?VVC
_dUc_PQ255=3ME+0K6G>N230]Z_KIN;F>X2=T[2Id6NS\3]<e171fSY^R6d1^0dM
;fA0.&#d#+3(aWVKLd)^-PE^Kc0W&0W2_&7S2S<be#DZZgB>Z+=@?](gd3CAT7JE
[/+8,U;/[J14O&.F-be^OVB=;R21TGWH<]H+.g-9<OBFb>HgM1dXA6MRXU4VA7L3
1<Z0]FZXZ<]?Y/[8GX=.OTVDgYUE2H#&/;<<T4ba23RPDR15-3[c2F(HHO4^A07-
,MH5f(6NbJI^J@\eVSTI4c0YgAN=AK>f-<7#@a@;LfeRfdE427N3YT+4#O^MeOSV
\>cNK>JIV6g+/33CLdF51N.5YGfH0ZWI;g]Jd(?Ce;9)G+eGT72Dc[JM24LQXQPZ
MSRI@7TaYN.f1fNS?QOQ<4#:Z(PLTHFU)Y9fGRB0L?&RUA&X-;I(]IObTGPLd9eX
]T9P18W7c6?<MGO?LR[T+PW_E7KQB-+Q@\2KBV8bHE[O7M.<]EWC&fG@)/6@gGZU
,gHAJ;[cATRQgRVDgM4)aWU&FH??2J66W?H-d#YDC,;YW#g)6ED]FN6#+1PS?F5.
geCaDHC_-#Q/6N4T5e@LX810Z+F1S5YK^5=E^[HH,B<;^J84&&TFU^7-+&.]+\TN
W4K_=RV/a8PKZc^C<,&gTK20?XV4VOVa/U]1X::Q[IF[B/U(>H.V99G^.H7b.Yg[
UH42E00fT05=b_(B\N]E3\OQTKON5gX>#T;9Z0&NPef-e:C7)2[#@)f(E73g2c[<
2RZfS(LMV6#LS]e=R+_OP1;Ig^2#\(5,4B_eXEV)\Za[WA+cg33_G].d>P&X(?K1
ePFF0OOc(RT(H/P;4@:7.&L?QKIA>EJ.;H>VSN1;]&cMHV+CR_3H7#.dM$
`endprotected

`endif // GUARD_SVT_AXI_PORT_MONITOR_DEF_COV_DATA_CALLBACK_SV
